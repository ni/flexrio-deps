<<<<<<< HEAD:flexrio_deps/PkgNiDmaRegMap.vhd
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
gjQxfoUVC1+c91Q8h6upBt6MO40asmyzYjt6VzGWHBbwm7lJ9Lhol80B+zuKYBmN
mcYXsC6GTMui+6I97KVF5Gvt4jM9DzHYcXhJYGKlSZ1LFuAbBoP70HctjPVDs1uU
K8OsbS55VyhEjKn15xiIvtXli8aGjXHeX/rfWqMfS42YUCbSyppgEsJODINwwOzz
1qRUUw2/jptV19c5D/Bb6RJm+DD1WPAcwpMfK9yt4tt5yY7aldrWUkuXKybQ3RoV
uy4U+pYfr3W/CkV2CFVLeksjTXHWQavgyk9MpfadikRr7Bbvpb8mmj9vgqfXNirU
FuwWU4CEB7Lj3xKCC5lz0AOsenn427PLgbpm5lFI7Vt8g1d76B01xjieSo9wQdsY
fy6xg7fPnBWhH93HJKW6laKa7uA5pPRIFnR8N6neQujORfa0mBLgPXva1p8X6n3F
/+uOR7CUBSJ4KycOaVs2y6PesbVc+Mc/+abM5Ivjh2XgJGj37Qvi8HySFfyPHwoo
WPADf4Ef0cA42gysrKU+GWwuP9gjduAkuSAig6wvduq4gofglrqhCENzBUIUINIC
o+mzymAtmg9Ko/NRgEPqqsY3E9e1i6Qo6DfY6J9LuZQXm1pRpxnE9atrhsZH4kt1
0bZWTNGYQoLyPNODFhj3SLHkQFax4M+lcTkhmqK2lJ3xiYTrJJMnLwoUGAXIRPOj
Kj9v7LYuadDGcgUpJ9jzYBj7ZfYLOUL7YWM5SJm7lhn4tmA3VcK+GvDBSz24MpfG
f4PhCJZ8DrEfGU5v7xN5ipIER3iQ7tOvfJBG5bUyl32B7JzdThiGHekpIPeSjuUe
g1A+cJr1k5o9HJYsZsG3taOo1C4mhKm0OIMqk/RUxPsyEx9KavytSFtfYr/oBboF
WiOsYQEmy27k2ClZnkTfsfzpO2F4b40zXoS12vf7DxNJP5iTkUGmuSenvyb7/sF+
eo0fT4R7D9RMLmd2PdevrdOMQPwVIB5IhL7tnmtgjtDHKCjOlBBP24O8ii9k/ACC
VyQTPB2eNfAceYUYdbipcU6zdaf9ehrubSxW8UC1Hd5f7CSUQmufGMYdrJ4lEm5G
kaU6Q16ed7oIM9zrWmZJHxPFiieynBGT+A/ONRlCU30htDxDA2d7llF+RSXRkUIM
KonFXSkysG5mV016JFZujiUHUXv3e+5vBFakIhwnyZYQwKvScohCxaQytdyPv+Nv
MgraL7UKXwqgACIRibVLm53JsJ2WlIyYvzMrTRzbso1d+mMGDilwVdzEZOyNVq4L
JqTDJjcsHCkNvQMLd8i3jYBiRqhO63ZyBF7ooOoicRK+Tq/afsRh9E3Ve1VDZjIx
ucli7ybR59rvIt5odT7GHyWfCyHtI8t/OEVo2GXfqurws09cHaziaL+cqDyEPGUR
51/VtiXiwSWss0XCdCeYOKm29bBzJlv56+65ql4E4hDvC2N7DVXCAxC3N7WX7V+i
9gs2YZ7dnCzKRR8t3JNQaB8daJfglY7FkPOkLF7M4qSjlHTu6LQyKPQrgB9Hub8h
fbTCWcftgFLkoUyIhkM7hjSaVUJ+xVkaG/V04pq+iD9HLNo9PM0I+19N7RWmqznG
7rifboZdc4fuOyB/aUoSVquMD+lZjKPo6juEaOm1eJhCLRHYTW4XqzjVZ5A5bvX+
H3aY13f7pbId7d7a2Yuvb2Ynz5dzhc6oAfQyCtJACIxkxcz9ZSinZN3YPKJTyS20
4DRTI4bVpbdVxNy6dIT0jA61pdiV//VNVYdIFYscUBz9x52MZ0ylwIGjncSLHPDa
zddfnpeNm8xgV/ouyE4JWZhumf23Vw+yUZ4taV+Wyld20gDlvIRmIoYw7lsTlJdc
mL7YQjWcqQR4cNvAlLtoLDJoItReMMnK+jdmrUSatayVDhNsuouQ8Y5/VOZkqUWv
rnb6ZATUsHFdSlD37LvGWtt6G9au17eX7jjWYGbUC0ZdyvpxI4tDmy3ti48/AayN
/aBxl+uPnzz7HBFHMeKzoGXaF+7Rd5gLuI03GS7Oh78P2Q9gopgIx9JPN/FVCBuG
4gLn/xUV1DVnXY/hs3Yf/Q8TEN6ixazwMCDLFL8yB47ucqKB9b2yrGLBXij2JG4i
IWFqP4s+JQ0Ckmmg7358n969/rgfXV+1P1VG5bwoUcyIRyedB50klNKVZfhRtBPB
M2shAFoCfK0+r2OuHA6Z996ZuljfvWGilLmflIBipEDPZgHoKPblnOPUW3oBD98y
pNUAx+ompypga3tUfVYqEkuiOFoEemjQ2TWahAC3bVEV0n0jz4j4LXmuVdeutJWW
N5l21cB2d0vIIDvNcITCT3k1NhNH8mJS0eq6hH/WtagDn/bA1qpDd2RgB13CXh6r
NJ3FGC1VLyqaYnqSmWdiXjGxP/2dyg8Gic4MtaHgqlCkSLhmUm4hZfOJG7zF9obv
3vf3hIWjRyZgx+bya/NKlowUy3ZH2hCLPgtbfLxEpwBvqEKYklBRs673/K4T7LG5
Qa1Bz3sMCPKmsMxiUtNPBf26y2VlnyTJCh+gZK9BbqJrw6lJmoYkpqGigjyESOYp
P7HuEmKRoA7JNshvbuMab9c/I9CFLPsP5iFtbYjn+6zT/BCACxU+hohr0rv2JT//
cFiorKuAn/idap+GiCzieK6OUdnUBPVfoOBblpJfHGrczLjsFz19BPjvy5dE8aX1
W/UJ+q6dN7asKRSoN/XEPLaf4zKHf4Nt/bEWBwVjGAwzs9KLwaUEVt27HyYhfIOq
FBGKht+4upzVIErZwB4Ftbb57xuO7IYUnCm3NbVyVhZAtUl09c1Ykp2eI4CsoV/z
4sAOHSGvRUyldNzFRxSrQur1B71o2lNhcaPpy4D7DU27jutDdlTdVhcQPv0Tz+SG
nLh5F+K9lZJO9NxzLqfqGe/t/zO8kHHVHoLhJetrGtJDPm5ybdJn8uFTu5GfazpZ
HjDTHoAvlBhhVLKmBtgHUjOv20AyxibkpbFWegFnSV8EfriuaSavq2HSSMLVT+ic
MtPyuxtUgVM25uTua1rIwTShOMAD9hkfeinq6BAGu/IBZchzRBW3dFl1eedgVGod
TIHHDK7cI2+RnN/bbWgZtMN3qDb3t+uIx+iuKMBke5zNElSB+JreyLzvkZniW6SY
jOspbdYKvzjsQ9kk3pt4G4+7cN4VnqrhLWj4YwkaNAV7J6wt9PnAqcjDGZNURiV6
jHI29x+/sL6G/8PNeFn7qg/w2LEkNZZs0/gnePNgsAmONHB8DIdlCAfw8/4To67F
dX7RNORsOkQr/0g2x4LY3aXBjTULGnfqvm6OFbYP7i8Eeks5lRQbtRkqiAK4winF
esegeIskshJISFNnpQ+Rcb16RKFzz3IexPhfuRPLkQQVkKxujo8Tnfo6VS04hJGx
LjGRwVMB96tMYBkwFtZhBESMbaGJQhKSDPtG696nt8QbtzmY2JLnszxCRCnjdQiX
LmD9VKyKohpa1Fu/V46LoA6+CXhaGcw/SCTsuYYBp/8kJMIJP05QhcTN+baEI0qA
EjCvw+3cEvcg6auA9FVYZDvgnpftHpiYzPyH9ylFNm6b6dRSZDRvYsiBcsOyjmQp
+KS9GrHG/Z/ansVxltR+dn99Ug0YtAhQdDYLHsxyuhxiA6geEbySd2I/JDCDsCl1
tnuE7gGMzu/CyUZ20kY7O3gMtiBH1VAl/wA2pvn7BswN4V2UO/KvOmcDyXezmb0t
UxREvNQTf9du2DPQrB3zDwIohaf/Mb9MtSfoHsKAbT8yHfVgW9DcjCWLFJRH20tl
ib4aWYORZjBEMm79TQwnXnT/2dne135NbtuCl3T2YB46vAtvLniaiegCTEdeJ3ej
sGVXB060JC16z9aoaZ9PrdA5B9nPWslcRqaossT/6yXGGZB4WkmeoGyrrlvOATzw
T2Y71mCCkpWp3sgC6gvp8IXnJvmN6fCA3WDwi73tqMxv9o0KcZsw707L03PRRE1l
jCqQUeCr+HJryMD5a0ex7Yh7qn2MMsz70Y5WyAg2QL4hZgO0TCkXN1KV/StvJK3M
YeFDq+YJBUM2/pdOqIpv5Cr2J5ueWKKNTwTAwMODvKEdxQ2Bb2iVG45QuVk5zntC
1wxlWkyedh+2Q7rlGyRQs8dtyn4qMK9Uu6WO0c+QPxdMtrdSCCRyfSBq41orRZ0R
bvwmgFZsiTYulaQGYegploNoI4fa2kUizwgynyf9Kwc5Q48iZ0UWWHovLMIR5vEO
673pvDYU+2M5GtbdOKQcGfPenlh2pyP7vMmcjUNs4Q9oKx335FuNfGHZNOIDyELB
Z1hkq0pdVM/cHhhUbT6slDmj6bccuGMXwdTpSjh+r+UYFJKcSls4HYxLTP0QPjCP
J+aZmvAIeIvPHv3RBoLebBkQ+8WuhnKUuFpuw4T9maWgatsBTQvP7A1LyZV3zOHk
sy9vnUwEALivicBXPPepN8PEy/qEAAAHmBBzfTQ5iGsKGIvnc8sxA0DvfxfCP5Ry
41k/b0MSbrLGAMSXacIrL5lWZgqy+cOX3+jYyJ0/ZLI3Jc9sza38G9/GQI2ctOBv
b5DjKPEHSFPUB9h//UDdJZU5iVw3gNn2IM77o/mpqN/HA8qtyau1e4Nd8rpxuzQV
CX+o2J5IImYQJ+I0Dki754w6RjZAZ3SODGH6Dfs7g8KpwpQ9co7VuKL3x1DM+eJu
v45/tMcxavIeyK6m9RMYt3rJjG8gz2OvdS23jN9Y1CsS/uCJRe3gohslS6A1yMoT
ZtBB4Xdo1zxBaQ18//jQNJSlBor+yqyTu3w8Vpgot8zhxNzI6ZWhznPiqNKZ1HZ5
68YxiEPapzWCCAKkh2Pa+PXSNLIKPhq+1BZfSqHM/UcLRY6ZPVohWkn5N7MIx59/
zxV8rm3WM+dvzfA/UDMKLhJoIfbLdR/qALOaHSvo7wN4ezl95s5Y0QpA8VU2/7q8
zS9SlykVF+sq1zkGA/Vx9ajwNoK3AX3hYjTGf3OPLgwxdnlRiRE9CIrgCS4NpoUm
shG0YmI7/iNVIBAj1j16X4qwTKOVc5rGRHvPqQs13y08Uu6Xe27pDZGrGp4U4bsb
NnnyA0syKn4Cu1GMBl0PSw4tIAXepvKUTfU6eCPwh9dl2E/BcrmPzGwQ/9yUNhyw
kap154aZsCphToIkxrQjaLwFh18EZBxMPLhHB1tm2jQACCZGwh8A2mz9JLUBJbfO
/gAMnO49MwTdC9MelmGXbiIBxqX4I/hnHOlLp1PY+F1HTWKiqnte8ZVGNLwgRNFv
h6OhyMYG1si6vEBvIiSB4oTiL1SC4Ra9PS5eZJmDD9VcsoEdW99ogXXjBZlwSZBD
k8SMny6h0hPvb1jGbj0CWNFuaW4Xcn+DuuHuuObCGW9H445GwbkT7soOW6AdunU+
Tp919E5Ol0s6A5BmKkimdFqVYhQPWMd5hTEzuefezbuIy+waQKcgZIeO24JF9fsS
hnFQUs9Grusw8fYrhtlT0doT/t6+ewbuoxu4wcVIuju8nu7OptkjFY8eyB9zumf6
NM324EEP8p4/8Rxtv5Gg9gECobCxGhUgNtj3YX1q1CRSxbePfgPzv9nL41Txs6mI
BWvDVr0HFcdXbnNeDss9qx1ingEwT5tCZArV/jfYOyUGp13Sr84VyPJOrrNqRC9A
a+uD+NL+61AGNeldguldXSka4pEoM7JKZYenOrsMWLz9eSqXjtWJ1FeI6QBmwYBN
f3ANCiNh+I+NgNlG6ru8qwGGLREabEK4aVZgcyUjVBBmn1ZvxSOMxspgd/y879S7
v0BjBVSlw6s0MGIDvyuj2FZoeZuR+UxBuhUTYlyNDgLtwqqVcV2ilwzBuvFarigF
P79z1yrXIRatfMmc2aRywdHNsV0ChioOlguSfbydElpLNKK+3+xMZSmo8YtVwi6/
mltacA7xEDoVOosU5H1TA7PC5Tw3vKZiJj/nN3dV6GcIe0qh05EuYx57miyQ1kKg
vfo8vIRS98IzqjXL+N1xQE6Gwhy8DFPXWi6Ys5U95zx3jT50Qyea+s4qmbpSlJ6D
kPQAZCaODYDbtb7HMm2vZPKSJ0gBg36GSEwkvOwa4UX5DVfnoX5dZ/5ehj7DDRDo
mVnKcuvFmqPY9bR4TOFtzfRL7fcc72DKkjC9oNQeetzmjWyG0/uaHP6kK/Rtq3GZ
/OB1Or0rnCbkhch+PVyMDqwb1QNrolgEnBzs0ZSn5hnPSgGnq4Io4hYx9K8RpQ8r
qAnXEbwVdOlq2tDv+uhA3DUV/3mCVwzkiNp7547fFWOAolVS3A5eXR1nXdBm2HZ1
msCNy/bp3brEIaaqMt5gxifN13ZhH4zXlWNyxhFslVLHp4CCPFEbsQGDhVVrlUBy
CXkOa49Rsnrj4CT6X/MD2UvFIaxQNG0WrQk4THw1ZmBkc65pEVmFFT7f8HzJj1gB
2Reakh/Jkmmy1j+G+KyqRdN+uwUTUW5oI+bRtrN5lCAEQq8z7bR5FCKRYvLRsb3u
H2Ia7rEDDR3z0vqBVkIxhHnaH+MTeX5F3UV2tuDZW/ZnErVJV3V+a8Rxci8b3ZMF
zKc2svHUKHXXhUpe0CP0B51HHtHuV6bcYw3f4Tda13iqSiOtK1VogOfJnuG4R9W0
DLU5G4zvT3T34oboO4Q/cdFsURw0OUnW680Or3o/akvvKJaMCIX2xGmQQm92MTM/
1dViNZhfRDqz+baTwkN4Cm6sv93FgiZ1KcytipsoY/cQf11gH9rDmzb/d8qG0Z5y
XDRXA6IQOYjs4o+riwat6wIdOy24L6LKrYh+R6U06C0CZbkEikQTlE6O4sRMoS3M
KSIiqcwynSV11+ll0mH43Reip7DLWRKAvdUyK0+//lu3PZOtBDuN/YHh++lnwb4d
jPKUw3G9+q6zi2PhbijhUMgbieSdQyq1PoiCJ49qnfjQ+34A9woUfvoBRBYVfjN6
o5dZzfKFcqNS2P/XQC+1LRO5R2zV2DhOXPPCsuYkOI/Ycab2giC1ZjgYtMjFeqHf
2j3IDFpp10ocBLwcTibM5iLPZa24OCpIbBja4hryNW6H1WVMOrDsC7eXuBY8X68G
D57W7PRUr93/JK642AuAF+r5PIaEvTb7LyLne2DSLAqyhJ3QHuhjAqSLxQteKikc
2nQ94WUjguwQX7hb2sxACcsS2Bj/7QiYYLb9v1K5PgI2KeCtxAU9sHCslAM5+54H
QBYBu7r9YTtyJLeUmAqvIsyFXPN8y+QovVTU78M25c/fgTXVn4sosymBhogySX57
pDqpc8vieN+NkVufuHVWmt3dfPJNSBivjwcNGZ8hzDQxvKYYCRqmbvnkxaiFQtfp
dvEPt3pALnyVfNpkhR58yUe5pFYrBelzGa+bbV7c3GBymmlWRcWRvLRdCfEsBEUS
AzkIDx399xNMLm8ZIk28BpsJ8jrNx9o6XupDgkvh1X9kS8zVkSeuEO20SqGfAObk
G6kwQhf1gVayMdPcnuSf9+UOq7Xbj9XOV82f7bEEuGPtvGHRyS17MHznarVrJiOO
aT+aPjwrYzeoPT6f8E0p9JqJMQB7Nut7HH7RfxghaICmiaaSOHQ+50bhlee6Au1Z
JZdRTa+Zqa/jBguxXgJF7FoKO6PujU40IVMblIlfT6HAHf4iYvchYFwGaMbzpR4w
nPoLEyc5asjqD4Pot//oBvVg6GrowokUDEQzn2g/NKVlxST6y0fw5cGyXKAPCDVw
OCa5zjGbj/b0twQD2lPan77NIbjxsk6NcRAgpISb3dtZRm+sLZWnuMGDoQkcOdkp
9iEs5aCAXbnOwjFCdmq1ricX/75BlLd4JQhN3BQtBTNhRecVY+EcESjO5mWFK7ui
rF5USxheYkRfaQIqBovzsJBuuzON6RWZcuONoJCtjVKh4Ag94v5DCdKnISWe8bWi
NNlcz+J9BnLovfV71gX81kOHmfn6XMldWIOrh73BQb6LdG9HKZE+VsovI0Y9YZ2z
tRTQq/sN89t/yy8yjyqtLkMtkrqaV0Ys/geQg2SScFkAf4QS3Ap5ICZLitW6qo+h
HQxL/MAdUY2CteeEsQbP3wDGhhhVoK1Rnma6mECIklvy+5Y0YdjWtcLU2TyxQ+cg
xpfTEoXTdKRAUS/CCQmyPRpFATxjAv+5LpcLhvKsejL8S3iblrMMHFLsDP7fGBQj
yGoMx7w+Ma9vtIHvra9WySgkRCOkPs+7VUeZ3sId7gcs1fVtkHY3Hy+gPC187EmD
fcQkhQJWUD5EuJX+y3nFr7RIWa6nKSNmg8TxAgnLNasVpJIt614GTzapuD/6OxLD
G/HczSGM57NhAg0+jxO1so3+vXYEKKCugZ6fUNi4u8lSEYad7eoBtt+DWQgrxfT7
xEOoBytOvt8Q2Kc1vidnSk99jbBL/umbjO9y5/aGLhTuwI7Q1P3c0skyhfcFyS8J
nUGuMpUfjl4qEav9YM/+utbfB9fopEfjK+pfUHjkiOMG3DB1r2enosZNlzV3YgRg
7c5qB0Bjkde7raQ+PI6SFV64zY9qj/je+RfqPK6qFYRsDrhOLL5VeZ0Jmk6VTsdC
37skkJlCRrbVdNTdd8SXr783EgcyaIaWKr0ILYgiNzw2LCJLd1e48bxgaiI2kGlU
7MNuyzdMANxMjXnBgQx9aaKZMks1Y/OoE+okuw7D0yoy28Vvm9QBltbYo/uAgQNT
B4XBArTkN8Fu4pFkti2WEg+gHrFRmtZvIn4uJc7G7xa+KmG1YvgVFUpGfKF7ZXMB
0lFun/HZlSjqpk4PFmhYqvq4xHIY3EnnHA4Kcct85VhbJ1437zgOQ4aqRhOn5g0/
YdYQO4q+r9zU4qv5FPvrLrnYIWM5Ghigen/wD/NVVR4KAt7TgePRmQcFB5pMUuav
VYsWJIlKPpasSQvRZtkHmTemmwZaQW4F9lh0052bGcPRiDBm8RJ8iEMqw6LjCxoD
kHSOPxuQLpu7CwgDz3UZiHQIJFdLvCDt/W+4e3DSOfLLxVs1UXGv6sIMVBc6y6xY
e71AhZ+mELF4LsCatcOWLBOcC9OxnZcrOoT5q4LfUoRckCzil25ndVHwjUuJdJCZ
Tsg6c/38229CuyiqRjRisyNYyflftRIQuGnPcDPO6AuJD3bWjqai5Jpc/H4enDXn
BuR6W6R7UwwIUcUGTrXso1DHnc5zJjlrt3nWjnZX3qXLiChDo/xvT/POpXCXHhO/
HRBeuZFGNLG+8toSMV18YSnsX7FgFr1VRaJw6LyB3/fq4uxWULfqefIH93rSiznq
wuOq8Mo1eKihVrAhe7xy/tFb3wHdsFERJQ6fPS4OCTcnbL/O8zZhLP+TfL+6AJpH
2IE9y9XyuiK3WhAlgyU5maYTUS5qh5NQwjZ5tMJqA5GKGwrvYbX8ZxDdGw52tmlf
VflnlwAdEtuF41+qg2o2JQodkz8yatCZS91cEClLMG9FDrHKKnYAGrfJvSsYBeec
2GmzLfbAFgNck5hoI6nIm1p0GJoGUwyoHIuAIhnsp0lFUJd91FrNR7DZvW+ail20
Ermxi8ehVf8ATVBQ065+lCcXwDK5nfnbLTtwHluS5ojn3oiXWUWBOGsytyT0SU0t
S4rocAoktCl/ULWbmtcPIp9bswTXQcgiQ88S2g1BZFLchnFFYK078YQ3D0kgxceC
ZBYB8SSfZKsMrU/dNQBLOeYxO+1sy5jOGWaDe75TTGXtRNshYomc6PPa/sZy4i7S
SdJ++jkY7JOLS/zvYoQOzIToxd2I1Lh7DPsqhstgmCPQgr9aoU14fLFxV2YPL9B/
nqlW3aAfZqctuTD6IHwp6pJU+Zq9V9giEgxEVGsLuD6RKOi4VcSp14EiwyW6LR6z
cjUKHbJ+jAf/rLqVs7ARs89Yj5gzICAjYex8rqPrWFxKswSPHs9mpQKkHUSVc2HW
aPGfP8wCcEtnMVD67vkVxbbZEnod7qLuWKY658cOgTQSev4TyqAZfLT8YgiptAeY
r20YD72lnvrCYXY/CxWg9h0BmJVsVLUjHwYfhgV/bqehM5z9zdWlhhh0rQS6BNrJ
NM6T88cwIssuo9s7wwbY7h3VSlQ9MI0R03kuFCXRY6J/u7cCiQISJBgyzrzl/IoL
B9X655nVMI9/H4hoU2FUd1DPlhzHM94+KEAfIu1WQ4uzW5epmu/ajdfsSIWnicKT
I0u2FKMxogvFAEuyq4s79I3CSrdN+1NbuZVv19lDv4QiOajw+lTKrt+wl+9c9Vqq
l53aBWBvEiFWqd2zOe8mG0wS88sqmBYZi3unrLqIrCr+mOnPOUcrPbEkiCNx27Fm
XcXCeqoIlmpoITzTe+YZGulddkSGy5fESB+yGFL4jq4LWhJY4HxPGMaJSdnayvL1
Iteqkic2L4GWup5Te3BlbcPhV7+2FKRObSFISFNQFR2PluBhBZx+kzmw6+X5b7v8
CRRizq4J3XDjeLMext/c64JnE32PXijy+XkRJy2otnU4HwecbvhQerqo9Kk7gzx7
BuiEODwphRJrm05Xd0eawDCIYOw9BmznHsYjsaSfZtHp+JTX3Hz+dIO4fDCqp4Is
rIsWdKZRZ7iRZThrCxMXHx8vQvAnUWEN4dkiQvj8K9xXx/P2EfYRcqPLN7veDj6N
G6YHfD+wOr7o6ZxUnKopAMAXcDExqCK6qFhA9oK1gg0wiFJi2caEvw6ovnXdWPwZ
vt/v+zaIoiHXjLQNPb3GiMA6BMX6uAt6FryUhj6VswjgfCB/vyjxMj3eCSAmn8aX
odcKfSUKvO+Ml0jekzGJBaTuu+guDEZmL4Z09myB5NeAeRj0y5L+PDeD5poatZi/
9Ym81hdExMHT9Cao3w3KHtW1IklVsSKsWNCWmPikog/12BEVQ0gvPolKYBrrbwAH
7BojMrWGPrRwDfmGl5mL1ayUUZrg9kJsDMs2v2kaPtJrHxdZvu4fTdwCiEd6UKl5
XZmSjkOgF+DMDvpvKEm8WBTZjBLP8iEaT+jSLPjaGoATumP92hqEya96obtA9sks
thpjUPjwnsYIGjJ3sOkTj9whQPaYP1IOZj6wg/3pLrYz2bQfdRTSD2nINQz6vrTb
YvD+5WklZjhqUnos5tY182pgaeLGwlvivdIVpF4RMCPS4I/2tbiQ7yB3om4bCzjK
yFDzdU1y8gKTUsuCqvCnN+pW1U/JAP/W8lLlWDcXj2jJGpvSN5OaoehQej5kqaT/
01Pg8CCBb7S+vlcMCnsyB7QmutU6toQ8bTa2UU97PGQPRGeKfMY2udrbhRXJQ1zD
k+vCZx9cy1cJY4Kjws9EMXdZu1G096npG0TKN7BHe8mU3xBYzx8BCHMQ7KqRxRbH
3rDkjmf0QweDKn2JUq7yZTjz1hlfkFykexS9KSOMqqxrqGEtMVhCgyaNhLLtmyp0
PggQttNKX7Z+fGQlL0BloByjkIAfRp/r7iVuF+gOxoGBb14zSF99AvVsqCit3AWd
azovZ836apIYe1/q5sU1KtTiBIxv122HCNjGxKWyLIHbq1V95FDzO+I19G7R1sVU
xCBXUgEjfQ2CDqmWiB9Yjdqx3We/UE+mMUf3+p0QKMskRJX/StNS51YXi4/TJiX5
TIYnIbqHDqTMklrpELxR6awDlvEhEXTElfxg+g9JFjGoTwOrCm+bvxPRhiXW0cC9
w33Y1c1sPtu5IkjyA7KE1m4VAYYwPV5nmMWwx0jk1h3I5+E7z2YVBCnhAAu0DVr1
VY9npe2t4rD+Dv4nP6oYu8nbM0X4Cvek8uvMnMP9ndQVdYSJAFWbAe5YVZrxC1FR
gNyxDZpbpW16YHb4JQb9bqxQcAoQk3lfTWXB0WbX4FvI5BBkGDnTSy8U7kcFlIpT
aNljyNLvJfbN22wG+ByHyu5Xy/DH9feC+zFldbmbj/IEu7VJUJ/vrddorYdmyfdN
GOHRHH7aT1kh0HKAgew813jgF7H8vbGgbutwgaHHIG+i2gzVRvsBpyedgmayuyc4
kG4B9lNIZ5fzX01PVR+GzEb7ObFrZM2DLcuORIMENA+QEz1sG4R4PHCnaW1jV9Yc
3/s2KhyAK6Z8DDZJJddnrFpTZbVv8igdZZBsFoquiqIbhmtEyRCVGAVsheSHTauU
zuo02UdW8l/EYiCohmxVVKzGvPKlXoMpBcz6/RK/r0QNmOur7yHbZRGAH6UD0OJc
HmoZTe45TbFYnDtP//3zmq/+K7nav0cHu74kxry1LUBoH0W+YyCm0ls/thr7Ms7o
rlQUS9QNeYHFKqkjJ8Eq+0j3+gKqvBlTsf9u4lzBBfSRnZ72Jv7AMF8U33YTZdva
ImzzrkZWVKhY0R/IVLlYzgM4+K3NFODmu+TMU8VerBlK4MbMuBno3aUt8CVTl0l7
OrErNFFrGv2MjNB83psnI4472F5vDZeMKdpWommhF27/d2wVoPuYTBsNkhmVH7yY
6t8Hxqr3a6eYfWw5owUScD0/Q/LTrHxbMohccscXL7KvAYCWtg06Br2W7BBrrimT
mGcORMbRYSLi4KoVtAKGTUclgpP5J8Skfyx3LfuQBIj3C7huD4m2CGXNtQIc5xyK
QzViUMHpCQVjdwJG1SGrHfQJhwGhP+KRV704KrFfz41Cee37RNrSb8ZaFUoEarVC
gh7+QoSlxKqMFsepBjBwcN6C8WE7B5t/EbCMd8bFlAHTcyVH2N0UAzTqRjzcw8d9
hVk97Hwtni7Zjm/O/3TKSOMMfz1bB+sfbn4sncnLiXviishwY12Kk2/iM2pYK6SD
xtuIOfbsLyUWivBHl3SJX8EXd4waZQ+fagZ6YgSW2BJX23ufmXnZReutJb0CQtLp
yVObt5xRFTBPO+STw8gC9SulW8Fmbq1zjrIY+AKrJYE/WYuKoqYIOquITC+yI9BD
zZdzBD0rvAmjv2QDySgb/yNhPBf11fbKAwX5JNgWd8vG7XpP84Sg2z2nNzNk5gIZ
+ZOlKDHFvlr4ZvmgQn+v+ViWiwQesFoB1lv8VGBeGnT52XPD3gngjwupJqx2wb91
pwwC6KCPk4pxQFbrUxvsT1HUm8rUv1lflRvoK6BeXWowp0qHRSdM4iZYIE34Znzs
AW8t6nxJ+mSG2T9R9WPJCVCwSqij8zrxP3O/stWLLHJjoDSCtxIannuwQXd5S9Di
c3DoNGIbJlNRTKpyxSJRoU7Vl7h73NyWnt9ZT/80o5jB38FhuXdY+2WoGUMzH4Ty
clZyY59TfRe/ePdymDIwgAfrBG47fxwI4TmUtW9DNZXMSOC1rHIDoiodQ8kLY6DQ
PEXyXD8Ph3N3/EzrITPiG5Udie9ww9EUrR7oUmJ5G+xGvUd/HSUo1w8Tvt0HZL96
/w6osR1G0xglDZ+i27/jyNG7KYjVaquUn61DIxXrpS1QoJaWbaIDUWa0PjTUxLRE
lVMaIMZcLFiuQ3x9qSLE2WMyyLIIEAKGgq9wlVul3bPsWwkTE1AU+bnY2brINWyl
i4gZbTOqpPpb+4PiMhMC2JK3sbE+7PF6mdiG4WQs4o8gC4Ta5l/OHkrvmYqnFsGY
Twr2SvSM7iUJWTOinwtqzjGZbnaCFDoodSYz9VL1K1M/bY3JPO4eh/HQwUUbDWhu
Nc9T/BhbI/bpFI5dTLzcTmGtGm76bvq7CUKTQkXykRJod8ahAMWkrD5uvwXD/8Go
PGCKPThxy3b4vjVGPLy8cU3BJ7Dezmah7zu6zN8XkcVR89d8S6z6EMwuG+AMW2Qb
c7OARQ7g3SXAMxEhBLTWBcKFjFZtXvFuqSJhqRuWDBFEg/wM74aA3KsIT1l+/O+A
w8FHhas1EgvemTDrJCZbiX28P2NeB1LTV/lA+WfLfjuNtwoCsXwoCu7PPrY9tisj
ZZESYvY7hRpMf/bga3oThow2Q1KKAHYsJrAvYXYFRF7xGjsCQHiqfGRBhz5dTu11
YTYqjdGCbEBgMrDf0QqqtPaBbNQyPG54eHDCdwL1auArpm4SYjTKxDd6CvVicCQk
uJY7WEPc2kzPL/X1qWlJ8Pb3dQ1rP1G6v6mNjvTfDQ8qJ1SkUcD8f5PIq1yasYRY
aEaHGHKd75s07LqEjbOi/8uLn+vLo6Jm4HqP3ZezwNT4jADA6O2d8d2R4DpPjzcW
tsD0VJq44xHkY3TZ8OEO02vkv3jK7CIC8TikPWyV3Y+iKQDFZbHIzU+LrEO+Qha9
eJCUSlGyVhhKtPN9yUlEhBBcFPQnyKvWYMv8aQELPrEp7xc7htTu4c3YVj9qmChd
c2uU3KQJDubb2C2SfWGqghOtS3yxPkIc/0Teel11P/KyXI5eSyIfmzx4mWyKMMyi
QPaJxiy8vtPhTWjhEcBZAYxdNaZtqTDlq5aU6i9TDzaP2qtTJvm/G16sRk+fPv7Y
czRgGV7LkS3OwYhGM0CyNol6qvfPNBX7/colzx78eIAcq9dG7woWHaxGumDLWEJY
OanE3YwFvakY3SObMrNPrEqOlb5SLU7bThDMfxteQh55pVKcsBcgC7eKrFC9ipd1
eHSm49pVgOWACXS16PbCRJAmAoEg4e5gu0RgJjCDFafV7k45rI+D8WH4GmRw5Ia4
foYZRJSTCBNilhbjuBtflU2lh/pbEQY8TEng6RXu4s9y68hTWabGdzSZAXaAcva8
j2lg+Sws+30CdpAiOOYfnIcDEdYKKDuOK7IVqog8CLEJ0NcUQvTFxranA+AnXeZC
NLs/N/GU56839r+WK+IZbX1m//0VPGEJceRIomdb9FBG56yAmq+Z8S++Nven8xCI
GLGNYUQNpRMidKWfTRhos5a/ejOQiG0pghVgf1i22TZ/TahDjlkVIGfg9nOrsIWE
AuMJWKh7voEpEB2jBRfXjAylk3ahe0smlzEw3Vc/zm+rfoFLotsrLnHA0sD73G5G
c/vSOq9/w8DAhNJW/FOBEwkhZks4AxOg/bW1VGL/FzRtQe5mtIX3ymBeZIZdLJi5
cNiVLyIDXOD5dcswB4eSDCf3WzjUrKmnQVzcqCJqUPDCHxeH+3Ma7Cj0ROmojltp
0Ui6PQom41g2vyBHbPpM4y2Ei6NHGd9A9C36peyiFJ81Sj9b8xgWPZayUQYYSF4n
toKVgPLyWfjQtQadqR/sHeq9OJp5nCGNM/x5TCcjTtebF+WsP0LqhyiT3LC3WT6y
G6RxejaYhyRQ0HymdgPMfZw5gjTD902X/9I00DynFYNyLmOEu9fL/Q+Ygf05vWkk
XI6F0S57Z917PlAtyTYA66hS5TGumSYFHmtYywD7sRi+BXJ343tmseVwsT3eN5FF
rkRk9+sz/DUUCcNtF+XWObmkl61cPaQF7zCqdAxaP7ZF5tKkTM+27a+MmWcot1Ka
P+j7Le9Hlraz4G2o7C8tCxiGM2GJEVyvPlGQwbk7MLxaCcZc6lSDqGczHSZYUHgf
094tQKp3tBehsPm2ZVEVUBcXF8UrLVe7PFFVAZXpx6cSKXNbvdmUC1s1p0LwGVCj
Qtvu/Ot7ctxq7yjF8x53jZnehtXfCK/bjiEcOXkKgr6xrRSBruiNiGBnhsJBveD5
LREJbiVl7wEcx+8ICMGM0GQHExO1B26NDNWrnoEQbezbgy8bK+KZseRWYgSNvjSV
e/U0Wf7mDxuUvghE/D/lNcpX1g9Qp7jM1Wa1xBHxzLqQCoDCKCoxJDc5QMUR8ys1
vvVSTh2rpyczXk8vguWCjmFGcA0bsFTbLf4N2740VPrVoRZs6PfwXqG1UmrhifZI
AKuR0bfwP/xYeCBDr733yjmv1q/IpRmmZLGhwerrMUee3RJ12mqx4R9JJSCrPcGx
4hEaQS3R4jmexW9RbvmGh1Ed6qnOZYNbDHGSn/wdNZ3QiVWtlBJjlOqd/awR4ylC
hCJWUzCMHGn+YFl52WRdNTmX9q2HCyFVXZYAnmGcWG/hnAnLqgTSfhwPzri6iheg
hqSy+7scYmRRVOSf97noZFAjS6QxSJK4QiDEfgQO7VvDid8Sod0TUizyGM0uME7c
nW8NAoKFu5hiycXQ5TBzgtrmymHUr5Smt+VPdSAdWxc8ZNxu687HQzMYaXQkb327
RkfrFcQr0CF9XZm9vsksyaL+gzBX7P2Nswd+kX8kzzki4M5sL8P/bakzuOufJSyB
SYqQZNW0N/FEeECgKmBg4fVn/19/MYBtKBLWPC1jNcgLbVBrpP486bpdDZY9kH2x
yQO9rBKFFnFOSe8cpbAsLTiMd7fafCdwFePMzo8N5dBTFlycnege6T79nfVBCDui
Z9VRQk9tp7JDopk5LE5HUstlmd6nZ2lS1rSAEuZHnsShu/blJQSnT8NivjGxNt9j
Qs1NY/17/LJX9Md8NbmP+doiOy+ajLGmlaQHORzGxOEaxgMQDi0fHnzOtwLmtZlg
e8R8xpyRqsqcRat2XbOLmWVeoXYTRpM77qkBUeYbXtRFYnwImix/rWNsInhihNUW
a8pAWUtH6dK+0fAso5mK2tn2l/XWpSX4ZSM7ZXRlQOo9BAoqtCW73+behF4ZaiZD
/u2tLYPamB/SGPYk8hh5PNX/DOnTDLM9NIl7YP4xbanMRddrGnCfn7iBA+1kBeIo
Am4O19bij7oUiEbninSgLxQMSgzEkmPcdgtfv/p0QgAZC8MtbLHSXUgDfFdsv1bO
tF9BxjmcHkSbAl6FbYrGGiHGurTs9Um3bM8tdSi+4Fy0h+cu4XQ5aNL+3KhwwOcI
4h2Rf5RgM/XDLA3Q1cwkZqT5+xh2199OOZF/zzv0BzsUhM7vNdQinAltAiTcQxLM
m4xyB9dGswydnUwvMzX0w6+2Ads6Xrq2b+8I9wnUnLEroDE53CFRqqc5cDqz99iR
vs9e6FC4lyjps4Y1hTwVgVghJldBhnoHBNbbYBj9Z2gqrEGJXEjS757ZIxi2JQRV
BC6BNLZpMkNpKUZCJgdT1VXy81S9MMGl+Jk3iZOyPvGgr7+YPzJBgN5oIFB42Ndr
AVePxbEfcNNvp/1HDDx2mAEYKcFJ+sufhh7oIos5P3vusW274uxOPLs4syO9IT+M
vUGG2PXWDozBUXSxqZ48UclKBmdMelMfTR7Q0YZnr++DTS7FvbkJ5lWz9jYtDv+c
rbqlNnBDNzn+OupqX3SimfpQA7CU0IcnWzCJD/aJSH7B6sEw1gy09O4kGqelftgE
DJqr4JtONjBJy8ZwFSQQVyN8akH+N+otwPwB7/Qx1JbVRdU3PRu6bgAXitn4tSsH
gAUtTB2e8E+m180HnU9lilufqBCys6dRL/eZAzqtBAFf4AjLlfNrtOXsxbErsnzu
SBBm4OPHeGUM4pUszUI3cX02KpM0kFBJKdtZl+5ImZtVrqOjs2NzOODCFoY43pg6
M62RUvUDmGrdfM2ezf4BeQkKmUilZyWUPr6Hyp1TgymvgfOVv6mU1Xnt4lNya19z
nxdP8XsiH6T/TuLzqe2QYqoDdulZp9jUXH9e8Pl+LSeShA/7j9Fl9NsHMYCnxaFA
GXYBzKVyouGJPtZ1OQR/L9BVQJWjfqFmX5RR697AbrAEe99Nj8zHPno2yu3M/IBH
WXKosh2dU0acFOe2efaXIFMfdQJ73b4EZyQJ39+hSSIpqegljnT5oaXhpI9Wl9m2
Kd/rY4B+OXulwqW8a1w+B+b1SHtoh1qsItIpBw2svH1Zp7cImCdrfVM6smRmMUAW
CsEYoeisH3NRdJDmtr1d1/oiOjvsBLyFBsdYEQRWPLERPXdUckopSKU8w2uQxq2o
eNL2T0zUPXdswtVwS93TophtE+kzV3Tk0JTEeeJHzXVxSgnzetNNaenxKrvuw4Ik
0o+9x/34hS5VZQuWZRWSwLQwCWfkL05y8TMCEFbn24u3bdBszdPHtkGCgJPK7vjl
aaa4+SntK5oIXBOiDY6VkJGJpm7JHHaU6riZkFpwme0T2g5jfmhNDH1bwBi6+zt+
5v+Qj3wCgSo641yCCwgPvFbgTEEM2zNAjsAEB1Vdjy3+I21encb8v3m0x19P4tPP
05d6hg6fuiJ5a54TX3A1si6hpmwsCouVNrHIQqf4dUK/C6XzJGDBioExOT4BX725
I9gujwWWJowV4SV7XlrfwfjNniUmBhcN3ICj13Nsh8LUS9KH0WPXHv41Ymbz6Zrf
1a6OUm8BBRdeY9qN/pcHvRur26V7P6WMM+0yVZZhDZnoj4pJYe5QCPAn4p8yJN36
73j7DA1QB7uLlrHaG741GaGuadLqAvcEbDgPppFNc6kizM5akDPc4W9yq/KxhD0P
dpWSmaYn0xd5qs/HkFLJIyRCzMHIzhqAzovwlPOzcd9xptHsrwpf5/yJ6W/94R4I
XpqXdZXVtltSwV5aEQUP727wQOZXI+aohAS1LxOKzXojHX6Z7u1/2+FYjWjZGzTG
oYlRqNkjRTqlyEd1czYSzEW4NYacTsOoxeudRpO2++bGbKXFfXx9m+xuX3/xHHD4
NE7mFCOCeYuK2rFJG7Vg+m8TXtSpYxkuwpcaQBr8TMezkhNbS3KhntNnuG4g1LbX
TBxJlrzIwgk9u/yQ72J0aNlF3YROnmbI4qrdx41zMbyvq5cxtKKKXKPeFaUpnUom
1bGtjLjzyuWgYonxUscmMMt9sQgINuyICKgZmXA7EoH0kQzvitg2C1fl6YXwN+Og
foBn4eb9nSNWnsWTLlcXfYMdQBeMWT/Dy3eit6VOOzFt2Vagv9bIjSYmymEBN15h
1llSnYMNXJIA2aMa8uAnijygzYPjvP4djM1IlnSZcOpHOFtBwQiPLpr3trzQvZZ1
v+SDYZfXOqqhzHLtXFJ2BtDKhImA/sdO/pQpJ2nTL7U970OtCgN8a9laNCgzfCLe
aTjmQS3hSl6WOeHsLbti4Apn9Y5d82MsDj189B4X12A3/Rhna0OpfNuZptB8V0l+
Vtcfxzv7IcchLRgT5x6t8shZDJLYmfmmzVvAyLKfhiZ5ZFx4vlARIG4bDyl/sE45
cXVtQtkGSfG+Ly6SgS2WMUDKj2dIXbjoQtdP7Ifryx7qvgFAIFQu2frwu4SXZcHT
Ols9V+0FmUvVWwXvafvUqqNIascqL8Cvyk3Laqpu6J64kJV27HAjVUrKjFl173Kg
YsRI/jXuFIpQXhfgrSQlMRRsQi5w0ccXjn8EvRgXVkeOOY1EiCwCQmHqH6OvOBl5
KK8k7zF/U7T+JhrlvZNG4jjBJinq3vSWHhE3u0LLgb08PTHKU9c8AN0GtVE4j5kp
CNgp+w1aSA84JXR/1ha/58IkXPdiYLm+tSL+N3w2cKgdhygjLt/fqSpHW5k/tiqh
KOdQTrylb6S+G/eROhynWHLHnC1ERsuAnV3uvIGIkPs224Q3d6DhcnLMyEQ1AeS5
iKLam5sZJkY2ahg/AQT6yDAMuThjx0TcGaR02BI3ZdAwbMUALAn9R0DzWEh0RPpJ
kPOTNB5UipLMGrIuEAA6wLAegpuB5e1qMBENp54C+5hsmdp/41cVidXo1kvVqtlm
yGulSbhxx3n+7OtvbJRyEylRTp/cUeN93oyd9qxZdRmpJIAJkzMDwRplhuqZK65H
yfATsZDoY0NTDlCrXTZb3fzTdEr7MTLbBc5PNE3t982L5P5qFtzZwFKOP5AF+vG6
4ptNZ8W4UdXvaNocv54RpuQ6ICZXae+hbM/fXLvzXmNqVynJn30O2RUdTTCYDSsO
N8m5bw6nA3iiNUVJlQHVg0LAmyS9tlh3BSbJk+tP4cxPEcVclfcrHTKBfQ2S9kQ0
2/BZqpD5gdiR8Ni4POzapt92Lhw1zkSdlujxJXnSxx2G414YgpY5+hzGkrggRvsu
QYBpwr3LBhAPDaXWvbwTnv642uplOMYER/sG9RMqQPgBF+HjsUIS0BpVD9aXfBl4
Xw7fUOLFOjQZmG9PCsC9q62GIiG4RoKBptn5yEmmTKVGp2/1BOSZT+xAMrkI+lf6
Q2IDcPhAkmaJ/FbG18sN6AkdnVG1R2njeMjX9RqNXpsrcc8yYIW/3COvEn1sadXv
z4lhkKklSUZTOMX7cJwqXD7h7uogMOMrH6lVn9vPAba8T/6SRYptiBH3TChdXGB2
gGN/Mb17SN5BDylrp+/0A8wXMjO1q1iR6wNUBtNlGagbo7sXZu8RFHBvsoHiLpoW
fFRQlDbXZgAgQMB+W+AyMe2bNvJaiUZELodPvB+BX/m642rQLuRjnlS8LW3KXf89
t2zq+9n5BCmiUwdRvB5kblR97hIq+pcrCAcmHraJ4PWIRV0wnKy2U+d4ak3AbDBk
2i9qoHBDf//IuUOg0nnKGc/mBH+fLvNSey+GpPQcuP2ppxHdi6b2P/YV3/2XtBxv
cuDyGk6dRwFJFKfB05k5nNOVunbbYRbuKwwNS9n5aivpwFU3WwIAMqbT2higbP0M
3yyjTXbIYDNWn5A17HfQuPIlquTBas421ku9yhGpqNS1SeodCxMndqc0Bmgo9Gyr
hOdvggwg5FmNnSyUV99T2LtBlQCINHJgsHMB9HftqFgLGgoXmD/ftqdQlphNpT2T
0kz1U92DhV4LWeSTqm1A+NaXsnj08U7Fqc4Lf2YYcKYWT7+ynFDgOpTW0ThougAw
CAQ1BqfvTGxUXx2/CBwR0eacWXxJe1eEDAPFLbFXcWeiBzO3f944ONbnZAfeFXLr
qDHxK+yjMJ2anGKgcdHo6wgEJVy12D4SZ/SMpjh4dZBgfKCPDGvVUYzwV9M7yOoE
mPWB6Zo/OpJU/UrJfza7sRuHjDCmugrRWw6OeuidKfd1//cwQUT3r5FeyWQOGfRA
ZzmnMLzwJQDNEmCkAHVmzGQQMtQJ7OovexZUvQQVl1AlEYHYmDJ8nKKJIfUmtwqf
Un9kcKzii4M+NGVNvxbpdEkfu5P0z0tuWy1jU+oj8xL3XmToa5zCufn3oKK/KFZL
+qisE6oj/8AmJni7lNaIwlgLI70BYP/GdL2SzWgJV6AMRH5m65BVeGTAdsQ0XAHX
iJSnmHoFiC0CRMGbgcGRfB0Fx/6HtHrYPuiD8ehEWLsJjS5j7DHgnvhAKG9d5+id
u8tCpA4AkG1kcQy5RlsP7W6QvDCP6I88T76v+dDk+bR6E6CuFdhgGI3CeSzbrbDi
2lt/u/aaL7qfSBaEJ5i1tOumgVF4dXtV5x/Mldtd4ExVylVBG/zYDW868gOeEIBv
nn1zCBQtDmWF+yW8cK5dvYugrDLtkkLO0DpFtMdR4sOvoSYbpMuRJei7CVsWbTLt
aYXF3GB1j6W4Rvh3/nF3Jhpb9D1rvHNrev8nA5aGzm12pzAekf7N0NpREypk2WP4
drFLFyuZnb7tkH/xXb+7FtLMaCQ8skCxBztwQsGpoK+gcIqf43O3O9wMerrw/kP7
UBMTO7YkAkY10HDfAL2l/8svX/2w1qI3rBF6tmXYp0EDNoyba//ZRMmYFqMNGBrD
omy3KeZijrP9UAdsM+wpF3jS2cM447fhEHqHKC6Dzk/qkuV00yEpPxw7dhLB7GUQ
86R55K06OjDvNO0bBFcnZN+xP72n0d1gfz58TaoqVV6l2IlwlsxF0pUyQgwn4khK
/23CR1uLUInYEPhpUrZI/eaXSFaaH+78GL4GneLAozr5DCO3v8eZo84FX1LLQnRf
uR3gKlEIuIlvft+EM52ACVku/U6voTAOx6WFpZGzONMnJOIHXvCp6rCKeGXWe9eH
2xINqxp9Cr8W/H6aT8W437X0ajDv4fD+UwlBIqt7ShnhPF3wwDpY7M34y+w4GCsw
pCycEqSU5AoFIQcoSwPH+8AexsHmLHpUljUyelqiIsFPhfOs/y2W/3jRLbCNdcrr
nW4iqBqZDQgkhR370Irw/xt8uTwo2RkUcGyZPJzlyVYQ1vsuB2kjQyshX7FW8Rhe
2AV6X/GwkbQUBVNXbrik3h5Nhqka7MfObuohQD/Kq5Iwwsn1mljN1mxtvcbck4hM
HLeIyyNh+xSjnqCK1WTRXxZtMEuYNtjTYH2NtD4C7oeKzF8b0UJwJ47/GURl1of5
NdsfzQKf8VvNrGJEi7unlrmEOHl3hhqL9Cuh5Iy19bjEcSB58k2a3WRxDY0fnk6b
v2OV/skb2o0ZBepXdWmsVJDJ4Up7ZPi19dNHvV1GcsHG91O3JSZ/VSSUqgsSCZE3
Wj9j+2CTyMISDGjkvz3ALfNdsRqswImo74eza8ozaOrfmCMPwBOF+faRfKiFgghf
Z+9TYtnuKwPZcRK7Idm0MkIl5CUVCDMBMwfpM44DKj887fCuPW5/M6zHnno01ls3
jBuBD8zVHFQiiBW6rXu4xLBfXssj2N7xD8snL4mDAP++2fLsPgUEu0wzpzoxVr/5
Uepr3FyFXGXF9BqFtfcz7kLDvEpkGqf9XbKcy9C+UZ9BAvB2ubnjt84tJKftDrz/
KiJhC9Z/5r0EwWkUQOHYVEh0Nr58CUxsCesW8c93mFY1W2HBi3RSXyPxen6/CrSX
TGyG9e99463Q82vZVVvhPFRe9RHQlXJGNBcoOECdLopR0/vhUxQQr9iLmZffiFeR
1oIOdbbIVApujddU0YlVii7Gog6SAmWDIEA25/pmK9XjMd7vRjwPohYcNr2rVrPI
xlJSxDin7Bxv/AXBnRb1dwfLc7V5YoxP5XFsWhR3DnQlPnhl44qRM0c0L0BxubqA
d5vrD7SyZOhsWSEjbKBPeKXZJVXHUUcyiVDZ1KYqqk1ZiBovD9HeslkbKbsiAV76
bGkPxRIFMRQk0xTLG6zdUtKUCpeF9R34fuCUWoe+VCFE+nEk9xsrRMJtH39thkQZ
qTSvx10AWaa83eMh7+jP9KnOGDms65/WH0QFURb6wJvedy2LtEOCGVpwhCfiRioW
nTX29t26AHkXpz7LYUGmz4T0ct/3hhbCa/uw07OR8qcL3aZkPAtovrT0mh5UIpu4
22N9cVW7O5rQ0c1/rJ2IVm/vkud72yt9LnyrwuzRu2D94q9tfGgv4epEvqBvKAS3
toQyl6r4W4crHrmYdICDGSoYbvKx2FpWE2EfkMUKyorytGRVo3H1aXBSKBhVhp6W
id8Sc7DGtXg83EbxdCUq8MPCRH7rVqLhuc1+qtYj5C5lh/1Hqj15CM6trQjqkl8x
jUusjGB4NXE3X+mL5wWce06BYZBs7IkabxHvGSZLpOu54uH3sGojDEJMxcMd3ZRK
l06ZBwP8JJJiOb7afbnd2cBwwB+cE07ivvIHIn8oRTKuJWs4IHC+9wVNV3HM3+Do
6EQpTYNSuXR2UarB47gebGENlaSvP3DfUog/2YyRV4YVjtFeAwPeroeLgJy/jtzI
IZ7ENEhMBN3rKv/gUpehxB62C3EXUfS7V19b+yyFpcpqWLKSdkRkLdta0s3DCgsw
kFiNDC6t4UwtlsLwUvcf30ZbhfQo6GW8RcSTUp4fz3rVXZa17lC/xnft5drMGcEy
MV6NUvOJKgRVXX8XD2CLUqxzMVE603M+ag4H4+4TPrPYzFPiZKyVICsvjNc/CFTy
fct/f/5mg2A4iIu+rv5fVNBSsaOzqQ+IOYG9e2xG/iLJ5Ni8YwnbqW33LIkiiqv8
BNHt/EIPM33vqCsJ5BaFFNviOJR1vJwoKzpWqBDlhRi4Aw5iM+9gKTUCILzcK8Sf
+oa+ovQvoysY2qLNyYbbv8LodXg0m8P1sf41gvrs80yY3rRWXVuDn6LQ03bDW+Cc
b0oHdlhvSuzQuVnrXsRpZF107X1AwXQbJv+XTcJAVitU6mWJFzAmH6kstNIJndqi
7Y1VHLbSOwixWLjJng9lUvPGCdGtHeqFh8hluvGNDewCMB/jDFHMsMTQQ7eRlaE4
zLrj3jVFg2lJhRmCn0ncuvLy/vAVddYPY8y9CYTuCsdMXfjVY7AphgZM4yv3qj2x
Y5OtQwo4cJEr48Ws4xspg+cKnVbBash1MzswlaOm8QHfJxt6mJFUZ78DoJ1fWh/L
hOx0iA1i6SzW4BDE/98LFkGr+xUCe5/jXeWOrgp+V2rpN8uVbDf+ByJvUyAyhqgw
tAlPrX1id+roVWFYVAIWvUqr/B2JARHT4081nrxL5lCzUAbZPshVCVxoCUcMhl/A
ple9CK7IIV3r0gxGSvr7BT47mqCAH+uaSOOeO/D1vtNwlaZ+ZMDTI7eHHwHzlqKM
k1pgvuNNRj45awFZrRzbJx5pAhjBFCKRDbOX42/RgYVe7ebj8ePM7wWJPlx1XQSU
lFBzZbgN/vARZK/zoI6VCCQD42bWS9XfzSMAfGof8Ivn/fRGUd1mCEJSAiRikweD
N6bUlOAmUMEoDD6XthhKIhvh8SE6Ixv1Ov1LvdQ7WVzBCgitI1JJwgK9lVXVJd35
s2o0aVwjnKkqaoDqJ88je4rIfKmS3ecnvFqyNnN243CfyrkYyYgtLUwmoLeHCT9H
0TO+lQC5hNr17NciYBLCoa0+OhOzZ5jp/8dW+G2T3WtypubA5uV3DYqkCxkxX2sE
6K11VMD8DqzYw+Zld6HZfH01uuZ1KRqIk5CdKL5d828IBqR8XhjnO/KJgjzn66g1
zklPOAfZ0ieO0LoyhaCcPkk/Hov3OkhrgKJcFdobyEsDn6KsTxScMARaJPxBIE4+
fQLvpNGGWc0UOyaoMnP70t3MO7yHcyJuzOMZty6Q9jZhsSTnNv7vKxdKVl8h+ENL
YChZ6+eedT3DocTxenAidL/SwFRZbKjSwRIfTji85mfwFvi1DY7q4QuhBY0+iIcO
mTms7RdHyflY7a/t6/BXKZYkCvHjHD0QhmTnsKMGMsp524C9YL4r37gP1FQ3PhK5
WD8x4Gwj9Wnw3dl3i8on/Nrdq9XxY9fEEJh0TVmCqF2Kiap4VBOh8iRlFwvQ14R7
v6QxYh8hx3OksYY6cdekFfotAkYXc3wgM6Aj3v2Y1Bdfr6ARQDeBp4Ma8s1HPYSG
dHqrtVEFgZ9q+ijPc+Ss1pjyxI7B42Cvjhpim1K15ZItZhk8upnGb0ioABKg1B1p
Uxk+evL+LYAjE3it32UASEKDOcNJwoKbNyAF1xMTreTdOZacD9n5s6UJOpmf9erP
WS2MdQmKfIMdfV6Tpe65e3qhVguuUwZIlqjVoZxacp+1NiuhDXk8neNsM/oSYFx8
WnmOTADk2t7X9V8vA7btnzl7MPTQPd5SHHUVb3tfdGjDK93XglLIG8WYPnWD7luX
VL1g9746j2fP1De9iOnpkhgOZD/IIqi7mBcxyfXkPZfYJkP8GgE0+vmjX6KG51sW
TgKyuOpRstrV8R0zNK1oqEmHCUrBa/Yay8x6NLBEPp794gFmUTvQbraElpPmd8vT
GZmNfF5s1jYUnobvYxpikO19yjjz5xjEjs+kc0rmvfYfyxEvOXI42rYwMTb1MJua
XooCwrHkrdy82NC89Ysn0Qvh0BJFdl4dUktd5J3qn9at8pe5RYufzV0w2JNnblTj
y98QRJzJR/DlPRScSDT/ssOMSybLvYPaL6JwsUOqR1ME0gFF0LD5zGe6wdABDZ/u
aXz1N3YtfciGZ/YpvkMVbgWgFS4F5tEKCT7hkSE0gs1bNQvb2O+UmZZ5v74gkHMs
f47eGrkpxB9BHk2prd8Ahj79e7n2lRpxRr2yvLcDPzjo+Ij/A+3u6uSu5qVu5wH3
4JRv3Qoom2xyi5FNaeV1mo+oyrr+BjVAPz78Sg6hbRkMfNhKFrhC9vj1VHb7Ttos
lINCcxKGAMPTDv9zwxOU4y5su7G/51Ts4MBUfvr8qqZ606dZ0uW53Xce7bwR1vql
i46Exn6uUcijhbu8ieRbdWDZAwBT4ZxK7r+ATjgTQ43WfFmDVPB70DKZ1H5wy1dD
urAelhc0PeVrV+j44BvePEuDsMa3EierJJRjXRbrDgSZQsiy+aVUdhcMTsPGMKPf
uk6iBqEEPShx6YmTyQw4uTWVw8pPaVC5uyMKJDOLCk3gW50UWKgDGy9N9+9J8+68
TIqvAhrjx6bsWzZutGZ/h0LxdttFKOLtlGKV57NoLbPWrS8U9KyaP+nHp7/I0PZf
nVnBBnhHQSQOlUjf8W8EwwmrlIOvyeGsQVKxvetUVUrNonRjI5kJuLDpr79uH7by
6VMmY2cyYr6T/r/eECQlokcYJQIamvcLJ+7PhS/x/kwcD3GDax1w28P4UQqi7UM/
zkytaSFO2Gs90GO+bLdkEkm+5+FqbYPLzEkrNjEYwkCVZmqLnCwXJUOjm8dG0m6s
yD+G+aGqBk7tBhP+zkv9SdmvQmFF3DwkeZcBf4MCLalZmMahwg7AfCz7/CIi21AF
zNX8vfnmFRYk/dwZ8WSTHfGs7iXi1EdRu3LcDLr6CPMP6d/XYRAMeBiTWTyyFd2n
6pQK/2TxzUQz1gsy6+a/N0L7javv9RKVY9F4EGXohaXOfj8p7E1DvpZSxcpYGVwL
DnDFfJiCM8aiHobe/iBgody1y/l1+9WAA711wclp/qyibjf+kRXCdfheyLc56B4U
UrTcLyisbTHwUisazyzIp2LW2wjprxLJtQXNZ3G+rivfvLmaU8cCkJ55aGGrA8EC
aoca9ujok4zAmtQHeqqVYWykOiaZ29/okelg7rSZ4JT46mrT22uo8vfZyklVw9qd
3n0d+KlSe5y/ydexCxBu6OzwcE/PPytkF/8GL2BcpRqLhe+9BLr58NpERzR/7eOE
88shZurNspd4W3AS0HqVIxdRFLc8tmo5y1szCAMB2oUJPdIm0qaR3saNZL3KhpKP
mjzZpjT4pRoV0RsFPCGcC34HSKKBUDRDC9pCHyCxI6lJA1vh20vbsKbqviWvE4RK
jRIdk3E4nYrv3JLx/eR5kQ2izyvl0JYRf7sXj/u3famJKwPb+d3H/E6SfjZ38JNl
I9aV/W0ef54jUz5ohj5VbeG/dnKyd1oEKTOCqOPiytNMP17u2TMgjw1MIdbND0eQ
d3xWTIro98FzenswW+RvK/9zooovsL0zRQxf6EyOWxkqGqBB0JXDyezjyJENdeGr
Y2QLM5pvPCIIEXagJXY2sWkbSG3NaAwaZgz4XJOUXEvMdS2vySyhakmamZ22p8NL
uc1IWN8iwWYWR1QA9F0PQwHlMqHwgvvRpRHsxM8m1YrwkgaQSfwIFokrVQtee71e
uYBOQNIgpwCWrrjv7nbbQ0iaK5vxW0tOEynX9ZEJVOPooxAqtXCr9bsGTwpRbjZi
5gjqHuZsfmS3K0dToY8Y8wa8IWyXRZsrZ/N3kckVYcTGHs2Ah6lxMSNuafDZB0zN
LZaaJpTUfR7UuPQADNHGLIRCadYWaWY/iZUsEFB7Wwnhy7Ey5FfB7mw5DLUHv9W+
9DmbaEBrbueum0Zg/VAHIZgW7QakF2zFn/f4k5GiDNK+Ah0DUV+WH8UdsOpE77xo
rWbqq/3zH8drA2cHeUbeBpSXJMd+Gre2kVcOnwdLDvBRXdES4hH/MVtbXwlwLkCB
43MZAk/4+QsRVbULTdfnqsyall9t1Ad6W0wdTSFm/6laqg8YXUmLIspppY0HY+9Q
aZbZmbxOsguitxwSXgJ1yKpGUwr62wxcj48K/u9aT0ooLo2jPcxDLr5khfHueUal
8FkfT8SzB63jiqwYlzXEBBWMBStwNKde5kwZysiIt+ulZym9X+PRuSFEat0FYuOh
q4eDSAirW6TAvljikOAzrgkTvhl/92DP6NvArh7nzVypylyPwlu5VTaBQLziKbFm
W8dzeyY+HbP21NCtv1xduXklIFGKCWhVBt/KYMXir/JtIC5m98R59qWQjhidpxdh
zpIukkLCPWspRU8BpPUcD8/sTf1xnva1slCSdbTzhVWswK3Llpu32T6s1pAmzvir
gieIU4JmLJsMN/Uk+XQAZ2dfo1AtSZ8tZ+E+M/v4HG4kSGGDq0WYrh48Si/2Tm0X
IwbX97pIG3agcQyeXBoYNqbEQhqCD94TEACil41uVoO1LOYI+FgFmu7z1AbqFUdn
V4upzTERfhOYvjhkB8Qwq/uwek7pmX6KfGbHuN6m4CB+/CkSZZUg3CK0FY5ryI4R
3rE+AyYYY2QPB8ly4JoF5CoRB9SHaq8ujyNqe7VfOSWVjU8+SonNKcFJl60rdktH
uQ7EeTV7YRW3kQOhv5yWRy0ONSwp2c7NA89ewygtSJIDNf71ob5N2uAokGfqx8fa
Vxa76RdUDvf0yli5wER1tShtGOJzb6hJiQ2678RO2kXwwQkaGxCn2+gmf61avhSH
XKr9a/QiBYUCwGe/DH0u6UL5AI/zYnP6RtnL+0cDDIUT5MZoeQaEp3BNJPRrPZrR
/HXtQZq8uvT/r76jVIvL0QywvkPziJIAhaYdrQ0VaPXcGvtuy2rPlWaDvroHy6yX
I6CIEGfbB2F5kQtYegEkafKvZ5h+1PyKxALLremmGpIp7ZKZB7So40/wkxXtIcO9
ocjr2Mt7/sBFv4CTot5b9oiPz5k2m9wvtE4i2bMtocDjTDCNpiK62pM/DX5CUBvq
AER9dwMgMQgg7gzcPK4IPjkXkEHNkmdOC8hXlE1zJywoC5LYXJEmIJwamrs/gCgJ
1yohG6UamV/cspwst2cs489CFsJfNFwpbY7hjjWTDgSSrcvaWpKHm5kQPGWSXVvb
FAAKfOo0ZVav8eQTHQCizUuTgpIZQR8iPiWcDx5I+R5o/0BNcHyUiemue8qVv9B4
oaWI1yFOYcHv2cQEuAos2DT93tjF7PQd59WVlWXSnRQppWy2bcNOydndE+us+Dqr
Q0M1hutOTXUru5hnTdFk4kz7tnzejrZoPkXoMiaI7GOFj8BXT1xWq5n4R6CLa+Bb
QSzd81DTDAvB0qbSzuYsL47Z8iXM3AxpmVxrwOr30CpPI56jksttZpaZuFCgynCw
J3sUuenENmeoNNnwvdZRMxtqPY55BQmx2x27Ui6EyFSw257Rwwho6kS8voME6wQi
I/IROCU4KlP96Ku7x+5dM07lQGT8KpO9qV2+UmGwoSj+yIK2XAP9vK3kuh6gMklO
nHN8TGEokjyYbDOSZg1HVvYsw/8YnMPF5DDD2xaBq2Gi/Spe78pT+ISbn0wsEz5o
sCpEbqmHnfDSQV9KHtSpNnYQLG3dcnOmElhet2oDlhbnkS0l+ED8yOzRvWi2kUcI
7BoCFcphjgoRqa7QVjXZocHsVBtnCpIwNLXYxo4v1dF6jG3luein2CuZ0yiC7Qgd
jg55jNqokL8/OYSdQcP5p7izco+uuSw0ySM69dCR8m78sFEKPYGdyEKjpMDqPGks
TKjxECL7ZECe46o0MZq23hdqTr/Zl7IO33Do3hHplmI0/Zrg5BhAfIFmRrypHNxc
AA57Hof5eheocP80EEFzPzMFAC6qIKIkpgpPCGegJo9nTZqxqpagK5OflI6FdEsM
AhLK6oLoLlzkqS3O1yW/q284DiyNbdPwZkcom7M6Kezr5DHFDdAcujn0g2SKznhH
S8Sp5CailAyoDa8C+CnoYEJgoyP6oHqw+QULtcOwcljGNqK/aP9v7ICC3UaSuJvJ
zlyVpgR/pu3RF6JPq+8yIYRHJBbjdGKTX1CCxZ0oo+mPWv/LL0M/4V1GmbjBdLVC
sohjuLooDekiF1m/Mjk5Et3LEqRvAWGNgZPX5/Ehy7/QZjyESxEoajMmtzZi7z01
rgwXH+Q6gYGs3ORphE5LzrTqYRlPybqz4SZrojbKRMsn3IWiQ63AYYDOHBxq5Bzc
9cL39jr6WqtKixV1R7B+wq+XCh2Uji3ts7sn6FinZo1WyLa35ISjncbIWuxhZckL
BRvnWTbe+Mo/LEdTjNepV4FtnO8DIBOvVDF0PLXOlRVAiN46Dbfui6QklEUZ/6AH
s25SNs4floScyc75EfnsclxPNhxuBV048bmPHGKBOAl79M9DPUmmX8DcQCFyqkCq
EHUaiRwEvPPaIzXpphlgBUWtKLAUWBn02Fu8ypPw/PNzA0WNxqnuXm4dpduGGUr4
R6BBaSYHpC2cL6c9y4feW6HVhYFJjlF6bjfwtgEG1dITFuMpVBY/dGjYksFMvuM0
picsTJrbN5sEKlRTbLvmh7VucPXTeHBR71+xUNGJFTewklmxE8VnoNdLcqQCG3PW
DA4fQlfEV1n8MYk8A9hrs1R8fQ0IBAEPlwKj4UNkhVOddAhuVz01plbmiU7t7r+2
nwBLmr0abztpn6+UP3nY3Quj+BLP9DNU2TzqaBapyfFJ5o/Zfa6U5b9bntsIoGu7
sKHhX6iSo1CDAXPquJ0ast9vZ0V120S5/9kGK7W9uWgbMuD0/Kn2m/QYy2KdkcDT
jZDr8dNfB/B5TMKnbtbj+OMVnGlkA3E/AgooBbiAl3poG/R8bc16IzXBkzvj+u+m
pnMILMUAudO6ecTmMyII4pnqM9TgmNBgZ/rGdYH7Uw8Ajfp71f766q02FfN0wZ2P
up6iUjIUiSq0IWpyEJKL0J30FAG0l91XxEB9F1+4yNG+f14/SDMajv3rVX/Y0me+
89aY02YVOQXzcDdQaUEYTRR36/hs1OwF0JlC5ImGvqU2XAlSnw6hoiG5+QAABkFX
4/daPOYddnO02foD9aVSf7OhvN76v4YuCaXAmOfI+qhEDnLChCYb+Gmfr63ryANt
DMjxJ8jjBCDOMzreQfceFEl2TSm93aKe6jQs699oToIIARTlhVh/dssqqTgZ2xjb
kh8KVVfAzJZ0XF7CGp1WrumLWFvJSPBuBTfLl2uVeTJxb9c4UTCPScfGCLuXqr8T
Kw2ad3HqIkQQLJk5R3tPYZTZWXZI9wDQgzgDHOjQTZcHaXzTaddKVwJ+9DUVQMHr
ASFbwbs2Cj/vXt5RSc1LY1/x/PmJOefKryaXBkAauUxCRCJHDwnLYYLLtnBWDu69
lLv8p2S1KaIS/F2qkE0cLXoNoCRB9xV5ZfOJ9RPghkWRqcqmlsAQFIKQpFh28qs8
rkw3xOMLqATjfBQaRkMy1Cgo9QHC0K7FRCeOP/nJD6F2kkKomI0NYDTdtVgdYFK6
cwyWREYRib++gPQ8+ftMYoWB2xo/fmLLnEjhWd8FH/LNftk5PJ3P2RRU1ksDKfyG
sg1UOUPd46O11Z749pzvjMtZrU3PgY3msaSVD3WhYWq7NtTTJME510iB12lXb0ta
feDsSkgwYE8zPH2vagI1u5y12+3a0JXNadUnQiYQjcP/X3lknEzx65ntJlq+YPaZ
kN4Tv8VaMvGGHl9pQdKo1nvrwPZuT/tzkvTkfaObeDpbEddJrGx1KIQHMbfJe4mv
V097q0rJVhes87SnGhrzv0XLCO6+Upt3+TCgeWpKtDfy3Ge6+WyFDXuU60z07IRz
8Q35KMZdIenYPBrsD0FXK5aLR57OzXucg5jTwO4uIW4hlkEThgkIesAlSrES5fj3
ERRg85yYoNIbkh3JRFgFdVBbIaHh2m33JOjKrG/nBrOi7bC/xSSYtB8v3Kyx0rT3
izVJnxKhuY59Ogth2CfNidRKZEqm5i+fV19sbEPhjuyDdE7WNBb/fjSwDnf0xN9b
npAo1GjRJQLgH+w1vnHfHuDYKzJmg5IWH8cVUC5IEtWuE0UpSwzJ/qrZVEvhdc0h
4DQOqHeRrZ2JiQNgv9eIB3ZcO5mhT+SxX99VzW95/ahUkTEkKWeLKaAKksg7nem6
zZ5D6cDsHg5+42cdevNrQbzL/1hWG8q7Marg6VbWHEcvJclDMq+Bc5OdIFSw+IJ+
szK92pXrb+B3ElppFF418pglxn3073DKLiFgBbwKtZAxmD9+6liDOo5JVfIem628
vOClOebKFiGkM5Z9hpcaxtBZ6zWV75W//K2k8D2jQvVkm7g8FCciNO+JI+M0CR93
Aww7hOBUR8sVGZfrrwDTnZzEapBOg76SSBFdUeFGw0KND9gsXZhgahCNK7INSUcC
dL9/bZ5PihKmHeR2yUG5Qi2/oPLIWtb3NMmHxG9EFnHMAwUkuNoJTGyb2cYFBKHu
IH3z29rf1d2jkaVIwAYDZR5adnoJrd7OogeCa/RhN9UG1oCVUfKLqCbUixyTuPSG
SRysBBdP7eNj+VRWbxirFSc/ufporsmbHjmOYHLpK0fhSJp8qwp8zNn/nErGwLF0
AxTBzGju/qoUCqKBTZo+2zFeYcOY3zkEEhYDIy15KeaNO2co0Ob6F9aatCB8GKwR
ARVg+23UZVaEOXxBHItx4kIuYGSNbJY0oLURu1pX6J+KFZac4qPjWZIwoC2AvAPU
Ce+mOHhhoDd88G7STErg7A1ByGTZhX2xfxWmaOGUU90dZ9b8WEhh9TjWDixNxzj0
49IkYzLJ6zQd79XgWVpB/gj/R3ELGnQ229mnFHVAtuirTYrupncuDdCMC6WJRCgu
nBOTMkjOXdykaHS2URdnHKVQL0ldnxr2zgtuQ/BPOaOcjZpud0oePH4TEL7PzhUu
8M58We4wPl+DVueiEKx0gQruMID7Y2cdAcBZERZba6/OOpCxU9Uav81fTFa6cXRN
m9sulOm48X+AvnChoGTAeNejiiO/RYNQ+UhL94cIWVYy/LRKsk4Pdg1htxYRXBWp
ktH3r+Exhj4N6RY49X35qKumdzEhP4J66YPZ61xL9br/7cvDy04RqZ0lu1T7eAFz
R216mQEo5gmWPRXN8WGQQOek/spZSzpCuKFXin/Nx/UwqBnP8+2u2AyA7W1On5ja
k2+1eSkLcRTZpDyMT7iDy7dEAN2W8o+5e6ykKXmQIxI8pjlhCfhb4SXLHDgKnEDv
J+LTu4fVK0W7nzYM1FJ0k3D/2wshPLHOBOHnFr0MMwKUM9EFJjLBS+Yq8aRupicM
fadaHmqBr2LaT4amhJQhMktL11GbdgEyPym5psbDYVTRZXOkTVsXfPShAg/DJcnQ
OfA1f6+/TSzESd2okKdLbkUfIDZajFHVf/cCdfie1xBr5b2qrv3Ao1vaKTl3wdQj
a1Z6L1SV4mV+rGHYLkZlAILId9tv6uwGL7clAu7TNaBLgL5YEf9Hc8C5BQeUbpN4
CtGKZNVBpPgNZiwlip+4e0Ch5CH1/PF4INY/Lz33zJebK7erug9cwT5x6uhTPNpL
UiJ6F6WVN2SFlR4aMKA4y+v8ajkaePmJsQgfd8xtzyXe0k/+ozsXnJH2vMweRxLW
rZf/u0NYwI49gPoOklEIOuyI1qggFIhaYCNquGNJ6KrV5g+WIDieLACOTx4WxD/6
ZgSaJKJXPT/e2gsN+VqhtSs84HhF8jbGGfUe9X9CqNPnt5AdWNQg2+BYhnEdAk2L
B9oG3iiROG1fssW1epHuLL/ll9NG7OZ1LS58ndm0HauBNvBwcyQ1srFnb30Bs5Z1
XhedMrfnkU5jFVKkvewiUqVGe+aVaIFf+rse7WWrgX8cMuDQ2bbzJ2/TVTeYkD7/
yFScISmy3nXlsUb9k2KPK1RZWiSumRNKeByBRAYbJs1ye1VHuyVGgObdObTSOkrz
A4BrtTziRNZ0YIkRB/oQd3GS3X+XykfoTbURW+/vK7zgzBACRh88EAPv60La3Yre
eN8Y9WMmYM1OagBPCXz/5F2hoY/gooq2qN4aqvxVwWWrDtpVt/7laOKE2sJw2OTy
NhnRqqRSN7/1aFlOZHmRdwRfDDSK17IOBVkJgrzFbEFJNyYtQEx642/ljtIbATvE
FDBQydePKESNza4U2Pi8ljMxepAtz/jtQHF4aJJtj6TdwFsj17gIvKRYPM+QlJSi
xk/enaSjoy8aPv03/Zj6iaQKzKfJWCYijN06Czl3CAqagYvqWjRKbykCJNOIkBSL
oCoxssCNcRfhxjhrIh02fhI8WqGhdTr+E4XentbSBoZmHuaHdsKfnSSyjYTEXG5e
K5zacHEw5PgIGpL+fyubKoKyqQYfiq5turKMtZ7Y9Si+L+9OUEuVCf0j3zJorgiu
hV3+lKcmowgI4Qe7+R14jSdeVU16Wq3AEG7Fmrl2rNrMzY527rSOsXIBwLU4FQ0A
gR7dyBER1PxhlD0DMemYCkFzpbtEiD9Qgd7YUdZyIECXKtqRdTTHTWFIsm4AKGs4
imqb93hUq9HxD2QFkKjS8NqIjqfBLwJhCjMImy1cri7uO1hZCa0vOpcpcuNKJM4U
BYLr2G1BSP2YeRv0tV55lDmBKL4oQBG69E/nscX3qxMLQtTwQLDRC5KmZrKGyGA+
X8IoX1pShSkIc4SAy7aGmsDhFsd9VOKVeGMTRi6l6/4tL1G6kCz+Bnx9Kc+YtyL0
OFPW7rSYbQUJxlJJ1PeUjp0DZS69+Js3EKO2VeDQgtFUDyjKwQHsdB0hh4yjwqvZ
CPYpU+gPWuRLGQh3FXVBgeOBYnWxS9B6uoZipsmtJecBnqbafewTeOam8lyyCfwZ
uDgV53NV/Bc3rEZi8VuVFm4rxarfgCoZJNByd123oSraED9wrKZgMPBMXJ7EE28V
/UvsNTuWkpMaFfmz2+w/mGW3XYWRgw/Fgr+NmbUmpelz1DWAzuyfEd0MWj5f89+i
PyWknT3sVn8mGlK3Gaa7M1rnjMmDoQ5FUe13PHMwspUV5T2ihsMJl5uBJI5dBi90
NSn4kssX28VDDJ3to19/+JupTzQLq9V4qykyIdXkUXAWYHb3NSlumPFKv0QOANe/
rHrgxVAPlGkwi3lSbdrpVnS1Ggb/VkNwPNlrQoXvH6SO/KqTm6vFrLAZwQpLvIZY
YobDDYVN+h1I5T/z0tcvZkWlbkRjcHz3I05bqrEGCwdEzmU4C2n/aAphrRVMEX/2
JTZR3LVTCRL4sj//dGeUi/mU3m6zYyLcY4DZ6pBOkMEZh0TgTb9TWi0Orzs6mQyQ
Tc4hSH/E18uMSmkx2g55MgddkJR5f4Vk9iLbWURR3e0aDxxkTjwN/AgceIY6p6by
59cgHuFELE/BjqXMb8oNNcTD53sRlKx+fcBTENx3vB+aYILTjWc3J2Vycl8XDmRl
cvQROFVPTa8X1u5FPkmzttAQ85IPfSkkrE97uNC9HERxwJukw5kkVl81S9NaFKZL
j3GTwcKD1WRdRV71H5CpDp2utDYJ2YIxnf7GQVOkJuufwXQMj2OiABudeEjJ1Lhq
/UsvMLq2gZ+8FvYVz8n+yiPkoG6/Tphjh94l6+SAb1Wqo63NNbeG+qF/fZHXCnd4
gCQpxbynQ5VVVo5Itb0pYX3qylSUYErmt8Gjxukufd3TZommzOYr/prZyJs5JH2K
/t6d+2E87vCuet0bL9fsVIlgLJIE/tsST7/WEK4XHeBH8oMwWxGJjwL4GKdYv7lC
qhN3N+jSD2fHUvHbw7zbwVxKwNEsGmV+fqTodUqgjy49H+IW1WS0OFqQKg73eHXH
ruykLXFqUg3pLMlbnmLUf8VyFDs4wkSudESKFf2c5tmnEPuCOFKc0CvL5H1mUZGP
hrRqPSsNTPhKHJ4lMgJQ4Bnm/yW8ffz7e7WZANAxO0ygX1uWlqUzdJJdktj7AthG
SHj3JMzNq3ST3bLZDK9xGXXwOD55soCnmGW8O//PIAGGVHdyJ6vH0L6ybiDEdorl
osD3g37fxrLmZ3WyfQAjhF6t5IG7HlyQ/mgGTxXa/IbyBRCc5O7fvYQC+jKscmHM
jTfTZ/tPe7l4oaHUs3MW25k1N4QJSV7ARzM9ZY5JEeclZIsRHtbP+1af0VKaR0QN
UQNejr3KyVqSyJlM+6kSNeLLZyxjwdDi0FdGxqkdaLg/+DYl5C8yCCLTnWNle/H+
c7H+Yk3+NVVHOvh6xHhRoR/AHU4VhhXVeztC9qDTv3qqMdzObzBbjfGug6tMIU+J
+eGwZG/ZGTI0CMCM6mqpo5cclGfs4NhruRn2PZf0Z5IkUGKOrwTwyzeZWwH1GVsw
xGRoF7TKocKgYN1UpUQy9a+cc4vvz6pVs+h0o/g/JxZrfr0Wr6TSimZrq5AmNMtP
R1glzd/SZDOMbu1KxKHrUMuaXVfVsZBZLW+yHDaFuNfYRo66WFamPzzH07Dus0Xg
PsmrIagdaYURJjooryXnI+QVrLX0g2eZ01AOs28Am5dq9Pv+f15RM94IaIQJQ2/e
bZniu7pMo02BPub8ZAchqT/lDc5qkPr2r8P2jPqGM9J2i0mrxWrmPkJ0mXy+KDKL
Z46NbF2cL6lEOKYQ7zUmhn57Q9Rwj7EMRR5TF38HrlYI8K1GjHXejXyPGVsgWhRY
1KDM53ez2FxS0QFCdoHnikwzyhsrU/QXgpH5kYTiraIatYIhynCMxiZJy3KmjEd6
s49Gu8ME8SI31TpN9FbqC4EyohTqUMj+oLrnk7X/TumRKnVOfyRx6l8VebGdfaYD
GdoFpCX0It9UVSGKc35ZfyHURkJfr7DOFe5PjZjtCoVSqFTer7oNm7h6geiuEMpL
4414380oqO6INbU5gKyvTaPpbc43ZvDljU1a0l9+Pw4975wOltruKZvu2qgkctaW
TTaUjzHTlj7NMPEl8/MM3i8Q4MeCMUlk/KiMoDlPivdLfoDCCUpOUpr6BfKJhHne
Nc3zRsfi5dDX52e8oC0uLhDYOlUtxC50EcLQ/y3nqrVL9LKHpeuvvQdNsV7VdJZa
09Reh+djO4ivghuPQnGAJaqFK5aYyYkuVXy1axHP141R0r8tcbvwI70RwnGfD3rx
1vV8jJ0T+xqVYAPClK4+MKn3wquvMsw6wDNbjssdqmoj/MEsIQKwbbWWH0Mivt1p
+BU6u+VkP+6Gb3gIsnAQDZztLra/SMkWQcP4944Bkx4EC9DQW5WCVSF6QrGTxWw+
0FlCjacbB7QXbUtGY2IzPwuiRtBXangEvFMvIq7TA1p3Z9W2/cN15KBTGBrlS4BB
fxg+7skYTAhrbH46ZysnWUfXPeWTAgfvSi9OR/vxbpISYIq+FL0sNJ7IfamYyRHZ
Vf1YTnj6isFrPqpF8JY8zTW9cpqhxjTtrTWcBUVzBqCE+uoCZkE771DJf3Q9zory
kdJ7FmOAuR6Kmtl4+zrZhA/hXHoWURr+5g0jd32jFB/aZRvBf1Z3pwUI96ZnOldK
rnD5YMZfghNHkCkJfemgzI6JCuVb69ccbev/f8UxhIk+HUZxqFg+XrEjdf3+Uikk
VynMdlNn2axhhx3eWmqMS5XCZiQmpqXrAX/5LEO8XTHm1Saf66torKjcCMKs6Lio
uT5EPjVvfj7XNwEowWIVzaSbB/aBdtg0QXs6vamWPKM0ajRLrUTKnwrNrF0Zx5qA
FHtLxbayK6sUOux60T9XLVGCYpJpy39iZ90FfpQYAqjc8yricqSeJUrDnFYIpXqD
Qzp6rta+9lbFZeYLU+CBshCPsoPSwP4tOiAS2AQdAlS9EjJWOja8UUxcEjIbqfzN
YruJEGDn7rf1LFvMzPPCRNKZjZW86Qs1QXnBnjVxfIxNuBl5qmh4HpBlHXDCfkor
dx3Qv+pECe+SWWQmxeJ/YC7vdp0M0e3zM26fdKoJRUWys9G5tiPJ73wmLOZUxvhB
rZxhARrlmpNjJAcetYFKE60W0cEG5B7Ftqn2CWlRJnvyZc1J10dQgZMR3shRzNY6
/kgJUT8qjiZ6GXExCyRZw1fVMO4N2zBQn4b0BBh8r5NtRM/8bgDrDohde5G8zRk2
S0mMZ449/rZURUOAVsIbY966fvLD2VAL1WW3RSQW9qXI5O/wQbVLRl6GehC0h1L7
aV3QjU5p6LM7FpUIBTuSJ2S347DY8We2PHf0S0kcKe317SJMR6hZOJajzX7ulCNq
7DvglGPDrVMpHs4z7JCP2HeP0qRrhE327FbJtuwtUXe21s7nAHEZd9aSnUDPqXOR
IYA9Vmme7PPa9bwFhICdXtHErJRQUXIt6qBqWOQizAj0aBDnfueSrWCCUYUsjrCx
F30rm3/mKfb1S8WSiSX393wKN/4SwweSR5tMgxpzHVMe6l73ojsTU/BP2cQUbPvl
rhKiyIjOAjyvEJxiAVdl4hm50guE3QAfun4rZocMdKefFxD6QUgNEm21ps5L3xza
7Uv+YsBwF21MDa4UCcY9SQ312n+TSDLnb+GjjtTElkuOK2WbyoLB4vu0tnyRwXax
PPHE1nDubejcg/I3jk/LGnJbGCHwKSpNRcdrPX+fVZ6ij9RBXciWRXhR8+C62pYM
L0tpKPj39yoZGcDFnf4aATI0yb7aNJF0WYeSbomdG/5BAA/0JwK/q6ioaU8eoUdb
YHG8fHEAa4y7a4vlZqdLLPQjl60rLV7MGWCPKP8lYtRofOOZQsd0m/O34Lpv4kAs
4k+hkeqJuH+zuidmkI8rSCHI21rmOw1H14q1oIJDvqr+9CvzsJMxPkgbMQguCC6p
u/foWbFJGkFjdahkWUQfIj1ef8GgOk8o1nvYyd9W++SfhaRCVN/HEIRGYVWOUb9M
TJ4E1rJRxfFFxY7CqJSeaHdYeBVimQ2xMvezxvx89ibONNtDS/R2ub7vy+Lvs7FB
Wm9DhN2JorGL7PzWe56QcNeriiY/MeoNV2wBPAGtjGQRpXrSp4YkcgrFz9mLlOgG
ulsQkSeinSoVeLOMmi2kfNFdiM1iz1jJZvuc2RMMZ/YbUu0sqYargFvFqMFu4O0Z
KQ67HNQ6/j5OFwdoZjYtl7Jw9Ls10OVx8B1puVqNvIdIZadvF+VpEEjO+cFBcBr0
KxyDSbohhw9tvB7byeQyQf6mHxuM/EUPaEzJnh0NEy2Q9DGisMSsdfU8ryToRgTy
HGFpkNsF7TIU52IN7nTee383Pp4irHHfMWCUW7JTrRWKlBRm1CfmIAh2XEtf8NCQ
m1YxOYTAJqj0emhWiBYCEjDSfXhSWuHF7IRGasiDO7FdqQUFFImFq6jXwjdO1wuq
BLAIl73qq2BNJu9Xae7fe59bXv/wd75DbFF1CmSVkrrObiIj/eENMhLWWGkRn5Jq
HmASGchFuOjS/RYwi0jGnDX9TgoRG9tnJlVlcxnEwW6wSzhM1TE7x/yaPNn6kn0a
cHDRT43/l7zKc2TyRzjZVO4A3qpsbQ0w4Rzw3yB+BezHbc68jOXeDcqZK4GQjIH5
RTa4BQ3C5G1CafXa3fEv08AWp39K2R09yiVjMxymsJh0+MoQH9hq/ja+NYCAHetN
6LLAprP2GzdIzkbl7E1bvrHCPTd/w8vVy/qctGau30XabvjXfin34C75j1iLynED
tniLyru+YWyn2rs+ITugUIdjI7K1naSMt5hhKp5Y4OQkiOkkfDy51yb7nx2VtDWI
E2Oge2W2cV1NLZ+bfeiazcm4soRI84AoLEL7ed2wUi5lGeJLq9ltOM5qavYSrI4m
ScykbqJpgtamxBVm869XVaANGeioJmt4/UlnynZIdKgQeefu8II8gT5ufrjM2VKP
wn1R53C0jLadgJdnFLF9CePKFAdcrC4eLll6dB1t7+451Mu7Oo6ZU+H7usocU8iR
AUDssawlxTQrfPTrb6600WNvWhpCFJcbEiUajXz5B4oAcWyLiHhzxpifqzK/Z3V8
kl0ELakC0MgYTuMOqD2lzvtFAqDZUGCdmGB9N0UxttPpJcjzZe0eyzO+3iY26v7a
GTZF+m20C1OQU+KjG9Ml/wAPQMWX9Ujl91IY33vndVoT3CWOHNBuByDOnD0X98AL
eF/pqm10t9GM3WXB/+5TsuHTG/Qe4w3FLYSoSNcOWP+69KjT8eIRtNli5eXiAk3a
etv5WI/98KOyOIqn1oCQ0//XxZk6ACjJLaTZrGG+V9KqMW4VTiGGyQw+lGXnZs+e
ox1ih+bgNo7afvCT733cSbEOBOrxc12wSFPPIK29AW6Jr65zI4p5/8tIXf49kqQy
pflmceXh80EE/kJjXyu6noqAI+B0Ts5lePU6gC2ymZUPRElCY28Y/AWReRXt6Wig
BrpOfRFnBfDTZZ3apDu6klGm+byz/R7teC32Ph8IEXmlO19DtJdTRpMnub732YCH
hKMBEpvfc6XP4u19V+AhArxSEIdht/O9rgKQDd76w51TDNQFdxcmcAC8QWjZHux4
ZHjBjmo1U1PJVidl+jXG2QwT88ov/Re8Zpp2hnSUS9Noxxs530BBKPcRaQkA05gf
0loLqxQVx1++kOYjwFW0AbUXPoM76IEU6OJbWEILhTqKUhmnLBzuSlv2X+4fGjZY
Aa8I23wrLa3sL6vSRkPAi0m5CSFojFJZ8dFqoackg4EegPS3D613DpcxWcnCQm8i
Diq2LxFA+tIvNL046WtL/StUNyhZaAgWYxu0A33LS7MpIwzn/lneN4Y6nO+NeSEJ
xmOpA0+NT7RTk2cMGJnQ1Ckb4BxYfi46Gx80qRzbjQY5lWvKalKmqjK2TOMs9mR9
taqTNBxdbdLYxV/1sVTdCRTaRFsMYfvpdKCkws09ftsfum8BXpbMCWRDYvaCLM+V
znJGvDtL8OQp4EVWCTNq3JCllQFta+eutsS+kvvM7blpOstiZw1GYENtAVZ/MaOA
b76vDcKrK4TrvAVua0h/2AsqCSQjpHTCWYf+si3C4zQjzuHCK72lIgAq3BA93P2H
5LgfSGnKghy1ebeIYp7WdyUquvUjj1MqoztxByjvx9IoF/7o7O1ffH9pVA3wNQMo
sa5aPsL27C+Cn4EXQ/dzbmvxdBOws8FLPxVuP2SflCXhQzfu88Cu6O21ze+LhUp/
68rhkGQDvVeO7URezRz5eRkD6BAxAHWPuT1/7cqOKjdvE4zJ3//1orhHfqHhF75N
GZ5JqmO8pgYWAVhHtdmItFlxQGe5Y227d40Vmg15a50XrXkwepY9yffZMF6uRcoo
CigS65kpLK3zdQVU+UpVg8UQ67hAALCe563ZBawIy6dqXf8M7AsRusXSxuHopstJ
lb6Yq8acdM5RKC0BZJavO/5rF7uZCd+xD2BYJ1ujOsTMGpaU0dzgg7Sdgsm5/E5I
gmG7f5yMlD2xam6Knui1f9y6Nf8RXXoCPJjE6kmV1w8HdcpoRK6ayAzNyfjdvSf6
i+sD87U2euXBsc4UowDkemD8W8c9gYsxgHX7XwVQgiclvjhVoDtkEso0Q0i3vrZr
/3lgCN04r0hvJ0D3/Lrd0fsWJ/TR9L4KM4I2vD9lWTMeSUw1nKlJdk0ecP/fd9Zt
vrcqZXqmEtLiXwUtcbtmZv1ciOH8fNGazyIs60wHlgHRKX4wd8gp5DpDBVDUulGF
zQNtfsnT6GAVSVNKApt5ETI7OZkOTXWOHUTSQSz1Etrop0lFLRNdlHK+RLIKxEsP
HgWcmF6wTGSNk8Qm6sKDu46lomEanFZ/nVwiOrgdD7XsgzRIJuO/dD2TBdRMf/cr
ki+ehAfy93uoZf89MswD6KjpIh0xCo0Qe7KVmbOPxsehX9C+pGBfd+XfsHiZiW4t
rPTPRRovZZYOGUSTGXCRP5puHmAUIt8j2dr758DxGjIRS+1cyK093BWF3oIMahHw
ybFtiKN1dkD5E+3/pnmNLsvgjKCUvuSwdUq4kmoK8DW1/jqlgzleqgqNhO0y3Zn9
o9hD7okQpnC9nmx7e0uTq9Aek0NbsM/pgabNfXRAzO6oh7CFq3GeuzDTuFdnjs5G
rcyWdGnQOvswSyHlZI++g70dQACRJuuRcG+dNrnDeoU9LfX4Q6cAIQ282Wpb984f
XSeP3QRq6Pe+Mgt7+pFo5LZ7LrI21m78LspNdIHVFRldRSptJLF+Crjp5E2m+Xdm
v/I1cVyAGoju4e02a946I2tws4IJAAD9i5e64+cf8Mve05pO8AZLsIP+p89e+0G5
8omx/eeOZ4W+x0x9TD1pqeHj1xZnMiyqU9+JiBS8xz9yxC6q4tksY5iJ1sZwnJiE
MRE7DVz4d2YHYa8Pd92WGiav+yaAr+R5MR0ACv2zaWf3CkQCwu0ccqILciOita8B
hEcJpVv/yUPfOXV71Ttagd9la6Kl7uwXDX4l+y83Xc72MRV72urno9qKqZXSv5BN
qg3frgC6tulJ4/eqhL6yFpVjFJlwaIi4qWzP9Ut0HCuAT+K3+eTn0T+kF80n/Agz
1VecRONLM+Ss7ghX61Rkkkkj1fLWze1pEAtLem0PYyDiX6aPodW/oEMOohi/JR/g
T0PYCKimwWPiM+avaVafxco8V1okeghEIwX+TPVItyZB8GoIrMYv9iv/hevh1sxo
ROny85KdHJbEoN0rztUIaN4TP4K+E1y/uoIjajtI9yjke0Yoce74VDVyayHRiCD0
4XdtppIqHZEb/DsjF9rMao+gV6Ef3qZkzjNEaHjgTDGot7bVgiqgtPgNngpj002/
/0DcPX9NWniOMwc/CpQ6+IIqw9D3T/nQiShQaonGifjTlYPsFo2s8HsUorUFkErO
+dRX/d+DpYpjcTR++2MoC+OpQijWqrsnBmVH5vrPhyjuJlsNbGaQXZGFWcgwJTOW
7LRGREb4Aluh5Cp6BTIKAQDhzDYqF4/NP62rkvmv/63RPkuSGu2G0pxKUaSE+jAR
uLqmY+SeHvHlyIdmiJLd2rLNhCkOh7uJGU4Kg7NAjzCG9foQ5DSEKJLtfZ1bk7BF
jDR/3ZPdRT34Cr93IWdXHCt5/A01uI4mumWHXlnw+nbtfp6IbL8Dq3Nn4dmq3UD+
OAEjP0leIxexIho9r/MfQug/ZlHokoYx2xJXmEMroQidmEwXYXOFIZQWQ2nAw2xn
5s3hGh0sw6DFNV8aBTlNHR19k4WjoQI9bosBbEbI/XEPJOI4NSJjqEJfNUZqdGPK
TDZCOM1TJeFCoKomD1FOK3W1eWlaDyaVbeLgPy4lYC5+Zv+Zew7beBxee0tfuLFZ
iPxGrVIsIrPCvZecZgiYYSnQqFnRy4IVxQyFTcq2HE6S9Y/UUCyF3EqxqIh9cqYp
xK8Xe255t+zR0uPIB4xs3amXlt/1qXQ+Lt2gC6A27n1P02aqsnVrfPJStU3Ks3+i
4RPCIN/T23R79A+XKwv+8JhDl6ljIr66LmBAGr5tozlifz3CpulIVkBFDBJvica4
q8imuUWkY3rtTbD1DLI++5qVoVoI0/DvOwj/RbjI6eNWEkqGfkGdygae3W9KSMdi
OY8c7JrI1pctWibsQZflPUWv8L70E/+0Ax1ARc2XgB/t+trl94K9DQbCqYQQxhEI
DPt0YlUyIBlE2xJAHZRag0DB3sFzUaRJOZa/WzCq4XjBWcPpV7ozDRsnTFVOAako
lmHs/ML8IGWzWM6WllIraVGXCcpv0LRswVdObVDfaJZxcbj38ETDzFNIxq7C/Dik
9BbY/WWKoubPgmwRAnOt57h/WY8HhDfbU5irCkkWpth4ZRhMhV6eSRWOQHQl/ax6
zLgizCxYW/DHMiGPy+zKQHXlhmqycb/Qxz/eitMJoIyLj4uvGcPDsMm0uFa1h1OL
uh00EbqrBIinpNm5IEe1VOXd3Ot/98ECqx7UOnGUJ4FOMmXxELFUn4LfhPSQ9aYI
0cIwrzsGGQ+xTDphlG25WyW5gOrhLhgW45Up2hRdWh523xbhtU0TYaR1nUfKbITI
38vd5yShxNbeuhr8kyCJxyfDEvrOm8uxM89dOLdATEf54Zz7kEwKAZnOlo6nTXjd
4kxhUBhpBuiO/fHSDGJ4cQ2BNN49GyhSSPo80R8CKAy3DLGpzLfdE2PIht/6vQin
qcfegzHsPHU0KaWtb5VfHEkSf33QHm3PLI7IEHm7Fdjwncs519Eo1r7g0fYHD2Zo
Dx13rhIZc94wNCo/m6kYXsvaEl+I6A/TjIlaXYqdyu1Rxy2HnM7LanHC9Gl2Z0z7
aoi95jK2PD28DYeJvNGQNmNTJtmXjpZVNtse7QrYeWOTb9N270HJkIB0kPwRn34R
SQp86rjr8QrLm9nqlWFo0+aLdblrqKImv3TNpplTFFzz5vClVntgv50eyaqWnlTh
Dp/R7e8ZrETJtOAfRdSMRNNG6f1xgQJrpTDloAhaZV2lzChlJWbJYaliP7DElIcH
iieURGAAC0puGtP7s8/bmRCN4EUt/d98dCZ/i5MJK8Tlx6pJl2wMZ+WV02PETBiB
QohAc84YgPJGQj6DwWBOHP2HQePDIf61zcirlFdlkzYDGLrNdFfLWlGWVP8niAdz
5aUWg195a3A7y63ZqmkaYj5mByMxAarBKzbN9BSPo8zbakjSwBsWleVGGpIPUEEJ
LSgpf1X7j54wJq1baOSbJ81BhdX/g7nwvK0o8BB8QsIhLa1n4mP2vwVGrX8Yx9kl
W4ctWddrLTOX2WzHBiwY6FffEWTf7moXXblBHwf1rZFL5ozz5GKRW0ZDVbzPSMWr
f6LId1y+Oo1bHgk90rGWyM0lxKY+PtQBamIugaWT/qjbsu2RLTvo2FZjSvhNkN6H
8rKv77YNh23U4FlBGK+zIrh9mq/4F/qlpo3GH3klY63NxWVy6TZz7lpIWCJGs80R
DqV52wzUIsbUapM9PtWxu949AdOGxNph+mBUq/bR/Cxd0Jb9AEdjyzVlJ8exiRvf
yyJHQUNDPyKQXvgbGgJ+hlvFNXbxDmErJZz3GAbsE4xusMdzrMFxpdHE3NH4Tjoi
TAVKVpnbCUK1gOFZp0+Et8bhRd1eV01LEnUMPwBYaCsUQccRL+MVaKW9UiPOyNR8
zwFSeaZEUA+G7AIIX141eizfQhxYRcIdjxdm+Q4RDxdRwyfAtIt+xTRnSXQ4i5dw
qELGMudeMIFYXiBxnqN89JAmDhI3ABaesrqL1YHNNkfRpAjcAT7qTtUmJXg4nnUb
Mk/bAb6sziikUlwk1VQdpcUiImmhw8FLJYEDNCX0PzPnb6izAZVde0GXInOCZChS
OiQeqSQwdtup4S2dF3/lZEkinvyZsFa4lvB1TLV+NnIRYsptmxbQBSBDd0lB7h2G
ZbUikANZRxvpbP+LfuKDvkjYSuhoSz5YybrZPwTwkwzvJfH/908GraxoZfyNWN+f
957eDUAo41vwJtGhlYVG+PVmIJiGS8CPa/QYR3oVxXCq0o4xSciY50M+1l6OJ31o
twahPa5RtUi2CKJ3czMbwYwpyaLU7olaHgrB6eNOgy5Nr6VTSIihy1tMO49ygA4F
4HhdcwKHpFDnPf7B2jh86jlCWmuoHte3modQyaWyYG5393qKyXVO75bVfSj1ggOE
cmRAgFgXD6Ah2QIx2lzDopfFqWhX4o47xhc8vc3WrzE4AZAO5B4BjjvCV2jKWyrs
I83hruuBY7rrZgP00KJWRpWZLX+XmRtwd7I54oU4UYNy25g4rThjcRZxDA+eDSLq
Z4l2qgAgQAk6M0ycG6UbY0ObrXf7mjpcyC2rAmAVzr47AdSIg1jN4waFLrGATcXf
3WeXFLVvsaKR6J5F0M1f5QAK4QXUMkiwrol6ZD652CYh+0oaFhsUbstscjyM0cvn
3ybqKI+D3Inw8qDmHqifhzNePGTXsz3J4cfhCbuqaRJvd8Ye/IEQlL85WaaUsXPX
mMDSvwgEL9juY9x3BmGCI1znRLr1eCEKfDMSeNbHyG1ThBlEIeJoow6NLrzWAe/L
3uejO00UFrIF0nUjhbw+TwO5EPKPyDZVJKy49TJaB4p4SPCgHCTuvqY3dRVj98Ot
Yu9GrsvEio4RJNgicq6wtQnf+2wUs7GmoinCirEZIxa/UOO6M/FSHzq+fsmkwKit
qFmAyu7vwisXG8AjFHwP5LsrET1saTcb8yGeBkxYHwr3QkG+VhNL9xKdUBV06TV7
ZBhvfGYqV7zmA/hcgMTvZd9BXL8uadGXQZyFpKeyx67DGEM7x2dfRyA2YB6/I4oM
KonLGGe5ktkZIXKg6QmGe1FaUxxgLtpi0YSOPpFTt7QUH3YIBtsG2uRV40tOcSzX
w+kyyJHmL3QRPsfkan0URd1owi/CZTQbOrONuajhufoU5x39tsFuGStZIl9g11ff
3b02Mvj+Fd3gcM0kljFPdR12cpooTpcoBh6XoMTp4X3/qPULcLvKPR+9iVak8s2U
6iSQqlTOD0izc1MBSp7rWJvLcltOUwTJ2dn6NYz8TFwm++xRDIF/mCe0ak6+tGer
xwdPfvaUaqJtHuDkAomdpOL6XuqSwgKjAABHiLoW9COKGewdHkw5doc+rUszfTdQ
1S0i3qsPaD/wadYwdrzvbmS7oNIOoyPb4LJZ5LsHK2qOkYOBpXl9PbZmXzwXPJTl
fXspH62yo2ihBLFEndRRXCaa4YsoNwZgRb4AhvpLz6C7AUdvIcIy5zPsrSQdsFsO
S/UKE7xueHXYu4JUMjvEWCU1DVMj3cgwqFiuKWKjwNLdQPQSRdgtxYBL+rHVIdX5
BRGoEKOfJJZ6MX9F25q26ijlzyHzXQidMalMuLkl5vWnBLlZ3ycnBIxuylbkwD2F
u+3nCq4xX5pMb/3jdHi5mVQQ+ByPhljDrzgm4zZsuXRs7TLUsgwR5ojLpEh5L0iK
AZPE9pfNxKzsEziPMkB9tBTuCAwPm5ouqg+OhcLuKovb46s7a3L4+qzY3rNpNdUO
cQv5rtLqlBEgG+nfgikyQ6BxqMb8DP11yA2hDhD5eCD9un94X1I3UeZqvl3xJXyb
+9D2qlyalCVS8TIBBiNE+l6v9tkfU/RP/UCsx9iFXLKYmhRQRJ48fBwOcZNcmUTw
cz9nuHQGjf9Og8abf0vbL1XF2uVtat1ax6nbfdtIORkVyeGXQPfmpy3GFQucDxRv
=======
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
DyUmSSJKy9uR92lovAin2loE39uLBCDwM0Icz/D/LOXjDRZhmiAqq0Cmj+OdSIWk
x53eFyFiQYmjkEIXP7xM44iSM+K38ZCq4wEOj63Uk49RcjKLFCwI9THnPGxoQN8I
zkN9s3NgkLW5wFyYWypJB50KZulMfpWGUPJaXTMIQxyICqOSCIK/oxbNlxeAgtyC
Pcw2uhL0izED861fPI0IycszuQag3vnERKV1X4idEkv3TxktPXRQAg4Z++RplyhH
rvPmhSKvhbZNNAzgiVes5uEG6pLXb9wEa0TtBJiq54C4zSi7yFsp6GySHusix9wh
NOO6dhpWJ1NoDEFEBYIcAAANTjNzBwMxegd8C5Ye8vz3z8IQALagu8S0hyHT5jZo
xjiJgEfDL5Qi/ddPD86hpJZPq5V3SgoxO5dxMzxs824NzS/LnGnRAy2gZQW2+GvG
beDJNJxU/WdTCIgo9gO82cehaKdgn16EoJkkaeTgEn4gfZQldyU6c/C7csgpOWxT
wzbl8LNF3J4NLOnq3uPTg5tdjBJ7fXTYpBbNG635zDIWmOG2BY0QF5jkziBFrpAR
X175uTl3Yf4VvQhuZpByqfKqOi40ftf1tW5AEa4SYjQqqCxvuZE55h22BqS0wUZH
qV4BvioUtpBttBR8L1OcWqrWyOqgiUkpeloIjmGvsUGvoCCSmfNTASBYjv9oMjwk
UBzW6qfm6ZdQtzK18Un+VpwQH2oegVSkAgQLNiyB4o4NPJZf74D8xlt399ZZZT3h
1EkeFiSsMr87PxbEaIRiVnEl1GfozobceIbwJIcWs1LMOHyXG2dzNXyZhNAfzmaz
0U6YbFkkxdPs6DgwIPbnewgj8jLutSOAkF0cFAcBai2kqa9ojhtm7W0lET442sSp
R5tutB4ZqBQ6BmEpsHo/KsYPl4u9WzaEiDWmGCWXXWudol3lo4xMsfAXLOkBbaWP
uCoa74/4binQsFc3nXhabveHOwWs24Oq6yTapo76o2J1qTma2vsKEEPBPTTzAsfY
N27Q//sPpbPtAgBgTYFPaNRpl2pyLnO8Y8iocK4YIpqxjXnFSSqNbtRi1bLchGhx
OB6lpawL4bedZ/I99X9RuL90+9bprxyutJOtgqnYnJ32CtNDUH8JesYX0ISPw4Rc
Fsr+YtYdc1b+dybFzdAujrzEv4Iud2B0Byz60pdTC4iaBpIJgTqCnY/7n+lpjP7t
+438V/K4EtlkLrMHgs1Sej7c++W2EUfh5wa2HdaPfk9MUljKIR+CJd5dtcrcUnKX
xEM3gGfM6whYqmhocjB/yxzyw9RgCZonP69sW5aInhuL/c5HeBwIsul8HvMsLMqs
D+zgswiReQbR1R2XJnzXTitd2NGYj3iN/Jggk4uYnBWdEH4ayhX8Ix3ewynGOaTp
x6Flsn8S7Dik16FvGp1AWFw1eRZjfDPSOwiDCkWM+GPGrdX0hqZjKhZTCD9UP7/w
GTQgcqBtTGv90a53aEXIchY+kRGjudgApHllIbJLZFM+VJD/ixzp0zs0g7rlX8DX
fIqk4b1vcCRc44jX/orFHZwbCO1gaKlP1bLDVaeQrBOEz0VgtGVDNJh9hgfOfNx3
ngqkXDjVXqrk2NmFgvPJjYxt6ba7bx+/5mQHojHqjVXpAI7QHI/gDotpD1hRTHX+
7qI/OJJUJjqnSRNC+S2wVPhBliQVgU1/Woxkb8K8SU3ykRP8x1aP6kzShlYwNYmO
af4MKdXEp0/ghASelH52lC0vjpLOL7Vj+eUOjfj8awhT0nExcLr2PgCIzeRgulz0
YRj+2y5MhCa7SQZFP6RQx1wt1uGQR/qpcQ9+yBahyFGKF43ngTVyW56ODhJ9T1ch
vJQCJT4xpKzuyQpOHD00nGpZk9tY8b0GnCp2k9zPCzTFNr/EE7kzIbIloWP02Yq/
LkriRMDwz4g9goSgharGbK8VUd8ZX6wCdqubQzHmaVUBtoP+Eo62Fzl6/FjcxPRw
SHPpDRULlX6fC7giVbo3mWIcSqVWlxw50N7PzdAw1aKbOZLLcOjINs8J/CfVCvoQ
3ElABdePiZQU10KyDX5MKQj3iA1FQREQqGnbHjK/VF06RQ188RADkv0eJN75lRbD
/q3d0ZgU02SDcVfAhm1+SNsqy4eeoeQis0FknK9uvbiIEERrOd5es4wY13wJ8I0Z
VxVImC/JrfTM6xmRmtBEfrFsoer0ygVM1LINm53fyvHdqVTiEw76CGcM3RxIMUQI
ooH3Tv4GfoHb6Sww3lbam+FiJ7gRVJHiRxwT3IW/NhvOhsyX3uymTbqNxBFZfiIM
/CgA4ALCOQc6wr+TeBzmaBdGfyPXeHwRAj7NkQgh0e7E3V6kW8IKkGrcAJlAoGLP
Y1JU1g8ZrgVR8cwBxgaEBAc/d3MuVVhJmEeiLD7nj3tMuncEbtORduoEtzpZiw/1
xOXlf7aCh4Y2WZuJ5IorfzKWNLWt+sI5JM2WfXkPFYKhfYPnejdCdfWESFY8FKF7
r7GfBnqDEVfBuD3Em2smLqk0F2M4TElgcAQU9Y2b/Z1UW1B5X3IKkm5gF+tFC5eJ
3WAJL6ASkljNRFAWuH+F2uXQencQoG5bBnV1xmaRTyN50ydSDDSWOzOEouTwa1NS
76gUupy2QDDVcLHeZdQjsrb8TVPEnfvVkssRpmhMgu6bja7qwW5GWssNfns0wtAi
u8dsCQQmT247KYlYc1aX5YXWDNHSj2WRKxrXvrjBPi+2QnHl52n5xi6gjPpDsTES
7dcFEiQ9w3LTILc/RH6u37uwGOw50MJgo/ArWsZxQIB6d1ZwPjWBU5BNha6JVnY1
wLK4JD6gY/GZiOU7ufYBpAaaM+DQFifEFEaa0zjTfClRcwhXjSrImY8UoTxES8uW
OXWGoP3/57HAbMEVNdNJWrFOKy9GA1+fl7BuE0UkQzhShjBCPGMZCqc4B/o4MPXL
mAU0BREMHAUQrkQxxjsIo/pWIFMB7meTeE/y5TVG2OxfLMV/KPgJSgl/Dkuhryhp
S1X+ktC9Wq348BwMxmWRoFf20EwQPsHfJzFFClWHg+MtsWHeooclgVr11iu2VrCk
8LA2+1QiqwgczyGDb0sZuL2FEudlM507NAyf4SE0KsdkhLR94C1k4G5mMVztuSUR
ic4Iairjbw0ICbJVr/+rgB2ihyedG8hld177gake7Fy+sNAZg4d+MmvSH9/Jibk7
cuf7fCjqJDmWQgrAHXwRe1DWpcGvuFBfy8SLetZw0LHdPhY7mo161y6aIO+9nvgd
YsVG5vPRNtCAcpMFp5Dyv1AwoIOGB2bnSKWHZUuDRIC9QfUGrnu/JasP+QP8QRsB
Pet1FaQrSPoX3vW1R2bGOuI+WQyqxleK4s0iq1uma9ZOj0gApCoJxcMzxzVl7rJa
jnvNKQiMqT2NovKUUHyhXLPmi8onefRKx4VktXCOKjRjYykCeUXf9+jCn0OofNGP
gB4bi8lDQEWU+oEeE4e84m3Vn3GnAvsc5eLyuEnl8vtvbhgHAiHhI5x8rabnUiea
7pOWS5pSlMA3xg6jUorM26zzTUgiqAeVGtv+BS7/t2lMYYJLq2o40Utu5SDwPqGW
a9lJfu8GKNJAJXQlQP/lXTU+4MfhJTmHQGw2QiY+r++/GThlCrmAOGVWXANyxP/L
XPg0xacfZ87/d6HASkBqBL8heOZMuEyakx9KNb6ivkADwkcU+1RYn9TooQ8HJdCA
yMkak7GZLeZInJWLbARLxBItrJSCb5FMpvT/D9YGkppOt5+IPIFrLaNL7/Fp6obJ
DVAlmbeL1P0nY3xjbQzu9y5Yee59iN1dLsNXLyff11zoYqSscnbRmIsb36uI+f5x
3/bk2dxLm5BvH3/DiuCvTXmT49j+wvd1XDj8IRvv+wPNMcwDmly4dvrwP5ZbKqii
WqOIUeR3OtQl+OgtbpZxl1VZQvTzGXhcFMA9RbJh3JdeKg6077fyi6ehf1Qrh3a/
XQilAyGThh4eM/+LOcKYTA14VhKmikRnifLINWFsYeISNAn79Q2h+uqG2rN2zp8D
X9yHhbw42GnCOO2tMO6E2npnbJEd/AybtIj1hVFrChkvv0+0JZ99vOMUxtCfWHy2
AnjOkCJm9hwkPF091v+6+zCKuiyYGw0UBZoc2jcI2lqWkncDla72tudZaqP8Dne9
KHuGtCyBgCun5M3Sgs/U6xHuEELUdx8IfZuwX3x0HMXlHA086Qw7acZLKOM8OeiX
mK7BMsacYPPoUQT4gByEO7VQTGMLzj+iqeLBKM2DKRBEFWzdxWHn/e3uHBRWK6pI
mBToeVt0gGSA1kI5KeuyHYfkbISU9uTn4tY+V/8kQGhdfa2/LN6j1SJRifjTNtC4
F2ClL8zDgx/obzhpdk859WhGoEPRcavYDzgyVMpcfosIzemMtbsqnxV+4Nv81EsZ
JwUeAyuaV8HRgOjB4SW4phWhyKhUaY52dIAxfGw5oIPLQFOlYjY7a3UQlqjoPtOe
xMdrDZomDI1h5botjR+nfGzEiYHcu5PrDzoWbLprGrEzWnvaE/NkXoSfuwweQr2A
wg+9djwijebOhDDK5At8H5A1KTqL5WdfvePfO9MMvk9FgxR2mbzobASetLMBGycG
9k7TGRAshL/N+cHPSLCIre/fWE2ur4bXbjBVZpqDqLdipTz/2sG5i+tTS+zYBbp0
ydExTjDRCuj2c3oZai5O7hCIGQzzv6Sg0Y4LwWNVA/mskqDEdsEAmyHSPE2iu1Pe
KHNgG7QrmQFhkb3GlcEPU9dthbQTIowWSzhSwqisVPqGd1/6CSs5xm3hITWz7Srw
kIZrxegBdJy8ikaoE8t5lbFhtW1anBG0O6JM99K4qSOrAqqXKqU/RRrcig+yHjWa
0VsoMucoS2OXBqnt6IvAHLumIT7h2g4nzzhffiY+QlngUd5spZB6fuVMyH49O5IB
91pc3I76JvpIN1JfgFYKIK7nt/6zYBKluucA4HbU9Qe7WQ/3br9WieREGiZ9JdQt
0OIEYGrtzf4wIAmTs5AjaJyGS8rc3Rbw8rHPpVBG0MnhsnddlwK2rgFnyNA8tiBW
zvJGh0BgMs+sTCq5MUjR/R3cbEfdN2HPc661pE9VZMf59510FQmYBBN5zRzACvAc
LNorbFyfgAxLJo4ccMR0e93s/Uy9Zk8+4afS+d3AD6A+uqjGtcG14V36rHpWNgOu
C9MnqOxGu7Cvj5yuxBhlr4laHur7VyTthyv5x/yhw7FxFKG1B7n85nUes0iFFhkM
S3ygO6ZlKLAiHiEwJrNzxZ2ROZDBw2KeXnifXyaKB5jjVpWd9u1YxhzdsXNv30rz
otlRd/UIh0hdhFg1GkTQ/qScQRZSZlb5wjmSF46SQnqQf5mqXw6sx7u5oOJ0gCV3
2v2nbBBSCpvad1tenR0ya1f/mKuIHNwkIKe5YwjGMZcJZrMVZxu/mIKpNnRQdsrH
9nJIFtTIDyZCoZaTkxiOCH491OQkod+r9U3OxvweZC688nhF6g9mI4BQA0gdq5Ml
zmgdKSRRHjeIvSzCpq3OIHFiJ70q07cHD4agQE1VMphQ39UWmED5GZtWQxVaSAwt
7yAtJTo12/nWaeiEcfFq6GJI50SZ+M6jPxi81SiK3TdVV6atRYKlf+BixxlPZA8H
+/M71Xrio0N3E2GhcR3RqoEwzb9J3acyXPDZIEAyGQX3qUqw2FWRKW7KXrFIR5Kh
Go2d7B2BinswjvJtq8YuFvkSD5cYKh6w82iCkbt9OHdPk+eM5R/8sxDry3FYLsIU
pfV/1ZKKIIYX11PZ2H+pvb7VAnC3vKdOmR07nwg/K17Uj5AuU+v9hMYt1S4c/rHl
FEUstz3wD4/QEPjFPLKbyTmDDNc9PBLDTQPIz98KG0EM2lGRuc0qstv2P9tDbCmS
rkc0zMJFMXgrqnvxhrvGoCabL43aXFPMvqfGFjDWxtfDYnBOR9fOcYNvjdUTdhA+
0BdxiK86Lurz6O4SiiD87w/JxPie1rWdxIC5ImWj1p6adCc28fmIeFZuL9QlXsem
TsVBcuea/y7G9q4WL54Uk0SaAPQCOlJsHe+/m7ZgokV1Ad9LhYBcNCRISOhnewLO
zBJzNcg+1J06NmJG1S5mH5cYq+qtgHssP7/9Fq5Tm9PdCfNaZiOLes4eftBza4bO
GT3JR+pjdybuCGr9g5rh7/dOfUNzUMrElFW2mmYnpgjstpN1PwOvBNQGakJQQuQ5
okGuar+CveessBYc01oLe9sR1+qOr57EhPOazr0/m5aJPEJbV9HIAJlsz7Uta8Ih
dcAPCmZnYufr6Pgy+RDZMT23G8IGHn82PpwEsdDHv9Z3orhxj2somUOizGdf7l8v
WYbL8IPYKsfrqc+scUrqJOhAuGsyF8K4SQ4Aeu5ogsDcX/Cqz9DW4Gjg9R71iAmg
pbq+7OH/N0BXXdOvu7mJR2tvaX0VB0xttHcpgfxiiEMca+OUMjKzBRpdZt8gYDDs
tgtKg11QcKHwpxVwCJ7rMTNIT2KleWvC6WgBr+hwe895e91zXCgRdEuXrntEIm0r
qpHO/DxEHl6IpsCSuI+dZWrl/F7rP+RhvgkIPF//VUO7ipnQevFS2bFloHFzj8yA
APRmBrrhZLD7STN1hFNDhJ/FZJxDxRI5GF8a41c6KI/QbjeGBZkt1Yw5P0GrBVPv
WmQTNh640eDK7ZcwVv2F0Spzb65T+sq3G2DDGaoIeM7efyph6qCCvBI12cWHsHSW
ahmsg9xd1ZZ78Ef0SvIfuW76qSlaaYkZVef4aE3PIV8mVttOrVA+K71fiZabSLEp
u3i81r8zOX4abpgondrMP4aRICVEIo2ro0baL8LhqzhUahIVtrZxC6qcni2kNU50
kRQFUpGbBNMKuvKXkzUg5qsI0pfwEJCFhj3i1ENGM92GG85YJukRehTbTi8V3L1r
4x1+aLzUyxYBPm+BcWgMsB60IWQu1NtbSWD6tT8+hZHq28Tbe8ERNcHoMS4/Sr0D
4ty8MItk4ZR76igx9UKfJq+vsa6P417YVZlmCH1rTK3YSrOZTtvc1izTUd82uKPA
OOfQollO5fDOYzyxgQlQNRZOwTnlcG700pEyUpqbqzy71A2cnXwJt1d0O3MC613p
NAElxhhSCsUhLVDGbUdmv1S+QVq65psellnAMPKmiV0UpP+WGzJJ9swG7DGhlObw
2Z+2jJSbUrwUantVME45w+Dmr3VO1Sr6dY76kDQYGm5HkVVQE3KAyZ5Uxdni2sxF
IfRNS8WwBrUThwUIDHUKh+IXttg/hkLyzzXburQ7upJpFXwGMCW4EA+++PHrneHv
JbMPGMbjSwLnSu5Yj4qWnkDXqU4K727gUDE2oUiPagRSKbhk4E5liGz5za4RMV+E
6kinaugm8xznwNDSORVR6XdOeb6wjtM6BzW+vFSI6et9C8SwZl2I+qEtQNZgGDKF
N9f30mvZ3IYJO+bg8whn8lQYQAIS1ipbhlIDrte9URgyNXPiycB2B94FppN6YTym
j9g39hDJTsRXUuIihvrZUchvcHCK8+/jhs1jRVHIbCCWC8Lu+UPZ4i3pJwUI7Pra
Ic9UcBqyQNSoPTWYWi89+UHDzfSZMEQjQCYsZkP5LL8JMlA1CCQNsHcQEIfOnlAB
TsCF/YKo/XMo+SCgAHjzMwcenHwcBDD8CGiojQ29dDtE/XrUO0zfpr2dxT9pue3s
ePIG35leh52k03/wAmBaBbyOKRas0ovBsjBr2P9wdhQcCseo/tCHs3PG1cOg8R0G
V1iSTpOu1xx39nczWb8wpgaF3N429cAnHLwg5kw6R1oR5eMhX77EQbE78fSuYkZn
jdRozwL5Q5ZXAzW4sLUtdz6oy0i98cGuk5ufjBVTyAx4QcEzbdtKVo3Efp1euY0S
KSeA4ai84AhPJxFRsAS4PCPBEnerVFMp/VFrPlAZzWKEraQADXUuWixZAkZ+X6sQ
0kJ2TSL0LoPywFP18BglXwAWqnR8L88yfHaU+j1Xa4bX4ah0ZWJ86zW5Kb4qoCYg
2Hg1Ipg6Z7CmBrgJkvZyRkyF5d2yP5Zkp7iFYQhHXwIW74NjfTJs+OvmPVqo9vj1
wFuC2i2IMuh8NmrcnqNsUKIqVvPv1h75ezQXDR9XGYHUw9Oq9fRL8XPJp9EPowTR
8h4fFFZfFnUWnbxJiW3tesbzvPE947mFNKg/GWPcGwOB2PT1ENHNiU1gBaTL3K6/
z2T+tgE7VnUHFKQ1QIppWOY207PiCFNWEr+NvayrLRT7J1e8f683MBYXSkcdlFap
6ttgIFSk+7k4hPb3l2Q1A0vtdV8NnOKrk/0zbQtg3e1x3O80ZlKrm9eeCfcNZeI2
ljCGf3GPI+0lPCuKgNAuQ4fJsWMlmRokcfSkJIrnF75H51QsMdf1Xjo1zI9xzYdw
WdeUmzDDiUv5KPNzcI5sCehuKV5dVhmkOaLH/HSN/4oINsgll3Gz9AKprVd6fWpK
kbcyGpVR8P2OmIasDWtjNBNhDFHuq0P98PQrF49bvHDycF7DstG2zjKxeo+itGgD
vvXxVGevw3ZGaKWB/6p5yKUc9NtWLBsc0N6SrP5JretzYl+7LAlntKfZvWLYd5nR
Oo4bkkGnDNrNYJoQvM+aMVqzCnX1KJ2QavENOwcAtw5mEwG9nQW99IIiie7pkIQF
MnKrkZJiHioklFdfgmaQYvKVL6zjiX+Hq+EVLw3cpYdKfxXUfFzfV3wNp9ATHoP0
jn2fL42UBt0i3xx4LAPl4U4/kiW9l3Iy5Yw92aJrxvoQzgBAjKPk9utW8GAjwPCt
ZyWsHIkOQyH+84JCfhn48Nb5T37250ElWlrAKqej9guze5VguiFq+fs6M6eFBGs+
o/JKkhYBQaA2fpQaayOJ/exFGuglAfFKNV1DH3FLzVmB8b6Ux4lSBCw0WHoByrcC
ChRLm6FIFKB8Ri7PuTaX9QA2lpe+lAO+vlIGIrEeXOVi33lcy3bcCUbCeUuv3HqJ
nRP5/78lgVp5PSMf1Vi6Csjl3vq3OyGyHHThGDoYdIF9AHjKFsCqjNp6ihcbI9uS
r1D7gHGnzQGvgbd/2CTCFx6jFLgUHQAuazndAlqA2Ww4vv8/k3fcPlNmWvDXbjXj
n4DlJbU4R5OivUvpElkJnAhkwUIBx9ILTQLEGJeaVnBZYRWJywLwZLs+OjzYq1uY
aM+eQPSadfqSzGcabyml47QTiV9QIQnsmNJKEtPBVfBvnEuKm8dQpmVBCDIeAGsz
IyG8BVqhOjdi0w1xMws3G4cncTgFxPxEQivhej1cqAYTQbKdtWxlvNk/cK+d94rn
f784uy/qmpi9QQoajoz6vhkfPV9OfelPicYurHlfG/YBkIIAlEH9k0f4vBroTbtr
8vUsNPAHMbwo7p0ZMsaG/OqStz7RQfycT5JSLmiuUkse4LaNuRFswbNo6Gg/GC3e
4R7w2Rli6bBiKYCOhH5ChI4xhyFzsvf60kaVfEGpaYKd8Av+F7nGWovV4ZxZ7qpD
+wDGQxmLsxc3hZvF9kQxnGEFXU4+tGOLb/O/wdSQpmETpbb7Igk3KqL+g6h6oC/c
4CpaYimWGOE1mhCApt6toq5t2aaApOZJMysQ2FohJM6u/AOmREm8KfqbBSfe7EgQ
EH2n5uL1M9GCsilnaDpdpYrQEJuYZ3dRHmwje3mhmJUig7wpJvMLOZMB05Gtwhj2
UqjvvNC96MbCei8Z2CS8z/+3h1+gNaYz9N1r/6tAmtNXhZyO6HydRVs6c78EQJWg
K8LDkO2zajuE3pQNEGSgYJhu5nZbkj351eJeBaWGJp/PSc2W6HDf7NoW2Xl9cODN
LNSHzt/Mg8Ick3lM/GeFfaAGbDkprC8dVNtaNw7gcMpq/sK3GmPXqAxz3zs61t2k
M8M6c7KdVGrdUYJwM89naYUu2d/q9ggJ4QTFmFtwKqPccYFRHQtLCc78TQAnfAi3
A8kCSp+oyqiVflOaL22ORPB6Nm4Y8W0yzjdk++0RjT45s49Cd46xPjuao4hrfexe
+N+wJflVbpn8oIrpTou4GnP+DAgr5LGfd7UNFL5NGf8o4X1A1PgkHA8yH+T5issq
epdmaoAHs0pm6MWmDHIJyDnypDGfX+vNyfo5DG1b/7zEXWtwiqCFqfbflCYlsp9/
CUmp4geznuKYKtI94Lu4/x3xKXU31mRgRrB2DY+z/mlHjBcoj4DY7JxzLARPtoVd
xJ3sIGpqeK90js+6XY8Oo3+Lu1F1/7T0sYDO7bAzsPAw8bqusztY5a2FgMVa9Y5C
Cc9LTOozKaBiU0shvZr//+bsZ+561MmeGapqY3pu+17+klmoNpRlfFOR0ZSVQIRe
7bRxojdn8SIxZv39bbXKTWMfEiqFuiEhTsCT7hYEXxKH/C3m5XlMqfJFZqtenaZX
7OSr7VQytk67sxDnH3anwpn8cu3pX/Z0BxNL7KMwQyjeTQM8Uf4/TSnX1MCpggaD
YkZdyA5J4x13e7LpVyi+e2tr9absI/bbIp3hFiqN1dXQivcbmeDenoJREr6FpW7G
BxjGRjVtqa3X0Qi7TeKYphHjtyp7fNSJ/DKI61EfJIKrlTI10yYXRtya3fhiUiAZ
tuL9RnMDWM5+jyIZsscXRop/WXQRQ87AltlQVDr2+7VM0B08zGf1fNeZSOZ9PqJW
8HIgKN/iV8aqc493+KiwdRVYYjSSgDrnFGGsqWPgZgsO6JQQVBOhn+Qriyz19IVt
6UVlwX/cpZH8yshBc3qcQ7d80ShjZ10v8VCxo36XiHX710fA5okr1YaN2Y7Q3fM0
5pneCLho9I6HulyjIaAbXtKMixDX/Qn5JflxH2XJn7fvXIIxHVyTk+R00nQmt69r
tGu7vDLaBpc60FbWBJ/ayGrHk+DbvLuTuVmpORsNrAy1FfOmKBWVdqQ6a8luEKmP
bMrqVYnH2HevSih8Prjdy7ZwVmHGCkv853b9aWZN8bccZ5jY8zBHfBj3jHDxlnsK
jbpjfn28Hjv/IFIxq/uoBc9IQJnsW16Xf871Z319d6PqcZhM0Ck/hj+cMBgrrXtF
QKtSBkS1oUbBTsJe3N7n8/96uafINuD7LQnCznouEFiX/kXWMn5wvtHEbuu+9/Qm
P2cLJdxAU/QBlApeEew/Z1AtINoAa0JLXjUrM9ZemkkFW9wbdDe1wxVRpxz4laEK
Jh0knnbCjSIEDhMNxqKR9JWxSc6DJ8ML3xgM7dxobc6YhIbqq5iD6rEGicotOWou
9KLi+cDYz3fEgl6GOk06MuIx1Q7UQVaOkSnYHTbuZEzRpa4A0Cjux9HI6c0vlFmY
JSjr/tZ7nkCYkbePG22f5UVei1TsoxGL3FnQVy0KzqQUZSLzrMsSPVOGRZJwG2wa
rSkxqx/MvYMyM0rGfF2tbITZE/xcoVIIboFx/GV0dakyT+Ue2f8yeY+IgUsHQLT5
9rGOgTxSjusfBw892ezRh/h3mqQnw+gyM04xhvUzK+78tEo1ohwiCPGTppbBivN8
sSC4KQzzQs1B38JzPrKFRD9nZjOGhrQhN4I+TiLKIL5Z+VxaCHnTgedk5WHtsimu
i/qH+DdVzHD0TxyPEfFhugBOYY5D6ornemx50SjRGs2d2fq9mOz3JcqXibt7RFwx
XvSzVwfAWRgjVEUY8ii7QnD17YHkpZsGswuIpcBh8cO7QScmkzC8OQ+VkB4iGzuU
44rNEI2fuKHZrFXAOz5BwQ4AR/CFApye61VjJhxoVm5IQXajiK7EdR4jtStgygf3
28/dMcJYjZOLVcqgBchrTM8E678T06OdOhbn+SOqJ1RvsEmQXKtrAmVA2fhWvDPx
bNdtwsgnQdQfV57LBViTpXClzm4HI0NAM+g1g5+91WTSuG4iWTSmiQ6HJ9vrVFYt
DvE5fLtVt8y/o8J7I2T/QS2msml4nByhsYXdaGzyNlosSi051etIjiwHjfLzSag2
Ew/00Dt3hFlmMyaW1Sx1HsJ+lQDmd+qlzRKbpKYlLE7E7CefY5Oz/ee2WBfTyg5U
GX1xWHm54lZnLte8J50acLEEBJNMaxX20OvFakabnNEOXRkw30cnFIplw1AOR8hv
aNO5h+EOYEWXgDekAsG6A5QhmqsBBcKx0pzecfZr7j9xngkrU3twrSdTNWsLcJkY
DAqHqtjp+yETH1CCQG8azsbKz5PZPlV2aMv+VQvMEbaVCWVchgFMcKvJL4tR6Zg1
AOntP9bYPyZLvVyNiAERkBPNiefXiwaH1DX/eeQb6V9XHaMz/NruYtcMsDYJZQC3
WqJwB1cX+GDWG4K4FwmC3zjQD+j08zDRZZ6FIjwwhq5/7kTowMflvh1ewjHJyDzK
VCuLQeG1Cr4yvM5oygubLajWVGq2cKKMSP7EDbazd2EoTazkv1Ux2/jr8d5+vF17
611Ah24kA+wyUc/1seESnQ1E/BeXvB1HR9LVuZ6jYuAaUXiUbIKi+8cVUlIc0dZ4
/w0NWrg2Xv5PB+YNrzW6MZUOGGf0IPPY1H7Pz4XrqNDOcmZA1FHFsN13A67xMypm
U7JjRc6O8Y+q3LXEq7nFCt1IGBOeYfPnWG/k6eNoTfpSwSMkfPdQ2aRXdv4J8wVG
E4RMyJHXDChVn4ZtQvmdDJuf/HKVoavK+yTO2GBnCeA7CR6c9u8ahoIF0nvqW4TY
NLhhveC4/1HphhFxnzyBmSfZaOgrP7KicBTCVFI+YWYXjhNLsM9bPdS8fGzOgJ9v
THy3jeGBZ9hl2xr+lp9FVPosXMo/NJdx2mY1cf5vwahFkySCEmzD1cu6/DUS4DuG
bsLjTQPBqE9U/Xl9N5UvxfWLmIBlFEcixIxJjSrCN/B3BfzHzMdTMU6bsyuVF9Mr
bzh4ewRsk3fJkSiLlZOQ43px0RooXpTxHnOi36uy4kYOKakLfPnpdlJG0d6P8s6W
yzcszBMrcHRR5dY2DxbbP62RJ+csjaDG93LXFbutp0pIjt1rYE8VxVlLXH9VP7ZT
dTBA+BKkKevMrYSXn74OoMOenoRnIFTtOY0Q4Y/ZBJgcfKFIJXxHhlKKsNEcdjh6
yPccqsubl/iaZl6sOFMNRa4Nb93Aw8DbvhNS/SZhSJ1I/7vGCGeubE8je5UZZtlA
0nCOOI2gHWBBgvE2DsS8OLyV4NyL700G5mv8t4sxE3DBjl1pgNsbP4dspla4Gm1m
NIg0ouIC9F5fJC3P4alvBJ6e33ri5pAt+WzWNavz95iBC9QL+LLMKTjckc0ywWqF
Chu2GCAhDU5NEMUITNL69YFib8C9SUp5cvFDDjVRrU5zTGWD2rG3ZScuBSejfRLl
Dd2wVZindljJU++RfWyKwLDB7rCYuijZmqEl2s3hToRCNPVZzHrEgOvtyiQa8rZ9
cfsO/MvzzcTFgm+dCFs5SrO9N+zjLyJC70BYXhGCcZr6lu0QBmDKaMt8945KsmcH
w0oRqBdKTvw5gPyMe1BI69trdQoS2cE25z1mZisyjPz//ky3OH7ziVrIqp2YJXvM
S+GYwDfCX9js2a+HmULnBQ9pq9+0boHZPh5fURF94dzVB1DGxt+e+J5EYc9MPuFG
RTmZxDAHa/Y7N2EaSTaJ8Co3KBiT0ldMVtSicWH6A1e9MobGTBex0lWoT92m9N6m
ad+fdHT/e7QBJTWnnHsqPHv3uRFSrSsdh/ao/NpoEqDpm/P6780w6qQRNVgXH7/T
inTIKZKOahals/8Zprx6H+14lE2y4xOOaMGg8q5FgNlBcmj6SAeURRnikSDYUn3m
bK5OSoBz9z5EfjM+r+Xko/rM2OP0r9Zz/hfbJXAJuX1Luh5vMwqmSueBASuv4DCY
cF0f5SM2OkgNwR0ZopoEIaBqBRH/YbcsI0UYAc6DXZ6ZQZjydWtusAyXSEeVWBCC
r3tUxfGmXUaU1tK+Zo4+DnclokkmjNGI965mjst8FQccWZakX1Xn9+Zutq1ySXRn
7H00jBmDiBuKgD9MuI1M4r09cqhzKnlJERi8BOFOfNMrD8p5wNgydxYKMtLh2Id5
FZ/k8NEyydVzsJZlDi8VjNbiTZJH35KXssXVVxsQ8XesMrdj4xdoj1xdT7J9Tam0
RuCbdDvLD09cAsx67aTG+c4HDa6jQK6+LBKKKEoe93wOeZFDILd3Ctyo3ntt9IUi
6kwTgxqOZ86muKvOeiDWwwHihdvUYE8UMMRWkd9cgs/x19ShBi2QaOYfGxuetiEb
LUXcH5yk4nA38rF69WlLmWVnzWRjoxIXf4KCIKnorv718lpvS592otkjYQHuzarR
FGTTCPHUYk+6lQHRFl5FyHclG6u7EeXsMDnHNHXfnJTbbgOl7y7uNlH4DWBfLU4d
xyig2aIBKiFrrsmMeqsE97/f3rBOOiPqfx7BADYMaM/ozF/HdeBq2hJduyIM8hKA
/jWBqU7oBTQTTgbjnGTWoCLG44nZYEtXLOyzwKT/UN1047Rh6oDYLU8LwuUizpdg
5Tx6qx9r4NKow7M2DZPeLaVI8HAmSn8usYC7/IEsCp/X5YNipokWHA78ytftmqCS
u0ZrhWaxHC0J5aZPimh9c3D2k6osbWbem3b8jw3Um5e2kGlxIxVgeR4QkHAgb9Vo
u8Fx7qouRIqPIAWrqmdYDVxsgJFuffQdEs5+vMUDx6hItDuSGIxBM8rkfTEk2IUm
vEV6/nWy3BZv+qe9MItypsqhePGzPS7y6BfvrBKQuLZiwTub4Kbr9U01SNRzO96p
dqcUj+eBv9TnpvmGI5R666Y98kqgKnchYHKwl+82PTls6Hh21z6wqyrk0ZBKLHYE
wS6u8zUbjfLZ19x9zsDhWRU6VIqfPYmredmazT+WAcYyus5fJgv9J/4rhepWqxXu
Ot1PKMdR3ZPjpv/9LkGRc62arGWsppQ3dGJ2RqxPg08rPaJlgDQ5dDufTMV/R7+n
EuWZ6g/ttH239SMvRIqoIGVAcIULASfk0/LVVSIZg8aY0IXum39i9U4LSxXUXCmr
7RoTOlXqrHNPgJ+/gDbbsDbMjTTQBctRHeahqMU1HUEjDAQE8HF++3/vIvC1LB3t
iOdMtc2KC6wS0E6tfzV2uE9Hqly9N3tEAYgbuWUcizQ3y2frZhDJ56PPb1p1sWEB
Lp9z+oG54n5T9mWnkQM5Oyp3adjLaAa+s6u0fpaXD8xdprpNS7kMhtAlzQZc4mUD
CgowYL+5a/jW5cQVaKkdIKuwE8SaR7F6CvP93bmeTyPRul+gL3MibPqj7EN6RaSf
LbbhDe6SVx+OFSq2ZAxkpcGzE7yUupVvse59UJ3n9otuXI2qZgw+tcZypEEW/QtQ
7opq6Pa+k62hi92u6M4fAa5G8BsXDLMg/ldWqCm0V9CmX8OwU1FWGD/C0/5D6jzY
TKIIbiW80f23hwn6ptBl6brPsX6xvkklmtGEeOeEgzsSEKCJ0WmkTlhjBsF6bEEX
tC0dLbymrqAnrw9UBY9SEjI1f/8j68Cqtj7CEfpZKs6NbiWL8Vlh3WzIqL23fEsA
+3y4B0xaY/FT7xtPijqYlvSeeDUpXpqGOUQP+AEprsTxWFT4PF5tOMmLjjiTbmLk
sUfohW/2BJImf44i2sznGZMivEYYNW4B01dumUErBvVm31x3KiK0Fef+ar7G9pTB
xtz0kidHGnZmyhKpyhsrXWzk6B6GCdyn42nQChcZUPvApvtaWqaLnY3AbzdMpDWf
WpsVjJKc7jGRFa/EVvVG3x1dDVxJG3zSHM76NHCYIzaoeSy2kgH6ISQGKNmjYj1r
JmgVyUPg9faTKnsgUc6z0rNTiybe/ZXuqhO6GVlIKQntApjASj97/hmLAPqahl1p
iw/YVwjDOdOmxaCirdDEA8VhzU0zX5IL8WJFtlssXQQOuapg15AoYd8Ti9IONFg6
QBPMrWPQf9fCdj5AjZCuY9Uo2Cc+H49666nZA30YcKir+U4nCw9rY0ES88i2nERy
FT9a1Qbz1OoYizvkt0EwaN1ERfQJqHgyCQdQTFgakKmvhZlnK26cL0xPBcDkF+Wl
nA7dGo+kRM/rH0IR3J1uyq9GKtDgxZ41KzqiLJZadrbrTsi83YUAVgxbpi7GC//t
L2OAWMj7DW09Obx5LIAI5DoywWFCFKrIXHlOuhVxNgvrIWNGWPiSufWidDqrFOBw
/TKbL4VhTGgFV5uQ2sQzcwenJ1dK1XU3OXPw/nVWHx6RxJmqZTQvm1QFXnTzZpLS
A5RSn99pko8ghCMu9T/u70YDUidF8cujQUxJsIEuz30rUofNA/NjsZzFEwt51ze7
911JrcS3Wb61A7VWiZYPRALfe3y2F782egx/sFaPM3zQYR+i//MvB1DxJhFvxphs
iEkyCyTdEjhgeROIrZNqb/btpqP3FZWhnoByQtEz1JgjAz3BdWQe7Yy+cXH9exiJ
EZ4x8XcRCYocpav+p7ev6FSvQHeSQW7G03HB+QhZndYInSpQ+MbbNrpBwVtCog2U
PNF1YcxA9VcUBFK4F1RCbw4JGGnc6L0MlnFAvpOkx8zSFfxYfwUgzsULkQFn135O
8f4Nm01QJRSGmkym7v440/Lpjc2Fwd7QbmKjJGwiE9XoyzAARZyca9nz4yV2t/ji
Yn/SmyGLYYT7QyVz2PlmHffn8a1ZHxuF4XgwcuKBeGjMrG5LNxE9Wd4SHz9d+Fn/
WbcJVA9jPlTklk9T7/mAiIREm/p2A9SZ8ltTbMFxx5v52TEHO98H4cejmjpi24yd
y+Wb+l3syeciKeBcV8/oYD4+BRAcgQNJludCAvmgTra2raLmeNVtBlI9yy/ggHtw
88JmhndWAIocmHnUqZNKQNqkICtXSZYCtECLkzz4BpS6xTJ7B1hn7lLN1cSN84Pk
IAWYBAunz+Kn94ogMoPiIirjnzhnsQfifwXzH9NjF86WH/O4spKvKVKxeLywowO+
dYfPc16s2/CfqCfis4oc/gQK+aL1fYt5QnUNdiPI/jyu0S8zrxB6vQzPcu01e4Ta
3ASgayQeuUaVnvqx/QUvt1BnTsvDCQdDtem51SDEzgCSousZGxrFGVpBt/FsaqK/
XyIZs/XZFi8Z+xGwFdb+u6CuvYBO7rYHtZ9gEU1SD7VRcn2YCCihERc1t3OHm2oE
VHFayWNKcP81TnXHTcGsKt4fbDWt6yp0a0b9wuUWRHTUqWtIfqRJcF44FrvniyNO
pBpYNLcUhGdDnSFlSjJYuUdg/rLaI/yd9ezeLn8ylYLUqfid9A5CITgs797BzxPC
iPqXnODuauDZ4CMuZyg8+R/0e1ICY9OSEba7cPr9JzYvUpWtplgfpYP7qVr/O8i0
T+l0fz/yx5PHisTRKoXYVeiUKoSNkrSv9AeUaKKEaIUOSZ2kpliUcwLp8nRrHf+F
troWEL/LMIKFlaCDKYuSLKLM6zXcPmxjExBAUf8usv2/3/j5inb4AkInOOvnFyZ8
/9JmikY5o8CYvbxgY9nCZWPyd0EOtz5mH4JD1y7DSDQ9QPxPiFJAWqDmAGmd8HVW
5jwf+xUg2c3459fhzZK3TIwLI7W/VmbnjRxjU4d203lZW4yVq4v1mtniCJ45pvDm
4wbEJ83djEVVff3R6H0Gd/v/Tvln/QKCRBzCGB30zPKm/w35lKbfH1oFjrRBqVIQ
OC2DQEth5HyAWdLP+aH3gyto8giw/6ntwVlzxK4NzvuqE+aPNVZgqjIJZ+lm/kKs
U0JKk9g7yr5ZGuHZ0Wk82Vjf9KkFUOOYJjP5ln/PJUhYiTB+0+K0wos4Oc+dbZN/
0n0a8dApOR/SVCWdvJtT9q5YiiafwTvmMax5T7Gh6dWUR3/rRocNlG4jB9bSXrBG
+WSM+DRz1anRW+Pg6eB9uFt3+cqYaOIORuGVL1Fgaph5+49XSF9HpNXHlKMrqBla
80Ybz3USGSFi/eYfQa1AV66NjOT24zgSTfmuZKlQ5blkD6GlQ27gsPNJyf3cz3Sf
0E7Vb6LhLIM4s1QZusxHJcPK1KBgeTZNZevw4Jcp6D7dn+D5S+4VMcgWu5hWEkrD
ZN+Q+P98ifkh6q38gOWS+UyIsBRHa0Ybga1kqSd+LL0+yoCKzhepg7ctNsgs9tIz
6SuyPjkWvd35LXw/kkhlhYeSeJDCMaYTZ4ZsYKR4fKrhkL0VrfagfVBFd3fy+bDh
wTjUzWevQGRoFd8VEkRTkB/LoGqpaFUAy4UgfIBOLnqAdQm6AWdi8NeeFRDYvjkY
BXwmBPjft3O3A/kFZ2zZFlUj8OcQexTgtz8ZWPWS8IvVsAkEILSjm6FeAbuMBwSz
NXDrnQWN30XLO7tV962n4a7OA+MjoW1UMZx5dEInC3qr2DkugrvUzSfE+4nIbkeE
aTHOM7yJfUD8lh4xya99nM8pALALYjX3CyWRJeswFpAbj5sYfwAa3EZINZwZziym
4TR7a1ajoEhznM8zK4C7jUPEVmRGk1rEGazBi3/DRJn/IAlggmV491R/IukqH1bw
qxJmWXxcYJ9EFCOhxTGsZ+rN5iT9zFpylWtUJmlx/VYS/38Av3PhUbjUymw5SVmK
LkRBffkuHcjgUpdue3yAPVP0aHUvy5RnH973PL1YE/FAN12dr6t+u+ojjcaPZT/+
+uh1MtOHRF8xdJF/WauLE+ePvdQjuCHZp3N4zxDVUhh7nXfQkeaNwDgMeSaVitkc
gDaSh2jNL3qn07T3X2dgl7coyjV7qG6INTbtVQNY+TYcZ2qRHBlM+qx5vNPlzysy
ZrUFUCstLnhQEtINki7cVB4b51J0cXtsvupFo9gmYJPy8oWSeHxnS8agWG7rkcaE
E+2ssSdYYRO0BFhgdb6b40j5NVXhe9GuD7PiAf1IjU0k4oSW7jYiSQxyYxkid+YQ
UaDDSiTiiRMrJC2fm4WEx3nGz12HHq7u/Sr8pj2zSQXzkJyl9pRIWGHQA2bnn9Bt
h4itAyAJTO0zk+PpdXClkh6YMF8TCUUZ5/H42t0Kqd1A/OZoNS8tG3WKv16lMDkb
j8C1yzO/eSNxZbYIYB5BDXZgQbLgPv3QmgJ06LYsUiIiMlJb4z+jdoqW2hBr9gnS
OHE9zCpgavWPe6ZWwka80tyIXHeaT6IqQbOJ+uDf0fK/9VLy1eQe0nj4cC36TchU
iIyLmMi3Pl8fwBlDfZVpUcLXLuswxo5k6x9X5aLIxaeeSQf2eZnbNw0zTR4kCkXl
7+0UbkHc/TN40JA5vL18lr6U/obzoS8dAOdcbV+qeHk0Ku1eykSuxAHjqG3GbaEh
z1stn7mwdgtKVVdgyEsry7bfyuRF4QERlcmesU3zfwT9diOXG2rFhXF1y0IgcB7O
+Hhpf1j6UrltgVMMPnz9ahYgOKmpUtZnr6+eDzUX+x5NN0d6Ks8XBB9SvcZK9zgS
tMH3jB/pyXaSXJ75hK/on+IWCRr0MU8lQgrdjGZx5JSmqad+4rUGxtAf1hCbfDXu
FII4hFGHLRPL7VjyokLNW6YedhK0uytPn2ukwfHyZ5XX0w1e4E1jNxCk5dvctxXd
n4nnqYiP2yY/QWfbknuTWTHyMo0wUWCBN3pAvODxzxPUUxmS84bJIfBhi9RbjDGm
9x1ibVzck/WGWqXAQtlBEGK0Dbj0XozNfcLID9/qC6tidwXq5G8qlD5m82jPkalq
IOexVQtNskDY0Ggjz8vhBlcLhltyhxqFVgCcwB/PO1cqI6QJJkpZzL1YZquJWXwT
ELLpFOH/DIi+p0XA/zWKSF9Q61oY754+17ZVpAV9+EGzgn2v1i0EwWOoqRgJwLzr
B7+MkvQZQMy6ESdSPnW/h6MoP89n3ePmCVWMaJ9Q68eT+I5HwpCf5ObHDTRobZq6
mYBXkvjYwZ5VI+Jk48LF1/4LuemHymkGSBK1emEjucUUQ6vKJuPhNVEOSdluWX5k
7u1SJU2es+D/55dB2vqcfcx8RegwNrkSS8CR/ddnRjgw2Ngkf2CwCMA6Yyo/P/3r
Waot2lZNGlWYetPeCAY8ds+7wx+qH/hvWBQxGqyBOe0tdPL5PGzhDXndmNqwfuek
ukxE5zplxvIpiTEV94acUXYZttOUjJPaJQTrD1N/+KpyWx9LDUFg10LZOMWZmJTF
peyKRnoczOzpFxYb2HmMXPkW20/g9avt6AK1v57agvynb+DUznWlo1XzyrNx/n+m
v75th6nu32EDg13Fm4AANch8StoWQIbj99SnzLcXtko0+8OOJVDFYTTbMtfDGS/0
SVxkZW4X1HRAXZHVxQFSTfQ2+/u+atARjRuvw9OmMp8LraoS3pkTcF//HDVLwW28
utiauSnoxLek8CIJ2/FRV0L88lUwGRsMdPeaxx6px8exzsIiIB1k+nqpX+vyVfl9
0Qg/e5Vn0ZnsirPwh1U1YLemBFmcXldSp389UAliBwkwNtAXlp60Q5CIeC5+vjoJ
VTbjfkgBaAOPpIrzAan+y9FCSx8QXJ+Exr02XxZyuWbxOXv74eIHjTgwnPlgSZZC
dGQOuAFpa4eIj0dXspFfWcUvamrs+7LBGbYA/iopuOcpMtm1YBt0gYGfv7LifBgv
eaqHG/0GK+PJYBWUp+FcNwCxqfWiaaNthSiR74UrL64uzGdZd/o85ZjZ6zDMKaIu
sQRLyLx0KJRvIQtdp9fcWh7l+G81N3sUkH+xFkekFP7Pymq5S5qtIyyldFkgkenl
JRK0AgFYTumP846do2MTGdf1He8NlfuTZdhVisLzeAohW1OJRCgC48naRCmNoPnw
R+XZ77142dbRcMj8NH1EBxZ7+pvBWptmeT6bOaL6D760o4NOuTC6BP3L1iqcwvm3
zDBloSgSaJr5uEdd7zZgn29LEST/A3FheTqdAMDn0nL4Eh48y7CFS/z+nQkOWY1n
3DH1zOVKYOkOBkbqDdtaV23Zz+BLFUe0Akxaq/SOBvJB0HUIr5RJrRGtBtxffAFT
vZGSHSqoxuXlNDiJ4iIagV+wNlGeRDGC13BIa2olItRf0WZhBTuqQbTQ7nn9ftAz
JpU/xUfYTnZqZGxyAZd+BK8f4wyK0JVXlTjbdg5/0rDKUUH2SweTR4intZ/t5ZCV
jLG4c21PlXX7OtdWi6OwkHd3HWON4TqxBmKiyx4geqVZ/Yli3SOEGgirUq5H0osj
FuUdsYqFpMYrX4o8dX4zpo7x+7dy4ND2aQF6v8K0uOvkVdfmurNHBmmH52s3yW/p
LaLCTxvN5XT2fE1puNdU/HWIRevvp2zvgZVmEbZUKj/RKQr8jLniw98GdHYCNgSm
J2S0sElHiXquxQXo5FUJ0tXpUQHmWV34/poYVqFSfozjlj+U6HJ8LkGaDo9kGlln
Se6JyFLpMuB3y/tVvld3S30jCHSRAYlTmTiUSE2GCzOcx+al5GZUV7US0LqBY/IH
sFtQrBLWiCKd7PKruYPAAbPJlx/safrirfeW1ubfzY6uDKGRjke3fJqMJpwnEyy4
zD9gsC0wbcmMyMjIayKjC5Oc+whgr5M3BuN3eRBWiOJno2YV2IXaVIsNy3hsq0S/
ayWGqNMMTrA0qFLLDnIFpNHAhRBJOttzcuQGn4ujI9vJ9RejWdcNozJvJoYUvJv2
/8H/MXajsDIIPHxqVut11lbx39UnhlHz235Ctyybsw87N9xDvM2DdoMisq6zhYRv
N4eRaNQg4pSBJmU0KSeKDr90dioCIM+S0tFh2UVKfOxTOj+PP3/P8/qnvCCVfz2m
BhnFJBa+8j3fqn5+JLJTv9+yXKOEH8aLX2p+te4wSytXTfhdGr9JQKjoDNJ7UOG8
4onq37BiLZvj/5BvngFDKin/B4d6Qe39ycLO7D1RijuPSVcIuId2P8eRruOXoLcz
vtwIa+VA9wo7i2Y1FfhRXtCoQMOfZS1GbiC7YW1sVkH1/AKmQywKNfAgt0j2jqFn
vzv1Pias9qD7rlL74cvOiisSD782ZCWgl+7+ktMKby4K0CJ2Rjvg6ND7o3+IlqMx
qFbzzBWboCblPBtdCsFk06zCHN+rRf/WQiJV8eDcLfFv5vUS99eIYsMjRAwtqjX8
YgXtA142AEhXXt3fVrMmtf24Ce1sl8Sl1kC30GQGWiozcxyJPdtKL9/iSK+zEAW3
9XKYzp5336JY0VK7nRy0e/XRyjysm2h1DfsSgQQxhQmZTYnsW/rbWGAU5bi4oXVe
1qjwQehZVuQf0B9pz67HbKySdiqP9Uv45RbekWU54liTsholggvM7pDU9p+8mcnf
m2Ozn8BhZFbtJjwvdC8ZZUBcDuBh/9fG2KxkLv37mcH/lUd+c8iQdx/r7t70KBqM
/jKsxcveC0ocSk+ZPCrdzLiIEKefA1zT0si4TDOktbLIgCXYhbuAyaRP5HN0IfXB
HnOPfnC2dQkBtiz5HhaV5+q6UPsHn4OmsOQGK2+9hTpQGkK69JePOgPOPqGUK49x
tCt/3pq5IaldtT9CIQatVu9tFvpkNwcalzgwYRas7fUgPWPxqtBD5hS1xozS+n5d
JAVSWBF0J98HTFmwF5C0mXNPP8/MqhIEdPk4rTzBhGzytOkeOpgRb8AANwGavYMW
iYQCsX8rPwcioKfM45JKcUsF2nTzCOLTVDNa5p7tlG1q2tEn5Y78uIqvGzY0ZqOh
aLus74aLhD565hTc+E7Jl9Q7CFAvo7B6Ns2zHSQu0+C0mhidt++wkoXIEWp28H/t
ttrJIvBySV+ZoF/5pIC9ifwS38BgaaaPPuj1TKykytZioT6G/sFJtA4rENtvPxFz
sbuezzKmzs2FoZX660hhmxLPYvUbt3+fDiTglHXjFzTcVCRZ2YY8KFbMa5Vo7GIC
x3WYWzcFKs9Qi6Mu2z6xyfbHUp8dSonF+OPEr0owdMGmgkTSCDz3Uhvlz0w+ktPl
aIti4JVqMtooE+HFVLzxp/dnlW0oiQP8OoAaTqpmrnLRlTJoIMrgHVpTkdyfI19W
+c8OLJEsjLAd0L/u2qDmX+HECXLM/yoOx+dlqzP+TcSqBaNV1ybJ/vDGTjBvd4YH
D3Tm1wwL1YRr1KHUwbMg3f/ElunjurZK68LR5CypJ5SAtAQarZdJTYwx0vnE0EFp
OBjxC98lHe3uJ4WcMBjEuaktcjEpHLYWfAqxGHJG69xsFscTBzJZHbmCAeYYk9wp
J5VZHBT6jnUlGgPDbgJvRW/T/Y88q9j4Dx1HkhArIdOSYPw25YqEw6/FTj6cQOeq
xmhuc2hHrOLEU/Tq17ni5ULfm3t0sa6oumpWiYqSzvqszagsNqlLB46vbK+TdL8m
QoVoN4XlqcV2lxaPkx43E3/m4R3wTP7wenYkJ4F2C/O8l/pCcDDzqpk7L3D5m3OS
lJ19ZNerqoNR36VooWCWL/sxllNDp81Tt1HGtpMzYZ5r03fJtV3FYr8SfqiB3oD3
77a6kMP2I8V7cKoJN54gFDR72l1+UqIOb1k3OCTEIdxsQMLCEgvfN421Gh1xTahk
8l719yU30IhKR3JFm2Iix4GCMknJd3Afnv4CK0ubCXLmfTlPUWmDfelixPDcJg+/
aRv5bjfkMhxaVuX6pYwZD3FlG346nke+KihuiGhNmIc/y4qEh5PqDMMbsez8iyGI
Oit1wOMoCVzJfA7hqeHm3BYlaQg5pPUppsIz4EYiAs9vj9ZHPNqsdAiS/MUxOict
BA1Z6oXxaAfHjM9RFJJf3hDGioubtUkDk31FSSwSlt0aA7hU1yecawLnsJN/Eqdi
4fBZ/qC6O1uDa8ZfakbkJfP6j1QBR4gjvFcrMOQ52DS0hIca19CRYQTWWOOSgs5w
mVp/xr6fJQ0Fv5d0/lFldS/tU8zWECp1+ebG+RZoYs6wkn5TZ5gPxL6V9tAzELo1
MqfsSaCYkWh9Qi0V3HBYKh39BOSqQ5gpE6b4DbjF3rDrzgMn8Ol0MnR9ZyrQ0tyo
aOYQ/kUytsU6vWurH0CRzA5E2GwHN++vlBx87xv3KrzwJWFSBkCVHwtrWIWjYwGK
Euw4ME0J8j08gwferrakjgu2pC8GZ+LC0mWfHyM7e9j1bwjYIjdmYifFZuwBkG7l
Wz4QNCzB8+QvGeKKKfTkjVCehNotSfeMcW7iu1nDppv5JcO/pVXV9o5mwppAfzu6
dXbdZI+oLqxOWMXpzqOSk5K/zSYOZsrtoMahfHca6mtKT+G48eYpF8ugigOAtGen
cB4/YYX95HmFUkpCNV/gQf+sj3Hf4tI0WujvSWJRUdAMGDEBPApRDBYus7iR6tX+
sgJsSU1hhfSNNaLoSVEiZioUnMuDXohtZBCrT2KKL0m5weIplMRy0yQOoV7EsLeZ
STvJXb+GGjDkotkUsOMMxP0v0hW64SQyFyR7/w+QT+0bd9RPsO6c5SHryGAsz5w/
IR1n/nqqp7j5XeDYcwd7jGcBEylxIyT1v2ujhKbFyws9/jwWOdcni2BxIuFrWFNy
ZQ3z+vFn7RtEbO9ZkR8PukQEfdZl+DYQEQOnXgTgm8gTBZ6K9f6BHolzoDvXeP+c
ZLt9p+98Sjou0AMe73Rlawo9soGEsEgVw65n2MF4q7sh6+Z1unBIcX+4zC8Y1cPO
QFIJjl/79Z9XkHFY+1J+w60Tt+AEGAoczHpcVbBr/WXCjoeWnHxasA2Zy5u+EyNh
ySBHJWjndySV6bVTS/a5q09cTlohc7fJ+KBRNG+kk+/RHcioI0hdFLF3bF78EhAq
IanzCFgE1rb0fPZkWjqGqE/NfmvpVV8kM20nJmgMSrzVZr7uMgv/92/d3IMK7SZN
E1BbRKrX1v9e5Q6lZ0HNemlzbl18H48a05hBGK+J81Wj3j8C1168N7laoS1H3hw1
zc5siZOBiMm3M8mInbNu6FWA2bGNrzN6+kNn+snxyFMtqAEBBHijbf63+GfxsHWY
f+QBhr27rhIFkCRJjEPm9Hkn9Awb/LoRIWnl/iInkRN/xcC3O0zAawY5SE56kus4
Sm9iEyjADrU7C0Ce0zTQ4aH236OOhKAozMD66yZxPu4qUA1CvIUvmuM5GhVEOd7t
ZTWC2vZ3kzhKGufq8p/TmkbP1T0VPNvtLa7+WqPaKp/qP1yUY5EortFpkz0px8ke
RZvpGvUp93CT6oQTSFvS3FfU5CCnwpTPFLbOrcpYFZRjatZdRJFWXLRSkebkPr+l
JA0Z6KkZx71zPyaYYW7+XyqLfZFIywTL1BjHHBE2wuX6vkxuqgl8hL2lWDI9t6wz
cNvyMpN2pXdqAju4XKJF/2bB3Lrw4rwKsPlR439U37cQexHB7WvJWq/FfaYk/opG
ugYB4A7VvbbxQrk7ThEnf31HSg6tmCQBxFhYoP3OGLbIQvuznRHzQIOpaKCFCx7H
3SMuJJukKzBZR24rdbSNL+ZDLXVrLBLw0dnZqdKwcxsSPrSrf3CVv2HATAs2keYb
xFNVQS9IINlFj4q4o8aCVnDzlNQSKafqFCAlOWgnReZVIxHzhIIK7iQM1a1jrDxw
ieuftp/4qdkKwfSwnOKFV8bI8iUp+BfGFuGVCPI5LR8+Bmkj8KiQ0u9Ko3zkDo2/
M3+aGCKwrtUKY0zlQlZr3pjyMVZvv9Gc+p1PrsTWxzbZvd6bt4lwkH2cK6aO5ZOf
QZJGwnH+KWDb5oUQhzGfJflbgYlUsZxrph+HGSeNALHAFPu7hL7gNAC3fMHiY4zr
pSGw38a4MZNZAc9VzG9G1Qdnd8EB6+nu3r4yX989XKrZQoJQE82StRPU0GTE1PAK
3kxt58/zwHQJMGL/x2CCjyGZprGapkEfDFlTTtw5vegHXlX6pDmgFz8JboXBoUJE
rrZkwdPi/kL7TU+Tw8FLnmLMed2WeYJwMZZmd7J3V9xoZqJNlu0zKvvMt6C89571
3AiMCeWWFQq+RBiI5MBoSJjUN1qu470TzFYlHtdmhD+ctSnmUfjYlSWxuzn2D1Uv
JBytPfFxqhUtHKxCyKZ2TSyVsRIPlzNQboILmtTUkc2KIFkKz0M0GF6E2ELfoWBo
PYXfY3zKON4f7Uwlu2j5DCfOOuzlbFL8kR0KO1K45SY26h+JISLcaJRhIVKT3VCD
ZnV72hwboGp+EoJhwqNaWcHaTqCUz9a1z6H9DamCefKTFjeV/UIzJ7kReFqC3fi5
S8kl38RQjuAHDPPYRfJba4lyoVwn7OLyDrHk6nPaIPHc7jHDH71IIqPUw6eI0KHF
FQFpgvd6V9bjSqvLY84/VxGX7ICTSK+irWdRdhmdHhfgXen1zahXxns0axgL+gxf
+cGm+Dni/GSzUQfDVnzMZjZK3rVM7PyshV5NIAE/5dIM4I7oWlOrX1fYombEqmYQ
KQmf7YFucu5gyep99H8BPXQXwn+YJg7pEjbV4TnK0iFwQultQTtFkdmDqJWGAeRJ
wA7C2enlLYQPalPbe7cRn7Qj0QvtkQ7lOMoF4hZt5nMs0Rb6htdi1VKoD/nOyKaF
CDbB2f1YgaZzIXLKaIOEqZkU6tJulpO+QlD81TA0E01HXV27g0681M0c4hvYZgRc
gWTLUW75Uufxvx4JiP1+GkNCtdG3O/6JHmpBNMcov9MGXwR+fKg2QgG6bnlnpiOO
djzo7K+MVbfS0k1AZByOX+zfr+uFPvHn8VOQYc4tuli73nw6Tul7VuPeqS4axkiU
D1bf3ujCPZuPrJ24HBL2VMlJkRV3sy6pXsUOYoYDY883pUBqRGUJwZkcjYHx4pNG
h7k2M3AQl7i0OJe7sqw3Kj6AYXM7bgFLJqHIR9RfHFk4hUT/CzSr8gTYaBH9gD1l
Umh8/1HOeDEz3nNlyFHhHxVRGj5pcQNlIQ0wOlPdTBMvWgJVVJz/btFz/VrOPeWU
KOTM/DoDcorKRQ7QaMC/lPoxixjKA9UzeXIMOF3Wj7boUT84mXmvGiBp1gSL2oeZ
dOUnW6ESS3yZ46UBloF8Wj1xunawV8tnMWB5B8Cu/U5pHlogA7zTNcg0U/tT31Z8
RJXFP2sbjym8muckCMIlWl6frE/JslG9+fOc0ucFnK/jAPuhzvqx8BRVX2nYNptN
HHNI45EyKqoyMnHKHh5E1efue91c9g8/5nUf+Ty7mowEvMixIR7OfFwmLOIXnZB5
LFeRvHESKqN81CClFuYOdFoOr9pF4kXy2LW7AdKZ0TcMJLm+zpttqtCPsu9mV5rD
/7sT6oiqknrippWrbQdnSnGnqfSxh0FjdLlnVxTFbQs44Hh3GcsIT3dZ7wUVUfEG
pOIOSLb2aqGd/v0IGwokkmkPxjqlo9mFMokEXqW41h2dCI8c7mtucGK2vUI/9QJZ
YDMG3CQrdCJvLZU+QPnb+OuP0nM2DM0bZDkHWYd9wwBqI7EjfsZxtYKEDTOzsbhI
8WWxqf71HGz6BnLQtw10LgBNpcNDm8nA5gY9zbaz4ilmqFhxeRqg7ZyME5iyieaO
Z6Yf1H8j5adrFLE4jev1k83B0rfyAJ5zB6iLRzshRF8ybaydabBLZhA2byJFJKU9
jZYNjuyLe+dYG72obVaZQUlAHQFNiCHGOu4E8sPpsxplGaSvx9LtRf2vXmWtTBak
1RJZ1hb6nDUP9xKr5JSK4YvqSxqaGGH6NGu2JU55Ww14NO3R6nkZ7hZKMb1rS7Rs
B1DsLkL3zXchZYvpui7oG+ha6B61fg/T7locABzcEaWAjcgWvWe/99gAGolwFmsd
I/AWFBZp8el8t7RXRIhxGmHlvb6ZxI59hENjLG1pVRxQ70m0jz74itMAjSRwCleq
e0P+gkt57pk4W2HKoup6lUctLavVkq635S67EY6u58b71feoJF34pIMieMn1mhxN
HY/u8lUFNpiDawJxFPzW02Gmk2bUpuGH/RnIbR+qqapi5YjbrSZ1hyGokcHScpb0
+HeU7dFcKAJepWhJwEzuDUx0HTC8pzABMP0uEFP+MdC4jTH6/0hTNSLGuzH9UOqn
354SZurpYxw4qWRFBIk1jMIiDxOjNZwusF2A26+Xob/8nIUxWuw7SSrWM02AwLF0
xZSHVV85iqm1TP2Rp9g1ArltcAm1BaH/rwfuih2iTXbQPKAoqEcK12RycF4pvEK1
Q7Dx1cF3pgPeMOWcWFZwZeSjAkhMQKdZ+LVZhiC64Z9wVi1gci7pOPXOji3Aob1/
isB0wcxhKAAyeANfKNOcka65rbGeSeDinFUR5ZfaRXY4UZSQwEFeYKMhkty0U4IQ
I81ftlt0FRJa8b84VkZNUsCzq+PkQHv7iMR2n9KL3nOzqkZwQONNv9qdlfFb1Mm6
vj96weT8RNHzpkHPiDQ8IhUAx+QTYNaVX5uQZtRVFfNMmH2vAfQ+nsLQ+cYi4BqF
mUihw6KdjYR2pEuO39Vu6FWSacOlxkR38WFoOaZqoQSwHB4utrJmNm8dZTw667yB
UXemodrqDfDNHyjcestEhey4D1Rcp/GnmjB6fHApod2jhXYKztq3wrcLfctRapg3
JS7jWHlEWs07HMwoVltPNoJ2vEqew87N9PihK6xYj8JkuU5+ajYrKXS4nDJpJlQu
fF9w0mzohFvw/vpZwkahoeaW4EJ9+42PwRuOcRnBBHuYhJZ9+C5v+Q+Mwum6QWha
GxrlMk5tPHyxYo21MgG1+Am39EHIx670QfKzVY90LAx7c62GEx9ZtHKMb9uVSo/D
Qt/X31XtELpCWDw9b+dyLH3xlFDVSb+fxfk5qaahNMqDmiv5Ik0tU2mMjFEikqBS
7P67IAToyjheanLeNaWLr6rtbgnoyZo2t3PL6HPu8nZKwg+I4aNNW6s1nEdmKas4
94HbsVjPRCtt//PovNeLQbbF/rCGaI2bkebbM0jcgQ3h9BtEjLZtM557l1wLPAmn
81zjcTjg7DFx+Mn1pcDGK5Aa3wU0alAC8wgyLhVhOAFcnzntFGESMoDMzK3Dkf19
IgcNPBweHAapy7dHpdamxW1mO4Uddr5TQqI3W+RgxZsdjsQsvOy37PxXQGzhBw2g
mAtNvhtB4x5JnmFXWmZbTJI3BX+7x85ljEgX1OOcqdEreub1uoVgbKVmm1McnRFu
SdAnreFwEDzE61WBc09untGIK7Ll6bCXjSKy1XHpUJWB65eQZb4PgegBecIpKLI1
ANTZ4KC04eDxo3zKWP6nsGWUYtjpBe9Af76iZgz2qxP9IMXdj/y/kxG1ieKc3EWn
JQjDk7kX1E+Ygwo9mSYvaYTJFXHOPz/1S/O6YxIcXVPofKtX7JOpZbrGnh5CZFlr
qPOSBtlb8UP/5jat91g1boJe0t3k82D0XvXn2rmOM4tCnKL+LDMVgNojtziK94bt
ZcUP63KcCHa5/0/oaWb0mlYn0AD9UpFx5pMZzo9qp+BPEeB2Mc659pRHL0AWQ8lf
j6fzcqHF7EC1OReVmMZ5B5dJyWqARKrlCn8xgdyOib8sZckzJObI8WdRn+TY1MYi
hY62hiWRXi93UMDiK9TJvVTLnwD2YVahfHBQPiByMRhbnlFEa92XWht3jve1htIJ
85hXGImjhhod/L/BEXcXllm8cjEJfCdSjECecYodQR6r7JCw+67Ggr9ajAMgeSAG
reJozSw2VLlgyK7V8sqTtW5XHNSKlk/We8Vdtn1GM1QsE7pgFe+4K4b2tv+sH9R5
925rheBShu07/jcLVXrYcMZtIhk55+Hl4mllC8LLHWHU0PsISrk4J5QAnNx5Y2Xl
Y2lmEByxXxRLNJFXDY/KdkhtlHTqEk7zn8eZY6im8sszDIfpLN/OFLIBj+Wy43o9
i8e2Tp3+Z0OentxNrEyFirRxi2Z2lTmX+eg/PJW/rpi6y3eU2S6FvzoU77xsPoG7
vt+xDjzVykbQGj0Jqm2sXEt73vcCKnMo3tkivKfQAVQUd/6UNftgd3GeUT2inlX9
U7r/0xTeRmnyI2m61c93Z7jhmLjDS2cUqpyOsl9zQ1g/MVWKp8OJiHy4regPocCR
tm11giDwTy5LwykmCG3DwW6yTlAVRm0S1ArSLluWYwpvzFNms0r5RI0XUDjvutzA
BVK5JuwJrouzRDj8Qi/oJPFLhs0tYH8mwEOfuAxy62y13D2HuAxBYGczJlwwh72M
P0axG6MRbkdT5KrvMCokYvbf3TzCmzU70plRa7sNVTUqmHapre1Q2fBnQp496C81
Iv2sWnih4+fsddusc3X4W9mVcRS+txOT+bZgQ92hIBL+fSXB+TMEmE98P+RfPt0G
M7uy94S+oABbS9GkAfS8ldvizrPZROM7Mo4v+2di0PVweTD7nE3MXqKx+1oFMZO6
GIwyESLFHUEEStSl+D6LiwpUBOJh6YP93+s/tZONbGCTXFDV4w284xVnsr0YKXvI
GWXcqKCAnUWGNTJNH7hF/y3eNE23o98rySgHhYxa40AtH2oaL7DAyFOIrQ1YnwUY
52D6Jkkg3Ebi2H6GlenM4P91Xydtu/uxJ8XpUmxMkCpFE4Bsj9VM5kaj1KSG0IKy
6hf4CwmK9Geyoc5KsDul0SJfO1IfKATsDXTbVwQT8YksY+Hlrn8uNNV9YfumVEvm
ivRM2Wa5hG/cXShyOitBpXspSY3iCjvjHBHu7rwYu8CF2L/DsyhIcja4Wgjqb/ip
7OqZOgG/ys8IoIanPpaEb5OTBTOH+PUADBIKYkKbMA0S8/qhd7cXZIjk9KXfWgJy
wmaFdMakN/U6mzuKKOwQNlHwBbunyV6pGldPoPyF1f5BSsYrr1G2l5LjxyND1E0d
Rz75DdGgwkIbUxjDz4vbalTc3U+UOfn0INt/sBiVE0en29cRFPLiaRd/yPw6bKtQ
33bz2fCKjz9ltOhbUHuErfpHGm1A/LS9MyhZare7WN0ZhRgx9sU8ozMedEhBQYvB
sMk3fEdWbgvyI1v2kMmhD3ILd7SvCYVVIrPeONJafiSJD1q2LTN7KxlO5F5EfyYe
PJRuXS2bbEmtwBWFg6hzKXAvzSlxLl4mWsoyQZcQd0VLufjSfGJJNiOw6FhCTqEL
S0DRBEknqCKhrDlqATiFGMzVpMTb98EqjnV5UBB91zKDbEl2gOD12EM+/xQOmFLS
FDVRF1q88yqbQCW6VIYKez6sGnShhA3szIPra6ODmQ2dfuBZaQJyvjtiD36l6iMq
NU4RflHWW3Wl3FvyYCAqIuj/yX4PvaLlKMUrkUce/jEsTfktm7u+SzUzdbxiwrUM
C7Q2YMHDIZhbmh+kOpA9uQ6Q+n5EIyhWr6l56xptyqAaTg9I0filoMaa3H9meqEe
65+J8Z+Z4NnHV3KDEkY9+v39PT+J5yqZk1nvbV6SLfwbRW2dB1LAamM4SQiCMcdw
6JELbHNuytxqLbyzcbCBQ5p0V6NfWidYYoOPfpDGhiilGdFxcMzmjcgCm7gEk+hc
q5AbYS2NCMCW5xl0I8mH2R2uHtDeRtsgaIL670KP/jBDb3XXFlcOITyiZFTXd426
erSLFOT2qkM7t5BegHATNJEeGLZpGYr4r7VjTSIdMPkWmJ+clwEYrTkL21gBRN+t
FVJ/Y4zRvt7J3UsbHsBJfCO3/QyWLXCQUtc6qA49DZE7KNspML7s9/M0A6ksoh+u
fSv00IOg68Sod+bbhYe9IEoeHo1X2SCURJOcojUDZDcKiEUTmzz478k+jc9LYl/2
FYXSm0OgKlmCvO7jGF3UuPjidJvS0DMpU4x+jLcHyk2PaJlNKwsLGHRqpnfvREqL
W12cJTWgxOFd3aspROc5vz/c8iuH4viY0yjRzjJJKCN4HddSunTGfeAzZ23eH9+R
pBYUj6WbkMCu81LtnU2hvADwcoWrhsaINESJ/c1NJHAyW9nupSG7WJkbg/QVJkef
pdGFkSDmjbj1jgy6XgNLG3JRYENoI8pKD5xJVo9OruHJLJkZBZH89I7qu4zGA31q
34qoz6gFtcS07zbSlElfg9Y12HQXe8cs3nBlOTDs22WCFaxOR8sp631+KhTV+fCT
qDmh3DiGQ5AE6dvbvGNSaUemGr/cIYggL4CPPwq3lCilemXL2jtiJkYbFHQtuT67
0Af61Eg759QKFYTPORKGqU08niPZciK0uh7L2P/0Jxic5tE8gzTqEF++VyVxgK1g
1UlscjDFg27oO7dfdFDO3qCq3Oy6KEihWqb66X1gUxnYM9NUHgSrmotXP8gfF/8v
XVExWmMWxSe/v0Li93SUM5N74CM3lQG8eKK8niQd32fHVL+hgJRwztixDH05yrQb
h4rT30J/Mmy1zt91e+Fb7tDk1YA/5GYYY+mQwtFgQk9XlgFQbmgpIeglv2S/9Pes
Oe/2QCwGtljkU/Z3G4arGAw1Sh8VCB8Vu4Sbd0MTfnwWfg71G1bKtg58EFA7T9kf
qNqn3rOYOmwSehSnYSDJhMkoCsiENxWSbLL4wceTFbHByP0h/d5ZSwCaucd0vn2E
ty3HkaSdYoO0uhbs8oesG+GMQIDFecVUb6S49bUmkEU5nQ90bvByCRYoPvN18XEN
opb1cXT/vwrUq0hgQOWb9/wHY9zJm14aHVbnChU7gtZT/NNwn6FqYotbuWfmaki6
hrR6LFlxdb2JqBwjnUL4gDCcbmo6SWmMEnL8bLEFYaDilg8DQg2eLNgWQ/4vksRa
+o7i2TOdsxRgJBDyMNbL5onbPrmnlK4obvicyKqTWXyqgMtD4kLvGtXKwigEiSz4
72/Alg69Pwbo0MvSRyDhEuBuQab8vTo2Nhe69P2fcSBpgY/5NpoMekvimG1dy8QG
VPJ8Y4/EZvRED7KuSeZLy2HJDenKzacflmj0840LUewGtN1/kyEWpG6DSnonLBxU
y8F6L+sQ3dIPaYNxI07TiKtrmeiLXuNcP0iim+uVwz2KfjyrscefVlHgKe6NmaTe
U4eQF0vnY2Z/XyfDwPvirjW0d1vjaBOR/dpwyJ5quqOZaPjoG4jJ7/kpv1FQLgTH
QWOOH7Pgp0lPn45+qK5VcQ09amyG498shfWlT90aArQI7bBCI0a6y0M0Vqs23MWw
3Q+S9yIklIY/7qjDzf+CSxtHaGZHgvxrrYCQDvMm/1eIb87Ol/jbkdHU8js93/Am
6owLd8rJGSpHqwO//ZrsGAqggUExKDstOmPnkHEJO3l+5xr0WpNKc+pZ1DfGN6Sz
v5q0R6VJTpUAw1BKlivNKm4XEp8eVuvIvcYiawrPlPgchQc5eBiQP4zfQQ1nVOH/
cLwn1L56Fpk8yeoUKQOI0mJFS9nZanxIGfAbkkdZ+4HvnHM1ztZ4NHPAhuGLyRfG
9JbLtkDa7sYKRHONu75uWT0AztfBOw1M1HAc1xQqGDMLrIo1BpfKJwiryyuR+qLh
d+Qt7AnCNsOLDlc5Uuj6qe1cwaxN3FJtL4vH/4dCFF0FEuxalTLljlZKxLt3XjOJ
Xf1/HErii+0JCafp/YWAdydza6y3PBAXI8R9gBMh5SS65KfIvP4ogndtH6QZl4oK
zdb+hMBKdk01OVW3qjWJmFlc1MQ7pdauzaVoG1uQhdcKcPY7AagGvc6oFJw2LOJ/
ZObwhv7F4vVmgBO9bOMtjr1YJh07D0bxKzWzOCaE6JEbNmx2Rv5FQzuXGlWf3S0t
bKNOPEiPCM1QqFMkcpT1n6OQhAPfWD6WbLzyMLL7zYCTEuRrZFRpvdItWKY1ARCr
HBcjTTvGxYs4Wh2Vs/nt6CSUgWOvBWEC058X6HCqUevmQ26+x9rBooOOJfUeC/9J
OZLim1InktpXcUmiNP1fYhd3/PBL98j+luAGSWqS3DLUYnHMJEvCwIB+Xs/F4cZk
KWZQojRBqF4U/ePtiqoCXx8u/LersWNVA116OYq52KWRwpDkoo00Ero18GHgf0+r
Wpp7xQu8+Atu6hd0068zAw/8xzrG+XnNtDOpT+7Qj0WUqKvPrQg/B836Yg4o337s
p63aWu0lRoomEc5I5EwbwLJqAuHBIktOH7EprL8JupRCfr5YhwTCdGKBWiUuZVbY
ILZmtzk5mkYkEWaLEukcx4Z54kut1Yx6+IqrO92UoT0+wuNRFWiHOd48YtBPsUYV
MWiPDqHbYEVARJkTf7TKMrqXqaiY7ce7NG2rX9v1Gxlo3umBOOlQNXW68MUFVxbX
ez5b5chVN/JZMYW5dHRKt67Q2i1zQM5dPLtPMmxMrlJODzYUfw/j8LzvNORiLeVs
tZZVBhg+v1VR5ec+fpKCfu60ajbctF2y4PKVH3PhIZyaeeJ3eUa9nR0C6zkyXHpU
PQwk3Et11ogHK7gUn1vyQ8bQKsBmaGp8mE3PGMxppqjORj6o9b7U7ZK5sHbjFiAr
Av9xAn5BvFHt/nGywFO+nskPlGS8tAbBdUiWLmafKpeg5RwyopQlziQDnRDtWGKb
Naw8GV9RZTFHkY5qoN0PODL0dU7YKqOgAaGUR8OmQVkj4Ld8OGfDWqPc9hoaNjNO
rv7VfJPu60ZAc1+lWhaKCdbz1XzT7h1bwh5EslisMlRlpVhlnsXMr6fqMNcGHPkF
wnoMbm3xbI9NSbGuXPC49QVubSTp7zsjtmhtHeJusmztO1mzFIhWPkegsc5CanmX
/VXl059D27CKBW+V0QfzsOoYLz3Rp/DWPknBru+C7X22+3VnIgnyq220X32inWLp
SZ1b/K3M/opoQZo9dO6Hg/gAuHl78W4OkkU5sujHLJEyv6UP2EasXSmWLMLxcq31
2puawBdPqBzICV4S5jUVhmzh/oy148TKuccbjgtNG8RwyyK2Dmplqjj4YBa7qZrR
V02I2+ICEh511czX36auN3aY3/Azt0x/rwbLBI1tCSsV1WBViqwUV9PifddNzeq9
NLlbdrc81Zsv1Cq5T1Rr6yjM8lzH0X0V4qP5ub24SB3GLb6uMc+Vj7oh4YKRBF+j
puqQUvwVYdNUgqRg2FG/S1aDCCLQUtwrQbkKhGv2O5Aga2J5k0TAUzKmqEa3QBDf
YlHIDi3QsAezWrQQOcvlZwxJBoR7bJf27QeQJorq61GUA2JwJf67EpOZPsZac9ph
t74rheG+sRJfH6uUz+JFW7hn77LoQrfEvrjR+xbG9ISIrInTri0fpvBoFbaOio3L
em5Watf+hkxcpbQPCFU9DydikpiDd8Nht6wd4y2sxW+FtSWYIW16c/x7MDoQbIll
z39i3eRAQC5rLDS81dsceQerw6RU2Pnc8U5jnKwzjOYIunCA5YrHL+R9/XyjEOEK
6+8pDMweL4vVNegapvoUqIu01RaKXfmMz0Q1TlNdD7BGiOvTZ5HWWhDDfIUrvE2+
+e3w0JhPQPvJ0eGEBmH0ZApD2dghHxrOBuPp19hjh0fsizph3RjFVjt3LUd+dgG1
IrR2QpM5t13vkgtnqUGhpsfIg4UMxz/OHT/6uGa1vNbEBnMEih8l9OlBa51JtrKV
sIuY+byVbDNHIKuDesoLA/dcUprKLkwB93h76Si4ERXC3WKVMqYSTruiMSoX+oQJ
RIeUW6qLalcHuUX/toNCHnxoW7kXzR+M/atYfaDH6l2X+ccXnhXIZHIpcFH15ceH
7XBBXMggBgw+XYqqTDgrqnTOxJEAupAA7R3ingqYjOhPBO7q4UuYhJ6iS/3ZZHns
vB98pteOCdzN3GULu9JeAMAHMdazBHUh3ryazgMmCPDy7Xmu3cv64ALYN+AGD+kz
FqsQ9bPop2+U6tb6xHIqq0c3UXI5CqHfJFqvyjIa3wbFUWeA33sWrmR1uu6UQ8P5
0zoYFPrFfSh7PlxAIUB9nxXQ6fCiu5XMDGhk7SxyH4ExeiqXOsy2k9XSb0NNJIuY
7Or3BSrIPHm37l6vIyOcOA5Cpd1OdDa2cRaXoRHIOZQXWphbVJHupUMm6HgCZZR2
/8bJY2YduIkYBpOvxzRow7gyrjiGG6AX9u5EvKzKc+tXwPzPwyzoSkd7etuOwObU
tkiw8T1e6pJUX2f/Tat/49W8vHvpOHqRu1xxZXSLPgSVgHFQx0+Fo3FtP5McrF8c
KPlZFlbFo4QWmZLEI3kbV4ndJPjAJTPqwAk9Z/qpx9g8u6JgQF5eM+33a3CPjOvb
6UhUbPFwlreRWfskwnJg12cyqGwJcJRFRd0tPnSkweDnFOZCcaWJoQ10BQ315SZ6
Vae1DZGUlFOAVgyRQu04RIhXiZtsr7VspcQSHR3A6j0rUFH5tZ+gNHUM+qDdaCBf
fQSJMZGNLrDd1jgbE1iY0764XDRnRfS+vTEi9YarkqSt9GmnfqH/+pTZg0mzaRZN
/MeshGPosEslVH8lfYPRfsPuoFDVSz4RR/x4/PXug2wfMzP2SPpBds/8rvMjzc2a
pTF4I0fZyk0+YxO/Pq20LmycbkD/rKMlibZsA9lkNEV8VveU4GKuFWxLQyaTdJTT
pLf7MzpTbUVZksMLIqrnHb/Pj9dxUAFCKr9FacyQf1RnRLdkSs/lHvE2Zv5e6pL5
wgZTXS8q9sFEvzq7o1DMrxfXOPyYe3K3URKnUErPtffwqKioS+pnfBoX/uF6dpRX
SeswaA4R2iTuXas2OqTWv2WpnzEraB0E9gm9LZW2yZ1NNe0W+Ih7LTeIpNK+BDvz
0UthEj+ejUhG6OE3FIvjAgAu/D1H1g1hB9B1xP0vsoMURAlQWo0MTyZLD8ZncwXk
m+0VB0qFHKEhs6aNHH/Y1bF1j8rYJFEoUud3D7yv3lIjoLBF9zS+1Bb9xnJGrkvi
Hf1GcRkSUfdQsB/dnyWublGKJjSyMczHjS6DGTczMOalV5drtPpIab9xpZbce5FM
QNnasqAZOkdQ0MI3KyyRgvdc6/i+8P88EfU19KJsP2nWfqGR7gocQioEv+K0TDzB
3dDT0+ppwdllczJxFaF4UqJkjfTSrr6GyM8EXpIIvN4G16k85ZfTMYFWfmR+S1LA
u3gXhG1gzRuJcinkYG4kcvGjciVXHdGiN2c5HAYXhkGtfuRjrDzesknC5kGuxreJ
5BFN51q6Kw3NDTqYWQDEo7raL+jjBqGA5fQpJGwB5KzGNkvz9SEob7CL90jF1Te7
qR53FVu4NbObLtfVpJqK5IUJypnTV+qLSPJe5a/RTxmQ6hUpVA4WKLJOJlLofywH
Ji1xBawEllQtaomHdVD+HcUyYvJVC3x2syN39WCHsFXOqrnvuAQMx+MKJqgt6Pc2
KSlqTzLnoMyMzXomATIbjPPYcIa3VDSMBSwuZkHNAKDCYm2YgVgKHsQTTNmxomij
a2RDrwgf9BWpkqrPt3wSg5WzHSdutylBYjbHYpWwDiH7DMTW8hq7feAtv5vUIjZZ
exIp3lv+y8dGqdRXbgjPHHs6krwsttNBlclPM8CdMbtEuVKjW4XwPMRQJJ5uz+bg
FVXYVgNqxl8nDA0BszPXzoLVGGB9rEnNCZfGKuO09psuZpFDWxNDaTGtjzX89JkX
YLkNZweOPhnvXvjbY3ka1c/sTb3F/sa6LXr8tKi63MTsg2cvtG/XCR5gGB1+kCma
J2uZOm79wE+WjvjF/qoVqeDMplqCNzWTYPqtxcLpFt6nmpwwpt/nqqC+ijFuALzA
j02UOMEj/GHN9Lw8ddIDHq3PSbsoyRPW1xrZD8lh/ntBMmOwMaXpuicfuX02mfq+
3lkTMCMdWHhKIMEI6FiXPuA5mEjKgGg/wAMbkWEssko1o2/lpn/JDhlT7XmUYtXm
dPne8GaEVTRphNfFHWBp3I1IjxwJ1C06Kd3wLJi/bSU7vj69z4o2tjI7IXNV3fXe
LDzeYnPH5leNdH4kEXCOiWplJXsbP02iyadpaW5YvyRAnTrxxakYaq4HD4JNQV05
aywjEp+I5etotigN46Vb77Vvf8bwGUME3xiy2lC8DytWPmVQ1Ep+x9UFlR1zKNSH
B9i1GgcBPoChsQJQQPev5wMyeYjkcOJJ6Wnlc9P6B4ulPRyZgyBKaIgW/5WH+45d
mvEP6+5Fc1EtAJuiLbQR097673y/7nN01B36TUDD2sov65OHDcD//kJ86rDJQXUi
TFvdrF0ikQm1uesoF49ZNal+t1Bl5EmDZ6M8Ho7eIgydVbsOdsIMOdXkd4C824N6
gEhQSgre4WldQUv2XcXxgwPfn+uIYxY2013tzZLSJAkf1fTY5DhmIjpY8Q18SOIZ
yktVopfQnbBRwQdZbw+E4hSsq+28lZNYyOQhVoOVf5ecZvp6XylaSZbPKm3wLt6F
jW+IO0Fbf7rtHf0qS5HtK4hBo4rNHvimbDrUF3oTGdDgCVLWRhIwIpiaCDBR1p4A
tgfpzZvRguYhH2dj/3W2tCNO16daaPAFU5T3ZSa9pi7Zp6/XaU++tSg/1Aa+9gq1
s8Y0yrVtl1ILzRbZ4b4NBsenXmrYOUryqEQp0YtAqgFYrmWPfdW3QhstKv8ZRHxm
yOZ7ytF+caJQwcv5MXfye0ApsvLJuF9mEtxSdjJhVuWdF5BOKZ/sgA5Vdm2228D1
jtq8b2mHCXqzhVEFWgJFyXS4SC+ugHcCSYIsdGT75Nav7Xmrl7s84dogfs+Sg04F
szaiMeLl+/r/dXOzu8P7aCLwO8EnyFjq3H4UHl/o3VaqNX2G2Apha968Jzyms9bb
hpCEs5tTzCBmYoNfbwh05XPQtFu2/vL1PygT2NTxj95wuYea1fgWCKQAI59AFd68
qkBAfuRswYntNNew3tTtTNmPxrPCbapQKPvMtcYLSSzbsMSeUpgQq1bKxr3Hvjj2
8BAqNoggAtq6h+bo18+36efx6pzWAMyA0g6k65YEnXef0XmjVZzvroYdoyZRbeGo
ljQtllq1rvpbYGFFLDzioQKHdn9ybvWlBMaI8e8cGyq7Ijj9kQX/7hlILfeVQ9l6
DTh8Od+8x4IGFmntNhOE7uvFN/Rim9hXIATHc70b4mgLWsm9diYWdHraHecNjYPg
zsoJajkFqIg3B7XLBI0fyjVY4OujrDIGOanOf+/9UeBYtJDMDOnbkjocQAmKV1ly
ElPuoKMqgS+fVdvORugYt8K4yDak2YbV6eZp0UQsV26BabZODHwA6D9rkrazqV1w
WBpi5xmOsH0B5emEFdoI+mZr8Fp36LjpESBtzyv0jzjWQQfKIxgBuzu/pLO+e75L
/2aE2LeQU06U0dZMw/jllpBnHRcHGqylKlP3oQcbQaYCC9O4Ec8YhvlThRielNLF
L1YH7HCzTIsE+GFoW10/2nWO4G3HsTmLP1sY0h9u0ulYAyqCb14G786OlwSnOiGX
6xXP6XNbpxkXCxdZC7FxYlq3dhLIpZ/bgKl5wvrBUmXDwJzA5KvaDu6Y+05zTH0T
pDDB1OWrf5dVqVQwPYj8xFkRMok4tG+rlMVP7jhBi7ZXL3ZzXhpYNK9hIFQ5useD
DfntdyHWzH9CGB3JZikDds///U1chuLKUYCUOAWc10f5aNr8wxq+7BgwCHYNjm3y
YqSGkJBP9a7/cQHNL0YY8OQesSih2eyD6XlVYfJfgYIBjg3J+oT/izHg1ldAPBfZ
oEAbF6C0cElpoVwtDXIM2kOtz0dAUZT45WWypx2U8dJ7q+p+fHr4le56t54+yK6i
aqT1g+WTp1t4QSRzG/gfEFHy/y6mP7ZnY7pxpay+CiSc1a+FNgJVKxHnpTXMUZsl
pWvXuFu8+jzxEKKQLxEv1sJcqXgDdbyG58mKIDHksYbpw2d7oMCnDJH9EirO7sLL
2Arnx6Z+LE+L1q0Davs0fFA/W+PQYyVTvyFIWgNAuLL+6k2ALWQePIRGYspYbSxR
ZRzhUPwLKpTLJ0eOYCeGPHih7WHiEYLZLzVKHzgz42GZkkwls899V1Qxre8kMuo3
sdPUnf9f0UpsfyeFKTJ1kFxk2HmBTgyCZI9GmKDks9zC5jj8SoAwNTwkJujKV6lT
aHTgLLcGzGXkoETzlEF9nv1VD0bIoh/6zatOh3YaeqCabCCesduOT0mV63EaoUwd
KBBKZY1efTf9ZRCtNokVbNSS/PfqPx8e6M4M0ymYTtXaxw++QPOGOmTUNZyugNsR
chEb+U8W2Mw6Y71zzJ9l34sJ7RHYd9j0Brj/HEWbCoOLQ+LYhTg4VzYIvYF7Wn70
RFl88aTXD/hMet3fh2jvKreKrB2mYcmbreCQOVf0E9rJIFs3eVY6EC66Y7kEhOaX
oqf4Su6lL2zoIuiI+ttG74ZBzgebFyvfNcBIDA4JgDXkFVCy8WKjpfbjWcdPAaye
0k7WAhr3IYuOpLkqAG5OgJ4WeCmweE8Z7qCZQl0/2eRS1/jvdZt5qLcZVubDwsyO
RDSByVvVtD+0TiD3WXBVsSNQZwc6flGqQVwraOhURqOWthZYJAe01UXP0E2daWXs
tcKCNFEDY7vcmt/4HxwUp/BzgoxgmAZ+AvDbbCa4RCcxqGL6H1uKJ6wHnca54bNN
KbS36QIA9An2zzoNWftHYHVk/p7tFkbk3p1T4WL5XF6H1GuKFMd5W9R5OcRodANp
BPwsiOCYga7oIzGPAKepnA5gZ3v7n9IOzkGly9VV7SgRewtF4u65BLOs9EVHFBdb
+QYdjrRnk/F8mhKGsXq7ZVXvbsF1Phj7SddpFOyRD0w29bwuJ0YpnR4H/msZTDYj
C24YGcMar4fJZg6M7gZcaDOL2SpvdI0hyhnanSgvkuLItYgtCVJsdtlyh8Mt8udp
Bri0aZG0fjW4snyo8Zh5EjwDl+Bdrddw5tIoeDNooAY2Z2CrLbF1LItzunSyqCym
m3l1pVjTbw7D6KIb2HIjg3wHP0OrMCjOfRp84orJpdXQ7OwAsZ9karZL/mDa56oN
u69S2tLtlevSEt1kWcGUx5KbTd6vmhrhDt2mZkjK8uyAZ5vpNRhQNaKeYOjOHJtZ
5MfbF3aDn+Yq3Z1TumF3FpI9UyN78uzDBIpIiB68WbJc13HevGfh5HNgrpnve9Yf
80sPw3zNfgDfJLuWQAbSGjXTe/oW+W/7eVae6gsXslSHaTETZ8PIybjhJgqYjnP7
aVVEuWBEY7X6TL0sLR5aAoxlnQpJKJK/eDclq59jCbhKW3518N3gHLIZGbbuF+Za
jW9PSEcGugaP7vCOCJ7d1NJmL0m5DTwPEkTHS78NMVwWDXdVnbywnRmg3XsSkwKw
2EReIx/YaWQiDZBVpE8ow44TfcgsqwYaiCHjAEHIw5iP0g+WAaBUHCqWeXvR7ZDk
jy7qUkFEOBghY7y2c1X4/l8rTzK+YdcbTPFOU70w+NutzI9JsW992QIg/MkBtJJH
ykSV8T/vYnWHLcxGYAwqjtBvyttce0GPgxr9ldEFQc9Y94SfNABS8RGS8r9mxB0O
BUlnyzLFebQNSWis0sgHYbiOsYqZ4bUxd/9rcaDQoPLDKJwMrE/OfZSM+JP3o/Kj
WAx/5yi9mG9pk+6+A1URu0bLPTbS/C6rl9u2HNWBUVeng4mag1VD+v4FRs4yFHkL
kAt0ydcwxHALBLyW9b9HtfNchqi4YFkAZBAomGujttRbrvM7jYrMYHGquU+Cjadj
ZrJDGweQ9eal12iTVQbXXktP3iN/mskb4ktivdWwopGXyZZQLbsfErLdZW9ANoKq
qtwfoE8aaR/jIkL9UqFzug7hoDPJczzZBf0epSAYCtI5j/ThNMyqFs6/p0Nh5/xT
T1O8jXwa9jD8m8PwKZCRY4395hkijZi42jmOhgRGMk7kw7Hkgb98Y3LtZJCDdZTj
JaejdqIzrfSF/dMn4RJLqOt/EgXk49OZX1TbFY2v7dRnmf1tA3WeBcxTpZylqDaG
lO/LhZU3Rx5R0aLxGFMnoTKPriNgjNk7mu7fUSS0J5cg1foj9PQNV+axx8GyfnBW
pOeNmMSDeOFCNNyc2r+jHphycG1ezJHZ53Y3Ua+dzaD2IlIf9CQABmNIyjWdsu32
4rawc6qxJfU7JLB6qLn+KJwm8ngKOY/q/ze7INN/+hyV1AGhKNyyaA1vEGwgKAx7
kbqK6ZX/QWw/fwWyx6OZzBGAUqUqSMVux1b0DKACmTKdOebGv5zR64pob4LSpCV1
LBaf1PlN6yIyvErvfyJnWwVGLPI3oaNj6umbk7WUAQi2T5N2xdprIszoDDbg2YcX
V/oH3AhI9bjhuACG+ODRXN2fyg9JoJ3Q17iI8Kf+pUMJEw/+HjokIXBJRUlPvLle
On0bIPepBqYJAA2QL3eC8kTj//cz8ahzaLXNoMH0ZRLfcn0i6H1rEGis4eCeuxDZ
zpXqizddASjv4Q0bIrem5blNP7SwNJK7L6grCH+MGDCjiRUtTFeLcbTJDhjfHgc5
zbrYSYQx2vLoMHDV+DJXq1DUdxAyUJE0+ctB9jItGULAPR3EDQesbI6yI+7rE2o7
VAKTuEvGgDdUcAq5nJwufHyv4Vshd4hYAg3WZr9j9jsKlEyZ1tPZAXtk0jyB3iIT
EDlIRQgGPXiF9nB3kk6CHH9BR9hsOSZsrJinbIARVq6O4+fKzy4Xxg+Kv5gRT0BK
gJ0JXZF6aYQ7gMTwwwYePmMjpU/ViiYt3GO31Eo5Y6FZG3zTQ2gEienE7ktbm8or
9dxt+ovRaP+Y49F/EqGrXiCgHoZNtMUzjtCYuVfYJscSTTGxKy3Vt+RUeHrUP4BV
zuVGPXiEcoNRlvOQ7oyHWFwwibWxlU156k6c9Gt8oVQ+mAUXRFnLq8yWflaz9ciV
uNgvCEdk/lQLtdlN/Z5b9M+v2c9krY+CjqS6wreZw0Z60g1QNXxRXSbcEGh2zHiu
wdNgGhuWd+fqM2K36xy47VNgR0eHSuSVd6zLD57F/SFwGcqUeraNxRgD0+Bl07rn
HQwAL2UX7ms3R6Kag+68hRXX7CYeGvqv4H2qc4VfrQPgEsEGNpHRIRIQtFB7OTPF
20SxTAYOl68wLN3MqrSO0drBW2vDD3lBakGswxQYqOFfGe1bl0/og0vYzEdSaqMu
2r7WpD9R/r6UMZ7Cb9nLMGiXKGFv89Lb97s5YdeeoT/TLlDYUjtLzVnSqJL7EYlo
dYJ4rHNl+o8725w8ZTGeJVmsT+EG8+RK8k2AGjuPl5wKi5PM0Ps7dF6MB9wUlZxI
QsuRPG9WaLCYJVyBGYJm+yFEGwC96QnZegMqLnOVnqbFicab1Lc7vIq9sKxQb3F8
Z/2/+SxlC2qdP8H6X0a1zSUgduVAdUGNfTl2UpYOSJ9a9Zu12/WNCWHL9ZL5Tnz5
DcgAM0SI2VA88OHqZiVaw/ekYNyQPr5PzddpVyStrgPq5bU5HDnU+7W2u1Dby+5y
D9eL1/Vc6y7CxfD5Z7ki0xQ6tAFvaHrWlv0Mza8grGqcglGwQcBYBVuyzDHs2nm6
r5R90Y1jT6ziCvt4saqzikysCZaFrH1rLFmU0vuVitjZ4XDFl6RjJghos6W3x1G2
x6iYuoEu62qP/oFC58kXtAcX6rmLrEt3UA1yT0gBGFhDzBf5CCTMpC93Wu3674Gb
nWvNLxYotKPQBNkjt4jaaRV10bPsusk2lvXeL8XICdciehYg7yd9boOPRRIopDQQ
AwlAUFTABF6YTEygyZuGOdaue7QU6ETiKwOE2SKdv022SaO21+hfjsPOgXzX/drb
I+ZV92U6OXDRgrfLp3R39+VD7cgrDLcF9aTJy8wcHfi1TESOdkHorWUpzGSealab
szrcyTI4hDRQ9MwOKHy1QPYh3Kvz87hZ9U9cPUtI3oCsjmP4jj2+84wfhI4w2E43
3QReoH3RX4ICEZIceLuiVOPZhChlzx6TU8mBCytcLe5M59tZiQwDn+gKunION6bP
thGoJbCSOWwY000HevQXJPPowxRlAfL5V2rA0YrD3QHkpaE6tW7FkZod91cokJVB
NzrM+HZr+O7NxT8RDOQWdUABeewZWZAaY2RLp4km8QW4t35BbwyzeM91aacYgNB5
sqnCqhJ+8d0vFwJcoPn5PqESX1Qvv31q3H0qJOLBMYrGVlGQOWInrJo2UpImkQ+1
YyMsCTW54f7Q/EcBesCOyS8i0Z2XrlEVqTlBnvUj6BjLCVXV1HaIZiiKfpCLUuJx
bWel547HfY71UueOf4J7Dr7GLaeRQQD98MaRgme+Mw0gSg8p+vvM+KJv+IEvEYQa
MYmSRofnyCrazkUR2Rml8sDpopyjsNI3GpNovFw4WbuWKUL2wZ6/yE0kBp3UlvlZ
qotW4BN+QYOnFVBDo6NzHr5AFcuLptGoTbqVp31epdciVuM+wyXwK4vyH1smtpAg
9BgO4kSD32va1jdvdJ+FKGGZBxZ1UWFnIVYXorJYBTTePriCmJA5j58unOc1B1Jm
ith7vNgZYR+eNoynWabsndya/dS5Pl9sObRAqUcxPbwyEl6bcB+uEsYEUHSRzUVr
pk3/1nyWCg1v6hvrvbHXcaofT/N/Xn8esHO1FxaHBmk0G0TtVptJysS/2bkYMU7R
pknD7v84aXZKqrQDwCuHv/ZRI14Ub4RmmQ5Ej4Nlvk7IfPoE4oEXZdxDxYrIjAL4
cAAcSapPd+7v5gbc/oWfs5sjhSWVDWOEWlPhAGLsJBiglMCchCZx4nYLZ2OqO1w6
t1RqHMk+zHrwGkUDFJVmGaV0v+XZfBBP47cHkZ+0hUv8EM5rhHYOHXKOEfTgs+7V
WyM67+IzEx13259z67jK2MORoqpK4lnfIOrwhibUh+07BfVjdo0yEco9jLL3MbGV
zJYH4Vqs7ywSEjWXjOwMXotLQTFw8vLDts4hZeCDhpNs8LHmOlOdWg/2tLMU9BiS
vXOJQHUB/4LjCwv4QBSlNPxmgmghkJ68kJ/vnjlbssLRBptbAhxzmQSkOqHAs8fn
SXTDigWsZtX9NKhRCX1TZgUbuIeT7OLRHSOQZhWBf+R1GtmYv7mmYq4pKQxwNQW1
GdndEFSRgKsp9ZQbHRTAuD5KpRyA6WzJN1xTZO6Ye+5TV0md4vImYiSqx2Wvb7KZ
u4mwjC/nTqkLsr/N8/hZEv0zeeghL6yADDyvPiGl17DENiym5z3qdR26+835yBzd
EeAZtBN80POYDT+TsAyusPTx9gWY0dBKczTWonPrvDDNYKr+aoKVVh1WwIzLnvsN
YTUsOW5aMWzxx9TNz5PTWf6q+Xc0z15R8sZ7KWAEclwtAbsSdGhWkDKkHlIP7tXi
aKObr0HkTcwJbntGVLPn/vJKZrjGD9XanuhEFjeCnEXrnx94CbplKJZWIhM97ZLL
zeSsmCkYogPF+akhc4a8E7Sb2xlCeK4gxsQKygmn4RY03c2ncW0YiMZ/TDxWWF0M
zmJer1OlO+ynudxakgMIu0jn7LaUqKQ6oUYw4suvq46aomxbmohybZn2JsLLtb6A
nTCpz0OOSit/+yGpXg1Ps7VGEw8+wTMCY7Tm7tKWxAj5tjiE/71OXzu0ouUpqAm8
ihfc55EKI4egRHndYcVUF2L4xhy3h102MnE2KJAL+IVsALADNBJ2KQ72doC2NHKN
OcGjRIag6YTOeQ5+9fUaQwhoK9/5VD7j4tPrQEfcKhqlq/XAkhytLyVXefLxbJ3s
f0J8sDMqjDe8eLGKFEfq3bD09VnR0AyTztNBXqMLF7qai7bzjYw9Nir6KbGfX2ZR
0K++gSGLlXgfaKIdIg1cnYP+FgtBuzmPesyBamFfo5hGJaGskpHkZ2cxsuiGX4EV
lIoQ2Kvv5HMI0DU7dg3sd478+dDMrLriVqKoYYVS1om/JlQ8/eVqwO/mABPIb6SF
3EwTKMFL5L8iWhlndCY9fsia9pPRTdnuYvyW2Vf7Clz+KQjCnz5GvciSw1YsX9fp
PNy7ymS6vjoDPLLbaqRaAsaaY8b/Maa1PQhWioZsf9eTVnmEL1p+ek8tswruXLDG
1BiBzkqsKcE4JmLpZLi5Q2G5szRO67zyiRKsfeWlGlIemmL/vZXTPxT0KMgKQx8U
iszuIS6R2CGso6w0r9ZcjmLWqsv1/wVip5rDgrE9w8vLq1vMvr+iLkilMBCnQB9C
E3YfUJwCqleiRcV0Lx3QRYyo1Krl+RtKeJrx25uZbd5UOwvuwQqGFJrF9IjTS1Ve
Vd165nhexAg3koppE9WXulEhhL1jYmO5Zdtor2ZzzXDYHTacLrbuilUhP242zDPc
bw8Qe0YcYxiHXuGvFgdMHTOtSihRhNBMYXnJB3m90CgYeCSi7kIn2VlVbdllAdMY
Ub3OKsUiTMYGEHVJ8GB9j3b6/HsXo8xOjkIG3Q2sJmT+Gc5iYIA4cIr8N6Rp5329
/8k6nSkMsAs5gJfvTT8UEyRIZHZLr26wu7YD2+rdjoYsIbN4lnUgkBNazaF1f0uf
Fwuae5OYea90t6nA0n/635+QGJ0lg+jedLj1fyF3TJw3c5OmTF5Ja2jWYCyTYuEg
WZIUSD4tblWZYGBXH0h68Hx3GozSDv/ZECPDv1fodcsJEXu+q9VeykmDCMIZHIua
jLLFa2V2xLukMXa4QCMB+pUPUP6dLLmqObbKZ9HRFFDAec/GjeMcFwigtPusmgE9
e9Y03J55Y6OewlleuALho1p+DbRqAOP2H1m/lu88PMN7EYcHBkBY2ePH9RX6gNvq
D01+wjnUy3bI+8zCZfy+9/Fb95EKHR6eGpD01ZvuqqLGUocIZuVhRVl/+8/GZV7N
A/X/BL5fGqXuQfqk56ownwAc7gq9c5p7w1S+nRCeec/zqEv2NkfNXbBGcFlpa5FI
>>>>>>> 426889eb8ce467b9c9a9f74dd4af433c5046285c:deps/flexrio_deps/PkgNiDmaRegMap.vhd
`protect end_protected