`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 55056 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzglQtoUDWVGGBJp5DpeDqlkq/HZ0eSQf2P75Dw2DfRCN
S5s/UhPjkn4R19MzTPGTVRNLP375GCPQTEqqLTbhZSIW1pn1Dwbht3htmcMC99X1
6TVwDapfzVGrJXW+rb6cjT7xxYfM9EVB3t33a7qiABvBSplqgyvuTHN3t4P1VVUS
kMu7oOHU8+IgJLVp38SspIHssMEo40ebRWvYaJWBjIH4n16S6ZHU/cM1kvj/uq0k
i5cFNP30vMKJduDTMHoj4yrExp6Hib8XqXh6RbsyCemG45LpaL4RLspI9lG5PP8i
koUgTZ/15ItPZEIUXjvvSGsLbzr7IvDsvdotqwnbh5tbX4UgZww4retT1PvY3al/
N/h7F1EemrnW3sAyP8WQ+LAnl6fRclxYz7j1MXeGHkPHDu9SfOSCiyfMjrNd2X2B
4tlZ8WAflNTm6sUYdUMi4REaXPVhoE1nls6nTeRgafeH6k9NzZ7DIMdyDutEasS9
MbSsUGMx7T518dT4lbIXc5AriPIwHOPDpcok2mh+nDJWTVKhFu+91exJN8EncT0C
RRgP+Qydy4/+O3CCw5Goprfa18r13HSRih37ZQCJtjx26gQjTPDH/e25IpWzFPd7
TkF8XuuzxVSkBWv0WRcE0JUfWb+crKCbYV0nviGs7aj7vUFcWzIoq55cdntbYLgb
PitHGQem5vF6T86mjtVIHVOu/khDC89oOQMLGvQAp1WYHJ+4fzAwDLVcbKGGc6+G
mVzd2TkRJFW9SUYteazcHmM6l5quHwqdTeP/MkD4r8JlEvDqe0ikdKaPLeqDqNkl
OaYtY1DeS6setzmj5OrJiuqp4/0Df5wgneqAfeQwoe1x1gwD8aNFFUwlfuHv1cj/
U2swMVUlzbnw047mzsvj/wbaKWm3X2/zuGw0JOMFbrhkYmkygMqDFV3pZ7iuZ59D
QejilM47XKJs9ZnaBX7fFWtwN6mCRt/IzedQ2Y3VThb8XfKx6LsKNMey8ieXoQ7X
dBjt9D3A2GQ5MIhjQ0LI20bylAgXOy3zzHJvi0xBZsJY10YI+Ml8F1uRaC/LTZHc
Mwgnb7NnfNlepSXlRWBl5o+nbvHOd93Ue2dzNCxo/Be4CA5vdXp5eWagfiLfyquX
Q4aYfPf6x+yrLZUTHV2Q8bqRTrw2ZdsG8tEsXlCy1zFRejzV3MdYjTd5D9GuE8r7
ZbiZvq+6+Yw4L/qNB6XElwhHuLnxcabE98DdS7/ViZNLWBcbKvsOS3Pf7HRNB52W
d/qw0PSrT0iGudBSG1b0rXawabbs/e24UCuT3MVdPAS5ACVKanAkY6Iajjruzvmx
7aQfNTt2GhPSppJY0l+CvGQDmvTrXQSHa0hiC/soB7Li57j2oL6KY/0dzFTK8NMN
VjRCseGZnF2SK4c1eqA57v72yhzfIkNZWWMbVT8LQAOPK5FSjMt+WZ3aMU+XSNGu
dcnZFt+l3MJmuLUWpmJMo742KjU8q32JRAhJDbOLLxAbcnQfi8swTPksXCO2Ia8M
Vms7bANUv5xzuzf6SlVxNJ/SdtVQdx6KK+x9vleTUYevV0Uf1a/F2udYtfeojngn
w0CUx2i+bsPfhR5mtSkzp1h20SgmCQgh7GvcN2AWwxmFnHJ1TXwbk8yNtToII8gH
THlXoUhNlUyb6Isc+j22c+D4BMjtU9rKWV7Wa+0JS7a/lQ59V8fiYl42Gx+Shv9c
ZY28NXLc/Bf2zBGlHdIYQKoB08MTMGWPsc4Qz18Q9Jy4AjwAUmKjhyCBgUf2B9Hf
i3AfvSiA6dqBQq/AX6992QLp7Cc2kDNlmpARM8+SxYKRqkqkyI93LA5RzdUQj1VH
e8ZgycCZIJWJuDNI5a7UlIQdgd0zBR1uOR4LNpDg95KwzFEYT4Oywy3/LQ2aAzjg
TNMbO75fCCp6CjDkRtfaYN/DAMUqI8S/oo7mIOuAZysO65B2Co6K1F2i86d+jEiO
30wehzUkX7Om9auVRH4wMn/fqZe8fVvy786fYiXx3IW9TOCfuFo/XoUKGjs/tn7E
RzHMHnOotKXwk5v5Kfj1+RsRxw/XYoQOgRvYM1EHrAn2rdFToO1HzheMCCLPZRvn
HAbWfqUng2V3y8Gm7/rtiWpXZROJA71g/E9PkEJjHzjDFA2C0nsNQEoXR8yuvfGK
z5F5Lz6OBVZEDOAH+zQCNSbX6nT/QSLNMeUqqhhv8Rv7nTapQ2/OPzzx7xnaofB3
1czFhzPfTeswdxa/vf/GI70iEfiqQ+qgUFYMnWxxx+GVOulL5Tcwps8YjVXpFh8A
ZgVdrnQwBh7flPSsgmRXk6Wqb08Qc2ZOUDtXR+5sx0oAMqdTXJFeObFiLg2qT2to
o7YJUVEs2cs5GeOJqbqzMde0E5UdYluVNDsDV2Stzx1D58eMRc0jnzFW49iML/KG
z4t/UOMUJGAzVKqAPSq6UN+4aijse91PzPzKRlyy7QTQfxRnZMbbrslYor8tXrCl
oS4Zwil9HQ/7/nh7lB2SZF4VvWaJ9oQQu6ieY5sU6n2ZJ2q4QDN4zDg1ozb9zUPG
e5n6YuFWfiMY4FVTYb1FHriHBnFZHKTXTXwjHp1Gy6T/n680pujcWtbRsDSCRPJX
2GiAcn3TchTgMqad29KIWgsYGMuwgzZ10d4NwP+1Woc7vh0nomEVQZFnWEcNNjWL
4DQeCLt+lyFE8JZtQJ3ASvEeKJ9iInuVFDw/y0Qn0kwvjeQRCQzCkoKQ+Y2yz53v
b0GnpjEMBl91gH9zcxFd7RPUkn7Kw4qV/vcpHHFeKnbR/KtAgYco/Zg+0viEz3em
A3K7vbAaCEkbjSMdCXkLWd8ltOkhu718f6OavDGl1bRIrquxu09OrELtOjJnVRAh
Pbwy2P+tLE9m1uaCD/EIHdA/nPb93nxKzM7Aljq8S7E2CUuniLujRtgQiwfisV9Q
l2LDw2EGhrH0HNZ0hZUpMlSBK1ucsNsRMsaRVs9oo1c5gGB43nfw6PjlzUEQb23a
rUwsn3nI94hhJFQnr3LA2MLOXy6Ufe4LgzNdj0BdrbkB4wYQct/2ypf67xFtgCAL
cCblMbmeQEyUCsf+4YZy8TAXGboDbSySshr/XFs1gtdv8mt3XvPdihpDsIfVUg39
JDyuWP00LPFb2LFxPEOBtVHAQjFwkO2/Dkbmd3IPz+eoFZO5CZNVlpR2FKAIMcBK
gzTxW/yv19dtDw4kUSVDWFFG8elh6uI3vFo9oXnTsXlksI5WJfWrixXBA9bQN9Y+
7AlDWQO94D3400f/WkAaU489vu0HBS4i/8r+O+HrWGmABosTioYKU3CA5XT6h0wh
eAMNIvbNzIdltj81ggUgvBCnJO31316jBSrn/P0AicPVCJiE4ArNSMwo4CL4GYWW
iYMV4OjVwsqKYscnWYgRnUy/rtr50rGuVOy4oDzp70piA9J0zlAq62aaoDbNaomo
mKvxm6WwFhSycRLESCuVMZDy7+aVv0a9l2cARJFKIOlMXLcOjHjGEKMfDvDrUuQv
5enhA4WACraz8mn04iJW9z4J7ChsGmqAxZ/nhCEhV8caRmAfnIV8JTePlBoUajXd
6sYUnYUL3p5NJdo3dXKQfbV5wFLyNp59wLv1qcU+x7p7ycGOzSTeMu2TKLvMuzkS
jdthVKj7377yp0jEGL4DtdVdmo9NSDQ2qTCpXNIdqLPqeelxoHaLT8tlDuS/rhXn
a+IxlhnShWcHg5XcQDn0czzuEgYT32SpC80cb+4y24XIK1POiiou52pqX5ymphFo
T9w0OttB5OU2k4TFCZFaSQarKpUjnoHs+rjWK0+qJEOMhVm8Fn77ZHaEjYv97g4f
Z7z5XOEL7/LPyf05PE0a73TPIIiQWc156/ijL71hYnDRksnFDlX32Qnm20qDU1Lc
cU4ohITu16RDp0rxMJKL8HEUD0coMesNMyulGEOA/jvl8zc3u6hZ0XQUlhmzC5Uh
LJtCMDY6Prqr//CN0Psls6CE2bOieu41YVnPVoz4hsGHHX8ejPrAbHx1selqy7gB
/YQ+iRqKIJhkFHM2LourB9YSmYTj19z8a6tLSuwpzT4nGWzqSHiFXsg7TrYgtMd5
dJcxb4/MFY0bQWEtqaPKDl79/Ofy0L10dsTJW7fXjf8SPY4ZevZ8ywC0YFObUx+j
6eO1grk8+SJcNpUpAvGkuiuklaAj3tc0MMqF2EQksTpjvrwP9h+GiUlxfpPcc7dl
TVD1c34WR7aYlDQTAGKL96h/x10qLgl5Cd3Fdyk3M+JMblf5Z7iUoWdbubjaky+P
PSEQomp5eAgfFMGNvpx6aytyGwM6qnt/Dh3qN6/k/DYGEM0iQTCn0sXLu1uPwlAQ
r4ahbstCCI9EyRoLqxgv9utM8r56xKmxH4/z2dr5yt8AFRJZbaHkm28nisDnmjPM
PlLl1lnq7ca6oux58W1tgE6FHpDW/KHP5iXL+IbD/H1x/4wK5J4280W6BoWSxRSz
jDsoOUrg54E4VQ8kvloRfGCe5OzmUsbEqhMKfQr83sBYLHl1qUbAHbzTF1FLyWkQ
hw7O96mJ56qDmPIGcXD/p8WuyNpY+JqRuibxpgQhUEvB0gC2qDgPWUxS1nYX7gyi
8AtiHS86HaHNijAoEIPy+wc7pJWD8eUZYE0mSYUY+fxDWt/o9G4Iq3tFdSwtJzCn
v4HYOWUhILpMPym+cimgCStpKzmp/vyoJmr3GTeriBLLlFustiYucWfrVETLPWVB
fwmGwcHDwK6YRjGVot+TMk2YwD7czh0acdpzgo+GO+f2wvHPOna3bYfswMbo6rE8
K5IYLekIHgariO7xktKQIiDDCfirz6Mk4WbTwyLhD8L3m+AHqMpzVyRHIVqSMlhI
SvzpsffvjzLeSMq6lN75VpEo58qaHRsBCmGss1qJcf8CjcfLa2eFwn4VPOLR7MwP
jTyJurgvGulQm8oaBRt3AX1/Gk+DNgnIdqEc3JXqVe0Y4dw7QLDYOzn9jCI0o8C7
C0DtnFlrz+suYvH6mq+8pEUcv5DntsXWq2c9/2EBwvtooSCZfUMu6eTuODmJ9Crc
MxOQiwSAvLD6RnNNqOQD7/DHH0RcK68vz+tmMJ3GKFvSG6+BxzCnstsXiy2TmANJ
i2mYzm3vxo0RnJ5/vbjwCIf1FDufkmVxImo8ikN9mp73paWTzg/TPC8tGejNNdW5
YbapeFHiHEhD/GfCQKL9lhreUdul80TUbnvGo2ItdQeQ6mKZ7wSeCK7I+KGOSAzc
/LDiMZJvtzrtbXvUUz7TZgb1dmOWj+0U/RePfGFP757YBpJGVnxJ1yy97APe9ZpW
3fhGnogyCIIneT5lipC4jJswGfEA9B+IuQAfm9Z2aNPzjJNId7TcI84uyxx+RDCu
2fd2B6vxh548VpM30d0ztHfDaglo8wYqUUpnR/NAykbHfUGw5xH8T0ENnE4d7Dc3
9sI9y3wMk6OWMIILN27nnnfXTG24MfQdahjIL8IiyLnmcRV7SwalipXvwfx1uTPF
uCIDM9mqfJOmVjytH2Y8Ncr4R8I4hoLC7wk2z3aWBdwEtjiw8+eBWTiZGkjZIIJ3
fy47J1xm+Cn8FbMss+wK9TlL8KGC7aQN7aK3fLq9Hy2Kj4RVl4zzhKJOdat5jNit
SaltST5kzEGaLubA28AKhoHvluNfE8m4/25V/vS/+mG/89s1OlMjZz8MOul19AuO
9pr+HJcMPZbk2rk2ZQFdtfl5Fxg6f1mo2p+9WJtOFbSY1OQOP/pnSA84WrCW16Mn
B1+5lAehjrJ6H+OxODK8R8R0v+Jof/6ngRGA0rOg+iR4dAPjBMR3hIMjv7JgZkN/
389yhgwPBQ9CSDfk83RpfCFVjfzS33a8nJiLCFMLT+th367eafGc192GuBUEgj38
+9a9GkiG3Z3rYtUhWaQlg4sLwXkKUfbW8QXoYRmVJp6eHRv4kZZkOI9fipVpdY+r
hfHLVzNORD5JbrWYoavjNkLTQo/p9KgSHL7HqCtLdMNdPDlXQQeH38akB7liQafe
PVtj6UQ5dzjanS3Q+XY56dFKW2U0NfooRZ3Vpqye/WItX7ZPal5zHh56QxCrR7xD
yqxRul9zphoh/GJBWdNN82HhCwKHGvwwSpYO/v4xpXkqic24U5iUYKyQYHJjVUVj
fJWgrRuaoewh8QggZfFjyvwnqIV4y/uJ9jSfIShRDtHCJ30do1mQ5ZJ4r+GU4TSe
6KX0QxI9nwpOlPSIy7hIekDf7FnzlAtuIRv7AL24LoBskjiFNwE/QFNx6J9DAcgs
HTEezhe8JY9558d1byUDjjNpT9maUCTm1aBwLAWhHillxlLLfzwFUKo0O+bBptpS
xqjw6syA1E+dWgacSmXp4ovkoZ+7hUyD/mUPt22zb1+ppFOTUI+LViaKYlADAZHR
LjBk/Qx7aYR+QkxZ7Zar5on1O/gSYVNBpT5JwXWb3H39z2JhZHTzUc2MdUHLl7LN
I1figQ5xU9YTv72d23B1iR8JZHSaqSHkNet48vmDbRExGgZuV+o/l2GJHv3aTBGU
M8UAnipltCfQ+eU/u8n0T1vOlzI/0K088E6WKoSRNIaBVNTyd3uY5jVtzOpiSPHE
UMDKFPhqf01QDXY5LGDZK38jpkOfOasM2BErNUqUqBJLJ5/9UxVK0NChtV6BTOIY
OyyRwSUDAAzfYFLx+weVCFd34mbk4568MV4J8taQtR3iJ7g38WICqG0dxqxzSvAW
PxRPtTsN37B8raWANNA/nPWXfKHIU6lIkR/d85F8mkWbY75xkDyh2RgDuerhNDJi
34zY7FyP+miURkzQhr/kToJEL3gbSnzkM6OGwcksIuZhnx5RQ/LKlCdZ/KarPWI5
q/QZlpFFfwzIBg+dEIsxmoYFphEG7L5xFk2n1nU1ER15/GYE4YMMOOoxguT+i595
ji1HaLAM16VW31Z2/AL0xYyUjrncUzi4LGmOFbWXIjO+an/bCHNb9abz2sIETdm0
i/2qjo1z678q6xr5h+NSeHTya7mioh+sduZUdvF5r3YznzSClb0ywJ5atICBDfse
lQ5K64H48PZE89HbjcOvqqJagyQOrc/JkTzvWGxnuJRY6CPHiQpbPJERpVCrvMXZ
b3mah3N/OdTQmh17G+QaImGGmyqbyUz0E2gOKk14pp8+7Cr2NkiCoa7Nhy+JRtcB
WrzFNHcE94LOIJRzj05a8ZJ6gC3bNnG8kREVEsKg/huNAYMF+NNWEok/y603EkeI
mGnoP6nLoGlSjwe0zPqs8U0wIENxMcE8+/QHRK9aq9VMrdJUdW/F1A/S2e/GHrHm
ZcOVfEPSgAtdLHGeIAu+6EsV9sUFSmyjhNXE1flPRye/Mppkz561d23Odq9iIDJS
C54pCX4FLckp01JMMFWowg6Gxw7WjDqsPCgPa0hCCgEV3yNLOt1JvagSbd4H8p/Z
lcTIUdqqF1gqFSese4+gZw8WAWEE6Xs2DYC3RDRnWeVPTOIpZMG6PSV0jTju5vA/
U3qoOdE0JgDKlNi58sGDtyTZZUL495Avm8e7e4Hk1LPHUvxOyQS9k5nDpqBv2A2c
OzJhE9+tEhhu/+7x0IbxL/wY8y7VHD8eSYsVNuw659dgQvAPpqPKwZIntdfnTXPp
DPLbPrYnm/whVqC4bzIpzvDhVjWNVv9xUfZ2KHffepGa6y6/jaS9r4zAIzR5m0jr
mtf04vhHqnetZJOEvG8NLuI2b2bKisP33S6JBvbQ0XVkgGD7aLLQDFa/xmqGsrIC
KjO6opWHm4kAIKxRJizClOlMQTEV26CaHMQERmVodzTVbvpFBsmx8Kjr24g+mIxu
O05tDZdsN4mvikd3iIeVvHiFu9iv7jbYXNH5PXosGE1l1XI+Wz0rKiyLzqOi0Kr7
ODuptWiF82N95JiCUQd17Pt0TxsI4RnvRqQuQlBaFvoF16jGWJH1ARmi7vPEWuVl
yZ+d0IRwmOPMe3Pi5fzGTS68WJNZXf50BbogF/Zd69iw7KCTaGLNQCNQBWFIBHl7
A3SMfevxXLWHXcwUyUfwq6aK334D/ippg3awHbdVIEXIuFk9ELo2XmlBRdT2KyBW
er2XGX6ocMwBJ2oIgOdLP8/a/ufLD4BLaA3UQ1SXcPDmSPdAfpN/wgnFeQ9eGeli
5riyXTsUCEpvtSjQDytrIGQ1vXivK260+MO6VsbewB9e7lZma0qs1nx4jQ294tKP
gD3A0BP9ViO8EpdmlidqsYZffxLNBw7H+RPw6OJ2CX8G3JCNqmsbvnm4ud66zOmq
8JcMil8L1hfUySxeLXALpwRNo+wKClw+hhNwNBRwH4gdlZEZG0S73mpiAr97oFvW
0Zz/sfnlBNBo0ZkAW3hR/eBAssgRQyHaUCXbCIrC7aKbN4ARBf3t5MH+4kEAz+gL
oAK+sYyOGdHB423J2WFJxbyMVqNtNnfrl1K1Dq/SNaWEhoqnNJypqQoyK0GRXckS
dlIsuPs3XpsyGrjY41h3oBN57cpST5akhtLr0GQklFHPBdc7I1UJdFDlfQpYd7+k
vY1hkuvzYRozaJfa7LXRQ65wNAZ4Jl6uaikpM76FyliqgZa0N25M9+v1LkRDjapc
GuRfg9aB/RETTS3Im8c90FaUI3+JrjeDalWzZpbslO3sGzXnshxosVY6fSNW/G7w
iy20VGQBaVGRyAtX3fcK5pGQYLpowQEQdfvU73p+V/QcvyJ2qsxVFB8f5YGPURXX
KhdgoirhSSIoc3G177E7jn2ZAJojrDHmTvIiOaaSeQl6/r6cP6y6wkrACbfdcOyL
+Nstx32320RZ1JGYnh8kvB4mBc6B2NxgmBS+9cfB03LIOTE3TgQsdnn07DbSG/a9
J8w2iTxNMqV6vJN/wNNnQhnV9ZleJ7Cwgte4fLhoVG46ZF9DXxWJgDb+Bv4+rxTu
HCDxgkhZbTX3+DnlyNQUvN5G/4efKRZY+0FqZv9qgMIgEEXnbwqFqZi/JTo89oQr
Ncnq5UveHTn5KlFE6AnYi+H8AqrSF7+FktwL8rSx5Jl0vwCAMUJnGmBEk3jZIq14
MASgw/gdAIwiM2WMecuq2lD1ATna1qj9AcVVhlbfaKPlxZENUznHpXc/BndgGAEd
Mg5nemJZwA2qRBSIdg+qfGh5XoEIiJIoLrKXtZgxfAk1w73pEj97rIJQEP1PTw7O
FNP8VS/430lyBA1v2j6fQoFk66eOcgb35K+PtUvrywmHbssY+DP8wUQFmaYFCARc
LqxWMXjrqxefGq3NZhWdhp0ZPVLKSU0FRnyU6NniQwjoGdX44TZQDI/1wnWkJxbI
KS4JHx0a+J9mSf2i3IiLEWSpRRRJWas/DKMRRzjc0nnK0h00oDIc+Df5yHzDnizT
G1MrcwFpK8LE92OFQwDWq8c0unBws4ZiPKhsGRtlFSPg4tjKGjwxDg9mPa//kbK0
gZzXpVPbzP4jRrS90HKm/Sof9+JvvVxFSKT+H+0EvLmtZYJn7VoONKKwQUaPCJGm
SyQkN4CEILosMyRKMf+cA2cN9g35V573AYwlhF3Mb3gaJkqVXwhOc7I+Wg385UAD
065LgnWBkYclOEMf0FamVJxdScFnr5wtZiANKUhXKWkftwL7oBqu+A0q2ysGjt/7
PwRgO//VGthCoMp/K4AHXeX483LaEBfe9wTm/rIQw82g22CnqKbM+bmU3A8/U0Og
EXVIJSlPij21D+pj4EnxpfdJAY+vXWT5oPmk4CVCvg5XbqXdKIl4/oxyl0T8xCrz
Rf1CPh9X3mjJhy+D7B5Ya/YJV+CAH8juqc6+AZmtIWg3MaWOvSE7qDqGa2AvFlD3
nwatDXLiZYXMVAB0hFqGOyYphH5zdzn8esmOTeYr72D+5XlFzY9xReRKXsqwG+sq
7yKC0+53oz1eAk4W9FwsbdUwi/5QpZ5uNn32wBDlaqKflNwIt25DzjkSV4D6mvLp
CaSFs2bf+vUXtHonPIpnGKPluF3u7LqutP5e1+960R0Rs/hfQjoCmVfr2ofzuLFt
nhZ0+gNd7wSk6uF4WDlp63TAbQi+yW5ubYdnPrBWiMuY84UjjCB4hdncZQiJtJqy
kdr9QwjzOulxBsCq0+9Pw9cX04ntr5bk96UXCnOwAVB/WvgSQBtwqz/VtjtpmLu7
3hpFepGA4HtUbl/NudB1pKKYryIgJdQORTxyBkmxmtDGwbGNTfqIholGcYOCTZUX
5mRWOcufYbAuoqdS60xqfy/dD+8f9xKW6voXPbPDOuCPB1vHFpopF+kbGiMRw4bl
ZH4i8YgQdwjYb1ftIM2jm2rsfY3hilZn0+5h+bKX0I77g3iHb1tHWzc1jBChoFb7
+zGFXMZnwbQ2/DAhYp1lMBj0kURlG0CuGgqnV1H4RQTOYk7or5YTj3Fu0ql3GYd5
XhR1xWjtp2Zi+fC8YelUEF1aOkRNmpsY6LB8ayCneQbUbHthOG36V6HLWyD6l99p
6DuwxOakhODyTjqk9CEwbPmICmJs5465nsPYySyYCD7i6QJEphqmIO3TJFcX0+Rs
kLjIyhpcpKC9ikCdDFFSmsfuuoQQZDNcSMlw7UVVbNnXpNuPVZ7GuW+bfwH983iA
mPfq9mLRqfSywi3oL5pMyUcKbxitPj33pON6JW8FQlWbwH4+8fxIo4Ja1jV9BElj
eqcdHpC7b1j7235k1i5ikODiMf/Lrdnnw+tLr1RNMauKInXoc2eqKnfTZUp72S+U
7MvvOXatHT9+t9a04urHLgdmcrrfH51DfnoiXPdUpq0OfOPr5vSQMXNShf1cJxaX
MUHBBs5fSbJjWTVWQyZjVfmLUHaDRHXl3tk/VQ58PwHZU26QKYyxcqsiGnfjJUNZ
ZgAsuVh92mX25jlflOtamNVBgZhLGIvPMP0aZhoBmuEqnFvtwZ0SwTNwhLCLZCKx
hoC3/qgAOdeGUkHagCCl/1PsIQKkPN4WKNSBA9Y/Yyk4pOyCA6YWHLGI2qJZ5nJ5
V92SKdOSg08dfP8A/wUgwCig51Z4nZ9lGTu+S+ytGcjvIyGCr/o3lVDY8r/u9OPX
QCAGoNu3qWoSq3IBff/7atmFx1NK2c6Xmd1tCDBbivAXntyTt7hPRsZ71VmPX2WY
odLl8afJAj2ECjf7GHPBLIQjuJeG8fPszgxVaTLFqKyvmSt3jNgtnYpVNwHlGA0i
AbfoFXOEvIbrbcdkpijp4HaNIlQyPsTnlyWUAN3hYXjc9+9GNJbKdGbFe2Pvey4a
UOr229oYldlnece68q+mJapSN4ERP/bQD5lCyb6bq8mwp+HKqhxOlVpnouCh0BmZ
GbJJQFA11vUb6wh9jtSmzW7Q9rSgH20Vhz4IK7YgoMaSq1G1Mg2Hd0mQlmL4z68x
0aqpIYYj5J0fRg1pMSKprAdK9lbNeiBVtRQpcAGATn2/Fe4jwlxVmG7r6raFHnAO
bCzYgIjGi1mhZJK+Ur1Dbf+bK/Q9zZHTDyD1l4miVmwGWqS6CnTNU/i2AAFowxqS
qK3wUWtUuMyVIJKlul6qlQ5dY4YS90E2Pn61qO0jU3nHwxfGXjb++mAMJQRA/v4a
H8TnAzZlp9u8WSzvrr1v+uSbIHLPf7bnBkwm1R8pVtKuzbsZbxrXASXz2szTQyee
+k6nCUU1p1rRBj69W3A8fkhST+hTB1ld6i07maPZD5ac7Prki/bCRS+N8rdtENk9
zLBsrNVllukZeqLFx98YjmnQ2eChn/1WVtnrPJZhLtmoH+rfKwi8ZL0OBfe88Acu
r5TNtgzCqkUK9kR8BGH7jJVkhBKO8stepyeI3iQBzsAX+uQcD3cNATQY9gimo0mp
yzRsz91TFM5bIv7VX0zX2FCRikdbSn9bzopQm0rQ+MTkcrbov6UKLftfp32iiGrs
SePxyYA7BW7uZnx3wzPDAMyR5w0pOuCfKXYk8Zg8tK007+5faInulUDg3DYZ1UcK
DU3sVwcqcw2YnRD29A1G3hlTZlPsPtm/yRE08Vuu9oHlt6WytNg6TzfbcMmdgyHi
HAOZB7xTzT/kVxZZZJvM51RJGRXgXyLKtnKnd22gjl7/wN1fOzUnTHLgEWvsRPGZ
D7sCTBNCbHjGAtoMT5SbzW9IbChZGBzkJnRadEmZSaXHjBZwPdrvr5rDprqr9XX4
OmkMLy8fAuZfjLdf5zYa+Bm1e9nEWefPi5yHJTAxLbwvAoxNGuySgkUFGg3E2xqg
RxVFoBNarVJVJJ7ACDKpLD3cDuL9gtdVGSD+jQ4w28X9CouyaINuuc7krotBNe9Z
4STJvUSIR/1MzBgi5rpKC+B44ArstdItSq9nC3P4nsmFc6WPOL1LgmaoNkS/32Ex
5XRnWobMCsKKrw8oBSDimYCMaZ3NOjSbgUpPxUKkOcZoqj+P/BZNkgtXHG8L4y9+
xQkyoCp48TMpkKXpxnQhF6tiLQuYTwk74/3Y4k5G1u/eoyNm0Z6NDILbEEZBvO2Z
reiZTISbAbUhv6aHgD6dtjQ8O1X1THpaTBuAA7/iuYUKfIwOQCXTEcVZOtLE3tZF
Nop+oT4Rn7CrwjJ17/qDPyPFH2mSEQxZT8dBkIsDvXT7H2ltRM8eQ71WsYOdmsWs
kglZeikn53jYJJOS/nxCeWTDKmE7cB/9oWhQABx1G/bgj85t6yquWQRwNmjzO+Au
RC6u66A8Hi0l9DlXSscRmhkOSFXii1qqsj7FMugGVLrSiYQQY8jqH0Ejy/bWd244
LA0BGzv5BuqpONu5dnSHWA1fqSqm+KqvN55hYs1a3LLUxMesnZLa0psgnDpSYmYu
W8NPDq9lTZL5iqNXxOYCS/Gol4VoVqanjp/xruQuGpKUT3YDbMkroKjKBgGtBaPH
FI+THVugWdBJd0a88vMoDbLBXcR4vh6kL8PxbwPRGRLDrZElFfO1QlA2/CAQAOdp
0q/tQH8utRm4Xd4SVRfmUqk/EOvU/TcSwlk+uaHeZJf78D94EQV7FR3Q6CsYr80b
51/Qdq80T0GD5WZc0XHHdxz5bc+qcejPR77O9nTs4CtIIezREaVnBQDuq3pwQ10T
ahIEl3nmmH0RCvsSMa5HlzUqwoz9kjwqs72iPuVroxhoka9BE5hTNpY4iNBoI34L
4RzXwE/tHzC9g3hc4mXe5JyyKFg3auRsR1QSoO6/ClqORANVkwzKoV1GBNKHEyGK
E1ldWiaa/IU+cXTrHmWgtjo4rGYGo3dUTFYQWEde/27VnwfXyJjeQ9jZV2e4CXK/
z41XqXJ5/ieBUqKFU+6016iW5uiLP7C7mc/llUwD3VTz+8aBv8Q1Mu9wIbjxMsf5
yDED7j4BxrpfYkCqy7X4nxZvn30RYTmvimL0ipD1XGA62zYDSssK9xXt5p3wpeV4
c2S5nDR0fijsqQUfpfX7FZnVzbeBMygTjGzgBpsoHTY+l6eFoH0kk+jxG6bmgNGD
6b8PEFCQTJMtLAAZ/pROhZ+xxTzC9tYoxJX/OD5Zr67VmKw1UxtPbVyZg/hp16RL
etjXbEw5A5uPecoVKtsRIfvRShifp1MQwC4QiLhAvxYTawKXsvhCcrBEmpToVg6F
Ua2bFffJyE0kaSYNNfyirkA/CxZuQ3w9ESrSYL4M/jZJCzc9ldlMaVU1AvzFN5fr
8QU0SdmXV9xSb155anWytas4aXYqrY1sa5csiY+J9bzZvKPFFdiaCu8PJ0Tb3y//
K8wv0/0QvOl1OhVO6WggR82p6yOqFRtDg1BLNEmXOx+V2DZjcSeOW1HFrl6lEWN/
NUqbmLCW+AXyvq1zP6BCAuoNFlWjKQkPRG1+iUCTxt9ABQXkmiITjMlZWA7JUHNg
TqBYRq7auBzGEpQMK9+UmgLnraXo0T5VJ9Qtsr7+2d0+5TiLFqICPPwzpyfVlgqL
x5Snm799kWPgEi0di251B//+ya9GmdqM60qXtRbNpMPH2CjEJwlbpve9SPUMweZo
ZLViDaT8dCO3DQBlZ9vUu65ty9cJROuwP+JM7avadijsZxVGApqecBRTSUO/D2Vb
SCzD6fRfAqSudVcu2pljcAf2cxwNI0/nyuutinEWRZsrf16zt3pVT9FwkgBdZc9Y
6C8HTnIAJULkp+o1j8EY3vNCA6qHeZP40OZa+TImASS5laWu7ams0arPADKeqzAs
ISa6usfeMCW5VU11ZgPEwh0yKwYveINLRUZ6sX+ct/zK8z6z2qGJedNr1W6Y0oXy
EtNDysUVzNkVOTIgFe71Wa44wbukFOMsL7dabMT18BGXhy0Jhz829SIv8+wpXI3Z
V+aM1W1HcJDI16o5qtV4dLJ8dhFXdhUlI5jghUk5Rtbn8ZG/sxV3j3rmVHDxwLH1
melwCTtzME/qDntOS9lrzwZwTeV5+VPXZUANR81NJ42j5cO8xiSUetaNfZWgQgCd
dcw6DM2j07G8aAld6P1RvbDqBAs4XGRATgTp2ICpN3qw8pRLW/M158DDptSkhorF
UfYhkWHWgqxZWRjKi0P7LbAYim9TSn2scwB+1zXJAfZhpdN4vU7958PMP6OPLMCU
q2gqe9Tp5ulT05H214qMZwX4owWreOBN0OSuyX0+gDhY0yLWqmHy88sD/VdE/gxn
DiJ8twHgbFwzUfXQ9WDyAjDrQqLZ2LD8VY9S2HE0uZF6vNgTIN4vQfeTiFZaPVqf
T5NG1iy5v2UH+9T6ucaJ1mi0k4Wd2wugcuh+uaorh7gaJ69Dn1cB/HWM320sTIJU
QfwdqmuWjySgsVlEA/1rjEyi7fXD6w/k5utU/Gofj/YNhy0B3yJeV+JDId0m45wt
AMHfDkAC2Gqgd2uZ4Jslp3bNg/4USTS1z9Yb7aw0boDFexz3KozAgntOC7pevZT+
4nqKKw01QhgzG4KPb7bDmKnnYHTBqD5ahek6jQOWs+ZvQ5vBsyiD/VMs5U1IS/+h
2K6tkD2Fyp0h9NJxjKuPGHCCj1qf2SO9cQyQxM8t4xw9/x1YRQJWFWrcKNDaOWzA
3WRwcjNhc8VpU4D1AT/eZ2XJn2IDUsZhiPIofwjqT0CG6hmFr4ff6VomZAEuCcrt
GNIkkH69ZSF0raPLrhoFXQ5zRWQ1Zcz6U3ijTum0sVkhh7cK15kmY0W2dxx0y5U4
cwRtLyZhLKrPBBdbWBZc3asL1cdQSOj+khYtbX0npkIx7s3cjZy3I6CrKrAVG6pK
giP1hqWPPlkINnW/ynZNnzXJPoRebJ34xD9RSlHXu9A+lL9qCikMzPM6sU2v9Nrl
da9l2pTMn2bRtycWmK4RmEmjKKfVHvfhB1psDrX1z4XjAAV/rdX0NuSZ3Qr+2fby
MCMkpk6C4/eRryhETICPG+phBMTZgA45hCTGPQcX/HI36xnXQnbF3HcYPIiaHLJN
JXBBoIv6rRP1LJnXngTnD9PD4CHVJQ2Mli5cq/MCXSNl3Bhg/USmZC21azCI7p7y
cG2PGkRARiE/yrNd49gGJBYd62mAjPxLg3/BzleLYBXkYoBsPCjcq1G8IbswJrjK
bvUoKWH9XSB2WDz3VPDYz0QP6r5YcoUMKAVwmXefIR/D3K3U6PGnDu3056iefwYV
2IWrP4N3GlvMh5dgG30BUxRHg9Vp18HrIERP6DtAnKbwr7eLceaR3kUvIRKAj1z4
+bCjN5FcCFkBZdIiGha1xvV3b1Wb2Ah1mneznehJg8vy1fbR/RzSaGuuA/J56Uxt
RF3ERsf51EbR+fAiqC8qskct1S1q6AlV3xVSsicChA6ZBUYflbw2byUINHylkUc7
FnEHpYPxZ22vfjVUZIpJ8qeicaQNXs+yVwE4fYjePB+8hQYTIVL0+7kOnEfudZA8
Pn3LEN+mj3NQGNpT0/MjFTIQWI3juEO7yyK4bJlOj88wvbS0eLjvhIsNzQ3je8Dc
3FoLPKrMOiKfMguNJUAdbSjeZLK8BUnucUwOqVlCwJVnrEpJEHiqPii6Kt5rUgSV
9K/8byuokslvK5SjtfVafXxe3poxbo6AnKNJpQi0PG18c1y8e1PNMRlDqUbi+Tte
oLW3la3WE02N++P6JLhd4qETWFpNdZ3HFFPMC0qROw+yr+aBC2gq8CR56QdsLMff
hLjwp0YwFEEXZQFsF4tJZJk5y5IEwwvHLvyAPXFdjNOo6GsxZwpoN72s6V56JbQk
KNTqo1efqIiFWnN0D4nUdBkwRL7eL5krm5VfOZ9Ogx+IxHwbaEuImnDjOfkANvUO
W5dtIOzEEa2x9Ny+Hu15rH5/Lglk6/Y9gPas96qscF+J8RvCsCXOBpX73xx3YvZQ
Ss1lrhRUkfnHmTLNn+HcqIZBr0DO5ddSHte9iMHd79ELd25vKTS+iEPUrJp7e3Ms
A4ixLH20hBl5aAnEZdWyt8hNBtIPBEgFuDOFUuJFnGCkgATghP6TJzI1iEQexxWo
MJamUhsAyp1GixGnNKl98hbMuARpy8m6JLzGzlU32MQhoSK2mPwTujfXNTg3gYip
3B3RyP3+KkzJrhyWDSaG9KFDOR/RfykGtUhVBhdBzKxaSeLbaSFcrM1MEEEe/H8e
NxlXuuiPqTT5NDqqOKR4Etx/x1ThNsdagmDxQKFxu5jX2rBoXq/3yr0XnXmTleP9
5FTEndqVI8AqDNIsic2pIZH34Vq5i/moKXRv1bqJ4+rQ/EsTpHKy4eHWJMmIzzfS
bDWaCYP/O+aK0nASHBMHtaO53iRZAg5m+C17raVf1URkAOjEu8qc2wjADsRzhzIm
qL16ANO0T3jRX5b/xBxr8NqrnHQJYhBQ1rSmicfO5uTKFBvebOxV7R3dRd7JmjfH
7sj3TeGlmDhRTzqOVdMUruYO3FEU1F4EcLzlPkWYS6l8tsIckb57JHcfpJLlVzx0
n/9UrYQhkLBT2qGM0Zr6boTvaKgqlKMjH9JU9haoA1iQcdfQMFVwJqweRu4emjSy
21zeSBehZrkW70icUKCPBdZO4mvhpOIp2gm4FNglGpCbo0JV6h2ahQUFqAcmx50f
DvIQBiXTrZcsmmfvVUiYcabUyK+4xgzyIIvBIiHDKd0YoHr4qMHiZy2bfCkbzrvb
q1524v/m3D11P8A05XPQ3gpOFtcfIo7FpW/GJ2ibkzPC1i7NpP3r8zqXM4YZaESv
3VsLtlLWnBuTRoLz3p5Wb1CsPrNyHcjE0sCQ/37SGZsjJrWjS9YHn5q49T2fxAmC
ZkiYF5YvtpyX3gtlJANylkgsHYIhtKXZcIdkpKJc9UNlWc6+/ktWPMCj5lI4SoRZ
H3tDR9DR66reyjomYRPS1RBhp4Shs2DUnyFPoLJ7Q70RRJJMveuzYpVCN08zFw4z
8gOVdenbmZOaCw/4GERJm9ISnhbE7bCh1UoaJVfqDAebuzeAffG8/Gz5Jj+gIr48
kBl6rxHain3NqqLwZnUN8KzdmmPT/WVRtxmZQcky9eYhCfVIlg8xgtIVxlLc030j
Sii6FERLviVE8MZ9PhGcHtEiD65hJ6X/qx/NdhL0xnSAOb5xHXnEew6RTVe6YX8q
nvm3hRubdRcNFD3nfe8mT2cGgKleO5j0Gc8/2AS1szgLV0dzAbmye+zYaG+L7MeV
ITZp1+db2Q/zT5wJNMLiw2CQfXsx8MRA8qza5zI6m7TtMcNbJsEP6enRH2mqsakn
2MGfdj/HkTdrhnzQQgEZNhib33Y2dxepholywtHXwAH2vJUOINZGcdTQIhRKIiK4
cYPLRtFTqKVzIwOKtUiU4jTjsIQEwmJXuCHCFfn7PK+5IGf8DfbQAbi4geSmyqPC
ht0UAZPMifyA4Mo9/42C3kNalEwzaOZO3TUuYD7OVH/QrEL+3f2kI+65jlgdB8OW
Eie/vKfQJzVGI27s5Rdc3APz1ZhhXBC13eE/5OV8agfzYrXc+V8Tg+L6Aue1Nulx
d/7Du5y/hcrcBgUUp1ngpayPchdAJtf7LfZEmL+EXSKXEbvUs0gWDA+pVDxXAyx3
6uLITwgY4+7fjokcmQNmByYREoQb+OwkS7PLJdJj1w6U8zFjvvvZ8Xz6k1/BANNR
/axXAUrjtyGn02JyShkpek644h9XV1d7nb7q19zcN3NdOrb1DI3CtCjGA29LtdhJ
+Oac1RLotJYkD4SNx/t76r3AababQbYduFuETHQq83IsmBZjmjILkpG0Gpkwo4bp
QJkD8JmVLUM02HMzWbziNgZ+DNGgIyTLp27ACFVVqVxzazSj4th3ivB3w8Zq1HNq
JhiXS9NxmSRi06IhzTIPHSKoY+2kTHxY2Rhzb4zbQ8ZUesM68b4Bd4uUizsFbMZB
TUJMFJC8WumHjajpt7OMRgMkcaFRHGy1CgD70FDatmNIETVUoor9KlJhkzqDAe3k
XGpFYyUU4JeoReqYvOTDssmmnCwD4fn/41MqEe5vU1qyvj5iuW8NtbTkmwxCq+Ki
1PxqYugOtNn003soKzZe7GtdGZfJBs+HaeyU4BaJXR88gPIny/xrihHBW62RsB6w
kcoJx2muhCmrLaiy4vMr6UAWb0rfQ50ulP+zA30AZAU1tCe5kfHy/myvG7AMPonf
+seu2DtmajzGZDz3wGPOEyqYeROsIoNNDl3lUfnMe+RZ+lIpOWxpOFtSpQfLfV4D
1GlkQ7KPrvWYnHv7EP835wMLT+83mFKD3KtO2YH4swuoRrpDVAB0o4gjNSgwJW+p
c/hRWB5HyrFsG8fntYW/BTePrXXjfhJ+FCM428ojh1zgIlBXoGl6DwtZ7K+4QOIX
8N8KNJbyvwr5TfF3Kd1gvAxpYCLVWSHdZsSRpgqAWCIjdPeigqO8e3f8FLghAU6P
mLaBLXCc+DUSeeAFo1U9ovhRlwXoZYK0dzO3b/HVj7nKfE0J52tJM+TPGBsA2OCp
Du89rS6SjrxWZm7TthvYJKjoLblj9HUVDdRs4mLif5XA38eO+W0ZlUTlF4AOPYU+
GKB868iqtTLrM3dq0738HzuJEjdXuhjz5PKvMVDBK83gLrPE8vl61Pf54TbiyD75
NEIO4LZAkrVlyza1P3mXy5yBZgigt6gcxjqKi1isEXXpQ14uyK5UZX++j9t0fBi2
tlaTCvWfuEUpkvqQ39s9S14l0IgN2UIlHs3B91EMFxlxrwsD3EpP6Y/lm0++VI2O
sN73EPbR12yp+z0a2DjzNQ/OWYn7BH3SMYDvuiQMCaA9D7/QbYoXdiq12u55j6fO
v0VJYGOBoc1wE+wCJ6M2TcH+YZLNdbPcDVP8Pp+/vDnTBUNijpAPcOeMgqWFCr6R
nVH7wpwRM3mZiheT1rSufK8paW99SRoCwM+y7QK1G5mJTv/S0vAo5xSU9WEffL4t
RkfJyADLGhYR/TVeCoXQzCpa0H0zeeoY8PIacu5iKxyyBrkPrhb70DXmDNZn4lRt
0WM/HlXnRUO5hQpwobj3DurbYYsb+DdGcwS18C3HHz4SrZXv+X9Y4cDzLXa0p71W
OlfGeJ4iuQn4UPHttxpqNSZ/jhHExtLhUF57aEzW5StolkdbfkPDAPZCa8aM+qe/
USxMbVwvUbkvAKNgffKAx/llPlI/sLB9ujjUIndfN9uBdx2D/Hf9FRQ8Z1h0AVkp
FOF11rykGnloYTXS0AScF0uRNzj1aMOSjJ6epK6l/C9LapU4a0lVavq047dD0a/O
NG4xeJMcqU5H+xhFeSmI657oLs4cBGEECIBrdqqB3D8Rnu1UmHte0SdX1vv/4SXw
gpNUDiFPBSYiO6cASwGXd4u8IPNmHwaEdFESkN6smMYI+xYxWsnAnlF6PK2TGgaT
RJZMWZfb+ISttIYrOIHJhlkAxSX+V9CZE90oIQ98HORLRiGBgNpA2agm4mZBo68W
SR0i/TuSmLfgtb9W5OOKNFnQBldvfjo6uicr4VU4ymglaV59zR6+1mUrPHsmESLB
yjc7psZAJl2d6En8f6l7BzpHNUq7WGk3R7MS5cwyLRYY2RBF94uihjlU12vRaKCC
r/ICTZ5Pv9dFmPeRAmsg4oSmHWsq8lz5OE51HyhBJDeYifs6Zt0WKmOtqV5qMnC3
Kbym5zjjeWheBtrj1l1hAz+oQNLR14EW+B7QX+KOqB+XsUHKCM1+eky5ezuql9D8
z5C1RVDEfj51tu2wX1H9kCp81UiBnc5OF3YkQL82GaXCXyO+Vq8C9oagZm7UQxaX
0B+5GpEHWHvHVpOeAiDQ0qjeBabclKcvmlFumLubGK737tixCk/JFPii0ldUldkl
2NyukwbKDFY7jFzATsg3Ty/gV5nUqmmDXb487LXS27kYYpAB+98EaqUjcUEMIQ5R
IcBs858kcrUvVSATGCRRvye3TmtxjWHNX7hzJvDgkkiH8ADfwCL/TrvCZTbw0b7Q
rcEkH2wTZgJBX2zx60WvjTw9HV4cVcp7Am42PyTXrVQ80qMjPSdRHrUds3faMsXX
vjPYALaxkCI5+dC6Kf2DEmWBj6VlOyPnEBkEcX0FfzBw2SvadbMgkVxk1DrpzmrO
3egnoEoMrKQ+435moqBi/1KrRqtBOzO83RfNh367qZXyg83tsPm0afo87Xs6QuoN
AKb2PcdQ6kNHLeYunx6penK/8AaXVc9SRtKS9wVNCKMyKNtuhwRm8JRbefO3zKeI
d1LtfdoCHlGVUVEITbw+yCdo4T5ngCuUuhGXoksYbm5+FaRxLFY+bZOikuOX8tVK
FBuWw93OZeD0R4FKqWnpwgZHhKzvFWWUYEJJKisxRAq8da3XSiF8zpJtO0bdVEZZ
zoh9xQaQ5IK+4YKzHo4oPTspb35GOyJkeKRugZqwoWp5yKgK3htoISa/76kiQZ2x
1I0+Hji+sMGiukbOgjV69GlkXdj1RsvkBay37nQZSb64r7RI0mkpuGS6q3rPWwfv
eEba+7LKo511q69EZnMbWalwQZeAAnhva7avdXECpuV8sPC7rqvQ7Cfaa7+klphg
ZFyK2LMwHTEzv6Mej1gG2Abs7EJ5m6J/CgEdORDoksLqsRiTj72aJK38iujgTbbg
AQLkpJy/zm0Tl5bV7pN5r0k3ukmudyuOVcX1nLwTassiena05x6aX8GrYDUVD6Vq
GXIJHnm1dNmnKuNtPmyA1qMT3PR7bVKggueW4J1x7b9Oi/L9TmCZ9aCvQlIn7NdQ
mjVGdTIQN7ifhTxKqS1OvlOWqkEPhSDxtcCOnL5p0XR0mpMihWXT8ZrPhTzvbhIL
eDrfeNVnyN+bm+9vsB+epKAeJKhHrhIhZhcR+AB5YoG+41WlDTrpxJTZ/94IMlWT
jJxrAieagx0jWLIHxzhh2YPQk9efgpU2VzKYoHskLi/Oeo8WeT3jr/r7X4lmD489
ahLi8DRTHmDW9KkqF780UotO9hQ9NkZFnUGIudpKQypho+WErSLATn9o3OTpEIOl
zblPI4/cbvpdbsakyELTq7BHlQRJ2aMUF4fZGLrgp/ojZNOy3iyFuNsQAc39WX/R
34dwAe3BfrTfgMFzz9U/bNTZGavg8FtKSPMyFPB1Si4PUaZRv5kVjfOjyLdl8OaT
23JT6dXx2yLFp+v/fNXdzwB6vGZ9x2geyaT37ZLQOx7rf+bIe3fz1d8x5kp8iV+b
bBJJXGBDw1DrngRdL1YG81DQqW1Qod5TeNPhl4LLpdLcPvriUMj1RJ8RsQNUOWDl
GGsAZwpxFTIQuEba1X9/83EsaHfFr7CaV//Ims6wUmOkuFtsUBat8zWJbXQ/fHJI
TBeP9BT+l1ULLy0M3Fsfcf89B+5/y5qCZdbeZoh4yyr6OfU3NGwJrcAlmBlKfQpP
CkeKpc0p2CcA6ojJkSULyHjRBYe/3rcwaqLlyUuf8iIqooqWy60dVCIIcU84TRmM
dYUy27shsQXr5XRYeT7JPdBMg+BTTAKou1SofWLLgC0Wp7UKsK4HG3BnbYLBZlhq
NMm3us/vTh8d0sB4R4Fj9j1FqFkVisPZ7B9ZR+IcFe12t1VL3EKSTfgdXLT+LPjQ
2iKCo945RlWz9/mKTGz+Jejbk2vbsaEa8x3y9pD6gA4cofDIQW14lI5wyEnC1jI6
uH+nKWie3Qq4BjLpd4Rk+bQR1/uJPP7xAYRFvkG0f1TeILBPtPLhZTSWdVHMXCql
526X09kues6fwKz8rpSD6sUojrAOcg7cnRhx90JUpjCD7462eDNCpUHwaVqqsh2j
1yohOXxDKkpLHIcWqPs9UG4jITL5+POI7yClkyA7xh7h7kSUFWztRxkfc1HqNwcT
GH6wUXPEi+ceNfVh67TmWphlsiWo6iSFAzrjb5CLha2C/2REqJB4U1pLfp3BFcvv
7GJ6zmnlca8Z6XzsLAu6IHEWCrH9BACQi75+v37QbdcmlBuZrlSu2J9vTnyPZFs9
ICKF0J2ujCUJLvRXloNmhx7w8AZA9XvSUCc5jAFeUedhBtkX9wOCS3xCdwvse9/J
oWHHgjHmnIjEbBA8lAdgpNQGmp/uH41dLs5isA4TWrK8nWDgcB+eDuLabjydzbPV
3B4JeN5DDmAJUFWF07X3VwnGNwbJTUORNHiKtQhJQh4UU0uF9DtlP3Y3wQMr7Yh6
iuQgZiiVjTZiImB6TcOhXx1DcJZIhCmT/FFoNEM3wMlQ1Bd0h/Kz7mWWzTAiR3hl
drwBK8ik3zxATr0a+j6IlPGJMKBWFV3mpzQblLyDkzrLJgC1Ul5Vv6VBU3931fCL
625jzcfksjuo9Vw7DREuGCIe62CLOQ3mQzm7CzZdsu9Ez7V1I2qenzzPRIfqcGTh
I9V/5Bq0FVgvu9J/k7Iog3TC42pio/scsqkLnCTx7UQoKTrfkpMn2B+4b3FXuj1Z
NgDTGeAAXHwriaap3H/ZxqWcrWZuA++7YkyYTxVR4dEm8j10D0rlFj3G6VM4+kVJ
CfCSk1ZLFL79YpSz8NNi0QERsBgIXFMIeWOZhzdX5W9gf4fJHUhM8p7OV92UySmu
bG3eQuJ/sIW+/n9u6XxyXEOTVYqvQ2iQH771ec1uPeALhjPjMc3wYyjM1cpDZOr6
fkIKnLLxT1qSgipUvOJKijQ08esWEwc2qnhY/fp0PsQyDEv23TJ3PE0nPTzHwBqd
yGJpaEt35CRJHn0KMg9wEUpmzkQkd2H+guVYhraLIjPxUDThyZkSeAEYQfflHs0m
P3bNqBSLUUjPuUhM4kCDWYHcIIK9YBvgl2Amt8PB0eZWeKFgHMLEJjF8BtKOm77o
NXzxmY8YtwS8+I0UGZFLbjjPs/2pAfKYjGFJ+3wSJyENNytauCTRUr0tajtD9UOz
3/czTfNhGl4mrUyHA4UhX+cxiyyl2OpZI6uzGyGWSNjacWGkKOODcVLt0SJQMAZ8
GMgIZ1G0kIavrEDU0eMh/h95cwgqdam7nAHWBOSGJBcLm1wZL4c5dXqL6uXUWJcI
IcvzsGqMSPD+bHxY9B6HthPwy7ayoDQcyMl0JE60AgKikPaFbKzcs3+uhcufJNR+
t+SlJN2aIKMo6aD/bkDxd0ourYernlxd3fe5DPOHVOJT4e8rc70TWNX6LeohqfS0
2a0fcndrLSIeQTfn68+hhFPiSHLxhkqZ0hfW3d4gHOb4ymdDRZtRFvF9354zlg47
W15YBTQchq6m8oO20kk4tW9qB45elF+6AUBvKusX1bYhjdflNRCzhvXy39n2z7AW
YyaBgqJYp04XDJZsuvo0Tw7AmfaS+v3nWAytODwgtK/wj0jqzxDSKGAWME6P63Fw
BiaNVm3EawWx+RPs/YTq16blk2j2BNHz31hpfsXRXp2WKKisz5c5P+1nqrs65F1b
WGa7TsSp+dfY9vcHNO3s2wgrUByol3Gw1YcB8d3nXugfECPaO5UsaX+Bd1E6/ib6
Pqa5oVmbyqxj79BVAAeTHTU3LzVAhFep0jlmUoXp2YfwKOVYUh3ryJQa1P9osyeg
zcy+5m3aO3Ztbo3HkqRS0bf2KVHZ4u66QpNGuSbxnbgmsqM700OAxMS1+8GZZxCp
ALCSPQ8U+z9Adt8z6RYygDggiYjJoPQRDpRZQ3hXEHVyvOk017I6IEgF1PyJgRCm
5HY5PEANWj2GXQ6dqnPXK29i1vnBBewRoGccVzuz1rL4Rbg6hxaGY95YfkyZe5NA
dpKqmdx8hBLyJvWILG1i1KFxAwTzCHldGaogkvT+dRkCPDgfOpRPcFv+bqLworyL
cVPZ5reA+Yow0o8YiRZrqzh0kjehfbolBTT5Jn438p9/GpK5V6C4FIDm1mIyNqfS
7hEYCcbZuhdXQgIccwy0B4E7l1LhNHJZUPGcdij6ZM+anXC1MGmFsGGrOnKDUM/6
+ax+qDDgOcSol767bILSJZQz+ilufQyBvH+eW5QbLpJJLDBn0kLJY2209y3UYwpQ
X9fM6W5o5cKZ4XWG+MwmQ35SUh/PuTPV1bAsdbrd/rTHaWWGpQMGipf4BmdDQEJ1
sBJxrgBsKhtHaGJXFBMx3Y5KwM3QbzrPNZjK9RGK7wL0IPQgOm1XGDseFrLnD4Eh
w00S2mYsu3lEXiuuHdcDcm6a+S+4qtFfonGpRy/LN29OeKeKoymiyFjnYHbBdTf9
/lDASwm6XKboV5LvI+z1Q5ynNaU5AOyveX6VVyuMXZMgICDBKzpHndeKMm2imjJW
8kkGjtqJ2JJRFALGN9M680Ds2TKrrBi08S1yCkb+foLDHB+JJA9QI2yCqcfxkJfG
Eyxwz7TtjiD3Q5ZoRI4/zq1H/BNWBwpN43awIAiE+GwxlZLfYBC7yEkYssByUMqr
DXfudikHjB/w+GJM6rg5MpvGTajZHK09pdrjw7TRW26JfL9FdbsMF5qWhhxOfz5N
8Gz4u4gD6uZa71iyZwQvxYMnqEgqh7oiTKysYRphEMLaR0WGvP0otdowxOvuyu3b
glNre3aoja+omoOIr4/tb3PWRPtmnbnlChmTtEk4PnzNUd/rsC6fmWn3brBLFXh4
qceFH8AdfH7oI9MKM1bNyufqWkop8MqDrqCgdVq4l5/VlHQIEYO9alYsDfWMeQJG
O0Oo/xDLkwLxpzTdN9xMyNaV180pEexQ9nz3hoo4gccLqh1xhsOUpEHT6ki6itrV
dU8UAIo9j64SBQb7q6+V6bejlE02DxHTVgGCURw+wrWAUGrA1xKWugAqtUkRRKsb
t9mvCGVJiZfwIjCr+ORPUKBI82eU/YfgB/rPJD3eKPyTHRScuYxHlJcMAo6DEF/b
sBKTE0viDroqOZL1NM7MAVx4mt9bcyOXATbyDownq7YDPWX55t7WEY5pCEBS21sF
ZWgGW6m896KWvekwsMxv31O7hyfvKwLkzWsQELRY0hfPkA/xu7CnLfsREpy3fO8G
oFV7QR/jnyUzoUj5i7gquiMRWR89XpLRz6sT6VvrYEvANHsbU9fY+p7qCgVhx0H/
6CusqpNH5iQNUOCe3SWzsyysWI93lTnEJowPdOtHSewGK2AcIGlIoxaJN7lkC0a7
hebI06lpfnt+F++oFydV0f2UETXTCd4cxZYmR2MjQiVBzQ2fg/n8bZOPWnhBYkDc
cNxfwXg5xF2QI+oDJ8DN4bf5BQWY1VWThrEGuaqpXboiWa3totjP++QTtHW1bgk3
iCDj+NCmsLrpHqo7TkufRAFbIDh926SsxH2nuydtzhyK7gqBQGxTknHo9lcTKSnW
WhVI33ja9JlrBEMZra0Y13EgjQq09dN1uLqmlXJ/NcKfoq6758MQF2CEXudtfufs
0lI48fKYNN7zeS4mss9riLX7XV/xSZ+muCkcIt88hME/G5ZmzG8dOW4sTrLeoYmR
n9Xbq/FAwgW1zdiiQjHhZrHWG16NmvRv09lzO6LFDbp+ugxp1cjTyL/ABLjJMkOU
aIt1i/1cPDok4puVMCjVMoganj81qO2VcHY75r1FAiz98GZ3D1w0Mug79YI/y8XL
LksPAQr69Vkw5q11jUUURIELdwx2TZhfOwlk7J7glbnP7taWlFpg0Tw6CK8YbqCv
rXMIKciM/KTEdQMVrGAbmQs1EG7kSnS3Vqav6ksFOsdLiU8sxhDCg6S55mQuYXIS
vptwu6Zwvu4Z2iKd8JoRMeciIn17kp+JVPiRZwDG/Ii56FjDY205hsDQcs+CrUvG
r2pN0xxE28awoB/BK0++rJn3x8NNbs0MbAlFMJ9N2ex3Omol1NUDgo1IwaDr+YCI
i0oXFepJ5NfbgU2U9gGOXkK+pZv3+ta/meqkprvT5D5HPouvFGx0T8nNlbnzAMkl
46DxQ4Q/Z2MziLij1nXozggy4KQhOBvkeWEd5dFCQ6057LGEAXGqU1XM/+y1FNLA
/NYonBYf9WdjHLozjr31ssln2KBhqlj2i8winRJlbBl/thxA8O6puqeV6f6AMXeN
2Vn7qWGq+JhkMszf7CDGv4W1HVFyqlm8J9mE1PBgfmZmYyU12pGnX/U5dYt/b0lY
DYns8vinMlk5w9pdwQwJXSOqsK86BDCMt+VqRcV13y5AXXVcmUO8gG+7jF275dx9
jrNz1v/qzDcDZx2CEs139aftHx8kwgXIwPOfEXRfx4g/oE5XgBkHmXZ62LPnN6j1
juaL29JF79NLsO0SNseca12thYH3hIuckQFHyaY1EU4U9eERSpiAftochndhEbDu
sRkhreTmxObE/V7z2nWprjRDIEKo0j3YC7wq86cDnVjQYUCeyNvBNR0gFutPcCcZ
YowGETdQ9KNsiEbjV7uKVIUDiRq9sbsYZmF4RCnuWMNgWcQ2Z2wgx8cXBkrGTlVP
jtZk1a089lomp8mMVBMBZluOsNnJVDace2ysGb3QNylDyabwDMaXnmSmP3T5TToG
APFOGDBPYYmXWinlWnoUFBgYgQLECI5N7SvZoqbK/ULgU9/2p7FmEdZvYGiVvlKx
TTBSv04S9nwjAjWkXOoYfDOxaoJRq7hGlr++AF+mxoLW+u/+MDxLOAoHqklPESWM
lMyJBFyo3ZrfISIeciKYhtDz5RZZwgw5P5qbXW2nc9I0TH0jKsHunWktYzp4Lf1C
8YnPVLkL7tAy04hCLVQiq4q1OD2/AuuvvLHm9gFGhEJ7Kd4+vbJ42EvCKIsgBHbk
F01BE1MxHPbG+MRZprNmOLXcSM1GpQPXXPMA0n6mDuzNEBW7vJFSHA9ZGU9WW5Mt
JYT+Mv5kV67hsXZHbAk14qe+SWck5dEHGmYisoleoReTU0laEeoQc0PMEvlTVMv7
dsye3ce0IHbdUfvUdiAaQuEhtYBgcAwB8YgRZDLw4SwSRR0qJbRadnJ6ZkRK4A8Y
P1kxmRw+WQakPIHfddPVadxjcQE8TMd1pjoq56Gk/STpJ6qwO5OO6JKHvQ9Lej7C
sfWfGRVz63KyInS3juyAvkDQ+3u5N+whp2+XKqB58vSejl4BN5czINLLFk/MX3zV
0Q39G5mZgrTDzRVgxSxx2CHIJ1eSU5kbiu3pZPxWB4Y499WOZVJ/EfT34FKIIoc5
sXXyfF3JDuz7iNBIbIoAfopq0p/wTcLvTDgF0Qjv2lFrPvhSbuh1lkw0qT08w1Hr
B8X0F18zciu6Rwni96ljziuEPzUzLeGxK3xAU4/vm70b5Ie0cpGzaxsMOHvjeGYL
wpsWmXzT0deeaaWxMJelew0gcJOYzySTwE9RdjtunLMDEDmP/C4XUW0tBmdOtFq6
jzipByjXAEfj0cTNkr3BcXB0rSOItM3OAQiNaY1FWX7lryhAmze9BQ3f5409/FXG
LWxVmpV/CL475wIUzZRdHjcYAuSLPwnej4bm185rxMEp09nEvFKudqraEadb80Qb
NsRx9K0RUOahGdkKE03HF0qiTUzlXUwpr+XACoqXVe/b90VrtEIdkyoZSibV3Wi7
MBOkUYDz/tTAEYlWmbHJN4VZ3UXp7bdB8MEe4kBpAbOyIFUNzja2rYEu3Y68bYID
pXgwsc1DnDLpg9gEnA4KzcIM+6FcyF/KFe16WdwqD/Vl5mYnoITFWAjfmYzf00PI
n25HMGccpHDagsKEg1vqzm2Yfux3LvTFvdkj5p/tGSeH32Ndt7quheKwgD0ZWmm/
rLji8XI03okGAbS8z3MvuZwKLuUCuE3dZ8RLRWrxQ39dqBBaBbyE2kG3M9+O4aj8
jtWHBoar6PGfjzmYW0porVlg9zJZkvYPpV1+kvOfjsYyL7Fjbi47lXgKQgxcNzbo
77uFhWUt3XD4wCeeObTzLvRbLh70lwTtANYWpqmOG4f+pXn7jyd1o6ieXotgzMRi
TNYbmOMUXcw3AZoBLMgrylFOTQ+CD3huGnGj0PYtYlAorRnSM+guzvFgNDqNK2LJ
ayotF0E5euxx2fqBcCX+/u5N6CrOhtlHjZxx1stJ4K6xh5y6TLtkFm+T003kJKhi
0gKRf0bfpz0ZtsGqSvNFYauGNitq8ZKdHVd/sx9qR5TWE3Pw1ocwh6jvFn1VzuRc
BbupZqwUqZMFjkZ55/qtiF1DeHBSDZTq0fmQ3ZrZ0SCpTN8+LbBIcSPnE+yu+k40
Z3pV4W/y5nRHNEuW51E6PpmtORg/BOl/NV7NAj8y0HnXFnsZcqhkvUK3dMEKNNOJ
P/u24B8mBLlwdYdpmMK21nLdSM41C5nkL4WnHr/mqaz+/Gj4BRcyNI0o9GUm2kdb
9TYyCXVDCLDsMW74bEPvzVvtrL3+M1EZOEhBS7cBMkaNFnPLzyGzGJHsejKCE/EL
kMKx6Gg/POn6Jz8OAUUkxgpyn3nwSX2U1abkXFXka0cfH8KZIWUwwe/8VjBs+JS4
b7qswcgOQgAAzY/7MYpARPdJwIyjbgcoTZbbeUb3aPfFb/8ZoazZIJO5KiyN1B5e
RVakRrBij5hIPDxRsNaGQnuT7Sw98VGMKif0MpRq2AKeftT2SuxWnFbkbSKD0PKp
aF+kNxCvjXG2xScZeTTLs/9mIi87D+nhXp60E1Ivu1I2K9qWjkuAm/Ie7lHZcAdC
ezROkZe0DxLbbrdxiQIoYu18fgL30MITscLPIyUhFeooXuCW1vdezpvlxEmdN2EU
f9AcC8rlDv9ex7YYoi1pN8Jw7QglUdoMWEaGzlFE46/pOK4+DjKFefxUfNzTxlyT
rO7+Nej9i41ty3WA128NQO9xg/2/+K8m0SmFS8nmMFDWJ/a5kxhGFaZUfbPGnQA0
nmIj89J6NWAF10gwHVL1+16z2OwQpvmoH9aKowG+TFx7SVhh2KchKpEpkiylT+wE
DVVlGDV1HWl6/PUiL4aW6WtzGbKeaf6Mn91fVf4H+rTXBvQ5OZxCkKFMAGEhgwSO
/E/t4VLWIZjHAVhkcoJgG6rNNlHK/aobNMM8twRWF0wyT+fQ+TZ/sjSoV0o7V/e2
NrmPmNFGUhK52nHuWs5O7JHbOa2wUhY/nISNPviwWP3R/fozjfk9YvExOJcj3YSt
XfrrOWxW3B2Sg36cyfuwnQzJ1MP/pE6bV97nmh9WBjQiS/eumYS/ZpgoCeCHDkZo
Iv6Hr0jOJ9/Txo2sx/GMQnict/1hpNwCUYs4QkCFFgi15oF4ncZoupddp4HpJu/h
d5LyiWsHi/9QEG+X6mLD81xR09zl+oW5kNhYW40Vbg3kMrF9VlCPNacBdgVYNAIv
jjhDA0g0pZP+/EiAK18t54jinh6JHZVITM3Xk+WmVaW0c2IzwHBtnP0Wxtw1fLEV
Ue6kjI2sRuXPw0f29yMPtbbzY6AVmwvx+KqyuM/kOrMRRR+8uaxGOpYmnBW1gLsP
Jyd2/Sa5I0cbb97A+/JVARMC2h9RHVuhzTUBBcumaJDJ82+IzOv7QwX8e3ws4HXq
whlL4+S0t+0K/jUwnzrB4iquGkNXZt/dAEJ9oXUTffb0kQ4hZvwQNtV+6nAtVRkm
hcnLy6BeBypVR3JxNskDPhpgtz2+DAQEYTr41ZiNzYBKVQoTLGotHKAsY8VWacd/
NxUMWtDIwH8Z2+xrD4u/sZaJoMnM+Ds9UluJfBQ58Un3+7fBmVFOQu4uf3sh+1hj
zA6VBoNWuZd7fzzHPawonWE7+k1MKq/ZKR1K2GyJQpZztzLDiUcXLpubO/zo3JYC
J1xhtrY0PkNSce96pG/FHxf6irzaXPE7mMR5169CJKWX8RJVcfKcC6pftUNqpofO
b/bGFt+0b18B9/ecEz0238qXZjNnL6sNg9NwEPX+254W7ipTXNK/sBhnaScuoq1N
HjHUHSFH8gnnlRxeHEd0ny9a1PD+Bk/fC/5XIZXU9BQn4XINUqsKxqQdmW+MaECq
l1snhO2Nv8yl9QMj19ZDA6TV6YOpPjkbggd5eOH8Ty8MZeWn6h0aZdRnjbzXXhzD
ip9MC7fUG8nkHLh6ayihGIxBc08WKQjzAqUXqrrHyU5pfxlL2ckSXzNwytuLuHQS
SqBwtfrf95ZcPXe2pGL8nr5nRIDUGVLqDIREoAksbwS7v6MApiWoemyN1GPWFmbC
EEs0+eoUW92VDZB7S+lT2yiSiXbK/Lymb3koNvn6IYncYvkgzm1jmC+UFOpdb00w
hQF1/QugS7Tgi0R9eiEmbUkBqZ1Ov6MhP3Bs6HF5uhB1eHaVWOBLGPCTnyNnwHYd
pHO2rqyxdrt3niift4okknXGt1VcnqfdHmNR7aowebTh0UIK0heazZT6JhC8JJqd
v62Y/Mi6n0Sx2U5t9Szn5JMfCJ8NQc/aeBTjLA+euwNAD83OQ0Gpcw0OsuiZcJ+e
3lVaDoPeV0wkkWzLEWTP9yIbh1s69utrtC7CRtqfuKHAfDnBORw2tQz4MTYRwTVS
K8AG7Fvtpp1spBGhjb3xZ5h6xbMunbU7p9OM2EyqSiRpY5Hv6niuDhBmat1qy1qr
a57NS3K6BsgH1osXOx/qH2SOopGH6hm6BIcdzBtYAdrGYhKdKdL5XFpGyQKq4kPE
nzgo0cPrxMfznepPYkWa2tQFUclmLYfhw2652gZKyjvxYeqlWesgH5XQEp6jmM/x
1GQBog5dbnJgvoo3gXUmZ71HSaYH+m0cM2EkgYeBO8YH1F64wAovnpMaZLinanoZ
7RJc50nHFV5e1zyMLBofkF4OaD7FuEjIabxB4bhFf48fu6GpQrE2xGycuemtQRfE
2HzpA4DLTec5KAv4Hr5QTYNDsuHbIIuiVp3wVyoc5+bsLKFAw8Hw3d1e9rdxHwRw
1VX0f9GbTnBu1pozrwhanEgvAbPPbjLCTSR44kbwNFkpyMtr5isdLOwtnAwNuHGX
EeTnV/rI36Tr+MSTmskCy6wgs/OPxXjYmwQGKEhpcPkvEL/DSbox/n4JOAJZE+wZ
7jKRG7vLnLep/hDmwGtZ84F4uhodCFcBq0ZNLm0/DAHsvghlyXGPJWmKhXHL0ra9
OWSQDbcmXW/oDP8aK8iC6sSP4xC34dXF5aCUrIFvb59mMOIXTYbgbhkx/eu/DdhL
Llvo9QrAHPyoVZH0WR98tw0DUVDohpyFAQwHZKozpPhHViEDsAskWYAyVFgXBOGd
q3em08Ou6ok2qbEc/31lJXmu9WyV1OuaWpnOjpzerirckc6Z+qr8mPStWgaTW2pT
1VWqCPp25SHVQOVmVb++ZQ0gLJpwEhLEiqCm75Q0VRRvqQe6XE988i+Ns3CZgeoc
5wnXM9fCpznmvlPxIDwT/FMADhXdRGFgdI5uxNTYEUsi1VZ6VFgpgi8vgbnFjaSG
ausUh50syZvYwBJA+mtwEZ08vZf0WyXfEQELKZyviaUz8xbv4zlbWLg2q1J7jhl2
JMNzYFmpcr10lsUlvXHZ8Tp301L9DMTZFtKpKJFgtcoJ8vbiBQUmCNLkZ693L73I
FAl2Ax3IlRSmIynjPyIvDcB5zCZOQQHgXf7VvZQ7yyOwUWDUjeAjZ8uJ2hSI7p3z
hbhp+BgEkpQ2NkJIt/YLSJY3ktwEEyWf5DOl2AaK4Cy9/RlTic87qDeUdq1IWVvH
XKIK3ZNoWkGnwnUdVO/ABg2R9UNERTPHNJbb7I5pKaFcM7sVJVkXEuDYp4C3jYO2
bO2moqFxc7TPcQy0R1JCp0Z+cCdP+UVmytq+S2eE9Pd3kGfQ0y5xhfS0rexN9Kst
F0iyDr+Lu/agRdzGeIa/U8cRXEWLxORurkMj5E3RIyeFo82NYzNsVN0lGp5R1sxq
tCf9915nInu4d3aH8VnQS/UH9+w+GkNFPcS3YsaPZ+igPY1slwLBJOy3vaKV0bfB
PecOJButk9jt8VI7eRUR1ApSqX6oaGCe0mU7McCDV7+q99DiwYlLSQ3jKwLsIy5P
mmJgfH5rnC9TZXHTPlkuZwFRd4d6PQ9Fsm925eR22H5k/yMJJA0UvDBkYLAggpqN
tBVoEq/7EQTgtDylEbmSMSFiDqh/i67so6IGbp1Ojm/Bhjp8iTJ8SBeAPXlJ9Daf
EU4LIdvhJwn+KAxUjCJwqdPb+jDoNXDJWaVSXqk7Ir23NUf0wA5OTL0Og5qgGtTt
XsTyuRHB2B0lxDK4kTa9MvSDBda/k3Ke7YnuFvez/kGURXet4BshXvmL5dO9TEQf
avacQK0p/4gPIegP/raJoJMBZjGJPYTeXuWCs1qspBJwAyRVb8cpODtFgRmNiXUP
Ye8MD529k1Jt5mwTvLXPWhXKisgqe9GbQpW4JF5HkKOmlNX9eNOAHtgKuRycEeJn
1siz77rDoW/FerJOpiWBu7Y9Utm7xokATjg3gf2wUraIL+yFq/JCqo5MERDI2Ov6
Sg+yLX1hRINHcQljXU+0XEPRiSP+dE5xMnz1x6BbO/6ibjmqz6h/gCNo/yaSq84O
YUyzgp2654yrc62WzbVLVEiccpftJHBT/WfcTvTItEyQ3/ML7trPxkLjHrHpjjcw
hsUF4Q/ExHFDlxqipZVIdOZiv9dQ8UhagCIKvz1/YzfHOeIUO+Rax7QP7jVhB6B3
R/IkYFDtFwdxVbpi4rdkgPPNC17rOq9189iyw5gHTVQXghRLwUeKhm7HBXUv3Br8
uPH037ifB7fLDn0h3LqoaX/qAtdDnIvRN1w0t0D9v8Hy/XHFLCjxedLsDafnMIh6
6NudcJD69OXAcYxW9DKtMyHbkHJQn7RNEgHI4fR/yZVKrX/U0/7CQ1MeE9y6sazX
JT7Zx5GUY4BeoVBncUV1AY2h48x+hcvJHgyCzDouZqol/W1dptZOirdHn1SGP/5t
6+Xo7F7e5Azl0OtPGacq50UV7HXKB1c5T5ePBSFd1oG8P3SmiJlUTWUi9fryvi28
CIV/rcUYZwPmY+A6JU02rpAZlHq70U3IKfTjCcvh6FQYG5H0xHBfvQ+9dGXLXPfT
vE7fYRuWzIYzeK5H7MQR5Em7tWg0jKKvnTHsvy7OJ3UXlH8ZYF18/FsL8cjIm6FJ
5NmRHomYWxCGu9hqXHuS/V2RV17PtMKWCDOprhNuY1fHXG26+0GHOhXlubfDR87X
mke5p5MUTFivpoYv6ktScDZhLx9/fYSmsgPuhFagzmeqbtdnkxCAZIz89UWkkyuo
8pEFxqsmEStzRkkugY7ICM9B+tcTdX39NV8s/cBgZSv4ukQbyjCTaF7bc/UGzh2v
iGJxR8MsknXznrZSSGXe2nHKBh5opTDGzgDq0idSeRsFAsiQUwBDBrJ2HiLHheDT
wOIdFptRuEYljqVowakOxsMMQT0Vooltj/KkGfYWvdoBJKH8NA2x19A6Wfx0O3c/
RmqAqE5zD9HTCbpb1C3MxvF+JsiF9lMqHNh1uvXFsQ2dCwhgwfCRuxNFMOhi48N3
Xh6Ixc8LpPtAsAKAApDum9L2p1NxRxNQYTo7+BMyUEKhTplozGRn9X/pvnzMQmE9
B+faGFUFaGBDb318wl/sLN/IcUg4ksbz2c40lqDXj98H3byqqLyKY011RVp74hjI
x3jkOzPPq1XkYVlrYx32tYdWbgmTUnOXaqEK87hhShrl+Cpymhweh/5U0LGD5XRU
QJ9dKDRNnBfWoU0K3snGrSSEmWcIxQHcDZR6e/yALq+1bUqOBXkya4sOeyEN+D1U
XZEunuT0prgziOTsfrRJCVwzs6N8HV1ePQIwUYIkGQIg/ltVNlq0HyCb03vvUb6k
Pl9cPiO0xrApwCnxUeIQ5myOdZRIsy8sOsEgkdLa39PDb2jj1A5lCGJPPFZk2OvG
sgt9GpcOr44OvVrvJH0MnWI6SzOVujc5hNBVOnA3YPJpWL/vKLcfLR25t1S2iQ3f
eiiwBWbds/t10yPGKI8gHV8rsIK4knbfYsEcIObMP58X04J2WgWQF6kGuT+dmolf
ygzx0aijeKXQclkxXCRGWKaC4TbCXJlYI1OR7fZmybuRUQTUrVyvic19un0obPM7
hgt4V3JcZyIjannpr82DQ4Qs6J9LZwlLCIlD7NyLsYia5gZAfmr1e3pCzWoUz//G
5p8utc5ydqfwBa9LJNkbzC0px9WB5SGqZevmjoAG+ry4wIerHTNUJ2F21jj5aHHm
PPFQ2oMz6y5dKfnY9p6C0xvKnME360mvXZby+D8I5KKWAea5xKDAI4z09tfqZNzh
uonOCOd/mrYGuwd3aZYzfAcc+uMJmrP3tZLDd739y1663yzcpdSMrKCmoUL0yAiC
NmoQ4WkNZBLxYl9w2XFYn/CK+BkZqtUc6UMc9/5v3rM1qbf95WH1pX3idoGaypEZ
WvNiCvQE82vwkuiSjfWlPakEOcKeAZ1m27GIPGiHKPuc9CtP5WBI3l0XZEP9Tf1y
Gk1BFID8A2xS57uAL6+t7MdsOE0CFM2/AJ1GBR8e+1KHivtR7pj3/AVnAGV2CtlU
S9wAjfnycxSzcYCDTDD4jZrhOM+LkG6LiM6a15roYIwCncos94JZnIhkOAEPdO9v
xJXOC7Z1lIlNldl3VQC7thPycQcHHA12DtSVXee67yO5vSImrSWwYTbPBUeFKlBW
frV0mOExIbV9//eQAVHiN2WmSiV+aofvCRMih+h02PJrIdpF+wd1CpOe0OLhSVfn
bwxYPF6i5GSftFMcJI18Q4i0UQny2LWbjXpM8fg2WamfIiT40ytpkSrIHMHuG/3R
CqNb65afSmtSXAK4UeX5XUD/xMkGBCBw6EBbPaCdVYRTo+RAS1xYky7OWo9idv7T
vLT3715cdIvjBAGKXivJkchx11VZz1tm6QXe2rji7RDq951Q1mNthu4gHh7iwWE6
mvVhEF2LY/Jvw8VWHFHdpU5OdfX2MyAtsCgFnTbUNhzrRKv3aRWOTlxeICXMHJFN
6VgMKWRBRNJ0o817b8o4q+E+SVqm2+EVxcG60nzGfKDr6N014sUHCEZJC8k6mp18
b6Wi32XaXjx0rIbFjuk5h+pjbI1ba/+cnQ65+p/MiVjb0D8RYHWE8WxzAvYR0YLj
Ck0QurPKuIj3rBo59yTuTjW7Xl1iam5GGra1NTxyGewkQyGwFJp1CakRMaXoNzF6
m5knO2m480WAQDGRAFNVfdyRPgoRffP85vLd8TG3MLqCTrvHhN/O5Ghun6Oc5YDI
owpiJOg4feo5YAthBc6lCP1mey6RhEDAbNWNpXPD8XINrh6HZNYO0SGUPuIfiTbO
g44i/JD2CBjPzbPVGv8in5c8yH8xfjKT8Ya+8SX8iy3WZKqWmpY/C1SKVcjiEBvk
/UbvRcXnXiR2HfhNOQUFANdP4ZEFlihzGhdZ1PgYdq37m0F3Jy7tankAqMSCIcac
wur4sRLt0GrdS0LBBYdftVe1YsVrG5zOkicFmhTr8xS4UGvkg3AdFdL/UslBP2jL
9Bo/uM3TUTTMmkL2J7XrrWDmtBwkZLwUCh7L0Uh7NB4FTKst/I08ns3cFImPmhix
8ZDIkOlINEkrv/90cuGf5Uu3ejsTYwiN6hlVBlhC4Nu5IY2ItbLr7cQSBjlZF8pA
2Ht4qjBvQ6wogfRpjYY7ofOgrY2TnAC6nzZNQgrR/rBaZMxv3pVJdovRbrQY5Qy1
/7f6O3NvPIZJ2M6HAzTqnVDe12gs4XGP2+tmJa3/BVRvRqJ0iNZlqhtNfqOu/9V+
Ur3F88sDU4uWHSUz+HIy1FXTKdWcpaJCebC8SRCihyV4+aIWTKmjp8lP5AxGVw8p
GgtQ4UhZqeVGUYSoHeQ5dzHYANjIZhjaDL1KQtlOIwXOSd24WKKjSTkdmIaHLBsz
Hs7oYyKIEb1Opl3nKd2WMGjopl8Vs7GU6lY2ilLOUJV94UGpYVKFmDbQBcrKrwjj
/1nVoq43GTHJfbQDUcElAj7kiGjwcaLpKr+sDi0FuBoLFk399h57PHOI5H38QG3H
esPnmlMHJ9H+f1voaGLONmaiS64kj0QvPCV5j2X39uyDx5UYY6RHU9FnoccHbaLl
DqGANlNUvEoeHNu/G01G6OyRONsjcq6eD/J+uMTZBte6ckKFVO2baWTPaxb/5cKe
bFIMOEq+zOtOkIg1YjTZ7if9o6kzkVmBb43gzXs+nqSYeEI3XEIbOz+r4fhinQb/
UGbDKPUYflO8i24F0MfDhX1Gz8ESxSIhX3qsgpQKpAtXQ+m1NCP/BAB7WwoH85xm
cbUv75UD9cec2DsDHbLrjzVnXAxZ/yjnQbHBwlDRsazmbHy0Kr4qZHAtyY0KABhD
d9jpMCHg1d3UywB2jyLVAN569Aneic0LUpsWBsRocQqKLz7UOZZTOueYqGVf4JhF
7gu/ojGARBYq8j7DlKK4qpLjkEtNx0B4aNfMywIBsX0a9eImGjLj3BjenxCW5uDJ
qtVVZYdSPPS5ZHx7XER7SZDIiMnKtzti3xhYEafa0bSigJrgS1olFdHgdT/fypm+
lbuUZSxQ5K4wW+Y8nyvUKodPc/n1o3/L32lRUA66Mh+l7ONLqMxgBpWuZmIGZ8gA
2VoX54qgtl600/T+//ExDAEANbx8OWGIlkwNzBpfGbCj96eUtcMMXR0yrygMXwFm
FpSY678NYpUDYdBGY1+p66roRSaIhDMFyzj6hH3TlScAmCy9vncXOmcxpAyVO4/l
AfcozwDSFbv7WZy7/c5tsTDB2rBukaRMJtKiiGgOiYWJEM3JYAjKZP3V7H1AqGIB
Ht/n4gQopTtpyrh7pfWibu0FvgpLcA3tsiUKp7Bvxz0+F4zRByfrh+9sebgypeRO
NYq38/jo13/TOt33rhhV2D/IupSXi4IcjJwzXCKSn1PixvKYW4RQ/hzdrRw4/Wo1
nuW8rKcRVuTbfvjqoPbzqDS5afV9D+ahOZzB5zKob09RTLoGUXNCt+Un1OJD3iSc
XB9azx1uPii5N27vvAYvBwzTgQV0ZKl3a9g7AcC7sGdKXcJ89xA357z7j+AxR7oT
UIVvNMxkrPwtcM+MNmOZZUO+mgOXfosmaSF906hjWCNSK4bRp306lyvyFATEpkhT
Kb5sRfMBsQ388jMcGCVJP4qbvbqUHs3iB3xRPBMZKhMNvYA5YijF8a+TUa4sheLm
Ej7auFvY8lMqyWE9bJ+KAhBHbn1z2soB/2Xk+T3z9xvH/LrOFAp3zPiXF06HBfuQ
/Zk7HbnklsugfBcaFqBtMQ186kJYxN7R20my9FSbX86RlHCLXoHmn/2n4nQWbZdz
Ju+cvGZTAPZHJ+YUbXkwDp+f5IkNfqGHlCcDyZImLyp/567baX7tIrGvrsFVJLmG
ZTk4mTm4sDS7n4CTE5P29DPwVFJbq6NCiFQieMVW9mv48IQtzXHRXgQ/gNqXxn22
O5ZoJFm/kPnmLotmBDiz1MTSvWmACWFavPw0ppkMj0jyAG52fOCCRDETiClXBu3M
+tdeOV3w0lJMEVa/jrFPf/mHg/xWm2i15o0PHrzEY+ReMB0UOR1ATmt7mM/cqmdg
rB/mO3U28RH6y+ITU2lwTbf8/sYfAklH56oqdHPcem6HMPUx2Opq0LRWS8ydJBNn
X7VnWT3c1GqCbYgKdfNe88rWcbSyozyaKBymGMICL5Wf7InICBxn++lL2yxsimxM
zGlyzJHbSLE4azvyAUGrMBLVqyYwtCm96bKBoLBbd62q484ctHNY7FDT5xuO2fjB
JP5ZJZFeHatIjiO5XHhcrWlyPhLJijr8PQa+u0jFVqghU6eLfDbAVcGSmXwaFuht
XbiyBuGD2nin2XOxqeozf/BdK2IqIG/XIJCGVA5E4eb0RpG482nOLqVddNZtPmM0
4I0lSqRCZvn2+5L+l8w/B+oRf3uppKiYBi5OujyFO36p7/Q4TQoENbNcxuaO3+0X
elnsQ2z/vjbuaFqo6trBY4U8xGkxp5Ny8fiC/sLxJjupBHRwDLJjOrGwtU4ZL0je
pEv95AmmmkF9/Iwusw4TI4CMswdRgbtM6DOAae/oxljYcCqJfUxd3uuIb2TiwTiO
/x7UH+XMF2/l4/yK+DkFgnMOK3RLhb373KZOV88veIveCwLPDTwNEjPPJXRgxkja
Fh3fL6zAxx64ptSEttjzBYte+8gNpASkBlbkTfyaZKqsMCZ7nApo0DMTcUkL03bm
tcZ+nY8gNgzMteJ/2NosMac+RJs9Som8CQ/Ha0Q0a6XQ+A74rczscsSF3DxdxocT
oLPwNOObx5zCRYcQpEJzOGkzfNfttV69/hLck/l/MI5aDTefng1HhJsuV4oFxhZn
bdtQtRLv7bsJBSpyN0myc3WYWMmi//XlIIl8YIAQKGgMqmOuGbVLzm2erZ9juAHb
RRy1GPrMiiJTxRl469QVOinjczigJT4rBKGiSveOF4OCciKinq6MmCnG4w+kSGxK
hsEeg/vlk0gZoW1dLD3J31nSmzeVNIxtNV3Jz54bs7E1MYAl1914RXaKmV5agP9V
j0DrCrhOs53YeXqYWXA0Xp+i2NLAv/GX93XKi/DDFU+kHlDuQg0pTNdgWU1nO9SC
/lfK5Lac6O5F/4+k3Sh5C3ualSa3sgj8bYK5vr3Qk39RaRTS/usInE9fmGf8jffo
GaEoAyMEeHOhaW0JRBZVRjMvWYFYHag5U6Tk1ZHyCD6Ds9vPr7p5zONahRrYKGGP
gff2cKqTi/m15qwyqbAvteY92PA/oubUMeuXUjsar8LGWRCpGaTuw3blMRfCxzpW
1FMSXwnTVFlp+huy+8xq4aLnpLVyAR7hmsSpo0SQcdR+J9bL2YpYcJjOvtfEar2/
ECrq8aXRvpwAbIxKNRMal5AWLkJ5g64GDZLytkDVgbRzkyfxeMWYn93nZGYd0fuY
QTqAl7eIEeKbnsw/PZooK6hpakPl2OaCwGaw7ojX8FGCp6sLM1e2pdRa518DOIjd
iahmLksxf1ElZv6J/bV4iTUXsF6Q8GYlLvyQtlIFg7vGuDk029F/OIrkpqNBWZJt
b2bjF9twCtISLycbgIRTqHEhFDOPmoDRJJWc6I1KURSLK+v0Dxm6RB92m5aLZ23I
v/9WEkWlAawNjpZRTSgA0XniepSsNi1jrO+wBYzzfnrCpiBos0HSb7OcC91D8BoS
pyOR7QH9U/EaMmyu3SIMzmuciD73g//rHXiUsbzzq80E8S1sEL14LkKkGnFANsYw
9kg7+nu/fy7aLInYsSrtg5oFlir1dZjY4heeFp9o4Jp53Jxf9tR4zun0sJkR+3DS
tXXqPDI+BbxdG0TIx/QFXpzstY7bbUlLhcNhaemPfB1iKxVKMZUIcABdzS7KiT4k
GzxM1YoHfur9OzQBko1XfFuYjAZyHLEZltaVff3/F7ILMAzRXUkmO/kXdBbhZdXY
W/HsX2Qe1Es8sr+GwfEXTWs1hQCtUUwWWyQ/n4T0vP6f1NfyTxeqagAso/C3uKc5
ehwtJR0hHr3L9IDBzPjXD379Phdj88O7OjaKvTl1HuqSfmxrMdy/uVFVAZ28mdw7
ZbdqQDN4p57aEUKSmXAium6CovyTSRrOlVAPoeRXaGfBnq/Xy9ou6aRxmfYQjMfY
2g0F5nj+fL39ft8fRf6f18HS5sXqNjq95L1TZIa2FgFjDkH5FKaftgLhfyH9TBeW
pdcLt7E41qsTTvrALlNLsu616Uip+SE7dW83hny5xgHLbs7mWArxVzvHEAYM+xwD
esMMqUHKjK+H47DLlm1ObfMchwRR1I5rZSTEZu66JNzF+94LeCYkw0c1H61bujVZ
OpFGHULtUIn/a8PgSAea4ngA0g1XpbSoimiGYAQbrVUm0WljzUZHNibuoQpe0yuD
Ag87NELgYHfjCHFv2uJ6EF8ff6sgtbKuvQPfbovnroIf1oN0iP7TvPhvu+i5orNh
+SiV5WviXaIICPOMsE4jnsMIeEKMBWsWCqPC5QXcC7fs/gf+37Lg6IIv2xy7eiCO
FX6ck/T3Ov2PR07eBT8v/uvZwoOIQlgUnMrsWkduTy+BqHTQGhS1CbVBt3ODtSMp
L1Yu0qZqvMhK1Nldl2W7WsX3/CWKV8LKwaTYSioT2KbfPjgWJum7M1sKGnff0Apx
Hdd435EDRLlBkMAlOxn07cMyHAlcL8rUoZOFuscubUCuM6SpdML/63MRE79p4kTF
c6QHRkWy/wqawFZk+2ZH9amNuxjSIdOEzpfqS3LFGnftc7qxhGP/UQKN/2Ev3O+m
mFSlGu5dsCS52NdG7Bs+XgLSGmcqroCMsh/cOiimVfl8mcSTG9auCUTyo8lq3JY9
VbrivASFp55SMjF/C5BB6yXBCeHR+Yrg3ALOgAVuw+bpDyeEk/AkYDvTXugDpii0
Y0i5uH8A22Jjp7BWe3iwG6+RGy/VPiOziVVEE7+PEJHCPaCuxXACa5iudrK2DlZH
ezI/jaCEUcSeSao0pZtR1g9oWP5NUdVmYGdRr/249SuyfBxmXKuQGELW+5QV/y5G
I/4GzXDKKzkfxw2sKZqdn0nyQFuCd6hjIDC3STvImx3P7A0nA9OgZ6MptkmH+SC7
9CKHaQoA1eZ8Lv+Wy4shgmCmmNMuEW2N+OKs4LkT/J1DXU+v0NUdI7/J/0YHYZ4V
VUJGS3FE/8nfT/pHGS7nWk6HVGi9+IGFcTAlFL6dep97JjEpN+QBh8DKmAOCuy77
co/mmpgTWzgx58iOo6Q3SaEzX0F5AMBJlX2enpPw1fOqCGVw/yBjvy+UyUxpfdPu
zwbxSVfcp38jq4waHb+Fj78iTSwQOm4NYFZCeSOylaJ7Z+T5WKeqCK5iYsiphrAt
+bhc2+Msf+WQpK3uvKjeFzn5QKYxGrgjwAXB9q599I9qzASRvzoW5Aol1joMx7Qh
azAKHGQ+2vFCYWg/Nm62GyYF698jnj3KcEtO5BL9u9JgAnLub7JRIDnUSBxD8X34
mzSCmhWUy6BRApyLq8cmamkZxFgrIafHYUH9J4o9z7Q5K3hTGiVnHhpdSRF16AcW
L9jnPdVmytmLUCCx7TExBWwr4wyQ4jeKHOzZY92WIO1FCRMumD3SgsURjHeiyVUH
QIGi0o/7Lbk2jI5QbMkgYU1R1qYRe4KcV5iIiBN4KEq+yGt9tGEXWCS35cdGq4uu
h2qsFjUIyDvEnE6f6lUtvWt9RpfBVSI2yvGyOXSC/88id5qarEEsLPDNFRo5LZY9
M5GhkoP9IuIFGUuslAb/DZ+aSFARiNpVrs+IZ7Z2y+xlf1FiB0nSDg2WZNIyiR64
orpYTB7dPSodeFiG8/Iiu2ExUAGX5LDQP9fVLnIz44bROiIA3bTjq1cDL7pg2MNa
ZsL7wHDOH5ainGygrAHSPRbANZNPkg4d1fas10HzKsJhZC9kVCnjerSz/XZy7Ob3
qb5beSUij2bhcTpjes7qnSqa88YGkU+J1s9K6XZNo+ehexIy1K2nrQFc1RhsfKhv
cAQ3h1HXwWasT7U4RPqMqlpgYVj3PPiMUVDbAHi4cSJWt4qg9adajpDli9EX71lZ
nn4jiPLqnBXpG6tNH9aE7UxokCui8bG81o+/NOZkJzcR3BV0pnjI6yKLzSYjq7um
LwQY9dg9e3qaRERlg9VJ9P3NKdD9OoPK5boX2q5m48ludZLMY2MwLDYwmUfQEj3x
j5VkSNbBHmlnYUtE4sv+heDX3cOy6rp1DqqG7olxbzdo7FwHglKu+HmGOyU6ZBGd
3o7et/suupJkWGNA6RdiOCYU1OBR1kkedPcC1kmfOU9PZnqkhLolJyjsHte+wMux
tVIDqynz1LyRAFJ5NQiWAnt4gJAjsYBvzkulZHRn8Lv+1oQ6kxSrJX3kkJU3/tBZ
MANeR34xQm7UtXY2cJm0Z1l1UfTPHC6JHlXkTI8K2fGN47WV7NjAgy0/fGKJu2B5
ueBOwNv1lG1kKuCTFaUXpRoRnTEVtMUUyMTMwu8Y8PIRvuWEWxzYYQjp7oJZhIj5
qo4mc7FtGedpW/K79uidnxl+d39ihwvCDk5sFf54uS7nyugB+eTx0pg3cFB0ZY1w
dLbtODD92nCBABPhOGc3ExF/AJyvZJQa7FtOu0bNVRdpZih8ugePjybRPANcb2jC
jsh1zSfwSykJc4z8bYzf0kYSteCZwCTqhHVG4JzIbXg4NlKFDm0bPjLKqQIDsFW1
dGKgn9dFla6ZFT2N+eze74rVFNvcBgRkDHclloadyqJtIgOJBNY1F7X3r4uC1WAG
Fqevs+cvJsEHD/Ai0PaFO+SIc0LKm2hxQuIOtW+XeQlM0LI9wZRuGpIAGfkyVo/D
J2+SHLj92/QdbkdnIi8eKXMz3yyEvzbWi7PRom+Ku/TcI1YthdjzmD4/h3p91mSo
FiQ+c8YJjMObJh88V+8NV3/PxiXvax3fptu1/UdpKfflMl36sIzSNs7+iojzQB4T
2ESWnMFbVivR5D9sDFl0m4EGXBzeA0/XKv6JTRsOT/sbmALP6Bkw1x66FzE1CTQC
1UwLOzs23cDO/7DMkjykllidYTH7yQWS+O6YcAutdVTkzTT7Y1R2RvY7YKNUwpva
zIJJwGFO8YK4lIvAJH+Z9FcQOeLn96XprFazFOZqHduYFm7R+Px/L7S5NiLEVlSC
Hc9hR5OL+XUHIkAKsx5fe7UGQ1zZiYItvXI9mrx2KS5jfDTek9zYnM+unoZ98Q3p
YLkcqRwLmkzuQWZhknf6wLmPdNKCWDdOWXnVEw0hnzBWjXkdvFo6tOrXoZAEFxDf
yDM2tPxn7cqCe830M7Jjb9Ft0uAEJASUTxY8Jg+Wp8160aCaIUKWhVVBofuD8ECj
vBw1JoFcDNBaUalnWAoIsryLAMaB6lt1ltSMN0QVFYxaHfWvjFOThBb5bkVj6RC5
vlu6nyJ46zcQp6/to7SHS8dJfO3RsydOMdKBQzjfjtrfMGlv2aKrRHDvzHJHHIgH
ejqsciIuFjjbPYpRETFHorAyo7PJXbQX//MVbottt1HaGB7osP6zi1//QdnNxd/8
LO4S6x9jgggeZ70OmB3RJUfv00s3bVTH5yhKAMw3/qoiF4uowX2QDrJ715kqE4l7
wcpyASd9RcDSRfQeaw7vo67O/cUKxqBDbhyGa6eNhWhXxIeuB0JUi5yn/QrYst9p
O3L+POIrXQw1ojnNwtoAcEQCdTZ8WkeTGoPUUQjb41kr8L6aq55Fi2uqpEn6kfl8
wRbqT9Qr8kgGBqnzRTkl8myLvy5IksuIRf82BdaEXKVgaN4OBc+HInDqp8RukiYQ
5RXEm8XXvEsYJj/LW22aXaWKB8ZAm9F3RFEpLECM1cBlk5C/7uGR2RFYVab0qYPP
1kzVCaYhnPJFZGE/pwQtPu8W1IVrBCgEQRl8dBvaqVFhaF0enhZ1bIlpCuZg3ksg
JmjhsLf/V3pFzvBIPcsHkTBpteZK+vzLBmoE/54+2w1bjWSlkYaUkkb/YfASFd5A
hqgTsGTHFCprSsEPUmHWH7s5HjY00QVP05g85asXjCGvI395LX6DIVEF0tqDR1mx
tr6rZS2C1KdZXyPJ5LV6q/J0QlLjvwEJrg3nOgWHzIc45gC/aozOTqIrU0jgXxx4
2E6/YukFiXCk6WJRgoch5vmMnOK2HITL0f92bqmMlMuuZsR4b/SnOi2F3Rd/AMpo
AyS7ZRDX0uLt29F4wqLWd5HAb4cop+tk1gwSDkMjj9fMEr/onElFF489mN1MalZe
yff6JlbEzWu7vOtkZlquf1FuG+I1ZSsdUvZ7BEfUzDgRujfsKerfls/uI2jjpMLB
qmtgEM2v1CsinOwCI/d7WWjbpg9XaKlo1jJxmnJb5DmKEhd2/5SdIt2ib6xQhppK
N4Z762i56lVBE3M/WcdVZPzncRccZYwpEsAbHCtKdFvADMI5wk1kro1tS7KtqL4L
0DuHfD7b4x/h96MpWNl2KLmanwSGbVydEvPeB/6iuM79uRo4j0c3AzjF0lke/gEO
gMj0yOdin7oaL2wL7kCmnZAPdCqr7uf8uQtmD4cZN4LoO20zchFXyyrV77EtPYnz
nfmDHM0eEoa9do7V7MlxlG83T/i6dV4FRhbnafKeKVXCsbtZ6v91QC1Y0J+56Vbn
lWhJJH2W456qpzuj29vURQRyYg+G9efN7vBJHQErs/ZBh4X7IR+d2iid1FDvNBlO
Mz2YWwBepkNGPqwBjdqkLq5s+w+Z3/ArUW7tnKboaPf5O14EnFhbPoAtZmAfuqEg
+jvCRHVIPc8hJuTXLhqpEnw5+V6RFKEHz2lvQ8hApBC6yo+g0LWNEQVpiKbE9gcv
B8jPOUmRAkKT73AcRLwedwPd5GcWf4iLCIgJJ2WpW0lrpPcuZrDj0Kv1V0h0AIYR
Vcynsp9qdmbF82YGVbAXT8lF5uYZg0NFsQlhGHfScqzKyBoRIMtFWil0rHuB9lPj
RYQm4QD7Hm8oaMW6/wG6bYphI+nb6YeeWZR27glIsqlrt/0sG0n9G67b2PMdoRnK
dB+rhMREzw57tx+p2x7hyXmoS5Lsm8UPX/8TNRyvUCZoZzCbCm7qbh2uFqdQL+E3
YE24aAvkRzwPIIt0g3RqSR2FZngrI+mIs9m6TzhMSj3Tjx4B/TzaSdyPdA8ZZXS+
UMDef4/T6pn0HS68dhMpwI0lxhmJUufJcDXSXRw5/GGmaJOKPyf7HB5JXp9XygX7
yuh+AI+LeI/qpZ1R75YRI0uu0jDDckN9rKjc5vmey45Zgsq04/m7KQ934pDCAzv3
vDIiZGYGrhfI5+SjYvf7gjr6ihtlkz5cw4kLGGZvhZ9yTW270EOv/4B36C3VO8NN
bWL5AWhEVIu7b2JnBpgGPO2cInKA8B0eyltxySkSxpNJA2SaFB/LEnUg2n5t4IAH
obUa61VtmHmdVms6R6i7Y67Pnx/hxj0FH9MHQhWuxfPWTnJXD5DVyRwOzs18J6O9
DQutu82E9eAt0ujuGRGyzvHIYt+GQv0er2Dzbi9hNWbpSg00xr3korKu0Tm/F1ZJ
PBFdOrWN5hkxiSnDUpTweiDZVa6P6Lz9YVTBvhCZyx6bICdv8gtZtzAWtqIRnqL4
2cMJxfr/aLBpS5dyKphM77TV2fuRUTH1alrJcciYQcEuF+/ZOuEBpk9TTIMj2xIX
R6sXgXl1QVGdo7YjLgfuK2+AxCnCv2A4fEN2AhJs+ZmYLEOoOW3MYzq/loZiaoIE
iw8RAdfQzGoMRgJF/av2xSv2+CbBMkxm8k61jkuzfoGegGh+6ev9F0OGjwz3GdoD
26X1i0Pcjm6uqB7XXqbTgXvbiIXiGzOMTFnkNTLzjTbmDGo6mHjJntTA5NyWAAVF
bHcSvkW079n9FNpkZ6YUsogLWyQxN9fd+7O8UasBck5TrkvTOTEdHkrhyIvIIXqe
2uw74EghdA62SBIjoxz81RvAMuNaf/4SCdQs0XT2W5BNiWeaRBcmqzpYC/BJsqTN
xe5KMeGZ/Loii76gUGX0uiS2TyKiv5qkFYz8fTFRKZsyERorCoa3N4TCim3wtLhR
VYr+n7QQYdAL8g0agKn3JBiZEexlQQ1ePfZIZDJRz2m61W3R9s5/Kq37gNT/m9ke
wKq63GNjbyMSYVB1wy/+oz01zIPF2FaE/29M9XXn08zl3dLICOApjeHgypScayCz
nwPRKSXyqbXGJAC9oFhZdvqibCJafl83B5F0nWOxEJc4mfuGiAR35zYdw0fwlPfq
21NNeRBpf/Dw0JX2mtWDAa5QhDzC9VavRIR1sVeYEgM2qxKkgKy00Ere4dtifdYb
EApYOQ/eNSQSVR53gUbpMAnp+pcA6ZkvzbSTNYVA2l/bYW4gy+2x70NEsd1YzDNv
PzNikAyh3fonFxKTyxJ5xDNyp7jwRCJzTxonRI0L2DJTYsM3QSjE8WzntPr9VbBp
uswH3A6EF5PjEgHln10oNfkPnE4H9V0cBQGxz590UnH9JBOiYL7wOspsASLg5F3O
Hs/GFuuKFTtEutYi84F4A0tN3oZrcb3kRx49SlERq4Lf876OQoYvjs4CxanQWOkW
KP36h/422WYLjD0oN5fHOWIQgpJIGFTnLOVTI5PtbXYV0yp8QLeqKEUWxSRfJZll
WRxpDkbdmqzf/cIhF5cx9o24eNTt3giSxFnYoRx6lNBxHNrcjk7Bh4XpBRAlBUMT
8UI0Pb68b9yxwWRHFUqJSLe1lRAYc9LE4xxDPty7/WGrwwyzEzq+MSJJFYSe6ClW
+iktnzYIG6eiLPVbi2w5V7LQEN7Iw7uNJWfELRN6SQhjbEenkyJTrz1PQODocJcC
uhj8Lfg8YLu7YmuZLYcnygRywEBKFQFHIB+KUiBia5hVnN0wwm2D95M7Vev6FkRq
UZqT0BokNUA2w9x1pMoj6ppS6LoHg08Z1Lc4ptViKi+l5SwQe8+sf2PDdBIM5Xp4
7nHml0hqS9xbn3/lVRbIDzJeld0owCuQHCcLbkSED9nr7RN0YHdlU/6fGBHaQsIJ
ObQaQ6UYhFsdF9jGbGYGtzoZOBh5zeXfuP820Yr3ywCnN401TJfE4sfY7fTwv7lR
0kptF6Hzir1xhT4s5u7WsGCiCu2ZGjMsTobhmbXUBrVXt5sNPMPBOwfu5tl4s5sf
UWHwYcHQSdA7dfxe2RB1Gpj0bUZKt2WW2s9TsVYEZZKtA3rP50f36+93YVm6ukjS
zkrNSHIzo2QnihxOxEtTWlj6QDKfi8rh72FZvirDywRJ8Tb/vZ7i7U0YdgwWqyKI
8l5qFPyjn4O0AxZzhvJPVqzrp5l4aZb/+jMfKoj56zadAa6a7D2iGIG9BryK75lF
4P1RR2wyQsiPCclQPsgBmTVWvWbKo8CBFoKU101j6ALiHEW9vzxnR2PG3glkH23o
LIiZRr29IxyYbKuAKHZtWGOgh1drkF8RBrsg4/CyOjfFeR6lXRqA1x7Wao6DNlFv
mmdiE4aU97QS3PFOstqMuom0NcjBd0RtHUHAJdjK6hTVNEKbM+yhNY5ZHpOR2+kk
+CkX1/Bsc2JPX9t/sv7/yVioGHt0Qfvv85L8OfKQpwBG+pL/okId/EWLJOJEZNuN
EkolMT5EZjNGkJMMLHrhakZ1IWHm5YsEsVx6vkChF0Y/JmF5BMoxf01A7VdV7P5+
ebueOMU8qkPlyDJq2EUJ+0Nqfb8rsBSc5ZeH5iuUPUAVbAWhr/6HCDujf8bHi95c
+vMlaF6Jo9AyPmCBqUsVtD5mb5n5qo4DRVFguvUpnduIb85kLLyjCgu85xnIn1Zy
ihDHFUQnYcW2f36oVGyDItM4ZnnOUoU/jJJ36rjjmdCSDWBtKystWu6zglz30fRe
gulY2rEZRRHKANaBbRDV2h3S/wCHicLqnM4bPN9O5BqXrNIJpw0LDyj37TUNokdu
jsF5C12O15txsHxHjUiaHf3hXOtSwp/Q+Ynkv7gR470gKr+E03Cg1cDzdgiV5vLi
FATjKfeqd5XiQccZYg2IcA0ult6gmzf4dIKGNSpyUlU2G8Og7qNr5m1zVGiz9EGk
VtQHEZKvIS1cszzPeVDKQGwABP5xM1SsB3A4lJgZOlbkDEIoevz15iTs6Ig2R+gW
yIkosC/0aJ64mkEo+Fr8Cv5N7dvf4ZlvIDfIt11FfZQwIi9F5NNb2ik77uCu/Gzh
bjOG61ED4C0FHQgQ4CdSu9+iE8n5098b/mbFPvSsm/hF1NaJtYBqqGq3x6NIe0Te
KlCOu4hwTVrSliY1bCuu3BCPt2X1EWEAQV7JqrGtXUcJHgBtmVMiKquQmOxRTOs7
ShZKE+x/oAZ9Krk/nHs8gnOa8Ka6vjnDyaGDoRLk75cRS8/oAmeS9jkH7jnPeOkD
kVY2+psVzJv5/eHipM6DLgtUv8jDh/dgBD7/Ha+MzgYtg4h1A4WukTuCiGPgoKaq
H7fhhgFa0Qu0q3t3OT0E7Ig1GP9RD9vgDhaDNtMHhmPDDqkuP1/tk8auxdpyrAbh
JFN0Ap08HQLiA49DD0RmISCukOqTSrxqZQQD/00pOArRPPKjguxRhzcKGvy4zPTJ
LXE0o1kYdw5L9SW1jeSrEK0js6eflgV6c4Bqr0tJjbdvFnBqR6+RPkgVebDP9w1Z
yWDbtEvKEL2PZSjfsLvHObqAc9Df5LJTd2Y2HRsO8mPxiPWD1H+/6WiuZx0DPTz4
EXKWDL4XFhf/OO0khRG2MK3pj7zisXmJyaU7FOH6JxkRiYudyfFxusw3EH08lnJh
oy1X4OEYhKZbcPiOw6xcUwkhimuM4fhVRfidQ6SfZaDHMVKd5RZkEgZwDUwvLyQC
qNRDx7z827V5RbhQv/EeVqSQfIIRZVuSa2+oW04C5uUDzFwgDydYPZc1SlOeEZMl
SN5uVdehJvCpmXlRgkoViut2L+c53smu9KcRU5YOK6IxrKl3oIzBwk0/NwruCg/+
tH6foDb49pJc+InOBVSKg8/sOyNev3RFRaICuy5vgQBaniNBB5zqc+pMuHBth6+N
9vLKLXXle1rWTpWFeISYq/OCoiCNFxRNfdKbTqqOp2to9LQF3AzjCGh2yN4FitrR
9mz1KiPEcq1r5vrCpCcfj5xbKcFZhd/LT5xYO7S1Y2ezcjQBncJzvTMEwxUPow38
C5M0VXjAbm9TSuWlUNVtCUDOXi6gXdyU1Fd9HhL8vsRcjpiqcPKsnWrW4gzpA9p/
Tz3qTQkJKtJv02ZZwOkAKiJ9A4G7sz13QbJ9P7PTtGYlHsR7UAf9s3IVeihc3sx8
03gDVu6ld/2dt3A0iZs6lwYSAmRqYE5HjYFPTic/t80XJSqWMF/Cp6mkzvxcL4/B
I58hiBxjgDKeHaLNFB0TQ9OLutX8KFa4lnVhG42EKfqvuADUJYs5afXt6ycuh5iA
B+Pyw3b4fQ/axeETAqSVEvHO8Vl2vkYHatodyJsYnfgdQHq90ZowWhU/pHoa4dAy
bgnPi77+e/0m+iubT+hZQnCOb32h+1cmmk5sZudcvs3z49iK3PWxdGN2yzigpId8
mY72rcxjKqKx2Xo/y42MWVKdGRnNAtOu4f/Hz4PZwEO4rcBLdc9keZYHXbUogvX4
1VdbEoolzUUSfgECo76R+8k0prgCOTdhqr4YhNg4D4UE2zZafUOpkZ+BlsPkD5zY
OftGq8l9SyLpNXR3pIRsV1GDXqMPcxZgoc5fU0wx69PmjctGwsTXYFucDpGw9hE9
S9kqZS8mMYm3cCEAxf8lqU7ZitGuRoI9SPVaUCmqsrbxXryiDTS2/+nZYcmZbB62
c568UOfdu9w8U1TcECj/4oFEWADZnealEZ5H4b5R8WTfsykD1qlwyWMH41674A/4
aJvoN5YezFT8R34qxNoBjp/zIUp220S9hd49RpKg0ZS5j85JHIaDzIbR3fDyJ1I5
WN0IraW2q6V4G92wHPAqA85Jc1fL1UvSZllhiXXwayzHQFsIl0BM9JObF1g122oF
tzjVC1dAMIX5U8L9sT7EJ2jPjKcKoIMfs/KkR6XOQKjyyCESR0HwvMrDCIoNEG98
c8mmBGJ83AWZkSsNXwlS+jf/6ioGFnPwDgT7i8NPCFq2jUwr2OFn313wzyHjpRu4
fhVUKg38pwM965mTPDhweOAhEioSOA3yBNMQNpgSxNx6jbugHgaxAVBO408jPA0N
V/wU99FNT8y+hgyVGtwHtUwkiruR/MlLOcST7Tu2KiHJ3DJNjZqCbmmvcHDbs2dj
ftjvvnep9sqYO1ixaWUyych1enbO9fZj4uDvl1hvZ+7iiiDWQbaaUKJEFRXlHm4T
rB6ivS2fXvlwGZsv51DB5gDx7cUU+MUlKLxaXnLnYxvtdXHdkIUMRfDZxaKqxtHM
vd6W7/3588fpOdodJi0FR3wEYvKNTgK5iphFCGoDSVbgmOW3N5dDXwPBHApnwVXl
PeN8Z+F5xEg6Sr8B4UTKY18W+Tv5oLGwumNY2facCaXGthmkZVuPFKx9m3B4oaGa
qzt1dHTjiXhMI/xX6U8aLpY1IxXLg/6EQqz/86qcEoCsngPkJfT9Vs4rwR2T6l21
PNZ03ysVkgyO3QC49n2fqY+U+7jPZNV14NIzjFtPyyGcHw6ur0ZSo/ZvF0E0aiSt
kzpXbj7UBo0dNr3G+Qp5HkxD6SgfZnHuJo+JcSZHdoC0J2Rtq8WONQ4hPE1UNh+F
1n6q8sLA3LF/HOgJL3BFiKn2iRwsEVDn8/5Ey91LZAnAvZ+juhFYESHN1bgTPdYS
kIzYCRfzR5AVHNeUthcLLpoC+alP7obyo3ye0D2LKEV0CpkJOep155kUIGFKLD3L
zDy8Dg1b5uC4diKM2546ibA+ygwKyB6m4MOmifN8xv+h80hsbFfBGxmIf6mht5rr
FW782YpJtI3C3jQng4bBaljMbxSUH7rPPXnh784qbim6oO+dfyxmb8GqWzw9Fnez
PQGPzW1mdVxXQnjgtu9kEDKrNcoFfZ23mBYSy0rfzoZCmPaifoATPiqk0s7UNcF+
8bMvYWIyAO8mefSVxmca2hZpd2p6X64Mzu9+jFlWVwjzY02KnL0A1Is2sxjIIobM
AWNcYRvhl5UqAZlOEBm4npYf3fK360YBzjq4yFeJyVlkEseF2KcSjBcZQAcNtVS9
X3jb14VJy7NxhJAbWe2uurNcXJdfO4IMLIOhJ0WvqjMTFMBupyvmqwlnIGMrGz30
aEogHYaaB5xf/rLp+zQvPj+dAi1C5TYdg+t8MiThA7YmuQwhQyOfTtFvl0dpiTMK
z9rCu3LwlAGfVTK9FQ3R9M0jOGx+MNkpSeUpadwkSjqgC/RcNkRAcTJEybNaDrQJ
RRc4ddY4hXYZotT/549nkxgKgW61iOdyNYZGoVqKKhbA1WZzPQKX2topMzXFoT0h
xmThPWAwJf0znzHI1Qbiir0OGBe71UcwQYKl/0/OZrRej4yjlVzzNmtuim0gb0DO
4xXhgNCeBvm8nLzBQN0xljLLvJSGiHC6G40xzmIA/VehHuDFF9RSpyk1JnE6b8Kl
Yp2TOmruBhgLrunaI9JGMQzPWtHl8zQDfpRfHNRh0ow8UMdQaDOY0emmz7IZ4DqL
byaQEgoF3g9drYol9O1XzSP5RDN+FziXYDD1BFWu0disGHFtjrFo6dtu7RGdWrSP
rHcd5XMM61vHC2i4Omt7ruyyQ8Mld7GT7fvzuqQdhFrS6FpQvsdqz4EgUbjyqmfL
nxb42FCbZR0QHDh5eO+0XTaZIQtQhKlt3wS/t4dglqEC2CLVj1a2CuqhHOoD+03b
z0nJXvF067r+RnRdH/WhFBnKoSZrLUOCW5i/VAJW2GLqVjhA+E1hgXKBG3ZrsLW7
xeeg+++lbxJ2uUoJrK1pBH6YmtXUFKBWRzGhm9WGn3A92nI4ktYw2XtwOzGrcgqp
+JZrEo4PeT7v8nTZGwUY0LlnMNFGfjSupljyxuNB/NXCIKehtfgoBcyEUXK23Mmh
B992STNkgtoGhUaf/yN3z1pV2RgOawlsl+1qziJZZY1dLMgKuXSw+heG73ty7/Jg
g0KY56KQEEHsWsyjzzXSwIOZwg/9up3+5CRL4AUF6FXGgasZI5hZBUYehoiAw/85
gizjCpkkWHofAOhce5TqaMbVgPoJFa2pvozhpHKtQOusNZa+QKIakMECptcYcdwk
gZa8Nc27dFEpWwoE1RvZ09ekJW1lTjKQfY8TVpvAMNtRv2rynf0KfvZoAkrDGFGm
ciVug/I4t9zBuLu+F1EtDI7tfp9Ug+KdcC9WBSOIDbdrBRLw+QtbvXIPjLjS6YOM
gJfZZCV2ksiBWtrIa1iA5rw+iwhLP2Za6+NDylp1qA5VdGmmPOX0Cl4mIE8EHVRy
Ay52o0RK3jj8bFnhqt9TuCkGGfX1LoJObi7+iQjEg0rVkbXqp1a3pe1rUdZOMDdJ
HmXWshNgMHaxC2xq2UyGqf6HraAyb+UANcC/WTvGBo8KdS0G654K67gTc44mtws0
XSYuObRSoUuhiawxUOcEht6MSv1NnO+9CNfntYGmvvtMN3NKtl1biSkrmdKdBQDD
x8eGH1QlaJbqQZBg+KbslBdegTwW6ePqoAHF5OPX/IvaWngkzvLzqak6yEk/gQM2
HLotMvB/LJZkPWlSyK70Xt/vwBhYiXpV02sp93iqfDu24DT1Xi01glqI10tVVgnw
GWfJ1IX6ChBZqJ3Y+Q3F/hEwtpDqMt7/S6wKR5K9/zlkASwPUXkTzGhE7DZwyE5c
GhT9eGNMo6PDDSgaQ77oO7nyKsODs9vPdNfqKR0QzDFwaSyOJ/4Odo6MoGa6HYb4
SdFHgT7guJEe18AY1/MqaPpy7D9OgNs/6PCJM5Zyklg94A2Ym6keN80R1VTD3Bdf
dW7xaU2uWxgv6yTi6rxyZZb472rDwS4TNrRoGDXDkdEzwdhRBXXfJgJDPRHKSeS9
SUcb+8wThZG08dYcFEI7OptefTLZnRgaXSx0IC1uJEgr3h+SVsqt25tWTNLUVIgh
DSBXEZFmN8uie1wrLqE61Gh7W7qrc4rq9Y58hpGmUURKhz2MJ3AZp3NtVCZ61bjB
r4M/T4A+AmE/0BpLZenf1TPnVEoENQRsbgPdHLcTnTG16Bs4tQB64TxnrFW7ZKbh
OcQUwuoQg966fAc9z2fUOqHN63ym0qOvqq05ZjwkpTL9iu0apYHzEe9rXwLS4b1G
rAAVnuspOpGre+hC7wGDbi0EUBPOf/cL+HvQe8V7PkuMaQWspJCenajKnwbPy/rj
1h4129UkffcNyAd5wpTS1VzTa02KnEQ2x7XTky4LZUVwHYC0aTkyzzTHXIeQZDkz
KJ4svM3W1Mz7p9gd72eYwlYZMLqe1NOnIERce1F8w+pRBi6IQJuRaml6ed1jEfwl
OgV+tYeB9Iu2VHEkn86AuG+my3VBzSjUaELDmQREJ58nzQ7sky4/eSufhmT6xYSE
hBCMMnjPzOXv2ceR9KDzvSov12U7LVHNUPG5A2vM/LBRslu2gqfF/sEOhFvcD7Ds
xmzo7kEIm5YiEnror7mX4i2GUaLKjphPa2J46W+EDP9AGrIYuuid999eIbj3bQQ+
ibH/TwBBrvvRrkTnzeM9wjyQtuq4pjGFX3da9hjANDmjATjQPo9K7SYV3dBohj9i
9Op2y6DoglS2xMSn8JgMvewEZgtkqCtxgmdCrekYI1WzjUMkYxJaGjijeTDLLhFe
r2z0j4jxTW49lZFyT72EqdFMrhEPLVMXhQCLisyNz/2dbhzTg/tyxf2q9+eFG75z
YXm2xlRaTGvcZfsKQPnQhhl+ZWwbMxGAwNtGSWaDHruV+YRI3822iVlOThkuZ0zG
xV2VG6jp9As8mWXywD4aaWrmg07Tib+SNoWqIXNFlzyxLUUBxrPCHz23gQmP0n6u
lzEiAcbzwbZFANSpnfMfEx3/kEY+D9K7GphXWHL2OUncuGxIKWvtli9oueK7jqKj
KRehQeVn3v/ZtkHgwTkc6IBOMBE9TtJZvibU5i3dvhKMPWGSqcsthgtyH1I2Bkjh
JSR3VWHjpoLmfKVpb0GNJ0qZYvCxgjGPFQFv9ZA0zjd5c3KOhebIOryJKpk0fpFJ
B38s/H+zusYKgn+HU4KuqJGGhWD/QZFjYMNoI76XPiIAuVzhJc42816TOBhOSQ3d
AJn3Uu4N8nMtrJYzLbYwr15Z1XdevqlYYbftVJQkSiIicotbWWjacF6YogfdzOt7
dj2HACSNGc5m/KI/R8WHaMLhI91fZVolKDKbYiwHVk0kXIk7g1VbhrosNXlitqah
JQsy+V30nHD4qNtz7PJMAmebii6Z/mKuxcr8zznAXJmCCdD7il55knwqZrddFocN
kAe/toaQqBq2Uo9Tao4g2MuEwvqty58D2r4R/u2IfuS5Fxq9aCjaJfLTFdKTMI0O
kW/l0rIk36hPdS/o+q2/C7JOtPSFhTTwCmaUfwFVTrsyGd4q0Rs2MhQ/N1EXA+Ct
rZupXESXrO+DRt6P7aoa98NyE5euUI/nsOJYdD+tRTN0ku4+zyEr0XqpCZA032SZ
gfvLjgOvh4HpB1Bbav500BYxk0CtlIgx7wSvmwB5i8Fc2w173UZ4aKol+RZkYpmb
scTukQGuBKTe0yaaC1YpbP9jIqu6+0wy0QwCYNM7ZeYZYMfJzbezhcA/T4MNp2Io
c27ZSUUut8nQq86yt27CJyEgHDYZV5MlLTj+VbGHdI/05cpLYoLCfs4XkDZ8zMR5
RUrtccME08Jui2gnJMnzEibXr9d+OKhAbqN9vjLx5CcvU4804kcuSrjbTh/GZ6PE
zpqjqmhAG0P8fQhOTY1FNqNjHrDNHIwpCyINbq/RsezzoYEU5Z5QF+mUQP6RTh7d
G3rYG8Ysf4oIBuh9gfbSgrc3I5ryxA3RqTYfNDktPrqgwuAvxAbNRCdBpK8Ogu2U
5LT4XifQszxFEtmSeWCHZuE+aMvdPUIoSP+YwB9syOkJ9B0TU3pDiKb4ev9ZCUQ2
wWbFDJYPTl7xGxBbZrC9RnlykGnlWZbyy0IRPqKwfvyYMi/QeS2AhGXavuxlgVki
gD7BxrAt9ili/bbPdNIalMrUTL4XRWsMzfa0HEiDx6DgDQCMxDfDnhq5SI8qkRnH
ne/8HQo6pi6tMjw0YPJiOHpZ9gMwE/x083s8kB2Vft5jpFn4ZMFwHzRc8gM9/IGg
lFnxB9st63hynBqfEjWuA3nWMyNZTr0cGrd321XMuVE9DL9NR2wftTcYtx2Nu/S4
BQhJAr7Pa9ciWLc7mQNvcUDRbzz7kSzb2cfnHxU6PgZrmyf+07qGLitbjKRcorzH
0COX/YPjFRP1QRPyBKlHB0ZMAYIM4D0wGiEVM3oWLlNbHFQTaXwdnLNmpnJE3b1e
sLIdlPpDu6MUa16Z/EDTMWQitv3kV7ZaGUYOXnmMMDFEbxc0VilG9+2PPVK76CvQ
en9UAX0le1IK5JS+SM48rnM+/ny24bEC8cjaepSKGZTzVA+3kjcqNbuggMsqNIhN
qnWFRiTAnX3zm3Dq0KUUcmqNEtji2Ho3Ut71e/I0GU9+i0RRNAjo3W5MufwxwIbE
YykHsWq4/RClo1gyJDRWV1/c1+wGCTkrcUrfJ+rBjsQ3QHnHUTSqXCyVaE6g0Ty8
rYPL6J3+VlWb+o6TzvHn5ri0frpS3YaLJeih06BB3ZO8lI3Gp6t8m7eqFAyk309a
MSQld539M6eni9hI3OETk85VU3FAD1OFh+Q3k2wFFymVDp2v7+Rt+daNZFjAKoHg
QMe4i2T1h1b5WU58sOOflQgeTDgymsRfGePG564bp/2jdm7HRSu9GIj7jbOvGz+w
uMOz7tMFML0wPnX8hOs0A2OP4x3KU77jc6UNTdbDmD85oLwMo0g+bXj2EXHBl4Ee
kPt2JC40QGDuqvN3R5CEAw3sx0ucfojQZaqGcnraJRCsdT9VptOhYFTOlnrGYGbI
r72YnSycoxTF57pblIyIK2cbgjfKTckvNKeq+w/jYBVpxNCixuJuts7DCzXX6xAl
r+VzQvokDUcq/d9MWVLovQoMveaqk9Bvqgyw8zRYsNh3gbjbYt3gkzHNxijLZc8x
u65rApYdFS7LR+7FqZG8vEPYKCFwfNcP51RSYDKc7KMlsEGn8f0fy/2t7WSPOdqi
3b3HCCc0weRRo1s1Ai+cdTpEcPbPt/Lv+Js+1dFgLP7wbNXAXGYtHmE85PLr5LMu
Z/E2jZ4Jb6pEmPHTImRDZWYS5hKcWhpx8HVuMCI1Y5FooKbpywknG3wdECRUphy7
8X7zmqjfUDOTM0IjUWQhiM+4pUN4YBllsGPIXFZ1yNo+zB9gkXfhq567nmJwmtnA
1bIeCRLp1FbbV4F055+ok4LaazHIoTCPOw7vikM9lDzp/NNjeYY1AnbvqWZv1/1s
Jifp64SbyXgMBzf/5OP3ZYwYjq/6i+nrig2DaprnbRQvTmUUQ36bskBe0T2++dZr
qj/fkxTgxAiEGby7g5ORozMsmsNg5MY1CEyiRbAW+LEMtKobGtFeGbnntH9QcrnB
2qQI/M5n4MfYbatPjEyWvT8B7XLDlM8J7zokmghRIcqTeJ0MZBGw/YaCILdYnuMd
buszfWv/l3Oxw/TM722A2kaDAZevdzyLVrZ2ib4qMEVGoGaqAa8ZqQD5kM7h2rMq
4lS9v7vtrJ3ruVGZdzGww33efnih0lNFe99eEb+kwfd4OL8flMFZ/g+3x1mgYhbr
ko+3jxv4fTa5FwjAWsAn1lJPWagg34lrIi6zVzk0PCC3ZBIKHmPaXAGrPckzCjuC
jVo/qOKPlRrpc7OjXzy9/SMPoha91pun1C5LIcZoQrTdNwOYKH42kvLkQl5f4Abe
q905ADZrJATVOGYOcP5WnuKiB0Fw9WwiiYWfsyRD2tsYtcE0VLS0RshM/sgdfe4/
HduvFHYRWoufn3+yi/wxg1dT/vTMwDrqvivVrNv+TDO2UQwgEdUUQOVFQFEWzGnt
Qmg56nQy21hvauj5b1/NXckA8VGtoyDUFGPJ6b1q/x1UWp7EkjICgG5LJ4kw90WD
qWVGyJSHJSCedl944mTO4W4sKJiRz1TVVJWnyenT5fiXkS0dxxYw1GkmPRO1whfv
dnjcqFVGT79F3x+2z4uZCGaXIzwylon0eFv+LP1c1lwcazpVUOkuJEhQ/s/KcjGX
MGK/HHs55EV6gd4LUaCOVpge+Ku23flPocMcWabShlQS8vqtsbgqgqmPeof1wzyp
OY/OtIurdVMfeHkwfURGc3E3fEq66Z/xBIX0JWBVBVHmgW2+VNgHTrQG/QwgJ/rw
pNjMnqxMwdtm+rvwJ6ovgVpxvrSjVAvV/0vwiiO5NkzIET2Fdf2FLC5y6VM2DBGg
2K9B6ncOlPLxgn19yqLuwi4/Q5wh1lMLa5+sjsGaFXhrk4yqft/25yH6BpjdhCMQ
R/kfaX3iWsOoEISB8WuHyzZjWsxnMY9v5etnRmfdBgFrqRB/3rUyWffLth/ofLOQ
b5jIaE5kHmmIiiZJkH3yovtvLUSkGYYHwVlnUfZWKm7+VfwhHjU2Hmus70zTepZM
wM566TNHyA71aVbAUzVUYl/8HLlcHcJ1bp26cgR0b+pdkOIH6X53CT1MS2B5e7aL
ISb2cy1NSxQxvINLfo8bleaGjZ6HizNJPkyrp+ZpPmFY0xJzjIUXogc/5JDq9E0m
SVSWlF7zUaiAKkww2LkP6CR1hwkEB1fgIxY+SlwwLVretikEBs8W7JuXPWKwRzT4
rfyHtSB879D6M9dudUr0cM3JRycnA0hUEpUjXyc1XG08GCsdatGrMfK4+DK92blD
jSPg8Vu2ZAf3g3Ry+EsOYP3dGt5POEtogNLj54a9EpPtHy/6Y2ZrcGNF4/v3Q/R6
9iorpnSKhF7A0wXqP4CJRKaVdihucfz4EBFcFB+VQkpGiv5jFNhjUvoPjnFOKIHZ
902LKC/xhbCV08uGsDO8S1XJrdfeu7lCoaYslBIWgrMW6wMZrFmwicMVmmJnNAhc
t7sXwhDPADHRxBLXsQpyVkhFrMTkVItgCxaEkfSGZYzT1AOV77dmBukDsscJgH1T
SZRhyQresKUc/dYYru2WTVW2FPl6t8ctC+taACRy4IGvChF2hAwRbxP3MWtXKr+z
yDnaT4RzlVAvIj4XPKxuWrDOMON5D39NuNkSvVYe4hcqCOhpP3ypP37IHjuAeAb/
mQaADk3DJPCMjLb4+evuZNeBeIUTgyHRfe1PW8m2q/mFV2vB+3IqDATfFQL9hA1I
9qDH8kC6FBHHR3huMqBeW2vxRk4DtUREMmGb4+mMb9D4BrezBCYyReedZKIyvseY
STVrrRtQCx8MTOaOCwbizIYqQCoDTc4iJvygFMepXkv1nen3XiYzmCjRBxIqPAoB
scP7y2dJaByInDvHo3XEEZhCCV+PoMal/GmLCdlvr591kHAdFIp/Iq5wr+N4PVtn
nZqXcd4tJ/CNVEftZ+N3Hq8EpZfG3LS6Mvwqo3m5P5VgtBkGuaPAGaeoHgDKgsmG
G6gB3IDPHoV9wCNUoCvolOR2PHsI5maROfKFEaWc4QhvXdcb2RbOIBeY4/ccrGYy
lY3WLhm+qJYnXgyi7VlixWr9+pXRFR0/p7LcYfbcuZnQ+Rx9kGRC/LHKzEpYi4lk
C8aEPDdAI9wsva6bBYEpVuhuYf08XYBOMrvqmiXSIobf6UBq95vt05RFczt6fnrS
NxE5yIGWBM+zeLyD2CwvL4kV/Y3zKx5Ourd6NlrZJZR5gz4FWvaIBgKguxgC95kB
Jrm2ced8bDcuRz8Od5DeBah4qhb3qJld+0VYubSnebmfeRw/9MZriW3CLwQUcZ8F
JracAfRzrGzA7AO9W2z9fiODD6XOzZwCFpM3wqXfR6agh5Aa5CkslJU0Aj1jvfR7
Ut49myw4KiQjKetGipKZHGf1zs/YauXYKbSHOeTHaWd+X1Y28jHSbgLM+C0u5yEL
GQINeNoqjY08xigqq2cdpqyw6lLXOiTnA695Pbq4LvFfZvQoFUKuUeBbPe39bvw3
RAZZrsMu79Qf5e/YQuwGjXzx3RSlq8sp5ctTPg2cmHAwW0COeORMF1LDX5pqnWJC
pBySj3/q1RiLmG8LblS28sQdlbejXIiXCbCvp25oxUro9pUBn9hU2KJn16JlNenu
zPYBrt6GqmumU3Ui3NuOzCymSJu4svgKNVxKDNldY7c52pQ+eyIjZC9xoLs6Uyo6
kL0Ca7/28CYfsesOY2iRAjYLRwdfWt0B62JUN0zut17uArjUb9OIJbdkdPFSFZ5R
KkBfFatNA947FMvrOleumcv3la6unaNF88OvRCht9nIg1XNj8XVmJzRHx6ZjHwti
7Y6CxzJqASrATbIkhqj6pf0v5DGXx/oQxGgcyYpPzL2FjC+YuOH8XpT/8GEjz2Pn
qh5LLniWIrUYfJjaIJ2YqvM5Pzyikc3dfY4fwyLUpHrTNP7boh0QWVyTOnjScdUE
tA4tqHg0cRCe/wMdDaHLixJwOD14X/34Uk15IZqleRuC1MkilVLbQbhKmkunKpUJ
3FYFXaTV4tZA0ZTzhLnNrm6gn3XILsrFWyb4dr/0w/ttwYvAAv5OFvx1snU0RhcR
BDWfx/4llEmjUB4HexnykEXAjqpqqUOYBKkq0MHRiMJsVCnpKTlcEB8bzsepMHcm
0XAf9nw2mnMfti1K4Iox5Zv5tfTNILs7VgIuWOhbO+UEg3O//xKyvcK2C/vs4vVk
zgBDmvD0zltlWT2f3lnaBIag0vsqSkFX4JkmRQIeSInV2FQS/cxyalUqOcxFkYJM
L3ocTpzyrDx9i3JrmEBQT+DQz0enCJFyWJtpfQjmNMknR3HGhGcWMOzK3S3FgRvL
orguGBbYo+LLi+kR9nMjjqQ0qEAW/nTq+Os4Vd0cKifcnirJ5edOKEAU9tDzTDOG
vNNfeoCnpr6/PD2FwzO2uxO5ik6b0VcUZW5226Meaug5UszlXhj5R3RvSCJ11pLl
FcerQ8ClmJchIVP1kd7oCKatzrVZNQGosqtjiFkEziOWrRv4FDVvYdTCVwEbQ6YM
4eUh2JE+n+Fq0jFLNafoh7qT4G2eBkQ83RB4jHP6CcFBHrWgiwlEauwG6OjMWr2h
cT1V/+fADHhQ/g9EZUZ3GyjpCRb0LurA1JidWk4wcDiBUZWW1kwFT//NUd8Ec4SQ
xRXAIOZTmNazarV2eAJSHWluk3kEQ/xpgItDruAwoHzKqP94IoKbtq8TFQtXpf6V
tfHnGVSZ3G+Q4BVWpGMJXJ2bnHIJkKdgiMa96Xt4+wA9jbIjus8o6MlIL+6n73y2
NjyJRxo+oFiEOPZ8khKY0S59Xzlmla3NXUZ1AnWWNSa2HAJyQpxx2fHhKecDCUTX
7hBX74np1kPfCYjb3hvnfF2A/NwwUCFW5a/Pwzfv2FFcP/OvU+3mzl6sBOwox/cE
tV5YjhPw6AmWxFET4yXiwL19n/rI6pnJHujCRClPd5OzB+0fIvTj7PwHw9IJfZnw
n62FMmWrhf12f94eUlivwXq6CewaosgIbVNtDtQHlFojskCyuBT0ILPDaU4WN0im
UFy/hcrqqY5fifQQXbq1GWPrArEWkVBgNufDuEbDFkUmahCwx1TPwx/rOOElMWbT
63qJuuXNvJEYgoc1kebvpijQlXEGC8zescnmjUAFGzJfbjejvOVq+TirKcu9ujT0
oM4GUdoakukgvUnttj8aRibTeMapCN9YXjsPqqGXxywv1OTPbUwVxk8LsNhi67FP
PqGmxGbmsUlUxw1sh9ZU74RbrjLeqH4mxmrObwt280XXpgbMFgYobMjCkhTmw6qM
IHPdbvPOFD9EjFuR9qegVBsJuO47smkcygHwPOG4X537qwda0gmnl/ijWYJhMEHW
vSpQ7P0ZPMZm1LHbAAzUwwKCQ9JkPge20KdO+2K5aBPsUgmY848BHU/7LfrsdR29
TR5Ttiz4OvSHxMZZsXKpS1xsYS4Fji+8YyDZt6/pPPDcDtuh1RmzW/XnNe5Mq8IO
93Fg4SrUzN9oHGn6B+nvTFwN6z1hEBmasHCBZ7WEYV4haWYGhoxGtHrRVg8ZnN4P
Q1S22rDsDqDgmIuC4CzJA5pfUzp2GFG8wcW6JU9WYkbtCrHxB8lAfwXPE7jcxVB8
2dUATJUHR3/pAq51ygwkSbyk2vKTSOdm3pcPrj8b8iNSfBdxAq6zp7T9PcNrtoLJ
rfBs+7xmhzpjNCv2Y5dzHCcXkSOV5+JH2isTbWaGAyFc2O939sOEjcHbJjqZ2oQB
g7I2Eu4ZDsfHFVp7kxOqTQALIGI+j/3Tc4D7EobD2PDeYQWpUib6WSPOeFHAxJqu
A55Zrqd/qBNjdoLGZxmPzfDmUajlV/ONA9sdG8fZRZfh6tmV7d7cE0kXVyOaCQQU
dV3Us17HTK62ioWtKr1OEetKvcLgVO14dfdiFi1iZ31aKa/aBX/W/KsouT9HBx9X
UyrLwRcFZ3xltm1dWdoHOP5C2pXbtekNAgUp7jnxQDsnEyzuL4Sb8UwjT5VptsJn
kCE0ms+b9UhzC4u6l0bH83giCkea2mNEp3qHbqUIBPBj7m7A0IG0nKNI5ns+VTg/
geh78r58q0ZwAerC7V+TQrBzGyBTxHYWYoGJMbwu3xMq/mw0aRucZDgioW//bJDn
LL5f6OjvhRfNiIsUkSciXMQXedS5PPvQ86CUt8JGGDx61MKy1iP+QaEkbOxHBr5X
1tR61hTEwYReIj126cPOcXjCtHc9n2UTDeFGrs9OVPIjLI6kg4U0ThIFFr9+FI+4
Ia4IAZVzX32VEWibFCM95WqBfhAM8E0VSYPcLmjUERSvbfxos9l3QF3QlM3hEENQ
ctiQ9ady11BObLr6t0opqYu8I0EXGGBgt24/Q4txd9fO2GSIXAV+pbyl21QpXxYH
UT5iZpHwCAkvtAo51B4iiry2OwjSsRWoFCr8FBnHGCGeJcDgEW0WjwocILSaAW45
qTp9HYRGyQoqYNeAKgn7tFelVI+H77m2Iulc0bOSTTvORZ7pFcxlsRC/PV86Gddi
Skomw3ssbk85V2NbHsuylBtqZpVfJer0VVAJ2kFELq9P0lcV0IQdQLjBk/N25yJU
RB1IrvzAUbdcujKyBdJavPj9epPhHO8NMg+OAd5UHKV9/lNUfEz7MKno/YAXjS82
C97S0Y3I4XJ8IJMM7lSWSZe1Bn1zQSomk30QI/56+6Ftx7jQIxU/aH2QD0dpJtdy
P3BETvDHwc/CD12vDT5Lsj/DpKVJI/rns6qzbZJnG6eCE4m3bbOLYZ1GjvomlKrU
OS1zq5OzWGdoS5hZdrjJN70nUgMCUi+o40P24gHP/6rAPMXv7lsrX7BEF7V2/mNn
HgQnHPAmDyTEmMJ6j8OIG65MowfnJEG2vFH7Lf6QB5m8L4AZrCDmEWraLCX4hcOz
EGIk4jqGNlH5WGdeYY/m93Z6LFwgs4HFy/50CuUOegtGX6RZddBTeNKHYTBJlkg4
HDpDwnLqfMDYC9iqS/t9jmzEveGQDZ0tUpppzJdJltwANWN4cigrdydE5BQwFabI
ucnso11R5I+FHzcOETiUDShM//T2Nq5AGFTik1TQ2I+ehYjUTxWJn4ViHAm/tx4n
z068UHA7RRi86hSNtv/YY9gYtMYAH32feXIRVBPVxp2yOhHk0AleFGzq1GJrwCbd
nHpx185/fl4soegWmKb+EiWUlyTJYJrkPJ8wODFW5m+aapklrS4je6tgQrxjeOzr
gGt/NB9CtxBv8yvWhcHW7V8LA+Nh8TbFmlEmW3Z6qe48LLhlVwzBBlvJpqlZmHVf
0ngkkOJ4KubQ9VKr2L8Sc8EtqIIjUZrfph3CDCZFif/vgw0tTuiW+1fph5uCnlT4
ZUbrfiRUq8qwh6unREsNtjh+ONlTc2qZQW6TxyYutd7HGXUTeJ9l6X2CFWjjTVGd
Az9BG6lAVxk1MaFx6tX2MFPUT+zM3RnPHXg0muP5/c/lN9a9YMZXLTKr9ABCo4BM
AdijEPkUECRDNRz6of3dzVEjvDL6Eq1+hmz1re/qyn1UEmIKl768MmDu+qhgrgcf
1R2gPKVxh3yDuS8H6QV5WayAbbq+i+J3dNmEc6dR01cHN1uPhk2PtKU5+rM1BunD
Pwdb9/PSL4434+CB6X7vypbUbwDCzsUGs7mpKYato1VAWF25UKFKGYGI2TsQA/QF
Eu4NUiashMMancGLi66csECk+iCI6kuUoY3YzxmolzhYFh3FuFSMXz2ltQKuq8di
w2iiYSqJENvE/nTPBm3JbUudr28ITiuuzbqpKf066S/1MI6U855YeqKZe3DlAoQM
nLoUS+luXzDh4n8rjtQ5TVmNmzvClGpAmOW42/uLEKJyLluOfANK1G7XLvnaaUft
i8sqHk0FH5pZ4lbrO/TFtfD8jRdTn0rfdPQ6d2L2zXKsuGgjlxqGvQAphZjZhMFK
Cz+lsfd9vZ0DSuAdqSJIhdXc4+19TDgdUZYFNhxEmAXr8WxMn/N+msa+ScDYV9zZ
gISGiPiEaStfwWxhVUyx+8R9Lkq0VZyxX71/pHYaKx1TOdzMDddV96Q8HMZdu+R5
pja+siH3oWXIrFpHQEajh2DwhYQcnwwkGf7Sc9peFItylZJlnAAOTtTC0q92c2mn
mKqyKwOuerD+Z/p55Lprj30fP8RtUWeGnKJAe2wmRxNEeTZHhgmAQVphulPwvzO8
gPsxSNubT/L9pw3tUb2uRAVZ4zsRe4C6xYTZXFuTeK00b+QvoL50oYfm8tJ8sZ+H
xOz2JXroWhhwfr/RT8Lw4rmkHASLRGtshCB3yB80uMzcvxb4colZikIVq1rUTHdf
vNAGIlw8tc+zBM/K25B41D1F05vaUX7KhF8LK5dQwxGSeboBEiIJ5Cff2LHMSx8W
RLb08xEEzyJOHBPPqUxicRdfokQi3jEG+KEdKmjfwFYb1BX9iZC3wbsC2b7i1VJC
gSk+7mJTBQ+8ZiJJ4R4kzazq8kbJH5V7As1i/fK/CgnDZKDRbOMzfbJJfUjLAMD5
VFe6UvXKUIa+kAOCMr3IphrI+iy2j5FkKfWRhOI2X/5/FjMDNW0i6OHBColvkTRN
Nt6GE+/ljRUlsCGUywMxghKX3arF3EQIUSPAG/+HBeXgSzph1rWkFrBy5JJg8Yea
1DEe6xZyup/wJtUqrTC4ZL7p+zdFIJNUXre+/3jGU+IdmaST9NhTYZiQGASA/xd4
V5WYJ0Pu7e6UsY9JE9EK3Qb7VTYaIgTb8pIynRrUzfU2oaEvOFRnGEzcjfrBlo27
adNYtuM9Zb3TVmaCpFbQ5NN7M3VOPotr3yi3uC/QPZK1uDmHA3NHi+EuUXJeNaTe
pRYwNziDCnlw457yQOsys8rpkSN3hqJh1LwZ1untg4UmUqP4awo2+uEO0/cJgBHn
ImdhImsNoDI4z0TYuMt17V+tdUbF7lTelWlfmMgh4wGcK7VLeHVgYy+EKWR2fwhp
MKirQwL0pGofOfWmBZI4V7Vp2GM/kL1vO7cdWltmtbJZdvDd3Q2HVQDopMZM/Wed
77jZgkZi0KMyKE6NZaagL4tlX46uSZx47ppUwwpAmsEwp6l3nxprLR8RD4/tn+GQ
cMnqm61ojgyfHGCTwtPvDfUH8dJjE8vg4TrCub53PTu/GvMSwCVvFV3UkyiYQHw7
gx66Q5RvpHIhZ90D+eFApV626wNg6XlidgZlnHpTnHM3PWsz4X4CUBJYELHasqh6
na02NrBqD9eYDwA2DTpJYfBu+eNxxgwaQ4zBmRgYdVQuZUKOHX3IbGoW0rGgWD8O
35BzjzmLt+hi1na/9xCx/ohXBim63r8pgTYeGqvKogBA3ujYHFB1aGoGspoSo0VZ
URFv2Gi9nDpba1iYRSD1UH0PcE0RG1NQ0fFSDfLptjD6+ib5Pll3cu9o+4xBuKAO
8Sq+4UuycWGEtyZdDX1i2oOedwylvHiHpYV+f6hMgUUL7RmcoRz0GYpYPWmA7BR1
ZCHSLSAp7+8mkXFLQNdI3knFQtfACSbFCg20nSl2BwAGjlku4qWQ1oczjA4oFQgr
LibG/G5e1gNoqPE3bAEeI2XkkYKXt16HYPjObpvDT7QetaJEu5EkZGqSBRhcQtZQ
DS8LroZBAYs3E+xTpYVXb8vdvPIckobaaQBR6hXQYbOEnnuDC7Fd0ErlR/5pjU9o
G6B4FLM4BWSa55yyC1AlFTBsZg4VqovXQAvw0DZjgLyfUt9OOuocrdGyTLqsydJN
4cuLjqTXGSnYOH5Ck/8F6trpY3nlnHj5wvYLuYDOIpbDL4iDR+n4f+tiiZbG5gA0
r173Uk2n5Q11/nFVl4QyKbe7t1PcBbfVHWwRMVnegbyFz6UioLS4RJBA15dGiC2V
716m9Z6CXFbPK8DzHrIyjksu4c5RhSuai0WxqP0n/LicuMKK898i+lNzuuY8Dryh
xavemFjhlwJVoKIQzgzsIar5mrDJC42f7pWPf9kh4ROR92W+lxl2Re9FsdPhmOpg
Msd1JN7rJNEZzKhl3XkqOryhbSBd+eTMx62yN1LHRv6x7HCFiJa0rAkyccOq3iTF
L2dBHXNOQDnggvY4AJrfDKAFgpFl1kldG/OviaAMmfI97e7kbfDO/dqe4TDmjzSM
bc0wnixcb+ybKCfh7+WFHAhnvTZgT0wD+j48vPhdt1oe+TzpHm8fjaZSSjQOLwZY
fNXbvQeLs/7sTjS39XssCP77pYd7KbHCy4qcBJGCJdJEfEm+DVRpuqkhVs7TVzl+
Wq31cNWkzUeeRlHVLQeI78mzISrCmgRR8K7dxw/1ySZe4+xwk0qtts4kTvkWcwBl
zv3ZYG2KCxr9drxb734Lwm6CtOq/QXk5y4Nd08O59Y486aOk8AXPfbDzoHgXIqVl
qe3llaqFTH0AdPmeO5jGyE+RuysrazxscpxZ7co1B+JBUd9FtnOM7n2S8sPJpjNC
ujzVWx5F6+fhrgCFZSxbX1tsf+Yca3w7l5qDQt921ihbDdxDe08ct0eBYYKThCn0
nuoq3wIrhi1ceb0oEcXeWiNnH9HkzYc/A+cGrZvch1/Vqunjz3kP5I8hbnzp1owy
sNW1fBBnUBvyC6Mdh73wKF//KUjjmNfpgy2FEQ0rqm7uo3QBOnedRR9ReJBQ/kVn
H74jsa/jGRSBUhaTd07EaZoQk1vohoXtOfTyyK6S7Yayjv3D1pU++JHmay7PECFD
qseWNJ37JG0Qf1atyHjpDGOBKMzt9/Ngal+Uh6jKvIFNsLE+CMcIk+ljhbPcLTBz
FrCpDuiWDwlTtAFgtoVQYNe+Cq9kP5r36GndBP/GsA8lyG0r2XkWVnINov41c4FM
9ezm6tCMQIYt217Mp0+vl9qOzsQZg626F1lexz3e0hcIb0aU66p7ysmT+qo2VBWZ
VkG70xWBetuE7kij9fBzs43gbOfhmO5vKRw/8NES/d7oqsvtHvCXV4llTd9jjCzG
JWEolE9b9B4LZzxltlzHmJSOehdSKSLOtsIKgxtJNaLF6vEyFWJGQoyeKLDT3zHQ
1M2sOv3UGt5Fg/cJ8PyjN8v9vACvHwGIKj9ORcZRFHDtTB2GN3yYEaZRMBBHXq2Z
/xyBnpAIunwYPkU17o7i3E86NPIuJYF+sE+gsbvAEDER/BAKDkRzmMwhVrSSZVwe
/pjg8iAo5Cyj9q5vsPigYAdbqjEAvAcDkyfL3KYnha8cczDAh00GZ1zwZdXmQyeQ
M9ng7B2ccj4l/un3djXMplP5826mZoQRgpYLlLP2/F18l/FbrDCdpxL58wOx9KrG
uOeUvbBe3rsvlhDvUBjl05fxy3teqZuY/MZ2nmyYXI1GBatmVYlIkbolJJsVb5vd
gF3MAU79m+c7W48ZSvPDN1UbSYua9JskuBoVGW9PNUQepiAw0drXUnJQVi7oBYrx
h+T2xbrnHtthl+n4ytpURbLfijQgs0OhLubKp/r9gogloSEujw0e2bgAhZg0hcIN
P8Za4tgd/Mp028IYOWBZs2B4bou6PJYrdQYsqEzQZLGuILglrp20OL8fcQAgyq5z
7bArUtrJhsB6CB6hR275Xntoqxc0gZMkY7d8Fc8VnDGW96dd4yZ/9fI6t/QEe80s
2/D++kFt49K3faC3sYJaZANKlemu0liXgRcxPB7u8MKJ/9uxrsuX+29J82gWBIby
SFwaliZs70QnErQD/tRrurIllH+6QXkuJ3rbf8zaPgMJEhc8jAbCqFmTNh32ecBn
KwOk3QWJFL/kbGgg72aVlwT8ZLjVhiFKRv2UF7eJufABpvrqksRPoeG/8lhP2YP6
qPpVhEx/sGfgA1/YHTf2aF67dxsX8RcOlAMA6iGMx3PhzoK4LTxs/cTrR2/M8r6w
FYvx7AGQXFBf0BbX2ToV+4Ap0DpPXGmc22L1gsFJm2cJLdO1l2DyFs8zqDfwoowB
/4Kerop35yMfKRj9vDzQxH9xd3MAs6fGJoagghAcEkgT2kTkFIY+GGQTASbf01kB
h1eOsMG3KCHhVR4IsJJmdtmcusQW98faNfvOa/WIo0Dlw4mLKDmMNX3xA/JYG27M
aZfXo70h20VkvB1ur4drEvgsyX1wmoZAzAQkd5k3ahXruuQkfkZvaDLiD7vsXaVX
1yt3NxKATCrJ15RZRYsP18RNpHTEVteHZlDKlqwJiPTFnZ+Txp8i6VLlFQYrSG7A
aT7z7KoQ4za0fFi3SnRP4hH5totKmazlzvITt73sNprBHE1bsSJSmjjG9v8U+nne
hUNQn9Kv1EaEZp1D3y8gIMxBRpXAPdKeN/4YTvj19Wlu/QrjJu2ARPh+jV2CZFrx
JB+UodnG4coMi7TSk7U6Ziq7JvWP4TuX+WmOrA8Gt6xPQ8JOK8noPShtrwWrgoXc
bsq0cYylESfnyMaJtYqn7G7X47R0smMtlLpJo0cSHwGMCwleIfkd5BL5kLZnTjjX
eMtSnyAjRgArhxtPOTcmdQvpYphHR+oibHJmcH3NyIZzDgx3m4cFGV11m8I5iIvF
nEo6Ikd/+GKl4EwwMnEUP5YEl83UgpGqUe1ECrKwgjeVDcbSexn3rhF7upEtBDl3
0JQJpizaCeUGiDvSRWvbHRU3OpmVSi6cOEO736Q/UJDd3bWNWNaIAY8HyBXfjA5h
7YMOjhdFGzSthbzL05zaAt0JmykpiWIUbzm44Q0l5a+xCmVK84b59ihEnk8+u0mx
aHbhrFdz9QYG7k+SgIfrAeY+NFcXb7Ul6IRiqCiN4KtCTpGvaZbZdYU8q0UYNp+N
qH31cQFO8cBb3EG7kpeFcf6uVf30CuptnsUhLepixUDHgOZuWW4CLbMD3JHCPZrC
Zr6vD8H8zmbPLvDEtiQ/TG8VMH5UQQ85upTu5hyyhYeUtHM2cq+tnabOvEAIk19N
XgdCC9K2MqqInwE7aFujQ87o9F1xNSDoeq9oWUHDrRtcHv86oj8INOWkC4+snuq3
yswkcPzXLsTgZXLRwQRhwttIjrUVOrQWCQlaw7tNpn5VnQW8NblDigg6z6I2BUPS
B4g8YsVj7WdeLB2sR/ETobvIkgparLv7rOssm5oB3wkGxy33XCNYXTL0pk2LNjan
fER8WaLjcp9ZQQZtLMK2qwGridD3yRBqsyakV5v07awMtY+ObNr9CURkLLUkSGFC
TJ+LjvP+YKvCvMcLH/4hRiLeK7bV07r5HD/zhcp1YAnU6Tjt3uIAC8VFJTuA098M
p2UrfMYwnTqSuOxvBHs+sGsbObZRLZveZcpxygjPV2g80JrHRzboWXGxDU59qvEU
xOAB6xNjZ/zTNP0OntyVMnJ1Lbn3FZfBLWBYKtaEsUYvIOPUz2qNwfA9E/hZM7Qc
kUOprCDFqVRSfq0q13r9Sv22kZArGDRkfgzGDGKnR153rfINy0ONZWDe6b205SFf
HPvVQrlTf9VCG75xU5PYUtWnlVUQirWO5ZgO1gzE5g9aLs9wUHX603CZ4FHZM+xw
8M6HOBS+Q8K/WlRab0KTMSXCtdMxe7mTexWwc65JdygBeK30jdtym7KjE1y02laj
EM8cmkYERJ3KSIDj7rccZLXv+IJHfAwhZCFspcsrBSnyc3bVQAGwLmLAwD8KCDSK
9v+Oe3D4gZPRc5CPD0DD6l7WJrItyOh3LBNrb8Qu608FDoSvrrXZho1jS4pBOsxp
F299leIfr9tdnNWmNieNipWItIdkkU2fA4CSxT6wQ9riZK4x13/zc+oCnnwd+Jcf
eoq5SeoUEVGpREJxHXXifwwxjQNFKavZ07Wer+F1u4vyNdmt5ZN5BRmqNQwtkgJn
6LeMfaXZaebWEObj9oi5t4y7NCXnzCI5Ebiphw3s2tgLPY8Q9gUeo56Y530+h6/m
OJx4TYg7UltAqRXg34oj4rMSTasF3Gqryxh9Zdw6LD6QEiJ08+wdpy3ctZai7C57
NV7lnb2KnBprsIu4jJopgTSQCeVaqkXvHd+7ME8YlLpX1Z67fh7YGlDGbx52L/kv
Jxw+wN8Izc9y9rY0yOdWlIPpFJMJ9VEVdQ0bLhWt0PfRDX+lTSercwK+4UzbtbJr
3uUn/rtZ1tpW0n9gPbr6/yAM9EKyjuiTdJd8EGTLZ+9qaD2V8KD8XHpoGin6pumt
amNVYKUdiM6YwxeE1cQoAb7ftqE/QtSHAOZW9m3sZeWJwZIJ6Mt1kTLF0qbzpnew
ROHyhHspoJ9lKkubikiUJyF74bw8zJDg8occgMiYid7MJDATP3/+GxuuopdsP/sw
i7RDoImGXkhzgyVYt4qUcpmeCcH9q7k3G8EFvVf9hB2RcHUtwuxiuFn/fISGIguX
y7jfSiSkBgjYtW1uYN/GcViCjtHXMR5kwQv8ky+u5w11mR5KhKMqlIWE0HstQPxe
VvPLIBfk+0befh7MW2VPyTES9MynEExxqETCddXzn/SJ8jIRmhpBtSGuknNxxwjp
/Ua2BGcxWy0JL6ilwoEWISHHNEnCJgYG97UcZ6XWB44XmX4X+f3xs10u/wH1zfu0
Uh1Hz1odDBPY3BrwgfUHahofDPnSV64uf8bFwFcO6A7zqo9HcsWK7eWH4SYr+tlV
OmddoLww85K86hhsxj8IoCdC07lOS14+Z23c33AN3V8Kn/FARGdx5naPl2RZwfnm
mrdSdaH4+BgV6V3vqqV7DdVVjm1rVvIy4q+U20CT6nrKaJ4sq5Oi1hmJ6F4+Pw5i
s2GB15q/FdsJJD8aXtq+Hyf9yMquIH2T7NMSEzSICIz0v4sG8whAUOjGgrAn6Sv/
wnbYkA27f3Rg4bkW1oTOWWRnc1Oh+qRz4vBpNK3Otwlo4koUD/g+AddJKmS6bO1J
r4GMKe5NxTeqX31o2CGXhhS4JUovTQZ+aE6stnz8Vx20PiitPaChVNBSd/Vo8hb7
RPnxPox5ByUKLxWCkZdlbGzTRv7zwJZD8eIofVTT3qNXllarXs7VkaHSsMiI5Gkw
Jw2TZWCvzqLVXrqANXT0hiVQtWk1DP5CxalpB571+NJjO2QLxE+4ce2+ghN6nLAA
z7NUND72C0rl0mqo2GwQ++yblLpKDmLn2hkCXPBFcCAXtuyYMjRFdh74GoaxBxcY
VUwgo+XfPKIM6ObRBKqvJWCugAXDXwPmeKsT+gUbp+jgPmoja2fpi9tx9LbzaH6w
yU9QUddEmIhiJSuuaEJFAC9UckEdyCiCx5BT3UATkQ7sUJboJuOVfBDJMVjHS0Rg
mFxqvMaTb2JQ6wuf3IdrrL3BnS28HGLD9Q/JTLf+xgAFxOhjYs3ht00JLUNrhEi2
jKL+EpURnmpNdKEClz+6yq1n64Cjkse6XGfugLmR+ZMtSXIiQpq1Ayzrr35lGKc9
IDnmrAPVtKe0bU4nvZS9VwCJDvqavuBdZeVS80NxR5keGl4zxYLgl7L/qFVYLkvH
p4+8cmiv0EEkNvfrqhYUrUWjD3FjX60/GEeyomkWneZDcsQZps9eFTTuzUI3t7T9
/6Wp3PYLRaS0Mi55SD9oJIZBUMXjvg3SCiFga+GLIVSB3p8EqBqA4GzDXGkIG7G7
FfSAw4l+8G/SuHGa9TrtNq2BDyMsl5BGPIhK+LktBSRu40bEJTBGMqomLQJ+r/Bu
VHu9aJjSc1gpKgIDB/uileQngUatf5gbgiKLsoTPo4DBem8ZF4NXpWwEkDU2bPId
vzrebhmfdMJoJdNzM5FMFKbY+xIiMy1Dh2I1s4bo7xN6PfvyOtKoX2e/0EqIKoxG
VTikzzUwWDOUP4r6Te5LZtfPXHQk1NdbqGQUQDxeOOfx2i9jaEjsqZPTmD9Q1MIA
lupSk3rcbAwmZwPw2CwSagxqzyla6adD9yGpO3Mh+8K1J/Fpix2DsZomeqjQ+TzQ
MbtYTPPOHKNWH4MSuoI1+JgyfmA5qptKzVVaI5gDMVqq77QmwiHKSy3CDySrF6zF
h6JFuN3aen6ToMcDMRrFyCbz0x/JelMRUu1fs/Tpn6AubUIb1PZZ+IjoG1cMO892
uBMOQtWzHBHsMRVfrE6waut4ByUTf0WP0P7g89ElJUqyS9a/P5vpKJYHxgeI1OxP
qGiDEcvDPCNj9j6lzqv4HwWcIHW3FGnCXFjk+f6rKK6QW6gbTOBECanoiy5PSIYM
0JmKOCIW9Yi6BRtVQn0gsIUDEYL9tjVNcQ+UgF2wfdVcVEZVu6Z2wIegkNVx8nHY
IMxA8LZrtETtqrfpx+VWh3WM7Rd6TrdBlxupjpvQBwxHlg77CQ/zQxCQenk3pghv
SZxLas6LpHILJFEzLE8CqyQOHchztbJ4qbFpqj39CBIAPS5xR3OaOJdJO4fJfdX4
up/A8iKLfVkl8fdB+v0jcTwUD2NwgudNe91Udfsju/aThs1pO5BbDI5/gWrp8MbA
kAfcTIINK1g5NJaCkn5ktdV2F59TUJk973CNXtrjyXOBimF5ppXGek3Wwcmw3sk3
YVUNDK/9tnL6URGghCUCqNTkb2DiFrHR4Szuj+JlH6zutOFqmqmB5lgFHbGwpCfc
aUrx1Xd0iwq5G7egcihUUBApCugR2qqsn3hd7iKB2BpfKL823gV3/uxLR1PmHzbt
LZdxsJ/y2IhrOMMOdmmoLIo0up90EyMdNfQKY8kPRUtjMA5CxbDO2wzCJ2iyZKBa
bU028D3IDS0EoLTONSfKH4owvV79f9hx3CoA3WH9VNfErdFl2lP+/leQbf3WpSJk
LuNP1/hHX/8kKvbZ5+HYFYmuChPhdY+OGeLg9eg7kWhGBAbGCizrc7jfr8NZjWCn
qo6KdWFC6IebFEUYdgOn80mh6PEpPM/b8NltyuWGBF/wl+LEROKZLA5smUwtwnKT
OohyJmFtlaZlhPkWHfSStaOGXD+jMktFAK4VFbVdVlBjLFt+OzMi2wJUMwR9o3mC
cfxMJmXvuQZkb3yuxfNi8iwYOT6U1gFZ/qPv1qPTbhgqLRDR7j4IYsLH1zjmIfD8
8ErhhkhIgZRfZ22SJAyu2rXDhR+mxtBxOmzIPguo+S6Z5xQcD6K37kCcwNAWNSFf
VQkk1Z+RKN6rWMw5AG7fUgEK0c1BqDm5q4dVUV1nkS2iUDFhso2W5rgNfPikxCxR
7YDz/5wv6s91x/jP1f6syuKpM0PpiN/azTClgRqZiYygzJypp92mV9YP+NlaZUeQ
PPdngaB9Qt7WVgxN5Rr4G1hNr4WspgpaCEVU0iswPdbmCX7IZ2dfZ57qZQAK1J/M
CwhgfBaaHVheX4uraPdrbtHOchCY3+Z4bVbndPc0fVm0FNfivS701tgDFxgjMHm2
6LFUWZqOjIrpMV4c73gyr0DCxc2xi+RiM6rKg+EqGiMQcmWjObYfirETe9tWxofT
5asp0ktHbUMaORBJxj7Uxgxk1RWXNeA/H4bbpFv/8rbY9LpLh7tdT1RVP0zM0ogh
fhgYpELH+2NuVQGYJGczjlyQUfmxyOVdg/hlNeUvJ7o8FqpQaJhGnIFAPG/fJraI
PV+fXluW9mRgFhBVgQk0F7cvd8/bWE9RnyxIvOB1vr2f630kob80RfarEFtrnVPh
6RLZgZSxYOUH0GG6rqjlOZj6olJyYSAnQ/zEK+4MhcRqXkCCTTkncWTPIq+MwOt7
lSdOYdTZKES3zincORvfakufDIkV7/mSp6hcMpurRe/G3Qi36o9hC2zWlwE4hof9
M1Lc4omd3aSEt72R6ltGK18cXvvOfEz5OG1VuGA6PDQTkhJo+0rXLMLbuGl4FXXa
yo6ZRbYrdIl18UihjmNNBvsSVqgiK2Pb1BVOCSsymb/9qrl4wlqhT9k32T59TZFO
iCdgiM6CbnjTQDKCadiGgYVmWEZa+Rb+mdMKdkw1X3DGjCuuHKGLZJCWWLvsMv/K
h1WhFQ/eAI03pzxOUfBHH2LuuHeEPwYoIKy/nDdYg47U1ZwEWqDHeVrwnEPKFota
dFi42+0QZTT/o1IQtOv6Tm+C1LfzTYtHw59jVKykxOm9lLefGBc1FqGvRNiclIIX
s3dFOoVWcC6fugYMbHze7WDoXn8LFEbx+opN7lzTB/wHUNsP6yH3aGeO+UhDTcfw
31SBRUHHLIXISb1mQLzLV8kO/4i4e35hM4fQ75HSOFOsvmFjPSHL/cF0v2rTkiKh
yhKZNKjjk8Hkl/MJ2eUlmsOTEwSM37ghU6yG2csT5G8LhSdHAnMr/S1IRLwPBT3s
HeeH0wX9eOvXaH4SmwQNJg2fpcVQXR8ACMQYpAPvcgh9fx13CbZlyg9/F5IZQIaK
/eJ2WtR8qeMjEao2kzINIaR3lwcqKmNoWB1d/8LwIPj/ULq1aDTTeBtdBM+NpE57
PiT6l3sLKHIWjt3YvdGvmCom6I3uGm/R56rDfePthap5nCgaWwIcNM0hWliLCQCg
hQho2TCZ4PrC6jkxA6/eHyq62sckD93p0ZH4hnmiVLUrtdYqGWh0yjhNe+3vqKLm
Z7dx8dVNJBkfQ7t0NaaAGFAY6Rbm/5YXD6FTvTDRgcj53leWB1BpzcKTqhhkHtnt
`protect end_protected