`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10128 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzs8FhHEQ5k4Wl80hlbK9WdJTMjANf0gzDgzn67KZtbaD
Z/JeutdEEMGvDBmEIAyhmnmwDNJpSX5Ft2kdKHycg0brJsvbvKG1fOZajG6x2YkF
31ek1bGa4PD3gXVrklRGKuyGR9ox6EzvhoYoEDruaZm1TDOY662w+jT1fxZx2qwa
q4Rj2DujYRNWmsukXVPsPIbviJzT0B8BnriW7etyBHUmtP51VOFSx8YLDo6z0HAU
Ls8YPRoa7sqrN0SwM2tWB0EYYfPslGytvgKA0HIE0N1ZWCIPtF7NfQICCqsyJtmq
m6+n7oTO8QQ6uQL/IxjHKhRRC0NJUvqT4DY+V80EpXB1+EdTlrKR/vLHq/wWOQto
BW4VzmcEq+NKZySM8j6IaUjUXig5lJV+XHPW1PZRnPLUwtbg+1ZxtCEb30YMILEz
nYnJHSnKIyq6NdlDcJc4NOa29mu9FmY3a+gFcg6QgjDBihTZIDJ+TO9OBBeK9cX+
/8zFxubEgZ9EMf6l4pB5mlTuvFi3kljYUb7rELfFIjiWAo0tfkf++sxLmR/ZJSu7
3QYcwfA7F08Tg0hX8/jbJe2Dv2tXFXHo40xikZCEYgG6hWI3fWd+9gAowO6wayRJ
SqRcIHvTr4U9DuWJhLgB4tpDuMqK+ofuTi2wH03T+Q6W8hytlNgqiXWyRC59azUj
G0hbljsLnmlQV+SgvNsK3Pegf8gaX8l1/2DJPOG9A6HGxAJXnrDz6vEj1rxl+Fqb
KnpCw2Zy1agiXvJgyl8thEi2z9j7FRp4JGU443FYyLP9jIyg3w+qU4GbRou3kJ9/
gYXytZjwByLveQqrorLry9qPQTjotvY9nNeehqGI1BPIbjzkKos6GmJSUwmn78g0
3DuD8KEb0Q8yQp5B0oPmmaPIfSHT3IPUCKqipyWIogVZRyTERaZ4pMmhdS2CQtCe
Nbhu2hsBvneUXgFBRFFyxacHKnX/14gtL8NvozTtcGFTAr8pE6Vd9Und2lxDFucI
RnUcS+GBtb8wqbEC7VYtNwJ13Tn4P3E12tR+6GSrUKYF9v3k2lsN9Y8YvEwM+S3P
lcgomgKtcQRvGaF1feRsksw8xZveLBhcXMQPGiK7VipepaZmsFQZDz8Ehwga107n
VqCPIWxRBX9uqyV0Mq4+5mFtMZ7W6zSI3bQ1I6KfbacqGQxK0dt79HDICOYx9B6a
lHNbQFTHPp1r7ZSIGy28i2CA1SlugescD0ZfmMkUGCnXnSCVjs2/6x2sWsvY4C14
jEDJrCkOsHtL5q/uNPJmP3Ikaas3lLDgJQci+n57DnbzlkhRY83gAovTCL0VgGrp
FgaQehleFb2d2+rR0GGu4Qk3oE8GIs1TEu9CLCU7GgujboD1099hlQW/1LEZfD5G
OkuDiXGvD4LZEIxNePvZk6z61cPH+deKsOZ/mhuz1duLKLt71Oqf1LA6my73yPuz
HO8L9u5/K5Gz9My8WSngLBaiAZXtzTWSSW0FhlhWzjrX7Su7ulDDZoEA2LGZEcTL
heQoi+byM9sSS5WejduaVHIYPQMcnxIDLolIUdyp7Xlr3lBfaF+teJsu7a7MEBTk
gp2++dJ7A/jEwuHSMF1dSqsLWxjNbnU/NQ9n1o99MMr3FQPa/03Q1lcuYkhhAKz7
2Q+XybbrLw8gb70dJ1+W5azsVqN2lsVul5hr1yK0GcaxU1m+LajlHmtSDSspS3Rq
O/PGZ8OzWSEei9ArbF5yFgflJHlgX6auK7G75bTBfrWQj6Cv2BK8riI4jNxAkiFw
g0clefB0ckv3lnEP546JnaGJLmZJ2FXuYoFapSs4wKyd99WZkFN6TWXh5ibrNNuq
2lkILkAa3nOi3zQqscf85HnenDKykCPcTcgw7RuzoNtp94/+ipEstxbntbWz9Bbl
RYEWqzz40Q6U7z/wP4NY2iMb2Xf4swbWf5r0IY9VoIU51dese/bHjkzOQcavFDau
REb7gCiKMINJAHS8meHgQ7Uphlp9B8j+Ia/gdpjD9qvvBSZQcs3NYO3JeYJFyBgL
eMgEvWm/rZx/LAZdLrYbcNV05hO9DFKvSfPI199Ol9skhhaHq4JI5AUrCgR4MxlO
9Rdh1n+RGOhXWROtvCmv/cvuwfuYIU12KWmy5h0YKv3nvuYv+rHQWxwI91DN+3j+
yYHY10ETLB+u/96LzN3xztL9/9Y2UpdO+HHKBkwsdeMHc57pu7uMmGUSzR+9+L13
+uDw5EQ13w3E/O9+muRdwRwACHzD87cbtonGkZYSMHudITRxzobJdFv4n+1diZKK
lrwJLZG9G+sVKm+4gNXJbpfZWjKfuEVicOjhsu+WnLhfZnNSlqm1PvwQot3KuvLE
A+RcD2GcvGVubhEDEfukF/JIzEjI+vTc2MS44b3NRba6jA2q08qnrVoBCp9EyXzX
+BIvpMONtbECZzTQBiX26Nyb3kH0YsC3yYE2V1juTkospVzQxFd4WIMPW5CUz9oc
bq6dJwoiVCDu3N1BLtqYlMlzm77y9igfBZt/GM/2G1km71wgBH2GzhaaQLI4bXf3
2x/EHjankHP//6H0XIrsDddX+gNRNefXAPFkHWLU1dBjosDL1QxK7HbkTnn+NQXx
xR7J7NyPWXt5t/NVxO4d/k4YYbnIDc9XsfXNiJyHjjMUb/0Pkza9ckZI5XW9ar5L
8SHQ+V5xB8ey12LMMYepzvTj68OGzJvYldPUoqSSSbCc1UBI4OBzS+/QY7NPNU8O
8bcMeiDuwbBBxdljdTMawGrrZ7A5v3Xf6GkEcosReysP0N0Ty9g0/Li4avvj0Oqt
Kc6jj1GSuRj2j5LQS50gnmL94q0Ee5CdoqhHXGAGiAXuqSculvgjDgVKhvWT+mk1
b7oBWZy0CZ8/RrKPHIhlBQgfBseFjy4/XZSt4R5Vf7FpKV2hkuMpmd/XsEEB9/RZ
Q68BvQoI18tbKSQoJT6kYpM4XhFdEpiYy6YmRlLdNTZUaJvQRxW0owdUYqECrB5g
ePMzxL4IomLC0aYBF+ZKBKN9xTwGwwPU+sQlGIcVC6p6rRIA3XzXvSJNzPkIE854
dwikj41uEREuSA3TLtlBkqB9R+51gbyyi/600mHYVhOrVcBpMFII79GEt7+Ik5x9
qoRjQYheek1qfL+4kCNJ6UR62NFT/UQxJ1VuwddDEz4JroWL3LMVWvY2FmdC4lE3
zp2l4WdYFqtERWkvFyZ9YklDM7o/pxbpsi3oX9qJJi+dml5tRMRvhL6ftzqrFG7l
m8EDtrlerFFReB4bgBX1UC+N25OIE5rnU/4QW1umynr10VnNFMwYFaSOtDvxcsbQ
xOdZEDr1/pIZMRLKegMjU20dL150FkGmEsDyuLHuM9ntVCth0pknEsvXkV0rEvPp
2tELW8ja5KIwNNe2JDVlKPLN6T0jNjKMJbMZg7lU2K93B9ZGPPYW7IIrkyX2lvfS
Vj/E0WWOJ3s6AicoZqtY6wpK6LI+zzpp45yZwWobLjtty+wGrhxXPoRAggwCR5mi
PCezZbD7E0d9BfecjwnEWPR14ROZ/0j7jt+vPXTlsUtcfa5V6yin9w/OLA2GsJ1n
Q80wJy1eHNUjulzGnC+0mV7oZC6NwG7xe3yw1eZ2h2KI57H8oW9dz9i8dKmA06cq
Jt0NWpo0gMBMK6SclaU95+rhc0lZb4xcNRmNBy1sUB28Y+D0RVl6TR5rTdXC4mTo
KDFMDnDb7hNDk5gj4jwjWHdX67DNIkwz7ELhgBD7su3tNTFXhu+OR7kACCJ+CFsm
RdThb4q0UDBCh+Q2g9EkFgvJ4FrpgUIk+19u8HkyOQyvSq2qud3Br5sEaMm6O1zX
XTQi75uVmBIoJtldP97ezWukLxSJn2wHMzy+Hlx8iYQ0dw3T4MlpvsxbFe2l1q/V
cFvRFHLyrqhATqTIuA8oh0N9BGwy0A3D7PBSh5v4Maqc7HAlVJ86VQDiojB8U2Hm
QofZnM4hhQIjST07mtYMxLdLIuGTe4LTzuAkKP/G7X8tnupXmNl00aVlWO/lNnQT
JTuBn291PgfzejOaBAE/RTJ8LZG+LTVuwVQRnmCVXqz+yZSCJ0i2jUg5pOkU4ryO
c9lUPz11uSSB0HI/ULud10dJz6/3s+3qOFnNC4ArdzI2JIoYTgTws9nHCNjB9lVx
4PAI5FqLi1TiUeHVETCuyYdgbI3+3/xN/2C+MU6BREqCj+NgX19lPXEIISaGfYOg
fPtaw064Z4idayLyWEDduSTAcP9eAaogMgMTz34hznlvIgSZ6VGmfj4CZZIJpb4f
7GTZPg+5cSASo6operAzpMnh5BMF4zE78OH5bOdZjc97EM8OiBzdPcGbb9lN9zjB
eZO+D5rpJzqcR3W2r2f/eiHZWUCDNp14CZEZJ6BNVQ1eAvZHrO4HyFSz8mmqZ/Ou
zyb53XWK7OW1/ALyzCwO12a+Zh2WZOtWcZA+QvrBNHj2aciL6VzXSO5kpY3Fr4tX
WdkXSBg65uwc5kulabD7PHRa3alruicCRXi6sbWe1KC0cU1lUX+hI6J9rwLG+sY5
NoIC075SRZtmsI6swIOy1VICpi4oo4N8K/9LWnfvREWcgDh9VysAASzwb8xs7+B0
gvCWNPa90AAjSS9E/tpUpbxdWXxrhNPyVnQ4h1FXxFskCTFPba2m+3EAEcIdW2kn
1WjvXjzwnRohgoSqgzPEWlDVZVZ1/Bgx/kuT/RBbfGb4kAib1RiNYPJSnoNVfjUP
kknrkBS1YrXbtIjK/dJeln6j4NDbf5+X0k2RaKl2diMzV80nvXcWHfdUbPQdzexJ
+gZd9a3Z8kXd1I2mZEBqMewE7D6OswEHlmRBiclcRX1w0Y8NJYl99UqTp0IrmPFi
dQEQHMgssDqEzw+A8jdLBW+ecaUqkiqjuT0DuMfD7hHnm4cL3T2Y4lgA4rh63qiD
v77V25Nof+1zi9tFo5SRJ0rhdwJHX5EbfJd6P6N8CDI90fjcE7yCZ6UwHv6lKzxX
nLY0vG3nC6mA3UV8neYOVV+2QVyjC7Fv3Lg4Xx3FkCvbHlEQhHDxYe37S2mc65q1
PKNLd9vlsowRx65gUdXx5s9YLWiPPjc6zc0M71QfO6AAi44ygQD8CPl5FvlUhc3n
n6x7q+IwoWezn1MyEQCoUhVXbngSh57OOo6wMOa4TAr3VIUZFQuMgIBuumvRK01m
RFyRnz0EY5WfK8cBSA9gD6T14I0ct6MbQDAZtxChJF/BsasXmNPE/mG4FalvNSK1
wbDLkmTc0Z0Wh78I2WhwAhqsEoU3YYOUfARCYKU54qu3ugVGkcvYKnBn5kjBlKr3
E7soW43nABfVYkqWQxqZ2smK9lnM76RlFuB/kTdjo0mM7rHYb2DAqCyyksrXKZD+
+2xpOFI8bv0Vv+d346DSgUlmOvBGfzebow69DcoSTXJLOFG8tyiF+wzbT4ESsLiP
IDlN/TqkL9ybpyR1mZwufNxLG4RZLVehCd6C6mllMOiI55ehVA8SdsVlOXo79DQA
VulzfIsgXlH/9hhSJr76LeqeH20Ou5XkFmln0CgStQhFZkjLGqusF0ZHoSfYrFHA
4PFwYHL+ajhvBnb6fqNh3GB/ch7M9TRpFTKowdYqBVTjoRpr2OdKzvzTCpK2qlBb
J9YqHJR6HKXHL1+E9hcXfcSprX5UgMnSLbuJ+eDuqGev7ikRP4ZRp4ZC+EL2+F0Z
YGkPEDLcbtrWuizZCgeKp7qRFF1aEqsGe/xyJ9ITD9CudtYk218sHYJANeA+M+WY
B7veH8igJpybbkAvkesxxS9tHhSapRmrUgL8ftUm7ngSTms9I5QzrvJNvDSF2KTY
vue4GRCgr5wGcJHz2miK69HdGM9IS2JarhWYobQ1bemkuFFJWV3JAPYyvot4lQHl
2pw/BGju4LFGmPyK0H2tszBjuSNRvIkXoV2npan+nldENycMN7PsASinOnh1mgsi
Uf5R8ee7TqjT+K3UPw8qKyYH5ZaHvxfT0AeQhxVVgMedwXeRTC8PtLiSaMUuaerb
+137y9+sXzZofuXWI3z3i8UJdqCJgjR4ZeSURu2+5h2mXjVh9X/43q6wXkKkY8f+
PeOiZVPzfqXOyGuErivxsbbUUp3jKLMSoYAwunuaHEzioP7wXj3K8qoqzmVVlr7w
p0PI10RX1I/h7KHC9/ZjTtqfw7+iZ8DMXcQ79hZ2eKL4K74KAZdWlocrYfPbQmiA
hhqQOiqajMQN0WPEyYMgw0U0e2s2BUFgy6lMTazuzHd+rI9icmvKEE5Se32PNjSR
ZmF8jrmtYkrpBTR3apEMVngadGBcMzmDAnDJDu64V3qIw1rhqKg/YyzACN8D439D
g8FJMOiUeVI3OqWz+T1oHJi/A1MV/XmS+LmRxHlAz27x7osufPMuaaNbnYk4F8xt
g8RueI/G817baSNrQuU0MDw7jOAdmcyLzLVQ5UGysB/MlH04g1zn0XqX0/SUpX5R
ifYX4dKEA9kiHIvZoCxZQgLn1YxeTW2ZX1KAdQU1vIdDymL1GiIU58+f96dClzS7
hCWxGiHDQk3RPX6bgj1Ia15D9JZS+23PNAALupJ5FXB5hqbJas6Zf7iknaSmU92I
bRxwO1HOgCcK6kGAJGo+s4M099rekl+MKv7097lRK13v9/fCYDtY1xt2BRiB+SAz
CoG/P9SkvDOZm0hLi7ieSP1Vp/YovSER6cE/bFmqFjLRTE9DPvtAdQZlzU+vka2d
ThAfVAvT6IEsb85KsYJXEHWvI6MILSyW/APD4HHHB/V2xMbFD2ykNw3UTsRmF/m0
bbbrEt8n0npQzg/ljfd4mtc3dsomEWfFaWRAPfxZ4UH6slub+yPDMwq0NCYIRxXO
NW77RWvVDNRYlrfDbkipjNwaRfd9Q8hlTxqQq1WD+TTIA0me9GJ726fzlikJVoou
saqV6bYH/wXBFNn/bMOdPgthnzX5dEekEPCgCFKB7PT8AQYwUIhAB66kiXqdmXHg
/4nslsW5IPtB+Bfyt3fPMi2q/O3+0xbKbgGFMTcR3CjQUE0PSkBoFaovDhzd2yEZ
FCCrGDfKWejwUc1r1BZp/01iuK644zQ+Ug5unreA4jxXCf/JeQqYqNUCdGoN4iBi
6O7Fu8IiTb3s361Y+i5yQGmOKO7CweL7nQ6WBzxZ8uMrNL8Us9+0zjkzizV3U+w6
5vZXZfUlwIUcVo5TveWDs005evnIUia/MOahuu0H6d6oZ/NEas3ym7PERNBeT2Hf
OGilJ61dpbCIRfJeNNEJyIQXZU5+IrdYML8tpXvpXplS3LgCIV2HYDc7nR6UxfHv
nm15j3jg4oAJnfsp0H/gr/5d8wLdk5KrPCCmWzrNsQ0NaQeA4deVCVJ6qpk9YxAv
Y/C79OQjTHznfizkJnfcPr4T0QlHVbJsBzIyPbcUKKu+yAKluWbhEqjOlEuhb7aO
Y2nEPfL93fkVLj9G54M0SzuwcdCCF/yQOlLLdff6qw4SYi5gCbvysEUQ54ykE7Ej
fCOqy1b9kdQwzj0Mb6RLpkpo2vAK/NjKHRKJasmI6M/drZql4I4tfOWxluUdt5GF
itE4TfKph1dC/ADPKx48BfhF1RJ3WckHCj887YK5zZlUsion46LoUObzAI59L4yX
SC9J4hBFmlqTAhc4Le8AseGliYkGgW8Pp3To4sCQ95hchlIvweZaahvZj6Z0D6B+
7vw9EtXqF918PzKtbEjHl0NgvSr+SQLR9CB0UE9KSoU7sf0Sl0uDWO/HwyhP9AsW
TawkPJoMIWZtvL7QqPF+a9TctIXpN15vXAG/P5TZSwVH14rgJbbBqN8XbqQUr8hK
hRecfZ3kb09InnKfFx73DGQ4h6iLXkIS68EJ5cgYaGQxwLg4ud7sbHprQsIucYg0
wkYZiEqvNTJtXfaNjmyU8a6oo3gc9gmS/oIq3EDkr9BeMA4xx9hHop7U39XngOmq
CpaOo6YwI9TDbyEvnNCXT+qN35bbcO4zsJBpLBOVJkWOTpcwG6XM6pHK8Cw5vpq8
N7yyEb0vRn/+19Yja2b5n8lVK+6SChLtfOHsJwDlVanQb3GgVMwMoMvyCGYlR1uV
Kmxwm5XHMbnNZS5wuQgIO7uCTESCIRcqnS6V5UWeRbzMXJqt/KN2eoo6pR7eXZft
c2J2pRhkXLxyP/AUPgEyyePaEOMnufdeFrWz1BrYF1X0bkOShotaW7PpxYNCfoUs
ivRdUau26GZPF2FTvy2VI8CRzmNC/Jhu33Rp/LJ3rceXq3sjRx3xi+AlUtAGoSrs
eTyInW4yhsnTjdqET9FW+ZkhYL18PpgXRGuVsZB/JzQKVQW07Pk3UjxqWR4fUsdF
sbxe3IMJozKFmO/B9iuscCcnqCmLqnf0m7JiHzy6wEAXbPWv9WRkMWq+qkKPsgvY
CIucD3PwRcRnLQxqJnaUFGbgfS4M0wBHDRfdyJ1mbWPr6E7Q86G3ixTrFSJhnJcr
9v3JUp8XYWbb56PdymucHH66ZPcgpihrRp6Yufc5Wz7MAsiKHCX3OgfyJbTyYT7R
uZR4DJSwe/FefJ+dHU/Zp1lnisSuSJVH2vIZffyVLX+4kCX23hD28EMs3eZUSQqm
h3eM8Jz14UUl3zv2JGAxi0DQFgtNCF6gUTeEYnkFSxhZAHz4ae1nh1LWzp+pbKy3
+rA0Y4t3EDIyXarApcozeU8nqUWNcRnZ4hYyiWNURNBkJE4d/demeRbqnQVgd2pY
F1x4qk90JPkOGG4AhJBmcpFtrD9IAjvR1zEnWPCzFNJURm2+S8zCp6HEKzmBFLAy
0yOXxyxd/d6uqJJOOY236G5CRsSugokYgBnF7+jNsTYwvW13xWyex8ILR7H0J/HF
mNvUS0/we7Ip8D4F0OiKKCC013Qt/Zd1zSKEsiwlSdOYCq4fN7adKKRRZrlB3/6A
8ZMEgt3p1o039GqaXJ3yujA/xPJMReuD6aZ7R7MwD63psLFwEcqzvqIRlfeJ639s
+akDKGpakjoxoMMghCOxm2BJ6PGMKu56bYyOimqPF4XpSh/C7n25gELp+D6CYNCg
cSdSLA3DL/6ojTVewopnr+dJA4c/m2e9qvfijqojDudHM+L6mPTQjrGMa67qVSy1
50FZjWHBqYKEfLOhjhsRrVE5UUG2HKYzTqeauXAWuV3j7Mp+Or63hYznwvy9YOSd
RFFowMbDDj13uXHxsFyRU5VpTdKE34atUuLs3kfHTD6qle4fzoRs6U+LhDUdACpO
CHz4vV1d5oTu2XPW4QweccBGK4FdVi91iYw/CzJN1U/pStiKAdsxJQyS3m0rFiQU
EpgTSP+rYsb63KmFPm6DKp9qmVBbApQToyKIfRy9FgoXXuC7bRWD18FZrDzZzcFD
xdpsSe+EHVNV2kaYdl80Z2SV06NzNDBKFcn1rYxwB5rtck7lzXJj46vDk2yHgJRI
pqS6aubd0YFZRXUqnsSnmz6suRWeDsbKLo1jLxnojRwLcKdByiJ6heYDvKvMy03j
R8xqLRh0XwqJyq8QkF0zGrxU8L+ntvs494rJ2nT3fqQR0GOqKqmbAhS/96VPgmHV
bWIv7pdErNT6yPpS0YBdZ/rW8d4c4stedHFhzMyuu5PXd0iSSoDL3NbQ+2SEr76G
Bu1JvlNPUOpHeZrWJZsKdpZ0l4iR958FJYHAemWkklX651HcjBuyubQnXopOyl2Z
/nVA8283SzB1jyhkLovMfG5VxTSIVmKbMHX7bP7I5l5Eu40Vmxo1EdaXS8X+vU/f
xe+a5dTiBXJSR+PvmctW6LmfzhDcZmCeruGnf1gib6G6wb1Cp1woPVLRNMPeiOBD
FwDkcjxJP7GYwRHrjZB+QJGJqvTAG75aIqNtAzUnI/ZOZjsSahiYiDQwb/qHKuoD
IwNRxBZiNCeCluCJUMZ8m8obNtp7ATkORLoShAX4bedjMr372h77Wjfz48DuJ/VZ
QFcpRRiYP/o+HTkc1ErdtZ4ibdrKlNSVyu2co1HmnFtjNvHj/GqTAo5xygCmpPCm
QtMGAKtRFjoDzlyjuAzBh8h06DfSt9DkH+Zh8vZd+zxm9mkoz0iUBa8XxoiKTa2V
58LpsKTTXRDTNx334QjIcmh0g6+Z3yenA0P8nVCKQU8CrLqa1jV7RLPlRGY2SDXy
6LvwOXEdtUEhxBKqUYsJKDOe0ootHDGJw+/f9flELf53Uww0lmKHSO013hBoMM+9
5cmPRNOOCsnawV9ds5BTiZc3kOymrD+r7VGdVhHdFyCvPUpfnq56tmWQj9YPeYqp
3OWQ7Up+nQ0V2MHlUG5mEQYePOHdDoLHXHeoKpExhRIfd1L2Vl66z8d7hjftO8DQ
ZEkKWs2V0MAXh57sqPgSORxpML1NZSTk4TMIETtih4KNLd7U3rQqRlfftP1IBKvI
HqIsOhM/neOelDJ2y8wg99pX69M6ZlMkIih3oD583xTCGp0JEBueaBJUCHs+SnN1
YVlV0JFv+st06EwZwMGIQdzRGOKyaot+hd6RmFLmLVhhjBTOLEaqZDpAeqK5nJsa
WhlVF/fdQbOjcjZOSyf4Vrl80PHE/EVA2BRW/VudOcXQqvpaybn0V4sHOgl6HNwT
IurFrDWNIf2//ZCP/T/jDbKvlk6HqRTXeEz6P0xJeoWe67PQT3vy+oddSwZzd3no
XTwzeP7cbGUPG5rtF+uef/mp5SBl+414kcHtAz8BO4ZN3eYqmwxYA1wwLCpodj2h
WkdMs8buW7cMo1d8sVxm0mRzUE5Q60f5yfPzmjc04CsHzk1e9x/jkwJz4sju1+lT
bYO2CPWI7PLhSmExtETYDb3AAEEtoQf1HJAF/opuIhsgl/rGpmZyt/LbIUNDmj7a
aIXK7M4XijbPtmHfvlcqEINGPGTNl8/JKHXHE/lfzwy6XhZzPbLJfZQSBg/Yr3qI
FMQMsPkpR2uOIGwX9PSCQIzbIGJi8jkqI++FTQxf+jd0FwgeRDqLQoHXzUfmyIyM
oLMsM6xjrLR6eouqLdPrFK0mVsDopuu0yczEX1mh3TkSCm9/O1SBXhZyGfYOZ2hr
78c9n7tT9YYrKLo7bH8wYtAziB6zXGB50kh43CHTpFJDN6hvsvqYh6Fm551fphsl
wdv3wIv8Q9Up5JJnuAp/JR53eDOQgmDUJU1eYjHvmcoc4l192CgOM1CViqPitqGo
ylIvRJnFLEVwXmU1tj7w19/LFpVpWsGpjaKma/ygVqhrhluxw5t/EvQJi51szgIM
mlIvbhK5Ebw/4pxUFmh5+HNEwuUDTR0ut9HKdzbeZUtlrQPg4VrMlTmAouyt3Ixy
YiEiYyBPhH3JM6TvFzGc65I48Ityru5MC8iq7gsTl1t3HpDxmoaCIbFG+2Z84B2x
6dAL+Bzfrbyv514YRfIa2YElmIo3+grOUrSkAfWM58SBI+C+DZ1xS8tghn3DFdDn
BFvsvWbhv48sdWj5bii8/eGN7UGS7psOqDOAm25sLy7/HPMF9cSrh0Zksn6ctGUM
wZ+Pzq7v5Hx+cI293ld7uTmjQbcUJW3u6vRd4SjfDnHG9v0fN4DQvV4XRDqFxo3W
nfdfCUyTBCcYEff4C2NPiIj/9BSpOh7WaFZuVHRig6ebHLV6y0h8/MKLFstrg+20
1f2/dQHUEDX9tIt6DcsFKND8surRBgaEbLtWOZ1NpNiCAaj5chMD0IgXr3q8TLoG
AZhSFH5i/uIFX/W5zI7nPwDHdwsQPdo1W89+lrejGJFWscrbKf/17/hC7eCv/QsS
t2SllGtfmau7h5ZNUVbFiYkomLAEmpv7ZQlSrzAKow20wkT59l2FjA5UgMd73Msn
lcC8HYzgOf7duEnMpBbdqT8C2XZlwh4FRKWMIcMuQUfTbnKdI5Mlk1F/LlauM24+
bNlUfVd4snLAeoyYB19/drdPEsuYEMppBdHo0lxSvoL4zofAkL+LmoCM1Yrk1MLs
UU1FHjl5jKMmBgkbydcKdyOVKjGtknTlvCAZoWfMXnC/cBlaDgvhKs4hUdenM+OZ
TVAYQ1kSxwXcDDSBCW44WcU2uj92g5NMyiilSRUJnCs14+5bGkf6nwjIKhyigjhU
7o5lhSmx2cYbgPnsRDgiRHuzWOkZTIKBhB6QzvgIYy0wGO82Ne1lJCISFuS7+MSz
itkwbSwkdwyFdkp6E3zj1sn7oBskXcjy1ldOz/1rLL2iMogt6WuD49uV2cspVSos
d4Z81aRM7v+wEEqppPmILyFeF6B20ARDJg7+GIHYracDobjk1AEWnaUK/sOiFT6Z
30G9/n/f4AilzrC7i3QQyScUmbOyV3Mt+MGMjycBTw9gxIIEDUkxqEjLj6Lnzy5v
sUt9nF8r8caYK69KoGJyy8mKdq+wCybVnsbekjhhk7T5BZYPO06KIzJPO+O0/gL2
XC7wHtFxb6fgsMZbdy2yhY4XFwMzVWXcvR82NJ3B+9GM3Ix/kVwDOtRdHgC6oT+R
U/45Uk2iHfCclii9uGXYF5VuBJY4kEL6uiHsKe/HedwRbDDSUwHUJVDGiUs2URmO
7mNOYqn94LJ/3QtXJYrOl6o/SPX5zChDafFAbtiHcdeH4vfZ0ygGz/pMEIEVv4Ys
7zv1J8EMhPMvSt1MuEfyCIFnI1JGvUGRSUMBAYOAwBG8SCnSPHXQz3jAMPJxs6US
raRqDmojuVZeOowjlAPl+86jYGKiPWWiZ9Eiz3kupNw3cYpuBfWhr8nmWG670DSJ
aHVgEBq+UW1sfCZbb5pAP76M+/QflMO+PuQRVIM//8Ko7AUhRCjQO2OTNXGqKvxp
aTf+BZ9fq+s+Wl4WwnMBT58DlKPm+BrCDARcFvObl0Vd9MI5W+APOozAqIZ6JBXw
uQ14ZthJ76OwXL9OtefRBBLW9YtW5PkFvwdoK1H0kwr72pbuNT5vwulxPN9lBFpL
OLBHvE1yIcUyPXCjtl99uGBKHQc1LOvUbu6aU38v952INBTh3HNzTvqgJ3UYfdOw
C9veRy50qlmRwlH6FzttVPOWYH2hjVrp1RivE5JVKgUMsu/mC2N0uHy38QuI0TLL
rjX91T2TpLJbiH/VSWVKfJekTs6lnHv7w3TWCWim7rNYEM+j8FofNBOx8gEB59zr
Geg4/dEZT94+zLjqHq31dNeicT3yZ9On+bTp0UbIZtP4lbMxvcNj8+I6KjgyUokC
G834vqV3+UVeIC0/Y9vEuAFor1GmFOSNDGxx7lFgo2svJEPPi3WjeivKlbNSM/fa
M19d5QzMxlBQ0kgkJKzTZTLMBnroVw9Dz3UkBgooyO80YgG+gIRRoDU0LxqcWTNt
lZfgYT2ZQ65Oe29tZNf+n/1YM5sT7bTIcwSrxuMMd3OiBY7h11NNoN1I3NV4zUTC
LjlcFTtj6B2qUB2CG7ra0rOo5484oXRzX5Uet8SYw5cghopFUeJB6SdkNWA41yCR
`protect end_protected