`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7184 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl7TOuMe4xzV7rdHsSWg325trfZrlt/zHq38tHZh/un7R
mH4nP19Gt/yOeSNiUZR8ZQpgPyrYjaYNVRz/IkqB5EjSEF4wxkXLOKUtPEHfKCEj
BNgB/AKtQboRp/AVj/INkjBFLlALqLBTUmwsqId202ZkKmFRMUhI+H4TZkwTJbsl
zvsNHL+LyKDQB5fq/6E19EUCAcDs4cGjUzpuoIjAbGUOvLJfecAstSBagNdaaGxw
pGrlvO1Orm/zyod35ohx/WFXQKtn6jxuNPzGAaI/HMf3Pp3BQ+CqYqoIRINBQm6p
/xXRSwWOIJluFgqKyZI59qUkWZ/9Wm+4uEs+akOmgslOEjtYh0l78S9UCCdxRQd4
w/o4lnDKMHmvDLjrf2WafbXX2Kw1VD2TaXGDKc9CcHko24isNEFD19W28dlNG34Z
q9mVuZSzBwsRH6jctVN3Bd5PMv/LKuCer0OK1PfYak2pChOW8s2Mw3U2LuXnZDdS
fJmp4ZI6YOOmWKjXSOOXjF7s2KCOlIg/n3YpnseF8m3aLUcKrJABkH8YHrx429k/
4uNWd+McYQCXfJwNLY8WM61JfQjLZ1kYJaJIiXVcY79ABMyqwCCIOJvDF9oHPIHE
dokVVFut5RLNNzE5DNPGqS0RWhuxIukI1b6Bqni2c3oe+ILOSsbPkRyz4rBJIIzC
2r41CTP0SQCy1i6+rHb/g2CXeHXmdO5kVsOM/nJ6JZxJEAXiW2Hb0csgRC3Hy9v5
BLVGZMLWZV/AcWZN2cwx3Ul1UHkOvnB3aHGzZikruWfrES9ip4ZafevNThEQH72V
wBb77G8fbpdZeD5pMPkmkq1eT9COI3vSpAiE/dyVIHw/6ErYuw5OGxmjI831XVla
fypr3/6ur0sGzMV2asEeFSj9yB5ZkKC0A7htLSVjC+GZBthPZTxx8l4r+iFf7/z/
Z/LproAU+gt0AD7NKY3bEHHW1ZDsn3NJgwAr4yR1mUD2fGI5I2JgddGPnSUeIjiB
iBW2dXtHdyYwsvhacLVgKnLaGbjGyRQFinmIumcGDG6phIl9dL3NEVxWCUo5khFa
6c6RUSLDfpgWhIbsBfPHPlJiJUmvvt3Uyt12PTwwA8/cVi/tmrTBjBZ9exYHw9/o
wtHfa721nFiS2V6N2BX1XV6Fu3B+9E7jnfkZpJi67FffPkBwCImxh8pFqrXdoC35
Y+UgkDybW3XIYQP+KSSR4KfXpQ/JSQcAPnzbfIkSke77TGVOqkceT3bqge5bK3X3
Wv02pG2y4zj60e5Uy3YokFQrhqohIFqwKP3wjNYTmiCnahD4Ku5dl+uB+2i0zjZR
29mA/lhUChNIe4dFWqrXRY94+yhw1aZHIxpC60K5iSUt8BjNwymJaLTljAaO6asl
i1q50e50AQ/AZ8u5NMJrJDY0KYA5XK6uOTXjPK15N2qKSwdMG17CUAB5E5aPwa2x
NVfM903v/lyJz65yPeg/qOrSDnSo0W/ZdMms8+RShlRweQfKdtKi1Dbd4yuXmFBj
W6xBULh/cLqA+PWDI6XkHAIc2bcocR0lVb6deweslxq5RiQhHfMw4vqPp+laPiYD
B9GTs7G0t6d77zBnZuoAa0eOQH9mhk1Rcx6qMOFFZkNRbZETlKGgS+DWdCLl8uwO
627puzrFZh7LhBubnGfv70e+5xjK7szM3xMtHULGPBpXJom93+p7H5PkK1Oa+/QY
+w8y3xjeWj9FU4m37fN6QZXv6W8sZMOHOsz2SfgPqj8h+GHMFx1ghbC+1hd7pSia
b+ONOXiJ0vM2IeHWMw08OKuoPX/KqHK5YFhRAFs0bnInFCNl4PLZttTpUI/NjcJY
apR40szmPCeFXAPXAfyMbYc5mTptQZE0MYA4HgWmMIAcErwAUX2oPXRs8n65VRZV
AYs73qT2S1jIYLkWtNyy9nga9gfhNLoZw2OzOMdf3ccmsLkAHmQ53Ihq5Eg6UbCi
RZRQO31tbIoqqpliamiS0QQU8Q1ATxZUqhkRScg0ZpOf8GJoUDbcEtr9LvQieI4u
ukzSHTRhPT7yaMR9y+b7X8JPdXvdqW4Y5rtxdxzxi8oRcknqxT3hdz+TWkkTQFDa
7tcO86E1u0XngukHSJb2S0nVuDbIsQWBpvwR1OZQihd46oLa83VXGKjYJQ1GcA7P
ycEPMmrr1O63FnweNNw5a+/C02jfzk32B653UstHGEBWytCn+XhweKuYSk2DPhQB
yzZgUtpnUgLxP7PgWKAYcBX7i+HvWsd3D7aMSzNpTttEKpp90N7lqjseTSogxCVE
DBe1C5s41+ZBPGsAtTy3xc/7i/YoGio+7ZBdOc/3zB8BFTbvPU2u1CKBWoKcjxcu
MiO1EzLMoQAZkU7B+34GnRo+BB4psUmTuVKpCovQVOwG8jKeSHGmwSRVnJ9LczO9
GPb5p69yJ5NhcoUIFRYfVaxG61svPDar2qcW16dowqnpJJtYrAgUjgJKm8AfTk9s
n3FtxSrxIYhvi8GmaioI+V45SsM/ETHNTQbh7c60hNFqjM4jGvAtlk6tq9BQQAEn
/DU3TfzaBe4AWy8p/uFO67n5CUkCpK5H5YRHMI0z6iF2XRF1da0yb++WZB/hNh/V
BS9Dkh8WkB0Hf7BfjZAga/gWXsWTpVZpxtli8syCObFrz9y7H+HsTVYahp9vQFaG
06upO+qMP/NIVfRO+jzFmrWG7U4w4wsdzrlm+7VJk4LuwAmsiLyOYrNJ03/kQnPz
TXQiC1IU9lStgmtMESUaf+x/DZ0zWfewBFLfS/67RVEqQ09tPg1BZPa+MCU/LuGZ
QofS/iC41X7b9yL3S7SkkFcgwE8c9a0irf/Aa8kasfLBlyOUh74ZVhdz03Qmt+Rv
FtQzPtpu6tpiASFZna4G0pqM2Ak4E3YILozhSEcApG8qaQKkUw42mNqDxbkVTSiK
rqkZvwdrHeyGzPeAt/OSty/ZMxqTqSnJtK7NTTv5wDD+2Y1KiuPAbIreQCLtZXsP
o4hU6DdSnfgxQIgVB4/moqWjbCmH4TjfhE30Jy8DatZSlKcxTDvY16bKDrt2D9vr
agT8UmCypX7O+9smBb4t/H5LrL6epPyEyaLbcrEgIFWKhILBpOcFxOQzrkYY2Ua7
8Y0S0NWJVx+UjhDbTpXpZYp5O1hG5x6ZZq+EIii4yPsoXeDLOcdFhOmlyXHNYONQ
uxu6HDqdUqXEEwMs+vVu18d7/qk9OuAyHqXxSFmL/+n9ExTWppKsW5tQLiVQjumA
/7iL6coP1319FGB1vmRUmIWiQJt+aR5tFW6pfi0awAXDCkKCcz1P3gbVOM/yOJai
e4LkEqq09heVWKeBeNMCKm3nVhe3D3e7o83tQsXf/s+AmM4JGohHMyehYewIQi7l
1q9O6Y+ndZWro0Dq5ksaNQ1CluPsad4B42iP8X9uohIIvODU453czprq/KNsGI1O
N34iz1RFNloVa4FJX2AVGSHqsGOswpvULYagK44izSWn0+/Bp6RSYY/6MZnknxfu
vOUva/E8DDbRl52qDCQ4dLjeQQc5sFcoP0Jq0/Fa7Wr8uNu0xPX7+XUmxhITDXAB
O79M9qYaBL0Us8f09Obft6TXmf6QNorpLGGadUgjzSh/x2lqRGU5qUebwhaGUCdD
03RyhgiUrnKnRNZ6K98Zn23ruzlAms9zFNOOUxHuEW2hCXXvHkbiBtBBw7+XjpEL
EgIwQIbVlUJ63JATpsU+2/+PKUys2zKycONybMxnY4ezdf8GzDQp0u63Ab1aQD+4
kx6LFqdDIwikneXbz976hfXlPVgjr26zpOkEUEWanOzCHYSK6QSAPxBlOGxbW2AK
suJcCWlOpL1+goOHbRcn0jGowa349AypbvNkTtxdzGMBsj4q9PJzbpu4do8U4GMP
+LP5eNbSWh6fK4oxxWjhwLCy/pgfxBRLHs6yolNn4HIitbBVznUZF8R9TBmkyjeS
Vr44Y1wtpIfYYq39e83aNBWwdt+VgOWo9zngM0d0bymBq56NKlBlKSmvzbTCQpT1
wRKCHhvGTQdCCkx6H/Ltr0lVx1tsyBuP0yxQagWjzLzWayeibuAJbEckjTAlWz5a
RyKVvslT9/J6N2Aalv+LsVG0HxoyeHlQDJFO51+1HNsMmss4lq5Lkqc/X0UXF+o1
TQ8qW7meKiR1jUiNHlmtobFe7bB8kb7cJQeD4U3w226AsGkA+YGoJMfud/WscvYP
idJVyfuMbgvwJQK/TG7Y3vmBhcP+BDvnaA7Jv/StZtEmZC4atJiDXUnVEg1TJrQ+
uvoNxIWsktCL9Kb6J8X3X+zgvDaZEZhXtfYh02eFnWLIY19Fxo2gX9vl5/aMmJ+C
8Hj6GW/2Q5xDB9lb/gRQBw/H0dKLLTvp6IDXIniJDquhi88PUesekoK8KMoflWlk
t4mawPA5PrDkYTKS2DoiTPp1HlepxOPtrrxH+6kpYV14PDTk7qUzHFOpl8VHCBfg
LTQl02POJ97tWGiGXsC1uyZjS8Q3HGwv9UWnM2GVRTz93oTTgRAXlcA6gYARiaJu
CfPnbuSflXczfImC+SP5DYdjngw69GiWmWgM9lmxkZ9vzDSY59KZ0DPBQgLD60TO
7ckJ2UgJlRiT21ZedE4WSPvOfIRpXzHjYJ0JV6PeHkVbxDkIl1xR1FltLdjVZ8Cy
TaOkjsw/3YSM1LtWzJzcsUfBnpMdW3r0NoxiZ1IvnNvEv4DiqppX5GpEpu/1KePY
Bh0vQQXWDDTydT8XrE2xCbexHQ/EXzs4+JGv4UTEuA3/s7UE8uz8PpCZQi0m3YHq
op8ftG21OqeBckbcrkIFdAnVb79XxAMys/jEu+N4g4G5BIVK6DRp6oRAuE4vVLD1
TDY/EnNhs53ihu8rpULnbi2kXyeCggZe9EpvgEuk3mQm+3DaolNLHP3jSwfRDdFF
S1gyNBtGHCUiRQID3z71GEThMZpyGCR2tTZlwmkHhFXAfDddpx8l1rDlP5/flS5b
Ux+l+QKPyMkunMsT5ZD/hYi2iJM+5TwYUQDGEJ/aMCjXAIWAqojQh+98YLpCixEV
IBL++/CNERypaId1VGXIycbsjBzUtQRaNdQm50a5eJ+Oawvx7SpA7XQVIKh8+6GQ
TpeU6i+afjxCl2GwmZAHPoDuPDtWLIIsnj1j3QX68DE4OiAP96qrxgbIbvSMS4Dg
fnlKgT3WbvnEYrpCyDg2NSx61G3c2/hDICiUr1d1DM0n8h7CeuKv9R1DrPbE9jbe
+mesiG/5AzrhgtmKciW8wC0g5U4YDB6XxYkv9PVaMX/dOePKIbk7vDXNFdG/fJWH
QG6qLVMi7iSuixyQ7wVhj+sSMGHgnINLMR0gQ12qM0Vsal1/cGHQ8x2DGhi160Vg
lOGchC/5x6ApL4TlLdtMwQstm9q1adNaHQqVKxAp3Ld54zsNEnsz42vIE4I4FXjy
13OP/soZ+pNLrmNOzvR8WKJfvnSOAAe3RJj1QlQifViV+PAhACWKfvRP6tu3aYTU
0UxJakufAaZH6BH9FThzPkkLqm+u624LIqNN/tmwA7o1CjnsR8paA/st0m5Et/qi
PDw3u/lGvdvRDc98KwBayPkMpB0VN1xZ9ZT72ftNVTbOxzjPmI8rlnw8kK5UVMD3
6LrBIndQSU8cC6wEDR8z9+6XfBXwN9xoVj6gfbzz8mkauh2qVWlppO+zq9QBMnyC
uy//GI5YUiG9LpPt67uGsf/P8lCFG5ZfoXxuf9GE/UHybrGBVVHocKL7JAanh/6v
oGddktVQetkBytYLXEcnE0bTIHB+hdaDWykuRxM0pa70VG2JbXbK/RG6yV4EH0JF
EV3rJSIiOxwoRd9N20jnLNuXNjr1Je4cYlUEln7uhbOWGFoHLRHm7p+LSB9/ZYlL
qPcMbc0v0GZEc1LP7Jo3gxb/hJpD8W3WXlGioK8yhgwxSJwlolFIdQKfB+SwtzBA
SQUaW+AmVGp+WuxQzheJJPWkxlfJRcThwMXTQGVBZR/WF1zFCmiuF8aHMho/42zP
FUNN2S1hVyMKWv6a9mIlfZ6RtO1ths38Ryz2s3OOwvXqsGuKDA4BSlCn6TmvqupP
OIVz0Ij/zg9mTRGdt9NEZNVRik42mXPa4gU1YSW+10NWotOYK7BmxJdYCYJh4iHa
bJ64WiZ3PGgDT5G02oxTLnIHY32lBmmTVyMcp63zOnL8fGQkG2RzO8vT6zRtXCdc
Ke0JoxFwuFJcXTlv7X4uZK+ZwpOgDAijpYfYFjS7rX6fvxSg1Fz971mfT1hfx75b
s9Et3c/XSi18fqI2zc4w6cBWmOMNCfHe9TCxHe8+jyF84YUH2EQYAqPig2UuMuT4
xlrrPqfDbR8TYa7QJ/mxwam0DwDgOY2xtmQWTbn9D7Sr16T4b6Gae0o7u7ZQYN57
g1AHCcnV2OCoN0SyjEOXmrwnFZ1QdRw7w/eYJ0uxSslAfTD4nbydsBf5x0xfxlc/
Be1rUNZKo7476pZWbkD2hg7tTZxzQBDa89uXIcr+S8AMd5f6Jy1/aS0FlBjGc2B3
DeN2V2O79W+6BUR6yOAZlcRH8vogJxdCnn4o0WsNWzmsI6Uehy5AOHULmlEsY51z
yeKZ0bCx9Um+3mdpGWzoiGwhjyxu5dZDBoYM6BBaxqewAa5Si6vbeFp/pNwkDHyb
ZWqFwR3+rQbGEeEIDXudgE9fEJVe+1QJll3NGnXMRt9p0tojVb3ztGoNn9aGKPNT
QgpndIzXiLQr+fBxj9+APwLyIcZKTxQ6iaHReYo++PUr1fcPrbNQS3we/Fn+wMTF
8i2c4uZTJpeVNI5TnSRjUxpquRi0rQGmaVpGOrBysHgIGlasaVliM+RQEIFbc/Qv
E0IkGxfzY57NyBT3UUSfSfqLxcDXwxH/C+0OnDXq0IVogbII33jdfCFFVYFtIEqO
eWR0jcOc1nLNPp9j+lY040Hfj1x9/6jB36UJI3XxD22Ywd6SgzmXUhnW6Ith2nRS
ISWVW+WQyG7BWIELCn8jG/Ae0as7XP18pa7E87BXgFIMe6Yw44Jo+vjbFvEX3nh9
3r4YhEv1nYOiaCsagc8SwQK5J1LcZIObKkgD3gdtKIKfNBpQb9OKB0Hk5p6Jigb6
6GI+VwOTt5XbU2XmI37v28TS6NmVoXnfC/sn0ColUbzWdoaOOPuOJbt3NVgtBbdp
aD0icSDKGpzR+C6BBIHDQtmRSWIhtX/rae+P85H3U9XlhFkod7GrQw8kjo0azB3z
4M0/mhkNi2VoeRsNbqnTVwXZRZRJamzDQfaCzNu9n9w2A1NIyGzbqMH8GGffd2q1
EWvhl3j/JeXxw288kYq/2ZO4yI9aML5tHV3TaxegkRdKtPSYhAdL8lb6TK1CMloX
nrIcozsWAxZ0SpA7vxHnLK5hiPbYwdQnQnomoKGDBrW0bErd2BzmV9MGoqEBVrtN
LNVyNJdQU2fjWjCUlQoDzAToDlqFNKSbNagfoHFtLSom6Ks7SZWlihid+J9OcpEb
8rBTwec4FDMzUsH/8HrqKTZN84kzTWPEwnv2fSS5pKV3ndhMWCZvMjpDGKoCLyOL
TeYY3hja+NsdWk5PSVUAJhHp/5SB84HqcOF7nXd3LtloCYMmaqlW6l5jBt7Y+ZXK
0W0LrgYOgJEcTcSk62sh+FBwsBXUOMvhCiOqlekzVgrJRtB/TeXsDHaMHmRujgyi
wcdzzVKh1bg5uZoLYNrK8q2e+16hnwfmIJJlfdJqXVxbCfM9is8KdkM82iWy3GNN
wxOmBir1e6JNTo78HDMVFy0EKOtwcxxPweD/+wBFAFW8ElJ2wY/XFzzlMS3aKEER
rw0BkGNxL2PDSvci9YBKDcyb0N2WdbvbQJxTO5HaOFRZvMZ28Kt/VHY/mESHn/y4
oL6oA+f9DSPurjjsedI+hS4G4rOUN8GATv3YlXp5rpc8ZtQobRLK46LqgO7li+5F
wlj8yXFlc79oDmB83O9OJLbPISppYZeIC/oqmOSnYiGZ6Du09LueEbsBZFFV+YGV
BDg68Zcb+4dsTkiYP1PcK4goXtFhvvl/Rltw49eLQiuihJCvrQMtN1bpIkn/7qFb
NeGblgpm6ndVyii/ePNLtfpc5eJy1SyvP3HmohCxpDqLLHmL3oFjpLMEaA2C7Upg
D7KGl6oMvuPK8b3qXLZXWyfhFouGCOgV5NtIFmbPNMPpZu0vT9MoUbBcA9EeN2gV
+S5mrSYBHSimAkfxIPhRDtOkTFIJ63Z75hMOKpbBrMdCC8jYUoyC5PbZNlXMjgfQ
KvIP9mWR2F0P7itnN4tV3GN08hHorlVLLDjrfegQ4x/5wyfLKVg9z8wLHYjpYc6P
yIrKfqPsAsXVawx6FZiUmbXIoWBpM68cy+Iei08xMx0SFlYaqfu5q0KL0TSI4Cwd
FbKn/NraPtJbqzJKBnZ7EumiHv98inWmzLjytGHBObTLep8z+dHe8Os0LMUWl/Sh
nccqk+HAbAwUDeyKMq2M2RGWftrw8DTWL+UM1zySwcZ9e/vTWyXeY+MLmQqonPHQ
OqfuJZ6uUH9q+adHPtHyCQDmNYDuIHcJUfQeDckJfytKIfGNb+LsjtSppnAoA2Pa
qNWvjf6xEJ3dmzcM9cu3NT2lxTaXLUnqsLPp1e7ezWeM4vRKkjkicVjqfYXPD94y
6gZ5S4hPe1noFmyk41M0zTa+gx7vXYql8Ofjr5Zez3jUf7YskxkF2AvBT2KDj5G1
QeIH44VA/ZRv4/zFH8CNHioFcw7wo8xZD1JrFJvJgwWenLFWgE9xdQxI/DDNiERG
6pUNsIo/zKJIfOzMNua2xyf6l+ywJI+OQhaVp0ovrR+aO8VSYEGr9KyXzotGy9B2
IiPBbIGfpEoTauJJNoYS+tc4ADq2HKfNfMk07/y2Fq/c7D9bjZbryKbaaq3qzYhS
HE+9+S7f42a3dgZU7X3oP02av4dZ88tL6xdEgHkldpDkP4RJiTWaRr4WLqQz5SZQ
wR5Jc/Psohgg1UxcV0itARst97UAmNoGO3kGzFqoencWDOfaGXL0DObzLt5ZPvuz
Dl6tfnxIC521jQuxCafksON5dsMnBq627+N5H73j0C8YhKJOEWvldshrZzNf9Oxf
E4kmXiDX+wbPZkHTxizSBMNc7oX7p4W2sN49Cc/yAi9nZ+Q+cdO+mZP4D9ZzEgFR
ESw1K0n9PcWrAeGWTJXHxoc1k2ivhVrMkVPjN5ub7cjq5Z0UfFtxUGHDpmwoPKVm
SiHuEAu8Jk0/uQP+DpaDNPmuVN4upWmqvHCnrOWp8+kNbHOYSd2C3pzg/jyCi/4P
8nlx5W9Dur6zeVPITST1BSFx7a9sO9x39J+mPntlI5Hopta0tA7FulrZyUeNhWbE
Vl2xV3DWdBICag27ICl4SVHWToAXWLLw+bCiAAXPoeuTdigvMS6ozpATwMlsd5TD
2pl4hld/qMVGEHdnb/FYi36pM4zRlw7qqz+2KBBV9HE=
`protect end_protected