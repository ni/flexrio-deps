`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1648 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTDQnjNx0SkebF2ITzJhbjVKI0ZuOl6Z1TYui9qBgZYOo
Sj1n0oyKqufY8qMD+QgPAgdKOZDwRpm25uNQS60ybw9KvGYyzWh2Bhs8F3D/7kW7
4qYVGwgogwBWw4aFnMkeA5tmGC2rOJ41IY0XBlWahcB9lkFvlgqcBolYnHQ+5M6Q
go1VOgudjqKToC+gkogm+bMeGKFLBiP9beyBojPL9j05R2mU0fOCQ7kkL/TtPTKk
3o9IzchQ4zchb4GKP2MPqXdj6wBq6J5X3eCA4QWk59uR/z0Yw8CxQPKaq7i09Ncy
NS6Eewk6hhXTeGPDtVIIEjbxgkoKf2XPhA1jeFOmbv0VKNwB1yI6YR7EORWK0OIY
LV0Hy4rMc1W2vXLlqdiI93Q8ipA+X62G+nazcn8Xaaf9+dwO/T1HMXY7FUdpAKva
P7q/B6aItbjyZJGurbNNld/R+KivsU+kA1Tj4MnjaUT+lG7UnVM2ifzuQTu6LuAd
xvFnjBKiMV0Fu9nmvDr784R9OWAFr/MyLDsb3CGFQf/GVKu80ar0ZErqotyOoag/
qJ6EMKQz8MHOJ50YJhOPE8omHy6WtfM0Rtj63r5XtZ93fWKB64lThn0bRPZAFUk0
Ae99QKueRnF/cIuj1aTsUt8hbL32/URXFkdQE1GRYX9fEgdclBcphZdr1PQHMlhR
e9eoICZgqHLuET1LmxqpKUS1nVxDGVfD1oEUvq+VaQK8RCuVSv5g+PgVtPBF7SRg
F802ZwJo/WGdzWr0YLSpORH5/UC/GDTWgn4iu3CPCvpPW6DTp4keYKNgZigSx83x
eKVlFi2/EqzE/3sYT7jP6OFUWp/6psloqeS48KkdD0cF2CZxP0AlwMXkDjnweEAd
cyQtqJODQGIQuEoELO9Aj2G9VyY8pv8XVG+qHA+SD62J0fpRxcEZA0iXWKp0vMOd
rQ01nicdqs1bZOj2zbyoKEziph/g934FTppD55JJxg6skN9w3jiAjv70oUdLzKtA
ppBxi/4Toeu6Vt/Tq48gYOMZB+QlUR2DgjPmSqB97gsiJzOUaXhKpOuyz7ADrFVj
CGPvKhdHcHl8yQo9OPQOQY9DVTmtjkEXF10yBN0UkoFPTyW3ta4HwYeE2FNvA2fw
WOxX6LxusR6McixGXuBIzG+cVFAvK0g8uToxj0f5vlJyljf0WXqSzRjwpJB1id4x
GBwj/ZnXvLIExuoGZa2V6vQ+ElwN6ol0C4BST2CM5z8qg7dDJns/tqDR7YbA+w5k
+U+bXSM+6s1C7d72Z3Rk8/okyrcxd0ZEUii1IaDZFY3PhQH9wXYMIu9bCJje+3Sw
Wp72bHiuklN1OIMjfxKfnxPZLJb9r8xHzGZ1Ti18kl+IKJd0X37rX+3XcBzqvONN
DRGRTzaI5Fd8U8PMwO+Quc01mjsokF+nN6C5NiTATh2hF/OmWcLEuhydEj70gEqZ
TywyFm5X9ZU+RCwPzUvnRCyiulvBKHe6oUsS1CkubRSzuWcNjzdE7rcbLtHxEmP+
rdZFMAAf3egZ3gDT+8yznzN+ItAL084nHMOOrjVPbIaY5QShJLyakR0fICnEih/y
ywnYEkzGUa5ZPqbdvyx8K44IlGXgFb3L5tSVS1bRP0wCpg73fw62Q4IOALKM5ArP
epa3RpnhoRRO+f/DAQt8Wr5jKEzTPmEwDtnRyD1m2BgS3KJTigbneoLIdkQSkbi6
AzXW+wTHLsbmDQxN1W1KN9yN32yutShJJna/938n3peyE01NYYHStO/SsPkt8Lg1
QJYRmoYIzlv5840q8Kw9wS+SrOOLdMm2m+GAVtd/2g1DuUso6nftBU++aSaODaox
c1n/L/+QqQTB6+xv1CaajXRRjFH1A2u6S3mrXpHtAOyDNnl93isdr+cSSmHPniLY
y/xrii9sBr7PMKSMtf3MoIjfxPwmu71d2Dy4Z5z/XjAxuvK0qR0D2XjMtXde6iMo
9otM7Z5bC15C/0PD5ezXcP/0h6/Gv6mZwdj3ZunZRX5vZTl85xVJfWUBVjibllMm
IXkcf4r9NmwZf0D+y/daug==
`protect end_protected