`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
gMcHP74wBZczB0bB0IzoP2xg5wC5NPjD/GsvSQ6VQgzYAsanETMwwsWi4yhFtJwv
5kY07u0WerSDf8woJ0stqW5xF501W3JLIS8KMiCOd55RHBOnavjYiaaLeu7oUCmB
TtTS1R4sO325rP2zOn9YwRbyyS5Ljn+PzFZZUmkt5xMca3p5NGqKtZW2dV6Babni
5HlLuF20Au601B75m2nv+ZRoGSrpkNElxoTibONmX8gBflpIVE7BehhHwaKSucEF
pp4QQ5zZAZjEC6aplZepouGVggAulz5AahlX5bf4opOVlB1J7IrgyjENtw6ysQ/q
DzybQ+ipztSXBGhmcCVU3A==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="jAI3OJE9Sh00Sic4PtM/KZ4WjwT98XM8AMZrZsQkxWQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hyw9IrFLPQsjvXplweG8O0lkaSLBN9Ijv4B5VdTRt6ipKJT9Kzsb5LxCKvkQyF9n
sGPOd5i74hRHnkHfYISGkfxGJCa55ieOyFShOsqTKRLxclm4oja9vTIey6yFm1BZ
54IDCG9h3PqfDiTD847UCSMRvFssyycwv+BRHQMQlFs=
`protect rights_digest_method = "sha256"
`protect end_toolblock="BnLuc3jxknmZOyxfJK70E5kp9u9O8IQ8cgkXv26kHA8="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1744 )
`protect data_block
xABArkLxBOK6xG+7CdOOiGu0zbCbHMrEntFfAZEE/xRFxZaAZl1QLkuFI77OC2KL
XxG/mrHJzO3taVHgwRXNLDdc8ePbxbAiQfzV3NJLBO+gsBjmIymaCa480cPNpHLx
MvpLmpyOzKTdfClpwlkWJ+29TTv0vxT4RJ/l8KqlM0xnhIcA9QwRvfOauDJ/SrFR
QwyVNaHg0v9Zp4cPqfG7wSz4x8+vsvYy8tOhonSKxD5vINDNpVr/fS0d3vINLabO
XKzgT1JITgfpSz65GElxrZxQdMDUOjnWxA78eawZpHaTL1XE1z2QOXikTQoY2NLg
BS8pGfpAIHKbvbjsdhaQnE8BfNoAi45Xfuz/oQHwl2m6UPlU4Jtqaz/xMdOVWrGP
bzXI6kU8mrzdaM7eleQEt5Jb+GGZtpeOdEF4ScWKBk8enEXIsFOHCLqsZifKk79A
bqYOqphu9VWPOwzCwSmwGDRehnz6avWZ4gM/gBLVsumQEApk8PLhnY2OFhq2jZgZ
HczLxt+W8PtE2TqwxJZ8HDTHfw7QCagHM//BvbMbSf3DhctRCLfL2kYXRbsu9y4R
I0QU65NiX3VmaADXrtAZtxZfkN3lLn6atBFu1UMNLSO0sAZ2s+Mx4GtZxZkrBs3U
M7k7V3prLi45aedll5jTrZyUX1509JY6pZ4I4YB9aaJzTDkSR+mbuMPwOGOdxYEh
iNthtajZ7h7RWmBP0qwCK8hE+wqKVEW+u2Nknq4FjYemW7ogTAbhsR0+PW/APYZH
3uA+njt6VlyAilBlJ1PXU3zYGj49GfeCL/BLvWRR5M8Tqn0yIuWcQ+dLrXjiWL8K
gFCTZc4JU91SAYF6mFMGK98mb7ZEDUThnOV4qMn0vSWVjnJxKD3OPhEGy+Q/Eqhj
h5VIHKIAcc09JGa29e8octeAk6B//qGO5UYkadEkIvrPkWlcyClI+sDT+6PIMc1a
yFwEiqST4zIpb0qOPbRQqRueej/7HlzZfaVkuZKgeYKVprD4N09Ci2HPnq2DGRsI
PTDD3psakTIPaukFV0GPM/hHONGZhofZ0SkkRA1AxVm6oll8/0g83wYghWEX/d7Y
SU9gfDE9jior3bGXZNcAedoRdLfzfOHSt4xyv3NlVygSky4QJFGbr0WDkYmR0LwF
2TlyFD+yB5StdA61lvrI8Yx7iqSLhFyB7+iheTcaylziXiEoHPGvN3iH8RTKXzVK
G3TFThn3zCK/RZGkizVpOBYdom6Ee00w04PvmENB4qZZjHrHh8AzOXG+kJJqvtoN
VTsSkVDkpyEZFhw3eDblr9y+Li7dEtRaIUqXwZPEcsBHLEbwl+XwZwagLWDNzZD9
dPxVi0JjwTOsdUiW67lDkn9ml2BHa9/comG73uE0wSvU9S6wf9md2CR/WsDlMhva
HPpHERHx9j+nO+GVjq8cafTOSZZktmVyygODBpNyxetkOGdDPjfbotSq8jtquWMw
z6MY7XaQ6m6YVdiUFBCJ9fT4d27GdBHBfmtFovQEr9IB2MSOI1o8MDvWRLdOFmV6
7RR5crPSthcmtkt9s6MNEItC3j6d7shsG9s1zlTqqCPAMXR9guniaxoPWDepMveL
loLJ53h2fPpEhn2M5zG8v7kFc52Wf3S3HvJJwhfUd4C+pWsop91Kl7086nuDvOtC
qZwnPAbBHStZdzmfKV2DbM293fAx5ookXxDvyU4kVhcqk8wy9umpfJ0oDVZB8/Ci
6JPTp+ycDid9qFiHN869hAYPwV9j11ZFG27zKKiUKO8kRX7VnRviqpQ0B8T83hPY
cGMDz3/dcT/TeqdITAqQD0u2qDZ7uTFp5yyxDlowu+iWLAcvHovPU/T5FgmyNvmH
kg7QFlcSAOY9hvAjqKnfZcYAP0uIMV0JxDa3tfpz9h2aTq2uwfVhIZdpHsxxqEIm
kHX1HvFp7kqOLVoEXTMTs4MjqR6Ps23sMnkUczE7EmInALQCyAY1PDWlo0ooqGCN
ka9Tz5qDCds+jnuwUMLyRpuSp4/+uheBEcyZBXGDDNh/GPFHgyi118luQVLJaZY3
AH6AHp8egXNa9DphBKOQsrTEV7Sbak6s3ruAxjvKR00yCkKVkCDJhEJTZiXy8to5
Nzz7D3hO4WgCfC0P2G2FtQ41sVqAgbZkg/XkMPfbxaSTZHoHv2+kdUb6LmKmSBFv
6kTXfNxSCquAaHJyFr4+RE6lPJxWNqyHXsWu0t3iSRVI9ouD4acbnP15Bn4P7ACx
wXNP2Ueg8gzkT6BGsxsmE/HbY3M9pNdLwhE9uh3QcWOOW2/hf23WajmPtS7YpxF7
jMASl1UfPkpnZm9YMJjOWA==
`protect end_protected