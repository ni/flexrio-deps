`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7184 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1wB2ShNYedzmkmBWjqK4Mg3
8iDfXbv5M0vDNkp8sRs0MIcU8mAJtZ4k3nFhz966ecHsV2UcmBibUY6X5EoYuy5X
RLeOZGxkDPn+5rGawKtwGGwOno95P4mK1CTmiV5HRxxBJ/IZBKQGN9dxPJfZLQ3r
Rmbl7IBsAG6rCI54yFvYLssXPvylB8q+dodtv5kHhkcwOhWUJcmRYrqbKoHr5Sko
0Cu3T0jl0eWNQjClrZo6xvqL60dqk+2wmSWpdkV7bYAGFKmOJX2ruMXJuCWKft9i
Y94RvRjQC2psIPYubBC8iqm7gJkhuYL5j+hmWc+YyBvWi26OrICvd+xRjuyRA0j2
y1jzl7L6fZlyT9xIXHeGzq3WTKb4xbRTth7RGIFOGfHhkhFQTRT062wKSL4lD0Jt
cyP4p8hVHU5NrfSYVkkr4Sm8O/Lw+vZWfTGVnN/90ULNJYCeGV7q8o194DtfTy+C
Zju7G3SU/PNusRIZSEDL+A4gi+8Qp1tEB0rNvBqUZZNTQDpqwf17BppbHtQ2nfLU
f7THvRhePUPFcT3UMmZrnLY58i8vMXhzOA+da/akrZI3WyEZT8PyKa3btGrjS66p
BYRtgvTmJKYm9K41n2lO5XfU2NYX0mSIo2zlGr5LXsK6vCGFBmgEtA5nATyThSoH
zaXRm7Eeh2uoxt2BYQmSlqt6LKplW/RKGjIyW2siIVxAcxMirqgd34SlG595woEK
bzhp8+DKiBH2FAanQYo9Ftc1a8LDWKHVZ1lZYvSB50gmezMUSvcnQArc0iSdMUVS
/bHX/dH6Bxz0+ENNjPoRt/G0802K9CpuXHlROPhlbC8jZvVYfU3cca2jXrdGO7hv
kslIyjSkleP9Gg+6BXdJN+QHVVHBs8ZtwmQZnPsD/qcdGrVB1hHzV0wnH7P2eYoG
SIaUmOP+xhShS1YrlzqNEybSI8+NOVOMDfRzG8ZF2KLgYkAvqXK5fLpZmzdx3SA5
SP0cF9aNia1MZQN0sbazvurdI45NYKaMeMo+R1pJyAITG1t1giTU09pxsSgTQ+7n
lFoyvoWrpYIgHY1rAkrFC4uiSB1kT5gEIs6868lI6rrBLAgQhuEE1r2mbYrZILmp
9JzBzDCnxLSPiy6Q+AZER/sCLuR0RG/J7WHxCIYtSzDjkA9iKevS208ee1M/rPQA
u28FKsN0gFyCGSBHZmDsZzFXK+whTWFkNDM6IUP5bGp4r7coZU6PJFi1lELGmpiM
FVKwAAQxZtKj1+Q9aH7CWvV+DvoPOq0Bc17ayKvVygcqz1ZypcubUjeqyoYuhhiQ
u6DYgZxBYxUKC3GBEXgbvLwtwK0MndtZ8c3fhdULjDfVotTldTPsc9gMhVsJ63uT
zz28ii6bWUu6XMGwI/+cgVZHsbsY6Ix4soAIrn0OjaSQlJfPJQDcbes/NJEG4xwo
ed2tACUZ+Wxt84Y2a+tjMf8w9HpxTpb1DeBEFt3YCtSgDUqXhTe1OpSpCqZqEFnA
8Xsc17jOLRiCQK8ChqwBU8CDUE1wkepilDQk2DoeDFMo1KYtx4NlDRBvki011BGW
QQ8CmUggL6Fe9dL/xxP7GXnFaQfPAc8vuDc9G/xsl2lEsL49BlTkH16MPiYPEHw7
75SEbphEF2Xn9ZjWjlAZjaU5GSg6n9ngsauL6NLBHvbbDR8EvklUi/X2idLDTfJb
/TQotFD8Zw0/EItLx0dPnR+Ev0iYtbbaX04qxsKmY60HHw2iO3Ko7xsrnt0jHDt1
EXeFbAaJTdPelJnoR8A7ZdSFX+/Y1E4+cczam/hAwORBuDVNwrBcKBV9KJT5WWIe
6Cvs8LoOX+Y2AiHC4rFnZfDBFOSdQXqwRXQTDQ4cs1P5ijwoKVvqF3u0QX3IRVSj
lPssMKdFGnuQ42ppnefoDPikmYDXNtexs/8ySmRcAkpqLPGz2GWCs+46bwP3LEe2
fptCAUtN2TIna0VBkDBalb89Cbd2XK0Qkffx0tRQwGLM4TDPQ8ftwyjK4WlZA69G
5fAm7zkJHpcN9Rql6Cxeo9WtpqlE1Xw2HOOiZyU1fxc7RSShBwJwXLpiwv/70XBe
Qt+ZCAgpiuErGh/jozlB5XABTM7Uj3WZtI1FgT88/dVu4OvQwx6qceBhTsD0s/xT
PL1sQVb77ssQIBfIat72ZErcAMPiNcKd9UbVKsDKBNXygw5b3XDDCX0LQBRLhgMR
4iTcDyY/0g3+5V8yG+526W8IPjdkYd1pbRsWJ5YMz320vslLFglAFQno1w7hou9P
mZGzAO7o/lb/74cvu4no2tBPqGrKXG8khF0LoKU8Ga8Lyr1tejaBjUIubicOLf2c
54+WyQvkP5ZlfsVZm/qhD3ffBhuazuPaGaRvLrxJwqY/z/GryT49mY2MxiF1Hvci
zKr/fniJgBvYPmgk7+z3O6H37x/7Fv8zdmQGM7V2Hhlf9PTTJiu4rMv1CPtpRSSO
mtl/TQLuI1gWbKjW2T8h8+21bYexunnnpoDN7Hfe0GySLOx0QR4/WVqXVuDC8WPn
3CqIuxdaBtQsmHgzm+4ukdPn9Y2/4kqBbl4JeytKzrzmC8AHg1JSS8afxtTEEsX7
aRZK8w/MuXA/SY1f1ydQY7gODDmcQxlMZ+kPa/IN/ncoQj3HNoWqlC9l1TdkrYdW
pCY10ixL0m40ohFB7WCo1C3SMSml2UU+BcJSSx8Cm1S7Ny4aObdDX7IgVlNaHQFc
CZsGzwHNpWm3WzURck6gZnnv3yx13GMuWBO80l1QA+cTM8nzCjMDy91xPIPBnayW
m0FZfYfcOj0JjYufQsJ0nMZhoVcSY/KgNXiayJWCEQFsQfPUpmicbOtjV3NDoEFm
xrQpQn2Jfe0ki0EEXodmR0R2HuDY4BS3gZJCv40hYp0z+aZue9XduXix4BUhI+1p
/oJRmpc57BwJHzjL9TRj5lolaBvu3QjDpFf1XosCP2fo+oM3/myG1k+CmujM5UAT
/dIOof9k1HRrZQHb4nQ0+HDFnVrYmgCxda1DwW/vSoTjdknBPZRedJ30tL3vDtyN
lQY67d+dx768hFyV6T4TkuexJuUq0TUpCvoRwnGmAyhKkmF2zxrotgLsP5wAbumr
jJTOQzXhM8v3jWKJnFLcvT2pFD+AbzfcnLAPdXl9YAdUoVgwb35VZIN9Pmq/SFrt
H+/2yd/QDJbcdWXo6C5SpRxbf5EKhsJUt5wYEMIwbqeQExGMFwc4+nnpL4O6xh0g
NlC6WuRg4MiSuU5oHFAbMuysjmZJWmMyONAqXJ1VZJb0Bemm3MZecu4HjmMTQmc7
4LAEQ60YMqr952hORE6kL7sKn330AgGpu6hbcy2qtRSy/kK6N/hlsBNbis5RQCKc
1vY4nM1hE4pQDZuPPqdG5afTlBK+qwwmvJ+ymz4FT9EDZJvuDje8SfN/Xwe3VF/e
+l8szQ71mMQlUew2ceMkF701DiRb6sHoP5dVyCuKEMj44KJOEmO2T15B1eKe7gr4
cHo2LxGFrwugrcy+M6k+j/BQhnurg5a7Dbc2W8KwA3n9p7cf4nwXWI1EJobtAH4W
7R/ViEXu0u87A9LSj+JbyZGe0glztwUa53lBe1pNULxR4EMY9lxowyy9ymKFAc7u
SyyomUR0L8a1zicXTFS+p100RE+A917Xw3WwWY9tWn1f0Qim3ExwKXiTBnRPO1kG
CG+6on2B3doR/RqufFj40i2aiVsp0pyRXfuL/12WlW9t7qSWDD6EF1oiRHa+dGvu
t+YOIpVy8VJ4/mozemstGxlP35aL/jsxRyZqyIP74IU9VpAFOk9kAgS8tdrpiXw4
aGvqMWP48EB+dmqkHOwFb2DRZRtUqSBXGzUZ4U2AuTHdbx3AbeM6bOSb8ZufvJ7q
t54PgvApR8GbqO3Y8aSvo3ZjzpNsOvG3gqvExPQExDpVZo8XW2w/5YHq0Bl9o3eO
ROBmdBYN/dLi6yxueaLF8h42aNw+Grnv3m12AzPJHvdUb4j6yysh8M2GIlFuLTeW
2BvnspY0tPfi4jC3FkNuol4jmpsC36vleF/VEqD4eop9uMFlz2lysoQAy/gAqcmW
5ZLjw5fdjzCoGE7CJHBWgeQyVdK85mNZk82a9lZIxg8gDCQ32DZdULpuZ9ZvS+ve
r1fqy6XSFpieO2o2fyFo1PZTmzIsJ1PCI/5FlfNgImZ5RKDpXAid9sw8ORsQEzLY
b7muqBH19oH9ZTiDPo43WGHM9qzw5+nKqPdoj0F06ZHnzAWSarVDiokELrJoFq1H
VmhKwyW4GX3JNyuUn7DXCBBtBVk+rVn18Au5Ia7ZKtu2k7RcBlIe6twnQX4OQh/y
cIxrkmNyBTfwrOjwUpLBt0wCAwoNehovEU5Lmkh+SID1GQ92khPLsdMjIjlHmnEX
dQfyaZGxaThpRBl8gKYzTbqRpHTI4Pb/e/ACtK/BM98pH/NkfDYY+cUXzn63SF/A
FNqnjxkyU+NghwGe4RIQMXKsOgwk79H9hE5fmrTg3udxqqQEiNKFmwzYXGdUFzaM
9eXvRfqWq1Lzgeb3+BobPFjNUUmVTxExM+d3hBmfD9obcDksOkT61trfk3JXEBDK
87GHQ/m80wf7fhb2unYQIpW6PsUQ/To3sD0XeXFOFGNO8fTZaS52AIa5PqBiNzHC
RwtMMipOv39VHE7fBGjqFJWwZDQfpdooAxRKDmZimy8WLv6/r4Y7K6Py5WQ6pL6D
UmtuDuNReQG8f3v2ulwV20uoeRcaPyNfkrZzdYfNS0gfw8pwrfMzodPIP/PcZCqS
EYkqIQWGo9rZt46KFR2hQ0czxrCvoz/JBaeHUEt5kIYywqmJKT8U4mSSRUJzUwVt
+Xdo9ZRPJWaYrBMdZur1HsWXHu7vDd4KMNLf1dwv4xz17o59kbPIUYGfV8omQOQB
Z4wvHX6fOYZh79uhbVMR5Ly3F2y1kiTLDh4EHJLDmA8ngWHX4UiJkhcru1d+VpcS
d9/rx1HXtItK6cXq7ahdQ/GVJe1LJhuiVCm94YOVywqH4qskTwMIdrMAWlwYouiz
6xo4pEqwtV9qoD/GOVlAMmzQ0OrjKTeNTXzlUc3a8XHeEQJi5fN8OUCGzBk83Ptm
s0Rnj86IiRRbnrZzzSboH9m/oUfLw6sOCycwtKBxmn1bZKUD7Ser7jHNRk3qriCc
Je2hUFlJOHLtiigoXuF7i+IN9yqq4csnaQnpl1PbXTBLvkKOM4zIBdDxoAONF8PP
HxTKb1wWt8yUQPBVjNiGzlOKmHFReg8km/w7mA+crsMlfjVenEgnqxBshWx7lUXr
9xXUoli23G4WhnQ0ESUS83ZM6Z+FrWftQQf3LOc84rvW8GdDb4j5/VUr8nr6T2ou
FKScxE69FZ/ss0CYmQAcRPSdmpMmbjftt2SxMdHqQ0WoNgE4Xg3rQ753ehaZk27+
dSNDbuUaWKH8OTQcH79XdzE6PE2RcLmtNM21w8VtRtQuOT9D79W4/pBA/my+UOVk
O5iIiVRXiyHR30cg6nfuqqwD14zZia2nHiFMIR/ehGuJAWaLod9artjOb+ayX+2a
T1TaDzWBL0hPHuLwlglzOUcw+Zq7GWfn1tIvv1iUYH8rJllV6lPMIoZJ9ThUb25q
09bLwuYTRxFJpccqsgk2oDYoiwokTyoYwYV9ifeM0oNLgNJ6ugkZOlY3dtKnd3S9
UlA4PhIZRnV6mhFKkIdzOkBjioHAvw8yGD//Xhyh9KWirlMnVNfxo0oL4C/qMZ0S
PbhK7tgKzIeCXVVCgxoCsILQYonacb0uDziixiJDA0tOXPFAGtvVCquo1eki9RPn
Ry9XBs2g/qNvw0pCT0xo6diC4n3JC7vZiUPiDtFyt+OWMBboSNF8I1IYF+pYAHoB
4pVOiXdOT2KCIVOy0mW77lHhFwJe3PWcrWv6fde0hYlPbsCvspdhZuKlCTNEc3SN
0Gd6ViNvSdDvdue6Tc4EUzX+wldwlJLX0RK4kwLCFMQTF9A8bN1lrxSIBZ9fkAzK
Lrz8YsLgHQjoVsZP9kBGCCHeTaZxXApNChBZAUAARk3FZpqdaWRvinXjOT2/s8io
c0KwIHizfHyG0KlXxQkssNNLIMF8xej59MlnGAkOZXIIfgEHUbkSyoWRcSPnfGkT
Z9lupv9xWbbOrftdRcY20BqNWkR1u8kE6CYAlgcehRo1909RMyGmikiWRZpav00d
iniRVWUZAElzXH/yMY+kp055WWdt7rgWtZXI8gIAbOmZNzkGyBX+Tamqq5DcziK1
hNo0COsFh1ui8rNM08GJT7c/FtN6lb5ar68sEQ9/NFn67poWawM5bRWrM8PhyffC
m3ohh9ioYQq+3l1UQ+dhBnwnOBHDwa+8q3mM245Z2ssCs8q/UxG8M+RB7Yi482Ka
lo7hAdNNmqDJx9PLYW0tSFauwO0IkLKoDxTrWz0HQ1N5KvmKS/lpKFuuYqtZ8GL9
iHhS+5NdOVbqCr0ZI0vpOToPjIHX0/QCBjz3yShfYHxbYsMv6W7C0X6XjWkywfXg
DEuq/v0WkQ3uGdqd674plp4OiKqPgbmoWhGswUMCBrucX/3mR0Qv4Utv7iL5fbww
SlFPt+lutnhDHclLp/0J0I8YekuW2mG9ytLOvhqP4QCfAfeIeJtt9C9FdlOXHFO+
o1NmidYc4qJgh/KSfMO2Qj69IXPDHFY/LBFKg2Dqr+B1ZhQU+/4pkB7coo9ABaET
Td8qond2fJtARqsLBmQwusYlQn+4XXgOa5L+U/c5Yr8JzVnuy8UJNHkvIds/Y1Zt
xWDaAYYxCCLjZuXeQAltxlN9v3rJqZHTIE4zIs27ewGeKT/Qi0H/7lrIH/ypJxl9
t4K3fnncj75mTXTN4lzEc3zVrEjxcr3IGqVwo4szzIfb1A17N6Z0TyzQii4xLELr
9SYAZApAYmJfX+Ru2yOvBB7eYYYnXNaOhXN/VxCap2zIR3xZC5t4GDqD+k1mk677
WcdQN8KywMUbMQJlYS7AZQdfOOY868KQt2kHWC3tmxF1fRzkwUmQqccpJKdjx4Zl
UMn2WkQLMamtiDu3YFR3Gekd0PW6S9pFfUBSkOHQ2HRdusHKUZnwZibA2opVMx6y
5ZM0aSWhFj0cpzBYVVYHSuGehflU9oe11wbee34a9W4gozA/5ECAPEXEU3CAuH20
hN8Ps/GtdLs7mydAzutJDKgsDvOKOIva7fpEvrz6BrH3HGtruzss95OmZTY1qa9y
MqHmv+E9eUJcEOzPq22ikz/xMriJipJMzah0aFfXA9Y6PgHWsZTSPFmgjxIz5fJ7
pMuFa121elK4WaIw59k7tNmjg4NiXBQPLevxEQy806qU9qg6hiyZfUibxTAWewm1
zdUvC7iLo3iOETLe14Ddfxn0SrtG9SWzu1OQYEstgi4mfG6mK2XwDxI0ad2LEzsE
r77Cr9T+4m0tcv6Hd/IV5d5kZa42mbjMg38/uKPjgxIlO/cUI+B5EA3YXbl6DHzB
tUtw1yBD78Xonxuc6XLQG67TfglPKhRfZCHNDZ9ATdMjPRokRVAbgNtYIPBfsbHi
39AYRFVHPPS65q1jRC03hVbxfpE7cjuKozHsmtYrsd9oZVZirJCzQFsG4f6fieg1
T8BwDdyJZ4RiNJoxJxShGtfVjMSYWqFkHlFepBFoeAkm2r3bVERF6U5EFl/P6sEK
PmNufKjSsiUWVlCptIn40vlg1XxgfvELvV5/UgVM5Q5qgftQCHmUBM2IQBgZdmU+
GZab8XJhni7VPSzdbyHUk8032iXTMrMZm2QwhXAvFFu0F7JHjX55AQ0oggbHVtMa
+Lihk7ql9zrQ/wUKrEjOvkugpz1Q28J4OgnOgavqVkvrijZX6tCfU6lWEQVAsg+X
lwLW0uFt9Ic9bTcoQXxJchWOqHOGddo84ZJFNdLZesnuwXExyqDJy/z2MTTPN9H6
QKQSJL1IuOu5le8iDhmiqmA/DTyWjSX7U9EE0r4jAERUBea3Kwz3nl+KwKmTlDfr
mQG4JZSUKGFRL9YoBRSuRnVfEUwnGctgqBT2zIMTvVkecWW0UBgrw8pX3QO20RWh
ZJct3jarqpWJi0x5Qxl+CxsNleo83Ve5+M6+2U6Q/CwfXpeZOVb7WDmrDb/2ae9Z
Q75cgXs9v4smCoZMRAtHfKFm7eG6Y+3D4WZJ9Ti1ADntQlFwm1CUR3fu91P8RVO8
kOdcvW9UJm+jCj6j5uzK1k9A26lgmjrdByd8qEXibrJJJhFLnIWSPDoRxSUBjjwx
FGL7ueLEikLhyNpLAWxWzDBn1tXhbkV4KNyg1xvgtjyVXF008MvjP/qPzZGSsoa9
AcWykZ7Nz/sRGG5r89WLCd6qy6tk00aUsyAUlRb61+dhKlp2zysVXwAn8xVrUV5A
0cpVAPFQy1DpNJr8KMSf1Az46o5slqs8Kds5+/GcIMpB17+h7ugI2Nq1AgQo7fdb
X2RHnFtMVUl7Vk4y7CPeFP+U1sfeHTucMFGhowap8MezO8mu0qurTv6fHUoi6UIj
dZmnutfsdehtvxMCfO1iRR9VoFOA8frNah8ak3F7G7Bxy+k97ZHH3GtqRRSbWhpB
//7YWWwXz85GWBR1L2DZfkayoEuzkIthny++L6lMC9hwShblyzj9NiaAh5IFovrS
ialgoUOYBGCpJh5yY6NZuKeTbgC9Rp0C5uZjRFq9ogFGLFnb6gr7E1RkDOy/8rzC
mHGoRRUJeSOQZ1Dm4l5WJ6oj+8sV11WOAuMFhgaleGvPTEuhQ9ROwgNvb0pNPYok
yK+j9VVNW46e5cMxSFCbBX71JHSDcf+ifzBeMV3Fnk8/HUOzPbjDLRE6ZhOzsjdF
BPCsJNljwWJ66iSH/O6E6zJsS/CZ1TsKfzdLmb4XskxW2sGqP+HRX0B7+c34WCay
xLizX1hYnC49hPj77N9Ng7WFuFs9ROAiYtZuVisJRzkEDO4DmTP61ri7Fugzu90X
mfiJDylC/PBF7HtRa8E6KaM3a4sYqPfo+jnNZ9TuFd4A+f62D90FIMQUDDK7gu0E
ZYO2OsgiUydm/tLry2QCqCtf+BzeXfWQrx3yASdHwp0o7mMBS5uXlSjLLXu85590
YqNaE1Hd8EdBmLRH3ASRtALpiEsEl1JP/hsHcoL2Gz3KA55IMQW6g0S6dcozROBX
9COjMSQbSepHMSx+WVUe13XnLBCyFxd9P2ZRDl7q2fOjiX6fORB1oo+3pdJJD9+t
CHqJI5xFCho1dw8g7DC3+zzhlelSKvs7hMQb9Rtwb+cd7ewvq+rSPrIh4WqGYWg8
kLjDMSEVr00peo7ZQ9dJipinkmpBmVrp2etbCOrwAWSEjD4bYpv7Pu0aAkK4BW2l
wjjt49zn3BnHq3TJAWea/5ma84doCyciRCXYjF/Tkndc2Iynty+lZCdxGL0F2Ze2
B4sV6CtF0//1heFMRbn1t7dgAzekVtzoucH/5qbLq1gYeovNtaq/yFDiIhd6RHjG
MlCWBxdd/fOeCyx2fcIzi1BEeufcOKBlNgw1TCIkq7o=
`protect end_protected