`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
j9eMmSPGcKCWAR9PvkqZ1R001FU8QKTyJzFqNLn+qur6INyYDE1AI8LWcxAzfnTc
IpZG7ua3uuk5/kQKKQx8ZIPLfmv6H3t3eWjki8YIAtY/d5E7Gq8Z5mNxMYRzGGTg
TCMm6oOrOTVYlCXHE0X9AW696Z7UGfWirVibl8hs19hrFdeZKGiGht4r09vHR+Gl
FQQmSObM5aSK5wu5KOrK5ZUKGHyBhjnIQO5NnittDjOwxV/57nHVg0pdG6JUqyvm
tEgmCY36RCMRGWN7sekPtNHjqpZkmYrVX1T9QF3h73+8ZekZYd2xY2hpHHGYYeWA
t3+Fmb/6NUmoP8+Pt2hI6g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="wX+NBVcG/A5ruHK3pkDqG8ZVPdOz9TJPJ5saXZYSeQ4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
j/hqWUoxjK88VtH4QmjIrexFOSwtsLKOZ/LCP4cmrqgzmR/e71apdtoL+o8nlfy6
eZxDZMmrZmJGoazz2oK6kz7xJU85UCwNc4cxAsVxNdCP19vZxph/nCYZQ9lUFkLH
uLBkOeFP15CD3jG5/dp945fHP13J9SzB/L9PWvDC/gY=
`protect rights_digest_method = "sha256"
`protect end_toolblock="sqDZkaglKf+bDjC7VKm3lOELrT2Jlynh4UhPg2J0Q70="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
f9kZDbPp4NLiAOFOgATj9W35i3s4a7wbt9jeHjHVcJxMoXY8rb8laqS5bNUhXGW/
MOc7UNc1VwolqhkS7G27SLamkGClZZtXSbRcN1N+5kZpEaBEj1343vVznnU2Dre/
MYf9X0zKxDxei147N7THFKz4ULcgO0HYZk0BoJi8sXVCy8qOuCcWR9jTYL22npZW
gdVeJQQ1+iYPpnyWHrB9ttbMiXNoZTHrjvH2IWhkTkWPK4eBSkKjtnGugNazT10G
OLgGxVOeewFMagrIjJ2aYi2FJuZPtzPpn6PEpY4VsKyP/kSDKT6Qdn5ovSQp2yT9
3+IOH1chCnVjoKfyIvrFJj7wnkPn42ZCOCw5x7A0ysPKVaiXcwW42nk4v176EZyz
UO39r7B/8YcWSaIYWfO8fWxxrqEZc7mWTeNEUHmX6QVKEECRkeTA/zJkjyApJ5AH
j7zyi1GClo54qZ2JmPdzLyOP3R+7Ayq6Hn1K545gAEmLOwacFzLakawObbcIqo0C
m7z3Th9b3A+IkluLmWUZ/jTYYcMEjIkQuUAFx9ynJ/lWFGhrHv/NOXNjztk/9rwA
j6qT+0a3I10fltdo/sNKbc4tVsREg96DUtjZ5KI0reJpO5XwTk2OBeVPZVkVSI8l
mmrQO7g7j7Z+rIUC40Nwd8jyjJEc2DrduRj+UcQlZAMgOnJBGI9sM2QTICO8cVHK
ap4fPVP7MmZTZOMOEPd1epMNslv/HWdTEgDUe2W3FE0/llyNGUSHgHEB2NwY4Dp9
fS1Q1GNCPXxkOTcp/x9rbwf44iopEf8gKT8CkULYdeM+Tsy+K13OPJxB+EBbS3wc
koTn4c88TzhzmNhNHYzCELdsOHL3ciJpLuCO8na5QeOR37O9iovfHoVRUwT93WtC
xD4EM9nRsXf9+av75nDui8YGaKgnwz+rhcNST+VVKwkMaeehDcjCht1VEOuUCW0T
59RIlhzo+B7YQIot8eQhKiHGT9xSmHmAUOe7FTCqY3iHa/cTO21uIkDpGfR+ySC7
1wxhF2p8tnIq26mpclk/zNygH6oVbCqGJAxvtEMQVCrKQWLQdUqxV4ozBLcybkXQ
fHP+omw9iWG2wF+qtCLWDCGvAfQ7BvXjV0YzX0mWsK4ni/1FNjyUWjAN97QwtfKE
y8VG6zbkB92IEe+/6/qB1FVFz7vLFCRNhWPKF1JvIvRPBnzy8Abp6NvGnKB6WpWA
Vfz6IEs67xx7CMm3eKMt7FBa5V+P7Jo7Yv8TfzyfzMIEL1HDwycH4SMV0Y+0ftUj
qCUYB3MiH4++0RU+8Avwfd8MqCliSwHeP6ceJkhFcUiXK3aYzVJi2hR4nLKJRhTw
jaSE21QVAHRLj6HN6EElanDp5FN8lj9BfE5SXo79xBwB4SMP6NDvyAXqD+/AA3Os
lnQAiIqm2z6/XkYgnpec9ZdCwDYWPx0WFN1BFdtzCWM03Xow/iNVHwz9bOP9SS5e
jtPT4D2iQzlqyrC4bmRpBN3tRAMr939mXDnXVc+OXtgUNs0hGZI+SD6vFqONc3fc
iMsjSgN+uiSU/E76ROGVs1rXQKsjcdy1cRnzNnkEDOBqnETH6EvIbWF8Q4ZeLQjW
Nhn9+Zx1jwDwDggkhmRHqh+mg6qxt07PtEO3FxgmDBYzjTEVEgIj4cxi0LXa3lKL
Tmx6zobDSHjW0ed5ZwvWbfd+mmkSCQZRh27++IsDtmILND+lp7xgn6G8Osc8ieaj
NwrTyGah6wuJ5en/dAGB+57Os0evp7DZASzETDxP8h5O4OYl9g19jTL9L66pDIpV
U6/n4iAPb9lnEYFnyS5Y+eep4Ag8JSgipVxLroYAyTKwmkqOJSWUmAcs8GlPiyXi
MUAZAQle+aYSS6omnuX6XDJLx0Nenk9MZi3fu2A+T4axC5raMVGblIJNRT+O2xHH
i1CMQnrx62ekQEBCGpbCnBXe9+AJoTw3/BaMKlQr7Ns7Zfw9Jp1sK2G5Nw0tHgo0
5xkZkme73PI77vlLWu/ztFg9CJmLfGtInFO/f5DBqlVPWLBoEIoSM0yOAI2t8VQe
SHXtudU1NP8b62+WFYGlBLF4K5O3013GYW9awTd5OC3fRTnm/okMh6FIogCjqVFq
0KDPZDX3/n/HtS1aEiojAPaI6/LjDGaFsYSxdfD5AkNPlN9un/vJ3I0oDiy5M9tI
rorHg4e9wwG68X6WbI/TwPbTIZRC3whyw/HNbVEP9QpXMIdYziy7waM9Ap0Ur7us
aJM/fyw5iSxx/HQEKhpqDFYk9yRrie+masO64tzgefT35V74ROpY2OkYv2NmWYUF
VYYTC1tX+cN+KXvRJuItKgG8tvEGv+Hbr46gjncpehcpXT1quMpWt8CHyGUsSLFo
tcN4dpN1jB7qouTYjxBE6CmTWwypLEdFlL3/sIw2X5KP3bYC8DoHLiEAWboW9Uxy
B9HzSwA+Tg1GrR9WJ7i72n98ehXChdMPgf9Bsip4r0hKucBZfyx7rwa06uQFbywU
tJ/FU8elaqzEHpqLBWVXpbVioy0zhIM5jUSi/ebwjGfddLKPwZDxDGASsMTXsf/U
SIj/4LQYrJ+vongosY3WhvNOGMTco5TWp7mw1FGmY8/acwzODOmqe0AhELKmkvgf
I3qc/vRDD9iykoUkXU3f+fif5xQP1LV60A3nIVQ9YalcKC4esj97RrXj3eRlN1Vw
8/i4n3rpoLnLKPbohKi/naNzbcspJVA8hILPleG2N9jvG2i4QsIVmZZI6/5qeqxk
11uJuqVhWBHBTXKSweG/gCQBAqRjiQTdl4zQIFpi5ebJpFBfm+o9PJHpdumTiCw3
ia9E/Vu7xRQQfEd6FpT+fh+YWtLISWVc5Q6ir1EYa6B0Sh6FlF6ZyCpTM8BE26Bo
3neWrmZUWZvUh50IrkfX/rqvGpnXGMR14SyipRQsQdKlTCJFVQt+Kjagzuyf1pdJ
OoSrTwbbSGE52SDXQ5P4vDTnpzD/WKCOYU856h/mtf2av5iardq5/rLAbz/ryiLR
McMcxI99yk6eAZ6qkZYw2oP5THR+SS+GUj45xVjDKLe1UJhbSAnaSixtQQhMacAl
7EEVJGQ0fyeF856l9/sov+OJgDC1UHo5QHZe3B2mFwUT+efxLZIgma//f5GHP+cn
PrNqJg+gUI3mkedlOxTS1Jp21EmbCpFNKsps1fO+Oh3ESbPXSqvEYcHACKJBr7pd
Jxf60xuzAvo3aPdXHdakc1mZknrZK1TE1AOF4Glevis2feLEBUZLghcNfl95STZ4
m2ToeXu/U5h34x+SP+/eZdfGLP2cjoKSfKS03hYRdPbWH9AmQ4WDW955D63vLWk7
1s+6TAki49zh8yX6HrIti4kpPJ5STK6FchTru6p/9dxN3AQVB+oAifj4va1lNPFL
WgS4yuOtWsz1IBxR5w0AQKeZ4Qs8vIv93F7kE5eHQnS321nU6aFNyYS+uApUMD0h
7JcVZ2kYfwzLsQVohFxlZwBHYEgot1+2L2XirYPECQkwZt6Y0NCmgCB8DwcO7vOJ
Sj3bhMAvl9S4jRI6VtwAqROejEdBQL/bzhiu9WTQTpE+3ZbW+hicF02Z93hLwMcQ
3MUFNDvJgbPEKdXnZcJ4n6QyvehrNG2upxQfzVxT+JYnES9fW29e9nYnibAq73gS
n2nMQEBYGSiczmTpzD1EvolyoN1fKIn2JJBzvutWMjDDgORVEs2ESlyWX5ypSw9j
C/8mPXC1xRsCJD88K/p2f22AYRxE8rG0oEKUOgwVn7eFfwYjd0IECNYSbHVzmxaI
5zPx9JQ2AXdPSiMNDIyN84vAcxXKDyQsuJ7NtTKHpyxRd4AX7K0hj5tWhGNJgZsm
v5Xa/B1g6Mgkm1GVSzy9K4mp/GqdUTHe9E+rlg1n/uVCdmCMQKm4/f24MdtcY+ak
GorVr6ZGvG1FNwFWJqxMV88kI7dgzJvngJw4n3x36qzY/1hklcRVUY2UGOBVdK8f
10ny4zqXdawYcTyAc2swVEgC9lVgEiAteP47Nr8pnTDX6JDpD/mBYJHvhNFlbKUG
ePX5RLkPtOSzQWmBbcGaVECI60FWQLdR+60M6ych1VikprzKnhe5ja91179x44mP
OgKA245ZIxfRCe8OQt87t3lcW7e7TdJMo4WmndvV3soADDkhKILLYrEckSXt0Hn6
pFjwrpVs5pGookkL1CKBCnPNOz3p7mcn8r9Cku73RShp+Rn8WN5F5wzQQk7464mf
oV78eiPw5JGi9dBdJd+7TE9rVS+xDI9+ZhnQFG7TtPj1wHKGDofS28jud1wGxbJO
+tq0xX+yiXP80n6QyBFwDh2eElwllzmF39LxdR0mcu2OMh64TtdpFMcQZUYJwBwL
bwu2klULWA+KQmO9BWyqTaXJaQiyiur+gnuXsLRIMr4KeJw7HmfB99lcJOljF7Ry
AEHHKooLOcLkmc169Llsh2XVXhQZpLhetHL4+QZrYkEvkLGsY3A6yvtv1+k4W16O
V0cymZAstbRlNGrlGVBUIhdA2wn94HVcyfercjlykgFHGDBb92+ay2ZD3ilj3F3T
Gfm218o+uGojA+16+XyuwlmSbBz9TvhK71XMNRO1LKXX5CTDH25uh/DPrceiMx74
8c0zsytwbBwh2M37BO4jjT2EoULoqu0ErUNRcJa+ZNhLMcEmjq4FeIw0zhkrHo8h
JEwnxvTNzf3auYX+DGqWRq71pSnbhOQwyiOnrq5+cDxdVxpOUcQOImupzYL5SXZF
KA5e4lwjT+dG7isWCUUE+h8+jh4LzmUgwZFgB1Oqr5npKFDbGvWlvueorKxksnte
YZciPqLb7OVBDRTCBMdzfyujzcgLccUPf9nolMfcBbhrbGd/0Jqj73ZOfP3pfYZn
lC1mBXyQX1o86fjEGfHpUKqnPemXggr/131bZCqiJWwMM9k7iUgNQ1zIAYGOxTFg
STaBP5j7MznRU9CdXgLGHSMa5Mg71RtfLdQimhE8gph/IdE455DbRF5rCZ8DzYH2
NHU6h7ERbmoILN7sKOP4eGq4xkWuRpZx2moRRwIB6RcVN+tOZV3IexLRobtc4pNP
2fGKlqseChBXiNOncKTmIr1cf5FQMtCUUiY07QkV0SuZ9tepMBjQi+wJa51gFUI1
UzNd3KNIBdCMfU9UJM8/jbxUZ0wiC6DTRY1+BatwKd/vPZBqi4NhNEVUXr9cV2p2
6SILb70rg8D+BiKQBmxmcRL7ICMTAgFYfF++tMvamyHKtptMFkuaXoGJSYtCBGH3
5rwaMdvEL0ipafhB7Unt9fDdw+eyJslHZjyxY6yMmTSxDUDCUNwJx7iZYBUdJKtr
UosL/I/VIU5VXjGUiiLGImJ8wXKw86h22rFxJ9oOyDGbCZuZ1XNi8YTeaAicxvGr
cF7nDpn993Q+GMsiihmH1XzRt/rSfKwhPcyQzaMqudpswEYwN2ysS9FNHEKXJdWP
OtBaBtkvrrWyNPvSBrpOTTDl6MBXtmO7zmwBNJ4mQvaxUK+fi+YI1MG7RSVBfrs6
X9az8gZRWf9aoiD9LrDY223spoEiOPbNS4T6cyNfHBWRQMZNK22YoQgig61v3T9n
AJka/HZN/wx0smEkap2RfZLFP9n9hyp1rYSNoMx2dmLbxCenAKs8z1XO01aqlpO3
hnIuSWog0+v9hJ3OpWBGJ0aIovS32Id6LxYn6BqEPxGntxZjWMRi8JHbKFcpdcOZ
Sk22l5U6E9FP8bzplFmCKf8PRAuKqN96GTQoOVGSJ5aj+jbYxqQ59Cw+TTeyIv4g
BFDHPZk0I+KG/nXL9bh2ehP9ziU84/hu9RWj7UxBhbM08iI9jNERiYhQQVXAbMnk
NxWY8oLOs/uR7VMNo9MThvvKb5GcF9ZNKdTl8Ey8xeNKuInmt4TclmpgHo32MRd/
A2g2o2HCAV7ylq7VlTD2vS50pcWUNiIwkJOIBz/Zzuq3M5DZsaIxll9vZO3/ClYT
nryB+M4eUDwzDbESOQMmoig/2ggmRqk0jqwlL6TZLtzSZZ5dgfWeBqj2ZfiPxDu6
WmE0JV5HOR5DcM6+jsOTjnpb3uSS4IPmfcy3vnfZND9syfZ1G7plHpSREx2Vlkaf
SlOMBdJAEQcX7pMnR5k7QbARmmGttoSXw034r02nKUXIaSSkBotxphAhvtFA5HnV
mCzUouq0uboXsPN0Iron6FOtkS+T+Sm7HpuewxkYBw34aSk/9aVPjhsbKbXt+fCw
BrzDU9UIAWJ+j2hB1IDt9pi15hczAiibXL8KraJ+UQtC7XNIBel2MGqfarAfSl28
9NkcbB8WM1Nppo8mNxDKL8I1ageKVNANKnqW6XWczDhEjoJ+cVXRb2+uZSaRYG9A
UyH7uTwRIro+s/sDpitV61IE8jIuKbpmGrdgPCSPj/BQYZtRJcySVTz0yPvASBgm
yOk/Ig1PSCVitRAVUmlx6unEKNX9sjIFTqfSOwZca8kDcsBTK+sUjBcp/XoRXdyv
kSECnHAbBhMR+Emp62aLdI6DO/essGbh7o7qXhhYjE1slgJrhtrZD/ZU1K+CkkVA
WSlySTgwCOmeoxBY6uniNJsv+W7pNbqkdPkZD2YlMvlCNqgLFNsAIi/QNUEQwxYF
PPfBUo7V95YqWHYIV4LXaEXqbl9lsKQdvvpgJyvutEeNyO4h1N0BNqgFBNd2Qn9E
6AIPn347vdAHS+sEPzHNORgId23f9hTB1cDt45QhKkC7ik+DBXVjAHPJ8SORk1Yu
ElGbGTSE97WWISS5hSYSIMERbHxXjANdETO4lW/N3cLtTosDK8q3nz3QepXpFwvO
HgzXmzGKiiXDA6shR6dpfNUvkxXM7u8eJR6XeZILo8ftZb/8LGiFigw6RRXeSId9
gjjNZMH716cf4TLK39Iy8NSv/GoC1Ws7ahPyF3vbC8jx09nd25Jpc7d+seCNimlV
T6u6haKK+Ju2moYwoQsUGD5Xm2UgBvJbGLbr9nQE+uUSj49wNK4x0Fw+u0aXpIe/
F8Gp6LctbpotiNYXAjbvZTjiODd+Q7UVBTo2wwixgzx22QkCgDSjdcyrTs4p5cfV
vH3D2v0vYvrvgRumxM/dMJBPQZU6mKPWq20NuikrTHQYE75QzXOsp1krmrXohwzJ
5M3bdgCuZKrxcnU0Xq60Tsyy6dU5VL6iuU8AZIef3maLNLp+/Y7YSMEUoZOom7nG
uCho+1w4Wx2cI00t936SMjIyipY4Yw/XpAqHoHht+Qe4d8k91N3hyTFpCUY+pMKt
SCZvwZqSMFZuo1MEIIre2Dj2spEy/7UvYQXOyS4T2qlXpzVbtmPcsWmXASLB9mOv
iBXDayoY/ASrrheothq/E0scchHRg/CyEdXmUrGPvSRG0DPyT5ebxn4WhY7rHzbZ
mtm6GIdbTA+SmwL4NCqPQZI2j5VRAchodxzh7a5VpAj8T8TXWEdZt/O6+N/lBlD8
WgP1Z8lAMNf2sw+/QX/+54iNt3DE/nZWEGus+cIeAMPeYo3owcBAxRWIFEA1FPFN
vgkBeUfCTiPKe2QyjYT+vuuv4ufNQsBC+7O0Nt5uEM5XlpJq+0HESRUx3YHJtsHZ
OKVcwA+seWxjeHeayTvv3qVtDbhbqBm69P3XkQjyelCFHCF7L9g3qM/MbU39PaF/
rcN2KWvm9z5cJqYusZY4cVYw6mnDretpJRK2kiLF4Kl9UJUhme9VWOieXAmx1xr9
suQWgjOLVka+/hDqVUzZKgrNwDi9miF/2J2h9vdbPCR6AHiL37t9SPTolt+ZuJLg
nn4+pg7943RMx4x6c6PHcXSiOK/v/irpxa6AuR4pyBf2IYlo67t4LBVG3gJUBtrf
Xdn7XHZQxfSO9ohu+qkjCl8n8yMlSzVjIKxDWHzdBngnY/SnzrT0g8i8qQiZf95V
TNlRhWPtT+L0ZSgzQZ8Bd8AQ3WOa2A+Ikx59CDbrhChK2yqYDfNGfLvLdmRjkwkT
r0QrymcgcB5UctYNHi11AaTBADl7vNbPOldaeMN3vArLAuHhWSqE9d1QckXqxhwq
nCvKRPhyheksW/lzPpB3BLCxEcM0TEroNIjnyowRs44NvxnuSLgtezop01IyG5le
fjLSlRzZTuIFBrNrgdWNefodZZ6TNBQDpemJmOfYdoeieUotu+4PV/cLn6jsIAbn
m3BCoAcHFThGWhMXayEQ0m+xXW7SKoTHW0Bo8ECL9osI+4t9sDYOqkAy3Rnrrwsw
UtqS/OYrZnyuoRH59NGpy8sJDpYoLv5nR9Zf0RuyJ9m/ZQGbyQ0FWET7+QGgK/6i
joni9T2u/c/ekJjDf+5bGpjhWe3t50uPkdpYHMWzqkcAi+q7sxZJDJwC3xWUkw5k
Zo5JV0zEywkMWphb8ZsFCA9gSqgPb0ZjrdZKvkvEFa3Bu6culbWVeZyigy37dJxF
8JLEeMwBCAqu4xY0DaTFnTSLu9UkYt+z6g6hbd94a1/tAz2U99hvyDSPwJ8hLGMQ
48o4R7wO6JHaIDswJGcIbJsV7y3H7gi1eA7vZmAT0K8bcjBAmMTBG/WCFqonj7gx
liWZCITISQx2/dlssapnHBIl65qeRuoKXFMfhIxGgoNs5FUqcqtIAFFxKf3xNsWC
H1NYe6+2Z7DGbNo0RJFxWXvfhsBqg7hFIpCwvTKe67K6Y5y57dbyHNPzJTMWfRU1
TJU0/X/axIAtYLStlynv5vmTu8VhYSUWHv4setGfPDZ6b831VbC+DWK7wMOYFUCF
ZgjWXnTTepnM7oJeX9gyzx3To6XlAtVubfKpfNlZBkchPraTvee6jjjTfYBtlSbg
1AXPv4c5odGQzQDCL/p7kPrQ+p3FvRhXgA4tosr13Qk0vP5yPZCSLbtna0z8VTIZ
bQ52oUBO404SZ0lugA4jmXYFE4/RVignttUm9Vw9Ud9eFvBHk3YwHxlo/P/yq364
8u1aOm8X8fuCY6S/dzSKSdoEX0kO5DoUfkv2vbGRwjIw5T0R7UHFHLkNNDN+sJyG
YJHlzr3KySYjUQ39RsXDrnjl2dGx+KHI3/gogR6+TGyWhY+A0+re4YJ7RDLFyYZD
IXfCxDlrsZdXHQ4cSbLv0KVPtad03zacN6rBado2bTesxtd8/37zEUzRFzyyteBr
t2zjBj/SGQ0UdbEFzr0H7vGvoY22Bf1ydN28sMBOd3UYGtluilXaKeCxq6kS4rm/
eL6saKY7DlnVaS0dWEQOcD93Vb2jH825n2/kEb9+7S5LbCFjFKq2tGTLCQAUQU71
lHNcL7aGOHSJu6ZoDAI+iLH1kVHnoGjmYWre1zeUl6N5Nd2sZO4ZIhQmDw+w6SsB
Jwt2ZppiEZKiJ0NoCBgLl799RtIt9JY78t30oyaviNWO+sNxtD3YosofkoiZ4vao
/CC0Ut1UtbTPAGCVh/nu/0XBRphgDoyg9pnIni9ey6ayOjvHx00qF4YU13CTYnU+
QNN72NPI948W8e3aQ0W4SdB7PL59iZ7Tgz8kMskUBvL41KJNn6S3L+7dqo17avOh
vp76XNseBhJwPuHrOt0EcnXKsMOQo7MCTOfcV0Bsxn/lEi1NJpaSP60R1sJm56EP
xS+oFuf12aq5XATpbnFTe90K40yEOVZ25x+RYj1JAaV4PW00s85NNhAQWSd2q2Jb
+AZ9K46n/NycWNKceqz/LI4zSPily2Pz/L95ecyuKBeIyhRb8L6P5nZL8nL/QXIH
V3ZvRrD6ea65ppbOOQVSRc7J3VTGbgdGLVENvWLhzbhkIaQg4+ayqIOJw33uQjVh
phFxQr69/0/Inuo+5vtdxUgrKLGX0txhuOUWQn94vt0ixp9UYGKT2p+d8cEvMK94
zvgqUhGe7p5k+2R5F2jzXg9XYS9UZf3bZpWwzDbCBwtt7TeY8g5sCTHaXYuZ+n+O
27k/HQMpCTZFYHIuombvgx8xVS7j6yiYFRsor7a8JkMJZya0I+HNIAHcs21pnZPb
u27alEt932evL4kfwTzDMJHZGQZwT151GXv3bBHJe3Bnbg8n/cfu+tUuejgXkR6N
2+Z1egVrWBesR0l5wAZLzWaCsIj1yO5Rc4t8CP70SgMR3tUcR4CEqDT9ICJi8nuY
7n3908ZlKkk/MpiO/viHbxy0lUszCyg3/scIdti7bM69spTDaWR3qh5a5euqZqzh
NojCpywlUHLzsQeQm1Wer7WWy3ly4vjd+gn+/ViajCAs6DWdwP2/1SGafplvr/iz
LZXqFB89yxd5cWsKxHI8OQW7KLOUy9yYgG3wu2n7jqX53eh+lpv1Mo2w0PpqrCH2
8ntbMM9WseM8XGONawXDgqLZfGnL07B5gUnAJsMH5JGoGeC1tRVb0lBZ+LVZm0gP
7ybERxMU9hJe+NMYHMr2/HjWVIPt43zcZJni9KhegH6/lqu9eBByGlQxNlwIZx83
y6xF/uBa5yRLn4SnS1d3NW6yRyJ2dMEPeT70mKDxl69GHyJUtWtzOiXzksDGgBfE
XMf6pYcVh+Xq+eIAsVTyViO1/IsSs+dnsqGjFUAsVzdfbxDm1vX02f08UeWFYC/C
bY9EX4UyIw5Mzb5XmqJcXc3u8T99kQ7tXZ/BXr6NuwMoC23XLtk0Gk+a2SrCVu4p
GxQwPByrX5Wijzoki7gkAFgRuV1XKPVuZpv/87NaVT+yB0ZIZbrZnjE0u2WspDOA
2SXKxRvevii2LuJgCIp1qOsDWu3JYN+l1NBhxDYutRZv/jcY3IUEnVNSAyEgQHne
VMlV/VvqjnUfmW24HxPHh9OCnvXIqp52lDDB7P3ja0tcoZyy9ZTNpX2Ry4yhu8RT
UDmOpbZQ91teKogpHWwwZQrrVgM+nrbT+Bp7V1t2INRVmrhm+uVLvYV2cuR0nZ0u
oZDUsca8JizKX0c7rN6LMc+oO2xPb5l4rpkl4SeNhNDOGeYXsct9aKuvGijJUSws
c7V6yUPXYdMv5dIQpOkPhQ81JDI2Q7J2xo0qZH9/zfONUN100snOBKpyGSMWDVAp
jxshxgmxixGDowccp38EZ2IJElYxgB/OirtDqds62PDCtviUbXe3w7oq96K3qS0a
OLUuBkHY6fndvehx9emOzzYfOuhi8gMyseECnmH/nb94/hj1jX7iksYmZHzwjiif
FFsHAsfEgYlVMjTK+nItjCvir1+mUCIC198XBC3F+88+tLWMjEa0LnGcdIlfodcD
xdWjJjGwyov2OwJCHZCpv00nU+krDd23NSssCJ/iv7b7jpi6rONxVcbKzc0sR9/k
NrS4KdKEOdSLVsRlrvq73Ri7YPsGuzMQOXSjCNHLi7vTUYbSVcbHgbNopPutuhrG
fgBUiCsUe5AXt8ZOO6H/2UwGz1uq8hwLS1cpGpWC2QQJPev4y3T4NF03MV91DhWR
XLc2Z/heHs/fAZEIdQijU3ud8YIbjEKQ2+ZP0jOTq0pOTFW76Y2pNVsoyZtVgjfI
S6Pp3av40MZCjsZZIVzg2jkVSqQ9lpzgkYKlovdFqatO6AIhs9r0Vuu3yJlKeY1m
v1tiAeCl3Uk3CAIwRfRZzinjZzZpW5m3j8jFH0I/AJYWUON5Xc8nV7Cc1jYcbLaT
wForicvY6rh5gThIrXmBzrAgXybghVSLVX8eqXn0SmRuQ2XpJb/DYgq2HRVept6I
LUZYen+Yuv8di36alSBvU/UgterD280ddtlbGGUj63kW4lhxQBabovowBup3rkDy
Hb8mWEZyUai+W+PFP3vaW9Ve4AZ/jl2qAC3B4iTV+YR7SGoduo5tJwB4oQ/pRwOv
x9tmGbGSLaPEjzd/ZAkmn2G+d0+M2fsPqvw5uAKL4Jmf2cJ4fhdRMvTiVJY4abis
vrV6b2pCOOuiOMwtTTndNpSWZbVaiLMD7aMrKCC89JSyW6grWJTQERHDVlh6unIW
zXE74n8ZHSUFsl5C6+eC+0cqm94HbeZnzqooHRvzNFmTRd4xQV7nCQHHmS+AuPYd
JlFCNPDOuV7cmaCc5Zq3S1Q2r/HOU78QTsETw4iqRNKmMwIBPdQBSsx9JjmbpwlR
jp0Ko07FEEvh3LsHJYmB74mc3RWxxnBUp0ZmYjxQIobOSdRDlpj5MN96Kpv1G+ph
kFtaHxDmCLpocCu9LS5v7QWONQFIFmS4JmuRwBfFBKcw+0lTX76ttniMNsltgA/u
TZB5XS9jFASq9BoQAtbPR8POmqcaD6KD3gmJd8vSeDmSawScgKP/lJNpEG+JbLCx
Xp3J15tEgEhFG3FneTS0SaDOQC9uKPiKn5dTXHPWzQXxFeviR/euQERGNIDDVzOL
33eGzPA76U2w/10Y7BVfAaddrZG4nl2j56smgcnd7oa3xZ60Jp8byoaWwREgcCfJ
DBF3Y2Yk2RJQsmc0QfQzIRKj7ZEaT4m36dLIpS6LHpnosCtWvl1IyHYQu+1tlrsh
qJz0f0c4FAk5Li4D2ojT5OYIGEtr7CVKIpLKMeHWMzcAK1QEDkBAR6QuXh9z7z7F
kilsSuM4q4RsyGs81C4/sQuML5n21cQiNiCH6E3wRwSOYDyUoBo0KwHnc3oMxTiH
oxiWtHZHaHDQlBybyATwsM8HwcQB4m54d9NQXALuFzt4fbme+RPC6IBpRXvYS+6x
FZElHaX2flMn6nTa22KmpAsu+qfb8X8wzBpIbSR2L4rq/8mftjt2fdMN3tFeQ034
h1u0EjQOpAxgopzmFsdLHxNn57Vq0Pp+p+BuxR7UgN1PEUyOfMj2axiV29++QpOx
pDJ4DMiJHTZoMwwmAXCp4qesaRxTx0jRA+HItdtYHuEit7r0vywaFkkprLyLRK0n
n7CE58FbnNxajMs9hIApybe0FzfkwZVMbKY65wVHMTzem3I7wW4bq1gyPAxJ8VM8
OKTHaTUU/X9pDai4/n5t036gyHC37t5w+PBcDgfkeMT7cRI98CTp3hNTa8AOp49n
lnTIMpO83OfCGeDOfa61M8LiuS7SZNXDq9Ey9uRCAnI7uK3krsmL9ZHEhEtRSW3F
RHUH4TXg4DMAQCGASTgberuEIy5EMav3x5F4J5W600YzcjkjTqSK77Mu40Qi8m+u
U0KHjXHLjOUkV4G3FbCnw6o7Lm/pjPJEBwrsZQ7OM59QwE18TXeIFz4E0nn9MerN
PsgRg0Gx4U/ReAr5jOx1VtX8CD6LGXjJ9JNcd78tNjQ9B0k3xZ2p+I5vWROJpjUO
5AXA1V3urQ0oImeQsmoPwrmgKwn4qOwXi4MJddLBEtG+U57FtBFZWX2cK8mDnr4R
/qlKPqinUCH2vBio4KJdvWIh5423dhlQEnKmsKyRgnhAdrJFtlz70ECiQI4utuAy
zTpGzBJ0uuqGuYNfLPifW21lt1+6G8EskEt8Q65tfzxErhbaaskjssLCz/OscoGk
hcj9M2VTCejRQrOfACYnKb4M9EmU2kJ65L8hkx/EF1PZMWS57Gu2viQkjBPREjf8
+rkfnVHy609FMnvbJXsgYRZ6pv7mQ4CpUoF79yVA3aXFzTyV9ojZuDMMRpsUpMla
zWe+REz3SQ29own/Gus6qe+uGUhCdQCueI441l38q6ggdVdoPkZUNaihKoY1sIpU
nel/5Qk5VpkHU+YJgASa4YiwFcPToVEB76f7KLbgR9VtKoumUID7miz0Jo/LI05D
qjpDsxLt8Ir6d9CNhQGY859id4u1HcE2kFLxVW3HnM1GP89AgJXEnzgKx021ITPi
R4TeHzMb/wWmaY5ZqyNlIq4EoCdZ7vCSzUmcVRwutLaele34WdfrCBrCaMv/Lqre
To8ZrPMrrrx8x7p7E6Lgk9FzYKfSbDPjzJSUCG2+B+lEFmNXFypMxYixpSf/ubBD
NubB3JNeK1wRl9okvjYd0v59TIqAQqgMp3fAs7rTaFz5OO2A1H3ol28kUC3pye/d
5V66WMweut/HE0ORn3z96/3HoX+jtFJi7LwecVWGHCuDR8yZj/tN4aFxmhLk1Qjv
LqdJOFVI1y5HKWLzVMRb/SsIEfeJku68zBgFbCYNqxRUGZo/SdmA8xHsHUbA+A2W
G+NiP8/X8G0YehOmP7eUK2brjYpWVrtAuIkcCm4L16OIb4ILUr1hwjlDNBbn6uA9
tkUIpnYwB8V9ORQBek9pB3HIJZ5LnwLazcjUqis2lhItNDRSoCVysx2gTW4I4F1+
LF+QK6esZWjaZApfi7Xi9MWsNmfsGDnhcFSxjgOYlwO/+NaJEs2i2FE16f6xkybx
HUZFAU8lQnY41ZizzW8oS9fRnu+hkO8QVWd+iy+u1VjfUUSI3n9Ogfa+VqU+UXDl
KKEcU0kEyi8U3rUQZl4SMuK4E0fgVQA6fZNKl8iXNI2i8gWXsXt+2oXXJ8PD+tMb
fH7IXhgxxa8qItcIctdrcbSc5FX0v7xc40xB61Hqz2XiWHd4vUuJ7utjK9X4A34l
BLWpaG/DjjOm6ZVgRpEQxT3f3Nn/xr0JWBCAfV3PA6t6hgbN5n+5CUn1IvY4pkcT
Cj3GMeDgsF/GqpUWgmq6bBp30lSNgyJ3KUSvDBfBKQtpaRHsBqQ0aYGD8bYM+1sU
OzsOJomra+Ll8OxbUXJ8y41cj4qGXjP3uQ6vYv6upehvG//7oy0O745qqzX978Iq
uqmrVe/7T9fQgMGRFUthAW9Fhp6Lu5r6zZKSzWLYlgHgjabIcFAhiLIcvcTCBrrP
waohxYRLuXU3mvu2weBAybNoHuMnPK9BdgGEgfcNM9birH2V64S/OHJXmAihKrOf
6bWC1l3MzVxhoJG0rWWq85pdUEz5urcfwJUs0mbEqXDyKxGhBlzXuP3vXt/7C5xz
l4jmhVshQeWmGdSL2AdnLvv2SRmVGCwjcX4kLDhSzbBJgQ9J1f0C2rQFHahJfnNz
HcHjyy6vtHTcx/2lAl2MK9EeqUHDKY+5p0WvVuH3s1PPbSKL3oifoIr0C+m9+iq/
vBm+ABFDxwzpMf9CHHYcMrQ58rdYoNd5V0EwZy9NsMB62YEIvcBJz5qkfNRiblKj
eDfHmlYQkCmcL7jqVWmisqJ/NG3TJ7q6VY/d3ay7nPtag0XtMQuBT/wlNhxAaNJ5
/FyZslSMDzUj54ERZSyd6746eAh/cp/5LaSyBVw4SXnMu3t2zmXMpsoS0poCeAyU
8EBH55Lv30/xTsJ6C3sGYEOiIpu1OTvqE7Ui9OIt2LkgJWqOpxgBQK4GiIrbYKWe
sMmVMSklFTo6BolTXqAFqhmQbXW90aTrzHHD8tKsb2CfjjLGytOdz2xYPFOi1ywb
aNH2M/XaYH9ImaxvW7RC1rrI9Zf9ukz5wWThZOk+Rz1jIpBHwTucvdfcCF5N4qyo
z9Ssd5OJ/ME9Z11Fyisf2/M4PAyiuYsApQMjAFllHLOXCn+ZK2/lWb1yGha/HQ92
ORZSTtLOtTXdZ4HMJ+HvO4Kguc8bukEjHuxJfBzKheyszqz5ldQYVPUde1Rt2TnB
H765IYOv4WZrnW/4yHo614XamK/EK7Cn/2QKtSBAdMCj34FvsJvkOF5FvPtzuiiJ
vQ9hbYIA6NtdlzRESB7Nhe3uKEbR54ZNkUhH8O2/VypYIuCl4Wqm02SJDiTJpkZE
Ppbl8WrD7/EzImnSE/hxK1ak0yVg5rVwbS79hwqObkkrSc+NNQwU6/+etyGofMIb
1Ij8VttlsnWR2bFUcjKJCPpyt5kvweHHydJbTS5+ZPCGb7kXx6XDNl1e1TEgmzQN
M+8uDHP7iMOIF5zRYSYppNbbXEZugPeA+YdB/cFLuxMHd34jiLmD0TqStJo8jZ0y
36taEHcysSBS54QwzewhCH6OT9VCwMaOopa7XtEy9/TWtgRhXuiRk0+VSePYv16F
zBQSCS67g9t7bqIrcdp9Z0lb9rUZc+sC8KnPnF36VMlWzSPWXF193Gx+H8kWCvdn
awr87+6gymBNDDlA8l8C8o1foCM7XJh0dPZtyoCna2uuKz6Mgchg8utud+L8agoo
GF6/Ua32msggaBQaSf/a/5wOX5vRMrvPWICDgiCeyikyACKOb3emrcxf9g4JfJ2a
X6fhpweqVj20Bewe20+fzduVMDSDfJiJvVenrcjM3L6RGH9tey7X0Teci26fWQ03
VjK5GHlAMTq4yqS97P/I2o2znJiaOeq1Zc7J1fA0F9tqBFbFYVe9VE6DYMQIhrRN
wfKrL4hGIZO0WV+/M2ORWmiDHQpn+8jYUVVOKjww5xwd8nQ1GFPjFgwFyi8mOskd
oLg57q9aUmzV5rU3V0el4vTU09HmzYcpE8c7ZoeJMhWlIhpw8PkPQ/3iYpDog08h
8KaqCg6QcxsXXjfDYzOssINbfHuVhNZ+nqL/XpRA2ELYZGjGvMCE7ET2/wUYiFZg
x0KgGIoNNzAJg0B7xtVhrv9uVvdKArFF6t2u7d/WpucWqt6h1VyQoAhHpUAIoOD3
6E3ac6FIb1yIu0bJRB6/pguOMNvoUzDq1ZjkzqHuf1FOmC0ig47hK8canAz5/jfk
9/KHuY8R6AQ7PqU76GdOm5Mns+ML/64y5djRxJ7B65RRNTcdP4LT29ce8e9/ETL9
+jta7KR1c+VNXI68EImMgnCCFZ9hFIlwVmtqqmOTqpCgrgmu2J0LvuYGPISOGxJS
fnXqGRjRetnDROl1cpluoMlJ80nFPavWqowF5HF9ck6zVjar7evS61gKdjfKMLod
Z4sN/Dv5lvwwZbw+CURL/w5sp+/RfrmYkt3yb4HBFeOKWH5aVLGFWsu1Xc7mmwyn
Bv0hj72cW17OhGwl2EDvvVlZRZ62iFpQppTV5eFdtsnpazyR6JscHwq7DeFP7e3p
Rbgo5EJ1Tn5FATmnLYhLX4vZSVt69TnJCw7J09vlEK0WiQrTPH1sTx2rpDEZtvMZ
YudsLv2FboQXi16/01zpFgzwCu2BZIAzsFlFNuBh4RqyNqyk3gnT2l26ffyonPvc
6omcDxbVDj5DKTG30abtRLt4z+z/uwOi6aR07v/z8QH2pJiwxSuTpzhEN28Ss97b
lXdduoQbU4CsAB9pyageG2iXY5Pf6MYR3JNpoGfg3EABZEFJDDBLYI6INCkqS6wH
nUb6prfCrVbYbT8KyQ/3Svg2qUrwXe8seFpPmNONMzJdc4EaRD8x2R8Iza6NGLlw
zRQY0TvS+BaFKtz2kCOmq9njmSZROL/cPy3JLInsrOzGGIYTSY4iOkAeXigumfBs
SiHQo7chVD3q9Wyf02axLwm5B2naWpz69rlkrRVbRdRxbwG1iR6hiT54mHvtfRK9
mpBwWZ6Id6VYmztQtNvryDHxA9vOr8U8rU+U1wRQS3tJqFoPBThV7yX3wxwEDMyk
eGnd2mH6JpF7yN69Vna8QX8U2i0Bj/vWK0JJyF4Q1njd6ViUoxR2HQLyxbgB2d9c
yCSjJVSNrIxGmeU3H1BzwiSYIf+ysirktA0elQolrbQUtJPykfnleyHTeVPNDMkV
EG/J8Z5bqEi6UvhxkJ5Z7dNjAfrV7K0kdP9+Ln3NsRnKpn/RDwsucVRulpd95yDH
EyTaGCc5axa3xpt5nRX42T+IWOTFA/HX/wtxtBkSn3eMlhGNlAEsOrXZe4ADU75+
Q/C3viDiBxFcoDG1wMZiw5E6s25oSyyr4R/EaKIEAIcdlf8vPIDxd8pdtZzIo/e8
6aDibYnyxU7z91fSZu+WDmZOIjzMYUFHj1HDBUAxv3lP6c1Nme3msan/2iNCDdN8
DNKuUKuXUcjH2VQlyTRflnrLQ1KcPQDPP8ro7W40NUxmFHyCTHzEXMik3K6s1MAP
+YwOmqloX+U3H0FoMzPi6nvhNnjA2lLrPGwMK5IYN20zUrvhsqPVVBEANJuxx7eV
BJD6zYt3JpiLjM7dSdQMKul5Cl3OQz3z8MVEVSSqy4vTW/XDTP+SD8VU7KNNq+63
tDt2eEIQu5MNJc59501JZOHPeawRSgh+tdt1cS932xVIcyIqSIBH8CyUCacKTw6F
lFRwKLPpMRgHj8J65mAGbJBYOKUOHHGeXHQF3mFsdH2o/aF0332tCKILGR9+f7Zn
pYo5H4z7nNHf89CZmZdebzC8Z9GDAQ2+UlEXuMG2i/u19q1MAGHAq7dUbTKKbeyo
xaOv9C8N1OGpI7gWOwGJGjFEZQrMudmD20LOkRTle5BNMakZeUqhyjfcsDYVFGOi
jTq9fqubITDKGygkNG7PmzY3cxKh/TOqcsUXfqH5jmjub8Jc5MsVdATveRb662Xn
lMIXWY1fN6sEZOKBcPWbYsA0+pDaWslLjc2HHp7AwHACqRPInmmxhZqS40i/lo2c
ojoQXlJDZ3vrpp4lufO1Dqq1BO1dGVJ8cSbaoHjUYrTuKAuVCzoLfPAYq0VgBzFI
H9Pcz8B1Ds+7SYp+HQcAsOadr1kZenOexKzc1259hjZBG2+toljnjkS51s3RD1W6
gfES9GS8QVryqOtemT4UNUdty+G6+Goal7ARCMtwkcfE4/zMcEB5nEA4PbCWMd6G
6bT2BTH0/EriB8FoEk/pzi4akpKv+GF7shOyrRcYSlrv9Osto7AqjlBvHN30KIVR
LIwcb1zNSflWvfUXU7/+chvTlESD8hJKZI75Mv3tDtSFDo/nvXWy63vlWQ7Q1XOe
GdmxAmE8s7gaVEL5sYnEWU3SfJM8fuRTntcYpoRUiy3MXkP9oTkI/V1+ro6bne5A
BoHp/Gk70BBPxxKJLnCsJL2rIOpPmYXnOsGB+KcXpFjt+4Uk4ALMzDmm+Q28/TSt
PRm5Y3rZ6zhpAjBhYRdg8J8anY6n/qBsraFoyfoyHXJU7bQtYh5Z7mC3+qHtDwHb
gUXTvb3uqLc+tyRyJXFQDrryNdQMPY9XXn7SDA4D4o+CbPjyRdVj6CRxO09hUHcF
xpRvucHMD+1uWzILV3fk1rocd2WZidQzaU1gib981V9lbQyPNhtoFuEHFGfPxrlm
RDUGjMzt5GRlOuCtNJw9ZpmoQbo6mIkTCvp77wLFrkSx+bWmY/C4Wf+HNKKTnnOa
wHQ1+NBsoliWxYX1RQCFvhB3rhwPik8PkcbtXzDRK6/zzg7eLe4Dkf46u/+m73Gs
xfzw/mA09YwD5RewVQPabUz9CljD5h7Nu9s8kJlIg3tFQXo/0dpuVBFtowRni+nC
XuFVaHF3mn/+FgjhAFEHpo64jv2wEkRQzHxSRUzLO3AC+N/VPqyDa8MjkcMXxXd0
SiovbnSPxXKmeng4aeOwv6qx+TFF5jAve2rjde1vAkRq2BDH9s1wrlccxs3Oa879
yZRLZk8d5ilMavyU7XLxF/qAq5Scykh6DsZW3MyvsAJ3f1X5g/Amolqr2pWjSNDT
GosnkCK9NiCB93Mf//Nks65Z1v16Gr7RF/Ie70ZBx9HNqlMPnaTtPtXglvHUuZ7i
6umZK+Q346W9YCVU6eDed5Mljws8IyPWbUnJYXBonHjgWLmmyByGe9aCa4IvouKJ
mtv7W36QFLQgyJD04mT7nHVBPrgRYNvnKSMkMTOi5umtCQdWl3zpPUWTsLd1hkOK
ROhiSoNyMSPs2YwII87foOyXRVvUpOZs8Mqq/tkVzmxlv3XYLuDicV87hxJ16U23
S+gNRzGp9nItEaM6+x8Lov0uXo9aB8xhlYLlBCJOgPjDWN2mOSwgXDV6bvE4GeOX
yrRxxrlOdf3phvGtxVHyR8IifAZc/JzRt63E691yV/ASnblO4a9ACL/KBwWrcjW7
tc9IYm0QHiwlP7oqINR3v9CQoxY6+2WaxUTW7K3hIf1Srdou0GbGiCEC5B8tZdMX
sNAfNdrODcfFxVJdyCLNvWs8O18PLg4NLhcovWmufWymQtruufDkJHhk946jFOEK
lGDWM+6r2mxyQGeGmpEgQGv7dJGZQD9/+MLOBZDIEWPHXBu/UcGcEQAJtWDv52Pu
wci/4NYbjfht2pNvFShaNPUamVsGaQyE9N5tmmEBFsBGONohVN4sg0zDIUqMMOjJ
DwPYTlh5owJRHsHF2SPG1TKXzHpWHTPmyPPfQLxuNs60dbmF9DkHE6WAJjOZNRY1
JRYCnFQIpfFMFCDSBovPriLEHpGnLa+y9gXdl08OUxBpvZsPm1N7WFsxZiDHuS98
JLCbZDg3hWzyvpO22mK02xDqjbpTmS7CegzxVI9nBtA28ktewpHkg69fgUp9UGWX
zv0kC6ruqsjsEH4sdcCbcZcdAyVp7LS1BwiQjvWp77+uMs+h74PMefSwba20Qs3B
kYGU74WiJINvzM3vZ0Zpn9Qlxxi/LqYf9P6v+Rwh8EHtAqCgYha+AeMeAgacMrDO
0dESDEJN1bZoOiQpxpwbKDfkdlz+nqkubxG0wOlAbuXs0YN/rJ96o1KhL2TNRlad
cfpi4YqeGhn0u8JxLyTuxMFrZ4m1FZrGTyaiqlBePWiDqJGoPbvnYOdptjgUE3YS
64dJo5/1+DH3Rdk7xWCmf9XLXkN1OACrR1ERmJlK8cHOUQ49izDAMfYgu31cIPxR
IqiGpjuzkRYdSLfvQO5/CfkHEXBZesGcAVCSoH3sc2bVyyWCJpvWcIlgIi2wvWgF
0WSqFKZAjncbMYgjulmKOR5w3l/VJIF2OAtQZLT9SI0vlPYOqFSzu/vnD562z9qz
8v00G/z9CdMLYqNcmbW63raGM+x2UDt9A0ZYA39suuSwfCEseMPYihmdeqqDb1TJ
ehikxYRkqqaE5lDFbt6A0F1BZ4xHc9AGPCz0Lg9CYNnXzPYl6CYSbJkgbMOXmWJi
YjCUTreNwP+QU2JNT+ZCDam7TfU+/nC3i/xfRBlRvhU4zbr+ZmoPHkJTNvxGLtjn
fld03vHlllFaZ4VXTDCeGGGrv83UXtpQCBlHe3qaQOpJT1xtssEH+DWQCOJtUcBJ
okj7sLyXBjqY2w2Gw8IyH0+3nPhUpsre0aUhV7Qyt6tjr5OhxbPYBIwPtx8/sOJb
+YAorHFx0HWrWtCHaPudcdYB+5Q+SDkDWzoafvwOAOoZ+cZUqLfPyEjH04j1dx8U
dhvJP6hhZu9phocKPgylnXwteNHz/E0+zx6zyKQXXGr8OD+7HlYWeJ0aAzuQZcpC
C0f8QnwWt4L/cn6X2v/Hmi0ACYCSHkuEBfpkXtSUgprLmSJELuuuRxHkNBrcSxDq
OoyefNxD6vgkVJdYvR5AWXap8wUebCxGqmaX/Oz1Qoinn96iE+K7CPOsjVqAlwHA
KXR60WZzwGs828zwoEKSQvDSjv8Q8PqXkzUyb5KcR/70Dz4SQRaQIbpeMqzri+sF
vkGux9XVf0aDVdmDnBAZbcrJnFdeEsrSzrf1Ai57E8r9H/AubIqB5p1s719E/yiC
+RCau1eR9muRKiGEinv1Z2unWPljloCG4UtPb0KxhForVYC4yDnMF7G5cdWcgXTb
E3Ew/rIe4ke4cCQcJU8ulWYG831if0666Vw/8aiQHeNb+ijVDb7YSJtCWESIAreL
Qo428Bv8ZrgGnfPHqk9/rHKubcQKzJ2eXWue7da7vIMH+42ZriGgh52eHFnW1CES
hGYViyx6HJ3T4ISE6W3cv69IBgO2UD1DKSYmpPYL7BKB+7Jw098qD36a2AY5uEa9
KSwwBnHuQM6H4j2z8Qi1a3fDyxqfegxEiKS0FdJbBXZmbEw+pI16f/69n7I33sk1
UUJUvsTizuudd16msjQphkyN1X6wiesoBGfFa599MT0vfPZUWLsICLSyksxTKEow
to/8xmS/aZkmpO7NzodadGZ/ZVjrTxFZq93ov2D8mwC2fZ37xJcXRsADMF3yqnp9
X7ton3gw7zzLjdHPmuSoPF3V0my3gNiG+gUHpKSMEYxTl/3cNd/Y57yKNGVFyB6K
HoCxhVlUpRtpENtgrAisYwzjnDyeAh75R3IVugT7lSrfsegRLeSlT6KkEOIGLJa3
WNln4eeT6yCxXLUiQIUE26WfWtdgyRX48c4X2n/QIRJyNHMJCbz5p0a/lPhXnqV1
VMST3H0ik2iyTexewWtLXvY0jmJhjTzA9ibwONOi3uCxcY1n9u2HL5heFtYN/BdA
DsWXQICYgMlzxbVc8t9+2yjVyAo2EVmYqxsWG3oTOQ5JX4wm58gbzZ1b1AXttGWD
STQWsZ06eqq9exrToc7xHjItG/5A/jYWO4U4MH75OO4/cgt/E1fer8/TGX6PS9ph
8P9YWmjBOeK1Zw8KAq1oplLISxRUhcUWtJebIGbc+Ly7VVLvSyZaMEg74vatgSJr
ua7iVdGjUSyW/MsIivwFoyg6s6xLfXXSlnhOoK5Tx7DCj2g92ivuJwy+SK4xSCET
+BtaFITDwtRuw1zO22HgtZwtThmILuXp2EbdqW6HNOxyx9X6IP4k4jFBzolQ70WF
+hPmRjVmH+n8wVnPig1ieRvibrFwJpmdPduvYdoOdGKYRLi1qBnsqfYrc2zV2foA
3VpdZoxVqC0OFgO3+cabNYjulJt+qaIRl8PyRia46x/E4CKh22T96UVFzYfUpXug
q8A0yElHyTvXHTHhY+8QJdxsAbhqD35eVJoUPN2wIOODfqCdDjoUDLL4N7NBOVvC
aKbo01lbAlkB4NrPHPk5IACY/Y7tUBY7gzzccp3J/7bYJ36AJG+dmns50nWdz4B/
AF6TTF6Qz/pOVuXoHgS9Npst9vHwN7OScfnOaVyOcOeDWAfSkjijUVf5fKxNSQ9J
cJ/dpipv4gxhNDQ+K90GBAeg3IdQI64bXtyx+iadAkTAiO8f6IKoLoKfMRPOPiGx
V41rJ42ZnBpsdY+ZXEib3dELsUwMy1EhUcR/T1iaS+mwHK6plAK1UJ/li717Eyd2
nnZqQu/7SGPOV5hfrJf+0mBfwPTGPRqEYIMWVxDQn8LByRKv/SdTYWB5OEGYDbHj
l+D3Gyi/zDRY2Rg0Z556B5E9hoiA4IQJ/2a9Q98qdiJjzGa+YXoMc4Xl0ncEF+IZ
Wvhwy/juySP8N6UiElsRtqTd7hKImuMf7uWZPrnWQj2JJoS3uIMJP396HH4RNs/Y
r6PHsF9t2LsXl2f4gXHXKPak9+Sg9B0V8DQfJulSBtEx3TYkl/QoOefX23zNLrcU
SnLFadZTnD0f7uJ+TcYRHZ58oQbkprUzykYsWd03xvqhofGJJyTKuqC0CDJdEfQg
SEnF9FPaExQeSRenreUha1npcbrEMCRRxinYo91pgNklZs7bTbfu8DxKkQywmo13
nfbmcRS95/5GZAVebNQB9o1XYXG32gncSRTyEmIXNiQ3w/NRN6TvJ+e9tbK98BId
Us+5UMJtfl7gNoGH8VnUqmIj2Q1oFb3DNk0M3sX5GKsxB4dsZ+x+SWCLDqcrJUsC
LG0bHdsYJolp01LuNU/iMs1epHs66xviwuhb4ANfL52rZPlhW/MQVmZnOIMK5miw
I6mFmkHz20Jvq69NMYR5lWEF2ep2mGXNxU6okqBkYdfAB87CvOxpNrfLXsDfNa+p
p52J6zg3xGSF18XE5HQH/1zJ7HVjLeoRJJqxQS/yjKaQ7928A9VOhYwzLMUHxRcL
n3Erwj2wkOfBZSWOXB+GpPySKOruNXeDvsAD1zluWCFM1MFVIwGMj6ub7I5CLa/V
bEg90G8NtJJQ4JV1rdcrJqb7yB/R4aP2568aVu3P3vRT79yiZ/+tg4hzwMI5tsO6
evBi3GvRPpNuaBzgpS0kC8RDu07Sj/IToKXvYsY2SMvOOH0xjFDNQ9XAlA/aDI3u
2Ux4hx8lUn/HXqYrj42UieZiIRe6Ou8n+AGu5lnom/pgmmhQygwVKRe16+vr49qK
pNrzbXLlNyjF7YYJstLdV0Yzo/rgC9NQ3JiiZhuT0eT21MEtSUd2Q7eqfSog+p1E
pjqtMTki1SdS29IHhJH7c176nVSNWtCWDz52+R+UkXrqlOII++dqNGwoJ1rQCn1I
jjpE4ZJEsLFH8XpjI57f3r9c8cqgiaAO54PqGCsmR7BRjx3pO77BR5KJietVAZ9q
izEAK407GR1EgMFTNciKr8QkZQYrIkRjY09JhGY/4avlklNVcr/v4Au6pYy8lm3d
9Xw8ZOgw9/Vh6TNoAQu9hqi3yz6aRdjkEtmGY+3K9WiPlKFUA6ykHXvsaY2Pxys2
BIn+SaC9C+6FAHmM4xGn5qJRJqB5llqon1fj9Kx4wPC6Idf4dYsGq7YLBK6JPC7Y
DdVbD/MYQ53qSsF0Py/Ero80BxHVhQDK1KsniBCQw+b6I2RziwzUI5xiBxZMyMex
nTqnAFJ0TRthIyCHEAkx6viL/Eb2zSroeyA1sUUOtm89J53MrOxLnkrYIivH40wn
wC+oo7ShhmvLIaTw0IQxdRqZVQ/dVtlTAtvQbBLIAU6vDwxUyizPqgNal4y0d+7w
UwQgt96aOpLuLoJSmg4h2ieSJFZgAX6cGUuwWN8E+bV5l/iDtR9iCSPud7WX4m7y
JpBQF73Utv57+m5kucDuvrZfzjdpwJYLy0VXIIvlOWkuzJfctAaAK2gfjSoZwe1Y
m6oWtL7wBIuZUAAoo1yV2vokwGTNJDpm6zgjPsy/ytxZkPgC1sBuhYJ8cfrlAkrg
YKF0XHfyvSAdCnZQBLc4s9eIs9kEH8Mkf6wv+bs2DCasNg9IDZ/nzKiljOI9YPJY
6FMHAmBxf0DA8ecfs9nf9F0vQpALlWNDnfI1DCOtbK/6QfpSBZ/HIJNLLKB69iHs
0BobJMaWBo8Hm6ug2/9myH9Bi60n5KeUmTga3JGHbBFhvfjjDDLPsCb4GSeu/9fV
tOOovoGnabQvLzW6jCPfSRXIcpjcduLgwyHv2zYTv28PzO0kga+pCM02NIu06HlS
9z2LCeVgI5oOEvY1vYo5B1FpP9j8Ar07MqwcnMsjXhA2Dz6CLIviXk2Vep3KT92k
htwyPeWMM025GePk8qBXcEPtAZl5otIoGyBBReNPxbmtAFmhyqIUxsNXR/c8H2TD
xNUZeA4fJ2DOrhxVD6F1sbrTF2NiNoQ3kCqXHoDPbBLwJIjIw95D61BHkfeUMqj6
MfV0QipPuruYLuJG1ws7ba3s5zk2JF0IIcI7zLD/GttQkIAuGGdhQxibCcSeSTjg
N40AGlsNuz8xGcpisP8vzhKLDwjvNncei5c9NmEQKl4JjRJjo4nU282trZM099Jn
WGDZw/TIvPTrcZjy8JmF0dyzKVvAEJb3p/YZBIFIo5B3PgMcTol50Wydm30C2PuR
uZtVDSDYWYGqbvqhVNtGRm6GtqdQo7Los06desXZD5wPy8ClmiOh8xZUfwFMFsHH
/NlvsLHLPJP0EmUkjYQCzOT2GMvajxhcWUC5mGWfpOH29OZmjR+nYJGIpnAXuXGp
Z1ks9qnDrG/vdiAM5ecthBYNBYN37u7iV/jI+wEn3YKZdZh176LrEhmbwkIuEkAu
akws6+U0rjXWk5Syl6XXhRdjwnDtWNn/G9BXDlWHy7H41zj4HtscO4yXRMbKqN9u
v/cRpx/BpL0J9Y3ah9CukO6mQioa2X6USzZitlTocAqillftU2b2ca4MWXMFVWyU
f1DISpW8cyhKIFJs6CVdsCdB3KleOREbYmw3fhrBkWMmU1TRfkpdu+2gogqsL9g/
vcgMcDOWk0xRK/czthX5Nqcj/Eqs68tJ7fPvBwTIZNf3vGZxc4UvejNm1Te96V7U
1pG5jO8IqOqM2QFzPrqmOyFBQ2aaRk4Ij8eI1ixpzdhVke+udU16/apVuF3p7agU
jxerONmYu0crMVINP0jLbDzwRq5YmlCQUIc13cb+6lmSkCwpdQRG27W8g5yI3DXY
Wysy2rQrNdTAufe273vLadCCWy99honfjEb2qqWa14OAUDtj/734+PNnyyCPPN3U
NSNKex/Poe3KCKX6E5qNh89qXRaO8ln1mgLlI8RA3JQh+q+BN1MJIuYxWpUhlpzn
1ftFW3ztkikUOut17GzAYvAa6WgZyqrC2a7Zp+9HEdokjNofg+c6z3lHYq0RP5nP
6IXqghH8JhZlKQHafM9+KzYLVUlWVte7eyZNZ2hWU7+Gt9AsBDxrsbkvuRTANG24
cT5ECjsyWGJBmrx3WcVc65f536dV+z10eTsv6/PQmyY5GREHEAYFsXX65VoNxxHJ
suaZ1rP+scWyhEPKSeut1w5+jorFGMj3QSRCezljuyiGfDDK6fKEUp0k8B9TR33w
ZDczUrm1ppMRU9oR4+0FHXK9Wv8jksAJicB1jr+HvKOlVYF9csawKzw3/rnsqbB/
hlqZEU9dXLcPtRng1gPKEsRLKnuDfHN8RBSWboHp+uDe+fZnuAPCFb0GoJlECdFa
vuPFEDA83ROu4Ne2fjGjfuLGlSOKQIcPcrJJ03kBBcJIGybYSlRdKdNGZnTD4sv0
EXAdrTuYXVn22+IHSRYTXW4bA4TaWxWhQltWXho7Ir2TnCEQsOzMjdEMQexJyHTJ
i+5r45loCIEvjY4hmMrluGgkHWQDx6bXXBqbonHPJkpuzzljShuZKoRjtawtWjof
BAQWauiLPZTqZPlMjIPYUFceDkKKNzlqkr8V+Iky6VO5ZF1aLVdHXumxGYIVqlkC
SjcQ8QG2cfBRazPcfntaiASQm9zMm2ogYuSeSRVv04VIJwG1oXwtlM5J9T67XSdC
9dMA9NZhllrLkXcIHcaevaTi7Q1x6igQlulC02z58s7TBW/nBjK7s1Cx0kr4LFNL
nhKY7JOptUQh/BreNOJmjNAMZp5cWH6E02sx5AfVW0uUPz/yvw5v0hOA2KDMa3a2
FdypBsd5WhG5CKboD2ryPBIbU4dZ27VZHiX8IGUqT60G7bKveeo0w8EWt7tkahzw
z8uSColJMGc1k6ZV6sLqputjRuMG/I3RKAhdVQvApj/pQNfcCDLftlXZSOLXEEwc
idH+NDitbMLcfiLuDEpMF4JzSIdHa4WzF61P88rNK04ee9PDNdt8M8Yj/JpJ3Sws
CFyoy8nxbnZlCt2lZ0EZZ45RBP9CZB1TCksGiMNHpziQAukGlbV8KZNAdW1tQCk6
eTzqFd8bGlhJqdAunmJnjQUBV5ge82K5TlymHJmmd7hf2hyc/7aSsUkR6i+nxsrX
T5sEXyHxydw1bORKB4eNlsJiHXg/+Sq94RHp4kCdSuGW99/IL99PuhFd+ZTAhi3K
8Z7QfkU1YwcKyf4Yae4Zqd98btr5mF8TcZK/m9cxhPRsSoX4sQQ5pcLLvctwz2Pz
t59xyw5+sNDT/0d8ye5PoFM5Pk2H4XeiL+POf9NhJujTwAwsRy82nviVFI4wVKW2
CTxoa3JsYar6ZokgjL/3bXXnD9DFSICdjaQaI6pqt7dpzxX6Ho3vCDQBZoWit0Tg
LrGL1oU0IcYxUkKUO4FEHSyz3rNKxCjiaOO84uxrVt2F3PZqkg9AGHQTJY6Dkhq9
kptwh9nOCLN0xerDYTPdHqd55zIi/RbZQJCLF78WG3sYsms2PGATc7ZHXOPeaQKQ
e79j4EdQuOOLJn3FKQ6yauUPZFL2BHSmiwEEYFlKeyg/tBlRtPMbIfd28lAHkskp
25skaMiHvzwSisvaTJmuXkLZNl37UJvP4hYJM1SNoi6gu5dQd/W8hu1sG8pyY8S3
7KPE6FJCLT8FUgj0ALB7obP6i7WGmfymEL14ErSXj/aiNzkMjVevDENSkaPwjll/
f8TpNP47/RBiKrF+QL0iin2rUgqgIJr4j/nA1wBfdmOtCwZ+GipR0gg7USSg49nm
IYG5rJXrr3cjHzz99rEvz8bOp4wz0LTAVxqiuJGrGt5u7w9B15o1JhzCpBhWqlcu
1K/d60AkLzfllBTemihu5M4UgIMFEJOuomPo6tKu23gfCclUowZEHxjsgwuykC/y
MGXMcVverBtGZiCY13R84mzjf22TMwzpVi/ABFBJSOh2WYa/nP93Te8p42MQyFOe
jTI+GwMqr/LWC4Lx3nh+KzPN3seFOTuu3jI7MLrQglFbrZrYkEycumfa3iKlDle6
D1wVNh3KLcpYa4Q3cAVbxMMdVwZs6V/JRhYfRYGDLah/wlR9v9rQua2QSSUpGoym
9NoKKwqHkwzkp7wLnlt5wVaWajqiB4+nDA5KouKUySsUPOkfWEO64uSI3t5fovfh
1HH+/1LQt2sLy6VKMJpUbIcTwAF0o33hC+DekavOmBVihWYfdPSlkM4VKsi9ZVGy
Vawmti/RSZ20pBnCUJEIVEDYHx4HOLrfEEnezIzWd9l1AiHJ8H4yeuvN3MFhiIHR
nrYbNa+DE7T1f7jBOgftpAvGV3hEomzfcQf9VE0kVT2NvcBXib8x6o3c9Sc+lhjs
lNckkdflv3LIkzRFP6YsqT6Z/AejmbLqJmbcBhAQOarPwUIMYKy8RlLkG9GNloDn
bjnxXoVO1JiipvysoK8AC8ks8q2nc0QZ1yG3ceDImFiP9I9fVGLObBASRq046whv
JOMLXBkwS/6KHQgK4qh+5S27v057FqhIkwz74VE86LakbTjxXrGzmBhvnKdCMRTz
Hd1c9a7QH/ZyfWnE4VUs4P0Z004IPr2f6Gx1AxztfBojAEZUXn3OQ5ZyPrKLQiaW
z7j84q0xYXMhUg40jzTRhbUr3EdbyFLTx/BTSE3Rmmd1J1n5Pzm9ypYNBXJIWWrk
/J/ssB+LdCl1AsTVmQFv34qJIVoI/lyidbGxaU9b7gFWuZsLtiTKS9uPFgow7+fZ
h8ujSKwedk85zEccZ6sGQ2HgzI8KyhMyVC8zyDw3duLTavcDpzK2Geb+qgo4bB8c
k08ecODutozYJMr/QthrOvQQ4nu07YSA/nonVo1zm2CXpjh9ehy2HtW6J1jKv259
4a12k4uAhIHUGuG/jUl27OUvUU48oB03/ndN2RQaW0YEz/lEMLNhtGEU2ovE59AO
UXK/kqTJdJP6iBp1BGTKTmY4KPe9gN+QvJdAVKng+m8LAZtP5pEWv7Ds+MCJHQgx
tfJh6gQj5jA9lRwRtqWknbXRZrR9jdXVxuBcw5+i3nzs+uKZnoavkBf5Cy/AjHNr
cUU/hmrbHJuLrbZKRm4fXQ/SG7/LSWAjzE0fgf9ihveJbScH2KiJByAfcpgmIk3v
ruyCZSfFkN/2v5OreMtciAJnjW5iUTQK3rh3k9HDAC8sFuy0JC5+BLF0VzF9GdC2
lmdXlxGlGMtC0OcXcUSuTzyraEK8aA2mxYs0ExVVdYu+no7cvXTi3Fw6haRC0jfR
N2AGl5vXlTrkzEJcVHl92XwmOefj3WbCZzHfJvCFmlO6dVk2mmIbiSFWuuCrV48N
sk+dtAhTtuXjIEw8O8boiTfSC3l10JB2FOlCnkp0vkmV3L1/NazGssNOX4vsKe5A
MpXIDWsCj/o3XYwZflX1i/6nYIg1qL+9jnnI6VKnABJu/SV3CMzOI95VnNSqVh+S
r0oM5FHVyYlEQVfDcEakQDtwLimgCxU60Zl2kXcE/IJ37nDFZg/+AG2JX1BcnD2L
FQbb6S+u+Lqroi+S4xXCyZd6k7cm/yDT8fL9sFZcWmdKPKYuvM+lQ1OsqgTPSOfv
+9c+bTxQ0XR8U/DCaWhexdUAm6bO2KVRTg4BtIb4qfsJXw7HvaFgvgL+xmLPkHXn
ITdOJG+bDfnRBfYZa6ql0tPeZEJjVZW7v7O8ul2MyK9P4mjs9U3uP9RAaCvblMWe
eK4PgEN2c6qsHtUSJEhcAY0XCwpAA9PxSpVESgVI/+Wm7WtyRdx8dJRTJJAGyw/M
CfPC+BlsXNBIIPUWFWc0v1LMITO5+3BtnHBM78Cg3H2pdNllSEqab5vP6MGX9mf2
YBiHKPXPziPSq024sVW6Pdzppz75E98RLK0VE9qYuEDS4UT2pNAzm8gdS7pWR4hK
eij9okOmZRLSj676aTeQoMIC/FJ8mS6/KHylI5y/sfrXlwAPyamhOXoqmj+3gpQ6
mp/jdqmFiRKea5yfLX85Srp6fS4fUrM4CiS+aKB8iqbpbUgjX+jfmnKjUA6g1iEt
OMAhpSEtSvLIE+lw3/o3bQbP5n8+Af37AAaGpy01BnCed7rWYtROE5FEU/H3TeZs
64y38trfDi1vw3QoBcA82QEfvw9b8TG//FhajI4YL+LbvqP6yqiamLHke8L6lCmZ
he0s4DYm/PmpeHCHhKHoq9OtTWjFpTPsBENExrp2fBBnWNW/BcON1D6ZSnWGLNvw
bJ7iXY2BUOeXMLSdG1uJKkb7vnXdecWQMSQtYqa1W5wT9+QTXBKh8uoHed39SQ08
CfkVkpjatsSam8pEdwk9KoVikkKBvn8m9BguUkK5AuFEaY127uGwlTCe9jTOEdGN
QsqRgMPNCDoXJHP9WnNeJwbBSYx/P95g7ydvLAMOE95rEWDAlPnaaEaLLMfMc2M1
wjra53ql12KAH65CWlzSP/RH2ozVkmXJbaxwATNAPYjodxstMSX/Ij1iHgDlMG8N
r+K20ACdG+G4goYLjBfachgBQkpbv66UHiukdzyWOcsOCfCLvNziCJFlJ05mmQpl
bPK0UKjFl+oxKG7wv94catBg3aWSOjT2z/dv0ztVJ6gagQKh4YHiM2ufJ13EZ7/N
ukzLITUXtdD9asFS9mLmx+XQ8utZNTvofiI83aempXH/Hn/q9F/uqh3UFkn3x/5i
QGx9w3ZhMURzVSW0YJIl7h8kLJ4pwjgv242JZtvkQSKanlYtF8tDrki0ocQEQsXh
dMe1Yq82h1/hxbj9f7tmr80hZEhCgqI7M8AIaBHIm8RYqk5bHYMLTd+yZrIUbXdP
ir1ut0lDI4ofa55BjTGykAwgE/DJZ3sp9ezx6e/i/OXTbCq585425cbkMsCcbbi9
S7Lo/ZlKnIoCJ7lATlqL5mYEmc6Rb7dU75CwlM7lmBJM4zBy3ecz550qGzsWpvc0
xnlmkMOitShJ77TePJ106gj4aeEm6piM4p6Y6nQR8W6xDHM6Oo1BqSfc5UTp7Bkm
8Jof7yic5JoEp/F4IMibX9vs4t69nK+f+VB15aVbnbBlzMy7ZyzQwvyhHDEoIyWl
ipNED77sX3Rh1tZlL5ro4FD3hqtlPoW4hd7o09DL/3cKtXrPnU+ewrPx4xeTeGCp
WZffIbTitFHtGqbJSCk4CjtLo3KxCXmODAJ4NlpHqE3XGMnhFBZl4EfcZHbjss17
TL7/sA5pH5lFhoi8/fTS1H0wgDfUpqyEzs4jUFKvok2TCqjUvHrvXX0nO5XaMkgz
YshMwnV5Nsjoba26CY5+eoIhhD94OCe7YpWA47gQLsADA7/ATVFIHhGzZvGjESp+
7fUHq1CuqNE0tZsJ/Yj7dAKi6PflJvXDkq3a4XfZzjBNew2XThhx9yXrmWLCcJAX
s8He2hgJlTbox5ak7BEBoRnwip/1dE7/nMSFkvq2zSMbbxMz9C5yAR1cdhDp6oTD
eThC6A7TAKsnQpUNeH2Y3MzcO4di02Te0t0YONgkPS9mn+9o37y64AEadZLO1RZ+
Hw1YlWPYTW2sgjApTNSJDPfGsXF4ta+IMHjZuGWQK4d1a/XMUbw6D9nFcSQ1SXCv
R23f34AQvZ9p6Ev8RtR3uhSJQMsZC4fR8yYKG/T/R10KcQrm3din266lyPtWGXhD
IWJEfVzD3+WY8fly+PXvUCF91xKE2bx/L2kvq8F5eN8hZdn3yndU4Es8MMnO8SlQ
QsjX5JmuSSETXUMIIhkgpb83MIrbRyhOXrkj4lxu5/RwAT7kiDr8np6igcXMLgRK
`protect end_protected