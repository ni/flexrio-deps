`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15664 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRmRy9l4xs0tB8DLo+i6+lxmZYzbZylZkJdfpQ1QH318T
WITs12S2znaVMaxiQ0esp/5qpHDSskDhRML5GRAKcX03Uru6RpHzVdPatAHyk7kL
x8wSRsPVMUtHHA4MbLFxv+fsDiyG73muxsr7klH5KGX96jVapDQji9xjBz4RlZbf
mWD2nmbhabHcSguet6jujNTg4uqLzbBhAWqFPeM0q886CCt5vgYwZeqTPow3Nz20
d/6zx02nyLN6s4sciR9JH0clp5cRTzqJvszaCghpNuXQmR1DY+BLFga1352oO3RI
k7duAKhgRkVgWF8gE1uqzJAIeiRL6ls+2nIzt4nWyR55vcxBd/y4qUKULiGhDOAP
nA8dkywRVZ0UWgJ4SsbGzOLDC7PT6ZH7qL0cpC832nKadcRHqn3qT6AHIaNpiW6+
ExFGT/WK4n3ut47MFmv4UVcHYBcauWXltfQfvRZQQj+1IXIpS6jFcPnEa6GuJDfJ
5WoG6OlHylf+iTBNVLi1zLCCKcEbrUX9TlKBflP1h7EZjDvJpquWSrfbAWYhUdDp
vhS6t0CnhZE9ysQnDh4TGGTCqjLptCiDQwBvS+zkQvDWosIV5AUfKeAasN6qQCmY
LOnc2+1JZlweJ1HQk3VeOwIm++3Lu2aG7/KQLQb/pF+3XiVmZJdaIrcOgm8iw6UF
HFYegTQXyn9xUFqlxFQ4kZdAggDeUHNZw93aO3l4si3lYgTmSNZ5SaozA5wkuG+6
okifOfbDmc7wLUZ30yaohDDa8JSkrTsvsz9GA8NsOk/vQ07jZum8OQioQCNPm0qp
MRDeJTgZdDxZuVdXz5XfuQQ/g5/JG01KusYaIYdY/lkjOo30K38y5zrCpA0jMvOn
tf+wGXqYfxq8YWsYLZ6LI/iaBVrDWvXq+LgOsD54JDltoUhUKASlAN+lfO6xHmKx
nS8Wv1kWQqUAXTYwSTPGTvGrO3WeTeBWgIK6l+KOy2p7sexFQGLGaPNJivOX7mpg
8VCKLggopdLHgywA7iV1huJwJvCJSD7FxODYspIUGVhpSJtHYW1/fK008y2pK0hw
eWwCY5X/eCgb7meMUvArNi74tRRn9d10foGpkKCqtBYfdBoFodZldWASGxtLzjM4
meGjxZc4lJTOOvyvaj3NDMbENVQwzKGSDaQoa/ya80X9oUfsuUF/Olpi084WIzqT
qwSWGKAVrd7zZYZKKLYvMB4xhpwztfiEIpbJ8TIgbaP7xTPn7o/r6iM1rGSX2DI+
beyR2mroNnL8LwAFFHM6fklyqHxwkGt1LiXW7QrmmJe+NoTGSOZAlksQu38rN3gI
PcqRBjVRQcKpHWaWqrzizq3xNOYLfpXEYY6Gzn9k8s775yPRyVomnubOx9HUi/3z
GduyB9GX8v9iFuKj2nUaBtUpPO4TW4sn3HrkTzE+53qMFf5suM70KGK8h3/2nJC1
NYz3gFPG4PS7pcs4mtoHSix8MTmGh4te7Uv47Os0SeB9gvtNCsEEYB5Hs8UHzwh7
SCg+2OHNac2cqnL0jgY5Xa4Y2WhSOiIphHfFu5S1e20AIBidv08bEK+h+pPD0iSs
pwLAArpLjuL4SBlPw1NRmlNKFaBsiwg1kKIpyBKg21zs+I1eT0iNm+GnZ5K4YQ9Z
UGQUl9SfXGfcy+ys0gAhiHYjNczkHok7Oy2Fo5Cff7yKtpp3uaigWyRMND+7abMf
KIBY1mjIY/d2dXSuabpOvMKinRivte4bifvug+jRPapcH1SIHbii1B8NQd01Hcg7
BnBzvm7ImHidrtE2UCINiSyhRvcSwwgeCMAB+bdNh0GHwbyrTUqe92MX8xGLP1hM
aQMfptJsSwtAy2waM1ZpArj5yM2dPe92nvzSQkt4DBSS3zVQol0da/pvEruV3t+z
XFN6BkdpYbuqfNpsIB+/26co++puQbXNsFHRvsqhOAvRFCQkHNFwlOhtkejmSoHR
uRVEZ+u17xl2auhbAhnVhXs4zrqY9gj5/Gfl075EWeSovZVmxB4XUmpvbrTQtG+o
jFa28uJA8aBcZ7XPv1FJFAE0xVIcJvy4afTwg3pkCTWq+5lqD3b+CiGqwlPiJ98f
50dL5r/TK6WWz9H417kqBQZIKxo5tX1tCQRc0O3BZ+9Qwjh8VfooX18p2ZU+/WQM
e66vA95td+JJ/q8zD/GN9aY+hGpAak1xV3ad/HiyMlvBdmGu0D9mUHjtCuPseKzi
0Tr+wnFK3h6b57NXq1q1PY+t4QqgwjVbfkBv7cApEcUb6wCgLLHSqE7vrchZLev/
z0U1pobCHjBKx9/KGJHPmZ9u6K0V70q+2isMQUDWbgwInwmxtLxXk5JaFYAH0TXh
SWDwZvZ1h08TJT7fUW1yAiuykPRNz/5NeY9IcpOsKAlQ1r6H5cYvneMJiuLMCg5f
2z1ifvoYHjrcl6XluN8c6O6eHQjVsOkXI87abiYqlebQv7BV+UfBBv1zI7uXpXzv
l81k08TDB4d3hxXNE1ybIHR6sfP3SxOI3W4fr3wHh+tNeWi0gJF+Oj6HTiXlaqE9
P4LECrxtaush9jh8lIw4AEWjvJz/Jg6PyaQRFs78fqbFDr2LBwVHRMnJluH/qKjx
ShNcICvGcFAIXhecmo8GqcPeUFv674rhRkA7ZkZRINRssn2Rqlmc7ff0rcnzfeK5
8EogcFq2CNkB7+0fPt/5MjNgKj+czPVetgfxR2VxDuOEB5u4OpvcVf5b4AvVFgfx
qjjkv6nvACFfujN2o9OH2CeohE3Qq34mHOtmVJeMYGn1fZuaV9A80wc3RyhKb3k9
fBoyGXkl7dWVEBTaongnfWsxuR0mpNxl/OqrpGHqzXhVqIiOUYsD1uv4ETxaGTwR
7K531cDwBQHYj0LOG87gbntXGm6ls3W+tpzv+9dBJhY6clF8TPllkxePDkyha2kr
tPpcTWigYjlotLhyoip26zmUybyq1ewJOsYyV8SywcLXOX4/ckH4QLZhsiX/scgj
8hpvWuJmbdb6w+3MmoRktLWj+BRX6NmJN+5TmqVlHX5XCUQIPUl7vnrLNvrR21Oi
mte8SjMWbu8/N2oj39MNnMDR86dvddT05aiIZwSlRAtYcoRZpmrKddHm0hoIJAZ9
q327a9isI84fffZCa2iSOA4JTJyRoPm+kDBTTFijsA9APQ2HXMnugEwgfC3/tetq
UZpP1ghqehrloKMZdqHTPRG2KwKc3RDag1xIHZrFHQelZ2CZNnVg0N9XNJhoQoMM
NicSd/JMy9uSBp/V1bGRXmW3S8hA1j+jmZh6oKcdaTmFKA2Ur7oQALro93tlL7R8
TrpKflxV7dFLoCBOX9jZgig7n6TfucMu5+yWf7mWVD87YxBFyCYSlM4h3cgk9cjo
yFquhG4pjL0nSdFUVgaxESzovyMeMkNAazwterp5iF3/p3atQZpRZTaxCVyTva50
I7LLVhVO0gZpYhj8TpCfL3j8/alGfCbcrDNobBXE+Zcq20Wj0fl0fcwA7QqYyunU
FivzNNQm0OjJvhczmW5kYE2r5oaWO/fyFmvATyAqtKVm+mi336ZMqFsTkIBcrBWU
a5OQOoinfnN/bV1uoiItSX6wvqN8YMY06xGq+/8qISpBShQqpL9W2PsSWpmQdjMa
upCg06m5J4uenEpZ04J89DY6BUC6Lm5qPtrOW76rgu0iIUnVM7cYhr/I5V718UXK
Hwc83MY2KbgyHKbbyBOK13Op8n4znjQdhHwBkbORwUqHQ5QZcas52UXgDWfqi9KK
WmwoKsWyvR5lGy12TDPkd5hOU32vHmIkoxguie1Ky3frlTQXEUBYYxKumSQErh+m
AZq2UjOXk6hxiIZEZb5z7z4uxC5nHODqSiGTW5qXAtEI8cM4W0Pvk/Wjs6eFRDAy
vc/OHAaBFQ0u9XNq3ywPyF3r+cmNdVWoJSARZnoyaZBhy2Cn5sDS3pwMsJUemh7S
+BjqmkWC0r4Y+K77IVxgc5WbhxqAnM7ROClmvlNSZBIrTcv0r0xK+i4nxNYUbPk1
3aVJkR4vUpFFbN3PxT0T8NpyvHScyGsOo0xP6BE7vB+7VYt1LdeQIVhk83Z6G6rc
B11sYl8cRyQf3qAPyaPWWO8Lt9fMt+zeMntzeh/yqDjL2RfHCDZZ5ZiofeEMO1vQ
Sx07Gia3cYsUErAkTCsXsH4ITuXBiqYVGu6dpNC3fZb9r1yPCkqFG8NwECnoZ/FA
tE6iDb/XP0uRfkCHPCBVaZT0MS822LPPDB3lQIwF6kXl7bJGUn9BMhq+U5BGnOTa
m9LAtkiiPSmu4W46Ss1bHjFJHLUPzAJwf2hEz8+23X3NcvcCu1CMELcF+AXSZL62
VkJOOk/zATSKYEpS1GfO0FHzJzWfk/AyKg3N8FGeLIvcmNe6ir7FOYVycJRWKWUX
+LaoYdXlsq+knZ6l+DJlZm2piJ+X9fZZ0Q+hMjncO226zkQ1TgPCcB1YRHUgaIon
scDOlb3FiFWmYAlUvoQhwFiT8ugdMHSCChpzFdQvHfGh9nl6stXkks5WhKucLj6E
kYhxa7QgMxTAKvXWjefoufTUF6E1e5pFVneBOysLbE2Z4bm3ta4dcKSTuv0cEZ5y
wOVGZU8cA66comQLkTnS5T9/mTWyyMf7qzBFExzXXBPEKneeIeJyW7odh1TOt5yp
rC6cTJQL/8F36tg5edVdqVZejtCgaFL7b2CZSC/AlDXlVSo+FfGBWxmRnkEkt01E
fPq7qEtuZLOYbAglTYDMYcaxSuSHPh14hZwWfzedEG6ODkR5mSDwowi02DLEL6f4
6MUrRcHDDOM/bWH72PxJSWsZRw4D3v9dC6XOYyuDcEUXc3PHSLft0HIJ9QO06UDZ
gEIPp/ud6S9cTEfD8/mjiCVIFT07SzSBWkPNq60xK4yGVYTa/18dZBXQs+JS9/aE
6qI3FamCB7eTl8ybVQtl53aDSqOm3xmXsfyPGBw78SW0u3vXhV4tWbE7g1pWdYmY
vmQIO9E6hyiJgCoAS8RUvDvffqqSS79JNOxkuHm8lIC5qv32paL2ZCN60v0mAiXV
X81kg5qEvI2uT6NFSq7H8t4g0OIbbKa9YDceqSb/nUHiaV9yqtUAP3OYbA+4HF44
pyh4nkCDklMRZyOMDbXDdCXa0ZXdROkZFo/LF+FnB9VHAuXqARcejG20oPQKJWm8
vztGKmahocEV/skyBId+I/u1rtAYTlRF8PJrTEJR+L7IGnchLtpe5UD1ptmy2Gkw
NFhD+8LDVqSed0u1wgvTJdWTJ/t1IpbKHr3whpY0wnmzDLzxHHAgm3yBC3wxjkNy
qQ5ONclJIrtUboQ6xWFuJD8ufgDARAqQTkEIr5XUs557BSI+7l0WTxvWbwzKiKO8
DhagyrHLQ5gmPdZmTzftwuXX9oAYkoZluyDAsgUgaKMzCqJMFQ1Y7HiYI4vCooIi
lU3cLig8+C5bYyXS2Ssr63FqlWuyaNvpdNORXdjC2O1qqqdUD+3cK6w674FxtzE8
j4v+Mp26Y4jVpXA8poDGwT6fJGkFXMMmjT8CDoIKw87I9SWZpwBgffM8dhji07ZV
mL8ZlQxo7UmmUy++6LqRMoKWvWw27N0/hBwLy6HSW2lvd9ii4XJg0nuEOrqJo1Wf
ORu1Z1DRWVBQinsjF6vERVNA/7CQTtRZOVmMhMMqv0JHvPYw7M/2WvD7KxIhCdt5
yJJ7uyEQkBeVV+V4+RrSwnQ0oDIUbSDcIC5gAFg4RGm5wJf2v1S0wy9nm/ZveaGV
Jn2CFdxE748crYn5VkkrOkLadFtsUPo0hvccv0FE1XozGtAdnzYRO25Ryu4C3RNe
e7aPVZFqNzBJ3e29pB7njOnzBzsWwu+mPQ5aLpkP81kGSsmAF2I8zyA2CqbME2OF
HsIfKaKvVNhonUu6ZaCqDRG1VWfyiFYrVkEGaA+KXTYDAZEhrCKWgA+yURBEUCq8
41ub2RSL/PYIqrvsVsa3wDofHa3MF1KMCna/X8twjTe6vK5jAlmoltp3fBz0fQgs
dDoS8q1dbVcQmhY4Q1GwtHniAulkWUpOi3GMTH5XXgkRPgoTxYkN5KnCbMytuN7i
Q1mQW5yFec4uqz9UOsnFn6NIaAPs4ul/JhCWPO6zmIs6Snwcp75SXuj6deGDGb9T
LfEBn/A6raE1lRSU7ffOPG9BHXuLyr5Fe4MM5llSU5D/VCMTAMth0CSXL6xRtkF9
aUlC1aRao7oZosZ6wk+HMVO9vhSH9xirg6iTsYFl7Jjiw0RWBOm7I+f/K+30v0rg
xheWGICib3sL07hnDK69tHMHUbD8se/3LtBNQdjpz0o3jwioXhNIH2ieH8wRwAgU
Q6mfdAUrbVpc8D8elhFS77yF8cSjDkKLLzjmLCGTzXUTsvET7n4ZlUvo9bMCOFnu
447PPnmbczvg1cH747rXD8U1IknuZGTDD+BJJWcCqwMcDdBM99ir5OGKpyRLsSUu
8e5tQmkY4hvj4/JRuUWdjH51c9zF9rve+lCmB+MclPc+dHiEG6IfNNmeIb+HFfQ/
C6I9DSnzpQYCINORQFoSvs74oyco1zYCN/iUsExvU0y28jx/YrwV9+OIdkEES8Jd
XjubFb6dSk+z3iGd/byZBQ7SXfNx+6/mZRtnx2h55H6JB1iTaUUBsOkYPM2fm9UD
dPjT5Y5tu+b2NSzmPIIJBlmhSR/mvcHInwzUii4V3TrQV2ajbpscFlXGKc/kdAa6
cDP76dKlI7rSWqN2fjX54OuvRe5ntvVJUZcQGbcM1XqdKS87S8pZbpl5EvKKpqkb
Y1B9jeQRaXcpGz2dzeCdTUL46rMzFPywhGcPUQA5KIE3C4SW7p0G1VqGce3/mwW5
9mPPJLp2cV0jNZEbT0Dkm2sr9ExJzvlssUagcX6Tb1rxgmsbEgUDdFzJnfpMSf3B
WQZ44bL3alD9DEwxIKweDv8Zsda4D7maV9P0hCGuYTb4rHJFtaPmgU6i50C41NwP
vVlFFfPw9dSOaJzMiJ27fqbEWk8hCtpLBK71JGqb3Fqf46eI54z815x9GGwbvIZb
m25YqnLv743rJWpRJCV6kf/N8AP95fCfGTe3HrlJdsOgrDfBMTBuB9nr5OiqszKn
ckqVXv8t+eyIar8zx9cRWRtklcuvhS8ybE0oLpJDvcJdKtVFosUaWLBSwzxMEvE9
2/gkXxukjigZ7JVS9bExynNTgeEU1baSRcJ+Zq40ViZp/MutPaVGHZyKuvcatUnr
sn9bNgZuG7hHFKiqXr2GFgYSVfbn1qPEoSzSjfjqFuN99Mt4vwOpfOA5jN8v08wR
OdQ/4K4aNTPHRmvCMPSgIBsk4p9wj0wmw3KmE2uVIddip7RAD+rx0TW94hU8Wdor
55VYu0N+12XW6xYvK2gfgkKdMqhg15MTWnFWfCuwVjRAQVV0gmXNXOGE283NwRcA
dmPvnWb4fgiVScFNPkU1Hq9yidsHExc4blSXWfiOpO+PIAtJRb68Rru9u2HLP8RL
9fKmx43WTFq8/7KV1qMM5SxMtN3LpGUJaDKcktF5eILHLQo4ZMs5MQCogLjyLtFH
aXVGS2f+ALj84Ks2ygEXHqMjDDoW5oV0g5LtjQ2C4JUwOg35U0GGKJllIZtfbN/N
NNcgbe79+SlLYADv7IOeX/oBT5m6EG1yNwYGL8uuY+98tPZpsqCMnBPWhXun2+l2
UbL+RO15kZoewA6Apo99lJajfUTKAiuj/GfONAzMJHQD1J1+fwhwBEp4Ud07Zdwk
nkjizEaGZ6uWZcxpG4vWtXvx65wHWDjbfec03F5X62LLvaYGsFR1ByPHMJk1IKV3
z0d4etWpg9SOrbMnWKIFBmf902nJKy6+arnXZFp8T/FKJdlSk/ghW6oQL4B8QDpw
ztQeKWCKZEpaTs1Q4iHxgn+nEm02PAp0b4P6vTv05FTirz6B+467R5leUal634Bg
ObxyVVDDNZOkjsd2d6QOxkevHNkw1/Bc0kyTQSpBuql+ph99dy/IHkb1qZ1FR0E0
Mgc8hJdJa/60fS4v0+RGKCtdLpj0983PcMB7OKfs1MtEJTyWU5hDHkrQcy8joCGC
MYkUNO6ZxuZIyHecqwv5aRVQDSe7A3oOoFQwy9edgdSmidzRsYhtBHs9m+jEUhnR
BLGZdq+rFWOxTmLa9VMaVoHqOeBz3xHSK1bOT/K2a5YHTrlQB+Yl9Pmd0gvCWJ3m
sNHZ/C/82UL0YKyit4dsOd6QRFWhYOgUk7A+Uga2qdqfdV0qf6dmj/RAB42ELs9/
NS2oo9/2s8gd5w+ttNvP0qvqNdJHhxuUy7BSHQb8Cz/rYCW4LwLH09uVFGGDO52b
96o5LZy9H+1kug2roiMXeMJgEWH0lV2/DUZx9ztX80XWqEkTh2FyWWNt3/Aq+VAO
CySO9dn1Hd5b44KeARMVsB1g/TVs9UMMckMULrrEuG4Zg/YosZG8NytruQj0N6m/
y+TY7jb1uDDhp3BKuafdfoH7DhbJm7Jq+bBiqotKH+ExBoZUHH6voKTn5ryR/S6O
drFK4+DMLr49Y/R9FZ8u3dWSShqKFDYBhRyOnfLCClFuW4PBTJxCRKJNOiBmCDaw
CGNnI8wZ5XAVGkmdWs+4wsX+g8mBP33HMBnhDZKrK3JO6v7ljJmMWKfzPKRyQOZE
ddOrTPlBp5b2oet+Sh/ALVYAg2rUo+IrvBzIfYiI5S0Tu39tjnoTpdLN3ee941km
wujXB2XQWHaDPQK0wgFOPnC8rV9V4+I36+Es3jmMtzqsGtE2dJr0Ixrha18E9lRP
YejWk6BuzWV0fKfqIq/GjH5A9esr+8fCKBsNgLsJMGZNgJE50vk76TkfhnxJL9bp
EcNDICWT1bndkFw8DcS9dWs/YA06tOjeyDuf/SwK8l4rvy0otfxPcAGdVpNK7q48
RUIPaVM1aJvNSpUg/QT1tTR7aiVlXXGlyRCwnCiR8tWJ8rgpB+kgqKixjK9kDPky
8D3PGTW2tAgWxapKKXK783cO3V1JZbxksTcF2jP7UjAhFMAVleST2mGD/9qvA/am
J2TP4NAxbWmj69k6knZecbUe6M7+zvFslZz0zL2ruaZErt0+oQnCMCZ5XAt5bxY4
tpuxb4POROOUy8VwvWRJp+t5MWCqLfjgq77fjrrLmC5HgqBwLMmiTDMoFiwKPfaO
qox0mnmVT2WAyd95XWb6XfS9S23ZL/Z3YYxa4CVVl5aakstGLFkD0xfx3eThf8UD
bjti9ZQk1YF4ZV6G0AxEPZBInBJLLkFsH3/KGz8z4gIZNpJNVJ1zS+esqI2/HmSV
TWO9PNxjbFsL/8R65im9oYcJRRilF37dAMBJBgmDMa7PvNzkNCkYKFfX8hxTVKQb
alfx/lfL7n4w96S3TPiOmEY9f+eyAZQ9WFA7hhu2MOEP750e2fZyO1DkVCtaE6RJ
uZAHmuantOb8ykXzUUkgV4hCOhqb4qr3H9XSSy8TgMon0ednG4cxoKqWgdgO38dq
2QimZWEBKgzWYkkyYwN26SUFU1Lulp93xmDMQ8Z6Bw5zSnbXC3Q9TTWom1s39FqX
Kcf2+/Zve0k9hfgDERG+avIseP4f4E2NGN74Bq3gZAKdC8TWwx+VY4GDR+sSl5UK
XS+QbM6LcNbOExGCC2ZwibXBMloAFZeHZS1F37OSAGdXDVZAgLz+nFe4AbQQUz8a
rRnWhsu3YImCLA1UvyQxpbC2ZcZb/ihvQbxlr4I0+koVnB1NzOqaub6C9d86yzQT
72m+066ux17YOGvHDGXLp1QhkT0j4hl8f6694qd42EDkMaWDl5QeYTWhsbCDSPpR
E7jy1b9zdJUdZUU32m2Y/zgpm9zU1OxGkCWMJhcExqtIEcPRgawXTRIPxPVK6LnA
xgTUCq9S20b4jQpLKnVHvIGX3UxY/3f+7/dQh8xEKvHhghFUUGYlrVqtaAKBxa4a
UTMNGKBPmMhZlLrdfZE4owhbcw5eH1IfjfM7MRKqh3+bW5yMTFckw6Ys+9U8b233
8oqfH1m5MRxN5WnZ8uRqQiGSvfRto2ZWSWcskoroxS2eBDZLcO1OClo157INJZzd
cvh1g35G7ztZCGxBOE4MjQvOGgz3Fyk4Uk+oChNOyUXdvUn0KZWQOu7Alf4S1Xug
XSpwPiRLZTA/gSJp9pU7hLCy4YEYkvynR5GWpoNrSkTu+laTwObF69u7+jJudSEi
VKF44vGOc0xPB3cc4Urj0TfDOJdS0FeVgbuyX38+INs7YTO0iopddT28p+yHrPSl
23xvJAM2G9wSkYYNADoInVH0f0FImUtfvoX/SnhuCUnCkfaFPh85Zwn6eaQrFGOz
PsFx3+oZWsiu8hIZj/f9tYcd6OhmN3r6oirtNjpLXN7cBXkHJZkJpxPl2Zz49l6T
snS838KpE9nl3yGHAcJ5ViQHNZdllyygnDgSE7/PToePxMYvfHmpI3f3u1deO208
vT/m+rcll1GRRaKkx5l4aLrVS7LsXW+pQtobxPnoqhzuXYb13an/dwhCTzVRb0N9
ZBYV+6QasxIthJZzDN1/yPhSOwwRbIq+lkSAQi4niC2tp4TSbPi4FGuczDlRm7Td
ezBMVR/SUV600aBc9+oRvUkaJRJGFb3ltIGCL4MIZpBziRBPJdkHfVQPAUjImYOI
dURaox+SKPogpw9fgtm+v0ygE1/gu8oxXVU+fvnN4OXLvrxSBVBSW7l0Q3PVOE/X
Q8Hsc8Fa2MYetcZZm7Y+/8KhpDJgRBEd7knl86a52V89Mzb7KYv/ofnqUl5ygof8
xWnG4yu4vAEcQWpc3wXcJM8rCX8JGpCRnCvXnDXvfCSo/YSA9h+v4+WbIAnml9hB
tUYnmWI/TUHMdUFRE2XExOqtPP6uwicUIKWu7JMWPU7os7QiFQaeYi9vsMqY63wo
RXc5jwdv5lGn3+0wFJCFexCSZgkDD82aNTVeYJbEd9+/xCFrABzGZ2u/Kd+OBBNW
okUg9Atrzr4lRWcR3ny/pmbWOaBFsQBiPNhgB7oPYwbHOIBocdZhgtaNmoAKNO5E
6+U2vsDzsmspdxrgSg/HzZFZkQ53XxkiQ4ak5orCPg9uzAe5AY+e0CWlFJa4yonU
5o9IYZAxWbX1WIF+x136xtRsEJcq6nxGUdTgdncEVCWAqmMo3LqaMTRM4xqWTtLJ
1CSbfATyM37yGKicNjjH2JHNvU5boB4Vp4h0C2RWPo3N4kP3jfadeN/ILYlx/YOv
4+oWBXAFSj2CHpb050qptoGT3vOttfup+vFqN/v1wmw/6+gk88mhz1Yk6YOxn5jo
uK5e+QvF/Dha/YUopehxF5Lil5rf2WDSlnVWQ3bItZv8e4CIPJQqYSQFG9ClkJLP
ccRXiYsIVbvBWbVusvJjARNwG7OsQfTKiYneTvp9A6Q9Ny7TPcqqy20ZKchkFmsD
nhC6HCl8fVMCOzq5/xxrTsPd/XoxML/IxtrzBJX6ky4u/24H5jhmVYSDBklskbgU
JmtTE235K/K3xyQANfi1czGxiKxTZh8zBLyEJgOgaoIQEfVW7Jbx90aRYqIPx6rq
7emKpaI4pV0hcD9VcpuWNh4pFx2T9ka/ZxCosO3ZIDvALzV5/f/zo/nZLvq1qCBo
YqLjEhOjRWoZh31Il7K86ZcxddzzvUwKCeEeaQkUA0nKMzDoNR7DfscvTcLr1EgT
6NqIHPFkfwYcXlKfkzYLYWNyehT1MBaRvR9qOtYhduIncBKnzkP1lP3V9DTiatsr
cIscdXweBHN15J9b30HyTFLCQQNo3niLSpxZb8FOjZ8h+BdqNoh0PxoKkuqLWaUJ
30ZER3lneJ0v9vgv2oXR/17AF+Yg7fQoD6cZMxVn3usUyE+BdcSJYTuHJF7ayF7H
mLzzcV4DabqDfaEbPY6j4tDLLUgyk1jaAR3nr2+/lYaJP9hNyckV7e6iA+q8fPJ/
UbTS9LZbZf/MyZh5e8+yX/fxCCpOPwkulyu2j5nkItoMcUl8QrU538y6sH8NW2HT
MDCtXfUbtPRw3afI3/ciXZ5YfBGtpCTgPqRlL+RXrh8FKKyo49r6vtSTDrV6YoMv
9hmcGROSLeD0r4lYodYb4XZ71w1pGlQDPRNG6IGcebFUeauFpQSoG6Fw4RqSI+//
noL1kF1gD3f0pD2z7qdB1fecxPqMgxkCKh5pUmP74UHN/HiDnhu+RmAHp9ekFXiH
5Lt/37G5aLoer8dC6yfYQJR3kMh6zW2e72D+NeHa/czc6K5nPX+MADPsLjUbs/vH
euM5d5kkMj9l8E4h9Qgy8QOtd93dUXDa/BgBAdg6ozXKO+2M50dRiABUx3x0bAbJ
/0QFtw7P3o4ob4FJpCwz4HIafPHZSFMn7dTMgb2Pf7C8JYZEIQEaXLxUsQAi9ME/
Fr2PN0/nDg0J6GHg9gEszt682MHdNbX7BM5AmEmL9dxikjk/6bwasI3LJkr9J9dP
vrnuVChpdwfY/bAjTKUmLLsP6QPbRlz+DImhjMNHUQnPh8JLVzI08/gdY4zf0+wN
itDuY9XJuKXUMprhQhR9jMe/DfPpQ40ZQl+wR+GeS3O2lxR+T3LceJzjEqCWK2ZD
s1uIfd207DcIjo8HwGH7wk1XCGhsQFe0pDm3FJihSWEfORUpkXsKxEMSKfEkzOPr
lfTuHSAto5Oo1RkjWmivFj5IpPhUqEBT2kdh+v8uXZGnIINYYy+wg/DPHFuzayL2
B/9DbtujSQ6k+xCc8OmCnPYY4V1tbjTk+9iQ/wp06Z0qo9YPaug4cEkk8YffokPU
sV4wqsCTttavfLeg9s8ulDP3XEu1juBynBPFzAPNL31LC6nBj8QqhqYi/KvKoDdf
I/66aRnVph/CvMmy1u38S1DHrNm4gvTCT0Vm4YmJtoBHbSUxCK9TPLZ+Yzo1+RqP
sqnn898kuPlrXZxRqMg1dgGVQ8hu7QkZZizUWydKOI5y0L1F8L11L/v86P+l7wOS
FDIGQfo/8DT/ZBW4koZGBbF/AkzLnmfbgPNXG/EWlLr98bAz62IJVWEQXmtZo9dm
9u/19GErL0t0x/dCcX028qx/2L7W/qpbPGG7UBm3RWH0aW+21tqxwa0Pdx/oUns5
8/qX/oeAajQMPU6PUtw5tkS2OMy3H+XA2A8QGPL4P2yEMVFeXTnSyUrqDbpl+QbO
GNo2trJeAB1s0/LSk+fmLBsjLEzT3o5V4l9FoScxcqL46mtC+FuW0eTkLfWMsx0f
3R06Rdm1FbS9aCDExgMTSrHj3KBJdE6FvdyLR7DOmKWeIYpTQIrjrCX739EpwKNb
0W+omRIzlC8iqk7+8jPNeJv3P1z6wmuzNYe9+1EeigBGkwgEiTYarhaOacsktlyg
8HOZEXfYoXfSQK3jyNpGf3pUiexg/Rbjkjj29ToA/M7E14CoQtksOK3RC9Mg5W+j
F+p9yrmAnW1co1nk3br4oAxl5zUxSEKglz9ocmEQn9OmRPh1tAbOr7lWYeC6i5yw
TCE5DQyPTITfTTkIh7c5lepAjoAMqPXCl3zsdOhuJBcoj/YFjpStpaUFQmJ88n+Y
WPVACBIncKD7J8/rDUaa1UzBw5C7uY7tZoL+hPO4jjMrbM0ZT2fTJWQ3sqxIkiVA
9FCpJ2JZdkr+qly3RiNdAYKFMuLpRkxC/WnfUrJm567qUJ6dWot/rf5iKj2W7DxC
s7vOugI6iIiw0VNvyXRzctC/FdN4ym2xZTbG4CPlLbtwFLRt1YAwfP5G4ZxrntZW
69ZssXS80bbpmcOHv9MrE9eVAdjhywopNllbo1O/uT+AEYiWIxzzy/QHjlnNaPN9
m7Fg/RDxoLtqqikgOjWr1Is0IQ82PQU63+r+8hqvu0ZyC8pMjq5/XjrB03b+BmOk
XVsxTs+xRicBmXv3Gh+7RmvMotBxpAZioNM5ZW2l+6B9R8jDgcg+eWD85UcTuahj
b8VQVZuCfbMwfXvm91hbwggRMyJLWpAJeabk/iVU8hhMp2OpqJr+z8LI5Til51mW
03rsxuP4EfG+wPWYB5FyjNRUSNdH4uQdGdHQL2h0sqt7urm0Q38TRAKbbS9hvKiO
2lP8MGt9mCDOJIKQULLIctcwU44TczoiIJRnZEBum45+Bjyl+3H+m1yVli01wC9R
mpFEt1pKMSVDRIk0j0ZY4vpFbXDvvWOuR5HycRCubenw1pfomxqlUx2ROdBu8Xzb
5EYDkjfn/fP6wJAqm1oPUgqrQsmLuMjbB1URinwYaFFBcN5rliT5q5dSN3gpPlcf
NAw+DsBrEMg9FLtqFotehPRoLaIyAOlBO7fIPi2bNxiRCok44dNShZzUEyDUEiNM
J7S/ijLaEfdKoUC6cUigTkgyOuIVQ8QzeCjTjbv7NivjTrVnUHFb/tsg5P9v7Jwp
P/+lxo9o4JHxAcqgr4efbhQTJZYNCcnOpWEk++Uben0vI+qlqhg1CxQkxNqYEbdx
hviORWSmRo/5eNa1x22rHcuICaZAU+CGk+KRPUUSW0NNn6mGG8pjP7OUAecRw2O3
kTblGcrclVfuKhXEW+D+8zip384i/7/zUDtJaCXtK+1f/3K/z9gRu9gL1xURs8dY
AxdZRuo/eT8SZKKkA5VTV9ZxDYc5z6IYaI1Gfc31tpyUyI/XRSIsfeDcQAPlGy6b
S4gdgKj7ImHbTMaXSRpiIlR9wPNJnu2PyGznqBKew5nYqqwKASS+tctmVs5Wls2c
e7DDfQvbFApugitU4ejn3bzwSSyJwvJ/j1cv6y7bdBjKLl/VonyKSp0yl5seC+7l
hpR6kvtEUS7VNaWj1ovrB+UHh76mRu/VTYyRajy6qxyjuC+AQ7+52ptkvNWzURd/
N8quYOlWx/FI74OJXapyyc0iD97UPYL3VOpv4fk2z0clEh+J5EPpRA0tVWeROznZ
lh7/pgRobo+/a6gl8QJW7Z/ReAkgnhdptDvxJz2uyjO+BrItNLD40bQq2tT5AfSq
+OZrvsq8WeCr6vSOw34y0ZxqOJI6UU1GuiHnA27Em2412VM5+b4p39C5xosSQeQP
SBEwvb8rUGlq2y59wAaQ1sb/QBon8QSkeFruRdUG428q3nyr8SnSgp7yVETBkd1Z
SDykX+nk5WAw7XP7xjTRCzQjnK+9Ul+x3D6CmP603pPKQUWvdQl933W7ilIASkSW
uHnFmymAYUuzgE1+xlLN4m0H+jOYiZFBDZL0gvl3JZbTSoEmS9nP/OVj/HU1gryk
ciyR3zhZwjq29sls8/KJq3jAhUdlVsMGDynZdj5oSGRueGlcYiXFIupGDD+lz2Yt
uTr/O3njkHsBob0MnNlJPCJIUMURIwuJQtooXZUfTHUrHEYlQagrtp0XPcQ3I8GH
a3aPX9KoGc6p/ihYsCHHyIU+xx8117+bZN0ntNaFiyVECFPk2GMVNaRlaZHDz2wF
Bd5D0cWAVsKO/BvIce/3nwDnCsPlutu2GOu/QiNHaWnHdQUxKElNgrokHR17YbZr
M2bzY+oiQTzwRnqC+7k3RIFynAaiq8H7IeMRoPZvqhgtT2Rq35iYFuYxbpcgUCkN
l5x0Il330P5IjcJP6N6ZqFGu3ZN6XGPLbR/3araChJb9uDQbqjWZDnnnifq8Xkzx
4MasknfBiVRtgiywPtLAAH6eiTSTX7JKNjVpq/+P4qlnJs+UUuw42W0WqGzHX+52
Hr0BNTVSbfBXjMDy1k7E5E1sqqBQDrgGX3tnKYgsb4zvWnBignXUR3MUjZ6xDJ+S
BtuBVfS/RWvrrP2WIdJB+Y0XtKWGg7/4JPojp8nRiEY5G0LNsX//hL9tbDoUofWG
tXdszP+70W+9Y6dx0wDSa1eCzykx6ZJqA9tJmTgyseVSFW1cp26o4LA9AAtaUCvI
cKkqP2tvyRPCUDAaLSI8as27uhzvFKof4EXhcCx0V9yT3bXgB04Opgb2Cpyvdt0b
bx61RMGkeDofTVF9ibiHC+ByE+8Dekz00N2ji1DjSpNTkDOcmiPWp2smXKM5vzqN
uipohbtON/5FOCLB9S8HEbVo3IumPb8oDZQunynLqXy8ekXUzNNn62fdqMVhgjr/
Gc3PKBUMm68Om1zcsiFpJ9qfECcz26AsonO0Y12bxUfue9sjXK7ccD917X6fE+Nx
jZJcOE4tznJXB2OFFy7sCN/mZQqLO6nqDVCvNUONiMWFzVq7Sc9CcB9XV/Weoa7m
CyHTehjpE5iHMv/n9rL2AlwBUbOWsRBUUsM9dxcn6MHPkXXXsXrOmZD7V6ib724x
4o18X3CC11P2ypQQOE0eWWiYCC+++tOcup4nzUlnRQh0Shb4ZhdMfFGmKEkzw9Er
Sb1VCjNuXxF7A3iMNw52gRHLf/NvgUG01aeVHD5Gz0yfWAogwegl6PZk/LxAW/r5
4WMfcEhM1pZ0mK6SANtGj9iWZBKkjosFmQpZpIDO5aarjmddjCHtNvK6L8Ef3jNG
mtHMyV8nXpwaeiZCgNYXGX1eW8GqEAU9vpAdiigpBiI6WOFplFbsdnIJA6LKtUVC
Mmr8ouV8YhtQ3fJ6ascqXdJlA0b9CeFP0gDxuwetRLPimDZBruor+MjNIXn4QGJJ
5R76AXbJjYcmJgHg1/51pgIW23nvTznvdYqyzlbisvPrInsAQtDl/UJwqAtxedbU
X9JySg7zgACXxVhzwjcXgiobcXRVJm2WN1by3UGRNsNEJzgybuf209FBCDUrDvzn
uhN0ejCEuj9BUVSM4YbRkKh+MD23R5HEUmBbYByX7IZRQDYhj8YdQhr0A4UAdfeZ
JPqckACd1m3/EpOSoZUjO60f7qjJh8jqZEQNHDjKJZivtqUnwsI7pZ6/RQTXf20C
fbf8QCZkJx1oS5FuZEYM4MRixeLrtnCdDW7Kf4llu6yqdmwUYRovW9m37AJtKaDB
1UYtVIbAy1XhKc1ornKXmYdzaJA0x+blYdW/kizeZH8aCoMlNP+vskONTRVLTJdK
mfKFrcmoY6ZvXq4SivgocRlA3XPRUaXLf49WwIM6YmSIP2F5k8hxH3HrPe9h8pD2
iyaOR2577BPO6bHCD/EvOtY5DaeYhrF50ZWA5f5S0GvCnQF+9W/p5IBWYsIQbYqz
6AOEdd3vCOOcy2G7VX+5IrPIuS1jXmxDYlQcxYLW8Ty+8S/XeNZ3o/+hpH6Elc/k
4j6LDv9qjkVJCRNzTYqahLp97jfLm210suK9bAZH5Cjt8Q0sUp+q33AUF8BObsAx
za0cTs8NqaDUlk+TD9ynJCvHftySP1DKzAQO3O0VcAfLThNsckRe2dJJ2xNav2qL
HpEEVYpv8mHqjRx7sk4+Y8VD/Zod3p4ubDEx2ZJ1vnPxkK3Tel/F8ZEjmRVnU9EA
z1e6uCHBC7griVO91oQpPY39w7ghL6LhdfjOeYPGGKiFT+HMHsbO0Uku0fSuzszA
Tk6FZauFrPBMslor8S3ohwY7WyOM7rqWYsS55Ls1VMjHwFkf5Og8LLkZyvNtOAf7
7fhr8WstjD4mHDnhb1jwieBD/U6cpx88mOGiobYZD48sBqihi6ESel5cwbWHOoGj
uCo0Y3sVwcRO968opcnzQ0lBcaqBQmtnJOE7uHkHD/qX/rHzWRrJBeB6KjD0chei
P3KQzRpubR4CGm8fG/mshwwwYPkEF0mwZa5/XePuRfk7GkQjXJ9urT3mcwgIGNCa
WemjPgeY5TXbolVtgoF3PJcrbcNtlI7Ug0vobbqqCtkvwaKmzhDIlckVy2zYP43o
cz9b1s9tcvSjF/YXoP+Agu6ywUYqop9ikErZspRJ9TyqlHRyoXDaRj4F5oojY3kA
ZY+h0SiczstKx0BJzTbsbOGEKV/52xLVGwSpYLsVgoHbLcFA0V5A/RfNhqgPV/JV
al+NYhs6FhHkUzdAbqTvHne1ByWfPvk8d2bwQQscpxbxVVrWh71Q+CaaHIMX34+V
xEue7dlPwbEL/kW+x5PgIrcqsTXnH4BeLHolO51vaxf+K8k+awq8790KuIbHkLIu
8ruMxEhhq4Bi+N91UPiWZvNURKO9HRm7Qp20QO0cTcO77KCJa0ez9iEzGFUjrDSr
ZYQOK3kvwo5aI8k9I1RfkfzaxUjhfn7n68MyltdpLtprRr0013DBdybrFPAk1oLZ
1t3tBA+aAdtQ/5eVhpNeGIwwhG8I70aArKl/vXK5vAaR9zcWPRY0NsVoWwl8189J
ehO/o4TsZQ/dV3n0FDOgBFatwpmalNst5xAkWazzaJkHj7e5Iw05+Qah9PqhQH0L
rCYCkJenN/uhOg6j6g5mf7HDU60QzJFMtq72sp3bo7tL0shvkVbO22++nSUEc9Sq
oDucX+0VTy2I83dIJkO/ts/P8pDdH9nBALHC5WaLe0anGrd9PY8FfqBN1Xzk4yut
w0HysO/6O1pnY03mCqdKufKjIJyYu6WTLMBoLaM3TieuO4khL+OANK+5FZtI488W
sQ0eQH0cdKwn/wAwMJn6P/jEoH5MzRFcJmZ866POHtBMvZwPQlHAGB8LYQLI84Lv
arh+ILWrj9Oe1nTIhVhCmO/W/V6/xMT2eBB5YMWS99z9sCn00lr0W2BpzIpI1LRj
2XDay+/KJSzPMTrh8D/NmwFKPAMiAYL5Jtnroq5vbr6uEUBwmIOj2gUtpRnj8qTn
IBiI2T1wmlpIOHkAf4ql3Gl7boqgNq3f48U2k1Kp9L2iXMjYeYa9QpMlQIjdiw6R
EqYW48expT+WXH2kuYXVK5xJ3rUz8ihbTLH4IOZNCPSjDs/b6Bg6srE+y4DpDy6l
LRARUSyNE3xkNxpp6vnxyBZaFuZNUPpJyM0k+z5gJMDZfVKsoF7gzDfG3LoaA+pn
XfhdY6E4fGwDtqK8jPcbr5PscXiCBWafw7vkeWy5D6hJuW3tPdgLz147pVuNETbo
XPHFVPs1Sy2GZri6c5lkQWzu5NRvGHLEATbi7jueyVCx/umV5F34gVEQCmkDtEI0
vuGa7jUEGTh4lijHEeSRaBNOfpDXEOIXnpEiT001gm1N8OugVPiZu/WRJLcrGj3y
rfYRuexMzxGhVXtrHmwWnK++AwyEv5+dmK3yPW9DrmVFjygK3p5F4quNshAH7MUQ
BHDE+Ht9ArZDMxlDPKc2uNPPtPaQMOyCjQgccgtL7j5T1U74ymE/TPMPtICW4Sz1
1wKCdtDhqPXoGpYgZyO2rrBbI68k7uyC82mG1Oeq3+dW9lTv8A1ypMcL0ZRTS08K
A7vggR8gSY67dMHZhyOk6JrifpfdtdsUCQWqntF5ZOrPqteJ5FM6e/4AvdQPIomL
RS7LbAcxvVLWnfnGhaJjolvtIMxiVScSlB6XUDhjwIISovZLcbWkqPrGj2dcRyMs
RZqi5J0GsVp/KHr/6BeoBjhbPrv4eL2ivjjFicWR0AuoVf+DLJJZFSKDeyAZMafx
unxRUUEdIy1slQQc47rXD/NNMpHYT+ph5/VmkvYb71c6XvYtKVeVydVC5/S12cxt
TqNGBq6peMZ5HPVvXSPXH2zeSE+XGM2urulWBnyQBrGl5Os/q+0W8aNvZ7OuSzL6
HZzo8q/BkyAXXP09UVVRaIzKsl9DWt2aZk/J/fzY5bc7ziXAoP5yrFRMxh2WvlM6
5EDkpMPVkOhlGkOoUerp0zdfn2APKXu0+gkkcXEo04OkbDc/UL000AchWvq4hTOX
dAVjdoxBlx9KErg556jzFxgK1Rt6Tqbts5fX4+7FPjR6pRLWf1lBYipU9dLTk7hz
472O8aaij7Kof+YdQZxXWXBOzST9ze2bddkueyrv4+xJZDHS+jt1dOXJty9bxcQp
4Qjo1r0E6zzwTk39fl1AAT6+bCDjhYRJOBXZbh0nKyII3BI35LCmbjxV1KuYcTvT
y2UnUGwNjcOxbn9tWaAQICr/1fK79QF/CP1Jb87avkJ7z/0qQzxMu82h76CAs1qc
2vMmZhQN6uSY5tznEOyJqDlKyBOYOnimBwJ0Z2/Fjy5YE7b36KMdCL8PTGV3jg5N
uEVOHBhnVKNRfik3/TzAcdrgTdBGm+WfePBmqvbd38D6GtXTZz25/8chKJNrAmj1
el2+6ySkfyK2hdqU8REUXhbhl9zAHy5w/TX300lqc8S2PvlNciS04lYh9GHaw46f
Kn7FVMjf60/EUaOjREleQ5Lz30WJdBZEGXgjdkfCCQlmYNsaKWct2pmwwB2HHiN5
5VNFiEkxlbXMgSucVspm7OUlDKOjNg/8edbHAeiVaqRKfhvaPdNMErqN2Q+A1VPE
6JMR+CHjW+vROenjA2NAvn8a1554Hp+qSkeEgqUOMsivIL3sMLpc2SIsInwqw106
RNMOw4GPKPJNXAwuzwkvPp9y4Sunj3wVXLp7W/6qEyT2dibDRmzULrubfGztvJi/
rLMZJ8eqtBEKZFvsFCodByPK+D0/rGeZ+USp5rS52yiQkjmo+Hip1I6WTaobUQmX
bCscFAiWGk1VTnwe+DzMFTVc7JYJ32otLlJEXV15JETvWWHMYG8UUM1nHGmbRRRt
0T0dP2iRDgzHOiHm00BzDMwQt5V5psWkLj8kfs/qaeUMtUAqqsZ6jsxxT9srzAxK
WH9iaoHeSNYCYRbLP3ZCb2PpL5Lb3QaOvSVO0qi467KCPSwayD0C/9TOWkTypxfz
Qaw4uHUtFVROG2fwg+AiUn9GIutuDQX4VKs8eB9XZyum9nik6JOmID9TCAiA9slo
DegAvhO4+Ai4zRXikelwhjclRxwoEAgjS8TqMJxi9MSNsZ3hFAHsXHLzp0oUOMWn
a2xLA0kzLtCVZ0QRKiIJqYtiEoa8RoyYwHoo1oR8OU4/PZukXJyVyHzR8kKsszbY
7fXhfXaZDnR/N0sxHrelTg==
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15664 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aWGCC3/z6KKo1Lc3LUdqKyuw7cmOG+SU046+gUXzDtUu
Wg93nPKw+882cEJThJoh6USXw7ByP1KdSD9Bg6J2nbRw8LHxLqaaxfD1GgnaaxTr
SaWnlHNq2jXtVdVrLxjet3av1ZuG8KmLCsGyPpmWDZbwFkT3yYY2L6bZzx1iTuX+
NYJjxfHBmgSH91+9Jx4P9EYh9bFElDl6nAOVI23lQTlkECAmEtLYE+oQ2IpovDIw
IMOFjBbw8aSJ7dtdG5tDVh78kQjWWsyWftkGzifJTCCPKPRf7uaT2GARHM4bBZmt
wLrFkFFWcdD8XknKsmA/52TouGneajlfOnp+KcNWqwB8b8+l2N5CICgNCpjDD/bE
p2urrPcG0sz961XA9SoTge2VRRHOguDBWS4fPJ0qbhSQH37DlYADNh+ypUvHu9zl
MYc7CMIPuiavcC+/B6QhB399bGKgZGsFHx61cYoatFsqSgFD9S8+lnxXrFtvD+LH
B5NbhSGL5vewYpWlwarsxuweVw9UNt43MMflyJehLifM54O8S++p2ypsECpuXHyv
lscfgLAn3DXPolmf8Ly3osolXCpjaQHA5p3uf9X7//p1JEf3/zK8DYkQ6ova8Zdu
nokCaLlZDWupX97rwGFA8gPqj+7oO1afu2K08dTvEI/XFoVRLf8XXG3TyRxHgfdD
2GpZleOTFql3/ZEna6DI/x3pbsQN9zSdHieuOAmvjyL9p00W3r1SIMj4LTQgL6Nq
nuN0zaw2HMcVj/4flhoDEoLoNWdLJSKpkrRinwUujvad47zDMIlRZpbahF7D/APT
77vBJSykkxcmAUsK8CwrVORUHJtOLhtgX9eStJWjnQ6jIBEJBn/5w4Aq7VkfZcWA
sZAk0QMmEp4k/wFv1jJaVw91uxvjXvjMNErBeBudBieqvkjVH8GQOOUSNpAXgoYQ
WHDo8Q9R3nQK6/Zihp+9EmpJSrn3WdFs0mdSteYbANFczJGSIfbzCsUJoPxAy7WI
EEZah1HXA9rUQwCumLi2aIrtJl3uIEaCum4sqmewgr9E8BMeUtgNTjKQZsHWakG7
AZTwzytgywokZIilou8C7Sdz10dcTmXEwpraJEhFSAAYyIJYyGrAocBWwQxPi6In
dXM5UU68FRxSAxUGT+oy4kMlwoTufbAscb6JoVgPeDWRTNf50cx8riHAhNHiMg07
sixswdq7vX5H7oCFC6Ps8oUjOqKm1PGMY7SfO8DlxdSDLzL+CPMtRIgIAqS67Pgc
nz1wC7rnedVQAxi8QFkMECpKflU8V1quqJ7/bQETfxxSPdc+B9DINalSFQuT57io
0Zlr5MoUSgudiHewU+M3UTeMjVTlnDrsOQVSI77rckkCSvcsqc04qB2/6WgVki1S
D+0Fc2lDFLPQbd8Z66E/myFdPNVtQRL80ipthfVRQYrWKQGBPJmYmlRYwk48bxgk
u/DHrbPghg4wp+ofGb1uWmuq7NtWc998LLhEX1wK5dkdD71fLNESZKoq06w7z0Ke
vLFyOVyEL5wyH7iqfqakbnMU1wHzBrj0wma3xargLjFzNmlAltFeaNzom5BNqLFZ
W8riZphYlYLZC8Eq1ybzOsDqRDpk+2cpfuprHE6ZOb37ffXVz9apiHc9FDN9J9nI
23uNjewodvquqaWu6GGHd3nZFqXSW83cijy+XYsK2Bm3dEqNy+dmHn/NY4aKL0I0
aiB3POBJWYaHheJu24KT/uJwV6Uq4ievO8p2hgkUnDW0d2JDCi3Z+jxMZIEYZhWU
mSzGW7vC3ig6lqonH8HY451jBuZmJQYo9qH4HXWdsjSUQXFAoYYKs8Zl9vHkCWk+
IrLJAjzroSbeckqysaeMYxh7y9KSoD0Xlo22ri3SThrhxbXEX7+OrtmVVl4b4y5B
36P+XO8gsgLOPw3tMc0CAF7GLJfKHsFYUnPtBDVlLZE/GQlVYKrexMIyZwTK4G0U
i0yUcR85Cl0VnD4W5j23/lfmaqLKJhOEUOJUgOoUYU3GLm+thq0goBUZWKDHKS49
9gsgUfKM4bO60QT/ANUQfxld5hT2txaR1NLiK4Xj1c9st9W6W08askuxWgCpZH2k
BAZc8V3P7y4ANXzRz1S6zuBE6QZiNx32mETZDEBlTSioJKjjvMWRcwPCq6VLUa0Q
bzLjSVOZginHshg9siTo4aBAWWf7bJ4R2w8YNwofKs8rq6m6L/xUzXHriz596CVo
jW6pmy0D0v9O3CJ44RccX0jChLlVRjAA1EtU1pfJrgBOIupLFFj8l4BEsQxZi6kg
H03Phpa02LGyUl50lZ3TETDP3u1fCaduRu+SrQw2nJsnmhm9e0jTQpxIQyooc26r
xa6ukJZbon9LvsgdgqtrcFt7On3gA0fRsMjecssgQaOIYlqr87lniY7m9nNTEAbX
XooEkMAK7OOFrazgXjI1FFJJnDH/H5Hef/AtKKQLzH2eci254idav6mkIW+pg0HJ
5y+o4ZJS/tSVx+4XlvnSc/3GbU7rFhIDMNyLx0kDqcuwbLYdA3a5X11f2hp7nzjM
Oz8kGgLaabNqNhq7WsykO8ZSKIJj06l83i6RktYe0X8eRxzKdl5zYz71AkW/cKlV
x9Gq/040uJewo+/gDF5NClbMJKfbUZOdwLZFOkvXDXEX6GiMmRgNdlTXfGGWV6Yl
r6eH0mslsgm3LhcERMJaw+W7g9ZpHrhp7UhpUdahfhIB+L1r2YAe2CaVBcJSCfw3
/W1RMmv+lD8dD1Ja36/CtAZplPukjP0uLbHZUOjk2xt8Pebaz6ikKTz2C9Y4RRn1
SlRpvDzSTLcbl8OTMj2F09fBKbupeti4Uu2IJUDcbEqHRoq3BpnPzBtIOE/+bmQ8
QaIRf61TCDKN5XKd11FcgRxLgeo8O+5+LgxUusjtIAP1UhSzD8RWtKZc+J9ahpR1
qQcV+CSvpVie8Vt0ykLFBVrjyvHQeVsiLf8G5W5we7/CPrQBJh37jTr1a9ovKdb8
ClG2vbpll4sgQXhIffCdLekgih1a5T6QyjCawjTb2pS5/7FQt32KhxVStSI2EZrn
mnSFuXzUheKcWyd9gespyZlly4GSxibz1/w2ibq47SHthhFvjok5IdC7EzOP1Wx1
k5fp2OyaJE/ffr5hLPgeNcxY4kUv0DQe7Ds3klQYxAikE9/ggO8QvRxIfBKujpsA
hwwDnVkupggaVt+D5BlXnwJcJm7fetcJQ3ZupG84VFTIeyEZM6qTkrHbSv6YN18S
X4jM5/JFbEBof5RzzrXjY6AkqwZXVERjzzVXGDEMhqnDNiL3HQM34Cs9O7NiJn4u
t2Hlo54tKHVrSKXFKTr5TbCXWZSnaKoK4PbJ3QB3AP25CWAyLYhaKN3UxaTTFs8n
wx+A6irUdzRRzWMT9WzsM010ygJ3bRw0sCtn84Vz+V0uBG8oGAR973Yz/yQtN7Uf
O4CH/g1+xZSta0TuoJ1jJ8GhtYjqzvL14eA/I2nNH9giQDSHLcqTsCd1NlXDCNNU
SdMwfwE8Bhi1mVkYmFGyOkKHgnRp420gKnxHEd73HmyNufHQAs9N20i6sFCOhmbJ
dvGuxYdwQYtQf5wmVsTMOa9grKnJRUX3U/lWZVnXZa6SNRCIh1zAfpSZsUY9AuEB
sD1cBi4+4AgK7chn7ySEc1akFvM4bx4LGyrlnw9tS/HvVTcnX6M+Xq28QU1kMavw
Mj2cru714FZTlhlAJzLA5oWXaCT6JfjybnO2T8/ank5dQ/ftgbL+v3j9be2mLPEw
HshQeJk9Wv3/ndhQfNWdiAE2iUFde/G//wh16wsEqRKiV/2FFhr9snw00H3UIc0+
tBfEP2/DoxaCmHW27tJvr2rG+m/Ule+/TMNEkeb6/1scCi2hoArW0oTAReHHH95E
qVxWUjBxGmg+2CCfpNM6vRegFsrMRU1VKqch4rnIEGzzTaiz59md1pc7uDjThUsF
+E3dVJ8ozKrUD9HLp8rxZBMOXl5vwElCcjaN9OomjnUS4EyVTlFCbrpOQtu0vEWu
BzExJtLAGu5exNHwt9kSDGke5IOEJ67OBPgNjz33hFXows4iK+HSZyWKGOqlq5oT
VSoAvkHyvFPrnMRjn26ggPu9A6Z/2lLvEXCPgNLNf2AOXQgI/PCjNKyjrmvmXiF5
jFoZlS8jL1seNCqnYSPq3zPuR1lCig/k1Oao20Ma+7FIvPF2dxtXicfgwg+ZhAcb
Ffn9f1bzP6PpTvr2epnb/EFz1VPcjCG+ND6xJAFd8GGIn31M9XlxxgrDZ1AkvK34
HIBwk7/yX7OmRGtwB9NR0VFose6XZmxSK1mqjZjKDM3vzyHyyltSVBV1hI5YsDKj
nCsc5HtnZGCF2hff+3Uwj5HvGFzlQryd3x5xIjgBGeeTdoioVjbEK7/kvdOHjkqf
53xLzFqDK7wIh38jC12FRwHb1WpLilZPeFdFRd+9swaSJW/wOXsuPe+WWdEkCqPC
zQS/hHlCH+6dFj0AcHoM6q9W23og4y+M/tu9RFKo31PHDxhCUXwYv1gUIuYRCZsA
DaAvXAWuXz1lGWurYQ32m/T2HgvBm1aimcd5uUVcJRqusxhH8EwAlCBymljvzIXE
ks0BSYe3G84pW1lS2jF7O++WraWAa+FpQE5Y6Veyd0FAZgOG2jO7ghm2z75YBo0t
TEmxaPFalwAhI+ZaGgtMIJyebicP9h+oyuIz4V/nEfDnNGUZP0KKa+0aQ9XuKmTJ
ye1KWkreTJ6vQXewCzm1c5CNLFQFwBMSszm7OdNZuC9WplAefe11t2x8CH1hXlnC
XZKSo4Z/F6qrytCTvJtQLUU+jHO1JzwF7vItd489inLvye8H+Um22QiiGOqM4a/d
UygF1Ac96XkMat3gZXSIuMvzZDRq+IMfSBVUiXIn8ILBk9FA6ZExz4J3hZ5aD/uH
Aw69WUXDiwE1eKI9inlvOPxO6JoEd80ILZtbR3WqKyZNlga48R5tWW6+mijUo6tk
oTaYoei8KBabANTolSmnCfJpNM9liIjcs1Q+rJPNPacez7f8LD/pZ5ULIpuYqzhz
OWs90zCql0r30ob8wKMihglfhTqt0qBvS0VYsw9BnYbbsolu0Rucu+GwkIU71wNR
IZjKuhRyiWLQs1oaDpKtpxe5cxuu0hGKBnHq0jBSfwqzA/6yxHAh2nQCiZxKD2Ht
rZisWDCNY2d7OHBL7NkXwYRg1fUYF/RpgqTEP9EW9T+IEh6CC8p1iPQ/cb1QU9LH
b73PUdzA6rJP7nEgYhTw7lAKx3NkQBJU8murMRDKgEgjCuK3ybOra33zQ87OXXmR
cyiLLTRdKqRThP/HnTaZAAgtxL0YgakFa2qI0qm4B77VQmyKFmF9DHXHgEynErgy
079R6b3AQ6EP/sJupI+Qw40XzGvqkYUPG8Gxuz7QUoSBDTtp/2xvHJYtHLJx6PtA
dflmoX/esM8bTzvfXV87wntAtHgSFm+7d+I1r8+teveZHedd7NsKfZR3jpPY5xNP
rrkrPuAn7Pt1nICKkTns+sbFy2xviuA9UNWl/m5DBlnJacdYxKtHQYX/jKdeuW//
A2/YULoyGxTxMckFIYdVH1y2PTv+cPYmcx3PmZ2QQtCVH2NTUMlu62vqJk+9HAfb
UWbxW5r5yot8UB+UXjanWTCYY8UtnOK4VfmWFv2sD6qTjs4LubbCizO0NBtNBVl0
1doDF9bY5cjS4iONbDQlHlBU6aPWCa+v8FFCDaTcMLO8GKyqu4vvKJR8WZebZ+D1
CuVXW/cnmUHFW0fByYkOIbv3RWosDXviZNUKApicOalYrN1IzTWoZACdWSEyfl4Q
ISMs1OF3X9U5iS+zOA2d9vT4DstS/yr4f+YcnZNsr4SMaKYGmooMIPK106d6hzdu
4z5N/5gZQfrkN8HAAsdZO2/4ZHHYyAYYg3YwttnVbtm8nQ880qfz755efNC5PVnA
bZiakHYJENasua/t9nCu0P5yHlcN7bA1fO/IHMgJjJQj50iTNzwzIKguUHZLiO2C
hNoBkQKJrksNkpUmLzNNaKefYO5xU/HkpUGh1lZY0LxoZZrRUA/Lcfu09/w+6+oN
HMq8+3KwA5Ckg4OHC+Jl80+7niZyDwOBN1tY3WhZLgf6qcnDz3y45lBrBfQQgMRj
QOemONRUKNtuLPjDLPxhIbGHa3Q0vRSPfepIKFW9/bOdMS37OHnrqYDCJCxk4mvu
2qlNC+Y+KJ5EkrbP3LAJTYlgAo4F5owQ0YvEO+Sc1ow3ePEoQcQs0YrMouSCUPeI
z39TyBzQRR6BBg/yDP6Iznmh/98eNyk4lozGmb96jY8ugSz+WjwDjk3nC9PrPY6W
5kaKzzCsWAKvqBD6GhdIw5foUjSEGN441KOsXciPqP0HVxQw4bDNp//g1LX/dVBJ
W6Xs9ZZpLfMjNtbECM5xjHLhcZTanqADw+L5BC2ZiHSgEjUJR70o73WGRyedUBqE
w5bA2YuFt/m6Yl7iLp28uGCsJtKq3YPX3o9XWDzOf4eUk04cDzT5wm3WsQwWwaK1
eB692+ov4Hno2dKwfdGUyXKFRjtZOhfQSEkFWoWWwCwtl96oMJMYYTHADrbw65Lb
eX5ocaGSmbwzMJYIPyIJALYhluxBtKZ8iPfmjiR3iWl3SDzO/uesO/ObU5/VC49J
o1cv34bkKoYiukCfxotbpI+cA1D37htZ8yV1TdFflc1tYx+sujWRpn0yw74d464G
9+w6xLYpw2n7lbAs2FkSB5nCnWGB7OWemrt7TvGf4Oqjx0KETrtPXi0ZQ9+2U6kq
lnORfubs1q5tG5VAEeQQajkSrewey0RkW9YIpo3sMyLmqhl6coTdZmJA0Eq9tiJf
XiAsC5A2riz3XP2Ty0cQWhpVSm2IZdXOlX8YKVHwdmNGosV8x2+7NTtw3/qGClJO
Ir7Y5e5nfPVFUZuiDFhLf5/m6XL7bcbDYD5mvnVKIlug7aiFwIX72as+gCzfInMK
y7NRd7trQhrBGMtkDvbRTfFROrA3vu8Ruo+Zlk65FjQ55QB/QH8V9Hhd7mNUIxe/
igschj5LPaYLDNOq43WU1zJICk9dcN0v9ZTxKjM4S+vryDmVf/cCS2uHqBtX3lhh
pHWDjzsDGDAOR32/DyzUs2jTZ9VPA/yIyaxYbqeAFKOPj0MgxPyVMQn600cw7hFR
ucRt/FEp2iNS29fqNXeyfjOQADBucXb38uMThGZO8PylptWqXr4HGIZB3l7KYDY6
DY3vw1Y+ZjhYVeGnDG1oPRO7MZhkXnBXMHi/RIClJSSTzdp9mT1hBl/jb65846YH
nnPG4THCYMspcuNR4HQvk0lHkbxhE1c32UtbxI8qEg2RyW0ejMsH+9qAWN7SXOXx
x4YAOmZfiYvwKwFtW0oZFiuSLy8zaG04hNnokK3wkBahJ42yv7STWyJiWfDVKyP8
+oFyvsyt6xsUP7cOBRgnnr0KyqlTtUObB87CzbNbXF2HhAdl6QHmu/JjYuvEg8oS
ocqpmtTV8K1o/0vvzVq98jI4DQrYF/Gro5S39TfJJrWdAMz3TrfjhgMRhnHVFCf3
WgQ+HMbRJn5qOD9m86i/3M13I6dNzGxjPuH0JVYWRnLG8iI+wzKk5JFCwkpL6Jn/
GpOIsx/flI0ahyNhStAPg9uZ8sFYWuYIFMe1a9PEnupe7MBzzhCWT0t4KJoRBnQu
7318UiXsALwTXuc7dOWAx5rDDfaViVdg68S6++MgVDYbDYB/v5kpfquHfsAtFCpD
8NlkhfyQ5/eXl/by76WQ18G9trNR8SCmDOyb6xApjgmF6jb2lqhA6l9d+b+c5rxr
LZkjdvadGjloZPWN5s6Vuy/IVt++1lEUMTtlabzzm8lVRbIbfsqxhyxdh/mVhfIU
IKRGulTkXIUvKvdUow5J++LdrRzVBeiuyIf70lasuHy7N2qcfzNWuFNad5n48AKH
zZG0GHlowuDFxViLPZC8Sh+0JdfY/K0Y57jqZtMuUkRdFnPPcSsz1yQGGw4mdACO
+G4TjJZH/JJQSSELylUwR1C/pU+9HwnhAjWlg3I5XC7LL1Ipa9k/mPIhAV+C65eW
iBzq5sv7h3F+bv7bJZZ6LyDbKwet3NPEPaIMz95apAXVkRkres9bn/SWWKpLmNmi
H2OE222W/aYUBV6WSU+z9ZOdFydfQ5tzK+Xs4ovNfHwxvfHpe62l3cqiw3r+I3Iu
75FTvCmIUh3ZBP+1f4TFQ8VfJTWUgT9SVcg9apezJ1c8cF44BPKlBQk1P1CjbzGH
P58VqpymoSUGQRkRPQ0Sm5aO3P7F3ZXP7A74vb9CT1W7qN9twBLJPf5FCpgY8bgv
iHmxqN0LiOgBE0sYwQm+mv5gQpNE8BoKuCEQ37yPlXJOHfXvUGsaqxG87lutkiQ5
y/+fP+bWvcGr6c7mVB+gvW5iUDYjh4oERdDvfBc1KJuIaiW22M2qdccwJUyuwsvy
dTs4QZBRB6xrUBXqwMkzVYAiXji3cM+xOhD2VFCzQg1Cfl2gAk8PfbS0rN0j6QB3
/lyoQC7K/AZHGVAaLP6qTgD7iMpvSD7mcYZHxCCQfD7+0g6opM9KcBksbBB1JJy5
DXs1GWUcbrZv2bp8/XeRz9K3uVPYotwaNWcL4cygzSaFEI/oOKpaAMBtR31WDFx+
T110dd9u90B4yw8e8eOJlAvhqR42q07F775OoH4KjeZ8867FXgXn5CeJOfbFWq+H
6I6t/xON2g2udEwM4lnupV0L0Ngf1ScUrjWnWSGJFHD8b77CaHQmtfh7MHp9CXVl
rG2fFEk+OHOjXOy885q5drZ5vuXM5GKE16BebP2vUZbB3xpVQXhsQ3B5Z1lQWJ+0
gPXBY/vmGKrjktZPU4dJOKbRrGoBUSZc9B+50/BZXdoxkjndWc8Jg3zLLTq9vHeU
IOwEVqA3czokR4O2Ik2TyGxdjM2z90cEGdh/HyuFZvQ9y3F1yvlZ0RWa1Wp//thh
y7MwXSAPnA2CjckvcSFDohgUZ0xGIeDMHha5p9DBWllVjVaUkjcP3xtsHkWAAj1o
ZctkKvRalJVjaEH2MVHKp2KOW0uRFR8UNBJ2J9r8U32mHeTkstBaxVsDpBf3omSv
jPlDwfKUczBhvkH4ODIpCrU6XEmbEhvBhBrOsSX8Fsynxz7dJ2AxW7QHUG/bLHrk
LxvlZt+bdGhT61ZrEzuX89hPkNcUeLYEryBFyIlcjTJy/Id5V368zsbdEQjs5o1v
SILY9l7GL+p1v1s2mtrBrTsGHevfpJRdW8s987AIsMOcLjUG3C5bOpZxe2vzVAPL
1mcGl5KuKUwR7136CymRX+wL0aUckIXSsac70C8mEk4X14T5/gscaKCAzVNQHkXE
cNHLBHatToKLQAvoaoiXCaXvXuNGFM/eN+bBxKtrqkc27BM97WYCb/OP68l9ZcV7
wvh8pjebxlCo0tWwCFhpnVD/lbtQvQXqf+xo7TydDz/m5v6elTbtFC08Nt7vCXN8
AbSYlcnJeIIyeMN0G8iUxagHZDHq/fXSra4zlUbPzYOM+kaz1qYDYgBLBprL51Gh
PThgB9NMftn/KwpHx4BXacZnXZpTxt5NQJN56TAiUp/1xOcGHg/BZ7OyJRtlIzY+
45f3VyyqrA2QUTcspyr5Edemw5egroSz0PtmsRsKZY3ACAZ/Hb75wsmxv9GPKKt9
RAmhEOWUbA5TdpSkb3h1oQNODg6dkAjRdQ5+v1TqVyytPVi/Rchp/HapEA/BtiVI
aj8y8Drt/yNkqLDZRne9oNcyPDTzX52c4BQ74y5R9DPBF94YOCJGxzKXsQiI7Pr2
mmZGdrNaveUvcvm9Aa1QIx26beFhO4VBxWQAKH2wLldyCcfINFskQ6WFb8bXrpOY
T8keSsk84ReZLHSSF332leFbcIDOIzUs0yJzFGDatxCl1p8j5KRlZ0vKMPMQCtML
zY0p6/qIKTFO9kKKgJy9ts3kmXyPpxPUL3YkYHSUaicXjfHeXkKNAURCWC57iayR
HMzw+3rOt0TRtUIVHjB65MnOy06HGNC+RA33R54vRu1+65P/PdPM4gKLnE1HWzCi
NqwLOUeHrBhdYIwGRQsd17DD7PtW3LsZvt+IGZcA0xVaM69FwKrB6KdkzhfbZbbq
daaoz2w7bnJ8hZdfEiPaFDko8W8xKQVmtBMlENPdEZvaIAiYERpbUpud2VUmdItb
NQZjvo2KbB05Yr+8/njv25aDvcSUASVVLhqZcvH4kPwowRyC8ov1K9bJZuUlsySy
s66ti91AhRk8dpsMZXlsndhknkEOrrd1ChW7lZ5t8IbtYofrLMqJ5Ri7KsrnfiYu
xJab6mc5AScoPtbHs2aU/mGXMLHkOOPblNeO1utA0063myDCJSQw+peTTHI9H3xV
8JMEZjnRzw8/Nt5wOreJcaJP2m1as68i1zFqOrjc5hnbpv5M5ud/QzFuxGmWGkDn
OmUQe3DhbiJ/cgppTMt3RLZjs0OMcUm1to9JdwN2/q3G5EH3IAQEQlNZJ55tAGoN
oeU2pK/bp0ISQMWleSVRt69Lwn0TZmSozoEpo3pxuO+zgsvopxa4vwXeVEol8Mxq
DVo2MdMXSfMKBfK0O9Dt8jLUHnbgMTFkBXNlXcaCQ0KBiaV7uK+CT+D38dXjaeUi
1v7TeXYOSHWyKrfwlZacR9bqr1re6bnXKNzk/tcEkhtfMa8AA6BEjhSsz4F1hmus
lVwlX92Fw4f7wwBZA7OSsurOMMeAmAHPigvQK1La1V2cl0x4lsCYmlf2LKAuOV5J
Bkir0sTkWpA+4aQi8kjG4J16l0DHYUo7mU1ChV6BS/hTn8CEocdMW8LC5YKWJbQv
a38+xzIe0nTRGiSgA732DryBCorsbG7a1RZWjEoruNLcc3jOuH4tYKTXELr84cJE
AGiB4jJ/3353o9TkBaAola8MD6GI8nhcHfvKfcAxV3f47ziVp1mdlPikqyU7Whqn
ypgf7rFMcaMfuYf9KZ/Ih3YGkr0lMXxw4B12vTeCjnyxd3XkG1rqY2Q1Y4s4h4DF
fQI+8sRkqjDeKm5YVVUaV5WDSv2prmKPXK+ZAPdYJyQGkwyKTjxT8wvkuf2Db4Kn
sM0SNDEOfOE/1Fvj+ghi/XhkSxS72uvEkRSO1PshQfrPBA6wMLSyxHwdJECqYJ7l
AYFPRTiaL/m/2uqRs0bChn4vQYrhxWH78vDjifcOzisGnUQONWFGEecuO6zeMG9r
KTWD5sgDO7F3lk43/gaDQltYIVXgSDVKhCss50M0dq/eJxxJke5EAKK+Rr09YRxp
bTro42nnFKLpv2+/triUzsKcpoqsyP+BLdLQcUPUI+FEU0ic4DzhW5VwQ541y2P/
KVhcKs7VGI317Z0uPhwDjBMB5v3V0otnpUd+6Hwqn5kZjw+ULHqb4CN6HgMUyi1F
zxI3EctKt8VuFc/SeSjChqMA/mWaX34meXftg4qof2OL+mgoNwmURdo7nJyh5fmh
KeB1N85cCsX/xnVdE90oIQvkwaj5wEeIl5BDflfVM35NDu004xIfjK1LjrBvmK5T
22Ne7tNlwwh/q0ZKf+2TIGRtRRvbLJKj6xp5F0hnVgc1P+B4S7qxVBiD9tjnxo0X
Zaoy8Sl69RVeRO072K2xKRBM0ghnHReDzBc/r8ifEbG0LtYXS3NGVFnA2VMQLFVO
b0GJIfWvQzdYAPbJaLvNFEWXcGAWb9CZTiTNbHg72HAfpQSMJ39cPKocZQgJFvt9
0h+RomepT5yU41JPkLhP+0RJRIRUCgLsIpYbI37d1lgBhZDxmBWoNblQUKz/j02S
rkdQbqLf83MbACO3/yGVqJsMNu+yCOyu15rAEApS5hnPjb3lGZPiYOqLEnGVx17/
/zcLU21fPBpzz4U590GT4Gx6LXjOTt9VnLI+fI4eVp6sRih5UJmIHt48Y+seIhQD
h7gauF1ogi5kkejM1LuENFEhTzClqiwILxpDTZ56m2wFbuJeHrMag479lP47Wva9
FsZrF0v3W31VCHkkM5Ios9UvA9HBA4lPZo50MjSeQM+89E3Oyy/pRU6szxedVw0k
uKOAi1X4g/FVJ1f+kUvtK5TI37Vv1Y+qV45XldzDn39cVhHU8uTz1mfNKAoVQMqL
o8CxCOq3K6uwtDt9H2l1HPo32jAEl59ZuyVGUsx5LVnano+P/rTmVGpAe8lTgA0e
yuU0G7xCFFvJY72sqB2+Xuugj85UOTpufOTr+YqdItXwkYiy93/BZa9u4uNVilnO
4zW3KuxPRXLHqtlWYBB7NNVJAeP9YgVeL3gYHrX90dKBSKsGdO9bFZNmw7eKrsuN
LX7Mig3e7mIdplLU3FGA7/NH8gwXz+os7NASwTB0WA+ottTNVGg5y1ef7FdZMxEB
KTficD3uKaW8mI4D7J7j8ObkAhAgE2FFj3QxBK54beKYuUzB/LPrKd+snvqCdsiK
e41H2II/TDoLqSG5C05gM5ZbelxoO70X2NJhRDZEtEuJ0ARiPC0PMq7jPqe42udU
CYo49eUeE5+GW3xHoGhqTAZzskmMlZMluguy7l16pzH21CYO95aRqZ4bZPYvJERt
1qQ1hu0kV7ajGvTjaA9I4ZCgHIqUD8IUPz2DrxzaXpHa3FtVrsyCHR1h23rfY6JG
x+AtX1hW7KYJE8tgdccDm3AsboYnUB9Os09vcVCp40LxCxsP6Wp+pXu1AgJe1vFj
WsgPztAilrJdoM9sjKccv6skp1pqsGoWc/BP2xxRJ2L0tl3M5DvBvzyUbfjTfK+B
uad42HLNuhE5BKrRNGTExfwNP/Q1gSgQ5w4Ss7SCgvCeRp2RCEc0exF6fBJlUI9g
MO08w0wx2F2z/3GydLnpcAvN9U8yFs+fnGbAWrTLl4KX6g/Q1pLPKAZ0saQYwkxu
5A246925Du/2JLGA9JoePg391hOL9djPWpBp12N31/iI1PauFMK5HXYSyRjLpN8s
jyX5CYV0l9Di5rTOLlpAQxdEDfe736gfsLizFwTgLyab9uM793DFF4MNxXqiXL57
SWV1hB6sLvb93sjXXGoaNHB050Tid20fZ52i/ghJ3YI19qurJ/XblhpWxY5V2M8o
o/O71we+4DBhr3pdKUZz0ThWEM9+o03Y2ENtN1qwwVBqnxiFaRPT7Ahdbb57yRfz
0RzWy2M0ML4bIEEo5gJqNkYbvM89cCQIXrMfr9uLXgpF5nbBJYcWCLpFyZurXXTn
frj04RN0ywVhTF4fspzM+fsgjBmDVGYtkY/T26bIgXxodO3LGzrptHE6rfkLNKb7
fNbIHgth6+UBZOPJwGZxpjHJO57wUvNwGpgNQVSp8tDRxRDQxGIsrUrwKBFG/uWd
KP9oBpqXZIDwzFePKhXYqIq2nBUMvMUqTOSvuMEVRl1L+Thc6dg/z/M2lVx5OjvO
Ey65z11v/MgMo2G01qP5x8lh9EV8diJrg+Ieu8O4SMYS6FyRIFCFfUSXZ90RgO8T
IEP6JH8jYQucIrH1AZ//ghOnrY5JctAmUiAGIP6rMixQ6bTaSn09cWkNF3G1704w
F5u08J491jvsGFxwThjbg+IR3umX40qDV1kBPSsBrV+Qpwbh6uWBVC43TWZY6tDw
x+M/gALf0yl7dnBEvRumg9mAN7YZ1PnicAajqZtlOX92ZnASI9uaqXYfb+vVgqfO
CbDEJQQ/qxKywAFCCv4Pmy13cnBZ8UpNL688XFXtjpEP/6HfhaQYQmNZwfptLQrw
xLNvlj4Ym30/+Pk8QY6uB1NQsG/OBGgbxjqA9GqPLGEktoTwepEYc47KMd3JO9iv
p79sF3PmFrGj8LMELiaisHTVl0XPhH4O1xI+ush1OjlVmexjxG4TfgfPcqM8ULC+
UUhRY+W2QbZHUsi+/9O0kw7Eib9iVq33yc8VF5+xGkoUUUZ5MtoCILA10FlvLyyo
HjKWW50wIpVxXMAwSFTONkl03+mjHFgof6T8wNg8xi1wSMX0iRwNzE81NDzS3dFo
hPK+7RljqABrp2/4fIG80Xz4cnauk+N3v53JF0tYSi3gEtEpJCBv/9FfjOeN5aZh
u7C3hS7JOh5C73T9CStJ4tfbzhRP4hlRkQh5oo19WGABSf7ABKoXUoCHJko+eqjn
NFUMTQDvEKocAJ9OvHDnRKYXpGs2WljtkzOMlySWT4LFBcLnDaoV4rGsYIUi4fuk
hDm7CM9Q59kK28aZ7VmxihgFT6dKfh0+VM6qHc7d8rKzCnTS6OB2vHV6ss/T/2iZ
9QongOkz9d4i39IHQ39EPnRWOZwheoTRC+U6B44Hfq227xKT2hPOrwx51/ehR9X8
D1sD2GojDOBrLDw/mxtapEWh8pgU0HYyXpnIfAVgg6KrM+S0mtGEiJN8s15X/0X5
LWgFGnm7Zhk8sVnoyYJPkUWXjYfXPYW+OiI3G53jtX2+4W1BZptCs9eUEHuApJ2K
uqDcZV+035anwM370eMl9U/5by7pYJeQ1Rjn5EI29FkxlbRzSoa7KIvuH7f8TBPj
NbuO2zsUquEZYUjUHY/BmWZwVbslAbShjlWWNpQjkEo8sp87wHE22Zn7yhMw0nCS
dOpekEvVo9SqOF6nhD1Idj226xPQd15Ykn4f9kQt8QhMKE9JmQlG5o5O+DvYpRdY
bDjTAXOyLOtUy8y/ymIUW0G/65i79CzpIv6NZsWhqN4TRUVkQRJwhvvuqifU1tm/
oQ97s1E+AsEquunEYmacYYYUx3QhCDgaq6UwJs+1tJ0XQhuWstIedjuSrzg5q2Jg
0vx+glgkEiqsM1c0dlYbIGJsVWRD/S9bo1hjx0RFr5qSqQOjSdadwTj6AIxCPxdp
YL+sDQuv/DSLAMyypnZVusUw2fFhSZbMZnBPF0pwBbGrrpGrwUGwJJoOr9wSSoAb
jyYNzQm25cu5IQ94QUDh7YVmYIFozZUshU3WzCRJQsqsWBA38IIIhKZDcRZQZ5sg
kaT8CtdTJUZlEk16Qdbh4WB+LNSehAfwJI7PjVdIR74UlNNC1JvHN2cyCCp2loBp
AeNyQu+yrt1H70uWD4kPA4c8svVSWWMXaEq3ukfswmml1O6wERejj4N/xqPTm46e
iA+ILfSdtEwy31VIeQHv7zoyX4u22xKaB2kNwRsIfp9kZNweS0TFQKvK/6HPKJS9
R5FiCe+C1kQFAAStdU21retjE04Ur1BZioayNa5AksEeIgf7SHU+inEO1Argc8zt
Ten9lzgzsVdPjK+NgrLJ/0NtvkMdNcJvLWVHtcjPfJ0eVqVuGifv4mRb+/apmxGI
pMQw5p0RztedGu0xlgIR9dEhwTCq6pW8w0jwTzK4J8wizAySzi1ei11GovIb2AyA
lTeEskr/HB+t106qA4GxW9+eG3gvmVDJMoRg/c8Ewv32nQQIDnm4miUN+mL+YsSq
vhGdOrdT6DcNp4ivwsFCiPb7VlXDMzIYJR1dkd1fTeBSWqcQFqMWCgCbdNKPv3WG
PQFZibr2tq/9I2XYMuYVJzpDh6ROo+HAroe3nIObC5PtKdF+Y14qeUvTs5QrDNgu
V6JBBxA6f4YPGsDe34D1ggngUC3yqZ+IWsK2lStZhIEgafsSW6st73IAXviQmY+8
fTXP43ppmHjelQJGJvwLvO+3hg1hfh0gLehOsv2lmUH4+crep+E6B/ClF8HZoTsm
ing7Ddn9kNSVY4bNHgDIYWx4S+pfYury8HEy7DBz7XmJ586SQ5zmRLU2MMBLrNuS
M2wEZkdVhIUjMGdgEFrAzpI4EA7yBO8OS0DZrumD2aWNf4qS3JT4eA/p0omkvnmy
sAKKZPDXAy8rw2XMToDJtxEV5dXbeX9VfFMtYWuZX3qMBxO4zjzYYaXLT1YJIxcM
oWPOS8brB5WD02lY/HkFUuAw8ukMsQe+KLR557AiPQ6F8SaH0PKT30pjPkz8LxqZ
f0n2RhLlk2eYGUTCa/+ugZ45TuxqVLmt5e/5/wgUUQVI0wOEpON6GQjvfFCDPz88
PkHb9Lgnl2Q07Bt0ectN4ezskNbV3279xlFfDmgixm/uaq8drqkRGDmG6V/dqMSO
wCcoWy2RcFui/glxuYOd5joQQyUcJqZc6qyacbsi68VdF8ohRtldrG2q37V1SAjx
IqmuMolxpmIQE/4cohQ/R7Su4iJshgdMGaRhG823xCQfSeFfEaqyFVkOkkvx9dA5
asm5eBQzvJBeGvNQ4zs/LNxSqR/Byftb5OmRvS+ih4rXjrtKLEF/K2vKOvgyxeOy
x3AOnhaPOyMqCWsePjMEl2Xx8wfsEngUDq8d+q5z4dg4bUxq4k2hbwGa8oyVyjh0
9ueCk1voYhUNlmo2dhNR4xLEzngZTthSVKfmos9vejpnQCdp/rCn9UOJpu5je6TN
ZbRecBMaXCG/sygnBYpmZ/c0geqK8kLAm/7ZdNnSG/LhKJ2SPqgTIKcIo3QLciuK
1zqtDCSz0/ziBRquT9QXhkQS3PM/gQCgaieJrYptyG8IwLmhxjynU0cl9QFDEEVk
2K6eNfrP7IBNNgdRmr83A1rXpz33S0EharHWkfkRxutSw7NwOwd7SrtjGHKhEAwu
B3Mzq+R/4YqRMkbe2P5w5yivwGtDjAESsX9kWGytqhtHS0TxJtzIaVDp1FCDtMLh
ladp8YrG/f9rBNlMpyjD11Z2gdQp1noegzK7F/P+F606W36jB+weSfUrfThc7EP7
yv1X7cSzLOtR8A4XFptquBuOlPl9gaTKeIuU1tdPwcNoWo0WvoE+P4biWqS29R40
CcHLwrWL0anIfx0WpU5MsfyBoaqy82b2x50DpNXvxYwf9pC9WywsPSNR/M6xydXQ
nAWXonGEVRs71UCdkyjrxYDDIh/EbU1x5Wj8Cic6uugF8Wr143KCgOsuew0Sh3DZ
Hm1XmeJmRxUQXrWj0s5fsZfvh7w+/l8VoJnryTgns8nFV9erkFaZqc9shq5rl27D
Szj8vLBgzldeh6NAeYGuEPGEWdKjnE1uDErm8YhpE8FWwcpk2WOK0ZH9c9PfTpUY
gZt+qBTJTU9wL8T5pH+mouaTwQEsvcs58vb7kqvyk+I3xM/J5l1ygGJ3x1tXcMJ4
R8aTsSGroxsfRAqqOQb2PWocGmAzFGdpJ+q10kh6ZryRSR7sh+cnscSk9DUFFb3B
rzrLh4KHqJDmFRJbzooleo/xIWWjVFiPdJF0N077bu3bFIYlsDmeGzArdZhvTF8R
4SWYho8GC+aYEQd9Zva782JQUVx97G4PWj5ZYelo8iJU4F7kPRf3R4rCZqa8UNi9
C1ngKfMj7TETXp1wWn1DeTsXxVhY4I3Wj9IUi6Jr8F1Dpxu/89496VRefnMFtntV
t6gWHNZv5r2aw5FgAZB8FrxdhmrAriTNg4tBSgG5eHMQxgJE33Mf+EyAU2Bq61dz
+KYjVx0AbYKEw8LDBHrVRtkbHsJFCDSaUlbUJB3XzfDFIX6Vc93iG6cgo3AZLELd
7h+6eZsyMHeFBc8tlICwhAbggQ1Qe6maLMd0h7C99r8rjprduaIHorUjI9DKulW9
vKDw/Xp1HGC5knU7/zNcBDSJa1hfnVO/C7SCkNHxA5V2VqRDjlbdAgZMs11hboJu
MhCWiVmDrckZfhXAIKQVPil7yhQ7ihw1T6tVhmMf+zBiYq+oqq+bVgkNNxA9qnjR
CEpUeKhPXVGVLdrkW2ZZIlBRgMwpgYld0pJ3CxoD/K9CVoWrfN3k7DYUlW+qeepn
Tuu4C8OJ2syfrZy/qmha2TNHfVEgYLtDqct4br+Xj3CcWkabxAz6vz99hIn6pCfM
qPw44jIAbagGe5oNIbHA1Bf+E+KyvQxVEvEhrFQto3DFK5rSjx8TKU2mRlZ2eOl2
+Y63Tc1jwWyB2hpC9Dqsj212Sx3pV2rIZo2A1fep3FoOEQ/V6Okwm35Ehoiq/Rxj
HIvbDy4Vin1YkVMnRQ0WMTNUXi2EnY4K8Q2LmkFzGUKEENCdK9BJDg9KvhyQmw2V
o96FaxsIjNvsu0YQE2q4Tc/7JOMMEMuvl6eyvDQlcZzcWod2wwkeExfhG50l86TE
x0yY/5j9JMhCO6ScUDez8PZn5xz5Jbx9FHaW25xDNNHsv/rSk0Zfsfyl8tnhzlWr
OkyRn69xuTOdntJMU/Mol7SXMgN/K9fFsdWrj2ko4KB5wEggc9+4g9e73idn4Swe
CJWoi9Lwa/ZZAE4nVunQuS7Fy9cJJ9lRrJhMTDDBIhkdAJbeJO0fHOSyiAz/LsI6
s3K05f1U+Z+qfJEX44i/wqSS4BIYzRy5E3QOfARoSTCB1IMFd3CM6J3arwAHlKY/
RM69mw3M8t70xO3Ec7WZBd6xiWGtSjZhe3Ex2Z9qbSPEtjbaJ1vqfBfVwkukANVt
JErgG68W3iDCh1MqcZw0W34kiq9WmELIyuMXFsX8OvA1TPxqgt9obDFPn4Szuwly
Wo9VenhGMgIimhgfnI3UfkliQt/HTrY+UDvb/HPZ1Rb/g6G92doef+3ldi7qaTiy
fduGZPxX3C7JDYaM/O3xV3i8EKCNpBWg1fRAh1VXOA8sSR2E4qgKZQbloqkPxYLl
qonCZCfThdXLGLF9QiZu8xLSKhCaoRiedqeoqjK/LkdYzsfPrEsDlMEeFkp+X+H+
ubpsZ7hTjv+8SCeS0i9ePoH+MORfazYBenpuCPMfiFCW5dyHV+Y284xWLr3sVpZd
Zk0VyE2jZxLCkg22l2pu0X4sh2CW8WI7V2p9kukJVoDYgd2TbR2DEwCMC1jZBjDh
VVE8LmBQV/+lbpjPe/Fu9qmJGPKKMfKF/NrWca5Y91Wh4NUWDL+Ns+0pp0+EWE1J
bQWHc6V35Cm2zp9vST9Hbh3zqUv3KqV3X0tmn3uGdJwhbRIdOUOekmWcjxPO7Mi/
az7uQBR3dE8q8veATHiOaacCvUjEzfKGeRo559f8S97rKLv9/Bq2m3KMqtq4Op4/
oeXEi/HOaIhozavML7Dkg535nxWTeUSAeTQ5fTLY5zY7H1scYwSgqt9vWQQR1cRK
FbWO5VCh+KU2MDv5ljN3s/rdsXLhT+FOewWEQDNr797sNs0qysJT9dTXGy7ppsu/
fOEEqO5De6W/y8WCZ7FipUqRUMQr0xS4ZQzDh7z2Ig+V3F4TfSTimya/J3+pNWzE
xRYCeA4zemFib4NPXU6wX1+WvL1CIzpwPS9tck2awGMc3MocLoj9ZEzENOsI8BVC
+kdZ2zt0Mn1Z71bKnID8ICIYJOA690qCqB3axKYu4PKF0FAUPXa3OHtuxzAqN3PH
9PEFL4KsFlsbn56BvkJ5VW0KprFjUk2+BcDrqohWqpwRZfhoX1KBlEgJ/oz2rSXp
ebOi4HHrj2qvYNVqw/oXvxiWZP9r6gIi047F8VNiMFDyjnKvv+Fsvmya+dLBOrfO
zB5eieCY57Wd+NszDqm6N9YpFF6aIhzw+uED3xW/l9VmYzZQw8hgxri0namoAEUJ
gc1WppUcWzeleTjWn3Pw5oZ8CK8PTfA0EIJlupxK4Uy6bCuXpuPNIxScBDpzAymK
TzUOxjGLZ1NnexMYbqKMeTisDrKhOjFbJXWY1AT3zFi0YGa6FLVsYK6Fkm9wHldO
R9you2rv0VFs7lTlu7Vdzkb01V6/1srjjwVlO1KEWWfTuRR1fss7LMwOrj0buRj/
fiM1wDBB6mFLM8PkWYvsAuhI3W99zY7U/UHnoK7/0BQoPY/F+kCgxe4mQ4M33VBx
zidS1MpmwWDHANdvnu9tj9GkmAyUwyHv9G3TEcmLmn4lnxfGW1BMroSXy1drD9j+
Mnfiuvzq6eu2B2JhK/MdUfMPZ0Q+0UANxGh0VKMM8o/XdK+XotovUVIZFHvRBl6h
BM7qKUuYYjhCzJD4fDs3npefixzxuW/cUbSBZRlPYrBRUpW59iXekyvwv6Tecg8q
8cuZXpmqJwDPdZVTM0N5q+/1/ej9m12VolVgjzgyA5p/sGvpm16GJmZfkBMnNNu+
J/riXTJbFBilMYroVq/luJTiGnKXYv48F96DlRNN+CtWVwJ8XjPErOFljMPWuD8E
nPUdlLHY6281byX8tvmkwghvn33rV13YYUAvEj8RM6e5JZR+n3dsmyUp5rHrp8Md
ZrRcnp42dXXegfI96HiAxhVqRzTGetSaNTN+vQNvy4cMKLuVxbNo2D/2hRsWBG4u
rARc+Q7LW9gHhjKOukTsQlmX6D9hMjriplQrM5y7O5q5bKVu1vH3Mq+1GjAODtNu
JIzNDUV/qw3vyL9AHSs6xVOWNRDSPaJeLvO2vshbhFR4jTlRpeW012CcEyxWsjz/
FlJAad61Qtc0nyzXndNIIubY2ghId2CLnH0qL6pigFjKbFBtU4BSK4KZqc/e5Jh+
WiU0rRwrZWRAVxFGkFBdAD73+k1Po/QEE+GGMYqDUL2PKsore+gcvwYCjxaCZ+41
hJYHHGOerR9TKzxIM2bGB2TafX8ziyBDY4XqU2RtZngZFfbc9z6OqSPNHurNlBT0
hF2zwFheMa2n/w8QRrxIQyIawqDw5IyS46qE33eEdNevCC9qEFr1PS5ndm8dcXmu
+JdXl2i0uyi5q/5fVOh40EokzgqYstMtsTtRDkI7/meSNjjuj33Rq2u84NbQnaLN
rrdvSMeGRo4VtLAXzJtdYTMoydgWwQLiaLsUXc1+ooaPPdoya/W05Ci0NfQmZDBR
lteRLXQtL19OLGoeHIcp6PPyg6/Sq1uU5xV+PBN6S4CkPguMmhW8+YNCiNT1IS2R
t9bEAXCbpJVlmzdA7MUqV/EwJSmSCOcbBzYrH2+ClyXZOmMUo1XcKsXj6buLGawx
D4ucvTWUQ0z8Lrz+5UEL6Q==
>>>>>>> main
`protect end_protected