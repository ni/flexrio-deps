`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
hVdJHWSfELCmA4ds+csnOQAALbB3ps7EiTSHEDd//nts1r+JQrRE4d3bDPRJpiX2
Sl8d+xAK9BIi4i+3ruAzYvB6kuD7r+gs02Jsvd/1kn7JYK4xBxCjtdDFjVHOTEl1
sSh1oNiYUwLuwR1yKfP+xBhqxD2Dv6pCKhH1NdGilpJQ6cvivGkSunAu0tzP76T0
4x1pB179E7uIeRplfHWX03KzEBF+eVtfgXVp2W1BGjfAe43y1pCvNYZOh1+TY62g
EgAFgbo7pAujZxZy/YSiZjUr2mGp7o83qMXyusx8+rQ41D3X6rxfuP0RiId2pOpC
6oq5Dfkx04a1dk4s8w8cVg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="Sm9DkM+kBxuxXCFA+l3fFkxuSWV4xqRc4Nn7Ji3ukao="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
m2emGBqRy4AuduN4dffN8194qYvc9UXRqiQc56IrQYMiIVQPyh59I8SYabcDdspI
7AFHnvKD5YaF6tQfxWm+mlcmMEk2Y//aUjxeiGGs+RkKgbHitJF/K7nqg1dmKvDg
a/GaBCq4Bqh0EehlN4ntP5HxM4qcvSfh5m/Coe3drc4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uG91daMWA1mGkhgP3oZKMYye3UAomMWgG80HuuXg2E0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
c9NqBF2D1wSep1rW7utzHsk2j40aow1MnrccxUTvKej2Q1cyeDDbgAml4eTSXI8z
QYgCADtWi7S8BeChdv4B2VxKcS7CMq/DaQrOy1MKTfQzfAlK0iubmlTkljLy0Rwd
Niazd3hQVzwxL2j/Np2ydl49yF5b18gLl/3jD/2YZQQpd1/2K+Jxc23TORZ0xSFc
gqAHKxdcQeen7xSEfqvi/3XL4bUj9ChMGPbk90Tm1z2y2HzYv3rTYcRm/3bsQKcs
As2mEKpU0qDTH1SFbcSvt+SVLeeNr2WNWq5bXaP2K7FiUvgIOBS4w+/I7gKdAGMi
wkogqZjuhm8Kml2ruHeSlmgSFn7dfIyHns/ElilR+oSZi6tUUGMnAQRMdnXul2XH
RKHJ6J/SPUsaugfnrwiometJI+fBsijr2B/O8ittSTBZWkhfgLbxh6MM6jj0YzMN
/4JQuKB51lInDS6x04XDjI+lHKKcUo6/fVIBQtgU/S16KaX2kUNJ7tvmRFE9HEA4
iBFiUmed7VAIu/jO0QBqnAXPzbP2Vz+djc4E064qzc2GfW1wkdEn0CB87xSf4MAY
eW2uKJLrMN1uPCz86CPhXN2qzVwNSEkHu7jDqA+fa16YoNvaT+3AObwSkUilcNx7
ePWdvD8piRlH3JTK7mVDhxApL6iI/VNzm5OVUyQJ1xtrf12tMY0qnRjzggC34Wck
AlZkFtnIa08h0F2q0S/7MFWmVE2wQUjCb/bSVOWm4IGwyz7qQWRuLWFoNszatQ1o
ADvuItmSx2Qd4fuVkvwuGx1IMBy0zHxbCPXoTcbFv75AHRfgu357hD0zR2AkKuNm
FMN7LBJt2H9iHM74sB58A/QL8S7/aVgY8brvuFAtXQeUFTTnKFYpEfPGFl5hKFmL
T1LHlsuTWojtYQJsZYV7GjX2yI5BGgNqg972uo8e509KZA0voDiIAE5+pFUjKH/E
yy4J8Kj1hcBdC2CleEVSUSysGIqVOS38x3Lk2DRHJhuNECCEcrcSBA462MPYh7Qj
vkW1xcIckGSgdyQmLrIlCaeG/1J/cfzbLdjm/mPV7MmdGaljveRNWwkrzJT6/X0u
2uVOR94Sgf/ABw+IKT7Xa5brEjpSvb9NmU+pldTz7tc6UoAa6E/7T06WHuK54At4
RklSb71WK7Zd8X8cVLFtBm2S8OM5fzx9DnJD4hmjYQnNDga2WcnGScG+I3sM+W5J
KxZXHec91WS35/ucIOKwy+ZZZaIQw6Hk7f2o6bFDPJMz+ePqaE/SqGuAZ6PPnzN0
4uqhsfUt9Ina1PH1BuyIDOE/Cj1kahUIJaKLyhyAip88wpRr9qJVpdNX5Z5vYxAk
6w7m52n1Gkfao89wAA7XcUIfoUxU/YyeG7UuIprLUWoGcbRq5c8wX3NMn5OWAS0n
8DKF6H27Y28i8ff2XBaOdQEkhrckOiY1CUz/n2Thb+bAbnfbMS1FqPTWdXRsvO4e
FJXUibxt+ThCJwhRtyJk6k6aThIAHAxsz84rMmBat4jUxpAp/lIGG+x2TBG44pG2
QEYBkraASqBon4zFAYE5lvNMzLNZhsUxyCfFsSiT4Qq3rL58EZCpijYGW89VHxc4
gdY4A+wGJDw13JZm79hwve2g+PT0rXG5UZIEX/QZCPjO5ZrtBk+Ivm2SpaQUBsm/
6QBGsg3MuA8yTHQXjQurjTZDC5E4c+gd8qihIFTmc3SF16yOAiLTqVbJSDZyufws
t3xnud+LB310M9vcAj2YL5GgpYrp2bQ6TaBQlD9v9e9wjDEpU4oOcWwSlPPvQ/b8
Y1boO7xSvMGQ4VcTjMkay0jDBCmmPHCzuxe58f4AL637goO6aXrgWI8q56ADQa3/
vKlF6ojNRzXrN7x7KH5qgi9H5Ags8mg6jUPx47gTKPFMiHAMBTEdB775XzQnJyhm
QERsSfQgMbYxpde8metOaFDgFJsmEE7ybIosr0GUMmpOGb3GX8j9p4bGRHjB1wcQ
IcuSWDD4DRO/F+BR/x5cBe37AaDauD1fEEe3B3LEwWBnT96SnlorsBHBx2Eku+Rz
znEZvff0PYWiKqNwNFAfumQUoYG3xka6MUk72g9XuMRSWOQ5eQq3a2GWGGU9tR7g
qCeIWR2TZDKwkkBaFxTYYbGEQiTDrLFbngpiseKAlHqYMFCxAvmPE4wFEpAQLkVj
ukLmczFUi4/6qNc25tl2u5GIpyLIbPz++cRAENMlCnZX8nuRnH0h+zSg6I6TXpWI
0WLeVACl5gmVSQjBvtPFQvJvHd3PWFiZMZ7WVuK3eL4pwPP4y4dFuAsPzw5PiQOO
fTeeSmp8v29HPQGIvZEbL0EN2HUHNfB6ILoUM+mmRxjgaerb0zwEfsrX7gljVObe
diG7VgTlOMza7VF7tvYL9zG2EyF1HlptgJUE0Pq6F7fXu11xyGlD7Yh26H5/u887
k/R7JCrCjjCBZss++xZ6nPfQa6yiCoVAUfR0+B5dnfhvOLW5Yizfb6t03M1fAXK5
AqrRyuG6Ny/hB8qEIJYw22HDs+zS+0xz/H70+oQnZRLYDQZCSLtKwXKZBjArIkKj
gMTVlVh23WKIeKcbOM6O2XiaQrDLAq5KXewgKooUn/C2WbAwE0moVUCyA7A7+kl+
nx3wNblmebIJRDxFrHkcP1cqO/S1pienHwdcT7q8FLUDJuv3n0J59DD+lloNR7RE
/u7nFVdcnN8TxoH7HKbB/85iWn+udx5LtXpoR+i+u6TXhogEFvY4teL0vawtsPc8
Ssv5UUM/44fhb1oIFBkUDzAqERrIJHOeRJ47a5akEMMuU1WN4E4iNnTmQyaeuIOH
CNqxW/rBHE6NXfSQbLueizd+c0nqgmhLDeIDTkUzw+Yzmes8f0RZAIccfeRYENhq
6K2Hsqynvo/1J1XfBQvNGjovA7R8quMYmc5jRsKiF2IVp2oXk24yZGdpZMlK980f
9XKrZNmpu7VnTUyXc4rJXd8xo/kHdYZdssSI9Fx7UXLpBtZKlrgmTyycyNwsQQIt
yKS0yUpVImZhJgPvj2g89zr3xfHzGPhJ7UUTaHRrgZZ/4Bto2udbochDSNZK1Jr5
gfE6Tj+twAJHSvyUjvVTHYXf5UwopbBfoy4aHNRMgDA1zSYKf2w8RMAmSzSCJTwj
0W/v0Jec5Z5Z9qsbj2uDywcBFuJlcuH9+bq0BGG4AxugdqplR0Q20R6Mjj+LveEZ
IJZJetDEM+1CKRzVnq4YofR0jXagO0qZ4MENO6/T3mKGgBsWyuvaB60pA+/UE9xt
gBUoDSSThdSZoWua6hT4EQqk/pyTQ7aKLLjkuViOCPmtgTNIZhFPpWz132b/S7rg
CvzipvG/jiJ2m0L0WB3jobwlEplytrbZ9hFNAuLYSZvRUhdJhKNREwq4cMWZJ3b7
SoDP0AkZKuNTsiRBQS9j0lGz0gtTeA49ugEQImSSC0nONwp7t0iEzSJUtmdF61Zd
IQYm3MgvMYhTGcqSNkZPjloJ++0D05ICrRkEYQcXW1MpLtget0LofgVFPKBOkMfL
EScnnrwG1PSt6ZiMZsl2FaoghVZCVfQJoPCkxpwD5/X4nShVUMcXMoDkQyfQDuZk
3MnBrmSnKgmcQMM6DnlpGOGCVO2RSamMBzyDRejsh51yr1h9bC2z+j0uEHZYujws
5peLL6D5iHVd6hEKUyZyestVyfoptnqSjNxEoIlTlho0+x0MdmkO5on9O+aLrKpH
pHlg7cgyMT9jlalUstO7g+h2e7Vnux7qxe7r0fkk3aALBrG4IXEic7ogDl2EsuO8
ID89K2el0J6mPMembeMQaVKPh78Gh1tx2vmjc/fneg2ch4nrcV3a+WB25cJ7wmps
QqkOZnj+Iq2/L9Xlx9NIdMwkQjOUri0W1llHqlgy5rmyBXHmwyYG8OH9SMDbprwg
p8TsKgKFZtO/Rgvbf2yh0raIgDQdNdmPDETLzZ3QTfVi+NZ8o9miQKekTE4YjZkP
yo96y1boKuEGXtLg7geOK1Xe2fgvmb2Dfrpqy3nwGhDMJKsfTZy1ocu28Ug6YEX/
5xkiVwv6C2XwmXngtNaOkQOAM/hxWAgeADLzokKWn2iDT9EQzSs/gnHtdFLfewyo
orcSZSR/iAkB2TvWEf6rm+UdYLGdODk5Pzyrihu3E/DY0ShjUlc1uHrWQeTuPSgu
lTsSNZK8UpAG3gwFaftvMr1vlqKAVekzMMoYBH2fBRK/YYxF0TXf2OKizT2DwT/J
/TQC1AyEedDi7Gw6J7mwTHpBHB51R6R3yuJVxfLr5Nj2akMwR2oyOfF6VGYhuPXp
Afled+OEhCWNMJSGPSh//kwhqqzMmKATaYJTaUtjtqN4KvvA5pSyZmMvAFzmg/SZ
7j/qKvc7rcQl/ki+IR7uUOcM4nlkY0lCV092mSOT6Vd7Ig6RogDC3Nhjo3/6UpjR
epjm39CcQddlUBqPg1Q/tcDTvsS94nnR6wdUeDDWAHgfz7rvI/9TvfimA7PAaPpb
PvAueAj8zzYr403yVU7DGdyebrhHcAEbJSvg92vPDwwoDB4dOXFjmluDYbEJGDQ1
vv3gCQo7h0fa8UM34mm+rzxESaaBYrr1LYxcjVcvhRvTN1V8t6Q6YcvEpy01UEFR
BNLegyvcnaE67G3ZEbEVBDi01mW3lVZjarxzA/xwR2qo5IV5bCbNf6OCce/ghvxW
CF4Ue860f2zrcA8cCV/oU9mBG1L81RQ2AtqX8Pvf9BnlfUkIdU1gMuIKoF9XU+C8
1wCmvn5Cex/rpuEZxHG0G+3vnV4wke41+PoOp+zlVxUS9a8poHz3QLY9geIlQXIP
jr17YGYyg1oCqQnisBGd4xyPLnWzE8W0fn/MUSw85/AgKZWtusn3BRhRlbQVw6RT
lo7XmDeoxbFakt4kt/Hatro80juUdAupSuovUJu8aJUm0TD6KJly4Zvk2JKDjYJw
yS9C7BFeWCgv2Le4shSD4MLuz97J5JzyRBoP48V8B51Kaxa4XFGPX2WDmfdBmN5k
NTtcZ2tKMTL1LoZiBLnJKDHW5VswmeOpdw9rX7kXFPEXp3J6vcCReCw8R+TsGo8q
jQ/uqXTFarmBsH+zfbB7lqXXqnPFbATfbFQBc56CGcoogl9z+Z/nAKBDeSPruTX9
rXoiIMFlswyPdTzOO+KV6LvP5AlHtWFZwDPgBH9hrQg9c+IiBJoC+6UoT5KwJPs6
yqF+T7uTJds141O+jawhQsodM2Ceo7mTg9oBvGlkvKcs3HVbjWt3mT5l17nS+Xnf
ompWAeAU2vVCbQdqkSCwp60MPg0SMQnN608ypLZ8zXpEnw+nFtX4bxZ45ZaF2zwo
WtxrRNv4/jLZRGj133WRfsowWodJRpcMTR1a7MNiapLRAQTUFNCfF8Lv4nB99K2o
WOAILJ7mvakO9qM2e7H2BY0ETz/HDCddQjRHQVaM3PlihHzl/4ti9DqOEvbjC0Qn
gB0s8FU7ZVafVuV7NP2RFoi+WrpPg90U6qnwar5EwztHmRQC6IW9v9wt3CC2uJRM
Yqfxkm2Bt/CLDpeEK9eN3n9o7D4XGn6xatrszeS5ZXWfGugr1YNvC+OQ9uu8+C1q
5VL/+6K6NxaAlnhOgI3anmX7UrnxMILN2nA/uIeyiPNP6NPr4OMwx9SP/mAiYyfz
ZGTyhm8fDVpdOibUHTeQ3u6N2dev0aqZfNO7TYQaSTQC1w8K4aTDKV/GV3dYP6HJ
f1I+bAbeVk2sQB4vmfiLzYJ638ZokfA06MRDb64WtP4FsIfIpg2JP2sbgJdeRyxe
WXmvU517ck95rS7dnOxiNbOudmnxVLIydXHb/0H9edGZt7MlS8onjlKU9q8LIsKk
Lqy9jamO2rD+eLAcjTd6FSRRVaZqy0u/AXPEQEOIsjIZalv+rtEYZbp+NvqpNftV
shF5KTHl+h18IT1ZhJNwOkMJP6S/iSI2eaI4aX6j18r+JDmfggL6rlgYhIxTyvzJ
8c1gwgqtKgwoqyrL6XNKNcQsIgBsVv9e9O+3EO6y4mlcIIMH0GKtunPi64vcooR/
vTcECYkEVmF8APiXPaVNXIMZMUWNv8HSn/NWD33h4ekbGeuXQX1hPZM+newUCXrd
rbVAi6TUMTQoBUyyh3cNueCFt1igx9mfMkMa4XP2JbRH6mryIG/uZ9f5bsQSSowR
ell5aYU0F/OhUmYSNqtkGsgbp4zrhfDZBGtYp65Smaa5O5VYdfwpNTLBffM1ofnm
RdVMrVA5a0ho4mkrcRfw4hk1pwF7cC+pYC0ECP1jSNNCiw5/ePEey7iGHj+/+Q1y
ePk5/Gpo3LHlJmnx4ja2uf701ZWy/ile5YNlaGiz756p8pslLeE+66R8A5zSMWr9
Y2HF6Q5WLHuof8LX0HLRhjGf0MEEcOyzE05m8y4bg1S0eqbr0irMuofe04UAQ8gx
7NxanIb9fWPm52eeePQ+qcl8dFJW9/uzMys1dVlZdrelfZSHNPKOicEYFTPfdlTW
8OBwRNAOkhDsaYa+llCBd50ic5oF5tw54NzJdmkhVgqyWmQSW2i62AyiDnGrLaUj
eAWUD385DCAtkkqil5mu7lzlluYaZuH2a+pSjV5Fn6ZMPxpHXl5UInTDuk9j5GtJ
NWAg1LF9uNA2D+pb2k/SMuD+HHRuQQ46zWPfUAVujfui8PncaRkmz7mo9HHQwHlC
QYELFlBK1J1wRY+VTx4fZDYXfruti1pFcJWPkDLwTC26rHUVHOxUZGI9lciCS2W5
qRnd3lPR7AYKjG0uv4L1hW7/i5I1w+D1IrmRiN+TwzSrlNSpFy54rspUuQJFHpPz
s/u8LVkFQ/9nX/IASaNN1Ro6hhWrXGsPit+TQYRcsuRWwMQ5dUmZa0b+IOc3SrBd
rLKDiDnVsTGm3XleIuSQ0m6eNLlk6D+da0pupoGMxiEFIkZWoaEiKMv6blVat8BU
ckLE2QTNH8tu8d2xbNxnObgCOFX0JnbQAXW5hi8ZUZyRcGPOyQAIeuYzN+yM/bEC
r8Jutr7CPfZZszg3+Cpo2eErXKb0DIAzJZ9YhutgbabSlFvtGesXOLWYYT+iE7pe
aBwd8AitwFK/Lmkf6dORWFFCXycFhAS4QSB05iEvQQfK/bxUPXpYblAlslkAJNij
IcFOZChfr1w08qdsJma2yAHhsVy0C6/EwYJeFcvPuR0OtIapFatp4pvtqI5YncU4
swz+LIX8h0nfvqAipZNbzIM2hsc3CuwVKH3TACHIG3QCORUXCW+A8QL7cUdoSx+W
HqQSSFN8kXFuKwZyoTQVO1OsT6X4FA0DEa7pwMXXRC6tJNiNiap7ZYQzX8mEykBW
nJh5JHrTHl7SD8DncZjReO9llpbgm9GWsuErHzU7UDBkJsoDEJ+qe7y8yci5zeO2
9txWkVTJil4RRJbUBW30ooySjx1OgNMZjnwfGrv+mKnrTc/d28Kl//clCcgDQzPs
ygnzpo8GKqlFXgiMzFSji8uAFsjfJ2pqedNTuKb9oCCeuSx1Y7XWDuoLHf33fCRP
UplqRPi6NQiWoTon+17sfqjvHJ8Fyf6KCBNS2RGvdoQjVb7rX92IVZ5GXP8nPypk
V+dGwWKKQpsdaLPe2L+eGhv5OuiRQfUrhS5zzk57AotWNE+1HM63TdecvcigVTht
SfGHSEsmw1qBqK7z4uKdAWyTkzVo/DXmeTetkjYL87ARkBxoWs2p0Dnf/461AN+R
z9z+9RHBzdlQ0Lhox8d6US/mGv8BEMmFpYYOSXX3stg4w+PfVBc82kO9vbmCOdee
01RlvqalFLjfxz8XoinpFf5sLuAeZODW/GvLqTOrT4JAvYT0en8avkQ2CGJqEkXF
Tie+iy0ReKFTHI3g8uB04wRVu4BX0BsmO+P0sH8X2plV8QChrnOhC6gEjXHbYaPN
X3pfUiI2xDQDCCx2D/YKUNRPT4uVsl9uMqZ9VJHkmdQczlUzArWkb50m7hQ9pP0d
pXAwfAvYfauNhwoC4AUfkIohHgzMe+z+H8msucZyyhi6Pgvv+2oIuTXPXiGGqf6s
rYoOfqOR67I6yUTSb3fCP81/lSLzgFOOktEr/kw9X6lz7AFQLdN+tjKzcRHdvwdM
c0NVOZMkimUwMeZJLQQYzedR+jeCrDcYVINlkRXqoledEDbrw0QP4mJP4tm+aSWl
RX/dS9wVHQ+yyAbwLMjDnPSv8aoWYphRZuAZvvdUnqQa675ApSB85WHVqgdlwfrm
cByN91mWxAC4gxKAp85Ey5Iv+PilZYsD8QzC1xHilnGAQcpqJ16GWYdCwEJ5/hc/
oWyrlJWqrW/UjmHaVNjg/C24q1UbKweUfoFYWE4rJ/lY5k2+nOqCunmw4BF2B+EK
J/eTCq2srsAF4rkk/ar2K0yUQIHkP6Jmzb+VYRrb5rQI0w8bIYSwI+2RiukVnRAx
fn/gVUn956L+9+ippjxwA4RBcIMF6pboVhFQF68I6gW+EJCE2iqtJTdkYbCUO8kD
jn5LPcMQcX+sAdeDVbyjiAJnBz2gTh3sgfYJrBi76oxbYp4lW/OXqJ/2fWNszOZO
7MuZ2grKO88BtGwBqvc3j3j+X7gCLnPJ/XJvXn1irJ3IcXRFyIXvb3A3cfr2NaPm
slB4vjrkaAUFGWcm3RP/FCX+XOWYImeVMK5QSbTV7WEpw8HiK8ftvZZZ3rw4l7kp
NoSMm0lcV8EMkY2+Fr1vLVXoCCpR3SM5EoW5XIHhY+2aOL3P5+9y39s/mbqiyjnq
Kpgh1er5ynl0SW9kT7xugB3+Ks5UvLBiokpsEbSG3tXL+YoWZ0mTBkob93GZvMGj
6oGTn5pp0kPiSL4lPXMRbXZxQVQHhBIF4FLr80fRQtSI7ji+/0g5Kc8pMc4PShRG
R20Rq3Zbfsvaryba2MfXd1GubLDc6mcdbN6hBR4cdNEVfNhDxCrXDTCg31bU/hko
XtRXV6JwUrrkIE6yyle3oy1x8xM9mWFX/fQb5fNeUli4sElTr8ij1fXbViE8DaL0
boxE7gmol91n5rbeoiQOYVHrPixydXtUCOqQPYfYrKc8aQpurlO5v7UVXH5APGFM
KKXBLI8ncCHkXwc3hTIZVH8bh/hPh/KziTByxA+3qkAG/X4M4swY7OmR3caDVj1y
Qc6OJcBsk+9vJtdbm9sX0FAMAjf6Pd+F8HeRCNzTs737YUm1xaUWVd9emZJ6zFLk
SD0Nro3LdfFke8R2yUeZC40rujv5vTty92DuLazpw3zRabIOOox6a6SguC021kiM
T7I06KDbDNwvKvLRznFjgXclr58w3J0yhbokOhuaQGbqGQbNAzrR7AwjVO1zCqHU
adC7drmAEr/oHNDnvQH4jqcKrGSPS9kBSWyrk+gJF7cibw4OfulLbkDFAG0yhJ0U
oB6K/Fu0G0uaFU5Z+MHLKCq5YAMSaTs6JR69TtsyTTLIVQqn7+B9OJPdV1h02Wwg
f5ajmQzrSwLuDZAMsghti/Bc9mwny6FYhwWz0nFsUVaMHk/3UPRoRMpduIlcLp+U
7wjDXMb+E5PdvWTHkq7/nuNm2L7VTUr6uSIrpBqZaV61mhWYCvVXF3U87vZ92Ml8
LVTDdXwJlBt5c/PtQ9rYO/N/0IUcq/MGhr4yEaIQXXhoCsI/+NStfWI1Fs8JW5Sc
oQHMjWH+hC4sFR4okO7cFfio/6P8OBNIkSzOtD8i4U6vL/iepVfghv9WyNVq9PKv
IlrFVC4naLiAJTR51jf2faqHC300HZtv5czRCS9Rtd60Nh8bC6RHX1JuYNkYzU4V
IixN5mjkhAfJNeUKXmhc53mBph/ntQm/3es9zWs4c6hKC739VV9J0F0rJreUJOVn
v4Brxz0/zclPp4wd1MUrtfHmQBhLwhXi5eitklyNypbJtJc6KXYQqXe5JMgx43UI
bK0KusmKWLFFchIFCzcx+glxMNqZQXJ2DQ2lIQOzecORurIl7lKW087GkFE0LvyW
7fyCgjiv84QgSXcpaMjP/3wEI/ttbLytcYApyOWzrQut8so6nu2s1X6evpFjA8lV
23dIKkmzoqjL6+PbglTDKLnSSb4pX+vnBA8JK1tR/E36J2epK3emVDXYmHZA0P9g
IFNakzRd4z/z9+tZFMlVqWrKXtozVB31c/G1COX3nFzNhkW6Jz7l+2JHPHj85BlJ
hnI7AzRHBjFTVVry7wHnRX3tFwqcyQwdGXCLkLVv0b+6w3+WeIjmfRwOaxqZ+lvX
yaSpEUEeZgt1SSZAkwulM7JEWQ/0zsgsvrTDuKnJEqvqTt2rqYfQuyhQhGIM7Nli
jesLOxhKhnhZNleCnlej7L1XIxEhASA9KzMPHPuGggVzvjcxWh3IAxYCv9v6lYu7
cikoV7MX6/ZKQrRd5MsBK9kRGPOTR+EoDtP9NY2RDVF0eoYe1x6TIihjKaTCqvGQ
c2UoMb3PJCKxssszr7Vdc2ntd43raLzqybcGsvuzue/YvhBKck51Q9dqLrnY80ls
9p6olb1mMYBMDY0fhFL8IEUQSZc+O1srndxyLuFS6Vi854NhutrrnBFMVCvu7p+F
APOoESkbTWaoTqOT2ncnm6s4ZLYzE2PLj2hKKFiBSXgnU0ZpBAp0Q6YSV/JAO368
GXg+ib362tOsPsdhZ9Ckw4yGZh++exF8rDncnJrCkydZUC3M/2v83F5vdeD56rvU
WZY072gcETZV4mLMNsBTFJ/ZGHb7RX5TML+nn2jpM724+pIEf9EuWclaN7Q5B4mC
9HOSsG095zl9dFJBMRJCgDJtdG6UXhgfavKgoJPij2OAyB4O5Ud7YfD/NysDPfal
eLiGpDR+lr/tCCVCGbW04YPE27QITnR4fRGF/plXNBOeCvvswa1CpxxGMRRN7Mys
JzjmwGhoAPYg2g5ueWwPm04T3pa2+7CX6O9f//akfASgKcD+sldK6MGFZlUH+yhI
FgpatswD5agaMHvpTO+lLrWnwGQPfAfkl6LKGg8BKogOBpw4muid7jNdskSn7Qtf
oArIo2F1HaqAE0Co6adFfaU11gFzpl7hOrnQpx2YgtQou21pwSG94trzSjzcoB2N
WUrIkCBvW2UCh7SCX37WQPSsbVZvkL+VhqRNxd7b3NIYbTyZh57wbBZkD+fqx0si
3YnOYr2hpMRiMmuR+fLx4A8f6N6GulLOkYHeMnO5PgQN7+MOFHfIwxNj6MrjrIwg
3tbkv6ArVQZOmgLqDhI852r1pa9MpZ8xjXqtd2vUln1qN9wTFr86GnQbAaXOQZ1W
sLmgXpMdGg6oCq4x5h19QVLnG5hLGtfxWs6HeQBlBocE13UOCa7QTd1kNdI97co6
4TibRBVdkDIRqRvK5amqLR6t3jr7yHYN5ZIj1+mepcn6YsvaHUxNk7JN1VB9RmiI
4DrsdkIOL+6aGVm+SNfHS9fAakovUIIahnlKsvHL6ot1plWMyeeJ6Xf/gW6wkFMz
4dAwcd7iAqRwmxTGsFnvgjiEuaD47to2v8Y9EjiUISX/4af4y6OihwOhcuXJiziB
QC3ZohNbWFgy1hPSioJRSR2h0ZOdb9PHixDdC2o5uIUwz/1ngnL/JUUTEFrvbj5z
7I/kOErHoi8YRoiLNLE0bysV1DTlnan+i2EUy5cjVxEFXyD8Bcf/0q7O7u4Fgy5i
b1EGLFCUtVaIGd3iuzEqgNg8h9y6ar7N4fGopzA1at5dmAicujQrBI7h9rpo3RDh
nJPOy1ev/ADg+5LDrYQltqB/5MMUALYbE4pCCr5/8Om4TFUhHK0FAJ0Q2f2JQN0F
xRQFrihe5kC1Nv6aWlxzveqEplWmDupBWysByR61l6XNFBYY6YLNpA0rIJjd4ill
A84rHZXsECsNEFpIEbcI4TKU6Ghtnfe/7xqpfJeyyhybKjUZeXifyB7ituNbRLRE
a7UHxQLBwjKz0AbrJ5J69FGZF6gN/BI4f8gKBOs5KWTwTe/Uz2QmE4zLhpj+QZ3Y
Sa+aDGXZKzmwtK+9mPpFa9GA7fLTUQUuaQwK+JgcrNxY4Sj4nkVdpX3k2QQ2z5h2
p9Vo6APkN5H1Ql/XRzUf8LXcfRWOp7Lv9jajfydGdyJp5t5hLVpbdjhnFxJVElGX
ppOo1wsvdxWbo1eWppYUhv+E9cio7GR2PYrW6Apln+PbROdNBa0iOkliO8uXjADa
jf7a0YiVGmbN9aNf+AJp3X3sgY6k37VBA5zLUNGba9iI9bG0NITtwvlzmzUEqNSs
AgS4w0CkFff5yCjaAotIUGawgjjhEOMxvGtduzxnXD/0+SAvcys68jBLd+zs7bF5
LXtGJbToZGxzn25D+0ohZOzYhJJs/5E7QQD8ZTgzHQyptXbwhXqjm2MXHUdFl1f/
oD0VxMmzh0EJaSxDUxe9Crdu+aGDf1iN5wzr41StSVvPJXWgJlspdn98lujpIJ+C
SyKqH85YZzyfOHivmtMb/A2v38BE/ca/TiCqXHk0IWnMKmk1YGDAqOkd3JCjWCv1
7SKhMXogafG2QMfboc1vT3qKsqqqqFkSBPmQpitNOBAO5fjA+qmrSN/KA8dWcIAI
NQ82paMJpVYoEJNn0He0drnVGkZLp1/x0J282KCTSfvxHnWTvCFgbnZedbTi+q3u
+0h9QTcCR6s58UP8/mBSNyB6NjT8SO0j0r027uIN68jm5I9+1xnkJVIdwta8Ok9H
ha9K7UVVrhiv3449+R5iTxDfPVYW4CLssJxuaI0JEIEGJGWVcMcJcLtjfJcr5CEY
GgerRbTZh2DpMUN8q+FJee5FfuYGaUKhYOi9ycKuN3/T/WXiWtNyWke5w6NUKgBC
t890H2rJaWqFSqWliv9OS8OUO/Jdzi9hkIgoB41YBNDyAdYdrL65GPics/izDtGv
as5d1Gho2nAamO9vzrvJyDrsNcdIPTE0kw3u9LZUFHCoV+rKgWJkEgxn12jGJR8C
pfpQst/hhp0p+lHhtmF+G0yFRjnjMpL8mYQHeFSCDZVP9V9WxiEm/dTWJWq3s+Wr
H4iRWLwzcHniZ/0vDcPo0xza9skrzhUpBKM2r8a7O/tVkvwqKle+3AGuYWkybIM/
L8g5M1spPp5dB7M2GX/Px6dUyPHRZviwLarJdGd5v6p3m3Dvj5t2IqqubaxhMHTh
DBKknPiSn+UqhY4t5mmZvw+2qe2KTisRPOHA56hBdbYtL+aN2tdARRXTvXs5SnYF
ioVtWbVL+TU0HIr7Sv/4TfcHkKWSOx8E1zgfszNnzoSnbBE0sR4TzcJP8YOKtgte
evKskteaQA04v/yN9S28SUmmHd3ZSuwoVXMZqMfIabn8AaOvwKkFRaR8fATDg4HD
qgSD/lJiExc6wB9ZlFlR77WeF+S/NBW9Cob8wYd7Rx42h35VqBqo+qprZYqW8Qpy
oWGWxEHigTpHkL9An6WSaPWz8ytQXtay/qkbanDWLAEq3wWbDxOI/4ZSuuTGP15Z
SgvBs8KAKm3bz2CU8KCaHekl8fXFa2M7ADNim01Dnwkf2pot5TDQpdR9H390Qiz/
Dgj8/5oyQswuN36eSx9FDaNtTmIp1QpaP9OElZcjSy0d9F0J8LvdffofF0Mt8Y37
/LHNHbcPkGe1wyAwMYT3MMxXCUgk2WYjsJpEhUZbwLrTCz0fXMROp4+jUlBxZNCK
+GOJtHmozzT1UrqahsnhzodBaPC+M7HMJ05tfjuAD2eVEqAS8pNoL9OQM0k/o7+J
LH0jLOY/T/GxsqtkHS2RKO6d1vRNKH63FnkG7tebXtaUxQhLzou55l31Qej4xWGj
FqZ9zIR1+v5Hd8NohxQz3BY9GSS9/RYGgEg3rAsPfK2S+T9u7/YAPLIWbB6kAhRY
aBxkCvNaqXkG3bfVYBi0XZcklM+T5v4VTP5TYc91KIPpiBDxfZR0cqC50eqE0sT/
P+DE0QBo/c8dtOop4n552wU5Pd4LpKWKzItmS09TkNszNBl1vw1oNvwvOPp/xUNb
wpTQ0E4ZTtHmR4z7bYqM9j9VdeXJWJjumhd19NdJBCPU/96+rFSrx0Fuk0EOuYHD
JPOCDtSXpj+oLAxbRHGh/HqV3OelZRWadtNEuYfl6TuH6Zg7PycH+EErWclIhdj7
euCtMOl2o/pIdzyVhnJpAJBUKApexgBUgInmi9VTTQ+x399apVYzoTCmF9yLwCf/
J6xsmrV6zbG+SvOfM3HP5PfAlA8u3mR+e7jaxIweRzi0JLTJzd0Iayc+9t5WwKMg
FvH+QSKs8u8kSSDNG/Ye+2DUYOtj7HtV7VpfKTkCtusEtaGT9InDI1YrcpeuTxhl
cxo01temW4msM7R2F1XBjQ98FjzJjgUpn2r41YzoQVHamxXYaVot0A+4yNeOI0A1
qMzptbi3zaAFnSMaZliN4JURM+5fS7P4CFbabch5zGlScfx2ZsdEk8u3tQnq3nHN
Q3bYR9C+kenH05YRHUb4P585FWhqubTN2eIKpuKQV4EE1pAylEuMmlQ9U5So5VQC
3uKKORQcTH6Xl1W5Ml3qQwxdqRnqMLB6tjmZfFWxc83Rq4SS+lPf7xgbzTrF9oXk
lGIKvleV3cJt7uYvExCNRF8s2/iqm6TUlzDJLGze86+eVwqEf3z0pzmNVGA2pnLu
8n6wRoWfkPfl5hq9VcNkKYNwPLKPzLOzOEZAmxVVsQ0ayECiA/zmWBE+UKvSyzct
YSTPRY9t2cqzYOAVMNHDAIF0A7AVf3y5ED4W8zPfo7kh+8GHXijWEexn9OfoSSB+
HWuhRli+p7dpeESiI+rm6rOXOx00SalPrJ67wWIQiGpi+5eOxrSo2a/hpFmTwf92
0pr6mHItiSZIw2vucK3M6Yt/q0iuzgSKJlUxDE3WrLjOy/wahs1Yyh2KmScEFDRW
zA/BEQBM87RZnXaKP3RYCf4rsUoWCfYdBxtkHeyzyACtCz0BLcoSqOij7I1OITfk
r4BM4kwbqvIS8Hw/+t7seFbJfNBlWod6KfBxkDB3wegbQaMynNkCBwPgkVXMEJ5R
ogZUPdM37ZYHhAssMSkH8ipnYVqWiZQq64879R3Q9ZkFJYxqHDNqeCL4K69eK2zv
9B49z3iTBdwskSwSLWj5psEdRnUtJa2i50D8ofilFmLllWSBrXkDHOJxq2V2sUxp
zS4/xhngrswaKjs9rv/AnZ/T2jAd/Agq9itdkh8MCBeL6GNdYZxWKgUqGdesL5wZ
h/lnegbsYVJCCQKoGxrd4qDofUqfRgH6EroKBZ5ulHDMhTdkRge78TTj+344vm9f
R1+3OoUsZkcpw0Xdm9zKTMmq9MxUiIacK8gSij7Osjb4/60D8UHNyCyXfYl2F5h5
oUR9goiPW98+oxJR9H2J5u9pSV4By8+Ue3wzR9cabWoSDDbt9+jdlM62YtVofst8
0VajN0wRVftZa2wf+8oU4J1OtmG+MWXSql3R4SnGkTFvqNCivVvRC6LE3TDjsTY0
iyyzqQwaEP/hFT8mIYsPSCj/O+nmzuzHAbWkiK+79Sl4clqjn6+63qRGLykLT/pf
1khbTLhrn43Fn0GegMrKQlOZU87ZQMCkPXzNEdK+nwYJ4mcoDoQopzxqA6gUJ2/h
Et96a7Kdhn0y4ZM8Grx8IBc4+3OqMtYZkly1NQkrmYRQnFIncj6HNktr54R8mafn
nC1Q3wW5DgwjTEAgEcvOBGLzWH+WJUSHMSPBrLMJWjugJOHB9cwTE0R3axWSdsD1
kbbvAUwn66bJZS0/LQ6S4Lx6gtwlAgMtm1uykrPrL4ywVXU/ZLzJM/qiXVngVDAM
gh9eihfNhwkWOW75aEfgwxce1woBfbKn1+YXyth2tJsz0w30/9kx557uVc5qwvOP
l8mgXAZY1JzDYuucd8cCdYALVrjICqB+y4N+BtkL8vlrh4Yizg8J4Z3Syu9A4yO5
A4eIrR77Zx0kfA/zaxEWZgLg6zlfH2PMxTderKEUO14NSOezo0x/mb9AoIcW6iOh
PxfiXsaC9MF4buXMoCT+O9GuZGdUBcXVWsgPRXueFpLC1cNIXA1rFdU8IG99grg4
Kz+G5Q8qZakx+BfOzI/UUn2bbGfc3r8K5O6ISMuxMFpFFpcCvjJ1GGL3t38B/T7u
zZVuPbmJnMenpA/LIk7eYXwuN25hFOCI+gBrb9x+73eUA7XQChUX1hN1jvxtJq4L
+XWD1IBm4SWtW3bbl6LqLjI9YyBnwkt/vZMOYRwywtibuFyOEYlGaIF7LWGw07ap
MXsoJnn5/PN0Ueaj2Fy99qjdaXRk4sQh2DNlvu9QsXgrlCUR53WLri+uv01T5uRm
z5u3AVxWcS7pBNB5HW5cNY+qNXyWI1OFKowuSIWN5pWhvonEdtVXf2kAJd8HbWfF
pqJlvGuu8fNa9dnnl73KjISZQTkuH8vkh/OZg5JNA5IzHqo4mZG5MbfkCDQu9G/H
Y1o5hDvC+9B20U8vLGTSZVgJaojcWVhRyZsrIfYfio6hp++A1rE0wcSsm5ul0v7u
/g181jIU+OhOkrqU2aIrEYjvtgT4/NV0rSFlIGXWmFs7WPbfyd0Z6KHPgXfhJGol
bfIcbprw3Z3lFeFUTuhlty3EqYuPBwc4FmQs4CjAbzb7aDHKWiUPwdwIhpxBVRAG
DKPis57MWFeQBlKLyyk2wjkIleVPOU2WVIHlkpqrjGGxVAmpMdLyebdsNfPX5eJW
H8ZjQIUr8IU9nwBbi99oV9B5ip3xwQbt9kWNfGt2PalhPOleQe+FLF8XsttCZNtH
qjMiDw50isegVLGo4l/K/YBsoYsw+9ZK9yP6spne0zwFVw4bso+x+fJhETKeBXDg
6kzkDRBdJ9peOKakFkbdB0MkQWQ4DaOZpWpKtnnf++htLd395jIJ9Zv5NqK7Tx2F
6rCWOCGXBFfrjqAPQJq/+wEcbqQdwOPUxn8rG05OnVqbUQ9u50rmtxUTps9kKvjk
IpnWOkbIWex+MyqkKSQmhChEWApgzkaLu0lbRl8uKnZFqtAtJPODutqdEfsMTF6E
NjmiFFpV6mO3Hp+vRL4naar10Bv3iT5Bg4eHXmE9WrcA4GhHidLqj2/wUs+Lj7yI
M7Bexd1UkVJXuehlZ19J4xB3eTJDMwBM7E0xFBzDT5v8gisimC4e3tPMTs9ahQF6
Bp8CooaMrSHPHegHWW/EMK5pns6G1HFvApyUJDI+kkLR613WkyvRm6jqH/t6q286
8HZMIEsabqFX4igaO3Etwc0jnqM5Zj+ZGvlX02sfUpq+6uyoc5+MGea/fbC9UC3K
imizGd4vyhkfAX3lgbtJlgZaRiCMEi31LO8PiYJQj8EjGUlBBthsgoATzj7ekcY3
aLKVenFr2DEisxTKKy/JDnxHjHycT93YBZ/+0fHnzYNzyt7JI9sFGyGhQJEvekFN
ofht9A0G+HnyRZpxkbTs8UBBXXsjyuOxBgwXmTLHj9rGCvwSPEQ1ydz4wn3SvnIC
QCo2DPOYvXWIg1o7ZraxA7vmdv58WLz/ppno/uQt+IZG2DAqXiryk1WtVo+BLwCs
KeWsJPfelnD3tqnzJ9ZiWSJVKETDnlLDc6HRCs8IJQI/+W3FYk4mTRKxxboNnBh4
mjdFT07EAdNk0NZrWMc2BRJmcgZzp7Hk9q9pPHKmZbmqyY6+XVcnMm7O+T1hK6d3
o60GLsjDj3S9VFQn3lL8aeGcgZFNeVPQ+6ixG6BLRfGqh/YXp8j9I/3jBW4ajxhu
VFrZFOhEcDtYGLXMQzo/zRIVa6LOcQGp9plCyihT0wsEfs+yDqQ2vJtxkOCyjyCQ
043J7B0klbMmEF117ZXtV/narmP8sRiHxP2N6lDL+FAuDKlkOGkuLFEbRRxBZz4l
GkVyQyxfiJ1/RkwmiTiq6qz7FdEd4eg13JWUY8Y+f6EkBIZjRzPasPY7ChHW8siM
oeH6pwPkhySbI2ffHnNaCNsoGqLA7tpZlJ/PCZm07T81g7lKgHz7v8poRDSmLUv1
voKnkqPAa4W3tca9AodLdS4dwuO6JzxKsb1geJsmWQ8kQ5Sar5PbeqbzTDSYf6vV
+Fl5Ks86VpEtf9Hvv+PGaBWO3buKou0RXWlmKh3DzyAu1+C/FkPGqlq26vJGTBot
GnA+bzAPgBhLeN7pjYy07hqm91s24LCpRKuzTn/MnGrf10S0nP8CNUL5tPtjAuvh
fZv+c6yb0rmZuMAZ0cobzw+rtBbTLEq9VFu9EKIr9S1x/lTPqwcI3Gfyd0y9r5ND
lkootD/v5oYMzQZ3tGC/O0EM8yhDTuUUgaxIwUiSO3/ecz65/sMfIxoPCWO82Kpm
fBVQKfBqQS4wH/Y2gyxYN2ts0cF/kwRwuqaPUhquCYOerEWF3TmZFDpSz5CgbUJ0
jpA/AflW1X1Z1DA8hAjisSa27DLh/NplNhgLes6gTbR7knZP6yl0QKHIRyTWoVL0
1sVafaX6wf7roon8XnWpqgEiK2Hzawk4yRkLKpAVGOz9/phXcV1JZOmBC00WwpGM
S5lOB6WFJLV4XVVH8obKNhRmXGkTUbROZDiKpXDbbg8H+cyIvCz6ccrLR4tI8CwY
RLXh7O8kGlsfYQJsJbWi10NRq12CLIVq8CtWfqjO+cCj2PizoxeCMcMXGiWQefe7
jzGQRZy7EgPyUHcH1rnLVmdKmn2uFtJ1BVflmWBbWR+bshx122Hba8cEH4y83wr8
dYStY6zDig+qU6kCfn1SChiLbjsAx6xsbV7CW/RxhHPFcGyLxpj3CwDitqL4cmGl
FnjOFtAGVDeJruOBlr0Hn5aV6Jale8txtbl+RMzqasHUfS57cROy1ZdqHPFbdJva
bEkxx+1QbfXMihuT7lUm7OI5HbwmVi2SZnnWKXoaNqWOVVvD69nJB6dI0CyjZYjS
Yac3rBtYCvjMjMg3EwI4aHhpzL+offVz4MJ4xVWpcrRqrmmp7LYegOLMWK0uBxau
NFvuPjIaXFio8pTLxUAa+6qHZHUvgMvZ4qVJvr/KSngawI769g2Xq0BV4iodRNOu
XX6rLN+216NJNiRnb3TF29XXiUNrY5R5RLOIl+JuZ/cR1mHdtxl0F3cpNyIpupTp
ChGEzdMjPIb1Pg7B9MpW/8lL4M0Ans/UL458wwejSa464W8Pv51b+QPRxJ2PKvFA
8JL2WP+3cdhtMF/FHnG+rRoEGt444uH6FPiIKoAN3WnMyR/VI2baTlt8EUb0/FwM
83NsIR2UDfGrBMOySYSLyFrIU/2o7217iD0uecGAwmx6aVAI9Pdft9x00GPKzRj1
plG0EkyxCfZtLgatYtvR/9ufNHi07zIpSfTw1/zxvR+uVIwXjKVCnVHsNlGpQXpE
dSpK0UuhDC+CmYyTOJAd8rzopDtdQrCiAKshyLsfsZd5f53/B8o2Ij84AiAz/w9P
RfPxou/AefDWkdGXy1WDQU5XZNb8AhcYCUVjv7mMpL4D8U5LExUzvuv1HHZIujZ4
NdKqAwzd4k1uyJaCwKdaIdgRWOyD7CXQGS9/DP4YxFrvxD7DerfcPGtioU6FBJbL
fLVOWVZEWIQFFj/CRpzVFKVriQbiBPfEXM7oBApu6lMyZcabVaw3bVb0s+9GH0FT
khDI3rQtz7gqgVGi/JysC6sKS9s/lkeX9/k4I37sd9QhU2QvXAWMaw643fY+frgh
agLo3nHu8v+KISKKQ5onImRl9H+UGnbs2LsELU1+tBJJrruZ8mR1F/p6n8behoc5
1VHWoS2U4D8D1JW+lZeQ46ftIsQyhw7nmG7QOTAhWBHUhkuKQ8J5Abbg+iyTY2IT
Ph7TUIiE/Jy6gqolVbvkE63ukM9p/dIwDMkoh9mNHsMPVTbz59GEJ3fRRo5GG/5i
NjIOrSpmwB+TC1nmu6wNo1cTuBYVFYEy5wIPl7sAQbh3tT56kHdK0l51WnFIyzHl
GVGo0FhrsaSUi0TatyMGBd/qmjbcabHqv8iuQ2s4EkV5I6OXfVJEAKfjJnKaNPrA
of9iyhgdKNIrtv6f3EgwMs6cVtIQLXBtr33309R0z4UHoY8TNx+Jtwxv78pLR5NI
1R2aOs/kiunJ+h856NRQPRW9/P3R8HupqRPGhXPjRBESPcqIud5L0xLxNUZ2L3Lj
HxR2QCkcah3zayqM2cnqq0VzeTgxOeDsP9sxUAM3/OrmcpHAq58oV+cF7Zx85RRD
PpnTR6HoAFUBS+mU/Q9djqP4WPwg3y0SUP58cK9X2tUmuSrABBWtUYwqUKqUUore
WiJb0edC7P0au+U4gop12ptrKchmPqjG4avyzUhT/TojhKLIMpZuVP3YWP8V0Psu
aeY5gT+UPlj1f1SIftHZeBRRMUmhs/YVqkVTlM2aoaqQ2lavI1Mifko8KURzKnfU
gBYkQB+6hWj3zx9vgZVg95gG1cZSUpr02yPoQ3kHrFIJLuP34uLUxq46y0oQ1pnQ
Jsa6A84L5/TU71V8Km8pRBIzp8wHE+Fs2XD0CsV7v6YgCWhmy9+grqzSUaFFLDHJ
lA37YykMz3F7rO9A1R0XOqL8aF/L7txCNsL5of6n78Oz5ZSPj5JksSltpzA072YA
HNxXruyYR1tPaSDOjvPFrI09a1H5jHzbB8u//e5ZVM8SNSUUHLxNMLVc25JLRYv3
/WEmofDpCmGWozHkFCbB4nYlEdbnAX2tXgD0QwYg2J39TD5XQEElS9H8hEd5UDaq
YRmR6b9JLhYZ4znsqxJ1A4NmBRIr5LD7mO2naUK7I0Dzt0LCf/u9k7jNbkCQ8A8Q
sOL5iXeuv+bCAHqzr85SPkx0pGhvy+5Upy4qQZTXWuvqCGYsSK1fd5vTRssplb3X
cbBJRgpeIGoCrCvxRXRsilt3cdzdGGCoJms0T7cnBcAFRwLYw2FWntmO/98zZgc1
Iwczwr+96Mf7c9wLMrBt/DGXc/FxanVRBE+XsyJicqOGCG7olozeecLxW9R/NBBw
TFHACgwEF/ao4lm2leoJxwtwcdl+AaaPU94jLLWPWvZyw9DNuhx7RERq01l2hFrs
VuNnvB/YHpQFPMlhmJ4zbLEb++bdj3QFJVDj/aZ1gSHN2nbv4tFLbOexUBuQKAqt
nH1QJai0G9CCJq8ZR/6YBPF8iwLWwxNyPQx/BsIGXZVgzfZURDBY57mRfVu7YFiB
0li7pGvEuf0392cmXjyAJNCM5hGaViyo03ieM/DXyaXcgxxUfT9DeilsSOQGCN7d
S3uag+vRO76YEbJAuBewoiBynlwa3ZGT7zIO+bV3jbrpOmkkbIWebtdZJZSshe1u
TVwTIOTo5dPOdDcFbZkthYuatmFZp6CuBSvPoxqz5d11II9J3Xempyt0ROOFCC3H
plNlDyrhu1q1pTn/yTrUjmtEnZUgQD4krc5glx8BUfAMDkXOp7HWmfBmZMWgdGQp
6zeYUeN8c6BndJSs6nGBsY2YslTPByzjOHN6v3gTG4oN8svqYBdaQwGlnY4dbKPM
2xkDJilBPKhp0WnU6TnnO7gPHcSmRPEZMSKLIomUNjXl0PWXIn3IJAjPWaJU9Up6
j/Zd0JvSXQW2UVepC80Rzf5eyM66MuNXKZG1iJrKkj8ETbGo5CyH7Czr6zJynGkJ
NkuCs3yTZuMK4NFruygAsAGEaH0zyr2VO1K6KIy0/YThP0jyaEXdbYA6e7apW8tU
wsftX3Ut69J0oakmKCLtrNwKUu1X4FHPbkKlURnXTHptQxngKK7Fre+f/iYg0ekt
8c51O3e7/7KtVtqdsq0R7U+NoQ597u4md3yCtzd/+xFIweWnAe79+k8ZGQ9noL3h
nZSERhHO+zRICg9k6wVCPrjQty6m25R9g4DxdqRbMSNu6wfbhgFqUAtcfnqvrqlH
7XYViaaQ3Ffj/HPJwXSQMc1k9x37i7lfzbdmJSjmxYWNmPLpR5yPKeYCOdUyT2qj
heIoF38W170qFIYJtkTl1JJf/wFTXuuHk0EoAkYLDiQs3yQO5RwNz6WbFExXw48g
g0lKuqaQFDkoZqpniJBiinvF3JCxvhD6Hspu9BmUKo5/Uw+I3B0Vw6BMpfs/h0gC
bEWBReOnt/s555r3gRVrsc9tDAyWTVd7ZV3zV3KNZI6SVzK6WiF+cGHe8MJQRzMz
czom3ysSoEX2uEB3C+ro9Eoh70E9L4azBPCNyPoVUDMZWOIYPfy5BuuOV6ab2Yk4
QN5LKvlXYbrHdrUVxlraCmQZVM2Bl8ID0Ne5ImwkJwT+aODSHz/tdluMDJ2lMSwY
fWC7pwb0tGlt6hyy8Np3Yq6y4eWwEtPSqK4R2tWEDl1L94dsudjomylsj5cohamK
iX75nk8OlrMrfc8CAc95l0PgnYwNwdjvQ87QcnP9+ilwnd1SS8JdqlvUs8nqd/fO
mSvXXxiL2aOfjHzNvHfkklhxxSyKZsQ16dNi1c0FKP30Csp3jrGkcQj+iu16WZCn
+SherNPnuFNW65Q36vEMq71/FDUJp58tZ/x+vYz+6waqOSykTyIjKAScAWpWQgcZ
7FK7S2rqb2Rk6aTUaaIBZVuSnmNN0qKBdrTTm+qBNuZGK5ZcXuMpt0FzZ3eVLXkI
qjF9nijxxjKe8cSerKG7Z+bAPZkY23R4U9biatbB0KsUF7IBV47H0OVdicaDYVnT
HtUyAI6a1UnjKxhRgT0czyKxbu27X1kA4OiH3FSI6sAtAz9nY0lZ+/6zCboKI+hg
X7fG53YEH3RiberpedsqcmI7bK3LoFpMFGPSL98VKL7DGcafNeJgZsNsG07MKlUH
Sw6w9WelZEwxONO8f+bh7EpcdRcnGps1CgXTSbZTqOphGweWFL3FFM/Mm58ZpxUT
kgd8cr7PKNoLZsU0FKvR8eZpqOmaRuIVbPFDFjMe1UVHch+jvFMTRLytvjtyg4Cd
j0WPZFM3Ecd5323zb9Jw8MR00rOQZoozQwPCqy/rl2ao1Cp9TVF1qpTEf+HoRClV
DTxyeBzWpeQA+WJ8jqWqgwwsFtUF3wA7Gmy79+KfC9jPwtW85A+mChWlQHUsnQLO
yGKS4YZHp23wkZk+Q3wwMLq7pRBA06E4lQxqNwT3Y3aLYQIrrrdzx5ZFC/wKWdhy
v8DK4KxG5SyZhLE3IV2m2awNzpjAqIu33Koyz7LZbZ8xb7aci7/77JMPBt7HauD3
DLiwFktVvoAamaqZCTyNRiKe3xN0TqJWPxlMeR0c18O2Mgig5zvhXzNN9z9X2uIZ
OLQyh/FDJIlqw13T0i6TXt+88GfWm37mjULpX72UGFXmYKj/Q43grxYk1m2Zvjdh
Un22TCLVYM+sr1wpbLU5gKxhcl0ne3q+3+1ZZXw8YTym5AMjBJENaoa4ai1dLXTX
8Cf+Yv8rAsZnOVuxzZnsPxtWs1o1xHBeNPqImq8bykRNo0yLQvNOOPSxxrlsR4G0
QsWcLcTvNs/EPshsATBWc4ils8LQqdyvggq+V20X0D2G7vOuOkbR4uqM2wlHO2ru
/jU+7WrNwT+qr8DUD7XQL4cpG2WiHXXVWs00WRLJ+m8ThndgdI1QDs+Fe9Wwtn/p
2koBDmtFksmxrFJj6LdonnwuLMGQ4ZfxlDYt1vNu3O4xLebf2WLNVkcb1vD/qsC1
esONaEX6fKricQ6QU0bt9oSkoJf9oMRsVH16KKVTzqhD6gAl6yB3KxxvQOevujUE
OtOc7uGVPliCjtHGbvAcCz+uZIYRTFIDj2lGoFZABAfaB8wdzFXRDmpJEPv+mDs4
oZbsb0hPzqoPe+jMwx0y9TAigFzjUWtV0Lswe9woyoWHBrIoCDb4lgwBJ376wt7M
Jqcd77DsTGjDtWgr82IBSqTPp2M6D0uY2sFM6yvtVNxwLUJ7T1JTbHYdC3qM+1EO
SHdo3q7mo2an9DqMVZaPcGrTDkpQQ/GtmJMtR1zTjMEkKtNn901YSpPn3u4s2vij
3p7bhlfd8Oub2mk1+qVjS6Sz6wYelJXMSMovNAz5GkSj0GpPURCY+3nRseETu4Fu
xBwvjRzENq+hvCiTelhqcdevZzzddza6BxtXPV8Eo2u7lT93+QkoWgNMlkEtPUXg
VHPgleoO8w+OuWv7hD6ARlVI5w1kxqUrlZcnWjkzUCw8yF5AsJ3+7U6+Arf5svUC
EsUFS1g2kq+x3475rFakr9ujkewB69atnynubohXFv5nFCgitW9AEw96EVnw0WqX
SGESFnZSHOFyqzUW/0U6igVsI8OX4x/zUkzV1AfvtvbCaCrOfRqYC+z3Z79kzhuL
YXgFbXXrRueKbQVsKgtL9hhpmodrULSHP7zKrv612ShFeUZtnVC4Sc3GJWstrovE
46bzt96KkgRS1I/ezu886rGbCshXsNs5GfC6eOxC0k/6NemkUKEkGMG/Vrb2TeN/
1ebI7azPOAc4TFtoK40ApGXB1OpiPTSuIr0GwxVhsowJy+nilPG+GdSkTVxXJtr2
ump89kMt9ILfbpxEMO+/YyOpIaNw2h4f9yySGafq1iSKrj8R09UH8v6ExbhS4ZmR
ZfdlDiZ2PX50Q/N1Jz76kVij51pUZSk11+0Q6AjL4ALxJWncfB7hyam3yGMVKX70
1xEsQxsuEdixi3mwHFfDxtwCG/A7UjYDdZxHq7qnA3AYMUio8fvxKgsjc8EV//Qk
kovzHw/3S827Y7KDBO2YzMO2Zvo9bf2/MOkUlivKibuBKuietXxYHTTNmUKWhjiu
XOqralJK6LS+PPUpdA5r6l3H6gWWNa5mPTCDZctehOng6wDViupt3SBxCqIg476a
RZehicZP5zghhzPZur4EW+tN7IQkrR+awoyncjhybl+AAcli/tvk3uTnY2+pxUAe
rSw4O512ltbCe2PmrY3wnHUVJgj9oVlndBE4qBH7FVt0va3SUmOO8bQBMVBnLvA+
RIL/SPXTyx63Zr4MpN63FI9+emyXv5V+sdwVvXtBd7LsvnOQ+ZPS/IRKvTvAikLF
lutqfmRWRv6DGvmqhgViaGjQqoHKOJiLOOBZCv3+T+TOe8wAvYtwXlYroV30r28V
y9FeI//QN7Mt/wwDp1fUr3VBX0Wb0lTkVfv0OrQ+NU6ayhAGKb5GRCUgRjVDrN4S
KaEBS5IOOHnNGcFwLijMDzyMH8gFSk3FNEbRdIbxqF5JG8WvciPQi8ZwWMISUcVv
JwzNHj7cdWeJSJDwExfToB8jEs7wAdDnc3Tx9LBf+puyClg+NqGO+yjhI7+kYNC6
4tA5OpAKtIxi52FFAfLTzAiM+JLs40Q9mJfIyaKBuUf90INse0cmqbHq/H7q1VjH
8wbjJ08SWCL8kAKU2kwXK5zOnH4qtK473WyPy7GQBZd3856xrr3S/82ZXTWbudbY
Hbv0Yixao+mV7lueW9GDX4Sq2dL3ttcxJ5/FStKTZTDShju/vkFHFYtfSsNaN72c
tdqjbpFmCzJPORKRYcV3vTkEC2ZIC51vqtYGZVpkjYY2h/+bSihxnZqHgDXapira
C7LGbdYX/1uwieO6DorGnkv5lsWkUBrQACl14MUypWhXdtyIAINWwXKMgo4fUCGn
lCyjDOkcrfZ6gd6+ti3/grL0XBQUYN7NHsykfufpM7J2HvNAEoTDE/Rql8ocAc3K
XSinr8ym7K5lIcHW10InXfD58E616rQije9hyn+uISN9EVho4VzNaPMfbfASuQMH
U/Zbat7eIC6QxyX/8aoBr3cmU8RlZq5NDBfRDXnHzwROMUGKTYnF4gP/mZCOcunZ
qBWq3C7bo3Ja2HRsNSn+OvAX2EtsXaWfk5afzAxY84I8EiehhVpBWvez3GYBH7aD
BSgshb1qox11/iuQiRsnEAxwXb+5tuqfix5C8pzWvzil31RtK+Y4l/qFsySMUunH
soGwkAt4U5V6cI1CLsAs4Ywh9BDlJQBdLoT3XL+tZfR+jyiHqNot2nckK6Zb5DsW
ygWFnSUcEI+veXcA5x/TtTyry15kMDMcd9WBbCLisFl6mjvNbKKNBQT+u2+yvvDv
pCqVK7aw80IMdFu2jJQ7jjWtTiegUd2fiJr5tA9VeV0OtvNhsMEYLDfCXpLf/T0t
bX5DSmbJrDtfZDaTUzs85YtCl0ItY9toTTY0NK/dwtX/ZIHzrNUsf0MhFPPhw6Tq
nwPpZChHlqnjfotpoY/Ld6S4CoHd5mA07CxTwi9nUnMXm1Nqmgr9lZYhwdYYL2t5
ZPg0n1NjwAEo/PdpzhRR3gSMEQDQb7AN+1mroV1lglo1bg4sYPV42BV0t4Sn/ZEh
nORUogCDHn5JOfCsWCqZPeC/1pOl+gK0ivEjLoWdEYJOG+C7RWqZwFjzOJLXTe5o
NsAXbksUjhk3hKb1TLR+1KPW1FswjDo1CcU4b9tAjakGH5caSpfYkys3Bc5DlTmS
DN6bV8VBpuLxSjNdIT9m8XvCYxpQ60UcIxK5Soctb2yHqJwm68q/EUkkdktG6Wq3
53m+n6aTPnEPurjToQMkOBlr65J2o5kL0y2CkT9kYh1MpHYJSegUc0+5y8XdeZJf
3X1LTSt4vLy8N9NJKNWJQoI7sfKtTgInEKqUJK/bB5CYQt/t4tmsDDBqr3dHdxMW
HgkG6LRyW7eyli1QI23JvT9B15kwXtXeoRo6CPpppRxX2irqlA1QFPA2rJmOS6ST
DH3nXW2filgAWULD7R/tLM1O/fhPp062Y5lpg9/qTkwaLxQCqT8TSG1SDbIfBenr
ZvIuoIDX3rZkLwMe1OhBpP8xoaiAzQPrhlh8XVFyu4aFY6CYC53T4rRbJ5j5k4Vl
XlsELwXMXtx5O+ZqLAjQUR1SptTTJ9Xef/nVdO7WYj/rTwBkgiLWqakndEwKj7tA
M44/ovG0g6ReBwzfw1EQ5t0hjfX0zNvHeM+kOUAUm0wS5iOFRPmDHuPJ7keFMZJU
J2Psw1ZCZLf4M4zVhKAXaPJQjUYMDIwrTZAOXRFDIihSjE5qEAsXqJs4I4lw/R16
PQLyngHuUCP4rnvf6fkVe0vwqprHiFC7NlCvd2MycTPeVqSL/a4YX/5Eqk0r06qX
+4Zz43CjOWp1mZPpdSB6ssmkV38aINNENibzsPcWOTqbggtYAElI+y5uplx6Sx5V
Ix1DOX9rC7eH9zNRp0foizLoq2KoBXFvbpAxdoMLuLj2sYp6njKZSNunVxWhioN4
0LeT0nmrGpbA2b3lEoWm6xn26exzE2oe6EmJq44S3vZu5M9inedE36IJU907GvEN
4GrYYIbKRhCksF06xAoriMA6wR3u8H+eBdrrXC6oBiKzZVoyPDVBHNXNd93z0BrS
TVVNl3Qk98EfJLYusSt7NcseCjZdBxIKj+rHhiRl/WUMR34nVuNtSAb/pmw9MgYJ
MYHB1W6IGqJD6yGqZvY/USC3zYBwyI1R4aJeRfO7hCnuIlHcKghc6Ua/U8wY3npN
AIJCW4DjFJt8GoIo9ZM+auEm39ywm0s0BTIhL+e/lOvz5zW2Ml+jxboeU9NjHfGo
lTFIkI81kfWsP1EpzsajJ0Y3qO/+ZSg5kZY2McQZd4DtZpmQWL0umgrAIH+GxBCf
BMezWul1mYu4aeL+NK3qf6hB1Tar+LEzkScu9O9Vmu+iw/y1rp8CYN7+NDxAcTvd
XQgOFdhwNZTxJe9XpkeOCxAcbku8F0huPfaZ+m0dLtKmjMMAmlM7ChICyyJjyOMv
+L9q3GTqT8yglwS4hP33NM6OcUjfBgU1h2p0epzenqr5VoN19zodd16xfq4dknBC
92uKRp4cELKnDWnlGAhoV9aZH+6eGzBHtRiOZ+QiJBAtw++DEtOkJxPOrfWrFIou
puNc8gP8nozMmmAYLehYvKPS2SxuBxl9bwnyb/jotvKVcLMCm6hxMxbmYvXyC0aA
qwcSnuHEE5CqEOOUk7TqGyoKw8UxEmHptzCAw+Ss+2wuTfKrczuAZ+SNhL86Xvnv
7dkTeL82ew7m4z9b9SN4xtlKy0IQkTMqz1a2QCsUc7bzIGZANwbtwdfTxov3qRtv
adN7L8IZEeor2dVm8tDuAAsEn2rV1X3my0yhuO3wvyd1nIqgYnL5ArJzDWBml6uA
wyzYpJURstZuO9U6Sl9ZBau8ihlKzTfne8BbTPgsvXufbRotgqasM8bludD7O5+4
VwyrLs+c+brZRFD6xfN/m97Q1BmIyNeWw1fhQjW3AKczV9Wgk+70+mMw+k1JR0gu
KG+PqOB+8C404uyYh50psyEVHhjJ8qFO60swP05aqH4CNTfg+MJLt6VVdtm8wadL
3oo9SZWpoUNGmgCWIzvsLFXfCwDXc48jnjrPoIC0LmdXUFYnRPI/7oW3lU4Dugmc
osMrA8Qp67Pe/+ue0jnAqACtGSYhHiqYkel9ueuFTNmPC4yKi5XUWLJ5bL9S/AB6
rilbydlZG45e9QizitoZIu6kzWDlOz86FTPAvIjX4/+MDjBJkUbTpmehv7nwmD3n
bWDwFY3v9QS8lDEQok5Bagh6yLPkSeHIDLdg0LZas/+sr2I4reipQv9dgPqnAtiM
DqDMsJ4rLCo7ek2u6cn962GmgEko7Q+bth/NA4ZZiB1fOZVyZxtThTjIdiBynWCn
C64BRJB6zEC9V96RyG30Q5JC/fI6fhkZBctav09/RJiBFJoQEmSHdArzdWs3Kh2d
k295OrNBPS+WeDcw1uU3QhHG256Wq4iWW6OP7RPiAeSlhLHVqA7UrbxU9fOLOFmA
Y3h60+bfrOfxpaJmdZXqgVDG0Xfyj6gt0Es3WwELffD1cm+rWRGM0vq4/a9JmsnF
ijsP+LltxCC5vOuplbZ+tT96036rqN+EDPDyKmSVG1PIyfkV/D62gtqZDY8duI/Y
dk8Id+2pMYI8s4JVoW5EpV7DWkvAPF2yRSOVRj0q36cV/eGKzAmwsPDIjBzJK12n
G9/dTElxQW+F/FM3D+F8rm9z1YdAwvp0xHzKxG0JPpkCNnDI9RncVT41L/D3WRmx
qKw/U5TTYVdrPVtznZYh7gFXULD86jm216mQZz9AUM/oRWcKpHdbri/qJa46S/R2
Bscvxgz99rwAJSwXs8+FV45BTvHHWVcUTFKNYs7Skf8aFBG47nc/OgQaLULb+WzP
28oiGLhADnE0XRxx2GfJAwd/HtngoGLJSdUxXHcEY6dXKZQOaoB/gS3UMtpCGyUK
mm1RFgbrE/5WYq7hBFzKfYQKB5PeRHEkbSOr6kYHmxIvZzYkwqbiPNL3AOx1Uaiy
3FFAht1/xakePo+hJoK9kt34mKGMQXs1aRDdELroaXChj9el178myAPzcFr2liW0
dkeuNfYg0zQbf5PzsW3fkoqNUjNu+4M9wXmFXM0HUZ/Cfta8vowpEhbWRJfj52tQ
wo3xo3q+JEXMYvgOTk9GmAkpqxyOcKrplyLmaAPQAQ0UFEx8nPlyIDZkp9vmk0Sd
Kh6aG+s//NrljE+pGRC30FbQSukbmB6jK5r8aVwweF9HYvjur8O5zlbremppEqFK
vaNE+62VA5tF2qnJJHziHQXjSErOsY9VJVsIuSMqlXHS5RYBtpQSbCp7t1Vas33i
Fze2MxJaVzMc3q1nE3VuJ9THKXbu3IPFvVMxIb2RUIBjHWwee6bks5zkgbAmzqRZ
3v1ITFUx3VtlRrIbwpj7w76ryxnV7aF9ZOfPwVwRcu4iHU32cNcr1wL6e4oMImIy
6ZJliWFaxiIKzvVN6y9IXWwXCSZHCb9XZIlgNDR+DpADUGwwmTcnUTRpGkByi7ed
tsbi2sX07es/+i5vf5ZNLdNTdKEv3+QIAM/4PVWV/Lz/kPfxDmSNt8b4aICfCQfp
zhRPqMRB4GdEj349jNMKM0zHWqyCBxsi4Rc12gWsuAesNjS201hI9Kq4vt8WcOZl
XQ1r5gkZJRV6ovtKZusNJplEu2jOUzCGbNzm62jbaLWs280XohhKfpZjigJtsgU9
gWGHAWwBcyxhbY2AS0lGIkz0WXxtdd6+ODAejAorpSahr1a9Y0R175D4K8hyV34h
cHZbGHXq64/PbnNM77zZG6eT8uARXJKrGyDqKxQzFecun9Q2lt22xXyKisFXbjga
Wpe7z+SjKZ5W1PvDHHYj7icbTpFjvG6AP0jEWk/IC5JPsiPY2JG2T3M7APuZSj4L
1PnlMSse3eGLtcEKwEJ3A8pl0VhkUHmp0U/Dq/zeGrFSxkMSI6QMX1IO4IzegSdy
xXffxCOn79kZu675bQpwLeOJsveXt/PGST9mXzb8UR6x//SwD/nB6GbW2DLJMugV
s3p0OwU5n32BKN4AEtXn1q0f0JionSZ9UdZA7f3qwTAq7oamnFgH1j9stOmF9by5
6o4LL3kWgtpwquAR+3D7i6IGnByDHvHI4gFUt2VeYn1XJTsTL2wAwMhK2QKOJ9LM
w/xy3QRMaXPuI6j54w3xjLrEr1M0f6CEJpCphSag+l4nXpScUs7xXfcAZBhBP9je
IMyw7P/N/qx5oEPpUq4/NFV5YVz0hklVA3n5fNTqxPzx/qiZHbN8tXm4q2HQVMX2
pf+8nHfAD0t9//JIgp+RN4dHE65hmk5yVG17h9RnmpzDn2pXnWJ9dQUY33Sz3fqb
lta8ADBV9kkyyD2+o8SUXiwCd7qO1H21lVfNB5Nv/1cB2cFXW9TkjanEeg5VQ6Pa
DQ7DwETxrZ5Tyv2MRjBSc+rR6pvqfb/ayxso0sotNatOS3EbseePTvTIZ4CeYtfe
iTmh/reqiG9IBAx97/nOBWgwh/qOYxweAb6fvmNhMnW104g7M/z4fnPcXY27eOOL
zsSjuTeOF+JGTb+sbG34U1Tv6eMhABdMvAexA/fuHv7hwl9w6qsvvffUewgbNLye
rpKAI4ACzCdQVhPypQ8QcHy1dFLAkd0H+3Wds/ZZo79OnfSs4olz8HH2ve46yiir
DZ4R5roMmRY+ChZeuaXfVnOrGg5euXLXY74MHY7K2+gzz55gWacxfdBCSfGEg40q
9Qj2PjPYNflUe5agmD6VnFUVokjumGOKuLEa6CIdmCYsXw5RTf0EKkkOG1e4tani
lh8XQvpaJWQ9yjMw0v+tYLU3I2LugnhKrWn/WkElnFvtSzOWY6wPm0yJQ/+hyEUn
GmT4YKoXv9wedrKj5/272nj5eUS/XOdl8KmGvWX5kwfKOdj3sPKteAbxjQI9CHWA
M32A3Ukxay9H6XgmckgHoYo3Rb6+Ko5MW/s1KnzKyGkl2RvHRHOa+s6ILGNhe7Xl
2t+D54+PFXOLbunaByaDYZxxdI2szn6yr6tmNPLFqvXBMECSAdvJTSV7LC3bRDs2
2bMEzKKzMlHc5kVNq+GEQfCb1kHXz/P+dy2kHuBeV2NsX5r0ZMmXYCG5gfhX0c2Q
lKKNpYZaShYvrzQl2kfPEHnO2fMnP03gRzFZNfiDbyxHir2YZaU3YQg/kwGYSBOK
cRkaJsd2At2CUrNDFrrYvLfQy4tMOpKBfeLQrzFL+v/E1E5CYR6nA30jhUMPbtqP
Rizj3m4/sckw0LyCGPvkQl9qAhYnpy9vyLd56df4Fq5NRRqz3kd6vJCXA2Kauv8H
Lt4rJqwcZIQYspyJIn345C8HS7pVH+vAyrMH801Qv65BmgxnF2/q5edrQ0ZNL164
HKOzDtRw4bH4OMAJCnoNvT7OhzxhPUCCGXdrLvtcaQ5D3QTDvlTO+kjZ8BHOPdhZ
1wAfIHTp2a8ixfr0vfNGILQ50eg/82L+g1xEMUuQ7EHqgv+M3i7Uyy5gUcY/ZQDV
7yHHxHLS3dpBt3o97/addEV4Omkjvnql69INJBHC3rYKTUORBVOhce0Va2y6Xo2W
p0x7JlSKGW+lwx2TGH9wCXtzJ4ImSQcJahMFv7hxtS7KomDSFr6X6L5UALFA8PQl
fQj5IOoMTeNNsoDVDNeNSoNMhCVaTnWCPzEbA18w2JNLeqo++8JIRuhD+QvG9NAc
cEjhuz2gJNhCN9Fwr0z2VxMXoWfFn+0IZLnNKVM1TQhKnMNrkAiMddlGyWgUBNAt
GVwmJnUZxhWKaI4TiuENIrw8fY3gIpzfZJq9Yuq8uxx9eX8xfH2kIWCcX2FoLiPo
8cQUmMs8uI0I5idSPeagj4jwbcKJ8DO9McJOxkcS0TTu7z0e9btN+LCEjEmPnoCs
IjwWS2MK2AdGGroYhPSswvM96nNRtnV8nxOc1MQnPJN+RMiz3to7aFjhEyjnva+u
yv6hV9EPvIHu6l+z9qLRRNErgN93jsPA/ny8c/ANsSlQztkft2y+sMyj07fxoh1l
xHaXAF6mmomzuP6nrDarSTxsog3Geha8LMdjGcosu4sc1ux3yKQq7jq1vLUCJsJ2
zDw1ycKKcDPTt1qt1hceyzworsD7xd9/ycVTYBKZeXz8Ekc1kYn+ymUhcYK5vvEk
Z3ODlJG+RZILIqLGCP2E6wlzNZFob6xKuAZiCgLWZ9zuUKAr1Whfqv45c9L4A/OD
1JSGEE0d+rYRlCGsGC5aATsI/J8XmYvXiOinDBTHS4tcQ1glNIBw7uGWsUJk14n7
IDlHL7G4UlPmYuRdwtxv8Vhi7IxNCGu1PEP2fgIGNnGexDy+MwwYfKCUEJwEzzzo
/PBnHxaVKHzHDCloVfDFCpR8L3uBsqaJyyyXrMduIIeOMPQaAzLxqjetQNBdg8Gy
SdpUVmy3JEdgvW02v/QmUpkl3PeYA4ptiGQR0Pjwi8KeBltJEVXnZi/2KKDcYFZD
UdjHq2cAdlLKkgbqvOPNopyGziVEN23cTke436E3Kno9WCRIyq5oEDV8kCCay0Ma
+JHmtqXSviaAKeZ5FwL3/ujcX1ghlLb5j0lOqzrXetlcj/hBzIxRl8BnVPBQ7cs7
9gh5OsvJpVGzczHN0jOTDW58IO3diCuHFtJOSQe/Z8cwLiBCJdaTgK1qAHlWu+pl
hEgU390I65qRYbO6XFkPa3Nf+WiFal+jy1sDkASGE7zIGn+nwMy1046U3pSDJls6
uxpcNe9moObH2BK37H90UraJ6kQJCSzW7TGYz58ZaqiZ/riDgjEJXJoOoUyHFHzz
zpw86E4kQwDVMIXLNvQ63+PC9a7hbn1RBKC3yWaZas4MrlyYJUGb4XEzbcyWKAYX
y4FVHYRp9k1clDZb+wbMUNjR/bGMvuHrVgvRwpKhG1XBtNpYkU/P1quxjxmthMjF
594CVUC1PJwwjwqiKvO2tEpEdjxzD4q3jmYNpGMaJ1fB9v1ezMf0IqgUlQb0mPmI
bPKhnuT+Sm9sB0/HX/XGBtZAU5v7mwfSh5GsYS7ee4BkX08AW8sw63GxX/ih56Oj
FdhPcXvwNgtDwnUeD0iZe/2MQHvpkJfHLlmWC8UPz7fEMOo/Vr8IhoeMfLjTvlBA
EM5wBmqcXugRPK3/TYkzU+LRpUtU3JAw+pSQoFfrqKlKgvp5j7ISYgI+Vr+quVf5
IkWZaisbpZ9I2gJ/RBfkebYxeRazgYZZ5l7QPwVKQ0FtmOyoOSfJ2fr7Gv6goyyn
dp+Fy/M97gSy9/Ccy8BmDui9P1fqj0eZWEvASxkpI6o37HrLgEJdiIq4z75xnvru
olemX0wd72RhRs5tAASrbola7Zrv5CySXMcMSISuvXo2+0DlXEF9MuKd846NLxFA
cuSeDiYXLR+W4ugX4rxCOX4BeRiLXnm+hm1jFj5dFQSiVr67/oO/+KtpX/e8ScCN
uhmvRFhZ+QEqzkGk7J58a3GQNUYVLc4L9tbDy+epIXYQdfKTqHNQkqIv0tjIsHlf
nAEVCBjBpaYgRUJ3KAtFoRTwj00y3d3a/n1PyI9GbVi8R3kvVQhMIQeDHzWwY0pt
U5+dZZj66Ax2/LZgycfQV2osyKdbgnjBecDWrlD71965ucI1zF3YxwQZohwo75nF
OfX/gDGbgUAuBjd9KPURdWW5fSODDwUJL8QOOA0wMxgl611R41dCG9PNi31sbvk2
ddy10Nzn/DaPXoxZNjZ23dIVQrDn3Q9B+EoOhdi5PoNkbeZvd7pjzKfUbuuzLEuv
pW5lj2SX/kLWETWKdntLnthFZuergZo0s8R2+KffI+kZErgNQW5CbkcwI7k4IYaV
WkN8lvjkIGVXJ2st7sy+IKiG09d247ElN8Z7n9tfrPTVsUM7Nw/FZYOJY4Ae2BTX
kzPhNMMGrXzTyRPk0ViMD+gXYRg+sin99zR+qzs2h5PACM6CUk0udA8cA4qSZswK
MyCpQuYluRaJmq0PTgaGOhqlwJ4LLrdw16S4Hrt2txE/c7PI9ULE/+0NOMNOKWnT
KF1hymjrmWntlyWnjVp4UD5rEZBZ3Ol/zoNWhE1s5lwdOdWkepuW+FBShh2PkxTq
ZDP1UCCTGrq/qipkoWl9f3EAUBxLb3a61TEyTo+40eNdd/nvvODDd4xRfaRF2DCW
Hvuh/pV2vns45EeTwGPYs8CpOMbevV2POYt+00A3yWXpNyAmUW6+jXK0cqlNYNGP
cFzALb13hcudLl4sSIBPg3ytJIR41UA1Y4yYoQQ0rLQeUow6H7CRjlXqwTL/X2w7
xisOzlku96MoDEjCADoe4l8hSBhv4X9G9CXbcgbTBxOYbHliGA8JVLEjZXVrP4Z2
IwOqf4dwnxfRNA0/j5J8hGh4eQJgK2CE3b79awQI6344O8Kza4W3yK0vcjR4b4Yl
r7MCqQkHc6VMHQ8f23gT1NB5cyTJux9Jf5ic3CivBcEhSXhOvKXa8xlfm1LFrEgo
Q9KAzgz4dFe61WlxGjp0ybAwkwPUFy0TjniD73iU07FwCRvxf8jey3UauowRjyMh
TB1QrMzMz7nvBI6fr0Vmpzpn/sMHTY/XlQvWfiqODcYi0uJRdjFJ1ztVE96p0mu+
NSOZvFPbCjRkN7z/ABbQJYM+P5pF25XjjXVYhaNH26q+Zp01tiysLuLpT+x7CY+/
Fmq9iPANf+ylkOEWSki5esEs2RB3LMe4Zq5pWt8GTu6c4h7guyhnATnoH0Gs8tk5
muGS13zncn2y02vinSx9baNWOjA1IRmYQ/WeN4erSSiIrZihXSS1YHPYH266XTbn
O6BE/4US3MPVVk9+tKfA8qbbuPcdwAApqFsCKZy3rUmdRWKCJmXDCBmVnETRool2
mRsvaM5bqDWVuM2b7GeRP5RoD6CMaHSEcqh9/f3KNeO2yzG3+tCG0IJB76FwZ3Ah
RYBzTQeWzOoOqpuhXs5E7Fh1XuQf8R663pAqLhyx/72XGL7AOBKXhVqv18FSrdxF
hE3ta0/frQ19XhQN6x25NnINvLBn9y/e1+76VlkXn0SCN2cA3B9nvYcZ6sJg2lGy
HV4uPWKm6oRtXTTE8NTmg+RJXYDrlqBEbTsK+8+kZuL4+rPsRG0MIlRL27/rrBt5
FWYc8gmnGN/KWXhILaLdlmgIFrByjiSU6c6pxlRBOj7smK0T8YJFe+eqQslbhuQx
UFi6J+3A8/lb37LxLV50UMqhDVBmswUm0KbtWBY7N4OoNpWqJ1xqZBn0zij+q8K6
bpkT9Uu6Fzouk4SIiT7q19uKePbZHduFU58dAoK9GhaQX8fi2gWWUmelNoAjdcYT
4SiWSGHlR6fmekUDIVmZ7EfaITtplXz2reLKQDAwaS2ImUNoutq9ZYjLMUrSZavi
TSOZlpylXNv3KsW4nepWBWVDEQEus3JUzXwBWIqZfYhsLsDJ8QbBhosm/TfZfUzA
YqEO+KHbXXjIRR83eTc+MskTNWYZFrdezLJAzR0cafLUvaSeWc3Tia23f97tiG+W
MCKYFh8wXFMyxu+nXZ6iooQNE2RCryVfi/2V8JefzKPb4VKKdYp8RWP9nkJzGofW
JuiKQXJ71XH6IfSzX/FEktg7OhhyFGb1dzSPZ0v8EAD773afGocTAm/uyzizjedo
AUgnxHA7tkYglgODVWoLlvdSY/SkKubJyAVvyJPlq2MBBQvrTM8b6+5MWht/5H2K
zVLDo+iO3wWH0NM4lmXF0DxfRqpS0MNU1yzkIT5GjxthU7eEpKv4mSubuh6AEH9e
om1rNHB0ggzvo2vXhEzauobJXSWFGMqe3BS9ugXKCrM1pM2rPbbgrX4kGUoE8M6b
eopWK9nYIPynREiqzASfuaU3cQGSaH4TvqcJgRFIyFKVKRVCJc503P3zWFGHT6nX
xxCybUR5CGtwjgDDZXh+P3dp1YdhPB0VBlsMK/nzIyXWjBbvPLztzjgg049BzfLf
bbsxtGn4Fndzojr5O7Zb9uf0p3FdBRqFIbXbZMXgm+qsymVfbGLXv++4notKmlxV
0YhTu3/t1P2HOW1iXOUDDUwapcGkJYB5LNmEn0jJ/5CDekBgPvcEv16q/IvHsdv4
EbSDs3x4xXaLsEMn4f15IuoO+lVHP1BXYulFusk6P1K/DoqsLJkxHcQBRZiOA+H7
curwcMJ7yT1UV4tbMjUqWBS2LiSwAnkBHTxzlQMJLh3NCCJhZPC3Q0edEFaaKKbd
ORyfaSQ2I+dAV2Gm5USplU16Vlh9FoSEUoUBdeet0v+NbKC6nQjPIypc9n8biN3X
8Twz4g22reQro6NULm5JUfHj5gXEij/qtMZGuMXninuHHLTcCKZIZlutwWPv02J2
jVBvy0mB/BSsSPFUBPhdmdEBes2Q5C+OJICJylzLJS3/efGvop9C0EMULhyXM73F
MJ/szDnCLrJ6IygMFbSqgND4vTFgwL1TqRRGBr+CJTDvgZaTnqRk4dxnh4qAfwH2
+njMZ9JCm3XkodmYNb3usF0VCnApKYCfaJighKPfvyDlgak9TN1kT8cDCd1qmowM
Jn+NG/rfNQMBtHVL5+2+Jwt37Dz6QtBfFyEOs4MJCTRCPJTCJ0HurLNLTjvtMaWJ
xIdo3/3uFbyr2l2eFDas1D939jD7VyLGJsPDyUrVxqkYxLBlZVDs1E/cuPaKmcOf
Gt5GIwgwQQEBXy3ZONGe5GUNY74DgDFMghV5kbn92Z0jXmxp6C8pcfBLxLN4SK1d
NyyYoUolmkNRZIunteMb88GBXr0ntScPnk9zHXIWQDlYn16FwgXA6ZI6XtBwUrv7
Ps/Umx1kzgupk3z1EWXmfuI2+Z/JcwMEvbh/RGJkgdNsroYnUP49UgGcWKZ2oDYV
zqBAGJg+oyamdtVbOA2ujJl19JuNLmsK0NpASXgr+WL6j/p/cwWAFBe5askr9YV3
DDYDk5OPLmt5si9vxytfgEtg7RDpJJHL7QqryK0GYFKCHhqp/uR4zoFNzsedOMIA
IStz4bBrPucKVwwGFf671awfnzHiSiTLyKsGRQf44sav4TxdU5kxUiJxD+mFdqbD
lguG0XPdjbos1WtTSozhSpNnXZnI2zQWugsNouOo+y8hTREk+0aahWJ/8FvTntSY
4dj3p8Mvjx99P3aLetqrnE6wIuQLzuf9Hkwh94hNrH9S9ik22qB198Tbg7EtMHM5
MS3CtxX4a9JrT2AugHqXJ2qLGkiwjxyXkfDeGrWWZebWCns0nTyCycE3TmyQedXq
1Fkq0M6h1bZiuBScfoZ85dNQj9n6U2u0YaPRH76Dl9pHm7Wph0Bx2/PtSrUUidUy
KgLz67ZHzm0pMyj/5el8o2vLOtrhJH0Z5bIInk5Wm6BrVAO1XLfRO5212idssar+
09yt8EtCmkfkUcQ4i8G7p7AH8ZZKr3vtWO2GKlttdeAidDw5w3Rp/wsv4CiXBoVi
VZiIaiHUQIus5nWMy9IvaVUPUKfMKue/DgRMSC07HAqdFy4pHIWFVL7oRe/YRl9Q
jlvbi0Z18pCGOn9mHZXrrRBEawT3QHikGryWg9acj8VHEZjwoJ6BzUaF1ojBHaKM
D0cUqN47kdWL2CNEjkrOLDv7Rq2NCg54S4zZnU+62b/yqNGnZiA7W7+pbjURVXcb
kHKkHE7SgSsii+ybjJwb9sKI4pu7QYPaSTRgcoAyt6Em6o9pshIhhwqlRenwED3U
GEht2BZSTwGvZoxRxGXyhqTtNQVTCdy3eKd+ZIFo5QkldvhjTAYouiM3ehSVdUID
HSjoQBjvEYHnIG3ZzLsw6F+qMeWGFBpp1qiOq9jv8Cd9bEJ33N35J+oyPxZOyWE5
VYfzVBvgjNWSRJKXFFrUN4sWXVVNZo65NbZEF2y3858E3E9Iv6h56RYC3XdHhxoZ
i/DECReM7rdpmfh4IDzvyUS37kww/8MQ1czRryJ/8qAyZGP1zoYGBf+snxkR8QV0
towHWKQYOMTCH1z+AtzopAd9hzKVCUhDjguC7J3moSRoRG0UzMvY2rU5iFj/NesB
S2jfge5MxwT4y5zy1k+BwxzrjoJZjkf+YNSlX+KDlVU3ZLKiCVuZuGT6GkKBl4tj
jHBzsUKL74a2DDtZJs5XmakKgsSsFdkBsd1pPdQAB/sKyC59YzbqUrqyXizgEIyf
Rt6M9x3eCKPdntLtdWpxtxmf1puGvmlib0104/amZ0l6jj/XGTRSg3Pr1k9JF1HA
izz9YVzlu/H73gkjgwxGtrXgqHlo1SzZ/0tp6HFF59P4Y1IfDbcjZvqru6LBj3+E
68s/GOtHydlZAeZoEaibn210zC7PON8aYSSLDM7xGA5EhYoa8usr7RuUKqIniw3A
Gnldl7vhiFB5mXPpiCqZjGLPZfNtAbKUPruEJm4TZC/62RPLcuQTsbNN0YIbRjAo
j9UsrVsHwsmO8LkSp8aaiLTqMMExfgqO2YSPRsEXpkike4KG0v7sjcC4FgWkMk37
yd7N17ACQLMu+9wBmwAMi3ZhL7e2W30nlsDuMMzUCUJnW/Ipt0+mTfkbjxi2d3GI
f0qDrloUJotFafkB5RYxuUkJF6RE0QMpEcZ+k/AkJwJHPfoPeybAK2HgzK0e1skv
WlqIOpwpWGE+I7RpZeh46TGTCmNmdKynFnobKiLOZJnPlhLTvDauwmQCHEIBlaVg
b9CvXvZ6C0dMUmW14KacUwLVOtYgrczV+DgCuGQEDRNIyUIIavOsEz3Zqalft1UZ
N8Ql0vYddoovcEevD6mq5z2j0yBp6PF9OCA1fdtuoTSXqGA7iPEefgBGrDWJ+jTj
ZF7HUVXKYhNVJU1RCS95nLvR1wNmJdy032FZpBGYCvdmR3nEuz/GUv/5VmVwDsPW
p29xrPvGb12GGFOHGTzMWse3ht9x3xEE7v4cp9tMnzTx0Y3pOLYxRfPlsrh+LWPw
uQWIo0bsu9Ranc07Mzr7wDOPHSa6thhdvRDgi9mjRa8/mwFSOIT8OmVm8VRKXCNG
sL1eoXV8XNXG/ZIdf0F+QxzyIimXc8ZG9kJRxR8Mp88X8zIZL8cOBLLR0J4zlIVK
5ZWiRAE30fVWbywzYl4HilxN0gUl7fwzWuhrhILJFT+QrZHIookVXyzmXkaQcr6j
N4/vsgx4qs0VCbOMVsQEJdNhKKEbZ5jZvP+S5GDmtXNrB78G8ZOluqUUhVZAZ7rR
M5CJK6qCtL54bqoraoyv9tUNqhniV+OEClBRB7/FLASaEh0AeLfMMeTfpl5izXF3
8+ArqzY7xg+bJ1eC5ahJdmGI6F/NJ+7dKjsb7FUpSv/4P1ziP9GwFgJuUfCLD02E
pDgAsqxaHE6bNpOxSd/xQTs5po60d4vYlE9dCV/Ej6qWscuHoqt1StTL/eWje87W
PKNLPxdzKixuXyXdXO3mHZNHJhUngG8gzOAhBQKswm87IeLVjLZwmPGx94/AjKUH
n2nbZ9oUQdZZOfi0JXIbRGSN2ili6+kf2zmM8ejTBzl9/aZupeb51Cw6rWyqhMco
4iweBdnO4/lj5HjxWFNABnv2LAkyh9VpIjnguxQDa1yweEuHf6PfoRC/25+iyu8+
RgUbIQ1/2SWxCxznHkS023OGPD5tc+JULQ9M3UEo/4c3vnCgnm2NZhwID8wXFNQz
s1Y5BH15VcKXkzcFDgYKozb61jpW6QNTLY21+TVFt7pM0W+8cbjiBc0dVVcP9R0P
oVXnApAauMqbKaZ62iaafHvmR6P5n7Y9GIzybmLVJrbvcY5pk6O3bMLpJVNQMcRG
sEyNbf0KyJN+Jri6DDHPPHnOV6UjQE1EgGNm01YVDRMmCLdXoIN5leEToF5zgN/p
vs+S+Qo1TM4osAzNdYWOFbnoApDIqLmt1bm4105owWo/hHvpDH/LeB7TAa2ojAb3
A17J8ZhiYrJ1GDXMJaoFg1N/xUQMmpR7tpaMy1D/1y6i9diuG6c/QuZRfkH0Wequ
ydbjXNMhemt+8nLApKU4tr+SypAqTyIilbn7k3SuSsZYHJHJB23vORr1ljPLQykw
icK7bzMj30fnD2rmCvHgoH2Jdtv0zVoImVmigdj7kfxWPrb9NgWmuIO/mtpDnwcb
OQYb+J0qKtDB6jE/UrhIp8QDraIvKpWWEeg8T/X5aBcrXUxh8fjpqj6SK0QZaOf3
b+2jZZDTFoDzH2kDqQRKMboHSjWC67/mQnJjgxXMXLchvDPp5tx8swcqmGBbz0Yd
zYo1CGs2+E2rxBiur5ixTTOYUbgxGBLcpVISplbModBEeXLAkEUCg47bekbM0rxF
9JxGb/10AI0qiaU/5zIwqgSpJx+sft7xlB+IGSoqL81+EHMJwfaAFH9xHnTmGFoT
lhrIaXeLK+/hmNZMQKpL7wX8jn0OdFV6tN4Bjja+3zbXa4QDtKlNPriEv0cJ2Dp8
JfOz1nhhBuQURFVDHF2GyrO4wT/86FbP56USlpJ+fdtT6FpoO3fVdiTWKbhOu3Xl
aRF0sLVN9+YJQuVqdD5dA3MezfgHnERTHcHR6u13DjgtEDbvRtaPk/SZLSZYnwgT
NhkrML6+azXkoQLFkmkkQwiE67OqadCvYLbvNvK89RGR4fX+ypeuANtYjejCg8ct
YauAVXJ/91uz/oUoNvpZljDtWacLj+WzqnEI0KVk44GJfISdqP4Zv8+4ss8QDHyj
T3hfssfefOYH+HLkQ2P22pvcd3FgLfGnKrmBVKQb/Wh5VIFeYpLFDpS6fYx58SRE
vlL+mL/rXqbnUGCTjTrg2HnKXWr8Zq2HZXoFyDnKSj+tbdbjGNfbN3rx7o8SNTLw
Al0t/f6l3X/ntunKCgrJ+9weFJpAF2PwMrPF0ngX1DuYnCmpm0UGrEXbgZZjWFAf
sV+dbOviiuTEecOlZvXCZdRbI7BAzPFC40VK2WsjstwE/YAfJNU6NCh7WzX8nbLO
3VB1ZiAjuzW0Vxh21wGs9acKxFSyM0objwLRln8ICMcAEaE7kAP06aW/lZejJDXr
h0Edvjh7vYE7vfzxaS7e4KzsjtivmY0D+3kaNxpRDQsVn1Sfou09F/9BUyMsGnyj
WlFCvSk6+P0LrJEKEKZgoXnp47MTdwMpdSsDiGXY3OLHc3+tqgoKISeDBufl1sxZ
Kef/eE9chNpDCtWnb6bSyJq/gJdcbeQOfIguhHhYPuVX5FFgEmodBMMyzTpYlRl8
KY/CzAV6PqWpMSYj/+2DKrcyC7ogHN4V40a6/7OtGEkkb5CEYSdhQHetYA1lH8D5
Hfv+qFGoTDitYAYrvv3M/bLP9di6tCEU34I1uTW3zt/Z3BLqrEDcBnp/vPLW9g8w
uwCoZxXDhhbineHVCl7Wrke7buyj/JYqdOAgeYAoxcDOQGLR2cIW12/nxVJhx691
Al/DT0bzR4Rtw+98rXFTXvEi1fA38nWuw9/6v55IFjBaSM8tJIZJgOkivGgcFi86
yFZCj4EBw2Vfy4//XV5ywCZSftHXVNCta3v5LDeNVjUIXonrUQp++ttC83i3zFh3
89vFPNYw4kpc31lObhJbA/VJ5dBH5LOOJ3V3BKCRIDnrCpoPwJbBz8dQ3ZtQWrjN
UdSanLFU55lXFEbddqfnmv4pR+wAO2PpILFc7AFx97JqoI4BtVgSxmZ3GOrT7l+D
V4wZx23ueJkIvh3SLII9oyowl7u/+ssJ+wvLHRcc1EiUeIxBmZAv5u+NeR+eLXox
57EtVEKGyGMB4kaxZ550/WfQNWBnt7Gu6D/x7e4a6YZtspp+pJFhVU/BuenmawrW
vs6U0G/WjyYJc34BF2yKO+k9J2SwHpcazch5NdH/CdNdSECfsFeFPCyPJoBftvJS
4CK0qu5cQLi7dcFl6+NFUCEaNMx4vasU/8wCah3uGFwwu2kouEP3nNQjZxAQCb8L
cr2BnaQ+IWP35Xgk3ZoOUv+oFW5P/71O0R79USxQMQ6oTjSqMQkopRHGdO6GqaSM
AYNO8GCVV2UYG2OozRjwH7AmEUUFwGKkK/bLiWY86A1IzrJlLGgisgn5Ix+HY3nV
HBja0Xf0hsh0lMJoF/ZHKK8JrSS/Z38X+WZzsDMWXN/CkaXeOvPRpMvFld6DM7Ye
LyzzfdxoLq5F/82JqnMLD14NlgKW9D+ABZ4Tsgbh6oI85vFggu7BdFiFM0B4WEE3
tdw7B9VyyXHC4LY1wuI2Z43hITB8vBXTgP1ItGQbVQN9qBWX9Fq88sX5YgluFny+
mlY5EYj+fYB3+sFvQa4t7gSpRMxdAsABktglBwAJoG0v+wW8oPRc9kxrSoU3hPap
lvkDRZOUh3FLWbq8t0cRxT7mrOMLWpJOH8jM3aoJvXitJb9WeF/RDRvfy6aovz/S
lFlL1bUYM/T0McICou0b8MwuzGjIesRtb3AdnsRYKcZtqX8xHVgUKb/3a7wKXukH
F8002pYABlXisRtZPJgvddX2jgU7oMaixXqxsA7VR4zJCHnKXv5Mr9v11MlVEepb
dxESAf5VHYykN81n4b74xDpMaJPfIlPScZqwX/WhPtnG4UJL1Lc/G835cMnMf+8X
OJw/LaLxJN5f6LB4SsPx+3XpM7pHBDYRKni+tyH2ikcg+Mw8RSixbHDNgyB2z7Nz
HNRnygQePlg+Glh18OZ/hof9U/tA+vKNOEHPwAaoL4uTVBaTI8UqxpZVP0LqonF6
87W6+2RWCBGh1ExPYQmTh5IE+rjA282M2M0tcGzj2HmhecUeeoBvB6yJfN8h+cBK
a2t3xpsvcPE/7hQoBrwE8vENb/bbjiBmP7TZUv9ltrP1mUmjTqOptXfY2O8kCUub
JDQuyoyqUJQpmQt7vk4PC6PHb7ScxYG4RiZAlkz/ohuh5KE7ysGgMmP0hfn2xDi8
u/XtvN+g5NKMhmjaMWTx8M9NqICinG/5jh3IH3Uf46qX35DoV55/GI0BmB/6rRMc
dpP0setWD2GWQF7mc7IX3paqEHOjU2IHkslQ47+Ix1UBZ3k63otmRWzdBkaHOyyG
kRKP2+TOcc1i+Qnfj/RvLAVcu1d9ya/nZEeJG7yMFJuBvHRpeZLpP1FE7mR4HLFT
NpmOeD6iSudg/y1X9o8meOvXLftTLCLuBzF17VZ7dOsJ0BPN4ub91ijyVGyuQnml
ZCveM3JfhDsi4qAnOoJbsifqeGUy6X7xPFkJznH60WO2SkirhJa/bCMLA+WH71kj
yA5e+zJvOx1eBZSntd7qUo3iBQzX2Vln1nc4Z60yhJVYu74XSKEMDgnyFQU+mgS1
bLJhcDv+ZJZ8xBq65p+H1vDQw8wXyLgqW9LS/FEbj9iBtH/G75dTuWB0lA6z4+3W
Scp5+apSdIe5GwDGAqpuaqSRdt8fm1zX1uqtd+Ph12dE273i9eahfCKgwpGvTp+S
rZk5rZ5WHpAXwS7kz+jHZVfFYT+PDBklpgwvzl542kgkIeDxqjFlTgp7rDEhQunG
7S4+uFoqBQrgXQ3//2KVLoputtd/DQcFmgapZ7P1te9qE/t3VjvfjKqxjGZ8wgm0
AeYV5+ttdF1aJcGxn49sNfX6uhocGBCqoDMlGJdtvaDTNtUkVED+nWzglVcudU8S
MLTGfhR3IlNTR5yT/KbcFK1bqx4SVGvWMTOp/XJYsWtzFHk92xKPYn8JruL6GFjN
0iHVQTYu5Xw7isJ4+QsB2ldI7fYaIcIan2GRgfEXMNJwCUOhjyHfGXBHTlMlRi3p
JF+PDIcAtI7uMla1tt7mF878Ej/eG3GY39y4ORU8j3oxDt4dSe7SpdjkBvJZG/A9
0+RzzcRYSKEen7P7s0mM6HAzMLpakraANakS7PhY8rJBNkveRrnLbOw/BC1espwC
76ORJjrjt2U8dqnHz8Z+LrKK3AVdIvFzAagQ7Y9Y2MUFIg2QFSK7L5v8r7xQYxgq
aImyZkhpP8T2YWsX0xiq6V9qDr6lhBarCu6MUnVyfxhatp+SWcMRlXUFgJ2d1DLb
6TG4TihnGzFlRFFCoauSohu4p+rfiHkzRr558F+cR6XsvSWxTI+DQICNCZnF+/iG
BDrx94El8P4dI/Eb2dNZHVBe8lb8D6/L0gpzAEMyc9XJgyWRsTZdnp3AZCeDM3EZ
SI18OsWBbaJDWU3nj6wZUkB4y9ENR3vVoLyNnelZ6YIibOVDoImpTE4LtzbYFWrN
LZM3HYyJisg5cxqWUOWzPXcYO5KxMufUwWOgi2N248cLjC4J2jsJpeVXOIP3+/Zd
coSd//2Ac78P948R7Yy8HEbuIHZtdDXJUDlfmuq4DBBv7f+t/s9WIbKfr7UXvXTM
i931As86ogP3Fdbo+mF5Mukf97Qu7I0hcGpry+ZNFXgcfKcN/PSlxuycBeDi28ML
fJ/HF3+rYpMQQOI3iJ3D64SamEPKp0if+QVR7YlfHBeqsW8MDM2FvO2FpK/fL5UA
LxQFRAow1W3NF7+mDarwCYCCzIEFthOJwxSb8kDmY6FJXUVJmqoALVRiTdvUJpJf
NEVr1TRAPPuFkhT5ie5p8Jf7WYca/J7wsnBdFhtEK0TXSCPS0dRpq6jbwApD0+DZ
UK2AcTeZDB3Uukmir0EouZUyuN6oSY4CMYcgnlJEknGWO4TGTzdLixCGR5O2y5+0
gOPGYmJW02+gmd5ntKEppgHImqDuzQKazw+pOyZGIOKohHocBlULp+o2DdHaEvnk
fHShecWVrDXJVWwKb/0ZYM8qDAFFVWRKTLJKNGO6xpPSGhjnAhoBvId1uAiXsVbs
pq4PdiokodqlTgHHTrO1wjyTUC2mEdorAALwubuPHZj8RzrnU9uYoBh/mf5ilOBG
IlRHG7uA1wdNaibzzkW6d+26fyMCeo0ajfNWor+tHAHHF6gbg1ecBMg7dLRpiKNB
XLVRgSZAYm8I0mB80xrhz48ofSMz7A3iG0tlgN2/AX1hah33W9zUxxnUfwkymVlP
P20u3TXKkj1mDbp03N7mQhCaTOiZZBtIDtcw07RUYiHhsbTtEon16faYbOSj8Cx8
3vADLJbODcnciSpJwTINYX1b8ODkD6L7NpYK/nbYsUIJtz4Qda3KUzrdqWNrZpbQ
K1T8ljngorJoG4s8Od8M+RikmL8dmgdhOkkFXNFXSAP1VchjgeXX8WBI3Va34fxq
riwCcteam22rUezTHSAM+8uWH4OVkDVPFHgKnkLseSnpQ6OW6pqAuIQeiVlMfhqF
KjhsBKfhIlwC8bEoja1keGtT0Q69OBK7O8pUYEwHTL7xLO7mD+ZEIvE+OGAQ6YfO
71E05X2Nn4fRjUYapFAqt/VoN+8+Xoq9yzrTHoN61aYSqfL5jl4uxcF1mHpBlrcz
74HNxz1dfuu96JGjcPqYn6YgXRw6d4jzwMwi9wrHJmjjM0OrFgfLJRB/qhqELHih
UTB+oJnOOW1ckhbi1PdLwBWxWg55EYzs4xZFPq6mIDNpByxE+rLeOUhbPCccnIDE
4G1n8W+kbQFOBZnr69KnO2wzWs1Rl641nMEugksZPy10fFi2fy4koGR3sAIfR8JN
12zHCWFOAEJfkHqvgWUsV4b82uEJCye2cIN/4siLiTfZz59PrMqHTvLTpO1koBAX
sx+C9GbvZ/mdz2X0+qaQuBgDLUwwjz2WbZU25em5dh8CxgDZYP+ArYoEtE/wJX3+
jWHaB+wit0D13uL5wtmRJ9Q4yqr0iRRlmhGcJeWB3Z/A2HGKKS6unkpNddLqd2Ao
8XD0CYKQ4ktU8lSFec7lsxAUCInxPaZRQ1O7iC/rnNnGZk3URou9xClyvXVHCqw4
bwxyU84Ccr5UEI+/b8aCS9X1L0s0CfWAKR1rAqGmGynUDmvoFd+OUiKUkbC7uy3p
601kHq4K3RG9d293WCKdOOzZtEZClVgFQNTr2nbqFvxAI7en3sYAwUbE9b+40BXN
N91X/bIDkB/icSQRsztpOfxUD5dpFlwx8kSqgSidBRqm+VATQnKTyrtFXZ+i2y+6
0jVXV/R48LuuIiB/1nf1Ld/AHzfCTWBedmsLQrmjzkay1wli2CmCHaLM7SjlW0Iq
VhiKOY16x97L7vrbpK+CowZ3WHo6HKhDVaQDM1T4GSazbG/SJD/oBj7T5z+Bgy8k
8EahmVy2pevVx2ZAxu7nIny9k4hcbSSrt5/i3cQOwBZAz+isS5/GuOGfLmF55e7n
b/BHVP72nhZVUna8X6r6lPS55G9A4YSnZ7Z1oGMOTYlhWbeQ5gjlFdf29h2mksaF
oHtFmlCDIi7sWQlAvQaLtwIiHO73I+jagpGQGQAdrjpHXxfxiFvUMGdjVTvnaPVb
lVuwFKjC6fgSDC/oAfXBYOrB37x+H+7PNJ/PZTdkVS/6njO/Lh4gZ/T91xl9FrOe
X7wHS4BVWGwu03XY4dhVBHtldM3BxpcRYFNxYR23EHU7CvbC3Xwq8GvRt4gsvfoE
zyRnos8Ofv8Y4gYRaCah47oi1brMvIlgCR48HWlsMv04VtcbEKXvruWyYNtWEYj5
`protect end_protected