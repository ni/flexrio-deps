`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
N+AbGUvfDpEoMIf7wLov5TLS6K232jp129EYKy0xiRWgVZvvzMhtpiIthRJpbZcl
F263Bp6GauBYx5qAJg8nn4jmzWxSQf4qplGHmrbXjafdUlw4d3V0E8aw1c2ZUMXD
8HNVOolMEcgwWnxMc007SFGcJhn9F6nyEbprOe9d+imNQQh1oLQeO8xXmOy9uHlV
1gGzEmkYiv2GZLIiEdNPkjsZGXyc10d34Y4B7bVclxzUjKKCBhs325vpZH73Jk2D
nRmF3Q2pooGsWT778cD4Ip16foQYa9CEKCy/F4csjdbR8Kc1YeWYHXV86eCBwHq8
Lu4AEWTT3OQAlGzmf4H9hcBttpe2lt8sfAY6tT9qKt/0lbhtEsHI/Mco3Btir8ri
pg385Pd/sLE6wfzO/XfY+rt64Z58bQMWyIZkVvMJvXNg6azjsJuU6enCLK0sYVyq
JgmD+/dXFjzmhaurRRacXQfEdW00Cfj90ziGrjHHGE/V9Hg9o9741f8oMwzKH2Es
+8WyhzD+CCTeRd2DdIZ2nd3MMjOpXtWM4zEI3Wm0Rmegrxq5flp0LPkkYKUVXE+c
JJUVx6dw0DzBAdpNZQH18XwpKNzc6uBhEY/cqo9Nrk4CkRX7dqK+zgJRWLnZ9sz+
e7ywSKLdIEe5FXvoMn26TLClapBYYXS4U7OJb0A6FIYiuDZoi4Izdlw1gCNYuiAe
PV6Ov0bw65yqaMi3q62d8kePKR7hRDLA4XhVQgm0SLezS40J052kUk1Uzl3zdD+g
8CgBgLeNqVOPta6mSYzFnXpv9YYMThPXPNALCakBQK0Mc/HITTS/9SsvplUwpTDX
/O5xv918rJTsO9rusm6zd1tA8kvJe7eHDXgQZe+AmA1uVxkQ/R1IGj8gbmhRwhnv
qzTEwIXBbvgGTYlZ8xhOSmskEONBNyjbVxNCt1Sy5kEc4XnxaiMSPsnboNTi5xW5
EDMbWac47oRbbEn+jbjXH4r06g8oKUu7+AUXv8MySohcoRzvYW5PxHaqunQCMxFH
HC0qxa0ec5rLN7Klx2dgCRWO/tJ7NAyi8/ns8XD2yOjhYAZQq6u7zmjNlC+djBtj
dzwS2hcmTbmAnDU39i/o9wI6FhPJ06LHo6WMLsKjt6YTULEweXaUIna6PHy2sOL+
fnJlW5Deauc0YynPm3cDgwH7vWOfNQQxP4P4lQT8yoh9vUi77om3F9kLSJ1Y2NOO
N0M6UjMobjUG0YhBd0K8HpBXRRjJPWPq3ODkxqS784vPMJruBVKDacpEIfElZnbi
UQK6vp37aYrDH7xkoD/jw+ycAAYNI4SQVcjG64LurcHbpsV+vQT0Sp0TFUiKYhVT
PmQp70eOeTLXTK/q5dHgGlt3CBtkzKoGrexzvY8WsBzlllYU9rpcKkeKPGkHuXC5
Gx7uCiiWa8WVwLrfC2JCFN6RpscECp1fbFWbyw+Ct111atdz23FkI1llQcMI31NI
nExfErwWMyvKAJwGvEIZ8juigHfKrfmIebtZxQJRqsYS+LmB3DT5ioSurnJTMvI1
nCzX5TDWAbJ9fJfyQewkYiZOsAnuooesY3lgTmP/uhLGLGPEdczhHXV++IUutB4L
bh50oYWStoJWGWC8gcxzOAQszUo7F2ETi60JBIosWtTEwKEb3qPZLE8C5Z6OkWGr
8Uy7A3Kf9eDds/+7OpyXmQomY9DOpRbhDbiXnKpedb3ot36Hb/QY6LUyCsqZk5Zx
+ek8EfoK75HGcHi634pgNIN6HooyoAtx0yEkUMbj79AfhQwPRbNPCYxJO2EUxFg3
pxpcQgfvDaq8V8innf3RCMLNsuHUn2DbbelL+lvCjvvZrxtXv9yN+/9/fOyFbOg1
VdnOZ5aHmgkOdket0+ARLU3crJtGj/VOrWNTjCpKnToMgSkFvik3k5ZXFi2mTM8g
iQI7EUkNgR/r/Ue/ItGOsVGAPHuGVgfdj/BdiztyT5NX2oSxx962uZQB3HQf6IGx
j9kOXS0ac8S43iXGMx8CklLYi9dLIpJ5Xl1DAmwrSVE0LCRA4taR05R/rfMws7zl
Aib5yukaLu2Ba2rWa/eEm4MYAeSjYm+YTb1VrkXj4Kx42OmNLEOcxFc/HKwzT0oX
Y8BSgTLMec176z+KvumuIoEX4y4zTZOIjJ7PUcFXL04CXeX6kKiSbjMWtcfI5rBp
o5x1BWb4kXkHr+qxoS3tlFN4NrgkpgUBKcMkEnvRhMMNucQVr0OSiVj069LHqYsT
1/YJG34KYdOT2W0CyfjhMUhdK8OaxkcPJajuCmyqBkPpHeW7Vh6ShmI9BNG5hJ97
2nPP8nzAddXE05OrQ83WnfK0vBV7p4/GReUfdJ33gTbld7aOeP9gIzNF0dUkp4pZ
ppF75pvbVaL+/UnWSI0e1oOdwJQLktC5XE5JVK38Bxp8CDpvMdtqpmuOyI3KYt2H
ypZzlnxncu26GspsvCSYmdJI5HKLCbM6ZO29dpmdAzhXhKCphi3HLrkF2kcbPIU7
x7IlG9xzDCfQQH7GpiSMbd/c2SkTPAuL5mbfarKPrHwyiRKUvMeERUnitDrzepIv
vPYIJdP2AAiusXnL4eOljQuB1T4jgNuLK9otTUhu05Titc3s6oy6XpSTfP7yxsXK
pz400/u6ZZWvPNso5sHdkXcuxfDkBDo82RKHDcLS7oPyHPdw1fqwwzcIgdeufIGl
OGGqDodKs614KjjnyoK0gUvEfIsTX8jeMa1NgAbdPjlDAX493xk7QcnOsmQBZfaj
OzT+GFEJZSjEDtwgIsnFHukGHph4loCooKPeKA5ibnGYApNuoQcVAJZyiy416QIT
v/tyE9st61vFVVtCPzxm22mxY6ZvEAWhAHL2AWbrOz4FItPwlKluzkJXezYJEyKP
Pe1PEC2One+ZzuNZrIL3sIYtUJOOirRrP6ZWQiNwcCkQMDlVMigL8VOPRw8/2ONW
7Hugp43wseukqiRnsFhxjnqZc/lKog4CFSW5zorMiRskZkDIcvx/IYLnpR/vrwI6
bd51hCK4azxkNob/d+j/t0P5sdPq5TtbQjt2QFsL/atvDUR7KiKnDDZb8G1MIrCd
OD4sAeB8lVAzhiAsPQGqzr3lEeqBfp3lQH8EmFB+FuNCzApqc/QlH+sT6qQ/3GAi
iNCiR+E0HuOzU1QvGG9+iID9G8PMImh2mHxWaRWl6UoRX9wV50Ifs6CX7Tfz5Yzc
v6xjcxvIYsLm3ys/nPu/5tUwIMI1NaVJ55xOP5fLysfN2ubP0c6+PjENbV1wbzeg
DEeGmfbdXQ/EG/Lgbw9JvLZko1KGU22Qe3SCIazwzTS2TYXaqSe5USFPK12SiHwS
1MscqKl/iGzQ6hhhHeiGkNWbaQvS7hYhmbQ0EKCgGB3Dvzv8bM6zLgBcgCv79/Oo
1UY5xct6QYM4/s6A1Nm599HWZhvGjbF24o151H10nx/KpYgQq5wEgWWc0u0hNCTf
bi3ZKEqifSPpYxw5XzMJwpUztAVO+k1gudh9We64KM15OChEWTAW2dLXzOX3FCuE
I/pxL3ORJeIC1q6Lr3wl1k0Jhon98yUC0aLOD74KiCbjQPt4XZMZxaIaEK7fnnrf
aT2c6sE3+88a6SSTsZEasxr9oQFKQG3t4csjkJPhwrc26aCR099piKv1nFRPWdJ5
W9UM0FW3QiwOuMGC+0L8Ik9NWR0ygnTEbIpwXrwazDf7Um3Nx6r0c7yVZG6ByhSm
kSyLpRi2sTCDtWkrBUm7r/BEZWoQwUvwohC7yz/N2uyq21rgybR4D3QnFqLZao9N
GHOFfwp5HuGNtxfZLnww6VNbH7xlTwjS/jnoiF4OIDfUCwu/4Kn2IojhkxPe4ziT
I6TiyfyA0eH8pG6Ub8aCXimtJkt5Hy1HnYM7+bSXUmgIox/x5AMwWOipsM7Ginif
mQT2eqsWCzoFUr9Np/ZTjqQvApCKjLA2y0G28Libo31IrXveeTwlLaBv21x8eTrF
KZPtxMNJQh3MF5nehlOlSoOR55GVkwMsGwz2j7kfMr6KFGx8f7a3DOYlM333282D
jW0Pwzqot1fDA8889UbZ93vuQz+r+S7SjmQ6RwDATbkTkRR7D868/eDDCpWoHUC3
B+rjVUJ5ED2kU6CxCBikMsmAchcNgCdOJ/vJuvNzP0pr169/9rB0BC2pbz0HNWHp
7sMj57rS7wyl/eNNjRGt6LOV0o4wOVpZf2f6SVgiz1IfiTdV2k1kuC8UGR6jWvYX
ne2gXwn+atG3AEKY5iUbW1lSLPlJzBfqk9m2EReviG57cagLBWt4OiLwGCdnGUOW
dLT5i1bfnFUfbdF8fl3q7U4Rf5GOQ2ZGfS8jYRThfbeErsDmgOnch5GDgceRV4pi
LhyESoYDH43WsrGaiGub5F9/bdX+jNSXvhzV0IqOYJWmhVm1KW4jLfeN81oWKvAM
LD+jIEDOPdd2udj76XIWYaY8CGTEAT0ZrZAOvkmbGkcc8Kd500RMg93iK+tmlcIN
l2isl0kj1YQ2TQEhLhgUoNsVH6hHPQ03RfI3kdJuwWs+7r5rEZul0K1wjZcA8cIH
ZrxA1Xox0hIjTWwpVvTgUdUiDvUamDQ57Ke0qq6Rq94V4Rdzcsp7DPNuwjSWq3hS
KmYLIroTwXOF0pY+CvkKJcxac/uNVopMJQnyKujvcg+BPbxJ3NPhA3PNPr2haH53
djBCbybRm/QKuvtbKLKZ+rjtkjuc8vVfp4UsnF+t7B2B2pXd55kFCd+rXp2rhhag
sRaTSUhRJ29PGHhidyyIGlu7SRumeOTS3zXydOfePXoznYZNnG1SYXXx0Bs0K9Eo
O0Sufj8Cpnl4GN3oR9u0CIXe2jLsSlUvsBLg+/xPNXPj3uuA4JPIZYYxoRWAho0x
+piemxlZgtZvpK2Z2YD2iCD5YryUGMNcFu/NMm1KD/dxIqjjuonXXdRWkihKQ8dr
lMAux68nMP3ntkc9F+ctvlsMIL0tsB1dhr0SWKH4wFI3v9MERuBDECHIRKF5Xo1I
Paetneh+PFElEsKcHNWE7NnSuYRq+EeE4uFVSuJxNYzCUuNi2yqL2TEhl7wes3Cq
dunSM7kFfEtPNTKqu/nW1ayKAYK4o+rTEMLGESJqcKnekItv+2pLBC+pqlg8eO+l
rpAEjkGSsRocYI4yqp51H9wilth9e1/LLVo72JbWo1G+dzw3iEhEYDgUmF4c/c7X
lRq2keugzJ9mACJSx/Mrs4NI1cTvE/3LD+CwNoN9RnUhgIFdSAr3I5FtMBrTz89k
uYVoCRp8z900gcd6QeGAYboi1U49im+oVy6i612+t4KUix/x69HCMJtWmHqQuAsH
b9w29glhf2rWjZinxvQRD2o6ERrTuUVFEfh5Nj1GmLeF2n1Ilxo0fz0Kjn8oC037
k3GOz3LymvflLedMCqgt27CtagtdGP6Qx4kIgnZW3eg0NDwrQ3oIF3XL+xWiKOv5
3QYkJ8x3uJZgeRvT7tZmdMf1FZXfIs6us2U7yrkUNqY4sR8pNwgXqEgCGHf07rUM
NQ4lDOM9ETDuqq1GmRiKhtqgVBVnzPyDhFZpOLKTPu3Bf2joZapHAM2M1gcmsFub
tHideqZ8QVyaiWn9kUxuVzk/L7nSyWkoU1iZYQeQcWTr+7fJvk7MCzHXJRqZ2RNR
rbjrcnl/WMTxOJAD116J7/7TkoIFpFuRktG6MF37jsB+ooGt3QEljmqMD5mmcLWw
m7CExjbcmDw9F7KV4EFT2+RwOi52ONw0pi0wiNMB6So+SHNNmWqwk8+VWKDQXAQm
dFhwFH4t80nHX5p/hGt/SAPHz177qcRFcP96mJIEt5xiDPkCQ1Q1DhSoH+I+4H/d
3zZXvXQDam1DO+oYevJy6fShz8/1Zok91ojd+kgym5TK+HVWGQ3CA+ZfUD2I8iXa
abDuCv1R8eq0jF+v7T/4STICnWrtVnEY4juyzXm5G5MOz+Gc0uySNoTT6xJB2D8N
K2d/y6drZ+17bjpPIBUZSN2SPagxLbbEdQ5hOrigJF/HwVMEbxx/3KTNglP5pc2s
XrwVRi4Px1Bt1rNqAStnxBqmH893JqMx9NuqCbYl84brwRLhIsLvog6lcjgtKtdu
/zw+iT1nMbqlrPIZYSsO+d2HBZ1Scy57lpl6Nc20KE9n3YpWZiGe5fGP2zYAdmaK
TKg2aLKXI4Uk/2a1J4koGPAggKmExXlNfsEXzsj246sN5k/OAStafIM1LDbq4NVk
4OQLdoHiOp4AdR/XDNs2J5efYKwbdEPHYUB6Bbx5HFQBaBLgbjxCJhKZ09jL6XMR
b6imQwBdBW8T4MKowrOf//RRLfgc84O35WrU5FDMbS10h41hEVcuk7J9bMSX0EAd
tdboEJtDHn0lNw3w52tKkOXfW888EIzTpXiOOuPtHTzgTux21+JjgNIrtGtW7gQA
6xBqcSlnsEr6IHq1KytEs9vrWAnc5EhqpPYck7tBOak++4yhdksuD/zgMBWrlh5Y
ApWk/tIsRzpMCepw4qM4bgpN9O6IhnP8TA8/ozHr1NME2phKLFH1oeGVlvOBigWW
l14aWkOKzzS5KvKs0cmcyjx/NJ3u32JYoat0i+nAYmz9zlquYe0HPFOY18gdGFmA
C/jQ3OevtjI4NkVbXc84QvkIpDbjWfGTohe4ySqX7gxNtQUVcztXXFZV0o3AlBUl
U4RIs5HyxZDzMYZGIK5bU7LFFQiC69frmUg1OUXgt1HWJgqteHkEbwXucEaRh34t
PCxozQA15e2rBOfhE5C2TggJgBeD2rxuH5QNAlktpFA+8U7KdBjuNhDO6njsRvWQ
xjYHEK7j5MZwd3+POk0VJdAu2vr0GCalA7+LKeSVBzz0Z2chs2pgE5L3mvJfVazX
TwazQjbYesrxsbjza6iGwVmGHDsd0b5RSX2eSPU90xQyq1yKCwtMtlkDun2I0W6D
mULzcrGuaVm4/ozRu8ZvS+O8EGHSWdut8dpERongBYDGnCOOXtKubExr/f3ndKD+
U4GT9+b70znMWvaUCRKnjkxB03z3QL3/UNxjQfsYop4aULwT06n/jGVe3ItriOvm
ZhF7h0dV7968ciMAFFOyIywk+LPIJoRjGitQPGdIM3/2wg80pEchVFlCbFIf4/OB
MBG5oXXjCSHIug2DBHlrM7qdR7gwIrI7OCSkp8FzbjfSTn9z3Ko+YklxNXV46T+G
71fOexZcYOCFPLD0l9MdNRDiqTDlHuFQzuU6XnK629XaWCOmejOy9Ogv5k4rqi+M
nqB3/3UuutoJhmxGeT/0FGFS41a5lyPpGedS1s4rLVAVRRlPaT34uNoIebc4kJq9
FEAWsfkl5CHfe2wJ9ofNyQdX38+lDBa7KuAlkB9wFxZGdXsuKRv48JbrcytvasJA
PVKCCUsngRl+inR/6qgu6SUUoUWe5mGKVhjDnKsCma9wUCdSHK0HTU7a9nqcn0Ct
VDbDeVqIdKqbQ0Bt2zERfHn90Z3J2wjQd5n58gv8oLZae/xTq85Z1tx7bK7NGoMR
VFYTkRcxlDIM82E0/XRRgoEitA5NJ7Od9Awcx6dmYAuQ8k5gbC6Bji2npWqKIA9B
z02g6QJfujeTc8u6BZgSm5D0Q7lbq0umblEwqrkv9a91zLpM1vG9Hn3+FRgPmwub
CcysoY0h+lRtinWv1HI2U6WDSDNINHq2Qyzl0HhFACMffDD6hAAuINI2WE3YWJFP
3+BeIjLwN41sRseJh8tNgtn+hD6p4HCobyPNMvazqGXiA5CD3RBveiuNdrtrxjEk
V9veomaMVYLSFl5d8ktUCihaVJlgS7I+K7Bh93pMi1Qq+8A+KHl6UDoShmFzUCK2
QtChn9Yerr47XeZHapSkj5UiiPWkT/g9pauTW0XOk0toptrb71qvRQf4CMBCFjLt
F+bp8Oy1/DMQNdvn9Q8jyLlKXZWuPwSIGKTcycJ2kEtGM/XAYKOHMLsNMvA/9Wik
3UmYOdBKqpqlgcsjv5DlbpAVPsXrGzXwkQrSOorM9C3yP6pBLdJ2RXgQesCBrSzS
50axDAUdiQk8sdLrAZVQ4+OY7MFmLLYoSYbi/b2RHYDLVTDLQUNBA4QQnF0yVK9R
X3t4VoLDTVdldw+nwgSPKcz6xUouG88mTrqlsA6w3AVlQtKo2BX5ifhbH7HJu+26
KqNxXtgQf07kJ8NhySdmaDuwr/8lXvwgPKy+8x7gKgf2WmHSVSyWqAE+JM16tx2r
qfVbaAe3G15YGXSnYUT57doXJMBQ7fEnSSIgNfC/+bAd0vPmfP9rHMDy56xHLFkN
hDMhg/Vx3lEEFBs3IqyY3EhJMSfOLfE5sVkV84WC2PjISnLbyHLpiyPPYNEMrOYB
nvgFBt88aUDgaNKHAytVeEPzgxcMZshnHYjvEZPSMiVgEZgl2Djf1uj43jxCB9gw
L7EykLVKfZyWaUsQr7mFjVfj+0XhbfqW0jVUCgczWhQqv4fHmylAkvtwX2ntUXvY
7stCVW/2tGyduS+a0DzksDoExft5mCARlmv6qol3SltC+zmgM5bcx8Xn/VWOd3Uq
/CdIE1jfrLZiANsyu24uDJlBu6vnPpu3toD4Ew3Mk+m5UGM5fQt/ETivZz1ja9z2
gUHqcQ2/meEVxGLucHTDnzlGp3FN2s/Ma6JPdFyFhQoWx4omnymOfYZa2iOi1X/M
/HXoybKq9Yqcd364eBf9ykNdVV3/Y4Bw+iw8375PDi8o2o3YSDU6oTL6f5zBhtsJ
vWNiDmcERY/7WXdWsnuG6L4HYhpP6PZWSL2W+tbf+hoFcQpnhYkXDIpQkoZg6OR0
XJfrVa4l3j9EFNpnhgTHrAJcpXCco3t0gy6fYtBCVAGQyEW2W2PuT38EdwBaZT5B
PtvjA1ahsZA96dyfe2IJFc9hlLKhOVMTi+CfOkYzTEZM1ssWtY9k0RZY/9AxJope
PzUy3dF5VswziLw6RC5EJd0xxYegyzC6tfWNUbc5/d3z6rs//RpunjwOM+3X36cx
Pbl0Drt1XVBDaOce8P669DlhgN2UKWIth4ks4hynXWrWeBwu6TfzCVHGxQfHWRBr
zj2x1410mz04JeGs2FhbfcVgLCZchjsfPQjJacTQ5z6xzr8Y1+VMBlYL1LSRqLjW
H00oudf7lbUnvq48+FMp3fmy55doB/ehrOeu5Wcy3FKSEYbgxYCYjI2l/y+lP5V8
YLJm3AStzEb5++XViv4N+OpQSWefYRxdHFQyNxsHOqb8DG3gI2ZwdMaLprp2SoUX
lzJ74mfoAO9v0UZDu5G1qkAIIzFKfLhsd0Sge8Ffuu9BrkIJNe1EeCZueokZutqK
gttrXVRhF7LrkWj2g66oebZx32hThvXblQipGuyF5brxjBwQkrmklM80AnuPsXiD
89HvHSuUeo+B6lT+XVDKjibkdYRRvynDwOcpiQKtKUEI2GEXyGU4+9PHPogv70Dq
O/nNm65jCMU5wp1qXSQQwV1JHpo1Pndbx2L+Y1+62rc1ns+v0hFc2PenW3Db87Dy
V/69wAZJdkx8EGPF7HZFX8LnZFuqlwJHykdGOY8x9lHg7Ehf6tnxW3z3VgmyDK+i
HjSPolAekw5VZEC1Bew724kROnypjj51A39qoP1/oWnoZp6xva/yPzJJH4lWIO7T
+nN1K+A7xtZ3pmSMBdScVQYig0Wth8tFn21OydqauWBBk6DtjPioTC0RhmWPsbUA
fLAFjEj/KC2ohh+yizIQk0FTefXI08krQoSaHv69fV49Q1+4xr5cqlDLXNgGgOMG
8erLOQwQyAccanIDQOw+2zpYDPF2vDzGVi64ezwufDbyBoSL6lMZjYPZCBLFLiVV
L+LrL4Q21DSpOWkgKs7An8btA2f3jE0t3oEbTlYqzGKwkUnMP7M1M0IDXcSxOZVQ
RIF1V+7DbIBCNBzESTu9jrjlNE35FgyDQ0yQTYtD7MJg5pXV8pz+nY3Md/+tK37R
7l16X44alZe3edwmj/UxDItLKdBVAoMGt9jiUa8zlAuMZHqggYrLLKgVO8VzD7IU
uJyP0EdOYN1dpHKglWeMCgN6pXzV5OtDQcKNRpJIhDn9SF1YdxgXc5g3Jp7QPtuD
lZXdnBvCTl7BV/3St8EDD/E5Sgj8HMjqyyqCafxHOye1kGVjDMOai7sJDGiaI9uY
lH5p1M1LKgCbE9Kd4PBUcxGAbOmSr0qFe+2ZGDjRMLJz06k+rJD28HIxsW6slC/g
m+R0RtMGDgH4mHs3f6MoVQHzCSf8ZEsuJgEs2SAUBvCUYjrf44ldAEEY0GXvEkUq
PY7aSkg5JYQ2rqAqmSMoBi/qkfKjozdR/646d7z7vepEOkgurqmc2lWK21flbhoM
C2DD9iqD58C4rHW/6nnavXAaC/FS83Ss18ajpYT4EYTbrHmwxPEYs9BwkfPNip5R
QkjncZ2emxPr9U8JHVVfoAL3FePMU7FmtMlZRrbGU0semKeFpL8u9qBG2CrCrNzO
vCTWcJi7q8OsrAIK4gizh3GGzCnUGOR7Ul9L/3p+cJl7l+iytE9AJUiM82gSV2Te
/NDlZw+Ofir4FIdOelGO1DJGo/rb1+JkyQOxQySjpTnlCBeRGvWq9l445POtxO3b
eLYUDKtKMDH1jBiqyfJeBBGBpZmLAl1i5Ela3T4EuOaezGDflw3j/fs88hBsAnxj
IfsrjVUkAVCroWj71cBuKqRbxUyK7gDSSUMMUkVi/fxFyDEiK3p4IB+X4guAuRqk
m13cvKR9ZE2rK+S6CXbeIPl3Eey4obWiaeN5IFHE90sq4i0umRbVG1gHq8Sjqpov
BWNhoALrO5VsvgHAUlkwWcaT9qeHw90/Jxk90+nUFh1eFFsSKWlse0ZC0ncZMVAK
MsWXN2kyMFc0FPOqrSDF+qBe6ich2fNuSXkqyzIk8BAdmWASyIFNbrj48Pzj/w43
PvJuIsQEWfdBBst7MMnI/Pjw1OA0Y1O6NBKt6PHNFpmDNGXqJj2MCJWjTMTdC2W+
lKE7NFqBelw6RRyoaQ9ezbtWS7722wp6ljNlGcD3clkAz5RQyjot5lvVy2BqytZj
3EBzp7cbiH7DAJ+PhWX1Mm0+6S6V0E9n/d+gf0d/gxpY3eHuk0HBW91P+KCgiuFg
bjeqwT6z+nPE6eLZg/+5b1DL8d4tsedR7qdY4yCnAH/Coi4uovZHcgzJWUlS3NLT
wk7jknBQdDU1jSawd5yaQwWvr4or/dDub6OjWyv1RPOIYRJoIUab9IVCULVu+s1v
IAQpwstY/NkzwU3wvEE+On3dFUskfIfAwGNzilVfNXoZOYG8VB8rzc75BiOZpd1g
MFaZHqpVrL/WhIFjvYhGSS/Z5QSPBql5D0d5tNyYQ1+RFS0GExXnfFlLaQ3W5vxo
q3B7SNMMHSTnHMQfcm3n6NFU+kRzG9WVWZQk39iDl0/1E1M8vLRVP69quYExy84Y
QnKgtBpkDoS86iZ01W+FKcs693BTnNoGAe6en/sONzzINTicOluPlxsFS4FMEIdW
Eim5eVz0PYGYA7Kvv5FW478g/GYI/m3E6vcveQOjarGt6ANn5vPAf28M49MM+zKW
KHTQYYVpk9OLNmjw8/gQa+v3LrxjU0pu+Kxc8kDBbVRqr8xMXRy5BQ4VM1rg4iAJ
sP8hVCk2vOLQJCQNQLCb03OHkwR0OLK/HC1tjJxmqBIypME3NCgI/7a6tCVVG+Ch
LOB8y/LT1kA6jyWc/FqepF1Gi19ISuPkIGz8fjVW4/UcFxGiSZJ0vNQkgtUEZuoy
IIrR6HBv2/ltDKkblq0Ydr+PhpQ+SLfExozzIto5PK9JHVoycrG40D/HALBy93Ut
8qMMo82XxrGEegfnvA2/lO+7K9+ivh5duW6gK3JXVXna5J1BYJtp5wyQ10rkkdwK
oMBUaFsDJ3oKgrhJfXejUBQKlFjIwHBrYma+LY0BIKAyo2jFVWN9nRfP4Sk5k+NJ
xPQEieBCTLcv61XlND9oo29zhFRsdGaOSPhwegUPRhQmec/K47K4NNbR8h6KdQlv
+G8hF8rjEzeCF+4x1qYElmtBa1kP8LUFON3jhZa8s3w/V7aL28uED24phVndKa/L
sAvZVcnphaqhlzrMahYcn+cyi3Aiwzi/1+LlozIUq74QcNYesrI1KVmQjzk0ERdT
6IZXEte9VfxdQYCNVFN99BTN8O0eynY5y1aTJAWF20Labp8QHeYxXxDS1KLded3s
quIPbqb5O65niWRmAsv6MK7zOsimwWgLN9gG7+SUBLnPdDT8MPzq8De3HVD4xbhi
4ycheRDWB9sxqdit3ST6aWqFJDqZP4VpeuIv0wTVj9PRZVkAne5uOmgW/3a6eda6
5fBjaO+sobaFuLav4lEBtFw2caXcQ8LWCPrbhpxDo46V2cnVoJhyzRhqbRBCkuYC
06j5QBRcWakhP3LSDX2mNfklW+xezrCslBjjeIucvXHOMziubZLFOqLZ9J0mNP8c
BPBlGoGK0VlB4hzHW82xNhcm/L/P1HRgtJayE97ANrw6fy+gHFWkQBmJb+fwyVe/
vmZnPDIcsfOC+BqWIKaZHsINYQeJwzqd7hCV1dNK2FTPokLLE66N5D7VfbXINHTx
4SSB5vEpdnG2JsPxmi+dUfiFHgrdA8L9Y1a1nOmbC0t8pM04Efyg88betoBharK4
ntgtYBS0UixezfyrNUggWH/HhXweW5aE6nylDrmKmu+xW4/cTQ98uHiQwWxPKqUH
kZjQ+GERTqYhvbKu584VtqMho5aGL8EcT8EuEyn3JGzSYLwUHJXZnwm+LDCREKNy
HzcbmZzHrxw/2arLK3Yzss5EpoH89cFPym+B3NsOCVO2Ls1kO+KtSL6T2ojyC9PK
g8tmAHN8O0B0uBo8xuM7hQW9OaTQSGYPEFuNm7DLstqtMdhmV6EHGtCqwVmNkUER
kra/wIlncNocYhIJTT7eF4+etvmv/lY+5Bgg2+4n3n1zAdoa3064ZO4U5l8jSZIt
DjrHXCSqQYEUFSRq6TlC0SUlieV3AZgk8722X172i0FsI6e0G/d1Q94hmUILXFwQ
MK2NrV9DOLTzDXjThNpZbU2pE7QEDyEtMcXwsTofRkUwE12ODB1QfOOl45MQv5vq
PuYtjrLna+3AUKiIGkMbb4vEdXufa5OPN+W85cfRiVGhWGb42LLtB8LeOCto/M5K
CM6pcuEIDe9RehcYhTRnNaAvN9DxwfMFlCCT1jm9nh7OAeym9Bh8WCL3+EAS8h8o
gt1H0yTQp12G1CRz4FJh9N78dAlmZ0LIwOx2vZPyfeSXDC+Ub2HWudvtk/jrmqg4
zRHQpJ9vSJdkJ0NJ7uOIisXuQEHi8gYchdNW1rPNFdGqJrHDUrP1SitigmbMXx4C
opI4+gaiCjkQdcuujD4StKpmuJUv8JCnH75txzGcJKFZPjvIalbdTJijBc/wONxR
XLVF+IgOdwRYu9CxnFUKjBv66oTAzLvYAqqAbWKt3O27YAjv9J5Rd1zXkPdiMDpj
jEoOjWIsTsZesRYbZQZndB3ca66DnCeAzmbSl7PIg36tTpFfkbg5Jrv44DKoZsZ0
GuV/AilvtbHXXwuCfX9ZNcPIkBLtrJQOWEAPuBYVy019zOX0V/JXBMx7U7RPa0mJ
3bIpy4GhKFk/RBXcNMd3S6xycfYCx/jFnrEp3ICdhfc1wjp8RUu5cQC+4pSTAVJU
n2A3Lo8XLR2+A3KOOAC5jGLFmGUcxnMiGVdchsET9BqgZQ9Pfui13xSk4HwzV2hY
GKolcUtYh84V8OnW53jjGEDP6KIW0+xn8A53BnvbbVULlZWuMNatXarKxbo0/O0a
fVUCqWvzFToC+Py+0P3+EfKoa09ANQcg6FjrmSnGLuHbG0GERtt3WNoKD0pqhmHd
ktjycPxJ+n+Y622vZ1SaaTVtNaG++EJ9r31Pd1SyOQAVCP8LeuTxYhWWLrCqG9/I
ByzEAhOL6rJ5qMhuZSEniRH6zVyteOxks8+SFRb6HDJDcckG/rFpL1pySqs3zyLN
XhsvRfbvYWaYeVsazX7P54sRnOHvMmwHB/VVHgGi+TNXJLgIyXK+pQ8zNqvLDtOb
jX67zy/YjA05h6/rbnhDFhKr6RtiFdgoirxN1MRmeQRZsZoyOMB/+wWyYXfUD2Ps
x4phopjw7CJ1OYPCacpMCwfCUZh3e8dx36z7YSJYhwO58rnuXNWNrGFxDEhbiA1s
u9+D7VEY58MltYrmfWpP/pco83yOmNSsHteoVjySaI1IYQJg4J5HcjOe0Dkm9aSr
YU3rOwhrXnWexubtbCNEMtnzGpyR39RVJuBjrh6n0edPheTAZ8A4kBETMytDOY2H
99vY9r26PDlYRFvg+ea4nbtCizhjdt/3rWjqO64SgaTE2+jUQPYTMLBOhVW2i8s3
mtEcbA2APSdh46IWtqNsI6Jnk2bjwvq2PaLzIGzDfvePN5xj9NBMullAIf5ZXysY
3CPkIvHuD3z0okFJZkKnKo85HLCs9HpyYuV6xgc4uG74g/C699klIKkCcqC5ZtKh
4+QunkeSsXwpnjGQrOAjbFblEfGkuZLbyvScaYauQyVxthz5v/omqeOZTkbl21FV
b/Oz6HXGuKef0HJjZpmXXV01aie7ralItrwex4e5nmjIXoYg0CSKk2xwLVdWTl5i
2F1DaAKPMnKJsyVCKess6XBM+Vs4aqVpMWUsK7P2pvKTlbB6F1mNuOL0qupKxGes
13Ou1iHYmw2M3kQWEt2yliPAuqWXJ+a3MxEtWH8WWxmLhwoTKzHD8Mn7CG4bjNNN
CT7Gwv1EPwvfYk4MzYCC3Ep08jonrp8atlZrnaEg72IqJonZC6yZzVtDfXEChUIR
5FDSqaxbWCb/QeUE9KGZ1MG5EhUQpQnuR8P0z5lBHKMg++U4przYia8A2VF/mlJK
+oNMq4C6JDZzB4Gje0dygnpYT6rboipmhrC9rImq7E8GMyApaZ8c0ve7+mKTPp2B
jQ0+hVfL5F4j/AAYtekskz2T01nXOHdtk+svyImUtXktmB8b/T6Te5WuNkuPW7qv
ISQAPE1BX2ma/WYMGPL+PQnVQ8vM6s6WoByz2i/EiTzmYur1PXRaG4qK8zZbtm1M
VzVMWAi8S7L3Hx3ZLuUt7p5eFFjAH24jLhx4Dstn5kmbF70PSu1RqTwlXJccYGW8
TtbU9Ywtjzijeq5lkiXsGjtdwfd+rrBpUDIXWnZkvvFZ9x7HottTkRgZLtEq3YDd
zgKjYlA/BFuKlYux514YvkNcVSoE5MlTdy5NhK7AmzNo52ucvwSuzcNu9XWZTZHw
vtfgj8gMaqPb9u6hnCwQUUm7fLwRMqNgrBhQCo7zVpwiibiV3gfBWVcGL+o6W5wh
GjxsyucCZbAT6p5M1lb7/wWQ/H/KR8Y+8kmE0Zif+iWhmMx48tDgyySo3ab0ReZR
ylfhU7ryFwyvKtgRy+uIc/+e/KicfeTE2rP+9d8gqNTUGV4vwGoXisjt/UW1uWV1
Aip9ZDKWfFEEK6ELcuG7iAH+/IPSXYk1YrbIBBDhe+XeiPS0WkBtyqtz+xQOpANw
0L09u8Ace7ZQb7bST8ai5PQJrDhuqP4gKGTV6Elfc/tvvrw0En8ChDPBfLu5n96o
ps6ZM/nSY9W9FnyCvGwXoQnddhj1DGiO48VtrhoYRKC0xid26Rjy6FNgLiR9HWxE
fwqvJrAbB+StdDZeHaojMetiPjj+sL2s6xtc26OpFQ8HWdLdSnn8OWM+uhFTsvEi
+yDmVR29PB/5EBTSZMNoyntJMQCe/oOlscptbJDk7db4QjXW4oAuK4bZzuX/XFVR
kxRN1BIbktqxy0MhEvn+N7Z6dnggzTHrINZ97jxLWJ7VNISyuNdTxz7fC/KTxfSV
R0cppLYOqjcF2pvEbTPIrOK2By4RP7MDiKH/B3vhfS+rosRVkFNNkXH2epsFMvRT
yla0qbKJ6vrvZru1maaAKgTBYMlpdq+YgLeeAtsqXA7RyFStICoMk0ao3HM7Ktiz
69oKGPmnUyGSfKJF+ug9SYul/egaByDwFtwDCXqFkuFWD92jSuB2psJtMbIx+OJF
fry4pk7NguNl19dXlSI6Yvr9DPtTuVkQVeE7p2rEc4oWuaa5Iwsr9xY40amL38hM
P1PnGLzg7/3UaYCXKcQHKiT6GLWoPwWfdAy8d08wzqUjy2bHxITiQZ6/PR3QlPA4
Rwezf53NUMMXpTLa7F05Mu6YQRXcgecsQPI/KoO3u0tgLACRkoGGaYKMgpFMFKHW
sM+e+BgMyxYq+hFnGNwxSkmT0xmRRiDoUKmbheOaWPVVzVMKYXE9bnSGUJigidrk
byfCVFEEmAzhvrAGMR2puOtlVKheSSObZOVTd/piT80k3pYyYIBtZimveQ5u7OHQ
Z9btTcqAw9+fr21l3zB2rNb7fxuWVXVM0aRzT1ZLK24s5DriDxTOj6imUsij6Pex
WF59qpgl9dwV4sv18bzXmpsWL9kOTeoYYAbayBHtedNxweqh+4cKCvyDsEczk0XG
+fUkhatCPF6YTUKmg5oQ8+PLJa02icOiliWjJI94Yo4OGZjYsZBM1V4YfJY0KUla
6nlPIvFaPyz5276Z9AdxvS4MiPcwA49z6X0G1CVJEvYh8Fxy+eLVz0+J268FMaKr
sT382Jzh0S83MtvprgoeTEwN8l50egfJ299IziOwgf78Cqd8wZUgdSU6LSe6fPzr
fBl2uYZfR+Yr+VvTsnBbmt82MdVLTIzCduqf8tCWLR500TIx61RVG7qWDbeAUylZ
zPSKirBLEbAsE/PAAmlvgrWEFE45yizqcENhMnmvEEHwk6oNuSZG6cWhYRHPlMyh
+/6A3btQ8wd2AKruVoy0M74hd5nVzyFwwoLIIByH2tQTEHxTgzs2+rSC3OrZZxTQ
Ue0lP+yDiI284rc3TIHGvFDGnxbO+fwkgaWaZS63mJ172EUS3LOL9kopbdPGe3Zn
esWAUmdiuQmBdz87tSHpfsqtU+qFddv+gdvDg0ohmIWX2bUes3OnxMmt/N9qFBHi
LkfA5nc/U/y/mWkr0i5Ch7LEsxuS/ObrTxYDRSN3mIv0TwASlFPJJTgL9U+NRMgW
MIMZs7GuPemXGT+MdyvoJmSAL2eP5cou5efcm8Ti37wHe6W461Go6UV5/V7prBfe
fggBCafsSRuob1Cv3dV2Tm3NIjnKk0bIYK3YWL1PX0SFCO6ZwGSrVYyQMgLfh5Tu
xYjKfk4MlRV6A3vX2+PduBAh0mecy/ajY805UT+k3fl5K8qV+D8jIOrVLGWD+xGa
UExoPpXrDcCulYAn8f3/onI2n0ItWUX8gQEtWff1CAA+1kMdcoZ/D6wz+o+wXJ61
1LoCKr3Bw06G35qYsYrLPVvlhMThAR4YnkrhJqX4uoyPp/nOzqu5ObQeI6njrkvM
w8E3/oQlXEBf93lBJTwynlkNYG/hOBaKMs0I98Z4iShBX/pnUx5TF8ErWsZSbtZx
hvaGtn0IQtZjG/Yt0Cfg8f1ZACtn22Dx7BWOQvFg2/KzMYj6ADzrjYsl6H3RLLHo
+bvY2wk6muhiaC6Ym0aEdLIXxla3xEN3BZzlIMJ3DWNIG9RdRVNSX1mSX0Xby0qa
P56MY1ZEnGLddEDAXgkPJrSBxCwF7N7KBshIHv7s/ivVm1/ZIkvqbe8vI1LOfe26
WwIBtGbhG0Wmeno+HFxb0R48uF3hYZrlSR/IvC6B+IhDGZaf4F3MpyTDQsz9R6q1
DJhgYCObXZdHtzsUAf0Lx1oAphYJ0xghwaVAsM7dsKWe/ZvsAAd5o+qCNFGHF+7i
Uig/EHpt198rPSC0KT5Wa6Z2LXvrq0O80DPlZz2697HlvtIRKOb/RpyzPxlWCLvQ
PSJFOVo/6H/FGOu7wfQ9YlG4K6o2ct6hvIFHd7r0Vr3jnGbs3ffd5VU/YE2CC4HT
a3+1jQbF+XpcKvpJHWQiw5CqDMsJR1xFLfFySUkv+l5+J0fapQeoKvAxtKrzW9fA
ks2dW0a+XHVQTnXFZE6oQX/KCk5PaI64qJRxkLV8DU410pqZORSWnqPkd7LLSM2X
TytvwZ1/3b4VA4Yg3XZ2oE0VYtRPqg4gg+qcDRsi9RR9UsW6uQeope3dFfuWsCdZ
5/nP8q/memSNKbbLIbHO5qyRph1GTkDC4HiRnwKfw9yF+qm7APq2PlFCjUrZHlBk
KeC+Z3aLmjJkGIuHa0q2Daffr5zes51aiZ1YitknzrElktMJ9RCqMFYHeFhEu3aM
YpzYeumhjZNoJOJwMudfwzxww2JvDY+xsz/R58j4CoO7X7bk7ZOONir7MLQyfvQk
r+A27FbuOgGtoLH9cUv618aOtnBahT5bLR24pkDb+sugeFJQcH2H34T9jsAGcTU7
SHdJStpHAxD5URkU7kcdnHnqmnr4QGwRbVohPdORGiL1/ZkzxcJbSHg99pAque0F
nuuUfME8cZxsABAftxdQ+9dfdfWrrLuCWC8cTX8H/oo4lyo6HrJhoaUnPm/NJcbQ
doENd1HJte+V06VcpWW+vnkX2+a/BBwZXyxAIS1TLJqRwXJVLTiI3Gv1hVawgHDe
bRhWOX51k87eaqiVNjvA7HIS9+DhciKfKdX8x+HswFttTNfhngNt5zYGEa94xhdV
pvnx6c8RfQ7Wvac23ENogCHoqXrmo9k97VDdRLm4qRqUzcd6pDp25lHI+CN/Nkms
JFeWf6Ymm+ai2xD85ylMnd2DmAY1HMGHM0hSMuvJR4p1iIaFti/aDRTITnGRmWR/
YnH4sZePIfbWCJq6DPMzsh2aPUGLFhcS/mEtV+tQtOSqznYxBkILGyF1Do/daJqP
8B4L6FoCU/3UWe7zvbEV9H0+quPPNmjBGK9sPR2j/Bh59D2bUbw4arw+GqM0w0EE
CBpp2u5JkQq5IUOXBmVj4IPQrndKdJSbBJwqR7e8Q6qSi+Sd8L+1Y169mZCpN1Bh
ICl0e5nQvqhxjlQoP/7JTVtZ3qq0BdKFnthP+JY9p/RvwMCUXHJrTXoZSSGePNLw
kgJOyZA3QJPPbCi/EAnKmhz6OSupqY5FYAOaXU/4Mfik15lK9nsAx6OxsO+0ucpQ
vD3rmuuFX2RLWq9/VvWiAILeQQcXMrcGILQflDjwR7GD0Vqvimqex5eP67RJIIOZ
B5yx3MRjjAeUNBAfaotfakQX/RSEcXsVSG8VOxdMb1VoxLwllbD0RIBpovhb0AyV
fHVHR1NZ7cQwHX6OuXBfPadChX4rMz58oU2TkbAAz/YZn75Do5chDfmw4JRuAHsN
MlgK3h+J/chIA3CwJswldSAC1+Xwq233eSaGSRkrQignuvGvaKHPO+CTEL5zZnJz
QlKTk0x4Ouc0aVfmE/TVpbjboqHm8FBJoYrgdS1ARX76PuOWH+clVGe69b2qGbvY
RAQ/cDvZ7Z1UitWK4BRqbqugSKxV+5xRgKsmfIKeMQEQdjXf2ZMgLrQk23XMbZpN
RADhA30RM1+ys3CEKjDGVAeKg5GYe+WTA0QBKzzQq4phSLftyFsTI4xeU4EcamhI
1/GbefkCB5NlKiS3MqRB5CAkJoxWWgiDj/9vCjQfKd6F/yWzxfgs9FHkfy0ONNJJ
q/OD6ABvj4EJdBdKs1lEj2adwxXvIGZ8NqBiyd8l1IdYWW94tr1iQ3Xc7DwLcTjv
tTBiihvR8lQsqNalcD8c2IINSnPs9/vuhpO/L8P6wjNzbFu3LSJRHwtlEcJ7YIht
E2GjDk2Joo6QfCVDmSsZ5whn2AKb0E56uCiIpUE7wMK/sh9v9GeqmXfmeKAHdL47
qcK4fpgPp/Y+uZVIEjHeTnHkgpDfdwhslmX6wKc/xzI/xKx0e2uGgn+dbW6VTtFB
Y/jMDQ79b5bTJVvUHdlq65t/nkB2O5eqBxPsjJ2lK3GV0zyuDDWlU174tbD/lAAP
I/m/Nt25bVjK3sE2zQFyd1jJir4dZi+Uho7GTP1xRweb1hlyLBiNfp4lCUKnMfpf
ONTniL1qwPNir533Vuqs8FXwd4sfzLttGbg4xK5NsWwU/8LvKzsKKVhzjJu6MxQr
SwqDzbq8vwmDg9pvPvfiOcIfY3eQdZsmOW0SZPCYrbw0SiIJ7e87CGg6f3zIKytG
mmm8MTIydDspFCSmPMwCgi2+OBkZb9HazDT4SOjjfzz1tz/XALyNRwx4gtWOM1N1
JF9rYqqkYm7dAefPICeRohMXNqDo4bw12cnAUfgvHmd0ymCU2rkg9Up6RUjzMVaO
3hre5b0zhcxXZYeZs5vmRHZd834vrRIatBtM92JM3CiP08qSJyY2szN03Z+Az1kO
qoLjvR9r8mCATzpXkLPJIUO/6e17jcvXJaLd6eHKC1yreNxCk49Vqq14qkdSFEOq
2TT53dLXUPUeMw4NkfftIC6Ed3PIWZj9E0Vtb8rUakLjNi/q6m8f/enCtyBEMgYR
PnDi3v/e96KZz7BlQ5ujqnm78ff3hpeF39hEs+NuKvm0gXQ5vKNfkARKBkUr2Mpk
tqk/xdWEV3QdqO7jhO/OchBMa1YwIPHqsDwFaxVxDznWK+XAhmhpBOMHpsPKXlqk
bPCCpZOluFCS3UyUGfOtlQJkKr3Sk2l1qUOS3OK24hSlqiOIM486Y/4Hbo20TgWB
8mACDohbZiQu2xPPusJULzL5ieJ8Zhz7F/KNsFyuiHTurpaOeQB16u46D06go+u8
OXga/psOSp0pYVgnBfRJdntSIqk+g/bY96hbrjpv8rHbWP1Q2JpCvT9nrOq5pKdk
utr1ytuD7XCvp8MUg0DU4o8E9mSlf89EVSUxNXxxOIgXKkbk/NYd/0aIr2enJoZs
RjC6foqmcpxTxAjH7DPTV2oYyY0xByvN7u3gDvdtc+e1ggY/n/+2MgEd+sOSPZQq
Ky9Hi03AEn2geuBRA0GuiS/thQmLCPtlUAwk0AMS/Orcv/qCbe2W+cHQOj4fPfBD
pPAdS6SirXZXGffxumvrCsdxl+jwhCkztJ4B7fq50xoArI1zl44U6FLIlRFqqY8n
kVe4ODWabYfTCtJ/zwXbKfQxR+dERyq4p3teGOYy+5j/0iH162YvQuMYDQQCsG0S
cmh/f+hw87vCyUjWQJKvlN5Te60uaDX9Wv09couyEJ/8ew0wEb+h1HtillY9U0gO
OlKr7PWBNeKMaf7plBa+D5vpZypR/Mtne39s670rHFQqLn9kO9v3RdX8EWv/tdaf
UDbw4XwCNrCMX9O65PhBY9eygK3VRZWPjA8/qNiqmwf1/IcbACRDYhby5W4cx61w
12xBe5sYiOzVHIF5m3EWzGxFCt5FoJDQIpLKB+qHESeOved32cWX4HLMKU+uzUyc
l5xzczCcGe0ZoLb70TkFqbMaFEXSmycWSxOeE05wtwSUAkSsknu4fIo28WiBQNGq
PSMAcqdo4tMAfwltDpyTfwzAeTlulijAeEzMy81w1WCr6FLX9YtJbWVggK2dK2Gc
z3veniatJHKpO1Y524qhP63F9wpXqAQ3MLWizTVS2Bv33SC9a6a2OH1Cq5nod/ED
jOXGz4V1suUKSZho0kxgJLa9/+k60N1mBEZPsCgxnRX2l5YFOPwncDWLXwH3WBpe
9nl9m2FXD5MRbuBkw0jlCEWdaJQNNIGm+9EavbrboejF1kPT0p+9c8XZju9SA6+d
qiJAcClqXGXErJ7MIbYrx79Mfih8J0Dl1aiqDGmSdTWLyoAZS9EWCG1gZQ7xBZoV
vYCOAjbGkoi+NKsEEUKSLwMo6vtL0Q9iPhwlwDnvBRBnPRHkEJ9A/H/6iangh/sq
qVzFXdmWyTUZjMiUakF5xBoG8VBY6h7TYTqniLGMKcRbdVbizNFm0jYtaePL2+qZ
v/irCiL4gVSQFNKAtlFMDBpix8nKQNrRBVuWtTFJlwVLNy433dczIJrw5Pq/PKV2
Jxj9bKuDl3kGYYGXZIHhOPt9rMjxGvx9FTmO7cc/Mumki40zEivm6ew+s12aVKBs
om0NCelw3zLleBh/OfUB5n6Qt9F7rDkbSxziO5vHIszjPVWDzgWzjsCgxltl0k3B
e6HQ4qW8wB0xXRM4tkZPjP2zQQjxdAuVXgCREEigVCVX2oe6SXN4/Q3z/I8QvryM
u888kpttEBlA+pBeWzq16ojkToGeLORF6vVdj4IrWO+8Rs2XxUqFow398DJ/16dE
TIwwor+H7CXhit9kVU4G7gZ/sdiTIytPXmumPv4WX953QKlnk+1cELUg4XDuLBwW
VbeYina7W0jjptRtY+Su1N+0ywQWi49l595eVrKxsZs8BMgFgAR7LKZhZnFhXxFR
EZ/TYFXUHEoANQL/4HKtxQJO9kLIrbBss6EvmmHhaLcK87qq7jxS5t087Xi/y5E3
iBHWwRxKRFv11uais809thVUqReW47Z+cDCtnzVU8W7BFMoVHSzBPuXCX1Y0VlSE
vzzIeyRldljiNWYgl+C+Gz8wLguzl3XlNOrLqkFybcyO11a1AJpO7Sq5l7iLgFAX
1u0c/mSg1Lt0ttkHVDd6pLmfkUU084A9oS6dwePCDF5ywVnhXMBP5kThRRjrO1AK
Thaj/o1qk0Mk+vSlZREzbJK20N4f+r6puZsWWBCknVi7a/asRqiR6K5K1yWu0xgr
oACUUFeyVJmRL8zRH9puu1fv5Kwj+4PWjBwMhge0veIt7SIGcPBPfiS0dpC+Ag+U
M9JJ/gvh0CyJnjtabMbY2f/efF62xCLAbgyzW0Y+L5IFm8XbnTLwue08DNN28fpl
1j3XtcBXgqh9fkHb0IPxvcgTCHf0lcc4dgUNFoBlOQMfef9ydYnkGrCw6xdDIljn
zYN5GZ8HV0thczrzCZPhYIP3R6sHINwRTHj7lKtIPY989qy/O2b7jnK93JZo/zk0
jch+YP2npGNk0tl93Y75c/5KRLTerKrRuNEayHchWAZg9eECfqwdEfvG0go46Oh6
mxiQ85qnO+//izPZG12ysL1A0mca9PSQ4oakhlSQNuhyUmYjBvWE6Sc6P92JwXTN
7K1e31XLuzi2Z0WTSVlImvq9xDK7lmaWhds8If1lPM23ShsiYVQIyARH5xAdep73
h6BXE1TZ1OFQXh/lkxxe+i2sL9e6OY8lri2I3h3/y2cjPEx7s7s5ysC+GDTgFGTG
nDx+E4u9sPdBKPLqC5xfR9s50/1X/xJcdzmOmbJWCRg/t3dY067eC8DcRzIDjLSp
dgrXyCi3/7+GbYqJ4iA4iTsoEAdEaVIyz8UhOQcwPqDYwct4ZgnvjHtBIdiQqBJT
8ekYfZNtn9Sm7l+ZroxGsvsGF6WC4Dkw2TRnFBpTapRoyJXU76JDiMMZG6KIOhz7
d4RH6ap108IrTV55B+sPJifQ+ed6MEeLSboMRpjx9H/h01m59Z/RJoi2fj5VyKWU
chVQ2f6t0xvC4j6b2G0AP2PwhEoqwivpj2l3SXnfm/ZL58o1O3SdPM+RK053NvjO
FR524W7evzMcq1qxmnZf3IzY+8n8Q7Q2OgqAxDeX490dbix+cvPeP8dd2Ma+Hns6
VvqCVdvn4GTtxtpXUSNN17yDephuuR8MTo1EoIn2ox1fjttvCz5z+iWOJi9iww/X
9H7xvVsKM2O+stUWfP3Vy/oAPhbuIZNT9ZMvoVMI+SRDlAwMO2oCFj5p9lL0ShKg
QkP8oBYD6OZ2NGAePL673NQLXzWDB2sTisDWPHLvw3rSNE04gS1KuaP1WC0IO9MY
Xe28mS/8hyy+XuhWCfJGb2C2xZovZ7+US65KS5cQkP9fjFP6YAHkUvgpKOKssiE5
e13RqdnE6iOwte8IielngQdXljD8Xz2hwndZRC/pgK5toGV0PbSD99EEcHIGVP+1
eZ7ESaj607f0lDpcyrxnoiJmgpV/rWJXtiV8/vIxR74diWOqYt/+/6KJPHbSScnJ
52862JPxRcIKNkqFCVEzjtYdkdcHWAW+uLStNDTvh8EvTCVH9mBX8EV92+uynMXe
gGv1lUNapP4n0irAL50zvnmVtsUiP4U3kES6bP+lrtS4zXiULEqfFzV5r8XspWUO
oVrQSVOy+yDAfQx/LaVppTclreUU9tvMsdAda110IYjgkLCcSX5pU2sd4h9fFD0/
C+aKP6t4ocly5W+kGsbAoymeqOBrV2Wh2Duzgq+3b33P9H4w/BuCSDM3fmTe/EZU
elQchMRjfTfQAdeXg2BFHRteqCxEMwPzRL1Z6dq0tgDziNClHHbJuKMXAv9MpyZL
gS+NP4BL+TEjcL1EJu4k9Bk8kmaeK6Q1s57IHFJZKjDf00IKEB5OQFFM6ak/tip7
5uvBJuYTw48XXT6fNbCkpbw8HS6Q9a0gBuK8+gm4kVfTxO1+fbo9Nbmg0seahx6c
XbSnKfx/ZCoLdC+uL0XCRu/jGomhnjvmjunuU5pM6LFyB1FYZdqQ1Qz9T3Jr/wu1
Q1m/qJIM3OrmTFXIBcYFUDl0+WkYsJj/NC/MnfH4XTpQgPhaF1s8pKO61TorAijz
XfcFfRxHcwlQtH7Izvthp3Wo4kuZbVp/1E4jx8jFgww8nJlM4XeAQmFAo1/fx8Vu
cm3p1+jrutawyQggh+k2eKaANebcRGN1CVO8sSvQSvXbDXlqINOQp+NYakzOC63Z
CXHYf/qscRyACB/iS91Nw2te7JkuPhg5LQqUNND2Vjm1GbXkyYywvMTdnz/7PQmz
AJvd7DCu91q99iVJcaW1r9xarHMBvB82ugKTy0Ql6tAoz3v1LgSl1PH1clSWuifg
oteQlL5KzZMf/UnG/CmC0RvjtpVBWZYuVjKvUTY67IC1A8sAlLQw/lu2dg8CZ5JH
ZXKHO4b8VO8wnMmXIpVsnbFsUSBIzoGp3nOjJbrgDIxlkXaVH8DJ//2OJ0tBxAzQ
7j18NTNXD8C5GdHiMoKWNSPcGwzPusqTL0qzJigMxf+IEsK3BIqBneUKeHnAYKGh
nLZqUSpZAbMH0EYZVLqtumdTwMjPQuZuy2PnUtJaznKfEgmiSQ9rysu5QDjltprC
nwTNynvlCJRrOj/q8DlVBqeeea9BwW2/an+etUjn30gjoCFDXxnAlSla2gthy4uq
5rJhXddqr4dO0+mlBVn/fb8ayp0I5edY8+5VHsaxecM7w9eNVEt3vOoV40O3E6VS
1tFbqW2FVMhnTsawbYUlFeTehOkbh0At2byY1m2vHUHtNTtEA4GYaRXQRKfpijTE
vNd3hx973Re4MuAUugIU7jqTbsk18VAyw8qJiezbZyhZJlsGPUNM/PvXQyPvoHiy
NDrq9B+elMBcNrPNuQ1rIU9W3tcdokkYA9BFTFLgkqTWSJ/uDW9suZu+W44mt5hz
ysW9+oy4F/FNzzUDAIyaltQR2YXKyZUCYqBO1WvD21ygUiel7dBTrj839xXn6Bz7
x8hQi+KBANLBsFBSj2WXwpW6LLvYYTu3vZzvDc2fdioDhVOK+m19h+LUObf/1vkr
D+0TS8tmpfthqfeTrQQ85LKORTf42gxdD9A4s4XcUDq7tyZmPrfgXi1Cg6uGtXy3
1BNPjbusUNSs9aKfe7Sxw/OzwRlxxZ204Pkr+J5C0vPQ8T+0K6MsDTqb0q7IOubk
n5kxMIFB4Oxgm8sYjhvgcEC+YiYhWWP32WOXe8ExIXYEHwWfOlLPPHjbu90KwIFw
FtP8wH/xfy73v0R0JnfP+Midd2Im59OXC0Gn9JYOXTgx03JORAUvL7dgwClXvwbW
S1/ptzuLi8vIH5H9DJQbnkWEd2NPimA0qTn9irbyrcF7hY4IbsenTO3EETnO8ZvP
k3O1k6tREvHMT5LcjzjhdB26sElNUbwNEFQI3O0CVwJ9fe9gvetfNgt+rZTmLoH/
5cYs1RukzMjBTuDkRnH/GrQ4zVPYVjyDpbK0d4aCcv8Ui+HCm5bGrSHCOWCNQlQQ
XRrLCKigRHYV3TDb6i6ACHZpWR2ZDWNBbSsBPRaV9k7HvhmhWWBFcrCtsL+/4UaP
Ltan62uf68YGrXUXvfGcJ/l/52mrTAwhM1GtA/i5jrHSTYD0J+Kz7Fd5Pivfk9vb
seF3ErwFrBD5iP/+KPWjGNp9xw4u6XdmU61uN7OW9KhANcb7IEOu8qMFrq8SWrDS
d4rIwsQ+lFnpoAE/yBEtnwBG7vl+LjU8PW2srhb47b+XaB6bHWuLmpChX+u+oIR8
AnEhJ9noyVHN0BGqUah6XHxgE9wCHLoTqm28K5JC/e/Xf3pcdbOi967AzOKi4+5D
R9M57ogha8IQo4fkxt5lhwqNggDks7baBy9OpSZ/aYvk1mAAlHXYEg7/FEunmzwz
IaCr3HqCsLVXp9AmPAUR7se4gyhkkp8mB9/ksyA8HzUgvyO3ZshixY8QkJnknWef
LlN7N5TuEOb30GUt1hPJlHjCaDXcJJYGXBijWxhSR8Jiv4Pcjc6s5ftnZum5RUpk
EWx5DlK5OnnI8buUEbS+rmHdIS/H0O3SYSGJ5MhGrsjaXNhOUhZjlEq5sw2Xagth
WOLIfPhFtyMNVcIsbzeLpnBSlkq5y1HKGaFcmHEJQlkm0B0VKgUeh6EE+ROlIkSD
sAao0s+1ixjP991s1bPDJKLTJHrw0SQej+t4StjzGwxZe0tBXP77njGpERT4X0U7
QMARngemnQ4xk4xSJLtr5f1Zjl1NdJL27OnPAiRjvGILl22ZYMWGRUGlqG9GM96t
+dKpnZybXZ1jCP3VNWbOstASIHzSsUIwe6ero88pld82VmrZtxf69YsImVH7KVBS
ErP3g7TTGOrIFcDQ0ycAB4B6hQNqE7MDBORKiYB9tMH+O5DLfqt5wDZ7IwBA951y
/tnoj3wwQXFWe8bz2XNr4UvP6EOObHH/LfJTxLhrPXMvXPqccYo6zjhR32V6q72Z
GtBjk2CE6rhcKWlufsHLDvjqheNlZVfL/PuXF/r9RZtR/XAErPpCnydbfRtznkMO
QQU2CcFW5O+o9Yh7fka20iXJ0EHAUFKvbuIamRf1mwXsOHUBCgaJiZDtQs3ycJFK
SCZ1accjgwmRU1AgBGSLBZF8xkBV7JSHOlNaXC9zCpiAhOsXpzlYuBnoPvpbBNHj
5/Gh7xEQJnMMuKMFDRTPBqjm9BlbIw5RWvZexaEwDY3MBv8507lPsSx/H9uXghhC
CjkKsglUZOIZp3w9zLnt5nONfp3eUhLqaJeCXUwboscOR4rRKCBrLBj9MA5ZaD27
lD1VSyVabnZfpP5OL+iFHnsGJyd5oHVkk3EGHelt8d6OVC1suz0C5n7+dfEbPHpf
3z9phx49imqiNecmhv7L+Xfnt1ufuUY2zD/r4udzimpYnoTXBIxE6H1+OE9xH5oP
nknRC7mCMnYaq2lU4uRxJmoLc/K6E9HWPzPt+HMyYZveKuHuX6iIgsqICmuXyJUu
UQWQsjHqr3xm1xsIUaDTxQBvvWNECbWa0lJAJN90/YxdGT1GvvSl75SEmjfk4WtX
1vCxUa2hoc4/I9kP0KlIGhoZrtnKwRvlquBi9/FY4zfCEZTzI/NFfCMFIPxPDeEt
CwRpSGQ0rBZB5kwkZf8J3SbrWU6+LXFhTY2Vq7YkFt/Cn6LIpuTn+eGYoY8nSvU9
jdOz5vyAZ7lQ+6tZm3SaU8/zNjM7EsPkjScrdHRqWTL12TpaAYxkpsXiw/FLu6g9
x/7o9E+z4e09ZqS60QQIXgIho068WaGlCtajraF4tHZ3eNKOOrIPgZ3k3EZ343ew
r4KqB9VLGhrcpFMYWNXwSinjr90PY+AeoptkEXNG+zl51LbTlSOICaShPLo7Ycbz
zilRWnGIGY0CjCcMaAWvDH71pJ8fjhrd+sX2kU+D/7Lh1vigfMgU++/fOqIwAPdA
b6TOExV1gxBaMzm/BOugHlj1s4JqCxusDB1lIMtmGJ8OgLab4/G6yRXfDI9gEnm2
iQZszdWNGxQ/3K1IcZA3bcwihHaQCEnn7BHuB1V+GATcX3Hacwo849YZ1A1/qkv2
NfSobKwS8jBThWMnGNXePUPJRWhDkyQJb8h89C4omt9DDk1g2G+Ae+7e4JxwAi6y
cddSjmpz4G6Nb9iCkSY0YMWMTx3ewj03AlaVU+r9IWXHUGcc1J6tMqJw/JN+2jpV
RPlppVN0zjepEGiF4f/ofaDvGvQb5v/i2PjUg7pgpPnjsrE7vvIGovc/0oZV1nvZ
5XAg8RpJoA6SrTqS1/a/V+Nal1B5hRC6lu57oACfW1nBt24S55AFE0SPNX/0i7xk
ztTgymio5VsqAZCvoEj4meLdPODOayesGiiR1bBkUankhVI42ke6HeG1a4xLKY2p
0vl0Dvg0fLZU1mGRR9wthNYr5GH5rc5O9u8Knpo16iHPxcyS8pRSl/S6S1KR09Qt
HQyJehD7pT1IdBd1Q9uBIW99soyVRpXKHcN1M9t92WPzweVkYBZdqsYzNnHo+B3C
KbTkDixV+o0hm8KCLTt3ZvljZ60juf3eOJP4VKq4c/cAlLkYcH9l4XDTHtTCU0Ah
YV8OQfL4qFgxWUrQz09N8wUanRmCu2K4eLGROPrvlYCr3KOG285YUDUuHmwNqsbn
Pid2aPWrBc/ydf+gkWE8RXBJw3hKDcORxa+fWtwCLoiNFCS52ULQbQoty2wQQSAZ
uOu7W+WULUr/8Hh7gbPhJQEarrnc4qn1i9gO0Mx93NWC8X+C5iuFycByzwlDHNgq
OtIlh6Vuf995K/O88qus1vVgPoQGrg01HRD/rD+8oXsOfVMVxD7rzg5tPyR58B0j
7XMQ5A0S/IsbRh3ULKPRHIqjSW10/M/i6moZY3GUg6XqjPqKLf6V1m8Vh/V4J2jo
6jMT8uG1gaKGu94AO1KNPjZGV80D+OCkYZ52FQfTtb7IJh0tojDjhKRJE8khfx1u
BfFbkPwPgofS1x0waxhEOA/N5HNC3ov21WTjW5mOPFhF1M8qWkYPvt9t9rEcSXZX
/Xa5piBa5/pZDStuxR8XrTrQp51KPu6Plf+mLIinwe9SKy4IrvJ6hX0qkILZMCZp
SD64Z/6KjUsEzvAxmT5ApzTHAP52toVOnq/PtwpcnbMCdYDUtATA5qjtRmcVeHOm
4So4183pRyrAYE6+GZ8M3989zUlJklSiOKoaze0vGKYK5LbPbY4SN796Jtk+Ic70
plWVMVoM+wvxh/HDPogf/7e1x0rKKT1JTVOcRoh63VcLMH8Der1uBIqNZzhUFDk9
rSniYZwsSwBeNfkDvhWprvwzonTYS3z/buqOaQhfRFljPVVKi5hOqOHAEnT6IrMF
QgsPyOPnNqoC+EZXzCA3B0H2s6ZasQQ4VBWXpTbRZvwVvnGeYyCHy/IRDizR2WmA
jaDKBEqfp307arxWNhNxPVHk/2EUCjLtU9avoUMxBsAHbIpFMmZS5r57AFAfZ7aw
tOJZXfN0f15JIAEnHM+fGeM/9ylFZjgjW5noQsNOQ6liJmzqHOur+Aevve4i+Qxf
tvtak3nEmbKYD5aO7qn7abNFeqYxfCOUeP5xIvf4Ja1olqpju1Hx6JFWGqsajJAL
6wjuu7QUhZSbBPd2QuAElfGElUtrNjFfReRxyny46kts3Nx7nna9PvfvGjaNIot3
v4yhBsf2j7aD78oeYc6mXFxdMPCrDtC5wAK0l0r9GcUpr+s1yUN/FrlDGt62H1OY
BiKfaifCyLFemu2zUb74rAJObapRExRc0KtcYu6U0/7yJr3Nusppv98LAKpN5RBi
QOZyoYxLrbiDBJFLWsxf+NezsvkIX8tjk4oNIHkljlYP612hf7oso2sjHmwCIh40
tiOZIy0TplTyvjCMw7wHkbWi8TZXJjOytfqCmzK28N34MudBJtf5ET/cSB1NZf72
sZqb1lOUIJTgOo4RdsEcgy/Uaecu0wcUGdi8BiDC/p0vxGzgA1Hur8ovfjZyyeLQ
AUWF3m0KPnA9zl2tzgvIbPR68pXgFnG6unrC6mLs58CTg/8r8Q3Dp5+EoE4PoX+M
DQG51+pyu5WEmi3F9Uz2Nnf4B54f4NvUdesmLZRAnLK6N/fPDP3PfmFEVvfr745n
XMCiQ0w9RdK6JD0Ekr5heQvQkOdnhOBNJZhYBJJn5nZTFStrz8+jLnRLjyp89XeA
g2S4CJ3Z9bZjlKCVZR/Q9Gu24Jd85eWr1Vh4tuMqYOhfptJw6vZQvBe7FKmkcmIe
70R5d8Q++LcrZPyZRx5Y98YMd2+6CJNr7qyv6Qv6zwHPFhh6FnUoTkIqSRdeHT3g
3Kr0b7NfwMLoZL2jG5YztoQ0ZlCsmazP5cUniR5mEwdio/tnmFTDs9uM92Zl750D
sv3sQ/JxU7NML2FNMjJLNFAfyCMXP6Ysg+OT1eYkBti/h+UuQNzvNuUCuMlj9rLW
bLDzMQqZOYW3yEj0BzQbBclpfv7oNL+nYpt8yIKXbrDnHHvgwn/9va8UZ6Om9MU+
WsC/UpaaoegSmIaTpm6YqHQdNhcVnYsU7vjMbrOH3cpNlekl2NwK4W4xiBET1iPh
VsngoiSBw8Sn6EzwXS0IZsTfJ/dDqJ+4braWjmsODrFM2AzYKz+6QnOcWBCYBKsS
yav6ZeIrc59d+/DNbyb5T7X7J0n7XBEcOjtksRx9Swx5gQ/XO7lqFdx7+LQ9ll4n
1xpaUPmO6HTzzJFolBpo4WAgv9krzvySO5puIs8sC3AF2+lns/2CKs2k9Q84hRbc
HpYgn6WR/OActCiq2VVrLtaT9u6b+/nbPBLRB5p0rhov6B0EkwIWQntGPwqm4NsK
BuPCqBzcuz422/PgQktLh3KKnzEdQVSiMBU6IbD2iug/Om4cZwvIX8dIe3PgtEXz
EZaPMvXuFuse5q8eFkppXbaMQ4TFcNeorIonlU4/WnGcJw7aW8IVeSXuKHHWj6i8
JgUFfHulMFJwnfft8JAWs2x/gQcn1U7oI1Z47c65MPoX2NTANpc1+GP62ij6KoXa
En1bj1uZtkGqQSMfZ1aYes63L5e/tbKrdEx9gYY3ltYNTiO+nnt0DUvq6+Ant4yU
poy+/SfOfsgk/btROxUQek1Oxvhje03SyM61MAXdq8rpJ0sKgUcEBDBZEDlqLcPz
o500p3bU8lVPQLf5earfOjE33FESlcma1CSqAy3VTxonrfeI1dbv4CNaQJ1Chxw/
dZQuExrCQkStuJKtbsGZwpz0QQSy+/3K3nRv7GEVz3DAxffbw6NyIIhBfcP/x3/L
RRP7GD04NAi6vgNzzpSruXSBsP98YiqAAxmYu2uRo5Xb/EaS+1MgD1P5THNJhIlr
iXVgn0dGiW5RuuufsnXpzg8XxIMk0FeFZ2Ka97Fsi0HGaaaLCjqLVYTtEBXsIf1e
5nA6vrNxGKZ0jansayriU3t2Wf/VU4QGcDdolzis9qMnMibJA15s8bn95e6lv3D5
2Qjcht+ElRS7PlS6L3a8CVx6Sr8r47g/IZTZkZ+goqKljWhbIkPKLGm6DMK4/luT
TkPtw2FZ9Oqm3BkPgCRXpZu+szWEUCjnHgQ3yv/pCav7d5ALPEa0dcb37zzirf96
7tQ7GLcpiqOEwMsuXyMv7NaFGzlqV4C+bTUcMX0kyPoSlylPMgc5fM8jHwkVZDfx
mtSYXQ99ejGbNFHzKRuuNp8yGdGiDBtAYdZhIPCg7zZlNqq3dSe8nA7Odx0jX1ZZ
djzxgM7vDezML8/RnwzfQ5m06BDAAUEdPitOuIJOg+HNADiBb0KJON7mZJlkxagR
JoZ5+TTuG4yZxdCVX+/13grR84a8E3gdHUyzqpV7SmCFwlCL/BLhQK0DVF1vOxD6
vyzg1bCwkBwn7f2olzmrGe6WtI9b9gOYzm2n1HIb5ShqekNJ2PIKyAbqUeM5VMCe
6L8prhyiA+QtBUX3lMD0yr6tHa1M6hA7Cab+Ld6H137hIg3mTO/N7x/TsijnKY5w
BqHpzMSj1zRcQXurSIkVh7PG1SkV5YwkKUXS69muXQLdMSs0/ux9/JWtwQjwMzt7
U3iaCic3v4TY7EcqHRe6Azo6/l04Ff3C4USMCmsBW/DmP3E3gIz94iJrMIsRXavL
y8Pv/HRjJZEYjiVwWN+Q5ApQbk08zQ0YH1xfCAF4KyZx5b9n7D1nwdXiaKwEI/BI
gE2FIkJTZhWgmq9G6EtGD5l6tk6EH3Ls0WYLhxNIkcupJBnymBkfVTAzEcevTOdt
/TaHRVOR3l1Q/SYGVcI/kKbpscNe6uingTqG+0Wil2kuGw5MRST6JPS+73Ooh9MQ
xTSHvENul38rwc0N+CJvhbo3b7Q7D61FHGnQJwX/rmJA3a8x72QWm6DJFGIdqGzH
UcWVg3wkAymsWa84hrVZyTcl/bc9x+IRc8TO82akLsgLYqf314hKCc8dgwI89fuE
zXGLhsIh2lmtPp94RE+nxNCBD4ANjC/VH80FX21FvY/R+0f1YaPSDMkhm15dkfn0
3ShWlZhVkByFfpVoyafbiXAdsOzxfw6dv7DpVO0zJ1v/++DWlJXg0LtN4+JmVE24
0j13GdR2el09s6HzoqPgvwSSlFlnpzD0xONt9Au7t7fyiDd3N21zu1X0XsV8FTYZ
9neinsHrpBAhx9giWbH/NlsM6PSiUdu8uSAorYwa4LxXbEhV1uz+3oeLk3uhvqYw
49WIdqK4Oc6woMGDUI1ol3OMnA3VxAngbhiHZSwUiCEHl0rPJLcBJA+py7bXCW9k
IT9ut9TbVperN7OvMQd+SqQOXVb75RYPVUryycw0lJFf6WLgVww8t3Uzenmnd9qu
U5Yz0Uq0E8dgAWowopMDJtnb9DHFNVxg46sDy3RlFahKVEU9AOzl+hIN41A7m7HT
hiKW78elwT1dyETfHvG4WbvQYM8bNNm1Bltf8aYxs8nA8ohLwaj1Rq3iKOK8mJCp
d8vLU75KiUQuuZYwmKOgLhfqeA8Wj5ZLOadapFDPZ/usuevvu5kdQOnM3biQKnMV
wpb54a1GDpKrkVMst/IHK8MTS/6tni70z7lO4oibnx/qVG/vIyzPgoCd690cj1yK
jnN+jE6u51NPhDt87YNCjAGXVtXjZwVLrEioeHMZMg0DkD8MkP7U/WwOV+INOf/j
JQ0swfisH5m8SMWP2wD8x3NfFjUM8Bit9ZI6F9NQODJsB0OmP1Mzy+v4iBHddVz7
DTYkHQ2i5ipThIRHbhCcJ8FduSLvBDWWg1eNBjE2PI0SO+YCtD4DlWvQDvaDXLgr
6aHHIBB49g/9KaGWo/f98AVgwM+pgctwzQOGix3Fj9KCfwfD/YYckC2LZjFve7Kt
MTwQuAEZ956LdScJq/xk1xsTCcz+j4KD2WCl6pAm8Gu2dNmHlyA5xXzYQlKMD6S+
DNPEnqFN5AUGQVowHtgCWMbu2IPHHvFSZBjxrs/JEPDzDAKeBvSTFt4Ku/weZnxT
WvaBZmhCevwVBQP+J14ebtUNV/T9M1Gnifpmwf5d5o8S7W7Gr/TwAnDOdAqvZCDN
BryFt/wfWFORDhvnTI0Tt9w8yp+shHC1uZ5hob6SD0C8IloSweiDJ2NdOz5OimYI
/0btEZWccIynnr1IdNvYwHnxdaUi8TMVKFwoeIfZl3goMKW6P6i705zCZhI1zrr3
/l1YYpXyp8+bsK2Q7L+DiuITgFUQP2c1Ncc3zlrKTJPYBLdQUSQsFMPBc30pYtun
dFojsK057KaZuVNbHlKA6eii4ZnfXFD0XIdquEZik40M/7hTVcPL8P3OMYNVCo+A
lLpsSFDaoD/+892KYOgs2HeHQSgqVol47u3SHEJ+G2R3Pvu1ANZi/RJdDMPZ4zEx
fjuh5Hqky9A3g3oG2v/Hh7gWI5k1PYnWueHVmZx6q/L3C+7D5DzK1kZivkfPqmeS
sQEugDl8uefHu+gWo5zKYq6WPuln92+H7VmQ9fikCb20K1Yh5dnCHoeCytvykz62
QI72a4BYsuoOhR1JnXsP/A342dInRAJBtUHmpyyag7rgIebK2h1KUfSWRQphHiFi
3UMPIC/wBLdC5P4slKC+AKjcvMc+P1o+5Ln6E8YYIptZWSEennOk8+H300tDz2BA
hZmyKydhj5LdOZY1QMQ0p9ritVjbYWMnSJsVZ+E2lD/U5AX35jMKWxvXc4EnxB48
WEXi5iGMc4vvIxmkrMPjHpKHLPPSI6RAFwJoayVtLDq8FGdqv3Hw5Eo+hiEsTYFR
sEovSJRHeIoMZ1FUGFkOQaD0OAhOB8LVBlBVLEl9zw9yVSkYB6ge3FyxRVElKJb4
y8GdR6dnbOl6W3rP7dN6kC8iCovuRd2HA3csczt39lKEavMaziBL3m9WMnSr57dH
SqM5C5UW6KFDQYfETSORUP+vaDSc9ezh8W4lunOQ2rP+Bn1R4m1FbzOxLdzgdbRj
G/7EeDrULGL1JRhwT/mQki2rTwOuruCzXNy1p4bN9fldHQMum1uPHGRI84zERhgj
xxP3nuSIeDRV/Kx4R/mDnYa+PtaU20CPZ6PfXZ8ctplyU/r4Nb8DRLFQyJE61mBX
cgFFvxfPjobQE+Zx+UPF83tDOfTk8ZigwU97WTkG1uIkfDWP4ldzQea6qC+1Wphr
9hHGiT/OG3nXOzy62Ufc2AotC7lxmnZ+CgOpuYAQK/uL0XOcpcdO4HxTR/ZtYFBu
TwaCoAB1AuNpbf/0iyMOO1tY5jJoiXXjENr5vpS+Z/xwMv9BMY9c9SBgFs1rqy1o
d9qP0012lqsNpA0arGv+QM+c5/C3FsGnB+KVYEnxdrOvE7Y1qGI1c8hmb0TM9N8G
JLGgz/avVURACxMZhEqfkKgTf7u4p6S5gG6az/zwgZA6w3dASQtUx4tM6uaZAlQh
mjesIbm9+9RQgbrVQjwbeXfo3hSVMCpaKiGybS1WzJKwggGCwSJSTpHaln6+SAbz
bVv50SWdEDxzFq5/XmHRM5JHttMLtajggt3ihV+uNwzaczjJrxfD9OzVYnJ8C5AQ
mQGQPOp2i6hsibKFMv+XIVd1eEuWQJ4c6RQEziAOgXsDpnUDDOZCkHTZ1cNWR+hF
ox81d9VQjqRbbXoCLje31Yezao4k9wWGmavK2hK9L5sfnudXhuHIjgscCcyE+ETO
mRX4rB0RLwRNHnQwX60t3Y2LKPUEQd3woTOfHLdSU538UfnQpDDOSXaY0tPK+Ckl
36SNIMOoHxHOWNQqYj/+zJ+zRGp54HuJq1YUrJVkWIy5WMpvGmQGY1MTSCOPIRcY
DNIhKFiZEPE+/9OiZAexX8egWbOeFbpoGld9BpJJZNrCoo/JLoXN8c183cz544AZ
d9S0b53+op4j78vd1DpFYMjH/XvQu9mlO74mzt123gKQ9Hn3W7eT/9AAkmxfpMp2
m9kDmjWwlA3CYRsHdOLd8sevzb3W5XyjSljDzMXOMDqCbJ1QsP95KzgUrh+rhg18
I22p4pCw7LeeZkh5OYf0Dppm6E8+JNHFdkvvulo/HjhLIqb+wAyxEXQFMMOCc0Da
kDbnoNo0HXV2kkTSY3WBtE47nFZfXfRQnJN6q4y5hhlbb6awCoJXsT1fOba8kn5w
G5+BRR/oHn9/ZkbwxDJHabPoro1UrB3hIWxT8hDbUMiaHuqBx1ZTVqRrcTh8AZCb
P4fKvrvN6Soebl+B8VL6S/AVKqQD9gb1MkVwflBcc0bEtr0nqYk2u1hkKMuwiNCV
3tO5/MLZ+xXW+fwbCIzFdEayOkJBJmIUAfHDexrBj3BGd9P4C4VJCrhAqaVQ+R9y
jqjZ1U8Vmcuq+6p3SvxP/83F6mmnA2s4VCezOSxKqQq8ZqwkHpCvvk0fV+anPJJB
WOrDX2QII1NkTnmXK/ZcX4bbFQL8feWZLcj//rTNCit6Xn9Y2lwMzOZatbJGvYlh
09F3f6qJ7+78gR4yP2xGkEC5NGOxvzlWQ2oUR0NYUZ6gssQhXaSYfxCva8pbLYcD
bvoZeKr73Tx8sHaSTKoVSzSMhbTY6ul8cVJiRP/icqTVobyuceA9UCsfnDyjsxuO
9tRG1ShEC51OAlH8Zb40nm+BC1dp6MJkL9ACbZb2Jr+6VJA9mRFKWaC5XFQuQmXM
7KlzM4nkCTdggODU9oN2cXzJOppTQzw3wT55xRBcjgGugp57QPRk3FTN3yR2hul0
5Y5hyfqEexmNF8KKCqj1a1HzVozu5oB5Hi57lTGex4niHmCzSVYSfpZ0ufjjMHCT
lZMu1TVOBgNQCAR2R0pZEOZHQKxTcFzruOu7flRABUZArSlswvBUHFk2NZSwTR/M
/oLTZdWeXwT9YbIZSo8ihEiAJWUcElSBEz8CmAgWk7wZUt+wobx2Ek3yeoCS1GPm
M9C4rCWBaHN69xlwnMBlxHrKdQu/VYPoBdfXtbwK+oq+C3svEDIOYLmfIElJoPQh
EYXD4YXh9yilcZyQZo1l0DCyVsus8Tg9gqp0iFFfdc+D5/e649YvEUCI/Y6w3CKq
RKpl1LEtCyihxP6SN0GKqcKzmz40QYm0BSOn6mK7qY9yb7+F6mqapysbufY/UjYF
TxI5qO/FexIK9zvcgQfLNr4dWWADjr8wnxwqx60Pih2DFpYpZ5EtDvFd4ZJrKLDQ
FjPJbeirjeeYDxrgMEEaQOU6Wn+/9og5Xm8liuhp7iJrcDwqCxXUI+glWO1l2vSC
t39yrmzKDM9Oq+tVH1jGPIwZvwwOW7rR0alTXGBQCq9r546K0gZDE0t/6nau4QRS
PGiH6jZoW7nx0pKFVUC1+7wRUqcj4cuFYPTtaoMCSFxY10DBZocIBZAi5eAhRnCn
1lPctcyRI5eAmgbtYO1M25UQjbkkGX6GYNLK/233WViN6rTIWVACToTGr+A9azOt
XeOArfcat9Cbl4+yVMq+11hBmXb+SE9M1kUoR2X+GvhyuKgfgnfIpKtqy1KwQ9Rj
pWZ2Kazheg9hhvMLpvy8mK2vparIs3eo1OnOm1gJ+UxuAgXYUG7i6KVq2Yhmj6aa
VvY6HdgBh29+GF8ysjQZaHYeYqAeeSxR9olAVmEt9H39NDj6og4xBnB5y+y45G+2
fIWiME9/7OYD400Q/FiCs2kzW/JU/TSQeJhrmX8rGX7jNCMHsU7CIQ6/JLn92CM8
6xji4kMkS5snrAhkq1HpB0iS82zZp19yXO6MSdtTuO3Y81oIreHJuFW61PaJ50HG
wpnF3GYKQZxZjJO2LF2SEndaaK5Mh7QIJXGmfHiyEnkifC75U30wQq/ceGCwTMgI
ApCtf1x2T7cRVLTysCCSOjW6tqoIusdm8WzFCD0p98VQvG+H8iHhtljwNaL9h5pd
alVytELg94TvfyQu+m0cGswPbT+jS5XYN4OqLqLiul6O+/+bhfKCaczEDU/Q87aS
UjAIUoLnbJJMcqwjNfLusM6ZSlB2KP7KTw3987ntZxSQcvt9qz3dQ76mgR3shc5T
i3B2jwOykAHyikdKhwR4s71yQTXQpl/4+lX9sS33q7eB2rutrhvQmxseACC10rzX
sf0s9nkZ0XiVUtwL698VcHVu6TIGFqwaU8rsx22hsOO+NW+vyfFuP4E2dhqycawJ
cn1UETMY7Z74fg7CaCz+jNcTGwNh6Q9S7UJAn8AT4cBFfmGEUGAyzTjxkvh1zjYs
XpPJs7TN6vyGJlmfA7aBFwYqY+/u8+bH22/Ggdr/R1SzccELgqD3w5HQKjI7nK7m
47pWaFb1AJA/VwHz6EnevgaQPt65ABVCaWvpTvNIJ2a4t1OgdIPXzJChxNBQP5ZD
MwK5sXPcoNkjpxqWL+/HOg7DmpUQLlckjjGDeAOMqNtG5Rti6rwCfmc7+f7oid0i
pBhuVoH1ldCOh5eXOsrm/EWnO9yct+/oaShPXz1Vo2OXheevigLJkba/9gWDeW4d
0SIiLAxlJN8fV00Cw8/Ji8ZvCgp3dlK5JYtn1QZuQklt9ZSWJVh9oPeCVjG+ZXIb
S7R/7kcmkE03WmcXdfPXlp2CQzqYJJzOuf+5kOZ3gu6Fvc1ttHQYnae6RWul9j9/
pBDXv7Av4reFX3sIxnViWWMTmGYotTbDqwWlknyOlFFQtiYhTNixWNTmhqqCc55U
yrf7ZTqJ3ogQVIk+BumBkcRBZ/ukYalKm4mNbH2dfKSqOrpC5OClFSEe7//b0c6u
fapkRjeJexetsHLCQKrDeJdLvRnjm1lACaOpc7QSG8xpA1jvoSued3V6QricdM0R
KExCpa2zK0u/zlJ6ei4NzYZwo4IjVMwJ/AuV7e2O7WgeMerbGnc6DX7SkqsSv81B
kdEmjA32R+IfrUJ8lYzHo5HXrofhsI4B3pafst4wyROrbVi4kmj8FFbC/1SrndkI
IlnTshqH2zOsQ2xOddYCyco0gycO5o6Eu1qW/8X2JwBVwCwByzTMJlLu6/jtATl6
DYhyLYJdQR3ucGQ0FV11f68MmrsfReA9usCFaVotezcVaAHZ/zsO3BaftGHvcV9W
M/ANrmFpIUSxtp0//urwdyegVVa82hI5SGV90G8k1Z986pCefGgNhGl1wSv7pJgQ
cIK4FD4ilg8q8qwWeA3Xtk9V/hJgJiS2VTICdRSq6XLB/F/uCa/cG3G/BFptegmf
IpgAc4SVb4fGZJlZPW3KfnSHE51TT60tJ2inxlkgyeMfVdOEqeDC3MnO6E8F2DLD
ZD78+lUNQi0OXpfNjD6F0M/AYMJ6Jn67rB4eliOMK/YnALrBgJG/M14hSnB3ahGc
sufW1k1OgaedtkdF5fBk7vSEG01+SrUbZrd4dIVjpU2Lpw3ypsfGgUR7aSDgnkgv
20/9JP2UIGUaicyOoLql5U7B/x8+omjNDDhOVW894gvpDvzFs8gEgmMRLnhchDex
kS6QGrTPAIQ+Qv/tr0qyz1mJUG1nz3BsMVazHT/L3tOA+Cf01Lvg4Y8AndIyooo0
7dOXhkfyzROM/tH+tTRDBote0VZnD3MUZvjDzUMVkpCRxmc8Gxcoc3ABuj9/g4Lt
EaE9MrmTq+lwL6rgx+TXhBlngC7khcH8deJXZGFA38inQQsaOY+uUpv55mkcPotg
jyPvH4hwTyEAUQg4WK4k1pzmsOcom6uKYDcvOVPP70O6qlRFQqmnYQjvY+WiZYm2
ky3TFhtshGtYcnCddKa8NCYSnS+HIB51+HRPmyl/dNmW8GQu+NAqDkyytVyvrEqd
nzuV6NiRfTMWi14io/rUr1Y5jrTWloilCLkSQHPgwzEBztuscmlN4fq6fEfnA2d6
++W5OBHfhZC0rFxnAJyzZnkAlKVUzmuNDFsjry00A2Kf3iim+DV+Y1e7zYcDTD45
loE2VFoRrrXPAiMypR4geYD8laaXEBF9kwCMInY1uz0unaOrZKKaojGqovdqo8EV
S9S6CDWwQI1joYEwRa3y3d7olP6BbB9PaJY+9HhEjS3FYzdwPCEqsdaqk6R8hUOe
TUTRgP3bGNlb2BH8FX/MyB7FjCDN+nb2WS7gecDm6pjnekwjRqLPQ5A91dNYuChE
aNDDctXjf3bAmPlcDw75lZ/dKZ1VV2+TccmCoC08AaPW7kiYN9tdnkEnztsp1HLI
3r+sm4eZlUke+EMYtd8+WXOeZCqi/9+NkXGULhfo2Lo2ZMU7708F/fVrP6NLXJYN
BUmpnUcUDvWJgJMLaV7UC2S7/gkFpKDmUXHQyue6J3ZcdbkumIJgCnASluIhWgC6
ZcUkxwx53EBbCRI/kBUEbDv6k3fd35q4EPIV3REkouhuNKSrLkafIt/ZU/vwPQnN
fHUxRP0o+sudxTOTyemKmfosoCydPmMoQS9btW58IBRV53uhnIPI7s7TCrwMoBJ3
/ElbbxfXKGv/TT31Nt20BYm+Z13kdsOP62azZBm9lgHs72zLmFLL9/KYV4y/JgXN
QqpotBaknJHh10RuLEyErzVZK1CMKqruL+RzsQgcc2oqDu9ZzdLiHUgG9IJ0tfvo
XtfBpJzxW1/gObALaOPmzYVeCpPe0snT9niyI6Q3GCZ88xj8hmq3yKJjvQyo6PKQ
pRj85FSB01elnTlEqWyU6sssK2Jwt1QlmgSeWBo9Q5Stcbdwnr6wkPLDvIkrV9Gu
YWilchMrz5znqnSQXyXFsgLZPjEhMHL1lAl/X0yDMLJfdZXVeUsznWt2bYmGGHWY
pfZmf/aASBhmfA79oP2MyYlnth3uW3TUhgqbA07kksn/lcgLEfuVKeg2H95v+wUX
JekFstzkkQWoJJ8mPhPm8xYZyBX80dO8VshIwfrBTnQ8CFyvfZXCKtah3MD9kHPI
5GOVLBX8CH/7xEkuyO1JxPOVS4tT/tH+cAJfUWg+V1jEeDrqxzXXEXl0Le5Zilz0
Ue0kqi312VCSQbN8VEUpZe+9n5q+tak6zgC1yDyEev6sDUq1+ohu4f9Q6qcU7kS0
KgE7iFLrGzBNaO+0TPyLjLXF13G4+8PbgYWTAqBxvCa36cSwJmHRju+dBgGMU3vw
I0M3M1YdRmDKKE1M0qyitBbxisis1eMOcUc5ZwW5+NikIW6tlHHtAur7eMXkNtqt
T+yuJC9zCnefrNvy4tBakAcbSqm1h6GJLIxti2Y15oLFAePmX/94yiDOp5PGzqn8
bCz3/HV/AFpMEop72m2uQyKiIvC+G2wm3FNVngg3UE95IBoCZueWYPSeuQMKYJV2
0bkZQpinTTYKUqLGcebf6vzrIbjMCMNdK/rBskpRxi+FnQ5i+Di/PAFWODQR2C2v
Vti3GI0MmYLa9vY6D0XkLAiHP60ZP6gyepC0y3Gr9zU8rQ32++RVI8qeVDRDmwgc
5ieFmu173vpXyPZ8Xnh0MPkng7LaVM67GUHNrUPvggKS9JKDaJUfCyqsNhDX35xz
P0iQ3MX7FMt/rNOuqNAKZO0u+i1MK9U8kxJoAu3lReVtNKSrhzyee5IV0oJOsowI
CdfRTmyj4V3iCRba33tZGSDZzVwE+EqX2owmVUEsLKt5l2q4qikU33QRDdkdnjW+
ptnEg0WaJRwOB+xEGKN8XsNdm3MoecoQ3oHSK8J2JStiXfPgvEG6AHhBpCOhuRE6
rxGRGjJZcau+YFeXmsVf79emGvR3XOwpbLNYL/PCtmUgyDDQVYvw59NvTl6cR+kH
ou6/kVC6E12IEgzT1ewe2jZ9JyzqAWfcXzVfnZNKd8tJamYaU12MeuXjkckEKDnb
L2rzWr7JZvcEEvx2HHEHBHR5m0+mioK1LGZdlXgEwHs+iBZuzP+hQ/mWGYqcMvv1
ELqw527lw/VBYVKvuofWgBeM1ZjWSKAcD6ZpSw5uCRJceJQUhNUwbH4KwjI9C+vW
007grZuz1jIlr3N9N8CgioutSOT9LNxJ05RzqMnuMNF5fwMZtpwRPctPOneC97rw
QUc38bHIr2vtC1zl5Bkq5XHRcv21ZyOCPsXVRqICNtm/QtP1+T539f2Z2b9LrSzk
jbfjq0WZylsDdPUkkK2NvMp4t0bY9G9wu43YiriN3xd11zrEqfFH46nWagski/oC
aTEu9uwrXI1msvN/Md5AGu426cAItCR6HNRaIwi9yWRHey+FVPivuplBktAGGn05
RqyKA+X8RygBs5x2u4mOx3luunZXianTqyS5MuHHEXp9z6Y9N6clzh5uCjGKTCUR
vaA+qhIcDxOWxGLXo/NCcaO0B35fm9xIX5rVjxoeh2CTI+1ssgAhosMw0YCWpIj9
o0FJVL16v82E4ZUpgsz7NUlap8pRZqSU2rdi8fw64oMZKyWXl7C//hjafTQayIQU
uknbZq+lBqEwVG1FYhnj3RVcWIZbnG9AJLP1KnKaha7nHTH5Z6cGQhVm82xt8T4D
La+Q7JRryXWggoGz/tk7WR2vBkdQWnaWqiyTkxSdUJoSf11Drto5W4C+xCQQkzBN
CppXmHqKZDvSRh5A94t/HXHMAtMAxKddarOHGIkbHFwDowqCft1WkIF60YVzgtwl
dV3GMSSLBpgyvkllVqB3EorE2/J9scvg1BsJrdPqr6Lt8YHixnW3hXBHQmI+2cD8
i3iIlYlKmEkozmLEls5RcAXJ1Yc6KLNu39usWgW5Is8sQcMm9lPdcMxB80v4Yk9q
SmDOcT5aq+LdZlbuQbK0OfwU+0722xA3mk7AxlWiBJKDU4E6xLztp4qS7hwZwBN5
KusOUy6qAGVc16AVsQxx6/TyCU9U0k6Tex3nnBOoAuivdKajAy7fO3ypBfuLoR0P
Yz6BbazptcZeED1MJiUyONaClzRbYjyWe/UFHNA3r1MS+2HWIpo1285MZ+m4MQwg
Dvim7A/xgo/25j/WRGskpXyF20NayAWlIrDWtNr0WxjspUznaYnLAAoN/gP6kuZz
RsgBkhvVbtR9xc5JTKT2lcZ/K5RZvEGmwjieAdpF5ez0NHZRuLphTbvTHz0laHUV
kQ7aWK3wYdx1phGLu6KZ3sj2oTC9hhhInfM/UrQ/YoDU0xdwq/oIx6WH8jx3ugGJ
QACJx9OIItF19pt85wj/wSXGdjiZb1FS4HZSTqR5K3oDkrm7uaVJCHvhs/TU3xrU
OlXHn7S8inTBYqCgWRog07/qvLApVAH9l8Y8SFxuT/XwIMPVxQCW9FAOjGf2AfLg
noOh5SQjpVDf95t0+p2cN/oNFBNfxl/dTwMOrGsv6NUNtsX1AJMGo3csOyG6uofe
Y3CoGbmJjBrvAj5hJeYlRvsZsOzl+PEPg2Aco4+6hdOirX5gF1X2DaI1wvKNPemS
Dm6XmwsAjRZdza8yf2ozvYN3Lmg33Qr4otJEe/EKV7Lv3r25mjQ8FoY3FahDDHGr
nYBEk2ejGw++B/LVjJCg9yUO+eszU14vM+lZClXpkBE2oq5qFVD2c/L+lkv0zaww
uqRijWheZxxCREVr2uqq957fP30gwAu36oC90VG2GRNDQWMtg9xbCBCYu8L0Ixmz
uKoUbpMMWpOIw12Ul6E0n0z5cbm7RqDZu0jUX0Ro2ZNKd5wrudUWR97JzBnlzYzE
Gq23Iik3HPVDz4Ox88CKAaaDcpmZufMSOiOXRX5IlEjOg5AwFTTXXLQFZ0z2I6eo
lnMR+PgJUjrusYHi0gDDtMx9yvMfZINc/4ZJjM6N74TDYdI3mZdiZpYx3dAVkHhT
3wOsCebH2Tu4bTF/s7Jo2PV2J1MI8jiBC7tK5ZOEBIPvxrOnqx7by5pAObHV8B/c
y0WmrnTYbo38zcUD2OtlTnBXcBtGxFF/CYTHzpnBZzdoGARcWdsSnHFo1nqGsEPT
adiYC8lcKey08tJYOo1tdt5rHbfafCPj9qrVA622y/76gJgcVGTyHSXIxeryUW97
0rSKasV+AMw5mODHhc0cmUM08J1ar7Zr8DDK3J0VTK6YKMCeUEzTsJyPzau5BkxV
tYpb5UpuCSQQp6zRQafrH5o07STQlVu8LZHfI4IuK0MUoZuK1T9K8w/jn0Gjb9f7
hPkrhJH9hreu9NkSfVnB0snIIRUdI1sH/Q8MMplSZcFelx5m5X2ftqoJ8l+gy3gj
aFwHaUsqE9SnyoazO/vqZtCcJ6mCRQ74icBkuA42KzP50arVi313ibdiSTZ5ADv0
tec5iH7OPzd8sYBoO/m8qR5inh3ahF/EW+gZM6STidbJkpkjytMqRYRCswsxVy3P
cjH2WHFW07n5UMvIuEiSpHymW6QWcEScV7zQouz0foV0kQU/VTidityp5NPXSi1W
4p/ULvpXJOt9SorGz0zca8FS1MaPw4fxf6tib7Z0FyT2tIjZyTv4YQFD6glm1l6g
ipCPAwxvcQnclbD2jys7aGyEkaoGQLwTB6odrGlJS/sqhOTsTAhpT53cfnxZfzjj
5Ge+WxHijUEpNSZAj/v37+pzVIrJtnyDb47Ul1YtSoOx830E1Sq8afwRWRUC4mmH
WB68Qkv4DmtarJHurNqKfP1hvVP9IJZ3ctzIZfuKEcQ+dyPjPp4zKOPIXFOuNjC9
+gCbaY7V9c0FJqSK92n1g+r6NX+FV2MxdoBmRINk5XQC3cY2vTi9Ddw/mgvu7o3i
ci0h44k0xj/fEsYSoR6HY93G4AHwXjMnh8zbfdQyMR8r9r1Y/djIqKCPYYHaU+jP
uZIg4YG4zkcbKG7pexDJsA7BLPqIfV4yezjq4oKyz/KAtNeXLu7Nn7g+p8Frb43C
LfCTRTy4DCsnd5xen4jM+2oQxwJHchK6yor37G0ZB3VA1P2OYenJYXeU0JkkujyU
dECnSX4Ld0omlD0A7B+hWImZeS5eeS+ZfV9CHtX7rLXA+SuKkR6LI1TZOw1/QI/N
/vBdiMlpczTORxsseE1VoD4HRaGgksSAIz5t95szLSQiRM2PH7LGTgtaBX6Olzvc
7cYcuxKLi15gEUM2/zmiRNJOyDg39p6G6PusjJrd2PefQykn57b8/lEJ7aMsDpgo
ZEXfJFgHQQPSVNDpLXg2OoykB5EIFF+P7tWYslkmGNtwxTOtdjjHcq3pAbZ4YQ+9
pNpT1XMTAEYbQjkYnzBXVEaZ/39Uta8/hHv4SevGv2p09dTnIO8yM+1A4ql6Oj74
Rgvx9jsv0XJNIdIIGZCcK1dAAhYbqPijt8VEZFWF2OKEDPjsBDe1JxacGllz9eMO
PL/pEZ6RBUp5WVO0fqD+XTu8/aY9B/DYs5jmjTFZj/YNXVkgqeJ6XtbhXtfGxM0g
sY0F2LUksbHOHWk1UIBgd4RtxyjQAcdSjFkR9q7rd/P+6ET6xDZyZd9ZQ1L14hHV
5Wsq01CCdwHAojeGkQynljgjwK+G+C9nQQ8UVGW2qz6ivT5qMst3pdVhahN/WWwE
yXiybbEhlFPVB3eCl6l0uWTm0RUO+mo25eEJ3+RBdbBOaHjTzpL/6D1COzhefvXZ
mr5m2FQPoIZlWo6itHC/TtTjsGzge87sdJHiKme4adTUQnK0LbFJ8W4JcaMWX2OG
ikHVLWhj2whdQeZJlrkMpjvWj3PDxFzrz8h/RK2NB/At+/Mc8bvwG7Fk1Z2FQV6v
XVzsu4m2TYhqFXwuGGvS6E6N4BelSczwmXfo80xjS7+/sjC5dDGbTgIZRF+SZIAg
rJNDjZ06uf9Ln+hPBtYaPm6wnXQGp6e3COTncuzY/uKNa7+DSUUkMTXp/TbAMQMt
geAQUATJfOxtpsY1TVSTtLbh7UNDOTCDk2lBk+UH6k2Elgt8MDDFTYDHyIeqkAO8
1WTO9kv/YQATj2nSPABsELPkjTLOhgjvdsGc++1kv0dyvXiay9Rj/SVW1PXcwf76
ZC87PpoHmv2gHahoppwYs6wAJ3g7PYdu1GCW3hGIbtSn2BcWl/GKYFlyz9pN3Ien
WpTy5ZjU92DUe/La1Zpg0ux8kNavC1HeJwalW5wVc5ir8XUfrcUn380kEvVkHBJc
nsXX2Eif2VWYrJx9ymvc58F3XrXXvSfUFdek4Du1vEQpQjmEIrI0QMu2UT5yS0QI
xq2JLo8lWSMiF36Ip92VC6/8RrKVCiufzWrzYQREuuVj3kZvZ4F3lNYmkLDZqvH0
SSx2BGD+uSWY3DakONdQFVSsY1oUHtX/cnJj6cViwwYfzHIx2vdtc6QJ5uwNVuo0
6VcfoEJYlCFtZYBjbLYyUPiIUzrr+eJ56xlydkVhY1e5HXR2GdU2+wvEGOSPFl7L
gT/w25O2OObdRUd30OIDlD3CHChR5DXeF7rRqRaka4g0kkUrVXrN5K+IopbUcvbu
4iuB5MC4yRBqjq+aj02gpgdZ0ezSr2bWCy4I9q2EDtSnGQN165zLkj4qmCYxrzYB
xhKlm10A2QIVFOqU6ZAfcQIdfmB+XDBGeY7//SPG/WGnyRltUd+3Be1kDgP8faZT
IUlb8d0R4fVOMXQhS2sBaga3QUC4Qdqxdf6WgeMrSpefZF4kinmass4IRY39nGnG
UFVlBtDxwSEpYw/Dp2oyfn7TFi/TFwVgs+Z3+DeOTSjB+bKPqYTOZ/kcIPU6FQHD
VetEP+5qgA8P+MjoShHpPDgtWSSa082qoEmM73b/ZrL6av1paySMH/+BrpqhK2Te
j1EN8OGjmQnI+kp/w5awZ8amUjr0ev79HvcNXMMe2zIzvJ5XWHqJQIeVNHn24g9S
HmgLocUFrwQwvzFjZTi6SZrbOujdRxZUkDdfc0B4Y7RRV4EatZLlv++WxeAA1wP9
CAUTjHbQQyA4uMFIens9yhLuulL1ejHCabPE31e3zJ3ktDIKtThN7HZLldP3PQdL
Co4GcnmidvZ2yHgFAPsc6fEZV2V+JgB8byPnhS/i1DKJ95oE2rHs4rSvmvzgtUiw
fX00rtv/8v6o9iMTHAniBqBRNLNYQmctMN+8CdRQJAh5CVzj4MRmuQNXbvh9kWVW
Ei6dFjVwrZZJKkvykj8M9ZT36Icf9Y3JEHLUmRr3isK7c+7Bp0GA6AXPB33ofwW3
JwiS0IjGWoC6FlKWKtAjpn4oh4rh369AlQ8KOKQdElImR3lWOVvZ520uV052QJK4
4zmazAOSq/6TzFwtQBEPbrJaU7X3fvGdWZW3GKwiaie4VMdvN+4OkTq6btF4EPYU
`protect end_protected