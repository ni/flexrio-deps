`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
Cvhbf/y8gI4/e4EDOkqWwz9761gnhfqJEZ2ywaa+NJeVRJ1x56aM+7FSras1/1QY
H7HrqCxEyEsrSW1MrpCP0rKEYz2sW/RZOzGrqGj2FL1Z5lSMdIpZDwJ5Kji3MQGV
DYCJhZacxDv5BCsghcZjeT5YeZ1UeiIed0UPO+XwStg3YRCeOYx8TwEgLHnR1vd9
8c+bVBY+OMolRmXgIVm71un+uaYMykoyU/j9jBTVIZAm5CLougI8ShSGh4rkH3uj
3f3bm7AG0u5Qb8KlnFnoJrm9IRCA3m5yZyxD2n/N97hy//pa98REuRlT+PS+faqm
/fA9O88xHQ67P7c89mR4GADUD/eDBpJ1u/5gXUa+F7+6vOEfXk9Ue9tEzqLV5sPz
GlpJZZwoPNY1EV5kJJi2NdsRWMNCkkyZm93bedUMn9gDKlnH/+k/vI6LPVyjnnER
Hl2E/bHdncPW8fZlMwAhSGwq+zTHQjxigwgXMrcfq2GofAcPeEbndOLdXlH4ae0L
rL6Wh3qC1snATIPgX7xQJUFc5lVxjE6aEewY8VBtaCh/xKOjk2YFlGEDpzGzs4Cx
oDMJ0iiNrC7QSxOQxz0ORrE03iHreUk5QLRIohdglmYV+kIwYa1uvNoGQO3v0QEz
Br2oNWHw3BLp+gKQNNbuhqDtd84A/bFsciX3EwHkzFxlDmFiUpdTT8GYR7eHK2R1
8NfrjRVzlMrnxBq3/MN0o/lgCM3OYA7lFnWCHjB0FFln45VWz3CKz7Hk7IcRQg+H
8sj3k6bLhYnRaFO/O7+ryvAw1qD6ei46jSIR7Qz9q0pT4/oWMhujS0nJf7tfxriy
qlFwjcI8ObUybTSSLcazRJHDOJRz5W7jpVY64JNy5SZEybTXM5H1zWf+KwuzUkQA
ylIFMQqPu3yr7Q9ZJ3W1cBU4dgSF6oe3NVbxNoWDNPdNuKgVLjcpqqFpxc8YXDWO
6DMsTBb/a5o/LGKDuGCXq0T3ZmuyRxXgTgIIESDiZBGkh/2B4JkBhyzsPwtndLCK
El0UaTOnIe0470B9K4z0nTNDCvKQyCxKEZFcUwMVxMqeThx2jQ9q1UH2wYaiRi7L
RuJBLMSEVfT6YFcv/Xlou6xoRWSpg+Q+669DToY0J8lxCtR0sr5h0ApClN5WUmga
fTjOfBPXlIwqM6M84qwqw9THmDPBpWVKNsrzfMy4hphQn9DKGAmnxronaRcEhQAB
6vORVCl+964Tm6OTx59NAEUPNU1ff4cJEh6jXpgrOsOh4F+L8Gw5YQ3Q18JVjos1
pDN19stm8zpuWgd1YzwQysgY5ojTlGblfcwJd25YDjZdaQLSTSm2tFjO3ONSpQKf
JVZ+buWrCixQiseTWWa2kjeipvP0OPEDK7rwxnVi3bnm91bQmv46G7PAUrPl29OH
TuK7mdtGmA/+2hLM4VKEj5oqSe3js+L1n++MUlE7UapmiA9LIyIcTyN2KcCcU8o7
g0RgwEXxGQETvXvF+JVPUQ+2hbEkoDe/QdNy+U44NlrX4j0YwTsDvLsldg8MFKBa
/2CIK2sHAUcqjk1DR0ScLJFiWV0yfq+e1aALcrAX1IA7EPK3l3PDEu9fjoddYnyj
kHbSNztI1uHRjzmqTzlESKhsjy0yWLcU4LKn2awiFGm8RrqzcUIHmbR+QTNs17qo
9uYNU/+c1tI5iTXIywKCYXUbujETSYDw00ZhtqecAp7szVHT5wntAir9xIiji7d6
fON32+Ae0OnpUV+HqyMP75rrgdFDcvNXXusBpxGlMw3hcwy9uE8Ir+XHDSDpo1uy
FYTEA+D3Qa5JaoJqfdSDuVwG+3lpsX8Ummhj8ABhU3ytZ6WUx+dVZERGuetrH+Q+
SiIhlvbqVjMZyR8mTIPCrtd/CFAkL+yL2aolFJUGlaNTsWYqYG2gb1ApfuanCh5u
rldoaXPCKmz0cCXNHn+f+QO1o9oKf7PWPd24h584yta6F0z3gRsD21AnM5+T1b+T
XeFKGB9smOTBNg12ByIQe6LkO4vUfD0/TNB7udIMdKBF/MbOfjaOb5r/e1Qat9Zh
avAEa0Zowqo53KLtBeCBFyqBlQPJfq/lFMji6FgDXxqsD1eqQLyufqhtOnCT8Onw
gXoN2ddtVV+45zYZutySu/4tIuY+PVwGs0I7fG3SuFDKbUgoiO04wCQRlvCN3lXk
iGB9+Q1Y++5WKspv7ap6CJIfuCvYmwuR6ha5ehh34Yry6LI9kJWppsfsBTGLIIfU
8Ry0lw39vQCFjwK0+Fom5Xv6uiDpEeK70g2tb8QFOQQIV9gvQ+rFt5Ct3fIqLUvM
9Xcjxl7bEh+Z1lSVxGkM30eNc9TrD/5at6WRmHhCnVobp7sSTcGW9akv99coASTo
FX1KmjrZ8mKkvE3A/Y+2HCr3z1goxhIw5N1G7YsF5NsHigfQq+ATdXuciOVFu6Qq
oWWLW07xaLBhoWzA2L3pCwERFX0kzLSd78hfHBDBd/dU6HKZXpCi8GpgpIvFhWq5
d9hKMtMG0tkSb6HGMgSG/rSEki3kVxjkzQjb0Ig1BLTCQgbt8R3R86l5ILuN1Or6
zi6IA0jyRHbSD5JM3sOGOTtApf9NqNia5S5h5TI3hD9ggawyEEk2xCRJ9h3Vdr5g
J1MLaWxHVZWHEZCfCkY+omIx4igI10yE2a+5Gkz7aHOCAZvCIw4VLCGAGusgpZ/q
TfETTSJEIE8CIHTopW6+9RS3it3Lg9J3y862esMbcBl3Q+sCKAaHGS4s6IDTZMbX
k0U4211T30/ileWZC+j3fCQOF1cOEzWt3SEBSJZMIcANrWxmie3mR8gJWsiVpxfx
fMOTi/qmu9Cco+PgOZg7rC7mDVLq17MkKlF3oGnyGrKxCiFvIuwXljCnpeS0dktU
TkafkhkEWIUqbiHSdLMtbcrSiUFtNH4yrLGWb2RLrkOgGENhARkjg+Q7Wyf09YEF
zIcsXbwGpuKYZ4td7j3s4h0UYfGAO83NnpEpeX0oai9COMUSwOAJ2McItNMWAG/N
Ad/WjochpFsGVHqH/B6EYtc6T5+OobSnCE4zAXk7VoGVQXAYmvor1La2Ru5Z8GBk
4jkUbJbNAEECCUFyqv8NCLbcUQ6v1jvRv5fSzZUNDB6EMmDn9xf7MF9D1/LRgiZn
DYK7rOstaSOeOe2L9xSn7oenDtuKRjoee1cvDXI8mO3/WOAdQI4qQHoRcZsV1ejG
3vi5Hl6UkybiQMHWq10U1Am0LPxT197siNm041KZKAmm0hXC0ciCY7HIbCH1lxAZ
LA4XxKI4l3AW5AJ/C+LMxUy70QFkBcqqaI0/iJcx2hy1P6xQtNiAMApMaXKRBdUu
00vA4e9JJH8EjOnl3BxgBSxVfzuQG7616jsT3MpvaXp2IjpOjCeM6/7nbNoONR7s
9SRIJhAiCIwVChyocoOkoW8DCp1wl9Uapo3n2mMRALNF8WP93knvSJHEufc6L3Zx
82llazzZdfPiFlSuU+/5wNcXW7DMumIuL67uxJ/WFIXljn4NPsuv896i0oV6jY3l
glnE+2DLJ5oiCeT+HKwBfAn6Y8f6FqRrwglOTgZdW3RCRveWz5sJf1V8U40a6xx6
r3j0tA2KNVrmTQJB20mybw8fpqKT7Hux9LfHGQnquPEscSZKtzAiySvZilGRoVHG
yX1b/cJW2r7wxRTcLl16F5+htO5nhEVlrN/LXvKSNLNmAv+9FD2zGleedfqmbMZi
sxixtsbchT8JfxC6qTsJI4kwXQsIB0eLq0A1Vwe0p2swMQ8jlinHZ9f5ZhVZ52kX
Jf9Ti8sav/QP5gRSoRmMm/BlmnQoCh6Fa25rCkU1yUGCNBWZh9j6uzGcx0iw0cTS
Y5Lr5LorHR7nZGJiG/GnQa2/m5+Vbi731B6VxyWrHhL7mQeb5VdWaoXA2/B/wjSI
sxgwvGKZ0ux4O5DORVpufJzAogwZJXPwDuXRHTYuq7qbvSU3VN1vamzxuNr/PgGf
LOSxsZ68viHYgSHET74G5bW7TmWmdfY7q5Klg+HLL0RHHs2Tmz7Wvp0HSoFkhkxu
HlqPZT09Qc8HKWn/qBTmGL0P/rbJfKRDTPV+RZAaGA6noQOtlOufys2lfp10F/Ec
XMPlM3+4z9TaVqVJ7n795kkFo6kv2fRbMTQFSm2QUUh92rH7RPYmXTdp21bMoxcA
KmKcJodQdYZx906cT9gByh25tcE5rU+lpD9LIn0J1a5yi2d8pT4sCHat3vVWxcl+
gU0D1tG/UzEzN8+5rpD1ftU6Uo/cUfhZfmVc855+0zg+3363dcGjIOWmBRu2qr7L
SboNoi4lNJYudE5emc1ZpG5EmYG1RpqR99gSSxAX5ksp77MSesC9RPyxUkor0Toz
oWRXbyc8uyzNgj3ie0yU9tPNPy4EvUTI9hPybTWEYNqTcjuKFRVpmL8YUzd0beAO
Yk5KG6YJHM0YZSprHkRokdIECazJX4S5rWDu+/7tTmhxcITc7y2YcChAUrCwHJ9O
O2zjNQv84D2fTVDvIpcoyHFnm1dkJNby8gLfTr7wpldGze04Ot4njtwfvFDzXBLw
Rbv+pFjvt9e7hRbQRlgXpjz/HfOJgPR2Drltr8SekENHrVWotFVsNsbrobEh0YhN
hO+M8cUyBF6kjWGDEteIkcjx2vtZMaJOLzPT5LmpvvEGcwlxA4NkOA7j1NnAA/BG
FZfPFLqG/G65oiaYXT0FmFOjXrWT6VQ3nu+iioPkilBF+/feq5z5pvtHOYWeaJiK
wTnn/5FW9KESCcW6hZCi/RpBdyc7woiGA/5kP1VG7ZnXfIniTgHCJiDu4vGv3XSN
2JpBrNBqPM1TrvC/SqujXHIoJ4LkAadlOHaP6Y9EZ7mXCoBn/PGU+moU57ydJ/AP
focRk3Q3a+k8abuUCPk+hV4uFH8JXW/Bgvp664yZRJWZYt02d60uruUF6/UUM1qY
WVFLOzhwDKhGuYDqZPSVsQj9NICqKnR8s+qhugOZ7OxYR49Q4RKPCOQO4aRiVsNQ
UaIGiYC2z1Pk5hGa/ENJXzr4qM4vwGXY/xbZG9ovO/jncxWj3l4eP4ak0AVOSJN/
WxqwXQICCH3kBEacdlhZs0N6kC6CuBoy/ubSA7SWNQqxGv4K9hDwUV4cr7Ujoqj+
5xMZRZIlgT5O3gumF+ro7c1FjP4hzVNzsFcQZFSlwiBtYKehuRpJqY25H/+gBAuY
X07o+FaCNEb27PCSag/Ck1DiSSO/27bRIY+hrtxBbQPpQ+komd4eD/1bEQZABZv6
hBAd6Yd+YQOEZtiYB7ZfLvLfk9u+W+Vo4LKKbyqeffX+3dD1GLBbSkDwzGMI3QQZ
+HDuHW2p3YIpeHI+RNbnUVD0rfl2HUvKSkZGA7gRO0JupaUzmBdX8mPkYjXwIRbK
4gn96sjnB+LDFpCrCSRiMqz8FXl1mMqfSVtNxoYnCDzy7ZW4bNS4gqelfjTqs9pV
Hcy0klh+HeGJEgLU4vT/y+XdMz/fdmlmwugXi0UXwZTQdDkfcit6dgJjwjrIly+J
NR0pw9DutGIEquI4kAY9yvmmaNBWfmLE//7bFglq8mDkHoTpl7C/EIso3A3uAZiR
Qpd2EXwoz2JWJA3h+yzwmyZJpoVHX1JiPWoXuZifurZhoa9qxUbPKrVogj6Du2Zt
maEKHxzBuIjWHS1lkvSSp6hNYUei/YaKLUYCUwNwtL38OmlUlREJPyk7IranIDf6
gQCgPDqHzUFvyUFGRypEmuomtnqYKi6k32ekiRI3K/gqSgaab/z9jBGw9vKzBizz
CsKDEB2AUL4osRzuEqHqPiWUc23+3B/guUmXUc8m1kReouE+LUN9FpzPWjECYXLZ
4xjWiRo3qVYwGFMGIvGRSy7orUIDcQ1p9NkhqzoqWgGfe1/yOm3CB3Ab0hR2u1Fc
cXJKFISI7IvNrYPALp/ju4gj3SIKFHaWCbgTMx8+JDR7obr+hVeRKA5niWlaueDT
TS3fmWWnDHtUmN1K1I6UKpTSWeilNTz1p4IHxS84/V8oYzEKNogXXlHs5EmYzD8a
Li7E1W6CkFekMVZjjOhM4KkmhCPmxDCj2lunIaS1kvI7NGLv+IiUcl2WzkCvR+0u
cVTaLw7Xx7U6KiLgIICRkYvQeQzSf5d1Fwf0C6vUS8GDvrxNpTnO4ySlB9HobPvf
bC083YMS54LxVS7KbAQx7R/j30iePWSo9M6+HrO3ls1T+7uZi3Q6oznvqs/e3iF7
L7NC7Sh9smz15BK5dl7jYYjD14sdibp05v2alC3YDoXQiGVVfU4jiYSc8cjZWG3z
oqhmIUx2oHGttS0m/A0XeJiluif8ufPkE3kXiUJDwxPKfFPzZl7FS6ABKFqEOi/f
f1ji2mqpHlnRK/5k5izdR/PLN6PMcb7aY/mjLMxCcDlS/9UQMtZn4snKWrTMeS4Y
gY9OwptKyIW8UEa0cPmaHKpfExLw7G5dQq6VCDTMQ89f8qhourqXfFDt9UMqhxHe
XtB/pCVa9mt9dyP2tBYkUK0rXKixGxu7YiDbQFk2J4VQNwY1qMrOOGCyt30XZS4i
jg2pToVt3N3lyAhldWAHotZFQpN9UlS169LQpUuHO4zDAT3WJXQMTAplXoniCibg
NSLvaLUrah4mUxEEivP3uTupi0Z2FlRlpefCg3l8b7hkzuB5zK670PHgUO01tT1z
qCa83ljcSOM4zC5Jp6pjF1b5u3Tv6j3/F4f8i8+mts5MzCDX+v3E29S3bJ1zegkT
8OESrAR/c2Hme8nf7WKRfTYq0vpAqwvL11L8k6syb0mrhP+LAByL6wJAa1r2NUOg
xTpV5Ea9K6BYuN7eaSylJxhxxCba36MeoKuvYQ91oZpUz4LRQjDC+X6UOWGKHTXg
ZsSKA3rXw9kotJcY5BjsAfrMhA5Hy28YX5MqmD6lUcDTYDKXVYjvBAMdpKqeA8NA
SuEJo33gf08tjh7Ja0NIdV6xmvrK1dZ4g7Obtp8IRINZdfIbXReWYuJI4+XR87Je
PRTRQvVDNMv0sykH4J8Y5Ad+H1RlgimK0oH6SQnFrngFL3wrijovadlun3Dga19K
niktkJPbj60HOaj7mptcXEy2N6FAVJ0zv1x8nYPs34KgRCd6yi3tmlxBVst6JbMG
LtepA4PolmUcjpj/9MV2kYAADKOiyUZTXii7+OzJdnlI9GoPZlBZ13y1SiOC5sbr
iXzzgKWpUTsg4eFNUoOZIowJ8miju4JUmAWStUMEzNecWNjSQBs7/sQxmCzdIuTw
Dxuj4VbDZhEgGJMawn9p3h/K3q03UaRSceOSod5spjP08wt42IPlAMS7FJzDYCjQ
9mBvL7sQEdRJL4j928zljjpwB4xqC6UwGCQe8Aysy8NOEGIvyPakZzWH67+jXPcW
t44EHG4YcVjfQGBv+bhY0P3bJDIssNibX2OxgFqxSoJIH0mtlJGFNqObc6VCZGU8
XznqHLcc8za7yeKCsE0WL7qlNZ4F0YJUpNs5PinL1kJU5mOutr98gSyjQl3+KD5S
g7dv7NlG2a+o/M/1k+bfweqEF2GCUNwCWzXC81Ms3xMjv11F4Qdkwg8bPqob/9x4
+63Lp9srk+ejU/ex3JYgGHqp6C0Ufhqa/PmqmyjiiyH1ppRgDeDCWniBXkoudl06
+4dlZqTd6T7mDbJosJ5l84yox8/EvwE2/dX8Re0W+slI8gz8llyAcASScFTbDcGO
QVliK6JLCfGSQbnEkRYJGMnS9OHW2OgSHfXWkWMSVrZFbcnrlwZJqSNvCXVwUxAJ
yPucStTfDv5qetQzuXAEsgATMW/8kVdWB3vDfezKd6efk8HHvAuD8AoIol1sJUrZ
bQA9hs2+74gD4TEhoaSQplKIBY5XL+LI6Evvcy0F8NMNEDm12gkptuG5DFn5Kx3t
7vH2aQYzwpNfkbMbxayXU2e8Q31lltDVmfwdYgHWPsorKb2kfMDLpzrPE83l5HzS
5jUs6PUJfHLeP1rlXy5cBqe0/+nPdMfuO8j3fo2h7OP3NwZBZZFNeH0XhCOg8r0x
f/bTBZ3XO1GeNMk1STD6J7jk6Zs8RN/mFtUQ7ePOttm5IPP/T+N9yWPwpEZQJoBn
3AF4eJ9UfECOp9jXqq7VQyHyzXcbsP46DDQJA05vInSYnoGRHBtEgVkA0Dhf7HEo
RJybnRTXgExYT/jKRvLi+BMNovK0FbA74kKyWEVz7hLajw98kfLDfncji4Sogcnw
rRWyhVBvUQ7Z6KmtcHcetPIQQhFw6d8uw7imoEY+Q34dWfM/nMhUe9v6JMso+Jfg
iPqNTRCNJ+Tv7ZjazZa+9OEnv0HkkQvp7lwbsSAGHifjRlgzRUlu+Be/0eqQyp1n
3ThR5VI4O4oIOEiYEocwEBE98kpTr/8l9r9VAUGv7AFUEphN5A/nwmh5QmkSio7+
AbR4AQoO1q2x31yxjfdbpfvNUnwnxr0RdKmTlYuSGsB0h/iMOfPxZHyjICvn9K2d
i9MFuCWG9IUSO/RCwVziCrQviZhSbdSk6SO4+Z39hjfoeCcnc/QRTcVcQ97jfB0s
Fp6ykLoaPk0RznaTHxB0AXUPmae0/W5Zp5CZarS6YzCbP0j8VTkup0Qcs7j/v9sZ
L4yRcJaUtGxk8wTxxOtgN6NCbhLvp5c/g2Aj+GuZ4/MRkaAsqZ5vpLzAY3mIA4NR
TDRDyJBr3t2vw2bnZvNjAjgbo5AqLIUJi6cnEAO9vGTTNv5TTHlFUjwQpm3Ezx9L
PNBPxsk1TMmPaQoMvE4NTJEBbhuGeSi/BamvIrcc1nMLzgzx41Lr3VgQml5lt8mn
Cdm8BOM6t1NxtKS+EzjLsyU9+CErVbn7U3JH1DwuzeQeoyojsoLwIP+AezMU8+cl
GVqW/1CZEWT1YQ63PEwpjZBECjRTA5ADmd1ECEy+KAagJcBNr1qXACT4S2VHp28w
lh/KHpH6IoblJR5IcY6+fYtAOXNNnsELlrp6NaLLvcrJ/DYhv3NNb2m7Lz5amgyw
/o2avHsmlJE7IkLkT+Lzg57+aTPyJ7D5gOgStgj/C7Af3fHKpl3IIrNhKowCd5uR
n25HXBZKbn3NjAkzVcqWraNkUi7strNa6s45QPABxDs7W3y9CJCCv1Xq8tCkzy9b
5S/zJdqTgsRl7f2Wtvl0VmgAIfFVFaBl/XxquZdttbC5kmQvFQiamrNjqgJuPYKP
e9X+E4yg+zwwcXbNt1FnEM4RksWJB4XQWidegDH6lQEGt0+tzRPhv5HAr6fRlEZt
J68Kpwfqb80Xz5VGEoC5nckJrWtlFlaZ/SWgLb2EOP05m4UgXFmOvGpOZdCRjyJz
Y5IoVicIr7xu3fLLWf5Oa8/7WcsUKTfkVEJqp39Q4qsJq3ZWh6nfMWdRl7WMdkYw
tvdYi4MFFZ8CwmjUqqYwz906Cp3MRSYNwY1/SIzkhpgk5CK8LsIDRkrxnUJUNAh5
WqI9RsIa6OMaVvUDvgUkn8uuc8I8CtiZoPQsEhkk68mlweh2Cf5hGb2bHI/BXyJa
h7YOfMURfjh3TvE8sbpq0Vv/OmJUs2I/a6d7AAddAWv68VAzWv6q+7KX4J/taVnA
dtrefOzBWJQRWc5b2la36YEoaHM4wMuAy+J/lYqljNx1qX4xjR5GzVU/1u9T9cNd
0x4a+1S8xZgovBpGxr2MWOuhGvCTP6ClrfeseVyUmra0Mq0hPrA0W/Yu+E6Nad8Z
MO9AzY8CMvdv1vH5mRmoAvX05dEJn2PTxDl2r6XdfoBVo+OUiYm+VJ1Qo3hH1W6z
m+jDLIgRWz24nn/DDMjhIfPUFaTEyoidIlbz5F100brlWIHc2b2LEsPGTPLZ66JP
mGSK1J6nqRuinjvquf4Mi+5fJJJeoP8DEzrnOR89L9+u1kmotLsimEycCA/RwlCV
Z4QpdMCfnMFTCjTYkRg89d2+2gEyeiol8z0MBteVVit64Ehs018rvgWLf91bUf89
9ChbakzwTOpmkcJyNZnRgSnKnB3EXmSzK7d43S9y9YLy7BSxSTDLbM0DRvFNc9rf
xxnVVeaV++Y1pezIwVk9emK+XA5Fd4pGzZFUXKP10wF4g1157L7PyHLOzfDfI3ev
jM2xIGR63GJXyfl+1ZdFNopmaqIMlHc9Yn6ygfpBZSeYdZWhPu/2Ydi81X2eEakg
IhKNv8JvUBCrzDspOWEwXF4YoD1zqOreEeaJbE5QgNV0cFJVaDvW/+EQbzlgldui
hgh8GNl9UdEgCF5+2L4U5SiB+7RX5YeTRzGaL6QKi+c4zBNmeN8Y1ed+ve4KIVAm
YsFYeYpZzJofju0IuH4rKNhWUlXgyYBqan2FqarvfXicNNjBF7SjARAMmDxgUoCn
Ta3vH9Jpcdjoc7oZxwv05i7NiC1KQ4yg/NMFukE7GMiAzu7bOKyYtWT9VrFUEnW7
ihH0Lx40X+swcrE1C7DfO+oaYLkwgugqYD7dDHb5t6zmH6HGbcf0xzCoNS/LbIrA
frE0nnjsT1A1EYtzOvQGHpDgXOWop1r1BAby7zmnOHvKpL9Dy36dXb1aX53CE1hK
3apfehFJgcmd1dFYUrWhVYDtkjzVu93aKpjn8LV+J/71kVSaMvbOac8t0dV/JRY0
Eam2BSfcDbwbtos8L76FY0oEw8SyYhKlQ3nzcnVJUwSgouFXkw5NcmlApkjwmPQg
Ye6M5e6mcY4CDjYvE5HMYREyYmD3366RBLHJArJ4RuL9WBsJ3MuvHTwz80QuwGQc
BZu/mqw5CcbInyerBxFv2XZrDbqng22i1kjeiGcnuEb36S2YGljZDJFxPD7fQ+dD
9hY+djdqKQoyiTGpo919aYszeXLkIFeUo6hJoT5cql3p0RqPOsLdyJwBxUWFSSKQ
Sb0JLrGq/RVuSNS3arPwocyzKAwwN7ErTsYbAQV87FSgHJP6Qxncu/Da4uQqUic0
P/WdbI3z5LzkjsBApycK7li+HN/MeBNZooM7muBkDOc7x/Ec+A/cXA7WHygJWFly
b4YQumUPakozQrYi7fHsauFw/KWDSUbcUkSIcghb/J/yqbeV1bcyXN1AoQMUbTG5
Nnozvu9OmKlB2tvbeh6E34v8YJcQypY3rp6jjI/TYjoWewtq+Thx42G31RdUTJpQ
awPXxWB5ANTgQYFTNCjb30jICoAflD6O4U91no4J2BP/uDWOin9NLQv642amN7p6
aQOhefqUxXUT3rZpk3WGKZXbWgyUgmXI71talSl8hX5IaFvzdJEbGROjtYZm8IBa
VLNY+b2MlQwMX1CqIpP/1c4Yr+wokYWEiT15ZmAJpcEIqtSH0LTbboH7ky4Ue5ri
wIG99CP6wXA1NsmQLHiKedREVqYyfGYsbRTJkMFvlmZrAEMOhHjq4QgZ3oYCmq24
RzXJ3qTITWpCXtMkfq2Mx1vivwzAFFTo0eEhRyYJkzEZVBJDtoob350EnxyZucYq
ZmX2Gh67bOwIjCcTT4CCJwUBx2UckgT9cPcW0ewoUx7AWJ2uKbzGVeja/Tp/k+55
ezdM0HtrRY1D3gEYCAwZpER+AYg49MeL9oGptle2TW2rq6Mc6FIa03oZMh5159vp
us21VkXwse2CXCSOYZ74J+6XOYf2r8F3KiNCc4kfcKkGr/9lq901a6GGOmMZb4/d
ARBfeUO4n8DSAtCFqpHUf4+8ZCsNWP7cxZWBF4WGMI3WYby+7JakUPc6Ugshfjql
Nv21HczTsZ+A03PllE8X1cEryByzH4XTdJDDd2DipIYJpCK/GQg9tcU72Xvs+C5u
yDUTXABQqijSwabujf3BCTx22Il4ourRGe6i+qoe6GhZ1CDhoWTA9hmi6xXT4GaI
jwm2XAcEPtQhK/GkIVCuyBChuUDUzBWoRxU2v+m6TTiSVTkCL+p3YbyUl1IAhaIM
VYqgx5jQplJ6hlgWrmXEuq+OwiyHUIriIYeCjuzp9Ft/ehQcsY2OMda7mNNoD4f6
dlD7AErn2UAMnkzpaaOmSc1GvdXfOfQwG5u+PdJN5ZtV38gjiyxFxvo2WsrXsPC7
pF+v/ca+UeuloCC3tnEMt9Oef7fCp8ca2NX99A0mpCQB9A+hCv+Nyk0VMjanC5Od
8kh1Iav/+d7rcLJ0GSaDqPJJNar5UcWB202D4to5UUTR0Mr9a4XGIohSEYe6qiOc
ghvj0hrxSPhQljeJTzX51W0dwwyvZLqyBW/JHsce9speuU9cAzCFJssijarl7R6P
5VBjmaljSjf9qEEl+byGHeBBhlrJKZ0ZXnOCENgPC0byglpyYfojznAYGbwgRWJd
aiAiXTR0KcVEOkkeC2M1hUpe3O6PtOhjmrW6jeg/BYJd8XQlmKOYndzGZC649N7r
4g2bWS/qFNssldNOD5CN9mUuuG9aEHAjssER6MRzRhiSl7sCKweXePsKklkCUs82
gKkpmjPQzrVcZ14XULAkXlQ8M3NDRhtU/XbsVS1wByq+B2oie0r0cTCHdOJAtovf
KtpeI7/oqp8EAl3SoIPh1N3SDsShKEdiWX/KcJTbQV8+54DMl6JfjcjqkfPDIfAl
fGKyZ4f93ko5mDE3f5Pr1o/kkDNmXwXA36UPjpjbNbjzjuWqJfv7KE8uePqj8bOe
lnpSaAitl6MEz0tRTYH2kQDq0m7/y8+UaMCSWyTg10bSObL67O4HxDELEd0xCHLt
NNNCPfOTHg/Ue1p4J8ODYRiqb5hNYJ3+zRYMuBoK4BNSuJafqw1KCGw4Q07syGom
v2wEt/wiTuAfPK5TA9axstYcqz39KPvG4GT7MK1eRUPGrr/8spyO6BvOeeWKsRj8
No0BoY2noeRt07lDV9/NYGIsw3WcJVcjwssppLGzIBTzKP6j+1AA945NlIysn0cU
rXnmQOjdlVkRAaLIhVCLeAd3juhK3e6qGZo3eSRuANfwrjA6n/BF3HNz+rJDxuDH
05PfjBZCyeC9s5U+TEThREgjYLW8ZBmSxaBd3NGk35rxnBHyu0kSeOiw3TkiwK8O
shOYnCpcFcMsuBmZSdZs6XRY9aYmz7ge/0HDroZrj+do4I45sKqQPnC2AbKb/OWb
aP/BIOr3xzAy0s6ZuUpFg/c74VJDFosp3hSnC9j8PrtWvo5oXNw/hNpSzeOTmLpf
/uI9yjYxDRiTnbas3LVWO23pwNEl+dR0Hk2WIeH0xAqboUwLqdQQeDDHalrpj2V3
rnJAO/qRBEWQOmnAPbjzanWRqmOWooWKBaKUrPAfmtoSafqjJLxAoeqtxg4x1ZWU
2hiifWKkd/6ZOLW6Rr/2tPzVRlBlV6e0mZZSpKAMjslBkK3beNX/sSb85Rj17a0v
sOKhS3xIK4BtimDEjKRHwq8SnoI70UA8391H49Y8wGKoSVZB6F6gcyGFaFv75cAv
K82IrpSd9OlJ0vS5CtBpHWtu0xhldC6+sgCLQ3iYiGojvTKwI1pAvQ99PgrSY3Nt
8wohS2vhc3hC67UPj9mD965V/LDGmdv/IOVqon/ddn/tGgwIYNgylmItJK4Pev/s
6lZGtGeqKryZBs4M8Wu1kkt6cfnOdHkY1A7V9+Uufy0gdKhB6Ys3VBZVdW188y20
Vq7pWAjqITZ8xfNR6IzS4vrkBECOzMOQR+uHz3l3E3UWLX/c/wD8X4P2CTjTvdvZ
vxnm29+HSDdPWIRB/a04JhWX6eeU7kqeh9jG9SffojNgFTC9mzQVNJWONM7zDWwa
yseX7jUPbf2RS6NiKV/XguuMlhJcMU6HgkQq2uHkesoinZc8gA02ws4ccxeI6i/Z
eCkEJnvD8o5ud8XODtmmPMiqYz48qRBGV4YmAlkerpnTGtFXLoPFs9qB+RoWLVjB
d3XyUPOQu117xjx8wqfc8TNAdDcCRl6g9jEUBLJ1yV0nQ2GoTYlaK5aS2QSpgDtu
UPO1hecOm1xUiK92KnFvrcdTxI/74C+JAaDYgd+s/n9W1L7gsCh57aOSGNIAhqa/
ywJ/QSwVjHYrboFY64Nea+rmtlOmVN1VOje5ceSuONnuawjHAUpH9EX5yl49zma1
bse/PWTmrUB9skiCZ/iwSls4RWH+bQ6hYxjYypK/CN6Z+96LD8GjLg9t3X+BK9jc
rkqE7TSJ+ywQ3Ob8F0aG0pZuOaKuSyOYN5KBEUQbBUBDOOCkg4JQybqYyWPITIqw
+TgpEPJ1WX1kzxyI7uhO6DJFMncTKXEN4DnJ8riH1/7h6YeklkLYlboAYkIn+zM2
YANvTDo/+u8lNMAaHU/cq+GbFi0Jkx9KmhnqVDG6zYUbzuUZmbLjyxaD6N4zE7eZ
oJUSbFen+/4++RD3Zz5jqBjVZs+HCS4G7+K8l7KtL9pm6EGuLxJUI0mGc/HokSQA
yhno8KTpV5Kkn6ER8obo1CAdhwqV7O70m46HOPpg2a77dmQRfejSiBnGJ+3ZHc5o
uN3jvYvizUWXo7eNqqH1Lh88C+l1TNrcXghGN7J0pXWlvOGihramuQehlGerFxLm
dWQ9vTAZOb17R/wdq8nb0q7hWdRuHXry7eZGfGjBjTRDAIkpF8qeElVulkxnd1HT
MI69vbbdwY14rnRG6AWIYpttsXJAx5MCAt/M5SMjwQyRsHMGj+K2vIpLxslyc/YL
k7oE0O70H/5McHsXyIUdl1uOkZSLlinO8uB90/+7E/O5e59HZS8G41Vi2aSCXesz
lS7PQysLI6D0yyabZh8BKBcWJuRUK2n3Np2FQy3ZvSzK81OwQC2JgCGTRe5xg3OM
wUi9UQHVy1Vb7HCuTvegTwFNunyhcUQtVjhgfOl3vJP2exNPQqm4s2R1oXlXqnzz
DfXN0/lIb4gZT60EEbkCTKNqMWPr38ewz80wUALxiDyiCS64BCpv0smj7zpiafBl
2u05IWe2uoXr9v9kqZBNok9lw8B0QwRb6TsQC+q2qo5Oz/aR1bLCHLeWe0ESFK0O
Qb25PjtlhaPRIrkbOjvSwS5Kt2Pa2YEVmHx9GPhf+MHzlrL/hepOmhq9uQXC7lhs
BAYYNMjOTp03RnbO25IpWsRyMhhTVXjcNG6ERUrWb0sJng9wgVQP63yQYt3dBqHi
iG1LY8M0KBVS/QCLNU6h28qieD1eAqd82WxbUWg3KONOF1qrhFg+XG4/Y3CRcr5w
3KbXKHoVOnuLUekiaje8b7sacFjqUKsLwK5wn472h9EYAHZb7h7nXtDmG3075LUS
AWSqg6UTs9fhS7BCRgWH+yNjH4NYj5V5maqGcJKByIF9cTjPZmcP16fkop2JokP3
TbYe9Q+Z96y0RzkomhHABWuI0CTldYqLjATISTB5+ADGWRegcq85AB3Z7vrSz/CD
txSKHCLGSujgC0v3L3R86D4HN37OBMXlnSysXMDZu+VWqln6jpIm5x7Upya20x0f
PrC6PWXNRC9qey9zI9Nv+0PcGhPkcE3/2amjp+ol2rNAQLxmo/U/6N7HWGF7UaYf
GcKwvYRJD/peoqn6w/HscrNtWPCxgv/PHua384rl6EFqynaDYDWsfCQ9T/kAmnwf
iZk+rBtJUNhB3CgM9hOMTEUH8lndNZ5mB2M6IUgRSxmwIWVdID7eLkMzCoUjTUHn
9umwbEhUKI9jTH39cRE70P0Ii3FBygGTOTc1vKXXx7b1aGFn58gS6Glanu6vH/5P
/f2AFn80FfSW4Wejro0faW3rQsZVt2jDh/sWCWZHiGNCQ9zjeDZ/T6Azejcd9zTy
66qk3SVjiproypp1mZ6ww3edWjvkq0M1OEJOCBRQ4feWPdmbcE8v5r0BgQ2418xJ
0+L5qgDSqGyKN0NRry9xeOT31TlB1JgXk6ed4A9h+tzQrbwQikuueRmL0aCRGNYs
SHVeecyj/46mmlCx6Zp26cEkiwvVL/NaIW/bWN9IlO+KdGquMg/ryQ084kXTyFM6
HKBJTVeCBD/Ngaf0DPqtGRkg5G5KuEgj17oD/oESlOcveaqPqZw1ccUF5e4lnjrr
tm0+3z6V7ZAmawZ9ft7GAfvFo2zqempCnk2AQIckvoUdyWXTYB8jGm/SrDcTEsg+
62MtbPeeo6CmI3Mjic9JP4KQWqrUPJnh5Y0O4OANhwjgqbLaKlwZC3sdwzoAdBQ8
OLjHKbR3HV+SFj9vgK6xgeNx6EDd8xujWmPfNzoct4eXv6eCuFyyTwjR4UUkgOd2
SXdUCDglJnn7WJnq6DD1yiZ4T4UypCk6bK5JLbDb6sT7LZ29PhlSPLtzow8RoMgO
PmJ6GLa2YsUK2aAJizZT5MgblDw9299smF0wMfBTu7S3NlV4h1DfXzfnijWk/0le
7Yuz0cMf+lco0aBi1HdNQ3wFQDQ8fqbcXjfBmTbeb7GFyTMk93NqQMrcyKS3PjYu
tSMHHV2JTDbiA9q3JAJrtI27xHmvqU2zQm5twvFMAK45RlqcXz9kdn+hc/q2K1VU
kX1VB5c73kvG2JzMyobjTTFtLwsJGs34O1ZjPUE6iUYL1UkhDeteOD3KQEhaNord
4/cCNHep71YV9sIpD8B71MFMn1OAhAlt84XHSu7bLL+ED7DgYJB7Xr28IT5jTh2z
UKZAElWTAV8vzBr+6xJXFzBvnbaD4qfRcujhqeII/18MV6RnNpJRs516XMPidtKq
k1wUrQbJQr/E21Y+vavK9lGajUsw1IP/Ah6xRu92ch1QU8XbSaz6ljlTNbR0I87s
eY5CqBYuGO+0n7joQdm/G8CRyynAQREkslFc8rCa31b34b52yNJZykt3USejYOx5
721vWSWexL06+aVPJRod+yve+qNR/S+to2WYsKyVCMlovnHFRwYr9uuWBD5PHj5t
fb7Pmmuu0faOuAsxWXqaF8zqYsKZrC7BtwUZUPSiv7LFjklcmmFYC1AfdA/tUfnK
93XKMXsjPPZo8MOIllGUVyeY7eNh1r7jJ8BE3nbos2expI2iA4bPtLkiTaJUaIMI
lp7q25k76W4mmjhAgojTWXszpekvRzpVBnFldZFOqr+OT/0bjZ/taV6adRUaKic5
/TKeue23IpzFfIuONE12OlKX/ip/n/OxOoMEjqzAbU7ChnLSxXOhU+DJ4tkMuwIv
wj18SuEW+vjhfiydvFY+nOtu7OK2bidJTbRbr/LZGDFDwaaAiL2cqHIVycZBNeE/
6lb4XQ358UNuEiGbfZ5q5xyhVevxP7YT+rWUD1nbX6lCwoH32A/XixHTyIBZ0XE4
A8zxLIKSA/q9OW5tf3dLBbP2NAk0GYznPFHeSMjAGgjEJRmJZYTYCOjvYdi6HTOv
1J/QquCd5eiBn/9Oc/gQgTV2euOAc7K0bbg57NQ9a7M6xPKVom99TTRTNq6xo6ff
Bag8fp/kJWuS7YqEM267KKVCMJGnToNo6PoX+xQtqVlse2gX6jPuX+O7sqHstPij
xQyqS1gooSRUtPodJ7qbrAmfhY+cGV67E9ayTfnCGEY3m9JBOneo8ub1Glk9JsE7
TOH332b1UtFr9roDSz36STzV8x7a/C77JOat9pO60c/H2byZuCXqSX9YieHjdXsQ
epzBl49dpj0ZIu5wrBk7OaanaOkV+V+OEyIyoxYWWW8e86OML1hnbmCi6/VKfmIz
50ua1GMz+aOBEoYpAXWyN5KBlVmkzSOxUIVMAb//4hmZZLmQh7frhq5Wv4dqLdLr
77lHdDFHmDpnTzap868C9UOezSzt2Y6RiniVLilal4Q7lFhMdWpPfEFNBzSqgZzt
P06lGkIqD8KgI75eBXzdG4rKJ7cv6qivElAfDK/esSrq8RhP3X3W0u4hil0IGKSN
IIiUyQppB01vk34ZujwjFMyeiOpTaKGxIP+ZNjfST8sXTkPa9Z1N+SyH5eTR6Bas
QLAIGRFmJUXludN7Wg3ZVIMFGdkqttMHgzwt8+fc4yv1+P79zfroQmnlLf/uyxv0
7YSp0+N+2N96J4rzKV1yBHMNAnkx1bXa1BJrXfGJQWTHMmuBLihpOisvnRTBYs3H
ecdjlZ2kWefRN9CzA+Gcv5RVareYWEfuXv4N0/dr8R4aoQHVOGoTHy7RsNOJaFd2
Z+Yz2kszoAHs4/CaCNZ5ifFTUANPUQWh8gXvTPNu0YicNkBmx7oQJLzAr9mn9ImU
cKT5Uskx8BXsjnAODe/CwYHJ2VI0NZcD991M0LfLMTo2b1TRzdY5Yw7b20vRNrKh
a/Q/t8f2xjKECfe3yeL4ibAAzOXtRO05eps7qk87BalzHSDmyA4V4ndf757JfQmm
Bk1z3CJVYPypugLzNpCvdO/OBnhZXa4cK58aLhtli5TFrk9T28kku8+Gj9Uu6s1A
sJCBr9lsIn0q+V5yZml+/2byaBOBR3768cHY05vOYfLl2twoxoqBksI4ryJVRH22
N0qQEm/hYJZzByl4cxd+JMVLWKl71YDF23jjWXxQkC9QssyYlbC9pL3Yk0ADpgRZ
3EBKCSw/I1JFW+iL3CO7WYikRPO2sGkOHLoWf2/Qf1rq8hLPb6pRL6VcYao9ndE5
eSJm9daNJ4A/Dee3zTCxmQMZJe1UadwazKalEnNHgBx2+hvylGCzCKCHPJAedqyq
9CKrWmKfLXCcleRNxQEfMXkCagOJdR5KxDGaGq53ikQt2OvrWKwEM9yI710YoZbm
PpAGLk33P3MBZ7RVaN7b20E18dzSaL5G7NvvyDqBYMlKx+Q6LfMwAwEWwLmkBIMk
zYR2zysmnb4kcXswBHBvuHFdiKpFdw9qtYtATzZxXWgGG6F2BApzl4cuRYTv4EtP
Gz+WU///xRFm8dcBVRxe2ULWvozfEJimguyWjetv0J3IXAtG3KKUOJ/ZdlQkNLa2
k5Z5FhsivdQFhSq2NkdVw4n3dU8CWiK4uwWuXIt4zQZRhL8dOm+i6qaYUC5ZDC40
JoiHG+PJIEyfe711JjtLzYmqrIbN+tLYKnqtZDOkcNM6kg1KD42dinKLuVESvCJX
5pI6aHnhrqQHfkR0672EJZlDk1Y0nWg4OU0vlrney8HqISVfHpZFPbYPiZNOHGvd
R4+lQCyADBCGR9dj/k7yU+yddzuGpPUb8x1BGB1Nkvgq04Ebq5wL5j88+/bIRmWW
oHat+YTl+qqSd7lidyDoXs3nABh5bTJsPk7zWE7OyWAVYm0yH1HIxR0MxqK/I8oz
N0A9hYcvtae9mkxRUn1Tnl+6mMfFh03dPSDt6sbm/5qUzlyl6U4MskbzkpdZMnqZ
x78Z+nZ9yEkasY8z0q/DWtT22NhvaN1Kp2uWX9vAk0OydSm0Sc7rrehALjpNOeIS
NXMaXka8oTBrIA9gmjvp9OFFTUM20CpAsiBObVz8rYLPtUhGvVyfh3v6l5pHJp3e
Brn8zmGTC8j21i0FKeXxqIi8y9NC8ZuDsVog465lnL7+8bhgU8GPOIprwy30rOCc
HCslqG9nnaRDmWH7EMGh6bsInx8/z/awqaIM83ggQzQdY0IGLft+J+aUyWfFE04E
YpHpOh/IkWNpNX2h2lImPVDrcZuF0TtM2TjiFPNI37hWCjZc6siWq/TQW8zZPNho
ro8HR7cebu7zOxlSyej/mlmuL1QooEsyjUbEbMsR1Oj3DyR04dSIEgp9maOTZ4Dq
4FPkZN5/XuBh4S5m6AW5MyaNGAomSag4m0jVPevDxXVgrCxdNGx5/UU4OV1YMCT/
BbhRE7poJTTalV/AtuZ0UXJ2Th20aDyc0rt2F2FuSDwXa6KMpliTUekG6UdAIq/K
fyeqSoUVvJrIdAfPdgt6hkW/RMDQ+iglLkQej10e6oSDp7nAGsJZFOcmxLa3bt2H
JKs4Y5FmYW9wNbaMQ6sWHYO/oXVeK/qP7+IRK1UbETb90etfr34o89imNeISzLRU
TZK3lk88UBPqA4N/8G40fhIlT3MJUnMnFAXU1z7GAwncIC7o5rjsVryfzMyxQfEf
bszBvrv1gW7pYvrllxpn4izGJZaVha41Nzf3zzfBKOVBaRMu/LFzoJt2hIYSJy2F
B08Bkamgm4LIfmZHbsN4Q4NuLcCkvxeODM4r3BBJ1BgnOAol6cJG+FDseKc2o7Jj
PyqHkWPd8KnetYA1LGOjDp+CYAtetd+k38ytopJHWNPhfkZX021s8Rkhq3S1CrOi
jV3AwBnCbdBLOTr+oF9sbkiMbNysgPS1MDUMWjk7CIZx6iUccgeoGU87w1Y1Nscu
dkAeNvd+mMepVPpt6AQJSuwswSzQlLaNftITB/2raIHUqDONy3hkgNNUFZpHgCg7
7C/5S/qsIzV/VMeoyEJrBHN4RSvR+2Bjw/+9ZWLLRTzcJurfwQHavBMXmVru9Bek
lcpCrktWGcgfU2dCjQxuZiuWAj3L60oH5vwXKNX1/+Z7wIExNVfaAL/JJ2mE5qLr
w2LZL+BRf/KJfVnGNyE+U+ZvKwTc4YwujxQbF2Jbtsz78PYasueilSGIiJeONulo
6+buyMmyBNpn5n5nOdypVFWM7Cy3pYQxvpOlP1tRtW1begZ5sH9AiBM7d60PPZ7N
RPQf7wslyG7E+sE+sGjYT3U9zAEU7Gb0VX7y4YuhQXJYts1Shgv7uvUANIdY9IOV
JiqSr4gMRTuDFSLd6u6GT010FPc2gVnoJG50pZRZlOPvMjlK5KtCmRSWp9GbSMTJ
bhnRz+XJ8XbfyUFeZHP3CUGHZrgZJCAm+9k3amQfT4qm9Z4aZxw8gSaJrYd65oXa
zangwFfYc25KRgc/yiYbFAgheih2E7SZMmOLnP/NDZXPV1bhuWeXWr97P+e2CmGE
Vozxxw1n//tNz8ff+2ykRbJbnN6ZWmqkA9Ba76mqOplXO6SQOmPHABevLw9IpmnR
6+NuDGXcWZP5N0bKkweoGNFULEz50a4m6+XjwnqFX3hlPV7WSPvc2JUQXwE4JiWQ
4wanE7gwsMLYiDn/Fv8psasc3OPDILTuG1oewbelyH0mWXLVuQL+lcUiGkj6xnZk
eIEMwchubPdp9w3NBRe6nvWGXCqdrqKlGy6CNEUNicq+jqt0zBChd350usTIytx8
xO2UtzyJ2rNq8oww89/Y9bw9a8PHzpkZ9GrQR4OAVaAe4F5oqvLzAhUbzFXPH4yE
3dXOWxV+HTUkE8StIHuNExU3El0TJWqZ9FS4VhqrdQjOwhTkVrZdQfUzTxvNwWSk
zhgFcOlb9VrfHksukOaEiNF5eIM0b9AOLnwj0I2dQt5JYmSsugYiJGjgQYW6WDAp
RffXyCTWW9QDeW+dEQTHylaCxIkLltpt1UySHIYcYG+nRK6Js5ElPUVrJZEommYT
YUJ+r3BV5RzEayJ5I7+cXOOqcL6RMbMd1XVl4tOuhFtu6g3LzkyHdcL2ThZ7nOZm
6IED/+xntePkSO90laLsvmxW3GjiPIUQbJ2HV+aKJoUeVZdBmhjKWBMevsjqW1Ww
FjTCZjd57NprQBBkJ4zOySeJhJ5H/CdHqxm9WKM6HsbqRF/Dipc087dTi3H4X/tZ
kzOChCFunXh0GLdnjjNJ6j5Ax5sBZz617WtnwAcVDF8g4dj5n3sblrQrHjl4xPHl
gG3al/X9/nmP8eyCrUZOH9IrSw4gDPpeTywkkY46p1yXBkjRQwXIqixCcCSacgLk
64L2LvMkHWK64IJN9X1Zy7VMPzWLfYZLjUFFaGRZOu2XB+mNIPNI50E/mU4chiqe
HYv7lAkRQWu+rT9nlD9pmWUrB2armKuGBlqjkzBJIrQzQroe11MzyBnkMx0RyDHk
2FlcS/9Os7nRoeUPiKSNAAwbOG0bzk5vZ+BgZ6XuiZkysnH8ptas53e8SJdW0/13
BE750CbfI6SBzbDs1vXznHaL8rmpCVy6udONTUePlLEOab3GYe2CQWlp7HGDjxaj
MH8y7FYkW4ECOxGdrGauEnuVyNu66zStYkc6/xtEXE8daNsqKC/xCvwVcQj1MfJd
k9XRaY37tcr4C1WqR9t4vB9XYqp0iBWo3pbmEaVRzOQNU0J2LQppBV+LwOjrD0rV
e1q9URXy2zqLvahISrE4MNp2AdGu2nmSbmjxXLbUMJ05xVRfYFciaypbMLMA32X7
FrFZrPcvNqmy9Tit7UCSGU0SpzhJQuMKiIDHhMn57pTp0ZH1cNJKqb5H4N0Vqky0
Rai5CpsDtnoJz49DKzOW7PobwbyOTWOm/nbPoEyzgOqP/a1KrffouMCK6BMM7RWM
vAPwuwlnvwugQuuRUc6RD8y+6+cKtRnpp4agepc3idlZotRG5m84NUxQIKF8HE38
J5MCBRGOALSclaNuq9QHe+mghBNKNZH/9+WepFlywad7/6qk3UhvZ9gZfpLIjhiy
fH4Xz6hlKGd/aIUhZzLnX/7Ctj3ZSOVk4Lxm7wyizpuanIWKMIeEBZ2mwKrZRL1O
TFlRfVnJbyoc1Hp3JMEIgFOu5IiVhxEI+DNGkaBMkk9/j1UI/a+JXG5Af4XA7tUO
gZBU+/bQiw3Fb/uvbaLnu0u7FjwoW8jWw1ZxiPa/IKmb3AwTuavk9NtTCr3TVrq8
/IpVvnSzmAon8hF5WN+ofA5DYSyy501bgdk9rMW0U+OH6XgHRN1CxYBfCdtQxbRT
Xc7dgNTrUWcfW5DzxnvVwGnNaPIwqtukNON1CwwykKG+TPL8xXW4GBxAL8mdRG2H
1AstYnkXvdq/aL6yPLLFfvacVHZHz8CMkbPwzYAYbrbdeRQCWjPPgRSqAUxVK7BF
xyJIGoA6uLgFWOXdhIx+z0RsHk7DBjzgOCQUwMkmURvXrBh0m7ec94lI1IiORNeg
PnrA6AlNoECNvGiFrGsW/kRp77YgZIt+3k53P+WStYPk02fM4WqiHJCXAJkGHSZj
zfeizYIakQ8bdUz1Y5OXZZId+627k7gArUM17a3Q1YxRppWiyGFgYIrmvBM9O8/+
75o3bmlb8z8D01454hQJfJV3S1sOnr0UM/rFfFaGXooUjBl8TwK2V39PA7IpC63Q
sGP6k/2jqfFYnS7hMwCIx60/Mn7XJb3umVY0uhdMTJ1v/YUqgwcOasqEvUjmwcni
kmamXCPJhf/SHdmPC4+NEHE/12PHeXYNm2AqVPz8MbbbYWb0lvgDejXRr4DRbva0
VPJ/cAnXQBq8gol4ofDhTUYt6tLthvvktU6ChaIE5lKWQabghRmnmo+NbYz9ZaF2
q1/CzOAozZ6FZc76NwER43937VH7uU7IXMRtLQolr7LxAv/9/Vp404rLpUInLqrh
X5Wr/IiYVeQWYjYO8I93Bu3u56yj7Rf0aJ2r9R2jnfPj4JK+pmBgwqigXFwCer5z
ZaPkYiwvRMbK9SmjXHfF2AEIZRdBuzDfw7ifxqOPRfUwryDplD1lGc9K+Nd9KVpI
quoF0gIXc+FQQxSlx4+GvJm45F4yQwKaTx8Az3NgVrm1/HE5GHuCqgcT2iIWnNQu
MekOFkhZU5APVccc2kfL8vvT0RTHKkRh5UOgBR+GYwJKSkuctCTmBmTShM3jUq2X
NaeW/3jy/KkGtKYch38XSBmMHoe4fbT6uj9KUtiL8sjWGGOgvTe/fVYslHAeguxZ
ekNO+LhZgHkVq/mym7ZvgxF170UwymzCJKcxza1Mmh9m+UVnbmVbp82c2/tmw/m9
H/L2+PGA8l4k9j/R5g3TTO+uSzLZqLQikYLcrZH0or2/MrsO9DGa/ACbzSLZcCf/
LMdxrqOqWO+aGyQQecR7fmyfvCeK9zqMGDo1iXZkeZIxNfV7F7Sv92dHIdwGV6xd
JFT6j2pGSDbJkvKlGc+pjFVhq69PPXKR6QoLqNtiQjGxXpdhlQeoodpxRidTCY3N
Ty+MjHxCzARf/8+CDjKdjx9xrfK7u5LMtPFI9aw0mLKUpjFDJvzfZeQkfn6R04rW
bE/p299Ytfp1RIu8RNRvASDxurxWHzVIcgejIfby1ICz6QESIugITvzJh4VzhDH+
ToEGhbx/QAsE1cWkcS5D/h7cwG1aW1xh1ryFIbwdVjohg3SeeqpLmYnquZY8+7ff
TVA5eYBkGeq92ievr22lAWe5erASLrcywz0GOuAp8F+anzKMmrQXGv5KNQ3VvOsd
QWL8ShNVPxdFyrhXXnxxgwewRBJKDK6JInvbuEL4HV6Fug7W61Q1F4LaHrZw96Na
DKRoc+hgaNlX/Kaj9MTFxdkUAbT7VVECjPkXuxw8I+47Vi2F98l9g73bp36lF+Rl
uL2S66zToaRyjN5tFI7KxWPUph6qEBXXCT+ZRsrFp4ce2uEEfRQjyqoLAyLfxCjO
eIt/ua3+3YDZ5snTi96SbwvAQ7AlvPAdF6U+QOhMi1Y0vMcWK4LV8VWJ1GrtVcJ5
LdxTaPIkzzFeSiqKaPCYvdWZ4boqQSkMMJg/SCQA18dFb2DBGaw+lx9cTxs8xGqC
ZNf6N7u2x4QvrioS5qGMSz8bb9EuOlaaa/dWDETH8FZdKFVwgGJ0V1LxYj1VX7/f
BWZOTLDZCu53M/zHvuc7/mlNzE6zGDn5fsiV4oN3Xit4F51WgEFpxPK2as9mDTeZ
OwwALbOJGo7JNL5H/ctIdIsAQi7jl3Ga2gJaKnQAbMfnX/4BNyD/KYL6bU3CLFQ2
/WEgU+n64gFIefkXriUyLCXSB2ogACCxJ2PAAoe57EDXJwDl/I8PYAiL03tJneqd
kCx0c0/scNyc4bo2PpAeDA1PORp8gpdy4i8Q5M6cZtytr4zPfemnupYW5+lcAMt5
zniqRwu8YwjfFtz7tfClVPngHNp7VXvLjk6m0gUOsaHRGuZmI6obfk2/2H++JcQD
WZHHsFf56IUN6akACh2KyfViSKJpvINS+cRAX+V/3eviiUuA9k0Nt5mPhB2f/lE9
vIGqMbcIx9WB5JoMA1ssa03L1NU5Mxp6f3kXLl06A4Eb2xqqF6Dohe20wbzlwvXX
gnKOjCmrT88yQBy5e84Qggo+bSp5YDBkITauTKKyl6A2E9+97CPcAPKX6kuC5qlW
ZL2BqatAXKRQu0KAPXMAQbcCwWVVOWSHjanwfaL8cyxrxlUa/Pbud/eZbn4SAcrg
ZBMqQ1MBEehQkzjcQbVN3eFCg4mNS9T1YmvlkTz8Tpanafkh70BX1GWiZ+j3fMap
c1FPo8hWEW++cLcHeAgqaLThA5q9aqN6nn0lfxWhUkyDaH03bht/BCAuXzWv82od
AhunpW2wvX4tWcncaveGc0fjxRja/TRs0NigbdGBztOia4K1DcG8XU7teqauZohy
zGIO/toe5MeDXDa8QCKTR32xTXmCQV5ZjprCvIEOU02W5CJPTQmmKhv9gQP6n7JK
dmt0kWnlO0P3hO3BQ7W86VyA9BzyUw/oh7/+h7MvvLOGdOJlnMyWvHF3ANZ4gxr6
dVsDBcz7s6CXmTC7oWbDAGnIk2hOWlQjok4ttVSG+Z4Wb3wlI3Ndx1WmqJjJnaH/
vTlPU896Kb83NkmpYO27y+ZhVGBz/e8Brhg8/GGlxd+yldxUfRfGiHH3Rn3r8iyE
QkH+1ysTawOMM39ULl1Pp+bali664aifJoHB15O+NogPh8cjcMk+GAtXt1N7jzIy
I5NjYjSqXMD86/50fUKWt6ohHXpd75sSrRddPSfbCsP8s2uwLZF3DCEWkrJCk7GN
0de4iL/KAfx60q2i/QDH/ofQzsuXz47REWJkC7K9s76bTfKjpQD1DZQE48mnXW2h
KbHxljpWl+TidDHDUhEPAnWfICAWPwWxhOhEirTKUnqsS2HSitHsfNVnLyvAQIh9
B492Hn+srRI6zaUcCs3AgLvmA+ZE5QmLqHoiBCEejr087xlZ+DhSK/96kHeigmwT
FWqUhv7bir1yzI9FTKr2ezeymjUPHTAAkOSvQ7iLc8gI4nWgXeknltqlPbYduI8Q
Bvo+qpp6BTlZlDaUs++zoe+Hk8NWx8xR4fza3CH2b8ra+MnO8ed1I4oyi3qdTFiy
7RQ5Y90lDJ+jGLGJbMzpLtoOXzSW0BjMaZsWb7EmyFGvvUEAnhx7Ujxj91065MAS
Kb5oWP+9zKPaenLZpAbqBeUxNEoHwxvlnp4qijdWDnMdNOruefIhWoA52Nph/s6T
cBArNGyQu7OHnHQUcD2ht8MHRq+4GzpxuMPgNvUeUCuuEXweBepFMrBQkeCaG4Jx
TotuQSiczKU4tXDVwrWG73FMJhbaFU/9Y1HcX4D9l6+Lkjk89nd09zHRlCXIF+6d
Y/FKsfyBuPC+W2UZQ5r90KMN6rQOrcYn6gMtl1+iow/ShFjT4djwLewCAsqQB71j
TOyXaUPzjtzr05gOx7ssf4etn4mnyCIF0MEoX8k7/WMRZtOPysoqU0k21msUJQwq
5RTc7VQa5ltzm0BbpLk3VHMrh4nu7kv3AA9m2DPX2rhvlFSB4oDwEtzs+hfEVa5M
6DPNs89GLSkjm/pjolXZfaQa43mW074SvINPOUT0E/0uosXfd/LeMkOEfBupyz2M
tt75Q5n9Mt4gvYfueyypTon0cxyMFGyKj+GN5FjQpbfjB6Q0mCyWEY8mk6KRPHP1
uUzUJCMN86ygu8p5EHx2DC97698S7Trcfc/8Xkf/4u1dJoX1l+JY2d4V24gtJbKj
AAqpopAD/7ni4w/peAzB5OZ/xiyB/4yR16D1+RnS4mTE2YG59nzEgGAMjwvmsbrk
SpzeomD2iYKJyqBgAxKWtXaj818Q0qEftnrfZOOcPPOCbfmsUoden0UUEGF6T/eR
TU4+TsnyOGE0oqT/F1Y2Z9g8NlzQMlZNsZviAvjSx3B+6xCzjViAIqzG+Uenp7h8
Pi2TFaLyE+ZoIBcusFrksboXjI+2wGlztQ4FFS94mgnsfviicgwtIANhARuafKNS
RQoOr79ZnPx54EsN1wPpo7OQJqr8zNdcYz24s8VZgcIKyVU+l/Duq0VUXeA8RYFX
0APxHxWNnxScha8wnidicoXm+SQ1BVfdlLMqOxAJo0iAcN2sLYOMLi5beEp83CI1
FWQpHxbI+F4fCUDPQO12fs+pgbJeu3QLTyWkcAB1AK3PZWp8vBrzAA9m1hjNhOe+
/QPEj6BHsRda7ttKJ2NPwKqb2Gs16TEYCksSPmFZehXyXnAir8xN6NWnx7LYWoFO
FqNHGgERHLcVSNImmh8JzycbXk27l0riTSQdpC8W62KROaSrmnHW8xOVsmV8jEj9
RWbqNyeIM3DX2m5NDP9PFVlvbul9mhFCWpkLh9v/lLdYQ0WDjol3+U6Ulnk/DxBq
1EkEQ+TEy6dn7bRzlDy0WAqJT1/OiJ2MgdGW3LZodD+Azj8Kknut8N3nS06iiQPB
appyK1IXDHKYD11n/t3JlcdTCyXYgP7O+/AxBr6wqZaxbuRta8p1xSaU/u93/psh
26ORWKS1lzeUSr5SQ3rSYDj+DUfINXy+O5R4nD2Ic+1ogFH0LnA6sYXyI86GClBg
7WLrVmoBJWvg/bx9qcbR8XLAZd7EHiZKr6AFRQ9oWY+a1Hf1nTxtZvxYx7PFaQ+T
B6muBzppzsq7S8iw6eL0z/lxZ0tvERZ7oKTfnG2A+ZYiP+Ee0ER1fox6jjjq7Yr5
OrH+eN29nVcHrcvwafD2uuDLqeXKBvG5zRWJH8sMim8RqCyFi79JUNCetug0IqjS
NsUOQqXg3CZXTtIbOrmalgt5KFC83MH8Ou+QStnJo1Lbo9xrWQcdOe7sUNVRLIX+
i2m1fg3CWA8YgMx7owAnucKXzx7BPb0JHwVIn9XXKD+mfeFTpycUq0NMCaP56jcl
XwlxoOPgyB/W8r7anTZkX4HZg4JAZYTgmPs+cGqdRoO1C0IQXXYQ+JZxIv4sZ859
NgjD8f+qEpc+IlXR98DOBb4HQUZpGpvl/IZSuMcnQySY2MbKlqCrtRYryHkq5Fbk
nDpOohg7hEvQxlSqDtJ47KDSf0QB1xN6j+yfz/T6gix7OBt4kQSa2rg5xmy69zDV
BjXd96GzMdwJ5njrZ1cbk9UugMz9aN9zCcGbP0vhRaO6v0pKr3kmJ7MWzz0d+Ggm
jtvHRySjQLmHUPsTAXEPCM2Vjn3jnQtYhM/BMcnAEzXSuJSw+7TSPvmzaxDJI/lv
Vhj0+dN1DSSjUR8IqpvrdNg02w96jgYoj0BvmltcQ1PLDJbaGMvJIwi0sBv5ABFr
kTvyT41/7ak5tnJR1XsGpNDx6h2YIHAGSxMfdte94YYKM1oS7xBnTIwZHsIyibfm
V5tjn2ALhOB0IfwxwLQzlabBd9252wSiOK6sFRGMa4UxxGgmGrebh65gcEgOCxE4
sjVL12sQlHEEsMd+UP0LcD77ecjha4nQj+LeXLEjcvuxtIq2a15p32QKta7QNMyu
zIqDvFn0wIlZBx6N6CdA9lc3saBA373g8KOoOLEnI87u9VTVgRAH2Z7E6ZowrFKa
VTAvEklyij/Icvmqk/abFLRiwpGAABFGvxaPVZhb2GzDYZ0WBGSmTjttPOPkRNSg
ogEFNyPDpEjTG/rLkcJT6XPYXF9YK2lCIZE86QV+sXnyZXtfPIHKM83tcCKx+aOv
VDPOAOB/wmEe2rcn1KIBMFxe0XtA8CetX8XNRgkPaeQutjadgzn5TmRzTd/UW9ai
kV2UbzE4Ul0EsX5to1+M0Iut4aPwcW2HrSy6p+TODuqjyKKOPazhGdKFeLBDn92S
l+uEflxvhnFFmKJ9Arlz/cnPZ23+HdUHyhiK+SYbtA7irmknDndkdGzd4gNKJEF8
FfeXaDVh2InBduU0ofihP+fTNDJQuyjXQmJ94yYJrBotJfWFvZ8vAg05DsI76UaZ
tmEPR/afiqQ/TknkiEDlFmCaI1LANeck0gh/NLkRPJSaI9oDCFhd0+yOnDuZbNOt
FqYFPwZnwrksDFYvq6az4H6MQnSmgntcYpOg1AdmvYKRBbgUUpO3JsC8ErhlTPvh
MYWfcKZfuSDYE30kZG0EIyX7th5AnKfwzAtlHulBrsfWV1BsB2EqXSNID4uZZJej
hJvtbXvxu/9DE/+wrRL+7ttgBxkIcsxsarp1Nr1rKXrPCsyJXgPQBdJcTTHcDBtS
0BJJ4S4lUzZtr5UchBBP2R/jxIdwjcKsHK372DaC9Fp/5iXjhH8stldo6jUrOU4V
D7ggXpfcqbEVF2mmBXslFwZy+M2N9hkrud9y8Uf73Zy//tcpuAjvHzYVPcqJbMR7
nibiqmSvevc13rX0Ku6oAIc6ROOB8lQZTP3EH522qFa3mKSa+QVPLsMf7cJzB2/M
IQrXGhDmqN4+bPZEu/v43ijMZ6NIcHm4vLTZcNArdpqMb2aAk8ybA2Q/onJw5y9x
AQCmGlxGu8YjBjKc1FjemtJwi3sbUBOnd47RLdA02Y8fr6uwsK4AadrEr8iUdCaa
crk9vsc7vMd+GFkdODXU72G9X9x6vlUKTKbx00Vb5JC30f6yLXGE9woMAJ3+LZLf
vA+QbC0kvcz38uGdP8qQk1ThgTZypCZRNGifPm/q4xTaNYFiBSUBisyBrDa5HC9c
aVeVkFd4sEHtVeF3lskDHLhySguVInMxpoKkPN/okdsF6Xu2jJclTs9jlIlx/mm4
AmaUbX89D6EjcRVuTwcAJMaegQGBUartzISq070UB55dt6EKQLu1pkugtQ0NZ0mF
5Tyi/UpdHKRChIfSSnsMQ8z1ig8NwoBQrUnEKGS4uVuMl03/wIT3VfLWzBWNx8Ho
9XnqB1hMDeHvLINF++hls1N9iZlLK50LZxzsQlQeaZqu/F47IsuWs5fM/T4QKfoV
3FENIaUwBDZ1JfAcrnw0IBgfYAdnYCclOU0yzpdMpR+z0eHmh/1IoVCJ3BJlIIrx
4gWE3rIl3bKwqGH2+qFsReK5m/LzYp59EzLqRvgqwxbj4tGi2Jc/3ti9JaziabP2
20WW2agLl/Ty8OP/YqHvZ04Jd4OxrUNvyUaXrlLP1+8VO7Nw+Ocdnx9vXjQQdOS9
aFENHHgVuG9C5w6R5MHTINs7K1k/ZCK5CssEVw3MX8zbSpke3H7vF4i33zOsu4Tx
Q47ujFW2kHP6VkCwUnFGBVP4h/tOwBCF8BrbT6T9rV2ux2EgrkMO57IzP2NF0a+F
avlIK+YiHlSDy1tYL8tk+Lk0vPfZkws8NIqeMKYe7bMTX1CRI8MtLF8SGvQ48X45
ORlCOAovDd+GWLE70Gzl5ELdZuKR26amZEiCtbqZP0MYXU/xcPi7U5rg9uwGqqgf
/MaVVmBTjhydF2YAX895lkRw8zojlgj4sLbD7SB+yhttPLpwZxE1Y45yhNudpWBu
BMPyVQiLb9sxx0af8tLk+E0ydJFFXeIx2+U6KHJ4JvK7Y4Rk6mTCQaeQV9jqrYYl
mzTW1O+1t2E0QJWF0sUcNl/TUFow03Om7gmcUDrmKdAYDwc16VlY6DfT2OF6K3Im
HBCl0BN5l5G1zmU5LkFrrDq9x/dD/VXFvGlLmbSVO9gk6QuK83A4slzO3e4D3UQd
y49Xkcu0YYOSDvh8+QKW4CYtx3rOQ12qeiEV68lBLK87tJwXfjqQ89cme3Xddot2
8d+/NKkENbGVpxDfjfI8gGAn4ON+ZhTXq+8NDB8O1r7wGDDec9dlX4V3P/GtLo+U
IltAUX3m2Jd3Bi5Qhjw1WZGV33PemjaJ8ai707VgSMeFFWtby6Lmu7vbXaBRTl/R
poDNtqNe58uidZeCYVmD3+25OPTNl0TLlZbum1/id+6WuGAkg4DEKlOkxpsIzgiE
QKqZYM04CtWxer3/p0B4LVOBxCujlGkj0OHqFa4evvBXhduoPTw4498OjopLCtLM
GqiQakoccHvM7VgFYKp1IjosFuv7Bq3yt+120aPb6LO5QbJ1EO59cEgYWkAFxY6T
zwtvnWQ0BQhMx/BN1y4VLeOESIXwQ3YZV/bOAHbiRFXsBLYdpeC68D5hDLg6NgAM
FiKvx3WU+sEHUItQcdwFoUxdO4GuDT0aNhwk9DZ5N4XHaQU1Nxgb0oxSDgpNd38B
c/0q4JUXsIe9CbDJV/lZAvFKfno1DRIZlks9X4oxY3Df2mAKgA5yCOhNsf1QxRw7
tTO27TE9Elvh9mvapUh7wVEaf+Xd1kl4HFQGO4LpXusLDt19rdXxuQHlZeGK2fQL
yPLocbs/Q00S9/XtnHrtATKM0A0y5epJD3mx1IJQHt/LOdvmZQLIyKyC+GhFA1Xj
SLmbnxXqSisuhi3odgsewCqwqF8Ro1SCulFGtjM34Htnf5lwk7muyJzSbYsDRKTa
zsJVNAR4Tiohk96pEWDt06ployjkt2tv006A8j8ZGJE71csc/I2tAz5gD2mzQqAT
i92htj1u0d3I+pGLx5ioYONDtcx09u5fPRqclJF4oLeOR46k7iWvfSR3tU4ORE+p
NeFSssjf3I+DKA9M3hVQ/EgC3ulTfs6RB6MmM+Bh+4V6pEWk0KmIAjW2hi6FWbZt
fIez3B5fXFponk2gQr6mqKt+t04WXBkdO28nXwvv0bTA2b/ay2huEJRMyJA2imJy
cs9gzPWw7jUVEGZRdEVt7TO40htX45veGFvjZl2HWjIhEUTqE8veFI3w613CKsd+
f/ZsHs9TswgaIogFJhSyebIu2v/8J4KhRpeMGOejdq+G87UCjxdVUAsbfkddJgRX
`protect end_protected