`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
m7OJaCYG4D2XeQKzWhbYg9nukT2Tfck0vtR7DyRvys9v0FU1jT5mWp4/1v2D2ITt
yprNLDSD0t6m75WLNc9+2ywsaQ4nD+B9zjg2SMcZj6seZ2uuDCIqcYtAz2epoWoq
S6VhcC68PSJN3p0vgQUxBfE6WQa7+nsk7cnTddGxfXczlKmFiZL+N07cPweU73Zn
jIxHmmM2Le05yrP8hB9HnPJvoQthst7KynDTCsnhsyRdLHlRlDRCZbsEWWoZio+H
MLLT8yImOTeCPHL27kioQiDZ5l6Xhr+0suFGjubLXpyb1edTO4VDNgWX9K4LyJDM
yX9wBCagZnzUsPoDDBbnEgg7p3uGnOQ6eoCY5BMAp1+P7MJa6DfxgbwsLdVyKZ1x
mLmBGCjuoK0kTVDWO1oMN2oXnV7pqOYylBOTGrpe6PCmcH106d8RRet5BFsaAyNJ
4UMU+IkyulwmlJlZTSvXtCOSTV/1P62dGwo2H1MhzkKGabtEChrxp9creeq4S+ZM
NIUkT+4RBn3t6RvmulDgP7VbCPb9iHvk0BbxzUs/uM27m/F744llkTzN2pV6FnSm
B20KwxM+GqJe9Mxfv1DHOnrkOWa2baiZgak42i2BA+4Oj2NevEQQetP1fk0GTioG
rMYn0m8KV4KAFVSAb7vYGpReYe4CbUZLr6MhYLyDpNqynXGS4FevBB4Pxxb6LWuy
FMmyxXCNCGp3V2YR4G0qMv4lT6iYWMrX2Dlhak0Nb9gHUPUHq7jMNslji2lKlANx
V5qIbJCNIYz9goI5doXBV75Rat8gpwIPj1GqkR/6R9pqQFiMsfOenTRCMVAres9m
g1AWoTykoJqv8ofOvukrU7SrezXaUpr4kwNUQ2AE1lV+fF8f6+IgpvrmxDZWQFag
vvmhX/QRI4evOaOLVlzaHKdNayzSWiv/LWATsNdfPKYbjVh4fWucfOHV3av1IMG6
sbWtzii9WPlkq7oxhEDRjyeUaFNgM4YNqSMDmdDhsc3bARl7sOmw1gd2z5fNisYl
e3qcGGo0MoVfTlNOsDSu6/cOIdTbcRffcLayCRakDEunPk8pWJmlTDzVMdKeKGN0
cSa+rky8QhPrNUsmZ8YQpTw5ig9eYBXqoAN5i2/ZqLiEThBL3z/MwFXSndHTRuUn
LsT2CiB7bLTCaUyGrPcPnQCaPij6VCGtLWpVEmA9EezdpWDL8DQWWI4pwwj7dPWb
0gstT2w7/SaEtBATIunS7abRWNdpLCu9whrN1pYi2fN8sqzvl+OzH1phoUZntCgd
ARN0doaFS2PVg++vSyDKKjyOBMpuEN6Djz+25IVmjkRIbVJbbWOL4yI8CfQ6ELVe
xNAOgLPFWPShjYQDDxLLvTagjp2Xe0XQ18XMemP0zIznsvD6KegIWbLy4PTQzLTH
h4baGYwDSwt5Ii5/8wPGUPcmeZxAsHbKBhrv9l/qLZrScmEP+kJAeemujgePIcEP
8HcMFT1XKhlzKHdmfrIqGJGqe5AxtQfL8uouGDPR1Nu8mTlrLCPrF0M8NtqPEv1C
oYdd33H7CSVxG4unmSJdYRf6phIPPjpce10gKdgwepylz6qjaIs6hMYVR5OtlSwv
r0KriUxtP47cyk4/yAhq/H6Y7RFgALI0c0caBfIg++Icq2T6U0uzOog/shQ6G1Xk
A5G/tVuEM2vlVpwhksaV1orfB2vU+EOYOSgE4Vbmu6N7VoUFQI6yM79ozIFcX++y
USKREKpNFBzX33fwtRNg8JsBpLQ0Bxqv6bqGhpSsO5lC+CHkPJwFOjEV4Rt9C/7i
TcxPasSSVdgBUEptyolIF6gGeMSQ1hYjxp763qAoPTxFluO9vvfkpLZ3eeoGhSB/
xqbOdBdJ/lbJQFQZlJWHyuyPu2jzda9l10tJ/AseKLC81wxB8pl20aQN+TfCHtqK
Eiu4IL6hScEjv+tkff4u10RZb1Rrqc8OKQJU5X/+SP6E/8vtTZP6WrTEBUWKYQ8r
M8zvKq1UDlGipSo77xK/gt5koqhdrVuZ7q53sSHTVuT0Fs6ZcFs0njeJibbzmNN5
gWtW3M3cbVXjkCrqtcmx/40ehOA5RyL6u+Torp2z1frRw2t+gNIv0hSvvZ1sDK3l
Xxf5ipNkLFm7vUutge6WhaxFnpaLeDKLbR/Vb/aXG+heh+p7Avki7Eq06lDicLlQ
gvlPV5Q6IrWVAT65MR8sT8O/sgznUn5pD10MDgcXR5nUGei2SJmUVdKdlmwk9dJG
FXumVYIDsJ6J86ELRbNKHaHwgylHR45M5nnuo40mk7LzhDStZtXzFEzjKCDSY+iL
7rnxb9cF4vBg5R615cD0ToYeAtvMFS6/4I9m1/LiLJNlV813rllhu3rWpTo5iUPS
xhi/1qgBVUc+mzmdeFM5KLYrSXR9ay7U9xXYLWYQMf6o1XZ9z4UXgTDltzz75SUt
nQ5wuwFPFH3fcF+c/rpNHyuydlLsnfGGUni3SnUtByNnzUEMTlJKwCigfoAq/02C
jWiExdQXht3q6xDge6nz3M+3xaMHOBQkVaHq9b0hHG12IB0YrlVYJ6vddr8hd6/u
`protect end_protected