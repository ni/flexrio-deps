`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7184 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nn7oC/bbltaB6y9f4wbJdgh
0G6WvBg4Flfb54G2gjKn2xhmS1OPDhzh8Q6RnaYECbF3NigU8H+tUecmdmydVHec
utEk4ycFg0f26Jqa6ZdEo/NvaUasO4chDnXUfJj2SdoeV1J/H7rNXfIoZATn3cTg
rnBrTDeV72sGarA5Wxu0X4lFGxOxwysmSq/Pzq4rl3j9IOTTh1yKY6ccVkofqB/Q
Bk0mJMhnO5dWxFwr6PzUDzzym9jMqEEeH8jumsWPSmIvstfcekHbpPq4OYcQoxrW
k9zcYWR7xLiF22OmDU2/0W/Le5ISdUsAru6xeZLHxK8V3+PPdgGHYvGc0k1ZvY15
Evb/01WU7hSnPKuydw6+y1+nEBBzfFnG4R+d1EalDIxyae2HV5tPfUdc/pXlaEUQ
l07vXWLoY6Y7yzM30vkNN/Ai28+5cA+YacJy1ryHRDWVBu04Yx3H7q+brwQa3UpG
EyXooPgkGIeL5kaVOSfKQLmVxEl7ztJof3Uh3kS6XAnoSR4efGQCd2rekt8rx8BN
cC/sKMMsrgIJZElD0gX1WPquNly+kUnxmuevyNZ9nRoCuPFuH/Ted+pmmBuM0+mm
B9DUbB5bbUCtaI8yiRDILz8SpkVkOqe7avnrJNIsI1VQVcvp5rblV3VVC14SRb5Q
Fgmn2uk/aRT1VpcrepkZrEuHTZdq2Mxs/j2996uLw23GfV0AkBfJasdr9L9uu2qs
7iYVNcTAhEN7FWuU5KrQIBTQXQTZB4+EMOPY2he+a6+ufY7tP4tH5/u+5s70yFN6
IpwPCSeFGGPaxa8WXTmySnP4omzKUl9gnQFa7YONAj1dz3rzEqKMxy17fbh2630/
9mA9GjuotgdqRqDcwozP/hV4lLPt5gpVetuDEa49ik+74uVUmOh6+/I2tQZLL66a
aSIkMyeFWGd0NdgLqTxNV2uX/WtrW26QgtHPGCYri1LOK+VWSSY/yMDZZnTqvEEa
by1mqgMafenitOdFwx0KmlNzedpo7CRmpo8ZSvOOXO3h2BQhCPYoSQ9F9+aQ/J01
HhqyErnuHabvptLUddlmSD1gB9ectXk8pDeJP5aRcW6jWSR+LjN+fnZo48NYTfhM
BGpaAiRKE+0DIjb9ijsDnVDX9332JYjmhGbfohuQF4UckogoL40Y0v07lIEbrAwX
ODJz9YUbaIOMp+0dj6jGmKlzPuRBBaZd3ZC8hJj4QDIMzGKoo/I0o87outpJl9t7
XM6biQXZrSxKHbj4HZ74wRzcTYr8oF8cItgA4u2Z1o51+Ii3NCI902/mIwqQoj1r
oX/F7M1SEG9RpIetZLAeS+IDXeRXbzsrtc92cQnmI8TPJmVr57FUac5SXtkOsYIL
kjopaQmACFj8F5TTyLUErfPjFnCJLOeDIS25ckk8+c9ZkujprSFdUq3oxxP8yU1X
xSSa///fxcDsoGg6SaHl3i+qtzFIKaosFJvQqkZetRgiLG3OLNNsqxQCcIRpvvwv
pmtyF1xHIeJZsqhlX7KmCJXzsu0yXk7OQUizYh3oPeQn5drj4b8Q7+/CElSFTlaC
KTQud8KD6nSmpEV2H/TpPUgf4g+PlbY588JA3k8Z+3tdHQCcyTyJerVhrY5D0A7U
Yo9vK8jBWYLU4k0NG1IkKjAx/TzH7yepqnUir5BlTAn2P8H4A1dF/mWs6m+h6UJL
pvosV5dcdGmN5zHU0bRn/mP1tt60QBoiWUYverzIF3G0Gp9e7bhATyKvkUsPllAG
ydrhexwGs9s0VMyhA6EQlhL2+glliHRE5TwaflV1TpMVl/9FcX50tlko7GGjB6ei
vBV5SmOuh2qh+Bj0Abx2v698IutYX9X96hHr3wce7ti23vdFd6AZNzTcGL9qaaSR
9rvKomNeKzmMELbaHTUBqnOhX8BXEGeZvCxg8tevVxEg9nrFIbeJ4W0RnzHD3116
a718fFj6/u1MQQtPRfEZv+q1ZDEqoEniNxp4jHIhJYYvy47cpmDL4E1lddN86AEa
mSuCOTgljtIgus+jkAV+a86F7Pct/2yLeE5R8ymVDlhyiKX6HQvn5OSkj0opsiek
6/LvbEDNU/ujaYVm3ghNGWb/7sCFNDtu7cX1RfcJDYscA00V0Ve2ltRkD57hOHAf
habi+1sNgRK+Cuxm8fIzr2eqt1RPmI6JFLjXjVfeG+pl/uz6oHJcnMu8mosIS3/z
g7YEBLmivTSXW8UaEbVvAaQH0vSHPIy1OFmXj0g3q8PNLad5VBQgXg5Asci8+Fg1
dSxj74rX18ikvgTHHiR2TmZTgcwqhmhByagBLiBnSlQar1tFApDoIZCBMogXQTJg
yWWfP5diUD4dQwcIwjCEs2eP9ZSq0t5pSbVblW+N8wGFw6vJwFZeuyYgAPXBCQ1Z
wU1KE5AEhx4nYjkasGNlZhqHMk3FBxghhcvQbAWyT8zxiKSy1KKQqsFRUMd75Bp5
ccOwgO1vfoclw3GiUoXyP8paPPSHKnWPOneO0o7Kl9BOfRz/WZyXcubMKGoWJHoa
2KWXpLvT6mFJeQbma/0jqKY0oONlZXJPoKHMu1S+lMeY4LrzMWNQdF0S0o5UWi1Z
QXPhlrkfQ/YwK7eJE4t2Rj9HKRijBSY2ElCgg/F6fub9EjFFNLvtuiRsf5cQEHmb
3tL4OnLQqYxhOmhq6BO0c9vn79aVeAW0StZo9o/8k6tMPs0sLAA7pW+OCAveF7Bs
baU1fuuDpkALBWkd71Q/el7JE/q4XGv+6VxzpwBFXtckCALkduyDSMlYmfkCeIiA
CF0gY6h3rWOYDZm7Z5IQGPWJ09TFqHvTkhAwCDAznGfNLni+41++Kwg4yxY1Ax2g
h3fSftzjDyC0nB8L0/evfo1jcvvDSUnpjzfOI2fSJHFgQPT0+qJ4pT7H7+RxBsJV
UIf4MLES85b+Jqxm/t4g1XFGGLMJul+rHNAWmd03MzCFFkEmnhmvTTjEk/iIIDlP
pvx/S28ArD0nuRUQjazXfE2tpQJ2t0LXJD1dgNwsPu/hSJAwdhop+58b6u7SVDQB
SEn+T/0yU8lyLVodJpxdHJ6kVer3pDMbTxkHO2/I7iWU++l1KVOQa61GMvHh6HUE
8W2f4sABBD+cr3yZlp6zOp5yAUC6UNoeBXzu9uiXTJQSbbkEzFDUBBVpU1/ghKsR
80jJrTMAc+HMnrinqgyKZ1m88K4PGYQEnC50Lhea7z9Jjn8WI8ZctGzIsEBJ7OL9
askcXYlhoH07cZh4NRq4Xwl7l40r57QGtLZQRtFRFktaAMqkff5uYUdASuDEjvcU
K/LgUpFwjVHAidAuFsdHktkTuoYzTQCunHofWZFXvd7Ki5tTRs02vdp+Li4PVROc
LKFf6vLP6kVPpeKKTIijHEaBeNCgy3y0Ucsr02gxIsSQieElaGB6vSvGx6A/oXpg
5PY2MbHGVW0jOzP68tnQN4oE6SKgXptDEcOJRj2DaKtfpb7tFXdWVIU0tUrlgZ8e
uJX+ukyBH2QypaDi/QBmyAz2g9ao8EhZUM4S5gLwzr5FeqGJYd8onfrc9AAjxPIp
upnL8I2Nu+RHNWu2Za2PZ14B99BkKQ98tuH3rzE/N4BymwY6uB2fKfdLEBfk3esP
DeUhSIG6GYJJpvvUZmdRg+9kbZDrfCLUf7D9MaFAVofMn3izH9e8NPXdZiE2x3bx
R9pmYLlGrONYHEZI0chdmwrYH17npeZsdBD2tAL0Sp5OhKnvyoQR4Y49jxUtfvIK
h3jbsP0B4HlZm/AQ2RWu3jRH3IvZycL0ffFKYKil7hUOej9VNtxV17eV6P73aJfw
ET9V4QzFthYCUh3Uo5Ju3WF+4/4PDP1Lq3W73koeExPyRvRyiHCmEiB8dloDbeyD
1LWBuPV1TuWcwdU+Xt6gOowLPMQ8P64h8310f34vnlmMd4z5ec/m8xsqS+l30Myg
D3QgnbYsyucmsnHi7m8x58zw//0dt9R9S/2ZRdaHnKtDTozd3cORmYs4PL75dbuS
UXS063gaqrIXJcL0Eb8ZWaHHtbH2BB8Hpg3zlF+wgsPNSdFt6T+euLT8CQShveQW
mSls7/C9HIrRjic7h9qDRWtApCwJTyXwZgMHHyb1ZAbZbXIQ5LBwYXW4K70nT46Y
aQucqcFXa5uR9NssoPn8Lbyjjx1KSnLPPfzwMeTf9hGVtpDhdplRnzy2qXgF+zDS
TCYqJuxYsB8kLpqenhFpb4sGtUYcsrL5q7qRRh81eDktb4+BFXD+exKtRL2GL4Qd
LzjQyZu1w2N/I7d9jWrNxdVXQQqAod0bv+59jaJ5f2PBx35TIpWtQxACmWM0rUdr
6+FeqpVYRyX1ARQIyZE5qseda5fKfB9/DVk7SONdZNx/PSXTsTNoP5IMB/dqmpbK
vThJBNe2UMtyCk12sE8asF0R0jq4m/8i8H/oAedtthAma55aoN3KVWClKE774E2r
3A77QdVXgNvDfFe9YzOWW3d2Lb8hevG99wIoyw5cX21GrxKk8hdpf3BycbTBB4mq
goC0WFBd0LTPHce7PXcwKPBNYKADSF3x4TuQhwnKHgzcCEm0eb2+OMSf/A1Xq4XI
HI+0u58d32Q1b7YAAklPeehHSkdFfd5DBETYh8/qLcVUK+keps/xfBV2ZCraAwg5
yblndonnTBJSPJWABfxseNfC+j54ZedpXDOMF21bGrFMiD6Z6bijmmu8vSEITB2x
MZKIKY02Lam6GLpZUpaS/p+OPNSbLBdIN8RwDn+pjcaoVq5rfYSVz5b6oYj8QR51
UiOcQ0AcjY3cgLDZHeLyDqhDvC0bDKQy3tZdW5tmrsQAkH2CnRUaqqR3/SdRZRkG
9DFDCb/zFE9Q9HLvMaVqBnzFm1MRcZhaawiIf876nvAHz5mgSLRbh0nQEFWCdMtv
O/HznI5Emu46LHSJwe8bRJfpC8NOuM1bKtbv1YskNbFp+5kDtPIOzwG1GlW5430X
o+GfTK2LWhZLepiiFWkJ99pCpFkUwQukiKDGzBDZaJ0fAReTuWV3xRkqSGMyAu6o
qiaoJ6emrJJCkiDVZXsKFUs/dANmGitefzE9z4T3DzQ6h8/BRa3daqmwcP7ULYty
PeDWEcWLxNYSxW1wDmvuKjqVtI4OIjhyOlwDUyqkBgJ63neAn80Efm+yeEXb0CN6
ki41nWd69+A6FjgsptCMflLetNKWY5w83sQ9tCdqsxHSubCOhkjOQkmhhFhcLs+U
qiizd8R4RtQFOvP2gOKisKGwwhAfHt7ZAAcwLOEqOmdv7T+cgkaBSlsinWvAeQAo
F0wNhCFY7/6cxuc0BDhTkQuDE+A3sDnfiXSjqjOv0sPRF0J7ZusVUOHoUsJ3+vrc
jwcCyHQizG7DpkifgWrZAQksEOgDQxLx8vwK2MBSpgxJrWZLBAFWAP1NYUYWVMBf
wH3HXWcZmT5YygxtSVzYRix6h7m4iFehyFutct6JF0mYISP/JFebdfdz9JSLLQN7
18yXy9IuKCK0XKvMrxZcuIaCIi7PhULKOuYt1/Q+iUiOrOFZwp3MPVjY+dTx6exw
W93cZz55Vg4B/zOo7OPnhsaUFQNk7gu7f5PNqpNIpEK+PtuCkOLPxuQEVv4ZMcs+
htCXdOHFNoOGzVWAQk4NbaHCQWKLosgOz4AWNY8kaQGIRrzjEjJYTXXaJG0wDUTd
hxkbQyREU8iaWbzE22DkPEcrmtJbaxavWu/U7x40mKPH1IXBmMiJjRyNPXJZRqJN
DZxy9pBoF90xBOcqUy/4KRLRzuVOLTBB4zl6J9a8ICvND3B04tvaXq+TjCKvwrFz
JWX92iwZ+duvZlUmwocKfBmO5hdGbyhoysTRttpZ8/Oa1ypPaLtja1Y9OHNA1mQ0
ieSaU2T1KGaFMTTgPM38HBDv5U2ojEMpKNYETQTIbatC0D8diyNV1bWsX39+90es
DVBstp/QwFf3+8mvuI6RL75hF7mHev3S/eWpv/MkifxhFG72X2W7hC+6yAQgYvYa
3w34biUhDSgjcIABDpvjkCeMYNlrQSUi5DtRKiKJ06xE1vCYSZH6bJwA+Fa6YPeO
M8BMlV+32K9cKkutBJcaSStrtWZWLk8AFMcbKjUdxtKk4HTVvfScrylpHMRy7lmq
gvE1BMCJhm9q29eyYNyy6117+Ybe4rEg0h8vNOb281HXuGpDXpD7kYyPS2epvxVq
TiaFJU2aDPVk+lrGSuSWE+WpICTKpPrV1FUU7Q2rOoeG0teN3lNvNlWGV7eB9JcS
QbynnGDXBF3VybVCbZarI9ui60KAhuAQjJXDM1XWl3AHvpjyBuB9jyAyCwrFaFkA
OzU5r7gsssfDe/9qdfukZ1WWgwU007EEDnyTIb2JTWZlaqPpx8WYCGvKku2F+xGF
PnAL6TKjlvOooxyWlP/Axcbnf5yRSbLqsV+CeKhhjKi5ZLjRqsH5rwaLxFCQlXpt
xZBzBvdZfdlZPLnbDu/pC+0CLNe1y5StGuZBJ7kC51eob2+YX/BwmtrXOtAjULHc
10jskzT9q5hh2r/fwfSgb03o0hN6nXrtBdu/Wh8fbcA5ObYy1cE+4qN5CPvuSCHA
bUMcOKUwBavZWnr3VCWmT1UCD+jvhRli0FkkK0cZ8++IeWikBMsuGaqkyEcvshFC
l+Atz0jgTyV74Hb02TK5vVo4PfuGE5YdpzG5itxg/mJpX0uQh6PbAfr6o78JEwSK
gW0G2nrj/TL8j1uNRqs69dVZmBPaQ4iiKqFgFGQL40GP1R9f2m68JgY87ALW8fnC
DnszwYsn6ovXK4WixAWGlevvlBX6okbN1ayD89YUU3DOhrixm6eNsvd/IRHvslve
I401g6F3qHAJi+4xh4eXncQa1gr0aRQ/syBtzZncAJx3xFPJ5Ioe9QOHnmfH9EGp
Tr9CKhLt5juZNpXvsP6IbxbbLZ3snlzZTw5nf3QcUumgmJNfqMW50yB3U9pVNfOC
Xvu1k2fnSBhHASLwb+b1q6XRTgthgqqEd/dEDRe+M1ncux0BDEa30TGH/bIq6FIH
FubDkXK8NJPPxvyE3uTmGoHuh1Wxpu5olQcXyKAs6ozTDkHEc8ELTowsdBkLkY13
9FMHoPwhOkdZoBb7zmcD1wVYI/ulQaI7H3juVwMEWFsSRotRVjeBNE1P036ST4tG
KKDWpEYq5RrSTEGKzBWp7d4O6Ox1D2GUl3QkcDEw1tzx7tjIlkNFGXIgxTQyJQfi
YVa2JOD51/yPsqeewvQvXY2w6hqrjOkqMJpTjDhWOg8v7srqJZfXlRhdHLLJnY6S
B+j8Skvcuwgr4ZZSwYMw+/ovuuJ8YjrugrD+xn54GTXAkM6XkIkrFLO9FZ7hKBHV
A86HNu2Ruwdbd63m24mAXTHL7snhbUwi+Vt6M5zzNYdl4aDBYrgz0kVrYP7sSIM7
6r+f+t0ccrTO3PMLCJ4Ne7GuPNz3DR5efejsh8bAoSK0oK7RFnU1pjjsDEu8OCfV
rq8T3Xvjtd00NI5YGSYgqtXwWMcYM06Pc/3moZko1OfjymjWZqCIzQYdDobQrfw/
6zVv3NJKSUkh+smnbo2SAE//6T9HqZKZGyI8NdK6+IEIpl4ajTHPhip0PCn69PwH
jKCiRnPAZtH3lVuP8zhwTROimTIeEqCnth5O8QwPBIpaMdJd0e8u9B+lDUSrFInY
y2CNF0ao+o7foB2bLQZdC5tVtgdJIxqmd/mlVCZZeP1/GDLtX3dSvuvMKl1LoTIw
//Y+LS/JqHSXClPdFpO/LrWbEzluOGGbqRBY8hui6uJWjWRxz8phn47A9w1Msp0E
a+HNunFORCcvmIpFY2KnuPlmjRdSCgyGOsHLKv54+2RgeB/tNSVocHQxgQclq36d
tBHJ03TsIIQkRHDW1b8V3B5hu8WdTWjYll5exeg4OyjKvTZu6iyJ+olTF04GEZA7
gFXC8nptJyH+wgn2qesCFktlXCg9sKSDItc6RfiU+mjrie1CoYscKnzO/sHSxTpB
fvYQ9oLdLqc67/8DisAvqOzDfbAxKrmwqbotWzxKWwm649drh7ZeRQiEHZD5VYn2
mXm6Iu96451EHGzl+3eHHu3mG0oTwcmand5c+3P8/obi7zJx921Nxo80vAQfiRB7
mZ7PZtd0EQzLsDsXerx8+NXzQSmBRCl7de2ldbGPRbPh8a8ENdPtAE7ezZoV7L3Y
Ba9zob8VZTtwNEV4LrDGLQplJ+2+IY8ky5uVZlr1pxmg5R+wNSTdxQwdCBaH4Cc6
DYY5ruiAfbNb9UWZyQHekHJ+NlTvZUhUeQ5k64z0GWlZo2rXbc37xWA7YISMmU5N
e6ZPwgXeI/yC9V/mcxw5gJrYKQZ3jEj5wbVAx9vEUgZwuxnprV/kEmbf+IQezQbL
x1jSSQ++B4dOE8ETzFZoJ/SrIUq45SZkhSAvP0M/CPOZdo4n4XYkYeOg7ZtrGEqr
WEC7XthG4UrvCH2Rh9brxZ2TSzyKw3qAX87WsRIzuLh9pJzt/FPyIXTMZJnKsMvu
w0rJTJqYx3Muo13JcO+gtB1nd9KFVX+Y/91sSv8gBBMpH0GxM6CP+B1Egaj9IxoW
YaqNguVs7SgtP6sWC0wZkQkbSyV0JS3NgWnwt529lkUXJN295VZuf+8fDXY48rsK
h9qfL/WfYcaxRKChqOQp1f3sAqVbAi0On1ot8qclp1pkm5H8gRbb1zjlw3SxRZll
7X7YrYc38gnKtmObPwq34qXPT0c6f22WZdR1MQLOp1mcDWZ0Epm9XPrmZiMk54uB
xeE+8DqJo5b0jKmnYuLfjCJiwRsX3YiBI6jS2hT+WWNFvFJBceGotQ78PmwiJEww
ucDLyapVn1+JSvXSvLtisaCypHHfu1IBXS9HF/K68r2WXwUoS4zMEiM9ob009Kem
C4M7iEnxJpznnBVDyK1a38vJDx8fnkrd+FP7WvLCD/OOHzUHlxAgxugQaOI7Wsxy
+AHga9GFwzahTqrtmXS8UiblHjQSHjDrNXn6UtJTFWczVn56Puyq5adw1UuGuGjU
0+EHLM92OP16x/cKTS58i8SNqGKYwlJB0fv6+E+PfdBuMIAwa7dE6/NXomXMRipV
/EhnNp4hi+B8xiDQrHUNlQI/qlcg1epChwwxChSol9AI3IfLoqUEiJnkucdkIQOa
jRVwMyTnwozikP+k+Wh3SPWNVBvIm6qAnUNaQnIkjXcggcIBXqovszpWEzfI77NO
gAZHJx4G+ol1DBP1MQDgeAlxsNdkT9USHGpxnmR5cstPlulk3P6RK5ctgQYmwEi7
SSfI6h0zuQwu0bz6iXDsuzIEjfzEplzknI2T06Qo5RdsOdB8IsxBlFVRXWMQC30J
8iVn1e6qdaX+njWA0ulWDW5mEQLMr/6kXgnhXOcixBmDmA2btSHKY3WMBlF+QQMu
i9ahhg0/Se/ma89m0uiYpRoQmfTASbcEVgX7/3r6tGosUVRpz9JTKLkjr9LUrhNd
20V2RwGZUoVpFrAklKDz+GgzVBMMv+DGDAkFQVxHOXU=
`protect end_protected