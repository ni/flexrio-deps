`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6656 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
C+Ri7jmn92TKTC1Pq3whklw3C19ShUGBpB2SNfIcOQmdr9r47HmbE06PvEbbazTJ
dfigw5mnDs8KGkXQDF8kB/OfT4d5uQYN6W/BHkTq8AdieFxNVHeGkcUa8Jz0btfT
ibAwEi8RCRYcfkD9jbrujj7ZGV7OlKDijyHpWr94gX2QKUP4v2n7mB4dtT5zVKxr
1SKYgnZFptQP0wFKHBQXlKXWBMeEyd8Yq6nyhpJ9k25Z8tD50LXTamGVKqYUYRgu
LZb5yKrqVt97Herxy9osnnRuPBeJn7gJuQF8np8QdlfhTWDTQa9TmqT/QnkLioua
QRRw9w0qEeko8aVc0cZ7d+in12+UqDcblvZeTNyuYIZBSzINbGJyXrvSPUyH/GOq
k2C4Fs/91Z1RE2oKCq432qbt1FNFAbpa1Mg/mc0Emhel3mdOxNodPTd+T32yMmX5
yBenOnBQKmX3ewCe2DPWHPoJxZaropKpgZZHQwtHWTtHD4FvebEm65f1nn5Ds5lA
x/Tb3btxxOIjZJQFYC7GRmr+uFWYus+TPFdUWSB4upNIXOjnaip6scaC5VJIxbXw
kwnrYj8heJqx+etQiMnIhnBv5RmcBjSJuPcCx87N0eNDTXkOOuo9sgN4A173IpNu
cU6OWTTBYupuRRQjacgKwH6vMYSthXKI7aW3Tw44sTN92keEmEk02aT3OfxRkhMe
YiEvfBFy6jRNRJXnipRQjtxYUAq0Qf2/WPameHCwDfcPCB4BaaOqHRsqrue/wifD
rmgQiiaR7cEztRTuOjKrgLhmrBPLlGVh0uqgnyVF4yhZ/EFnGNtwLUZC4Mvj0Sx7
pKUeG7SodCO0waNgiWoximrnBPhwdkuVUNsHZiwK99Ai5y7zV5fKrx2+HiV/XTKg
k4DAn2wrHpcYIp39jLaHYQT9LZNZbSL+UE/xLdNssdJCE1bN9v1D6Jqih+99SvEm
utn/CF3qz59DDP90lKJK3vAJmDin82nt8IBtHRQdJ7j3xMIsiFXQQ6co2TH+Tp4L
bDTxz4PsllewZ+uVLDXX0bSXZUhSEU/IWFOVEoTKCd+gUFlgYVnXJlE2a0/EcXhc
jqlzFb502R+WAYa1YLgP05DASDUMkz79wsHoHOkD/8IAo7+A7eelmJBxBdbMcXCN
ILm7M8al47GPc1Sd9Mi22ncG+WrEiM3tvldiXAh4dY/14nSriAqH3iDEQuJxEKWA
gKfMDfdf1P7pLLdu8dYxiqXx7UjLyk6NzNBMwyNC0gOYp4dVQZ0CdQM6mQ0QJNTy
KMPq7Jn/rK0liX1QsKxeXp++fp7om2vpR6cMVr14PVFqe4SD8oDH0eJHvSXTPOSM
e38fcXYdv6TIriBW2aZvAQCw5KdPj71l0tSnV6ZwM1/wQKFmIGQxPstbD5dTE2dz
NePQajuGx5hxMn6euxlaKcIO+wJUM02UidNv31MKfZNUkKoqKDQjvQ2hKmhPo4qQ
zjHQi1uEvNXWKPxHJ3FXRzizIjN9Mf/tlR6j602ucLQ8omrTXfkA8KJYW5eZB/C4
WlTsrf62jTxqCdbqY5ktnG7sWlsrBBM8nJGTE6zlNhvqlzqR47MGbyoHGs7ITSGY
/VJ7yl32wSgqPE9v0JmN7vtRG5ziEsj4emOTJlkCH7w/Wf5SZHFdu6ag4gh3x9Id
4yTj6yebueRNOcZXihJ9LhIp8mbnIsfshwgqw0PZKY4+VqMPXsYU4BYqdJ6gnKlp
qtYO/Xu23Tj9DIirvB8dRHHnIkFQw/A2Tbhti//uWAqQEn2tRAexgj2WnVw4+6QT
ZodV+X+jfhmGQM2cKM1b8z01cEx6dQVSXntAwanOpbHIZJlDIZWcHY0F4/a8f/bx
w7MFgdgft6eJtqot6kRvwbOOWdjIjqT+mS5mv/19w0KYAEP5rSMTR2exUJPApAvG
GHBhX6m9rMZZ2I7bmObkwcGPPRnXfXGqLT03qkTy75oWCDjCfSDphT58RLQVmxK3
68EnKcZr9X0Bs3pqq5NrtebVAZNOCbPmxZuZQZNsllhHREP065ofHIU6F7oFHz9Z
cXifoZVucew1pHcc19BSv2/ZJcNjWnEWI9w6w97Lruz20mZeHke4a/pVtzNw/zyV
hvd2Rc6borF3HRfa0ZRm5aUKlzn9fNMl2uyWPlW7llmCMHtwnr8SmUZ2IZGs10ap
u+0uVVYLmpG9z1ydW8nRSPzBR5yUGwflBVxPnN9apPXypSG+AYx43OY7c+gYLW/J
tpIZpOLHt8gIvFD9N6Mk8Eqq94m7XYHoxso9Y3WmL2KzSeUx9/Akaz2eS/2orItY
TGMXXupZrPqARjqoMpSNj3H2oyY1J7YZoo2kxC1tZ7ZW3okgvPr8MRkxfRaL56sP
x+IQawShrFklvyWwx0pADliDUjIhtdf327GkwOmH6OTTWVgfLbfvVoj9qJS10BWj
ieLE2BTTXosiPkFbEPWo/WiQeQ4cn0s1fAv/bcayaEbPyXy+3lKBwFbbpEZHKfb5
oamIXz8DFd5jBJM9fLNCkYwbVFXKkKGyJoneeroMaEkzTOg2Nif3W0tMjMiNfmKG
thIG4G+7US/b/7qpph0VuPw98AVF21zgFW0d77Xzzmq2D/KQTPyVEu41cJR2WkyK
/24sIVtdqxvhxedbrHSkwqe7fSx6UkV5bpSuTnHt2C31FKOSGwACKtFhP6nwhkkv
k2HcrM4Ccq0xC66Sv0JRbZAbH/+IXm1/Szb754OrLx+rDCBO1dQ34dJrKtYJ8wnH
YjWmffs4/U3DxV59OaKSxmYYFqffcYNU9svyiem8fcV7MdlYEJ1lwOx/ItBOmY7g
1OngreImLb2IuOea+zIu/1XBjWxlRB6m9j/x+eETh05aW8OajvSQxiGoMjMp98s8
6VwmpIup6/ISRIPs+LjKqOkgZfW8/hoOphhVu8FFWXQrfAoF9i+81AiOFvKrgO+J
h3su+hN9bWyzp4oIIFoGwhRRFMzefP6t0Aw/fD6SnHO+dHl2dUPvGtQIo2dWjba1
CLqZBaDOnNaAavNZCNmbRPN6pCnkRgdfJ8IVR86yB8MNg63XEQDg4+xCVoBG6FNm
PBKZgwiNUOVOIXgfNo9hStxtYILDMGUmzLKygo0zhYoQ+PWW9APuZ9V2wuty3a19
1kuUHVhMskvZcT1sqoHx7RRQQDvpXNIxmwiRxUyK4YM58F1EeGq75iqjuqMmqiBL
zFeBWZN9M4pDBemncxr+GZHShFJyro/vmGvzh/IJR4DMgJPyZ8ORoReFRxrgayEq
jOJ1JWptnlZKL2y9aMDaoRVFr12Pcnth8fcvBzkeyKuI+t3dLpdCH4wDiq8Yupqt
pSvWiuoPPixlL8tSRQlRLCZDvACEhj0N0x8CvUV1uUEfq9cmXt/Tbiee2/I7DxSK
78N7Psy6nmXafmtyL3ix3EkBT/CotUNLVJBM7UO78ZG1patWPcJsAuVv7vbN20o1
8IrPK0AfA1RB2dF+W4Zued4dol8Nj0ZB5PfrEO/Mdgnz35fR1iV7YDMkItvPoPuc
DSpqCmLaI7Fm1n0YzbV+9Ga/9tEAGoH+rje3QjJ8WzYyqCFuihr6ZOpUGpnI54rZ
qVrRu/8ZPQScFr3v+gX++sfzZTjyLRZYWy3BfCLSPvAtO2nIFE9aeAnXXI37aYdu
ETUeZWS8t5chEWKT5Kqq874Idx1JS4NS1ZZumB42ipTQbTxMqsshYDeDFDt2GEtV
FjeG5WEVXeJZNp+t/+XkF/TTurRIxNUwsx4R0tRYhEkLZS4ZG2V4krx+e6DwDnVE
7WwS7OpS3p6+6P5J+LMST6dPXMgQP9Vr4K+IBnmdz9Pupqw3U0gBLYsW7FpcunDy
9ZkMwb5hHfILbLNzWAqk19SLISx0VwMPDRVWVs0VICDiF1RKKpRm0Pzpw+eU1/h2
LzNxP5n1visD7uetbtb1d2Zva30s/sdeJnmoI6vVmxrr1Sf8zgN5E+aKQthJ47Ar
f+P6emGFmdG9TnOVRzdZ5X7eUxyrY1+TUPTFHRkrN/H6/16HQ1Lj2q2vhO+K1/bp
tWhunnQzlQ5+fbFV356sytG9YfzwUCDb0lVuG/OEDsl1ZSiCGIBIAkVrp+6gkr8p
UlLAK6acqT6JIG57U3Krvojvwl3crw54mztsslTx9rOlUlGvltTwYW/ruMYmP9eU
HFnnvk8pV4a5AA3PIcBk26aREP1yye5lnQX69TS/mFbe9HFlnf1k0jFJ22QMIqZm
mhpb1g0mRzkQL3UonYqlAxFud9jMM3/aH99RzTntbutRSfa1wCHAXefsOH/ZbbHB
NOTd4L9/F0TxKG90+5R8HiVxJq48QSfnCli0X9dYcIbFH62RjLYkzZ6cjm4NfONu
cPS8q2SnFF7fXnVLOVCTcZmprA7Pvv0pZSPXLfk+l3gYzgxGZPj2Iee2v/ruQrx7
NL87+HDfHYgQ0mMXzdxN9kN9wwDFO5Y4U78ODMRH1Jf3FQOaKin8a9K5OxgXN3+A
Pq1ruvna+1kD25HndocU35RB66fT2FyiQSIY+SdwymOnHSXXRTb+bB3DG5czBEvv
WiUtE9BaA0GZVuGqJxN8Sz9vQdVaaOyqOsSYbqWcu1lyEs/vQ0ahQlkGH9LeKU3/
6ZM+1qpZBOn2ebTpdnIcyTjH4jdHJk8HeOCPFsSxzJDX/FpWf9z9TRg3vm+AoEOI
/NykOPQq6SWXrXZvmy+Nu5lY6a7cgYJ+4HjwMqkNK5nZJNfCCQiFABQjsdrZHLWi
lQClNUtfhknNr/4Yw1QS4Gt3jBAb5/2P4ZE10PJ5LqD4l2wSPCOF/Gt+096uo12X
grQDsie7uc3jEMoRQ5gRpN7jSXXdrPuabc8ecuW8OTiaoLdGX+cyObKYlZ4w+r9X
9/aQxEgeozz8u+A9O5+bFw23UZMyt1d5UUhxdQ5aAfQepuyXcCgobj/6TzeEFaM8
ireD/E6wd68oQy7W70f3DJQBVxvGH7TKwM6eBMMsL0OHiH/ilQVSfAay7kl8LaVt
DykfBVah8Z5JejypKdfOLxwTN1KE3ad52TPEvnIRpbL5NYY954NuY8hJUJr6B1Hl
sRwPQ05ni/xm3zZlIB7ZH2/tQ3Ul1RkCdy8zdhmmuGQKuj+rrpTEjwXL01AN0jWS
q2x6bsWjZ4CwZUGOYOxTRM9M8NiwSlV4T9Kg2tdUfj6ZqesWhCtHRZgzb4KBwhOP
0i9jAFuN4oZzqcskp7DLk2JDwqDRRX4vOjp1c7ZboWClZG++btvTcM0FCt4j2+T7
3TWn8Ith1dWpWN+xo8Gku5kszr8VqBPLXSNnVGiwAU8Np5nmYxPhxJ3c4WXNupvE
LOz8Yk1qad9EfV7hwV3f2svOS8sblZ0dJW6ZuTN2o5UOqBED2aXOB23tJOvKdoRy
JC/YZv5zzVBlhXGtfdo/YJWe1gnn2+ZN8kuCXhJMpJILKbIUogT7RzMyfyEjIx61
EO3LGPyGixdz+LNvHavLENC/dRQU+CZCpJ5XZbvTiq6sR1XjyquCamJc2A05wk5/
VZay4gxjw8bmERywZdJObjGHRkBtOI3Rt0JmjwkiTCmUYGgyugWwNxK/fO6bmWbe
AeT1Rpe34+2bIcgY3giUg0EiRv94rmHX086mIe4ELLz7/QHs+cdjMHW/RCEx3goP
98WcSrkm6WoP09XQVupDgqa26ML9eI7J5mVClLkbsvE/SqbaR4BJ5Q3lHcTRGesB
+sQdRI43Pu1fVdBgpOihQDSmmwVoaA+ih7GbgZrwO5MDMwLcL++0FmdVeZg8LDHX
0L6c0B0ix+4BPqjCTiHNBn1MYtNXqGx3DLvQhcMXOFggBGLcdjfZIRNO/+E3mNxQ
pp0L72wr9pJihIeZwiNlF9Fl02YpEaomQB6XkfpyBz3b4qNtAfJcc6xu4bO6Hu1h
Q/JK4BBCuu44J/aOsQ+uWQycgI9ciSgqOFOG903Os/PwgdK+DBEl2MTIjDSYFZPK
R5heSdAjviqlaqnlUm+TTHwu990YRAopaujS7BvyJpBiaz6eRO4DuixtetMWByMn
kTf1OiqVLCOTqhFmTNZ7LVNG1JrJKfrYsGTcILIx0bLrEmZKNQfV1KCKrsQMD8/U
q+8oS5F9vnLM98Skw4MNBEMvtmDcydXurchWZktCyaUSu/abKtdXV3w/EtfKLDnI
VdPm7gNkjNr9Dl8O+zt+7A9xDg74V2C0mE+xJRMIk+Ull9BEOibU8nA3+skifNof
K2qhLta7WQlNslmnpc9kl4xadsQLgPMqNZ3rQMcinZ92VT7jmbvAyjzMHxXxTrSE
FQ2XFjO40KDKkiCT2eM+vMyYMGWgM3pZXqbJjfGFORzXx8b6GHMwFaHPCixBLpoG
6cHxrR1iA1aj4fO/8E3astKWElJj01h20XTQWA6QJsulMH57byGMAiQXx6zp6UHE
sqh99xNqLDYPajgh1mHioZri7HEsSB8xZx7sj/qQOuosh48yOmQiuQLeSHVe1y4T
vV8aD/cwXJDlrRZYslqmKGp4yE5yiVvyQiYGb62z7XcCPYsMf6I6sTzNe/yQO7hK
kLwyZ3fGn4mlIcSQU1y58YmrEryJ03u1fdSa438mQxIP5AP3n6lo2VsEAkM/6QlO
O4yrCXdxph1JiOQXkZsvRngzu868iuclRnyGvB9G6zo7axBpqndmfZBqP8/yBiKm
v8Cv7rKWcsX7ttqYaztB+fNjT5D76JUfiv+9/IGv8heOc5EtOdKoVS0dc8zkRFQR
IhI07ts44Q3HRZ/KR/1NxoBOHEJDWwirvPMWewumvTQJ8PVuCI653f2mFcs6t5J+
2+Ja/ADNM9vQd1Nlvmq0VF+lNbqATqpCquMsqXNrC/YV/Yh3m9WzuQDpnuKXowlC
L18AU95VmQGVssa+7npAOutCTCNa8QRBjcqPQsnqpmmUh0PZT4zFEs/Fq2AtKobu
oy+JFvEo10QfkDQPrDYW3Mi3FRHAeKj1hKm7UTkNOJRqyjRDF1lWIoOdrKJQqEhb
g++yQnDLoxyTpos5X8o3P+SZP97BiGyIYottcWE85/0MHTWZdtwJ2rp5sJ6t7tfd
b0rUJlnWe3RoEkjAgByViSFuSoDUnGoNLMWmHsW8e5CwS2KscSu7ZCVR3K7/Rdwm
eudI0Zg1cqU3Hip5Psd1AlfnsQkW/0TRY10pPcGowHN3PsVHjgHVrkQWFabyQ/dK
BZFQHO97KJ2oGH3gZmGF/d5X805i1o8ct8Wf9hN4nbSodB3+/UwyQTVahn0WDfkh
cS8p4dLZqMz7PtVg6M+c2Brf3TyPXZX+DkDjVhx114FVDpjBX4df3R7APR1jACng
4E+/pGibbfbzQOgeVJlVT89l6Z86ueo8OBPIjeVgcNKMXdARuJS4fodNHpEfEVPV
oNXElSAg7B6bRBA/rjNFp+ofki1pdbKqf1AXIg5LhKQsj1zQm6vAi0kOblc7qhuK
C2FyhRl6GkLy7TWu9yxZInGvNbh9Sz7QFPh2muDF63QPUl+sUtlxKqgmdmNV/Svk
vpzNizNo4JbS1xngX2wv0QmJvHvHOC57tWMZLXGB88v3YzWnTqPROwk3vhNaHqVk
8o/r67e+5AEeR2n0IwXBoULUXIG/AQQkksLBlWg5dAjx2//mY0ndH8LSIlw7yxMg
2jwEOv58Mo/8v4PSkRwlG3QREG8m0wYLbafSqkahRbAB+ZH8JPegiq3+cmGTEmFj
OOFY13/JrJ2mNVTpCwd8itwSq6Hl9LEzzBJy7+6FYRxxQoGf8l2Zpmof7DU6FPab
T1n9Otsm8J6kXt0bZvVHSMCKRUNZwXSUp01ubkVEtdPenRu4Or8BGFQG1f+/IydV
ZNCiWX+8xwCLGlFUOSWp9cY+d1z/XYNBNpHDdE+eXIR0GLNH5QWPwEJ1XEMtBzK7
lWlZRBT6dg35LzeEe3Kc/uMht/vnhE0ehj9ayDTrrMZXCRmYnapWtEkQLg7yavFL
31k1HY3v+0DlQh0MyECApNBfJJLiYlm1iwi+I96/t8hinO3go4SqUEi7OWF3Cj6W
Uq88uDmzaC3U/h4ZO3jId9bwQ4OsLUlBFUPtQ/lzNdiHM8t1YVHw4DiDjoxC5lEl
MJ+OYkLVwbi/OSipQq8KDLelCXr/rp3EkvsrizKNi4RCfWNvbvpyod5O9X6dNv2r
V6kW2LoQaCiQAiCfwycpr8Gf0I3epl0Hlqqq62YFq93XRUeZLtMCFpR4i0IikJOV
90WQkdskRrTVnx47/Jea9bRoSDN/Of2AalQLipnGKpk/QvVDjCy+OsRvHb6Q9VWa
jqapKPQbB/OstaCq+HV7CrS2gvqx4TDyzYvG2RUi+QvLDa98tgRC2sGCaKCR+HC5
EZTFnMGrhN46sy2xXaO4Tt3BbWVzAnM/DAo+btDrqEXqXSp0lSpgfSDn4ZNfHalM
HcevU54iVzr4k83eBcHJrSysaQvdkLh+XmDCw/KxbWh2CtW/Fp6CB58D6HexrnY7
Ot10rdzJC20GyC0AvzIijQfXHzijhZR+mb93vHKq6/03pxrhp+5NxiJIAK/C1XD3
rw41B4AOmkG/XLQiF0lvseqB2ZxSoAINhwvnOduu12yW5+AMnqOQmOoULPqLzFtM
o+Wt2H72YVFFZjhgi5TwR2MgMEOEIowtuyhfFyLV6C+24dI1LBvi1wXA2H3QZDAA
N8u3f39+/PRyKdRES/DFQAIJFtZ/9X4DFW1PweIZ+40Esk9bBUwicdLf88l4LU5q
6Tk44lDuLZWpvn/qzOgCDC3PHsh2k3xad4fx4o0Ekgk=
`protect end_protected