`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12064 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
lmOQgIOM5jiJrGbWpsW/8q2c22QVGMe7FjboMpP3FJ7jpICQXeVqG6ImT6jXSEqv
950UCnpQF9anHYCGLezhLucdVpxC6p6R7yVU19tg51BVIMp7mh5nrwmH1qbgNack
mQEipqPGlHrUftmi3qvDavBDY70NeIsJHbA3oFBLPD0AAwD93wipGzpTvAAZUT//
Yf8k4FgL85CXdrWwbgc3EqQiUjm3gNtTJuUPiE57pMohH09s+b5jOIo7kVTa0rhC
PBoHrFoR2YGNRmLvivBket/BpMGCo4sZ7vzvJ3JmNged/9wDwIreVjqo/0+EZIqZ
v1ub1dA+Y4YsQQvuhY+NvuKOKvAE9KOOWmpWDEUfaf9afR9Zp4nFzUhkGAf5hwEs
pCUs2X1ej/VZM+SnS49SSBUGlo7YhQJXVgUe1rQbJCVHnp1tZxvcZ44p6mWoDnKN
Q4OEMP6CL5ZG6Wdj1RoONbqntaaB/7AG8aobLKbhnFJpL59bS0W2WOZsdzo8KJIk
U2OboQyRAWHkFo4RmgGU+Cdj6X05J0dmkALBXClHz06t25AEY9hmTgsB96vnH/Uw
D15JSSoPoGzYB5y8geVqzq0KmshVUzhvGNEPIjlO0IcfEYzlS4WnS6PUgoLfYeJ5
u3bwG/KSOuIXACi2YcoYxavTkwnlmW14/1fWyW7pUsWOhhQtZEMxc6t1nq0qBrml
unbcBsGchyVIi7SCOFM4ypMoIUJpXg+7rLiQN0pBFlbLtmgL95xJbCN4j3IBiC+D
kAkWsRp+EmDROG2sPyPKnRhD5rRwcWBvYjgR0+V6tq1Bcjosslegk4mX9Wno27TJ
yy0DbFz7LnUkO0SISYf4owkZbFuw3/4G92I31tFHdDjc46JtYnegVt7guFDxSvWK
71Jj/e6sKoKSala2+IiRKJCqYbFDJ0itHQbtWwAC3oBtsrEh98Q273j63ft7tPs4
R6oys15lioPPuqqz4KhXf9hzwcB5Pdt651uKa8jtq+2WfULF5cLWRa2a1+Y3E4d1
RPcHRA1r+wFAaWB8hVdrIQbblEaVw8bLP1L2MZwTwn7gMVaj7nqmqfDCF8VGSVWA
SQwpLSG75ndcRDgZG75nShYhgZeDmPdyGkc4Liq5F4e54CbpeOMi7MbDWwCMcIwO
ggVqq8+DImPjIKtRD8/jO4vo8FSXBcxNi0Q3NODOqqBH4K6ZcBx3OqbeQ/DmTbgD
qmgGzvkc+bnAfDWr71q5yvNEit0y0Dts3uvpcg5mVytOMVYXHf010TD3orxlmnXB
mXtnwWm2fFW9XUyyrD06apmZOWjxczVwKQ5DKAEgKTOuRYoW8PKri99HkH4+1D/P
9zXc9Z495Z7Eg6E0nKuyVOV0+rUVg9FIgyPT/UxxJfneTFlb6MfIRi7y2WerwjMD
OthG6AkVfnJv5pKS0UBlI5JJMp7yOu9zXXMd5kFqoeQxoIFy6cLti1BDhWvsw95j
GxVQIuuxqrXex3cEs2F+n/T9FVZlMDrfoX7Z18IEtjFon+2j0rD19KW+mVbezSeB
UjjePDLYSmeKhY4S0vUUX4oqabelpa1SnpjiDx8cqaxLLX2RBikaMYf87pqW4rxa
YhDZn1OxSl781GRoOUIF8RjDiteedc5LwC30YFWsS/01gPT526UFVkYI8KA11pj2
CPxp4Rdfr7SCmHkHenKoHRrobWY3M6vSkqN2nUFEBLMcyujetKoajayg/F4/iT93
RNg7InD+Rr8yGics1pmNEna9RbQ3IFdB37XiWAs+xP2hDebChu7PmmDDPvLSEQ+R
4ePp8g6nXAzAqDVWRAGuxhYHrBhLbNC62uGaeBq9ooz7gCRBG4koYx937vfRjhoK
7LCvW4QWJCE4Pp6tI1w3Em9hnys8JjMVuj5NU33JXp8TJBTmxpvwlfQ8Pp4UrTBI
7aXC5itgcVFrgbBGA3O0RxT5j9vtjMt2mFIKqKGrSzb4glQjO2nwJrc/LP6Vd2KG
pehDu2ENYW1NpJb6jotaNTFg4T5tyQweyK0TBICE/a/kXNJSbNe1reWNHFr608O3
B6INaONRHNDoE7mngwaWOqeSaeJer2wLbtOnO9hsJfBXLLxOsGLsqvgTbP369xsE
oeL2RfwYPOa3M4laTHfZ5p3qntd+Up0o9AGkPpjjbV3r2fyTbc8cU3ffouftRnWK
hQgIcYSEEDfI2EpbmdtNkl1t8NoyfgIm6kZPLw/lmbCkhrFkSBZrnuyXbVx63nIi
umKpdFplnhRRiXZ/bcA4InNMY+aGFue81a7h2LcgczBHIiUvjHfP3UbCziEMCiKr
d6co4vfzhzf9uqejNnR0cub3kGDaZNheQFCucY323rOCQKIhg9AZmnnpMFh5Lwyc
rUTxleOfEYIOUYIS6jaNmlHA8XGUtBsN4gPbtV6u3b3gMbITXCTR/ksvTjq4lM7C
rk6wSPeDsd2dfEE3wUa0DItNIgYPO54WqhBvc70AjQX3e6mBwGwTMuqX0fxAJlVC
nT7cVL7CIqm38uEDuGoQ/njN6P/CpQICirL3tBjilP17vxpEiRwCG3KA0HyTl2Gr
AtJpbQvoooVX7QdOG05RkOdfu0lX1VVftRv/xghL7+oQ1+upmqSH8iweNbiTKA5i
kvtFlJDdWZ4nA4KRtmoVi/3x69191krHMC+Z3JrAlDDsBOUbAj5QdsFdvBBTrf2S
fpQQ8BKe6k/9jIZ+ExuNmfawx4zpvTWYrdqEHJ4oG7VXVOnBtPI6EUVnfJBWxcKU
/9jDZ6veZzac3iMoOuoBzNzZ/IMw1jXHc9wUgeOb9grEQhrcmNFVTf41uAxYaY/S
CBkjPAo94WzXRqBlwGi9ZvevOpMA2Z5qElih1oakeZw7WZ7T4mBu04jl+Pc24BGg
L27896Py74pFO+C1sqnBrx5+u/KfH2I77hwrPSQmYH8DxKYOFaAGksQzJNVXqVdK
MRrhynA1R1uTjTN0UP/mFXoNgsVcUADF9vxYGqnWGQ/6SbA+2pDSuiCa2N9glPDp
xZEEU+4xxTGdqV1p32aA8xkhuSubVsM05koXBWhGKyYBJNMZfBBsVLHeH+vjxWbo
FuyIZkOx3l9H62oEkRsG52+2f594s5tDVpq4JOXHIcKNueGEO5t5Ca+nOwbBsCG2
iJz31C6qkYuBPYqPDuLoIC30YdxVYf5hiBgtebEjesQkIs8H+jvNxo6u9k95bjZ9
3Dn0Q63IZztzby7OGuwugBINm7oDHDQSCSVDIVIeGeDkNvivh0FseByloMAHJInI
NGrZYpEjeKUgNFnYpC4NPXl11T4ckJiLt+O2sQS2gxGchdVwF1Yczf4ipCSmh+fk
YbrQxSamJrsSDmgEu5XL00SErA3jOW/eJ477gYjK4yz48LxzP8YSlVIxQhuyBmzw
mQzw5qczF4rzzkahOVuUz49y04g38A0wHaBSsnKOUAlGAp/Ql20JUtgG+CeK6OrQ
6N53lFGURhZkYjbJ3Tvio8iNqX6YOTeoS/Nuc2pWSiiJKN5DPi5LxB/wtb4oMmO7
lmw9cUaPnLHR2gfQxCVZqB9RL3HWecfasSMUHQbAEfWDCn/w+Dm7IoUWTXrhAL+8
I4uTbSvRmemW1F1bj721HOuZLFGDhUVqvkncMw06UhgHWA97dxPAWCDDiaujZimP
LAhKaXt/02OZvpjUfRpw5MazGB2jMmA9Tyow6HnKeqNPyplfAYuyOZ9MtAN9CSVR
LdQfQHcvvioaeJAMnifUI+qRdCeDQ9wnIaFaGT24FbfFPdrGYMH0Eoui3E8MvavT
ucH/4BTcV5SP0u0cpNUBqNcn7uu+2DQqGw9mVJRcKW1J8SZl16C16+K90qn90/Ex
WCztrt0W9QvY4qkYaamPaQdpW2U4bZsvXhiO/jTlCaFZ6P2ah3OWlWb6DD3bQLTb
23YR/fABqmuDpCSl86BuXvBdgYs85RSiT6OzbfFpRm6A+BY1aAbBr/xBlATuMsvt
IYz0T5sVBUwWYEvnF/eD82ZkxWbmHW+i/tPyIZ73AoXVFk3vJepZD040N69duCPC
WOxQx4T5DKQkSUTFS7qgIh9CvMcC20Lz1i9o1yRz0W3yX53jj5kuOk5oSjuMgTGV
ifqW0Q3iG7tTrZk1FiMCNcM6UAFpEed2NuO/Vp6aY6yKAMIMyAVvJiRGi3xayid+
4L7mgv3mboKFjgEY8sbyfts3CL6osx1rgbryDAyk0fSAjKngV5iijOmCJBORtXyh
QHyQUZDnaa5E3v4GpzjKPXBxdOkkNbqAst65iPHbgNTeHP+HEroDKgEi/hHQ6n0i
OZRrOLqYkF1cW8Pkxhk9UJuso1sHnKklmzxXLXZ4ge0CmW0uxEJYbr4f6vewAKK9
QIjVVo9zcArvFLwrG4HM0WkxrVpI6pBaZ777eb02MYLV3VGtjMXJ97lkxbmjAIks
BbXoiEhi5xQjDkuoETFg81hKCyRha/ls7LyMOccERMrxi9BSYDHU1eMCRrZhUXhr
LGA+H90qUllGUEZ7SAIdG+dh3tkFJhrjXICni6CvVSdhwW6HzutGiVHqD+tQjjdj
06nO4azHkerCWeXvXwMVypwR0lLQlpCsECr9jWEVeeVfS98VUJxBDpwpmZFuDB0I
KNfz1M+x3524NWPJZVRxyN0/XY0Yz5n6gZm+x504yZ9PKBnNg2V1gw6j0FWKwJqH
tKWXCTrtB0gm97dwagG/1aeY2TNBad1XJSG4NIWE2sTga+EyBvrk/I/jZqmx+zZu
gtXob8ovAghDeZHGi1Jg1mZegUkrjoNDy99HVe2Ge0tGmvRfS2YU81bYjN8aZGhF
Yc0b28OFnbJMpMjsA4FjUdHFVV6cxVeOrPVSjD4P7qbzeB1Rvlc7tFTLRQ5Rf3De
I7iMnoDkA49LmilH3p2AqT8+KSjJXZJb3XftK124xj1iQnz8snVCW/Ha2piz3pT7
jqwjmAiL3VjFPAkZYj65m4H6AltqenxtmWlBm+zzhyahQ8qxu+3MmRPnOWIZEavv
sCssWJ6yUWku7iNzVYLEz6zmyy5qUzXVLPk2p7tlWVImaFaUOOKYzfbf8Xjp1loD
sMJMKLUY61gplvYkgcwt4TFJq3h0K083thXKOEn/WgZxY2BQumyNBoRe4cCpTV8r
ASpoijuUhq5FZLO8ImrEehB4+QH9fL4OKXyrZ1tz2JNHItJNgpH84I7gQBNbZsgR
wSl6aphz6toPUHtWc7zENI3qjoW2mnJbMAfSI5tVDMaVRK4aNt/nNLWpGScG1nWE
/F9JkJC1r4Fcz5y7rxNzF1P9wabwToemOgav+6Bv6WQ39tlRUs9QxVX0It2xMkR7
IcmjNao7T9hz8gPlJrBSu0XYCG2QQ6t5V2dGyN2y/94ypWL3G9QeP69RK5zbqGxJ
Xn0495TUtcDrHFRUbEdN7T5o+zLWUMybrmYu/xq/ops84kRXZG3xxyksWgkx1po2
ykm5SR9tmuXEhrcpZlJPRO0Kv0GyTjE5JSmuqhLYWAz4B28VATfnWqlDSSfajTyz
iPxJnRKmsWoBp8cWcDrh+R3HCcf61N6QWPw6duAZdXvdN+VU19pw4y6gqgu8UdFb
LiqxpiC+OzNeT3Wqe1+80L16MOkL/oi6XctI1KZMbh+Z5iTdUQtMkypQDceLehXY
+2VCBmw9SqQqJLj3xdKUUBOJPNikUBYiVIhFGSTDrdOLOiCI2S8Ove2CpA9gEkWo
shQ7bX8iR5OaODR6N8CUZYDMYNfPBu08wreNX6r8ZpywGK9q2NRVpje07On8WPBD
l1roIXOgIAzDprmUQ3SV17FWZkHTyDGwkj6vRW50I3vN5puIViwPNRvuVvU1P/SH
A+uP0rbRQ8MwQuVc0OYEyuQX4InQDyJakkBglP5M77v3DXJWYIpI8kW1i64a4d/w
oog2DyIUa7JbI0VdyWV2IdChfQ105s/oX7LdgEwSd7oL7pC/AWWzOaemvH1xa1q0
UqhFoenF07tzGLQMXSFGqRcSHdwxkR7dlm5FNOGwp3fBXASnViiUvdZjudxeNMWM
RtmxCvEAawYdlnonkeuCZ08W78RCarWbjl7P85dy/I3DEzCOeVTmVVQU00E7d5YH
pUr+qObkYM1lMWKoepzZC1Mq5j5fmnjb5uSrq+sMn40xyTnAxaKxjWH2QV/CTUwq
UgtB6R0e+ls5VEPZaV1XH8EdhQUDozYCJIZh4pK0L9Pstx0RsQF0bsXdPuNzWvRJ
biwNuS/qiejHn3gz0bypULv0TUIeeRE2rPCWFGaVmnr4Gnq74UWWtLX2eLnQuMpw
K4zA1lvV8Fy1JjS61yYdaJHyQJw4pQeQkOPIr7mddv4yfTrOfRg5PS+17Fno8Mvi
zCrOzdR0iWm9Ba1ZfEX4Nb6uVN/e3RBcR5LCbkOCX/gBnIsQ1XsVHFSpzdFo44gj
W4/NIrc5xWAvCXsMD+gmE/j4mtpe5/yquxv9j41yLyfvSv7GEKRWVL7mHt0wdzBP
RdAHW/c40b0d2b3Hume/8P7jbuSuf49UMGkkKbnloftSkSwNZWBPDi4sIMVxVWHl
PAiXdbpBRgZ+eHKb40BLWaKTkldCfYBi3O+AYLekeN3lB7hvPhGJypJNQmCQLwj+
qbC/FhdmFf3ThkxwwziDFG96xefVt1laHKTTgnFnbYSoVbS61XrawCHVJZ4s01yn
QkbnvLjHEOkyuEWSlJc2PLO2+tTyWQuYkw4rqTi9xVw4KkZ8Y24bLm+LJBo7s6YD
NWlO8w1A9pZQcDAYKAedgoYOzBgOmqGjzQ/1bMOMrjOMkadxwBdXXcjAc6t74VNo
/uzvPFyKC8ALZdgi8cnKcu3pI8PMbzqHy5JcXyA1cbb6uduN1sjjvWtqpgwzWAZA
jdFvl6vmxZIJeUJ9TaR3jsHawynTVbqz9ofJ6wLyUhhS17YkybR7ewo++murUz9p
xOyPTl7cUgiozMqWQ3qwwWX29QuQ4MI/eF/hjFEu+r7F4rrxnJ50s9rm4FWB/TYl
TAUMMI+cntJsITk9kwUMUtQgiK2K+Pt2fDx5LneJuaSap8c0qzf7jyqU7zf5RUnU
ItiZ2C7Efp/JAYsPQn8NFkJox/v13zt48Fg4e0bD74aNyhZ1KvSZY6q1OK5F79Qw
C4zhyw3/K0EwZGBdN7D1qmECGzgfDBMA1LAqsb6iNLXMPoEQsgoJbceqIDQbJOre
GGBZ7BkYOWsp5ioMQ3Fzo3kdxe/sRd8+Gd61M4Fv9sJeV7pMVXPA8yKiuSfS9KjO
KqyIo5qzsQvgp0+L6xTDgv9JE1lD7744a+TLlkoKj1ysFo8n3ZLM9ZYpRiE9gFa5
3hO6yLic0087e2GWv2eTVr3QlLvAIkUsnq31e0SuKY+E5MBX5C9kRrdMCElQKz3h
zoXsxCn+cSwh9joSDGrgarbSE7Op8K81VuGI2r7QagMPGJ8CVRxgfdHZi3qZnppO
wM1ZDUYKNeGIlm4RjjwaZIc6Xq2wcRp6eYzswn5Y1ncxF4dleptisp0ulpF/wMeb
XZvLqiCX9p3aqjQbnGouUqW1u8EkR2qmIkz6ecKqe9YYoOmAuG4y/PnUD0VfPjwq
SX5C64GZ28VHJm+7CRpDBf+ZUjzkAn19h35OVHKc9glKDQn7TO11h5f0h4JJFmFH
SroyNHcm+1aPhsLHkdP30XV3E7f41K6kdbPhaIepoFzr7XCNAfVo9h5XfQ6mrpfE
+1G+ioiM9qFsYU7qbAIyhQB/GrtcwaBUDaC5Ywa9AsZ4SNRlvd1cmAJo0200QPHz
6DHM/POU30zu3XhcHrAoWtC9oc0pfoRiHCsa5Ro+tdFp5xsLZrX4fswn1Vn6P3uq
Llyrt2gWphb8sahnNOmfWnSNWWzFQ1mDO6WvWn7XdOVrJRTilnBsVVpPk8dmZGax
5woOfcisHm9ADNAUAS80xn+xwgKpUYrjQPp+vmDWdgGjnhO4UQ57kIuZVArdZ8tb
CqhxARaZefTNnQ9yZhkckAJlYEypysVty0F3e6gT4Zs7Mr6U1c6RBtUj/wwy/Uig
UJT4MWHhRIR10qKPqsK3PjonKNA9ZgNzpWo7LrnrdS8wuzqeHsTzoPvm6y7zFZ6Y
Ac5c6zsUBumxn88LIVznqb1+I4+5/USTMjsP/vTfN4H6gIz5aVLvGCqxQ62UX+2A
H5aCFpXh3EaGWC2biQXdpRNqUheTfVj6k9kPhGW7sAsfvzrZRFyucaUbZ/h1j8F4
C80wzCuLjjc9eeftXwPkM2QXXRKc9EqtqkVYlQVMpjXoIJwSeZBOY9c2Y0qQ3ceq
I/I9nvkid+R091D6j1DzQ6XUwxqTw8LsxM99A4wUdfun/AA2JeOrZMTwtWlp9MSy
4PVGYm5aNr53xfGbGbZfO4ddj3/CZsMK/6K7Kn7Zlh95YO3wWAudhoEq0pX0uaHc
08ESxOWipzbwzf94MvQ7w//DSQ43E+1ZU4NtFvjGKSiF2XXR5+RixKXOQuRjaDDW
ncCnE+rV9zINJWZ2eITiTp6Zps+3yP7qEqZE+Lwj0RZD2GzfKd3fwGw/CcdCOOBy
iZ4N6qj/lr6zbOqc11NFAR4T10bbcvtS4t+sGHL+ObULL0bjyGp7o2qsPAST1kvo
LSKueFBm6V4gVPGOi/m4SRZk8u07dVs+hPYbGX9OHDKpdpBGlAzCPXY2QU/Co1MH
UD6PWSKiYG0UuxB6sF63l42JRAME6wlE0s2DZ+I6aNjbcKWUp80Onf9ox6DwUa9D
61zC+AIuYPPYRWCcrRqU5NzSqM5vG/mJ7R9d9s1PXll2U/RAgisk4DA+9oBsdpFm
FbxLicxhSH7Yw/JmJEx/S6oIts/Jx8hV3Nv2hYIkb4EzzMD9GQns42rb4L/9pSl9
t/1OphDIDL4f4NzHpvskbxlVsPiCcACjO1ZlkrwJh1s1XAape8B8vW+KHst6Y5Ak
8CA5D7lLAMri0Qgbj3uPNxd5+4UkzH07Of5xPqStRkZC1RnEVnYEQXkQNqTZkNKr
BNJgwhY05gqqKvOje2tub9YmUFd6K42mlrMYjof2bVZ5Bv6yVbvvsb1kfl4XR3H6
VCrCj6wm9vYI7DAprS+t+d8pPg15Rj89+ILyZGw7KFkVUlPMHoq5tDoMzboVg8ri
i6h0CH/i3GzI0Sc0acZKnu4saUxhm6A4d2+V0ZRKXES8EkdpLIEwEc4/4LAOP9pP
kxgg7f3IagBC8SLcix7iu5GHAKtwhL/66RvjEmHEXYGv8bBXtTS/heJ+Rjg1lH8n
FZFxbyrQx70nGjkG1/MSaxV3iwsR0seFVZfFWV9Ms1F9RthQuIAYyoSPR3BLFUNZ
GaCGJnkSyDBrWo4wNYqMiOfn8tlJQ2qUbtFkaDUlIEzmOHytbVAROChb7P2fia23
ya6Tlxu29ER1GbguGb4kXuFQzr4a+rr1VPdrmNdJtocYeY1lfNLz6TXb3GLxgWy9
j13xutgbTMbeHMqZ8LHKjvxaioakEGAU+SwcMEs0vErUC7PKtmDcCjm16PEpPqG8
G+O2LLnoRcDnVEeVJDeWHanKXW/H8HfUTNe/B24VfEtLKBobAiEf4bhXqz6frGGG
qyqPDc1vl/zUi+XOyezNfX5cdnmUTMBJVdVyTA1la418U40DLbsbnzVZebyh6NBT
0e+JlX4mtbIS0DXjRBvbkNrfhg53Uca8U/+z0clY/R9l54fzECf4vJW2g/OyfIy0
suAygSAhmVbOx4obuTUNeh3j1+wbWzrEv5OkaQ9cRVKE9HCNfKQFR8QPhKKHQM8w
V5YMUHPxR1+RK5nDMWYYk1V12sY9YPnIUsMLX4hl0yc7ReUVFA8h6S6pH5Con29r
csNiz0r4q5Y5H5JTcEmbPlU04xdqnl7P1RlBTZMvJgf0ge7h299xMeMwGQ9tz2Ho
N0HY1XmBTSmtr8qcm1OJ/sC4VP2oS+xVR4nCjg0yTIFH4DGcW1hsT2WdAckLI1VJ
nZq+XvVOK7o8M8FRZ2DGDeB+DFkPTVRbddSLdGtcJMwvV9YsoGjv0F2C9k+3fseF
LaHmRszUHI0JSocf/5F5IdCsuPvjjX4Y6q99E2LAbO/W2TJdAX6Tn+Hemer2jhvj
53o9e2HIcbX18OM3zTdC4eFf/jM3A/I6QYhFAvO7raE+o/OJUovqNI+e+gfje1nd
EKdhCgdv//EVLOkm+aI5w5MVASn6ORapMcgp9KYs8a/mAQr3B/GdTg9fB/KnNGOz
fDV2wihW0Iw9uk4SggJyI2VGmiC6zPtW0ggwGCiZeg6h+R9oxxVlx6KCF6wtkatt
pK0WJA7hwke34MVwfdDbarEYSQv7kEwOvGjdg/vpQw9ikxJ39faY7y86M4OzDZKJ
rbJw/9yak7AokJNZdZi0pSErxnJOFbBc71q1A4BPUndfEtxVOZPJ6H2kE5ZYIKgN
7v6R6QQBF6HOJYVEJSWw4gkF+x+/1xJnBufg031PPkGkC2wPNs28a+Aa+4lJUU0K
xn8MsBC1i/O0zgBJwrsuuqbyDeqVL7G4gOqST5qPem/4gNYIShszfL2FrW2qaqH9
NgUvjZJQwnk5H/5pcY0RKfNB2ecWU0Ue8rmbI9oXSOdI8wOsgkShIl7lo3T3iCqK
TO+CHzBISp8dcYVo+IU+LFhA2TmeW65BOkC77g2R6p7JlK5Fog0hoNQDTIdfDJAK
E4vLJ+4go9/HgjESwPlywuBPH6qR9+tluVLYx5vm5nB7cf2YmTRnL9iwD3mFaG62
AmFTB3//eSC4jRE++ay1DLv6OuH6tPev4i/EVkcQFPmhVrUzC2ItaTEfk7AZaF3V
aymdvUqYrWoe7iEGaMYNVyeQKgRZgl5bMZgO3Nr/FuFoN1hfTNZ8l6iqAb+y6UFY
wvtY7cWHjObGmYaoU+uY1XjD97WZBJ+vgfB1m93IBDMO5TuPNrQSb3XD7QhoONf+
8BcZWuz1SzrKSNe8Puy6wMclE7n/ICAy/aPA0s3HemW3KyNto6p1nyuzqKwLjQ0R
+xu8sop1WgHoUn7ezLaf7s0NXb+SUN+30gWDVxr2ZTHkZEE6YZNK8d30cpsSukHW
93n4QxCKSXRzm7cVHxzgNpoy2bZ6UyKlGp6VeTe099chg4WtIUqR0FhWjTeGmTt7
6gT9l/KRv451EZnDMtZlhwuGwIh02WEtnxH0zk/u5G0DkbhapmTvg0Cbp+tcTFvQ
6ZzYN6GeCu61ZT6L963UtTE+HjV5gbucC52+nG5JmKS3mGTovd7/DZer8+VXjotp
y3YWJyKmSL0uE23fQ5tW0HE5IKjoZp+VRCc6QMoM4Gg8RKms8Yq/bFi0FOQR7OMe
CELhOLopcTgG9cHDsA5jl1WZ9jePyiQB1PqnVdYVhUBuh9U2sJQJ5zqI9x7wmWk9
tH0XHUuhTBZULCzq+ty1gk/rEiK4kdg6GIuS/oQm22fe5RPImLvexht2tV3g5xTN
YMsPI6ny2PZ4tDZUwa2R92N6lGakekIh4mkSu8cBERBHKwS//6+se7J0vA/PALUC
v969/8asBSiT+K90uTAGKiWysWQLFecRKHD5/Zluu/ErAYrFHfmFkY+/ovkGddH/
B0aaZEyS+lqhL31p6ckT83h1lzFb0aV8MABHLqKkzNGmhAq/ClWiMvIe15q3Ap7r
2D0lOdJSlIimeySCtXhZk0gRP5RyOsc4BR2w6z+pER/qVvFNNdo/McGSqYmr+Rjk
LHDXlQ6q/YJ2Xr8TY/+t6V/hkd5d9b1wEYWCf3vf3gSEEr4isI4oxLKKj8trzISh
Y8ZFgT6HigHk/eI/Kz+F2LleXAQ83yRPNxRITyxL+/U80T3j/RbjTh7lJ5TFnYzd
q+UKGkvFKfi1P7OZtWfFhwRX4vxeHXs7PPz5WA26FGS3WUHylrL2gPD+yS+ijeSf
IUR94vxlg62YVxQhOFTqWdjdEpVyJyQrjEoXrShhXdG4DTpNxgDPA2ht3OwFggXf
cszS2nkdaOAnvmFvkOEoSnKnQM4ZoNP3z1MB3NL7PQYwqOHnKwhAGsTtq/3zGvnF
yShuCXBApeC71SctDBC5D1DR0nD10VTPsJp9vHdGJc0n3M0BgipsiF66zZo/ohNd
xb8ziz4VpJdm1tcr4kj7Ct9Kyvh2P0RIaKFj+BtFrpr3XEA3dpQSQe2lcw9bkmXn
5SBxBSCu6JSR7NT5YXAYDM87RMMG+rl+Mu5VeQQBWfrmBB1UYDzz9lbz1i5ECaM6
st2wWh5f78M5GBi01c6nBOnscsgMcPcZVDh2eRtgodFrqIKcvngkIPDo6ri3ycpj
AnpO2XOucPK7ob36/P8SXeXOw27tbXnrkTvDBEo4h9CF8hBZtjjQze8oqjuT3aGT
ecHztc7em64LpckEKnkYqBmFaRt7eR4SVMmAwS5FxbJTQ5+mr74YVQOvdIpFO9yH
LjgbXnGFFpPuJv7oNH+rIMZTyzhMQCeAJaB940Ud16TCw2FoaydXBhGkfSF9NPnm
YxfJr21DQeDG7nqelqvBWOyV/hFmM/WTbAmlNaLeQPWtECLEKcQ+wNEFDnbLeAwM
LFkO1vXWnjjib2g2O5T+pUf7kRtN9Hu6LwIFkmSRbWsB4wOxQqzebsP5kC9C1iN3
td//kzXc2qn/Cq27Kguhfi0yXO82jUjkeamzzUhukr5PFZ9Q9zUxjmY6RiMNcIeg
lH2p942BvpTt3ozyOgIhDG2J0Yf2IGYZ8JphzkXDBWYzmXz9P5M9gnoL1hr8Qbm7
FxEmB7L6z9yIAWcBu8NqiHzQ9Aa3Sf1+CFiTWLkZwX1OagB9tsrsMuHIbVcX1cgy
Y1YOj5jieZSvls7murdadVqTsWylGe3ElX8clhH2+p5u5Tq5KuyXd4/FEfxa4NKd
u84theuGNOOytONC/ftfuvBFDttE/Gdr5WaLJCfAATvynEvHejLHXOghvbsZiBNE
o7w+TP5yYVMiF1WvNvbvfFrS/ZZpbgU337e+WyTfPbDfH2ym9BtTJiTTbi8oZnM5
heORVWpDUu5bAU64nA3UNgxzkriFXZZPUE/vEgQo2Opx6YHEEqzDumF1EEo449F0
XYAYN9g2y8v6DdoWvMji3g5ZrqcIC8E3HyDm8iSJq3Nd3l1uM0TnAmfJkJiifMzu
ima32DqMfV/2SyHehFyqrfsOXyrDRFK1tErz0ON+QuHlAMTUo/xQTM+2oyNL5MmI
TCaA4ojkWbISK3KAEIAX0dOhxsyBDNLY2vC6u/qBmgTPcrx60DP6q2jNCaFRQSQM
pvIPMWJyBeRD8Y4k/X48cZpPyXkJUl7kHhZ3EAjgrFreslEwgQrjmfCH2V32YNFi
07CYVVvax9FVzY7ElYq+eDDiSSK6mr2pC1irtuMLZL+JCrOhirYW2nqLgmq+0+/m
FLka2+BgBd8MBMnaZu9bm+aQL3lvh5qk43uexLvboarJiagbqvIWj4q4zJSS+DO/
XOw7+x8d7+gHEPIB6eBSWoygabWsZ2gJzbB74Vj8AQaijtUwP3fVJfudZutEKpqQ
SAOSh4pNvC3N6vSptQs1KG9wP9cR742gwGWg9lQuJzon80IsvR2bUV2RBo55IB7S
XIpjfWmbbCXlBzKbCqtqmBS8j0K4yJmBBKwuC/ShCwUsKqbrvoP6ycwLE9HF22vW
ypeZ+IULIcY7o2w4V3+OXwQQyJ6FIkWfLK+01jDSTSIaMDyq+uvrco1FBN/wdRSq
P/w+7GmrMWPdWVI10pbmgu4cqv2wi07TxcwDawwNNV0Bfwu3tVe3C8D/KEiePZf8
migh/iSXjthJBPVFVtPrYNEWWfl2pvmYM2AtxwyW/7gLQG+h14F1rJ+dYidzy3FR
P7vuGObqkiUAZ9RsmUPBlt3WE6Ai7oY9++IEmMdkK+qQUvIG/6/KkVU29jpydm+j
0Oor5urfsdPaCtUmniP2mCuoGqNTeXCUS1KxWEiFYhfM282PoueeZ26txu3MB5dt
tbG9IdRs3HzWjeXjUG9iNQw34H0YTQVe15NFqzfDx7jJZYwnE1dGClMR4sTKqQNl
pf6pasBM/n90d/O4MDWdHIvAdlxko2sDY623CK7Whg5H8G0WUzWtwgtnw9F8kjUs
qRjW3sE0kpsMwBJALWBjjU9S//OPBXnbDanQmbNBjXcesRCiadWKTXd9yVddFRXI
rcnvCZDvzlorRFGM4pIKcu9wSs77u9zBDAa8IaUP8Id8+NWI5SERc1lJI2gOE8WJ
FNpy2BYlAa7crsc70Y4niFvtau5xT7TNJrHkP8bnCmkeAT5yU31blIyCVfFoaAyE
26uhJb3PZIXmbkBioqBWqwm7RuSvBdAgB/U0S1PcG3vOQuAtC32X9jX8x4JvVAji
xvroMhH7gzFSkAjdWhLCtVzzycoWI4jkTFsD80jvL1k+n0dem17gGqOEg9Uaw6ju
8CuV3TGd1+aXxWsUmAoAGXKwU2t8IgeulYmDb6sPwyvXQOIbOg86m1mhkVyCPKg3
dFUcVMNk6b6fAw8Eq4d++d3dd3roO5W02Qsa2W1sjmlrY6VBRIgEvvtekiYNcNsT
YLyhow3wo6oCAQyd+Ha2LzyqsK52jOWRB3JRkDxgGGjvZ/sb3sF1MrMLdIRyRna3
lDlomuLtJN050rlxRqGmfB5NEklPzz65sDnDzvc8umP4mYQ7h9UWRDoWjKOgPkOp
TQo+TkT1cs71w/XCS6q4BFiA1Ps/5WHuS8A/coHIsqjXpadOy5lKO3Genb9yfIkq
md/KfMphI5B0DZs9BdTpv4FHy+0gt+0HKMi6qjC6br8vmCFKP6XsOESt+q8IprsB
WKmThiam+4AGkJ1hw6RXljnraXKB1yNok+ZCk6cuKT+LOvLR357GX3Rc0E31+bo7
vpkSti9LLCtJIar0ixsK2Mca2HLWEUSQ9GmBejT1UcmvTxWrNdZCUIk8yi94XkXg
ODndhhL1U83BDWc2c1Esh2VBmgoM5Uy9cfx/orDklR8LGNoGI0lBrsrYjm+IcLbR
7gRLqt5DqP3HZJPsgDnKiK31GmFoNuD8Bg/s8NDsf4y9qmW3KadL97RlkpEnKI+X
b8iJlvAEI2ckPFU3mtjoj3lt1folZ77Yr2PfoCxEo5FTQsWT7ynaZNqoCmQxoJf0
wulqVQQKC2pLsIg95uxEyfXXcGfp8rDrkOWhceJG26aT/zr9kdwOKu3NHijpWgKM
d2aTgX5UZWqXqP2+f3ZXfVRYc9KMYoSGUmJIX9Mv2oXFbsqvF3tlddnGJaF+sTyP
wK0Yrqwyj//ZA+Knz0vlKB1+6J9ymnu+9oVGZnAZlIySL//UUnFQExXtN8URi7si
KiTRLi+IgfD2n8p8YS81JeRcfa1kE/PUco0Y4baBWCFCe0RBDIUIgEHLDp65drfB
AuT/M7xxAjCEX5SGS7MqS7JvAL9Sm18E7uR+3yTnlbWocXAc055nPXHkfUcnxhhN
MQ31ERHgf0WqKYTrkiDFKVH9eZvIMwQHunh83ocbfHRTo8tqdwpM5qu+2KF8qJ1o
lox9zepM37mAnJshrf6BmCo+CBnivQWEXo8iyVAqLK1Tl0ONl7LL8Bg9yWEPc7LK
2I6rMOS+GNPmfq1iKlHmWoV1dyx/jUYPFITWEAZZSNZ4SWHLQjo7GNVOjPJdeQFD
lnknd/uXe7KtRBD6pD0gljWN7fvqml47pX2riRQC9agJ9ce61L4Nq5u3r0FAGguF
woRvw4b98yAk8HEP0CwpxPR6Ubi2MkvQeNrGO3mu/plOraN6gnxHUsV5yCSHnrEw
ct5++EPbSHgjsmwMEzBV+2109Y1OEaVFDJnpv7CLYv3kBnuoTV8QIXprDnXBApiC
J3zidjKy3Vuf6XFBZbOZV4gGG1K/U5sLDm5u1QXXXIhS2ByM8wR/ttg8BD75FdOQ
P+44oe3ypFT+8W8ySwEWtwDqa6H4QejvHovudQb51LFLHz43r8tQJGXzekZ9KwxO
S+LH6NPBPhKEydhtCmQGW+uxooSGYxgSHVN3NA9ks4ug7wEcxF/cu+j2Rek92Aro
2PJgbdDAc1Rgv1De9VqdTQ==
`protect end_protected