`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
5UzYaoC3tfpGCmdkAmjlgiHIXpDYKaqWJ86Vovpf/3AXsrmPEcuTFqfwQsYU5pax
pEWcKGwe5JptPSjYsayZ7FKTkTETGPj5hL6FJ5FQ/358g/em/to/rEAxjkIQNRFu
vPlgpMaRX1BInYka8/MZ5YUxYjNqtBm0lTA0ZUVlxSHfenwc6bHvJqSsV0YJ83y+
A6YFqmLVTql4Y3W0HRJWF/svVzq7xeDxfMN/+9QlHrTrWRLI/3Utp+PLS4ey1LgE
CC+DSymtsMu5kI3GqGwlEcNmSk+PdFHoK7ekcdhCYlhvw33ihwDXLMVISH9vcbod
+FnZkvStwIN1L8gVn2Gk4z1zY6TjakcQnN+McabcqlCiFys4QvWJuxlTJ1NtsSyp
u4rMBJcoScH9XupFq7E8eA6yLyR2R98i1UoGLd3oc7O8bA1qUsFGV1dOCpb0NWF9
IabsiUgW7D4r8wWbN8PKXD4TBTroUjrkIWm7x0bR6z1UMcDxdtpFiBgjaCAU2w8j
0qsSXir9Q7n0N8EnDikC3oGjROIEvzkP280NFhPZvTDEqlfdgBcnIo/5M7USPN+g
MECYlfVvy7wwSOeYDZQ/6tYECyoaevByqVz6dJVv65Om0tuxAdskOhiuzyQn+F4g
4P8d331msHkS+eqoXClswu+0TSfRYdNqoUyhPiG3hnE0X2QLz0HOjWHueOSH6qyN
f0PJfOlT18lQZkVVepa6YGsqKUsArR6ss9M5F0eqpwAxlx29Dd2KAmeFS1pxIWuA
KptiAHVRF1w3HIR1PGcc7YgKWZxQbvtG1ngxAUmRwxZoWc9aaC+llqCKaNCYno8w
wATViRHNpzEJOunBhq64YMdIfmjNszwzoXOUAPI/kNz9d9RQPZlPP6yRxaWfFjD/
HeyT8vuAOiTTwkeJ7zZcFIQYSQUMpnlUCyfStYVTYNfx/2lrOGdpFZjs1NciIipb
jUat1UhwqcKv9mWCX20lB3YJ1Sl7UmOEXNt2r5qArZTw2ZOSUFq+FoVQHzDxRSc3
Pwb5cnTSi/jjUjYxqFmtluvbC/4mnsgQ74ZuzlawYde0OzcO7W7DKWWTkA8Hdnhy
SWNhHqxzD16J58NPH8xlUFKMSg1ETtVLZcvxtLT5zEKHhAcivHCV0WPbG9oexGtW
TA+KRYEVNHzZ7LeSV35Jz0AOLq/lY1vENSZwfL9WLBfr43Uyj/59i64dQrdDFqoH
S2DYJ75niDbZEUNgESpmhJ5UkdNp+ATa5VUNT/d9GHTO/9O6gDOJb0LVSNNGmCzf
S5TZEML7rgWJY1jy2tYond5VVYoNwYOChiuu/BRFkyjCWGLZq9QsgyXwlnsdE8MC
GovvTclNkyXw2ABWrVmzIXA3m2BAiTkqy9kEUTfHviAgC861oZz5noQ9T6DrkwqR
GDAjhr9b1jJb7PB6n9bXYEfZcHtXJ2uMLo0vpovzPWymqcbrwMwLwvC2UCB7mgdE
zFssncNGc7eoSDxMPcDKovpicd/VR5EuySPjk6cryPJ+CU4ZYQhnLwihyJCxlCBj
8VzXD05S1xvtra/UU3zvwTfOG4R/5E+jeZuSE3mBf/kOEkNrg2Kf8ngWij+Pm1k0
h0E6logysKcnceWdZY+WPB6i9Ma2tZIZYHZnqi00cZwSyIXgvuvmfaAS9cKv5FPK
T7s3c+Ho3HK0ARJdAoi2jBOHbD/5/VcELF96fyvOiyn0zIe4PwwQstKctb6uQbfb
JMMqnCRYOn7Uk6eTzJYzhdNSyB2ekzK1RZ/2QQrM6bH4Sgstz3AbvvdyjlwWpEJ3
alACWWMsiWuEl9h1r/AtKzF8OnUwn6rXb3KM49Aq75jPBJ3ezRUxU7wkRuqPdk46
QSBv3QWxcp4zUNuA2NAgGCWH2y8R4E+5cc7pu49brbztaob8WmU1+fmC7Fd/4QGw
eN4VXWHlYbXdMtnviLSLEjkj0kuDxth4kZLC53XmWjyj0KC2g0c38YFTzVv0KFC+
yZ6Z8rTlwmtTffM11TdugGByZeW/EgZsvy9f2UJ01Jr2V8DqP3GGvL+figvEyy29
ot7qyHyO5p+m6figTm6LRYrgzp8+IcgWORwDJbqPgEWHjLLI4AFiCGZBbrpfgfdO
GWx85XvUi9uqze8Z0LpIARcCXLHmL2SL+gqpo8D0MESPnfDeBb0rdcBzJfiLCZA8
yACY5hW3Sm/aC+mCLcof0CAS5IEsVCxSRBiru/twveEvTY8hf24zcamXc+EUxb9h
jT8rVInPd/Jl8RBqRrYtmp1uwvH7NLET3QQ6D3AfTFG/hW63hSFigdyjrCuJA2zJ
0tochoap+GphdOo5/NFKsJfO6s5MvJYEyS8MgETXPRUFCcy5HZLaW+hvGidq78kr
gY/+g2dmiXL0SzfiI4BHFtdzKHMoCoCrBt692hyMMhX6oaDAi+IH46K3egJbWz1B
AL0U2JqmwULadPD5FjTFnbNwdCcVtMUqd93/xq6zJxOJ0lEKG450u4UzTsM4G5yn
bqa6SG9+GQsTScrsAiYBsFgJ6s8ReOSXCMlVmcfcDlYqEujlm3Cc+hZMlMVuJNhI
`protect end_protected