`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3952 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhDB3ruPjBpbjY7601ZaNdHSs618xFF3kDHo/c+eTTl/4
vhEAmXo5tmy0l2ak+2z3Y/avO2YDsiz6jSBGXe0865xkfjDwft6EslxCsp8i39qT
mdQzwHoHQTncbszDxdRMGKW3zdnCk0lN/gmkuOwL/4wp9QS/L3vhv3tz+7wQIgl7
HaQOidshJjqrHuBv0TlFMpCP7tQMpt/cFEdyP/L4WJ2PSe4CP9ZyhCNkqE+0Cbgj
Ywiht2XAT8MbOnluJlo2GjTom8JMNlculisLqr0pk0DeaXSg6oxDXR4S+JMMdbsZ
OBPhkIlvt+T34IFRC5cBLihvXIACRySHenuaov6mmZdJwfl+rwCpVzxi2jFwI58r
7icPcwziZezwuCm5neAD5Zr665AHv/QQAJRLtCxJh+jTw2PqoPO8nYJWNcr/7KuQ
PHhU6FyNnQmt/xgD9MxEjpB9P2h3iw0za63MC7teqwqP3E0Dt5YKhzpqN9Hz1mqB
4AnoWMNysaUEIlSIdxKC9W9ge2FdwGItZVTdbp/TMV7IPzGSiKRDAAv6mO5cI90+
Ig1KnSLG2v8mLBLWyBLDjILUlXq/DjhdfBOZo1LSVeBY42oCj1b4Kghc4fMxGwe2
izGd31MOwSHXljL+bUm4QGJv1zJmL3/FLWyvOaldSbKMK2zApxiVqEU/HcmGEn+R
N1CJEfytqi+oPbf7Feaou7n0na6veTe5BWx8ymZyf173Bh91Op/FcF0ln/MbXYZG
9BtW61OXkfo1jcxxCNNq/+9kCG8GM0tmXIH0GP0VWtNHrWUSGOxvQKa6gWjMY/Kp
nZNOd68WAuxvFiOiJ110iOqrT4IkMQkEHRL0VJ7RhFI6YORGGKmBgyJP8S3N7zQL
MMZAIuBj74MDpNmPrbR9Co/nJ4uLuiLIJCVR+ocW2LKK1TiK+nLP6B4axz7Ri1yl
FSD8iR1yB9ZeB6sG8MN2nHpkITpFI0ktG97DLEWOaYaYajStom3KkopYzeAa/uBQ
5GERi0tuRqJCBZQYdgDC0RP8WyXpKYHd5XC4WxqMawH4M1fFjFPXLxh+Yad2yvl/
db9VmvEfsAYo82Mcp4YjqLPz06M0Tfr+hNQgVT4LzsNSl9nF8nXOQsz80/PLE6F+
r2KzDHNv/bcb+pSzHPZHdPDYF/uZqTJrYe/nh/G4MfYQDTfkUidi3vSqpukYXCaI
4FI7DgbX9f+bCn9OmkT2P4jeeg61297iH5SDNEFbvsEW5QTc7wEDmwsvoU4RRXvS
VbHv1yR23y+tENgElynMJLvP8ihq0zP77QiOfhh8YffO1XJxipjUWId46eXEOyAX
paUoV4mhEkCLIMGiLXmWSMFCf8++6mxsmUfade40+/43o2zUV1shPdte9oMY9BAy
bq7dfXyZjzYC1g8e0j/9CuU7jolMsQM7FmDpf8A+hHe8wQ6qE3WIMSxHWLD7Qawx
FsEu1YQh7g46ErMGrv30b4SI2ptOKE2CwW5p4slwpxYxMFLgYfW7qGUbnFjLiwoO
GHGBmm/H7sy8um0J0I7tFwibMW2peSlppQinT3fqWfEurjc8axo6QnL/gDHu2rNf
v5ERPH4cI4Lkpx1QdfppOJhNaBpY5GYAUFrqzbsPpYqjRDt81hRb96CTIy/I+65u
ko6kP7C2Qg/J9Kq7IQ98a/1Rk8bC37IjhEb72pEKSyHQ+hlanzCU5IIP8+PmsUuU
jFMQT9l74zSwDJe49qoNIE+Y5gk9nTrLJF0/o9yrWRTficyFawu87mOJkQmS0VxM
sUxiRPSxxnrEd4wVqvnOHRYyKXCc6eTaZhKhFVL9IF5+YTExsKt5YayfExeQchew
I/jrJUFiVeLSSJPBNljj1Be3d1nMdc4Clj/66SEHHgrWQ/oNjeoGJB/zFRGGmObO
fgGTGvYNFJtWOItD8VcIMG3LlvYEExX92JqZJ9mlTFEMOZRaI+cR+SVYczdkKSFx
c2BH4A+OmsaZWQmaKkjQa7yZ9evr5Wmp4tCD08dP6Fbbr5jWifQxr2l2xonuj7zo
4ajbYYIDLe0pqAE3owxl2G1BMWk/FGvT4K9Xl2MpQbzyz09jUDm+UhRMZAKvpJIV
hJitH0AjYlVMMYRyOqz7pLc1nMApzFWSHvuanN4sR+ARl+T9mFKLJ7SalaMcB+kJ
YQeCLz1tlnOdD2DfVvFOs4VvVoIR8ty6jv7I5+ylXMn/EuTwzHdwrKp6VS0+xrHY
Xz9V3QQ/K8sJ6yGfeyFWD+yZi21IfgBXMeJzI/INRCxgwDtcNkr1qRqgdWagNhx2
7CBAaIkPKBhk37UNueU9q1NQZL8fB0XLCxoe0efohIe009Bg8cj3e4jFI9AGkMNQ
ZSskZB8oD616bjfcN+qpfEffkZEoQdXz6INVpiwhaPPt7rzjUN2tUihqA8RbS55f
4YU2bBsXucT0IbRyMsMmeeiLCUaGSIFFj9mzifayDQr7mYCJvtGmC4UNEtvEg2r+
o4IJxtxOYI2AbGUgPxM899/8fIG3CKfwslDBmBjOT01sTX6s8EAGEGYnsegrWYhQ
bt6pVZvEmV+4ka/ky3R96FJlV885h03G4IKZT/VZSpo1M7g44cMg7ZWYVDPWjMK9
zENmP4xpEWGKNxbCGZQ2OwG1RKNCKHstZP4kLHAlshFGeicCInVfCOpPViOx2JBT
AeeebtJylR+iZZoFDQZnp2J1YTvQlHwQ6KnYoJ38rHKmBx102lVi3Kwg8QECzBk6
+LsHATx1TpLm4H0krspW9RrsqPC+wQMAlD+BeYxFMabDPy1v0lT2vA3LBbukeJXc
9zyra0siz8owQkOojTme6+0UazpRlpMR2k+CVaUDMv6irXbtAdC5ituxmw48np6u
lbHbJEGhPqi+PaKnt738tyclaT1j+/K6JdikXoLhIKilVtAnwQjVB9kKRyX+8nV2
Sw4z4AJ445Ucx6Gr/xh38JXjmYR4ApOk9/7jnaNYjUkOuDUB3ZgqKE4K9/6W7NTc
jkM/jxeebVMI0L3ByTqcOLdt52BGcOgC+GEh715+uoCIMk7jHrkGqfFQpRQflglv
5yJNEdSrHclJ2vK0jDPHjiVjHB/V2mvxar8uwcJ+f+iIq7xL9wkLi6inVvwIZWyl
jxym1Lbnni+UZEE6zBBptcABv301pkV8BkchqrslVDRm9Xg+6WjUaQn/c6Lbql5D
SSmXW7dNxQzNyJY2bcLsTtjlttuKBHm87bI9/2BgZu+gqdIgYdkPjjHbDUdiH9sf
rEdjnHXYDDtFf7it88m9cILPTg6Oh0+qPQK6VA5Cm9TgCg0x2VyPNElHi3OBxt4b
YT7TBeK5IfI67m0Lz6sHmCsfedRadihqfAXVFK7B6Q4FF2F/oBa6TXk+pxHSdx/E
vTcOc+dJb0TLE6A89dQJP4SVf9cH0QnJyfs7Ewi90R09KlM6rvrY2hlSXxmu3yVA
ebIQNbgVXX9Rfagewo4OcHuoD7EpYRrn1HtMQLZDbByZnYImwgjxfscpCuCU3lCZ
x3CFYNf/5iVfbn3bJJ5elzk2kdNEAjujnc+SweZ1oTuB/uXKh1dJfHbMxIzEAzkL
CASOqCEFqEgO9xbSfQRpJJUC4mtpU2yaaHzUqSSeKmZ8P3Sy9NVBGQH3tRd01sRR
Ce0cMBI6+bJk/y3E6inu+zKapYjLCfo87CpP7Q/h+O2yxtp51+Oyw3s4P++W4S+d
EoS9Lybg3kWIQnDSO32qifeeHgU6XG3di7Y0OvBJOT390i4BeWlen52fRnXyfCh1
LSrPPd9ELoIXHG2hJIpzEu1eoKaC9JCdAWrGwkMVZIlWPaKP6rKu/il+Xy/6tgLx
YILNoASXxIKfKrCTkLzzDDso56xW8u+7RpyITofknIsml6u4lQkhWAiGwtRVsN2D
hUFyPzBLaBu4ZZDoKNuUeWi8IOlMXzj3RkVWn1rSdoNXecfljLT5jifX4F42eigJ
7LkvV9G6B25/zO7yNIKFhQI96I1LvyxPb/9NcYkzkAwhLCU/UOp7TWsV/fmcJiAM
YHdd3BiEVsEgrNJ+5hUySYcgn5bwqbrVT6cSh3wUFZBYNR77KZuIQ+2A5fY+Cymy
ugylADHMnWOss3RqfPkTOq2Ix0ZTg/np7rY+Kjs+xeRFgtqFZ6HEqDBvkFSu6aFQ
X4uBM8dnWe9z1LmLnz9ZuT9fW6mimmEdtde474jgfkiK/n4CHzMULg2VFlexx1MF
3Ld/cj/Ytd6GFQXMwBwY6FopUgAFqWub3T0jLBkNduyLkKNOBCXJ4BbNEXS+23gK
2jNtSD4i+LSx9TsBxHe1J7k5bDokQwsVuYSNeIviCcKK4QFnbXgnErYMslcEURlE
ARC0kUfrV8dcF5ewVuW1CowJio8yCZYu7lQoS630scrGDQ/D4RYKn7+EdKtk+e1I
fYZ6VFlZOq7IsDQrH8chPvnjSQ+ubgcILSH+W+rfm6WiJJlwVOgSDh0NCm4fk020
jnzEK9Ggabr8feFu1eDDQOTqMZFe9GSnMcSKBwDgn/8LPcat63JpSxDuInDW2H+t
D+yBt8k1lRLNIjEMfpJKZ2qcgbv3zb0c3MsnO7aQI3Z/Rc3f9OccTxSHgDDzl3rO
xRzpEoOhg4lQwPz2FPJXyBr6ORyeuzea8/vDRe3vKauU4/Ks1T7dwEcRPzxG2IHL
75ROIxMJ/w9W3PCrEGbV0Z4ojxTS+mgAoimmkyjlOB+5e1nB+9TeNyMVEqFJypxW
lNSlEG0H1QV/yo7nl51UBLTmvE9SMtUzWL98D0aJWdqkKIA/ovP5XxsWX4Y9TfDx
b4KSOgNzJh1CCUHS9MH8wsIBFb2irkhKFR+7QOPEtNMyhwcLHvlvF/LeEQwA5yGv
lCQ1dOoZuY5VbKbN/yPWcc5k8rkqtvIvoCsoesQPc/mUrSUBuDNgPc/4AEnJzoKe
kdYy5A2U6PPCmI/Ohf7VjxRvUA15+1Z6V75tYp0D8pCoEPb6DK3XSANNHtSTv3F0
8BAfTayxfeyh3Od+9P4C9OPUX6tU4M0+Cr+aWGcu2uKr2Mi1Xx+UTkGoNIzpoOAz
rY6x0kDzjoORBDjKWkbFrhKFAgwpdry9lnPXRZ6+Kh9Q9wSL4DOP5yxlkN6h9PA+
ZQh408uEp2egTX6JHczjZA==
`protect end_protected