`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
j9eMmSPGcKCWAR9PvkqZ1R001FU8QKTyJzFqNLn+qur6INyYDE1AI8LWcxAzfnTc
IpZG7ua3uuk5/kQKKQx8ZIPLfmv6H3t3eWjki8YIAtY/d5E7Gq8Z5mNxMYRzGGTg
TCMm6oOrOTVYlCXHE0X9AW696Z7UGfWirVibl8hs19hrFdeZKGiGht4r09vHR+Gl
FQQmSObM5aSK5wu5KOrK5ZUKGHyBhjnIQO5NnittDjOwxV/57nHVg0pdG6JUqyvm
tEgmCY36RCMRGWN7sekPtNHjqpZkmYrVX1T9QF3h73+8ZekZYd2xY2hpHHGYYeWA
t3+Fmb/6NUmoP8+Pt2hI6g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="wX+NBVcG/A5ruHK3pkDqG8ZVPdOz9TJPJ5saXZYSeQ4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
j/hqWUoxjK88VtH4QmjIrexFOSwtsLKOZ/LCP4cmrqgzmR/e71apdtoL+o8nlfy6
eZxDZMmrZmJGoazz2oK6kz7xJU85UCwNc4cxAsVxNdCP19vZxph/nCYZQ9lUFkLH
uLBkOeFP15CD3jG5/dp945fHP13J9SzB/L9PWvDC/gY=
`protect rights_digest_method = "sha256"
`protect end_toolblock="sqDZkaglKf+bDjC7VKm3lOELrT2Jlynh4UhPg2J0Q70="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
f9kZDbPp4NLiAOFOgATj9W35i3s4a7wbt9jeHjHVcJxMoXY8rb8laqS5bNUhXGW/
MOc7UNc1VwolqhkS7G27SLamkGClZZtXSbRcN1N+5kZpEaBEj1343vVznnU2Dre/
1cevKNyx4kKswjhZbozAMjEtZb8dp0beGoH/UIKMqDqUl7me7z29yXAgltDhxgKO
IELUH/d0CjTcEoTx2tKl3z+q8dyrWV48mz/tuJ6viR1l4kADyhS00FhRjwYfEKY6
l4o5EY5Hw85ehlruAuZP+02eXLruNC39OV/5t+WNwGBfzhglxaTKVmmaCozVYiPI
F8aGHF7Ff3aAYdUeyg2XiFUOU+OHYpcDTpJkGlTDq9R+Lx+bpN2WIYBxHYUQ+kN8
2To1hVjdvkQypj1/WWNmUeZjFyjz3AQAOV1ac90qBMY46UgcK2kmFgMuEjmeF0Mv
dwwOnD9jUydedbxy25wVDlDF0FVG+OvfmPk9/Gkg7yhf25hbcGxaUdR+lMHJEWbF
2dKqOkWLn8otVYiav+VT24b2owU2qOo9+Hqfp9Hua3X8Z/0GXb+CgU/Z+e5IAxKq
+6YH3VloedAeyttWkzrPEFR/UtoCKyjPtF5tdOpt4YEd+Nncybvp8SONKjFLImL/
S/gy6skvWugJhg2jZ2uZOj6BaBcaEWAbYkZk8Ryhys1SfvpHBfDVXs7t3di1erWW
LYEVB4jqBJLM1HfwslbyWEaDo3Pwvva82tVvmhi/r/TH24a/tKp9Eh1h3d0vBYzp
x7RMNYUfEND13yCh9svYRXtGjmxme0G2Glh0T7mxWcmyjl6zZmUil2wQp1HEhh2N
ZT6z9kydC8kCLt5n70cmX25ox48625+25nOD8bSPjMhARHWpKw4NLvdmzt/UNEtq
rrF0ETKRg5LP57k7loycOFWnDdhE2TaZ9+fhR7uDw6jRKZwI611r95b2WeG0EZLs
Gd/5fRpdDvrYgIsUvvHNlQl/dAGPS42g1fTvegy/Q/6ARLEVIsMsjquCr529i9Th
FxM+LejEtes+oMUeMBqnQl2SoSuFbF8tB0ON3JL/uvnoE2rHQG3t2R3LHkm3wxsS
S5h5VePETPqvN7l2Cj4wvQsXHlEN2cRDdF+x46hc4RAGhwrAo9EghWL27t9jxEI7
lLbb3qkuaUVkTNcqGcLw8109s5eYIS82LYsrT59znkri9gIAjrgI/Avizyu4AmSu
jgwB3TKFNgP0gO8B3wXln0BQTOh4aBlKFBW2JG6AMNgORDHd8h9j0Orf0AJhx45p
bjAQW/eofjl9E34TwZ5uBYW6QO1mZEOTJEYNeLXvjXlUaSPvAF4IlhxkitulQuSg
ztqJzTkq7GvFO7VYqPI2L1whjMAFRTihl5myuykPmoIy/IctNFKHxmC1c0cESTj+
Dirvee+0Zemg6HZmpJTNxTpEgfyt/xmHa0Mzs69WfUVXiuaCygKy6SNWKys1d8Dm
p/ClK45iuavDuOQ99I2slyA8+ZNUWHsBXUAxJzDZLxHNIKF9o2z/9TEvHBe2Qs02
bjaKOCoMdDmSKPvlxXS/q3Q9jYGSTCdlax+a6SPnRilzevj/tVbbdJk1okwadzDH
BTcft+Fw4doy2VgXkSzZp5YZy/GvMiwvoThwuYxw57Ag7Xm1O2oNdPHiTTxMQPVV
yWlIMgwn17/MzDcy8T1kPHNFIF+HUTkq7EslHv1qgsFRWj2Tx+mmokVg+t38pYxc
56lNwXfjcf4f/MfO38cMHWfMPud3jp1xH9yizLH5YzFRNs0OtMqSAohdWztsTbb4
uF7gPVghVNb8yWLbMxWkpzLuE0A+rzoH27MvDrUKqxVJfECgfkNzBM1URbxoq1F4
UGI/LwDSlTFv9bWZosm9APIZwUNgKasVTyoY7Shpm+TTJiFzcqAPDQVFGDSEI+/i
jW5sLoVx4w6XzWlpim4Own0tOaXvdnpcOqb0WpFNeaKGvDRmEf4gk2lh00CDPOco
IhySSA8NLGNEs5B+4o2NBCYQRisLmuHuTAdL7fU02KAcqW1PYtYaaSyiFXWdyCeX
iollxaK0BF7zi4eDqasRZgifX3XTAqKH1iN2z0knmeRescTMNx0hm3gNkLzn10C6
wu+UQvWtYsmYwtJFPkgnU34AJlN2OrbfWM0fHL+jiKaP1Ra6K92xtf1aMr7cE17k
WyibzZUuQueYikPT+yXHqJxFWjLhgzBwqbzjlOqhcrYrNgXiNXzAqlAmTVxccpc5
fT2pP8B4/rkhRNi36LW9F5/DH9amfd3m+dj+F1u4sLxbvap8EmgIiqUegz5ZZogE
fzEgNg45WxI0W2XoDcSRSYKzTxGz6JA8EnOGv01TG1dRWp2BsuUUhLIsPGpN9PHa
abHfKOttECsdnfsCX7Qiy6gmuvA2RXALsSeGHHUpefhmRTZ8bVQVNfkeYj5WNQp9
Vxo791tVKmzr/t56mkGCcPuEaX5CNPXGKlprzrtwhm7km0WKb8jFBwr+jnLJi/IV
2TFZoJ5MVnk2tk36yy4KhWPFDpHkkKDzQGFab8Ed1QKvEE+oF2JYrUdEx8dcSjth
Q2y/AcPRXUcTGj3KkjXYNp463sz7/vTEaY7nsDL/ud8xEusDzuHU4+mlFWM1uxI/
ghlUg1XlamVEZV9snx8EN7xnMUyu9vmTto5IvWn+0qE8MGbH8pxy5aJpUSJmxvzd
JZF2f2a79dy8+9bV0492DEtTgoqguR43OMAVA8Q0rH/Wxsu6MrloUtNk+atIEL18
XWhrPAo/hauFSVdYNb+pGgsBZZsPhig8AtzCdy5GgreyJ5e4Gu8jyt+wcAIhqtUb
lc0BrzL/1cT7QIAVSof5lF43f393Ib1lnkflmWDnh1ry2lk2fo6IXvnlSFv54+vR
1dcY+KQtyD3DbRv1H5bjUdFTmfUwEC+w2ISFWvEffuPKXhl4EcgbOmbt6vA19CBa
8wcT4UM3Ch3QokNQgQrueWm+IvnSXaSyVV94GIn0OmvZIptfQ4o6lV4k4ca+hg5C
04q+3d8Qno3/umvMxEJN96Z3a9RdjOByCpzGesvLMTcjce3HaW/m5oOFfAwKqc9K
XySvKmuNdOJTDCYCGw93vwlIVFQFiC4k5YNCPKLoNJTirGOGzyX5l6yxIDVlDizD
vBU8W+K6UQoz/9GAmWeG4ZjNsyzNAbXWJxkwcEI3whLe5DI17as0BS5L38nFXs38
xh0Dqy+a86Gg1MRe0eoCd36oJND0x2wgBHPzbtVz1rHmeMv2LtEn70E2o703UnAk
vFW8GbRl9GrE1qMGzqW0Kc3qqeCstPS3Cv5LmgL22lWQnev2a3Mlwjya92oljbyy
3dxHCSgHIpBnK/uMCV60ZLcqEf8/VQQLnrDoMj4M4oY0PSkLgwgC+anbJchrTy/E
7KelAEeso3wH8TxMGRhRKas1oUVugP5HsAJLmgCCmzBL0M5ZxAHSh4xTTYp8tQtP
CN67k2W1JA2XJYnpWel/x7esGHkeMpwL2LjLIu73do8EGaFYwAyAuZEsDe57aY3Y
/fz0mjAcSLn6+O4vLBG2JhsNySDazEEvy/DaRrSkys3N92pH4zQl8tWyiqq32yFi
PlUJ39rv86em0oSS6XAk+z6IDdFV4t81bkMWsmq1phNKXKfYN86+uspoCjqz4wEb
nnLbdnliEfSQ7k/ZG3xn93oLrX50kQ0Yb3386/VD1+HEOZE6MpYTT2IRTW/Fb5N7
lT4LqH6ipWlqLqWTTVdtC3m33aOuyti0LZdl/ZQWYrMO2FpJiDJKm9zBq3r5y7Nf
NMRAuyaiC0LzvAtNvE4BFwxHmUdGkpCj0VTpbWB0bkcfCqtjTnrWWRykwUWuDmSo
Q+dvNuyPz++qeJLmV9AJchbIevoOnCalXqwqbIOl3RHRF+yjIQgbRyrFgsyorTns
z+BDthNvGaotjo97SJ7v5JpHR0SIzTGnkJCPv4he0mDK5GcUj0Zn/JdUi3xYwsVb
F6Ygq3SWxarGT3e3PlBUFtS1aEJMnvIBAEScZFm58CMG735dfIfLeoEWHB41eiNp
y7CEBlh+GaAA64kMQ18hwU9olffum+vHYO0mTtNWD/wphxR11tjcizC/1SkO6LmR
2noCGtWH4E4cVgeQVhepeR+Jd40KhTv3ChRyqcfVnAp2+6/wpL6Oy2P5HSQNJrPH
AOF6qxf2DDEhAKlKhRZqNY9MCB0ujpj5iaDKnKRUPoERPGauxR3qXZ6gpKGPSRju
M5lZCWHB3v9+vgbve6cJD8zHE+sf5dl9xYcWMlFxczB7LI4uyYiaHL2MvJbvjDpg
QNowUIBrtPQ54+e/F0GO/em5ved2c6AIR8q4K7qpI4xv2yNW5QLJe2dCFvZHtFRd
IYINSayG5Dhb+VAUyh7fDlpYEcAooAr0iDEdqkvEZr5iYD0B+0tZUPD2tESR4zpP
AFciYUCUhPeL5VUXvk7HtlsOEnBP7vkhn1WLMZA2nyBVgOq98etBJLgLofchqHtc
h6itRCbfv8K67PstgJIJUiMMkCMHLpPTl8y2xGTLoWVPPkuK3pRcDPIln1nBz91F
bn6Vjp7n7ralruA1gflYEQ1VW+9OvORFApDWXRRC4H+uEiq7EthAgsKAgUehjrpD
Rqe6Pf83lo7DMGZQKGrM9Hmr2ZzGLaynZRrlBOSyGxn5oQb79A8VSQdulEaiQpBc
glgc/n258j4Wp4wMWd7oinDTbBEDTpau3gpIpgj7ElU0zmAIFC1z0DKhlm61kykk
jzmYfs9/ZtAu/lz2EljBkfUibeToGhBtpbrD6yVSQUg8Dw6IIi8JDWg0lQymhYN2
A1TpEn6/L2ohmekqWUmsysMk802KHoyyvzMTdYT2bvhcT5h1ZXXxDJNGYTkxbgdG
fsiobfCqOYNYCCKWmgHOEzpecjE9EIHknROTyreCzX7/hXkCz89+WJQwIoLBiTLs
aRTkyvYbLXDV8WQe8vFx0JQNBTUn17BVhK20rdc7+HcnwIEdiWv3YyFcCKTQDQ4Z
j/EeR8QwQqGSHIhNWBfd6xkQsdILCfEFFK5JJrsanCTnf/YPKnWYYmzlGDp4fSj5
rx4zcvplNESO9BKq+oN3c128syuOBiqOunuieR3QWnS6AuMjasj26vqHfasAlty7
+GSeH/ZCX0adDDNcnLOG058vxnLXdeZ2poFh/VogM/vq3W78XsYiTkVSNBP8AEUC
s8GIZUsDR3YC4dDfMOSyhIdt3/vCRWkF/sG7r4TJ65c2gBBo3xgxcsl5ER83xEGG
DHpiNu6fSQ3h2PRWEWyg9Gk70oQm40g6W8sq2mb39LNASe3ZTy7dPHbbhKQdnH92
aGYE3bSSr6yC/gyw0uXgjhQV3C/j+/ouLS3JbplrBIAVoSb8KH2q7cKEwACTj9Cc
ZGLq2l09IT7cCjWdhQPhxEuSsg/jFZWY7EkIBywKBc5HBXtIVbpnyVJI3sSvBifC
ZYGnBImGwieKvG+mzVHJy+vaeub2QGx16oL8sQvcoUGccWIqXrKY7kzd2ssN9VbZ
qMn181uWF8/6odRWmqZ1dDltC01fNfJzFMZj/rcQEHSp1qkCa6ht0AO+zDOh18l7
zPSV8EzBJaXLY9YIgcDnMPgZv7LuTHHwkFCDl9m2V9xdQOL9rzVnSwMB53cChmyW
eoPAiCDR9r8u0bWqUiO0RYX1VZk4fcSEn3ZlxaGaVATDnAUMWYr+Af3QCNZ6DZJN
CDW4xINmho5qJ8vXlnOauMKkwbJd+4IbAXQTPObswUljKdNitBN9V60vP7g9KPFq
FYpvWzN6tnvgcOJ1XKZExYB5TbmqNDF3dsEjW1tDHXSHAgWuUpic96MzObOUmYXz
SJg38/SCK5HdwuoKz2kTqWmwLZurUSSdAR/z17s7vbbhOmvlsmdU6DAiXxyil4cy
eYqjbGQhRkkun6HPvthltEipSvFYxKUQDBDKbkBavn4ZvSIwDSXEWLSYUajI/qIM
xFTEfQxsLUXlJd2B50+aivfPHXcGmY7zglEEuOcaHLvWemsiHWpAdA0HVZ/db8PY
hEAmfFawRIUoht7mVcyx0NdzUgVe/qxiu7GSmdwKGp2fldQfxLcIpglxXvGqqrB9
USoJ2VedPfGKDKXis2hg0NIoOsQ10xq7ut3X59mHIX5YJCsDXWo6N7invjpAiJKT
FTJM2yLq/z6Pv4lrmCfIzgmwowX447NT8MoYTrOALS9dg80wAXFw5mO/0IBznATp
urnTuJvup0qh3P98ndzxsxBtOoq5Ayv9AqvbdRqY8cdlX9rBwtrQdo4r/subi/pq
+HdckOc0JlUn6vbMbbP7MBRGAjQw2UqeVpkBA9TMRwi/fy73+LEKHQyE9I+RlnDn
72ers7hQbYgX4fRO+uVVJH+l9japhgRO7eb0O20ssf0XZ/JQi0o5RHMMSB5Yu6O6
dqZACK/tPtxSmu35xzet1+V/P1kqGhBksPN1D+Bv4qa22k65EtMJiy9NoVNAc25H
+eMXNiKsaEEngARGdvNH+x6E1Tqh9Nz6bNczAlWogbwkWc8jZ7wpE21LNbVRF/cs
PKywTEFzdqYPv0OhPBELtmqvqpZL70TkOb0x2taf52xDO2A6+QjgdjQrWADanF5K
0VlfitZBjCGDa4YOj7lbqNcx0KqIFEJveaYST8N9yhDXZ0gzUKpk2xhblK+YBtUN
Z66PBu+qC5mhaPCCDt5H9mcmqgUrnfrVMXbBSP5rpSEWM79ZPQhrM5hVsSQCIULg
dhpZjJPhWRnfo1vAtIgJSYQZGBS0bUPeYdFN4voGc0lfcFb206CeS4FOjUK9sE6T
yfxDtDM0hF17d8fZRTH0v9afSQtY7VG6eqdWU/JP69ZjPd3cz03hkebFy6QwQEDL
YwitCt/eex5aW+4xGG/+hsKUXdBZ4y+UD6urmpqOzvfvgln+lb7Whba9FYuE9fsI
HXlhaIKL7CihYT99ViiXPU9IqDkYWW5aoTxMB7MZUaVH+xkI4YAAXulwIzLl611S
eO9jR0HTKN0EWTHkQpTRD8g5WvOjcqLKAkI42c2YGP2cfRC0+ExW37GBL709KJ9s
Dn4EKgEICBa5XNpyby6H+/llMWM03xe1JRJAvKPKT1IEo6jb/6Ij16h8ZAtyE2Pm
spqZKqJ9nI9KuMxm7I2+O6yHnIp/vcd6LeSxlecmVZHuBKhtVirBFNCgLx1z0lti
7ztOQ3seSyeOeT1z3ffdZLscpA+jZW2j8P5SIT4fjyCH4aHjKGQnZLgRmuOZZxur
oqFiRTbKGtZ5sfSsK6hYqoUqg56jBndMs7gSZ8xno3bbNPHuc6MMeuzhD1JCR34L
n9ilHskO2nMpLrRIOpM8DxLViI9VJXviXb8CS6I2brMgMnzEcfT5/N4GvNkGT9kf
xwLni8YeaFF1tYpevKRilIoWyKYgCr+0R6Y9jVze2S4rw5y7812nmYtqmhfdSNbu
wwO2/4+VexM0tAaPWbWKz6cNCaWy92GTgmIIJJ2fZvCvt2h8IKfauIWvzPlA5ctt
3EkmV6dwOXJn1PuCpeSwBZ3c4Cx7gvfyXgf2GndzRcFJzdvgC9gkEBQFhmbBlBgt
Bxz+l9hhZRQq66mPODOIgY1QAfvJakHU7v/lRuGPsVE0DSmu/9gw5IgiIJWLsana
rljYqQtPPDO+s0zy3DSgQ6sIc54wsk/T2qEV/FtoVijZnKunbzskutXH77Gog7CT
iigcxEMso7Hw7hDxMiR8MwlXnEKFHrxZ5llcFMPRCO6QQVRxu+jUw8LbloqFD1Zb
rww9aTDzxet1ZlGfbp4sshRWPqOIH+b0vBrYOJn6ln8eYS5tXN3QYXH+G7pyhyIR
mxIxn8HGhdaI6xRGfXjaJfywc7QZjHQzoHMFrN3oWPXJKx6SiPR6nNOUnraxyKBj
Ajduod7IO/wRDYKq4unUjE33HiJ9aZQ7hd4ARMAInSCGnZuqld/4yssK/cJEzjpK
0T8ji1CU7aHm00saPQyKiWOC7hVKe2KSnDw/bfindnp+XlLjpAAzOtqiWJxe7y+m
DX9QZb9Zx889y/kzGPcmB74hLu2U9hK6XeKW77B2R7gPuM3GcCgPqdUxbVNl6n/e
ZzTxzKjZvQxHlITtZyL9EtQDu4aWIqk1h26LlXjUKa/aWV4zm6vHoZGthiOtJGUX
B+j9Ci5QvqD1pYMYwt5+annKzpjkRg4FZ6EHGMLPn//sswN1ekzqDn430P/7YN8I
UZ4iUVgtRVp7VweJPvGON+qL+q+5foFBReYbiBZY5/L+BX75HO90RVEYH3U9W1XL
c1zQWB6wyM1jdY4TPFjoGngEc7dt4/qr2NJ4+8zWFNNfSFWrr9jVKdnb2wiKftf5
HnkV/6AOMC0814fRRfIkqszbOkIC1gZg8pbgmDpOlE7Qm3WTQhYxmOV7KHncZ817
7GzzTIdVTgzevRKJPpcnliC8U4YOdhHpuPsaPLFcaNdBNqbsvi71DC47SN/q6WwE
JIr4tRAaloZLuqm910vmSa7Td3FLNmMJc9xLceQA9X+NOH4IhZfsbcmY0R5a71ND
L64vMvPNWXEBAyjzwJpPW/9P+CJ9czDIVDqpwiWXF0xbamzx5yxqB8ma4VoYJn4e
+smY61jgIAnakvgRKs+TvW6e+KRfWUBUv1LWN5LtnsEvdW1CQAVVaFhFVa0Jcq5e
GcnqMbbAxIS9jyh7rs4DnwCbhOiaJ3I7CqMOYVqT/FzEtpoCbz0i2pXoI/2oJtko
9xE41LjVVmO6zMCVLWULfcB/77uKEDgWs9v+OEcIJFUNZlao7QrTY3QmWTU3+njG
D+UPWyAzVQGfArLZ6Uj6h1umCG68hJHiDYAnF/PjEc2Gs2VamivIJNX4GI/qnD+j
qiR2b/246CcQKM6lqgev5MsGYKBj5TOzBNjifnCA9Kvcf0GvwrV9bLXgWOmaCFQi
vyN/1zssxhkK1diTtN0Zd8c7jZJRY6SfZ8rE2R0w65cDXlM79fGJ1/OUVQIfYmuO
jq/7sS2v6BLCLEWINh48/mpOcsVqrYdSc0RU2x40ODspmolo2qMpVoJH7kIvQ4tS
84P9tO11np6CxG5PbFYhA9/LEUQsszypbK2mrpy51FcLnDqALp6f6n+MZqv7hV6w
YZrQxSH7pyu/gocrmvHkrhNIhU6tJlTqUFSLWtDXjIujEASUJ1lKDd48AP6feVu3
4jomSSo+ygEM8gWAZloM11V5M5dJ+Ud5YWcIUwmpSzt7IoEIxCjfJdQMDjXD2dBk
Qht3PDox9eqyTHpI+tqL94qmYf7/rO0eKjgII2qgilKPdgOTKndbttRZ/eXEp7C6
ukifZKLfMGb1xZaUg35yc9ZP8YA17+wgf3NCPxcQDI3l/b7wqWBT48G8Lq+NvA0T
QjDp6KFVSBJZ/4MXkPzA9huYVF8lTLWyY0NQQH0ePZf8fWMIc/gPdYLhdih32YO4
Fbg10zO/Q6SskEg6fpAfToAyoVm/p2eZDFLJxoZZs+zIk0GrCRHB6yVSc0SeNWwh
EktUdN7o6S8XOjpp6TcYKzpTQwMkVfbg8HlhoMOfYdQ8YOKcUhP9zRvWqe9XQpE4
fdprolWNMAoeWsqUpsqReVk/pbrKLT1E6gWL8Vp7ygg+Nj3mk9beco5CjyfO/QM/
DfqLzGO7PQnlY9AHYWYZsppjFtFLvsmBeaINZlWRXhS5NSApJ9Olig6ahCUyMiEe
pH/ot94CIpQxhoN3MBJHYlEQP1cHtfRn+ihdreQB2AtbyawGrwkIY3MIDpSu2ASS
Rny/+/FuQLAzz4YTerzhR0Y0QU+Jag7qFY/2sTqlWhZFzT1hFfjEaKhvTNnh/ANV
v/teKOsCGzKeVXNggr4d8KeRnC6HTrFb+HbDRQD+dT9FqKZSNNG4+wjy5y3M8MOA
xm8UaqPdjDjnTTW64jJe4OFURy6pIPWcA9n65f4wmOEBJVWl9s76L9sCP7wk1AIb
mkcJmOkknGWiOuCuGul/BfObdZ0XtJxlz2DLAcQ5RhELIsqUJhiUFKfzCmZreF4p
w3akBD82rPvhS8P/Wx7c2xDmhIEbAS/7mciYRJDaGti5BnSz+hneBU/y36BplOtV
YnUE1qFttMxCgCh/Daad0MXhJgZDfxkVmSfZ50+ChF8ri304Ouqx7DdbFdnJA8mh
CDcBhrHnLv2Z/NyNpNOimVxR/xSuLOTAk8tZuDAaONAY0URxI3NWvtnkWqUoprQq
UWqqQY6+JkhPT8T5XoSe7VPgKttxLDn72krEC6Rh/nhs20yM19rdz+EMwB5I92xg
EPM1pk2iplpnze9lUyZ4yWQiJieyCLN/yN6ZC7/ktLKsCwYAjE+Xf1xEmbbexe4L
U1r2PTQn7TX2z4Eca/WId+sDZVIGD52yEIzGNSxm8RPne20OXtPkyfihtFpG7xXY
ZMWOqz8wcNeHdzM0Ycic8o2XF4U1T1eDz7SL3N+weqKHIUEkhAofPBvgUlioL2/x
n4hg2vUg1X5U2qjXMmQPFJe7nWtwsOlmMnDWiuY7iWDDasvZyw1qFPmjjv34ytOr
gKMgjERzCIVSM1hmGt9HpFDkv7Gus4OvDDQPGeSSZh0S9B/treyWKHeDAA1OvIT8
UYGVyLihSEE73X4bI7GBhz5/1KoDbH9OAG74Em4qHlZARiam4Gqh73LQ5Hc+2Az5
qcSE8PyEHhyq3rOxfNSSDQNbY7IxA/ux4K+Q3o5wM97zWeavLXh4bCS3YtteUxdt
EJZAFB8J+G/l/b0VD9spcraOZ7WfMrLlGeUkAHHWCMfRGMoz9bf1yeN0JgNMc9tN
bWmtCXOBqWHa2ZM9DkOwb/QfCa17+IGb0aOXT2YC4mKiMWczAMCa8Mo2VFBk4+Px
VjRPDNsjsk3Y5VbC8AmUcy0kIs4K0Qh2AKs7KQuXrZ7xjr4b7AzoI6EOCsyS1+I6
whYkix4GTSOFUw+JL4LeEwnxFDJRNxOC2nGt9edvfPzNUXyW9iB+QgtKUXorAs8l
jBaAbwHiiEq+d6fWLbNINEj4YjhNA3LR+2mksFqgYwM7cndagkUqo9P5Q89gWoif
g7VcTVfLVZ94ofhVuzB9RNKhABKHcPn518mxTGsDSdsVJ/hY5d8jFsSHeQFLQnoQ
HrHRG4Q/z7z4oZpjSdc909sib3AxL/etlivZTw8egERPmyNIYVcccstV5LMNjBn9
BtIvBmPqtVPj6S2oVaNSCMd00HW4vyTIPh9adkM3ARKEN4TOwYyl7W1kXR3hIgEf
IaTWD1FskH+qczuKGIgqMYt7PM9BlI9AYLnAdnSN1MmlKueecPhWjwNwMFPOJFyw
Me2VdSqvpCBLI10R91nJtGRCirL+JluslTQ3CtzX+gXFMcy5DTyHUagjc+1crPGK
eYst3E/jgKU59I8j40z174TppF1Im20pDggRtGRWEcghEN+K+Db2Ujz/KMIavvZ6
q6KKujIKXa9kEpFmMLRa/7qhmIESNSHFDUsmHxsRNYLU60hzFMc+L7HKHDZNnFZJ
Iwd5mTF6rRbievxSkeBIxLjq+fdT6RSO8RnmCj4epogJxXyGNBvVR1pSj4CaNKUx
HpBmWiV5S6pga9cSx7Q6shxm9Bl+7U1HumCiqsafYH5x6fGjto5jC//mRDxey5CA
aSqMxyI7mkTUFhLOl1VJxSAzJ1C9fkCaAa9c6x8ondimHYDIAXEnX0VhVpnafj8d
Pi15wnznakr4dLHGdEp13ZkFdOkfjUe78rnH3fBBA1+NX/psT5VevfbW2WYtcwL1
8ZEJ+dodpda4Lzx9rmcsWWtL1oAXv++6Qp9N1PMN9v/P90Idvu1isaVACxTHb9gQ
UX5+8XEybUMHLIEuIMx2xRU2+Z6dsk+j6+l8MIuuM2ZHmXxobfnOcbN8zFM8gzWN
6F2ETX3A9jPK1fi4VLhFKkKGC2gr7mFF6zEE1QFl0eL+SsmuuhxhW4NSFO9dJzsY
tstP+WLbqlI3DaaKh7X+69ftSkBBlV0gLWi6CObi84p7/i2r6sYPTTi7z/YPnxIp
wg6+YKL0GY6HndxAABhjAFRwGbogwQJjrBE/YRXu/lWaqZ0gHzsUYqlEgl+Y1e3R
oQUDh7/AJwwm0Nnz/MxMgJkzHoK3ZVqsEhLg+0uCukTGXpWf1M8NvJ12pwNjTyCw
7gJGpea+B0uUmIWlXSXq9X95DN11UjSdSf7PaYpo8CFMBfx6QEPoJdv7Y1Hzhuni
rPo9OCquKcUdoFldly6q2lAVF2LZmKXW08TXh/589MG+rugEQoZKrqgYY7c/3P8Z
TiHxJVZEmVE7q4OQSo6WpWmOl6rdo4NLR0U5O4ep6Q2OlazfNmLDQuhF5Yq/QtXN
uWuNsmBWpUiMJ9hXSLWke2DkU7lXAFTh0xXFuUXU5tPyrxjeykzydCvbn8lx5S5b
jRvsxC69jTWswNiH2zjlOO9Pj8aiF4CA97RzAjgt43wOX3X5Dw6PFi8lFrooenmg
D+pXQzCK15IKHp+s8SVCdEYWS++lb+/RdtC6uZ2WOUUab22GvXXO7hBmP7C2aFSx
srxBoicfWuiwveOLbwMr5ZLCKVDSv/DKaoyr+OqvONgV76L1VAZO3JruBkaDxd0Q
69aAVGu0uqas69UYKo2BuD9S91QTZKu6bXNHJBq404KZzmWW4Mubu75SzZn1Su0+
whaeHBEPqJ7F9ycxUZcD+WvKPZ1hv3ZH5SAcqNFWWt+7mnbyDcDBotckYGKnkz3f
boJUrpU1xgvjWTnvds7Hug99YWJyFYI/XwYDpWK6gOFzXWl3FUyWaHGIsPDWfWRX
fI43RFmjVZYcXEO5qA4vHIZwg2Fp/9+fYiJikXSPaaLUMfcGpmGiyoAd6Rmexgxz
rzyWYUcPqbEt+lfdsyvLOLcQVoQDTf/Qcb8v3aw1unzlFNNNGRWKs8DeqVNK/ITK
l0Q8S8DoZ9ydCXMDRzb+T9Xq3PI9mk1PtjfYnnH4i6RzB0Ss9lx/0R3LQAzgP4Sz
LMt2/J0I3A1/KOQ76C3THp67kB3K31Qje2WR06I+ewPyAT1WN9XKqv2d1n2gwXFk
pFFcjIhjhuRuZJTUHrLbgrGmBiHqR3jxs4t+1iETu8QX6m/VtBkXSyZvP0h2Q7+x
cIW80/27q4+sH/TdJnpKUQT2+LAr5j54XlOskedNvivfxoA0c38RF1GEyuLwHYg2
uspSQJU0BRpUzN1OHv75DMwTfvQykRegCZWuLFDNGS62GTQpWl8Gkc0tIK2fqapZ
P7vBxtLiRA2Nqd1Coz5NIKd9eEHWrQsu2twtDfz9iVZCkn6YqtJ2lahekD9GLqVW
kCjQGnppbugEylaDqeEp0E9cjoZRvVUYC26EPrD4+yiFF1yZjTOSJPOn/RJoZHJE
hWUE9PmjaC0lHfwGdkeAGg3G4oYeoDCTdBGHxwLULdfFq9BNf+P6oX3dkdbnNrGD
jOBB9j2FFQX/R6yP+Q+AudQucSGetVlu0BAFwcZVW/uzV4QH+RGipi+LyXScKkVU
n//ea83k/ac6iM04FzTdNUBhLkkRnvFvErW3REVLA/x+q9sy6QvrgDgft6mqpJic
Msx39OZ49q/VmozbM3KlVng/qAWT5VsLLinG9zTYqjxw4IrEY0DY9qpqovXhF4t8
5tpcdqziovGrH/BBCBggNr7CusuLvMFrIvV5u5tma4StIpbMahde0M6ieWgcDk2Z
5v5R/39WtPICdrBWLLUHU9owScDvR3WIZY0FgluXt1oXqD77wZlhACe6Fk6e9FBm
Vun5nraHF+TKQLfahoyGhYK2nOnhe1y+ue0SHlKSvLTCbcp5wFttsE8wkJGjh31H
kA+DbZhvUGvwIjchpJfbq2xj+/m9KmdjlDVcOsOpwckG1qPSbiUeAMEgiiPfaXGZ
UFEgxMQ7LqKUDEZLg/RKnvguqVJrJKpg5sf7OYsqHm/6rO3KMarW/nInA8FXe+NY
XMARaP2FOIhD518lpBaGqiFEEv5RLJV3wr+bZQeHdbcaIzdzU7G0VqwKvH1AZJcI
suDovhOlxsduhzc+Viv7kTyOPABT0R8V6mvF60LB7++nbxVeFhx9BhqQptoHUVnY
l87fKVCaEnoJbohhkCd0tbRjHfkQQ/39KepOV9f/5zzVhNmJ+NfcRfVgImm2qPfM
X1Mar5W6fg94lgezUWTGV56Pp9wuPxhiR26IuENGRAD81V2v+G+gJp7EpZn67P2C
NXrE75oxz4IiuXD45vDqTr+P3DW1eJljVm7FQfmnlsmXl1HcvN8XYh3GH/a1XnWh
su0mnupfkmTIk084V+Sxuyh6e8lUVMioNGIpVFhUYkSTfe+s+fZalgLBjflXIiJp
YBRD4Y3c0Y5sfaXESA1SiSP8jSNuv8qrjoEKjRkk+/tthlZHdjiCcYOlENRF8/T9
fALQwKTC9ZByKH01rBIuBEYQdH4bUESjtOmbe5wbhZILqYXCucfb/z4OKm2ShYHp
fcUp6X4uWPYt25JlsZXmMBje2Ghqfps7/6TDqH2ZRhKZUS1meffGcEMeDGzYKIL6
eQsLWiQhzvfa7NLABuS73K6G0M9JD/zJA+1547s6JhOTmcFQsrkVhnCVh1FS5MYl
dr9c0Ph+GoQFP9iVdmcZniDyV2ImIkGU49aH+4V/h73/XEy8VzGtNEigQ9wwPX4Z
bQ2dfS0yGWKFu+Cg09k/1aFrzivISCZu25wSpKPcZy/h+ZKPOZkjvBStbzq8hjzZ
G5S2sDLPs15bXgwCTblTOfDqkkk/ddIX6PWXnJ62+AhALJdoXniC1aIu1+M2WiYm
aCOzUPcpuQN9EJLNLa8YkjTnxW1B3lqA4IWpleyxtwXf7q2L09y5uRijYS9lx8dj
YFrj5oNj3/QBvdtTxMJKqN0FvlO/T8ADcQZ4qHiLWEutlwchClOk2LlI6R6mZgF0
29wrVyZil4mwFfWgWxsm8MWOC+Fm1mOVxwWSt8exTzolgoRRTn7Whk9HhEe2AL7f
4jL/9XdfqhI2NaD0fp4CgUrKLba0LhzNsFQHhC9nP0gfVa3BX0yohtdaVA+ai2tN
FU4v+qxVgng7NhUthREmbzIE8gJS75ZtRqIgL8IcmHD1q28zQ6vBQns4lqxsTDgW
Hz/H1Oh6arRk8BibkckpQwyjJFCnJXuguJDr8jqWpuipeECHS4NanROUpmaLsXAg
cospvZrHEX6iy8r9ybp4ZUkzAT4zCcqRFFEB/AFzJAntSwS1BsrJku5KTorm/bk5
i/1bMD2LZgkJ45mE2DKYI0vQX35E3zhAC8/Ioz7GKkJudgv4g6T/6fYjsFImWyxt
eqhrwFCRAOPfg3oPprPxq1DL6/wTpw/w3yt86DVSvjxsQASAJ4JP6jPHO3eXsaTQ
P4X1kU+qtFsPuF7+Z19KbbnG14EZX+u4eLSchn6kJCE/graB17YqrPlnH5ApbLIq
Y0gfHZ+5cKheFC64chSuB7x9icpWltDbtPYXfTpWnVrwnZG7vPu3Tx0mcReiF6dt
+b98oEiBCwMQoo+kUsPdsuKa48rjC4C/WZB0ka2gnIob5pbA0teY6a6dtpj6Mb2j
+8i7GpWZBYwC2idmnTgycRFXmG0tQiD4QjDryX3lCPLjicCzKJJ5FmJWSocJ4G98
cZaBHYq6JJe2XmXvRH7e65vJYWtni/VNnO4oDbwULELNOy37fpj4akYE6iYuu2Fa
wYb8WS5BVD52y66y/EZt40dM6TjXG42p/eglRTYrfcABzJ0K+KaLkCD+LoJh1Tgu
5gXVUa6aHlaAGf332pkMKmzBzbx4IBKerAXKYidOMIzzfZw8g7i8CY5soZFkLl19
BblmRTUor368G+RYRhVGUdOtDKq+nJyqgCRrxwTZV8r7oZ7iZ4EUP9TYZxw/aw4I
EspPwTqi6SpoKYMcwElOtnlKnjpV/HIH+UrLEXGyKtKaOVL86dZeFhsNxL0XgqiJ
Ujj+a1PVEwveLSknFzIzIo6ix1CHX2iD5+IP0eFAN06DW78EYRevzv10+TTwqk16
qeRlAzVg7abclY79eOwhHX6VEqGYxs44Ylm5zFtc6U8gIe2za+yyRzM9BsJGGVxX
GhPTpbZ4PvKMiMDQp24R62/tkI3brt5meC+DjpFobE1xhn1r0BFCCignoM1xlqBC
LeR7x/B3qSIcj+pqT6RKHRxXyWanmlkbZy5j7jmNtHV9CTDl7KIXM/vwH3w54Hrw
vfFiqKtyvVpyFuBJ5KFtj7sxsNdL7U1vhB7timdtmFB/2P4tUv3McoK/+PvhK1oG
N0pKr2Dn7nLSu2kTGLwNUTYfBZRhzn0L1KEszdfzPdLpVpkofFF/Y1ld01kr+8yi
83ey8ZDBwL1cKzV150A3mjvvk6l/daP4zJkmLEtnD0kt29PTyjtu3yWbpcTBtlBb
cNCfP2lA4agU33IY91eEvAf/To8kIn8JBlo3FC/w7IsKypbbbNpvMbqkRJW/TW1v
kUmYqv8g7GgD0NyxSXmtJ4vEEul9pcPhnaoD1GpPxbzogaSqRKFOleAy+Ri71Nw0
mrGn00Yfgj54ZRlSYCq5+czf3GC/ZxpBTWU4jmzjgdmIznBBHyi/uGcuwuphLgCR
RD50/j6SaKIbNvcJlg7Tk73mG0B1+0l3Nj91cSD4qBMuzMQxGwwSzcXue61rj9qT
uhnSpxrjUUlrEdF2bUbHdWkPAtH3JZtlhLutMat1zeoP4JpMxBN0xDkWITOMNIKq
Ztl3Tux6kvvtch6KDxt9eopN3q0hVy/4kkzW+0xJGItvDReaQouDIzY+63M0hyhs
iYubefzYRKznC8+jhsDk5RhO6ufW1jpUyVpPf9DvoHN23+eeKOQlttK4obMSxeLM
ecxeDZiU4ZcNciwPKXYeGRHwi0RqUiUlW9a8Y3Y8yEJt4xaEObt8lTk3ZxH/BaEz
ZGET8Dh5JbMqxBfRI0yNdlBZcTHpjA7WEEOC8vJhHrmkdwxsIzZih/CHXnva9kwK
75L/MPVy0rSHo+FixRlKjWIXhDKbTCBz41Z7DuJZmmjpjEp+kQTsqPuRFgc4cwRU
HU6HIJJUytnUZjqsGG4OYtbtOFeFu5h+iDr64CI+p5sgn5KPKglM6qjxzF4QqvAm
aMkw3VJhJr5dN8jS4GFA+L+eQoJVb77rR58yqmA0oHJCYZG6txsvhgjogaWCgyrL
Cc/JGVZoQk8F+yQcwpCRf5oKJ7tuXe01PForVE+3fPBYgeLW0N8dsWmxsULlYvvH
iMgQ8k2vspgYxGONfR1iYVC1gK+I+Ygs5r4Wk6owwl1/tBTZpCx38/25aORYndFn
aoBbZbW6Wgx3oO/fFNyCQXxGCvvRmHv4+GRubPLGYQPMRxAl2jtNx11aRA3dm0XA
Tp+3lNqLDpim9tFV+sud6Z8UyKqfs9kLlGknLsJPKS65cV5wg68HGTovo6DJW9bP
oSbpo19MqfQlvL27EZVyvJoEgY4WbEvUHCNcQ4pMDUSkldyMx9bIscEYQeLKNOB4
hX1AN7tqfx1N0cLzCl0DXFf70AKDW95gsalvAu6TByo2HdxWmQGjcfY775BXPzKg
OvGdd3iFGv+1zzz9HHAXfBjtlMMf6GVyc1U6d3Ax0y8DUAjijoKqr5AcpsbBdtLh
1VtRFY/5wSpYvu7cn2bH/HeNuxkuz5YZ9zTes4/dZGeI2hIhgdtThOVrbbCaD5iM
DCDHiOx+KrBT8PV5Gz1+FR2hIBngBsLfjz+yqroTuCNIHxgrTm1vX/UpsHw7hyjk
HQqzZyJ+5gM4DVsI9OQin1zf+blxXUZEppMdHwBHQAxIhLukVjEhefQJ1YdqOYJF
Dly8smWafs2G0hCg5RzTXnn12fvU1ejboFrflTiKfxbI3WIH3VFbJsSEQNIG6+at
TTzgh1hy496oeiF9RiBeikiZv1lesiE7cenO1bagjtSM0wufwDXUCFqy76vKg92k
UrP3WvfzoYhFUJXITI/vMpI6CpuYMMBatGVa7HKI1Lj2Xa84o7/Z2QfhgQyjKX4s
Ol7WyVz17iSVxDr+dJKzioFEEPLqpRDHGJI4sYJdYDuGSNchzHYDSQKIpgMfH+c6
ljIKNERdlFoZ3CG+/6vFUiEBAqxFtBJbIiUETHG72EM61gjHB3i05012k0gyqT04
L4lMxTjzoIgV2ISXxY1CLhNxJtpbTSnv+2VnDhLk8voJWv2vaNUP2CSbkzBJa8sw
rhMeIXe3IMm/ushTmifKyo8WACTt06NcTVEWXScGvZ1vm0Dtka+lOjFZj8LGOANM
D7UPmOLD6EZduikYEveEA74Z9TzjuRnEck76CEjwPGeM2HJ49RKq2Yxd0T+G0Byq
AnbcPh8bV4GwtK8ihII/iw0EQrr6F4UpwIP8tyMpOxeHi06GA2591Jw7mFpc0ow8
vaSH/pKtKFhovmPnCdPyDp/KWltugDRo2HtdPS7kZOvvBgSiJRy2VIKjUcjMvH5X
k2Na4q7vutc2/C5BYt4MLQVNVsuenUTTKRPjThb41RHKPlPhG11vjCCq/hKfm1F5
d1IzSAWVQTOygbOGYSDtH2lTY4mgTdxPQzBKUTn5C2GVJswLwrbkVlFPLQW9oOhO
5+yl5dVEUmGAwLp1xKcnVTXGsxfVo8U6vkXdIvGYt+Q2V5yaqhaRLUijIyVgIeqQ
/gKWZwdYnCnaFKS+XgiupUmcFwofjfjaKMTKqmyNRyN6z0zcOvV34MuyON6k7iIU
iclEIzpLhdiEubqlbhQ/GPizMsc/GyVACa/gWn+9v4etCyyGGjbpz2oQgPyd8vLg
wyv5kmvMxs/wHkvWlrGZXyH1gqBm4Nb3klAVdDowZiwMq9qSwasfO87P1FpjxaAn
2ueKZPQfc81o67dDvNIV7bVTPEMCjZs+9momvdQMNZkUgoLNhd5r84vCAIqqVK/v
pAcClQtaN+6qabXpXZ0+FBS2Q1BOM6nz38eebDl+DkIqYgO0QYrFmowxK6DKuLk4
FzYq0DjWTTxR83m09O7gtU/qsen2OHidh9nnGSlwCKCgW2YbezHoKAvMPvZ1fdXG
l7XL0zRkjb5n8XA4bjC6sB0qaK5gGvNKsMgPyLfrgL0S+e+dcLNDK1CnXi7CwJ5c
f/SPvijoFSyRKVpKZ+V7iO1EgoChMDvPxlwsN5STEc8YqxvzqaK8u97qwQ1uT/a+
gHa+n8mAByd+URjlrNhPTD4J15G0wGNqXJuLMk23FnXqyTTFuSmczo3EkRJm4cTt
6ZnS87N9dqhzC8a8942cRzHcp3c8GCa0GacvPvMsqobLu6iGHdix7XTmjql5TGQr
E2FOieuUBi1wVvDugbFakFJIT9S6tSCWiM94E70bgN/uhpQyc2vKtA6WHiM3Uv0T
GZrE5IMI5rt5XBKKleuuRSleTveOC12QtoDHTJqotauWjDBkXCBS1ree1yZi/MlL
AnrPJqRsE+5BDFU2VCVlWKjOWGhgP0hlzg7BMy7UzzU6kvRIdv84u9BJDhM6D3Rw
DNGMHfEHdKDMyc0v6Y1op2eVwQl8tAuSKM/j+dZWIUGjpNIeStoB1qLIhqBXSB5Z
y1PshjtbYBfw5J8AYOfQ2Mt81ZL2AVqrEGR1R0QHllJXasvwqtzO3fAmfVoKul8H
yk64Ah24KFokzKrqdjcn4DFyL6vzWrEi4Xaho6Z+4hrScC/xZAIbMOmcnVFRkKj4
ry7d1zt5qkxTYQirWn1YAMWKkAzXk2aArqzSysM0mOkO+SiDyTiMEJIjc0/AW8Ap
c7x1B7mLjozlNPifn240ankph/V31jVhmvfWF9yve/LGnTKQiZ/CIG/NHJLhZn0I
GGjXjeKSrTZnlW+ypE0vBql66m2wvjHlEwMBqkyRznSuZJgB1UV7PLCg/xjkuTYX
7ARXMHEgNBwMCpgpu6tDtKZqWe1YxTLdltlNqD/keZ+fRYMU0YeZg5y48fIvhg9o
FbkHml32jpWu4T/4kbrBIUk/gaZ98LGB6FQUnNzm9tgJ2zjAM94PmCAnqPuo7yJ+
a4ximCmm2iQp+EjyHfVda8p4dqzhwAjHkXId5A5lYD7EtvTYnRam9IZj53dq94fz
FY6J+/9iCJaRCSEkIfGQy/OIe9ECtLYBqcn+vtijKtmJh83kqZ87q33VCP6Pj0b4
L9i51HzqVJTDJE+wyrS8blsrT9/e+9+n7vUOEwhEh8FPeSCfZ2F2SIl1QsG/Svd7
qUMEE7BSgKVJrLvYRyahctX94is0olGHa5JcbRtt4hX4yjUDvyMP4DuUQXQtlkJA
o+y2juwodz5BkAZwYka3aGM5flESyKpXJI3F3Y48nG7/0iimHUqEykzJ0aNyXkL3
Trkg0I8YEwMNABBx2el0D11BEWj0b0WVaYfISyOvtUFtVjzudo69JvR5OS6gZ8Qw
PD6SwSUTGnDHq1oYFbROvqu2iL7staqTLjxJn1MqzvnmRXIuYqGx9KI+7IQTftLI
6ZlxSyCzxc4RkBkJK3AWzIatrM6Npfx9R5wrq4aQ94kZLHff62LA4BOPGB/WEpJw
2klEcV3H/DtmcqcDUbV82QrW5yNb0X/1MR2pqWxpxwz3MbP5BydUq9XiA6GtaKtP
UrgbBrafK65CMqU4zdcIUD5OM4JIZsdMJM9RctECeq7z0p+Db13RVnLvykeSe0xH
np7RhNXW29VabHCLAIcptaDq33IuY6uN3SF2fTdzhaLL8g1ZzWdtTUt252xRYa5z
6AKn4fs5mRjXvubE46ijKjqTR8sLW5v9jf8hpFozA3pbCzEb2WDw2g9SZGhmreIR
1K/JC15hYJlOOAbaB7LJmXJ0tDJ4vpzBTRS5DqxfAJeQ08ha8iX7AWeMJGJkcrnm
rTNEa0yptxv7K7ohtY0XHK2XIOAZnqzog4Wt+d5nHYDOm2E/mczucBF58ok2lUwq
8FPtTTpDN1HUUFMgHnkA/uapB5nmbYSIxzMZMaY4vglUGO7u7hPozXYJ/uqTo33g
2gqe/Qzo6CnT6lfIKth0PpRTTQIe1RSP7hDH2gThNswoEk6yJ4LYWuYwuHsV8LnO
dKU6WBXLa/lNFfo5pEqNajrWv1ZLFKXE/BoMZV1XuFq4TaPOiVnzoZqJEncNPWDp
mfgEb27/yQ5+9D74/oW7zZjQ5MaxoSHY2bF7fdC+zZ3wctGdX6sfaS9PPHE5sNGr
3hO5Pz3NGeZtjiq7p6VN88S7eWDeM1qXvXpUI2MXMXvrlKXa9k7JS+1rzBtAxWRZ
vADSbNKqolIQKJUIta9sKVc5zTe6zDBzXFNELAIL9kVpQEvQUcDKhVKah0NpAqm5
zC4wfHrwQfh5ABE33SuQnapFKofVp/09vwGMy5+5cljNXye/Cz7PndrcvbmXnh4f
or5DCUFf8imJ9sGOgmPOE77QBfdEK3qMWnRWX6kDXmuGOvprVEI2Wbwv1olmjtds
vh31s0Afo+ClOgeOtms4r45zTaF55SnvQZ7isZUMN27EAuNcOsy3OLFNlU98jk3t
vA7apZvoexacZ9eQvOaCKG/0VlJI5rMv74hlu14pkh+aV/ldN0Ay1YmUggY1pHCI
W1kxsskk0H1AQvYe5WX46Fq4eQtnE7OjvzI0lb5QT3ULeu/s61u04TdD6/cnDLRe
IiZrGsKBlaDgXG1IrR6yW7zm1LQ9nhqb7bhO1w2Ja32CHHBASXJCiOqlNMJA7xu6
DyivfxJg1Be7zg/+bqvEiusHfjR7vCAf2y/H/ul0fMc6+l5fFyOJICo5RkXMQc/e
cLis7c+PsQnMJDmZDXHA8KddTEkQfMFvF79Yc+AsKWMDi03MfXX0jrBAMhTSebFk
kpYN3QAKvjdxHgJ84l4BP3F6MwsSP9GmlgzPgZFV4v/r/qL68Q2asjDijMjHlidV
iJIQEHMDIyL4Ojh2sMxV14DNZoyUn9QFSgMC2M50Ke2eYEvbQiEzkEpHYAq0SfKs
4w2AA9o89byW5m+Pt0G1T3EnbWLYgNTDgurLhnv+S9nwijk1pI3/R4qgAhocsr1+
WhI0pQX8H0ydvYFPDy5peUv5wflEkNa5LvTKo0eyuF2ZCRznpyTsMScv++vcg2tt
P13KThtt4V9Dqh3exSpaPYLf7HE2uq4LWCqigJsNfhvzaqhsa36nUu9mD6bttsmZ
/Kkchd9EqG2XTrizwIXFR/pMueg+6hkvbuwlWKvV1gGo5wTywUAqvBxs+vGX3r8I
QfaDqRW8GRZSIbi6xhFRM1qmWoupwdfu9cP6DoTqeOlAystxxlnh/WNIJIZNArXU
J1s8vgQWvPMEAnUJ2Dpr37aBC2U0NUqisI3XQeJrtAOpjOlV8KP9fL/oDIrHX+Fo
YbNrSbAFWx9rL2RIdbowUWRLmQjZSjVbEfMaNuaISN16KMYhGM8z6J+58ZqGspnN
fiIz1rvXYG7PMf0Hbg8DPRcE5jgG8mT/vgWWD+oTP76cUiqgsT25GJEOGySmmS0n
/U9GSeS4iJVGjS2zp0QbiI6s1gqx0ZNZ+8zCijAnq6B3RsBftert1SdDMQaNuJqR
JIy5VNSKTASoIsQjEJhr9Ii+Jy52hGxHySPcK1v21WpyTsLHtESt6TUBgyeAbtYZ
9+RTyrRB0AisXgqknaUYYcYKYv7RE47Zp4Ial9rrHxw0T4L9p9cmtquV0CKIe1bu
JPspdYP4Wvn/fWPmgNQFHsNEbMBJ8LFaY5IYJmA6XE4E8k12TPSGsKB1zKzdwDsD
zJ/pjgH3b6jOjU6PajSS1R2ccOZsM/6910crEZZP7WgDJ339W3bFt0V03QTGLsUL
5CJuJp3ZTNAtRgyfKrWQKPyLQ6SSZ5/aRXCvSRjfn7+dolONntSUYKIHO+rivItW
dbrHTyZxAlpZbFMnWtqAGM5iBbFmG8ORIS+93IjCLRwJCy0b6lVeE0nyySq/svbd
fiDygxc4QyLi7e3l/sNjao18nTmrnp0lBtNTHtuQwS6xIJufmnVM0bYr2VaIEfSh
ypW6z8Sy953mVTL10SZjdD+LT56OtkrntMjMc+4epOfbh7GWdbf5fKCSRqotUZJ4
oiz4Jy0H8QgHIX9rUGQH0aYFLXGVs3wytG50awM6Kgd1+QRQBaGPl4NCgEkzyBtg
cZnaAtDcpi6TYlgOC2HkKGobH461BTpvKLb1PIBINS5yTekRmrhgvWmHYhitJnkS
3HZxf+hBo84EvcJQIahz9oBEmfMx/7JU9FwtGYG0PyMfdVM/0OtgotoKRIHnq/hI
wSlPFqjsD3pYfAPRtUqth3JRAm9Xbrm+otBsMHc8sA8W/ts+U5P72sM4vKAWU+4o
ampkTA1m2UHCb4hxDuSR+lIOCDkxyha4qty0OOmiFBapIns6O03qS7c6w31ljFa2
pbwT5Q8arg5G3MHYpgkO+ZmB/u8UQD2g03Fjal+XxFyQ3d9FYTWA+EmNGFi4k0t9
ttIXQC9eWlkeNlTvtMJ87N0gitMfSvRoYyostaM5v4VA6DzQZCQ+Rrm0al1G7m2q
+PnsYbqN6ZQAshxkkT81MZs3/+BG4quJSkjNMySLOMe6nIMT9X5U0S9hPWA5C0TU
JSBJdG85TEKCuZIs9BN8DBgX/eiidN46BME3Y/FrXyVuc3OttJRAL+LVe7LXdqji
md0cVb0tfZ+bNtVuLVY+awBE13JjL4pGouJdDIDu4bgtxfmu/pZ4g5F8/MoMfF1O
Yrw0VEOmAFQMmitzvvgE+CdR76KZt95AinJ1TGbXne7hC4TcHOB3X/vF18z6GVM+
LY0JVpMq37692w+krCYWc3uMDybZuGSS6fdQHC8YmI7V4CKQzB0izOgyA3tBP8wu
dFStkA2+gwNaoEBa2CAUKA0Ilt4ffZJZ+fJQbBlReCZQeugc3yb3FN1p94cG6QA6
LEq6tRv9ik7gFfpfjEL30G7JH7hif0HlyqJaY7ldHBnraKKd1UKkrO5/I7YJ6UR0
ZcWkUeYysm5mxyDHaEfN5fbSryKQXhvYUvYDDsnb3fTbydGub9joFHFaJHVxAomH
7K8DQxf/t1pAqcst+h4BCIL/9NRJq7I6vMvJDFkCzM+QlBkAMqcCimS+oPh9puYm
OpR4faoCLIQR59DW8C+IGzyYSsyHaH7Ib0nzyVOmCZFGjpd2FC9oWP0hzLF/6baX
OTIMIpWYC7h/ebGUfbjnsl+MqiHom+ZHMp5IHiJuy7mgdMQaiBTu+IPaSqUGvt2Y
0XogMCVEq3nf4qeHJf7GW2Lxoc6T+uIkNdg93ezcqbYLmNaUM0BG2erUE7o/s5BB
/vhF0vopq9b40osrpwZHc7rdIrOfOyIB+KLOB8AXY22/7ZswEBlTb+07zvU2sD0J
uamhDmw/4DwwCqpQRogMEeI2Q0+gdwdy97zEpfz8u/f7jWsB6PwUJ9GpepeM+mua
x40jOurb//SOPjUcH9L9ajtP8m9+3Z+Ftqv803I1zMewaaLXK53JBX/R+M17OFie
G4dwdorPnlyw+sYnEnLMLFhK8mESkNC3zdNl3iW+Y1zxZNmV7Z++eAm7lh8n8P3l
MYMRcENDIw2K7DhP4QcgjdQ50UvxzdD4ZVsgweT8AFoA/GZPNsD836VTNbEsFHK9
r8pQDRJGktm3nXxi7UHAdOWTuy+QU6yYS9nw3tZxripXjN6/6OBnGLLgRUuSC+s2
lKksowAItD03Ii5PMKmlRLMyaLD6OArZcOHvhUMuXuNk4qH8BYRyh3IWNvM3vj3h
J3l+NDpBe2naEKbh6BODtktey8xn88bjMxehU5b2aYPLwo7myk9+Kkw+2CM0Fjxp
gV7mHOtLbVMbO5zQsnodt9P6VwxSp3zAzB+7RlTCwKGcNJp0gabQVgfQ048ykAH+
Swq7xNQ30tz5EW6lHX1091q2+/7KZ3LIZaASX4trEMUp1zsl/dqmHa8QDeqefskS
FQUwqPfsYdEIMu/EyytyI9vzYUawsiwyhhRq12y77pLTZO6ODjl+mMWwPeX6gkDm
wP2sFpn7rWdHu2KOfcqNo94NcApG6X38wNdCywgJ5P+CC/Y7I9cfcG+oAPQ0qU6h
yZMHXh+kS5slgpDz2j7DVaN0y86vduU0Ja4rTlwLgTSP58TDDDGtzVCtKw+RAD/T
i6AngOpGlLuVO6nKupAzdBc8puGqUOcW4RK22MY3tLUJ7C44gOWJLI657+lYM3Bv
EGzCeqRyXlHIkKzOMneIZDhPuN2yBl1HJh/C1qiw2Ff06yxsxvAncdtOpSvyn8t+
8f04ZyNcNvhfAnH+dZhekd/I/C/X8mSOhkA7GQEyWUqyaLgoCIbuPUMjDcNXFhEg
3mH4EFHBqTQJd5wjXCky0nZ01bK7BS6/rbkQ1pT9W2QpHic59gYwwTcES69wq9oG
zcMpDnAMotZ2Smw/1tMXdzV8TWcwKxaZB3TyTcdUPU847z9uosTR1h3rJ8N8Esuz
mwVktUNgij/3rcrj2iJUag08TqYpBaNkbXxZwt/eT3vC6uz3RSNIyGyrIfPEpsFL
rjYzVz7vSXtGRPTGY5GVgG74IBuLCKy3jmh85CO7y0BNUFfQyTNAtK0AO1rr/Zob
eyUzdQAplDpJJAdhBwrjI1Pr+sAia6ZfN+UZxJXtqImrHnuS1SXjLPaq5gGHXb7C
0gF0OKq1yvYO7OfYXo+f6c+FBIQSRovEEx4FlGWJ69DozCmUCUn4y+GEUC7xmfId
T1xa3GfsKYGYywnB9NFfy8mr1Z0nmjYmUBSwenWLY5m6O2tITg7lYRTZt+pwWMS6
nP487DsYMZBHtfLfCIxYQqZiTGlJVb+lj3Fh3Orx2AMHND8yi5RN47dDiL4SaAvF
S7kYek9UqzH+iEtS5XaR1pjDhFycIe8pPanOkJ3vTfYes/dzOuMdL6qv7q5SK8rN
bE5OEnvzObHCeVxF3K7e2meLn9dr1RtFcGYQGkY9pJRk1ver4kKDziW+hjgzgaFE
voSlelvUTS+7WBp/jRXpplVrgIyVvoY/7syzs7knxldNesFXte3kp30/1F9ds46D
Hix9FdhEK7KJqhr1jcB53LFHzyIGnaKa7nV7Vx37OA78C4hM6KBA8WD6MYJ+5jW9
GsCv1KcEi6mliNxPvFt9W0JFQcD59mylg7DJIdRVZGAfE8agP5d+ScBLUhgSYPZG
qKivr33ioDnmRRZOoCnklZNfbn0FEZefBp0KFC7k/ho3QDwXQPogsJ8z58D3Tlyg
TxcSqPAO1Y8VGLjZBV7iqBO1LJhuXUqcPyfZBSip2edqgD14CmfVF9hRRxmHMV45
vwnhg86iGKQZRBV1lNIYhEg67U8drD65wijWwJvQUySGVmPxU5lp+JTi0pzRAMNZ
P2Pm1jejnVWJWMXOaXe+dAhRgfxDDRZANvFIzuJV9scOl+wq9MhRu/OxVqWlYxmR
/T7AXqxMF7Hlytf6Mdx/9YFDOrzSSPHNc+6TC9Xho5GsN+mQl8DbbdzAbyQtcBKQ
iPo/tMEfAq8LUkjjL8I5uyQCcwiPWz70MN1MjP5J4sqlSFJ6SJ0siNpG6RLo4D3E
xTrbvSYqcAV/3pYnoMJulnDEdizc4FlUSeB8pO2YKcFC0nro6jA1WBsHfg/9wTBF
nJlua8zuiNm/1CdTSaReon0GASFSAfTmf5yDyajroupi/3M3OHQbKcJnl9fhf6hN
tdPc3whLTlPNfEHN/gt3zUXKAgQfSVAdN+p1fnZYwdTjk7qmJAb2JA4CbJndFgCJ
oRMtgwa+McqRz1sE6dC0r4NiKRkq+/7hfAAPd5ZQBGQaXqiD5hXkrNFZqiPXPohr
bwh4QvAUgz+8fVR0JjgSHDo3Ik28OU6VZc8JNwsbl9innPqPi1hPAc53L8MmkQSN
1uc2jukYNJQ3he9jiSk2ojLLylbdwq7uxoHu7ilJSRV3HM5j9usIkO695qBkiXe7
DB3OIdEJr1u0vhtX1KaMhLNp1V8CG4TP4NZlYfHky3uxVU/6f8fJYVUwFPhDbCmy
nr5omZyy44sLf/vO2WMsEuOJKhflM6GWqWr+6YKmbvoEkvEupNjz8666mq5p7R8A
Uwn5kQw8Yp+qnVv6nZ4+TWlPIoygEraqW6Uxydit5x4uHi/x4HFXiNWPbcUPcXDY
fYh4MvCi3VX6oB+KeDpR3LgzSckCWWEVwMxZEQhGrXpsDxpbKiPXzTvU+7WbytUy
5HiUfkOKbVfUsjshaiUV6J/wiwvm4ftFtK+aWetSVrw897V049OUB95Gs8OzzgFx
fO/TTXTdaN5hgKtVUW+U7+pf8av7oz564j52lTwp7fvWAkbN0ODbxiIf1+1VInfr
+b/zUoky3Yh0WcFpgsGlDasXL2qMna+5AzJln0149ur+Vaz+0dhcYXu9HU+4BzCo
Qq36D1WGZKZXbmi/oG8CEZl89vh64RGe3e04HOFuHBnjUZXPuOGq9y0EkkM2cXZs
lMvBykUQirXeFiLhqPVL57Cx2RUtp66fB0+KYDCmCIlKmNUAWVLP9zESJ88GWYqo
liAvWUcL3XIIebcNN1ngucVsFP0mOLgxxuzzfh7KApQ6CWuJcmmIeGGlWL1W8cTq
I8BTabADcl1tZ70AsIJIdZE/MxMVCMundOtrIkiZTf3Qks0j2eeLT7EPKK8sI911
dfVRSIZThFu2qH9FI62+rwhSwCg5pGVFWV++5Xg91SAKReC9s/IwS2gIwGoZt6gQ
aRx9V1itf11YLqXk2PdnzyRGlfQ/kmbxzrbCj7VmncI0e9CeospGZRAaioVgI6OC
UQWT4rboEo75877hCTigBaS68xIQNwWiPx7q/5J0gZyeEJC9KABwQbRFUusfP7An
ENJ0QAtyYGRphoW1YUgp7KmyfonT0TVwNrf95G2qciVP2ovs1DfDDi+J5CFKZpvi
19RAKclLHHTauze5/WbWSBaBRIAQjMp069eB3pKT/U3J05may2iQfB4zuSdXqzUR
leuBi5sooor2Edq2EJjk3W7GUs8WILZQ99kDWM8/ujzZtMbO5AgBseJsE6MRZMdQ
btUfFrLkp6fJzwgzU57fn7ixNq61Gy1wUWrU1s8so9lSnYtdeRfzaHsRXItaXAMB
gW3BN8Gj1BIail63GADw5eXUamLwFuUrcvQ92skFYDHdtDK7KZMUaxxh28kUqVOH
tZ34fx585AYX6sPkJYIQpeKsAf92YZ4iaMUZKgNToQNnKf5eZmuIR/sKwGOtYmCO
lJ7NPIRE/DFdY2yLPS79gRS4CYZhFtxFD8XMgnRNcTxnIbMP6aCgI7P4qHcelUmU
GMHxwC16b/ZT2AwJ1ngv+wFRHYFhrsdMhhcuW2eBoDt5fWUCVHEjj1+mWEmOYN+X
QAaG6InmJ7houCWcxav4Skjh0rQBmEM2R/jWFnG6TZdy8zizpVrhcs0v+QZBVk7W
xl7aWToZ2gWpMApU4JzcWK+2yCRac6XYhMWlVKRlMNX1IByt5MLtOpoMz9PJkR+x
YHOXf8i36Uw62TJEZf7DPJ90dBFCyZqbIe5vLGyxQB+KexoYhGoj29pZ0poycdZB
5i85fE1OifrN2EZF5GM9KWxYxlu64v4pjjKll23Kim9VZE7YEOKA3AHKOcCHXPAf
9pcKOHWj/wpTN6/HFq1y/H+p+KHzeCdZnEg+xp/utMheAXwGCKg2/ZFkiYdnhv/L
82KEBdPlNGHvQeG95kZ9VfSmIwa76weHxbL24Uge7k5/56XYfvVbd2ZB+U0Ae9Od
nxgcKoeAz6F2rSp6k5CQ8XJ9XPAdxWIraa6f2UVd2s5qYDdpHaAD3GMNf5BkRRGo
MhkwiI/Ikr9qfQEZCHJ1Rk7LLEr3q9GlkZMN571dUOzZlazqoc6yrjdLrQnvXmBc
LexC6z/UyLS28VkxOaD35uJh9LfW2vIQV2QFaLYdx4DYiBcSU9X+pqyjzlq5OLXx
aZ3u4edIQXzXbIzrFUdw3chSKoL2tbHfCxVx1aURug+PdXCOkIQvyqgHJJA0beJh
v38TzK1Q8Yc9EIxxwPMp04uhLEJEoLIGzmIzcWQ7tXw8VaoIJF8R/4XjAGErHl65
XqxNLE8y3aMuMtJiSBuGIh4vF6yNDrQef4SuDsJgQauosVA27UbAenytaujwah9G
BiVvu0wHt9ySDar01r3KGNO8fXBpBPqyvLIfAKE90hZvEWnWSddygVyaQez26YCz
+7Xv/104LujmfwCgfO5HyUIqPzTKC+GoalwEAAlGcLHtiF1slI+DdODyaZtc+rij
F6kf3pavwvY2IMp+9+/NvJ7nnf+RTlJrGt7XQZ2eG26XsjE8pCyz7kJqw1wZ0sKZ
bDc2ozgILDmRJDe8nzLqauSJ3AmIAgFzDm9zh+b5vkQXE+vrt+VrHr5zUsQBE4OJ
Z3xtHdkvfKMemeSfdRJZH73X8JTetp4+Q5D2jWudVp5qTeW3MpZomJVpr5WPgKxb
KZFoVBdacA3EL9CWvaXfRlclujW4zaEpk0HMiWOjpexHq6vRBeosBSKxVfJ5JtkK
7uQE6ZuBLfiNBekEsc01Cg/gWGgABE/xFLdc7ELd3wMKWGNyRD81aF/NUhEMYOGJ
ktno87EfbI7mbHSp4/U8Fjsoj5rP8xPr27Z9xVjR8h3iwpMP0306vFcCqqzXCSrs
Lon83IQbrEDnKbI2nSFPQjQ/eILy+7Jd5vQSj3QuCEVAlh9aN9Txto/BUaFDFUc1
RojDcuaI862SS5Ou14VEkqA8uWDJmGTJGuSDWLaRJja/UKnnUjDxpw/lRs/xRgOe
U1w0u/OUqbntkGH3RryHVpVtxPI01cu0LeOTVpCA/O6IvN+WAMENI0uVvT/3wNYW
A/nuF9FdiY0MiUK2B/Fmzm9qXnQXgl3hTdDDzfstNnrtSWrIK9rGCh73gwDqfj5s
yqKl2Jv3O41LaRQeyBfnTe7Jl1NaDVNW2V/0pXngG/gv135U7gieMsQNVvNDgjpa
bBCzR4+LTX856cNvJqDRFymDTcRoA8T+BHW0QZTjD7CEh9dJ6LoCASC9dyXRaS8A
j0lFBKTHsFhzDA4lpv/O06Deo+Y/qeQ0yya5yNIJuyv85jQTFpgKFVfRocqLPCPx
jZOas1ioQXm8VaPliAiBtI487ie7MoTMDM3MI9OEbWtuMsuhTxr2PCFcxaLrReaB
A253kfLzL5YjiOwLPsUMPUfEIEKalJZoDiOjHfR6E2WIC9GCmAM13YAuGjqEzhvV
mMjmZFhJV9kfGO78Z/vNrkNMT3FhlTODV42g8PuwjmKZXEXlJ8S6zyiUyXQUh6Q+
vT8w9EntkLSCsHRCZSYBOXBuiExj9z6k1IO0h4mHDcU1tSWfxYWVH7RoHxH+Bugb
M0ew8y1+E6URZlNeMMBxIA3qE/p+Izrs5Q8N33Pu1yn9wRgP06zxzQLOljVyB098
S8+7nJ8qqUsho3pedNfTu2EPDgJ3TT2OWRKnjNnU9YgIAKv41EA7fwViRDwqIPgo
rntH2b6eWr4boMvVJ4cSBgqtslDq1L2Mr+JCclBqPuwD5oFC1V6obOLiW1OFW30N
r7NhaLRC4Tov4WayJBPNgUZDvIa+cPfdmDxNsG8aTZZI9hOvapiEOhceKPs0jVwL
mHgCaRVd17GaDfiGy4p342E1F3/A3BZp2zXZcmMFMBC11lvg79tIbaE5GImFftqj
eTw+AjY+qn3LuMj5HcMt0WEsaAH50StOHB3O6oQ39QeMnkq3wQnEnVfN7LUkGvpf
QIervktDdxEUKKW+DSKSvI9brY1olY1vec+CePq2c7KtvQAiNm0JWkUwoT/+FDdH
UBNWK+WSad8IqMez/pCbNbn4V/n7nyRqIlGJG1B2e5/6veZ3GALcIJWp9J2V8FiM
kHSglizUvKjB+eVR1ZN2W9aal4Ajk+rpY0P0avv2SbfOhK3rEdFXZC2phug5n9CZ
D9mrCM1Wbjp2WUqD02wk/hoQj7HXD+vDJRHl2mNQLK5hnF3meux1WZHv/eX3br3H
EXVRX9io5gxlKRyWxtigXTc5yL3JbeBIzNpqLdKtBpIQ6nvEJfN8LCJFFY68AAjY
bSZ9C93opGS5w2ThNapwbprS2OOYnNc89uvBQHokh2+GU8iKEv50VPJnmUHnYn+i
dPOsATXTpO4kSzCxgA36eW5PeGGwdkvOFxAojMnMieYoiSaNWiq3JM8epB1n42Ag
9a20FCk27q4+PbPoiR4WhIBrSTASgCnYgeh2upmyqAO2B1wu9VpvPKESBRmwzIFK
ptwmOQMXsCpFZ0BqTxaagCC4u1OqBebElc/18M6bOYVN3kDx9Bbv3wpv4GG8DTn6
G1RV1kf3tRKEiBsixTjOggeesNlqhAocQS/clm0qOin2EFuBO/LyCe3/MnLT0h4n
wl3Z09wDXoCrRIQPv0XPi8X3kis+VSup4K/tqHuLIXrWXoecE0GR5TA1I/XSpMDa
9+QusH+vqrIOdjbNmSgxcWlM55xRbLemtyXZYU0aLZRe9Hlp3icFPYaDdQD3eRNL
akkE4Zmf/Sd2k1qARmIp0WPGv5OpPb643YUsIKigl5FKolAul3uuYUwgcOf3WQL/
D165qZ6EAq/hCXpEjZ13W/arTeInMXINZBED8RzzjTb7y8QNN/yXrV7vHSMMelS/
YbiqVwaa+JnK+TK3DwzK0Vh64Rk7OrUL0crKlYU4v+Q5iCwxDZ9OIhLOsxwlAdmW
kALNw1bCkQEMpUtKLIkBcDiEvAAioOUD112I3srx2BCddT4WcolgTksA4TkpGuYS
MVr/NgPvpl9rAu3x2Ciccaa1WjIxt3iJZnQiOfR7RDFtTRmmdOAr3MU850h/4bgE
0QEs2uyhrmlRsd7gvN1qwrGM4bu/CWmuU5B/EJ67dAriANSd2JiHwhKcVaSZ+FA2
YqKhSkxPUMoeCfzYfRZJ7RlXp4Z8bm7h5sj01WBK1y/qKrXMgnGVt8eDamaGVhvT
UucHxJ53WKl/xUjUpNWlbYNQwiZyrnvV9PrYSKgCUcjWAGPjP0P5QstGAHAevn8O
d+1/XaqJ4RdJKasozwK1sqW08BWV8vWfaJx792/ikYXKSrpMpP9jqD0Rfkh5mVGY
EnL4hLyk+qWLGfmOjoIzn/4OaHhB1A3717DQ129EVX9Y2yq5unbFPoHky65gxXLM
Npk2P7/rW8mzh2cYuLkS77LDFGSaet4rGkqSbTKk3chJWHmTjglY1Gm/Xjm3NGq5
IHpPOaXSREH3Au5CLDOCwUtILkHc2XjEmCj4Kla06/Owvqwc5MCiCqI4zboYzBWt
Yow7bXCqnxLSBT8H7SU2ccXzi7LwPdQjTwQHeKGudUEyL/6bniS+CHbk5HEdBQRk
5E3L2R9auIijMUUFWPw9nf8jZd7qt9P6J1/rzYwDWeQGeYpzHKyQOXRXpkWKytcg
fb8FuWdqaxpCFQs/lKEKePJFxyejmw5su/2rjnaEuECDcSUqrBgcZl1ojBV8Vo59
+MGEa5DnVDZbI3Tcqv7QLFaBzjMdId2WWRFR6yD4KRL+tmmUL3e07wYwyznkr6KF
jIkf2mfbrDRCiM4nBNgEmT+gH+bHU19atHyY4kbh/AyhLdIeBGNc7n3UrbhzGljA
2PsjeVzEDjg+FTNdlhNxs5E+Dtvlk5SD1PypFmNrabaQ3YDgkvzANoWBRvgMrQCl
D/aP3pJgCD4RJJArgSFYRySBnYsmq3NxTUMH9LyzblvV0oI+q+aIyuL374q+CTbb
0f/3baBoBaaiJ1PJAukpxLAPUb6T/yce2aXGgdm3pUJMnCt/qVVA9j/UeW+DZBK4
KZL70lwk78V9H2F/WmnLlf69IYRq80k3goBOwP+5nRffUiCHod7NbKKmPQXp+NLf
7W9CwNYos3ph8hWlmjLICdqqaOS3VIJULR0M357/mQ6tDkrNj7lx/zvhWHgFHp1F
eKUnrOyMwS5WZZg+c/0nSbR1cwyEki0aGkeMfNFZaOqzauCv4H7Q2h5+O3aOfA8Y
/KXkYcKD7kUqY6pQt16/df/1iUF11tiLes8CS+BMJtwi99fm2+I5ud5UnX/Icxza
L5lZDhU1/HPvsofCcwh9Vgo+SDtdBb6DSIAeyDTPxoc0sQGRfeX/ZA+KL8l0U2rv
02Osw8YAyOqwMPAw8fpAAdoGu71LCJsQ76J9MxEUtJwmUInAntFHnQewFLUTH0vA
7XRp8rUTNbKtE3UVquIb7+Sc7jtpj3nnEkpNfNS9D+HIm970d/NdS3iS2FukGGn3
O7Fae6AGdPUQoniYeMv/VjsG1Xw2LQvZsa9WnN+Puy0ihgaXfR0xuIQMY+7Or1Im
7TMUMrvbaa9m7YhrjeSSurGsgvKrjuuhmLi07IAz8BhYtSjIrQb6PAeMwn0X03hy
K13WYxZHrdUXf7v7guzEHKi/tfsOkkVMJWLJUfeqeKoA22TIB8G8hAp3kaBKVRXm
q7Q3Klb7jJshju18dgIw7iGnkDoWKaxnNpdyL9w/Ak384vXdbR8olCUwgwoMgbSC
bcz2uLtMXoyfJ7dCf2UiI3u4ILRGA5v2JZZA+FUq3zrOcfG+uB/UkuKUJd6ephSr
gSfMusdqEwfL1t7OJbyuI6sVc2G8FBiQB/xO8n/T2cfsE2B2RxjkE5RHN7U8d/qf
EdJTLeHsyzWQLvbGRdH3O3dHHho1mZned2QXbiJBhhzG1n3RooQoj0t+0GZcF74y
IRyg3TI/U2Gi0d6OgYHYoiSj0sK8l55vNJpA8zYfids8mt3zXZviWuidMLoUASlu
WOoXw/xaxk4o1A8xE+TlyxM9VTO4s5x4EjPJq4CihZgdZgcZpCvajxckPY4uomLb
Exe9wF/pczUA2KxWgKto/DgvxjLBJ/Jo14Hqki6MApHjgsI/OXIu6J/1ZWZ1O+z1
SRQ2G3zLwpDXwk40A7Heb00DEoMO1kogf+voUhXQetoNwBTsOA71FSBCT8Lv5ZPi
Bf5aQdqiJWCQoMvu8fRBiQ8lcD71Ww/LfX15Ss7JPnLKOSPlmDoOXq3XT6tKymr0
Fl5QVzWrzrM3gGbffft6lWaVwKhELdIrGpE94eGLtfMPwbjIwfCl6KvDaqmkLofl
u4+Wyaycklie+wo97EEScIhZ+V7pY4hAECzyaZ20LtzUPJslWsus1n3Vtry55E/x
1xd6BNwfD/v9et3UGloRgEB2q07YpvtyIg8pWFoVrIsDhaqgMn/M0hBdOpQyLkXa
STziyceneOALY82BZwbvzML4OXM1zZUEWkOAam9/+88WspEmbZzeoAE6LpYVHArg
ORl41eJ5gbcVOvmfMzFCvNQs/ZP5d6rhMHAr9EUuY+foaKGa/DlNXQkAjRiQFBj3
s7wcIG32p0634yNmHc8xn6MaYhy1aoJ+7PuPmoBrcIbePGNCkfE3gewKuG0VFv2Q
AyQfgbdojmO3asfMFkL8xsXXiVezkM7q2tpoJkTibvqCAJmn4DbyK20uhuLHuN63
rketS791G9Cesk0Vwl4GbHDvczotJO3eWW6de7v9VOtABMvnRJTqYr/mxi9Ntheu
CmZtvDppS7pUcV0XI6bFoBEFlln8YckQo0E3t4fRLzjxqltEctIJY2MgotcfltuG
J0kFv+Cb9KE0ZX6kqqREsnCDCfY7ScB6RkmuDE0SCgIgz588byo5Cc5Ne9MMEl1D
t8Cq5WIrdZGCWOnRjr/9MP7NdPh/sDH1yPiaKZb3kJ7O0/51HQn4/7QOR/J7WPF5
uS4e8odvrWRIvCu01RPJfPQWsLVt/8eyltm/SoldHy740KrVe44LFGjF/rAEkv4H
naFAjyC5ACfSy3qjB7kSmRoV/slLhhZEo9Keu2Xr/kEQpzz3CeDk/mPcNTeGDnAO
ZygK1udgkztHswHBzA+oRHCa81zKwtxdxr/OMBJie2c+dLdv+ik6KekTrQ7JLMI0
SIBtr+XYp0Czv8pO87Kqh4bEWLVMnObO04wh7bGGshyWREQ6JXhAVju2ENsAJKWQ
Y/kuqUuXFTFUxks3ADw7sg+x39QgXrHs+2Toi9E6jUCndTz4TjD0rBOEUf0EOqTu
DztoenYHH0DkKshGwHGPMAYSQKKGyguv0N4m7S2xtYBpPXW/+q7CY+/OOagBCvRu
jjJrN0xkaNWenZ70ANAF78qSRR3k+7l3YLEgx2mxH32pJ41Tjnxvw1RrSZsQOb5N
nK6y++ETTxxdhY2xRZBaMWXiVvHBpk8FAbyO5wKaJa29/JV0QtFRyk6QcCrSg75e
tSRI6gNg3zptWtvyyZ58y4faFt3Kn7jE26XcCgVIXHAg/Hp3bvZucNe8WpAi0sK5
yescUEhazG/Ymvvdnc3UuXS4qtoTAO0JhyTXTw4VSCi+5xEV0hUOJwXJPCYNhGen
0nXM4eDtdMyz6GSxpo1XML1CeKzlpGKScN9OwU0fNO4aCox8uGxUdrwLYglc5sVx
cAGhJ3JzSS8TewVI+F06h+Nk7UiknxPIrPLSDuaDw3ReGZcuKH5SCnZ1u6A8+npC
qe6kuO5bgBVAEDemIhud8NZemidoOFryp6RYXuDqmPivGB+fALZt6JSVSGv+bUzu
aTPjVKL/AXA8xk7HsI8R3oLsX3kKdBtWewWarci1FLKyFXoLvs771PavwAqZS7gP
3W1EWhfb6kHYyda3l3xmXFifxFru24aVmrZY2pO2iZOtcm1wVtvWCHOIP7Vv88Fb
YfywRw6cJ83PWw7GwbEgXdbbj4i+qnabU+y0lxPTSMezoqXdcQ6hsz+1wtrxKPe+
5/CX6YpPUBrWjpL6rGA0U1A6n++fsMLbs+HZknrAGdyCK1cugCKO+/U5fyqFv+MD
eJ4TEfXHo/MnjOxDPdMrAFQurCgLNha//w4mj+RekPFmMY2KWu5UH9TRWMaqcRmQ
IBtQ0Is5bhFmZc77vt9vIwzMtM3cjXlCk+gxHENtuYbP8dk0q+mbH0eUE0g1cVd0
GbXPmoW2NqiVTCRH0UBEE9Ujz298Sz8xDkCxKyIx1lWFwtMLuWna4GogpyvJRUTh
FFdGyuRSI/Bg4LnbWGMozDdeYdTxe1RrwbUSsC7k8WMWdv77K46L5FKE6Z7IvgCU
j+a5hd47Q/2LhkhwkmnTQhIsqS54FmjM9hJzgKv90wIJk0Q8Pl8eWnfARFf3EJVx
HQLyU0djTlPODjXMmcf0Znzt19prn85t6zI1BYdQMtLxUO7ZAShHQGwxCjQ5ksGo
oEvOl5q1hgzIxTxEwcT4+Ds3nV/gyNiNyDsYwYu/bkuRiELMq3+RtQFBpph5pqR1
2//vCvMArlaTPK+HxwcWGYj7WpfbVSS2vwqYplYr2QbFAz0Nqzy333xRjZqYTNpK
X99E0G34qUMbK1F9Qm21opocPVvinOZzca9iWU+Ifa3aC+1MCkDICipNMTYjJvCi
F9MX4yjUftsZhX6jQq2FMj2oR2RNwvmV92eLIEx1I80DruaT0m7xMwfGuD5SDEXJ
TwW4elBrjj0yelfkbMb5d2bw9yr5W6QVT7KBTLjbvYMp0c6nF8C2t7Uhqy50HLkT
TNRNCMv6BnYNkE43JahhJUf0YfFLGCBwGC3c02EL1w4FA2KUuxYqgRfW/zfpiycJ
2X6D3e7fyqjPKMTzPRrOeJTK31YfRwnHEvkO6dbHj0cdjK+Q3KMe+kWeIm4DRYRK
7z+uhtswOled13+2hema1e6ciYEofv5K1c2lEv78Od+AP9xjGQlX0WMAGPS/DuIO
6sEUcqwG2PKOESZIYn6hVBRWDWV+W9oRslmwsxtxku3NvxukxCltSxk9AapbtGYU
lFVGHKAOcnFy0U6G6Jj5twcOxDsOPHpn7R/wpi3gOQgLkmTlkD/boLAYScMnLPTz
gaN3y4SUcuwpvPlsEG3xZS8h8TrUujvl/bDzVXZRS/XXw5XyvG7nQERXp3o2u4XZ
Vp7xh3RIxfZxnJqSzZRzQMQ074Veq17tPW1/F2nhzXNz8wsMf08ucXF3xg8WWfcq
JUgabztfknAWsMM4Btv6fD2/NZBzpgHc89h/UggMOyWko2bIUUCrlVoT31xCCRVi
9SrGl05NjyY+zHU0Gswjc6ssk7hY7BJKGlkjBG2LQDwMUae6k5bMRcFSudoeA6V5
pfNudjHDbPv/EXJKiDDkpcBSpAzfAq0B8v2sNxrzYqVi0kJw0lF3C2FXlGieLjvj
hnPb89dcOefI2Lwr1kCni52Plq7SVvjhvbSg2Q6Zw4k4OCc0LeFu2n2PNO7sP4MI
/2uL5/wvlpHewKqQp4pOvhvU2GEuOh8dDsADY3snoizgT/zcZMtbwBujwednHNqb
N1NjT7WB0hTKkxsY1e3ZUFGoCVvnrUY+aVSguc4y5t9xjBd/RY4Qbf0u2x1Ep9ws
+qnnPv4VC77PXki1Ds7uh76Al3EfrnM/7Ov0GPEX5A++vsq/ex8tivnNB3RClfhD
1E0Qlsp3UHbTlqneeJr4rOKYUGmStRjIEIPMj3ACe51ymtCkPlgbsdPGZgLPZbDg
s1/YOFOyYYzwXHJ5tvpeRvoU8M7Yp0h/uiSCfDgr29tsnLCap65hE6Y7cx3YiBkk
PDhnUfyRcwP1ZS379AwoZWBkd22vJ6wQfkt663qgE2TOctx8K3BUa9m23qt3CA5F
gx3nwZ1Nbtx7zaKgqYFK2Q64D7OLS15WJisETEmTv6oUVcKeQIdtsioMZmCs5Mol
tRIDdIBwy3kRDcSESIPF+iMZc4DncXMrV+uRLaGbOPQl4fyzfBougko+wbolQG1U
cDKW09L8JaroOudIZLJI3krdCCS6ibU/sS2RW4Q0JEKKNkMU1B710aLyL08MsU0g
Pd2xwVcoDTZXun53zLzdFIhi1QpMnWPNyXvbiP4M0aFCKi+9lKgc8uCBqhwiCKBw
lXToPJ01wATNdxw+nVa4SEI45Sf1JbUnT9lxsui2JXsdP8WU5sx5HIht0saOtzII
qdMVD9zzjS1mHDvFwXgRPH3rUsimgfBjx8gjYN9sOAEdiWFWa2L1DLUAf8ZOG3Oi
R6GVvw/Vd0j2+8BR/QhhuCK8lV8+vxDPf0J1w7cRHJhYHncHB2VenFcjnnkt2d31
PO4XmxZ+qQuXMwnoYCVnM0qb1JeBA4BzWwZI9Rp+9kHYXn8oIeYqyTszUN1DJYRY
QXMhlqLc6HyPxRp2H22Lg57dmgNV8eqWDcQROPaWBWtlfSRSb256DFNmwUJDYnjz
po1ZBNxlZNWBA/WoAXiaDDx4OF5zpIhWwJPyVohy/Y0wwBvUhtvZOA9rTTWDnFvj
Ss9JivuLtAOczOMiFDaMetmOn2Y+1bcV5q11vUJ9lNGLYILlypjS939pawtJRSMU
8NyzpmbfiNZyddxNh4ql3ykSlaaWvpfH7fFYTxj6KrtIrUHS4tn9mBrB1JzyXNp0
j3jQl8j9SGCUpKZtv7cO9bJn9+6pWSDQPomcj+xReQQing/Irm9dwhad1TATLc0T
AHp92o1G6Ftt8QeHhbSfdH7e4zR+VXSSdQUQ3tmYsURC1urdh5nbqcUqsXoyLrv6
L2QrqlL+uHUYcLGbgCqzz0imTJuq+KyNXGUjCXd4yxhdQuYTT8yI/SnFdu2cHglX
w4pBKGv4pP5UnQ0BkTFn0phU5y/0IZC0XfhjQQWBEsuSpjfIKQ8d7T0px7LY5iPm
EhVU/u+1Fw33kUTykgaS2r3cfJ4DAZSxyv6bn4FvERSM8qcCO6FdlX0lfpQumY8H
0UyWKNGzKyz7BSZ8UHWI/MgcKw/iWUykDUGHUWJ6UNNz58Clb26DaACupVuDbZjs
j7u7Fzi2oiPYRJtX6UkIl+v0OwokTUxq1D/Or2NmeFPWROVtLfikqSe+fg3/fhmE
3C3rktmY1tHxdGoe2V/g5UzS1rYGMafBIJF2PLT0uAsnm7VTnuHqJsUAPsyMJlSs
fDTK/GXaNnD+EiVUzA8rR7K7KQXStM2OKtjHb639ATDAJAVe5mPWdp7aN4qhfJbo
RO+TEmXDRO07J54qW/7bGhE5tQTGTAEVNXibMG4pD4abarn7GF6/ovuYHWtgPwOZ
3BgylsOpymOfjdtljFFXEKnb7cRuZUfRDVHLts7qnkQPmxa0aIfYJRk3uUdIE8nD
0AlAkU8J4Nz4b4SwmKZiOfPiPBQ0o8Ym7DjFJTNCsnJDZ4Vno1qQYMpwTuscGX32
faNehAYHXRxsGhO16/BhIm7xGITdA1KKkjXQpCnXMKqyLGd7s0A6pA3AHVMh/+oT
0+sjyM0pebmVlMJcFz9Lzsb9F8YpVUIkTlHYJWcJ9atGF+ifXrJknBVZgtlT/erK
TR6dbSMptxJKByMqhfu+MYwtmnOBZhdzCmcPy8wKZPHz3MScl94qXKFg13QNNl3x
pF+ybXq4jwK1SSoTZh4xzIsIXv+OFUsvzh9xt2NSKFvmNROEiGef5PQTpq1wFT9W
4XxxbKVf3ePZXK41Mv1ByWFA0ESxo/83R4K0aD6u9q1uDJdwAV2xK9X+IHh0pRFQ
kRlzS7YySaCzAYa+0UQgW9lHio1hahLa/WSHaE/QivS8X1dqIQugE9mBAsKwLe3K
WVS6TP7QVxoKgfLgkjUbsegaF2uuY+LYMNGnx1NJiMgryXIna3jF0XX7jrf8wC90
c1K3PyC5OmmCi2kDPMECvcdJbauCfgqhvFxDFAxqHbUJTftz386Htk8fYhy1zmLn
S6+GsUoSvj8KtWAVIUPKR5f6x1lJ3s+DWLxiWWjU5xmWtswIsMGtWrlLTqucCnIs
cdbHkBQM0J1FFYb4J4x+jWZUsVtbRewlSfJ2wrqKbVWF3UfhKCYaOIB/40H59+U9
ZeJEGQr1EvTXdE+0NGlzZl491MN9WaXJmcEAr1NTPS4EM7l35LDZ1J6EMmAP6STp
rfWdFS/1/pqOJe3tkcGwwHukfy+Y7/5jdsNPmRglz7xGE4D6+4cei0KDJSZnVf62
1ELTJpk4QHpWHKzNpdJmF4/jFRiBKUgrZbzkZVDZ+SYTNRyVV3xgpJdjGATMQ5CQ
U/NqBDnXlidKJnqcTa1S0RuhKb2SOn/jopGTGl0Kiol9Sja4P6ukG37xf7hrEpM5
Z40y4aJyTnrB8N9qGbdba9HRDPEQNgUNgbLDzofOypnkhdJY0U+QsFMy/kZjREFy
mK3opT8cxDjYecEc/R3R4PUK5YGbqAcRQ0eNFiI1gFxp1QUV+SelTo2Xw2YEkVyC
YMKOVtRlFmIzC2fQL+XcN920k4GXOfBHr/4ExI0WnaYehaH9lrEF71wvrY+8Lxb+
VZ/Rmhu9uJw5O0Nnm09sa1HrOhT+CGK4WyH9cYhw7pHXhPTaThH34tUXT2U3TMnd
ydnD8FiO0pEBLYEKlcHP45cdluIS0uNHerTdoqbvqNcWAZkGQ0u3YgO8MQapBHLj
2q4msGaUT/S8ZsE76h4Gdd76TbUFU5yiXcPC/xwmFslFh79LI6H1Z/Rqhc3QwPAm
E4X5hSod2DNwNU7TKhhMbZgxO57Ut4Y0w4PVXhtg66PNfDTdvb187oUQtFZ2J6J9
nQmwDva2o+WzAoINOYYRCrGsGWqh9Ik/saIZcceqhZFN69oBynfqbv7qa8Zwif4y
+Z2kPIjmDp25NhcTdLHdql9fcyooDcHcQUSDVBr0DG5yDVsrei/cuW/5Gb4A4ybt
11reY9ip2bLuF4F0XIJC8ypuDakijxFSp0Dsx1qfGA74vdm8RSI+Z7EkFj2jFDgd
C3kDFMBeth15UEjCiDZKLOfserOzGgiP/8CBa20zG7OnUvodx7NVad8XJrwH9wC1
ripiB2IkOam7WNv9Id56LBQoZpdx0c61IQWTe6GrfxOU9KHu+3ejY2HsMkw3eigT
cH2Uc4fCQwOJVGhg6WDvSPKqgpu353lij1eZDjcifa7GdcGlNGiA2nzJI00kdwtF
n3rtk4VAiQr/HcxY73ZOaCwlJdNow0DuLo69UoL3N94kMuFtpXHhNmnqKmGZYgXr
9irXkeCNGZP2ru/m3Gw06Dkl3b5URhXcv9oX5ux9p/GEL00LG70T9i8u6M6sPvUl
tQTCSvtTIXhorODnvNjYKxNsqD/3nU1AFqvfSOkRV0TOmv2eXX9oDxiqRzl49yhF
tLXlEXYAztASppgWrG+9CJdmeQ1u7XsxvXT7uq9cLT5WSxSN1c0s7Bl9MS829G7t
cGlcXblMcO8qpwVbv702TUZxxknlBvz/jjhfItXZgp799LAwJBShcksnEkAmr0ls
IArGm4ZF0NaWds3MmA0yTd0tOUf+2+6QTnbb/MnJbDFXppqDxGyZaMqd2Sk/fHMT
qMwe+Vuxy7tbtItvZ1wbvgOREvT1sl/6tKbwRXApjQDnO/omx4/SzI4tigVzX2yJ
UevOiJAYzOFepzMzr6+oHgL8EUbCQ7Q4bPu7HKU4CJ02Jvjij+OcgsKE4LbNDmQm
tTxwS15k4Yvhskp8BMbs/Dhrgvo1kcm5SjoHRSIVauLJ3v7hlAIbm62Mgpe4agW1
/EAnEd1fY/ILrK4EKP1aRoytx4TmzRNn3a33xqvHCsfu5vsE7BbL03vARBw9S+QG
1fcJAKRvwRRKkk1BKxshIgooRLQkQ2kJVW4OC0kJikLVjOvI4cjTiPSwWdRq7ceW
oCAKpPAwbr08irB7c965TM8p4mAK34jO23jZuaJaoIcrC0MWrrf2ngFbsl9oVc/j
7DOhRoe+irTq0Gkk5TZXun3+cRj/aBS2CNncVzJh3InlpcWERpqRb3irkpUZQH6m
155+rQWc3ASwE6S6w3dKyj9rc+FtZbaSMMiOWzwk1YpcBAxSE3Ly7hl07DnpW0DV
Np1iRB4C3E6ma08fr+KrjstWCgaKr13vpAj8tl5ElGCau0pV5fEQcRKQZMSd3vwf
Xz2sIDzgepKmWN+2TIYmrSIdMjZ3I0TOZR726AkADwL3z5gwE8vuD6SiPdQ+Yv0I
PmTiMtQMxMlvCANAOSGwOa+0OG+E6sV2S3Dv1yWMSJntlDq2AN8f5mg+GE4I5Xon
oVCYMwofAg9K5WneKQJ9ZBIO7hWByv968Hz7m1McazXGf4DWuXu8Gz8RkUmYYzW5
0wR/aWiRyqsSLiSflYaFAm8q08AdY8mmqU98z5hKSb0FCzlz5UOA+6DNy3hf6mDp
1vTpcSrzcRDFtfLDoF6jzKTN9KtyUTFAj+i1Ghc5BKOHakqjCNkgGbP82njVRwhZ
QL7CBTnbdJA6+wLLldvURFnjyUQTCDlI2AUFgL90oUsuF3aopeFQcs3Xq0aRbgCM
FGKVNAR6XSQ4MFGEob7O0Pi89qV0PW0oW4XILNSegY3V7o5tWHTuQZF5AE2Lq7Xf
M/GRNRfQhV4TdCnOVS83AxBwxWPuQryfygCLKhZrT0I62uKAXb27n38AZTzatcF2
9IDFMES1Kks9pUyHj7n+9PAU3vn0+YS86foKqWQEI+x0nE5NqGnPCe1brE9tZQe/
qICelBcMF3wMH9JwcfARD3H02H8KeDPZXntKS2u8HxVqGnMYz5IRXq4EQG8YGLVQ
JlDf9z5/cokapJ5h9DJaD3gGvRo3al/oDF0MPJUxi5ZXjO3lazCqNfjspxOVU/G9
Zl5OfcR/XHh+7Xp5I9KTpv/RZDZDUPR6GDx9L6yb/B1qEgJqJ2rajUsHZ3YkshdI
4wBaL+z7ZzkygQsYZJZlfFRYDz3RIg4WUsefgZ22yBdacNWt62IaoT9pbffIZMTp
tpgUhP4ooFJCeaN/V54iryZ8WEAsgegLiDoLtHYJ9D+4RVKmfLa18BUGb6ILUUK5
/uYXtzRM7ZidVamThl+ZQomveHHEI3SYOQLK5bBQ4AgRiA9LsAdM+LyYGHSi/LHK
XU/kQr5FfPgIBT6BqwM7/KnEPmve/oEe14kCrKaOke3usNfNjUnnKcLUO0frygL3
bH/Pm/oceBIaPCjtDNDm3gzzxdO4HZyqN3M+sheH1uqMHQg3UAYVHb8LcXX/wWET
4pbQV45HBRu1Nu2FKSy41OeI+meuFmjieZ8WBHiIZ79M174GqyWw5WK2dXu0+71n
R7YeIOZh34PtidQIE32uJr/yJyQB93DPwYtbRBVgB+zKAmPoTQSHgupdG1hBPkBT
a4ma+zOxU/bbtzjP9da9lSbqY1YnmERmYBUQxEV0WA2prCGfBbHFFUkOszokRUCv
fRMYVFvxg4wgKOC0zvVLZEpZQ7cJZhLpkcAgoUjtuKZlIUr7UjwRirL9f26T913t
/X0wXiR4q6Ngkq3kNXh+kDSemFlAp7vNEruYsA4SGARRI9b9/3ZNEJKP7wYV7zUE
JKabofTRTOXOiZYRbLKVQ2OTDJuo+nxTlmdeNu+xr0UcPT0130FVo2hlHjCVhYFU
fIuTNE5IiXsMnBS2zOMIgeC/2yLaXbOrjpVxwGb0jOPm+tniyimy8efLz9Je2w5A
NGs+crl3Bvvo0sQ8w+cKjYVXf2hXo6qa515QP+JChlEPcFkR689EZl1W8GebZak3
pb0HtRlZWzxbwl5LNFwPAPGb31vonzS470ffk4lNTyzQsYgkXakXXVpW+5uIJGiv
08Wvw8LnJZ14fgGkI7Vupcfc2BmxpWHwTtS7w92vexc7gLy5fdPpTr44h1ZGU0sa
y/evnZ414OINcXuOiaGKg/XXsmlPj0k4dpREHzJntTItjTOP1dj1nXim05YqFWHJ
xCg/LrIPYjqaABN7Wtoi8pUIGa2erfDFKJv55X0wMMvEzDjb69MSwgETwBSr41UU
asnxe/d/V7bTyI5eLA/9I7U+X8dGgfLcuQrYTQQ2VNpAFOjdHoe5jQvR2fAZ8gHq
K5gmS8GwIu/ji0VnJq07nol9RrFcgN/tyTdhyIoau/AJfgxo/g6tb5KwjbEW2nZT
DdXzW38byVVPeqzPMP7/MvQz2+a56Ilf5lWy5+Tx2GZae+1Fqw92ttkznJsKRdBQ
Lva7JE4gW8RcX1yvhBJf5pB07f0Hqoe9/Db/2gv9nFVhrnpGr3wlaH7NiEfMolKy
6/9AF7TKwDseJLArCoq0Od3X26H6nh52s5SrV//fjO5YlVFSML13sSjdwpNr35T9
ng+eJqrKwdftZeIjmg79zxJbAsi9Gn52UXsMRS8jjbBwa3G+s+s7qGchZv4+iU6W
KvbaKicHgNw+q/F39qfZhxPp8TWGnk9OES7cvo6cCyn3BPb54XG/dFVvzYXbOsOT
aLT26J81uiSB2a0CRD7MH24qJ7cFU2f/50BMwaeSugPs26sTF0EWYP4v0u1WYPp0
7w47Gai1UXwo87c0OaRu7Py2wyKQJtSMCQqi+7E7KX08rlxHA5LHCB8wLdcSPjFm
i062jugpzh5TlZ7cZyUMy0r/s64kxkWB+NbrpPPKmCf/YugEEkcg+xOxGXYZeSlh
dZ5ONeHjyCZcApplN1qlb40k+tRdumDtLbvq7icjio5Ce4ZHlBUPWaklFleCNOU+
Poi99mHj4iuX2FV5H3BDxKWlFhJtv8IlO+7IYKwv8l8zrg7KnJUFXnqp9MA6PXkB
HLPvANuvSlMFSlflwntBu77SaZak8KhOA2pu9g3KAtxEL4xVv7E9NSkGuNvRtymW
rlR1LXglhJf4MHRh0c6OO41cI9vDuRtWLGD+SuJtFfZRq3tB2jT00jjIrNnlawbb
q9QoUGImx5y5Y1UbJ9djNqq5afrS/Z3Mb3Df4qpxYfHwrfjXVnFXoedRJMcgMybW
ZXRss8gkU5nlAveNbUBMMhPSPPxCB2wwhz32+WMLfYlXYO+2co/yJk9gWW5T9C0x
dIavCvMQCP/OKwwX6Jbjn3KgVBweZ292Eco5+WeetyPQFIeCtjlTYyy4bRJEo/iw
AW5QLe0ktemqU1eNx+KxHHHJ2MIQKqYkpxrLsDf1FOJXn81rcTeMg2Ep7AQtCiAw
L3PsW5yiHpDGL4YYt141kNd0vuFX55c0V/I6PyYlVJAQo5EUAPO77womAMuNg1Ki
9eZuQ5fIwp2PodG/RGOYo2+Z64guac5I1LciNXDCNZV68iNWaUchQ1LM7CtD6vlg
V2tzeA6b7H9WtXVuBoxxOWw8qM3/pJBIThkpccqT0OAMJoMTnqN3YiUzbmPHam8N
DOXTkJjBWyoZ3cehuSkFqcQloIJrlT2Gb3p1TnLxDeyUAr8G7BN2EVVUOBHqOS7n
gyAU8nk9CqpLVyllOv+5gsWOs4ePMP+Aa4V0CHvoXWxgkLec6aPOVyD8lnBj/2C3
HZG192QcTWStwZEjc2U+7+Cja0fWco/SxEctQlxUC1IXmUz6sJ/RSTzBCJqiwrUM
RXT50TBemq+XWiIZIdMHzDqFqKc9WygcWKRiFT7lrjtVH3JmLhRgIvidQpr/VbGK
2sVE0p04dixrx6bp2Ez70Q0Xt17oG3aPFiaww4h+YO5dTnsTuzR3gg349t42UFhP
nhtBMBlGFzLPAQUWjE7D1nEVA6W4uBFL72mHW+dOOS5R2eFRzlZ4/wAtSkaYaO80
LoIiDCS3FFRHAEXL+NQ3rlF/kcrIiGY90uaYT2tnnjG+VgrOO3YfkWSSLyyBeBRT
Y3remZvvSTlRWyElMz9e6kLHs2UiOCkSXJBxeckX1NG4sV+CrkGudWnMIuWKjTVC
NDNzbRkgu2/P5mhTHX1HyFSxY92jVP4Hst+v7o0dVGpu0ixNND+nOPi3osUVjeRZ
5dUjQVaA1Ob2PJOPc84k1LyNvW8eLsbD8dY8IahtOQc1DKS5dxBibF6w85Vc68XV
v4unsxoKneDiHxD9Mx+97Zcx4WyenzUskYFbL6NEq5PsimZ+JhRaWN/fC86+QArl
d7BvZDCng3J9KEX4hvg03s5Kh6d7WFnw5cgSiltb7c+MpX0blXwKPFZ95K1pkopx
SL2aWtaqIjpOT3bgNVP+2b0HY0wEsDK4AeL2BGXFiY32XWD6+JCTlcpLSj5aA0f3
dcr7EqeXD9hOu1lIb4a4SD4XVLhr/W633x9r6OV5FnY/ancZ4WJR42yToLNrHyoQ
WGtE8yBTLZ2ZYnRmBkaUpb4Uqjb1c3bdsP4IDNvJpQE+40YZvWMTudIvo+F945ej
jUXFdydnOYZZc+iqp0EPa4GLeoZgizSEMo6JC4LJ+YePNz2TsMlDGoIOaCvNtuw4
KTUQbe/5JS0CymvJk2e4mXLDnN4v9dm2FfLXRUk8diljQi/ZelnpzHouwFdn+dc9
svLGi26Il/WSnPZOTtUgLd8ye+KdX+zbIHBgjeLDRRr3m4K6bKVkfipycfx+im0F
6zKgXAKr0c3pLXKszOk1qUQ340XSs3XLKe6cLXuFVhLluSNsJUIPmrzoYqVQIMmk
w/IaCTl4dVCDDwpbUh4Oc1ap/z30zN9lw3lNUL0amHPejsHRiM8eGT9/KkMp/HcL
re4obpIkGwuAZJ65zBokMHtCKlf638dEWmTz87a69HR+gPaIA3Qcurn5N4BFrjjg
7j6nnRlNSLq6yRZ4C2CCq73Iol5CzhaiHibXqcQ1lkf9AG0G1X4m3JQw/Ff+XOBt
YxSOY0rJxOMl/0HzZC7fmGUIY1PfhssZRrMbi+N9wu4aWkYws/STYzYisImJb/rf
yDeGTf3HQEzeQmNxnIQa5y9JqG43TAm4XQFDfby+oYvwXAtjwWTJUzLDmvHhLxF5
`protect end_protected