`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20704 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
VKWNRQF+vfUNEEp7apOJOYZ+3DIAZ8xzuX6OZ0zKxuSpMu5/zkUxvS4vDXiRCFct
mRR1HpTR85/1VANsjfZvFVuEdJjZoD+nD7pXDnxeIcHWRmlpTmyV3t74bOtKNZ1I
ifI1OYfAa49+kD3P9Edq44UdjeFRIKko7kbS48E+/+g1VE+EmXp/qbBRLSeEZj4j
JPNr5IOybJcfKBmAAWD6CmR+Ll41PpxFFk1bjEoAHs/7kq46906+yYEArkMSiu5a
NFHvcUvC01Dnu8tHUhPfjZv+Bjcr8dMDJxjmLn9Mx8I0HNPm4Lp7IUUSPxyGW2Lb
TWQKaSjCn8ZMzrEviIyPbCiP5ZSrU2xyalFxO67QdHCn8WGCAaPMDZBHGxhhhO96
qrCgh6qeeWdqJOk6wARe4WW8WKNs0RyNGsW/uhFvaV6KHQ3ldeqeXHH2OF9SCrGc
E4Psy5e5+u2TxSj4+GPWHPQM4QDJs06HEEE83ZBddYb+fVVls2Dtk1SAnvLD1jfb
49MyzCJkj7bWkRC3qdrVZYH5rHmpDwrBuVac619x3jsY8lh7RcyQIiOHbHP0HUz9
/jSBorRCH6f1M8WSiF0wf952J1ozEkvm9gKRUNhosQRBckKfKNVOUX+G2tM391Hy
1eTzcdxu8INQPZF89dgCp8Vhf00TxxLcVtYzh+Y2IKN11CgcEttHF8Ys2uW3g9aS
+pLcpduUviLewlCgTN2Dyb5Ye0Jw1krLt/jgyrZrVDzvG2Ej1gKPYx17XBq1daQ1
uX8MRtp6XXaMSUq4dBRpXdaG8WFUM6XCoW8L0GdxmN18dWjKFh5AorMUpSb9B7KZ
uBanxEvrapYthbO95I0rzskocF02KBGmtKTffv92qybWMJOHHKGBwWfZx4WpSmHE
o8nUuNbQvbocW0eJL/P4lyRAG7+a6s4WZ2600DNyjV47bgDC+h0EYz8OYXT8K/4b
4/R99iQGfIjAr73V+HAa3cQke7KkKB9nBlnfC5fbTGCDWj098uFyqYcZooZLyNZh
7UYwKkQe61sCpBlkJhC1uIEV1dzNMEes1WstkiiCZLRDt0CO0GhGHt57JqwspSwl
cABVXm37piDYtl+RfWztsg/0alwEPtPz8ZapXGSI6eFUyxK22MwR8FjkorSX9UIW
jCiVHrrYjm70kBJRnYxnEIQULaSKWybPV5NtMqnbQzJ5weeSbHonK4mx0wEcfyCC
IL2/AIv/mAFVdp3J3EUzO2yb2J0Mr+xJFHK7wjA6S7Vor2WDauHzepFjpnK7Wjeo
Lyw4Gje9KsF7YoneBiOex5z01ThXwKpWZRQ3X4CMlMrKHtou8TAyxe5M4Gd1+gDE
EuNaYO3P/ZHsqZtpvOVOMhLwrnEk3rlPk4BWMwopCIdG10u/xfASHESmkJLq3qxB
xXu0qeP2QAcjRm2TO8iCFOeJlvTbZ+fXT5a4CD3aYf0scVBPn6l5HnZ4w+LBjnOj
FrUezISj1UgwH/2tAEioIlv1HisbDrvbN954z8blPwVVXzCfLGZc3XCR3VkNKwCG
fshbTEZVdmPK4khmrYMVIXdNsi8cXrz0nIfAJ7ybdKcfOr90ovzgQhfZUG888VOa
/VHg+hYRGfpv8Zld7WUFCEwn279nEeJF4H8fbdsVuxWiIoflTw4W6KPYuonXV6GV
X7UofDwo3uXqMYvvr9ebfLHrCiHRj6JsuHre/gFWL0z84P0ZVsIhWdE9mxlbsAan
zEKb5paNEyxqf0L/lVXoJ1Jj7cKgzwue5yIHfCSFpkVkPTOdI1aGqF6jXhFL4lMM
oQMjF4UcRE1vYhMYFB3xUZBgzKDZ8i3nMk3FNbyg7tdO4DsXuf1eXOoWWdXIV6xp
WWDrRbeCd5fdVGiIow3Z6ArUfqt2ES2R/X7R6XbhYSSxFWfjYwiRYjjV21wLU8U1
qxXnpgY3GCdIhMG3xJFp6cEoLHXa+ylUlk8fKdvTrJQvBkNqIRRhX38LUST0zFAT
49Yez3zhRqoln3wYM6YIuWxEGUaMttsW+s3/OxXu/VwtZjlrMO7oQwmTfiJvGys2
TqrVZdcU7VEwiqBM7W220fhEQdG4N+QXYG/p6wr6BdRn9BFDsQFTQMJxCagoGImy
wvMwfwegBtJiAecs6tCxTU4eKybnd2kZOpaDtTSkpNBiM5FB61RXpjjN1W3l3WFE
XGx6ABwW+zR7f9UgVdF6UEttwZJ0nbgBiXaFWxXf36bxHqBK6LL4icV8FhERrkCa
Mc8wUDjXaLkieN08yjBx9Q7Q4ou80R16StFdFBKGOSI7MFQ+ywJxwlN3GtLkmPmj
fzAs7yYzVXPzVwFTl7jlfYp9HxOiMlkkT2YeRofEBlE7kYITiywnF3R+JkilSvzc
aVL22EVlpZxQexCfkLHx0/Ne8t70rOM+9kd/43yNilkle9kS0Y/9aDNidBV1CjXJ
ecLZMefTAODpeEoFyWjAqgtyLZ5riTflBJt/dltjfQ0vZ9oPB/mkewITu4U4sxK4
7e6EfPq47bcQt3BQNGXMyYz1S0+USfgiCl3eFlIIRKVY8Kt258IKYPDC+/lcqDEg
eDrk5qR1uaPnjJgu1eIq2RqvLi9ZpOx+KQob5vr6/BvxSjwzwoN1nmCACUMQvliL
YMGFzg+pbITG0Qp/jgLpCMAZOOmI1fpq9MQxNDj+GERvGIoinXeANp5tGmxjzfvc
6d9ckir4DVNLfHggG8uY4ZhZ2Q1w/EwdDJdPKL5K1bs/OdROIfcOwtipUYlvlE89
9xub13FIfHBg5RfeSm/iMbeQ+fVmXTMh1VqrVII+BN6MAjGDYsXZ5AKtlfWJwUOb
t0Cs3F8tu3gPsZbvQEv51FC/iGy2QSg6eUknQ2tuIHCLvbQPjQBcVZPY5OSV+Clm
CGW3JnIONfX8aEkdWZw8ML/O67tnIgXDJE2zVIr4BIy9LdDenvYGfuHvQW2B1z1i
Ajywk3Xpz4uI+hGRIYzzVG5+2dZliht0CPg7TxnBa2Ly90t3QCdquPZqGtbd5j/a
Xx8i97wtA5juEr5TR1L6X2AiGgn4eIiVg1rzixZ9i/MqwmgPu79vBj3AYligz2EO
1STn1Qmgj0xcIPiMEl1N8A375bHQyrtCGiyXhiF09uRqmqQCz3Erz/pYbPwkfFUD
WjGEFmjMDSxIOAmou1JAjN8e31petz+LFP5s72T77d3A3rSZvY4DPMRIeKPcaB5F
FXlzzLAQSO/ud5ihVYzoRTV3wNc4zDgAXrRJN7vSUoK3k5+PGVmHmdEXogkFQRuN
IE8LVLEBXCiFmqX9ErcTm3/YnsFfbq9pxI8QOUB+GQ6Lwwqx8vs6aLNkjSPNsjbX
6i6bdQLYtj38jE18WpNZETTRgM7m7vZd5W/yZF59aF7xJzSuRjrzUw3r/dcTT6YT
X1eXK9o4SzcLyiLHMu2sNwKgGiTtCCIAaqbmDdz3mCB+sfldyIBT7fIQaXnp4KDw
258NgjqivDX/XiWYOTt96qUwAE+XgQMKGcUIyjzn5ai0xEp2EEnLVhWQrpj2BB05
maxOM7aZpFnuGjVHuRHNTRMUucSfUFYwMtMxCT0p1L1nz6qYxU3QgRkkeEN28ATf
aDIrcfJkyfNGK/EbHIBu/63ks4WTGJT0wSbAXlSZCp/QEcygTkxARFD6w93StmXX
kEqF1qc57bgqPdyGEMR36Yzal/c2lK/jv+L5fdLLmRQ0Y6Keg/ouvlD7ddZWJxK8
3ez4IIAaDFuolpRDVAO7NNxUJ2lb9By9njSAty4qziKZz+SkpJmkx7lKSsK/47At
COOZZdruMqsKh3NPFv4nHLglm5V+zFh96xOELY5Ro7h8/WzlMGtSM3wOdeDkSz3J
0MMbOSnaza9bnVcdijDcVnosrbRnhIzrxP2QP1RIjVY+f6orbwqb56/86xJ0RSnZ
L/VxFuj/BMz+fD8n5S4ULZKl8rRO61Ig0exD6Hf/Swkg6rWp4I9wlmeZCCunhpmF
PrNx/yTD/mX+6Cy+/sGJwOAqyFigVd0xcIkNVvrKKnb1/HNLikjkamsIIBHE2hDh
eJvp5Adr8mPFWUHCA+kXHsbbhB5xFyA3nUBhdoiP/vhVDwyzeO1/Zb0bniE16FoJ
UmCYwgQGr4RDWgeom2qWyIsAvoMOj/Lw3wSS3AKwOvpC57URPqwZ86GgArq5AbON
pbYyo8UQUZ0VUX8JLLesFBfGmZ9d4newxDqospk5BQ9J3UN/SH7TxQ1/F1iy7U0u
JxfreL5rRW8h2Mjtniw5M/B9kpuzEVxtfgM24c5D6jYTNC68UhExKJF5KtXYAYJf
wR4QcK8Pw732WycIR5XS+ksmlM9CegR2jvxrJKHd7Yq3zN9zkWaIvyAH3H/ptM7Y
v1cFAsCS2WV+6XncmVKKuVSZnasBxQaYN5GJv707vkfov5kt6pjWTEBI+m9+iM45
RAO/JSKbpjcj0/P6/x8Lt6hEojYijpF4FrrydNNSNNP5/adbzjp2WFMBS8mYFl7J
AKaXZrfDWyRwxdloPhPGmrBtMUVAwtekkOpjP9NKK5j/R+IbUP+VxJAdQQ9GwELx
fUYo6OAtdZ0OvacPpuAcQCusYheM6sA+zv/Ka9sMrSNlLrU99tZkSGPAIXMonNhO
NcDvWSjvm5F6MC4pwy4TqgLBcfiWcBqyaLDXyvp08GJQD66l3Jhm6HVVZxsA2NJY
cvQDvDDWqYe9zFM8CuAdZ73JeFzQTjpWjwruRmcSKCKAo8q/h8bZ3O9Tr7GFb0IT
0xy4gP5lPXJpw7RkOvOZF60QEbyiRXaFcGCCI2osSAd5a2FygXdJF/llwFndxKPQ
Jrx3YKFW5yoa/1m8S8W/PKRWGOZcjttWEcOe/bwLdwRB+zGIHpWC9Ao7YFELNstE
jSOvD+B7xHIwbH4rhho28MPqCT+3kD6mJnp4IqBmNbeX2F3jDjbIFx2RMatvJRLO
4AAAGMddgfn7KjW+sQGFIHqHu1/mOI8U1DMULDFTfw3j21Fc1E+dqkrCVsmJrsNs
PuXOIvVOh1h4+mVxdPGKuOrKyqoTODta230zJp0f6WKWrHRVB62XV/uv+FRAPwYO
/XSBTjB93QTz37q5DKA43XkVSSm8JFriJRdm4w8qJLs4VZ2fzr6JatpZ4rMICbfD
UygvopBdq5olLyBrvI9Z7sUvblaRLQQEvIxNe08VMMUoC7kxcDMQB1wMvC2oPffU
YUCpSCq1ry2V7I0EX4JBSNE6pBCxmscOnBtMvspOaPHWCcQVaRnyvsxVlQV1M/X9
hrpK8IXuaF4rHwJsNcqhKHOzWCIGT5l3jzoL9+2MyoCeV2zm8hOhFTYRXGAEnVoK
34fyTUR84qe7eU2sGFtTW8Xh9siL5IExHCYplfCmMT9TjryyekO9Z6frZJWk3uIs
jyCKIQSTSaNI1bKq17YTrsigZGir9Hrrm3cxkkvDAK56bt3uuGsdNvSmdhg/1rUj
KjqPoEhh4o14S/Vu8bAJhigvXTHB3cTmgvFAlS1Z3GL19D47fmg2VxVxcZiQF4Fl
JYnAY+ojqvFeoHkIu250vi0UNIgTwFdM62J1eQqd+WjRDl0b1qxlz9wnyRQGRsM6
tIHIpIsGF5pNoZistpKcb9HCATI3jxynMAxSN/6nWuaob++Uo0q9Mw01q1LgcXfU
uj4baOlsnr7Qe3FZT/FfCbI3TZZ2kjCgiT9fW66Mo8PCQdBNm7ct5kUh8Rx10ldw
Kat5fL/Mpccyycue+KXLRFjI5JPiB0f3sy1VS1Wj1dY5NzxXQDZx/jQ2Nio31Mu3
FonBBERAwO8DmI57+sIc3yb5EM60WuCUF371BEiejZsN3eexBGiOaMKZRmyhmwl3
ir096YYJH9oMMZR5LN1TUqWMP4a4rAu1bCLmSxfH0K6eSkGzrR3ePW5qZK/HcCaB
u0a2M0sJQo2PwkCH/8H3UuawdmYk2v/Rlog9BZt0xb4+KsF3cXUA4ZNBtjxIj7q3
/mjjL7elNUt3OoiEWjmWgKqZaWh61BWnccq/rHaAC67lX8yRhGopdi9Ybu7JEUKt
T6VKkB7M/dKHfhQROE63YaLd297gBfh0teCjD6tL5qI4P23WgsBW4IEeFXraE/z4
lg6a78RKHaVal3A5sYYbnPoYlIm+J2qisYFlIKXaRJVq6ul5bb9eYdLlx0XF/+o6
rs5MAji+epfcR7qb7YzpmGIm/6f3HBaowBvNkrkR39BS4TGj+qH24AmvM6oRNQBT
BzfMGkrbyXvVUoNeCZCsJDYKMALnKlfKejPGd53ENfSrRikr2lqoxELAVK0c8oVw
ngKDpRRZHHxwgE/8N2gSQfjMzL3nAYmJd6ULXoBF8CFNk5FPMZiEG9Pnra3h00EW
dUJawHXJd3n17SBDVwu1YIQBWP2jPHHdnbeLL3LzXMS9j/pvssrAHRM6bj41q1X3
XwkfdReBxetme8YHjXoXLHmFFEKOkP9WgegzOZZbeU2rhexxQnw09cW5gwfbIkvB
JUjQJqKg+XpczthU8LKvz3Z7ndNYk4V0zQv0WbeTtuhrNQIF2rcU+5owoNYROPOa
p/1q0G84o4QShQ0f9BZI9XPVuZk7Fi9iB52FPD7x+DTXnx3+w9g1tx2ndTJhGL6t
ribc1Oicrzq7CEkzLM2YUSU5Zr/+N+xqn5cAzLX+nU1Zmpii49g4zl8csK0+trwg
yM9wYgiQzy3kIfYRrUTiG3H4axzw6ELASWxCuajn3T4iuj83WQPmuy75S6RuUm/P
UfrdHDwKStc0/BlhGMYR3AJiMbnQxdHfES6qFJStG+Vw1B/dxqTFcVBSWH3ku5zQ
7n2n7zNwLhcgok236JeYt5WiW/L7Ehhvw5T1HhBhrs2JcP3cHLZCk27QJz6d93R6
oYTy/fI45Ic5nW6NfO+fsOJ6T08hWFNmJNtKFPweRB8RNSMoBriVd674l27j5MRU
3OLiuQmoa2Mk72a1NT8MCvnZrbfryOjtkDZHNVSUceH2bfW5KbDHIWBsD+L4mWfa
t/Nj5Li0FWqLtCyH6cWv0CrZTTjqjiva2SkNnTANz1cyOezatura39CRU/JGC1/F
+k6mlhR15VsSpXYVgwBjnt13TTKP311lzMOikanSrhVRVda8t1FYoJpPWQUY/vHO
9Ju2o3ahNwdFTNBk4CFz6EDrB3QrErtl7FvqIR7Gj3wip9AA9go9tlOG03A6iWvZ
8Bcg8Vo5D0wAHnSCmmP07rOUE9OsT8EoY+xxrADtpM10U7oXVxW/0mtUEx1iGHx9
UKQ5DsHEGl/S9IDr80rX80PqLrOqBFMsIokCIYM0tDheHS0JZkWaIgmJTLo7jnFC
1MZM8ZIh0MZvLAnoZD4O67XF54rDKjF4l+kNQVi/4YO6MBMlOWHOrl4FO2/CfYhF
hQe74weZmFFh2Z9GRtC+qFZGQEv1MHe8DUIFU5osxDClSJg1/GOBYhIij+RX03Jf
LxH9fjsG/RRxYSsVSWU77CsWMsuZtH+5wWxYxXIRyi7/seBmoZ3pHfXkh/zgJCuZ
u3nqaZoOTGp4FgG69ZiUs4iAtvwVLd2uY7uY3SHJdEbqF1GssWQcQf672kVuEKnD
fhRmqgwNBdN7Q9mcaJV7Oxp+AzrQd/qhoPtzikPjwsTGkcur+e2zavM08bR5KhbW
AtVNR4TxLNsnaJYTkOvV0XC/tpA8V2wjG8MxVfpV6FNYFhJCnXZ94e6QVRz7OHIa
/ydce0/HQ4p6o6438v+isDP9qvs8emhkZXoc7m0MDcfxCz3LKh2S4RjGp9ZbqWQF
/1bJjb1JJBIDINDtQKcOGibouAoxM6Qf35eyGvlq2DP1fyPwgHVe/SRmkYHdjZTb
JfQ51KGI2wYXKjVSFOra3CMgTrMF+W0k+qf1CZp0ZJf5y2ydRS+/hts1MJBuyzUV
jxMIO06x4Na7iYLUo236C6e839gMmHrTYsy6rHfGRbAUkVignUpLtkkDCbF+LDEQ
YpKzmllJCxmHxHTAI4EaSjvI7TmK2nS+HAwKQn2PjIKZGjLmuvZDgwbda34E3mbw
SkSt1XqlMc1WwRrhJuI6kIhoReQFUH8AL8ugMSprQPQViHrxXQzh57TJSydMNavn
i+uGu+eGBxyzb1Xe5fgQrG3KqcY0mN+2fMRleCZQmlqrbDdtsKUhit7n12sLAzEh
OI8KE3qJqZ6Z5NuI82Mv99RvOaBpStkvtQ9ANIbflRqr0iz+XX4X3NzAlzSwB+pC
MLzdvQdI000x2zj/gjm/bGQlKyCTF3FO+ieQ9X6i/2JBUK9DjJG1tn53Dkr/YNSF
stFYX6iGID+TpEmdPyriTm82xC6y3j8i5D6E9OpHUNVoHYj/1rZIkmIDJpAjCcms
NKfrPx1Y0yzyqKaZkk9t5e4H0V48b3tZhmQVoxfJpEjazlHnYE6BJOpKIZtPEDLB
DGz0yINr6qpQ7URxersHVdoW+aagjMGNcbMUDVOCvXfu161jTURKNIO61dhYp/+j
gxJ67M4BnisQ32Sjf/FdpXhsmpB2exASjYVem7pMLdPewO4QiTlqR++qk91DIZ9q
jFtGvrJe8faJV5gL80Qk23o2PqDrak/4R54sYUVZiignKc7dvF66ZVTmoITMMfQY
iNcw9lXd5Z0ByzGHH6Q4o2EG1w2JbTxD57wQPDZDtH471qTc/2flpbKVyI6AI3js
N6eus6A3TDhHLCTA63DvPFkMB+iHvIZjsrfbnhvTF5jx+MIubZCagCmsJhfJC9nZ
d/VFl3i7A76xaolvkHMpUD1slzah6IBxpbvQJLkeulD8wJtOj2AF+BGJaDJEvhQa
eotz1TOygvA+yYeCNjEcIa5Rm42SqEnUfNQ9sh4IagpkQvdNcBN+Uai1klfUUiZp
LPbjw5/6XiRy1W7ghVZEky8MRSANrhjjaFIpFs32gw1EMOv8zVpv9we9yDQsHnrz
+k+SBakk5GI1zxqUBTzm5p/1U3HC2xauQQ2K1JA3qvInVZsgei2bF8t42zqq6LXu
eOd/TErivzgiSuWJejeEDtlJnlO9y9QxsZZv7joQsM7UYQN7IsR4C8o6KE3Sas+n
HIx+7NiQ3R9bDF193hYkfY4AUVlAC7jLHAZHT0Kvue+9zERLlg6FrsraaVTtofVc
RutR2CKM8fqn6RmLlQVIishJXPasADWJiQ1LIkT27w+NxT+BsDtexbbZMbf2sFc7
ja/YJ7eqXgnb4wKBZ9ZApBxbs80xdlkeEAzYE+5IrNzZhLarTsIszFYsakMHLTWz
+1Vb4Ib4W0KjpHa3uehXH8Jw4+TfWt67BbykULnhb9abOeMCg9VSkAhs4Rp5cwUm
lhu3kbFFHgZQ8PM5Wizy25BS/oLE3mlkq29RZkgbmceSAt4DV3uja3/DfsIAqw6p
GjzTH6kLhP+Kl9xnwIrj0ClOG4H3Me7wRM1Td3lshqSg/+sw/oZ9/6wV8sIzbQy6
WPnskvWjFyV14j7zsr1O9sO2nTBsBBeHVuJztmQHyXKXKJawImDiQ0rYn6fQ9fxE
7CD1yI7CTI5hxOMY9CoRw9u7mDKigSS34Q5VzOfpY9hC/8IVKNM4T5Z+MXoqfn47
024fQ/Hb5yVqxPJsfPtGjsb4ENSSHtTTMgOQdG5OCOErm5EN/ieWMVcQ5r76mjgm
pX9RZQ+tzKWevzMBogl7x5KLprSU91JaVyYyFqkMxVq7GPvD8Cp23ChETBLP/Svp
pCX2190IhVRjLkz612nH5vj4DVArjIcXhM4xal5dPbasa6hvtHKCH/GoVedZbRo+
Xh71e43BeZC2PZSXgcUwsI+x2UWDU/9wI6clLiyMo9isd/v7NCQZSlXErzWrXoPt
RFNO9MickhENM+sPoAv53fQda5De7DDfqi1WHAfcC8noBfDZ/tS3HriBsipbCFHO
3LcEU1GSY0OF3oHCcehc7HjnTCIgBrGGdEYaEvvNvaG1BW/QcbQpC2HRzTnFDkEM
+jqnkSfOLXNPRS9Y+cT349DMzk7cgSeD2NwuBwbs8R7y+eXIhG9P9C2eyPHv7/Bv
eWvej2vm83hRr3/mSmbxMHOBnQ3DnVJTRiYXl36s51nSIllfEzfKTN5S+p2c0R88
qC1HZ3bWf7n1lviwIYX/3OhJZ6mW383ieiIDlZCLVDMJUFNOLjcCAqLTnIu3JhPk
3o7cLaMiqStrVQp6qYcSMm7Kch3mOn67yiQc1SEFIbISTBXrIqfCva/Lx0py3Tip
XMXtfnjnuWhaPkiZp4zISL2Hzko+Q5dAQzTnGapJrQd13U7tHVSIT+1BwN+Xn74h
JZy9jlsyH3FmnwQDepzdnL5mNvaqd901ChS8UG0NRufwoV7jHp7dp8Xv6xDFntvv
/abfkx8tHmi27BjKSjzxjOsYhaEw7Cg/Kwb1fpc4nHj81+UM6ckyfrSg87JjNMEQ
cE9R0BfRq8xEY4JmzZCRKN2gO17kHNl72jhhx1j9HUxmOB9k71mA1GCK02ITApfL
F6UZoQjK8mXy45Af5/bNQdOPJMxCOcFT1dCUx6mGGSU4aKWeJDZPhEveUQYu2prE
Ng7rJfpFa9RTXAovHgr9R/eYvfcpoD+Nnyq0KamRVZKwBxzRgySUbCqtQmahISY7
6XUtQwXCsLZKyrAhAIew/3Ro9Ua/mTIZfTMGqF5qZIvEtxuICgFAhYOauS4o8cu9
uY2JBF6rD/8R1yD7rJFDvQNDX/zloFcS7J/AT2HmnFugKtnw3eId+DNMxOz1B5GA
7iqOi+gUrBNMYTlOJQJ3ZUdhPl+INVQ6jOvNf0dB5MCAxawyRuVsorKhXv2hnyhY
+hbZNKHDTIJpalvgjFnSHWMYI3513biJr98QQ/jmzeEbTVvqTUBOL7QEoq1cr4i1
jZmmZrOqE3g4NahdsATcH6Tm3JbDlc4nefb0NKmq+aw+afEUWWCpkev6LanGkgO6
jiSHR39/ElfFDw2YM3GQaCpJe1rGMSslWtGPPwoDF3hZ5aGzpmmdD42pynysc7Ge
P4mejgtO5Xb7n5jLcum1QbIL1TorYKzOeiTCSuXiJhrpE+87EFzzE4r5gMQkunAs
Wi5AObE9i53UXJe6KX9vPjnc8BlWe0lY+MCLWBSiKkB1m8cqtWSxBik2yALxAyBX
7Ar3Z44A5BMhFL6IgR3qa/RVyRPSee2krmhmyShteZRRgRwhgtcwzNJyH0ZiZHxg
MnvmP+j3obJFnyaWfO/UL3dIuaSXAYrVNRlgVWkyT+HLCGmR+jgWesU59ErsSLy7
+ArbEBKP40IM4RSXvLzuWffT7s8mtBKs1MlcJHgN73sJA0IxQhGRCDJ7bvk4yWFK
Vgqc1T5rRXcBeUJuXTeXgv6kLpKjS0Z4+zW6WQA7/yNtqXsvmKScvGCxYU59SOnx
5Yq/JShJ0fe8z0TER6jGPaFoL2pxxEd9A0W9ExfyFK/VsH/WNHq5DvkzcFuHXybL
8ddXqQtfgQfwnvQQgGwV/amZICtJDqpxVhR/Sfc7h+IGIs9VJ7jZ67W0A1dIJbU/
LjlRwHg2VTTpNlh2lWeffa5r+9uMPGUTBt3PsTSnIuT9BztgEo8HQpwruvF4pPPa
CJ7Wk2xqNRzAazwtAtloVEPzwnM32RTYrG1F47wyp/oEa5gLBVFDvCue1sBwtsOj
+DgJSwBqHV8Ti0BJ7uewp+7nrqtHWKFC4n6IOTzkdI7Xap5rGZahCo4yQnIdpA43
PNwjMzm/X6If57IBFJ0auH83SfrgOfXRvvozbZmMxkNKhvdHGWypmIoBRlzv33l9
Kz/z/F7MXyH49wtpMVuOEqMuwsvbmSvFMY+Jz8emM1ex5JIZmjZ9kUS+IWpiKVvn
4RpQMX4ScWc6UD8gx2OsGmljp8uazjFh+do8/fmpRvEGNQceys/lxmJHFJVzhzTz
mZa/Pzm+J6CsaeKL9skwfRhBrftdHkSZY8v9s6aEtN4PxfUiJbUs7rIc7dOAvf2W
YgiCF/5W1oAcrb9lgESRp/crn3TIc4y/Yv+FOGs+jPgm6DwIZpdL7I6TFEbeiWPR
+RPmxybG4ULL8QQQ6XIll5oN3ZlS7hegmifp96vSelYWjtbAmOapA50WEscwuUcI
+Y+U3u0/W7390X5LF7ZVRH4D+Aqy3Bsj07B6Z8A5xoOf4E5QlvuKr5N3lHzj99ZH
zAHtUQ2bprSAchAMm9IuIfm+Nx4NgiccMeC8Iy8h63+nJo/0wx33vbEvEm47Y9tF
aJrCmyckjwcQ6ThuoCWT7tTAjKQQjbAaeZBfqm4eAnT6pCYj8wAx/uioFF5p9G2X
BkBb+T4NR1oQfPpJISj0+OGvn8OE7ZHuiIcDYhaNqNrnVJCPZWOk3nlQt225WAE6
jNNtukKcaC1d0jH3mu78qQElEpRbqdMqJN1w4taTSrigesfdKs5ZDIk+4Kvg7jcY
+ZgWZJlwznVR+VX+smCzBiB6iiXiqPifi0R+5I99YvTehojeGZx4katUJdbSEqHO
VQf5gYKF0Ezum89jtH1MQuuHNLX5vlHgG/xLmsX5LU4+h2qvidprS0/Whsc1XUjz
7vV98tU0j7Z+w3grSKmFj1JQd1pIUbifMQGu6ha4OOX1kn/rwSNUnGLTzgDvbFw/
fCNkRtJ32VbPavDb3Y7Y4rsNice7Xwp6JOQShDi8B8n04Qw/FisCCd+JlwUU8HpY
8FtvJt0LrGqtuyUH0kMvLge51tBgd/dXhKmM8FaeErrtjmcvK/HFYPSMyOpA2Oo5
cDaLZGz08dZhlvrj6x0iVPs99hR5xPZH44HQBONXWpiSWIgfeVoLFvGwLnCMxZws
Ppi41S+6kcxRtKNtcc8j6ydQoYaVIVpJ4dLsVbF5vq8mYUO02BcdfCTWGCtdKxVT
rAEMLGo1TLxs5aLHrNjHPB7sPVk3ZFkzqzsqXW46FLNuVhb1OmJiNM1A6kvZV55F
eoxlCEuk6/tPGKs+o/LGZvm4LSWuLCTng8iJPgQU1yBvbRI0W9leSU5ab/7aJlTT
OCFNe3UkOt11BGXwCUscYQyTZkJYgauSMgoJlGry8uAx88eOaK4fiD/Pm9sZ54ME
GYHoHYPjYAvEzPGL9fINqocDiWWpBU0P0pmvlcCa/PB2lZe1RfqPbdIwZLj2sdeu
ETMLQlPpj4vFzgzh2zO0mBorZWrBP6Erv5LvjUysZxbBLRMQub5sM1WolWekKfUW
Z1YXfg79sFEenXEK+idfYJ7JLZU+9XStqexTB39SV7svrjGmndIwVek7ZLxQM+6e
fbVC37wYyCvZKEwf1kwrqVa/nXkGKMRUI/biuUyMc8vQziYRvC7bo1vgoAewon+S
JlhI2RipWI8RbOTk5qzXBUAcKuETRQrS1H01UyV2Eax7pp/azoacoDWXjzklpwNi
4NAr1opSA+lkp6I71EHAZggtG0CqQzSUaC4MxOhJ7By1e6wdoFOtpj0wuzcJdWgc
nnUAsKoORxot3v+fpd8jR1lNMvXHkYe+Lm8sgGBSk2OcaWtucGuM6X//ZPcR7RK2
OTH0YhmHLiiXdnyfAeU3L0LkCCLomQxzHi2rTugDnss1z9415pw+kd7FUrX3Tqyv
eaOgk1ixf9K6tW/ZARrosDIu1MvHPzlZ1BdNmrbKNa/4HBIwQwHHvYz4ThLhrfMR
I0rFdGKHrrbG47w0Lv2Xgn16hkVruLkOxIBaC49HmViwuOdb5JRm/FnbxfUyc/Vo
dvQf8Ei6bMUJn0kaYr8ergCAFibmgSruVNU0viSmp6papNIRGZfO1h1NNhjx3gWS
KOPKJ+ME4lQybM5LPOOgq4r6tSGTiMMdlx+foXCNUzZKPzKRXcQSWDlAjLtFyD0l
enfCvPFphc9F0pdXUWxsvBr484wcZbRb7+4OnqlJJLDQTv28yDnO2/SvxevcJzsX
4I6WBkQIS6CRQLiEqT7ou0ATDNbMtSPxErq7jnjeQuQFFDvIjH2k1z0OdDTQrxD+
nk3YeUSZvaO5KDFjs5BFbZEkZyFiSP/Hgx42Czg3Afkgm94bwl+dDl/DXBCXhu5c
djiCYepDMwdkRKbONkWn6XWhSyTn3MfL6Lxpeqbfs9ICeEKrX2PNCZT3oUkEAe5O
eY+N1hY27T5hiRIK1JBmiksgA7CYUMHwi1rNi2K6w3e7TSoS1tEhNv7zDH0UIJ5e
LPZCgJZXBacMYnFgfLnJd0YOE74Y8YIp4FNQ9pE6NEl6AUA9O+iBqTeL3v/6cvjv
bV0Eeo2SQ0HNakjuwcX4i+BQviMs4PjD8Q0dAA/IGVHQPqfztKXaiVpD9VWU20p7
Y4V6sqljXo5w2rTn04yHGNfVILxHowPm7txvUYFmanIevnkFVl0tCNWvL1z7bOAt
6cAgE7L4Lr1QGJ8IGN2fx+oOktYSMxC5lLfh5PXizSkXPh7yb7+XDYGjR8LFMtYA
CORkXlx28pzmP5yhlxWmhaWmvQ6+EPAMZwpObL++5ZrRLxfNuzgDg3jEQf2cF/GP
CEJeZ6H3vJCq2+u6XjMXLldtpeQ/i9JL9dTreF3Z0zPF5TrK2UTGmGuVIQsixQvs
rH0s+OgYVXJmc8QsxTkwaBb3n8U4SGu8PWcAZcvamCcV6EDFThQaMGpMQGmChgk+
ROXHVea9MGBu66ihGvbn//uZhSMW0rj1UFIkpotgK1OCNCJ5c+yPb0q3AcvY5uJq
qRsiFLUv6GKfSmCGgrYH+U3CNcLOc1w6SlLGcDdnTwMmK96IUsSiqK21BYfBkpLY
ebEEx2XkFxGDbp57toovHTCwm1Cin8jWUW5CRZhxKxpG4eb7hAO0LroT1Gy4tA2u
Y2HGCM2lfoS24xlx8/C0ToBEAkMkh99Gdv1PjQEaDXS6HUYrC0dN058GEU/nq7G1
4hpY+XkkDoTvI+4RhEcaBL7HQ2YDzhlPjlfCf6nQEFDcAzeF1v/QY9Kmz6aGdbIz
2IdMhBf7bGlietphFJ58AaKFgt3RJOJ32Ngd7wHF0GJRxTqCGRsdOVw9d7JmgJyn
wAbp1D4uLAGnMdE4a1bbO4Q5FKf31x5XC1OdzxtYP3qAYbX1BiSsOnaJacBSaOl9
4ZoKoUwORYDKuc7rJZxX1n8yTtS7nyPcFI5vayN0V/x2dVM9UsSrCJ/5ZYPa7juJ
9RBOFb/wYykBki9ga5sl9txxEd5dTIZ0FzXnR7pi4hd+mwF7eTgQUZ9Rv15L+U9A
VtMco+UZy4xiAXOUS+T3hSzWNdo95THCyR7tV8DpOdQf8hiR07SK0OoXUCYqb8cb
RwpU/IBHHNrMYuRhfmyUZJbiZRCxQktF5A2a3UUjfqOx2CPWn/lEGR9bopB7pqmg
HnWRxSxxoJA9lgDFl276SDHctgLHJWoLz9aAZRnTYjX9SK7gPmK4sUwHiMkoRn8x
YtBuKdt6pcGEbmnglHbtk+Zk0pG8TdlidhzE8hdKiy7fQPtOVRPf9XW5G/BhZz43
wqZ5yCsfyoiYd5bz+/NsFY83UBtTQL8eRYkrza2WjxhDIx2k1wUiJ01uFQwwgGOm
lyghHUWYnWEUd9QkXiA7sg8gEuPYkK+GKQEBezlPZ0xZuszoUcL9D/r1SzMO95k5
tVish7o6votjka9FVgvzIwJFMSFsvXc9JJNO6e/je5wlihYzj0H6ziUKrdAmWc2/
KKSAWtaXB55XG99ngalD7j6L196KbCkzop8UcE2qeIfDXM0eOqosd2LczUt5WTss
LCRrFu6/YMQboXIf4aX64gAYJT7Ls1JCIX3Lt1yOYA8fB+YLttcT6/CVyY8jAAhj
Tu9HXzSNyEfKetJYIfmAFd5KapQd9rW1aOFv/cWDwZ4CtAlphZ/bN0W4bJ3pmooz
iKjjPUhfyh/nkSDnWh3gXfaXJ+HWywbmeb+VAoUMuoSRQgxAwzxIRWoGqMmNxpI2
siIdrqSl0Zz7qQehPJrBt26JCqRrvIca1Vw8cuFoi5s583wn2UUTBArPhDZtkrKz
CpghJRNN5Qvgnre+xxUrqSS6HxjK2k1kDS3ektbuTVDU5LwjuLTr9zVlv7nR6hpw
i+4ND+0d/7H8oNdkNpGZ3Qo7vJe8cgr/po2KMqN1w+q/oX0txCFwH1iTUaKxmsjA
NcMK+6sr+9ChfGJEyJ6GPilZF0ll9Nhpn6QB7qTdGoh+Cs3OUBBVL2EvDkxX7Ps3
EoTWiysU7RzHSa+1m9cI8cz+dFiqot5H6ZkKlM/PlTvMP1zGbmVRVPKHyXt/aSnz
HUqczLyo2W1B60gpbD4PcKDmsibxojZJmMI4DUc64gWFQIWJAQ7YWlLOmpjZwiXN
/BcsT5G0hFw3/E80rEVa8h2xvcx/C5RlJyOmQP8iRz3qKSUNTLPlRMmdaommEZrX
Izpdc6YXd+zC7uzEqFsxKz+JWgJ63kSkOLIHhNuz6OXWhdwKmR31U2fSFmnZgoQl
1bS7C8bCs3N2vy6dvUQNZ9itY2dRtZRZKk/F6Z2kTxIRSpj3ieXM985lfMagQKRe
G6jhuUYD5Ap1YHdIkXeAt5zgiASMqv88MUvdMcv1Pv1uF85tQmlmeloFbcRs4HGY
YuDDJwTLsim7hqKMvr4KGrh9S1quWSk6sSV4DITfDdJTOLAPQ3ihIOz1ikCVTd0O
oos7oPZNd5Z0hWi1bc6f/q9NopPWgGafget1PNnsDnJW4CLqtsMUiNKtgXE4Duwf
9V9yHHqv/lqzU/QqtqAZkyKWceIz2D8dp1QoJbYj0STy0MXg4SsP/1OHvGvwT7VU
fww02mFm/Tm3QzGOjkcnriFtgtq1lovVgGLaOi40pDLAv2c+MyBUgxFE7f3X04pY
l8JJioy2rxy1o6eUW10pf0+QY5GoMTvvlNprU+qtOOKqqC8mU/wWtmV+0ZdDjxeX
rRO619BhelPN2Lgb6Z6FtS2zkt53vcgxf3nOc/N6V7dsUmaiLKxZ9Vb18Oi0/1M5
XWkL0KF+Uu1IJHA4HCVytS1sdhKgTdOKT6fofnvlxspDLsEUu7g7K2s+OetuWN8u
uNJIbEOZWDndtGWEwPXtX1bjXBOuBBrR3StdHIt2tkEvtlvZ5gFaFAAG2G29qYHf
7RogXp0+R9Uhp/uCbubEDttkzUpXoVcAlalOcNW3NepjHiaT0BaNliImFSta6FGH
Jdb8FgXi8DJLLV/Txw92WBvmEt1GWwR/RZrudbkW8LRKpFy4bVgLDCoePmupuHjh
kke24D7vYWX1uQnvrDQ/VFb6mFAGBh3ot8CqsOwzAWQapCWKb2UXRGmuXlclqRHK
3TnAR/VnWq8zjH62ZhVicIkxXgPltBS9G9hmF1B6wdZDfUfgoLNovvPmilW8ZbFd
uKz4YKfxC+c3967RLbXoSa2abH9Gv3tsyGAm6puc2lFAxxCJH4qyq/MSZjhIB6X2
j1uDo283c4Fk6A5P0gjtoKtAT5ob3kjrc7e06IHhrUE/ZmvnFvTrRZ0kKlUgRWv+
fqSpFRE2OlhbiEN6muFdYAtrdnXQJT4cRgpkl9wbSaRDQ0ZibqXnLjb6qa2OX/5C
5wxe+pF3EX9sZRpFe+ggAVMdq2264398bkRgtpRnNQRDtJKJ2Qfgw7p+m7snM/xJ
o//8t/drR6rBHkdz9td3SIvHj7IDRpQ+r7tURxjw2vXW+piNVFO/JfX0hnEQoHDX
Duj1qysbYlgVccH1T+1VNm4Pt4cmmSgcGl1xCpLJ08AcsE4ZnIJItYeI54IXS758
XMqrPehcfpX95YVVtFD39mXpvgufbi1x8aTQ40QhmUiNegCEZmWw2a8bdWhdnzn6
D1gq6aw/dRo8mqyNxDgyQf2IeCaxyOcig/91lQelgxGqurxjAGaMb/Yj1K5Nr6uI
r1YhfFbCN8JN6Ql+Q+NnTjnwNFOK4q8AXd3+LNXac6LEvHPmGHYLggAnPgKkchk/
pqHiaF9KtdAa/+ZClkBUHhLiDmyAibZAt4ufe09F/jG28D5K9Q3LH1dkhjHVtrpE
/qsNsw7dyztLcScTHuO4JMF8Ao35Mt4JmmesOLHjHGtWbOLcZ26e5bvHp2aZUI0M
WclkEEhYywHw6MW9HEIBZvscnj1k6BObMZfzxtzxA/bbIvs2ky0JdtTrThoZSzVA
BFFquBGNXnkpdPLxhh74iBl1bEPC2eWA4fl+VN9Yw3ucpheFeeHyBLjJJRtMOYii
exZ053OyKum5y5mkEXzD6xhsxCtuRDzdzZStgOK+kr5B8Cur9nVTYBXpyZtDLTSy
Xg9Dc7qtWjpllK28p0B8Xx53AX3k+j9uw87GUTvFV+PqioGaio+3JT1VrzF+XVg+
wt3dpGFTNSmem5NVHkCbnID+eRR2kw6jMsCn+L5kD3IjrlCkhRJjPjtuwaJDL8Pl
wkGMtu8QKGBQj/1lxZLZQjSsOMIU4ms5jeAsJtigcwzo1eG2YpXqXLNqSKicEIaJ
6959yPGmM1pPh9k0ZcMao88GOSLgs0BwDmQ1TuYl1xsdFQSwHi4n5OGNCvQwjp2d
oJ/SpiuvYnSnMGP6XcWAWPpV+Ziv1XS4EWqArfDVNPXzXrUD1WsAfATEpcz3cUhV
a+dir55FBf0ERnZKFypLXGXNSieAmsO60afMGhuzeMZd915BDItPEGDPUlw8I8ro
6hCodV1g3MT8hpoWsxzKQtFk0ljkvXgkL777SAI/FnvuxRovR6bSP5hIjfsTjo2C
or8U/1jZVQ97yQuedRli81jIbwis4p0O7E5WDonK8mDVn/NPQMrVU8TrlKZxGB1J
NSwWGwWjKFLqnOiNAEou0L53XNeSRxyj5Uz5zKwIM+3AHWQBgVNGkrw+AFxzuKdM
o81Pyh01ELsdKvntsOHcfEmV5f3a+uY7Sk5lh9/hdQXcA4tgTf8vgWcKJuOhThoF
yEH3HBA3Dp3cZ1MH2a6imhm0Iyu8T0ydCxJU4sZlzygbsKEfkpdB3uwhS9swL/RZ
/eqe5FskfsxQsGYEBl+hvedhRO10hB051seTATsUuaDYhoqPPbbZETshT3Y0L1RW
es6v6yLkTakezdlIRfBzGDXEXA5hY7iDdnPALHzJPgqtrGGWCkvA1c2dyED/PNY7
a/ptJuLxnhrr+U2dWOx9i5bL2dvtp7EB6OZHfmjxwQXmo69T/DmpfLI7riV/Ge/8
Xe2jkBDbMUHJxtoi1INvb5i9OGvnYlj1tXTyzIgivbQwZLdpGaoevihMqOKcSAZN
i7M87XLDIElOZ1svJ7/5cvupdKPqWz+7lum8fm0tjLMEO1bc0JL/lwSjiqbui4wH
fRXexSsBWCaQxZanyVuXika1uDCZrxydJunBesbvEXu4dhBFu5BpFQ7crdtdBbNK
lC2XZG2eGFDlWxne+viPBzNd0/o5HGuAzi8IdznSlHS5Cv3N4P9uVBC0Mqz9U0Fq
iSFBeXaCEEpSqdkh8r8VvkHH3E6bcClZ35G0TCvAttc9Kx8rX5kraeWGkedaI4j4
xC9MqJwh9YLpWJQZxTxdJB1n36bTpH+AlCnEx3OvJ1esQuE/YiC6hUbTtIuxc1Dn
HfxzF2cyMhQyclsxPPQYozPkw846eQgI6HOPI3Yf3XIyrPHMwpw/0cfJExFXn/Rx
w03X+zLlkZnzPrp9ermgoBVGeAYFA8ucuAFVzNR6H366/q/0sbcjbjsaG7G9xUFa
8hBVfo1+zpqWMkWzZ7+WnG3jFTe/Fk5Zk7xUtXcchiUONXojxZlCaFitd8AwJYZF
XxhekDqCnHtWj6PWc7xA+yMV8pXO9RfWR7GQ436sZcok5/GNev06aUx4lOmieWdG
iPkBx52VEaRbeea92fIgcwiDQP5FOvbotr7Ho5EYT9T9UxoFFDiwgPYQ/hbo8lB/
s53eCpLTqDlE7ntyjTJpICY7e+sT/wQ+1rmr9BxUvcbNOGwWGTLKCIaabNwErtQs
85Y6FSMRSYZt0KC1pY1SGqVGeoyDslD9nnniqTCRyn6P9FQRLNdxq4ecqDXk3zYG
eTQZ6eXt76mPvtoH+iPndQruGAy7uExYNw6VkKehmstHDYEKljg4sX2c5K+OLIIV
2/bp3VSDvrghd6DvtEZ75/9o54c2htOuQK7AJK4kaqrbNpiIlZOidk7R2baoB1i6
cX2OP4PIIxERHpYz4zof6+FBL9YkIit2StaHxQ3giZQaC/PV83z0ZhYq/wT9qhHt
G6EFAIyRAItuX5GL4Cg9SBwdXC7JPkAzPNK3I+JZDYZESRDK0Xqj2UGJLNt7pgVu
Gnq3qZxyU9le3m7/OGWpDjtn2oYjY9F2d2AUQuBiDexze58lyN+XpSgkOe46DGMn
NhgAWbE/Ao5701amCiFjdiUsPYfzioSQaI/OCuMtw3+csDgrDmniw6SS+45yxCJc
rUUNHwA4tLoBcPhI7Iw/I8VHPf9CNdhyLg9pZgautDqWttfqvGvDelJo8dPxW386
JJ7OimAlH95j7E0UyouXVysbaLn85ASG9pxlWaoPiblPV83Zqd4A+PwWLcAwGYiF
o5fcA/HWDmJRgxTR6aBv63XLA1IZU4w82Y4w0jX3X7fY6Uky8pG6VuL5e1JSB8DO
zS6PiuCwSeBEnxBRD/2TS69tDsyu7bfwCfIdiw6RhJm8QRI3UTwZ2Fy5sdoeQEwv
fZgdHhDMA7ejs9gQ6FCbc6AaJN6Pp2rbBF8jXGpV23FRQ4J4nzWpcTj0uKwSi1m5
4RowSOUQ+n+QT0zyBMlcLyGEDinG0RuFaGTZkGegQdiWFdiBHtQJV0E0THBJb0p8
2zFHZ81cxBdStTercP2KyK0K27l9Gi2ZReYvw9zP5I5QuJ6w0I9f3hLLwJtMI1fj
eJpY9vSVgspJerYYexzUMQtmZL6K4tih44R9d7uMOhB3F20MpUThwh95iRE3xAzh
NuK71IcYqn7VNG1G918sXp8q64Np3hvYfitq9JiaK/rl6iIEmvir3g0v+bf05qS6
yH8rEg2pX0SrRiUS4KZdMldTjKVX5+xQp+a43DFN6H2zEdxoQ6koesQFffbm5t/A
VboV3LsW9KrtVUQkSKY1j8QIhGRg9CfMuKAMlObmPStMbhWGav3wmG6L5NIZXD9Z
KwqpeBmSVdnpamw9zxh2fDjZTr8uD5ZDz+P8F62TwrkrmIq9bERbfs/R2bhMRKYE
f+pebWWUJgikS47dfNUrtAJ3t4A7yi49OKCMjY2DM8Gt3rvIUWQ7zaw1kmMqGOWu
KXzV3QN48mQ9o7/2g3M3BwjpmKBYkMRb/M6VSOqi2NLU/O3/mfXbPD4mQ+xrwLJK
cryptz9+zBAQRRq77Xl82UMxyM6FuaWUDUCN5JiWTnAdCGEk575or+NTSpBx3BSr
wAfUEugwc1v+J2IlKZjPBc4TmkDrnVo+TQ3bCr91OUjy8Vk2c2k/6kt2qwhOr5E4
2DmDe+K8DisEmS6Jf/YIPVWghV3KLR+aeSMdCu49U0m5q0wiuK/ZXAPBL4pYVAuq
YgqeVm7CjxKdbM0i/g7dXvJTxF/91MMXor2WybNdz6BD2UWyMoRT0J7gPCxG2a7E
7QJNRABEvar+It/CSYzNd0p0yeyYSjh29xTx8pbEJ2POQ9KUwtuH641jwlZJuXY2
X2AUs+y1EyVxHaKZ/oU62cY+VRvxM1L7qZerppDKPwr/rkjPPYpmilb2J4ekKrQu
tm65KSkNFS8Vlmy6Tdo4qkOjneqhKsE/jb48EPjfr6tIqn049PBkiCEUDu+VShR/
pWum9/J0ui1NprQtulxLPubI06ImSoGCH2qB9XhN5Jjr6uPZw0j0XVDr4tHFF+pC
DN39ySU9H6uNvPAnzKwxtJkhDfql9P7UxpGJg0VVqJXJBfLMyUsbi6rqk2clBhYp
8035JZq/n60OJTXSbdcnvYITD18BSSyvhfbapVJf8u8mm2hhGGBFfgdzDSudEp3p
F9qvVw3CodMUhzSRHiKZUebflMWQ85QzIMYbuWBPdr5SWXu+Kv5wtvJMUbRONYua
hHPsHeWb1IPYb9hYTf5CX48Vxf8PpWeGuyAFdVrAJCWYr3T2dF3kED/zLE51VXLk
aPAmL8al3p1LVbHuvU8VZMQKgt9+GQGWAA0AYLAQ7z2WE0AdcZSRcQkYSfqxyUCa
GXxSH27mgio0VxYU+WRYppfficvyJOzUBaXArG34v1xRGmzKSYdvyR3c59aR+HKj
rYsAu4ZXJ6Wm60aAp8w4I4M5bwwrztE1z/jO+LOJ2wIsGKLeyiRyWqiFVgsvvmDv
LxMTbjZWt/182Ew5ynM5U1hfvGtjvyppO8HWiOmWBt330rYxlPcUj8ritrHdPwya
CZQHIH8gyRuEeHqvEmHoqTzWmB7H3unB7IEVHzD0udG3IMobguff+/tyXMwfduzZ
S16qu75/eqNWZLXoUeY7eMgV+KJQtd/nNTf49DhgTPrHdmX9pYrdigCA41e9qa0d
gG9PDgyjju3jwz4baYc1pKAVd55UX63x6K2/a5230kfvldLDDnWPhJdeqsLgQamz
E+BNgQ9+dxE6T5PHcGhXQWMef+0qoz0kg3P+6Wu+/FTiIfdjQGnOkgRbtlN3c9e/
2mzKOxm8q/oHIwI7B1QsgkkrkvKLViYvd987BhG4FDlEWEBlvrBMricolPNf/ri/
jP/NQXlNsg8rdOtPSMCCQJ9UxyKIww1Ng+kQeLwqX9LL88bkseQAEhX2PYgxScRU
vVc5F78GfLC972hmp/2WjkHF4+pzbdaZd3KMFU+Jp88zzi2p+5p3/5DQfq6atRtA
TE/bo7kvB1pj8Yc7aBocdfy5JWL9hABI0OLFlTm0WwVHwy9jSdBHtbia0Zow51C8
d2/o1bEwoTzG9A2AcjTKJUrQO6MyRCvRCK3WfQeTzhwXBcE8ueiYOX1bE8LtJxL4
rdtHU24MqWjOPffc3SdE97cNwKUVvmjEOfKzH2uOb1r+P8JwEus1xor/KMr5hEPn
IkgBhjeYmM17QAZRUkPnxlZedVhdTj+N6OV0x7QsdwosZr+xAnPRsBgoxLH2PZ2D
17MLrff4qfUxT7RtQWrzekLIQXetPunm+ENp/T6P9oBkTNZXwM0s1POXGRN3MdE7
hSSqtTB8+QqmSYaoaNHTYeQcvcJ04KlhrHyAvUT7KOMASQTX+ubErJvkh4W/Zqc4
gE169V2d7ul+yYFHz2gPlMAmIKJzEFTiNVuYEUnfECbSvOn7nohgR5nFMnyKwYC0
6EzbAjlbUnrU0+UGaMkSMXTzYza2XJPqdx+sRX42Y9uP9ejpk2npPW2qemkNuOHq
c3cb5q0PLsbJ4sSDkI8+tfsiFoPjbuqXA9wq+WdQPJww7ZeRa/EpGfpl8tAOHe0z
f2rwGrULue/+tfFoVc7HkN/Wq5f6/vxKb7he+ZQtmHqpVZ1/F8oLJAMnImyG9R03
UyWC17cXEQ1fOKJL6roaGqqmHZoeNAOL/wAyjMpQShsUP0WPJgE2ZhmEgnU+5U80
eGEnIoZfh8nFrqSdnkbAEoa1o1udpHQWrZ5gp5F/FRwDroMVmZcDlmaMf0ahfwix
aa/mKW68R49B2pIwu+G6x30T828H7FcxJuXR/ERtQs1vFJdyJpr2NQKS/82EWVZ6
+vxQO8cHrXFdGyamT/tpxxNNZ+O+BA490aflWAPAXCr5ekrtQHI0gC8NRo0OAyO8
Ki2RKNjWhtI3nGwKpWInhTDofRBiWji20SVj1341p0Cw0o3/vkmCovbRAbJgVvu8
A8LChaRGRVLuxLRSarH2xLhAajozfETwW4eOj7liO0Nhp6Nq6R3Ui/1tEi0hm+yS
CWXu8/RV0EDQOOypLpQkn9v5Cvp4vIz0+hUgAD6hcrInNVDWepQCSy/UvA3Q56ZD
zJWz9oXbjxu4MK1GWSIe7AOSe1gxfzFGxCM9HIBRnR+pJurYjbQBwF7Gb+0iAhw+
OR8vELQZKB4YEtqheNEvLssegEUszYBe5BG6ZXswYx7FNteM7Z7tRkcPyomHtcdZ
kntMXqE/ciRSUebOERqCUSwkYvRL+dhRS0Q9Uc6f8q9wEcYJ950RDKhxzCqFD5bG
+iDjXijcT601eNDcpO1qMGlACI1KNtkIs85Sl9CE21WK6CVwswkLjV+Xmo3DNG6I
Qkr7bBeHuEXwy/zxO16u/+EeWrhu7wyEtKCOAswwh4F9dHvDnp+l8ffzY25VTxBB
hLfj4Sxs8cq0QgMmD/R98gtrDtsR9V/ZJ0G4IMzHka4S6V9eL+mGFsBzj1xOrVci
yBlmO7z6rVpMVETRve6jvesMeXzVuvMIwSyp9gy5Wbw/UiBIq/65JdMf7xMtBkwl
lQIzeFo0GT44xRLxkclJjGBn6nXW5eeScKcftS1H0eR1EOfJIk1dLrib79bWm0+b
0tJzaO82CN68m4sN0TG+aM0CR40PvlgGpvIWVwOW4aBN2O3Tdd/AcPQsfaY9ye+D
XZfH9hUCvWhNAJwWJSeWcWZaCrICxgP2aSYPPgz/7Qw7vbKvCk7hx4ExeBefKepP
HBPRmwft21DK2ldyhU8vWijBWCvC7Iyz+LVRanBpemPrapO4u42pwHMjheAoCY/m
lUg3SJp4MCcbAEf0w0kVJgoqNEVSucWiYOf09c96YLoBzUfYgV0g2UlztnIRF/YO
+nU8iEjHZp+9Hy2P51npK7u54p2OV7CN9m8Ct7IrwFQueRyOVYnwV5SI1h0eH/PS
28u10p5RI/UN6YJDNWQoH5V/WWc5MlDhFldVPF8hs626o8EfoFWv3IG5zgUBYAmJ
K/PIAsRsbGnE7zZBn+/4RNzT8/xCcmdyirK5yeEl4keuTsmGhC6/8W4XqeotCgnV
x+JU2lxhPZSWQsjRSL1YM+T2QVhAvYpkzoQiwKOrL0mqV8JddvzLiuWxn1+Rlxj2
u4o+oYRENdBkbEXbmSbWjwTzyKRsATCkIDJSQTHaMkd6+s2YeMUSDlFO+IR2mqSf
UCSSisFxiIAShgJ7Ur0lPFgEo8MDKtKGTKS+U/iagci1yAjAx+b660XPh4n8L/YU
IFGWMMgrm2nMdIy006iPhpjC9gd3AcLUpWyzrfGbw+/3rijNvSlOmFSNtQfrgfyb
xc9oKfh3ssNcjx1IZB9Xej3EMFLT/ojts9P46eXGZJ8eHoTtLgbsiPzsAWt4SL+z
I4bpe3TOSE34avNKFlGCz4dPL9/7xobipHalwijI+yU9PGpO/yDVyS/z/SSKGlet
Q69AdxIQ6/H1D8wQp2K+HYa1+Xbk3MwgZY6IzVfB2cTRHaY2B3lkJlRfarRHkS/y
pAgDd2BLQwQY+gcLOUo8L2HzZ8eWw4Q2ENetnHkOaQsZShXvoZE8RhXh3RSpwO7E
O6cssTRXmaKWwIWufbYObtvEwEQYkJCfQVXby9qABn0aNm28meCaYhIluHsVRp6O
mBC87oVWhte4UpQgefisnXJ1L/btnEEkRbF+o6AOuFEF8sFDuCWrRJpZspOMhL8X
bjnvGyPdppOBM+DKlp69VCeeFGzEakuOZwZxBAIgccLzxQWhRhWU+cXG+1zu2prj
iSjWAmYmXorezTbkQo12eyiS83UuD9bbWJs6mNBcaRSKtyB3iz0jl2gx/DmXjD45
BdhjBBlBbLQwiEiD9JRbJtnIbL6efdwgVqELYHanERvz0qOsioqN/vW7oqel6FiE
dH/NLD+BkLlJioAH7KnMt4I5dOjSjFVgfopPNm6EglfCYBy9LDyPUYs4asuYI8HB
g/8gsF65fPjfZ0e4QMlG/Wk1goHI+cI6YcCxf0aVuhtizVe9zF7WHYXwlWbo5CA9
6oa+oHbuRZpB7UQmHdlYb95IyODqT2u6Qfwwj2exRjGzLopRhOZ3xQyg1Gmd+fnx
hww+nWExyOYXTRtC7gAQtyI2d5fqRO7RhaJYWMjkb+6JaGE/skMQhGrHsG6D+sE3
+QN6HtgdggAYWJ2HEsTPWIrF2gVSMHpUGoHD/FkYZhThOkuNEbu2H5A/BUfnx23k
3D5rJpPSaAzBLDv3a1nPMAuOLl96voHZKwJQJAsEwjoCWkHIObhQ0A4m33Qmgc1v
gArVMJhWoczcDuhg5dyrDWwX4MTqBqFmqLjJzUzqzc/jUCU2zieO0u6bgC9CtA3D
xDEJIiwdc/TLkuN/78AMjbLEyP7J3lDBDcMNM4zK6294hhPXDMjLduUFjIvRIj7I
BNj2o7fiyc7fm0jrJ7InazaPZdMU7ZwEIJG1A4zY08cu4F8mhX38AKIXbjSjzu9u
9RF8aokLZpYhrmwCsJQcUgtHSngdi2ixXCthXIfKMvGjYzlg6ecwGXbW/Pts7eRd
bwRNWQXCeZOVI3lbkxJJiWMGxPTAc5QLcd/yi/mEnPAXag/JHQyadHwArDla7YWR
ybQTWMQXzw+iVnoMnpByWZZuWlDi+TZ11kWGZKe4N23/AfvcUKoHegZj62ofQB7w
iiCbPRerI89KTnvgQ6vGp2Vl7Svccv/H2U4x2xyqArAjyF2osKeRboakmIvh+xMU
wLskpj76J3wtlkc8SXB0YEYSLwbgiGgXfCGPg5LPaiVphGxTekxf/N5YZysvaPfz
C9TNUA0+8XB+OibIJ8DNE1cB6/07iiFoIwURHW2Yww34Mv3LakNBvOx4S63lhA3O
dWnna/S0wVVo0mrHDBUW4Y6iJnw9mo3awDljDNdeDhY3cRtwDY2LdDn+XKyVjDSe
NAlnFcAvOC1klEvHY372tOgsMhJdYIKgbKrgesbg1f7pstDf+Qxg/BpMYPrWlljY
aB7KfRijbhQCvGvXvd8/VVm1SADLNVWmr82OXMpo+uliC1uv87AyK/C9XPNT3zr2
/LKIupoSaM+WhlzmzYlmzSur6fi5nPrqxDig8ut5Iw3r6eb/dK9DrbAjiM+/Xta6
WRYF29hB9LryTtRNtEHztaLVppK+cIxIrncm71k5h9Ba+ysuHrIQnHSGP9xIHF/D
ICR8hzPxHgAshXCzlkhjeI31lQpnXptOfyBZtjG3rvQ3nF8Gevfd6i5MhQhbTHeN
HaiEffWQ/DwaxizcV0rmMgngWTZO1ck+4NkifC8dH0CNZKb8uOzJeU70xhpACcRV
QXS2EEJ7y5G+8a6WQUQGxgxjLB1S0iOLcWSdy/RitCTJsNm7eMxDuGud8rgHPxVg
KhGeUKS/4+e0/oH/2CsPjTvMuSi90nVhl8lCJfd5VPZiOjCiKJvE7i1SZ/7HfFUk
FGhFc/+rbo32KRXtU6JAMfkqZyRf5yDSD/HWOxdC2G1I11kcieEs6+CEkjzti0cc
oKlJnEREgleVKyp7Uhj9B9Xb2mcJ3aVLKq1xRY5BqdFU+WFWbc1Az0/B0qrvzmOR
t26y0vuvcQVTVMsNSPblVcBQvOsRSUdYzOlBNZaZLdcLKO1M5MhQ8DTAGHGa/BP3
KpayAlDo2RvCQDF/HtVX/B/tVPh/QmHpGHg4sBTIiNHKecbTHmDg7VpT+3j5//6T
zxdym3GZdCh3QywY0qy8hyuvq8PLXdPXP6UbbO34B8AN46WfRf6wNugNYZkXcHZx
NfHfcjJQmywvCqNJxpnpml5IOzca0TmeruUutDyBsKAaKA8qjzfpZkOvdCbe7lg3
I4R70oGqR/Rh2ZxeTQ6mg7rmBN+N71gkHSkbEhS2sTHKYaAs43o2PkvTPycS71S+
xAJLPzgrmZ94/K4E7cy7FA==
`protect end_protected