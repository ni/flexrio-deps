`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10368 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
DBGZtUPdvgnvgIFp6VMrQayUS12cAbQy0qMlMffENAXIVOFokuz4nzHnaiJdalKh
BLozzVRsK945pB+Y+OBVaW40S4BpqpQdE6RH0dxTgzns6hKeEm3SmpbAGXZ5ZP/R
va+1izYPShd6fqE/tbH/c6NQ95zIX/LAjswV9nzJjR+1UfxWQPeOBrzithS9lWZO
LCFlUjvD59D2JgvnBjnYl+UhkDGC/2BcfhDpZ4zPSj9NVhwqbytc1ge9drk+e05t
jPHaobxbxfETbUZ36a1QacZyB7d91pv2oVDjVmy0Y+UVslo8tQo/ysg1XOkl0mSG
p2iWQAW+Q+ZfJJ5JrgJK0eYMUcjGF0xm14cqscO3yIondzxmn3+InDWzEQ3QfrlW
G/gfLm/PLQjclkSZWADCBNDXC8zlcSVrMJ7je6bqDCacOke4Hp4zkkZk0jFRb4nB
7GdB+uRcHdwN6/D97zjpSsRQSMwFW+Rv2OA7tGUiHpb0GbNfVZYoYx8h0SgpblY8
IpgP1wphgqinD+/eOUnVtjZRodl5wakRTXm+TLNrCy0h2WQi30wK2W1QLTQ21Imj
sbDtukknDOFaXSGJ1WuSFnnxrBlyst010LCAD8vizy3ZqyoFlsubjwfpacfHYfPI
za+hOD23E8VwdcZFCGUwZUFejvC4ueDSRxbgPjchXxr75CUj4hnNY6plIxHqvkoq
Q10J7cyFMwcKlr4Lx7hwqsIntTZHh0+fasdAEAdR+KzETcR5IfU4WzGwe1ikAjVR
DaN3bsAvsuVJJl0fiTh0XKQZrSf5r3Q+O/fpxXNTPRYvLcwkEAv9EBisuXkcjxC9
TR5eZWGUSAvVb6U0NnxgWW31pfZbF+KG+oJFGhw216O4ScjbJvSDUKWRwlmoxf3V
rNDsKK+291/OQC7nSVSdEk7hU0tffYt5L6nyKrkMfWGX7dHzDEn6BciGtWctVJE4
psp9h0Gb957P729Id3ir8bn9LBe9hJ3VHyJO07hwV2P8jdVlyNW8GLQLIhze3GfL
BcO/web1T8gEB5pR3u/nZHD4Chkzsipwf/m70QQFWWCU0+VXjDfZkDD0PQmAHvbF
aLe9/i/xgBgUKZC0DmfIY+f7uXjEMpi2VSX0fsX8HWs+NC6Jh1I9Gt2EPlaMAM3U
IZmOt2E5GVa3kTtBxLdKpuudkId3fVXelxG1/8UnVP+34PLTv7Y1LimYxIynzIY/
15B8cNcFu3qbKhzUID6ADRh5CBy4eb2Dv79a+yPQ6DWmWlaqLB9Ion1y+ZGsBkhM
qi65BY8Opt40J8M3LnG7B2rkz1Tor46W5A5ElbrzSJUJXZ14eaQPRAgNSHFRPCXb
QMQqYZtPZpd0reZTH2hyuQelj+XLkS/lgixYaS6GCQ6adzo7aDxNeE9c9KDycGuU
6ds2RADhi9h28u7imLNsWyLQHEsE6WL9M0oVp7CFqHrZGQrICeVmG7+6FHd23Z1V
XJjBvEPyvlilWrhxW+95nQ/Emjp2ojWVqe4mxJSFy9ezwzkQmsCUiWH2j+2dFjj7
OGt/LqH9L/yGTD+e9hLc5hQHgWMeWIzB1/NM7tYIOgcNxYBtJjh2Q+eVAXygMK94
cJXQHU8Lw508QFbiRyo22/VXkVzJZXma5dfu0Hl39TgPP/G3kMGHaRWPncgDiusO
9u1DCEy+XaFCa9VR6qsPRkx/eLQMA5fiPpl3YITWOpE3UnkPGo+SxKdJS+ES0f/R
Tv/Qsc6Ha4rL+yAHSQ9CSHXxFaz4zYpEkI9YndiI9rFJ/OVOCU74E6brY5TFis7U
Unyc/ZqeDzBcW/v4G/utkonmY78l1BrcL4Nmbv8AZScjBldRw9Ej+kCRkynJ335j
ssix0mqyFIFirmc9pYG4SIfW5cP1rIobRKR1LTDe1FCfDUkhBecwoAELOM3vcIfh
erlqZRFoF9ok9RFIbKLOa9tB4S4Ao/WdLQ/6OtXwGX+1nk2bps1ss+ysTEy9voPo
rqwi4VPVbfiJ9BgeKX/RZvrTuUD3J8wU2y93a5zbbXiI+PbBynNfUKpxL4tzcN3m
yXNw1imYkc6ORcq18i+c1zPRodgPWZP7qeHVFCPjH9nQZ3pgF7J3j39ahX8JKsyJ
l4rFz4BQ2xG2CEDSgLEzWrPnQFJnDKB+n8QRf2aNJAkMgzowwNzuWXO3YETn6irA
70a+H9AhywFyd1OqQYMEjRY0NCJSxqf4+IBHwBssVs+GPJelAC5FDFivWQsNuiE9
lhakNX0Vuc3MD08VholQKImdC1bca/8derWB5Hc11hHSjZOqYqvPK+Panxt4yJI3
qAzn7A06bUfarNNKr8ABgPoNuCyRei09E0pscGVKTzJTJq7EdHcD9okLSowhiUGb
CXPQT2Fo90/Yty9tk8tPIKqMG/f1MwQKD8jWSgKu9R0eVbtg57ORhKHFGbTKr7g7
A7Z1MixGj/bqFsXSUZwFelfCPMbAPfZdaodZ1PPpcLFPrHmw2bn9wSPv9VDEYK21
IFupUd+WrzmQWV0jc3oooZ7pN1SVReJj9QcX4tuiUn01owj+wui5YzjrJ6u9yMCB
QaGI+NMLvfDBTurBfV9mYwBsrjT0iWAN0cN2G0lRcaHVHRdMYDUT4gWMsgDKfqZp
VeH21YB/SXWVJqGwFKOvtwHT5OBtG//YONxyuMMOKmFz8hJww8y+NxkJquyqOrtn
k/tEKvFxqUSNoFbhK8zlRT8sLPeStyAXALea+uTuLkfYC41KyIAlabshOGzV4Rjo
lTVIJi2xX5CF0nIwoif94MERuHpRy4NwelO8JlkpL1X9G9ZkuYJ8hCzFuIA+0sBC
q3VCmSyFI1dgjz3ZF0mUxhHNKva7oPDLHKfdcoqsAo8WlMwhxiKLNA6dalTk1hDr
AAVmu5uJFBOPzW9S5HPnQBjvZk7CYd3BVw+xaMXx7Lic3eXVrF0kOchMcozZpi+e
DDPYvFFIYpDzK4CPKZYHeMszUsdtzGYmLo3cSKU3qKafD6sVqXD6xlLdy+CkJYDL
j+iJtEG4IL8liClu5RYip5lL+3vfAteeHQLf0fqdctHWu4XN4g8K+xQN4spTJ+SY
mLdaEupMbCvQvW738Nc64q1/TT+ZDhTxwJVWr1N6PmwoHX8f0fzI5dZLDLLpDOId
UEEwYNLj2JrTUgcK99fXKBuWExjTp2Iy+LK7YSyw6P66q8TyaWbXhp7LgTA4U6uY
Lba7xQOMR0YjJSDSFnuMZMbGXTzkjZ7EzPljAbj7QEDLoDNDsywM76hFcou+Q4Al
7khJFn3zt9rAZi4WnmnRG/awaPKoh95XIFmqRiaAiSSLLZW6JKKLVGiO1XmtCmXL
jQ0kif9ibTHL3vqSl9CR3IuRM1v4cBNf0x3gXynPXAkPjkneW5a6LDXTgt6c4PGR
niruFHj0wfa+iMFyhh/XVG9F8d05McUR4Y4jxtnuDHEuySVVbc4e2xRGKKoFQsHi
yrztE3pL12A4fMMat4sBOJKPn1N6/1MfC2w2Boz5qVQGLeaGWJLyjK1/vCDUqlO3
QP3dnvAVHKqvmKo9LzVpvKzeg5IYWqxEBLgXhl3wwdUNtbTuEwVNwjSdG+5PjHH/
vjF/hfZCfZMWn6CDAIINytECJLtGa5crVzxmiVOtGnVutFVlB3jlxEOs/LatqmgB
eJ9fw8MsPFwmgBE9i8Ba9zJOTIC1myp3SkkjnuIwmKfAHgvTk6uT3KaIaSS2KG3a
cZl/i1bo0lATMEVq+9ZY6iqKG3rd+iiyBH50/Ji0yySY8dCmlwa8iDh6g0h/CU6I
3cq3U5QOr80K5Y0TvpK3fUevRIX0u1PRJBE9lzGw7i51B6dVuvw6WBhsBnKelo68
8Ca11kp5eh3bl3IesthaXgpJh9862DmA64/pnO9px4il6bzPWnr3oQZkLikqu2Sn
UwaCL/GzufUe2GiNlgKfS7Qfv7MalB16usOJLoHqZrYrMvX793JgKFViLAg+8y9x
WRMzEDgRY0ELpfslSluUGv9DazwhGs/ArTCpIR0iUaxl/oCwO8U3H4PW9fv9YH12
gLJo2k3OnVA4UkXQUsXYXfWvG9oGLT6U3DHD66qVSPwwGmBSzAIlX01Si5P2v3oD
M6qYV8h0iIZvRO24ACNewWcrDsyot31tuWM0/QrfglFiLjDDT1LM8jgB/DKd1JtX
W1GOmix4gmeXgNTwwmASbCyoBiJJv9C2HBuky+1TyjwVZVomVasJnE38lZMNLt9I
Kh0FNDWinXhP/6peBbpB7InpIesesrhfYnO36K7QkLb8zfWf+5CIaKwXoxXX97Bq
lywnTnfmQsyQC04PzNxuTg2RPfKyUKsZEhdFsvEeV2kJEaXxjG5gojZV12P68gNh
BU0nA4fWUPR9jgjprKV0KGwdXdAO0teoOpjMXTaP7OfSz7n0Q1p9ZO+Hzoao1PFI
zXuAOLTRRSYA3/4a0YhOXwiXskgMiBx9VJE0GpVYjaF015efClhmyuPxbm+XQYit
KE2R15t936lzBIOE8TqEbpppGh61MTcLrz+Pai1YPd7pnWpRD9EFU/uY54LfSMYB
rrOzThxcGoo+MlX9tASd7O8HZYS37US3Q1kOod20rQt8kczEraSkNqV74gRcn5iL
ddPM0E9gKljndEDfIVZNRjcb//jt0fJNfojzpUlfypB5KXdyhnF/+2h9sltqQcaC
/+p63P8g2OI+yx8cTwr2kkOZqRvRmYX/LQ5QnaNPFUr+l/tPy5s4BzOTwh0dlPQz
oyYn0MegX6+I/ObBDvLUi6RXQMpYFK00oYVjYnL+2NxoDlm2E2q79BNHwiFLc8f4
6oLDB2a/3+54u426lwitaNtY1yivDRY+wB4LmGhLgUTyTaTAUhHt/0wcHmNyJRX2
XTLWQVui+nTqasCln23QmQz+Hln+VP9/+ccuAOWQrljUhXfpwTS4QOzBl903SV6f
rRi6BUcHeLRmo2yhB54ksm6bbzVEuKYWQeOyJ6ttVyqLVELaBjdnFazvLslSYoDO
k3FBNoikbYv0VQ4tsFmxKGdx1+thav1Yp698B4Hd9Glutu+5WTwOu4+HxvI/YVLP
cd30X9XRvM7K6+bddkawes5BLpSv/XXozkgKEE+72oiJ6LIxKqPQAMqjJUheZLYU
18GO9Eq47IVgRnoqoYDA5NahaAzz/H7z4drF3DzrSaV+PBmJhMPW4xfYffkEkuws
HEZTw6twOUFppu2UuseridvZ0I4BkpL+LOlq7wlPY3VAcyWr9z5wC3uOQlUkky/P
zT4ZKP9oru7gzsKoB6hhNDkBAZjDv5C5+3Edgmv9Zk0MG8eeURHQY20N32p5Eo0j
EWh82RBOT70jy2zYPKQP8NdOu+RDvQfwuCdL77IZZVE8el9TAjSssA7BbQYf2HhO
8jmcf7xixGJLTtkKKggoytBMcCsMsvmWWLbGQdkLNwlUcilMtbGwUZI2BzwRJU6j
QOsq2P6ST48iq8acsAa+x/1vd6T8QOYOxmLT/nqqzpeOYOybOLfFU1Q3EgFGOCZ7
abMMfXKxVTNdxSJ5u+cQjC++iR6R12verPMJpSuxPlXLRfzrE7gY6By1TwjsbxQP
6wtAqASdIdQyPlCasBdcHtzdJxkIY6MVD2SVT8frDGT6Uyv+HZDlFJ3jOMaJ06y+
9lhkpNfXG1cG15Im0+ggB5iAmlgSRMuTc+NGiDw+ZPOiqJLvp6e9EXbb2yeVrrzX
TFthsXeunCXwYO1kUvnpje0NU5s2NasQoS2+m5YMDU0weoAO1m/eeVzKUFamCw8C
88dWN2An1cznQln8US9RwzsXFGt+U2O0G1k9PqNCMDa0+q7q/T8lWyjWFFip4Z2E
geVZc45B3vn1eEUuf+fYUeCfw/QebOiky9ETJThH65UbJMUlxna/xBezwJdcEiA8
0dk5nVWlyuZlTV2NnfIx6lOGoZuXzvoUTO4aZxb0lkvBm7Y9Cn5/BpgVkbAtVHvE
j9fZr/ngArJK7ggtaSoPal1sAODrcl1xkYnGm1xrbE9LRL6bF3aktXjCaI/BJj5J
05gsGei91BlAlNK6R4NSY1TUIBssTEO2D+BGOd8jAmbyF6cnTSr7iGpaqFm1RYyL
FEL3GI4SNmIir+gXQzwDMeQzzSszUEAzq5Kyh82i5OdxUpyuNGIrSB2R8mdAnHXD
kKDr10qhaeLm7dYoeDDQNQ3prnFhuXxbHAYV9VR+uKTMDctEHIWexPE0F9huyZKL
S7/CJSUUkloYR2xXk0iELjIzjhCyKAo9MAn6IOx6cogyZ6QtKMgDBNVQ00CXYhe4
BzHj76+hR5Q4y00L6IlfYYEXpFlbRjwgjLKF/HNZhSXohOcZ1sv5o1fOj8LLePsw
ZNdb9wU8fnDjYwM/7b+h/QHpuWMl7TTca8c3BOqt6wh7Dp9vGA6oJSMWLFyIfZm1
Zgc7rF35M+U+Cmpn5CgjaGZJsyXfxPyQuZu4PkC9zSJiEWFe5tozgk0DNxoP2Njv
ypEWSmxEO/P03b2A+BqaIsAM1ZivFRt7ZdqvINEes8TZIEkaaAbYFXP+JRH4EZpG
3JyIFH7n5ZfQ6qqEeJlIWv1x1mVkLIgINveDA/zQ+fNWnOXWQW2kVkyvPsRDSZaC
VkgYQSFsy5NU+LKECJ0KeKSCHUMqYIYGUupObQ1cm9PGcEzMsTnIsUHrQocLjjMg
B+jICxwdNy3irkgna0pZ8wGEJZ9fkvax0GOtkcYeaxgaAZL0wKUswRUe3u6RNm5q
YyW4A6ewqFOsdEZ50a3eRvyg6IajP4cqx5o28gUiL3x/sgQZxZ4ALb9W6jh6HLqN
NJptHOiPgG3Ehwud9DNHgqGEit+a8g29LJaP1jIMoz7xk2IE6F0rDK/3uK5GVJDo
UcrzA9UJH7JGCx39CHI8BkW2ATn5OwO8jRAMlC+L/xAAR1Hd+IgEFZv2vwRpthN0
hZUIP/jPN7zFBuxClAPboKQmtm4Bk6lvRGykWsrzgQzmq2Rv/nNRV3JeP9wHU4DS
aIFrtvYHBksQ/mpTiRG9rNaGRim1dlr4r7evjuI8sEmIfXMw6S/NE0EbSWxzuaQT
2F6uHEGGwbsGBO9NqAujmJYux6PonWOMD0SXTL/Q771FsgUeOmlsrkQkM1V5la1e
CqiL8km1fpz3d42vKdL2SNaGkQTWzW6pcxzttWTQ8nnnzgkYCRDnhtwqfWmnhzJu
5/SRlsdrCotYa/F+TUKhfqyFIjajXUlnEBTpGCrxuA9RM6+hrUOhfDn9fJ/JTQBA
0/9R/kYbdMbUBrI/xSPNyBZUN7xLJFIB+M3Ksi3FGQSbRUL1ySJnXzk3aYGoWaCu
KZwTRs5dAeEvYaIs4D8jh5Haxtv5llzy9l0eiuiaNg9CIePDswWO7lQBx1shGsN/
25NryTXAG9Q8D90KmPvhFBWPJIIgNtfVLRYURgdLEZLWMx+BjZUlKZcsGUHYn/lg
8pJSCsMonnKWwCxwOBo87TGFdbMDF61Q/d1BoO3oBEHPU3JMQ5pwI45aqw0UmCfw
SO5odd2xUaCAISVKL61IgnbPM5Fwkp94bM8v0YTgGi+0ii2kRd3BPH2zyEbS8YjT
ZBYRfWB+wlP2Q935yJ3PvH9UDxRNCFz56PXH7OtiQiMw/iOKEXDv05lvaIIWCsnw
AjvDmRahpgVAKVcIjkaT40G+nbWaZ8L+IzadmTvvnltC6XNTK5hsYC2Sh14Ou8F8
WdDM6/g+ZZ3wpWOhvmADHQ4FxUeBYfDrrSWwH2+LfWN7w3ynNbDtM14bN4Ri++9o
E53xihwfgGodfncRHR4RBxGEB0dX+T4oDyZSVhi9KVim89YN9wIelq88YikEunK9
xct4XyCeBh+WcAXOmX2kwLiqvdteFsbjrrT5sF1RDWUMDUeLcuZNTzAg3XKi0JLY
0R+36KAR068Gyk6Tq2dpbtU3jQxPwSyU1dqMxl2+j1ljsNNgRDyd1Y3WXl15+drb
m3MewbYe14KiUFZrmaKcWdtLAx37LtIBj3txhTFRkA7HsbCiIzCLZExf1Ll/Xza1
viYE5L1DBropmsHcoScc/MdAVYE1uMI0uXbD9OGKj6Ljysb76FrvD/koZe3XNP4K
u9e8NRFvjeuBLKiCLUkC1aJDhWOvJWEBJw8PhHC6rL/lAtPRAx9o1M3t65hQSNPw
v8PYKuRcMx0CfnxYSDyQeNHDZZVxtKvB4iJZOWpymbIDMjI1W/QpqBSqUpLAHpVT
FySoZKjyL0AsB4lNrt/TEEDsOu0C2CANPMly87COejhgISegkIgMOFXxC8GhRd2E
VAygtAL8BUwBTnqrwRmmnaQRBU01jLO1G6ZQkEPV95VPn5WZK9r13RFXlDAsqvpW
df/8RUvuyFWt9C+0U3o5Pcc0Hip3/9I9nBLDcqX3N+Lv29p1VVnj5jkL4RySnQNo
aIe2QYo90NHhAf/ZWsVYuKsj5diGYScAVXgvPfirG+3IW78QG0WcrjnnoDinKKfY
e272FQLr/IHbGq0LKlbyu4y82ID5F2dCXvBe71ITP7JgBtT5VE2ispA44HVF9Rbg
BEhxAepKXLzoj5oHgmssEdPG9kFwdjBbm0AfV7tmYmFvGJhXfC6lx/UDYCWrf8bc
6elbzAc51vH0PPQUiQlfrn9dVDwi61FnvdaEWJY13JdAn5IFYDajhGZJP3nvUrJo
2hVhLj8KXQK+T4rbwon2+5sskQu8dgJJ+yRf4fBcXZet4jwuyu71QoKbebH5XHiH
UAdbWgX/XipJz6Gvf1xaXOWuLAqJMbuARbP8Uo4XJ+jp1whsUgLfq14n6T/d/p08
ootIHydqWh1QORM1AsTPnlDLhDydl1EfvWRWowg1F5mMtpQQL8A7V6bCBPegUEdJ
SDACJJEeI5YBnj/nauJHD6z9+Z5mMsasw7rzL4NK0Z3aP1kPP9lMOqUuAzUDeTbH
4EQH9XejE2Kbrk2Fwq/PcfcTMZejSSeI90FvwbMnxOFY0HJ5WS3Zm9u5sALjPhNZ
i0nEdrUEcGIuLMvfm4DTXfLYaZGbhuY+88mGgEKx2/C395d6qpdlnakx/Tb+WMs2
4dyY6OHAOsKH10K2wT7psWrTJCmfPTcE1qQwDbDOVCZp+cwbbK2SnwpfiXn/Lctg
oblJETlvc2oTG8XH1J5Not1eJVALDo5jrq0j2CgWBBuG2awnEH8y0Q/iC4Y+J+mX
wdm0ZrRtJ9CuTBhWiz9H6fX7l5NGDIwwxSOYaBUPYY9U4gBKy9WarZdkRufxyaJY
xl7GkT0+jnUNJTk4bJxvtX2blomOZsp06BaPyZEG8SFdAvJMavCO+6YaUQteC8ZM
/uUj/91vJ4+A5IuQZ8Ms3YCHbsRhCr5NM0V1LGz5MCAfEWL/n6H8CbD8n1ZATNrv
WdYttW9b8F6Uqe3u32aMD8C6Qs2M5Gdju+gaHpcOwhxmWT1pgeKUvkLYu/tzwe8F
mOd5i36v36ZX2gzi1UlNlt09G+PAwQ6Zjja06WqvSQpKmSvDgYBr7tZkzKxYpCRx
QZ8e2dgZQ0FTdVbq0Qj4UjU2N5x5C1JTi4DI3rQhPsNmcmqtVrmD/cq3p+hoW81Z
seLLpn3ykIh1aK8LIJw++I3JSmOX+bE9BYfFN9S0NmgZTflMSwfNKaHxZ83OuYnf
geD6SqryP1ufwKQ2hdW/V1VcnBnegUbxgvd5nm4+zueiEqqFi8E9iNbFhL2XMlXt
WHpqhDmSt9P3YNdVSVGqVp80FWFWlT3oZOfPbC4Sh850Dl8ABLM0VNe/X0EwdI7O
IH1eMIkZQ7N0xFEtD9DUoAfpwPdAUIi1i9lEAzIkhFmtvRWpsGazW+RTUbLZ0AdP
q8qVEX68VT19XJqIKvQX/zi1xphCKCYOzM4ii1Au+2p6J27hKJ2AnPb1NUlwL2zF
UpcCIj7oAw8w8d46X1bVL9/mhLbgrrtDA02xqjF22/Vfe2iergsxHRgz0h9UBfUv
vk7ihIFIVEmdVNn1H8qboQNQd7D+lvKOqhcRYMK6eAkyeHKZkxwUPz1ukCrK/J/M
kIvH9/CYMW0nym9o626vLjaw/YB9niVyC9ona6Qacy5V/D++S5kRMSkW2zIqGwQC
PeuYvc8Gdoq+9jBSRXdV0BxovFAAvREEg8zvAeXrFZthLblzcFi3Uw9YkKlRYxyl
tn5izvjl0bZ7ihOX4UZ662fmIGaXdHjJ+p9kjEDfGDcMiNLRlWc9x8EdUqXL2lD5
SJ8KMCyCCrURkb2mYITVnTfW9wBuV76ipe8rkZuAB46i9AI7PMUeQOP77spLbSlD
UWIH2daDsiHiTd/xYGR3ISyfO/kV85iTzjkhJPzaUvyvidvGRQia9jb6NrnSeDK4
pNCJsOBGaQ3hdheMZGbToAJAZ43DipBS3+xCfuhvpCJrZLa3rZ8G/s5vjdTgeeDU
InlQTkO0Db7H/4gTkcuAm1fmBLpINeN89mcZ05cJGU1POR7Dah1OHXCMs5O9Hr14
g0zB7gvSS97zQXlMe9/kiztvNDtLWLON9sSOLS2fs/y82wMhQveeGezzgaCjlHOr
gnIR/ctiB2kRApwCKnSsPsNWaBcjACY/pbgjInfIcoENInq8G7k+m1qiWIiSetGr
kZdHLXTro33DHZ1Pad24TYP3WR0RMP7DA5YvZpzs2VVuQ/IcQVN3TO+SLcxNuyKz
JrhxKD0UKJDRQ5sh2vVE1AFVn6zdIdKH9yf7930ew1yW0KhcpC8OgHZTWFcwIJ4k
KaJcT9ZpFsgpZ3GxIftVPvuD9OpaDKJwmNywHb8RKcrrwBO+3vEans8byhGlleXj
m8BkGS8TJQwol+7Pn3teGbUJ9AYjfY0/7i916Ab2nqEzFjAtf/FKNIWxKYvdbogG
lK/Hb5bA2oQuMkxEDQETaXUipKH5KHmnNN43GndsbxGZfK9U+qOmfLXW5rGqXxws
T8+WRTAErGsypwWsAAvWbA/rCikOCypCn+NQG1PFcUh7/Ia+iSgm1XdXCkWkRWHH
ReNpp/KkeIvfja/rhk7ki6eYOgdCX+0+Kh97PjERWtzXD4qg03AGR47YzDNJImEj
1y3mRNLrIfCDIfPHcuOMSGYA9P+8ap4sr1PbMvz8PEIVKTZQOx8VTetT1FtTgN5s
LF/nvnWxtXtiH6vrlykE8jwtP5AC/+/h3S1cZBniKe1pQTrloh3ABTLaWq1IlfbO
Gr3iARGmke/pd9D2U8zhK59rvnrfirYtiPQSVRsCXszj6Tl8o2kxNF4NNcaCSnVJ
/i9mDaz3pM1P/Mmp/Wm/KSuDid62f2gJ9OaT9e8yTRPNGNqRMee+ee9Z9zciMJ3+
ilA2RYK00vBY/vkUgPetNWaQps4FR8ktVbM3swiRVnTUSspjHYT03JYfI8btHl1o
Rq5WpScpM1k2TC9cdE4tfwl4EHZqp0t0JOYzsmemo4qJRWP+SSzNz06L7Jn7vahV
ReILjCeI84UWrRH4kIFM757lq/rKd0bMyqqvq3FK9yKSEQW/07D2CncdWJFpNt7l
JqK3ji4+v4IVHJB0wEnoeS0nDfrsZJ/rt1Ql5ZcaWTYGz03Zfg8VIlVpSH0yfuvj
PRQOv1wbNqL8MHiZseT4K5zncqtgqZuI5dDIfamc3tIvdamrzm4uKfHvPYhmrXTj
gfxgqG31BKDl8z/ct41G8LkVYr8Kjf4s/rvzUShoUnTzBHDYZ+UP/ki2XQo/x++z
vxbAUm3HpetJWMjLwjg0w1/1ZUDrwnW9eIG9v9BwF6/rjyKyU3xeHR31/pXD8EcJ
UpsXglWCIP0sMhRuCmQX/ENCzWjwWJ2BFGAuEHUjmlauRqDapAHlBqVXUrA5zsAY
72a+Dn12AWK9YtSlUahYykRsNPkx1pGy2ErDaDIvk/Ewg5EDtqK+LSUFny/H98lI
iidroAuqNmIb1VCgrfdjiGt8y6LmrWFRnXfaSCoNag2MKR1q6PWoc5185PhawQHe
UOkvETl1ouXsrnKKl2lrOrQSuczLhTHjapKYWUCaAR0W1meBnurUKO0+jcbssIgO
QMUNmx/YZOf9J+x7l2hSo8yR1CKm/z1yYeWFsW+GiuK/AQlPtl90rxxRBBMAUEDT
Pazc/hFi3xITvEZDo/InEhykYRLlQ3agKmPJjkZzr91Jj+5MCN2YBvSPF+DMutp2
fHrog16b7SGxmcDfyShmID303hf+F/KEXXbd0tyq6u0RpswTAKsob1Rbkqr0Saxf
NWrht3p9yUhpFW/k8lAFIM4PAylK+zabYESj5aFpIuGF3ibjQjAichC5J+VymFdF
UWIA6hI0biRLDCBko0zZLTHC3UCubDjSzjMyyampcV0SOoEbaCglgtGn3xFc0ttc
tNMNI5NK+byWfxINBfIa44Al/gIvo50CF1GG+gbtcUrlx6wwqeza2Zy2csIDZrj7
ObzpGWy3hB0E0J0EsSZE/XIdQPmTcxFNxPcqKTgQGKJBUEHtlCmFNqQYWi6E5nmw
ai+nE/uP8w/B2oZHOFq6dRV/sWiWwatLdtfzbYhA6H3UXUnBKimY5lXV4KXB4+j7
ktv4/pKTen3+viTtKmKiPJDIK00zOEZXQ9js+G8iJZA074gFU3UtNfqHzjxZB4Jl
ZP6dY3PshDiFfgoldxcbAvk3FpBjdo8ieGFxUuswYrJ3GzCMwnTd0H9L8kTIoI4C
yurKJkS8ZNwWeezypGXs2USrlwtU+52bOgeLvN9w7Wr3vFGiRSMGBKB2DZCdLMDq
2kCJVhJX1s745eA7LGoOlctjTC2UhzfmbS28aoGJAHMzVjJf34Oldxwnmit8o/ZR
+Jsa46OAvWU9wF6IPYDKPRVyzluagbBXqgdGsnEO1bAxHllshJQcvLedQuKcdKug
zaIPlHO4E5GL5K3ku23oK+u80rtMQ/x4+3/l8H1csr3Juij24VVJxtEfuPpmJWaF
EZZOu/fBhECJoPHcgaF2PziRzzzSTvYvz5ko8WfP5zoi8/kqiysOWhi1J91eFzRI
MhgkE65vDFVidzQl7KIvQqM6GU95A05WYHRjZlh+wQ03uYCPbISyxbZYRWXlxxjm
0NNzdPJfa7+3ajAY9486MMg7JGhotPN5aoDNIXhBBZ+hum1KBuYCFUoBMuBeb8Qd
CZaBRVfF1LQO++KH5u2HzC1oJBVQkkFzfEYhTnAjoZmKZknWc/rM7sT6SiuAF6/k
O6nG/E3WsQCblE8op6DZjsVOmbXd8+l5V0QPlxnD77/uP9Be3y2/OP38tlZvP0uc
deqWog7wgogs4zbqiGgKmOnSuwWa0LGRImNf5HJITWkeSGnkYQ5haYk5Ije55yPJ
J/VPu1ybJsYM+SQHF4DE73sgtX+uc1Qd+4lSexYjOLlE5cu5o+nAETclhtVR4SHW
Fuvbj27lOENz4HKpz8ATbRjbwXinFr5h3sZuKrdELeTcFR2Ge4/Cwr5smWZvrCaF
LtuZVpx+q27KYtlh4XoyQYwRKYDcV2kgFsH2sbuy86EnBdCr+31GQ7UeZ1jVF1Wv
7lt7tdiYLvP1IoRDKfox/z5zSKMDlCQ9mN4ppvY31MVgUVVy9lb7WzbWBTqelOjt
VsrG7VxG648STjOxZRzXpVyf8wtE4G98M5jEKBIswCzcButGwtyMuAE/HRuHYoPO
gdq1zkMBhRBIT8QbJzKYTvs1KBTsIwqlHoVMZgq0Fi6vVJsgpT1s4HutZaHQ3Uu4
kLHZNsdjGlFzICLRUIai9idARwmkr+FP5e6lA+4WWFKLkttTiEqeMqDDuF8r/1it
`protect end_protected