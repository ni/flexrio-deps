`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10368 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
GgG2UXwpbWAyDgGIJC8iiEUFn71cG1bxQH2TmDv1l4vBvFTI7JW3TRfkE/WHaCtV
y1sImQnayQj9HpqaaqM721sXu/a5wlKocUNpfqwdkBSw74YHnrslPmsxgCKDwsAB
gmmf/8hVQwIjbnxKE5z8qicb6wsVum7OnMK06BtdkdrYJ5tM0ro4R7PiWhzHIrSx
of0RVPtnmaaXJqR7fpWfq0EuJme22/LMs/Hx2WAvbR58AS3PJ7UzdNMw6Xfmad8+
wA/kz+oFqKBRMwXr9E6oRgotQSJfr4ys+10Uiw6bY5HD6go/WPXMeDUx/RXk86df
WRiw/1jhtPaly5OJRv8m6W0SdmIB9kP28oYcSKnlVHvF0qQZiy3LKCtBekL+bvDl
xegKCb31ogA3uBEieBvWyZaWVbFaKWlD4PFEF1hufupBB6kHf9UNL6aV/EAIIIlF
kd4H/NtXs/vgxDq3z1JUKhUQoc6VzbpQKYtRQ5RRpdc5GQ6yh8h72gRJP77O3d+y
HYcQH6zUqlRVHi13U9IgBfQGlyZ3BBvdkdrH7JjSycMFmNkisudDyPLtXnPMlOKa
R1/ziOE1RJxm0GPywuhJOfALGcvetBuDaEl7W+9OQWsJxMHo82z5CDKs4K5RL9Ua
/Rb2phBoj+0tnzYSJRcopJza+ogSW/O3dqjq8iu/kvdyxspu4OHyJ98+QwQ9y5+w
gOxoHh8KBXaTcxUDlyNd6speuEaj2KLZEiVfBXvHNjMPmO0OAexmTiL/0iFuAuBl
MBFKsXk0e/0sn6fWBtJ+OV3724601lh2OZw+9Ngt2HstnYTWvm0otFzwMrG79jFA
M5Hl3gcrXdBZxoAkTp3lGNwbPnDdO1/KqMwU3/30cDuCHOf+pLOCwnwjhhDVRvHp
GNxI//m0WaauNfkjY1s+mfjZawlJPl99wSvKQzpanY+9npxoVvi7ozcy7Lr/rQNI
gSHHKLTkRc0wo0G2WlCxHfOjxXaHrlgSaGyQW4qlyeVtWVgKevU094FeJ8YpXJOD
metw+gLARkhPeNoDEOUtjhGiYoHuVRSumcFj26hpmQ3LOzzgU6lPUP+EX/Aj9IHz
KhRPHRxysnVR5hnFTKQAF0NG0JxHw6Z2/xP5CNJJfXoEcgnmQv6jzNgce1xXrE12
LBy4I7F7Uqcjk/Yyqp2GnCzmuQx2XoeJKoiYO27Qb0u3HkyQD4EClLmg2fJ83Clj
MsvVmkbc2C1+owuCiANote2051trUYxn5hhhkj9l4THYFyx5sstUsIXVVGHG+Pv8
GwKLEvk1nE27DQbk9WVWyhwPJ2+pwwpfy5da7U2NWcelP6E8HpemMKspjtaThVg/
zrisQGAoL/hMyq076Skv77wuriN+7WD7SF+ZxerbZp7lkAYUySO2V297Xa3jbTCS
V5tx0GxS9lz9wSdgegL1kUEKZ9tntE+AfkwJHWL8s4sJ8EPXqGFoLJfn/Zb4LqYo
6/CC7JHWeH2nPmdBza0/5pF4puOx2QWqT6cv0/VYwkfvNbHHE9zB/KXrnktLn1dk
cAN0H+3VYjp7AbtznrDGnZ78RX8LsfcJ48gXIsFkFgEsbINS3GY7WFIZI4/6kVBL
1rhp+eG4ZsHuMjllbQSVM7Im1QdssrrHiS6eP+HPwLK4I7qYUmQw2kwIt+xlWWUL
kvC45tlX42gROPAMnqXMUU8UprbBziBErStHojIZAZ1xTC9xXPvk9l0uqcRYnF8/
Tj02kZJ1STMWUZb1lNMPl2lJyl+aI5yyaEOlrhJiD6riUviL7lJ/B9IfmJuEJ2at
IZCRdbKXf/YZnf3FNmYi1UO5/tmQNPvg3x7DBC6lG0ih4u4SXUsRyYnz9HlYRqTf
5RLeZ3rf2yRtWuzsLrD7UpV86aEANACGpRRySpMYrLydQ1YSJncnWajBgRzv8AXX
5XTTWvGmUQ5PUt6pB+VmWpwB6wiHiytAQmZ9i26c4zaawpQJ/zGlbG/MrWKGNGnV
g9HKR14jhlW7fycgVJka1lMKZ+6g6nvxfS1B/biL4jsrt3vKQnz5VTKq0B4dmke4
zZUXU5ZOFiy7wKsJHypuw3DHqIZ/JY+938EXkC0zpadxcQwpDu+6q0dxoSGUdj9C
Pm/yQEWWyBm4UdFS5/hhLjT/DNW2nIuPBY04ZcrZQ7XRIrZMhNJcVsceQdKAy5rH
Ss7HkUSjZlX4oWcXrPdYC8ekjpp12pN1V4YiBX6GM64aPqnoNpPI49lc2i+iNvax
WjDRyyGhaQKFHegTxvbHNKtdpvalE9rcd1ciRp/81S97kEJrebkSy/U4Y8AbGjoK
vHAkWAGgu4MxJeN0CfwJEMjMJfTXwjxcy/25K/GqOP2ctPc6wdkoRF+Ha7E69qfP
dJEAIAlyjK/pOdH1SPKj95u/m8XuEzMc5sBL1sl4UElXvp6l6aQpE2pyvoPXY9am
/94Lf0Ju0p6GrMy5XtYa7R2w0eONtjt2K99Bu4cyaSbOaNJCwD1cM+YFuNl9YtWq
8xa9VGk4HlMiXP7GJj7WTDr2+8h6feXPYq4iAGkHjoM5sVhX56x+hRtmXX5jXcte
LGjJ4gK4AdD+bqQz4K48AYeTkG5yQzM0fw2A7USJ0LmfHq2s55PyBb6xR3gzuiWA
HfapBXu6QDkpqw8P5PgsJhKeXSs9v3VI6n5UViYIjv0gfXdKw6lPTbqdE4la7O5g
4mmswm9Z7PF9u7o7O6Hhfz0vqW/Fs88iGc9LuvA3dXbXaydOp6m7AAVGi514oSg1
npR3tbocInmNlSn1isyKPRntcjAc9aFb4DFhyAa1HwnD2OtPnVBV5KtSSgcT+aq/
ankuqR3Lb9hxV/uCDMW+o5rBGZkZq2w/zsimSrGj5aX7xiSorWEpPkTYhie5bTpi
H7CxMe9MhwTdEsU48r5ytfTth/mhBhPtA73YMqINfOxXhQUAQi+vP7A3jjLw+Pp3
4WAQZYPHnXMzqtnPSAk28tNd0ZxkLphSsKtsJANCUL+ENgwy3bNt1InXJD98tcQN
wHMkoUxx2de/VHSRZm0f9uGIVGabpUf4MD1Xs4h445n77fTBkIyGbSeGzpz5dQRa
M3kdOjPxY20aAhQZX5QvaH5dgu33MAkr5EtKx8BkWnbCnRxjRbCbl0tAun7YsXOc
/9pllU1koUGNcizTnapBYSV0lTJBneFGxNYaFLgZ4qOUL6q1vTiE/2Yfgdl5xEx9
iN1XSkxEiwFcDjqjPVl/OnwdmWPk+tb5GLJGAijD8ntIVlgYu3ym9KQtTL2Fizih
n9/nMRC4nFQGmObIJFl2z3w9WQQ+hlaPx614DvsmhJnuAjWbUBAsRnRXJDO7L1Rz
ZvdZBGbIh1EXpnKTlrqa+IWQh9RZhyGBwT1O6si0/xptBrHmhjG9BdFKSXpjxnAw
dQ+nVrEZhwzAqSW+ePTfVvV5bLsob1rDP3DgP8APv4q5ffHD4AScG9AjwqZr0qoq
3aYWNQb/wGQNuUJ84+ayt9f+aPPl9X+SBT4p/sbQzYvKPo81pTp5uxfDX+26mo3o
oLd5yPOmq1r/SPK3T8PiZ4C9Uwreo9Q8M221gwCCHqgP+MHlCpI1KKelGP1gByGB
pPI0wcvNqojgtIefZUncqfH7M53R+CIwtTkhxI8iWhh8AyHAtDYknAZHU7oqkZso
BXUBwjQ8E1JL1Gb/AwvPTqkqccBAdoHO2tTOM7tox3qrJBueiwxaL8kCGc/PIc4/
UZFsGYKTgPMMq83vBmoFCNW0EQWtGJTVgOL0wHHG/KSeLlvziKivMvCugCYSYPhL
sZyj0saSfyhRdEmHZ8LeC07QZCL+aLhK7Z52v/PkWrbzsiBPN3yBQK34XE2ZxakR
UhiczvX2NrS+cDXwb7Rz1T33taiiFy6vM3BgHFJNL0nmRujGylTiniE/ayn9Mqje
FYwQK4Ap9EJ1GoSesXQQ23OG728vzTbL/K1PG+9DfoHXVUsauS8SBeDprlV84sxi
hGyU5QXmE+Av9FT1zmKoVm9r3Zko845jEa+PYua/TRdg7W8ptuCJupXa5IPFFoda
Tu78yrzt56any2D5qosb7P1XqaqHB0/vzNGyy6CqrlkML6DVgnpJkLKIa8hlhsRZ
8Y5v/kEKtQOsUmC/VEtKkvW5m+nFIDrXTzHdf1FiKw6hiu/9+clug8lpUCRekfIE
QeAa9IdTQfCK/VUpD02ITqWaeG8jjMtpzyysob09xfrHA6+maDC/GqaG2N7SebWl
FmFsBJl6ZvhK3ezBIsEBrWN1xHMMgVdGS37RcEhdCJ7+06YLmB4qUcse8HyuXb6t
PKZWcfamwhGeGLdKGR0Jlm59lMB68FHnIPBcJemm2EW4gCtEf6sdZKK5O/Ynml8w
4y06JqkpbuAno/Iz4+4E2xe5//FDFCbmazWnSHhiMAxxmZvQFHGvkUxufBpeZnnQ
3K4XtHsfQHeGZLJyO0TmKIdO3jcLdIBJ8MdLPClnRl4K1la97Gd9b6Wiljr/l5Ih
nmyf2rK8jzpgzPdIYsLeBmtNKt0vwUpxfGj4PqCID3pja8OeaunRCFaOwkc4ZCmZ
6OEqUEZ00aJqXrgYUa4z8Y1O8xETcuVaolIXJo1LxHdEZR627mGBSJnwGpxjMJpp
b6BS2GWa2cRtLmyc3EYuFi0eTLAuCdXESVEs0cJSOkq0ucB9ioiIxhEuCypPZ8Ox
Ax5jXkkhzRxRTTm0zYJhjm+0CBan6bqTP49s/n53IObmfr8Zn7vvq1kwkCirZFJh
2feDPpexYO/i17G/n/nNEBbKMK2cKEgDzZlWiFms4Pc991JGdiBQlwwvzN85hd/G
3991w4L7XyIF2BKy7aFgM1IYxyysHi4xzm9iiCAWJll3vetLrxPOR6c4vPWS0h+F
TdLIiAU2G99/ZaYrsp/HizA+H5ANmyE1dv/fhBFLEKyvl6LD/+cZyBTATqELfE8Z
pZ3RmCFuoiiORkT9aQrmV0Qhs/aceTh2BlvgzrnmXxl4XhE8zU4mFZ36M1Fq0lCD
QThfF4vRyX7nmsLyE+QYAe1W/Trrz3kJZJ9lfJF74RawpopilvaXq+CD9ZfWPKrv
LZ/lEbIyt4i7wW//a5ITSBbeh5NQ1EZUZ8ZzkAGdkvyzxwVQ1qg0d/JGvhF/uqNK
rIC7dsLX2FJEe8lSGz2mKyts0/hdib2sUnHfdwGENT4Y2KodyxszmOYrwgV2hyfp
XPPauVaR/jULE7YzN42GpkWykkD40Qzx0pTxRawNwUac+z+IpczuPYaLwxwfEMH4
w4CrrAElmCJmb3e8CJHeHNjqc+u6pVLPxLdtKALjBvhK8H+LJqhwfI8ou0BsVLrz
cB4Q8ktBy5WX3Csc9pXFJku9dJf6MDFVROmqaaF0WUTpn/7sN4LRKBuYC1gC1/9I
MtgASOOJgRzRbM7QV2vLp9UnVZai2HVhJxMZ4nbuDKOZWYScZRCsDaKqoXZZ45E/
tKma8srgCTfKQYSQ9AK0Dbv98C/77d3rN2CnHYTAv1j/eZl61LzCtoBMwnGtBz1O
Rk+BZEoOq7SPY/YxPkttaueL8xKvWDCqUSeQS474wN8Qz5Psj6ChLllVx3ruRs28
VTxYx2EI+sC3gOY1TMdxaWhDnlL/sYNvfWuNt9TxZl+1QezoNxbpqL2nVN8AlbEV
2jPk+GQJM6mo3Laqx31WBK9lCPLmkhVjBWcN1yeyqawvQr3970XI4n9jt9DTuZE7
NjzBo+bzbRXS/Cq9kDJ7TWfgqmkmJeSGEHhpGysrejlHOO2IV3/5WX3fl9MNb0K+
yOx+EojK86k4In/eaVpS9n0+wy73hseoAI3+j1OTc0iH3h/9FLI4WzneEaMMeQPl
P8J2jL8oKuoo9A7I7Ydq4O4x96ReeJ8yFKoX+6M5MtOAA/RGwbFstZm1CM1XRgmL
jKoZj3yMn76AqmkmQFck9ujFNw3l10d3+54SfVAAEIbPUBtGeilC642AOW1J7z7Q
St7PdWTCHGLBJqPhwG9DaiKVSSBJILtmGsYdyutlcxgQehd1uwSkreGG5lt9ogd8
2gMqZzpzmVoSISoEmPiUYVk7HLYlPp9jnLZdOwRutIh+JD9twK3ti9qGuN6sdLcb
DZjSGtsY4Uzx2ndkTeLeGPNa5tZ1UU0PZLyx/UBShrbpMV2YxTMVbBHmn+0+xckI
aned5wp4x1E+rXxKxjzIPPanH0QT2Ew/UpTDDJBvtCnjOTkCO/zMnEkz/7d6WV3Z
KBH1KvVb5tJgGueMlDPLKoqFDVH8Pkbf4lCDkKwnYxpBTbysXbfUKySLb3W1nYox
f2zBBbUlV3KMm+WjKef1mmy+msuWT4wF7OgXiNFOwCUKdORozZYf0/bWkYukKFkY
YX7SETFENEqTLBEwuT5SsUHQ+e//OZkP2rAyktReNl6QdfjDavQLmNV9xSXHiHmX
Jd+lU6/LOdBBFfm4RrpMo7c2WwSuhse2sqqRYDvoq8ZufblcoicRpnqqTFhd9lWA
RDVCh20nT+ON9t0p8yo7JamKre5PFL7VuM4dIrZRH6Ujfh/TKkqOOJ2+LXSHItlh
WHyiwlDSTIfpwticK1H5S+eblmHMrzLTXcy4sn0XgDpJ5I8ZBf/O/t/EEYuHhiZb
ok5Kz+BHd4ODxvrz9HNw2C1keID+uvbxgQxWd+PEz3V5EX0zztmJ1R2CPPygYrAP
rZM6caZRZs3rHJJ7xRRmnlxd+bprDwoPgzcZu/XbvKITW8YbGaJxrwY/mvb6/3IK
npTfkeA7rO2aTr/lanXP+3uiMHAkONGS1tbaBIk/dEXl0T3Qyyl1gZNT8xyfujXe
ndAXTsx8icf2C3TtBtrViWbwyx0IrzbUA3P/VqFNmQ7g8BDiuaClpJk+hGKIxxVM
qFXCVngukrASeWvZTqC9jEQSShTN717yD+f74hAA4KynB0MG5nEQ6R3Bwik8AlZE
oEWWivhE9vZR4KLtePAQgT0f7qses9GGHcLlOY2wU0sz+fQlguyGolQ6RWx6UY7l
GOr1t09NQFr7ojuoUX1CMtiRtFcMTXXfLKVQDkOTG/qhv5HxPdR7AXw0uaXNSIPt
/q2QOOsJovXMP9OS8wZeZboO2uBhtsnZNrDP9HcoS3ej0uGDR7IUDC9N+SCbbTIS
RXHVMW0ZZLg5lZ1WmY4DFVCm0IK9r4u6FcBSb80Ku2ROQWc76X0moLC8updPCShM
yaZixav38ubvQ2frGXsQvJVvWuodH8h4ZxS0M3RNG3nzojWw/5Z3yPosaaqK87Nw
L5UbxEcJRJ1KhgLcmImsU8946umUvc1SjEb+7dTJLGrdkRLeuV5ajSsvPAGBX4uS
jUIF42AeDdMQ85PebeHHOrsCpdikGgYhB3mLxqn23c7lzmxdSPcvSEJvAkK1xeE6
gkBXTEKo10AxfdqLQdk/4P1snodpVvKaYpoQLk7V+RhHLiKbxwZTbxxBNvS/Egih
wlaSYBYIX9PQbku3WExiH/RFb5Fhzy1FjMwbO+eyS69MdpyaJzCmQUGP9XSrpb/k
G5hi4i5SlllaQEOYbj9PyG+hsopJIKJIA0waXHgPPIC5mYryDVxUsDF8JOWniD2K
nktXfDCGlijlh0rUYTzTvNIruVaNWaYUtFjWQxzHxhUQo6b+zzUAkmdfZZL+oA9S
IClUTcDpTL+/Od3jKpgHVCrX7zQuhD+RkYX3olENtDglcK3QcI9fRWp8pExoPRGX
A8b5vYehs/wAPdmZ1xJH4fWJzBVkthduX+HuonKD496DHnGIXSI9ALqMmwYkcQV7
7F2aG/T9bXYwhJfiyzhjYDTIkkgDqKQ83O+0WXM7PjZFDBhe3u2PRIHFLzl+U1qp
A905xrSQIeF8XnaxzS3C+vawam5ZYFJ4YCS8sxt/aO25942OF8+CCL7pPSYtoSuJ
HyP7uhWLxiksFJMycNIP6d4uBdLnJFBDEaE6n2FlQTGRlGk5ByzFlJSwVHKA5mnn
KE7s8Btp3mxXgnanyN41u3e+pcgpp7CZi3YQ9s5BuI4on6AnQg+bdh1S62X0+onX
dmLV6101iBcfbsR2LSEg2pl9eCFIwAQZsFj5ZUqZ8pHNOrtpMwlQdjPOO7g5CrrE
yADgI9A6WQZKqUzdWOSEwuOlEn73gkHdPMOW1nU44yjB4wKZ3bgxTv3r92tVh/rO
cPW5sKs1uQHbbW5GPaHJcBEiPbgBltH/Haz2C52ck6AYi0vQJBqWTex+4s57LX9P
Y3DLNZbJlrAhAbsqmRfeZ3IHiv9hxRmoxGoReIIb61l9FB/bo5mjgSWJojy6asen
gOpQg6S8xxQ+s4pXRMWo9nQWPgyK048fJ86yv5TFZNNOw1r78wDTo7FPoMpL2BRR
f0vU0qGPCPTsgn2U4xT+McWtl+1fnIWRqVFSLWCsZWW00jY8QC912JKsCRsco+mv
pp9DgHA5hEHRvjQ5FLG+lNn4cwphf2ReM7cWngMMCS3J7UeXFT7qb4vfNqYym7bx
Msil3kKdT5CCUO6JQZ5+22JLrc41MHTwQVAbZ7u5gNpSS9VSrGLy+OOfqppDhAyu
ltVlPBH08a3JiaYDP2mHJNpyUiwkZG/L8sc5X5wCR+mR/O1DNR7pX5dPKgojBkdD
FO9uwHd5J+Tr/L3ipSFkQcPQHdsY0OQFpF0Wgwcm/+LFZiV1Y7rgIaBBOea7qcF6
247UD+GHFUi4GXMh4209/hJAJHzpT4JwJcpByc2uz0asgrIhYeXHJDZbUnLL8BSe
aCSdZ6bfl4gQPsn0upFwJCAZ2TNV55l8y0GRlbaI+HhVkD8Jz3tFtV6bIB6RhvXK
gK7vWoaOwljEhcqXwa00m8E354BBvJH0yZkFJ7NijaCQIilkK4WUx/tqQ5SOhX1F
HqazHNo/9Xb2Zu/la7y8SZBk4eUGbe59pqyAJItGpCNOgjKoxvi1S4sDfJndx1xI
Ths0uEXfM6WkIq4aGJySZkSHUmD9og+CJAfk0IDglZ48tPbGCgnwqNt4N720tBOc
0kQBXFY1er8Pzq12x6ZHP0NbBQBCtJjuZYGLBAy2hOh2Knw5SezdljiQpFdJAy+s
+OL62i/v4q+gN4BunkAh7eKE3JDiFscSQAVbGgl+XdkZ3qncumhACrh2lZRDchxC
TFSB5RROsNnGO85x3GVyuHH61edUtnpjmwUCcpRo1+t/Em4/y/vq0eULbeloD9a7
h1ei+PvTuyNUjM+o4p51efXOcL75xJrRN9uoDAtQDs+i5BnSkTFJTP5Y7tsWLvEe
veAvJtA95ZZnBC9wIOkVRk9swzGIv3kv/U+DQxMr9SfV+4XyWqR7Vo/5JpvNCpMv
BS1jrl3omXKAOeaNnLnIWYHa3F50oACb4Qqeeq/arbvpZ3dSXQFApFcQsrtWOw0T
xYiZ8j4ofoA/rK/4Z7plq37UbhanE0tMyVhQttBqEQlnruZIVJjU1z8SmWWUQrOj
pVUSi+rnHGYF4r9meokAbjgpRoxO4Lv55+4hi6vX3R1FCq0DQaoPpqU26wYhwrHC
ZZgxJAtkTfA5DoS1yxN8MVhNcbDvQxUJY8yqgklVhETCb0tfCio57yFg4xpe26ut
rbMsGNuS4PzGF/UWz0kZ6jgb9g8+6KqcyNdyGqNDlz4EYhX76Mo0w1E10xqnSc32
ztp2AtxgCKyCfptXpJDP1XHwN2aXhxzjucxX2vqxRqtsI3/GpKPrXYKBOM9797+T
rkXtG+WwL6mNcOIukBMkG0xQdaVv7S6exNsHhiKiTEO2G83nOcPHWNMO0Vu+I216
/vhLbAn4rVk/i7VUibNKaBoJ0fbKaqruzu3WG9lEgPg7/5EGwKQbHkDmTptP1KXP
MdHqsXhpoP2HChiZjAxQ6COcHwEZy850P++V8Sk7jXAkeZxrFQ12ysAVNx+hoWv6
JaeletA+IT7Hn9EjTNuLFzHw7mtsFWeNzo6+gtpRS9S9KcEKhdTn95thTp//Aekc
a1dUDMjJjyk/S39wESbw6TPS7LF59+w24ikPZbyMYJgVMq+ri3CCIFu0zdotulIn
W7QKnxreb/POiFAzW24FFy/eAM+WLqV3AT4vpUOQCBwINYg0oCwgEXITbwol3Cvr
M45iPpXM0A5ZH+THoj8LKMvKXCpWfeuvJjqIOo/VUNPt3Pra3If/5mg/ilJOcm0G
88KewBRrQGiMNsT17oDodRvVGyBTYjpQxHxcksLKmnUXMmy3TV2pq6bQtsE51Nq7
IqqpiKyzQ8tT8ZteWhnZT9cTA2ftWcsSkCe9y2/uVoJB73Xk5Fcik6tzhI34EqIB
FTHPmstZJTRfSxB5Qn/sdqiwH4g/dzpHfw9XSmMGCshhlmhCB96FEU7AuvHal64H
b615AZxt0TtHcLOcRNSH9oOcS1tv3g823g6IuRXsbqsQ/om5Yx9JUT8d4D5gkV0l
7Ku6l2c62gidhV7v/DP1m9sHJKNFTD+BmM2PgLAX72W7H6w1p7TCyp0iLiNMPnyh
D8k5nBwxsUhWmaBDRW6q6wU0Nt0quGF0RoiTSjZWgTgJkpirib7ZiwHTZeAbEOjz
VBrJjoEvjHrkCqQg16JY2ajMHwRFDJZkTTDnwEc6GKYMqs//yvkCwoBUcgu501uJ
cdZs895KWpKIvk5Z1zEo/yB4ittEUVQZAyBRnojpGIqmVjFrT2bpbfskXVY0sUxs
MepLQBo7GZI8N61/SzmJYuJGOfMriYa7YF/NpwyHHzC7MHUY99h82tmOgl6MVraY
vQHg80l3PMEL/noqJPBuDgNSTlcsvyeESU6v2IqwTVB/ucpwbv7C5nj6TbGn/hwc
ctFiKF2mC+sGfUwPaqttA9lHt+UsR/5p1sL67K4QX7htsuDIJcGuZ3g7f83sekep
o7kp2ijd97Y0FQeBHASldq9TVWw9rnAPgCGALVS/R6c/oJbe4i8F52UY/NW+OtBL
Bjbl20I8cIIRvMxKKLbb2KrZMWQhiZUzpG8UI7c3is0ptr+AsGmvSQdktCVsTSzU
lO4hhCorSIIjyObfAcunkEvwXzCdYph6pHU38qaCZOuP56RJDrhdBtAYDoSIuGII
lvO1NUu9/mY/fNpG/roJHMb/Ir31n8ghKlucfW/f/C/YPAOxyMHWUX+YapYNhyo/
8WYFXZz4+eNVKPXbRzWLVEb8k4E7C8EAue26OHJf70JRWEnTnzjueDM0e8dmEjZv
2uUQ1Vfd8qVvjJUnrw0y092IEejTHs3YIIdqH6HvoR/bZxcQjXM5twrer7z5qbgJ
fdRdNXNWQxLPlwwtR4mcs1GI3/dbarPK+3lIcnobZuUHT2YKr9NRkpVypTuBgkdB
IGNafXHn5E2zBsOZ3VhnuRoG3edlp3lmj374CzCNp0o7AzQM0OOkmCJj5S0p6wlF
9KmSluT37gZTxPUyno83sp4qXHTitdIxT+G3uIWfstzzacipah49WeXBuByUmIoU
PR6gdLhLBLJmblvD7jpMmVgWDS49Uvh8L4lwCS91xSkXUlEV6+WDDarqc6Z2mDvQ
6gqVWuWBB09njMLUcK6JUBfMYKeTc3WLIzoeJ9WjfG9TEBsp7a+xduU9CTL2pSnH
yTLhgHiTW9pKD7bdVvLkeXuB2+csSEE8KlEd6XDtL20Swmf8TQo02Zp1KLjfeMTJ
jb0L8cjusx1UahTG9cU7rSxLQyPW+cACG+2b0ApYwpm9PVYLtM+qVC3vCD187uEa
HelAiV3HU7ZO/fmqcPyVufE1s1Gk2kU9rNqad0urloLjS8WQdyGMBy9Bq2bwDK9i
xZpPBjCO5aysCAvXaoeX4Jq/1G/qyof8+VajUrqI/R4ZjIvZG5ZZMMwyeCbC/XEx
P/xaoxXWiwaGtGile+x5Cxrg0EzBFbY4DhhVr+q4VZ1xsDX5LfUDhm/uMzjCqPq+
BODTkhHSdagoJ1K1ut9iaHOut5G5CYq5ry6v7OIvSZXEgunsIGKWP7VWoWXhmxhu
ZxX9L+nBQlV/bqfdzH2Nw7LlnkpZdxZJhYlr3PzAxOqCYdjBHjBcxeT95CjDZk6k
eWmX53k6yDeoWEdvu16wCnVrftQSqEsY1iu8+vJySaoL1+pGUMBjPVIYt6j69evF
RLon2pZGcYT/UL8QW2Q+N2RPJHb6wzxJAB8nitR1YIl6r2BkUDUflY3REWKDGCpk
23MzcoZNbKghRd3stx/6VnKD6MzUBsSMcWD/4frIkB26MBRY2e7fSufdefViNERd
6YMBexAHwAljbxD/HcAcyEd3hugfC39paMPrkRu2MPxtGx32ffmxc97lSpayXKQX
k3+a7KmHpElxw7eZc7k/nRxbrpPjBpl65PUA52xKDhzyx7PppKrJZoXd0BaIUolm
4xh1xpSkI9OQ+FvkJ81vUAto/9NFuMTQmWcN0geLMvhdX1MZLeL3Vm6HQY4voxGq
n2WDkaJt5L+MCcmbxsjhA/7zmexNQnHtzM0dms20RLm0Tk0WY7ltXYjycLutKNnH
oZWPY1tB4tgR0QO5PkZYhmUft4XVy36xFJKX9czM48n3ERL/mxP70zv5PgauLETM
jBrCotwIyUJk9u/69Z2smwu9DCaBBT3jgtgoqR/We1W+o9AVm8YQM75nl0ywDQdC
zfjSU2hFv3lQcYgoDJAHSsdeeAex6CEc5KbCzbIiKDTR0EFVNssoufv2kWochc95
L3Wacn+9hK+cq2v69koe26QnZkP2v0JcWR0Mgm+ggEKVO5vgBS07u+ydYQcaCIse
VdrH5Aty97WUdoSLaXiddXN2phcXP9d9AvuQjAzKrxayciReUnBu3kZINbHCn0kb
Xp6yX+R1CrASCLOg6rcQiU6wlq1wkVn6hqk54hr1lrgeO68CtfTvJ5qVEW75h1D3
d1Efg0x4gsIW2JGkjI+zBfqgNuULD+v2KUNawBAjfENfDPrD9fEsJXIiTjeb5XAM
AEsm1bB30GTudTQu6/yosav50NGyae+dtCNoNAMzxpWqRzbKdwIkRtcsYGlVv7a9
0UmkjMeDITJg+coZsxKR6NaKdL2eUj+hbTo+ZtFlFPTBcYlm9JQZn/Meo+Aevs5i
akh0G5L1wANeZu48YwxH0xIkX6n8AiTwWHAYOuwvpuvaS7VWofiMquPXzU0J7sS4
RLnZnQlp024DtlyBE8QKvmPc9BmendXDJb7pPYdE5Jjc7PdmsVi2a92iAcb90eS7
Rjzggh6h+tQfgn1+THJlbNJWpAVFamJaABDlZWWuRcvM2fsftnYpR9Hc3N1HqbVv
HKYlRkxw7g40bC11I4TrStxBxPAS8d4gEqXRxUyuECWQF5/okfT0qSV6mYqLjA3k
WQtRvpv3wkRkDYr0bYklI+X9ixjZfH6QTzZHKOqUQvkiBW+247Rky0X3EfDFsKzK
DBQXx37ci1AdOPHRQWt/3+LOibk3PGUXRTbjXX3QTMpRH5NN0/VSPMqO2NNLu6nI
1CH8iJxFIFy790vW9niE3r9Atg1mRs9BdvCiBEB4ix5sEDQYw3b+udwosdav6oj9
oiFq+uNIIvIDUv74w/WxGdip/tL3Eu+u2+UmK8I22N4/ZaKKkGbadRZfZeq2W3CK
843EJ68O3FQeXZQ3+1roWIFASx2qraNoiTP9Fe8DXOEwlJ5v3baqHxrZz3DPtRTQ
W698WgFMb9NNukXKbgCNERYH0DHvPEIaHbP9/CH74gcjWxrO+Cm1Z6WN2wuuPK5u
+W3dn171qIwdwiLxH0KO8L0yZs+tpyWby7qRkVABa5/p4LefRtu2AVHxdEOUj/bH
`protect end_protected