`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2128 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
JoTcvogRvquVnxbhrbrkfKF/5gNYqZ7VkRA/f/A8iQU3QpAcnRr4MOfABtrUjPTs
7KCsSTUSsZ1rNW19VN7vDWCwC6bRG7SFZAG9lqqHpKLloh7BWV0tnyw6vlQOEfmm
5MRLbsxN0L/RuPEqhfVfC6+ztImtyleHY5QZw9ZD5old7DQbevxCnNViRmSQ6Lie
mmEThkPOm+XF+ZBwTDFadOw6yY2ZB/CoBKzI2s5tVX7BnklVrDu9a5sdfHF9QuEK
dGKUU/Y57E9yigpph0Rn2gYDXz8tj6GCnn7D1/guJFRefl4O/ipYke1nHG6+G6Vt
uMAZqty6O7ujdfZiSG7mmC+CGNcs1jUZriZ63yizgHgaR20MGJ5Zu80idUbrIReY
5jTqmqkMoPhx/A2eTebRoNzoeLDsCXPTs/dCJvvKEZ+YW4YyXDqY1yHe76CNlYcm
Ql53ayC8DC1/35vYHpfyCQrEgJte1xPwh5rO8R6bEuAWWI73TFtMFZNAqaHNtgNU
AdKrOwltPV2R8Bl8oyDn+1caAY6qFx9CYiRLNujbnJ7LzF92nRL4vHmB9A8P0+W8
43vdPfb4NvdLdd3sR9EafH068yqmjDwUOltesalKeg+8CLYHkzcwAq72VIaG50vb
0i29hHJhqkVryGsiR2HMbMM0qlBLI74YpyFd1H5AtOF95eQewI+lPcIu0YugWVKW
0RgsMG2SsWYEL0NXs4mi4FP4hw+5woJ5uCMooiNaieFVMHrOTd7fuClht2+veqlR
TjzCtW8w/3ehxer7u2gCeLhx7DsdJrtz8LGPds3GvojH1/OSgor+E8KXp0fD3vNj
Mo2O7PsLUCPePNhj8YEmie2Pd7Hb02X1JlKRPkPz32Ua8icB3owuuHUIfUOMCxF8
rLT37lUXT9kabKQLTnj8ch87GpkkFEg7FMX5iupvncmUIfOKFAX+jOvC4ico9Tif
9gRmIaye3q4qqZw8AMA9oKgPmAabGVC1eXKAtrbipnIFMYseo4+Pb3Agg38cY/FZ
8urH4fiyt3aHiB8fxGymnu4nUsLnD4XdBVbXvC0qhVLukrpkLGLRPRB9VpMuplQh
B3N8+1lABa/R35bKZCaa5af0Tx/wyxJWDWNMLtM0YOaYtJGhFJq1qO94D2BG8rrB
Oa7qwA9yF7Bz6i7443RDIdUjq7WbviIL+7LhW9IZHG3t8VttlQl3+RqJ6obFYh5e
Mulp+TVnMVkdjOtCARHo67hH2o1vGYNI6lALHCyluzjBC9QIP5hKfQKyZSJ58q5W
7BgN1hK+VSX7Gc4DsHx6+DA6vgX43DpSRGeca9KTY1kAnTUXgRR3GqjUn0AdXziI
tpCfB94JHS+fuaqOiTjO/ub68aKn0FL6eRopDC4fnAgbdGsoOCJgvjyMNNODpnxU
HnXe+765uayKumv+zOsy3TkV4yXngFkvXKfZBq0l3AVwSO7rcL/H2PRrUAyUqAgN
EqY/2l1HtZh+a1bKTt5iRHOO3yLSIWNDtBaRpJy6J9ePOwZTIx9vRqQvc2En1M2r
nrE6IhgJLdIVhZgUb/TTYbEY95CkNs/ai7REM/8oniysffEMNrKJctAXPZCwmysQ
NEJZzcjVeaIGyn0MNLL/IvFYCEjBCjxHbWNlDhY2OR8EjJqs1XzmAfeUfBCI91Gb
nx22uxpGxv71qL686JmzMIsQvHAM8a/GPJTqPYrIkgE6MsJELuDE46TKyRTRd+WK
S8pSRxxPl6fSDIwgpRNnozytNB3eMJWochYyzQfPHS2/d+9J2PhWWjvW3k/RO1jr
P+O3D0Wfbdhr86Zz2uB1jc2RdiVtxCWtUFFNykGLPT41D9ccx95sTda73N0BWuHt
HOv+NIBxT6+JqvHAxmVreoY7vwosQ97iX0Zlt0oz7tln6jNTTW4frtSgrjPPba7q
gPUyNV9qbI9h22SalSOl3kejFTJIJH/fRcLyPrukdu8Ab9O5RMA1umB4Asg80jK7
1IJuxFZUmgcoCtp5mpiC6r8sU/dr4nmCnLt2v1x1D2NPfy9OVpyjYfPn6tBzHZ7b
FyDhM0vdK4C+tJvpjC5v+m6kG5rPpEwLRr6pIp5ldKH6OZehnI3bxgknKiPrnifZ
p4V81EhUvYdOAngaih1CD1rqwoL2ig1Y5UwEBjJ/hU07pHc9aGeOwtZlr7OX08fb
fwvGtA734dQis4w9I7VufaBCkzswEH8zuIJN6WzGw0jEfHxTVjk/tjW3cJAw7EwI
4uK0Naw72VeZlQzFMS/wE/6y0r0LeybGD3vc49PY3Aubabw6XGyPmmGq/b87zbCf
m3h+UoG03CM3NAHxO7sYfDXsBcBdvf/Rj9ceAcOhh1jJ3iSlTF77E5XEN7Y3AEnV
NZNk6I9h/pF95aMmaZucv+BGGuX9SVxah8JV6kr28um/cH4Xj/6B0+Duu1cXzDay
7sUvbgNRkJdJ64TvAOM+s8p42bjZkcfDZVWqzUqEB5YJlg/u0DmZQmUyPzRtvOKd
8IvM5ceVJjqo2fid3SnSLOroWVx0Fnjc9qeybnjM0CYj2cb99cvFZNKkpZ38uLC0
fu3NSawLpZ1Pl3pyQk5kEDL9+Zdfpzcf8lRibhpqndWI0kny299605sa9HYJAZ94
hTkZOLm4zI83QERrEVLN7H13lasSz+YiK2s7rXbMQ6XtEBvW0iK9cPGDnPzpcfid
n7OFdBRBuyqpfAXroVWGeg==
`protect end_protected