`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 43504 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
5ak8DVq41YiTdsbEXvarNyT9AsKyBCu2roejenrWhs7GAldWBMvm2SF5X66m/5ud
LWG4H0Hch/6PMKxjoMYp/8VDFrVkZwQNm5v4RazZoFvZdavfVNcud7utWB7fBhkZ
AB+PHesjXhS0tElW5t3OERnkvHhWe7pWPzQKQvs249SB5dKeFH3NWAFWLcQaIE9V
4f8z5yuENQAeZeb1xRJCH05SZdFWeN2YQ7Dvg/aMExSe+IkzQQrKciIa/ZyVXfUc
owaWZw2gz/gwvJ47eitxGSHCt9ZAeq2x1mMalg3HHXj885+B/R0zXYjcqpRaNU9g
hHkNPvdV2idubCQZsBBn4r1Xu23C9FT8Q7Wu79IkrlqW1MooAH6UK8RmnWNflUy3
1yT3IgRUQwNFQfVnq1KLAEvPlbKr0mddbcR3lVJ0pyecIes3xQYYTdjAzi2t1eeh
l2IdeVSLjlWLUUd27Sfa8eska+LJ61LT5phhykVoG6fU87vciM0aiuBJT0B4bFDS
TiAiQjyLNoJ0om4DzDpEG4pOPZjnCnWiWYOSB5YgiRsencDsJwaaYhv9tDGmjyR3
dh2cRKTNsdAyNyWx27wtWI1LT5mXr33Z/1ahed6JvuiVZqhTN3TkQbv95cNNsHe5
cuQOvUKiSyE2rwSYoHMxqjopiZLDE1W8H46JZy82XezFZqokVVUOf6n4lYFSu2Yt
Gmg2nf9Ad+yOKC3eKkr1mlDpVJi9QxGRYL+TAng6RK+aYFxBRL1mgpFI2mLzZHeJ
zqB7QC3nfUp6vqZnUKobOFo8y6WI6P49FeqJHD/nIQUvpAbdhqcCXp9MlgxDcmIu
3kpVnfwEfGejlVG9gxVIi5Ta5Iuw7b0EW/2bv0LzGgEspD0jOmEdp7QsD7PGByE4
N8hO+ut/XoSyroH3+SM/ndGCcAyae/YllHMOEteqqp9bH3eyGKxhlmjzsiafu1gh
/CwNPBKBJlIo5LEU6ieNDsZpZJpRBzlIlu3jBDXPbDnQxJlDMb1L0icBtKBaXa4d
JrIBp8h43kP+JvXPSb8ZNA26pTFN36/oeYaKLn+no20MKYr5Ynmv5THoL2qnonx5
uCzejyPG9fXaNud6wKX3JJ4EC77WUMxk5wblTlA0Q954nSJ22mAJPQmqSrK7TjdT
HlZvAkxvrENpLIW6kjvY1Nm3FIKxBrBBIv7+8yB5h/5T+8k85SNPDv9oHF24aNwR
ELQi58M3nzPI4if0e/kdKki+2v1TkkAbQKiEvAra75diAjjAEtvqT6VLr9HxiR+p
IUkQAlooevy1EtrRh2ewq8HjAuvrIL3xj3Leg1YZnDZQ3DiyM9cvO+wquq+Vop12
IgAcZJ5wSIhtxZQWEEuBBzZ3PNGfovVG3/fRaQy2xXhgulcp46hQirqarFrdV8vw
oAVD5W5y3pAnUfHJzfylfObnLtAL0ORdILb9OEC5hWYvIYeuKZxRK97sIrCCKx0I
bxkIj7nCWG0vOtoKlTpPLCgUs+uXDJw0SP3Jne3ltEhi09mrJK91BgQvGLPmCCev
5nWk8d3dWUc94ZbYEAMEj85RoebAq8S6q0VeGd4jVBJT10kFDn3iOdxdB679E51b
LrerRfH/likaj9AXogjZn2sFGTUZ7Vqu8nSHIaA1dJ7M5LkHPwRegK7osxccDhRN
BkctIO7XoQQISb1J3ja6XRXA3fLoHzfxnDp4OmHpZgupf7NrNi8eHwPNtstc2DJ2
ptL2TPMOOtFREVOf6DLSjV48Y1JEuUugm2Da+wXEk8XohTkeleZ0BuvMt8i79yXo
YbvV+h8gDOicX4xXLwmzwrspy6xxL8mvmZV/byBUFh73Cs4zT6XQZXHv7HVFWNFM
q6VOOvpaISp8n5+Z7SU316P8zjFOA8aZg6UHy6Z4NfXWmfHzE+OIiuiL57TT/PTx
/KDikoP+vqDvDypmZzX610HDOt31Jktls8jvf0tfW7YQQ7bW6/3mXmaMYjrUVLTl
3hGmoIJFJWEjQSgDHrafahOv1AnFVs7vTIy0WWhmbnpS3DjRRoGauOyVTVVSG/tf
atrDeHisp4LRpo1Du/5I+CkgxhLCO3P9+M0ZyD6VtKROJOAQgbFLdmOVfsfqAEUp
2ze+9jJHoyVuooKyflabNCk6lGwVL/mbXhl51n3l215lK7EIAGaPndJLkVixVJQT
/ZHpuWje4tdf+w2Z042oHsl6GBHkFjY2U+855rYMhzJuatoW47c98ZVyGqtDme4x
pULdk5590an/ocXH2xFvr+7rQJuxboPCz7Y3PFaax1M6tJ0Ht2h54NG993yNYH2y
Re7DMJ45hDqkj6KizwdyXJpQ5v9+uyaqVUb4nm33ioSRkaBB9QjiFlTWYSCHrhTJ
qyiqpoS7i0ryRjKtPz2EvoCVfwxQjc+Iw+GDpCOS6fdOLY744RKMpPI3LzBl0E20
hVxmwwaCVjhk8exifb+/auz1mVwFppbiw5SG+GO4HrdN20HUD9inQO18UGKCVeTE
H1WB/u4/p8iA6k2VEqnQ4f9P8uiXYw5PBKz/ojMOX/5/v5UGYA2mchih9W8do4uo
EgWt8fZCWIuXPmc98Utgzhbw/jauGid5Ugp9z0uPLu4qGi51GguF37dYx8Sznvn8
LzRiXVubAa69AbdY1g1HFFAjEHYlD79z36AGYnyaAyf47SQV+M2K9LJBTne8xz96
hDKKh/IkemotQGZCTFjowA4lKhwm5eUCF3ntP00ZbSjTOU2dPouRNhAtMIpO6tnx
D47plXWh4i1aKUpPHwBDOo1J3RtMtLXfsAa77ziHlDQEZi4A7kOv4ChIIOm0Jrew
X93imDVf4svSD63g2mt8ZZ8lMlhINF3ifrBbyJpIikxSB/2irZNiV5Qsg7OxrX+E
Ef7TpF5ewQ/NlXWkehfl3yxjaHQ7CZCozpXLe0r0+1f/zK/6Cs/dDYfDAFqIO/VM
cx34J8ktEbqhLeErpOSFPPYpOTAq6ug/eYfjDDOVKnJfrnqd3yP3ZGzvHtZzKrKU
Jf1rUI7zar4IdrmKs09JVUFrmo7XU6nDbZYZXd1xOIrUcDYqo7Av3eaYSEuyDtoB
Exs5/+k9IxqIjDipbK/h37olcP2997ngO1j9zovZllcit8+Wf2w+qrxT4HWm1/GQ
dTff8jJWrkzPdPaR8v1wk/+mX9BPgvvStpD/3arL0Rt0u4evyZxubOIKIq7Y5Fi5
vTyskIiondOcHkEKAr5u+IoAPIA+AkpLgJEeZpUEnxxXuFB7mgAX9vg8cQGPjVEK
Zr4436WR7Mxheg8/VkNFodOLmjzZRa5rV77u5XsoOE1j+XdBJgGvy98o5F9vrABS
3mts/i29yU4oBdpG1KW3BMeA9Drv94R+isTtYqM4oH41MAw/5m5aup0sW0Xq5hbn
47y8rFfApA7sfUvIB9Gl43p9YRGIsKRuWLFAaInSwV0mcxbxn/MWwctecnzx3rtj
IuSN3lVliuIbnbSMPqN0meZWQ2mfjF6KrR2n3h5TOGhOIk/jiMKNVB3+/0vUN00g
U/epfS+ynBgPfnwBRJ0FVhc/fY0cdtmTh9CMsKvaFUgZOMMIO4Mb5AZUptNyJGGh
oFTpLkWnpD96XQ6eKY5uT8f7whoySffQE8kMeILDdkbALVWcjN8Ow+w+N4ODE0BE
NLeLWTORAJ2ptA/z0n/dySPbhjjWh73DM9OmKVwCH+vVR3HKvpmz34X2SBpQXG5W
gt7AN+lqiONRHzhoRVM89BqE/V7V3Lg42A+X0BhwuSHtvcaLvhdEX7OawQAFK9Cy
7KTqqPPhnPkp19T6k40D2j3IGRQ5if+cFyGYwCCrRQ4KAW43EcCBuu1E9mLLdCGl
S2olf4ZAKCRw5TeAtNk+tg6t/MGQ//8Suv81zqiECTWJn80RSxeIWcGA4GFKgseq
FQ6iGA7up1F7KGBorbgYIfmjXgvraPSljsax2aebm7yzlD6Zcrx8NYALiDbnudIH
X/LrFZ+b+TYfYxLMFTmyGn1pIWFU7BkPQh8IlpnaNNOPXdjixseYo5JYY1xsV1O/
71kj6YqlT61tcHubtRxA5A/aiORlPX6h4gm+EVfATCBu/to/yKyP/U3wC1dc/ygl
Uk7UWliKAM25e18ssrJbZMt/pPu/53wsH2MaxEZPInUoxsVlMht8oyMgctxwEeoL
yXWy4AfQ4cK+vtHFhk7g1WIXptDY5wV3ELCYYuVrzZmm+70RVACguOYL55f5YAg0
q4ivTUFHt16WtX3aBQ+4s+5q/PMyi48aAnSaoeT7rSHj+os2Z8RP6KzeDpRkxKeJ
diBLkLufl9SjO/yaCyUFqDAYmblAb3QBYLC6p3vpgClTsG+Er+I764oYpd+eEme5
hwMwdOeK6sOlBR5tPH9MbTUljv9sjqfdvLgmat1bR3bO0OTV49gqpTA0b3ABr+jA
FJb1zQhyG7PyR1GdZamaM2IrCPBWhlPj8acQjcRLyFDYto/Cadbr/PK/c8HmKz39
x1DqttAtJXXV2jJJXouuiXmbW+hgrzakbxPxYfi27f42cOjDe+lTU+NBP07zQ8KI
6VfIHgDGfy5RWW/7NK/LSxXt0DrMe04FfBWneM7V1qVDvPKHqfdzNiDpazWV2OIr
3PUfvuiXhq73gWR3Q+oSq+bzgL4yrybJehxQP6YwtsxehBBIcc/lkJo4iFdRxTDW
3bx6aIEj09rS05RvVO+Eop99OZ4YdeWCkPl7q7mvLi0121xjyyrh6BZBd3JK3Xi6
3tCsxicu7YLaDlupsgdFTu0N27ENwhDRE0/cm6x2al9i2nbLO3HqxgwZpULw2fu8
hM48vt883q+MZV8hDoU7xnWFnOLj0Naly1Wu8IIttpWbY0kTWnob5rA4nc25Za8g
134qzaQLTQ9SKV8GlyTG6G1xi3xMY45Oko2hXJKGZyARFUARs6iRpq4DRdr6bw/s
Rud1EOW0dcyP1Zobl5+GdwN8jKZAYtazhgNXS3q+5dTCpO1QQIgPPrrfLHFtzfFO
mVpIJuZqz+5R/AEivIYvq2mgpjVQEc4X3QA8q34ux5izOIZR7HyuK2+gF0GND7Ih
W6yRWGTstY31nIC+GMhO0hyRTlsPh65qgUarcp2kr5GhkhC6RVLT/q0UeD/btHdK
Kkx2B3wfq3B2cYZIpWy5zxBp6/jrjjXKPpP6xJfhXaP94/vGEAnVmfKwuUy+sTmM
aRmJELf4K7xvebeXNyY6AO0DVixZoIYQlMAUZ6WlYR2gmjIh7KnCWri9Ptk6HFi0
OOhsJyJncMxu2Z79qjX1bfq1901quAb/RjCPd29TZL+lVWABmy/rMSis1E+4ZAVO
UJi/cHRhEhWBO+HUZ9BGLjJ1gK7fAP7nWvASK4+6noiNQrmTk8Vc8YnSCHc90uzC
mcKM1RmukVv8vBK8L2mvxanNLs1SQ4D6R2wguBG3ZPsBGXaS6uL1MLhIV8U2RY5F
8Ok9dXNvnD0Kz7NtLcTNG/lkFC1cu0tSuJg82+X/spsURxjdvgSLcyXXi81J5jh3
jjRfSg1XnCif6NKKL7rcUkxRWboguqeJ/iyoTAWoO28QQz0kidw33ph4xUEM0AsI
GH0Fa9pPf9Uy0CQb3RRiSTCTdE2E13RD1z2QnAz4coMy+/FTSPaD2cNoMySq5ULl
T7MCH1eCenQ/kK3M/MyLbnuKIPuujfkqQwB9K2aIMgZWjLhbFMlDxFS7mTOHUmQ2
ndhUrQFFmoZltIS0ccg6NHB54MTI9D+tPnmrtU9NBKkyNYWJJFroFZu4RqEMoT+1
YapjFkGe0F7HY26+ufSEaOuw6WYoW+02b8XLCHEmwgf9EojqTyooQdE8S81YW06V
6uC7zkzYoYNCfax1o9SipG3UuPptA7k6/xemhmEoRbZQIe9qMZw6rVfjTxaQ0X3N
nNEJlyQP7QJoA5QfZ4NOS9z9puDpvJlC1jlhDO2KjeX5zwZ/wuSlWEa4DIzgqmgh
4a22WJJS8BdPgSCa39kVpqbEtLT92VyGbgKgEa8KzDeO3dZXLUu8csLzWmYxJzfw
c4FSf/TncJw0xFqlHZYmK/hBf9yPwc1+GeTHeYOWZwiRhonRWBjca0EV5bNvnWkd
GxaVU2jm6e772AA4pxwrYvSeQHSC9IhVaGH1JTZ2hhZukmSl/SuvnSw38wt/Z+L3
Usb9fAnvx/9P02kYfw3AvG+lZqrVf9WdMQ/qFzQP4RsPWDpkFxeFdG0X0etdGsqr
syN4tfDhMgJ3Rzjg86coUqn29CXU8z3z5jlGYCRWRSs7MLPUy69lhxEGiuVeabsx
M0Fl8xiPlY7xmbt1Qzki6eK+hn+PA/TmnT0JGsLxqrF98LoOsJfjw43beseBocXJ
s51gMQw/W24qPwfszG1n8oq7V7KCTNlZhzWJtbVA92APIsZ649bogsRnah8UpQH1
4Fhow7r904XL+a4BtLRqhSPf10fgaXtC4cmDxHPCPqQ47tAAINxiRNvP7/gcV8+h
++qd56wjMXUq6gIT6MdCGvAXaiTUZsQKkkkfxkSKSule6/Zonx6C5BmrNSjrx0sc
PER/odPz2aDZhsSrhMDDbsv87aHjl3/481WioVsYqh4gCR3S7ANAFYOGWfol3jc9
7mlbcUFCxnzLYl8r5sLNI+B9dFhTli2n5/ScDiWZEwKWKpxcdpoc/yOFJh4Rr2K/
o9XridyGDeSlbex8ZgQoX17TylEwaluc2lDJo9tz0i4+qbDiqBrtIFjS2QHmCf34
Ppwir13K7+EkwfO/iI997cmwooyA2j+t9l8NZXQbTK88radLD40+oc3NL/Gy+0Sw
ii2p01MAU7IgDsPEE53T5lvjNTxQdPVyWZ6cFHT67xzUYzhimX0johQ/LHpwplAl
/kY8jUb2lZFMzbLDiO2/asX7+cLNPFXO8NTUP1LEUIqFfrHbVOmg7790cgC7wS1A
1RBR9F3XOOJDO09VIdyALYKHlIZ+84++t7bE7+0t5L2yrlJBpQNtXzb4tWHiEbpK
BGMTlDPInIOE9NfXx8EsU7RuqkUtQkDbZn4hZ3KTkGkQa+peyWXSnLiukNfIjcGU
TeoSuQo+EdqVCFuvMloYhP2t2D55UUawWIe8qYsonXdU25dAn+1UVCTDwRwO3M6S
UOp8zEXO2KCvFXUbNe+PIJD3ZkqCUt8rVUpKMy+pxo9m5SE98+EPtRoJXP5SqREA
G3tybd+UTKK23ya2QWr5yocts+914KF5UI/97DrIy7BvrcipkPr2PUw7hGanIHFI
jTxxQReaySoekSd7wvhO6IuCAp87pFmOfTx9gPJUV67CoqUh1VqB3178R8//E0yw
GzP0aV2Hah7cbH62xmkaXxd9gSGg6sTo1eV6V5GTdQjiT0YfSXoRAwH2wA8R5hYB
3Ds8Npe784mcqFPxj0YOYfXVBcAEFsW1rXVgMa+zzTo+Qj2Rx0siOS5mIbfZsIqU
Uz/4//M3gOwrsqn3P/6uJXzIkvZXGqKwuLMcpWt48pAa7Os9S1/hQIYmakqGXcHx
RUiAm0EmR1c6RMmcbZ2JnnpxlokedK1z07/kAlCa1ZuMKaANwUXJ6IVMmjNidK8+
4jImokYSkeiUZOOappF/Ublr4se3MQxsfTDk6Becv5m8GszEqHaGRmkzX7eteWxq
Qdj5+pKrOKUhC3UG4x28+xwAXg2VzDjVN7fGO0O+DT8CqFF/L4MXgAE0wam6RmPK
YBvRNWNLiSo1oGfQ6V2sUGVc23csepF027ggx8jMvnGKr1mHkv38XWrlVNxofwWn
h0XdsiIEMc0d/3SBGDxK3/nMzK6UudADOUat39JcXaN1P2K7bEJEZ+Oj8TlaQyt+
3cbhooyZu97u/NtgAdEmc7VNZfCPhXDlFgXvwEIWDER+jVNXFbhTioL/f52yFWXM
evBCUS5NZ3Qfu3UgrFpuHF3k+ZLI+43+Ektxv8WaHRxSsuqIhjbOSzN1X+LkKKoN
RHJO6WHi0CcrWJQGxzxIVN6WOdzZ4x8chhHeIDCZMrCqw+feBO5iGrwy19yXVvnG
ZhnbsTrAaIgV4hfD/MBkv+VgLxP14mjHjukPFeMvR+4HKr7Ec90b6+DV2zvaginI
p1GfkcOadrlD05ZmClysBG71P98ybk3X2qc2g+IIuTMXDnE53bZYtv+f60NVWVoO
8XxuaZfKGwgWG5dOfqZCqfM+ap1NL3LHpT7PW0xaWxXTWeYST/brUXyeAzRpysBS
GDdHIt5Wc+Ay9txulYZksMCA3QwD+Jl2QC3L1Bqsqra3hqMVSh8Stu5OhddQ2MrS
H+izBzheb/3D0Ge2FigCE1rWxZvSE3+zO7uRAsw7fXfIFDgE+CGz/lEmPHkXd7j5
PCxABIObkOwF53eq7n9lDoLi4ktbaSwurpYhSNSQ5LjVAuJHK3IlMz6RZdHsyMAw
DEu4b3kaFPjr1IroDvqHhVv6AQnJLUVT1SRDvT1blzy8/vAhI9WthMetIvykHcgx
x4iWDxrIhda6svGLTK1pKwrT8tqa0WvuKj7hSncgMz7+FsL9kB5884hUsEyHQ3wZ
0lqF3n4AhydAw+AFRPs6sjcmzYIMNwbth2ePwQgjHXke6oB8GwtpZbAfr9SweoDm
+oIhANvUV2aaqj0s91cMvc87jDKbhyBcWaJARpRiPq+bt7X5tagrYbOH8iUW3IvY
dOg+/Lc+9Kq6dvdcpJhWG9uwx2eh8ALyGSlbIRNEL2AbHKvHpRdmr4fhQ86JmSJD
ZIe+bt3st4dJ/dxYTVe92xtob72hNTJ/m+0Szq8y2rkSEGz6fXTC5DQvrY5Z/rlL
Ydbq4TjuqmVhg2EKilWAFer2j8+hlf5aF7mrusaJ83kI+yselqKhVw+Vg1pRrj73
yX0aZQJjuoQFlX8rHNnQssXspDRrN/TyLLPlDDNR17T4cpnc3mq5hmYS94BckTsM
3VOkRlZSVHN1q1qgw125TUd0orvJQiERSerZaBhhwIOiSa38ZHzw+Y4gnWNki/40
BONLdwWwT3rxM4XAlcYIeQ7dsIisfjc+zgERLj8Z0LrFIYLJVhcr7T/Obv32WPrR
3qvhaywort7oa8D3wDft2QKuWiKq2dNOceBeVkX1YQOCNm2HHZvp0JzFEWFb4KqT
YHvfIyu5aUFGiwe6UsgO5p1T4vT7B96V5ex0hIjba7Q2+3/oGaWkiG9JfZKKtQfq
f85ys36wJCxwBF8yszC3In+8z7kf1l+mB9E3cqVrmTnT/thAZxeG8j6sMh+ntMh8
Mug0ZN1miLzHiPd5cTV9oTpk9ukId3hcVJmP4ULeedA6w6ULP9Sx9dOgPnqQKh9j
yNmQVwD8f6/UDxbV+PuBI7CfD9jtfWL1OAwtmO1q8rfx3UO/yWtCXykJUq9+SIYD
fK2nlxlqx7p7hx95pn2prD2XmAqbQWGIeGgF0MtO54a7vo6vYHbEUZv5SBmPhrEh
mB9niAL6M7iMkdJcGnhs9PHU8by4q7VIlGlf+qlZUO5P6g3jxcciWILj7Wa7letG
ruxZwuWHVmkj7LNYzq2VVJTTAcnCOQlCY3HQIy315NvvYPMmHt7qkN+iMm5McIAD
s1WnClEtiKTigYndaaOaHS3jBCrl1lPCw3ua26JE0X0WTyxjvHbRFT219nNN5BS0
u8mRE9rvzdUJxSfP7Abkuog09baVZqURwY3KDDpNGrW35GqvL/i+bn+Dkc87gQ6x
p7riZH97JaYkaij1GVA7q65W4mc7/kXwuY+Du3TziaflGOGNOSnUYoSWghIK5Fbs
xU3ympzKuRZhmsz2/ESKy5/6BSE2X3HHKJKZ7BZT8g8Dx9DXtEfduvdi0g/JhnxZ
e+vKT3/ZFSf0O2or7tUW+SbWM4c3/WIzUzGj6LaRalu0AzlT7qrb70+Xhjhnt7vE
oKXs2vAex7d90S0AyZSkyc+k23VtOk+p23MJP68Dv3iX147xP8aHkt7J0MKsF47N
PO6vJSsZOZgrRMdqwmdNVPzeyRlzl2gY6DWJki3G5o1aY7i4aCC9pbs42y439Lip
jNUomyOt7bC8/DjGfZWSUV1SM8rPkHcZnBCvwTBp+ofJIyVeQzMd2952/iVb2orP
mGVMTf7TMVVlUXcXUdn+FRk+o5U9fRXBWjmlOdnAjIZoLnShNMeIgRipTuKA0dVV
yNELlWaSh2nedieMtehf/SD4U4RypK6yUJwg5igKAg/HKcHmc2W4ZImpSehlC+/l
oy8BKEAVpRruZ7VyHJ673eyvuML03XwP7R6RW1Fxl6bdOom6BzjYe0qs68hfzNTU
4Xc3OZaKfAPmLqxNhQdsAIsu+EPCOUoqzGR7m9dTZgUK0tp4b7oQzU5qz1tVXFdj
jSBce6pqGBm4CuOkIipJIf3XAnJ3Q7S6YKFpLXlgYG62E0AgRZRCY5cFv+GCbycS
F8m+m/cQ5HIXSfMv7XqSDk/v5owOGIZAGVLFMc1Tc/YIL0WKOtAq+lLc7FXotHv+
FVlPSwvXoXSe2JtoUS3wRxkxQxtg1zGdA+Z1S9Qe7PdZEFK3qUjs7BLypetaQM/V
S3ZbzNpaGfvmaRda9CMsdwwUEOESFStzMeCORZTbT0eWDBm+e0qhqL8z7UioTC65
ByWXh15acXMq/rUlLkWMICI+65T62zn8A3pUo4xMi/g+GtaDXr/qTo0wQWToEcGh
CKK4RF8BOyEkLNUUpw0JaXDMmr8k/qH5a+ehEFbc8JvA6eIgmh7zOglwffzAjP7k
U5Sd/04WOmr2GE4UE7A8F76i0P0VKw6TawW4r+d1T0wz55OqVIXc3lQm9nSW5HlV
NZXgwEuBpd4IkBSvo7h8oU+o8cDyeoSQ5J1Q9jj8k6PRYRqPpx9YC5UepB35dVNG
GsqN0DYFequRjI9Xc2P6Nqp+/ma4XaWx4QK+Lgv9IJlhS7P5SnNay/G/gqgV0/0B
Wa/Qwa41Xzwj23yqIWvSt61Q5F5pRA+ChL2hSuX4ZBd4cpslD2ULpUQj3vxXteRS
FGy0Xsi+3O22dVp27uAoqkC6N85+7BjSrCkfLaNJ8GcGfT5cLuPl/9Kl5n+u7Y6I
Rl1kqOjWyfYD6nQz4XZFdpmQ1lnPuhE1KaL5nrluFFwPlb4a1S/u1yrQMXAfqIq5
jT7ShuYgD5I2P9q6tKcnyoy+8de4GFCeyDXkajVBN0rprEoe+0f09Jd9E/pNM2Yg
WsU5XXhUznqCSYAKkyXJ3T5KPgT9tkAJghy7mUUsX9FBkDOdaO1sUIZZSbTsOs33
DaZSxX56KMNV7mhF+rux1J9FfyCByRib8BpXlI/ctLQ/4LJcOao+JEhxL2xAAljG
nQQAzFHg/JdEwzht7/6oWIlFYjkOi/Qnz3WHQ/5ZozTltTxzalsd/6hrexvdcWBd
cMIWSHJbfqxrEYfrA6XQx4Ogjn1tAJb4N28dXiPGtSIAFQLDD60IVsI9XVdKZGCI
sxpCNe1pD1B/fGF8XGp+yOYHa/kYAgiFKSbtNNMWfribpgXP7mp5ZQrSs75Rjtiu
8kOp2Q7olD3eihst+7dS5r9VmD6QZ7mTnKQCOQtSBzvrq+x0WVxIFy1BSM0K/pVl
cQCgwasBtv2XP8pSvR2CIxZVVvuZUeT7RgHN9vRXbhWfaAr/tKa27y3ZrJmJw6s4
DL1jcOTpoLCRmhE8DnnvlfQ9buM5ZDQfPUTd7wuH2jh0hux4gimo2GifHZoQuw9c
2n4fjRlmmITch2jliicqeWq6h1E/7Hy49lAI/4lBJGSYb7gAk0ybpk/DYyvCw7PW
g6xeJvLTjgEtaZ5X3S0rgUqRmg7UIxdaH2rQ+Sl6XE4AOvP18F64JyhI8UwRLo5o
foz6NqtFkcAZiW9Aq1wmK4mIz/KPOZvu9mKPgUgz7gQ9INCeK7384EgQ74yw4fUZ
yEDCL5GTgdKwD/kL98ioT+ehND48TAqGaqbvHNZaRQhryJ83wswwa/+JQrNft8UB
rcq0gmAZIaV0XffDYn9LcZ5q9RJopRqmt1Y06fDhdB6s4ZKZSFD2NZOcrO3iz6kN
EpbuBU1CEEvx2zUI/h/7gBi+4GnK4F5qMUfmmDPpXB5hGlTxmDSx85qmdmK1nLQX
PbnudVvV/3mBAqPuQkAX/5v5nejdZizzijwHl6ENHqLHaT1KKRp0yQI1QAcVUL+P
ULbFub4asBFBlQdnrbkNcPEj4fs51uT1aMzFaTQdy6888XswFk29m7I+vO2M3WQe
Fm4xp+3+C16WI55Z/1BI2OHH50+4+Hw0Yv/7uQmqCMwri0Sl77tyagH7UbcM5+Ec
FgrSLMgqdRYu2sfQvKBzCg0EE6jli9Cb8yWcJjL/VGDoWfLH521NLZvzIorc2CVG
kmEakyZMXd8U/ITbRN6aJ9OYnov2FbAeI4PM2tuyKwEbV5KK3uZkqQJQF8EN62GT
9Zv7yIEcn/vFxTS0m9Rae5YrIbxxImvCEkj3cZt4NHo3CV4tRQ2ni0PsgIK6KPqF
5rdj2Tyf9kKITIXFhGTCgk4C2bnqSk0QQp49s1j15V6NOM6B4T0XeMXcWVGmY3wE
ehsZoBx8hq2IxJHRoeYXMB0HlW4FjGbRQmcc4YaFCkWxV4H9/t12jNx89zSg+u8Y
QS2qKM+P4bkFA22iC9JtrVKgo5mGEB2Nbqkmu3BWPKEkv3EBPx5185MjABIcsZVv
MFRpxFKg9/5e4SMDU4CxR2yxxh8WbHiWW/SLGlnxRjm3as3f9Jo47d/NXcEfFLEo
woWS/+G8+EDhqITTkcrNjak0Vwtxdg23bJ2lh0GMTDyxHrEQxYK0H03hR4cG4Sio
bojwnXB2z3wOUP2Y4vsNOwE43W9qzLIiHiSf43Ysnj9yom/l67xK39swNstGczgy
o60iO1XFmIDn0Vk9FiOhs/N3O0NE3JLR3ZpFLSFPagYkxhMoak04KnUjdE50tkBr
fMfkcZHWiuXGx+NOTQL77QWR+kHSYAbek3suqpCF/AiPzRXWihczyIfPjegKDIg9
85giw9go65FE461QwSO92QHLeKVM4Ge+YWWxc/7wu33S8lCNn7CO8hrHzTLZOj3l
HAccvePJmBIVqwv1Yj2PMAlDtlBfjt4e27MzIhhwZvEOyPtREYcxIYJ/lbt+gG+g
w6HBzOkJ25az7oGcb5Cp1DFp5K/t/2/lIfDwt4tOrJv80ViiEM+K8Qfgd4aXgJ9K
C7KE9sGphPZuMTsG03YHWEdvBEKPf3+JSaf44xCPYr2zSBoHEKtecHb7xG6uAPmT
ddUa6CBq8ZHeNBWZ7uS+gf+WvEgAzrr6qLWu0tUQxsyJfa/x54On7r42Sy0bxR2S
HytyjuQkfxUAZaW1Um5S6l61U9FTQN6LaMA1loOIV7v+4y6Mjd47/OF2N0ibG2yP
kdG+0Oln0+/ULTRBJcNLTEFYWxOCvS72fXQofxg2eb/FpqKtgHJzzmJkJoZPrEuX
DL96r8QTnhxoMa4tt3Ikuue7hpNXOJIrLtIRznnsM9AcgoIdKOZIqOq1X+fX4vJM
vn1HT9OggclY7yhFFaX7Jve5GTXePuqR4beMNbhKP51S4d6/LZBCIRv0ttiCQ5TO
TCxNHA8xc33sFi0xVl3U1rW1btWtJ2t9VbihlSAYeRupMwRJOYmlvNpYjsXhqB0N
6/17/GkDKZqPzwPlQTz0hYgUvE0mrFeLbPdbMUjPzT5ofS7oL83D4DOQaxOTrw94
BtxHXFH0pjGe7zYYpIl7WgP9FyvnFUR/mqu97b2fdkOZm1H6xVyg/ZLbYI3qRR+7
+Gz5dW/gknpQ3z33N+y1JGNydALRpHMHHG8QuzvquwkVpYlRJXoKo53CB/q/cXFB
oK3F0Wgfzw9NRSClxgoNmxzr9msV2k1dpIZYiS7MD6mOHgCRRuosj43iUvm1uEzh
aPGpkzXWSoBVg/ws2dtmfgfvj2Rulxwj9Ek3OsXXSU04M+ITqNhYp8tLk26bn91o
74scRMcpy9W57OJEH41lpUFQV294V7l+YNgZFM3iedWtkrwjSHiwCC61I4MtiNjz
lhXOQdUjZmPwmcZOTWWpG4XZDmd7QD+ziWSnznBygqgcK/mil9en/wUJd4EHPtwO
ssVzE4ZqYZ56J/UAARamWNlWqCXdYbt8J3jhHqCe2BO7VstbDcWCcLcP3G7i1snF
mdfyi8cM6A3X90szxMeE5IyJpt6q0sPNcwWchxqer85iPrw+tjvW2RT3IbT/2Zbl
aArNiMuJuBZlwCVnyWj0Dnf8eDiOzP8Q8SIUyiiQ+xMRrvGX57lEyv45CkBVULqX
d4l6Dv+tdb/glkLs9H1MpMSIa/4xuVpTxeTfJGBNc3t4C66N6zO3pw8yf8wSUjNQ
7qgEVDlJ3A7e0HRF3wFn04D8/H1MNtdPdTwze0sCHULCJBTVC28lYsqgabEkv3Bt
OVOecj9bilhiN+vFaQDL4T6CRpkxMIzQPGqmYBBdHEDxg2sHmHgsriGV4BDIH1PH
y8050Isfn/jZQzXT6LsAjf932wt4eT1oQ/yoap+aCjMdd8Yd8xvfsssR+VzIjBaW
/c7IvCID6WRjIxB4xJt07ADvxK9LP+5+yk+pkAbjWNWnTd3DEmbD2ic/yotHhWg6
e3/fOOEaSL8RTZhMQE21c0aNarmDDH2+BjHs2C0wflAeDv9mGJLlFS+7WSkDH4vv
1Ea15k7LxTa4pxk1XJDPzSBH2MPy0jHaLal0RFULXwqgTVaTzPUmS0z0pOfD/kOH
ggnEEN6S94n8wb9hbk3FHuIQ+I1EVbG9j6gwA9IGe4PJe7HNmUcn0f8DedKmop68
lB1g3fJzoOnkV3JRtpABNlUwO0i3ZXeCj88jrE/mBw2hN/JirFHUyVm6zAEypRsx
UmygLQp8dqHP9DwhGB6BqV3LoA5OTpDVNQH/p+N/mb/ef0hlliH0MrLP6MWiQqYL
O675MQtwTQuN4EzNe6NcPxtppfldnVJG90qR32dIO3YEXY+urltK0w9/ovmuzHYN
nxKzFbWcbGy8Brz/FxYdLYxXKqc6E3ySLCnMzgDja+fL4v3v9/O+5RKEqpP6YjQL
WZZP3e6NAw4lMFhedJ1P01ZkUfRAFVmMfxhimaGixBe8JZyspZK1RhBP8SIx8nol
y0CKfNF+IqRq6dBREfsrThRfnwEtwq5ag91TYtC4S2ml4ACyAA5CmvTiH94mcQGQ
wk4LMCXq874u+kkbnJ4VAUqiazIOwEQpOZvr4xSoY7EG0r8fELY1XsPuThmUuXdJ
TzgF8mnhUyek5xR+AsGLgfEm9M3SaIxcfSGYfH04ddX6rJJFNslXFjy22qavDWdR
KBboKWpr6nNt4sVxfgXUNXmZJiO9yfNgwZlrkRdJzzKpWH25t8ZgTBlldRR6p/83
+QUfIVQfRTPpL2gCBUZ1ijr5UnN5oNXyXuf1rw4r+IzJVDPOptsP1DD88O8mTFbD
+yLXYO/NbnqRSrCev2pFcpIS4KG8lKa8PvVx8CZKH2b0uVCy3hagzttzAdcJaJKf
CbIZZEpVd9NjieickXlwLPODUBr31NN60iy2XnB0LhtrTUZRVjoMRHSa18HSC9ko
bvuUrL3XF3AnsUXAhKWJtBwsu3CrAvLYKRl5E9ug+nEKbNpIORO5opbAo4uO6odM
wkA+TwfDPamCpfRDNEs7xQDeUfaMYhG1mNkw8u5/IFBO0/02hdjOIHnoGnwoKZIc
86pFNv7xexAjYa/3gK+oUu+fE/ghm5/xXP07QviwiNi6eqTC4O+L4SoQN7wU4sei
TaQfbAj2PJoK/M7tDDlLHibI2IGXWyotGU2j5Vfq8KzxOWBNnT168qn3PHZHKa3S
Rn2zgmrMEz45jpyD4S8srrTUjXprw2qaijnsRt1vSKbv8SnqY+Myxpmn2+D+ZzpK
7yne+WDJ7PNBxILk7KqnvcINK2o2happOgdK9JMSX1JOteHG9/5Atk7WgdIkYMR9
L3zXYEtNr2Y5/RWV8uMyCmYcuYeTvJW92G9Y9+vnceuosGUUFKmfejtu0zaGDgq0
j4N/9lMXo2YU1RlSqErFlc3YsmTAqUAnVrIwLFNIeYY+K2+pZqOePIv8opY7g8ct
Z1tEX0+GNQ0p1QSehono/4Zizj0JjylRphak7F9qsdzTcTB8D7GyOh+CFri9/WfZ
HXRp304TZzHVX1BFwyZgg57iRCF8//f7qc7PwMGOurAlAaLNbUSdZmB1LQTFkqcZ
X1w6cwR4s4wxmERfHL/FA75Xtfk3KTIXNLHrgVA/OthWmNMQHgrLMt5bHFuFpjAt
+S2I3pv3A8J/7G8b8xMMOXt+bkbCk5QKimIr56OaskxGbTL6rO/BjT2HRguAwKpX
C+xHW0OKpWkC22ZQyGdcVtRz3/4mM+yw0nR2lYcrsX94taOSvK2wEERz661yJf30
mZtBdtkk3uuKmx4JGwvxb+z0Evize0Q9Jun+ZyVqO/12d4dBD5hjp052r/Kzoq6D
txXiUM4i+ZPWh1kQ1uo+WEwj/noXpZbqqi5F8ATzf7TTcMi61/HnjC/sLl5qWYS9
Xpi5227V2V7Vqx7NRMz+FLEOnG/XLWRvOBVUDwcqtTcfK3me7eV6lGbbaHCNXcdd
tWssqghxL+2ODW/aUVEQIzWTYYnxCHnhwpj1ekIKwlfxHqpd06iEBZmo7CuqUHht
+5Tfwrpe1aZaxq/9k3Av9vxLpl2NUt9yzp0XVgbDSWCTrc/76AlFWrRFLiqUv/1k
mbVA6hCvhrHRO5lCOApsC820I1v4/I7uo6hKquNvNQHzuzBwGDPgCDDI/BH73cL/
ftCq3R7fVAPNkc9FuZOpNep3+WdlrFGcVNjBThWsHm30cqGb+xD673rdkybCpVno
Brgb8lbRStrqiDRBzOWBp89naj0AQAPu59ga4amMcPUTMHZfAn+kOC8TOlfAYkIk
zXmcIMckOiTb1bi9f8tXmNiK7pJo8BeTqbhneRHLqfewjwQCzqU0JdJX/v7JIioZ
02pAwrOaw8u+iZwH1j2pp++lHPzFXrBBf7tKPX51GDl4qyh7mOY2C31s9DNzH9xp
7B3oCpEm6FWS5/wFvg2DnLmRqNGwnEqZa7iDEJ+VMbnSd7zWRgrUJliFv9+z9KEL
YBT6pqM+Zmo9EOX96KkjdaTZvI8Xo7S1I0rZg844V5LhZ9Q+L++Rj4FFdogf962y
Yl9+ojiT5TNTjmj4OuDmjVlFawvX6g/MsEk1IrACD/ECf67NLXpw+DigeuY41ihg
khxqDubat7I4jF0j6tRzmAujTl0ezxisgb2G09NcnbfGJcxFh9OvMXnsTw2GkyvA
QYJn0S4dN8dzxPGUek4lh2/mXbDi5P4OMMRwdPOjqN5UafnTLONYLL20hEbW9myW
dwH/vl0Q/cTzjyWjorPvl2uNw1X5nIY+OEsPjQ7kgWHMnZYOMwhkkPhrsre+ySun
I4jwJ3pYhxD0afLvPaXyl2YQALdyXE+RbNjx+LRdu9zw9eRIMzb4tdVb1RaMdVqm
Tz+nWVNFn5gluGY4JsAbx1qogEP6TwOm3dRauXyxuXTGfMBs5OYDnR0UpCTZ/c9m
OPeygevJiAXQg3hDxzEMZLRp0OUARl9kvbJMtzZSefxq9RqMipHFJxBP7pZHJWWQ
GLjtNmLh+HvH8sbX2oKnVWDKazx7sVHGE2Ek+zqH6zEFjd5V9bj51P6fR2HpW0Hn
1mfU4oPjRNr0kPeXhzS8hFj5QFqlDqiOMSOi2mXUXhNmGOKJJYtrcT8/yEClNNL5
hnCiu5JbM3P7vruS0iGY+BhswaVa7fQP5tW42fwcrPZ41ILE2H2LoU0mszuzsFBK
YGPGn+A0U+EwWfgqoNDOe7C0W0jWpb3Xm8Ipbul6bUuGjx+fR0kYkHWoqnoqVvF+
BqfT1V5cHTIaMHPUkUyBngKtPN4Zy14uLiWhlrwS8fR/KTQ84sQQ4vgiveW7vlpw
Bvh+57dLN4kNoBk77R1qJkoCZETkZgrf3SbggqFkNKpm/tXTiCYbRAlVvzzu7CAh
bexQJRsdfvRJUB8f3fkFvfrOgTHtCW1S4AGooqYuoWKYkOCgnve3FPZ7zdtVarNI
wPFzNv5pCnp46171CQeYvdnn8PpoG9iigSvS8v8TKMJ1WLY6uAwVj+m/NSJvONsJ
HVtTY4EXYxydIn8R/TtS/ohcd0JMy0gyCrp4AK0cFdmCCqSy3q6pngJimWbtoRD7
exCvKEZrwCfQTjnhxVz6eSRvVwC2yCnaDpwBNuh+NKRYLi9NTBeC0E2Qi1aY2IWm
+9k78GOavK5r4ebQBWb8xqfrDWoocJUyA4BswLtZQVx1JPTJsIiM3OVTTCKLNWHQ
A0gJVE/Qkq2MRhro0vd/9Pla090uDhw0lGpMah9UdvCJP9H0PT0LlUtJCtOtMkag
vdMPrW4u0f//dfsTXvsj6KDK5hIWOT4XK/Y6M3PVNDo6EffLfp3UMxN2TLk+XHJn
3R8kgPkJSbPVpLYS3M/hx5aUGAWM2kgZo/F0GltnA7MKG3Se3BlRrnS0yKV9W7I7
A2woPnrhLfXeYVMrJy9stEXQlSh+70A4W+WXebzWhJp0boniRfDNdjrlNNVkntZM
h/EPSjKqHfyK+faKVWGN7Y46kTqIrI6aO66WjfhWyXrY1ME/DSyuQoWcWJ9TpaBp
hv35yLKeCA4asc6MdecrNTdc55YOZ11qOQ/w3fSTDmUPJ0jagV6h920h2HkwAiL3
nO8LR0FoR/26tzFsrW1LW9PoGRnsfvMMZgZrTP8z7R+eioZKNyRHIvPaCnZXk1Yh
gmL+KqshV/CXNCBoE6ID7/fVdmVdt50002TVd+2y+wCCF2C3BNpJkjeDbG17TJ3F
llEdB4KcmANfG0j1eG9imHWyJgiDrjkDU3JG02kTCR1+UFLldFpsEsnKIZHCJHbp
Yk757Z3LzR0JFn8wNo0laMDjVfOhXIQ/R4F6sayjEFFMBRvFs4EGU/36YnQZRokS
sJsUfS3zGGRzroTkPFj/b9xoovuSlFOcpI+E8ajTyA/G+i75AGgJ7tIP7XoaxGHE
kRwidX6OhMFJ5qA6JC0DvGGCbzs6GMhb7mCVxxQyFGG1Y76u7DfkOVPlHMy0R2PD
ixxevF/xOWyXpqvFqOzWxJrFKgVzkS14P4IhO1JWuLlKVgBFxyK+0uA12kvQlUZA
3X0XPu35xOlJUymmwcWwsxxrlAkydQlvfJhwkUnLfYVB3kDUVp7rx+YPHCjgC0c4
g5M+dxoigEEQukTgWuH6Va8t0Ez29KxC43v9SmGH545AMMbW20wGF4ChGaXQDugE
g4anUoiMudczUUjpwT12Ult0EfoXkokr8zSGdIquzV1WGggnkytBUo87QB0Praw+
1MD8rb42Fu7P6PUTjxmu0a2lbLbfdL6DvLl+HZocu7luSyA8dOlKNalViRQ3yThK
902qncg3OPCDAX6k2bJgryodrPpPdP6KCNmX6+ZE3jSAQ/fmxi4jpYUw62SXDb98
rVPtMZopyK1R8QI755dyhemZhua127GFGkRIzF2jXt17KHyn4qY+zIbs/tNaYVk9
rmYoLws2vsW5Sm7f0gYH+kuxecY4jZLdoTM9RHDXI/lRWKUAFQiweitJQSx+zCF2
6vjFU6Y+LUXTUtQ9r2M0DZeHApqDlOw6Er/lS5jOtuN5gxTfhHWgBQIwAv/i4xne
WAQemHKJlozwRcnAcJGy83C/5dk+tddogNLRikVbDx7q4EH8xH75Z1weG27AECHE
UmoRR1gFS5i6Y3FN1XXr6238KeXQ+O3eCGkRb1yvbgsrp8TMuZLXtKgJSQwo2vpU
AUuLZT9MxpGdttNR/uqlNRxF7T/XKSnN6mGr3YJduSUVH3tnQr9/OyIjdtndSkyt
50fAlmCTAsDCozGCa8CIKeXFQOET/u8VguGB4nJ/AocaqA/B2XsX+fwwUMNcLbjp
etzQXQS59TYI9jjQN87Z4XG/iuxBnA+u9ZKEweRBg0n242wo1en0+gOcGKd+/J9h
OIqjIGoU5Jlqx8PV8C8k2Wb0rvMozlPeTlfoHX6XFlhkC4CVZUndO0KW0EFOi9n+
QAGlfXP4CwxYG6cELsE2C+uuZpepRr+Cftp4UudnzKoYvoDuetoxXgjnnlTP/FkE
AIge31WeNz3KDHkMHYgq2SdekerD5nPqf+GUI/wnqydudapU13HovLSxZXMJSPXA
7PqvsWsQ8d+/ucXC0YTr0+VeysAcbGNEVb1urMFPA/Tk1AJrqdOhdO0hq9gYqtEk
VIHqtxS+GbogHSROdaX15DUoQpLCrbysLg2LRECkBIUa1+gKKFljOfk9usO4e+4J
jufbp9T6OSg0OpmnGx9MXb21jPGH7gJcV31HcdYoEZzaONA6ZgBQDZw5yQujOvv4
ZGAMYy2wQ7u06Gp0teyrVv+x/NM0yOW30ulU+IDd9SE6Kh8im4QUGBdh+yDyNo6X
e0SjOaIT52oRJV8Nn264lPc2ylHZIvESHRG/uPP2roxngxQvTggdNMDagaRiqe9S
1+8+umcsfimno4J5EQ7x2SqwqtptSsfcWaMlF1mg9P8pCC0LbYqq9qIyzE+fkdg4
yTUI9va3oeB4TC2TmVVFn7XcCDF0QfaS9NlgHdlr0AFA3R6IS84pNRbXeBZIcgOd
sTjyN8pbU1kEIFvCUqehUtiuICPTtp2/rf43dQKepAYU2somTK09W/7muQbVGsPk
z5rzkFdODfNZajPquduH2COkF/37Dhqvku0N80rtrN4Ceygjm6V6eVA9Vybx2GWi
ywH2EeVEU/Sy8Mn7ANFrj7zAeDbpUuBbszp+oljzY3yEuyE06NmeeksEOb7cjqEx
2GPek4ESGomaiR0f7C1HSZ+pEuX1KaCwQ1dCfljm7NSGOlWn8NPmxXOyt3LIMEt2
WcCeeolrtDBxdfK2UPKF/9+XQxn7qTTBHivRnp5u/6DJSNDsoS/Lbd0eVWWO9xSF
XAsTuXRVl9QIC0se5/gjVz84FxN1Iz/RppKDqvlh2g6ux7xC73SmRvxyJxuStUeM
InTV3thVSP0uwvR/wjBi94qYy/1+FkUZYgttXS8pZIMb+JLmGqqu7hV6XW9Dlncj
YM6wie1nhnzZr5fb9aq44gxd8mjKmUKY8xHOWTA1pNM77H2qYMXjMttey54zDzxE
Zc3OgWgdB+15+A/khfLD6DZwijSHRldLMpWbZ8QIx3ERckQPri+lvC/K3OGdQlVL
kQDMh2zTch9hJnEmiNJFPYd1mw7AzjB0falTNfc9mrsfemiyaP+79JdDF2UtEjB2
M8akI4JadycDx4nKEmWneBAsyYegMqIPevSY79p91RJHlOt/b3Fb8TYbTTxt0qTP
7bu/x8x8C99oADa4bITdsrTi/YVICKJ/FU3D1T8xLvFmIXhaGnDjwiw+xNF5xJ5X
DI2A0krL3P843cocki9vIoRROieczHPfy4vcegmsG3Fvg/V1yQCIPHFDvjZQb+AZ
RsNxK8Xy81P178I27ZPndbBR7g4PXxUBREyZMXuyk0z3S2YGVXqcmPqDp5ozGhwW
f0DB3VOQnr2DKMhLrBWN1AaLkVtqizXQVefXfi9q6uwby1mbhXgq3BbVIUSAIwiT
zqVM8n9u8PzK/AxBbKxdXnPknhCRviP35t1hNltKdZsDOhDpMotsbnzBCacoVp71
oJTqpKoDedfn5zFnBGxSjelk2ljRrlvKGeP27bTLEMyGb0fA1FRQubcLnN4KN2cd
r19aGTNJWhRwDEHdO7kYVBHARaVEY9rQC8iP2+moyo6MKw+GkYy3fr1S9ct5quH5
C1w7YH851n2AdhVet9zFu0KjFxMi8S5WTah9YOLerHMdx70fSsYvjYP4gVhyZDqq
MeJhZFO+CBTnS4jLPkiVcge3w1K3JiokPG1BlnfWYOmnffR+gKcFCFpI6TT7h4Nw
49d+2QuvMW38T0P5f9mzsQulu5P65QjnJBW2bkB2uDkgFcR2IncyYM8dy15hV6U5
85zMdAKY5v9uBLf9/qxQqw8ZJyx7uKorUucIfXho7qH4oqcqhl6pEqkphivhZKHa
OUuo5Bspu7Ci1Ne0jJxgJ8tlDfx9dPLc1ydFycKNzdjA3MpGxYF3uoX0wag7FyAD
st9tgsL7+RVU3lIu4u04qidKpvMCdvo1qH0z9nN0aVsuyFCUgUtVhW7KJqtIZPzd
nalKHfHZnlu6ObGNdBOK+dKsrcjxEHwQCUjS0H/ceQ84bVYXunCEip3bvdnmt46s
8fncnLL1JtNvWYVkhWo5qXxOh5Pz+OM0qROfBGaR00pCVqzja7d2WH5vIjcKk8IQ
SS3vISkwffpP1KmOZ6bzJFgrQpdStuy+LIehRbBHJscipdBEEVicDF5OnBTbwiMe
guqb0w3289M0PFHYBAWJjw080Cv2q2WgjKW9K33q5cu9PC9UrL6O4MUpfE4f/6Rc
DqhAjoIjsZyqchPV1W8tXa7CZA7hgoOQSLAe0iPF4JqwnIS+fTJF/PsZIeZnOUfx
JAPHS8WXwVD8mtlKoGkjIXbXDOuKPQcIMgBPoRdiyHjGizC7GKYMgH64pdvTULon
L8ZQboN0WyjoqBhuecnBniIhwHjPPrctgOuktXLCfLLPq4C4NttGQTcpg1L41slq
KxqEyIiOdaTaM4caUQAgIX7cNKYYVBE7XDHr8zp1U1NB0eqC+IXtehGRzVLuuQ1d
krTlzjtG/aKEc3VtMLOO39n+hXtAf0/p0jVVZGKKXf9djdVGuyysOSnD8IhYIEzY
YQNJKzoUagXSwQdq4YUvo8j+k9AzTZs/KfKeUvsBpnWPu2OiIjzmW+Eg2nLuIdVX
Tl8CZQdmbo887+2AgHXu1H4pbMLrfArb13HqFGQ/VYg4472CplF9Ag21kVl6L5Ns
CXzfp6mUpGHC1UtbTZv+J/ZvOQjsqTWHNR/DZFRUU9vQSwUrEhMkhigqzsbhvE2h
kW/iN+vq/BGrkf24GKNgrUJoCJBQ/IUYpXabXVs/Htu8sW1MIE/vwxo8azm1bMO4
FLDaA5+p96DsCF8MRoLNeCqYOBpTl0dyD7QsNubtQFqrAurRnMgPAvSKFnYOWW5l
OtEoYxJ8MpVZldE4y/kB4q/+d2AEzhwK0hjUSMP4+odYCsvn3TOxdqDAy35nu5Pv
TX3fauPw6KupvMrgvXYRf60gPRjrmoC/yLlrN1QYouTDO+sa1T1ttxTxKNvOtbRQ
/yvB3RDh2j1dF1wQsfD9Re1h3W26i1PXgpj8tYwOjn9Qqu3rRNxPgjucRFn+ML8v
rB+WbH1MpuHtBQvwPCOI7xxBPOLQq97q+pyVC12m0kJK00pdkJtYcH1y7Yy9AVO9
TlHhzG0cgCxZVvZfrJcVR1JV25XsBvGMX1NJkaKvnRLRje5tS1kSZgm9mcRlKrY4
5tLRP4czyW+ILDPM4RdezSWf7rp1Nt/e9F2/tlxs9vcQNAUCUa49oI8p36B1EsIk
3sYWA2MKVWbZ/q8TrtYJ7MwsxYEPAfcaWcUhAnBnQAy0mmWzaaiGP/N6PFq9ZMwD
Jv33DJerE59nsZIETsPsxIjVGPPLEFQJu8OasHDl0x2Kbi4Qay+YjNxoHpvFrqEY
zZOZJXGKfnIDFSn8MMUE9xXkeVGecN4LjzOJ9Zatfi6ulLFQrrGpcj+AnO9qYmGG
wqOL0mHn0SZUjEy08zXG1jsERs25KBQ230XN9EDeDNDejwm8zFkOEHVtNKUwlnXg
uxvcctkm4tcJxXNu40Wfm3/2RnJM85tNEW4fLnX82MlmbfufgFsmWprZfbpHPVo0
YFV7sQCTLBukVOY1qnkdsuWCszXmbfQ34RY3wBcc+cgrF/jdMTvIAGwtSN4nyo1s
BhLzgJhwNX7I6E0XlHDZOfj6if+O+4CRBnJY+5vyCuE1cd4LzonkcDIVc0cxu9kn
GYqck4TW35yPNJggrKXhO02QQYq4pRzTjcidf0vRCNWiOqj+ouCIcEX2T1J8BoMs
Uagwt2kJUz0qP8EUtNGvVH26tHU1Dd7VDWh78iUF62x3J+SZuGcGsghnhnWp/zV5
4BnR5Q/se0CricNmGg1Vd4MZ7v+50dxrIkopwgineOJL2MZyc3JlmuKzVblsPT45
GigDs6aIexIeQJ/Ctbgg1hqC1nhq+kD7NeyNAfQaED+e65RlDFdSIUBMXVZUmAls
UKybRaq3MD7zCxl49LNjnBXhoFcvRnHPu4CHx/FZo+/8ga7dLO666LXINbnbg3i5
02dpjquKHhVeSmNs7QHNlcHkyvTL8YKyqQ9G42oYW5PHwq9+hDXmmKkQs0okLyrN
KPHQFlFvsPqle3MKH10WtHe8C0/5QACpUnjG4nT6TlqXbvkOAN8d6htJcA/DJkU3
3+DgwrCfPiTDWSqpUvuhHsns1vvON9Qh8gDRxtjmsWAfGL0it7aV5ewlwwkQq/Vz
vxdrgyDheS/5ET8jfD/6zWiO/OvLSoI3xCoxTTBIABXBRT2Fqb0KLwStPv+A+Nqa
rycF5kojsJILtxf2M5bbM44VI9FbD9MEk1WWmILo3+Fhh1u3NmBl9qtZdX2Hh855
6NUX+5lGcnnDCfVF6+Idv6s0ZjCXFWhdJ/0ppHQJ7YS2HXnjZjoMlWtcKQ+A1Wgs
za973cin/vE41NpS6NHW5ZCDRUtV9OKX8SFPdYo/ssRiIm+L/W4UQkhyp2BdzY0S
fYPuqwfmL9N3BCRejSiiPv0Es4CuXxbGZvHyWC1Efq07a28QkJtYT/xFxTKR9TzF
HmYlWMtf6SZW3U8F4KLXWnAuMEXKxCtiQT1NZYyTaPwropvGB4MBOAD//KYdUB4n
K4RYofcCEUCTYKvUs28SHX7IS55uB17rl82oHhZgjWSYfcKYr1uGN8RvqbtRBANU
F2B0euzMXfArfD+XZSHabcG2F0/M729XbPhjLh4ZorC8+FRLsz6BxsGWKQujbENH
5yGcPGHHGryHtt+daIAsyY0B5wymnGDnUz0yTFuQvoiDEwWuS140HAZIIkK10Gog
JFMBng8VAmuLsPXahQNXm/PFlHSN4jB8uFipIBGuHuIHB8mLai/KLqe8HLRs4BMU
ppYnWXfGB0lVWMDEymyHToifiBDR2MCrC+d6Iyvby7hyjjVIAMx5cQsLiT+Y/Hgb
qAcFJO96ohIX4xN4x30oRcDXkcN7C9TmL7ADNezYylhLZ8GKraWeX75nvTGw0vWe
kxeChLgxa1q+af4zpxr3+dvIRN6INbGpKx9qhs1vnYTj2A6njI+sCWT1svm6Qfyi
/xtjimIi1h1LpDt0/i2u9bkL8Y30YQELmjF4uh7H5RiOyo91TAB87m/xUMzQ1tUo
eN/UuBVMife0E3a0Mc7T/d4a/mRWa7buyCTlX1nH+FQnIK8Vhk79BkQkiF9zQDy3
2T+z9CGRI/DPr7ijEDJ9lQC53YQcHkJEr0zdVQEjid94tYRIHbQVAf3c4PKpHkN6
d7K2VyUOiu4gKqOB0lH4wtZYTPRh8eNRDfu5+aJsZ5H861C3oGN//AYgebkOvfoq
GFIx2OPqfh1I8D1eURFjhX4ox19eqLdYCkfEowzaxwIbxG76GEA24ELEtpIjbqCh
0BTl5FJwLdS1WNH0DbNL0OX8rmZ9feP2VthZ5lf5lrqsfrtIOZP+Y4sNtb9G/pDm
S5/Dxv6HpQh/XmgSGr87uT1qcgmQDMANAew/CR5w+9cD4H9qEyDyhO7UHblgyCVI
p8WWvGv/KGRI+R8lojG4Hng3RzN60Pb37GNAMVfETXwXbfn4JO/mAN+9IpjDQLqT
lmAbYIhMRWNYwQduNLASg12gX+qla9yrqsG/ytmqUIEN6QMBuzLcrq7hY5E+Vk3r
wEClLeMAZA5AMF1noVpGDIzky1dfgc3V0yN/XbbbHjdmbpZUIPhrnNUJjAOsxOjS
uo0/byFRzV9n5L+1kHKQyD/YUQbj8lvEVWrHR9ANw2AKUecXyNpQXxH5Rb1IFPbw
1j/gt72msx6S6PnWG9Zfc9Dk/83hZpkci0dYr5WaWp6K530CZq9+1aeEB1vuwHd7
pclPKasdOZCCvuPLb/EaY80ZX302XPZnVzlg544a5PcU3fVGXcdkFO3HFlm22mko
8IoTmjPhRVAiFYELZ1zyF0DWneUTxoV9AhQhA5GcW00kqB3LSSVYY7VAPs7YBoBI
wck/SqHlYKn+iMyV0idzxTu5adiigZyiKvmB6G7lBN1rScn9VI5Vf3xUwp4N/bjo
iYp9wRQSe91MPReK5+QISG3eEK0C84g7EWUE23/4qOQAPyw+16QjeTWzEsnGf9WJ
ImvOi2AYx1ip6k23oGU5XlaFz/6Z8i+caNdpMjYa56eziSW5EtsoHUhJwITInDh9
FZrscD8LL/Jy8TIs6OzbVoLUoB3y3V41LIXf5wpodeFS2gudciEVcnYa7GTP+RaB
DpVetFst5+XuF6u25r3e8QK37ztVswfNB2D3BBZHdHOE0zPMJTlwjJMb9YGYHx+s
WRk2U6C+LEOZefkHz9kW7+UuS0rAX5xB3qvb7afDNAwv2JMAm5NiZXeJVBXegAMS
VJAi+nsNl6YF/9uVXAAHMdN3Eweunj9PoDMuttrK4aZAholxSUY3kwS/EFuePDEy
Bo5pn+nUUd+Ns0XTh6qN8GHwKL/i/w/URd8DJBU6jcyHCBQcjbTlWCZZ/W4P7+g+
Mx2WQZC4CxU8Qt1HqcE+P/v8C+jXsn1GFHIsLka79c9x5MAWJ0aq0U/S0EWTIqxS
7wkGlo0MHjTMTdub2mqkgD9F0f5AkoKc37Gg5fOOSayUpuPPERXhubdcpjmMc9ws
ZMSzdce8/CnmHAY2zuHOxk6T0A20y9qlEZcd2Ho0sjaiXlOV8ds5/M/aMC1xcAPY
orXk72EhmWxpRTmpHWgGkibRci+ubT6f6Nbo6wj9RMB855iYlx3gFG6X0oi/UW4T
/RlE5yIBO5lIJxs7PYhO/H8ydz775MtWdqq3Xw11FofZ5vLApyk17UZ9pHy1CzcF
SoaUjDqDiYAJD2p/aedFhSJBgblCI/u8DJdPemoymfEKRMbzDMMvQnTkDnMAo3Y0
0r+vFmRyjwjrD2XocsB2UdPmjViaFdlJgxUke2KDvNGo1cW46HEpbA+OzpYmtdA4
WjwQbu2TEFfjvNIR29+5B6qQX8Xqc3OA8qG6wwb6nmkFDHn7C8W8SmyZXElX1mdD
jzSWWk8zbZpzzdYrY+khJAslN2SksV0IKX+nwN3B3W9ZoMbcovgjgW+C/eaFeZg6
I+CZjHcyA32qGuEwiZ1fbhEYd5mbhYcR0BzoJaTkCAslSYv+F3wfVpGKNJ3/GF3G
xvTU6dr4rwielg1Ne6hEIZ/ADZeos6CrwMoUe5Qm+0G5DfdND/gAiPDFXuQGu+8F
4bniBW0McEA+FiupcrQ7wB3F8mcrY33DOneZHc1UU5uW5aiMUUS9PAcaPSQ37lyu
I9qGlmljtEq3IoaHHb+U9dezKIgXkaOpTyKjYg0UyZ6STu/l6uMZ2QU7nFSDd2Uq
BS9l729gyKjIk/KgLy5fuW+TnLbKwa24s7A+oq8r/tt0oxr9HT+DIEPw3Kpmul41
m+x4hwzENpsmZvtnZ5NWADk+l11PgHC05YlfiC/Dj2JpMPX9nZxmqdLYuhhctd6P
4iQIeNzp1fAQLFsAQzCVN5LHNil6ofeczryr0elubDVAOBPVubz+Zac0yBwgCLkR
M3NcV9Jduv2ieajD+5wwX1b3PXuVI5piMKfm96aVLhey1/3nnjvew5+azYEQTAYx
5VJ6SKKKPJ7RFwEJCfgrtbaZfVj0cPqy2YQwa0amzPNz7GvnDBX+XrrQgTH12++X
1Ge31mvAqv5DlQX+Gobl1AHIqfEhXI/PdlwxMHE4X8I2MYC/W5Ff7F7RJ51YVxIi
ZLRDd3Hu+F5BcG2zuSVzDozXm20Pz2EBHn8GPqYuTk1CjNZR2EUj2p30Lg39gw1S
CCUIBGQcOH+sKHZjq1UoALRtBqh0nUYSfozz60W40KXBGGiucjU92Py16HA8oD1p
w3SiJsVzewqLbHqq5nMHm2+4KQiLbXo/bkgoaXxg3XsHfw7p9cE9Pvye5SX2fe0O
+u+Gvk92Az/c8fFBn9U6efttroO8+XIPi6xGOpPHXo4fTz/xZsgLAtQG2ilZXwH8
hZq+yT+kxriHocN9lieKy4RXnm9Z6PKo+ZzUszj3PyL7GqoymN3HJ0tOfs910Eoz
pJt1AuYeJ19sHT7HqKJRIpUcNNBajO9UfF29IBHPWtS8wLtCcva3BZiQ9d3cUE7i
5UX2pCPjZztW9o4rHvS6Rr/KRdojhLiIFHKiPta1CjKa6KuSRVMxqbpDOqKV+5e/
n/25broaTFJpojLgmBYRoK6DTCkyaVCI8FfqZzNR0k+kHI10NsaMLB9jsPTSsWFS
y2NDaY5OVrBnTnCgOt/+fDAq4bFs3cVmKG5bM6T2qQK5R0I4b6QWj35Pv/jxb5lr
2PTJ9MzY+TM5Uw24TIBun9eMglKyVUPLJr1xL7t0OBKY1NMDMUxgJeiF71mjNgme
62sO42CY5xqk9nHktWHreUM6OUUg7ZA4Go5+B5fZdFPp0UySppcEDkRCmFq+4LTp
pxSCoT5Vw6SUsrWGIIlfmeD4faDCVZfWjVeHudO2jV2lxOHE3Va/74nteQDc7n26
uHvOPxvvyGJV5WHZFVJ+qhtGrDty9m1xfRJyddOm2SZ+m3zwC/d7jUwD2VDFky/v
NoWehpkbC7QIyCHCKv9CvpQeqAQFuLjhtRu3w/CuVQK7QjKczLL0Qtml0KWBIyqK
M4MgPfnKkU4OWLlqTN6+fXPH45VsW+9onUbkJuer2gSjMm8yX3Ng5m+Y9xUiecU4
FS5tC6Uk3vASdE6LOJs5tlc/zoAtnxfZ+yNmKBmFrvOmd2CZzItVU5V8W9K9pYXC
eOv4J1b5mD/nCrofGr7IMdVEjvEMXoJ56LfEQE5LLAn0hsmQ4dD+3i+Ny77B2kJT
qJoSTEGk3OcK/2GcH8GNpWr+6LhJ5A4T5f4jeoI0ZxC6IZ9Xss2ygbQo0LjpB3JZ
oa4LFRtNATs+jn28MwlTZ6kqj8BEttZUISogw0goLxSi/yFibafyOz7QHh1/79O6
sQViQVdeV0d/EQC8CPyA6j298Ku+uWVnYE/hofPdfnCvGLCxQl9ebeu/XUyvJt8l
frh2GYwz6Bzem2+ndfdXofDTTsI01wfTi52GrgRoabJNFO7CHRgglbHimJJQIpE6
bgfaI7xIF5047CCWgzR9N/S8x6puHiFi/XhqMx4y3DOl+bEDrUJkJBhUfraU9OAV
DmOlhTANPHk1bgiLLkOzCWbv0IXtE5ZHxOjj6P9tdXArvDrPDyibR/R/GK1/ybjq
aCFwJdXtJuSeZy94xcIUFpUcatkbC+bbXJMbWS9fnK8c/b/qhcX9QRvP6TrWcHsU
dF/LD+alVyVp1S/N/9VehujtmswD5t3hH4TdeYqmN9KVnC+EhKQy/Y42NvyMkA3Q
qzk2PvqA+y2FF+UqIgKOq7uwCcH+6yIcG6lWCqXIE4XufcI9Xvin+dwPCdJZfy6n
wQ9EnZPIUg0rQAr4b4zztysVUE/BSbbaaoBVfmo78UtH68Z/jvJGoVJaCPv1aTlW
Oy3nKV7lkEm7dGm+fXu4e6jkJjphA0qZ/BVcv2+v6Gf5/BCaLSee+d3BAYdzQ9vs
uxm+ufZeYJPG58xjHdYoDDOaGP1gvxXRjzB48U4w7b9/bdlM97mFrqqebmFiqlDP
xB/7pNRu+mv5Nw9yVQr88wqJYZvPy6f1igs62bnUf7JW1lFgT9+ghbO/B93O7u4O
Om2NgjkTkJg0gXsNqSlQA4J1MKasdLEbvgUMUnmnMLQxjSzfothmK7FFY9gisM9H
Hq9XOv3i3Rr83/KhFRvPgmwjmzqYttf6AZ7ZSHKu7IfRQCYjr5lFbCpgjeUTt+CU
N900Gvm+D/4x2NJTzRYZDEQKRcx39RLc1FpCvzpuhEjVnfpmwTemdcXGuelq7S5d
RkXD9g6uUecs1dK0ZUEGfG92JonwMmZqmZrf05CpAQS6r89eg5CMQLP6V/aCYgxy
PjItWYp9qsv4Hu6Tp74PjrvUADi6Omehr3qLthC8z5i64xA++V2lkjDmb7uVAlTL
7xozwOQJ79wh5ItnoMowWWh1ncD31ySohReVlA49cHbiD1U4kbM2pS1KbUAEZXBH
eoxZ9FfLtfvAjwZOX5jbYvCS3oiUfQK0YLEPiieXZEpUr0vOmiDkD+CKKPATH30f
v1+amSw/H1gASNCu5jJHlMFUQBWiYOUq134i258C9n5IjRee1x2c+ZH8xMiIJh4M
dPI9VTpRydHBkmn/du8CuHh6ss1FrlNw6Tc8HCK7/ND8dbWtU/JEIqWBnJZVnG5M
vtnxio9TnzPvr9x46fiiysSSHyznMF3DpuZGvaJs5FhemafPjTamQpcLhw07NdqR
lj9o37449qjY4RaTBcwxokk/qzfYZrdVG7oFw2gGsRVQ/i/KBPVwdYJ6dL9+eh9u
nHXgvS3RtzOb2+nqKxfAvVUBvmmMCnIyrjYkEc18CfTGxdCxWxAZwtrFyRiEWu5R
zEtCv2PCfydLSx0q0ByZ/eSG/16OmfvgnqlIT4AuCZUwEuAbI36E6YHsqgNRrpLG
T9npOoKMDDJTaOytCJ2VGi5F2n/5EKo/a7f9043uoAr4FQEZ+Xh+OYvhZo6eiDE4
BiwH3V0c41XBArohXczxsMQytsUxwML6uXHN9zBXUzzGRRBfqqpGltOz/ZfdbzQQ
TnS2/CkYavksdM2WjzuotzsMUv/gTlK2BihDUfHXtYETSPIAITaU2894jbbJ+6u7
yZGtJ/5dMU7zNmIO4J04t7hX3YpiU7ccLv8JPrTtoDgNWvlXEaBSC4buNfLwwqdg
dL9XHc6fEvead9lQBIJoc6H4EggOa9zv9lXed4DmA9OL0PtFtvDUWql4CP45L+p3
XAqFmm+oHMbU4e8/CfJ9snFFaoBa/m3F3kPGIIMIEtmtoLXcvs22+bDaTH20mNa4
AHJyzJqe/vD1HRp7zZAEFMpMhQgP36ncJqZOKZYOm7n83DmnPzCBtjYQTqub3fyt
/Sy+3Q+ooiwgzqZuWCDjA82mhOCv7cRQmJ7i6dEj+pN4MXPCsATEQDX7rRbgrUVZ
HItzkpB2Pvkj+2KF7rRSqfcVY0X17uo5dPbe8N9DxmKosc2EfKsxYxcUhX31W1wy
U1fgaDFi0Qa/RMkSXE0v+rOgqGQ+TmtdGzoIbf58tWsuuwg0XrJE13DcAE/KZ3es
RHY5FZKnFng+YHdmGWeO86XBmno7QA2lkUBexWXuC48U5gMbjptD0hh+CLxLlV9/
Qi3OMyaBSbdmjOm9umtlCZqz58/7kf3fz4rIphRoaesWFbq0Ma+8/Rri/pVtJ+Zq
CjmqmYo/7wfFSHOd8PUMJhQfHPrPp0CBi/HYbUurSpnFRjGfQJy97Dn+7wZZSoN4
qurSIEtN2+A5tJ9aZruYBEQTRYIMNoZweyc2/66eGNNOynLC2v38NFJRR+KGviYC
QzeX6L840jsx7zGXktkl9kIQuaXf5YD7Gap3vERbTYoMfNm6ovE9uW2xhopwFd0u
Ef5nYlCroDmH0XaTAHN7pHN4pZj7KkAGXN3lzjUBGLcLy9u8nA+jeHbH03DNRf/t
Lv8b1wwArrORRrxcdb/3ixcnMqy0hQ9a7fNQzz96rEiHLuI0eV/JFKl2OccTIGTV
ivVHp/wOALE4gsnAv4lgSKOXGYNAujD33NTPPkP8JlnSh2nVDwZ5PJNfta9bheC9
GICOFCVNWUF8+zuJOUpww7wcnGftMJIa/D3BiChrfCMwSqaZPd/vsGzwuvVaD9Ug
VTo4W3a5Nbj92coWUarY53nr21OLjBBULCDVyAli7mrNzzH08d+e2u25MMhTbj3v
mQuA1O8/WIg0bCLvkvXGRw4GUj0S7x9bVCsev9F0aVdhDRAjopULLXuTcVRdHN3F
fO0xvnXDniE8rhBNS/qQ6ox8HosH6XwJ4hUOuRx8o95tUePKWdFMoWDEt3M7i0qu
Z6IdUwTxKFKemuH9B3SMsPF0tnx/vqY0JfpMRduUkil2KE+/K5+8yIteBTYVOx+p
afDbpQC6oZLMVdthzydBc9yMh2mqcTA0XBB/TqpLS58/p5rZPwc9dhFU+VqeJMww
T6ZI0dU2f1GQCjXcZK+ze7i8kWZ8TDz3R+qFaBaRK373ASJXis1H+WCqvoJ0IfIa
dYvdQfSOzVQw19+9ES9X0ZCUB555WqedrVkA7uG/NMJJPSaRZPMyFUAQQxVtVycF
7Jh4k06qqfq1KoZPgi5TxasC1z03xaNVXC/J6Rb9Xb/Eh+BWgYnmj92wqleRbXcw
qdOItOesjyp1QyyZ2sbUI3a81Pjp6odQXiz6oXljIMgBAmV5S3zJ97wbgGNqsHzb
syvY0BDyvt5Yfp7sZfZJo7sqjlycm5wf4D9jUlNBnt8nJ/ZY27URTEPZrsu+8FUy
8ZsNsqzWaT2cYoHtLv00hWAjecSGGYWE4FJTm65GDjNsRx6xAW/AOX3IepmzFW5l
mbE2P7DgcU/u8bpekzxwPpk8ShT7OAOz/JSBD4hJ/2ye8SpwVwCCb9y/wSfUgCvV
tZiXcR+Q8MPeCe8sgbsYRHmRugVjbuBNZGFmdS5uMcOIFbmUBgmEzCtQF9lwcjvd
DDZgfl29ymwCJXqzU8fBkO+xSpPuZO3p01371MMhfgS/JuLTzEv6ABd/rxb9hi5L
IHDFUM3gaiAE2D+04a9LKQeWUIHYaeuOB9Vmrzz+knjseoYdtEo24N1u8YMIde2S
/jpvgcVZYKunWQuF8JxNasZl02Gh88ZTmiCfo7yQbF1+xiAU+o9rKb1XFukf+A/n
NIMAw7POJQmtUTzomE0hr5mYtQ9xU9uYihU+BDu13LqSQ3e8yoq5eLnwXTTv6Fci
o3to9lNOkAhh3i3R/+SyRCvu1VZ6KD4F8HExAqt+cmXu69hWAg3vfNWBzPYGZP/4
z5y9tMuXSYP2ROONaRhULernzPnrS8++z2QKdZqvfXjjbZueisaX+HiZSXssizG9
R1id0dKmk18xbYcGQeFBJeJHnpAlNnp6JMaU4SvaOueqSVh0rSNt3q+hMQmOciBF
Af13VQHxOZzoaiVsOT6p/aEhNj11EdnPPXN5JwPGIzAFQJEXG0szWskzCu8c33BA
tGxnAtdhmIshZush6D07M6rD8At/o+02aRSTWNNqcREq5XMNbnLyAxwcOXUwyQgQ
rx/HmDdfhrlTwLUC+fRcVTOd+RWjjSoO0kO4yN75yII83SbE8l848BysDKGC+kvQ
MlItZ+0s+in0/euK28bknGX/rNqLeEmMovVKbyRPcUYJVMMh+hz5VgWvMffP7yhT
rf5JC9din4bTrrrF7fDtPDqxCBrVajXY0bO8ldpFm5E1zECZ7LHTUNrjxqWOGcID
msRQCN+U8yghcAcxFc+m5h9sqExWzLE/vsz/WDy4X+p0+jsrCz9+1A8G6LadGIDE
8xTPh6sAPhE7evUwZ9qYBTrVJz8EWpTQBrbs/VweXxEXowvzmwUPIjYGqvqIhDPG
AYxTH0qtUUlR1tJlw2/LGNXDSiLoBA3X1SWALTZ09q6G8lm89WRE6QJBBrcgZdhZ
wLh4LeGO2BEnf0fcmifVeJocWfAT9ybw34V3tsX1IrU5BeZYGfzaEcAPTZpBDp4P
HMD4g7GHHRUwNFjoOxyx6oCw78X38M0tt22Ib+/7Yva8B0cPe9bsHOW3Xy9e6HIz
0AeCRTB6JArZ+5lJRbzGbJHNyeArs2Wp7J4VdZZuqgWfS7983hLMst6TIDHnkcWG
8WWcIMd9kq6LlTP/syIxH4MPnG8poHMRfWlCf2AnYoHk2tjkftSKAzT14LnVOJjc
NIxIu1TdCw0Gk/JQGqvnOZSOa3Kwy/MgyT+r7zg2YVDjX0t567A/ogb1btc31cm7
05MS/0VFTkmoIEBAKRKwSsR9KTmYRd8vS55JCRy+x5xYy+te/BCA1hqFXhOfkl8E
NQ4ZM0HjUHXRq0avLNBilEzNX4H+MoauMnojtI8cW4RLUec8FF7I69p8G1gePwsC
fdajbwhhOb2y0YCvL8REn6BBNxdbmNstdQa5nZjlE5UM3IIv7EW0VHWgt+sSHaMP
i2nJZUacMpI6F//tNy6Z6sozR8XX24VewJ4PnY2TXtd0Gx8JwmkSvNscKrmVqVj4
1mKKwq9SHKc2+JkqelK+z3icunCutWbVr1aFtvKbHPZUBbms40+y+mogrD/okd9R
IHaVgL6JIwJEAO9NAvYN65Sowdc4CfdjbyuwzXYlvmbP3qNXGoihT4Cq4bIRWa0o
v/oEcMcvLytsxI4AqP3oDqiZCVMTLel1BM7bpM5BRwtJfuE9oFfRqtqfQ53dFzue
Z2wSvEsRFA+a3OoHgNTO1KIvE3iFC4gYZqMFXxjVrKOplU7xDPBwZtIR650Sx4UT
y++WWATeW5oCWBPx7FW9PEEHsVLYwT2VJk6L5/byHXt9HjUHr5jrpDbzd5TAv3uG
7biMnEe3PFDAly+wSaBzA/5c4l1TrgsO9yFrZS3zlRxYo8bKUmLuCR+ztRSxrBvA
5mmKDlwo9GFtkjbrNia0ryiXUbkLVjROuleRW3L3PrUSUHXnOLpbKkXASC0cs6ym
Wo2IpPdprdZiHOg/HgEePCj3D2XbevaT9/gL364QJrtT4+jduwKs0WTEcBgJMbP0
7qA+d8veIxiA6giVNnQmGDOum4f4euQadqbCgZ4vQ0qa0pGJWs6Vkbb9EOoMMj4S
oHTM2jFErunxtbVHFNnZh9prv5DUs3MQulf/v3ezzwod2C92sortcc1CroGEWyE9
/a35nhvxs4eLlufjSUlWNvIBpIc88PkRwMUrGzviMqFRK9rtZm1E9mbU7bLHhxto
Cy/yoGrxoFCIT14WCh/V+w9XUGc3UlX/gNOAiWE9+gPn4Jl6o5ewxwrxUTrwyCQD
0VcXnuIAwNPjiu076q0UVDgPFWqYIHHT8+SY3dQC5KTQSFZP5etFj3G2srs9u2dy
aN4f2NF8ypdbJLCsKZ2crcF9ICjxoPSIYHmIiiQOwdiE/saPeXA4FC3cNF+9WQuG
CHH4ThmLA5SmhyScRiaeAeyrY1FUIb56P/nlfnVRLigFrmSWd+r/JLj3I497HZpZ
36XBl+FleE6NaOriut4XBnGll7NDHEQDypzpv33kmr6A536KUta7DBKSxnID4syj
bIBA1bVaB2VUPoPaJ9WSUlEMfgrnT/KC6f1dV0ZirauqF1NGZ4CEtRNBx8Q84Dij
LQAX8RESBnwrmcbtiGdcoFpzSTHY1wfvBRziHret6RAdRqIqkxsp64F1czlhEH9Y
/OHcVBxA+QBYUJmautvZWf4bsKa7W9o5JpzaQQAFFJ9PmHbhZVZOZ0g/spB0ILwm
UGU03fybblqosed8p4BL0pDW5v8Uylxx23tFYU7h2rn//FFplv5OeX77Vn/zIryW
zQTGZc3HnSDBIrdTVHSn5ATH2/uDnHUxNjg0M9wzKbVhfYl6fntJyDpWYgwcuYB2
kP6MIgyJ3ebZRaVOB6PaQZvbNG+CvRa1lMZMykamnlh/EwzvzlhONmEAjhIeaM8T
i9uaTA8ukAfnYov/WW++uZ+voWyOBBwwsf7U/J25Q/pJxxqF/Vc0ez+VukzydMSN
1lfJX7NKOj7iGPJlj4TKBICJUWqRSaXyitEUDCzUjDMiCjTds4bG+Na+QtD+kQSe
0VXDbxjJ8ocF2EMAXjYfPl9XGzZzXH6UEL6nQrXaamarX6xOXvGH6X5sLHzTcXng
eNr5jpBTEXB/Z0cc93mytzraLiVQyLIXaT91xawUCgfM/oixOIarXXsJP/wQEthl
x39UyXox19wOZafwE0REbOGDdQQMqd1GOPBgH8tX1RyE7T0mgWvh9B/rPDgby0XI
gynXAWhO7ivEvhrbo+HqhMLbj0ObVkjlrMjE1/K08G3f2WST+izCxP6GcNedymY2
Bg0aXAJpw4anysEqci2bVcIJCxQZg8aoCeSSjHd9BA6h1Ch+7grtfOnbXtZmRhJb
MTx3Ln1loUZlQcHoX491/64WyXsBiLtkCVvl1T8xa5k2rOv4jfkP7EM1/Vtwgqrf
0HaAFQPgXlouyy2DM5AneobbU4lk/kfz5kuyyiesiByxymBVq7SZGYlgdDYy1Fc7
MidGOgCq1KRDGvtMwFjv9dMXlG/SQBAV/46p9BHVow2XvpUg8ldL8lywUPHVpeIm
b/HVnAT3Hf/N6tKCwbL65/9eMFpk22JyQeL9p4NnCIRTSTdfAYu9M5KdeMzu7eFl
qMdZBv8/uhOqj8hKAnqzR1K+mu3YiDcUELNd5qQd65xdxmmw7wllCoph+GOYe5ii
y0SF0Z2fEuA+ZoDLQjdezYm+1j220CIWidqYL4iwZMOepPZJ+LAen4XXg+MsYaaU
PgSzHTv3ZlT7iB3SJlsQXhGHRmtR9zlwHGxqi6hzdoiUbS00kTsUKOxLEsx5ObVB
TxeESKFpMA4ogkC86tJzgl0+DLGcYzdk/DLDXQKf/bPdKgKgBYNED2IcJEjEnj4I
3Hw3akXrVwLcv3dVxuK0eXzt5AcSAyfcH47Q/eIvkK0xbNlBLNmQqc7+lzwPKr0O
1yC5eCylz//V9oYw4MYSdoBDnvUBpgOfJSfcR0lMB7rZTndDH3jI1Zw+AdZUy5gb
M5TVrClmw+C9zl358q5YBxehlc4Pcbst5s6KP+35zNpO5ASKwS2x9WVUMOz426FO
KX8UgUFfOYQwysz/5MdT3EWXzogpF3CZVGNWY3LEmSG6E5JbGwEs3H3zE2kNTs6S
BwyodzSTl09am24ZWkirFA4WiPcZSrnaSxiMwmLmQ7YmNE0lzYs9rTioUWgOzVtD
/PSAwCQHQ8tpFApklEMSATac6j+eslLLLf6ZruuqfqAYPDE+/Sd+CBeGpM3+YeM3
J3XSw8StLLpzSsCKyhS9RAoetlzZkalX1bRlHx9z/R4lei2Rf88pVh0d6e6py4ns
60uGMQCA5X5UPe4QASu9AVLJyYit/sMZTh1cw0T1MhoVNuLbRzy6o1QbkacSEocD
Lg18ygSct7XZAoaATQX9fgk/5uki/JsEaSWgUSXABxFj6mZ2D64HtkUbivKUQlXh
nljmAgCBvbdhVn/VfWrocQ04KhQO4nCmjg26yggKqPWXPxKJUdA/oGmmX9xfqwB8
4xiMusfb0CypA4c9aUYd8LHwizqsk9n6rRbVFlqFdK/YHtdmqg1bDhsPfhsqmdvT
/Jl1bpMpGF3++mbwxfhiVSsq01XvtMSYFmmGBksY1r6G3oiRyDMkzqxDV5e3kCwM
cdO2sLU3JfTJa2lwOV6FXG9/R8UIjh9PqSEgF+cQoJLlVz6+zpQkGDseMqeQQ4OJ
ADdKuZEDwss70X8H6G48sIFZ0GKkr57r24TK5vdCHm3PVSqv2M+Emc+tNz/TKXzE
r+TtlqxxkmZnBK1DCsaxsSqcOH/XjAPeAXw3RGRdli2vRyLS7BNESmisDGVm4jjl
piBpQVDbQgCaYbLZ6aa/Aj8cd5YaKU4dppNJs12RKot8kMFPcRMKEkUuQxMMEhgm
Ftg8942UE+iDrO6swm2A4ib74A+WKWKfTWZv2Iyg1wpyLGn51/W4iqYtPjuaRro/
yS/bTsPNfJfLzc5GFPVB9YBinwN6ImTjiljUsxoGA3QjTgIvF5QfeYQJfyms7txO
L6zfnvzO9rNQGVO6GZEVfpRZhQGcu24Zc9/Ni1rS2JJIKF7fUNjv4AKqT19Gh+MX
9Yh5GyGth+CWMSGdA1PcfdKMx6afMZRlSl8BudDbwbfyEh1zobFrwBgXqyNuVZzx
2vZID21B1N/zNRTUUDnyzd2B1rJLLyw460gyCV7goFHL/dYMwfZ1mnsaivc5k4Ym
Yd2bXsLrToQWvQnCt0z0L8HWbVSCwvS36B2Ia15Ijz38h0d4sLBp1ucTY4daAXZ0
rrRmBVGVK6GgnTqwAGJ07w9e/R2/v8GZvOjW0Ap2GLLH1kJ5IQAbb+JhgHFBXBcD
wpteG3nmBDbcTg9qktAWx3IiwTG4aTwvv0pFitvTNqbTAKJHnR5TzgVCynFXyj5f
pSCCCfyOvjLA2SmCWWcm5vTIaZhM6eX7dO2/b1G4B96/5+VabiWzjfsQElBMC+4/
SbE4kPiDT4lDHSo9LHTZLQNyFERWexZOcQuU1JKvdV1pj/ssEs4V/fOLFfvPWEvF
RjYKQJ3Cs92wRzdye642imWnRHfbEBZ57bUGc8/b8OW4ErhlT62zkIseOiC68X0E
womSqPhY6K7+38xG/kaPJXQIfV9SPyJJurFu+u0EORlk8mPVuWUrvqlrxtl6WIf6
15o8ldUMydg3O/chB6oEKLmJ2NzbfjrMSKAIPtXCpD3W5goL9zxYU5DSTgMJ5ko/
st9NisQtv+SAkZx3rYDfmX8lOU/BWHjExBpjERAJkXo+LC5zuiYIQWHIwAK7t74P
skBnYAzvGv7Ucj56nfGUS16EqMsLIFpj6nRyuzTunaL41MaqM49xiWbvi3s5U6i5
z7QXCWmGinnxrecMbM5nvoWm8iHQrOvJupGJmhzDPcZ2WQ91W/IQmiGAz7IeFEea
vcm0VRovtlxI+gHYKUHSIk2OOAvdwtnvhUSDucqBQWVXJMFe+TMWUAIMHsx8kVVl
I6eLvhzaYFwssWMkyOZrNbGzQysjFqZ4TFRZbNLCx0+B1WwEfEb1r9t+KDALguYx
4K7STFDWF3W+F/vfCrny1CYDbmVlopbEqRnrG82W38ZB8rAZhidcaqkvp+eMZm63
7Yk1/BM9r4EuYPnVT9xUYu5VdINsNeNFLb4BWLTybpdIq0uNTFAh/AQNqlpNJ4Kh
sy7RIv5UWGfbb99NEuc1O2Zq0t0q8HiRdjw3kYZTljOAGPLJKNOgaPJpnHkELO8s
BKbMwJ0ZN6HrK6eNv3GRrqVvwHELuXbdUuw5UVUgLext58EOMNkVvThAPjy2nZm8
zNEdKvQwNTCS1iePdcUAE0jf8Q6gLBf5RXnVgwNOXYROyC9Cxibw36zfzDvaKmJy
wbR5auls9FpSaHgmHHo1KA46E7v4gkfkNbN6Xc07iC6lLhCs/C57QuqXwqcF9sKD
KPkIE3XGE2wFrhkSODlJDtoAzwVrlc0XH3A9sIxKN6X+Rt8bTMAIVJOXX2TSfVrV
A/V4CHMN4/SP48X9yzIb4crciioQEc8RlyMhbo37ZNWT0edBrd++yq4Nhe0hv/XA
iRzm+wvuMVZhtHbU2NerU8sjUEQdON0ONGth0IGgARxikJEeA+20g2q/BDIpK2ji
/4+/fOivWJiMpeoMZNwDV8UrSK4ESoFpY/fAoTqI7BOSljfDtSFIHiurHNw82z3K
o82h9L6poUGyER4ZDdEauZaootXh7zPHe/uxEX4MZDZcqHmac4/z8X1wta9TpDXF
AevGpTspGpJPSKrs7DDbYaS/hbtt02Hnt55yhqO+aDwNFdyUWFnSMjWqpO7KlNcP
QTsu8YMX5aHnxf3BUS9TY5oRQGVafYIazsNNA2W3HZPZQWRoFs0AlyOKfcuwsoRR
Gz7GLlPcm0AWpUaCzn2HfQZVglDS6FiInVDkTIBxHHnBl+MAorxbUTCAoo3++Xgz
JZ6FZyA3qEzT6emUoz9aXFWTgb5gGz8MfWhuwZ0xvLROF/y+VEFZ+9wp5dRg5X1f
ovWZ4km5HtUBynC1W7dwOVq0r96nHL1XTdGa4UvZaX/tj9tKecm8TmnbzzxpfNoe
gZujtureaI9dXfsFkX8kZ3WNE6h79JiEDXy1Z6DSb1kC5SMDZUw13j9tTM1CSYfh
UVuqeZAjIcwp1EgvKGIOMkA2eFAuZqRkX3LcMOPfP8YaoY1ouGto4ttt2v7CZSHt
lDXiAl4zYI0E0YckFQYXiPkVYzx5X79SvCgz6D+YvdQhZDC+lzDMTPwD+PLZgQ3E
FG32E6ZDxf2HNXaXuRV6+JwqF/8OhfoNgVK+zsP339d5zkbBvO/KnDylsbBGhs91
+XTIMxbAPMHVV/a+DMYum1MyTq+lLIu7xBM9rp22o5yebhElJjoUgaPwWimhWWBZ
wq+RRHyCvd4AHBZBeIf9//aMThEvwQSJbhw+nJP6KPgdQJYxeOKQGJke1gHfRVcr
Gd3RW7iukdk8Ua/iLYAlL8uAH+8tlWf8ihcluPO0yMtmcvwV1K/HbshSCxOo0H6U
BlT+/M+MzcGfKgj8NJZ/VPBLlp+JY4ilZS5mO1QPmHEva4TWzkRcweTT8uD9YR6R
uKDCUHCK+MFCB428V9hllSZE54z4mqhyUGNos1AO4lVJrDlIMI7C75ZSoEyFiik4
JVq8hWJ5xZB55ShWCfPn7dqmOj1IcgRYIijyTL8FJglDwbNjF8fzR2b5E4KM35s2
4KYkai30R0j6+7XoD0FzjG5v1CQZ0C2etPrMawyXl7asdqvGQprYI4DExHn6J2YE
8kfco/NQHQDqdi2z8Ui94fL7wIPCowH6OZyQHkdNiW9QlKh9gz3NYxlE5teW8cRR
dM4q3dKt9daOw3KRu3g6z2w4gQ3Cx3GkwjgJVLhfundtRXTugir9LZv1Pnd86t4D
w8JaCgnhj3XKEzgZdeJLpLWO3bl9bYBiL79OPfXvfvzXENkaVT+7n7S41e5FCE6k
ExLpWIE0Qrtl4q4aOFmlSiUD8T4RxEDmk94ccbFKIsVfp3Y34/3PuZa2lt0ym5BV
yhuhhmgBAx+eGBooNJdwkaLGOg0X4gAx77XTMf/JDkP2XiX3pj4unEcV3sEoiAnG
lMLGeSD3wfVqUAONWbgaNpKcw+gaBXxgP2X4yw4j132eFxIptm2Hv0nrG2ltfO+8
c0EJascl7AtbVacFMJO3QCmmcYL4k9U5DIryIikNLFe7WW5XcjXOkmi5M6ZcK/hk
ZtMw3od/BNoeuCVOoSbsFT36n+yFjYAO2mjmtmK+D4TMO6Nb6ZrRYjo0lwrfmQYm
ZRPM7KEmwoEHuhBYD0AFQmd6Hiu/IELF4mOqJZnUT4kPWiSrjoNXnz4A3gyOmuIB
L4WmDJ+ZVTnBxyUOrGHChFwwIRVTPH1O3b3xd5hvQvuuBxRFTZMSHs094YF1LVFw
q+aAi9RSb6rJ7CU0xaNqV91y8ZweZ1VP1t0tJZvtQbrF/zVWQPNx3XxcWnME1NYW
SuBbJPoi7qj28pTnPo4uFmfpiRZzihW4jpKVmB4lInpYhJW9A9SCEN8UytpMQS4L
A4kB/ZcCDIFjfdG+mztc3jO6D7SBz4D0LThZbdzPC74/TLR2a0YqQ8Jw+EnQpA1y
4KwzDObRs2Y4R2xkMPjma6DulUE9simUFWv3zVQCNxd6xO7GtSKXxWTDRd3zkABv
Ocg8bjdJGXV24YnCZuOGIpiZqblM1jO91YTrHOrrKm40IpEtcKTgpRkLRhmcDCk9
cLqANAxI67fVC/3TkkcuQeznMN8XV9e5eL6oXrIFeCFhDf4VK7vKE6yvsbLLPjKu
irdgeHEqy3PpR+B5leolgUHG8ZdNXC1cnBDMMc82ryLvUN2Kh5j6m9lqexKHeOBV
tqaDirYV/Z0RyLbyZPRXMBlrW+M1cqHu/hKhH4Bysfr85ESm/MBKLZPq94H6DUiB
Si2V7O6SEnY+eiYc3QslwCgZ0jOs0HCv8kwqZgm2oMH4pq0PNtHj2DrUOUthtDBV
fChM3HNtBWUKcyTdpwlvDnNf/+hgwLzZCk9s4OiMgZ3wqm6hvdPLfXF0navbvuYw
aN5sJTP980dyntOn2GtWzxZFyFnZTKUc89WKUxAIiXThRd50bJdmfvamedUctQm+
4grWvkHJL8dQWZDcjAdPhNrirNfzGdVxvdKdj4LI86PMNQZkusvH95tMbi67wJXJ
R2tMkIzRe9XgsU9sEOtwdyPZi0yTg4/kSFFfqEEtvqKttaGj18v33ZIXQpzHen6N
YcBGh7kqZdrQNRPwlaXF2++Fbf6iB+SWQPicXQGDA3dnC7DRj3Qj6H6O3pgeZC9Q
rP+gnedUAXoya3I5KCyfuWa1rEbrceVIA5IGsbu6/3F7z2N4uxqrOgCA2FVUNQdO
zLXv6u+NnXIMADCgWS3XcsoUA9wBWBa/NQZWz5Nr1myehZFOuoU08zDBaVHBA//W
rhRGMby/DKcbIz3SKNJ5rJBpqki9dkTPmJUQH4unOIk7OXUst9gJEJMWkQMpBa16
Sj9ZsBz01Y+R+oGPwxDffK1vRrVpj/aUMwj+piIcobF2ySIw7Ns4iE8fW9TTR2pk
WdKLAZsYsxS1akFrttLQY5H4p4c1VLfIgdsHc4nQDe4d+wntTasJnawXufK5hSEw
wNXkom/OthaqwxdGN4b5IktvdZ2yDsPIBuoeEQo2mfmP549BxAbkhT03JDQ2BviF
HObUwsrK+ktD79rohIdrzsvCMT7niOVGILRFcl6k5Y+HmUUdPGlK8vALZ+PoLrgk
bIqwMbVcu0NFfroInv9mOASiOn6oRZ4+XHB5sGlmt7XKDCPeZevZok2be9LWjbY2
RkL7dJ17xGG9ByhOp65oU7MUi1cccz/iohkGq6r0bfhf/yFp2Ety4mIozTacHvgU
38gADh2xSggpV3GnOGCyw3hHrgfBNfmAZyA4xQD2JaRAP5wZ3qsBu0j0U9Za5oDv
iMmMu12KQBXYIZNf/IMSVIs9tBqOlsjIxA9OSW1tsW0puBu9PPs2TXsywXFd/hH3
wCAHBrsPhaM2hB8v6oU11CoGVc/7Ot8CCMrlFU7vVzR+uyweydIHW5Ihvl3zud/m
TzPJXbGRPAY7tqn70sbyFOKF1NyAiMJvOB7Pg16TsN89S2A+528veovklkX1gfT1
vQ8oKJ7Wx8SiaaKA51yLVy4QsdxRXwf+1LFTMBClUpx8/C7ziZtLSTJPGJF7fvpG
S77pVPF89InCC9Eyl21M8/rmcCMxWh15G7Xizx3yjMjxfz0CqWydZFgIXeBvbcIx
bdrw8mtCEP+CekZBLK9jwg+sg7NFF/kj9EzUeKj1YwFeihqg5aSiWFEk8ZLJDe7k
bJEq+7S3XZ7fGE4pFkrhad/3HsUhTFTdCESB09Vq0OfOeg+cUaNmbSnBm4PTSz9t
FjniyGo092MDUrlXykSxhsoeiTOEFQVDCmi++AYruO8+A9Yh8R7iT+moERKuiTS9
m5uHp199of4o/mN83sLOpUYVYoWLtts3yH4A/1qlXvr/YSh1NWiFSo6lW/6EnZY8
acNlZeHx+dQ1a0NAzoO+RVhqi9E4HI2rKjD4kRwTiZ5OkGZFzVgN/02v09E4ARWy
ZKWJmzTJo7Nc2TomVy+hT7pGkr8/1WgS3+Xer22OiDg8DTWNHVtkFM8CGYVldNx8
eGRSTP2jN279BQpZICgfBoRIvNL+J7AMrRSWsAMvAimoU3IDhRdv0Q8l+oCGX13Y
/3oBww1ii1t+V7L8pAEq2AyUlydu7BH1ARuYEUyn7TkjNFE2Mb8ifTpt52Ht4DQC
RCn6+uSf2bnKtIJKoDmjjnRduLDVbtzd3DOGuKEeqSUXK41Fm9EPpDj0Ex7BPyBt
oz8LgM6OAIu+Yn1LZXcZZPavhZ7may55shmE7KefccP2UlYfPKeOroWm81QBOysU
pa3Pfdy8aC5QgKXwVCWZtHnDL4sp6YESpXxmQEI/k0ssfoGoIf1TVdxaoZDee8IK
qZIlVYorqzoYmsOi4m1BoryKuBSgisf1NYZDTSTwgMDTwol5YzOYVanrOvhXLt+l
C6jBF8VUM6vJZg+FJpO2HqdHrLTK2zKZ7/tJ2URDWzUNHIyjSZRFvqoRJ1voCRQ5
TbvWnKs9Cc4qT3rDYmTDQTJFxdl1o+j9lZlvlVtZ4qBaEwyMFEuh7STS8t91b1RC
hr2Mar4HgwAzu5HzfUkheg3kB1UJlZsbh+ZZSB4bCHJ4k0cP3C0wRgCpBLkWdFdv
a1jGiolfrKkaHh1F/yAk69iigAIqwIXr2lhm6rrDw+lDN1m1AcuzGwkYiJ1FTMO0
w8eIRVtq46D45KSDM+zSVmW5cWA8QOhPMxNxQ5gO+ij9wNz8/8kYfXGGNTQQCuvv
EmOnp9UT/fNGVieJ3CT0T6IfTSX4YtiqTg9DX/sZw2XBxpUleUZw3zMtctOGNuBr
65pKZcXg22ycQ64QXy27KvtK2lDPFIjnsNRtL+pGjU2lwheHScQcWo5rwhgbibF5
GAOyjY1PQXsEtFj1Da1vt2M8wa5aoVyIlHdOWDnEQzXCnBQu2TLOO3YsU7aas7dR
7aH/hFUTD2Q/bYiOKpj8SItOz/3QSU523/8iDn2qPOlmF6ibqPwrwTK9F6gZ2s8s
sOoyU+xPg+NgphitsEyGrNx8x4Y51QLC7u2PbxKngFkGg2GLCfJpRvmpvcqP/Rwb
gCVv+nuI5VQGF+GVcbbMbt8jKfxL5kDz/xmaVQrM35ZAxktEF8DfZHEO0z1tnDji
mxJktoTEGzrsqtHyCyNKRCYkMf6tNEn+1KQY1EnIFjPCWZvtvSMWRA761xIyh8Pv
A2TrKZNlVqXRKys//uq8rZhLTt5ZL9hVRyP2IqxTS2vo8NjnnDGgiF3NuEGGrQGU
cyP2urh3U3Qx7nOFdiP09yEr0RthKQNb00p/cjqOxnOxzEJKgCkUcH24wA5X2evp
YZOLFebaIp+oTmg1UgGoqAi9cFPk5auNo/PzvvNiXddZzDmL3W7MnjVYcgk8fH/l
U32khHu2wNPAiMmMnjLBSS4Ng1YOFstzWj/9JgCrg1V8bKxndinUgaWxAugB0JOl
hvtf5FHqvEkb2BowCd2Zdb20pxMhK26cg/Fxc2DgdXHB5uEttkn4nH+aBjQnk6Ny
TSDYkNtSWxI9QkoKlx7nSPtTr+lgdmu9gohTVg1DcxxlQaAHD3kRYQNx2+eeGl+E
9YRFBmu2gFH2Q2RuqEy07h2Z4i8XUnA49gSJzKehCRjpLZFQK3EqB7QEHQQbiwrY
wGjep33kUkGRfgxpjDeANZpBINZ2N5iivMd+Fh4roBtKNzt5w5N4m9bz76Hlvqvx
sFTHynSpia181AlO/Z6vS1vrfBIoxdACmojhji2LWcDN3b1kf0fB7GdEVM7Ckkda
srejhPXcGLFn8OLyBGYaY/g/6aGBjN3L4f5htVFl/CkPqpF9BNKgmiAf3/Il5bBq
WTwpGQrsWWffHCCXOO49bItz4B4uqZfOm2TTDSj+V+KpHrMHrceqGDgev+5ShgAC
qI2fcS3/Jq16XTExfUG5+l2qY99VVEENueMHPvDj21VVfTh6lBoprEH1LkImr0r/
vUVjKNQXfsLTj9Kpu2UsdEvaVQ6VAD4ze4M3uwSI0dNUq+cG75hL5fwgmetpIc9L
Nu/HRu33mkkAIrQy6RnaheRRnf+3F9eC26l3Waj9Oianex6v9/wt+14LyNocNF6N
vAehIBm7DWqCSlh36MceURZZdBUlyBp+NQC8hm6Lcqe/lqwHXr5hvyqePDajjLoO
+xCGNgc29YyW2XNGX7FP/8Qyb8AQ4Jqr1J6MXs7kgD5y0wAvoUFFcRhI/TfItoRG
rMRGTpwLje3bIvkuV/FK66a3x/mecQbTJrnJBp7DqodNesZgWGSX3qCaZq2FiB+q
U7GYZeAoL4ZAfK7/NWlZTT/TJus2cn19qJyL/+DeWmmvPz0IxrSd5Y4IJLNshMUq
0A8M8TEr7FT4NfwGthgIBewGVDcQypOuKehVk+z9u2iDotPfK+L0uXGdC2ZcI0yV
/2Huc/wOhp3Tzj+if5YSRYv0IXU/1qO3E3T3wKYCfhSwSS/057DFV8aP8xodl9v2
bsjvKME78cmgBZWjwlUeUWUirBBE5F5vdgTWqZkJTqrsB0ERJMXgYM+i8OEkIiE4
g/hcp2vLWMPnAWwrQU1wa3xrMVsAsb9P5KvMMBuKowqSQFKoDmiFMuXj4+tCEpOO
PUGGOGHi9v4gP2OkHG5uXimymNjS4NSteKLVFZh9ck7ZuzYj9ojb+FnYWSO8Bfoj
6rJgKMq908G2KkbqlrH4walB4Q/k43+htMythtNYAu/+hq0S9IrbTb7whUqfxgN+
/xjCHAIC4+aFyzo2f4nZSAC1vNKZtB7gXB12jcY6dd+B59kFUF/u9lGznJMaAorv
fY2gdUGm4fbRcWniiu4zEjps06gIf0ZEwJPySwG9D1hIHVErvJcxi4g6jotJUFJr
nbGR1F5zpfPZCFUHTG9VADZvkYOyf/E5vqb62PW2aqCV1yG/4d34qwx5/Z7Cs51n
9CqRp4WInWSR3l7yn9jrzSzFH6fXQryXtXPhBvxwQijH03Y8Pu620JOdyrlI69vp
kwh/aMAepyOQVgbmKx1wCWGWRp57ZgINfYl9nZ2K9kW4lGqz+tZw+QlITZp5MZ73
idY+vAq6Y17plg/iFDzmSylbjylExW/3XCFYktYdVHn5x4o+cFWep8EfbUQKM9fE
Nj0XtanpMTwkf5qFdEUbfZYjc9zvRDqAuEyJm3DtRk5OypQD51s51hDgto1HcjE/
A7IeTPE6H1r0V3XCAk9JAjnVhCiMopymgYpIQ2UhJtzZAH86tUPS09J1qEjwe8qG
Th7S2GW+sCXP4WNdL1gcIkBifYSPTplPeQbQ9JnN+6/CWI5CekKnfkRocpC3ngv2
yITEPU5dAfqPdOEYt0cXLXBdo9Ob0+20AFQ58Fpub6HIWJzDITxQIL0f5776dlyj
tV88JdClfo6HFZXdHzR5hxyvF3XTLsPKyRUZlF4EyKdV96S3brP7fmUu+S6FuBzv
6LLiRsk001JeFm3Hswz9Uw8ef7ehLnphY1z3pRnLtoGTYvIjza5+VY/sLLVh6JSA
JXfjM6E7vuhDdz+muLugqRldMo6crREUPmOe+b9GeMuiNqiGgeVvk4FcSAzHiWdp
cYLFH8Mfe3cROnvc5YU39OVKqUsU440dnyhqn/4w0SGXZqy1mMDYwbmVahLkZosJ
ikhkhTq8iGxSLAb7xCqYdjPR08kHUXroKYJJ+yYlQE9PyyKJzPXNZifCCfGls7YK
JpfQ7OAcjh3Fxhem1LjzGEMQcodfJI7quC/A7JKUV2uTTYkmVYXg5285H7VAStW7
xSo/oM31L96fqIN8uk4ilbEFV3/tu6QNeqFtFIopre1lfWykXT+d1PZX2Def6JD1
a3KVWTpR5VPI91dGBRd00mkMFV30iXEMCIOk+mAwi7OSNbyVGlK8Iryl4q/4G+vE
Giu6vTPdt0hTM/6FE5rDaGQDH+ECuqjA3j7wm4FCdhJDThRlxzHN3tvTaQx9fmEl
s7Ixl7Aam7/yYJI+fD1S65ElyVrd6HGaughrNwcC8T/uJ7fPWoIKEzS+ygDXyJI1
qDY15UtejmvTcxzXZTIc5eVa2O+VA42vngi25WUOZglWh+scWFzLOEgzyoLsXTXc
59ID5cQMrrBJAAvAOtWVvofjWis9w3DfDbt71pJBXy3ZFUGZzOCHuLM55Ko/ItDO
klEMCFdUZt5EfWKFTO3fQ4ADu7jTzKYtk97RW5dwrMjYwhAQC20VuReoZZVYk7lW
9rrcfjUr41cfKRKD4ObTN+/zn9/OPeR8iwm4KSdhLHyS3rpEjYVhcjfIeik94SHc
F+sIpN7nDL19PWgYp725Rjb4VghkqskzelW3rLRhP21XifEdzNlSCY7biiaoNXF3
n5PJkkGHnuOW2SlSYHseXlSffula8wTbeem9W5Lt+tfTjuKQv4aLZfZfqwBhMWRc
NE3WcRa4adpjo7EpQGYjUbfvpFS4w0Lw9fr56J8cVGUO/1YVLJenP9av3dpLmgNl
Sf7RCSIxVd4r3JQdbdxsckCIyT3LuM8nU+nU2II8wt2V1xj5zhvimerq5aLTJ0Kf
LCxnTB2G2DKGY06bcSQf6C/l4SSDS4WQncN1Eqtz4s2LMQiSQxfvD4KFUqIah1Ic
MN0prPMpvjAhBCFUMazofoSFuIUGW7F3VXWXXtlP4fVlqRYpyTS9pU+d9ds0R4ut
mQvaqyH08ajsZ38f+RbAcTvwv6pRkWw2zd68nMitS9oq6zMGPofHhxY0LmbU313a
OwTx8OI60gSPH4M+Is+FyGhBtXziHyWw14JvEVq5l0SptP2IGPbhWEu765oyhDi1
QTp6EmMjA5x8G+l/CucaQPp4eYchEvdIe9eRFOcjPLFF7u0lHrl8Qa/lzT6W5LbI
4iKBOGwyxTMQzrH0OnkqoYtSsyj2gjbqDLoJU8ITBBCcxoDFrzbHGfR1mrmI5574
12Jtly5r+ScrLrPnhdfC4goh4kGP/r/P1jSyLfhVG+JOwacoCTuLATBQT/cb+OEf
JBcxDTs/FvGbHgMat3C6Py/yE3DxX9HxZ3TqiSIA6yzhOPtZfCvradT2Z2h6JIsw
Q56MXntM2D5LQR9G0eU19ESwqlxtXj4pK0mdqcCZb/UEb5LyKI7I9yAP09J0O5zb
qBR67GCp4Dg0zs0BWr21Jub2IG3Gvu7UJj3S5l+msvWVzjmIzAXQ4psouzFXvh2d
UOTnpnxaV3N5lyfqM7JPFPhYNGuzzEGbq1ACiTI6SajS8B8mArrOcAI6KauuRWUf
euda6G274cv0M/XF2FdL0603ts41uOhZBs3cGIihiXkCUyohy0hkRn1qAXHPFLqa
KZ4+GjFVcSGcnUbWdR7FmoNMwJEoTxDp0yhNG/QOByWOWr9YbA+Q+B/xem5HmnCB
EF0q2wDbKyY146ptTHjsckf9KR3WkxgmVCNZom8t6X8PQ7Y+5bajeugG/rOdVezO
PUTwZWSyWDPTi4OpjnqiPakgauVeFFQE91a7yUCiIqS6vTsW4Q3BZM44Xcg9v6pN
IHb2m63oQXIC57Apq/TyfN6dkRScAJp9UOnCzMLxrP6IVxODdGiOtUaMvVqjeHaf
B3vAJMJYYHXXwW3CrBbTkHTqZDD6j7BZ74p6qf+y7RfN2N79cDcNODxH+jAoxC2/
zf7qbXeiZ0/Amgo4AOKXjZmGzkgOf/KvB5ZCLhdy76ZGkiXKoVsfajPtXT+FRrvG
e1gEOwYqtqCYIJ1A5iMw5kUi/wh3K0WMCGh4n6TpNnMoPSB4St5T/e4oRx+1KnPG
W0TFwOkHTUsWhIYl/3H2U94zjo9aZpxCAYO2TrmWTmH4hqmHdHHNbE5bpJFlHipN
B9zaS2erLGnmzJNYW0R78/vMr5dWZKs8m5Klq+XDytIyGs16u2OB5ud04cqjOur2
t01quMsspPgitxdVgqGibhADA/GGVJr6W9qqbSJ/EY3+SHcrnnKqnee3EbaLvnt5
pDzqSnQN7BFbY3fSxEMSwuGiRaIxVEBTFxLyjRrayy3J+oeK5fGC+/DeibkbjchP
LX60ejo3r9lBs+F0sPFiIV3bm8tmi0OaQ3ThzdyMVc+j3Oz81s9cEqyti5sXxFb0
49Yj6v3dNVlUD5lw0kNRuEzILt6GGj6fAFhsZhca+b7EGnzbFFtouUkOIwYIq6zc
YNYMy1YG8fLzD0TxXJqYZ7XrGsjkf0bx5Bvfrras8cAF1Y5eL3i45NAwSmT6pDxM
mxokbPy8HsrFEvMs0W5UUrvhKX1S+RNIOoY80GRt8NHsKg0sAmx9WfjPwWAXy2sw
+D0qmuqZeKOlVO9u4MtAKBCM735tARTSDAz25ccBTUI+y568RK4aQW1GE2jdTElH
+8+Cqa67bYEx+iLqHv3hmd71C9uKv4Lw/x6cRIaZR4WvS26VbizLEmzrqQL8o0UP
pPm99G0WyUnpSSyxuvBBkEI4Bv+FSKomkXr6j85G5hMYA19cBCTfLp9eh8SqKCfk
qoUBZXJ4yj+jV6QG498qyGSXSN8WgMwxwRsP7Bh5z6PmYgTEJYqOVzw9HfGw3Tt2
IYbUD7Cs710RaYYt6atMbfqGsIrkEwl9iSEyPlJQVp1/0DhPpqLbSLooH7kzouwb
cCqy1X8Bew+2/pMMw4qm2Yv0Zl/ydSntxJzGIOjLVOO/xEjV61MdDa1TD8gfRbOP
sWIXbeLu6kYsRAa+lWtb2CLbd9gdDRFY2KUFPUnpy1aRYIKLQYY3/wT/fla/6AUb
ybm6drQTRL6lD3bxhxMTzqyBrjb5QnTBy8QVvR8Ym+s/DDCTKqYKDtxb+P0BVrsM
tz09KzutI4GW/C/2ScvpgylEsiZumDITvwaLIuH78LqHyrL1JsOmbW8TZ17lbuXv
poXIPtxCEMYDRopQVuen6WpTrogcsUFmxrpQKKkus5s0Q3QGGmyLChA3FkL+QdUm
6WQnRzqRiaxf9B6GeoIBgBzpsN9UPLS2Lb/lCroNlF+FtahV7zi3HKLNNsWwvUNx
alVlAU6K9WLj7Eu4vkCL7c8baR79UK0e7VOD/ZCnl5Y+jQz5hyTvzSg5YgrCksXr
M1feSPUueXgHXntZskLgIxdbwn1C3ATL3goVcrxaQmLh/8+UwaqsBVI7KYnTZiYY
5c7BtF9vfeooB1am4VHAg00bTD6FBx1bGpDgH3JKYhN5nroEomGreyYdlpvdkZCz
sSJRdF7beLjX45b7paXnltY6ez4sa5aG5hsUyD8G9Sb5eNrAARvaWRsmQ/IWm+B3
+RWVTB+q9tY3W3/jF8ay+Qv7gTgNi384eysOMih1/QQ+o0pJKZI72jroDOadzk14
fVvRwnnp2p8W4XrGGTMFwuGC0nWEa4aiiuyiC8iQ92XQXj+BYdwzOrvevJewVKLj
SVuco8i77rkXLjpFCAdzxaUifsA87wtQJuG0dkJ+JflkvnopIgUIQ8Fb+HaThwEw
LAJMQrmowncvjGbfecIpok2Zlppx//c/DPAta39tfyqAjZB7KpWdPwX7jDsWpMaG
lE4I/ik9cSz5H1+YovWnUrIkfLIFVidaWuE5GPXrRx6tA4V3mbqSuiSMgvFkdOOo
1BgTc2YDU2z6k2vhir3DBEJzt4Igjfkz+KXUP1MGWwB55RRmcilB0D87ld+AdwAp
Fw0x3mzQlglQMK7UQQjQHT+cU2IfKKBe60W1oeeC0fnNHC/LEaFzy3fDXda5hqNw
FPcAGcoI6unMQ16HYPgc8VfKR4SJDu0h2irpN0Y8fZGLtYLuf8RFGak4IQn9BxCG
g22StxlTbtwKGKMK5KyIPk1KEjwTzZF40kX+H+Gh6M5Jf3dURjmGdQ775n53F18K
DadytSX2WJ4Er7KgJz0D1CXwDOlgiUTLJe6Ly+DMrGjfeGVq+GSdRp0ah5AQb6DD
lxz+mE06sXTNzp1dLKpDDZP5qiiIBNZK9kt0g2RPo4OJBxzKFQfPzMhTZqPhKUbO
aPLyk4GLlsWR7QiPMAo4gNeC8xGabGQuH0oYDZRIgWlSIF2Q4jtjFfLO17TKqF81
DmJHVDEkgUhb+ylg8CzvuWBjlvgfSzOvUTpOFdJip5JSkvDkJ+WBqh3pLx96FzPO
aBS7WJdoi++C3wI2zDwUY1b1AjBXp4DyQ6kT9+QbnZ/qa3lpsbrFOUCfNlqc6Atm
6hSlnfxX3N3W3PMEwLIK3VD0K3M9GCCcgjS+lmD6hpu9D1DnA1N8N7BBr86+BRB1
Ujq8K7treEQfIqAkaFlOpd5WpW4yZNhWIZYYASQe760QfX/ifcxzCyHaL2IquE/p
ekCPngqmx4FAHy+zzg4yodLFbr+wZcfufS+o5+pZ59QlCzMrvHxCOd5Jm/6AVzsB
j9Ggcbq4EMI6L37XkYAwBFvKVLXhrJexFJSe8Bk3pUemd9AAopfaxp3ujehmGjZy
Jv1OAXf51Cl6aR/h3NjLMF31Kwu26birZg7lhn58effeBLnS+5SxuNvIAPdu/R/y
LZDEg2vPApnxVDV1oUBY+OD4QTitg0fvrnqfeHA5DR6Pzz0az2viRv0WL6xiHiGU
0StrndqbXNQu0TAEuGYprynzA7rt8M5PqdLCojDwE9DVBrSPFydJL4gcvyY3etWI
c96TUJ8pVDoVBGzHr8Z21dS6fQdm5/5sY0fkTFYh9zLVkOX5irpH/aUyqMNsn0ww
1qBgzfqZDgxWGiI/0G3SGG1irZx38sMlMw0QX7AugS9lu9oscEJhz2ZWJpjpvFNu
pZve1fC0OgwUbXLQc4uGn9d3U5yQwTuGPN+c384djIx+ZVy1IuzQ3VKG2g9D9jOt
vCfdQTauE5e6S+NHMMfgoVY4ZweMJ65Eu/spG6wzDtTnz3n5F8qyH6++iPgqd98z
D93z3KocW6sktX6PrurG2ogs32Vn3Qvtz0o/VV+bucqN1nGTWSJByRvT33o+jEkx
ZzlJxs/e2d3rdnJfuOG91n05TvJ7a4pk2TkqBUWaK7ey37Huy3I5rQvIkZi/GZpb
8MEP1/1Skyw7dslhuUIhWEdFdBvsLVTglx5EJIsYzMGHq2DibRXO/ptxqEynZ2/x
/wx7URk/b4Hz4gtZPH1JNDXN+g1hfb2Jfsi6Mjrzjhm0glQs3sEaXyuLfIfhrJ6s
8Y+NhgLS7mN9sECKHMthDnK1Deo+OY92axNF3UdEtbfaBZ9mlwuUf+109gJUBURC
hJUEnTkVH601zTu54iZQu9F7xZeCgAZTDi+hhfJFPYUGiep9sJcKBLohLdDtHvO2
EafO1Cvn1aAX9EeoMDhG3SYqxfiCplhx71C2rZRU4Y4rRASfS2/gVGc7Um0ZYGxo
RhN7we19AOiFAL0cTrHlBq6h0ED42SaahFr+/bxRIJQT5c/3YY/lO9YJF7uVYLwH
H5GHQhduAjj51HKLuqor1ZJMlVel8QPt8HPEU4Q8Tfh+yNUpYs+/I5+lZCbGcWP0
3/rZiXc1jJji9gUTgnprbPOdBHNgC+XA9nmLrxe5n3j9hDXdrxl7AzAP6Zrgm9Eg
2ciiBxsVgA/VhNytHqnRrheSJpqBUxRuFewple77mlsz1MoAPcqVH1zRA7Uh7AGN
RoSw7sjojtU2fuHMRGkO9OQ5V0xE6mQbC3ES0GAYeyuqx+NLeYpJHHpAFCga+wL+
aBEAA/MCbM2UXe4Zfyb4J5KZ9eTwNpYegXzfK6A5+4WUTBMaMQNxdrr1XqSN+/YG
whmM7VH410CsrBFbYLjCz33xj3my5JJ3HHrfHOzrmJpDjRTa0kfba5A7KwB4N8np
j5EqFJ+RwLHmAnQAGP7IXPxA5s4wZXA8KXgv5Xdi5Vh28BdDtPOqB1Tzezdff0Ik
ZRnsRQag+2olBG7f7hwN3VKlhtQNUzFSpXyyuyO1m4pKX7TfDj1Jy5RJju7pReu1
zy/+56o5n9UbXVMIXBe6fXzXWnhRkDc5eQqlW8W+vCDhpWlc1TFyRZF9rrrqLXDA
Be8T+CI13DRjNQ61sE6zCHPXgYJViTn8VA973SnesMZ5Xx56NO/Ildy3T+lw6/FA
OBYsu6LsTcMmlVyKBrjm3cnM/43YjSDzvTyPLEMA7zpgG7XOLgg1t4ASXDEqxopZ
iqu6b3fcGyFkDLuDP/+jlZEYp3RClLv8TDs1vuDjB/Nr1lulS6IG4u1GsVCo19WJ
LqxcnTWfdhgjgaFOtKaVyBN26y/yJpllmUeK2skyazFRFaGQzPlqvIYzHBbDR9Am
wylkPS/eih64NZFKardxNENLtKOUqQzMT4ZOG9WbvtaVw9Bw8onhUW18SbgtH46W
JTLZPZGjtfnI8I2xcGhgzMo0sAv9QZWVli6LLiTqwfma/HCcUs8i5lt7BENM1+gW
b/iMHG8OTmA33KlMSTRoOkdzdn9Ggn6F7f+BeueUmi3vmxLHYTLuEAQdGZ0jMgBD
aY+lons8Bm/rZVVlCk5cosm4jpk46BXXMAui/LJFX9G08uvgfQ0LgPgtpnBqY2xC
Qcfby62e110vJxMM99NbFOqn4guFIHYdw3JEQ9G4v8a3CT16HCN0qNZ1gaNyN/2E
bWkgziQ0HBSIku9McXwsBz1+gMESMOJWM2gh/gEpmgGzPQ5PPFD7RrGZB+HQ/+EQ
+eWmK2xaDHqeuTbCqiIvYy8x9q/8RY5eODrhuOpFxwWMQpgWKn7+5tdKligpmXBB
z95DqsUvZy5xM0Qafq9mlI8xhyI+vsmnvjkfC1qAAVgBzmUUBzdXJ6VscTjyeP4P
1Qv+Ie2itWu1b4Y6eEOIaML/CrUrHIBM3Znc2PiHQQ9yt/TEXsk2xY4IH+B4MQ3L
RnrmTn7pyE0u8wuAvl4YA9te9lBkjJ13YjkNiFl6I9vukht4IQN6GOTeWskn0U8A
hfG7jvkHZwejzlfFUI+NVAUZ0X1FA4bKGWjDVSqbEtOZwLch0XKJbpV/fRSvfZTS
TBVM2u3Ol0MOdBRpTiOD03Ktg2+TsmXwJj4jxUB+qzsuFwjY1Wjdl6Kv2jLawrcq
/m4mxm7b8xK6layOAADcs9jTgFl01QWE55cZblbyPEkw2UOfMZAoeVPTRqOgPxWW
PzAjigz9tHlTwWe8wxtdLW+HQjvHF3aFrdQHg2EbPJewk+CHEK51MEW1alMDk+PP
usNFwIclFOmX8P4u+ORM5sY4J7Cr2d/UJ3Fk1e+rThYedq2ShkluRXM2mHCypWD2
nAkIVoTjGgltH7kD4pTsZfeRJl2zvyAXDn2rbaC+VIfNb4ZgW6e8YiNfiggYTvFJ
0zhfFNLSuVVJFR+xfpV2gc3vHvhM3i9a5MjFvwcOUZiPLq96RaO5tObjZNq3Ovdf
paja29irqux6UJqSAATksrixPl3ndMFW0JQ8bPZT+G6Qmu3fRrPQIN5cfqPzrsLL
7eB83movPIoRlHYXUvwjTUo0Gtzc8jXbywXyTHbEVbsG4eQwOghIX4sF/Y2JnUSH
DwNCGiewytN4DPcE9TzsH9GEGdkfSyjTlGqFlWv9mo/IwqjCNK6164aUXElPH+X7
O26uxIKSk4uUyBdaFMWuA8fza42FaanBQmZCe26EI+KbuU9d2MeheeA2cBqnTYwC
DmKTkX+N/pWjUTWqos9xM1OMB6U9eZkGXyXGeqa1yPJ0MdEeG1PL5GumniZe5KoN
OP0qfQyKUjsDsIbV/gTNa33eZkhP1SMv0v5PtTeFzUtk0jkC+sGt6FUGMRz6qzY6
0bcyYPSnEcLRrlhDapI3hSEpVST3arg5nu+mQ9oELJVLApQoT1imeBERL44EDS7z
TU1+q7qwX8px0HC7Q3/F+9lLcQMmZzjlGzml0n05cF2CxHP2Xngk85iqdJ0DE8Qv
7MDfbdCDv7SE2S/YgT9x47YnyA5TUulZzU5yzxfAB9AO9W5GSD/TfhnrAamvgAUr
Lyc3Yj953rmwu3u889b6r2ffgW02Y8fssZQr7wOgPclfHDhL5WvYseiZZnLdgX/Z
6lK/4XiAIwzcI4Sj7t6tHHsosmyTjqaPnLbDqA6aXn+Gj9q24h+hxX1muBnDNhLk
yFR/Zp1I2LdbOmW5uEdx4OKY6vsvs2EiUz82QLX9ItdflW3cPPrgniP3Ek9NB4mK
pN3D5er0zALLg0PU3fKH1eKGByRBg4+v1JpNRokCp+J7r3iuD28IeSNkmPuns2Ql
v1CCFy54BWNk6Zr28SxU1Wk2p6MaWVw/Y5ruYfIY98W49xQjBLXs5tld6MrwUDMD
Xr6taZxCDyyxazehsZM3p7DQoDqiLRJskAJP8kNn8+klLTHmp+/8Y/Fzovs2/F9C
OWMQ+COkDZIfyEkYwgD8vzAsfOE0KBqz92GZf5ZUhgk/ZshzOBbd6zHYROfB9r/2
S6Cxpj3cIj+q2sS4zxW7XJLYblxQVrGvet/0csRcLYBYAKPv/B9BGKZ3NatLd5Pg
x77DF9P8qV+PjN88O9ACPfASMlWD7siA6pefMA/SpVHJu/LE6PmPH0XIBRAoRgKg
H53V6YPAG1XZ48dGLSp5mjDR1MUdX2bQZGSXTI4S4NCy2CNGaGQ+UjDi45z+7rZ1
wWqsqrbTUORSfPGoskeMo+8rLdbBz5hdIlEmIh6yt7VzPaBmU0hxSRE7HKF3t+BI
Y0pcfPeYpJfy5nfyOUz+t4eE1Ms/WK+Dol/L8S+SZ9Bdg32tVXn6Y2VeZ+EZQkiQ
dTY8J0DTvSxLYHC6UYjuzC8XxooqiJT1sf0GRF44KzIuEDgsfcc2s/HnqkaOVx9v
kX/Mk0rTrPlqeNS+pWbDBbRVNwuB9dlnthtTA2PhtlGgWe+a64yIEdoMQDilhKdc
qviorugHU8a7n3C4uA5yizd7OqkRXW6W/JHyXI84GMZeJqmcwWBjNt2qGNl5lR5C
QqmtKcKoa/4djgRm9d4ugvEGt+9yWsxhg3v9uCnvnxS+bIRzGDMZMaX1LJQh77EA
U25a6eDTeNUls7+QQMkD08CuYUWFXpSxxaYk0bZBt53EECxcaT5ypHE0l1DYVcqj
MaL7aFpEaQrFFwJPGQixhBugWGPYaY5DML0sbVHLnKCJ3WIPi8ziaRfce7ufI/L3
vE68PVQK8l0ynWgdUApTdbJqnmG2hPOHVZzLmKsweNXtKc2Y7bYNQBde5HdVByuP
Y1QVNXV9jfd1xA0cum1l1KuN5KVaaLmXzL4DzXPgt+02bEhREBCnuGXUAVdw9H1T
fuYfR1TBi+vz54043oLWgW5NA6VKhixtZC/ZpGMTk1FYNsAG0hCdhxYdPrxJ9nmK
iJrdYLEe1mpGUrHVDC8LantsxiPNCcaheKimUMa8xtlxFKi03KKe0Uj35sLpnBdq
fJ1LctvW28E93co6nX/ONkfvomJjjkLzILE+2ZmxRMx120aZV81QHzhypAaldpRL
jzYUaDTx7oeYEJRTLivqNcW2uC9c5fNqOgWE6BPRUJFuc8fp7vcdGeBBMRqonwi8
T/M+FcMdduBo4lExsRlz06CZgTIbDVLyPCWAqDPYfm0w7qfTUuNleOdWExRESTTC
NLIJImeVZDtUUt1b5l1XkH4ALR9acpWALDlGUVfAJE7fQ9sahrw5E9qINSz+I4Ae
r236FSgpazd17wsDDJ1bJAKc305pjUUirocLGu51I1L3hC42hEQBzd5AN0Qd1WZa
zh9cr7pcJciAG6UbsU2IkixHDW7ct1zkLB69xjRmNKx9Wt3+YLSblKdCwq4RkByP
T2u8SFYaEuRpcNSflm4GJ0H0Fto1K3iaQEUdRMovZzYTDQlQGKxAiEPVYL1eBWLl
JQD8AvFyIVagBKIRSbK4ueq2BDFAz9vvaPJIid8Z9HWzzPRRs0x47EUK1BMHsR76
YxuKScF4ZL3wFlXzGvjk8aQIXdyTk3VmIbOM0Z/R6Y5BiloHlWJcaaLeeGLdccwd
kmfF9Onf0CEunHn8U+aaMoBnlVMJKMkYikq33J9BwhApeHA5775wZCubsfWvmqNB
MQsFNygBOfw1jYmuvE8ZwrzBZu+UuO1zdByili0RsulNuWZ1AYx/5ITPCr00Q0Pl
eBH/iGQa2kxvRPDUX41VZb+MEKrnpb4X3lxWNEYwVT5pppIQzAugu9gOUzDIr8o8
juLROcoUgGCVjuXq2ajqfNPBIrPtNwq213sQMGYXTTooVgNlasBGo+sKwmUtglhg
Zmm5E8QjuAsO7YP/UhOHHMd3Er6M7Pec4hVUge98+0SJfOXK38OFnomJlTpMezba
q71m9BsaVDm4qkhWWfX4Zh11nDC8oE675qhFUugnqWdJJA4vSwWoWKgU8d/gHsT/
e5jMVYDpr8saUwa43oRY/Ww9p81/SW9EuApgp+fo/2SWKkGO6mW7DJuOHbNE4H/n
oSRm/2+dIFKbBosUmdDMQ07zOldVoAzqkHcONa3T3hE10JAzy+FAPN1SRpa2gK+Y
4ktiLFIP89ftLnpz6128aibHjmyBHGGz5KjlvoIC/8SQnP51oa4pvrVPdoMkWfIa
TfTdiq6G/wB0V+MjU63LwI2sNrS/Ks+m8ve3JZE62zqEcbnP6Lp/69pKt9W3XT83
2WYesApDXP7NOSitEDZsgtuFBbiWw043iaQOcdSI3Q/sNyj/3lmlExYDG95gi2oi
ktMJDP8Ycog36/F3Pq1FzqfQBiCbPAZcHSI+Xd4UGasaObxHlh6DCxj/bjOkRgGX
txUV24YQL0/bR71hSzotC9cNrbYLEnH/kC78wY8GZxdpNS4y9UUQdIxujzRwnR6h
rlcIX5UzdPtuMIF9eiF1SA==
`protect end_protected