`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aMReDmrPskJscpWYThVKVItA5gecPPZO1R595p0GoIq1TSTG+UxXhmmUXc+VYHJ3
u/C3EW5qePLufxmXxmhmDnr9U8/cYC1zLfk44v/2OPb1TBrTsludEDQZdGNWeV9l
cPUMSIfZ0dHXN7L1M1E2XtgoTWQxf3VDHs7B7lU2y9Rdm/ibz0fWMow7op2nWdD8
gJ4QlNl3f9Oiotp1p8vz9RFzzZOF5gBBslZxcTF5+z4qO2W7+xLByngthWm+exIr
3Pzy8qyUo/m2DDwOz3VJSvSNm7RUq+0/yJNOOz3jr3j7ZyCj5OqT/jDAWjJSMH+i
2402Un+wDMOQxi21JLo3cA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="5R6K2aWI3OdbT2A+sz4o9+2XAInTqB1/cSw5W16RnA4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
Gm/2BIZF5/H5qen8uQizPH9RftTuEE9mgEOF0SqeOKegtP64CfvEUnIxj/ahmIpA
6xUR2v2l7E5duaLZh39Mc1GYsfqE91NCPU5whLaBPg0UuX4cgTkO4cYbW/7yvcrd
4wavUfwXEp2VSiN7EVxL8RcZTSMSI0Jr/aojiilFqVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="TEmQtJ1Dsm7TOzpJk/CeTSSFx/zKExk04H6I8sT4Meg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 29664 )
`protect data_block
nvPqn26PC4XWLLQG0Fq8XsMTlhB4evbpiwGjZroFFLgtNlE6bBjdtwWsB89WW4j7
jNfYbKN4sBv0hDeMH0AAR+8g+TCqoX7yLdIUd7aGwBUZJr6FdDs2wTUxRkXFYNTL
pZPBKDWpw8SI9CeQ0UEeISN7SA9JsEydseM1JA8qKKEA3Px5xNAH4RFUnlgetUIy
w8TlBBYnFngUGdGAyWqmTjwHULzW6s8fmCQrOpCX2YtyEHAcFfpPVjX6wol3L3O3
4NU+GsVNtA5Vig5Hi69W5OMzVdTz35aNrt6296y0Lst5IjMRFHt1IS+IvRT+HZEi
0MWqn+/tGIv5YUpQazK7BmVhG0Ge6EBXSO8PdVDHlPnpjQGo1KUE5RmWtQZbIavb
1K+GHIYT0kd2GZZKsOnW+iaG0rjYrdHIZ8Th9sjuzIIs57iCrS43Lt6/gH0KYxVG
ZBWaNKCOaCfeuGwWpOha5U1Bkvmjdg7lkPUubSbaaHwjBo98i98le+4+xwyFcxNr
FuFrAzyBkt2bj5aIUYJF5BhPsv1ELiIXUkR3lTnXDt3eUA3xeqRCuNaxz6q2Vdgj
i68lWlcu3yOXNfaQVnbarYYBNmr1NCQF1O9ND1HH2Fygq6ARwpNoXZGxjZV5GrN5
oSIysg0IjCF3U5AxF7hCzrsu23cFJi26jKG4x6ELXJ9XylXXOtAEdkv76iHeC6JR
zKydYx+vD8Pp86BJ1ttYwNzCCtFbZkb8ZMXbCOwuOWULXWqPd7fJa0gwKaW95lBa
mLjYwsK4ORhhPR2v7b+U21E02JiUT8JEOyxlX/tCLi4fZBB0Se2Wu3v0l2Z2Nr/x
SNl7/4x3RY1V/oL7wTHcP01yZHtq7NGEbRCAstsgWFXn3EwRLboRoPrL0CtSxIGi
7Vr2utInezVmRwFsIwLyGrn30Q1QxuJOWn9Ycve6teedMu4eWin6vClliWngxiia
6SSvMMbHE8Spghu72h/8k+zuxywmA8+e54HT51MMcJNEsGWwLHS+b812E0sHKwGU
+YzK3VLS9Oxa4if3Ci5nb+9H6RIExBxPBYuDt2TyUN8sQmuJ8DcrhIJ7KskZtJYM
QjDMO/snSS/BJz3c73wZsZC5uqq8vmaCj+YeKa7Sgu+NK/Pp8n1fb5mK0RgY4e9A
LOqUf78pohxwNQ3gIemloxlrndS6zZgYjbqZufxDefLxROUY+WGdM23UgzKJ1Vte
4S2Yhnv6StGE/OreOUtn5ONaLNU+gesWfLHAulsbm5nxqCH/Qkc/obFk9riHck/Y
VgeQ5zOm+YLKvMqqhhwwMK5QJxIzYGdGZktJEnUOx1AVrvV89qLn48/ZSifhTza6
QiRJJyTJabRNKJ0kjylFI5e6p/0zYhrDKtr/WD6WSJKQTBnZheiw3Exr8m6Paxmo
NfGQ01wOEJebNJECiQDHO5SmgKl0NPfDDgsNrFzxetSt2RonISWUqPOWwO2WhxxI
vjpdIXj/bh4+XwQnvXWVXsllX9P87FMckuPcDCa2yBhlA8jYkykUm3kLNA9LibLS
sI0dEmZQjpDCJ1mZekwvAYlIfJiXIxz9cjnC46of2JIZDa8b/uJ5mzvLPb4uk5LL
KdBVgEnHekJk74INDryfdD4cIdRR/o2+xRbYVgIn3KADEE1Q1wW6TJH2VazTM9Sz
FW+0yEb0TBn3fMkcYuVdiG7hMuWbzkrGEZwxKp6sJ+zEMwdoXLjcpXISbv0CJKpP
oQjZ0HUygdy5DSJXv2i7jyywIUqPNWYET1m6Bp/NU8djzE2Sfh/cv01BYZFwhvBV
h27dUPL0nK/r3Gb5PkAIHWF1qzM2SZYTvjlLPWAGKKMSEeeRZpYNd+Wh1B3VFwr8
Eec6p5ohc6pDJG+/Nik5YQj8SJ9HHBUtv8KQ4RCjLtMrZozvZb6YVAy/uNOxPaFU
/Dw92Na4JNtUMfWxadntWlPtnDjgeYO3CYcvZ997XiZfVStYBKBIsuAYYkdZg91i
da9n65nf+DP3tKRy08H+8V0rsVq0BXcT330XOLlSiWc+ZcSF+jXIR0D+W4ml2l/F
tscPVuuYJp6keSdY4RM3iApwGQw2NJYfOoJBbK6oTJHgxNnABpoqSNc9y3Lm0tNw
ljo+8XU+FaGBlRthxlV0p46WbIMrJ4Zp1kPJmvaCt6gf9N/4pDPqx5vpBB2ytl5Y
GOmHNqWtFdJDt1HHOqDENy+iyvXPk+xuCgftEXub70zmOorS4JsfXhOiTdESMk33
B9Kv3G5b+2XrPwanr/jWmmqtZzFwzW6x+fssP8QSJEF3WnHWF6rVIinRdnBOuBmK
JdNnTMQvKgIS69HWiKr5dMA7QpFoycM/+K21EyGJAHB+uuQiIao/wq+1gMK5+pZe
m7F8v2LIovixyiZDD/C+aJUThqAwqcVDIfEBZcYiZLlON5z+jkmatoSVfyiZNu5O
LCeq7/qfJGK078isBRfLmrTA5pjgHa1m5HG/M3lbhkIl0MQ1iP6O+4vvneWMIl9T
IYVO6s1TfKxfLW67laYdKDQhTgSfix2/3LzaF7pzymh2txcrHpIEDi0wYsy7ZZe/
g306wyzJ/2X5qHaI1r1qcSX9IVIhhTtIwLxRnRI+Mi7NUgOBS2bhtVN0g7l+ubQp
g5A4zFU7vb1km0OL8yI+woNHQewqadgP+qtO9JaElOkfiqx2xQpwVWAid0j64jIQ
2ZlJNsNq09CINbhqTM5qWI9ngAaDNdVvLYygj7BVrWtloMXb9RJF+XgdiMwwqoS9
kegG34zEyCP9wCwU0CE2VIoy9FrBfeNSainnBkJ93TLOIghT7HqI2FODcUrbIscc
5Vep9tdsa6F0c2wG10sRsfbfievfj9ou3fkEM4cLRQLyVnL5B+C31RSnQAtkejJI
ggKIPamjK0pZyDE/Ii04LgfvkkB1adEGaCTb3kE4g0J+xgddewmFeNk7w42ubdGv
stdD2CpqJCjkgzATp55NjO3th0yhlC+rBaVE3f+VWu07VRx3zde601cAo1VF3ngt
7XRnMi1yOzpaIHJB04U2oFeS06uKms5xOAt1JmuD/HFNQsEiiA/jE6TukCI2H5ei
qBPyCKMbQ7sy6/YH0p2j/n5XEHLQ35tRPH2JiplRcxM40ppOeWwIVwqndOd3UhT5
86eeE5x0ux4SfUVD10Ter1l6jYmglCFcr5G94iCdWg57tl+6aduCgmCNkM1e+UG6
cNtkvy/Dn9vVdMxMRE4nVUjCkiikqS3+FmiFC9DDM7RWEoWlj71yEdsHbWzPMv8e
IRE1HI2jmwjwpaKX4CBtwXjnVoMq8ceP1ViBlewDG9IvWsD3qgGErW1hDa+nCpvJ
8UtDjJh41JqRhQQVhCZ7ejyTYTvy81cpB8hffQ6QJs/+TppCoiD81Ih71wXrg/7f
sghwR3P/sFpTmrXuf+icYiemHlxTNbMqVnpFRXyLrEVmFNYRFEGV2BEIieeFDj8x
E1b7pddcc/R04raAVVCoEe/+vy6Oi9zTbyAtzB/Nv1+TG2m8cw/08QYx4lzDTGhP
9ObIOhDulyFyOBNE5d9NSjdMLgUgPbUORpqfjtveooBDlvxiRIUdWTjhAFCR2ayc
weo3yZylVVJ64XgUzfbR9bqf4aE2rKrKUR3XL7A4ohKhj3x90WtFImr+9nGI8PHW
oqsZeLSuUqM34EKBPqRTe/R1rcAr6qrw3quNyRON6KLgbuCyrCsFGsp1gv1/uPY6
wqw+mR0s1ceXcKyrmQSXnVCFO1fBD2LP6afhyQUZmLQgYm5EwIUf22aYPTvDk7oV
QPihAxomPuruyVINWgi0t/QaJfXY5PJPKUQ9YxT1gR0vbsb4XhLTy0GBTPtExcgi
NuqRUxg7osBhAsUQKy0bs9iqYMTmz5D/GMKghJJylffnRWlLV4TTP5d9U7fvYgVr
bJjEl2DnmpMqTkOtUOlzriOutcDzsVlV14QJjWq+hfsKUMkt+CQpli+oZMvo0OEP
WOd8LqB+ZKB2Mwh8fuTnCZqVfR6hspzuZELKf2UfQEApLF+HzaDfKJOaFP1lpeh+
xA/ZD54zUJ6F2w9Q0udb86b5kM0t/xCBghkx1/wDtqgiGhqFFfoB1ldHj0uxlGzl
F6XMNN0/SNVimfb9nu/LVqWwX89SlRO+M1GJ2LRY98Qqe8fTuZ94/mlHta/Y3PLv
COWv6Xh6AsEWawFWZaQhjQ+2mrAJ5NOyRFtMP4RrkwjQhRHM52fbKV9E7ntv6ubo
E7z34i2BiCxkbAorMUI4ezUINwXoF7H6WM4Nuvv2ugAVKHcV5j3PFx20AfCxWCqJ
yH76TaNWDhGBF5vBconffKUp1QYUKsea9kbwnkXiIlZx8HVj3q8EJir7rupDIUJc
uCKP6SFoYZmscZ2n6yYVwMM+RcGJS9M7elXF9fGzjXeLGEcqveRSowM0zZm9x0Tp
jc9+d3kt6IXJas9LV0WgXphr3niiceFcI/xiJFQPPMdNxscylZ+Meke0OT1XUc0c
e8mnXpQg0Rprtjq3edUK3JMz0fH2unINQacVTwgKUcfEbV4bPk7CVvttMPxG/5De
Jr3CXFWTSMEi7UuCWS9KgoXCjfwx38yoyUrXrUD2nn+SqmeXGdE3WiydM9TnPJ2/
pKF5LBwIJyJQvVxIkt++HGWDxxa209MNs+BJRuEQxE57ya5R6JoPm0rgLd9conGP
6SS3NXPgxJOEHemeIfPjyOL5JEkUROPt+eAoH2qz8nTTcLsU8c0eUvQ9iQHQ9e7Q
FjuC+WII15uzD/mlKKF8bS1zrAWaX1e+I75jwVfencoMVfELxN0U2GYNJHmeA247
tpaiTIG5Y3fWoiifqZFnl0p5hgK77LEMdNj+xMlu7di5mCSfw363OMjX+0mZreGT
2gum4/lccu74xMUbR37nsUuv5sYNqeXgsaQW5/Q3CgAO3Fu0Dq0nHqt1ODl7Dd05
7DQg4eH0CMDuJoMaumnFJAEKQvCJpclEx7+LpuddGqBwNyQSFzsIJ2Ii/myOXTdp
9PhjKMnguvf5khfqdOKtseWUQM6nDAA25KrbR83y8UOKrKXXbkj6QZPOO67fAw/X
KOJTzgi8TrP5QAwoEYJLPjdiU9AP87EguuPMq8j3hhp2OR6ednmidAYDZ27916sK
OnKrrRvbcNhjycmIBCl300m41IU2whNDPahtE369eDLgx36iJMbfXGomwt/iBh67
gGcwYKeowc6j7iHMRkb+4JUOB448vgTKNiT4ixogPvlDLSYSeeWtZDlL/pmTEHtH
wZrFCwo5Jo7t9AGFvz8yGUhFEWZYTL+AC9AD5lsjcfy2zhde0Lj8vYV0E0VeozF9
9QCs4jlHgC+U/ndOB0co527mSb/8/+lkj9U5V1KLKjtrH/rG3LX9kHbeQAyuAT+L
tgQ9b5ZYjNCrnlUNjqpZCcBr4tK2eaIs1CN2im01rl6s0jYfyHK/uR7+kPWmf0Ze
MYGWgefTZtmVIEzdwAWmaGDnOc1qj1rkPiRzhw9MzSCUXhCjRm/NvVOIkYwFCQRA
IJq9QM7M/35mpT4HwaJYktQJcBzPWJnAPMRHHQJPrNv1V6r/MINaYVERdRGvcQHl
RtYp/kfpLzhsvAesi4ilmZog6Eu4fKV7//doZXmnsYGYFwJfCJEbUbN5qceazhPV
LDACXgPfD/278tA7uM43ybskNQf45Ww8PW5hINZvNRufRIOFNdqZINlbh8zKgaOQ
p0Yv/Ql++qL+EdqdmrOCw92G/lMA/nQfsbSojHIrecCws7fJoBYk3ucNyr5z55i4
HzaXV7Y1TEXM9qJoShPvNjyGpbOvJZAH+EYATh0GbIKXDYuqRd/xTJkM3C8MJFP6
yCAhvIszfB13BqkGbtSpNhippmtLzE6sU2vhLjfbl0zWzp/XvbnT1Eb9h05d9bET
XXsat5OgXhlkmus3UEZePEFhYs8syvbjbhQpqdzD5mEcHwML/VXBABF91sQv1p7i
M3pTuULrOQNKmrfEJyzL0Hhr0BZCa99sSV1cevbEq5mXjWYZEelRsEUxS2Rhp33Y
p+NDjC1gRVkIa/c1F4ELxOcZlKQitGWV6bd1XOlxfLVc1WJ/0E2kpjMrqrjqlrL9
YNp2C9uHliEXZ+hqZkxzOnl/aGrUHCRNehCNa4lYe0mbsd28EQGAU+cqbP2b7HVK
lO91K6jl44QIfbWhoim5blJO1CjDOxqoRa2FuAVdkyUcvmtxM12DxnelDJzBVTHd
7UEN5c8rFIMRq5J9aq5Xappvh58P9q69QBKESaHQvYFsOJ9XJH9Is35oyWuB5CRf
Vrq/anSdtM5YVRF33CNs1WsnWjIpEVKKvTxU6c5aueB4DjDLI9q+KhQ8yMW5ICbG
wfcKF2qz7aBKu3dllWR5C3Zy7u0Ev00Q5frFt9rJRdwPCtnrbVjT5fMTB8pjriFC
mDHJeRGpxw06grUgS8EWUB33WMMtdjfFbGxITM05RLhWyV3G1O1+GKpBGG/eQm6f
xK342jzNIFooQRtTzZqjFwb4MLDnNbui/Uv50hyUCcyGo14xqVhkHR/93k+xCYTp
D2KAQ2JoK4CjFwffeC1rJ/fgOgOWp7ldky+XKSZ1x8+UXeiA0PPrHQwkEFSkbfXB
ltu/F+64GmJuGYRuLZSWB8JbXw1ah0YLpKwyxcAKSYC5tIjdWK68GVJlGKGwSerk
B6MWY0P1ZppJ6SVtz/nQNosqfRMPN31B8y9ia5Kx01LU5+w3gvRD58ZDlvqvUfcI
USUwa0j/DRV1IypsiC3jD5fwVwdxchrhUaRKFDELxSqKP4H2c3VmkQg0YNZPd4v5
9RAryhkGaFsLUqVO6OSCAozj8E042FBTAmMXljZv/RJWLwpAqEGdaklWLbl4fDCJ
5+wIum9J+lUpI9uUwprFHTtyQVHPSsK1BTdyqjcYE/CxIJ7bjC3UzQaSvlRCVGX+
QeTHcByyy+SYUpxwX0+ACJ+JbQV+gcqGV13+cU3pbnCp3pse67dJNxkQaK+Dzj5F
+leqPWF9TFkyqlfDQJ568RCfJTg/qI3vLb5OUBwnLalRLD5sFrE0zQDn3Zoh46Gy
sSS7ZfK560Ma20/ULY4L4Bo4mRBjrxHVuz8Ob8Y1nYn9OmBaHtjxEvavOTvh5SPe
3twHnUeGjgeao6vSzWesNbBB/7MGR+zqGb0e+oM7lIHbJlNTaTI96/w+m1soN+gY
5jgi+C4VEOZfJhZuLjLqfTKmoJtHntYzhhYji24KZ9y0H1LtXsPkKZ7BS/kOMcVj
+LhufkfftLIJvh0EZaqNZw1Fh1KYy9oZDsYKO0Si7LnGwOwn78upTn29FOPQJ/f1
D5H0MsIxJ7c4P3BWRDjxcWMPvL98yZ0rK7RoVNl1JNvtZcMruT1K5WTAKk2D7ZIu
bSq3SO71piUWll/tRcTodPDiVo4jgzCjMSHeza8xYcsPo65tN246y1eEWduk51R4
UJEsWHTwL5AfQvnneHKceDWnjz/5ACzQ4jPNJTNURDtJtivIWi6pkF+cQGUo1d05
/bO3C8CH86A4jnE/BQLQBfdu+z70Ag4H5MfjvlPr7oD8n+J2CmBZmj7T3m++C6SM
e7j7rGz6NqecfEF210NUVk+J5v5P82tYHg/9NmnjmDxoeekO8je6TPyrT9NRAp/4
aiW1eX1Wl3ZwW+DLsGLoOFVSPTmXvr+T2QWuwyUqbWs9r3MLruAwyWb8dQm1qU58
us3jAUOImT/w7DmaFvKJ0CwagIcqABMsvUxR3PufsQdQPZ4c/d4ttsmAZkRqG3qi
NymnUACD3+bhnuFJoKanUOrBdAtfaG11C8GdWEu5dsl9Wou356p++2QUqbPjkIHY
DZmuy4GDOLP0gt7kYZ5d+6eutQd3/PpfKmTr+INEm6bipDtK8Rw3Ejeg1v4Jruq/
0ipUXyPXRpjZ0p62C/iB4Xn4TPsSv6PwnINdjG+WSCY/JKMqOa2Cl3hhFm/prwNV
kD+UHS4Dt6OBU+DKsAKIc4XC8tfumvKu3Z2I+lqPargJ7cBgy8DQXKhgjlAHRtnE
S2LXf55CZd50XQkTvVGnw2wYOYo2G/+2DQxCyG16t5C3KD8X0hY5ZOV9iPco2dKd
XpyvD3pdPM/RNYkyGA0U6aqAHgrSGvKaZySEbLq904aZ9g2VsNzZGm/unoJcPjjU
9Xf1EC2WIvV9uh3YyYFISAxDnjrBbBHznbjIGPbtDecuHP5hJ7I8zXFwx/2Cnaso
OaJJaWh9s95a7KuDD3KuqRYlqFs3CC567kbZGOjgWMHIXVJCPqbmxHt1S/HBZWpf
i/c9EQ1F4KXoIV2V53cNr7t9mhcBW5T5r6XhZNhC6msL8dbjIZypfSycWQsEnsMw
+zdq26N2TQqIYawv7LmJm0VIf0b17r/TGdi1dIh2ZmvFB8f4JzOh78ikY201hFlb
2Q16YJr/jSbpbjSCiCIuODiIN4t2b0GEIatLasbNsF6nm4Le8fSKU/y0IxwKMoBr
Dv+7TjLr1GZnCmLKyddjqfIS1le6KW/sib67Ds6j6o+A+SWfMHbh63kUjv/9UgbU
0rlWtKi04DNuLA2C1QFnEP/oqXEV6aEGkLChsW/W1SvYJwwwwdbbJflB76NMvB17
+YQ/fhg2H5sBurhtHcn4Fc78VEpPH84gLgLClAtNnvfMiCd6dHtOu6VL1rq8AS7U
2xAs1Zxyk59VM+UEoYyZ96Bd5sdJ7uOh/MzaebppgSbfz/UOcdMPMAAcahqDemGu
p6BAvNs30yaOboaLgaTgj1fYikaPzHDiChvL89TSmCRU/H6ZKBgnPnGHhJ7rqBS/
eyBxOPNY+/Vp6Wx1X6gZcsSlDank90GoyX2G6IWpHWx/tP+A4T5p1s4dxSkyqKWF
ukSL/gZar3Hq0r3dK9KXdCalQGOWx4PQPn2IAQomBLjV/kMq1Kzwf1wn88Jv2IaJ
bxHcUaFTP0oBF7Weonex4+FJiggLMsJULyIPauP+jPf2fyNqNQBn7FRcjQTLZ0Y0
Rt6PCpaTtgQIB++pbvkK7Rz8M1CKVzHTZPKyTWSHaE2IMgHgNvWWm+B8jqfXAkIC
nfDcE/77zW06NWDRGq75vXJU8+UAUYEI4pd0b2xv/USVxENR60MrLLP+pQoWk4g+
FbQE608yRiNlPzdV3T/Lqbj6rQa+Ef50q+SS5Vmz9QhCyicOh9XOEs5oHCklrq+l
tE3o9Z07tlYgnx7nAwPmmzRoiJf8WST9qbKX32ZqNBS/flvpzXfAx7+4jhY8bjMi
Aat0AAbMoU5Du9+jbm3WKsLcxOnxs7UDU8oWya2NtMEd1Q5Udy7kGL7ptOdFO61v
gznfzfORUW7qPeCZAnFLPggGsJTCcTcZYalLVmZnTE+2lCimCXMLsqxw83DSuxtA
8F6wko0im0SxOwZ3ESe8XpA5CoRRq3q3VMRk3isUNouppTs2CvrheXaK+VsN5UNh
1PWr+8LJqo6qGrUZAbVMaTwIcq990JufugZayEPT/ZB89B6KalQ9XWB5sJKp2ZD4
SDDmZ2930lg+WUZJ68J93z1prtGZezGs9zWTLCg1nF02TlBqQXFyz0dIIGG+w6Sp
GGU7Ug13zNqymSXIO7xq+2HeT/NHu4hVcAGT5d2BUkOSSPLkdOpcxyjF/O7kjpYf
dDUdcd92xyXXerGN5nVJAsa5QHE7Yaa0g5hlodOHSVMZH5FvZ6PR6fBabLIEjAuS
ryB+liOwO4HTkorjzz+awM+vzqtuG8LD0BUTqQjpJWT2ZfS86lihFj79apmuuL85
Pwy5lmVnnXzs7aOAsUIzy90+KwMGCpRljkfnMsHYSefTTUaT5YPdvaEgKfJLw+cY
Ssf4v/ygPSvPXnt0BXvRmNkBgNUZXyb/M6JIT0sJmeZcW2AQHgnqd42ziEcx+ikd
j+BbEst/ur7GP9hO/9jsgT2xGRpGV0VAuvie8QKXdOhj+zdtHdn8n9q4P/TX6/Qx
3f0W4hTxgE8JTkoSAT3eRfI90XEQRu50dh5pwpyXnaWUF6x/fAyYKuDTlH7l2its
3leosEEkK7qJ1iCXGuD74SFlc4IbAG3g9mUCFJrVLv7GjGe2c9Qtljw67qVD4Kx4
S20btoZKyMlJVjlAsWZSeRFotH5S3BnPP3e1c+E8pOmlb3/kzp9/DeDPNGLd+EnU
Vndt01XY6VkNkMxb45yX0RcQJZX2iCUv7xF39nRCO7nwEWtt38MBF1iQaZzek4fx
ScRAyksabACnlZmAFzF6i0j5/XB0DcQM00tJOoQrlZ5KlEKkHFCuU7+ZJkAgQnDo
R9peo0VNHfRX0uSykCrVSfSmIHkhea9gVLRurF50zbBatCOp1cvm3SjnBTEWaNBC
l74jloOGR9R9HRT2ibX9O8VspPmQAjT5iFP0n4JPjtHkhxwajK4E/gR/Qbfq5diD
veRMKgYmnYihZwCG8+2UhQtbs3U17JBbmFvHZrxcR23I+qWzZpIkenlLB2jRvtHc
e7wC8cIFfFtPQDBWneTCW6u01p7Y+IhrSceRKZ1Kkg2rcfHK4tIBKynh5XJJfaS3
0rci/og5nqw+l0xm+YoVK5xzI7gao+xL4hcGzAteFG9egC+Yzq0OaxAVtl46jljd
sA3sk6JEwqQFXVkZNwS18wbWg7AEvWim0CAzWBIZ4n5M+hBqIPFCi7l1pSGD/WWH
rRZcthi0TecApor2Twg2yD6YQaU7hZLU8a4yC0DyEEqI2NY7aG6HZuOwyXPPslUJ
DNHzy8/qt2wBQBQpc1A0ie7tdPLla0XS/6UGOi4lm23xtG6m1Ku9FxvICM0hVl9t
E6EN2+VaZQC52lWPQh7JNBWUyl3arcVCvEXwfFJNhLfsb0EXW/TheasEOBJ0/e2c
+Lr245+Jrqbc0QOf8i/tNfhW3ZLawFp3Xybm1tTvKr3V1Xq+Z3HBCesBJ5wb322W
a3WhOrchLB+bB4pVy3nxUf+kIGDSiJmG7AtR7rkb9iAc+O3p2n7PBQTP6WBES/Af
YQG7ZyUGzhRGyEVc0iOJs8W6kMBtq+Zxl7gcx0pxNLxMn1EH/5UlZ4kWn4j80eKC
IZTgBTfa0kowno/wShu7/iOT167PerGpxK+jHDFFZDWcx8IdwcS2sX53TqG6Dpo9
UHBLxhHtQlSaoWLL2VJnC/8L3XsY1U/Y/Pqkwb0Z9y0iwkYf23qK6eV2fwOG72+y
o7REIuXjR21rcSNBQAYgyWU19pCwT2xQL/lqqaCIjvVWcuZ5+SDRnIueYo6bzGkJ
L0cB4dXCSNzET9Pal0Td8nvZ6FAt6fQqTSvbLAZHXU8YWZSpCQH0qRj6SO199dPv
FB6L7l9u3V2d9bhePS+rzXoVj0Pe9L86btIrVfkd0+9r9WkeFUV3NziGgEGPeSaR
HM1TmiUIHF45AaxMwAMhPkwRUtvp69tHdkXhzZty1+C2BE3uhIlbmhXKRYkKN2+n
21i3W3shn9Qlv6bljnigwORx1TmKVkm/ngIEDi9EwWe25CSias1ifoTgaiK51yKg
Q/R68zb+TgU0Fvb3F4F+kzMPP8XrCjfP3ldz4XIOKFQo5sFkK0R0G3vCdfkvmLd/
t3ZrOJnTO/noQ4XyCy2NlZ10Fcpc3tIZJbEfUo5Mvt8+bYWF9jBEyM2Hql0En7/N
1m4z1Rd2sUXVhr08cD345aa+PclZImSXZ2opdJPMQXAx54bS0C4QC/q6gJnweSmJ
kxJOQP3VaAg+NR6daLnFXS/kWez8WIlHfOFz9P8jqsTgvq117B1QzWgeR9Oo7Oom
DUQbZGIMA5zNd2nXLbxm/q5VDP8Uk4v4bMzTYogxcarK9u6uYz3PRapKxrYKO85G
MJrOhH3ND9hF4SmKttK4/0ond96KeLyTJsaG2sQ0/c10xNsdvKHuNSF4tI2xP4Nf
t5+jBWpR9PxQoyykR96mkA6nveVI7fLsavLY4FCyIHciT3weUBRhIlHgeYi6faRw
e+FM9/u34IeC6PcVPsMFlbkx5xT59ZDVWzTlajkhazMiBrImkN6QMw7aSoGyevQf
vT1ZfQ25Vndj0iubnfJRAzTL2+wzHeZrsHHlrlCzUWrfBol6dAb6l3pPmwmakkiz
8VCuKILHhTJajUHk1I8/Ivm0PISmOlrbAbqBUkdw1LJDQJS2ox+wk2VwUesD61Ep
UtoKS0xeOxgWWN4bBIYjAzO6OqfU5mspnpw00BUVVHYZOWKHKuxDQ4+5F8LaG9sT
odg6Wx0HFuPi4fw39kXha+SFdv1ECfQrA671PEpQqkin5AAHHDC6G9WkuLjZZFzZ
oZYaPetKz0HqtB/Y9eu7Y7odQMG8SBf8SP8HkirvC8bVlSNsDMOaLNxBNxgmaCvn
PYuUyA2m6+5l4YR4CClrm1T7KwHbEulet1StQmumDGFne8KQhcLS9SW3imi+SafT
mXHocyvzBb1bcMf2osUtzBJuOk3cLRnlYg1/Fl/SynpYN9FOd9wHW3ECKTniyCnZ
rovdEENaCJU9RSv03fC6XHP5Jep7mIxRKO+0NoOKk1XEx4zHW7Arag7tcaCjO0xm
MxTCmpL6aGoePBQ3e6h66O7EJzjsIGa9glI3Gjjypp58Q39njpuMimx+MW7+uTeo
+TUUW8iCcYqalC1+Oi9gsCsQY3cY9ZdRa0UDEH3lgTuVn8xAJecRgNan7GkSkuxY
C8Dq7A/fOY+USoAjzPCUCckjHHnqIMm50sPjyNFLDivEQKifXJZG85xGPdzfefhL
fE2tvGiWWrIK2mwGCIYYSmupujzOG/3v3OmEcRvN6PZbFp9j9y7Zo6amKRuPIgR2
eLcFr15Gd0JgFX3zeMO+95S10Guldte7FgGlbUpoflahrIaFJ34qWXHHM/K+n/t3
AWhwyTzcKwejPB1D9rg5BuzzWA8ByIeI3piuxEqoTPhudtOHl9yYZ+LoMnK/JuEJ
iZnnnnbZxlA79U3TV+OKCNLF0J5DZoRbdDuVAfrpUgR68V5nhpcEawTsjyV15/Ox
ZTZlspLOGYa9AQZnSAr2ZLyjKjE+yJiNKX1oFTxeMyHsxUqHapAnefv24zSJehtF
rFcDZqDI8I77xRHm/+upvoxlvjg1sUl0QkMnLuPSIZZIGyf+CdhWWFVZa9Wp6VZa
D4jl3r5gVskihs59PLSEiDDoMFXXLtm5r07f/VWMRCeqpt+uego3n9yuoP/YKmhM
mgxnmAdDp4Arx1JW7cDubnUsge4E6bdml5v1o+y5UD6hu+uCcPXgl/+oYVxmOWvw
pZsbMkjqy/t9PI7pLujKitHD7r+6iVA7jIluzsgkWWmzMs9YGYKdoykaEC1m8Fdt
iZCXqcn35KEfMqLuqVRrq4egdk8sT9Qsj4WwQMr8uWCMFMt0vDdm6UJWsN9vzHMg
svpXND/A8/ZSk6ktooLqJBJnJaEFw2Ai96qL+6/kLBMl+8yUDS45G9JBNNwwzBEM
ORZyuK6dMZj4k+T5E+A5ri3N5UFCGmCnhESxAhwUyI1fAYpR4bAFo+9U+rwWDK2f
KwJvSinecrte26Q163OHahLr7H7ZTXSptXHwI2IlSq/wgjIm+OVNZ84/yUw7c2at
bFwTxUFsabjTqZ0RraS8dCdY/s08lw7D2cuIgYbJ4KyF1YnHZD86mL76e+1YVo7u
fNC4wGNAxzGS7OjulbsDiXPwAmELq04EulgH5Oa1MWCFMZZkyFpGyPfnpNZUzrz+
rpmejbm9P/jBVpJ+CKsjBmoh0k7jbSYyIrj5/rmddB24nAmV+G2EAfnXqjifWEFj
Oky46Jm1LmpWhDDjCTj4CvyTAwtN5yujIHl6QWAmbyzONr2XSqGB0o1LWhpZCaRD
Iwxp2Yp2JULM6+9XUKEkFiICn8HoPor2Loxr6YBkymmlLvJg14Ow3/LIiELHqRAC
rjrwqTD3hRSBj3+jRz4AxoDAfR1xNCZ9o1/LG5GWhtWD49EMkDyWhqd/+VrSSMBe
50jPhU6IpvywJqpAyaRWHAmU38a9WsuiBZi8JHpE3DR+qh5p21/VCvqVCQiBm/Aw
bVBKc61pFTJyiZ3KGFfdhWSUT3bER97z7gHpjoLm9X21VGF9PkIf8kdW7gWmL9zr
Ct2CESCl0Cs8ipm86xu7+MvZMkv228i2UiHhqNMUbOVKZHOxUGPLyB5qnIOfq9Vw
o2DAKBfnIwGcgXQX5HNzTw368ZAmbQzCYhOhcb0m8ox/3YK6rkLCqiePZsRlDdWJ
zv5+JKXkA7mB7lAwfGNXVTne3lr9L5j6+Y/6kW53c0U3aQ20ZR3s6Gb8i1qcFZVV
vdEmsDqQindMnzRP6pD1bkxdM04HqJ6W+xBsTNR1gq5T7T9549psQ9FveKeZ4HFX
sNpOfaAhl9EmvtHzbAxSGB34W/B8U5oZXMLrRdVMDkDCXf3kee/77A5TQWgo8e0z
dhPxBpttg6Xfaz1tR4eKZPA0I/Px9GRB9s942kIk5279SUVWp/GOX3Q/T1mIY596
wfuMjnAmZRzAGed0ZiIzwkF8Imm4T/hdH9tAuZbyouPGegPOgzq/7HUVQkyoILIu
P2Dt783JuQAVvNLOVfjJusJO0JeO/TLFEDvSjoyZVmPty/4kank8eK6OV8ONxXhg
pWB8gP0p76FLPXuoMowRfspRaUbuwz1aUBzwb3MsuRaP7ukRFpb1QlfwuE0dMc4V
irdrcIHzagTUzw0gIdyut8nw+jj+twclg2zsWweC/Ap5TaF5y+xd58/TkZlu7y05
qDhXytF2ekgnri8rFKLe+XGaWDIXOITAjUCGUL2otyymTWkqtTJfeYAVeACwlJn8
r18futpyimt/L38qyt7Ml+SaMbapsl6aPWlXZzdtSdL909zGOgGGgKonnqQ4MuVe
9tTuQVTH++kQZg4p7+s8YLtyfbsAEI52DAu7bKMmyykbwzn4GKzLbqy9Ooym+0BC
cDBFtGj8GmAVJk9EZOrrr5/u32X9fVxBhj1Bf8e75ypNhHxQ28MvVrCK2nFu7tEa
dBA5pF4S9wNWNx3i6L5Fd+DPjY9U5hK334ovB0im6EuU6hyp7hwl8T6i933fp9J/
RT2Zmgya5spsmRRu1PZdSsSvzmLMxoDn6L627zRYHW23m1OUClf10b4qgQkN5rer
l4szGvA1P2yyju7pCcye6D6tZJZmobDJXyj4ax8p1CRE7xjki1Mi/K/6J1rJx1un
TXqK3eyz4DTBiFoM86VPSZv+XosF6uC6VzFO6LZ/ojjtWpO32x7D026nWJmp6DWh
pqxq/c32qFjcAKAaACsJ67IZsH5LT844SGpBzBYbufbDQ1/vCAzoI1p/l+aK20qC
FZLcZv2yJ7w4hO7DZunaWNwtV8dLMIqAbejsk3fw0On8DnT47sc/Legv6t6dUipL
oRmI1bOJYASMRXjVYjiEAqxBNWIqknaH2arVtCi59JaFNR53a8IqoyTFCOVbboVd
+tpzAcgZ5UN2KURC4QXrSXad5fXVEqUkFqgAazq8w/QilYr8JxTLj807WIko4HUi
iGuJwF5Djn0p+jIJuqK3yvj+7tn72+NKb5p1cr81tCNXyjpH1gHgp5NmYXqCjgbE
nYLBRrSnQSvUwLK8iRMnOSLstSKksbai4uWRebyt78AGoELW32QMQYMBdhVfz4EM
9q9nyjts1KtjOzexFXBbUS8uap5Ys8zt45Ic4CjFBtgA9eVjGXCC1IpW/Mq2e8hy
oY8SBLCDiinS5zb9j3gKMKDRuGh9iD+IlNmaWqcsEBpEy9q4DiNaSTO7H3/473pg
+JSISkidt5Q+dnLKU4n/EDEytphb13zPTFjP374f5D9iTvU/IvQn2sAwVEIG+ZA6
b/LW90C4GAe7924hQPcmcuP5lFQbXUEYGwh9nbD31uaCX2gZ+imUVoLYwkrFvvO/
rbDvhI6hvym7jiYnH3EFJaD2Q40Nwryepni30/UhONYz0VhQfDN/N1HLNEFWv4Vq
Rwca58hLxfygqb1BXz1BFko72lLZaJOD/HB4Jd52xr6jT+XQb4zltbDtgBxdBVpB
+kIBfWdGtFIx10hXe6Y5MyYyuSbuDWvCZGioIEOiCkjGb/hkN/C6v5757sNIMuCU
7oGBTLIXINksRaRdGpZ+IxXcS+kgYTNtBmGoqepDgfhm98lrfy5gwEsK2yfuaL9L
ioPWWG94KyrMk6diY0jn80M2hE9IQsdLyj+zNbnqecAZ491rndYEftccwZIv6n18
HGej4wp+JrL9hI6+iQJBs41zNUwu94j3pSH2zroGjDg3XTdobaEsr2ZrAnyErmCe
XA3oMYDPaoEQHPmQjvYj9p85lOHAdnsSlIRMTqhy3gZ8zIDZG6dSyNcTXm5kgtZL
fNpRpaSEoaL1MPk3QlZ6MSVwaHcj/O69FEp16fo/Bsu3xcci1hauHJh+rgL3NbTg
8rFyATmqpxp5J3f2fO7X1OYt+p0ghDrzqgnmfaT83AjT/+izwzZWlNevFQuiSXxT
rUJlUCfHQSIDGooMRiXIIzmFHLSFrj19UrlhaTWpoX6mL/Mw5T/dUV+udtp7S/RP
rGtMMiC5mmWFkTYqkiGJfo6/zrQG94GrEKzDT3vUxAiUNuDWmY2LPjmCp0XEtS7/
8S+ViqCJRMCJWaTXyuoZP+pvo3EP1xKMGxdbJqSFWaN22Q7Sa1kCeto4WDLb5OnD
AC5BG7TtVZnHdHnHyarNW8I/5i97KaStg/jKWp2NEkTfA/NNnkZUh4ywtNCbqDbt
O8Dty10oNlEuwN9qf7wVUecfuVGAL0RqBmPM2KG3qlVhm5PPtrpw0ZaJlBadsavN
TdubhHWxqPXT4F8Vd7dspx42805k3Yb87DgyY3lWvgr+s0GcQ8fKn8aE1Q3XmlqG
YA0wDo/wcm4XZs2cxs0Lrz4fn8cKq1IUxNFrM57PfJA2gAT5AHfR968XZ060ZP7y
B8R+krZ1h9eyMYzzWzWYb1PIXcVxmJNtKaJmJd5uo9EN+KcAXZALYizi7mPrmreH
V9Q75QMxsCb+8HW6auY/xZ/rTt/gifrRN608PKXfP8dRD8OPMAfoXRR1SQyJvSKM
zsxSsb7Se+EBUum73zwfj8DZn8kp9ra3pfhGMnk3fvxG32McYfcdJD3hSE5e+BLo
GeYQ0o9Fj13vXoNV6yLNtlNF7r7TkumAA2W3+ARsO/0Zt2GwGVf+DwxQjVtyeHmq
naox0A7anocQeZYKiifX305QwWxWnR/FKxdZzJR3I7WovNz/FTxiguRDROTRNJXv
BJnWx4EeCC+8jZFX+6k1uv3UJvaaTSXS/SgVHOWYMkJ/QYBkHR7/3PMp9q/dtzT8
yDEyQewdogHHsrxLsv/1EeertJnDV83XyQj0ZAYghwy300UPQ8CVP42CsF/059Mf
cu4WoUvy9sY2t8nVrcsVm5SvvCRHm11twRQnOCHv8VLcitfHSqsXUHnqs9bxDDIH
7J5ufuYd4ZzyJqxcID/wPHaMd1sNITtIjf6m7oDmIExzxh1zTp5X8xozpEE9sy11
tdLfL9yafA/UvWBrtrmQ0SzXkwCJ5rtguvhd3A14fb27N6za07dyb8cOYU6JqJpA
QLg2CDlvkJsX5HLeiYvgHfXuWdNScRbawJTpLx1Fl5gS9xb7TZZLqqPdcTiNufAN
XWT/FvozJ1YZ5+F+I7koqllLjP7UgjaA8Xb99RpQNzn90twfa63uf2OhnkDfv8xh
cJppIhXntAg6GyfrGB0hwEPWUi8VRPDvenGd78a4h8mz3fIj3jzrn0oP1IUtYdTB
/aFAJTAseIrS0sbHMb1QOUBrpcnwXn09NxyE5x2hLy7ue22Q2KzNkYULUWGr60wI
fB8hKuftfvimVsiLEkF9DA9znavumYCELARO1Zqu44J3uq25b2n4nEuFuTW58IOw
vURoqjEyhN/HyAv5Yg9HFBrL9jBaGI4WepHsvaJzB4aRcWzlcpeZ1fE7Z61H6FH8
jQpEq0BvA1sXkAvlmG9rj5q5sTAOg47lP8PeL+XAuDNCaOmW3UJpUPpEB94d87Bi
QfTsKKgo2DWdDuy3HIAWYvXpLfobGKUoUUWxghBKSVHZRJX1ISiLFxd5ccyJQetj
iQQJl7jnw7TZxIF8vkNMMW4VJ6nAuEHphgTAi/eiSMHYs3dOksNd4EpZtmgD5Wv5
IrDexSTsS/XAcOUBifjfgmAfrVqFaFnwjwZWoNI6kRkelWHQ0Ll0N7GULqXVNL5g
t6S/zVbK8pp6U0ffqQ4mKqpOXn22uIQNUZGUPaEodZ5JclLjECq4krT8n4OBz7kJ
/78JUrEcKBNZDD/HYwsxaEHxM1qYTR9mjYWw1gpCzlhYUXZK3l/oVTVC8meC0Tr5
X+pT8vNqRzreYQisSh2cQDrdGw6LxWukDByrGsIv/VOxrSeVS1telFLVUaLg/9ny
Qr/e3JnsJ+5F7afQ5My3BXzR02MesTBm0+tFv3NTdurezcfW5gzgagHVE7jKI09e
/fdcEJqJRFxUltuwPem+I/hg9eQPMZdPaLCdNxQUeB1OdaMhBXcJMM8X1uljruz1
HhCeh9ywP7bnCHrDbCDedViJPnAqVayVQuU0aZ+9itOTmFrX8yuon/IkBQpyCf77
92V1i3kxT/XMrCl9gM9pOV72d9rr26re9TueRjxoYvM19CNk24G0QOSKJYvIFTNa
kI6FdCQO5fjtxxxaEF3O1iZ/GRmqruwKtpI16CXHMGwY0dYMq1V+dSsGV/V6IO8Y
kz9gbeaGiuAGCkmxQj4Q170qEOJP5AN9tKu3CjG/UEAe63wi0CZjurdvug3+Lk+d
5HZpyJpIM9xpUcij7IszFu8jb4rvPE6e1ApHZWr4Oz0fTUM1Hom9ZAgf95znS3Ew
aRhjfLSY5N/95jITsPBmegAdZDtm41KQ94PddJ4NdP1mlsMOy0GyHwDs8hKE5FTl
sXjzhCs1L278+ySykvv5DyEvP5X06QVW2RtpmjU2hs0+Ex+iyy8swrqXTT/x14ts
HWBCrO1OYfnULS2rwrZSNHzsFECfHavpq18v9vOXbA4RioL511JkUzH7CSmSMbtX
ZZ5pQ5hAiS3+/wxcnHUNCwuLwnor4pZf1oMtAAKWBfb9XQ14hNm2YUjD4VWqU7nn
5YemR0Bir8at0cGq8gTwgo6xvPKzGsq8M7Us2gtC5Zy6ftvvyGab4kDXAEyGMB9P
vSsVFcSYcy7dsvYEyFZmTappvXlEMjxT5KbW0A7sO3Xij4rIHE/W+Nv1extd9i5+
A69KAmmeUO4GmoBsJ492CP/oCWYPQyoP+xWJ2wWR1sxKmhd8X7MOevOHuIpLkGka
dwNeXJ682Xh4+TeSVVx8wV0HtpyHy30vWu+2sb1qVjgyJFZbZatiSOmtmtK+XE0x
L4Czh4u3S63RL2cztlG4fRKm/s6/hIsTGsPtmFS0OYTdI6etcDKVNG+pFSzrjLn1
p+E0tSYmSw7ARZ/JD3ZxBzeYfoAiTT6/0Lpl7HrdrIy8kQCV5RQDMhNkMlZ2EBip
NxRLAV1Jml93hF6Upvwnc5bxRFv83gLpuKcEyG+jWT8A2/SfQDn25898iDshr6J5
MCMUtH2tCjbGlWgBmhegHX5QereqcnsixP+x/dkC22aSfWFKYVN8JZioLcJ1c0xI
VGDI0Nw5h+jqdGTVq8+X6tVYu7Qv5HaXtzkp+XLCU+bF9u3boImWpLnY6TK1Cfa3
mupbyyDQoGzP6nSxVKmtdRokP1g2phbBiycz31gZGmIM3IQuo/BjIq4mCW3qU/hb
JExRqij8RSVRfxdN6bxb82rdYbFtIj72/mo+YVXOWn/MdsF5/6ZOAAJyjQR6Kvew
7ilO99pnvrN3fKN3gb0mpS/5tjF7TzDI2lH9rKvB3/lgi1wmZ5HXGwn+qwErhOrh
6cpLxVsQs0SPi0Sa96h7yCIC+C5qN6mdecVptsfC7Gp5NkozggoSO6ztgATFWvZx
ZFYz7dr9DSeCzkDORYQVbG0I42AAYd6SGWjEBFdoIJSdRriCU09kKO1gQnkx3Xxm
DRLAjBApRqgktF6NnzxmUOSTLDROk1le/38oxr+879RP++lUUUJ//HY3XnVagrEi
T3L4+lbviagpC5kShZfJT4pHWeu5sfpSXWpB5w2WggxeIdoFDpZbcCJtxWP9fW/g
OjoG/UGmVTxQaiGF2tpgpiPv0OVwHgNzTKAKVEYVSDVe29JDf3OIWHglWNOOV/kz
aVkQ6SGYEuy1ftoUGcK1hoqcuHAKsvpMRhuVlrDRXVfK6CtTnanqt5LlZrN8MqzM
n98BdIZF9C2ieX4Ruxb4pnxVfwFw2/EF1YPeeR0Zx42DMZ6a7I4ZKCebM0u0U8zZ
r82VgLn5bE2k65VWsOI8g0BGWimb3n7cfpslzOcEuoGoDyCX+UUuzy/xttsN4SP/
3bafC3AGf7jPY1ibDFtaxfj4n6fy0IzNI2GuA2+cvIkQqCz3P3yyhzefB61szlJO
gyen/9jAmQ9nr+gvV9tESXYMjbCkjzyqdthRr05CDmX2e2jNUVHjxkqNlaueD+xT
6ji0LRJFb9qEljGYnSReBl+ehx+ovp5d7K6fQ+zoyFAT/DQLVK1ZqLf/ui0GeB1n
Cit0p1pTjy2BtAIfRcaEgz/LXTwtFjv1Rb9t5oULhVmZvscVqRaeGDBwkgp7j5tw
zXW2hjtUEMRNaK38bg1GEXQd2FSgJn1KCydAyjpAG7Y+7fEze1k2hdkUqWGTGmiy
mDQtDym9L8EWnT2KGlMU7d05l4V59veWEwpg0dTI5VWjZcfnELxr1s1zYc/+J/1w
Uzo3MzGBMABWFc+UTRtxWkrMFuqDNXB5Z/OCEKPWJEOnNlX4inBxcEZfhwLPydw0
V80UZ+N3Q/PpHGUBrwfrj7WLPaNu3HKfLRCdy50o7jm8fCn3M2gYVtbL28TnXdFg
A7pr3Ma0U/nkNePP6y4/B//qLgHRfygCUPUC/XCe7Sz5Wl5RU3HA25I5Sdhtt0bJ
CtjxUztI69nAjD9HxpqxuiHnI2/rcsT67Lra63BVN0ZqGCH/uJpXkrgzRBBptts8
WBJOd+h3gTP7nEalHmaITXats6Xs7Ife/nfVIuvfaJQBsDsvErbDM6XCtG8XGAqY
BS6Wy9yhZPTSAfL23n1nQbNWQZxtx8M727SVc+KJKdSdcfH4RNtnBoREu3WkzyZ3
rPbnbzAQEZJt+3QfpgVaJvEZF0Kn/zpkMh4hiqzQoQKv5aLE5Uw0yz6tLB6n1mqw
AQrwCrr3/ehQY+tRfu6lIBZZw633Dz9gJtgxE8Qu8H70g1QczDJ3mpPtWjWnS+J/
z8tgR/2GqtrhMR+LQl350GWTl65jOObvBusO/rxkQaBgMfbnaWsc016wvyHqvjYf
Ww3xWFeMzHkoB5z1LK+/fWXTV30Rrz64vVj7d12pwp6mQAOBS2UCqMs5oyymb56M
p09zGglUqZ4NmlsPlLt9diJSjknYjpdT6ETNT7AwQrjaQYuGIAjLOSGSuSv7WgYT
DFLy4sTFgEuTwjkgS+TAK5RERypFXW/ApIqwn9z80TRzddPRZLJy/+NjE9RtmUHc
B3NqV1S6S9iJ3c8NwkZOULg4BtXrTo+rFbLfIi9XxTP1eJ9ZJYElr+U9pWug6gm9
vyVmF3BI3Ori0CxpTFk4O5yVELrtSI/owgF+E5/EKanwkeZPtH6Xz3qRNM0JFFeM
v51wgL9RNVNqOZEBS75MWFJci4mO5pyt1KY7F86caSHvsf7A/SxyE0qL0JZl6D6i
3xANzx27xZ/VeKlt0QvEp9T8ADaDYvg2nYHbR5gGD5jI94HsTFTWUaN1HofCZzow
y/GDayg6tOI8ZJnTaZr1/tMH+LvfFvX8qoO8E/Qm+BBwcnZ9hLioBDRQn2ZXT+QR
2+dvQnfVuKEhPyUnq0Ifvqv8UdKdKSwZd1ZzwmBivN1BnoA8lnmMf0wXN50xAA4E
2sBTaBtuI1jLbpZHmQMO2zURnXTU5VJqG4jwMA/dkMsAFI+aHPwgl+4by6AVEwUR
bILw1anLUu/LbhSfAjKW4C+uF9aYHFuZ7Pyc+RkPqM/DMMcTQFxkwNcoWDDiQwRk
0H1e8tWrJhGcRUqtnjI4BxiPSv5EKS7YajHxGLHVd/PojlXecFWgT0JDK+uSGiFX
kGi0OvcJl4M4nvjIzN1DXzBrJ5SeUwIPmRDY46pWMGvndHyJBeCVBm94WS+FxRXW
wr/KwL1vF/3iknIXUVhEl+0POiOf8TjAN2wlKDpBE56ZydwIQbKwY4lS0P7TCcGk
fN+aaxDKjCoRyz8JP5fSQ1A6lv1JfonfOAvuoNdg4K02z1LOl+glapdK5uV7qlYm
XEv6aZq3GujPlxqe9b35CW1FWofCCGNbiECTmwwjl9ZhbOM/i/6KeMgmj7OK0EKn
qPmX7cF78mPwesez0eo6v572CehX6U4YPF231BIqIntAKSXrmvYJBLJ6ovJu+gQt
/oiEkEACcfGFOMOU1fzjW6de9H71z9Y0ZoHWhoUvAjE1EiuyvWEOO7xapP5HFbv1
ngHzYnUdnA4clW54HQ2uhmYDLvTzJLUvJtcRj0ZYP+ENTv+EtA7dSs6MgVG1bfHL
YBcOJ+ypRUZh+2V3/9aapWuB8OdnDhYlzxEGWO/yTXujNAMBQ+ytEgpuI/HKvQkP
6VrE3B6l/zfnn4uGeHfVDl5OQ9WWl4gxBTV+syw0n+KPg5VYt228+2+Weo4uRerI
VMkONLgSLKz/SM9Tvv1oqP9becA+nU7D8nRXCfI5nCvdy8pqr+fpbIe8F5I5ZMbS
Rstk/zC51RopEE1BYbU5HiLgCtucgf68b/pBalckk25HRYPjnF053SxTovVAGreC
9IzROTNDwtMaMt1U+knBrzf+I6UzWcFVu6HjEHTJmz21k+YU/S58JOkkAeYF+Y7b
WksiftN6u1EPgKWweSp5udfuStmCJIGx3txkas5R4RAIa0XMSy3SDnQ9ctgiFvvQ
o08wQdPptfe8A+3bCGOb7jqvPlz8P5YLiBGs1aswaz7n2WtC08JTKDsJRxvCMuoK
p9SG/BXMdUZO11Vr7c/uJAIGUFfmsbkFjuqQKD7bJhmjJoAl8utydp/uxkTeqY0S
fv3wEdnqVY6pFlHtiuByq5AAt5jfz6kfImNBhotSh8e2auhqRBQFP4wlUYrN6AQH
v2fBzlSzynLHlOCn4W2PRIKLtB19VOtRSrU8qrHDJS8/AVakNJqHZBq8GjlagTUa
q9JBEP7+FghS3vSO+rwiOojisBGYvUkAM+Dx5H+kONjD0R7IL9AFtw4tziOTEQ/c
Jz1F3DfxsqQcgwJRBC2S20ziqGeOP9mwdL7peus2NzhvMDQah+NB8jYjbLXP93OQ
p9mgthyIK6O51tSwtdXkEZwUMKPsU3uh2dolBKkScZGyqlS8MH/cNciibcK3lUxo
bLE2wOiYKe4cDsSbcUWVXCsJww08ALeQmr5sJ1CrmpZJNDmVPT1ry/ahXgwS0ka2
ldaobS7diAEfHeQLP9A6RxuMGNRVE7ZR3Lyi0sKERBIt9GKG+af/cixB5O7nF6Nw
eBOBNZAYkkASBHYBnj/0ZhVl8gBrtC3SJ3Rk7VjWaN3qHPjPaSvO0kFIfCF9lZG8
VXDECjJS4KCXrdeHIzJf6y0MlHYkhV5mrSV5UOXmZW7eA6Q66TEOFbJMBMCLHJzk
M9rzSE2e/hKXIH7SJUdMD7mCi8lqA2iAx4ZMsI4ai3r9F07seWO/+ehpE6I0iFcz
Z0Lkbe/pknZZJ+rBU/npx+468g94PVugBj8vxr0tlS8ptvgRfVOWOcKjzaalq69b
Nvhss4+CfJHNAmFg4cy93iLGZHYts+FVbxDaB1MN9LUO5JJ2LgAldaHvP/QJfGuu
sm4eCM9bk3wL11T6GE1pGCO90t+aZJLlsDZBm2Nmxq1X24RldvuPf/aqj8WfzoJk
YMYk7kWoSNtiQFg3dGfrOv3+KF2PXd65GIyWuGv93ZfGJJNFIJIz+vx+1Y+227Fu
z5JH1iaosGpDiiw+mxACzqC36uNfUr8uyNsTe09PLgp8mImCzXU7RsDLyAfh8bYW
+5hwNWY0i/vfW81dvb0zsyH0ykLhkHirhKINzL6sFOq4UiXeA4cB1hZBUNWtsJV5
WF9r3Zfa1bH2FZkarMp+5G+bZzq93buJVyGySiQpUWz0X9xwOjcSAogHE4hKIsaZ
AaWaKcEh8W1QVK0NpXtpYZaWojeFSIEEwChna46F0aNdH9ad2xS3NQEGneeWq5a/
jns+H5vMlzrUbljSprJGZn06Ux7pJXDL9mZkDpxRMshO3DzH3AeV5c9P1QKOGOhh
DXzpbXw651ngzGdr/r6fLxKx6tDPDwKtL0Ow1EEpiMT6E4qw9udt1xGkyPm7J0ds
Gpeyqwh8NjXWeFsIKvPvDVOIOCvjNFGqQ+YBSNbrcGlsXtmxDNS+y5czap/UMQfV
X+C7fZ2Pwv5nvN/PgZTf+6Zqb7xtVBYBZKaRRzec4hCC5ROeRBe4Ncnia6GMdufC
0MZzbatzCK3gPgBRYT1XWhN8Ek1QbmtTRsNclvkSToksjfu4k6Hf0fAIy3JvWIRj
L6JeEns6/rBw80qL8X7/NYqsjJaD0jJRHbdq5l11ZvyckyukjO3Y6skMp8B11+zc
FqsG8+Z065lUkp4pJyeWb+2zRrg8336UcTvNaOy86NZX4yI4TqAiW0ijOcs3BnIW
ExwP+W+dnn6atWsLHe3hiIDLJ3xDMSfSDwkqEA+0F1RqfT1SIFi0zjZRxVkr1xsp
UwmZTY/r123JfaqvJPTe037XeQW3obzk2OEQ+A9Z6/qtrUTtd9dUCw/ma4D4U7ti
u8hPASplpC3aCOh+qKUoyFsRznps1l+xuAWX9ZEGnxZwcyQf5+sGMHKjnLYpMXeL
PRoJbgPWLkpAAh31BYd5J97J7vbCgnIqFvJL8muMA4QKBtyGsTS3BxjIk3PhU9cg
wyFxeXkhU81d1dn6r6K22oCm207TS7pFe5KgE6xWY7jicDVY4rMQItVvSHGTiZqV
E6crRrxHHgCiwVl06+6YUdQZqrYj/uhv2CpLNGn1Byc5SsPqLI1jIkCazhnWPcXv
ok22c0vv/hP5kY8hTGgrNLRp/Bk76es9BlBgQ228ZI5ZlUpDzs3xQQDufXaamAwH
UpbF2OywO7ZWVyj8iRMF+sVWxSCyciuiABIuWr8oKQHk+0/Lr54Tcv9LkDiXJBy9
n90iD8xmanqf7R7a68Ect5NDCuiVEJu2629Aw6REU/hpEJH/3H+lA5s5/Xf0n/Mk
OJvNJ1qdT/uCLVk6Q0ZQ/EbhQnYaGx2rUv6Dji6TIAKIdoLY2Uns9xhVFtucUkU9
ss1ToiYFB8t36hShyi32dVu3Jy1QeG259BzKlCiNwjkOuJo75trUPAQFPqtM2pCK
sVwMz3qXJXFLAjRJxmh8qa4FA6XoW3WlB9NB97GTyIS2HMM/frI0KekGAhq9CjLj
KncZkE4ySNVk79K3wohAbRAljE/fr6+cJp55n3yjZXXf0W1cje5/u3uUWAvWhurK
Pz4VEWkx4wPYViOFdUbuO3xBadoY4ivFKm+xAZ5warcGhQNHFTgCW/K5UelORKLY
dq/Dp5Je8AOT05RiHyFd3zCOoUTVQ8L+tmxAAAsIUHXITxklvvE1mIFHO2mBhDdG
yNHjOxYXYKOwVC2bd2q/dha6HjSffLNpAKe+Xpqx+FHYjbXRNW6lJuB/23v6Zc1S
tQBYwSSTdRx2/BDchQHp8AUBuFgaR7+pQlUuefjA/7v9KElijoReRhfQb15Q3taL
QiVZtucEFfw7Yi3FKK4faPxqv2pwl/b7Rqqq/hEvFpC16A36XTlyUghTdXGNThHE
AG9WaZtxZS5RNq0eIeIiKmho2+UtZtZvXR30873BFXyhlr+NQce0+kO2iGtKvt1u
sb7hpe7HJHlS9AMpckNkGvFQVPNR8dBUg8v3e13hP8EokhG583Mowc8IH2Wa+srd
JOJ6rkbvgjLy2obpkWyZenlPG2kuXRFSoa4FGMdrO88IhyQRlHEGVY0/Gd7Xhh3R
0LZSxPb8ZdctjECm0UDg0SY/yURpWdYFgCxrS5V5tfHIvWWEO+8IVKysBA4bscN9
GkZxZQkALgc1IGybzNrnvmumaGQ+8GpJLWxcaDmoJHP3kFo5uSWD7LJHpFuPYCUD
+AN/Q/G/ssKjZUWxgfQpNl9IebYIsJWEnlGTOYqY0JlkPJhDnHdRBdNIMyqMHBH7
Xy9nsZI6/pL627eOJDpIHfg/JeKngsVUGRXEoH/AAJDhAwJt0bQ4A0T4EQsRtRXB
Z5cFCKJU7MQeDy5xnVPFzWjmk5+C0eIdkUq2X9IdsHZheAubmawenDV/8l+u7vog
hQxXY8ztINTVzq61Wd3RDSqL9xP891nE7+Pees7IfsK89q3agrtU/WRm9w1+wv8E
vv7n4DfqniaaiRahlRQXjIX5Fs2OCLRbDv27AJGQSoWe3gD6tZwr0KIud5RkrZsM
RvOblqN3BCYKru4mPA2FwJXPGKbJbUGCOU0qevEfoKXPcfbngHnM1r/rdSUCPhFg
EG+bNFmxtJH0w1bKA5TBvKKoQBEwImkvqxB9Po9H7tQ50AIevd4/eevOLg37oLE6
9fcW74yrV2P4ZKYBHv2ZivHx+cunycCbjVfO8dkjzQ36Qj9YYd/3cOZARjZszsRc
tKA5GzTFBYiCnNOtUApDyjfh/Kr5vUiPG3JI6dG+Y2wM4Vg5/jXMMKh5/Cmuuu+N
qFlak8GLIRYrDdNWWjS6GrP17thNmmxAdnS6Bjrb1jw0lo9wa601jQq3tS+SVY1R
Z5y7JNkqlk7Cl9Zemfcp6BgWmgAn26FpcGH0zbr2HERPWvXManJqEfBdcAwACfTj
DbslhHAQQMcFpzfJDlmKRZSn3zyUY8nUGkIHsHD1fGV6Y2VSwlBCPazMZMC4CYAi
lMXqxTeqnYvH9O3T7VY3rZd7qrLQxtf09wynXqFXL189g/Yyi6BtfK98wf2L+z8H
/mrhbmm2vzB/hjQM/mQZfbbEsivRBpw8hygepJzyt8vmaYmcF1raIOKC2XEtyCOn
5SE9BLZSKVDB6wKVfq338m3opyUnyRA1QTZolPmoxrB5/IpJSLdTtwveGz+bLd8X
jcHuKfLRqi5DmWphR8pvzWqRf/cg4jF0FTTnpo25+KpluRoRjI4E+gE7aT2AiWCz
/9woeuQmEcnS7xxEJMg0zWsIWNdtFiV1meOD548zJViu8BhbxLQUT+AmyAQhjPKH
ZBPCdPbOGXBB/GUUmQe5Pt9EZ+z1ThRhMo/JJPZZZ9pQO/lc4esJG8nY0d2la2wq
T4ph6NDAY+nCyrDcdrURMjwnnsqLF9o7yuV2sj0t96j3QbzkmAV055FFfRiz7a8V
mUsznjxM35r0JrqVfH/0u72hb/JRDdHtPDS3kefb3WUrQfaakBJJt3qfPARU/msc
DuzrOIqtU3V8RAzXjdx7yrFoU3EGhwg9tnny+FqIXwFlz0hnW6Txh2mviuEOs6wd
YC2AvyQTmPi/ehrLqxXB8f8KomBqDwvPz4MeB9oy2e7BDlufmP1H4Ytz1WuGT4hO
V68h1k936dysS3ANr290uK/de2+h132i/3jdUkSJyXBFhVag8hiQQ06lEF02vBO5
LrvVXukI7h51EHB+FyuvkqFWuVCcJvf3SQ2vbgsOqBbVxUtBgk0ulhay2GJEVPFj
RK8n9uUJTXKGd6VO4zW83v/6fHk2Qyo1ggHqSgyNSMDQTQVqOGRyhsiiRmcYtHyy
gobrq5tzT/zjDUs9pSHl1x56VaQoyygo5h9ZhxVvTJPpf12d8QxQzOK+4p2OsyNn
17M7p0tnttW/4FTQggxooXvvaYWAhdkvMAXg8GLWvV/3l5jZ2k3sRE2skJDV81eJ
seeNP8FVxSUIltqXqkP9CH+VVg/GSTTz8XvUSlmJvm6Zp5OCrGg31RdddRMHiZtO
k+CuyheC2twH290z5iRhQiGbCDR6+K5KUdwQSnWzEuM09W6j6AOlkuzeyeREPmcw
7qZaVmMmiRZagUc14jhcd1J16LlzKLqpwrHCQBhhp/loQawzlAIRwDd31KXcTv+g
Zq9se2uwGF5jaHl3QULCxnFdLt+9LV5QEigRCup1CXZuuk8r7KbMOg7gLpV6FEcS
HmmWB4ldLDEwKpp2Q027hMepnOsTNHJDVCykEcyjjJw9VF7puGdK/MJSxORWMPEJ
zEcu8SYQ+X8zOlpTNYMOq9ESFo7zUQBiCIq9NwGZO8fJugjPeY9ZAhpst+zUhe+I
XAh52jWZwR02knODioRY89IoimZzuazb+BBUP6yt38yQLEfHlWL7SEMgtm2hg/ED
Xf8mpSB1CHlTUV6HZFZbDiA9TYxH8n6jkEMiXubTPsUgESHLT10ChODya9wbQYNr
GbLSxF7G5DJ34WoDkh2cvLdl7Q4vHEsCdJVcPgmaRj+BYomXOzSB/ROC7vsNj/5D
zOK/jDXgM0iIiOfiFLsN5+YJzDGJuV2t0SwkJDOVRIJ+8XVWWeLSeboIQPiilyjk
6OGv6aDK0SldNvbPsSBqSkuFXeWk+qJ+yvKD8QGvecbHIvchxHI82OWIgr1LznM1
+jTseCJwwGk7PcDXxjGVQrLMgsjihzK73F4Rgjv7eneqAzgIwziVZ79cnzaYlSCH
8V8dwGF8QJXAcwBP0dvXogzuN5qu4vnqgMxoh97EVanjGZL2+7S/GqlA/AKj7jnU
lVWrVnAfnO9LbNazpQiBOww1foq09LAFnpv7lqomd0D5PybzakfjPlHcAnZYFOmR
jpOO7H/J0fWAXV387rxPFok0CWwfiMvqNEYDilgYqZkiZfC1J9gcBjeNoGWS2yXj
149o7ie/JSOBj/ukiLBOzpttGlQ9qLqRgi7d1XaNMe+dD9vGu61ZXeAcsRgxp6j6
hMjNv1oW4JFe+bU5IG5yyLjjwz+rgRQg/+cfTu4KUVkEKGX8/wzgHT+klAnVo9Mg
s0/Gi2bJK2FHDZy5HQOZEWwFe+ZU2NK+fGLD5oweQ5+GDPGLBmoLr6txbNhsWuw1
b7tN0WYQN2/VmbUWV8nhbHItqTSYeWVjXAPPics1LGAkEc2vSmWNt7dzBAbKlhLt
qkGK/EkSaPQsLtVghEWUzCWvK3JiJew81QFS2v/xRQ8cN5TYUkhgJ8xdxQI/8a7Z
QJ8gPctSQ7+JjBScIe9gQmiOXW4TER7ZxDaXKxyxnh1RZq0iv2CrrRttECwuYpTm
GrCPkW925eJLr9Md8TZprkSt5Y8EIRERUeM4nQVyJJolr5llKqobX4t2HrNtujgr
C5mu38rJ/zN0zLzFMZjFdsbcoiV0nXz9NESb50J6TUKxv8xT21Ck9S/bw2/8PzET
v3YRDlkqo84evnywQXbmpAjtzM+RRQHEkgrA6wQ7Z2svS1HnZAnbJhMSPVGAtrp8
mOAwR+2WpVyvIUItU/9iom3NfSHaK3gQsZPVeyvL6Ux2bMdD/2Wnmv3suZyBlL63
OZAiufYmUlEn03uVtEkxrawLLvh9KdI6SCSoa4iSZZnGQlbjCbhPvkUFa03YFXRG
m3IWyy0P2Gr8Bp0O0QO+PS442zrWeQww+77mv7sl1O3AyynkMh+ELGNCYIuIcpB1
fVndZ38gkqSkBvEu3xom+OvY5iRAsj6uqvKlX9uL2sj+bx7M8pibsusfCWnyWNN/
dkzV2umyOPWkWCbUFDKHX8xg2+SCSDEFrQBraR5uYnRFdezMCm45qGKRxteqp8LZ
jiDYkEiIQE3QKUC9VQSIae49iX9D/HDQArvjk7x1DBNplzrSdUtX0cNZmIzlVBX/
sqg79mHIasf8pugbufLMic6VPb02jdPsozEkqB1P4/zZWzUH+Txc4tuZDC2jLrGE
pmgf4dOSqichfooNNFd3avHnOS66gCMO7Y2dCmGVqTel/JKPTzGhkjK5Q9pKivke
iLZ5KQ2O6XH+vOJJ2Ubb8L/tQXIenNwFEXO+cO4U6fevkHXbiBociCcYbO5L0bQu
E5kP+8VgyLmJ4kY8f7uCsqYeg4zsw9GHl5hPCrPUyNhPcgrgLUv72ESgn3Y+UEdh
ombbxqvbQjbIzqjmXdr/VxsdRz2JE2gYR9B+M3aoFffpYJ8Xk6AcsofU4agsl3rB
D+tkQi3PoskbgkP6/H+BYrKfKsdweJl5Y0bj/MX5r0bHXVx9ifr41COL+jP2xGD6
/ei+/KLUS5J3XusE6N/7a6m6HDa1JabLLk6bpvLCoDRKZeMBpDDcf+1OdEcbouMx
t10yNyKt9AYjinWWjH1fZZotfKrGjTPfMp9e/9XR7PX2eBqMCdIqS5KOrp+tPDHk
K6SQd/0B76u/E3NzGvpX6OuYB9A6MxukSELcODBs1oTgSf5D+tIGm5u78RayT7Ej
yiPZpb6ZDE2XWVhYDCBLVrm66kXGWk714iFfGMUoHr1JMd7nG1Myp7TwyzEKbGyi
giYFuX0dpkVXKZxl49ujxasf1zMqylAd8VEJBIoTg1vTGGh35SFwjt/A7I1Gmbb6
6Bw/55tNXG6OoNhYcfHhhIQ61mPZycDrHRzfGScfMmlcQJjkEJwqSvPyqgs2NzmA
CTdHlEnuizdjcJzIYRc88RQULjep3pJpuUY0YuHeSmocl2pyVZ1ZMeqgaaBVy50J
RncgvkQ59BmLu3FhQgzvimVR3DLyIkSjeyCboyN25gVTftfADsNEMekKrV98hbK+
n0lxDsMsWycUTlLa6GIScMT9m4dDQmboO9MqqEwMi3urzbToKzOGmONCeqFVZLxH
GDBSHGX5p4sz3fGVwbqZ9kIKrVlMvHUkUfc8QWIXfhKLk11T5TtDagj2gmLQ3If1
t3YeT5WjTaAJaMLKgcGo7NAOiMrzix+chgO8m1rcbhwuIQ8iWQBxdwKGtqBlYL48
2bbElvs0BiacSPz8m6QOiiAkRRoI+SMVvyfhhDOrZHc3jJWLpClCDO5uPW3uPTEh
oyZvcnKh0+E5Af05oU5K8ed8jSalAufjBMGw88zqOvP+XmnFStsNMf2VpkMpJlma
Cao5oWxXrvDkp831J3rKy6zSovHfwBKeJ4WY6+Gu4pZKUw2BvXsM+ZAH3qt/IW4r
Bj2aGQiWtgxYHIVrGAi91qbK4BYC64I+J/aJoEUJFllzevZOwqhAClvhNK/B71v5
hgz0iBJ6X9NfNH5gh8VLT+WoDLmGkmkKlgEpZS2diAfBG8CdpfVRnRo6YPt0Fy3V
gL1TvUGSiHLrFASehbcJPOgumn7raAK3fOCZ8u1FOf/A5kIYMjZAbvNFIt/FyUiO
4Vs9pBq4jHZxYE/stfWbtNLsW0mlA+0O6QVGvKhtUTCw/EdtTKhQrHanhHubOjec
UznyOIwPNSk7OnOpdcKj+Dn/WEI2A8UeilJdews/yTNXFzuNR1J7yXM1kZx5TuFL
uYL4725lBIOFViJUFYs0XdZBRwopoq66NKspBqYXjeLR5uDOf+TSnjCJbWFnkKEX
EY7dIZ11Oe3DwXFmVfPV/6J1XLsI5nHnjRzyFnbe8ZBsMWk62g4IYpH95nVVuFhw
mtuXCMj9YyW5CTf50wQbG+spUIR4C5IAoJRWyh3M638/TOoCk1W+l+AbifHSqeSq
Sgrs0lFq8/DFD6G/3zGO3MtdfgE1Rzoa28qga4wA/IiiV5YWsrIY/hXzH6/GyUcr
+EwO6kQWJZSFlpD8eOhoTMTSGoeuumdSU7o9601Yd4nkKIsEbZVk0V8ifA5wmSi1
sXj0oINj68LOTTIO5pCRnlISxO4gqqWk6JbYZBEKEv/YpHDTqsnX5WlPnIbmNHYX
acNtoRNwGtzfT3PgwEjdx6xkZ76LEIx+eebcvkeNib+ttSfAPRtn/ZjqsGFlWUyK
+g8lJZz/GT4ifsSVjDXxezHCUYDGRKna8Z8dcKudzzVoJgU7rLbSCmzNiHLUmiR0
cQa6HO6qARrJU/utn2u9xEKIcLJq9rp7H2VMmmxZr/bBuIi3PEYm5a6Lh8YJlfmm
feIbr5oal2aC1gYwYMwjpCEvsVd3SqUF8VL8Xiq9EyQkcY2Seof9/2IQ89TDUMxU
3EXtSp2tO2myFtnymov0YmOd9NCd1e/KtR43Xc/DymYV4BQROTkx2mbRmtZwmQ4z
+DtNNe97QcU+vwKiIiowVpXMM5MHWC3pNZ2AJ+c9qQ1NSFwBqUuOnvtBqnWqZaZ5
TJqCq7ZEBufiSYzM/0J0SDCntYItdnzwbLY7Qba9gBOsdM1iTIAyLfjWg62DILe1
ELwO9N9pwiV5t7EL7C/nA1koFGWWud+YK+mzBIlDFL71ML2XjyQjY+SsRFqmLXNT
KZEhnfK8VebYNgjNuDHyNPa7UCJ1jZYkYzTgQyD7/wczRIngDUPMvQmgLGDcjO9f
11pnCWTajKO2lna4Hkke/vbY9h+rvNfz+xM+uUA7zIlqiAwgPyPrIdRT4Yi6B5y5
dOypgpVD/TKjc81tGbKC+v1YsLi+CVQwVbfAzL1hkQIWmhCq+VcXii141fvoe34Q
cdX1B8S1HcP4+8ewBSMg7z3dCvnjZ2SxyRjcFzST8oreewolv4GrXkoQgXm8xMz9
0Q9i06lT8gVEYKpjjd8v3jLhf9JXb6uX5gwJ8/0OcnM7RY7P9YIHjuguQ1Qut96I
qlwit14/B0xBsNBAsCmC926j5mesPmQ7bha/RLxof5e0VfNmM2reI7G7YnPHRkZH
Z2a4q+bi9V7sAS0zzAQ1w4Jb+UB3B1dlPjd1oJwRG+FX23hBaXFJUrztDedybant
yACBzJ76qLdiGUTfH0iD1lSlZgyAr1ConSRfOFbd++KxBzJxtQ2Ba6jR1C1TcOg8
lJIcXw069Fjr6/c7r6PE1sgmjeDzfVfOTdHTkGe38cdrYTowyCSSyOHnUaS6pGaI
0EkBt8J0SbxVleP3H2Ff5qL7Cn4ZnYo19XDZTgA2ZQvMmXtXQjzh2N0qntxDTPfY
hTMIp+9mcJfrIus2ta6aMdVnOEhvoLeibla37l/lg/fcLQaB5wQpAwLB+SJUfvtm
emukHowQJQyHXKVg6Qi+c2eA15Am2ShMvb40qp5CczTQdPf2wCrZpO/cEXHiOAhh
gO6iqZNQ+jRkZntx/fhyV8VdBo4IddlZa/PoFbN0kSLftO4Jy9MO6s4URfw6a6Ur
2XxQCIE2U68XRT1HTdlXg0Qfn9OJE/bEaa4aoNKL9jYMukktJBWodINv/qCAwtYP
ylM3vNGmavIWc2hNoFSFkSb0yOJXipjJ22RgwoVI9BIsXkHxSzBK/rY/D4wOXlqw
KykGq7feWDCvBy5MXvz0aui0XiZl2n0RcTika9NiNkS7t6fLiVQBJsqHu1h5iRLb
p03edE+rj2nZoM6y8yyhkQe7OJKuqNzVgPED/pvmos/ycGVHuDkgQD3y8Tex0UPo
ZlaOG/iU/brlH07lx0cxMOaAYK9VXlMKmUXyisillpw+kOeTCKWuO7QAmp90ZKmX
y0AbfeY0BXSoG8awyjuyJNRqrGFfVO4sRfevvYObs06taC0+wf0x1L0k8w4IrU9S
w0ncX0jWOwlfn8Ho9TwHPkfbE5BkHrek6M99mSoVwfxW930hUCXCKZHP6YQofyXX
yTdfopTtOlbHNZ71F+czOekJzKYt1gFfzN64uDBHFm+OXJy/igPV/+hvO0DXzkAY
b8ojKlYGjfvczY5Qfs6JL9yZY/rD8ZH7o72EUkwojnggjfmALe4lkSdYBYCK1k8m
8hxu3u+bf/DSo2EORddaJL12U7mUEMZ7jqCUuye186SvASFY2LTfuDLLOq281jRE
ivIOmft0YDOK1ATykfIox8mOB/vwN/m0cJs3CO0qWATmKUB3SRyG/FNcgHbpWJbe
LpIqNqQ4ckurqyBuuStKKJEJRrsDPkkqx+jpBhJuhLOqO4ye6Yo2t+xSMu/0XdJY
wRHPYfiAm/TuyW97vzZ2S/Y28I1DYWC1Gmy/+4m8JPhCyf15Lk//P89uD1mVf41r
jkCv3ifhhLu5me8fANCUMqb/SPt1OSshM2Kq6bJuIaaDRCfFdNmER5xaPkJIeXMO
3eYW5X+wgJ/rQWd++vuWK0I0ETxtcKNRkpA3+VqIWL9ZyZcYyRbrZpb2tr43NPw4
N8UJf+tp51U1oOoGOaWcDsnJ6ufhYeqXgUPg0BDKxfEBlXPsXSxDTMXUYRLoVzEj
TvYhRekrBIpJNgu+vA8KdbC5nX79UKPNUUsPqVY6e9EIX5hYhUUVZPFttjVR4Jm/
4HpEmJ56K/akaQp23janlUzQ233PcDmyckIX623oUsfzvmHMAB54jlnwDResbirl
JRTU1XNOsl+VmskLnxz2y3bru/tcPhqDHhkL76Q6IId6QyiTAYebR/cRe/uPDMiW
zhZuGKrysMCB5ZvFtY2bW5BIgExvxapYcvQ4nMHajCerIkwMKs3+Yhw8Wdwo6Llk
5w8U3tZ5gYjL18pTx86e+hSCN3myR1kC9nlwJfgPOjbFoiEDtLfGuhJtGafadsCU
JnsCd0Qo3IXbspgfjWjcl2kFb8+j/s+PJMETpdgT6oJ2a5+hcP6qIsWweQfstU02
kkruW/dCsHW9bY1H4hrh7L/vMOSIvOdtSRQ+XqIH8lPixACtWvPk/6OGceVNzlXe
IOt4dP0F90CZNLzwYB7mZfhN/V2OZZi9UeRWLxSbwJ0zY7knPxGFbwUNLc/KOovx
ds/3t5shkSjej0nqBHJAswngnpLElGEfaLWjNrraz1go5qJKRIS3TfYXRq0NCY/e
kmzhb2N7MnHsxJzDo0nwmIBS5EHjifi7lzxShDQY7WRb3AmZgiXiKC/vB0Tu5gBU
F5oIS2yTRfS+u2Da1wdT6Y1RxiWRnIbFPAsEmT7CGcupj1R4ExXnM75g1fHrmn9/
F8kZ8wesSm/sH3zkZbrJ7kZ/Z2svk8hmcK0GdRm6Fu6HsfWtQgbe44TiW9oyQvNh
fTmKF4/uXL9XnO4rWl+QWndssuO+EbAPquksIw0sKcz/k3v7d24WaIvk/fGYcXCV
6yRmp0D0cgK+FqjWd0XhE4CfgQ1BE1nz50K82dwBk3hfBp8qkod4IQjXPbuSeztj
IwCT/i16zP5emWrNjjqu7T4z/dswsZKsRchURp63Bj/SmrHylMEypS3CwQYcdHnL
aj+UtHr0RwjpYyW7G4kbkPIUWivr5C1LAe+cZMzKBnNX1SJqnl7YBSeHyU1JHVOv
+99Uh27AvTtiT9Vmd4gQABvjN+kh93TRpI9nLL9CXXcyiEb1DHC2Va1iNgmVdJCa
vS1P9Y30MOP8vEhXctVXUrgUrMd6q3UKOr6hI3rIuIDXoN5E2MLvBmx5oygp+L2X
lEE1sUTN2Zn/FTS7UhSG+Iopry8cuSNQx1TGBcoyKTyk1kGc6fiBkSRLZfpuvcRS
wMoiiI1AO+cloZ87ZPaBSa4TVG+lzO5dHfvY/L81ueNUT2aRYEESJYZaA5qQFL4w
5AsH9cGMWKlVTZgIrQcFzwW7FmjKUp16C1VJ1F8QQ1htsZrk+es1JXs/JrnLr3HP
TJ1bOQ+PZWZacWcbki2E+EIOv1DXjudZrXHQr4ZJfUmu172EXiKjs7SLKbGW6hKN
2dM0O5Je/kKSKXW4ciBFxmEAI+HB5DZgZrlN2cfTgkL0BzYCY3l3iwONqXHgANbe
nZvqNKQSJBkoS31Ybmcse0lwlAqhw/Cb9ko/Ujow+5wM4tZ0FV49RvnvkhkNOEu3
aaJY8KC9zM/jNZX1RKQVCWmj0Yjh03M7atf5H04IdugyHRCfRnevuBx3aBV3gzJ8
byBr4KTBC83T1VEAY4yMeX2XkJjx3GOn4tik58ll9+0yK6k26qyp0+kcFRZHipA9
zteJG/lhhMSOUqLCGYlbbVFn52bpKqIL6PKhDkWAJT24E0YrPn99Y0tui+2iGadY
erE6sVWziiDU2X8OzZJVq4ZBIfD9la2RNhQYeS8iIuGCpzUJ5ZvTB87hwOiMOLCv
XT7dnKzdC5Hna1DdkvfZt6MosNsEZrwOAxIAb56lWe3NgVOwBTy/pIHLtP6S3eod
PRdlhX9puCDwFB7oyQCw7I5kqIa5ZCutsTqR0o5pXvVNk1ySCHAf3t5oQtNDFyaS
tFfLIqMXEFp8qxwvlGZFejIy05YM9DCob27Kp0fGuQS1ye3NsE6JPNYWhMcnV09e
U+3/gexBIkI81wXJ1tjni9VEOOQCKI/s4+k/A8HoXCvUl5lPY4GGvqEJxsN0TatS
29vJxqyps0dLt6pNeEsivGDpH9vPdAAIIOLKm1wiDVZpWWg9Eyjl8SeBa2NbwZnO
q5PoBr/fMQbMLfYjYOvi4C9qOEm3MdMxQUnUE486H5jdC4ewwVgXZrivmmJuB1Iz
pMNZyL7N+lUYLNvpk6qgNmmXNdNImU0u48x+yBEvCuvR3YLO/LgDvRfOKa7CwL8W
pOKdV6wBHsTdMr5Bfi4HZGcgWB9WakSs4ggpsfeDhRODTcChuNzegcKa49sgCEIJ
ZM/emKhkJ8LSv/9AkjzcT+F0H7yvGx87Px6abIctnnD8DdtOgk700tr4+DdUWvqL
UkrneMedEIhsaOid5hDktIDUZcdhEzPXLBM5d//2vhT7qPZfaTdNNvIOeCDxFP96
VQTaEiuh476Ch/I/4Owk5xqlo2PRf6o43LVJEAbgJrh4dyUjc3aWRzr6EtebaGFz
zRO8Me20WXQtCKb/D4E9JZZGLOQ6KgHvuUtjRzMWfCEfDMQ8+upOujUieVzqGRzw
QnooyMx6u0V5RxTkh+4xgRsA5Nca1Tl0sTSnwSEjkKjzK21H88M5u0MDFsvLZGBy
yEcE7wI+KkCUCkFBMFerIdYuWOAU7V8bJJrAeUU0wRlTBnZRwnA7uhQMAqkD+Wtt
b76F6uQe1LSdUD7J17rvS5Qs7ICUZdClatiHf8sWzyzcA4BeOyOAruL0umTR8fUk
qMd3IZpd5v5XZtx5mVETF55IfWHOO0qY82wGB21lRXemCLcuClrh0ef0P0DrFiBn
nkmK9oMw13Hvd7c65ifKcFnjgb8OGWhwaL9W60JaZyMGY1RE/84hDjZQBlVVAm0U
FaofWHyql5q0BaRKNqEVxnwrnjmPXKiW0UiSh/W+YNgAKAwf86x/svRBK7jlIAiV
c/zymbYxa7BM4SOAOpwuHj6TukkA44ck64FKFcBBGz8TgE59k4wju0+ZIWQK34P4
D55Br5blGIyv1aDxtQBXhbNvtSMXZUcvI4sLF3WfY9w9LGvuhgkK7trzx+wHeJ4r
XtzlpIBYfDi96WiJxhyO65bOVOeWK3myN9WP9o0QzAwwAnjWTu19v+Tps/vRn0pv
YnZtvm09epR5LXPDqzC1q+3QGMOih8aSLbRSD28Y41uSoCYRqxZIinDDOjhwpaIf
av12VyHRwcjZ3nG1gbm7su4cPAXxS3uuQjzIndm8zlLHAZEI25iigCS4C03SNUOg
WRZ0eUtkfMWpjcoApnknQx9gDMwMZtGOsjpbPSpPyPj0wz3vE4upopq1fYtikeuZ
4U6JH3Bx2hN7yEPRLJUFIp/cg1Dzo67IV/ZD1WY6y/31qwzqRz5g9CcAD8SBxCYT
EJcjpwNJMxwNJ+czNk8LiBvkYWSB+XTnEFWFDABFAexjdCsZ+TN1uDJWhOmv5ICF
4ylMqgDU5vbWDCDkypRqaWWxl4RlYolWNggSccFoUyWyzj47M6/LET2Pe/iaM/Kd
svs2ZHLqP3x6YN0wWIR0OlCdikjdVsPX18AiGR79lxwpQzHIOPSWtgd1tOXkXfFf
fVeWlS5Tzc+Tev1OGqu9CQg8mWX9Xrw6ydyQUxX/QLL9symlgdjmZJxk/vX2TUf6
21btyNAaBWN3kNCclwwUnJH2jwpUh6Yu2zer9bUuoRnH51AEYMnzhStmb4pIAoyw
t7K5KkMVDbhBJ5FTtC5jWa/cMaPXK+mtDMeMJ6o/MweFprntzZx+x5WYesoPZmLf
zXV4ga7he9TtZBEw9RldMQVMt9UCDtkiqAufkakB07tbsjP6QorjFrgp31ICPwIx
dVeaNOIM3wq9M2JHJo07b3htmwY6IjpvccBYUfXyjKtyfYbJV2jV5Z26nIyJCTZN
9CsorofQzM9XxlXqRZJCN7DyloYSOc2WBgefWd6jw5+gSP8FUeGw1AEmu0tykb/G
ODK3pWykzItvThlwBrQq7kI7vsdkEFSu1oMQ1GFWUVB03kR4OibGB7LE56lMYIHo
E0SWO8Jo8pERVfXBGB+1lBTR7AIphxAKML9wyc+ofyVu1VYvHdfg4iJEM+BQ5sHK
IuPP1pwPs8osN0nRtfnLtug8pVziNyUxiKlBSkAp7uT2VUoNh8cAutZ9OgxDqQwM
GKSEILIzWvQfaZ75avdEFdEG6+NeOmlkgwakIJi33ks0+NTBFrP6wIPzmHsAZgV8
GPtxlRSCHY2Sk4vn0J7nUbLX8z1zykGAZTI/hmQ6t4dsc27icxCY/f4HFopDqZIe
6m5JfPxHYLGTgO4REaScZDV9bp/SMZ/r8sToFTRfgHA9o+mNY0lc+THx6HevFYIF
sVBd/kJahI2JyedPjKIVddgxUQ70Z2H7galkFEKyjDMrxtVPcQOmw97SegDN6bx2
oc2ERU375EfCLvjh5A1kGiC7PRLuw54Wl9xl5pCOwPHLvwv8i62+Cjw6H0Gsno1M
VU3t8w5Yd2n8vxjcCo8aV0Lr0gjUdMOuYJ5h1H+tnGr+rh+AcePxCDJAQ7ZzfXsv
uv8IaQPwqSuILI3u2ibrCc6yZzCcT2Ca6ksjey7Z2zKsCztI1ExZ9+baOtlc3QHa
i6ge8YUEMTreDXPut1r1Qif+ElQ5jU9+WkBRfnPwoXAHiOVlMhjkTwwiW9ZBvr7i
Qi0IQ5HmEUBmDdkhiTtaucyA+Qd9CP3m88QG/Lo2F6LAXf5zL82G2vMTSTr+c4oY
a/lhVqTVyvTKkYpbJDfdJWu6B4TMXMm0jaeBfp/brjO4SA/k99Q//WYmbf0Y7lhw
iBezxONDkMVA04StaoH2xJTzWPpuyI/l3AjrWswwgpglHH+tmRkwNTjWcB4kKccL
pnmFNohEWdab5zIgv4VCsK3/wcLV7ARv/Xc+K4+sV+tv2jgKhsFfCLMioiQrBGLk
VWaA9hYJN7YGZYC2o0v1pm3a/WxJWTyH6Cdix1JTOuIu94ll2vhfIyRZCgIFISSa
WFG+oxlK+YyyWcYGzYdaG8sgDJPB4O+kSGdV3QlQxbiWvYqRRxz/T5s6Snf7T42f
fKddXA7e1XKELAaqidm4FjCFeL1kbZvl3LofTWizlqnLY9m4W0J0amg8/3QV/N+V
8fQW6ry8ckSMte3V1twaeTokw5n1ia8oyBwXHF3xGSR5PYRQVCA1rN+HGDl5IDzx
XU9UoOUGPzB0U/CmT41ntMpwFEvqi2UTlIhy4oswNzOCzCg/K/klQZPyFeLqZDB1
XiOqc//kdlVDrQzIujLN9lqzAhFh0yT3OcYEOZe13vyA88rRoGuJXMvSS7coLCC6
IoRZaWdsl1kuGKclCdniXB1KJbet5/vNnEn/cs8SsEeHsYWml+hDXFzxe5QscUu+
eqOMtEojW+hQAoWTV9xCYUBXn6IQGcYT0ReaCMfM+t5ygQ/g4VejAevJm/wfIMk6
j5EeSjaaFStppDg9EPH3tk5eBh01YDoFxmD0hitHpvUs/FwnWoC/hqANNq26liiU
`protect end_protected