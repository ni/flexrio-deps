`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23952 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzkZGdUrjzQR9gfRaWjj8jjLnC0r2xMGuH5Hj1kHcXX/R
0TP8QdAj9nl4wBWjTYRg6MrcS3XMdfxmc6pmcGbOs1YODjhT5/bLC283lqyoVxjK
cSK0sWO+l1cxQQ+B6/2Dni/g2vHzuMsVRD7eXz1rZmPnGqeQGapmW8vQT9JKTYw1
nVOYDYDcEiIrgNP+Q0g5zQxrJ9AcgV1iLnVZ3KfxeTQzUqnT1oGUx/sa2GZgt6fO
5YztWcQbmiVh+E/R4Hu2Oo493XXJz85dCKJlxtSdBtm0AS/8eWPFBU9a2iXtXT/j
H4wH5OksFgc9zomgRqAz11LYtfBBCyck59ZTWuVp1Dvk9W75bKFogvVKWae2y8IT
bgb5qyRklebo860IdmVsz9ceftFobFpVkMMqfLUY+glEDXgOqYKrFpNohFoqPbYy
2UmlEyfBm+Jwfemse9VDTGtw5Mv/ipVSkN6Q93wTXqANbjw8FHBAcGfc9idk6pg9
X//t6xzONEuzdLuFWWZQ20YD7slCDEajf5EZQZIN4INp90oJjKeMycuw4CfrDP5Z
Z0bSXhs5EFD55CxIy/RDGIgam9iU2vI5atp1srJh1I0PUAxRYQTRyb/HPQrJXanl
aWDH+zaR1Ie7qtLbbWLjAjVF01zx+jriF9WomNx1vom4O+QcNsReJiTKPVbT7D/0
KAgwSxXqccgyHK82G/g3rSZSMYaVxFgfwNyk5WF4tDHiiiWLlzEH4V8T62bLsQ0W
7HGAPjeDZtBhqWv7QgNXBE/13MSVLIQNr6xwNIfhI0ET+GlcJx6af683whpa71Wo
0Rf2cgXVxEkb5m/0ySDiVrFcoK6fmAiiEprfkvbu1SNbbe+VYdqJDEzqRDXi0AnS
VMgz1GfrDyv+mE39TyUVLEz25D94gy9FI6OJmu5uo0XJD9bUL7eDyBnbpJ3STcb/
tc16eTCczzJ2aJ2P7KedLsjw70+NIRHDAmwJfjgdXbJ54SdWB57Dj/qcm4sLP1Sv
5B4pOLQ4CUKEJekTKSe/A/NDlup/5twa6/YQvwycYdu2QhAwhPHPCeuKqVxkiEYg
3n4TA0k43Rbzpp1FwBXnB9VE3tOSW9STFHzYW3UUEkygOu0sXCC8wvF0BXcro8+0
UJt9yVm9sfGAmQPJW6G5OX51lZAxiXZtPSIC8vHPNn82HOZh8i90Vk7/fiO8Az/L
BZzBVOmXNavR0fGlA4dhREH9EuE5WosFkme349FmjHXjREGsNPHm39UvdhtKbsGC
9cG8opGs6Dg7fzYlUJvYj2Wx8t+0hZgRJ3NdRWkSNHETZfMmFNOn8vAvoW8w0Ngj
Q3WGf9G1Fx4zwiNTNKUXmPOnYcQ5YpExwiRvc6ITVrRnwRhiGY8mPBNhFOdDLKSC
IioZSxGzbiP+Dy8UhGCqTQdm8EFYP1bI5Riz33FkhIvBy/lO3sIAXHJS86jDHVfi
4jL8/Pe6WdU8I+lEKYFNBI9ooMahX8epe4ZfJOlZug9lTQTz1iRbdGzaAPffiqUo
GBXV/MLF0vFOssVEYbiOHsyj8lJ2WoR9/b5P4ct3aFdaFDwxhEKJ/bQU8NMQTbgA
TMACWl2Zaq9OEPM9XKut8lnAJy6FP2GLlZCMG9YgeRy8HNgD85mHBcXZF/apVJZ4
pB2RKcYKDvGx1yo4Rc8KcTvSBznpJ36wHrwURnxBksu0mplOtz8LY5DK+DeuyYFh
X6LSycIhVPLNsg/PwgSXvH4YfXmXqMJfHjTLga90xA2mY0xzY2Ns3tmaW825EkWw
mSbwSz20f0KldhbreH6d1EQvA7OrmaO0hWFFFsJuXf+2oreli3agDaS4xFCXoOFP
QDB2iaxILoIC/ObXXNqTVd/wYPqNgrnVn+68ABsAAnQhNw3C4pwSi/Sb5HQR7Cfz
JHlQQl+xjYXkOEJQiUh5YKq9I6NFRGpyaLi9+proYf7BhM7KosejQcuMB2vOjJkk
yyATK6DHTR334H+Ek8BllS9e724blLYckD4NVKQUpVbrtehsCZqRvMM/mn9o4nGl
4di/zkibfxLTguNZT4m4+ZLwNBNjIaT0fb9Esc3na+92MN0kufKaapX0ZR9IR/3k
SXVV6ceEFiwz/XAJfbQkxjX2oOYZY0VB44mN5GcK5abbdkblLtjFQqb5ml3KexS/
KyifnU2JuJ1ZpBzYbY/F5rP57W0pzX6BxhqC4CxeFXEfDCncSMp2IG//KXHrFD9V
SppQ/WdNyScVqmnoG1F2vPbpUUYqtDWinsnZCTTvjxM8Vb9cD2+707tIXesE9dbR
TJ66Y9GWvZOrPjMdrpdYO7XGUaLxme+Li2+yXCN/5E7OkWgVFnTa3Gfrb4/ym2b/
DSazQyq8SLx7DYDEqjLKIjudSTyI6RvE2Cggl9v1M8Jq9QLYaTubtXJRruHRyyNe
zx+nKguAKcGad84B8Z66LhkpwYFjucKSPImaAgmNrgpFKfZuMgbsx8531zZEol94
InO1J0CVRID658myW0czYBPv4JR3w+Ij9uvby14s0wfqhJ0bPpsX7YXr6WyYlqSp
m6bthCEQfDWKfiHU1uOOPATv0G74Ai3YAGTkAC2csyaSDmH+7VXJnUOqxoIFi9GK
8neMl/qJtzawTU1aQwRMIPlf90I6IRv+pc6c0QXtuA2TwkV1GyHE5dMAL9I/yy6f
pqRcyk9noBJYX1g+VP/E8w3znNumZs73hTfPljvf6V8KrqkG1HL1Ap2TCVVpgc/l
rK0/l7mQzomf0I4n54WZrsiShZcaJgkhrpvGP4rLPbG46Fd2D1TL+WKcaOU802US
Jx62VI2J2ljzqxBn1kIMHpJY2Du98Zn5ef/pmiWhQapT55m66JepY0uICx9Pnryc
Xg5QGBkmtKR5nnXgZgCrzhxv1Wgar9hS5ZF353T9p0+GeajJxsRhY1wAWhti5zkQ
l5IXYGbRcAPRg5y3uHCKpgNM4eZ6Mlssj303dsPsPOittalwLT+sgRorKSmVkapz
k1tGu/mT/Uu5U+PvyhenliXIyaBxeUwItjrlwzgf1liLy269XinRJXHTqGMkLhDY
+1V+C9LVQSaAK6HIyt5SFoBdHVMWDh1+c8qt2rdrtHsGulEyFies7MOVMkh23kss
wwFrbzJuIqGPjt5u1vo9MybPa15wR8Vagpu8nCus9VtbQqab4R7Q6f4IX0o83Jo7
f1RFBxckgbzCv0ubZL+sPwhkb5wzdJAwzo3DKHtcA643/wH5eyqdgGQjUZX/kjnL
F22y77/lPAqFiXZ82Xzb/8C5XgseqBCurZGzDq3B7KG20PtGnImvE/GoGihzjJw+
dacXvLXpJOCynx2kVWW5/+qxR0ZGVlULDfs608CIWMosSGy27nrPVS7/mYwzqx2g
+TvztdT7g+3pm2m4YkTfbkAxC1Y0zFqLl5aP0pFjWcf2LFzQLrDlwKmJv/gEec8d
tZBup38+vUWXP5LSOJ8f+SOq8q9c5/W7ihKDTQ9lcVaYFzjrPfEPd+88JkkcZjT8
d5Tk6mdBdU6cGduek5JeOkYnFkdZoWJSAxp5vHe6ZziKl83KyTpzd+3oQjonWpka
dCpQ/gARJMxShTdsJu4kkPnGrycCOjsDjXWxEs58gTZ2YLtupLhh6Phsd5XmgNQ/
NTPURMd4Ki5E2A3HbHrjO2rERSQxg44adfkJWaj11+atTcAEx/REaBORUPWujkU9
3zKhhK6JtJ36bu9L/WrhZR6CgzEwEltSmlQ5aWCHnetDVXSo79piW06MAA0XRh2d
arbrXGyYWALwPtCR+Vg8R4jTKJfluWqkPc9WPlTobdx2S05YgY0IYUgl8GZ1rLc8
qAsvdlmBNcmYDVZgGz7jAeL01m8r8dk1sNbcWLPU1shFylCg4OYIh5fsMIFkP+ws
zWj0B54YYuYxXoPNYnJpBNaG2HCCEb5QWeFFJfBJkneTVGitALes8NwC6C9t8bss
3USwtPlqUcueVR+QVN2eho0a+Hola32Gbtuiu4kAIEevNNwNGHk5SNh5xJL0l91B
osvqQoZK13RxkaIRHiMIQzQCLLUxRtyHephlzPruFoPqoQitQpWesHT2dnsc0mI5
is8ynxYJ7i1ZgahpXxgTHjnuzsPETi5iL/DHd/txyUWhNua8KMXLSkTZtqC9L5qx
qNU4doUMZ0uf6OCgQ7YJ31Q2XYRglz5NMgX1+9CS1acxffYumzqV+AwxjxFCKhWz
G03WanHONK76/qhZAwyUlr3SoGwk/4EnwQlCOoVU1zaW6GcTPx+YIOczGvN4GjgH
QGva8vq3hazcQDKAOmCAt0dDiZ6lpuEAsz/A6S8yFCJnZNDTULnCvgF2ejMgBbIq
7vjqpXFXm8wqLWWq8LYTJXpRS28MqEC2Ux77gYdrH1LQ/Vev3Vhza+ZwzPk7oSeH
BJ1f62iFFKEzz+ffMDOhEE1sAt2BnMbPH9HBGu7BP1QSllLvRjcDs5VZICnDxR7N
7vUQbv7DiYrHtKTV6M/lOPsfMsFIWQYNTVFB/X8AVzAbr5UzoG3S7MP0A8FgIrFM
vQCabxLh4U66FOSruIeo8CtPVLlkofRn13m+Je7RKI6Vu1A+Wze6TUHufDFkULY9
uKcmV7NDAEDu83+cYq7pn0MwsK/x/Ne8SQ0eq7f2eRADdYUw659iuX7tEcalZZpz
L3+UFNZL3zuD7yFO+ZJpx0wwjMFG9ArP9XCQLTBH2f0TqfLZv5sS4QiDglsmi2/x
3dJhiA/JQbGKH1KINYxQDrl3tTDBFusUHV4i7UyEA0SVmRK+CX8/tLwHipx3at7g
TxUe8ZVL09yxkf3Hp26OodJoGMVZ+p94e6u3rq4/ClMnR2chW0sAAOLs/zcbIDf5
K4gL7dciIHQIVpBneIelCAcdQo7Trco1mG24olcbVE86JLHgBYPBYZzbHexgERbN
TSB09YHMWnRPglBsaJaGb0YQX+QMuFvGpYYjfQJwC80oiHObDQRIUP1+s9gd61y7
gG2cHFb7O4/WshmfF3JJ6UeBJA4M1YvhXIeRCc+RWpmMKr666qx1IXXFh+rMhZF/
W6Oj/j5pczCMYF/T5EbQXP2og6GKjdXkqCjSfjg91Vnl92WRoa969savXZMPp+dX
oY8CpAQNDB+8JxWl99EPtCXhsR/C4fM3BKr8xIhsbkgV22jsAS1lN5YMPvsOLsW+
0AbxcgufRyZs7j9BlKmz/fVi4lXKpTCOnXLwbijnDdKb969CSFde9yINkNTv4VOG
/VQn9F+KnvieOQtxexN1x5ZarSlfnz7Yr9SgafaeFqV2/zJgkEHl/ACeF9m3+whA
5Ia9spORNqbZzKGPFnek0sP7znZSsAi/loABOhRAnwDRs1qf/z2egpBQXPBTX6VH
suJP+9SsLZQq/Hzdntn4jJ/3KF3ugUz0v30BKhIZszvEjTsYHmPzqdK7VfdqfeEL
NdDJ3wtZmMjdZBHgvSobPtTCgNSe5/jqXH6Z2kegm3/iL9qRLFD3XJi8t4z4hrKb
fvyWouIma9d5iLpVX1l6uSxaeeprUnOztXwXVWE2jFte1wXKQxO3BD1HKzz7TG8/
1ooDzWXJSiVU9wHzx1m1YfbvxNt6HCb/NCMyZ1QNMI+o5NjTP0NjRo1XdpajdbUR
eCubWLJvSo3eKyolb369JZn/IKBKZAslbOAJmZGfLDPLtPNSgMVt2IisubiFWHD7
0WUrlnmCiZ1O8LRzucvlJY6vXOJi5mNBgIdrUKoFcnTTPAVAdtKAqMW13uh9coPa
813EnwOJEdjXWkVfRk97jND0vWa5nBFC3zeEmyLHjsjRXj0aWVbQc10RvQEhpTN/
D/pxS4gfIiOqe1n0qH4VeHK+tSJkTNsWShsuyO4VT8KfPgPshP2/78WKzmSjGAis
3H/ImozH7KQxNfV83DmcsMzCGnuVU0z13PrVHPiRWwILxYsbt79DTo9jrAJMqXlY
wM9vtL4ap+CsJIJ4BQLiB13STTCoHD10uRyt9fa28HqTuFjyDdaKF75cU4I9zBm5
NKAQCZEktHR1BCpYJZiS8bOgXTML3NXllyBQQRAvj+xT0G9bL3a6mwOFipIaI3ha
w1dhYABVBPPnU9qL+eWshjk8yNSdjWdCbC14RN0lJj7UVXjka9LZCgWOpXbxgL7V
1ridN2ix2wpqSXymEXvUDw4sn2thdsdKGeOO4nsCWmweEP/BNCCQ4x9r2s+Cs5CW
4Yg9aB3ZqDchCGmESwn//Fp/C8h8Tmrtmssy2ovkw+HKDMIQqNuK/i90f1YuYXjA
4sweYUJPPgil6yJ409o3vocIyQnoRdWEkULjQ0ezW5oAVnRPNl1TevrJgVom+PNT
WfUq0Zv32qAFyVC/RgwrrPesP+nL3O8JlJr7b184U9ZkLqOz1P+OYH48RZSy3zWr
eMEVygsh4Fx2DBWb3eWtSNkjpZzy3WA60TPeHbDHS0O7Fh3naH8aPwffiOhUJboq
FV+Ap6Ve60vLy7e6fzu/9BEEBoz+kCjJQrRbpsexpxOQ4IEXRkaPEqOMUCMWxE05
Ga9lqsqFzBFQIP2DkQlB/n4tPat/5Bfm9A+tWV+HH7g3BABOg6a5qSWrE/HQzPBL
FvHgtvMWivI39WuD4N1H7/PIFnb8baHAK1WLRvVnFhoi+ntsuNGwzYw/Bc5mJRWb
V6Cqx/xp1MPHnyL9K6L5bHkpbS0RGxulgDRsuXl7YSH69HTO0L3HrgPD+kG8TbN1
+DFSip0lDR1AqrDGXBk8AKvsz6mvlGH0Oq6/V7hpCBOJYdMRVi/XPFRTw1uOGGg+
2Uroiy74M0Kg3SNTU+2OqxtJeS0oZN/CTAIzUT7okb28pQO2aJSqcY6sTelpOvLx
rRkgypSHv8geaN1ecucYSDhhEO0wQrtjCfU76i53KIpghhfNGbKghbHuVReZaxzM
t6rZTyU0na9vlW5ScRNnMVkvYpriMLtplsVGmQapnCAMf6M6HZ7IiLaewNviD9ta
UY5YrkzrYVNICgT5poVvBEXJJWAcYmBW7g+N9jUwKdRwVlGXYYx4Q67kOuy/iiGH
jNlrmdNmMpvsnXOITktr/6iH9y4EQSvZN1GEKNjb2w+j30t7CprChqoevXfnGNzM
57FX/sqAsNoVcfskV3N0ZvNT4/f+gaj5RRLbH63eBIZRDTc/hMV3cAzPszQiAecj
sjItpl+dQIWmgBit6L6XQSTY5csZOd4WxVIn3h+ySrEXjQNarVznSmCd7V+HjEef
9q08hUy1Fu8sBcDYX4Zn1AwTI0y3PeZeatFZyQeeI0fzj7WoYP5vFx+hpKm0brIk
tQ07xHZ1w+RPgIhpvlvKgZJ3MWUWmTIA9FlUCVD21UdZ4siVyVKK8c4z8Rvy889N
znJOZVbG6W75jua+NmZRwyPBTKh2U3XLQv2bg8m1eP5pjb0mtAFeiwUkCzdrVcxk
SUuR+x0ca0MBifosl2ZRPJRoJiIMa23/uu5XBLnPYv1S7KidoyNS/C5OQWvdyidp
xLn7qkNHfOTDZG4rDlaLTV9ArMHNpCpMUcfXqvojPfNV0ZY5HVEpjyjdI8a/w11Y
isBCsQFvF7oGouFTFFyWX6Y+mKt5WomRflMqtXvaY4312SY8ve7+h8xeIp3TeHWO
DE+W7D6gIXnEut3FfP4esiv0mkGpPmZBjfbPowiFvFHbQbiHZgqcBiDadpaA/d9F
w5V9nAuYO7GOtMi4vfn+UJvLc9JzBK+R9YfEo0rDLhMe85G1kDEHq01eiRYO9bBo
D7T/5ZpIxdPZsFTeEnDFsY4UAFa2xxu3pEcoTuLEcBFAzt54Xs4ZDsxnbGFi+40R
tP4P6g6/HDOQEhg30qGWkQk7ms6M4YZPnA1oLMr1AeJDUGXvFAFKN2ZA5jIn1L5m
GtVTwfsG11cU+wIF5y8fIZorfhBSuqL5O0wKNC90K2E1LS60kWdu2Qt1x0gJMWqO
ngER27EuSJ6Z6AC9ZzQNK6HeDwJNkuVfVmYeOFU8Uwf9eG9feerZbjE8giES+PoM
4tXZR8aLd/DH2qdIqnUO/UFMa/IfYKZ9uLRIEIdVp3yydNnPziF0XLb/deelbUTD
91tEg0L1bRYYiks5SFN8l+JyaUdy9l0JvJ6D1YuDIZygECOwpN3/qIQwV90/y/hE
BiQn5279ulR3A+M1Jwmae1fWSef6NhkeZHNbueYyB5wDPlfLoITbrGjSica+ajAx
x2UDMebMuzgRlWaZtlrgC6aChPtHa+qaUz2mqK2/cuNR8kqKC09L/6q92f83kNZr
BEQh0CrqhJ0ElPVf1l1ft0AeGGJa0zAaTjmkraLdUkOiOteIakl/zhfbk9M70qNK
lDganzDV2UqgR40T2KZM0eN0/yI1UDhn/JWN1LJKlFmND4IpxSS4j89wf1aTaQzU
IVgZhxogQJ0ebDxJer8IIYHAlzuP0cAEoGnTeuZYTlvdNeQ5Lo/1A77R7anyuGUb
w/bLyc5HipZLsf0in9/rZZk/tUp5Y+YQReu4NthcurJ4o0UT+XSAe/HLLDc94Yah
mmLjyOa7Yn8KwchgK449yNDZwlowGLSlqpuUWo/RVFh5wywE5txCMO4ZejyJ+toB
7CMoY1c/yKdAfbbqZYcCpQrVrfJn9P0TMcc7HmkTEWj7lIbSFQy9Pk76COFC+kBM
q4Ogru3m7dMEozcRB9chwx+2JZ8Fi6GHcgiCKCejb7wKy9bBcfX3Bwes5Q88SO7B
wiZ+qxRFMpyjbawK1e7K1gQJ4+NQAF3dnjnFVRuOz7/TjkcqO3x5dk64rJW3mDFS
RJCI7C+qv/LobadWCTU9yoYGKZ/fdWRYKG/+IwKC5j3s0szYkLeewEvrIBq5jpkZ
sW51rXMCd9v4VBz1OuwoE/0Rl0Cr74LBvRJfK2o2dgX3dix123Xr7f9GF9OEqk0f
cgmPwfqFFtHcJVMbqLDlt3e8Bihs36g7HxUuOOuZbY44BcMEB+jA80TSI+uCdgV/
dwdd+fsVMKYp4260nYmposBRTtwxuIK3Au5ZHv997EBqdeMrRGJm+RSVxXlA8Cq4
YCJzNpBbTy6jsdiayNRLDcdJAiedTvHU8ZIXI2AdsK1E8/x7LKtsIf8bpPxf37fS
Iunq5Phd5y5eQJz65iU2SiJQEw6Tdd4p/X1yu45noVUzdcrvyOua1WV643TEa7nD
icuL21EDLGe6VPnJkzOt1PP75nToRqo/VuIAnPask6CxCb45at3NmCyww1dvyhjW
Dg33aFc3yWChJ66KgQBbJtSyUL6EsyIrjYhZXLGyojtfKstfW9wg1m5CHT+U9+F4
nB9eFhCzW/486U8hvndQ8uk416jnmyDzRbxEVh5rVUmgBV1d9b/LosgJXyRauQws
hyrVQGNYPdIg0SfjIkRdaVNioPdoxN7vfylx0VOH5YhRI5HVFQehSh44S3oFbLCm
/bu40beS3ozGsRAxyLh4yDFXyGqsIkyFbENPCjBBHm3gnRcYhoDgjS7gcvwN3Uqr
pYnbs+zjwPCVdZqwttZhbO7cx6NI8Az9982H1SNJk9gsTgMRePdnXbPpT4HuMpSh
BRFApyIUAFgyq1BZrsypP2Y0DxmnngWEfuV5rplSciQj3husukJ1g4/exXLwQQOA
JGBhSu6Ix7eajHzHwGnk4igSwLsnsLlHy3kBo9WVGr7REK/jyJVyQRSDOETP+E7a
eemjXT0ABTKOz1Y2FP/jJRZyGh6e6b2AWGJIUzrjYgsoC8kV8auBVJMPhaYkdWBa
ltR9wDEW4ZS58qOa207FlDFQB5Y2kRJF4MfC8q6OkQm92Ahs0Mv6QscegzGFTz3Q
kQS4x5kf4Zqkix1u6kssptucykbTcTtjs7cakG9fAmkehn6HimmS2Y9SCe18QC2Z
iN3c+zw5n2XwlUYfOmCWMVpXzZ/1/fVtvGKmgphGnEoAvU2WIiINlNDUKi5x8AuY
mBz7eQCG8Ez1mzLC+W/awjZlXy8UZEoRymYc/toh9k06/FGq7Ru9eu1xUCHnU+mW
rscI5Qit8nMDktgwwv9E50G2OQnOEkxfSXkr73tEhGUH9MUsKWWSqhgUp0XL1Wpp
lU3kpSNgIjwoJ3CaXIbnH0+zd0B6fgCjwvHyRMplbk1i0FFDMtblEDYdVwLmiTMc
iEd4I+A+tqikAhAIsYDw2QoXoqK0TwIeHWr3voZAuOaazFt+gXL93T4cIVhT8u07
dpyxbePnCkysK4W1LADGXTWzj+w0mOlf4hBzCWE0LQAKWPgzEKM03rpMwlDX7ChO
EfqnOYfAiUtWY+uy9p50XyfJ6Q2K/uRH4rPRRsTLksqrwEGsLqXGhMEjsiGOBVPm
90uUpphjPKpPkBqVAyfGsOpgglJO4ZXfhUW7+VJmk4J6obsy6pgmGefPY3VWdqMr
OJ7aXsB6Pbk7fhzrJW+AJ46f8qXYKkYw3vWaKsWvZ+zrnSX1giNcoRvDGhkjYfLt
GP154FBQrj0hAVrL8EhK4aDOqN7WvzN18/qyJsjyAKant/MrdRcpFGf3171n67k1
uSmdV2gfS7j+U9U7ghcmfni65BaX3b7gobOLql52pXnA/qCsIq89OnbHpChReYod
z1Gu6rVYxpp81tNf8J+IUlvnhB4BMVOTowyMvNV4gWzl9vNNPiK0L3qWFtmkCOwW
NStB56cYGlzK+3cnqLoJe6a3jXuis6l//6GY7P6OpMuQU6GPj6Rq90I+g1DvK+Hb
JSAiQBOWJShlLd2JzCZPuR1h0D/KgJ9uE6Fo7UfmmfgxqJZllkDWKQuKj6VBynXS
R179YRgNq3NntlhG9E5w11KG8ktSjh4Xsnbd15qhGKfDwq4uIqaX/wLVuzTmf0e8
wHYZV0E232TiyIYQ292lDTEqlJFXWufpIIlL2UvCMQkQrx6f8CzRMSBWTEGRu8aX
k710gwJo30YFvocUbIUqERuIdwtIIMLcV5oKnQNK+durtzJDDAHaetr72tfdeFgK
AlxDPpvtzKezzEuOUQXm10VHTr9LJZoGcusC9WVw+gZ6jRP2C/TUaRuW/0d1e8GN
svDlQpfrfXp8IE9Y4xPB7UnqJkdxxTPWOGoWWHCMDpJoTAy0pdMwS1vLRtuKlW6c
dJOacr1zfanTO9vqIvaP5yO/wYPBDsL35g2SnE1a4nA1k82S7/UawA/A85B4FtUF
Vb7ALwEh+Bk3wtmNL/9h2mZ8J+3RgDDvxhKLroco2niqA5WOnfA/jPkYle6Nyt9Y
ZBJyW8ClMWlL//IwxFLwhpQVzPT+gBN8LIKdTl6k8zd/qrDtzsL/Ak4RUpJKxna5
gyq/z8teltyUeQRxCI0KVoFkgb7ubRQBIJnD/+BxC955qn1z+ZHmhVUl3REWTihZ
or4OLCbTqLE8xYWatvl18eD6DQfMD/EQ4BOEUXdzGedb5ooLmFSGMOUhddZTjapD
zZ9YrnDr7VqWEf0L5XyyAOkFu2htLEPVck5pE4+cStUpXqldL0XOG466gNtzNQAy
8tzynYRfsvsgvw18dkaZaW2XBd79d2s4HG0x9hHQpjdw8p8oaLZfj/SE1rP1PFGU
FhZoyrjwlhCnvcxK6/A4QFz8j3bHdeFUZiyMi/sffHPpr0G23FtDbAN7vxKyxaom
1o+1tRZU0YsMS2dZwg2CoOnERGjZ5tF5nF0cu3LZvforar3s+L3iQYVFXPuwDTNh
m0ljuDa2MbMIArv2SEeHb8WUC9m6HUtpHx612Td+lgDLgYgq2E+cy59qPr8rsEf5
HC6shjuUevSBEH9DKtfB71rab8E2SkAtxqhToM82UyO83olqWvGDSOPuqNBDss8l
HldxQGgsNQ6LVzzDeroioS86jr+gKQZ8lMOOuovZ4xjI+s2ubFmxiwLp25LJ4xAr
vckXLt40MT7/WZav1PwtwQ/21ovpgxSikPBID/3iPpOovnBD4SorP3anz0wsqyV5
qlgUSooW03Pqg+9jbi6/o7VFpPcIRArnFCa5NxS+phrHJO8+TSJEkltTyDLMD5qS
y42AQXqZg4eYcaaBO4COGeJ02aifYQQguLi4+hEzZJbwNM45Be++5YCQx1PVSnlv
eXZUegJ/fNN1Pt9cUuw788DCcE/8KvlL7oV+hjy21qiG2tUrUgXDpaGaU7QR8e3/
b3uJY6ERjI+564l4afWS79Hiwyp0X0oB5wWZCxdmhTLFYcPlxPBG02QzVFfMmazi
7V4nQb1qwFqvKOhldzw3FP2cu7OL4mpVQyXNngtGBBCMju6DQoPYZjNGMp1NXgg6
I0hqiCIvJZZYbhrm0/5/LGddPviCcS6DxfjQsIKhTTLXm9hC4rerGNp8VfAeEhz7
gJt9bJ3RXrv09x757XrBdbRpURtqYt1zV8Ab2nxbdXmksnlnZhkJVCqwewkkSq6n
Zr62reQ0F/wKRsg6usVyravSFR0TF5ov/MGtCw930AD5sAaUeGiXvBGQ6hTcSliI
+WE0NzKVWi4/e4sB953/P/KexTW5+Z4y/uDJR/NYO/sBTY2gsZiKfVpoF9WdREy0
V380tPjcQ8OERcY66/Etg919N5WSboLLd1uYv84QcmyszdLhS5s1be6ubY7d/X0C
eFzBCX7ovShOy1sD0e2Mk3ij4y00fuSKH1Paz/st2TaXFOhABiEp9yQgOw/2uDyT
3gJLsko0gjiOOPe1a7an3Gp0ybCJeRMyZf7yeJMsu3PeWM9x4f/qIeX2XpcGuRdJ
1wVYoqgmFGOkcMGevL8FdbCYk1H6ATcH3S/ARWjGmyoSkpXfOOY06HCWJLBfrDD3
31kRfo0Z7aZNSNHtsre1B6YthCVGQWG9fgbOsikw++As8a6xfaOfV55emzs9gY/I
5K2p0xPkunp9mpIR/NxAFBax0iySKGNLvhiJ/C9i9vxOGuE1tMGpQDpzD7M2ZZpt
MpirlKpo8mBfbxhmdkzbeqkgEDILcYPjN0JUq8POL39Pc5d6P6YOzOtt3L6pPeq9
L+IDctITCFdm4ICESYmwpSNyKGVy73G8zZPDjXlcKKOXXlwxJK1tHUQpILVHVbL+
lcmG0hPh5WMJxDQr17jNefQrdUe1XzufkIZ/fZzsuvG8aANimgM+H5UjuH+4M+Ug
UdRg7zI7ZOak34S5CMsiUN5U7+MTubKNUpV+SkZzpNNCQ0bHWve+EKy8XmE4unxY
VLVFR3TRUdQIGZ15AqwJ6MgiT9r26CGVVMJtecGJtRECN4KXKXgIP4b0K9Q5OnAU
QJ+hSn98H3k8S6W1O+lREMTVlMFvKnkH0UC38mi1GEPT+j8Ua3CfiCiisF+6JGMU
GTtOykQdlo81xi3ABfgJFBDavnZGtvxwmeoQBh5MMNOmJ9pVgcoxl0nQUxi/bOFL
P+zRukmkhc1j3UqC6nxtm5zLItlm0x/akjPchD99NV0ZHRetfoykqDYoU9Z2d5S1
TIbPz8oZ25SPAUrVCO7iCkVac8ETfgfNp3Pyz7WUjatAbYfwpuq+8CKyBw17hWtE
NLqVXdNjsdyntO88rEIVY1zNPgLCtdQi5q3WElf2Fq4g0zi5OvOyLxhZuUKdyITZ
KvSrlwwhlFF9XMzW7bZKmqiplExc6iXusF7VJ6+9ItRooSj6nYO+kI/33iYk4Bga
z/OH53kXy3+ommkHlRTL/59XpSjV79Db+PB9AXqmxKp2fXyQppWVuMm58m67RMXl
m5TG5Q1FDYiJuD+ZIPUhbOc0e+eFhs+R1RzJFDfgtP3gUbfkEkmB59VanAg2dKGe
f9LZ6AG8ou5FagvT+tX2F3xnek1zPatESePlDncLyg/HhlQQCo52KFug0jgjPQ++
H2/VDmGT9MLJaTPAXaNCii1JQyQl91uL/FsbPx3jdIT/ig1hJIQ5EK/ov003wju7
Wams305YZEXcl7+/S7bAq/9+5Fb6m8tNbH6vvRceWAC7W1s2mZNczWE3zZVwsKcM
/EznpwtxB2mBB4lDLtQsGxlkZPFGRoVgwfr5HQg18VnKdh2Vz/UrIXSDwLzJh19C
aoPL5eWsWhCdf2JuCaoKULHHFetWSLqI+t7IiNDGfNkEY7h8sfBcPgUVfNEbbeso
5WTf66NazadBGUTRsHx1t0eHXrqAs/ZKUzNc60Vlmr6PCDEsUw2q3dMkQdpYVYEU
VU94rQQpiKSJGYha+BF7vqUGmifZJELgaSXAyr1Um8ANBfQ6i/m6CfH27wdDsJ7K
gYsbkJyQ2b/El81vN1JLZhR3hCckykGokfhmp468ssEpSwjl1dGGK/mqt//WBbXc
yBU9JE4BcyF0X6acuK1I/VFiQwh9dl7c7BsYeUV8Iv/yXwQDAx5v8MZpk086btrx
73f40GJMTYsUSeWRYJqAuutEBvDLFPNHwXiyeqG+1i0bDEM+EpvyWVapC3j2WOtx
gqbuvu0QqIjPjPr1bv6d7W28v49RwknAMZ2U4jAoWhVLde6pNbkoRcCbMvK+00sw
yCEs5P92TxMyK0PICStfCTEm2SD6JFEK2B97RewvlRGEgnR+NNPlnmo/Up6kJ2sz
U0q8XHhpIuzTNWPzJLLuiWfygmZwUiHlkGHNSjCrClIpZgEpQvAqioRfWCEYb6/t
PqzyOsePA6K/klfx0RbA6bg2lGYsblfdtSTsvLp8CPjPu3jsLS8SV+D8qMUyfigy
ag34DsQuffRB6rYv/vUe5Dv6R+PlTQJa7FeDTjsyLG7VsElFmThn5u5uEVWg/dAJ
PVVvWRNkZwA5BdUUTVYOIdxrWrKglkhZtQ5HhoeQ2CzxYYPXeyZDwrP8uDrd+MoU
7g0XCFUf5GQZyi3bHsjmz60/KBr/R9iWT5kKcJf9PTWOqtQ8YKmXZEeoILsjqzRg
wUN/7J/WoSPq2qj8dPy4f1jL4Ae3mw+RVhkNhzADmhKrVSZxp1MaeWq65nRYYxpV
ZqkDBoMslbsz+atp50GMcC1Imo9On7t103NcJ3fatGiqbfe3bY5drISyiKSVB+jK
8Frb3NkVMXEoJgn+ney2scXbvy4DJrySnyrmkLk8EyMF1pmusd8Dx0o6xhQjymVZ
RbqqfBu3/Uv/Fw+ndfPbjsv8YGt3EpUoQMQW6XkCVYeP7tWHnvfHuEltmU9AzBlb
5YHhyLkUVhrQ3jw16q8fJm5uFoilGkpJKd5I8RqhZim+EueXXIUSPYN0/c58BOD6
xZWssRstFH4rJvMgmp6XF1SgOBtyR+LFHtG7x48c7kJxXckRIUisyM04uBS3doMX
OI3Opk+pkVk/i/XEAHzUJ1gGOCehhcVOIR2KHp7mJ/SkzwaF2rg/uwcC+OcEQal6
+8qBAWc5qCTX+lCKF0J0O9vt8T+Xu+ENyWtJ8yGVtCqJwmbkjiK+bLZgcwGScMhl
3aGvs0EY31liBzDEFkqmN47tx+5/riDvXJsDfuCupcsoT24+TyE8yAJVQk0u13Ws
JNi2YudCuCzyu3VJPyf/eF63w5PHQUEZGJjZAZGPGgT3Yx3nztNGzk9LxaPngd9c
TnMir9LkBrDxWOZ2HIosQ8W3byQafTaNzW9x07dDEzr42v9H0ptnlN4H8QGa0Oa0
1dyCNuQ79az6aXVRq5bZtb5BLtSLReW7s6+qWgshHexOzCr/0Fwrb0t7xC0kdwIw
cKu0Kp+dSHqm8qMv6GmDJ/c6Y00YXGQWRQzFYidtg/rHvR26ygBSZIi/7FMUV0iW
SSzxt+c2dtVHaDn6xyQp4THYJBI7pJjbMSh4bC/MHuooE3opHEwzWhlpSgKBLYFk
+EgxzDVcvfqIdCaPiQHxya+TWC9eL5Xo+JjKw+jNKZ9a0clK7YPOdaSn6oiXO6Jf
3EOOaHqYCEWOb0bIx4Sz1CzkVMz6L6Q8DC1YwNCE3FSFkB0EjD5hOCZexh6mdra0
LhnuFWJIbVAHAt6rvMyCA3IFVUXapclzcYGnNFkl62JLFwJFpIxgVDL7C95fkt70
8G4Ax0pemumY566urGDUDFsRp04uI6jYBx/QXSah9yR7jmq8OCTNWiBUtcsznNTz
GZ8Ui6schnAgiKryblifOv5CUZ1uXs2jED/4+sQLu6yVubEwtY3tAOJKn2i2NhVB
HjrOkwZoRmMBep3T8EciDd2B8w/gP7uvovaSSIVhZFdTQ+fLR+YicFGEBVD9udvY
5sAWFQ5A3zY0SLHCruJq2R3HG3Gplm+rDntHK1ves1v4sEUeRTDvMdyAejPoy5R/
CQPx2cytzB1h0Qzf+VfkE5mWD4uhbBsfEpW5geAwmqSbFwygUoq6DpEQcqwPu2HD
UILEe3jlKtH0emVmVBL+SH/tBLDwlZzEYscMP0CSY+5+d76mLkBUSiPx6xnJ/Kyx
lUUO0y9iAzpOXT+qiKqm4eiz93d1RHmHHCfvT9DbMih6xV3SRjSpnH539QfHRcFZ
Kxo3+41wxlgRjTMoBcDuJVs2YEf5UovyZpOa5cNPDxD83kUV7mn1gmkYsp/ishUa
z/xh0OOCOzzOX0GFtxBafpLPOwEfKiOvlzqPz4HBhyP7I/c8mNXgR4Is/ns6UShB
8fJI9jflJxeUG9Y8StB1A7DF40IogWswzshRN+EIEBQcT/BAwZq32Rksoeu8XrKl
sc0J8m2+ryAT5XH94rKQHNW0vROnzZuubpwth9giUa2pwfg38giUg6kRAOiFIC0Z
oySbNSmzttN3G4NIgi/bU5Pp8t+hAcMBbLF53A7gYJ34LTIanZq76MG5KZ0zTgWa
nlulKbSfhyEythS5+Zs8+ttpcTXNsUMcsorZrkbmhrT7ioJuPWp8eIzQQA+UqxrF
DrUmq19OjK4DqjafOXk5v9xzw3KalBXzco0oLiu4GdVQQ+G/3j4lyjMKNR1WH+5g
z/EVpgj7KJAreqM8geHc+Gl4sUrqeJQ6o9mL55e7v+hrfSEu6spIhHmGTH1KmvEz
F99KV3uMLFzOVknWxXC59y0LMHLcGrWojNxoXN8ggSZNHsPYta9V/E6u5zRe/YAH
r4YgQ4++chfmeXFN79pcTj2/gNFWt4PitT+mucyLWopFlOtAXQbpvCrXxyspLiXI
sgWRK+WKuFj1v3jKCzdWUx/6Nqb9TJ1RW7zC56HEJtqq1h7PcBjiTNi9SHRgXVdm
ml+YF0GbinIOgsAQ+t3yl0aTK4NE3fGAxPZoFao7uaDg6C73MxfGTc768RdJjGsi
XqTyAG8F4AXLNQHSJAJCzcBYgVQpuFRNaSGpz0o1J1pk38Ls0sRSUVC+t+ai0EDL
uSFnqDiA4X0rI/GBXWqKXl+mg8RXz27wnhEF5gjjJOzolzm9q3fHWXgYAttoPYWs
8QM66eNpoHZK/cvi2XB1pRcv4FrdhKa4CLclhuHV1UTViR6TbnYuAYH11I19GmuJ
aqblNzxRStwJ9WTsHkAc+2Hr1+9ejiArxdHVwcnx0dz3xWgrbZDBqjtALVd3mpR8
iy5HefN1a4TMsbI5mM48l/Mlja4Sxnmf38hZX1VPHmluE9vHFYqtgfnXOqszenrC
omIQ1vmnvkDiigD5uzgNkDFAPzXsRt31soL+dFwfUw7aCBVe60V+ET32yWkQOPmF
AGBvRcUkzHz2JdW5YYZnnvfYX8FgVyu413H9IIJw87g/5GYARNWbL+b9Fez3vVdc
bxtT2b9J5aQ4tM6IlHCHudQzWEmyfVAuKpgRketdcGSKzNW+p7LIBGcnYa73JdMe
p+s1OlvjCxHL5kM6EZHgaS8cdR6N9KhEVfqul8wkchl6ohCwqUev9diZbnwKUJ8J
SFFn008KUat/6V3TY4wu0D7U0ilcO0xDxMWiTtdwGwZX17m/lnWKpDPjkmiF8dEE
NwzBLkFeKZvJFrhpq9n+5XQ/RIkx7s/qoA6Mas0Pp5MZE478xSCOLxoTKNctfxji
1D8OmkmUki1AZCPSR1JL9nTekxkYEyNh4z+rkmP7Y4/CNhyrV7/Ce+IbN3Te70ig
YAv6D+O7cIIKTZteUnOs6926zcRYRR9w44hs8u7CD/8d7VfU4iW+an+AEvTZbqBu
bXHUUthnwkBccgrFVdytwK3+fXegKbkDv1l8ougw//Z8HwHSLq1iFoOePKbGmWca
RtimkfME2l6uZg2LMUPBToPA3+OMSbnwod91/7Iz4wXN7iSxs53x3Nfx6+hD/QkE
UgiCCtCFaYvwbbkEJIC1/WHq3zLvDndL833IOr81usour1d3cs1AwAeWDBRtpN5P
HGMKz9dlL4XQ/k+wmM1KSlxi+mRrxP7tGqYthzhZJ3SCG6DCsNeGTq2LKPTrBYqQ
rHj5w3ghmNsYFP/PtcMVhLUW86tHx41/u93/Bv4W4NHmNf9Bh6dpLkLQ1F+4UHCk
mF6qF1LsyA2Y5DXazkqyhII/PTfUrFZx64nQCAEgkyPr0NiBRij/j0Qx6SWd5W6s
kO5x5Y/KVsPqBjh+pJHzEckZXXj6RrM81L58ZRG7YzRQbzJTrZZ0TfyArxdVR++M
hD4wxdOv31VhOm1m5+0fpeyybviS24XFQignMBY6hxCBC1sZREX8nETHVhsiCBEA
cIhb2rwEZT3eQ7If8+pnp++w8ROJk3CWIYwHcbg6Rdh3dZwhjXrX36LqEW2DGCT2
64GKo6O24mHMAhkLNAmH1F7uX891b/E79vZdNVgjy9rw/YfHqR6WZ2sHLuDVuiyn
H9/b5Ras6wkpQypurojVJOn8pekd5BgmPABmRVwhBEmXNcikYf8H08EeIW2WdHyV
fG/yK9/KYwOs3ck3P+OlL8JnlKJFc4aAWmjzu6ogEXcDqZbnPkAqXqssnYiUa7Wj
0jsWDwjux0GVtUgnjy8s5HsqVPhGegNwqptgHE1q2ULQ7Um/GXwvzKKUOB7ZOkzf
5JSizC6Tt8VWftc9kzm2r96cI3Ik5uiUik0jkEgNX3Ag0OAutjRh33PXQ/vnWm/W
ICl3iTRdrQrnfH4VS1mjNNfQ1RIEJDN//90mbnP6WXM4dYE6HXJmHHKWpJKS6R76
HonChZseQ9CwXViMB9E5b862fVAHswRPp5tOsRsJs+cgQCY2KD6JOIlCbSPd4VYu
4+Lp1Y9h+ze0WVzfqR2lkPjeMDDE6q/VpmDbsrWCSq5w/h7pkhV7IHp5P1B4duWA
KM8fT/MBwz49ZltJylrdcyVTMiqNpm1CXXtS9xBNWEelLCezoLKpTMSW3/pR+Zwq
IO3eSE84utPvO+y4WUmc+5BAoqqLYzZaBs1K4TQbpfKGFmqRgNpjO45qH49iMcR5
DWUfHnX3E/o1VsfdtBwm90m26gQCKs0cNVcjAB0zYnbwXrzwD0ed/QI67SJwc5Mh
Mid8csdJY851yZnryNJMTRwzIuv+lvSIABvoO+xaf/0/bwHosNR6+euHCYoQ3ksH
6+Rw/hdFJUcSIL3ZUncLD4ERv+baMjPdgF/3fg7Vis5KKZD0SZuMyw5abF6xgmfE
213gWX6wG5E4bHaDWhS/pQffhrG4SOS5/cSufXWe7D57Fc4aS7Q75p6qpxCgXoeP
Kqn28Mce5tTGdEi7f2sRsNOW2Txo7JGODTr+KnT3ns61Yew8ccsz6pKcEpilDg8O
YI9Bl3Azp8JjQcw8hDVoMyOypNWlz03eCZkGYMIrTJJw70i5aAwY9HY92wpm/SQn
REJWvJqB89Q3B65eoEIy9KUrZvySDhzkCP57zzh6GdMFjFeD/7oOXXLMlPB3rxGp
eq7U5fkFC3uaYUUeB7X+biY9qv/uK+/O72qYXFe3nbrI0nI/N+JbfLS7CGDDnUm2
WEeqiyHbZ9wdaegEekoMa3mdDeKm6qRzlT5qryJ1ImtAbxHtDTCD680A5CyOKooC
cw07etnxx7ijHYYwD6aFYzpH0agRVPf+XOtJi4hHzn14wkH55ledR/e1MU7w1H4A
Zkb7NqgXhj2XAPb51S4ACzpPqisov/Bb4AdI0ExsB071LIPbLMavDzYnDmV1AjdY
GW0tfk7pX2xPxjd/W5U0kCw41hDJ+RNo7ubG2mqYUaBTsf8fIWUtZ/kW908Y9zaq
X9kyU+TrV1A2WyazBPvigt8T9jbTJvKPivvwbQiYbqyL5q+NUDhvG2gQvS1wU/HE
JLYGBtLz1xvmQe70G1W/sIPRI6DTTS685yTukRf1q0tx8vDzQ4AOkHMxZ8JeoEaQ
VFgAgz2R7ciCUYYqmFqhsSA1bBE4rEMZ9rY2MDnH9LnJfzhctBcjNibbOZsC4qX9
A9S3UXtG7wewLyRpmaGZQizvlMj6FMwfkH3VTvedstuoyPWg/93MKgubcmoGJkXV
DdmBriZkU6GliONOuTSTK5twBGDLyM+cGFqUtJkmrFuiBws1rXk/VVNhNaKn8Z/m
exgQ45jpTU0JAIRPUtKKANW0kr1g+Q0qk7Ogc7Rg5Fs0J4MHMndRuSgq/NRsERVb
YNxKMx2kIeDyJ/4gvOTCywwWBMOvwxyvR80PJEY+OX9NtuKcbGtphNTqctCNGuLE
ykliQGQQe4++jtYevIAfK96MJCHCEutjKanP1JjfPQvAZQk/LhHkjgCoGCSS0Uj0
HagRKI/iXaPtsDmOF9fZ/ZWSuRMlWlfcakSASh0e3+ccTOWJzSNgpue3p1dg/CAj
cT1SrTJ36AFzCNcpb9efhQs5Xk2pkgIyFEGk9sbG/n+iR4yh8JhakEe+FvRGKIPV
aGbwf06vuVQ78WaaIvfUSrwr6gXWEUt+d1FzOKvnkwbAmuLdEnaXbhWkTqZCNS6j
pxJuc2wmlhXJFXnczreDe1eM3KXNcvSYPWOWmtKEwwwCmINMa/FqzpTL+EwL8gZL
z6HPLz86Kk3wqylbWww39Sy6wg1zNeE7Nh+eNpTDMzaUOMADjnlkCdcIk60FNf+X
6LRg3mE4FHZ6vFOpa317alZZomWFh4vBbqE3DlfHmbSPe/8swG/KcFnkW5hfpMb0
dCRqlCJ4P7JuYjliKojIY3wnykTorK31uysKI8ANoQD0zWycl7/s30Ho25b0fq5e
y6uFpSMq1V7eWsmC4VZluGoyY6QQPwSmHg9hTBWSNiNkdK2UzaQP0623IRd2O+Hu
lMuZqOIH9geWVe9yJjnM9mggrx3WPNqeZLfR1ZzcUnWIddBS1hWcB5oy5zUF2yLc
lhL/8tQjM6B85TPLo04Q9lBk8YAHKXbMb9rKCj336ET4ZmwupUFlkv0+DZwdBuQB
3klXF1E1vdlukaAHSl7cvHszzK3a8vrMcgqaJF4j8AApZO3AsXLjfYcc6uz1l5sL
o5H9g3ir6suVBHAW3BvNDezY4Z7Eqf3sByo01ZjLcWQ6DtasYh369cFesEJyh36O
myvxy5j/Za/QSSPYfh6TZq6O0KyU6Sue2X5OJb6KSBdn8+Gq/HpzOFsNqXCfI8yy
zSOxm3D/HiEZqUuCK1gn1nFyD52DuMM0lvBhz8eBcrBz99KIbriUXuhbXS9ET+bl
95RwbFZDT5ngNEr7DXelHsiwnVX+KxCWA72MPVXbvHjaEGOfkTu1al75fgjU5n1K
uS2qlTwpzTIgcsXySbWep9rP93K/pySh9v6LogOR6r1nanSFE5HM3c772Eg7rlbM
/bqZO/dK3oRrBVg7EPQ6hF4L1gjcUVOJKT6OLF0SW5TE2bLfBhypqRcFB+h53gAk
LQ7AK1TJ86Uzl191igi332ham7vPagHbo40q1JWJ24LuVx09fV+XkC8OAZ5eEeBI
it6221jk3MECKbbX+lIhyrYMRXL9HG+ShDZ6LuG8VdVMyR9nawVC1iZM4A+7f0Lk
aFny4lB2e1D1PJfjnUlyMGYcOkjLnAcSZqQz1CsyIi7PI6RHHnPw6Zb+R2R5r6GC
RSsx3lNPGzDAAXd+y3rlL2z18oNwhYaUxkMdRMdt+Yk6E/ayEJlRssnzw/Z/SeeG
rqXd0MWE/tnZ3fM6AULzYckl+OfiDRoh7xRQO4XxRbMxF+qgldwVIOMw5sugkqZZ
d6b7dC7evO7wpu6LFuKDrx6aNhAEy0wd+it0iGkAFz1LPZTa8TVQMX1cTi03/a6h
6hJH/EvgFbnIt3Pht4ht0067986KrSFQvgh6erfH4yc8m1CeE2P4zAx/R0Xv0RkY
Mh/NI91FNMyzOpRHXGbEhMZWviOyzJ2M1naxulIWT4ZmUdeiRFErs4xbRqldAxPg
fKCXeBnTDLF1jt/81tRm/TbkxSSmY63IiV6I1IWfQJIWRRn7xwsoRJCvF04lijLq
4tBHfl35+Mfts/sw2OfmjD1KgwCQKvhHCsHJaMda/RqH9G+kk6/n/9grnY5joWan
G6XNSgfVVVC7GbJfIuE5Q1U+5zNHA4Y1se8pN8hIkCNEtfVORwhvrTc3+kadvE7M
LCoOOE1TWDbUP7VZviVaH8IQqry8JYFCbD+hpASqXwyD2sDRPNA1GhBCe3BN/lt7
RP039tSoudaRpjHJlrdplujfL3HjKxKi9G6rsGcVWah9U1yW18GM+Ja3OOkVBDar
WKMcX5qn40dXWpHnz+d6C2KXyIg4Ow+VxnlqPeGrns/Nz0+/BgQVZCfigGa20SbV
y+vs1DxwqDJnZm/v9P0alHXPyr8qDMIxZXPxsdZzgq1EAYPCkXvaaP93R1B5hnc8
eANJbz0hVAsvCyB1cyz2FrdgA+LKK95IZrDxPZmP9J8wA1kFIpmG0tLJNZTf4cdM
6oR0gvJfiZK904e0Kh4p7J4KDll3AuDUi8yXTJrBiv3KdkGYiZpbPesI5qHUdf33
FGNN1XlqOmllkVLUM877aWIO6lFzhY0h6gFoJ/+8N4H7WW/LSmXPcQmia2em6XIU
ZYXa6Mz0QnVGEvoI+6bgckX0OrMv3VjAx+2xx9ymHwdneubKQgCJ96mtD/S+TyKj
3juEHddiA/qD8IiD73xaxP0TG9int91Q/lXkd7JRMWWrk8hzXpSuzpA7Hbb/1PGz
q0taPWs9+tkahoJpjMxSowknGqPduWWMW2OiF3LQKRm0dK3OyhGE4jydKMcuAibx
t8jWjuqHioTqDxEY3XIYK8mF+KRWw9EWKtgq+8gTClwnBh6ksndWHSbCvQnt8RrC
lZruKA2xgvoDicWsGZ/sMWfFSMaGkaurK7uQgvyBnSyLi405LLfZ/v01wA29qjW3
8BNd/IcfTxLV7HfhzQL37zUnMR44Z3E4Qlkf/EjlaQa1MnH6lTbZvdT0uCCoI69U
xuq4r7YoqPxRVQU6Sgimge6L+yBz3q4CYbyUBrRmyQXhmSsEQmrYAtmACkivg510
xhOBlK2+8C98Zo3ASfkH4nx2DRbn5RzpuHAU16S0E7+CA04Q3tFRy66KTP41q0bp
IVOLVIw1dJ0ghSx4Jog3wi8bKR7orYJdM+TSgBaGI5qY1GE0YNBd+AGaTJGq2YLg
SAjbB7kGS1uJnP6lhGp2IfM76mVUYKeiav/9lL3edm4beXO/YHrdjC+wzr/qRokD
v2DDIMqW93Sd/wYS6Ej4w+Js+eXmXGFLTYVbCCwP+5oTFwzxxgRo2BmPAL+lbdo9
wMn0esUd0dF+cG5Xx+kigayBNgHDR7jL7TOiwsSnsyuuYTr9IYEbjLgTBpeBVMRi
jnf4nuhrqhTfiLinoHpHoksUwOyI3IDAYxKbkq6sunjZwrq7pDcw3k+qvK/VjEx+
l7XYRRlkpNHcznQOP/60x/RdBRFfbcvGxVspnI+3thEQVwHMlc3Wec0fJ10DHWMf
oumo2WoXf6HcNSEtBdVajVZhjBQ40bO8SYEfa/bB7CAVMp45jhvYL8qQZEyoSgfA
8v5MOmTi4VcasPn72vlPFJ3s3Ik5WbQS95hpJbN0QQtB64NYnVPrRuULfeWULXhL
9pFioq7KFvL/KSpRm+onhhI7lJjvzk5rJySoETIw4aPMnigKDdRoM4Zww/qu5Kmx
XA6gzoi5j0okW4ODC4ihLWwb8weGWrr/fU8PSxzVfWZY7s5AgRsavN9zkGtBhE0o
Vrku80OponDJjCRZ0NlDXKZzXAkItuemIb2l5xiglXNQzJ7k+JsUNkXPpyAN9DcO
AsnMPgBDowluRzHugbzPK6snla4agAm4pO/e8xqY+Od60dTdDTGaDqd7S52ip73s
oYsI20IE8R4j15TCjA2anGnXmvnCJa+adRjWDmRTB0tTpfbCAzxdOmn21UltogCh
kXIu17NuEMfuwKxsPny4dd47AGNVoqAJdTQ2nJ6P5GLdlb2Yg0Q8HCNi8QmNSIN3
U7/JNgHb6XxR89zxNU0gTKDTbGznNK353E+/PvxpZ1Ej8DvwDHlY3AeuUn6zK0m7
RlMYabuFpYaA5HBSqmmjWNll7XwSiiUJ/vsFNor1MfJIGV8OVD1ZYfnCE+u3KvHp
2A/3hBydceRYuWAQyR4C5VS69T4/2rNLlSC+f15l8dAoYdDAOL8LYgeew20s5A8A
eBJKP2Kl8zEVFJHgr6flA2ey+3j5em6t9vjCTUQ4IaCErOj3oyFB0qNt+fvMW8fU
jtQuY+5jSKknaiwe1K+PaiRM386BT89gmW+3eQUYFc8O0T+FYWJWx90s+QQ/H92n
wdM/9UPqVGZpdYD2BlE6Uji9eAWhZwcKiceVN4We9NnUOBsuk1ATI1/Y57uoaV9r
HvMEGs6SwzOu7UBGpzfxvbvCdY4Nihdei9zcZRfbKbHBMsyO5Jb7Tv0ZmxpK34IK
zQq2KTVDD+mvoLiCJVwQ/58HeGlTwD2TyD9TtNXXG1v+uS65NVUhJDc3o8hpDgLf
DLh5Qn0j/8tkf2XBstzIFkT0lw5SciiHY8Uw2DVrYZW4bb612ThVOnGgGxuqhHyt
ZVF2dcpNJ2H5MF1Syt7dCSV4zhr0wXpuEAJV4CK8QvVvLuS5WG2pbfGZafRVDGMX
Sth2vAW5HuGerRolt1jHo/2a1es9Sz3jsTHLKwv17mRG/i7Cw67D4cLWUKt95rDE
xN3JkH7s0ndxBaqc2fZsFU+JTIuasbYlFHY3PQDzKOmRPmJcIgstSBYxx4ZF9HmB
7XRy039ZwrWjipCne7SvG0XHLIsJ9cGg9+B8CfUo1jsokYeQpzr+S2Em4ta1jee5
bj+fQP7m9CUvS6mSPtYWBBACX2zBtb6pngn8PL0Rm2f3xv+8EHzOqqUZZ7PdUdUN
m916fXftHofdTgK8ZcIr3LklRDb7LCYdpOc8JV+W5c7AqnkEzQkd6UYwz2vEkSCg
1HF2+aXmY+kMJsY6VlgG4+PaRBGoX+BK7IEVWVAYmE9N78vyWwpKxDClDQBIfC/W
zvAh3pV3KbXG6ZIRttzjSnqTPFetlk2t4k86UNTFq+vTZcfT4FEmDKJo7Vh9ECVE
/AnZ6uXwgpY7ZfJQuwHqS8EXvnZopu0qwTt578FsSoCky2Ivg8Kgsn7hWjYBAh1z
T1CghA0E/u6QtuwCw3sJSq6IsGBaAbbdR3QJ9lMO7Eb9T3alYPBlpISYjJs8XAvt
nHuCSpbOZOb0vIZG8wQnAWlktZDdOq7oFCoOHiaoTeJpWBmydeRH7FqPDZTiQC5o
dAoD2iUBHlv57/HPvjfOtvsHcEKCbOVzDecs5oYc4W7wULvDvzlgwXtUq2luuQoe
AqJGXGiiH5Q6/O4OEYqUewAaUUYc81DdVZ1MiUcNfMnhleun+uQVPgoKWX28EbB8
CvCKjoSMvkh/bSYKApr986SCwfXAzHeAkf0gOBmfibf1gWsYL09PBpeuNJvBN6Gw
TDczyu7eH9u411vQ0UKhmTJl8v7zILheTxxcE5XoIyIPn7QliiJA6alaJfXV/Zl2
mKIFACEkE6rsQcOGg9rpNPVHterkdm4JqAfN/2cEDBq/edp2Yh3vRRtv4NhJryRt
cGlKW7c0MG8SOZceCPrMtLbAw/lt92MluGB74+lP89k43b8Y0aabmy4WEWygFRcy
HKaruPBljHIjSRxsqlnSQM7tLoEHYFS6Pm38JvLvaZ3mmsxC5cV6bz5ffjj434GA
k9PWzucOmp+gWQaEd/Nf1Ak4wUCYn0poJ+7uns5ktUYEf86ye3Kxg10KESz38gru
ky3NYcE8IT4cghLPMTpc7wwwWDhDXNiynO5gc+2YRXBnMPyLlSHyh4ciC0HwbcXN
F+829YQstG+hv+DLcpbDaz63JMg5hSTXcA4/Kx+4itM/kihPA83wVsVf3sx0AXYn
JyYOW65Al+wrvudxtX6AfYDx1qZOY7d0StY7czlcBQI74m5QnBvZiqIKZKDpbDwE
ROAi5rG3lV4inQnwVQ+3RzihMDLw7u+b8ibhXcF9U0k/e0KycnJrRuLFlEQ2EN9A
Fkhd+RIBCZMLPRbxuz2VowvZfh3IS0xIWwqdMUx82rtGo+w7ZsJXcA3M9t3kOs8r
PPOT76S9dsZTmE/cTp96TxwzM69JwzWxoTsdrWIE1HeJ0/RuJfarp1ZZ7sE1bsdL
pPKd5wKsiPhVKQ7gRHdf1LDeEGuANhnUGPwBvuohLO34oG/mbpz8PwRz92J2GwZL
NZnh3KCILaSzIes++kOKOGIOGXZO6vq+yExTLIJ6p835VMppm00fp5THJOIsLm1v
wp2/sFOzlWegroymoIQPf9zz8NWKm2l7iB3NFLNGqNqegf7da70ngK8N1z9twuJ/
VsQbclTT79Cp18kC/FZcNsV29HhkXRXJ5iKbpK5B/1qVmwZDZvduiwHJwPk0DUlu
H5Bh+vWgCL0O5eZgv8lvZbahc49bi0O6XeCmRyf0AigDFg0eurJk0ZguJ3wkkF/5
M0ADWubO+gJE8o8h+GA3GD15qNXBl390MaQQbsx/ReMqzfzrDV/roadJu5hcLesH
JDBupKmp4sMnUf0uStrX7ZwyJA3d1Y7kREAp9RO48Nj0dLBewvA7h/LwJNhCG+aN
EdcY+6ZcRIMudR0IgO69YBB8+hu4g6DqdLdcEen3E5GD3G/FKgXhOOo+BvvZHZUs
3X+T33ByDPjTnJdq5/jJHOXL2Les2aabEwOPUOVl2ELDuWjzYikgzo8gzaVl0Ied
gSaz/+tVraHR+jpMFrSdaiGEulYMBmTkM0g1pnxopbHQTkjU79EAUYO3qm7o1ymh
4/JOliZh48YJLqFOpFjiR9dXlSLWLs1LTXL/H921OZm0WMQaszLQiDdIU93YBFVx
LBlCBCn80T5ilqgfswp5G7MAT8f5AsTFKonH/pO/WcHKIqFAHm+Yj3adsWXv4Xq2
z+uiPvvK5G6lPRyLPtFoutmFXcs6fI/fooO1g1k9GiT7TpuFBCmPHlLrlECF5ikj
7/GGgUouFEgfPCp+iPZeL/YxBhRiqlpk2yYXyFMKoHdRd91iH2B2DLCW4ykhLBQn
FtC4TcSWq/ZZwsrnmS7ArTSYLllZwG4bjXjEMTdV767JhBHqLSV0qrFzFnUdVQvc
7JzGExmGkDqIIvRRBdow3a+qbOgwdMQTv5a5UXF1nwGH6lgc3rG/qTBFFGMKxg1f
r7v2MLtVhQDF/LXBkOkwyD2P0s/0VQyBFX3eT6iNoaSkDBfT3i4RcoZNWE+GxlTt
ciyejuA+/NSeR9tYysdV+W/wxo8dzh3Gsf7qV1ss8aCW+OvcOUhKMHwyFepOiodM
KzdldnlFEbMs1UXbiX7lXmNwLEocEi6lZ0RCvBmuJC1ugNpNZqTdHAengUP+nVDB
JskLwP5R6r9EW3dZY+FqG7+II4qTIHdAPEgQFytxIGmCOY3YxeLhJvRxTWVabrN/
Xs6ND8/zf8N5wl0qqxhQ81X6qBmlsMMAr2iAIYR/G3SID2rk2pWGDSBHVAoIK/3a
OER7l+Qg2iM1AF2g7mo1F5m2YT0dKheKrYHnLaZ5HKDInBToV6Zpl3+7KxtEFqpg
ofJWVMOHFXLVKcaknnnCHxWIaoPIhfn7kE83N42UAsxU9Ac9qxnmRWsGjqZO3Q0y
hxcmiLpCLYdVlw/jEwW8NpOvosODjbCt1v3GwjyAEHM5PtL3LEoD7trNkxR06VFA
fkip+aG/nJbye4qgmTgoFLdilgyAmGCu5vm5UxJ/av42jt4Mq7fM/LDYt6s0SeLm
1CRwUu95hhleRGpW3jLsxH8ozdCQjvmGTflqJBffYS8jHUIW+N6FNBJDoe7C6Io1
ZJhyu8rjIf2m8yDBR4VzzSbLAiOtch9rlp2swc89i9M/jwbSSzn4Eglrdvqqb2N6
pxW3JwY1B3wcrjoa1sOnrNk+KbMmUPR0cHOg+f1zzE5SBION7EKJZ5eKh6sK8KLh
LJyB/ay/vBY/mzlR69oHd4PjgCZyzOKQf8ef6aHfx2NNJOpizcbW1IS8Y5/wsv/E
qAyP30eX6u0roQspd6aX4+nXPRbuuJ9FEum9oO/vSNCcSY1Astv2NuLrsVk7AR5h
jQiQdYHCsCfAQN+veD5Br/Xes52vrwysAWxcpRDBk3+nW27TL51AuZUSRW6ZDIvH
iagq1+ptd2W2bMse06F5+gS0RypEzO5qUAm0M8V7mi3CC0jeqWkNpV2FbOdxOtyd
d7XYbqwyzwyuMmAVieRZeM44nrY0dHh6bOZEPzkXJh8TUomblBDGj9n7dsyGYTha
jw83B/v0mlzVrGKOj9S2I1cox9ZKeHzkQpcKqqIud0zdYOaOOWhJ8HzWLlzU3AwA
YYTi6G2wE0DyzcB9A0MpRfc60izBAmAWjzUjp/n2uKLWzMEmGL+X2nWIkwH+LJTQ
D0ru/lbKpFSAsWIfZQZkqzbCEPrRLpFLqogn6MgsDqX7HPu5xUMH/Bi8cbEawNlv
sf3cLcqUl0ElYqsEhUEALhifZ/ezwiR2A3B0lvS1v2P2q6ehnhNDl977CO1UgIeb
wRFCkyyduwQ4p6wlW5MtVCdFS0nuOpYVytvFMJQWx4TiaNwusFAcqISnAPMjIrjb
XYj+DEGnXXzdTXjDWw7t7hZOnqAH7DFPqV3CP0gvDethOh2ID02sTv3cDluHnCtB
pGyDWUaYfLBHccAukOqEeQ/SkCDZw/hFKZU6spOVQwO18YEFiy0noANE4zsPqmbZ
WToED0JAEqNS7lzfxSrs9Fe8cuya28mFv4K1xEFoXyRWXKNfom7DK83AnOX0DxS7
pdc2oWiLDITeuYVX1xqUplC0A2XdteV2ESsrDOcHjwT0zFZ25HcOtdNe3r24quq5
hYC8rCnBkm+KtS6SF1NDSG7s3iQN+7G5XFjZldS4efv2rPAeQ/zgS4A5C2uMnZ7m
GMsjLo46cG4NgHCqdiYom2lCmrWzw6fjXSPQbQeTetHWqbzrMeudcJkL4d1/5TTq
vDRTrcdbD9XY0ZiqEQh5JnJ+NvPBZjfMGAsZtL66OzExAPhygJg6ccFGKMxK/LCE
6ZOjUZxJQG6Wu6YmZviiF8wRirCgeLPcUSy5g6A+i/mS9MfjPQ0zv04O59VKnMDH
JyIZBxqrLIfIcfqKk8MJJcFLWuyp3xXmBBYgE7NGWftA+ck/z756VoWeJI/l5cCW
OWoYyAgT+XaiFkJtQrB0lKgDk3+aeHYyYwBTz2jKcElmOgHsAkRWbvIgYImTyHWb
DIcS+f6gV6jaIFKcnyEZbQFBrznhvWOt6NkAwpu07llTFppNx2LJuixpXPiaSkqM
7y1OD002KvILQiIDAfRH23izxzZlUviqg1OQtvKUxgXboj/nJIHCBpu/si8cKCqr
H0C293Ez19+GzU3cv7lenrRwZh72OKtKNXHtZ5/2kYvj5DI6t81Bdj7jKuVv7oIm
3/C4G6bSgWYuCjy3VkT4XremOGmuh4/k1R5jdYxg+GSZDSpMpbvADVlWT5wHcz4d
H6iEuxI8GFmZXXVv/zQX7G0mUQkxf6M4dAiPOCNaJF2Xdxo9iAg6ZHGhvb8cO45B
7V4ScziTb4D85VaCKmwb9xOc+3MGqIWaekgerzh0eOLSBjpZyM6WAFzJYBDkNEUY
t1LL8RD7+AMTafftkMZbDNr9uoydIyP7eKcs2ULUgKX18u6Y8uvDGp0IH4BOerHu
onyshr9hyUu8w0q7dt5et4zDfMuRXT1/ou/iWE984wF+KkhSCHHBm1U/m2KvADXt
ICIhC11N3jyNuf+efbFGVBgv0gOmp4yxezDlmPnoTtB+ARNKN5GdDyzHHoUpVja2
vVkGkfMiZOxgfrUt7wacQ2r/hkXdyQvbz3TT0hO8/WNkJdmHW37f752U9AsgxUyk
pzWIEqONglMGUpMiYQw3VKxdvqFdkbYktfSpG1POqLjOUvOBQMXuenyhCiJs+u8+
ab8MiCuCqreGjZ9mMxcHV1R3lLyR0/tpRRRGfAt6OuysmqAIuNIdUhes5Gj/yx4p
lPYZIiiI+4rEyWjDRl4AVwb4ZlOnwCydESVp7C9eZzLpeUd5nVpEcB3dJoht3fxZ
8Lce2A/5OjywGqKk2Uv/qmGRNaFoBGDHpEJ0LhVrAGrVec05uack9vd/z6JblhT2
em18sWrmUZSRaJDu8exTurOHzyE9tefeK8yfmPNaXEo/vmtO0TFOQk5HsXVjWg2T
JGWr+uD9YRuuA7by70qEbq87kWhKvkxnz499v71x3fO2l82x+m+dBlcg5uEFkHvi
I1v642mwxH1iaOo+FQr6CyfJFATSOilEyfYNB1lcuz07p/y7jVpLO5vaIaHBxBjo
Zdu509P+hjYojMSISubuuaGqdZvi1kiJw37F/OzEfvZdy2DZyvhj9IXyzK7od8w8
RRfrvfhQxUHwwNDzx+W2B/+2Ihd7GqtKu64WMcC3rGdsbtD4CUiTeIggW2RAaybA
8f6EmhAKgw1aXTrW+1OEI3hE5dbTwASVPkK/heaYLJgG//LusYlJUlSDKM9ridpz
k+oscAZTPdXO1uRNzWK+y57MPz1YXGXB6rK0B1xT9ZgL0yjkJinf4T+43KoIwbgG
RFpks+FIwdyI5OB3DaQOLn1pYPVFRd1EujXbP6PYvxBwTlc6eDePRjLymRcr/xul
AF6j3udclvLevUF9O37ZD+nzY0z9i96r/CIBQeD9Mu76FgRwSaOi1I2g56q49alY
RSGWSQlh4RZjMalUUVyGyPbdkUxtzZicrjfu6siLho/i9JZlqa4iKi6c5YknTYj2
vd/Qj1Icjv6eVvYDB1ZI1laxg8sZkLSH8VYrEiQDbaBCjqk7mgPg8NdjhAEAddh3
qaPlPrB2kide775JhSyTc58OsPIt40MO4L5OP4nFVQ0YFlmwONdQM/C981UyoaE8
l8ClV4yFSoqI305iWB4lV5Z2UYnKkWrX6vjIfePB82yKX8PSZkqkilIbxPLJVPy6
/JfbCDcrlRqzrFrP+5iteAaFsTCtGgqkkEq/DHFTmtmFMBiXvyFeVkNxN7woDkA3
FIqrNhV69Zaa1kvvZFtVzV/Z9/E9wOG9pwAELNPJtlVYkl0Eu7Q6ek9g1ChxU/D2
qCM1Zq+zyXexNmwaciCKbT5ax0ujGaGFgE40zotQb3K8RIaNe3QVXEN7Dus43Ix1
Xtv3sW8U6MHFuGjAe5GJfi1Qvgpu3y8Z/pXz/iODkfwCvmGZZQQhr3bit0gWpbUe
NxZC5Hfw/uMZEpSU5naFi6GEUlCzTO9l6uBHjTai+kU519M33hQA9Lcjg5b42zPq
m/etBJzvHMZ8hatdD1/OfkW8Xse5HQh/oWe/2BNX5Fo137XL7arz7CSBwOkClxZx
Adl5b7mqYfJnEIgVUKs84l8JmHoy/5VI6XZQjemP0j6ilK5VjgNTcXYYoXk3/eqt
LIwHuXf2/7IqBGuoi7eXzxIb5sIsH8emXNF1Ga6Ydulgf6SOLW/wl//zoxsqr7FE
xqhUng/4Xj+1S+Xv7k+jaaOauiRKurKlpnvrBKqr9IODsXQEqRsXJDS4EjE1y+z/
9PpHNtxFWsPEfBypxABOJ9nkg99XflL70YCWdcmOapTniKAswbT9HHMuYgGlkYp8
UjoEqzMwNLs2SEr+o82u6zDBAfFq8p23wpP0Lp8JAuMWZI6LpXnCThjC9ASpZGQY
Z+4WOO6C28p3FXD4Zxez/nkHbObr6uD55DYvi3DzVcded/uEeRtFokkUXZF5tK34
`protect end_protected