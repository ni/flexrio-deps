`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13312 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
JfUWfeA+KKoJK56uw0JKy0brr2yAtaxHJVPp1e/rl5bH2uF556hiEAfsCGWxVlj/
+xMPMkmI+k3araIRc3rGy4TLUMWxaGukYnXfgyiQAFHcWhG/cBlXog0woxtFuqV4
OTZjcmJfA1KDchIm1Etx/XsDU6Qob7cXuHEml3buVgoWIQUtpgGZCmu8gTnkVOTu
I0K37xOJpIdy6gulpMqN/NHyudLAv3IgrXh/AZmDfZMEPlOftCz1k+V3Fsixsc9M
BSjh9/j1yAlLtIk+UKD54eSIrwbuS2nSEVKHcebX4X/nBL9THpLId3IbJZLxCBST
XGUxr7F3mIgS20PrervNIlcFsxmXa9+pWsv4i4p3s+1J0s8YEtRCgSHRHuOT+fbx
ILTFmdWxgSaPsS42OXChTVkgK1JSj2PIkbAs66wr4chaBuTGf+w6ELM0nd9abB8v
ptKXbTWq/u/ntbIOSb9ad4z/ggajquzQNvfo8WRA6AJ+XA176oda8BpGVjCllu5n
zVkh/sVQmJ/gdKNcE78SiZ0HAANwRTT21jx9eDbJY1HcX5rMAvMoyWvne8+RE/aD
ULViq6Zb3oTcuiyjbUUCOlPWNYydRCjU3Ce1ZWpelln7fcgOorZCxsWE+IXWHLHV
ieh1xEVUSIG/uUVo6n+XiiND+GSF4OmOcZ30q1yfS+iXb0PZX3WJpB+1NtI6D0iO
VubhZmhzPSameXinLE5KltspHvX1qrplOhcrPXDbXylgPLnFy/AaWJ8gktuD33Zb
yuuO7JdQCjtWjSS/aBqQErXI+ms6rlXXVPlpxPPKkL19kTtfkwp62Gnsmp/gcQxc
8lgYbUTXy55nKFkG093SpFcSt7fyI6luFSI9R1QKvZzgVCVEltlBuaFs0XS1Ur/t
uAWlTZPa2RnRVvvnmjM0yf0WjfUI3pUxaMx0KNJsgZHN6Gzxp1gANcat76ktjO4Q
iAjUXbIG3a+sPYOC4YZlPlsP66dyuvuA4Ruuh8mOm05bvuhAnHYJGCJJVlj/1z2z
kBGWCmHO6kgVTRfVHhRr2pZIcNlUL0xXgP4W2yW+5eKWvseiMq/QjHnSvDz1vkPI
uWepfCnHiTkl6MqvcYObKcl8R3Hyr1A5jn0HiWpKkhzJNFaUoKgBus3IGVz1xt8v
+qvQV8fOsDt+N5wm3u8/Koe6GzegSpiYABvOKskhCpb3QRMEwJArTriSKt5aQ7kI
Mh+xFsYM/nrhuVZlrkLkEaSdFj3adFnix5L87WbJYEZzbz9Swe20+FdO8zvd1DLf
gDjcNgtkL6Zz+bEOJ79LhsfIVFkZuQ8+1IAJi7k3QZde0P/fNGee14oyTwtfvTeN
/DG9fT2xz9UyxDotCZEtVhvw+t6qLc1eJIbhQV18OfX/eOtvc5xhpgCO7nKihnlB
J4tx3gKiFzQoT7511moVacYKrKP9culBfXiwZEZttt399STrk9+oBcYPsR/19x4a
ZTT0HaDE9turHTHO+qjofL9pQ9Efs0h77a1j0P740iXorDBderrjKmku9Ifubf10
i57LooeGEt3OUFClgMcZpgddLL7jtPx/7oH1bAO4CJZ0xIdZtsNSbZFE0XpIBLQE
GOfF793p+Gmkhzw5x/bvEgSrcAu1Ug+FW3WHlB/t0zn9iLxtL3Y8Rv5G590Ujo4F
gA/Fl+zpb+NE4BKsAOsT0xkqZJ5HJjIQR5RW1CqpVYDic23HQYl4qxj/Zkzaw2KL
ATPmyuTQlwbjkj+nxR8pLkhtBkhMExfNqc65fCb355A5cAJEWMKn+JDfUKmHNh8T
COKz/50RDZZDImIJ7lt9ocueJAuDmbFzV87gglF6knzDIc2cuDG3Knienxt45CtG
/dtE2Scrgd3mso7w54v74AF7pwzQAqk2Rwt8K2rbhPZPVhipvTr4E845UuBviigJ
gjZP5hdY7mAg3wWBLCTbk2/xxD6tFZfGiDho4vbgEyUYdd0dOClZChYS99kjAxva
ZBLoVz4vH00+3pLUlpiNP5NGFv9Go76/VqhUozRNt5HIEkfadr5EuEP218yiwHge
B3e49cz8EObvuP8ViDlh1Mjs+ms9sNVy4//t4IIDboSZ346UXsJDyKWQJAZThdOM
6dA3bXr3j58Gbo7bWbH0HEZ3uIEyeJUIWEYl/JVfy36PoVw7sdXreBVR+Viz9YFa
OidPiegwBIma2JfrZOexM2Pu4OOSgw4cia777VwN0T7GXMavTeXCGpb+0ft0MMxA
qnNahQqxeMp4UtcUfr8oXZon5BBBlFo3yPMSFVZtchpL0fD4T25NqUeDOVAN9hm4
VA4JHq3D2Q85vMzwmW/OeOo1fXGyHhZYcCoCQydpZ+YXf9Y4EYy3nb7N7xdbFXOO
DO4VsjAYQ+FiKHmIymyERjvz1Yl0RgxjiJF72+aYqwpXJbeM4yhQQQAGvBTn3mGN
hdqJ09cw3WXrUAO22UERGBfiwH6eRDVSzZHbqanlxnXlRUXOKhKgacviSvPvlNfu
RaWokYSscDlNhV3lgy3FSbFedVwwXfskt6xoRfbZyVQvmAyc0guCdabMk8ZNlb6v
kz/NIvf86KwL/PTRRlpqBYEdG2Vo7qzh4cQu0N9jqnE3RCMonQj9VxcO1i/mG8bW
u4jdaJazj8Ln4Tz2rfqndFmPbhWvsxjc5ERJTkzAIzTf1lqr4K88qysYBNwruCxQ
e28T19NP0njAScn4MrYN+ZHMyEh6hywmchTwUyseBvS/kD9HC21DYzB+9bAVOIVO
Ej7UdTD2CSkDsk0GELV+ZH0mNb6JeCogjoO9bMlB84v9kog8DRlEe/vCoPVtUqRh
0zjc9ym35MUu3J1rvyDS+aLmtTlegTNJA1luqYHEOj/3EIwUVM67dMid9Miaa++e
TQtb4MbLE7qfp/HMvDnTTghP4WGe6zeJlKdVJ1FzFu7/oo7rnj3gQVMJBph1mg2n
CstgVh8SzT9ixVE9uzQsGyRDH8EJe2q8pq8ch25tedl2bS1xOm/X78bbt42dT96K
tZis9KHF1lr4oCcslL/orUDt7rM2sciMlaYOvbdnenGtgRMEG3en5S7OY7Gk1GVG
cUE9w+xyPjKuBk0ejkwLsDGkwz2SVD8wfpnO1d+lDCcfki+kJiJ68/6abllgX6xe
f3p4UlZX8uW3IBM5Fp6MOmFaBHaxKmexxSDCpYMR2ktKCPF6Jv69PsgKTQ1Ek8Pl
xzw+5EyyaSvUCmxnuplTYbc2pR8eVBgGw/p7x3YviemlSzoNZKXNB35drzPB6Vy4
V39yWZhRXPLNjs0aQUOTDdLQH8ZI7eFsHLu+MNsro2Y03Xvn21cj1n1+87REaX/U
Z82A+FjSF8VyHoqlGHEMJOy3AynSYlaxv3dD2zLJDxwVILlyFRoH0X0LDemtm6Oi
42xk4p/fIQ1Fde5h6tm/n6ZeRFIEgcdNUz9nzjMg3Fgs6ps2g9jPjidooIp0ai0n
LpIuDF9bWQQJ2dnOGVqp0eIy97qNijqnsSC66C6DUQnB7le5oBu819qg2X1EVsIU
mpScaV8/cQYDYgeo/zmmUns9wIFAAw/sKwZjLRJ6zzgoXX8NBK4n0Oae59jOtaMT
EItbKUh7gEZYQu4eiKlHfpG0gU2cKq8ki+fw0HtEeJkGlCpkMx81FGF5BaT7KW7X
n/ZbIoY8CuguTO2u2Bp4uaHQvjw+rKU7CgHtA+ak00Q5u9yKuqtoNhV4+ekD1ykY
i6Gs8Y6G73cTz6WrdhQFs01WkuhBEgL8zUGEsp9qTdvT2ZBb2bBVuU2ykMHVCORN
Gm9utOqQiKsE2f2J85rEbaLMvfR9/pPP8ghokcClVjZV5NWEhiJQE9cBCcyQPkDR
GnI4HW4QXlg1xWrMiB6Md7IYCy+ZJsN65vkIFTr5K7X3iA8JaEU9RC9rIsqH/AHs
jWFVvm7Sy1F21Dg9zjOh4+ZgSoXmn7ednKHNr6dH4kmj9rwE6kJGDWWO21YRQMmo
SW+PBdOUYH9drVPom+ia/++MizIffkW6JCWvwMQmWCZ3XTmmJibSBz4sKlxZTWxf
SUfPC8FdLwh+XHjuQbzMN1cQI6qdjc0HM+QU+Y6q2898NiavC5hNDNgvIoyNsTCy
Uu840OEV+NeCMgAs1tH+Rdbn0WMR7LDJqkdyr0ShqYWtjY3vuL8N1wLqlYgMZbEt
b39g2UC0IRSPTLeWmCG5pVOyvvIc8yroOHTxCOWfudC/M/fXDzHxDLOjuIcLGHiF
qYh6L2NwqQCVEpTeD/2MWXke5b4rXO4uU830KBWdSfJxAGXf4HDUqYp13k2qlGqV
gsw+ZSYDQhdfgXrdd+k6bC99OU1cVgY5iBcZl6TbBAmBDBFB88ebqhS487Edb/yg
lcbN45ts/nX7VClc+uIGurgH19PI+kphDdnucjXPx3TH/JhExJ1nZQuAGgmxl1Fw
NcYeuRO+Pj4LU0NvfdWZzKKZIbb7Le7uFJ0waDESXGQWQ8j+wG7UwNa2//5lHaUT
Pr2xwjOlsHOkH/h7zTEo089R6o6KObBSr/ZBgvYptT9BT7REyiXx3RSRBm2db2x6
gyl2Z5xrx4u49QT4T0whGWujf8BJGkLiK7PWSaD6l7iY9Bv/v04lQ9IUys2DjuwN
UlTWzRW0pDgKTFvaipZ7v/JsmFBHkA7oKgdl/asUzjD6e8w6UaS5Xq9or9NkqL3F
KcEVTLI2m+VOz+dmUOf0bsitiRCBIbuIZM11N6nUUO4XadKmlw3pMZ5sj9Exdu+Q
y1Hc17SLQl+gXyP7ltvA+vHWFKhdvkO1GBzbDVjSHv+1CXo0R0Dg48kGXpx8XGvY
HxRI4zSXyN5odAdS50OfzbyHnCOY5h3NFO4uw5qyKtJUtnGVlqfR15t8SlXNpDLO
jjYQy64d2wSlO2aF+UAOW0sYxIW4HIzt5y7axu5FDZ34xrASXL9NLI6CPQ1A0+np
coZTIch32HinzAl2Ffu7X2ASihWVmmFx++JnkKWQsCMZp8xQEJezIXKGHg/5Z1ID
rb0zJ6lnYT+QwIxFY6/jtnFlit9stPcTSiwhujDFUvX0o7SJiE0uDctkCLE32usv
jNcHxt5UgbuRPSk4yxk4XJGFuvOs9Eyh7T03Uq4MieNCVPw3hLTKm6CDPtREq6dn
+syJIOsFwVa/8Z/I090RqOyskv7S61Wdnq0viqaohaTf/3niAr91aES5vNmGuws5
1uDSwLTZw/H4a21yD/Nzcm4hUWXtn7ZQz35eOi3ndcyUhX5GaVH7XF6cPvxViXFF
LXyKKZR7BHyYTlYffRP/U9YEH+ch7O+E0tCUHNNkNWALvvnvTRkgBP0R1Y+Hz34I
SglXti1xDm51hVH14+tOL62pJF0oT5zeuI5BcOs53b/DoKgY6FQiUUXEZadC100g
eZmHUEeqafY7F4NdX1IRqX2wttSsX1ZtiyPoez6N+Up7ufae6cS6vO75PxbRScT2
yyVa/z3mcgjAl0t2BT9QoGMGgrpe9T5eeYoiFqvQckZrK5roolNUOMOOSjDkCW8k
AN+dyRpATl92tCUD03avte/Mw8Nee1IuGp4wYph2qmiflbOJt2M/pyPea1D+1weQ
AuKpPo1XSbJi4fdtt7QTprBsqhGEBvMxaVYv6gA558Iv+fFSpDpkTNL+MFDfjuSx
bCK1XrvyUJyC/UEu9JecypCx/neVg/Heb/JoqF1IppYh84bTsVEjq8QsX6lLcmm1
Fw5BDI6vpJHsFmiHC/ITDiwPH0/oWUJXWgPGctMQ7sVenqAVvtNOBdbRbiLrKk5j
ThOOTlZQUNChZRFJm+v7hARGLKoVsS0o63EfT5jslxfaA23frQNJnF2di2m35ncx
8NCGgyiZrA7zudHLGB+jYedvMD1Df5mQCq+KLi+Pk0p9W+mo2W9eREAkxO6ZoH8m
hyXeZw29Ua9XpmdzpXQ0ZrXt8PyP/oS/Ir8/xLHlyEVP8GaiSOBglLinfVk0Fhxd
8SmQGn9oq/R08HOYPdAFNZjsjPi/ji/dcBOuCSHL2XaF/K96c8llmkzZkxG5iFIP
xjUZt+cXkn2rbHILXuCRf/8Jsba7yhuhzimiC3ATFSUJrzaPMPwwptZ306MXDAjX
tkbuzn8avoNNRarVv6BXEycIZp/aE5Gq/e3iOyfSF0FReSnJk/jLtwKl1VatmuCc
I8rOXqOpXw7+AWwfcQ59dIhQFA9p9F6Rtyf2XH/03TH7a1fktGpB0L97Ya79FQkB
CPHSYyrpvnlNT+tOuGGo/aCFq2sccTB1CCt0tAUBUFBTWBImPvzTmX9IFh0CPckM
WPHsmSexP0C1KbuOcepsnxpUnmBelq5pQ5bwK4oEKS7luoKTjcHtip/9/x/ie+W1
hfdxZSDL4+ZDJFJs+OGBl9jFhzCnBDlsqVafS9HvMwFF2y3vh4SM3PpJs+wBzSuG
49scSOLrRTzG5wH0PMXbCx0oQ6A+e10vyi008SMsUHtFRzZ92to2zmMUsWlGEntZ
4RsLxV0uz9vS3eIdIxDS/cSbXCazGnxrZZ3wx4uaqPmp1JEAdu/hNgGPQa97Wm6F
l+RwqijWHSxEdA9qm1dcKPzTPbiyi2pzUjmtldA/hOdULKW1nm73DAAEw7J5NYtV
QqvnOG1T3SOitEVfoF1aEKdbXEeTop6ZH2d5eO8kKQkkOBLGPNZ/X7hHLQF198/V
0eyfTCYEjGYaya/UBFlROksdyUz7gzGQ4XJ7DpjnYwse7+vb4FvD+EUX1ZH2Ctct
TeknNcndR3L77LKMsYpM06G+sZxOIHqJwDoXuK6ESoqHVQoN3ziMGJklTuX0pJmC
ZBuUow6vCRqrJqksP/LzWPN/dYaFJy4hhvON0XYF3Gq9iaqqz3vN7L/hpwzeP/tb
Pm6xeI1Iew4jL+egMnf0GCU0/H83FQVnQedteV5HDSj1a75IMxpn5EVi9DX6T4kA
9ebub/pZN0IvPtbDNkKfokIiVwvjHbQSQsAh9WyXQVbcPWw7/eu9oboZk8+PxUsS
QiRGCiSoJkcV9TKStJ/ey7IvmXjG3Rdj7aqtQvMIQB98yI+XulSzJf9qzW85FmjA
PBvbVKJ85a25feluU/+DugZeTLqLuzQLHM1cs6Iu7tkDKVj0YxZg8Ll2t7w8bbnn
Qcb9hh0yVRsBGZKUPTf+ZseM33u+Vp5bz27DsIXXCyEbOArhAGA4EqEDV5n+doUp
OpeUPT0SZN8XAcmBPcNdIUXqAHA9vuj/jALXnwVFaLxWyaClB5fCcE07OEqVY1Yn
E2XdS/SrICy5MC22u02tjHsH3Suo4Abkn9SwwfCIYofZCrorNvV0ZDAeZpaKLuom
SPCJG5TNP2s69BLGzSeLYpRch3advcuhNsb1WCRUqPzLLxvxOvYwj6aNC9xTAvgo
4EDcXT8b/bc5pLd6aQ9dcizkm6XO7v2zcvGhdcCUt847QfTXz3zHLhtb9rCufkLZ
kBEC7Li6HmK8q85Ebsy292g9Vx8SxcmEn/FsJqg4HQafz6hyGtXwVnOX+G+qG6Oz
w6lXGTr+DS/dkecW0EIB56ifvrLaghngRXC9yB1t89Y1Y7P/lUC3GftaaDNdiHgT
8zMlrHP/oobXnnM1bmkzIPwX3w9ejrNnPHa0cqKovNiPw8kYiHH0+HUe8NdnvQVT
J6uAl2rfPGoExu0X5JyJHJVI0GMBter1q4thjIZVsPY+l6I+SI3Tt/vkdawGgsFa
oZOnGxuuH+P0V4PsoXK5ulRmRx3pN9ZO7NUcOFww6MzrTZMj5RrkM7KdCMdtbewS
7ZfQDuWjcEYqL/KyFM/+fpS7q3mSmlpGAO/Zor8zYiHn8U4uZkLT9RfYhGgV53yY
YCAjwxUuk7zBuXYZEQ/JhJYVsT1kUA0fxz7fON0e3Y3F3edYqF6OQcT4GpQ3FeQ2
iFQR0899Vz/xOEBdY54N7TpTlOM7lE4qBzYqfKUGSAxpHJ5cq3mphdCdiafE6e/g
P2ASoLDeRoS7owFbOIxhSSxVpaM8spvVNSelT25VvhTXbAXQI4UDZDkPKHzS+NwO
k9PN9Tq5GV83GF3DvPxTjyBBQAMhCCO9GdJK4c6FdDWXgoWFcDDKcoftSKZy1gZP
OAFRDDFVf5cF4CKHqNu7yPeuyzZzBQ/lfRmVh16PPnh5dBxgVup3XTnCTcfvnZc2
cLYhwCLKhxPQb22a7ybw+957lhBroEqKg9F1lcY2YX8ph9IMBEn/3la8MuZeq42e
YzLcVGPEFa/zwCFkbqBRVtWILI+V1g32Qvg7oCGe3dX5ZcSWM7voRC/cLblmylHX
KNNvF46gc+SjIOhlO3hk8uZhxKOabIL0WX8pwUWhjEJVDGVOYB5c2ZUfs2yqvwMX
mqbuzWpwccGfPNW3LjQ6MjRrwrDYacwXL/iLoadeSUZiQ0iyX9U2Ji53f4Hwb+DP
AjogoieEGxI3wvszRvvIWSKBegYTUHrxWTowYXpC3bU2SbIcpy1gpDZdcfq7rTJp
7mOl/CdgSHp3ly9XPIAdrw2hXDRZ6RZ86tgzl2H6GpPb4fivkofVz+e5ZEo7nvJ4
zfwN2NyLm7exOuT9XZUTN3goJzEhnikgpBWCmbcsEqObOvWxB0RjV0lFvp4nQhZJ
QMvww22rWdAJFwkrDEjJUGjevJIdYzlqlJlAoa5UX6Uw+4SKo0IuK2yP7gc4IXWz
qn/3iusRZrK4mM1er5gcGuQAUTbP3fgA7KrtWg8HcSkJUKeLAa0FgZMp0//yaNNX
+e1dDD6DNE3btymBESrjIdAce83rbWAUNI0FsprxhNVNqjaXrHCOzEttQcHdJSI3
qrEcjn93TGz/zGeueMbxHAnkkhYzSSub5NScmORohcfWd1qOHFgn1vZK5c9+wco+
05GpbOGEIQL6roVXV5F8h6KMVWc5AXPmGM4M581ISuxYj4+BqywkKpJIweO4hCKK
FhHw8pDptwSTJMOALMs6f8Y+OcvLMaLbiFe7vA1KXqhDAD3CyRs3hjG4n7ws22go
8YVpyfUqhvcmd1nvpO7sLJF2eHW/doxkJG/kAgvj3TwRQzJbSntJbnDPwc+VSrvi
tGQLU30PUyp36u15lkI59fFh201z4OviebSIci6KBG7SuMsNRjPSNyVH24CKJy1i
csyQyumMK6yEiT+qDzmk3Th2oX8MG3jxN/E1g6JoQwl9+8ZPC9JKdstGoWyis75G
7ct5rOUpFJ2iRYztGgU+HqQgM6Ik/dcYH2YBcpNDWhyE+Vm/5oe6mjEVYMB3tGcB
sqaVLrRuL5Vu5IG4vZAbP0iLasplsJbTeQedum+LolzSwzuzJGPZOerPyrYu/4Hs
4YTuyEeh0zL4e2PyRxKXJ/eFVmvvTU1XqUAuBbwwpQZf7jg5HDHwAdOi+PweoKkf
NBz45T0ORaUoBm2SL7VfwNA1g+36oVCCYhW+t7Bb1L0PjC9lhXcAjjY9sSCgqozO
V30itH79YzQD+xuD3vKFwbFAFgjMdSJ7X6zw/WcTqb1bnYpqsgg6zYhzt3Ty2Dar
ZCYGy9adQkHeO0Nqiuz+h74CoqERXTaGQSKvctdhxw883lTBwLiok2UnEND2Sxks
dgDRVyLVhqCJGAC4Ckce8EYcNRPXcIrEk2eXEkqnnMHhkOJ+YMl2lNjm/OMq+b8j
3J3WQRZ+26B/jt8nq8J0NGAKW8GpX2fKFjXjxK7SrJVkdOhEnyGIE1junvJvZcJr
F0rxYep++Od4IUHeXzlF5kN97THNi+vj9ZbtrPRHG9QIBtQivTfd9YdKNHwb8TbD
1VcvWNuwkcioC/WXEMwCZ1H4l96USfta8k39snbGnA3RXDl1pX5DT57ZMt/0m5A5
JGaZlwZCsT5I1dVNZlJCZO1sTkN5r4IEV8064vfRWLWZtOQW+vDRFmTuI9qY2zBY
3YGPo5OwfnjlXVkel4xfxtWugg6s9iseu0yyUZxRs5wEzLG0z1NWoPOMi1k771JR
IU7Rk/gkAHhzIHDDuz2b0+PIOKByYZvhEnJF45YuwFCjCgDIiScIBXhXDnLrpbp9
L/wlbTmtq07RFkmKa77HLr+L5erKd1MV+E5ubgCucTnL7zZhSED7JyEIinoO5JN1
QrCvlDHxV/AftPDqCx9PB11UB6JI0lk9Y0LVUDoUyzQOWyF0aHA03Dp2/nBbshe1
+bB/MrXe58aYcdJ6XBWThhznnoFDcqZDGtQ96S8Ok9OxIfp4TrJp82KNkNKmMajk
QYGMjy4Is1qyOajuFTD+cXVpYAFP6rGCUBHD5AfGnnxksFZIql8n8etA9yxazUpc
KFdCEKrbPHSG+TDlnhqqTRc6+M0aq0Rr1rv8oUEfdIQsHuwzyO5STN+TRaFEmDuJ
abTn3mV+mZIsMoXc7/ewDQ4XzkZ/yQxItnjv/s0S1ZJDrEoQWhVoUJiRmIpBnTP9
mDTr0s+knHOjMr6uvRWVPLHO0ZEt1lkvscQgkH7L3a0/4a3UdO96HOh1C+T1N6ew
6v1L84kYFt55VnKwxVZIi3E+WFH/NA2S21Xa6twN5NrIaZtIQRnqFEvra0dhQr64
2qO+O0oUPRPkLUFlGV9NTnfMkeKsp7vVtHt2S4VgiYniRBAeaumJR8eh9Lc1oAFd
+ZBniXajciiC80Iu4pRQ+fTe4G1quD4qXw4+EsX1miWAG819mToDHIRfBtgIFAm+
ZSILe2shLNXCd3wyD8X6su3+E/3eCRL28wcxd7fAr0yfvtkrIV7b/rS54u3ZxMXQ
PxDR+8j+Q9NSyY0S5v62a1ox/JHVMIspReUK9+L0u2/gZ2ZTTPVqpCPCwrEN2g/e
xHZt5ymUVRvKSqv/D/PNfDNbJa6IoZNY7zvYOQZSUvLQwzsj0UAz3fqE0lCELX0l
HQ71V8T6cBwRX5cIfMq0nOwcDyAeiDgnBwZXkVyEoJfblFeBjLSk66ipU3HuXXUG
3JXcnMzhzuuTR9Sf9cZK+5Jxq923ZxNWcZ/LfJC7skTlB7B2d1JlB4RfIWFFb351
yWcRQfOGyDZYKBMdFqYPTpaUCQzBPtGGujwwFKDgyM6KwPg4KnzYrhSwtP3XxFQ5
DjVB/ytae0r94uUq8AYfKgYV2+fgzDkJwVrCVvq+ZJhgvaO5Ea9UXgu+5LdllimF
6gto52h+8xbDRjattruA+DywpNJo1ouCakMG8TpAogXaaovlAq/F50mDV349JOrS
BajxDWyzGhuaOdWXzF9Qqq5YiKGmUE+gjmoJfqiFoby526i7ZlTC6AMWxA5IY/ak
qonhnUYy6J44t1mBx7sbugGwJSWj0k7lgmFg2fNiZ4aX5tmfg4IPVkRb5llGulX0
8y2n0cFPEhaDNaqFFNBu7X+XCrlmhzKi5g8QmIzSF28J624gOleWZ3rb2qR1hczx
q86strFouYC7CERS/7zTPuPLF7VX+hQKyTYdkbm0FmWr/isk2AvVXBFuyH8s9w0+
L2ynRpWnJp8pTOU0bfO3/gQGXNjb47S9t3FGewJ7cGLT8TCQ5ZGvcW+/4YqkFZZP
bBCZHYjZ9kCbkOZKb80BhhLrMJPS6UavWsGmGrpNCBJIt5uRH6FvytHZBDQnr46E
y9oMFeW8vNSldG5Ur3ucYeHm5Ggtip9HYSitOecOPWm0gEC+cTdYVLrWczgl9tK/
TNTUu5zfmCStTIskSi+r7pOw6D89tlGsHcPJh7BX3uVLFs4msGh7bhmvnomY9/yY
hl/R4/CYjvATa1X68pDjPNWp4+bkYuRgha2YCE+sW+MjM7WqX1yIFK3uFVXLg6XM
B6c0kl7TJ5/z0hr9WshMRUpOWTA+I5hTHUihiM0vSEnADcChZdij4OYBKKPE5Mdn
CY+pXCZ4FpzR1JvCSWGg0KsS4W5u7xhBTudFOPYynfE4tUqPH/M+Xe7k9CYffQll
coGWoGfubIKIz54R06sbKzUamm614Ab8UkhbHZObveQPEegXlq2lWiMPQK2/edGv
elROy0BnXwujuPlB8mUcMdOpkzkN+XvLB4Yg6exSS2N9JM4hHtLS/te3zHqoKttO
TGcAHXimGC98j4ifWWEyLCabbCpR/rfr4eaw3CI2S5oon/Xw8EXZ/hG7oIQ66ONl
HtDAN/ompH4FOJA6krGGJUO517O773t6MlCUqSftz9DAz/nTkzO9BQVzj470enum
BJzQ5qZrMP50Rt/D9V5jvcCT0czzoSfzCVLzVIWPtbNr06qfOI8GbNA2jQDDrHWi
MEEVIfebVINfDmGoA6TWSsVrS5CAZD5ggP2TQ7eP0zEotPRu+QnqqMafinB08KHL
egntpWn93A3L0F9mNGTf+/baoKGf+9G0SWY8/uZnHKHhwUHRB6pvgKyeNmHSZ1Oy
6aCq7ZZXhxy869QPQZWCotiiSrTSSILC9LLr9uuo5fISk0EaAiSiHElvT+BTeygU
6nSyq2kuvad+Bew8NJLJ88DNR6OgSn4U9VhRooeJEpGIGHhl9DDxLTvSCB1xaUYE
DsBPZo+xGdWX3bDecSlI7SEEkImHN406a2aFtu8hdlznVqGNY3Rs6G1cZS3C8fzi
k+uZz6E3QaykhmVLr4FA1FuL38ppG8DLmClMHQN8thq8gFPEO+WX69QgLjWjRfcq
cKUh5e6uwpiSNN37iM18mwN9YoZ0OoDuLacuuINP2/eqmKyLS7djMelLjSC2dfNW
FitdpwFiZe4OG8VPjTbnsnZo5+0SXXHLiMZNFNtadNfsROBb21jOVMVt6IYGsjX1
JGwZlVj6r3jQh14cU1PkU50nr4KG1tIuyiGqlpHsP1U1iW0YXzxidZzxodf1jvvM
xkZ8GCat+BGFoiaB+KFiOu6ebTOhaDR7XokyKqWQp4nHHm+UYgOy6SGOWnBW+QpI
nhABg/HSwQkKJQDGz2W4MUgx6C2b7O8yO423UbYKJA1e1SpokuegdMMcJKzvA3gf
qInYiadIdDuJC5OTOKPFw+yywRXg3ED2WM43i29/JxQ0RrSMYA59QPwdcVvZdmJb
Z5Zdygqq/zF+SP/St3ojp5ZfXRjcN6p2E5+6Ndcm2c17kc0BkEF34Nl+LoivFVSp
yb1eHnSmr2FXuQtuaVcJEaZfCxWEbx0WsUAcxGsr76EPfRWdgiIpM0jAMk3QCTAg
ubia1jpm4WxyziYko3QwO7fyVJJcTI7iatBjywELtgaaOco+t25rxG8ioOnO123L
IIV4GnAfrkipg4KyF1PIhb46IUCm0BRjrClZotshniB4tVBGLHUKLhe9V7bG+NK+
ot8dcoXg5hSy3KqfwnQPbHEHwP8+QYF8EAuqKOrguocfHNz9x81pnjJso/xo0QvE
WMzGzbI54pDHEP4OJWLE/TaRMWO609nNk7htRWvU62uGn6zuGjcUfi6/ZUwE7oEO
SjqVbN58hbLv/eQHPFEPW7iMBZWPvv4Qp47J2uwAgtcfDFp7c8ylZHhu8fhA9/QS
yjqj6hC44Ii6cW1LkIFsl5dJAPtBbOjWd8379X5VxITA9gggnNDsDl4B4POnJHg5
VzE1rQkmnQL9E37mItQ2QibR4gH1dFkfb/O7MoTDi9oQZ9Lx7+nD//G00NLmT6nN
7r0kpxQTMg6PRb1u51Y26sazDdZjqhyQOKP57ZvqwZEu8VQ1UWABtqevTOF4JafY
eyYRNfSKWZUdBXJWAWPFocNNbS+6tlrowMhlZUE0RHw2jE0vumPeKo5BBlb+q+D2
9KmQC2l9xXVUEGVVdUFbZmSNWdVAxUkaY9eVqQ2wmatbDMzKcvBIUmgZZK3yPknm
yfgeac8Ifpidt9h/XtIzZrbRDhhqMawVNKWqssoaD1oc/5fKx0andFTbFzJBR0Kh
0vUHK8Lp6TzUrweqrnPwu/7YTJCgKf/XrDrB4ped9nAno7fymQr3entoi5ARo0H1
C+BASWtqKSv23bHit3cE2ayg7dGEE1F63s0U276CcIJ8QyDNmsXku/e4ZdBbMDuc
on7jS2Sq+/L3q6+lkkhEd5TvDsLy//myzu5+AJCnNF4YzgWqzvWvEuINH9+qnjFS
UJPqgtwsZG+yuyRi2KvXgQhNnG3sybaHvP3TlCQ7JVrt6Ehyt/fHc81PrCTLLGvC
SIwRDe0o7+1hBbhTeViLrhlzcMR/IPJYoTgQQjVCuDSJNtWFUV9lIw7MmmlyKHG9
XCBaejEFX8iIivA93D8ezt8Fn3xEpNxx9RGjOk/iv9brPjLygMjxoND25KyOM+M5
qZnxaMghMX060MLFLqPf488jFjmQvzBELx0eI/LupTmFLlHl/6G7y0TqPmvUxCpe
GVK3V/txZyYxnG0+gjwZZ3Z/Q3F9oKH9CBCuVOC8Us7EvFfxBgIFq+o394WShi5P
d72tfFoK+ldQ22cWCK/WJSmk7sGf75QpLQv5QzEWPllNtfqURrGsLlAs2FMH8O2B
aVYjvAbFjkmLE8Ic0A13R3T3urIljBu1aZ3wJhluykhplwp9GekVVq6GPiC1koPg
jCoKZl69W6F2MLdLUBLGNeM3gFXrFCsQzjNSHVip7Km8ufi5UMvbYGzQXwxCBmUJ
8GbOupXWIMGALdsbSwjn4VrQaNJmCqSwSyE07gg0kfu/Rv+HEbErtHMbVRiuunF3
PbmAT8OHTmJ66PAZc5gFbfzQew0DTdE3ywg4KFpDWgIjOBBzblmjS9nksV3+U5PW
Z8B1JqcqFU61VR9sOvFNBEH/H9r2tqEtVjLcB8DJgiYwZMkLJDDHGFLYaIeuxOUd
S+Gge3lz7VVpLrUCpYSVF/xB/S02ZDG+Mnu+4oXJfs++Pv53zAQKB765YghMJ/33
Rsz0E9IP3P1aK/jCQTWCEzblXi9pjrSzUbS91rqEzl9JHP0mAtms4FvZoTIrFbA1
FMYkb/0xuGTvlzHXH6CHYIfFJpSbW4gZWd5SS8YNbrtyLNH6MV2U0Zi48Q1eu9mD
pFLyz6F4M0b9LXi94lKtN/OzGEOT8GqLFYnPgoA6tuNt0eH4ewpF783zPN893rgs
YlnIZy79eVJq31sUtK16jyyzr9Xm2/jCNtqOb7o7BkqqWxTSIEe/ACMUg+JX9F91
UzLVlS3cBPlWs30ly6t0TwpJz+l27mg7XLyLsKNd30OV3Xsp1q18cK8gDkhvsF4S
sjP3W2aG2wATvb6loj8A8ET8HzCF5LbIlYJZkk/hzGCPvZ6eRvmdviXRIXc+rDJQ
gjEmdK7Lkyyrw5/hnHD76RQqrOQbhvstCyjy9hsMpV5ZXE5qlxv/jIiA7VpOVvMr
r+hiPdTTJHB+nb4bJp6TEFh4RuBQROYZ74P7OsKj8w/d1q4DhTh6A4X2wOr+QWaS
2N9Y3JDygs7oKmrR85e13pKdy8wlISfAIiGdyWYQ0lsWBEn+VhbDBOMd1vfkF/9H
iM4y9ru2Gw6ZbiDTu+Zl3C8+bMHDKyIpTdXWehJv7fNIGYOvWrFx912lZFCMj9tC
Fr3Oi2NepUof7FNk9eifq7+uIoy6gzT5Z+x2EXArInPj/hLKAi+mVtDM3KVM+BIj
S2OJm94J3oi5bqj4jIycthCFrJb3YyDEbNCTsLq0t2CMx3P85YH/GzeSGmpn4yZa
q9vXAQF2F4PzdmuHb9FWXOfLWmcxHoDDPL3GnDIXUAVit6Ujuz8oJNyUDm7S4KoI
NDIm20db6VRRa6s4FNehO8EjR04vtjeiHcfIeWviPpPxhhcx8L1aCx0BXdbd9MPd
uy1RS2+22HZGKXiw4xEbbyoo/QKhZ0SDr8BZI+NeHjJzmqrogPSuUwG990TkqXZy
Mjh69MEYCxJXtpZikGNqMF1nMguKTjRzuY/GEf9IR7kK4w8R4YfvWn8FPmhRcQDq
Fe1REYjPKn8MaB+8kDffLQS0RqAlBH///lj5OOxLXuZZqPb3IbHu2OBkT+D1TOhe
y7pBWWQWO+jg7/KMnPuddNzbgv01XAPiiKWSD+beKKCDAxH5V9Mzw+SeqCNAV+3s
v9JUibMDNQI2dfu8SoSIyQVjnkqVThTvhR+bx5KQU7m6UzagmC6HfvekVjIaoEsN
qd+I4sArpXmfPy12AWgYpRlFxURaJjJEQZ47+mlu9d6K3gEZbm/u01mNsEHTfxIL
0Cr/tF/UB0r+MJbnlBEn2S3QGx0jJ4AZCWQAvpI7qb66IBVbD6ec8s4pjQwMGWXR
HduVtXj4BMWDMTWk06uJ/+Q1SG1LckvUwOELRuKiW1hXCe0f2IyzpPRJJDI7PnKg
Y1yNDiAmumqHfirfDwGdtKVRuref1rkdTE8goVyGqZiw/qce0PqH6qqM7+3xTkmN
nw5qsjt4CRvdHg+u8cfSjZzaBbT2D+IVTIWoL6LgpBOQewKa5nYF9LQUI7oiFAJb
dW1khVpJzllIjgvAvxTrWWUTjRRQcuw/7QitcUDlIUAruvp7tRtyXKlzt4soGg0j
vsiMJLsXBkOWN1QqC8aIu1O0+Fe6lVfqipXyH9cxlJjVcykt3v/wzbdzy2FLdfjB
CdXzi3seUJzStCi0GbRw6vBvr0XyZH6x8iMHC/1pme2Jh64/FvEpycwe2kTWvTLO
4UR9HrIyzDX3nmpT2ta1ft5U3yEjt94zq0QthAb5c2QHgFOMICCKCwRiYu6iwLsR
yhFx0DsGH2fm4jvDXb7qCh2uzUz1vq+4Fc0Pvyo+Dw9f8/wllrstl1ZXjMCBjxYO
bu9L1+UrQwGV9/+hOxWKm4Fd7U13b2mCM4X5GF38IXv9iQnHNCGlhnAg5eWVl1jT
CJL5+XT0f2dLB+Kd76E8A9Qjks5qINhjE7jdKOWeC4BpPwL08+zQ7Z+02h837bzF
zNl3t7ePxjc8GSm0h50L+YDVndhJjKhtzKGqwZ+YiT2L+yIk+iiN7Gv0X4SUjOuk
cFjeiXu550V1XMRqYi4mKzS4nj+zjthg/Kuu98gkKBjdc2qs1K+ZmT0lstrlVSda
ckMCJFKsS22YDx+wf1WC0/mesFwfloZoblIWeR1S+IDNB+pBkT5VydMbcQ8uG3OI
aqLds/iSGLE6M0ON8E242X4X56YAyjegM30NADSKq5ySuA+AIa/vniqkvwLwsisR
Gt1gp+WKNsTxsdil9qbmK3JDbrspn1qT2BqhPuFKV3ikjMAu0vBDa63XJ9LFoKoi
xLv9UnunLyPLLYUyHJjjPxLbIYLdZhyOYiz4yXXpJvFs002dr64X8/X8lKX8Re+m
ZtJHSypESVnJZrPkt3D7mocOaYL5xPWj89Q5PVRSI0kAP5anrqKJk7iVfb1bzreZ
mcpWzNElIzIh2wnW/NR7VS+sB//reYWf9UvU+Z+Ch8i+BbByzyD6KFukFVdVC7YZ
bcmemoF0jzZFH73PPylAIyoS7P8L8HQGClm95VwhuNtQy7gYRF9sgNDFY5QisH6Q
qFrEbuHiF5pmfAmyZXUqXo7Rk1NQKCdYGg2fbQQjGa5Hakp0lEQaTcQ9M59T2gmM
zolKmHoJp76aEkNgM4169YhIolbeFQq133O7a4sSV9GkaLD84KonItlqHB8U1CUV
ZsPdvjTHUvObv18eoR8mrRV+zSL8KROxKHS3FtsJbTQGpmxnt54Ep7W3BIRW88tK
LPt80WZlZEU3Mho3tXNZpjd0i5kYVgzI7uo03URxqZKtsDQnDoknlAr2YFsrpdJv
IQbMMnNQwmye1KzzmTu3rv4I+zCGZ0ko6QZnCSxnOmZtqqlpjw6lv8PkN9ehLsrP
Siw+M6BadGNwf6nEZZcNSg==
`protect end_protected