`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10128 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
VKWNRQF+vfUNEEp7apOJOdNMPnd44anEzICG3liqT8gpFhH8LWbLG4STT0ufgaWo
0zZu1gkI/GizCabZ2zQ2Gc+wpYYTJ5Ho4+eCPH+YqGfa+rgHisjod/Ecu0VZ1WQr
gZigtpTF4Cco8KbjJxAxgWUZZEBTg9zih3oP5lDZsrhm2nmBh3MrXzFSvsizaJHP
DGjiES2hXFScLJCyMdejAFWnelZ+Gcurv8rJa2ncGCxR27ZNi0cP5A6yh40KSBEK
yAH6kgphcyjq0C9LFvPECSQj2kRjl+Itt2Gn/AeF7tbSo8FnwkE159etmHRQ5odQ
At1p1CYZMi/IvMl78lQaIGw4ApTXa0i53MGrtrPZfTC5CYRBA35+5IfFpljfOw+j
pry9m/WXBqY7CxMBQTvd6hpffYjtETZlzNC7bd2mhcvJpuBLNMYhCUsxvVhfaSoG
pBI/Oe1+9xDZcmDeZ3IXpWJEkP0ymlSKy5rf09V3NSPIJvszDch7sxKNSDSh4SnZ
8sF2SOn/4vtvEB4buQBC9rS5sduIikkJyf4mNR1nfKfRCqKYOzy9pnDV5FqufWts
5PhjexC58d08K99APwK6SiGar0S64lBpLtT5yekNXgDSJ4MT2CH0d3MucZkPEERi
1mIqiZIuSFvnbVlFC/Sdk+8VixtUUHsidj9jW0ZPUYsRc0Ub/Gq1nzKwTL8eRosD
1w4V8b8WkcOf6RC/Ri1Wsp/xsFFkmYkU+IFyBjEpKWExoML90e+j42iLHI/2O34z
n6bVGzi9VuFz+tfebCF5nMPep7ir0F+jbZo1yK9XRNs53GW17df6ke0VdPZsYxgW
8z4VgbmFxIBTG/ErZvtUiY84tqjpBhXdJmWm9OC1/FD7f0NSNXEUm3T32KpkrWQ8
oWThCicSh3gh5HidqvDFBHE0fejVHOPm13ZunrS8OKNIBZycdAC+iD71LGvy9iG7
3lgU1TKsbEOOGFFA6qRqRxiu6JSo3LaB6uhiJDlo8Pl/7kaDRKW29FsMYDJww04K
rvIVf8cQAycmwj+eITbasO7XnWFiEZ8Xg5WcQDOZHInOdRssZvfTqYEScFzwMunj
KwxUgGs/9c+9/DSzsR5i2ESn4rJW4PlYoBKQTatoH0EDLcfa+53f12DSo+TOQpCc
gS7soIgLEtP0IGOVC2kkmmwU5l4RR4ToqeihAOvudfewDCEveTCOINwAekPP+wU1
q1arPlRWA+t0wuXb79MntV8kprTrvg8vU0rhXyj3/crj4LEmZ/LAsaYRssP+agOW
K0DjkClHo6pjSJhts2AUPbJtONw+icuCF9ORlc+BBl46lC1eq919q+79svtjNU/d
IHfHOHG2iW+hSQVgPYm1LhOEOcQ6YJ6FNvItZCu+R+qy5NsWC0X+7H0o9MDaZflv
X3Lz6mpMGvOKU8LvrrGfS6Pc+vuI/vbLcmQ2YNr8j+jcqsTVOINFzSujiYns+YJC
ZWKeLcYqnRO+UPQgxfdML/lTpNwDXM8OLvgKL30yhNRF6f2Fz1niweKGIOvR3hsF
bZT+xPZdyTTNhfYEDDjrHvxw+TAtoImlGxaReeThG92AFKzLPUxBxM3lPxaXl2qa
VMXQqoIse5epmcDqA/6qlz9PaQsTBYB9KfCgEzuIx/Arqh19s6WnMsfxZeshRjK2
sMPg7CyY+Z8pCTlGyVS6F9FW6n4CazmY0jQk6d4d2d1rCzPAeWcV6X+Di+okamoZ
nfHNiktPOoISWXzCPMwPUpjYoU+n5GFFsaX1nbIznUgvnPHYWLS5+awg+rl4hszx
DzGWG1ofv8QD9x7NuXgMjr+7UZWe8trLu2r1pF6GQH3NEwWw4X4NcEJ5va7S0bbS
H/AaJuPzzL3dcvLFagxlsVWFX5uXzaF8MZuo9POi4XA6SYmwF9O9yXYY6+HCb8+j
BcyzXTvMV2b9vSTquvCXSXiswVwmLc1bMdIDeT/WSS2J+zXa+SBfqcOaqRBlP19H
o9dVE3D2U0a81XcdZsRdMDPGtk+n3i8is4XDnIzrl8CoBheOvACtE6LzIXA5obck
aivvkkNcTsp1KUw1P0DXYx30RyQBHTuWYYxFOBsY1w6QWkato36/UQxNnWLPT7ue
PW3RPkJZ+2Jqil+mbi9N+IiiI5vbH3cEIptpFHUM7ga1BIghL6OyRSXTiZjJ73gW
2QCOmYWjT1dZ7bBFFL/EiySEoB1cUy8b59efdM2iUhNJM5f5UMSAvK7fUv0fB4Ne
1d6Lro9omVsrPt90tQtdwx2LmhBiPFHpXVUfOL8DbDMdUvYQBh8nc+CKln0BMaPF
2S10QGY213DEnOT+xr0KFSl0B40ngCzmRDPF3lj5Mrr0rET3PQ1XldL5j1H3IMV8
09aayL7y97B/U08fhiEWh9ciHyPjMtB1HQTjaqBOBuwLHFDwq92t5/R0E5yg5PHX
X6M+ww+En0gFH1l8Jp/+/V8a1tP6JcNlTFxBGUt6LG5HI5lsV4/q/5/iFdcfCZpq
WwmmOo2SfAjT5ruxP9T8v/Cm8y4ChSHlw2vC4o4E8pnImpudMYe3NHSCjYTGuCNI
fGSdFEpiAo9fAM7AaTMFrO65Brbh7Be7A0Pn5uLkXYTFNXmAnCKDMl7x3mRhbuwe
xN9K9xPzFuFx3e2yZw8c5RAntODra5QhUDwfHaqIXF22W2/m7Pn/CRDD9mCisX9Y
WU9yNSjCL+WXV3awv9Z+0iXweS0YxHrPYa5zkH6BrCFq02uXgpt870DVzOMoC8qd
KwiwcICkTFyid+JmUZJSpCKU11+AfZNojFnKifhRkmf7keItmo8bO+TZ20tQBVEg
U4O+FWldpDRsbWYtQhnrAq30ixuYMbISmHXc47kxaLEnz5TBV3PNDmiR7kCD73rg
IfOWylontzx3MWS4I55fY7VycW/GI4uBJaJgci/+1rX9ovJ9QJ0CK882Bdq6GZxG
9QjwOVhyuxQFc2CREyp4TIprDO7X7e7/koz79h9FyTnnyQR+tl1MOcT7G8FqDXka
2fn2Z+4iA9EFZph/sOnN8WDiFHIbue3QUW658VtAC55Mx7ptHNn2PP5lv8ekzFV5
MYSLsjatGdFAJZL/PG0CHnvyvy9xW28v+ylOtn3DMQYRc1vFf/VdnX6g7You+Lkh
kj7J+WBNxMs49IIbDZs+rEFWgGtbD+NY+KA0s8iPRR/jKV1JfHbDLcw6EDDn1X60
kpoN6gi8+CHCs6f5gFxXnjUnKEtPo8LOxVFw7jCVBDSpnMvGH9Oo5Gcrb425uff2
/m+gaQQ8upyaMEtq6NZTLA8BfnFnOTvTHg0WcgkO/yG8UuAp4iW/EL8I4EYRVyHr
KTEtAEs++VE2NDO6SdRe+zbRJDxMaxHe/gzNm+TImnsM41fKRQ/S864+uIOGW3Ng
VcfYlV9etiEHC0gGhZJKXV7nJg8L0HScaFutztkK59P0/Q8yoQV9v354B78sIsEG
UVzODj7CrdIjv+yIQX6sLqw3iq8Rk4qGyWh9vRIAmwqXOocAXO2l+NaQI6JWDfng
Rl02KpMPwv/J3/aHHXZYgSOh6rdT5oLd6FrL3m9XFEvFVsXfTgL/hzXE1izOV2ge
pqWbz3D/3RqZG4SP6v6cPNNULvKs9RbwLOvjYkFZTo5qEUjnyvY54FTpCwZ8bQsf
+RvB70ebii2a8UTR3ZNm40mM3W2/fKLKnvOZUvUsnrjtMUldhClluLo2H255vn5p
euBwpy+L+uN6aFDqAoM060cFA/rOOA8ZaGjlr5cySKuBFkn0kTMVEElZQWcrokNh
kXhdZ/91WL9ACCAegnMprlya58H12Lj6UFn07PJwuDWTDt6Qe0tvOdv8g5kQs6ad
cKsbS5BZ+opPTynKLU46dIe+CMYVp54mKnmrlX3NhsWVVeLjVgyJ/lpwbfIH7qPy
XNjxVm4/2p3yNj/LsX1leeRFIRSY0Jgx2ruPEX+0E95xKod7b49zZarRi8GIMAdq
+zc75hKbdCeyg5W5E81GkgCS071qIIeMPhDF0784mG8+U1YE1f9ncua8w7C8DW+W
gHYpwP0gkT/ZUEFFyAD3pSPOEHVpMUXI/HNSf6qTLLoiEuhRgRNwzYlPVYomnVLg
loS3uJLgX16RKwWguMZq25/rRX5wIAhWRieOn9f4T5O/p0+luUoBILzBM40DnW9+
9dG4m30MHxh6Bkv6U4Ad52Frd77MYqTzg+A5OPLpH/KjMjQcXCmVprZHFm1zL8ew
TfOgS4iX7esed3YBVtY1ueeVVnS/XnKnukWTOcSb2rwfnXkKr+H3lFKurMyV+Wbv
bd3+tqmV6XIz8whLPDPASrJArUft1VGl8HGupB9B56d4Xs7VXhRzuOdErViCk1PY
IenEkeMpheOhjGrMEjmoN34Y6Jd0ufzHqI3xrHIZRcgMjL8GV3IecbsE+d9zSGeL
rShff3dILU3pVjT0nCkbTY5bjMizW/Vpp/3/i89x6ejlsSNdRTrZSCT4SPWAkibi
UD8sczscfEFe2ycwQbA/aOTyRN9XatANVEo3/I0jmYrPyOkg03d99fetxeqt4R4l
/Q08pK6UDZL5EAwcuSJDQrHphRX712LcfGh0OmwZz40RePJy5tGZpcNKhXPS0GpZ
Lf0HscwobGjVNT5tfj5hEd9r00zNEubA+QaUkCHliM098HaI4MwISDK0wBnypcJq
pl8cQy/rF738hdU1B03QBL3jCc0SxlSEOUYP6g6HfQBUwywqty6+kMpgmEIZ8xDh
RNKcJ7C06dPPehNikOj7FBvNQcpAnkSYxXCVyBrUDkWTRSEBgI7M5NJN5sbj1O0y
rz2oSnd3MJShrSfCzu6lw3cktxpYKTZgRQfb3iSUBifYV5HX/3hLCxNf6dCQOvkr
FpjcZ67Gx3DW+jT+OM75QDy7qCtBOaHsMyiGz1xrJNpsaZAyAWIIfIXkc1kvnFRu
XMBw4JnNqTj+3nvZxTDaElOgGzFPM5ZAWIXkVAMyesV+UpXr00NpD40xlPPPQqTC
QxiFdRcK+SJt8guQz5ISPkzsItvwbMqV08lguieYUyEOj5KSL6JNTwEN8hWSlJ1H
A3o/RCi/mrGuWmugQplTg1Umd0al7/Ir7ZkWeeHVtcp+lXTDy1KjJZGnBhN3cJlQ
N2M8BFIDUEKSNrLf9UyUPNBshwWqkOa7WYwq68ZpvOa2ao2Vze4ds6yEvOCgn2UN
uarrBnxVBCQ6bBCZtryuBOGxEMkP70f6OwqHfqPvMwr2hs/ilRiGXq7SCtQBJ8Zu
y6H3dNgGxabnG/GmyGZ2yIYtcmSHr2jyFmtnpjxeuNoeOC4Nf8ovBsFMDiJOP3Or
7bFixZR1hXyZgU7HTkCAMV/Ah/Vx5DNyBDGR980UaJIO8n03Nxs3UvU5AClsaFk7
b/c5m/V1tnXUmZ1P8klNREHZ+WdTa9Mqa6cDtXeKJmmimK0WDQB98TpMTmeDM4Pq
JGrUc+gHBib59ZivOWEqj/rMv92pgWi1n0DsNMa2RhM4AGLfuENOOSkzPjGP5S8a
adU7AChcSTNKCb0WFK4M5I/BSKjIcFtAn1CbcpTC7YhdM5JqpKWQx40LY4VEckG+
T5s4wIsacs86mD+pTLZRK+rvRoeBERcboUkFWXrrxzuxEq90ffgAST8R/KbmO79g
R66CATAhCheKeVT04uFY3WcGwyR5JSrBvbeEpTl6d5EJ/Uohz0JJN0XShhnQ2210
SXr3GqEeWsdfGLiYWmo+weOfGgfDTn0MyCI5ge7keKGiuKGqLCx9o7wpEixRnciY
FeEuO4wfwK2wAry6dXuU7xwJsYwlU0i4T5VMjAIv/q8B8YAXay31j+I5BXSMYteg
KtslfW+CAwQdvQ3UGoxOgvjrNkhjkE+lzhIV78+qK5A8Wo7WKU/cs43PRNNrF3G7
AYCCtqxVeDW0OAAtjLs0+G7peegEIpihYHveLJWqLOnXknKauddkHGGV8buHRYZC
kzQ2NUaE/GSyMnqEpdH6ksaMC8rThNodJiI62aj7UOnuvFW38jSDHIsbDbBbR81N
EkHqc/pUL2f4Vt25TiUe0R6W47o9OWzh/GAFROaqVu8/ARI446z5p2Hhb8nM+tAK
3ut/d3Xkjnhhjq0SETcsCYEuUNXA5D2e/9wo1ZIuQR+2KE0f3HJcRe2E+GnZkrCP
Yfou34DX47WK2Q7ULKRdrsVpsjXd5vutQ5FcA+VB3QBgLh5JrPoz7tM1w0s4SU6D
3lrLz8enFdYhq2oieSE9R9x/zMv7FZLGO1tlpkF5ZHml0txwfBjVMoErePyfWME4
CdgGjzWcC2QNQaSxRlcrRq4FKgaO6ajSZnoufgiT7BzxOvedTrsjKyaT7m6N056H
uB724Uuhprh68RP+UPiBdrdw+df4hmW2b0C55dUaNB7aQLDluENkT05/joE5DrSS
cjUCXEk2weU//suan662TFhty/bh/lokF7YkMNpLNuOb06v3+6rX5+hg7uFT+Ali
DL82ErOMmiuAmSQePqmPzEGMY9x9+1PRniGxi4lL4WhBsczCv8lt13zXgLJqNF1K
029NBfER1W+dE/cJA7BhobAU2GotFyDPOOW9103zrpjEr3yiQRI66G88HXrqOhh8
bzrmlSwc12+2RB9zQ/29yf7F1bhAdGoVqFA50a5WHjhv/4xol7dmTC4fq7wCj9qp
QjeU/OrHDDRdTinukqcnBj2/QpcMrCcgP3b4zIWnbm84oKH4w3ludgZuTF6fJez4
iHsSAdDfqFVr12UGO3IvT3AvSu08PjajgScckze57IzciIE1MakHxmbaMsi4GWhS
HdfNOQkQGsmeBuQtOg6qj9Oyu0qufalI88/89gLnX0WirvtXW0FqnU4q88XxKW0l
UlRTQA4QDvyxiXj9NbDFDw8bAJIXCKpydcVVtB+GW2xqjXQO8yfPVMW/hao2AdDT
QTUuD8OJyGueomAaIXi3/09W6MPIa1Ov8mv7r1Yxsi25q3oI3XcE0EOQ65YE49E2
SrhpQt8NtddsS8BPnxS+ObleYxxfyyXEUGlcuM1dnOaOm7jKj3Ip9RaSWSfc6DZd
OTJi1puTUozitNZjqeuQyYPrPXXpUcPr454x5u84tc+2M7xcHC0e7ZfjOY3MDGrK
5saJQNgQ5jB8aTvcgBI/c+jsAGF6NXVhfF+F5qpIDM1IfO+jHS8imDU7d/WF0iby
BQy0JVmtW6KnR4gHYk+jotobnjbkV8e/vtkqdWY+qv/mfXCP0AsnhFwTj6q382jk
vaI+ZJmaHOyi6ikofIjMKboHmHsnPlaGLivyW9TmqRcOM+fA3OtPhRCFjupFlLUH
k5tEVkwgbQDvr11MLGSC5LEoWU+nEGkT/EgAhV10Lnp2GWxEg+gas9jcEpXlhxqZ
s240ZBafSgigrFQQJ/l2KonyIKxDLDPw5GCf3j3hCGmpyScOA02V+S4IVTsVJzsy
K1BwmG6OTjZRr4yZMThLFNqivUQ9TOH9Hv5NqbD8Y2IYVCly/RKKNLKwW/gh6PEN
q9U7oAZOo0h0ecMEyZYATZ9UPLsJcCdK+Ihlm1EBM5MYFDUl2vvc8NFwuDZ13CkF
HzCdHO1vRXmalU6BGc+X6UElflbnBN3jiiH0sDbErbz8quq17B8EhoR0KBmr3UYi
/rJuxFFeHUUmu7BbATRVD+oPPvRu7Q13TJfl4nye2O03JxwI9Gh7BEdI7sYE7u16
+SCd+i0xPO047O5K3Z/TWbmTWwE8dg+08zEfiOoNw+3SUb2Gw9z5nE8m6E9t928d
es7nmxrRAFPNRI2yhI7ziTnRYArhWrzNobwHgCUz1eRfcOQlldw+YjsIvo5Js/ns
1+i2YwsiVr3D7QXw6okC8ncpPLYqNzSpQ+1h/kXGA+7Tp7SHKIf9HhK2OzGCeTzQ
iGHb06u7GTU0vAHrQSCb4Ip/KVHzp8A6HWD7O7gxesK8oukgOQdpzaE/1WEpgzFx
X3Rs3cYKKvmXhE2HCwo0ugT2vofm5oFaS3oCrcU8y2vWpamWWvlDoGKI9sP8joaM
LTR3k+QQ3TlTL9J4Vl/jHiTFp3/uvle1iTEHw2olUzK1QUWXAXKc04c1SJgemWRZ
EPIhhf5Vg0hdjPeSz2Gre+a/mioS3dcTF1VAtGDqVpC+v5Uc/YI6SPk77AeuEuoI
mueRbWPBAqrpHqfmYvCWQwJ+iSlpVtA55TfrkLXZXZyiqK8Od/Bxxi/2M9lByOp7
q3NO6nI3yn7QCBJBEeYjEOsfg3wsrQBJOAeYcyyrHBxXnCKX1ZLpfZ9DnlJMSI3+
NQ9ITBRnGmb+N5brMbr4gq+em1DaxC76hqTlWVy2qkmmB/TPnTYi5JK0VMu+2ScU
6e46sOSOoSLGs+lUR2F/LNWfENg+JBGT+1b8dfAvSVmEVleXtPGozter9ImYEPxY
MahK8dQx4NXiJ0wD7/EgggQaosa5F7W8I3EyzvdML3ta/99ocbakB90TBzjd9AMn
GSkaWg9jvuWmkkMbArehg9T7bAkwQlRp+Qhwo7Bl1SrDYNj30LOwNjBujyMsDyhf
EkYmYMh7kEzRyE1hCYy6gWGPFmWQLX6XhYcd4TCa6sFDxTObP6hBeQ66AH76ZZd8
CMCpVaMhM+Sfb3Ss2ATlLbXmP9XKizgSpfD3Wc8rGmD0U4TcxyB0xMa1gvvx42CT
rYkV3e+Ue1KjPO1QPfPvvUGBdHi9k2J53Uw8S9v3G/QYkfR4gJNLkYQPW07WKAOF
C2tSC3Tx3GMtUCMZ/o/HuroW4hPE7Q3wIrnbDwr8gScW8+AdtKbzqdXg790ao4pu
txxNKhTBNHPA9ErrlrBsytcMV/5njRWFP0du1xYXx2MrtjUyoDkR6RIMEOkmyhQ7
6qNPF3TmMbwOHPTNNOKGPaRDJKbjXrh2PgB2wBHuFb/rrxqOpyqNxkBDqkquvMWI
s6/M6AGgu4bQADfuUDpo6LnsokTrNGbzhBGS/neLMjHI0S0xfHCfhX2/v5yFt4b6
kfTAjWpMJttW6Fi6ldBO3ozhRMuY85PcWfgMnkMGQlTXgvKuc2ZtEzLSQl4BQWv1
HybHpzU9Ir/P5oWN+d1TSePth2yR6cxVSR55WZfPCI1AnjSqaFTV5gGhyDNbu0oc
ZFXORS5VGzea9ZSuyX1L3Uwy5aPtbj+JByfUCThQABdPKBT13qvXcr7s2wv0VGVy
Mb3RfCtTcJs6J3MsBOTfwPCg2wzFjZzyYayQNtjAo8zlDTIr6A/K7jM5DN8YFC7M
BuqUEAMV4KoFSO+zBhv9iAeOqLeoET4C1DU+vpfQvQDaTPW2Hehf0wBd96bnBPvB
Li8vBUAMbtaU9gRAhgzLftf+kOCxDOZCuPqsZqTr5+NUhcLQBKGJovdzh7TAOYQ2
NEzRq+QzFFmVM8Fj7QIoLukozO1e2TNyOaE14o0L51y6R8rhRyftuy5LEXkpYoll
F46ZkK0d3ZtKGoS9P5y1ZkDdPU69L/zdhk6nAz4hiOXxlTA2Z3UBlxdfQVB1jkf1
JD4yekVRwEsmKcaf/fbXztA/ZWuT9AV1n6nq3UrOEKFh86Nlm1F9Gp8/m4D2DoKq
6wFZyWvSKnIgeRnWfWwGII+74c6c61bIt9P6a2NFdi513TqqZhMgbsvgEnVxIqLO
vhZQS2eLDRh28ddoTHAXAFamu+MKe+AOvorKBoGHRkNg9FzZsLi5uPRMfbqgz7i3
4iErRv7SbJjTFqGMLKj4jUw01PBEwQvUVIwCKetnZLJx6O4oj0Kx5/7G4d8H/i3i
GUpIWEWyqAZxH4zymIUn2FMZi68CXXRZsN72jGD0eZX3JrYIaOTcKVpV4viYt5p4
lJJo21vzYvDsJ88ABxrZrXznv3/4xuV9R4vVhqxq2WHTzgaEwXVqtHA8NvMgWd4n
UCmeNrPkxBHE+6hs0qpBGpqKH+/NTHYPCTB1E3oesHa62N/OcAD8AHUFQcziZ1S3
l+yGVwhJjMF6aY4ncHNvFSK9jNJos2TyeYUuGnqgcrb6nXOQxtJFPxDnInFRmnmn
z3FKi4QLURSw+ZQoi4ulBt7uveqXTlWPKWrqYW1lCg0el/hkwXuCZxpexg6rlZ3p
vKGp1JLndEgE3AlmERBvKfTwUZFrEpovcK7oVGZXDHC/cBZHqIu3heZnIFK03GoJ
ifVm5e+wSqLBbA3+lhpt/i3upyYIcYwfpBNFCF8E9sw1Dd//AcZSITXHvxAcT8qo
N0QeZVBuXuHjb0mGi9tREvxXi4pSTeeXKFWuJg2E5uqlJMXFtcCQM0wfy72gpPjU
2A5P8ocYLZaAUfBBJsQhql82dqJtxTjQw99wCbR8szcbYxdE6XZNvmWQUj3NTRuK
dCmZUttuK6c7WghNHeuUwvXpoUoqYoyTwQCijvlktymCruQ5XuNeoVxqd2Yzw+e+
5ug0bCrtL4PbgH+vy9rGw/A8JW118VgPz4kj5y3FSCPc6i1lfmVBI9o7vP3RIoCK
tdlJlZHdR3Zv8J/fwYvck0hA0fU21H6m+ZMaD3huwJS7a0wSex/t1gcsQaRn5EVu
QX2coi87+2/8jhxLgoa1ZEMPNfUyl0z2LcL6Gs//VqIO0lqc48EOqfC3DSIIuw7z
RbtGkIIMjmgATYOoGA+YM3ZPkcTg4DEEPJ6XhoSqSb2Jr6/pmlcOu2X60QFd0c5n
4juCqAHv6tzK1IMflN3LYYgQ/irSbUtFrhVkEiDxodix/ielJV5T6jmbypAV0WZ0
yA8Iho5emw3Iw9/rUilpdmPyscAz9dcs1GKGQHrgrAK3LkZsP0QhOsDpvyc9HGdl
DdgVxX3o7edOaGUnKe30eb4R6ILNO15+eZA8M+LAKf138RRCAaZBv302KykYbQyW
jaWv9ky6maKAJ0/5AQQrTz/iZBY9wmV39YN0V63xiOg56INLCekYvrag5snPsPLl
aLZfMoeimufcADlTBCPN20EOU3j1//lmlhDXJwerE+tbA6v0mk0DU5gToFQXaulc
Cyp5vN03nU+rE4ZGL5wHVKj78c6U5Ok5sGEeEESOccBHQgLOZlwHKiRwR4jdNQiS
ZB1/h3V1kdVMQeeNiG/IzYnq0+pUqPaCwOdEuQyxzGVfri9HAQ7uAnjpzfQSs6tj
XYTC2laaA4ylhreWW8GEeNdamU2TxzSSNjmFLiHOdE+fWwgF2m8TJmqS58VVs//J
6zCCnxwuJ3kEQsO0qeaj8osaKHG8/rPzTE/3sT0agW26JxCjMd1r8XkG1rpejV/A
fnwm4vkDh+yXCjfz6mpCbdTUd+BkN4FCyqYyvbrYrydz0xQlr0BKMnQ2zcytVoQ3
ELaP4vnk45eMZ669g3qFcBaAQEBwU+aF5ikMsa9AePk1Fv+m4YKPqJcxIWTPYZPh
hwbdAF8yfp785LtqcE04r4AwSqwhexdGNOIZD+yQT7a3g4RQ2fX2bsj6VWB8WGMB
5bKGdDEMXU3imofd48H12J2hG9zqALRKEePgkJ5QkNiAEb13wrm5AmxF2I0hYhI3
Ze8jz2Inn2ym4R+EVMGkS04V9+cfgxqP6US/Mvb4H+owxfzmsWZpewMgDWwOu0vZ
giSSdQ7wmP5PWyppDzGmmSJv1wtzOFpOMkr51n6U2s4UOj1f3WfPqLD/gBcjw9A2
tcpJJpTkiu6ju22YR0GMCqiFKbvbcvzzZRwsrbqhdVbubggimDOkcEOESAR7I3+e
os1yQOzRGyg9ie67qGAdubNvjS5ha4RYEI8Y/gklagohKGC6rqFlDKXA50vlPCX2
i81jPEQjPR2pGvXA+gOxWuetxOkuk3xVNSmns3KkZEXNfExa7sbkBhVb+ynTkfdg
IlD4SMUSKbbfeRQZgLpzSNEiYmsylnQsRu26twkkdaFUUYM6k0bEkT6p97UeD8wf
+JwxjUj23mZHlEKXVxB/s3VfbwRHLjyfW+enYMmR/k1FgrT8C7k9vaPLB8HUJjn/
Ix079zB+zZdLlCtExe7MlhArty3Toc5qtRwWmHcpz+6xYMEGW7ys8czjof/hSBi3
M+oGsYiQako9rV4MIwCNv6zHj8fsgxqTyG05XU8WdzdMC6+jsdmt4iZ/gegsiK0p
HWJyF4SsHNIKbrBJR/tnOmxT/Mum98J4yNkf2y/VEKpG380VHh7iJJj0btvUoUAh
O99b0RF18xuXPonP/8ierpauVSrQ64xKKY9Hxnzmptk7GMSVOlaWcavm0CakSAGS
7PrruJqJSAz3forH8BhUmKCoPvGvb3+3ierJ1fmXVRCl0g8UVNJ8CQ1lfPC6UhLu
eZc9qqfOoFm0FOu62uymwfsvZprNISSNUbk9kWWaQ4MPAB2y+/nL33pTTw767AOA
7H5YgFC4yeCrPuKX/XOGMVCumUZ7zx8C/P6stUHGTG4LEI0h47PbLRgi6OPE/bEc
9MPCqQShnJv0pO4wMcMVShUSSzKypNFxxT+1aam0jz3nCyK5t2MlX0UFBgrjCRFU
m0fgdkkDzeHG2ZJTd91VOH8CleHbWLJtIrnnNmfT4a37p5RMOzJSP1F72w5Xwof6
YShX7JOwHGcC5e8lR9jyDyks8Imr3rnroibEfgdwI5He+EjxG1US5WAurZLcV3XP
MD/j8ewCgH7Tylepkams4QQ/QmdDRbLsvFz8AqiH7oHP5+Yhp1YK6vvLs9LdpYNh
iX68YbXXAtu1bmPKhBqjDSjicLji4o3a7BKUVZEmABbXxVqdh3MlHMDr455XviQD
u/iYEG1xEP3btIl5cXSPTqxHtgOJswtdzbangJ9PFpgSOhi3pjPQLYURuQYnh+5w
Q4ozx2btuy7szpvSUVZhfkMuOQxtG6X8e+wgFGkzwfbdLyvxtq6cQzGWLbW5/7br
7PdaaBvCUjmqHuCwwA9lEPsL0cytQKLxOZzdZpnbJuYC48QdCjKgDrJIid9886OB
ZidqgvLDVBEHM84IwEpALtNUiJgMtPmmeluXAKR7LVKFeWPHcrKvF7EWnlwdIngP
GUyKDIUZfj6nSvIrr4r27sO9bIruuC4v412CP6NXhuFELx7yLj3POuqjyBBSzv2N
LK40YIEywvvDRp44UDGFXA6YoqVAfQqGYBaIhe0Ty8GCDYOWbaVhHqSjghvtTl6y
HzW2ZPW6ddTcTeMC8+PKdKDLKDMOUlgGV6q9P3sgDZXkYjQJNEYWcIGclN8a235s
Z65ua9b4Anpt57XvNN+VhuzFKDaLqGdz3HV5Qz9NqlCCrfIvJ0cIQ9fAnwa/7FxM
KuAnlv+vZ02iRb247Z7uK2yx3zUYMmxTfBD4d/pNTjIg8ZWwS7JXJcwRgrI74FXg
HkpYgF39zxEzuX+zmF2gCRRhBenzLJyHqkwYTBUm9s7IaWOyIfj2GhVnBausxrt9
kQswXbX74YueakUZuZ+vSDk6VEFrcg4N2Q63PvZ+O3R0zfdjxIeFoPeysYGVSTIY
`protect end_protected