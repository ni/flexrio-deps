`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5744 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTA/AOCNY2uhRA+k6YI0pBYL3Lu1ov/T7WuCLarL4mA3h
cjOEbLV9zw4F74GcU/iuV3w0uzCzD3aXUCI/knJ8FQiPkp/snoYq1mMr8hI6uoMR
T0YUuEhAWAEno3eQGsDzXIMHJPc//hpB0x5P46NeIyS9Q4TrFojZ4+UT/rZpnRHA
fPRtZwcZAQTWEq7sP9teVcDOIl4Hj//8aQNQLczETOGwB4x/4hcbfbQJf1HQLUV1
u+FlA75x+C57hUkPaFtCRwCkYfnY0vHiaSnM6r3fAKFZm3nTH9b57LEatbBQ5EM+
645iTtG3og3dujBB7WJ+R/aRYt9lfuFONdC53EqNdWlTC37eQOVObXIYjXsHesUg
TSKAskcnENQc/JDjb7ev4Htb2GL2Il/Fwdugyg4P3sdXqgeZwPo3hCkeWhHPmV8f
2dYig2RNl/lwbVeWLTsf0cZOCAFDwUPiydKCh7n1GjbfndFuDAqX7587vbVWKQEV
wqxrvUNzZMx7/Nkwn/W9LR9uPr/rQGFIRYD6U6fCrMM3hFtexdzrFbWhPadZTqxY
M36DEHFHKQPkpKWD/ICrmx2arZgwFhGFU+n5Y8ckz6fsvvjSR9ZOtQBapZfKPQkn
0dOFpw8/JfZA3Y9lKz6LHfJewookDOeXgnUf8Zmt5Ouys9fqJkM6GpBZiu6KNERG
RAe3DJW3M//9XYoy/ZrU67pfmz8PdjtBgJat3IwixsjCT8cf6ZKNCEiHu+lrYndB
c80unIzYYdsIsjzMDD/1vQyYtk90tdWJB59czNAkvqA0F81cFekwB5yFAAaPv2yK
tiDZfSs6DvfdmeKgsgwZ5K1bPqigx1sfCMY3N8A7JfQc+ID8qar0qES0Wdd/PgZx
NJhPRrAQlYb2sNbfof0bwDBIuRDIp+2V2t/DViouGicQPek7IQ9DPCstmwhP7obp
1hQB+q67PO4zL8dT3hF41ODAr0Oy0a+LEyKUVrVqyRmSz0A5Pe0KdmnaPXw7Ks/N
BB7C+j63RegWKo3bMOr09jRSiQZy18dq8Uun10WimaX5KbpPocE1Cyd9I+P9bz2D
vqUp1V0pxdPRspsG8S0KGnul0dsMW7nKM/l5zKbEAdYT7WGn0Nsa8PdqD4dKRcNJ
chwrs1nhDtmk6mMi2W8RH1WWZ169yxdvaB9jd9nH+zFikZU3gBgKWghCNyk5iLZZ
8cfo/ImTdrFmrGMiX8Pn2LPW8DI3GAw5h5edc45DlY6TjpBOiRTewQKMfEU6QmMT
RKh9jWgs3Rnlvjx3QIKYoAu3ziLSa1YjMwVpyv04h1J3eYWD8j8Pg3L0qSO2PtL4
gafP7mxbB2aN7DWwH29fDjZ6cFVYTJ9P8lPu8p2fq5O5FnMwz/BsKcqal/1570j8
XCUOcRpO0HD7ux2OfXSQVNdcttcQMSQTOU+qEab899WFPBhTllVqe7qwCby5BPfE
mYyrnBEikjTBHsHLGeGa9xyprv1fJr5yKfS1F3FvfAQ9Ju2yXeOOPALuPgWr1bgE
7iZWwrmYEBwq0CUBOd94D73uBsbbjyDQU3//9e4kIkswWGIChmecDJfNkZSB9/Oh
eBLV2foUCybbvk5eEjQDjJ4ygoU3qaRrp7R/Vx1BPMRlnSpMAPn3vm0IGGcdL3I+
WM7nH4JanlZDYcNhaKELdgmpCIlMsNSWv2iPSMnd4RmcQsHGKj61MpwTUEH8cAPA
nBUCRwJ5LTFcQnVBHQg/TWKBcqvgM1roSPIk1krZ4Nl7EqHrPxw8pEoQlUU/dO3s
s2r6IW7COakMRrLgGlx/Id4hQmtE/K31u0JpOlTTirSpOjph60jNIp3MMVS5ReWS
d25Nc2N74I4nZ7vgVzH++FWnqrgEajvoITEsDw2ferH8IVX+Y++cVb1lyjRUk/f0
1Z6jCVGYg8qwvycXEGBcoBe6zOdP4GEyqqS2iArOGTwu7nFt7+rbT3EQZkCKAufL
J2Z88EBG0sK2Bf44jTesqyEY3S9mk3MfCgeEWp0EUPzlD4AwY6nucnQTjLnjOriH
zkwnEGwlc/6hEBEf2gARt5VBOyhFe0x7J27VETdb6GEccab6CZN/DD7mwOSH7M9w
Vrynx0KDoSMpUZfRuPXkHUQr56Yy+Dkpk/PgCqWhdGXolohmmJnLIroT9q1zsfS5
T6NzPR4ulFr39NofrQZMGwvDNVTfhHi3mzEm2VCzueWCrCKVcvNcvJREz+7eIn+N
o8wYAwPa1pdBcEHheZOKdIfCA2neLdosJna0HFzOaOm3bjgRokYcZ129+D94wJSl
KwDO1DCPxyNNiYmTrAGoe5u2GR9bqTPVjugoULINJ4DpBAA2kkTUzyzTW7681/aB
KrwLO36DGLSOS0TGyy9VDK/K0uJrtX4DJRXOWqP00iAA0EfA7pNkOMifEsdttp/w
DauafhZP/JHkdbHxH0Hk87GbhCgQF8T8KUzNWKt2EO3DT25OuF84B501EAMsRUqC
eGzN4HPLcHSUN959qH9SRovp4dyYRRAChz3pXR8T0fSWCRPQ6oR0gvPEjGodmaei
OuCmtozc+1eFNc5FQy3O6rikq57leX3RHj3dPIdqqwAVhHasQsMNxu2S+Xw/5AsD
LDUZB9E9ZHBQTjjhuwVy5kvE/SXgr0Hsvq3jAp0S9MGzntI4GFP9wmYXRUHLvKoF
/kPXgMSst1NJvPL3Q9MkNnDqbH4U4byMM+6qtpSeht1qEWu6C6pzFGRVwI9eQUWf
06WGRg+ps1uFt9aTt3z+k85USMYvryMC5uac5+VaVLppsX6HZ0IrI6JiKpV7xkMj
j3pke3T8TNIzZ3kunnGVKO/BhidDZv42zvz1uV/q7P5B9Vc3tniL6TUbSmzkcYjA
G2sAdyPKUZIOIy4KJqfNWO06p+Cm0uqFljcsdXoNH9IUlQymbb6CTJwkpJlfuwD9
iBO5te+gUtGnb8akjuYvVWP9kq7OedvL3z4+K3O1dNCw/hu013QHPn8corLj9JBs
qxyI2hs3XqT8G1g8aYCLNicU+vrq1BKn9i/jIbGpVrns9pKAEf/N9MQ+/j+guqZb
G2T8KkC00eaC7tzbrVmLv7B5Ho/WeYMsC8NL6MCNkf1lHbdq5AQjPFKV2bse2ooM
bWgDccWle4nFp0tlo6Vd662FgxhZ5WPgoW4qpvPDIVaFsDm5G6e8QZ5rHmaLWO2d
06geuJYvgANwrdFx2RM9VIzwm1ufu1+k6OhJpTfYnjFpWnbUKlV5Tx83QdJyckSF
bbuDRE+Xa9hwsAlgUnj1UaoO0T5KsYbu75LCKy/SU1K/M24bDmu9ypDVgJg+EZhh
SLJbyB7gNpNkI/epfFlhDXmYdVqEf4rLGsNq5R96pfjLZ0ufbpFwTmNHk7UAsjD3
vLMLLP2KGdkrpV2/PDISeH9bidAQ+SFLthYhOcqJPAixkAhE4GrKFK2nyp2AUgGr
OxcccDksaEVMGqOsphAqZNoWRBzyiLMcQ1x8vKbJ/daTIuKXIOMhxqAig9Zc7DEz
eXqYuaJXf0P8qpYr3lwwCdZ+mUMQnm8zI1gSnsCsqtjaBa1qXWR4KT5iauJ9puKY
OPu8akCrDCq7D9biNb334qPiy1wDVMU+ft7jbvuIJjbL57Wcw4BfrwjsOrkR6Qsn
7cAqEbq//60Ne3x+kskpd+dsUB2qISUtTSN67WEAaegJXXL7xEW6C/X7141/uKjs
dyu80TbPDxpIOwZ0d9G92+zfFpdSO8DVtbOHv2M4RFCgHu/XWyJYFJKxY4WvfLoK
6qTu+Expx6aAUzwv5lrcRY5J+6RpxTi3RyJSP/5mCJ569w3/oNzTV7fyJKxTRQzk
m7SnvxLYryiRMoVaLYdCEqDfDp3KuaFbCabR3FnJZXaF9AIgXCIuvcchqaX6lE3A
KDKbdB3BUrpVeHsFNBSrTFmQ9z9D977QqfRKjtD6oBOs5dyGLQrG/TDGoUfqxEfr
/V5RsvdUNv564MQaPFZcfo+DEjxTcDRJlmKvilL9BGPErqGxjTP76aAQQIyrEhrM
V+4Qbo/pFluOmjTs94MY7ynsdcS2lSevpo0oHpAnC1diORhgPCIUrUUFlXGL4Hbt
U3JY3JPNffWspdPC5+/z0lcw95D2VmpzAcg00rjpU/oMKOoOnV7NAetz8GkEBmRm
JyEJtjwmYKnZ/EQBJNJNOxLG6/gpVqkQC3XrAQAVBd1586qlXCA8w86UEyGAUD3/
iwOfKGewk3WQiCQMu/i20qut+OdpRdHuZtFhF2SfR296J3J0x4+d4t5H8psATmVF
nwRjP4pKS6h8457iSMV58CkZJP4/OLon0MXopKPv16ZYJxb2tg6nVdfUdRyfqyLK
e/lE+HuRu/5+Tzo/n9n3m5yveOzDbmcdd2OEM2ToDYYMuHvtsdTrvSAvmuXw91nD
EbhQSgBdnolIVOf3QB56NGT6FOv3Qv5hcmwuLno6J/KylI9c5mXXzJJPWbJfhJDq
4G3tTP+tL6GmNG3dRY7mnlFQTBMy8sJYk3qwWY7AleLevAyOdWk17wb/it+Em+qj
AQcDBm+0E8DAeRUtqsWvxmd/jDrem4awzsMNEYNEJ1Us9i59oA8IN0hQ/Y/O4440
3AsgdThAEccYDIveX2HLYBdMkK42vljAcZUQLpQYMHq7B/TfDcaPMo9RvIpUAJmm
4Y1AYHNMnxCji3nInBqmLNEeTWzc+wd02np6Nef7/JVB2UEJEEkulbK13TIv5FD7
X/v2dhU/ck61+M3SNtc4Z6cIM9G139LU4z/7qXt6xNrtkEQiPaBKVy9vUASlPPaC
KgId+ieSL1E45bVrKrS9m8ztKqgT35Vwha9sMwog5lVId6sKnpEj7IwYwrA4g1s3
yQJElJ3n4vPO+A6WSd3GOwyqZ8T6OuuFcwrMnKh0MpV1fIptaV6g3mQLNPeBsjdl
UwopKVWmaVkVWvO5lcYiobYBh8edL6RkEIqbpWlU4USrl5FJPEbCdlbT6BS+eEsB
heASwQbvq4ToDTVtnwTHPV20mh/fgBgB+6GS64nIdeNZHdZYAXumTVOY1+aaWOUS
58UQ8a/p6iOQFauVMVNhGf0+U3O44MBQpttuONs9SREc0YwemoMhGKinxXoSiPCj
gUGCLwNzd3V/l6caNGvw8qxrhjPl7kauR0eomr1kb4iFhkEhHqLhj+kiiTAhOevP
iv0Lwi01QCalzDXjCZobm+O+sHyxa0LKp4UhrX4yzeaiogne+Exd1stmF60/tmCp
bMyYSvS5zFe4jfs7oFhDWjAZVhMzCfv5vljwkXtqWWULfY/QEmjYNAGcU7q4cwV4
kcwTWxnM8B+T02mSf6iaZhZnV+rOJHq1vN86mrgW2U7Kn1xnCFcdzfuz7Ldt8GwT
SIR3GqzfrnwTQja6sxkVBmi4fuyDLREC8bq7RxNjTu2GDyiEA1kVsbnrMBmko91f
RpNlbQobMwIuaBXLHBbji51Xa33WNPXbAwcn5hwndBltZFFstGbL9215MFPjUPWa
T3nCqc6ykPM/fA7GB6Ec4/2esrTJNPPnxfDyc/EkNTDQwsh5qXeUvMeQqMFuMwlc
RShegS3mQO5FDQWCqKnad/58I7qtES33kcxSRrvJHTNi+fPDQy7FPRI+id9Ts0OA
D7ybeNj3ZZf2nD+mnFQaOTLqpr39aDjnhSESKNma2MKKNr87peoRL3U/up+B1x2F
iB2f53ofZNGi46LofAWrJi4AlZJGO++J5qY9r1mlLsza57AnDQ1FvSR6TWBlw30k
ZSeU1F+YvSXtkzTSD+nXzPCHt78JUWQPKWob/F5py2ndOWtGes73WBVAlddnTDb5
oRXz62n//whvJDiVrJ6kJLPEQpwF7WzkOepkISRTGoZgevuwQfwptN0itoG5Tths
+xYxzxHkPPV3mmONSUad6tlKhK68xQiaW/JNCJZDm0Iixq8mdjBXeelC8PbvkC2u
MNpqCUYXfL4fGyBAdPqQFarGZ81C10HvjjK+jXczrTfbMZeAV/FVgYmHwyOIrnx7
gCd/RrKovp/EwAp2Q80QO5b68V/yLZVVsJ7Kc5Xq8j46E6YiP505920vVhbWvmvg
Z6J2mN8r2KdjGl8RhtSp2w9xoPcaV+4V4wmBlxcqo1IHJ2lSsIxxNcRCsRDCo/q4
tgk3ZnxQ5w/NjbhTEVYhUhzlfCQ9Vb+FmTv7Oml46uaoVSFRcQikuNHUr9g8OrCp
Hdj5d+bkTs4x5G9k0dTw/8L7DDWHdO5wytnzdVG5gQn/B6/tpDDhqOaFNHOkgk4N
2Y5fy4nG7aiBMA/vGK9OtSJ7yr2RRswfa8HH/NV3zfHmI1PMs7Ex9KQzbWNyBEa8
ppgQHHWe4qZ63YTvtGMaWg2oaDUygJJ4B3xlOBYP0qXj/FZqYNywdVVb2A1X4kLA
9msokwpkI/L1E8g3Ykxar6cBQIxb0jrQEyx/P0jgDNlvkUaJehs1Xyqel5N2eTD5
DVDqY/khcpyZ11TJXncNltudk6vqy4vBetOg5yKhY0XynArR+FtEV1TX0fvOqbOZ
fqGRnuHwTp7G0YTl2XS+Inf4Uz2XRRgLWBrBrHXtp33474TMocDinnsDzLKz86eU
4sv8nXjUjFI6sXzAfDdbrF+pOiy9LYAB9sOhGct1cWUJooNbTgPmkTazzzcTjQFB
Xw9YA/3IuAUVg32ljCLKGpXNm2w5FTXzwgB/3qDczWbMTUuzFuFBZrB2R3/yBhox
ZoL6CSvq8pFLN0f6DusodR1/NX8sv2fzqeKCkHf0yQ+NmAKrndKcYFEqiDE9YvaU
OCGdEt7q68w9YzDixKF5X1ZaTrQs3HF2xnwUKq8dcvzyHDiXkOLmicOaj8t9TF5E
tsZ8ld0gjHhrqsdHEMzzG8wuNyFcJJspDAEuVvFs/T+2qUiaRe7RoDEBJ315eM59
H0aug3Gk5vtRVGcFgNlRuvQ5jQPdg2Vw/0kYR2Ss7fkJPBTlXqiSDhR8nXuf0OQt
V0I5yc4sG52b0wk+qfeH7FNhi+6NzXIJaGzMUM+fTtlEIu7UmS86srGb6gGgEOYQ
loNlEjvyrx3BQ94NR4ckDNNLrLpndfCtr3skDT1DNVqKNoIl4B69c47jerS236vc
xMOjkoTIoVeDyZ3dlc/zgpwmDacpMJV0D8P2a0TN8oKwzadfV9sY0pY4NJpVfMqY
Vas2haFhE6RyAt8o/awNDYo38PmC1ekXk5HfU2UiuC1rdZANsmP4m8tIKD5Rq7ur
kOPMrVpQniced6Ksjphj3qVfDRxRausws39PCajye1fo2LgrOy1yrdlgjTQzqMLF
cNYe+77pJLnqxzFnttBmVz6UBy+K1OM76p5dxe7uHL9gE8p7lEL7EvWD9V7rLlA+
bry+lhCaBwnJr2SwnjwWSmskClheXsZFhoKdHDeO6sB9E378oNCdC2U+GCiLzZl4
D6ePpFaV6FRynflBOtf6BwnA12/fHKTfWJuM/XVHH4KTo4MGLME4LoYEhdWKDlvT
yu27lRFMmxCHy3kumyy2WF9QQgV6B6p5KHKL0WzJJq8=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5744 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
lmOQgIOM5jiJrGbWpsW/8lbD8Py7oomdr/mNjPh/srU6WVVjB9OMYdVMwjpx80uq
zUlmHVxyeL14/dnf6+SBA7eIqI4WfhHGLAhGWRXZU8OdXlIv7tP1RDRx0qhlLkwt
Wt5/rdmD0+gRYX5bEWIrn0q9Dl0QLTO3/NsKBlkAS5HbrvFzO1JR8qz78sF+XebR
heluRZAkMHjvypWkGevi9rGAqHHhY7pjL9DlFP/dgXR71iEUYJZ5B4n3HXanZPv+
REmlQkYELXxtqBuuqIC+0crjYz6fW0XNsKzYMr5c0n0n+oQydg8yDtQXIt8lFd7U
gF9xU0SK+/l+R1ERqMh1KV0j0xppYVxKDs49NkDtWF81OOf+JUixssjwoA6KU4ea
Mg6umyQmGSTADFAjaBP5IpwN8NSPRS/TXF1NBIac3lQt0ILtKsl1Th0NzgUWn6Kw
q+hs7tflLZnSYVgf78JFP/4uzSYo+w2XHmJSU984aCpZ86yED5jhLBX1QQDQcw/K
fhFEK/gFeRRfooQj/LSCeiz7FsXdptxb/6XjOXES99/8UCWs0FLmrjcLT4DvUTJg
7WMkqJ0vDCjFMzpJ5sFs6z6bAckpFrJCJGeuitkD4JlHhh2Eft4CsWfJpNNwxzgl
vsGf6zxCxVmlWHE4xje7ZXQZSP229xKsYuHoVMZ2o/qMLh7whlVN7I6YQFo2Cm7H
PlghlA5O1R3ZbPn9l/ai6zc+g7hgAGhk3D7kzHQWFBGqnY1bRFYQqHaCEnA0e2w5
d4aEagrUy5nVo0RFki+ORzmEBS8j01WCT/unwIRxWqPQ1DjkTJnD9fOJ/Utn1Kap
a6NjQldrV9b0elTqAMY3ktUA5umYxo4jIsC41YYh4JE9ohi4ffqoe7NGQQ5hBi6p
6vWnaQZPwNIb3w5dfWsHpV68RJazb9pD1HAnpalkzMsbsthapkb9T6X5UqJuASLo
2oVIrhFwgZiA1MiBzQk1Y9OirHtiyyo62T8uKRFomNQP50qePoRL4NE4jyxsE/cE
AuTCI5k7hddY/zWX0FqFZsxINX+P3Ku6DIKrMeC8Qa3L4k/rkv3Cg1UxTgp/y4XZ
TErrPFDClsdQvoNGVTtzU8rQOG9z2/R433DNXnTJ5fDZU0EZhREjxnmtvLQrmfsL
nrOEQz8oJprEkOEuD6a5vZgIYknR9ymVLG0+gQuVyBU5hF8yP3vKOSt9bjeY6MXI
cYWofgU/EqjXsuDdv8KR0wKJtFmIypFnFZzDtF7sL8/Ggb2/B1nnmQApkn606P0r
7XMkWdbH918nzXYnYc20FQKJeiQrPjQP1+N5CynNQt8jDeRG5DTKpb6pMTmksdE4
PjIOR8UHUbGhJl9FiZe5/0htgD6ara/NX5oHyAg3KAvOCgwizkjFvsTNhThtrKBL
Wr3Pzz0ckySxbzAedR7+/e/uOEV4szyRakRn56pBH7VGjpu+BWOhDw3rLSq27mon
Nk6oGv+D7tcXTd6VaJ99hWAg+w367FWX2UOGLChfjAwrrNCndoASTZcWCq/XIxhH
LffwddFrZDwrvbmyTYZLHwtYYFC0ZDZmg3Akvsidg4YNrwY40SiniEFy1kwmvbY5
ScfNqol5MTCTkImvA35a/bK+tAIk4LYEAwkR1UHmbc4RPevdLDRJ/NIlWClJ0Z7T
VFdyGD+Nsj4XAY2tX+pub43LsrKf9q4wdA/4xFlaZs3HiG2ZV3szyhC/TusovK8W
L1WnHi0Dj+Kz96RPv6hX6VToL9wlvp1txOnSXvOVb6iXyygBybXMu7ybTlweY/AR
b3j3MGUMML9kku0q2EbeA2bqOZ55dlTfExBAZHwUtd5ahESWwNj5WMmMKZLL3lZz
qK+F8cZJoDzMCGA2SDrmDVWGil0yA4Mv/N8NGnIn5YWePjOZlXQyYQTSeVDEWMl6
xmY/BVJtT9nGGE5v5pmyIwIzbmKwzCpz1mRl3DunA0EbAMbztO9erUn4oRgZVJUm
UOhBdsXzO4zvFFNiqV5pUQI+VDymVgOfzzbvhmGDazoLwThr9/SvtLRqxWsZZlNF
9TsSonEZX93FHERB2fMdD01G/ovYAdnAtNepWx+6vx9dwUbvvxUHgLoOIF4rsXpU
O4B9NGEm0IEWX/it+hsAii1BzNq0hSg/qMBfQWNdWIrrHBiFIMqEIL9ZwXu1oJkA
D3IAz/4rbSNhp4nVUamdl2RKkEmraDz7cLOz31qK5DQGf2Ed6n9yxuhcuNB5XDrh
YG6blVa1Y1AaSPKlZAV1AaGVHPzjuPvSeWQR+iNtW8Y3mrlDo7rTnU+WJMQ8ZsL5
X977KjBtIkV2fF64TC6QNFh5Gc5QIG0Fj28rwfTqbZwnxJ5jEplCvgoqjC0IfzLT
ofbKd9cu0vTegUn8T58AwfzD6bSR1u2GHXz4PA4qYSZykd3koTzyHbuAsCUjUC06
ttdvnOJbI3Sl8uHsNjpvbsnOVnkk9N66GsE4spcofukG7j/f/znaoz/TfuPTk327
WRYMQVceRarcM7gQ+ju3JK5G1l4UmnXdPoaj7J+gktMXzCQnCCPtlxB44gzLxDL4
bUkhEooRHvNbHzpq2P4+4dJO9fC83SNyGiPQSPdwdAXoHLaVUfI1wHRShL/FiayB
1bGZhvWZTcfsJcv+9i5XS5nx6AceUlid9nesyEW0CvyXhrfcWbwgjsP+AVhi4O4Q
J5RYrhFJktZb0oO0Iz4cnmv1WwjxVgyua/lqozFDUSW/dEhCxB7zw2ddWYVg/Wk7
0nOHrfdgEA/yByoOt7lbq1Jj9jiwJZZeS3oRnAf6GVIA7IRxVNO2ajYeZ9DD+jTJ
iORa1T2ZXfZV/yQ4xplZKYSVMS8/STSTptcUGBskUNdtYuNvOzR62xCTzGKzbqhV
g1nRuOdNhBanTrsb55Ewru4dM/oC5d+r14EjgNywZ0w0IAC0AvLMn6R4OnHBdsxV
cC/OLITty2EjtbeQak+HZll1mLVTuWE7GwC68vtRs0B77VnYbGL9KILbbLSHnL8X
BgFEacDdyuewK+k9xHHPvUnYfs5Xwul9osB1HsQ9Qa2j7xghVYj7QSw8Mjm8yORF
9DIaJ9OZh5kZc9OoTjkikR/wz7WgdcfyRC9Gq0YnR02yQfPRjyW2PCUgjTlf16eN
uNHd0WzfH49qQVp1VjCI8hCcp5h42RLJCrBe9lGidFRptEcXgR5HiZinHlXF03Gc
KRY6G7KDqbGmLWLB6zERvS6MrBSX8KUo8WQhnQ21Iw7CZnFQVY3rtJuglybA+8Sm
n4OrFDN5mUtZf9tXhxc6ZzRhM/+6mKuv3ZC3Gaw4kE1Gki3bs+SgkV18LwICmRja
gXxOliSG9nEmixAoVYX7SxIx26h9kpk04BMJWpgU5xSbqaZYJN9FiIcaOMAx7lJL
RKTLxH5hqT+RJXEd6pyI1/JaEg14ciHXO8X2VlnJkiUVTUfozjBpV4vNmVV/eVp4
VboObRH9GrS/SzOLNSuPX/8OLbA9Wt1KcckWs/pklXtHQT2fd5m7pyeXcjOBOiQX
+Y2dIJOU46WHrvXWJ4QQnl2BBuc+EJuUH92TTcDfKjMZ3p53nisEtlefJMVIoW5Z
lgJmVgBiWRhMQb0FXHYQytqfVMB9nfIm+n6YpI3FY7wKtggciCieh9lCFJE4pZnw
2vj4gN+WOw7PXpiDPjN9CXRVm23oQazimwJ+0FoRJqMwHb1pCAmz1WAjAk2LmRVB
2hRK+lT9A1MjP5bPOrX9P1VAa9r1abpqxTEFZSfwoJHF8p516upbJc6dkWEmlZqO
zxtHC4D9vnoz2vGNvuEIDUcOdyvmvTp3ORfTPJbkwaYedM8UVQcYSTQKgtt5KeF3
hYfRfVfu86b0mVOzlOF5xg9HUNwwILhXkeEbCKPmWF4yvM84LvQIMQDCjfvbTT/a
zrKOQNTWmAdpaaE6gw8pTjciXrHenF0dACk+Vz2YTTUSl+ZvXwc8QIQqUAceaHsd
9hPt8FZE3nAiJxfnzJeavB9CW9v253Lp46nHTQQsUgmfX+9iFyIY0rfuSlDCatIK
77wI0P69UJU7nVT2xIOT7nfIOszF2FHIkPqQ2D8tnwZsu99qvnfyx3z9UFw3NXsJ
wX/rukMBopLkFL2kA9BYsklNGOdQrT2RwjxuUWZVOga7z6DXiEeM9JZovbYb3gnU
4RVA2PL/F5UCT94BKP5xxFsXa50Fm+3aJeVUSBWLt+d/3RoUgwOIvDg1ogAlGrXT
PiFSzDkCgHOzCOUvcxYWhtCLvhm9QtZiXOPJblr0alDPUgjFKjdfDMU06aTqreHm
zIwl73XxcBhmbE+Azo/p5z9NJWopahVUeFrVrvDIXM2RBnEBQ2gK+ivFYvc6+NzA
2Deiy3Hdub/QAfVjTVKZHPD3P6kebIR9FBZ+NvVcBi1phr/BkiF5Z5H5sge8aee1
ke49YdT3zbeT7pmaZ8+qyY/YW/p8MPgUqdhca0dTXdyuNmAQfWmCsJx/FLeqrzvt
DzIUirmbbO9Wq3Gsw4W4r0fXg5b20YjUhZaGbu5nZG0ZNQ00/XG/foLBP9KbfpXy
Jyuc3wRvnROV1UvftSKNNRQEE8o/YgM8pLT21CpE8LrqIExguyLcWk7AmsWKTSmH
YMXfsUiHFNxc07WkiQZk3/hHzhM6DeAbkwBMom4cO6LurhGhlO4C7vSj0uk5xy4v
VckA89C/PszWaKjxGEBhcy852eLKsdlrC8aMssp3Fl2M69kSWQ8YAVp4o9jFd7RH
ZdxOgm9yUTQ/s0Sdu9P8uBd2cYp6m/t9ADmELMrH2GnyWWJsUBovLrEE/W/0iej/
e4oGv0xmV3QV3d0vKv4FVonIU2yviHqZVfWLk1qthclA4799M1JVAH5XlqyIlkPY
QrXmfuIjltjHIMvgV2Blo8Z0Uhd3uihmv3+ZVMQcfUPVg470MGD1w3KXtwdfo74Q
u7KS+OCikwPM5LvdcBfDiHnlPO86Mrp//15tcw8QE/a5mveOBIDusPrWqDVQUvTN
jMqMY7cOjrwuThaLRdHq71p3OGoX92Hj6rS9ZKwrn0/F91c/UH9kfy9oWWvf0iwP
JG2PjZCAAQLZnocRg77aGmcPo3anKd7tZwxum9CaYi/ujfW06tDkVI+hlawGlqBj
IlIWSDUl4zQzBgSVoVwMOZoCiZpw13sVsv910aofgJPc2aI/qforXkrRlUCNzdTd
T82k3jFkRIu8vUQjVU/hwDb1F9ifbgJIK/m64CvFAujKb2xpHq8LsajLVw3QUD8J
lm8JrDgFPjfEdJD3/CvNfW7c8vpmSnjceuEjHf95INajstHVu3JNmnePBDEESWzJ
F9daQWkNLC9scV2jB38U06qOtH5C6yRSfvVktbzz2KLvGglghVp3xaJ36OiTUGH+
9yiIlbCrH2eYyBMOHK7uNiV0BwlPyhWOVu8BPqA4iSg9d3Zv6JmW9COQxdz8RNfL
LsBXPx2x/+XqBZ9gnG4J56VBsLnW3JwB1nGzPF7U7+AgFL71sxmE0biLc8kXOAlQ
oLPXITO+0OcAoHu3d+oQ8F444V+YIeKtWuIGr9KxZeCUSyBbUNRcFz8xhm+/z/e/
/fpnvdSKAJq5w0bGR5J+6Jr2L7Q/F7WAIXq2Hr9UxWdMZYh+U/1gq65YCGk8ZJMN
f4XaT9+PQGDwPFwdYq/olXNN8wmmEgqMy5hiQUhyJWLHyg2nk1lJ4AY8M63Ivofp
2E9673IdCEj3nQyQVYbHBCAmEUsdRo0CZ7JCqaEfwska3JoTpUYwGngRgfHL6jc3
lYcynV3VbCNG4aR3Xxlz2Pqm4CmVajnCYiglafyO4BQjoCh5OSyzPNI5y+24HiL1
/Rlx9vx/gZ0CCWdRGs7pnfoysvNNiDScuUP5MHFF3oyB/9tU2hmbHulm8t/ciIll
n3uTn3Zujv1LDLyi4/t87cFkI5R+u7hWI4yVfbrtg0tkzG0qzIDM8yxY/ELhebEU
OUB8toEexP63uYvSj7nL6MecoQKUna+PHwGRzFE1LqWi4vITi4Pv7grc0qcwuy9l
LlXq6jldns5j31Y7eCCXLSYBFhOUbW+emwL59S6QsST5C8qr58haYfmIANFwu28v
E8Pl2ghH90ABLcuoalwLJHRlHCBet7q9JVtajjbdaTkJ3fHSiqNhLXiNMDp8qhQm
IKB8Hn1Yeo2MDKn7fiTJTBxhfWZOEPDhnIw0n4o9LqbZ/lix7zZRRn1Ezj7Jrm6a
C2jNcV7cLV5RlxaQNuAG55NuNIpw/v6EkwFkJ1EbnkByCYl/jablT+V3Vb4LZL0p
1vxHz24W7VMg4DwvwHg/0ZO4xFCyHyWbja5tlURL8D1RS8fS+oWKRhaeKsd5inOv
jCWISo+m4V3IA99BP64dSN3Rs++K2jnIIGtICE2aCJvYYeX2Z2YNdyxu2X8pwnvB
MQZ6Uh7zXNRrI+P3IiRZKzH5rvh2aGv/OqeXy94MGYskgEHmkeDUAKcql7yW1aNk
otF3ifX4n2HwbCxxptst7ymykw+5JeSz4BZKhTz/yiBNLBqMTL6y2Fjz+E05zD/r
wkYCVKKJD+AEYnKCQslJsTtXmzcMdCrOOQwOmp+xIgvSXnnwvnie32GFaFfIyKzv
8EtDvxkdUONJiP/RcZfAwdBFRqhuRXuAtPbrbofUiKVHeKBJS+WPNPkebESWEo0H
sKVKLicUjhP59gNpQHwnYbGTjAKVFYirqLu9hBNFh9/BUOFweIvoeZGQzP50+xb7
QmAhkBCrlEFonLc+5KHADASSj8DAhyQli0INX6DhBwjw+nvIIEnUgozBQWQyIUGQ
Fw6Mt7tHomIC6mELaTOdaAT3KUWzkUTpTNHUYfL9ZG3EGiddBHcHtxnFJPYp7CKv
2aYSt2B9Ch+DaB4sPSt2b5z4n97bWTKGLE7mRpXwjq46oeMDIv7Fuxy86qgkyP4Y
KK3PB3N22FSO+iqELMD2LAlKOcCOXqcVzAvzPHZ+3GHidLAZyH9PIXMZ5o8CCgu5
BWmHTnqo2l8llR1Sf1DJEqyoSWjnsarDCd7jKE26sxY7Uk7FUzf4D+pR2JI8LE7l
LDNeQ70ePXl56aXZ8WY5jBoBU+CIrtpcZysykv2mkjWiT0JnYcdaD3AGNWFGgaHW
ETzTxNE5gFGIg5KlYSJBrO9LxgKq7qP2sGUwZaNPaT4Wx0LwgsjLDcL+MzNvfh22
rYKjOn9yzNHXMPK/+QD3FjikXS+E2QGeWvTLw+Np81NQlkbHFctzVDRX3wjIxJBK
pIQ+SPjmI4pkS2VDjrcYiW+a0Px/gnkwgjT1vQmCL2uB7Z6cUeJuoDYlSVK1jZ4X
3BT/GPBGt9Ef80p+kvXw+Yf3WPO8V7tL57tVMKWdxXTH1kMyr/+Vzobz0TP1LWO7
4kZkMoBsr00PUy4Mx9S/c4noo1ydXNny/Kyz6QKMByZeH/4S6IQIGKJKVuYkBDtA
Gdj0khCiYZKTEFrPOZ8ne/pPDh5vq5sy4ptUUzzyabNJyIHdyTg307wDRhYD/xa6
7EG4tPW+pEN+VOw1gd6HHhkU4AJEvFn/kSnfAMllme0=
>>>>>>> main
`protect end_protected