`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aMReDmrPskJscpWYThVKVItA5gecPPZO1R595p0GoIq1TSTG+UxXhmmUXc+VYHJ3
u/C3EW5qePLufxmXxmhmDnr9U8/cYC1zLfk44v/2OPb1TBrTsludEDQZdGNWeV9l
cPUMSIfZ0dHXN7L1M1E2XtgoTWQxf3VDHs7B7lU2y9Rdm/ibz0fWMow7op2nWdD8
gJ4QlNl3f9Oiotp1p8vz9RFzzZOF5gBBslZxcTF5+z4qO2W7+xLByngthWm+exIr
3Pzy8qyUo/m2DDwOz3VJSvSNm7RUq+0/yJNOOz3jr3j7ZyCj5OqT/jDAWjJSMH+i
2402Un+wDMOQxi21JLo3cA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="5R6K2aWI3OdbT2A+sz4o9+2XAInTqB1/cSw5W16RnA4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
Gm/2BIZF5/H5qen8uQizPH9RftTuEE9mgEOF0SqeOKegtP64CfvEUnIxj/ahmIpA
6xUR2v2l7E5duaLZh39Mc1GYsfqE91NCPU5whLaBPg0UuX4cgTkO4cYbW/7yvcrd
4wavUfwXEp2VSiN7EVxL8RcZTSMSI0Jr/aojiilFqVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="TEmQtJ1Dsm7TOzpJk/CeTSSFx/zKExk04H6I8sT4Meg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2688 )
`protect data_block
nvPqn26PC4XWLLQG0Fq8XsMTlhB4evbpiwGjZroFFLgtNlE6bBjdtwWsB89WW4j7
jNfYbKN4sBv0hDeMH0AAR+8g+TCqoX7yLdIUd7aGwBUZJr6FdDs2wTUxRkXFYNTL
s0g6+xYdoL8wZliYWMoLx7GJ8bAe3/UR2L3GAMbsON5VCcQtw5ZvvzuBf6TdTMVT
E96gLecYRDXV3lTjlKnd4DKWvRZyUuViwajQ2RGZ4XMbnTMmBXuhuFm8lN234DBR
1eeYQV0MOQnIKjjVhrgjWFIe3rnkXrbPwl3QH5GRGlw+xVmBy04TEqI6BQ39epD4
KGcgCL2dl/LQArJP3lRX8zhMRMkGlKEESiI+vHd0hl3gy72QUfswpUKZSmd+YXnH
2Veri3zgjVKf3/DrzDnLQXdQCj0X2XtyvQTg1WNim5FJvcpRPrIbC4ewQDpVpwX5
2yC0L/cRz6MmAL7j8ljzwoxcOKudJerUegj7FKejsHFTwx5DCa/H4B1DY46IFCR9
W76WwBkT+2Zkc6W3aKmr6MhhvFpczRL1PXhKSR0gD/kQ4wf2Ji06p5tA4rdpi+7v
EsTe31A4EmVkMWbaCjiwJv7FcnMXKcHMuAGnMaod4S1WQ1zLyuV1e2mwaM2eOk4/
bSF4nGJtUjOWT/emY3QYC8NnO/gxqXfvihFDzoLcmCaYmfJNTdyB4dpNkxtERd8m
XlPoJPbnm3b0Asa99HNQ7Gnh1skZpcv75gJvKUEO2KBXZ2GBOmzxIzez1CT/AVL7
D6EaRHwjtQm+8j48HsXPuK+qFWVNWXsW4cBXnB7yC4gGFM4d24AsyZ150QGyVZqa
VIxZeZ8FTrG06+QelH6m7uNOivwBKx992UR67qU/sFfhPAR6MomHxgeaiKMB7IYn
/sx2B8YxlKU0hQH3j+FSfP1ck9q5JGPrcMn7qq71u+Bk7Jck30KUfs+rJRuzLWRn
fL5pJVRvf4wn8eD35vGcSc6eBVCUK6o74ahJxz73fz51jHwSL64o0M1xYVu6U/W4
nsRUxJpadnTq6VrEGdaXGF36IEXM5KBQx2S0u+qmgZaTatYHJg4XBOmlCE064IzD
pZHErMhuFoDfAw45utKIrEoXDwNLiSdv1HHNoi1ExqfBy6kFJxXow0AW/GV292rE
rVm7ttPtePNpOIXTR2nK1FYLdFVZvg2I5RzclTjS7NhW3nNq/ZWl0VtZQGQF2STt
SlAWH2tv/SENaBlu9/QaJQUT2C+CKcx9pxPrXr2HJEHkw/lu1ZUNB/yvStCnni2a
2n5Yzt28vFMhprFluSYij6gtBTks+1pKYecouzHspEBptjunl25M/WgKwRIWoBa9
6BtFyqOzSvc1t115h/OYpVCZcXold1nPzIdclQZoTXhhD0JVbVhefr8J2MysIQju
Ici3oRC3ocrUmuVVXAQLNY4lF728j6lstdyAeX01Ihwe5Q60x8eqB73PBdV6jHWx
hen9XkS7ouhZ6P8N81I1XeeCm+Y1MZtxw9XM9uivtOOGb+hv2B/edhaYRfGMmf5K
rFmBiFJvRmp9wzW1cNM7gvtHCiReu558tKnEMyRxYUdjh1cc5BiKIpCVAgkIjnNl
78po+oG185d/YxdcJI10TAslTH3pNkIwPyAevrqmbXIjvIocBi0DpJb0q49Jd6W6
vJeQQPNFhg1qj+QCG/Uy5k0DiTK91ljCLTNF3bCYJxnhdHdMlHKnN/BYl/NuSvto
wMIie0CAhNpaGZOexrj67gsRNE9kFn9zYHIRDlRdhuhUWGNbF1Htl9ykuUzUNQ1e
3NfrEdQyKlPzhVfZubygICUiYXcN/gUUScOsjTWHOoVtjn47kYitDgIbO1yytbAc
ghJGpCQ7C/ZQFkrDRmJuR9uLEii1/61+UhANMS+Dk7OUbgmgpZJa4P5VTPtCJ5Jf
Gd0Ytvu6AQ9FbIRhzubAD4fFXwcQ54OszkT2/u/Urjayk+4qIFpsBjRUoGFJ9wli
3M82amUmrH5tgQZaOKITSrVKNLy9OYCkZ8enQrNX/ZZK5+Uu+LNY6Vlii0ysHeLT
32LXZwA8p0EK6H4FMs3qLVt/gH/aflQwpPqEOF2pxr5fewElZ0joAmwoCeSyraHD
7BzXOWNonqSjPEB+2Um7hsvUvDKgAW+twNqupohUkVMKPrsKEiac4cMVOGKq9Hiz
rwfj+FtHKAjGoW5+ObTnKrptvFC67+mnVMF/0WId9qM5xErID0bOa+KPgdD1vk0q
4PoNzbowLMMc9DXOZ4l1nhMzzG8RMiFXgZB+QDjqni5PlM74wvrYYBe0o5V19ar9
8uehlWlhWPiOMrHyiBd2PeyFFIHY0iNvRPVs0n7xYa0N9us1wyvNRtoGfHp0l4Ye
rK97IvtLSB/UQwwJtpT+yB5rwOoQF15pjvMAQ7JIWANJokOiPmqGA+zPnIYEMCky
KjiiAg3ZCmfnEH2dOu8zAxBZ1dqMK/ZwOU1pQbMxB7TXUqg4qnxIc2uxHpdQYqOo
ghSU4cB/aW6JWTjId8mZrtZ+Tjf18WgdtfluErWlbgxxgh8C7zs+oN00Ki9tsawK
g38YSTV8v6jlNTYrqRfdQ4uULV+B87qWrWXAR8UUBgHHimLjl/vC62QeCSegJqMS
javodbg8lYCsLSQ7Tnd2jgSoWC2PHRyKCp+qSxm1O9Ln7vjBaSlIxlnEnAoj1Z/W
UkThmDa0VssPAWl/q3b7pjBGfvr15DWllxMv3h60C40rmkZTUO6KGhgRp7a/bMHF
1e+28A1yUrW/lMJ3lkhDS1Pk08znobC4njtwRRgUBOM9OXRRGYkKL3PG+Ra86LUm
IakCD3Wgpez9xj+x4a82YZ+OB2NFcg01kOBOzPP4A6WfQsbsaTsBGMee+zcDXdb4
b1uZzvq0Y+oDYVnaO0yfScv2PQgUka3J06nwmYklvKBYHziLF34W3zzswMhot2n9
giM5dBNbV3sEk6kharx3RW2Q5b/Ot83QXln1xyePZYUeIK5hy+vuULv7w+aUaydf
hVQJZR57YsxGd1xkZjuOWjW2aQlCjtcPMP7u4iPgxwWmoolr2Q5UghBTVXkbUILv
OsI48ZkIURzVHlOY9Zo+zvESs/qokR+OcaWDgEQWjquJhuEb9b/4lixigChlDjkT
oPr69wN1YGf8azOuc8Ag8ADhAd+vr2zQOriwBIOekH3fKMez2ntXsAPq8ivF/6O7
oMW0Q45tawpWMWe9ilGtiB6GDi4Ov8g62IFs6Fx7zVD9mfartgjXfkKMRUIjcb5D
8KRByBaHez+ErvXeiYTqmXJgt4DDVEMbm0d8M2Q0uecx3puVlOByc/se3RiyXqcQ
TPpA/6nxhgzS6thy+9s/2hgsuWSLN7GC4e5tbUF3sCRPiiLafEvykN6C/qTcC50T
WnnEfbmuo+jsCybH2OAj8g470eUtQQKuJDVtMmm+sKsf37PrfzXPGAgTA9i7jEql
C0aeto+j0uZvd7fUDGPnPk9SI2L1b8dTsdXDQ4xZ6rQzTTTQqIp6RLwxjn/f4ZsM
UUhC3xodeT50KBNda7uVBSMMzWrBUXuhfozXlHyE4g4n63VwMbUCueTkj0jx6oAH
`protect end_protected