`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14192 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRvp3o8+RItkxKTewZIo7szbhVt+X2UhePTL3ONuIIS6B
jS4QTIDES1AAvoCrVfQXjH/RAVW4q81cCPWznEhaUUNEa/sFuNrFRae0h7FffBzX
RUch+C5EskNektRcixlp39svVqE/rLFNHC+eCm9cPbUMIyMqtGqIX0OvfSF175Ko
HjF7yrXs/PQj8A5rLPW2FPKbB6GmQZk3M7FKncgi8DmAuDArhW07UeymrNYudH8T
6iQ2USvmovAP5/2F5XmTqqpxw59SS4NPSZz1+bDL7NnKWoibn60M7GT3j4A6sLyf
ZHzZQbRyTGPBbV4ELivNycviEvjmcht2xlXD5UuXh8P6UFZwmL8uIDAxvb9Xelj/
dbWYVRPOeT0uNzIVGqzoFZZ19NQCmzkjMA4u9YhRccXZEVeLOJk+3UdfOkmLqZKD
tjP7GDtk+w+mcvfH9ESDZpURuc/BW0waK8i9JD3gQ89V+Xc9oT4UNkNDNnWl+Xu0
qhjiXmeCv4ZwIgMUnj9gyGd1pUgbPCW0stU7cuoLcelFTD8jKMzYS20bNJBADaam
GWAnOh+PmlYsMuwcHRVC7oXbYX/S/JgcIan6JWUBTuW5SC2UqGCZjW3QW131qive
s1K/SsrEEwmVmnYBUuFIsEy0WgXKT+5MhdudDm+H25L/mvGtgmML6ck5dgSJIIhO
RbroVr4OUg8oTkF9VFXLvlo1kcbBmoHp4bJP35JfgSA6oO5z09ugnS/oaAfKRUy3
9EnAr/1hmFhA5KQAG1IeYna2NCukxbgdMom7/tF7ws68qIpYJtHXIvgJZN2YSI3j
YDHJ6ccoPOozJ21yT9ioAwKxvvze9jH0vVNZJu/UigVpBkk0h9obKzyyZften5aI
yLCSkk8oODYq0iotszfxmXYmPcloixEPzqEh1cJy1p+u+zppqpDZXKfIZet4/zLW
SiI67trpXdZGGBRSJR0gQUt5Ie5aUJqmrwJ4BEY64jyoefNvBSKo8jjoWYV/+h7N
lQQY56q0NCKnyKV0fsx++CCElJtjvyTZK9gNMoBIzTdzplFvKeZ3X8+a8XpQGjDG
ISrLZhlByTexfEW2BO0l38yfIfOh8poImhM0d79pJn0iDfWCq4DJ8n6yx52DBouz
QtVihXkzLhHtoBwW5RUfzVl9rGOy0JImZ1id0ZPR7a4/AuVue8hiux1Jm5VgdgPv
ZMrI8pQBkdY3xHUJNav+VfHeEYFHbaLju8SjiQMxq0ac/McqSVL1PrXDePIzGxvj
BQvX5FD1NGYI8myBYdCSa1v/Y18GwGvdxTYm03MToGB9iKVXHCksGcA1FWf6h38Z
c5RkG0v6HgT6Qvfc3QQB0GBds9ftBfdrYLv8gxokYMzYQ2adpEdoffLk5bdsshgi
+iXY2QlqgGT/WSJI8tAKZgFFG/ZgFG41WqRaNQRTxc2Ghh48LZDmJVgzn+Yn46Od
Es/gzZ3vU+HtXeQeV1N0XruJJ+/P9jDUHgP4MVDbVwIq3qRfEeDJ/9aRz23PqjKd
5dMc3ajf4V/+1JOrMv09FQlRyKqB1p7tGm1oz5av+ASbgQu8mCgLo8W8Q+YpUTh7
6uUz+R70y13IIIgn/rahAFdH2lw2qwfhwnUL7xGQJLAde/3A8X/ooJL2nKTWA2Qr
P6Mk42eHS9Opcq6Iu8insk40LFCq7ebMoCOMcZHTBGagMWAlus4ABIsR3WJulxqa
OQql2YhHgxLrG7tMqtY/yAsj5upaBsMBJOvF+0eqbfqlei+tJaFwyOt5BN1O5l3g
mfhJrouCxgnkkUF3ftRpdcn2XQXGmRakDuwKqx5Dd13yzzxPGj8z2R5jJz3T91SE
UedsQ4CEFX/pO05RBo0hdc4wuk1Z2iIKHGfw3XxXDwf1DNXSmfnxQqKANbYZHwkC
D4lqJ8FNnSEqeIC7QZyeao8pakOx+itcDwd59uWixWDwJAPxFL/ft9asCNDY4nDr
OtpFCbM2Fo8eeVe1GhUykN8sdedqHNNdHDrDiz//YVONNKD1JHMAedkhNXwLpfx7
BjRRGIKyZRXb/SeDSDiRFQXjrVLHimB6HI4x6ltfcnjvKbfz6WsiYGxSJboSZDA8
bVel6k/51DQxZYseUlkFBHVQcxSYcQHV6E7VQDFs0k4mZFu+vfYZCZqqRY+Rqrz+
YyxRiHW1NbU0gJR5SuyBMlxwNpwaBasKA8gujd8YBi1RYIHeOczy0gVtUU/SL1DX
W3D69tEFHPfAT1lZCQxRyP9cbERR3hYNPpkoeXervH1kFiqoE8Ax//PFH6aVh724
bxHLq+m/YwIwSBkLkLykghqcMntkO7Fr/+e3uhTiR8+lRhyXDxw7y6k8uNhtkPIT
jw/JHF2Rtd/iCAH3Uxh06EegZ4duUc31y6EztMYjnz9ElcinoOXNQqyylaOnhZLc
GNgjpnfvVlmV911h0wFnG9bZQlDUHFuw5hkMB8vw9o/AaW9CvQLt+KsLyhW9deWc
kcVTAEWg5tDqQXf8xdfISetgt+jDO42vVtp8nxhlfR5ofGagMxrO5YtJ6qSFgzGy
gO720jGmzHJfvs5InI3jSmc333C9D1ltxY4/XzhBr87T8w64BxYK8nt6bjLd+K3s
9X6zwZc5xuQ7gTri5loy+I1BP2gKlH9MbqpiHAj6mBLRLgaaSaQZODGBgaOkQvHP
ReMZCTByH+meu3Ig2PFqC3zWjB6f9dHwovLXzqF9J+gfIgDWuFy9mw01qgLFAd/g
WJ7w6lUpllbj2OGegm8tF8EFpj0mGLk4ncwLo3C00A0UBZzEHVN0TCD76FMVVSiv
pKCJM4IMiH+vmrIULHmae9xMfRnr3v4hv5he9vZKzNfhTGQkxNlBU88Qk5cn+WYM
blI9WP1W/eaFobKXqQ3s5bHkfmpUd701aEtoL090TUjVPNdpRD7aKeZ3POAUZuho
oJMdGWiwCsupxWnMOdNlh3O7r78IkNGKgVzjjdvlSGCel2czjCqHZR3hVDneEgCr
VW99HctQCg/Sje4AZwhABottDFm2uc6jFGMe8mkf6AlZosbe0l0+4rWPva6k7VGx
naYzw84s++9JXeNIB0R5z1hbOO8MNaK3ey/E5pLt6ImqnvQ/V9IcgeCfDqkDT4Yf
DwcfyKRMrVas2If/44UzGfmZmo//biEaaQFdMXkVWANt/HaajjhmQUqR5tPoTUMI
rhUE0WDNKJWQ0DxRWrvVPBYIv6wszTNjZmspqFng4iyMNy8E2S0oREM6aCWT8q1d
O0D/qiKiaWsAoo3tfULr7QZ1YvSeoTryS5P/unOJj57NNb4UXD/egqRk+P/RVkgy
bOsj7Fl5qukYDjiauzFsUqtIPdt9KrFYFP/UlOPaJB/uMi5XRDyyY+Vw7JjEsqjR
/Xfw4ZZQZK/GJIGu6D/dJfVwPe6wrSxfmy3FKDXkGnKqYqXXfKeZYUl6TD4nvXqV
ftJNp2eJJtiGUPkX/gNB7VnDQ70MNbym6od0X6K9s/L4U92ZgahJ8Vn6SN4XozaT
DLqMZNsMdnjeTDQjD6uN8BLs4Oq6coVNVpXLL9ziadMMGFY2Hwb98v4LRech037w
mtg6Ki4zoRp7R61PSAhFuXZdzNfaEFYB/rgDj/D6iiGuKQRUOEu0s7x7cPViVF/q
zP+WFosy/qYgvX5SVo/8nPp+wYOJxQZ50QYii5SaAAFG7K3bqkuI9e/svgrtGuV5
11LKNx6+K8i8FP3DZw5NG+R47/vtSlmFbB9Nt+iavLYMc9GzQVlNDAapIL1dGxxx
Bzryu71rBRYSOIPVcchBNPdDYPazzirSP/CJm9HyGfeBM7vRJ2KSgjIfSz424tjx
kBNQLocsLsA0K4i8AVhJjO8tmvwAA7fl0sqz0Fgrcmbn41Sk1t6+QDpaZRBGcupB
m7UQrSF/+PH8wfjn5iHDJ8KZlVE5Upf0tMEOqnb6h+T5FqCp6Vmw9Gn77GD6FliV
CptNxzPWiglucsGN+JM6OB6uvyZ1psz/opU9UWDa7XhuKNPSxUvPTQv3DWdamxY8
1Y2xKtUKdPjD2gXFKnTVxGuPcrsg+TI6fLnYGhNevf7t79nwxhy2vWuhg88a307X
+aYktDqrLOLEWd9FpZLjwQ/RlqmmGRilI3N7GsT5BkvoJtedk9E1G+J7o/lQln5o
fhmAp+f5EDlsQrWdT9p589EzJQYIHzwOPsugefyy5ryUCk0LKe0691cngFV0wn0G
ui71Bh7rGPrmUmNu/O02Y5PlkDogDyIIb2J+hLnadtYQqWmIdEoOz+pAEizTh7YF
Vb2I/USm16+rfPmsYNGg+nV36CfQnGrqczLQIeluCc63nQ2bp7xW8/++gLZG62/8
Psp+Y5PJAMKPGnyBnySUpLAipq+/0u9SojSVqawHdengVkH7W3YDYEsfptTIMNKG
ESaHx+FB/4MfyRGBk+2hcfJFayRwcH4WGoSdKIgbdUvYwfbca9WYuHkhLoSOp4er
lKixB6WQgHllqJVcVSkYT2ZsbFlU2aMOHJgpVBXs0PpQiYRjLS1qYkv0UYPDvD8t
Bqg97dr0LRXZhzNvj1yYtILnuX9cnLPatP8A2HuPA8F1FJSVHPyAEAxNIRD2X6V9
hoAE3keEFN3GSy2krDcAH1z6QBNzhO8yKeM6rMiyiUYCpIu7cgUGUCUDZL2Rixr9
1ExRpEBc+rI8AQmOK+kPHpz+SO9dhOQPm7zAgAws8UPTBC47aUhxf0Z8EhsFZeAI
AF/WrFyg+vVbA/x0X+uswjwf+cohLSuRa+3dGEEKxwFVz/+FN2RJ4fA+NutmXHUM
ycGTdpPgzmsIU0KjkFE0HoaF2ZBeFy72aQJZmfroiqViRZ8BgO75U9PP6v0u//bm
oUEepu0/QhmuXyaRFpjS1c447vCW/SbjmVf318yQdYeOEEvgXKgQu06IM5+xyz3G
46mHNzblbtfPSnvWdC5F2mEKagXVV1LMtyD/zNvbwpRzlqEqk3p8q4f1z/hvg7J9
D1Ip0CcIj6OWHdAn0RQhCfN4sJODTlSxINTtXyg9+7IiI0J0f5ZOI2+PLlkRNHpa
/jspR5e5TmbYGeghaN3nwvulUpIFkZbrjI0lCy0HdMdcUCGBGnvW1uL6VMExNsfZ
nBIEgoAAlbEQ19sb2rVyjSJ0mjo7HmSq06kUYtT0514eRYryZsQD+5V2jocJJmX8
XwxjOS4HSnfL8gEFKp7bWwNBJMXFgv9IGXNsLPYNexplOL1uCMrPsaVydX4FtfIi
QorSB2vBet1cEmbCso/vGjpmNpkm6TN2VqnChf+fAgsc64mI6a20qLV0bwwN2mx4
ITbh9OtF+1GsZxRn6hl7k9UNHTKEjosTa73PjWrywJUb7FdzwkRYDhix8kY3k0rx
aX5CIIExNqjauub1q+OMsz3zatchX4QbgDFvm27YHsEI9N9JubuPXwazWQlM3f3i
K7O9p3DfP3g7OPXn5Voxkq+kAb+X8fFBr5RVaW+DacuQkzBnnUDdPvxsNDwM/KvI
7/425LvYX/7AID6VHuooo+pDlFI4OVu2Nnxm9p8fO8cAqXPTfQzcLeZerdEGg4oA
TzOREc76Qoil9bZ5B+kmxGZYbAGvxeH5oTPlw0OzSO7ssCpWS+/MGT7A/UHd/w3U
jIi2eC1a+koPPxXtafrGLMEawkcSWMPC3NCGpcc/egT3beLdZreheJXMoaBRTbZ/
yylqPSExGTmxwfTFuEcw0FFv7jB4QXa7oMJMTU5QBkQI4tQe20Jl/8RMuEh6iUdj
bnwpphMP4eWg6FG5PW5pY+ekxtB9iQhLeCXAlfvgnrhu1bUScTg6EbNL1O55jd1U
2vkHrUPNYdDcbUlEC3ru3l7Zzp8vGoT/rjSshbb1Dj9LuaG79TyUHUhas2cycn7g
aSKIOt+Rhp9r0PsvxxerNW8cap9eC5+neIs8ZS1WlulZ7JeOfkhnfU2AFXLnrtyr
unqH0jOPyxxZ27i0x8KsEhr2IhGUHRLepj6JkrAzGALQxbXIbx9iAVPuRMvBTyhc
i/l0XlGmFawnr9kautt/QkU7gb6DvAT6g5t1cOah8BLd1tDX+KV8EQxDnutbbps3
Dzx21mbsdxpMQGAmgoYkqMV5HUhDygrEVFMpKA8Cm2KvmzqtsvD7hd8fb7hEYoX+
9ZwuvKOvt0Rnz2z8mmqZQumMZGkNn1MtHbLJnBLRpbVFxUdoBNviPkBqGlCwn5L6
7Fd+gaJDkNJ4mMRjOTYDrUsDVtWsqQS9KKllomnglwIBvU05D6hSJHCd4XwjWwJN
yNDwnt7otO2VmDkprMjcvePmZw4yiunQcMSNTTLcknWMB4+mCsbSu81BiGtRDmxj
4m6yTCz0UUWuHp40tHXTeGYPXHA6yJQBEyR9+mlPofA77qgtPIHhJJ0LPxQ8BwxY
fSv+OG9kiUmGrlNTvlbF96tUyZPOr2zhpRji+G3b12swVrVgPSf5a1BK0sq4uWzm
I3yb7zeacuTT4xOPpM1giyBH6LcYZkILRgp8tnvF7opgGxJdMCJvUjaXXIjkCKos
+VMgU5Gwy9iaCzavAau1rFm2/cy8yaut37f8hQB8S7YNS7C+cs3BqkWyOr8pHlk0
2/x2lukP4AO93IAaJmggumxHDPU2F1c6UbZe94CO/u1+cu1UHnQMx8xBoKooxGqr
f6FDwxQfsapimRFk2sLIVkya1DyRBH+56te8lKatr9ZIvq48Hs71w0sSO3DEQkv0
RIIzGn0r6nFvtGq+RC+82TMUb+B82kyvb2rcT5rwU9y01TMQSuCF/6L94onCQjfu
WkDj5migtK/n0avaqwF8ZBMDHhPYNVijlng4L1anBijCcU7gkNTLYYVJKZ/qTboF
XBlEgN6HC9ghIstmbCjnGm0vC4LUTGN9lMv1RN4bA9a9iZeYzJOgpd1h+pvBGqwd
rWZQy4ac4VT848uR1YCoAEKy6DJrJiSUqC5/958BrEKTH8Peo796yD2awolqq2pq
OkwMVu2dqAtih9roT0WPP8a/l7Z0dB/wY5HAjO/P4025yFG2jUimGB41Vjro6/b3
7fLSKvRI1uKciFsng40V1H/n35pzHXQY5xbZdoQtfag0pVVPj/kRTRlQ44TfZjEN
6fZNfnEVHLOpdINHsscYF/Z0jkfUjuYhV0ZI2l/22Gvx8flhSIJseNjF559aCJMd
3iXmrbQuOde5METdh0x5f8bSgNtLGje418quPN29J7Eo3n8m8YtiBFlDLinVKJ1p
KCPUGuBT+hBMbtgZfgI2d8uRa7f6HeVoWT719Khtwp9CAKPyWPhxIi8gSjo2e+7U
JEM7W46XjTu9G5/LJzsx0tKhgR6cCbukXOdhpWr4Q19yxx0Ed4ZnQcyMZ0KS6wOF
pT9ljeXs7gNY/ODHV2NuuWKKkoSc6uBL3D5YXRq3fLfiL/V86V9aHlvcoUEltO39
Lcz9L20q+uwn2BqvgHXYNxTUAGInxCIM09BhlN14RyubnhFyRFeOFsvsdsYXVCxj
yXbn+YbkTjFPoRV29eN5/CODXVEiUUPbbyM7rJHq7m13FM5uvzHFAa/B1ES87RZN
MSFs31+otwJlH+bA5489mzZCEnLqVfRw8fvFu/tmMGizeGFFn3Scv4HlE2FgbRt0
PONxOcShBTbsAVnGZi4lgke47lyHEP74F+e/LkLAVeISGhgRP9whtTMr4QHTxTAj
qikyV62VED7IhGm0aZQJT8o/ORl0arrqvpVoXNCF7qKqiLILU41qWGko3J4JFfuo
swroUtXLXWBsL+rRF26iIL9a4Lflk5lcvMwnbD2xey1rzIXrdF2a4X688SksPfCX
8sG6btqsMqj6QyJSHaCCEmc+t6CTpqC7+BY4/jDmF/EX5Nl/zXnM8DF2Oy/3A6CA
7kuu5MkmYHVQZvtvd0cA2WqOo4KBM+vEkcrY1wgPz2KB/SrLKH/MDEnD9oyamVbM
a5NfqRsOCN2jAE3dF42hv/Dfd0anJ77ijIrZMUWhxQVnBSmmVeDop3JBtlqotxzj
/fyJ1tNm8o1yd+/Q2scpB/aHuClC/GBGr9NabLF85vMrnruT0kiqZo713Awpt6Vu
lRyVoY3/HIAVpjRmAp89lexuUOjVsxkLMQFDHFOiBBU7L/TzRHHmb/bgkK/4UPDj
uUM/gXOgoDADmGlpWoe04CyXUo8wxTixtbH56T6mA7d0qsbUquM5EhbcHuwBRIXp
a/ppGNXzKPpG+ppmayeihXNg6qoWZu5LezYwHfSC/0EGansHTdfPpBlYRB1DZFFK
EqK5u4PDWCZWFcONHu8kcHJ7ficUC80FygxrmpjQMNpnRqpaYBDLAjBbRRb+7vOs
FoeqSsJ25Ux3VjZT8G7RC9hABxMqjIE+wKdTgo7RVN3AJF64v8y9AqGDz587fN3M
9sI7ly3SGBREQAMX3wxdavUotBNNODYU6HZN1cDksHw9SD4qHz5hsxntx8+Xmz9d
vnm7EFfAdAU5WEBPNjWCOaumydQhRm9Sjy5qvylfIFHg1jnA14t+TnAWq2hj1kUG
OnvfMBt5yYoFgYlTinAX8GTQeLZ0fUcTHo5fsz9F7kWjc3MKcaGkh0WCBGTt2P7B
/RddRXcVQj+T/npHfLPPRL8q+YsHtV7WrxjKwRDrDTEoczijNE0+/a+GjYxDArt8
TRnA8jzA9+Rzmn4Okh2wlpp76u8Xw+z60HditKDxzqn8b7rD6qWimbaQ94knoET5
UoDy8vyohYuObtDkKujW4mD1D+i4o6VAIC1rtMiLVvyunA6o+wyru/vUFmfbZq3Q
D3XY9GLkwcrCezEasHUk4N8pAYf6y2oYh0iLYge1eLtopOh4jHsdG0Ldxo7KVuR0
ETBor0F57Ih9rhnKdo6NKBZkLObAXft81s74etEyuRiOqo3oku2kxR/UgZZhO4SY
qJ14pn0HdEiR+CdSS/IbdkG18ztnoqR1DHcBgtO+R8pxMYAVT1LUCzXbd/CqMQG9
g5muJXi97xrBq1EW8tj6DlMZbVK8fFLftucItAvFklenm6AYyfIbbSQybPQcYM4F
kc83AML0oz6UPtdWuuWfoyFSF+QyOWWYhMC7Hlpa9/wxiE3YRm8LoHY6c3NmlfK5
oof/CzsihJuZU6M5+LbeDCKChBAae6H8RCLn2xRkgz1d3+x/2K2VB57qBgCFrQ2e
3V0/09CGuij1oW9YYoO7Bmf774i8WbN80ikjOsxF2ngZ8N+rE9h5p3ZbcGGc8T3H
4JzexBq8vBNgFqjDoQVaqzpyww45lkbRQkhhxi0sqY3bvD8ly3kkc/jykIYJt9eS
vp5IGnAhWzIAF6+pBDCWq69LhgiICvW8zykswOVkVrlGOq6Bpi/DRgB1OxfYIVCB
FRWv5sxFKkwEDs5NFs01u7Rcee3803fJBtnuS/zvgyIOfixTdmK4FBN5Wz+E6XBN
rn5PEpfPqAQ1qAWux60dP2fYlDQeLchUjuAddqtzc9Dsto4C88uNMA5Ik6FQf0ju
JMNUMp8gwk/JFXsI+gESppYrPrwdxAwn2JdKnN7Q57m0wFHWqanvhCAR/RUrTA/M
g4C8bFgmf690iO6BbCxaBoWTKRlIqyj560WtxPRCopUj3vOApikI/Q+RYUCJHBei
77KQCf+P1vqvqSb+tv/PmM4LdDc8cM2QvcYhjd0HljRw1EDL7ZN7ckosY/wF+SA5
vlUGMK7I1jyhtBytZPk4nyo0k2CxOgkkzVdk+S4GCska2KPxY7eozwVnqIXSCdlk
F+0HT733F6it/tQsM40iycY4SGPDoxf9wa7BAbXp0Dgem+3NBEgYzi0LuedasrUY
V3akGyOxEPU+LNQrhx0/baURzbqKcyZ3SQajUdAcmdXwemBOoG3v7pIG7VQgwS1h
3zlKFRrJaAKfPAsHC2RtvnQJ1kYEV3LpZdF9QBAicMRYHLRc+KrZooCev2fUIxQ+
GtqAHlyBBu9uO5Aq4FRxeyJ9BkUKa3gpH/xY2x2Oyz7ajU7pEeLf4Kh0bH270Bo5
Su8SHgYG6oAEeoycuzfBIOCmkLps4Vuu08mMB+6iQ6okB9d+nON1aGXZj3oFsLlF
iXr0X2+c+iRbnbQqw9GGL7B/p2Jp9uPWBK0+ZywacpTTosswcChUjF/e0Jj509ay
8FiqXaJrVP7dr6wRHHPcX6Bqs7vEqDBy35O5Nxf6uW9brLP5AvxRqe/87EwuEd8u
Couvw3oeFN3RUsgOL2lxMytjdcdIQfHPPw/AZ837SofkNgkDU7+duKm+WtDj7nD+
Sv9/6dI1oMyTe0VgGWf2KTwb8cC9c3/9Fm5UcVIjbZo1OcY2lFBZyK5l6D5j5TqA
gD/HKN2EcrDi+aM57RkJRUAy6zVy+SgJt3E3d4d5JQ/LdGxC8mIbEkFmHO+6Csrm
p4lGYYfygvDDqZ27IDc499QsGbnCsuGDAJjX//X67gK2bSGoMf7j44IGSgPcns3o
qpjwKSIcQk7jHJ3tDwHQqVkVRtxpKX/LTc2kntriSPLXFO0OjaIifez8yuo8HeFu
wrgz/h1rYDw0dATQHq5VYufXKKz5oFlb7L4ZLwGa5tEODaAENvzqjywuNlXcHKt/
+8s193Is/Y0v6/accG1YWbiWod6tqQVelfbxekBV6XUu5B68+jt43q6exBbj3h+X
EzpfriA8Zp9FtUj1d4Yyg6UG9vubE11adzgJQfIA11A80ljaFvi5KMroLLOGiI1y
Bgry4+ocfccsLbrZJrkZB5jEeSRAWsbvv2wjA245TKWREaNdvbBEayYqyKV7leNW
1eop6rI1fJAfm0F7KDmLl9Hv8eOCU4LsdQvImAJfERAv/P42jFk42QS9xkLSrtdw
0XsHtyLPf9l8iDgpayPixAvP0+COQE8+Lda1pQ+AcfsjTCYn7EALdPUFv5CphN7e
EosXteS7AlvFe2DdSaw6JwZ86eu0IpeBtX8R5yzIHVDz2CyVNkRswmAck7lm9X4p
h4wW1sj37KbqNXMdoO/Pl1jfxFEJ8O2sJdFOR1/Qy79xas+qKnP2sLgrimEKDSBI
mmCRozjjgR5Kq0Sd/Aai7sB+SZ5SC6u0CFkegmbDEecdHsET39YYQmzDNe52h3R8
d1DUtG+kMzXK7nMvacehhLlm0v98WxrdY79BAcLnPisLx22vvHx21Ses7mkGk7bC
VCJZb0k83gYv9BFGS8tluRD3nDtbXphhcFsbT/eohbZJxikVgN9vL4nrR/XYlb6a
WcNQifx1ZXgkl/zq+1wACjLitwb9oGIBKpeOWF1IE4K3Vke572lTSlsf9iT3utGa
HQrIIM6Sin4R4R24af6O/GEjlJv0fJTIcZCMtaDGUyRjOjs+4z44Q7R7xkWbdiUJ
r3derVvu70F7wKTs2zi7ySJuoycwzGdBzXfBIUfWXjw22sDNvE6/xFbqdG0pSgMT
tlB0S73/n+u3Id9JT39u7SZyje9p18ThmcFMohDLOtMFfGeenipN9HZlssy6+evs
LxJkEaOLTuFg6kKNIYxliG/V7Uvw+4HFdZwTZdwwjI3/M3ci5IkFPuNvBB+Mal6h
RZv0uRmsKwKJtd9PXjFinMTzw0z0VLI1QEuZcNGwokMd3hy8/hIDQyDuVF1QNdej
3pCtYcrYx2d8bHUV4vYVJxH4VFKQg5dLX2AF14l7nV15mUUw7XcoJON77sikChcn
uf7fm4QDYVNsu0YKaZU+1KkxtHVsQsavf39u0uJ4zPFBfEgnYHxOjHqbc3W3FNRI
rAJo5fhhfwUYNzjkqI3gEkUmRXQ6r3d0IPPdJmClaE7GWthRTgYKcJiIyNre5w6g
XuvOBKXLmfGZzpAKBnnMT44eXdUBARZ57DWmzbZvWfmHGNfH59tMl4M5BbbSYXQt
eojX6aJR2rEXdfnEZOOYboTcXkCrOC7eYQYVOOJlM7LAmCqd28aXmkkQoSef2Dhg
/3h5Eu5Wj1/o29dEcoyh0YeHl/pmlibUj3cUF07vTo+i0e5UWAUiTndjTtTReTou
jJAgjT7Vs/XPoCqfZCmEE3Xj40P0aGKKs8pbbPtfTefiWrpBYRDnB0r6gWdlI9jw
feMC8MeCBKZ2n2f1DGfAlZ1Uksyw7l+iPfbIT1V8kHcIyFhvyRR28se7uT0h3QB5
GBbBkfjuZE1lhLLhLHbfOXmYkPEKiXoYNTd5yRCyFoPlnHC1Cn+jAGwslyQIRQvq
lFcKQazAXxEsFCd3jEt2XQqULWADu5O7+49z8O1oM4p1nJYXLEjr9YpOJyEJ9rjI
bxo378wjiLxdtbrF9re1lQ4nz/1S67rC9Byv+eQY61vNO/cSja0jes7BH4aaUCfV
08pgW9QnkcKQBD27YYqCADjtVqcgiHL0T0xYtFMUqs58zyA/kK2COVcrzhndPM2x
w2U5J6G90A/PJjPqN0w/TRcXDjkkj0FmYNAWMcqFOZUKToctagh9e0QUa9+Ik0il
I7iCTX+cIcKfNepW3fiIh87J8Um5gwBbPwFfj1qvugtpsI8dd/3c5H8sBawfrPYr
N7T0iEi0Yyg8VWWlPhG9DBSE+GLqs7X43Ihi/PUjSgIkKLyoJd30Y7I+pS1paMsS
736KJGmJCdeB1MxGSSoS7HJL5YLoLD7rTR/2NFlRlZIhYt6aOPpq9yZ8A5dM4QUD
fWQSaqG1MPXPt5IFYkK+oTtKjej4XoulwCX/Cs2bloHWwNt2yMrfRKn+G7CPrLhr
H0B2m35x+6zktR64viFRl2dUijtKuGMd+nJRb1Fi9vbxwGvSN45dt0cRAMDVtlUW
R9pTec3C4fa+YdMFCZtvybr1PdXNwWmlJFUK/PrWxsvoTscaOm5prpfUN3J8rBT4
wXXDxAZ09eeTLGZC3mACEvysILmLMrvfc94U50pqKPSQNcSXRJymCj7IMFalt6A7
ijDVA+HzYRvey1lY2hIxKFbTJicxZZPi3rX+a6ppzbdsup+GighBakpwwdbLgpiD
CiP+LTVSh6aeyYBhOtJyxKKcYhTfKCZ7bRnb8RF0eMXJXgkxGt1P48jvVwyvIILI
R2VXBMnVMgDD5QdWaOPF2TIpplbieTDcLwzyTHQFb6fzzjoB2Q6KAm5JNdM04doO
EKHI80K+YtRjkplYJDOX5q5T8Mm8zgvi3FI/4PQHZpPxLXOJzUyFohNg27JHKiYV
AeBKWvY208bm6jDI0niAEwtA8eF5tzTT08BYmD5SqvTR0qo5V4SkitPrfKajN2Nn
0YwDIXoO0MYsMIl+j12i9o7ON4xtKXROGrIMZrKQJdEKmLEuXDX0mNDy3CpilIo7
7xsyEg2/uczD123l02aIK4njEJ3VaCY93RU1fSQ6dlPr6+iJY2NcT+3LvILd51hP
2MgyR/FEt4ca6avM2Dmeg8JHnfvWgGe3rjCPfwbAm/DI1JtM8FRjj19vIStikfXh
R743NhSk7TyC4oM7zD8UoAPOqfVSwhf6oLGNlEEEzZDrdffyaD50vi+ZYY7X31qX
1EbeBT2wrLjeGXp549J5JwzE9j4ADVitzKBlQL0eZVmB7S98lvytHLhV53QjEAn4
pRJyBk3ZJMJmlKKg2W+VWU7BiEQSPC0JnJT2VR+fGRuPM5ZdSk5Ty61IcxO0gNtJ
EQI2e9Ygp9+XiWQrj5blWdx1FfQUdu+wmYdPz22j96iMrWnkAG7eN2fflAqrdL9A
kN2GjNOSuhCP94SLvs+i7OPELeSbYdiO/15zX4OLyUlr/DChIqB1kdbLbcuvBb7w
O4WByd62JMn6s8q/Cse98lv8jytpdpon1a2szgQLeIDTcRDfPqtlz6b5A07g6/xc
9vkawYuFC8ecTn5AZX5SpEjeaZG4EB/CJFUIBTUtsD4B09ou4WodXGbvlee6xU+E
qmmjTwHb1vo3udOS+OOE3PDqWD+L4ZzrYl2LWD74Jrh7lK29QAUSeWZ9ef8NG8Jb
uZYKhjjb8J7E3Y77hybXPLiU/jmBX76+EvT8dECjQmlZBfO15GWZhHp3YyQhrtEk
lmfjzdmf76YrlUCSwLBCBlpMH5vGR8DIr70QOSe3xpz4a+JIobai9lg1dYhVfNoy
RpZMkAjAitswFcEWmzfARvqpJIsalvgS1bukJIrOPeHACCoV8ZnJMUNJ6j/4oFji
ig+pJ62IXY72pmBExI/ni4fnQL0N01iyrg9yRqfsLhBFI3JX/nT7Jm31LcD/jPy8
BQaOKkqhd0r32E5uEpUmUkU02+hrieJgVWd0ZHmsQVf8gIdt+jyM/q39jLCq46j1
2crlvH6H6oJ0EuyRMIvdU8/UFbOxGK/ig0vBZmD5Ubh3klcIact5l456rqUw4VDu
2x5Oq/U731Y+zhkX70VOO7gsAgFLOdEge559HcuXKuxi+E75KpFdnOEe1vAMTUuy
9+p3hDq74ZhY1ytUyFYQgiSfK+ypX6HcFmTLNIbvHBw8xmMV/KhBcUgrzcP4Jsx7
TLal9pjkpoPaklMtPv+DBGcxadTyZg4eGxgW5Tt+jQkHk/DHsAOqfMQ8N5lZMOo7
kV2G15rDDdvkKRiZ9LB0s9y9ih0ePGZNEkh9o2nmPpAp5CTPrs2tUMfe/t2+lGsL
cxIHgVIzioZEvn+VS8/XpRgq5/XsqXxrnHSs6Jlo0CL+8YgHS0TbSgrs1Xu7ZJVP
5TWCx5VxQLD9acNS/po0TJ9sMwwd59JWQwIOmoKQeHOvTvbFYcKFZqF4/YQjcrix
KuPxwTu387KFBRPmETCQZmKAW3XNQbEk62Fp24ftpNyTRqKxw4xcNyZEd/bVKmay
iufMM55ggvQVIh5VZPXVv4wIO7w2+tcidEv8QRYoEZJ93+wIO6zewFhyc5nkiMTK
pJ9tty3jl1xrDnUa6+hUrhuJGSRT76KbnlwgkQnyOrYYuISzjR2EYVUe6TYPgEaj
K0nbDZoJl4LqRWdEWINbpPRRhtZOuL7oBGPt80n23OmX1faJ489d48cMZTDdxICq
R7Ff3w0jnETJrIz5aw3LScrtLd3E8hKaHHyc7jwTH6L9GOi5s3J6g+jFksduDRqz
ckv90+qpjiFqOBq0HpK0SQXWHuTwXeB3Cx/w/t3vvOPVOl7eQVuG82g1+z04ATq1
WsMq4blJcsxCaHXq8oVkQBCc+j8YJ6tWNxobuMjUJ9nBmHQXq0CUch73yNp7VPnl
03RkPmSktht7UNj6RXOhDIbHQ4EsoxFJiiHl13CPZyOQustSekMdiuMtL52FfLIB
PSOOLQL3KIFPDqkeb07upYgzuSfvCyblE/iK8FGFLaWDR9szYGVXudzavUvjmVqT
HQyYDwX0j0gRzEhIBOIxEJ+OTW5Cr+j1bz0lQf6JBanz1YHatQ9TtZTbbcxnWk5/
SsxEz9Ld0/b4CKZ8Aa/qt1kTez7aHYI6bljXqouwaWEGT+JgTf3fv7rQzr9wZDZa
1eIZmtXtY4TnBCyAMt4uzd/7POFxdsT56MKiZt1l18sbwkZvT5jlxjfpDRz9pdJ2
ReBUS9Xf+TIOAT3Zet6QSuoC9yGt1S11+N0sj+DM+PLrmZlJDffG5WXtV3yAt81g
pGW5leuhPjBfrvZRn9DhW17CREkZAvun1OcpbOsApy9K5O6gpZeYbvnlNEII2Ydm
0F5qM2A2TS1Tf/14THCk/7/B6LCT1E7mG85oTyrAoke9BU7tMx1mmAGJEOjgzP/V
oPGYs043UzX28Nd+nBfTUUCk1jRTGoSNqzw+VeXO2XYVd1TKlRsmh45Q49afPd/7
/G99emjfUoUPty784xUFgvBxHeEgZnLAye5RvQJn1DTv0XXxtPVMP78FYNiLMHU/
8JDfkyKztZn3EpbLo0vnmXBplwk9HOUFrwsHzGY/bwfH85oy7ijA9evcKCNKCJpE
9B+BRzcKTsipyO6jUsXbNlGrT/yXspix3InjriTDFAjN0PWNkiyWT1R5eIj6T9z7
ZOQUT+QRsspnjtSEkMKd+sATdJfjbylD9tAh4rATTJDFIT9FRWvdd3FU3LDP3RBy
axC6wo5jn4q+aXLXARO2fUNJpM0Qf1+pns8Ccne4T+dYh+AT10MHlQBRpSBUSiKS
nhRj3MmDhvOvDtBIeasAWUi3SmLoZcXP78yT2iDhryzJvc+a9uLKHorKJeHouhJ+
9MM7AQhJa/4x+N9XcAUkF2awZbbgH8sGDjUzQhP47jP/wSac38UiZi1F20+QBbmE
JuAOcbhacFpRkXJLQyJhjSDc+5CQkee4H4Sx/5UofxmxthLciABtdnl8Tk0uGUZE
Xt0TZY6gl7qV/x7FpL0i+hQCwGjjiyU+VJZrPZ6n5ycOs2FKG9UNlT7VbwvozXGA
O8VffljSpeK11OIBpT4ZPKIdkdynPEDHhUhHxpCN/EnC5LGn0dOEennx6c3UsflN
bY8dO0ZiSTo3HQdCZRF5EViODkz3Mn505a5q8mMo8CMP0su3pyd2uuWkr0wBKaLo
B14tEiTVSJQ/LNnhrHoy5/+F4VWz8zEzlAWlKfmk/pNSRStcXBEjBjAghkYSu+Ar
mHqF+Sh7gqLTL5UcvlTRwWiEJDAzkin8ue7Fc3JQ7KZ0/BRTekuiCYy3lM3RwmyM
GeDFMn7AMrd9Rgm0XVSgseezwmFN5SF5EyJAWAykthvFivrOShbKW87kWxZdsgiC
1NVPT4kyCtRmQ//F6aGAs7ml321rmIpIeRic7r5iybs2S7+dHlN+9qxSQQ1joW9+
4d9jfsEO3HW1vp50+aYpG+tna+NvkIR8yFmP8mgtSHrYlTySu3D1l7H00YRPfvIi
fUKYT49YroMVfEB/jih+r/llc6RQFGdsaDKgMuO7ciN4jut9o5VrjQHpNP5/UQLF
LoIZ9FMq2xPrknp0g0QpauK3A7xnM5TK4c6XVog3BzsDfr+PoBrZIxnNQQoa23fI
qr9LfDuiLCeIUH6xkhalK4VLGGOGd//kzh1q/jLP8/X+FAuScQQyLmgpOaCn4epW
x8mVGnIXFCht3N1A/aiNzPoXgP/HI4icCrufaIixwsNCrxqnZghxSLiAmIgZbNYc
NHQPsvCpcSzgMcUyHHx6EYoF6FqvttAs3n9suetH/iMzVdED0AufsvrL8EztiCX3
/fkc5cK5nfUR6+x83QZsSphACPDQp5yi/W/R1gNO4ZeDGu5Ir1RxmKj3g1EVwgVW
LmcrqHXMED4VnkbR+mMYb5l6RZfs9pRUN028aOPiCO3vRJb8dIS0x2uFeFrCf7IG
L/ChgLVr2MkxqDdTdloNDkyPLYbnk065x5+dJ+WFoTRxHQ5Z2RoW2BKrZ2SlnC+F
3tjwred/bLM9I5vYbM1EMpOIqkSsr+ZlO9yklDHple7MzSz0mgFKPXOmzenuSj0x
5jwlWayujA1dBZERxIRWoFptX4xytF2CBWNlOBy2Z0LnnRWQVXhtdsq9jO9zrkbf
zBCKY0w2YRZgOiEteX6ZFs5ILxygSn2KkXS3n7IPkEYZNddCpzZIB2Z3PAXPk504
PtQDc/xGGPOrsrFNBnCAqX8wH+Amv50e1Aiu39RZuordhVk5rxuEqkxqFzf/mCYF
GOro0IA01MpXYxAz9yc/I8lnuen5jSqE2Gv20VHQva8lTy24M1oSXemrj3S6N2lC
Frwb3ORgherXFtAeGd1HeVJYDxilPJUNf+r9Qev9UT0+KMTlq2l7hy7FLYMbnEGm
BQp5EA8gdSuvgeG05QOJlaNnTMxzV9e1YLb2MXmJi+mQBzPZvoM+jjUGcAQl+/nL
a3kizRPHhlwPLCbw8hLeSxlMnCsFP5rFLnHQbyO/ZdqIs6Q3Bac35N5/g3aR15ba
KEaBi8nIgvK/wIh4QFCCcKD7JyuSaCIRHcA2X13wS4LWhak+LxOa/HVzziOXKpOi
4IkWifP8qMlKkuIG0wd4s66K9d74RCmglDczdujwFvraMOFYVDvzpCaHvgpLpmFq
ta2uFBH+eVVg9c5x8JNi3ihPSFqhCkwGec1BOYKq/liWzSA5ChtHRPoSnKFTM1/Y
Je3d5N/zaXfyJSqPzFk9fLwJtyOYQf3ZdDtXIfgozAEahFqBQXITUikydDgKLM1t
0j4azrbmAJnP3nbPytCWkby4oq5/faWjOiRb68fbwNfn6+IJIg7gEWfroZtVp+ki
k8OX2TVVYU521t1XFVqV5xxx1+38D8Gra85eHSzbXu4Zy4eJTY+7pbot4JIxXZfR
HPOdGnYbjxAW8VoMbnN1IvCECSapy6v0aILDlBIclnSAjvt+xcgGl7CIWtrM5BIL
ViDnATyJ6EBymqjSUHnvSTebkFQV1yfJhKFPOi6dbco984gTWB7JfTtNETT+dhmR
ENz2RLmSqEgd5CgtVHNVQmHH3ryL9vYZJSFxqQUtY7EYU8+Tj2ajpuX9ByreAIEC
F/qAW9QSAKxSui0S4/iU72P/wieOuGEBeOfp6qm58+POVd5X307Hf1cx+RVZacjl
z4iLiULDqBK4thNRcDjo+ofLieYj2O/bdH2wr0BGfRrcbVg1HR706DgICM4mlD2H
4VoNi1QGlY0XOBvxSsxRGByaVQ9/8wMmeogelKQ45GKw6TUN9sQNvdd/ZcJqkvNr
eeZwwDpvkFhTh7JgmqhGPvASUEpRFONTEghOU1v0W5p0kxhQNA813KYmgrnZsPb/
9S6WDLIW+HuhnyeCWwjIYaBz/aRetIsRf/o/Xcu/aixdmecqKjCPrUeR5snQYYUM
0mdQ+lWXDMzzss5YYcK/ybRvZw5TM/QKc3toaSyUOX70H2kcMFWqbwDdKsIrcr0l
z5kqnjyNPa9rxOASpxBRJ9m66ZHTGqRSCZ6Lj7r9SJJRydxiOXLVTav/NCsK4fH0
QHnhU3FyCbvLBWaXba0DRJo744QOrAdRONSMBwGk5eA=
`protect end_protected