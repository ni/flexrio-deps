`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3824 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
/vEkqJfyK/81z5lf9X8oFdXiMosQ58m/ChBRu0cPvtaaDeicOQ6LYqiBRJBiG8jd
Xvzcl4LMEAOMT00vY4oVYyrSfy9Kc/8bBkA98oLKdWC2ZiO7whyFkpeeiZKNTCpz
ca8UfrGPb+IF7ihHdnX0ty4cY7T1lQNDFUPhyyNnJVGwu1ablZbHM+xPPbv5MczB
DqxIGQUvTy99NxeEXspyjvtX3kYoQdueMN+A9qhMfI2sXJvZiFyUeIw9Ziqq+iwx
18wZ/ZCN9VcdK0UQn57AU4qLO3a3iqK6He2hr0hxd4ZuZZ95eXEz1yYuuGNcny0+
xmqQgZxdez9jAqnPEmYR+Fp8XI44KuWr2v8bQqrmjDCSXwtF9AgVZQogFYFEoUUP
pcyTqUefdYdHqB7UYhsQ8BrmyzPt/TsCypJnCAe5c43Ogfc7/DaC5prLkBdSvmNW
8a/Yf8zb/+EoRWXeLQaTcVJRuQDOFvk/3pYaVj+b3jMpGNP1lsXryAYyYqp2sUDH
2J5NWcqDWCR+BG1UPRS12T3ayZgJm/gZeSJMSzXZ3e6mAu9u/m8pyoxlODhZEfQJ
JylxI36AY/VfQ8QWh1QerRgS6O2aV8nm16muyf57vUZBbj1W3hNjRjCAnajiqR3t
7/lPzjhxbMbXq00KIvRepJYnAyY5wwKUiHaXKUeUMgF1jAC4X14TkQ4MxISUGRTI
WKTsO42xH10qVYJBuAMCNwrsi50+oa2cwgmOrCKIkiQSvAOGQywz/cEobSvYU2jX
ReJ+j0KuUpjgclHo1mFa4bWOyvUXZPb0MZjT0kwYwcUeC19PeHJHs+f2RROw77fg
3JyyLw00/BFFNYLqVxx9kYSn4v55PhDgoG5ebtWsqlvt/qu4zHqT3h7A4JyXl+bP
y5+JD5W22DumgRLfDvBmh0lqG3OvOTODPG78pjUy4niYxRyxMwP7S1oOhTpGJecy
jACelmDMQF759LIv27uHYpVl+wTkpJycKITBGoYofwswdjNMErlOL9RxSlY2+MQI
c+DQ7wP09C1TvzRvLjT3XicBlbE7xVykyTUvQ3dOc0NyCeEuTDGGnAMmTyoqcFUC
6BwQ82hukQ7OJgKGgEgbchIqtCVn2wZD6jS8CQ9lFc1bmbIgtBEW3lH7xGaxbrYJ
RT0IslESHXBi80ZCe/cxnrBOYE+KWzyV3q/RFoSh/WjFZ9I2SB6N0xVOSWn4r+ON
UevNIhwGT9GYoYmBFk0uESdYywyOk01HYvAC3UYgWvqsrPj/I7Yg33ol0vTzEcnE
E6M7K1rHHzqKlrbb/VO3HHNHCcfBm2Er/SmR24fr3OGAQRFgLDXtap+evtUhoEnF
zGc6cTCEOcv5ojSk/EjbQw0qWL7NrWDyYphI6s30TPy2dxxr6EdIqXNH53so0Mba
xI2u6Y2D0UdqDDQGQHDT2k8GvlNAe14rF/brIZtOabmVw5HYEujpIfsT331c2Qci
WTjDy9dP4mEdoXnC+M8qj1ZvOZJw7Ycx1tF2aY5LcnL+Iqb/W7Tkt8C2AmUplZtl
AfDuu9b9w1awCnwV56KagPowuGjCXhUaXBZVnx2bH7U7VeHuvV6969Jn1rLngNYT
pfky8sCSK/EDQDkAlFA+4R7s3Sv7hVMAXxp5JW/jeq2ixml8tFACrfcUlijk34Bq
Kr0qsr2aJRTbE2tbgU+E3TGw0541V1/6sziLoFtjmkoSK/2QY7Zz4C5k9q4yMuYD
DLQ+R5lpui7/fjV/o2cnTL3WLSp4Nw7HDBbmCfv5pLn3R3xa6EKcgCIZ6Z2gwfVL
yL/S/lTtmHDuvhKjYhRNTyNWeR1lxkmoQGMGrFlYjnfi84vzQU4M2KqZ0YcOlyeo
csw1RY9Pjlt2v5D8Ji/UbGlfBqw1bOSEl8JPe/biBcOTYkKCHnjMM0h0WAfM7dQx
9KmKRvTU0vM8ykia7+mtZkoOUu+DX0m1Pov1HBBTbCCejomISqUvMT9VeE5/QfFl
kqR6tTHAQCvhez1Kj70O9C2zjw2/4hcXT26KigGK2s6eaU4X5CsFfpwzT2V3kZmI
LHjSjrw5RC+EXEeCuyJb2sNrzIGjVYSWFBkcWCiS5a3KqqEnTrC1dmvp4e6odMhn
Tu7HBUWnJE013GuAsi7Z98CtQAFxXKSPwOjPgQC5vv84yquo6SIKOtElLAJOSKhO
Zm2AphqmtN7ljSW85JfvgunEVWXuDPKRDtHxxIj3brr4jdZX6iiZ7TRdrnGz4wDY
Q9goyO8bjV6pM0pMNOtrj/5totbv5vNyDfvjX6S+3q2RX61NSjLKLTmOIYMRMriI
/YcVrWp4fM0lOXYRy214Yo2ruy4ZUrXpmKRFf8iEwwJDsj7wBgf6plV77eI21pYE
++0iX0j53tWnxCYbp9fS8V4RA6c3ppF8anJUx1USOgIVeqGsMlgTQkWiglbu78Nk
4NIauBCma9phNgqXcuIuvFQ6KubXMcO1Qi1pceM0ckkMOTGHNv1fSWCZ+qH0JNRt
50CMBtbCM/TLxn6l/i9PfMUE5QnGlGFMXFHQdqjkKCCElbVmCd9hqmdapMUhfrDP
LNdwtsMeJNtCp5mbapQKbbWWYCWEsu6SugCjK1Z6ehkb2E6HoWEOiHVGwA5dYA3Y
k5PWZcb6YtQp/cvMExVbEKu43I/f6CGnQhwHFs0cMeAKVhEkf3g4WwVX/VV4IHSF
rBUmNsiFJRaKoivu69gigwTCDZywY/KvkNGIFG7zV7JpI7Ihq57Ly+h1EfoewtJJ
81BE68NMeMLIwkKT7zhvhE8Z6vUc4peZkSPn4tbEs8XdTA5ZC7unAeSFfs51x+XY
l2h1RruehVY06PaXETPlQ+cTgRJKfiES6y5xzcSf1j6hkWGck2ClDGPpnHHhAZ6b
CWj3n8r7d4qV5HGXSX18ebj+YTQI7LdqueXJxP87uYeyGhmuxjx9Oggdumv8Fm2w
bjkv3C8jRhawFXkv5stHFQnFlm55+tJQU41ILR6YiicNdRybKnrR+kCMWTZuCcbZ
WlI26upa3B5ii1G/t3vm+4G7Us1CKRFaxkDuvCsLrk65qSG3DZVCaJ7IcE58drOW
rCrxUillyVdOVyB762A84F8e9ELfsCdwVHtBovSnejKJtI3vq6yOBqxkTVIrsMp1
VLSvADR7wyQF+wLTOxwErFq9Oqk7c6c159K0jDELCpSJGDq7JbhxZmQCYNFOMLp/
7rEOuZda5jYss890KxXrR5Pvb53GYb58ikqf9ys3HFn0mQwc1/+EVa1croAfYC+3
8o6Bn7X8siXkNhCd7u+In2kXB/7n/Keq43ylZGKeydacDgtv1m2obVf1EIDeu7xs
ObvloANiyWDvYFAJAD3E4/b6RUTRgvLDogKdUppoGBEaBmDuRBsEdDXwG9Hjsx0M
OxOiDnHY3QV3hmTBXvZAjlFjGK0wZl++79/ZAzPZB0S33A9Ql6B+ClI7gcOINI5z
hFzBOLtQYjqZXecTc7R/yzTBYMGVoRLCT6u7houO+bMZscgcVmS2prvse3CI2e+e
zjqeqmYCIO1ehskV13HOlz02hpdtcDss+1u2GLpebbBevEYr/rpw/nWvB8FEXHul
BNgElMjXZIexb/UrkYmADBUJOVeEPUqYs15NmVGkdA6df9KXr7COweofManW5mGx
IC1xdPXME2sZoLYfJzA7oRLcpgVdXBXT2rc3RFwQ0CLzSvgBpwtfIVmVSxZrGdr+
j3jO2b6FYahpnO56nH20SNY/sSiqNf7iMKYnit92ZtbpcMx5cGNUOJWHXOMQa8Jk
JJwfcyQrOaENkfKp9Id5tXeC8cNCNkuYzuvMBjjoCAO2XKQys/RT/6vu5wdTvLMh
RQBQSjPhl9wNU+yimZqmion4PyyHCjOe98e/8Y/uit+NcxHyuCu5Xx98NPZnO1wN
9NeEhUGMaBxVvc7RJwLs27xaFDAPlu7N3aG4akm/g0/YgzUSE/IBpcJ8UhJWMRNM
P0AkSsauFrjYoRD5X7lsF22UxzUuQwOrI65Q7hw2psBTOF4Av3Q8R/gfD0UVX3w3
xke0z3oSVL78UEjvYjRrJkQOHShV1KZmhi2bAswVQ2wUeUAZXDfmc17uKUuvnzxP
2TGNGz8PHG4kVp0kG827+QdgBXe2psbb/wBeEW8897L3sGM7WopuJqCWdrRWDg96
ggH+ks4US6K8fHG7yBacaaSn+o4EEHL12JMrlyyopteH9yGEfDKc0eprkrkTDYbC
4Oi19H46A0Lkv5b9OSfkHm1LQzA6QV1IJQUT+tZ9LGtu4ePaVq0ok7L3OcyhIMPH
2UQHvwtx68Nis2PaxSO/WtajmCsWpLJENlau+3hh20jHSvc31T4FBRumGXNyAPKF
i8vJh8PbkD6lXzPhma8ALEdEh0ABSi7guAIbnYhb1Jf/gFQXWqlSSHEscMpulWaB
JYK7/OA3U71UN3yRX5yLdXFgX3onZcsWYFhGXsi0cI1xTh5bqKlZlU74y9+gZqjj
ZCv/SRlr3goiHTorec4UBOI+oU1w20bfCgHyl0iM4n87L+K8L17uX/UCwLeSAUs0
w06NTG/oZMfmd6F8qjzaKxIh5s42SJXUjhlMmCA59nI97cotW1S6l10QYulNvf7A
EWYHV8HJTk0iefUSyHGOZWw7DbTVEWXWtMTlSRoIz3ZpnFviSSUfKBVnI3jehVLR
0cTQ4vh3//AfUYxc78lSEDBsn4EgHe1mvVng0ilR8vIoLQRZWQYE9LY7pH4Z2OhJ
po7xlp105G0FcAj4U2qnf3I27+q7DO5yXHHM9rj5EMLkRhWnQQcxsEYq8jYuzH0+
ywPEFPPq/UDaj16yATDsnxj/f/ElUSkt6LJqkMIJKgdQ8VVxHxbhvgl8Fxr8TCmk
zzDjwnSfiRusp9cO6t+Mkp6livYGDlpiX6qA7yuRPlxVauCT3nQJHCCIM1tu2DNg
mDe9TgX0UQzmcFFn0YnMsRFHVnSKAxVls3FTxDnYfcs=
`protect end_protected