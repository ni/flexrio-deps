`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3328 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
VKWNRQF+vfUNEEp7apOJOfj548SAgouC4afqmlR4p1DUPURq4UK/H0Bf14HmB07R
8I5sigoQ/XnEx7tnXsOn6Et8pkObYalbDBt5f5fxn1+3yEJ75nTC+oqS4ixUuTeb
Yz+UotxfWmQ34J62JeyAO1rUkEaLLOZkCCIuIaFZ+m56FlBd9movObT9mk1UW3U6
eJ+MJHfeQShjaTGQaXUdooKlKI6klOGqnm8UYaLXjZqjdw8gisWAsuAoUIw6Mekh
BszERYytXrBeB+GCArTD2HJc7wGqY+CnX6H1TY+eYHCYGJXVyGZeeUSODkNflQjZ
hXCoxt8YSVPqYugFQatGVAfffC4myGhbKWROSCxVnhQTVQNFY4BmjBnpd0OpkDeH
BDVURV0x6JmNxlKxs9l5NlYpSscbXoRb5RkX50rY4xSG3HTjf9OKH3SpUBK8ZiBP
P8tR/8e9BA0q9KF1xAE1cdd0dk6MbjKc2cT+XX4xzGKDyw0EzoQVZrRc5m+1JtyA
1FujfSja0W3DIuSzN5lKVghElPa4EiC+zRG4uprJYBJYFKh8NmnlX7zpPbjFQM+o
B6hnOvibtOYXzTDfJiBJF1evlgUN/IAn7SxxA+5IWXDNUVhwQTb8y8UpXacUP/ZN
X7zSs3V9EG6O3PeVTHge3cPBbxW101RFU82ZHlS2Q7ULWE0zhLdWEIoPV3BjV2Vu
66NS45jhrYFsdz2pSlS4lYtoIl4vooebD1osmLSA/r4l6YBPZ8N6eoC1/Wto4lc4
6Uk0yEOR7qfGTC4kjwdE0WZ3i9iZvJD8DJ83bSHUuglm83gTCG2II5Q5m0rbKBcn
tZT6I9O09+CUmbW4m21Dp79sOth9W9Jo0FeMLN5tmrcUb7o9mVY4BQtRtwHy9Ng9
hmCpmjRLFEDrbw5mJApKoZG7S2ImyzC/c8paxev80y+cRjSuXKMV4IksrNoVofLM
hLuec236nR2rd2jHejCxyHcT/peIYEaWareGNHLl4LXbblepy5Df4wVJqRKDxhmS
DbCUZFXKwKpGtq9Szu8y3zAAYqgAIrh3TsGjGcHjlaFL7Y7HfcRYB8gYf8kfVDTg
JLakf1vm3k61Ou4PecW6zvZVD/JNAK/+m+BFkshT1teiIf8WnmCsGTHOA7EYyPbK
ws5vvYOv77pNcmv4VYQ3//QfjzeenVhjK8xIhftEJpZzxE6e7nuZMqszOPmEf11h
0PS3Q1MQ9DxD+jO+3pX5iy0Uw+uh/44sYFVyit8RCpUtIV11nOXeFjHROex/TyXD
AKr8h1heexX+MCM/XuooEtRse4+t71CcTUC0fAxDZWJBsRj4nPdODm4/lE1Q+Ewo
8RKaVaNHr7vJi8eu+vCM8ZDnRbdp1oQLnMh9QsoyGorvYHslIONxReyV5hyloKNB
99EKRtxEBDBLDPNNrIrRv+y3RU7MkOM/fyGYDLiVDIvJBW2tjAjKDfW3cL4twSRB
HLnUly+fDwEVU69Bx+2mHFi8NhWJaYRrWSbNIeE7QC/ifxs+3x1WVU4kP8fahKwY
kiuDoaZUW5YUm8DHQfZVYtM7GmtpnNH0n3+15kGClFiw2ty5IFhpfGsvwNbXfsNg
lzCSob5WMv7hsE+KyIbd2ckz/J+JmIi4rJJiZzA5CGSJtpk74m2tRAqqDnPd3T4c
FAT6vckv95UQLORzlCGsWgi4l7VoPlDRWq3UTOfzi0xQePorw9oL/WMVuJhrRhO+
V61qFjbj+Zb1EyPit4Cvvtn1tUwU4zMIOrzir51BBcJccYX8fw/rEnTCEo3PlkW4
UOws6tM/RrYM3rVsQ3O9K8SNHGx+VNAV03yR6pIDUJxq0Y4uRxm15oGu+bUAg9VQ
uOLlmZRgNENhYvkTgcMv5zfPE3A13nzW5qdYfpgKIlbXYt8IjUi6TCNZ/cBXj5ip
q3pWMqoyOuTCBhHULwckYUYphtQcII9PqbD0V9D28VszZNJGuxA9Pka/g66gFT4X
ihfdUjQBX2k058kBKXwb6UP5SPb7iWDDX67PuRDwFO+WH8ZCrYsfez/YqY8hUX4S
Ezsj2auSLOfo/Dohf+8WYVFrntWeqibrPDRdakqD2jMznB+0Fa19xl1A75cr1d5b
cTV2H9EdG9H/L/HTiYdxwVD01KLoztz3SUzq3y8H3H4kzyYIIQIttTA4JPEaOnNM
SupxATaqayv3WxhI7do/qmB9252Rjnk98wbSFXq9UyybjD5JxiS2tQN+uu6iOzes
pbs/x4xO7JK/pJTWk1V8zmQGKSVa6FYGTEBTnimuSmp/NzS1GRojH9+yqSLuEHNL
KwzJEajVd6P18HZD+ggu/h5BjolgDRzF+2haVuidLTLrssCv5ynULxlVckvgWT29
/+IdY8MSXJl+ppD+zidbdUGz58O1ZsVodIzE4lyquW7VIJ5gTRRNNoZ63hdwWHHx
ANtFCDGHL82JoaKfXxAvE+9SKukOK4AEieYRGzb49AP4+kBq023vnMnXiQYCk0x+
X/arYDQeTxvoAGTpzWY05m6t7vkhyXjabrJ78qfLnBqwiSZy6DWRcpWmoIFYLqHR
uQr6ZiLANYPux+PlOwHucof1zwaujCoG6xqI5mxdi+lXRG+BSu6srXHIYN0v0bDA
7RdEyYkF1sZiYr79VQNdv6tsHK2xlaUBlhFrp1W58FU2LCfksmzsN7bBd1wKFeuv
0iG2LYOuzxMo2XMugsGdhLE0Gva4v6a7Igp+6cvkiJlvTMAZ5+sfDFgFSDfPxx2O
PTo5/8SzpA65hyAaP+AYDI4jvcp4C7kIrGvOe/1J8fI8qPtCBsFQ47b9sq5wbHLI
C/bknZrvoflNQQqlaO691oCQ5WNk0LywqeZhpLCL3K/tcRAIsPF30xLKGtYaS74F
kHSq3aBArSYyOV/qftN9fQX+IYiu0pCmI5PZqKXnGpcBHAX0UxJBjlxhHi0R2d8c
9igcIzGk2IWZJ0I16IX+7iKwjXZep/gV52Trzrf6hngy2lWICEUVhrcrHf3DGRcJ
M/oS9L1h9JDlFmc9Ul7QQKO73LHR0GXdrmkPmSpHU9A7o4CBXO+fzRbgUK3bSkc8
pehT8USC1QMGa6Bv6V4Wo460HOzZxEosPEK4KlrV01uDzU0C/Mjwkx9GVQdkgCWs
DfOz/5pbY+7uxd3mRSd/mRvM2aDIAIwWfKUnH+mtC5kXdV2OnvzEKkQQc7mWPjMf
M6UuPeUiRHtmJU/UaTs7Pa3t0WCUNciwgxeWNcl06Mp6HZrZxVIsuC4SbJg6VmPu
A7f8OqEpiKcVZ9SXceGJYMIvXhRCShJ4ZG7VCub48kG1/OuysKY7sBQi3TkGwVo1
3Yt6lCRqP70IrkD0MXzTWTT586W7ueM0mxunrtWCCljdqPBr9mZC0YiysW7AUoS0
DmS2Bc01EgN+uoLy5YfuldiJ75g0TViMZrN1bCUsEDX7mSVDdnrx9xavGJVO5Hvg
0nYcBGzOV/lhElfTxdxyjFkztgHpKRW8zpvXjcKqorCV4tth66PaWsHbkI+hzHa4
N7eRgipJdOLFVZwWFiSxit+I9WyB6M3o6E/y0SttlNdzI/KumFZnqYElAeEswA4n
HocHzzN0BA0UdrlAiZYeIutx3v+eoJp22KnVUSqGhR+eEb+bLoO5yHp9XmKoji6A
z4qiehtDYDftgWH2GGJopiSO7QLfrPQEcB1vSQOsZtRE0OvhAHT2OSm9LPdQXEzr
Y1ythTVVU0CcegfvCw8R18NH6uA9NdTZ62q0aWz1F3o5WSUcD48G+uPHwAE0mg18
ejzREN3eU2uWg7K4njr7M38rltbWVkrphFNYSQyKQSFsg6+sHvUjYRT38hkgAYGd
G0+dLXsvWwUb2vmvh1RY5652rtdhF83DuYWiEXyk4XQTeItrhGdm0U4Wl5YIOtUe
LYCo6PNaUfrKt3HQnoMq+P/VsxWgGe5IYXLtlz++trGCAcQ3tc9geBTM4xzw9Boi
JrAZEcQJVARUqMsUNBGQ1W/44N/GMY8CoAXnY4SXrzm6mctDu4VviP3dk5UWUz9y
FCHy98RpZmwnIBzGI2WUv7fbxtO1Z7UowEPIpAmtahWAgBHBM6XBasRGAICCR1jm
ZkAFQOkOyqpxNh6fn2IAh11pcz7cx2sx744MSlsRhQpqOvwKwVtAdVe5frGYISGq
tgATsu1gkFRBLYfpE6y0Z67Flheu1e7ntlW4DNMjzwlTW+tJ3JPAk62Wk0T/aGUZ
6qL+5Vb0dXrJC31c/KKaLxcLOhiH7N9TMTliby0scwFTz+fNAXj8rwPEQkdSVivy
DBac5Nke5EdXidhG2OnCdQ==
`protect end_protected