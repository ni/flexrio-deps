`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 55056 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRvqr1Wt3HGpZB2xHiQ13wU4siyl5kbTMtRk5PYcPSgHq
h0kAJTr1SeKcLUrJKvxAg9t5Z0fBfH+ePxKzmQ4wrfPNPQjIiVzlWheB9QYPJhr3
k9RgVCMX+CxAeURQUYwir+UOFjxYeqcFJvrp8ThuF/tB8rvWkQroCS14QRQ27hc4
GizUlR4OKUTUSitBH5e0O1n84llC/7z+gR6PZfp7+zB3uN5EjLWtUS2uoPRizwNw
Zq5lLs9Ii00EHrrDMw5UvfGs4czN46i0vUaEg0xUKaNhRDEMlJd/C/moRHMQXi58
ciGu87TJIJD02fRiHJUgyVnqBu5lEcfsBp9cfope99z4N3i44z3F3HHsMC9OECSh
jDBNGMrN/uTJBbt5icE+yo5vJoF27/1YFYJ/YLZqs0AnhikW+RCTZMmWxgqPdXeA
k0+zyyQZcg6W3wme4+MSK6moZsT7Fy8rQa7YEcYrRrg9729e+IwQuxmGtniS8LlL
e3jxm6nsWGqAz5fdcvn5G2oUGK+49bwKZ10Ki1DvzR/y+jQbfXko8N4T1m2uHcn5
Nkw05cBknCkHc7LqHFxB4XaFcwEx+aEu29MrcT+MeliMk1T0TDE2jsKhnWAyVMRi
klHhhCqObw4HwKTbBNqSKL66soF6QNhTb1D6SIp7TjdFd1ZxdzWDNTR5To0i6v2p
sxD2C8E6VxrZ0u9S45h8iv/rLbs0e4pVtk9p+E+shXlfOWUSOlfKpyKagF0P0+k0
xd6zPziW0FFpk6KzUPeR75crT/b52RKUML93OxsAMN6lKnFuWJfJomKejwFop0QW
XHVsqAyG97bsoHIZuJEMYCcxYrLtduZQv9JZypuaBMevIszDttyv78RKjLl8w8nB
1s2ARQoXmYP37non//Elkd/jV6VIExwHGumkHO83lTezeRMzH4B7rPfcFyQkVInG
5bSvv9xoiY4Jxj9LjzywZnFkSIuyCrB2c/dxH+zX84dyBDNute32sGTMxG8sOj2V
hQVdbF+8afx83Ld+1mGV+h3hjVJmRdFD2H7wUmncYNRZXWkBPa2WycwalWGXxhk2
XxvSI9b03qgwBacThK/MEBkexdU3/WFDq3sS7Rr9tblXK6rtcWs8U4ys0m24rStl
IyE0hn5hBpGi62n9frtNeJvkMa5eHzAQ4+z0aHbM8uJ8PV3l4ye3gzYJO2cN9+pY
Ut10JwrHzm5qoBWMou0AMoJ9+NbtkakOU+tJv80r9l7ZAfQu0xAk3oIz+1Gg5a2N
r9xKxSnrHxQCIP2k4Xi/5W3HcLKHHD9UZc5ZufjRt/dvc+JdiPbjswy7Mz1/91ZM
n8GFRy4z2AIP4Gwsdbf6jrQK3mBw2AEtz35dF8akHyBRIBh01+q8zZqIYt2zeuCX
XmFO5cKfqhdlacjNCeY534RV5LEwgd5XNt8HxJtVzqDNIjRtZ3HsUTz7pLeHAsVO
r07ITOBBZDZ/YBqkDrVnkPrldUcc6NbFWkE/jBWBcwKbPpsRFml/5gBHXUMEpwX5
cQkhGzsOhH+7HIqx5ixbRkWz5GbB38QGLV4zNIHZg+538g22quJ3kuMZpMTNJ3lf
jXXQwWH8fkj/4vJgDkKxQpsgdCwOTTmVdTdQCcr6hWpFz6V1D7Vdm1S8wZ1EZUXt
hyvySa+tLbDJKQSnDJonsPMkJSsSG8hPr4sRJJH+I/wBmGdM/9yHS54F6Us17zba
rOap8AuxJ3x8jX6iR8S4GP+q8JYv4DJZ66eFkmeqgdbTbL9UqR80UMotD34VbGG6
l+UEcMTnlb+uVIBTDgOS6mChoCHuLO+1vwcVXn0xStM9v8OfR5qlkqanDxuHdMlW
jNiPfq4YzipbHbsbxatXCHj7CE+5SdqVzv2uJv5yC6DLWgZLl1Gs+wYhbBGzfwvT
2aSY26s8RtLBd91jhPR9mFfkBDkOErGSEvaYxE7RI2Mgaw5+q93qma/7aXxMgbRU
tqLuopKn2D2kcBVNZp650ll2REo8p8vVbQ/5AzGTfazQZNRDFtEQx0hIXw5gkJOw
Z1ZXFROQEowO2M/claMfuUNaxqjepqVT3WMoq4QyuCs5Cy6jQDbRWaWmK/QmsPEp
LjheaH6rYd69hV18Jhv+mDePzjgxK9a6bQkQdqQuN9d7ovdE/DG7VRe4/gEyDxNp
j6f++n4w7mIIKnFRQO8HoIIPnbhOmsOilIes6f2Tk4jdJ1mktkXcNn9LqYk9oZ5/
fiGVV4Wyx3mefooE5+5HQdJ5+erx0lfv9gihghonf59QIoLLZoDuQk4uYJIsma4Z
q2/a74rdnU2/zV1h/CngYXU/qvuHfQw87lsFS3Bc3chQzOCvl/oz2n7PmukC7CGg
IP5RcOhSMJJnh+XS7kcxZJtEZg9r55bMS4pseedZEnBeEDXeRKEgfgctATo4IP0l
hL5M6cN9fvZMJr53GK8Qjr48w2PCqHDGCdQ4PtNF4x/3AWaSQAqdUxx096YB8gEM
Aq286XNYhqubCeHgj9740/e94P80fAartnlkyxeY6mkST5VxCWzPQELSm1O/aHtC
M86u2houDToNgFDxMwzzymbAtF+5nzqrcjio0VnoAHRUHtbx1n4MIARp3kipvdyW
oEDfZAZTUxh3c7eHgDt0ZVxOe2m5f9D+1upIWhUMdSCmznM4KoU0lr/eETnw6lJA
zIuGeFVeZyAkYc9b8n2fXmsfLrcvhic55Uvk/fUxC3D7XGfhs0o98CdX+oJW2HME
eRFSeft6XAP/2qVchw2S4nEWFzHVfKuvnRKzzjy9ZPVtPu8JiSScpDKfzF3GXmfR
Kv1LLZ/8XAnX5ly0zvhmbv0uX47Z4j6/xpskEzozJcmRC1YLyVdROhETZOqKklPs
yg3Pvsg1nWyzoDBZ0aHxg/8vmSQ05fuwb19ZH4RhxrTWB9uSA5xrW6cn0wYIuxzm
GO/jaRAfE1+ScAPH6SfCqharpatxu/hqhnSiZhGspemHRes+op8WwcCOdytnYSRq
V9EW/4l/1sf96+oV7CgLZHuzWQBW16cEGkssT90NZNGLLP0RF5gcGWBRTAy/KJw+
cq7jkTzInJQnW5MM4GXzj9zBNXu2v18tB9fsX7JlocTsAiKipx1TJLjbAO71EA47
r9M9r6DoMfzJ5mzx2wD7JZEdktrwb0cEXae+ccgMK1Wj5Qlgu3d69H+mNoEgsQoc
qvUUiNpD7f1nnBIhPZgaR8+U+fuJT7hIhKHrWKUcmTIYXNTJ0POOJxN/d4ulkei2
WPkCGIsWhZec6vuCv4fqvazfe9+E14fwVUFg9t49UVqlMB1fLx93e+zwZbiBFT4A
MeTGYn+mzyHpowGbzUv9xZU6JUhvdi9XGGnDvX6ngG+sOzKdJkpVdX4uSGEUSu1V
pKSRd+rpd5AIfvgdt1jocXwkPuy632EtmE+0AZghLo+IYSbgx6JnVEnFcqyf5GXk
SXvtO4jo0lVTxgjgO8hLy4BwPsVVvrQBMAHzTxrAiLHEdF5hgqAjaHszXRMpaDOS
M1At7iq1dBhuo9kFSTzqlYl6ehH7QKv/ZC/AmsoiMhXc//vFE0U+LuOaeok5Gyt6
xCDlVU3bg3jcPSPmheybHJkjxMZ9y9x4Ymj30rAN4WfJRculS0FbpMPnF2PTxil/
AfR5J+oTBXqWxCh24Z5c4lUdU4Zz4XVcJeqWCytah8ibdXSFAYQ5mkKkJujSt5d3
QyazyXbl4CgSxIZAaVwciJHwGVP1UiLL2ZW4mbStK7TkQyeqm6mWOL3KMQw/t3x3
Ztv0NgN5LJWzOt26zmbNV5tA//0MzMI2H9HXepsguVdjXRwB+J6RJwgmqZfskIV2
+5tg4KGdf83xhbJ5afIxnM6CXm2hY8a+EtO/JrG7isOMIMIP9z6DZBWzu5fD+Ko1
BFyI0WzxTvBViM52ASz6ufffI0sobb7dEQov7FX07Jym1Ct8Dcw9iWZOXGsm7f1c
58WnCTOXNaZPSg+S2bQKdQFwRcdM0Cfn5HpnCZRmVvs6gpwHSS8fvbxSB566hUWH
36n/T7m7D38KDKgvWmEG10TOHRp+SoZGTzXi7vqEzPC16KCoELy6EnFS+8GrKJ0p
UAzv1hcW5NFgc9BJXiaE4Xxmqwvypq4E0zJ0R1MuihxaLFhQKjdcektJVBAuI56l
59XwSnSneYF+6cSeQomf/UlQGq3aEjmRjuUfnPxy8lFASb7qo243HdxAEf41x3Pb
Ca+u6ONzh0DC8+vqQ5lTIZziygMU8XWFS3cAflK7AsgGoWuMwA7MQtCcIovfNlTw
OXohu1PTLgANHTzyDH6PSACFX08Pjvt4N8pOodyy3S0u2PJf8AJgb/q5gCVzZ17S
h4iU8OCcbqSza+5ckaS4vCYUgoLczzKNZggS3saX2YWYkubw9KUuyV43kv1n8uc6
RHHrTmJNxXNGgchGhUHSKvOqAoBZhT3+gBeh5KWFOIR012dXqagAXY0rW2PBnz8k
2N0Fp1KbFZYAbONrWtiYjDXLtrmWzk2ymyW8+It65vmuN6dF6fBknf2Pp4DPlmEk
oB9raEIVxdSYhC+mcwQeWRiJJI/CdntS0kzC0z18MqFOkCJeB5XwmTH9oUOtW1Hz
qo+EpxkaToXPWJcSZeyRQbVhPGGyrVpoye1AmtR1zfH/DHkbd6eghTrpJPWb5O32
ebQKuQKO+zFCCAbpGxSSVqAO6ZuXzJrebLyiXYl1bAl8G07abbSCMp2XGS52Gw6a
HHBvlmRu/PBcnDZY8OvINf3PMldcDPh69U1BRcwx8/zFJh16Oo0ZpSYiOZKBrVOP
plt6BtQOcaBjGpMXG9JVcufuBwwVBPs4V5K8f1w70cNnNzOk/82H0U12PwjuzeK6
UIrzH7OawEcSE2cvXV7K/srAyendAWjcKqiD6DhlX4UO683ZUQ5HLmlf5nmIOMzi
X9sZRXIrxt9qz2l807ClNaOLgf5oFoDLQXW6xzujqdgryY8oMID7NQvIexll09GB
QLXQeg77u3I5+0EjMmYdx1xPhblwsyCL9YkjSHYgCREEb5QQRoqAIIUOBlOdBs/J
ZR6/HSznCyFO0HgBS3pcZLb8GbKdjEa6MnoqKWMDqXHd/v78HWeeV31oU+o8hILf
+aPpoUWJNgm0BrsmgGUpzSzvbNjD08bNr0NhJ6L70U8tFz/4bAxl3fsCIziKQOVD
DTgjKCwwh+38D269nRHQ8hdFtdWmucToJNbG5ZWp0wkHRSO9Oe4suKt/YbCdhuc5
zPVxRtd6zDX0X5uZiNzcD3Abgv+ChCMZP8XXPhnavqLdy1E9idrbVNwEHlYE5Orl
E/VOUsPbjw08mo41w5E7qDTN7b7yqadjm+E6yo37cx/o3LW2IRD1N3z8tvYzZTjj
hOrTj/UB9wk6v0dw4tlBJhKwvPJo9i/EsK8cUXcs0wEOzcp70dwD6eiy33ymKj8T
HtpBVceS0iCFf0a75hbCD0vy8mohbKE4tdJjCDIDMlMi+Z3kt7wmeUyJucfumSgU
yLO3gbv00Yb/riEMYtLijbnyI6YK3Y9kAk5PZ/cXVcsoOD0SxT8We6LvNkx9ZeIl
2bY5n4VL4tVJW/K6Bh1AyI2dZNsrVJiHh0Tn8ZzbBH9D80a32NX0RszDYSmgPx/W
4uIiBQHXbpgdr7F7N4btxEx6JwmwZAA2O8jWsssuMNmG0x+Zh9p5SIXQDcsvKOrn
toE1YOpx1sdoqCLPBG4S0Y9WDK6YKchY6oE4Iv2Y82hrPnaGr2Q9R4Qa7ZQIVEAC
P/1K8GlxueI0OfVD1DJQZekCHL225XSfboo17x/XcIcDHVHaXULtt18KbXcR/1C2
vsVKPZS4OmJVxuStsd1873inhvcUkCq6NXiPu2ak534m4ZOIO9mH95OlTpYENAXm
NVTJyEDe7vYwHQndIRuLU44iK5QbT6EH6D5EN9yyiy7hm1tSkGxB7zFDbYjcy+pd
VZxj6X6VxYYpqXgoCt7XDhzgAcGJ0H3ssaKdu/x0g258Z32nBE+c4Hhkv39BcZ9f
1UZtaiU+32+Vrx4iSQ4lI3wRM2uN93nusTMWxmOcvIucicdyw0Xn4wf3zpLGWdGR
NZ2tOGVx4pyOvYI+09Mq1X0beDIbPwWxBecd/QERr95gYxJUfBORX07FQ8O7wIJH
hNJGrXl5YN5Ijv8iBEAtVWDQw04i5MaR6qok98Xub8smHpmp9EKCRUE25wF0IHYs
RPB7wYtABab6tZrn3UMcl/j2hnEqEv0+RbM3XCZn8NQMtSFfFpmaAPspxJVIHSIK
ufSwYwYIKv+LAYB1FIRdBxVxwUH6YXeere8YH4E8ErwIfhVyfqCWGO7yP9fbEfAP
e+09fu3sehWJIZz8ZbcGLZl0DzXnXbNTAplDZ3f4UFavLJ7DwAYkFuF8CO8pJGDK
stWM/e6V2DL/Yj7ReHYZuLW7PBpdCLM00yxppBA1AEHqh+PTOxuUpDMHGqhICjU9
6LzscYCnyU5nECz1X9VUpu/DF1xHRFxcFOrA/WJcmInHk2gjYovHscgMfGYZidXE
qdjO+QTgw4Lc/Mtlf9oKFxo9/V3yk0T6GlJdOLdLrUkR13QYaBRXi4ZH0j/rwyhC
Obh8OnyifT1PXG9as6dBF0aLFhoepJTwnYOboHBmV6e8FY8Duacj24Xn2SyGUOw+
W2REi0hIUHN/ScX6HjcGnA+hN8tMjQXCXkEKscSwUeA7ogYkxKLF5i0bAOtroKZ1
EqxNxCUEuQKh+PRqxLNXHBjvd/qSjGHj6JBbiQaPnvb9ftt8qgF9+sFO6TaFK6xC
/Se6TxzRxIotN58rCTd/BB/ua0jjhBbNrqXHony7wDINSl5yBy0V5II6pRYJoM26
umY9T1ySK3M4+p0rF2vOn8Lc9NTyODC61CrDGtvD2Ld1aciVZeGeDX0M62vu8tx6
t07uzeCPUD/QQ1zVysBgu/pQkCRPZ83ZuxiU22KnoSDcrcute4Xh/1vglyg68lBW
vlkK4Jgbdnxl428xDmo9ovnMiPribwkk7lo3Iz9hPw+HhFkTzKOL6zSNdSFyMFQv
4Mg6Ild5P/GK8Jj/IOWQFlVbGAS9JsiOuTjvR+rjgvgeY9ZIj5GmCs8rT66Stg3F
3xcxwZkuvcmsDWPEB6qkbX86y7nJQXED7U+1ztPZORuXgiMRs1s+ZStneWFH3iiG
e/wRBRXYoVqpO5CDP0O5GPTCn79qoi7Dpcm9rgVpVcH5nbFaXtDE/N5QKo+MAvAo
hRcxHLEUXKUuL06Ny9Tnnl10Eq3z3nB+LjxBMGoPqljQY6mv89DE4DlayQ0B5Ghi
oa3PbmfmkFC8KJ3yjlO10I6MF5kaw28N1GGLe6iYeV04C4OkD0oFw/btGOkIrXIj
P+Y754KuNp2VPFHq99cxtN18qGt2YQbMhe4DIgY/T6VnrHUQoXhwkfCTTRXYtqDN
udgWCcnGgTfoWA/R36fLsl+PeGfRcl1o2xDN+fOd3J6rQyQJXxWSj3A6nLZu8sWQ
acCxEy5idbd6y9ssxY+jwG3DF/DzxGfoBZqbNWBneAdaIDOCOlgFzcISN86xhz+5
12+CFstHUNv2BvZnVr1sginz32SWi4LQQTG8u8UiB+5LCHtaY16RJKwiXabzchq5
PjkgpKGQhHcdjQIFsRokHsfulv1SPomw/0PUi8gP0Im2T4voGWSGow61QnJgntyY
QKU9g4B6rhYgbdEtQHgWvF4THSVMW5tL+CO0YRXiXRhlFRh6Z5mBKVNsHM0tqwWZ
+whaLp4Ygse/7Nf6EOz5Z5cV4YWvVmpwE/YvaXBrrVsLPYyDGcK5ms6j2A1V60nJ
eldOMBSPP8s7rGZPO6po1Yb2cIOQFKUdbPOLQ6ygcVH3MtksELT9DDrVbY/uZx8R
n+ugLhsq0kdWC3DI6SWievnoYWuPFyjeOhyDKwQqIshUsuf26PV5aWg9h24P7ZkO
gdD8ZV/sp+puCnblt4c1P8SOEkdoMXDVxVp8t5nRXgLABg8viEmAYlzxmMqd99hp
mj3Lw59lj62gA0p5JG23ahX2U+Gp3Zws1KeDJ9McFxm4rS4UgAUhKar6WmICC4Fg
UDYxUqqqfp3V2DKg/dmit9h7SIsig1KKtCes+bsjBiT7ZjV3eLV+/0YwwrC0S4Sf
mN/+Ecp9aRYIp0J06ZuXkZKsxTLXe/HznI15DNN8ujgzSiobEE1YSVTF0t6KgKN1
0GiujSunb76qK9tUgXmwyY4ksgy6FgMvdRcY05Hjg0crHr4xbPF14f25Ba2i2aPA
/cJG/FrH/MfG2BJqOeGjG7EULsnL18z01gOCIkxIHrOI9kFd7Oq6zZsKNNfPyYU4
KqDT47WqyW5i8KkQ+jD9ObKaPkG9+su6i8NJgMWLYp3l1aPaOW149wyJvd6nfu4k
upS9Yt1Jf1HmxF3J+9byPBcb/0oq1Rzm5i7iTFVcrBG/2S3tp4DVOBqdsokOzUdP
ArbBNy2cBXgDfH9CJSrccuUD3uyQ1X54t3c+pmO8JjFUe7/E/OZV8mV/Yg9HMpgY
wS2TCYi8Ok+ZScO59saif1vsu3x4basnAG0rmM49liMfD+M+DE4fh3MNrzYWTmin
ak31gSvEI9Y/tRlwU0hKoN49SKgOs0uLI8DUUZ6rc41XL/ZmVCS+Z1RcUx8YHF4n
zCpue7kKl6DuiN/EJvUNIEg14XBiREuRn7g7n26eOlC5b2DwWMo+fKu1vRtSCbd4
eiGFaRc+8JThIRr54UyrqbVMujG7BBolX4Rqv5YzAKBF6V8loQmcZ1HLQzprlZf4
dMVkUvqjGXo5RoIVvtHg6G0+OaPzEBomLrCkoFJbuejiGe16mK2GN21J81jLa5dS
biPh4s/8SgzEtA6430RNMNJuUQ5TI4/aNKVJcD7+8HrZ2Ffl7HlFUZjQq8IZwh/R
eKiEOByKfOKjwKVhAe5mGCDNQ4rED5NGzSbx3NazukIEqB8aoMEWMTlO/Y282vL9
NoTl85ooi2dbMNyRuCd7I/7I0ztvjRImbcdz0952BOzPK4F2lhwqEAhHnIbUs6jR
dkZ+Y82s+IrQsXwjQlxey2XPEW2P7lQuCzpgBXKLP/0AgHPf50ABWHLIb+dCGDvN
CG0wWuk3SnStdNg/7dX6dRY9MLxC3Bdxn1QtZa4Puabqcd7PTGagXCkf9hLvmrx7
r5nkraqXrxKdaq1mNr5UAB7KFbEnjq37MozCXxs1B38GCQ3BMTA/M+8+7pd9nQiA
MxA4Vm5sn6uwquCBs9ImJ4vT6FTfSjy/hfr8zt8ir0OJ7ufywWE2eOOFTeHrWHis
HjvcFe0A51jkPYTWc0NnE0pDLUP3zpsklabs55w7e1mQpuVUzvX+qnwFcigUlNAb
NSm9UWXlRCnw0HeW38KWdxH1xiQ1kKIV4uGWpS+gP7VdJOnznKAG375P40yxFVpY
9UvrldFPKPSXZrTCVt9Urmewlmfs5+SQg8tu3Q4WVyC4EfnKaq00FwiBlsfawit6
kIDiXXdOk36zrJ9BlOZ0Saw2SRVEQeY/T7B3JJi5FHjqfjDEqTVwLv7N4gRk8U4j
bxNWEB75NOiAxqhNWTX3iRp8kgcIxWtgABiPbGSRAiVGjeIfFmNiZSe7iIc31Yj1
1df41zCFzxoec2+twFDRq8IQyzOcHOiCrQfOPTFboBjDUfUp0Q6d0FlRRp6Nbd0z
cSpiRqBOVsqpSdL6ilAKUkxVl068V3EN4FzKDBVasQ15pwKOWwQmE+uztc3fmxVe
xsnm0xYO+j2uKFuaIusEPzqpNqHUj18B7WNythEYoMkDzuR0iLj15r8uZGT6iGq2
R3RsOnrBxMQpV3SiRHmN9cEY/BJdlBkCGjYOiRZkkTzLRiRwhwSNLCQgKeyN22Uh
9BbXSvFxrcmNFCt9leRK2AH1CIrBCC6I2+vnRvw7qTsCh2aCDX6b/B4/Z/MlE1C6
L7xHqPYSAtM3Cw1e0ol4OvQa0zLKzw6gyvxIjrrDvjNTbQ8TFvKlMNKZxbtm+tNS
d6HbMWUcU9s3yaQG+IKL1Mqc9+BOfC7kfxJU6of7XUWtpMYIysseSxQk8Wf2kqNr
bAhVmrj7fv6LPpkYWeciv7C1KW5Cp8XbZj/4lRlo2PJGCHSynvdjkiCpyY3sB0P5
I1mag8NJ6P5YLKPNqE8M6GvlFmNTx2CVzMn4YTB3E7c9cv4eJ1MP14Yb/J5szohj
TMoL7GsXhbvyWNpPIeoXD0X4jl/hGmr7C/2tgA2+Q9b4X6QR7R7fkbV86Euk8n8H
IfgGnpuyMLqIV88a/9eCF5zh5JpATTDY68lEhV6pfyUdJ5BYXG9QlNclDqrVMpks
BBx/XcrFoEBXvmxG8is5k1SwYX2sFxhJ78UNU0gLa11MxwfO208d2TIbXENNskA2
aYK+0Kx+1RNjaceTqDg8a0jH2pV95eYSqxpHkEKeC8mGoWdJMpPBGRfsYEKkhl3Z
4pWew1eq6/8GvHJkrE6bGwhI996ysbY2S+H4LiyXiQbsiDyradf1Z08QLjA2KRJD
TjHQvN4JvcHmOTQ5hhl+w6Mp3+wt3PeLJp++4TmZyZmzXm/NKz5MLKmf4tIHzEEs
d+wbJXv0+J1isZsKqH6/mF4mFDbP/OIRkEXSGt1iiYwIZZ7k707ojGMBMPH4Q6wF
T1vwUClh1u8J46V5nXIlYjCX3whh8SjDxugyrnmytz2/YB3vQZNZrguHqMsD53ma
56TPk4VZ/PEQgIE30HVrV2K6oKjXTyXx0Ew7rMW8Jp5p/lRYq7f7mZR+8zvqoGW8
omOewQEqy4QfphPYWjyEkIDEe2zMIscKhwRbh7lNVLF2k44dIbZ2V9+e56xzAZPx
RbokzZnA4t/QtrfwN0kYQyjf36FyjtJMSc27mA+VDPUKJbEnQ1M9rhgu+ogU90dE
CeifMOY+zT4W3LZ8jygpPFB6KT1GL5nCH17/Ecp9M3QXS+AodtVC9BccUgRixDpX
+9p/jgLOSlW2t6HE1QYgt2h0AdsjPcQEMEbH51Zp9NLI1fc/5NRJtmTPS/bbjVQx
EZUQe7Gp04LpdqU3mAzZf2xU1e1tRpP88VAh/1PuQo7CW+5+pI3rpkulgm47F6TA
eq0ee8dU5lcaFi6b2MifwXGQ/hcvwzznyJQE4qTrGDK759WDYuslhoEpNGXoi0Ns
9egY0cMAM+BkGJC62QMQq+xGX+7dpDZRXZOy67kqXNwSgXNTsgIB8h1b7Ek/NRK1
L/fHdse6WmrjMlLPAaKVBJpPlqOn1W5atWvBIDT0RZ8AybFUsOMqzqIEiC8kk0st
7FyAkPJOAnGD+IlOJbEyexqWvf9TVJlG1Trg52ZdvahxTK/9yYbqb9UbKw/TU7uj
5/B82CJ1qw6YbpreDljqNYEA0Z3u1+oo1OIAeyK9d3afPIUOJEUEe7Q9jMyIjCQp
P5skNust2EG/xccF6SxRQVHdT4losr0JbpniF3/UzjpOj7WiHPHtHd8rPozw8Hxr
4+BY+W/sT/twmDYca8Z4OgEKK1snLfv6a4ItevP7oDqIQ4Avl4BtHl0bgP/vkock
RS9bOycGtbWF3z/MW9BTlQjJKAFkH8rZbBRHdFkVXQ0Mn+3BqtLWokRbeVLw2WAm
EguL3/2w8zMfuzajCwos5h7eCVstPfSqH3t+z5KSAyzGYb+tvK2ViOofKt3aUhTG
+Fetl81480rVZL/XRb/+/DW8+PMII+zdvtsVZEtgEa2svQteMRFWm46xuqjNo6Pd
PhVUParBRYMjIObLdBiH9yrtBdPS0NRb0cEI3+TufClYGdXrsP+rJZu6idy72iYc
3okz7rwMX0UlccsqNXLGM2dCMfttIm90y7O1DNL1ydST4dVSYlCkjxHCFd17Z1My
FNqxRydzZPFINcdJY6+595VGKWZR53/jhecEua7xmMKyU50kYtaEX3CYDDd8EZus
lfmSu5Ia8lLp188X2disNDvrosh7I54B87qbBfBZ/jZCXVcq+vXtHNdUQ2BxIW1n
Ow9saqJpG3RzuXMf4hHDKRrrvCp1RJ8J8ZGNPEjR5YZLglGhCS3gckxMhqMJ+JqM
z1vl6z038b2f1TQ2LlrhiNKb8mCixWlFetNoJ/0Kh8DTGtpYyrPn1tMarCRhajLR
1a5GTzZ2wFA5ZVyYu2YGS11p3D/BwYd0jFl/XOkAoNj6o7f16nr0KuBn+Q731BwF
H+5wlvwBC0L5ChPFOMkW2yWmuGyw+FpWocd0X5fb3+I1EKsKwPd1KJ+OFadG64XO
MFcmNCiey3PlkQoaTOyAkuUIeHT1zt+faGtib3oCLXaUhcLfPxKLvqATIXUMsdvR
uqScbz0Cq0fzVjKHPZDONL2q41gvMSJ2ua7VGfJQfGRFcxRf4S72OPVtrrNNvJjz
I9LlVG/x5yal/Hys6FVc6hGC8yv0wmCMz9wFo30X2KQIcsNZzu0T/DG1bD+nMUca
DQeFnZ+ACjkq/Fe+Z7wTyHddO8xtM25vc+76+Y6m6QHWExMvDJKT/indHihzN97f
NR+h8hfTNTcBbnYAzrxjeHiqo5s+6WzUae3fWvlf6IoUHrzoBUEh0BWgiXBaYXKn
IC7rOEmAXwfbcdXG2owYny7c04u0UF5psaTgRArshgifUEsxf22S2fp/NUpmTEg2
XDkjBQmfHU1kPpkSwfccUmSQUfQZJA44Mbv3CnS0kawMPbCucP/i6IcVc2xAago+
P+G6q7R50anq6B+8HEVTFSchVKxVPQ4vrPcFWGwtLEPp315viLsvEvphgjImY3hT
a28/4Lj7UQBBjR2sTLQnIssmoOV3Wpc1ESXsGCw/BGwdaxk0SeiokCBeSQkQzdsP
0walYDj+cEqMbtMwyFNAu2V98mVnD6Bm89O0ZnZhmB7g4ZFhSBi0lqxb/gg2qIyb
QtSmN6B75aM2OTakjLYgaLswBHdygmQ4V4Er37iR0Le9MSv16BuWniDGxUUz/wPj
5bPg8Wz/CLtIXayCXRCknAXDR7/Jm76bWgPHtIFPn42Dt5fMPZigOZdyZZPE3xHA
MM1tc7rPBVK+xZSLufJbGWi670ZwmG833z+TX9iU2CDmdbq4AS1S0CWGTBxVI9Pi
IjKcqyVsF1k5VBrtVUNTK9jHM6zx/r7sWCNUwx7QmOgiPR5AkPnG3mlVnJqNImY3
jg7c4SnlVsUeHDI54mvlt3RBV9sDIOEAHqfX7y+5lGdZGqMbnIYoOX3ihBVUKHGU
zHcJWQLEMGRpI78ZHwUSDlFpB/xeNcn7Egd+GHBBOPYpmSGf/0wYKoDtN6Gs8MrT
Jkfp06sBdaVCZJosiEIXIa6SyClB9HgWsrut0Vl59aVFsf6RBLVlBsslsSoVO+dk
5C2SKDyTfW4F65fMgpAHIzQ2gIPXE5torC8gCPL9aWI9tTqo+HJ+GxAvW4yxL93E
6f9wRyfDRa7oiFOqS3e78MczInDx7gX/EOvw7LdahA9sntyLhPRrk9TdrrTRW3as
wJ/naScVV71XK96J2NQ5zMSJAZbG3U0Ar6Zqs0v6Qxm2CRWkPiR2rvLjio3sgprJ
9h3wIVsJS53csrh5GFvygS4243e9dkPt39HHcaNOCgrTg6P1cFDn9+HXpepZwgOU
YEJz1i4OcGmeiV2cPIo/Iy5vr4jbeGfxmlH/JjEvilE32LHxhoBa4GoY0dn2NBUo
7QQ3UVIkuflHb1qCwbaVcNGLlj7lRmJXvfw5P+xNLd6YXVrHYIPQFFVi4xoKR37e
OK7W2yJvP5v4PmA5DHenYy7emGwYoclh1+PkFA0hg66b09JhI8+FAe4p0n25H6r7
9NYSAeDUEsxAmsRhJqBjDGWHLJjRSPwR+oL0cZ1orW4mMIyF1bqxMyKe9S7mHE2l
pGk/MgJzr85q7Fj5uSraU6ZjCE/DsUaDcSmRoxaLvF6CbSxuoEXVnXCXFCPh57oY
ZRoG0NOKUY7qcTdgPzxWrDnyOKmnnjWN8h5K6KjAEch2tVt/nE2fyEgxiycsNuDZ
lPx5CODsNbEawMoqU+TxiLD3DtjrMdok3DncrnPAuT/doj+Y0+8ufnh2r+bn515V
/aR30MhpeYzX8oGxyZqJIwN7su0Gf6v78GY2rl2clhlYajx4avc4lFqJOG5y67/I
ihy++rKPmQ0Euwwx0QxpFZ/D7NE803FFdM0xyHgMSX/1maTMBHS27Rx1PQk0EO7f
1cp7hIV2o7PrPPtq+LA22Kd6c+kMbIOcl61DQTp7I6pra89guxTfu1KbQFQPnnM6
MU8akAHsfgQg7xkow0GecktJ/nDDfws+zQf8QFQODDME5AcnQy6We+kf/fkuAnxg
yZaqYxhmFwVxAOVM85ok+ugLjFQ6dgnPVGFZP3EUW391A5sIruQ4VUI3ekjdxTKl
W8UjkE9madG/8FsPADxc6R3JjmQq2PJFz5uoPBt0DIXqKFCidDYPJRyR/TIg8jtb
Vr4XImOe6zzm/XSPuCgcUCQWyVcWdRb0dcaR4HVb6lEM7fnEKE2ZG47k3jVzGFMD
qzv8ShNvDPuuyeqGmgc8T2s4BcztVDMJhP7sCKKvPQWjQlMOPuElm2AFXQaVgBzU
qttTGC/z38HW9Hug4CP4Os0ftEZXWrSTu0ndL4mhQ9+FJLUWlnD2gOuYxbD0v3p/
WZtySf+MJrG71kQ/wLkAB6GWiydcLEtc6YAUdizeVSpA/D7EpulduUfQ1VN/XVSf
tT3MjvEv1FbAJILSbv+sILlq1woQSGAcjo/5gl0Jh3c/fP0i+ZdS5wusl3zqGHZD
WBBEXItgu8Tixj3+XzAjvWjzAx8Ws0sPrB1HaLbEgcOmaAiMXwUyULYF7lOPpDbm
3F6Iz9ykWT47iQICI29DLLZJQ1MaH3rbIKYsoBRz8H4jpDK96wYfvE4NTyytS4di
FXLAsbxu3KSBUsL6SjHpl+bCrj8PLdQtPFIC83VqcChMKFR8gf6N6rHVEnt0ciPe
juJ1BiJJWfVclQc582FgYqkGD4v/UPGxXukXPNJYJPPaiTxzU/Wn6uLe39uLBiDO
kpL/3CM7B9Z1pnL5K2N87yvfRHoEcdiPxe5Rro53wOENEPLLJy1JHF5ZWt/WwWp+
rUwTT5dAdnOz+0Ivh2ns3d9gLj+9SKaH8lho0wdNoBOzAZ44oNTXy9GBULvCfJBt
B5Hrbdm5Be49puELaXANRXA814X+YNyjgXKF2KK2B0LVPipFDcrXgmAyCxU7PXOm
9ECOPk1Qhv/aJHFFddFTj5xN+HhHupifuBjEiYo1wlWG3felfMor6CEBAHaXJh7b
4MUmD/nvs5WmLqMSdDK4FMzZRX9Y+yNcwz2lcVfmr0QBzRl5dRAR3xcQMAPdjZgm
JGb2CdDgg0FVTN6t2GBaFjHSiGY8owfmtsIT5ga7XpfnRiEJRzp4W+fLkSeyK1ej
0qzR4Z6WwxwiN0ww9+ESbcV73F20ik3rjIHMM62iU132JSxc1LG+v6wHZ5uXAbIG
/HeSxpUMslIHfksVw9mHcA8kuS3MNVouzkFawdovDKPjW9qAB3kSrqbtu0Um5skU
/vxJbEuZM4ZoWJtulclrRIxUgpwVww+DxjBqg9dnEPc7AZv7q1UwEqj1WnsDdl5C
obNJwvtg3HiCngKEOvq2jzSblcr0MzSpytQQZjalC7cFNzBYOr6yA5q1zTp+wJYb
2jG5t5xRdnENdJG8ByB2WFNEqUprGxGnbPb9HWmkLqxdBtWgDsbxMsb+XVfhRotY
0idHXC/dwwmw9SVS0C/UltUAYhbzv6RM3vDQOt/mpkjaK6o0+Tw2ZrPEdzqpeAlk
GnI46UBahxK/TObVRURYVhe0BA5JflemnOhGX5kMNbEMBm+7JsabEGww9mK6t+5y
xs2EtoAAv0FRG+nHDiInn7t/wQNxykGU7pM6rNXXyX9KHqmofM1INGpGTnutquSZ
nOv6OvQw5r628ZdGcF2uDdxnrTQcubHaUUS52vLaUw/zMecx6kxr0Qs9/hNzCabi
toUPGB+8KF1gJKJqIHG0RTmsZ3nDA5S+3i49Nj4sS/O3Fad2+XocpMpY+UwcjVxM
zj07sC74nbIdPRMG9m8rxGsR4wGFwpE28Bg5Zw7Ax2qDuBVa47ZM6iWkQUE+kL2W
bRb5CBhDluEonMZQAvl5yCyvaxOa0xKMspR+pKwjfDcD0UbampaThqiEqBZZ5xP1
q2yjcjtorpedOmQJrVj4vuByXsb9mXpxZrriJBka/+Ysm0Y4SPxUBbfwPvFJDHp1
PAPftNT0dfJxkZ0RO301fptqhwONZmznTmbfjYp4xIuJN7OmJ2mVPEyrekWTtNt1
h+aTunsZffFW1hoBXFtEtC8z7bKc6vPLQ6iv9bLL6FBWA7iJW+MninjRrNndt+7T
l0rBDrOqebuHtnv4RMWXpkufW6bdvW+eWDLga657I7t9EeGlWeIqfzNAEjn1djQM
CCtPzFj3OXjNy5IVsUWJljTPSWQahkK20oYAcjd05sD7wJ4/KQ6+YKgxMa/94oMo
kBjR2GsvRGaSlzYotg0LjuoD7AlwbMwW2NCkSH0Erg72eLAyWFxWAqKY3QNPPBzr
XpYap/309gx4bsM8mJTgDUdmvol2Iyca6uO5t5aafXafg55Ojrr3KW+9DYK7d/zp
80dOs7FzCArhi6BJKnr3OOQvAlHX2+E5qQ4DsmIpCXgKjJf3qOKTfbD6GK5MvL0u
T9wRiHkn4RO5RrfxFTBV6avxwX/ZPfsFtFZF4dRcqT06T7FTJfXOSPvVKECbJ7fC
QWzPjni02HNLmvZ+sfarZ8jdYqoiR0j12Y/2b8LFjY/8y6Vaz0CReZi+NPHIH0L8
Cz2yIA2YEDtWirkRgLe15jNX8y3LmVRvc09BKd5078R8TfE9DsJ6xaUODt1OYMF3
oOZgd6LfTT1jpmzA9t+5p6TDQK1aH0n+PN4b/g72S6wGT5RfnaXzjdHpXaXa+4bO
OA/jTMHblpa/A/OlBf15qN8L4boyh3BehPzaORvibYoT5AgasSUl+z451iyeVk41
8WumDNf5r5UpZm4XgQ81sEBXndPlV4WNFmRPnwOYr2nKeyF3wnw0GSZEMxmB1RZb
7cRrb+ccC0n3GaGE+fb2RGGSAo+nACGt4DJlOsXb9bs2MUZAxM4pFjMsO2LCABHN
7Xv2XLyDMGzYCQ7eb+6mFspIoZYR/MDtXBUFaYvUb4AFtYaRkooT68OxNeJhC10Y
mcEVoAePFlws2bX2s4qSJsb8gLkBvdxAfNJTkCFqo142A9YSDDpu4H/2wyTD2f+j
WnFuwKJUnR90UoV5fr6GacZuTHRyR8rDk/ejL0MIVYndmk0LvpotQ6zm6cs/Rxv9
vKsOgiI/jf7k63qO2EZuFqqcG+ZNzvaHyPeslKo5wiLPsFyZQpA/d5EuvwGyZm6T
i/xvDiT4IryzwpvV00XtDHpiLmiqh/MYm7tTFYt6Lt5Q+fhrJwFmjSk9/qeyrHWv
luR9uZL7WRNdiYkc/N1uqEyQ87oWKJUXEPou2OpGVzjHXSRTJJSdL2cX8HtiM4Vc
uV1RneGYqwf30ygogTjbPyJGPB2CeWNOGJLuonTJHfiGgzQvqG0I8ga19R4kQgeh
5LG8ZJGF59ZNngFZ0pxTY6/cw+oGnheLCh9lhaxqK+2eK5K3oJW7Daup+DVkkxaQ
7GIFoWQ1bfFrURIb9/JmB4bPDHPxw5umWMTIlqovu7ljvKUi8Xv+DTcBMiposQ/y
yY30c+jVXRn7do3e0DkoSTi/Qll9YBrAyO2JgqPzClneoksKAWw3Rs3cJyA1ogIN
QHE5AZ10UiNzaAlBSQ8Q8oo2VG6ZqFQ++z4oxfmyNXvIIdHcV598RqamhZlElKQA
1zl6jRc5NTSvVXKuYHid3+h3obRrETj7BRNzd5ms91IWJ+EGNRneM1TBB+VxqPR4
r4/0YYpKAs2YNDUnv9exVv9pGRuUYhptzMafMmyi6qUCTm+CHwVmcjzqjhLp5bBg
PQzC8dA0Zy1XTUU8ohAGesYX3tS4cv8PApGv1c6hhfrfYBziPJq8PuNVtdNg8eN9
0hLve35OvwSFVzgylw8IRswnx8SYngh6UYfFata7BILh72NYwqtSFtXXop4xqiX9
D3TegG0/GMnDb7slGKWx1AYF0BD9s8dY3fp2tKosoC35wSbbnYAQo5a/wgHMBkNj
KqWzYuNQKhzbjGPc5rG4dtqF0zRQHZYDR0g+EzDgwJGyT62WhW2w8STksmZyUOCP
VrTyy6cHXVD47aQTE7iLvEX1s2LfnzcR6JnUKn09/3a7I6QcVomKfkzvw3T1+wDt
pnjbL2fxcWcgRlVFD2jhjUk/Di+//BIft9YRUxhD/Nw5d3kSR9izNTMJnYQmHtyx
wX1K1QzlmigEEMfeyR+il7UE/7RIq5lDfb+naNdcsKWgDt1TSep2fTBodJju1sAp
HFOUHzkcECX/yggIYLLReYTjAcA6Ya8QXDIDj57Kxxb4zo92eRiBeKGnZagOvlJt
uFIRB8THhV2fNFcdXA8MRBEUGzJx5G8hIlQwYiVDzjnBljFhm15KOrOkQw7EQ9fL
rvPCwsQGwaAdnufpj0HdFgKhti/PKD9gXaanEeKdUGyVex95MSY4eNWuhz4Kn1d7
Mb5JYlPsxl7lmCZGDzVAznr4PtUvean/1x/Bd24ZhKfiRZ3HpS41UAU4XTFagprt
4DhwQ1S+JdB36AaTCcn6+LZbZz0GjPEbSO0sJMJcTZtUGvoW/nWw36OIsEAmVDJk
DK66jW620hFj2wcyGEkQSEPKplohTf1wjs8NZMhTD80scPynibSmHtKpZ/335IKB
EjdxXjzDSf4EiiArtSeg0T0c7G6miq1lA2ZKkb+h70cJpHBye44TVqnQC85DcqZw
7/E/kpmGPBHr4wZcHT23eepcALtUO34TbLuxJ0S4qr2cKvRJChqQ7Ou3vq+r+us0
md20+5aILEW1EfbTQjgMOMZz10kpajStFUs5/nSnVli/okZAl3l1NvnJWFME18pC
5efigX2M7/eQbDs93sDFc1S1kq8Ogx6h5/yUBFhDowCVTBn2L8MQeZAVUvEvt6cq
xy1fXTASPleTyw+dNnR//DF5iQRFtil3GgouEiRprGCppmooL5Xdh44pPz2suCGK
e5YHdrYQMkAf1P/SPRRVSfb4KGIr1NMfjAIOUrmdeiM5RKEv5EtAUJIiFxHRfSfH
ERn4s1C9OG+cHpvxY+PqoKsoX3hOx5hIk1YKayqhAoHxcYQiqWb6mpSrF6A8CukB
Oia8Inh+6j4TkjErMugI5HpwPLgnjEZE2JXGPM/3yOQNfDT4aRAgoY9z0YpHPRlc
wcVeQhGfX6gkVzHG3SSnD6qI4luexk/3mDuSJKXbvwvFrwFAM7VypWYRl6EbXDzu
htWLb6GUBOtLEGMKeE3xRRZHH+oyUxnZ6bIqvIWAlkBtkl1An+spGGkb1A5CLBDD
xSjTqeeDWzw8sPl7Sf96IdFqdFREDlU0LJZ5ra8GujSnoSN9LQfRNEeC/AQbWl3F
MF2Nsn5YIn3SojjXsy1sM5OXKgG0EYa3OJ27Zo7FoxCEAp14PF4wx+CqdTFglkQq
xBc12NBN9IrZxggHT6ytAmvg8BrSY9xtGqaKma/o9XcIPuPxbzCBYMRJTnh4vd0/
n4qto47+U7XLqIcxRnS4DLYRVXD47Ifs504P/wasWZ8MPkuVmCBfxucr8r+nE5W0
6RK4nntRw5QRVetHObA3jJ35Hyd4qgvT5odu/0HPU7Zvxvq2QP3DfnUlknWZYTiW
0wOroYMqQkwpGKtomzd0O2O1pToYXFtvvPKlj7gkUfiOnkXMDrYa/nTEYQoNI/L8
Uud9VBGc6wRN/PGwDOSaot4lU7xrLAq2n+3uoVQU04hlOGF4t+5QvSNURIbRZ9AL
eQliWxbtKywkcSEWMrbkTrC53ck1GZy7e7cAtcRhilGwQRGb1wI9hJaiNyS2fQyo
ODBJgJTGAso7/Gk0klPAngizEqQvB3WfSxD454hMup3kxVUHEKLeaWDvc07e3OEz
j7Pnx8ncVh45/1otkoFAdJgt0u9MXdglgHse79ziQS+qeZCvFlPHkf90htfaCGO/
OiutntG6RVmGgLPniFiNAMimdxs4PgXafw7Fjbfo5fEe9Lul7pWhcwaiWHuXFhgo
TOTVwN03S1Wl7x0/8CMEUasqX0QljeZcStqpA+VJAtGtGiGI3n9JBB+LF7inP/4Y
9CzsTiYoyp10K8Bk/YwzVa0sW6LqQI5l2JNWzeP5dSP3AQl/0yl9EmW76UaEA9Ev
/v8SCHuJjAzfWcTAKU3LSaPH78k0fZDkatl+zdjNxsYa8u4J545jhE7QUU1z93kX
3TBcWMfIaSX7FFLoLuaJu3sl5l2wxi4yYKdpNFE2w1b6mKbnSwZPW2U7eaPAhPF8
L6+CrDH4qP2RtuLd4ooyKTHP1CdkWLwamAWiR1QjAYI2SlR/u3VbvA7Mt87LHGYH
FtYHUZhfrDEe2B0VXZZdhEy0m39lV9O9JPLGHqPFiNQ0CTZIkQJJN0vKvj8jfXic
h8arbTrVYSgRJlahfEuQvQtUGgAap55nQ7QD/oeJmsq2/SKue+XW7ZpEeNhNsZaX
lrxqhpEboX9+/u8wMGlXb1aYo0LGbIYlR43vaX3D2B+JtUOtdATYifV4HlyTek41
JDtbZhP2ageTr0hUgX6v0OFIc2ZthHCSpHCrn7nL1PTWbvlhmjpIOV4nhpCt8oRv
YGt1BaXx+9+MRfDfxr2y8Jeo1Jab5kIhROVVK/lVneRuxi5Rf9nxuY7aQvv4n40R
8AuTiJTvew/8v1IuxiB6XTOF6oZerngF8NnWGJTnZE8UVgPOqPcIjzhSEQfsbhZX
se0D/8IFyF7Fqyzk9Nq4PbnkEF+EuEW4J8tQsHxTF/I7Elt+hR8Rost549ls8aTP
auT4lXfpfljWsdz51FQhQnWjxdxA/0urnkuJoPUCeXBJBLRwzQo8oQOQ48/C8fU3
4xNSJM07jA2+GtJzIeLgxSPfXmq0w0mojaKSrfx7dqQI8l6t6sNl+v6ZoYG4xqZ2
M1n9na8vI/OwiYr6uf5HCV0FPkfAMWGV+jXHM6muMvzID6n5zKFFFv00oGEpviGX
bue8QfkiZM/nxGREg8mk0jsyEHDVFsXn+LV7xvx/25k9oHey+O0C6T5I2sm7heTN
UZ3NXJi9uckfEgssOvAikjUTPk8k/9gwzzcpPKz6PU22RHArC/H6XONqX4WFVJd6
YclplI5wsbnticu1f2etPsTA2EZ7DO1TGkJuczrAnVf29tWtcDw006xIvII3clTN
nFqWjE0uNrVTsDy0PpZBmwCFn5OCyVcpTMHvASbXym8L6SIHEC7Bdkr00Ey2K7Xj
R6yLQT0jCt0NyJJZSyKkS306NBbffCiUB5pK9W1TdjZIVu32lHv5gzad67kJLjLC
h69KUuUPE7mHicBrLkaPh0+OYdJaQ8Ak5RWR0XNH+3UDklSrLjM3kSUHoMEwtE5y
aXN62Dy5rvHigNahCo5iV/TP2mi5+SqPqNPNnxLQ0qCPx6pt3ZFLRqwqgOeOcAqH
u9ck+h0bNcpUegUrb4aj7jH4xQ/zku2HS2jaYfb03O0fUsUL47M9Q9aCpVCJ/4g5
WDeCrU1/mrhJH1XGtlzEnOTbd8TOzSc19tC0R2kZxOFefhntDF6OoYlQ2SpxJoMR
oZDy77+g5WNTOpYlpBX1vaM0YZTEAiM/EsFtHM6GvhTz9hnevLzGhbG4f/JDN188
I4v3rs3EvH9y8q5dJytxkYS5Z3B3ssUooBauX15BZqoRu2tqcwhLFo4rOckCJtI5
G4ZaBPw6pLxENvBf4Y5zhpNb9cXghbaDDRG8LpL9ELyQL6MoK/lBD6V00lDIEjCW
vzivJkX+MhVDi/ycwllW3mMVf8h+Lc7ri43mhh3xMWktS+aL0x1gOlA/7jZenBsR
fxpDAQ2RDi4I/y0amK1sVG1HsIJl7/QVanFII+X+Z2OGYf4FeKdHRJZu9FRTbWDx
yTIaVpwIV7/JmFftQT4+QqpLq0a1qfGJR8DcvzLMRWeh+0sOuGuRcA34JRIAEshb
y72nKLegnm6rp8F7nB8hskdOiG7TNH8JrtECL4UeGm9OoMXoeKPF+7k6TUz9GeDf
M/FOzei6d5T/ehspzRt2eJOCCPJ3DUfUw+UJDNIhNCywBE1HA6kpqsoAMo9SzpqC
2/xOtWm8nRFlsLQi77gnQdJNQEoEsVAg69G+cqBMjQXIai0xbIWpXluRCjNLDYND
0vMJ/6iCSBbHShRnz3MezDhJarkkKGfsoImjxDqKWKCw7OwRkdBScOXU5bne7HkP
G0sBAKjG5FEkS/btATvepwyi9gDXtCnP9cCMontvNaZs/hNwMPt4uvntJW/jekI/
zxwlRM1sH9P/XLMPJGDxBMi0xqE7NqxSl8JyZ0UM3pV1fss+acWZ+VqoytLcoomZ
CR6AEYFrTdjVo5NaGE12+ojgWCziis/zcgklcUfzvFrWX+2zks2GPNT9cw/n6uGa
JQvP/SjI4ujSM1PAB0tXDZ796VVpepGJuoEFl1P4ISOyPzM//qAWWfWnZUvw+91+
PbrrqAiYXCjDnKglzOISwrkYO6cPcOrKaBwksSFkLEYftdNmaBJXshfMpNe6zNFZ
NNaXBnvntBO9KuttR5B9EtL+2KP7mDSr1jVEM/YbAWpbbGQZe8lH0HTsfBRaBft3
/Hft+aT+HbZ96Jn3NCkYC5k9ciECXTmIM7eH7P/IzmAMreIfdiiKJpba/Qa208AK
+q1eqZVUnBDTig+a6XpxZl7tvvpSWx7dC5TDNObEdw1n4TelMUQyWITsaScObbrf
t0ghPbZ3nmvKNIEguOm+Cc3jeBEMzw7jQyBZFdFUEtAkeYBhXTaP0yXVWE/4VThX
pSu4Islbddp/p9pxQP/NxeMkr8CO1h5PEoGm9hC8xcseC2onvjQyOiLk1k/k7Rzb
od9F4ZEnY4oRVUeS1NmogQ1vwGGeulO2YpcwsvXA8e07oommO/d1fEJ6JQXMfMSK
Y7bJviSug2VMfN1e7nxXBJbGgqgCZZiuVGGQq0QqHlFb/7ozgwDfrc+9LKgKexuW
U4SiaazcJhnYaENO1QHLc9aunSkwbSyUDeErFZdjmPJIwQT3uinQd7vOig6TGUbM
d3mq5vhn2qIXHzsf9M/VUurELLktve4dC26X0Vjy4RGDF6V4ANpxt+zSYIVc5gHk
I7WGHO6vISSgBudy8Styl18qSWukbrDl/yueoI9IHZfYkugnZlEKoe63KMKMtQ0g
PdXmj6csJDb48Dm1bFdOO8XOBG3EvWcm4i6OxBZQtfB/21uZQUAn4GHvaQMWABas
dSki9chbSLWUJZZNM8MQxGEfnwna/hmtzNw4RiBD+Hwtp5+LpkM8Nzd5sutKBDXR
TC4aECy5cDn/H+WXOv98+vZG4jQunJYF3fWilLD5QUEoyDr+WcqKCN4yf3AyTLrK
U690pBaxHQcv+S14FbJqhxtewrH4vCvLNUinFS2s0C/h0FMQBC8ZJynEV/zATb/E
VzGjEa1aXd46Eh+LwyeUhTD4+ZTytk7nkVHZ6Ndv07eQxpzkVqYtt/8UePms3Aah
U90RP/9rPYWhIW6sYl0nBNBnZp4VmR79Yqhe0Pkv2wfSPim9q0lblWvZP+RhYJbZ
NEDSkU/Wj49GFldN3UmltmhKqwKp0QMHUvi81f/tTxKDFAnBGz2yj3daDtGtI5zd
K1TS782rog3FPA+0XsmrZee2GmMlob8i5HWS4tGfYJx5rFYQXHzVraROlWeK0l3i
V/HfNocHn+ZF46ClNk4msg3jbEsjbt/Y2SsEAn+MFws49KKleZr5OGejGa7XohFU
nhS9x/NfW6Y/3z8Ax8C/9ZF041S/H8ngdfEfMjZPStzxwHpTMOljpZh7Ekmg4g8x
AD13aEmxS1OlGxwO2iCize8EGB+y0g8IvQk3Z6zyYP1WPwgtR5CJXBNRP57W+eGr
wDyQfQQQvTv/MTfxBniYOQJv+dLj956xfq1eNxmn71Gl/eRuJCLspU3PfBPTVH3X
vLbYsG7RQAF4Wgoq20HYzh1qcM0JaZ07zDoCghQT7p08+FvaJZE57477iVXTEyB9
9ZUyGlrdjGJKWw9MGx9w/87gDVW2YKCi5Eu0/Fxv7d90qiGqrN4Qgk7F5oW5Hwfu
diY9kjY7yGOFWPICniqtY1SkqrZrOiGPVJgWSku+OkZDX98K1URo2Clqp0updNs3
BdhXkUEzu+Audk70heodrojj85TJUS31Z/Ev3VfcQ2vG4r4rkbbzdFlPBWEMhtI0
AtaPbGFkj+x+MFV6tKC23xSpoOXbWDeTuAxouNKKHlhFC6TmLcBmFmujwHlYl0ll
wMhSBcapY6wmvldS6Mt0EAkj78QqPei8Ttyk4kBfnR+cQr8gwDPxIhcN8+/3syzk
fSWdhURxtQE36+mipKWlIGy29SW27znkziajqp3G1bvZwYV4ZZwD2bcFecy55wLE
6qkWOTCY4CkFW/M9U6bxk2ojjGtTrNz7M7GwPeubvirgWDadDqel1ha+8y/kXdRj
F2QlVasRIkLHKoEiJkQXE6nGW1VGDXKfgg3PXRX9RuFXsVv+YkwCnxrfinspwG4Z
qmqT+P6dDbvlJRiwRTtzRsSGqVhJMkT8itH0XEuMpjad5L7KRLVa8cww2rgrLG3g
Ssd9BopzfJ97arcoPhOCqHp9I6mP0WdX8b4wXQnEanhcOb4opH7sAA5v8e2aR98E
iUTZaI9RnGOUd2AUMZvC37lw4seI3QwlPj79ZHcteM1R3RrFbAzsRl3ZhB0YTsjT
XG8BB1Ui9w8o+dQXEsiPfAg89GsaEVKezpdiYi5FK3cjEIu/RY4cEHiD+Y1Shg5f
8X2GHkTl65ZxkAPyPstPC04ZwV+mbTEqJaqA0pHd1WITWdQZ7IPSPvonFhb4UJpt
urXLo6TcGGYE86oh8OLabMvsiV/9fMlbldKbpVN5ppDqEdloz+6NkJSN7BOaI+xT
a9al4yfzuNzS4MHJDUgPND1VQegewfshPO8WTBwatb/XGKO+QvmJJ/RXVnfCOul9
FjCVqaHounqbF+b6zymwzzvJsAvizRwyIa2CKVI5vQGsdnMh6F48Ti4zemAWiE5f
Rh7sbFjBX8eWXUX8PvocJid7M2IJuq1tAhyIRFx1V01lOjUGdY6fp9kZys1irAvM
nEjyYs8CW6TpCyEOQrd9a0uCzunrVFIY1HD11cCanYa+iLE7s7zInjATDT4EvUjl
gj74MIaHuF5B51oAIWGJS8sovcu+bjTvyScIWO6CfMq/kIUQsW7E5bYvrnxzEncs
hCKcAdeUmNkNNUKzMrhi9hBYWGXXiE5vmjLZx5U78GTfxSH6xk8Ed769fGdtyqNA
i7ilCcSt8lKDtqtYgSUZiYBiuWJ84UjTbxmQ1odLjU8ud7Rguac+CRGGgySlNLOj
NY5D8GYew6UX0+R5aw8c/EWcJfckn9Bbndre6iqFyQTscK7AlSCvvdoP1aaLnd4g
pQAsZLvXP6oQl8PLIwfoPy1ok+p77ifcpDL4darC4u+43cKSZKLgpX6UO1Epjk3+
siksqf3/PFnW0ZFGvH8s0+03kexZyK3S9QGVAVnQzdU4aNR9A8zkDutrhtItD0yc
YrGLfNIHAtrjlu6vCQPbPWDYp6HWbdQQs98aRE7hSI8TdBRhynhs0jQq2STs2roU
LyC6ajf1NpDgXKt/5boU2CvMipvVNkaFq/Gzg/sCG29gQTCWc5iOXCxBE1FaCA39
x5ftqXh8hX/YkF/Z7p9gdz5SL4i5jxY3YbbBAw6TOIjzsylv4IWR2LPhqZQqSAW8
tstJrCtzg39unGGWL9We+IE2tIuoAfP5083+cK+dXfwFZ1z6s/3A6iFI/qW783Kv
RkQXyOjmqkHXN4MgYhT45LID8IXADChkNVkain7AV8U3yVWSbFcOq27WoEG5RXgM
IEXrooBLoTgBiu2n70rWLY5+RFMdqgIRxgqAih7kLPMg3J9zO4T55KmT+SP9X9Pg
L8ERHOSImAbuH/3DTyQHUDwOyEDA1Uk298fWIxTOc3d0pQovt7Z1mi85K443oW5U
8D3Ly25OhKEWGlhoKaR6Rin0Nj3Fzsbw7p+5owaAThHQUbuuoUUbWUY9uYt9dG1z
b78sK6O2OcUYAIFM7hvyRYMHZM4B0NT/854iqe2H0sYBaJBDjUj83E8gja1XHp2o
lWrzQqwh1XUkTWWlyeTZ9YO8Xqx0sFF/z3VL4SAocG/9FF4FZ/bwAmAJrXwLOJD6
//Ph0l64aODhhzcIykJqODaYDtQ9mNVj1gbC8rGFmKpxaQT0KR/4ZlNaj1o+15F+
+UhUC47Io3IUOaD5JcUyX2ef+jm8MdeBRteI/ZAdF6yo2ktOCFqa+XTxtj8FDLdC
tA0o45AvIc40iUMQPKBSAdfc8876K/r6eIQonqLVOo2OvZzJFvqb0IOdoBSZ2MFZ
WR1pEJVsA2SCeaKLa3WEz8o5hq0gLQaF9xp1FICJWJEAUIEsjegHogNlRUUoELG6
kbGW+Tfmj50felHiayl1VyYDpHqHL2J8JTJL0m0xFnaasHCPjW86vf/2M8+mdkZw
pF61jFu32srl2AJZaBal4aH6TYxTev692kMckmNHGX7x56T1x6+lRVvudUHBiega
GGCQo2AU32vgzL3Yg8HhW+j24Uv5XMgaiMrxXjKVUIljGTR7YXrRF9rEgPL/xycF
th987w9vsFVk2E/26rLnwvFpOELBsY2/X8BZlCwmsYx319aLhKPV8kXzMUKV/u/m
D5rAQe0hRZnCI4zY74Yq8V75U/kYrBunlyzc6b8UqmYeORtqJRmVb+Kkbr1r0RiK
SPTVvu7oX+ZAGby+QUDzkYNf1MhnWkzCcY7Q0z3wOGXN/4GaUIxXOaa7EQgB17yd
iHRQz/KjOaM0Awx3dRhc1XQF/LPP3BjaPh4uR7sNCC4h/c04rC5LlJdTqKAc/G0G
ba9YRvVuVB88kQIf5I/98Q98VfQ+KYAJYM8GVfSDFc9+6E9z9CL/uZDlJjmUrmO0
q8l2FklgY0VNYeaZAONcZnUrmjm+1rnH5mYJOpdS+KlV36wNlWykOy6s62YVzvqP
XkSDJW2AEiupS835HUAktXapshPoQKr6wSUomUGWQBNlM1bkNjIoO2MzaPSixSrc
r0HCd8IhikF9K80jbmmr340i+frVWaT5Vz3Wb8vVdLdQq1oVuUqpo+KcuxUzJnFq
/DUUoUdWkDObRKej7vhlFo4nViVZfJpitfLvgiqwYZL5x16eoSTdHZ2bDM39OXKf
W13XZ9jjiyEPpsYVdoxpmG/pQWs46PbOgwEU30AO3253xl4shPoGbRWUhexUX2aq
fchWYiWxh2df3ax8iorrZoaQHjul6WxlmXEp4syLAywZto8YnvusW2RaVJacqBH5
k1HfpGi+1MjqNjBeJXIU78LPQQI4gy0lDTUpQJtdT3oBQhUA1VTXbvYHxMzC2xdN
mo01xOfX9hmNn73fzV9GfVvLRwxfas/z0h+go1CIwQss76LlOS6Wxby3dkty6kBj
OMVy1lHKxr3wjbpyZqo4fNiAGQ+8xLdBZg1O4wE9+unwObMsI7RsOLVxYGbj2Lxn
Xq4mxpm2+BHQejk3/I81l9shT+Ro59vftO/Gcc5/subCtXZvudVIbh6MF5o+4UKf
nCtB60CfY19C8RbQGiG5V+6fmemmvJmkVY7shjC1TTn2V3BBYqoad2zOW95lmFJy
tKEvzdFkgjVGf5+S1IFepJf8UZzHIstXMqmZ20ZDeHhm6hl631LktPq2liO9snGK
Wr+GMGfl0nL6ZmH4Wj3E4gAipME5KUpiaSkOtvmL6YJZcO5n6Q+aEshZ1ici0/T5
O6SVBAnY1e6eV3aZ+/kpxJBHsKMxK1w1GrYVoqkY19ahr7AY+4Omp0seZFGha7UW
6k7iXx3X16bC+zSkC7ynKQOifbMy7+f2Dwmk1Q7J72ACAhIFmdDRsfsP4hDvUQGg
HqvoOxu37TRUidiKhPLvaY5IdBB6JjXJu75r8ZKGMAti3VHjYz+tW//GddcUMwMR
EQAMh0GECCNlt7KkvNABxbz8hmmsNIRehgLwbPR31JOAAqJfcSPW9PxmQoLhyu9a
6D5OuCmSkgx6nTLtDgDhzTWUrlAm91LvVHGOOKsUobwviRrU5dR6REwCTTF8K+E4
lLPjEjoYC/3QuQKNzKE/mRvrVOtkedY0OeRWHfJqgYrMF9MC5TLHpTzyBqV9l//g
rsHaisbpfbdUK/el5v+X2JxGNroC3NhODWRISNPYJ1qO8JNrukuqwg0z4vuwxaPP
wfLFvyRhbk1jM3BkPM6GLCi2wqlFTTkGZ3oeYJe8PoUC2c3u5PClHxr5IxZAa2gY
JM3VB9pRCheWbARR7X5qcFU0GJPXlfPmuHvoDBE50f76mKdVxzQCOjbws4jpL1+2
ywjDLdSVCmmurKRYTMhsQNNm6ej2vY/pap8wrLqN0N0R0Zr/ET00VSrD5Rbnb3Zm
VpO9T42Ymz3TUbgQFk6ndyA6hh1SSmCsF03urp8WM/FA7cb+I4tq1cKgt3G6c2Z8
/K9M+nJFbzvcHpqvnf5QheWDKe55XrVFJ252AmlBvcQsFSuDXI/6UxvP4HJPYpIV
ZaWD5jDwu32XiSgYA8jV1Z+plOwVZCbRG1eCJ+r6r8gCcXz8nk5gNEuj1dQLB1V/
SG+yvnjnFDCAOq9BFH1nVWw/z7Lu8MeQWgWO0MkSHRQfAJ9baVrLDY4EYffoKo33
NhNh01m9+oPVVQcRiJGnGWiryYhC1KXV0L83+L52a4d5k+4Iy9kuNDdVd6hTLu/I
c51j2+wlvwf6e4QscrWXicJsuYqtOKw5D0dGBsLGaT48+PrY249Tn0KgGzILdOjK
syy56BIAB6wzHLSiJgGyaHk8aGeBrQHu9iao2qnH3hPqSWMQ4FW3cIevhbcW1mXg
YXKZhJiu8YMunMq7Q3JYMQZFjsiDR7i4Vug7Pz2dahHE/6DDLSMnIzDxtFrgdrk4
6xHUWEztJwHjmQeMSkBczh/iobgIZvBkfJH6ua+vSxi8sgCPE+rJB8NazY9EpRbK
tXDGpgkxQb00DB8GtuGLf1iGNZj0wiMAvLQuSFRMWjp8ETuF77TxUvqk9RiEod4r
jLP0ElY+5s2K36lZgnFA+48H00pWXHjXR3XSvGr33QH5I+dnr/GIK2BkBVy8z6nv
RQ+wpC8UPXOIOgC8bwWOA9dl1zRIY9Mh19H8fPUDQkig3QfLZIkef/cIqLomWA9Q
GpxQJmUT2QaJNWyfSNQkzOVk4BES57ENzWdrw3kOsIcMyC5aTkZgsAody9LPF6R4
HugWzHrzFCEidoBey4/S+xLHLPzRq7gjbiYpReyL4h5At2uTkUPMBb2kRFeNL+v8
gywwauUbwKmMtWPykAVE7NJdQ9hiGLoelRrU8YSDcMB3onK27hm234f7H8NGAqHw
7IhXrNERp4JpIDzC5V89ZGtEkTQsEvZiyl/8+Xnc84j1F3H6HIHKett4AbIbN3Hp
KiN1c6AJg2A0oHeeLl92omN/n09iQrHe90rB+VQhOTjgY1gvtOcBIS9ZU5nPiEce
Pr44DXXTYbMAS9Y/RFC7TUqRmYzBC/MkGAqS8ihP6zHEWNCojMSLDDJ7C/bqdedG
oBN5zv9JJYGXaFCcgj5nYAK3Ox1lzA1G0QyUWepq3jOF9UBy4/s9ZVhteEgldAvB
gCmh3DfJd/p9Xi3UIbSr2wP+8zTl+NEgY5xl3ZPtQ2LIZFT8mW7mDI/RWV8LGf1k
OK+kzXB8R84o+LB9rK56WDVGKg7yY81VjpfBLwgRHMbTvtLsHEMiCpc/Q8cMCuai
Ay0YzdQa2ZpbwczOQCE6hnlb6ni3/hF7KT1fNzHHcAKZ9O2M8NJQpr2ZB9ajH/hp
m8TTjxwtBxqW3SyXuOQKnoCa7AO64SJ1lATHVLDDKsFFo2P4Ki0V57pjjesCFehi
P7ae4dGkzVCOrWl2N4rsBy0sn/40yrCt/e6kNbXJbQGMC7aEM3SjFiCEu4HkHG//
Jla+8o9e+yEf133llPU1R8GcanW7FpNqW2f/2XXQZH7f5kh5ynfpKRXcPk59f+fp
/MbyncUNLHVBTRf7+pZ5cljbw6BznYi6LXPwZpUYgYqcEz3DUSME+F/LVPqKXtFP
f7u544WjJbn9+ieKAxMMx5hUDIt8MK/qaBTf46kLoskITjwvVYdL7yNn9HhNWOPv
V8Q8O7k80dwx5yZpmk7XD+i2l+s49eZ5+RSTSfbeBkdj4xR5DOmto8unF/PQiNhU
7giKlfgA46BoZ4D5YWCEkyZosgtpNtIxcrxoOEjgExrYXrvnlGcnxRGY+3PTS9F8
q1WrK26/A+fLKgI34x4p938icbpn5CxsNCix5J7O6hZjlAPo6IiegVJjKy0xQSPX
leurdCLqkw3H5N0dzSXbgh73WabDIjthuPVHE3zai4tpP7QmKylhj1LYagkqKYEr
V42EA6ijh0eku9RMf3O3CvZT4m6XGusVH1wiDfz5VOk5v/jcfBeQl8zif31HOHs+
ey11992wx0rG8YghAfFsbQb2xYMhxvkc3UQH99mg9IR65ODUPMW0yQMpvXmP/CRr
cOwf19uJN4A0fYV6c6Hp99TcaMAKXIJZ0t+GpxgFvhWP+CSprxvENcBXgVuw6xi+
e2rsLyDmuEY9YFn+sVTGUxZhoFn5qmNBRyrk213O25yGX33dsbomuI3LULeH2OTB
Td28cGpvTlXR0UlqGgbenXbovTUi6Y9BISmJ7Pqqe2BaFrxz6smvw+epIc7G8mA9
Mo1hHnvVfq3jO2kBpp6L4fRD3FtOktUtqGdqhoMjiMWFjYryP5dKLOt9sDCgMGqE
XJ6R1VeO329xcFm/R/JkQBMPPVwOcaD2s1WfK7kH4LdX3lm0A0d/cK096G0c1nnM
GExDxx1vcjLm9s47c9kKXEQKma7IZD8pyvxn4AkW0nS+qat6yf+cTem2DyJP753v
mVlTaqTXgNIPxN47WImtjvpiCgEhCpo1RpHYTMJCBIUAeiTqlrQrAVZ6CV4aKK0Q
AaKPvStAg8Crf2V20BpH3IxroxmAl5FfF0BYj457RJjSNbeaFeDzssz3RCyf2OBk
N1TexeISQrnVzec+YszFhkzYv5fb3YACxkhKgSs8nhHSUdKLLmZ7vdvYaFwaky00
FXrblUIEgwll1Bui22BAL/naK++md/sgV57muG13qo40ejD1PHeZjXgTK6Q0GgTG
EOLStq31wSrUqdUzxESGsejXzeEvP9TintnWYBETMa8nSlfkXCsZ/gAPB+aX7Pxu
FuPw5PVFf4qcV1gK53yBlwF1CsNkfrINPHbsMkd0nwOnztTBiyq8/PWkhmwDCpIO
GWThlOVUdkn8iL4f1XoLIjtSTjFOAs0l0a/39fEOuEDltgGsBVydQazTtLr1vHCv
aF4amwkbKHOSwlBiVOhvuRtYg7tPqGLQ6O0vdt68mvIfqRw1z4yR1A1WlSM7788H
9PtR2wWNvvrk1gEgAT3FqOgnU6JT4DuSuGVM49JUYAktldZyiNsxV73jOWUtvOeu
RkasZs7MbQHXIcQ9cDL9iePO2v5N0bexsxbu0R0cmOH7jeNBCeI6qa9OWumE23uH
mFnrpRIbZs5JgGssEVqaUT2Suh8BhBGo95JSi+DtxqAN4914DcgJBW1nThGb3e8V
O++ymfBVmjq+EQK6AmrGEEC++yCTXrGXKj6zulm3oow9vhIH9kQ0PPpeJ0uK3bNb
TmNyTCR9liqm1O9mmbAlrK6P52PPrLnWP4g5i+Y7tlm7VJssePLX5SWqI8UbH/4S
RZ4twzCr60cnb5vIoFvlTMDjmAiZ/CgQfKxyybKxmZWARiOPeH9MJx+JWRCGewwH
S0P12XU5td0rkV7gAltJ2dBTv5V+uflimRWP9yYqZUEqMPi3W0VSHauq9qHrBGl1
AqWuPgLOkqcvb9NyfEY+gG8aPDH+IluWLhtempL1S9MLlOs68Povrp8adPU6CadM
CPRbCzNfiYqX3Y7u6jQTRc3tJV+xTH8mkusyPQeEyaZ53l62exdqNz8LN/0E5XtP
5Bq3swqhrdc3LwtQ39rS3oPGHMhDFH75ls8/csEwjib2iuN9PGAecQTv65TOFEAk
4RIRpPy4xQDitilyAFLaRka/S7CpGzh8k3KQShv3YXCtDQCxRKw1Cfc2ZbJFZqNE
OL3MqtGjelqovWIHjdTk6tmOgvhuj0P7Pax1NYupX/geoCu8tnLsTUa/tJDSVfl5
EQ5FL8VIZR5lPsH/RXmGyvNEdPw+WUb5F3blg8ipxg42X+OIXOqnxpbttIVSs2ET
subSFtO0wPR+D2Ppf0GFmCk27IYrb1J02xEfXr8W1a6M+GYywfv8pYbBGIYsYhEH
QoDNu9Zh2PU+cdYOP7Shh9jyiCGTUhyAo3kiRzr+B3VysZsklvta98l2+6oGVZlL
U8uus9hXJ5TPyrm67/K8LOaULBoPFREKLXe+i+tm7gzG1yRe+Qv9CXk4aRulFFP9
P4RZZ/mUVOcDUVNBYYo8s3vNdDeVrgVDFu0TJP/ppq9uJ413IE9lhxVMUC9m/sV8
7xu9czTPD4ZLsh5JQR6vaj3s/KEGhwvHeH9wG7Y+V7dBZPUuseJ24DzLbISHc79l
DIwggR9E/zuuPRdL4KL5POEHOqCY2q+2bdsAOrvXFBN/AL6Jx/gwG8HFc61ttyxq
UpKlKJNFhyqzNmuq2xOdONJyGJL+X79Eku1PT/LjHhunVwGkvFBuj/27WUh4vTT9
ZiaPW+087JdxPPXE+GR5g9fhreZ8SnZ7nKocZMuD5apsxvs8UPwZ7o2Q1EtrWXKh
XEm0hMDdpqTkKxhlkf61EFnJbr5cECT3kdymqv4CIaWR5sCbpp5ubiRhXUzJ1pSW
MVXVwpInSBoxlYOXQNFgYs+5K6oVwklvAvS2EVj36Z6ewGM5MKDwMLeS4m2IEoGR
ICbUWvgALtWDzrknkDxciNgY0IV+yUDwztWF9bEYNKzSKkHjzKkHGKOx4kwZOsTY
OctmHG6f8LsFmKouCJblE9+DEbR9Yo3BE+G3t5Egk40KGLAW28QfBsJcSmiDs8Gn
mRc31QPdKwQdmL5TbHC8yfkVKCmpzRyE2I5+U20cn4cSxhU+6iy6aFgqvRifD+SX
YVIVqXfhvpOFNpiKnnny6/SHNMmxjelCDe9R1vPk3Sl7gxnrCDoaV6CqNzFhUVEu
mR3yx0xW/42PIZnJw5aepJkSo/FuxbqZ2ZCluW8W/tt6jNBG0gmb7zM1zL0r4izP
JGrQiG05jEqkjhuQ01y1XxGlBlb+NpV7p0bbHklwjw/tNa+trV8MJQmaf8ullyIZ
1/+NURPXpBvG4RBJHbLzAWF30gINhEFnceL1hA5xrGaqCi4MecZCxR2N1+YMwzUf
Rn3+ZvSwmhiHPwI/lmisOhTkCZx/QR6YZpXld/w741V7tTnGq5+0SxvQXzqqbQXB
APe2ZLxKQ2aVy9CMK7WQhonUvMMAU2Xi22ALehdTibE3FolrkBfsNsPMC/AY26q8
Rt1yWCDxgsuA2NP1th0Yavq7njTWwzQgWPaK4OLgq9nxnqSdBSgS7F1ijIPEqJbR
L+TB40nEZs3NoQHd8D4zTJImm3jp5YrguNRHDlvWaOXvtyBclgB4PhqmHm9+HvDx
OUl8EhNHOmKnjHCZQztb2DXwxQMBYUQ2oldklOjsg8OMBsmUuo1CZ37/M4dqWUQM
4HPemR7wiB/8PsOjUBd3/n2VtQMNSWLHakJ23u1P6R7z5pKZzXkh58mKuoAwmu1S
zPT/ussazBksevFfGMsLEp/DpVfi54emFPwJYlNVTEN3Zq1iz2kCWdhcS6hX/5GT
xjSN1yNMQ2LGX858fizjMyfdMR6log7+VS8f+/tfDmA+QKy8PYjLMKKalR3GAZ4/
Xpt5eeGfE2Fvk5zje0OMiHw4inW+B1ZV6UYP4jGxiiVnOiA2TGGD6AO7andaf5zS
U/2RwpoqRyW8VhVDhq13TOy8FWz7G4lV+kupYIoKRv/89wS/FecyhY8JGAuKyPTr
QuJpeP32yNi6cbGBDV8jT9wz6DNywUjKlniiZnRCGEckluuS+jbfDDyHB9R/l2fc
HK7eN7SdOiWtAE87Qo83G/JELZFQRg064y/PKimHNcLSFGpLLw3Z2SB2AiV7Le8Y
itlBqAYDyzeeye0qrENBSEX+loiUH2MeJsbh9hIxO+270Cx+0wZEpIhYh2zTPbi0
xqbyQlk1bywJaqroPEEYXWvGJDmMJHdvvOSpFZgct8WcTsEdoPhC+pjtUcIljrOY
opPKVGRXJtvE0bWEF9h/dRvUh/l/4y4//zbZDCZNfgGFrvN/EoEWbvlMlwzj9+T0
yhTBFat5krWEEd21yAGT8fd59hWwbBFH7Yr0Sd4uCQQuT6SiKDc47xHLnObgWjJ0
Jtrv5uGnaqLqyiei4YYUmHuM9tkJwtzWJtVLrQet7K+ZhCfEiaMc1t2i+hU6oXZT
8CBEwsRaQMrMDGXGf71aHhOlnHp1sFT20n0v4D0DJkUAPBtWvREmLZezZYvxuMDn
hY60dpLiwtd478VQ1yEEPzQLKqOmCofdLBr+DGr0qczxceW2Mt0M4flSagriwkpU
60xAkxjqnwrU5UuCednSHawtXB0bBqeEl2DOkW4iPEb6NzEOutsvyWKE52+J+eDc
kgmuqXOvzdzbl9EOOBwWku/OyLgHc/IeJcj5yL0HZm8XDFVPXs1rFmGMOAFhE4Yg
c6PK5YPAaLCUFQBtltnhaAAA5r4kgi00kyJOpeJvM4O6g39VErogjwr1Qm2awe9H
/c06S8TEeZ0oTqt5c7rmj++25XIGlonfb0bE9b/J6ivmssPdJWkran0fyX/4FvWL
+uHXfTrel1zfmmQpFZz0fEb3mZehVbPYrSd506YZAlojvwbSdOa0KwY2OekEP4th
09ZbeKfD8ukmaQNcoSLurayLql0SzjQNALS0A4KtuEZm51fdwax2c6ZNls2Hb9TA
p+V7oVPB+zoJbM1pYp0DFJiyLC1Ep6GwqFqRm423vg3c6FAksHBIYIfKFLGoKext
d8XxHf3rLyANeu45N8QsA/xfWq/PUq0nzgfRa+3qO29PRHa1wlCQ9Y64xH+pP5iN
LKZdiWqJ28q/k+dR93/xmY6+TO5JByLWH5wUw7ndubTIMfj4RNxpC+CJmjJhZjiE
0wL4DS4Y4Gll1PrDLeVGodmevUdFltDDtGYx7JrKOCd0cRYOKKjQ1+cC4WfVmMFL
ugG2ZWcU5Cmnmz/8EOXolgkZ6/Ovv/oF7Z+ZIdMKV7/8ipB2srpAq96akRtus2Rj
z60VPi7MhhVFj0SS2fOtFPxg8BqeT8HIsowKcd0fpCl8XVPwOXKa6871YSiSuL+S
TSxIVKdsqaQplj3WaapTyeCrWX/dOjY4CD7Z8xs5zSfwiNw0kK9LvKvCv2O3WX53
CN2eluiw5fT5rAnCZ+62ZQPGaqpqUejLc+wOjViGrr9c/RrUBMiWUNZtCpTl2kt8
uoxzj89uIHg4vZqOOHSujDz0mjvJgwCaYaSPuYWk2PO/nu9e37wYfOkVuHccPTp8
fURLrRh4LytReOqy4KMGNbO/11CZglOXDEX1oLyqCdUxVk6n/EEaK5TFi8BlJIc0
EvO1vTJA8NlMnWZBhpfJwSdxlDrCJq2T7DNM581vO5sHCzTYwljK9WktVPWbdv2q
7ys3ktDRR1nPhz38K6ynlOAIMW7gY8xXMu0h0BVvGA8jW4OWzWMaGAxa7Bijj6rV
J1V5PvD/BBNSidfgFJm1F/Fxt9JsFf9uIOynDyqtNsqmMnFW2bNFPWqaeJtiZjbN
rc1u9j8va67eMxJj5FZ7m99aPeig52oakZ2Po4T8DCb8B2LQ2zArg+tUva0LPW6S
WfYKF4HNeYuntVwSgzsIlZ9L+jlseMC3ruv6f+JM2/OVZYaBAe4PGPCfOnX+K+Gi
ZbTbtfJCptYrJ/hAZudNaUy5X9I+2bcY0x+pk60jTcSxaXPcLyfgqTFPOACqI4a3
L496MFB7h3cRlGIg3ne/92LumJgOVYREfz5Y66EX+fPCM8Dm64UfFKsZHVV23mFo
OGT9cOrSWolqZRRV6I+g2TJwmbpiCICft4tBaSzwOvHb1q+yc1tLKK6nBDebYN+k
EgAfGhCmZOozGbMhMA32vJfu6a4msnfZukucUWEjiuiTAjyygFb2Am6XQ+x8b8Ll
04sRYN4B4yCioyKNEiuq8Omn6lZwA6a3GytZWCoUiP8BQ3/ymwOJaCJC8wmrcSnO
k4qIca6uyjjV9eHbAITCpkyHiWCh+N4JZJHbBPmBvuiA5l34v0vbp1e5Gy9sFvml
7FWzsuigP7Ipow175jLZyXlpuFFcX1kT/StbZVT2STSR2nXWEFDmVRTcceIw3DDq
nknC28GnWYkqdnZsiM1QHjYFS9htsh+d4ts1Px4naBtjFiOXvnt9MuEC5zadcsON
+ksCuxZYzFsyquLOETEtD1yZOrG6FebHZhO8pfmtvxiVJmPidyghXH2amMLSGciC
u3L4BED+BrRepXfiK4YbVZElrfpVqiEuJYbZ6Ly8zprLkFAGKByMDKB9WmIIH5eB
X3jTHGAoiJNGyPwJblgmIxSjv89vX3YzpJHf3ohq+zWETHcJeETdhqYXc6dkiW7V
VstjJZRVrUcM9Y3szxWVQbm8DkMtCRMJr6Pew44w8ZvJgZZzfsKC290aA7mmbGAd
ie3V/jB58adD2VBf8+P8o+HL8rxqZ4cX5iZFAiEyHKP2oST0RTs55P5IqD5IKmtK
+dOn46O9gXdkiWsa7eEJHoTc5kfhz4wF9+bvAxbqhbhqwsUzKVPaitAp2bGYuwuR
wggQzi5S6C/Q0YIwERAgOAB3rWYFSwsudzkYQc91Ct2IiLkw0eLD4wn3sSaz93HN
95CbnJmJbFCVPrIBUuJzvff3izHmroQVAzXiPkXy4rpUBDZTZ91yUEyq8nom+KfZ
fkWyocinrrLspwN4o+ExHaWlIuz2DJPffotiN+r5a32tdiHsLgcro7Gxj23bZrD3
4h4wNBHbeo1U1EiLRl3VaxnYpJZIW0FEi3H0YXZYsNtSvzUFxL6PMKe+u722Vadg
KHFJLtUJFR2++C2oXBxZRlXBeJPmLT3DbLtW7bsEtLDRd5rOZgfz7oDjCcHiB2LO
qJ5DQJZwDD43706KmxpuU+HjeI+kuycPfbJBqdZesJdV9ULohqxu/kNKfIeqQIC/
yvF6DXkDQyk3BWkdsDgY5+0J0WGhSw8UlKwoaZRsxAPTgM0Ag6fJHEZ+UFxGwMV4
5k4HhcQcOyQ7LC45jqU30ITtoT+IHQOM0tVxZrg++5aBHsD/iajkYy9Eetew+TN4
bFpf/67f1ssGUMIs8PGvVe+8qcXMZMR5mMdnQvjit0lR4dWf0mHaDYqoqSI0xN9l
c0PIcAcou8m0YrE8qVYx62Se6G5IocFAQ0lsIsBbA4TXiQWe21vpYWpQpgtboX1M
PFJqqu5blAWsu2WSTiSZFonI8ghu0ZwPqgEIhf3KEev7ARERDZr7SldTlQvs1NUI
IrdPV3jiAoZEuxMavhp1qJ9NIeaQu/MUpKbBp19K7D0Vp7PsA9zez3vogshUQG6J
/FXyoJvibekEHqUxp2mdZaEHGjMwhgh2mBRf1GlYWqC1CahF5cT0vIkrKHIDiJpn
L36HaYYKdiUncAHGqSd0brRMEdCGWqEXGdDuE3mspCA+uGfAwBFNEb59IjM+sJxr
km/aRv8GR9Gy6d1D673RIKl9IakYgyBiyu2QlUL11inMRmjtBn6+VyxANJWsTmkH
yHOO7XmigEjPvhn6K/W7j1k577hA6dNfNu1iQYkh9Km+4uSuyZTDrhmOG6S3sgJr
Q72/8DRE03h2/sIgAhX6b5QtUUJhWypXA234uIfs8olLLQ+7R8iGjOccp5s3IVO9
TwwAXl2vPFCG00EJUxECGqqam/f3aE5EHnqEMtEQwdLZYkZIMzR2A6vLVnkAfVqt
7ENTP1Ty09j7ajfnzrgMlqd3wvObSlpDQa5k7m3f8VNoN6XufDN7BlB9Pmv8ESS6
xmsAgyXrN+C/RSq1ZDNuGjdHAFF8bfTTKqKEcXZwwtykoja3Fl5UzQ8ehjLlsu7n
EapditqOuX15EZffO1iza+IhlNUTiWXA/x8o+HVNnXMijfIEfABcqN/zYiFEWi3h
trh9xTu/xsSI/z6iWtGqfs+zRBv9hMCrCu3FaQ+I1XMy0ej7dU3jgbAvzoVEU6uz
9Y+u4Au6nTQOaeVA+3ucDetwBN0aEyVILe7nVyU+zfIHCeTznhe5AmrnrHK1szxV
XJbhnk4jNltYS+IJalNvYsy9UDjqqf8YkbUx+jU09ByVSuGOUJO2YjofiEprRZp0
RjW6poST4HCAulMeqrlt/dCVjuW2jCmoBpIr8mBZdVeQz56LwuH89ftiydiNYcVD
z2RrqpxMkz+7HBVGiIJHc47Tn9Tuw3HzJlAwsLHAkzoN23Kr9/NiwaEuedgwLGoq
dZmcEWIZ9yMVIIYbtmOlksULDxd9WFpESgXy3cPf/qxT7oIrcBcuHiAYG9rqB9F9
7jdZCapibUDlNtzod4RtoZrNkK0iOdrA4YO9nfJ+ToRTIjv3/fqI7ONWGdmKOC1u
8IG5QJv6lKap73ZEzO6SJtAmDjnurWiq5ikkWSqcxXxngEjJ+O0k+NkPgzTYgz+p
r/kQIqwzjfZ4vJG0wF90svScGKiXt50KPLJ5F7M1IOXz+WAnE/PItSD8KgyhRj7o
elZp1NLMqzG060ZUKviu33pF6uHnj6aYmDxB5vvToFqIGP21IOVBL/AEFHxvIC2E
C9jBevT5NbpAmrzFz1om+4469su9KsZdksFGe/keBRZa9ZJAPwBEte2lQHwA5mF6
1uL0hEe1ggO/u0+M3DYT/qkoYYyWHdggWBdr1Xf9dLH0rPzGHCO39Q2iwup/TkXI
MfYzA8CvUfoZa4KokD/X1kr59GAvXFpp3e4TpqdNNgeXq2+2SQHl2ADh6DEimnL3
G0wRxDmuhzRIirAlZ4IS51RPRV8/oNDf/qC85IEm8CO2fPa0Xm9zx+lcaItCYrpW
W8mR04RRIk0N9M70pTE+UGD8OGtqlnppGzjjt+pilIG/EdjQo003FoOVcG8U5Lb9
IElGylBNqmSbTJpiYoDBvTE+v0PtKyybBAo0kEhMLElGQZP/S9000kTks1Z8boUN
7zBWCIC1voqjOYCV4DqiE6sbCV+stU6g/xpgV3ADBcjRNSypzbD3AzD5fI/cCWnr
5k2I+iyb/11cOczbnKAx4pzRxs11rpk2o2If1CuGSIefqCirDWOkKeVZBumH8OUB
jd7FyLToMsfYFA75RL13iYK40tqqvy4JZAKHoZ+SNlrsnUDVPhSGwPABeITmhB+e
kerR1g3SYAllrjhpwKc4dzjqjfAbPP6lJHotZtk9bnKaQPqVOuFE/SwoxJS0zvPd
NRRD8KMfIBhDpSrqOgUcAizIGVKRZJtMSa+NMxlL7T9j1vrJC5E2KX/xZxMaohHN
Ms8zg0djaBdh3vApFZYj/kgEQlpB76pU/0MrBQpbKHzqbFq4wHQIhOUWrWmbVC8U
1kk+2w08o//YDP6gTcc6S7XPL605O6WQwYa/wyXVmuyMgTfOC4SuTKbkpkzcxlrB
CIFi9W3ljRnvJp2V5ZvdAnUf+xBF/ZRh26dnyd80eTSo12sFDFPP2XJXhPo+3/oS
7qo7d/KOI5ISiQBHZauwohWDuQa9+TrlL2rzxK4ECP7NBbP+baVuv5F09wbKumFd
oEuoXxMA+3pD4JqYrlFBS6K7MwGxZ4DRBrmzMM+5H5o73gG2A9/oK4WgE4HxKGzF
y/xwoNLIYOjbeO6YkQT0+of4aPBLRzYlN4bg+IMx78PBeRfhQDAMOB2O+inYh94e
W6c8bKMeVVYnUkQ5H/MU3HLt0NNDf8yajFww7Xl53UoTUoi1a3oMXRyBhLdOCZfJ
/gD0W7npm0M15h0SgU9H9hpRnJXRbD0L6PEvudZ4p4JVax8docIZWpfSCuJHmkIV
AvZg4fsbapLYkY0zGPW4LyMrY4xO0YEDjpW7/DN9VD2iHMyTHmkrI7CVr4DokYpV
/i0u16AqsjrLNB3/9G6fhDn1v3MYZgOAuREA9EeCZzZxc9ERh2mLQhgob4JWZwag
Kx/t2NbNQlP3j7QdMjRUiAZaSClvUuIa9+G5ZgvHJ1/Aox6pSosRmc3EW3jQeOry
0qqm5N+8xrzP3tzqBE5P9I/W4cjJg73H4dtLfEiQsMRGM4pkSfOVYvexYnM11RlI
yVIshx5Ft9o+K2lLLguIWFjHmqyv1B2jn/BCgnJ51DpauEP1WQPFbx8r8I9UP6RK
BjtVzKEkHAfFpcMncoIenRL+30+JAXDVxVoxP/m+tqP/743YxfuycmvdUoi7qjRL
kAKhz8OFMUvQ7XcIiKUoI4RItN4t5/vNcmIT1HrX78h4Hj/bguexXVLDSa4rPXai
B1C1gkR9rROpbovyOb7o/tWllMLsK/4GIUFMmZJkNcKb/O+lFU+u7p0GaKJWwlyw
/kPyyotlWwcjZ2HSSknfucPoU1OuBx4xhbHIkDgG42B7MK79dN5RaDGvH4HyS5op
AvRsC+H5WNo/Pj+Tx44nabkpqvc9GP5b/bLirbzhVOHZia17DjDNReMFLUedCJWf
Lrg/Tyoxy+cnOcxqaDA0cZLu/pDY5ETkYvjuRjH/yZByvjqafONmaD+uMclY7AWd
DI4yQtMf0/xgGUfsVegdxmjqqjw8b205VIifGogvS6MS/jpYhz9jmuzzb9zwHts/
sWsWgdCSCRyvjUaQqjhdGmu09df3Cip//RnvkFusOdfmOmCCW9tONDbrOBy1D08U
ot0obbx8u/C8OCLAOOaucV16kthKHX+LaMR0LQ8gWY4RfWZk92j4tIzzCoX+HttQ
kmyk9VLE00tTyaqx9losU1tLPIE0oo8k8zFqKOz+sDU3ED4VaD9gQfqO1jR1i5rq
1uU71opelx7L7NJGkQMDPZkUYdha65sW0LuvSVSjMYTaGpG+cunYXiLuc0ydF5bl
6mw5bUGqOyaoHeLLEH3UUUenqf6y9Me0BFqb5rVDHbWCXAbAJTBanhIHXSB0kpHd
xIhs7VXDcHEpwiHUtZALKBfV6mefBN6dUAJIDjcAFrljC/XEmNX04xX83q6QvZZv
T0/2HkXi3s4Fe/nUkgBu5S3lw7P6vGFjQWosXRGiKBOh9icyfNCu+2thLybYhW32
BCTTxKbW+B21wTsg/4MWSbR0jdA4Ar6bz8ZhJfLbgSMekBVoElbHLJOsrfNkqerU
JDNq/g9tQuz5S2TE3VgSW5TyWrTA17hjXRNUOWae77y3SykT/SYovQA+wlO22B4f
a1P4clMBzCVWmFI4wTjuoy0fgqxDyIdKMu+VIBk2i6Tm+FaaPLUq8AHU8MuTJkfk
UracKyQtZA9EeKhHvPRSbeUrXN9oSg1v85U+e6vZfBTH+ROdDKmoJkXFZUieCII/
DCF5/iijU4B9jzbBfEsN0iQuuz8IlgBw08jVNkCcszX8DvZYWfie5n2UTiv0vVoW
cYfNjrXjI6AExHp86BHloeRhmR/48G0f7dSgNv7DXbHFmdJaS/G+nrDzCj/o25nw
Pq/WQksN9//ekt4pH/AgFjGj+kdYg/tVkWXb1h94ZsJW3pHS+rlRbHpqOEyzkt8R
WU9oFP+P4Pe05d5N3VzJDZzlYLxAkcRnsHZl5RcZGU0ZtnSMJ1j5WXOBfT4kUddc
7J9zi3tO6rymLDfv4cHLQiJS/5UR3aDKF9b318x33S7PfmkFREH7nOh0IuJrehea
NSCirol6gWXOHt5Mit+jIfZtGepz6rVsk/wLjtlhKtrzV2Lmq5Ix2YBCUs8uShgl
yj9CuFN8gzoKeSIWLnDe3VB60qUqnT/mnk8crJB3PPmbWDtjuSljs5kAcjbqVb/k
2ZZ5WPE28Q77wNbrxkMXfZoQMvAngIJSNNK3xHGl7kgsLIfIVpzAgoqvThbNB2O0
RR2icgkSapRLPzJ+RHF0w1utaltQhFTOF5J3sBAnTtju3RDiuBnEKRn2PeAUq35h
UHuftN2EcWGAO2PIHAUvWFHs1lfBU1/T3l4HlaNOaiFLf/e/Wi4Dg4WsRWIpEw2M
NVfMoAw/Wn+go/k65akvuS1FQc5TysuM4GqJERnq7d60jLsWD8qR3nSev4bJgx3H
/5DbxFUS2yIIEkyIz1VTNLPG0OR1zr7c2E4+/DxCtl9TqunUArJ86i3xr8/sSMl/
mVZSlULcOhwt1QHjz04o/JjOD94/1p8FM2+XZCrJHKNbwtkieojx6cYyn1d4ay/O
l7vgsnZacyk4lhLKr/K5763HstxqDRG2WTMEdzMHkIFxmu5QaSSxBaqqr+1LC6iw
IYzMzISoLVVxGSGPsTyNFiLzPmiZQLmJZh0BJP5zLBBsWs4HUPN8Dq8riekaBLVK
/x4BhQm0g7KeEH6PJwhoJVrwx+ut9zM70QsHGf43bgcXq1fHPsYBhMXyoQyf9f6u
A3ExIFq7L5sIDHvlUOALNCMw/xFXh9HK0+bja94HApFWF1tiQfzyqBu6e2xV8RRk
Oqi04kyC+H61QX0FUPz9HdsIoerlpqtfhI/cgqTiPvrI1/I58BJnOUorS2lT/bU1
BRVxv1H81FObgYBXMUzdM5u6SoLcQNwrFw3q/VWDz1Q3Be6kttz9l/dfVXx8Fftv
7VUTQw4/A1qDBYRg/tJDVZ0GS328onpFY56NZXrB5WqvHBuSj/m4dqyOSQuImWwF
aHiz+/F6y28rpR//5QDXuYylhvhD56YqpmXt64ZfttHw11uA2RukX/6FG84M71fU
wMqHVGj+H9LJwiqGMRBW7SYj7G+E4MCySPNc+kLnOA4wN6UqbrZl7kbhTd0mgZkr
vvHh+GleALr8kam5In2bTxSNVki7xlEQA/c0m20Zh9Qg+3Xg6W9tYBAe6zNAsubL
71RmrDrWpoEFh2u2mdpa4KFTGQEvMAmHG75BEavory0qqDQt6VJRPfQk7I9ikHP7
S40gSRkbsuBPI5+PVbouF8bG4XNAv3Z9lbKEWdX/UgzLd798Z4jLAWDJ00l/o05v
dBIWvsBTMEiAdLWElx9JnrtbyUczwgRA2dmP+gyf0nAhlJqGap4NUBrkMdCVwky2
T2LNRWUq177FD2/GGNfCQ11FfU4f7MUi7UfCVEjkuxi/Kr5dEms9roy3IagzioDx
rPQkky4rRFOSvBweKXUgpRemW0+MefvkSWh8g3+hh+WPtDKeBnN59wUnufGn+VXX
8aKgdg8rqa5rrPyLGhfDIcHpnFaj/XGngu9PtO1zPv14uMi2u4KAlMsEg05PAKeC
LV0ai/r2qcF4kZUfFF7VqJDWs5OKLf5H+uhFF8gq/Ojgl/7FczbU+jioceGPgcLx
QRCRaRQfCo6PARMoPZmezF4oGn1IyToEqc8xERjMe6bzkl2GFmaWKQc+Zr4qxues
7SdLYr7plN0Hzzcl2XKx1Uhy7iDE2CmT1DRkingFc1rHJ7jsfA6fKJSqUHI8RICF
xJOTTxdctu4pHxMKDTOsbUWoUZiLoZmkCKroFCiY3PzQ6hlkPkwqDyku3SvtGiMr
rgOYzdcYby3Tq1hiayO/U7cX7f9SIDiJGQLgy/36p/wyE+7v1zkzEzY/OZ0zxpLT
/gSkm9pK9bjSAn6ydhDwx4cBTYnOpoCS2+lwC64eDUd/nHRUUD77hBJqStaPJX5K
yCc8WRH+Lvkb9XY4sq8okooa2aJZnswpxV4aId4HqQkS5H/ER6kRSuWcRLB674ce
WZCXIWJgi08Uu4tn49qrB7dSnu2tf5459U5YS4Av5+RAVA2z8E3O3IMEdH8YD3jz
JxqqoaNE63ywSD4xkj0hnme/yq5sJsZ1TtyS5IrHqXxWLdul1INvG4jhOdFQUKkf
JIeECkce7OFNK3ZDIA3D4iaqDGHRwyV7rcS66ES5NKKKoMas0D9PEz2KajCaACSi
GtI25X+gdz6JGFrdyeEEUlhiHblR4Yfv/WmxoXYS43U44NutIUKPbGo8RD3iSNHw
BCaApHdvxZ5djYEZklwxwBxcbNutx8EZq/JK+vBmZbIUZ5g91I+apQ4g7Q+O4w4x
jJ3OSWgr+mrRr77wTynjbbyqRIgUupjkQFmzlZE9e7DAPHQ2AyKdEe/1nja4Nuew
ZpU5dBfWGjKgfbIN69eyqSWRLZwWkSB5PoRrWxQ4qXDzxXf0+SeNdXCBIhrXIy/D
pUHa527fueGMBJvP21BLAs3HjaO7Fhab5Uy305XW2wyHXBel5XaKiTpAwmETYTop
BdMHxS0zbXpZe/ypxuzZqmsIpPMzJbrYZrlYc/FSQmH5hImGnVSvaenuD6XsIKqe
3gV1i6RaVPz2pkhZN/QSqs/Q+ia5gbbZVx7hL6YqVknvimBx446IVqyywYvpVIHS
tDJUSysw7YuUcttBm9umiLxh5OZCqjnj31fAp1eqPfC0nCswDqILS5LZKLyzPxvf
IsA10DqLZ7NeaIUeSGp4wUgF5EtKirwL8AdIisuY71VPsthqdA5wHIsD8lKNn4mB
Z4lRm+V+C8PVRZOgRbxH6W6rqE9ifd9qM5252AUgSfWct3WDyFew2cyp90PYuTnA
zlMGVl5iiFJWzalyZXGQ883mSkRMMkJ7Em/Im5YW8w2lTpsstpNSS5vcgJ+S8EQ0
GGontgOcBFMlUgLKPlCIKBzXx/Ri1lPmm3G9zG79omh+1TJhYq/Wo/32lu5AXaiH
/AiwcvUUJlkbmi60ZXia/ljAHeIn6EZgx8qL80y9nHt5JfWakB2RQi2WGrmbHKUj
3XFg3Rrx3dPwUTyKeKIlVFZvcyLojK0rxHGp+yZPhITn/IvD4ZC/yhIB7P463RlU
dD4zUZVpZmRVHd9HnVAtoyNmfFM4bk0lv2f0xuCSfgsjTXMemxJqu7df6p9dgRx2
wz//ZCiAdP2uuG4hIstMbjabDU9FpdQERduRlT6mIcxXSIr8bqHRh4URDBUWlupN
jT7sfTTQiNpWvMCOjUam2zblpnwo4rbBIwjaq/mJxnivzpU+xe7ONVZtRHyEkAOo
GJBTnhiH/IZE2PLSmnjpnYvdgmDQk2xWNZPl8F36OMF+r4o3NtSIUh/ZUBzcG5Om
zxP3OTnkwjxPj82Lk3SrvD3jBNbcRvYJpk/XaD9LS0F551uXSrp+q/Ofh2MYNKgu
fcAHd5drM1+NEhEqDoSS12+8Ze5TM7gjuIJN86Z4i/cFOEnauJBOr59Qj3w9iNbc
CWbQ2qxjidyapkN/VLxgWQnAhUd25aWcJukDS4V2i3r3dp5+uFOIpK76AnWqzC6u
vUGwd6/YxVjX2x0Tl+8cjq8NYV62L7rRitZNXThJ9W7D0pSV3PXDxta9ncKIZohN
zaGE2VYnMCiGBpGzzhxB/6MZ65nZfkS7WYxfAyIfNDP6OgBb7K99GkkEuJ0vup2F
eSWfFqLBbtc1/uGlqYxquHcjqFaktZABxnvyoLQnIH//kXZGNbcwnPxmWd0kEnP2
aiEa1U7EZoPj37WwAiK1mwAndIjzDnce5bkPIICepcn47oNgz7x5fIv7bBbd9V7E
2KaUueSg9eBdNZM/R27DkyVQ5G8ILnbFSFjFLAtGakoMWgSa6Z4zAd4x3vkJTm0C
hrEz54eUy7rqmVfcrpKr2e643Wb1WODVkTraBno5Tb2F09jZeq9Ohw2Jxk5RYLSf
pT4m6PKwwCkuB032uE6QB9EK+06+T9StuCdNuL2XpwFgsWw95ZWaibwJCwIH1m9E
WdBUGB5rOrT5JBxu3gKZisLvxjOshVHK+R1KiAL7kANO4l3oNXIfE1jSR9HDwJhO
o2QapnArxDCLKBf0+WhqR3mYbMFYRHDU4W/w4t3XiTNbSWtT8/r0vTkbFl5/0M2k
UX+/wjNXfuAlnBsnDZqoJrVQobsXtukBBxE+6NTN/9b8bmZJI5XSgngnAGtddKuO
8JpyVaQejaZh4iMBmBS75+YW9H9CXvypjYDgThAm3/K8f1aHThy/2RGugqU4TBMa
TwhZiA0/mIYO05In3p5zLd9k9o/zb9QKLQWNL2p/tFzEUT4okPOqywahZk/rmce6
eC61M5PHGP6yRwvdb8wLjxDO+HCmCtRfbhPA+Va/IiHPDKhHp0ITslvMVyHLEW4A
teHiRoy32APvtPsXA2EqBp+Y6/mPgqnMK/sstys/od3XLO+0jhOGTqxRmqqiTNby
R/iIFOLs7aXVSobjowiyJS5FqfrT9woTV91fAuDbQY1QIIPpniFuS0RrIbkaz6MV
FHjcS+7YqQkGBACnTPTCQgqC2msZ3fTSnu0rPrrj8juIb9tSbtmD/bpBA85a3rQT
6+9iWPuTKtyeL6YoqF9erOVZpvccwf/ApUsRKLEtd2ylOfJRT7/cNJHYyaVgzLC1
BDFRyCrwxEXpnqQIhLB8idC4T28gcC9cwxo5AhDpynLITz4+8RE8hBmA5plgraX2
/PjHkbKJX+M6QA1J38o/CliPpJ7CK5xkJsJoZxRP6HvLJt1c5wKbB7UiyqPMWdl6
ORuRcOsVxTIiaBy3YsDoZphc7Ockes05vAWtDFct02QprKUWh6MjHcXcOvsbB/W1
ib2Ikz7cwEZgLuURdLjUjAVuwfws1+7fMCSFgPNzO9TTe9Q8jfAGDDW/8xpvy37S
QQl17qIvFcaJnKA04LLmSlHHUulC7l6lZz3pAIARqAIG7iYdQ46j0nUtbpviCHL+
6TQxSiyjX0j+nUaVfElNC5+MwSprFv0fiRuxe0oJ5mI4UH8PuQFCpFxLicTuqL6A
KFF/2h5CMPMCdkdGkAMQtK6JfqUTC+p9dTlshD0wd0CrYiJ8eUKcJKpjdcnczgbx
O02aLFrdjnlToKe7EV90rY7cgZVqGGvhBxj+3t+3AZpoxtV7Hphh+hzkLyfzPaj+
mx99sYvUlDwqr0jRdDzner3OVSOXXWu3p+1TEz/HlrAbtPU+ozmD9+fpIli5zewW
XaEkJG7o+/SOSa4Af0JQxLvbY7KprwuOjP+s3Zwd0QP/nnvt8WROoJpNoUaKnnSt
08AdM0XPly01VAFUQGy32RcOp9bYRouAL5Ov2apdVCKAnW44a5gnvcQMTHL74hop
n1J6jBkqAE4BNRH5C0xV9iqcB/vWopvRI9OCTZlv1hwWtoV6QeWgi7S/aHBilGt/
Js46eN41+Gu/yhVZuzR76HS7daIYCRjMc8ljf0AikG6F+NEhEt09HcIO2PLtP4uP
lhA+zt8x+T+OSvopKjYXKXu81bdUoCqn0yp9GGQk7udFIx0o/UOiu06btDgPzC54
N4q8FsKJP7hAdU9T6WHCbzJOmeS8RN6lNegb83zPjBiucmYHt7OaVpfc/h88Jx1d
+0fG3SFEtqa8b+c5OntUsw5kxOjF32VHNm58BDDk6mrSVpfSAhAGEGcjFdpV2wTp
ASIbptTJ78MGfpmNh/yoduQwaw0dMPajRdO4STJ4QSxh5dfxfGyVGWSRLaIjK9bF
EJXIo5jnaMhsOMApd/KuwGRs3gbVyaReWd9MjrJ4N0IoKoQyYx7aTRdRVgQ+qB5k
MC/sXeZzzApP01BKDo9JUzamNVZEkiBtWlAISltodRtG3dRR2QAdRm/MFVYPz0Uj
tB/49UrqS6SjqdxxI1ivb8/quit7uUeUWQ3iXtJjBBEsU1DbKM8X3UMs47zrAQ8f
8G4cBTFu/y/2EN4yl5KqbAkxZv2EfBfOMiXN8XM0sqRwDlJwP6V5y/uoSfvR46DU
X5hoE0Z1mXAmj/bD3RVacrQt0YdDtQ8aPGLdXTgT5h8BAh25Rs4EtRboR0lOirHv
qWi9/ixCrO5oWSPGMkrA1PDTJIaILBVCX0VSvyDZM5+kUVEtNkwaucghaspUTD2W
ejY5oO4h3ekaeAYngBDPk+rD7IZ9KT+SrGwiIFQe4yWCPXg4Y/MccIFi3W086KtH
61wdTvfa908BpsjX6pXrT0unCKWvRW+hzJGt3OgsvRtutS+/hedsSsWc/mWI5ult
JQjqS+Q3ZDxWLfq/TSbo5mTrYbAfSN8klTW76CwD//CAsH7Ge30pjFHMsx1fxIcL
wZKr+YfvW5wDwT3dUg7sc/MrhFcsR4Uw+4mxMwH9E8ZRuPj0J0dCPQjnXLHSkS0W
v7u6gamQsTS4lAzkfp7VLq4tbcHcze2/gg5p/18bBGZ31SeZ14AlxkW0gwq+du7C
qJihKEeGToSFEDHRSOHFEmWGPMiKD7lw/m3pgAwZL5kZKJQvvA0XoQrXzw7YuqxQ
8GKqw3H3cQiN9dab2kh6PFo3DySkFRGbwSyevSO8CSapsu/LLpgJ6AtfEjsQs3G4
rGM0i/0HWGo7IG4qGbfwEigeCS/CxHWYwnM1c4B0l7I9N1boTEL+0mIXOANghFbr
XqD18x4iEDRZK2K5yahFExDY/zdoiFl4jDX4N1io1xU3OaZDYSu9d9UefK3cDSPD
wBUs+3ZGIuLN8hD/h3OmrWwzOwipfE1XHkgK1Z0toeCEeu4InUWkeFqsd7XhyrBf
7nBuSG+/QclnnkmzCu1xAw8egRd1YEKfN6cnz687AiMA5BNf6clRqW/rXFb52xOd
iqPngtM0K/sj547bYF3nEN5EziKTHFRAy3/kzmffzmcXJ4h+b5et/KAKWgV3C/kx
+dipD6zN0vfSjN0hz7xagy9RECrj6tGZRTXsyD1TBDoRAjMl9LpE4HT0omSdsoWp
Q4rzI1WdpgBmiC3slcSrFmg5nGIrx8r1+oCTsKFQxmvrvwTSQsYnDzrqboWB44PN
aWu2k4sMJgDAHNa6PQQHBLrrDSevvv3GhwUlOUORtiYLpINj8QBKLD6aMZ0H0slB
5VtTV/txG1xt3ExtQzxpOl4ww4TPaGZS/hFDEtu+Tw9EBWSL8bC0798RpxY9rWhD
gaYQOX3UlwXHSUTvebTDxAGhCySR7BczSDJGLDTihODNbjuK62OFjpIeaBec/Had
C5LTcGMQOfjKZM2b4Cb5crqCQQGMMIyyQTGBHlDOkKo3Qt9hRFkYT/zWnGasCJ5I
gFL5bplKAHmkFBHohBuBJbarMIxKtGRS4AR8ZIeEZu/z7RwjHNkfIt9YuJoAfdc+
xhQH/JDWTZfgcosmkPAepl5DynEGu9xrbDNraTvK5vE0zmm2ItMdCr0zy9Gzj8AI
j+N1dGSUur39t/ZmS2IPe2sWV/w9+CXKve0l9m3T2x98o5AbJX+7usYdm552hap6
D9AR9Gkw0KBH/Y3TvvHXq3m306nlp9LuJuL7FO27d5GGoq/cUhKw3kZSUB9V2FU2
gERZG0Os+Zsk/EGBaL4WllM8eW7t8bGt4jze99x0h3wbWmd9gKzwl57hNHeVkbwx
JCDVKorDeP4HwoYcWcKkUKJTSE+vdF9Ol+hIlFB/3HWxeDuX74LECCdlWAy+qstj
4I/edno/tFKYVzxQ/PEIsIpYTVTsEZbiFKzs3G696tF7Mtgpo0c1YdSE98v2zgSf
fg7frYQrwhu+Jju1z7A7ggTytsYZY2CqOln4JS5/3eRFN3paV1Nmz2arH6G0JMk8
O2bsKuJnUCixapBZcS9YZgQAtDYqFxaRo6FhdMTAn/mGo2VhJPqQINAyxgyyc0kW
HWxTGIBVNyyHAQaC1eQlSvpW8TCfUST83BJIGKFH0pbu0st/vreCe0mDV0SKnz95
1/JFO/X0ZrbZ/j+bHjqIIt8NU6ug1DKzwEOu0i+6xiGtjUI6KveincwbhlwN0XDV
JQB4Ze/U0BQ7MnIb0sRt3Oz4NKwGapzx+PMlZJCOMZNGL0d2ZJMFBwSSoVm6gsRy
NYjU7Pq9anla06qGc8GqQreeqGB/NdxH18hqY7tAHk63iCEyIzlcZYYcRqqrA3nX
q38rwWZqe1x4USIrXwjGr4Faxxc/uQh03cvvG/MYVS2jVscbHtGA8cxHu9nLuf5i
A0tvlAo94k+e8YgaAEH/tE2K/ImdzTfwWWBJitKsNz0pDDc6RN9Ws2srnNF2vIl8
DTm1WnEYM/tPVMvVpdNRbg11eKyLV07LpUcjx6gBW5xuuLfF7slvVL1dYx8yp0CU
bKkOAdDCGqxotApiNQVNl11y0Bjtu1ztPGOM2hVW7+I8C29Ng75TrEgHjnUij/aF
VwzrSr9lpG1kLrb7LXfSoY77n/i6gcEy5t+JXXmpW3ATRxwg3gKJCB8y9ELWcyCH
9MaVD3tKKuK7W5azpRT1rvGZw2Odchqk81xugkV7v9uzuYFXqhw/7VTTZS/CGJ4r
PSpiektulg8KAbVw1Khi5DR0zQPNswh5lGmtiWoYl7ng+0twTja0/16FrFH+JkFm
Jc9aXR8LO6UiU/Ii6q4v4D9ztj0ZRegPRYxtaN6Y7o5528TQTIPfzsVevvaYrCok
m45K9ChnoFokieZMCnx3/57Tut93ide+svyso3hCvwPH3cCO65IeYrZEZU6Ee5N2
/jd31ZpwSiZXkw4HsXTgBb+IVfcXPxlsjZ0zdW5fOnT0B+sq0QAstPpKyzxlu3Y7
MkYhxSCDpkv3Pn2T+sC357CFO15yNJjyV5Fkua4fosdF2gA1Ri9o9cVOKC6GpGFN
ehG/UhJAWyYLmpj2abeFWLWAevP26NGr1QKxidA1unDD2aTRt5rAnNW35S3klNoi
mT6731qj/EfTuRik/PlWY8JxDrngDs5rCYCBIia+moHyY5yQWOkhxOUs5qcvCRbP
dsKwT89pILScWDtJV1YWcl4EXtWv0+4poCTuXVXsfUbTcBmWXw9qyDy/jLTn6ijP
1Cm7CLrdMHtqarLR1KzmVpZzMINlI7tDC/nQ13PfNwohKG9XtYPgcMM5LkMqKlx8
bsZeVpJaFf1hbXhK0qbynLZ/bHumRmM46WxMiIt1/WkgPnWaqlQ+Zyg8EGYi/YB7
zDDhOrUBJXslsI7FLlfWWQ6Fs7cIO8r23aDsYocfsXd4AqR8A2L4M2Vx5HnF7dxQ
c4m4+LJ6DCKgO0dCBJAPcnnGe3uSdkZqWqZzdA64X3AbVGrZ2vJ64LkIIYUL6G+u
beN3MkjlBu9pOkighJRtbHaceI/EXW4h1bs/bm4N6GQINwh9K8q6T4QrXup6l2pt
bS6/F3QyRxjc+H/62e61FC6fny4oWRFTSxzR3rIfdJl+eD56wi7RyoIfQTzUV/z0
o2WUlRbZIv1Wxs6rw+s35VphnTv73xkb+BsyKeBoz6ecjA+tYsCEmyyS40B5Y55/
Z+X392xCZYkK4pizCXNzE7CATOJgE9cCT+5qQ8h7tGsLjGCBemiNrC2cpjFfjecd
nz1t6/xY8/nFU3erNtq7sgzG5ofRz/SOjyiFBARVjKwtCmzKioC/DSdU6Uru99iB
oTlBybwuQLbZprgib2YujRYuaCoGD+s0x454Llz1BIhDf4EEKvQJY3rYxhBaiF5L
MQN5wU7lsmZQKrcqcm2J4SRBhOWcnaclD8JnNB05W30hh3zmUYn0LPOEvDooc0pa
MQ+867Jp3ikHafHDkJTjHhw5H61WZ+0LYUc/1DSby5UOrqeo6ZkbgjZSlu6sSXca
mRvhHxdwpCglfcWGc2TzjKhcoT2NqEReoxDqY/lLPrlvxLG/OQ75oG8qbIvp2NNm
Uogv9vhV7BD9F+oC2dFp4mgna/Dr/+6ud36nJRk7aueL+72U10fVWp0VHezutL1N
K76LhQ9ULQ9STsskbZnID/0+GInseh5BsFkDAGQZxjF/sJOVgnlq0QOIFZkik5Lo
XJFMRqQEIiGQMhqN5o7jzpoSMohusZZ/3kNAtjdhwdMLujWTId3Ws5U90WZKhgDB
ZAYf84gMQQDigqlaW5xnMzjU58YmFnOz6S+LeLUcnO4C0XmKChNZfWrMxhXTT3gI
iiU8T2HF7gsrokCjZmqaZhq4z5fAwotQZFIJ8WToy63Kh3sGiBHwmBWn990jfnhr
WgUmjJlGAjnB8vcPRRW0myYq7R02fBzOjLAroq02Yj9niV/VkvEyE3loIMtHLAxE
D3wW1TTanZcRYwCLOhMD+wpwLUobmX7QxG9iTr3WazWpt2I32+1cwP8pUjsBcuub
8nWNrVHw4WYIWthmBmBAUDvza//nOutJrDivpitStk99nCNPyddeBybGQ9pybf1x
RrJM8dn5HjL8Ik1vw0Hk3yEE6TL+5Z6ugW424HWhzUY/i7/R6KGFCBDxu6gtxMvy
IXostvdjuNAcv5CwJ8EOC0XD7qMxM/tFk60S9yV/Ksuw1zvmmpRpgFulelOF7fiy
EVaAY7Og1yvyXRZO6IGgisVwQvr6hNcgcbwd/0jNZnx18K/7NAy1wqPOG4reowGn
tB5dttp+i58CyneLnO9/6lVg9c8Y2hrdDr/Fl0OI92YoBNeNBLYKhfXZXB1SyuVJ
OiMRkD/vsyH8g1JFMxy+DeSd0zu3NvWBpA0KPamvSRBlOYsRYBowFXXoMZsA+uVx
P7mg3bAgcglQBLVIF53mYiyR2Y2p/wkOaPdp1vp78cGpX83mSDt+9odWjQK9F04R
28rbsOwSwGyom7bpwMnKmEsNGdZLTL5wFgtLNHg6hYxJrWQKyo7RaSN1Wbn43ZWk
1azTlf+7FN0FvLmBJHU0jJhTuk6NZ57Qo8y1XePOH86ZVQzXG1R4wIokhFNRfnmZ
rrAmp4FJtRW4hbrA+IYRHWGNiLH8GQj07+hBw1MhrUAUsJKO5ixGPg/8SUfQA9KQ
BMKeV2j8tbUxx8gT9uv0ZgneIur3iRP3pB0sGh59Xh6SH4d/Z44+VmZRlRtfHBIP
kx5ZrjkbXPzu4aCG/7uDuzZLNJsaXHx/oJS3xLoAu+NjZnKrAqkZsJ/UdkAOQhi6
wCxKNNSN7C9DIU6umA7/yQCDg7kRjEYfVulIaHuTnQR26uedkVObIsUuwr16COye
rwrauX/d9VBHD4mj+1gQySOk73qxPG/5FswmJTZoLDkVFzYHRkYKOs305wO7Goub
dJEiUDpVXKnmt5EcaHnxYpEC/uhDpeBz3MHJWZyvPiS/UuLLhu4Y4e6ySY8J15ic
MWnAytdy8CDrw/W5Hlgkhya+ozL6pdPpn3hsGKTGfru7iGZSiWKF9G6oD+ghppkw
huvia6Zo6hXRnSJ+zcpEVl3do21erSkzFTJtg80JSEaXiBnflkhgY3l0tXuGS8uW
d+EcFWf0O017ta+Irg3shYgpcK4ujfmFu52hZcFua7Yxsdl3Se68KAd9a1+TaCaN
juJtmp+3s+ZexacS13mKvYaFqz1VRzm0Jv8cT8RE09YGUpqTQp/03QzTh9vWNjWK
E+i+BrsbnIFeGaZ/Fq2BBMjJ8rpvROBKOJ56v1aD3y0I1ouwg38xmNU6Lqui/r8i
7eR9kyInSAii7QiQaUa+bO/pfEAiROanqQ8fI5PiT5HmJXtZC9X/w/8Jqn8EpwE+
f+HGFL5zRNGSNYC/zHXrl9KuVV1Q9tj47wYrbSVs0/iZCiwlRWNE8YLfA66uUHl0
PcNS+ewUzpZBGUPpkL0Tlt2knWHa5SnYEWkbOZCBPv+1uUWTqBNlMtqeXukC2usN
GB87fx+kY4gJ6Mqx24yOJ54xEzr0t5Mveaik7ALYO+ZzG5VWxbf0aardGtCW0JTX
5JYWRm2+Q/+2aWxQq18iO+PbnMMgKnPPREawIsHY8Ah7QTHPfidUrMk+uD1GMaez
fuD64v4uBvKbvdJASv9B3AawpGkKAbp+01Bve/amDObsx6tJWrGXgsm9ulcT16kr
E9RcVdUPu88jlmu4M09C6HIlAsMISaz/3ocLU+kQiLlHUkIHKu8BY4gjYMJ24RbE
NKtjE2P7a5PNYjC5A/83uFTangRXt6MMJQVbvDxGM25hA3SzWmA62Fu3HFJTIoEb
fIoQVfn3Cn3QfXRl08n7HbEKtGFUTLMBmuDU0ryg+5kKedETHr/rej7lnKrEE4ZW
g1XLkGI+ygijNIiuIOwQ/sdVVCejo77RF9UNxfmL4kwzDpkYSNc9WFjEYcEMtCzs
bFNwkJMbRs2SJ9vPl75PENJ7oEhWts9ZXacq4PgFhmxZokf2vBb8nsk6PosQEj2E
vtyVh/qYc59u/sLfQQy4A7MQ3F09e4CTbtuOpbmNfJssS4WX6jzX5diiZ5ijR3Fq
URVZ7/YkKsYyfhUAYbzHla2ptjmJfIABV9NXuKTtyu8K5g0YF+hz9pE26ZqfU+2e
uxDycduQeynBI801AF9eosq3hCM5sq21saWKrt/tkEVHccU/f/TVjp4W7uh7Kt5m
uucN/Wp2ex+ju89ICR8OFR32Ju4mfocDNHYtz+C9jxu9MsLTNM7f+2zUAuct26KT
DI9F4G9IurwwF9GKuSPOJW/LzwwyIs9TMX464tlOFxoEdZsTFDtGCaCt2gR14P/Y
HykMQnUZ7BRzHK273Y9E4DXWJK7t3sawP11yk5d/BRvBfp91x7qSbYz9R5jbEPKO
Gz84ZF89yh6nQhBKtocOMnvhsQZcgzdG4aGdypYQ2EqxTdo4+NN2eeFp3NV8K4ki
HdIQT65ZiFxVT1rovjkMrPWyNEz0D0+JS+metem5EDXQXd1cT44WlhY8a87QbaIi
upgaQUF9OdwSV2TwQ6MiKz0RldyO4g8tgqvWKweGWfGZnKWf1MscJUuG7nMTOD76
w1K3fso9x7lEoSnNOCX6PK979/xiJXAKH9PGBC+pDt5/p2sfpdgmsrOJaNDUM+ci
Ktep5tM+4BGTXo8Z7D/ib6wOqt3uEc0Gc7kaMi46CzZkf2Jys6ThMG506rmTlEoP
UGMyK6vKl1fnKOZQ5q24LXnalP5QGOjLaMH70kR4X3LoYf+cLZd98bztbfz7K4EX
TEcseto5HylLbaBJMl7Pvo6hkoJEz/pyaog2dPXZdF976+pGtFX2isK830riyo+0
86ZmgumcEKnVX0r7cnGm4RtMcTvzwokLTsdOcv3GIyXSz9tKKaDOfKiL9/oncqYa
MiaM7lYoOKubISQE7hO0mNThlAN4Nxpqhzs7r+Iq66bB2Fv3it3bSFemSHVQNVYY
2Cygo5ZZ/mZ3QE3IXcNp0AUshkvnuH2y6Wy270zRidhuhELHQMVwNBnQ23h1zxt/
SqaAvqjWbJkPDbvs6wxpHkRYdbY3fRFOajEszaMzIZ65p77a+dPR5y8xN6hWZX3z
XxkBI0lfFKCyfOnPFibrBCx9r6b8wPzOIGlCWe+Ua05lDT6sCyRPKB7VnSKpy0Rj
REQD1VsZSvmwt54HN1z1ryn6a9KEkYEZpCAT4Fb2fg7PUsnlWUWw9SgduGccOsH3
g+qX7SCJcgGJLN+LmifII2pbCjCkbCtGD/cGkv9xdtT/YtvnIv9aBJXCB6rJzsA8
h347JQDw6bX4DAfK0kqhMgsG31mJXwHGv++rV/zFg13d3GTzimKzzt2PWoWm53wO
hqEsX/ihrPwWxd1Muj4l8rwIaFGm2Tw26wHN+DEhRPehRZsjimeQ9xJcPL3nSDX9
gVeF0ZkdGaDMkE07MgVF7XkItnzwY142le5teZO4pxPQhO38mOBzgd6VmbvJWK6D
MWqa0KgTPoZPZ3QivvuMGis03XrLiSDSBpLl+aUuCAzhqhHFqrs5V+CnAZZN/cmx
Fb82YfRenwl3i2oVJLfViJHgi1YW8Qwn3ZGMG07T+0kHvkgbhUcsijp+wHRgOII3
WQrHCVA90ay0RsWMueq6YBNhBa+TlI6/75L144qkuVjTUCJYpkWJR4VJ0c4qRGV2
F5rSvsiWXPoEexjTKGvaigEOZRIi0tSGCodo86IH8oBS353XhySJmaypEUp+L+/+
2U4sItaa2h1a1u08yOJTXwpUMLimDA9LxV4wpTdAHv72tpRW8AziylKTRs/qVJCy
9E38MkI0MH2BB0CvxVVS+n7xoVi2ERAv0ovKxd6kK+HyR6fi1d3LgrG0qoZFGQ1r
fP9byQBTdyBzDORU/ecnxTrY+GMys+HSz38Q+MLYHXv7611CerGJF8uv3yHPAT7h
TMLyRD9pzX+tJ5yKsoi289k3h+m0dkBlQPS2WOPOsbRdQYAQHUnBc1p6jIQvcnFE
TgC/IuIlldpmhf1EgcgdVwhD5RZDDlPUkuI9Yn1QmCT+k7KAT1UWhbCDF75peGqr
0B46sX4jhyFT/lfY7Ym/e3oGHOj+oQA6CSJyIJd3mm26WHjZtTpuCoMuVx84069D
cLZnUaZH+QoW6rfJFT1YqVHwlbduHSqujYq9yHVr1AmimRldVoNuDo2fPDkCI/GS
ejpZM7/wGi+unbTQtJHGOWy3fQT/HzhKAy6lxrjXb3zjBFqNRygFCyoojjxxnDjI
TdFRWVfBSi6nOVxC+unSW+Q1IzX3ftbzsQ7l+plZKpJu6xuTHrdZVxtYKKBf+ego
xl/o7HdGzBqeJgryqjKoSdGKj7Es/4e+j8chGcJd0b/6R2mta3kYrWw6IGUr5wlF
A05imQyFMWTYLWt9jsbA8BkO/GiDBlpDm0B7GvyVd2+K/p7zP8M/akzQ+bTotfhb
fgwrAlLKXHka7ERMNMl8R0U+e2coI8IBXyG2ElOyeO3ftqCfVWjVy7zv9R9iH4Kx
QaDdoeeo8dwxopNR2Zx0Nup12Q46HaUmPwIknSQbRiFlEx4D7Btdt/BoGasTiQqG
pvIQznPceboxuxBw+OGP5Q26w81ifQa8JNs5i8cmefpRBtNqbyTZ1H4pf1FpOgT2
jrZSKOwKof6wLKFE16xP/QAOtxU4rSbsd/zMEftUheosVcURvIrvtRRvij1KPX7z
/xu+J7oGwLbMOPa1/XRrB+aqD4Ptxncq3meT+jO4kwFh4aQR3qqHgKpBnOrq7Eul
rOddQwAchydvZEsSimzaK9HzzbVcjreP7dv9DlQurNw3pNDWiRQFo4Mf+zWyWhv7
JllDDpOyo8fK/2qffh3LLBr0jqOVgIoJs4OfC9pqP+5Gsdibb5h/5hsSUnavPxfK
SBwM2mbVfXGZ6KvD7YxCI2oCysnhbyir6x7v+OQ1yBzVh0Y3T3xgmymq6RW8KUCK
PQ4tl3/BXLJtd3rwPoMPHZoo0P2rMKNmXF2Bz4RpOrCD/w6MtGlTw/SCBd9eEsmc
yHVj0Vj1xHYlrDnKr43jjgEL0KlfEg8Ai0OpnnwcfYPZadPVStozy77TgfVdhhCC
74jOvua1gdWLNf7E7m8eSZ2GQyIfn22ntQYqZOJzLJePzMaYRx1cBLxd/8+l7w4b
xCoEMNtwb9e83T+lhehWB1iST8F1h1Y/WbIfgX30I4Q9avZ+3C+aD5tekb86F1dT
sfjnMRVdPL8bJo5ymwe8mchlQES+/BxNvb3C/BlF4g6eYnAj5BgYMjVANUPmwKRM
gL7ZKaQB5DMd8eBWRrM8ojofO5eXCAx6tO01i5OCcNP5PKyAruTvbo0UOT98sITT
whJ4PJzDGr9pL+kWaBffE2al0qPxi0eOj2VxVVDSzd+hx2m/lf06UbdpiyRQcFYQ
+UyjNA7YdfBYkd0MgRKktI3uQSiQsq+m4F15FRGYO85GG7T1xN5WUGgd7upwPzys
MtThRpTS0aLhmjaU6fJHs1d/iReuBXdJsp79PFlN2QwJ2bmQ/89U/DpajXH9O6EU
7nN6d6Nn1TAjpAohMb13H57T4J5XDRMjg3bIO/AaJxIEUav7WPQt5bgWOZbidW9F
OAzJv643uQ9mDAObnUqBcbpSS++STeJ2OmrPWSJ26V8r5+g7tXMQcc6wVk+vHN6j
0uSXG0qbPKe04A/lPRo5zHn5WGMv0OZfbYnY8fiReEE/GAJsFVhOMAgZzrYqFdaa
9m0+DidQ9bE8qtm6u88ixy+TKQ8U6EXGtxwOa5sb8zHuiIf9f8PHW7ezG76IQrVd
GyaLPtCFHeV6+aIY2S49E31l9Vf/TVe89pXhPM9lq8nYajtaCSsgGgB+NlbAD00e
qTdhA9JZHkTiUQuo4WQ6zEkEBtkinGxyN7OcHQNnKp2cs1cMnWUChpUO2Ihknuou
jaqBIJRDTzZQ/dGmtZm9sj0rfp39ODZNm/a94D4PIGF/agGm3BoCCd07k2Y9xcML
BqHg45E4PeQZ+TaWnw4aXOi0ZKo3WYqDKRX1xlrCzAA4djYwCdWTG/H8CBK7wF61
wKJ3Bg9qszwjJyevTUowUrLHZ9WrUmcUKlu9zeMNgA3DTyTGCauiBIZR8jQKiFs4
klThPzNVu28Ttyu4qyVDuokKcjjbKpJP04VyMaqgVL2DAWahvjBqR+2q8+U9Hl9b
N9B3HLfQJ9EIyQgtQVSRvGTYghFZMLM+cGx3oNRMSwFNyb/5hmzAG3nDAeznrP9N
awHMJODiQ+fUu7vmklp2sJFrd+jOe9l+8qnaHDgrrHq/g5Z/8hQz2PWhM3tcRfFQ
Kdl1LzVj+3eCipw/jTaIWKVGqobWpctozvpicDdhLegvMBdzFW5VPhK40p3gCrnX
lhU0/c50csQ0HXXpCJST8sqpwx+j3ewjkmCwA0s/tGeq/W7k9K2yVNo0wLnLs+g+
QWh8n3u9e+9m7tKWDH56dglD6M11aKMEkTdimFkEyOGq48cbkdV/ugZU4lnSEbiW
9lRgG/YvLGro/4LW3CZR4v8kYWuVvGRA9f68uCoTZlPImqopxz8cHsfkk6RgqWdq
iSnGs5PVwLJVlk3adlXgBdQJxHhPQAuv119suvItheYvaxFdGNQioJspHbqmycK8
bl3LMspX9qjdjtQewcgS477mkpAcENYABCvEF8cMyK3DKq9PY0AZrpqdPkdI/nkO
FdSx3IytAppAEtzLUGkJLzNpZmT0wYSId0OUAvfV3rdFPI2A9DCLrBcg5MqJNK5P
2NwhPH9jruC9z9RYiP9Kt2t3gGWE/GCjg9FAyY53O/V8c7yMicysZgfwUV7zsq/H
JQqp7srEGR5H5j8Q3q9IugH49GIt+O4eSx4b5a2Xhy1S74vrGhB6dRwZJEpH7yNS
mgrCUc5XiyNWYm2fmCWwuGhFLt/tUZyDHi25p+qyPbCoX+rqKJnmyG8b1vZGudLd
QHAuqQ423NOqz1EE3OXPZThlOk8Ya9nqwhxak0GS30kIDRmqNcwEjK/YzJmziNpe
12hl9awySLlyf35Yl2t2BR8MXEAJyxS+Mh2rEhwjeSKKfPg3NQzWN6tYuv8THXkP
f3n1bZ2jTy8sJAOtO1tydXZ4Am9eDJmKps3MNfay2x8BIILgY/vHZrAHhrUS4pFV
FJUixMGIQxD3edSEgsPFThHcXSwPqE2wDw5jnZDm6tCkTKyI4TcP0w7wDinfsve2
Ga2CHRAIuhsa/b56H+9kupoKudn0/+qpGwmuB0+8wkfrasLfWLCPd4U4wzsNxoJg
VED2J8+7LmrNF2Ba2ZRJc1YDPaX5aysrIennQqtyM8dfY7oA9ejd6AlJm6Xry3/L
+pd26s8K3jSlIu4rQgCnl9QZb75VgQeS1fMBHJfJUvgbHwfGGSXjF/l55jYmKdmZ
KawpHrnCkV0tcb0BaaPGanNQ0wPZmaMUUxtLxxtOJZpP0rQ66SDQnnuRWmZfTgge
nx9CHQG4dVCFvPsr4uTvZp6PP+2az/laiCue7tUeWE1teDgBy1kaFwJJ5CGjkb7y
D1FhDFA83B6yXVu/0INy+O7Cuo0nQy6or8TrgBpx00As0KYdkWSz7j4E1idOeYdz
xZbE3vSQpnPZX0SxdhZrbHbkcvnErqPT8veDdXY+QNExDEKHFmNYmEoOUXxJ3RLH
/CFUrNjGxf2fr4T1kIBFv8cJGPlvTm/1iHwfd70e2sS1HfyWM8ygaJQb1rjQs5+y
w8y4q30tslMLLtsvn4iEU8tLbTX06jFhvplLnkCHMuM3FIG0TUnINBPrqtvs89h4
EUQZfRUiOO+Lg+3DIqECOAQtdy96A2lV7JL5uhI0ZScbDjzhDBUBZiDcGbonO/aN
Bc/tFASn9wI/SwJGp/ttN9ogWf5O1L6IjkvyNli1ukCETBaoBj+H+maNMSS4Wz70
XPybAoDETbrQbD1C1MT08VT2GVzBK37L+xLNaelOVppO88hJ05BRJQjLKz9opsaE
UewEIAFBm0axnK3MKaXYhI/JaFWPflrJKI4bHsY4DsZdCOADqK0WvTwRPwCH/O76
EcE+zyPjPclV6ZcBrXP6QWIRq3t6IFNjB47b1i79r5N5jdlFnWb572bKX9fQOGuT
wQ31W2I+nqFJ9yepOT9uNB+Wb9kEPX1wDdP5zICIGU9TPZ5PQyvQw6OYqsqNUqnK
HTrFwNFwHPHD2nio+JtEP3Tf0ST7k+Ji9uVfYNlWWKVD5FrZebS/QOHrmvC0yIVw
C8juMcxMdRO03MgqOQqrGNwpRPZHkjb0A/WxAj46L+3ejS/HTEV1zf4WDxUVcp/Z
4r6jpg86HVc3YoGdWH2qXm7+3Pb+nr1CEE0r/9FkGWQogwTt3Y9UD669TB8lIWz5
3fr7HW8jGkDOevLv++DJ8dIMcccGaQ2+UKNvKnInug2Ekj5Sn9qO0yWa16IOd46h
J7gGjcmh6bSwzB474DPeg/Nz6V4kbBkazMvIWHMC+EvwMq2KsvujjusTvPBID2Vf
Jmdi+W1amZoPBYXXSLiAB2p5h5oMDseo5AZ8BF5XvW8teD4zhPEWMBWfRFfXslAP
vX2kWpMxjntcD4iwSHeEt/dyjM76uBMTs9g6aGnC7o+OvvRiHx6X16ptclP3yTEC
JWPLB9SPLWR3BNZqEn0rBoDz6SHcriFMv1rzkmk3m00KWxnNM/oLAL2JVfL25UPv
8HTngdqP1pJyNs20q9aVFS31sal1u0DiJf4cAN1PC99U5TQsZhe1VcPWS5x2wAge
Vb8W+MD3WiGr7LI12BIP8aQEhKwHktvSyvacHCoiEn+tH3kXKKDGvpNHcRai9e9S
TaPeUuRdtIe3EzaKvlT5IBK8SlqHvXagrfkQf0sDSqqSrsf1RdXXb1AaemNmHoOC
+c4pD0JjOl3agq9EpvAYHJhTAlQPS8a6HogaGYg+1O+RRQGM8pdzKf69rpGPGFE3
/CtKjh8QQKmgw74Bbd0WpB8dHPulypL0PO3cVL1+3VaAO/zO2CIfdhtf5i6H7ozd
lZsmo+zg1OQG6uqHkWonY2D307WMY1AY9RQcecaKGfXodm0SQ3kCOLRWt1x+wxbs
4RQmmcYOob7ly0v0c397mGK2DN/xI6uqrmwF3Neg0Lrc9x9TxcYS6om2xTugqzu5
7WWiaLJkurmE+m1bLzH4ygMVVUrl51vyUzNDIsjFoC2g1hr4CCsyhXquSGCKG8DM
Ba+fK+b4Z8lnAx1KOUUqorNt7mkSbfMYJnyBlkoexb07na8smeIXPcgkdsB2fUFb
TKUBkv9fd76HK34pNzkDk5Lo9UpFyDQBR5AS3YVeM9uz2zKJlWmENvmjwJX39m/g
FhP5nZqGWfvQCQ3k6UlEOmtWkf8svGnHoDSg2WT/WuMIi4X88WkJ24HBmaqLmpQ2
b5Tqx9yD9NCzzWzixkk1OD7icmDUE/rqB2dG+rWyF5Hf5Gmo+2Irqy90VpY12xiK
um37m0hwN+WEWoJkPdmt6h13OFDkx+Wge1FTNC5zNgniOgLcU1MOkr8a1nV9SfEr
Gy2jkV5fjay+iKgJZbgSKV7HqMwOqwW6cPY9jZU3MAufO3A7R2322f8JWRXt6Vzi
hdnckOkXa8kP2iWXbUgQ5XHx99CFAWT9a1wHMjmSvf8k/K9tb10XDbXZ3hmuRiOh
dwXe0bYE3sYW2OPbLnN/wK9hjoP2xIqwOcbcRLMnqsVi3WTAWRsordMTONP+40//
Jlt82EzwDZJ9LH3SFj+jxzCcEz22JJe1YqCtFIcwmlAsvXwprs8mK8MSYBK7evOu
hGEVKcN/t7ZQWYXWyjC8L5vO+85DiEHgoR0607q8seslJutEARVoKr0cmfeUzEjB
W8o2DlEIJ1+hlA8a2Qs0rL+4dSnWJcjt06jrn2jwhe6A4a5pDGWpkCzuJC5atwTJ
N4AhHFqxi9YYxeAbwpw1xCtWQioUpcxx4d5C6RNBI2HOkbB18FDP1yqe//uxarzN
8nG0Mz94CUE0z0tR5WPxCGlNHTaN2IA5wg9bgekalFFKPyhPRe/C6J5YbP+qzrad
41M3kj9ZoVF187wJATTdEsalR707OaYisASK+3T9ScUQEoQt1yhxhwZfK2UQ9zG7
DUYxWfQvQVFnBSNR8QO9N0WYYR0SNH3OMxRJQpj17BhDiBvRALeldm17MiKAqCwC
Vr/16UwDXm0MfJOJsnjYaZmBMibOsIPHJIdHj2dN33IgkUV+8984MWDMawBjCk5b
8d6yMUbNSqNTECOAtrME0FRRQLQA7/qS1aDZNdzAIugxc19XvQALOD9kYYhISeHD
+0N+YbOyQdqsWQO3f8sletdsEGWnmki5LQdmKUXNc+2zlzbTW3oHeLUlo08LZIP1
9yOFdaB1kYQLtk7tryhphTLbR5dvIwG+htZJTaVvCZaxSpXiZ9MHfgLLFBROX1ec
LWgxL2Kg77hKEzezdrgh7nrWA4RCuh0GIMKdczOvs8gJdmPsPa7BBlTOvsUcYXRf
J3eck+/ztxNClNKcv2pRDN0lqkCNeR1twytql0yv1jIQLvtJmEnqjxPaUXsurZzZ
V0UYg2GqU5HbENNNII6+Dsl6zcqBPPpKpInHzEj/gLb3NiHh7TqFp3LQqyMvsk9c
yFD1TsidNkv33Rw8apTiRQpNBk6Em4vgRc2DTWCCyWEvy2eb0iodcQUmJd3NTv3C
DsbG+cHuK8LXFxbVEsXzz21X9XfVaqH9SMsqOxCVeSTPTwZDCa3foUT8ueitfJxD
1GVNWL1luFQo68spjL0oMYIot8l9Q3Qg+9V8/Uw6tJtth6Nxr8aqt6SmrCkzroZF
zQvjvmFDKWi11IPCo92PclN34Ini4pv1dgAWwMENxJhkaSKy7Gnj7x6/YEtrinFW
O0mV2VZ04s/gzCGWNtyE5uEm+/cdZOWZqRmQ8VJfXz9ohLyEzMU7JuOOVdo0rGml
HAJoPVlP0U6Lsbpwg2IkJYVVGbE9mQ/QCgvIdounNwEXVt31aeo9bXK0Gi5YLspa
Tcrale/g0enpKgzso8AxVWdc46waZPiOhXWNp7VoN0juNxevpG2GVOMRfYmXc3FT
IXEdvhz9QW7g+HHEmVoii8Hx6A/5CUuoLUZ5DPBxtLp7ybmeLx+hCUzxeauHSDZG
sY1TYrz9s6+y4f5P2qvffjOqYKbwmyKMkyw93uAQ5bDKxUYOJAYxNrzLA+xUji/7
/YBeWvpZOjun73dqwPIYFK3xceWFHi4NfA/stptGfa1rVx5U33MNmWjr8cN83GlA
6Csb4lhoMnWRGt6s47gjZXVOw+2tWHASK4wM7GkLhkJympBNcE0G9FLVTWKkf2/3
9BDjxN8iglxj/Nh3x7TKgC6WuhW3/ftwGjZAym6rn4SL6hJ75JCmt+4OOiiwTIDF
m9dvXW1z0UI0Im2HZ8164szltmqBw+Yh1ghHyjdvVRysZjEd2AGYl3FXeqC60Erh
kdFtQM9YKLNbCui4+cbgVSf4dqXvTFNOWuRYWRJYFabiKyFQAYKfbGNS4/JWmKGL
OI2ecDO6nkqeoJwdd4wT25spD7Hthqfk6PZ7xUk/SBucTW3oPY1pktkj+O3rVs0S
HmXbroVVYNgBbPHn7EeZD7fGuH4+4pEozA4Y8/lUeUtZKEtyh+jWSRYG7AyWAnKF
zgQRqY56vsSlsaBkjIjoqDT7PCuaZDV2IfZKNQE2rucOMRo6jPZun9/odUQaAKhW
2Fbfy9cfdE7E4vGXf9Zc66Wk/hFleQlv1C/DRSYmJjTpPZOxKtyuEpncxXd8+VT8
qPdxFAUKYdjjcc0Tk51uPZiDwt+MCYI/6F9nt9/ggBDY8gRnP4UKnX1CM9J60+4V
dRePWDB9YWXQ5j1yZfl8RW2bb4jt1FzN7EZhraidkY+JTFe4+AJ7EOLjecA8oPk9
Tm6LU0hhat9+3cAZqZP3VPEqC3L8vdfFYPOhqv9rpHBKt6bilg1eat0MbO32TPYL
DuitYbcoYTgyeBVmFm5BYQYKoRQq2cSvSCpAySHL7NvN792UWJybZPwiVqTgF7+e
jwYhZd9B6QpIZ3pBfXYfi8RG3p1/bLuGxjKHlWh8SHAaG7zeo5q7AU6zoi/sZR7I
dWSS1OSwu00sjl7l8HK7roigDHRJwhGDB+X1DczOE4KEd/pWEmaBjQWNCVhc97Pj
g90AsNXGzWn6WnDyQX9IIzKbplLIDldOvAIk/GG4gYiNW5YNuQFJaDC4RHxQoHo6
sZ3S2TwGJeIGEUWtZYXqi2DfFGMKlEFst8qutZnpqGZSLgOY7YcOkMHbN5NZSsJd
Nx9lVeht/EMDFl1ed0kQbrEA+TD7knGczOu+3l8GXorZ9tPX8ter012cL/ViWBde
0eSIvmF2Zk6fwVNsJpFimjWN66ZXnWWumuKhNnNVA9LiFVrFXWUJzq1N6Fp7jJ+Z
Y7isv6icaBJf2qJRqoAvIfXE26973QFDU2siJSrcDgEq+DTWpmv5EQXBLFIOlxoB
PY6D7W6F+dPtqmiBQJQRVLYDzlOFP27k9bPts9WwxJk7BQ9Z8r10HoSbJq8hnmzB
pkmxiD40hBveeC9mcmyEfS5s21TPPI4nAYWnKzLWQ2bYeHQyJBRBQypc/nKxN0bG
Z+bXogoo3Gl4tvoYiv9AmJkIm0Wb3TVIkdoEuyL8Fctmgo7bbYyt4nQbTp6CGhCV
JLKQNhzoEFLuibr/HdSZJV6p7VPJTAMk385vwksGm0cF7Uyew8uZXmLPNBOXS5r2
63nMJUBboLIklkMPYhDqA+Go1OOZkZ9y80ejK8yYrorpIjz6AYV7A7lkz9aoWRLv
tYZ8qrjMiU5yRAcvaHi3GjR7UNdH1E6LPMCLx61I0l3do5jXv1ujO6p2oNlhjHPW
pg2qJlGZR0Xdj51CfytPoYceUISWDP1djB/HCKHOtP7SKDoH0Hd6PJwdhE8GYccT
iGt58A9zsSSVoNB9Vhp7UWYs/Jup2Chdp46651QD2c2RKzWtdrmFOVxkmyiFx8zj
urdynALAKYk/BnZnM70PaPeAOTlzz4o9T2tGvwYp1iplAkAzSjAZpVKfF+KFjd73
Ynk+3SFrnQ/mN36VFGX7uhLN+AhNAm9FgtOvPGP0q06denT68T7RmQvTfelAT8aw
UG5K6ffzZsgmisFfZo8U8jaIP6cHdDXAL2lz68u/esA0wPk1ceMnggUbI7p06knZ
2NGt76dG6Jkd+5tApy5AWYVVjJJqaKyKS/aB/czAW4hF11FbO2vrGGQUAKf0lCZZ
j/56518fB54aYIdw1a/OWO9Zrt8oSc7x3H2YkV1+2k32yszfRK3JvJ6fNuZQSlRb
hV6ZKYtA0M/gQYxs3FGbi6pnyd0esANho1QZRG/F57tGFP7+q5anUTg2AZIwIEf1
fZclM0QPgL9IzDmj6kXrFAXyJkHGo1B1M0BEPtSrX249EVkvauXDxGjgvbcEgd16
w7mab+F7+7JV4/hN5DX202ufjMVixa3XZrvLtzqcSa1VX4F4x/N0CKeifacGpeSF
QiZI9ra0mAUae6u8WoDL1iCQlSqg64T166ezAFxe2K/7oGbmxFe2SCApwpd1p0kR
5No4ksx/Qkm4fPAzgEwlysJ1Rl2uGYtvnqF7RlFxdqpdcCiMpXXQHKAUl5XOg6CI
L3SJDhpIsm5RomZb0rQNHGvJhT4oUNcfQBF/9xF81N2ytVYDkY1790E556XG90D9
Gxx2qs2n1U1/jT/1hCJwi1R7aYvRWuFLESESxYyAhgA17MODWpoqY+cL+VPf1Gii
A+E03naKceL6KAjblsQXFLWnyHqPRvWp8e9iXo7SD1beBh60FqJWMc/3TsdlhptV
2p+Gm+3NYsYNBXhkAGxCVGJ3MQhHKeFNHd2NW+3jX4VX0CPcU+ZTrJQ226xR7Vay
Jaew0kE29pZYKR2+xPlUkvGzU2RhvgJPo2in3Yvie08bJj0Zzikb9xeGS79bgzr4
hi4p3icoCW7CqFfgCzEpnSgD5zWZ/CIUquL2Qh0r5iMn3vyJ33z0et81fqwo16Hi
Y90AXRModSC53oGhwRR/Qq2Oau2QWIb25q00Nu6ETOUbqiNxjrwBuqvZuHuILFHI
M9pGl35tv8nYdbqVos+NTwpZwDnJzKD7SrjiQm7F90JayGfRsiIuBezBUPBqWdcC
J/nQwwTK5uduC/Ca3G5Rs2FGZM2aFQWM31G/xJhALfMkFyMS2K7oDMVpkT9irZj7
PNyEtGayKaQKWOCHDmTSPPTwowDJiXmb/UM+vp+uPmM7shtzbSmLq/QguaHt/xxu
j830272XHynxhubaoxMYuy334rpBVX+cRiL4sz4B6MwzqO/VVGMRTcf55hBbvgS5
zPZ/jfFAsXXURaOOKW5ps5JPNY5fNQruLJ3OsZd4ddvj6HkImrN8/BNsddwFnDTk
+84GIwhrAAgCvmgy/vEDL8sSifUXgImt32SxgavveuzgFZXa4CMLAnbqXDEmRzi4
80hoCEdHMyOwncFP1V/JpcDtqSf8p/0CT4jbJev9hqYoXKQLqhSNfO0TUnFatSVW
yytszZiQhyQROQaKxPhsRYgkJIMuoAoMAzBn6B35uGRdbIvAjKcNdm23mWZRYcef
/2boIWNuxd5GawT6ZR5JTgmBTJYZs4SwsS6jfxcJ3hA2bV04vEwiS4V0vdcNIXbI
05DvFPHmiOKwDcYlBeDk4XsBGMQXgkHMsyofsTDn7SdDt6asZxyZFbLbUZFPxF3Z
WH/3a8ypL8qGYToo3qTxp7/bgXvGhgyyt5iP11J87DZjYZcSsrE8xWxpHFZhiqIN
SyRlQXGGaTQ2YF0UP+1bhbpz5ZWUrohL0KFXJiXv2X8Dqbt36HAIAQKcq74ErjJU
luF3bnnrYStpm1wwqAhDAl4iUvT4GenCd7v14Xrt07hXXSgvBzw/K+TWiH/IxtxL
1ABi2T6l46LsSGNcG3p4K5DrgzAw7z6t6ca9b7/uJ7hVAQja47jSGgoWzcQvrHcg
yR2G7QKfu401+RS2BNiI13ykGFUJ/oWMSyIqCsyKL3dYto4CJeayzSlbUewWXKkt
HYjCXhoMcUEhWBIXTcwVCKJTOTrypdbs3SU2bP0FN+jn4+p+vfjfDIe2daOZhXTj
XpcqP0WbcVRx9hUJ9EqgqFIa1tFSxyyve3I2HMgyBywG2uKZsl8LxhbLhoJJatOS
YoTL5m6n1je6lwi8c1y5VfTckjzJ1JXVJdYmJiCV53TBatrWz2DEtxdSfFuWwU9m
RzVw5K6Qgu7AY0M+1meukm/WUuRvF9umLfyPWzBrbloLDHlZ6/jdV5mkVUFTnVXE
UJL3CKZjJUXH5S00x3v0+7PEgpS089MMCKi3Dln/ABYKVmlhUDgsRgqNQkWDIDmF
UT1IR70a5Y1qNX60P3yYsG+cXRCUtwmS25p2pi3ULUxpyAIUrdaAlgH6CBX6STUm
ISQM8VMyR8WvzIgxxv/7yhq4gjEm1z7Qe93G8c8ynXTBHx1nanrJ68tjy47l7OcU
Jap7SocZlkZdV93MmDqX/H8nULo7jew4iNWk8p/ex6gbeG/+SoYSrrD8RCUJ4T4d
ETiZ7XtQ86sonyVlE4yMRyQGL45rjUx6TKAwhUBQxi+RA3qL5NSj1IDC/RX6nUNu
zLExZFS5swsqh51q+jGtpz4dzNweyw/gQIeBlNm4x4/7k9RiHftkbBmNc0y9DEZp
OhqZPJ6fygszTbG7sfk7zVBtsJQH9leC5jCQt8XlvXb1vop22EB5Dm4AUS5laP3M
rcgRGsvfSjQy7JYjQNeOf2ua0ZVRm0/PvGK2Z0pllDaijwMKofMaqNpSRU93rNdO
M+V9t4HBW78uzH7q+yzVrbnt0JVCnjUcnRe6jE/aV68HWjp1KihsBhkrl5DqPn1N
eyabegs5L4xEe+SOOwDXsVl2Ss9vu3iEhheWObgRY1o6rU4HZRtNIVwhLRFGgvt0
rmzs2G82hPyizmMH2X/bUj415yy1q0zep8AmQbQDHneO18mWtFpVrlDcC3MoCEcf
+bLHiOVx7M9D/QhY8Gy34u1RSv7re+uu+2GN7KGA0mcEp/E72HnltEZeUzHNbIQy
lPk6sw8PCcif5fzFMxxq71P+RhCQqNCDgLzuhMNLVTfOSu9UlRzFvoraNqLZrqv/
P/Vy7JfZ4a1iWnNtNKicgcEGfNI1wkKbpD/yhHUgHe+QD3VRQ5MSHX7y1BWwVu33
bNniz9A3rtyUUqxhDl5zbZ/QOKboq4MwIvO2unVkzGZO5zCSXetcVX95Cj22sT3/
nc2RunRGQyrUDudbyXis1xTUgPYFOJabNe3OtGVqWjhHwwtCBWL8PmPfVzAf36dz
836Jd9jB3NWfKhivHyHFeHaaZIa8AY8eb5KIaaaUjteQeqZj0a/Zt/8ffI24yqM1
bSI6POn0XbcU00tz4dqFVdHpa3g62Vh1n2AR+nixvoxe7E7cf3k8MzSTEVTBa49j
VkiUMtFlV8cp1Ew+ED2/11Znwk4LzGMdW9yIa1X9eDahpeI7B04PMZxigys/0/ZW
x5K+SWzxpi9GJF4/+s9XLMOQcuep920jPmvzeLSLBTN5fcL/YOKzKGUqVT3SPirj
r30Oi+67KH0CROWFXBvENeRLGTRQMS6+S6ePPvT17JWJW2HzOcR59gV21ls/Nq61
QXlktkyDhyasLOlFfUUSG64+X0yq6/+v/imqDVHZvC808CcYJjfOEYALooZJ01kA
KX+6z+fSRHKTlo0iVv3Ty/iYJ+V6wU0PHMnTk75vi9t87k00EBIu91814R6On+AA
fL1S13I3JODN0XhJGEGioUKUH2LZIpBr1+z3/c/Y6olX1kW5PxlEWQJMmAzUmv1H
yGEcGmgXk/82p7Ow4fIWmJNPkuyX8XK4lP/LKOqfjwy29ded3M61Ny1iXGuDjY+8
uUBJm/taf3RRi1FIO9S/ueLnm6NsoW3LEud8pQhCmTOuiGxRyLr+C6P3qkMg2I6V
PNBdRAw0M3t9ZstvjwXOIeGfKOQY0VARO0Yg7UgqbLCVOkwaOjuUoah/TEjX3pGv
1BEUUfjfzM7eo2XvoCCnKkuxz6We+i1rXZ3NPlKmweus0aYJBIF5wIICKBZsyT+A
Pv+0d3VKsqBYhb5AHHBwUBMnXFUyQq3SSe6PQsL6paSRWntT3mHyxh/8UdZ0Tk+H
KZPpeJkRIUgO8Mf04I2+yJ5a4k4z9teFVSn1sreTtBlqguwzdBosym++SU0ogEtv
sSO8jUDAWxJ8scc4DGfWbyaMNBSQzkNWO7WMo9oHdgHnZrgPNj/smyMpSIOL81C4
JdsSQu566dJGtfpv8Ud0XgOu3Dz9s6U1AyU83g/C1rK/A/13dzQWqHJi0lrvWrIU
PqCutcJzGKeVVBdLD7LQGzhad9TOGZqOphQnrHfg4CWCoL6EXkTWQ3iPQYty892E
E4twyNMtsn0LfJkqTOw4Ydag8/h7J9XLTlF259Al+OIJdtOh+TS9wG/olCfePFAZ
q619YMXJffWZLWtXW78WLF78FL40W9B7Hk6djGaJC2OQMVmCXRlLLcrWrDBFTfq0
ZD6UQ/iGmENq8qAPDbaE6T6e+qOmuvWFNeSFwxo4PWykgmycGacVgtaN1QJnhRi1
2tUBzi37XNkx5jOLIEiO9r9qM3JGxYFSwXsG7SHgUGQ9l3rdWV3HHpvdeSqxOCbD
fhmOtQsm53uUjub14WRQoegKgItqeD/Fc1mX+j74qRaJXm4O3ATRfCBvJG8rt2lm
0uoek0EcjEXX3dJ2H9Z1UaVZWgSsOS7dlRd0wODhYf1soN342rWcd8D5cxWTKoF/
HQutJrXO1S0Sc+qLLPukaPUU4GAyRXaW+S6XM7i9WZw7usrdTySatYYQQNmSaELY
E5Ib7Iclr1XwRNavYPUtxike7ayu67KZbc76H+vwJ0KcpnzgLzs25U++geLK8yfo
yKE3H/ocPKL1gOk3/7+R3fbqInAEHDmK3kXWhXnNb1t06R0zLC0e9QSeaF1BnQh7
EOmP8GhNilHcq4MfBPydAjNvIrZBsnE2nercFV7AsZTc2kz4VcRaq59qeaT/0Xf/
z+yGVRtTIhLZgNy046+aTJEXAD2O9BSD6JDG/+VflMaxbyr2SlaooCu+N0HuhHIu
LBTEXrsBuRmXqelPeWpd7TMnmul9X7rZTqImrnJkUOyBboYL+gqTXTvzuZztZ4qc
BUxBJcddr690q7b2T/WgJVffPw1dpmhsZFDdfBRQPdXRrPxMnRgvPAv0liNe1Y0O
PEUOvMq057tttsccjJTxwzeh2s2vlciZNtijt3gHFLZYDJ+0dqM9M/Lx3TZYaIgB
V4ELPN37GavBS7AD+KpSTWg9usUqzTmMBw6o5jkI5tIqy8slB1lvbE0ZP46S6lRs
zZTos18+BmQMvoRRwshLAtUB7sdrUzrTgTfeJmhLvyO8D4LSFc7rZbXuvtK/PO0H
Z25aM2sgdaj874p5XVYh/tTbKtuxFPFx97UsW3A8yNg8QATV2pgI2hBZbIDTOlMY
hlZ5SIP15AXE1kYSnfufD88YHj/G2js+BSX5ZjB2wbRxQyoCUO956opvyU5GYXJp
3aRe2YK4F8mCmPebsYSoWH9GHLokng9ipRYyZnHl8XGXjyguhgv5RtWWLPQMFzaf
nd+0UOO85eUdQXAwbf1c5gY/pmnFsr6C2Cgmd5ADsdOkjuXdeWQnn1u3EdGAh/FL
aB00Iwfj6yx4k5zpQY0d7q+xJO4jTQNhClytP8J7F4yq8wYqgHzGJ/bQNYTHlQH1
cPMFoZTfnRCA0JWSwv31lHdw5CMCO1LbOp1ioovkKK+L1bAwRDlrczO76YpQCXW/
tF5XlI8GRk7ErGmCSW0ST+RbYish2Y7sv6s4ajOAEYUN4Co+jYCYwL0+hf9lIw50
og7gmrG5TtvUifXsQLOr+zYxr0Pi8RJ6UFST65+IzBt3aAVjgOYFM2JgtZf+OHJI
Lm5ch9xTFAv761d8iM6SyZOvxEI94y4NQ+T7VySQYMZnmKKKKBwzBDKeiw9lvoOp
1PSQe7F35C5sOKu2+/Up7hqUxZpMCZVWqMMGFkmoEY2MsyfoVQwW8rLQDC0YDIyz
v2olWnVD/Wx18vlP3Phhfzo6eoxFaZ2s/qofBUmk+uLyzFSFlrx+3+jsSqTFkpTX
o1S8cI/Ssg7BGxVJQZ2z2fU+2NxfOlDPqz25k3NMFapEaVFWr4YHckHSJRjNr0UI
8xs9cC4VqlezievJMIcDXQdiA73nnNsi20yQG6zVxQf/oBwLkJ8v18WFdV5tXONK
Poaw2ik8p2FpJXX2uPO+NW/YkuqhnC7XAv69v5c/gSHnEaBg4yeHkp6U14tvBR7x
dxyiYxGlCQzKjTtiOXp5gzF3Q8U2cpriRaRBMRWPti03LE7hWa1aWivZvGTUEn70
CRy3rLehj6wEMB6qHF+7fy/WOvVD5F0SUgJ7/MEZCl5iCairphJueDMuIIT04rHy
a2nRaSPAT/onZEfSjs5BGHdHJP8MDsYBxmBsapnWMwx8ebOH57kb9bjCOfxd44rm
cixL/w3dOcSU60JvEei/tfpPzXXezR14ZWTFxCf/x0OyOBR1Wg77tIUFewkWAzQc
auKJZ/QOvjSC3UijFivs3a5K5Uyv4/h8QU9sH90tt6vd4ZTdQSFPM6UHDU9+IFiK
Bv6glq3zgt+Jap3+e0YB17pfTHp+LJEGzYrVqURLbn1mHYYFG3rWZB7YL297SFcm
lZmex1W9W78t1HOuCepywHkXDqj1ZXWyy1lb4v99jd3jPMnT3hPn0sxGv7f3tJAb
PW/kbciqFjscJt481wcyg7LPMHIOuGEjYDaV3QCjBsEd2EHnQoGzhdgq3DvXqGfy
pSE4XYWBceou9/UEemLsz0ovtQdXwmw+VlHrwfp6gCyp4RaxqyL+LjDf1Tc1Ky+W
gJrBAxRciqA1wSK5cAuub8sSIbVnxa2vFHL6DRf9WbHMO3XOmzNJQWa2eV4vov+R
/iaUC7+RqkWzpgxUIixyWzfOEbpV1+gr1nAensSpISd5j9wPkXSX/VaqiBNJjU+D
gKNChmYxKHp4X/RkyH+yXyM1MRSz3bWuRaZN6mZha1orpSOjqaaNjH3a26u8GY/J
xVdUoNJz1ik/KdM1dSyjkjoMQIo+fP4/tszJaJJNTtIzDe4zcM5ixqtgosMvA6p+
CxnBl72H1BDaT4sPy/b0I8NyKF3zyoG9WLS5AmgH+F1HirHygV6v6q4g+fJQwIy+
Tdbq1OJHBiYk2PWwX+B6jTs9vLIK2sW5mB9JV9ab8px1TlJgc6mN8vCVTQpYRgk6
izMhZAf1ah86+AnqggZ2HwQAF2fgHG9/tKG5saFdXeMNVz2aKYcXKEEu3Ttmx036
m/er4NZphxNTwlI0O/WVD8A+MjQppR45sOgLrwsaHEqNDO4Vwp52ji83j9nJF4Km
MYu140REV2BETCMptq391hHNDziMufArnC8wyOE0DrNduci84PGwhiorkFEiajiE
bRZaVGwbPwvNpN80yaKF1WUrKAZl0YZcFseJrhvZ4lMfErzvY9/MGG2vKFvdjZxS
EdkK+NyaVU5XgkVxP9PR25j8It+KhzVE8x933C+oW3Zg8oegVY2aNo4oZg8fYTnb
ffaynKeV2acfVBGu9I0uDQ5G+QsU6kM52inpfULbsh0WHwCMjhuNpNwF+8Ggp39r
I4XGKNY8LjEN3KcP9/yB44DUXd+dy/1Np+466jbP1Xvq3/a55hkXFkSzPWarHPeZ
tPiHdIJlCXkkoA4jwERsClnKXtUpRKKQZ1FzXYhHtvzEGfm6zbi4x4OdJHZn+1T9
PTDtm9ZbUDu6GrsMRDC+C2Y6/dKTRsvv/8EfddFkZhXxabCLPj4edxOShH0kEXL0
q4DL+Xyv2NqB52DDfCcGH/xlcqo6LT3EnXVq2EAFOTVMic34RTY3fCZqNlSNDznF
E3oE1pei9TkW2cCgSYk8lWUsqakRnGVZzyLlrqwVu1ot1Nn9E618WGQTkRv6MUsQ
dyXhJ9OzxHSRoBjRzVKOJ4A2/8PTdWhasaFnYcTKBuHXoSkIEwwu8NM9Vd70iaMn
kEz5b9outTpM2nYJsHMcT3OVM1DF+ALBtk5r0nCVob8xJpOs2pFzFG6Cd6S4EmtH
lnJSk1j/ZJYGvvzI8v5CPIX5PFa/qChKWK5B57xX9Oak52jL1hmsh0NdlJJEhKIZ
69fiITNGqZBBzgzezLYy8WVMrfmUm4c8YhaD6R0IzmZcmB4RQyfcdXd36INZ9GTR
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 55056 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aVlarhe+WUv8WRJlOJJnkAG53ou2yrz0BcDB15W/Sj+q
0SA+EygBYZmRAeXS5ded3MNiPSvSdZW9ELoDC8vWMWb0yKCQx8x/gXiWu9XhWO8b
VXQz3mfh2UblQjz6JpUa9I4efgvRQKrLVORhbi6rd+qoJ29gNdI+fEyUToRet18y
ouPHi+bAzQ6axjf9KyceSwhmNtb3z3DQaBu5QTQJd9QL9gUpbfH1Nq9hQgWGYcDj
WRCPLWs9itMPjc4iVumq9VMllP76HcNU8nB0qnYsowBx3ajWvT5awgUYbByH//h9
vnxqdfQ7JVv/tuF4MVi5+Ki80WaSIpg8akb5mNNPCYJx4XoHJXpLS5kWRRM+scsO
tPk2eEYhrsfMllyhRpA93xsOWdTkLhIDNr0Gl+K1hCLW+oDm5BeEFenk5nfcPnVQ
L4d24LGuekIWcdEZ48jT7EaLfPLDCsqSxzDHzuABOjrMSGi92DnA+Ridso8Xo7pw
0luvuvvG8gDYoCpeYSfcy0eucolSF82Y+Kk0pNrb5XV4Rs6LQ7IWTGasct07fej4
kZnw+IUwWp/HOT8uQro4mdoAYWWnCodBoTTA3dG6Gn/9/PyMH2sxiQ9B6izrqih5
DkzI8c3HNuYbaPMxjpRcLhFagfEt9lwnXoOwv/1tSbjHt1QdcCexxlEAWoqOWoVk
WSer1/7v6vQ8uiP4e+rFg4r3z2AfPdFk/pLMrAqQ8xvKoXzljiI4/PTOxpTKNCSF
0FC1ZCsy4Ww8XT0tn1QlDdkHW2YEmDgMna7htfWFyqHyRQt+WrF9/7TKxkgcfDNd
gdUFjztdbPMbPAQoA7EVhqpNT/dMMKy5RINQjTNO3iXORwL8hVsXk7CUpAZ+KJTQ
6iLNvdXfBdla6VF2jh/Q3lCHPWyX1+cTbbnswRrkw2pBnIJGtAZzNFFYcWN0ZLzF
ORuKFgFPOnwQRc67xTnSlSlAFNDGRIir08p2stCjLH7OYchlWblqe3laVm7cx18E
oURVWJM5H2Yjtz3v9NFQdQeDSaVyVfI1RdXcotd4jLyHqcT0HCe1EXDzSLPVs0L1
WN2bGk6cK5AhXeMNG01kxplCv2zpmJ9Tkl0y0DPrBIy03t1gbPszBA9q8fcrpZM5
tO8c8LEhilYGTuBXNmrtLkbFoNdB8tibVU7BUeMhMFapcp/YzyoYZpQjkQchSaxu
eZrqmBRGXcfrVyBcvm84+0hTQCCAbTcaCApHn/5Gj31DeGyVoSNeNjsUqHIwVfNS
I9x0Ean5RmzdHPTNo8uJ/SEPztL1a51udtRuBUGJhac4plaQ4PTNOob8sM+6haOY
1hsHHjMsWutJysBZ9dAUjDn2gNT6EGKwNSIwe43gZPkSMcl2yd730GH2ZIwkLLOs
nqAAhU4aJZQIu4VSuklzz+RYfOO0yLGolNihoxEsKyyrY+wiTxu9C19Ngb5bOTF3
RYBSKVprRZvJYX3iobbx4mfj/PFMSzgR0ryMnTDz2LYosYD3YMdRoUnIgncZ9e3e
LajArF3CJftRPxzgLfcaAAV5P3InhBBoHGuu8vV1binKLObUJJR2ulqWS5g4BmKH
aq6fAK3B69DcRdcjiPcm11GI5QMRTYobK6s+tKXA2f0WW2HsaRfkUCkPY96+7sd4
jMP7QQN+Wl1IUFxXKd5ll6VxgmFFCMD4h8RDRCI3/qoCBKgR1e6hg2r3S4aN7omD
kpSpahouvtVJIwA2toltpxr0EP/I7Rypklx3MAuv1rGCfQCIz7AogASUFeLodsz8
YzvMxvvc5IzynzencrlJgCAK8MHLHgrxy3iyE4hWjSsO9r4rKtQhb/Dz9GNQe1nz
XAVAuS6ND1wWcmU7TiNnvjusIExH6Cu29URjullROPUDSVgqV+hc+sOZag4eJa7Y
Z8csccLwJSre/M/FXnv+cJ1y6p1LDask+yewfTM61hzq1o8Bhv53JhZclPgXalQz
1fuXzTwQbC+6HkmnyLIlcxwcFkehjbPI/jeBSFQnxet+4S2R5T133HLLquRjJ8GP
B5dmUSmU5JmDtLXJFBBFCnOuqMPk0T5/QR6vCRtbAPTnDE8RR+JPV9JV1mFgIeoH
ZFR3h0eLbvQx04WarSAoP5OohFj/LWufOJLFTQxLG//tgvqXZ+ivsnM7TQKlBy0I
EutCnA4++XNAhGIild6aX5ksy+MrG/9hKDJlA9YKpVd/Od/7/Uj6rdfDcgwZ1k6K
gQRcCaBr1RLSCQ0EnzCEyfG1SkdSj4vkh+vsk09fLyKqCM9fYFJ0sUVY4Uo94w0s
KV2eOuLCPL+MBuYznL8xEQ51ai6+U/T87G1/8d25J756gTXSYsE+1YxFFsBDBTZQ
+k5BqP92oqaKiZo8YIw/7lkY5LWTU8HakwNWESoCzrsRqb3Ltf+bH6RZrhGBG0T9
728VpacY45aC5TwnJ4fFsR0ivfA6hUYAgy4LZAxUegMhYJyHp8oYr/mrRiKUzI00
FafM7UiZdBp7KvPaKz6kECs9RvoO0ojLDSrxM+F6gH/c1TtK3NB0tQoKhYCpBYM8
3Upwr94NsM8MYEmk3n/FaXtVQzqJlFebCxGfRvol82TyTDdjk011udBI3jT5LQak
UhhoVyDbNrp4FSsPZpQWqiEidUbwhk9ZwlAOL16HL6YX3deceIFbo5p2P1rDug1m
JHZe4KJ1xA1MKUd9Dj/+99HD66O/1cCqP6cBr/xeVh7dPRMX/9kE+izXWJGcMRfA
unTYta67f/0qEDGWw8xZZyL42HLvUmXV7WlILj4ys/PicBqnR4xVgShSD/Bwnnvq
0TF/tEYmc2QAf2U+cA5yD6BWKjUHc8NpSii0Cw+lmk+K7TqmRmx4JkeK7C/V0ify
Dh27VDbQ8hZ0qpUNHBpDpBZr7IRzqagvBLhHqVphS0FV9h3ucTbHE0nNEVZwKYNG
wXrtIq7P2beLdD7aqP1ESssgLjKlzaDVnE1wwyoEuvEXk5KHFQ4SF63R1D6dm3yU
NIy9alpAYmDgY+mwJECIs66ti0SfHTV4w2Tjb1GMVRsQbZliRQcPpyvrNCSyTsPE
xEIEyGFY2Z6HQahLrtCVZO4tGIs3W6ZjNc/SY8oPKRgAXZ/vk29lzJTC1ihOh9zu
CE3RmWBeZDiwjq3diyzgu8AGXyfyPWPJUs/l+3NI7l1nYgHk5bTde8Xe/bYQbBIT
YfCbHILmw6b83E/rESqk9KVTzTXTPrcRpitJWgXtXA9Lq3BExGXjxoTrXQv50ApZ
zuHjVG+uiQZG9XDzTC5TcAxQeYuDGsvLtKzEe44uPAr3+RVjvoDhD5iVqDzw5VDA
Spa8z+cLn+S/TISAHEvGfdKAPckYkI9otGt2LZCJ7JUlZnVlAVog314rb2BxgMxz
MljOFX8PwBxgEXu79HJbqjUYQkagZME56gknPNjljto3ZmVGq1x/Nlg52O3wjzvA
RTjlZK8lKF72E5ghOFcO8B7fksONoacuMmgHlWfusqCuYCA4HRiZ8Cwnalj3vjGY
8/8Vk8NbhqKg4ABW91JDdVR9LwrI2BxeL+uLUrUWTgvVUJO8VHxBX6+pVhO46Os4
hHJ7HcDDfqmPC0hlGUXjnNWFQXl9eQjUR3b8MZE6Ha1dv389nFGUXhE6xoT1Tqqi
yNCNnDs7eMUK/Dq9VgxCWfr9gTM3f+eLLJeYgXEdQTYkneD9ofTn1Q3w/92bIfD4
XrEj7d5zA2bKiDGhbpTMlmJ780NEhAFPllNsD7PjTZqQcfCZxe7rySEgM9ItemLw
ulFH70Ic/SgqirY46cKnXM6oc1DSqs4Nlj5vSjvRmyirBjrgxfL7y2BYddzJTZK7
1lhvxVXXiCHfOYK1+mZW5YkQgzAxEJvWd/SPE7V6QKQkU5hebOGbqNg8Td/XUjbs
thWDbSU0/eQ3fp0PVPluEOaiQ4BmpnTR26VpTi7Py97PNBbxE+N81viQCUlKHyl8
4quE4r+L8QlAwpRWIVlrsi21CdcZdRJ1Ti271UtDynEJPzVibwWhfFwAXw0cvqo8
o/nMYmVQeAuTs8n+mYmpFYTIChFLTlbZ8eTWqF99tLZuEubnqZlEdlXto/jnOE6j
BlAFJ1ldSpBed20cWxPungKgWb1kDX8IxcTLUVQBBvm+YYBjkPLSbBGwB6rhUaA5
yPbXSFVIPlHwMTApxORs9X6Bw/M2xAPnZm40c4P7qDSiozpzplYCqFOkxdQkjcCw
cPmAVPNewuONgxa7HXVKzcZelJ9BjnjIfkENmmcRoxuTDK/+HOZintpES4eF94ce
q6Qd4GSC8ptxR4/WxtBAZeAdUzUtgUARSl2wSjggqnfZFLjYnqyzuqLgnapV3yEV
sVDOctLxpTRFJ4SifNYaUMzFDoRy7ySHLBPXDaXcH7oWB9TDjFT8mJ4S80CORa36
IWYXx4Q0d9xH31EDYPHRNIszjffmX2r5CrCAaU0Qnr5V2awHyfF6NAcXlmabQqmD
ElIabvezOJ3Ver1xEkT+8mgHL1VSDjmS8S7XUmlCZ1ZRyFxQHx7c4SvFq3n6ek+l
RP4rk5UlmfIKC3XqSclq/LrPleSV2TWdkx7pT6aAJcZK6g5vCQMphnuoCcNFh6cR
227YQMMMZmRncz8Qq62JviHFR6iUoQq/RwPqH10zboApNbLPweugDmGbGY3MVw0C
bEckdp/Hn4HlUpWQ84vfMmAuI+JFP14Pu87yTkypABWWWd+5kirNFgkDS6z/LsjY
VSFQ4v/hqOxCQUhIl3AIHR1XjOqpdl5HtckMZMOt9OooMILDhQ9SqGcVPFcWDyb1
xTwu62zNmDlrUWlDZ5oQm1xUZ7t4sePXyC2voao0cDj72FGK9goQAxNZ45Z0VG3h
EThDtd1zsmbWzW9H6eROtsN6v7kH3Ql7432BxNiZR/OUv2A6tRyxOjyZJUHr1A48
f8PS9i5tk2XwhAhTDEZcew+o0mQu2gd279UDFNmjU8gi70vJ21Liz8J6g536P6e0
w/4SlpBJmS+nHWEDAXzVkQ0JKpCKNp6zsxbhe+xvzqMWbJejIhQa3alkUTEP/REA
SNPyV8JhddnFpzfBjU/IDt7iFIHQOfaiWAiyBJz+gOlvZWWlMEJLlCXVPBvuEj6g
LVntf1MO1uiiyxSHF6+iZ84OSCfWp6HPLp6vlCyn5zOFA8DIYXf9P+6TMOIya9jN
zCTtIYJwBnWeWJeDqV3KYz6+8oVNRH6YiXa1av7pYT7zkIchcmkNBUu/ny9GzLmV
1uEshgTauwemjctaEJ6uHdu30SbKJLOEm7b/pFjNDvNiwVag7ogRI29nn5nYYW72
uRqsdWvB2as5gZWCHHHIZEUagKZkhnzP3jSh8DAVsJgyMLhG+gy72IKQq/MTysMM
oDOZVKRVLWLdbq957dKxAnxgfLO4Up9HW+dEE2bNnX0zOllx+ixmvTBuUCYHdTHh
+V0rm5VNpc7mb6cSIfOlEnPNKEkNOhC0sfcC4Hb2SgO4ujTfLfX+qOZsNMhN+QQd
ioLcn/KKSPIvxrxZ48b7PXEuBtJDLDA/bsrIw4CnsQB8Ct+x2FN9PO94nm8P9ecT
dWgLtiJAUlM6eHT1uKHfQSGXysrozPM7sGseCtcfelBSEcJQTbi5DnkLX0TSQ+Us
y6mdDMmY63J+FdKRkYUkyCuxk2doBXQHAD+qpQeh2IEr5DSh8PDAHoc3O8Tg6mWI
YaQFEuUMCaTrc9JQBkAwcVOR0GJe5y0VspX4QgIOlTLcHeZjLhJGFLClAMk8+4vR
07DWhK3psLCaWDNw7BW7q7tCUBd5RsXsRp1PfJOuhYrdsOPVJqPBqiFryEqE0kNu
f24/0xeM7LtziZe6Zdj/L2Oohx3G3KoWgr2N3RYys/UAuR8ca8JeJBgaWTfyx6Dy
2/I0ZwywPtEjVtowH4aADpcQ64A9E6BxOTFMChbXfjfoQhqjXasnzv+akWXuk0/c
HjCZqVdZLEPB/oBCVSSkN5VpECb54ji4RHC/DSTXHzIS3AZxjxMHcujwi3jWFoIo
OjkgSMxijLkaAlBNfNWCmsyZUYIhT3/xP4Gzkv0vpjuk+maAbLzFvoQ1jwPtg9FH
f+YjnfDWO/JjugDZtQamGUs/SKvNYDrw9Ja8LuELZhYVotWrD1GHmkIDmR59+7X8
wuWt0rX5WZ98ERHJzGmznvPHtgFaSGt8QWMceRV5V07CfrZwXa21jXAH6WoED8WA
DWldebwB/H3skxS5vPJSe8D6pspla9J71p+qaOOhNFa569ANO/GK9ztFjk5Vphai
gVqifKmsQHSxVlcoO1CZpSd/0TwEJmaPenSAgIFeXS/bs+v1e0NFHi0C8gttUj8L
gAicYC+CYZdPGARyf0uiHUEOA8NDOfYn6AvaD2JDrnjHCgn/RSjJXdzuTukcid8R
n3HJgebhM92IJeuG1+q5qaMTo/jxNYSt9dCLxdX1z5Y44vtUsyoPpbQY/heTnR22
1VaUTmm0jQrf/qNT77IN4pCdwCgzee1Gb+2dhqPQC66JdueX/H0g9yAjOMn2JBit
/BXoCJgM7U+I2SoSIEjlVfm3AKVbkYv7n3Kl6Ctc5QL5AMCGqpfVvLamhk/UGBZF
RFrKs/H+FYOBQwNCyQQI0UutwC0YBxWFP0Voe/AhBYorvuPzryKZUYNsHPLHU7Bn
QSH569FmtgIKwB1eqBnRiKKiSboqkcG+rQ7D/t1agGRnDWc68K203B4RVej0nht+
cMvefe4yez46X6sEcH8bU/UGpYt8OubVGqnYY3NFQgDQd6ZJqPvx/eOsMjkVkr56
hoZsZLUcyW+TmHYFRtXrSgDRFUeckK3f4wNeHK+/J/+sq8fS7LcszKGveFvxXwXp
bPEembmg0/JjAfGfcA2jusJeT/Ps1Mu4C0oTysrCoVzAz50ECoCki2O2yX8hGExc
CXzKJqGusGWcAav+/luVeEXLeiQt1q1XR6Fja1kR0FOqvfimDMmellSYtFeGp2Eb
Zfo85MxuD6ipMwyUyzy7LZLsZnpiTDj7KHgR54l9XfUj4IpoplbfoIFmjbHoS11C
Kh8nZRyz3vipGR4kMWpB97u6XyYFtPK3ozxZxKq6leuV5zTE9DCPB6vV1vThWkp2
CWzG3lNEFZxO+rs3nx+SqHCbOgrb+YGfoTOOpECVDmYODZA29lMYfD+/ZdapPVI3
YpfwVUJUYywB0rdM0MHfiCb3NN5JmlGskHO9bGO3TOwfAG8JpRYjbzfMvTSNIzGU
hln2z53PcsZTbuyQu5LMoXbu8qDt1I3jZ53m2k/+pnS/IRYVBnzWgAEPg8i6Bskv
CJ0ZiaA202yKMj3fl/8RYYcW0FIhZ0vi3VGrq1Ml941MS02IcQ0h5YKayDtWaptC
upiaa8wydDic9r0E1CcawVEieRPSNDwMfw2GwKZFi/BIpyzeZzAXrHt4fcrnhiWF
4VH4XgxtOYnRS3gV6pRt01L9AFl233Tibm+WTzHf6G3N6CrXqKXQUBUgmdb404x3
P2N6nULKFgH8x+zvUnPjs6BADo0YbtiPNfNsMmC36zFEqiNM2K5rI3Te9TBD5Wxz
ogOPkmymDyjxIBxIckAoWpHElLRlkbVCj96HBWLSXmuoXomETfwLfjgV2JK0sgGz
5qVACrKoptxfu/c4N0mH7yCTZ7mloJrMUFI+9V3QKImmf/GlmSOAIXW9K9gueupW
x7DGNOGGxYD/c0bHtNrfShnQYJIYJ+AGMlbuJiTMMAVtc0mvi8BBXR9N6PbUE/G+
9YcnNhPm1Wamlc8eoMN1AOaIGsAEidTiYEY34M2Z3FSEhevFDYegCvvwLa5Nfncz
aN3hg3MOFYRk8ElD/m/ahkRmP8za65cd+XfDvQ9nI6RQQiZe7V/c1F5llH6meyZy
Jbc1vqGLBIXpt0HICCRRhShLWaYZqaQ+OR4ZVR1Kx0sAGP2FUCkHTR2HQ2IUF+QP
SRNBTZtGDW5tXWntwNAWf4miVhHg1wWMWD0Wv0VS3MsBC/eWydobCcAKoqt6b6sh
YlTngNLlf/ifUtaw04/j7/VMuD0jx3ieVlHm1l+O4cjPNmxehfSst8+h/qLly4W1
oI258cliidywlWj73yBDQt1EYU3kSUSStGiDE02AwJY3KORWRFMYFxNlMOTDD41e
+m0lVOe20KenSOuag/6IuEuOfnrXvfgtH7JsPyNKPlSkqiE5B3S2vAMuW8+GHKgS
vey7vT7ZwTAyKaP/k9kMfTRog/zPqAEqys7jw+Dx5yBgWYyRstStmtsVitVxRF7g
DIeN30GEVFQqmqkQI/PyBVZR6iqZ2BF/SZOWOs2nyMeve8+tFiPgqNBcvl7Tm8qh
aoEWSvOvP40hjCibphtB0+Ln5YkVTxIbXwXescaVp1iOiV9Xwxra2MOgLwvDdyPV
+C9m1FJKny++VnPPk2Bl+Q1PBZba2dKdbeCbGi9xO1H5Ucw8OKMedH0HVEB7/lJl
ehqZ6vvVIx4Dm8sZfGXD8xq/GHYlNLBYBOQiDb24v/1waQVncveF+qDMAOZl/yIM
nouljXs9d71nOB49M9jPlDjZ263LrwFhaKb8/00qewXzNRtzHt5g4ZkFCzHmCgBN
v0MUqhbmkXNOq4Ebw+ooYdrGvyO2AZsTJ+rlGQGcE25aIcR+TcaxbTmKvzNEJvhJ
A7grGBk7Bb0waLRFDesNJ3yjk1Rr0ZM0s956682WGMZSqlZFOKtoRiOw8YaeZsqZ
2ak3uZ0xz1k3VNB76rtuOrHO4+VGVt3/erMy08H9jJe52N9TErkyP1mukefOdm2v
WisR3CeRl7iLN7wbuNKHIf/Zq8HTOWIpBSgDQp75r0/jMf9HawmL+obfpq64tJT7
3LKCWCldIldEVQYMQXiqzfhe0SR65UDr0+dcm/GybZBxkJeKkHc4yexmaUUFBHJJ
h0KYrsG8iah4ANrEDCGnY4cQcuGCXuUcJzpv7UXW/pU4ZnVvVgVocTeFXmQSq6cU
YrjODT+KrSeRs5cbsd7JOzVGEp2ki7i3U2a5iWFD2U775WfVSlKp12yBENhoGvxa
yMWqSHjil1QEl5CA9z9AwFX23xdaL9qeTi2xxWbFcjrqZa0js63wS3wHbQtnPcqu
ZUpAFwg3CtnX3x33LneIF5YYrwTpTgoilNAxWfCVtSKYBiS7bAguWZPH9t8N+tW2
bn5Y+LbcXPA1ALX+vrQ5OX0VAJWSIjdiswMIvcCaBNzFnwWjKF4lK3vfl2nSzqmY
ebQr1cnhQzIJqc//2mexQ8qYacRoKsHaPpQiZuhI3su+ql2rk9paYjEzimZWvp6G
WFetvNNlt1yXCYRWzuc9nHSlibjR9M9Va3+p+waauU9EcuFmU19Ww5R1ssiOMYSI
Q819m9txUDjWI+S3cy2b2HQt2nEJ6UALesb5U0SYF2VXJqVu6QPNA9X2sGFrzUP4
gxTahoWoV4sds+IG7jAD1G0G2GPKsY7hDcLVpoXP5vNxJa1Vlbl4HpPbablKgNIz
Z4yoDhnYNg2ltTV+nwXhRjT6xJIENf7vrkubZ0Zob9JCc/h1cedpzxjkui5WoU8u
HiFv2a39hjpcHurgd+eXWe7+xVRe74onLaH/kv8ZBFCjPCME0zKeOIWvTksYXFLn
vjl3QupUg/BNHxalfQ0tv5A4l4nq1BHpTFvyvr2UHeiLWkbgk6uZF44E+PFChY7R
15HXB8aBHQJwxmEvGgwCPUODMLd9Gic/O0bp2irkV8fl5l0/ykuFzopCCw62SDS8
fCKgikSOp3yD96JuqCfDfPaFYI28NPFhvsoet55JXyFKoN0vtxuLCpsaklYd0CdL
FkqWmZpEq37HxOXtPQPh3iaBSPQ+VR/eFsFddVxdTdh++uUb3iCAooewGbx4OoYL
ftIxlgkmNmav8BMyqMumDDPZRNYZq9z+Kj+WIMZVHgUfbz4jrpmREqlWrQjDsoei
ZBjwCneMONb0bCwVgr01gOPzl7QcpUrAIy22dG4DFY8MiBkCP6YKYuekrZzcgDaO
utUtdyeZm7ZogrofL15F39hKdSqGAlCR6xk35Xy6mcfP/N9heU3/p8OTH+VOxOp0
ys3sOYw/SLqLjIsZF2e+HUiRCNGERIXK9cLhusLIh3E6mu+7QxtPBeHhpQln56u+
cFpx87nDk8TvbR0BuR2TG7CFAV1GYfrHslNHMmJs0crFVo+jLRqbsSJROTXDARop
0uv9qiZYSfWP4OiQEOTg7RBR/cS2Kvaxb/+22iUZEQRjc7cwjUcKX0jCw7Ck6wRx
DJxZWulXV14KkYoNNJUYZHDVvEFw+by2/dxfkoFrXEdw5X0EowpDvwz76pALEh9v
Fn2JH7AB54AUXo9vOquEVOkTAp8FEZGAE3N7PjSIXl9cMu9gPCjvHjhPOdvEeF4c
MngpdCjhhkTCxdebl2/1to0ukALYm4/SA9rHA6AZ/vATJp92uhWpDqoJD1AFFtIe
Vnftst58Xk3Br/V8ozzYSg6nCSXg0/D97DAAzn/FD4bD2QPe4OWss+2cMlM2oCut
5TP1wWaL3aXID/MAhecSLBxxaYEdktLu3mJ+PQ4vyHwBbo4OW/W/npg9ZFKyRhre
AKd/idYKlx12EZK4Bk3jqXMJfOEz5yZ2G66CffONV4yaNUukyzHcwwImtPGKVQCh
BSZZPZRdZFKzg10UlZealXDvKPLUSBfvealrS3OLYe4GI47nRjhzaMFL6p911rMj
YZnpei7x8nT4QJZRs+MFSyPLbBZEWe8zpqSDIyAmFNh2abPJTEru6GOPRSXtC/ZR
5cDOfmhFuavGklXJiJzWQKY7hliRVoL0GN00NI21fMOLOoA9L8ZbfYjmNXQqRA2M
t3GZ7xobCqXPMxi8oHE2RnbgmIbLYrw2cdHXouw0SW/CnPAtAb54hI8g310+rK4L
waIoTocujB78d1PPiJDwWXrJm61mzPRLP5pf5i9WpjblwFkU+CUxR+jI6BsLAr0X
jGhb50lWaSNxnFnUBlwILH7bGBC8h/XkFwkExr+HH9sSBOoFfgmVAfG9v+9IYMFx
06EZ5dfknVprbAbqrlLDTo+601XxKzS+uIv+9MRXlJ7ry3mlVMegcVGO82b/dyXZ
2s0Qd98PnEpJrcTsVJOtIAzqPEFw7m0zDT3L0Rqk9obK5ez0Pv/XhzAr4bwyI0UZ
oSrO0VkyheQ82J3IMSQL5HsKWWBWF7vkDJI1bIVBXNrwAdiVXAGTrFrIeQCqwbUF
NaCOvmi7gglh/Pw18jjouF5HvnQD9psNXOUOWTX1CCZnqqZeB4ofDMQ3jRR2zw+B
Cs7qv/GeZJwErfyboxdLRoWSsIZKL4HoypGrK897NR854aasD3jGfArzYHPZVX+S
z/e+qlpTPEmeBFdBKyZalkEGH+Rqg+4MqUIedaNONvnkbUGXIQNvhJNdd48vnner
zqUeGJeIE9GZXGUgPhI/zPhv0dJgKi3kh/WZgwRQ617zkfgtmrCB5xmhu5x/KQdq
UPkpWO3QcEiT0sRJc09AgdTxMmx4+jvUZglB5RfRjhIX5ZJxQxbL+BrZbeZhLQod
DqWevK+4ZHoqmT/fmIQ+QdH3KwhmB/OghPeDgLq5aHKS3M1UX3xNbja7UbGyI12O
ptuFzWBYsi5TrC7S0a1jDU2I//wStok3UoT/3TVV2bkvBh1qMvzuJ65DXm2M5OzH
pc3s9yIAbSzC4BfUbR/7wYrhvmkCZ94m0fUp8oBrePsF8aly/EBqaUoaP+u8829Y
V5j0gXNfxd20Kln8LyY29Gk7TeeYVErIIxCZiiATnHEjPLsLeXyCNrSZPrbfjJAE
M2bNdlzRUpW5AOZAu2/zfRFrMLDI4CHVLVeeqYLDM7zYBxEACMgjSFaaNGQVnG07
pBWsCfp1wqgFbXi6hoA4q89gg4rUTErTGTwvYqOqOUU0u7moYE4o8itqKl09Xk6t
Sw+vscnssun1YQVzIMjTY6av4H5FVtKdphKcj/LVa9s+48cKMNZ8xhi844SVaXc9
cxRbHPZR9VjYz/BJYL/U9ECtk3V1TL1ino5DNsSizoBVgfz6hWnfH/zYIXFGnPjs
W7Z4vZ9LRNctbHxpn2tq+N6leuIv38GE1ApCZ6NFkaoZ44ZmzuF/ADUp8dVpRyha
SsSSBpGveHl71RkF2Y+HqZw1IGfmhbRI8jtSBb6nCXOWsyxJsOQxsCBmt5wQGVEx
RsrHL5OE2qM1VOIBXArU/u0JDFGn/jqiejmZzkR58brEQ2bBagSqc7S0xY/meJoY
AUTKZGjgbvi4qZWON+P47nPNHnV6xCAPl/6NapbxET/n7ws8LrRhbOXiuOdu8ru5
XEez+rYZeavU86AMjGYnd3a44Z5miPoXJuM75gGINF7e3MtxJ3Rcc9hLrBVXS4rw
k11dASWTPcTO4ylQlA6805oUgEe097bOqIQGBmtb6xJzCEX5+WiERNlY5JDQ6kZ8
c4gLTjy6b6j6nQKsFEOYxN+m1NbxadKOQf5h+3B0m8WtBuGgQEjpK5UVlIQi/f68
StOKIa6WMlFWAW7Ma4U+Dpp7/ncYEdZ2GpizRdpvm+n8vdOsHEUevzulB0Fh2dUn
phk6N/NdnxnLIoLqgnDnGxPov1XWBHwXkR9C6Fr+6T92n9hwJJhdvEYXtaj+Id6Z
SIUjpcS8jnb/mLWYhsTkkITWWdyAYn7CQV7oGY5CTtblymIlugyGZnWzYe13AcHa
JAoSb+zy7zG/zfbpev60PtvtcCz8CnzCUhsPK8uq4mOS+5hwWYeCWqhPYYcUga/a
nEIsDeA/GJeBkPltHhGmLsjH/Xn121Ryoh4uxg2jbSJO3+XdC70/lrs2R8CjHwLn
S1KMRRUokqiGVz8b6M9cCX1NHxlUpLrU8bCqH+zxA744fG93SpPdQWUtvgDW1ZXB
dWeXpAEJ7x2p5mQEyRY6pj6oM9/Np3IkkcMzQBtTzGs+78MqGFJNlAfKrOXhyqWC
bwaenxgsIu4LRT9PVpeQ9A3H5psnM40Y8tWJLbnfDGczsVYFGrp3kS8K1dlFx6Ev
U5h3RtaccUtu21JahU8cU/Ad6Rs3MmFUUV1ZVdBVg+ZPup8NF5L7a6azxezRKACU
AJZD56TH75l1EatNnJUF9Fj9PLhLxjrGvv6Ypa9IvqV06XuUkPpkcD2xV3EMKjI2
9okmm4Z98NYJpbPnvyIDjTkQt5vOanEK5KdkPSlts5bXbM3YyRhm8BhDjr35tyQt
HnmaMJA1RLFUgUyH6JMfi84HFuh9QMOoCayWEhFjyGFBRKXdN8brjzC2Cl0wHJws
BAXmKAIRCSCHpClT9G+AJXAL8cj2TOo/cjYa8gizHOXFF2SedkQOd1bh3H7Lj35w
WQuCWW+7V1U0/nWKlhKpuKrYZeD7LM7uzeYfEJHAPMwEyTtY81wwE3e+h4QvLB0G
usHkFXojxFEwaKy0zowOLjENmyZmh/OK7NQlTrXNm2cPzbEIaP2Yu5UcFBtMXiVs
1wMu8dKrDsGsRfeTMhDwaPd9+bJBAlUM+gj979fJ5tpwxiahWCYDgW6gntyY5Gu+
bSCK8phF7MoeCFxIe4jKlJbwaScwIPk2R6B+5GC/j6hLQ/5y0SZ9/dw3wSH5N5Dq
NbFm3w3qYnWBwwU/uREl/4UrdDyNcnjclmEOyOTgmrK7S2ylCRBk7P6rMs6h8cFW
M96gQaU2+DqLtD+ScMNXBzfqZA9BgPOOqzoSV0ikQAf79W/h8yytXn+wy9nTIafs
biHpE9yeJqunAl3TGF2zi/PMdqfPcqq2oR8iZwU1G9E59j+JVSsieQiJXmLludwz
siIeAl4bfP0j0x02vNOdPoyTSIM9v3z76rrMnx0PX9TwU5WM99QFBstOMGSfTTWA
JLhDFB3qUwjwjVU8yy6KyV3oKVzCLS7BWEiLUMxJ8xLQmc+OIj46RabfffvdzySk
tEtBEmMEUYTVxkrWTufWJ1tnHlU2A67QoUY3fammWzjfuabPzVN6voggIw/qyNMq
3iGnkxpB44MFkwUt/3KEAw15cSxnA9St1Y4fs9vFaAyod34y5MfR2bmAvPD/namU
XwBEwa+xZbvewlX0qsS6DAf9Npv7VnqHIfYDmOmpY4VJLUQyJAIER5Tm5EIIj4bF
x4xUhgqSdhA9NFQL8aTuhVPCOXr8tUXtzXOHGdoRo5EkwFpEX3D18To3uS6M+eVP
/X1mpix4nQ7GvVD3+tK7nTrxdOdwtrRB5TeEQBNRVUW+AFdNJeUOLbakTCdZ1vrn
86ULM/WzcDrmXKUzxf2MWPVtwBOoOi2yCL9+WF0ADb8cEnmSQ+AceuN0vIiGhL75
zYs2ZjTCeSp66gKmqd8MrSbMi1qXUimthWBoFHsEwo6f9BAJG+Ws5su1Rxpjtpw+
3m34FQi/761ZqJlFVGPyv20cXBsDVUNyW1ABR+1GebPFvknBoHXQhn9Qbg+NdDaC
DCCYUoHZRqEuYR45rDzLOgTDZbU0RahkAMAQLnF4Z7cEIm6dSmSa/oXl53JWnXGn
0Uk50UisIZAXyKgutqJ4fvh0jAV9Wz6o6VUqPU3LAb9q7UBhU88egxc36XquSnUY
kRNaOKUNDxc9lVtX6hfLvbbLJbi3mTBRxp2tYuPDZV37G2ibXOHXeagJuvgeZMzK
4/b/n6xW7XhxiPGnUwGERXuCMFb+BE/wo8XOCwZ1+9CsBs/d/4MIFyNygZM/s8Rp
uakHXp5ho95qj1FshJKuYsJ0XtPkO8P1eIZeIerHzrk68NzyNzxEj/nW4QkvevRx
bQqWzMEPnE6UA4rWzGXkuhynT5afj9kn4EVTmnoEpabTDKEtpBwdjMaHMlk8RHlw
UOxZsPFYQ5jcL2Ou7/L+GyBvJPU9aw99pD/gNJXN/cLqST6gfXEQ91hNguZ/ustz
e9UWIUNG3YBPr+Z4YFgwyl9ijclSslZCKKYpYJtAMMeMYNvMwUr/eQwlzCd1F7uV
UuWQ7xuIxv4+x9W7xD4jy70HdhVwVS5PFunhHsBYbqmdLBPtwVrNwPxNiCBOf92I
E5Tuz2s0GfSshIUeEztBqatRr0BoJ+vnX1L+SyEvw/PLtxRqYj3GP5xtOzsB5Lbq
E9UEjVvOdVteDTWhL5SV5EaWnn7VA70gwpKqmHDoMjYT7Acr9dYXOIZYK9KnaYt5
KxF3i7NTFYyWkxdyTTejBAPVQ6yzIUCeRwZbOxptvjoS7D4UyBEmUh8QVpRq08Sj
Goe7RS8TZXCoC3nPBIEx1Z97JQFMK6TXNYmZmyZym1+Iq/hlRbuq0VrEtEFqbJik
TYb6y4aeW8lW6aR9yq5hBEeytd+hZENweeA6xOt2b8ENRA1Cg+o5R0gXWWLY402V
NQtYD/X274jRybaipyzx3XVI+ecqXToGElZ4wj2BCTLJsmffduqBWIZzKgmKlcLz
GPl6qUorhasqMZIthmqfKHd9SNjzV0oxSfjP0p/NK9s1ifVRbIOFl11V/JccY8yL
yyn6bgKM40V5zj6cthjiTeDdpEBbOb2u9yDYukviPM2IEVMs0IhFFudXgM6MhuuA
IvFRfcH1M4gs1fRStNPqtD8jQtZgFlTwZF8cZfl98WAO8vJDECv+vmtlk77heFLk
AYNJTza8iLxgDyzqRlzXn/8LWstHiinTcWIneamwLblqi4StVB61AOXU92GVsBSI
clScKOVNyUYEJS0nLWbhYUhnxmaQZuw73Wn7aZ9Ttg5XaSPtB+jbhNoSO9ZJkQGF
M0VV81q/CTiNldRR7BETGRP01nCrmu1oEv/IHQzv+1ipbfe8x8AhaScW8oiHJ/mk
fh+TTdzWwz4C0wWbQxbqKi73hD05GwqfeOblteKHcsvGUJsv/uhFHmPi6MhudSHX
TY/1jxEGjsDyh5kZCQjf2n2qLkVmVvUDUO1VxU3FKfrcK/vI7uLZ7kz20WDpJVnM
6UYv1dOBZS5xTUL5zmL1QlNYWU2rPXP7wxuG2gGE6z9wYGinK1v4wedRwU8EjKb3
cP9mWUH0tcYB7KeQUnOajGGOvAasy9ryhwINWjHSEWthLCn1J5rdWH4zd2F6Agh4
3crk9Br8LaTmOJPMXd28AVhSYEW7XXJFpHXF0bDVvacvgssUvH682rDiknI2ege3
suSM1NPoiK3AjTgIkPVXuWWbNLmzHhJOsm543UWN+iMFf4u+GcuPthl6n6V51WeQ
aDHXiO8vSek5Yg0WEeycl2HWLkpeuRd+jo0G4TEsGWPfrNOcPR24ULmCLk+ncicR
+io7wuQ9f4fP6pbsPGZAbwGFo+bTaX1R4L18fiGUXGPJuEYgKxuO73hnbELNFEWe
9JKcx++Fbi+S/abS10p7YARRZECjz2oOPZm+ln80BZPP145o8gSKcNDN4bqpwmYH
7t+Fvr66H/oqSbmEDKKzPlFQ/yM+v5/FsvPSbkvwKyEgir1EbhHRkvgG1J9ymWkb
Vkp9YXIuChVjm9A74KrivV5cmhW50qb8czoR6CsvYQz0GxQNYhT2bCR3t4qiXilL
7IozG2Svt67T+Mp361llYSULkqe8ElXHgQI+Gt5cqL4kga0uE/HJW+qYo9KcI4Sf
5RYO905NbioQQfy5hp1t6vcvWVc076wBM/THNfejee5d2TB+AMtgxd+qq77k6vjs
r7Slt/7sISz1p8fbqQkZpPPEN7p03loHe7ygSIIzqsbwlJvmlsjMq/rtpvfo54U6
rD95d4+6HpGK09MY7ZGpHNxL1TMzkovTaK65uzJWmzCglQMgj0bQPJYqE+300aoI
hXepQJz5MApLt5PUGyeLYqJ/Bs9b6Y6Xrcftk+XBwroN47dEstCXr5Cn3RU9XgRY
Yei/dUz5M6biHsAhs3ygIuUGlHFI2UJvxWPM5P4a1ZICBbaR/CdLeMC+FrAW8CN7
wQ/XYMX8Sobwx04RzJPh4SfTk2BSDe7yK/TTOkAlYbhVI+kNKxMxp29+kicWXpNP
8NyKLrvBubGutuFV633NaTVmh2tlYL4+f/QA41ZGSNlAz0l+eLE0aEKWbJOW9zwT
72rOfz/nEqxIMAp7vgkUZQ226X7oGvcwu3IKHBbTqPW0vW+b1eYBFfTyBbOdomTD
1i7DyjDNNBtCWSQdyZuoVyu1+1UahX08Sm9fB90zlEe8OhdTBE1jOaRpGHiGhK4J
jbmix4iXS3frGTMEUy2pHg0X3MrtSD9OB77rGh6Mp1ODtFrNcJjq3Rm/E6WMK8zK
ntxYSSSc2NXddyO2DuusssqBO97UrL+fN3WXLVK5+bu1ZCwoNaWhWZBqPqnQcJ4d
IQDVAkV0iubXw4tmEDEFVAav6jHt7CumYJnKoLLeUC9vVSUAvZ1DHRaEaxltoF7u
Abvo8Df8DIJ0OLldiFriyiSzEoiZCs60l2iugmdKMoAMvrU8bMTLXAXRDLm6ICSG
KfdBMdXDbe8g3li2vp2sksoeYQ82BXNDAOI+BgAQbXu2CbT7/PSgnPJDD6eV8wPL
oESuShOAbXrqT7O8D9niASG5DDXtF6igzeoz+klFcC53lqSspyiC8jqxeLH05+oq
2HLkWwm3GBW4IXOr9YkYXfyqVPqFGWBmH/sUjxn/WHVf4P89dU7eYXl1zmQ3XA0o
rXFhxHMBMtXKFQN8gtqTBH7r0cbfAQzchaznzEeoQ4ETdY6koaICmgGioBI7fWCs
12U7r7d0TCTGg9gT0beidmkAJP6qSut9PyJZVhgHMj+RzHajyH6kQJefbLDyWRt+
zE/ntBpSyBTITuE0O5YpgTKOtSRVUva8HOlgRsrhJkIPWmjEh2i9dZ9wcS1HGB41
wYYreEqLJ3EpStRKo7hniJMLH1G99lYaTGkiQhZhJsufojbS/IijoNVb98WjAQMs
KDqLPae9kD+m8L+55m2ZotJzMu46625nVRw8xaFHBSAP6HviyyerAhEWAU6xyxbc
mHGXXUcF6eh7ahXU+73sW2OR9HoC/FYNvbq6OD5fB5MiH2kEDV1YcHVJ4YB/nmCz
5LA98HN6GTx8vwDS/SjB2JYsSfiCq6Ts5OpTDAbOnAmRJiSabvEmithY4dAi3JPT
cnHyoxWEaJlQEo+IEh9Ry1MRLUL+hpoaJaSDuixYxefIBn+v2ozatVoTjlKgmIvF
45+uwrH7R/fD+hl6N3CucWX3wLZAx7VnsOIV/3pS/eihgfwvjAcZszVibdDd40Kv
Oxl9DO3HVPCIZm5mI2uY6kLWxqpmqWJAk7e+mtB9gc/VznoXYebdL1po8gCrFZnd
+90BSErfKJcOA/zHxMpoa4wIZvxEiWOqh5DLQ654Kh8OtODOlYAWDuKP3WPkzGxr
ShONXy63HvgxtocKRI1tWqSJmS/Miu/vD6isHoQtN7lsn+jyyldshtCWGBY0dwxM
dtrA9KmHQYwbe54LvvXosFnHJDqlCKOFF5ldyAohmU3th6Ixex17ay8LUwtdCGSE
cBMJIrPNE6BXfh2cjmhwhz9rGtnmbQsZwLp1yQDR85/z7C25CG3idtBg6lkQx26C
IdYHQzMqzQ1ULch5VyHQAd3vfH8kgiaznQelWap9D6yFdwDHe5OHfEQq+mZNZwZS
pe12E5ExPSAl7zjfVLbK9/JK06vltyIQmaL+kUDqaE8v2tt7AeA9URmlFBlM3ZjU
Tki/+u235c/aiGUCNEujrhUw9ky+86NN9XmaTUr8VXiT500z8FBrkq9YJ3K6Et+R
fB910P1G3Ck85mF+Rcc/LeDLHasS84uTjNdUr6TAxDtRu1tK0DyHQuFzGKP26lbk
235rTiPlpFDp+/qQCAS/oqexv4rWsO04TFEMSlvysAblCxUQBDxhI++wthk6h+du
revHuO1f4C2wfjT2SFsHagTprJmQESCYTxJYHlcFZETdCzH+cPOQvEftrULLNYnc
UuZvndlD8BFPKcCoZvEHWDlReIYeBKLPrYVZVHQcDVpv8GJi8pgtFdr6MjGyg0V/
nIrZMUhiSG65Qe3rytL56xstZfhQnCJPqzj+0KWxdhN7TyTGoo4SC2UeiHcu9z64
M95PAAHixQCq6b8lxWeUUgvhHkm/tBqusRBONSp7slZlmsUC8wnxfKeIDPNee8O/
xlGHnba/t9OdrC9tjukYh5D4vV50bQIFqN8SDa4oHlU8E6iXkJiaPlHCqvQVDMTV
R4FajG5XufUK+FLbIO0pxRlHiYnul3cM5X6PbluEr7C9PZl+0+3Oi0gOZFH7/YRE
IVdHbaHh4Tle+OmnwasPPPdh/ZuClbppMZINib3iiYaYstbBxMOOE764SCWFv4lX
QFtJIhivbjeGcf6VEZNvmuZXSTmNoWm3frfXi5nYtanSuB7AZxT8o3f3NmpwKBGP
irPyr6FfGRl6CAMuJLbYW+XYjs9E08K96nBLIr6WnaiZ4E+LpJv7zoCsuLWh8BVs
tziaiN2Zz2x2gCr53jPkGJwHRTAtNLYzMXgnCexi11JrJ0WGfY6aqLDAc6kk7OOK
H9fBn5jAfaCN/duEVCRg0hqDVA6ZSfHKiXkW+cWozeRJwRjYS7kUlbiqeqOlEf5U
CpnK1ypIbVpoyarvUihgjnaxcWKzOR+HRufMv6/FAZCF2kcGp5HBRJDAKWl4bWhn
i2E3hC3qOnWyH2CAEFIh12qMZJe4QW0ODW/Q6VA+hxklDKnCS4ySA4IS4u+NXgHx
Ti9kW4cQLn7WsphjR9tc0R2zv/ThCugAqo5+CoRIpIZU5GWhS2PrwOOgKqfZAJKG
35FCah607z8/dFyx9bT+mnqAQycbasawfDgxxeYsAE1DXf3lQ91FIr1khRfezcKP
DHjUVbmgRi+z33zJ8yBSKkWM5wXH4ONT5tNjEvonrnAAyW35kkL3n/zfFyhz4xEl
TSgdgjqB3+CyXQ1olJSy35V6cbWbYWCUCkbSt2Jsvx2aJ129J93gPBMHT5eZnLIA
3lRkhyCWBiBPRstJzueoxaxjImmDEBfbSwI17gHaYmSHKdC6ybKJyucWl5AH5/E7
EYZdZJy1fnN4eNMw75XOOUpnMVmH/k7FhrZINF5X1MeVIQpS7mXuOCJh3wmoCN9M
o2boa9tkmongSGBn+1yS2PxhzLdV/e36P8jn2Or0LSTcEmetqgeJPqfimt4FaXI2
9iqodqaiUiLg2L9ZVsu/rh6m8FZ/cba6Wfrg8TtAOxvVtHu+EKcVOKQLFum6aJMo
wJYEsE5lKJYerrtoNXnWw7pPXTPS7p/1CSUQZL18msgc7ygXDUbKyW8Sfj16AHo8
sqq9pYK5TawdibbE6HCjHdv24gx2tNUBUDBAJV+qBAyuQPenQTuYJutV3pEqiWnz
sh+7SQ6HJSMVULtdmV1a2SRc71doNEv9UBYZYRsTq0+92JaUQZXvSuzS5HvT7E9E
hIh04CcYefoezqxJVMcyyiTgzODhJ1pMOPGBaEuCSY57+fSUNCsRckGzluEDJ9wc
0zCvYK0WWglYbFkMZ+K+8xSuUJosV3fC+0kUk+PZYH3qsb6OuT3l0ba4jg0nbqnx
/U1gHSuUh9vMboAHW0zGne+F5ZJTlcvMfL05AzFjk1lS9lyoJ94fEEtn5IIyH/zU
213RWJ7zckoZTpOh1y/2Mh7RatJLuZcRr8nXjRbfWv4QqcGjAdZkP2MNkBljV/ec
Pf9ifaWfu7WPXlatT0WiSUdor33C2bdeqH5sTWP1QdrwgMu8BF8iK88BpB6zo66h
ggotiJQL6iwoYzUDGyz/XaCeqyX0pjpv3OSELTgEd5N4Cab/AWzXQ8FGBFRLXeam
uONOCew5t/FN4n4kEWtJm9D90wI48ap/RRqVb1b1/MdjVEhzH8VrYCYv/UI74Igu
Btf72XpnFXwqWWvkSEJXP9Jwo7rvgx3Ycu47/uOwqNhPeylj34NgL9EbdfJuQ0Lu
TvJ4cWxHQT/vaRbqU5HdJ6eniJAQg4kzHKOcTAEGaUiirtiZwq/w2q5z+NczDPx/
vrJ48L8FrifVo/tlNW4eaDDX3HWvjnifabxEY03pTyTBrvzRSrMCaGBYDIhaEb/2
RbzhJ3Mu1H7DJFIjCsouf9AlNFtE1TGyxh245cVV4cmMTOMMGuOPQUNbp3g3ttDh
qMF0kUJGYWg3Il2vdhQcfQUbZ8NLAlPXA3rcwZcurIT/HWD+Xe11sxhp7Opm4STX
Yji3ei5jqygnhNvZz0gpzgl8IIY5BtV9zJnADxvuuf/ZUba1LW0R18tg8g2Bl9re
zOjpISfLyJJMFl9lTnroYpx25mVEv4nEpLBe5xs7HHnr8wfNdnSoSDgSYv70Yf23
NRTkSxolV0eHGk1WhY6m1CcFaXWYu95jAdXQeFS2b0bGbm1W3umUaywl0cljdcGY
/mqqC1aL0psw9e+N10COh+VQzbaQ6D54jeI4UafdYqayDGVzIXqSU7z9lTgNUQz0
T4fbmWEcHss4H/S9AldsVdLuL7MOTBBLonYn0e2hLKV8lawHmUU9nKfLAOIqI242
S+gxumYeXHsMjIBDMb8KBeXUx0PdIPMnvyHGQ6loVawNmxfqLiYRL8onf0ZoeECc
N6l0zLIrINTJ7sVizi19i6zQb7hA6rpyHXsD3wg6thVbyGMjeCVDrUD3CAN4dKRx
sHNja2LmwDp+Bzm+uCv/xuDEO/0EJItOQjQeCMWETHjFYm1u/sUsU0bx2BV/qsQA
Ef/LU0b4KgSITvFwuIPphuq9nAX3sZlBJeBnIFV2c6R7xNrw6LTclv0KonR8geyw
Lbyg3CzbgYa1q3Un8qAj/pPPLZUEosI/S/uwnNbTuhhbJ4xH32vgc/JINw0jnRRk
88R4iLxi6RrwY1gVqBJtMJFmtlgCAkXbXbP5CNLqrJT7tS4dVb/7uRMHvV3EG8Kh
Lf8E/RGuvMbPk0l0q/Q3yqdINJSJrlnUsPiF/nMel4TThe66CfWNsD/b0MmkLDti
tuQcAwFx/rGd2lEkDpTh0jusiPMyK/P1n65ZECe8GeYiFUHGXBK8dWx6MoskfsXg
H0gd2uCMhBFyheqDzr9IxAJ3F3+D/eqPNAOJ0ObXXodSG+SPXcJpghf/tfyYOpzI
HY8ZOcrDkhSxpVZ0Z2xZ/KMzEpRQwK/8z+uDLkAnL2htOD6CApRnfKhIJ10ti339
n4a/i9A0OwC2UiFEoaPgdYrvxbAbCN99fvIy6MthflkgNTV7c6SEOmFUgMltlzgn
5zqdgrYASCI35UKLDZ3WkDVWVfIzlOXX+kzd5vffZGq2TIDxST+3ndxoXhRnspPN
RAykxuXy2xmP9Zo//rdZcO4gTUcS0QE9no0Q+UJMq16XX5OlJ6HLnBPW+/OBB+Pu
1qRvhLXiChu/FXAUk2DJSKS6mJDMNEax3qSIim/COwMQWki8OgcFMyjkgrQ4hSf8
UupDdZ3SHjWdVzcyaqi/MWY6jFXhToDKQXA7+Ld4Q/9fLpXtmxME13QDTyrNdM9U
+gYqAcDDRC4AaBNO14J70UxSvi4dpg7b4f/5l8GM43ftzH+hrSsUK8g0qOqvf4wp
mDBwu1id/aHof5s5GhYd1b66/UAutF7fKaF4jX6lFo5MLJ37OxGWQQ6Aw4W5MZRW
XdCTmsg/7KuzQvhroMH8wGMp7zFGBfdNXNxjpGigC5Wsatt3U2S2ApuwQ/C5Dfh4
N/g8kfKEO2ZWo0ChCPDDNG38+XBhWcJ34bEVdva3FZydNz7YEB/ApyYyYJL+LnAw
zx6LWig6HntoPdrOR0lYKVaT+Sz4oKuSyZNFh1+4chl3FsSZYa8sf2K6fryL6Ukz
DR7SE6AE3OC47QxlXSVgy5Q/B1K+Yi6JfjJORxLB5LwUQSqDo2aL2YMsaspjVJgK
6a3a3DBNItSrxUUHTfIocM505Y0Zbl8FNcWj2+p1GyWnn87Uh0s5U77eUqjDXuL3
prtifgUbkGASQVB6nUlF1EeD9s3sGr7q9GGc45CcTUH2282/3EqKXTugDE1r0eQW
tmgVkL4ZYULYJslor69Wu802dsamuWRxA85J6BJxsFofQ8pKxfwOXM4o4co9O2dZ
xy6hKSaBO86lbBAdqD0z09q+SYTivy4OZ+h7rzo+AwOPX1Vcz1ZAYrr+gX1RRCZW
1b4s7o4lI7hfePEi0omx3Qdzi1JOIZoQq1vapKwxTalS/40hBuwjRuTDaddZIrzQ
DhQe8l4AfqUheTgZY5bKEyCGUB81Dq4tez7so42TTIPximS4BuAxFxAm+qNwWunr
EMMMWwl7gn1zUGLI/4tkPqtZj3a1RD2ryMQiLwGrpe3szYaYpJE9DZp3e+m6Xm9Q
Qzacw1MzAbxYL9eAtwg5wEsP6oiMEoi8+40tuh8zaTRfriIYQ+WByxhEhLtM5RiH
Vg/JqlMujYkGxzWSNF5QfuE2Rv+VDm3VrKRp1e9lpZpEDU4Uyv0kDJoHn5IYNp9d
KwmUoXtZkqgzg3ATaOvWhdPlxwH/cb04ONh7SsbKmJkL+U6xkQExDHO0wWQh27ax
1xuyT4FuEkHRUp4K8BKrdLIBNLzyZ8IqOBAdOG9lUlKgpkGP2IJbmFgOcNnHBBQb
KzRznBb/+3z++8MrLipO38NdWh1w955C84JTSLRTMs0IJXmnpEPO0pjs99gWK5Eh
1odtmY5wP57JnnJ5Cg38UI00Ud/utAPOhsejSqe5PUIGK6b9gd0YIXzKKCSf8ka4
XwtbXAPbnvAJNSd1vCHWtj+muNisT34HWc1rIU7NtjpTAzHpwAAgrK/Wkh/Mx5YZ
hFT5Gin6/LptxhZczKiCRZwWfbcyP+EpfKsT4gA6eFfwUWRNGdWFM/J/b0dKfE15
Bmd4rKIeHXUu9eiGgRYSVZoThsr/UNKMBZ64+giNXXiHDTNoazWQb1vlkKNujoMk
brepo/8+0uyH/SsWPkfKti3Av+943B5ZEng+BKSUnCfaEsCW5COyJkGoktn3QCTu
a8xkmFmIJ2yIBJX8JPqhN+KAy3icwuOOsrfP3Qzf3zwe4y3908ekYyFC32AQ0Tkd
HaFmJXjhQQ9qh5kouocyz0Vc/m4uODzmgwcDwbY8xTuJ5jRk6od2JvEBXlBfCEjR
G3IQ9AqRgqYuqTqXOTQ5iy+4ecwfVrrGm52k5cZv9fw7xoT5+2e1B3UTIfLalkUC
otWvPsxAeQJHTV7aV1WuVBM/GxjR/HUrTiqQb9cyRz0PsNla7n9e1ZcK1f9eoak0
a6CU2Av9NzW/2F89FVecgVCrgevjzyZFEbTfATJG4OB6+AW+M5RQ8/3aAgLZKk8J
Yejf8tmJycyoyRXnkR/qmz+ayJ0SnaOgh1nlXBrcvycUOlaYVGSJsGeXk+rw/wT4
VMm+TBAyeOu5UOUz4tBUMS7PRvj8gRT3C73StydewGe21jPqNsBE4A2CfZHZ8NsR
jTV2VuAtCroGBdVvJsOQ6Wu9wWzm9y82hozxIemx40UVss2dqPj3CQHhg9O2qoro
LcLzMu3+5+ZbcjZx05Y/PeqjIEKVdQbn9EeCShoRpnkUxaOxqr8TNIYD/rnGLSMV
Txbc8NqlbnWrnWEer+zoOOVU4MgaJXuG9o7ZZYcCpLrXufRR62RbpQ8x5eyjYwrA
JBpYGWKn2CLX8/aoLPfytyKwC53ehUeBEmFALSIqtemTqZnOxu/YYgLH8k7Iw0fL
Eg8KLkSHiDn+sX3az03kd5JQZo8mfiDKAzi8gn/zpbMDYRZvz7dJ3Mi1IjK67NrC
4Isrz8dwWLZS0U/ulImyhG7286Bh+PLDezSyit25YkkYk+m5lCfn2y8cu4p/rOOz
yUG7iwZ8Q8PTApTmA0NT6QFpPbOqCHSZTHFliIchWE7c/mOlXmlibTPNoh+P45L6
/k8SNOdPFuNRan8MFeABDevJHZiZhSyP3DSdQN0qKAAyBWUncc/4SWVYMZ9SYs+1
fPCXixc8IXWtOJwaJuUNMuGSOjJhtlMSo5OfpJTtNjts+xGCxQCNKSQX3GnfAjm1
9IQwHcRIxQGmBpzSyMC0Y5E4E/Bw6ryzVtux84ILR2xN9fwU8Nb9M7xeUPwsmQWJ
o+vorU8O2Ifyz2/3f67lCF3HuFm2GHbYhMgM73KGlCtZ2fgjLZ6tyzCzM0hECf1U
V/0CXzOoNfOz1K4Sxq/NdEtzN5ImMjXicHIntCd2V9SwdkySOAmLCKzCIo7lUpCc
f7IvKIUDif6F5nVT+fITAPMGgJ/wO+5kmwtq9FM8A+QPpyjhuGdfjOwpR+/t/n3L
YUCnJEgXpjFHZbwyOw20tMZETs/Vb5rgY/mwdFzoOuXy6k440K9YYDgC6aln14SG
hylilSP/Q7RKojkG40tBd8g6TLDz9bsXTS8VBdaoSrnx6b2EX/VER5uRKihi9UWL
TW0/yOeA2tY3SHg1dQMZNymwtSJJqRa8n95mwGTmt5z7jftD3+sI2kV8DvS6l7VN
DYM37dQI3toohhVxkFWYVzTuivM9jp6laoetlnkXoawg/p+BtDt4euQ+NwVObtix
oneZZhxeIjuGFiDUpmVZQDIZkhH2pBX0tCTFkY34beoWqLfC3DkFZYlkNK5Z3wLH
Iu2N4u+OoAXFbnPcNusl41Mjqzx/JOk1vOFtbO9TZ0rZXs8wZFX+3st9BLJ22aGG
kpDyGHC1hzAsxkIrgdSp+rlbvsr8NrPWAB+o6putI6hTMPrF5xS+waSqLJduvz9z
7QabfPjA0BfAsL5fIC9w3iK8SC3Qb9wyCnckV8IhArZtWofr88oa7Ox2wiJAfBGj
9nqJawrstttv3nXdZ5kmgf9MDMDSqT2MUj+CLOZ5ikvv9/25e43VyRr/GO4jjtGq
6gHPw4iizSwT+yD0vdeG1j+r0uTHXp+0m/0ubmmKDcTK6OVefWul174qZcx4IzSm
fH/obj2BU0gO76N3631+w3spDICFv10VPQJf7Q/XaFfC24q1pjQkdHqyyeQIuNzs
t5Exg8VKpii9PDqh0DRkx20o/O6wDnwLVLLVlKuccM7o92ckJAhXAr5cM+xm/Dez
kbyeSiwKL6p0/hBUFROWHujy5ccrz6r/RgEedcoCC1GfF6gJ5rXeV3ZeGhb8I7AU
L3y8cFGMQkfJuaJ4lW5CHL8Qq7TB1zaALH8FqbkhtB/it/TVnC6U92HmoZ3FMY+U
hbSukwKbwJ4Qd6PNCHbuCjO5w0fy3uFMNgZr0X5jZuq1Y8ckSWuIujGcjGsEe9Vt
cVxNvF5gNE5Tf1fEG4ifO9LZxNx8EudKi5HZyydkmlXRFzJJfVoLbTPwrfixuCer
ohCFkI2QG0EvlPUhRfOXSnVvZKy1yzuq7vYArgIpjHUAl+EAj/neNs+8v4Xgc01y
hq6X6bQlghAW2cvNDftnrFmiZHWEW0cmXSR7g2Hw6Z/hUIdZbl8XGTxBzcgbE1pc
pJ+InTMrkZgnoA1azr1OSAbmAcZYBgjxQrd3nlFU/yDfHeCQ35dce4Y+nno3C6s8
CL2bTGdBSvT6PWByTK1pQU055f5uoXVPkVZdycnBRLCix0iLSOTGsP60/aoPkKnD
oUFgHEGc+Y7jqIinc9pGxqopLA8eXl3SX/2luo5hhCV+NgYS2/PtfRay5Ip8DpbS
JrsWWyxBxWcdKoWM+V7iWwx/hsUAXiPW2MDHVuTlMkgi3N1k+97CRukZg+adqyed
xwjExxliBGksrrQPafDWlI+v4irPYBLQ8xy3HTkId1gbo6V2x8E5kLrivVsmrlyU
SpwSztn49L/pDHPK1PwQQ7Mf9A140O5LOsh1KJcgbYE1SXLOZj/7OlIFh+QHkfYV
HYODhf/e3BMFGUW7cmJnycPxuPFHlU6LsU2s16baJj1EMEd0m4TSjhFsZh14ddpY
ZIy3Vjr0jK7pUo+TGpSAYKaAXAMpHyLQwAxB5fhHf0aARcQauZKFtsiicO80fYEW
aMENJVCeopjaBRN+bsVW5X8htuF43/+5Y0TEjJjTea1e6ZdZMHX7LuVRUAEcYVKS
KhLXa9uEvNSbSijZMsqiq9KaAZTsvpuPcaP7aZup6IdbAZyBdyxlfONGHqmpHwYT
malRujMFQbCf/PTivOCGG7d8issy2AOdvmEKymZoeTaWThANdP1HwIfX1hwJHbSE
JS0aUTxWY0wBnkwEEqsCsGPavprEXF9eAME2F6PaJWAFoEgv4SZ19az1wuWZhpaw
HRLm0tnJhucK5tqcBAEmhVpSjV/mtSaPkJBpdn4Zm+bRTNpWIR9Gei/J7BqWbHNG
sI1wHNev3jo2DUcOdBuFpcmkoG7JrhPBjtvl8bssPW7mPrJMnXuq8/7w6eEmIEYd
LzZYlXxq0lDPbOcsB5fUMoX0p1vBVSlDHTuCVyGnlorzHcmndzHD1Q8wLiXkgbaP
Rl/RptQnvLA9Otj4I8vLAMwVW89kLZctChZhfZLBtHNnFJYMDsQEfNAzMFi4V+O5
GzLm2O59lt6Y42FEEFh8/QTHTVbSb+sWacS3yjW8Q0C3fhkn5vwohp6+TnLVFI7s
W+E7+1ZLacsZX3OAIIOLBnDp1KuFgdeO2t4nHkF5dDolBIk2XCDEigSmeH07lkQR
7XLlj5BZ6BswNXzOHPpf9apA1imbkpik7XZklBek+/ZHzwfSB3AZESKtH+MT8Qos
WzZjVpSNX1NLTZZoTdAnSnAM7aaWesIReFT6H+peby/S/nwwt8Unv34iIrO7g5n0
tqkhqsfNMlyZD0YfwuTzBHQvcau+V79Ct/hShKCWLd+fe6XB0rkMU9Bl9gI8FUXn
SS/VgHvgvh/N7/Oq6GnsZG7ZfUz1t0i55woWBoz09u8o1IPuHK3fI489S2LSn6qT
o1KUxrZUTeinfkcwUWSdYUxktZcUQjY3xlWMmmzyVyVEwjoDV0nU0g8+72WU7cvG
rURWoTJLqUZsziQTRlZiVnXMtt+sU5SxtiZYJuw6urucwh0WRB4s8kjzaJlIV/RZ
gkVrk2mnjNG3qxpGvRK7XnV5c7uTB2MJX7rMgk3VYbdfKxI562PdbJcga5aiRI2Y
kL4nlstgZf7Ok/QHwulbU5lT26Sr17YurQSBdy0GnuaMNkRQ36ue/LV5SMgRYz6m
RXgQQlCm9tc86rdEzoYcxgBpiNep5zpZfsy97OJ7Wk64+joYMwnOedwG2ZwE2o5e
64Ylutfl+m+er8O5s14sONWM4KecqktGQzUXpghjKe1YfuPF+vsURE6zD8pOCuHL
q5oVGL+Hkj6g7G11IYtx850RPuI4zjvIay0d3GD3hb0iMApNfZcd4tQ0ZwI+VeBS
gR8Zm8lmsaX/8oo8EQg+bl2fNSIQvlhbMO0R6cNcmOEP9tgh2tKGMC6t9VY0mNlB
CxCq9I6xhvBFOIoDfSGiXiKMI6ZuoiJfDfKmm6J+BgSTszzFvRvTY45y0Fe7f/Qr
Q0rzPz0PIpe/H63Bdl3hg8fG6MLmJcUEO/+ZrHlTSTMy1CoQMB0IudGrIlyNqLl4
846nvdOdlbK3FpVlooQFOkObGX1Ujgjl9hYfgnJykUiSL4rbunj25lu3rNwIpozH
Xm7Cgb7dzH1CzZJbyZUiy3mab0kJumx5dzKtF2JdoSkv1wxj8YiSsU17hKWnSftE
jJqvFgzyQP3VmbULfHF3E3Df38hZ397BYq2Ir3SfpB5K03du2xK34+1SLLnj3JTq
N+isIziX1IYpgNQTCsHr9BHB7VDn6IgFBap8ubRpIlIsNTGZYJKETdl4XcyaU8H4
eUvS9S0oq8WEzY4sX9/eY0T7lXMSOGJiz9S4wWQt5o9xgrcI9tw9Gsj9sTvXWKvh
p8eUb3Xz9Pbq+CCvrKEJJzP/hnN0ijBB0t870VfRfu7A5EWQfQ95NPQRUhcu6NtH
aZCUuW9S2nT97ehfWnwYM/+yLFQApSBopZJ4t+KKCPkLMzivkjZ6obUwh7GTnmPm
qj1a1sL+YK4P3PhHEqNUd2wNjcASgQ96mKg0K2c1gY5nucWAgTFH8x6P2RvxYBqX
uY/J5O2nLB3pyFRMPsGdwMvi8PemKfXTugRbojkk38iXJ2PECCSvVis3/yphWaPn
orb/lISghfAd/nPYIKcHp/CK22LR3HxAJLczSl+c+mZBEjnzFxPqsgaFvRrOWRFe
kc3+Xrm2P2aWJJVSBwyVSdwd1HXjYmqh92uA+EqHurap06fkk9tN/YD2ojyNJdQu
mHkL5aieiIoImByJGn0viE+rgQtgGUdo6ppnowVsfYfXDqL4Ljo89qJWnbalsgQr
4yTVDrrYN3TBA2wtISAdIOUTyKYb7v+wp+QeDytLq/tvMBli6EDQFHDJVMqV3Azo
CO9VIgaWliC8NL+AgK1paE7fnsvnmxn/QfI3JDGhyQHn/1wQVxaAWE0KISu8NQ+q
RMeoa/mkn28sRJQuZwg1NiANMuLfD3W5SGA9T/A1fsaFPnBxegOcGW4omXZb77xB
YszXZ4DUbqC3kOT80QLIk7G1MeE137umOFwrwUaRMnuWSeMwByhc3NlghZulXqse
bslVXcFRWZ2QOLiWI6wgFogxXYxLYw7nfeNLyF7kHglvXPjzVdh6csWS7Qm9z/Th
zt6M8LZ+wJ4K7Wuvg+BY0yicbNnck8Pl4mFF8943i+gX1M+1fk/NgwEIo+I1khDn
wGkulmclfIJxVpNa6sW/uKdFfcivGw3QZtPq6JwAyelLKgankE5cmF84yKDCWWdx
admFfAqQ10GizVVlU4qLAvI6rAQxSX13JOEHTykzQ1pKrKKJ72J8VyHVMZHPffsa
ilSkZdUGrvcQjBcVy3kz7LfAyS+rF3aArKIHf1GWelMyfawVIYpWMvCLSIVhDSN2
Qf9xbEQyQ/0thOR16FnswlcwOtjpAWIT7cDoL6yLQXTil2ibd62hTHJ4/mBEWHgx
QYEa5Q7nD38ocGHmRQesD5guah36gkI07EZ7IwgMclPvgv/cpn7mJanEZGp/PJrQ
tIbiXFFvJV/Xb/rRZSrXc/Ku/q0nq3LYt2xGUAxXV7rdg0hQAEboSIpaR5YiyVFd
4/vd78hf1dd8ZNLnfJUavRQ0s2lM1aQchG2Opfub1zrlEeMGzSUW4kJpSm/4tjO1
YKo/2vYOXFVh79DkJDt3kwanL3Jz9S0oWGPGAGO9pgriYwdBc9sd55Yft4lH+wQA
XwyMWHZcuTWiIZJDa1UjH/mEhwLkAzP8oslPslpFlYlxGDdxV+CpfBpsOFnc237p
OW6Fp5rckvqp9sHs4lRakdXVllQ2aYbvfE2ld/jDHLc46UiPJfxHP/nrILms+rk/
OufUxh+mWpyuIGKWpilk0RYf/+TXtgRRZsQMEHDCMSrp52l6Wh9B7xndHts4aYuU
REAn1k3bHtRcJrEJk3EnNgTli/PYVdCKuXasgcIuCyBosYzwoxRhTuaxiD32qL64
Kdeh49/Mb93P6Q1xhSPBFSEqb3AEqKqPFPmlKnIw9sz4d1RDmWdr0ABmm1nRjNrs
vSz7NeHcS6QM1I+0ZYlicA5YAz8EbD/9XrXckEbngJaHRjPAg0sUsqOWMRe/G+vK
0icK04YxWvIC4n3+Zewjd7VI+kxe8KR8jeQsS33g0LVzXukEWTw5TfEwh33ve9qH
OQ09vYvEgHIjUGNLCj+o7ypXms2IGTbUVM3uEspbmTta/0BuSy5FkjrKt+hFgBY4
KJJwsY1cc0TN7MZpVcXPYRvEvntDgXQkRx5cDx4RVbIYJwxa8UZ+cPnj1M1ttBeW
h3oa8lxl2dPfDKimVSq2PUU18CEKbzqMh0+wlIPAMnMRz092T0Plm0PCWRfUN/w6
HsjvNl+r3Gk+GcsIWuiQ48/OB5u9XZgkaGd2df4eie3ah5a2WdP7CaX48g5/+BeF
+t2j0I88W2wE/8X2Vhxdv6vwsl/coDlfpYy5EjjBp/RpPe0hF+OY8Roob05LTYu8
GecuVbqNMdi/RA6rXVN2VYFtSt37h2TQQtWLDQnKTiR4miAz10ik2VFDGImcp379
K3uUOXHaxoPwcYO/nCh0v48ur89jEbNIsB+FIT13V68JCK/qfbc6Hl8Pmop138Fv
qk4hXr2BxggxVpSSHaJUwK1Eymyv3khD9qmfS1d4iVlcEtSPxnFxt1n8QVkVenNu
JZ9Hxwj54/lW/O4uKT28YsAfe2XpFpUrf7ivJUzmoAfow1tfpfDeSC+UAJr8T2x4
kO95JntJY09wv850ZUopafjKXEz+lQgSC0E7sY6SWgHtwckkqzgN/NLBVxu7cBYM
chZl1dEW8reU+P97zs29kbN600QNCqrBB4TqjXlet1epjLMXHokmU+QlPToCYpP5
W3iY1tT4ohztrZsEhZer2LrBFFGcwZAVw3ihmPD+ugvwtIJH+yua9zNCE3dbzVE1
9kz+Kd1dAHt3avMfpw33s6bShlwhC3LymJgXAtwj/W0blLg/OET9N45q1Y/euU4E
BSFPdMrUd3uadoMjb7XWlRbI/WdlvzWqde1keJOiAxOh/MJ6LycZOX9o9P8l0EqH
rbHcNQaekTIC8WJH6nMrKwT4jvpMKv9kGHkUw6r/7hMK1hlE4lNLh2QnvF+qCMhK
CthjGQAFXdKW/5y4iuPe3cFDQLxjipoHzLItupd/eWb4/P1JY1ZjRs3M317V2SM+
EMW52mkh/R3ujqZV6M/8gI27We4Pqm0J5rpZOv8jF1UqNtuIxTmlFk41f8myKeuP
8oqS3++5o1taaXbRdZavhTkPgECDbixm/vm8z1eR6667VkoDRG6YFX47EvrPPBgs
LkOkfENowvy4RjiKbKWx8Et6eCJDHOak642vfLzMTSUV9QuvgDF9+s/BQHeQO8xi
LxfkLPLLJzHT4PPAYTUqI3IyETAGy8VyRjRaaqP1N/FNQj1OrCIvh0+5NrSpZtxY
9IdwVn5HGwOC2rmj+KcTWyq2CjvyWqlFpLH1uJc90kxoQmZBm7ElxjB+kchlQnKz
I2fYgbZCCAdleNXcHbT++ekVZ6l0ModqQWtjsQh8fLQ+7evK0SsKyLT6vrxG50Vx
LLPMhF5nFtytWuiPTOsMjzlajR6al+9QOUtVEdmKOcM2yBfRmFikBL5EVJM5aDWi
RvJqON1qRsCjG1UXVPXwkcbPBN1ooMZ+zpQyMqFVFlJWjEmwzFwkICRZNzw913cw
s4RfXXOUkxvQMR0jVUPWLX2OYWeFkuEdLcZT+CDrAi2I0X4QRuqUUWnTFIiu53uv
oqCTAIfQpHetENg6hpKRNnYRmbnmpltqhy4teOlLOUWaGLDW9L3lD6pNCB1OVviu
+uDvTbdqzVzTMJxOfZ6XvyscZeNL0emayFhMvHnOBJaCJ0D2jG3PnUwq5LretRdb
7C+Iq8zDldl0DkEA/6/VuBR4TuWkJiRxtSUKOax/Y5PrianoIJCxoy+j9dtkwLAJ
u/xUf8p3n5H7hBoJ2OU6xBqGMRCUf2KAznwv8zkURkvC/TwLR5/FMfECrjige2YO
j1hMtupuRfe8xr1wATy7mHzExG0XIZhFMJMd7vxHrV67A6vIeVZ8bMvAhYnawInC
/GAhjs6zkARIkRi9bLejuFv+mEBZ+Cay1KZAOCK/d8fF251vLVMu2jo/5dP+HD/x
zW9suOIBjoC8wiG/47Jwy8CR/2ymFEIfjW+UZenmUOxiIX4UZ9YrEG+HGxEqKt+m
p+eK0n3/NbaivTovVvy1My7ojB+A8DdHPhkR9GHbwRFeKSLj0afHPpCsECC1DCF8
+04OMskR+h8+IPXG/ZUn6jw4jV23j2E157dUSti6af0KLbV/66iAGSiXeOxtlA+C
jvkgYV4S52qCZTwk8uMKRkZooAlohfxVwS29QTOXgO5QAS8IlPP1sJyFqXFwo5D+
CFTCeC5vMF5ntQog90uLhPod0516fSos56xRxGNDF5w7Oed21umbC2rsCsHkrnhr
ijJL9ykk5IFYc3TtcfNgAbYOnY9qDqBz7liltyXJI2BtnDKcRc2LTedRlyEHw7d5
mFzdUYig7z2vA+3//fkNujZK1DQVVwE1x1YKaHW7641tvPFT6ZbpCFggturjgsiH
jzYP2n7NTD18TVZ/VCoG7n6BItLu3ICmRBP1vsg3PauC4spRkXCRZ4KXMFZ6xgVk
oOl6hTieWHMISx8goALUFES/9d1zwUwwF6MQKpxuieZbN1FI7O0mBkzIDrgU+gC6
tzukJZf6a4pR0ZTmaPG0QeYFZ1cqTQrDUuJ3NiHBfSmaPWh79k7lWYU1Zc9XUWlB
KcPd7jAmwfmhx1Kgbh86U2bXWpRF4zRcITQt2P+VNrfDeB6P7wOyeF31iGnAiwDT
yYOVchQwYoJW0yEulEltTeJGEy3biTL+n1u8suqjw+IGDO7dFkiX76ApJnzgPET6
4yR/88dJvLVXSNd4uTtj9EmOplaIsaYK270rXYNeXLWF/gOwVNS/3KnXQRtq+Y8I
N/mmwJjoMib9B7Sj+DS0WoodhCw/qfZ+NBEMPV/z8ZbvEyMwopSFeipsT2BEi1hv
L9Qnudl0NR72v9nfXQM+fdWObeU06wMBf2wevtsH/EzToNi81epRjo40+nGoj3wl
QDVWC6KoIMGoPGGOPyQi8VykoKIvUcKvQrCP0MKYCxBZwru/BVdkayrnACTnYFCx
xXVxh3mITeXaaPP7HaicEgN+PPdDDSfI7u0K8i0UYhYf6g+4moLtpWUs0Evr21a3
P66Z6Yx06q69QdAhu8IZzQXZwYbgWudhrzs7i+8fT66yu6D1Hc0uyp9vGXHb468W
qfAFs6xlPQR/dA7GzN74WqJt7Er88EJM1gQ1s/dZrwQdOTNA1p2VhFh4Nh/SAgrk
O8ul6u1GYX0oHJppcwLrzu627RJq4Hv9DvwOlKVeflEXY8OAan7Ct3wPOghB157w
zkJTmcxaG6CWVknuXpkr+gC/CODTmEYcTMkNr39rrILMJuCg5LES9C8TKkNJOuMI
1n35cr/Z8Q5M572uD6OisMM63K+Fs+jmDDi/5z7DBY1MBunFJTC28ryFzkwLmq5h
3X00oQkoK/7Ls/9DERvJjjSZ5pHOu84phwHL9M0996PNq3XdHueUSJ27cOymtf2K
NTVTBrPyu5+m0xFpL1zbqH29YolJi7sfhkFso7qthM7/N531QkRDjSeONOOethcx
AMzHB7cd/acqyZ4QJFzGQZdD4+5vwTSTwaPp/wXHpwxELwCrNE8kBXGsTxeL/MHp
kEGzzVFebfPigoW2mkOt0+7szarudLccs1KnogvThLn82qDg3z2jR7cj8JosWYBH
rQbYJnKHtJXFse0/30BN1iXq/5iRN8jUFhYlQxMosG6WdwWLV24kA4aDD9l3gqXN
UH/CZd6V+YE5e+7SmFE4/P1ZNgfYaRDHY8NFpP6CZvdJN1K324FTLafyb88uK1LK
DJkkKcTc6sST9AK3qyBYwZoikTIP5RBig1XJZ1A0xFxkVgLtKpXshoY+L3vO83Bh
ZkQGsEEPz6xRJzqNO+4dmT6s9/qiUs1ygw5pBeuuoEQIVlbtJOP/72HEi9cxpiDV
e5H8DbqcDC+QA4VhXtRaVwJDZsEkZJQ+S0xOiYVGz8+k1Ri6Wh6NK9iGQIOzTl3I
boj/6kDYm5yzd5NgfbTb6n7Yf9vXZSlSRknyAH9qhNomVg38MxGSzr9P0R5xPfUF
Fts5UmuQORa2wLGk8g1tZgNsBm+yGJXvgsUmqPPHXHXqyor4WcEPNyGL3zi1OFpl
xyrQZC9q3xhRHHWtNRJD0lBjaR6CptTdFsJ4h3+1LXePZkXYMrRh3xJkJ20b5wnL
Sc+DZux5gS9ETi46oCDLjySkzzjcyzjZfDbLMuYzBWCP18Oli7sj9pg2jig9QCsy
IOHYpNUCdeb2gWcHWAHVxlo9XbR9KcOccw2nMglfK1oQWSbfPTTm5rggVKtNq6/4
HNCNf7djRNvGM8s/riMsLX45EZbDQAh5VTWoTec9HQwjx4W6uQyyllEcRDm9+xxF
XOc5cm910vHZYgEQz/YXKSZWyArFBEmzVO4ma7Z6hoch1kifIbLzX4UtLBm1jHIz
zETVTsiTMk4IM26B36Bnw14/fsFHtkQ7yDb1NHbqyeWxdRuQUt5L7ISFMAn66Kvh
KrZfZeGkxThzbB7PvJGDLS1/Y00uag3M1yTJolxHPT3411irOXKBPi6rNSx/XYZk
Y98ZIN2wEn6aA1mA327SVZ7yFbFGtHwIfR1lIgWKdiGQ7f7+V9v1wah3d7iWtiqN
6gxhV5pAcXMfXWe1BtwUI11D+St6/gALg+uBZW0Jvh/IqVYGB7pcQkivxFEhxAYl
OUOMgl6cfR+Pp3gFym6/cpdIOJV4Ilx/aMaVmy/0tMFJpCDrUoL56oy0SM5Zf9nx
3MMwIoxFUlTmGbx62bftDnz0nZ5YAygsmaKzAAAGiMLam61kvfFBXL0G+SBLMQQz
olPogCTP1xCGdzJMOoJ1nogoQBT98jbVBcp3f329ZYjrKPbO6PZ+l6cuxjLPMvEm
VKqW4I/ypHu9vzmK8uYTD2Fcbw/uc5P0gpgEn8VHNKT+dD4tdW2UKKCNDMJ1pEUY
RnhM1ilMwXoARbVP2gjsezsHC5HjHcHF3kB71sEr0MsY6azm7xdAOtUfeq6+AUDN
SDoNur7tD/eN7eVfuKhYWM7ID0sMXWTKe2VjjR0RaVlCDh3snbEzJYBwXFsAGNpW
JFX02WgekI9RiwDL46FxeZ3LVR/GE5PZAfN93Ppg7BXqqfAkK9PBjFyiFcyCfljb
Z2ZXNqyVRiMQOoh3GOylkaSWnCRd2muf3hs+p+Oge41cxw9bio2ZzytwMYiowETI
Ev0fewCGFPd9kIia6W15OOoSHUJ9GYqaMDNwX3KYibC/DJweMCwQoyQFRbBJt7at
fuSfoWJjkT+1gUXwGZtYuqpwGwqYO8ZN/2I46nfYO7H+T8gztM/mTNZ9A/zOcfZj
EqZBfN8UyxA6UbL2n2VpXUR+53nDq0JOsULI7h+hj6Aei0Z8hyd5zE/DUvAlGl71
kaCCBwVQt2NwkvMIINRy0MfgOY+EPye3aKoZ/P+iArp/EjnaKiAqRaajWSMYjG9b
G4TqdNGbunyMV4LwgBaDRlbCmYI7jYCJdiCNjgUOGUFU/42I2/dhCIB6qMFAtecR
jLFIl01KcRwbD0JjugSwGBdjDIhrLglhfgiUxZAbz3fKMeBZ4HnZ8juufuT5+laK
MRPkgjHJaa50krdWZtMjzftQig5SjoDKSqIrz3W9R4y0a9eAFk6HpjWS/W4ATFLp
fVNC0aQPtWM+ekvbeyfE7Koyz+IbdCq6txkf2hBL1My4+8Q8U7lopMzuIeUJFiHp
iGxpqAs7YJFbBRk15hvLziAVPSsxlmqDm4fQc8N2dtZhmQ78DbeZquY/7NPuIzVq
tSrFm5EYfocNMuOJp/gjwRwvCd/8EmCuDDUTKiE5GGwVvqujPjh+NXccxYN7Cn4I
g4ihMVZlqlKK3Pil3Ugk2lhqFORpVKhABbapE6DA818TKnedsK6NZAMTHMT9cxEd
CLoLfGsTa9madT2e7FmL47q6r7CCwc7T0G9CMj+IUIQwfp/YDmex6T5k+8FmVTXr
NQzsqB/v3Bpwa8zQdA8na8bitdHkQKFZQ+y+SSWSWFLUdJzaCs2LsS6Y/4o/ouG0
g5eHJSLVtoPq/C/Dtgf5j4HUIaNqmxfVOsbenxxRXR27Ev67dxz3MByfHvvapp9J
B2pz2WGPPUKGTz+aT24ihKekJYGszPvDU+9856A8yWc6PfCdKmdMQQQfQcpapVXl
g9dpDFNqIZdNssafmA4790+yGF2WMQ5UCzobAdm2+WPUdXaYiuB6iXk4P3xs4MHF
bVVN4CRjyhDMQryFkq0zZolhdidIlEMLsUL1Dkk4IkjSCG5DH0yVrl0yh5k7qJQo
Cm1v5Tql5fbWoZFCACfnWEy95noj2d26+L3K5bZ7TZdgiHutaVLuRtpVzhc83A9l
NpNER9yZWRTXNs7Cx+E01M7kCvmSFQa+L/Lk9DR+O1x0QihwUZ0ynldJKmXbr7Sv
9fOE0B4RNw51FiCzXtt9qvdZoBSRbCbhZC85abXda+hcrYoexsnIIPRKHOlcmnm7
LwjuDXj48CQtFbfxdzdmxdbbftcY2K5sQuw/cMqPt+Lt7B7usypY2dODODoodYhN
Tqaqs3RkeI+fIP2mPayR3hvJ/SiXJtZopxYrcgCvPygeb80j/fJxcrCMYaCg3Pwf
dFbQY7p1xWBUCLDQNFg067fZ0eFML5nvuYsBiyd31GOMf7gpRImVjSMithvl34ok
iZ1ulyEsYb4iCAJN0ZJIWLLTHgqK/kSZkJOC628R4UgBshi+dcScKHq3OHR7cFYk
pL5yer9Q/MrCDxgW7LSVHEEKhWFW+IC9cPzoKeP0kUg1qzkmEoUVVD+CeDPjBoRL
AFXJHiQBbCGAOPmGHKEv7vUV7YyBjCBWTyl28Y3b7yCUuvzSbaq6aJpS2VU75Vcv
jvKgcCPS4o/ftmX/jSY0m8IMnG4UBD1I/zqi0lNRW4rCLUptHxoHpA2GXUqnP/CB
xjUo/Nwj0hQcKNgInWaY4XXETw9Te+bfdWGCdq4crS71mmy64+g9cRIiKLPdzPsX
gYf6Cm98EM/2FbffGvSPhoQB7b/9TPCmNH+kHvqOY0iRC/nvJ7oazrrkfX7jSKok
3kN/jSmW1+suFYTOqJeHORFtCOzafL3iVyqlm4wiPH1HVfmBAnLjUTX8FhJKUbKs
VKoeeRKC5vGWACl7RgnoBlqWc33zwIG7fjIK1wu4f47WpSNlQct5jOgvTWUoyoew
rq7MQww56w18+jdRikt2XtLyGQ4+M7wJQypRSCIZEAIaZ2H6pYjVBZ0S45lZFcG2
vhto1UZRQI/uZu/v53CuWVJ3N8/TD9U0AArMTtKdiBchRcqvrhERFONhwxfT/6GJ
TU+TKkzXUE10e3b5xPm9Y2BIH824/FkifPpXQjI2EMtL3uwWkoSjkaucOMr3Itwc
LCGuXTdL7GMT9NnVS/OLP/mS4WrBBgG4opp0vmy5+R0RAVyxMVliCSTTKX3EsqDZ
azFzW/IOTOCxrI+/65KeSRFTpSbV2/CnC9K0gHRHRyvXe38wnL8BJRKdsEbNFZ0J
qszXLNqri1tMhh0Zc0t7mKN7VWrs7xwALE0FNenENHNftGb1LvPvYB9Ef2SLSUgo
YsftTyy/jOiBdZ9a5O20v2Ebs/AawciJ89wdD3q2R005dBbJ04+ZMyONodWoFcXo
ftvDhd+z6ZY0337bmfYMLlpVRgv4MayrN2Zs78NdmN5YNuOjSaleX2Cb6UTAtoPp
WPc+hkgVa4C1/F+R3jeQdJe6LfrZnvk4Uv3f630Y7FDYTeHjH+F/Dxk8Zxchg3rj
CzFH2kW14hM2AbykgUl4cATsxbIKdiKArz43C9+a/PBMlNhNC5PflG52W2f5Xo4I
6RYMVBV7om5dXPQbP5x0jOQmQ13D6xB2ueuF/jfcFH0KbnOwps6Al5u3QvnRQPdJ
bkdiurc8s7NQvIQsJNkRSKFrUhRrcpA1it3H0KVFGaCLYhg/zd0l/qXiS5ZcnYK2
38S1WycGphYOTg+aK5/XIdzwrf3w9Kp83az9hfFxIoit5AiWtRL4yjt3CrAPEstP
0OSsV2Pl5wmiYUSMO70ruc7kupREzVU6fFwpZYZShu61O8pmYYebCIE7Zx/yL3Bh
+HNVzugQQK/0xd23IFTDN2usvzyRKRqfMuQB90jgV9E9EVS2xlDr01xQi8/F+8jl
Dm5s9OcwZV6txYZqr1Lsun4mIARxAxSusNWatGhMXQkdZBMg3pcK99e9fDWvw9Dw
WyJx8UA+W8Jl16KMivd9qiiZ83PXNLWwR7y5xMCdEtaJr9Ybhor/WuAYsf7soZqQ
ivB3zfPYEH+Ycsnn3Li+TvFXeIVB7ZisBdPzFLk6jphwEQpcO/E7SdoVandBEJuF
hBsyYVip48xF12RqXNiEPY+1Qgimzc92zhr7MxzsVWwyHI8hP7k7ADZhOzJ+U/2r
6AQiKBOHAIS9ADqdbti8gRJ04T45/CtxLI8xuYOchp33+S6Io0O/vp3YgLQlLPom
Vp8fqwJcYL71D9HLBtayg9zazv5DoVKz4FNotOpACQW8sM9YaTXI0G/whl38JYit
eGniG8eXAzc6XNMqxyqSIUluuxwV3JJBF8V92U2l1Xm0LGI0IrYYtFW+nIbOAfuD
bXuDClRHzDfsBNisop9MVbNguOkpVazuxh8zcEq+5X6MYicdG/Zn3M/I5ay0ehuG
SMNbPHniu1dy2PDdzHcjK9YsjuQmOvncSocTLBixy10SBD6eGG1oGHhUccblpwpo
7nXIDNx1UNONAy90ZXdvBwxVWfVmyvfq7nsvy1LlhfiZmTxV4tTnWtPIlKIdIKV/
A9xhPvz7giv75lV9Zrt4KvwZlTsY/BLFBZAVelXVvuakZj+M8nrsIO3PusJOPQHi
Bo8kxR5gYIZFMj7s+39iLY3KL8ee9TnBik+rFPoFRkwadcAR+V2G/OSAX/ycYnz2
TOY/MUulHk1OIn8LsY2RgJkzf8mvfqejiAPGEwBQknEO/pMRLzJYngYVEHhu2gDc
PLlWDzCgjG4J8M0Tx1C5WNULUO4otb3oTY8/1Bi8Qsfmv0rkmASdVR+rPXkVsbze
SeYVTHp6ZkVJ6tBNyYlSP0N6hIFbmvomXkLfCuIysmeJ/DdaAqJNjwRtFr4quqCt
koMoa194AkoDJTodLVLgPLsSyp2L7D0V8seXg4iCZPLmrR2CRdz+aGUxNzQ2CMVm
d+K5Duvr10IoeUmzUgCkL1JVuZX623sXOfNL0UudgGiBxHW6VCL93d0N3ErMD1y/
BfDZypSXrgH1NnmsrIt+4SbzPVH+8dH+R9Yeui+Vbx8m0e90EQXhlQl2NqgR8PC0
/8VneTR4bemldvmnlzcsnFOYWqtqZFKX1Z965v/3raagcexJbaRHL+pQO5ZKExZM
1llvxq3Oh43N6WXiwEDQchekLCCnW8IhkqYoub+lTynLp7S4TCdfM8XKlvee50FP
AMNxP6/0J9NCPFcopsb+pXMHlFibRbLZriV/X2ypEvrWpTTUdsBq9GmHhF37ppZD
tjaJuVhfEl5XDNTOh3Cv204IAkBRbqs57m+b64v4sfL/wDKooKvbQxSAWSCmpk4r
2Axvh4mZwpmane5IYydSG7tlRCXDyTq6VBMtsuid8FlV83z6oFsl7EnfsgJSc3ni
ZiS7eDusUxmSa/DamlfbxWSgkvG4afNHM2GGi24C5fvVWnCrWN9nKIyzkSTpBcp5
hJo+wIjYxGioYoZsQnLTshWodNNrDAfbSnN+5j2sGQ37sDn5YeYkSfPlLW/SzMVs
5+q2M/QI17uwqYCYs2IV/DAEQeS5Lv8BqlW2qvIHzy+gvLxV3DMLi+opAfro12rk
pAxWpx6ZfZMfp/vtGOUHcQrFY26/KlURAsWQDqSgI96lncGdZ8L3OeF2aSTC3bT8
ifntRW6KQMTkjdcp0ywXUTZGRZy9Fva5XuXLycgfGIku3UAgDCxF25rZ0Olld/DO
OgW7pXJBDeWtYpDZ8cwSZX7NDoBHT1vOBaFa4Kr9yE4POdWIpc7SxegULH2zGEOb
H4NRJmS9DasyN02/YRtDqWLR49RcPFFRo/zS0862vE3PSxL4qQGrtpN5jua31Vk2
Kw082k44d+GiWENKeVg1oZHtUNBsvcDGj+S7qcS241zgRK/NHKcMKxlLAzFc3X67
v0F3AsRAViPlGntw5ylf8xR8+La9VKxP9Ck/Ni03bLQVBBJy4tvTVJ9s69OrwCnT
dReeFGpTy/BZOkWg+2Yn7U5nCz+imooHGsaOlnUv9jdO99NpIQZFulWZ32R4ifGg
4R+V8cFqozyKaMnFe/ZIHO1RiiCWxRAVfyLQfB97R4MSRc761Ro/xedMMK6tScPn
EwafjPSbhLKM0Zlv3KGEkPXla27wPnjyuqcPaKKej0/uK2WTuky+vQwshSFWar/g
/TSCQDEBa7y8dVqKRzBl9XLj7H2RSqeZys+g3rDt21xMw5nqEXbwUgADMjZOhb3r
oIQNEL0Y0w6wjT2UJuDI0pDRsJbTWqwuGlkxRKy6zvTIclK5fKrRB9gBeICecZqQ
2T4Sd9gCQs1sugeHciOrTI5D4dYKbdPmhOZbJW/o2h9N4kuQ055VnTB2wQ1UxGzi
MKrLqS8UwsowqCWthLFxrBA8mdymnZbWA23sS46YODOx4hegFveq3P3MheHvCl/C
w9fkfkCprp/VsDBhIqY/gFiGf2ULi5qxL0dxoMn4dbzwasw9li/pymBL1k6eSAMk
xv2N7QZcBXvqGxWK9/9swF53TwHOLUf5JipcVhRmGq4pqBIEtZZYxvEpxtCJln40
ygRj81ZuiOmeX99HWlGk/KusciXkBF8cdC2oYCUsKtFZKpQrZJyYD2Icp02pnHGC
O2ubJKmxKm1sF1vhktPWkYRzeviRnsiA8jk9oOD6XQKNUL1s2a3sq8fkSAMyGvwR
RQjqhAkc5ieXpnclPIdsWRNdbN9QAGsULw6HBXxYM7X9Ri67a9KeGUsK3urc6mFW
uLne1NtVN0fDco/fUxikP75k//cT5yMwPth8nYs89GIuoy+sH9XorzaNbInNl2Gq
aYI1Gd4idaQ0sOrr0BVGZJLithDg0qWdDg7k5gFbaLjr9D6ulSQKXUInjZTNhQeG
D5RpJSMW81A9MSNCfznjpNPXprtaNfiI1zCcpB85CyyiuokpdiVtv0+bgFk0t967
rMZ5GEpVOi6jUmzdiJQweNwim4Xqb0tOJR9P44NqB3jqVuPmXORRuhe7z4IuUDqp
O/J9miaWmhrl2y8yTNSmYHMJVmJ4WhZpabJOientg9BjQ6O/HWt9/UrZxQF8SowK
BS0e8tMNEx1BCES69Te+W6vJUvbyGrl0KXciMBvTxnVM9at4bGmF9JuVuiHlT69j
MJBE70bdbr01WXltk7RzrsA5dJDmCO8iVTzRcH1iBqTbd7yD01ThloJydH4fH7rS
2udxsy3xT8xkLGV7eVElV5CUi7U7ZMV0m/h112B+E5jSYP2mekXdf2HMv5nzB1G8
0sapYkKJXmRE/tCNgTs40OxNu569YUOC/1dfNqo45N6cmh8HmpVSIxN63/4/hjn6
yb/1lxqb9SwFoz7hOzBaOQXVSjM8T4jbQaU+cOIoQr+B3+y2XI7364o/hzeeCru4
as4EUKaFtABLeD0M1CBO44YPHgO5vVU48cgx+tAup5n6GXQKREfME3NMjqATxA1f
m3pPHRFeubmK4Zm4NO6gt7m2N93rIIySUB0w0giOrVUTJKk8mp2XhyHZKRWZZX5T
8aRyIwqJTgbtOQZHQrmMprbQEBk3eEkFJF+JlKTPM7xUC/+ocQOC9w2iEmoyCXLQ
Ca2nZRB3Hnj/afNffY2hGGz+ZAKZXrdcb6+WHD4iTPUReN4xYLGSPg3ZwXs5i8hQ
okyT76RCHquHEFd0vMip4kcBvWJZ0mmHDlL6X8AjHJWqQL5JGoIDFsVZFmzX7ZSz
iF0aqdoAse97AlLYqOJjf8S+39vSkrOJ6rwh+eWFcRSBgLvZwiWK1BBqwspPBrQT
J2iE6B6OOKf3tss8UU+Tj46BpC9qUlTDqadCauw8ZNkmMmEWw9RzKCn63U/RY9Lc
lwoFIR9HLj0TFaB8SnjGgq6n6GbkcqZn4eD/Wd8dffbhf21xckEI2uRLqd6iV1hY
EUo8XFVYNihm4eeCdFTayWUr/iZHxvfZymOLd4ecT/+OkTLs22Py/ckdxI4P0Rsv
slWI8KCHdSLaqRMpt2NNWPseXfuhNCscvRmDGoI7jeMspMfrNmZaPcf3Nx1PmaSf
5iRL0vtGiCF8Bm5/MAh0T6UvwsMjqPUh/tYP9YDv/Vei4YmXAGmP2OHKnyevpaYj
o34v4oT8g+NuTGYIeYU6iuiLmSbVlKTJXsXjOWxsF4giBLgcuJsRlSGtlE1Mlk0R
JV9URwofyONpjmJURdBj30vgzE3q8M0PtfUACTGVQemB8KiXrIBQ6KoEAsby8Szl
3TtWBLIigbuYMEG5yYaGg9uorQHaFljXEuB/I4f3oY4NefBMh+eBS96j60Qt8G0Y
Jh8vkYYFm/yG3SgwXlSF/irDWyiKtoZRB4nB7yxP2Qh/zukoIFHzEsOV8/nH9X4v
SI+dMwz1iwXsdsmwov1n+6qhJ6ULnB+cD3sCDFWxRJVHjTBrvkLgYwNztT4hZcGV
1amfmCkUAKNdoiG6xHs1uuZf6ZEvgGz0CAK2nXZZA9ybg68qoSc0fP6Wzf9C5wPI
g/1JWoPCb7qcUDGVXifnrTg4mAGVNaz4Galt/dhR33doOkZyMTch6dXl7BV9Hcda
P/S5s7Y1gyWQFJEYcaRz1tjEN/SGf9yMUxeBn8H4RJ0m+SHLNkyjipFW1F0IqmcW
TxBb8qrj4RC6SSmOioXTSQvTXdsPrQXCqzKOofeWKnBb6YDJE+/uxz1s5yuGEj0w
4ZdQEVauMT6rir5WHaHSTN196J7evL+l3/Mix8bOCEIz5oZlJaL3ulRE3pJm8ICq
njdUvMYaDeBltHJa5K5aZUcoKx2XYxllO+7FnbU69Y7cq+skfigNB2ykDSdJbNIQ
LY+S8xJOc9ka7vcCGmgDmywUvV86dnO07l6OttVM1r/0gP0WSd6GxgDHYuHOfyqd
6BjCxvhRyF5amCMYoLOrxvFaO2tAQ+zfPa+yKQ1dls3mw8muGhDp4/gK7aVR9be/
IeuKOP/+0mbH8gsZRt6XRjmY2VIXj1vemz4onegvbqsphnCe70hCr29PsHQNxZtC
G3BIYtASvmsn8WRsw/butM441I3v6GGsoMZTu1fhHhRiZ1odNAIwliYDiamcjkpI
Dm80F+QfxWByeBAOjKMsbZs/fjJhUyT4h3AU1Dh2yDqTbQAuh0MlwI71AmCfz3y/
xiPIDAgEC7YVozDdD30/+HWKWKeVQ3XWMHHQ7vViZyArTB2tV1Wj5SA0UN6C8Het
IY3E1aowzhzoxOdS+x2k73LAbT/SL7f8a7pqL8pfp2B9dn2vZMNNHWb0em6WDU8b
hagYR+SykF/WaRVqiiTMDxIPcND5cgwX1Lkt6Hf4SxWyiydF/SteCI9EB2cUFIh+
fqrI08bW78Zex7Lk3rtmpMjO/y2hfYA9oyExLvUDbUgFJpfBe1N1lS5qOxiCBJEr
K2aW5bpUg1hUKQgULn3MkHuESf9RFziXWllThQ5aYrBUhg+8uf4gJhp4Vb0VFjOq
z5gC0/DsScQbX/Etxq6RtLaPyc/sUkcYIp2eSTBTO/TSeo0Unnt2SAeQpcaNIput
wuphIo4uAWnRppuMGtnJK6VogonWZWAP3KzWN1a0htFhumqq+gPrBUW9xpcLFacI
7NDyxA5g0g3Y1n42WBGnr8UHU/5IvehmuRM9Lz4l8X8dV3yHIdrJ9Zn9gUOhGulN
qL3S09IbAhWWe+biuveCxAwQ3rRkRL4+/yjZrrQAIxyy/5S+6cT0k6uknvByCNJ1
PO1qWR80ZsLCF9XDyyaYuEiJNMaJ/8a1QvDFzyuVzUWIAM95D7bUGcYb+tkPeY75
xaEU7O+VAEzYu6OJf5WokzJA3H2j/nVodPL1RWtPT6GlWm4Xlw2fosxtxF1Ln7fP
TR34BF9pEiuCSPO+c4fXkJGTW/RcRsGzJDO3z6RR2/cqvlE3j6dn7DCL0TExk0L7
XkKpElipGauWCnnOM1FGa0T1KzbQcsOwTNK3oAq2oWzYOilVVk6zLK9XMEmlMF5J
enraJ1+AKMLevyDp1LF3Lk4cwZ08T2VGaoJNJm1CX7Rj3ALj/SeLDwKMg16+4PiY
bOMui5RmBOsxFNX/DKkysEmXnAxL08bK4R6yJ77bJA9i/JTuNU5dPrJprIUG/ZR1
Bx0rf+uiCpTH7pD4w//dsfcFeVtk6MepUE7pL1GhprgLwSf8RMv6cL3SKom6+JWT
J2zTDAMPqzgiqLKOZYpF7FPMk7P/rFfyS1ZjNbHuPCYkYkXJD4kfmhccUbQ9Aa4i
p3lSjBEQIZ9DICKvm6SyOY4bAIAz+zYeNmu4hRyNrhkTK9ilTwcYWWvJFDyOekqw
zVELrQatNZJmJDvR0KGlP/0p1cf+5R9qTcl7K0cqNknjpDwlv11S+HoYHgDiMMeG
v21xhKgPqi+Q/GDeKDAxrK2e8DneFpevVSfw6aWdCkHbVFPu1OxTRq0nq6Wqk+JY
zg6rEnyxasrqpyhsgYL1zpRhMFexsSk8IIygKMHwoHQ5KDu1l3/WwicKAAlsLGuf
4dg4ufVdVPCZkbsp7R53Z4C73GQfshtjiWvp6jnat3YfCSS2W1Uuq4sN7nkVYu8n
nUsJADlnqmHzqr9XvL9A8OUlFsbgGcI2+FmQ1qU/RPabDrLgtp7m6I4Ls6SUkd7c
y3tt8Ob5qnUmefTwnaxMXUx/oglt0mZQhx9dimE2Ji8Md2WcmBO+SVVBNxWWpoCX
sxKEkhkKGYDfPP6x/0uvnWQ6lSUwloiibOvi8MZdXNPJuFDhj2R43byzmZfEyB97
FFBwRjQ396cugZ9IjdP1GGGExRg4xIsrNjPKB7LggxwYj5KiYaomih/f3XaiQYNV
jfkDkIGZHM04uytQjxmGgRmwx4uaV456GSnUXePn4CH6PBajRadhk6Be5W/PhKZG
wAzsPHE45K6m47BMlcQSFTmn1gMNt2dAEh3F18cyiYp8QU+m9pMUUN4dFDoJ6HVo
9bZaVk2zLItb2+rqmBomjVghrIy0r2GgVy06PuPFScvEC7sao7gOO1kKlaoJRHHB
g0CFzsTErHavcyKu2LbmOtggQ4+/iVHuHul6zi2wwrgEI7fcOsiLlWp0Fb89Cbys
WZKgNdnSyGeAw9tQwz683WLaB1QFL+02nPfioxHOcZ/yW7ZEiwYeVzBRxuLR1TLh
20hAon9wqtzyRdKfL+RcJyEN55jDYcgauIWFKzKeoeBA9pdTNaHCBodM3BKZldgi
rgL96S/QOBvJJdCMkP3HS8atxaomnZvnjEhjp/tpB3B5HiygdFmsSAH5aPKzin1C
hgrahy2x/Y6KT9Kpf4Yi2swd8fz6K0hz9mNQ9bHefXuuXSDnpN6BCgFiHkzFz/TR
/VagXOIRCHzqe49LH/NY1m3d/3K6UJBNuYFT3L3Oh0Xqa+KUX5XHDKhf5TBxGQLI
WypPCFDnbjH+5Ftf+vPsm1izTzBXW5ffpNKL17v+F8n7bnfH5tYN/z3986IAJi89
zF3ZTGhPE/YAzFvinKDNYbfdEwoUFNoFqFx5pmj1Iipx6eakvcgcQRjKM6fhhdBh
7IBy/AtbG2nEvSzy6aLgXxiBqErWP15lJLfwAsC+oOyjxCd98Pk+pHgQxk3dHeRX
0D6tg7HNMQPooDIGBnPgv9j3x75vCwseBNbuqKmrST9syjn7GgUItmDxerfxtwtM
KCODaZMqA0Tg4eXlr5GoPv/3MeL7h7fDAi+jmRJLgw5i2DNChrb/tW/Jazo0Bqu1
o6p3eDlN5ECWJQxdPoEqAlqbQYr3jcwFluRU48eLc9M2XE+vQEIo2SxGmq6UXSai
8sD977JVB28BkM+FeFxKxxu34ASf0aOpRWSqaH2UwvZAWW8wTp3s1482jNZG60rT
whui9ULZSNLULvzBvm8RarmhhHm4oVJxRH9MNA2G5SNDLzWQ+j1Rn+wEWPGuA1V0
ylZ9dB6Z72QLnQmdlA1VaHDGmdqExStEJ9XG2PodnyXPze+ATitvzIpSMen92cqZ
sCvZ7vKhnaPRN/GFzxeeyCJTwxNWs+Hm3ckWrc6I2KIJCTKZaxHttIXtYWrNrQcf
CFfUOLOWDN5ooCj+CPQMl+axl8BPYSx89Mu8d64aRZyJgYZodi+gxaADTcyo4WOy
wN0mHmhqziEoLod3jgN1s8n7CWkbHs7Nj23nV5HGLPGTj01FDLurBchML3tY7WWM
WiJuieuL2985qBBbBrevhOT/KUhmadq886PGa5mIKoQyWR3qscaHs4qctGOVBxpz
cIWsm83y2sUqIR2JOxsyz87QaA+nPjq1PjH7BVZSXqktKjSfpwbmqTSC4sh0/HIw
TcIEOpX08OkdiQiGDrPMysn2dXjuAmuHeVY3R/rwSnUfFofjxYyFydpxvGC8Mvq9
ZlxAXbeCTkNxqOs/41XdsP7tkHvNrG298t+AlFu7+4zDj5+t7tJCHQ704npBqk30
3YRf8OpbnpnVbe8V9nHxpnKHb/BgmqdvdXi156YVnvF3fxUeXdEviVwxO02pIffO
y/Yzpc9/jxeNkDsxzOdtUGnC3jQszxKU75DvEXqnZa7TPTrikwLL2O6BAeJgewAI
Cr6Mu5mn39/FdpPP/nHNDomXFDROKzbgYhLw4VJaj6EbTohdYVSNNho+ORe4SqlF
g2C+JKEzxgq/SfNPxVMVCC7pbS0j3z1+FPkj1OttdazQZ2BkKnkTuPyIWEvAfGoo
fZTU9keh5kUC1b4lalm49Y/hCdndW3bYVRsQy2FSzgSZrMfpykhxMxLocEYmVE8b
BHaD2AK8j4zmNm3y0ugD2X9e+5RUKwI5slZ8Tc2AA3alISgvFOv72xNgjGlOERSU
Se7wbj4PkPfGjCXXLXW89wyWOxgboOQxtyQKZoaZBtZQq/bYqV18xHmqkAqn4mzz
keKhnuq2TBDhJwxE+xi1H09fp9+eymMBgdwpIOKeahUwxoqxoWSrQKVboyHEMfAK
yvUrCOJzZ9RiFsRGY2EY4QcoDiU28DWRhPy3joNQ9e8YkeO+L6l/EzAXTYdxk/mi
mFhMCjlLn4+9icoLkZswZ5bGnI1Qn35Z45XOQiMwy0tYRlWCSyvcfS7F9Xs8S70i
/umh1oyHzcbXwnx+wXQfLXKZjZmFCnQZnAoMdnyHgagoberQqu0Z6GfvQM8a6y8u
NtjdHr9Srx6QkPi/UhH3xcSPYxK1MtR6uCAXR9WkZ/zhoVqAa1h3AUsqsZ0SGQOV
i1y7WNcG/E2HMzOQYqpiGINZACk4UCVSfhuRso7JDtt3YiYbj7FaZcg0Nfoc88Ky
rFMK1H0CfIAr1S56NoOH/XxDCvatZSM1+mSaDZWSnshAkjT06jWA9yghEyTjCWSE
+KYOYmZizl5k3g06O34KP0YSc6WCOAEV7GXpEQHr5bMYYEh/gEusNgSQnITKHCRI
kONoByW1U13KB/VdRVGdws+wb67+aojVgEXtuL2zdxszJmkHE1e/4WObV6clDDcj
0taUvXdMJeEYxp/N2m0jBcQkNr7LNCCgJA3P+/rKvHo8pim3cFW234AXJ7YwqwFU
9ETbfBIsoEPb6tuADVTQMmZBIYuEcHl6wmDGQyI4NiEMZWPn67kO/OA5VKBZQ8Ed
HO5OAfF7BX9aHqH/+JMg2biMpMawOAQiP4UnLbDk1x6scBS77nwTYICQpMMhdLNs
DiwiR9qf0MGw7GeZNnnmeHRjUTv9suapGsue8P8d592o+NbGNWa+tih5eQopFw1E
LYZiRTpPfdlQ8gKszlQ2ltHC4hVyP6DY8ucMMin8B7MrgD7DX7MoJ44MHLNCJSYd
X2bFNO2IAHZUoUx6VDhdGvwI4L+ciLEeFv8b3DuYIDLMUeQqeHdt3e1+h8rMtdnc
WAQRq3ZNW5ejyqk4Bsz6q/yfSfkpsAvVSg1A07hfi3VmX1vZ0zh8cxFpkH/zjl4U
AWpC71WyDijUjXw4X9BOXH8NIYZpoqB46XbRdurTMY4X94mabwCzoZBGV6Z6Vi4Y
Ee1oi+42YGMlcQFjlEcgdjZ5yDNwgKQ2dRRZ5Wnxh5Q+AVhlcbCI8CO8NtxSH3bp
/IeE+4awvo2ta3wU6p5LVYZfjC5vCDBnOD+zAJKX1W5Uo+f8ShMnLzPRCtEI/yYE
S8GJoEWJWAzSWIP0NVJG7tiWfOJaF4s29fTJz5bZlh1GwWeoD99GfKKgHcawWLIu
JmXXjU/7f7vs72BADGTxA+++wxnSbmhFNd9UrSHMu0Wo6gB0YkEkBYeIAuRb9SXw
ZAemHiH4MVURWyluEuGQqluH/9ZvXwnkeZSFQIX7u4sZdVAiSmcaGEeiURGW8ugN
4R1jXKUHrub+eaz+lI7UYWWvHCotXpVn9u6b6Erj5UMgbIRtPWay4RKJHIyd0sl+
1uKzZAS6hHiV+5emBPcEmlyhj8nC7c1BzI2EQXNKpyxhrn1JvulO6elfJZPKfKgG
BaTrwZMGTF5wW2Nn5lVtJcJi7qPbRIcj7ZauQKmjijnz4f5HCMdTU/jlosNVlZzR
cKRsQSolCLjhIjVl9c8kQCZyTECjNgI1A3cJer3BvwvXnBa6ptP7yG8MOVjfgHtn
h3G9w5iQaLLs4MY00ccsMhyH9DqNo4HEYASP55IZNyet0zs2ivVPIz2hUE3pj7+L
wgm/3UI0WC1D1tdARqluWRMqO1AuvODZexTNCjruQEa/zypIco3Kk1l+pBc1lyUK
j3AHa5XFGuw3V4QeEMJRUuxZoNQFEzkAlIudsUsGjVF16dbvmBQGjd0B0H3CH46F
RuAF0uuxcdXG+f9BYbdZMe0ef6xwMzyZnokdurIBiUEioeO9JdaCItGgHBRjF0Ah
iKUoxHncSvtOI/9S6g0epcw/9jdeJVdx34P9t+GTi69jPmOZ/+4EJUax378TwM2r
Dz9KZrAEGmv+l7/1ToS4++GjB9OCp6buFo4xiaH1Dwg/ccbZNGCSQd+L7JWnSvWx
9BH6y1TUuJXe+gRafo9NAuygBpaVilvETzNhKcVtBPvdQyvzIwRrf5/ezznt3Wsp
eyJAbS73nHE9xdezdYwopEIcJy/7KtCDnV/EuWgXFc2/pQM1Kn6WmkoOwH5jivDe
0eTonRhCAR0wNYA4oNITKYHR5V04zLHglS0n96FG9xYM4jjdhsvpjnUP8/ygZBav
vT2xJXvciKF6R6EJc+JeOKX0d8w4Srt98rdiKyHkzPe2LoUu9YsN9Q30H6pdQagA
M1hM9/86vKV1rKpqW+K4LEAWv54KKrD/EfO/ibf+b6zZ/NCkHQt5Z7kviRd5phIc
v+L03vBI9CB6/Rs2Sji0QyznCXl4SIBhRDGU0LZqH2jr0YKddO1YftBkDHpkJk+H
emImfwt/RB1WId+4G7PSA9kwi+/9WPNuXazA9nGqXLwQP/XvTVVY8AFQlxtZq3iB
eVOi+t9tj/fgzKqCnYR+34gLvAHmlHcXS/Gd5nzlWC0cr63hh/B2PwZYVhGJn7Y7
Z3ZkZEixRphZ/f5d6X3fdjtXSTqBMfP8UPXUbZeo+X0tQsVHukAgqJgphd4iW7mG
1/1n6Sx2O76I6hetSgYcJn5kQBj89adoxZ9QB6tx8BMle4h/EqxSQDF6gDxO1n6L
qc73zU44+mu605NkWnzGBRGUKkS97Mx49FRO/tPZscXnLnP1ec4Sf1pars+26s0t
oVQu73egl21W6G/yewrZn4DDmm1WQXOykiMtIpyqhgF5H+fcdAsjWLBJD6SvRJXa
T4CZfA5ku2GEXPZ/LEAstAgsFQlJYhFfWaAUdHAB1OFnx6u7ofk9RzSB11Df5XfS
8UM1MVEebUY7AyxyWqy5oF093mc9hhH6OuUb1XcXeT7u3rAGgA9xAYv57gxEg6YH
/c+5eAxDrVEuhgxBFmFLW51RGkDk0Q0B4IBXffUGpaeXmydDeewf/jHB++dlnaNo
F7Xe2MT20BKGca+NMQVrnU/Z9F8Z5Pf3mPj8YO4c63rqA+8kedbcWZeKXJ7qqcpM
0HTaQVwjSWgMA7PHGGYXvJD8e1YPJYqIKWSCYo6p9ltN28q+zW0qssARBF0yhM0O
Mx9nscv8RTQactfTsRNG1xy5yaekhWOQYI+9hKIzQMuB49I2nseL9anNRsMswIEq
SROf3Sc8UjLHMTh9eQBG6HUiUCXPHZiStTwe9joj5+e9E3OeJKFJHKnbdKNYKLMx
AdhCRuY/ExaJQDVE2oM7PcX38LB7d61rZEfRuhzrlh2jw6N04tGIO1S4TLimcsYt
dfOR7JHN3qSbMJGAzHR9dSBDK3hKAhjgS5OqcZgZnYRqdwl2gfbMDBpiO0J1sA3M
bmODYJ2++BBj3BD/mXg/qHwnMEhLaHZBzMbb3tN068cwp0lCeWZsZibOPa2S7Eb8
fIjb1fbzl953lVtTGrTUIXibINhtfqaBlYbTe3yh1/DSkcSTEkwvml/Y2sxg4k+n
A7CbDj7T/B4F8WNLc7KZTEb++MAKAIgH3F1+rE/dtQ1HRiV4ic/YYT2cxDMsU3d5
Etn1UQ+HGQTm6+RQdwHGuRyPBqJcvnICOiZXNW2OG5EW5DrKm2hewCK7hQPMEOZz
+vcKlDPF7vqSTkXU4aNTr03e7HLiNN9P3FED2Wae18cA6NILvwJCmGmA5w/cPb8I
fRdvok/CXXkcQl+aJZruZYjj8lMQVhcqTtXGgJrxByT4o9QCfGZ5f5AXqVPaSo1A
pWrjYMVwE2fCpU1HnYIrHsh2XFBnTrlHkeQOXyPoBR1aymbCpBSTkIlbJ7HLMYCv
i9cbfZbddQ5GBcJuGUobOuHILLHjxw2WCvtX0KYrKMxUYcN+YHB0EwZN2fNZQfCI
I8gr7hwnTfqk+aP5Wn7G1siQQwdVp22EorkE7ys+TeMAuanyFBJwG37j4mTBt7OB
L5K6xJh5yLPcLUWuVimQfnuXaMdzPfYDoBL4S9QKrSuR2HJ4zp7pRdkkDDu+Yzvs
soCeKfWvYWXNiur3J80gTROkidkdJbIH6YH15ARJul3I6/e80DOV4TiHMdBTQyCO
ghZSAiAujGKFXzF5G9fuc20STbzxnsYLJ/+vAUYDrtr4U37xnORss/7sVm4vFiFp
yIaiMUZFFFB9n9AYME1xp4cHig9QDfy+8AF9IpmMQYLlUtKjVezCumY3S7tKB9PR
s28ZAE21iOvdLHIDsdwKiCGpHruQqYUOS8WCbqfbIBU/czuV3VjHfE4fBPxbvPql
QuK5its2k+L8mi9hrFEWxfhaSpgGC5GqCDnPV9uy/Hu0YLxP433bCEQOcf4WbhAb
n37z3pkcyabvDkMMiaVMdZj22JvDuGXeoNyuT86ww1HqJkih/LNowG3TIsPOY67C
QwCnox0+vEJIAwEW6Ei/YTFWehWn5RCXoGMrWN5gmgIu32xzqvbERXUiO7ODDy1b
v+34TSN9G3kr6lWW+Apj7fTkiu2XXbtrunba/1m3B4OrvLnjPKdMikc7yTvRIxEj
/x1kNiO1OpEmnXTi0ii2GRLBxMCEqBWQ7/M5fkIMve9pV5uXMF6noOkM7q8yDFQJ
68xalttF3H0RUH+vFOE3zvCZbfkturzIA8O2QHxTq1v2WuE76R5ikE7pFJV+vZ6p
WE631egFADKGCKxg9qFLDPgiFjQ4ALMnOTprFIlG1410QHXEvoOhfSuVREgLwwUv
SoT9rxfE4CZV5/SQjon80YK986kkPqirsa6tJpcxFG8EvDwbsB/8asJc0PF61cK+
Xf99+c5dV9+YxFj3tlTFVSr5WhGcR5g84PHztGKfjN34ytPs0KUid9BAKVzBhhX9
6gW5wpHcmqwuzkhuyB4R6nYjFlEppKkDq8TYzPjsSHv0q6mkXCh3NtRr7BQ4XTZY
rlhEWEBjkygBtKN0hwKfhepeOF6ULjr8jA2YX45t5C3gna8KWCuO2je7eQpTtQGU
4J7CXwdDhOOo/jIrpvThEiYwAl50wFCQbo0I1qHy6oDFrfKjyYX0mUG/HVEJmnBD
bxY/uUAzfR8QXTUzan6JGWwnyKK8QRwSfnKIoNAOmtK6IBx8IhcfhqNg0YzIeZmt
6jJZkCHH12Q6R4aNEOYkM76eOxahqjFMxZyUDXQv5fPymwyyeAdIy07Ex7sLCXQ/
fs/gbV57zXnY3jYgoZBVg0kqOPgYNMf5Ox3Jg3njwcfXUfpKvl/otaiHO5iqB4JW
f2gZwQ+3MuhQ/uczQNkwMYgxvG6eZJVb/pqiQNePvypoQv9cMPYPIVKoVLoW6h3I
MI1M8WWJ9Mf6u0mutSfyb5SWBuwOO7Rlnpr5/XYQiKphzeWgarxQLE4xpmQvxLve
LaHjG7y8+tUKdu16MhxRzqLlbh3FvlXAF1//s6kvnpwBnDDQdd6CcnRkyAuMKaqa
2VAaR8G+Mm7RIFuhZoDh3clyuA8NcWPS4TFzkca8o37BzZf1q3G/K2QyJj1WMqLP
BvqZtjCwxgYv3Bw2TbJO7xlvreTvbSmeJTcBUWE/SNHeqdhDNmkohSucQnQlmEi/
cOWGxA4LAqoQ0YbfmJotRBXM+kLAoKqy+pLP15YMv+rH62ilV4T/r3bOWbg9oEr+
Kn2NaERnVjgZ66udsRhiRSSFJKxSGhYJFrSlrvvOhikP7C7bIu/f6SPHpvbRCC+z
1/KQIiPiEBAUc9I/FI494YxoaWyzKLX+4cVvpf2dJAWvZUljxUQmOFQe0ujA+tFH
C2HwTqSmueON8rSfLKcpXYevDvtWLZTKOGWMtfnkSu9sSgF+Foj6uWVcbdCA7PFt
r9aH64fh+nX8uRTqH9unlV7hqlkik93mJO/l+L5DSNrvryZ8Cy5nzaXzlyb+f28m
ihN2tJdHisATMynhUbyLnmG3PW3KmKMUBYXPdI8VOoaoebe13Pt5El/osQ/UwKri
zH0Xz30XolXnNJJX4TJGTV5eqWhmXTeoHH0jJdW9oLEiekJw/SPdvMPKSXNMGwzP
Hmlqzg8DCAqliZZw39pE6MYwARu987oewUlZ0jtIZlKDbA2bTzBJzphCt3zVTzqy
BqUm9W6+XJEiVPk6UEeP7lFENwnDBEQLVBL4tijq+kMyA/VzYcEACK/j83VuTeRF
hJFanqNEUAeiZLrubXa6ZpJFdK9pNUcnMqAPRUo1dIC+PP7wbXYh7/gl7y2OoZ/W
33+1/hd3qVyOx5CLzF55CoIq9pAApI74YiUrF+gRK/P8KPdoilB2JMzHuxp5e6ig
8891RZ3kiGlyghV2MHZqd3R3UWufrNRmqNdkk71M9fPkkGcr6OgoVQ4z1QhVZZq8
Afsn55jwDLoSYj/uhLGe1QGa2lccIx2p+/ZP9COHB5oZ8VOSK9NJgpQnYg0ZqZc2
GDWl4prSbifyYs/TI7XKBBjmMEwNwyKbcS2XNdkFLu8KxHcvFjp8SqMPbPUHH3uQ
p2qDgcuRwKTskyAK17uSs6lEVrCUYLd7dEhjUpN2dW/dHdOBVns/J/SiOKqaLEJS
2Io7Lp010a5oYqDa7eIjLSq4b1lvz0IH1aq6hbmWUQY6YaRALHlHkpFgGFh+BneQ
oXYhWed58SNXVdgOjVl7b37U8KK6wcryXfzYrBj8IXnHzN3TzbkFzzfPwnryzdtL
eXWbFL21R5kdQCTkK7gmiFA40nnyiqcfQ+phM903KimZOSpQwi0pvdEotACU2RBr
Aza+irG8f+SOvmedsTaxarFFcfu3TbFkgQ+5qlgutFHBEXl5aO5Alf4I5Kx0N+WM
FkGrGXLWq5u8k3xnG9CazML8TFXSAwmorwO59/duLCWRjby1o2yPh9GHAhUZFBIo
EfMnt16JqdERHI9q+7hRjCzX1GMo31U6MFzpnXab4XWEhD5kGL2Nnyr7XfeL10nO
SPVd2MJa/lbWkvZD1m9qfCsWeM3V4Q4+2RPzjLFtn+gbr8t5oYCCDN2ispOJUnSa
9O76YnMMcSPcE/EtF8xEpic5WkEviChAqMeHfXVc8lk4ES8F6JnNXCRyquk5iEMs
HVeOE2HjBLtPhw5vsaFIksj/bYX53T5bUGG+cQ4hLbk1L2AMXSsqU/0qb7Y34tq9
K/Ie/hpBDGhn9oLzeF30FiT3YTmTSHi3nPMkYUr9NPsiKSXpyMRIzdUhV5qGyqf8
GfcbJVlZSo1Svh+xN7H3OOv5oJLrtdcYPb5DHBXhC/fh/8ZloWX4HIe13bxiLuHz
r/i8hQd+Afw8L/PJVL7k3ZY7eLjLiGinB9XUadSX06PGYUsovQd6O4xSJJSgLx85
QyAKNg2YFyV+Fbzv1zB1cv/k4Wgu9D2EHS+JG2+gaRiAYMMmyfkQ88FeN/vsWRMk
Tg6HokL0Xy2VgFLGkdqmUgsOeLSXFl8BbeKmQ2BfFSEB5qwt119aO762BjPzYZN5
4dEqglgPbYeL+9BYqt9PlsbKXc+HOOJX3ZgWTcJMeBJEvpmkYySV8ILFT6WY3xxu
a/Kjm4kMt/ARWKJgU781SrProE+wA/2rxY/EHLRFdCVGnt+8qxwtKT77ntnEuxR9
dz1tC0uK61uMi0E2NT+sTGp3TCIfTTX2IETbImpLK/40ofkwsCTuZsFUEmAhKDs4
f3UJ334VsqxDm116jDHMVK0WWebuaJXQzTVS6oxU4YTsWV9OQ2jD5mzhBJxEKQ4O
BRr6T8n7BMjj+PtFjE4XAuBBchzs86jyDnt+on4rb68vVm4TcWeLGirhsMQIW15W
G/jHQZ2d4dq4tGVaXJ3RRazY593A29bZccFEpOyzsIIYBoN2RGYBc2MuSQjdTdMo
UGQ1YQe01V0ALfvw6hPgVHsLlevNpbRcDCI8zaA6m0WBx5SSfR1Ll5tEho+Yfyww
jE9ISDngrXQbDjVX+3k+k/JurnTGDEOBfktgB8XaEeRp0MEcY2G4G2i1a2H6udlN
lThaXq8BsAhf6hbP4n92Bbbb2ugcSmZC7l0dGoisEu6DyY4nFHpQ38dZPXSzroek
Z3Kyy7IY0B7XzsPHDr7uq6+VqxfiVgBL3BbIU2UxbJfJdffO5iwq1VD36mp9IZZs
xQnNHl8hM6Z8yFi9JbF8Ma7XYwuHtlwpDn8CX/mG1nnNdpcfEhVk1OWRwgb4zhRD
xcn4a+FsrDtXwWdMtRb/xYVe2DhAsGoeK48+a/53CK3PYIthmKQTwH+/PQskOfM5
ZB5BtSGuO556PrlYWBK7UXDxm/ZtDrxvnTwe8kDKC+hmOh+5NVROqFLIY2z3e5h7
ZK7Cft/psiAlrqQXQSONX4VTPqsijfGMw5LV8W+3kbxbHOErVsHjrMkO4NwXQ6F+
ULXMkkbxy3jzGKef7nLCA9CF9jS7MsGVCuuxkCYlK9hc+fwArrevyJCHX7Qe+uOy
GdQGkRBT9Y22D2Ysq8+uLBPGhyOiJ2ofmrxyhaTzF7s9oFFuokQR4FPuRb/665gL
zp0Gwow5JeZVu1Nu7TpVxwDuR+OnH6+uY4+FTYNqP9f1iJJCbGWaRzXLswufpiCC
xq1t/xy8UkSl/O0w86Hh9TLSpSsvRd54LWcOHVTEnuCk9KFKTlQt4GnipKxFNZyr
u3c2/+iKw+DBVAFoOw4CxuHJtLnUPQ0x6oq4hAmT6Sozk+n57QIRJ+EHe4V2I0cn
rDrX/d1HEO9kT48cqS0nv79I6Pla1H4qUL3Q85I+CyCwDFVhtPjNYCfcvxcIZXTS
o049Nt0GicyQjgKhR1m4zHbLaQ6Uzbs5/69ZMxrkyrM+7ilI+7S62ya6WOF2oXE0
0NzOx/NlTSj38cJnkg6RswJk4zwbU7eo//lW0RHX9wKosRFjLxrtYEFyKIxPqXPD
cSahrI/vnt2S8pEORJGOr0R5oVFIm4ddYMThOoOXxgLjuIU2WRg8gibVBMfelmGu
iKAHbjxzjD+Q1jb70ovIrqMxrcekOfWclfNLPm0UjpJyRZMm4Mc1NT5Cq54OxHMv
qEtaG8ghBhFqFIa4lpA7lNFnXFgBItlPrkPfXihXGg93pZgQdj9qMvdSRM3AvwEN
+k9X9v1B0Q8ImH+gwM5CJtuYSLtrEVTgPgNTJmWmTFTuuQBt0XTXY8HX/XFZpRRU
jjo3ViIRv/1X4oYQbIvSsG6Xaut7vL4I3gLWmAUWeAfnyn6Yzqj3MspfxJ11QwS+
2sGSTd23olioOhkUoxfGAEa9s1kH8p86b1KNZ1umB/tFHtY+yAgBOSP0J0JAEQ8R
lV33TRY+dG2AlGuCqvGClqenBLrvn0w1y25jtApHAPbm2Dm3TiYNS4AKrVK5y37x
xYM8ctGOxvP1idqlihGBSO9W6GAdCIc0GMWPSax0MG/92iEKtfI/oNx+yK6PqJh8
tbgXQFSp7paw/DQ8PlE8o63S5kx6pD1zela0VKIU/NHI2Usi8aW8ae2y5a2WhtP/
3d/OW0BcJP2n4LXGKt6NIvUxUS2I5cbQD/OJYr8nngSHQm0ZCCcAvqYXPDXlh/s2
H3Sr5ipCG/cStZ/2g+ATAT+vPgoM9eRdjwcb7tuj7CCcOqzB+OOh8rtuOHdKm8p1
52De2Yh/WSx85bunwszTfPjEqOMeZsZZAdpCjKCp4pBIz1BAKLGj9zjxhy3S3RwO
cReT0TK01mChWwjvGD4wgyVyb8hP/0sSv6A3Xgr0/HYtFUhjBa6reu4/QSlpnR2T
wUT34QqYaZyJKEwsX8KYHkslaHOV3MvGUFbWJfxPC+FnvB6X5X2BphE33HI35+HE
vfdakzjeQfDJZ0eBXojWd7HnLMhqV0dExiXkuAypHbd+0LIXCc8/ZZUoHz8XlvOU
jEO5J9In/zdqbg4NVcD/C8o5Fd8UafxaEdJBrnZ1snZhLcQnCnyTE+7oK5FVrDpb
ENMcMH8VZXFnzgP29pRMNSwVv4dmznYok1RibWD+goonTXWX0aBeUZU3YRAZvKNM
kJ0rcRw5rLe9OBhaD8ZHmn2PfsMkTfYzyjOTmR1KTMQHBxxh2XHyYPdDT0ULniYV
WjHCAGTfqUl4CLDmadfWmGhzDvqyr/FEYPWcsXnYPOJzWBmED6/nYWHSH8YpDLAP
BCU5v/7y9JUMkXK7BlNJzJJ7XDcztGHJGtXNYV18bKVYePsprlQU6M8KjCP8i5mc
eIMe3uQcRolBVqkPFcATErhhnUnVu69648lrxCLABkqoKSB2Ob49EcULKlWwX47N
oi4BGNTDLBmpGT5susn9TMsMJjAto5zgygwQzOSV9SFk7N8j1CV76Te0hKUOb75w
392uL77jrjzZo3/KgLUIvMAhIUeeFF9UUd8FrgTNosiq46f8KQH7WLXfKqx6NJbC
xAVZDzUwzyPosVDfxyJCvH4kYvGSYp6+6GzgLEy6ew/LzikUT+tsj1OYp6ikR72w
gEY/auVcsH8x0/anhiR9WUH3tHzWZnkmCnFkn7FfWyjMHZOwmC1PKU2qzkFdAMRg
yDGACnSgQmRMFPtFGF5q/bt1JU91fwd8KDCPLixRW2KXU5tvX/rbUZsK8+GU9VMz
HduUm8RUADAFElTcZ3TtIgoGqfM6SptKndNw4Z92Qg50cAcd9c/nQsN9lit/2Lfl
tR2SeM7ezUclH8CJhMARttZu0Kh4wOVqQz0GPOTZe8ZvY0Vz4m6wUuZAeypnZXxu
/MgHMGwqmtDjREbwOYvuJx6gyiO/Q/bqtEwwwdjNEeCHT5U3sNYNJs1h2252fvYu
Wfwf3K2dY0YWp4gnnKiLGuVU/xYFDmnEiqBCWwtQEcCGjAVJlW4Tk1AXeiSmW2q8
wpTUFiRps9XCQIm3N1EscEnPqeecaukYWT8l4c23JddbsSP2MWCL80vgLdka0+kt
WRFhOIkj4hVBFpATQX2QZUbYBLH/U1m7ilf4e62TYT/DITQrBrmqjgWahlHKtPer
UhpwqlzgW0v0YRodhylZxsBOrNlaZdSuhP2OAob+jSsOfbfldZpS0+YK85iunvTf
+1TQUgIMjmc6jL6Mc9YTWf5uoXrLYKUHkL67GaFXS2kD/yghzKArWgtjcZEJAD5O
05+oV42mITOZqnYt2Vt/YOX3MN5oQMCtMa5xZ3MJk1ahDPBMSY8uXVvkm4wryk7M
6fOwX2ysRxHEb2/Ep87QZG4CHXNACRQTf15eOHTsw9F3DaOl+Vne77Jw8GgkngSQ
GM/iCr4nCttHhadO8eOe3ZuU5jN4OQXPJepurT+VGPnvPi6PmuY8R4G+UtYvGKn/
nuHj8mTHnW2V8l7j43h5A5lDZVXGSp2+TwIsEBRAgPXmzIxPyfVtMDtCQH/uUXt+
Ki1cN9ZDFsy4Ao+XWJfSVTOO/dD1vdwKUXalL4Ev64XQMev5H6uFqW03mdX35A9b
gAvfUzqfhEE6X2v8qUChNIt3kgftRgegYLYfQQVbAs9D6S48Jz5xgMM4obRgNx7T
q+5Lz0i5ZSIMUVwpVQ/aEABW0Y5bESZ63oTWBGZGfkNS33miyoVtvfks8pnWCJOJ
0ia2p31bj5qMHsbcvcXteRMHSiaO3iq0bymE/x6TYGzfjG8+Vz1NH+A0HmlCXMp4
eDelBFdmegUC7iCZZ38Iaz+XuIbStJ3eHeMSdCau65rdN/S1rwdiRdgiBJl9HNcD
MZm0P7G9Hc23PwU3YAHm53Z8WKSv+JR08+6rIPCjGjP1ubxUzf0YD6vjWY0zBGGn
Y7SpzigSFhD5GmiI5eX6WEVV1mKD6aWESXL7Wux3oW5rnGitWeT7l8GonkX1I0ty
Dc/BcPUBGxE+QjgmBFRjBF31DYjgeiqqDNyvC9lZcYa1rxyI0vDQQAMhHr/hbM14
ATHftW+WqA38cWp9poQppD71wm6AJEYiB1oEh7QzHdpVfHBdMrzBEytpz0s/MR6u
l7P6yb4EKXfwGQWtSUJU+xYHhDK7n0FH590XUPR6A2civerEUKaDbnRpKm08DjTr
pID+CQA75KHOuFR6GWGgGbDqX2GJeuXLZ4XLpvjeXoplO3iUFoqu+YaAZq0AvM5U
XWlp29bry1VDRBi/70gATrF+lVKQQkdj33SRXRGfwYBCoHLzevLa1S9g1+9lLi0N
OuM/60e/tlMHUhD89O1eL8c38QfjUPThBPHdX6eaza/fcRWZx3tTXHjzFDMJUqhr
KsrBNdHOvAykvDdXi2pURTnnxQ2SF6p1v0c50/nAxs2BGHHelshAIIA+6etnVuGe
6LqIttvBO2B1xZWPWb9nbJXnO7ViQOKE/9/5zHgf/XR+0AWFoOpWTcK8vPPsPH7L
dSxbhgQxnF6CqrDYY/2Bbv/3bFgTmpJS95w/1y2nWJhQ+XXwjJSTMpwOZA6DZpPl
0Fniz3dF7enO7kpv4KHA8YaJ1p3a7l6hz407JIFkGMwbwr3LZ6gU4BBbOtFHGQTs
JfjJUBtMtpxJmhg2oiRZxmL21NIOwIAIvPleY+8V1n5mC6pp1arJ9oyIGVmjDs5M
qzcFQvsR5xlzlVbIW9k9na9f3KiPiFDPd9Re1/CyJwkOdt5yojF3nG+JstBMswF5
AfTWZA44t3kldH0t9t9h9ZlA7DBDI9i5ullFiw2Nfi/nJASCRZ1+g/kUvrXVNBiH
SUCX9cYyCh5Yz7j90/Fdh8/s3jQRF0iIL5FbHq6pU7fzbohe0C0zF4FmrT3DB4pk
ZHMSxxyL9OGppAGwDYMBEtFjKy8w4zVoJH7Q922O71G/i66XJnse6BwnX30GTTLd
y8lMUfHlnGgToHOgHcn387YUGa3YBa4CiQ13z3mpNdy1991a2epE6oVjpKdZFkfd
yz8nZ2eFm9vATVROY51XhfacB0vst06zwaSB7B2/ugaIsYsMcAoAoP8X++oHdCgC
YySAkPS6Rt0YRD+5eBAJb14K3qOipOfiu9XkUdHKiqwDcibqDI5SwBFAzgGa42oD
yA5cIVUUMDoxhe6uBKuwe96jVV2PoKI1C1HtkxKz3iFyXhgJ7xGPMwI5DN5Um/IV
iuajazcwCYgSHtnrxkzax9Db7ihZt3MJjxMWEOL1SpnS0uSA/yxClNa7Rii5mAph
Zidrlz+8+oQZzXTZ6PJjqiA7+AnAMCoM5JkTQcbwLls25C5OR9Tz80+wHu25XuPw
EtjLuVdsG4D+1ibXgKddtAoNzgMOf4c8+SrXUljlm9YcqK3jTuvmuBRdt++p5bi4
LEk6VOz3NNQHIAf+wfTUU3YVz9pMwgm4ZmMZVE1Vb8arRxKs1147/qbqEfHW1VT6
qrdN3PXblVVoDdBRZsr1opY4W/8+3GKqY9sGJSKWpw9zAs4SFB3NdzSAW6maPww9
lhgyaSbJlQ8k0HiTv0WbuBuzH59Byl2UagRP3ok0eqbFiEcxiPKYvp4ByFuzWpig
9aJt610oWPoOEfBErkBG8fm4jIkg6MM/aOdHQcTkFIoVlI1a58DV5wVg2CTIhAge
hotKqOf5VwW5ikr+RerJ1lCzPBv+BmDxKo+pyy3k+Hb8+UVvCjVqSu/wMgrT/FSt
oCp24A1uZcNetteiUpwJnqLg40NlxpkKrjswaiLFQaN8fxv8IGhJpRfu0YhWMIFB
c1CW9WAM2PCFcb2qe55jRZEv4Wc+WO+mInKlVYVCDnfgKbUtTtaLP8IeBV1sEFTC
srspz47R3uzw4Bi2r9cJeE+0foavH9DlS6WR9Kb/OmLHtEtW6gnpSMPIgNL3EE/z
6jts3hgy4tIQ042ozKO/nXuUM7/G7fIWQRNKTd5ITfQ9qWcgQFrurzaCD07GkltK
RveV43DdTlH9hQ0f3NMuSrDycVjSISfPdur3Gk6ooZ5duM05wg9OdCI6LVmZ1aji
XwXs+kUDpXozT80U87BLJaeyUXJymqmmROL1lVhjqbyZl4hMMMFzeKizTxZxitfc
rUAt7UD0l6Q0SmqFoAgHFN5b+euZbwtds4LOZ14Ulbc7gF7N+aJS2ouiu7BVpDif
DRoYA1UdU9ReqXnQOTNLoW75aoXluDGCW4rn8m7H9jlbts+JqjcBeWzjZ8RknJrA
t3QQ7uhJg+WE87RvTqUJwI+m/ouXoeLANEDGzP9Y9J16gGFWESTBPbjnzTeMa+D3
jqibceys6dStT4MUWNDYKI1NzwI9veXnCjypcjL2L2rssXBcGPRYtHphEWQvUUet
H1yPZ0RyiuKQcdLLWxzzSPgE9PXJMUR23Ri/3sesKtchFk/c0JJu5Bv+VfnWZvbE
x7y8BKAAPTNwJaeAw7sO2fmeCA+/xfZkPoDcPhNAycgqTTG6ZqH528bnqdwHQDkC
xgvhLzYZ40vP24HhW2+JPFr+iksY3+aKUTQMSVmbDd+2FugqNDajTZTYWA8dQIpy
+g41PdpTGKmmfRiuRGt+S52otmtp3qghlOnLCNYFTfNA02V278ZeTxUDuoEiOMgj
cS5hGKhn5fwerel1GBkyjnC7Z1UBSsKBvZ/NgNWGJbXCsFQSRjGulInBtVZcTZBq
vBiM7KrF4Y9sel3cbKbLKYiDgUke/a7X1h3HNlytePZFJIsrMgyHikKSxSRds3sG
8P3h/cKrlz5VF+/PwEnVnDVKKSCrJTKCk7TGw9bWcSCf84J66yB+eT/beIEBxS63
q9VEzSOuK6fHUCVIe4Xyr8gVW99afCjZuJbCyR/2jX0enf0/NfT2Sah3sr55zfrh
Vu1shrrdLYZqgrW96yyJ5BPvkp5TtvyOR6IoFXvVI40EbRQjTTuIftvwf8ZjV48N
jyqRDyGhEb5j0EnYnc3xl1PqNiHZBr321CFyLOX9d/EB1uhDTnNb0B1yepOShHnc
+GSovose2S14nNe+j2RRwWstbi++y4Tnjm2KabRxbDU58vEur8OmqKb6/b/X6ona
uLWMIIFcV9OJFYnel17J7GQYGbV2f+V04eJH8TBiSb7TtTqqopgb3etP/pUU6S7C
wWYHRSxl9busd+ngGZI4qTsEKig3tuKkFDa9l9dGG5NZq170T3CkqGgwtqkxVirV
zcRsHZhDzDql1jaKW1Wyo5V5dMOqMBu4+PE1+hcX43L2itzdoxAw9g+8zitM1vot
cMRNDHMWdMC5uBuRckFA6uPYZqfzA0DFA9SuidyCM+2V5CbfLtVcexji56KHd1h4
YfkKhT3qiNfDTiWHNfEiFi5fx4e2qJmHGXlt+961tP7AtorrlgtP/oYyTA/uNQ6j
L3c5WRnOX6reJLZOhJhUhbvoWKAwyILIMsSEhD2adPexmuqSd4kkYjBrV985y/NO
YeA35M1Pwz1TYDref45TP4qTwl53SGTPwjA0ApCvNgU6ZOFjeF4ewfU8VQkmy0AA
fWkYzg4GxwjuQ+3FZe0M568/x3XhTsNeT+AOslSoZJLddkvX7/jqhezIZe6jtDGT
u5VZ5ynwRr9ZAldnmhB3dDv1F4JYkyP/IOfY3x9/yV8rGRGhgPtiZBrV7b2i6KqU
aB2Fn09jZzJOY3eEkixXGijlDy0+0DwL26eYWXj+xPixiOv2OXFRsViGFFJG5tZq
uZ49XyrZuLyHMHRzkHf4nWRdvn6jTaCJQFvzUA0GF9a+Z1JgyXqkzbD98cPd1kpn
ZmvT8T+zSaTdMzN8XACVfbZshAzUqI7/F/OkEswTiMY0sWWYLGcJCo7RsQSgYEDc
rdx8wpwQiMak04UzQJebdn+1CkZxY947kh1KEQrjyH3TQ9OgIqLxbULYLLzvODkx
PUi/6mN/RadWmAJU6HxEEhn8OY74RETUMY63SX+iD1h0YARfylvkmW6ZDhyj84xQ
1HGZU64LqHOJvLgSncCoc+w5FY/1QbKaciLkfFcq7cBqrJszPKct/tv/WAZHQNMO
3othyJWwNlT/+pv3Iw05NRmzGDZrzQ3+RTTT3WKCk1spkcU3WPQZ6/jZvGgWqUai
sonqvoHmsqo7pwyhxzirr+g8ufvJ8baloNCn0LywQzG+UC+puua9pQ100aAWBHgd
TCbk2aB88pdBQAuL110iR3vh7GZKizO2Xb8/OwSPoeMBKNRma4cE/TA3oTVSGkbi
a7Qt0/jCAqj62gpvDj3Cricn9inKPxO74uuzWYLHKBhf2AmQwNIy0z7/DIOv+khy
pWpxH+LR4xtQjj0YYb1KsOxQ1tUu3Pldm7W/D2NUoYy79fMK8ohouF8TdNsB/KTE
s6i9ntdKhCfIHexkdC5w09V+pd7+9f75nZwHDWTpWJMUgSCvBdv8wBymsnm2ywRt
FflfpMMCExsR058VtputL66R9nMogPbMCVCKQWq5BU5GRF9+G4vux5Hc2BrOqX1A
Pk9MGfudRezVmbt3unCJUUOoq84tW4/d2p825zaUUVN2oHVq77JUKBBDzoc0MKOd
S3+7Wh5kuB5BjgfCvxoQ8rt7H4zDxjsmtVShQ5jmCp/nZnyeGfwv2D+6vcFMW7iW
g+E0uuSRUUKRwMopZ22YniJaDGsAsMg0Gd9JC6a+nKP2MzznE0UvHz5GPh7pydkt
tYtFLl1rQqVDBaLkql0BFZzGK6aB7kHxLKCP/U2ZXlkcuv2XGGlyyDGwQW5uFQ/y
NdtB13WtzwO/L5ijq+7RoaRDAc6GHkklOqOGTVjQPn72sHObbgMA3reJMNf/VS9q
axhaGk4NiZ1C0OtkwriqbyaPSamHo6rhpeZCT478g/ZDmgzeI6VQszAqcZkyVadJ
sCQHj0eJA53BA6LTCbEsBuxjylDOb/agT/la4jYxkQQ2jtSWn0SqmLAaWDf5OzeE
lLIdzhlorRAgVYdGov2cPDJRXlZy+0ACMoFi/oU825hOEU6/KJzfTK6elH41F9Ek
+PRHCts859DyZmj9nqn7SoOSzipMQRl3wa2J72s1bMkniz4q0cHOicof/wLWG88p
znMUUUFDZ10qkAG+KQ3ZFWyjdKik7dHaPLsFwInAXOVVtZNBQmGk2kDLzwX9/CMb
/0yf0L5nkN4sEwHZr0+PFPTJL+hZ0liAxEkFRw11VQtlYmq3jmRoNnSJwdsYB6O5
eJDwPkcS4CvUXZ7Q1v8moK2297TWuhrJu3CoboWUIZfzdX1wG+Ri3mbLE0BBCK+3
i5lJGL9QRlOs1FMH39Ox5ODzJss7PUIM+mCoGnGNExPZl7br/JnC5BDvTHfxSQ1z
7Wvy8SCYXc/fZhIfm1SLPeHKO3ZFsjUe2FaiCuVcULHEhehd1oaHkjE/paT468B6
FU/z7aQO7E3BxHVxcp41JckW3iMyqddn6C5+4z0zAp0Fl1m9fRGvQbDEXlaTs+XG
2MR7VYFqZ7C6iUQ6rLZWpU6SO2HH2AisTIS7z+Ds8Y8FC5KYV7Uv0RcZla2xaizi
72i1qOP8VTxWJmaXP9KeVUVorlxfPmEirY3lRL+sIOC/iUymV8j3qW7S0EE1fGss
aRt10hwnSJ6M0X2TPPcvBU2U6ghbYbxv/sZkNakN1Q7B1c1LKM2i0s20xASLXpeb
ys7gSuC+KLiOXLNGhbpbWIlvJiDAqikEmUG1JLvi4woSQqWgMaykYrGzV6nSY1Ae
BWKatEX+2nyOaCa5WioSkqa5yygl65MwjYCoQAoZL0B/pnQj64TvH7Fm31vNPOek
QoSq2c2uCCREGFSWLd5h+OYsA7xKzxglriE+WqyS3dOYYhiwznNB7+r/Fek8Ve/r
/IT0Zxg82wMrRuB7j4AFTmhGIdRjlMczXtgbWCnVB/ZWlJP21g1sw2K8+M00zQ16
crXQBjKj0hVN2NB9WpXhLQA53Tiy7qRdztQl1euIRAN6qRGDfAqRVQxomsG0I5Bn
e1b3WhqAV5FEa7XpqeDQzJOlCpbhc9pum9kscTcKJh7kvvbS4DietL2jk2YYdzPQ
3nsZ0yMoD9LSHxJT/u9UbhZEYvYsDH+J09V2acbTHdys8CXBeqx9IjHAmrlCbFBK
00Afao5o3s6+FC2UU9WswYQZlR4cmniu45+94Ia6MeTu2q06Ono6Uf/tD7AJxEeQ
MxlouMjd5X3UAoNq5Gv3Qg9dduB8NJ5w4p/Xv85a6VOwB309qL288HVnytL77T1a
Ox8VbWlZfj1HW9Qx8WXL5yUxFHivtqykhhuvmdCF7lnhOTI35VIlXMro07KB8xfC
GKavqEY8XfiHneoDUVFejProh2qSy3VotJ+Vsit2T976QqtD9d2n2rKo10ubMd2E
6TMpSuFD1AxKtPPRU/rxudSHckWBuPIFh3zYdv7457YP+lWIIaBn6I9Uzuja6XHu
ODk2JlQoZyAxWW4Kq0tOiZGZG9UqUcO1zYLr71YyEhM4v7jXvvWiX1gvp1M0xa0Z
BGl/lq7aYP1lIcKO0wh3p28/Oti/C0+ofZTIzT7bc/9bd7eS2VSpoQiBp0YKNA1e
vSP1ZMVTZO26NqOBSx+yhrvTOCxAchXxXkfy138CVCC1W5tDe0uDWnYWCz68kcnh
2ZelHZpMGGPyJE71gDtn1Uq8fAUlx/7C0LecMwyC3cX8WSl6q9GLN6ft2/SWq+dR
SmfqMIjRT0kgosI3xlWMVIrlcKKyHvjs+PXb1KRzazhjznZlU0ict5YAwrHTVAkR
eba9DmhCd3QK6qD0x4vZRHQs0/Jho3ZMbbDIUzKGIt7BuPSVcP6G3DjDkqO5OME5
Abgi1A6WUZngQg0cbMc84JaCx8KgELwELW3Xkg186OlLcfD3mhWakJxX6ZaENObe
8zTWFcsagwjfyIgAn4gTtAH6hp2yxgg0S23eASb/dAKamiB8dMRNPxZhy5KRFRfl
k75G3XOpKa0f4L8CdOwWrgy7/HXkp4DjFZrjTHf78WiITa9jWXvpYyEyMQhpmCTH
DLaVsnmpBfPubBMJfmBbUKSVKQziz74rSzSVuF2iP/ekHYYyLZKZ0CM6Qt0DRCrp
VDSSH3kO4uqKgDG5hTwJ6t85gjMR3Cj9kZg4m5TQtRWJADMa/UH/UmgYrBspgMUF
Oj/wxjLQUehjGn3W1E/82azlpkIxxV8qgjHie0fUL461bwBs+q1sDFtnASolSK9i
kzqTrjVwOSQyonw5/MZtkzQGQgKNkhA2Xr9WzNfWjpe19dsn2zuSi2g4T6Zbco2j
WxlRe/LIaByj8D+hIHN4s8OGbo0xuXDrQ50srf8NUP9SC0168VuuyNvrUlew89i1
O4UFQgaA0bXAbELMGaW/RtNVNACsQoQHK3XHU4WarKk2GyBzfEczj78HJ+r6AJqG
zsTpP2EeXnAZKJlD8aRU/9GSJqOIUkcLxlKBWHgWsWqdk3ghO2ZsLudikdzTPLl6
brl8K8SzcODNTASP2x/SMoDcyA0vTI2uyPPfXHrqguo9c0iPJihzHmiP6zK1Fk7u
cHr094WL5tCwsG/oJSaShx666xB0NvFmF5ez90fIINKIKyUOSzERKFGx8Hf92JIU
FcSGzYvnN3AdcnGaxCnjWZ7t3tcRWpaj49hgDm1E4SH4Q8KpGz7gH9zHzWdTpX7w
CQ3wurrvDCCPDAdeXY0oIXEaNp7ZCSkSSXmJIjcuXpKDr8ojnyNvTsANkXID4xr5
8JJp7sT545+fseBWJOIeS5tN19jKQIsI/YAhoAqSh5E0uYxW9e9TMi32aVwOoQOX
AuIzskop2sDJs9SOehclY1rtNg/SpxiTPx22hRjzM3iyK2be7ucy4ZxJ6N+EOZyy
ySDQYgxcxab9ySboyGGjHtPchATHjmcjMCFmuMrfx214e2fotdqiPacP0jaN6RQ5
tS6xMtv3VhfBO+ROSVya1gx3JbcsJmW3pzhAWG52oI1z2mcEWS8PRXsi43wICZG0
0S20y+T3dpeK6U/UW/5vZX/ObO3vbhbtx7RL63UazhXsmO54Y+/7+Gwff8FnpJxV
pNeP+mghitVBcNpd8vdrP3EnPh+goVZr3re/JSGKvLdaLrOVm7uoQfHood4+FtyK
nqrj0SsitWxg2ncLY/+WYltaUJBPG6cPOTVSm7urbVhExstbvLPJs0OepWSLXi5K
Zw3bOlXJ4bYCqLkjd2QRzFuJGayPT4mLzSZZjLqXDk0H1TvWEskf5ZMU0z218hCK
p/BjFcWqP058olbrKW+KgqiZT5vdgqCbgYzdcyDcdsng3dnzqoO4VMg8dzRAlrJE
BzboulWDTt5coAXBY427dVU4xMEiIT3gkhcE6kBCsZ62KTXOwHMx8o5NRHm7S2t2
CaDBe3a5zypiqc+bYn65zOnVtbnm/XyixOG1ns/13bgry8qWrOVvVJAc/4HWp5QX
cSm0sr830/38QFMHL3v7/jgQjPgcxH6cXV+NKNmgxSa8lq5SGclx4vA7FaDpSBzD
mESC7tfNgk3iHO/r75JtH6qduBMbkxsGS1C+8PJEtyqNFdEF9Pg4J+3/kZmAphHO
Vgg5ahv1A2RVEAuLmjKIvOSmJlp02QlUol1D54JzI5WjuRJUne9WCxrc3n3kihsN
1F1ZUtkeHmgLJQlVgw9I6UObeU2E8hgJT+U3VVJwxbvEv6azoTjspL6QCUQQ2KeB
E2BDerE1zUUdkj1/xYcE9faHkgxAwnU1tWDf1lEBHEKSHwZSOxocI0Znm8CST1S1
TUglSf7wzMqyjIkm8S2q0+34L6bTQBClfBWeZ7/VYwcLX/7pgJaKfe9Bv5wR0Rn3
+NfrKNq6TWLM1PK3t5Oy+/5uxSxpWDX+MBf4w0UYpuItRiDFscok1a5YHMszfqJu
/eX/YCeaZxpmT9eVIrpd+kHhHdqTGtkTwmsFLe5BFOypsX5H4VNorWp5b/sKXv2T
ssJKn316pvak5m8pFfxenLM3S6i2bw5F0hJyy6GosNWX0g8JEpGE0MWQge/z7L74
mGA0irgTKcY9xbkMM4YrH66eJpNZQtRibsj/I4dQlntZWF9VUrI8cAv5QBMp+9DS
jOQQJ7fbd+A4cDsYmIUjnEscgmxpq/HgapprfyZstQOAej4hGgILXGAlrYje96eV
iwmYZlk1QFw8L71CkZB4ZgiXXvI7hUOb0zggpmDJOWeM3jaIBbpk1a+dcWmhKsaX
OhzOkpa/cyNjhmxCcFQYDsfduoY7G49WZ24W5GfZFij1gAZKKzV8CytWjVZ3k/Lu
COmiay16L0mcbmGKwuV200j24reoT6TsCgAQdG5yp3NTsCFARqdG2yqiO60u04FK
DxAfDzvdZJaENx0uuvmsj6nKQfChCGgSHK+UfyJhfcqy1EJIu6J9+DA6Nn3ZKi8J
W0EbdphNfCYrww8m0PvIYeLRAVfZMCPDW7VAgBi29UynJhNi1Mzginun31mOKL6S
DS+Mum5IHy4qaAW8yNhHW9So8KGw/7ufjHBUSLQLbv46AjMqxtR6DBUcYQYMx27D
YBtTLo34azfc5nMKBm481/7OpNgWOR9oKRL6iM5e9C/AZjDlgRgM1dlgdOec3QUr
CuiPXrE5qVxVjHsKwWdc1iY3T8Q9gOpA89RtlALUPF3F5bRiaXNmz9HKOKSHQqUn
20lf2RQDkbBxfXm243XbtAdUZckZGb2+RrFsNwll9mN61KZ8uE6eL2ldEZBy0s/j
ejLKpnhCNXNKSBLtQR2Mb5t4LdtEazPAD5/Mi+YelC1TEgy+qP//9SDyJRvkSx2y
B/IgyHh7FrA9AxKivQcBXR+3kuk95JWqASYaHEhj3MKor05JUQDoXnK3bL3EOWk9
QmgzyvUtv1UJ2soej4Vsj0QgZ+xLPNqbNAPinbQ4Wro+Va+wJ6tWtsiojDGPtfsm
GyBNvCQLrHpYi9A4294WVKe58Tz/gsv1F/d46R0PE3EP3+PHHuZjeCFu4dcZEmGt
xrs6h5YEmT9ArM0oRhYtsGgQafTRJ4dOS3iNBtlRU7iwr4OJ/NjfAPjOBaL4klcw
+G2ntHWE/pUvdFFDQiiu6jAJTGvD1cWIONwRE/rUb33Fn1UcMM2wXqH1IExKs2Gv
X3e4SrmvcvnfVHgceGwu1eLxFQ5noWdIePpiV/BEgX+3Op6T1YY/03MZpM/Wmyut
1cylwEuuwsgWrHkkR1yf34VLI2rvXNHtRKzGCQlIaBy+lTKQbhEc23TUHckKGT0Q
xH8jgf44tFoxHrTxLqjuXKagSv6CLz1IYLC3h4BanInuOABZwunfo8fLIUL8K4g+
j9fSJDLgbDafcb83A9vwcR8677TqRlbh7sc7+1KXY/nq26Jty2cd5oZLFrycsN+D
FZz6TE0hJy/8d0H4jPvGBJnbUDOQyi99RkTvM8Egg0mlxafSuXt5GydhKynUoi9V
9u6n24o3FcW3PaQ14AF9X/boEOq60PXCN3RMRtvUVytrU0zpkBzJ06/TIk27ASQK
zUGV5scx3NnUXSt1EmooppkLFetsIA61W+fDYaKaauUq7su6Hlu9r/c5ksSFkeJT
7dCwTH/jx8mNCUKX/W7EjdvOsaWhjvv/0eoKL/yTMji5SSFWbqGHslKOrIjmnUsf
onK/3Dq7/pTPBZYEVcHMlNkOoilJoOVgxQmtgh/v14AI7hkh7irwk47KwY8Ot5uN
BYTNmlGOTXydD7/gCeMgs7VVCptWhyjSxQeCbbGsjm+kD7wfNesdOBNiiu7CmtRE
NTm1U2LkbF0Bi6N2qSGC6s4VJ+1A2mjX4pDF3rAOvXEMJE/CaxOuA+XVhiISV5ap
5Bw+fFwuK3FidXJXHkVKM1gitjW8EDU3Vzght0pZL0lB5DesGNVvuJAb7wYDRXMu
i/+ZXOOIEvR5D3jDJpF24K4TTNFAs06wHKWp3VeNyOYpZ8Lt1+/y6e3roT4Jg7i3
pcS5RVZRttoxIS0rq9WI9zb9zENFto2JK1fbU4gX2+KaIU55ofiTrIR9ZKW4q31C
iHbb9K+1mWoQ0IACVliILS1fxSIvOYF+iHNohL30odlf7nev6YGrWQItwCt1UKET
Gjd65xBM5MXiLhz+gQ/ij1BUbdHT5gU26772icuz2LLIcd9aA3v+wH1wka4f9urI
BUdXY0TTXfipetKeaFrkdaF+IvmvYf0cZUjn5U2MScFoGtEyzp1o9sI2shekXWRl
AXa67l+DvrvwTRggZi86ugipR2lVwBztzvnzVR+TgiY4UKy0MhGt+8YlruY05PcX
g9CpBqQd4KIkynft957VMuY3MMpaaZ5h4Ww/+5HXFB2IoWjanYwxz1fF5Ps3SkbA
gM86SramtZ4bqjWG4xI2tSWdGcU5Yi46lI3io9d4s7FMpyXLIjHG4TGFCDfudv2T
rSgLW3734je6YknHIN1Z8RNSIDxxmmghhwqgdxEmpGctJO38Neo/9wiIjoqVUZs5
M6UD92K80C2JHBzC6bCpyDhAvr2oD/n+KF74JrnJaBNYvN9IllrhGdRfrBfQbBNt
Et71p8norI6NKE3GUXZPjja79Ca6DgBUo3FxXJjdMTQIUU9mKJ4A9M6CuAotRz9c
0Cow1Gy9obpe6JglccIvIoOkvQdidevr+ysMvsg4yAEOE9SIhAwEbbxVy5Zq9PDE
anE2Xf/i689/y2YDN1fpGZ0uAsKTDaOjd5UJzgA+zDJoqe1UgR+mElaqlW0J4qme
43mIa4HHTm5wSddt7azyM5iAw4005bXWNlSyqh/KlgHOPteMBc98QNcgRWB17PSs
jlNi+XQFMmQ5WpnB6Pb6Cslc78TKjRk25T/AiupEx5hdnGT9Qt6DgLa8BGAWB23T
G8uxUVS6Vg3RLjUoXGURM7OHAR+u1TuK36rjCI6gU5YOd90LsOZPxvQf2x6fUpct
fV7fHLWh+Nv37IEoknbV8DMWNnFok5QcfXJPx/yfxWmbMGjgDUXNnH00Bkvp6jb1
JAf1XUSGeeTeFk1Y8UYyCC/IRXNs7xF542TxFJnlsiIOwZdcqsTn04H08kBHIV1W
UXm9XHNudXIo22yTEcuB7Hx+MLUNucjnMKjtvIQcOTKUaj4ESuAb5Iz6FepnbCi4
+a2Xqb7uM9ZHEd+SzgR2QzTBVZP2YpZ5MDLB8VpQa2QqfZh4V9On5hL53XNB4JZn
Gar2CcH+tky/JpkpfdsHxP322qnhz8+7dzNT1yPuNT2+yli0sXdvk+ryTMDKDQQS
CM4Ou+lRST/8o4Cax5+jtaCqYFqfuKc3FSevXYPEBv9lk/b4SkOgvkx8ZMEU9ot8
yqMS1F89LecWotqJJaT3u2O2hyXYZpCDl8NFtThnkTMJtur4LTFJdxeQ+yV5l88J
oL1K1UcTOpdoHEa0saM4a4skPeP1awz8cRym3sg053WJk7yJY6VLdyYy3BfSiIQl
MQfPypVI/jNzdLyyQ2i2tLXBKvtTR1BYdiiKyK/A9AwNV93pcwAyA8WfmGFs188t
YLX0HfeDZevBMCc7E1121rEZBOwrh1oECPoSz/PUQV9kQcN1I7x8ocCdCj7Gc1Cr
ZgjyWOqunNYWMVRHLuKTnICSUFzrOgwCWNN7dr2xl6WBb6maL9j88DVat9b7ktKP
XqFRbrrM8xzETSizXdIeRnzx3pRqgnoBVfWzEnY5oLbbdfgAZpseElYT9OSaZ+3o
7ZCoCLNhpEk0AyBIRD7iMl8YbK6SnPl3EaNz5SoB1pb7+ghn/TMfN38zew3f8Qgq
7g4w+DEY0xQe1L/0BzvthcxXf2pJrCDdxfk/7RrgD2SlkaHCM0k1k1cyLtZ6eOgb
nN3t0fY9VYyfLNiCvgSkrwY40RIwQzDIQTAeDUtkbuJfbQ+Q5F/qOTpEckCI909w
wk2XWcgFCxFUtUXHdU+maXSThh1uWqsSKc4a/PX9MG7GCqI+RnnFmfT38B6/G/hl
Gi0lR7bz2uzi9hdVN42i8GCYbRSggWlqYMHqA1sjM9pignchlVDeI4BWw5GBdddR
FGMGw9101DHPcez8ua89cxQ5OARndut2DcSPw7D/e1qha07t7RtFvb6m49h5thnO
mnXrxj1cNBucLHCkzXg7SVNnTWXtxhqHZiL/zH77CfWiziDlMCgfB05mZeJ3oppX
hiSyjVUdHMs2gnde+KCQPuu+rhSZx4KY5tOgJdpGikeZ6WN7b/rzJWCWilxBA8hH
1WaCiJWI05o3DH0yojAP+4FAmGXY0th0vdQaGAxBCh/J7/ICW1a7/6OT9QGsPNTZ
mz5Ggr/BhA7sFLw1JIIHPoHMwMN5l0NyNxRMQR0fXc4HeR8m3X87LlUn+MyHFYls
ZAqYCFHzp4Mwu3RV54I4D6RUUiCHjFPAJF6t0Xfp9HlrNmGHIMS/AALW+xpM5Pud
igxRj7HDKOantQ3oYV/HC+HirEBs5uTCXPMEEIs0YCxRGgbBBcT5CP2Of+gXeRZm
4Sy030qOaqtspzq7VZpZKxLZxmEdVf7+hDLVmsfnQoCPQqUSdul92xMty8W6aPQi
v12gtZrRnafwtJ3F0GVeijY3m3HcaCK26sXoCspiXPBdy3n+EK3r0bEFD3/xSvMz
OM3ZJnxVH6MReCY70dUu9Upl0SUduYIRtvMzgdkkeSpuf6dwjhJYtOz+6cFR/M14
qbj5UiDVRdH2SybEnVONs8wDCLrAJgXjd+a+A5hLPleF6sxrj4/7UIbV4VoawqT5
7Ic6J9x32y4kL4bdhiO2BTn4TqaID4funoa4VmZAt8fVdRpdwRHhz3CP8hJIjWBq
HXYzK/w1cwIHnyxydzGn0M/VEdCZbYB/21kfnPpLuJakjX5IGVmMHUu9+ePNPaB0
py1xOd2y3CjKSaueAP3bgFFjFLp9wVPijWnRFxIuSgjxTrNE3jR+4yeRHHoxBYOT
8JtUW49l4j5VpK3MLgrXAQlYAOL6IgjYnZMB++LbIxL4r7gc1mqCyDt7N4jYpLQf
HzT5ZGtRjFHdyLdGYKSTJsR0JsUBGXtoQA7Rt6oNHbsAKd1UnUKVQH+H+h5szCrA
S8bqyvElzJ8mS0XplilyyFkR/nkG7wvNvVu5tDlezHnDxxYEHd2X9sh42xEs+UIM
wncCoOOH74Ck4uYmQ0B+o0TqV3S0hA30B4cAgDlKqomIfFyXehiDvaZ24sKfZXgh
BAMKlY1c/cv0h5VCukZNfK4w3dxXWIJ6S29ATTwv1ucQ/Bclrj/EePHWyy0jeo8S
>>>>>>> main
`protect end_protected