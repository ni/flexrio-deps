`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9776 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTDCo+dgLeQsY+vdYN8sJUP1HReGyVpr8a3TTtgVHLALl
xz5uSiBt5fNelWoMkbVekG5f4tF4sqR/lfyQwlx+XPWkLuZir1JDWRYNgFTXKer+
LenAFy3XC/NLNaF9k9B8uNoRJ2UCkeQT0bMo/OpcAEnNOoaBHKzRjeTfpAUvhKcM
ebr4ahVw8sCXn02nGpC5NXCQG/ix+MoIRzIdxDNF5/Uw3JvXE/XUY/wb8EzsWsWI
giPHfaBPffHxofEG11W8OHSsCh/8P9nkpoWlKsVtiVX6oiH7ynmo9Wn6ID9QDxma
0gJphvztFUi/clGeWTWFCE19EjuRHl3oMw+jNF5Nr03B9DvHzGZFoa93XfVkAGMT
+lvf8tKfmDXxH2njj+A7PBankRtWqv4JSuvRwakNkTCTBJO8GQw37k2NA2Hs24m2
W/fLnH8oPDDOErsORvO1jg5CFOZlNPIIVzYhjItylYOljkQS6WsGtt0ooEalnaEP
tPkApr7GlJGzAZ13IsD4uizdMf87h+WtoR0QDZedX7qiEnvOtl2d/y5rieF0BksX
2qTa4P0mALPlOCRsEBAi5rMxm9dMIgKKRC6XTrI45N1xMB0kgvzdnJrXWVGiwy/o
Ql03o61E1b19CWxDfJ0ruaD3kWAumK4DUDNqYulG7e5bfymXevb2e5NaUPdoUnMH
d1bCbSkLMXtCwl/Zq2TdhpL7Ci5DEck49AKe93gM6G3GBX6AaBkRYPjHQO9qfc5U
S+yNX+FLf3NhhVDzHHj6JmGSiG4SDMPpmxPW6pyzqbEECxcj7wOkuornU8LKtTRp
9cyUOdCF6Ycq9+Tm188+1pA1ibV7V0NbYVOeVP4Nofer2JRFJZbqXl4C4riuW7Pd
Hlp/1aHJZP0He4B9NYfoG0jViQw1QRW5ID/BatNhGm7mB+jtRcWZnLXu8t4hklgG
6gcoLLUFsDv8MzC+wbmFMwzyIvjK9P5fzMTG0T019t03+xjzGo/9luNkUb5WxT1y
+BgO7qI1mOOx9Q95s2DfmaVM00e2sVJaYZ2xj7Gc2a9nuT5IDePmM8s85rWGn3GN
aFr/qC3NT8n6mGS+oM5DwxrLOV8Cn38GOVgAdn3XAhsZbwqZuFsjkClq8+oJmrr+
wQp9Mqt1nEj7+r7rwQK6WmUstZnHWu6Ex2YdRK9GmhDMczxuoh8UkW0MpRzx+1+D
tAaPzg9zssl0Uqf2h+xwZDPVhJHYY6p1iJmZ+asyjzDi3exn5Yl6VIHRsBQppeed
FHHrvP8kNsNBE7qb3iBTBOEQkJaZtaQC0BDehtBUCm0o0ke3fTFOtsQdPhXjJwBU
NwqOY7Mb4lm98yoUlQmspx231Eg6BMjA/awmOkQ7NKGsQAGToOs1mDCKzR9a4JQR
jGwI0iH0I7NsKTIID+gZ0CMM+dlBFUA8vnKTTCnkNLeHMNon5ze0LW8121cO4eEx
hZnWFrYi55Gs96Zhjg0iZwQ36BIzjwm+DxhdpJ4yx+7IilcOMcDmglPPt2sShnl4
HOU//a75m7FNj7VMQr7VKW1BccQ7SN8LRSoQQpU0OYokgv6tzL8yobCXfTTyEYWY
SzC3oxSQVvJN5n+rpccI1de79VKQeHfe07HNaYte5PbNwztj/FjU2IUohYMNSTNp
Hne8nowEm/AdP62BLFBdtZBmEzID/A+In38SGuI7DSxUSp4c1OwmBdxSqBI3EkGh
lg5JrU39W4HvGRgrGQ2NR4hzT/xKPoWPjDdqHvD2TEDutTVYE5R/qcI2moYkiKTP
DY5qcrFNRC4Nf0D1vky2s1JhV6EzyHXIyWoiFSiy9EEXTv+jhekjuyO7JITVLZpF
/n5sOXLACJNBH5Mheuh6Nuy8dGXfWLIthfKcb2RSak2yHbyoHkTWYELvk+rIvh5N
S1ajFgs29pIOq02JOiMuyS2FYA9kdEJnCxysof3YCm7NwePJvDzgQunEOnzPrzVO
3lEpRRQYJ6DHmsDVqk038ArgIlgTUPNMb6clZk/Df0gJwQX303Ri18T7z5lJ1Isb
XDTdIUXMCquAJWVrf0VIYDRmSXPlchiCyBcfjMey7jpY4/8lwxIdx3lkYsqPT054
6qc7CVNIvm2DxwjweVhgfpV9QvriyyaZXQw6kytgb07ycjgM7UVwTYL35wr/ibuy
DCfgrxWKW6EqQJ3Q7Fv0NOMkJJyhoudlN3W2iIU5JDasaXVKCJeWp5mv8pe3KnFT
8wg4JNX3vPnsLycFgrh3xyn86P4AjDAUxRK8DxatreAxwAjXEyhQGkSni1LpLtpG
xAy4UCDYED1sC44/a/IJE2/w6U8FWw37qEgf7mmbu8eWbf3wUlciCliH/4VNbBCc
6sHk6qLYhsZulZYiPSY+jFpx+lZ8rFP1bIXNt3636qMRSJWi6+NjhTIQ815czOei
qmD5AvzLLC7PuOdl3gTEqTSHBSaZNNPU+UuCseKQMsR1IC5t1bBPoSoed7N6JuMi
xGILz6a1pwcEn/e2A4XLCBBhkJ8w9QgNpvXtHmmLpJGC3UYDE03PeH/ugU3BiRRT
J/hElLWZnEsveMc8gzfaMl6Jpqw5tFoMe2NvnmeXu/2w0DeHLqyv0TQCMZGJflmU
Dz+g2eae3emEOSZSWuUvi6LK5mdToDlKwnuM7qoDg3e2ujohwRf9ZfUWA8ivd8mu
lcTfRFUe/3QKlhnm2XzwcYAe1YKYHr/OnahGCbS85PYN18VRCoI3w7S8pmVK6Whu
DCJ04qVYftMlPNSPvHw5TeT1nOnSQQyWcn1dUeS/EeQNp0T3eoTjsqsaIwS/bged
yV/Z6qDw4WSCK3It9PTFp2FtDDuF9VwyF7CQ0nBtYA66IsUSZKIBkfC23ks2cx0V
v/jk7yjJECJ7C86tWetB5qJ6r1Fdy5A0Lq3DEGtr5Yny60rn75VZ9PEJSXgDPqFZ
Xs8/A8oQ9bTZ/Dnj93rPd5IlxYxyfUyJqPD1jZQjUqoHBOytTfHUauf0EGW8E5Ch
Fx09ypCtfG1XppnziyDwKTgaNIbCGPdNax2aQmQjan3qMXLTjueLNfppbzicvu7X
t52tjk1KiHFoaiKb8bESuRNhtE2+gDhKBDgUX0rurDF1lFcLB4PKLxeA54mPrtpm
Ij6/vFpwVjr/9cY7wvjgsLDBOWtOmGeVvEiaWfIKnI4QGJNEXpdeTebRCFJZ5t0V
GgIUlC/bRyqimJ3h2btZj8Y/O+kRv8dVfswNjksQLV0ZOudlFGk3E4klLWd6gn42
yHsLrKcodqk1JaksAoNt2tlyRW7jA5ubPV01G3w2Y/Jy2koKxn86d3OBrQ3JaBul
kz9pNnGeDXwC26D3wpftwLs0BujkFUvsxNzcYs1UVEGGTjXF8eHMPtr91ss5hL5J
i0brlOZQkCwDFd7ILwMphIQYATml8RhrcNb+4GWavAmf7WlHwfbipuGGM4Vxw/Qf
15m5cSzTtizbiFEbzODTLezFSLfX+Ektp191LnvU6vEauapXCJeZkzu27ySCXM+9
WLVhsqtHX45MRxEQO3/lfWsNkXDTYSWICS8XlWqLjFrkM5xR9BHifMEJxfVoaxNZ
qVInmxQKXxgrlEk+Xym9RuWENk9TsG4NqvfNLQJQOR/RmOCkwB5XEh9NW6jAiMJ+
mxaaUFh8/PqmeOB9frk/2HtTwq0a8PlXFgOYFJlDrFcsMVlB60dIIe9+1g+d/c1R
mUl7Al4G3HQnoMKOnFOPkZrUWMyZEhc349BST5IT0X1S5MqrZIhqCuDdMSHMbAdi
ZctsFvao+puAMT8QfkOiDb7lR+6gQ4sCX0joS//nsWwW0i9HC6Dw35zpaliVqJUS
J+J+GYItIPeYj7j7yKBXN413C5KIFmGHCTvfTNkTbBYS+HSNd/rmlzGMdCS7QNEi
m5BU6eKlxzamr5nF32KsYVqZED6CDgNRqweDuM7PxO1cIAp0iGGpjxExXQ0iGjtx
e0hKBNq3+XoasS99BwzslTVBu4rGjtifVzvtVn6AA73uMBq7dvc4aam1kwI0bIpA
0imV4c+qcG7jS7OM9zmSoBfoPEclzJxpeF0QttNhCe4p5KxSsH3ydcE+0njWO9EK
iAjcAZ51uK9h3Vxad8+HCk3XHftCRWPW8eu2m87X/t0FnqFe/9T8ohe1KWjLrAy2
3dCo65YgALDht6RgHcHCI/74VOtOrv7Oo1P6lphbQloxgF/yPGiGExHeVh1dqjwu
Lpjg97FUZVUY7Tz2GI/F95cAzq0Xhbw2RbXxxff3bEYOruhto6xi46+WcYRjAXE5
AcpnXpjtZiRgnk5ZAccqQTKbtgjpekx0mZLS2MA4kbO5eGnyEk/yRTm/HSiPwI1u
rFbEkmC/L3i38mQYy9maUwvjXYocyTZPsBvRMFYGXw70wQ5rbCRimDyIeOuBbQZY
e7m2e2f0qjYoYZ2/R6kZbBiRYsQVnZTSOHTQoAXaslNKSscZOGdlioS9Julv9Hm8
tU8kkNqmL4QFVHuULR+Dxxj5FB0Hsrd7p1SEtiWPtED2yqceEPBdnpEE0jXNeQNt
efynI/VooNX+4OmAdZ3taya42pMQcZangXNM9EIJE5pko1WdnUdSN1oSxfbSIJ7A
smoyUg8O/ZdHFxwIcYA29pH7wYDyUoupLLvo97tRy/yXRgTiKCVFMZuD16v/Yczj
I8l14rXVYnCVIXeeaHnyM1ElhNrryshaHUx7dfyUyTRqtTsmq1+faau5HtZgp93U
rFc5joTyN4oJkmHvdfJDn6w3If2GX2T7DIWE2LFWeUv9jNUdgjm+TrCf90fIkh+U
1eDN2O+9pIqHBM0TW9MrM6kEd6kr2SbOJsaLa7L8RhLj900Nd67c/dYPH4pau7c9
TNAZmP4rw8LI8UZaBgQrUbKCexN1gw70hZp0LBgpQcmI+qw5QiyJa4FQok3f+haz
FGgO6A3YUB1gEHv5q5jY/lswrxpyfzwetQryib2GJyOGARPqBftS6PXpTFNjRf7v
jl/QUUcxKTnMB50IAQmEfXORNOAQWBd1he4U5DA2JxDw+vrYb9LHV9AVjr1pvO7B
1u4GWHpXfRGiMAzeYNCS06L3YRGu0CInTcE9bz4zH0YYE5TnAvLdKWr6DIqh34nO
1V8/bERYeS+PjetUQflIj5biEGnsFgklS9/BV/3ASgBdJrIY83Q2y4Ehw8T1383Z
LwQzQImOPZkrDTgK6Iiu+L3tZHt1MqN74Yi2szhbBqzEqidASe8Xd6blzhj/vdL9
mg97fjrJlNMpBgXHqP3KC8FZU80rc5uss7LBStq9i4/I6gMewU9DMmuS4BtGzXXi
OhYo7M4W1xCJxih1fruGNWbZRa6dms4RE0PlMmh5ITAhoNF4m1d6kKPEyjg20/5P
XT7HlfII3GVr92vVK8cialok0ah+eadzaLzqJuxeGZ/pSjQVV/jC7si7dU0zwrv2
0BcKeocFiaQEnW/uswF56AHxbJ6mnso43cp9lx27z9w689Gz3+O+Qm3LBZoKkCXR
DyUWZgxP706iV8RxTIMFMx9yviEbo37i6GldJW4tZMqQWr8MHHWibX6l1YmiKDRk
JQng5f+MEajrD/jiOBp72L8xv+fesP+FayTfyrEaE/vjF4ZZecTopHFP8WR//+pG
YAW/Ho7mEghUAj6f7eyoBjaLLiWaB7fNsj28a22GWSNQtgKjYtpBcWP5zwN4vDxk
SuSxE7QOlITNmy8GD3Xm6cGvEgekNifev8eiRjd+NEY39rkri6b8Wgb3TlNBzZRR
4VIHatM0kwbKM3Vu/m5GNgs9/0OucNYYWuhg6eG604bCCT/xPbPPOZERr8NlUlae
jA0juedRCWpJUS8s4tZleBcEx09jFlTwwlPecEYsLxObPyKfJfM9u7ofo7eUFpk5
lZyBv8bk9V/uDWT+u6X1eEbrPUW95eX1fkh9OTd/uyLpsIPHJgp9B31xvz5XADgU
T9Yv17S85DG5BLLrk/Y7UGQg2jEjyssT0jKsklC6X+5hecz/dCamCE94OVzt5fqS
kvDhEiwifsKz7XfOBlXz7DImJ+5cYBvQxMCcskC28OXb/vQ9B9bSyD00nHndYvVR
aW9XisDR1j0bsm8e2VqVa40VtynoSsBlUsUIy9+3oPFcQoUr03grCmsMkf+aXF4r
CqhrWRKvp8+PPpZUM2lr9gzbK2a1OXJ7X1H0oaRY6m20agW0ynPLMA4OLWoLtAD5
hvxzkxux5SYzKyB5HFD/CpXOIbSHB0be9oW8sLIK8/VHyCWTtiXIDaCeZT4VKVz7
XrO9gInIeTp2KGLDb0CkeDXpDJrwjmQMvo9A7MAuvcW1A/lBfwNiWHZIHvt9albr
/fSlZ02uG2KEWq/f4UxFCa+uszggxGnCUvZi4z7XySH4NR5XqV0zwL4+Uv7NoUKO
ukDdpP+GN3Re69B9o8LFudtr7JBIui3cBrHGuKt/uVMsSG+RFAH77JUrda4mQPf2
5ouuPqdq8CI7xNzE/tLAKYG8e1dlfmY8ndjKN1unqx+DHP+gqs/3ObvTIoX4H8Vm
Oy8MAcpxajbaOeEehytVUpenr4WrzyQwqFlQz0uAvTk+a1ntK8aABFw0O8abq9jZ
LQvobZ9VnAaAQAw0TQVwFglSjUVi2Y6fkdbU9Lh8eBk5gaXvXWa2gGAOzDZAcNK7
IUO+YaaX9aggOxeKaqKsLQkOlafuHomtiuv3vhYbfE28rCASgGWkQ4MumDKcjPpS
sWHWV90C3memYoxBjcKvxYwsCzHsu1LeEGowh1kTNqPbkBFd15YuXW2dOe4HX3g7
xFM3PmkkuRPkKytNFGcNDiMtJkwdYy1u6CQUW8sgkW//aZ13op/WpqKoF+Yka0KY
urBAagNUfnXLlOeES4GMkF04fdY+XnITRPsfd4OEMfVMqg7ruW2UGQN0oRtyysoY
qhWdjCO0QjWk3kqDoNfGvExiJlBO5VtDU1hBC8igGGIpF3A+lEGy+hUDEfyzc/d+
8z9+McER3vemY6KDYjmqKzXbdmXK0kmBvb8U4nsSESdGUpXFj3zY99by3GbevIp3
Ja+t20CjBITirtkP3SZiIoTSgdGZd/zVZyyg+lKEVlGXtFS3FL3IQXqjhwZYG28T
+JGc3G7q8Hk1n5OoWSKRmkzVrsoOXTsf7OdrTn3P7UyjgOJscjZzf6HWR5lZyl/D
2zA+dguQc1p/S9TpM5B3hktieLEmo/pchY3+Ybccvod/2s7nC2LMyuZ0ajnoD+Cr
TWKFB17KV3YtkE/ualMZE+U1TlJzRo4CfMa7lKzCuraSRwNP+kFIK302hFjdlNfw
byslbUkMfaW8I+hvM7mZriZeYseSlOB2n29zlciebHoz567O4kqIEDtlpw64SXj0
m9S/6omJKA0CAv6HcE2RWspzKC69Q+SKtwP1qHk2h6FQfaR8dnAAsOx5Xx1iWku7
zHCfskYBS6dU5CgAUab/wVMQ36gDZjr+HPcSCTd8soP/KJhH2aApg7odCMhK/ekB
ENzoQ0J19TsKiS5Ziq6jgc33cFc3tWW071SRQvm1tEBdFdOviFjlQZZ8CV+HDfnc
v7dv50Q1NAAwMPZyMEbLgzzEfR5bSLfEJCGzoapc5FmWg26k7V+3oUMzHwy4vQ29
ULDy+t24o06jdzx7ATxmfMnOQbPLNGunuFy+vNbmlvX1qtta2XlMGZYXjd96N4jO
Y8ZU5uP51dHxgSJJFLNLdme1wAWeauboIYHMuTF6NYTmEdyZplHMal4GaeX0iNlA
F2jcv2eNTagbh+/zinPez5YG5pau/rBqS1BetMEj83C4UMyPc5ctsCvRG1UY7uDc
9XQhA2s1XrL4o9HFsuEd7tfcDT7Hhl4UZxEIlLH+si8o4rXefGNCMIlTxFq/hHas
kdx74nwNsOV9zg5XrLaPwFYFBMrb8mdoVvekMc9kxyMgc0XrHCUS6fQP87cg8pr0
AX05e+POqC1EQ5llETkQe3CQn2A4zscyxEji+BdjS+I0j6o16xeysPbZYNKf1qyD
VlYVR6vtAYACOyLQ5q0Nc9Uu+m0p85KS4aLrsnjufwCzBDs2WlPHMnaFFJxteX0i
80HctVZI6Ik8kf7+irGQRsyeOPCP+TrW35LegLw+cqrYDeZw+fr345RbgjIZAd/u
TI6i9iA0ikvZ4UBCl0EuzS5TGxZabWbe4gC7vMy69pciia2+t2NeedbIDHr4d7W2
kfCLrjKcqi/MYzGAvrQLIHAXnRXihtPRDPaq1bQF8ccWjA75Mq4aG/3nSQZNEWRv
iwvGHvgKE58AVa+rXNOyMiVdIgEI26dYORPRtkZst9bCAjqfGgSl+KVByhuD3cki
HOqRaEM8V9qRH33GL73ZQrKT2wVHRkenjjYgp0M93dwSt5qfzCulLuU0tjVBL9cf
i1bYgtpaeoU6LhiXik3/djbQl3z9uLfzPR1fro1zN9AJwkHNG0t6ERvDz3+nsb4s
+YbUJyansMJ8PQOHVjfaDHPgzaHJu+8Fk8XEdpl56eTflBRBBT144D1bmUDTfw22
BfZmED6jYNHfOEFTQRw0tdhLWOQ0Ol8i6Ukyrco75z39wh6RSzgICURGNsRTzTlk
MDJpyb5wV38pbelek+CqaZ+rbdUsN7M6cFGDEtTOUWiem3UIgqGi6ZkdA7g4hUyX
+Kj6S5Zc7y1rIeCl9YQM4pYI8EH9STYg/C8hBP0epAF9aK5iDkCc+ySEUpu6sKzn
tMk2lpRuKEga01qvkWiSDfWjHjU97WseQripq5LZ/HF52SQsMU9ssT5QXoFWDMGy
OyeZEaYCK8A5pw5c29RLKx8vxGRlH3W6mt4QDk5DEjDkMJwT97SoMpizEuxuZwGS
Jo7UteNdkcVLNLF+M57hzwO3CqI5S1NHzXiupHaP34uNKwGzzmIj5PTJRR8P6i9n
A0MAXlhpKTHCQvYzL+W3eschgKPqkGIoRvDMDzv5xoLbe1krJWy8qkjQAv4NohIK
7GPSFb08jETagXKH1R2B8NMwF24WaRmMK8+H35yUsZ6nEubuYAgXK0ug6VpeaZEW
jo8CjOs0waDqyLNgbHDaDiRiQ3omlS4tjFKT3UoCFNkQgICVhjqjXc21hTPcDwUH
98DbywxA9A8JN41ygr8shXIHNOTiUgnLl75t7fQ5vunaCdBTZLLt/+hDu+heRJUq
Q7cR3g63xZDSouaBzmIEJJpzoWPZdvEjgc6pKvgmSUj2I1sPR4tK6h+m8U7JAtP6
UHYaduKm7qgXUx5KDtKPHXtCsgmNqs8vrdAIUOs5mmKfSEPYi9JqRgkhpcBTUYl6
74EywbSsBE1OTqJFBW6uAb869pq9RPeqA8jXXdwMMd/FSPA/5s3YRnrTlS0CyJTu
dGUVGL7WtEAtkkA/8oJjuxPalx5POnE+dWmj6a7lrZzuI+wo+M5k4xlGCIhfjEOg
vY9jzWJWC6aEDqLfNLBESFF0VtUm825t61SlnjvLNqLznQ9ZLsV/0Ni18qhs/AKR
azZiuCMO+ndx6qYVdh+KcdKmE5g4Q4ja3/MC9gvjG657OEoKAG8yGWyu7uQSseIb
0phVnpT5Iea6FhjpQ+8+derhB1YITgjzZA59ohdbkEpRnQZX+H8GPDkyup3w+AQX
Fr91QhLFk1Vv0u1dtcf+v/RSESAqFLe4Ht6m5ybNr4GsV2BbUWnzEMYJFVDP4MOt
UFUmRzWAAgfMVtuMj57ZepSL1Y3oC0I/OgjK/oRrURz6b8FymLNEWyawyXePi578
u/2UGGduo2BufivLt6Ygjpf27EKz3Fd9s1wIBWubSvB7eH8qx9BKpobiTtBAcc8H
RlcVQZbuJhyJye4xn/jNwzPS18OdCpzUP0Xsol0nWPflGiR4/2gHCuAmm4F9M3OB
ut91T1Ve0bDDoA7TpnYHQQNBOQfr9cEh/cfnZZvzqQUlEdaIlu2+9eQfzc1XXGKP
7NzCp4YiXHftnp6sBaAMVFj0LO+a4Ekv+26jgPjtSTahuNiwbCEjApLdgHWtbwbt
hC82lTy8MgzmWm5Ts8WRM2+X3LNtX3YVT1FDnuLYoiUP5FCz0VQPrCV+Qw3twnQy
rdx/+gBIznPxKRVsMZDSR5MRHJTptBLDEPlIPYVgrOhb6aYOeJuJ8n9At0bMXLJi
boQQCknB8KDayc6lz96DSET5/1iNYCzgv6wYijY3PHGsDWBJQljocODHaszZ5B3m
s2DBQWEFONmbg5a6L8wm80QhAxs5s9XJxKwX25JpP3bwtgkzOAfaxSDcAIpS6P5P
ZNelnyIgo9I9sApRiVxDsP1n8l1iKl7Rxi/1McwSKK/rkAR7aFXl2e+d6bqlA2ah
Rzbdg8NmHvg1JIOaYApuJJ8lYmqCKG1CHPiqAJQxQru1yvciDU+5ZlOE2VrL/A+y
9ebPTRWBGgyzlADtiV2/jW0HfQBoRi1ppqvJVimLiNguspj3uJ+1tvpPi0E46App
eVT8oJ0Z5tuFbs9sykt4JPyEd5hAQ8gMVu6Mb1a1dPTKdoqog4XpxYFmbwFDYyQj
NsTUQ7xhPISxAnKxfU63lLQvrTlj2Gh/oQ88bc4/Cf6Zs+48DUtOP7s5X18QJ/hR
edvwtfon5Tz0tNJrhwIpVlJNtITs8a7oBo7yWgT2+fPIKjw7oWg2/qgonHidrryv
U0SHp+xnXtw43iwvkyRth4DkASxjjPtRwMJynN4FkYtHA1kAQHqvUNE//MnlmKI6
ObCTP7alUMuxpQG5wjPs5Zge15lrnY2+Xj8h6spCQP7s47LT+jXiGzcWVz/eyAy/
fsCzarCsCvdt514X0QXBT2/NmSVrphcF1GFALJWpo6pb0N8i4ZAlsKxLpIkhu4LS
9GQer1ac+ElekdtHafmb65O59obf+ZG6gUr/Kuyq87Wh+PSRskU8byt7wDu5xnJa
EW3jRmVO0eXyr96BNqfO+d3Z57gOlQaEZnoUstLZwop0hit/3VjRSupjz+radiSA
x9gIb/XUyZPd1pKk7GkOs1bkVhCPbwcfe7NkW22Cp78dqXF6xSav1U2DC+8TjEhq
2xlHV8UJjSwQD9Jo/t1ROHYmw6TdKNIQsyD3l02zd8laup6mzmpT+cL+3zv5dOwA
aklV+g8AOQfJFQ60USz+kIJtJnkJ0ptmaATbe3N+FfvOrS/GhgrHscz05WlUQ8up
HGlldxWZLFB1pHjAOeOxa/f5EjgwIz8yjZTqKB+D3ov11j1195Tm6q04PgZKecYP
YsTCE422SAcFuo6V1EIm2Jg5nfI7TrS+TzrchcgPtUAThsuynyFgAl8Gb2UJLdyM
vJx8rch93A0yoPRMYKy5Vq0hPtNUxx2t0fmNSVjQ9ZWldS1Bn1Z+hnGTidh7+3B6
WGzJxMHpBaz1l4u1mf2MeqQNA5qdyBX1T96Yo6FzDdS6WFLtgVrGZlVwptIhWbpR
L6MNYxEYjWCsPuADxuV0DvsJMbgrGRrFFOGNqHkfSNPf17kltN+HeuAl16LRmpXJ
dtFfWa0tw6FsnXGP+gwhXRT4nV1F+ghcJJyfLGIrCP/qcA+mOWjjcDeNLp3mPZ41
VKeOKzL42MQvvMsG+RWIQwvSYfo2a1agKYj6YRK69HITRYkr7mk7VDPQLJzEyBvJ
ruw47f3rRJtDfJd7v5otdhEZdsJz174gCZh5a1G8uCEzD63/Bd8FWeyjPGRLMoZp
peAHlWr4Rkx3RxY5VxM0L/YsUeyiSF0P6VQ/wASxlki8oIDdn4owr/HAUkoPCu1Y
HbvRJOfjRwTPy3LAs7YmLjDh52tjN9/UPfgZf8iKN7HsTPvR0dTzShgRL+e38cyC
aUS1DmI0bj4Sgncbli93wf+cQGuCVZMkVKrombW4P598FDFVOX+d8Qn7iWeMez02
sm7Wx9Dou417X/oqTg2h12K9MLtdruupASokZnrzBa3MGgXsduwDPi9XLxAtN54S
MNpzTqU28zevA6qZjGYrAIm5+Ff5sEGThMq5XEXBHnXW6RVTNHoQA+0pAB+3WzHo
i5grhgH8FmsxyR+xk3HP3uPGeafW6sGr+LWaKdi6pkYgQk/ABdd4bwAqf5oI4c/I
1DTZDdVwLvQ0OwYrGALlGTtM5/2ASOxE1x/OjvIRFLlm20PaZ5YrwOxIppPPsuwO
j/CH7i6jtBkS42NbHvgjolK/2G7cvRSGyRUQ4ZWG6MFXLgHSwmOJgJcLfSgxzFAT
ig+TQqSQTm4GwclMSMaKeaJ1C+x46YYClmnLUswyYPKULz2LzZAdBBnV+TsZ66Kr
+2gDTUH7mHFYP6pH9FixPK7oAj+3XgYwPlFTPl23rqWVqwp/Gxyg6iZtTq4Wmoms
DdVhz1N0yZE0unXie0+iLt0vbSgEwMag5ZUur/t2Y/PeDth5M75fiPPs9HrYzn4w
+T1C+yGmcJDBKCCL+LlYobr8ov56pGbOV+i1HHKKLYm4SLbT5YpyP5ZV1h1kG3Vz
eqnXS7qkif+QY3laie7Enz/gTLbr6neqyFq91/lRsYYDwTHsjDPPPrroVlKlKE9a
L0l7osCCjzCdQqOKUniWTelQVJtLGmxhD88OtlgNvtI9xlahzPclFVWWd3JvF3rg
XrZ2MBbJ+YBGfgTYg3nDZKufgPNNbOMI2pFlwhM3AO3ALc2k335wDtXyA4BTL/z1
4s2psHdsPplNfsCOGusyJMVKbPHdyuVuSDWfOl/mLLKouGLikEXsE1kcn7IluSDt
i52lI93n6b5Mp4B4xUcPZq4oJdvgY/pJNr98x1/2X1hIHCmIuTkxyWHgvei8h5s1
mMeQ6A01aFIKW8PFaI0VyPPcePcrHA0IF4NsjBh6cISevfvKVDzf8QQw3yY82T9C
+qDCu2QrvYej/sMb/nuCQd1ZOVvRl5195jnq/jBlYhTUT/5JhMpxf1xdQFIyAaVn
9wYY/wuLXjGkID06NQbmgqQWAChN/YpsvtNYFN6e/CA=
`protect end_protected