`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4368 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRhittEAvl1oG6OrRaxW61nyEgtczdZV0JI3Q6Jk/TZs3
rrHzkPZ3ciDWXIH1wFEHwuQcvkCLxL13qoqKrznCbQ1Hf+7eTidCAXPXDfAdLY+I
kM3z5ueMtTztFzOOhuroB9Pold1flPkozfcxbvuWkQIGFk8GEIvLS0t3IkyfokRV
kMiBkBzcax/l52/lDAS1/Bx41BftJ3Wus+xk77W69hbjmGVjiPn6poQITYqF0Boe
3JUckCOPeg+24Ta2uFPka8h/UMK/nuLSOT6MzhqxJbsBCdt0+LuHuxVFliXyjSFp
nzOlm3UHN7OvJWr1gWFo1YXfQy4ijCxGIsH+GfI2m5mJJX/ozB6ceq95XIMFWfp2
RQlISB3bIuLQj9aU5CcmJpA49uh07ah7VAfoAHjEEJ1wA0ogpvFfmkvUZOeiny9D
AEooP7UhncrqVczSmKtLYwKv5KAMKLGW8nXVRTmQcXWd/aCYlGaARS3JbSA03zmx
lXmQevWKz8j1v6GmzuVFBBJ82+h0HVCFm++lkp5u7iU5AFX4+rSuRU47hyrQy7F+
XwNNMq0BukifM4w5kct1DqaUzVMHuPj1kmwezxaBFyUtnBBImjRrDdPTrE96nDfc
CxvM3kwtOm8Is3uKKspg2xSG/0kO/R9z14RF0j6XsZBOV91CLmQJvyEcuk2MCdk6
5bXN7rfEieync+apTsDcrvj5hNkyV7v+CRd0Tpyo64QnmsroGKqGqkhuQlub60vb
TWAKLY2gcLuU22CVudY/9Jds1IFD/5ppns1ALcCpDy/3MnKzt9z6UzWYhF77D+nx
AwSfVgMXEt0sW5m1PBeSKopKZloyKpJDUU0FvIkYc1LF1wW5zfl11/Wp6vRsDkAq
KrSc1SPZ377JwtzO75RfS62tH8eJ12X1UmtksdrTYDmfYUSv2GQVvjwClA9qY/Y3
y8eB5/P0bP3vtJaRJP3Kn3eMtP5sh0pMgjdqS3iBVim53bvJoTHazQ2Kh88Br08D
G25TeAZZjC6ZTWmQOnryVHc0fDY4rrYQZTnx2d0wuurWAxzql2gjfsX5R/1n7BwB
u7A2HEKQlnw0p8dTiYE7WoThmdhvRnvmY5YfRjY1tcIZ8ht4xYJlcFrdCqb41NOm
0QxR2MRxL32K1FIXReLb88lQLqeBYDFgzwYj+glOJHo6yzqSoSPHwsXy5W/GlZvX
NIVlyoHFDxlHi6kDnkqIpk7yDMeMK7RPVI3YFiscel/pvU2BxU59vfZ5zphBeEXM
m5qQk3TuzjSrWL7Qh6+Q86Zw531bd16FczHWizrHFwfDtiHdfdzmUqxBM6l64qas
t6XM7pBpI1R6Ldes7iUBjqtqkbiLn9xWxtoNPALEnXxby4Qu1kvJ5zGDlUyO+NQQ
2/zkHIPu5FiFSlurb62MjE9F3UJKOIy69C8rA/hrILGdoAJhDzQCtRBMRAf0hWQI
F+jlI9PkRLqalsCOA9aC1Ojka+85WsanlPCfJx4l+7afG+w9xh+9d0RA/UpCd3XA
ibnDsEch/LsT/MUPHFipNitSKhi4tD0kCt3flPEErtBMzjtuBxTXy/xaNhlugzmU
6EI5RaJ+pxvDMq28RkhUOWsBnjuxGqbzjx/i6wkLMJ0IOkJMRxkROrOtzHaywAQy
pRaGm2Z3dWZ0Btme0YNpzLQ0S3DNQQjRx3CeB7wYf4KGf4sKfrNQtK8s7qCekgQk
lyEgRhMBI61nsd6hidRxTuFZPclxkRmvxMSKKZmaia0eg9EZtGBJktHAkIrXdbN0
aipWvABG4mjG+8tHZhF6c03lPlC3O9ZqnX369YpiFxc6aHvEPAhioRxES4ZMUNfK
SeIzQL0QLwIBpQuxeNsSKMaHQMXUT7hN0DwgDqo/L4pxaigrVulZMZj9Kxm7woTi
PEsfPZyxmRokeC4cN0Hyy6w8r/b61PX6wUpn3KJnEvDND3BJZE7OFGyRzQB69IGE
Nev1fi16lgz8GRWsOkBr0xA6deKrm/Mu09Rb8OBA86Qk6nQPMt/vgiiBiD8hRAKV
UgArS7SQAGTeyjQnBwn9S/Tg4wYCU7s5WM7zNdUQs2aMsTJjoBKK8dBS1aq6lfjT
vaRcs7Qu2aBMHZNdqqNKMUqRvKr8FgIzuizI1u45aiciyfT1WTpdZZ9r++mOrPme
IWh1eF0AR76fQBPNgN2xyeFStkKfHaT6bF/acD467Aix7n8+OV0W3Sue4ReSooU4
qtAUAKMCvSnBzSMp5jZSaN5PzeLqgvhSq7+a69hTnAgUU2x1Z4AMO7wwVWJ4vN3g
t0M6KbXpfg3gpXiKO2XsU7ktvHwV712jnENCEbfAGzOl9/LqX/4Sa5WT1efvUDLA
lMyJjnfFTcir/dltGXb1a4Mw1qN0PPkfD2SLZVLYmEQ7TymigMldNRjvVam5ecYD
vlOUAhUgCqwqwGRyiKCga7mSxklIOyjzn+oLdn4rjTiyXXEbP102qxlV9sfmHFQH
6vRZATHi8/2mfIq0qxZD+egDvDcoJUDutk/XhY2hiaYA9OJoLUNSkv+WUFAOISQc
0Vnm6ef1lXD27h1eqvCxBMoeEOrBfjw/ziVEHuTMUgvEGORss7haBSKiM3+AorIC
1IfVbqSSjrp25ZMMQkDCJMpPk5IvCB64C+K8SzYZqVwETt4Zwi8fXjd7OBHCZyMg
dezkIP3a1LhwdRjE1dFa9nJ5eg35zNabAGtO/FvFTydTQBtclE4O+gCFMmcZwLaQ
ZqLCJ/x80E7yYESYQx5hjqZLGUAoNDJZ8o2pIAQXd6QvQC8vY1rmCYo7xFBQRTUo
sMlLptcQ1dBzy/cD/AmqDZ79FfEqDnRTXLE7DRtfTFJ+DL0tAdCJzSvXkOZLqKqz
CLRxiWCcRNJWBf9W9OwqiDrxcK/S+XHW33338ellxbVEKXFVTxz+zNUB53lAVDsz
99LO5ARlarPjvRdTYn2l9ZHx4g5XEjeEJ2eglGMp+fbMkOSou/mAx4I3V9LQlyyV
vwaf6GXp+2yc1Dne0O5uvpdo0s/TZYYcy6cvyA9LO7tueCrmc4w+jSHooGBI+WWb
HX+83bGPbfFVu3I2ftg8s1ZmqvcuQXXF86F41ypZHUSe9FLwF8I800Hbz/Mm/4JN
aFUs0/Ewt1fiBQ7wsmUuGbRTbYrHyjYUMnEtvO71YShMPnoifirPzt7Go6KnJv7J
xUhosICuVwkxhZBHVCUu++okeo8M/SFeUIyLuUh30QQ8MGdjto2Kw9wp0PCB92r1
6X0mTj1+aOOjjTOWmQam1crebvJFzPvrib8w6PxRB6zLk/vEk3m3uTfhlDia8SLM
HNKu9eDbz0AbQDBMuXjrSlvo/P1sdhueu2ci2IF2c84nkAeOGHauUfMLXoZdSN1+
52tY7VFI8tUlzQmozAZfOZZKAwxuu9AMEvVx+6NzNvcgd6TkJgKF+9ay7gpZtcxb
CRHNSUq5GCYKIfFgRp2KkigMttKd/3g/Q8m7AM/caOcl2fa2O8vvhCr02C6CDgqN
6e7eZLPyMfQuyBOjhKo3zu00NNOTxZ6hcuXOtYPdIWT/AzFVlwt+7xN+zMPM1aAp
FHpbS/B6Moy64MV8FkR82ekUY+RIV6HuIC3FpwvQo03man/6hjv5IjbJXCGNgxYF
tosXYNwoBG7xUsbGXqOvnc3MtxJJ2Tg7p7SgjA32EfnkKTULcnogub2kocmA5zPm
KcnrXQuQN47UW3R4uQTBnGqpseYuF8+5vpEvI9GUqjHAVJSzlCjUpXezzsms/OCA
fFGi268V5QeEzO1Jy+csiNcCVhCUiRqgY9QlfImucJSTXwdDudox1gy9WdhLWMB1
cRpWSJqAaLjlZvI2cB+y+yqEwh+CqN/CGRO+ar7gbzXDAURjvMThS1m0xh6+rqFT
qzZMATQRI/Px1sM8bqhQ8q8HKQus/YClDID3eWkYOMlrgEXlsIdd3tc97XkQveur
7pQEQvoiIsPwDIT8e249jR0pfovE/URNIsC0PV+xovbMHALsj4v2Q6LgYykVs8N4
Txga4DHAO/mbvF1C0nfVfDKD+njZUfMMLDDcHTccCw7W5j7lwaJLMI0K1keaCeA0
qql7pp/BMWTPXThMwd7RoP26sbk7QqstbbCJdS9wRpvFKQ07xOhYMleaBaNWJwx3
ZwbQF7Wc5ZUe99sobv9Htu6wq+jmoTFlBLcy1NWHoxbBhxDFTXCQanQ3SvtFrjch
yD3MqGlx82oxFNB6OzHALGPvK7jzafiapPibgZauoRd1HZvBSagetwXSeBHDgqyp
KqqWyc7e3JdrbsnDlWUBcG1Xmi2GFBhCx5gNsXFEJTZWTUuv/t5HdJUbXl8oSyoq
f0qpGGtmielkUiRA3X/TwxKgRCNm3+eBPoPsrRhP7+Z9JdnT3grsrwu+zbILzUoD
enFkRsSzn2oz/WKmS0mC7RyfkNvpt9Q0Mue2alBMmraiE+91SU5QcB+nTK7CPPYP
jdc/EGXSFnMryEVPMMQGS9HTGzwqzo9kvZ6v2op8orfTH6ZzUsApgpkFCEJdO5ZT
iyPTHk5PIb7+xzpYIs8LgeC5kI/olArFCOxbuB4oT6nrRxJ3yBouK/Pq40plgMnL
cOnqiI2K19ncG6EVdbLWFhRY0zMwEIqfh0tKN6pAuz6jWqbj7HWjDYLURZ9QxBSw
v7aHYM0UlAT1kIDzdWY3XViGrQuw3dGhx2m/sRH74yFyDMyCZ9DO7Gh5JHVrugka
mbMlcqboEPPrp00Fmgv5QDHBo2FtWRAhbxOApNrzdpG8Wui5/33pwx0Kba3yc2UE
N4El5xVRh+b1VnWXMwlVBfxP+Bl1qQXIXgQ+fhtTl5COd2BdrbAb9LnEoDLoyLaD
kow2lAwLc//KhDaFFP5cvpUPVJX7Vh5ycmue4aPA19Z8Mn9gujyH65FKtFQA12lB
k00cRyeTaZoOicXR3hGh1kKIaUTQRbcFCFFuV2OJde0Gvh1qEZHPcTI+nmED+6nh
Uvky6mcGyGhSkhKu658s3XzcSqg9MyYKdjFG/8H0SX6tlYQWgnftgsxo0yNMwvkO
1RNE17NG+V9/TGlAL7rRIdjTDqATHEnKlUfCimg1Yd4NXv5nQdDj8h/yUea6NAOF
fgiWhiZawGg0XIsvFXLWBiLhVqSclmJt8C5pXH9GhhuOUWowWmJWKPc5text05qh
VaupoGn+ZJrVwPV2cnJTAUQvXioUYjZS4jPhG3Gr1lH1rEWXyKM0w8L+57Ldv5Le
45qVcUZ/mvwjWtxPd7P7zi3HN8SMqqbS87urtyRceJ4SUwlphH3nlGqTlUFWulks
a7ivWX70nVadsdaiMeEp9YtUooHs0mb4k3ow069M76b8Bk5gU0ZCXpKh7SXiORAf
Rz3H7y1zYykrSMe++0gF1K1oG1XApJ4v/33x+swXZZGTGhFkzvNBTakfV2iKLS6x
+sHoIicquCZjsUBPulOrlVPw/ZlRmwghCMA14pjykivBsRoMkrh0/TFBJ8BDvA5w
3AeAdshxAg9AubWw0AR0Lsf8erPJWZA4Frx/B4GvmMO2vKjzaoVk/y3FIlxP5B67
29Lj91PkaaOaWemMNujfhY/VcdGajfI5XsKmY+tJHom2ODLauV6DUU1dRTbzGlWI
PfGAJVTVkGp/hPIPHtJA7D5jvyo2fdJTZBx2EO3vntaIllVw5eir37yW/wNBhqCK
`protect end_protected