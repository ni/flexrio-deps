`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4064 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1wB2ShNYedzmkmBWjqK4Mg3
8iDfXbv5M0vDNkp8sRs0MJn5uVuCCS78EpvYsGoFoQj0I6NwtHpFH8QNypeWXBHh
B1AAk2N02F0k7Sjj32nzthdswVd0cABqQTCChVJ3ImgmdUOPxQDF2Q2FIyutSODD
uwhXGrx6nOIpmPS8q8c4HFENe0ASjUkAyxCX6ijr7ed8ZdOCLiCEKf2YS0y3k5fl
8Bxj3pAo7yNGq0XVVkr7nuqXCM9F3ERx0ZBKfO6gLNc63iQZXFZ5YDfToNMTWBOU
Mb233Jy/yb4rb80bqTsQs0qTUCHYSB8ZPvJBEEii3D6FFnB8DyBR/CD1Kpobdobm
e0S8mEDx3iJ9ZDRe+Sylo3bZoOcVHlRaZl3w5P5yQkDTmzEUu+J+lJ/Nv5ilYXFz
kVtw8U41cUINWYIf44tWpYRSUSW/Y0JQZh5RlulwS+wUA70Q8EEgh0yrs5hnwE/H
TZmOAMhbvJuhSqy6J8GYSDudjQliMZKkJLwxksyh4fHmZkBhvlZ2ahFCHtviGnIV
cqabHFn180RFUU7AbTmxJCGhGCApqYKd+9hDp2PIVtIZWuH3AECxLMeZtzRr171s
qGVWGJhVEN8bEpwCvFOUbbdwrhTeJTJXrzkihCCbSk9bKaK1QZCbVyslTmUL+j28
qy3GaMpYFGW3NqeXPi3ii8W1Xamqi82wTmM+j+iPPyDZGc8CuyDhcYv/bY5SZo0o
UvtgMGIIILPWjVW1GShfTez53eDwp47ozMP2C3wLztfC0w2QqLD8JkBS08alSGOi
5C5BWP5EfvevbBJoji4A564WDK9yzmApBaSaBuvT/0KOOTpkKfcBtwpZDiWcd3yb
AxF4aJkflJYQXDZ8qxIK8TXM74uOdPdZNEZnRdyj8oNDt3Iqg7l21XFWoPp1knZB
+EqFW1Ow1FVjZbmUJ7FHqCMLeKZT47/Bf3IdE/XhrjE14Srl01svpueX0pkoWLMi
b9eKqp0KW3Zm2APfxERJjPq5rtdBZwfMt/OxxuroazuZ8ZlBOk1VSZUI/6ILUjBn
KTbPUH6hYKvW/0fbh0FLH6cwXVFQrb7N30yWFf+H/u7fTqEufEhqBut02OYVYGDy
0jMZ/z9qn4AzKmNAYW4E0pw+n5yHZBh8zi8Xnc85kCkXjJL7ACIC2jzEokBtNxP2
QxvlEoVO/+Avmy7VjIoeTLg64mXxbaR3Qgn8df5dzeYqmGjEAQKhDWIuSSnLfVLr
M7jwIkGxDlIqfMlX98+jWWHONuYjTDxfhEd7DbObSkFtIbfqrMdrRsDmuAZ7l0dd
gekQte4VGHO2RsiFxN+9dOB+H0XFqgSsXBcaMwq3bFgqkPXAkM4wMwKu5N3Pcwvs
4X7jJJ2ueg4ddKR3Ot5lkNxwn5HDgwvxPieWSpz068Xqa1DEe/SMipUyflXgLJcC
DkTg0NfwPjKh3YQOc2l+/+iNRLNyaNdR8NpQNDiYG2Jx/wm0poVs1ist6kTiqgSQ
k/0VHgW13FEIAE0ztjnAaB2jn+D6FgrY/GTyYLk7sej2zmPHICJWBTD533Tgnpyx
Rvn9pWQBdqDt1Y1JlZxWQHkwKhsCJpnAIMbpoWjpxrcA3ExafA2F+8vcZ/6fvLvV
yWlxCDvndoiVC0SDLwgVAaTJXQFT/AfgxOrjtgeY4WJFnzDnKXf0oiTsEdeh6JzA
yH5SUcPM+znK0Jt145dKaLORKyoKhXKllE/u5iQAwqr7tbMCDdWyQoSQHRUReWQ5
/3FCozxOP7gwXvDyqnuRCBBJMR9j0CV6A/3bjkj4pTXpIodug33sxEcaK2viZsiw
PMoK+2/5TmjfRiwW4QMi3QOmBEFUK9OvOekJRjxEs7p7oWZeis4oFxVSa2bmvLYg
mXWbbIgx/DYRgQrhD/JvFmhwRPZPOIkxQe7yJpQix4ARwTkZ2Zl0GYyhacRA/z0x
hdg+9wOO98eeXpdG/8AS8nKvM3AQHQvaYTu0tGEmRzzmLTPeWogerIUJYtdzxsNv
A0K7DKg+CFpGSe2TroCQfvAUq66yPY8OfSCjIhTpj+XkyukxDYu4BG96ly9W3+2Q
uRro7UM/O64C2g+b3ah8tMJX0R7BJh9EGc5gSKXbCgXi/8V4Q08JUblfqiIhrGch
JUNoK0fZ/BTO3rDrg3fTmpKyJAKYLVqVJO0/hJ2FNjKVOh9gDHQKzVwyFr/o6I6E
7B32k7SmbF4qcxULplL0NF81B3OKCFpL+rqFhWWKSzHbcRHmu2k5ZiUPfLjKCRbM
Yx6MnHDN0IouVMl6pRovurlaNXDkfBqGcQjJGZMS3PmZOdfmJHqrSOl2oL2iusVE
GUf7ZnrDvNCLdL6UTmY/Dihfk9fXWtaZPwSJmWQJtgup96Y5dh45cDfS2CtWSjVB
c6XML3jE8EUL2mDIblEsWbVN2hdpIyT+EqGscbXOxIpWlObbcc7eYWx2vHo/Bc6l
pxc67SLvQTFrL6yVzFWN8lEpKJyT+sLnvdF9ciLRS2nC2OVmCNcboYLwOq6ur+wy
g7bw1tNVlbMKRcTnIJFrkpLt6aJ7SQq+0NlhkY68/ZpqJLZa6QpnayJ2GIsmjKgZ
MBvCHyHTa1AoaxYPAyxHkGULZ4vbCJ+epuNgThFFGCrG5/SBFvkqCqzR+VrUdt61
keAjiNjVyeRe+NhhPEpCdajVh3jjpWDYCvH8SPAF81MlMx6cTLTCXKyI0wp9kgrv
JyJoc9Uhiv1E3ppQ+VAMgIMn1+7ywX1MYDovx4a06EnaWakIKGje2lVRMvp8bCYs
2whMV2SCZwsBb2InRhaPIFX2Yah7AnUHmHR9GLjOUW5FqVKBSJmBxCh5rk7HpETT
z981Jl/3+zq8rXQWdqeH1GyEEMl2oa6S0FrxXbKLhN1XTk+vyVJGSiWAR8OqOAt1
TT9QmEMbccKyK7udwUsNZzo6isUt02JBoLANjMULQlvYJvk15+S33SUA4WRahCEO
3Xjwn6BaXYIa2umQchHOAWbX+YbBID3oLzJ3O7ACNXD42ciAHa4TbGHht+pt/6fV
FLvf2mZPEEEqgnhnfSaGDvYhswolODav7y7FjhqosbpQ0965zBon9cr/olz1IJIQ
sKC/45x3lW04qbs+6oQUic1Za/pHZodAgzFIlzN47HJIVop6X//SbDHMZRQ1REby
Mo4P6wyjFOZWozXALkurVB/4WmA5YED6Af4AFQVYTBhZ00UpLgDb/bm39tdKpP3o
Jwou1qYkXwjI7v4sBxxi0gvKiqv+NCRYCFHf2SqGdYeurn7j/kh1liBNUwMND5CY
gASs9PaZ9KtC73q4HgBnSe+4OFe/8+jqT+O2kk3kZd0fnHFBWw4xAzDHDFvrOPb3
f9B0scq+/0S9u9ydYfXn6ihzRF8Mchdt6grItskpVItj3Qpk2MT4dl6zWVHulJu5
nQKKECSHIIDe4dhb1uT4upJYM9jyR4y8LSR+D2cdvFoWvw4qHBMOHvgPSwYMmbKN
z8tz/mBSGwKF1DZl1rwzGW7+vSu/WbsYUpWppuzMtIB11lVBQvmOMRHCaf6Y4xnm
ABByFIklvVkoYYT1pnWMr0cP6LMr9ykNnkM+oW2EOcZFD6Y3wx10KQfMwd4nhiSH
9nmfQEBRW9NI6UizIKX63/46envcq2OD5UAZmVmEXyOOlDDo9Aatpki6g4Nxztd7
iz7Y06ozf1EbFAbwxMw475wP8WnmBWontGpernJgUnSJHTqeSCsIGDnUEICWWF5s
4pnfLJI4lZ7a8BiZUWR0Mhr8AXzCSTYRxwQyWDtDfnchot4dm/ZQ5qNqNRZ4oBAk
G61cprOFfFya5TbDLVq1w0NbfbH0stTEyQnKuefWtOu+nAQ0of9xMHm/5DpbnwzA
q8+bL2SMpgPiax3JhvfkxPezIOzuFWSZ/LZcie5gMGeEw8Me9PhMKJ1NzY2iTfCS
Wg5cvETv8DGvubISv04D51my5gowWE9K+mztAA96OjZrXJmoFV1DC44xhb1+Zqz0
tnnVFYMx1juNTp2ZNl58PW+FSlmUDELGSd3KlL16LqnSmrmhAOuAiIxcowrjP5QK
1tfnZjgoqwcvsPZhTwvWLg7rOEDV6HVNjr6VOU7pwoSJ3H1FebXJPSKKPpcaBSm2
aTNNQscUIOa/p2RFlDnN/eKwOFZPwOisKgSKJr6qVbzMYV3Nk177lPs8914QM6gF
BFOp2xpHR+9hW+VRIz2lu20+d2oVkns4SZ7nT+Ope5QGc3Cjmgx/7oIzs1qfDlvz
ffSh3iYjugjPsgyF9yGSLXnCCjr/ha2joiOEHMa6CDzvuo/Y0PmrqxAUxeEM5HaT
9WVbTaR0EOXICW5sVm4U0tZPZULG7EznCOkZHxAZbQN2qvDFUeWM3qQShW7KfECE
9qyEj+MZ+oWBBmB5/qlaAhSntBUcSos1jP8gVbfgs7cFefagobxqiaoYBpkVmNTB
F1315dITWbccGJ0yKMufkxKl2Txfc3xDhNyJZjBIb7S3DBOe66Ghx9SGM0KtdPWa
34v1gqsn+FlVKvQZLgQO30bH4b9404Io8NwGGLmvbm9U7njgLzyB6p/48LSoKmI3
1RGUWhzSePOWTWvVj3Izh3zjP/PbBUxGedjfjGzJ3Qcc9YevtsnK5jcatJ/eYap2
7DCxb/Rlhv564WtQ4LzvXj7s/eh+Og77zroMgT+FIUGRarJIywRqJxCDnTg9B1XT
fBMdkVnE13AFUd8pmkF43D3PzOH+Nh6hxiIJQNC41cYKa/5iDvrA+/AMKg5ragHk
JPOYXC4GlEjOP83qrvdQbeywi6tiLoie1qtrDWzUtOnDgur+iio0zxpNaRdWlL+q
/vGXY5UGzoV0evjW4VcD1lxRi6JlHzCVoryqkk3phIJj/kv1xmaLc6Vqf126QEDt
X031948uEIRpIjs2WRSDwNFqFcW44JN+Nb9AK7QCYCRtW3sl0OZes73jyV6ddNdN
v1ouKyEfA84wWEgtRzbAPVyLHMzsG5QKJde9V+NzT7hSzSduBUab/y3TaPRvanHm
EaLfnKu4Fl8VWHuenoDGjuh1Hy0r04TfbUV1hpYpwZn8ZflFCRWVQ0cEPVME+sw0
5PvErDR6EHqfWlKvwSzEPWHS8t8OpMb9l+UzU9/fgOq1mySzDzxnAllVjzG3A5Pv
r80gH2cZQLZvKfK2eSB3UCzAQ8kpEEmRZN3YaZS7W6ULWT1StcsOimVkqzldNeOA
5/22D4Dc3Hq4PdgfRKRHP3diEnc9bGmMIjKQVoDVXzmJ4oKhOvnHBuxpjCJvOpI0
pklVfKVTi6kxeo6eSIUl5PvAR5dIxVqAIMQ+l0fCXKc=
`protect end_protected