`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
K1dgx65eVu6lpj9nEzu2xogy85+H13/M8k4NT7aQKerHb4DtN11h0rLZEeF9nyEz
jw6duha5ai4QsSxfvrIGwIicmDkKMUTqD5yn/4B5r0x+gmjPE1PBEYqY0zUrJ8ke
PIeF0VG6IGSIg1Tat43KQ6MU4ipLhWZIvhOBeX0Nze3Mf3KDI/knHu24Ly531/lx
zR3BwxiU4+NwVDugRIMSl87GI2EtfZc2mfFoDkHCTjb5cVsBzkaruAcpO2U4TE0h
GZSRUgpYA9YhU/dig4w8R2KgXfcpsNz5HJfJ4DURnodBVABy+XVY/Sy6BbB7NfBx
HLpRYIuCp8GxTnDQZqUSsvVgQye6iUZVPZgQN0raugFdFOo9T+3ptj/STs1UmQFB
wKtubgBzPVYH9JKMzKkxO1yeoomT8sU/Gkthm+M0iQIq9/n6Jb5uOkoTVJAh+YAN
sSXDr1R5kxA6J9+ADBUyFYoT+aY6Ix6zAWZ32c9RBDJO76+h2QKDT7AOvzCheuiN
dWdfINf+8Fzt4srWIP/CaXCTcIJ/BRy1Mamimhz2I14V/yVX+VQc+DI31SgibdWW
PTxetN8RRHxzQW2EGYL0AXdM0zV92X0BpnqsidpIjTVsv5JXxHTABEatwXGnbDLv
4UlIeDB+m2JWbvGEuKbh4+NhJB6MFOjsLuOteId2mS7g+Mq3JOILysFCzjbBFQoq
WvBzO1e+eoi0WOnlLvCKh8Vx+UzmzSa+V/s1BPJ/QvDumfk13wk6myj6Aw0gVWUu
pZJuxCC5/8T15GbI6qsM24V6gfpyGF6jWU1J7BsEC1jxIaTv65/hAYcoCQZqDHai
lmi4BEI4yu7BYVcqNZ0CZ5k2sQNxgZQ7QhHfoDag4VUP0jKsG3pIIwYmVJgmzSjY
RVFPCnVsTWovxKDzkrwAgCNzncT8wmHYA5HtYX3mw6Pez2QAxBaOxA+0C1LnMy7j
0ge2efwHPSDRY4KMNAQtCaokhINlyb+RXp8ZpiS5NEmELf85X3K2JuwwxQW41FeQ
3auHG+RkJmvi6LohvbZ4DVWixJKfbhDSclubFaq2bhK+rNbsLggN7DpkI40ohgim
iZkH1NgmCwsOZAHxFvcBhtEc2CmDzJa7hJznyyXDMKbL5Ygq8SoJOp1XXw6w4qfY
pin+2K3C73Qn4dZcmDOaGuywOlEyFz/TNuW7Q/Jsy3orBeGUngo97rICfcN0iyCK
u2KJzDciYogoGUeGd3zKQMQvCv+L/oDpl1EazRbbEPnghQ8Djter9qKGnBm1gmRh
RCHQSPbm9s4BySS6phl5lyYIriHTn0H4cjFzm19sY7dnWOgPXq7WF6QzulCHUtL8
fFcMVPmFsyRS825t5LYNlOcLY7i4RxP/zgRRwr4smdlQXs/4LUW/QsKMyIKkWiI8
CaTsPQoWIpGjRCApOcGvV+CxVCfyIYo944y7CLA1to/wXdtPlBZg2Nxnscjjtycm
abaGQ5dp8vr9zmaHVCxCG0yCuN14zV5jQ0rYUagccoN7+q7MdddLniojc8NIs1E1
LfXQiWDdFUwfE8D6Ev4AV/UhHPZzyY2m/fHPzUZODCv322Ku+FUJoW7a0zL7nwtY
mgmq/A9g3PY2oYfRwIOmK3xbqRBgTG2w00/EOBg9h8YIVMx3DkvxJHakm8McClB1
I7f3MLeVHYkS9r5BG7cWaS7GgU45+yU11Wlc8cDRDtSV0UKJR8Y8WMN/QlL6OXM1
UWaaTQ6OELoURURGpG+U9qrH8ObWPA6miulfgHenGBnrUKvxzBbXYGWehBFf7WTa
5OeZONqn6v/223qVDEVH8y+1ne6f0hcUJ7t7GwuEQcjcCvkmJtr3j0XOLZrNZmhN
ofuCOgsdFCUDvL9g5Ld3dml8GwR9EQRS03n/zf4mZBlHKuLeO/e/c5DiXiqL5Q/5
hQ0hKl/F/daDSppgID7aUE0it0jIbI6YQdaCXi/2ofxT/8ICNQHSzJ3pQamIfGyI
w0V5BhvptJWE9TEac5OA2US3lKcgrFZPJykbwrRfRoM/hglkZy99VgzIxrKIJ2Wa
2mNR33qUmnZYjbR46WznUGzplIIrHUGmTQ6AOhlFd4p7WZDIrfK4Gy6tfn6kpDts
LE/+nWX9NjE0bn51f9ZLPKonJK0kwT4UUiZkXe1+yG6c8OAvAP3o7MU6t0sSZKgL
54FU5fpfhDk4yD5bNLUdY4sOOu4xKiG/1e9e2tCZKqWZi7nfKYAo6Fm1HHO9QONR
sLeoDbzTy4peY4hf4l6HHP12sh/gdv5phUEt1Cj0SdKZRDq84peHOZ2Kp2l96+H1
+3o0co+Se+6hajfUx/igLUic7bxkNB250wVvh9owIn5US0howLYzmv6iwudQsqT+
2BqoNAjwbm182fzkvY7dHb99YfYwivoCRGNwQQEl8UV30ezv0foeP/Sbk1rUZmc6
LKuHhMSiX87Dut2/LnBZlGGnuOGv9RpzrnUdzq7EQzYTKZj0hercrksF2+ilCXeZ
JBuDpOXgz7KoxBRpvk3B281qsVW0qjmaLoRmO6bMZYXEmPDV2tsY+ZsXa1W15s0y
syP+EldRLeERP3ZZ2nlTOK0WsgOhaPa+XdnaOqNiE6N0CP2hdLYQ7iTTHz3qVIzW
nwZXvAa1f9nAfFxKSrUeI/WveaDq69vobREUTQdvP7zSh+d4KvsWfAC7DMIQRXVP
7J426NGOeykKImY7oFJWcFL4BpE7UxctJpGHKnI4OshnEYhieYr9VghugW2kpSIT
7P0iSVYnBUbWHj6B27NSF65dqXQlXf2qga9lXHC6+Wj2UVVseR1j4aFQ4akXIHyg
f3nOiGf1oY5920jfHSUQ1tv9PPb48SSUVS6IcHX5K7DgDFHxp1iIyjGVOR9KbB4u
RAYggpMUUvRvOtTloy6BvkTVzPf2eLFRNHn0/fTDzNZfGYl3yLfdMRHfHWk+T+FL
ywd1nX3aBBncw/Nw79RiB8ZV+HM7pQxKOaqOLVju4I6xW62hsjTi6/e5WqoZrhUB
PQZKzOz6T3R0SmKDvpFME7N2Z4nKNO3naXK40Tg1Y7y9Gr4TjKaYPRCZy8leO6R7
LoYuWDj6A+yS45ObeMY9+muuFn0Jiib/KD2Knd36TJRECiTXaEBLTW4/e2FoTcDS
XWqrvpTggTTljXO2K8e2jVPSBjp1A9leB7ZSzsohcKWtXYH0E4iAhlrh2XnylrDp
IJqDVQ4X9P02egT0u7MUAaZKpXViN6mlAxCYO6Bjivjts8EZUHlqhb6m/vueLwby
hNHRvECyN0iO2RIlnKluV6cWTEROCqllCWbhuFSXwdFKrQfdPTBg9bUBHf0fcCD5
DJFIb6udUDOnpfdXM55F2QKyNU1jmkGfQvRe1WYO51aGZGsr3u9PUTGA8o4DxWpz
682cRvpTN1NO5F9LMEL4kpmfG/EaLaqNHl4833y78vEYcl0wnllNw/LMFE4xKt4k
WrMIc6Pyjju7T4PM8hauHmR83KEcBJEHpYZlz8FBke1TPR1Kpo2WQlEJJcDKT+20
usK2LdEFFJA+oKxVkNk3KVUKU3PBMs8h8THcJvnA+T7hKbzQQIywHApjAmHdi7+7
iALjIvmCCdcwwQy+h/S4FjEdo/J53jsTCKaDf07U4Eu3R9XdQd+TOlUvxH0JDJro
dy8XkS0sfidFEoigVAtZUmFEvT4X/Dqlz6WglRUW2xB8v4FJT45ZCzyZv4mYmsxw
uLygATsJ58SamlqoY/nBKv7y6NKVCO35VqOWqPJyLEs5BT69pFysVn5rzgu6Ca2f
W7ElSWl5Ffm0BC7yiwlfleUrGdYjsWJjK0VrEsR4iebAq3NZobLP8hnwRaPEuJyw
n5a9WhVdmsjfjP8wr5VEyhMGw9erkNzYT6PpRKC0++k7AcESQtgXbXtGHFemmSy7
hegH8mDJp6BoLlLr1wNlzfM4NozsJgkuE+S0wZesqlQecSy3ciKWTgjEI1gL5L5h
AgWhO9DQ+4NC7Da+zdwTvgS+QvtoW7wxZeWJSk11UR31+iHXG0nZqhZtpHj1WJ8q
ZBKdl45GF9mP4SnSu1FQPqxlNpn/B1VD/AEC2ReRGh+qUznSJ+af03JedONL86Yl
+8N2TgpWwSiY6o1etPp4/nYBRxHKKFr55xkYEYdchb+KxKby/maNVXV8ziR1jIKt
Bb1jj3VNOgqlMCklkTG0Q0MHLRt+IB/bDCmzpPji19ciz+cH3TFFlqt51gMyC985
8dSLYwDbYvVntoxnu9oAMLrk98MeOjLKY5v9e6p7vtji4RN2a6rukRIv18+yWCb5
2O1UIce1sVd6SM//4NaEV0nswfscAQx+36wXGgfvzs3pWqP5KLtUvVqLPSYGRoOt
FolBwvUKyjGbQiWihKhvBFfaR+LB5AfEny23CCwbTx/Gr7Vb8lPoCj1AsUCOOgVh
AkYV+z4FiscIzFFCJeguIbYuRiTw0mMLzfZOu72HRHs6IojoZP0lpkRCAWSozn/n
kmcCbwusb01bpssaXMIOR5i2AxS7qhJo73JRz3f6McR7vcDcm3bZjmzejyMJZYJk
Fj/lJGjGYmuin5S3JiyYJRtLnNe5AD7A+MWGntvWFLUWEQzQjTM5QN2t9qNF4mqQ
qAaZSBlYZ/2m6Cu83nzd+6rlJne3Uof1KwSbdzr05Hkmg0Yf6D8KGvecA2yUcpxD
iUWhQP6hDNPzQ4sCnbTPCuDZ4eleoA1S5IygtM8ue4Jb6SvACvT3JQIhOor6sSOD
WuLuDhmdQqw19f7zZxmCWCpGGtPFHnFC8bWE4ZKtFszdB789zssJjs33v2qMWE4X
G+H0Qc7Cmoo48/YWEh+IZobZkQaSswrVS2VNa7wwCEGbqDWibabKiFQB7Qi6KibU
GtFyJWv4hF+VWT8MPOT/RF3vykQuRNuvkvi3ND9Clqp+j6ES69fWgN11ECKAuAmm
i8FYiY0NANtxyGeOEs2SM9Fs6qgLl7HLa5Dx+cAHFYjMfpvjmXwT4X9qGq/CmHTf
Tf4XyI/lJCtdcBKDIzBBrYIFcqn+j6ce5qirK2SVgogmUl8wIZEbxIudMngUFJm1
JbZ6kbVvqKaA7egpkJdNytW+OjcJImO0Ulbmxv0PjdXEcxY0X599An8cB/G4f9rp
OCe97aD9MO4H7shD5Kkyx+gvCv9Jeiz6tubED8zpx2SgkDti5l2gWPK6n9ifIZVQ
XvBP259xrAxiEHTccs9hporQ2wlmtHM26N93zazsUi/rt8vAlXYK/XZSOREG5n0S
iB6a3IjZQrJwfD8sdBDpfEmqwerBWB/NqQEmUS0inwLSmjRM5JTWe8or7LH57rwl
uT3s3xlbIu90+Ok9HHZG5OZf1+0WzLUcJLvjo29BtgkDcviwUEhnOiblhU1p2HWs
4xeRuzcYRT3DdSgdW6OP13+CM4YfhYE6PTabNuc+IWBD2L9/zZuqDy5zSs5CohVG
WCFVpRQQR5VFADGVF36WTsDqH2vreqXao92p5M8Eeey+fLk1zLrucWe5wPc/C0B2
cJ162QsvhIfAy+uHTZtCaX2J2kW//twRqLpryb79N9dH4aorI5iq87J2uyUd6NPD
xaTN9H1LatbVe/d3UlyYuNBQkTrM+UrsLY+Zz2WtbEuU/+tYGPJIMm4SKGqIg2Lz
tOoS03djUNdJo25zeTArv+S9fA/X4y6f+cIoygMSlmv+y3vyYlSRbCm+/z9DokD+
jo6hbEPs+DCqycqFnGPt/DWV1r/ImqzeapLxuD6aX/6LkXRpkBwnLH4bvKzQUVS/
qlNwN0wtY9ZWYrGXhsfnqXmkrYFhdWz8gray6tXF1WFw+3ciewk7PxEdrZRSryWU
n/laPsQAAJJ+x/Ky7L0pj5plsnc9G0XRTjIF7PUQowHLch6IOkxHxuFL5hQcWdS8
ehVS9nUk8a+Zy9RndXOiW7QtdRONoN7SnOfdzdNj+MAT9oXpzbg6yZCjqEF9Y1un
7rBEp9f+L6hTAvvDeg0tphf70cSMTHKt2uHmRBTRvY4g6JBjNCWJqZQfhdQYVKL7
+j72yjVvjd8e7HRcytZFlGfAOXid9X/Oq/olHnad8NjR55NQtFugNnjTQf+AfsxT
aHFZE4BQYPoylaejD2Bbg8FqKqk/Xn8OGTWzhTqCrrAXzen/lgL/IpEAme+7cau3
kbG1P/WP0PzBChX6lZSdMJ5v1bTuJL2OQ5MUblsWTACIW3ZZ8aAuxQqCWV6TtPzp
F/7GMC8lc+BPTHoOvCRkhJdxuTq24PQGLMpvyX1RuYqOTiQONv3ELNVvf9sBrkdR
ScSOzLL4sX8/dZyMDgpOhX0nH/iHnxnKLJ8MqWMhgKdVlJW7iYjx+XDCJEBAPn/E
0ulNxrCY0nBruAkI7jVri+u8UhVoCd6HVuEYugYxim1fRKuUjhEYA4Vyaqv0kLtU
mZjB1IIpeCo6MJMB3pmATFvFyLnkcxGtCbCJMkZzbJXOI4gLPA/NcumOqmfDS6vd
YQy2YQvezmBi3llQsX4hbq9MExsehukhOAKj4Y1CVzDiguIE0evLDKTWdlwz3S8o
zhYG+uUGIGQAhJD0afZGka+XqRfrxiJtNG7Jq+oI2GQoq2M/DWt+0pN/aWKxAAxO
TtSKMaZd7CE2L/nXu8AnWPrEjnMOouLdII3RMN7fLGGt4zepHgei81XrlAbIra1u
3NWI/uTo0olUfisyqw29odXLgdT9FQmlYm1LLM8AErYKssSnkb8/87MtVTWSySDN
eusaC8KDXqR8OcKYneYr4HGS/xzfMaofYatxczz5IIHfwWwOfBlFf7BErcQTudS6
DrmvexqXlvxH0+5mNIN0mu9xTZ6dlYfhbdWwp4kDmEjzqsfDTwNKwvncWkGWdD9j
sJrGSS1prPx6Dln8LtNoej2ksb+mVKxqQrxqKkSipMGj+Cw9/RANZ2I/YCG6Voae
LV8NoBrQc6Bj+SQ0UAd8s8WL6TaNeputJDawP811YCwBeelA3kxPgXgJ0BVNNl6Y
4LtHdkrIjpi7pcDcK2MnKBauhVMHevWJDMUNE0QYiyYe8KhFm2oHE7s0GNEoPRN0
qTsPp2QbSAvAy6IdCFBIimJs2Mgf3MF0iLhcp+kAQz0YizpqCVl+NYtl1mO8PHyL
dvLy+xVb3U+ygGUXxmd5XUzrfTgMSWEI1drcr7NVihZsnsBn3upWjQaje/IcC1wL
w2e9+Gy5BgxKt8zvp9Jyvy45znU/m6OhHvV68NXGSE0NpPjYi1rLpD1RXYcaegQz
1rsnred+PPgiy4lDpOecN4wuh6e8k45ySYcWjEEQymMoK8rG425hUkOmdV+KyZhT
Svefwgstr5eptewB8Ryfs18Szijr1hajp1N61SpKBr8H7CInfayPQF8a57PupEMq
UvyQ3LAt/PWJsCwSmcLiEu81nqtBFw8quwtjJBqhQ16ku3sNuMDFDw6r/xKF5vHj
tygrZn63Zg3t89gnj8xqice38uNzipDhA3vMjdtEf/8dxYjJZeGU6nriUyV0IjoI
fTD7uX8GyXbFO8T3nkkHeZlkjaUZ79hkAV3mN7LRARqic6Bp3cW3ZfMtOQ2iuJFl
LuIA9iigmdBPy7OYuYyLuz1D6Jf7C4PpdEp4Rk7s0+pQSUd0ebz8f0oJphkBnuN8
arxVtNOLhRoa/pX3FpBZ7pIpOwGq/HUOt7xCEadNbDpHgeUF5SCdpsJnMAs2nGs5
9mJUIVhjstouoHOqnLPCIRgMmKXVtsK3FLRuz5+FRquJSFjzMP7aDl6QEWfmhoxK
ql5dxi3D2ZUJz412DAWUprOPBETIl5RD3usje+KDlqU6h6dvt3Y8SC8mQn34c8GR
ncDtRExfS6VYV/27SO4az8EkAuvZDgi+n5NYGmTaOXoWZA7WjNwYsqzQO1fqCXxU
Y6SGo1jkXEHeaOsWUt4NHP/y5Imarh/BYpB9xyz9l9tXHyXMLv22K1VgDPP0wQt7
AonPwFQDcnKeAy9RoF9PFg2n6UZ8eQDKXTUKulfdBpj8f2QmNZV0yq6++X2Ic7EX
mhAuljRg+ti3uN+i3h+IHLJhwfZKVQiuOSQTQLi711Q5b2o2tRbASyonSLAMOtxO
rSw8B6jTzkhOCOuu5AjmYHmw6nGvlCfzlSGq9XYE68CRt3cwufiglBA7QuWvF14i
0GG3OMJIrnom6cPtqF3jyAurZoVwUK5Lbf2UcH7+axu+uoi6ExODggjsDBHYROu1
BVCc0gpL6+y6Ci54Ra9RQ76kDPy/P7bIq0+NcurMKl7jW1XTX0SuafH8p9o6YEd3
NWbR89MpsNHl1uB0xqgyhC29cUkwEQ6jvH5kZh9popdJe+h1+CDS2N/ZeNahQyzm
15KcHFoAj31HSfNaXGQ0e2SOdcXOoIoURo+QnFNVR6GN1KEXZRDIeCv0MYXpVEsl
0cx/nzC5o5/YzbVd+DOv48aXIQ+ndgLnksmp2J8J54UYgesP+aQqVg5xRaCpTkZE
8SG2BCYwkrvbu9XCgs/uywd86PMfLqbM6sVlOIocuoRIW6oxP+Mz+q4IJ/gVqEQn
pKlbIuclJ9i/c75WqkzB2AjdTE+DmiHlJO5YJag0kwJgLvwHhuOn/Dhj1zSKRXBe
UnwAcXJ6kU+MpfXt3EfEOIfFDFqlHOvaSs9X2VAUuxvlmf+KNyh1G6w6F5u3eTwe
3UXmDm2jb+GPA/FJB0y/p4dvyWt7+4TSmBqtR4FvMVLmth6jIke5Z8IeF1hwxWID
0Yt2tRR7p7uyuxGtxHqZ8lup14T8DFdKya0xirhwANIgx15EtL1P81v5+d8aOxfs
HLQGjaQ2XHjoWjxU+gShtE5TXI99JBbGxz2Es8I7Ur+IMdLtvPv31FHizKm7M1uX
25PRGrFHiGsDOJ6TeQtL7JT+9fLeJjlSCY0cB1TdVVADOBctNDmhwfCO7XiP1sSu
s/CfyICXqJhZ/Ir5cTJQbhNqmwUuHs3XAsJO4bTXfGcWqL/ebhTcLSdbaK2C5q/h
h5XsdA5a7lgo+rAJ0NK1ALK05gVQds029dJOmsLrARcpAV4quL+bDL2xnWyA7iHB
/0plZMZ1EM24e5FkrpJXw/nhvA2CjGolZe61++pfTZxAP0/S4fnhpTtsxri5wf6T
W37GhGM2BYPhmer0RN6Q45kyCOlt9/1I3nCXh5GBcZ4W8fTWMCNrFrkPCxhhPGHf
uDW1DBf4M0paCgvk3fXuOF4LMikzOiZFJXjDcZ42jTL3KEtPgeNVJIRlbtgurHE9
9JhBFwnm69IktJyZfva8pZ9J2T1FkhPplOlbRi8fAWhYu+vP0VaCkP0VinJla8OG
w6JwXVR2Pmo/Dh1juCYXR3HTBXTduUYG1tltf9h7rF8xaXxKHR+I1cn7sKj9gBXx
2fkS7/tdaj90si+PTVw6qgjHLGyvpXim4T4qr1Em774SKHtvmqLxXOv1PWmLG0FR
nWLOCiJi0x1LSIZabnHSfrIKgTRHKkHKWkRbBP+d9Kg3GI2rlXrxvkSk5h+tcmxx
hozRDSlYUz2z3FXU3AhMfimKqmFXXyWAeGVv2l1C5lhCOrP5VeiiWmfJDeUw7NmY
0FKeY4izVkApPPTmnI2MDd5gX09Wg0m/BwKpXcVkYyeFeaObe4q0pegEpa6Ogxmy
exeTjGHd5uaXVF7Py0E+N0q5LHRjx2qDbeoCD1368XeIPEuiTwZlOWnH6Pxt8vUh
zPeEq6zOKTFfQ/ozuL15FFW647EcKGR224ZhGn2JKCrCLtkgxp637hT/gDfZrcvx
WWkGk9MT4r1R3N5Gtfept6hETYsOtoNZhU/0/iSOU9NN+s2tU138JJJ7ZYOJ9L6Q
qswwvMjwiMQjgLUG25XvU9qe453ny0a4bRcvEpgfQt5K3gX+6WBoxUIOUW4YTO/4
nZptW+ji/v9Ij6RJ+5pVV97tOd6ap/bDpqqyzNYTG+s0uONBFN7twJiwTQx79J/e
DWxYlOK2nsGAhlEkB/kZdfa2bERqt2e7dqTugjz5cl7yfBy2NA1WBZbczwAE47nI
/OWMEDdTrVXa0Rpd2mEG4vGQFaedcE8ScrfwlaF4aJ9oNtNItmIVRkloRswCzO2b
ZeJkV0myjpMHsRv/1tLQ6bsaGm51Ftkt3cix5cJVcYxvZS5u9BDzWIlxv4UP+Hsl
OLkAPEDUCpN8oTNhZ/mBPGKlCHmvRQwUFhsckXdxeMlZMrkyX2aiSR9tpif/DuD8
sY7/KQ6ax4pkugAZPrVkYYqf5tpxY7wb3PTzb7UqEUsTr0oueXeAeAOBs5DvvIT/
zE0yXhdJmKSJcx7YZu/9A5JLqrR+fs1BWd991c/M6SbSKnhyO0L07P3a8zhEOraj
KdkiSy69WeZOb2Qc501lsjIVTGKaIWMoiw1uxqiVW7ie6tZgPpT6hDDhOsuqFRZX
GR7xOjZsECA2S8bYsUgZEwyC4m2F6zJJvKV4l3ZB2lBWBRXXIYS6mL2YHLBagy+d
0QMIvrLr2+0oGhL8xe2kHn7E+w8LaSmsEHO0pPcbg3itJqFJaLxVrIxV1DkdsiHF
W/0Rbkr3aYezCu1FCJEOSGOnZ0F6zdvZSGJR0uOuOonL0RvTQ7cug5GWlHY68Mep
xb2ZjPlV/2BW+ZJxPcWIaF+9lLNcOqeE4T7Hb0FTsVNkXWahLGB4fLufol7+gDNQ
N6BgYvoISP6Y/kIXuFY8+54rImAeOGHjwbCqpL76vX0tXazJIHFESmF33wOoSNLp
zO6vItHOphFiDVQf4d8dvnG79TbkXGIVo9QdKb2A3pBnHI5t7Gsy5rLSWGBbI+UT
YWP+JFE0u1ga0g3zbt5Ik4jm0y0bHLZkGssFdPnx5Ata/1Uhr1gxjO7JanZtOv7t
Kpe7OcHoLVEYOjp/LftjAQWLK1RXiY/TMkF+lCIZNDzL8Q1RyVKPfiO71wT/Sec6
hjMiIY0exzLm2/r+8SpqdLP/uVWK/P2BxxYCC8rrL+N+q7RyfP30uwureg3xG0JB
4ia+F6rQTUiRIhBHYX03Agq74nA6JPXwD5+wwthiue8YWU0G7VElBgWIHXikGeqh
2UdDO51Zr9T3agJeCRlF1GG01L54muvhSUgWEMmN73pK5HqVwMzFDE8reHdL5Hb0
vKq0iLfu2m5tRpjw++kjvvHQ0D0PLeGLSknIdEe31rkC0J0f5DTFpUO9H0/5cqVp
3AYlDpgYS31y5NVfqYY4DuKsq9Pm12TehFx5eEAYT9JP/vRx+5Io8iezhyCJ486E
T1hNJ97jZemiMyr/U3WusnWpg7OSTEhXLBn7y4NTu+Pm6NCEGgavLaf4UI9ILuGk
+RReKIZ64GApQx3SpkRH1cG+dRL1G8XIouqKgRIg4iHzxc54vT3O6XjNLOk5g1Zk
D/GaCnMWTvgWnsvLRUP3WvmFDBogCorpjxsXePqE+1lE34UOABz68TOfwSFANNlb
bvtnZljW1TXrwEQRs1FKT6FH/PP0SEN9wSkTquwvgOMs4mDJ05T3e3KNzPZvin7C
R72g8/aVFhSDc0oIDS7KzJwH62xqpQlaMcqMbsnzjoH7EuAvJUHYTqzD6M740Rjq
LCIWO1k8jTnahncfMJObxyU+YCHtBiP2Ep80DJsGnR1aSMjk2GDs7fZjAPnrq7Xs
4n63iLoKdyeA6867/RduXpEB4xoofLJoUQxWRTJV/N3/aU3C6UH8j5tCjVxHqDxj
qYHQz9C2opbSOzxMJlUP7Aie7iGhCBMWI8PwHkL9P4zN/xK2KyJuRAgqlUnWMXbx
nitjckoxn4kZENqDdc59E7tNsEoEUGMJPX+HLNx3Zrn7kiKmqT8kPvbdr/reOyAH
rrCYtf1E5OUQOah+Fb9K3Rz8h6MqeeoRwO4rU+Q3/DWgS2DUIPNwbm7Gc80J21XO
xV81SMIAbxQvPZYqGSopPKdSH4+SYICTv5ZV7Gmv//HfYvWl+knRjadLxoLT7qcv
+fltxAYe1jZNLj5QR0+NYsrdoNjdd3qLqgUJY1lkQpPiPnqeDT7FVIuSY/RU8YJt
NOBaQS+z/v7q7jJ1P6cJxzev2cHJe9n3isxmJ95RRaEl+9tcy7vSr2CaSoXOG18B
/o/VsJXZrPdT2D2I+7d2hR0E28NOT3J6NGhxLm3L82xG50SXBOEcK9OJNC+GsrmR
MxUFsxj7unvwtdvUBuD22joXeo4OHQu46PF+2fZr57uU4C8ETkP0Y79HlhEjpZ8k
jbkC0HzS7wrLZNrj8AqK0+iZz9vmvzVlLZlC3TLpcOUvUFeojW8hyCW+JGqhEDA3
sAJJz4l7yrAtNvEfu8KGNg76uKXyjrDS4woklojdu+f0bR7w6W0mP6xuzQfwd49k
vJI2LD0aARxzuDPZX75HkY+fO5Xocu7sQVuOsPnVBAz9y1cw5W1hgDP5p74DXqfx
tO4Sh7G3fOo7YSaFP+6IeLm8/bvqqNtCgmfpO618GvHj2Oydapmeu+JwylCrL5k8
5du59N3X2+AnF22lYQ2ccZCPwBvLtFilj/mJPMcOQwQZFcJo8BJaVLZjCgfNEJmJ
boOGEkoG5cJI+JS8CsIHD86V1U/QN+1o0lEqa/imAgNXe64Zm5celNxhDobn9CC0
+sZFXhuVJ1jczzy/MKVx8ShGXwTRTicXyPUqrEa8HKda+cQrGuzhyR3w5tMeTUwX
eGn+2OY2GSFe8GxH9lsLlB8VXNudEpZzWUVRAIu42P8azYKVOdWc9RNbNU6PIAgz
RoojpYdCAif0B77/QgtXyikoX/mCRR/HvdBuPwDixHGCTEPR/eyeGMbXNu7ufnx+
hrIhsQ+ep0pgDlnKONx7QS7cFGAS+2tBXvgADQtrwbmMZAPVIbti17TDWVYJjnlH
X9tajI0eu5UbjBGjAvuM05IpuYRQV5qIn1dVDV4bE6O2+JYAxfizeclS4FzwQyzw
lr+DhCKGP1NGnUeL8ecMKK7TQso6rhs4hGZHFvGY4N2ferjLvmLWqjx0WlE+3Cge
G3fflyY6/CM6No1JTP70uBeCqZkehR0sWQF5dIagZcIIq1VBMGjLarrWVtxAwjMQ
hxWk7uDZNNgO7n2qJfuovlFx9lG8rJ16vH8TbMEGRVg+IaHRSL3ZCDGkZ0FmgTgO
Vqb19DGr33nKN/hXUBp5pmfqfvHMtgcE63znVAp7rBWG0LLx+jWXApy/2Mvd9Qan
P+4jAHezkmjfW0KFdYmodcdVXwKmdPk5bQF3U2z3GsRrLu/lKIFyjq9nb0Fseebw
VpdVaWED4ME2+K7ea95PAd1AIpNSN5W+Y675DvfO1YTijZrNBj1+YDg+20L7M9AM
Vctc6GD57RJ7wF83i+IFqMDkUaDPNmac1LLpnWTHELMmFWYQxcikINmzi2RDUbgw
nfIaIngZQeX4G8yWNm7BWZ+1jNCCv6CyiM+9UruHqkEPspAGBdV1Z//wY7SRsSJt
RzEj+Tgh6iWlkJAqjGYIabpIa+qR1IxIYFoDiSvVS3+QPO5Ljb5RIOilHMW3ZvRh
NXo+2us9NSrV5DrYb3RjEJjo4zWEAE3lWk8iCgn6k5FmYZASCsyrXYHLqn0zwayX
adx0rcKZu1NLir1git6Xbz/NhdTzyHJeDKxvfM2NYoxzGgapAgGXP2Y3/K9Ukhuh
fJqq8L+SQHVKZXPhqtk+BGoYCfX7/FAvV6gVOHnRZA5ocstPmAzOkxjOGJIX/ctx
YgqmpLnitVHVWdPBed9VVv3y6Q1qFXCa6fZRJK7WARsySZ3nJ/G4Y7D5B70xfpjD
30dU4Rw1a9rF5+GQRIrzw68b7VNJYY7rgZwq67ZSBORbuNGikOlOHd2n0x10WgtE
uhJ1cHUZSZcb4jeOXrvr9rFXq9dYqqG3B5D6q9MMaiS45BGdDD79t/IBCpHInG3+
eB+DEXPjG+g+DvLQ4BukJH3Z/mxoKhJq5DW0R2idNL+ogXSYhyZ75UYslJzzK0o1
uY5i/iiWGU4woj59m15dXBA3aEN2jxBM2w0doyWaZ99ZN45rZ6B54d05FcT22JGa
yeXT8v0SEY2SzEl88CM42cYgi+GV6xpj/pAzkMQ2jN5eMKO7tJA4XQmawE90p+RR
7YUHF+WhoP+hdGEH0jDdHfCBlmNAwVTvn+Mf8E11/98H60Y0NSTSGutc+5STWOQM
8pIUow1nOFSafRLCWOJ2s1dG+0cswIGaNrxU+X4knCdgdxcD5fkwSu2L4nacQtLu
X2F096Yek2BIEoL1ZCW+toiKpMzNBxs+O3SXIId5mIY5p/VvdeqGht+/nhBIqITR
4442hW76YBiad5fDFlVRmMjy0eiOid8IPDL1635Y1fYWRRPMuCYuyD0rtYad0nqf
A0E96K6+R+AtKyGbyaJx59l4GzGHY/6IyfWQDFmo3p5sL8DUFS6tpJau89Flo72W
1qQA+3UgPILVqsv3rUdiDr0wN96kV8T+4BrSRgHiMno7qan5DuaG59g8OnpBBOgq
mO8wtYTw41zF5QfdtK2Gdt+VVZmt07xE6NkvPCSE4At9IVOSxgAxBrUswijaqM42
AaxEmGzw4vniOENMcCJnvu1FcXznebl8YkIe2agvyrBkVYf0SIdXhz0okq+g6C8F
5Mp5b4ciOWdszpunVfMbNSiScGwnBackedHX0gPefu+aNCYEKftXNmr0B1g3MWK2
xvRBKz+0uKv/D1GhcFEv3jOj5Tq6CWT+sr7Mub4cSyIwQLR5iDqW43/UH3j1+ghv
jywQyNdIzPNTLJ4R7fihjlFqlKkm0wi+myHC/0mMm8ItYioaBQYMDhxfLBE6vV/9
DHLLHEa+7CzKXHePp3mIWyveWjRXpDL7jbSfHNbDW0G56RvQMApu6ylV6OBqhO1I
nL5ws0SU4jzJIMe9rTKVUUh28X/h2n4hMUouRBpElzCcIge7WFgAGTcu7sOYfpDx
gpvqZEhpE8+Gyiy6Vr2JK5EFPCEtRwrFaMCF2UpHo6Iw498A24NuMhYcFd5ok4Ha
Vjdxs6qG7nXjmn+z4NykLs5p27/34XpWA88wSG+QzM0uzoTH3JhFuHSHmpPyujAR
JDL8oXdDJdQt86GiNyWq7SyTLz3tCMF2gvm6906fNQ7bmoNyUt/VhRvotQksJdfj
j97BcwRM6Ow1pjphgDyCumkvBQC89xnHlI/Q0fNxJrT3fwYwwSVKt//wtaQgI+ww
KCo0BmIvmFCpVNk7zSnDcMV79rEBsC42YMcrjGrV81wa+8jH/vNsBDTuElcUxrG3
N29+p1CP73NU/ZfWszh7IMsX9Cf/ypomULn1W6Yzla1ejBQm0PGZXEnk8uXOKbhB
rZdA+frFwPR/oEQfNXye9Qsj4xlVlnPgn8t9NI1fktGGvw20NxH6rrI8JVZPUEE/
/37dBybfrZeiqBCe6Feu7R9m2fajitALxDfnFbUgm1BN0SrGjIoU/78uG/ajL3Mk
uvF+4VM7EKkQtY5bv1Rfz547FKRRPvHsdqZlglwfFiAhtqvIKe0qJAP4S+qdUDEb
kxLm2Mdo/5bFfaG/CdJ/14NJm4xE7Y8lLw1xL6lvdGgqp4LtuaSenrVnW2F75jhS
bJ3T73mATqSB3SXPjJsU+B+BDCiYE3G6uS6VC99lkMrP2z4xIAWo8VK7mrRlarpQ
spaXDHhIVso30y0jYFXATV9JxBYGPvlpgzgVB1fb83X8kLr26+vti0x0eijSOxpA
IBtIni0zb5YGvgVzGs0b8y3HN83EbN5MZWUmYbDpujsiRsg00AaoP50WuFo8au8i
DVTLUQoBCCv7sSFlNDZmKT/scKnq0VECLM4sr6jw/A3UdOJDZZnsUFNW8gyW2+7i
3mB8YPuSMGhjwEfi9poyyp5GoMnIoshrRDCJYUcEoNMBlQsKoeyatXf0lkhDTUzs
Ia87daPAzUbw2PZoKHJrIr3BemBdoCFM+WCym4fgKp2EtACkHMFe+l/zZc+I50of
Y1BB0EuKLi3+kPoqFXZeVIliN+B2VA7PQh7UTlMCgPxXLa8xZm2vTuDCA1+wKpML
zkANF9+t5HknOcvz6SznybZEtekTKFWuuMtlhMaKo+7L+Yilnihk8KGF0/glx3HJ
9qKrcJd2KmmR5dnjaLDeePIcvP/T8gikRABwf9I1GheXf9F7SG4Cx205nPYaYdxB
ZKdaKuuyq0QbBteQjYmL80ZzNEHjuUzGj5m3SEGQmq9xzHXoMptOnvqUN63PRano
B4WpMIAAo2/QOpqRuD6BMjkWVmLw+GPITpLgLAW3qABhkJ3zv160Ny733tuHBWyq
o0b6tfSe9t6RLlW9PTEfGHqT/neUWC5AqPRUlqgRuCroXZOXSXeMTuf16a1CDRkj
IyYSmpHvB8Mn07pHI6ROVcKMOguS4d+F+0E7DOpz9c97a6w74y40Nz6hQ8/doytZ
+kSp3XGkgAJ+LJ203kNT94I9865UJC+89/lSd2JJMpv6aM+mpiTEpnasJtV7z1MI
cRlNnElB06Knh9SmUMpxPP843lP3gCzY1GLjlZKw+Xo6tIcXp8IJfe546oCvXFHX
0U2dD1pM4EECrlupDi+AODU7VC9ixi182/YRbZgFGG61rSQ2DMArEii5xjPheY7U
RizpndTRAMrekbVw8BYp8ysgp+quzKHHc5fWP2HdzNjwXWKB8FhZ/4KI5GX25AlQ
URNpzhhhs0rVdKpvv6QKC51za/OYUB8nPDgfEU5VWT3e9sWtVkXpwrPDJr8WR9tc
Csb4Mvt2Y7Pi8TAU50cefnlcfZv7bcaTCNA80F38GnLz9eYqaPdsNVFv57ww19oD
dG/we0oewnuvd8OGnwX+9AouzVtfStsDxksedbjkH84oBlShO+GLcftNH+TuBMa0
U0uTOEFZjyM125jbJ5e78gTYQe2xKPF4NLgf3EtqPEqFsy/v+VCVAA3olTq5W/C1
hxcuN1fjyWcLo+MsbpvZ8f3UzoyM6XmslPNSRYFNXF9vzf7Rk1ezBJR6Tj1gHRTv
R5rvzOA/6CW+lFWoGz2uM/O35bcfQcwww7jfxtcCCJ7dfl+OSGWKhFLxuXjOu5+F
HVYu2w5a83mzClpvvIQovW6kY9YavkLedtlBuDaT6bqAv08TsO3hCt3E/wA8vWYN
CIvvXfAyJPbsYoXD/LffwYc2PeRmQj3ygoI1OKfqNG3b/Xwb5/Ct7LARxtPCODeI
mPSO9FqCjikPRLn4Fw8E/KHl1LuCpVzF2WVTzGNaHao1mwF8F43d/5OQQ0YELwS0
jRFWyWDWFdaoYj9zqxvvSFlpkBotDn0AKnUSMBAveaJJzzgf7KsPkWYNlh/MSTI+
1UjUTUO/iNbaG5gIbVP9DBIgxGYcZSb3T8pcGLSYxCDX/M0OjU+h/3QehHuQDB3O
qeGjBtZUWoPpwrNhrpVZcXZzX8RwpDWyi/qCBZd3EJC5Ay28EUjjZJAd5KXjCFzP
eCZWvyk1xJaGHbUOvr4xdtzOPE2694J/M8xhnDHU0Is920LIa27M1x8pzQKZ2pFv
3wtlgxfIf7p0Q7IbwL1NNtY+TLufCQm0TDBX4XyVzVH0AqrDXY8Yr1H62nxgkvvv
zT+jSwJlCAaEDWEkbniqN+Tvq14Od2GxLDECxt3duJviFOUGxcjCrIJpy2KhQ6wP
hQiG7BMkcN7ppiJnpMzA89Skhu9ruvHtl8qBx2ew4xFiAtKzZDuaxYF5vPEzCkv1
iOGEsnLIWZfVzRSWAt/l6YHr2qTsr5v0OGX8AEuuBQyV45Quz6pJl6L2/PrUm/Rv
ukFcFtrMBbpz0HhYXyWAEjj6SMgnifXj1W3FB7s7IjQITsvBiloxkYBAbOPB4YpW
bt6gIp/Gk4QXWhf+HacTOQA6K4UTUGW57yJ+jYbrV0ylnoOhGxUQmmjI6APPQ9Bf
dnq0hzfMteD1tu4QcY9goNzxMJMQToD4r3GovOgiWyxrkRbrRfnE66BnqGyQKBn/
ciNAppGmI4hbsDVRvJPUELRMuj85L2sPU+vEWGOvzwE4XO3YRa/piGqAQXuM5b25
nJYPGqreST6rGgSQ4Er90uzYDAv+YNqj86DDtEAWAlUF4MwfRqo84Rf5K3aSdgS6
o+28lT1C0OPSaqnUXnCn5musQpsT+HcHsLi2Nax5i3Y8ZH/T98WbxeqbA5Mqo8CD
pjJz9UYThI60B+KCe+5LiLF/kR9a2C2adcEigOGbyVS69JEIzIv0uc96P2oJ8wef
PPH6cxKJpbb53DhnmrhiEFLjBXSWW7Qt16ZTK22NjRjRfIzFlfTkB58M+i0a2TSG
0veQWQ/HtsPHFyktqdrbM9DfNYrHBf+unWuzga4ETOhPJD6DlcGuA8JJPtHk/ztK
FRYVW161/j6P+tUIk00kcDBWyHzpxjwy5z7WeFHZsyGARGYTMu1seqbj7Ct7i/GO
o+Ff5plt5r3AbtI5EussuCLwDIVpXxLZrc5h/aTazyDW9k1UKoSD+LQPjuKFeyPO
ITZHHK0Jzf6xhZ71BUK3BHleI1s/PLQmoY3gMZMgWs+h013rpbymjIzAznwP74BG
u9tcKKprzJ8QVAR9Qcx4vvtlqmHFCk36/YXFmU4EqjyWcVX63P7yy5J+W/Cm9F0P
LpICJDr6qNkHNr1Wn0+15fSC+bGP9X6nwTqjlYr/6L941LgK6yVFt/JieyeRcNsC
zIZMxbZW+STQ8ZgszMHoqxeMRnXdXLSgh2HZnD25ihqJXIU6f9yqxF2AxMLPvoiS
8xs5nOc7YQ2o3x9w2kqy0aWfp3IexL//KLCmOXDaydLcMRf19+W8+PC7hTxcNSnF
JICqejkDWWLR51z5gwtyuG9BDLwFrTWV58lyZ8s4Nh3m5KB24tQVxPi4CgZAsJF2
PDZQG6Z9OyTFDezL1nyFp4r2dRYYuuX6MknzeUtlY0hU7eAot19pySwx3j9ZBa38
zn547+h/Lz3Sb8LlB7pBE6Nx6DCYZ0658QBjhZtxh/bhDeMN257/ztCWv2c1UiNO
7rM/ml86PmBIaaqVEcDiF/VR1OcwWq/V5se0cMC/GQsKwBAWr3CB3KDsnS2XlPrR
VrSqFMdnIgZNN6R59x2n2KIEDm8A4wOrerQ7RR272UC3Cuf0mAWHxeQeUR8pZgkd
2yeA0rmnjTivpNYacwGVvqW+Ar/jB+qs8A1Nsus/aBMKapcszjfcUipo86mwkLRN
siM08TgFf50J5Lo3EUYlmd3a0An6cKPiX/CxPLTvgTtivo9Qgi9oYgNn50O72lym
6cl/7m2vXpcrrZYpC69eI0jAy2LA0oESQrgYiAmtJ2dCAWGQMcM4+hfzaQXFlUj1
K5wB3q6IuCtEGX8AUwBMC/Tnoqq72gClrHk/rjNBV9jyYBGwq8vPHyjduC+0hRhu
Cl+AlMJdtRNkvdjDMHvJmCdVQcQx83X2WqHyu1w6UGB5Pqk1eXLdgQuzi9RAgMw7
qyQg8FciO/hjtdq4W9yATLAdeRpAMEmvUwnde3an7yj9zPsBAarYJyGzvjJNzmXm
mJEBvks6Z5pbj8TOKmreZz+nvNKE9Rxwj2+KbtCn0N+4o4Hl52drUZxaSMtnjmNj
xa0lWvCFwXLJ58RVnU5lQOSop03WFyOMXhNC3lfuWs9DBX+868/o4SeA3AURkrvY
DaFM9TLN7HJ0eB7l78aXhD+IXYbARMrgcbQn3RTefnPqGr+w3xqRoZHnPm8LcWT7
dzaJSlGrSFGRh8W88kwVoYcRFeGnpzO8pf8o0Zl57x/tGzZb3DFcvwgeCn1gC3aj
/6pBhtdD86Mh4+zXn6b+OjZO1YtA7iXM7EXr7p5VvSrNKoPlkxXwP6CbFgVALZqV
FU7iPuhheGlpQUvI+0oiC0jP4sHgBJfAnNMRf976Spsif225OwptPw08D56pmuTl
psL2F6UP2LAlZJYvHTRZcqfhrDBHlTP78Yp0cZAsX8ieblsGu7Q7C0UJ+DzdDxWG
ctGl3ligSjUb6ryzkj3jr1qcIVXwEPObxEl56asnINxPyHDfccB/lfd8mDrt6Y3h
9xkX5tkscUbO73t2BxBO0iZ1dZQy49cib1ms5YpZsgkJja/AajG7pCj/2iuhS/Pv
vSOldPNpwQYCfLObCkuSwVFGytB7xGhNzGUSQRscjT5hpC/4S8IQpLifhCHh3k67
ca53aCy3/ia3P88iLWXy6iop1Cn6oa4E0Ai4+vGd4+JHu/I35YGtjddZ8w/q7IXM
QhG6VZneOeWoXkRlwREk14jDQ85qcyE+3SBL21S7Z/me7McR3SN7F7q5GbGN3e4j
891TrPf0tJVVRZt0Dku8U+lqqFc9XS7hZhxgk/acUFxqNs4OgFyZ2kjrWq0hJiud
G3/tagSr+TS/kh2nFmNLu8QDK1MkMjCWRoo+DCSLke2PNO32Mp1mDfvHHIYeBtop
SK0NSZJmt2BU3MZM1Hyo4mgOXtXlyPQ9U68ZNGSJN+RGFbtuo9bD/jCMO+J1kjr0
VcIA82xJlo7Xux9vO6ZCVu8T19RPUIKeP2ZI6KOsqhs2hSroV1IqkbDs3RoJINtg
x8i5a+sQlSXEyk+W/CpR3d5MnVucmwMMxzz3BB1w+TypXMMCdUk/KttJPXIJZCsk
sG4zNOdSUfko7gT8vYNPMJUvQplo2igSzgQPjLuG/Vjvo74V9gLPRtkA74IAwekV
F3tyq/ep55lG21zi7BAkgb0E9MhBeCixeso90JkkS/FuT9gogA8yPrHI0P7IJDzV
mXC2VRrdmSKfmX/mKWk8A6vcaKSEXfUUtOoc07S39CfKCqYio/we7QddFiJLGep5
IWapqjeUbKZM+nmeDpRJp9ert0IRnUFPUn/pG6pnDIVWxJFUcz8fLZF4L9fEUEqa
mTyja9/DxfPpzF+IK6fUlRx6hYUIgoY90Lau64V+d1X2sKZxVxq6ffHjnKR8qDJz
dXbk+yioNX2vsuu19oCuvgjDoaVRzEHsVc/3yYCNZKpQ+Cby8OuG2WB9vp6P2Opw
A25odkOWNXnSGGm85cZlh7vXoJ6kxlYPX1iTGHADWSAwQm91QKVnZN2f/b42rTo/
OCIXU5UMVlPON5PyLS/+cOgyISBatrnv1Yo7tAcodiXDPxbdvua5a3hFJ0L+lqH1
n+gl6ae60JiDimygofddMdiVt6knRxleFA8C39jRWxeUhTAjnJN5oE2gt1sR7/dy
78SREVnxxcf8nsn1erz9igeTh9k6iBIktUOShN52rLQahjeih+G8k1pD/toTikVv
ZA1qdSKDk0+0SyxdBWSGdwBYqVgLnf3bqxdsSvsguuAPMgloWKmhOOfY7DCLe83P
zFFPr7GPsUkxK3ttEljswN8GhXCZQQWqhb4lJGWs3YQhdCrneOVhRwUmeZMRiYtc
rzJ8VsI+83xH36qpRM3A1iE/4K/WaC/r+UN5X7hsWpcRa7pJ6X5YRUKsBdjcO/99
M0lcuzhWIW44fJ+Jptm1lfoDYntHaXXQ+Yc3bjWwkqhS4luL0vyuCI5G6hNgsn8S
1EHD3bWaDQ348s5aZhCKwpWTveqiR2qW1dPloa/E7Qs0STPf5j+YvFG6Nd87pEKm
5Zxz3+BLcR1D6iRLAY8gU0CvybWafrE/R23wOib5gIbMmlrVXvpGpFKt9hveOw7s
vu3ncvIctbC9QksxbI4JIsH3Ife/VwEITUsphdvVhlvtjBPh/tyqTH28OEtTJmhS
qVJdsgdrgewfU+DJbrBk3vVVcuR2du7j/u6wTWbDVlmRvWwpt7oMQO56OhcM+XLJ
t/Z71As2XvjeATFZzaMNuWRYm1NxBzNtKYGnq0W4jcDh8+jZLuVPAj9r30mKmNCW
3LQhUZRv2BgsdNW8GEQlZAndjqtHdGeVHiwmDmsWYTtF2sr8UUpNrEJxEaq2dy/i
8g49bfRsf45+Wh2AyliXmwiadBNXxSlJeJ9OsmE4fnr7pLVYHhJpjtE2xcTyKCFs
fUCYlheKq6iVbO2ckg0jerop012+9USRLEzswhsozfkTYMC676/3yWrdp55U9yKp
bIkkmmvA969yK8bEumkwDsi3tVLP5eIONhe36Hz38gkXZ32VInzPL/gLHIgAaZE7
QZKeMe9EFgEIivt1KvjexMDJtCnmc61PS9tF8H5jVwVo5abJel+Hn3qVwPSSQzCA
I8L/dMLq+3elFmsjjWyd1kGtkRBCTBxMr8D/JYyHDs0a4Jc+aw7eBOR812+gt4hd
BockRDZrPtV4XjfzKGewNB0Mi9mgW/R3c3sdcP0NctUSOzMXLBMUKWTuojJvmiF8
p9ehOSjNmcuqTl44AHUddSbyp/6iwBDRHf572I/GfFfcxrO8js0+aWKpmoD/kAIR
KW8ekXo6J+1WzMQu1ROsygrVeJSNmLryGTp3s3p4cCr6nNQaGOPyIB85uopex6IE
j3yyl8ZE6+2pBNtTTDzQljpDTvSwoqT2tKH0gcnppkjePjHmzdAIlFCIYvfLXFuA
1e45GwJAu5MGRH2kzLtEDTQ/UTtw3HJQ9msYkyftXe/upzaSBrd/j5XIg5Jsp+Rb
DP4oi1j8M1itcdsb02cvrTyRhTFCr47oozeJfvhlFlWlyLsa5CIuYq9vzBPAIH21
YmBYFL7QdrHTMhRv5sCWlIWwlZLGSTKLAxfbGpSJ5eQyeeBmTbdbATVRLnpdwpr2
i+xxOeIJdO9DWTkIFvW7jaHOI78z4pgrBHr7miWiHku50SkM7zHJx1Gav/lb1cyA
a57a0jy0U13s6DZXig7zdPZJo4bVB54RF9xMe+VAhbYjKvBtifobOQXVwjw3g4vJ
P5+6O6RVX62dJYWLBKjSHriUZWxWkUDeTIXzO4b3DPpUT9NhVnTlmGnQOLOxO00A
6RLRgBfn8wxJr9YFXAV++qx6htKzIIBDAcIhBn406SXq/w1HqMc95O43TlZQqKJB
05YroxVGWCOzpMGltycrelPDHX+MHCoKetXkOFIroVkg+9LipuE2Q/yT1hTN34Na
hLV6tkC/Q9SZIzpV/tdzf2i2slWKIHzLLzIPuL8ycxGOHyRFD0H568gBwkhWj/gN
Nd/WLk9K/NeL6bSV81NaIM/dJRRaTNjseR3Oz+K71IqTG9SLM95yW6JRAoW1CRYm
oSBmvUdLDxpsO43eYZ2y8DMhQH4GJ4wJALtd128dCVbewfr8kGErnE5RUr23/hxD
9CkoOonoTqS2uqA4HwVDMdR+qLcnlj4LN4xnMT0tnubILN1r7dFS6FuuuLTUWM3L
sF2l56L40tkRb82AJ01FFQ9hYfmBKfRtf5coFQslydmuBQjRhipVQ86bJ6GJOJIy
Z8AYNrM+WjAGq9zv/WomGqk0YBbxsRAiMM7FWH0n++HXekPNDUh5o/k5t2ItJTl8
GVkU1w5u7TTMBm7GiVAUQG7vwBLGtER+q8ftQI11XClNtNR9SgHY1OBkLJiUXf4b
8rTbgFAFikedKo7S67nofkjbGIXq4f2hRv6qurQOSjnHwERafC3zIEOjuwsNsI4X
Yqkdizt3WBr5p82FbCkf6NHgJ/RoqbCNs3ay3ab/Lj+GEESCy0SJjYDfC/0MwKyh
7U2hgcZ1iRLZt6pXiB6ZYupF/SsUjTw1MUFcPgyQfW36fPmDKVG/Gok6Qa9JjcD2
KjDj2YX94WCrSh3cS/6lzDXHXAMediTYkUiclysbjlJ4EOVaoqT5gnljmT8DvlKu
rFnEwKS7OZkDM57/R0l/5OieMsbBmX4c5LW5HDMiVlJR3HuhipsjgM3tKXJ6Lwur
fwPdUF+wNReywIGmoue2eeFf9Z/J3+2h6fMx9CwFH8qfpXvq0PIMvXRba8QmgeHg
Io8HaYO7bHuXAaQ+dHHe1KVVi/g9fwAjqThfP2KWPfYzjwULLhPzOWoTC4ebCTBM
iindQiCc6a1rL18YdcPp9gdd3DBorrtvtoV4oEsGp8LOYlrWOHFL8duHVSw9qdns
YQby1qPo6pSQCbIOZbx/1g5m4jfhzCJDx7aBGoN9DjpI0SI/exCuGE9bLd6VwnTu
HAxu9XSwk5kdFAstaZ+SKOpbIJQuZQdVDPk7LfsxajPoqnRkZxmmBzemoMQCN4Jp
7p733qJ/9UpGKMQ7Vn8Ip7cj1U3rQB/nZNHLeJTJXDc1TNbrd5aAt6zmaaBJ7FcD
hBQU7maWCuutmv1AzEBA6jvh+5SK0tcEUfpQQLGfgVc2pziUjDOVhwbyaCeALAKc
EcgfJzfENi20MoNmnTURqL+c21h8rLEzQKdNFQk/hXoxvpGTIgigOz6O6TleOZQ8
EZE5NhITsJC3rFGwo/DKzc+dZ099SanSuvQaih/7KoqRwth5rF0sm20CXQ5mMXUa
zXNDI1ufMTIcUDAKZ41fNBotVCSNVlKznmz0d76UmJ8XB8xKf0xgNqe0U0hPOXQz
urwY8rW6bepnSeyZnK4d6Lq3gplP+eq0V+Na8hdM9KVMQ1v8MKi/DbKKY7QTil5C
7SAGqTaVwk1veNevBXJsKUe2HDPYynodIrWu0snDqdliTwcgHoHZkW46mfYunzdJ
ZfMJYEwIE5RRDaFSg36YZAdzuWT7LON5DIYthka6h0q0mI7pZDT0dMKDoxHIN4p2
SCO0fadj/WiHsnkTPLxqy9i54WGPJm1CspGNXWXx2YWCOUotPmidAZnH/J7ZeVC5
+1D8BtR6GzjHZIF23undjylUx2U/5Z+fXgB+B34+j2SqKbS7yB1oGPD+FwwbpeJy
ZzoMST43Xj2YCQOsH/DZ3H0aoC1plXBIGoqQ97eJL041rful/hohW9gD7JDkIrrk
5fmjO+iuLxSW29JDezP2sZHkpupG7Q1Bj1i7UGRPMazgua3125BwG4jmc3d3cYyp
n5yi19Yxa9b4atEbVnPh19LTQvz3F7SMhmaEpEG13bG0EEvYxRHOI51bYZbpXv80
93afPcA41BggWF4OorVxkD2b/9MVQbIYFanIobCb7IsQ49IAE73UvlKVe1bjOWlM
RggYvQb7GI8WotmnM5Wji/kcNhOrEv/GyYFG/SvuHDqCaCtEqJ/APn1PvlKol3Aa
grP4m9DVQ26KFB8UXD/gJEX7UQx0r3cN38+OYMAp+nLDQPafrCsAORPiXx22dadw
um7SXxuOiAJw2TV01dkWmX3ByxPU9qqz2+Pl7wWDzb6PwuuAWTPnHjE7DB08HYlt
RM4L/l05GImdB/STo2qaq3LoXC9tbdYp6o5WglFbMCBRin0ZoD+1DqX3bWa+x02F
Vd2YQpoqeqN5GIFK2EiOx6MoXwRwTEOBeNxF/4rJ59hrdiB/DbvXRM2hE+kdpiV+
V664M3fIKSoSwajISrQWKyIkkLwh5dVaA/H6vSZ4LeMjXZPFqfwUNOq5y6jPXyC1
l7TedAFLCY5rlgtYQFwgaw4Mky042L8ipPTC6NPX6l/fXLQhpne1EVo0XsAAPhzy
Woyf7iqX6qeLCPxf6WdtiQtg+azPEmF1YOxfZCQYPQvwMTg1xTidm/zWeJNNhEeM
9UxwILpvnCOCfZW2Ue8G0ZthCxPSvQb1eYfR9kKBtx0EBgZs1Y/EUr9BFZwAbFmB
1pMbHVlraD7WtF2gJPDZ5jNA3f0QD/qKG/MUBZhmwphhMppzRu8Ob6rZF0LxXg+s
qlCXY2Xxd88ErjLK+i09lbjfcLtb8bj8ov2/tOOteKLm2VRPYq32S+JdMwPF5kgd
Bm+WhTeF3qa1ED01l385BXM0EqOaNDlcU9gph1ipwyc5IO3cGMh8/yLhm3eaELFi
gv9ynzKe0+HTuIYuSOuptkKWEdRAe7Qo4HmokG/AIbheiSava5KwUjrwb6smIAV8
MU15dJlj5DFyaBoIE4syRT8BBSrqZiesa/t2hID0+Vz1uZHsvuWu7SGjtENn2pJ1
2W57rJt+kvClLF9eHnalUmnP3+E1SL6IpECuYds9JcznZMKjPjJkL7OdVRedhIJH
H/buiCpifts6w8zF6qK09a8PD9iw8Tpuu5J4Ts1zouSjix5o16V5MRPTfpfg4VdM
xL3t2dSorBuOg4TMe5Ao+Q7MraLa/PIWuXkq7+DAD9PmNUrMU8S3ImRYa9GSvQaG
+mmXnlTJ31Z2R4jcx6jKLLJnkUnbr6tRBkT1heu4E2tqpXTiwp69V1icqcqEjiyk
5TDS8fVFYeQ/oJ6PcBL6XEQQwALK0Ca8dx3dOZjKP4NKKVVspk3CKcXd7dd92H/A
cMLuQ4r3x97uAfbmiHIX0W08OPFSZCoosMrPHAXwfQfv7Z14V4RNHHfsrFK7ylO9
zNkPQp9ZWdeihIzUej5ZymEd+P8HFU96pWIPInIfLlO9kUtS0xVeS0Msn51kWL8E
rlH5eEE2CK/CBryTUGsYKxQX+6RoHkuf9jEkieNVXzrvwe5aVrU4n3kA/dQVkk3U
OVVHdb9dIs2mBwQbhgNsaOUeb4hc+d/am5TBqIprZf/pMDk/0/AJePbSgesCsp4T
Gf8ZZ3hqcW7DT0L6GW5inFPR5yIRejKYS73TSfQLZj8t+Z72Q+LUbkVBN+ZSqPQF
/e1SqMo+o09njIRLzak5vCqanepFuolzhDHS6rfu+lkClVNrW7++8r5fX5rO5bL0
3q89ph/D6tvdZtc+WWXDGopoKxkZPVgWIGqI4fltYVoseNDfIpfD5aFNYVdX1hWU
UAKm8IIznU5YW8YmMccd1auxmuFFVQNnl3/enPhDKlVjM6pOFiFA2R0iuOF7TxTI
cxnmLcTQTtyqaWlUgi+Q1K1bTbLVA+xfYC5UiNkYczTFa7ppSIG0IXp+9ljFPZoT
fOCw8eUAhyZhfNiimzIGJ/WvQfpmLEyjALCbboLqpU8vstJVuJ6+L0J2hQ2hYxaQ
08/UqhysR9CjPPPZvS5Lda0n3745vIGZCAEVlGxB8L0Y6fELJzaauI/LlIHbuPjF
LHeBvS6fGiJPURU62ZwOXpbR3kSYVABubFBrtxNmPK7RbhSxuJ/I5zi+AXHxM6ju
e7FRUjjy5vxQvrxByhZz8NqxYk5IdsWsn1kHAaqUUHEnAga8X1BdnceiR0rYbVc1
TlVvlecaWPwRrbDPrsTut1xS/MU/OncLyEDx5FhdxaeLcB4n+uzgQMynpuU2SoUf
f4ZhbZYcUf9enposeEer3xCkIXm2qpWdXPaMAFDZ68u77dxDdkp0AL5M+xzw6bzk
xCDOYJigIXzjTeWb9VgZNHWuJ/mt3Jx2wbY3xMn6J96tIiQfcRxPVHbhZl4EOtli
5Iv2ORWtsmMvJJTwPrZPH7isNnaKkmq+IRqqPqA21YqC+hie/Ig4HC7bQo5hZ+u9
aW5VycAbD0YgpOl0zer5ZJDRM+9fDc5YdRxuSm8weu7fv7pBVTJROJTT9E+K1G4e
cUD0V4Da3JKOF7tLQQ6dXv3i1caH0JcwMEvop2lsPPGn8BTm4enBvwiC7Yo6IUoV
9ydz1wFzNI81DpLLdLqo/VTjZ971rF9Ln/Wcojm5Rok5D8FQZk59NlLvA4uBXb2R
I9YUmh832DPfzqeBbVx3LZVCUk9yBnOGPIi1f/SQPWj93k2821y7gSuRtDAQYTAd
VXGMcgPgpRY/Moa4hY51cFx82q+MaKVmWluVdRyXrFhHiQDf0Oikuvl5WyGJlk0s
6gxSrfP+edwKGHocCEQIBHJ8r+6zSqHirf8sUPqC7isVW7+4DeLEyph7sdnrJh/D
2L93Z3vNvrjvMWAqXBdnX06yKNLrxbe9vMTL6K4ttu9i2uJbbYENXYyikbz6x9L4
z3IJfLtp3LUY2sdSsjmD6r9AR0E6NAf2C9qg42+/wpOnsfFCVxNbdcLn7oqZxV41
PliyP4ZauxkMdsoyI9rlULL0aQFxA7IDa+r/yMXs8vDzvxjsNMe8KZfEjyh1D32Z
l6jmgAaRALxaWdiWjvamZ9q0LphZqejMeBydv2e+nApuZuY/yCpXixo42ggqsXGX
8dPB+6iV/cIxw9qReQaxAzbwJudAvZ6rWzRmFh6CTgwJ85BqJ6XtcWbZvrstBPvp
o64u8DvmelQJ8wrmOeEyRE3kNDg0uHaX0sGVrVgifbZblMdO8KIvSbW7KmKzbI1Y
JABHMDdhVFk3z53KAnC/oyWe/gd/zDa2q+shVXZqhEDTfQQtAB1Kh9K0CW5bnw6k
zk/PQ9qyJMo/qVap8wa9ldS21dSI2wY/oX7qM8FUwt/Tqa/LSblsy5fV622z6QWe
UvLRVKYLShVqJwq/6Zrszv5tGpNJAc2D/c/kDWIAwW3ykx784/B57fiTj0F9q4H3
AXkX0B+RpqfUhGeZMmU0bQTG726vPaffU8AH47j6sgpjwwPeaNfcEUaFeIwree/u
cLZ7mzNyvhVczbA1Hnuhh6f+CeaY45Bs+qVHSuv1if+n+PfGJidnN3UQZqWhQs7O
Jkgk9Ab+tQ5wbTPCbDqszlnvxoj61DPZ3Mi0mgRbDHCsnxdsC6bJKN1W7kLGwLpv
eDA+a4NJsin5nwGCjhvJLm+zb2pAqXIk8V2IqYoxURbCuyMhuBTSUcDDHWeDbWgs
PuHZQuSgEr5FLZNYyFtjPkQ9LBCo9ayQE1RZfjD9TCnUwtqc8d2xRxD7ivv4xD4F
w4zyqLZ9alpQC1Au2yhjjW5kzkDsRnDUeF1oZhZOivww4aDUjyHOtCDCudh8TLpl
jpJvtrZZzjWEA2UkZ0wRXDzajhK0TkTjeycuPrQfabuuqZiCpE7XcsRBf4c8JUBL
rlUwHX8xnhJiQx+0oEKVWXv3Lbvb2n8FNnkDglLyrna8lq3vRV53oKmp9XxJwJ7r
TdvMVwGh74G4By9MbvnigOq0QtUoCzpPh6w096RjIRXXbvmPuzIT05TwU8igzY89
pB3Nx6p8/06pj/bQvfJqSZZBm+40D7VEXpAvoz43tmDGd22b6u6XToFmUFMslYBq
vMpr8MYPbcYQ2H29wRnWzsIsK1fgyls7D2ajo3QscMNY4iUHpOsc/pOoUzsCeiot
3iRc0GlNJPxNAb6rgHIXkY1hA0eTa8KJRcfEDSD99KZRdBFzYpqTJlPCuZg17iVa
rWmlOVAQo+09f9SvaetuApvtieDBcMdM5kr0VSkBZIM2K9jazY+BAQPkqfUHeMgf
H0QEVHEBwghQ47gEkH2JkB1JrbCSHhiHgB/OdpTKmIsKYJuGktheYH9JHYtFqZ9V
CeMI2Pf6QhyYX1X+yGZ+jyayMuY19x/wfE0xvJKqPZPZi8+QkWP2LCOJFFLFNIy3
OHEHa8DZZSOIdZN8tWWICJQDTIDGqHQdQehU/vW4x2tf0ht9SwQTYW9yi/W/LQ6D
0QKOGb8068Nn8S8Zk2J4Xafko8I1jra750f2m5NDDweQL4fdLsCHflCS8C1B2z5f
8WUkJHBPCh7n6riksKu6OkT+mbhJKzs1iJBED6vMrdyes6BZ35fy3cJ07u9it5+3
Rz69lE8yMFqyXkfCiQnrjyVWgyrgzVAnP9iqpqEJCTep5dT08o2omcq72Xwn9Feq
htTy6NuHYD991U9JaB+umMGwcTZd1MdRljFNXyjuHHm5FQ6bfhKpDt196DAKwWOT
Or0v0v9+9Bg5m50nbzG8bSC7ZQUA7y5jXSypLIHrNT67yWTlimirYF/EKl4uvT5q
3JTNTiFjcvZMx8tvICZhSu3ORiTAv2byqRtKDvupFZnPFHSZ4VhtHSs8r6Jcjw5r
4EmEyHkKOijgn6ZwMAG4RAFUnASjlfNdSom58J9ru7BWIOyku0YJiKiJE1x7AFix
nw8NvU1NRyNpaIdIe+FlTZRBucGZwPY/7QdFdGpS4Sj2ho3VAeP8VFNk/RR9ig65
DFvyqsM40l6LYJFOKplOnMj+0f81MZ1mN2zJHoA8Wtvs4QCGzPR+aOcHXCUnq0oX
yt+fPgz8bBr1SVh9/9o4pQlA8RVNeQrgBnJlbUQ0iUiKsF0tuWX4gNz3vWdXAzlX
t4MVm9ibZ+8f97D5da4i3J5s7dLGClQLQTz+IJy4eQcANK10ijm83xo0fwJQQYkN
OS5yyia09qF62kZh2SPDNgcgDaoFRCdA6D0Tz6efHtWBkuZthRCNUDWJaN68M3uP
PO779xyETH31IF+vS6szkkxHlZ+AopddrkgAcH3TQeJx6H12ZSHXYob5m24bpmnR
99CVB9eZH/1oI3DUKYxwVjQ+hGsmwHNEMz6JYE+hoLTcPc4UgzR73i13Rpm+GgzW
5W9ekRawdMX6m8qRoc1BXfyvIKr/C9m7TM2plZd3D+mgLaW6i5RlvedxyGo+QlYD
Q8oIb/pEqWoC6GenSMnA6JjBViabUfeet5mz3q9ltTWYpnmQLeDRQGrFLHJs/Z+/
nEdfO9Al45+cGCPCQP7lhXYePsSEbGlrQEL9xc5VPxl+2oPA3SD64smDIHxfh2qv
6ZHtbvzdAD5WJjxR+yyP95KpzG+kOURCFVUTjxKB9nOVA/E07NeYNh7c8qdOHHH4
pncV5aUJqcC8vaw9nI/Czcn3HJkxlbVTFueH2zC1p3Ged+Fon3QhXxWiPSoH//Xq
MZhDS4UGO+ZmtwY5T03tjZLIwSws4fX5iiuBOvENP7OYjyo8vyw7jAtiRUFwzPvb
hD5qyq8OVD6OZ28+sXPsTFKTU7iFnMnX3gGmxBgr/hGu+c1SBs9iBHOUl7CAfHAN
wefCtP7q1YO1yZN7Cqs0i6j9ykm/molw8xnFDjRBNBXG3YdcvMccknbOELoT8Lvc
5FBNfRuMOaM3KNqg0nhArAvGiXOLO0+SMgK1yRVRzyes7fre/SX4BXSbeQ8Ko/mi
BRy5Iqo4k/7I3qTHFlRvvZE5QRifLtK2Dxf8Ws9l2BGNreHWQk0crTC9O6CS6U6I
tUqUe6lO6QPsyUlBks5QCjS6Xo5oDPTpxL+r5YYZ+IKlFga1Q2a6II8SsSVqBEfH
4ugXV32qUn6bMdPUWLpRa3vuzz6kSWkX+NnWSgbJqdV90eSGI9kohBZSpu45CFog
mWnk3zwOjNBB8Ry0Pp+mfH/Qh0djnjPpkKMR2t80vn2H+saWDrrXPTe8n+SapU8y
jMA5S/MhC9exTaPaJRgxM/elLytcWJOKHPC2ZRYpRhIR+Tv9o7ChpTPKLJm6l8I5
qHQMDJZLhcPeUHQ154EO/OhiPfSpX1Qy30bxy+TgWx9q5AG7EQ24SxiBGA98wxgW
X9X1x4gJCjkCDM7hFaoelzgEt4R3d9/E4mpTiNbHuBDu81ZXRcvuXwcOYtP/TQgE
wI6rzX2K3kHG2OXIxeaeiaGg8mruW0CzuV5PyHSIik4j1uRqXftWQC9vpQHpvke6
ZyaC8itfhHrDwpSu6iqRHU8BbpszAsAh3OXZA0zA4piwrvda8NUkTICsUa3rQxT6
M6RDDupDKzZXrEBBj+czQemVIosiJCUScfZSD8o1claHIaED0ZnOgx9f6YPj8g6q
y5gAeWh4QMh186+9aG9VrUuXGdkUfcak71qztUuNr53H9+ApvztXpD9aPFOY6Ren
ULpJOXhgrHYrr3dRYewMn8wjVoiLn993X+MZtuw33+czIhu/KBBuBoTcSRjPC2Nm
`protect end_protected