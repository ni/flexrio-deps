`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2128 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
48M0DPGCifQeMesWYlY7NKiBDl3g+diOldxsgC7N4ZUSqhQb8bEvAH9IRSmAQHHH
+2s/zzi6D/dWboFpL7DyGEGaiolFAfhT954B8y1hpzXUnF0N9UOZT3LiOIK9/zLq
MFv9+8onbreXc9Kyujx0CIgc4KNF01ty5JMC/ryoWmet20p0DaXwm/q2kcmTlDKu
8s9V5ZWnN06duNC4meP32f/jzpsl0wEkFwA3xmlxMVMb7aGLVE6rZr6OMHh6SwFj
/jEkQctzEbfzVua/XuafQOPHRrRl/pRgMui8ibdw6GIMa9NmyXFBtSTubQmGkwwH
e5pJz5ILFVVHaY2EVHVO3rd0WYx7xoERfoM2R74fAB46fWVstKHasSVWzYu1sJsC
xpukpjQ9h3agWElEvXNPn5XoQGoF03CzmrpFjVwpDMZ9ifwVjaSqMkhFeJXMUTKf
7nIqsO9femhZE8vjKuexZBlTq/XJsD9OtQ5F5FuPgvgrY8ApnoIe63A2J+80mrK6
HZaeURHc647XMV3K6fzItUoUTopu8is4wY9fWu6T6sHgIlxvc1RrhEPlY2i0wMM0
5ekpOEZNvFuKKybBXQktuON7Gn0gYKk1MAwYq/OijXZhcFxO3KzCKZYjlv3B14NI
jCD4FhObq2DzqISH81P/qq6ZYIrkIzp4t8cNzhOXd6TxJUy762lo/yMhK8N7ADki
q4guIUcJmxUKPKKjraiC1OrDDgcch+IIH5xkipAhVC+TlV3VFsewETMEZBqBkEjQ
8xh2thNZi37fId736Z8uK01vrwYmy4krIBRdKB5fBukGoCHxxBX9oT/06ilynyT+
JAte0wU+SqDxyuH9PhlPgKI11/xx4zReqOHxAeQGsV6/MEMnYdiLt2yfEq7Mf3Qk
6VHnIdsIzv3QOKKDbsJJiTutsAiobyMFNB3zsGF7B15xl4w5QR2R2cB4/6oFeico
Cx57VwZT4JeqIVRr7I+314VT5gF/a2RJJhA0V+YxEgQyV7mxuAvDiviJM9gBYQxR
0XL2/0BeEGrrpoQHtn+WCza+Mv0kP0jFU9NC6c/4gLYr8BEepHG0e5SU0o2LWxEM
HGAaEIUEpmZ4DUa6iYUKHIhQkGBTqAtbW6L7ySBwJGi5qUYfzrVPTwYMOSMK1oVj
/VRWBtp2+sEGa457b/BOudEsf1qWO3Cunb5zuLjKJHVw7rcgGJ6mH0XvBA2EZzsK
gdlgneWwWcog1sigqeJ3uiR0zNwPP+IGBYKeWItG7RLEopIqLVg9hT94soZc/FuU
4va9LH/JeacVScIc+DMUP/xHd1EDW+T03ebIytXLX/1ryg+donT5H7FrJYGaedzW
52sFBhBkuDfdJxF8gvG94RbJwt/Ivc97iR+sjVps3qXVQvpZrCyCQ63E+QDLhDRO
+3EX9JWioQQ8fwusR/ZBVcvHTqRtKG7980JvxFc2qXrh/Q1WeeNZmVJXlNcIGZZa
Q9YxbqOGg9Dv5Zn7CkKZZCJHd8vy8kNDnLOo9/TnufJRG415dlO6DK/eDsJofBmr
/Ewwe10vXTggkO8LR6/WFp1rOuvkg9Qo7Qh1PSb7EV/BmQYlui4KFleQFYPPTMjn
7OATfMTtwgTG/bjLWUJipPJLhumv+3E8tyM017/DFb8ukRqYvpfiC/GW7ksa6vuf
jJYTItBCq2CpDdIq67HBIO45daKXvS3ac/SNCNuJFi/UAF/95Wdvn04m8bqKKCVu
I062nYpNfTgXxpVyURjWH53Bb28ATArYeK+Cwxa5hSsUwzUPr6rK9N7wuy77VzB5
aGYNST+RTKJhUscfpsdgWQcU8wzqoka8XPXSE8MWWhXugqa5lFKQ+35pFPO+ZqmA
x3iVghfBIuB3SfuRwB1cW1CYh7InLMInPNaSarMT1jsu4XjV5aN1OBPb8pt234Vx
/3WI5PhW7ssmoEfss+Cy3l3AwpgLFQD0sdN0IHGuOmGE+ThwXrufmiUKtRl4aQ0o
vV1OiD5B7eiO6jAAhonH2dYymGwoqtHVblcGlChI6bZHR9iF7JTDkBhKZAfCv86/
b5MMSLdniGzniYToGW2IYoN3lAF7bbbOMqPKyx1atVCyCyJENFiEWNar/DVc8BKx
9jnPh4clS7FaIDKoF6PH28qt4vCw3kjO74o7NJi2BPfn2SMTU3C3sb0L4vriWNFo
jg8FnQIcw+n4TG6lq8iUZ3MfUPytw6HTebryyslFfMrV9vHV8px9rMLIFlNNEj3r
cUArgYbvidjTdV7fIC1Ogh3KTAsu5o+weYJfvzQtbj6tThXh2wjP9bxqzk0eNSRs
CI1PVT5slY/uk7f/2xguIvaUChl3mueAgSdO5NCcdEqIhijDDfEbp59EdmXoWbqT
snaQ8M5noD6u6sayV5CrGaGXcxcDj9b3pkSmu5ajSTCED6ogNoqm8f6N7n0uTG6E
N/yjEOSGNj0Zhs3E8lBG5POWrTuFIdQwhduSFH1HcOLB5VBhj9ebCWcJ0XA6YHwy
YS6P2WyP0ojsuSO7ZJThCZaRBTt9QVk6Uts0XCL5Cob3wYohhuenP9V7vPcUCzPH
7zII82SVoarbozIiVz0hmgYrB7KoWCo5T+dhF/yzWd27qZIBJfZ5OCyqtYJVEX+E
j+QQq3lqW/EI0yITDYyKs5lgfmMDLmbkY+qnAqeDG9uhEL73DNnID0+RPp7olomi
VGTesvqgO2a3xyElHLAUxg==
`protect end_protected