`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1456 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
CZ/1hjxIYH4XUI6J5JyuXRddsBBweHNq+CQf5Jya9s/pwGt4pbFVRDPHKDJMHetx
ki7ZYfSCLs9Vikhaf7C+8kxr4gk0ASm8RG14INNa/SLVpxDBVDmaMV9K0sCu0u6J
3jXXI1SnR2c8P15vbo4RfGEYfVvoooV+pDy0jRzeKeFmT5S2pEOLDZBO9q0mO6EL
NewHzsiW1RjrYqgSXIPNtiytn2TPiZqg7YAdRGm49lXf40HRNvcT0UwJdHPyxu2s
tjmcnyYZuRKaVktPifhmVsuIMU5a5Qk4tfFOnd2c8MDdnQvFqNK7tIORimPk31nb
Yztq/R8eRTK6DigvQ9PXWx83vHDM1Bt/aFTHn6HSzEu2CasauMboQrcSZSAp6295
sl0dNORCDNgAfjQhqs782xbWISMGA+Sb2uPzSd7/4VttwoZf0I46FX45wVbcSoMU
MOMxn8eEVaoAqAQjZOkrUu7CrGnNNH6Pf2qZKFBwMuSDf6GTpr92KC9NXZ12+qoo
9rDX7tdj3pnTySZKiW5UHLICQxDkjht9AHBtjCTzdD9HBs7cq8Vl5tgPAy0T/jLA
LQT7w1dl+SYvUAJOSERkDwDRTwwk+Q1B/cuyF9eXVlP9kSKpI1fXToBsKl3fanGr
23P1KAf+M3zgUtYFqSI0SQxt13g2C2F/wCWSU/7KvBnnGJ2YOgPI3QxIus2Eaziu
CavEmDaOQ2dIvbWjZif9qFNZNkIPA1PTtRuZbAXn3QpvOXtwSO86zODk8qVE4PK/
q3qFymKSaz68LYGHpnNWofROeL6hr5JrWoNWbGbgUPCKh5/9q1rBTbafGvCwIxY3
tgLwEZ2Qo3sT29JkZhL4aMz3XUfaVmYtDpYKndPE1xak+ym7/LIY3qATfLyzX3SF
eRjqjZA0WwWu/IwNQ9EdzZYZHAv6cno31l/E43a9W+IrEEB9/Qf7wlwpYfnrBh7i
wxzy36x2lBPhCGy+VynXq1ynqa44XAAjqoh7ekcT/LeavPpNhqg4xvvGcT1LzCCG
NAaxtN81HAkObXNYfFFB81kJv2gcpbgikCUPOERW128KpxJ7zg4nCt3Xn+QB1eta
GoL3Aa3L6QC2h/odV9GRiaxDVBmfvxr/q6RZtrHawO1Ilpz2KeXHfZog7tsdJZtT
T27DgjVQWAzQt2m6FwwDtexotnlkvkjlWR5T7qXSkHkEGd2BKJPX5Wx3RB/tFk1O
6bqLTXjmfmbP2YKKoWF8pXApy9eycPFCph2OkOCXFU8PLRlAqaceZJtVrx9kPJW6
/BOhNy/sle+7gF2WQ9UIxtHjnQ3Zk8MoAlE1PgdcrwwIXJr9/g97I0T5j4wcHbSe
7vxxcITCdt+dT38f7mtBhe9tFc6tXd5HQaobq928uACr4vYEJJy2cs7KjBiqwv+D
JytKmDhJial3e3h30f7Njhgkvhmwrgpb139hUq0TRiUx4LezToJ0rAsZBYHFO2VR
EmCzC32hpB17eYTkU2lwZcXm7L0zWnWzbd2hQJfNgqtf8OptZkySUthc4Z5IOVI5
HJz6w02VHNGaB/JAIAg+f9qx5WRibN0sO6Pn1ENj37gzDWyo4g3LtvbLCnBojsV5
qo8wARvtjbn+bmJdpAdC4CC19FZB+5TMeoZrphNzpUp5nHY9SfkkIibbmynJOnhM
zYhCoya4QJVGmJg02k9aMlCdz1D9ziIbESbZegUtrvkGPQkiaT2id6FgXbPIFuxj
Ib1wzFNG3014BIS2VGd5mFO1PvSD/HHoVODQtIJFQI0IHGiddJpFHWWJ1BWu3FzW
tbKtZfv3XaLCQBf5LT+M7g==
`protect end_protected