`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 57664 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
SC+CoUSbxx9YOJ458hhD0y95s7LCj62IOQ+3rzw7vwajSzZAcqmHUquHmUF97Xz4
AFXemMoe9BEXvCm3tldZrDJ3IRcX98HmBm0QvS1dUBJL/uHf4LV5vEY5GBsKEjC0
Rej9x3t1QCT4HEBN3eBMz78sWOPJZCweW6X8ZOppm+Bs8gklOERBcNelxmwlIadl
0pl/tm9IcSyKLAQL+D1r52KosY3+btnqFyqSsIjL+IriqqnIlPAj2JePbgpr3WnE
gzYZ9s0IJKuDT/bXnYARC0vYtLIbL1MYyyTEEPGxIR5jRjcuJvevHmkgPcC4WPIL
WJJccGPjRF+TJmfvIhw+kDdMrx/2F2cESx+yNciD1y4vdQygJza0eRwLWteylilq
WcaSGFM+iDEqGggz1ef8QKq/v1DDUwMOAXgfX/aTf4fhcVRbkENhc3BNRmJIA1Z0
E5suC9sMjPVIg/IV7Cgw46xL6YpxsDmqvmjmVAZZhPSCOLsjiNOc3lMffs7j0ETA
QFRU1m3GQCPp1Ul+LTDWG+xx9Ff9i4g14uzfnpH+DkuLceK+PnmjOGF6xmil8kZz
MeNwp+kdk5ULgjRwvb5hCfcAEP2CDZfMzDT43cFSnw+QLEJAWUy0c8jza+PUOhyH
DZEJYhekGUeEUV2HGWItHZoEYpAg7OKrqfsKT40Wcbnpb1HN9AF7sJs4uxNDlfel
Ey7zm+ZWB9Hu8pKniCoUG3OJHq0j4PNBO45+QN2mO/znMnRhwgpR2jX4OoBp1Q3f
IrjuzLfAgXU61eWhBaJo2tb89RtyZM1SUKJAamjZvGOJRoDwi8WUAJ9Nc6mw8ddO
rxgYlqYKeL2A8vhs1h8zJnHntA8rS1tCDm+8iPIdgNh506kaYT06VNTt0EQLn0Z3
y7bBWafrDsBcO6HbsesCXUNt6yApDUSdsvK9HmSO13N82ZvnxMcsOGUikgxUeT7F
0qwxAQaVd0xaATNhwvKEaZ9BLrhSMQM6xu6e0csStfTmydwYiga6zsRIHvipIHQz
HAu0+l00m41DG5XmKK86ksgHzCyFS8hTA+vraruPD+/CNQlm4hJwqVarTgl/Jb5u
f3CJJVifzNOlXFRtgy0Uh1eA2o2vmeuh4Rt9kYB3Bhw9zHMJ544sdIegI77djfqA
b9vi6TsCQN5MhgZeezX3RXDiAwHPxtFJbPovThj1xuHbsv8JcwFqdV/PtOHsZZN0
1GZVyeKnNn0tR29PqMW89a5d5AwVH5frtMqv/tb9YXxjoJ7ZvNr0u+kk2yEGNpNc
C8mVtZTU5C3/6Mph0HdI6n1nXv0CL56YRQT8OtllNZoeNzmVPkneYSWONI6SONqe
6CCxy3szweXTcti+U4fsiGNKY7oV1wPieFxhn0EqRMdPq4OGhW69xkBvl4ndwY/0
6A5RXdQ4FN2FiM2HpMzEBFTeQZs5gsEpVfhYCC7tEygPx1LBnG9RzIam/CJhGrZS
Jsifrb47OHg5z3ulsZqgCh2YSgBYShbizdBqFcGzBAjddpfi6YKZjrXaqllLgt6C
naZEqw4Ezl1hrWYJE14qSqIGrvDHYbQpMgLxEJkwZfMYvCMqUxvcyhFC4S4IHdhp
pOwsQBqoPqrhBXv2zmArvM04LUdysTyb1R7rCvk9ZO8h2Y0v96RpC4/oZ9Wd5Jnu
dt/zo2ckkvLcBXlZzJL2SdgTEKgIs/dAyGRf3z+865XL/yI5Qm3UKXECoKHvCN2T
ZQY/cDfCmheN9XIdSHmYzvAjR1k7TpWZlctaakWtuZGXRwbTv8CtK8O8LvAxazku
pSa/V0kgYptlU2qIEZ9kY4eF9uLbNiv+urbKK0CWGP5HHoi/kBXM72SW1GPilI8I
efx5pZRSaMWQF4o18/zSDktlB/XDcAFnv0PmMLuXyFqR2P6qkBwoT6JI7u5pNwip
1626PrMWv3D51LSMKYzN4GOlc4+Qjp4ksLx7zTgIEhYhevz1nRBpOI6qE2wKU7U3
mkG6R8KTH2x9cdaoC7s84URZnAGjay/+oXizmDmlPmgqoJts2yf/qVKHG5x9pEoK
rKXJBtuOpnBGP2t9hv+Sz1qgEYDUxIfGPY/Rgo76S0Y7t7dVEYhmQ/Pk3XCzCSSM
wj05Bxa6qw5qGcwPflAbvM7NGAtgKlfn+zjRKvazimEHz4g5Xv/GTPWp3lYEly39
pnaghT0zZGt1kmJAVJNoJ0xywFlACYLSosm8NFohfFmgI203K7KeF19iX79A4Zb0
uWM/JeYJ005MCRQTn7RsSgPEIyHTpzacG5MunsOI+u0enAFyBgkQZGZ7tnQLhziP
R6Hlp3zJSKKqpEWvwu8G5l3+wJ9H65l5heOec8osK7wUIcQ+So7I/02EHdQrasZx
gypKeTxzrf3YMcsqQrq+2hhM/cj81TzhviL06ZUhOgXtcnScq4p7jRaWYlEsz7y3
7DxrYP/Gsh4fyIneUB/OY5P1lCvhKKMPm2P5Xr8ITbTmYewCpn/xj0bzctU9C48Y
wQvXCvDDFdnl8iodmQg5tk9HsMSd8Ok9hRSmURPI3OkZ+CybkH5bcXqsVDhTeXgq
Tdvqs+I1sN1A9dkPi6i7DEtxa/xBSh5Yr51CNBhuaMhiKCRx07S2o6dzvOCvM2ox
LeoZcoWVIKlEOniiwqQwnzHsgaLpQuviOhJGAI08uDQZlcn6ujIVRqrGG/v0HJZk
OuGJKFz1lE0zaOcqM1bVw8fv8cR4nDJljfe9DgLdMCZjNrq/dI6PW/dpjomUQxFi
1nB5l+TW8TkKnQSQ3XN5hBEK1BRjWnfqMeEb6tKx/853dTTjTh0H81Ud9boWEJvK
jH6y1agG31nqoU8qkHU+ClaIMH7hY2XRGVlkzTs8KgGWysZoXICT5qmkVwOxLgRl
zWRsHko93Jj7wFS4dULKPjJ6zlFCmRGVMs5XBUFaUSzDM1QFOFec9758bFfRLjcz
eFdO7Pa5RRi8uRJ6XOUWuzDRXpIZh/wYqFH4QCmAe1bQTvkpfwZEiQWuOQxFPtZ9
xZWNDh4pUxwnmazGuyAP+/B0UaOA55jxkxs6JT7zVQwM69JKPvj63UyKoGntFmX6
ZDdknWG4KCAgyrDbrMIdC4YqpvjJVQ5f9+9p6NTMOam4fVR44z+cLp+VEIyEkzYW
r3FWxd010V8gfficI2hAl/HXERunbiAMMzuq3Eu5zK90JJD5ow24JGdJUiQQlpHn
KKSL9PcYz02MilNuKaW7ENE1HcIxQivB86qEqAcHQyDok+U2YhMkb7v+BJD6Flp+
uKrQYDeERd5NmMQpwra/32m1+fsZeqD2TzwQBFzbe4aeqzKn6KoIxDtrys0uxfoR
6McC9h9AZ7xcA5CJIye0oVTx2zDZiIpBK+73cAF0W4KXt/LbJrzYO/hq8tNiI0io
M6F9ydvXp2E1zksnUjxvpy9FgJg+gBzwJBGp5Yg1hC6Oa0tW/39Zvw7qye/nBQOA
FbNi+hZxqPo+thkI20udzdbEWoW7+YwEJbMbBDosgIFJOVCv7ttzYxMpZo0ClqVD
Rq7tb1z6A0NkHS+2uipdfYZ+kjo4Mw8XH878+A0atj4zL0WMFlGePVyvGRHD+F0K
OqCmlxz1qfs6IrWuqd6K1gxAlGyqEfZRZhNMuiIpt1Oere36J5KwPMNGJ4L+lUcb
u1PjL2rRYqCzpXBlTCsPQGJR7HTlHRFEmuBsIk72dxlDVWZwRJoae3AN4r1wFFlN
BgZ38LAqNr3pGfqcyij/El0njQwYGBeL3thYAsjNsUnFNI82sIagSp/C6bjtOhpQ
2UGHHnE99LKjCgriyV62MFM9vUWNRRESrO+/3wJggRpPTQ1IZjpp3SsLZMNdyyac
a5k9eNVAaxaAJcSUb0CHgvENDKAUfdNnXZQAN7XyYYGbSiaIYI9yvgqiU/oQTu7+
h3S6OkXKkNhuK8SSpVo+15ftSuawkTFEQ4mcwzze/X9B9lWklw14TQxR7F3QrBF5
LZ5WA4gNtM/ETJ3zJPITYWgio7RyyVQ2D3pj6kOIMr1CxUY2ZV1hr5z1UkSs/D6D
zz8eUtn76HG9RCvh8mWBbyUfhL0AZlGqxqfp+kkUV8dCGg2h6eF9AjHqF3cAN858
iFEZBO4k44h/9eiOJRrez4wX2uknFXmnf2hz0TWRIEzQuh7mJOK3+146HObvGyvs
5xeWGHiLx3ak5wSQcz9TYFw0l28SkJ07+2ArTQqhhMkl9Ig1cZe6Ih6/Lhd3FNFt
ubGhcxHb1mhGKlmaWmQ++eKZBRCfm+w1wBiVBomCw21nyHTxdC+Vs5G2HxpPrJYU
AY/ISLYONLz27iO2bLIOnFUsGwI7DECfx6an53SATzYzQyJFf/xl4QwygvwkTwWg
KsWSDcdJgmeE2pYVnMDpfbIeHBzZF/j5KTrfha2VwDVM/pbfuyJGIgkjzcMT5K/X
0jroDwAicU4xio+t/IW+3D45QTqlQgWIBS4c0XOIN41AqvncP9FvmKw9Q/cHqN/T
+1DNueF5Ql/yEEVz3voCvLhfU7Q9OvFsCzjoofvfNrYgQKFvOmVNrUvWPXC/1L0f
giiI4V3c2xnrBXkH1SVRGCtjxMDRe1dPd9ra4e19lskYPdeWP+RCEO1JM2fSR1O4
iobdOJLjFEwxzxr/wxXC2GLOwiDbrvszJyKv0LuAxYtaSZ7wSKDEAVdga51NhJRc
040pAvPiCpIbTEHie8hxeIwZt4WLzLEmLzZKrndUGtcZl+8v6f/hUqPUzLj1Hkbf
mj+JCWdRso94NWHMumunziaz3xxv1XOkKnneH+k1ZkSce3329fq4haw7O/IIb7cQ
Q6DmfywZMIW5L7W0H8B+TBYzjNc9OwpodLSB6W7RJrAg48DKDS3Wh+c9k1FCqxSq
Fs3bsRVXGz9ccFBzmLekk9+e1QuSRUc0lwnrkm9SlfXilTTfinSaLVUFAXeh8/KW
iXa6T31dj8YC0YtPZOHeAvrzUIyG9X+NHHKFUmoS+Dk6pQ66t5+zxFJwTSpWT7CN
3NuUOpse5B71WY0BU5WZ+Fhr+Gnk4ZRA632UF28ojutN7/gFDx76kVkaBAgjOPsC
P0BiouQzXWDMxizH9R8Yf2HH6MsNOU4ChPVVBSnmJQLrNScmnYnNU+VnnTprQ7w6
RcYT8pT9hS/LBQKt5d2NFBsiYF2eDi3pk8SGsnaHVZBNDPkPOn9gDtoI7oCpnc3T
JP5m3utGXlskqas+O0pDbLfgRsN61ASiUOxShYuP/WmBp1YIPAq4tUnGZzUHP6pe
VVZjeeelHCg7k4dTqBOeKtMOZA4gfgH63d/SmUWXYEfMQ30FX1nUqHcu+cPajLQG
b631E9Iqw66Re6eLM1n3j1tGD1jzy33zBXzSt47wHJXWYmoMXBwfkWtbjGGonaVS
QNnfyvj/tGCsoadcrQSTAx7s1XukbNZ0XKotiDwohDVT17lgw1GFF7C+qRWJ1Zbs
zXOPdSdp/WT4vYTeVmixNQwXdYGNw7OCm3iypCPsukgetHewvANinG04glYHuqA8
xrT50wKQ+rI08ooIR1yOev9AsZ6CfRj3QgNUG+QFjqcNNoPjJo0p3FOIoJtWb4nb
aMvxhLRXLtzL0vTpXbEJUjfLfFm3YLeG8wYvY2UByjDBbS5iWvPjcJYVvkHNEH1z
VGsgox8Cbe+TfgDZ6uc4fCSpWXCdnaSy/2IxN452WXAcVLbMHEi3I5na76zwPp2a
VHLTRpE8/ixbOSLKnDNxjmWys4uRk6/Q/m8bIVurUAoamzYV9l+8xRHt0daM6Aa2
xWOspzEN45hjIIhm2HcAof3lq5DOn94+uh1AZcYwqV+uaZEpr6sdoh/n3Bb+rEIU
9PmqDJF785USxPyeg7fjAOV9I3pRvVgra9lV2VnsQnOg6yJZ1oW1r+1GMQQq9CGQ
56LDmMJ8LbYqShI5QwnCUgPZw5y5FXHZOSFdDhLoMoCl6/7RKFfOOb/Jklr55jva
UKzOTBrTX3J958UaOdE/oGm7bmTz2Xim24XM/XCOnanrcqRc1WQT5YEcpwogpLQy
uImmqr+kwraPZJXEJJkQot0aiK5c1+QhQdpD8qDRt/83CCIN3HgSuL+mnSQjvbmU
vaCJiyO8GPeT3SgC8MDv8h7FW56azyQZs9eCXxsWBlCg7B1/nZn5F7NevFfwQhPW
65h2febXVqN4eCLOo8fmfZzx/K1ngOCcqgwqZpy0JfMFqFSFzm+48DM3urUfkH9b
7MzXWylEiRSONrNl4lW04k4Lgjr6TvOdYyQcmGbMxWzXH++UFcMYr6nNHy/xmBKW
VbKxm4QHv9gjPPEiTd4yPb42ZrlN78+/gyjZA8Cm4C4yE0wESyZitaimWiQsBBai
jrcrPd2PGc+6zrvvrfjQ5TO2G9bXRCloCYHl0ytcMVXI2Y5GkwDG3xKUy3w77mM7
EqU1IU8qBVKrGgk+VRlPHO2OWk/1xLYx1DAnjy3w9pMYvviHnqy9guKf8whX2kuI
ug5KjbCyHJcQvj0Xu9xnJmHJShRHZJUEz53vZL8G65mobuUk+Gk6J5q/araASgPx
Oy9KLn52r+PapUKVxvCCOwx7YnCQXfv3nqi5tjbKoNWz75Z3Mui+NNT30jc+oxJE
F7JGiTUYYl0nHdbU8KSl+1Ljz0QezqSYdH6vq8W7oTFq4w5WbN17ER3+NiN738pw
OjklPTYnT1WD1O7efYGQCQ9lXNC3jO9TX5UGfrkXFFBI3/csxoIw37I4KF3LqA+4
8M8MPGUheAYNs3gXoMbA8+ghV3zIuxcHvoOYVnokuj95u2bHouHCUoVsMDdxQWYj
PSXfCzlMp5rA0hyFZeXMGVCAmahg37a6xzzC+muRdVZVsxXa6EZIfqmeH1ZpkWXw
yNaVmIZ1avwFR6lcMpGILEF/53bFoUE7C7c9K6pu0dpVqc0oiF+PMdAJgJt0gQ4c
hLqqWjzMgfvLpAJfncTz4v99NPSbZQsleEo1f21gQe9fz7Ycrv5o8Rx6FYuVaA/h
0EZAWInSULEBTd8+RKwCro5EFmcDlCjQ2PtbcKN+y5eqkWJsI+EsyCOlriBRnJUt
fUwNHWd6cSu4jk/s7JDrMRQys4BKA2poluTpaZEfAcG3p69SD1UPCDpnew7WcyDF
iJmNdQEYtCOTALOHgT+90GABlrhdZBo+Tm8QMWppM133F85JHH3+i6DlXjFcKf3J
65jpb/OTjXz3zaJLWsGDxO4AR5/Jeoh2P+/XUKLS8OIhK8AIb14UcpXeUG+so4pu
Qbj3hk+5M4/inUPxA0o3KMUrFbLZTNh3Mg4KRNJgQB+RAovbAIca6n/IVWkre2/k
14/bsU8ax+dFmGmR6FKWeMT3uNrb456cuWNPlZYoHnXh4X+W/rjEUHM3GM53fItb
P5h97YnEH0J+ndWtf4MScTACMbN7YIDpiDu9++eZA/44W+c1lGaGkl0+Mlk9TV5P
q64YEWjd3jBPfjImlefYu7vYgc7n23apvyFTc36B+M0a5Y/m/ChLO1bH3L7JkvS1
j7xrf0BRna7o1VfRwCzPxrLNLOHKUaIJnKOQxUhAjeqO9nXM8okrJOBkuy6bEVRi
DRSqe1PIpEHYN5tgiEsjCfPbAEFSQ51HR6oD/LGzVrv1eAbR04DeH9JEXIbPp4d0
2esuvxhxcf3Gu8tWmAOV25vNfgu0ziVRxqlR5Il+crFlImjrBUisFDEIy3tYhBxp
eGs6oRzE1FTgmIjk86hclvNtk+xysdIouFNT3mBGyj25qParYbm7rmH89IqW+xZS
9t8PL+boJ7rvt18FLwbHmlAV2+BZQRQFQHfW9gL5KBqYSkdxjbmcF5IyXyC8UQlF
yaNCmI6Fr65IuIRvEmJrZLyJFgjba9JAB34K+uCOzljCy+V61isOuD8dJcxmwtwq
WYa+XGEp96ZI5pFHQWFWMb36bkZTyFLwyHAGvAkJz/3MYxHbC/V1u61tig/39QNe
EHS4MztyetVsNwQO8Xr2dnHlOEjc41i5dO+MRXYkWmIHHpaZ/YnL8q9pdFcqXlWJ
IPo8Bf/YugWte3mnKpWFLJ7MWddZjbjMZBtuhmHvqvibzpqEefn85B7V9x71wvGM
qyehXzhwjpnohfpww6mgl8USN/LaPE+AKoS0qx2CEUDhhZIZxGIZOEnNOr82E8Qp
nY77/IU8sQ5XiPPnXIoKoUFej+JJXPHS8Rwgb/x1/RB668v0z1NfrXbmMrqA3yDK
L44B46pPwfX4Wuxk9TEs71hpKIJ1FJmmRIch3Gi8S0JsZOkN7t9G0L5d8Eue6bgC
bA3PoqaXZnqA96JQuDyQ6DMQRYRyWBuqLlI1/GcCDQyQHVNWCWP/TPBI2nalh1FK
3rYSusVyaEBHIeARZssJluVCr0OUj3fUjnFr7290HD103LHbAxzv4iEZHkKPskAB
L/uvIty9SvkMS0AzGkgfTt2QyiXyMNzCqz4gSrt5xQoFyYoE104FUZDKBkLZNjJP
rRb2KYtit5oUdWE6SAGtyIvXhu0l80Kszyl4R02ii2BRrNBnfRv5V4mhfluPVYs6
ixSeIYofVJQKdrpNpjU1VvJFwURzkyAWq3i5aFiZTyyOxkGxAqADkYQstJORsr4v
CuGA3ewvPnV5+RpBrlfhEZxz6bRmAMeL0Lqtg206SpXy0gBBZ6I241PZ90lBZRc3
8zQ8c4SaQXVdO2qTJIdlAcH0Hb7tQbg/byyG8iqieMTOYqNhLGVoP6anA9GNzDYk
LwmpDdcrz3fStTyAHW3yRKGvYKyGmX/bD/Uj5yuJRLOA84kieMWw+gTVVznTvTRZ
b7KGF6ge5NcVc/FSTRLLgUcqWgZnMjcGKycdkb/ajkaYRACYcvmT/wVJTpAtD5Iw
tq2ZlwpUjhJ/6RPr60SxONiQ4jrKTIZwcqKNWeMzGKIiTZ6O5M2b8YbqqhEVbXcM
3AG8xRbrN1Ae2+UZnONEgpIXqRR70OsvO4ZNbMPJAP+4r5OF0Hx2WZVateBKbz0t
zubT3R3yF9Z6BMDD133Y5dRcn5Sr8aUznPfo8SXmBOyn1RPk6jJOWXi/rAe4O6qi
0pYzUUOxgxFsJBh+vk337BAMAejKo1bRI5F5zbtt1cJrpjRsYEQd2zXQV0oEGyMj
AVDd5+mSN5QnWjFQEZy+WYa6oIMaxE/GbTpduFKTHll3GHefb1j+NdeiMjo4hRHH
iu1HVsAyymyR5hYmhoLL4c2hgt8FsmxTrFGVoRo+lqKR9aoIFxwdtyrQS43Gjh/V
+abtA/3Q3tSdFarJ5bBKOEJtlfQSqcEpHkOgWnVNtUf3eMwwG/aE3zE/iJvYk68Q
fyqPBfcj7aJiSTJD8cB2TkJ6yvex8VyRhwKv+e3DB8NoW5KYHhu/wxc3h+Vp6nlb
MkErbTxc/+j/Mp27QkD4X//XhHCEzn6vDJeqE9WUzxi8wgpbJaFY1uNXnZIz2f7N
4iQjwi1+CrRzMKCWuSHXnpZtqoH7DOwBQJ8iIaCHsJ0pwL/PoC3Z36apauzps31F
qPocfy/5ZVNQ/6ajs7dwal18wyFhOg94f3ciLLIz0BBPGcH8+CvvOdbMFIrwrs8B
NKefq8xmakKoVBcwDsxltGHBrZ2/tkCAGeb/8pZQ6CNC+O4VlY+j/7nFIeW+/rxm
U0isICH4jO8TYTPDjfBpPGp86wCtlrDSk2vA1Mhm8OKoGhlG0aW8HIMwgG3LYH3H
CIF8gYlfJ7Y9nZUNmxUkPFlyrKLmi/md0NKmGh13wYbN0GvGnIGMLVxQD2k0u9x7
Lw+EXxBDGu8tnYryT2cvD1F2hZZGfLmktuNlHkIWxwixtXczVVg0zEGkK0Q62caN
FMG37B5BUEbd76BYks6lFA4oFkBqDalwqELiLlTW0VbJD7MvonsqCZUpAXi/3jmj
4O3jTcLq6I//74LAt27soEB+1wjULpyQcPY43F0kh6dVZjU59S2SQpkwd7xkZoCL
xxWXpRZVSjKiv4hz8511h9nhuvxClrzMqR1q9wRpKwl0aTDZ1YsDvv4C+vcn80TU
6pTX6L+kXTgJS0RPHMqixTQacO4ImmPJ9ZDhPKzzqueNqElA9l7rc5xrNW9HOHCC
dPWeDA04La8WgcwsMK8F0py5fNhehoMDk9l0/lKyH+eUc/lr/5honn331EOjLtVa
/Ba23n+lrkK7p9o6sTVSy7zFqPdGiHoYwqc96bz5NquAGYjwgbYdgYzeEerPADa7
sn1O/EYzsmMNOHO+TNwjcIMuHiNkwP8awXDSdMSDkR81ap4JxBmyN4Aftrl1ZlRe
tQwXc3ML1PKXTgft90tUTTrmlESUdJevyOyqeL/GisUDdlUvThwEfcud9vB94CLD
7DvtKFvmKZ4FUb/3jBQ/PSrUAst9zoAHvXl17gm9cnLYx4BN2Sn/5qi28AccQ40n
z97NzEg7dGvnzObjOk7Sq0en0qReyrReGDH+cKAqBLJd1+Ze8sCuk2MzhhIn8A5E
HWF4i7YXJe6MHRfDrBFNG/IMCwC0DUDcbp6mcMRYJ+r3dLNHhgQ9x87y9RJuBJtp
47ccU98J8tNAPDnUYfejQX1yPqZR8VkPxKTw8GXum/udJRJxAHhSG85nyQ9F1oA5
SobRxXZz1zgg9OIPs1HyygzroyQuNJ9kplMhQGGQz87AJUkOSO6pvAb3uUen3Wib
ROB9ACbUPtuU2txtRQJmtj7yHfnd7WnJiQIEs6VLdv8lpXwpagbv2Uh5NlfotMhm
0hmW7SHFnuMARmsIvIcJjWLqRqF0GyefGLklxBgvTZM/B+j8M2N2MsfL51CkwehK
VfyPvbX3uRM3ghCAUYD/4e9GiyY/i9m2ZpJRjTSnALj082KBkNA/EYcdugRBExS5
X4WvLh5skNlw9YPGFVNUi5ixF79eG4PBM5UBaH2fsEL3O0vBglL8VBzvynTpmd31
MYCYeBjuutOtkySvuPyEsopFibID5hfrnLqxWD5I6IR8j95lGjajpg1Q74PHPd5L
fkHDOGOtMHMsXR4AxPgOilZ+2B230kC6AwjIL5GKfeX8bs2uJj9UXJUYEDNK/HZ0
+WQLQZpin4Oe5SzlNG3zTGBKRjCv38IHWfBu5CBT+yGmsiS2Vo7H+Njf3B57TlcX
sPAWXRTPASgB8dpGeLu9cWr+YNf8iMmyULz/Aqg1EGHUC4R/RsKPGle+onaaILu0
GeVCcziF6J/e1JayISLGwQ2DWB1IykqAZj6vfuFER22fdKh7nX/tC1OKACTfp+9g
IyrWaaQHsoGXSNggvmWeYr7JmBabWY+5rm8C++zk04NTgeLfN3O7CYcUkt7FAjEP
1sdFmQ9f3H/T2AqqQEe57f4PupR+kj1FgvWb4VMrYTWAMFlPtERyVNsstMBx5FC9
mnwlq1ewB2VWWsDFXLncc1T58rYtyaL2StPodpAspEkPB4KIi2kcxV3hcyQ5SE6e
5HyfCf4fNBtWBBjDnG8V/JMBKbGmmtl6uLlzV0rXHq5SA/SaOH0Us91fTFSG/B11
RcH489Xq4TIhjAs6onevjyUabndwBXW0XFroXW7W0a5qeoi1vPZPJhxUUcQcfRCD
oMzVpJrjS7HrowAZjf+kcZKhXqb1Qa2tuQUMktLxFYgZDgMTwmsrqYGzS5v1SSxi
JXIzzaCIgX1/C04T7gRESjdImrIFA2j3Ar3qV+SGKm476t7ZXbrkD9xlTKCZ93f/
9pFwaPIZjJw0T8BWcOXEEFo5gnKbqALGUcwsjhj4qkmQ4IhPrzhm6o4AQT5VVfON
25CoaW6jdVjTJHYSeMepCmts/DSUKdqwiJtspDOkzWzxVu6331plnUSCDPCZsYHS
OwGx4zrXAjL4MKsjvmYy4i288EhiD1iIlNgyW4tsyq3EPmIiXcWEoZJqrbAdLRC4
iX6qqlql8Gnlt2axA5vvx6Eb089d4NPu2E9KtRdRgcTpmVjU1QeZuSTYx9EaCSr7
ZbViS+v/Wpma07iDr+lp4JVpFMDI2kqSxywUuodaltI73+jt4d9Xeug6W10mYS9A
/0FHh7gSBiV7LHWsKjaBKnSWBlmCmDsvvZVOPTh2dpaXnTE3+wRcrASIYPHpeUXJ
4uJKeyC5knQy7EWT5ICoRC/9Y2UjiFNxUMQwHUzOLpI381yPLLs/zAc7l3EwSgkK
lumqSi0V6mWk+Gsc+dTXXmfTrjpNHHZFfl1npTgOqgFS278kAasZItZFHkZrjPbF
jj1Xg7LjdKqscWJqyyV5iBKK9gcucyOngOZHqt3ZlhVQXzp3vTwSBViB6AbuFcrn
7EyjE/qXyrrIBPm/KYiiAqEgyvXCkJ87AxxJC4giaDy5oiA5MuB8pOy5T1iUBSMy
HtzRpLJpmPebcQynTsQjBy/pTETnlBw/RqbsBV4gUQt+whlqlK8Bl7nKsTA9oTGv
b+N+wD5ItEgmTXt2GcLF3E19e2L0WRcgSnRyrciTw9paJ8PZ3dB/0ZtJwGkjelh/
nmeOAzb3vH5NzjOODlCUZXV5wItp/xmgDTgzBEwBtwS3c1Pr+H4DyXZoMR0tAQK1
18JbPcLpyHv5zaW8n2+C1wf57+JzU/Kv3/rLU3WMSh0pllcuTiUWl/dalHS4LktN
lUJoUq2dKwhn5Ve1ai7KBdcGgCumffksgIqH8Te60fQqkrRQ6e9czIFHzGQeUhK4
Pj1s+gTadAH82Nh3wYmWJELySnNugTyhbBVPkowx3Aa3q4lGi0dZwDmYMVjdCrLG
qd8FSxG8dK5/u18fTOXj8SjF+rtRYbVNV4BhRJRZRz83M8/uFoQ4AqS6wBSe27iy
dpLSh5mDK5FAuFMpT/PvFH2CPeFMe3BcUwTKeN7BmsUcxFZUBI3D5Q6qX805plbH
nc36EYDah3PnIik5P0bPlWyhFubSTxipxwSfND0xlGSr3MtEOPCYryc3iUoASJ5V
+brEH/KT7qsNxMp0EUVuZ6ExeNFB9jukKeWB/xot+IvA5al0xcwY1ue3yF46/ROU
Ap2BblN5ygrlC/hpJbe/nklkvhzlsICndfDPYvoqFX4k1B/1XlfVMyVAoRag5Ykz
h/myX80KG5joTB+nS6Gh/ULs13pALeE8lajiiVSw/ZQyrp/L9gsed+iGx5LNMySg
444N8nGtLY8hhOHksEhDucLBomevG7Afxi8EyaMhxL5XhliKva1oy/OJVYtKdtlu
aZ+FT3tTG7I9WM6UAjSfYuHKpBCgR/0BKRkC0g5OIETti74n5q8PNET3zdMvLIPG
L4a4H7OwgTG1iV2CDoGypOml7qaMqHkfLlvWyzwr4mu6G8Wsqfeu0ojRFaw8P4cD
H7BcEQ6XZwX7F0ghXxrxStIU5r7r+w4hpNVCBgfRdbOUD1CjB4KRMn39WMPZ3IUa
Cl5FWBeDg+4pDs91IxOZVrLkhQKsr7BZyba7qY557+xCAWMdGXZi+fAORfgPNVho
mVvuFsqBT2ZxLeqz1e/jyByfUKF1VwvQxxk2EwcHO6z2Wyv7dO6hDuIQRplQi29m
0zyZY7OKTgaPI/mqikTzO18Gs/tJyvTK2GNapH49SJAIt0zIU3UVh3RUq4WugyIa
LltVf6XnRB7GXl61WxSgDNSekaBpSIpDVzOR7BmkKrUDknKAoFSgU7E7t4eI+Nkl
Dmh/YMwLjzuX5YSzvYg+ZZKWJ9UPvj1JTrxkMMxqf16zdf7NZAgDUpg0sUWuAhxi
5EACxfwCurghbXrVAg+ctg9bg//8G06jahnPT560H1oflZ9mbU50JkVvZUArK6mO
Gpd+Lc4HD9WfoQwbmDbwKgI9fwflv7orSnD4hGDsnlLnRhww2cEvdwfEaBmCWaN2
lxhQIBIRODV2KYxfeQ+6UvAYQTfTFYne9i+TnqBReeFNy+ReKMv6G02qis0nlWjU
8tUqqIv5YJVrxkyyvFDMAgQNRaCJ08Ji9oWHTH3f74oDeF3NO5KY9zlZ1Ggs8XUl
gXJy01C6FdZh9qEz2fhhzM8XjKBaGHR3WH4x5xR2J46f2mU41boZow5CyJBfLZzW
LxhQxgA8wWxntTBQ2I06u/mKwCNP6qMqWBuAQKqHo7TcYkY10uLy1PouzFgGID6R
pSo3YRe+nh02c5HhCI2vXRvT1ARRwNeTCToqyAzwwE7p+xM2vuY2SJpxJRA563Sw
GLn06TZmQmtStuAh6ffkECNs4m5R6dws47geTqpP5eL+AcUtDw7hyNNBG62mUWkV
HwlulqQb8DgnLBzZsDkYly72hnLzRMm0U7XZHFfgvv6cH4CPFS5dDUNLhQNuNjOn
8yIXSJM4kq4W00d01/YgNICb86QODIJHRBJ36ZMBuWAKuVdGFKj7zPq/K3TPYRp8
g+UWV8gY7D1QqRhHC5q11l18d4Kki3mPm0Cpx4gxkdKh+KFrKiRov+Nr1h05gGB6
sO8R2l7l1h9hK+DzUYa/V9wVeu5UPSiu1cQsMzyM1YejcZCk44fT7lO1k53U4MbP
8tKMBuvLVnD8OMIRyLGc+wP/n2QSeN/wgt5M9iThrL2IsQG8Co2Wmjk9r/Oi5L9f
RT28S0gT4c+RMEAly+yVoERmlUZ5CRpm9Zf2dLkgzgBSUJ15W2cMWcNGS9W43Bwq
o22Dyl6KxfYF9tAsw5m61KxT4hFOEDLOMulE7oLk4CthgFHC5ZdDQ54bKjZ38Z8l
OB65W+CuGwHxUE71a8CRQkykaR2oxyBTFo1UQt/AQ/enBTj9qfPDexxrMT4Ew6OC
4zw9P9nWD0WCmeE5tUiieHwNQXwJEJJnCVUTi8tD/pinBu38SEY6QePEtG08Lzzi
O8FxinM/bHKo62U2Zh2EUvSozHFIKwq+dyPBNZAQIqrbSnKT52te+3Oyrgm0sYMy
ymYRE6LNP7SZU4XGTOBfdeELZC08px4NEIr/wMldFOUJ3JblUNOXykWqKWeLSIfu
qOlqGT+YHB1rHhMXADKpEUpOcnaLvPA0BNdeaIzc0K87GlvPUVTceIN39Q+q/x1b
L2Z/Okf2pnLP52D2vy5zNjJrfMn6NFuOUNQ5PRN+AbG7Mg62yBkHBeSgr6Fun9Xz
Lw/qIb8rY/+YPLXdzbzFlNNlzgVK4zUfWj+Taf+t1DY/mwtahwrp+uBcZP6ijJvQ
QNSpymHJwyYBUr1xF1t2KHzioCwBz4kxZJU6Jxb7sj6qZrRCF1zIr5Osrv5JNa0M
SUkaXDyBHJSkPyvCxLZNB70hhT/733Bk/WKvVecfl5Lzts6sMCbVGT+fUA01JRCb
cAJgQ7awYTVYyOrxOZb+zqkt7LhmIaPd9R6ev/kwOgapvjG/nfL9LDqqlgnKX+Sd
DJAwx+ZuGQ/H40FPh2AUfQoeLioNlN/Hp1s6oaFqQd0WBE+vbkpQlH5TofUM8Mci
9hstSxfS9eyAJiXZKXrpIyFLl1UScCtBE35izCf9Q1fyjSApBFETnmC4j0mjBunz
r7oILBXqmCnlr9RrBAKgyLic9D9Tm2utaIzFjUfuW0PRIpWIfoCILCU/SqwiJXeR
69nuso5V7SVX2x8SIALTEnArm+nEjYInbI6W1e26adQ+IefJPbioAQcXFXkoHbyz
B7V2+JIvQSvUyp9iWAr0SZv6Iy95hDlsDyEoyasvCs+PXs8OWjRhUCnAkEDBOkex
JMulHeEDY7vxZmq64U6AjzEWPoHKMeMUtRLwMsCjNAF5omOokzymVhEqCzkx5x5K
rrG9gMtdVYzaMNTaLEN5ZhV3GHcxKMimNyAwAbTySoM2N/aCQBa3D8vZslpiWSy5
iNBYy5hh04iS3qZ5dg+Gy/uqHFImkgZHieXbhAcr6hHrzJ+i6dr79M7Vuuzrbeo0
KMQuI825LFUsX4lKtAGXQMde0zkeGlY+M+seqpibvE9nK9it+u7kWiEkWBVQXuAH
9U3ZD1o5qlEZ97HwnOeSxiv5/A287yYHbNL9+GV51nnZNFoa1RK8rAE+p1yUHLnv
QmClyH2KpX+CqlXs32qGVmRWgAJutYGJ1rtmMaz61RmYsl1CJBRbXBnQBWfMVJCS
QKPPErNFD++iA086n5Amgm+K/aleiQCkpIYBIYkVD8tb/jS56AxOAx6HJvf+jsgt
YBpbwwmeBE03sTAFhpZnNEwA5eOgo0hrH4ATR/X00Sm+h+a5lsEVhAH+bnEERkuF
tcMrHy62k/+Xw+h3CEExyq33XyixzCASPJo3pQdrhrMq6p48qQLThPJYQ2iUpag/
/dsFer09M2oCi+lGI0bOtT+KEyC77eATWubi476V6jZqAIVvam0rvlDxEzeu2ikB
2DzuFGutNklpIAo/kRJTZuYPjLQywHvRTU5IeTZCXVMt7glO6Z4nw5rcdUORgAcJ
FaCqWVBmF4cjQP9BZsERJdPxErG0ZDDrxlwMfEaCEzi4oHveO8jXH2HwgHORl8U0
D4DvWtNEHdevdgEb8/WvudOzWnF2SsKnTW0avar3VfV4Ev8iapVRbZRjrKKWTnf5
nHRosWF3PorZhw/uC1s9TzuPPneWf1gaGMlolTIW2/5Ic2ireM8nyVjdZeQMaOOg
G0u0IuP9ldsRIcOpfHGflh2BBgGBedl25DcnZtpTKGTVHIC796w5nvrwIaEtPuGp
BiQLzJKwfpQY/HaPiE2oC4JEOwFp8FsBZofy2tN9LAZbNEPtZiyhYpVXd2odoHv5
J+6CAOxpkKxuFxaQ3c0mBx4Ud9PR459kdnE73ZeMrn97+sYFtIQ6EpqF3Rm2Ghko
7ljlXEQ5sk46p7Kj8GB67YR8oQK73l1mPwfeNODmwVCG2QVeN3+QgcsH3SOvdg/Q
AuFdfM02ESFgzpBoxSfrXjEDrzCwdqLbBMID3RKmUmwDoTp/LYvNtMiIyMD1gHjy
4rd2RswhGNIM5NI8PfdTfvuESco9DVoOqvCGDYRKNGSLR1e+kc6NDjdAOPBZIPuU
7EKvj1bfhAn5L0p79M5dfQW8zNbZp+bRfVdiKh/kl0giByiIw+TEJQYgaxcDdleG
AbHT6D2zgC5qJ1LUt758aok9NkOPk5ngqyymqN4ZJcQNBnAIgP4xIDdahnXIxNPC
jLn57nzAnrCA5Yxr4NuO+EuTQXDABURwhBaTBu/gXcSAt91HC/ikRXz347Ank73U
2V4+yPplARNSLZmXDig9VZse5ekFhhNdqzYFUS/Yg79Be3ZYdcmpscUDEJYyZiSo
w1jJsyvhJ0lOUElHbQDpYQHj1bd3MvyuL/dhlFmsvCM0xosiwIthBAF/ertpBFDK
dM3di+v4o4YiQcWgnrfr7IlxNZEJsU8D79Q4wTUAys1pMtpRkqqu+iE/ht8dnaI9
aBPscV4XHqufHTieccMtQLix2Oc+tlbMbGnE5365/vi2bd7MoB9edUWJRmXC+Qbp
6wqZ3H3IpIP8jpaBiFdFVHvYFGH6BdFHt+vD85+djdCfPCGCRVgrj7/QW7K91AKg
KEQ+qe0oQydzlil/bRQFWKxiHmcPM31+GSn4QSNGxqpbiztSpaIp2mEY1NoRofpA
yANRPEdSyChnWsSkWR3ePTMoBjvupcduXHGhed5fy1xL11/d9lDZZsYWG2yrGl0o
A3VhDMiozcCpDnZgnuococym64/5LS/8MUlefN7mLToszOR68vkFi8aw77B1zOJ8
3jZxLkW/Jfb9pjcBuH3BshKm589IBUWcGooquQ0ab24z8qjfHaJKBG+xWT4oyyYT
ZSx8hwH5u//qZz1QJReFrSTZR9RFdZfSL6h8CRKLfdePLzRHpAY+Ia1p8ux4gMvz
EluUssPXTINLxKMnNJAIe8+z+YnVVEYK5BcPxjxrgJWN0B9ySrwnWA9A3wv8DSvQ
vAFje3zY1cucWQapP4mJJdYUQ66GYkdnv7B4zL/2LgWFPuhuTAq06Mw6G/wZqjY7
7iOJaPWYL7IxmDhPX0S+ZjsYvtoDAF4/jw4fgQ5O0ue0WUy0r0Ul9mTv489ZLXqr
1vsQhMQLqpgXNx0hTylCFbgOPVW+5DPKeh28rJbJ+709lLsJTRA+6Sjmqnod0rQ+
pubuzb2otkZ/VI3uEm4VqVG2elCIQmp2QJG3cDRUD/COcbcmexH/0V7Ufyx0PFNy
AZ6CEbu35IgfifRno5NAf82EpCQDTbwPxtqs9tkkiUJkZBxI+mvuyfFcdMMvrN3b
Cy4TrCNkhwmjv6gMI4xd7UhE2nM7kMG1ycxlI8gDnaDtZ24JwffNju+iKCP690e4
SbliiRkHTQiq6+eSyUHMjKQYAPCWjZ605ot4zo5Z0fYNMrYcCkhj1biOBBPyH+/+
6lz3R9i0uh43nRJZtrviU9HmDGspM2Itrsj0p85sh3ZMoNOal8XX1so1IH6lipja
Aq0wj95LR4wBQohSq0AeVC6A0SA4yHfZXwOn+aLQG6V2OiH6qG4L1JLKZ8R7wxb7
PYsnYWKQfAQ3QlNYYibs+pn75HUgwPYEK89Pa0RCBZGNO+BvToXqupoeb4gOpJwQ
+gfQqn4oNboXMG240UyaKQ/y9h5vze5ElRWAeRYnD/SLFMsQROx7uap3PI3pziBm
uPFyfqMt52mhGicISOjwPcUSeT1NHQa2Jtoc49qwZmOx7jhOn57mJTOzn4MlKE1Z
ZOIDM2ZtYktjICQC4fSFbUN6MNQ9oJPj3kixhS/Q38k5QEymK/1MuVmQfh1mdG+V
G1gSi66fMIBhGM/uSaRZCCQEF5ZSx1ewBn35UwNYUweMA0yYMj1P4C6fPyZlL+pP
mvFnd8iF1g91jK/sSATkwNBrjKwDgjHBlVLGrH78EliKPL8zP5IUDrGOtU4Q/pN7
n6cbyszrbNptP63qM7PdxQD/u63XGh5d1Pe3VJa3lM/I8afJHAiXBhnRUrDlX6Mg
1GjITHwEQsbxIbop18a6Bz75xp3jRoAMi8uvzkoAwD+eaUSmFdjM+ReZN6d7DiLd
+zCQxnaj+eFJ8hhrOms50WyObPdlw23+ytRVktkXstjGbmRIBdL4JjCiQYJG2MBq
n3HMi7/aObJfHfnZ0Vwh1Ko0CoaCE0fB1Q0u5PPYvXa+mhqCjjxnypCrNTFJ36QH
2FXTKdXnRoGtpEBdxi08LS0yUG/0sasR0dy8uNUzLm0dgtAuXwuzuxsvryLQCHPy
nYAor53EFFJx9FRBMby6tY4KR03Bj+4NAyKP/OmAn1j2fINSCOLhSPVXgoyiHjg1
9KvY2qY5n7ulIWIi62/X/Hj/ZUBmxKltbBTHj0Y56E7iwGhsqeppGFDAA36ONkXF
5esJAulelqSddGPNxpKaS0+zM4zcxe2W7RLaAHnpkFAGTcX72b/ouWbFj0GBqTFk
ZP/elmmVR4o0D7m4F9obnLbWqS3GS33CWQHSj/pcQMCD+cxl6WIbcHm9GqSpWLTF
rJT2n4Nf6ao+69kxk1N+LLWZu9Chmq7iX9HPM6Zj0K4WUIwxVX9sfS6QkGv2PwKV
shfnQYo2hZTpYiBvMRlpl35N57uXk6Gugj5YKkCtKVCn9Em3JqvzmOGZ1NMljWmc
ki3zqpBKeH/tlCkp1MVtv4TLA+W6q7TLIPn4d2PU4S0XgVPZ9ttcmEmZvoDFN0W+
EgBy7IiT0csbAWSo1ro5PFO60aiO50/SyOT9S8eNTMU7Oet5wRNSupVzwATn5hif
hBmmnV8lUqQwMPOPs/hRnTbCTrA/NQoK4/B0SAa7AocyKEsUQ6FxY/vMlo8Cp7ek
/WrxeLIBmcd9kTWSrE+QtuwiVEEzzXcNlPff5ce1uZ6pYSg6CHgKuA6RGaHkb7qO
22tpkfe6vZpx6N6OpxI/TN55vy8pxz0fwOIEI2uq6TQP1ee+67Hg34LmW0w84inX
6mq3ZbKo3Dm2K7nrZ2Vru1aegZsEUvN+9RFoLo8QTj5yGuVjxSRpoNX/IciFmYqU
Esb98KRSN6OyD78oRmtalBnznbQzOIdd/U2AW/K61pkv0xoox17t09fcqPMMZxrk
SKN4Uj1fpH1XFZuPO1YvNv2lLCx/fu44IrDgKWK3rIWaZn0zwttxP2NGwzqm6C0y
jqTtDnp2477YZNRcBa/8uXOcZyqc8Z4ztZIW3flsZ0mMl+r0yPQxHQG8sesDy2A7
XnbIZM/LVY4T703OmznkArZKPeHv7fsMuuOxlBemLkx9ZkLOyf9jHhE+fIIOerpn
wZcojfvwl3xClp//6K6kR1562omuNEopJqzi5bZo7jnDTnWnkUFUyb5IOBwHTi0U
EN/05xMHCwjMd40Obb59ZFUvs1Ew07Xgsy4PdPBYrTjPiA8zbWu5HXz6H92CUgo6
baH5VwA2nM5+62I+ozYJUqgLvzO99RJvOvB6D3cpmS5ACrQVfnyjHvTWsE2TAuZc
ctDiFyVMnz0ho0KgTHhf/zTn8oR0vtfE7D4kyZBahkcno1kalDPhf0kimuWoEyik
cvuYzwFIGhirTG/6CAFjhwLvbzb7jEE15ab3GF34X4YC94GhY3WnQ8nmgx2cHnZ5
Bwmi1FrdC7YYusaRUjKCVz0qpMcaNq3aMzjewCcOQGczRdwzO5UXqDRiLAd8GRrZ
tqGuLQjRbxIWsS/zprfaa/HJP2j1Uzyo2fyGiePJ9uMp5cPRbCBv/r+YjH3/lo1D
tOxUN3fC8VLVDZq1pjeZjKNfbHaqQ63jirTBNLFglZzIrot3u3lSdfkAVKxOInBE
eweYl7jwp6JcZkgDm8h1SR9d3FSnEMzNxClcif9/TvYAbZFT0CfOyCq4yotShai0
GK7JlWGOcitUN5OmwGPhzMgaXwFLhqWQVIUA0dzWrZtiYTaVOA+g5dFik0hsA1US
T9BDh7IXJUAXuGCd+Iaz/+YKobzdORKnW57crwdqWtAr2gz9z4MEtrc3yPQQdK0l
mRgiaZKXZRy6rh98U9EO/5/ntClf9cNr6HzZKZ3cCVZf9SpiIfaFoZItExxcdb8T
aHYa52EeHuBhSyg8Uh3zp8O1czPqZIvTVkRwYGOR+P5EOeBFwiNiUzFKKm6JpWz0
zQ1mHPXaLeMN3M6auXdmoa9fDxKh0+UpTL35ptOn8XbMEEn2QD8av1xMR3mTbNKy
doITk3oezDmWI4nP8FZeG/8N9pL2KpL+G59cEnQcuokKVGzLdPG9pTYtal3fupm+
5BIrTS2U6b9rhE5sjStctuJMVGzNbtsUkok6aw65vKs8suVnsg3GtqqMr3hueqJb
dnkEuM7bfcsRWu9kbIBIeNVZKkTd8S4Vi4N8MGdObyyjYnlszVDzAb2SFSFF4ixO
WHjoW1KuaV2Au5Ol5I9u+N0E3xgF+jI9RI5Kt+98a/v7SRO3J7INBhtWR5CnJxyc
nbGBZYTfyTrZbsHjXLGfM5Nq223qxDf9we0Ad1d7VIw6/hGSIAnFmebRFRf+p3xr
JaR2h5HU6Yxtj2RQum9Ouo6Yk77RLjlH7dTzgvBFuH2bxjuBEYnAYw2wZdh+N8AC
W+jWmP8XnHQrfJy4DDx+B7T4lO02RByXzpxB10J3KHFgQzKu1lWwuiI6zMfeli1m
i09vBmLNfQhd3D+/LwZovv5g9YkpBtwetJuyI2baszRfs+QB5Ss5CEc0ccHOMEdK
TBrJ06IrCCvX+Aym6/XqfTdfDoTL9DRW8HwIh8Gdtk3REx0kTzkg64jvOXhltJTs
+pNBbjjU0zCCQKugGQao27e4ZVcyuz5iitB7H1t0N0X7cxGzuey9rQCCLQisjZ2p
Qdi1nmq61JfhsdmC4tyB4B1mf5MDPZOo0LJXqupHLX9dwiT04YMxM5Lkh4lV791f
Ke7WtJOeDnPIda2qoie4dQBmvkP4K0Kr74km/phjsgvKpssCulyUu0KRtfvaD8nq
V1qkRFWVwyotP5F6m2cyGGSwqGu1V7g06GbiMVGvQKTqiv6pwAF9EWQivRQ3+Oxr
U4p5JEAsCQkhCUI08DgYcbI+pcHiJQTwNTe5iyWojcvW/ZdnAkRXEz6jmR5cVfN5
C5RsgoQd3QUEP35dbO6n3KDhSQm9JSE/SlnITbO0Sl6x/u57CpzIabQHLXRViKry
/hmfdlqsqW5fqkrpZeiRqoLjZMqQr0FkmkBUj9SERebXZr4BQU4PRAqIMl1XjNqZ
4qie159om5/pARtBCdPHXwbDNgSJqYvKkIF7p5FDVh+TjdspbPQDjFVAY8YPPPHY
Qvw4FR8680keFN6J9lrr3uq/y5Q+WjIUarexaNzgS22QnZqiSrOL7Kbgfj00H6+8
A4YtIgMVzUoA4+Zbyksb0+hsANtxD62dOeZGCH4icZi0iI5rJnWdvLvUC60tleSC
vB2zMTy6Y1Lxix5fmOxZj2ewUgJtOqatireYpuquK2DmzOWApCbO0Q/wnIvabpqM
l32e8kTt25lLMbeGaKiAdNV2kMzIJhmjP5Yi9UJNAHXsC33r7REeIXKyZsD7mdJI
IHHSEHyzB8s9b1DrMpy6RRCW/MA7/0AFcwyHqNTTSpaJM6xqKiBTRWFfjMrr7L+g
mHS38D1t9Fw1Gr6jz9+wPA9LYuPqYWzwmdU6D8zT/XSbpEJ/Q4yG043EzLPVXGfn
KqzrElZOQgT7tPdarVHgGJQFB1fvm8AeIcggFZj7+Rb2m7vkhulBu8ojkNC4asRR
4/bQh/6XwRMUlPuUamjRRql/cpk5HxALLoxH36XOgbPi68drzFdk+0kjv3a7jTKm
USBwuC7I1WYHGbsU4jIxCMUZwf6739STI5pVHvz8L4d/+LKKMqS/RtehVE/yO38u
7bcF7jyA3I8quk6GWH+m2ec+YUdkjzLRCqNx6UyKlcIdE4WJbkMQIgAzAxlumtCX
VSilDjsolVISNrwA0FbFfrHxxrJv/HI/bSP7BRfhlORpbrEtFp6cfjjvSsEnSDgs
4SYs/3e8ft9PjoNDAI7x33lo9QnoCyjXuOng5+5BHdjK1kSFS9mLGegA74V7GeEW
LtnEtRXLTiWjwc6URcQgTlQG3lmqf5OnZvFdqvvmp2qRH0KI2nwZwpJPx4Q9no6v
GWkumhtjka1hbQCAMELQbGeSrI8p62Oq9H+xKSEofbDJspRN4ndvo2cPkEi++p8P
pnsFdtGFsaX4s3cm87UiFl5KnkQSXcyICJy2xKzyuYC+lp7RjJVm7V4eWHs0VbrF
o4s6QXKobJgiVN46pyblggoBxPNZcNXnIGb8L4GuhNKvSkHVq1+CN1dhs+zwOZWb
dBZKVt8FO4wiswP7CPJzXfyD1ESkXcsPjlJMQVNUbNOtCMMCH19hunR8w86SerTX
//A+NbdXevWz+hYtbIakuGc8kcfDIF8i1ZfLatZKmLqPqmdSS4UmUoLHbtSiCdnN
1OnsYVs/zrO6JNLa2+ud2cNfWHqFvLDX1DBjzplXzxvFVu4Qybq/QZcEKp4jbT/J
R4s/7ajIEnRdpgyh+h3OdpatbqAjs+YupaoAr0CJllL4flALfy1zomnnXpNIAXsX
1RryszPmyHCCbzpqlY1fWNh2dvXru7P55bbjZnzJ/zZFZvTUhDOp4eIc2tRPZz82
frUnFFLTHHf9TN/eLjNmZXEIJ7JxNGCBN/CxgexvWY9uwxojiQafyv4qjSzdE3C3
qydFNAhJ12ry6ZsQQ7X0B5ol6QM6RDfGz2Tp5SsIJUi1Vy9cJi7aNN6404z5yQIq
vQKLOdxViIJH5SwP6ifA+1IL2bgtDc4GAzgYEkL1JuZhXQ1IlE1GSVdXjwLg4Qsz
Slx5vBKAN3wDX9WMGQfJ7UPKkaLlJay7XfQ1jfOVXnHjryje4UUsXhm0Qqgdeeo+
lSGghnms4eoGZy3Q9QlCGk805QgwzHLwefIm/2JekfXp38JQRn7mELGQ2wqt0gNS
eMDMXDtVHdR2GWCBpRasu787V676Wn4mUapnpWU4rBwhCE8YBk22zSzg+GqlqriQ
CiKmCRhNVvJRIxoUDYWu5TXMNc10t1t1US8DTBdsHI0nl2XPeQvfOvnIoDaT0MKZ
MQFZtxoDTum4I1EhNrPuSXtTgwDrZGhxIUne+PoZFkfBqsKM0oFMkPwvykBIa9Vy
EDUcYgte9zWojHfyT3Fk6zyhjPmO1rQrDBYx99+gLNM8dGvHJIABz/4RqD28E649
tQfy1/HsF+IlgEPW7t4AsnrOcV9YmvRUfRvC7iZ5bNqs8Z1So036b7PGOFtsIac/
bg6nS/B3kXcr09ph7MxIT35Astrd8fCG2HbsmJDmom3gOkNLSNRb0a4l4JvaGO6z
ag1Cszl7N/GfaiiXbkZON19nYEG2BsJsSHNVcKQDc9ZIZIiMVX4B0N+SJJ5Wv8VQ
QEld2wPEGf0lofPjaHfm5y0Rp/PefPsb8ayWk+eGnP7Txgpxjc5Ns9n9kAvXL/bM
Oo87gYQtgBsZ407Es+jFdmfJeSWp0ZndVyRroTrekb6NXDKifpLGSTfBqegTQwaF
wWXsN6XenGgZo4Jrj7ZpvzXCUqrBNJExMW/6oiuOA7C6wMmm9lIH/rBBBm7wnAiQ
A/KzyncgAFVYU7++fpw5Io3kFlfuVV9mOLR5ORYN8wlEEscSQpxk+He4e+fp7x7L
V8g4B8TfifrclOs5eS8S6OhxhVKRX2WcKo3an2645Tz4kuBobmVLvk4IZWEMobx7
9+t5WD4P/R36gSQBKrlGNiravTXHba2iWjP7iQxRpGTLeShW65HjnCNenxk1mORV
Ws7UOAY3w/Gu0ve7RLwQzasHfnBOA8o07XWmnjxcQWWHtkx2yNlKS1bap8NsRMig
PFqJRQVEOjEszZVKXKGcC5e9iJzZBvTJKijAOGyo+NfrulCw4WwsfEDSgZi+M0Ra
Det73/PxSb8vBavadCiGI2nSD5OciCmFkJa668ZTOvAEyrE7xWn1y9NejHNJtbtu
By5Aqb6TXmKtpuXxG+YxmkXFwAqBak4LhN7FtgR3nyalLS1p49i5pi63zoQ299IU
gD0Wj8ZNqcDiYEvOe6K0cJGzOThsTII6EZA0nQK2URpnpLcxzy6JPwdjzVioihVa
21kydF5UE8F0K24CI1/SBDjH1KvGi8A+IYBlNe6PMGKScPYTjmgC+LeQgsCF6yw6
OreCsclJKaFVTjJ7YoubzXQ6mkmSa5KrJ3HkS0rjog817xaFCNM4QW8iIqf01Sqr
iS/SqziFBFxzr3f7qEK5n28n3u8o/y3Kuxj6UVb8k6Q0C27qCt/P/NNRS5bZe/9o
UXqGOQTU7KwnXgg6jjT/MEsV+bBsf3eqQCNPgm4FdWHt+ADCHiESGxyAfg/2/cp/
cl22eI2rTHaylFReWNA81da/kcem9V7vbRRYccNOc4cIOysuQ8Cj6Jcs+oWr7kso
+G6IIb/nkqXdc4BDEe76PmjTsTEavrrDERG13oOOmotMyHoEiDvT1nftTM803Tjb
FcqBs1Lkv6mWg27SPKlIpR2BLFNubLyKsIKimq9yjTPGGtXkbwIM2IfMZRteQbMW
8xN+dIUd5+9UEb0DsZygEYXI9h53TavIP+7KZLlgFJ3D0ITukhs8WwbIe2jtwFSA
NRWM32nGeVlSki5pwEjrAnoOP5W0RBpTGF0UmZuwYo4nSNcjwlnycYVmbi83B4Ka
hQxONdEhKeVuAAwUC5G8S25Ryah2EF3sSz7Bu5gzkToVRB3s05tn3rLQ3MSxrTE+
5D1UAq/eqcZIx+9iBl5LBBdw4HVAeW8p/kqZDoBDzKyVQ7O4/7BDQcgfWwKePvGv
piFDndoWSK3lKJ79HEpkkjprsMaaM5+kldP36cfeh5zKJIKH1H67XQeB2zXvhGXi
RB+IxwveqmB6Z801f3+EaP2bPyBOffeMM+7m7OGJ1i52rh7GgMZ2cKyvr6VtvGHG
I9gUe1XGwfd+QqlYvSVtTivvVOZghqa+Xx8upKrSJEvgVXw4Kx1IJySbifsbmWUn
QaPE+T+PmLL1kYFDQzr/TyZY+6lgClQPNRV24SfjvvnOwErNABdvv/YetkE342ij
Ohv08x67P4s0wgvWgCyw1rJlkwjTIso0ZoSiNvsy3u41UDEGJDcEfvkz3Zrk9lBV
cp8RtN3H/Cv/AQ/YCwU5GTQH5adggNrpvotAV+rYfewBdo3WeOUhglKoltY2r5Zi
0z3+S24RJf8QVKkjq8uh5x2S3MHTG0tny6zd1028mbxdfD9jQJLnYhQCO3Df1UZO
JCS5+mE1rqSF4fFV/WlJyV7dsb72wketdrS352BjTIrBCIhAfB+PoLvwW4jE7lck
bKPGo0Z6+tJvFIxylm7uhJq67JG7rASVKsuJ4VvOCpGhR3gm90zlNsmL+xks3vwJ
0TZj/YiG6m5It13ZVqRUoB5p412jGJgcrsi8rohSiJXVuLXAdDRYtRB6qBGwdrtS
4Ns0scsOZYAyWmY/ilLPRzA3XtR7NfcCpLbjD/ey3o1L0SjckwTd3VM0I7TJ/Nnk
5AYXKePZFTGpff4JfQreDgMoVE/zTS42KX/X2eTDoIL/mGvZfMg9azy7X0kt11TC
UjJij5YkFKJ+Z3PU2vbH4GiWq2/2p5rv+7ynAbrc3DG50UaKxaQRc0RYSL49Bd7t
DZtW+MSsoMM5eA71VTFSWkcD3/+rh0rE5d9+lOWNT8cGKZM/xV3dvZJoD5urnSB4
ERz6Mj4X85V3elcwxdUrhHktiWPYA6ow1+jyxgfW01Y540t5TuyW354GJrOechjf
CUUarrXtdkALHq/kjKEAAvrV/+NMiCE6/yjbQ1E+6XyZtnvUl2kUvi1AG4HqB/84
aqJgIFZvHtKfFhncgthGncsf0cH8Qf0KI9o0VF4VDAsvzI6AFnxgTCwvj6FOV1sO
sk0WgOdYvKjxsiqwKoAmHsO2Mk1uIjYf+wt7GnTIaL2f2qL3vIjkJF5AyoTuIw1B
+ybLZlnD1M3iLvm86HYY7scp4s4rZpK9ce4jWiU3/ApgCoY8/yruLAh26+zo98UI
1ScVJsr7HWjdJCwCM0d0Pe2Mkao9ERquzg8shnbnNNt1CKRZPEkTz4V6g3RWujNR
mQWCvulOsZmqgUSQNcJZXJ1EjxKvVFtmRcf0O8ZZ3RZ/X08tcLQVDYtiXt40xs3I
KpZZ2RlpfN3kHQJSI+vnHSNWWo0L/QI8wB0+iL17QtBAy/OcZh3hElQ3vUpEfISM
j1o2z587n7rgjqT41Z9VUFLC2wCLZonNK58gT9LRuiruV9qPDc8YN0ITG2ZMVQ9+
5BaWL64CWq2hdVsUh9QeeT122q0LU6GOPO2PuSh+epqjfBNMo2tDq1PnB79tTqxJ
CrCzyD7KFOtufWxochU3o5oGEruro4YL/SzIoynDECk/SVd2ULnTGZpaRY96MXHS
ziLU7hUeXylsiJhjc6LHWTdLXcBZNo2NFR1nWCNJnTR1AW4Py/XV9141EQ5uMrUn
vSGh+dbPf14MVtkxiNExw/WnxG2VJYtrALhMYfwPNp8x+6rWc/7Vj5g4uC6yxEpy
po2XNQfERege261dg1ufiJIh7gnt8wB8uKuYHLiI65jPMJyJCU0RBlzncR/cWTXF
sVrjaWUTF58IQnSlf3goHJzlPjgqUOmzgyg1WNRThb/lPsdQRhmIocDpucvJpDZx
Z/ofJDvi6m5JVfrIUEVvlwLBT3G0PvYJUtmQGLKoitGFmYFsbKMJrvMbYoYYtjV0
4UveyIP8jszZN1JBK0oqGWK3GRyHHcRYFQKIC90rj/Uq12UB/G0jC5rg6uzSaVEU
D2fhYXOS7SUnenJUQKlchL8TpOJwZvxubuWUgO3i8b2p83m7ZkBYLfMaxRA/hNVd
CnvovOJ7NGCeIyL0c+MEfcnQsMJHAwo+XNQBZOusl7VhXEMpQ5c91czHEliZxio8
UrF7zu/QdbnMV4a2K2vsG4q5vLqIblBvtAR6oN4FP6b7Z9EZPdRSQwyxgXp2cWn1
94tbMJzZ3WYg47nZzH/hy+LEJHig1B4GcNXC0kGU2eSE31PvCwyzy1KYMnu5HcOv
+IgQEhaMZdkFHD4M5NBYHyhMxWKC2GofTb26Gppe5Nr4iYZA4yq3eTYyv5imEgoF
YneeNi5areoI+c2uJn/7vMK/b835y1PgkwaDdJS9kBmzR1stnoW5i+dVKrtXVS9z
93GS25HCrIAvJ1Qpoxnsi5KvLmcDGA9hDciTaaXT7spmT3V92aJXUiZ0Rvsr/AEa
zUVEOY+eX4U5ykwaUxvTeAqEtzfKlVSMAhvosqHRI7JnL/AUvkV+KOLjKSFy2tej
KcNYm9v+SAN/R0nV2VtzuD17RguUPsDICCKhfbVmaaLXpuwZE/mWJBm/21v6U5gX
h6ktfIDiYCR2X2CQ1PrT6WJPfsOidC8ANNtCRYqGvUbUVXgNCaXhn5JyBMToGEUn
fe/jLQBVNFztBh07NF7sLqogrAx6LyBZ4bTYbfZGl0XxVv1nGQ40KzMFuQROlPxr
/lvKUtguepBNknDHacozDeR9TY1aVSfXs5ai2WL3ID+GZGbjFzkNLVTUV0KCF51v
7hdlrOrq2Gg7b9WSIf1SQ7aHR0LhtNt/8EEFPpxH1B7gh5NpquruV5H/l2veTp/O
HSTIVQ3qqddXgpO5A1xQ0V661BGW2RdQeztkuClbBgwi508rRrSu848m8BmshsqV
YRyGA7TkHruoJmbwduUoxowmBGb9DU3tCiOyiir2OuF1sDpWvoeVCIQdS9mVEWDm
dwiAH2hwyg97cCQnLsS6fLmTZm272aIAH02puy0MrPBDuZcCVQOpmKliDEgYm4uO
U9n0RA3CsgkwUCZaiD+nAScafFqlIZ60i2hbm/DYWxv1y5PL/CnNw2LVOArKFXty
OEeL0jv9NPvoGn3RdH8qmGkki+r4pqGVvora6muO0dwQ5csUDJQgriY/01hLXPaI
fLkeo+Aiw0TiZV6kZ73VkFnNhJt4TpHXl1MuXZJKvRss4kGc+D/6dyIZAFbK8Rjr
NcsLmKTPc0KbEoswPMm/4HXHOGoM7MYvukuG23vXqwaNY2108egdCMRoRZk0uZhA
DBq+pcvsRfgNzR/ZSm+OKKz6EW8EOjaGBw52a2GPHejZ+N7/4xNUSbFaGoISOUgw
M4ysYyR3+0fRUnaVaaa6H0bQKJfUHC3jyCUqg29sQxsFAQtNv+EEwBMER7vf/gjL
I4VkPQWfydxdc7ShZYB4xM/EOtSqqC2Ib6MZk3dp4MmuDdsKFdgjLc1OhUJkZra3
LgFkndBs28H457ULvxyTPdi+VkGjxXK+imkYj+TIPa0Cd3tciCRB3qdVv2zo1cNN
CkejkrU5vAWEQCmlBu4GTXXLm+ERyQS/okWyGyopguTClJd6Ib1uno9QpSj0xPl/
Q5al2xBnF5qwsIbO6NNU/98O/a5xmdr9ZI2zgi+Uq2zYEaYVPFIuCKh950fszboG
Gyyy58dKXlLAQYiQArcHohy7cm64M0x5ghK8aDVsyFYRteDhP9O7Ibz7txcNtYnu
xtfcMN3t4Jc1ZDzHMYfEhUwnF2M6iRomVlpznYUDGgc6F+/DiuW690/fx83vgjfB
7i5lorRSq0rGD+xgbfYbPBm95vQOszBCnAqlxTW8tFMvLNh+yaYxG5JUJfF+LncH
xKGE/ahGm1beYxs2rj1C4WHekrMenLfd75a+dDNqVtqjM2cX7CyATih7gkLf25mm
JjUksChNxw/275cLwmfqVjvta7chU6vrY01ttmdG7WMxQjtECnvyRYMHThH1Gj8x
d4KJTIz0O/cz49Ii721KWC5wAauYyRNIFdMMCorgj7YIgMsroJT9aPutXGEPp533
tKav1YgYhYivhMgkB1FdRo96TOOF7qCYlTcvtgYHVPkfklNGOPcR4ryAypBrfup3
vs7T9pHkwDK3zBwiQjvLLP76LSs5a0lQ9MitnoZpCUZULj/mNyZfuO28GCRjHbjC
v8mpBxPQalGnz1bo2ifk5Mv/VgnhqZ5ArXVerNz1z37HbWJxIDdEEuBVIL6tA6qD
XkBH43Q7tCJPDEaLDT0ngu5cU0BVR0e375x4Ga3+8Ra2UuswbHrwOk4a9HDlQ7Cz
RVjEs/Xe5lrOEAg6VSl+6LDRBuRx3qD8jnBcvKiTN5SnURzqGTQvbbUAUPXbIk+Z
eKwewAyUHg1FRsqIoIANUrIYSbwRE3N5mIrew/AhBtcqQsOcOUNNef68ixuppoTA
fYXZVL8YIv3Nd7VplWmA/r7qeS8VKWQ5pyAd4DpdOPqngxUv/P4cDe4OIhxV4mql
0js6cuRzrvcizr7xpzeZn8/ubKek8QCQplgQKclW015ypwdP5WOKPxbmdZMaGXpn
qBT1QaTW8cOMdtdVrCxE6EogyKQ+dzBxxC6Ogkv7/lBzMEHXD9q3dLIIS6h6nRSb
8lq5yDZ4rJ/qa2wBrl10FTr6nC9loCerw+bpUSXx3dO4Gf6A2bBjJCAEHBMH4fzt
JsWF+0sPifFA5Aw07f0tre8+xpPxGSMdAUkbIpnOpO9ZgafUzzKmy4GNxEqHyrnL
1RPqsOw2PCoT20WDq3hUXM3Fc/YAdwgYZnA7/9BK2PvNhaUi1O4PQXxW9bJWuNaR
d/x1X5WBaavPBp/s9GJOZ2AnpA4Rj550YIy57loEQdp/EarZHtvHoX/XKD0m65dj
WBMV4LJD+TUJXJ7CB8P1HM83rR/ZLoJtEIA8Y9ZQcfOEphBBcWRSIC0cCVU5uEB8
2t1jIahrdqLpOLQK3ZdkQu01Ck8Z5pKhBnc8fNMT4iuE/ljJmcFaY+1I+Rkd9Apg
dqB0n2c8ybEQUzFRhbgHKfRGo3wSgSXEjHRMYHnoZ1I7jAYnt9bZougYA7ayw30k
XePdIqKFeHVgdmjlHF5hEgufL9EQnuILZR7y1ZWYa9t4/W40f6kypmiiLnWhNbgw
kJs/I90zvGZIPGCrWyCyZ/r9qKygE9ORVSqkpaUCXmR86aB8uNYUOjcq4PuoviZs
TmXIa/6NASqcONn1ZtHH0DtYzdBgHtejbqSegWMrn2OfIt/Ag8DtY53TQRrLa1+j
GHgw2aXr1gCSEsjzt9eYLAs03o3gE6QG3Cdxx0AfJAv+6rw5B1Z7uyjh3Qftjhgv
s38uQhXtc2oi0KKcRarlmoaU67GwVC5v7ZBUlPORhwDmq5NZpbHHDQpTfx/UIDIu
kcFrQ2zVtMfE6socIqA+khpH8tQzSkZDndsYhrrNMrGJ5AIVN5v718G7PNREm1sf
jAgcJP8pcdk1BteptJd1z7tgEKd667yw3gqngjg+xMfNghDeerCh9BqNQ9sDNvHs
PmLDmJdSAO6C7Rgw/XvgoPhWl8Xqlz/IZQd/Bh/Pr+euDhoYLBVTVzPansChFsvU
B7d4XzqXq7/B8jIwDZDXygP1fRhgh5y0+mTXuNlgJrNWhg+HF7ee3SX3xuOxf7eE
stQ5Lgwy0N0vSlCopozD/oBQBH4SfstgQS2yFiu9ZylgQQ9UgHf9gp6knVIoTlKh
ZoIOfAL2tSiXjOsSTnlSW83kmgb7nfrhqkeeVjWEH2RMW990cq75EVX0a5COfRBL
8YqLdlfc/Z8Yc2toFCBXVA0Neex89FatmdQzSBVWSDt1ivsVzb8TZfFhmvWHwjNw
IAOgfRGg0h3n0o8i+jalRljdzYiXXuUVv8ULFmpsT/43x1WrrKnDhP25qQzQWtd9
h4x2rAdTpgelkS+zMmCC7x37PbgEtQZM+pmOEzVtB3/ve0jZmCjsK6oBGZo5uhHR
i4kgMKCR5GDfAUeq/dTchX5jIHU8GsQG++peimaf+agrvqE7D8f366tslnoYdIjy
UHl6xzpxnCkqDG7L7p2F4JVZYz21RNbEyHS2g1KCvnrnip99B8ZUC64I422cKmTL
m9PTIdTceppdS6FsoSEflnKGz5BtCaR2TBJngCrvfg8tc0nhUUNhICZLYhO4SpZE
gJ37vn/wWzo3048cGRfH3gCRruvEiDkf87nP/0rC4DQyMbQZtjArMRCqlnAhCCgj
jBgkNyaQvTfPaf9gbVXRt4gr42mKHz1sy27t4+Quhn0Y8xwXoCB5wDTagsAzBgaa
vkibySQQsKgksBQzzv66KSPkbZ0cM7waf3RVW/sauwbsMVEPkVmDBUXYmUPxvdti
tlSB/kuzuZc/7GwjnT34mZDM1/DBG3BqAyiGRZkoA0plVmYxyug1xYIiTy5I1q2i
xYP9jpuT76TYrT6Zbk4BLVvshWc+81LLsqaMGyj/8bHrNGbEXyquykSlUhgJ4dJ6
bcZhMaaXDLBXjZ2kRun9bMZzW2ZDaZ+O1pqQOhU1cSJAMTPxJ2vG65MvbvbSDdys
+NKtin5AsL4iWlichJ7PeCoTzCotQMaN6PGmZfjajMKNH8B2PIpu2L21l/S/qi4f
eGHI4QoBUw1NvsJ5wmFUbTxDWnoAYztaSLGnHSPkEkZAbfgG/QhIg9uAs6m6l1d1
N+RIDAC1R323IEvDZheuidpag5USYF1OrgyMuqX+G01cJ+43hPIdsRUsxqMdx9m9
L7UAx59g9BXtPypJckY0hXPXGuDTEMdkIn0znEHy7xnvtZI1jBUx9vQIqdAaNjpk
nNHjtx+RAKVXoo3h3BMfF8n3ziBbwq+WNvuXN8McNO+aO0M9gou9zwKx0+tkrd6k
pwCd1t5gEgExM25egS2M5gsmkPC5yMmZC835qRYAL2KSe6Dj4ob/INl91poUpAWT
ZePzBrkAqoDKbfr9zM0h6Lrdi9oHMCKHDi6jXlJnl2OhobPQ6OWAOmzctOOIaQ0B
F3n0aOYSJDNE520XQjcJtbJMewkkx413xmyyx3Tz6YbFgwm+rGxAOWNMQ/RC4V5I
767iGRf1gN4MBmbhnw4LHzQ4fyF5vU3YvgE6CGZB/LjcpCvNRQDewyg3z+p1oSAF
q5KtbeHD1Ko+rVhGrGwmoF+lbbBhNu4nAKCmU2ykwGCr4mcSbFCQ8mcwfPCHjSuf
v3SEuUrQUueDnEDhaepaD+4SYsI39/joRVY/eUXNLLY7JzDHTREzMEPtPm8zIwZL
SuZPkgY8FEsWY6c8N6ImtYB18rS9WdS0ZEhNnAFG1cZ4ScyTlV/t+gQJTjN6532D
drfz26sbFLmMkI+CPRmx/TSaEdaAi0AMc1bf/nEeF+8DJ92s++mpl4YNVxIXCyEC
Q+HqO9jpuqSRzEjWadS63SxfbDZCK7UVCP9qmkzNxH9/oJMCV/YIgg9JVuOl2C1j
8yqy4CjFqaD22hO/llOv2UqswHoaDUc+VTNXB00XkztCzkWkJz0sU/JEkzORZ6pD
OAxgvay3FjA7UXZMwjmy89Tgs2Bp9oTy7Wc2jBEVgoZdZnGsk9Ca0NNK+qyXzh04
HP8yi/BCZwwGqQ6E4n5mhrIvgJ+iRG26YWHEsVvGw1Msv+bPjHiLSbB29oETyG3q
7a4EzaI+gY3pGoqhpjl8OMLdyBDDqAtQa6TbLF64riP+GU5f4ATN8R/PqJJiwq3M
12bC7BV5Yk7kiwLl36pmwojHLWSpfTTP3hxS4iU5R/UPXHjAlbnNy1bfQsJhfHGS
v0AiZB4CG8LYDu8drzSjIETfsT7Qusn7MLBTSQkJ+1UhMeMK7R4b6i9PVZ9Pu2ON
6u9i10WJ+9DyKi+Jgwv5RY9FytP/vXMHCHbOFz6bJcYAeDtibYTyZuSIjXDaUXA6
rSDI8So+RlxFsDfL+HhBzllU/n6mm+tGZyVC2QXPFwI9s4+LxxS0jXoxXUcHGy1H
h2cOIBN547dEmPWTObcAKSzi3DKojCEJJHdxD8Yp7jwwlW6WdjCx24q3mZDAtmwN
lf/5TCVeMsZxuPRKwWCIldCwHbhYDybTe0Gj5/yvUowpdX+0abJ9S4XorKTO/8Ws
fBF0WJ251JIWY1gqNLe7AaQNvrhRXvbfLxN3ThvbX8xEDI8eL5qY+2Lylo4eSuPl
nBM57EOURAwjTQeGL8Png6KI+eKrDp1crDNMxnD9lMUhQw/6DaAzhILCR8ZwWn7z
souYXr8O6fN9ONQ92BgVDs+3j5+fdYs5rbwobgcI30mx3xaKyYoqN3nyyGDWGHkx
UAXfQemxLIPSPgDnLi4pNzFdDqt93MGQHiYyxWDjJ2t7gZ1B+DaJvLYE2QUwLJ8v
CN80bc4uoMx+TrHDMAMAyZGSgUslRQZQUQNieKpcYtpJe/HPUwWe7ADn0g7Gc37n
h9ttiFv+Gu27XH2k6xRm5LvzuqYdpPPHcilgzXLa5TIHf76YTwPn9FiB2APmvVsN
B1qUrSN+84jEEjaO47dT1EOaTM88vA69WROYn5Mz4peHblKR4iN2NNEPRoNOYZ6c
lPS9YBUQ/xYZehTh50MgUMN0IAzV8nBS2i07O4b1Nngk9inq3hwYdQCRKMiXSyWC
J6u9QP0YmGp8AX7S5itXti9DJZJXhis8WH8aEAZqLvI95tqaYyU6arnPWBQjidn7
66IUODqZpVCnA/rTLtuwJJA9nfd9WSWmijmWWSnIBX7FLMdvNBCHScGipVVoKjNR
k/Aa2Xlh/wsDCwzbeIbYkdZ7JJ07FPTUx5cj8BNSIxV+rocJgUDsi4fOZfp5rkzZ
o4kUwbvJ6Aw+z+8si1Ff9DuBQqm1sFFQADkK7x3x2lbBxL8MnpW4ZElhac+mUzKh
7dDvavBJ8YWpOWeTNs1IayIrkmzaLo48CpcDhSzmbD2DTaKQGdMjyeFmT7aubVQn
HyDAZJ3gHyojjMWerker/n2Y642GkjQzX739hl6G3trRAfmVujuSSysXMhr2c6b3
DSRAJ9HrC/Rrz9FudhE9F2cwtitdHtai3lOEhABtAXHo0we/hHDxW3F4nB9ajtzR
IxxF+jI985aD0M/u1z6kebnk97PJYd4oSCL7d6Eq0iAajmI34YEOfowZhD07im0G
sV++TX7sanE90iok2UtHgUyJUkyZn4ovC5xcvUZCfbgwdQOHzOPVr+wuaqwrI+FN
kDBh9+ZAu6dgfQuBuguFvuObJcPkI6TEF7eO8EAhytZKb58B7EMqWVgtINriaWJi
C1mvp2NyevbuadIF5VbFciH0NCuYWZYvUoeVhhIN07EyY7ZDTjertncIfPH/JEon
T8FSUBTCLGDl725NjKd1e6go5e3hyvj+aXp1BRyXqAmmVorgkaHjpMpxsWqH59Rf
MlW5N3K5Z0BJY3AOmycMVd9q0dix9XqP9v6Z74kSz64vKd7foCRSQZYPuavwG5Qr
ZinAuf9pzCbfPH3Nu+dLHtIhUbO/2UzWYkDotk81dS5XixfmoVMyhDyB+YOAAXXq
pD5qAwRMBl4lf8gYeThon/bgzXPpwvNsN8INbQRpX2DE3MvppVnpQQGX6ha0CWoN
OKU6buin3oWqqkIxncVF3FhCi33gH2Fc8sQ1eHYL5zBnRpzVbuuQ+ucH8h1sfqq3
plKW+lpRZ3hq4P7RfJ0ib/wZk0gsUDBLx3LkSjVbLq4OcT5e5YQT2omD0bEgOFuJ
eK8IAEbLZUFZkc0vtpzZOsA3/p7FDsCPWHwxUG8wbfXPpo90hrISO5kSTHhxLc2c
NIlptjqQ2LCRO+54VYwJyHIBpaA7JGtRWrR0tOsGDr2B+PegTEmuPBKT+ig3EvW2
Db5njYLiet2OZ3mti9aUm311lCwh3TKFYBN4DFBAhbBTJZ0UzU6zkZKuZBCu3elx
+4nKfw0rtXUrRLclifC2oo/WNi68XH7DsHNPWPmTE70V3sQMwJXmCR1DLOrpbQ6D
drm7+80b8/45Ms9ElehK+eQOKxrXnH6s6DDiR12Djmbx6Abr4lciQnLHn0YNXF9Y
cGngPxe9WbSYiNhNmOya7M3cnOxM9y04FncSUdg4eg3gy1k+A178/hIDKW+LeAXU
kmAvG0+cDvavV+RgfbLjKg4Kljh8+J8I2TCJ3b9OZ1VTNlN3yZubvefnVYHON9zO
JBW7HuYCyzYDp1D4l+8kBLuV4PnFdPCLIekrRBrVMBqo3cluE6/weG6+ISFTMuJ9
6Jmv1Q0QHXbHoBxKAb5RufW21jwqjjo3euLZxYCR+QgGa9A5eaTEeThTzs9yY+fz
3ZOcup+cU+EPWswYFL3JBTrmzpfjYIcnFuMFVyg5VteOw0r4s2/bfAgv0vCM6Xu1
ghvXfB99giBnwXqLxuXy+auqIOZ1zZhzYWz9nQSn2kkS/0retqvkbYDrXSl8Bytm
wOrZ4XobY4vzcKty7JJM6RuR2yYLwcvdcretrC57bLx4tlXKcjWoVdbUOyocoEpG
xud9RixcW7wuXGPI5AdQsdn3pBHBFjMwZ1SPsclGcBDIyq1ORCqHq6x5p/ALyuhW
/diIlWUX2dQC++c59+WWUFyQ3mfpls87CQD3+lJMC7W5PQpI+ZOwz+lp5oA+HYXK
DS722smMYLNyOLTL89jj+TGf4/2tW6hjRsrlcMHhgT31DbBrbn8yEwlgzkzURW58
+73FIExqd/UFpw30FojRVd1UDqVR2hFx+JRiyzPs6SToeDQc6DOfmZvrEx68xwdl
vMH+1IF+WKDPCNZSS1OxHDkeapqLNrOGKLXMBIG9r41SIp929stUbFHEgarJ8Ve0
hoxg40VzvYct4tYVY5YQuHR1dk5dViGXl/bCzMIFRLvOdQ95mKDEvpzrDNyibFRm
+r9KlUaSGnXjK6NtvLT96Ro7Ar2424ZC86MT596mw8mxgwPrwyhlNPrtag+6Ezix
HOJRu0dCZuOLERpxY13l1tkbetczKebnwILrhsEy6uWnsQQd1PcWvu7dhVum21nd
awCyRLM0lq+2WKbHslP/IV3hrV19cPaB77xuaolMtj47OW9Dx5vMw3D1U2n9TVYO
f9kKt2RJGBWeOSkiLUVs1GcyMhBrwG8Q/BUguqKx3RqZPBfo/tqkq5iau15qHo4p
BBGAq7uT7kvtXpRZahFS6UKFkfjXbtKW5s5e1Zllo6VeQWa+qPc6feTucFBB9ICI
PaF+BGheyD8a2T1jhRX54+o52fBv/KI46gSUAmcBYZMJrMKhKKRXiu/qsfF5YIl3
LmNk/NU2JqMbuC+xsXMl+/9YPgny671L3X7HcL6gAKSOOyXbE67/2zjawtKChaCO
vMnrccfBTJgrmh81pdKuugDTWI82RMFljhWBj2+jr5iZawjeBr74picUYPc/+oOT
pAMD3NDeUyPH6/GHs0mcf9OO800paUJHzzW9CJcdWKkrW7QwiJ+VEPCdaHcdFEvj
BdfgQzH1TAqRV0m5d0I0E4Xu7TZCYq8xkS7P0zzYQfE1/mHJGSREkXF3LE1JP48W
xVaMQxsrvUGEEGwuAShVUhsYXQJeyqz8ueGffe9FvxErL8pLgVDQMqTBb3q+RJ8S
jf+2G3MyN9Tv+FywU5NlHWvuN5U79iHtJi6Y0OSj0/RugrHJz7j3JDF08UieF+vZ
C4GESSrTbblqKlxDyjH7Y4Ct6HHNA6V2gbRNfPPKboIhxBu3gixzXtwS11LJ2EI3
FXZw3h7uqF+lV0QhUFpDabkJuQP+w6qWL/eqCUtkeyv1K+VJBcX3Wf02O79Jip5W
4k7nupAddj09vQoIjluUdsMliiJLLMC9ijFxquY+NTKqVCxc0qdS33pwV1PBlag8
SGKYMMbVE9T07ad0zcMXkRLj3DDKHk9LL82WXmVBZBYx4VZWjYSpc4sVwp1gn+Ok
hpfrxYE+QvbwWa1sDGxpC/lz0112DhawGr+OVaVOirRd/nXXTRm8uzunm8DYe4uZ
Zoe7meRsrSyCJq9O1j4A6G5B0tWOY9JN1TTAgETRKMkeHgFEpAwSULqJidNdy8rB
sm5taa2OH22sBZc37umq/rauts/eW54S4WinGBu9tLvpNaWEISxE5odewbJXcqmP
AspPJ3tCNB/o6IibL0KnD8IitCTAgyM2n390Nh24rUqzKFjCHR5wq+X1jWC078bx
DsKNB3G76aelLECWJgj4cwviVJACxPUVY0+IpPRCaEmT9Stvy9zHKd7y74LUfLNc
vk4BxRvNyjTGpCP+BUdXn+9tFcf0rld2yn8qzlJQgB6pMwVlimDkPCsCTwjJPlQq
n2ByCBF5B6RnP3+GVZACLovw/3snzRdPgrSn2PBYiIvc1rP1yZRNRP/+enefzdnw
R6gOPygotQ9wAzZQcu/iuyB0z3AnWQxX2HQIf5G3neQLmVomCAH40HNhOYl1Uy1T
9mmKeOTjkokMz12a0s4KNiQ5FFgO6+7UEpXUgn+zDBssFpK4s4rTXryPAfdmy5sU
QREG3meZQ/JGOLKKWNfmdlSm/m2/xldc6RyCmaSZhpNZH++GZBCyasMB524PNMzr
H+/ixY3wD59g10wrD7TYnThsFAZ5Bynpsco+bR+7vCjyIm0oSfIyTyuRwG2fc4i8
1+3ODkW2YOYJUDIaeuB0Krbjv1p9i7tSEGk+bFqhJLT0/Jsln01mRM1pQEcbU8Kg
OIM00XMm6P6yp7TNJT56qBVEzGGUf7fjiAeP1v35wvWqga5n976z0MkRGKpZ7Bg9
scJmNP2shU6NZ0qE/6BoqVQcXZUWOk38Feu87ryHGlRI7KNAcLi5g0m+RwpYhpVW
lx/jBxF1VGZvbyzT1lmqMNrGpP1oUVrnQvwn8X9EfFytr4uqleeg89t3sqZuk5UL
J166HFKqWgtlY1nCQPPToBwcau9zbtZLh8YjIdBDGktZY/LOJfwdykmoE/ZMboS/
iNFA2hC3WagkqZOSV4vQ4Cq/cjUXuJ+Hul4r4EsWGPeFMrzIc4AfODt+Mfy8NSnD
9kyHYNUP1poBzsbGta+catN9CkBpmCXp8pWOCR7laUFiunfUhC28FrJCRc78YPtt
LtsA4EK+QVphhBiVLmUgZg7dQP88dMT43qLfgKeIdI09X03WWWV6chvJe+7IquGl
l4v4Bf3iGFvrLnpjcRfp2Y4i77q5GD2VpP9pHOgGQpUI5poNMK3N8JnoPXMLUA+0
bH6zQsXg9++L7sRIJ1nROWH9E2f++m8lsS54FCAB1Z9Fq5MolDWRSUy0/Gc+zSLp
tERlGDCjGzEc32kXjkN/NS9ewgPPHft/FKJ/Ogi5qAOBsm/gu7syXjEeUpDCHEAm
l5CQR8K87rd0NWdN7Z+Td5Wbra4UFObmYevkAdL8KPKZgCKWGEqGRT/4B6Vv1ozx
W0Ud7wWFNikNbUNeV3GcbvdWpMP7akHp7aArqDhnrUOO8ecfJUTH8P2i+DLIb+mn
CuGbbzUwSH4lxDlTDjZvmrAIWrFuerUHeWE4nWZrGghQg7iNxqm5BTbXBz7TKDNZ
pCA4tqCUcUIucU/DRCFyZ8g/vIwdpvBOUpVVWVCFBsmX0ef+Gp1WYE4W0bR2zW53
tEPYQNkEE1TJCAtx5OaLdqKsf8/5wGQYcIiLQZ5RR1H8gfyMbslS6tq3grojG2bw
GdEP9MeMbZy7qnRDOG7f6tWTeWSsyQQmX/TlMMoNBQ7Jitb3y2p0FgYWssvqHBHS
NwqlzoFFH7CtwAPxZBTZgSZp64FVgPoHLUCtx46IVVcIGBn8vKfDtE8vN1MD6RHG
kY8GWcmsrhee2INDYf3dqIiAgc5cajj8ONbDsfNlGClB0ijCasq76uisCkZOq1Kz
uHXOkvnKmSWHGeAfXDZsVUndYaBKV8AGPV4koIGqb4WZtF/NpgEulup1CwKpbEQ/
6L5mQk11j1E+48tOZio2E0xLT+iKLk8M+gT6J4AuY/4qKKUI5Hn28bNogiwyIvo4
0sWHj5dLFTNaVoTwntBjC9+95i1R8zsfk6ROYV1GTJeWXUOpxhFFuj52qZO44sri
S/P9qz69tVfnV479Ig+KZDXC5dWjZ0BgKb7nYXnSEuy+KkpiClp71JiwKpGYpqce
aeactx/LOko5SX8HmHcwEz3dwjiivSCsIlxWtsk6PRqSOBd5OjZAnAwmK/3IicmI
EnjSPh6BCoq67QSS2pdxsm1Wix9oj3nvaLNm3wv190rt5BDB5Z+1X8PbOC1sFA50
zy+06JnVfsL5ku2fvE9VUizDuzvyIDGMbbnwNqcVXPFO4JvlIMLbtGpQoAVttYQA
GZKAYkeds6j2CVRPKQrLisxfPitVC/7+aJZ263wMnCXbLs7timHnAmy5z4xlrSub
Brxsc7fe3gJZtfaRPIAUY0+6SZIGiwitvUGpdTVsWbO2+Bx6oITD+PyLTYlRlcY6
nHDMs+vC2SPMxlaSrrK1zcv7OfeKQs47TYZBjMpcJmO3Ge4zC8m/V1DfQqQ8pzwE
XXB2m9VlGnR7V1G+zS9HFh3Ja/vxZQj+2ItbiCEwUXLmOtsFtXHzPgF5u+Xi+6ih
lia5JVcIhrqJAkOCPMA/mI+Q8goT/fiO+PSVeAlOXQSHYXAqYdVXgJ3S/M3zw4xb
ksKHNdJ8mMdXX/J6D97mDZH1ZmPO0b4HHJCHZODJwEFVGunWHhgRlTifwCIS4+P0
xtol5O+WeOGfXcbFTXeGhU9GlcSRfYhohQHIjf0s2Ny00oyhn2sxVSqtVaDN/r8Y
3PschKd2uA87Q+zsxZYnIhY2HXzpaMUEA2tWTqrh5EIdxFwyOE3pFIwYz9Q5L1HF
G6C52QAwPPs9Q1a154Jjz8VmmdalO0GgTcz91c4lvSnLnlwUMVAt7CiJ9U2m+E5F
DrPZeprWr/rRoFIIQjts7/bDBBezzad2xxcRAvgeAILzFuK5n834oa7W/JH2wkU+
rffkb5uKBOSyZk1eRJc+Y2FJn3OpEuhvRBX96tUSjVElRGUXwVIjFwDim6YpCGNw
SV71QN2NbewD9wK7OVXlw+WcK8e3QwAhkhxu89vIjemCMHMjXoSfF3/6mxfK1UZq
FS9p12ej+tsZ9aoUPId4lSLPKXvK/rs43Rhz3rDIUXlgR7ZH8wXwmorUucQXNkAm
3KyE7tMlmjdoJVc7pgHTFm52c/eQYV7r0JZCImy5j3GgiDQKgsIs7MGZ3Y0TQ4fL
SIKd2qGKu5hYCRc0qg+A6Ji/eay8RNO+NH4tOrN/wDLEebNcFPU+nQVvJhGEcDe/
a9tm8m2isPZdKhvp0FygEPab6eEiHAbPIZ5nu5XULTjPL/DYTEEi4zSF/SV9KvcX
zeK9+er0Okdx60AAmqXPz+iBisDhhpVcT+cQJqhG0ZlsFj2rnWUQpbIxXuR2vWTy
cTDFvdeslshjSGzt27vJjQSsDERDMG2Dz2JU15h+5AZf1G6rENWPnXwAEkcDbPbQ
Ixym0QxW7cIPKttEGgpl7FIlAk6rkAlUJkEEGH6g4B/r3YFRwZzpFFXSgoz9FSh1
JbIt9CbuYWomGLME3+oBOBMZ2iyuBmp8AKzvtY9TYfMYYzdp+LxRdpXTNDDSL49M
BdjMZz1jXWI/YaKMezYU/dfRCSM7QNDY5ib84MiwIeiSq3UW3Vz7qLtYvQNQgW3q
IY5hUQ5MwtCvraWO+6m+4ssD22tpveNs2PRAxeq26DuZR3y91Q48w71Gu/7sOrbb
6sI1X9qG1VDhEk93hPx9wSIdcdIZXDQ36PzHW4BWelgVexY5O0QeSDzO4fKX7Q6F
RMzeoxMRjVZfuGtCYd3Ie+vbnXQvZf5pFtGUM7cz4vmCwQZ19W4ENzfVqxlSMkC0
bTv7gtXNyC2pu4+l4mW8uYgXAikXhLip1NjluGsHTvRaZWFf4o4kGqEFRYtXgxhJ
hvV9s/U2sF64sIwaiMH1Dr0oqGkiYMs/+juV9/p6cnoBTDiaXLwE1Y9rx8i6fxPo
/gMmEYypsZgU9ZCkP+nm0J0I1VYT1M+lbx1bm2iyjgjy+sgzQWemM2zJPe92Ssmi
RcTFGzuQC9hHu1VZ4wfPCc3vsuqqLOfp/MwCCZPQANFvmoFIzqLcGgWbbK90qLHn
PAKZHtSf08FzInzjLAsrkfP7B22QXKkNON4H1K7IenD6/Z9tNJt3/OlR/MoLxaOQ
2KiVbGXSbeR0YP9TJm/JYDPTlURyjPwX4cIw2ki9rkoJ6UWdjhDwQHT5HFqqqZNL
QjuSum7ddi7MzWvrU7SsoNPCp/SwsojIAbm74+ZLlqAdzsqKU4mLQlc619QH7QU9
QzrU0Lzalzp7lPrf4E1t6fNOS78jCn240Mk78mMP8csfl0H0y9zm3W7OhJA9x14A
y2+s1zQfRPm+vddspk2Cquk/3EFv9ym73oqOCdSe+LGeAFmo4zVpk1dgL5z0t8hu
Pdh3yxwXsqF9sjyr8bh05iRoYgcL4LRWaV/GAFHvsymiZeLMbMFVrCVYf9a3X9b0
6obVe6go84DwpT7UyqFkdLA70OVD8vt5iotnXEIp718IF0vziJXBcr/pzFyX/7mL
vL6SjiqPkOksf1Bn+0qitg2yqmXdNOk3h9HS20CAg2zf5DsDTH5F5ffhzMPB7NSP
DPfxRNCYnS/TBrrudyaZ++gP9EpPxbZVYb7dbH+iMYM06LalWjq0LVMTO27rBvZ1
5aYTc8gjnnUBLVePBSmSPC7qk59t/tTSNbFe8fOcGvYRvwrYMj9AR3REll7dJTzW
jVbj4vSQ9ARJ18jbscffQiDpttIDRklLLcNPabJG6/eCPzfVy9Y+V5XUYQO2DJxp
sioO/iQoIXnN/ITHMc9E2AoydsAQwRu6yGIVU9tXvZL+FAdh4hcniTPIDn+jrAQp
NHE4jsZLrGabFeNJoNkAGFjSMKuyNZEqPu9IBJeH/gSwdwzdE5aFLSHhv/ZYFBnD
2RwAVuk1qPTwhKDuNvzB6ucwJlcGVOMfngBxLTj1q3ytg1aKekmTF37cth4ucAD7
meJs+wfLR4LTou0ugpiDejBYbCBOD2pauJtpw7AYkEbdXWFGw3JuTi5M4ZFTWx11
fYx2zcBDgncX5n1SG3yO1GTcn9KT4yff+pvN8bBF23xDLBfSmkIwGW/MGUD/wp7e
k0lUIpssK8aVtEGLn/R6Qe4o7o017mIok+xMeyTRRQbgLpkko/SkKYpA/r05S0If
GTGV0JR778sUE4QLfh02H8AhgzFlA8vYrfgLcOKvae5dm/MJv/cGebGOC5r3LAI3
9I4AfmMvtLHkRU1HWphKrkOwiCuS3mpTOMT2lH+kCG71egqotOQrRfHfUy4oa/+W
GC0kb8Km2DdAocxt/BVyXV6XXxmWKt/5XaIDmkS4Tl89t8HxkrnSvSyNh2PQVTCp
phfY4EF1/y1h5R+fNvAAhXzzH9R3DyMkkh2BZFYCKYSTD9V2O/nc4Xa+OsbKe+yI
/fnoblCRwj7tpltE8kZlNKb6iOAwYx1D1hcV0NYbEnsvaFPemlW837DYvXpvXyHI
+/eg/KWXBS+IE20lBn0RAo35bGCjF8F9AbAGp/waWd8IF4gy0BmA9CbpTDNMlifm
xy0fjjxrsB0AAg8y2UFZ8ytAqQaV7l7Mxc2XDhYolKdBKM7+OHBQMEaTdiZ0mMpV
gsLZO6fS17Olj453pr8NdPYVn75d+NPN2IDwvuAB0nuORn7x0IoVzzNIMLGjsBou
tk/YV/2LyrEyANz/R6FJnfahN3vMnpxRkmtw0rku03EGqbKUFkTJhgrPuad1qGoU
ExPz4DQxsCOoPiayiERkFXCC2zmDyL7taR1BsjjF6eoDPEhZgrlOw5H0zGEa5TAo
8ItFMwx0w134vUXwYXbnEFguHkrkSCHe02lbFBRNEECGsLatiqPp5SfsOKp7dlEe
dOaG/kyU1sAgVJ1FmyNuilU4OLltPCaxc68pdyv4BcOvWwsUjnmqD1dsBg4/LB7Y
fa/dFbLO8FIKW7sLBAWruj0wVHBmG4gZwChdB3nqVQnLsR9h8B6f8wnCRzbbJFGA
lvqLthp1OFdh9O/G6Zq+kGn/Pti8X/tBl3s2OZswS3eNWflhtlH6j6AmlJf3803N
dXmn7CNN+8pUvLQjKI9UrcnqyC2yWk42zlW5pJeTQTiFjdVqPl+mZo0VT1iqq5yL
sCCgnYhOlvT3SKH/ul+9W/kyVOAlqULbNDi6j2ERB7Zzxw9GZhpJGM1PRt8+GsNm
DDn5J6QmD/6f5UqqGI/HjJ8vYE/8mPdqPzyXJSzEl/3yFxUma3A2sJiH5kp0uVKl
z6lNOYe1Evlmebp8+LenHiTwUmeTo9/jPM7HFQtXAOlANxSxkblCb0YqQaT+a6a1
qugro+CbCaW7E3JNrAu0Riu92/qnUwrUnWax/q1ahMnnLx1a7kKww5QG/NXSZE/g
1tcMXmtUneQ/O1NF73fgZE7PYnNKUX3DmMkCSBmKgNZHvNMpG02O6HMbG111Lp6w
TX8eldStpqG80eHw1g8tCGjmE3swf5eSxkU51hOo4O+bLdl1SB0/5URC+khsphXQ
3Ani8VVntgWGOnzVvT1puFS2jOT2QduY1RkQre3lH9F1zWNnAeZc3cViRyAPrX/j
phiEh3V5hAqEsJZcV9iK8xvn590WvC67Tz8RhU2vPyEcVCYTjsVTsfbtADmv+hKd
dTs4SsoN9kfMxOs3CMNctnfk5LLVHgV1Ft4JTYS2uONAqTF9gLoJKJ1qMrvOZPNl
kBzk8uw371FtfLLL7BCN7KJ5LnULxnwkfLm2/2rgO+2+4H3zrPgJ4KS+AfZ29FmY
zxEPa5fiLQv37cdpyUUnAY77LXxRzBECQF7nTZaLcW2ARhyadkp24j1qnyu4R6Op
/hu08OoWsHbjCmZIjBT1w786uVViewWYsxRGfsPiqxOjEu44SAv5/lGWgJkHi8eK
cm9gxOxWgjWFdPOQyVVuA3N1mGogJzS0HLl7y18LIU0V+h53gLQeBzyK9srAQSAT
KWKZFVCXAxKVZn6xL29E2/g9ZiJqrQoaFAOHqaLDZ03FKVMBRRqZguGf3B0+S06a
jo9ah4aJAp2wJ2aO9KAXpBKkQY02EpP3jjdKsQzBLgoHrPQfxDmhdmBWY/I62O9g
NgZGO47zA0ldpr1shvZ3gIQ1vHAz+dPtTM2UfQjj9PDXq0NmRRhQDlSEm3OOh+xL
dGQvJmVVIj84E/Z5BJDis/g37PkK7+zvEb5tn1neOHCcJVAaL8bUnr1YDji+TDDp
FB5fcMzknRYQINmLYXkrH+LrLkm59pRncVYdlbIJDi6rYvas5xBRc6PFnrcQxDCR
zg0CVyq68K+lnLiXawoAwj3pv0gKtOXp0m5zfpWLzKYjC3Mt+xL1otBmCvTMXOg8
zQZMcxN0za3B+atAjE1Svpw98uP9qOudVUI2fuD9Qpn1aCgLTUG6sB2e4YvQqFS9
GHZRjFxCrddmqZ1siMkWAVC50od5Wp51LegHQgKanKcKLkfVUjU7kpJmFVnyv+8I
sSHL+BBmbywgdL482oryWAoA6hZ6vyw7Caen9IfZv52x7Qz+koqIc+DG01oasiXw
uXhupTOwyAwa416GprOdyqAiEtH7yObmfvEeCcKsA51xJX39AyP2loyk7xYzQsmC
i0+XgNf5NN2Nog4KAeulIanA44RNHLKAVHjmGuZ/orKOj83AsoEhNB4m18r/XjLB
u9NnyE5ogd+zKmsq/PO75La0ilNHWjvZlqpaJW6cmsqCwWPsKjPmxnDbbH3s9TBv
JEJkfDQNCehULNSwr1ais5oDqMtVoA6UNcCuxfRNKSHxjbHMOq552MzFeVp6KXit
+DjvlyM0Idd5+Xhj177KcNihR+if0KHora0Pihine2ugqF4yGdmrkZFjWu9BAvr2
GTjeol/XgaD4lN6fDiYRjFj3PqdcXl9Eir9iG4TqtACK3l7DNjjoxWO3mG/gcyQE
N/puFBU7sk6iyfudlb4J/ITm+XT76Hcy7xqbLTOLG533K+aNO5T5Y8hbYyQdN9Mg
ak8S/oSjRl7an1xAZk79TiHjPduL2lKMitB9FRTjwKw7AT+U6ht83dxj/+Hrillr
Na1Q8VQ/XArWOy8zRimjVrbJWeP/I/t4N9MydDmaigbHGX2guRWSosZT9Wn6RFYb
0LyE9ebp1ak2EMInG780s8l3UI9v34JP+5vq12xcM1ikTyCfohy1U8QuYR1qkokp
J/iO/dS308oJl2KiNVfoCxiHPbzH+Czy6VMNAMtm4zt62NJbFlp+yglrKAYGQXUD
tN4WreoWwGhqsSm+RyBgUYf3sqCqdt4JEtAv+JNUYhKJ0AAn7ynXPBY7CdUBse4e
8oM7U03+Pm2jNDgpCmcYdCIFOIAylCVqBRJ5SCXzFEIBM9mQxQsovGTF9Zqd3Cox
D4QYTlT/H9mpZ1bhWYrJICZXcAPLL1RPcF+HasnOynPZH1/uVYhnkZaYbbyqs70I
h2PjzIe8YXXSGAYXYj4hoqTbUFD9Mqe0N8iRtDS5FhxBhvd1zSxNZPcLcSMyDK0j
vhoEuyE2ZHpwpIzMPzZutZa7AEMUBywXpe7f4QXSli2Dubry1DCpIt2IXKKoJK2p
tZutupYlAc2Fg05Hb/aP5E5MmiCRYCxs7HEEs047U8P0QshbFESGBgCk4Lhkc0Up
hiRHR6y6jGp2MESP/urbFQeeF3Q4icH1qwk688Sp1hd33fiK1ccFtCRgbpas9afQ
LRnbinz4kgCi5vUod8HCfoHfZYgiKiCiyOtnCp3Az827lD1CeySW8LjerWHaMoxX
vPPH/w261ilyu/GgI6/s8UQmQl2GswGexb12PYpxYQFCxxtLU3IlUTMyE0gxAltk
V1rYvNiyKa5gzv9rfCGd0BMqZRXmfmdnY25q1jeuprrNukBXqHQrj4T09HZ5sBJq
6jRNkdGIKr72sNwTlOacfJ3gUMamx3NLSTZ90Zkqkydyq/Z2Xui2xMhCcgsN2xcn
YFuRw212q9cMaLadjDo8Iu3yeDKS6l/UPAy5V6um2U8JU/hCfDDb8Dzfyxu4Kdx1
cU5eSnEtQoQHMy6OYLXVoR7F6P/3ZUWXPIphcukU1qeVM+IaEe2TzWn7gUekw5ew
+4rFYaeZLhOCW+uxMF5a7W32Q2ZUjn/RDBvjqqZ4BZACjxLOFmtHpbSnsWDtw/pZ
EeeScL1Jm2kvNoLRlrzB2EZKp7lU2YkHWr0Ouzed/38PyA4NPt44EcPvylsolHw7
0yj8NLSeAnVkygbpcM5KS342NXoVsnfyPYCVv5AVhFSq3kCz09rDnuOlX7LJIYjJ
+qxYYfnsuCh9/MnkOeDj+JK/jZi4OdohgnYrk5jU+xyeSIR7W4QeM83BPwZDYE0I
3mWCwsEl/YKNaTsQDofLcJzKQMEAw+BsKnh2MIwx4o7F++gQrxxKtSEilFE+URK+
i17eUljTw02qWjyv30Hn4eIFmFw/ItGYyFcS1nxzqopUK2DsDcEGGfN2CL3tkRKN
bK+zEumxhcz9RN+mUF7R6bYMehkexeaJoibNylGUJ9bV+8j7MdKJSc4r4iWIZZEP
YW1o+AG+dGSE76YGRm5jl4swAaEjOdfeu3OY2iLvImr1E9R4GRZo7k8IMwQiIUpW
+eU8FlLpjpIKdomtxvfrOPDrmJvnejKwDOcSIZ5kdONqMzJgFWvKyQVAAxIvXu4X
MLqo78bFNQI5Mbhwb409+O4pTfDYYbYRrbLLNIrw5LR6r6xxJzlz6sUpEjYPvhOq
SXqb3UYXdIHE5Pzz41/PCdQwA/VXelwpyblUM5rOU5h2q/dBqZERY5Tg/HgIbcZf
p1MYPfEgoXRhdet5/3KeXJ4EGM+CNIFHM5II1HikH8mjq2QVu8bRKiRD2hG7gxuG
glliimG7dCftMEVi+F5QbTlBA6HcyFCwbdVsJEmEx+VM2ipFpYIpck+HUJ/XkeSh
6nAxQG20MG1weP/C2IV3kbX62XIyKf8Dul3E7XDmgwRNcqi5nmrQNFTBiwnJ2Fw8
DoUGGoWB1JUPykvhCy3szrlDtVDRMRnnPW/mF/orqHy69RGOk/JPUE+5ksJ50oDv
0NDyqNWvT0G6f0Jil3+xVLCzLK7EpAW7udfMHxDEqtqHHRNLlo7ntAeW1zxlBkRe
B1Xxq+dFra1ZS9IB53AAi5gXfIfiZ1Or27QFcRlChTxdgqiXa1QcGrtWOrULLj5k
d5WeT+19r9pnZp6LOIXLRi1VTHe9d6+qNL/0qHlNVwY/zz/FF22oIS3oYZ3wcZ0A
3MI9oYZQFFWVvoeHw3Ab1M+heHtJ4s5wfEb1uVFQwQOhTHUYHMzqlDuv+5AtkC3c
ki/trnSTUPPRpj7gfV7ViegtmI/M+zRs/6Q3UaJSWWY2nru671lmggNmxT1+XuzV
4RduGlmy90oKhHYpBYpP9GHr+il5CqBXrF1BWWmVVONu9EafXLKBfszMN6OjjGfT
z5bBgrRN6ZxAUP4kbyFqaFTSeLqmnYWLdyDXgeGseaznX6fIJ9/7y+Mn9mJR+tU8
6Wyz6tKFyaxahhCNEgqWJu0jRctI9CNr2hOk4Fxa2ZFuySSvuEuMJhWg8QAXdKZE
8Q5C7BuOoKNnQNGQ2t5nSY/hQUsYtMJosQeeGEnDs7h++d5ucWsUbhAV0YkRpaKD
BRkG0wlZuvZ7g8GwwaoTj0R9UWGiIcLwsxv3mRyiLMraHrlF9DzeS2eF7Ab4wATg
YVtHO3gqB1BZPdnmo1F+VVWeR8EotrbSu4EybMzDvaw6i52H0JjzOJxg1FdorIgh
nVNyIDpo2BAvMahXkDYd8zsMTjOSDzGwcAzb4oYHw/iGZZEtuL4LizMvg/lU6WOW
Ktgoks+2hRqqyd/N6Bd74V8rIUn8seB5aIJEi+FN6TtrIK+0v1pqIhchCV189q57
IOMaJomUBx79Lp9E8EhpI78Afp+MWp0t1E/JYY1rAyDm4sdnDkd+g3/ttBlh58Ow
XUxkuNnQbKkDJyfpdfXWz7+QFDk1a3KPEInyIU8SQaa2ETMGV0NLyadqt4dBE6cn
HCyRqVYc06MwoyPW0FdnorbxXU+o6iILdpCcfgoPs7X4cXDR2PRSSrsXDv24ZsrB
ysyWKBGtSAOYVueACyCRYYamfGB2D9kxTYmAm98dfTkMSnXO2qgDsO9BXRB3jFaF
cKAyHxZduZut51uhxe80k2Bi+rp90gTlblzzQR52ww2G+YmFT0eMWZ5mKNIGD1Cu
v/wt+vk6MeVqYOpDTM4rgPZOZj+FoHlASxbamqzRnQe7AWA53WkQ4Za90DJMhxGX
RbZItG56Tyue4tDcUcJZIKARpfsz2U/+7758F7+kfq1tdQn5ji8f8o4vD1qPse7f
vH0rNF0yct9X/LgWushu0A+B9+UoMwI70zZAaLsQ5rMjgJD3QvMKbh55v/uNaOed
GXnZ1fC1o/EaNIj7xNVS/YAp/xgjh0J9anzyB5cNxXA6MDM0TYPF5nEDjpC5LqIc
XfHjgBbMkWITds9aYGPcOCehtt2NKRF2jOy3Y98m9v9urWs4EZFYeraEaBRxOnD0
C2NcD3zL41owvSTOFPazRO5WdWdqYgO23GgOlam2AEwxZyrEGkLgRRK7zamr7J4N
Ng7CTowninW+wGMdAwW613IXjsEWoknvetre4TflA95Ib5dyh/KAg24wSN6ddxAg
JvBsyqSUdDgrtqDbYj23/SC9iNUl7BqI2iytA5mjGPEaVMgpr5J/1egE85Vz2dDC
y/z8zjr95qGfmIjlV76UBD8DPsiGjA6MtZPz56cIIp5j9YdOIq1td8bh1+3Qu9A6
wZoL+5diqT96bf6Q57+yZHioMowoxuV6w9TUYwjTqaQpgvaNVyWwYKhgW7UiaUP+
F59KE2UTdmq0ECG8iqEjCHSg5EDrZvIdYKGidZBaHgxtY/rf7U6AJgsqgfMTuWND
dj2bicQrU3xR4QRjx+gNjFZ32IHYdckk14naCjNH5rpAMsZZ4dTCjAEo9GbtJ7ic
wY0n7z0ADXILLcKhU/taQFPuaLqa89rbP6fllXzT5yZllEgGSKSa59TRiS6duphT
aKiQ0lT5Mo0jHklHp5IMj7/lhTamGLzIeZvdhSHgbFtGQyiv27Kef8ix4yB8YOrL
EF1k/5nnSsHnspxukFwGB9TK1kQrw+/X1OOAB8k6AvKSlISP5Df3IDC2HekoVQca
LQX4kAR0ZiRxOO/Ek8qnp0ZeiEwRWK13nU8jNArDfExsxr4t9hr3SYQA92bmlBMB
qsdoBMLAJLa/Tr7U5YqDwKSkhUg1maLrJUOmVXcHnLsgpg3kk/ZFSBqYTX4gRMal
5iwPG+5XPib+mpXTk/hJi/SY+uT36Yx+kiICPwfWLGA9uhw6BuJj0z8qXpVjOnhk
0zD0IcApsGUJPQhHbZaE+0bqwTI59LUeBKkgn6uwT169I6ggGPODo/TwSJ7Oiy94
IwG0QH9xWDZYYGm7/AJWk26J2+3+yFR4du67moacYArYH09swWf0M0risSLacqAl
PtANFncVDOkFEhrEk6okCPyT0PVBK6DECTXh8eE6/c7TaGIW8t8ZQH3tFj+ppMbu
L6q4wfSqrpV6VF7M26ts66o/gh8tH5QQZlIwuLggSjoNNkSySI+cJUOzV+56hYka
ALVOgYYay1+ogc9xnVLXfBy9Tlmg5x4lvnUtA4kkmWpvPevJKnRxbgRorgK6IiGr
O+9g108aymaOdQJkeIjMkEfQvQiRj99Si60zYG0gcfpRcnZny3POlqqK5Q8NE6Zz
pjTttanY1SLbjRnoEQyqMlw0hGdd+/MC3qv8OMX8AefRHTaHav6lPol0L0kI31SB
KckpMBNxitl9ACRw5+zPsiR0aEPQUEVoSg+qz/zb4l5x3iEm6lYxnVHc9d2fTy25
4w4W/VJkGw4iVy3tp/MtGLSK6n9JzXGDdNhodCTv1xtbone2GXtb/R/qDnR4kVxh
RCXTTtdjlwN8EANbgobyZDOk4auhTvkgICxEW1GMBDcvO6y24caAXe92si+K9G8v
y2mBtLMwzKU4mSyITIW7Cjy4+cHPylqJllmv6nIGpt+TCag4Xu1o7V5iyTn2VkQS
RNNXq07GF1gecYmLS2D2BrOagFroTTnkw27P9Kj8UseJ8OVC23USwHwowiAj3JuV
FKQbWUg7fzj6LWJ0kFChvp7PEQpUUzlbn3vpwbDgAwGIkdYY1dwmiJqd48q0pQIL
DpG3cstFKPlixK4QOf1pOzckORws0obTjkYCyye+OKQW+LwHoIPPRUd877vFrgpg
bL5prePvcQxKDIw3/OWY3aRBZ3B/1iDZIumyCPgipjWf56dTHCCnW5qiShUXHvvC
KtQGIqBlrtXP/CmUZylxz5CU+MQnZKVB8iz/HdFAKcGclR4UjxbVMtn5JfQvJqKO
vpM6kNoIdB5uxC5vZdKJmbZsKu5qHJpTUhiquNG3N7Y9letMVEelO76UrJ34HsRq
gmZBJmGL7ME2m4IZrovhuvfFk9F68NqD/fM7o+YrVP13tEONeVNtL9t14Wdni7uQ
mgy3Fv1MumZT0NKJvQVyNOSem3mgVQ4TH95z2xNyPvg20mnMakbkMkUMfG5hOSY4
LjZKGqSaLkniKnQbJWJsaRLLFuzkdd7IFidJwW4q970+nq9IuEAYK5wOXDuLpK9t
B/lOUtT3Ef+i5+9xDj2H4gqWXFhgr77D6brr4+Py2qelqCn62lrr9rUXhomTD+VX
4eUUkMSW/+/WGaHJ8kRNts9rObz0c7ZbtUvhkVfqqUTWwx9qbz1H1Rd1WEmI9/Tf
uMtuYDXExlKGKA8CoR2D7pGGbpuuayVGxRAYnOvm3XVCUiH/visoiLCEe2tlq1l0
geFNspqgYFNiB3YwOhzEIp5qhOrOvv46mpn5FHTryl0PpATynN7JsJCl7nc9jj13
hYV7NIdmZGVpNvDn+Ro5raRgMtd03GqB7ygip9/otiP4BlBINynXcw51uTDQzT/E
jd5AMBs/0wGf87J3qbKsMy3FgIdK1/Uy7Q/qwTP1Rn3IvWqh72pdD+l32Bzw/3zE
tfY80cPYJ/bbHgeDjJGR6FLpgxdOIJf6GAkFdg1kKZxo73LqHTV5Rp8/Hk0F0PWS
w81trdNd+JrKb8atlcHIWNRzhhdeiNn00UBMRZ+vgOnvmHD1qZUdSw+kG/BwpG0p
2pM06wwS/bwxwGpeViZ0Xkc+zjOeJ2yPZU3s6bSas0Kp8reLUsdcPtQ5tK4doL1u
GTmY18YHM8MRiUlOo6pG2McCbzxi0oMenn9MNoc6vZimjbrZGTU7My/Bxq67owmf
daSZgq+9GApCvX3kFCRBn7ZNL6TwXs+ddMqnovU9kyzv3sKcUlaCzMktV+TgW9Ec
bJLRVI+3L3gTSDM6GXfne0/M+ybI9IMNehGYz0T7K9CozeKpvgaZJp+OYduy/o56
Lnt6DVSOHqBatUPQ0IfbEFt5H6w3PiGzhfSCU56YexeCl3BnNd/QbQfOYVggg0Qa
ZYY288enpb+KeQqw2Xd4TEPfpfGsXro7Y2XvxAK8oR4Y2pgbk+dIy8RmYKdouWOv
HVJ6ApDZn4ck4EZJiD+YLv3iahJZH9XO5f7EtivwBmjlH5aX5zR60XQxAu6qIAX0
2s2IwLv+7s4Jqwfzri1TUrlHWP1w/l0A76qX9efgImLVQaRRlkdQUJ+0UxFJh7IE
bPfnIwjyrJXKrBf7nKaHdHTkQA2henWH35L/uJVFYqpKE+FJMSs91K6lhusaMImM
9tXBfW+sAG6NDhyMjOe+RABr8S5m7hnzJ28KO2e+Msj1623MXRiPMslmd6XXP9hx
D53zX8dx4YZzf/2GBl5kyoNKkB/DWpZfWPWYPxt98YixbK1vIB4vQCvCMjn7l2vA
kTzo7Aa1nnFX7qb0nchdjmv4eORgEtukLU/DXAU7gKFySyx5yZdFqv1+T0krx50M
K5YTs2LcD3IxvEU6+k2wxMMGu3b74mbDlAz0ebtFqaAfKfMa2ZlckOILJXE06AWt
if+SQn4jB8X2+t9XFGOo0JcaQ0paSWgtsljVcQNZnte6hhhX0+yFTVIZx0c57wAU
iEvL10oO/1qQ+FVIPjrU/nKsS+EHQkPKmDr5lXsMiELEdngDYgkac38eeY1K1Gsg
yvovlMfk8gbBvGLaxw2bYsiD6eXJVYL0CrrDfojvkI7IFvV0F2BbZq2kePbnsFba
AECdbUbJ+t4Jawr/mMcC7uZZVVS9pX8eaI+rKXQzM7rw1+NEtANlhMbc8cfG3MRe
/6KMnJXI7q0cwELhYifwK1zaRc+f3rr0sYiTPM4PtIz4OBWHjI4CX2Tkg2i/DxHQ
QPI+aK916fD1sC3ITHJSv5fBp6woAycp8Wclv/CNn4GSIi8kTyHlpJ4NjSQPvwgI
7edfDwMdeVnHfZ2m4+zWgAc9Ty5T32SaKKzHN9ve1aGug/lStG6ca3f4dzn1gsUA
bdLuh7darH/ALZ8VRAJLI2+KhiTJHsLsNc8BOaiDc/N4aygBpokB6sDflWneYsxi
7nIX++cyoce2ojQ9WbXHZDlYCjDYUT+Yg9tUraaNxAhardEagszJyvvtR8KxGguf
Lt0ZM8P6wBlbsEjUWN+c1fMc1rlTU4TpkycepxhsSi2aruv/Y1+CG0cj2/wQysKt
tUr7wLeTMxjtbsyB4kEO+FNJOtHcsYVVnl3dEVt9fb3f7peg7GuNPHSMEhulEX7c
5AvfOQ4oEeLmChwW+f47uWm7Tu6xJRQ1QdY3kOlqmVbB0rDPQ77EO9lt4Q1Dbzkq
zAG3Jm+STORpnj4QQ5uvQAZJ0/AQDN00JfqDBzzEsr7lFN5pIkUXVioU2uouYMz/
y4/8CYH7C34B/bMBpeoaZgD9A4Z1O+QdYUC7kdXGGxxzj1gP5Di4CyNtLdC7JWxO
93CkextLxx6icYMLZBoOdbq7xTwAfIpWOE7+mmQf+Mpf72dIDxa3Mn+4ZHab8Z9f
5OwuY05+uBj0ao07Wze20cbnpCjLEHU3p1KzZHaQczqt7ZpYQY/x20xI6WnJbs9C
bcVG05jyXZvC8CyEUxO7kXP1oaDUxTgwsMFIA1w63ORp2Zoi/FfAF8qBiWDCMQUE
R3UXfDkR7KrsPEABQcu7699G9+S3m693x2LFUKdvSWJ16ygmJKnWRJn8yvkaJyIo
ImqCBpDWq2rdhjWs4Dx3YPGZIkJdB2YHsiUS2VJ2YJyHkr3AJ1alOETpqrFtAZv7
7avJv49AQvUV+AOw93k90sztUk4eCTaOpP9I13Lkba6otJ+nX2tn5PJqAkfU5R2n
dd0yGaoBAA/arCuu1wk+GA+ca0Cb+VfRuN9/QZYs0URisN0MlNmbu+D1/HyhixB0
8la3CV0VaKhYQ3eBt/N8sLas2wYeOzh3CQXWZQYGpMlDuzuQ7oPaAGKTV3bph5N7
P0zIQsszp/GbjnfgsQDJGmMJ7ChBdTHoQF6B3fIppM+ooe+dsWptsbm1oSZX7zEq
m8id1JniHeWPUGvjEJoG0SDvoyrkwMLwBENwwys4uhhTXCL0mRauhbciY1tQZm+t
tjRyuO7lYQo/46W/O0bnXihr1yJHDnpyl5yaf+t2dd5ocRuLgsaE4QiRgVBfakuN
MpxO1sIK/zXQlVOfn5sO9awu/Jfxu4/oIHWceV6ZU4gLDHpdYOBVHNZbvUc9z/+s
r/Yh6G6M/4QPsKSO2uo6Pa8C6JQD/o6MWOewIClbycB+zk+eGEVxV8Z9H1KBv/gw
b7X3setBg7bvGurXxwscU3sUg23qkILm+AV3mHWqCVW+v92E7fiqbTfzrhXBADjk
evSSvE7EHXx2Yk4vdC19C+svp6PnXYWhbl/Ujv+EqLBX0h+LfApMbRKmfE4WMuRA
f4QL8c3geC4aMRboeCv/+DpH9eVNGDmBafM4DTJyg9V/yecx3BtMNKy2s29hXNmN
nIlMKsyF3Y0oO5FGefqMVMbUaLb5EpbrWyC5xZZvUDpf2z6bnJzECPvaZOa0nB2E
kY1Kfedl1DB2s9LE1QGlqNHDHRgvRT3NO+VJ1irS/CM44t8NbJsZYq4DpPVtO6vO
TajCHv+v+o/WTg6Wp2K37bhhaFoUSYgeAgEvfg2ghCrWx1eIk7lc2H/4mzVktvIX
gjGbtiXMg/pTSu9b8VcnGlQOpAEh08gkXP1zr9VDgMeCljcQktouNZtw7Y6XpN7V
wCCFkMEiw3iZVBgnmh61z+P1PcQtmCvo6YyotWr8kzmyzCHdNnf/jbvzNqxMLgBi
GSPXQOBb7pqWnyp8KbKyDSIFax9sSHVp/sG1FUlabVsItksl9zg9nqBTTlpb4tC+
ZXGBH60WFGYdyfv+8vMFKIue5RTKrcz3JMK6PnlQZrBKiRi+SKb7BNPgk5njV1Mr
lOtYs4d4FuttwUpjgy+fEZse1W6EKOVkX317a8KeiuEJ1a+3PrSdG+QN4qawoFSW
8sOD8tlXLIvhdweqBLG8OcyGXgSwBeBiIHDlRbejuF5aGXHap57+nlYFPc73ah95
fZ2glaxkUJCj8u0jG1tJXRUnamwGvLsuaDkbOui8xQPiNJzA0TuCGs7QrGMxmNwo
NO19dUXnJgZ8ebZHMYFRFPaaUXcmeKK/Z9sJHMPnw6GvLwJilQPBUoKpgc98Vu8G
2KkiHsd8GiCtjaRY10HeD1ucADmYeFdsL+kiHJzBPEuFMQ11Qs47GJYuSiRv2VDD
MO4P14lL72j6Uy7x55qK22an4gTr/tVaBh5Te80sZLQmh8scI7dOH/aZpqVATfEw
6XAPytluGSqy+u3eHpjzKNs334XDsDA386MImyhpT78NsCs2Jf7OYZOWLj6hO+0O
ZYG2nD0CgTUrsxBR3drSvJ89+4Z7khtPqz1sramf9uJs5BTeG6Z9ZckAHiNTYYS/
Tl1pAZl0EacIFWwJMx0Ce+sMgSUMbteqMaf9+V0ScfZmjHvJfqTb2X/3DdKEpZ0/
+i/u8ZMjf0Tms+n/d71pR2eNG1k3Z2mCQT5n/nRHVDqrewqKOfADWE9SkHgFRZBU
YNZRD9boLeoAkZ+zQTDEQr14ZLsxfLakz+pFsEIUtWALH+nAIhCfouTGdtKrEx4S
RMzp5wAfUWQByn/yFcN1bG4Hy3gKY2h4WzKWYW9hSQYfcKGayyRCqFv+8M7eIqF+
pYXYVgMS2WFPVDRuGe3w0klI4JK1NuFY7ntcnAa+P1SB6ndUi9OEvsdmoaKrJjex
yad6K4Oo8MWKuEm3YCipU4eufgGsUsEz/gB9N8QiV6ZlU7GZsGkjp9/p9gf09S2C
WMKZaMSBsF1w/1sg+/JlsJErZBF4fJgvdl+RxFNiUUQbCsMaZICoNVcDlO+G7Np5
VzoHiqfZH9dXBPefXjrS3fKHIFG22rCKtBix0A5ST4vDrIBTWIXpmK8hvLAESrA0
TBzz6nKo2eEb1IxSQYjniaIADN68Mc3KG0yHfDWPa5PbA1BWm62LdUK+mD/eoZxp
k5bdNU57+joIWOlqkuceaMl6yp30AtQLJPFivbfXRuKZ4YFaUnT/6APuhfQEKLhq
lVMjg17ftUgJR8GZ2aeoPKuK23uveh7IC8tHZ+zTkfMEX8SHvEzTISlWiDVf4xms
8Bnmt+ub2BRe2lTbsByBEgEOQuHXbu1Gb2/CQfZevlr0SdN3EvEVyvZqSneiuD/Z
6/sqyl1YjPFoB+pz+cratZ8HIhG71Vlf9VysQ+JvnVvGTEN0HlofMc+bDUVpxqz9
dIABQzh4mQWFdHoqLoLkdzHvisXkBygGqu5GRojsg2PWCtHpiGGMp/UQWDYOkp75
hHxUQyxsSlgnsX6ujAbtPSuKkbKu0LVfbDBRJ3yKZsXJBD4oTdSWS/wkAvYG7EWW
OTNeFjMrk5mv90SWb2jQ3QUv6xkn3S/ql06qr6ML/KFk+jKOr9nbdv6F6wgXzonY
QGXQhnBVtvetZ/ObdheTui8Te4fsd2so+OOwyN4Jizbr9pDIGLNzBl5rC7fZcAb9
gwZa28gc718xhWhHDDEGQLy//DWiTb5G62jXtV/8gfKKx4tFLB8e0CLJqqABLT+C
JETUbCm4PY8yEu2OWEojcDULIM3yUB5CPUul4y4XBLNuvZu5/6iEVD9H/Y9QoOPa
Z1fSbY6LOef26Sl+UsJGu8fUYJx2kk5fB5mvrKxT6tE6+nVn8sSYrAxFJv9B0KVM
Z38Y3d43Vifyxn0oGaioN+j/7yrZT0XIKKCJehmWRrSJ9hl3w9Jx3y9kTm86uwk/
9qscUkIw9qX5aVhZLlT5CKzD+FSjbmtHDmSrDgyoqsnDXqwXQa1hflBQjDHzS/mj
vIqOdrIgcEdZjBNxv8jnrjb6iDsxR99BRMMEWwgeu6+QLCWTMM8k2EM4cVsVJR+Z
HQLefoOYMzJ2hmoAW4tfUo2kmLzIO+6gHhlebZycZgx9sC1SWRs9bUFk/lnie3Oy
AhJ3W2kn41OAFUSgjY2kp9KRSgh9u+4i2IWjF+/oxPOFQ3aiphQDC/nBryTp55wa
dO1jqXBhbsRqJmHhxHoj3crIupjnn8uoraajzUcbJoo/w+MuSAtA+WfbrVJZ4l6C
CXoAq+2sxkjVF/7wtVAZr9qWOjxjVNGgKo6+KtvWZRYf9QCbRSamElA3MiQ+sHsN
HslsoqPjp9vuO3KeGfzBpnwKsttrrzlGKuVwEJHUnknZ48zaXI63GDXAgZhagW8a
Mgb3EPq0/0OO/nAI828AiXlIVWmEbxERww0bUZRPk09MG3/OZERrltvtaZ7Zn2V/
myVIngA16kmuBNAvAzNxv1xK+Rg3E0KyIJB3kgOmGhlXjMk3lkvE10wwtYCOmrOc
rRQ2jz1g9Uan/kz9IVEPVDIPRUZT3f5V92VnMJ6BDZmizZpXO4Po4nUGdyyOXkr+
Wl5GF00rwuUm8Y+sFSvWrOst25uPvFMXzwbTAH9jClyKHQjr5DHesyuUYWgdZn5+
2efSBu8lX6LNjgoPSW7mjeGsYh98BZfKO+VdlFrFnU4NoCVe5rgJYHOhhOLwB3rT
MbA1rsHZ1qHbBNuq9Wkuva6bnUjI9g6krefe2Y8az8NyMoSOqNEA1q+KVagh13Gp
nKm0ZQ3/OLxfkWKPmGAYdhbBm5LHIURuL1o4piKYU3RX51ftpMposCWEzYdBn4Xu
spFUBJZhAay4N9aZNDLA88TLeKr67sK07vLSPX/B50BIdS1EgygtN6xfrWOQ/C5y
vlAeWs4X7spFIZfOxkCmvu9gB1n5SQMh8PeiXqCli/cldpQOowxR18sipqXfggvF
NqHwraSWIf1P1kMel7FyJ6LgxTvkJK5RuORQa6YyPvg8fNy39zBZQkGZ1/SdhIOH
ATw7l2Uk+zSjwI6/VvvLxuE64Z2y0ZCNU2jpvx/NbYjGG2tvbRX6crcgi90SscqY
uhb+5pymMWTbsF2rguPRxFF085D/AiEVCqaNhI1lkxqRmIE2OQP0RSUxt3NVCOTm
PclXATjxpAIjRDACaH8cHP2UTQ1gmwG+DpB53zB0uVRd0HonXD+07rpt8ZumqAMB
g+2KvsjIW2xa/n7DryqT4mbjdTEc7QHl1zkzuoG+t4ZgdqUSAia44osFdCi9eXQI
HCE9McyYnc/gQiSo3DWFllC2OKP9VcLrrHdiqB7CF6+Qhqq0LkbTOGEz4giijAgv
wEP7cvNRbu7K4oB9gHnHOkCMg+BYHDngvELnyix7WydI8wjWv01Mj+F+GdN0Dgcf
P1Bcb4vSie3Xe5j8I/1EZlHzNR8DW8Dp8v/x7/vkMsWIyH6YmaIZCLV4ICMRN+4U
Napib54FLxqnI6PZ+oc6jIWmEvR5G3r2JasGwvxcAMzfaf7erncVqOfmZApUcvuo
qtx0ZVBanGfRIognWR1JEy7WdxPxcc4hrLji62M3yZNOLCetlo++W2UVJNqCj8TA
bFtO1bA9fpH9C6h5rIMF2x1vJW+ZWW9we9SfiOJtnT+3c5SWi0qc4Y7eXw5JTReR
g3duImeZzwknVsThtPaz868fZZGCPxByEGfCbYVRSQ7SMIdW0pfN3X/TV8mIvwJs
CfEkfR/UbjkMqS3WR1EK+ZBrFfpIH2Sm9ZOdgVx7UDYy6jhHy+XFKxtVuCS6hcBA
EWwOLTxJieObTx/4bZ0gFYZxDTUNRITwDqNEsE6YDy7g8D2E4gTcsSJsQNGvqjWn
AbqyDKDiOVfvDVmU0JQr/qW4yrW+oPZq3F9aVSk5YBD9P7uVc4ENWDWJpYraE2kz
wUpXLRlbSqhqwEo0azMwZkf7E+gpn0g7HdeNDE7DwcDhgR1k51tL59dH8JVc3Krt
rXSJkzXDqnCYZ9tEI0Q8SqbUkgdff4TD6s39X0ZIu5STHB29B91W0q9XIASaxMB4
Uq9ezAEatnOdvwGUJ1nSQxs4dUNJh5w92D+lS+1MUALNkxfiRZJ5hFieYVSjk253
ak+Mm6I1Qr0M3ANWgSUjCR3JgzaXrw9p3LxMJVZkctxtUTN9C3PsL1C+OtSbZdkD
J3zY4liAtTvQzHuDSPRXXqGuVdCfceokHoC889DFc1Dcw4i16WCfrvSnAYLpW07C
gYC0JiLpwMyvxj5QoA0gda8HJMeDGbZL28CCb8EfwwyNazDA7iTWOpkZg6K9gwpU
1eMct66ABi+UgzTD4UKT8Z98psY7KDfBTtIqJcI7ApVcX2gDR309ihQIjxC8Q42C
nGoMzSPOiXdgYFTSMDy7qa9bCBTt+gmaxWRPt3xCcPILpp9mXTcdelss/leGDdB1
aTFcy0SiXGCpUkbPkPykjF8a0nRdWr6VGjEmNp3oFa5/hcRT/F+PZUcyDXsltO16
RaHt5sohUoWdFWE65+qXWAHg7GXNsgkLiwZ6/mTz7Lhp2oRPD2UGIbIiLhoN4cU4
JWTo2RK0jSwXxK6wBxZItpdAjNcc1bGOCQjqz22wTGyzu8YPSQ3yVlI/FFzP02nL
iPlC9RUEyuXm/STcxL+JFedN72BWOvl/qi7u3hzyRSrqktDHP+v3w648yfiJnpC+
Gbf5zryFU0mgOAvScLV+/hVU3JgkTOQ6IS8bSrBTk4aUTbVqNyz7GGiBL2/thd41
XF0BzqzFd2bvekSLPM/YjheSnmuqrT3obmYq7SpA3gMfeV330ESSCMZ7IbWg+lnN
Y4aQ8MUYLIPvLT73DrlJyPdFlJpI/x3fjw4AWJqoNPe1Ei8V4+PhTdMikHeTWTNR
44g4TL0O5+RwXfgRmZJPkkILgZL0yF0Zm7EfDCJh/cv2pXQLELxxaQ5QI4ZamFec
TpNlG92L3zOuF7tSQHUHL7MaFrVDPIdNoUJJ3A7ZomAcqx+pW0C5iYdEsHJrLlHE
Cr2zOMenYEv6QWcVwtMCNoIhCAoVhRjP0gse9XnMj/3MnHlQpab935J4/5D8RVMd
0bc0Mf1LUE84IVQM+nTGkSebdcq2sep427iWaffpLM6aE3sh/U2L9sVyj5AODdNL
8eahRHvf4XpoQu16RKAI9L9cfUnqomXbgTIAiwjZnpCBwXnj7nwSlgjwo269cRh3
YsctIwliiu08CKn76m7JnguaeS9f3uYX4eSrAeOkaLinxYlRSsejl3ej2IHT+l5K
+YasmTxFCzBw7I9bC4cC0v2rv8E11oA6XTeL9J4K7wh6W1DYnbVDnNV74/SqdJsS
5cGtwVO/04yt0zAgqb4SxHDT1nkzI7QiSM21rxYDynqYc6Itv1Q+w+mOK+IkZ9FC
xFsThHnp4KNkWarPqDW98XXVB59ftgdjiDG9ZyaXBTeJ0J7t4xM31h+DW4u/87HT
FjRpczxZ+qm6Rh6Fbiyd2OSri3j8c708Yrk+a3ftGIY7Fj4G7FQbDu2JdlFWDXX7
Y5IL2AoMq5vV73F/qX3gNctV9pfabDuxoV9WaMRd5JrY76VXOezMDbXKpY5RPt16
9fLIrFB+oXcWOPDlhW5B+DKeyag2FmfCm+9zolTVUTdCyUrxvfCNipDhLGywGx3c
gdHzHXOr8tSuZvLgQ/joqQz7iSO1JfL5myXj0W69VdU6ziB2hcbREizumAIwzDg7
T4c6lXb9PnEpxjlwsw/K78TYd3eBE83lGz2pOvd18m4T4zsWr2/Botf6DvqsjqOG
owDCuaAekikeAMVAat9LnpTzVISNy+6Q11bLfS4vG8SIgWnaaFiagojfrTX2szDk
vRMeriYjpYFrpqDi0GbC+Er6cSzjFmA7z+QyT2/3ufCr6r4TGH8PBT3AUJOEuPMG
JF7wlzMfTM8Qarj1RIajjwKMK4fHCfDtHtx1ML2Ur++rKucf68SsHPda5VhIjV4H
1Uexl/dCKNmTc4L2n19ttbrMrngZs4Dur6dPDyLD5bKKGnSz/ZZr/HO+4e8TiJk5
n2Xs//yIpQttY4PqmkLMhff5flmB0QMVL5D3LYe0FlJrgmdU3YuRSgaV+5HFd/T+
4OZdmrXGvEOdLYSFTPA6sW2M4JLN03bMdvi2UGps2rwiyl/R/NUhS7ZSrg8t85gh
jljK84bovMhUXPftcg9PlqjnEm5GIAIWBLI3+LatebOz0U9c7dwvDTrMTPQPIx7p
7pRnNgjKuWpFHOuZc0aAKBRjmNGdF2SoehJjEzJdbTzREQjoTzdmESBoKEXvlORr
jWMJGK033ctYpLyXeUtWXQZSZoX2XJOj3RiKaRBuTyzcMi+XjYr9L54PLAtlIaBa
pHVlOOlqzOGMxIj1nnE45TXX0CbOWLJF78hvCl0ZXSLaat+xlETu7ZtX8iKzLb4t
eVZC1tVj8k+u2M3Wxam85cj65dGeYUxb9dInU/6CV94ToKcRaUXzLf9rdija2xDZ
qhLiO/DGr3ZGgdYqdIv7JkrX1OVHcxtz8mr8OaAAmoNFxaqZZ7HQswK48wFJRKwq
7GO4k5lNjd2IvC+J9RZ2+03aqfmO04EUlsuSpPCLmLTpDcM2PFmTZMuPiKpUg0wO
zWjOMqIqdCvdctSkPBdQvLAg+pvDz7lsnhs4rrE32SvURam+J4/dCWfqcrhsIB+g
B5XQ140o8fTYn38D07EWB4eYbEOtCQ4pEJOxIG+dxDAy9xp4HmMZKy1BdT7Ot7iN
ybFYCySrdnMKYNjYvvTkYJIDkkKsysT1EBa7KCcXp59f+UmCYxCD1ziREBEhmIXT
MroYKV6EK0WphU40eoHjLdfWGmTPTcce0QmbA55Glm6/tDnUncxzWQ9s18ajc6L/
Mt1OGIveRng2c79r9pZJXFItLhlyahiqk3psD/6pwUrmKcCTtzRTISQeyDEfQFnE
QBP4c+LaZCot5iz5dnNK1rFtMw6AhZYWfSkUzhCgeE/9uyMmalz1PoshXaa4xOBb
eWyOzkW57gy+AO6Ok/ciyyr1EelY/0fc4fCrBnTKbFGVKiYo6twi9eh6LZx2tL8s
sGg2EYL4I5oHAymt6SfZiPhbV3qInFPJAjpcaBvxc9pDcZYbNGJNdweVbCTbfNRj
XCvrzd3C13SBelEfCwQPLI8kjqceDO0V2ugxLt/ly1wPhcJN1PNB/nSX3hOsshl1
AwrD5scJQxLxtN1/rhrioEu9Fa2UiGcPVKwoQ7JIU0B/zHPMog39gVK352fcTolI
JvyBz31Ut7CxWxniXTNrHZseFkUHowSQhRFkcsoGtpsG5LeMLoH/yow8khfPpRru
FWv0ymwKZJgRgL/8JeWSpsBtCf7b/uWbcKWwVe58aSQepoLq+Y9ZwBY6L6ZPmjT1
lvhxPde12o9DSqW+vCV6FbgLxkCbIfkJCwq4CYATY7nMAq2muFmR61io/ATNrcGc
Epm8yPRkdcOFQk5cXlMTon0KFLeeDU8MnGx/8mbCkV4UUK+NUkuJv6KAg6p0in94
1mzdDEOWiB2IO8/BcpXPdmU/vhIHRDMlMHStpMEbmrR3RSzCOb57aCqAc8tZ1GvB
LdP9PxUTDVg6UW2tfpzfYHp01jVgrHcRSAXabtC6f8OzAAZt6clesh5uvb7Xl3BW
uvLE0F/CYf0GtDd/fYcCHfUBc5sT7I8/I52Q++tkC9dFgFOHSAcAaGC6T4IoMCS0
t7+FpsYSsaz54im6tHEgcKi1fhXEbAKvsrpsbZCX4bGmoq2HZR7FSEApMnZw94yS
sZEHCyW1sO+b1EPlzqcS92uZkK6CqzdaM5erXbimag+aVQN6od6o4z3AwDj92cGp
3qTwCCBV/nS1uFyEaepTfRu4r/VLQkamZVolYwaLKte6fGLzic/mW6vGFlF9yXj6
06SENPSwbOXoEwJJfeql+2PAKP33pthfWuBXrVMk5JohSgEW4LMr0fLnnoUO/WGk
ToS/RTKckSYHrghKCrRzm3Lua/tttJyfTXZCYjIENWr/4gIZ+ZM001m3egtkcnTf
OhURChP7WkJlaNwWUvu6yACdw2D7BKJ1FRK2sunO9avU8le0+p/sxV5F/Vzaibf9
yxoXWoKBvSd8yTogg/Uj9jX/Fp8eSxKaf9eFYpVAsvNcOx72UCHjZK6hXbPUT1Or
5eSAtVE/P5B2B+ZUo9ZU1IKDCkIJrbVILzMNTQfI38sdOLpnWtw4Z5JJaZNkTtsN
SKSaAZvLe2Y5OceUmlGBr021IOUIqDoHWi8o5pYAZs2rZ0mT2hMe1YJqtH2ioLj+
WYH438U/7X7SFk3ATqx3hwU/ymV1TaVlL9yb9AJ/b408IRX2k6Eowz/409gm3L9e
Zy26mgoHi1xaSwcNUuxSQ82FH8c2cRMJGLWXNEicBW1PIdRXjSQyDhA897m1GEdR
MEKoQ1NgQniEjmHUS7owkRP6oo87yADb23ApToQr15Xf8rlJDyBatSn/ZxMEjXzb
Hb2UTJYUUplEK55Y2goIcZVYipvGKDsTjve8OuY7XB8OBNYInsOMyr0RQDRth38U
Lc0AfrxA5icwMo+8oiV1bvMxguGV4evEHMk5WfwWCsRZy4MrbMk8ge9MKRGg/9Dc
VtpSG7dyqbTmnBsFIQcTYyDr8GTtQEb88EZIS0ZYBFllvzD/59jcvRqvIOxGNVJP
9KDfp8Q+JOb9M7n0r6PMpQaANRHMmQF3uSEdrAFenNcL0lD8XehtQs0oUPUDt5on
24YMWAft/IpTnVmpP8jEsbKoSqrmFej89yjsvgqg+GgOa0cOEf6zww4PUfTlRA1T
nnmXahRumoukB+RBJTLorMINDBcBwPbRPGCPgycS2k/MAJmdXb+WRGu47bMpp6rG
erY+6EK9O8tq4HUHO5XgeTIU4dFlmyEkImsZaO589RhnkB8/IbY5zRXZNwd4CbVR
Bk8lbXkzSa2wMNYTnI+WBEJFVK90mG2n/CMe2Amo3WnjHGTPnXnLIloqBT7PRzhJ
3dC8TcJR50UvE3s/qDEn006vZ3VT6KXc/XK6137Bv1zv9IzTJJODiZdujUyptE9/
ZytW6EZtOy9K+aYHPdhex2Ple5Woer/6YqRIVQe4j4PE7MzdW0EYdwBT2zfQC0gn
Yc3ziGMcqM2kzaj+u82l+zsFod32oUUYMrltfq6xnkllY6znzqLXbDzkgZwcRgRh
TCxcO2v+0BLJNGW0E0bWleRzqU8PVUnJuumzo/6VLzR86kEXBdC1C6AUTmXLSLod
x+ckLbqCnva3h+27L5rwrR813EByYeneCo8qekEKsofNsNZO/AFzefrVw33lxKDW
hBITIgXtP4T1D73MquiTGDbxYwkLDZ3o3msjVSduDz6kDTa3Lx/6F0AJJJxae8Ld
jNSY30gRXPkB3CEL9dkGl1WO/G6WAzHfWxauKNeYfUL7n6QFrrsW4S9X7plhBxSO
RPfSHJaBcYKAHlWXevmremVxXw3j7kDYqveW9zDj8ns30Ct8abOacsyl3hX6lKB1
kN0Fd2zDJGZXwogO3h2GrpgalgJ3szEt4wL+f61NCmsUtzpDkmQKZ67xBzc6iBQN
RPsZ2FLa1HrmMugabzSj6OTpBLqG/sB98M2xw+g8ZoQfxQFGbDHp6SQ7AKfnHVUR
MfkXfrbWp3CxU9IbGME3zWDcv+DOth0G5g/b0fXdjxBTA+822LhhvK44i3spzg5R
Y7tRtGNurS8AKP8HY9xAacO61IFDo6Hu3NWbby//6z3zHH9JV6sa4eSlMhBZ3HWI
Q1mj5Cp/hNXMTs++/56RiogV3f9e/Jnrpwb/hULzQCDhAtqm3C6/pus0jHrsQfBo
nIoQ6jp75/2eHvglOUAIa46Rk24O2MLcJj+HGIAzOVUr3to/LEUusXq2UMSbHh+E
HNWF6zfE7Hy1UHjj8aiKGeQrRBROS+ojdExR1O5S91/FRAv2Ga5awyfZaNOGODX7
wdAZgo8ZQisy8Hz0IN7GaTYR2Hub3z4Kxukkn6Ohtp3qnaNqRpWs+8zS20aT7QZO
SolP+J6YDKZkA8rBg8AnZgnqTz+9Ks7sLPgzp/W0sdte5GOuAaVf4uKr9jWjFins
xzCQrql6SQ0OjY+vWj0CDxvM1jF0m6Zpq+JTEzb4PYFVHh4KliaXkcUw5PtsSVmF
CKMZvXQsPHMSB2/nRHG8rCzbfJBQAz4hj4U5usPRNwhIrww4AWufx9tB3XQs4WvI
Ni0/2n0Zn1HoFPSCN7ojcJqPJ09Zr5t1FwPiWQXD5OffoMeWhUy/Y2EW1cI14iVu
eFaZ1wRv7DxvemhwqL1O29WaduUbFfsip7sYvix8Jgw/Z3gdPbYuIg69gy/2TVwq
KJwOIYrCV1zE7pMDhXk//3EI3Ul+zPbAGJRhGJ1BnHjTZ7Y8OH/hRAI2oQhKvlJ+
h8x0MUCQjuG9XpsF1YcjI6Rmpy5E/51mUUE8LOnC1eajF5hVyLkfZ5crztbXtRIB
CxmB9Aw+r0vXkt3UFpPz03f7YL9cfFaX0PAG8OH3yOIyubV1Qf22GcCAGW2nAvse
reWJXcUMkVmQmahA3o32iQrI6CQDHjsLfleYilVvx/CZ83XVTtfoPgZU4DZoQQNJ
+4MUkzPwFL42vABre+Af2ozjTlP4bjhJLT6PwFldvotwrWiUUJLir/QAuVdY/8J5
hhGDxGYUAeuOgPPcdpJ7IsqobQAgLSDiO6VlUrRi7Emy/2wfZN+J3zeefjVRtdHd
EvyTwge58y865ahkmSitur+CozxAYjHASK03rztnd/xntTEyqZ1xzN+9gZTzayT8
La7LFu/zSfN6rVKuckQCpLgI6lJ7URjPnsIdQeQvfjXm46ozAdTHB82TwOeehcqI
8x+wvlbKqpk33EgErKP1kNqEP/QzwLhuCWgkS3aUvTIH0FMASvhitumVN3XM5BaL
0DcIOHmaWIp6v/t0AG2uDD0zeluXx05DdzuGeDzP0R63x45GRZ2ruwes9VEC6hvj
f6MIfpY61j9jFWM/YjLcT7plIJF8P2tjUAHe9bH1FK1QzojoIHUTLjRrDtZ9pAru
YpXl7KLhVoU3nSWCPC6NjziOfAHNXLYA/Nr9KLH/ZJf9Eo4kdEHlb54L1UsjIvQ2
tr+gEdthzhi04P8phDB5WA4GoX+C5bey8njlDG4rFTe6B2cdpNB8gfhrnUB1VkOC
S8Rf9gXjtEjLmKsUk+kIrQctYWbMke5FZtAPNiqS0Uc5Ng6lLncoe1oo49UfO6bP
0UUBonV0UHxEiZHh6/tOl2hlncc5PN/BoQKTYvmD/ZbUVnSnNT5y5bvq7gVe8W75
7dP+qOnXYFa4m1+g4jS58p4/X4DaQhlHqaNN1d65T2oRySNRjHqqhAI+5yajOPxG
hjdyAtoOO4snuamL6OJJClB8YU83K0gg9m6viOvuR/0lAZjlDPLJx7fG0fvYGHjG
STrrw3nnAlvK584clj57+orilLjJBEjqQdg1BHmUoWoOfmxu8Iv9VuzZL4hwdzcV
Nww0h2iB4DvG1c9o5V8W8w9g2IagH3ij3e8MHkpVCE6CgO8rLC9J7wYYgwJa935L
/gPQLC2mlSEqDrtj65l+nDVsjnNTeLnxNABGlNtYXgeO4WqWn0cbF7+e379UZhRd
IgSo/XkKXDVBJAJwDcE+S3P2Lx77QInlsKlIcBv7V6GL7agxfmCyw7Rrv32zqRrd
BG5VENU9Aol/23gRZeDSTxISnbghLPZB2xH/NVl0O/WhNQWp1RtQRgyKgqSnNi5V
qCbGTxmMRXaB2tZ8QFMQVoq2BJu15b2q7QvitLZBGLGtB5DTIdj2a/NNOli+QSeP
xImzRTOWZ6tZwZs8vYqP+FaSIc5I4NGCuirJ2EEuvAlpfUdL9odXlRCXNP45wGY3
4K6VIfOQmzP/EGgGQaUezedDMkXPS5V216a8JG8WKBPqZjzQ9S8EgBV2PrOdPohE
j/rZ+wZ5qLYVSRuJ2sT1YNQ+NvPGQoiZSfGSWfosdbld9akJrqx/s6ORXhMmn0dm
XuzJW1992nRW578ZeosB77SVN/AQ3nYxVUwboKBo00XSC3Zo2bvOQT/TljR5bR84
ePGpGoGMO7vy+r0rvBagkfdKnEesT8HOatz1AS8NYqzPzn2BtLKdQ7/6+Uyn+OaK
89D7crlKpwQ4inb9NNs2GF0PZWrh6qFFxlvsyLF03KY1vP+eA0Jow8VSwPaWQbrN
dAxjo6aLeiEnIYwF030QhGIWHBMaRv4z8WPTl2K58R/95wkty+iF9gyMRZOm1de7
rSCwRSUGzGbajicwn+l8N3ZYYSd77qaftwOj+YjZSuvhP7OeJmWcNCVGUjXjGxr0
RxXiDz0hh6SKjNooEze8/PWIuYZ6N1ZlUQ2xGZWsFHTCKW6nLk7o8le6Iclz4K8H
eIJCy2HW/vjeYznKEQncv7OdlWvq6EHe3lHW3fqOfuwf664XNawvF00O1slf3I7h
dfhSYeGH0uDULIGH5vtLFa/FOMTPe6BZdpswlL+xB4J7Xb8SNYJqG5KuzioSLdCl
IuU+z97/XfDknRZwW0MuHU7rjXn8IN4HUdQEN3zaJ0axfRgbKE+SIDniZETw5emk
WUnt/DGaaR6NeaYGIE3FmqQixPT8NiZOdBmjJK8tDNHwaE4PTysFt5UNJWxWB4fz
OUd3oLbVTDcSXEpE13SD6z05f3D8JA+s7QKPUrVzIYY54iVNoJS/0Z2N6lFR+ayl
72ApBMSogykfeRP0PaWcBB2aVMr0H4qd+ApITFf8eIFcMZTiSXj6W0qhaOpL9kN0
gF+RQa8aLOTFviyneK0olhma8l7TfeKPB4pqCO4XE7tEwRiPj0gbZdMCcEx+BQFO
eNQppzVIkpdYXLc3B7WLpakBxM9SNcndRnWGSzu+ifa5KH1L9J4qb4I/wY0/Br1y
tCKdDqAr+6i2mY/g/Awib+xqNyNaeA1rXpDYO4SYr4VpYLGJoBCJRrIQ3h4LvHKt
EeRztvqBUDmfW2OOqvgl/577GPaa9pTYdME09jhfn7eksP18prB4k1pfZ9q5fHZQ
6hhzMxXlRKFDqeP5vhFmuLtiazYnjZvoXhsIq/JDdUCWftC51FoG3WsO0mOF4den
9BofBCihgDBx6ChZPyCgqqCnUR9H13qqfHHAiElxYsvhEnUGGfTHrWPYGEBp/e1f
L6uAFyJDGMh6rCWD8Yl2fp/jy1CmwClq4Kk48ZnmO0zLHDN2qMkhzYsaVg/Vig/+
N1/oBKdJuMatX5O3xdTL3I757D1qubsf5tAcPqSgRgqB7xeMy1VkO5OXkPPINQQI
oAEV/lzMQ7jBBIks54UVarwnLFmlqqdBEtlwYkUAoXRskNLbicPRBouAi/YxS3i4
CQspa5EeZgeSgd6MDDZVWYn6SxlExcA4lchn2xGFQqyheRMoIpfJMKdh67g9OfYn
poucIjCDOVX5kOQtGX+TyNMcWi67HjE9/b6dhsVdT/CHkIkZF9HIKCz/ieEnycPf
gqg8jXVePhZr1m27i876svxLgHW4pj+Die/Za+w55fm5J8DLAhtSVj87Dxl2Gt0u
GEuQdjRGr4NeEuYEqhRSU1HDzoj+oc5aRNmjBZkknFKA47LbYztQ7QZ/yQlqdAiZ
N/cEG3lIaV+7cU+miMZsMyOloF0prwUkzGAa6GCt6Tgoyq5NHMicNWZ9Bl+ydd80
MEC8FFpc4XwQxn4IGt0puYTdpaViTmk/xWxQ0c6Epux9XnjHdesO4VJHLHQ6mO78
Q7TH5qxghVtawATIpJOFzFlUAyKMH0Ng5fQPTxEmQoKWhy6HdOZflEo6WQ6gxnCl
OZY3//qCj6jqRa0BCj2axe7P8GnBa31MtySEiopq/7o+KpdpOcS2Apra4sGcExCe
+IaIkdtdQJ5TzlvMKQQ6tZSoQbdUHLkXxbDmGoCxCrwoBpOjH+TBNccS6rUBmBVl
MX5dW7UjlEOtL0XZVqwV1LN1nE+5Z7giOUC3Tzi3IGPfOCLQhl+AJ1Xb5jOohxbi
eCEtrxGJRMr5tDYTlLVk2QnXsp1B+kyD/kXMldVuoKqccjL5h3z/QFfcPPonwSkj
IU19mcnEs5TaQYENcBINnWx56AHHTGqOKm2dIp8FeevutTGRIQNnUQlX9iwVgFqA
A2PW0lb1TnqM8WEgtHQIo1wLposE7bCSS0w9r9vWgBj9Td1eyV8Saj+j9XegP726
10piPaZYeWozbP+CXCEWyvvWwP370Vzu5iSmNk2qNaIGybASy2qcDD4bFXl2PHWd
a6awpRYFrXvKUqjaa9Vc8XFZYCV25nLDDG2Fkl4uxMbv59ecJLD0TXZstDWvl/Zj
Pg/Q0EsfYOOzfiVq8qdEs7J2C+7l/F1axp09YFLykiuHy2FCIAytZqrC/4Suldbi
YNr2cwff2aAy1t390H3ybsxzrVyEguELu6vQ0OHyKuf0LwzkKQmXPuFJ5YbYtYba
ZGVc2mhQzLNvb0WNHAa0ep2Vq3ktMndILZxOaibiSTVNm0/11WFvwfHJL+ZclG7C
o2gF1wW41+ak8prmm9TNChF3DZUfeSL2dx6WPVRFq7NdbSodYM2b7f5BzQvpDEaG
jaEkkUnyhRgjp99eG2Rqu1yIWO2UhbPRsLrn/GJpEUKr1Xl1M3HfWDIti2zD/Tcg
PjGyoP2EfIYEQN5IV+C19UJ1BVpGhYWPntkdo2+G2rdHWI4kERvCFyMBw/CKSk/i
e6C0qRhU36qz5bN1/K0kOZkPWos6JzK0x5kohSKPiWx8fClmlijp8t23OAz46sXN
DwMTLyb8dH9U0qmfCLEu//RJC5PW0hCBAoq/N7MJ4O3mvl2IE0o8qId7d9iLldTk
HVoVtumhG/irVj0sG8TiE/RCRD9K3q5lQyulSjE6Ypdrmrf6g+NVKiHCnBfM/6uX
p+1Hhn/krX8XRZ+YT5jjxUvx0UQ66NfTSWKdwK2131QFH6/0CRTC3yyugc9VJWn0
GpS7Wl0RiV8GEE6LXCPiwVc5vKvsCMMIopRMD7sEHzBLcuyzeEh9TNPy8orY2tt5
hGrt1vQRG4Kmtft/X4hOvwmafUj9WNp7X5cqWdK4xl4J1cvLkyRC5fYIr9kCWKQX
cusZDql+X/21AwIwXpbF++2j2WPFz3JLThunWk/7raFpbwzvzdlQtkbyjfX/UPkX
UbnLNyaLchT0F1EcImQ02VNvrpTXGV4/S3QfiB/R4FhQiGaO1lM+Vp553e232pEb
bQIxsCUn77vH2hJnZa5NBaIa/ndDTeyRK/K78DgfEHd4b118h9I/VDiLdArtDrTc
uJQ7xyHY/+EgfVY1fplTvfkb+segJf9gg6aZ+wrIvrcs3Lut43pRUIbklIttbgoy
nQBy/GWzeChOsZiAVvAYE5DEfBAHXlYMMbTu8chIacaw1mXIxycAX5Z1ejxlJnB3
NiNyj27dCCO9b25x8N5IGqVCpg9mwzqRKmsGZ0KO2KJiViE2mdqbItxFdG7HeQZX
qTlz0i/ZyPlYphi9VHruTjgaChHZTkU0UHoQaR+e4yG0x422m125Xl8BB9htaKhF
mcGo1XlNHBbmFrTo8oL91nYICcr34CCI9s1D4afDhtfmUkJdf5lUB/lfAKz27xqT
SYawuEku5CmE9DYwFi0LINqqFYo0IOn1mQ6w1fzxOdvAD6Ct0KY9mc70tLJzjZwi
iQ3ZGKQg1k0oVuyQDnjKYqOgyZN9UwvPH/liCNs3jvzKQho2wNQTOUGeVVvkHjQV
lp63AdJ+tpDqzAEDNplSppQ/+dIVXK/wlcgHc3nOW+mi1ZBPddtPdKtXPXQQB3RA
volpNDMlVk8irOtLYW1ZXhoHpJe29q/Iz2XK9e+U8S7GzKIjuZB2sSGUbfcN9ehw
A1rW+KUACs1ckF+O9T6CRR9YjeMpxQ1QCXGmDHMBsl18i+17T97aHeUvO7CNvLVU
q1FGkCJRJzP0wsnLsPB1OyogKlLZu4H+y/XoSJHw3hrOA+u2Q/Yy2+v/Ez4I+6Vm
H6VdTAa4n7Nj870tXRcHchAMjopDBHdBuZDGAgiIf1IsSg5Tp2RkOzW6bCqz3ONc
BtF2upGsUkyecsXz0dErrJtNBZ9DWheV2RArq8JzJfEzlpRzhteurYrqm4hQucyL
0bDzkbOCl4If+2Op9bGSli8tZYFHuxGLUb72O3bdVGxR56TtEfv8Y9gs22gVybLl
gg95i2F5kUv1QjBmAy1IstKmKLD2hYCnrk6Ykk4d7dkZdBk8pRmHu1z6AnnWrgpz
ORF3UmmoNgAB4s4KN+nbp8/Ve8JnZompldSfrxyYRj/xJkpoWZ1bMfCAUCPtxa07
LORxOpCaoxWSNrrsrp4YYAoK+W9Kg2v/utx2oftQ/vccbFXiT1XNyaT3pRG3fqaK
rlVgmGa1MC8/+8o7OB+zu+eZ1k0+i12gpexWGHiHl8XGAZUYvkXmr3h8qgti4hLJ
H86MfCYRtEzunkD0RMaLd0YQYQyw9+J6WdC/ZiB8AV6CNjjINV8HZ0VgX1eYajcj
hiXu51aa3CFSsN7VE7gZ3V/8eNSPK6NU1wEdDgpo4puIDQPcKnoVbdPWWiCsV7r4
zE3HLYtMFqY+d8rfD7sV5BOq/GLqzl7XCCKngQLa+CxMzAx3qnjAvAkZJBcjxjXC
sssfF99QCqcgTK37C+QzT+UQupl/mTi8YTpumlIEez508u3ejjlRlz1Apdx+Ivaw
HRp7Nbne0TqL9nweHaC/QCNhD7bRqPvDjt+g3qDazCpLoIqNeK+figgjTEfO4X69
X9bmFiKZAy1f8H6pUF9qhZYgaHWdMCWWpeZf/ipyBA0AQPvRp1YOZXy4raOV3+TI
u8fX4Qmg4ikLtd43uvFiC3TTmHzqp+FOuVjuVEYbK8QeaImWTJeiTarHtQCPP7FQ
estaJhUbg3Xfb7pc6t4tqncwJzHm8Wpqliu8Km8u/TIGtNqXvzPyBjooMzP5xKHR
U0EhM03pAsVaURxYtArVbl8IjDhvcda5AyoaWoY0yaY7keqqphbA2GeNe6qXvxWx
rfmoWBZsiQrtSWiHdUwZb5paYEXt0rwxm0PhBAhdaWL8MRiKKPEHmgItdH8Zw/UA
YxxLPQJFJ/6AX3QeUP4my+WH9zYdDdTQIGCqMd3TR07KKFeIh5+Hpp4NDtSLflVg
s+8AUPVwN/78E5feWOoZqvzs4WAyiDwHWLDiinrMfyvivww46QYmNwQxX+suZ/Xa
NVpGYV6FdXVo2VxhNivVXnYXSYpl5dyp7dFXvaPluFBQEI11ArxufF09bem5Ylbl
kUU5LEj8wcxRB8UbfJb50dJOSkIw7UAxucThUEaSrYwBcMWRpHTlEwnM9fRa3Y89
JMNLsAv7x8qRLZjirUar8vwq7eV8YRE8B6uVNhAvDwo4tB5YYpy55RzOx60EHD2I
Y0rwgUZDOuYGwR2C+UWevpgRL5Ya15jQgdSnlZysY3sUjZV6+vr61f9PaiN8CxQ+
sbCPMBBIqblPTcbi787Ww1FJApd4doI+ozdCI+dTCr4dWEDbs6M4r9OoxRczq/6r
hpfiwTdmmMLh3KowTKxk5R95TrP1GHxr4oTkP/7FYytKqJWE49FLJSB28G9sRvDq
13xagwwC7TAiBE3tSao51wjMkViF/+3c80WJl/bnwS4J07hkshDviv7fTePtcAH7
NwyJ52wJVlsa2LLdIRxWaDGJ6pOFQuQwJZp3QTEEAbpOrnIjtioY31SShvwTHQ1s
xerzSf4PHKUzcBtiJzwWRQw4idlmhmLM9bKyJ0sbesUJngXix2p+AQNtgQ+upfep
yzzNSgbY429WmG2zXNALQCwAkwop46NOFjAcX8xCccOIbkMDEnSQkU+zTU+RvV0I
jDY6g25qOOxshgoK2Pr8ebJ/ViGUk4ElsE1ZncPAs2DEZR5fiQaUsn+1iGnPgd7I
L0ONh1ceRSbDYGOv38q4xUY2me0VOCE6uVMpV+aKBWS6Lm5I7KHuiYXZXSOuBaHa
I9QWwKKe0K9436TD3oqWAlh/JMpYmLPKPKh17wwC5skGh/8Gw9PasYGICapQR7Ca
43K5r2qtJDc4LmxVtkzWzpcOqoOJn3xMjGo9CSqpJ2irfEmMwpqgfoXTBpudVynP
ZvReDlQc9juAIxbaeKUxKuMDGz5rkoAtkTdpdNScNCg2wz6OwB5kdkM0aSaKt5JL
MZH0akigPbv+o4vVve5nP/fVngP8PUm9awTQcj72g+JaqQN9Bf1BdlpNoH3d3vMo
Id/1GDJP84/jOxtwZgKQUOLtTPKPeh4k6Q0C6jEeah0gfTVxzhGNvBzYI5z1b3mc
4bMmDEVOQQaKxF6BYG0+nwfwr/b6kSkJCulJ3KEhKoEynHJvc5SbeegFpztw0BZ8
g6tG2mhqRJNzvxM5h397nejYhEeDyc+u51zhVJZEFNCENoeLYsQzhLkYKoBJe8GZ
hAe3RxUcPRTtHobweM6aTkHw64hCTCHE9mHZpNBSaIqlrHwHXJmK+jArP74aQpMk
tryf41SpeKz3NHsfp3akUC1HCzdF4NKPSjvi4B86SPJFl9Ico5e77lA46lPledCL
FZS8FnIY2PAqi7XBaG9q4/jm2Kuh5oPJw064QfzMWUKVvFwTNC5Es4JkqK66Zxud
L1rVL++oIUz/RshNAyaHqcLAd5HA4X6nu2NS7UPyw2BcFTsqlUvlj/sTc1/V0I3k
AIZ9181XgabKBlGLDJZT3owgTb/eAeSPjDyNVdfeowfabCSxZUvE+fEEPHQdBgVz
nLbnEHz8GAloUkk8DQHPuQTLjOn2nrQk5aYbKOp/vUyPdHAzh0dnq6f+aI9xoupH
vS0HF0qqa+S46SJ6poekqLPWDVwM0wHF3/XR2SwnfFQoaowv7A1O73YDLqg/HZKK
xQyyZwvaSv7PJ+QRrMsyE+kxGET55Fe2sjkdlLQg053qvQPAzXk3RSa+Wol0ZOPw
4wQCV/qMXheZnvWZrsjpPpR2sqovqqORRCQjinT50u1xPwhOb3UAK6vhtFTlLQPC
628CUQIMCLbI7sLoZexftr3bAur6QK6ymAsjfxxGSJKtpywQS+oI7ysMOrtamn6B
aHZDkHao/BjTmM+aBVv4HFOJVEarYubGSUxudaS8pMHUvJuQGg+Wv5pUv+lin+Bb
0fGoRu8PR4nzOATZ1cW6S9vWsXsB0Jv7ft6Eky7OocuRXRhNqL82xmgfuCL/vIdi
oioD3c4+xMhSybUgqr6zUolnMmKv5spApW7CcQYOdLQ802OfFKuwG9deRnvrQVnT
b4AbTNBIu5n1mw2HtSVaPlix/jy61/9FO2da5wkOHtNeZixO+5vXsgp0qO6vcGQu
Adp/8L5On6lhNysI28lYx2sJPJ+TTg70qMWUdctsz9CtQ/KpJanhDGgQ0cKPcwOt
A5daSKKNqsLHW3zWXCzKjLAbCIFz3dcLiqtYfY9yc0LenqEGEYc4Kk9ZwOZFGaTC
FbEbGD8Psa8TMQQVDI1CSRghTI//kgv95DhZzPDFSa1I+aXGkAPYpvP3jeLzPuZg
mjswrA+DZzi9CAeIkfExynCw/ZQFwJbF/4jc1sI/NzCZa86LAXPaWrPDL1Xc0o5Q
B7QWylYWZIsomgyzU8dDrB99rorTJ50r58hppa/mLbieIhrh3+adZ32Nu5/GzChZ
l2vG/OylmoxQ15r+LRhOhigDwCKQhOubvHtsIT7DWpbcwtOcD0H5itkZE8LwMB4P
ea00pEv/UoCFugXAJ0biEM87aEhghX/XfbJL6ZM0bMuP6CdHlp9AEuE6aQ6DiK4o
KeG4I9gMFigFaESiccsGizy30issXjRfRkm53ZoUh3bbrWJkI+BmE/4spr9cxkDs
zYPO9bSK3h4ogvMwdm/zlogoM2cyAUrbW41zdnXRf2w2Mu5irC8T6qrymo++W5Si
DML97/hpQfZ0G9gIxsemfGgaX/WyCNTZQRp8K+Y2o06hmm6T/x71voZVKbvZZ3QU
qR6N2/Z+9965TUzz04dB79ftJEE+Tw4PYuE9QHXc14peNYfn1StH3XilchPFcYb2
5M4F3RfVFKR2607x6kLGwLkjwxmJUFQJ+0/xvRBc7TFKksQDwuax7OcqI47yQ1h4
vsgVo4QOTd7bCBeiqOiftq7f+F4ulKH4VrIcKQN9S6HrDOP2XT8n0VD5XwxvPe7d
DPvAMW5QpP55RguLMQn00qqY/X87VFgXDC/Jbv3Te6+kFtEDevAgS6XKK1s7IWST
1+TbIAD1HoCRkrz8p2NijZnAzFXmCzIOBY3Y68KXUJEfW2cEDfsHbq2splCUQoZN
ZO5wnM2EGZok7fhSrj6w+5iMSSyHnR5Qj9OHSlJj/El+f3sQu62+X8coIoPsBz0z
zf4OdGz9gGf9hb/6meY1ylFiKfMN+V52DXy1stOSzfkEMH0Ui3Y9XU2yhxRs3/4N
hD417G5jruv57RLppr0SaIwrIhf6Xf6NmyOBtkk+3VZguXrQxdQ8SkmcECF4TKOW
pnpjhhG/krQR+QQZzgJR71EDH4E95s4HsUx4N0k5+cpAV58YGrNB41wea9QM7CGI
4yhx09LvQfmdauxPmMpT8h4B5UEzcYwGVH/TVQktY8dK+EKiJuLnFf7CmLCuUeu8
jFS9DmRYaC5MsSVi6QrqPreP9bakLuIDM36LSJnyOC8iyViKz+IqqhERW7YvqtVT
N5rjncsEwWr+bgZ6qYy1ejwYud+841WtW2aYj4Q+5oVA9whrEymGTvc0z4v7T/PA
k0NDZGK/uuWDCoV9XLy+OaOZqMz9AMRka57fFhFuTO3dgqhZw48yg+64a4MtZqgY
6/XMeagUCzATKuC9GhPSDac5R4Dq3vWWrElQyArzXyGEH+oaFB/LfqGFRd40umQc
GuVm3Gt04Tn6A255u5U5NJV1Bu5zXRoz2mL1mhwwCAmOVxW1GV0egfqLx3W2ggy6
RJNuv2ynk05rQjWZhKqLl0huzKNHwNhVgl4DAs3EjGFFyAvOVPz+UDlvCekyaefx
PT2XzaIakbFeCcGlwEf1HxPfpF65Sfiu2lqS1NOmIPtH0kr+2Zc7DbwQe8yMKNeZ
AhRYEdHkWlUbW1m15BbmEvWIXqzBMmvMOnujoyctpPF+Eg5Q1x5+UBZhYJf/OzNU
e8oqIC0OQOLPkONVJBl+2SCW0vUMBmcNxXnr7HTGDBYFpzXzOtL4BGbKRdPCvhrj
56pz2b0cys0SCxyNsrytqaKSa/ePEgMCJhoc+b6m66dvUCtvObp2BxLppymJRVRt
mhUSvoVIcDlPaXDG6xJ0nY40ziwLlXUWWlpR4cq6HxfQlUDVjmltna0lrCwtKcRR
kLQq4WRz9+xVl2JW2+7jgW6C1qlHWhXWgdPnqOSRJQyueufrVUSN8Bg5C2bCNqjn
8SkCpBc0jQC8Mki1He3MFQKbuG5HoF7ebnbwatoFEkWp+thT/wbTV2kyLfDsnIEP
pLXQQ0PYE9CD+kFczvDKhHK7AOuerWKPHAy9MXVkELIqv0GuaxMQbzl/oea4SGoe
nR82sCf24QPS8l0Ly/21ymjD871hVIbd6Wl4/fuT2Mo3efzAgPky5dF/7Q4dbOYD
0Ma1ZDP3v01QFJA0BsFetjdccO1VGmOlVUq0feVgb7vYk2nDTrT8/g00AivB8glV
jIfP+qrxPwQHZPbW31iyCFyShQ8Jl0yUWbBTGO/895a/RtFtifa2XRC5skmOdLSi
0FZgT1JvaMgA9VvyUEdRCkxM4z13/p45foDv9Go7I9/VbA2+DPdXgDQMaH6F7B6g
bALXga4F/xm0IG2lxJOSwvJXC2N6t/mRHKo0O4hTjey4K1cXlfRBUbJcBYgb20dY
/PWR7hAVgfnfk+Tqj666eEMt8bmtBy3Aubitkc6X/bCsfBDHTqS9R8J3IllWEaFW
ijkF+h+mvvOqah5Kw8DA/mcAY3cWR5rOkrHwxdpKpjJiUnGypUedrtmQUpeq1JwK
lUVRTu3vDZQOYBEr0AviK1F4PdTyUbg4fu9UT5jAPOvHPnWrtPw0DG5GlsGO5XcY
1FElUNVWEQAnD6Dida2GKENWXAd4dsB08DDJk190odxhgapGZfhYapvYyUqJc/mC
2ADSWAIgn15DdH+eXdeORQ==
`protect end_protected