`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7184 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhBNVMbsl6PTB5/ApNH6uD+ABMea5lxpzbviLFCJvUttO
BIcMUyRwD8vshJLkde6WoGDnXl5kkAUCG7eC3nYQpuAvSSF6YZVJbZwlo6POQ4I8
znPuuGUobykC872Ow+D0RwUkzABxcaNqoDSqR/tibmOHVK/zPU1T33rlZe7JqIMU
w1Uzx8I0KCFxp/pO4mKN2YPfc/Gc5SyMF6tGdKddp4D7/B0/y4WnPBHePhYM5II7
hnDSnxPPMWkQncEOByO5df/8KtjKDdeEctWo87a63OJECTd7VRn7fxV/ToU3ex+j
gbCP5Cht58Npj+aQI+yhNmTxGGYdEX6eTzepYLflHO/tGLfhCNqvCvcEdRepwnxO
gB1H1xcT7RL4/fD/IYsd2bwPdh68kq30uQgqn6WOGzrCJKWhNyv/aoIs3rRsTsTx
/Y7H+8CNjZorxqT9UdR11c3Yt4DZ1scp2keCtzMb2+avm7iUSKmWe7cxOmalDn23
rJNyBUm1L4ctPUts6ex0/RYhPW5aR/n1ZjywHAonVBmjC1QPi23XyQM2y1tSzEoV
vgnOX5pbJF2RE5MH8COjAFaGD9f5FPuJyUnxOXc9EB9RXsXjoBm4N4JP/ZkL1A5h
dsVKpL6z98sb1kPSsfLWYlMqx/Le19aOdmT8MtDRWDwkgN0tkqejM3I7Jta9NyFZ
dRXLdrNI9efV4wuJLr+cxf7lj+BvAWt4MMw1Ag1N9yP72YfWHz/4+m+EJpwH883v
Xw+ib1nN6XZlXbQh8Fxy5Qyn1/J18Gi/1MjXSqrAOgH5Ot9Tu6d6rdFUu/dPBYNi
QO3TQSIWwHYxLPCh20HccMjPnsx48STHr++NixN/D2H/cHJFr/X29vmzQxVxY074
M9VZAeT+CBuPTiVsFQRgtC39XwKeDCQjuoLp7cfAZfZS27LeJBp1oLOtaMF6h5Kc
ZGXmJtcbxFuctMvid0n3daPQCLuhX+81QvixOrkE2/3/B6kjIa3AN1vqcZD1UKH0
HqKsCc5m95TtAkdsYdMK4nhNMNx0SZgLTewjYDq0cOr8ZlrWUYpJnPrv7hJWHnT8
Tjs6rp6yhzAMXKUrlToJGfnhcHMNXBWavVgATaU2KJtdObBEbKRiiYgYN8PigeXk
rtCNpwBE6eDKaYOiGS262Bu50EFw5Gcr8nbtajZa8yu9P2NbtmhDdxfHfkCvjWNO
z1OOKKu7bUPCz2WkSbQyV7NxYp6kDAzsQ+RwkiV2CBH1MDYdnb7YEBdyEG8aHHNH
SqxRGTtLzBm7/6kATjNVHOqSmSiAt3CIQPoFeAgdvgmWkNR46MNKTd93Vfdi5yyX
4nqy5XRJol5RfcqtxTXb1JS3cGnQNFy4mbURg2iRRmK/I57CzjFKubQOlkY8rLur
UFFgq3UbZidd4duzCSO6vrF5aEhrlJdstPpqT+tK6IFHjSrn9MK21bT0N1Sx3Eum
Nk8vw7o97/ji8Inm5ZpmYIP0T2CjsfwPM8Nc52fYeDZnNN8r9mQunASRazESGs0c
j2EWw8jC6A0thkA/RHY6Rts+b4MEzTqtJ0qP2YNl1AKe4fi7RNXMK5V+5QPk9EFa
zG/1ZsoU/u8MY+svwCeZC4q9hBJ0IbpgoTUd48W4WlYy+xrSMhdGcAX7WRfg8nG4
mgG6NVUlyh/RuT3MrNegLxfB8uPS9k0UZZKvbr0QsNLX2oU3i6yYGrgiGM97ps9g
yxPbrtgJFm8kwJzNBX8tg9qfvfroM8lJdoNEcCiGF7xT5BuPnBSGXl9/0HhCmAKv
+durS9PcXQSwPpQNW+ApOSFlMWSK6o4jwOgJR+ZpH9yF6e2rVF6m94YWuzguG64f
PGAHUCkIlnPR4eB/DRuPtQdQXioBVcarTpx3JuzU+cwwMB6eiFqqIOBl6GiA4ky7
sK7hyEMp3RT96T42ZWZMFBiy4O1FAUy6UAWhZ9FRKGQUtPmtTU/3w7dOVpwKNCZU
XIklOPfiZEsr9elAq81bd243tdlAYEaTN4wprJK+vNdJK9u7l/yVxJblO1AHo7js
RHiN+W/wRUHK2fUGHg1tfG2cnwdfgCbkJ6Nxmub9Bz8e3iSbmdFcKzcovY5PLpFG
zHVrAe49BLYwZsyEJw7B7GUam6mhawuZIxJqupb8vGuMxeMN2ZrcEz3eTVa1U00j
SAGzba/6F5JlfUyyUFuLBzseuibg2c5FgQWUscmzz79m1sNyas8xpKRK+KDsah6i
NT5oACVnoLBYSX+q0LXfY6IsCCzjXBZG55kAwG3pOZPE1TxYm1SKU6EzeHrKJvHH
G0fSYK9HhWik4sxarI4GtTgZpmlYO3SHi4A1LKqdCxkfWKIShNSg9+sLNez7sBXq
Lc2/TKRJsyguPv8denetk8ELgIIGI23lNBqRRkJlvvZTa2fO1WnTap0biGmEf4p5
xDrgDrByCmuyFOUA9GEBbwYfcEZYZw4HsobUbLXX8V1w4eh2ZRvDzj0jqZFsecIe
8SWxjyRcRtZNzGV6tQww2HOmhuCw8jfnfwimgqcBdw9m6JuNslDOYhs5eHoOtyW8
gIpLKLNL7IlwztJDD29ntZW8worJnIVjCBHhQSttvyizQ72KtxuhQas0asY5suU/
tmFlm+bye3j3hSbe/y3Cfkj9piaKnzMsO+nXU6p+AljE7GIOW8YknQJ7lfd7TmZ8
uj7nBqiu+7hSbKygQzenCSGgLrYraAuDIhtBb+lA6q4Lj2e2fcLu1+KUEbmzdFx2
KpNLoFiPG2pdxdmXiWWqSRqUajDAOsIdxlSSgXFkkJRhRZ3cPWG3/1ZTygbaIYpg
uwHDl0LiSTT97YBhtwhDWqPUy08NHuskCnp/h/y0M1mn5VQ0Tf+nvNGoej5BCaaV
/kXvELBS1LHO9Cpn7L6iFTpIyCm4Qz6TmLMUhIGSnEW8GQlGr1Ab5R9Ie6UGxUeA
KcK+BLb5PQqkeKnAx6KP02oaREz21CFJcA1tsrtTvuA2hwAN95MYW58nw0xSpm3L
jsuDN8XPCBQMtJ3DeSPt8mml6o8GvjOQvTvPEyhRDalf+ctPw8EfPOnPbpoTvzZJ
LEHJ7leZc/LabyJL+MterXQAtlNE4aRlhglEDhPwbOrkTr7aodrvHo9Dz00wPx5E
RGhRqmXyW9EtZfJVYnZySEOFOb686ln09lHCTUzyDJrIPdC0WLVykj4tdDw+tBwB
Jm3h0x1QjxJJb6NoC6aF9LZhYy/ULd0iAIiusvpNIVLlH9w+tQnmlJfg32NlcSVQ
SuEgSV90/YZX3sh3eD6elKCWPmrsYd+S/KSrwZhc2nn6PwZ8Pw3f4f4ytBC2e64W
1nvq0LoGzMgmUlrGPc9+pNzUIchT8jfPJh7ut1o2+ktfP6QF4sYyAfRr1d3so5EB
b0tMJYXwsOm4jpaS8MENXc6Qyscha7ftqYE6bNHXHic3UIAiXZ3Qj7EdJWfX1Tgx
TN57PpN7x0oHqZVHtWNqT0VU0M1+SMBVEIxGPi48JWAAXgjqc7NGmdPPirGS5bYC
6a3RI9lahFHhC2PTTmtnjMPA044hmY/VMdeRQyVYHy1caWK1fK3rY3zlw5OHvqs0
o7TkaX4tuY1+c5Q/xqpD+oETvAqFtH6PcT1cTy50tQEaA3Ag6FV0qzcnP7L9o3x2
AsRJ5i0ExIRvyyMacsS1+psVdGt9DMx6EIxH/Xbkoq4lUVWvXjK5cxImOEcJa89H
tSbngt+HnmpS7ZmjUJWTn9tKWZPkD6gdeYh2gvENHMNNmK/DJvvCfFij2vSKVhIE
VXAFO77jN/OCvsnzkk0Xu1a/kOgTwk5u5v9dzcIDhoIqeo2sQ5AS5Kx7QGaVRAu+
6SUJ2zMtKhLiH1iXKuwe8r6LPfHe4W0U9QPoiT5v2rFTwvT3k3QdLXYuutIf1RuH
xemS5bKM67kY8LWlnlpk1lz9TTp5w9uhfNYI1L97+PDwSLxOxohF2DHBG1kZrVJX
ukSx4N/STix3gujv85gLnVdCF1du7F2Tsq6rhWOEpKW4j3uyx0quIbBeyZ4BUIQo
0CQif4mqEup8Q6WNW2eEQGzAc2AypKa1N2d8HeqNDd09IuaNcrhXY6W3IKOi+13z
PWYEBRldZQP/5bqflirDjasbeRXswPx0avRc7lfNWaLKV2EVALL7ZKNptAj66Osn
waM4HNrEKoFtIRjnSC95fJ/I4m0tLdLq5C0yhA6dZ2BEbWvRRCZJWgj4b9FGE/sS
R33zyLh1v36f0u+39xMCm8WUxVymvOxIMIhE+DSDgSLhmF0lVD7AfF+qyrQnEiQL
1utcRQ1ZN2P5P9R1pWeFHRxZMo2ERV/4ruhz3zKq2mIqc3KHmhhVv8/g7a8w5uuX
TDXFtesNyGqpayQnIGfTJjbotd4jwYb9T1+WYP/n/dq9hbUBOFToTjl0hy0oASfg
mPh+Qd2OsYLijiR4L8Cq3sRDakoChKZsd8wSApnXIKcCONxgASpQ+GRHbnQ61uwr
qyYNdcDC55wzeMrLB/L6i6Uw6l1lNHdGh0N4tKphoM6uJxUyWyUUlAzgZ78wuDh3
RpCsgQsT/CVsXo0oRFP0MaLf5ApjJ1lU+6McUqdVKWnz/0xvQ4n+mhI3/2xAE0I3
lHrqmtYifOrOkK6SX/Sc+kEyKyNjdoSu/4ZMoN0YbSXe9iUi1yKcMwuJ9YvpDoAN
rVgUuIjPnmYjBYcuoz0z4t5NgH+oi5OI+oIzpN3qi/9/Xk/NBI4YnXTliZ/t76J0
nVtiXOWjh9ECHV6c67Lg24mqO9DQ1Bnn1lpNe3GyVwBko176uicz0n88dTJic9ni
vQixSs3wtdyEqRZHjD2X/0h0WKw1IKdNvM0yUqNWRw5mn8pXKkkluro9vY+2L1Of
3l2Nx1sFU71pCch/9gx8VUa1BfHt/66f0K00X6YDhUk9lRVXZgWl5eI699S66fcr
iqPz3N+9Y76FIapIhHmUxZe2w+XMHBnjSAFhvFjeL5JC+7WtmeVXkmXvanvYVLcR
mhzm04/S+x7a9FY9APkS3NUVLAkL85KtzDXBiHwDQDyvleoYXZ1n+LETXnKK7SU8
pGWQ0YFEwRMvcFH3jfbvVUzcaUQs9ZJOsNj4WJJSQp78ooHy+7ekC5QgY6AgHrXC
F49xyucItSMCuUCevYppy01T96d6X4AsmPTrAQjBx3bQUlUFwMHE0WMPpdZpbLmj
+enCfSgPpVQP1bq55MfeQ+XrRcSgZkvDq4MQLIv5/6rpsRmkJyPpc863tj95I1Oo
Sj6Jftwy6zrtSQZE3U/0m5WAV/TwYfvcp5z7qxIGuaC1zhDwmJQWeKL9s02V0aBv
VylabtTW77uYCGGNl/quePqwb5e1MFf/IVh9/iUuV7hwC1I1dFprOOHWs+Sjot1/
dDAKBu9AqvDyzlqK/yPWcItGIWQx2lauwfWVQW8F2fKmTUW5gP1GNJX7Ek0yJ/CN
ehr+K4i+QZ98iPmCjW4mlJEEMEI7eBLurONYIeIU49PP1bzI/P5Dy5XPWWlC10Hk
hwiuXXSan57PthIcmpXvFimQ3ouWAR5DLtC/hXTADq9ikWhNKidNXOOJ9A6ZNn9C
8gkb4mxLxRNHSsKPnnZCO8lXgIFG2f27P+MMq2XjTeBf5gY7NXSeb4+ApeWNV76M
xnjPJD8aXytyY/qwEkUirjV7LjJAbzNszqcqBGzYGvqRLLlBJj1gcm8IR948bsZs
TpIyTTTaTPoy8Ljt0SXmiVTkxBzlBSMMle8PpVkIDwU0dpi0BGwNqZ7zteb3+PpN
rQ603EtRLG+x7Fq0wH4MAtYZxaUPOPcEN1QF9UMOAcRq0kFIPrwwBqabdE93Daud
2Tao1O6ImdxqNpNcBqqp+bW+0Qj6lxMGhn0ka6lRKBFI+C+pickJzS3NF6x0Odlp
udbHOVzV+DCaj24wN/7WJU9iNxbQtf7JHr39SdeSgo3szyMiS2tGt9m327vOwCEv
Owx3qOzTWIDVDfTG+kLFrJKba7LU7WbUTUmDy08+CD61y3YcitBwcrwZKEiY31RW
UsMTMvMS5k9AaFERx/PSAempfu8iIPJk/UXv8Wstt88oWdU3QNPWWb8nBZ3WGxUS
Nn8rBgbV9pGFivdWPg58AbW4Qd+cEkI/n6cFfJX58qXiSxL5qsVfKpOwMLyE01Wq
CRTG7aSQLQ/yHZ3Hh8oA8w1/DVa1xNGfqYrWNn4qYbwcin8ZBXmIiEYkCc6hcxAO
6+7U/0E/9w33XaSS+EpKFTAGVjYS483gGAMU/sX/ijT8WcoEcM++lCiHDL+gCYQp
nXYIO8LO38h/nSxTkLOBZh/gQxBoAgu/yq5z60T0RFgGa4UH7S/2/tGmx0/W4XIh
dXkpt5qi3Gjb76qX77OzF+zmQjhpqAB41hOC8W0aAwS6t0oSpybd6T/uxVE0wFIz
MO41fiVn3cHyAdv4SBhxQJN2RBbvGUK5/fiVKLSRTXDgSn0fZVotofu3ONSdKMrB
ErBFc3AFYQFZuyN7qyYMnfHRnB7VjT8QkjWIN8JcXGN20AB2Lix562vS9CtQJKMA
4ilSQXaHPaZK4zh83Y0b1eVdloDbaDDLSFjGWgb8mSg3Pxlw0Pr5Ydp6qRSZJZt7
xK05I8Ha9Cko60uH6FgJiBhX7ykRsknVKxZJ/HSK/V6mDRHGi031JwPUCJ1Oex6e
1Qx7qCveKTT4NNL3s021xCsY0rb21M1I8u+sdPlWWGVyz/GOQZQJNlXFto5xh15Y
eG6rNPWo/fF7hksIlA3xQdCZJzxThoOfeIoxWMmOBfdOI4n8MQU1oAZdQzV5Oql/
gg4/WPCMP2eI7UmZfzXfX1jgIgilDzGBxQOTDHx9PFFGxYA+iSXmeBgWw4JOW9Ik
yLHRXw3AGaM3YdFV5Wyh6PM1mGIKCCmcCZaVay1KmoWZILAyxhGf88BEEx990y2T
dRRahu4aUSQzOf8QBcs8Tzt9iVonAI2SZycXbqdUY+S5zofskaWMBOOvcl3MxkVk
sAj6eLmlIK+LYNTguLuIyFBWjz8LGYC8g9MDLonK4yZ46PATlaSNVxwT2YcUBpd8
/xflTTZs/xUOf5UvCA+IHaDSaE04TLD8WVRqpbac50D1FAOS6X/IjY96P+Dsky9S
95xUNtzst79utmjmu0S7wqM8R1Ay12zg2ZGpZfNYkwR+AVFS6AZ0Xm5AEyG8a8UH
XCpw5B7vp1FNKDsr/stz+7CHawqs/FkwUWeUt5FSLkbu6nx14GnYw8K8sZBteTVa
jlbzG/V8rkY6yWTs0q7gzgWKFPH1Qu5Ospm1NcZH4rAqZusaZt2ruWiFvTolHW67
10gRICCi8vCPlZmexZtouYghxZaA/NUhULlOlpYVqqQf+4HC48PDfrRixP/wCRh9
ReWY5TWBJQSlyHcICGItGxHpJjV5stdJRH6E6udJxlf79VpNJS6haKZ5NgnkqdNt
Fz/j4fFXOv5RbjfzVcaFFezp2zdHLuajbqHdMr2NM/+ZAkoQ6QFYk3qzhCMdLiZd
s+h4Nei9Na9sDV4KQ/0R93DhjLkezF6D726JREqDVAAxYAcyZiWLejMhr3s9Q9+U
zRvcfE9+NJl492TKLsienf5mFBod/m7JUfDjpI2Un4ckzsmRbfbb0eJhOgti8tLQ
TL7SlsAhOBa5qG4UN7Gc6DJgzIAhNf8WGmPFs0DQdYluM0eU5/k47XDBivDlgA+a
SFd++W/jcJa9q7l+Ht42iGJKpBwj3SIWrbvokg1KLniKI5klWkkErbwNUjKjKbJL
h6eb87dQpRQDmdBe7lLLsW62Qmz8w+YNK3ie+6wyJxRQ4jjtl2ixunR1Reamux8C
s2wfsHvp/br538OG+G10cJLzANNlkmTZh+HB0W8tbzW7XphhYtcfsL1W1Xwj6rKP
49mAxvAvCjx7zecGtt5lOexc3jf7gl42ctXtYB95X6IkpP41kAObJ1fB/uIfjhiO
OnBH/LFUNKiVcTPLAvAewMt1IeU2cZ/shrL2qrFSunhQFfrMc4SxRg+ss1Fj39vE
m1FF001cNa9VhVqNzu+rMPRJ1Aig+WfvL7et26CVrUPcYFNYQ6eOAkDcuCMgrDUa
lQ6CUq7k8UJiC/yI71osqMX9g/r9kRU9ma8BnKfpUUzu2xTppiKkHmOyU6f2rHht
e54pVt7PCc0Nw4XBX7dcf9rDggL97ayiV4d7d4RZRHt4BsFHLIV9RNYeNjdGDimQ
TIuJNkGbia6vX1O0c2fsfHT71rvnEQ2TBX71gsoAsKHrtRjv6sQGGnqgz0tGerhT
rXTIkLNkYX3i0GfVuvPKLHAzSv5IQlxX3pCwuvFqne+I9Y1gRU8VivFbZhS4w+pI
Vyonu7aVKw+bfPcE9tkAKGsJD6LoW5a5LWt2NQ1+Gsf1HEdqNTysuAicW8Su26lt
vbQKVipfBE3jYVRz3fxnqO3eLeM4jmBZEwQLc1QmJN6ny3ZlMSHDUjIlmZJ1qIuk
sFV4KwmLyONRZ+vCeBCboYBjfowK7IqcJE38MG9phi+oFaHCwe3x14kWVauSobDA
jRLlJ6CsPJA+V2OwIQV1mQ+A+g7q4JejHUnwc+o9x+8Mamuqa/2ufmx50UbSJTA6
qZ/2ZvHBOB6HdQw6qNWKKDpbQa5REBRCdaTZ+k7sfcptQoFRe1IrcklKWIgHzn3U
2BPXE7WZzlV2APiKu6+9P50wVsc0jFjXyXu8ONuc79uq7USmfP9/PbBUE2pDxSup
Nh5fspuVur3cR9x6OFiltqxf56qYlLF9+eXjDaAMxBaYYOBXRhSSfkzrqaYJ0iKu
5BEngyjPtkGJQEtL2eryKIjxhPL7suI6Au2ZwDEWEv0jLGmTdjnu59iRNNZEfrKA
sYffYeAmOt3MHczVltUQMEXwC6bxxXju+dD87x+DY1MGN4TvujLXRfCAVEnw8Py8
/AtQIXUtoSC3JQOJAT4IKUU7Z5jx66ZUlXJmOBrSO3Ci44utfDQBZUtmr1x+4ZPK
Fvj99rwMP6dVT/P+5jVX4mRSmr7JQ3I52daEPsbNgbaWtiefQMetTkuN8HuAftEg
OQgHSg9uOSwCKjXOlhljjyItRUXn4VHSJKqdZT1AO1FcefIjy8sUxOs/7HZrTPZB
m0K7DPWio+lYl5a21sprLpaKlNEvn7/CD1FGANRvvFtffD+4jjxcagYOgdWCvqqV
EoqNMonN9SDeUk6WsWSS+bHnr+Y+fdLBgS1mA8oBm8Dp/draAaH61NIBHeC4tRAu
OBr9X4dVypYGc+HoWZ3Vo1KbxiOKgRFm2nGP0Iu4TbnDhMo9vtjw0R0BhE/dMQ+k
X+5qLsMDpaYwiI3buhrqU6w16C29lk+1LLVELApTbSKsJhDSQu560jkRsrhd9Amp
zw204bdcC3YzaViaCyk5+FAHkyFYl630oEKJ9vIbFLZSan1bS1QwGKbNwhZcZgHS
G0TJJ4f2K2T4KJx63B9Qtqosg8fWBQBdOrQX7YaY4Uk=
`protect end_protected