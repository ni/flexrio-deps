`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6912 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
xKvnjJmWFP/6yhXUuLZs6cyFXOkiDpgEOoNw6yCs0aVlhEGLCz8JaMd4MgMa9Wnv
khp70gFAgTImUvdvod2D6yTOSDOMS9KpnUgTxP4yTB4w0sWA7aTiY1zETroMW8n+
wXr9Su4/dcymNlL8n2gq1W8+SR5QoOZNY4lZmTDJOU8DK1j5DcWEXcLO5uQ3md24
pb29vAvw7UyN0leoq7oOmbkUlJAsbw8KD3rMCrAIcC/0xMM7hdvj2NfEwHZug9Uu
7lw0kbEdLsO+q90uxYoSC8VOmkan6BFfdeWEcvbtSloNyoABy1kx2RJNQUXuzdPF
oEjlzjlMG21uQKqHivSEbd8AyHrsgP/FnEKmQAxkJfeMBHvuzbMXzVYL77pT15VL
CkoD3zxrFdB5NtkiC5S2/yknIM5FEAA6UYQC/bY1LXqQNIjaiWHgln1sT3tnvAlL
x3Mr5jzaBhU3jrpoYjGWgCB8yNdZYPJiY4Lr8ck5Xa+WtPr3cMjJ/GmqgmRBX2xc
HQP0+pRR/mNSUEL0VTOy1W8f2Y3JWkRZaEaGmuiTNgzIcXtKS6K34JdH2+JfizgS
Zy+Gzfa9W/pODWYqIqmRx5CGbWRSmn82V3/g5fEtUMKPHNJB8D6x4I51ziBFQkm0
h5uzVsXX5OrM8UE5VMsSnvOublvYfbDQOuA0D3NpSYdoTC8lOHnkZe1a33rI400K
iGn+ltwOSMzEVSXsY9tOE9Y0rQ/5wJZALMHzs55d9K/g4JHaf5YJrhOV/ns0kJHh
b7BwE+o4a8WGabC4c/i6mdgcrcL2GedrbLVAgLCcB9D9o4MlJZoN9aQZYzDNZic9
mNi48szQjJfXX+k/UVUeRcKk7So/GvaiAfWURDQrSOPZPrY9xCvm9vBL77ANlPni
1HZFWGEmJBdGdE4jOyJA5WyT7zthpO0LIqsqcWpNILyGARie09pozzOrAWbkG3Yi
61SDMZ5uOAEoeGOLusy+P6XfSgIAaOZgRMTZWh5SXeF05l1kTVqgL+z6V971fIoN
/q3NeLfw8EYZlYCU38/iqN+LBgNpZCc79dEHg5MyIabENAZGItkP9eCrE+0yJS0Y
o8LtCWu7O+Kl7BvbL1ZOnDr8iL6rzbYtaM5rD74eIr7JZvL6UWVyROTuEFxOaeYF
Kh2rhP9fr5NA+DhTi1bXwurE7WV7rB9qJHZvvgivdoru+IvtZd1mFQrHHlKb0hYY
lK3f6yXWWRjYmcHnz96A4d53AxD+uHAQKrAeEuwt8ymF7NPHUsx9zmrPYGknn0f1
FW+T+D9R47qxmzj3FD77/fZbQImWDS1stAQcLZLJIqqisbimsis1Cf3TUdjCsLh4
ne7EjRSkgtXJcJlynnMGdrcDuMpRa4TdSypvALqIpe0pd99CvTlckzLCiUVsedI7
lGBrpEV21YnXYQJ4W1RnQinHdF73YkeXTzN/SiVvvuXJtyFNeP4/POZauGV/sDta
6FZkST8K8qPJlcI2YNjEX2lpaomOI22nB5spnOjTB7Cpi5hNzdMSCd2n5SAdKJnR
apD83/qB1dkL+fja/TIjbx8uq7ovdI+bmv4tYaLhVKo4bNhDfvHBWQm9JzDs5b6V
TFGGGO+KHtAkViRU0LXPxkI6GRv3Mb8+nPQGnXORM/mrJvlcIv7QzL/Zut39cRmG
hGrz53lxtsuGtbJybpdE8FBXRSE+xFS+b73YkfP1pA9isIyAYqU2655SJ4y1NMd2
pIcHuJEhItwAsGtrWpqiffUCJot9GvuHvwis8jSad3WoVihxHuiyhTMksHXhLjot
Fb8UeHQrAxDh1zfSi6TxowO+Kc/m7Qepvf+mUyP9bRwx8vuyop3N9hk++mcLx158
pt0rWYqJXxeNvy/8rEfT25nu5gxcy67DGqW+0Voh7JyD+TMyv7zVqnjvDsFxGpB/
a1/1miXhPVm8/Dps0iMM5WPnJpahDgCJ5EuEynCV2R6dwunwUnZe5BGIe5G7dwxk
iG6SudzcHhqlVj4Ryf5cEj0hdh8DVVM574TEzcH6pTq5Yk1AEihaL3KDgm1owVX3
eJg4Vq+7Ortq7QzAIeGDBYK61KXh58QJvp7SNPRl/ww9rvqyKI1wIiHmnhfhe36b
3aSItwLQ6s6aMpwMFLPKiePkR1AuKGvDvuildq1UUs4TS7rvA5KYjW2muoCPVIJi
N1cCfuWMKLeBR93O/MMnDU4MnIh/JW0Lxb/kK3iDNfmJNpd2K35ohVn2pAPHqu+V
BuOAzz+Q00wB8z9FARGKYzVQV75WxDsviR/fqSfkNTX22+6FCpFK98K2IFFa40ZC
04JwcUYPK3BFeFyR29xOJkYKg8/dyWSfbMoC13Jt1ct9+6XmZPu06DOwNY95xQ22
sQsOPKasGdwXFbkfxqRmio4me1RWDfVyRW1vrYHBEM+yw4+W8x4gQf+MauRdd5gb
UPDdnPuIIpNxI9IuLHq+3G/o4AG3llChD1yXqSG/YUdTbE+oAGMuQOMqhcEf/xhd
Ys0SV96kPn6uRaUeNGeOwX4xnYVwSPu6KPpPT37b/7Hm4hplhwNwxqh7Gsr20fNs
kioa0M74uzcQwvQs3sK13CStseNjfg+vRLA8Tkdbuavwfklu1ILcoNfK7O8cHv50
LWuHuL5LpkrFDAC1HEgSgpSncvxLlgU+/3Qu+O2I+rKfv/RmanMcu4QNPL/+LXjz
Ev8xQwpTVXEZadRl+cPjJvCs21Rp6i+TsBIfczenR6Npa+ZxxtrnwXEfqz1ULwN2
qKxvQmcezzeEVQJHNpKXSJEGKLCAibvMBorUKXnITEeG5OQ9UMWGh98frLrrfRwA
+yYAdq9AAhcjN31QTnZZza9B9WHMuY0+kpv9tM8q48pcTp0/OYxkfk5PdERuIqDY
ydfvDjPi9nOdrjpmq+2iNT5mz+/kPu7QH4sTDL1gjO06EH0/X2UNsfXkuacxtL1M
u1BFu8CmasgC5f9RN7QuEBeO9f0WJ+YB8DNWz5TdqMe4me6yfelxG0kehGu6X/qV
sCEbCE8mQ03ZpOZZjhf3UPgryEWqlwucGAawNe/2tqnf8uFWdzJP880IE2mPXY2F
O+9LN8vaychVwGABEvYyonUBCVx2vAAV+OywlByYo7hbABPOC6RhyFSm7icDiA/C
9IuvcwDMPeLRtim7wv/KBWpCummk6h3n8jwn3ZUJJiaGdA8Kj0hstKKyiVBObaqE
aB9Fd1zUX0/BXe7x6kv1xYJ+YUTw7WcincNMFD1lV0Y4fVKxVD45FAksWCZATWZ6
+4LxTECyZN9SRuA5EJmPJ7S35wjRkujtLLWBF4MlsABFkBokYGr6EnhY/jHBbSgz
jb5tBuFWN84VEwgT2Tsf2HFK7ZeHKuew9uSGBfCHDzLgRrb7NeNof07w+yPxNzqr
F+ygTPVcPJ8dfwF43mIjWLqRkddRYQ523vrKdeYmEm4TdnPxp8nMPTfs/rkWnf3z
PmP+hS/2+S2JWBoz3UnhUHLmZGlRvzXte/vPVSvn5bzGK9tPrPwvJ0pRz4ls8y9M
0JIaZTjJVgii5X1kC4LuG8X3qbyZt0b7OU2eIlZQe0r9hNu4iu2w8EwCCqvqZQUm
UUJeCeA0eipUIYe4gc1Hvdj1eiboserK1xL6/OIgshuTOd8zTVs4SKzwXmqcHDIq
qzcdnboJEaoQHm9SU3fhY0drXSP0R/p9nFdfi4KKcQI60UxhcDL+9gE8Z4LfwK75
fC1lhM5Ek4KmH2IfaZVwZihNVjDehwAhjVCA4G910PTGk7yfN/P0IvOIpvUbdHXy
17K2LMrkphV762DnMcGpFSB+clxbLcSVDLaspYwKfrZmJf3bVRM81/IT+aRmdTOF
DCeMck8Hm2V1F6/o/EYd/fKKB98lTvbmmRA1EjJo8NCKzCA6etAxqXTaxEzHEyL8
fgQK46fc19Kb9YkIGhVRfin4QhjP2z8X8/k+XybCnvikceyjaO/o7eBQqvbd1Yy8
fqyEV25O2BiNgdkXbshBjOEYGq41obP4YqRIFCoNtsPNERh7XZFsndrMsIl5di9Z
uZc5+KS1fdnxli7sLLnKkmQO9YHWg/jjQM/uKVvx8mUcgPcNistVKfqLmKacMnya
Hcj69EAyPs2Tzz6xw6BJKm3o2jBGL/vn5ORI+B702RajLOD57jWJm9/Fs9GWMj/z
hGsPiV+0BL9K/9j3sDappIYHkWmElwKihModarfdjfXO0/qkOgvsoPU2CAV4wWIk
lIYvvJrQnP5eSzg6o540edze0IlWuYxA6HmafUT7oBR9rBu+XMs8+76vx7R2xP5m
qqwyu44J4bBMGGi2RpOd7bRls5S7q527QnT4Fc0CQ0PNI1KCAc3Jo7t8iguX0ROt
8/uTUkJaecpSyQyKoshvIesOsVjK2YkhXKiXk+l60gIrarHHj+QTYFUAvCTwnXrC
cy9mVK4pwnzFfYxUgl/O7hu0skgwTA8CIgFSPfOQ07sMQH/FdxRBHiuGCC33gj+D
wUEkOlv1WwYS4RHviJxvAc9k/0piWEhT0a80JC4M4Iek9uHyC4/N2UW4eJXh/FQl
1z7eQ8D3NDPo62repT7l3ZtfXshQxyLPS0ewVUpc1oXB2AP2QlbIwqL2cRx0Dza2
EXhdUlGgRgiTE6+4PlN2CzP9AzgeXn1w4jAd4SsUVSALphX6+XpV8K1FbXqqYLUX
tXo/1nsSRfooxvC5LnTrsKt7ObOZ84Vmq8gYczXD7TJcMizhaaUylb/m1DgFPCH5
k0xJngy89xa0IelrgBq8KsF8um1OOoMHTmKMQ+9shPu/LdA7O/8cyiru5fASRrDm
up6rvGhfa3PEfEbBdvVHcrIEch+CAubhMF8pkJfNSfWdKRlcVbovMDywc27M+W15
wy/iX3p92rDRHxAAQv75DWQd5UCzWDSHb2/oGF0kOqDee3s+7/Rhd1U79M6Jzlgi
ZEHL24ba2dyFsmMYuTU7D+5Y1uUrbbD+u0pQn0LcUid47RDRJ4wMQK+mjrSzhiQa
VdLCTS6vS6XxWGb/JjIWQGh4aQi1EpoDuqNDQgxv1KNS/mvx9gEsNlsr/zyNSlr1
d4ONgcqSuHBQUJLtwYu+TfIlmt6cIAU/aQdm6QAUNKJJrNQYXKGrfV0wafuwNT1h
PWlBTDEsZUrjRkBA01d0owSiBQNNzGP+GoUPVrvIbFyr2uPGJpGSMgN4bNUpnBYX
AjZygXUEoz4BXvDpMNO5jgQczRVMnQnBwRSAJ9c2cEcM5sDiljE1XCVI4litcTLS
J3Y9cjh5pnzYq3ccaTe7wvAFUwOb6h0hPsU4kn0t18OeSgUsWOXc9yLcoVE3H94K
fMqeChFggNwoW/rjn2UG79h4kK0G6Prmv1hl9p1nEvXTxh+7XlMBmjyxcsm9+F4v
3QKsK7g3YFU0s+gKDccg6CQJXYJ6kvD8pjOwNNgiM33lKaEOLFm5HnCiIx9jmh7S
gK3HMelfZlm6PpiaPMYt80X0P8AbaY/mQoWWZbIldbc1++Ws81nWXDBkq8TPg2fg
NKV2A/NwWrusCwxJoiOplhsoHU0LYTEWJMCUYX5jOTXg0+5s/qfk6cx4IZLTDH3H
myP+heodPZms2L03oL3J84BcygJNaaNGfQDb1Gyu6REnupvyG4iv3kqalcIE7Z5m
3FHkf2njLplF8nQZbCyBWqySrQYWFj5QcVqA6rHc91jdLraJ/Y6rhWm5F17JbUuQ
1VE6Ki3kNEpYftQqt14l2ItDzL+QFNLuRrcsSulK7kZpAyeKcXC89Vfzh/xVUa7M
dCCQo+XboXAR869kdqc25Ka6Sg2jKQX2WmrMVUu5/jOL2KpwoUm1N0v7DbIoZBAN
/ghhaEE4yGf99dF6stf24gepGN5kcOjGwRHEflEzbluvR423TcdmX/3q8YkH7/Fr
PKe/07XLq0WwaRA77fdVoAx9V3nS2XKCSOK/vi5O+2JevvPvRHIK87UO8OaYVoiP
6psInO8vRmrgz36vl49z+VofVGFAkLnNHXItBlLOc1RWa/tJE7M04VLhZasxAyRU
QXBNcydCy/mWhzBcpt3asPLyle+aBm0XWTy7mMpOnJ+M2m69EH/5AYVc7Plv25zu
7GY8to63tYe3PPlEKaZm0H2RKb4yAjPxMoh+orl8FmmURYRuEzlmWfUsM8j2sqjR
fOAhxX7sXO7z1hlGx3E0utg2wpEGGOFpwsl8sAuMUjGjSJR0iGMl/86DRwjqjOz2
P/Sg3VP9oaCl73EjBrOuah7sXgUe6bI0wk2RfNbDF8/ckEPO73fyntM/42PUO6Hs
BKTWrPSnUzvjKwCN3EL4eYdZ40lac5fP4hWlHBWJvh5Kw7h4/bZRUDOhMugMr2Vk
y9NKfvsxsTzojNjbpWArFw1/eBKuEEe4P6hMUEIQqg1e+gPTYG1uDycRp7V5/6vP
QJ722RZiRsdtYY1l/QvAjqlfgpuEE+EbpKugoxVd0Q95CtjqH/DJHzymJdLhIQLW
0QByUYGZLtgNTc6mh6Mo2TZgIIWyCQexay9x94Y86+Iw1V+OD5Zmyh6zLkJFB3AH
qhPP1NixuND3AvzbU1Hr9r3hedO5asr50Scwy39k/15LIlWkSbmciI++hbWPWwgz
4pIlXR6gj7tKo6eOewWwX6fJWp60/Z7VnS28VU/RAh5MNa46WQQ1mscTYLdKoKwZ
/gBaUo83XFR7yQvfFOT2ANwz8PFTCs7CcMehdUOcwwKouL0REA4QiO2dUkzQB+qP
IZUK2t92HCubjPI8lc0NEVPA/P1A1252zbi0n5OV2xQlhUMslJtZ5JZEzCuujfKW
EaoXV0WOYrEVleQAlg8aowhMpzoPf4GcczYSbgmIdD6bCSwU9fIYhOloCWHL/3GY
76YPWh6ame4VEfVNpxheW/iMo2lraRUdm7ghms59I8p0iObtAPD1YdKINTim7Lhq
YcegcS69w7AJ+x0paSJa6PafcNjTLLVt4zXNcnwTRfIYCxWkNGL2TDteJGeNxplJ
EdO7jYAKfXO9KUqKIECYRArE5enCjnQwakVp0hngNzZqij6OqmmrWrglhTn+y3j6
vKztdD2TVKpgbynoJf+Qi5ryCZZoF/hL0yfDYd/WwEgiIM/bzXbBJ7fB6jCUa4sd
0NYZbSsIiyFJTX82qRw8kZOx8c/5bPMY1Qw0A+Hme/7Dv46dMBs4We7oGTJm8753
nABOEINq29IFV2sJv+pzOSWz3Hq7Wkpbpl39swNcUXNzpCs+agMSr4J00wOU640t
TLP3fm2VGFJ3H30qYT42+faV+7Cg/AHIIJ5LRMg6Mdar5LmNbpV4hSgWUcw1vIJb
paAF1gqB7/6pWvlzvetRoxOC8Wkze1U+ErhsknBFwNnUO0BknRiy8GuTzj35QFsv
Y/ipxMf60RiGbgKVSTA75TBWqbietpxjzvh3qhg2mG/N0dENImaC0+4eBgjnT19c
W+B9/mp52t0KmyVdjsvZAkrydxC3Bh6D5e2AkmjLX66ptiM0kSpOADzGAuTxkj8/
/Vf0N0cJoofvZlaP4hhFJ4tR8S4HD6t2tVH6C7B7wx5N8f6Y0aMNZd2xuzOJ6uea
/HLY+d0KUPm90fp+tQGx/zjBXkAT5r6T59AVMkG2aFSLfC9bFvQDng0u04fOmsk3
nBd6Cfd9CwLP4EJT+z1yH9i9CaXG8csi5vcBagc/V4698cYNl/i1ifmk0G/uKnup
eAIbL9D7uamcX/hJ2WYriQY4f7NmU1QqeooyMNIBmia2AdZqmW8b6ZLWi1MMI8dd
VV2FkIYkvsbnTEliwJ0dgvtDyGEYSBtqJ21plxFkOVKJdP9gxPdLNZmr4Quj06pF
k7MqXKLNDlB81YcH4uctNlKnote1rhSBmG88G11adq4CuiJQ3c8MLpa/wTehJqpY
TtkJHmUJumycnKhs0H/aJc8NyP1V1fk4xtc/kd2d61mGt3Vj4GQ/WbbXIiM6A/Aa
cmqMFot4VmaQdzr3NZlhiMtMUmIGlWiLiQQyblvjP/WrEx+OQh8If30ExzOdDAuI
qE8voSKoHFPXMm3Nzq8FzDXD4aW8QXDKbhioEYjdh4H+dDrXnmKhn9wf+z2ZLIH/
hpPcX6Imva9TlpplOl+coAIzjSznN08fgeB6hKU1HA3K/USi3UGjddXsOPmJwHc8
LpwBYf2RA/L2j/7rW8zkwZnTYVwrz0cH5ae/FGAU0o7rTVamZ5iTx5zaA6+S7ZH7
RFEcGjARleA8mYL11yFAdlCMRvF4DiA3zFJ2sqcwunhNB2MD41Fq8akJrU9lr+5p
Ttq1H+cKGRp3+B/OvdxUWAKaoi6/MpDslWGVHYpVPyGmEzxGbP+nixWC+m/9rbUh
2T9OF+NkAVto9/OjwrHhobb88FlRL1BoXeKUEMssAxtwiHiMQgAzU/rvrKBp0qO/
NNFtQTfoQDUaCvVw8iY9aoYuuF7beuY5mwDXjVoNB39a9ZhnLCJGUJVOecAcul5a
hKjfrgAXO0vvJd+lF7ivG/ZP+WObDPs5KHYzUbMD8s7Fiayb3NaZ7cRTFNL40GDM
2JzQR4dMaaMvxrvchVtG2Kw0R7XUxVG7Q7Ik1hPg0/OmrBdyXw3HF5VdQGgkFR9x
YfVTo2DE2NW/ZeHL4d5utyj8sBw4nING83LoZTyDVZXVAn2o/nPCvJ5cak1oJVgX
PpifSY3304vI/QXGe5GYfyT3UVPn1naO1l8PO+3NaZPrG8+3h2dNQzRAwrx/0NYt
+bVX5tiSFVy+Z+dgOTlqZB6C+jg5tDzLUEv1ayRhEbURQB9W1IMt1Y93pg8e78+B
rYmV124rFUdLPViEG03SjDPPs+DQhG00fYP0Hhfem4PkSBv6os+NrYSUlxquUFSP
VU6xSKiCZzYVLX2mFO1zSj7fpkJr9V22qD8udbtG4htmHXIVTm0GV0/blUnegTUQ
Lgv9+EI9kFxvzXjSny2dctuU4M1C+753oS2oAu5+NUqSCR6zY4uKVvDRpBlXCUsL
MxtbngaFUXO0iBGSf5g+/gPo54FRFnaCJMYeLKAA7nmng4JN5Q8IDZIh1s/laeoi
8Ng/0J3CIvOg5s6F5cTnjrNJa+k5ScEjp7TVSxatTB7oQEeLHWvYEPtHDrH2v3zN
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6912 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
DZr/8BrRXj0KUruQ2Zf/9sOODBm/9HDMbaX+5gKOC78Dpjm6SRMzVUaoQy4UCXr/
/BrwJETlmJpfex45YRdJCsmr9FW4r4K1F7ZOdJmai6+ac5lq39wfL37/so9dVI7D
UDcy32uKv2VuSZTmt+Tkas8P3Kh7sAWD8lbRLhF8G9bfT0zpFjz2ipe2/zcxi8Ma
yThwNnDp5WU9yAUrrRUEP//NwrHuepMFIUhOL52Bx2B6GU8Og6JO3c2JSZWa2gn9
Mrc1bebUo9fGtEva1bZOSjXxNkChkHpPrImMr/iXR/9TR9nMqtMkk6HZo2kl7yyp
kBxFy6ObfbZyVYoxuPptf1xmjOqa7/RHhEJeLHLOJy50kXnnYO2a5cS1r22X9iK1
TXcYVg7Tdd4MrI210TOxVPJQuK5lWhQFamI3homGkUeE+JaHcbgu1Aw7mt+86J5F
NYZypfopzOnk8qJIEoXw+23/r3YleBKheskxu8L3X31MMaT6d4vAC595BWZxYNIe
Ty3CvJaP7T6o1v3yUIpvejDSbvJmVlCd6JxPVT2pI2sJO0ci0/03/3pf53braBb9
FjnuLDtsYJjV+rl9SeVpHU9ho2lNfdZA2o+DADZyv+SzTH8QI+Hz3K/u794Y/Nv2
PYO6P+XRn21wuDoTJfMpxpkD34eT9fdmDu5lL0AbuJmxGhtJs9mhO3uYQUfjb7jd
73QzHFS7kDfVOTy1xC5KDhg5zhFLyoFBXsT6ousTXUWZboQSepbxj74SybEFuZ3e
bd8NJ0n5exhIqFaRuFF6UBNDhRNzxgzjzzcKkEc0766G+/R/Hvst6B4l/+o53AXx
Sik9zEnYDxcbHIibO0HK9pcOKPqE+n7oz8UTgX3KTmiHF2fl63bSE5QuMkt2D8du
iKgTRRXoBMJdUeuuKSs9/FY9MshoNqv5Euz4RLvIOq5t+RP35vwuoAvg7z8GAqU1
X69aLenzZrD67zs/KIikeEHETUQ2XobGMQF9O7Cce0W6DfmqMaGtl+X3egDdfUhm
Zy79P0b3QEkNG2Acl9v4nCoC/rO2Ik43ZrUP/f+NppF38OAXU2Macn/9ua5Pw6ze
qVpvQT4n8MroVIjrLhis2AvPIej49U3MRnorCaAKbV9TICgbKn9sl/uiGAo5LhWT
l231P6uRWdrL0PvmS+oear6pudjXfZNl80qgFFFsrslZHEO3NYzwxN0ue27397xH
vyhGpLvW6+Jy8wUx9M53Wpw53zQ/sr9MqK05Ps5EsmWmyK1/JnjoSomRnIjbZFVp
fvie9m5FLT0VvQ0+3kuVn3t1NR/s1S+DtbvqJNsjYCFbkQncg1I02b/XKar3i0pM
0fyAWksegAoq/YgMZ/sqvutztO5rDlk4QjXzlI2uKJEO3vFT4G8c1Mf5Txc1okBd
UiJ97GXmBKmvAOQD7TqS3zRi8k/fYsdVuq85jipH/XywT3nx7PSpjZHbFM6KNvfN
hLWlsNQvCI0GHMaJS24057Kw7PD2uJJoiBUdMmd3VgYkLUt55BYUUbSAG4b3H+jX
O+r9hCxnU5TQjcHl7f9+dbHGuAznGYDJRJnUELeSwrw3oQs0c0kksauiv1p/rlaz
+hMuut9IUgTcx9EB+8NtU8+QJ9uR61B8/9ZHXcXeDbTR1sSXCxSt2xiaDUFnlSpy
YWeX8PUV+ouRjp7Ui4pww4dYQTJvCGlNs3LPKEHgPObOBZ1+K+iSwbDsMnsaAk9V
yli+IfSt8w2ie+Xfwh2+syHy/gTpewUbQ/nm/yc5Owfwg46mch4Isu2q14uqdxIR
ljLbVl0VKraZwgm87bburyC7OKtjiqVBY4XWtAoY0+BkqSexATGvHrwv/4DS+idU
d9pfdYZZ47/Yn0knXu0aII76PkS1RV553vSjkmawPED2o1Kv0kQhDR/j89BxIbM0
jmQBEPFAVcGji0eli7HFamb2Dj02W7C6xOtSNx33/pW5Du+jybEeR1PfyGLE9srt
afZNdWIoR4e4Asz06b6QsTFuBIhgicxbUF8QuUno8+urVWRpYBEodvhyfDPevb1w
MhH3ZYaTCrSW9JvRP8x08HMZk/24NKGDpsK/IwYDodEqZ4ABNA8j+SROXHehhPrT
yzHVnDuKbYdTJyBhT1pLjJzRN7UFg7L0g9bRJXvtSqDCECX+HmJFEoNrxWxGSJsh
mCiOC+q2Rl9hhiOMm0OAofjN27fxkt2PZh670Oj4pPxGzd84QLoMlPAOmqXfHks1
1OfQcytXKa9yQg0B1kDanc/PmX8gRv7CfzbTkOhc3GNMWPirmLBvSVE2AK88UE7p
G2A4CTsWrHs04IfBtXQsqajWkXJt5I5bIymDtN9qzTC5YVMIC4xWMtVmjvaRGnC8
o8t94gL7acmT91MzNnYx7VEKLlLOJ19Me2wa+whjirnpZv/GjtGcuR6Ud+GGCM+G
jfk64NAJrMDGJY6opkevNPU9uRrdI9ruuShAeCC3VHh71oUnLOFYSxTyx5/he06J
pbthMEhm7FwlwT6cLw271VQ3pK/+BOdFjnijimnthbR6Ca/FN9hzZ16VXKqQ3LTK
JHDY6lYszmVTh/1eRrIKFqLNVynnNYOuxqdyoZiUWgOhL6aZqxpyXGIQTdqQ1EZi
r1IkY8qvS/feOy1YdOzTV2OoCwEyZhydNo84l/CHQyl625pIxB6kYe41jDPLpnf4
ztaG3AWwq9xRm1J0Hfw0D1vqEzKDJfPOvJQvuOzHlyauTAKlhX7gStXTll1FDFms
coFN2cMEbsa3wzU8IAggGmXkGYVZthUNdGBgdPxGZYGgPMlJdzA8BAuy6z8gXc18
dILFSoFuNwy9jJ2/9LA8czUwuDN23Udlpb31q6S6pcUgeQSHqdJh3q2/kZCIGVHw
efluk3lF5UhIOCvBBzFDUz8R/M/tyJq7wink4XGCrlhG6spscXp1win7Ym1AyGp1
5YV4ie5TwUMNPzLvXBLQIRL1yh82MDruylhSD+6jDYWdnFSYLgVY/8E7RCnFXGrK
k2PrEzQiE6KxV4B0F+ci6nvFU8ZJhfDHlySCjtEPxXacOKDzmfR/bbJLEyDKGZgs
Kk2d7wcbbzZ7HO0MXF+k6Q6tNUg40KwZP7EZAc49TLL4cH3JGPwQNg9P5mFXvhf2
/mRHjcIEU1A3dJODsgeL+kuQZRElW+YFnGTmFAzD+Z44DpipLJTfkVvJaUSy96Px
bea98tzWsiCzqne7ekahApR2RZbbZ7ysaFcwSM2/G2Yp7OUfL6BU7HKrBH43Dvye
eIrr57JPCLBfv9E2mTZHqcBtrfSv2IEkWwBuX4DnhVIWT/iFUwIgaz3JOMJhleiD
AO6YdTfXrTAvLK1eXSgSzKXfmbE5SnDBkYvSVMEOtIWz7rbumxErG+suecFF+n3Q
lESWL1aUtgnLWIL3FxmbrtFckcjfijrAi194dzUYh2v7J8wwaBXfRgR4DfkFMg49
+a4VkMeriKZfdr+mzO6ZsQVumx3A5E+qFcQLxVCR/PIDUZI0PJs/vV9l/UvAVDLL
D+umia0Eq/ZyVnnT2VRkHL401R4ZM5mSRNmkOEzDNwfTKX5t9lMDqXdjNlD49BUy
Ps1WFAhWdyCKcwD0ESyBjQ51pC5p0hrXFmrSF3En679/rjl+vii8FEeeqIi/MSa3
iLKyKFroXp70eF4GSdbFrGmRJYJM28FiaIH9fccYiN42efdmB6U6rlH/nLv7PhZb
RdOzsrrEPUwMvB6VK2yh4yNrXLSJLEzmU6v+WyT+q92iEnzxVCD+rVgW6JfFhMt1
kpqrNLoye3K7u+oz2KBac/Ujr7A1fSQFat3W01uRkcXJb9bO14HyreeIbqEM3O8M
pusXD5epI/j+vhoiZ1JmcQ0MdMexIAWZa+Bg8iEGcExHDeZdVXUmEIOqljn+lBXB
yF76Xz/y+/CEsbY930xC8hcs/emjgnlX7rnjhLPM9SZfCzcvJ4UTV9Imh2pde+Lj
MNRdeY92DQQ8gr8//XzSyLEZ1X68J2kgXOM3dgNmRujtw5saFNZ0zW5i/OgzuRek
KX6IQw/ynk9lwGFF5acMMQ8JrF/u56hi8u/IFHe7No3xWsHBkSBzruYYJ77tvBm3
NHagqUilgejZVykW6ZK62LJ1bwb+4nsIaJ21qS9b/gFa2pDW1KFhIycgpB8wnLZt
8rFBFbuB8jHqxXgArQ+kGZSz9vJQENsZdW+UVf1+7tlo7IHUSaAYSKr2ckqM93AU
H1S8zTBC7T9+UkcQH6qwOdHU2+ZtZK2v38Rb/NwlCLqEQ5MVQsqiNM4JZk/zUTxC
rWer9iz8Wwz5teA755tK98p/fZ+xvTLiTAZsAqGV9mDflr/EDTIJkRGW4kav/ZDC
qJQzSSVlHvpPA765tDnO84PYa0gM2vHhM6iMRR1lVzmL1nEU9T6/CUbMfCAF3qRz
2aXHFR79Ff/5NhIcgkkGWd3VQM6SIZ+u0ugiejzfRH2skXJfHhE3bTGBbW6IX2zD
gMDD0mw0UkE9+CPxOb5PeNG6cHjoOjKfs2yVB35S1AvnM64M7Cpw1hnpuucKriIT
kmkjBh7XdidRjAWphZpGGFUbf33M4hSp5Fiu5n3A7UkWDonVK9I/cGQQmchD2PCS
9M37g2LbJngUNJ+knfvVwHLW3dskrrrm0tSmHiC+slBh71ydb4B+k8ihftZ6enCR
2oCxyGhj+21YhPYfl96hWE/jTzNItg5miDgkjxKQMw0gDdlXJ9dreQZBC27m/FdK
akK4ok/u7GKsIZtdy4L0SVnz69LH2StN2ceFSdta676jrUT86U0ERpFOMwx5ZERJ
k3u6G0QRbzAfFr9VgjJ9DyNoCozUq0fqdpbxhrqCKFdYpuewgCsqdiINJvcaD3rY
HhQcOMqzaGg1qdp21eV3XqvxyU57wgpw3P1FLQms67A0Ykek2HCYftc51rU8AJP3
W/XDIEXq9p+TVFRxZaeySjl/tUo68i4KD4DZxTiMbdVVf7/qNQ+onbrf+sYuHOjX
pJ65gJDgyviW27EY9FKUZgfXk1TD6k0kHpTBLS9uUycI3FlwueudtzZHFzGn0dVz
i6cXvPlfgdQyNUvNbW7/p+olQPli4XaRrvqAcQiXBKNteImOe/3eF2xMdb3U9ZdN
y2jua4YMLuVRogOdZheReodPMLgQxroLvHnYnuLcYMYma3xmdv0iPC0ODIXtSYX6
Kc2E6obKculeYAsejTAxarYrcAT9yRtUwYqO8FzURf6MOj62J2xFiwW8LwFeKJj+
/5tbYZCFWBpHEp/UKZqdHj5WEFWQCYNkdgMi+QO9lFvwfv/stLnf0zVkf8qmlVPp
y0eJts3CrT/JqVuNkP1p6QGbEILr0TOqlHpJEkbtqkOouv+DlnlPHh3btCDgX5r1
2nl7Kx+SFyDaNFcPCooxym2jKJdsasFLYgD78jxQRDWIv6VRyrdNrFr/W0L2wn57
V8Pjk/z9SPygVTg7WXU0N/ejqpLsV53wKDk3A+ATJ6hmgikgkekxvdXTMuUGq/rN
HVYEWKPu8tXwVSFU/Z2x6NGIcHpgBxZQMfAvvogT7JxnDXXcdAOasImyk3zP+TC4
TcM3FyT94ENxx34FxUvsXp72n19sauR8WYHMnu3+YMpnj3GZLfCtVb2bhJKjHAkU
CV8JtfsQyplIWAo2BpW8UU6aqe/C8n2SaZo6rbLzqRxAcDq06d3U/423fxcZ5C9f
TMh6/SaKZBaRMxoojd/rrHcN83dEDaXbMPQB5M1vfHcAObgoWvAkGeepIZpQr4K/
4EeQVaodL/y94UsIPWUoFUpGDkFRZ2BTkom8fWdHAG0V6AzJeorOu5Xxs1kOHHG6
uui5W5V/wmPunxUkhm9S8c8BE38IratOmr+Ct9D/peLBRlKDUq/lWinQ4XvLwRB7
tD/EVFnb9M+9QM0cjgVtt/ZGQ8dGybmDJPRRgfjxaRnIK7Cj1ct4uiZhRejYz9iz
/lO1a/lWY97HKMVaeQ+yysjsxYLjA9F/M9pad5WVKm7S6G6JKWWtnoveer85OUL0
3Mqmo95FIVHjcKz0Rx0KMBWAfH3jepXaA18kLChfk6JIW71F9DOfjpPyzHA/KPdX
DqsWcBfMkhzsbxhMgx/4nSh1BCZu+lwsBEMrh5ddDWITZygj9yrLQ9LeFyvyvTXy
v9CeaqFZ4RQWY4nBuJWudEDwv9HyuYHtJm/B/EpzfTl4mxxle4q91L9EapdTFjV0
l7DQWLRIJzbcu0fmac0bdqnYBzfDFFsi2n9YflSEG6jCi9tU1b+C751sNpifCp7G
/oJ1AcHQYbo3qUcZpbBjGoTvIt3CZF3S0zfX39T0bwdIgFjrxZpl/k9bsthhqmnZ
VWM/00M/tE7QIc3LBjAsFJc5VLEYNwWSvWxbzHvBxXgd+RRAfh8ErEDvuAyhb9Hz
1uJRGs8H24HEHB+vMoCefl6MGXXPq0aNcyqCykGcCYFhwOuJqOqvhkJsm7e9x6Mq
yBYG85n9fRtZH9Hq6JOlDDr41ESBYCJZJJdxevHBjJ7OoZuuBgBl5s8oOep/LBfl
qSfiPdjBmvWBg54EbxSKnG6NcpM8U2qGrd/KjpBPWYu/f4F9Yyqzoxnop1GeEMC5
TE/hqBeHNHmWWxmxX1K4rM28rAJJypH8ZDCkDb2ClM2JPauxskefB3dPYkZE57/b
oBQG4n/SKOs4flqufLA69LHAM6hbb8OcAeHL9gb2Ao7mRX/KYGBCmfAn1gMsq6oP
QbgZTpI9JpUTtD+r2v1lyAoe/9wzwbyE/5XaMXtEtAayeY6IzHdT/K1lwYzPaAZz
3nnXG6tYi1dgPQXN/+KV2AXdCQjFi3dPB9qutf8Wwlgi5KJm36FXYfB9x3efWfGW
Pkiok75rsa78r4FqMLhqWUdrnVjr2GuBT6BIvqYBswIALIcVWYsZq/lHSz4oJdLO
CayU9dV5DZe0/zreqJ1ofTAtteB2vYUlYdeohd0IlwKTltjEi55wmvrzN6+DXQ+e
59qPFQtoDDK2G8DkcSvxbNfHStKYhdZmgkJjMiQxH+y1+k59nyI2rBJJpAvC129S
kkjZyJ1S8vHrXUwwU3C5RVNZ5gGfutZ8APnkBmmyPCtXDdLMDyIJUykCgVBorpv1
tFM/oNMSkOKmR7/4Kcq27UcSUskFY0bzsMH1yNZRtsISDYcAZ11U5eKhwWcVaAIa
u8Lf0oFZbvUyt6bgDlm731Nwm02fuBgh7UCSlOSLw6h6SYTx5s5CFcQpIZWNBBbC
IrpCAHaHzXhuQ8fnDXo6plT9yx0emVLjTVSW/yjwv/yC1jXwQq6T7/hw78qG+hJI
hF9HQ88YU/khDIp5ofcCb9VZIOWaQJAkpYEU9wvZQn6PSrDn2lLVM4Wgvhs2f1l0
oovLSkN3oEL0I3whvpmbJcCZ1RNVlvszVMhrTmZhLyP2QOFQ8zgaJtWCKgZGThHK
YOJC0ThK+4PkZdpECKDMdMikdRMztwVO6eWN/fVRiKPUXNXJcgDH8AffKD649eCj
KalYMvmUgZxc4qlooNh5GczJG0NrOtmV7Ldx5eVsh+fewFLgzFh8XaasdDUxv1BS
qRG/yBp3hzJjal341kO3nj75g9wbogAvqcxdeSOxwPyq7xSgX7L3G7e0WHAMmCkm
T3O81LCktarPratSJce4PnsAJJ5byke7wiDPeBH0ddTbMpApquu4PFhovSvSGD35
Yi/f7iPjv2jUJCyhhCuQbM6YSMaSTaXjkkHZVdTvSaBRcTnLfMgM5xDbT6MdYgno
5P5Roxav/+hImeeNFauauMgUnz3bj1LWy0lu1t8uAWGBJcqflNUwETfimXp7P8Qk
iKxQXqgSvaQ2Pk4kau1uqAqDuKvPhN5axfyE3r1WgYGPAnX6B+JoRZ8L0hJAo/L0
6uXiucmnUphFuGCVZJcHTdZ8Xv9MjD4H6OBgIDzBwZg3e81mEPuRGwKLjxcdVwSQ
BZdfQd0u4Y24ro9M3eewvpHy6HqxEj6zH/TMMqYgzNVQgO6DiGO1vdfCS0GcVc6Q
30iMAOLR4awirKVPhfSW0D9C/MpEWfiK4hRrLP8yq6qkAe6547C7oPFzkDm6tzAN
g8ZnASP8+EII3+/zDh0v9A3h5HVFpk1J3vVccbL2W5/gvXMA2UjQ5lOA0YdUPxP/
lY8aQ7XpaXFrPBUegNENxZTmpQTM64Bw3vrB9FPoBkx8RekEaDCbuMDfDzCafMic
sZ/e5YVuc4bhwRulRgS2q2wGyCoA7rRQdXcxn0yOrMIfogYOoVlNYjGTN7i/Oqyf
FILcc9HF8QJQ6CW3SgZMraTTi5CX1qH48dF9EywvvXro7qJjgaXLmCP0jYpS/Cvv
5WB8+23Amf4Zx0O1SV3XZCemokTlkxrCovyFDaqKUxRqdZ9PWF+hgSEmCfcZczP2
06Iw+ZQ9vHbWY+x3xHeky6U0SQEDvwdYk4pbp555AZqHKQISaT9b+yf/Ap7T7Em7
oxadqYfFRkHVCBvWcHQZYb421laq02zu0Gtc0o6S+lYQlRG2bhcENfGyO3nAnwRT
THvSHuXnBgjbLK8IO7huReprK+77t1Q9or4feKE2a48iTyntZXCAF6gGZjtPplSo
mZacJWxM3yeh/WrtVX8ONn1aPjIHpnI8v1iL0BzlHpm1fZCO3OchzuGfvfmxCgEY
zKBg86p4oV8LcQR9uxAI28HN4DUCD9qaP7w8Rz5loqrVOIFzBnxbsd7K78v0VADn
ZpEK7r9K9EsBhBHehGLASmAXq4VfLll/FiUCuf8EvxeyMFHuePszio1FGtKFd7pm
TiSIIbb+FB/hOlSulJSggxeYKMC/rmohbkQhLLq5EMjwCDc/JOEdQk0ycJ6YZzDB
1s8Ie/HOep7+5zZcWV3VRXMiE9vhmamuX/nmfYi1pDD8KjTyvjtKqWht4ayZ/HTc
gfP++PHTGHvuvhL8WD9TIab8NVVNb3P+dJOs+yp+NSer8l43Va7FtAHvUcyZTD/3
GGOedC/YTOq0nMAcXpsAWpKaOXai+bd2DTz/tX1eG55BDy+uGcQzVfnRpzZilPwO
mr6EP0YFJQ4gykjwm0zqXVj06ico76w73UBzsLy3GXq+pLlBgL66bSS66NhcAZ98
>>>>>>> main
`protect end_protected