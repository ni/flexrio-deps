`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36768 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
BpTGUlWg2cHZljFhnB3CrNuEXgmNxVhLOZiqdeJY0IRCgmXpEfbRJWMiEQArkdng
Ex1lKFG6wZw5l+u1ksjQhHYIeWMu/rEppjPpA1J7LI4lyxuZV4usDomGTY8zfbDY
KvIzp35WXvOG2JSy3IzNKEGt0VbBTsT+NX9dcfDRtwyMJ07c+n5T1kRsh5Dhkq6I
viJwa8hxOJAzyZeR0ikhdcOXj4NIGSCKa06W8WjKp1XRav2r77fpfbFoDXTvL5UT
rWNlLiB/coirpP4J3lbxHs3eoRWvy391EvHPmauukF1m4Qu+BCxUdGpxWCpsZdl7
XpfZ0Q8p/DS3UnHp9NXJUz0f+oeeyuNLpEVNqwCNQETgIT5XODClaXTGHYs1AYx/
blQxzQoZn8MFxF7THqC56KNuINrjNk2QffBrGf1x70PbB3gNwbeIh2tFQmBU9Uek
eu59d2w5DY/cv0PHsY1xx9dEXyNWzOR4ph0eCLrrY/bFbZzAEixm7pkydCqmt6Ik
lVOq9KXLs2aUynD57yYLdKw7pi4S8CaRt8EJZnYVx1g+F1JKFwIU53c3sMg5Ab1i
8WdEptXE7qedpFdy7q8nf8YRi/ZE201OoUAo5DH4gVUJ/ShoMvjx66O7HTYVtzRd
I6phXGZzt+mmv/uTpsYwOm/eK75EiWxWGWrxgu6bQ15BHYt8VbyOXscdssRiMsJN
JtChMAk1pBozosTIf0oPFL18ipg/c9Fsr4PEarIyNLfDgXo0LCnWP84KMOpGjnsi
AReg01OUbPEZZFZIpe22mOycgrA9fkmogcNYuhbpdHjVRYST7LIaKUZ3BNJKPKwo
e/PcAEoR8Brl4LyswujWVBnRy1Xi5Fd1gvTHrgtLLe/zomgJJFW+KSP65ofo3DUt
LojEfrZidMFNxNvr+USsKZKIm3mwG3xXkmz51puem7tjRxTYH+wM6/yxXUZsWpcH
evWr0l5iuv8VKJfB+rV5dhC/hAH0zuugObR3I1UEPfnMRklS7BO42MVuOzC3WCVi
N4g9eL0utePGCbLMkVHTxzLYejU3YnBPP3jXi3gkecEBwNuRZvH7b/5g10vvimLg
z6f9LxDBToglJzKyxJpbeOrABit1x8giAscY3Y2kGO/hEvuZYobnP3maaJSyQbGa
6sEuCrDp4yF79045KmJAjQ+YSPv8eiwk4csuXYZHFEbtoO7GwldguuvLZJvn2Qct
638yKJCKnKk26OTjPr7zTifwGt4P3vrFjFoEH9SvtZ0YmW4dGv1U/ABh+rqQStXt
/jmuNaBGsE9k/udkSRCM2nHPRtMVYEbqwJzn+YJ3CLAaJhHjNwZNw24YFQVHO0rU
gVS5p7rGWhLiAOKEqrLUZN+yt1qKNjTV1rjESoOYgplCAbrCX2wb1uswxruPAe82
aQm8YIVV7/lQewm1lz3CDiE5PMO2RQTrmw0kIvUgjwinyP2K+heyPMkI6OCMB+qV
tLb+P6KmsyN6ToREF90I+W8m1ueesWUz5vyH4hTdaH3LaXZkHYfUXLLUxxBg409D
m5ejUIJlIkvmQxLyLV5l3KzuZ3kQcMOMHl408b7/wT5kEky9ImgujBSraVQQ8IZU
rtp99FoA2QAEI/CdMj2BIAadMxWI/RCSYawe648jJiXKeOydHUqPDYaahDN3GZ9B
VcKq2LzbXs0zgXKtUZcKbr39p8FGIb0xqWplcFirGD0Tmut8hvHJhG8WGB5CChpH
Yv7VV0nRjNsJDJuVmMOyz4M5qY3TKXy1fgGpFaZWyHQ040zlRP/vy+4PJhBZmPFg
Byscvb3/navzeoaAkd26AYIt88hAeNj/eYsyInDZKxLph5sep1TF51aOGorQmXVt
cV1nR+ckXPHdxhG4RmruvCqj5EgMtTjeXwJQneewm1PVKFKOm7OvSikvlvBCiWOm
EmL9Terw8r2XyDunZc7pSCOLKmkKFoTCblYcI1PyiBXwjqrF8b3MztiR+BTkW8gc
wNoH8ZBbIX2PkGF4oDzwQg/giI6SZ2zqw5C7x2t/0MtdQKxAUrZtXruclk8h/EWE
Snx1AMhLRA75nmam5/kS8KfMjAgsvwSV6lBmQaZWgqMUGIWMLCG6evteBCUFTmgL
ZKti5RI7dSW1HCziO2EEKK6vJblLPghe0y+6OoPTR+dvohZ1Zfu4x6ZgXVvM9ppk
3kJ2uaR3Zni6zncxurKBRYxc5ggRRzsJAlZTcRSzZgN3VWGbp4fr1qyQkhFIPQzI
IuCYCvS9Nb6ayxyp6ccy+ntJj24OtazFTJDS5OHxwidaOdBKbqIkzAJm0vx8xaPZ
T6Uq8uZuJy9u7jmZogjBfjFqsR1jVTYy21bNZzntF+Z8jbs8Z6CA52RoULYkhzXU
OjT0bxsnc1rRKHNV/9lEVRdxvVJDZFiGQeM5bHEha1bbtakIMWhnZJkbnCY0rvZO
zcsvwNvqtlez7FJBMzx0RUy26UxMf0AuuPjI0S6SIlut4JuuW9ZuiLuypTdD6fei
EM0+OPasPXaPcwCq1mNY4tAVV4Nz4/nsoykKrjzTtaXuLdqbhay96ebSHlDGd1Yf
RpB3yZaO0vgFILCXnuppO9MUcla69Zpx1x7hMCKTwtcAb9uAEAGNyZHtmf7ySQv2
osHZK9rW7ieiEg9xk2gAHwyZuk8PsHybRaOg6eBY0KAxj1o/FYk60pbH8GU6ms5Z
omYZejKBvIv7lec5nzl1ZTvMHidTjqGteVtMBZlOgknmQKem/PgMidO1BKKBGYOy
tySBwux9TlDLZMftm+WZ/UpRNcnJphdXb/bEB7mfbk1fLlG7ivGdEgUqEooBj97D
kakiMr7MCswGfQS7yQuNA7Sk2OjuUEpxmMzIDalKJaZK7BK/ZLGdk/41WHLrClAd
lZBqc9IGxgq2G1m45cT+Jv/qvANgRp6du7FbqwfS0YP9Zn52v3aOsAK0d5Wefg5K
KLUteSvNxQGw6eRFWtRBIfY94mN0sNHVKGLWZE8UdfknkjBVOGCZoZHR5LZL4zPH
NJd76gd1loOWLvbe7v6JaG9bEZ/eBN+KbSxeOJXzkpHtInV2MUD0gKIIrzzqTgXz
KTVbKgsy3luKHmO1igEmZn0RdTT1XDwQM2WXRia33RCCqFvMl4sw7w7rkjbgCEsO
2ki17RuKgybNmyjlQN3h9DucD12kjYwyd9O2zf08LRljfhBnZB8TmZw/m5FEfEh2
11sIpinWkc3V3fm+cP3xLXghY0Qx6mbcIEjpQ6wNUCaNZ9dXpUPh7n2OKYXtyZVD
2UINAp08KWqzgTfZWCitiYC6yUV0A49WC9YzCWee3AKGI0K5z7BAgtlzBSNOnLia
PUaT0IE5vktQa945uVXVkSffAqubw2+p73stP2xLnQrCWYBGmsIdoBWr+MhUwijY
EZSRVBLVAHvX9MPt1pngGS8uTM7nCqQgJHd1fu+LyeVkl8izRg3BY1QvsnS5GcDj
20PsbWzeCWNqX5By0PhxFSfhFiFUaeULJsMFSdWMboNDATHBlyTWBzDMXp0zkTxC
JMBmLQbluR6joF7WqryIrZuUgzXTWhmAArUaWB+6iAe8gqTxT0rXxp6OyCTPf1HD
Nti7r56sBJhZNvU8FWDYC7Y/O9KsEDhx67GOHM5RU624mufrl7arsNWqATm++zd2
Hj0CksrXGybfejkyXsiNDyHMgC5fIPq02rU0nLTSEyXStPPet2Pm2q2v6FlHb/FQ
+a4kvawX9riel3sT5AfxnfLhv5jsDG7eLVZG/1q6LLSbV7NHc3CFE1Nbd85FKS6t
LxkU7hRtvT7l8v5fLvPxr5irOZCSD7Zlon4qtrr0WnKtPxNSW9amky/O+QHO0FGJ
ddupyRPKG4WRKHSWnsD4w+wRB2VCA4dmse/hMG6jLFl+TseE8cgo7xiiGudJQmu0
CkDRSlQyrpKO/VJirFrbx/oMrSMkyHug6eUZVJnmG65HdPGxMAzv2142PfyaC+fQ
G58IkF/stecwxCCSf3JqfyLrXGWvVNroOrTE4btIzN7MBfLSO2Nf+1Gi/UkaEVlt
3nIo6JPu1EvwS0qkLyzJiU0LGe2vzfbA7HRYS8aSxwmnxHGiWHqaRXnD62dtfgOg
KlvAYinX96hcU2EzWRdE8jyYr8UQ8JmNIGwP6zcodOJzniRhOTVr0AfOx30UMGWM
DzgGglbSKAGEu4/1d33K9fYNv9jwKEVRFwB67PFRs+Wdbu6t4DrGUacq5+q4DmUi
fwN6OJgfM4JbyaqeAsAySBMXyIZZeT6+YnUWLpxJlCfDCNMO/8rx12diKwPXw5PI
kSr9xf2iJ3hi98toTsG784mElOIX3Y/ks+x2Nec6GiMJLnlIzITkauLEf0+2fsRc
XHSbl5taUVi12xuTJLK1c7luVlt7VQQKDQ/qB8wUuxOdw0GKKi7YKYtOAWH3JquG
1ooyNO6VzdF9RfTHDKu6imPuoKwFSMK8XHGwUJ22Y5Zd0++hrGNh3dMQqWY0d3S7
sBBtup4ZkrB7wsUt2P/rVzv5fNplPG7OAvSyK/8XgVt5XpxkM8s+QW8Y3+AhFyd4
DbhwATxOvUJejiPWvhlUcPwb8vdLae4/HbUd72VdcjV51b2qvppAfnFXj4660mxE
w4QWi1YoTbBj5Q9A/kT17HU4zVOiL/2BJVP/KV6kqaMQcJ3yyppVFRc7jUkMhyhB
rpQBV2VYayc/rcpknEMEK1E40LIgz7mU2n+IbjsDz1NYGrOdspJmG42atxFjTq50
ZpSKEoUh7uqgP/7jT93incP08s+lbA+ncwVIJdfhi52IBi53UsyV3DOS0Tl3fB2M
8NwHKWGOJ/tAbxXjumu0nPSXNt7NWPobbssXT1n7qSP9VSf1D7xET2YSSd0LnUCn
EwRxhcnIrNXoZjq/yFGLgkjsiQN+SfmFJeyQMyumrlzuQxIuBywv1akybUcBLKmO
dFWCnnMM11MznX4ZNbvZ8Z5CwBHFURMXt8MV0MfxRbew7pzKhEPpnpZuhws4j0j3
+wi66xJAJLRK4lEVvbtbIYSGNcFMv9dist+yno/B6xEs7WcqRao3peohYBMKkHf6
IzHy2V7YCR49fc0mWl/uh5gamrqcg75rfeJOQAgA467VCjYeTfGasnm5GD91/lVe
+4zcdsARt8vEAEQVfamA1rKb6L3lp3/88s+omjxvSfLbOWYcwgIbHtMkaqNiuf4y
LJUcpxjpA2yjd/ViJ58DgY8fp/9I0dJHieLs/poNtOwmlB21dtz5/CUsrTsZ7Dqy
S+3IOEcB4y5deQnsyyt4LoGTA5cyGJBxWPTheyGKPol78hiGZPB/7lpdiHW5YfS0
+rJPE8HfvsjBGhZjwesBmycAj+kWx7hZ9OHWgqqZyRkBsRM4ffcN+bh/7dmWWxqM
kMCQxSWGl9yrUEfHBblJnSga+SzD7nfDzxAF4NWB2d2zq2X+QoVU4ViCLOFGXsoB
IN90idnSgQJzuIj57Z1BdVevjAn8fyDJejjg2dR2ccrrm/O521MqWnUfvdlA1x/7
5WG08WEUSaW26kAU/TfPxS3usqPnKqO/otwrqlseccTVRtiPI4tKDq27a9XJhUGs
u0e9uxOaUDbxsdokyXXxWYfqs5TROatAqA2UTvJh8pMj7WdsfEExCqpeOrY2Bo1N
E+44/5cOH0fLeDZPjd1tc9L9sLD8e9gdaPdnaL1Am0l0xz9qTC8MTZ2OqVEuaFeC
zlQ0VkClSGyBTDGdTH4xQSumse4maO2DQA2xkC7sct4DP97wNtUlHCquSfKkuGvT
NTRZ74vP3sXPk2CmsjTHSR/WLW9y1oBbvyFBQdQv4D4+g+yE7UZTxY8ck3KHvB00
bsL01HyLbu8KzUOEsp1gTE+Wk3/W+7iaqb/l+h1SzwMCOTgC6M1BF1BtVeGii/4Y
kmmvtVsmZcuBu4ohDqYfQ9HsLrFH0u2eo9wXCI1nHFMS1jUWDbOWfVfSf9a3tMGa
cx27GAGbnyK1G1x+c1EESHJLRlhk7o191iykzY2wi6j2lcNLFIePtnHfyRo77x0g
yZKa/HXd62BnWEfOZgZdT7EfSMczW8CdvsIc/P1zqVO3Hhp4l5+mP1/JKXBoTnlJ
el48IrcH9EapXjfcmEtfJgi+TDmK0MMrtQdPyKjRm9ygcZGsrJ60lGlIs+o1567Y
ozbExFquljpe9ttGFusaYe4w8f5GYlzdidgClcw1wGT3K/gA3fXCYusz1waY5QI1
pjCeJCbekIKF0rwfUkq06EBQpJ1y7SK7hReLTbY/kwtY4bvzU/ZLAJ6xohcmZhnD
lzvs7Dn6WqsW77sJ7LOoUH3ePks7pfIDBD517kk9QaLYYWDmuB9ohsavOiMnbGfL
EGpgE/0lFajV2l+DpvlReP/iVEYQ1pW7ctvx9UJFlk0sk+vAP+oSFr2rRNNFBgri
KfIY+i5B9tMpCUXsIEdtsWEtk77NtSxaLSaGmxZG7bMChq/ThaOZzzL5hW0BGL70
i0Dw+slkvHIwssaV4Y63BcmdMbymcpWe6kqX1yo+Dv2fSymQhy8CTufWEr+oB2Ad
yv2IvHwmNPWZ47I+GsPsbkT0levSunX21+89k/jn+BpNadhVWzNo+ctWQ0HWZUGh
4RySUBZUmh8kxKMuht8yyzHXk2HmzVFe1MsFdYsuzzLOliizmLsoKjG4yE+1mRNZ
41iy+ZVLSHLWZ1pfe0N7Oh37UtmxzVM4rwBbm+pknMskF3xthouUHzuJ/m3NaMA+
2X8Llc+BRXWkjaGVFLzuGq3gFraYLJqR2C0sAcohJ5iYdeooRsVcTnEVQxW29QTb
9ZnnzkhCu8UrIzwrMPwDFF5pVlh0vwjqmYZCgrbVIjvbESV+hpzBOIGhe7nb9PsB
ZJaDmqlKRi1R2PXIrlp4fVDwVmuaBaaqY6HohshQdDLBC8CADFqKznEV8Nk/I6Ax
AzVxZMUW3dEd1QIXVzsGsG1+EHmvQw+QjCzYuLumzQBhfXVIScjH61b8wCf+qGju
+nl8v1Mf1cZyPBhdab1ZfRBos0x8QSH2P3ypJdkCqH5dyvLndJyJf0z2mBvTdy4j
mZUXGCyYGiWuJtFRjVmVW3M7oxiVcSkq0T7JoSd4CR//A9hGf59eOHK/QOz7uQQV
f9LgnbcKCSQOwJ30fvTeK3quKKXZxw1vlYo78s44zfGleAPq3qhxqgJtwbza1E0k
GIB2wl1/XPhkceccLdYe6aaG6wZld8gRWVZpilu9iM7X54nxQfT2YQQdEhKYYUTv
/dbcmxkkdcBxX8upllAjoEUmuvTJ4c8Ut+IDbvEXeDWLGVeQHFbepjREUIBeHi4b
uUQBadr7fteI6FCEEZlTeVnZJ6gSwaja3fPV9hCz57LUep6oLVSiiQCypsjy+Ypl
7dFhHMPxnmJuDTukiUZ19KiaX9D0W4zggnFEBi0C0xOAC5kFIZc2VwyXtnOKjGZD
mwLTj9wSRlUB6TKmdlRmCibp4uJBTqOy/Fwl459pHuUBbdA1bcnSAaRlN6Y6D8Lk
6MoDdr0xweX36/WIn+2rg7BLDxrrZVJ9ZLF1Ty1gNOgQFhoFjSWApFeWIgO6+yuM
Vfelmm4uOJrP35DiwS9uOhmHh70hljUjLEzEEJt2QFcud7GF0M4KDjLDZMuyxNOw
4oUsz0vIIfw4uJw2rb6SG583nqIRQGWlffNrWBR600Ap8GqpgNNxPyoplbYbHbKt
Ec8hE6TDRsrC0Ts4WX4EKbr2Xv3Y/ZL6crWisHir+acVxPq8zTdYm/ulfbB3rUJ6
kWaATmW824fvKNL9wB3m5JTOacOPWLJcaCEIABk/74a8GEE++O/g+CrGNrCjV5Gw
5XWSKDyqk/1+gxcpHw7/EwElu0qeOaZVW+B/Hi6dOwZXqnRuVZZACAA4B14MXrUp
2nSIcYO5R+/6Ic462IVCJzWnJY1PJh/i3QaHM/gmeMEh9eGuGVR7Plv5QuN8V9rI
+F90ydsSbks+85pUPTiIgzDJJoblA4iJOVVQW4fDtIILpmU+UXoDV+YInOIXDDdK
6pJ2Zsu4WHVwV1QvVDTdIjlmcOOxEhMqdrFQBbfs1JDX1GKb70V9Z6eohcpaCoYw
8OtKLv8QhPdBuGyNQiU71yUfnLBBIrypXyGBFyAfC31Ok14HGDytaRiba4keMOL0
TIHezcOIMizGRavVQONV/anff8TBpgCoVkj9vgZkZ58uy7I/bT6JGFFD9w7HhFvJ
jV+t0QAe2RT4LUr962qnz5Znyz6gY8b8AE5QK/PUk5SxdeBGQA7dRwQ3nssYQ2j8
xDIeLXO1VXrKxAHoLB2c6bcEJKKyarnTe114dHo5v9QC3vJ0gabERvL1afyE5PZJ
aKf/U9kf1aaB9lhfkKPlnLhEchrZDtaqUN1WK1OmMbhO/T3L7ETNMRmkVXZFPT+L
abTL0Xt+Cfr9CxaAi9MshrTfptqYuOijiEaXvrV2yzjPFSpFh6+ydQ4f8ZRgTsSL
7eX5NXPxaeN8GQT8/TBpIxbeu0LLuAcAOMDvYS3dOzu/kJdoFvnvx6L24IOTPArm
Vf/By+I3Kp+xnkwI1BL1/sH4lGw7nlryQ6d6373tZAYR/C24SNt1mJbXlS31Icb8
MbBkYbk6zO24uEzB4DBdsPCUAjtexAVkBPlqPEddlTInSv0h8uNMpqQn1jbNjBXJ
qPEqZ80i49HERo+mDFX5cEAa6yMVYWeE4pUuQqGSPWJ7QOuHqNuepZvVKhc0A6LN
eQKoLTV7qXE26ySgmoLBVYD9uf1z67hkmvjQ5eDCgWvRJqw7YnvRVI/v5DK0JbJN
uGbQjqKNvocv7mRs7Jf2h4JS9+YtMfGr9UtmB6XdPYuv9OkxMxzfVU9LvFAzBW29
benGHb4VhWyATMR7c3XG0/FaTR6KJvTfT3rTfi6+AqANz4Wj2nre/5JUOzY4IGB8
pimpYU4AIhL5uhQrzgSWj7AUH42aEpXh0QzO6GNxOLQdSEq7JAJS99vHfUHlGgnI
vFw13dDWNGCeLJsDKVsm7abycagRz9qdwgqgPkkJqLsHkrGQ/QW9JTJSH5aJTHqo
uob+BIfXOtQv5a0be2Hae3Xp0LPIZOEZcZAJCXTVjTuOLdusV+EBKs1LnHYAPUWx
0/r1zC4F+1A1o9piVAedSGnpmzbTSJLBzoMiMDCwYZ2P2MzEfqvue1CZO3Co7t90
Y2iEbbKBNf5i3eVQIilLUIkLm/jPVT4Twd/oYqccFoeHzzk22cfP7uhzcgX8LwJ7
KsHH74A5BGchLEjq7iNP4z75083I98apAadfMdpw7rlgUj0Oo39VmoxKj5qxH//c
bf/Mwmj79pJTc2hq6aPKSg8GWKLchU/c1HnD09dKOyAu0ojsOye6iGo2XGNCE00t
Ja9pxZniFfFG4u35chncq2sRgpnHzH37AqTqy/nDe9LHoukWjfMvChsirATeEQYy
toQVhsyp6z5thRxvTdrli4Ug3IC03+XKMpn+7kEKNWpUQDQctzbD+uKTY/kZMBxu
uqzKCWYyK+riDDqZrVJYpFMXSzMF663t1rg0b0z053UX30w7FldnjY0Nc/d9yItS
L45PXg2TwgOA95TcTHw+f5WEeNH1srxrkGjgTJhdRkuiBqyIxDwr64g/7VBPgChm
6EJ9138E8n4qMHDPcM825nY1bYYMbb0aJJFpC3iEQoCy6ps1aNmAdy4Z1pcKv/8V
lhrOrfDv/Irr5i7fbXneXVCrTu2sdOec4rLT/NjIDMTqWRLK0Nw1x+sM2zcJq15i
PWQdVf+UblVYGj3U3PXqpGAAgHpOR4ijIAYMlkIm2gFTxibQhbsbz9Cx9w8T6xyk
3gol/x6EmWV1J0YTOk9x6IivmS1SMJ4Hkv85amCxbJVy4Io55UvqsKVnPkni2+QF
Sh4K+kVrBlVTMKJTKs2qWpv3JgEVXrFHN0mvnM+m3uLYViZTEGKTA66Pvfo7VD9I
wJeEJE3ToKFSueuUgvCYDHDIiHwXTiu7MXwvyaQXJSDPbR5eDUsoDI6xaWElcyP6
1ltTcG/Q/VnywBO7CvhyQ914ypswdcHf6A+SfzShRqnaDvqClOwhQCTDyQ6jHk7D
YiATJgOEViYbAzXUnfxVTOBbMBRpj+bbfAnlk6v7ogBU2aSU/l2ITWhcRImANOBv
E6Mg/MJG7+mGSl6x4fb26LlApGK4Zh7jwQ2f/mVg0cSOesN+w5+KzpOsIJFjdlfX
p7p0+73qzOivdD3r5Yv4mUsyoZUrbJaG+Qfajxao9yXvOQP9umWnx31DAasAMTBG
UFrCPHTKy0kS6ZwWW0RIC8s7CHxLXPtU937o/vnJXa8ZIyi4DZxzjO0+FdmLsncW
a2NligXnnuoQmNt9comK4w+SWKfGBK8lzCNtVyfBYBOIiVRt8/uvh0rX9fiBPLC+
/TnrXrWTUs79t9BuNdwgloUsttYJJOtR3VvLP+7t3V4XSXLYIHvRVYbIKNLb5BTK
kCP3KXUZowcLvIYyacJjXRITDidqQEKoYQVA7JbgwDqfOQriGUmy9Tm3KEpiOZ57
dRxwTcxYHGMF3ROdOVhOaNxi3jVOAyK5bAN36nK5SjxiG7r5JDU/RmGhNJxy8hw9
zKttRmmazfbG8ws/PPoPjsSK6VcV+0zm5NuWsaZcd0+4S1wYWL27Z9xcvfBHUQV+
4uz05WWsQbYQCkrvFeZHjkXLP2k8Q0IhbP+kMq2jIQ6k0te/89G1/wvBOPXo3GHC
LCOu2iqeCITcK8LXEwDnhqHW1G+OPGC6ivFelWLtMtEMhjuIrXc7HMvNCWrEL/ot
FEARGwAAalSpbnjtGqi3WD1zSzvXqdyg0cr0/Kw8EDOHe5PcSVwgJw0KrnaYs4Hj
T3y38O8axOdQldUORuf90GH3PNIeBgDmcswSfvWacWK+nwi63x/fxFig+N2Kva5y
gl0Int2lSgyuOQzFfa7B+x1U0U+cgj8IPEKFsTyHUm9doiEig4rrkjhsT5kQ+g/P
veNlluqrRzl/4eWBXOe4Ibx+t31qlSzK4+ffhwKZLBrezYOM/uiOqAKsZ0NNCGJI
MFV/DATaz7qjPwB2GUJLMksq8VahySCZ6WVew5ka0KUfzqaAjVLa91+X1fcutU4I
SMisSkhffXoTfGzAws+XMZ/rEj+hF83vgejcZ4jKDdWTfIQ5ncoFhWcToHXLeKoU
Rk1wWzZ4Ai+6ZIzGYdS25X0s756apDJrioyg2Hir6j2BYdGgqh2ne+ObP66hdtKJ
ktLRAJejcA0LfehKO2RKO29nPHgfkhy/qfbrHomht8MhBtGagadcg+8uFvG8yX1g
TW+J4C/ySe55vjTpL6ernvUu4bz9ad+cRaI5aXrTSGXoCsHe1VwXMXfSAK0sfU/d
qPn0w0dUx5uR2yQWM6BWsQtdMmiJY6ctiKPQg8ull0icjFsKWMJ8H5L8fJJscKop
Ofj4iN8lV9Xw6ateTfxGlkfWrxmOgQLmka/o76UTAe/Y3wPM7xAsM9VqQvUwCbTd
leAN1EgIJqZzaj/osAOKida6x40M5g6oJOUZGaPV2fpa2MXRpLE4ieZKln0/Dssi
Y5zbiXLndUCUwwANxwMumgPjGjlOYkyx1lsqrdeTrC5NKv5Ifz1NAEMj1uiAFIAd
yPmc29XNi+6iLInbYejOFmIDvUCiiryLb4jCbS6criZeIw339l4pdZXaN+BwwT/M
HprG7REPT4/Pf+KcwZFYldumfbHSOx3kOUis7mc32gggk1qDtTSHeo1zfho9tBWT
0/bahEgrwAZaplDaCMzDcVpEZTLNepRXRP/VH0YpuHh447UZo8Fd53tMBiy3NQc8
AnfpAOPBVKKu8A/jwqOZbHHLmplBGeqA5fFu9RNiKYKwbvIdyjm24Plr23OgO3B6
Oh9YiKTxZ0oFMRVSKy5P0NNRR3v//vCDW2YQkSnsK3ruABKZSiVcHOxV/oW7V9R9
PINc12OJ9Yd0baDxbVHZlr00amytNdyehbJIEmPRJtjZtWGm6k6wyDXMnpprj1be
jXnPGKhBeFRGiGEGPyZXhhvW3PE1Pyjch9ehEGSyE66/nnR2H2gZtGLunyFxRLIC
fhV39wMMSa4kqMjr8Uk07K25I3cgXkQX2WV/esh+7FWictiMYlbtaUSgUbzcFder
hc8ODDtyL1RGf4f1539FVRJ5pGqZ/KL8r9FpVRs+FHkKLNd6q3WmegLJDHf8snyj
J+WiuaiEE+3cP82LRqYOeDdB8XEcJ5J5WsWI23DiFtjsEsskRRXTdkyVUWAEdI3w
pVXcv4gqAzmP9DG6oxIdEBKxe6mmqIiAb4pnx6S0jUKMra/8cdkXkJoQczWMy96S
chcaXfKV5ZLi7V9AiB5wpUx/CRU/7GhCIwQtAoM1oQBixpR5/WbeR8gGOpOFAteW
uLzJgJmK+Si+afGo2xbVrUlWxddQL3MX7OltnLgFzOeTIk/3nl0PyKY6aymVr1Sl
EaYuL2CViCGZiUNl3WbjVkLs/xMmgtek5VcNSyp+mcMlT9MyxNMXHa/tdytX+a1X
SqvaLpJTgU47+Qo+03I1IP87fISHsJ/PTG0vaShs7Q/IUDR40DzGEra6aVsY8/Oq
ueNFvHa3Lr2+anuRcXZ6xNjdcyveBs50vyyP2kpPYDIMrV+VqXUartWkIDcosDoX
S4Khl2U7jyVlQfrLC09hSiGtTybY7PrsOWX40afJ+W5SVIP7itWJuZ+CAt6XqIWW
mFlcgskASftSwmz6SfFTCnKAcQtsr/DyZEYyyvAWrWl2f3xDbYdDHUyL7XRi1CkO
eVkFhFMmZfY1qLzx+rIC7dlXqy1hixb/x0Aq/BhHlOnRWTYrSWgSscBFffMOk45e
FIl7cE6YTazBxaI+Je4qjakzQwdmjjSmPEQFG/hQIQCm1rjczF8atYJv7zehqtz9
fmxeEEX2g7oYVewedkwNEPyLydjLwRCW2L8PLZ4JWi7UhUddbnuMdwe8HIWeDe/N
NqQ0QqRoTM7tQRFAeZ+sNx2tQSUSmFE3dJFdvhxm7yOjAoB8X0IDYZ1sstKgQQ2w
jLR6Ey3WM3023SNTs/cRl3OoMmtiqRfcm4Ny2xnNRaLZMAdHOOe11QHAg9CFeFny
lJgrKHt86yItYukR5Z/JN/RdS+u0I0mJW8hSzYI7aBR2rF+pIk4KEOxIziYOuSTD
/6ml4vct7lW6XMxqHaX4HQY7aSfRc4wPOMJgbU5Nqy+vV3YQXWuIH0iDwDvjuHPG
1rCS0/kCyxizlTvjHL7UCebLU5GBiCqYbNoT1JUXTGadhYlAHLdHaHNisDZU71eq
EnHrc1GTexlEn+C48zEkgrIHU4xJu2Nu8vwUz0SYwfqaN4jB1AwXrcM3C/XkU9us
BJOwTbJuR7cI+k2F8Ygy/Pc71ne1KsPcyb6/SLRMmXVzGePhUDJO9kYcss1F2yBs
c+SAzdb9vUo2RpAGQ5Urfi5iqV3UMvDC2FUDiaaAbd0BG6vjxhcd8pYbd5+ylZGR
eENixsleusjTwKbkTYKPUMUsoPOyEYEuwkTVc0QhluMZGrjCHICNQ19+3ETKSgWz
MoenYtytAic7SXDmKvlG7giJrdhCQJaTVTcWFPh7529Qlss2Gk43BTbyldVq3u/z
NCknbyIiKro3mhHlstCaz+meOdfCwN7c7Ehvkd+4PkNwZqbStWlF/ku+tw9ZFPYJ
4pLrInNGgyHifgcOw3SsFpLzzUzr+Ew16XjLEpQVy1C3wKbq3xWP0SsGf+FFE6+T
bSTUsdcfxLThTrw8SsUKPKOMyf51ue+YQo1EYhVQiopCXtDR03aqJNOyObpU6pFI
2rLqnhmJ1evigl69zjePR/3ED4HbWr3bSHX4aHDr1NMUwCacfiIbPSJCqR0WaK/L
XoRsgOdEubk0tGc///LC+//Foq6971d2gwAPC4mNi6cqwmGP4vns7aJlBrBdml/g
dyUb0F/wInKKj/yak+9wVPuSb2tW/i9J52NlMwBG1t6Lk5wWxf5Vs8vd67f7AEBv
0Jr01FitClSaIwGWTAsFRyg1zQdAWHB0ZdmRPPQRiXwxdUhzE+MMcJGS0HYgzJ/O
dTeJxTtfvLeOd6oI+bzb7XUgLac3sFi5ZqBGV12101a7kHtk/0b3949Y4KC+8QUe
5oLqoePGlzKqy0WqdlOZJiJLb3FMK29m98hBY8p7yp3dCgKVlcGLj2StZMTfKcPG
uJ1OFY/jFddiXL3dliakEPnR6SYZ2Pi4zMFgD1In7lUXJtH7V6VFoPTpDREVC2WT
PVSZ8pi6KmW9BlaGShendDIsj4MAwjZGaz97UbTd+wAMXfkC3mHsvDeu823WauDx
f2i6n64k877YnyGmzMvybz0KUBzAmmvsBxwNFLUJQE0vmNj1cMfVPQUEanKt/G9+
A4sib9vuG0X/5dKbhSDZZORB6+UHRHNTWDVnloVF1YjjoP+sAtaJtvjuMhCfV0FB
WL8VzskfQh/XLyrdo1CrkzBsGgIjZvatib/8XJUfZhCjbaJXoLy4E13QExZTUZ9t
swo+KmcQAFg/VPPYTcojnj1mY5IfbSEdbnhHO24FE/gE5RYeRpOOtlitdu75PmXc
6MRGknWAjVhWpcbTieIhbYhgb+XL6jppwhXNgLHsYszLA8Z1bVnJel5tODbEagKE
0NldgOK7a/kAMZjqsZP89xi1eBz1Q0zvo9FlkLHHPc1pIeKBI2P9N9bjYIwMwZJY
Gn9lvOBh9LA3gz/Ji93Vq8HCYkwy/3UyexlOM5Obx1jZDwGAxTRva7dCq7uL9P8Q
64X0g3dltHjzk2793fcd7aMOWV+01UrDHrzjLsPXOWEdNPIvALayCmRuXgaShN17
4L+fBLmRB6RfLg2LQ7dz6cF9xEyEbZrmwbnBxLQ7nNRqQ2MXUgpAws5DcpxhH+AF
3F1LltK9uWcHxexTnNt6iTABnowloLPmvktGyDEPGWDqxnZjgZdPxz+/jzTC1MF6
zs8xcHcpzV+QN6A9nwkS8VSMyOY0jUFcMGtPzmv3sODeH1EmKgzLIzz/nsntJm9i
4z5YgZSCML/5E3grrUPnRBR48i1V8xNTNJX7YJKEdfYj07/OyX7zlQQsqQXEvsEL
Y51fnLvxhAZQxH/baaLRCw7lyYPgfBMwJu4GBHUB0D/5a9WNWMlOkfJv4sQT+0Zm
dzXHgM8ud+GBK0AyNjgatyBzOueSCoze8DeSIcxxJojIE1zn6zW1o8Ywzi7QitDX
bM8PYZFanriqUgwblHit+RXLTQZcz5qouTfKcUJcf6vMzBTTrAEXNxbCsno27/N1
DnWvXOj+oCPRVA2xM99TMRU6Nv49V1N0ZxptX60NQTCm2YqS285K7BSBNqxbgwuO
m8LNOWIEIMiMwaxDPSMYfGM825EABdEVkqq9s/4rrjXOcEEkGDdHS7jzjic8C2pA
bq6piZAJhVoc+AvP5uv/Ragk7dF8plgOjA2wCN5gt12kCijtzDQ0jNW1qLsZh88D
Z/bWztN+Poe8vvr1LdJURIBWi18olPOuc95ncrsqJxoWJI2XE34/G1wCn00RrePu
3CjLDxiNvCUbkm2GJKxdc880svQLuLD2teURCYtMKnVEKywErVCdQ3HMKPKOyzPF
G9Aky8/VnWBWAhqwUb/4wJntlK0OrbxYROxwTCqydrCDh117VGqgJO1zNlYAc2Ls
CvIE49Te3vE0tMwjXdIE5fjAwPfIY32EqWg9LiG6pqsSQ7MEJsZ+CYCcemPxWrw7
ce3eRjd7pIqguh+tDYVDYM4jLEohalw++wdoAUZ75ZG9coiNqZ6zLBhUwWOeB5ti
alNcnpSBB8t3nSLUxQ+TGMYWsrhG82m4iCUCYMMnG6O3WkoQE4XksmLjk3zLkBxd
JD5/rXNUXdqnFqDo6il1Cu3qC4WX2uEA0MbirIyi+VGk15Bvsnw7QGLwO166habA
gZ/joEpNkb1lXfD9w4feith//XYXuu6geb/Z8hvMN/UX7eVFHYCrw0BGULiPstaQ
ChAeocNRYBA6iHMkozzVm//5SZ5dQixZYYyZYHBuBfzoluU9dWhf3yH+6BGOHxl6
/vWfR3ITD549ovptSzwjdpERRtHcsXcCJheXQgMrTZgmSxGib5JdrNCkhvuWcuic
LQbHOdYbCK+6jpGQCWnUxh2Mep+jq/hFjRSv+cXrd4xIRDgwSP9YvqUh6nYjkJFN
ddl/lMKzp3i/0izfjonNKOyhOFY22xcn8bdluoWeq8fJ7EAVybz5kwzZc5FoxjlM
bOiDAvmXF0ZOZBl8F6TsyhfO6tP81TRSf+oGbWBUm1x2NxFjtWXCfPV2gR6Oh94e
nUTLh76GA3SdXiy3QEOv28HSbRdwx9/G3YhdQjPj4ks8Ow2qA3cTjXez4tDXFdNj
Q4frKyKGo8udtGuA9C6EZYWb7lpt1mWBt5vDeNS+Ii8J5xb2rVnHbr0k6f28aPUj
CjuAgNQcrJxKkwu+0vutv0A8iW19j5eC8ynwe2VBBOwcLFSRcQgS+bKybX5skRc6
Nfp0MJ33RNwyMoHQVT49iq2LGHTd28Tcqqe9vJAr1yGoffcoFwDlgAx9d0Hh3G9w
IgKkIWL4L5LrjWpS0Ar7ZXPTGbnwmu0U4gPBit8B0jxp5r593JhI0wiqJMoRmmgs
qrg/NXregpRwKWXQXmz3+597SMPn521NqEm0qYoOND9xUUG9dFE9X8DMo5eclgcR
Y0C/NxhEBXINDOjce5OKMU+T2/3JzUtBhNhl9otWaQTIbyqpaE1ot/Rzsc1OTABO
YNokfC60rfL/u5o5eaBUeVjuMhqPClkkfkY+04y6RZZnr6hOQtxmhzEAthV6shN8
Y+L2z77GnowpxTxolSuYmwscbMK6ANspFUQtfMvz8EtJRDWQ+DLduwuC2THKbe+l
6cCmld/qzwG3y/5Ft4Af2rBTjI9smQiERk4ZTxijEOk1kAV4cG16rJXt4HyLvHRn
6okVtFDCYR6QTWjukusaKRQeMexSsSWcJB4YnQIlbRkvjXo64lJhk6YVg/oSBmBJ
FAtF/IQYvKsKH5obHHjXd29r6sJDMGGgo7/FzIFbu1XpAAQtPwsmgMmAFhmCLiL8
x2Vb024ga0wHXto0EhralLKPt+dP2e/13or2CIDpJwrXJxo/D/klZNnQGwDNBlLY
hLKfHZGCYmdldNWI814GMGN8j5J1sW8zq7Zx4hrGxzgAt/T7xvPeA8TDw9DLpxbU
aZMj8TiioUN3BUNe8A123LGiwRDsbTnHB/8cmhO0ZdnLY1Tc/+nRH0twaNj+FjcL
3rdsBC8VJ+bz4vEia+Kr4enfwbTYn4wL0LhU+D480cA2OT5n4BxaBOYKAvWW+twI
e269HrssHA95ewFO9lGQvnh+4UfKrIuPr065POVPpirQs/mJkijJEGysGhOfXH2k
PBXpwMVyJC30+BImn+yGELel0ifXxJEotlV4TRrFQwXmsNA19v6eC99f5QHLl7JK
mTQmrn+VucjcTWlBpPns0VW+VpCkFxBRqUULYHL7g2sJ3GQ99xyHMpmTOglrJ7FY
SmKEAGTg1d2HVYz1XB1et5i5X+IVnt+5RcLVKe9MTGVri3tEOngwxbNTu+Fp5ipE
LB4hj6Fi5/NeUtEPtAIj76VVn3lu3DAKwwniMN5IriE57fmf6t5XCj7YCCfGY3n2
U5exoTdPJaQobJ0Uim7QHAjQTSAmU1m7h+Yv43SQvexAA+dlv5MfYtC1l3vz5riv
UMkip52BB6ibBLWiZIKenlRG7VUudC6m66cemQwmZaGYDHOEUYSwydptqDLu3Dd8
u+R0ePKQ2kdx5W6n8UsjvaixBYsLJjMnu0R+CFbrLQvjcUhp05P/sLn8cDQqAGpR
Wi/4iH59XjS4G6OXqtceYaRmumhoYfWE+OqquTyl/nZj8F8kt89//NmdeYlcMV/I
SOggxV8hjp+pFLfbJjhBn2jiQZevTdmhWXPlyZyVJk6IgWFhnMnCPa+kjgSQEH0B
w/Qai+uTcNLKPH9Rc352Lbymne13O7TKom7eT3VqbIV3vmuXXQEHwzW2zsYald0A
G9JHsSqL871vqcRzB4GIGmqDUCb2Os9rQ8Nc6WtN7raoXq1H2nBq3PKbb+4H+EJ+
jIgdhIcOD2RNCXYHUbUKkJM2WyL5ZQWklkHGIXUYd7RJjreeT8kLqmcQgmNkmeOI
m4VeFb/SDK6kCyMPEayHw5Pw/Xh9jSpypmljgyuIb/nETLvKLMtr33eMRycO+Q8j
ZFwzUPj6dQJ/R4o8wQpCmeOFwjbLQPRCNuCEpQNJWTOvmKlTYLEs7vCdfHS5KLew
m2qQWfDLOHQ32TXl5zk5aZVHXUi6QtMIZTfiDbf8gc683tY1dxnEhPsMoxEGTYle
JZ1XfMU4HAzbjoBj9H8LhaYS6G/HpG8aTgdzs2PWvZjfY/FtB+GOuwBqfh/Pey3T
8LvY/QTTJ/2cTWMc3rtXQI+l4gyALbxT/7bBHc4G5pOLzjo4w3SCkHxTZXDy6D78
qfS/WJHToPBvmOrfV/86Y+mtmFSw3pLKkExTG2/u4284s3fm/Td0BUmjPDvTT2gz
yJt4VYC/s60sfkoYBnn6ONeccsVLRmM++3gfNFrMcWnuHrGFM6xQzwWPQUSx5+Gg
AAsDkiJYzpWy0ohpCRqKHl+YG/xzlQT6lnrmmOcOrKlDpB/Hk94iaR3i8Rjfs5iI
dU7sNB0mmOl/Y/ubkuHzsmRtoJHJs6abcBmd5JiCStnIgrE0yy5W4qm147axliB5
oMUBaA5cVnxJobetxfeM0pwAvd+Fm6bxT0lzeP2VOTGDaIKOAg5ZPi3R0m6Qrq7R
Xn1eFYNNvpdRKtNDbwQuDuJ2QUTBO8h3UlQg+kXQn5dvPsVhEbAQXQK5zqYLpHtQ
42aeF9vEKjCXnyRyrUgCpkYWycTArHneOoxNnTfyQ0Q8qbz9ZiJQ4SILiL9DBZvd
3d6iL7C6ocbgGU4ZWfwetW8fwZz8EZWfw5oxcu9PWrUkZGuGO5Ln/f6wDZ2vTFVt
BPx9IBHU1Im4t0h2TMtQDhSbBf7d6GDTsW976es1s9FfESH/o2MnMMsGeM13g5VL
VrlKZ3N0Oau2nzRSkd4uA0rcIYDVGTJcG2pEWLgWIyImWA5eBKeFI6SKdcdeIxFn
soXZgu+ZpUAJBVRevg2+qmNsPNB2XgjC4YMGtAbHvbZP7y0ahboAANgEZGzY3L3o
j695iC2caIaYAHbnlql1Eqm4g7KQ/dt8R2iTtErQYMMu/khFwPDb57ezpnmDlgub
ZjA1B1+w0iFwJWrvoCQcuNX8q58Ncud2nVpQW2pXnwA6Ei+n/KCLIV+ErceoB6sR
etm2TFwSNiuD7YyMU6cjjCB6Jq3Ui0HEYJuHvixBtRTO2QodjoLSfjmptypy00qb
7/jV9sJ1PAw4i+vZj9IyJwhuFn5XTu7wwHayO9uaBUz2HGsaxdiWxJswvKfgy6Q2
K0PVycmDDxPkjjWK4XhfAc0HfP4Nd/RzhaHa3x2UxxyDzo89Ro0iOblK7FgbjJG7
VwfZRkjM9cGuqnFy4ov7jeuRC/gftapK2y3MpY2SNfqROgqM7xgDWVe+3+ERMDse
abs7nDHDF1Is27V8QENfG6baEjTNmZbwySPgJ8v/mAkWbNWjylhigP8IBlXhw9OZ
ecFM8jz+QBoxQpwPiVjGh6yvTN42ZCi3p8L6XnBQEqhipDv5ZlzR8XDgSswSegkA
0XWn0hNvAQeceitv3fzWAvWAYDSXHCBg0tIuX/9UiK0DiI4HgrT/F770F4jxu2Uo
9TF6Z1tYvAmwSeGXHLF68OGM4Lg1I7Jga955gX3lTtIe5P5Ul8WBFI89Ymbb9697
JrTwJte6wCZVnkm4IdlKneutOi44Mny9RjdqeZBu3Ll+6tQNSQjE5+CbiUHHV6HU
3LG/xruO8eQguuwOJm8nnhuLnLSK5XwXB4EcQGhZPQtyrQ0IXiEJI3K37UkmeZXR
j/dHc1yJb23UmRrPWzrk7iW0YIn02/WdIMzfhaTFGSRjQ6gHSIsU46Ndk1KizfDM
IV0Kgqx9VhWyT5z631Qpe/CkfD3AaXlPl2oNNPMJ+7QjuH/zmIy2m+/XclnBhiWY
b5PnWmQ56LcqzXj834ZPh9tscOUVj2e+fCmxEKlnE/zWd2wstXd5i7U9wEMSUdqm
jMvdibNTk+QXB7PVCdLOutU18DjLAkf5alINHnBffOAmpKTUNTmBNxDRcIAtuApN
NnZgGT0sro3zaRalds/oX37aFKNQi+6/1rMdvXp3dV/Valj1IaOhhKF77e1CtvRn
1uZNObtc3Mm0KbugKIetXvoqcIOjlbjkTcz8b5m6BcmJ2flSdtzCM9UAvzPeylcS
IhfpRv0dXb/+MjgSfZibgznVcyLZPMViTdJameUBUIArRaSki56qOGH8slN8ErsG
dvP6F9Vif5lXWUtO0hqdOzow1AvSmgrQgiD5zKm1OYhmWo8qv6GYNgQ1FLeEb/lV
fFxEIngiK62Xpi4kdvOYpoy1GMK9KsPKDLRjtZWN40BLsLUabhwNdlcefStJnTLu
Qk0izRw2tj3tQTooN0ZOjtPwCsIui2SGjYPtaGwBWniKbuU4u32MAjdxbCvzA9cZ
oiUeS1FCu9zwR42p6eNbEXyXOaidpxtEPUYz3B0S+z+YwO1prpLjYO+Nx3PhZnrM
6dh51EaaJklbGzHmrWwpPmywaXaPFTiHjNuDo1r0W6HX0wqzj4C1MsUL9thgCcPS
G07GbIyECU2DVXObSwPw/fjEzKb/FfHFfi8f+/jFj1M+tVMhMA9JzVBkvOJDXx3D
e/JrldANVvF+gLdOm8db3eW31Gmeibf+hmcgrsjht9l22EFApGcYeT8YWaJ2bImg
c005dML9FoE+ioEiKGuvh6OG+54IuXPVkww6cpr/w0D+FZHloVqIrMzGSYl/o3aO
M3Sd9pVWSpoXvj684dKFeXBwWN6zN3BgxL7ufXTcSwEogUm0B6/dQ3PQmuHM7a6O
fJTbTpWZlya1JLWHWgWjop+rXBZcTREXtkTxq2NXQaaE03j0ehJH+xjjb//JiMVp
lAVh+fp4dJKzJKahJZaSB2Yu/tTXJlXqHBR4EiccuSgmmZfYsArCQYlK93q28A8s
epZZYARCtc3/v163wJ+1qp1YgrfF4GXQV/ngUcFNNZWRjQEpDRPxEvB+vQ6UM5KF
93d+//MwhS9Q54ZLI2DbLwUrPxcg2YCL6WC3zazpjxA2danJkFFVFx2anvmRQ6lG
x9F3AXg7FN5M4Jsj65NHJGfkh760ZqfkuQUGy94QVTd37h1783iEytwrHHJ+jl/T
JxP7b/Tx0BM2r/3eed7CrHtuIynktKVDi/+hIy+R6jOWQT90NUDhVsrwMzroYfGK
KqAaAZ9VWjcH9F2kqzEkKdcKk6UHrd1KyLjjPce1XRcUHelymuV1cXA87GEwa7fi
Hz/2I37PlGA4GIDGPdW2TWB3eQCrBvuNHgBLEQOoldaHfQwNtrhwMK1qKx3D5hNe
6WrQzq6mIsIPuP+WiSaKRneTun05/KggajEmjBe9Qpcx+gCALDniqpYojnpi8eL7
Pl5F/xc+53NmStAhjqFGcrR9YP9ZJT/SW03ht54m+IH4J/NpNDcIRlAlqGhEz6LG
etn0HOXX2z7rfD1jvI2oCGs/FjKgmsor61UmulXf7WTfEop+L/OQiOvzSFPbFvqe
FSm7jSJlZRVpNoClAp2+2hCftiL8lXUSJ+VUhmM2cbPTEt3zwP563P7dEzmVzlY8
JiGD5v40DWTUNidFO7un4bFphcNaE+sv1v/8s+8ODI+yYuY0teaz0h7dulkTfYkG
YcZsmUXwLpZ/9sk30NoAOdvMIdUmNvmL+Jzy6hjrCJn52Ns+bLdYJ2/EGTXgv3E9
RxAPynyFIqjYwUqi/95WPbs0ULzHyHm+JRLpFFjR3h4jJyMYLCgEOjqvWldtBSRb
SOH1eh4MFuDnCDCBFmEwp2Nvxhbea5D6gOXvQhoe06ZNxrfR5+w8BRVs57qsqhyt
CKi5gzW0AtA9vaV8DCh3qJ02p0LvwkOLaEG6t9Vsco1Rs0p0DuC0fL6L9Fk0gOpX
zDZ5QFqHauMPd89JXH6hP8OI9jcFwCSmChd8KEYZooyKXeCSKkpAcy7kvZvNsUzI
74ktKf7L/sAHeYIdlok/JALTnhHY7avjvaqKcOak3WmmhFta0mvQCAMa2AfKrA5p
ccgrQJVto3LkP2QciHwZWzjQKmtaBjx5ezDHMKGDgFqgTLYfmxst3sj0F/4KUpJg
IC5NQXUD7xxbWg7ovI5EdCOyjIGmmJB0IVC1UyAzgvFdcLwuIxqB4UDCO8JrSgWG
GsPV15DyyqFSyB48h9E0xpbD1VM/xThe2EYAlteGXcpZIdLvmZ/2tEaDCyWUDRnM
7bJQyxUG5NLd42T2VWNi+5atqeInwEYDoTpMcYQZP+4RvQpQ27OGMQKZd8rtdhPD
WFq/3tRI5OGfrwspsZvB0oZg7Ws0eZOCETS+/X3MiZgoYLzcw9pHAUX083Msh0RH
wudttQREl4SwxVq3JFuZxpeO1ORfN+cfyAirLwNDcI6DII4jtFwL1x3xrHif3uDH
JjOvmRFxEQ2xc0rBW21PlqXyHBil9qZ6t3pBltjbzL5yFufHPWjoGWGYnPngpPH8
/fQ9//gzQdk1bkRWvlZhFdUurs309fjVkx7TN5iYmWVjOtxCPNTJTrvcuHMML679
JE0EK8YLnLRBGUjHC2u8CFJS7ro91nKtQ2HUxGE8DjyyndHrQRJNfZ22cyw+kE0/
hmhwYwsuC56ql3eRIDUxsc42x8DmX+SPkRWwaIUTA02m1KqFUXwqIEVrrFd4xWtp
tZepKBZp+0D+6SFRqtwsltUa2tdgApot16UYJsBr0mkOTlQOPmDm6bC9iexeOeuo
ke6LutsYAkaSitbPonmc89hN6UlfsIgqeLmRfJlIyqU/uJBTiYjeZfTKwanSWTae
J4YclBHJwMPaSG92vFl0SRyn1E6m+VHPNSomsx0rlu7duSuG2NSIWPMEIg6JLr+o
4wWSL7mLNg8n6J9wWuyXVw5SrlR127EL7kpQzSW61cZX5qSvdfEGf+hTzMv+zKg3
87nNoaLzRRWQwRB6Ph4ehGQxMR8DbksdF/JAO4zUnhZRZtgLLEDEhKd8vNtQcF1c
d2OqdQGsYyhBxQF013yWGaNZS4V26xBQAlK2AMcyxxUXzdlLS+77dze297TM4Iaa
w2ZVMQqSp4mdUdF7+QNvt/w6Cb0O32qwhiiozBv2RwmjQzwiMiHZTs+j3SeDYiDR
KHfGESsm4peCwbXTt5Gc1/y9HIWOrDxmiSBN9YR693KyW2LgHMjpEK6qucDKz8qY
/CbNaTw8mDCON5lvnl7bWd0qlWOR4YvQGsiHavvvVvumxqBDjkp7HqQCUYLkQUK+
neG/2jgG0EVWAq+iqiiu8w/hGl9IS8RPO1X/Ccr8VwPRONZjFgJEM0V1AEUUgmYj
H/HKjKkpT3CL3aktMDJm2m3of4ssxaevFiIFcu8RRnKwsOQrwuocz3LgMByyOVqp
IYMQS0EygCu1922MWo8hHYbaBvDfeJ1AKzLPhpUwu77WmC4gWozvt1os+G3oYoR9
h/pL+t6wDaudV1AVeph92rS7Z6EJZ8oFfTdy1rHHg03QxAlD2ZuX78H81FS6sJuq
WRfT8JdxQ7ezW4sLKYPT/AlQMyYtTaJs8SHyrVQ7pEFBnvlXg/sQwXnsSg2hzzKB
UAFLFs4O1JKtVRVdHswEW6fOTfnbyhUF7dqFZil168G+r4PHOTXM9fOavxEHMjjf
X7HBq4JXy9mIIgqYsEJuQlgbOmJLd76YSkfn/r8xg1iiOXsdGZrBtQdGvAlWxZdV
RNgLB0xGwY/vqXerBaGnBwLhctaiorOCr6a3/yDafwFgE1tWi5UUwABT6LV4Eib1
tp1zPeRYYDPU4xSbnw22lERNCPr8plMvw0nhpCMq87YhPTeFGeKWCPlyEzgJz72w
1IYukCyt1rJYe3McbOP4iAKej7EMQTnGZunaJ/psftQQvCmfsTsp3She0q3ChAqK
1ewNvKpzjbPVCT1qpnbnyTO0+bxOsBO/ALbtXyFcvJcg3meWHop9590SSXEW++PA
FgWtzzPoFkCUKMjcmgh7HwvVauzbZWVtCYJxtnoCg53gx1ossRmmksK6Q3pemWSn
sjbqpNFKUxe6Kb0sT0JKs0ecQ/3WPRrh1+oMOEz1m5ibUzegO+v3iEUYREb8EhHA
WQLB+O9bSILDIx+8Um5KLn6w9bzbtLZzGbXoqNTDFOtyXKAVvY8j9fizw4739VMS
zCRF6IvgAwVZOTUUVcKwCAwibmZlFPCRyCowIRvu52bcrgOGVawEZqi0ic0NDaIq
mCTa3d8K9E3R5BzsQtm1AwtLQKsO2bQP5Q2NUQnz4uxNjT4dCY4l25I4IWf7O57+
3KYTuosaRy5aWLMHJd8DiskkLgMMItQNdMh+Q9hHjeKefxA6fg8h90oLkeVwm/hb
cAM0aEsE3oPHk67t5dVCuSNsKrvuQ8vrzqahekTlz+XdrJHnayRlfZk1rvuLXQDH
6R7U/aL1KIxg34aqBj7n6LbOXUNZLw2xraeHIDNYVcZAsZ6j3FMHE6PHaDQV8WhD
3nTzJfRNVUEN+5BgJ8wbVE+DYrmpfV/ydkDILEHPU0n6uzMA/qINYUApFyHztgot
CstxkkHJKdnOoboshl7ag3sG0szt+gE6OIr/4+99fpMB39JzU7iXkNbpEGPNDcWk
5UIglZBKBX/J7yEcBgi/2NEereV5Wxik0ScVQk3QE4hnLxQ3rhGtERFV5a3n7qKQ
Z2bl3UvJftQgayPiYbN/CAsEMRLnEtjO1i08P2Gn5Gyl5L4bB7WxnzWEqkzTPQV8
tGllf0Ewc0DL+xzNxfTGVff6zAUhssAbs7O949TkqlTxvMBpliaQvxTTqRvDaZHN
ei1M25+t/X8ablD+OvL46dg2HWDNTRtq5OiI+UOrsPpzUwJnI8ThsdaLn3vOoz0y
+gaHZ3VUduZzsBfBzLtoAJusxbiK4hfNmquN6IzvRxzzp3Dgdx/h0Ngg3E5LX6bc
nyVaO9Zuas7YS2EaI1DOhjeU3pc6dED2hW5ykZZkJitx0wJAm0TBCiWzBl6uv07T
FkhgAPw0GRpX3WW/lmWc0vZD+aN6HQHsLhb9qqeiqykXn2QhGKEKC5yrbD7H3AJo
MNH/PEwplJ6dsLGKWckLN2/r7PFxVX6yK/0HHLNrzugpFnR3AavbFHdlwfnckQUY
I0Mw56CHMnn5nT8lRK6/OEnMQxcQZ+PtCy1tu+2v/iYMRCT1r43d/sRv3DUB13lM
F3qKw6IREu4SsJH1Z6tupqBYKsdLdM9Yhq58sQU7/aWuQ91oW1+qvPYfwoWmR8rv
+sXkbDj0NqWNSwGxdlqpdQtKItQ0S/ZxPhgixcMnbBatdAKYKV9XpaMVwas3WD16
27mcEV5NCxPJ4oNfw64ZZyoHX49/wqywyP3Wm+yU47RhQi+bppglWh81LkqhV7CO
yIJQzhT6f+TUpZTzK1Ks3NSTq8RlE6uYMwsQ+zMZ1I5a21DCx0FErgipw8lo7I8C
aiferWulIVdI82cJcl4JZ+sRxHTMdgnIx4CBuvCJZQANm97TkCXNSnFuJPjDL21z
zsOgZoS3F+ERvebF+FSh7TOT98Vv8eHN0FYfLV3fYc04nUS7gQRY8we5RrdJAzyn
IVFu7SGoUaTvnWdyd+b50tWRD/+UiGNCK9MB9JgBkFORjhDj2zujthePTK0QOfsu
h29Pdk+80p1FLaLp/DaLgaJkscI1Pmk1/MUlGhivQwBIoQjo0BtapaFGoOOB77St
Nxzoi0zl65x72e7weHE7kRMz5VvDGcbYbNKsNtzC4wTitXkqp+/xgNkoYP8RllDY
X+ovXraxkHrelyPAuwSPg2sc3j0ak+9WBpBMOg9ZBFP/vRuZjLMWuJCDif5fMvwq
20xCsswAAWTbclwTuxwbs0Y2s2tia9W8jBa4hR3sbJrg0FRkQ7eeQI5dlvpIbFQH
or6wT2/nnN9qWLTMJ52SOu6YiBLqZnEhqCXzT8Fe7EsD0GmJCLRsiCsJBKvsZlUq
/4PJ4RgfkISNx8SkbvkjniZohcjrO3RYzn/1BMIt9uqYHktEuNYalQM3vAvkB+mg
FvZfZm7rf/3xG4bQ17E8cKlqOI15U0Gw9ilgYuGpg7IfyZAKUont9OieIHRW5uF/
/tgxCR+CV1ZTCV39EwUY9QFsMThLlnAsBYLDGD84Kxt0/7itGT89QW7G029ng6sy
MTs1AxFtlmnL74qrO20JeGQrx/XuMrsMbizED7ScCwNybZR/pJgY7BIkjdPA40gu
H8gVVlhG6WAfMvl2Oik0LP+FZITwzd3sFLUBTZsZYqrXXlhdjitGYy2oquPKHxGo
cbyok04dyTmWINbeLm38KuJf8HA464uCTF6aP9rA9O0nCTwOyZchA2OnFeKti+fk
4+dv1VVHgjDBcoMkdqmPMzYc84kZAXk9wpza1yRlOGonhwYg8BGGFkyv9mwiYD7I
G3Ob4PLrGGpVCnGwv8jsCi23KUAaDD71M5hVIpP7In35bhMChP37wWWI6COdTC+E
eXcMMieLPpb2bhLjTvcwnDc84KtvHJzAa/plZ9lql9HovGhUOt+822y9TKoVvs+k
PEHbywKTucbY3CNH2VxJwiG87GLfF84LOk67Pu3fMPMfQN3ElrpxktbTET5s1Bw6
rQuyWP8x3Dbb4F6PnduLUH/GlDWk4kkc37hfGKUWp9QoaROy+kLp5yEZ76xzDp5G
G4xZMH26viUPzt53SLj7SkmftGt9XeIp4Rhm3BF8q25dNp8w+g4ATGHC2FaeVfL8
Dke9+UfGLaHK+/TYJjR4e+Dgu6M5WW50rAl5FTvPmJGCTeSokZYi2soPD2CdB65K
EAd9Wkk+LAPP+XV89zmRAEga2Kl0uS5OTx3KGSabl4tDxFbJllYjQLNMydNriYCm
CRj/Puapf7ISOKuIeBJPMOqjGHgmZDd0i8cfh6850fnai9aevKckX9CgQeqhXOkt
B3LwvYxa48hC0D014DOzMUzVbh3N61bWgq5XFK+d/78NlVgZ7C8nsb8IP4NznwZN
y/YVBKBkCsr4TG9jHvXAyyGQS6vnqTWI8O2+iT7WCDq14qW8nnSQs7/AYRVxJ9uZ
Xzknu5TPTOJItbqvF3ZUanKtxhRgRrVKYflumowa5CKKSlrh7MhRetEfto9hR+Ov
2TZSTJq1xECoYnHgFN175FKJ1Ux5T75i+8mVzsLDXDNz2cdEXDAlOuuV3W3PxoJA
zVBlVpzC2l3faNzfOTX9lTMBYiDZm5PeCg1X6+sgeqNUqwE0PkOzlucSP8GuA4wG
DuENh9S8KmH8OLltK9iT68ZD2P+1n7Ali9w/fKRsQnB2jghHd3DABOHhoCjBq76n
I1wD5dsGbtPHooICEzDzIXz7XBqzlR8sRjVGx+28fA1ELiHSZYf/twXBHnC0ghDM
/VdXu3cV6cQe+Ba+uHPCS39af6DKCsn8WId9hnyNq9Ia5ODV8x038lmLUFGEtAzH
sqqpU2GS+rm8L9etZZfnXWDUXh+xxFUxWZeEjoR6QSWfe2YxKXVEtswvc7rDzMSf
rPyJUksqAh/iamTCpdLdzDpkHbGCdbHRhfUlB9Ld/ClgmBcszm66Z2AQJ7iGMN63
6LawGkI/q7ECISd/16dhnPSygkd6EnDOyt4tefEAToWxZvr3u0IrRMv9agjK/Z+Y
evzdxJEaz54kVrYHsNlht7Pejg2yHAI7qnEJRvg5EKWpHPx0/RPi+pW0Q/ovcgOI
IoH8GbYozCipNtQRX4bPQWXeLOP0z377H5tL0McHI4Dbztxs9Q6TZollMzQW4QPb
trySU7LhOcw6ky1h4+u7y4GEkpOHW8YfiBP3wtRfuXMfv5P3nLzzyfh1fYhcGoDQ
JBJOU/hc2fSD8FzSU3ypD2VWPePyCffbREtOpicw/1v9/5XNOk1s7UeocJh0IoAX
61LeW/P+F9oAqQ0/NcHsTuI0+p2NAN5l869h2lxY+Bnz++Ss91jrGsO838RJ4oCo
JjVmDlMi3Hk/8HyHgifL6qlO0lfWKSKMR4HpU3ZB1Iz24NsgOpxXV/kLCJKuDRow
DlObkP2nCV24/NHkMUmoH3Ln0HaDAnoH46pvXwp6QANxdpW5/w+j4pohliFV5UPK
J6o8so9xxvODprXMOYrxhZ7VUdJ4GneSWRm0qPvu/lQhUmGpbZTBKJ1mUUip5lPN
JxSVFbPrYI97cUHB+pADJEhsECrA4xSJpIhnUQ08uG36syXChqiKWJkb5LWYfD44
DPD8c+PBSRvJweT+uo1OhF8WSAJjBTKhCD7bqXIsxDrR/5lO6eiSPVyAe8Fh3z6p
54nGjQ7BWkjZrLnDZeBCxFcnsJvZ3aFgXju0pvcH0OCKbvsVRIvficeiFkLrktFI
kK/Lt+mRo4mMhZ6A6CcABxvUdQcctrNtSymh8uk44TfaEOhu1mtq7r8ZvU4yawKG
cG1nny92k3zx6F0Jgy5t0lFjQZFBosc4jKG99Z5kpnrsVZM/lJ6wa6dEHIFpEJ78
zghs7pU/YkP0I6aB7+d2+em2btCsFPot690L7Zt3E+WeyC8eYeKIQPIIG8d93af7
OZV9FLTGeXkaR+JOAQUU8DaKCaaPSVOnQF/82hoDnE+x5abAUPinJiSNVTF4Me/f
+nm/YiVJXQuahKHT5IUJwlefjSgiiiWK+HoUjomPUOJdz8qHxWuXFdQ2Z9ejrmEI
HJ8VRUxODnsmE4g9ULt4S07jx3fQ2UlUmMxowldGgY2uTADIky3FX4pOlifoNKWw
thx4WiiD27l+fV1M5WZ24SubCBzkBl2imjV15rxSyv9/Htzd5zufSPmrcKhlXoqZ
GQEiL/DdcuwMcWzsZxPU3m2MB0AYfJfEhe1MUhklGbq2ZB1egFseEdalHK599wLW
zo60vs8KMWQQ4LSCAWyP35q3Y9lVQ/QgqewnSDuXA7fzo9xubrQ8OQzxY4fAeB3Z
nnJKW4FQML0zC2iNfc+1Yt/gicivJRhcqPnRXWfVcWs/9iKp2TcZpizO7kpKty1B
xeikvm+mbePbvUT6uVEZo7qTlIZdpCw9ij08joquG+93L8YBmehZDe4tfVCUFpU9
3kA1CxrQUEqgz8AGHsk548wdfsWyHpwKsWfU2HUKYJ8ny1nYQAgACwhqCWdF0Aho
RyRru33nZe4cgcqIpEdFXeqhsSYG8VSRm0DBCxRA/9DfEk/VHOYYstcOeanAAWLF
nONMjlm9VDV010dE53FYAg8tPtCSsdfQEi1vu12fIkM2+VwI0adGngxWTlSXkrmU
fT85/DZkRtLQePJGquKh6v//sKlXsiV4I0SqHKNaOyKhQ9c5u5neU3FX2H82IiN5
Jw2QYDVu29k4nxNoGHWLhBdYGUuivO21NjHjvbn14+c7bBCC70TfZeXne/G3mNMc
hTHBBdLN0At6xnHSRzIRN8M5e33Xc4mudpD9EipBSQatuFFLengppiPAQpXmXPdy
KAL0Rm1n8LisHaonktZbJVxg3dns0FKHBuYMeOsLyn2S2rK3rRjkk5ax1/3xqmYv
JLUcDl/pkOPv0etbu9FkBvGOmmmO5px8c04l2xRgJEmm5vVfXZ8zTzWFaoeQEPwE
mz7TWfAB5rCiguF+rZPvFFh3qFnFP/1Qu22n+TRhZ9BXLqMwTgJYhXi6rOj4BhjN
qGdGeQ3NHBHmUoD8hUk8gcJOpoaU4tQugSj+sIv7D0z81vz3bgJ7vLpZVq8lXek8
zIcGRDUJG5xb/PPhiYOZIKkrs2oITDWhdWdheYH9ejIu3rpBI+9q9W1QtrbwG1V/
1GThymYAJ6TgUChnxDrjw5fzT/AeS/7rLtEyJiSC6T5wYKSI9Mw+tEXuSSYAU5ID
R7T8s3iuvPTAHChiW1EKUTeNe8x0aidmrXzOXa/lzvl5MkxEPIbyR8sQr8gjdx1U
Q4Al4DVd3WifasT0iwXOI/qryaeAwbWlyVdirlUPeOio4U0gqAsOcZcMLlE//iEO
np5SmaLXP3wpPEKfpnK/PRQbcjvJ0hEMSmrb/lBIwlP0YQh/XQl/FOK4EREc98Ze
/cyCcQpn9LVq0gPfNN3MEdHDuwwfBFniLgvuCusQwlh3tXY1j75JL7b/8VqeR5dD
08dV/H0LbG2XJgm4PiPj8bCM7xHJiEgN8l92gFTrbb+Siqgl/Snk5ExBMtDMsL06
R6R377nQqG2dWCPrU+iKnCMhyCfPVHrG2solNjH1BxAWJXS3olRViQf1FFiwtngN
wSZ5DAOe4jNTrsvEo7blGT3X1ebn3aucg2d8aOVNRDCKv6mUftvlkcl7XJ1RNuAG
WRIl12ocZoAyWx8bxb/SnuoQKkskFNcOUD/J/3qW8J7254fddqq36zTbKVEgZKs4
DhaeoqrUujGR+8QUvh6bvQ++uabu9AjgIoX0/I4kPOy8NLv70hM9LxCyh3SU51JA
PpUj1dRcre31QKsjcy01LdW22Y2l+8NUdpnCWLFsgT+WTo/JgWY4ZWvwcCKodpKT
bxRXsMku30tXmKtyTYDhX70ilGVFqDHfoIKDgxb5hvS91AcIEnODrjTmbfSuStxA
SEbxsh+uzVaCy85GDR7XKByf+0Lq25pimWTzeCIb2/xSzesGOxf3zzCbPnkU92ET
PYK3yfz7JOPOW7J2mmY64IHmM0R9r1OxW5lFchUhYZcyIKH2nyGIU8+9xFHONfdf
VrFE+TQYTWxBaIXUTEcQ+K9VV0JwgB60SxAMubbEVHBsCYdfW9zOMlIffdR7i+kL
/QynoPRbS3sG+ZZ+qDNYN5zzIq6z5WeIZAds9oCMiDl5gwkrwbn8zm4fvHpAAsX/
TQcW1g2JdhS+X0xLgVF7zKFu79Di7049DMf8SbXQS84s2bsoETodmxW1IJg21Wx5
+L4MTz6NWOUP85+xbrJOkwRLfiQv/f/VxLTg5AtZTlUK2LOAaow1Pdf1SF5zcJcP
j02lFPBRLCl6Iqy4rbmTF12vOkW8qKqBeK7AkZLRPZ07EPC13FM2dqeoGxgjB6OH
y7ln6F5QfYURS8sdtax1t4ttcpTHUiQnkd7kPbtO5+7tnQxlyleY+fMFooG3TtJz
gM+/4Xo8P2sbxcce0OUh4V+oC8xNjA8yED0EJ6UUjjgwi8SqGfGcQUyMmlhB1I45
sqnw6BvPoXiwmCqe96hv8VtUZBtlEjFEZ7AIcZCpAzrdqvVLsEPxWkoGFsxjPRrn
BtCiMf2wDl1mIRQZQ3YbIHDHIM0Bq7LIHfXegfVpGe6McIQnlGtCYiM9OKXVD1O5
AvxEpaenWSCvpWRpLFir9kd5/p9FZLVrjEOquU/vJi/Sx5sPlZWDbGTj7xC4Asr2
IGxXzji6Iy3YWo+Vjx+nTXQftGUhj4U6qCGbI8C3iRscIWJ1f52bDMXQ0mXJQhZ3
D7/HCTDWYLmicRQMjWyDb/lY7nomZ5TEsEJ+uRBIZGUk0VPNr4aHDMMTxezTr+vW
uQ7egzKdE2HmZtYn2fwHjXlx1+QLJF2mIEH5BLbqbYN/9uiCA2gKx9FpWR/C7YIp
miI7OxVFQs1GtMgr8N3qCdrMVZruvlZ3vlSuLVU2ovr/myOO+zvxnv4bIfnY0Wwu
XpXRKSWne4b5WAFFmVmyddLEcaromJhEo0KQJSZRSUhDoBECNF0e8+6cROMQ//vJ
bwPNLWCs16AnI1EiBcAldeBYvM3dzj1yXs6DcxsPUXtVvaVtlCuO2j5jE5/wJ8B6
xZ1CrRaIE5reneJZ6OPsmQ1f7KnPOHPj/iUDTrRjlAcD7Zn0T2p37e3NfwJI4+ck
GZkP4IR9HHyKNJ7jPcBNFAoClqL8achjpeNbrmK/03MGGnhx8oWdzTtw4j8+AmuU
BNO6UMU7m+pQaO88R/345k02m/O/DVWAxc9JQUcdt6+sRwFM0gkBNDfAzBiqIsMn
ssEWtdrDWOnCtQfuCfbk7lcYTZS6V/AiQf6rZEY8OQa0dbd0y8nlGfLHGAsZ67XU
rLiyeitoZ5r2aDn8epLo5QlW2viiU+o7KKiGwwlsm0mlslHaWDqajE0wrEHJtAit
mvLTubrxyKS2MRE2wxeq4g29+qDaR2eJXKRQp8VAA9G9yJ/JA/A8v3PR/mydDaC7
snrDWO8LNHiEaW3YEsk+FdLGatAa+clghMzdNnzMl/XCC+uIR177N2bRjq+jgnXj
63jvP7hQy+m6OavJe61n8Fc3xPFKXe+QotOcmWab85GBf3k7QPYgBEpYwOzpAd36
57mYkcOPNLEg+bpWaZHeDiQBrDDjHXpcSKbUqt4eYta4OL4nJApcMiWgeozbvqdN
NzXRDMFEN3WXDGnwur6uJDZk4ZoSWPRZZnnN7RtwaajTWKdlG+aHc3IJ2dk3NoZs
nTTGbSAdII5lWmdEptJm3qwSi+WzaFfAPX0AUNTUrZbuDwlVUPZScyAW1WcjMcLj
i0/MMTA0s0VQy8UO7b+QmFmvuCvOtab1rzEGZSDDzdeXMH1fhpZH59BBitoa+0uX
eA99OiIrvFAdN1mmx6yXrfQJ6AJVtkwBcwXqhyh86NMwl2b76KH70CIeH0GJGNxt
P3xM6dXkbZhDwVZsQHynwfPA514/DS4bgsIti62QU0isAbdBwmQC/3RCLoDO2FJN
BHvxTBsu1T+pt4KsH97cgcac3zAFnXziynO2aoF1OpGp14GT+yKVCcRwGWeW/lKW
3Muf7SWu4tgJKN1LsDkXrdkk6geNCzWzSu1iuTo1C2gvrNbEqhR9pH8cNfB0frLS
67FnXmPcF97btGgkCQkg4Bnq3I2MYeGnEIx/K1NaPzM9iJajbe/A6xkuS97diGv4
jad/fdPk1zt/fcZr3vT/UQVPQTRTguxUC+pg3jvuNPXgEbQBJJS/YOreHM03ljQ7
5nLWHwMyW2hri/MuXcYjN2ARMD6G5Uxoa6dJ2QdP0+bltzpcIH8g5YCXnmweqHiW
M/haA+HcXFj5AufMt/TGW/n/wd27GitU0kQWV+JLacw63G757mI/LmYbvMLoHddP
yxpWJnjhLsbh4SeXEGH8UBWROnv24ZgphZcUb9IU3Cfel3mR5CulRnfzqQ9u3+lu
QEI21dWPGXTzJ35/tV8oJ0BaShOeEbqrUHBtg1b2N+66aw2XkHhiD0wXgQYp9Mup
Qvazi8wWTogInyw7E48AJvz8pxM+VtdJ7CcOIf72d8F3bZTl0cziiw9rduhZBl5r
AKMdLxhCykieM6ttYtLaOl96POwdDB+T96uUSHj6kiRFu6W9xibxoUeB08r6fkvw
n8+v8J23LXJ/H3h17BRjvdVJHrlHdBx2zUwWpfYd/G0hKnTkLL0bbH5lBUcI6YFa
ze3EKrKAl+ZBziDAiQn8t79mggDSAxenDWn2wBgcdt/7Netf5/7sCDpQCBCR9ydv
QwcGyS2jP0c8M5dv2Wui9KjjaS6a4vr3FH7ZsggZrtTGk4lafq3AkT4tTfnJI2s7
WYBKbm6DJ4zvwyh6gGWiMJqYsW5P1FN0jY5dHAY5PyVKLXduRhlcZ5HrQt0Pia9p
Si3EKAqFhIowZ0PZm3NnVyqxJzVIu0AuFls1i2hGv4TaySB/yA+4l5qur98faE+c
pqsEI5IRqOQ1HmlrYC4N4/rbojJg2RpEKftwQpLPurN80PECj+51Z0O/Fsb7lRQX
8WY0kjgirNdrTcYlGtcDfGcsEQbsFg0MlAbs4ScEjszduNTVp3j51gomSX8xa5GG
kDgf1WlcosWmI7oPnmfK8ZF2ui/Pi3lv5MOe8rTZnkEUHcnwiUie0MVzkU6AZEG/
HMCbe7Tt8AnWPy5iqceavUsr0ZuCZvyZ0Hti6gGvqA6PzGg2JKDzxv/am+nnWeS7
x/gGkIlDdOfyBm5kSXK2Kd9stubK9/PTjcYO2NsLO/l9y4+MqCFenwWeOKOEGnuN
ogj7rrDD0b9Fu+O7USKNcqhDrhYJaeh21VQOm6LPHdJV2t8El7qbCZuGspmikIQa
CzhIvMKvdhAASRk0YpWwhZ06FIMTJJHWMddWilWqhdjHdtZMlXCcxjMmILN7+0Q+
XFPnLoPGNU+h111exF7wnqj6nhHBJXs/qrTyJ3zgjIn/KKDfYhPURrOOmh4lyBBP
tFJLBSlCBzSlxQQtD7c+oxs4HcOXjihR8G86gg8W2uF9CqwEtoS5MMfhkdItZXIZ
Aj42wv7MMdDx51K+fxoH/5jE5fH/LIPQFq/vTnL50Y2BSVn/5y4pLItLhqt4ygDF
bvnoJ6cPkKt8bjxBijC38UjdAzVlLfKCjylX2rEap5DJYl+dAiLoO84maEqWN+eS
067nz/IbsGt8sMqHINrnXmYM1Rlq/MbEHt0pL3nCGnfjnhyoQlCCLKoscs+Em65g
2Vk6XjWdlnvDEzRCzsWuJRAFA/2mKO99+cXcM3M1hRgV3c4tq5vStWMv7DUDvXqj
m7BrXNa3XK5eeW4KBP4MqzX7DAGg8DqJNMYHYLNqKXAtH+kJv8LEi8i5BOiPZSCZ
uK8sutOBNWVwD3xLz32vNkwgBJPHYOGMNWbeKFRNvnnbs56xyu9KJVDnP0jnlQaM
PDCqjx5OlRM57lgcxRU5dS8FdTDxoADophpJR2Es1IqbAkj1rQrr7nHnCKA0axm0
VoCUVpRNoVyXXue/kbf6hWA0JtYi6eOn5l33VFHFklful+2sFuit4SRqXZ5cW8G6
Jx0ueX+P1reX6ZAMzN/jDuwgcbjrEVpOqcT4jVChyvnG6ZYV/0BmhdPEdHjnIQCW
wUhzG5OENJNOTh8gQnyY/S3PNue/CeqU0dGzTAXBShu6rB7TkEWlMwKYS14Z0wdx
E+nFNlv3JWOzcqQEv47Ntu1UkiDVfNqs0CMAOym5U2TdN64qEJzvDXzScQj0HXCV
BCYakWU/I5btsOoyv+rjE7/LXwT5T3aL/HAm0FA38xOwoIEqRJ9P1rmzENo43h50
BDRE0uAEsgD+sjRp14Deqg/rpF/waUhh41GnS8A9IqCORhfG2hpTToJ1qr+S8g4q
2aYYci1dE2rQIakxn7i8CdhPERgtDXhI98hktEXdH9AlW0wTkAxdGMxdpb1xwDJW
yXzyImcBGNAPO1//IB2zl0Q7rn8erHHRc4Mgvsa/KgqvIvkNciEup9cif4qoxZup
XFC7iEurre0bD7voQvYXRjCLuvT+P/r/5G42Q4L5FCNYshRgUSdopUbp0irDaiuQ
IO3HaOWYnPfSDw7Cz5RsjfY7wHlZez/Xf5EVO1z9tDpDleUrBqeqI5x+c+agFptO
CUUiGjKcma+kI3qV/a2/lPkYqejz98uqwoqNAnM6oXZhfvOz6nuioZbvHj6HRf1E
5W230BknPA1dj/SSO1MZoG3RZbVjJ2LVZf9O4mDG/SSrg9e4Bda1iYDgh9WKCb0u
RRaPM+GRAF+sVf0mzNacc6IsKjxhZU8c89YENgtp0H9ECIo3NActtgNlt2zKqMg9
US7t/wgVQ4vaWFfyzQcohfOciSSPEb+IuCWfz8g7F/J5UdBIQp83YnKwPCvpGEAF
cwJtxaLf0jphoap8kQvtva87Uph+7LLGUk6ZsVVx7wAx4rn8V2JffGdmyAI/ReZ1
pBM1lJIomxD+RyPdtmxWjy/x2AGcBP53jmZPGozQz3HTCkOngMn1OMdu+SOaZimo
6VD3P5gctu9AIF7ZavVchqGrHh8p/HZ8XWnfiZjRHM/9laYwI7e0YdFdBZDgQQeS
jRza4zuGMro2LnyWysL7hmu/w4Hu27ArTYBTcyAzGksKW3iX9sGLnexCgqKI1IRU
/JMO1ijTBitlFEHs28WOgk/ikUTJ459WOTxXFgenfzxxnU1wBC3IRyKaO/0hWXmG
VqHKJyoEBiwGqFKcqC50jC3qbXDLll72mmYCdCAO+RbxIv3x8nk7UL5Vd7wlpY+u
nybwKyJl/oA7C7aIc4NxuDjEC9dPJ7MY7NtVkzjOGmQEtlf1H1bXoNauMbnljuhf
Grk1KMjMw80j2KwLVALNr39uSCuv/ykusMFYQVG1PYhoCthd1UncstRAXGG/d5pl
rPxWOXa2zgPrU1P4t0FKndg+gC1azocIbql0Y6NRg8v9W5zxrOu2B6uV6sJIIFw5
VJ0t88axvrg0LSW8aKT/BmHYN4G+hOW7Jpfay27qsVSovtF02qqgdFzJUYaE972S
itjWrT4S7B62+Zc/UaJwgtFZhtnOj3/rtZ6wVa2DmvP7l6Y24IiTe0MnSkP0DpMi
FpPfLbZt6RuQaX4xdliaTZIUDLGLnIeYvfd/BDX+OyStXmHQ4h0rNAholE67RKY0
QZC30nUEFV1Cuk80n+4MseYFKKxihtLp8T5S+q7yScgVFg0eodcKnoyZYhcwsYwQ
W5dJqd98+oCzdN3SbYVzgsQoZbsiulusObxtbKTDy+JCeuVgWUe1VKGlm2DxVs9o
72gVmq9ilLsAflQwTvaU0zta4ugIePG9hCFqhWJF+pOTW31CgEXNRiILtKqvjWEL
jf9S1/4Bl5HVKqo4RPiUiy6Tv1OiGUaugH7PMEmlMIvnFV21ebio/BImwP1zt721
7j0cj0FbVcGEgZpsbsZXPXWAAzN5MKZ8qIpCIOOD6W00x7/W3yyW9Vq4p+yZae2s
dfmjrM/676aHrS03E5I+Uy8lgehcp+ETObuilJVjVPr/Bg3gIMSgBIUzSeVP4VUy
sHUvv4uUlY7cANFwGns2O6i8seasQKdq9xcUogOWSq2ZnEpoT7220qSSZb36afnj
Kd1UYi0TtvpEhmQk27xwAAeT9PjkDRHIDEsUYIQmqpaLxIq1mTfcm4ibTm43JRU2
/cX3YMKTYwr7lP+Vr4bOM7dB+3OwnBIY6okT5p8ohv+SmAb6x7gJ+IzEFKpRojZh
hwWX2ZwJABe8uUwEpIXHc3grKzUXYWopf5cco41GdEeR24VcZFQ/oGJGLBJVZfJy
RW6v5THC002mQVyMRun5CkLM9ETF8fGB6MQ35l3IaXNa/aK67x/DxmCMzuLSJfzQ
bAm5YvIr8sAKr0vvVu3MoRyBFfO9gM/OB4L4yElxsX521+BvWbs03OVR4ZOlEN6Z
cyECjoLZ1ho14GFFxiFzGqP4H4mwIkjSA7eQacMXeS7mXzYRHY11ZT/k17zZ403i
eZy+n6K3uDpWG7vxY0TV62XKKA5DJ7V6JWYOg9LlMVaEB3u4D5hbZjOa9vBf47v3
nwaLj1MvdAKgZH4szdQlM8ZbX/IVTcYpBIvgNcaEuXkOXgkiB7Ju3CHHeppHBD2R
nvlSdERFALFsRZxs8w64APmwmMzjD511000JcH2xrhyjhJ7J9VN/cOUjRMT9N1uY
bOkNwlo2po3PZWPBzhYSYxlhODC1bU6tZOTU/m5knzWQeBLKdDyzS8AOvC9smqi6
LDgWGzUbUlOX58Xnt/UDfupxYadLdp7h1PoI83hPyj6uqKPczqgGUXidVYKDlcdZ
wS+zbQWckjnKvRo0othbEnPqmgU7MloWloNbNFSGvObdpciCDKtujxxQLmpn1E9Q
sCiMAUZquhxqMhQteVsiraUaaTvcW1qWQCuNg4cT2oagN+xvKXtw0BfIISgdHE9Z
kCQBwtiXHXzbV0bhIva16NZHsipGZ1LDcv7TRFmfHxJCkCD0TByQe6FbOBBuVJQF
i2TUTF7woCQ9OfVvjCxYNihIyJk7Y6cmnNYiupcKCc1c9MReENhyAfc1Uiko0an4
YBGAXOe07ihMVIROyox/MI/pYQ8EX2TQtanXClUqPq8YI4ZKC9STmSnZc2y1akok
OWAws/J65ZJwKzX4fqBsktCm16S9xQezSw2eZIDKjSOMUPTx5ddAGip2OdfVJ/4B
laVrXmfUtLR5Hv51gczG3ZF0iTeCMFTSahZLNk2Ry2oFR65gOG5c92KT5GSJbG4E
+//Ydi1JHuzfQhWO4oLKLm35w7o7S6euyEXv0q2C1ZYZSx+ySZoum5V0p1vLpYrG
ZqMKPT3s/Q+XkEIekbe2ms0eTjN1KHPb/2BOP9cKjd3clCBKLgNOYCM13NQy0gN8
JvXMB6S2j/rhIScmsyqKVemFUy+KKuZzSqSL/dwhVAxNwwo2V57Bpl3f9+ckQ+sB
diPZXHFyV8rS4mxGtFZOHBVI1wv53B9vC/t8DYx5riK8/wUsPfcdwcbDQBeq114U
K/IeasuWVID6KeliPz+XEfvDpiLpF3AsRaxfgDRaFaKo3JN3Fip8tcJGPen/W4aK
uCKplx1JBcVNL1xJJ/d6Snn+6K/fu0sx5wJQ1PDX0v0Q0psjOVKefri5wSb+il1P
/s2ZhcG9fQwDQIJDvhdG1QdI3qcjIzfIpfSBEdm1kGUfhLdsBC/2HZIM2ImsCf2+
9ujKVEzGDiRdbXn3+Z5DOXNgpByz7igTOgZEKM5qX6gJthjzcVyaCdmPCg39qDqD
8/ybxRSkJZqI4MIiutXkAUOtvkd+5GRzYmOTlnSW/InLuccB8Xd+rA/Jdk7NJhy0
LM659wybMX/29ct4qc3qzGEWDOFX3YsQjwo7ELtzd2h6Q31NGSkpf34n9E8cHU0c
7zu+dkIin0QMRfbzDHRKZYWbSZ0/7MT7+yXFjW8H2HuhnYAEWnc3d4pBCcng+8Vv
i0cqfoI627Pqpk4IGAmcdawfyJ2RbwdJHvrGrLgvKy5tGVgteOCwvMzNKX+/X+im
2U7oyplwsHy1jpuERPif4f3W6BTRQGj7XAy4ChsweTa8XWCSwr2fFkymGtgrpJ2S
DzgKHGta3kR+RJpp5pUwQmQgkdKbGy+FnTUcu6dSbLXlR/QRPx1a4xbkrZxm19KL
DE/+Xijqdii59tA5pP9ouvNIJAYZY+FH7ULoDwkLLJGW9mTZyIbafHnpbcT8h3Av
eACUTa4HqUtozSpnmGe9eXI8jbwB1741dGMeGzK1n1jF0p8t8qcalD3/ZUxIL7j+
A5vcbgjk1GI2K5MO/44dJQyF7Vb1Y+p1PtYtDeqjE10n3YX4R8s0nQ2qSrRXxsGY
E39rctuhI2Y93TaHT3ISpbUzbAEvUZFrTUtVOiStwH+neiFbYIDJVEwJ9gh1MJJe
MrzOtXYxaMJxAAcAK4k38koTRxbLYiMqQrOIxoycjtGA4MEEjD7t/TDWcaZq8PSW
3KZzFjGvPGmCO25wHcZ2Nkfu5GvS9NL1REoe2t4WiZ1Qf6Pd4+VE12x52oRmjL4O
JwTRtoBZKODbIUUTWaJuGzsBvG+W2N8Az7FGJJCo6NBuCRi9HXSZVLtehmHyMRZ9
3FRbiQia1YUgJvGhqGTNJHu2XZcZckpRhJe8cdxrlTNKBDx0B6nAvfckLV6/F9jV
dDYSdO27feX525vSeWZko7GwzVFplMrtIpTrnzoYd9Y6aejKHAeqVcePFNZeYoP8
d7Gu27ZI1HdXU6O0esVu2rYthKzMk/dW1dpqujKTnTx227+KHga1SHPPc5bryaus
hyEcCFyuRzkASeEZzLHVJXPObZ7HuvvunD3CMkIh+w49zHn2dAfrW/ibhJXxkk+/
W9lm3QkL8J/D9ZdvAsCiCWADRIQqQLy5uvg1AAr8CxvMynuxFIVrflaeptziC2tb
k/7pA2zMg/reQO5Zq027uQBKQC1s42b5Gr8gOADNnm/czMafkARHWH0lW7aMdFUW
5ahPv/VDUGFWH51yAazfeWd79B1D6ZIZxG2EebDQsUU7MHUNDPLWvRFcEoWlikiu
dg5veTdDxt0nFz0rhhaAX5hp15JCLREr6ZnkfynUW2un2NoZakKV51DwwtfofO5i
18QyUJQrKZZAIx4+Fv/2SMoremhq4Lxn1Dq09Uh9hdpx1A6TdH1aXERtF6uM0vgQ
cFEQuyy3ZL6EeAx/Q2sg+gNy4TFsmRz3FYsNQEs4yS4gWfmg58xQ9GLFRdbt5IQZ
Ds6gkSSDIadxKdi3/Y65XR1MQ/fGSPJbSJz/RRYUJQNP8pSOeosDUGmn+PZKgvfF
1I8lLg6yUfo74zhyvBmQWBLWBICNIGQNMHkS3TquamQdR9mneMka7DrUgHcXhKiz
45yZh16xt+aUHF+QY717cVf6xUjyQR0X3vkl7c7aPYn2ijVdmAJjDDtwZFvtoD2n
lK7xvUY/kzVaogHkFTvo+3E+pG6hSOtKvBIGf4hGeIPr4e2tLWkSs3+JDubvww3v
+gvxGGuSB4CYX7+7wY0pUuwarWp0Zdjo/88muRQSvcUTcTH8iJiyOjOJuIXws/gW
eSLYN6HmDeLESyPFexNnNgQ/VJzA6ERrVNNr5VfZosQUq4FhjHlDQxqI1ToIVnE+
VBC2caZxL3RWmv/4a/YUpnGj+ASCAC4igGkI9R09wQcfqALKly477tIjpwtOKvu6
qcDWbgaYwxrKn4CYfkiWeFxx1MaQvez1hraags4DCceNF2QCeBwhq/oFowwmpcxj
voGE3FBDu1VKL0KB3Fi7omW7QtxftN7NkBHY0rvJVHYOzbJewLnkbIlOgXe4uTq8
pQefFTOz7qZiv+UvI1mZTrD5Oku8gGXDvp/8NQ8TQd6Rwd683I9GW887W1t8dnPD
wOEGfVZ2vg1wGFDfDDs3vItmF69wSMJf71F8enOfBuoujHmqB5t4bE2hTKSSpQXp
xVoJ+w+vEiJ9ibmlAlmbASHJ70WRqcveuBHDbzlUWo4UlrM+jqAWyiIykm2nhmqf
qm2MEfwKsA/NA5CNQ/78edJslXAKcyzYEeA/e0IL9cwrfAkRu0YAGvslg0NVnzNz
6lNJgX2WbVfjhHb0q7mb51MRzu+8Uorx/WAp3y0wIqR0WmMPJCKHsI16wwmCiby7
esMY0dqsmcSAJ2Nbs7/Kb7d1UFZ64BJeFdXDEoSvnR+FE0Vgws5wVSE9I6uQIAf1
ZnsZEh8z1opDJhFRNUgnTSYhVk3xncjY324/wDk6uPt1Ec8uYQVIaekeSxGZGmr1
iWt+DF60z/0yFLQq5Ur/HbCQ4FbOuZloaFze7DpZD8j58koAPGoxupM5iArqnSDv
e+M++Xefs/3Tbj8Xg0DoQ3HXTnDzpehe/q8gnhPN2ncP5avxwTQ2051Z59CaQV37
ZFKgIn8hFhO2yWt3hIO61tUCkBorE1x5guk0DmYMkWGRfyR4tHnpKKr2YveJArUL
Aloo2SFMwqjE8E8VM065e4v8jayEORfz22Uq4UuxN2lswzEK9hhQ5cECbZz9B+FN
rSQjC/7UByJYw+ydCIBRDLvWB4sUsTTILhRpfLtnkCQ21wo6cL37QnVkCow9HEcp
YQc0rxQgdJDlMQ1HNohKv6nhfCyJQ+r7wsGTvO3zG6EbpjxNB24w++8aUrrCelap
oD29R6y50/jZvppcdlSuMpur6jTb4CuImpqUKshu4DFpfIrA2CooIBygwEMRdTMC
dWIh6l6l+iO+Z/EOXNt+Pw1MCj1Zvffp5hmdmHo6mpo60aJdspmE5Zfu9O4YL+TL
WosBQBA8QTKNPu24tawsLzU67RaOQyd2cYjAyvZ2VaL7+gCZ4AXlmxq5YS15VOQu
J9XOFQnU8CwUCjMe38h6gNSy02fXU026pnxsyuWDzuIwLRTcAn0ULVt7SS9H3tRR
kYkshLKz034Hz/n47W0CRD9PiAhj0bZ5tytgxkzay5rXs3ZjXQoXYHogsCUKipL+
RKfC1m6MkEQi2qKbQqiNaOnrN2aUiU7XFXiAjP79TzaX4seGKxnHRZNn43DI3WJZ
DGHI31VL/JIi8irBtftsCu320B1nh80SuyyZu8/vUmWkk9MrZwymq6aNXcj4VyWV
RNJ/SxnHHgfQFRAqzckeAdFhd/l1M5uSFYn466aHZdJKt3sHjXOYt/2i0FSlFw+X
CGGtwllgeWR9to0JWo4EhEMbVcOw40w65pD5ibK2DEhpnIfknULOmmHktOa+RGiA
FO+8LzE12A20TH4zX8fsPMia26MF/eX/1TUoboyXUioDbJ+e8Thk0Aa9htOY8m1n
CRS5c6YjluFGpDXb3ZtWN85WvdS5Mo8t8/QeoaOXyyAaojcEdLbTeo2+gUH2CHmh
iHrapIMx4io7l0MeM3E70s3nd6Ll/5QM1dtvSc5b7pc6LCJC1Vb0mUrEenjopsIp
fNJ9suytZi2YMaNeMRHvtSV8EztZnoAdA5NktGPlXEW29e77ff1dT/huO1oVX3yP
PAXSm1kGdiwMmcnBeALHODTwYLap0UUCuICcpn00JZ4lfaK/lmE6YGePBiD1h5z1
3+BeoIJT5aC+3Bu/KeNqPmWTbM3SSNCYXENPz+Avendqv6UaanT4EdTWKQ2jAvjM
T2coFURRjkdtqjMO9yRagIFNGfKIaPCvPadLV61u8Na53M1koJnyjVAdqY9C6CN1
gCK3N9jeXA3uwNIBHWvIiJb796Wj1IP9il7z7YCZdh35M+weZSeOcQZuBOHKihxa
HLWifzQwLfLpfqETnd8LHJajt39398nfetIm3UkHOopmFdenC+e+U9qdIRq8bXvp
T0p88zyiaVJ/a9T9FSr095jiHbiej2rJgA1yB8xhPhCYwWi0+/kFV6/pmInkZCRs
A3+omMcv0Gm2muPUqE9XK/h+r56nk2GaHrduU9grNV5qTtkrmLrvwY5MPl/l86Dy
QrqvEUmNmbHSQ1GpSTZViCKQDvR8dFT7FlyHw2CvZuwvjeZj33gmFYlL0Z9b70TU
Fb5lx+dolRwCj9DoEg13WOeIjNcfbHAHvcaehdWNA98fT7uhtdKjucR3rni8lgNd
mprv7fm4ubBHil9ddON+Qlc981DKpc5QEDHgqp7dzYaytykLriAyylGedWFca/Oc
rz9EIxwrOGYsGDl6b4Fq7B7wUPCcVXxrCa+SBXIozAPqrf7MX/KKabzDEZJodQL2
JwGZ4dwzTq2DD/hERStDtI6r5rCI/QvCTjvuunlvW3r1xzeCbdXLjc7liF9wwyDb
DTx50rIuyvcksO1AakxlTJZfbmm4uFVKe4jJ6dEFZKVe0PAu6ipte+5KNGwz22mP
GaUQyo0+sUzycBE1ZpePwTb4oFzW1KodNCOvO5fb6Z20IG3Nh1kj8Po0ornmmq46
xDQWPQiYPMWgl8z9ifrTGXvrgC9jqq1LUhgTu0lI304qtM4aRMlRJGaaqbPV0c6j
6/vvNxt3QAo7ffoWcQbcdnXHaWXYWOGb8D73xCyw297bBseuauSMvdDpqLCyL6ba
8a0iV6vimOrBVnj5vHSmmZ8SriyePF6GsdTkPkBsYaYbc9K9cd0Wtjk/Hfy3JaPC
3VNLppfMCCmWzisHlS2Ytc4ROnl0xQmtLkY0vHTm7zCHE+Xy0vZSzBWjJQDCZnH1
lI6NU54QQ3jshbXmY5Qiw780eICi0DDvPHoXhXgLy5VDSB6aEUcWTQSxTkMDDolB
ppL46VZHhqTZXVw+aXzBWkJtnirHyjnVk7rIpQeAE1Dcbp8FMpCRkB3irYk+0S5s
2RAzsthBMbaQoqs3nXW3gb/w+M7AUh7hyawOoREDkTO9BrSsrVV8WFHHHn8cJQHj
exzbwkKbFNi4wBnyX6t43mfltn2iZkefeONgSUNuPQzyBMMygxEAZcLahgxdtf6C
bzhrsl5Rt8L7SC84zYd53/+9rw+/LxO2T2lUPyEbBHIG79a3XxO4sEMHz90XhEDK
4uKSHog6nyzkPHA/cqCj1IYxtuRGWCpeuFzumJMUhxqMjRl8bQDzlWym9LA1169v
wwgU5VUcXOPDp+nGGtiycdNVHQwBDwxRdniIjj24UXhGf34hNRf3C3FFoglsXnZ2
VqbuJINOSDPVMu56tWFjlhsxaQCokkWSvwljWbPlZu0OslqBc1jvU0DUesGiFuqt
pA2BI8nGrYim3iDTU/pPDKoQRaon33NLOO1DoSp4ZQnTMY70SJAupBi9vYSszOHO
/HyA1MhlEO+FFCXKtdFn6efQJpHYc0ivvMlHyIs81ZjjiUDNVYtfnLuLXEdm0QD7
yV4wRRJqKrpdPgn1P/yS58je5xwjTJHNuJ7Ztv5evBhtBVul+wW9k9U5Aqt0GGNW
OMEE12b6jVWL9vS4FdG50/09tH8nWKvKUScvpkT607R2dO0fvVjIj+5ZbngxV+8X
W1iPC44/iE4N3BFvR2AytkOBr2O7X5e7L5/mMGVg1NmZLPXlv23Hrq7+/QKBiLI9
m04e38r0zZXvY9XUmlknQSSHEYMrBdArXY6m7T102RJIIMWAce0ZlWpfUSSdTKT0
KxyPv/qF/0zPdh0LwdlcU7Okd/pin1G5lx4/oEdgvt6/p8gXZ7LF1eqRRi7GGRCA
tjU8s2RibyjObJm6TsIdRz0orNj/pBtud5V4V/LhIpryHQLgFbgLv1QEmsaPVRRr
5O/O59wwYlJK35+RUaI0gnJWJDFiTHHdEwP85fE5q9JhCTNukf2YXXDdrlVOZ1AN
vO4ItHe0s3eq1tkcPtf50XR8C2MQ/kgmbb09VGzPga+DuPug/4vLCdTCzBL13Cq/
xR7TKyKkxkEOqmRYXI4kPMe//q5H+mXCAZK5i0vqgMVw7KxBelMe6Ctw+L08JUwv
IjqQkSxHRMx/zM9wkVMFOsyk7mTZC6qTIncDNPYIJGDrlRtbDNa+XB62JDTEI8bS
mxaI5Ww9gIyHwsQntqIXVYfb6afg2JxK024M3BUwjwR1rYbkZTpPf/Zs3gbldGUb
JeSY5L+OycD/H3snNwVAHsYDrzTZUb1veZ3cj21GtdJGe8yh6AgnDYiGdnv422F3
aMTqUi2HTTtPFVZNT0JTHRz67GMg9g/D7Tc1rLaAWbwL+LJchM9DfjngJSK8Vfb1
QcEjmOvWyt0+sz6fG0g3tQAGeqWs11yOUT73hWtmeOU2ZpZbgs+M9GygL2JkUmgi
FH7FUdtIrXumEOWuaIrXFcz8xohuMWYVUeG5gQyLaPkW5E+dPbgsVGMSot/g6G/z
eOYCd9Ed3KJHLjT6Ogd5d25zo6imWyaiqBLRQfIfOO1v/y+XwsusyYay/hvnFRO0
kZMDE5FYJObGMHj6O/ObKy0GODg/onSJIDeHchgyqGz8lN266gpOUW32y7eqLGAo
al0kdWH9klMoHhe6dRzWOfHWdxzqqm+llL4ydzGZX10akr7eyxtA8jXFbQ1Bok8H
AoE3sEPR6588eitw6QYMCD1VO0/1zqgcsaIG95rxtzFybKpEFJK4WoKXWmob0IKK
HJZwrmouj2iC5B+JJCLGulGK9HFybHSr2nDKZ48KZGLYScLcEBh1pnR9aJrWJLma
tIPyCKqY+5Q35fvoNzoXWzmGhhO1lbm2Jaax+MvtQvyu0qrWVdtQZpptx9MGNEP/
4eVR78MDxq0Q/5E/MdNHYdc/ox3eRBKkT5w0/re556mI9Nm4h3aUasZxBtvCRGtO
oUX2gr3FSFiscTTeMw6S7LmhFaph9BQ273zaZotZe1aVb+4+FgKC2SG0z363pvrO
e/Ez4BteWdxlMB1LKAOK3QAi2/HZRFvwQVBLUkZrVXiHwH9Wl3ERlbmKLfC0/DKE
QaQ7vuTdJy/kFpMvbeCR5uqXGN7EdmOSqfqaAuQzGJi55OAfvPss0Z1JXkk6u/ZV
OcniXtEfXEZES9/JRdu2onQwwUS/I5dW6DgAljwVf87Hbtk+UPZvbtXdqlVgWVZA
Fa9K3yTdEkruNIZAHi+8bH9zC//dTUKa0t6O78dq8HfSgXqug6icH+j98i6p7c4z
OYkYh7MbZFd/Ur9czGRMfOnNFj0ytfZkQ5cnbwqqXXOgkIPe5YxPP3ZSQ6fDeTp5
mupY2GetJODsLG9q5ch5Rn/2YMevkg6FMpSuNeBBYv4T+UeNnSVJZKClrmmHhz7S
lUGSkczeUYdyHq1161AP7iHCjjx9dqh2Zxw1kPOORNm0Iie+OpjM66vfiBc2+X4U
Ld4dP30FIWvb14x1Yl6z+Xt64cyiJeeUHrPPdiNYQx1yQRSEtLpNTaGnnFws8KVb
3Eh+XMo+geqvJNe+T9xH8u0XzaLbS39HGXKK56njIyX51YsBAkeNp5Yz5MPvgdOA
HSKCBmkfTugTqo/UlSZaNcANZxj5HfUN2zL74XZWOpIBURF8xreaZQ2Q4agRLc+4
66mb6jpI1CEGayugBZPMcMEkgBjpvzvgDjbcc+KxgjiKc6lQVLcDK7VrXIvibUbM
w1ATLF0rSr4/iabfHgELNp2F4u5mI6XY099mIxmyX06S3MXkRLOkOhnCyTfNVR75
SQvu1Djiq4E15xGYEIA4wkmVEE6XFtk5u+lCGm+nQnp0lTMIV2iRkXOo8diiHLuZ
tbYEvcffsv8wYu2gujJg85mSz6OAZzmtIRbrs38HbEhCSjMgCsgkuwILgnXDAf+i
bnRJYv7gyM2ybWekTokJHaljAu7d6E5Gkm/LSWZjrVUm4oJA4Sjjl5RaKTvU9bgl
YV28utMyidSvltzqxkLV7UwrxwMxxYXPpeTDnLulfTbeb4iPFqJ9s+Zk6EePDcMe
3m7dV740ksKlw/tbQC3B+c1xW/MS1iPxxVghaRIOZcSLKxZG3AxX4YJE/QzUo6cc
fzgYkA+2nrofZzo4jt1Ookm2gXmv8z5fbtQSoW4It+h2QxkxYwWziMMwAIiZ0SnF
cRAWHpPZOUd2/gXw1EoyIIS/KjGMqj2e7zRPFnUzAB3GJKSkA/wwIWEDWCvl+e3v
xH/4OKR3igDp1yqrcG6kZVsz0WXEilJVr/S8bmoZcrwVt+3B2LOwk9n2Ut1WD6fy
hesDgzWa8W3bLW9niZ+WkkR1EGelEHXxEbmyMHqFE2Cf/5QxbbLXQblxIsAPQ/tl
DbxdCbx9DxElcdQEKAXnISkx5evsMCjno1lwQviT2mmkYA1ZhCCgAv2PlK+9FIRl
BAWctKxUja2H4Bue1IMQ20/1zUh9ms4TXpVRI/rYy9mfNmkDB5EtLj83z1vpG/ab
8FQ4SnxE7awmFgCHe5X0oK4HCFUe2hWdxFISnrq2Fswow9hw6e/oZhpyy0D11U6l
0Jr5SN0xbKa1/Y1E7GLWuZw3kCJ30UEPWe8b3QTy2hk0ydHDiBplMUzNuqv6iUvk
z3ivb0K0akGE3oHSnAz2GmPUmwdDIWNJ79bc5X6Is/e1YH5TbVEsS/MazhsuXyEd
xf2TY2EFnkw2BHB6mKTMpPO4m8c5FdRoSvfkiAndUm7OWyAhKnR4CWw1FM59wCIu
nO9dD39hy7VRUFPKwJtCPNeUA7AqVfATxuVD+NEmA2C/PsrNWdu9qR74UYnxxxQy
YvbDcGRmH01lpAnG0LtUs/zhmNqIbbGiArK72h7cpYuVPWfIsAOWlFxe+lR8fvip
dzRCkHbu8HEuVzoG+CuttI/B8VqEVX8VHX82rYNLbjZvGf4F6bahl/2sQWMRIAky
OtwqlLFQUs5rJfzxrJkvN1DHrWwAhM/VL4/dAcfIHqkRtalyHL2WOXXrytQw/uNm
xVFwrNPoPjvMNblXGDESjcyS3i1MG7kzq5ufoasyghezF1h6mgmuw+3hYamLb1oN
4GKOMbTvxSyNtoNcUDRmDLLO0oWsgmRjdJJi1pK80XLbMiJjJUpO7LIoOLtkCfuO
O/QSz+qe46fXQAj2OGwWBHSn/FUCszD8vw6NSS0Wr2Vhc6ACpXvhb9TLuBlkw5xc
svnEdWoYt8i/ECNeXgDlfJfbhi7P6Drp6JSa6pbi4JmCC0Z8McXNpoCIkxg6N2wJ
BafDm36hduOvjH/XyM3kuQ77FUS4k2ygP6PdFZXn1t2apHDMyauxMeeeBpjrL1nQ
3oVJU9hkC/wntDySThX1QQH3pXpCvgoYeOKnEci8cVfoFqek0MdopiyzLq02Inpf
7gsStpqF6vXJikbLFHM3iRG7HidxxcxpfdL2kaOZz9vwzvkFJNEPx2Q8LHST3zjs
IxUu/RjebQNSIBlv2lgLu96LTQG/U2GdnyXHfOEd+E38jtw9wVqzKzWPzoGJhOnY
auH65juRNm+bRGRXxJZJYM+nveqnP1tOHDxFf+7QxT/vTKyhRLFClhVXoLJkzeES
0wLA3JJAHR9r6BJ/sNyo8tZ8rHLK7qy46NIc2j3CYOTW1Q9Y4WFYJCZE+ros71sX
5tCZ1BZtuiidgH78ud2PMf0+07lEFaipto0D4W0GcqcQImQKUJrpAjINoTOMe6T7
FH8sq1Rd/8DxXNGA7D+CuolI0p/iy4P1ibdE2BDnKOD3HE2LnCIOnmTBRFer3ICG
Q0a7Bc5rW+VBPsLHwoj1x038F9m+NfpPOMJsBtVJh6pcmFykUJ/9hJwIP9AqSJU2
jckTt6MeBqUz9RC8UbpfWaDk2LOEC0hIeVUQQ6MEynOl39ld8p1SLbvXoApjV5yx
Em0+otP78Z6mrQFdJbCKcwnY4hbdzhFYbH/+sQo1v2oy/4eSgdOUbahLosFnE1cw
2r0k+uBeeD7+IVDZjXNTbYIxOc2bx8kkuTv7FZOG8QVILJN6Wnf4ZAzgLoRRq+xA
F2QFbYytLiCBVZQZGJVNTazq4K7AC4L/7hGHyraQaLSLLnOzcYrXozVMF7yzxUw2
NsqjRXiF8owO2creRUMCRcLlbApEjWObWW4RehMv4XQVnoBhOPtUjv0w13Bsr86R
CXwNFMUmKQSSpy9jXG6t6St8irJYaZR6Y8ZePYm5+WyiV8cxlD4WMclUWryUeQaW
t8p0V3CScSBCKY2cV5DfVaEtT+5lcQEOmeE1LhDb1mulxPojYD76TCzi5bVJDM+X
97H7MifOlP+AP+eArqbIX3Wrh3aAFhaeVPnYtFyA2S/6eOw6mdUkVVvmeq/kXlWP
CZR09UU7Pw0G9VsWlJ0t1aaytJTssplZ5gExfdUnfFJ4VQFOCPF2fYu5agHkTu2K
bt2gSvfqiKsKN1uiZFN2hFwVFII5dANrzOEhudU5lpTU+xSOnVUhqk6k4F8kg6iU
BK4eaUvOHVZ/HbEBNYdm6xgN9LgfcjV2o4UmT1SBzaX4HUpaj9ieWnZTd4rCZO1W
`protect end_protected