`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36704 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
qe1+t0GXQ5YjcbQQEHGgOYi0TZd/WF19sJ1AgVIdFvfBsp+qlYlkup4zsWoPpDIX
D+k8Kbn1b2edmiP8ax5syu38mBndf5dhhPksHIJ9gYwM+O0UPzw0eC8ICjh4Maiy
y7lu9Y4dxogZxU5wlZkrOFLg52Gd6KJ6OfokEJHXWnvccPLr8UWrQb6EwWdVGl5x
zLfht7xGAiL/gm7zqxAUbn5T7tkE0kvMbq9lYCxenBcOyvuNm9lSUGDDu/W5bVNQ
y04Qb8QqiRO3KxKohdR1Q47H+1Rxua9NZRQyCGATnDoMbTR+f85uQXOX/BaDS3cz
TWtfR5OTtpT1yte+DsN0/JQI/qYrEC5/BtjCd9ZXNezseQzHLtelZ4cgSrvrU570
VCuu9mYHBIWef9khVZ3AqNyNLeqxWy8BqlNyI2bpWR5+9WeBpCIGFeR+kSwFIGNv
01CSf+/oW/uNCQKJ5SmGxwE7AR1+mdmt9fePgCO2vr609xV8iRt4oHhlES4KsKNx
tP6+nBeRHTFc4ZJuSvoQ+VlHx8UO3iUvOPvpm8EGGxMcg6DcZMpguX2HFeX45FxC
1lWLpFNXNc4jGgarY5It+htlncAWjTqCkgeylLz+J0d5leuw1QwI3Bfj7sqHHiRO
6LnQjAiA7n1EBIQeq8zsk/ZLVZwszxihSzX8XP7tfVHGWOVTe1FIuHS0Wc0obWDb
nk/oESo3XqdZCPAfEkRUgukoZmE8N48sTNlTq7vifExT6qGqRyvmy86k1F64oNtE
ELl80nUgFcekxTwLMfg5hrMbbLoO5zQztKVWDB+05DS52yQJ1EFDqshyMhuFMO/y
EAOAfmjKjd8RMnwzYwERtyuewVAlPjp0bq4WiGgKwVloQTcabbcc7CgbITvR96Ni
BPt+Y7e3XUFThmzhFsKmWx/HS0uwbdSIttLlX4rGJZpQk5LQ1I16C25Y6gSz2nKD
I5fXIgH+/CihEKVRbkwqx/0y1ABWcTgZyJ/F6yx1nR4XEo6u8fVQ8U7qdCip2XE5
3a7+qQgCA87Rfw7GjT0NS+YiqnPbe8GMmsIkOGKE6x1As6c7pB5ydQkYcLE/NTva
2ww2n1uHqzWsSSZZ7ZeXFVQwn9yn6N79Le9UVcYt9Zx/zOT4TBeI5vpiJp38G0Rw
7+z5wGcABS9OZ7PY3YUpMUhEDI1QsJPT8fLOI8D2UgLwDQTK0kh5pPnf9OULvGTT
U3UkB5F4gXpfjtBdfhomqti5MqZRnS2UTSdgYRINexSRf+RVBzh9ydQLNkM6Vj/e
oKnVuIVgVDfi5gRe9eIeZYdZMhum0iAYRlBIsvMo+61XC7tsiqfbCvzksPSb88xC
+Bvm5lwR9wQOV1Y3ydvAy2pE+XfMA5QaXY7SpJH0ZJQ2ShGNheDQb1cS7+x3Q5S4
Vqe2oVa6/KoftLSTaAPQAuSxikiaaXF5eletUIjHOjNdFAcKLlyn8Z5Jqzxc9tBJ
pGye9HxcuKF/A6eRfXDoCuzmdXlhcJVSq6NMh+nc68SwxJXTM5gyr703qsq0TMSN
8wyLsdAjCVjdh+riIDeC5Sf75BKOqZ6vNVKPJJGej453vEaQnuG2YiUiMKz6UAP5
oO3WRITfTGgpvAWtVBLJvkNnp0+JDHiGtec9KBK0QfTGw5kN7pdvS/UjP+w5rXWO
gZMK2EjijPFUT6Gs4Cc5VhC+42ecK5zcTPoTdNv+g5w9dZrPF3SA7p4G2R5rVruc
ICR9Ulb+S60CVOi4T3yhqtz/RxUnwljPhpiARpJQRSGaGM15hCsZcKkXipxVRC6Y
JuFdNoJzhUhp9QlsS/qJrJaDbawLn2l0qZEGDwQQ0GYmlrFm269gDoPl2j+0L0K7
xLvqKLrp9lbg93Bvr29RlJxNq/uskAblvee+ovDVyLmADRMMvJE05/+S3PQSKiWk
Ov/S6oiImYOAsc0p2/q+a8F0X+uC3DbfBPiv9oCYG7iPTCbLnFzu4BUpJRqSxaSD
j/Cvl08s6wG6uCEkVPpxamVHrfASGWVDGiJZPWA8DS4tk8DsVBVyfIfRJ4xdpEeE
oodvPNYXAUdhGEbDuGrdsg+Z+f+VyKLguNn7rTaPDwzu/dkwPjS6sHUYqOgsomgz
osvAPr3nos334srDhlwmV7vCicpg65/Fjw+7M/1GUKMcXji5MjULZT37/CNtYSib
xyKutQwgPXom8Fjym5ECV13mduMQVy+t/O4UiQ3M7aM4S2cnBQWxtjP2A+tZ7afO
J0DUo5WgOp2iIzIqutXfVZHanOXetWhg2H8K2XkkOa1C78HMvGX2qnk/TZoEgqGW
0Jk2gD5M5FxEQ0ynxqqWQQQcaCEsZ+wH/3AwNJOUlDH0nJ5LI2oW/zrPqFQKr33T
mnbqd1tODbk452rzs04iJ9NOZ7jflvuV3TW2272/yymgt6jKKz4fiRATAdlkJiMd
DTtN+K/cFH2CFtt8kgbsW2tg9dqiEUXrPqDPysyXL9B6ay/lO0qYJWUI0BtWaeOC
3E5rPGr6ynzSi+sx7ru7fL7eKwek/7xx40fKoq5p/2IOJgkVZNMn2z0vk2I7xMd7
+WI98L+K8wU8BY4UsLbW1+oWMB6O6LDnLMS6M6Lm6kPH8k0hxpfOUZnAj3Z/y0Ku
kZmcj5kVklEdYI89cfzjUfRSIZ3c2v1xaCbH8ValWr9cqV0Oc70B6+nto00gLJZt
23faY1aRKoafIqEjKXP5mtksmoqHNcNVB8HSdBFxNRGbdaSvtThDCAEBY9HPu3cz
sifyUMJmH9EdwOGfNuVpVGxSHKUIODMibJ6mHEiKUpVcU4bhkDvIZ7lH3j5TMTFN
bPEX+h4ayNNGVuAxhUXYPcsCW/giyFWQIo1o7rTw46NBKyBdZF0BPVk1UiVOuXP0
X0M7BOz1eFTCAgeBXRevaZP9zGwuRQfciU76nrXBFVcAHjY8g5tZGtPEL3Xiybxn
QoxD8Zq+60nXXdGlsMnsaEtcDIMvId35vou0xW4l/fIPoytRyI1XYoXGEyiwxHxS
MuDw1WfSSxrMI/g3ssBsb8g3G+s8zhOdHFGpcMUstz8dCIMi0XNt56LDbcy/LFRb
fxBb9Mjbplrnafz3l1yCL+7R6hq209zZQ0P+cIc0eGbpHiVKqKAS4+M7g5A+8MUL
g8O5gfG3o7QCTRThEX8hOLEHosySDSP2Ms8Qh1xmmMRUvsSchw85Z9UUKFge6w2J
f6qiQJYs24KUYLdwbEvtaxj5pLLQ+0eUtNs9EsMM/aXGrxX2NvQjfJSKbztgoYvf
6fjnQUC82hTQsqwKoCkbL3WvAD3c/H0/J6K/KzuM6ADKEhSrXuKAGnE+qpRkV/rH
dz0O357NvnSB0FyssCkcio8PpTHRpKaVFSb7Mmu75Dv9wnibrxybY5tkpq9qF+o7
DQphQ6IdQIoEOe1rxVW3O09ST0TWuubQ9ez3engHl56EbUxx7cf9FvkSKL6AOIRA
HEDurgJCICOe2GdJ/EdizJvIHmOf0QJvwda5I7lRKkAuP98hVqLafv6/eVRQXIyK
E8iM07jz8MTDx/xmc8r2N+z6Hfzn3jO/IBcllTjfPdpujSjJ5HrMNiMU+t3VN5P1
K8jMu8x2W4ZnTQDBnLnz/nJehn3gm4IsQPQ4881W3G/komeQRF567TIzAJ6iwUsP
rmH1yevl+TrmTiqG5nHkMA9l3pIKUknxZDufByGICW4PBL+DEFmUdquuIRxLeVXL
MirPsLWt+xHHsdrEb/ZedBf7t5sFfnReudDRN/x6d1qvaL5D75Ydc2YpcYOkeOpE
bKTC6w2trrGH7RBqMLOry6r3Po3YSMJ73/t1btV5S1xsx06wzebygXkv55+qCQhS
4NLkKa/ZUkcT7paDdISoEx7AEG5rQoz/wyvw7XbVQ5M0jSQW8O0HK3bCyT6y6dMv
eSGR+iw0xd0ziS9HoZWQdvv/4I/+Zug8Yli5qQsg435pCJSBqcdJ3uSxHy0lD9dG
xnMA+gi7mI3POt/ATKbcg8nbNdQ+sA0SIFaZ1e3iimPK6y9YmuMDdEi4YB1hvMGT
WJPgrrXzoEAkXAW2vsRgWy58Xr0h740rGtZipKCnef2OzlmxTptiB/7I8H3TV7Sf
69zyFB33Y92BYC4Auy6b6q1nQzj3oDanw2ESnQOZy1gnQs8Y/5lJIL2d8zoOsrO/
tHL7br0IYdQORB5O9w9QwGgm1zkvqHb6/ixggsX7Og9wmNNUuAoAMijRYzpLgaP9
1m0VfallKYc1GymIj38aY6bDhu8nKGJ7W98WUrxsWMVKjj1KBTXA3WgZcDtPrb07
1vjUG16TcNZE2GBWytU2nktmJjfXtgQdEXQF4FjfFtD+4+oIk4xFuF0Usb+PcKa3
hOMr70r1V0J7HTGnphiG00i7W1GtIP6JAO6u34m6KrxxoedFzAw2LD8NRGMZmgBj
rhpX1S6fsf3Ooj0VyrbaZ4OOrtc8jDPdr1kI0aoL+trTR980PUOY1mmfBuNYecgG
OlHCcK+DMh1p2GPa7/WwA/MnQcFTttsSS9PB3cQOcUcr4PMIbX76o1o/y2lnDr6m
k6SUTZgapXPzTkZyyhF4dUDiAuVF+PEUjfNxRGamunHvbl5pswTlqnjF7FTG6ElD
mLTmjZTUJOT6aBUBXqDZg9YvzOpIz8UEZRrPcmw/vcjlPnj3m9VrkR/WNuv50giu
sMYBghH/XJTo15TVCmE2usF8QdoX7mfgeJayXVcb0+Ux7W2zHpGLXxKWIWwCXLp7
nfj8aLsHDOxCwfm0hAr30FcLFexdkEP99glsSFy3Zheh9PBJv4466Tr7GOYmg4i0
OJrWNXsU5Lk72O4IvWuBTbeHoIkwpXXdFoMo8E4c9IlSsM+buidbix5DLBn2ZGMs
1scwdGPpa5zuneJOPq40vxsfENceokCq05jjAKVdWnAG5zEVbzckPn9IKAanlVqW
lq/NwV4gh6hY/cYFczkZRBQi483cDaQlK1x/6qZ19UfZqW1VOQGLYiGnl3aZ3MIb
g+hn2rl+BWkKb4QfSHrsvKpbjaXtiZ5g1rWqLnZ7qICGmD5ImjQ75WytKoIaYQ3E
3X31L9X7AFLsgkfHSIrHvNyLs/9Hh0MW/yZ4DZ+5cp68TypdJYmHgbyrExvY6kU2
zi1FdGcTxnOc66N0bHgmplJusMLnzNOF6CJSEd5list0sM5AYPn/Jgn5Xohh5WNY
R3WGVsfva3qymrchfhcpmZR7+vX8Q9hvApAe/drMEQXa24dpfFZbnCJnmny9yv1p
TVQe9K7LIQJ9x2Uk4q5kfV7nK+4j5+pQ80XUr2zzIiWHvtJjc3ea162TU5/T1Q5S
A2N9qDEMJwjRM5OzKoXGGJdH1cGIAb/7I1yycKXn8Yf39Qq0+u2EdFbBTDmKEY/S
CXz4SUXtnC7V9DbBk/5zJtGqGh7p+ciDe7vjBErXLc80+5pbtsy+me8y0HDBlYor
3dX941YSLxFnW4Q1Jo7ol/yOeaSLykr40Uz6unUZB4pkH5J+kkpCqRVthCRdyj8x
KLcDGxgAEJJmFPApi1ECylfoMumRCELkbkJbRECV/k0kxILOd0G1TZbk/iQfLXM3
bYeJYUneQVW7HKzA1OVDi0dCkD/KrARCYu5HhRWosaEdcxKNgaptcwcvdRPpS+Jf
EUFAWIUtoeQViEpoXuJR+E/HyA2jb5/U7/Nl47Jqrq9MQtmlU7PZ9hKDTR8lj6hd
6OuF2y0KahH09TneNIcXhIFqPo9wBDXNVEijaCGNelYmhED4gLoVXemjwC7XEX+k
isjBBeiVfD+2UzOMgk7QQC92vkPBWJbe0M7kBAfdoaUHnQuOcKwNL9sJ+qeON16R
Qn/cDHgoCp2soS7YoH9UfOq2gbQB2tS1BMrIDbf+3WwpWRRR9v5kA201SYqNphkM
p4g8jXvFNVd+NeaDdlg12nZjS6TjboqdRQ6luFsSYmgBnvBM9XbVoWOSOtI/JBQF
xG3Wb27wsTVzN+Ju+o8pFOYqp3UBD8yA+S7n1Ur9Z6pZDtwWv7hfNyjuN/opAHKA
L4wAUCN5d25BCDq/W65BhUpvvzLYHHkpHEr1XrNGX9mrqgbWXP02+JJSzRn3ESAz
o8Cq7d8ibuQi/7D6oiiLJZVatFGA8K/5231bPoiXSEEGnKqGm96URj3tQNYxOg7x
Etkl47qOB79+WAXUBZBOWNaC1WZBfscVoe4vlDZl59aCHkA9QojkjMcaWeS6g0le
9O6xdDwVBftV9DqdLWtbPH41adGBADWm+UuhnOTT+XISPNf7XnlWi/MmfgSQDq0p
bphP+tLL0nVB0oB5X5sp2KX24wwRXXUlU24k5Zla1jKM/N9hFqPERZQhHc+6yBI7
jdpLqCTnm9+vnLgYIwEB+KHsMYFbBI++I6SyMJSYXZ4C16dH4yzQ6f1bU+rqIDjg
0cWWETud6Rl6qkujWPqfHN6Hn4dMkTSFGxC17c50VkFQXIyZ0FhYu31T4L1xAOn4
pZzP2myFjDGrV60QkogKAbE5TTDXBdGG9xRDYDSzUiN2dT8PfZPcHLth8LDV1bqQ
WPo69maliwRfMKOC00FIPDMi1AUoOBLDmsn+6Ir4mXoNlHhmoRfF4L6ijqW4bOKf
h14R656CAyWu5sbwOe0pV0uupDaq6i/Uqed6bE6d6u9TLZjwoy3ml6V1qtZoWB+l
zFIVQwu2jtjU2IOtXPP/1fawyJ3GZTHBSLS2zPM7oYLFkkMMEOtdcAjVlvo5ykUz
wQd+v+DvMslBN7NleUl41+h8ut24QDgAp5JO4ImXtdklKgc41VMxUBXTygBIf2jV
SwaOQ53Jo5kSuna784XtYj64BeOzP8UcClLcgZoSpAOXt1jpzkqx3qWzEN3lB7R0
doKjI6xC1WLafTkRPiCsteYPm8JK0/SszlHN3hHhko7hHZRz1/l/uS84iFbwvc/e
Mq3AQX+K6G/BEl8GiIXw6ANAt7mNGdy+rnXl5hVA+0+h2aqDxwtSixTyXlIM7/0N
QPlJWSkO4ZWYXVPU6wcDnLipNh8hUxWE0lVPze4dr9GmVLN0i/ru8HiWG2pz1ruu
SQyTPskmucuki3muAz4Qx831r1LJg85RJ/UNVVuZhxHm5nMRUIVnRIcnrGt3zLzC
m/7w5MJaeUCbyPnt28BW5Y2ROge6gqu72p5cNuKM+cxmXnw4/PSYdy7o6jGYU6PD
wtqO5lGs4u752XgMsbBRPFq3WI0L5lcw5VwD2Ov4IvApSMcL03r5HnrIPVHqGEgx
TcLZMKmnrh2EzLir4CfviGp6HqnCi2Z5xLLqDmtEtGOgtInCIQCNu1i7KCuGBG6a
YqTiKDICyco1jAneQEk/LmYNmpxg2XWnbGNHotVeehx0R+XH+OY7ayRZZbgCn6M0
b5AEN1/ZRWClm5O3LJSK5wNqfmvJSycnlDmswbiS/nebumNTNoQTqIHqR6WzrKvS
o2cQdEmXDHE9p/5IcNeYn4Voyu3UiAcqCYSe6QCdxnF0dOWJwcjUIRcIcKjARdNn
R0ydtT/yNXxBwkTazx5Zik33uFlqrv6jeaeOj7a+LXsSUnYX+ji6qK/Grg51d5Rv
Z3ouajMqdD8uK2odAhGP1fnEHrsz9F2dozKY+8ZtXZl9UIGQLPX53EY6or/J1NrS
fkFpdCnsc24LoERJMjCnb6/MGxNy13oUELljJj6ELCoCUxwgESWLL9n6017Ngjz7
AJ8bK8gZJJZEqJvquTzryxJtk5RHgD+y0OQD5rI/qFzEaPcXLGqeJ//y8im5exef
fvI7nrAT+//siaOjiEKhS3w9kz8lXqb74p07NQoABArrdNcAzx1M1L0T5Ndr+2mg
KS29HHC2alG/rAZ7dNqcb4DGFBDM2QzODGZNSsWuaIBiScQ1o4l9SeeMlB5Lhzbj
Oxc+ZQgjN2ZSXF/50XyfHQVmzCBkWS1n70oUmXvnWRlaGWKFPMOyx+J//U01tGCx
LYWMnVppD+ih9AquuijS7MH8SrBD7XTQFzGi0n4chimLlR/JipRNmAv3HWIhZnmR
R0os5fp2HnjSENwEZIVomm/ZNc17eVDli2lmHVlwJx81qf/cXPZrglX/eyB89DuH
P9gAwdaeeMwzSsOLMdtKfc9fjTYSPxZ9BlANZpwW6JbWi+9KmkzYluLlBJ8xDWs3
zKK15HZtaY/RKcw+ukQ+5Z3a5EapcVPWqz9kwAzWPXgyIeWvOKs5haw0gJblorSQ
K5MV5Ay5dk7pElh8L/9OSTFjXTr93jMZN+BfJA4wOGTr3IDA1U/HRnEEB030eBlS
PaZ66oj60zqqVTGidnMIVRiv5TD5eG96CfEd6DlrGohm3/YXFbvO/A6F7u/VrhGL
w/+PRwM+UP+ePQvHus87Cl4ok4oq5siRWs65yQjDlII/x3gTuQoUivmVU0SqpFY2
gxbdYyq1EOIQNDido7T+XQ1a8cjSh8GxobuBCYXaJ23TJiX3VV0PFV/j8/Mn45RF
0b/iTto5CD+Y/ROi111JvIxQH7H6/0+6HYEqVnRjzZF8X+QlQ/IAPHXkim3DRZ1+
Bt+f7r9v7iZPm3sy8J4/jqAt2r3rH4K4cQ0k9gH581+0iNpPNbJ9TuH8H6Z93Ppp
ycdR3A1u+73ZbnszRqTU06LMqzKWx9mdgJhF8f4Epl6afN9/RP9rKcJvnfuQ4RlX
Rf1YFiHAarVL8bN+k5AO6CP5K6fvdgC34xDwfu5xeF3a2ZVjDT/FevbQUFcy1Jd7
SX9j+ffrnuN0ER9KjrNSZroD1RYjlsyWAhXRSqB6AhktjWspAiHGtJkfT0NHvy3b
sO/t9FuRhevzY544nAFYJoH7RFKg/IoqZwMprwVrK1yCuoagq4CVLmqqqjVmiF8B
U5daHn9Yg/hdyduD/bRrSD08tZp3FR46KOb/A2R3JPa1LmLY9UcvZd7woc4iTdKj
gQgSwg4XB4M7BBDwtFhxVqVbZ/zLTWSL4sioVNojWKsfkaGPgGvqanOItCnCuI7n
xi8tmDRBK2mQQn9MrSLrUOxXc9ByJ36bufUVvRrunXZvfVg48geUTxD5uzH8WgD3
8X6nbc2hH5W2g7YoF3R7wmC6HWTQHDlFuSn40a5sr1uEX/oEK1h95tpHygQsOBrO
I/R+W8Qt94MGNM5k745AGPtnnYb3M7TpGXpjEgB0t44Tr1TZh6fb84Zs0QQ2OO2f
7kgOpvyiKwb2lN3StLkupqoTZqYgYMwPapsaUSAXlhopkUfb71g/8Pa2f/gbnYdf
5F4MAk2lIJ6B0xXy3mCjzBmrAJ28KBYkKihrOegre4y22m5nYKHm2OvGhU4WWZo7
vWOhniXDvkRUGw9/XkFLfOWvFT/XIZt3fwWiSLILtYioo5jlcw6H778bjAkm/8uv
VepdHnVFQYnAAQYmZ6VAtfmX50mXEnDDMYnWNqL8sIMEskAQ2JLnOUn98iPiBsqS
LOFyp8UG9dPyHNlNdwSw+5rGaXAQ4+As4aW6a4fHPMtayDpAiZPtUhIVpKBFs96K
vMitYXuhlOEvWvhLo9Hltv+CHtFEnr29+Di/8j+HwIOFF7JtEcYcBq1Vykf6jN8y
EVXGVqhor/WIOBCaFModpV0yL4RUfeOI78SEZWN4QnVkbV+Upp6A10gGtV4RdYZ5
p+5KKDwdRWd8BQj38pMm99JAYAFLnRXPtZ0hN1xafUO77/8lbcgFUg6NagxWoXlK
Gy18GH/S0eh5hwgEgoXIFpkc3S3tyYhXNqVO2+i69oSjOhBJa30K4uaIIQF1fimb
94MfYpKghw7/TCtZISCFs7ZC4Th9HsTrHwBP/ihm7+x7TBomsUFH264SnddTOziE
+IeCl1RjXIIEkdwn3X+I5Lyb5mtLEtw63RnzpPez8cHVLUGE2SwhfxHtZ4EYtlP3
Dc8tf8ikkl3OVF/+RSFi6h6H9N4InC8F5qCljTS3VRfpWaOfR6113Nab36gr5ru9
gUWhrzQKI1hd6K74KddyUdQth8vyb2wbvxGxFM35rSx5peyLsZhm7wPexSmQATtb
ifStAAoLBI7NsBXCWiv0ffvYIM2hFZQgeU5IffZhhG3nk/1B/7b6Yq4uyPb/cKk4
NsHyymL5xA+jlWa4IEQ0QTw7EujCPz3km2kHhhOBfwNp3qoZujdzWSEI8u2J+nOT
NzEjpUCed49X15JHxKQg+upJOu57xcqnUgcBlRcyorzaW7cky3Ld5mPhRzEx3Yc8
OT4aurxx+7cftdUD4goG8P0PujAWsd3CnOmbXT/eC4Y5Qo6+e59bc4A+w07OkNqN
F/xCDH+33yEM4OaivZQ5iV5gEk6TzfKnhOq68eT/FqJLHotQ81WOYqVcknRPSmHJ
bCp5qAJianNcm7AMUG9ubuQ0wgSfJKPSX2AS3e8c15jxCDKTUj8VjVbLDyhaxLp9
OHhgLQ1xYtKXyTlc4BDlvAKl2BFSrDAoJn6lw3Vyoy69DhimrGw6NEUvTcaG0Bc6
N1ycUpRXhkvPD1bESRbgnEIOpNGJx1ePa+0P48G/eRB5CMXQEndO9KfyBsgRF4ei
LFk/3UKQoIBJdVvtvHDlT7E8Axyl+ZZCx64+ZeKDDedPp492QlZwQfDYfA+MxmgF
pwm7I0mUuyQibCmExD4iFUdWst0QYz95MKUurjFX/EB8fkF0seAz4IFa1UL3Lnfr
YZ30k3vYPzxHIvO27YNMogqS8TbXjZv/b19WGWioBM+S1sAlSLWDQJL2zreB5pL+
Y8W7HxdJ/quQXwDK2504CRi8l31Ts4SAoqYfzk7Z/M/G2+XU3lw90PdcwNMzcBL6
z6MeZn7THeCSz5ZlUhHpykeJF2Kp8anbE/Jcb2jio8VU1iRBz5mqi6EF+wL+l4NA
xR3YQxD/CwuKTensstgiAFDKKLMWNvnFuRT2jKJIwZhPQCeiPQQ17BIjVdG0E0X4
maZGecnttErCIAZrqMBmoBZWa8bZHoT2lYopWzNMRy0b7l2hP4LMgTC0CAHUU29b
eG2JRGEy+6qiZdkV+abqwV4+eD7NLqIWRvf5qfyaRr6unIxz7dM9wqwfgyThfhOD
LnrwQCS+dhFeR2bLMSoL6fiDGJLXdpqw6a6GFnErHasyxD9ulffsfOODH0Fau75+
4+exZ/DkkqjweZgqkSLKvaB81ZOeg9AQZFDoznxmpH6Bqw4MJPt43Qryrh96FFM1
mRI30P1XEEjQFy7PUe4P40Gh5CKGrWJJDhu2Oe1IQz8ze53180lTbnpg205MTdGi
j1FWQMHBGoVRRQENFbAJtRS6PiZj7tOzOPGDRVXBFnac8aDi+85SRPIbD5Wm/3p4
vRWzX3e31B5l0FD8DHbf5gD5VCbpopckRJK+pAVEg6Ru8vwqJU6FmwMoupIgCQFQ
fEQKznmo/3v1LirFQA3DxnJfvDScztl0SbwHmx8Jrhv1ieDEYjc79WazTTWcd5qp
wQiV7HrU5yROQI34FD1KK+K+UDOG0jKaAu214aEisbqsoCD/utN9dc7T225evikp
wZsFDmVTSZ3Ntfn/k5AfzpYg7R7pbw+dWV25h38bVKF5uUtecutLHlqZeQZg6zyl
l/rYogodH8tKLHjClIhVaODa8WRRX5cEC/jqOQ/RunGFfGjXQwmbMPlf+pZL4XaA
AKR2LZM01AySpuCUnKbb/CXQ9ghP1zNGLZJ7WrXqHR+blRynI1MRk1Aeu8K18v2Z
/D+quNJHOPt0SpiwvflFJoXf9LfEHpe6n69DxYtbewdmkDHy3dmmf/wVHa4eOzkb
OUKu+vfHJi7oaWV3OWAqEWKIa/ZEX3mmqSK6mamg94WdjIhPNxRZrfT069L8AjX8
Ms2grYuN5wy3GGlWCtVSJzUzLjqCmuJgcfhig2e4ZzJcjIysS1aipZak9UBtRJQN
qHMugFWKL5NtRJ7C4mxgpqG2Z9fC8qPZ73xNV4WmML8csXfeCxQwaQeqzXSWErE0
ARaxbj4vumRnXNi+qgkLm9ElqAZxx7/n7NeUIimJW4Ycd6An76GZGP/w0tuD+3zT
le3XGCIrm/BCCcjudBx46BSuPOLA5nUer3X7WAzwSqX5OXviJr068i9aINGpF/NJ
XwBLF4FUkOXaM9I4SXCjxzVajpI9K8fWnug8rDVQpVzuMER6AYnyXhkMbbB9A1Bl
4AJtGjli+f2hB3AejdDA7Ri9NMjS7pxls4mVfCLfNRni34dJAWWuUsso7TEusj1m
qbrMmh7ccsMvoor4zEZCzf5Z1LhDAuH8Nj1KZz1n9NVQqYjaC5I+OvGfqhqBlew/
B+U5acvNHhK67eoLM543MSZcaPTbtDVRq9etRbdu2+WuOPy/dR9RV0RW5hLrgJmS
7V4Z1BlZFgUOah/gbIDfcu1VGguZG/bEMxZ3J+FCCVB1u6wv7dGz0G4KOkqRdetV
tcJVA/CXGPXcOOZw2VcwH2iPhdVsP6YuDoxsrrA2MGNYFg7zhoDXKAb3z9JuMCAN
mft8KbJvUZBFX5Ut7jf6hEGeKsSevkKtl+NNG+sgcYJMCR/3HlZgpHGlzIok6zfL
C6nk6f/w0t7Zi0q5ZAeY0eDK68WHOcxMO4FZov2JUE1HGk31r/VLqrTa46hhxdIk
3mZbgEubE1jWdm/6WKSkhhObLVmyAgz2qAzSX7X0YHyfP3XpkRYz37qvh0Zhh1Fd
GOILgz17q24NPpQFz2nhINf2bP3KdkC+wYEXAs+WOSR+0ipykW8UbFmAIZrikUa1
WHi/fBrwCGn7i1vCJ+bjuAUL+6DrFfa39mMavgEcIwtPGFO1hu0Th8ech+no+WhC
siXq9bnWpabre0TChGrdgZphusuCnvqY5HIL0AKJoamK0wAmeHkSt107ktaBaPlJ
fzeyBvsjTVwSPrgAoNRNxG0JUk1yGPXRs1YrIBudnlz7yyjNvxImCHq+vpqv18Of
sLcPYB8SfEJnX5rsvuk+8+MLcCOTJ6hSSFyNpSe0ldj08FNQyid+uA9O0AW5GjFo
+u72mw8t/SMFx8BBuj86+zwI9g8eyML3qiIN78W2uI49zfvm/S7Heut4ZgZHSTOg
K0e5+1BXphG46+O67K3X0jN2SNHqC1OXd1SBpWq92P9ptmRZlCKE1zFj4E0hYMSF
7jHN9pC9n/Mc2sRbSNTP6s+ahDBTy7H5zlGq4s1/Xasq37fxZ+cLd0NvNNAMafYQ
VSw9gpyGZib7VULwv9is9/z72FaiBz7Lkkvf/sg9Ku/0gDDfpUmx+Rd8uBS0rZ77
vPAVJ8APQxPppX3e14yndVy2kRvEaDKKIfyfbAiS7pyF9bmtgJdE5tClcjUPKx5d
n8wNIPjVvCu9l9RsM9FHJDb7MDr7qvJhomcqBZRygU0fXiysuzoVLAbeXVFZ5e0I
NS1fOrkUQU8uJbTqMgTSQHZNzg9CQIwbUgR1zyTWNLkRkOAhh/6OeGf736FCELua
dhwkrtUhqUHlp5T8UEyjseF0JJxcoyVsr1mF2BvubtRufNVu6XI4eFyvf349NvtN
YRq93YEe/7ZLJYI7zIZcAoUq8+p7pTFHiHYkqTFsKW6BqOREKpiQCZZrcwYB6Hv+
WmQCoRfbJ7nKya5k4W1UtUBSExkAFkEFZOfRtwLUV+Rtbk9Qu1fNlFgA1VdLoOkQ
g3Ao2Ekf4rLOvsT7lGs6QbPBPcp5iOul3jM9GtZGMmOdT1rZtPL5xkzj6X0uzEmI
o1DE6aYBdnbU20HnZnpCIkqsDvMA/NhuQsRhdjROj4OijsjN5locaLwf2WinJb8c
NJh2ffzTMfD0p2+RbE0O01TeF7V0ekzHWc+gRIo4pV3TOzFcPKCm7FpT9bwXH/KC
3iGUZQNexbJ/fDDKzjiMyBkfnu/09mnmXWhckwKolgqrvJJWkptm95EcEtUjWwKJ
oMMvi5V+fuBHksMh0abCk4LzUpW2wmGtch2aRPDaLUCuHKNx8UksXCie9ibLgg+R
06DloliBUO0pMwu/YcOuiK/dc/XTU4MztEySns68dybN+O9Q0Wwk7BTB5mkEPMUS
CZbPKwKxzOXDzKhTprIXDya6qmX516zXTw525h849o21S/85PWl7OWMN3io+BAFQ
1F4xENOY57q1QAyR/u++/MuDSjLOS+UTahxigkjEmWMyxBvusJc+j+lM0rbDeTpa
LQpUlRvhI+yQ9nLjkHCTik1PtrmA2Y33cJt1dF8/u4+4Bz35+ot9X+VPEocCR1qa
x1z1meihDnXwXMu6PKyszDvwm8OpFacjhmdI7DIWJE22KPicTFDUpJ+CNOODJUCT
FStAo3AtgXlv8bF7gCY2l0fapg+NYI6o1uD8Z+niqSuiEmd/Slnf2ikstOgQFzs4
9IGKztWbZ/EvcDoSirXCLpgnBPNI3/0p6JNTUMXb9PWBjvtpokYMG5umIDp5sOA1
THS90gDVtoB0vH7N5GJRQeDDTN/cQAfcjteSOV5bP6XdMkUhIOkXVvR7C9IZ2LCc
fXmMsoZ+uRWWbhACOkctOrwxiHQymo1H+11kD6O3oy03hhPH45c+rhj+dKMEt3jH
trL5KK4URmxirIHIWceYhklm6YE8o+JtKj2BJ3xZYS3kxMozhLuG0gi5ZC77OoFK
jpDUziISVdfVlwd6pV/U5rtfZBamt1Q2UF20UtWujNab1zEDTml7NThBBhSurO+j
WFY2Ll+5j2SdqNRQZVRTWkevd1qwsA32boHKsrDathV6MurWPal6ISQsMTBnwPh5
kHD36L4G9Xj5QTeQrCw0jBSa+XLVlg6GjvfqCdv/YBw5jWaKLdjaOi0pHCIS5RD6
VFvBXd/EC8MkzHhW2/Df0FtV5GTWDFOXChyxRrdqRaNUNk6IS92yEDedOUzLMRcA
1mHg16fFg+cqV23QgRSo8VGmqj6KCE/KODiZNraeZFUxVjTzc5+Z8jDTqJ74Nlvl
ho81JYPus1wp9RI5fnKuXTD/Ncu1nnuw2AdSSy2Ls9SP7w/SLpwfM6caLWPfpf1f
LbZ8UE2zcikKcS4t5VEyvy9f0aD4xMSdBxIGTjRwGehrDtlWlJ1Fs1lVDxxp+bCv
V4leUqtOFecB3DWv2rjxu0KkXR0QyDomTzX1C8hac54iHMiFcn4iYM/I+qfpgbqw
tzC4BE2BJNFvFVe8dQliYgTiuOzXzyTvtTKDvZM5CjvBEgZueM7dpdPRKWWVinva
Lt4jNkJdxYYDfolFbGQvrNTBI9BG0/DI1JaCikGi3eOuVXPsFMye9L96O+O9EpGO
JLVY/zx2n1e5lYcWM6Gf4P+0nC/qtACUqbgvQl5WN3FN/9d6FgC0gUxk8P6EQIhS
8/6qW6lAKDoWATl4Q/vss/yAPVQmTF1sXI4hVu+0uH/EieOkNf293R3yb1qP6w97
ErqBHbWeBXYSbsK5Z5X6gNi678fRucicVQPixNHTI6xLU789i5Z7RLXC/F+zgwBl
VCN7H87CFpeA8kBoDCz+QYAFVX8U8ictUqw5PWP4zJsKWJgc82LjH0J0EuLA7g/3
R96VRQKgXatTYC9FShp9fDMk7gcXDO3NiXVhhnqlxIC6lSjT+HP07i+xFal2W182
id1luP1nyrX9z3HTEPmYc0uFU1mN36fQ72FEmOla6Hwkj2ntL70RnYeEYfBdvpaV
HYT+KsPuk4iJEEEw+aZObwfUHTxh+F/WhQDWASesCE9Ra72hRA6m+Sr7y2FlO5it
KoTf5W10oqzGh151aBtibovr6GnDJ63OTYAqkH1C6CIeADdFqT5PbvJThVgK4u+S
cDXmi9Hjnzrs25DxJzd+HCjidBmu24LdLik8fZXqjS2VTR67m6sg5WZKttPzvNol
+W/gJz0CNBRt6hoIXKADAW/J7gOwDaH9gByR1/xuiejZXgcQIbefPgzHMvbClK/s
cTiIOpsFhxMFiANtaU8oeW+xMZwAdJptdnSjeZeo8You4O1iR7AHaVcJ06yFMhB1
hUjvgT1fKFNy59Jhr81/U7CF0h8z5CQ77zX7NU+OZz6yasts0PxPjEZSVDaBGMsL
c9Ak1R3OQH3ftln+hRcSNOoDkB15QTpjiPuMCEIMH6ziellxDA+INx3AaGSBd0dz
61g5kKzdPYTfHSGZlfQvJXhv9xMfGD/afnujCMcBcrh8+pHHnrKcm163qEPwrCLc
ThRNKtPEAtWHl/PHWY3erpCFaEty098OL5U2kTtU9PzgSjvgY8Hk9me9XuFgWxiN
usXXHARIpsiQfQx7Wl/fcd7oPsnrWQhp6JAlr1feqLW/2531cEQTCLCUM0qh+oOR
xinDihkrPtHuMnPA83HlvEy3A9SM8KCV3HzBxUnjG2bhSCSQBRP1DPt30a8hZHy7
qMjxS5SeqvHleEe0eQ1txecSU/wpSvSljD8ce0A0Q0CAHQ5/u5V8q0gU19V8RDEf
5aiL4Z6sAg/O0fT/BGTUG/Xd1kvwpOnHCSzTVbgrHOkd19hSEIpuOluh9CuKvXAo
hsQkiS9TYMAzsSwonm+mlUCB7DB3t/KPCEsq3MdmLYTx8MEiR4Hrh/QEnFOnxZsU
odA1CUY7zKJis9iRywACHi66sOX+sroDVRlaKbgRXby+2Z41MLzFQ+xLdOanmSvj
vH93kxtZJQ01DK3RkYNVUduxQY6e9l2nO9eYoeGoSCuNI8yw129wIhN4WG6f0LRZ
PEzKxZPiq+Clvw9aYojKhcJtqCUQUWeSDt3xquXUD+oAbtb8ok8T7+X6BddZV3Yk
rPZ8rT++sudjjScWkJ8aRcFpT+3zE0ZBETCXDVvpk4jtY3eU7AQ3OrF5p1BpilG1
yxKkp1IIwW8ck20WQv7XMEkZdrpdtFRcE2xA95nQbokX6ceIM2FsYpRn180jHeIX
/XrOF4eGcCjiNCapQxNL8dcViV1s6U+5p8kIJkavc9A64INeHtBUVuBogxdw7Wrn
GcgMS9s6P+8aDJ55HtuOFm4U+Q2t2Hba9UhG/bS7f4p4f9IWTQYLeKIuryGE2pT7
AR4mvo6eygjEaxszH668s350PYyd5FwHmg4EoAQrYCA3BOChHXhzCshITsDM+3bx
PTGM6++2pCkYO/ABGwnoxpgHoZfU9NwEcTupLfm9oswhCeZU9C9Ak+2dgztrP156
i0tbhHnK9t+l/Gfonxi8oLTTsE66Fl9+vFIlorDll8FIIH8jwm9O9GSKxcLH8Ewl
a/aQHhouxCiLDarzvQvgzN6CGK/8jzu4IaCw0tchrLa8kAiUN+1lxH6qciNQ6ucD
P2m6BAOMRKfpNiqDBxo+YsuNvI+SWLleRW74l4B/OWvJ7AyTaCGcC4z/lFsCoELg
RrYK3o4eYxk4K+0t2jAJy+z6zNhu5oc0mdBqB/AXzYSuMckzn/JPgsbbvXokzVlv
Oh6nKLNkcuV395Hpbwmnb+NoHfZPu4ndwL+OCOuYG5ftADkG4+FG3DnkKGF++3FH
2EoOvkd+PPzcEgpo2wgiP98VppbAgwzPZakW6dxkCButZyGqRBNBxEkDvxwGEUUL
XPX9kQCd3YtLQzIK1JoUQujAyqLenj5unthysPYLs8FH1jBoIiEv8mwnAAflJDtz
fWyvoZPI4RvuxG54fx+tGwiAKDxMMg/2oFsWVyx3XQvySClzh5VmSPKC5eN8+3b0
L6R9nYOopbwzUPyTkG8w7jcCgRzhsQpaEEAm/ubU4nMniRr/a+anQdC+vHtDZLHf
Wsi3NlgIXY+iUG6dCdk5XDXKiqG2x65BJSUCeyUtO6KazJsuat5dH+PyhGOueFGR
fwdjjGZgQAMQDIEeOuxB89+1t/R218QT70G9LhbZ1BYtgrsVJqqnIkfrW+QBNJaz
hhlnuP6QouFAVnmkCHwbcYi1iEmfLPI9XJy5tNxQHbAsy6ZHIgSOttM6LPI6aiy4
XComRyiX51KGkrpIZhnvMMQv1icxAT4KQ+qr50mjgiOJ8BChpyGhllUMeaSfit3T
NdBH/4c2NxAVV+mnVxEJjQSl83maQbRuLg8YTeDOjshNjIOdITV9HzInbiURFN64
np/UfGY0hE/teeWxBghFl1meui8F6eVr3P7mp9Ry98sX0DG7b3TKLkc1vZLcdjmr
fv1JbR+XKfcMhf1QzbcIgoTDmw7ZV05i5ceMrkiJPmKCxoNpFVlaIoYBaNxlqS6Y
JEgscu7H9p++u45k+gneKFMjY+AlZoU5gDpvYtwYeBck/3jUIKsX/sRm12a3doXI
E1ayRIl6w4cRpgLPYfLkithqwOFW9tMUGwcihKnNG1LYpj8O6F3QubVx4DJt1XkN
dUuhKR+659X0elXhdrChu39ybw2a7Pyy04zh7t2iHmFd9mIpfygdzs68tIX0wS3M
YsaXmm8Imlnx4qsoyVKCAWnlePu8XynIX3EYCNoW5GsC95kLXXHAP4qmXFbAOSrQ
xpj8QXSK8GcVS5CCwJs+SuF4hKlxZg0bY7wgMzuYvVy3lqqviUmVjvJkf0mfM+Wu
RFxJin7bDtUZ42XeLGZpvht+b/VPP0oUeQsrNGLir4JSZ8X/4LV2KEDOIEAUCoL5
2KsJzKBcR1TGBBS+OkYMy8l+qc8RlFrtZc5d9XthaMKfLZfay+qm8OoZJCB5aDvN
vQsJ1r3+RYQtBgI5TjEBl1Fpzq8wlTIBaCy+lG9I+gPLjaQRdfhES1IYUwZ4V1Tk
ew0fIRRAtrc9G2KhwM1H9OjtPQXAChchxiKCh9VD7yV17dxypX9gLzFr/204Wxkn
9wdeJ5YskmFCQo/poB5RRzn3rE5JnmTGfbWO+K2YDLA3tgrvDMWn5WbZ3OayZNCQ
OaGRLbzPnAMRGPm0Pp/IcsfpoEx0Ivo8/Obcf3weRmPHaliVRW5iyqtgz+dUczMD
dOMW8pOr17sCI5O3270zVLX/2gdwl8lrC7IQG3AuvMdzGAfhAA9Blzi8Se/5AtPL
vL0LNAOa1QhIA6M/GF+qpWSEJAyWHn3wwl14wx8kncA81+PYzZL/WN8/+/hN2gRb
y0s1u7jK4R7upNYg2ECAKpivM9z3mJdw2Bs1DT0NZzud5LWnwDu/RR+niBHMCCO6
oWqE5geERuRqk//Awa+/JkxX7XtyR+1u8oNEmG0B+8c1kD0WJLQxieCZKeirLLMe
Sa18F1N2T0tAGcQJFg8zTXJOHGbijvh8u/VgGidnOe6RveeM24c81wRrAmGA9tl3
34NUou9WS4ZHv1h5N7xZAT9/Hei8Md0kHE/7q38GoHd0SbAOv8T0bcclW+Y2FAR1
wMdBoJXy28IWNlpVVre8QWBxoleUgZdzheHfu/9gd7VSxY8DFSWJaOI3+RtsYCMN
Rvo7cRhL+2wz2f6HMfWJZ06uNa0dL2YonIIqDjt1OeCc9bXRPUB7FqCJTfEwwgVj
6WCiOkQ8oTYsdAr/Fd6dpKmUHljHjdv9qTGj8axuobB7SHT6T9PQqhwAsivGMclh
DdcUK/un59imuGrCw+U4IiaEo3E+krLuSVAmW+wFg/EePMEwZC9yhjmeOdM5GodW
y2c9T7z6ahPy0uZ7ySTkg3t12mtmSfW3JoFktmYNiTKX68VtCPLeG+JQ2ihnMc6K
UbJHTPj/MsXqlKOi0smIbPkgpqiCotaTz/sChkRvaB8pJpr2UqCGKvrPF6eyylxI
c9Rcqzb4UJWp6yiNj/oFkj8jMQBaX5LrAmfGY42tJC4tqhj9PB7of3D3/nqYe8ji
am0G+Z6BaqUphOOoci5ZmETMjiUlK3TS7rW+Rd2mxK8rf953xXH4YZWZTYSncFvr
asELBadthnhgtOp/ZVIfVbh92e+OyoPOEw1NLV9DT3qHkVNNrgXSzyOCiwYOQoTY
rCetD7tiSyVh13bIvRmHJH/6BUf8ip6zrTKphXS008j0L74VzFZRLHu++XiOxpEW
MXjphrleOvG53oS5q+yCf5qKO2lJx9kL9dr2Z+3bUI3BGFUqCA1S4qjYj1627Zme
6ITT/2jJ5zCEHrUSqIsIPO44iOQ/KqPFM8ghhjZEEslmkKr/f+vg2GQUrJje+5lR
VPA28OGgqdhhrM8q1FX1NFHsv+ftzdU1cnfFHzy8nrlhphw3BJfVEo2bMo6maVav
JHfF9Bzojz0IvPKcmx+D+5ZbLsMWS5cVLeNREtAdi5LFjGxeScHYqAh4lovozIh+
QvKMJOjiHTXMfTbgG5729oTioivIzdD/Ti3+WXFAA2o7LjXdd0jrvGBrbu/ZrTzk
fhKfAedXdC4KzIJrUaDEAZDeVD9AbR+FduxgCkdQUb9+MZtH2fSCVTZyZrw21pIa
GspDS8Ptj/7DgKiGCSX6IsjbjeoI6ASfmJvgQ2WF8q7B9DG+cF/8yqI3qmrPofrf
MaEVDvGCDCs9xMUBXW2/OhASn6W8QfYgf6U5eNTmbEWOB7qSNeSaO6rBHVwZS/9K
pvdMJfiZewymfGx4TFb6nNXG1EsiP/6aJQPm/001Jiba+6pevZ6ZXe0W7cjBuPNm
M1rek8wMNcusxSJTWyKD/8BR9HWj/3iA7WRhdMFC2S/FVgmIXZedwhAVzyPzqd2U
j3jpH3uOpCeIPTFX7cRYiCzbAMJTeKb64Xv0SsxcUcdXbMH15dT6QDEQHskVdv28
U1Qa4SRnAPM3VQe10R9wZH6+MxaP4iIJ7IxIVfLD4uhGZt6M9Az975dqJRzZ45qJ
yeKmCXjacPhXJvIiEo1tJNo/Aob59zJoLs34p69zOYbxGRkq4SECqkz7Q9houV3F
Vr1zLAljBruNf+XykyjvuAjRJ/c2MFYb97MXURHqn3FcrPP1dysCeX8NTld2oYmj
+eVL3SLFuL6lNWAlDNh6KhW2C887qoru1hrx44PVfZJj9qyN2SWUSVx2MT/N5WY5
GCHRlGJl2TSYVz4fWWbGcPecOMtmyRJ6Iye6/FvzPfKJf1CeLgiyPaN1o5ir32bc
GVawvm8NYJCfNeABrJEG1WwME3y6yG2s2OykuSGq8kWLY7GMGiEB4XQFytqnftnj
2eTWJ6S+hgMaYHSQFd+UW8SgXy+PGnOk0nKvdSm1S/3Lyc0jfqDaEbuOd348HGnD
8NMU2nWpIqOKlNflmIIRQUblXi2bspTNwRAiLjf97IyZd9uv2eXgaD0UuGZsKbBM
ZFLRpsqCHtyCCX8IdzQWBPj37hdi+yzzfoBawla1aDOHK4C1rkOgMpGVWoroD3Mr
xeotlD66JTVwnz5tmCfJhn9erD8PD6wysw1dTwC2UR7M0YGr1U/hYvGEExnynOUG
SgTfd5nyPVXCobSEiOjxp0t2c5YnWhCN/fetc6bPSauUTJ8q2GKCmja5E5ey9VKR
emRIdIwmk1TexSfY92IkxjfDlpyMuoQIsrK6pU5bTJFF1OEIMNzHa9W/fXqx9Ul8
j6e0b4AuFpBkZcdkaCAXJuYhSV9CS7R2pcwHQTwzlgpf898/m3NuEXOMYIM9tlsW
uriLZ3wZGLHZvikQohfzmm2FC0cdhdk0HezsjO1X/AAWVlVtrECMriDuvNmn6x3F
Pp2w6oh+UGZHvcZ7X6Nr4eHAqTxI2Iz2NDIhGmmgsgUFePBb6dt7oSOKVF92B38R
+bp4jHIUKxx2F8G942c1GLwNUYin2cnYm3sUWclBeq6O0PEKnlDLtR0q2k0JxtHd
6bcbg2mcE5gSdc/hvWml9mt9oKcHAFNx4/dTJe5G+hM65qbAwKi2hqj2uSw+ko1v
uuS1AAzjmTBaRRC7e5kz1lU1JAYBK7nqobkrQroYNzPnXQynn4GwVXDcK+yD36ry
XkSLrDU69GrGCMfI7L6b/HQns1AZFpyDgQZv3FA69EyEL224BZ7cDGN6GfO4VwZB
v0syPw4/eSmAjlU6oYeWAOcPALgNCGPlwN6cK0BYpnRLZj27abSAFG3/PPVjuqG6
DDJl4m2Y+CbudZbwEPEPTuYBnRo24uzw4a1dNqjtXIfc7aYx7t8bhdVzC+fMR5gy
V1F99OF6Rg7eKc9thnUIU7lXAUUpkBUAMxn+wZuntU5RXXQv/lsiW8L1DcdlwMwT
Bstf+MBb39FQ4Ncs4QMCtgr8sc2O3yO1XZCV4aiFLF2WlkIXPV5diNUQFwNV2ZrY
iNWKzNnvfW0K1LQZBJFV5SCUE43uHf50Af+OVVE8zts5cAKi4AnL9TgqFAiX9R8b
za7aSF37//5LGUWWQxLC3HK0qN+N9PbtZZLz13KixphpbVnKpkKEQfe3nyNdebpl
kv9eA7QwHQxk9/Wm0dlqbG35XlZA+PHpIGA9pAzGpxv1vCjP59iV5B/iCFO2Ev41
5V5dRYKECWW9i+erl5rYxBpBTK8yIpuOLeGHPena6LalFcA2SEhQo+OqdW7HnMct
X4PqROm0OHdIbufzb8V1tN5CM5iNRjJDu+dBYYklDYpMPc8o5DB62sEmhe02gqLh
LqckDIlq/FvVo2BSIu+HMmN3mXTYNwvPYjKF+7etoqdZ65DG31l1/WlArGri1lA9
CLgoTokzZ23so0li5YyndM0FokP5fDWLgcl6vWQUJIoKh3lh1VUc+zY5Sk2BuGRB
4jwB3UxuxuTBS/bfD6bIio/1SPRBFGYrqlDRtMqWG9z1+VDSw8S0B7iYljhLWoti
gXPI8n/+HKmq2J4rS8SWfe51V9CCnCwEkRVSsJpCtcBvVMDPo2c/VOEqA39PKj+T
Uz+vWxwERoA57L8uHM/Nk39DsI3cY2IVdpIIA8Z0c/rUbfDB6hGN5SW9CET8OTaM
Hs43+bLtD36GMqBczcvEsm3/RLFbV5sxbWFpdnpE6wZ4on0lnMEyUs8AE/PDgAvJ
Be2e91+2OXH1DoLe/pzw0UsOYkLlaXJGnBFVySfnRViOscXz4Grw9VfO+Wspkjm+
P7H3dxCjHRly6MLu1tzws01rpbo8xvgREO8qXFpza+t9S+rg9BJHSKWaTjX3pf+b
nmJKYBIkTTFXBFTGo+0M64zQqIVu0AVIs/X8e3JrVyS8wGNej371SftePR4WqIs+
/l0fReQEr1koI8OGZ44EsmfPcYQXdoLRePu7ljZ+m39JBCqt5bBHhnBpu3fVYuQR
ZvGl3Ue5Qea8REpL/2g7Qdxxqs0wn2LumjjVUfps9CIE8NsWMpulZDbdCJWvgJUR
MsXCk0PBKPnHBUleajU1YQciOvEc28DxWlzuAhHuGfB7JH0mms8P4r2cC68PYMjJ
+VYfsg0Dd8w+CU00sDTa+/4O546diZkW+MScN/M96YWNGs5dEnlFtBooPR5tVxf7
2ANT1T3ZTX29Hpf2WnsXh63Z5h5LCEtFJomfl3APXnlzPOfBaNj4Lp+EssC+EcWa
IYfkvFhOP1GJvIgV7YucRLX1MBMiEMYS8PO13MWF61Bp/Hwz2LuMA0X6l7wzfzZW
CpG998W/Dc14xkuBA2bx5XgUm94gODc7XZLYYNDFOWimahUKZWxRYVfDZ2RyAi1d
JWWvO6XW4gACcfDaFsPQd0gebmfrBBYwGuDsW78VZpcuFdoprkh99LPhaLvg+uHi
U3Cz3cnubnTEFaPOHZMRfBOpQ9bHUrms58cpDAT+vJfVL3rAjdP+GbwaKIEMoejl
6xn941iTe+DUFeG769aXQ4GS5cXMLxWMqxkqdqI309+w0g/R11kIrer5rkcHAxK7
3LrMR+5FzpTVyXPJIozyxvL9qE7UNOJUFGqLVxb7pO90qouWbmdipFHLw05mwpZ5
YgqRf9S/SMONmDVbvbilx3lAXVSIprGvr6PPWotap1cbPz0Lx5YjDqCAkpW+lLNy
9pAkfEwXgzT8pcQGzNsNcNPvULUXyjTA94igJ6oI/c2OjnLKe24/Tm8DitQ2dHAQ
8+q673tXnEDlZ0trLVKYYRSIROo5FUn99Us0IJu549+6LJ9oGn1szJDDeBz0Xt1u
NzTnKtFSRZaUGMsImgC/9GnfobWGEKFheLK9lCR1vewVp7/OHfKX+2mlzVyiPV8l
XpRr4ygUf1S1mKTUA0Qv7+VQa7ueCvE3JoTH0cXthbgzdecT4VXA4YXRP6s4cGFM
jwjY+Y6rAsqda7mgl1JSJtMOsALzAWBgNkO5kdVaoTaPnf/9umW0NM8mh+qFGToy
i3w0eyeiWTgiYsX1nuR2u2uVGFfvJuopktFcr4H+IRDs4GqFHDIfd1HK2IR/pIwi
tk5RT0BHHyww9k4hTqE4UH1tczxqCjNAs2S5Kf7hFjXfmMPBiz7B9HZuxWe+tx2M
vIsxMEXo52aGxnbuVmWMuHZD3E41shW1vuvo+gw4+qnK1RQoAzZTWJCip+DL+NrM
dNy2hxqwXqYvRo3HGLEmKJ/xN2sZ33kzKO0v629JepbGS62QQsmADND/6thIWa3d
kDWdxYAgKd7qe1XwkYKHCPL0+nbe1VY63wtqrny9kbdhy5xoNrVznZoJaHd8Q+76
lhjcXM9MJbegFS9cPG26k5+E3KdAA3aiuTfw2Y38uF/3qWE/txloDM2xopltamso
Rau30fNs2RGsQTW8ZLt75CvIDiIjHaDLV+ZULzhe2thhEsCDXScD6FPEaJnpoUBC
LZmGA3mxmi0OMjKOPUXCXUnun/qqeMug58HTsBkIPkKwsuVy5/cmv4ZlV81bfj3p
a0ZBwO8/XiDZKz3ZtUCyQa3SSw0X7oWkutU5ybkAbDAabPjGEqjmPEgJES9ZmSbL
j88iZbqcr5i+C2rNf4VPJ/Ia+WRF2miQLablWfLuvux9m99IQmleoSAjzRqqdSGr
SWWgt17OwL6IbARzojwFqTunpxVr7oosh7z1t+WCnhCgmpm0XFfH/LjXvwaRvosK
c8lj7gaEMsJtaNEH1rqoP/4Ku5VJLbfOOhCZC/TAlwDqf+dpr9Ne0Q77cSIfke+L
r1riJ9OFwl1D6HgV9c72YaxRqIkYllKszWpI+3XP3Ihb6gWc2QIJuwisw2kJrrPI
I8eaoC9THTeSw3xr06foEVZvXWi/YAFc3iKSTRBua28fTTlPSD0Cox6XMLESjrp0
iZHJSkGuuquBfVXAbr7OUXcEcgFpaQgtwHZvcf1i3/trR4F/HNfSqx8LpkjJwWji
5fZQdGpP4KX9Z9OJvysaTQvQsBD/lJZQ//EQQKnUQ/jMnxsmfeLNKmwoxtnXkz2j
e+ckmILX1Qsww87HzlzAAJgSLkCYqX4bu8ntRLO/Nrj9DOl5AkecKRBU1rX+XUrU
JL0OqqbsV/FguurEfjBqE3XAOnSlWefLWRJildo8GGyDAbAkr21eL5Qo+rZx1GWg
Wb6Bz9R9JJHeURiAHRU9GhYqLDp2zkhP604W68Vb0xKHJADiPLANZI9/74r8UHD6
PX1HRfXjY+XzF0VT2jsPg3+7xWpij/4LqgfAtNZ1iRc8R3U6/HjXp3DTlvxQQOSX
qakbpG5eMYA46KdeRBIrDCO2WiHj2Oq445gDOA51AJ8kP8gZl7fI3KzQwxhFB8HQ
cDjkxo49xEYj54uFM07JN5XOD7CvkLdlGUZL2IrDW9O6KmQBNwJom118eT/QGCfy
Yh/pcGLZWWnRyXJHu08hnBTUkvXU2RbXLglE9hukROHruOAqtN15aLg2NCLvMlte
l0guVqwwbBckoQZ3rD0lZls+EKiQpD6QQYK/iLVu39Cv2miVs+j/4XPq9MDKa8Ht
j0jJ5JO0sewQmuidtcON8wV0aAhTsTqN/J7nu4pd9T896Fm2pwQPo1ETjQLb5wwf
3AOXhvzv2U02rHF/I/gz79MP8GSxCKQUccDIiykf1t/rga8H13i8RQ2mWEjzVM0S
W+6xkAeLkoLyFx3+9R/vSemNMHnSQK0Q2MJwtXi3+F0w4g0hSc4KyMzgz5hcgsdj
6ypcG54a/NlHvon7HlMXilth3WrlXs7MWwjqhE/ofQgpuKSNUQIdQbJOfU2i8eRF
KwE8yhYXXUNkf1CxSaRbM20QqGhX6wDuj4u4NqjczC+lfFbZCr7c5vHmaikoMfTl
7tjK02zhGSmpumN70xgWMa7Tl9R0ac5JnkNW4krL9ZRJ3iAV6fnMsauoYxuFIlLm
ovS2EdL58iJ4bhsaCVfuOgqTowA4/9aw/HaN2zvHh52Sisn0frcYPyVqkZaZ5Ppi
cUF+6qPde8ntf+3d061SBDI+K2MZDwJ3jUWgHUKMsJwsv3YKWvucQyAoCSKk1sJZ
+S4XjYur3ke1av6+WHmtEJ4cu2SSZL2YOI9i7m6Aif8YRtT+2k8lUpx3e9me+Etp
hHMCIM6r0Dy4Ssn1WdOa7JcqnP+opMPDhWEq5S9I40sbRcDWVFJZT0YNpK5AFFxY
trGw2V08YWS173TUEl3hvl+0EzDYwEL0EVu90RqlY+pVvx0SDEX7ZoV2n+v12Lbd
MLrhHu1X9F0TPQjwzcip5AcQGBceXrzJp5vHb5Vuud2IjeFRQc2o4FHKnJfFyhAg
B/n/logtCf7PnbawRv6yjlCzfsvSTljmzs/J2G9K7pPnCiUHO+Nhzo8bauRRgYXQ
vb584aN7kG7s5n5dIA6rNRW5KJZax4rKUyfHIM3hUsC4QhxbYOXCf8HWhFmdUr0q
PRT3y/YUcRbK88lskqFRj/riN5lbdp9KoOhSGUkcyzeW7JNQrvKRi+x72pomRtyZ
aOLeMcYpl63HPLDi7KACnmOUgwsUslutKA9OPNlvhctOp17+10bT7qX70uP//X39
5E0oNdlywooH09o82nv2X4apbwaX4zZjWRlZiQj9SfmKoRg76ZtszoOGldX3HHHq
wFCmNGtuqE5GS01S8FMMLm8vKWOm0KbpVhAxNYBfxFR1eN0JR477NZMPe/0Y+W01
gAGqvp4xxgjCR8zeXRYAgqWm8MMt5dDK/A3YVqW90IzcKe+Mz4D3eSeTaJtL/k5P
C5S9O2zdqz6Tft2NqzJcbtWDL+8YHF0K1KvHYzAqOR2OErEqx4Mqx15ZBMIHP+DV
X2yYXR9IxjnPL2RBADCnEgU5SfI9QcvN/osc9wUyhofngj0JW4+wRc4VxuoV5ipo
8eFngyUD7xVN0ugPDbXmUDpwGbE6HdHQc7Q3fyseA+AOUDUruA3f6MAxgCZjEvb5
SThfVonhC8pTnjB82ELRBFmsNey7NJSxYfk//Ie93fwb9+RnU2uStgMQpK4RPTRu
/d+BQzKEr1DvvLwYpEIB2m1odcVBy3RjZ92hgmROblaXO85EQrJDJSS6Ouiwf5iP
F3UllLy6AIoefWbO8cLV+xz15s8hvRy2Ul5r8Kuu7zzYw3FOAmmFMDY7qjGbRFk+
Xn4ZJqP2vrJjo+niTiXCAJGu7I31WpRkaBJvjjpuuKd3b/XcJ8xH+Xn27AO4Pzp5
DCsdCoIWgzP4Nw4V62CCowbZESRs0Rn9mv5hMFJWUWfR3qu3BcK7Qsj5gRO2w36U
M4/36Dg8ClQ4TJ+f0XxHNbTZDRIH0Kpa9dyQhM1QzPmH3SB0dtYS2u4+AvzY6F8Q
eZQOzweyojnHGsh092Iam6VZhwpH0TI/j58qqR8oZYjJtPGZadsT3o+FH5++s0ZX
kgY9BGznO0x/OBoTMhUy12OGa4Sq1hU9L16PXvFYqy9KlqmYfXl0CxcQt5gaQLSG
vfmzUFL034pPpEgoL6upOO2BTVOaxUgynjvdvu/ivlWs6eFLcfQdmpzz7NUT3zXa
9hqmZwGzzrPRl3h0YB/jplHjMQ3wEeupWXr1vzdT0JthJENPgtzLfILYR1KJYGs/
xFWnijZ4ALvDn7qQ30wcbtONwLwIuU582N+rwQUsitP6cE2FyAaEuW5UurLw4weC
ILZTrWPEnaUsrXawFXGK3Ad0oYBbeENY3hdF5M7KZKRx7uUsZe2FoF7gg5zGBpbD
sKVpfj8jlaPxSP/wb5lSRLg70LJmKiOzp+fn2wclvThjjKH3UAeLp8iJ8SLvVka/
StDs104TQ4dRurb7L9LOrfZ1wUqQB8hDPKOK1AdmldPJOn9cXF1srSdvGBr2/7gZ
z6Tqjhw/YpTuTX0AgKgthMTQ/0RyaJqFnNs8U/x3KNkuTS6YKBDfB/PFDpKGKSGf
2zVlNbjcAUbY509CLhaVTm7nF3ebgQVIJUYA8mGRD6n8qMdSSbu2wucP3Iesux/3
xUOp72AePq9e5lLA9SJCxyuy2bSEoI9Lol/zeEFHijpKGNKTLtYKAaCUE39OVpi7
66g4ByjMxrNRIVQjTvctO8KWwJpWCEJ5+NHgMWDFAcXjaTCgztv+ESmUpMxvyjV0
dEqDPbCL6ST12rUBx9ekqr3HdoZ5oHJehiGR58EM0r79bHaUOTNS71pFmyOyOGJ4
d7oYP2lDmhi8fHhiVge3lLVI/GYoI4bhyccE0ILjx1z+EpYj7CgIh8kWU0a+bARI
0dBkE1Toz3bTazAuNPkSxlYxWECEb5swQ65UGmfn7gj7ltIR57QACE2PouNKZgaA
3egDMqsvhJ5Uxalvcwf9QscAePyfzm2pM3rWLvFrm7qwlI/ydSmnLAiakjMaLVcq
m57Ocw1pAXQmhM6mMUDC6BEZ9GzBRzTr04m8Ec743kfOcDu8YT1DxrhT2NM0nUIZ
HaSe0T88Ts/Vq4JIVNJ1PDPvUf3cHc4Ntlev/g0Wo0WUw6y6f7xTDaOLqcKEip6J
7nMKnBo1BVpEFBWtUd5+EdP/GEeYDiuo5ki7ejeSXuo7cP+zCYDvMwHeUFQNLeyV
2zTz7ccS+ugHw85JojpqtVuNamCCL6iorGrX9PMWGfWdRULjV4BgWVWPbSbv4RlL
f3Jsu+SvpNJSmtOAS4rikw8pLz38qpg82/+N0juIdp2TsGrmqKHO88s3+Cw4iZB7
1SDqPqRXFQmFGicbo1ttpJCpjfI2Qmle00YK/mWJCNS5WSVsZ24/LciMYjyrESmb
bZcQVr62zo1r29tfG+EANG1oO9YLU9XFZKzNLZmiQ+wxwFuDMGHwbt7x++uWEDwt
gaK4DB+RTTskbR4V1mgWdwioMbxiFtA6eKJ3BC68YzXHdZiomwX2HK+kcveRK9ka
fkb6GKGPvr+3tWLQ/hueWJiZd03roS/Fyf9KkqLj8lLE1c7M6LinGRXFR5PEv6Vh
Oq0vxh/Mjq05LU7X8oMI5kxd5bQBeqGU8Bqt3bHaZO7+SmBL7N0nmairLZwWu+yj
yyaBRQYArlUz4BzP6sOBue8OH9mFloHgHdPLaoX/WYjdmNdM11T5h+G5Q4h+QiTW
J1US29A2WfIXESEWBc8EwwUjmViVJvD4npHfZWIAVNXYOTcPA3aq4y+0IT/eI1uY
sgvZI+8QTI8M57ciQUikqPV+Je8w4UgOlQwn6eRR/dP/qTTSl5bdc/tK9U6OqcBW
0Tj4mPufiUsUvQlgSrLR955Wo28WsEjjCe34713xlJJTPgurEbN2CXnOvZXcrfq0
x+O6Yjs05KaKDKMx02g6HcxQn5uZqh9RDLSrufu1m6vfKHj3lOKWvS0o9D0MT3/f
0Z+bfjnZ3WUJuTK4ki29bLkbrxUApFVrkwImCkZ51FBIoRMllx8O5OKDCF096/cH
dtqM0z7dHUcx+kuucDsYeFytWRyMJfq/4E8RrYCItDqYk08kNBXHiMGGZg1ZsGJq
xnXZzAMPFqeXmAY3fJ/wJILeZ4YrbuuveoZKXbUknd3xxJ4HuvySlrpWl1pq2NJO
Xi/U78qTqd9LHJVfhgWvp0hLpys2J1SPIeBKL47s60Q5KsuqosxPLpdosB2jTgBG
bYJUpFKwjybYRCzn+C/zlGmhEmk56xi0Eg25XsJPO5vENRApOkUVw2YgAkWFiYK3
VqbHms1IDqpyD0g6r+MEYlWaQDXtSLekYGtU+WMXK0nwtk30dDx6SgcLJQ1maGUJ
YW9vyshbz0fZtrQD+fbKCgsB5mgjjpSGeHbHM/jUM5TKNiK2tOVEM0Kv896iI4ix
OPSyXTTUgmIRR8EMWVgnQnkYjPs2U+rPEkmsOBuzhqRSKzQmB5F/os8E1GRYhmuY
Mx5BRBjRm2q2eN8tyFpf2w17L84kGXBL8CkEFjvyidhpb7CEdh+2rTBet/YwrHtO
YOzBmw5PkFriCgGvdEq/tr9v8cTiUlEn454zNMzwLoBt7CgjUNainh2ITdQ+AXTs
kVa1Ip34qf/g2fqt/KMyu1s2TFI/QKIqJWrNIMV1VhrgrPfyeBm0b3tgVS+WkN9C
CnWmJz9LNhNh32Od6mFtQPSCWnTZvfYBaUemNX6daQ6K5LtD4wjQBqDfeeFS7Ymu
e/BmcskctPY/IiusKC4TgtuFM41HZFM8N8kw5cz7mzWydqnvmkdH/ex/5ULifJKM
dphhtUnqWB1rEAZ3EO7n6ax5EtDE5Ek95Dg5Ij46O/F+FCpyQeIusQ//0Myba5Fd
V3lPI2lHuP6G0QQcODYdyBnZYF7m2kzbOVUMVyGgmlEw0B3dWE7Svaenx6VPy8p5
5gd9mO0iKhCGVuq6tUPa1YBXutKpQd7VVIdY0fXAhmboa10z06IdhSX4rGW1Dt+K
4TIIxZbJ9i+Akj1q+QJhqYbvDwB4lKsVLsIY/fSB1A6EjTe6DFdXgP8l7r/Tn1H8
yRaVsyokSsqLUx+r96vuUWeuajW86PHCvioGde2WDHAsY3WwGEZXiqjjIQveE3BS
gZk/9BETVu/kL+WAN/3kf39ouHDrIngiSPB3bFKBlxCNyVVeq/9+8XJ6pFkqbfHd
6m1pnfzVW0S9s+qoV72eAvCEYi+tAs7TI7KjczrW0ND84KldNL3JEtK245x68KRQ
r5dZcl1bMNEaEYZbaQXImAHtvqqDX3/7sC1S4+MrUyx6uyvQIiUqKwXhthy2CGhW
gOceUKDM14Fio8FcU1tNWmaRn+r/Qr0X0qrZJU7hBET4t/6cj8xdZR3KYT23fD+K
2I1Mz2INIG/byffY97fSKj7gsNieUKgFAeGOO/TTOIieu7OODDxr98rAyZhnDTr9
Ff5BZG6XmXqxpkDFCUgdQEZwdLev8gPxhfzY4cePB9KXYjvXOU3MEpGowrW5/pRB
OLiv8JjdNdUt10Cb6mhFaUSJUMehYVg6uo9USNA8oVEWLNSGojJsY9Y8gSXkcrFD
wguyQLksbZS0yG5xFCBnNtMsyWujjuwmUvQH5MXdeqTsIItlgdwBPb0Muju4+QtN
B4eKMxuoei1/DunZ+RDlai4fX5eMYrtyDM9UWgw2qUqWqLqlvxZRzlrmw1C2698c
HST/Szu952T6k5+sfUCf4dyvVfDwf27HUGAyiGwJSDU/8OzbjjLiBku56MXd+aCn
SwHoetD8cIgUysEt0XMmqv2xkn8o9Lxkweylvp8FiTW2KMbJNdR/Xflh0o9adElr
DGl0YvVfDo1tZdJfu4DNcf7IEHNePDUqWO86/SX3ajVF+xj2SJgEICuTNXtMpBGm
WFCRGdHdfzeCUaB06F0U5Dbu3lCmib6KQEvzrs/WV63Agh1jVDGU13PP/454PDON
pDdGwMTi5LRsfzniyZDciTzD0lSsDqeA+11bpZEUjrOVpjBUc4DrLpHYtNOKrOsS
Z8+zZ6RpDpkMnnS26IPhHUd1n8iJvL4CplaewSkVy+Yfh2lhXpLnmTtRMNSTpDmj
LTTVXI87ip5VaVsa65ZwX9pKWDRge4mzUt/lc03CpQcHbBPKEBkJom3+7Fx8QNH+
7B8Nn+VKLykVQ4VqL2/axp2PqrZIRVPxIcF8dPmO50cIW32tas2TZvWcrw09kSmT
r9hotB8W0ntTkywFRIHxmND3AvVWVYM71twE4bWUNAFpukkvZmHN78mK6mQbnrbU
tX4QJGSr1OLpnoouT2EHntvEV4a2SclBsrQJj7Jne2/JvKHT9htnw9VERlPfc68h
98dZUYXiNjKq8/Kc/QpSvBVnG9cxg7R7slq0EesG7Rud1LDIviS2PGZDT1GZ5zWi
3z5/00D43ejjcduKSBbBTFmZAcRlUxxQyTOgdKo+Tc601OVqD3Q5rrohm2C+Qfz7
sB+oY4ZFU1MFt4usNW+Tgz0bdSw3fafkTdkNc6JDQDdL7B/P3gvC69XUDRnlpRdV
PlUDY2xwDMZyo2r3Yxckc7CqiMr6DUUpRKbvSVPfM+DD2KQbwqowmB+qlbwpyp5v
5yw6ZonxzU6anDcQ0yhVIp3MG8xzPppCNTxLlQFnKIFFOXTfz8h+5MY4QkZft3Hf
9rVqXZgBlXkL5u5fZU0zK3fgarJwzwldFEpXNqj+dr1JNt7qlD0TEa9z6Cc5B57d
CIgGvZCM9HinKptKn+gF4zsyC3n9xNHZ1k6u7EtVHZTgXAoNjI19f8WY6FpF16x2
GII1Cdu5dderaCIwL18gDVd/vlJVeLJ1SMh+P+c4oBW1hTqCSx1dBHzGnUeM8rNm
n2d1UxbvJR9h40L9M542u7g4ODXlhtmG5KAphVi0aPiGEdPqOuh3Aej70nB9vEOt
mJFls6HRmbfXd7MUWeNGlUH6K6/aeucK6Of8uCw5SVNNCbCQUBye/CGrtt8yOtkF
hpaIV+7cPfzz4E40SV0D59dlLds+m+Uyg2ubuNUe3LSHyCDB/XrCU21Z+DpkJvf9
1MU7koibH9K5OyzhHoAiJT7/qq4vYHN+eW11PJMlA0fFsgYFyp1rfIYsnJbiw4kY
mFgYQkr18KJ2YqilTTc3m5OvZM8nhjgXAeCrxairdxNUaPKISja98CTB0bUbGsO3
AGOWHtV4P5dUt5IpTPnNS69UfmPC3riJHDFCCpv1kyF1ZU5X66rEyZpf1E0TC54y
QSzj+uzJ/niNctwcUjb8ywHFlNHOIDOGGHmIuzW01+sT6IiHQXo0JXck7UGyEPJQ
70ZR1LE9edQ8yHx46qlTAVuhsKFkSkhI6tMVDGZT9SiMdmyzl3oG00cviA1Hkm28
O3cFHPzT/JnLB4unmoQMWfaiIFwZrYG6PTtyfZjGHquRnMd8RJP+Tbch2OnPNftb
6eEMeqW+4Nkx7PmsY1MLv7MhnFIQpEbts8ok67nHNyi05PWaVcYDyZJl++fgXx4B
PPqBUkRfcWRvUDEmZE6TCHyIeTCb1VEEqF3Dq9M4HWvuxaKbMkkZIuUvIjMxW32N
8dAK5iuIZEbTYVuSX+kHiBNlxXrEZ4F1npuUxv/CCyfGtJF+fU+mwOknMjJ0lYuH
fKuqnB2kKyn9+/PzXvjcGRckhnH37lj+CcaKMFBeFNIQwixzd6veEN/IdSMaTpyY
F+683xJW35dbmjoT7qnnWpilMicAEkrxhS4WfuxuHJV+uAun6yTO3+bdpfWZx+VA
KqRHDrx6CJG3vLhlP/x86Qw9D1YzVax+E44X0lgbsYEY49V5mBFoS4gjiS0RtiXx
SgOJ6DIcqJoMrop2mh7fa9Kt8TXvI70weK9WkoMc5W1jB8M3YAShO14T+b9ByAQ7
Ps5Erg3LJ9W+Qn07XqtgUYPpp6d3fPHZpyIrvIZrYOAMroQ6tka85zL6XTjG97Lz
Hromjx8Bi6gvoQaKTRAStIqju7L6mKYjrKoirAZS6DZoC/AnXrtuFQhBb3VqN1iR
XrAOfay5VMsfgiM8bFvMoBXItDeq+snO93nV5ykQu+VZJVb25Fzzaxb4zI+7FZEW
UWXdDM9lJK0yh646DvtjR0h/ythlzARPipgL4phJ4XBVvEoElluIMTyLpXXheRuK
hSx4V+fFmhVYQecxtovlxyDoFjqdUEvRai2xURjdsWfFBuwvt7M5mqk3ODmB46V4
pBL72y3dEx8im/NyHW3iB7GyayFkd5viCTFVo27beIlf/kHw68B6oTc44kLWiqBU
qV+FGO1vkeAOYA2Yydise88GddRKLvfvmyg6k0If1iaqrkPwSBI4GWdt4lPjqfdw
zK+HYS68vDhRatRN40cE2PjfWM82HpUIzb9UjU1UWgOBUxWyxNQ8mXlLtsbvoAo8
d7gA2rxHhPtylQywNwPI60G4cMffn7zbahtqvczxm6DBgyFqNsoNyTghv3VzG+o1
+azRMpWPdvEITXZY/tfPRlwGkxx71eoPjGiSNW+Z3BZ6/qvts9oCs4nd0UER++sN
q3uJ0tjJhyFFF2Q871XPslfZLx7BL7vmJNH2VAbJAqmvRNYmj+FxGwm0O3Wz8qPx
K7H/f944JA+g6lo2qj4UVd4MzGQpoha8SSrf6P0GwyLRz11PwWZWVhO12p1u6SvK
/zaxH7Eu/8w+z84Rqg0h+taWsmTllGzCgL3Mo7f+DSZqH58beODXfpspkLZVeeO1
nmCVCW0VfbY24fzRstUcbeZbNcDWHPRLOAWCvPhvTndh2l/6lMpLEf8bIIJQYTUI
W3W5frvdojHd0kbS57rFbnpOh+Lk7j4voP/EJQ7lzO6fwK6cCR6tTp23nsfkCW08
TAc8zMhfJBcDXDtTkBP+RjnsXXKQXglw7ZJu0NVWSH1LWrY2ayi3NF273H2s1apW
mhpvtOVO1oEjuK6R/AUqaXEr6Gucad0Qp8S1zyfnHGjeS5t7lDsl5dfRmYcanjBY
MnXijHDwQYU8l9PWljewHiH9NTxedeDP5jsGQeZDaljEFy+XlZlh2TGmSq6VERbD
9QLPR87msnM95DYRJ5in53kRMN08HVXUt87CJy+QPr/2+SYbhPVXkUUD3wRMPwMw
mLhWmyMkCVZxxR2VmX0CYsnZA8DbKIa33kpMDg+VNsTN5sk2VtmkWf8YCpdKQ4wO
Gk3W52DgF5EvYqspHmjWplL3HL5No0oo0oXMjC2UDIF+nJ4xyqa9IFEvJFXk4zO0
xDKOJClay87OsH0JEIfK71ef2z87N3Tz3SXbrgl3yDCPYctDC+pIaPjeUQpQ5iPP
r15/t5PM7yZ7xILJrQiE/P98LbbC2VDI5awGkvQFoWwaEjwQNtAaBqE1ad0eu9DN
/+S6k6fKRiOTBLmYko9jMb1G148wBrLqGyMcquw7c0IUg16AyDjLSi7XXKub0Zcq
ONT3nIUda7pG3jUlT1+XqUpRlt1HQfoOz4BwdTGLUwZCBaNFFZijQmaz/clD1PlA
JGJaBKTmf5DMR5tzNmU0js7wdg9zXHjKCYRzTWR4offCgaV6bFVpyT86du4dkHcZ
n9ObaT5ac7m9y+5wJNSs49Sr7kNZMA7ngS9EdnyKPHfqByxg0iwZI1BeFg+3kKJL
JB7AgjvBf3XKgXx1jfmJen+JMfzvymTKIb3SsBq4wo2LNDaz/3A1efR2PC2LoS14
fdJv37qPIsq5RL4mJd+ijcIXSZLBTqgSyA0q4Or0/zTlSbXnX34bKO8f2Cbqdg3l
FJenzL24LF8IQeY80/cdDsxer67j+yysk+BKIxUytTKWjjw9z3dAOYcJCjY4Qucv
Dm16QSJ/gJZWVFZ+slOY0UZJYd1jNXDzhRbqFQ5zujM7k2ICa0KniDFOgs+GOrlq
sxDo2iBDfPCI9oS2Y4JmWD0knVxhMJZ0mJLmr+8buVZx1zQTS1NyD62q9mYnwpPL
by3yKQ5L3S8apea9zNwW0YXjfhYe6Zp5Jbu/qRpnz8S0rMKvD3nC7DObkZVXns98
uwNKszndiiGh4OHvjPxJz3xf+8mxLJc2itsViTDjU+crfdeV9NcoQb6F6jrtDhXd
xk1Vjtm2uLISFGIYilf+xoJbXbNcsi4+K8ilsbGgnqXWpyej2XHORkqkgT2jlleO
DKsdYZewPO4rZ43bUiXdE7oG8rE68csRyrCoGPg9uEmCXMbHNwVKCIPz6xR6nx3U
nRzu1Op1dRW68mkQUnNint+9ca4koMZroGliRgZMvjvlzf2fMvv6vey2ys3wf8H/
XThso0t2VujNGFhvNk/cR3IRXV5TUuTSvFweoOSy9zcGusAmMHToD3jnjSEL23rE
43j9ppw2BSk0TrK3TeBVsbHmkbzv2lX2PGD4EU8VTGNGBi+NmiBTU6T2YeDOFt6d
7veysMJu6xLS7QFCJnKkYColMPQ1rpKkLFaxX8qP6mDb7HmX9m+GLTzBnynHkOVN
WhhlY7f3SP7cW/hSNMb/ZBX9gFBoK9vq3xiqMaAG4gUge04f4WBywat6LhxDJZ3E
wJumRi/hrJxoqmyImB9VQ9Tv2T+b2OkPiUq7cgOq1+7JPlzBbvX25RBhG1oRp7sg
08RamrKJnOm1e5+2anjeI0fwSkoXebQqjboit5yaRhzwirHFauisNBEIB0lK0zU4
K9aNkBlKZxSbMvIs4DfBgxcb2LSfJmKG9l7yfCq3awJ87LytUKRjlfXnn94peV1d
09fw+aRrvJLOLT5F6YjhIMAOpYl1GhWyJzRHBe9Iahl9kzPnJbPAdXEO54kIRzQY
IIX5DyWVbFKABwHUm2TbvvnGimGBidEgO/xFAXY2JTrYgycwTgy+YW7wR7VDdPks
sYjKOZZOPF+oyIYMBZPMBN6CpEd6pn8CyKsfow6IEK7+fDbZNgDrXh4MCBvq1cx2
RbW8VTT869NQblytYnC6CC556OQ+lqdtu7P+dnSlsQQEt1v+Hvz/wHH8MrR+k0h6
3EMWEMirPGN/s8iJ4PzcawHadstpLHbgoOIN9mhs2avfBbfaZCU7j+IOE5i1dKkP
bCaHh0niiMNCqAnUCDl8zDEkSiSlO3XLfWBZnJnpfvBoxAjzAj7QK/ZRCOfJLp7k
S8RfY2exNe7KrGAqoOjbnJhQQge2vtI1BOGpTyha3Q/vBhEbxdFOtY5sWXRP7Xzt
gymNW4hXxoYPfBO/8++VmJ6CcKiX/XDfx3DeXuhyIL29SzFkEQMZnQHeOWCh6Tow
Lu/SesVDuW3gVk23aXVLq4htC/cjhz/MGWmO3RXTzuL7JGYX3vO79MTcAdRft/js
xnGhq7DQuH3qPERWylFl4iVwLqbPKj7vwWAr9vdwJdjouY8HUn/+vX/YZbbOeZrZ
F0BSqrS1SeE49+kxcNDNXEhgE4HzWcJ0odhlZPPHNUuHN3VFGvc0J8nx34WWVswe
0+IlKcp2XfYfop9Ohu74Gk0Sy2IgameEnlMGuT1/+IRpQpf56VC8HD3qaR03AG01
AJZCopOzDIqFe5/Tvgw4bBUsnBPO6pQ85yZtDotyEwCmpCIZrkek55HtUAL1oV7D
6pATnDT22by1fAZPAdKu2V4nMLrmc9g6iAZzTwuuTHJAXIcUKCqnf2z/Of6TbexO
tt2krGUGDczkeQZRC9goBLMmYiUtCQWdeuxzm1JxP8VTpXpcPYvrxE9+n+wxWHYl
/MxpIG0D327dxnurQOQuQWwXWcvZmnv5rSXZ1zldG8lsYfmQWsIdw0YUvbHrRu6C
QQhsm+2OSKYJyBbysHNBAN55tF5nttmazlufRb2Ei/XmzSlHXbAQNh05JTYTIg3y
I8i/AlmQsh6/2cwcUMskswxkuGrYlZzLXZz00pgvGfcFas2ulXAgN86ZEvuY6FsC
l7zuzOymRMrPtPoFDeyJD5ixUGl2cYw62vf6Ggoi0vbxbeLbFDPLHlu2jhCLng0a
2RsACYMVq5bQirgSudWC72+5A9Nst1HYgo1q+DMeS0hzq1PI4Sn/HrknXTXMugHs
KCy5Xg9SMb1pQZulfHjw2bngToSRNvjWqUkCmFtFHgF3QLMw8yW/e7QexxVsMr1f
Ta1mM5LLiDmVTelQOfpy7haskfNqB5R+XUWWduGgGJqS/Fr+LLRleXLoKgwZ5RdA
lPhW1BufmBYtWRvxTzfp7/yh0f83tUeKZPRxeCa/ICT+mJ5t7axVa3xvknfVw4Uf
W9i43Dhpw7Cv2GEqcUAXpj1mS2SRnr7fAFoJ5QEF4jjNRSo3cRIcPEq6SczlF5Fy
YFf1vmLcL0radOnwwejppRshYvq1UenjrVECZo92vUC2X3xlzTLqcbC1F1JiOdUt
LbF3cLWg6ngf0g3lKxNK7hu1IeaZm0eZ9dytJdPFzvLfoO9WD8MJW+NQUiSPYGvS
NaD1axqecsC/EbvF726RbYu48FGNYPiUZpdw5IfpXqj+09Z1pKy5f3F3G90pr13s
uaegjX74ePqISBVLZxwvqKNtXdT9qeGFRgL650TvpTaZ8WZPJyQyqdhp5ON4S7VH
L3hbxyYgQJoVKOJ5U9K76QWSRWks2P6YIUGNmelpYn8UoXJMiU4oSWJyX/wWSXCQ
WH0vKpoKbfoid09gDHpiYZ44FBBF5EOaXwjPz+8PO7iiPsr6qQ6RRQesdXnilklI
OMTqR+KQyz8LSmky2oNk/fhI0CL7GxmdSoL4/i361r/Xim4+2zCIVOul5hsOWXhE
3uiwmQQKcK7xIxsVA55vZZSG3A89dGhQcdDFcQb+Xxrua7UrCDLdudI4RCW6d8TB
/5AnXo73P6Wkg0E9Sa+RxpExyPEa/t8LddmlXETBMVLNNT4dwF+A1CVsM+vEwk1N
eUcJoLtBvACfQnhrRx1DJ+cOJ3S8lYurtYAjbCFm72UDb3Vbs3vIt9+asDC9AVIb
XOvB+AHl2WAy9NNtcF1qvwIJaeNmmpolA7+l4Lc2bTk+y48EViu9QbFRJwQT2q7Q
AEsea3vhBnsCcW9yUHV4oj9Ur/cLg29qlw7EHIzqQhD4txTG9OJVoBxgWJj9S0Y/
8D+Ddjm1DOO40hExH3su5qm6cGwiCsrtqvQSJXOSki4iA5AWGhW7hxHYiRSmQLfP
d8RDYs02jO0Rv/a11t9nvWKDRg/db0479ywceuPcfwqu1o5oqWr784lOvK/xa/Eo
3aCqFya6ZdbJ418sPngx42KPZGi/VI+XWbRssRq2uLb2GVdDEiEoEVNoqTO3N77/
9Mt4uj4rnfG4VIrL1xEiVPkttQuKSOhCZYd83chisPc71H9CWKFEI31ZPaaGxF0x
DuDc5rmTBy+U4phHNkQnWpfXKlQlRMybZQ4ffpwj7PQOUjjpwZ4MCmbnFx3xpnQS
2MzGg6sduPF9c3WJbT9nPKq0v9Z55rsIJ0Kz/qaPVH3jfcJ0yAzZ+/oWJVLN980n
MBG0cQR6SKJBi4EJAfntGd9ccnQjjGnnwd1b78F48gssNwbtyJbysmwnffL7xuKP
egNg6Rt6ekwAc7vlf0MtnnsqRXPRh/Pe/dIBHJ4mLhC6YBkZ+JvQMi1WXRPUO1OW
Kfn+Xk3JkA2/5gc9F13ulOKOEUhSxu5H6qbwlb31XOSjIh7R3F+oYTMx4iMvcgkH
6DzJtfsZ32TboJqrV+++QYo/HKRTfuFbhBDv0bOQTVvCko8EysXIoFt9fMH/i6nT
tPOcKDh06e8wtrgF+X9Z4E/JglGhJZmmQxPy7cRrbKxuC76AyoxPTQIlX30Vh6p1
vylkJxQIxa5QyqmadZxcMnUTbmUiIxniXA8V7gXI2RKpBrsYKnM1xEE+DKYhDjT+
vlFyBCzPbl0WVAWS4zx4uosgyzjpunJqb+yKaS8LQJVkpREENhnKXvx9WjzzYQfM
V6wdw0rUmroug09boDmJcOEYcxpMepNBEtXHRoRPvSZGUrYMIxNM4A9blerARuHm
IcQAiEUE+YoNz/GLlS/TJ392I4jfiJ/vhUVWHWmZRuhpsjGymI7NZ1409SXELrNN
wcCQ+fWR6zoT4I+K/shccF63y+cXonWLZx3A4Zu0U+Cwji2N4yy4sxfey4hXZVH3
8DXqBXWA+S6fsdP6w44hMqGIwfmSRU0K9XmlzS5yBP+BnRafxtyav7hl/0wWFLQh
bbcUcyECm/KuHf+imjg6X+1Gpm9wRRpI0wBGF4jBVi5DprsdhobOFGcmSr6ihmvS
i0Row1qhIGeLb50lI9Vndow9/rrH6dYWdKHjptBCSY39sttkvsia7lUtM1+rLtNH
7Dq8Qt69Mnl+l63EXWEg4f1V3c/+1gErWXWzwawQEaBeIpeXlX1EAQFfExPtocnA
XLEuWQVp/mUywFjuihVGNcPDN+rS9CB44zIOUTrT8/kuqV8Q2sRHrNOcY7TmR4OW
ktQunqgE8Z9ff7ylZ10blj0qOcmAW5Rx81+DgmvmvjPI8RHsnqESrayzEt8yP+Q/
Pto58fnmDGgsircobM4RaEXAsvXP3tRTa9qa+rm91VPgCjrYh0Ok54MyUsctauoQ
cYJldZLORWONuzwPvvil8uXDR4S9QPySWVQqfRiHqC3gskhBYHysyHktg12r2OpN
vBfhFUhh5ipgVIPyz1ZwP7PDxH/1mATbPQMLEdEuL2bN3s99jnKxtKnl3jxNTw5T
msFTZlSSMY3USNpwigGsGCrrU67lIBcuO7xSOtvP5nRslrIlCSfo9ncgH+8cRkcM
ra0k37aJJINH/lwfK7G9TwmqxYMrpd2SG7jW/0UzHeqZIZK2dhPcYv24YRPFFpOL
p2+uqVvc/xKrT2iZVLJl4/MaFHVsp+Fi59hJC2SxGlAJRrxIxmVmhYMgkkZud6eu
i1tW5VjKgRh9IZAOgxNGcn9oFgd5g48TjoNwUmEqD/OoPIpowFb1rq26F2oBKPlM
RCQK2bzV0QI38wO8WYPlsDzKaaCBatX8HBhNGsUuA+z+R3B+8HAQgtG9ZvWCu+Ip
s9xyh81olUgs95vjQ4ISLqPDOAr6WNdrjbxZ0D3RkFngtUS31tJmShbOf99hP4uf
St7EHnW6XX4uVOtKJw2WCP4PtyMZN+hffLA6mTZArMrwfrPj012Zt+vU2Fm/BBpr
yLD1yCEXDg7aYX2iHPjp7WrUWTkYUCBQf67GWWnpVEabliNix20hf+T0LEQTNrgi
nb93n+5mjg4RaKXyJpZ6Bxm45D6noglPstwTX2XMNbiCnd+hNcXJbXW+Iw6TsO3I
LB6iGdBfU99dJfdSvY0kcTflqxMUavvWCfQdKFfB2y+G9YlYAC/zv/puX1UazOAO
J/LYaTqeSTwfA1uZawv4Uwp5Ws35tUR3mrU8CSDGWZW3n2cjz6rtVQoPVmfDVThw
cwMBLclkFpnjYZ07saMsjfV0KiJDAzWJ00C8seMlAPyTHBl9ctwbIeq6NJMVaBEm
g1YBp6a+IGzoCyNS/ZmLHeXjYQ7blMMGit1VgQsMVCG88Z1/UUMDzYHVKn+JIzd4
MWM5JKS01KxkHHkGE9JzOzk0tsEAZzZ/QbzjSbIIza1EjRxA+900YssvpPKKEwTj
R22BrTdsEyOTzyoHM1kS+YJgd1k/B/gYuvY9OyeGfRBfyOhwnwnAhYkQPH+WUQKR
VweKVt9kWSQ4DBGahaNa4BUcd3NJ5ftZYYhTnMqfqoHJCBpJCCo4NNXYuOKhDPXa
QdTF70mX2zJNyyUKiiIxW5OiOKKNoTD1BujVRQq/PCbqE4TnJGmzCii3zy4UzzWo
waL4egqLJ3eFWRuOIqQfQ9eSzo+d8EbBhMDbrVktndLvmvrFqmtjwDt1mhZkCnTz
7XQpTiHdQmdALC3dFEaOj3ZQ6jhGQEhHJNjgv5kFFopVWsBIHdMcdXd6Ducheals
ghZdINXTmjGGI7SgPBBbiUSCztQ4NcnaSJR8oQDrjkZIYtm7rjdPN9aJKoNmptq0
zsVFygVO/nRQZx+14KyJPQ5GpFE8gBeTefevuipzf06cv6WRtd8QaC/wr4Gq+mZ8
eDqdHb8UTEoIlIP7xnzmS8J5Rp9bY5IYfoPwmt+Tn731O82nzwYh97bJ2MxG6K8j
7Qp+sFVFNemuZxtadgVO/Kv/jsFTJ3MLYMo4BPBf965AYybaHWXhRFuR7r2ZO483
gfp07oyHX8t1k0E7jxn5mVIQD8L8MpVgJrZ9GPF2wjegXTHp/Li5vHlgHfgfDz3G
A/MzmaXKPkfKLqhtqUFQBP7DLj62ACx7QJa3GJJ36r9PLMCg+73oTXEjIV4/lmIU
AOiDosKyNpZHb0GGyF+phwqD81/bojjmcjY5MuwHm64vn1XSom7FgO9G1DG2bJMI
+5XOwPwJPVW5UbGHRI+SInP4OOVBRNXdm8c1Wxdv6tduuqmHPLtD3wIJDq31d4gh
83MK7gsH0Vn5v0awsZFiuyVdkCDd8cJChuNxgXbukxOsaku2ZWvzmaQ/zJQTfI6v
2jGo/TuOMLsY1v2ck4tcLNbVxXaoes0EbvK2cZdYeNoELlUh5IAe2QeDtzLRDd1g
PiCaj0XOXD4MN1MzdZwoGgTVwcygbMoy77xwQhtvzvz/yI8I8/uCVy54t+bdGBcO
5iWuG6Ox1kTaPDlm43ZLXtuLFjc86gOBHJvcM8BkP150b7ZN9G/4wFwwYDnF5rEi
NE7Oou3WhmMLc0zBct4v6GuzC0fM3VTzhJDgrre5TEPJrRNL7ChqdtN4Ined50W8
G6rxTlEwgCY0de5bb5dQOiB52DbTZnuXGlAsDGwQrqZEsuA3uIX6TpZm9EOrgtbm
9fwSeLf+kqyrAwJ3jemx4jutpC1b6hLaOJrPZbhrP7HgOc8jOMiZpmLEpBvMjkPS
+eVXBq5u3eQKDbTxJSSWribvLx0suQrrD6ATyNv91CHqIyNcP+O0vJLlKB2kGiPv
Vb+VNp/s7eaOd/P/+HRUxu/hyki+WOf20lRNiGqpFe/H3UYcXAe2GBiMmhph8ijj
l1Tq/7gzWj0D4nfN04EBL+Ff/37bCrrcNZTIeNUQkPdaAWBET4Va7epJjFs4a7RM
Sy2WwM9o0OpOSzkqK8hfz3TROYfKpuRX8mu+0SnEa1I8cG7GQhsRhT+sLErJY7O0
cdGgDa9HmxBEZD2NQjPsKC7ZY7IhaUuh3/+5YBEYkGvDwfmTRQxV+QxT7wr6LIdw
J0y/oCSDBDwe431jZvJTbca+K5GFiQkY6umtfhRuBAuA9UMBtwoa63/++gJrJVW6
87tY1AKkhxf1+3hRqn5bJrkWQCPp8s7mjOtT6Oc8o9qh+1ufWKagsc8gyWXTTt5S
R4Ly8/ZjffWLzt+lFdHN6NCdLUZ8pcyAViYryH9GGTJWvLup3XfZ3YYl4HoFrHL+
KF4SGB0hWa+Low2hgkgRTvIXcLlf9f4IkVnOwNoUIKapgZ7vhK01Zk8daVo7VM0/
/ToerMh+SLYS6tL/00Co1nae1TnH9hUed4tUO5budN0+1iukF8b34BRbIpvY4sbW
IEJnmv6bOoIMcXaF7o/lx2CWpOVh/HmIs7oB13uy/POm3PzHKQ1mr7litwQ7Y0ww
0nn+oP1m6+fK2nmkrCM5F/F4KQRGuB7Vws4XZ+1qommmE2Z2lG4r+nNi7YW+UmR7
kq2JUZvnqaFdCwj00kCrSViID14/SlDt+vatkqjspLUCmcRKIy15tRNzmXEDz5N3
P4RHLWJ3Vv9aMd4/6EpolToofsSxsNiELr1YmWjwRzUENPcEIPo1uC/Suqm/FHym
JkdwHHzr0yZY2BMyMykSkhYvfsSsDYDXHZd/MbapeJo6HJh3/obXiSEigyftaFkZ
hW8+ebgQYByYvoMv0rRdb5C6cG8ES5sj0zzZCfY1+TFbJRVfE0Il+D9kUKiV6/lI
WV8r/C7WRqW5P1ZacpSlPkXGw0trKrYa+/+IXRvHaejrx6LPsGD2tP7eHnR0kMOv
ZcYZA8NFbcuLpkGSGrj2HyBL/fBcUJ1B9IUKyPq8VsrdB2QWc/Tj4XXzsT9+H1aD
UL0lotKiB8/WOVIzEO1YHE8QEmsj2Fla+MHjP7aST+ZYuImYXdrruv7X4G3V/UOO
kBEQT6lI+Gb7FZDxsc4Bl/2BqmM4CnSv0JGnlJmdJBE8P4HnU//XzwNg1Mn0a8YM
p7DAxRD6a9N+hPzy8zE4bEixA91Q7iYALA50WWek4GVH4MGPY+U12fXeZ++pfSw0
tdUDDG4xZSdlRFHY9j+TQ31kc4h+MdtOlGQAuXITfl43XbPAKiCTIedK23ON5+Ar
nx7jvxELoWKfZOLwCxNgGRyX3FpK0hnkGQMubnpXRl09+b/h7+SXvDrrG1CQHC24
PsKsF7RUkFvuc47yk/vjNi5yCcPt7bdvrBOS9qxvMLnGgmrCv29F1FblqyUksTOo
m+WmRzzHUoev6zg726mU1S3Z5B2kL2H8hMw6HDQOKzAPn3ecwBNbf0uqBDRO7hlP
xb9/lgLLHQqZcj+60ze4Ro74TAsnMQUQFIFmpLoEtTjJzVUJxFnHyqEQkWNOPhK3
N7lqjzUFEsLkOcGHVGn5GASTuvVuar9GXUNv1BG4rEPUy8D0tLthTlBv6D9FIwqf
KoSfq3rZk+Yrhz9L9Xy6dhfbRBwnL719Q9C6VVeNvNC+oHtCbqRaHAWKznQ8wkT/
kUEMGfh+sxcQafsUQw/lst+8cgcKscfoSX/PF7Z7jfX0l44LOePt8qXsd28Vw5i6
uMFe8N3XxHVajPAxm5UXWRL8tTH1YAdWTux4HExGhm5UY9Lnpq2EW/fLxSKW4H3x
4R0GKvWDSLID0URJBNw8lj307FAA3/qZQxarCQsUcWb8opBThbold1pCrIcXdNer
WhWAvUOseccHRd0506SXmZbe2e9wWQY/+duLJdCz/mIZ0O2nIsRUC1I/BYhFiLNB
E+y+6oeMeESIVTi5iaYx9ekbLQKyqGhGDpz49OqpZeRlFz9qXVx2dDlYnbMJd21L
LPKFDV2SgdWv6ZgDbLhaMDrsJxWkkhs+ohGJkmniNpNjDy0JlxIbZL3sJNjTPTJs
UVVkh8toVFKzt2LiLdVBdAXrALIFen2VoCPBJHpO0Gze0Nruv1Nt053uXf8t+Va1
0ZyTdRC5cA2rxiaOsU9HWkjnlWSGqxIGxBSCxeVAEXutZA8LX1fHfooO9Kjar62c
C7LC2ab7hg3bTQhVo196dS+OEUGblHqUoy8bMt3rI4PYVv9D/82rK4WaSrprwaYv
rNwSNynVsePnQ5XQhZ6aCcDEtKCoZnpcZfqFjQP7AyCBupuV8BrlMA+Tx4ducg21
Gc9zxzk6TV1xQrTfBJWEeUUC9uoVNVdWJX3MjN+paYB7DzZ8LIs9oPEXGl2Y39/O
wIvSzTugq5tjzxKX9YMuJiLcKgYaxkluAcwTzyDVfGj25824X8I9tDgOmfuDJckD
fUYOyDs7p11BsDfDnSlMxeRHJ0pHUiXHwyxBk6BN5CoOVUtE3jCvFc4vdN6uLfPb
8uPNMNczG1+1WJ6RpMUrXHN62wW1ElIEN6zvszYGf00QkUhJa8JNEBuYtg7akRTR
KIkTujB+lY68u8qjks0ZMXGEoTGcksbUmXcNft+LeBUudYkvUSK+YdPmTM8HUUBO
X0yEg5z95xCXzoWBpfGDWTDQMJn22ZbQRsghqUWc8cSWqv1vZsp3ftJv3CsdZu8c
P4BQ+amfbrsu4FqNjMK7W+5qKZoKYHK7M1mgwIXsgvOTfF4czbPoso9YXIZiJZho
HHVH+k5oVnnLgItEiqPw1b48DSpvdnyjxfckN++LUxiKEjzM+bzC0HkRlZPMBT1+
itNkBr9XO1Sa9mWuVABvOrKsQ/xR5pu9G1WJ2aiPpyWq0jfdBfizDDK3cgXuKb1p
QNGNLzKCCS81uBfapst7EO/O4IwQ2dbQceYun5aLtP69gtpVKxQZGlW/bHJ3GO+E
p6pkCgIQgMPKj3ao0a9PAelhyfekrB+86dNN4ImuMD3VTqgvpgQYx+EJBfCJskcJ
Yyqchcy18N/yYBSjTytWtnuHwzDmIdCyQamauFy94B0DBjdhcsQlUm+nSMamDHkw
oB3U43HODyoe4iFuvKCaOx4WtwkLgYssZEappy4raB7gUG7KxgVZl5C1BCcuEl21
N+IcfFXaobC2IRJwssgj6HoVVn8FdC5COeunDfsqgqxD40F7h155k1gwVhFvr5dL
CEXNtfQKEZODau5uPjLFkDVOeNiZq5mZDaBmxrPJQleFaVAyDk1GCR725ITgm+BH
ooCzYfdgCWQpUJulKzMRAc6M1K4cUHWGv9W6jYGgjhcqqcQaRGIZsVDoMj1ZQ397
HicU1/vyBfruo0JqwTNZY9ZOD6I8CkJ32JPI4A9lcdPXpZ3afFDQ79UpgcDimxa3
caxi/vliNbY3fxiiEhd7BXchBQhLgXtcFavdv8co0cFe+240sydNNBecj09o/bW6
2jux0UoTf7ghCMx1Mqd6OdIFQtWNHHtqWftDJVgBpRc05aKJmUjTzDUmH3BhHJWk
sdzveW9MokcVgB8ZV9P841gzI/lsa7lj6LIqvNGqgbRWa5XMeaizMEogho9GyQwB
fIcCO0BPCQfvQC+R0o8zcs0rFyxgbEryj6aV8sRrw7anc0jixZVs0bKltvuFhc0C
MLhOtu/wigW48+tkV1dRMbrOM5bm5EePc+91tjtYKE7Kq5y+HcD6O9PnJiKM0pEH
0s7HEnFoUfFrwJ4Lp8R/rGdyh3V36vWfohecnbhT/tEdMF+oQ9FfZvVfRg5M1YhR
69t8ABz1cnj4VFW0AHc+zwQyCvtlfcV7VGvg+190MgopSNs3+vkyWala4XB1dh02
wb0S1YOTTKhAdw7fveJBXcqgWK0qq+IoKGAuFltggf17Kg0NBJLmwv4TTmcXEENS
JvgFjn6EmyVTVXey4p3C6c4Dnpg2UiyCxZRc9RzoGVtWpwFvoc4ZZYgSE8FIjobS
nAEFoGTdsr82WGgMkAjKepdNUB2Hf8dbyvSf5EXqnH3WMbuCOXo0543hPVbOLDKC
tBzvdUBAw+epv3/6eo1VSRqs0TPBYAKKF2DvcD8jNEqbL8xU6X6if7uhw2VSKC0F
8eiztQS2rjN3VZDafHGYPMPmzRgrfdbZwi+q4ZBZeJ1Vvw9qTyLIkw9Ypu6uBXkH
TWzfJU4avp4xbU2aA+YehfPomFNf+9wqK6bEUPeGjX8CYE4C/UInknv6B5oIyswo
9qYR6vOA3qTdA0Z9XOB6pd5lIzKX+Xbt16Fx55OfYtwzAuwpVpuX2Fo1f3iuORkW
7+3STqCClaZ/BVljzoifYyyNrHAnvvFfT7shuepLnaA9eX/X7PaCGNuWkRLJaka6
ySsnoCf8NbGdENIw0GVuKUUFj1F1ufYO5Pda1Ktp2CTaYmExxxazL9OnLaMKNJBB
vbB+u2buoBgr8llNj8QH+nbU/KE9tbcLDJGys7r1be4zEsx64ITNZGQ6PBPnyfLu
fPGQd6RvtHxyuzlr0YFMsA4CqSbNlnNJldAb/VptK7gNkih+D4h/4N8B2FBTQVg/
8Pa+u6e/N2Fvtme9Mowg4h7vVUUJJX+JUSsV+LkXaYN4lQJ3OmyJdwXfY8KNvmEK
+iwhHn1jgAbYXBmy9SqOeqfz7yRITlrFSS7PYrd7gEvOEHNEX3+U5+kovrb8oSaY
jn4x7G0gVbr9sfrJMPyU2JFlLBJha2HD72Z9VsFHHUVpgLsJH4Zu1jVlTObUkD7J
viCjC+IpRgP9BOkqad0Vf2VxHHLFlaCF9tJk8VD4qvenCiNUQriI0Co1NpwskSXL
pjvCQ9J1UWaZ2CIJdW6jC1M5rg9pgtGvU+eGnvtty1XTPhK9ONGkmiQtnNqb10ZD
7/NHFspuyTvZZUHFBdd+jefO/1raIS/wPx56YlxQOq1EVg60JIE3MMZyofCkkoIl
d78nF0FsXjeJy09X5QYBueAT0Bj6jLzdCDClXZsYeqWuHrlRIrtfzMgEcXRSPswk
8AKkkby68c5JvbDabwacM4sdi2fa1EhcQSG7YiIJWuiZl6EEEkUv1C95eG9U8Dwq
z+0Db5QMLPyTkUFASk98aSXwtqIHqgVVesEy1uTxkxQ94NXyXHnOy+xSsTSC1LNX
Nd4+Hlx/F8HBMU+2cV3xWXOhu0HCmfJ+i7f+h4FY8qFxadqyLR3BvQe+n9/bNUVV
wD4DGban+1ZQWN30KWQtz6xiimUQhkLlX3w/QfJH+Yo8VlVkukp71EDWksSTWIjl
SSfUjL08IrY2zLDzRJxLqqixvKHDQcNo6V3/8xUZdXX6lVFYBRTSjlUAnjm+2hLu
q4Ne/pAg5b/BiAg97XCa9r1uElY6OOiTHVDOGokpZiqfsoDbrLbz7GDLLBM/wLF4
BFVFgNwBxpqzz/3aOfCxH2SCqSkbrpBEfvLIHHHkFpivDUzs8W5wqvfHCyMb427E
SreJFgz3LF3pY2rfQPA3CkIpjA/05HKEELPFL07DxPbQW8g6SjBljljKR2Lh6FLQ
KmnX+iK3UsJqw52DMDQQCHniEE8x3cy+yjXjbEFaidmFXWVZ25O31DF7CMFmfLJZ
s8kYmLjmF/IP4zzUcZbu2FM9+11vzzuCgG+GUsswX3D9i5tVsK25f8xAnwSjM+yO
SoXAJGQ4eZmfnhzjQjDGdrNxsjLN0JD0M973OI1GuCF2INStnr1vEy1sAoaigJN9
MZ+WOADQVMKdGCe5oVDVAlXEJdk4vJirG90Fke74qxjcoghrgRDKuslX7EFH+HZQ
hr8wjnMXMv3/mu6NODdE6gPxCKscpAzbLzp9pEIoJyihzwIFS/KP2NMnBgUYNeI5
/d6Jw8WkI3LgCQyriBSCOyT0t4801aPdgrbzxPs3t4/4EYK2Stbz0WdDb97sstSj
IaKWH3dcFpApiF+T2BsqX0X2zfXl+ZtWwFcPOXYBp4MTf8+paKlY+Ltyi/l0gQcH
s67RC3TILJwxx9fe108Jvm1z0v8Vg1LeJsdb8iO4Wr6iWh5699nD97n68iQyVgR0
hr4NN7mawVcQPKLaBaweSc36y3X/elkXysLYnB34Uab7BjuP3b9GSmqdtAhJKltv
rJsDrbT7SQqFWuw3NbnWCgrxfyC3S/Eo49Z38HqtsXqiWFdj4T+YhFoCE1H/HAIT
aXwa/mFj8bLMPuT58u2qVlItBPPWztnGxAKQq9WKo5OHEe1bs4/7ofwyki42ieoG
X0WzT30XBrZ9nOLyD1McZ9URvbpdD5tIzwBMieOxBuPEJ9SqlU7YHo4qE2v2BlZ3
bhdSu7O2zR8OXiJJH0FGSnlUaNR3tJtzdKQ2TA/GFciLKfbDxEm4hTDMh22237Yk
Qwouo2Or6Ws5llqxyTgmVJdcZX8eopr0XkwCNzXk8vodfzzpNT/27V/zzXbhWtTW
zKc5VaCKmP70KYs+pIkTZoCbbCacUiKnPVUY4YSTYzJtx4xv7OMeK5p918yjUlVT
wC+IVjLsiRU5Qe2veZKzJXNNuAAQqlzmtudIfeqB9u0KZF8J9UNI1gYnvNC1NGPJ
ZBm1QhgNCH7SaL0GdL6UH7S3/C/r5HshrF5dprcSp9rwXNSFckOB+G4hX78I7HEC
RV6u+AjEueQx8d490nAQp6NJukWgsHYBw1icUBRH9Uw=
`protect end_protected