`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aMReDmrPskJscpWYThVKVItA5gecPPZO1R595p0GoIq1TSTG+UxXhmmUXc+VYHJ3
u/C3EW5qePLufxmXxmhmDnr9U8/cYC1zLfk44v/2OPb1TBrTsludEDQZdGNWeV9l
cPUMSIfZ0dHXN7L1M1E2XtgoTWQxf3VDHs7B7lU2y9Rdm/ibz0fWMow7op2nWdD8
gJ4QlNl3f9Oiotp1p8vz9RFzzZOF5gBBslZxcTF5+z4qO2W7+xLByngthWm+exIr
3Pzy8qyUo/m2DDwOz3VJSvSNm7RUq+0/yJNOOz3jr3j7ZyCj5OqT/jDAWjJSMH+i
2402Un+wDMOQxi21JLo3cA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="5R6K2aWI3OdbT2A+sz4o9+2XAInTqB1/cSw5W16RnA4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
Gm/2BIZF5/H5qen8uQizPH9RftTuEE9mgEOF0SqeOKegtP64CfvEUnIxj/ahmIpA
6xUR2v2l7E5duaLZh39Mc1GYsfqE91NCPU5whLaBPg0UuX4cgTkO4cYbW/7yvcrd
4wavUfwXEp2VSiN7EVxL8RcZTSMSI0Jr/aojiilFqVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="TEmQtJ1Dsm7TOzpJk/CeTSSFx/zKExk04H6I8sT4Meg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
nvPqn26PC4XWLLQG0Fq8XsMTlhB4evbpiwGjZroFFLgtNlE6bBjdtwWsB89WW4j7
jNfYbKN4sBv0hDeMH0AAR+8g+TCqoX7yLdIUd7aGwBUZJr6FdDs2wTUxRkXFYNTL
zJ+Pj1VO7cmUiJL18xlX+Jculsg488x90+6wYvbF3oYtFITcg6T7ZmYrFycbN8Ef
SIyaQo39RbLfVo/MNp+PErbJz+fcC9MOprOROVTsIu4UFt5RfKQcjO6tqwIiXhNO
UK6Q9vUtSkYHqBF5lQSWVUD1gx4znq9cKyKbhaonVmK/iwdR57LhxuyBHazLh5Cv
wJnUEPYuRCVpt9fetiCbt3c5OR1WBIwYwWkdmAtRIbS+m9N1xe0kQhLVJLTSNbEg
IPpoQI+hYS3nIBqaM8EG2/kiWiC8QZsnkfDJQMBB/hpPhmfgOZWWayiymMiCSRpK
pMLYjtHT2u1NFT/UTWs7zh9Jual9yexFVSvlLujsQNxMcq0+oo02qOCGNrcVCXtU
KSsmOVWioAzolVcIrqZ8fRvRNoEJ9svQr/o9fn4CTQJJWGJM4TfHd75Wqt051B4K
FOjJ7Uqe2yi5+vf9KRvsNP+FE4kRs8U/DjD54V94CkMSqdUfTTsLvkUB+YaGEzFm
h35DjacApGGNn9nS6+eAyz5s6BU6JRcF+PRk+3SfQqskBxoraBY2xUJ6BvDVeyIZ
uPgVGIS+0LcnU+lQRcQ1mh5fxTovSYotUg9hDB6RGT0s+JI9SbUsuD4pyttSQ5vU
jVIVnfa1rj7yI6OZEC/rRRoX5MSoa845IAF9L3MlWnuIIWECUaHsbk22TvWHE+My
h3P08YAUL74cMzCZ/kG71twA6ILzWEdiW3cHvgsol+JDdFAa6X5RDbNGr7yycFYO
bKb60PoV8wUUgmO8/AnZfd9576TLC/TfQBdIRvdFgBAXUcehLSwP7OzfyUhwjnZ3
umnnAcuM6mf8Mw6FuKjijAHKL9VXaMewk3Mey2cmnOtwRKMEC7jRagpiT7ofOTqr
Wfn13kxm33TAEi+5I9RFGLFrG7IfvSqkfxcJ5mVDXttMa8CiOqk5/DtIK9bTs9xP
57VCSk+wfKzBu5CqCUgfG7AVlIOOMgZK1LR9zyzN7KI5CFV+E8qL0tq4TxVsmEtB
tcbZ1Sm7PxMR+pxWwTDpxIXjfIcaoLJbfQVRDD62eH6TM6sNcW+jT1BRGV65xwG/
B5oW/QotfYQNwfMMI1ahUCI6JMnqWy/HZygxu5CARrCQVCK26wrg189emT1BPH8f
sy5cdvKB14oHBfow3ktfRpvb461ZA0QGXhbFRBC5HXG+MjhifHUEPg1C4Zo2uSet
QKnoviAHuuigNRtttxDpN/RiDCOckjoHbvPLCsz4J2yJgPS+prfg5T6EEzpMYOLN
K5kEzMQ12j+gppTeWn3vm6g8/jrw3TZK+J2a0UD2ffe20EqnP3VDwOvS3vOev7Df
//7KAr7gKxqxuduhON7h5w4PxJeINgFbr08rVxh94+RY6Go89eVDdFPr9L+zf1zx
5rCq/JzCWx458INrHV2exD8GVOfGhnYQNKCorZYWd69VPROSOTg6BWMpMufIO2Dm
9HA7P6m06rUQ3oKta+pTX8BcFD6BNxq/y361NDCuLIfUFxlfoSSRoz/dI5Ej5MZp
/hCFSR9rUlIinc3LQwQ8ZQ4Bg+CLo3/jdzCgrS7Ha8Ce6m2MP5BDiix9SRpo4XtI
7lw+Zj/0n5BHaPFvA695GCRovhWPyLSNTM+Lc8RfdJ9oiNjXlw8Mv6ulvtQ00xmw
NTkXTlB/Juvz+TEli/T7DofrBUq5QuGNy/E3QrDjqJIl+/Anh8kVD5AS0GSZNpex
BJ7+INzn5UqEW2I8JMZ4+H9a6Qio4EukQRaGL0A03TDPe9yA2duzfNenRE0WfQPK
312Nn6U/DJB4METL0TQa+U89RxPBGfw91R8T/EWgMWgUjBnS5YmZrmd2ntY3OQeJ
YIDpjwUwQSmSB2JG+BWHnv4UaHRQZyLLmp789SYSfaqjumlmHxbpDJ6j620VXETA
43DvmywGYSIJ9vplBlA6Pz3CT+Z/z5gtIYY9lt0YxTgxv9Y/0MgwLc4K/NYpaGzU
BQ7lLApae8jX0QrqCjcLIO7bUNEcifxmFRadm1guoHCa9gvJoyIM3eiFFtXODLi9
rJizsKIH8UQXYSaZxBarsE172pgUZqAs9j5NSTuuiaIpIL8nsGQsWO4v1BIAcMfY
QTVrpWoA6JRmgMVh3ZTPhqNPt2LdWan0k85vOOfB8qU=
`protect end_protected