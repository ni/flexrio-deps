`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1648 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
GgG2UXwpbWAyDgGIJC8iiPKHN2h0P+peQtw/EAJ3UD+Mo1acXjTcN1QpzghS4Bp3
YfJRjT1Zmd6uaqvTc+hIPlJGG8z2axyrrHkSuSYhB9k1WCRh0M4D2szdMYTIHiL3
GSzguybU5iUyYXMXd/khnSVkb3D20RfV/1c5xZCsPihgY9VukkydAAgfo06XrrG7
YfNSBSIp1GG7SDeQdT34UrY+V7mUaj7DcypZp4W6tyQXIJjkNi01tesngWG8ad4l
zuIWFIZAsHCJw6FirZ0WiMsQKQOrOeNsxQACTrLDDbyfEB/sge9tA7TyBPti0EcI
WDe6ZsvqNum1s3rMu940nU3sJIDtLBlNnDJcCHv0UVgzi2oWXoExGDt3onGTLdcD
EiSyzmTZyrA96ToJvBA9JiJjVuTarRiDmlMFuxTgG7zVQTjgi4aFH0gIkPivTjuS
uQ4kOO1tJ5sUcR5kSoMtk239a2R9KiLDm546YhCrSMdtqugRQfsIWS3FzgJwvxjo
ZCyeUqZGfa+r6M0kXi7XLXVaWVTpBv3x8tI19lQR9XXTlV47rdAVtaGh9pu/nTVD
wjvXLFotZKpNk8wPuhiYZOTFUZcHEe87lMXLu1X0pKpPjGZ8AzA48yDePLf+QYY9
0S2s7pRo0jUG2bB9oC8o388hcp0L4219onKJKoQ4jRNlyTa86woipr6gBjYgxKmu
h1RN/Yhkm9BfqHCzAsF82bgZ4Qgh3OQ2QMGv/GTECPgB0uKLZdYtIwtJJxdhgsap
/1zwB800GydwEGHJENGgP+SNJNLMWdzBQ7mNkXVAPx+HBb4vvGJY75N7ns0vtwd9
wMNOAoNqbJBqwPZZhmsusGBqithv8jq/+D5T/6pPvHGFPOYcyUSJna8SvorTbN8Z
rcBjcTlA+2yzjFc08dNhobe2G2SCDsHw4VctVog3dMX/xAJwbUuHMVfCrzJ6qtre
YwAvkhGJ2Mu/JDfWYmuryJLsegUPCh2sociBnucSyRMT0Y53bNNz8+LhpngQKcyd
44cQCy1DDZMqVXzQSdJnrM3UEOcD+9Wn146pFO2DHBGyK0EeNgVZtJ+OaVCs/xRT
XkF9HQ/HW4pR4t3Ss4+H9bffEzNpv4XqqIAndfAi8ePuUDrXGyO26rJnp7IGzdJ0
9yWU8SlkBGbT8wNKlFb9Vu01Yt+nAPwfPlnjLxtqn4QkC7w8u6YudcvZxfr49tcS
bC40kwdg8Zv9qm/pUd1A1J0+LqwBxfKXXR61R0H5dNk3h09MLIjKqq8onnjquTZu
J2d3d+PDFp7Qgca+orWddhwjO8QK8+f+n3d9x8uUtUHJFSeJFo8KLfDcYt6BzVJm
EAy/9aCR5kQfCwjjPVxcbN6Edb7hSXi1q5DraxlDqBJR+kQlv6PjgWY17BT+t5Er
OngA0/tGYFy2xq43rSd40fEDONFwm1wtsxedNHZDwwBu1Gk+oKF6xsBlBb88H4OC
WZu6FC87QLSuU0lN5JyyMpp+89X6caHYfsrqPtqUGFlHDvb0dftO81lTL5e7+285
AEm7kaEbw2p0e8SGzhvgZw2zUSo594PLtQznDIc1RpqXaoBDAXq8iQVjW/XxXORR
1ogEcOZNt0FNg9VFgenRc1o7+NPomRV7T1N+0YvyKNZ505z78bWHYryBMjBfHnwz
eByjYkl60U06KCqzq/wlU0khaMp1dJX9A+nuNeT3rDnmgv5+RszsLglx76ZH99eI
wYjBJ/86uk2+lNYIa3B70BaW8nWJeFF1q6H8EulOwmNjVxffkq9uTFbtUIMbajSL
eij26rLJHK66Wga+XZ4p75gU/1zh4lYcg6Jg5A+8oBtTHVT5Y+h8NbJBodO4ti+m
1ML0SLi257b2sd2rBgzatXsF/FtT00ri8+Cgtp10rrCqQUoyvoZmTvIZj/XD5EXq
XdlY/NGkBqKsPUdL1Jcl1yV6qrDDga1JtVh5saE9EscLyPCEa5NkrrPQQOr6ur/9
XbDQ4VWAFkpbfVcVZWyiuY84S5fOjWjVjKuUiZnLc9hsE38dgLY2RBqUPzsqxTxo
YnjRv8gftzrFDaNPcMVLIw==
`protect end_protected