`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14192 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpukXuDUJ3ozoHBU3zo44aVFEil6IFgm/mAud1E7fNZJz9
cttj7Z3V9joCmPUc2dytVKsazbSGQmMctVMV4q5xeW+TwHuCpQMtu0vrOBCPoQ+X
y9M3LrFDiZDJxwW/5i1nLyDj08SQkOYWycaU5DbsqnU8lmtzIteiMkQjPSvJHYer
yCQ09qIVxScayBqKEr5E62RALh7y45ubW4Bum8Pa+EAgaqQWw4brMBLqfcL6busq
6D9vMoNLe2CJNvMgJuIybVMbJV9Ie0WrhikgatLzAjilJxkCKOEFPANK46A0Imzn
KZKXCOr+Ma8OMXQSJH2auMMmRrS9oyAqk4zN6MPsiqBcfPiN2iX6ItFlxxZjxs0s
wu47IEgdcNtBPV2iAgzoxmW1QqviXRN8k25S90mfWKH20Osa8/5v4iVr6IW13ZwQ
cKXyp41ao8b3oy+G5e9mpPTlVARh6FDXnAwHmT5WBiUVmwIj4KPem7XWJTCvSnsx
+TNLGxuaRrgcXoej5MHbKlVy/Kz6tOmZrwg7tzLg7UnMJ46LvDqQPlkBcv8WsHeY
RKdOUJ0hdYYNj9ayoPEDDGGxxTVpTvaRckxk6KlBytGM5OMTEH4FGEwBr+5IehJr
pAkz+q7OIh/xgTgBf6WLmkyzul2eg0OOIpgyIMhicPJHhpk3myv68dTBAado2UMZ
k7a4UaTNHPw3xndeCoUwWnj5ez3TKaNn/zNWgbNQ58imAZLQiD1zN9n8xg9p0H8R
ORoc0SjcnUF9uC+kZf3M45ywtNWzpoPQYZWFdIWpyG0IDsDEI5cpv6+ehwUD0QZQ
7H/09mWTF/WRadm2PgJXrE7NR5Kzp1qyBdvxXOZGhgkVdIcEHCP05ldmCFx84fNL
pwnx8PCA1bDNCQG86K2DCVhr0IVFncI4pkZSV/W8MCMhHKAYNY2RcHlorac5Nuel
Ukq3A0wZ/AOyUv2pnccsaUQyCUFuQ0cbMakxR8hjgwZKtkWjhETFp2VzOjhNMYT+
Sjudf/1RXvuxlOs7/JryMow6uomBSRPNVc+fkRgbue4s9l0wtumP6j5lado97bX0
dDmkKl5lCWz7XpzpHuL+k24OBvazxa6R13emk1SXlimZCUo5k/fzdzWIGC7RDoi8
Q6CvS7VKAIzb1fMIpyWoHI1aRyIXVe8gxBDDVDH9fBA1VQVK5kxlIzKtY94kgmyd
mk7n4rYJ2EmB8kKmVf3RjeaHECSjVZqd5LkeOYlRlgOXNbZRwmM/XXcPFReHYPg6
9jYfY912sZPWpftUxH9v64DaX0pSfQ1P1FP431gD56Ro8bvel5mRevRb7+gmC73p
nvw7+BWMejogd4DnogdAyteoWoDJkw0yDEJHlMm4m9NT6Ps0TSpP+qm6wDUAPGrW
03hk6haHen4E/5MWBa904VtAVy95gPcfhzk8z53/5jzHZtNH0ny5kUWb7KYc1/I2
LPxnxf+q5eXMxjMCkbzIzAOlGd4lXxjoG8jwd7QyzpZF/iehx5wEGdnH2l/354op
QWkSL65WQ9s52+k77RAZZFWQSpuwrr+9ajroVd9G0sNnZklopEMgTYiqY9aZLy2a
s37JWopRyWqnTPHxDmjCirMVY4x+a1q61c7rZucEkLXPuK8Kjz+9UkfvDYiAKmyU
byR/4Bdu+y7lcrbGsxWelI4d/SpeYmBQZsBSgzQ2RwN3j2vkIKMd0debm9Ts2Oyl
voHwKRHBUQIDR5fjzyVy6W2SragYdF0Fbpi5uyhU83Y472h0f/GG/NbQnA9GUwNT
40XtarQUF47XDCiuvX26u9tu/fC6fKeQ4M0XXsoGhAOu6gZxvOZILfPDfyt3Ck19
XsqcOFYgK6NZKHKh1PyuSeF8/BavnZ6v1td2DJwvk58xnIUc94M5UZryNMC9Ow/u
O+mD3Fd48VDsE7IreyIqNkvOQvyQyAjreFysDe+0IgsNbLDTBhzD+A5A7Q+IhF0z
aAgdhOlSwj79SBlK4s8MGlohtlnKtOCfdG9FNzFiwQK1Nho8CTHnENHJzYC/Tt8B
8DFRwfw898vRqwUoqC0ZduqZKGtE8BNjdHE/gortOVNP4jjBeJWm21YHLIHSTZhx
awD52S0GuojPIomY2H6oaPt/rsYMnBAPAdl9oK13Tr2A7XJF6qRm6QgeaKDnZ3fJ
mEoVqYUD1Le9gHReFYOyk8WHji048fzy8t6/k8L/5eZ5hDg/nGE3O/wyWb/U2K4E
DCYqNd0F4WqURhrbCE7oJur+j2gqBHnzyqQ+3HkHaOmfv6MYgRC9GmI2+/tX+00b
fYwJlAekTVOdfYhEToRNqjNZ6vCwix1BdQGdfOsJJSGdMwpP5BagLTTBljmbw3Dq
SCJss0JD99svHhfue+/mWSMpQNbjyCz6z0X9wU9/E5UXWvhn2KwsLzr8QjuSxY/Z
hA3VhIY++4MQZF0NtglihynV64DaW0vRz3iFt62j14XzZV7rs2fhzGJ5D7gNCpI5
4phrR90B6Yo+qIQJIYyOIeTe4vxRFu45X706aPOMJrFGoK1hhIDNxEG4rGpw5qMF
866nGCiv2jbYsgzdlpudbQ24Hko2mO8WBqCrzCSvCuV/we0WS/e5lewVW8M/t93l
glRoRu6td4Kiq77P9D7r09/lXjbMu1L+4vUVck9/av+xBZZ+DMOIiR6f9gg+Pls2
CUHrDKt5JdpFwuerc4tQXKaXjiyqBtduGTr6uN8eyyh+JWwHukMNZpmY7nYNDuQe
IBukisdEmVJJLG/XZ97UymDAjs1xkdMoGrRrdIy4qW6gqchHbUJ9RwOhRXciwK9v
3h6ozSiW1y0lqUDLeYpdG/nMzR1vblRg93C++pOkBCrtjvVcUNGlA+BBN1y7vwIv
+XfQUThmnR+IJX9uoaANXkpxZyzQbtPG+iVvhHSXKF43XNwObU2+BN0L+9xiIkeS
ufKY1BV9VSuVs3fBS82SpbWi1E8svdZ3Oyuxvpx9/VcIJ2LpyllS9Haor392+IMV
isR4ifJno+kqA1jJXNooN6LuiAd76IcZXb0BQPrvT2U3V7jgCyPy4wdosf5QE9F/
M0JZ3boinUOeYS6oQtTeu0ocwaioxrDm9+4sVXXtW0QypraP+6q6nPNdPHFNhEwZ
F3MDuqxaPJzjQNdr8BpZQLOKuFN/4oPy+qvudMQPoOxhifKqaEDTkREsC/Fb5VzM
QeS9P0kQrK9uA0Fipw2yv3tWEOJ2Qlh5M3AKkR6eg+VnZyfhIv+dA37fHxaNEXVh
Lz23qxK+kUH1FdiU1iRLwMEIU+QgIkb/55+mStfFU7E8ALT/qAXmrO+BEeeYjTW8
qP+oa5SQF4nWanZxIeaNnQvHt3BpuIUFIEncDpZfAgAOFapf0D0hUv8aeoZQ1uME
qywUkmhdMdophXDuSdwHO3Atd+xJU0tXNr0o8zFKnKKbjX7LmIgOmF+Ben9JmypG
+xyPO3GWnEVwNDL2FONyQeEngOg98nuBKSCJZ5tDt1awSyiF8AkG6mb+xXheEipe
H1+5lviywZSlIhDJgT11bkbg3DpzxfEOKDTFuY+fVNqoKMIO8sxCZAUu9GpdFq1y
l6o+Ghoc2ypGd21J72rY+EnvhWa5uiBTufHW+jFCtpdBnYr/H86h51Gv2NQJAdpF
qEaAQZeyCdkEXILxG3pPPqvYu8sOd7fNN9aHt7AhT4JVWPjyKT0jdF3OqUXSahbc
WYfv09yttT8K6uYXKVKzZjPX5hdCeigyKTYZ3lGR2HLK1eZBXe5+E96kaB5SzU2A
2+PPMQxbELR58j/Tn+0H0Uj8Hx8wC0mqjXwN0x/+4UPR+d56yQQ9UmMr9DE4NEpC
x2a0iWUMegID7EpUr1S0V1ue54FsihZmX+E/dX6HExl//IPTUuSCN88gCEuj3lzS
/aT7ktyOBlD3uKtOekhGDVNUd0o/e1oRiCHLTkg+nGqNhrwpBzR61X1lZDZvc9Kl
w6UXiPAQ05QRUOTzC8et6xkFkfZ7QF/tQE3a+BawQfb+z5omzs1tQBibhDk+20aX
ARJfM74a5+kFhPP6t7TbrZuk9k3gpkmi5c7EpwxPhyneIluou32qW6lB0MNsnKQ2
VRc7RdVh47LgL6OsbM+Gur3aPuJP3wT+BznYrlUwuurYZb1CHRrOFquryRpt8RT/
zZBJXhNDTesxEOBQu48ieUmphUVMmpvwfNwFbkPcOYWbeqbnwFIP8DdDg58bsHzn
eAFD0DaoCN2RaPcKD8KCv+T6aH+p2p3J0ZswslzlwtkcY2hd6EU5e2Txg2VZodiU
BjHkpuLiTfiSQgYZhJXuKreheKPV5bKed+3mJBthbL7C16N2SoJnv3NOifK9aSHk
x3Dz7uPCeOQH8GxLuWlaoBZdAGhayDXijDRGGfnZVS6SfdAmxRU8oVN3eDBxGITR
LjdUnHmn8S1u5LDYK803oBOJIlSEThB5VPEpwsI7ykPcOg1p1z35Y3ICxzxxtDnQ
Ii7+0ysAyGMMFWklI/CITeRX1tFwzMgwKvtxIB5lmjoESDYNmg4Gd283f0SLY5R/
A+VU93LItuRRBg+Nq1QeR1dcri2AInmcdzHHszeOpuGJDuqVjL387q0pon+Mp0bj
e/84Fpg3avjZM9skPoymAd70SXCyRkIw3Ha5rJQwJKYCTUIdyGkbsiPpZanvOMNP
emKNyu7IGOUQ1AeDfh2BCu10EnfBVnL9X4sDbyMc6ECei5ZdBpqPKyKsgelWTjOW
3rHmMhLo8EIt8lwt2TQf3ty0Lpj/Mp6AuqGktd8xqC2wI122+ktGMAxx/TujEtPm
nKhYEzjOkk9EDm8Zzh+BmFYNIjSwsxSw6YU11D4XTofsqpdiD7/I2gKXmIP+25TI
TMn/p04q9CfT2xGGmibrVA2zAUN3CLNFmBYOCmoj8AVGP2LpsLaDaMWnjvvimnA/
jRlsWlZQJgeQA1h4oDNjxTc9jEH4HNifieQl+4ZVRC8FcKXZduQoFJ5qpiF5d0SX
2z3ZJtf5ALJ3ZpoONkYmKLRGw0eokoBBXXfsPbXxGBeuq/y/UxZ0fW7qwYBRUTn4
NLVZLIEXt1A19esShyWzed81qRRxp+KXJ9CrDvMfg6d8IMus7ABHctbxsm1aAUIL
Dsx00wTpA1cfjA0UtErpkp1KHPsL9j2BkZxxur7YEtEEA2CWAAU8AeEXx+qJtX4a
ofKn5D8Lk0pskjoJ9qqRVzydegpCj32J20a/tR7zebdhjx7OHVkQRh75X+ULeqWA
BQSuzYv/SCJ7UZHkOzIU+V4tniW/iZNCepIyXcvUTEQOqh+2dE92ptvVp5tp34bn
U6CQoJvExK6By6Ubxj/1540hUHsFPe7w1Xm6VSGdrc1SSL9pcPg7xu10F60oVSKq
oHyBl3N6epqGNxzOeHYm624ayedHKGM9hW+FWuE1rWAoOOIBzNYOmpFsvt/HvtMh
9WIkyuaZirkvVv+DiDHL7EIQKFF+8K/Rf1sVHdL99mKphVNGDwIZxtygC0eka6T/
1kko3R8wpyv/iC1AV9VbyyN92cdHOMA+ulN+yvIDv9V5lMUF3G7Lt2jl0HbKmWeG
5x2RIi0jpU7R8ipuNXYVwk77Ie76KlRkQenp4Lv/yzeebhQNgLw871NSvmcw/V0j
aOxyKhlw9ShyqftCvK7El8SfI/3YBon3w5Fvr+/roBi5l8RhT11/yAEGVf55shUW
CPgPpivDFuJr05o073R3+f1xYwiUfGaif/DG2pt5I0D7+FE/AWXo+AJYewi6/beu
p7FOdxKbkf36lFYtFBph4vTpH3Dauutxh7Se7pgeC2Rkf6QbGXVp03Py9P1+PzoQ
2PK8S4DBLPrji9ZgwGZwO3XNop7YlP0WrDwktJysVktRbx7/k9fmYkmVBYQNPV9B
2mWo/7R76hkW2jeZ6qlPYLu3r5DgjSJTPykz949mKpJPxymSCoGfph85UJaL+LJg
7t3bSffKcUYa/S2cPvmCCZE9d2f2oTdsCXxqtv3XjhgbyNt+ZQBcDWl6TaUUBG06
H8+BglD5XQXyZ11jKsLRbPl0uISbDA3DpazCls7xGN1Opxxoa/aCj4DaOKUTETsd
PKngnsuDYTwdmaw+afCs6uZ57bDPvM82Kx69NveLZu2G4mqPocqyxKxt92iKF+RR
fAcfFMf4OovJnRFZk5yeQQVRs+YvSp9ulSLNCThGRQyHWTXCuIRBsWqzV0Dz90sW
B609GdfskaqaADWudj+hsogoHYs8n3VwWvte5a8fxlIOuQ61UzFj+14YchBSvRtP
4JvNkYuep/vwj1hjtHALDECJgkRRE518kKO8oKpc5GTRFSItfQp8wnAC99Mb7LtC
8v/BAyTH62/8zXtLz78W2ahMYbDf0EuNmbUF8xKvYbbOGEEaj1D3Upcsxkres4HM
lBEbyFgnAdFioAJGN2tDIlGehC5qG6SOWegNhzKp/XRSwP1h/9RFoQHgflNKMg8J
/sg22sU9CjR5yJpCjn+DGe/BwwyTpTntdP4NOWdIcP/vMWNGzm4MIhIGo84kJtFl
FL1TOpAL8YVuwRJ8ovjNF/cDuOZCB4pEaPJIJJ+iip/hxTCz4dIkFuREHJecmfm3
mHBDG/Km9td0oX9hkMvp7wa3hAZwjXiC2TcepZv8UvMcjSGAIGps1NOVgGRK3OA5
alPnUEq0KLYuAxKagEToLwZUhdYS5remeLyZt8GQ8JD04eu7SYaCm6lTNUU4SUeS
FKR/6Q45VhfYDSwtoqXh+ellGFzfsp/q2E0lVGcSxpwC0yZEFYnUFa5v3GbCtHTK
DtjGnSrdorg0ohE0DA5FqCKLuXnyKMAa8VeoqrkrEPklPEmupukEGC7RhNZUmD4u
+kc319BIyAkOJc0VvVYyntoec9AYHxpTdNJB1mqVwJBd7fi2oQ09FIfX6NAFmM8X
q8mCTMJpLyLpTbHP0fXpdtcbwx1jDiYUsl8UgzP1pdbsOdsnxFPxX0+kpv3E11VD
Wm1FzrIHlCrgIQIN6kK5iBuFSFrUBowI70/+iUkRA7fy3RUOlSO1gHCBj2CmqMwD
I1iYOVkh3TBffT42k1CYxP701hzKS0TTn2zSl7Chhjo+n8c0cVGsunCfFGH4pDTd
nHxchcgeRyg8t+Leqqqb5FGne4Li+yYVIdSdyavuffD8B2nA45lUM0Abe7IgByft
uTc23EbPDC826yIw72gZhlBnk6h3uAoTeQcXTQZ53L5/ROYnZ46Wu9dbMjsCR9f/
nD4xf8u1bkVIcwfKgOvDx8hLoFRFIIpo8aY6Mqkm79j9vzja6pU3JD+CN86wza8f
0QOp99b7mbkJn+s+VqGYbclrBG6oHY+cnY3FdqvwFeU0UtufG5MXyNr0fBr5TzFd
oPATXtUMUe6vR2zReGjJJv5QGvCnrBqnlMut7xht09Sjrh7URj5EEzrcy9mUI2cZ
wz66tR/LRV9iAz3D9CXpKHGP3hI3qo09HiV5I8p25/ejIudbNt1t7z4+pHsoygaq
xnfH1uLUbQBvIUyztch1/TI/v9pU2+8PzLk+CVuDBYj+8QDQPLxqkpZ93j/ARWbe
kS65EIaRX43kCfWSKUNrkN9Ni0CJn9vVkAYXfUVVj+uuzHe+eW28LyWWzJcy9AhG
5BEsFPYSoQI8ZfQGPd4PxVVSHbX40NqQTw+WaCB4DEAqPcMG9uFe7mzTln43rKc0
/N3vT+qYFp0OZecqY08I3HMU+i3Pz4OLJIMZ3c0bwqcPH/UY80kWncxUJYz1DUvA
hykR1dGT4vOQvbl/SfmRwbrDQ265ML0eZO5PfTpGQNm2mVm8C0W/b6BzrEWJ7F2b
G8nPl74Cu4f3OEPmv24VsxvYEQ4GedKcyNZXulDcu6fYKidM3hx21JaPM7V5rkoD
ifTNO1dZuj+oAvo+g+Pnr7Xmd//3nBnKGpAulmlMr+6yqhq1FpRs9sEGDkLn8jv1
hc2r7TbarJv+uacplcYAUiM2ZgSzGyljMdFDSys79FEl8wt7DBIvs/70vu1RRmiS
zM1Gk38/+iA89Sc+WgNr3GbXYmInabaqsL7UPVRo9IUtC9Xo/mdkZLLXMkL11idL
vvO5ujIcEItqNjgnwh8KmzG2Eyv7OhxNizSMbAFwyWA4AeTDX1JzYZHElUHP091q
QGDDHMrmWEhLfTN5Oom2DzyjRlTIUqOEesS5oWs5RxJgfUi6UAxjORchh+R8WGuO
9zllMuDCl0f+WldELp+M4Cieo1xTODCALCG9EbLzLenephFbcNk2x9Om4a+zOYwJ
J65/Al1POZFJlIZmN43aTzFBNP4GQKWK5kYPd5K3lc1fK6PHeGhmyqFzmnW9HDxt
5rpxYz96Ojyvv59qbwAhuRZIwzxLK5RlWVt48Oga706F+zPqitAG3PIqrHLJW8vL
qoikfUzBF/DhLHAOWfCE07po7WfVIbLLz3TUYyD2wyxRdzPaV5/sD+HuFx7O422w
eC0I7mgKp2WSuu3C4tfDITr2bHi6AVttxVu1v2IMEuqe4DKxpH1M2wavZjV25u1o
zGW5ykIQ3BCXvxmMEITZbmSskHdrPGdvqj2U8vmGkzDIpkzMGL67y5LLS89F7xJ9
gCFXCDzFfluIf8u/Vvnbjj0UO3lrCBO3blMB3GjzhA++HzMp3YovJvPycMgpJhgi
UYsb3oLH5FKhoOOYTOq+xjz2cSVHgUCctgxCmIeT6F5BBUDYS3NVKsOpP3B4AlCg
eEr3bTOZWP6RErbCTC6zf/ZHD+gWMT5NVxHwdFRFNg9oInWNPlK8Z7dYViBFUDZj
JNO/E+tqeW40e3tbnIIpI5+P5s0aoXq9kTsexJKytFSgLOr3diMyyDAwcpjcFGmG
6ke0PY+04PzZsxNAwipGUr+LfgoBRHqZWKdIGlPgU4ASb3T4jtTQa1/rAf3J2zOf
BJ1+Gn7WwfKRvhI8ctN4jsmf5l1xQ5VxZzX4vl13FaNClG+dhu+34b5i1ffD2cVf
lNwqyHJkh3RAO1wLt2Wct15jdTiG7/acPGvPN3qgZR3g/YpcPUUkRKwaRgGVH1Da
ZlwrdVNTnxhf45ja4p/HcbW3WfBhjdQT0cSj8b+kugFnttXe9wgMXNYtsSO6tfb3
oJ6Jl7CeUaqCUnOzZNIa3DjO4l10IOaxc28GzI8x1k0b9wDtHAEKZQjXAlbKI9+p
mgL2grp6fkDCMvE2vVDw8O10mXje+a6IiPvdgdJs4l7dH0k6G4Il5tKI6DJoEfCI
GFatJ8H6CFyyVA7MgRWQon63z6SJQuRNfL4ks9EGl3PYG2P/3YaL210IrSSJAoux
atdkS2R6sGR1+iyPeAtVRdu5C4x+aNmQm3DtZ3Ase9UZIJiWmti/xMaUiQDjDtXf
n6JFtWSx90zZYbIOo8ebYpUMDyGjYcDQE0AGJDNfaV1UpP3RhVwbq2JLJqvwjHT2
nn17yn4RdYbgWmtiDJgK4+1zh+pfBmFvq86szQIoCbGQm0MhcvgijJqHqLeA0ExE
nlQwTGdgv3B68sCmMOqV5tRxJ7Ne2h/V17KvdmwS0uJcyj8Zax7BiAbe44ipztC4
LPbSMjl4ix9mub/OnNBWWN3K3XXheTEIAJOfYvqZyX0/67ns8LKO4iAp00dFxIKr
Rc/jPRUrhrRaUl7cyWnUg8D+jS+w5KXmKHZDhZbXhadCfPxVBZQewsjMaqSy6YOS
U2EWPVj6o5NY1DZsDXYK06hzJWFf9V4p1da2T55J0TzfaTy/RKJC3IX47QdcGLYO
idm2OOIiZnwrrM7JzX4ueh0dthWC+3iV2GUcljwKY4WANn18x9Dej3NDaWkI9dLn
EVmLZ+gbCRXfMOvQKdoU6iCx0+oQQiHYkcs/h5DYRQvvYMpxnmELjX5WtWHkMRVj
OmHJ3A0w3hnuPWZF77VccZI3UGKUYq2oppXgpwZzwj9h741hTCOcfwbMo1vCNvin
4wDjiNOCeJIzV7YhxIOB9agoW2/0Vze+brNZ9BSEi+NKJOeEranVE7uyRZGeRgDf
jSIHjlCHBdXzoYnzwq6vVhqm3t05BxZzthkAd3kqBGBoK7VVDq9tKCqr+cT1FXh4
ym8WLoIT6xRsMoYEk8ski/hslbhd5pF5IVysFCIiBPlcUFnvcBy5nbyTwIWRsml+
JhA28r1CPTLwLiPwjLd5Oz1pxT6u4oOSWKf5eIOpajjM5P6E1k2DCoyHd1Kad9kf
ntn/Kh3FFXorhJ4emIBZwz26Svb1aG0Ue5Yl2j7NSE2w6zxPNNmnYrJtDTbqOuGJ
dsi1SK+64o8xXz7D6V8XSPmK8lXpt2kqNF6NwPWajVN0jTLzxcVk8DHqB/Fm8F39
S459op61XrKLm5VirzQWCTzwYMjk/4rWZL7aN4SfXt3vX93OCag8tD1GhOa53xh0
6c4UcEYw9D2yroD5sk2669Lz66SiCbV4qgIlzMEifbbROkpcTWFCHt6OUEv1QKne
PK0QCGftJGJjqhmYJ8VXrLp2mx1Rz5Ume46zh+kgglEzY1jJwj9R3RfMOQyDZLts
O0ixZyzj1BGpy5ozycD+eOJzZPkOGaP1Nkn9pl0X+1g1SzxgdVX0CsKbMNODiMiR
15H2P05mjPnM63kolooXBRtNSSC4nS9ElvIwR2jnrCYo36yAb881nUdATBX3icoH
cMxpglsSJyd1G0e5lXc3K9KsKOWq6mj12hGxMmLfZmHA4WAawaX52E0VDLVO5WyE
22bEf12mT+fusqLwyUlY5FX38vj1f03hrwr/t1at6EmtXQxnx8zFrXPDr9DiXkID
lfxjscwrB9itZ4rTt4THMAT/IHLywafNu3igj1kQS/WhRMlzPEn3DyZIzmN753I8
bgZllc1dzCeIpdkX4yN2zfIsJXvSVOaIz0p1FUpZimM/H5iJas46avOCyZVizfqK
74/pfqZOL9rvwXcjlsgpkYsMqKsepwvAlGTKfTNCGzIOyAIFEurqoEykQespQkh4
gUM9WbPg6t1W8y+joU33dZzJq+o6aTdnV+bQIqCp4Nuk2X3AjxsAf7yoKaQnA+en
jFLD0DAo+mNgDCYKUydWY4Zx+LFcIHerIwiMhEyVLqBGhL6xoO5Xo/owKNOwazhM
yozru/7maTQN8yNAWGrdqXLNc/H0Imq5dj5LW3Dtv76RdBboa20DzQDGJS1h3vh4
9T8HUDF73PkSS7N/5mR8jaItqQHhnlKsROeWpVkQbvzdyic8GVpxFMRGpJufGe59
B8rTFi/d8P3uCTnSydrX1n4Xb0P6NhWtX/bjaENsEV86TaPEWo90Mq6Rv0PcSDFv
wOEMdKwdWCwJxyWaQOyn/GZLrZoBQb0zRIT2QTipxuaAa3fRGYosqiMpeljq35/y
j8YA2ZeZAuwb5Z6H9NyIIb4gzb6Nqneuj8AVUpCm4iY533d+oPSrFifw608kWACO
U09+3oPwESet8SqrpPzxxIRqnJl+JNvh6B2bpvygSBNIkFGIrcsIgkCkcDLNXQ3N
E8+TPj6jGMEIQbxxJwf/UFyccGgnAujgu1BYAvbdkWSfqBlozTemL4XObDM5G6Ma
WUL+aCMD1/7voBkzeC8RLrqh8V+raI5wjRyViU4VT9zxu7Wd7wEgGxa/N2vCdZ4t
Bgqk59movGheGvAbrXjMOnwClhGXQuST7RtlwyfpKmbvGjk9sN878r/8axKTa/cw
wnYtSSB5BXyLr1Egpbb1ltV3cqcLNO3QZ3R8QHx7FObnd/AsQTBgVe+UXPIoVjfe
IgLnIU4ooITu5AK6D15xu6dSwCWjBbV+YNupHG1mpIp5bllTSpSTwVS1qky1uQmj
WZcDlicLsqJ8NroH2QAq8T862XrbQuhhMzBdem+AlmXro7Ns457Gc2y7KFQSKQqY
Ds66yUvchoTqsyr3v8BDLdaka47SDHfP90IW3D43+CGnyMSq5XtkezKur0Ikx3WW
W8lwU6ijyNpmKq8qtVbP2WsT0inDWOSZIBfvP2wMNep5p5P/BLacd0psxmf1/U9v
qsc66eWRd2qaIqjL2/rHNXV7ww8iV8sj/KEiBFc4XV5tpj03AJv7VfSm6+58FC0W
jQaTZJvDeGOD+hR5rizyFofX5+4ytKJt63eUBF8Q2XlOxNxyOVNQyJfdyV3uFOUY
LagE621JHLxJB2QKqsloHzr1p/y4Cz5t+Z1xO5vehhbM78ARCFIRl1FGUNfITKnk
14uHGnO6B+feXfjuKhWZGPlmew2UQQLEyceAC4cn861sC3lLctUmvKglPV9QmS+Q
P4O3S6aBWM78fO68/08Gd/BSdOXypIFOjHr1Kall3foJ22jkJ4KAgv8x263expPZ
6zWUNxPjZS40W2aKRZLNIT+cHxDRGU6e85sNrQo8qDAv9YP7H7xtjkjKGVhjwsf6
I4VFsd+XVLOJ7IEz/h+H0x/NmIbh6V2ztUSIy+7FJAPL/O54ZAthNWxGnDglk7G/
Or29fDiW2TI22l/kV3z/g7trweM+p3+NwHZFHHJJjkr6E2rczkEnZCKFivFLXKmL
CRIGoB0WYD75cyL/GGFrf1jWZ/mPgfQ8kki4FKkEr2rSUHpAJseKdFfxeuJHSevP
g8g1x8wfd+gMo4dr09J4SX1PcFJPx/UmLAR6TdLmKLPLhXuNxQsOzgVtI0bV0cTe
1eqhwVEnhkHnxfFPsWrvrAUHfA3yxbl4gLC4MTra8pxL7SDc2HSMKlSzFpoJsbLO
imeo4WVVzLVijdtep6fiCgnNPpS2Pqxdg/m9SCdx78iOq+EWkOfOJlpaKYPC7+tG
B/iZZEUfg3TtkyqPBUofQNGl+Vc8no7S7n/NCJFhBaBRpsdtmTRMQWZ9kz8/MGVg
js3CMNBiuSUwpP40Zyx4ZZzkezJernkvVLYg652oX/2w2fp0hmLCYyuA8+bXMnZd
T8YbDuhmTQuStp7dOGHWt0oFNCThAljW6aT3hOXNVpFUKupg2c7qcWG8vLSqSScu
Oafoa96NWnhvjc6vqj8+P7TgcqrChogrbmQJ0+U6n0D2sq14tkeZXi96rrOyBuGl
b1T5mPGmYqXFiOaaZEcWw6yWSQfpb5t0iVdwVmhmPlUDXDrxLFoBPeej3x6Rqpat
sRTW0Hm7PfImJYuo9qY8BmP7DE+D6SwRSX4VN4WQ/4/k2f0JXAjp1ttVez+p1XDd
gG4Te3FWSbKAuyCaplBaZ0I9bjJhQ1CPCdJsZp1JIkvETZQAWqI5SVi/TTH3t3id
wEVrazN+beHHceu5ZNxmvXE2X1xZ1ZhRZcia9L9D/FGxRmlvwJ2mo5aMSbguzeRj
+KyrKYNg3so7Ldge+X/kbK8JRqnJatXh655bUveD/qqbZfk9tIjUpxY+/ADfNnM1
l2FSkKFafOXGx91274ZmpK9XJMb//Q8mHwQN5DsWNq7pvoh2LVFRVeiHW8pYBwD2
8PpLjKzGhnsxar0zYEL9WzBaYJD5qSD3sHeapOqc5b8rPzOGZmL7CzVW4IlJrsAD
cBJthpY0zoX455zJri19o7URhY7ouAjwMgmUQhT1g2sKpPZ/nnARnSfYdqSiEj30
c3sqdez8uB2D+LnZSQt/5OBGN/6cCeN5Y8BTkUh0hFYHJW3xqtZA67xaYW7p7lEi
agskpo4turqvjIouXxFGY2vfztOZphDpOenrOsAAzLQO4yKfveEs2Yi7Gy2gALGZ
wVUKkCkzjn5dPOWajFl7E14pGZ54pPO8cQEduPhiKVF1tXvUSPQ7mDLgozogCdJe
QqZakgo1ozd583emvF0lFVES6BesaW5DtqH+Ighl7iGPpEOO96wD4HfZAcOa2+az
LlecJxuryfv+oSUIVZshFA/JxD44GoLirCPYnetN0mVnWKjATqrSfoxudvngyk7B
uirer8GeN0BrYsF5EhaRc1yzAdkKo16z4j1kFeORxyhYnCyWXpbLCaqQKlabBzUY
mYPp9cQw39EJ3WeSzPP1WKt9NT3HiuqICnv/ObgRl43a13XD+AMI8RKTGsr9iwf4
UoGMQts3aCp1cLWi+w5Mm9aKVb53o4gEcJkCSLZ4fUros/iy2qQr8C3MYkNi2rxk
FUUwsxxg/IaW/8WmVYNO0MZU/XeyBAGaEXIFmPIGn6YcMWTPCYHAGtJjlKAmEC3C
2bU/jxhQKN7/K5tklCGRYf/tTaoi0jGm7RY+gNw+Ss5laM7NlSC7t+jX7KhDKHur
HP6JlMQJMJ+tOWXfsUL26RzaV4mLECM8AAxt1sp3r58xQL6qin3RJbWtRIX9nsuy
Xb7RzWgjJMxSne8DbLj1wUWDguE5MruAsJMEeKO2nyG6TORrNsXORxcSi4nRjjDR
rFWp32HiUfl64L5J8yQ9qO8O/nZ7mneS/hD1pwhncYPSjRnEuiiPUyHA3jDu1Wz/
hMknCYtdfP0gTAqnUk0ByexdTS5rtJ3rVKRivKi/sQPuWTRLDRp2K0Vd5n6fWRUb
5v1G7rhpexfAbVAc95sd2RMUq52JTgTtQiAhG1sQ08k/M1RSIPSXkmJT0D7MhHKJ
q3hxNMypSqa6TRNdNSA/FjxL9jqWYqtzf09xFwyKKQPYCKLt+vkINqLNOGPeWsKa
IyZZN9SBPCm5k/94GFOKwPu7EBiFpa/dMBpJu0i8LqHjbEm8a6z4tGxN36ZvbWOi
gH05+Bjgy7LzOx0TEpTa1f1RdpUY++pI8iR1kn+Z8STkuuriDbeJHJdRzHTwmvb5
x908TDDiSw3om7azNEvF2mMf2fWBqDX7zSIZ0TNsSVQvIviedMHhb6d/9I0crKKN
3+apkNvaR/aeKnzlyz925rbnO04pIt4yw9aJs9bqHx5yEbFRFFLu34grSIZ+vjEh
CxaHcS2hzsaN3avKGpZzd0pS/dUAwPD/KZ4r9A3udpfhRILkxvFSPzTwR2XU8+Ge
I9cd80REcULNGFY27Cl6ZuVSIzpD0rmaZvN/MKMJyb4RiVJ+ofIHeoZ7dpWmZyhq
MBpaxsu+rCj150wBryct8q1E16l89M92GH0Av7fZCOrzIm7QI85k2KyfKid5hO3o
PAb1dwzAzYXSwTtVvXJwTf/Iio/NMCN7RVVFGqc22h73Al9FIXgyL2N+0eGfEISx
sOj+oNxTQdWRvBVWkCkuodZvUjNHbmifX33x5Gva6BSebiQUyqMJIWNBE8bQM0Cq
4PngzB/d/mG4VSJxhbZMByLkOKGKYVZ/Ixp3i2104ctsNzRXpPGbaVvU4upamFvb
a9OsKYS1YoA6yMkvYi4st2mnUE0d4vrZ2I4ZhQY5or1U/PpnnqtFlHXnMpDF3Qr4
LmYflMffsPm+Aany5loNb9W+9KQ5WNbqB3vtk3Jf57qUeueiwdBoH4EJLL9KkRTc
fITwaa/JRXls3VXNQdcpYu43K64way53IgANTpZvHbKdSRcUBbTm/hEpVAji4tYS
VmB+zwqCNdNOks0MAihXZApngOGaY4gGokSJb5c4+Lqy+1Q06cvbk0eeCebe6wVW
e+PigB8IG3Is/mIaHKITTkMPtjo/wvj1SWpj48KADTu8hY0Dve5DQLK44nltENDX
mLHwtvDgKm6oFdC4RAYJcvAdvBb/raSniNJpa6yFZ3uhgcec9iPBClgpTXPqbynh
+fwKwZTasC+osCIovUIoz71TQZMY+HCO4okC45XOmubm5JvJqPMWETonUmt1JCmA
jplpQ3yRwVqfLwcqWu1GXUdbY4BIPRwt7Xoamr9lOCowvEomMdqEtUjB11u9DPYn
SYkEx6XqQmwfB+ciieZHGu8m0wDPJz0zCbNL4tOwFNEGXvuJYLYAKrELHWTghoHs
Msohiwl7WDUV73rVg3KJQxpPYAMNLo0Qp28MK7iX4TTRPhGKwSX1UL9g7Jr7U8Zb
FQK8mfqnEmK0kpBREepoNT0h76eZDvx7an0KbKREEWWuKcTwpSpAuWH7eIYv63zL
P1QNpW60znRhVvKaaIElQGMk7prtfEYGonq0WABM3JJzyjpe3uNmG5A37zQqa5HX
rclM+hV2y8Rv1PfXAtIu+oHv4DCJV+Tj0IuDVLObZZASDPMMOgPAVojsSROxkElz
CyCybiYgOA5gexJaSzgF0J2kg22TYHRdDAr5M61FkEG+Naw0NJIXtfQjNdKnsDvp
/efqi6UsywqVtCFHVTieAQt7qVnDbG21sWdNYq3rXT4DzKFF7RZtgM4Exsl2LGaa
4YiJFvMkoUrsOT7j7KQ9XAKSAW2csv8k0+3VHAq+B93J/9RIOIG8vgwh/xazOiz5
W2d2Y4m0QQ6+0QklQPsTejMaqGzlwgp/Lq4wpHwrxw5L5fmlugEYieUR+P8CuFTi
1TZxBgflA887pMUqM+mRmKrP48Ab6PYZOCrYCVh29VwE3Mp+CB05FpTN1U4gygZ7
v3ajeeo+/uyRIoSDcPlClXR7AE+/k4Kul69VecWvNcoPfqubIOMB45BB6b5JsXB6
svMuIsDLV34A85RqrRI+O4dQAMMVu4xwKSvajkAvJpTfTSRFk3qDk9mj0HLIZm4p
vUf3JlPTeA0oF4t1hFVtwY3coGMWHnbmBg+3iTB2MFhStc3+vQq/AwY2rqstxhEN
PrPr5zEiw+T1LH27KgDGGMAlo4rnVbQjEXZnt8hsb6wS4THywEX+uO5NO/OKcLDn
CJ+f1Ol30lvorVju/gwxKl7Y68+/cLSpeWV3aQUU7BuvkDixkVMcApn0N0uraUlW
I4b+MHG5jo/SA3CfAl6fnbsAuD+Sy+78V2P5c/1l9m2cerWamRafWm9a+kCW4Y1V
cVuiYcZl6IwRlFzGo0P3dfPUtoLRW90W8pgcCv1g4Ti5sOjkbcRC99TZsA1abyoO
gPbyQqTQhOUaPZzvr17O29xUHEu4H/wbY2VCuoJz/C7gLBUK9z6dcvI/ZG7KwM33
P9IhGrblOBkRqW5faGXzbywkfcmmV4jQ5PlIvfzjvInIX6pstRmc6lRTNMuazFpM
AiMGt7EdjKWYIqfct6Ldy7dV0WdiCSm/tCcRVYpKNyu3yWVUjJtr6SYS/pGCgSZO
oYpUpnxKiH2ZOgg636IIq9yUByYSYwHCoYPRwGSC2YXkOSMZU0JmHH8YGZdMMBsA
qJhU0hgNSKR9aRKNFiVnuGfJETq/upe4qMJV0vMHxeGbViH687IjiLceSe0QHQr6
SH6WQXELjc/3oCsOxd+FQ/Q8lEtcg+2btykYAPb4p3DiPbMoxLI6aKmXsNL+cfmH
ysIxiA/4flhmiC1cG/caobieG8DsKKbECYgFpbSA9h2rJbI2nCw+Jvp0jADMsHp8
mhQXqBddiKsrWVhxCLIr34pAwrt5sBN7yUI5exoYcMJpXTYLrZ0SermgYn9jZBOw
MdM8+oFG/WzLaojYuTAGHVmLk9c8J8pLFvlrlGZrAaefcGYTT1g544wfLREUnBBh
Rne6SjdvzW9igBmtZFaolCJFRGw9fNmvGA+rO//gBnuhNdG2vETgXPbqiG1DGj0H
lB7eI6etQG2P3tTpsaqXreVBjuDr5+VazVuJkcDdL4r3e4kgUKc+5LOaHiZ+5TX+
Og9UtgvBAYaBIvd16a3riHOXpiZPPlZ8N5AJzsEjzObvtpatEQDWVsl2RRDv+JZ2
RPWA0CqxrA0KJRw1CuRi2C28VKCvjCaYcdD5iVjJG+YabBkCjNgivqauQG3bJNCt
drR3BkfhngKlTV076tqiOIiZo7TqYdcR4ICwC1dZt22VUHjDrzU1PTSOHO/J50VM
UPxouDsh8PpG3m+s5W5ctv5Zcvcndiv+wSZcMgFcFZIvaWjHUedxMJfwNRNkXCuN
Ck5o3MJViO3h26xCSBXMcozQ/jAV7tXKPm0AOQ5TScMwgnfaUKCsZQr0d9mpLDEf
/6fF9hYtvQ6KWQf5dxq0wb3mAo1moQSwqxK7qYIhR3JShAnqSiXkLIEc81RVHk8X
RA35frCgQBnTDFHnIMqpu00rcHIBL9utM3mAeEz5hcz6PNOKMbbUaXOy+qVXzUyD
qJbjt97CpUOELjzZCL5WCU/5rs2Rqa1YqyQfMU+sTWxuaIPt1RCdpk86Yxs3S4PM
e3/mcWsfen4Huk3RAO9pYg61xpymtIWRz6jp6uL90nQ74+Py9lLaZPzZ9ASJcp2m
4BYP7zIdwn1d47EBH2hayK2WKccNh2IerdVzyy716wy0fA9Rs97RA1qDsRN5ExCc
cul+p0r+XchpZdNUzWWEw3njVlRxLY40gJ7Ei05BbCG+Kw9+tCULCgEmcZu41YIs
JrxDH30qHpNkH8HJdYiVRtoVyA5iI67zWr1QZsp8P7hqg++GsQlisQA1TCC+Rpas
seN1H+wh94GuHA9fBHolMJEfIwfSpCTtaCNftf/VTtzSZ6RTUEj0YZ8XdchyokVy
pWsHGTwam51BJktPDcqVvBJe8HZ7BdXg+3mQRRo8SaGBe6CFZ/JEANjKYpu9d7rt
J6ChrkZeL5Qest+EfueOO68SIBfUlemgp44eAPA9a+10+HVWtHIM6hUFq1bmALcF
05Cp1sZsbU3hCoUHM5CgRMm3bac49mB/GNN1w4aYZ4Z6uSXsxKSjcs7DhneBdP9u
2qbVimg1dk/39enmBw6PePkwZOmsTjGD/zgQqsG2SzZXnytR8N78vZkS9n23JHPj
NvPZ8uQUAAri3C0VAhmrujwuJRJnlwQeGRF70vr52f7JApoOZjbtrNQ+VFEAWL8y
Qt4beJSb6IM8U5ADdzROiNPkO3dGXKSudpvG9fLmVWce/NiEP2ifmutT6tylWDeI
b95pvsGqSLtIYvLp3ec9eWDR9ys9m2zFQxGetGp/D4/eNgyemPkRlebXGOSHjldW
BcjiVXiPX0SrEz0jcTPnIOoBvMhJSp9kGiQ1IhawDcI=
`protect end_protected