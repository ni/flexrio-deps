`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 29664 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
FTGcP7VlpSOhasofAJvqcAPB3wm79aNDA2CysYS+mIpVx1fTxhDi/UU9njHfeimW
MgEKkkf6+CE/PY+7pUKIEZIIxZIIU5fPzo0qye5wK6HlKz8AgnR6ZcmaNf1cZQsl
SJpNZmI7f+ydRHzWeja/2aRZqYLOMgk6ZQLa6CGQ9o++raL5LjB/PYPY5IhDSxsz
bUbEyeE5Z+xpUnQ8cK3UR0FoWQJsTtXHZkhiyoXkfqwxW892L9Zd0OaGtjDuBQTF
uAWY476b8TiBkLB/XE8TqZkZra0q0xXrpvH+6n2eys2hNzJ2E1JCbbxk42p2FPtz
w9VofRhFT9EMBBdjgy0pSXXS5uF1tAsNHt84cSaahZYDIzWDcMMMrmX5nP0oCAY/
46ou9WAPQqlZ0GWDj0n5xLa1K801m+GosF5ycU/LRyllQQ9hmDA8RpiEk64bLahX
0uqIBDmhrBcuSIR8+wdkBw1zBl80wNA4VChWh4S7D6gIAegR4KrDrz3LopK89aKi
yenHl2vT9kh5hxEutLPpvWLsHdWuMJlRhxopvq5BhTDPtN9VcAbDCLDut8hUuhnV
QEQVIm72lsXcgA55gpp15HUKfJhPmVfSy/7VB09as7tfQl2RQVS9jdOGVXfpUh8C
PV/i2PyM580xVouD093OZx3HrbHFq+mVBnhQThIHwb9wb0Ks9tlZY7as1Mq2DBD9
JKU3DqqlbSAmueakgcNuD5caDeA+QH8ZYtB5ha+aVEdStBMGrZxaeCYCANyVWmzn
WSicffUYojhvgeZzhR3ay+UU4or7hv81N1p9V+d+nPiub0BU+zB21iMQHz2+3FYJ
+2ZE7NiONETIKs7HiBpGOHSnsKFz+GHX9r2zMeXUeWBkuSNcsbZOAyJueLqsAhOQ
fVmkyBMBQ1f4jlyPXpS7HOeHpwGGNWLerXr6V5d9ni+6JeJQwu+BHyv4sCMsWHyo
A7HITAFstSqn+1qigj9wtJeuP6qmfxy5JK+iWS4UenzhfOWCk1P4BblUqjMjXYaW
E92o6dvbo19jmZFQly49b4C9+eQnvJqY5R+XQVdyyS5FmHXcZeSXYZvKtsK5hY1j
hLHl9q1HN5yqkp/NX7jHhLKuwTKwUaok84Gts0v5E7aqfXXxUOQS6y8+OT1qJdWg
VrqNTggEOSbgFp1/euP2DzdKaDO0PqWUyJX0WJMgEk13LC0u+JN3CfIE6oErdTEA
o/5XfFzE7+ba6WICCSKHdiAaQUfGGg/aScymg2JPdRZNW8yXvVbwaUXosHOmGvOs
dVGSPUHZHjdzoCpH2J3wOjJXQ1BoYeTXpEu8+gfuWKEY9enoXqC2RTWx9+ydZNpU
2N2JwXeTAz8qdEeEYaT3D9MD/Wz9DohVqvqejaZ0mtMcdZVYGV93kSvAGcCwfUIg
1saUjvjKaaU+Q/qBYLUZytQFnsxPhGBtTFkxtsJEXtlLz0XofBSi8wuYG+N3tckV
evzGRKU0FY2Iy2tCOWCNsSm1eraBJldpp5bP80ScKEkGrntSxA6YYN51wxlEwWgM
hYbKuxlahEbjBOQf9GYWJeJbpnlCQ/UWTNQnPeJeSelG4fc8p2ok55qHow8i3dbd
L+TWeMZLhMwAr3hK6VrGidXmSRpiOGNzvLt5ALTdg05dUWnpMP6Q6kEXiOA497rl
O+Z1a92R6tTVkZdNaejIKsA+ig12aNn+2D1yCXsglKyHz8uX7d8dRUfWjgM61563
FHKAIWAgETNURU067BBwSqQU0ajaBo2DdlZO2mPqPyO/XTRmbxerHhCc5Sb2Rj1Q
hdFmXoIPSqT1tl7tTT868LZiKPs8Fdj/gDJ92Ikzl7EkBpJLesXJYxdZ1DKlMTf5
+9fFTlpBl2FXmjhB662O9tpm5FqKE/aKY+bNZcfdoQe/yk5kBZ+C09Aer36RLP+E
kGfDE/aNtG1begKaZYCZMTsXERcaL4m4aQTNSKyIrVQiOAQ7QiiCxYBYXfkyUh2F
Ut7+2BZylsTiiQCGJ17+K3qaZOSZKFSdmYU39Haa/Lovx1SmGRcZTZOxFgIFZys2
6oWY+WtYZ+uuTDqn/wudr6gIQNlyyVhuteLukug/S+FR/4KGBwBe5M9KXNsFk4Pl
IVMjKm+8hZBL5jDF8sgilqSgCPbH9Xfk3bLAQeglD/G4qDxBDvPrIHjpxnLNH+O7
5+rgYQUdOpttvjG7mMNGWmY52KqXkVBuiLG6FpYzmFRPPPSfp4/ix+rYlWXpXrku
X3m0OGSS0SWtkHzmdUJcPVVsSzpVBYO2n6eRqcEMx+KJefNvKaNLbZQi6jmBb8Kr
TngECWSqF8ke+GIuDisE6Y6Ua1rcEVEsns7P5F4wfJnvW1fOZT/Y7cOY67yOeTz9
Svo8DeMgLwv6WetLT2A/yE6KCLHSwyXARvu/cAXyfU/1L2O6GcnH4DO8PYTV5Oyi
nJvKUX638U8W9B6fDT377ZB9hh59WNbU8cGezFZRq+N4lMnzR8B7iXYE8lQ3N770
v4Z7JJzRg4vriwbThjUzJFcNg1XpvgGVA81PuQUjE2FbP0qdbo5Kbb1MKknXC5uG
EI4TWUiKkkH3DESFWt28xi+1U5NS11+kg54KBW2xbEYSCgLd23GuFzOZD5SWTYHF
t3k5M6GLT1LF2/Xo+Th8nxJKWLI7DQ4SRTRgT7h855tGxHbL4MFROJeTyGbxR3K5
QyXrF7HzhPjHUTVBh3wm59Wzcexpk1m8tZY7of/amBabziZ3xR3F98U8c8PVD9zz
YFaWPlxjA2/w+ujs9CzCTF0W1A45NbRxkjQz4kSngtW50pBH6uFrRHuYpeWvpILg
qtNztzN14j+9Yn8WC5oLAOPKiLrfTi/BDl1j/+nh7FBUVYJwy/TVwDaJA2ndpngX
xnXCnymmXQlRvXEHUjDI5stZr6/jBeEx4JYeuj2N/qiS7C2jtJnc6wUXecOK1bHO
rtYJTmzseGjCwegRTTvNOLdiNPaJvb4p8lokGLmjS2+qEgtLD4JLU/WvikCM07lG
xJc2wk3HmcMC90OR97zEdTOTX+0pIoiGA1eRJQLbFaBZOSBlY29jqOVBuTPWgufe
xPJo+1mg28iR4th3uM56WoKUOmPUQr9ymE94r/axtIEVuoYQS0PmpEBNhUXpgPjC
myHe9WRXJ8KGs3WncWJDslL208564UY0BBHP7+cQEDlhjT/VVbY9t2rabCLCkI75
Fir9z8153Gr+3ZFdldrAd3KshlJXeJSdbvqOO1bQShgzAryQhb6xCXfSMx4U2yWL
toymLxLgfNRk/wyIGI3s+IUJMQ6VGHHHRF9EvN1D07FHst3p/mDfKBu8WdOtVpPN
b7AXf1vgoDAUqd74P3zw6SYeqEF/5wlkjqotnBS7Zq5+2l9C7mBStB2z8X6hVZhM
6FAVVaE6OzpJS9H0Td57nuvR2GUWEP/P+tK6y8IBH7IS/txYWQpAy+aCUzfDi2NW
w1u39AH1dyoxeZ2/6xsCjEYe8BDrowayI0fkuUs8zXo/00bC03+aElQbIAoSw5qA
BDhBIVLmy6ki9uCD9UJ4w1XFmNmNyMinuDB47YtnyHgyC9FTXmczqhkHiPb/nFz+
PxsKPFma4Eibe/HqMct+HlexJgRvoCJk5PlxlleTGYCf4ZVYcuBeQG3Sg3RfrUla
Gwg43DMRVbZ86dH5xQHwydN7XYh1dgpaqiH3r0f27T7udOLN95TcH938BxCzFRHQ
rRJYUmDpZNY2ER5cX6CC+PHsyPZjhE4UPuBaU1W1tqlzpNeL/muvgAd94XBmAF0/
s7ee1XcHagkm/v2QFTT0bNv2Cv3X6hqY7lMPRbnW1lKLKFDAXo+X2cLU2Gf9rSL+
xjfmOUB+kQUvbLg0rjHroccQ6HnjH3skblAk8iiKzYygUi2n9zoaFxxke1wj/RZG
fREOViY0ASfirFCP1NySQjptvslW/IFWpEY8/mW87DKQsKAabeNdHiqU9QfgF6jr
48ZgQZCl+wzkk2+LFBYdcphC3llV1P1aqcFdykONT5vavUgNzjRIzJ/lc5Lf4M/0
nbAh/Qw1XQo09ERqc48yHos/1kY9wx8pg5heas5WaG8ufIHqrp+UNtl6CUF2sGIu
omhi87CSgcOjgfz1/7dx97yV6o9YTN/OnMbaZ3drA8WixxCBWHE0rDBRFhi7LaBd
VFsoy4+fPGwOceiyV7mG4CkLtHiNCf6BtHCMTDrSPyXdFSQD0Qkz9qQ5IAXOh2G9
Ai0DzzJPUsOuzWUsZsRckPeY8r5mEwLgbGfcv4OIsu6AIWNVkjiQOgYj04uyt8aC
UPG5eWfWU0uZZ+qlksz+UPKvHEcMktTfex6DwL7GhgAoQlKVxpuZiphMuqsmRo6f
58UFOPKvlALNoe/n01lvntiE62JWcqp0C7Lup9aM/ThGugUYnLEupKz79EkTpItS
l6mxo702j2KbXv3l8fRKGwPb3OWktfunXtbMUnA1NdhtSS0A1PiSU9SEU+0+Dn0e
dkzYsJRF1BaBCq8hjEPGd3ZS5Hr8kNUo5ERMXjvXwnxMU7r7/hJXNCuOlLDPLVDJ
kfZb/o66r1o0VANHpHDU3jONByi3h2z3mguoRQSmT4glooSkOV2lLxxme7epaMsD
F5zvxmixsFH56DZplBMXnweJ0H67E0TlqnYH1Ju4tt2nkxhbYkgsO3M9bSwqda1i
h3XMy3/e/5V63znXsFyFyXcP3Jftf9UGwQOCRgeI7Xg9TYyfJtiY69CDTPh/l/xQ
OQi9zXrT/jqk9kvF+fBApTo2pnS6WO8QsBL4LA4Y15jlSwrXBFKUpL/cSQFAc+m5
kocA2JtAPCizCBSSMDCpl7jJPFTyVEGzJyEvjCMn6QEGyMwh9Cr9iVZEFDl8hDl7
fkXGbB1PSUmVK3n81Hf3o7mg3TbKirMprrT3J61hdOAIxEMJIxl7IZSeZ/N2aQVq
f8IRp3g+0kgMuVggmlyfLd4gGKQDGzxzPjcobqtVO9/sdcFs6gMU4LZidO+Cm6xZ
igbNttr233xAug2R02dy3j8JcW1s6WZECc9MXMo3av19Vofpv0Ob2z20FoT9Jm9c
BQE2+67qAVb0IuXOILSe1neCe6kEY/RrH8UfvEmMBuAsO4/FEmEC2dyA8zFCzpCi
Gj+Fa3Rft9JLkgBryVltzAhpg9LHDhTkAHRVDyLqvtMo9rOEVLh5Jq+kA/m4cDiC
xjjFm+RW3o2KbOdrQANvY28+FSHFCuWV4ozftxcOugsENtUvjnvXHv22uBTHljzb
tQfeVraSZu574FdgE8Ns4RJeByhRv9z9u+b66BVEPRZCwlBfgE/eK3s/QCNRNqnl
Pc0llywLgvqXUbQtZwD+tH7O2zz87MZ4DLI0umKL0rsa6NPCrG+27dJ/fgA/tD/w
dN95J7bJI+vI6yk3nBddtW6sLd/Zjdq6VRUP5tFm8s/bLk2PWIqVjpGFrmoO8/+x
6cZxfUXXR2AoYkPY2ahYl/IRi0noz3uZscH+uODgEvDu3HXwTRMx7+iq8zm3VhcN
yLi4qwj61/Kuv+fsENtQ9Qz+euFTFDVRDXOtS/JwrCufXzhy0+zj059tq1CgMB1G
JwN7USVMiOmijCYGWkY4TJZJvKnZ963nxKfefHWzn+yUf7PBaQqmvcXr4PRBo8yi
WRagBojJwlLeYzVSjDthhADwM9x9su0EXsut5JIo/wgSu4AlpbXYWNSaVdN2bC1j
tLhFZ5X81Qg54EPEuXW5vkwr8QlwVXl0WwMbXXVolMTh3Dym1v87Aa4IENwpD1Vq
HXmJx8qm5sebPHBmCovG+o4FwftchcEjnS/KER8//1upTLXJZ1GL+dMHQerHmbZd
VyXxMLucoAKIbd31jiZkRYKfNw49cfGXFCcYqWdyIZbRCC7HWX4RaTzEiHjf2k9I
aP2ahfAVqZb8nPK+FvNnfP+WV3kTVt6fhb8GMpsHG1Sm0z6LDtKvYa12qtH0yrpb
sFNwiebVIg4NDkcsd3ifXX/v8oYUy/MHlms3J+4ozdMw0iAwPtG8gek3oxtl0AhE
m9nO40m0Im/CJ6bzoA49By8RFM8bnYpZVymcr+hpuCW+x4WA4aFblICQsgdygYxh
xrveA/TFK1Y2CUConVHfb33wiuL9aQ8HodFRciDaBQEQ7fiF3oMpwUt+41s2CEpR
a/A2r2YUJILM+082hElDo0kgJl+q9GsjUIN+4RXCK+knaUgfKvxIk3PnMjLi5YFG
+SM+hcuYGJPas7DVMGaTBcXplU50wrbk0o0muf9+rogp4+2u7s22QBi7veJ5Nwg8
gDuk9PJUHuqs1p1VkP7lFuznC4yiAwRmvfrjdu7z6Th6IQtdyvnLYxHIxNKViQm0
6sCAqfaXlHpbeu/t5r6/ee7LlQSCIil517sxEgjzDQGfUW3SKypY8orp/d8AxApu
MJarOeP/Hgk/DUaGWTAXSF0XLrabzvd+Kjte/FLajoL2y1uUkWBxtYmPpUnW+yxE
RWy/TwC9yb2G7oePOLuANqbs9cd19GiCH5Bl936PICaULr08EKV4gmSbFTUlsgjI
8YQXh9oj6n5a2qVDH3LDWP8WIW/QN9iPnup4pYRgZfLEoGjoWB6opQRbuY75Xffz
lgys1ZjHVRFvy8g4Iz7n4prlKW6e66iCjvSCJ5mk5E3E4VAhIN8BXQcntki12uDR
MlANZpb7TMRdQWG5xj7TWTc0+l+GzIDLL/XA3FZv03Vw6xmqkmfrsF/cH+oIqCj7
J1prwqwbRjm6TU2nJwa9jgBH2QLWD0mMI//cMB+23HjHmE0woFXxkV4jwYqsQoqF
XFexYWJRMufAH5DDbtk/YvTpFaHXX0ZNV3zsrK9Na6b7y6Cijocmkvu8RoJapAPU
CQgv3GdgOM8c1xrC1Whc7quIA4U+VzZ1R9LXmRCTJ2A3n9XZPDnE1tzkz+Wvc96f
l/wdk/l8+AzxEREAN15isGk3HVQwbcdIKHYhrZ0mFt1h9oMyTkbnEXWdV5r3gNSO
hmHl5EnQGrT8NAwXi8ptIUn+r0fNcJagix5a+zSjvJryEXRcTL37qmbYc11BQQa5
fmCCJ7D3akNOZpmz/7L01/s4l64s5qhYSOIKTZT02gJrnino3z2H4uGftTHWbZfk
gGQ5xPCum2wcLbCTWHU7KDuN5zGwC9NeFIQaSH8CDULnY3Qa7nYJcMghhdAqxVbZ
kcNyyNr0Lgm0BxcDTZDQxJ9Uu6JFA0dHIrvzPeb37/ktRef5+NlMmtaCp3i0LnBF
J5pd3OriDAb55+FOenD1/q+pfJZIOFkQ180ci2UZoBnRWz5DB4zfphIJyZsP1j3T
Xu4s1Lx2Yd28reNwj2TIoB8STm2ieRRlMIAtqTCI0A5Dn79nRK0iC6QWm84nqDOX
qZtB8p2FI0NmNH71prtEGPaHxJYbRa49JgnnhgML08oIiKodjn7ZtBikueGVV0Jq
Scs4rYC11NRIx+vAxy2YY17MlbdOV/5H2qkuWV+GmTM/6ZK9KbLXFe8+igka/WV7
9b/g/omXy0z4c/QhVUWvjhaQQEVl/q23UhQw/nBoPVySctkVOnlHqAIDCtU0ZgKv
htqYeIaXi+VIQ+10a5x4tvUMsICL7WHgcYW/Ue3YA5jKjVY00m5JG261/dUwmX2w
aGXjzrhud+JGepL/JowE1KfvvzkZBmhEQQ0xVMl3Xt3qrk+S+GMuk8BvJG7vgvpR
HC+fEhAFC6H/KeniTWIUEvxQIMNInKHB9oAGWC5WjRaosZZtOJmMp4Tu1abc43sZ
+oLzhi8ToD/4o+73vXkkSuxGh3svMNmzDhkGTY0k8wM3iUpayuoIG9e/Sa2vzSmN
3xtSbh5cy4W0Xgfk93qxsWStyYWscaO4vRs69vPNPm/LPWnZ0TaKLXge4sMnO2np
az4Grjmehv9kjt0er5exzGytPArEw+pWdh2gRZnN+dw9bO/qMDWtXZ7a/AYxsj+n
wpuEda/gocvs9uxvVd3poAgCezDxQw0gMjUWYkAGfT9Nk7Iwb/MqOuYqAOZqwnJU
IDxEAwcIT3Y2K7hlCl2Oi8Df4YT4nzWtJfsCgvickZSh/hdyfrPdg6CgpQvCCJon
OkgyA+RyvLtdt8Gs0vVywQ2MPGDuX1y03IMao/788hRYyNv+O6EkQoVyNVgnV8ZD
WBjdzZyCZjeq5rPkhYJV+k0AIWooa/ZTCj+vwK3rI1N+D2TR7hOj0gZMNXTDSCXf
zz4GHmWdXi9CsmkYxksgxSnAZdLNboac4vamXrGZ5/qRM8tcfUAZRK+xfR41S43P
1lcIhuXrQV/Ny7kZSZ1MWtpLadmYwlzSXpTtskTpRJQVgi08i9r5/G0OIHPAYlHZ
mw8nuDUNKSHbW38jyhZEVqyw7U2Ytw06wlhdHqxMvA029nu6Dw42vlmL9OWOsjeD
16Tbq3AnsiX/ADg5D0TCwwpbo/FSGUtDlvKFIh0anYhCbcRaH27ZqNf8WDuXzLGv
/BEMYUEORHMxOjy/f9K3UoffW2oHsL4EMvygrkyZkAMCPDuClMw1BRkpYEoV1dLB
NU9JQ3oVM8nnfikFO/AI3u+kiM8P193AzZMnJ5DruenCZostuMgqgZFiHWfcXzsj
W9wnAREt7kdPs7R9wOxav2k3jg3hcdqy+HbRoz8Ov/oKklzyrFZZl62i8r6KGHyJ
Cox0KdcHKZrSz2k8evStZD5wwdfbp+D5Lh+DNHKIs6eXAJr2cxMOEtyyCG8CTIUq
p/aF0UTtcZdtGA+ouxDvqpdNkwfLwsY/lLrFg0B2jKntgXTvHb3XVpn7UziLq9Su
PeNOa0nny6MdykZaEgQAjbB2wLPSviNsHy9gaJRGLdJSMQddAtzBR7iw0YkRXpPh
rXYhOJOobsml2ASPlgr86PXwEmpKxHAK5UlSp8MYHCdlPq1gxOZWJL3SH4XZ8Ds0
TWmPMh40udqXZJ3NYf+0jumpnYsvsiO2UcR9wyQEK7ZKhGGczVvLac3mnKTZfsv+
YBfCgaTy50e/JmgzBH+kud8lbRHQleTYqBgUBWi6KpoB711h6hXx2eShTXbfKt26
KfbblDV+mK2Uu8ibgvMdiI6yM+9ywK4Pdg5OgG6wBH0f+k/VfJCHb4O9fRDWnwaW
HlZXJoEPyFj0bmOV58LhuVZzJm3LcfQkI7zTeP/oXzG6LVxMO/8Ocpe7Q1JOpIj1
gi73PuuFBJBQdHIY4k1F/dKH86n/ctEwehWG9q1ppNv0xQhlrok54A5hraoZN0Xk
mRSE1es7peV3g4De4ojBYwC3SYryG5sCdBKj2U2uvrhJ5bHLCMz2ztjEk8wPthay
2vGPquoYVHSKDvjHz58XdNPuPLUUZI3DFGBHYeSXpx7TQRAmDkllr1Cn211AdcU7
RDVRCJglgcsk+mWZVqoAN7a3Gg/PdeSSp0EQsZ5WJyZmHY7yZuI3y9wcmARfX15Z
Z8FAkXxK8A/im4USJBuijJxGBQ4COA3SGBLRZ+lGk0Yf7Ty4r/M6tBcIiKB+STw6
j2ezy0HSpoT9Ootr9IiKEtw2WDjVzBL8synRusVTjiykg9KBe3AdN37DtmTF7KO/
vj358PF1zFUEcgCndlDALpPlwYB4ioeU/gqg96NQdlUnezsdlqt6bI0wF+J4cHWt
dhIG7jFNPtHK0kCGAyvjGdOUVHnfJNfw+noR3xxGRb6ZGLp7Kjg6CQ9t6CpUfmlx
PzXHeyxBtCtBsNxNfvA3F3UvPlbQj2sEs6bnTrTok6Y418/wUvTaYPnk11RlYl0o
6obS0STRs7ZC4QTf/PN5OEFTLkdWbpF3PP0+1bLdAY5Cm5XvT95QpS7MwtQZGRsm
Er4HLAlElawnqE3zBr9X5d1Vl+DvH+s2K6kooeUfj4ort3EuS5SAXuJM44kAwolP
cFYmho/K3NsUUCEWm5DVd2cIe+BiS7hGYRHDw197uZ6X99ZW3Q4ZPKnoVdERGtrK
wSbTLchaokyan0kxyHCcWoUc/YY6sHQaGGt2o3Cg6A2vYCFOYnCWdLB3FCsPT3ax
dFWj9P3U1YXr8V+QR1jEFukMyqd0v+S1r6e0hbTeL4BR/c8Lszt4k5P3wmJ0RUOH
p3V9kG11ZnCcpRxHW4ATtxVnFg9dv7rqhFXIcYnRztvq50bh+hFCCOkeSilMEbkb
Q4wowlG2d8ynLvJY7XNwOJ9CzAn1vIYaQwa/AE9JS2FDFTffqF5IH+Y0vvdb6ohR
0FXNkzouK+zAoUXCtrEK39IBuehe5TObRCJO2O33guiStocVjIT5xhFwIpYmz+6f
soHks/272u7iqLNt5qZppXRr/VRcPKQicHHolyxslWmcv7iyUywX1IzMXFoOttsg
2e41F8act8jaTabCa+nFfumL44PZSExLg+k6wpb0HcI6XfV81AROt0TJjuvZKAtM
8lxzdmTkrXXwd47a6XHA0gajZ+xtogbdN8Ih2cocLKjUEfLPbeNdonyhXcIaMGFd
Z5l+KyzlNLKcDF90Vkhxl8JfSyw7q5Y8eN3/K/6cLCD454zsyS5pKDf+Wj3rB7GN
5U7oyjndBIafw9GcDc6Xx1Bex6wZH1hzUvOEG6RzbHVrdruiMMp3LL3CZpId8EHt
m6dU+2i0j+PnwlatDSkRWQWqLG4s4rQSYRq3c8IbaAXH1/zzvAB/yMf9UHzZouWM
SkeSZKTisIEICLjiSgIAHoHxfRFdzdKx2Gzc4erO0xlZ+OxCmoWM7IymugQ+wbVx
sEiR/IKofoTK/4GH+Q41WxM7UIW2xmO5xl6jANO87zNX2HQkc3C7u7ykLc5qwGMv
jUOs0WEL/c/HiPdbovKodCayORrSEkqVYc9tbNq6aSVgTo98VwKfoMYwlWnU+6Tz
HkWBeWulDNE8sMslNNX+VjzpUym+LyCT0c+F1oPv0NEQcCIdOidrzBxRKoj63lcX
sTMEe+FclJGmBWJ6OHBUlz8OPHDwDgR0ZgujnkJN9+zy/mtnZDlmNxNPRjwpl/5U
cJVDxduiXq8Z+1tuskq4TXZPz9/HnRoTHwXqLyNHwkciyB/PH+DpWY3TQJx6wZv4
MChfWDQcdX6CGVhzEbk9lLpMWodTQi8aL29IvuEzTcgEpQc+T2RGZvmann0/7LL2
5gxKKL8OJB9ydFk1MejKxcx762D67KLacA5iwPkPZJWHo9TYlmkCHlvKssTCC8zm
CAOT8JzmmWq3qL0uHqzQD4670vTKLhqHJv3E7Q743V+6Yc3tGaZEjU39/SqxQ8zQ
jIRFKNhfEw4okTwl9b5zIbb/zD0B4J2zMEURr70+LG9TEKmMnH1Yy6JZlTHDVLRh
QHimItLWB6kf3anwDDEa4ScOqIjR+HnbLuWlXWMi8w8A+XEfh3FIWM3oXa5rxKHO
5TI6vtoyavx2d9vTE2l2R0PLfAtoJxT+Q0prnWQb26km7KPjltA1pW1xC53GI/iI
XTU6bR+MOsS4KpequLRh4X+c7Q7EFP+s7ZMWiQiTGgFQKYEnAelOqA25yqi/5HVi
n+DhM6NhW6ZR7FqaCxTGXBNgLRoUCPq88Y3LgH0xyXqf0tSKWu29fi5htHkHAnGR
SxSWGvcsuzaJ8xXFvnc4glZXc3FqC+YaNmSmDw8jOsAIxCoDF6vmjNxJLHb9HQ0I
HMfhcHsOYe5YnNFfowf5FYNphcQ/SR7Ibo+HNM0m3/WE2EEGQRppwrIqusEPAWeA
GgKdHHTJU9+DJGGwzrPfZYxRoW0H0HiR2TqHgBKTq20MC8v9OBROQ+rcBd6fxpih
Wg2SRC3YGGwrd/Lx19QtzkZpnzmPpU6umoQ7BQcFhJ5k+TUMtUcXuVXFmEHjvJyL
MO/4kmipkQZdAojPV38zY1p2gJ76BYRAFOZbJejdC+FujWgLS6XftGE4NB1Tj1bK
uxZNg3+1y9ToM6KNHtEd6ZvZai8UMPk5y9qL8eMmcs61SJKLFBhtwsd+SSJL7q/M
5CziJtqJnYOk3/ms5c+KjS46bEz/5TYT8MvSZHMYE3vZzbDZ6k21fVt0Zk+afCDK
u/3x04MpNT1Ik4ochc4S9Lr+1dtON32CD6YxyylJDnn+62JNKwyUDO7/skjuRhz2
0kZ9MISpdy38+bVKvFYwLDnlVZf5p6UvtHzxU/UB3bqUzWalkR7P7CJVr31nFbZS
jv3VeiA7YA/0U7ZoyjufwsTA+vBfxsi7xRrwgIHHSEO2RpShyagu/kya6IRgVobl
euyWhNoJgXgxTN9SUL6lcA0wX1kASfL6e42JpVPkjaUXE10v8tbksmw5GxYiO8G2
9uPChiZKsqV7KjAdPmJ8bHZVDQoregtftPNFsaFRH+6NW57BhBYGY/dNlpbds/BT
LR/GylSmE/x3PSXq0ve1m0JmDyF8/ZTWrWQi78uDkN26bD0iE3zzTER6KFKoi8Os
yrwzXr8dVxXyEuARJTMRiG/GNA6o5KeRaCS8fD6N4nmRzcKbcxfB0T7flm7pQ69T
HZhHBDD4j/b9TX7JhFsmJ90Gq5g8nrJWLZRJn2/+6esdWjQVLVSocZ+kMEQm7G8P
DiSjwZv54Gchd9UQKauw8IMjsY4frHp9YNGHbu2/CqQH1kKsvwQyNAD+rG8/9nWr
r5DjBVoW6KscQXUpBKhO+3Q4eKpp2QgXX99EsGwM6pjzeNNJS53S2LIjs6eZBl1y
LPt/SWGdlUfCY815qPBsKHKJEXamnJe5HPhnxkTSOikrUkzESP1YhiSfV0RAwI8Z
7SUW+/X8U+slegvvWMUXEGSC3EUVW9j7Nbpa70UGQruCe3eVru/caLc4bmwTTV2t
17dcMqHQtVd1G5QhVWt6YVyJ3XjHpg6wN62bjpby+Gl8B8I09z0RM3ofsTisC5pf
kagXx35rukTEbzA0aBk3qi3jtayo3DjO/x7GNXbUJtcUSfsARf2qbUz1eYa/zi76
6UtkKLgBW3XxU+K9wb6Lf1KG502vqZU2rAfMYXOPTiSWrq2butprRMPLy2qacveg
7Icl+fnHwm1maJsSAqG76H1e164gFsKvqP5s1ixSeSTCOz55DOuZ5Viyx3uJ0QTO
fszKD16pMbhIx81F5yXycfOCnFhR5Y4/0f4pp0QCgRe75unfjcKJ/8z6FxSB0F3a
N/1wQzWJoFrdWZ8coSU07exDUPDsMFyKUA4ko468FgcHTL+Nuroe/BiGfT0Z3HFh
CyBITJV6eNt9rE6BUyLkx3ziQ50XPLv+Q7jw/np1jcZHGvAl9VIFbo0SRDRI0TBh
yPPVCzfH/XvzH3h+Knw7s2Y4YWqMTiN8zIWiOLn8OCqfCTAx7X1bOvrCW+FEhARk
E40FEij9cVDXnjmv1Q3Jo0Ua+kMkRVF04VsxmwMVCDEnvK2DPNByaYrRwJbE4iKa
K75iftHnLKHM6ws6FlgVqEqnJE6/u3yuABzjWdjCaCeSrJyZ5tdDz2YirWwKFWX4
1ldFHheue29DhjpYunCtg2K5SylN3+OBvclkk5/L//aSMaLM6HBfuCgJafRzgteL
R4kX8QQMfn9tPMfFrc98DhYVtDhjkgtN/xbgGldM7l8aCRIhaJRV2Sg62w532o/R
8tyV5U73ATE7aSBEXlhWkjU0C87HgL9gsjoexrri8ExJuBuOZbK0I0JOWMA7zS7I
q0yC1FiqGzu+nfo+itYlMiOIfnBmzAbW1MD33FlK1dp4rWCUh5nxxmPOOR9/XYXL
QN8vONQHHgdqyb+a/ZRWgYsQumTV+BUXXpXyfNR26GPoAvjwFI813bl8k0BspDFJ
Il/YMQwSCgVXLlTEuVHWFGmIr+EBzEJJkD7qAn/GegJjIX93ojq1UjNeL67G+AC9
botR+bEvk4bYqbI3y+rdI728Gt2TGdZ79OWTiUGDNpBWyCV/oW616Dd83qc45pJm
wZ8LCadiSXXfg3MAYyEpvcqvLdlYRko+thsxou9gURi/80aXyBqH+w4Qq0bG5Cpc
XkDGeiGXIAFWp7LDrpbUyvypUmWc0PINNxHe1+60Eq9kgHmgiPVOxRowM3GLCH4R
W2QwCkT6Ez9NLJwE/9xXvKeHcet+YWBaS2I22lklCFU8M8t3difYd+BkgE8SwyJT
Gs3fyM/yllzI8xrv5fb46gcmUyiZrJIFAiuOP23+nwjAYpqnJoYlb/35r1VK3/kT
Jm/HFLACFoiQrrfNpG/MmTqG3GV7EHyVaFeV+bna02d84J4hG2g6m04bUHOs5GzX
2NWTgEeJK7MbXDk8OofXFkEmoYOeP3emvh79oavzNMRcJFBqtwWBVIgLNe9pOI6b
9SlpXSUM+JctDA3cWeU8x4uWtNyXR5XSPwTI2XWu36jechSyl+ONxGpG7SyjDpgC
fhkHHuGqWybJpu7VJvG36gIB/w8ghgR+Vwo7Ems3IDklOl4jECLNzg2pEJm58XO/
kTo34mVNHqrJEsEhhAHUGI4XEr02jxlRbapG7MC5sl5vBCIbfPYSdD3/DNsNWyOq
aza0fpct+ickYCdXVXvE3mJSdUpwKG/OOm8laZcwuJsP3if54Eu0gEl7Hnp+rmDJ
H1bkZzWloxRQNy8zHpbE85ePWGYKiw3WTBZbLOoSfWnKH8gNjwTjwfgvMXfKcdYV
ufSoJ/uHFOfxyRx3dKdJdQl5vKpUGkL8WFc5A65vXMT1T3G/gajJlxp5D2hHfiO9
FPOEFwgXgeS9bVy9I9LdRrfZGFvbwb94wXkQRIN5QWqVBM5Q5r+iwcNpsDKtzUO0
DSxcK/mGAUBtaQXOElhzZk0C230XRvByz1gWwbRn6/i3PPglUwM9p9+s2aXm/egs
zdzu/70s71tf1OlxztBOS+KAJve5niv5pYu2jcGZCAFKGJ+VwtttW5ctOOA9y/J3
5EVyhFbFo4cwz1EmHtCj2eRq/fZk3gF957oXAJc8zEH3DviYuKcqLBquqisWgjuK
gejOydPrOx0rT9S4lghDQ90V/sTOFfjlDzc+WV4QbfxBnX8fqwoWSfPm7vof508i
mq2qu1T85BfF/1Rzna9LhP+lxW9XGaMJilptkmx7fvrjk8hh9tcmf49jcCAp3uVD
wWTtUoy4z5xEfQLwyWX9CxAHV8XYNNtrS2Qm8hJKtTWJuX89PtPwLkzHyoYT/qQk
fPvW2aGWff1IbvA/nuE60MSq/G4PkUbJj9j4sThqs3TrwXPbQ7tTSm18efk2WETy
sUs52+y3DngonUVX8Qs/1VpCWCADL+SCQm+XCsub8d3OBLIQOoOCRnsSyf4tSMr+
jwopqT6J71/mxSmdaUccloEKIZp1EFI+zAow98GYtxC6B34tAFvR8dgYXnvtIDBu
X7cNFXIzL28aUvA+MnUPjdyxvSiMBRnfi667cnO3JEYKcn8TcSX5KeBLmFlIZDT2
92EWddWGZuEii0opCFF1pzH40huEv0dhPDwNzDJ3eA+tRLqkIFcnnj8dSs82DTdI
ILRoPb44lAOiAXHY5if3CZ2VJUi0LsgIbXcvYPPsw95pDW94iNZFzC8BCDXk/O7s
YMjhcPLduxZvGzpR+zTaEY2FlVHKOsW3wkQWI7SLXqvt/P/ntVecFgHcorHgTJvU
eZyBSa7Zfu8xV2GfTflf34KAPcwsov/axxFG7WBp11ISMMnWJkhAHdXsmnyVLDfi
CiQ3f1Ij++Z/pgC/6DfXE513xgge/KnfsAKFfcn0u0M1QLzvZFJlVC8c0/QNAUfB
IXF1en+1UHN5RYELQuMMi+TCcuMl1bDm1DG/EeCMcAFGp3NGwg6vrmukfLVjQ0bh
J2Fg1Usl8EgHvD05vCv+ScgSnRYgrv4tQGpXkPTh2r3+iOJPK3BLr4MCBVe+rz6s
chIcwirxtJNl71Q799ljy0n/cjAZuVlrxX8zvJKtWDd+nhV/gOZ1FqdJxcw3Sz+L
4kJRVVuyiGNm16HjFQmtghgabw0BTzQDYmCFDnoPURsCWYPmtoUY+msRqr81aBcy
xHpbC4HRUoO5gHRJ/ECTy3vw24KBWtK55df6uSx4pG8b5XaMbpgwogi3xtrbE0V7
kpxDr3lDqWJV6LVVBi8jMw+mpsdQ1oCkQ8qMfX1fsEzBllk+MRdjNqtWRgb1q+m9
SofRxiBo4oapqMUuVMbyGCy+y0eR+F0+/oXQbvKVAXhxwaJ1TofFBQOSl99N8LyV
RMDnJJyfeIm6ggxgI//LFjIuM65Z5qwYjFzovnPUpJgx2sjnG5fCbCHLZN8f0KhD
ogZvwF5P3egDQ2pb80WPaCv/MqAnPNmpyuOwTEiRKZIbGDGKVNtsj44hSDIX9YS2
cHQo2yuaNSPFv65pirnL/4sc8ROv0Yrvrn7I178meoh5U1PLkxwZHHmL7yeKSZVz
nQikfYnzJyZzW53SzJdXDfqhE1NfQQvqlDLd4PciTbDHkMVMlicAWynz707bnf26
+7DTkkWkP8k/IdjfujuWNo/vuX/m2NCEsUaUzC6NrTCRxb1sC6J3jY1JXuP/QMBZ
ZYbIJbS3b3hsSeSj57zt/wniMt4MCkSFjNlSU57BpxWfp+vOuMsQFpksvEnz/f80
pRUoLTkFx6NStahF7D/0EHb+DnRvt0uthGUbKPNJq9QjrcWIpVox1Ww5UGTIZKz1
Asm3NKju6YvIuk5dULeWsNsFYi7twsc2ZhtngYsyRkHqACNsO/DMX+olDuW4XOAZ
P4GvFv2WI3PHCZcynLNomkIp/8XU0q9bgQouXFPWk9BYqbx2VixvVhEIG3kt+woy
sDuTp38UJqOhgK8S5Zwx4sOfn508l8mhO8G6QPrzec6/M5MfqshOCXqX5xruoMhY
gu/GlNAMatbiAYWiZQmcr52PoJtCbvdeLajkGBT8gzh6pxdiWOQvm1z4AB3HPs72
Llpkb7pVULVZ32L3ST4IU+4PuWYqF8uE6BKs3uObGDApDPnq3UfiuaOJ+B7Wgt43
CoOme34lA2RSYznKCb8Nkd2loeXnx52x5ZOzMTWfupznMILeSzI30ZeXL+ZgCt8+
VivaPDI75QXVHOPwZ3q9N3yix37oKPA2MAvQxV13EkDJmp2zBCh3dkhEsV2TAbE1
idMAoxbKF8LutbakpG+TTM9dtrCqcCUf5JDloK7u99K2q+3zq9X4Kxw9TJPHsisl
CBnFo4NsfCe0KxqMu0KtAsJ493XAnAkUCthWqxXeZ3dxSQ01vBq5+sR12AVV7JGf
DF3EOP0oTP7QOXgT61CDSJjUE1+x6DKCRK5sitJ+VHXUFGzXSxnSIeX/0bes23Mn
x7uGLgM6xk4+iMdvVCTRJoOqEJx08roqfZgW/Slq2v9RQpyur/sV8TM+whdkk1HP
gqwv04OawVf8O9PDx+5pz9khJwKFQOgymjzwFCU5mj9/AjSDBtwUoqb7UU4mSIb2
MkM/UkHbmOE8wCkpXPMFWffZC8ZxgxeQMMojOTKmhXcbz1PZ90J7KIlbhisrbtxY
wNHuWSZsg86dWLq/Qj/5v0Q3WYVksjxMA7LQBxEt0GmpcGCTWkf/s7ufKKP90ahO
78ya8ZBeVkL1RD57CxFY9qJDytJdbStUNHhb633ZhdiecuOuUXxeTK0o3DhwbQf9
h3iiti5NzLDKhpRWtbK82/wdvHsYBE/8/op2zZbbVkGT2PMyhb4Xs9ioJKJpEPHH
QGqWaUWRV4O2m2MVSj9csoTK2Np/7e5wXU3e5qEO8N4fcJNZpW9ipnheLMf4RuO9
T0Hr3N0aSqOWADGKS5RLZizd/EZ4dHS8C+MNbZIxLrgYU5DeqRH8fJY1WFUHozMv
o4y/+Ud00g3LX1uNWB3tZqk5sztY7qVv4m6/ooTysmfN1W0/rfftw3h0znnF+Tlg
d6a8QUM26TeldgpCCLfi9jiVXemoOHVuWliCZaxxFlpFYFhTbgaaLUCOF7z6dcP/
TMsTZyIHGXRGZgjYzvg/uvyvaNluy1WrWwhOv6BfbolArFqPadwm2gtHsWrkE9P7
XFbz6qgr0n8XAaFvsTUOesIff9HxFPmuOeXuJcc9QZ3YxCEMwplgW+Aanemm15Tn
BEdGM3koH5M4+OncYYISvArTFsadOpGlihxQxenNQEs1s1KRvf5cunfyHTZVbERB
HJbr3nPeipC8DyxUlFhUDwG9w1n5bktmUa6vbGWkU8Se5zlnGtMe9i5gbfeLWv05
iNrYHQNQ++7WwCRGbT2oiOLd0e2vbTlX4QI5xKd1NtPuOVlHU1JEjsXkH3QmNhGp
of61OoPvd5Hmec0Zsk03mwccBJrmKxjiBPO86JyoFk9jsqsOcue/0trmPwsTH/VM
c+FOvvT0x8IOxJie1zfA6hOqcmx70jBG5INVnMKfSfGpvjrNUHXjyKeavBNwo8gb
F3m0sTH+f5nB0eI8LoUIIhMLTWmjcEjGlbQt1jOZObUeilr3Sqs3rCmcPaLTWaOY
NQQV4Pd3zE9YMZrYEPToJduo99d7Tfab70ZzX7QXpX0rPNHKrOHpLD2KEUhHNL5B
1ISYL0jaaoXVyJDgg8E75RR1BPJP/waWALB3CRsHiPJBCPDFiWEJp16JA3V3pm0O
hVmDiEaOL1DLAwMPV2DnYQ6bv0FoMWWAy38hy2ef9YEZRRiZYvimrsHaTElZpdjz
YhzyuxbCdvxgi8G1w7CtFVJ051YLvcuzpIVRrXJg2NCCpyhdUchHjQTs7pItABzA
oM5TIO7VFYn1q6IN/2Rt7wc2+FDnpQXupd3Bd2/xXVYN3yA/K9xrX2i+eqgCwXVy
FksjszUFxZY82EpDbAFn2EgZXLef5DAx7UpsQL1esiKFuMFADFVv4YAGywFtYfyz
0WJpzOuVqEp/EjqUd2kLxZBEgBf3mM8C+pJcp9EYiYTeJkmY941NiyJSenHOrs+z
HgbiVe9tOwj5gx031/d5Y/Z7G+TDpu7afw3lPUIso3Gtx73pR+jVyt/NkMofcf0J
OWL8pu27jjWWArdAPVuQCr1aoX9FjyGefOx6IMwRnL2w2U+O5u/YKOznY4n7RVTQ
4gtvfLpq9vefWUQF48kAAHqhe0qtC8SPEagH7zVcfy8SNBqy7j1F0PLef2rkzbDU
BbtvXtTlOCSeffLaMH4uLhZWh+5Xspb9O2+HNxYUbqflzripp2nT1RLsNlgUZRrp
UYHc+/zHoubnUvdQ6AFwv8OTLHJqH0dIMcjB/mk8D7trWugJAxLdMT5c5u0dX6Rs
E5OB6gUCfHIX2ob+GarDu33UcQgO3SEtmWhL20XuqB7fUGzs11MjP3/n+f4pBl8E
4SPtgjXpC7/XkqxErDcaD23iQA5JRj+sa0reE8ir1rgFKvP3Fue0AXcv2CD8j7+R
qRimh8cSF15tA/Hg0cdY4blr2KBIW6hhWmWg9cgmlADgiToX7MtvNi3wHeyqAHLT
gTaoHqHcidH8cQMw2ST1Y70IW+eP8k0Es4XnJ8qTPzHdvzYun53ATWKMt2uPM5C+
+x/fd6S7iQa/8CuwSMfeX5h4GaKMR+vRU3N4SiTmQKjNUjgcf7tyit7QM3+USOt2
8tDB4Ou0tzQTFFBipOM2TESyPTWLbUbF3Dhb248uYwz3vDqy6OA/DBIwR5D5E+RO
tIYonaOJt3VAh9RdVijg7Dwfgp8QC60HlNMWq2DtVM1yfkCCgfO1yHOhI463SQIM
LEuDTbXmdEfLVwXjs+8H8lPM5+3CZCUhj1mx9R81y+ZodrqE1Vb3hn7BoduOa1TS
BiUsD7aSPp2/x5IJJwACPNq+bKDqlMklJEkvxFedHfWWyperQ5nhaPKoD9eNxTAn
66+MkpiXTX8eDWbMtTYEk/PKlpRl2V+hBq91+/v4bsdQE9BHAfbNKXof4IexqdHQ
5sHgZiEW/oBaFIn9ofA828Orij82Scr8lb9PSTFv3F2yRQ+b/uxIyySOgVvBqY7w
r2zEazo5oUFIO2WUpAx7z28n8dtKDdaRFdJgWUsAacA+fLk1tkQ7OgKPOnf+H9cF
hTjDpj6qnKni3DH95YKnw4O5IzkX+VRquF7qmW/hubQeuhR5M5IXHe43USVOUR94
SNb59PxZSlk2dagReeUlRsNdEva3raLnPlc/hZf/iuSGFf7otQHAefhqc2m8PmXP
o/JgJ0R28hbgEs5Htu2izESi3831LlWQeCbDNBGT4UdLXBmJZfo05d6J6zFOsYAr
HMt474aNHikpURnwNryz+xJhQ9NyxD5OKzcV7SviCnyoLU+C24P+9w4znPiAFa4c
Awss/HpVgJb12MZajuf9L6P5GKsKltsoDMBc7CYzerEvVsUIfuVrtJ8wqn5WTEkz
b/tFfc205U743JOBsA6GERLG8x/VGFflaj78B1ukurWy5cTCIJREui77l8SkHJ7a
f9OflJev5SBvCEyfiLffmUcfpmfxMY0bePKRRrp5KV4zY5+qxcn3twR7KFQBEilh
EyjSriXrLj2uoSB3sDZ6q+OXkH6nSPnaE0HS+3F/TfQS0NDo8vrapp4MAwc942fw
oCyjY0xx1WZU6c8gBZhwb6tGMVfb/3qSeCWEuFEB590HWNvo6mHfqiuyTMkx3xgA
IJgJ7MTtxxsutSFG2Gu1zgdapG6vxDzCyOd14c2/lTicaKrcgChNY1craXhhwpNX
8aL7/5KC7YgARDVnBk/K8Pqvc1hNFA3YJtqaPlbEYj/q0oSXj+0at1qSayvMjmLr
RjafV7w4zmrH8bEEIP8TiHNTjEYlfm4mumsNHEabRUumW7JwYA7ohuMhkSgqNbFe
aF9AvrrxDb4CkXkoxcWyCVE+9agZz2WFZcgVWFfdCaNLcaZBJ80dd0U1Ho2UbWW1
RD7/8CDMTb8YKLZ8Cpn57x93sWRSRudXWQsyzis1bkc1ipKSB19Q/xoFTd9i+cwc
/nOeOj4DzSa5LQLFUdktUPNxU94Yc23kKoTgdquXfH7h51HvFnnzO5/KR7u42sGZ
d+DETkoQLqOlOYty99Uo7hpjnAZh8xTqs1WVB3zIPeI1B6etpoh8RbuBJ2inuH+x
QnTLZq056KmsQXVGwgZ/pE/JgjoutSnaAj4YhyFQ23J1X3T1TlvT7h1z9t4d0OjF
v1xPO5Qiw56NpCg/KczvxT/QPeMrn+qmohBGhN5HK9DZBLA9DIriHsGkcW1tZAZ6
DsDgv5WiZ0O4Pko6Opipq0YqoYzi36EgFagXN0oAR5h5K/fJK4gFesOdtrNTMoFe
RHvYjZMYbSsT+ZTCnAMLTDU54O02Kn1fX2TfALmdbJHCLDJRndZnuuxUD1nh/9O7
9k1321BzF4jhcgTovqh9LwdZ1IudHv33rlFzvkElO6RpVvVkyFGsQVTsgM6986Ej
Cvv111Yf43bbvwWU4z7gXZeWDvG0nvoHBHQNK0XZxjLQFaXvRi9vXUk5GPAYUzYB
MVXb2S1X4WOnHKnynLUGG71xO5byR4AblyzvnExLmdymiVx8J+pCU67u92itSTpm
lzso5qnWY/UUhA1g5kVmbgbfLQiT3KBrOxh1+lG6umzCly+FIlpJlsHsh4+owSgk
6lPNjEOgiRmQY1DVEnpgb2qpIBSuzGPOt8Pf02nO/vkOg5PsPY6A8FyzOvJ987Rl
PePpRq9vbhS8bvt0OHdAef3aH9HdqtsaGptr5F4zvGraX0j12qOiGXRjg01SNqoX
U6z0nzbZckOmB1NrAf6G3RzVXFDxtedjaq8ZTn8TVCXv4XjF6qwNTIDcE5eptfzp
KoOg6jkvWsdQWw0apkmEv+Z4dcSNgqazM7OLqo3JEzarHpgkdiLrDyzE6OF6jQ2w
Rs8IuRMEP6ICJdyvJCNTWcg5m+6bSH7ryo4NIQFS7OKiSy5+Vkzx37QYTvYLlLvf
nPpOb1DDmibG1dUA1tshHfTVNIjiP0ACd4euJmpmBLOxGL/Qxo1o57yElAYGS1Np
2M+ORBT5otPV4cixpQ0OZv2B8PjYH/U5UaBbPo9EHbX+O6Kr/a079ifZKsKxAEXA
Oagu91bqm3Wdmgd4Po9accUZ3fYeUYYn7kjNz/T+hY0sqJ/gt4s6KRYYk43D3rjo
KXp/DxNXGbfxcDXbreFrW9MuuNTFzVDs2irNnx3lFukUqRJg5JN4n7daX8ixqVNS
kYFXrjhj9ElVP4KhCJyXOvzadoA732ff6bdNnOXLnGvzL68ViJ7SorunOdM15lE8
qFECx+6dNByplzA0+x8X1jmh53SphoyqpSh3Y35liYh53V1J4GA/QP4muGLvM4EZ
qnLfgP0V9Zh5bSp+KqbfqzWO+A2SDJaj5MeA7XDPxaZ1UlMd/ZC5h1kWybwr0l8O
ZyAnGouSz7qj41HMiEO0fQprKDnZ8uCLbj10VHdmxXhO1L2qNiD9cdlkQ8uH2dP+
FU6FeqK0nUP/jmC4rhGgNEeDnLIkIOixu8TjlgwB5x6ENbJMJZYjIhZzyUZRYvPt
faFtgimFfFXuf30iwtGMQ16T60UVi9Pvgnex3Q+mSleK8kaOYT8n1YYycjipkAmw
r1/2Q/4mURa8TdYrxc8ouSBn7JO6G6vW+mW5i1y1GjDNHX6QNEwEtzSnynfl+MyP
CfOQ9cwMbol4iW3QKMYHzE4UX60Yk1c1OECYb8qdz1T6clhfP65K4DaukoWfgCqh
TX98l9qMQDSZNIYyRiuK01z1QWuXu9lHPR32XZj4cTKdYcTy3k88sTlC1k0DAaXC
r3IGeRrzC7eKI9YWNWxTy6LDLBjNLBlEu7mcRDc1dHgg+DvqKiY/ZWxjZTy4kblj
DYcDeGnPMUWZ3bKUWrzpWdeLBNh153r/4FztPovvIBjLk9G2xOCjMbqrS3o6uM5b
NnKA/cbAYqYbpeBmzJV7tJjzGwlDMU/ACn31KA/zpiTBI/s9Ame9ZHraXgOswXcQ
HUJQCp4zwNsp+qyugIdacFcomPC62iPwZIXGJkvqhJpKBnciUF7ztZwtbGU3m5uO
AkZ6Sj0RA0QxA8CMr4yYC6YwVnqPLy6vRVQyRSGR6NJ2vH4PG8YJKyh4J2KMhVrM
LcO9n7jRzjAY02OGA0W2HzhLDIFxkHmupflwvaarAY3NYBOw2nRnsWAgEPd1Iwpv
OWz/r7MBmVdmSVtDZisZkLSxe//r1w72uUPpicbNt3Q3aZialOBfHJFkSmuhu5vS
ftcQt8zg/fWJPgv2Xgo3Thzh7BNQVh5ia9xCBZXUYGZVG/AS2+OOd4o4DGnGlU7l
3RTGXcFcwLgOf2DDpz/5qfsj9HUCFA0Zz7KVv4dSibu0CpfVc3y8E1aLZ8NYhP3X
o264/+Jsos8RObBhAn3ruV+zefLMlr9GWCiKU4C+bKjPaGcHNJLYGl83AbMikAMm
IhBCuGS+ZrASuPoaTPz0TWFUuSqthOKUonRRObHl9zuo4Q4Oq2bDHyvT3OhC1lZJ
QxRPJpHiY/0JeBG4ldytrMXNxrRKdqLABv7SN0rD5kAEuGXzHCDt59s2rEi3vF5x
3FFp0Zlbucg8sfhQC+WX7m9CAhogZFEYX9/0JofeaweBS7a2+oc0MEcU1V3uY5UL
xXE6XC1LG31BtuoQZJKNuQDEQWDEW/F45lcdLzHQg2Dnnye3Xlc50t/3V3E7KfzM
X5P3shZH9M16qqo2LGIb2piNS4DKUiP+LPgtJXJ8zFRNh8wFaA4XTJRH6q43xz5F
WuGzgwYIWbmg+1vnbzif690yoqt+ajnHdNNLaPjs5bqVzr64oe3YueIZWYizfOKG
4FMminsOtTAmgwCWseVrDrfnojUu2ZliUWUoLQj6cPw3kUfnpZJoVhlBu7vuUrii
9iD/7WToUfbpUs1FMnhm3YSC/mGzhIPCuRFGwC+59GdcRfkjqMmrK3zq6+IdT+VG
QNSBrurMeqPioTt9UOaVDW7kaDy7sFZFoxn+gfOSrUXew1lLAHkOb7xrjB/ufh7c
qlPsyx04Eah3nkxVSUZdhRatPk38zb23z07+E8idzCqLZop6PFcO2uNVTdaiI+SS
ZF82CG+QJrfXRLmQ1BTPOMjbX5xqDpA6YyH9dD9gsWMvUWheWjZ8V4p1FAh5L3ip
5QrnXxQB6OQElXn4GFO+y+ato3pmPba4VyPPIeSr3gnsOQxW8mij1boHksCIqXMz
WkE9rrUQMm8KcINrnN4pRdlLbdlAgnMe+cpwa96ebWwQ+AQY4s98j14sg9UJtc0s
OUcZN+6embqOo+z1lWIExZDyPAC26gX/vNE34nfFE7zMbkcYNr4gqbfjiSlyThQm
Cz9j3bPSIgW60ZkZLePuqXTrppBAT8yr7MiAT23ZGtXLCjgokyid6u+G3pNeEdBP
U0w54K29Vtxi8gIkD8TFqiJNPLrBGIHgq37IN2X+xQ4Q76nc7dW/Km8wBf43fhvB
7xx2m/sbNsu/7Da8WvWbfvGR05lRnBwBvhmm1LTzbW34l7aLOu/DyLAkzV2ArhbT
NKWOPgiXFZpmNWIUQgZlMjn27nIANNec9gqLyqOJ5GTAXjQqAzmE8x7KMns0z6v8
CHGBap+r837cuXoXvnRRCebnVQ51FgRvJOYxutOa83vK+cMuYLqQmL1ITaaSzFRy
VZz4iYhfz8a6dbvCJa88bMtFAY3oSaDI8qd8UxyF/alMJGH6Ay8OaT/fV2Ff3zcF
9dEGbXzJ+V1eWa69PUfM4Usixn1AQ/DLVeaNpyVIt/2AXjLT4sXDpkJeOxRcS/Pe
iAdHeczYL7zo5NzQ33aAqCUYFRuH2rHH21bKfxxqcxCELbju4PVDVospFQjMUbYG
sXs4F7/WE2K365loaOKJ9Jdl0wjsz7OqtaHijGlrtl28Zrt+bmH1UnvPOcojOZpS
z+ud7mN5wsNnVJ3FxMFIgEmxCk+THiIBCUNYG39mrCBCVUk5wQt4uVmetNtKWcxW
CsvZ1s25ekqTCqNnBU963G6WQ4hHdVxi+68HNC7xQ47I5FGxW8J7Wt6YkzgH2Npf
e/YVml6rrwK1KvOJWOUPdF+r3iDPY6gZPKjZ6lMOKeUBHaGqL+4N7zjIZHsr+BMP
VY53g2VFL90N7/LIjssClcOJONp2ve5fsybtphfodrtKjLMDQMXHBid6usWdLlX9
kfv95BetJCsAH0cULNtB/2E5ib3jOZk11O19VKSYAU4mS3nj5iLnX4IZnETZz6aU
g4PT0UL2gUrzsqxtQvGHkscecGibe63Bqv+FVHJ4rErJJaR1EA0UpUHbg+YHjk4n
tg6Aozc5hxfRIRDQJIh+1qNLKm1a8mtK93UURdPkgQEXeekx0LxBaH8YL3shEnma
OUl1afQlO6HwWYwXhurdPpR5VjEa3c6r6DqKfWIFulGcWjZcaWxVCc3yzMhIbipC
AWpFRmCT/OqaSAJdUmHELB/Zw2mKOHCIec+D2yDT6MFvej7vm11g56sJmm/I9quR
AKYLFj4pmIJgp3cv2zqJpBUZvfDh/sxtlHq8OafELSzelWgq29j3Cqn+UY/Jdyep
FMJzVZDTKrNgLmhe7Quex/p1X4o0KQlTccjpAkvpB/2Hl+oAmqo4MKF1Xm0IRjhK
+8AnZV9sASXyMDWhmJEZ8qLu4ThWK64KBOH24y25fP8NTJZg88z+1BCbBjjQfI2+
awbErc4p/rcXDudhGn5dKvvatSzV+yg7Ij0VfqES8MzxUamrAR2do12r9k+QmmKv
O5Pt1j6ku5sv8FzhhYzc9qn+k8jCy7jYyT7WX1T0Czi92v1epyHiGzmbCMVDqrBE
WZgS4Vp0lRG+ed+CbYbmMavo0EmYOwIDFh3ai7B/SsG8OklTGKJpqkh6+tsCaT81
MeRepnmiK0Rk6fYKMp1j8QG342UCS3uq35ABu+hlWjDUI5ohmoYnSb59XdvM8/zG
NIGTNTdkR6p4vPIaVQUVhL6Ycy2LXTkjse+Hv+3GK15B+jovFI0hR0NxxO8cvk/o
c8z0vj058mtQHgRz5rsdCECRqkgGXMKI7UtGkIyZpOf/jci+ysSD32IANwEf5EyY
ke6U7acaE/vmUP/SiianmRPStaKTI/orOY1XOjIA5zKKA3ea+33dg7JCSiKV8g1D
2vvDf6OYMCrqWA2dkuEBKvnPOMt+xB+FjV3ZgPpbvOAMJFd5mCtAES+YrJPCCeLx
cTBeGsd+YHhxCIafZxdHDJV0d6Qdp9FudhyNaqeVzG7Qj8TBpL4odgAU8qsa3zGC
5fgYva2jic48WxjOenUEimRqlvlwBeNQQaFvNCqU4WVpTydilvKFvNBic+QRS5Fr
58ZJ62HEFLx7YDoM1Wb3+IlslTc0NS+GiYHjvO0houXeT84qXIQgELBssBWm5ufT
2bAIpeDvDrvcyU4IOc23yOAgng/UGXmZTs8Mim4HEs9hDw5/7BEB8UcZj3615zQY
kX9TVyAv/VD4Y3iimIcbFjN/xPtgnzb5FPTSjGTro/Y68afHulnWFQEZkBtNDvqV
5IBwRz5SOohZly+X6bvYCDOavI/kMxRLg4EzOEnLmUKzFoOD/qhhpVK7LBG8Z2ED
b1ddbNooNG0UN/Q8sEY8S0wOSYlRh2nKDaBFvMCJZ5MhaftOWj5pBx1FuEnuqDU1
Qtq6gc8hheoRnwMz9eWP1zJQLOXRaAX9W3qn80++D2HnXINDOW88ahghtQ+clNJX
kRVa08moGDT7qhXMEwIRUjd14H0BAeEtexS6MQbGZha6rdaqV3M6HXoUFPDLhbGc
vVy8ONR0jdLx2trXgg2gnqK0WoI71MCAJo94h0aAU2gwsg+0fOryj1byfF5ms3UT
xq8h9e11Fkz9qBDcfWPHc0AHEo86f0IX/mYnZoHJ2fPeIB/erw7pIMLTjHpl0GTH
2wYQHbBnxjC0Ryzoc4ej6R/QRJAIZkDiesoYpx80IbfgrRJOAHl3IdOrLih5kJB4
JIUBp6NvNaEKecv40jo2x4QsaxcpM7EpNzt1InGqCwj5gonJWCXKRK3hvNLtuEXw
6H2bjeSK2vfk903kO9W9zvLS7TIXSJLDmbr+8dQnnu1P8cZF02IZrGpHHkzOk4+z
ZJFIf55/O2VIRRdFZgsiS60T8dNFfmsoo0Pyk+dsgxNhkl4bwfWb3SUoBT0cnul8
iZba+TfO3zdkz9yf9sm9i1aiy908o/Z8E05JiqDXebjL9dxVdS9W/2RSFJbsHRUU
A5/NcvIsiC6ZlKmSEjDqKWjA7acj7tt2+Yi25HTwoWzA/WjsC5VPQswJOvniW2vG
R0Ew2IgPzLXeZRQlY7byJum9Q6vwoozdSFYDl6IsYXUvEZmFiHlx5ZRLs3cVvLTt
BCfd1t1ghqAITNvICT4VDmjYYHeCqvDTxWQ4osVf6sy7wmeBeB5EU8qsKyiYK8FA
axDTjB13OYdB5vsMup517TOyhUjWmAUzwQL+xmVIX2S6pE1oygZE0afSLc71F//x
b6tohJyUBMBV4M1rTgPC/hFSmpm2/22jpCc1e82XEVOixRO8Vke9DVDQGz5vAMGj
ESY0gqWF4i8J2DVI9zKtEThoJUz2PZWYFt4AUmnm3epXyj8fl0Ijm+qVPzBL5sFe
dGrlhQ+Ix/pFz8oVyL1Cl7JH5IqTf4u+bGIpQQMfbMr9jI4us8WM1xNdkQfKAHP0
jvvPQgM9pSGLWKrmomGR4pphHPOQPghYym2BNB15+rB2ReNTmWwsh9XUgGwciF49
/TydUYxac1GeUas7ArzAN+Ns8XmpNSoIRiosRJEQh+BG6/fxBFlIxHeITCHPFLHZ
2eNORJklbLdO65vgUycOXKPZvFzLyOQsjIGGneR7K+gB8cDKf5hJxUK/QPN7sgLS
3oxwfAfJpkpOp/1pTLZlDQdSq/gxYtXkNT7yVS0uT3yPo+Iy8nCKefw85hdSZmqY
INo2dT5yLpBSvWDfHZ9/2U3W3LEWG00BWSkED5s54Rkz0fCiW+A2Sn9GZPHruNA7
RAUoBU6bIve5mIanv4pG7o88uIX1Ct3F+Maw7FKcQVkCEuAXBvmy6pB6EGJxvoF1
2VpXgqU1pFgxziFghN8DPLUSsw6oCZBB5Pk4tvpjJPqQJ/a4/QTo6LwjRL9z6yIl
ZIW8/0rxXCCsZzAPXIqkavOWYS/xE32KSKL3H7ed7PNUndDgiMq3zRpDe5RKhw9i
pLwrh+y2K7clowa8gmL8T0by7eV5hbAxuJgBXf4bZNJXuB0hi2j1KJq5IT8WLzBI
f624QUnWyzgTEGKjszM4NClb/2y7uHUBcg0dMjYF1c5AB8FZBk1yOBa+gey3yzoL
5QOYB9z8CZwqp9hNgATmtJY6IVT36o4aWDuNbdtFxWaofoJavzpsQzajBack8tD9
D2Mx1wjww62ajQAI1F50LQIyMqfyHKPY7zrPvQyyOj9bGTKmA8eD0ENTUcjqeCJP
h3+9GpXqmEZ3W5JWY1VILjaoP2eGOUQhXBzhMeIJWy5qq7VkNCgM0NhVSQVfbaS+
qssTF7rEhBJEJQblwsBXZNy+0g+x+lIY15bxGo5X3ETJqQ064JXurYUqA+9aOgrd
AD9Gi6356XQzreFSjknFm9FIKpZIc7+0RTzm99kLVM5rdTO1UaTwpXTZZUtqDKSE
sWdnIFb68b66jtZHax8mCXXlZV/uA/mjWFbHOXczjGoD9XszrVu/R85vl+dGSNyR
xlkx1pRVLQiyHFxsXS5Pg9mpBHDpmM3XKFV8A2cnTg/aB/vAxJdH9X8/rcaQPDT9
pR75P4os+bSsclhKaD2Q97IgSPHuvcP697VY2mNsx+Eykst/1uPirG13tTfosTal
m/24XPfvWkRUYRHNterB0XbH212MISTOkswg9v32aFT0FVu5TJM3c2z5qcsGAFCW
zn4uuc1/PRshT1hFzvgAzcWc5fmarsDkWBNuKHs4JZdCDzy6KeIbG/kvAssdrtJk
W+q9zPS0xphHWEeRlcwAARPDBLNMeQZVMtHY+xa0+LwiwAtWk/8Kqw8+6shIp1RE
fU5S2+5HFuuNBVU7Xsejnx5vDc3nRtrVZx6QPDJ5aeJGUL0Hz5nhrIj/ohDREHWd
k6lsi9r407DOOSLsgNppnCZTVX8rse10xQfW/5I3hKAhJsqQOKs3zT6ShGRvNRL+
8o87S1XHk8EgeMDw6BeHlvyblMmNjfs66terVZVvO3fSNsK6uNv6aJP2SZjTRlgK
Ub2P2mB5szglhwtJYH7k/iKdlhYzuwDyQPyvWIdWtuduJj+QnmrSUhGJqCSAw2gx
6LmWecRA3MF9MOXsgf38skv0Ga1RKklzPSocS5jBmba470GAKB0aG1idJo8kFs3F
bt2Vcoee3Za4TzIAJ1D+6Z+VnwtIo3lVsibSUP1vOdY9eXb10FW1urjodrYjhaco
xjiYKx71FEG01F2sZqCB+3I9qjmHnLkSlzJhCaCLDbR55MTDHCGtX82SbAiKKMu+
DJZkplel1JKToKcpfBv9Y8/IVqoFJ89awGxcYZ5tesnGnDv8t6nigxG2xa4eUeF0
Ly9le53gEh4+InglrExWaU+aOXw6yG6mTJ3xpIxHSrQ9IG1VxsQzMrhogS0M9scY
zCSBGWRTZ5crZQf0NlPM3FqEHdeJBl/Bgyru5e0ZjqunVLfDvS0KS0yfEWMzsbTr
CEJiK0b75KKrdoY/Z91mKfw61plPDqVusyE2GtN58DzHwMTC9ckxpeYr9j3mzf/t
lwaEOvkQM/TrZ/3vk+5sUqP9qpKAoj3aLfophEBnqL2tYuJ/XePZDJYc7xe7g2ye
80Z65RDg3tZsR6QQlcSntAoPFE/eyBUa98+/Wq+ohej4FkMEcOhq+wCCWGE8UuL1
/acevUknjiQXJeBmCpq4kvvSQj/ncjV6XCDViiuyHE9P7m1qcIjTOZRE/rjPsZs4
+hbPb6JPyTF6S9dcvRr48s6cngr4pKFD+wIg3rh1MQnbAx09yDDaUeqdT8HjC4ic
9x2LICWDasLyMTOLNkJgQN+2Qs0swfqEL6AA5fiYU4+ZbMnKMrNwi44NJ0gnngNK
gHO8wXceB4jwPySIYeXkvRbjs8QSEBGpnczHSUmckrtCrdC3+F9JkqIT3P/cDUHZ
eDcpXfNmNZhtAQswPFjihl9ZW6v98sc3eA02UDbXnHPwu3lhTK+GT96j3A+hd+/I
hnRew+W2dm4E/lrjPO1T/CkmXY25eRRZulM7n4sWJmdtmEPXH/Th/YdGoC7sbaP9
ggPwaZF7/lAkIVb73bHmUi7xBHmlgVP/yETJIACxGQ2rOAKe+QY1Uq6YS8D/FwEt
Uk/R/2WygzNgzA73D4azE/8a+Yx7EscHYG0sLdM2F3htQW82OQtyUm5pSf7lDTfV
V6g5q6rpnqmo7IhCB/skQLyBePsvyFxOgU1E08bAUZqx8WUDIvyQjhI/OxRPJejx
/v30yr8SXYg7xlqLwkrhmjFNDm0aWm5LmZiNyHD7AYEcpMEekPv3QIKj0YnV6q83
0LItsWX4c8i20t5LOmaDsxuvGylOqbVGz+p7BGu2WJQL6FP53bzV09OxUUdkxKoF
7z62ZD/UTs/dSekeX5gdguRMGru89DhWpR2hGO4QFwFNF4WNUObcjNhIasOPcdXl
37YBrzVyyVAw8DfNwNpQB73uf8Tl5tsKcEeNypBZKmDhA/ouCDnqbBpwZd7C3xGR
XgVwwh3wMWY/Mw87ufIDGIutxWc+Wz3sJboFSDbeDd28y+lZdD+/KEUOKM68oe4A
Or/BTtG6aTnYbq9pq77BLpsRxpJGz+oitB2iq//FbS2rqJUtJXSGWcppjlOcNVJb
EwR9iwkTT/vpGxZSWfay6i8v5MmcGPh5E+hl9gXU1BiNZxZ1aDxZOGj4cUBu6HuE
P2lRXpmbu4yR7cCeZBWlHoOpcRPU4N2/ad3WmMrOneZMZaFR5TXk49c1qJI5zXIl
6pAvwD3UEBHLJyGxTwD3MeOw7y7PcrzZFSZLdAmTDC0+6zA47h5KxX0OP4JN5YSY
uOLlgikhvTGxur4EsxE/GZGjWe4u7AqcouUEL+4dh67kBKEoBLQUhVH+9YraIIw3
RQNDcMDDcHDkAueSt2mHB2S02zkoAMzXX/heqcTQaALLDtjlMvzxGklQapuvP5+n
FxO9whagCJTAQHvmBsaESUvLlIiN/48OalFGHOU7unuA/4DeOnL1ONaJtjMK84Vp
NWtVO7SklheclLEtkHmIKyCcWb1oGGB+bNuINpuJzCWy6c5hF//2iDmGhaxEo+Oh
rewNjDFLPG/YervlVlQf3dKo8VYjMteB0YSA2SSYKy6hbkGwGnPDtflJPF2HUJd9
/hSv3Fld1H3lEVIGt/PC9ciKk2ynUQAKY9qkP6JsqGtAZDWmdF+7yn4PuasbnyXG
wR67mygBmJm/e+SQL/LF36MyO12bU9OpVMwq6nbz37EoI6z0RdWaPZV7v2MhjDjv
HQlzVeRrh4MNFUw6OH27x68aCk2fDY39zk6uQSR7LJNc6xKdLq1FfhHq4YslQ0KF
R1hKB98URCvForD5Wi2wOp1QZMrRUKUSl22YBnUJgpOhdZJbSkken/K5UbXS3Sew
0asNJ44yQXp48N0Msz8oLpnFFj2AGmXfC3qdfiORFl/CfMnCpTfqyZcapCptSlkN
19JxhReN3yw62rprT9BMNc5fjqPFBZIX2eVDRCSNcYX87dqj3gQTRAvbotqVQPNQ
Mo6fIINQmXDORPCMlNOPGC8GTet5VPH1tGE8k15RHpekSoIOYVReLmzMpJmi24kl
4oFBO4ULp2hWCIBtuaaNNs8gl7wtqL2Z8jE6TToMtrkXDvciybFVHDSqbXjYt0RW
lDWtAszxIvNbt9IwEUDInUCFFYHxmKjlykx5pE2f3t18RLeXxY8a06eNi84QiO+q
OoJ2RZTFmRLd9eSUudQHcgMyYSMeOUt5zZOGLLPVIahFYe7uByF7XChnYgBAB+yy
V4tTuLlBzvIIVD6qys2F2cv9iO6UnjgMEBx9v16t1kxI9Xv7UCafo11wGPm3UtnP
mFz200fW7JACTh7sLiNSjMLK8mAViNqYoern1f4nAeZ+PrVqizwIAw4ggNu1UDpa
/O/bUYYcqyyC8bkwn8F26EGZtYhNNd9Dv5XIM69Ho47sIpQ6pDM/8GkExj45LF+B
miPQs+kmmUYqzJua4ICFWr4ugyADcW3u1cMBT6+RY1JsUQPqnfrZYRWnYNdsIZf0
ls5CrWeQ5WA6bUxOzSpYBjotcMlp2rZe/EiFn7ondRNn4cZ2/ikRiH1LrwMxK+kL
4O/2pJz8+LA+3UpcigDairzfddTPAGZJxbaP8QDocDFjRGow8UVwoeLJTmdkMIjE
r9nSgcX6Jm319IAVMzKExLIbzare/GiBvEOWZNfITzc+DbxZ5cpYRwgnfZftiHS/
npqYUMNmcDB0BSuAobgPU31XuOyamvzG6WL10Ll8hNdNlWiYPHQWjAGXiPop8x4j
czPYgzxw+EJAG14IoX4NZ7fD5VWh8H3/cdVHh1LLnDHY+n1xuWsOjeb99NJ8Dp+o
YCUxznXhFamOdliRueOubriQibdW6QwxTCCHz4Ogm9Za1wCy29Y0Ef0d46yFS9ZK
RZCYP2GPf+JXLDyjgkOxrziTQFNt5Ob6XmPMjM6XI+ioqNQ0fjLEEL40tRqkdMcX
7Wg+rD3qHTh9zCnoA53dXj/ceAHc4PdopT8bDAyhqNKt8kZ3OGEZuvtddhMBwOQF
FQWPjn48wDjt3GAbG3lFLXCwtY52g95zD9viljoyXre8wRSRLC7I/5PdohcZT4oG
TSuhTYc/ki5JWz2pM8OquE2fk7J1LVQBqQa7QZME6Ur37i6nue19H8iUyqPAj1dd
N0+GDEDpEFW/4PODZo4HttFxxdpaoVjwvfxvCtfMUgILXJ55ZsGtTPoN0udqHWjP
og+gnLy+ksA3tkwOT6D0qe74gIbBHVEYYh52XsjWAmzpmlTumJqgBXhtUjvSxokS
OWYhRlU+jY4NirLCQVOnuWX9U5VcdjSXS3S+BwPctrmiJL/RGnai+nz0ye9Xivs9
IyTzdZ2qFv45WNXujRJmrk6d8kcPbW2+hw0U4gon2NKw1Y2HVlAr/kmzlW6TQTqb
1TA8CUDIphE0Gtovp2KKCIsQ4Ji6BRf2UxFp8BuXLaYJZgk3lHWvZFrDBc/9iFgH
tnCCIcDKWVXNSuuVtwgzKUmm1Ej30gaEBRdzaB2ywZ/hzdTZLT1VgLSfqz8NdoU2
cgDhwlXOjrsfw7y1xApp3s3tR0hn1gjUC6uRSoep+Yhv5rtSp2cnsj6YZgJcaGMq
qmo5GifFxNxLMLyyzkjol3L2rr7y888n2siyJ5tDP4VB/D2TwpC9XwMbf9HU8GuC
itacTB7TLkqFvMfSpmMtUhZwQ972hmRRmck8vw0nhdntfoPL7u3Mo3IlFaJuilOP
E1Rk2JWkChu1HSTMiebQkYlq+Dl2KfKpAm8qd9TdxPVWBn0nlSy4dgU3YOn+AGMw
Pe4WPgq8+aw9GqEed9lL3g/JSRqis9FTeB8L4+57q4SxwaAoM2jKozLDs5N+HSau
0olKfXsL+5Ev/HrXmXR/bB6nBcR/ZaIppuW+AxO0SPxoG2Qr0Bv1KZ4wUoeUkY3M
BnkzRm4lNOKLFoJysqXv04FoVWYZR0quDCRsVceyrWWzTWWhcrYFf3CiOfgh9jVt
IVmy9BCoIIt1gCMQtIP39oL/wy6NGsvnBrvM088NUJSShQ2kTd1ZPWpnntILaPG+
AT+lY+rZZNZ3dQ3DMREfpr2xpZ8Q6iKXrUx5YYXaikIV7r9fPt5tCmDPMIm0aAgg
FIkX3uyB7/7DIZAOnQTIRo5dCQLmK2K51rIaGrxZI4C0ZaSOVq8ytRwfZPaOh4TO
CrDHsA6vWZr10LtISau1Ue2q7+d8IgyEl3aub9gWduQ92sRwquZcpD8vYkIMHNf+
HYz5+6LUP4g56DKUYZfjPWBxMUaROtNytds9A8WequfF2PItmmMFaBc6M4UrZhfi
brFPb0PRJgsPMT3JdF1FAxNMlClXT7KAuYKKfxoRIj0DmQZeUlN8hj0cclCdZh0C
9nTmtK4RD4lcw33Mdq/CkxP3ZPK2Yt5wT/EXzJic+2HBIt7FjObzdLC/abGH9ug4
FHA1/Hx1dIeZhckODtd6LFwtzJexzmxHod7vNDBIYudmYCa34/ajLEb1bx0/kdHi
g/kkev8yBgX+HRSfO8Idy2C+6LjTSP6e8iP6rYSZ11bZDies17pBFf1/TdXlLC6c
78m1X8bw2axo8Y16dKttyYh4N5wDbEZPPQy5drC8ywvOYn1Wve8Jki+sh7LYmeSM
DzwiAG/jRLGdg1UkmdnIjj8hffd5YYd7JUPyNsjsKysRdm7lW1Qowyubq1DVaKtF
AhtJH3W9mNa17483WI9aZjwrqUSKG09z7byDNqVqUM4asfbTGTKy/286PL7/op0x
x0SZ2Kn2ukEM7ULMIQvHtc2gOOb3ZMxjBBDPhap+bgZM3ZuhqKetuXLqKLHObbHJ
5dlKvSvTjg1uLqOvLUvvYkYKkox7OtCEvn/6wuN0AFlIL1ZfLGzXAsuoapGrJeOF
dZWRvLWNBTkaZT7DchsmPQJTKywnIeA1E4yINRxNw7jLlPb8mouwIJuSDLKHFPM4
evKC4p2SIXSayJ1paZ4pT5YPoqZ0IGw2ISari8pqxI1GjV891STs7gStRQuo1tmb
LU9RrqbnMjdEDsEjc6vvu69x3z+5bKqszMZn6t5xrapx7T0Ozc3zXUfT6iiv1wYP
KJfsiz3poRXMH9PuHObXzv5T8wLU7h0AnNWGccifWNKBAhoWMOPBlpI2IvrRClpB
7aRGNCt8W7doJTUqxEL2QNsaa+lOOzR6abr7w44BFVz2C53om4j7Tm7DH09Yko3s
kZnzC1Fpp4iw+v7+iQ1Vprl+MviQUChnSxXFj3icq/jKRO7OWvwRPpxxU9cdOi1w
LzEoVR1Hz8JgCLh2foTcflPt4m+kmvYI43pmOT2DZi5B1fOWid8qlBqOUwhCe4Jm
ORJJyQ8gZChgs/qJ6egfzPRnCcSihYbMXBpou8+8bzrvCfhjWRUCbtL1hqdSLull
umLE4WsGnLg4HMjwhSEKOVOflNBhXmUO81gWh/WmGwo/Vaf6VTHKxgDc69s9LvY3
Q0sTnTL4tdlR+o8MtbmNFK9M8DD3AGAGCTvnzTlCeiPIgGg0v1siiiXQHL+NIoBA
labI+8G09MLze3s6cGFhvUBCBrMGRNTuP9/Ih1a0iu63pjOdatYnYw/+6cpoyRvV
0GDcMzAdkXYcaauhwrdPXf2XhNFfP6SBw5DmsNY5LTy3bLN12Kkg6DkDLZ4/Iau/
5ZSSDudwtd4zqY91Os/gcmbR/LZ+NNnsU27OJ2K53FGNn1SGuPAHAJFfx1hQzPKQ
DSYTsbdWwiyJ0mNbaJb3xsiShIOmFL1Tw5iEGeFqB1hk1P4hD7qlfwYePuVXzy8c
eDifA9oqlSNywHyKLiWwolr0J3/j73EMOVDecwcWWjJl5vKJ8AN670JcMkXEy4Mb
uKZbycNsKanOEMjFK4c1RyfTEnNL6eFQHiR975fv9xraI2Wps6F+6y+E/Rolr+r4
S0hgQODkrxFQL3O01dlfva3t4O9eKnLjjtseS8IPnwBYDglyXL6nnmSzP0uyzCt2
9VXde3TlGWMrlI52+DmSMykHBz8eFldNrhFdq/2WMfFCt/tZTSli3/bauTePjtPa
gM+MD+n5cEUJa4T6VLpypXGAw3W4HxuBr5nbG1w/xKRKeRDBACzHjtVBHELBLdaM
t/akewUojAy5+oxei5gcmeRsjAj4Xg/P0yXB+QS+cTgQjDZwRzwlp6g870l4IMA8
AE/7/2d8ukg48nBKGWS1Xlb/HO5X47CjlOm1xejaJ27pc5nT8lX/kVVAc31Wda06
X1MTovvGntHn1uzFfhVVsRfRU39kV7uD4FZ/HQOtbvIyRIHZ3n9q2RI54z4haCyL
uS/DoH9qtL0Ijw9QYhS1gJKV3stuRjXOiEdLXJpAdzyK3vbG9dseQWzhNX91YMv1
4mqi5LVeMKVlTJsjlsF9eOfsydKDkGcA1Zgoys5/OuDnhZdJjmwJcJB97y2cnocO
pIn6LuemxhhliBNOyJzpvnavmMWsxSw0OUHoQxGEaA6cHPnrInnoGbeL9DjEiP3R
iw0YpjqtCs7iCqXpp7FRivNDWrsKVhGbqlhdD3oCf+7jDiilNYxnvdHiT0qVqFwe
qxfLoij88fLFaSWh+njqC/tPPqJJIsDh3Cc17rnZJrdiFOs4pByL7TgzrdIhWiAQ
ioQ1+erRpDy1u1qS71+DVDiC2mhID7R6aLgbbgH7Jb4u8ceWImqdQovtuh+20lVw
j/ztLBDFhEMp7YkorKXJ9Fi9rdbwjxptOZ9NxKGHjHw7GbnuU5oGKoNKXRePUTdq
wunfmLo8P1ESJtqSvT6FHpDB9tHrK3RQxCdc+Zd/wlaptZc8t3UxoIIxHvwK1vLt
u/lav0I3DsnCDBBgSM2dS0QJXrbxvKxzs3Nf60ukSuK4rWhWCMsBiRaDiJsFkM0l
7uUkoWMcexIHBrxW9h3naXPu4DdjJRMB/zIUrUTVxmilJft1IVcs2z0s219av/cY
ReK2P0hv52u6ftvHdJjzKM3J5P91rJhtq+CM2nXTchmPnYdGu5IprHglPLAbQNL6
VNGXNxzKM0VKut0QxZKAz8DlXua5YppdxbJBDFhFEdcdYeYtgllSUepw+2MmjVZb
LeVkbhToFFJ40w2lHArf7skkbCWycyyaWSnv6QWl11xku34UCuQ/gbkicUsFF682
tq2vkv5l9jyHhI7m4tQuJbpIg7fNOFYE5TPBwdkJITZ34QSgC6Bkeln4sjp/S7i7
Us/bBb9QANM4qMJa+Te215cuPrjL5KBRliXnrew567fRB+uccn0aE06r2p0jNZom
z4zx5MDj9uE07cgJCEFy3C4Swx2SxL33s8TjNKGc3vJM5f/xjmbHSt80IyAOgXgc
4XmXOQFX/NSZNaLptM7fHOjYMyscXZE3I4aSGUjvevNUvrlEBXokz7Wx/sNYRCtj
ftVyXXG1p5ELX/4yTiviUjBebuf0w0cy3a47XzLAwlXhsf79b0gfo44LQgi3ULEa
ma2ZhmqcoQJmfCuagfN5PP5SKEP+Gp1fZyWWfYas0sCNh2eED2/y9ENxVKMpAB8U
0muQO0Z/AyUMGgrmdqjWdyUZK6AJPk6LVukYwADNy8rxNQ+WDSwtHeVofCOQIEfx
0a7/Lj0OdhULAKYo2SkFWuetxjQAicD9pHS4j17YMb8/y64a5c4YTwsJseCv94PM
azqVlOdBjx7eG1diZq76F4Ew9igHrv+tu5/3CWkQd4aXToZr/wPRpXphb7NMSuQj
Oq0u/dHBVgMfW/GcXulesFhSY0RRYb6TV3UpgFG3zDvtQYyG6+RPrz8QA/7gSOeS
YZWlaN5UBijA4QiJMqbhVqOT+KG5UwyojLVUORi6a4U+2ajc8Ph2fLBhTibxPgfK
Cr3E0LHMt3lBjXa/QCKPpHR1tq/WOK+Nr9pi+nB7+aSWGuXP0vIaakhvQ00hf2Eu
9cXyKChKArMYUuDVUzZ7ZnaAr3imnWxfBVr09Q4V/0rkDiJljo12Ac9b5dfZWsrX
bzWGtQtnxnE5PKEw6HAlWzYiKc+P84c09TptzDgkopR2Muy9A9dW+1xC7tB+Y2YC
41rkFXlfynGxf/flNsrtE8DdURpf9MjrIk9N2r2jvDSVmb87VO4J/rCqXqLCfMcu
jdLYdWQsz+B+jvhhmw6HJLfhRdCCCvfJ20AnAWJBpOUF6CFnUv7JBk2iSie3NfLG
XmqPxBqSK4UDosL4/6VClgB3xqdeE6PlmczstZ55mbM39tU0brdmZOEeSp1+G8Hy
bHfOQA0JxgNl81DJO18BchnVmqeFYF8Fae1hOLiZFvWYLKKnNDd1ioSLlXP0DLd1
E2WGmh3mZikOaKeQIosZO3muJ/kd0E0rbu/8Ed6SZO+Dv+Ei+Ws3lhRvjO2l2x8b
GMqMfUXcBWBBBQn/J5uy/4OpJD2l8eznNBfXhrb9N/4xQsmBPnSwNQja7+nC27Xf
QhUBHchlnQsaLDGo+d9tChJR53AVHN8TGfQv/uTuNAzI+AmhD+8bSzVOZr6/zklc
CaWS5x3R/nRXd058k5Il0IvgJGrQnN8opZEAbJ0KdZ7YmnxKYsVQux+5nhKQXIA8
2ZfIa/zlsh5QDk/baqucdPVceWgk5xSjO0xtBsXPa2bWKh1yPzJi2LxKPBQNJRkh
1zPGKn2sOf8NnYBpeG1pBcyDJCvBDi5F1NhS5cJ7TZHvkkeh4xrGpRzRy4Sox2zQ
ydPs3Mtv0zj8kXzr0qX5N0E1Gvx3T9roPnEFAQkuJHDkdAV+O/NzNg8Rv1isB5sH
XYQfNoLbFzz2w8HlvfGr6Rfhwo0B9Xz7l7A05Y6guKz9uvpyuWRkk1x/CyZr7vPP
YCX5Arw3JhVrXsJuYJWQhYcIWZXw7ELLkhJbVgcIJslyTzFB+QVHXVwZLS5VShDg
vA5jku7G6wWfxcu2UFwyRTy40YSP6SK7uAihQVez59/E8qzD9RcfO/nvkQr6SaD6
JHP5Uau/dszLAqz20Dc+pdfLeTwFrtkegeiM6e10KfWlGrywu7akRnEf+Aj5niPc
eXLqrFc2/YiCsl5imQ5mglvBBmRsist3oNI8GRsHCKWF2amnZbqGYIvK/XU2V6Ex
ONO6djo2nIS8KqIEhg0LBQ6raHH+QbOkg1Dk0nRP0jYn0B5UaDE56NuUFotiMemh
lWHXRXw0a1egj2DZXGBxdqmdPBh4aBEomwvs1cUpqxzV+jPT5wOnUZVnnvGjy0dS
gvzstl9wNxMthXVg3r1dSAdVsfSfTnPwjPEKQcA1GExAhkUPN5sqaBaFzH0S7caI
xgvnNJb8Heu7py2twPU0WIThWgjmOo4oSAi8mXOKQZTM/FEX2OelLGqSazuQZJ1Z
+GCi7G7xd/wtDmV8pJOXYxvLZEucUb5arbxW/ozkwdtgwNH27Z6pRI98yVyaFI3S
EiwJ/fIAkaQL0vkXDnLUXeWFjiY/w5GH+vZtD6NKWr0Cg1gKB9OJJ3qVKdVpEBr+
SLtedm1zwq+FvUYr352/piAxXoc4kq/nguOgbYjgeQ6BO5+MrxxQl5OpHmBzYko3
iMs6gtiI4aa0o4Gz6zBNHszdgZTX+TK8Ip8YRubSLkWJbmz80C4b3VVStO7Co1vk
CpDSX/yYq0x1u5APCHAjThiONeL+9UOQy6p1sz9gR5mWvTOrMaEr+tWtOiGJNJhn
rM3T/gR+TKvNZaQk/+ATSIrgOx5Fy3dw563yKxXiYlKYOdNQgxVU9ufpZ8Y+ECe9
HDasBdR2cZrrfuR58EHx4CPgzky5VYAXUJ9e7l0rSzdYEFNSfTe+p5OV/fhwnRMy
PWfUoXyZYVGwxZmxggqbgyOUW7J/uvEGt6r5bJjowigtlZtWL0+vJzeoZybkzB41
db37icc7T+2PiGug+buD3y60KNDlGCEiVu710XGp+INo629BZfy8A7/F1sfjFE0d
Jn1tPrUwxmtydD+KPikI8TqmNFzk0PtOLErtx8lWsootUcF6tMvuM6xDkwRE8JUh
5y9a/p0FAlQepGzC0IgRgKqnQW/q1SzJwDKTd2jt1dPKFuY/v/pZxX2ALqbQOYWY
`protect end_protected