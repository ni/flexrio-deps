`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16560 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10OtvJixhnWeYVQCxik57Bc96+XAYVSdkdiRVdRcuPqhD
KdUZklcVVO+PiO1z2YVyb3o7NOVTP0wVC98UiVBhuqMJf4CrvH15EeH6miysUokX
sJDSaTm3c5Mh3GO+Ol2r8L1yukaZkvWiehg7j6ttvXMXmHK/uUNEJvgJbBjBGRG3
r8m2dmRL3VQaT672FMihTS3xLVhfeMIfdScHMn7t0zpKQS2l0gByH8RyTgEF9LaI
03sIscqpUL0/Z/hw3wswyYMrshyjuCJb/za3ZkI0CR6fIbBF2jxHIFJsJZv9wR3h
iNzLaBu/2l62U6ZbP4uFyXOgH3Ex7unqA5u4mPVZ1UKHkp07E0jLDQh0wlNo2I+h
xNXvvqLmxjXAtRA/ZMlFkj0+z57PieWxhZziEexUuOzyTTJmBLRhvehxViqeBHcV
4DgDzgjcsnSCq/Dtjcr440V8MpET37FfDvMwnXubkXZZzC78g7kcVzXhDgeWXKLz
FLfJstErPXhk9s/uIna70Qqs0lefLg5Z9yDPVoAu3Rq2+KeucZWyXmNB9CACzhqB
Nlnaar9gW7WyxJEAHSK0LNaCwujI1yAlh/Dpj6eI4OrbP7R7y7QzhHfAxTabLomx
3moHtqWxUVNQzSaBrKWVqAziASzoCKERzLqkj/VYvgy5/PHLVd3V6sQZzScFiXMA
51idRefvXoZkJVF7laDiKjB2mOvEs/XATo7Kt+igqVkdyC4cI+ru99SksRYjIFqE
TJI/lUiHKNUDNl5smR+rzyd9E7JWP5hQ8vWvSk9THu7ianfDgprKGLrA9/fAiezn
oIMIWel80/6HL4RLIuuBLLWaMX2bMsvkHBMz/BDRFTIEwskH4mpiLHk7t3HnwSGB
oJDmITD04HKGUGbXKH9AGDzDHrm8h7sC7wKFjXASidcxpHt+mKU/ixI1aP6FwLB6
nBBX6W0+EUADLZb7GblACDJYvnGbdB3yuZPYtE6vwlWv5BOVnrZCOARzpyPW6jhU
D1xPU9ko6c3eT7SWHH7q7PBHV85m0qWdYYoXMhv75W2W1S8iRFzc+sssoIZ5pcSB
1kg8CrX6UIeo4rtYpT0zHe+81qh+uTzBL1IJL6+f42kB3nM5dfP/CCRJYWs9Ilmh
CPZRrYFkSixkGs7jBR71CZjPlkxb6BuODWQKDmZosmvk286101BsUa4xUJpmsdcr
Vy2Lmf2yItKeIiR1IgMsTghhsq/0YNV4juAiqHS9hMvTa2J/3FEvmo1xZnfPr1Gn
VUoSr7G2GO7QDp/K5OXjM2b86GO1MpVjv28Sd8iScMpx+rWhgFpb+IF0znEwnu73
+DTV7Mw/eksy5nxexIzmYrfZ5FuD5yF78JfalARzI4OuNgc8q/+l6Za7NkD/Xmhy
HUTtK2IAqCCp1jWneTy3yg6rkpSfsq4aWw1WN+YZlBV+J+a6sUr889LsxRsu1c4f
crERtz5P8XNdmWLUcfCzAn6RJMVGEynUjBL+8twPWSVvVSH8Uqo3zekz9tLLVInE
JLvrqlii8NF40eXZ55bypkpCTDhQpTpQgvOuOAoisPYIyIAuQZnNRmcgrdu7rTSZ
f7nTMYlvtwWhOGPmXuYOkmWTvwlTW5PGscEyX2fOmWsmK8c2UqwR5ginJ9rascFm
BLgdwbbaOa6gbt1bleGt2RHuQAMkjDdQS3b3VdglLCOBHoovdwRskafpcuy5hA+C
6xkqWWhfYdA07jC2iymGWu44o80svu55M4nQzwviM7kErHTHc5gnEfio0k3t3PRw
vrgn1KxYRHF3W3IN4oM4Wz4aKz2bnGrz652D8viAWkFcAuwe7UfoDn4EYRKZ08+H
lJSNoMSkXIqDYHvjAQCdO7oZPvF7nUbEDC2/GeqvjBWZPIMFYo7mognPt4ZT7wIl
J1GtGskYgIwKYk82kAkmdEvlScREqjwBeC7SHFoZWAs8b3kg/sSVdgpj25wolROW
KOurQa6NYSuc0H/Slf/fY8GcuEBHoOfKSaWMSAXayeOgxhzhHy1j+WVBMYIGROFo
6b2vNopfo+mpxnzASLibvbhSLFf2Tv0M4BtYQimUiQQagqJrNDvvUp8U/t1mGMwo
spPEm2w2FbN7znJhSG4JeW/OLQzB/p5F8ua7QoX7pbODp+TmiHvaVrJp5TlFN5z+
vfW1DsKD2lanqvVhxtHMgr/uN/4zb4KXO4WnLITlYCTD+c98HdgdrmwUZgtzhXRh
u0MOPV+stid+Wez8tXQzIb4gf04bMSs5zXCXm8HXqBEAJtMXALU+tR4CcKL8NKvu
glfErNX6QsxmvW8Kz3cgJCyEIwvR0KEOjf3+3+W7rT+1XHbK7m3jmvDW2sAVofUF
CIg089RPM1xO+73yZL8gUBGJs9/oI3LsrLjOa44LQAP3GfvZr8QwquPNjnGWrl4m
IVwYw3OB9rC4M8pq22G++jA2qoWDauTuNJM/lXWYdR1MYsNChzXjmUr6+xbKSFEp
27ogMCFPRs+P5nu8qU9XbLyNJHuAXHmGklVr8WkyvqN3sM6Cd/uMEnYUqv9soPyg
IlJYzx9TkW6IC/EQmdZFNlU5g9lKvRfXNkv2+M9jK8+YCPMJWzvWVmWvu2scE+OU
92IADwHAziBJFQmrzJBkegecjfHNC20jpjdoTAItGNRtBwhggBJIjnS0wYFdmbTr
J/2XkBOJ1l6hRj6h5FjbhIivOZ/im0XRBgL3bOsEgZ9xp1IovQy+Nrh6iumGFPoG
BYtOi1Rz1iDeeANBJhpxsGXtANCdhJQjJVliNiwfu/dlXwHmnTmCHVmy/cix7n/E
ild7/9dblx3SZwPwnWisvzpRs0vSyBzSPi584J4vrS8vMP2djZL+KBdd6+EyoiRr
BAQ8xaHVTt6r5bYHbtDwbYwh8oKQmpTpof7w5UHcED3NiT1CXNfvCPyKU/TO4qYf
69h5jSKjOjub1ndoHAxN7Km0ef/YR1mhvnA2YpNIOaqMdal2V4nuT6kYhHy5UYQb
gr6WY3TjaTnB1H2J30friU57ELCH7+i5erJXEam71NsFJJ1n64+itMR8rufUrHZx
beSUlYAd90Y/pmuPj1PTEiJLNCbZ5l8tNkEekhGL168defSD/N3kpoVq7LcH5ptt
SFVWO+Hl4EgaVoU8fSqbBaSC9UMsxfLAkf9fcsqVlikhwypRuYr39r+mDgh6ZA7U
6UD59Kx41upB6xI838V6TEhCOMQRsI1S5FnTIkoOXyLpZyxaT0Oakkzdb18jOIIJ
r50z4dVbj0/o/ljCasICOXZicg0jwiOcUeR6yc5FVfEFKg77A4IJsZ5oteWiGlUk
YkzTiBprFvgW045DnwlspPODeexa9ytd349mRPfb4lo0shPyobZdMJSTIBMkO2IA
nP+4w8U/+rK4W7re9fg05VEll2ioiz8SwDfhTWy2zptU+LE5Mg5TT82x+BTLKGyW
GESyfJC9PSBF/qBnDrt1BU6jKz4ARc3I+uZ9CIQSOFqpn2sBd2gQ2hf1cZHIsg98
FHQtNs63GUdLd2u6E1l15PTvg1ihrs+viSr4YXV8DFJQTiD5XsgjC8+Ed7LnEMc1
PRbb3nDVIsR1eluYsvDL6eSgJCdP2Rge1689MU62zKg44+RmA8aiIO3uWfmQpggo
5pz4n/5DiQzQlrGYJ2LabAwUbasZ6wKx7MXUBpIZZZWnyADzh6lX0oYD6L8oeljO
1sZRnS3WAOF5UZ6TjNLhMwiShpA2AnoVfIelnTHhHv0jpQofAK+mb7FCSmbcZH2U
VTPzllFFVerA4hUKpt1VExF0yk+/sSQIyTRXMQTmjymAp+yUc/o5NCL1ZlWdVnT+
tK+naFXzbfBTfhJtvvimQRYvKrFYx9qNHmMHWxqmnJOri78nvOhHhzsN4QXVkdQ/
2sDnBZ9qAAQFuRta3cDMxKV45VlU2oKX/jGij2gMSGg/AeaO3mrn9U3zDCGZfrZ4
Tf2yafS1/fDA12TNBl1bZnDE5dwqbsPxuFhQxhTN8V9ktOx88rqf8CalIAjD72aE
V9nIrK9QrPQsDUvMOkMFQJia7Ik6UlablTfmToRddyX4TJi7vyIS4J98ONYnJVta
UVKTERtxpq0TPVHSv0SzQBWgjTzmQ/+DPzvHsC+W8Ad3LxYNOJFTdrtdP5DMwg5t
igE3fLsWxDWTDIfNqlL/5Oku19PC9RTqRXzwZors8Z/zj1XBuwAZyhLjrYFpKYv0
IE9UaGOWeToUH7eLYEgEE52ru+fz4YvdcdH5PHjJ3dxLoH/Y+neQLxRYZqORAZLa
rC5bJeavua0zknmde5dKA+E3vwIRtqHV3cXSif/xhH4Ti4tBhCL2l1NTZG1hcd9N
+OiTV7pDF+Xl7g76ZSMO24r6M76iEUSCGj47gMlgiRPfoQyI1th16zSHah2GIV+x
3agU99DbZS2ks6k4FXpkj5k2JnAF3OqrhAQhFb/hLAV7HjkljNkgO/lIckOud0t8
OjHSqYYBgp6jlGWFofX6UorwfaIYVHJsRqx46GVlMNSVdbhWe6NpbMpHAUTqnw5g
231aYyKsQP2nCyZakZXHbKfoxfpbDU7vxBNV7kPiKcWaSo6aEgDYe43BTNxIqV71
87/12fHEIVORYhPNAW39WgOJjlEBaOmvVH0ywCPXB53QtGkECB6gGP9QNgN538aZ
3udgPF4E0GpTGlf70pf4xCnITNHppIEgX6jdmYvqMZNqD4DxgBUOPQMjgOR7McPy
VP8qn0VFoOs56CgTBQ4iZ0y+UjgyDxEzwxb5wxjv6KqkGfWrAXHZzfum4AqnDPaM
Jjq9hK9Vx2wGSbJ4KsUIjblz5i07OwBtSYpp35y0sc/B8wsgQjw50164OlcJVIS5
TLMVB5qPRDGX+1euuME1mkfyILAuq3yfdDnKC7wKlKed7COoYQVGWcUzRBYgG6m3
N6XB8WMegYVvH/bIJ/BJ8jSgqNPZdC+RjNYtEMb+QM3VnMq7wi7GCTSWF8vKtJxS
0G0zo3hfK6ZmemUmYCn8X8K9FngIGMqIS9FpQ+Xm5ydxLGuuLSt/pDPBLBfYuLPA
vnuvie9YUvk617xtySV9R6v9wd8hBuDiK68tR6oo/FEQ/sgs+j3wb5AlJCw4Lvfo
eOBxudP8HOT1JoXnMUMHivdjzwHsWHVb5VaKRgkPQ3JeE4rFWiPAXd9ejcSpQj4X
I06F9pw8wNnvA/EcWNgxs1uqWznSstc95+nkASofAURNmn0KebrEtZDXoVDxOihJ
YooaFXpuQJRn2Ue4PeUcoH+yyZ3wlFGXgZnab/r8wZsPKSIOvAf0VF9v3Lg3CPJk
VSVfeo76b4unDM0fhIRywyrEI17Wbrb+z6Y1UrsAPhdjtq+HvMCdlG3pMYlq2HkB
6PYQCF0Ax7XNNjQtUt/pNVX1tt/TW187SWKQx4O1wOqOCRNGzUEeWw46n2DCtODr
qQTBgSGkdh6sDHepAkXUpOAwd1MHYBlWdkLcGwHDi77gxv1ZB/uqP3DekRTdFBty
xhfWYwntA577hhyL5DG7x3AeUjndXM9TQOiS9/2wYpNigkGzrtjK2nWgYCqd46/3
1yBSu0bNlHs4uiiaoUigwZYkx3vc2V4wf3/ujFJlFfFbD47pZ5y3Jh3zTNWvGhjv
K7zfR+hFB55THlZWG/srwqRh9jlPhZQCp9UwubHAcO7I0I7reX006RtNtDd6gm/Y
rtSqxFvCe25+dK0qMEbNM0cF5SQO6JM17BexXjT4FqFpLpOPQuISb/PhvpPUwCyD
VDsulplcGbioKz53B1quFOMNtigwf1MrfMRtURTDMcGt2cHwSkYCCU23mzw+S0p6
KD997MigFaQjMYmcROBKz1dZpo9e78q8WYL4DaQU3dvPKWIglQOUneZjGzd6Npp+
P8tALrtlKMTQxqy9t1LQTDgJ6HeoI0Uzjt03V12NQZd80QUf1bsUlf2cS/tscsQi
uuWu8OdfEPJJCaHRc2QPPiyVqYuP3vHw5MZsbzqVqsb+mAY6ZHIUJDlBA2VN6opc
pjSjWaxOs4Q5naqnr2VvValzTlIteh/kQuuyWGRLFLw+uDM7ixKRQGMaK6HstU+w
sr/mq4xDlINvp26s1kQCkgc8L1wYWiVe17kTmGSdj2NZJFFuSsRmLKoLNE+ZJ9ES
O33jmUaNnwKCVz3u1hMuCKaJwh5RKNkOfYrYjhr0+eezzMG+uTmOHWGJ1lN4keR7
+ltiqNW5drkJbrNQ3Us7ak34pU/XXzCxQu1F6g6my5Eb0ejDu6gTZSVmGgCeA3Vk
84BFWa3u4IDo55c44evWKqcxo9J3FFEvqoNW11sISp/FFn3BUCTdl0ogOddtADXp
GsolM54iihrff8SOW3e75GokhOxUFDMj2DO+7SrsvX2ZsE+osjgV75oT1T1lCT7P
3i3aa0tnO9jax8yQI/o7JfMAcMVB7dfua5t/Dpo2H3oJhAz2v5VM29K6x0fNUhb0
FzcbpYq/Z0d4f6uN23M5eiVqHCnH3yuZbxLRSwwN0PeUT/UfJXgKA8mOjtpM+9jQ
OKedUY2CtnOd3Xs7km36uyC4vTeUdicWAS2KoLktjKsOilyyQLzmtl98uIQe+pUF
TcxOePP2fIv5HAX9U9mwc2JbisDvGe+R0oALzZv8xJM3HsT4xayAdyo/BUGYu/wN
JoiFVMySY05HqSZLM5nP0Oc/cF0JyYFfvF28qlbaiFEfiQhC60ycp6sW43gQcZ1s
cr/tJH87CeUvCx19dblw7Oz3gRMwxqDDarN9bh8oUUKhMeMS7ZGNecNjf65cMKqf
GeVFdExyZzn6svqlRjLRcO4lzBktBHWTnpvuvA6VnUAwnWdb33YkwOMqlDMkB0Fa
emPgDl8WV5KnIsgqzHyVqtwPCw4tbZ0sZxhNx4jQpYMVqC6moSL1fAUxMH6FKOib
j51nP696J9gCePG38xFNa0O3iuvdCm9lt11g7x7rHDM5PHPyzaQQmQ4tJUczRKy1
aabwZyP8agPz1k1LGCL/aatDPYlIJB4NLFolAI4wEnNFgqsBIJFgUx7Q1f6ni0MM
yMsvyGMDV/7nFZkgQwQq6KNql5Kof1n54kp47uczllEEmpig9P7hmm8o3ubPk7xe
0f110kBv1KZS3FqTvn909hIkSSha3A4ma7rgyS/Cs9X41EBs7Tm3RWEjMMm5QgyG
1wA2J9kRXKymK7uIh6T0G2RWvW+fNaF6rIBSO+ivsDNFpBog5lB0jMxRHYHGHsqc
WLXtJB5am8QMK9i4PpNpjnefz0CwtT5z/0Sd+JiCCxU9iyqgd+XroSqH6HauUb5+
pUAYA0NoSS2k5az9xukWQs4vegsPiM5UsgVwZGTHLyWErSZg8R07JcUcJoFaWmdL
neyBIG62drqZ+CKOR/RSmp7fMc18Vij1BlRIy50g/YRy203q6/j++FsFKXdZjrLd
K8OINMjqFvxmKtPiFXMVHQiAN99/JnYqBzc4oJP+bCqdXbcc9ygiW3lSwPlOd40x
lGK2FA+ll9F4VzuQ/4/RTsFWnFrWOgg+Eybht9mjGODcFXns7amYiOn+AK/uOetw
iqklbKqAYn35kJW2zSFlrC31WUaJImKdoe2ZV800elSnfxsANO6yioNfe6+g93BL
+fAX6AbtxESu/6pgFYNGvNa9QP70UjitHU7lyG5cJZ5eTd5LdXvjttSUnY5+0pYB
OCKc1IfgWrpzp7pogf03n4iNG5qAvRRzNLT5/4KbT8u38dtFSZ/NAjHyx0oBA2ho
oJ33Qli1VtvWm9nh0zhfJzyxZXR1q7DWxJN0PNCvFV3m76aojY2apWijr6JdfCOs
NZfAKVd0o6DyMDZEmlbfnXgy5MABpWwmV2aQVRxyLcweRSNfUmoczpo5NHKbWpFA
4/mjU8/IWTpIgKXruA9M9Ri7DKc+xqBkRZkYtqKCsd2q5Clrc9klzJ0SwuurlHZy
9pOaDgWY+ngSIirRWYAGWTQ6CDIVbtVSaqIcvZo/7jYw0smGek3voRkE+ni06KR0
5/CH93UQEVIVVpPdruK9ytfqohtkXW5lJ1l+K+Sdpqo0oXLEqeRdb/CmdrSCCevU
b3PG8yCn46G3sbwIsbKu8t6oecPj2NA1S10newf1E6BRTUSyAiUunzA7RSWzwbm2
kRnm7jSS6SoBIgr4GeWw8S/csVypTqrnEwGJn87+leJuB36j4Qp1bujyehLg+raX
0NvVZUofIFjwh9+F9bg9mzUWFXBrqnivlV8RbV++4gZQLrEJ8qC7LrzjnLTZvAL2
e1SIFfGhhRABNTF0llEL6omLqr5+impknVaAOFBhzJ8tTj6ECO4mG8AVgI2lX4S/
8LMRA1rgv6Pr4mU0I6CqETeEr+nUw1BlCwepdxCt06o7L/Stqg510HQh2TTzEb3N
HUW3cRaiA1Zen1SObKsVjP+kwxi774j3fLEcypLCio0/IktDSOXp6+ctMmkNbrIG
UKr+Y04+dkhCZVaUE+6xCbQ92uPXRGDwDTg3xFuITnMAfqzv3sPFKu8S2Ymlgf48
0/72taz9VDbSSchLGAJvtfk2tYKq2lwx5teXs+KdifXrO0wCnK8AOkRS9aOFKm9a
HXIPD8H+NOIGj8Ri18J6WHd+p2hp8eNbDmW6FtCvP+0jeWzTPlKQ7J65HGrNK9AY
hOq/Yoe9zYwiHsM2rU4P6eSD0B9tL2jL/cmx/GES8Z3xNcQAhL2OXXS/JuDLUKuy
G4rHwIs1orl2v0F8tTo4A0Z5BAlwVbdVrxcDtacg06KDo25DCDwHSfzFKow1GUqC
TIPM2l5S/XG+jXn8V8EP4Iz238ZOh+8Ff3zas/reEv/SqZUzbMjZB11JNmW3Z/+9
NRRbKX0BqiDMf8E6T6dsIRD1SRaJHlyJCY2XE0w3ubDTD4MEzhfQsq6nZqIhS7oX
crukamBkjEgun/DGcnKWuh+KyUMsM7G/5CLCDPe/oRcvFMuf2gozBDn/jYvrlWao
eA/8oDLzRX5OVVX6lLXVj91cDM10KtkpY1LwBjD57Mg5D/5yvlwQCCFHqDOtn3S1
vB2pwdFPRoTkOeGcoyf918ex/pwihpcC5DGFn2bIyG0Diq+puRr+wea2HSJv0eRi
1uWmwNMkm027h6UeagteTHVc7D1pFT++xjHo0XTdlw5qp/GNHIvtOungsG8hhqxp
krNfmw5t8Z9Wzi7XN5DM9Mob3UbDOotBwQ8uP4GBJIc3WoNc9K/nje7HZnj3T7ga
2KhBratVcSLVmDmYpM58Lo2wACu1fwrP7OspcaE3wNClQzGexNv5B7r5thjf9l9i
ZEq62XvAGjD6RGsA49ZdFhXlIms4lSP0kseEwHmT1buXtArC6KItpqJW7iT0QRaw
uGNho8gAAMb+TqAm06zZMf+QRnJ01MCiBIxrEZW7Bhg9wBUsl2hBQr89J2CCujmI
6mJT//VPlBdd7RdnoxYed1v3wWa/n68k3AOBvpcIDEmyItupQUFoydF0qNSjRI/w
FVBoGrKBqjhuphf5jmQIly7fpz0zBvsiAxFM9H+1xpqi8VT651eU0/eXHwkU/vb1
Y7rurGusb7Ogq9nsbWQvd/L4cwjPWTZoGr+cQ/6ZzE1dUaM6i01nkUh492KLdjMo
b7FMaEL1NKr7U4jNlnEIiWWIeHJEVx5+4AaKADxuzcJyywftpRGPpQEtHXedK2Pd
HLIiS04dNM5C3YPtD+MofUXFBvnZ/lklTLU0oNMEGj7otftJJsQTbnTQ6XE+fhKZ
2/cQlxURJfY/C+XT/JRX70RMsMsiU6g/Md0jaxeMGuY6ZII30WKqHFWbhnNzpoJ+
OufpPdoAbMlN1UXfZrk1xZbvOGkmJIJmOkDkWruNH9BWcoLxPwvxLfS65CwmLFm1
byDXeG0odGaLGUVYv4d/ToOWfUjEzNrYC4iIC9Yw3ziomMIYlR4HQNSeUscZcpzb
/4lpMCjOJBD3zMThRrMbwTy6rNDU+fW49W3eIlJ9saldbuFQMwsLwb9Nfadkg0q5
XUDLinEWOim0+iFczQ4F5N/LKqyql1KlaCeH/F4wui0J0CiZ3yFtJ+f6rVmHMfez
gCDe/eT8U1UraLb8mm1TgIBHtuMi/mXgYrwJm6X/tzMHbXynX6vNNMKRtAS11yY6
p0s9Qrb43P5RTELggwoizOLbfJA7h3VcY1/pzjNpacak+NPZIEVn0ggHvuc2Q7F8
b0XTOmIOCplk4eccPjB9ng1vU7ne3oiyDbLdfl9jB9nLzuzjUZPXJJ5k+mQTWXnO
zR+cRZbwxcaTl6ULZTBk0JsSyGvEJo0Ks2BcEa97/ymum0dHYl6TtWrqkC3P+rgx
rK7ih5DDurp+AfuoFhja+fz0GrjPH1Uy6F8mFuHDblgGAbk+INBiFLepr05JkURl
mIKreXvV8IcKxuypsx86hoHtksn0WUS1MRPlobYRvsxkSgWJHkyLbphtTBv8+g7u
q/FAD0g+6QE1r4gwssUsY3zdXd2+SkV2vC9o1sL5f+NjpC/H83AlAr9a0apv3WAF
TMLkry9cl13HKNhE4N9g+Cslk9JmrNoAUHQCyAam5I6PlQcS2u8EUsmj6fNVdihi
otISxiQifEHRJT8FOp88TdKptpTPrGP+dDO1QlJou1rMnA+Dpm2gAUgdDtfaq/Bv
HUZFIdltiIkbEm6H32HMfz4Lj/FLomdkTiGXFcZNc7oFr3Ene2bFvZVfNy4d72iN
NW2yIGKEgl7qGbsFNsyQbeOMYu9ko+GuqNZ7bEswnhjGz3tpRJXel52SEeJdxZo+
44sOCeMGwvjS1B4kwOrnusfl1aabkY3cApK1+ufBXAb13wJZ/3qCfuMkTdprPw5u
BSmNEwTy1fq71tLdt0K26DbSZGvQPbP1cioqecI5iBHNyUPbIhkZ3Gb++wfzXzzT
YaUVrhChgPYbs4C4Vxv5CWBgdvZSEJkvjpMNrWbk3xJKf/ppR9EuJD4X43RY4piY
+PoddeulambPix+e/fYpqEoDwd+7eBiazImxI5sIMNLXQK2Se1dnluBwgpHWjjk9
+Olp1lh1c8Q3GAHwY/+Ou9iocUkq2xcPjbxCfCW2u3drt4feAFjpBuIH5yWfj23l
AvAnbkGvjiwKmnomAW1OtbiBZHu8p/dIwuQnEyQmY0IDfrGGg5dO+5jvPHrEoZ2a
Yu/euRIR6T/knx+KW4Pwie2eQ1Sa8Wu8qINaputwquKl/LPHURFyUXGPeU/c/Uzm
6iE8erKDn0WUQKJwiYEaeDkmKVmrBjyuHq2HEoJT6Jwrd37w0VfqMrLtLb631qVA
raShlQ9hUbiW14NzatFtURmvW2ORVa3MpbVmIMRzVFW8mJ9N5sNms22dqpgxPFyI
dkGIADqiY+s8krG3IqXTfEatrdCaT6yDc9CgV3LVSmMKap7IEaYVEK/hAZY9M2oC
tZ+Sxf9FqUs8pKe4TqdWsbWr1Evh57yWLIU8LD4anJWSGY9ynWEP6Mb+P/7n75qX
BQXHNuX9gh09/IQV+iuHDoNbxiAm/9hig3xOWwjRXfJSZezEjkBrI302guUDm4mk
MsFe8LOP7UlrLcS1QsqF6/r/26nr0CiAjoF7jVOQSwasdNioc/dOSOXTkmYaGcCd
Y8thlecnGGWyU/ZjUPyyeDGFkkevzs40SEfgFuHkTMnw2B8yr5kQG9zwWaX+tCuD
O1golqXCQ3ON7lbQzVVsXHN8VICOaW5M5QmQ2+zNSFhFPNb+6gwJ+5J3gjT790FF
TFuUqHSfQjvEJp3chX4NqjKFY2fI3C9t8LDHwAm+2SHHkexsdbYTyHiiWImYhcGq
D3KC61cvzuNiMFMYF3TkApdJuwLYyS+tdo+w4WxlQ9rmyRGztqptmofPOmGUPOr/
7gglmCTFLZLZuG4CglkCK/cBWlmtBnsEbErSvf9Y4Jsk3wfMaIWMZ030seYwUdiN
/gcrsDV9BJ2yxO9q/0Cd4BBDO0XBVXp+IYcVrTqbmO4IFXUEZBwj0sFsjKGHTdxw
C0KSGr8WQ2pXUW9a29Wrjf1wwYq+hF9yheSvFwQk1YlcwcdLbb1QG1pzMQErlzaX
hUSThVF6u34oWD5jWTN0hmw7WhcZdrjy+kOHKw4jkMOcMnyqdOXjyBUOXtfPPj0+
VAGdg44YB8E5gY3YbOvNAt3xJ6YooKCtQyMdVx7INGNISNJJecgledOhB74g7jc1
CHqsg8ZoPLz5EGVZK6rPruBloIivQMIAlaJ0tpdTpU53tpD80rp4XEDvEklD6frt
J99QSUC71pwJ3Xg7jovNpt8jc5Tc7gz+LFzB35qYhMZgXuW/E6Q+c83tteTvns7k
9FLM9ECRgU4YY5msEVBht3CRZ+JpxjvP9koGATlsC2EOUi2DsthpDlxvyK2RYS2a
p9WKkk3Jx9tAdEsp2GY120TtuUddtg9onM1ty40cIaKR2WRTdNXHBpjVcWVROpKb
4nj8Zh0Otw0I/VVdskNOSCcy74jyfa9CGUcPq6jah+oLLiP6abLkf/mSJDyWdApI
dhpnvEk4hVatYEWsuXHjV7MtDiJoADdffwWK2iQum5DozTuIlbLYX0rn9bsz9N79
jV+MgJYr2v5yyviQ6h1MVF6bJ1qYH6ZOUuq69qztq3+mKUapRYAn6KUWBGimGlVa
F+YZjWbxIzb1o2wCrVa7lSk8bHvMfyHKDwnoQyAISqPf5OIxcJs3AckSiCR1JTcV
KlZA+xU9gFYUZgMFqXrkirVbx9SzwuQ9FNC5b6kc2RTC0p5kvU7wstuG7hNlZabF
mO7OEF0ce5QJ6SIh0tGevVo/9S9rpUHN6iPX6are8lz8elWeqPyDJ6f6VIXcyZ5F
pvfp/cEgq09NZntsP6BX+5jK5TnKcBJ9H2V5RcpG23JDAIWdqYp7xCjHU34V6Qda
3aWLZ8SytksUsFkM7pzRn/i6Nn7BA1a6qZkbEhs/zmj8YRiR251sheM874/WrJTl
Ty56eiHdwKFc22LiOA446emlWJvNTgeEhbp1pvo22Waf8QSKuH3SfP1/iPIctK4h
tWHw1cgbNWuCNWiY+IHV+vYe1rHI7GA1x3gcIM4Zui/inVLbSu9i0PCuwrmtNYki
LzNQHVNHEc4949EoPnF55Xt6iy2jwtNK0WJz89jC41Hdh/NfcCRQCQ/WmbuX6WmW
DjLTC/R9CY1jf8n64wFv+DI9aSRuHHIwI1uGkpIMXtQwMd5eKCR6Kqatt6u05Wpn
CZfOCZMaFngiY7xWhSodKAmFPjwj++Q0u7z4t+HuilcpXo/6x/GmnimVcGs1ztPC
9/OaT9vE+G9jDMM0QcVIomg6npSTWhEA1MeXDEoenuc0Kg59TuK8DUNZP+3N7kk9
gGuPyrXPhGUxxWdAV+XvltieAZzxoMDTvuXCUvMS7Xzh8bt2kthHPIjkaNJQV5oO
Kk6GYiK+bOHycb/cnK+GX/+bTgmJ5F5xl++4m6e1Ukxt3WuJfwaabyk3cuYmGIQi
pq6+n5wiAMizNVX0rBeGQdBzsgOz8MbFtDOvfyElqKy7FBPMptox0ewsqJ11Hdb4
X5vDaKkz5h9ZdaKXCGPpZarm3+RDW4WcTQoiynr26Z11qnPNH7fW91hj4Htztoiw
rcCrLfZxQdMnGPypZjcjWDlkeRyIFrMExV+kijP1ywEohZjcyW4DKs+PPYnclbiv
9aQ1MfbRvaD/v/aYhoeT/+e+PfpqZ9f5vm+L0dNTstiobV/QAcQA+6PBgMoQ+70p
iJPO49FIMNof1T6nQhnPT1uVxmGscQVI38kzMLACikWCzl5naBY6/EGFYlcVHn37
4TJsFtzi2aTL+Ovp5pmxAuBQ4lZRv07qM93RRj6Tb/JqVuIYvSrYr91nIarKwXVg
RqrVnC1CwstsJ6wS8Xj7eDxhS4nWqpp8+StBOsekVjWwU2f2Xrv/RDiU4X6eE0l8
5Q96kmSAw+4f9wVuPcOSW34UdCISNtiZ5vaXK1gAxeplUZxvuBF5421+CFVDp4cn
+knfeqCfIWKR3mm4d5J0ovKPmDe7CiYpMF4JDCp4Rq0xBA/RdnVhGhgAvTYK7guD
2A0PK+oKhJFP2OBLoOcsAgEYnmfzmJkJuNigOmnyp/upi1C1thYzDiwcM9QGzsSh
4Mxd3XVyggaafCsjx/g8zT/hByobS3xv4X/Nf7UjZXLn0D/a6XyHvFdjRcYu1MNW
geAZQ4s3T5o7sEt0ITTVdCPwsreZdr5fs+H64QLtu9fnCod5SeYtfOJ3Ed2BKOR7
NY2tuxgZsUYMOWrpOXEJdExQaS6jO3mTW54t+EG3T4TDCZhP/Dke33oIufrTodT+
UtazZ3HZdU9ncE7SlZ2H+/R4OBy4Dfnr1brz0P7mYcuKh+v+M79qjA/vaI9s9YLs
paH9M/C5weoming9Xz1blKlSnbYxkR6PCDdjGV0gAjzLiRT7D6lRBmq4r757aSuk
aTJ9t1UasIujfFDbVRhtMr+d/cxQW1FlmcA+7LkqZiL3+re57ssbRciivB24BMv+
xV+Vrh8kbUjza5LsGlzoOid9cHklMaOGqqdxdnN4Jj13NBKNtGft6/HYRj+/eQXi
NgGsi+JteAu6oNS5hM06ngUInknPhy37JBbjfV6RJhOjynxV5Esq+yJaGQNiAO+b
1GRs0JaCgO1Mq6k9T4Qs/7eFsRaRt4VT1oksY3tD9hsjMnrfqydZ3cJclL2CmJTo
hJ7ZlICY7xfpkDT2Z1mTQbNWvuVJOILJ/XqVdYnAixiAPb5oZdNoN6BulMv/JCeb
HBv7/InIiIYQaKP/TrgSDnO3IJXBa817usbtMJF9Ef7Q95xvOBbvQp6s3FIvmDeA
SOp+jKE5Um6SacjjuyrfH81ZpLBE99h4KBRdS8Fd0/KcGBvjHV8uqUHieWP4+zFP
IHVSpAgs4sO3iL9QSYAOlcL6Tl/wf4GQmwpLBhVXiDxi/Qi2N2h88Yoq/U4deZkG
dmMiQiRPMlwXzP7RWlGechUuvt9qG6JThLOvOKR80vD3GBNwv84CO7D8U7Qgc4ws
xNR1E0c3nDeBeOoEMO9WQeEjD3raFQvdXlfebumwEoBBgcn4ND89OehgAfBwrNq7
+/kNj3017Z8p5+vxde9OrlJJH2G60wQQSeq0agYDvesg3gKU0zGGsjgDQ8Bglupm
PrrJ9S3ArGTFfgOEyCWXnaPRiyrg6eSqAAt1sKXO5ZEvN/6xoXAVnm+jVksoScgR
63F9myKKhyLaA+bo3MhYYsEyRZdMwR0FBY2btHc8otbMJ4/OGhnbXzrh706unWAF
Y9wP50OnTlvo9Ep8lPYvmWjb1s+IVWK8uPdpygwVKjshdkJY2K6pI6UqtbF6boME
Vzy7Ayawwc/bvZFffribb4DX63pMOAKh3wrQb/YUz7Y5GJE8hN1yZAz3vajLJqOY
iku+LBZZFjViFjwVa1BxEcx1fOwXrjrWo39PgJD/vTeWxK24x5KQqdCTDC0ashR9
FxVtQmMjSr89Ge0aeJZTiS3GqgrvlzlLJI2CibohChUvLxYfUUf6MAIDk2BEJKB9
57tCMdZV4hXKxvAeF0XtXvM+vNbuSdnSRf9tJgHl7Vf1VDiyQtDvt4d/AQADiG84
jEEAZGsbFdogIytbGBmUrsKoZAoN2v45V1/bV13B/Q2U7+PGPdAxoDBq5paSLRDP
4+LRi5SwLOwCVzYsKtkhBxf1EYHVaQcq9oIpbUZVLY8AP+50umIT4SggeLaK1GoX
wC5dncHaZR2jEM2T9iTMo4uUJ2a2J2YlrsH0Y71G8IsAaOz+htHIzVgAQ66cXe2m
NhPMGnR+GULDcdxJ7iUIQ2Dyyk6Aae5HArqbkPYJoZ3fxPy9FTSCV40BxIfEb4XR
9MsSVpUSosLlzWTBIW+POZiGVP0+xQPgqmTAHBEAkiDUjphhWhaAjdBo7tI1v2h7
V31wyltlRFRM3ArVn0bfh+vS7MEsuzD2sr9B4mNHZ5tA9HV/2J3oPb9400WuslbS
Mi4fOGVw4vgSilxrSR+5RycHomRREDTKda/sSG+PnCiIDuPMQbz8zyUBl2la7vHY
YuhI6Dpzb/9Wa3Y0ioOxqpm+IlPo6eIorA1eAqtRGQEtdjYFz8UD8ru2fbjbGgQc
/sc1LYbuOhr1a/pcuWUGboRB6OeQ06bCv3uau66kcHJ41XOvzZ7HI15UWtKOvMWd
paV/QLPEASOUsxYrQr1O8Ip7p31hhYrlZMJ8rvGk3ifas7kTptHf7Z42r4T04C30
lwDmPshEUWo7VD0djH2+XjxAnArxeRzLQk1N8FKqxbPUznAYNlHgExRHyGhzaN1n
HgAxIN/86AouVxF6RVdtui26CdpyG3rXwdBjAYbO13lCWydXymi7MkjlHQBtwu/O
OE9XpEJAjvuzho68JRYB9C8BvcXan8vv2SlevLZZoYRKWp6jAUZrPzZ5VGs903DD
Kpgimo7xR6dNHiFTSnM2FeDlpY8atUtZ1qx4nYtXPrxn/DUH9HSSEmTAHUbipX74
G3jYHUI5BQf2PaYGT4XJT7J830nSiXhi+NNTqhuiJ1eb9hDA79LP1OalxPr9xkF2
9Hgq4PQfkmRBwGICXtNG7WpFOph+RBhwbcsFGCRM9oRYNLZg0+qA9xtTRCpbwT9F
EExE4Cq79A9S3OwmEglNm9BLvzfdtXk8OQf6Bvq+8+EBgsRMBwCFAe801H7at4gT
1TDe77uk2s4AHoWh+GsYvDujIFIB0cl29SmTgWCgmOrbVS+7wt4A268OFpXigGV1
xLp6PDj0GNwHa2eGhFVsezX2AjEK5I6tFQG9Q1nbVJll6BcN+9XqGen+wseR8qqq
opnzYFCJ6gm7bPVaZht7WljZrh5e94xA/lZL2cCIwQxlED96kNQbRPIFcOcuntVr
SgbbrBTT7FUu8ny37P8PEm8df3qzw79FcUcgn0pC6jOXhkuAmv0dCymbXxbPyxL3
nYoGlGWv2Hpm+j9gAqwDfxpg3CO06wjJSvc830g0tFmHjHQcnCRBR7H60XE/lm5b
SguA4HEjVfPfHny1GwsMcjJq42dWQ+xjxTW4TjeiRH+WKfdqBF36Ei10ew9WUsG5
S7ocmSrm3eRpqL4TQwX5rwB8nQuBgMw5xO5ONXdb5AYyp1PwiqUtgAAPrwORPV6b
ipDAOnQUjvWkYcXxk4CrvgoiOGy8dl4lyJMOWZYQRBcMSP7uwIb5f+jtljupy2J5
5r2zKxorzxg3y0T69A2/ZQjQuL3lTrkMpqplcnQF/z56D7VDtfh+7rH4kVyAAeXF
TDFARe0mDTMBBHUiT36SOJliigV4Rr1hSjuqrnb716Tudad8i/TU6wVlzmMzuI1z
UI8TFn2+itgNx1EHXHJ+5ak/UrDvtF5TJK7PJLJrI8pElu0uZeLv15gCMEm6Ms6e
MZii7PJb+zWJRGytrYRpqZ88alozJFet6jHW/Xb1je7TVi2X+WVM2DC7AQQr6bT4
1GY3O1grlIOSGaUVShHZu31dpMwSqWRADuhR3vOvkEsRwpcukxLHOSp11eJGVyRL
qMBYtsNNVnLlmHuvrYQpMZHl93JC+2R2yOn7Ab4aAV7eH7AyLW1+B9iR2G6Kjyl3
k/W1NXgQJyDE7EunsKb1CGRH5AXINJg+N4mgE24xnejR1+SkVBDMDr0FlAj90u3X
LPMKzLgZr630M9Da7Mdoa2LpCQWl0kaPk4HzlYEr60PT5Ay8kGfFZGm0XTSllbuV
GNxGlvvcpc0SUYFwlLcsbjQGEV85pVA3dD01yjE0z+kKSrkcOVkTntMTejXr1EvY
hmVU8sBN74VT+pyyvwgsKlIpV5aQIOYEhFKc/+DJtcCzv0ZAQKBtGz1EZU+zzvvH
OQdKfMsw1xvckBtUca/VKVOmKe6pRj7ltsYt+2VqbP5KM1+1JHEmciWckqXIay/K
nRw6i+cMPAUYqbbwZ/WEgN2i5knC7dZP5u7VI09q5nNlRs/sakszEjeoI9RcODOH
y+PhFn4SLHPbp3b04RJvSwv4qzaSc8epslyDvASIpO4W1wJU0E6ACKS5aSPmSK7c
7h47VBjtM3j8dSaPykR+epHI7PrkYVQpRqkQnKnHxYR2f/MBSMStud7b9DWjqjN0
U+4h7rEMPtwoZKGt3+7ywLFywy/M6W3SIQEcX8WRESGI4vZq0cF2oTH2Xef5ZlwW
wCdZ7E0mR9hL6DtgYn/GHkVtk9ZkJO32mvCKX7x+K3yeJ/tcnshXf+3srNPGExHe
08N1ONhgzJsPBB3R/tn6DpzeaYQpvpUScbNJUKuR5g5bLoaWcgGjlVnB+WYxZpyK
laq02qjQ6wKgbQlzHWlBSQ7rbgs7XHP7d1tbidKcQRl79H5BOgASt3ndwu/vo8X4
YUDbsN24ZfPMXxS5bgBYamL2FYzhJwLC2Nco4RiNK7PtgbUKhYxf6G44l7e/7a1c
vk6qxSx/iiyivHbf97YzWZfkcxQpRK4eNTRTPrIajYvMb9kpKrUERhtHQkOWH1Rp
g+NGjj79dUe0C5vofKEVC1OpD48EhFHGnIjxobiabgOdwlwPbyglIeVTASxi01L7
uCiWH+kd5llVbKsI6/DfkBYSu3ZBUdTPJeSfexUK+nLlIZ/fUE8cDVrj4C9ae9vb
KOkGDcDxcAGeMexTyPnUPdrvuVVJfWcvDvt8TUz1q7Yym5G7Ih4wnKDmvO2grSzy
Xwz2KOV+uXaZQlMCU3HF1gflfJ4Fqu3G/i/tvryJwoZG/1hvw4kcLIX40DY6w5RS
J5FXW6+559nkHMxRijmLexGDWiPyMU/XqR5IiLJ5tQOstpIJOiO8HwLdySp7FLni
mvzb0JxzYdwSP0/FDTdOvTAAnXURU42rOgKIjzNCSKhQkjVuEgzCpZXzliOAeAXg
zB1A9l29o/hoDUpnnDDClM52ifyOmy7O1ClxRdiAsX8rUQSxV0TK1HpLfkaQVtLy
pZ2IU8EiAvJKhp1NnRC2YTWrzuLj1QZxSbs/o9a41idaw0AnxFb6+NYOfjU1vyw3
R0ZJSVurdusw6TpLI5pcCMXoATvhvQqD/khY7KqyBaW+/DGyxb38bLQrNZreQRDv
g1wRmy8daaZ5awG1niFQ1PZwxdvG66Uq7m5nY2ffbSbN/n1DCER4fafwJagT7w3E
+8/F+rhVtAsdWWDQY5qEu+9YTt4WNVps7pVRqfq208dSORSyg64b1OWERhh86K9Y
V0TuVC+Lb7V9FshMfvnyveKX/GnGplSL+LiGJbd8rWuFUqReQ8ITi4eoX3Trhi95
1Q+kLF9xTvlZsv4t7JA0KCT3cGqPZILs9pU5ov9i9TyvLIh59hHPU1k9AtEsZ2uS
st71kGgKU6+yvAwCySYbNWPJX/PvzqH++4zZiOLJ+I5BN4Pdr7gNgeYjmxB07JiM
dr6uFYoF7Hzo4coSw8hhDYedHi7A4a3AXoKvfThMx54iG274FyAeX2hIo0jCYmWz
qMv2/Mkl1QUm1pMYxNU/5iVJk5AYwHRJHuK3T9uhCqEdX3iA5tzOTaKgQgULeM07
qw6Q9+X+Hns7hrM1SzdlNEs2Waf77kk4mNXBXFkruzL9xajYXwUP13Zs/VG2XwOC
g2Tg6SuJVbfrrqUT4lfnIE7wQJKoVx/O3E0oVLEgCPwvSqGYWzJyXqqjIMjVuAQF
Dx71s7Gf3G0jojRmIBt5nL1HTXzyPAp0rChL1oNSi9SHcjS7Qt3uI6Sk1TCLrfLs
LdRjRVDiX4trN8UY0CJd5rJ3nVNlPZJEci15k2w+jamTETpWyKpHQcWVgHbGbr2s
zaESFrPp6+QP3PAP1uGRS7FT7qJI+4K1zXgxP3KEqqN1km6cl4rV1of3XJ/eE+v5
N2h/QPhMG4/xcfydWNdKcB6O6HvtO1E2rHfhTFdi3U2PWcclV46KnEuxPiAeiAbf
9YsZfY6Rsd49eThKwTKKh3QltLlcH99ZEcpUle0fwfQaZBLOcH5FGgEMnEbSycYV
XYDsDKsNYOPBnyPQMFMu5sGrPlsQl6liEFuXAmb63zAzgYan+M+TSfJ8IH2wfoqM
E2USEqiwTtv7iqCg4X5mSZpsoVbZswfUjafacRQVbqt6i8mXUREvCLnBA1pPAUy4
qWUW1j92aOG3t/lglx9vf21/DXZngXtvg3SFBSScMhBgNw3vo0L15CPgrKvzIzsc
RNf1ZQSED6cXRd3zZs1IPnZosVoMZIhXcqKkC3jZfwnz9QVQ87E3jEJkRYVILDkc
dJe1dkZmgpDri+NVmx8AcCOxnlmReeV3A/aRRu31sY3oMoQk/zVxwySutxaG+K06
pN4MsFVp75xC/x+QkOJNgWWbV0KvI3ShhAF/yD9tqmedMy/RLHtwNFnacnxS9e7x
81Xh/nleu8XHf00EY5Hc+7NN7jcXmkDokHogKzTCPWM0UsZPyUp2DQ6/7p7EgqOb
AWLKNGBif6uMzN06pGFKJH5iJtbO8b3gHyaXpPhfvD/kSb9K2maTkOUU/85shsa/
ZC3O4R94MroxLdRk9URgEsDXMuJUeXNQgWsA6xWtdx0vf2DB9BQr6jgwQPcUj1w9
B70sz1ZF2u8/Skv2WHFxVTfDvuARH1vEpmIgXZchGGPyhwYyhNdLO4GA51xMjMWf
xCvKRh1XasVpAAg4dP4AAg7JBPwm+YeY3d0KGxrVy/aeWSU78s1Sk/mwrpInYJGi
xaNC+a4tQUAPN74+tcpyEU600k7M5jdMysyenk/s34XeLu2o4zmhNsUUPKAcGsnd
OZkmmjk7SoHs/FiDp1eiYcj0/47PXqNvJZrd1+AmOkeP3yjthf/w7fdz1WLi6Bpy
23uSON9Ahf7x7byCeCEjyBxicw1QxZIwuT2mbtzW1/XJdtIji+nNlOFdYG19Asp0
y+OwzKjob9fEIHjZFSU1fxgb7epr1Qtzz6rvqwYnpUYAyTrOBPgw/efVp2PAMqHN
L3XsVsUfZoLWKwPQD7jbJFt3NeIQNvwsj4VtG6MVMgHf7hRQlsjykJi4hk8V4AUy
ifaZ//HB41tbMjPTss1G9LieiGBTgNj7Rbu84fXazqxdVFeS9eBj9PVesB/YgnxO
1/z98riGnizDKWigqfAIqdKomCPfmw29O827afSNHGwG7xImbpTT0I9duWmuiQ5I
sF6wAF/HFeE/hENWxGMiRJEaI0RGUF+w2I0yLYT/TdgFyGift00C+qB/2z9LCPzA
0nl8ut0nwi0fcg3wyvX3UEkBiW1npFxmQSk7ydDOWP2U9KgDX9i5CaFHhZy6Nv9j
UDWSLeUf6pEdsxnyJwa3h/qtcssHQXMc4QCYlNVFrUVBP8smScrtMyH4aQDyFKMK
5UgXxU1VxFJ4C9fLZOQT6htJyulY5BZsFeVxwAkMnVzmaljAvg0BYzJqnMj5dIWq
A5foGoe9fY71FkAqZMHOpIeeO3/5DpjYn9lo0zXWcVix1yeuL6FShRy1TdLCzvYf
DZ+K0WCZBxH3uzJyNMD8G5gOMAnV3vTWcIYeomVgIlquJboSZSs6OJjOWDpTDia7
db54bK54vo1aJya2vmf+0gVSP1GaslRF4wRZTYZoMyUViU0j18mlvFeMUwSSeED/
/CqKcCTWxRQj8ACHEr697sjPigSBnSLijjGOmKHmVeiyvL8D5ce76qcf2HYBvtaY
+mYeP9xLiO1KZnBj1I/genvX+Y+n3ceHsjiMUPsXHn6ca7CqeY0pa2N6LD6Z4dn2
TeKsrWOmPraq648nt/mf5eH/2017g2fY4jZdtQu3fN+CCm9y+PgLoU6g14Wuk5Hd
4V2UMmcER3kmLAsPPWiZLESZs68GsrcEYhJx9HFFNeRgfE/xZ5MHcuaFSV6aVhjb
d8AlfYg2+oOMej+C0sn4kYxJeMzRsWwMLqlDty3F923ugGwhI4vDVA1CEWM1IXam
qIiJ00A19cAAnZwO7jT1lnH3HyQ1MdjWhvKWavWSMQ7j9XXRoDnMc44996acVEzI
rknaJlm70fPXNGixYMIfMTMxapqvcyzWW96p2q/dicllIuziDpWKlFQqiL5tA01a
`protect end_protected