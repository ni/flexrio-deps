`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6912 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
vwDt1LQ8llo1bkKxKo4n28ptHYzBbqLyhYPikXhKxNqt69yQJvAwGZR1Jd0hsQ6Y
MT3Zrbj9qBucdiGU67CleDx2WhCPgakPHKEOsLohrwgGOu2to+zG/JJS2i1tUCZh
E5tvTUM2UU22GO4iQzDErC2jMrKtLsIErkdfmPZ9YDpeHs7iTFZBxfym6zvsixoD
JURONvedHeK5DOkxtlvdl9X37L7GErq2AATOoSoZuoyq7QqtaG6S+x8nXJwmj9hq
4nQy8U6aKngKsoBS2JniJ4cyaiwGJ+Ds3xF7Uf8i9SgrzjJNqfXwgpLH2FTqTGd2
Z5bqIvs/sk8hAd0zgDR2km1FuN0Pkg0d68eftDFIoc5zuw+/2OWvyipsI+C2Xeeu
2fZcDvSbW7tw6jXS7hYqEp0Ng1+3lpRp4XMAH/mYECQFMouRXxtTOHJSEtyqwCRb
mL3RrH6wsSYsSnFTSJmuMImElUcvDuP/lKHuThy9ycT3WflwdPx57B1v07bViPqc
uCjfSK7kCJ2I/PubTrywVrw4etMmgUn+HJLXn/8dmP3d/gf+kpJUipdM4XOkwnCM
JCyhcQl5S6BM+WHspkEt0dP8j/t+38hxCMhzShfLS8kC7kdk1IxF6cbZMP5kuSL0
y2CXGAWgmk8ZD1fBZW02xF6X72SSqkZXHj3ezZhBKV8dvXjT0lifkqYi050W1a/7
HS/+ZBto7KcDIHv/aThG4s+TRXKz64/hKNtocNBNGVbIqH4WXSPyJztoh+nlR/Vg
4fG6cKYMuc0HozflIuC5h6Mngb0jyqLZmOU08apYhmy/CPTf3GGjbm8eD81GBI+S
NKy6ogNaZp4f8J1aSeKnjxJ8mfckxaCsQymVIbAb5KfgcwTSaCQ6fnyGXO2ekrn9
HSNl7AulSzec7CdECq97djIOPAtiZQ0Hr5UNfdLCQFdMv8CnEOGAv77Y0jXSDlrv
Epzh5x+CJMajp6rxw2HfBAOhNu8VFlQ2H4ZvxTq60IdV/1RZvZvnD42HALliipx3
Q0ZKlpQTjQo8zojBOYVALQTtjm0cRm1q0nU3Iv7wEOE0EDbtiIg5yg4ICOfznDgJ
YXQOliRkAjPSuuRdUbZCgY0RUhFec7GW1CSB5a0lyaWSxdOZesFTYdTQws5PfZge
Fu57taZQ/Czo6RENG0cWs9cVuX8wDOM0M6U0axs8w/k3nz+fZrodOaeQA119xnbC
3jdAnBziy/me9ytpm9r9U6LzCWGwbNNTliHmOwU35DQ3jwdzpPgD4BpTR6LhwKK8
oGV4Ozhic1gNLWJuwsdCsNvYOQ2u70VTmPCxjQXK6dhhDPDUNBY9EhRaG3uJfQyF
C3uUAidMUg6PYBMzr46LAdlsquO2AGji9NvLGyT/fikfXPC6pb5jTNkznBBEIWH3
DklZkG+4A7aKLQ7chJseH+2c2eK1JrNAl4pVDQeBCrfjGv8tovBsfGfYmQ4KGCtH
nm+MjBVHpHg/AI5PnZPJs/8KWrnhuQhq+B+uHST2X7VUbkuaTeqreD8M62VsOhbr
QWgT23UkjTOJtgRgx8SMPurIWOYf7IlINoyMrg8le73++hGl43fcPKkmHVfQZNP/
bPgDnMZMD8fFniVlSKnxpgK04n1Fbrrw0orXtdfhSrkKlwE0cg0PK+/aDJgTWPu/
57h1rcFV72PvH7BdZrGdeYHFEuZ5ja56IWXy8Vhc5/7S+5jMBD1dnKS4AwRPgXxB
v/pAOipUBzEuMeZqzFLxlnd12ZGphIh7VvMW9/A3TEUCw/b7fCwYca/ox/5AzhtL
cnc+tiVQJFkrwWfGewSmZqQss14P/nEerlfH9+aYfw2dmIn4Inaba/yl7a6f2p4h
ApSfB0GENtenpkB8MrFY5ed2a3i6bvh58FZhqMq/wTdFGrO8966N25XQYwLZ8LMa
84224HEULx9C9gwVO3Qj2sxePw19Vq/CnLTkHxJH9IWkNKH7mJKJPPLyJ8vgr7cL
/TZFNo8lJYCFQrmcloBHBfTC22F24b1U3oacyYB6isDSzGqYs8yuOmuSoIlrpt2h
cNtFkjHpNi64MkFmtZgw7dopiJELFlcs9QmWNXxPofC28wd+yRNgE64Tr/319T4M
x3XMkjwOnT9rTiDCnRfEY+30PpeFqsSQVIqpKCQwCDHJMKFx70H84/aNzHHBXkJJ
cY9PQrEFFw8zA77KHvVf+8487hx8if5x2nFgmy26wWKYzIJ+yUqiqE0hXbzeMNN1
B4xj0g6LTSVB+w0mxaBQ+zvcA31pmW0DNfPD9GtizPYtkUJnyCdzFbrfookgF4AR
E+XLA5kBV0IU85gP8Ndq9QHkWuRvMZVAjpYanNbRBM26U6T2KkMaStVcRNoDXPKw
VFD5+MaWtIdawNvlsecOZdreXlPgge1ZlgsWH3Wya5zg9eHqQum+kTqcNTjIW7b4
MFnWjBAEKAjyup1wlNxfIYZ1+xIaryGi5SXCXyvfoNDqkQjGQGhNIKQn8bVuMm1a
p3eD9YmhKQZjygH36ZNTsDeSpzohjOsh5mY1elDsKMbuvh748flMAa2+hysX8D55
PJZketEGc4XlsY9W43F7mVGb6MlhxOFPhlN8ScvFQ0rbZgySzJQow7X/++1nHBoe
XiqMoinNQ3FY01yNQFBLrC+2I/1RHLHm2HW0ffX6pZU08Yt/wOzkPZrtbXkNVJWD
/0/fCNuu/0maqr3JYWmb7I6kZgYmrUZ5Gm7iJD+ItMs6BAtZOoPij0yEQcitYyvk
LlI2gL0l93J+85mOeCi2wtmZQYQ5/eTTQuZKN0DuTSjSw6YwSgJC0VI0gr0v5lWK
LwwTPdtWbaTlM79sRP7ElGgLFBB0hZb0JZnjgePPVACWCGPY5ehZG1CM99oxgccI
BwrpKPEBQRrwtgLLhmlxoMoVf1Qmy4U9P84toMw/Ed0z5styTEpKHiW/cGDMFgsF
42sE+3eJEybQvSrRu3KpzwQGbdkMbeeZNMnWxLwlBpGPn6lruSzx3O4xyCQyGi+3
gBv/8Rziq0wXwtrZNRBQjon8oKhsAWIZpjiz4fvtv0xJt25wFUBWfY8cOXZf/A1W
oNY+Ku7XEC8a3VbdNNkGoVSA48C9vVpEFC2gqX+ne7uIguhtKhnu8O/dWJjeOovB
QZLvZq4xHDFcM4qCQ2HhaOwEWX2YciSI/3PXQcNP9T0Z78+lB3rhgbGRQAzFuiRw
eBLvaeNsTwhws1vRYM/NTz+Ml/e8Qp9c2xq61c47r2GYtVf+t+rRg/jYcDARnd7m
ZgX9HzAn/JZWimDddQEY3UwoxNZBcHpGeIU4QqTbxUPHwPtulft9fFrTkhyRDfs2
FXewGzvSyO7Ol6whheBfRJVb2uPy5tUFDyZp5NmSkyvee5phaYwpE4kpVtrQ+X+K
IlhSA1SIWbVLHEN8vLV64D8GZOa3pgGJFIQPImhxfUDdgF717WtTSMBzKplJ8sGw
QJOlBynuE4l27Xk2eLHrlYBAi9SoaQNe/Ast/IrFm04Hc3jmbxVbKNMHtRkdK0aG
VbZYnkWtdmbCo19hRVvu4T9U143XG+2aqWSaDuhZSCu2pYoemNMv+/0UQ1wfGqUr
CC2lQO5Bv8eklweiE8LUJoZETQNussSqnlNr3dk9YbTax7+VISyc4Xvb1ZKwQS5p
+YzYabSkH3XiRpARKniuA9Gq9UhhmF+gpiRvjhEBs87Tptr2HtXg4AeyecElS3cT
WfMJhYD/jFlUxKvW6aeyrzpwtzpv+5pCO5zBBCQ7oLzgUTROZ8APoxKG1/uFVsN6
TVlkzPDdcUzQUdzpVNP//GgESopDY6Mo26HXJnCmswhj0dD4WLsdsuEGBdtApPRy
wTrR4rn7suM2TmgKf9mdGKxr0xOsT2q+vc3cHxRhXCOktWxjKjsMa8nShfSuh8L7
Q4B+VEqHpNIjViXHpsJsSrIgBHw/4FziQy8TM4njlmUpikhf31RiUyUYROPYA8yf
4DMZFH/aMvYyT8/nkLPPwd/eCMxfkVVHY5fXICUQfoCd8s3xEWQAakPrghtq2D6u
X0KEXT/u6hmA1WT1juFISxxoc347tCRvx+XPTCTlQPd+h5g9IuQeYbeOe8tdOrwh
xA7qPBuJ7JlY4X/INmbwXr3TE9u/MOktYjfK2rjTeQ9KhkVAt+j5/4X50Q3Qgz98
r41gEaMXKIir2frvWgYOD7+ZSDAFx6kFSmxm38J5lH3JsoEhAGjC7ZB4KG8PBGzT
k4r64JmkuIUyo8+lWtIvcihshpNRyV1dwWbXNgkJ7T1J/ju+Ln3EH/uZdL4Ny7Lj
W4nChvJK6gnR+fCh2oxkswIa56zQzqYkUUoBx0dECbsSpCSGdGtwLdBu8qG2F95S
fMU3W1CVUuRXSxiRxSQOlPRd4jbi6vrIf7DyyDStdaNxtL7JyUEk74+HwcBzr9MN
YJ37Tam6lWAwNX8RmKB9eFYmJD+mIbx0lUasi1r4jMA/YyMX/1C5amF5RioGVGkW
xq5mVqBocg2hQfxMIgUgrD8okgrkRLr2WdlOqKcuPdEjfW0/my6m90+B87jNLPFY
iK9pHc+MkMpjuHe048xtRdOdpSMLQrDoJbgznTYTbCHBYTNyWDF36iAi+mZdzEBX
CoMRT7Nbw/CFXANlc8Q6MZehZO1MGT+e4ZQDaSBPwt31Tds9zjU2nt89nR2dFiDn
mej+xiYRZRMhK+yuid5tKZZm6WQKc7wKUCIk/LDz2beZzqbiBtzJwkcTwIaqzvNl
9vtvsSLmaadwUfhbq9gKyqh9omQUai2+sKM84+5riKcFRuEDeidObUdNLsrPWGsc
ch3BK2huQzlu6/lGtg+t2H+MY4JQgbn0INfchOvGMN4PymgWKf9V9IRfstX+vfUa
JNH788o+Ie3H4qnFTb3fhxMgB0ysCJaYqOldg8JHeioO8nv4MWsU00MEu0q5slJF
bo5GFT4eGeCih5PRgljK86qgIYw+AVAWjtNCMxkM++t6MuiVJbMXCqJ10kihbrNj
qPhtyCRE3UcGiU8UWP0b9WG9uzWDiLkp8KY8fFSePxMKxgF/dFxYA2DxDn5GVwOC
yirXt1aHUcWr2UkGoV+CpG7lVxpnAZgLbumNIkNLBqqi2rb3ntTla/xebJVFV2zd
U79YqXVcu9MR9G6LCXoIHSs03bdElE4g627ZlP2dB+bwQX9D3e9qfSIcIai69DOP
lglBsjkD5CNvFMYloIWv9pJGtav470C1iFWhiFeCTUWZ533wA4Zt4mfE5zPNJAL3
eBDkoWxN6z3m1P4LHFJCLeYqwCLkVx0IYlfzhtqrqBIZK2HhLoNavhCTWKIiUujA
KQvEbolRD32KPVbe5NM4AcnWH1MfeBqEQNg1xOFqE9ADjAAU0cqTxRRM/vVNbHsi
9F/rEu5RXQIveWJJPyh4BI3j4XQLjThqpkY7+1+9rFT+5kferMXnYRCBHxFGyp9I
l7BBP/x2EtQvMfqIEtN2VoUmu0yFgsjbG8kHB25amHFoNn8ylDF9z9EbSDvoXcCi
th+s1N3WAr464OlpS4wa9NzRs1pW2MF5y1Zec6oWuM4nC05cJqyd1FAHdWEts91Z
btXrBodG065IEcl2X/nsiHY4g3yqL6xzD5Io6J2F49OO9AGYMYWgGg0EexyRtPUg
QrsGIeNt1h+4qFu/8ZymJladVU49h57UyqP7evnTtSqXmShUqj0I6lx0WsAiyPVW
ylfWzKajDobYSNIbESeUqhkgUufefDrzWWlHJqQ8xnxAxlc1bZcOetmN3rg5ejS3
rQTBzbLXa/IqzNnEMzkMWgTFN1/KiH/OYq8B0EJd2k/Yer3EfoJ1Rf0p3zM6zcRE
9GfrX75OgZ/P8maRk9GN9PrS7OwXXT9mwhz7fqgwA5jDNckVZ08DACysbiRQkBwr
dEKexo7ymoI3UBNu2PIejcODO/c5xy7clv01atAlNOAVfpO1AWaT/sO1Q6iSYkMm
kQnXeAXbPJ5nhrZafufZjabwP0oa4g39HxQce8H9gj0WqTvb8H7K6vocE/5PqsVR
7vXTJ0mQh6mEBSpBre79NxmPgf+xJnNyu8GgPr4u4E3jByAA5wEzL0E0d8b0K4hx
U47aGu9d+vkZMOsdJeuLRH6V0er4o+V5+z/V1EfdPLOqs6mrf09YH6BpZf+1oAkQ
jwKrj6Up4GC0QGCFjcs55nnrVuSvhNixuwyKb8DbkLb7sJH2mX7DKPEVTzbVjg+Z
jOU4dKxo2IWGtzEsnMgeN17Ng/9TvHcvea32k6U8OUsxUkBzS3VZVXD7xz/HLZLi
Qryq6VfFrzlrk/m4lvUeK+KM7yCEY+4hRUo/2yoLBDkECU8pasihDjSjgkPEcNix
djdc5bqr3jSLIL9HeYwP550WwD1YdcGFHwBJ9oKa13Q+wMyROrLD5wUVguEMfGDB
738ayldt4wNC3j4jyTqQjw6Ykx3CnWxWoQQI9FGORDprC7rxLJ7StH26QmlwHh3U
/VFylg7g6dMA1BgOzHGAIcZVoWQHqsqq/Ek2xLc0Zyn3U4pEyHfSGZmRNBp4oKjx
eX52GOEKZXSC+8NnL8fCVXCUVmSf7h2VCvctaJlV9mNfKkRm2rH2UH2sO+VEzIHk
XA5E3UaOCEwbNPQPOVhoIfqV4lkYsFnQqfz4sfISSSF4dF+mfc4xeE6E/h9uEiKh
+Wc7EgiG1Ljzl7H3ZwOvoW8vXUYS3DO6RYX1ZK6Y8sYZ6qs/jRv+hizZc4yeC2ga
VqBdNkYX5tTEiT+AJiFt69iJQMIUGR7pRTeFy8oGEPwaHV5bypsNIynBaY0qFlxT
hDQIx5zEtd7J5gOPXt01IrmSEMBIVqtRul9buLq9q0AYcI9fWkKpwr87nQw1BqTv
h2Vrs/P275IgMNTQw2qzeZXQAyYXrcv6bD1HuPp2EEdRyPnkvIXdB5zdKjeYaTns
wdegQcw1qqbOEr5GG2SUMGyrSwFNTarDkKLfT20MK1iL87BSVJaT4zE19I/SxuYV
Us7Slb3zQ0PvsxQQ4/ow0nbi2hMBTGQERs7sehPyKtWCSPen5xz6l2mlPyiC39jE
iP1+WL0nAXvoKQOPQGpLDWD0geoOub1gNDB8rmQ7p2kv73nVgJ4diZibg/+nEed+
au+6W8Fnj1wQQe7Jd4D1NHP/aX9Q9yZ2cBEm57G8y2JlaAPDSpmT2sJfgio6R/Yd
OplHjhNjjMeiEwSNtlWI8i/VPx6x0FAJlKA6Vv8GyRnY0EC4uHHghXEIk9wWstfA
6iRMxD4gZ+t6dk8nybRVFJieIyPDTeLHv4wg2hVZoqkhurBNrEhJM+62f/o8ZmB0
DNNT+Zz255eUjVQrAZUV8TVVw0Lsz2QFdMuY0G82pIM9OdRVU589U+eB/c8kcffI
uVE40ckJNHpgVkQ7JlHPjY623XHXMRJxj9A9cDbjxGnmtgLuXnOXMjiE/RhcfyDx
iToy+zmoEFLaPYnKvCJbEknoOaZ2gzWPwm5KcwvXmgRTRKWvuCZxYPCMfVnSMcx7
z8F1EPpnFT7Hij5MG+rEwA4qm/xKF/PVyyIdrpwsVAoK+ktYRLISRXceB7FTv8ha
YKBp7aDIWm0eUU5xmgYYqAxuDpCyJc/mTFeREmt9VxSPNheTDptNsJNBXg5GpVI7
kfh/ruAtXdSpTDO4Yuv5fpATvPbUJDcWGvzSiDuNBJUSCh9EQZUiKwmubqbRQiHd
vGZpQ1tcqk3dNJAgUH2LuGaffRL7Pp5NZiRWKOGxwK5bQo8DYr6HGYKDk+l4zI0u
HbLY95dbsd8uulvSP6qGwQVm1uMvg1b2FMsVsc2PEpA/m1JJ4DRNDIA85wHUdU2x
iIbnO1dzjLuItjPYwHX4TWy0fj256kxNbAMTC6PU389qiWfT41R4Chtism3AFQRR
Wvjje8fDpMr29D3/4+ImtOOpX3+OODwG3r24/pvCTlssHHZfpcWVcZLOq2b1PmBs
y1JHZ8ZzTnf7WAqTSau/+FStNj6VLI59PPLeUPdG5BRM6GNFyne9Btzn8TnBWm8X
GZJUC9L0f23iSDU6LCPhZQr9G8nkQFfbSKDKHrExvEPB/ZYpryPgpR5H5pKew5D/
zkQANahM9sZ0ucPsvvlDMyqEkQubTZjOGlgCCQbYS9fjtj87On4LUslmz/Iwzq4G
LIvUsVpysU+6sxYLdx8rWFHc0Qz0K1fGxQe2N8U9Ryv47+Ho7fvTt/92uauDnvlW
SUFW9tevADGKqIXiXzmwvZsh3bHFWujfxmueX/THYvvANZFXoLBNuzwhwE9SC554
Ss/C3E8VlAkVFna+gothNp7v+Ql1FzqObkwqm/AvAuO6roSCc5+DvyHeK9bPNi5T
0bifd68mn0WZm782XQ2df2LTioykbmU1KFpZ72LmDD49vzuhhopAIN2UCY1syenj
sdDsQhWIlI4HSs6H5otlEy0s6nwTkOrbipXCTIJeBgZpsJ05Bu97EQYt6pqB6vz2
wfc85JEEwEqmoOr0hoflNhnVxGAvxJfob968YnJpttSb5bZZMFdjIqzqRm9Phmye
ZFcQqP9cQ0Lzvo6EO3j3A9e/DoUh+PRoECsQGZAxXkqkeYqO5R8Exi/BZmqhD9Qb
iGc5no7dvRyz+7jtl2z7VOFomFGSecvIrosr3YemYdp74Fs6LNBVsQ83dNMygMaC
NVshXaPnxGA3nGXdocGrAUsi8GG8L66rnCJAdTZx4WL+VMpRLDsJ0lqFq/vXYQEN
c4AcPU9jXDti6bW+JRh0DTT3vqC8Gl56sCd96CjC7Wrm/DpeMMyfBDTh/RyBYfqG
TpFXiSaMCKnks7PfaF7e8wi+kR3jD476ua3SjYYTPHnv2RYr/2iGtyu9AIWuCOjD
OxTl45rteqGOWdogWWlqiZWrl8g8CTg201YpPuxxugxoYgMEWgjaMtxHwtek3k3v
38docbErHO1GWjLPauHsouDoncH+WDjUrBZDcxddtYe8fbMzDZoaXXoX7lWat2zS
KnCTXC3gxU1oa2l9UaC9LFnDnxZWksbuorMmty2Fj5HmJ03RtItoWKtnMJR9g7b4
IOYWec6fLgrMxl8u6RdQ0zawnBkj4lLRMoEvWnsyNQpYtTpdg3/0jQ9abzlEUgbZ
`protect end_protected