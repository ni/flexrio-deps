`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21376 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhBNVMbsl6PTB5/ApNH6uD+D0J7Nd1ZGkjioM/q0trIs5
E/ZunsOVESFcQuX7N6g7zhp+QpEbTj8tAvEaMvDcdfe8WEDAt5sXLI4O0eXeih4p
tOFk9u6Qv7GqDWuMYMtXdoDBhYPIA7bUj1JKsJBlvoqCxwjpWKBFqKZ+NaN7bEwE
tQumPl8+12CRHA3JoOyxpz48K85sFzeQh8aOt5/3Mq0OSycFrfGTtYgPWuYHaFBU
G1qYL8gpxN8D/n/v7RCGhSFBlD7YLMl73ic7BylF0TLYk7Qr9GFf7znezLZEEb4b
PzuTjr5xnpQqc1/obfRZm+ewBJMvNCL9nqhefQYXcQtgHZNgWENDLzaeRF5lS1ka
mdgm1kqBHwSvb9IiL4W982Q8QNZf9qQ3h5yDaxPcDbsH5mfWCvgx+8WmrZR6OaQM
Hf1ZVzZLlbUZO7OI9dbtnZLZ30mlGnuYIg/p6PInSMYd//pWPcyHLcjBqdyDHnHD
ZqPIqxNGgRmAC0W1XhlEeE1Q1afv0AsI8nbMS+64PkPRI2lDmIqxUqncOmmQEsA0
HIkZnOzuNKRtg6wWf0jJ9/+4CCm/jQpMFYdwRbEC4oVfgYeyfsuHQuYhgoTOW7L5
J9RfquF/porkb8PzwxCwAK8aDO9F0+aPalnfjx+BjQqfLhOnjdQZBe7IAkbV1c+3
MSFi0Huzc/AmEWLFuF/0BCxERKlFeFWBhhS66s7bovWV9J/8ASGsTCmD3TZ7HtOO
fBczjbXN8t7bQEjJZQnhHSGpAcbCsajpnugHgwk381rlc/2ebwJ3HEia7uchvG9k
9MBxLB9TepG1m7S4tPbMdpEXJLNUH3HU5+dtfLJl2P8+QKihZFP9ssJbOrh++wUN
Wzwdw3mjzP4r62m7c/aPJlqlhXcomnbPHiHZDcZyeoTI6Xa1a0AK098CsAioye7G
5I6qeikWUkG6mGl2mTObkwyKSxVAT4sNDsxPA4e+UYjohipij4/zkWpnBr+5ODLF
QeVCHrydGd8ApJm9f19V8y+UT6Qq+IGtz5VtN4G9pv/rFo56F01BfBU9clWCK4o7
zXMn48osoCR+Ch8erghDNVmLmG0cgM+DqmiTwuc4ysFMOq8CIb9UhpBHC//7LpY6
R+kx0F/JSwW/7O77w/dZ4UCmZzWL/Xb1zH3b+Dccu05jIBZxiFtnyfVjJpDRorYC
o5dKGLMWXXSTEinbEIuEGFEqMHVHZv35oNig0r+DwNZUN+3RpP7ZVR5fn0JIzppL
wv2LJHdzl3AXriGnaVi+jqMU0Ds3kEEHLhG27QCHEpndkr3kOmtBiAkiuyr1/iZV
yU2bjnwBEIIil0XCvtnrcX9MaMwjsB3kVqHy1Cbe7ktnDOixGojzXuT7dL2y1fBV
plOSEmCl8b9/m35OPOmmFLks/i01OD+QuRHW1JbUp2WXgscThIGLagzU5ZgAKE6y
1zlM0l6rpCVZ8N9vFKZH4ANFsn3yfq01/TrwrCGwlKgC6AOsO730ReUT8JHUQVZd
iEMAwFBreruu7LYPARMtsfDJDt3rZymIjJlOJUVrN7ixuvO3NKuy1zDDO7wxoXsE
u05xz0VR4kCMBA4yb20UAOs6ahKLsgjV1EaU5v1qozIzUSvw5KH/Yzb/k63Sij9Q
Ki1pvfuMvQroMMr+ZjTRuFeLoDZH3RW8akmcIYTXsM0c3SRdP+tcRrXGI4GvBb8s
9YI2QKxGW5dObcios+iq60tirUvar55Ia4shvWofGWaa5RcA1HsMQpZ8vlaK5CmE
zh8MfvJhT6X4N6vOamvUZpfc+v8AEg3Q94I5IgYcz6FEMwebLMmIx+aepkfXTral
aKqWXzr8XqAfQohImUwdd+MD+VcqKZaqOjibxEXFAgnZc7DpjHbr+Z3iSBlrORsh
tjLk9MP0vmTfM0svhRZ1S8G7Zi8z49wSpVVHJFVHett0cEy2p6VgS/MmNoJFG6ye
g8RMmJzfWqKoV+xShSwJJPyanO367tfrwsRUbdpcG2h0Pkg/+3Cp5ClpOxp1wkT0
/hrier5bfL4TxV2688wTr+SRl/8KxcUjug0YUNejzEz8yEObGSckzw7EAIcQ42ih
S9Kx9l1XwCLk5jgKljWnTH/BdzrsuCOFRRmVYJRwnIo+DuVerAlZzc9Yl1bfZqCu
KBXGa/8du/mEIpQqjuJUBN/hkL4pUJ1M+IvnK0P/GbNOBf77vEcQfpgAnJAsKKoV
Rx36U0muzKvZVD1u80H0lA9M9uIes4TuZWC2WYcpj+IOMEQpKLuVe2YQwVSzpceR
bDaw65HSUH9KJjl3vlB8d4UL9dZdxDz28cLXhzpq7D8LwoQGoPHw1/SSR0/mgA+C
p1SjgXrSrxnkL6gYN8+lHKReIM8kCJkz+XkeChCZY2cCAEJb/j1NYCUC8zoDPN3p
xKD00NYhkoBGGKJm++kuzwVc7HJdWHZiz80mjIioOAqaLyY78aYXD9mTY2zbqnl+
RaufsDJcV/O/D7676kL337bwrigKW2nNxrvVxbGfbPdYfU2I6t21zsT/bUZP91tC
6ZYzDsQF3HCHoqWjhZ8as49RKVafFm3ffGKq2dE4ZgD631GINWCGKRLV6xEDDOqz
GCjUusuQOj9BfPJoGvBXBOzP9uWXw2wQietzwliKqmGb1wXVipx0uKONDgrIq1aE
GeYMD0Lo+2QoB1KYR0XuBt+oMD6ZRm1ltHlkWvYI1jyn9wP36d5JnO78LbEzn/E3
/RqJkDAwxld756WlLLbjD7Hx1nx5EpLvC2q3Vc/OSP2hZnkngPeJD2L75zZb9+9X
hbu/YWTx/S1Wtg0tWW+FhnVSWmMQOXPxKgN1dYu2iLquO2JgtTxgi845CLdKaR5O
47K1ysVjXBKlygmI0gFxiVqzR7OsqUFlN9Zy/QMtyMVyFRrc4ORkQZm38LsQPUR0
+q5WFmx0yKsdew85OL2LrHb367GewUiwCcXEGzHsWQZwQxbKIYjRbMBCVv5iJiUB
2fkEMsDfRbkI+QfDm1lkk02chkAjxrVlRQHXSjsORmv1pj6S4DX02nMAs8RID3qB
165NElQKW4AewedcoT2IU/tZaTMIdDffVso7DIcbjzGgYqp/vWqkB9Ztrr/Ok4ES
FePforZKngsWpAZCCUMQJMVxGPsAFsETKuRkP83llXYlcKBU26ysmwoYpc//4St6
CENgezczYE708tNTBHadpZ1lrjBqNCUp2hS7dqVwXbpRIjHew/i9TkzwnquBHnNU
+YAHZ9FnQjJMi0kIaMWHjw/oD+BJJHyB/UvjAqcoAQ0SyusARfozD6yukdnPIOaI
+omkyfk+t/WxVgQZhi6J/ahPhTI2drT2YhzYzQOYuJYb022eBUDlfl+0F4JQkwLO
A5hPKoGDb6OOIECoMqA5hoMe+hSjYuI+wGlInzWSBf+DPKnad3tENcmvYNQujll6
9sFQLkKA4SUTnNi7f7vs+u2aHUDNNNTyXkT2vJgDDgx7p+KFocUEQBiosK9ekR2d
jjOZyAjjkiVatLAuvRCu7VE+Szxvq2MklL7v6PUwRMT1+cKiSOampZ/Y2oHctO8y
fRSeIlbAUMAoljMg8rSxU9xM6/Xr0fbKBAGSQZ7lbBP8S2L9RheCFMhLw6jsJ4Y5
2lEJ92TzxJANrduFBOElVCmmPXIFFbNc4rN5n48UW4Qlz1DNbeT65Lq8bdTdnsVc
5Y1TInwU2OaVe8+vtLrUPr0AHdj2by0CvNosBrLXM9fam2Z/lRsUxyaOoJqkBSnR
Vv1qpgPfJmzdgBLmh1yOQy/kHOBYPa7y1QNRB155+n6lmUrhT9U+wpwtgAquYq4g
0FLYPuvHmCn2gE90L7oJXv2ySEIH//sZwUwMntZCw/8Mi1RjTpmDWIX808GwkWv2
A2IsBbqFFmqq0n33OALCBH3Ci/nzWBioC7ZAPyw5X7q+NI8UCwCFCI6Q8iNkRFTH
vS5gC4uf929GnJGaf2EaFKYt7P2/6gOh8zGxbsemzv9kGGMXq9nKlOuA+Z6oDY8H
Ih9CZ7M+hZQyGsm/YGuQAYg4xh0H1m6ggF2IUtERNbqKxvFrI2ndJhtyOZcAK21z
jBnNht4xXHwRuENPmp3sRgBWo3zB9lrIWvR0HcSrRCjJ/ufq5qnzcI1L9cdoIcia
eOpPQ5udp84yzyBvkMiADdLOOz79E+PS0PDKZ1t/AJsRURTi9S3lPFpHgpHVjsu7
F5ILitIkr2CxidtL+Lc4820KCMnXu5EdKSVN24tWCcwA765r+L5jRDLDICLBUX4J
MWYXPgkVGIJlKnh6ZJ18kxr/HcxKMBw6rctM+Czwdckc9sN/4loAk7ecj4BgE3ev
lXqIsYPU7rjF4kxWos1Qwngyc9ZOSAA0qMW74bitITj2u6U7EJUItNqJxwID/plM
49eXQCX5CoIJFU8bFjd0YdpC7/Xt/lGXPmAqfb8wdVNKO8OI1ew9tP6o222SAPex
Rp2CcRcLUyRBqGXe5wDIOG/BqhEVRdZkY6AsLXr8B4wpP1IKfooin39IX4W024GF
8Lk+aAZlTa5l09e8yuhmzdbuP6AB6tbnzmY6OZc2Ff8ZVc+z48PFQqWyrTXV3fNE
m6mu7iO8TDIQI7V2RHSDEcIj8Ybho/o6BRSk2lqID51tZ7/PCtEZLhMtbt+feWMi
wKWlMZi6WWqZI5eUpuiByW7lMun/y2m/RUe4jSkxNw3NtQ/LZclADS+z2RSHTJWJ
md6hjlmDtDA+U30KGjpKYj7VCIzbAsq2q+g+FgA8yVUxwfyoHi5RMvKb+0hf20Qs
U61Oldhj5kwFx/KJA/5cYyKZXV0i4xO8GtvMhGhgJjpKhhY4P4xFqOuuRyO5BJmB
FsN/2YLCjhWSUyGTtnH3F+lknzZxlGbCH5fQXbwo03bAlTjGzLGrWQuVzh/z+0Jx
AkBPeCecGVe6Scv/Qs9PSTnLDjS65rxd3NIxOawx8y79VKIykwYBwlCnAopFgXW7
UYI2/2idYE+1CG/Yax3Yu+aMf9u5azGRJJfMcV19ASlz7iZBXLTW7kOjxptWxcZB
NXo5HHEXrH/JNrclTsHfoaIJZaNfdTTENqDSwSA5dU2sg19oSYTmL6vyUPkdOx57
GXjATIxfwZ4i69MAAg+HQhBDkLJdXjaEpCaf+nxqBrBCwkoF/QRPNpS9G/kKnInE
JOaEnFGSg5cWYiUF912UaicjHMWeFdCcv9JdjNVpzeJEgzcmFo8DzfR2AjY7E4ab
dSfyYJ/M+lPYj/eHEU05jIrAZKeSAKGg2+xUKXr8a0cFa8iX1U8Ub5zrbU7XCP+w
Ags7r0RqtHTiH7180IMktC7jEnc1VsiDffyD7npoO2f6OYx++mwRT8oUhwr4BUYs
kIHzNTs1IFw7Gf+RcZSBcpHo0uvdIz9Cxp5wWzs713wF/YsGuQ7b4C+g5dXUVUej
jnXbyDByz1yywcy5xHZ12ur+xZEVYfHDz2l59+QBCBc0J1HHNULfVwDClIF39j5r
1/Ml/dC81GEjYtmpeNoDHHlW4arOgP0BBqaKY/UrbdreyrB5J9Yjh8VW7+pfTsQf
82jtYYWhHHWR93/GcUwHucRuuuHZi71XSGi7XOBoCP/wtYQusWeE7qZ94NvEBGSr
WcH881WlD74ROklXg0X8zrpGSHCtBwrRUMw9+Ar8NzICgFjb0xL+/MZKmZj1wQ9h
+/C9PfX5lcnWqs1PRzEM7s8FqoeYhUjAX4l0Gh1tsaqtQTUUwr7vz/WSqn+ejdaA
jrU5w8GV3zJaXcrJem33WoMABvRVOknauBh7VuL7wphI9UXxp7xhHb3dDMtBEMZU
BrGVIFrGyyMPTQo/vPVseyOzMfoVJaicGlYEa+lfQ5TpJAADXcOrEkALp7/UlspN
IgKbcFyIxN6JgvEL2SEGXXTCaPfmG3GXmP/ylw6pH1w4lVVNm7J9RDBq8eFXPrVD
yVNz+1zSaF9UE6SMN3gkl5PNRGquaAhJeJ97QO3CPrWq/nXpP+218w3yDGBmcEQs
izkmtsP0IJ+3JTq/H/mkDZXEWhfc40OH3PrGHyOgJXgW61BF+9RRsHxZn47RaARk
Q/rVLnj06Mo2TjOtt0ZTKgYPgjFFY8lFUtQn2ECYPIZ+QRZZITUZrDnySOyOMTOU
v4Q1LLdIo0KENr49IwFsIf0Ydrnk9ioYfCSXkAshnf/RPvEWReuxbDKTiryZZ8D8
yg+ZDV6OqfDOgUZOqL+BpRW6CvrHuCFUeF4L7MLGdHFptZ32Z4wpxHWWTfS9JeEC
+WFUH+zFSnJIrHiXRuXAf4gl3HrcHl1NiIaJzhAYGEp1qS1Ym9NM91JG8K3Qz2M8
w0Zq2S76v4V553ATjb8PCz/SCMtt5pvmvPu2g5jdgZocslnAl0P9qJ/BxSTck6br
VmZwuaUFGFi3dj9LcCH05zZJ3pjGC2vdr+0Aeb3ts4TqPGtgQaTCCGxVFrN17AEZ
F45J3g47Db8ug9KkfMvvxNkI4V7iDUNcXhFYTAcPdMTnKDjNjJDUjX4/g26gpWo4
EVeerv+aclGvJ+MnBewg6FnDYOr/I68rB/S71vYhm+wKobTPL84VfjFy8ixFh7Rx
yuWmonC7VgF8tNxjrxYdLkSlVH+xIckdrLlMV7AYpDdRe3e1eU0nR+6fk695PzM0
x8kcRvvIarx5zENUPY9o1af6hlTdXJ/jvKtL5VGzlC47rJ+tK36k9ipN2jg2/lEJ
0Ep0bEZ2yGX8v6SfWgldjKEirpP5ghpSwavuq4DRQHMGVDHKiy2MK9eUchH6XOOz
koNWFEOo1/hbriv5XIEtxLxfcx0MytHIhyauEqrGCpNh/NOhFIoTYSPpjCWyqj69
bLODagBNIndpUgdvGzuoqx1F6S48g4VePvnLYkdFTv9fso7hg9LURut5YbisPb4k
YWgh9Iue0dHhi3DjGYTcSiVkZjla/VXUce7zihyavtt0WK2qSvnRDT3tf+2Qq+rI
Wolr5IdLcQCioSYgYw/h1xV7BXZYr+1HKzNucXaHAoVcVRgR1CZl0v4K0znR3EEA
CnB7zv9rletgnkLRAVbrGjb7ofiCD3HnuDYZFzz4d9MDvcH9vd0/P94js3dMK8aA
nmp8CuQKHCj29LSGc861KZ8ancoSQkrxWA4qeQuloLq1Mn6oHcTXVpX78KL1VPCy
giD36Uyk2+1uOOxOgLQnELYqOIvT9z2zSSw9Wd3Y2vqFe4ttWsWPXqdufwtaWTE9
sGubcOV08wX9WGeq2bUWBNhQsu1HO6sE4iHR3Bbyj9+PQ4VdZ3Am6OfN9ZVC/YEG
NapOIV9VsB4QdhPSxYU8OwoAhNeBUiQ0Bmmm56Ud9IhvI2Fh+8yUVzwc3l/r0TPQ
5VX61PfWIAZ0yM+zgRL8/2I8PRHTNfhstlWXTdNTQpWmyfvNIqUfD4Q7qMhV6GUU
zeu2prShgVhQzjUo1IbKnPvug9pG8aIqoxBYpbl8AVv4Gy5cdP3dWrDXosIlvz4n
rqvy3rcJAXCu9uuB5kwqqtEC9JC20xWsgYbvEKhwaRsNW4LfuuPXFtEG3meveo78
6eCSMo/GOTUjNAwDUs5EJ6h1UfrqOLRbM9soX2FrIlT59IDPuRuy2pd+5j0Pr6/r
2STpVa9AQjRaDaIVZ/mKtOZJaqRCqa9wUHT4CrbeeRxr+k5UKQPUjssh7PHxDzWt
R/22wWMbcbR+IpgbEMhzfJGLX5C1HS/5JWuMFitW7B/gOGziGYZvPkNnsTCLfjVu
kOWmnylNxxE2iPycCf0objOwPD1ffP04Yr50PaMHFkgEUJxQnYoHTZFK836qcyYK
mutYc7nFlFgIsufzZda8arpXMOMKL6cEWKEgAbkWzITUwHuv9Rxf7NY54qYGeWm7
y39bYu1pYUC4bDVm8+aeG5npoRbFbBsJ/04bD/QaJkKdVJN5zjfhFb3fy7BQFof3
gWFdrpXI69SSoDbqEDaGN/g3qofyoTQoQsbT30QGv1sUaW8wCWbC05fxBqr1j3Lj
LhJgL55gUNTsrxb1kduHQcb5wHiPQvhrjkfFPMJXL07r6Fks/emU1n0fuQOHbmJM
9PUV88optwCYmww1QJMaoYdmnfQAc+1rII/Tzezk0O5JiYWMUlTYHsivS5LsQNIl
kyyCLMRjY5mhduHKOIcaEZoWQFNziA7BFPTjyvVYMfAtfWELqnwqYIxObbdIC7Kq
za+cH0HMArjhErk6rKkAMScKBIielR1mgN/lCN/MH1+urWW9rV1ms1rx7DqZOzKY
0aq9L1Br4MieF71DhiIJPQbtb3+CggONJAIvquyNqoFq3KbhJfO453G+gLuLqfMB
aPN2lSDuhk8uwxd8TeI0Tvuaat4+doluCd1GgH03vaMwX0aVpm9trthxFZ3c+v3a
Ac6A9aQQLa98ffWKdGiVH+82WVqU5u0gO+GPvIuLT/9fKC6spotFrtBC0sv2ilVm
Nc2OMbS4anp04TQuTJ+LRH3CquBqL4rNdhtg2an+WwJU604pWOFaHduQeHP2G4vO
ZLxQHm2ymKVa+VwzX/2FkzohlaR4u01RdS/NVV4tdUrJsQo97o6th+A2HNE4AMd2
ohOd/zd7ii3gmm4cA7FjNtDpum3HaVNzpmt0C/C3J7g5bfu8DehJw1Z/+mJWaSmN
gMGpuuUPchUTt5tTO512aniduT4zyZItI2/5zqCgScKpOwsvADRNYcYkEQ9gwYTX
SfynAfDA8ka/RMEAGNS38TRAK+g52OTtVcF8fuSbAtuBc21G30Eug/uOl+Xcwcpj
yWLsuY9Fqg3EHP24mP2LtdX32919ViLEkoLKS1gfNsOysIP53fZdCvsB42RrvuOQ
jN10Z12OIU9jPARj8jexb8x7UysDZbQSthi2mw//vg6Q3IZoiTrVO9IWJbBUx8NC
tezUNLxAAOTa/nXL9lqeG/zKJyUQb0XKxR2envIEEVSqNGvtr2H6eJPT9kLQvHK6
87wynRLvguXTkbVB9VOUVcdm4h1xc7eWJE39kYekAKY+JdgX87YDnppC9vYGxPGQ
eXYviUkYNoo0xSsMGtctjySGe0mbzmLwuLIsyFzm6kky+bzs+IC4agDiqrwI+pKr
m4hACXGFP7W4l8D3KAafnHi0QRX5KCbiTyF02xuWwxyEp91Y6cIC/zkBuWeIwXi3
rzp5lvGUsChjKygSOxIVH3RpLMvrDZWu5UsxfbyJnlTd7Y/s1zmQ3ZMotUkGbtKe
f/SDJbsGK9MAyv68GlhyAD0J0fI6EV335H+q14phmPpkp67FT8/PGHCGeyEpbO/0
Eaa6kRSEQ8FdUCtS3Tw2gOgDnTQ/eBtlqA3tyV3R7UfkxAOsRBcQn69G7VWJ3BDc
9SyqYKTTV30BhpKwSouB15CYX214yZOUVE2nFRxoOSTFxH6N0UQZ0rV3oMg0p8Gx
kbo0wjQOBtRqjr/RCCnG4vrWsexGPvFno7Bg+EdXTYJ996ZH20JdcSUnXfkL/gzx
hb2GvkCHq9yjeaUFrs5sLTcF6bFR8W5Ujw2aFZzS12qdOpQrsveW2kZKLXXwy8Io
d5vdKnHGK2WGm6zTZgBYIMARAtSAj/XknFRv0uzS/BGsMPdDPJA7KSRxckQ7BkET
ktemw9J9DkxoX1suh4lAyoT+Z+d/k34Ueq3xkPfMa8yGv8YdGQsoGDl+PDfk/onX
rwBfEgwzU+KpOeyNjpj/4+zw5aHyTigNX6SlWcSQEggb2kRTPomL673YyOCFLOxY
PLTF2c3jwJcJZaiNYBvXhYuILbZOZxLlJL903MDSpUhMiuvj/bOfcQUZAXLQVjhc
ffhhUlcsgSR3WOEcE+/ABdrGr3ZnPprFzmxzbN4DtHGtUwlQb037dMVhsLW/q/aj
co4T1bgeeACWXf+xC8ALj9h313Lm+mHkn87AzMRLjlkgbomzoWH7h2ONd+UPFOrg
wTCv3uGBpL92ZPvcPqscKYcUVnMBgQUfj6ApzvLLKLIJxvf5Mn6N0yNolOMGVIVc
3f3N99wQRbjTKahTsGrM1I1N0tP7tMVwqnlU+pu05rmdbknWPfgNtyGT+vnF3wC+
9U7/KiQv1hS+/8mwFuYPZKRMx2NBSqppeQLhuHm7Xy7P9+e+DiO/de6b2sGPQ8yS
Mw+8zNn5LK7TALatWdkLoeBAaofu+MrDWV0OoINfVkoDP7UG7d/czafq3v5l0kVg
Siq3xS3wlGcoJNHQ3Wp9d3iKvzQaSUUORTFWPgjROo3EvUZadS/fimTZjvgMHotg
cyJ3zAgdksZPt8essptTvpxTT5eikqVxuhv7izyNSKEaY24ygGLXpnpPLXe6GE28
qcOQ72kMqnpjtlv2flSi7TWvg6khtlS5arWVrVgvLO6aIACS4BGssGbNcJRDZ6xe
ZvgFJXUoOvo0X27pjHQdz456SP20Mc9ojfjTEt8UwylUItyKxl4dNX21wyDiQ4rU
Pg3nxQwCjzFXfvaQMzfty8q2EvlMk6rcFKXKqDlHosIl+omL6IS1/Pbx2tSOaLO/
1tuxkKR1x/sn72ROEjaGFruhDQzjm5NOYe9Rk2Y6Q/bpyQ2NEtSEQp4VEdhMcdWz
Orda4E7EsEYu38o2wGlXzGZUkF/6skFHt06MqNEjrlzguImNSB9KpwjPu9qjcKgc
hsTdDAwlbDf6La3UfwKl5ZkDynGVsskT/s61p0h74JU3pU4N6GNR4NosEEdV8BCb
VppiBwW32m+EHKDYwags9ZEILkcp7XZM/yvKwZPtVpt2cEEHrCM8iScXPy5qqdhL
gyAFsTWX7NLiFA+mT+zUrj/m/Zbd1YElHXQrKqIQBohuaBhOmF6sRDWRzYAY0sLq
T3hfwU127pqOO1O+aL7FZcSxYR7VhKaE0IFwCxJDog2kqSj9wJ5RU4QueytjXdJl
k0MoIe0amtDD0caPVRPIxDmk4VTYYyq9KrQVWoWdUp/qO9jORkMOfaGWpp+CNlTC
MZrfe8r/IaUDnmvEQXLFhHNC0kMVCL+frXx+qwHnEG2xfvv6CeSsFRZNX+KTknUm
eIdZ2cY8Wbi5lldEJ9ShVdO3Su5fDFBWoOpfGK0fJf4QbHJF063AsCm4OmUV/J5a
4Edgxp/+kVR+WFzoFwGW2AsNB7arnBrAwVMNWjBfvpzRYsym5ONJpDALrBc7Ih+S
T/e2lSBhlvc6/nl7gM2fITcnxJVxuI9hdnW+Q5RMj+LUfLBc30d+kT3pJjyjhmK5
sPxEuiVUYj8FuzcKpupDs7yAqLMuaJUfBrq613WO1O4RA59Qe+HVWyI3r8qkU/Um
twkZzCdIjNFCgwULcAjohFMqCmdQMzM37lhr7dAk3LQJVw94FBmcL4wYVhEizhre
boAvm2lDkyDC2SXrLvK56De7wZDJ9nAsEUyppKVnVvi80XerALQ+RERYAMt9l7LG
1mHutoIQuM37N5VAXTIx0x9dyE4x6E/31sYBVYIgnsx/65o7gisButcovUPBhouE
V7gNJMCVbieNFz5Gv8WUiI/HyfIraJVHEq8Ny9Y6PzVxfO51EW9EB3tafBG9guF5
HjHPJMArZmFF8z3dxv43/g6jhuA9JCgzTWSme3CptsOWNLZ2URvzjsQicG3vYaHt
ao/slDmO+CTlP5Hm7iXavxqzhimCNs0+UmmfEGtzavhAxVycbb2yx9pPu4L1WuEh
Ozf8x9ZgQzptI0Eq0N6Ugr7NOAk1CGgA6Aza7dfWdojBvo56wj8RrI4xCiWbe1/I
TqsPzdp+DZdHkBPTDGWcHn3kMWqYWZ5m5sh8fDIrml/YtwcfWEszfy54LpfUH7ZY
7CVwXaB9TzNqihVSxdVOOdHiUZBtr2PVeohgDYwZGNmyaJJ1LSlsuho1AxaXTVmL
uJQjwRc4YQ4kMjsriwBA72vvHA3yYgxUFqgwMgxhffKJVnpQGGktljWwISrihie7
jXL5CgIk3ed/YlQf03DRjU9MzsvCzK8XyiOWX6rjcvw5JTgMV9uzoRk4mZf7FSUW
8W09v2L12meRBjNq0y9jYigDfTZ/lg798rEsujkyJl6mgilyCd/JvIaczqF2BqLm
SvLhcrGlpcz5PVOLVbNKlr5SKq6/hpP+XDrxS38IqMKfsDiUgBggKa66GNqwh/UC
yhbVsJzA4/1KEugF11lC5W9VewV2avLUkJ/QaRbDmJa1/bKbqNNVThJneB36LJR7
M0pt7xMjPhyryyZw0litu2GquSSQKZs//iNUdS2OpsITJhUdJnMacJm6Vgc6HXMo
Fv+Q999uBTPZobASlboIH3SnwNLAgQXsZDIkPs80DRvryxCl34+UiyQmIkv+1PSz
XogrbIxQmzOH0h9xk9J6EIyXIJn4WXi7rBMfOw+btn6ng/K4z9eC43L96mP37Tis
d+iBMPK5++iAuQ0ohcIHFSuIBLZOoewuK/GdGWsHgHw5JzKgpGYKBiSqKpBRf2QN
I0L5hGVXFLiT7a/UtA7ySnBH28M08tf9XtRMRQRoNP0iRol84etS746XJZagv0Tm
aDBsYTBTzoCzXWXvjny1oPITUJvW52NdUcE2QhauAVaQsyfGeLLKrXLUZpTVCgRj
m4J9J1N8jZqayMUXo2DN4TJJIqQyVfdEGYpCWX9FJTxP2/tQ6EAMdLjGjMrXQj05
U+aWR9wsbDLRFfoGC3Oc0DmoUG5hafGoIPy9LSEgREmZds2bPGk79GTrhF4ZJMHC
4716D6/1w3BtMIh7iqGbFczAiQpo17bh8qT8AH9c4y5e/NhEk3WIzOmFKfK8KRGg
ZCRtG/69AE+y08kG8BCyGFihCQTGIDXOEmlFbCOG8oBD2fDUQiqFeFYToQ/4SDv2
IA3NmT4d27UAQ/u5aQdTAsZxuHyVl4nr8ZDpAn1v93X+lhZfRybFT4w6i9H+DCO0
idT4/mrEisXfGMY422qArcVUwufprvpJsp4LAXSAKGLUN7Di3kbeuPJITcVHGnhy
uKjq12yKiS83teh6qeig+mQDxJ1ZTmIzsR8tWNHfdQ8LtHW9wMibcUVHEL5oMAJn
SDnWgUgTdF0tCSdf7oHNk8tmmOpMm1IcLJOBzSUKVkquFHm4H5o9evGkoKlVoC66
/mOmdkh9HFf/3KYxSyFPAwKgYwETEpS4xyRMqWPoLHeC1QKY0CZTlVIuVFSBgJ2k
llBvCoog7lz7igdWxnfV0TmJyFKi4mDgPJhSJqE7kCT3UIc84p/2YtGM21EgjZEK
UgAKXeanIMRIHAdTlMrIawF7rjxavHctzvOKttEXrqVFekRivilLFyu3VubS8zvE
iEgVaftXPC/+O28mwwuOwxOPLsLYHnoKsC0NCIkXevX2XFkr8CQZvaKG20j0ErI4
oQSMMWW/Ne3iqdsaLgXOsZNK3I4TwXSSGikbvtdrZbwXbh0gS9q2sOLQLDHCFlQQ
uBmpzy23i4eBLGkzAwyeKNYBSUsNFV0BTcG9kROSYT252BWA7nMmXuMTL/mIaxmq
yEEbk5O0YRIAWHgG5H9pBoJ/E3nUaAzKlKItxvMgywJR3dmq35PB/hru6JHSHkRW
fIaK3LTn283fpxwW96Hu3usLYt+ROyZTo/Vra8khK0wIGzSSR6s2VBOR/1qfA0gO
rMnlR6ZgoXsmaSCQzQUXpzYcpStYLOYOUBQs078YLrEZzkp6qdZNba0sMHwsDRQQ
9NfxXMBTnAaIi/zbXDkDLrjiJGtPXkFz1hbpScCAw2M2BXiVZ5bAxV2mpbcMzfx4
B8fxLOSyeYTPLUdB0Q/3xDQJIuqkGUO/8FTJRRCvCPhVb0Dbym27ht9XSMrXBe99
7k/FEyyN4hi60k21WrtVV+3d9+b5htMtBqqXuvf5LCMkkhu8s9euzSUcMcxGkI/7
gTwsqs5zHYmLLBXriFviqKwxw2ezoU2HIUov3Hb9DF1snM61qyVpeKAJqcx9ZiwK
15wtwsV2r2brzpLAqI/xcDCkOkpFZKAifA3M7dtVZux6rn7iACb3UDhauGmqJR36
wNRf7aWLXWBfWn/ra7mSvBKhHLEa5IFxfLINOjikK6CnNzOX9nE09GjpOwVbUKiN
n9mqGxKd6VhpK9kO05vplcriJ+eJhu+eoC4alANPk0jQwKKCQ9XwBWJcMtSHpOhs
dcRF3l4cY4tLPW0yo1v52BRlK1biKtngYMkOY28rGK26+dBoJNr3yosy7WZXXlwL
k4AxiP1nj6n3mK7e8Nltd0gyV0HpLUaHzrXSncP3N8bL45jyXfSfsUgd+lDykjS2
B5LEWAElegPDtSIuawQ/gHhILtE9Sibd+1Ex5liweCD6oi0dAFr/w0MNWT8EVg40
7qov1M6bMaRJZEoKubq76caGWf0negLyTgsmxka4en50R9CnLA41aCQy3VWj1848
8i1nRJqwaA/IUVh0g1d0NrXyjDu6iAVQ5pwEh9J1D/vzOOKW+Z7qpAlsEgf7qLii
T2wnass6jGP6PsYsZlymKRwiabd69hF+V0gj3SBmsOmBxc7EcljMCEP2BHJkqKC/
vztGsNPpcrwaZqN9QZ5hUrHCcwbrYHkshQN3efoq7ppjj48KBrg6wYMyOeFW45EK
ShOwvhaIdQt1pmSL3kXm/uMosoYBi7KEve5GrNGDFm7isoz1t8wHVpfGqZtdPpkf
WhNQEcKtsv8w1tIF6vKm6Yi6QjYMzEwyh4YZR8DZYgm+BTY4OQIyyLOphPeWoTZL
dqaUI+vbHneGSu4P5ifagbZGCEo25MN+NKrT0KxBLEWO6GSo1KNSkiXytXAIdEY/
a3GoplzwggByfjcRWzABzuoeMVHoMrkQcsVMaFnGmI8kmLE5vlPJKWqw0AFAHSQk
E4Qw8zpcYsEeH0sREoQuq7QbILsYadd//TZm1DtN7/9YCgr3e90WXu6Pk8knc+Q0
VNMRVt5oghlzUym+bMGCnP/vtALUIBTV2OCTpDNMxHHTbG4Nr83mnaspzEtNYWT9
pxqw0qQhhniWLs4/cCMLOqOe8DbYZksk1hZNqqgEfA4SOo54KQ7yNXJW7pbco+7u
692KgN8/clWbdv60hb69w7EkjA5FyMKCOovBz04gJB3Ad7R4fXZTNmu36r860z5+
NkPDk9epEUp2IYO2xfPXsmSo5PlLqVi38JrZh5FnXV/yrhisX6Avgr7GKmw+WKVr
0acPET7l/IUOgsDvCaORuH6Adt0wOlgwbVbdlLrW6pbUVU6TVVx1aT22VOPes7Bw
Xfqs8liDUVpQqTfCXqp/iTlR2KqoGqOA/pSDciZBToLTBkoLj7Zpfm8UkGoycAvp
hXoFypYMAt71C1m54diQhAPI0dW0X7EcKz3gUBOuSU646Pkex0+kf6RK35SRp90o
1Nlgb18XJk17i5LHtZXVXtbyBU860UJuxulCSxRADFvwvsBs+VxPcjXcrF+6T0d+
D3fhH7Uyu2x7JvW1wNFoYS/VmeQmOOB8+L7jjGuOo1jgnga8+lRKig6MnyaaKUT0
OXP4hFwlyA0ProY4bw1RIIxJ9X/jtqoBg4JPChfrvAAhDOF+fzvYHIjNwGINxAQa
sdFFUPN/83iXX6QjMGyd2Y/Z/TvZIdfNSo+CKBEvR6EY5fTO9xXqbUqFHeotqxan
03wN8TXJUP8760DjsASbvCOuez4B4+KWb7MWzAk0diyWfgyZn9J/MHus1sv2nuxV
Zl/rAmWNrgMfXexhCZ9Xcbrnc8d27abHZZDydCiJWKuohtkPSRFCdc4ivMa0meMv
CsRE3W/FnfuL07yxUrwtlHP7cZ+uxYKqzMZPToYXIKSVq/FhiCFVRveWE9/7oLJH
q2uJQpAv1bxfftZRSEFr3+JQEkM4UismWMAHXVJ9JXPvXpS1VvnS6r5o16u+bR1D
ZmX5MC2pY8BU5+nql47sX7IrJdF6otG1clIJIeWuA2bqNpSs1lJFHTCq8vw3d7+o
j4NuhIlSk9CrgZ9pi6h9pX43Ph9cFpJcV9XLr1ol5sdescZ47aKpsDw+lpWYQeuZ
jlNjdjsyAxtXUjpjcpK78yfnSsa78kRc8qmWHGuWJPf6npF3ppb6dJtsWUn6AmY2
H2z0aQMUy/gNf1hAtXsWZ2QW31XxGIWWsC4zYV1wKEY70JGjqS07GIdRoP2Hcnaz
vJiy913E5lKaTIRXDYiWB9ZTh8Oje6feIcCSVfi/ixCLMIDCT/41jPz+DDHbpftJ
r7P6mun0esIdJ8nM4xIaGBCqnRjCQl0heR+EAC0Dh9LA0zqOav69uA5PeHqTippJ
M/8dUaeQcEL0U3+kWemZzMXNQWxc1qbmtsb6Cp9U9v1InlkXTfaNMJx2MGJ/sNFu
f3tKgcd3CqWjorSIxO1GP85RHbsPqYJg9ALN/dCtIXsxgwEVuRljDeOsGx+MHvQK
AtsxxR+RGn6wkUfBsN/9P9TCRG6q+kgfW0mhs1eELpzQtHy+PiNq+P5lOTL6ITix
PT9ccMIISOIgJDP3KtCYuprBzShGJ/FmnaS03LsRd+J74LqaXbGgBy8KKCNFdPjI
rz0ICQJD3crzfDzA0wbPsSzhnQeSH4zcrYMyq8/2gWBMsyy6ITBSj9wYkxbqRcQl
CrahTj0/zql+R5z8tVMmwvY7cNC7QNAyCoRKzVz+V5znmOQHuYJz855hn17i4NHO
h2mfJmbC+pSKdqOD/yEtVNPSh8y5ddgAdafUAFSA8SkY1hC9jeqbeIp/JfgO/NPr
SAcPxKiDIEYatpfnHIt/NRzK2UKw30252fyYitPb92hR3Ss8WmoSdZw5rDeZs/PI
4YwpP2oQrtyaocoEUN6HfGEIie1AqSGBAst32WBYIB+HBdrAcVCR5yuAD7v06G6K
Ct+7k24+YlFKZSdj+yuxXYmi00GVDJ6EoCntV6kOdrRXvuioBSDTiEDJ1uDmWhQ/
juCYH6Pw14ClXbb+z59sGB01hDbF+WVOMYjoxboi8zCcar1XPf8bYIyGtsy3FJlU
udsZVikFM95PuU+FTYNezadon8N/hv8ExPgPKOpYlptSUaqxcD5dHzhol+siqDMi
GermIlM7rCS6W14TspMUIf8JAlEGbIYJ7aop3fwXoKzVATb7icKgBlH1ARRkB5MQ
d8pm/BCADoZonfKNRvyJmzaWTkOkK2iylbqKrOY0EeLeh3FZX9uia1NxgsCBXwY6
ty0bLpHJXbLKufH8QQbU6lVcUlwFdw4t5o4qbQh7Zuv7aHAJtGqQpuZOI6df/jLG
bELDq+r+fvB7I2epOGnZcdFbyZLlWsCslTmduvTQ1cEHMFKD0HWsbjd5eO+E192v
q6Y6APkCcN4XayZvxoN7wGHuc8VsCJExLIbXxgzOkt8ytOeKYJi8zDRP4htJfRct
qJi1hektL9UWvy9xl0BkgVjqdsSsUn2N+dNOcWYW0Ql90NlEE5hFJ5W96AdjX9Ij
v7GQpIaVN9EnNglln0K3yUnie/j736lldDbPLdtyMf5VBvtIlUQTP0Z1dmnQqn4d
292AQXknwbz+Q6m/jQxFPmB9bvv+YhdA2DtkAiDeDmG10tDeVTgBtMmb2ktRwP6h
1+YCM56jPlRbX6p5VWIt244ZALtRq1ORa3/u563IXTVsgQm4KElmSDMK8/twjDyZ
SQMBsgJuBHC1Fonn/B2xOs4Ynk3lF/QeMZB0OTsm3rCHN/e8c0VKZs66CukOGxeg
q9ziXnjKrDO23gUZccdVnQbJYy1jrwgvU+yHVDDOUEEaZf5TUiHKmMjZvazeUjpf
9LWm716d0uATA2OGxjJEFZI01YFL/r2U6wtpOyX1haksZ9Jm32DtwLUUesXS6Qfv
5+cU8OpfFZoNCOY227P/Lhp7rzrsLIpF5rVpCmyzQP+Ra91Li0KqYzFybg6DqKNM
xMUmnKvgkFHvqpe8/MqQZxect80YKAQx2BERfILw+TNg4Cb9KSYO333YIoxXM70H
ld6x3pSAFzPBmppj5QWxR5fVHBdQ2Ykm7UH5WaKUrDuVAnNuvXN3XekFfjkm8N4V
hWYOGg0TwVE4XgiYOlTbSzSSSdUSyE5Zl4nUveSSVtR2clhPtK6MiOstlZe4ADN7
m/+/P4uZTIXY8ZukfQ3QR0FQnygtf0/axJHZcyH1R33a8EnuvU4MotgYiOswfwr1
LjWGuIU0VXGtkNOI06Kw7XLdVUWPqntfTlkO34NsXBzVloDBtc7TRfuCc/rwBdcz
roSq5RNpF8vH1PbAKQ5ZjUUnPuNQetIUFfR7xZncWwRJz1yyL7Ri2NdaOoxpTPmI
icf65WHqGFEaokFLzRQQcUl5hFWFjXVO85khaLXp4lwyyEuMOJIL4a0vNdb9Et20
MR+MWn51pYk5XTG7CLr9mZybRFLYvPc5cy/lzR2iGolpTMtAVGn/lUK1b1dr8SSg
ea8zBJ+USqWYMcB9njrxSUlBk98YPiAfLCPNLnfyeWji+PI0WKKb769xTv5YQsxP
s4lU4xZhwtiDu//J+A/r4e3HKvRkWVfOycwAFwm+cur+uK0A1ocE94ceEejqZ5is
vejEnOg10Yl/flgt4J3seAG9AbMA4ydr/u1dMiFC7hjrZpE2Z/HgoVFwaY9av86c
Dxnbxi1pWZ5cIKPklITRcQegBUgfJQ1OQWHxHMXlndN2izauzyJ1rNaXOsriRx2P
h8nXbxopWupGp5Q3WuFtdUxt3Ag6JOs5OQ5yj+KcnZfnNNtKy2RLq79+i1x6k6fg
8rvzY7RhOCBcgvhXjIrhldp2/PnO7Vz+MmGZq3T860TWM+1BXhzzINVdCvQZC0va
WNMDZiKO/z7chemXvKS3BF0SUEGl64XRxzsm/p+NXMyDUh/dmqSloGuah0mVnTwA
afhAx05cj90YChHGuWUSYNMkqVwB7WE4JBfjEuU4Ugmo822VyYRe0DXazoSVfiF5
93GRs9/3TSHRJDIAHytirZ6yVgE6/Iv2iWLUobPTXQoNPu0B4+gkCDOaiXm3EwdF
nzHOMllx7+g6y40N4w10yoU0jMr2n/lJQEn1U/+TZqmrDOIx/Rr9+NjoUwQGARts
O5ZTUQro7e7x946kDlK8X2u4PoeTR2DtZC8SIXhHBQEwZi+bV2p5HX1x5Ihch33s
OFOeB/rNlTNnSa4hmFgOTjlP2P1xACsHSsc8gBmRVR1fwYRy5iRDE+HLcNpVJVGS
iLUUT5/C9Njvb+L4/Iyl4AkajGMLlWBm7Wf1iO6qVJnoCFMOgzfKdpOZa6roq7QY
7n35C1svyiqCQ8GC55j4UWrti+c9OJuOkElqy77iJ36iyv+nwjSkXwmxionnsl7+
KZhXeDldyOP/zsR2NeK35e+HIEQ+lVspJDrIYod4Er+oMK9XQY4USXhDe74rQ3WN
Vlmb8dR7U4+bHr3h7qs3l5xoVLPE9MdA0P31SYiduPhcYQXcBF26HHrzd3VWmGtY
dHxLjFyctwJ+GGfs35S/9zwAXHS752f1HbZWI+ThfHsozMrKqMI+YZo8g711lVjC
20Nyb66qLuelo3DEKqowD4AeaEwAeySeah7wmb2r6aTBYRIl7lalCvLRCQ57OuLh
nIVLigO3j9HcLxt0DlHy0RuSOPM0cQBic71H8BpgwAqneCVjxj9BEpvcM4hgH0Fd
8+yzSlS0YoOeQmlkc0gLu7WykgB6EkHaa7PahI+ngTmG84zgqES/6Aqkpas/bQEI
cIdc4BT9KDzswK/Dhg8G2oHX0mC1dSis2TLG9fzhTIgdJRPAR6xtzIqFFbLTtxYt
f0/Jyy7qC3BCWiic4URWyUOS8/mXGbrREBAC3FE82JJVJZezPKPa9GrGE0NSVp7+
c+LA0IqVrlfr5FPQLKcmtjcZ51+0UNgjouRsAnDBRWBmLd3z5p7Vg3yphaWR/YQn
NZ128T1HoExrHRojlWWbLUm405AE6RcxDtYkSsc9tCsndzBEYm6x/mi0JEnnGisd
dje1Ov42kBnZQDfdWehr4vR7vMCj9RdpejW3/OX8lAZruwxdu6pJC1l8Cg0uCoiO
w+HP3zA2hKcpHvJxzKX346Kg4lYJLjXwwUUQgBjqvSiUNqgS8cOvM40mloP52Ua0
sZg47E5sWmDryWWdjsl5rg4jLVrjwZkLLVWfEX5CKDb5f9+Z4DmkETOluHI7l0h0
K/jdmBujAHyzBBfH3u8i9AIKLwiDx0vIgtmrKywG0zMkYKeY2AlJyX4a4vFvJ+Gb
1gg58tzSATC3rQhDpSBmUO/9grRKpO1Gy12FlQYWuCUVE+pID6h4rzX6EJgx90xt
u7cfv8xUnf2x+v6J2H50rDicofZWg3emiWNEkvO9tX5R85+M5P//Nluc8b/TA+g9
anUM8WJt9YjWK17KpZTtwD6hHyFbfgRjl6l6H6wetzcySuhauDHmrE4MaL+IEpN+
o1DRO7LWLGWqKHdPutl4c3iyZPC5DHM/jeOI5yX5r7JWdrk7dHib4Jho2dXX+crP
xbt1QUd438hAovKfW5uOaiCA8dvT5HJYFfE7Mzd5WcZkQQCQeb5X4HwpGprlFji+
eCygHJKUTBBu4ntPno1w9UtrpSK3mKG1M6jNg31afup0S8jgKKKH9raemf/kLv1z
ing4YfXg7hwC3Y82TTRg+oEE4O48luJH2gzbmodbKju16dDOh7JoKENI/Bf19Y0d
Sn97ig5Femr4xdx9VqxVzD8eEGaYvHdUauI70cZzzwmtB/+/97IieK+NNPthEeqX
nNTuiK4YU0JTBj5NhYFrE8PGvxpmmTQHQb5q8/XR0bD8sVp2AZDCw5j+VR+PK35L
BFnArlDU+LxqOitWhTQHeJLiSOS0EW2IzGmgRJxKj9LiYrhB+e6Zek+84nhBZti3
Bst7gq7CBUCEs+0wRt1GpAvTbA3Lxw9Crp17efuNyOyeewR5mcu8x3IrtrSjubyF
ldy+pr/yfvkOfffevMmS6/w7lvWZcG3wKYZ9tpkoXU+42X1/URzz0mQsRLoH9TO3
t9UxedYeB0UEqJpWj6cCto6AnO54zjyvrbBz/LcbMpS8IEIQG8CXkw22LcI4Niyx
/JP+UiPdyui1q8I3BFM8oGEYa80wb9jcS+bepcsFLwNb7uezGfZYe/9KLA9hlz7m
ysNI9TVuhLJVBSJP9gsOrB3HYByJYESyBo2HyTwjMHCkxHBW5toYAiUkcbvbgevC
qVUbPq8gaxR7xnXcPUspDwfehBufmJImrHMm7xRB5DU2qgfulCJH0f8NwP40iya4
f5KHlaYhvMQRVEVsDmW+L4MY/4q9LHb8Jmns7fx79GfEBQ16V7+2sIsCVadzSVVc
tQMuhlUqcOmzKltmD9dw9ZTCpHTDcnGoBXONLREZIHl4wbcoCK3OVctl88u1mec+
IhVMADJ85Io3cEh7Z8nPOTxOKmZYem1idgPGTLHo8S+1fT3iWTvlBsF7Om83S4rL
pA+Ajl4Chyhry/8+aNRpyN6jiW3FOfoBPVliZvwVfQ7vVkkpL44OxyjZk11fV/5w
+KxW2XE8AW433QWAQKWUpOYCvgAml2eWEv70Zle03HlWC3+eL66tu2604y5l8ZIv
AObmMpHW2uzoRx/Si0g6Tw1Q7cVrLqUdx9MQ/9vQ/DVwpXje+5RflTMJdpRC3PNX
8Ax/5W0umTWi5D8V9cC4ARlmYHzpZtn+i3JbwvB/Nwdz6aCf19arSNYmOFAPqrMW
Hx7J7KPbZCfagF7hNw3P8BAAU8JbeGzwXHGGcbRSP+s4R2jzYN25ZV9St76lWqsL
W5a/YeC+FWlO6cI7aK2iInWR02UbWLo6S5TiYJWV567Ictr6nGeZtGoUgilL7xkN
3EyLrbR5y7T04l6NjCyQ4BS6OmLy5Kg3MtAf1pol4cq8dIMBeu/rg137Gzul8eEQ
v4UC/HIec6HzkfBsKSG8pFCbOuwn+OToEi7l3mzOqcz/PGnE4B9V+1Jf9uq2l+PI
2QxlUh4ZMtatQ0dpuCSGW8a6AiWEvlUCViUXyVININvSSGn2J9VQC5tdz1e8R1i+
MEsjz7mGNZvnPpqyUN6qPGKheI6Wi438FRqB+dqFzX3/SC7SiaJfLmY97vEIXXzl
+KjXbxA5iWGOtaFoSd5rJBUG/cu+39QETIk1k19y5nmMO0eDPar48wu1CcMHIvCM
eY5a1soskLRTkzljpTPy8fAjR4/+3/a9aDWnMb06J03ePS+8uU80gK6ceCrrjAHB
S+F/tFSsgowtFosvQuADuWBsx1A24TADemw+v6GGfObfmnjeO0LbmJ5boSC+tWpy
CCqEigi6SAla9E1A5/WaOrWZBNBcKemPkhFhKnun98eMdJQMSt0bT+cvSjb6v/bj
qa7bkM+vy2Y9+Q/7oWH4Un80LG/c7/PUDOIX5b9pAGuawHZYEgmqDDmRzCBvlvfA
8zsqnY0o3x3q1KTyTFnJ4k2gux+wrYa8MPA3q48tsjs8Cy7gI+dadxtd9YpMAbi1
EBfleAu1ZztlA1jIqsWlt15Jjnb9Q9gL+l4DPl/3erMwOHXcP8STNlak3qTSkjEv
sXMOJB9FSJYnaAf3vsNwm5hWp8UoE53pmff5XtIn4htrY4h3SrJC5JCEmEmuNCyq
d2NnpQAWWpOrJWEDkSU3/BOqNeXsFpAOr+CeM1gHoXtAJ/+fk4lRo5l2VSnIkrjE
DPw3BQk4gJa9FvLbR/31WqUTZVmIwSyy7j4yFwb0KM5+gNCsL+SU+62L2fsnqc4d
SW8KAjwWksCccCb7AcXfbbf6Cz0dLQpu8dBLvhBh2uJaUEfjHgIrtJm/KBndpLlW
CV5ZKOEIPTbUmAMJLNLhJN/FTQc+/SPjDiusEMPf9YSt44UJ3adT0Z56hbEAhS/5
ol+hnDOtnQ0Sjo2946qG3YfdM92JG03KFc+pDoM/kVc0f2ccbHYnl1j8/geCnUjy
pZChoBBQUhiYizaX82dTqcOQgV+cjNVJOGfsIdwJc8u5HVePWe7gev2sGzE3imky
WBJDPnDkOLOWnlFkcYaJGtYVMDvmTxEpgC/wd1ZBg7gbz9n+EmCabuvHd6+seN9H
adHfXym/zD737TDvxQpgzRwYelUsja0ECV0U/Ar8cqUsEsYCXFBYixiEqnwiHNaG
xwanpsJMUgs53Vhx6xlxYGgDamVyH/zMBxiesS9EUFfWevqOwzvho/Pmjrc6Cymj
eCQidGdpVpY//jSvA6P+mT3h0knWIoNmtOFfHesXDEd+40VJAKQ2aEWUAx+54wEx
+0psloS+KibeOf2lyCRkI92hJPKBLUH/mrDuhpylK/dG82eXHSP7de7cYOMznMu7
RuSL/Qyn70dmTTHIRhtjz0G5q5CxAqMjHfEsMNSuv1s42sWnjbLLVp+kpMEmH6Hm
PPKHorDH6o5lJbJXOaN0bmMqX8b3mfKnWSEh8jz55Z+vwfwY0Ntq6Xjha4KdFRTT
oMJlLn4SlecYpnxu4m9Lw/tIUIqLhza2pa9zW2mxQ5RKgiJeorc/ZZ8obLqWgnjf
TfDdzjsU7Phyl0rkxwNP0zCPMC3QSJ8l65B07LYOT9+pNZ0zVtswMbyiz8ILMV52
+WhI5C6pRSMXiDjFsRABwOo0gLtUV/BOyDyRVQVRmiG0rO1Vesw4siI1Cek5jvKd
Xh/31uj0KxEviwaGEVufd6PZVlPuhP3FM8nn7lER4w6nKEOS2yF98jQIlDKmNWjv
5iWy+V9n/pPxyTKjQIFEIjxGRy/WUxZYYtoK1B7g4z0mQIZzDjH8N12L27EEiKSI
iU8k16uvdhRJwuhTOJonK9ndf1kSeWe7LasWLiKotLCkYZYe3EbvhPX71W/Qq+9p
VPjX5295sqtTIuARoVg0IuQNNhq/6cW+4A6I9/NNioVrIz/K61gAgTEPKZeY0mU9
nkQMCFurRAoy1CxVDevxwFukdGncb1Hts2b+O6z4nUu+X/gYzxzM9Bz0o6TL8ZXl
kOal9M4Exj33gRs8TOEE/rdsDG4Y8MUiGp3ni8pXyBMqOds5VsuChfxvaG8BCbZm
mlSKz7oIj8Re4/uNOI1ssnM5hYv2qqk1jYWbU1mLy0HjEzY6EzP3SEjOhWL92S+Q
EKCrrFI6f2JxL3Z+G/WzkZhIP50YIVsEhO401VCMKzPxZN9yUGVyhhVUU3YlZsIm
ltAP05X3QoID/74QSEvA/K1jKsv/xuIwN5TEu7ULBPcbM/JPlnlehCiiSrU5fYrp
BRsuHvAlsqzE7jRAbZBkaQcdsmmZUF21/gvU/p+KuLwAkzHRYdrDAo9FtIiVFw0w
/7Y7WKwmttxplca4ifxHU7iXFwOY/CH+N4YZL5TzLk6RycMiqxPyfg7Cz8E3Ka9T
m9IM2hq/H9FLscfbO9xhiwVtOXgRQMdoT7OS2fuo/vYlcIFnTwfmQA0CXKbwauzy
oViJ9Sr3puauDG2jBBXy/dOdsgAKtKCUyCbIK2wtHjMZR6E5lGGZNxJms+6ov2LL
QUwn4nqOrDyW0XJTboWBeUydNHvnRlweOa2Her/FeigCIkdweJOlTVy3FOeGIpvF
2qjMIx3nxACb/PiCpIU9NUXRek91NGo2V5v375CvvdMtsPMN6/uzrkuWkgrBlNQc
8r7EojAINNff683pnWXgOLhKGd+tg7SydP+Zxs/AQj4oHY5Xd5o/+wyxidtCpx0s
X2sQxBoaUWeK/TM2le3pEPmCe95mh1ivqBMrsgW3qml28VUVIPBG0UOD0zfRPp03
Br5NSvag62FH63SunjUs0tFHOtjqB4BMdMKWHKzeu+8aBiKlwL4fQDlBngoBnWnl
v+RpChNQ740fh5+nZshcFWlAZnj3cHXpnF8wwTS7G8LPKTuNzQiwgHiExnoVSBV6
GaZoFo1tSDaYXlaZ3b9vL/ySjl2xiztfqBkCQvkg23ycE9eUcgExx+OH8D4yZeF7
zo8JO4ZYZg2hbG0COgK0GjTQBIvJuICCFLQW/mPnwQQUfjM5s5SClTljfM/A9Ft2
X9TCnSJfj9rb+1txftE2cUid9fnNVE/IFsvE29KSFPmbF9rfe3uiLMS3w0f92p5v
nI3vJfNO1zC6/1vNHjVRu/fYvYuUepOmCBiRU66Zyh+zLNZOKYovoGAdWYqeR5wW
Pjm7PIhudF6foggUdgTtT0ZA2ElocuEwiuwdEbuzDvaUAhtwxpcqgeJyIYxiKyIj
pnUZgJHuQ9pG9POEi62Nt7mexEHMON2YHoHQTRqRXZLIeQ1gpy5AejF+N0oT7pDr
H1N9m0B+NsBmAsJ7pGe43jY9E0S7OensY07ND189cxiTLjWBI/73/qHqDnTcoqDJ
k2s/i6ysQGwPhwxeaE5PxXEGy9RHC9md3/O6N8E4qonTlyEqMGmTvr6Q3KBwZtTP
0dY4MGsFO5a62CsmD8Aq8sH2uj4NvhYGW8gAQ+2VJ+VKsoI2GZNYbgUTJZ5odCqF
VYqbIkqq2UnMqBw28Uz/yKF6sAxQrUbG7OGemmwNLjUz10rfomNOIFjbVXiLlcFM
rfuEslIHjylqP0HtvbrrT9fe4ekNqQMug0d9s0MaO8gi0umFJD8npgL5hN8dNP9A
bsvRfUbTKofqfdm6zgbKRtJQVZXOAQeoGXTJgGXjUIAq0TnpJPG2D65SCzrEgEPR
LrS/KAhmZxrmlIwiht2IH34tJimOkbJSzaSv9DXfmod8Xgpo0WiZPr+LpjHo8KM/
qNtFilsW9WBfeyH7bwjTC66oR1278y+LUQqkfNmwGRQAfrUc/uVn2jRkYlpibkAw
ae7UFaRpMWL/+/NiOR7t1v7ZVFO3bjo3bjYgxTtaQH86XAPf1bm9F84fwj3Px77S
t9FxDvEOpN+tAou7KVaASaZvCakz5A5blofLxMFUwAzaX2WQaXg/nW9pCpS3hJap
LILgmfnjwNh1JbIGA5lfvWAsEHclRLp9mBfGCCP1bKI+NpoSEEuxlFlAxxypTSFa
L//ey9K0LGAjPVyQClytkAO4urW/v7xfZh/t17Wv/UQ7Ff3arOAwa3/nXdDFuy1u
FqDzaZA9Vr4IijyhyLs6BMK/zvb3kAwTsXikJIc3g/8yQjdH+/bX6X6UpATcILOA
UwTqBKF3R5NfNPN5zR5+siaXDPL2ekhMZaNI3LHsAjau4JFMlkUz4jBEUe6Ds2m8
KpDv/ibY2wqHTj9/JGCrVLOLbQkqbs1DsILDUlIjJcCKE6aApzz31A+vKD+lPnfp
b3QecN9u8jEvFExGqTkDy9fe9oWmOFOMgmmbin4ocdVizMVoUd6LAcI4uC7GtHdW
m66tT0hOHLm9p6EQWIEZuXBPtKxLnnhWVxMrErmxieGrY0cUi6oTpe3zY8ycTLrt
8Fx3BSBsLJqCKNC08I2mPapA12awsvC7QTqsztqIJ+jBlWtYlXjICDuPnTjj7Ysx
Mq5P0x5NXEs7X/cYukYdReKXqljnDhOmfPeS2wUMfcB/OuDf51NbMmpGwXuEWRF7
4FeAzIIjthLXyAm1PWIAhYcQOfvXcXOmJmgzc8kjvVo2eUeQ1DgYbLN5yIlsxiQv
pez9dmvgu71GZcJ//eQtyAj7lSUR8+ttnRf1D0axrarpIcT+Zup9ICdMZtVhdXBn
hAh6XOB2KemEGng5okwrG3EVWpxt8/RVS3RiPs1J9EQRxNcYMGCC1JNAaaHxK9uc
BMk1w2YjBK1Xhi3hXAseadP0jsrSvnbXUKyN8iCTnNGqMuiCPpALzuf/cC0BK+xN
NKeNJegEz2FGnF5iIoyaKwmxzh4Q/MfkcOhtnyrkxTnxuMtLRSVz2zIxSZDK7uBl
N49KQQPRUzYKr+auRUGZKpJZ7kH0ZDu50mz9zs+6an8FR8Qwa367AGzQD/AQjlJV
nUtnmSfv++1zTMY5Sm6RkP0y0IMVJ/y7LXrQyEoQkuviSelbxCdO8p02cQ2OpKGK
uaCbKrKM9tPDahQkRWpNDPLTrBGXkqk5haGI5hkVs6XV4flaLXai0Ta7btmKwRLA
YyDJKJwqXzGARcE0pcSIhoEqDZSkU1n8w32TZiqtjxrdZcGduvDpXJGuW0RskSKC
7hx2Irjme6a0vL1tRu435NqpX2CkLtKmCHFpkOeubx584eSfQ6oRB16oB2zkg9lP
B2oHV40yCEwcPdi5Q6xq1ZivD27fV1PKLNUYYp/bhpesuJ/k8VNiDZDdPJwqDWUn
zxfhKZKBYrp1ow1uKd9Me3o8AuDbglNUmgluaTnuGLpLWB4qY6IPwSKvp9EviCYT
uKOYyOMKrA7woQbqzxuSpZAzl4nAvArSLks6W8wCQEjORKi2Px1/1Zkmg+GySd2l
z2uRc/5+r/xZHnOElVhupa/YWqgHrYEjbWXGKc1LaEqV3RQe7tSUTDV8cV19so2D
0P0Z9WAQ8uYYpRbx96yrWyDSBsZKhR+wHVjjj3j8ZGKw9Ascg1h12kY8/HajnIVM
Xwd8b7IVO+vikpArC03Ae//cvARn3u6zVysuMOjxhDJgHOnNwNRYnG/cEnrAYhcM
anwh9SzaUXgydnM+T5XmFJAAGIvbr/z/HEkRZIbspCJCQOAufesscJXfgpWoVR5e
qkV87ebqEso4sowzBAMOI3hj6A+PP/+lRf1ApR23YeeNYossLX46yIXi3d+5z7RH
jQZUYSpgpfNCyn27odQQTfcAClxPMgPPc2rmGtPvkxERY/C8iGAz/lSsj4Tve9Jl
REvPcD1Q14GU654CTI7g9AXv0LFQAuMzyDjKR+ESmK5u4axTnWRV4YgI9q8GssYe
789VvkWOAzlYQrJdmC3IKgY/FTfAhCmnzXScWFzbfzW4QrOvFRpTYFrggblQPuDE
BXY5F/IAp65BfCbfLIvimaEvnFxHNLdLkDnVUs94CLfYai9Vs/uxeRHtEyAgthhj
ypVBQfEOPQRcwue78dv4oaw4FC3bN/cyVrVPx603NsD4u1zyU2K02EclnjSUBwj5
ju7FKELWwDT8mwuYW0AoDjMUqQoFLzhgCtA2Yn9COk1pp9QuChSqmBWyMFbRzq7s
3csupmt56nrI7BJ4v+EFkJ2TGbqIS9Gp1UjD3reQ10qVoi6RDcncpZUG+OiqnbPq
YJrsbFO6haP00XicWEp3/1g9lGCRn9797EgI1JYi0RUVcv9DdguQo07Cqd69Wx7B
QaH8G19TQgXHwaFeoGhwBgLHkg2p+2CC2oxkCtQojhnwrLvm2NH6L6pNCIc+O0Ji
mWTINi4JvZKuwTH7Bd5u7gEi+NYqzJ2CKi9MiZM3WIcIkJTnDFN/N8ua0x6fyGEE
LzuPfsfBf5Vn++7rpZsBxRPRZLpxEdPjTSTH2xg5yNSCc8V+wSXRWTZp2j+JdsDF
j8X3sgw+JxgR8xM3SwPfY0hLeJR2Y8WiM2zQOH4hT6551tAwZqe4XLeE8VIkpTJr
Wq+k3koY7Yr5i5osLg0VBeugwfMJM3Xzxg9/gcnx/X6UDwe4EBNIInZhto10OlAr
n4u+XMvaF1xunjcb84TvZK7MSzH3Lbqv1t8KxyU6NYd35KDwdMP1WKL4wYLjW57l
XGov8WEQw9NU8IlXvZPZNg==
`protect end_protected