`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9776 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
Z6yALt3nnSw9nTnZfQBUNXyF3H4hW7iY/UCCECV1Z/+6EZ++KIqASFEnKLO0GYPj
ks0J3K8AiBqAWyCOvEpIHALsRnqB3KMMnkJm2+Hl8TuoVd/Hi4fv4mIszzl9r7yc
LcSkwagZqtDc0tFvRY1LbVy2i+YPB/YpFmah23vXROPjQuPmtDSihPNnZHb7rEdk
BoPzNXdsMigjj1yDN246gJIDo9lQqM6kJpJBA+a/4p3ua73uFde7pl7fv1NQMt9N
CXzqbmGOVCc28FMxkJVAXxE/MigPAVJGx26qeiTOqnXkJfiLZQQDgVBNXh2cvY7B
Adm6z+lyHUwbEFxvaQ/rS1SW0y2JfWnjdNj02b0mAC4TqeblcTaDKIi4JF4DQJBt
x/1PxbvajNCP0IBK6whRQLCXiFMR6U4JiJeN+Kugl6WBsTOk8BtrrMFku3181RHh
mwEauTqxYMmb7xk3qYkUd/Vu3y+3o2Ks4PdpquQNGv5zMIOGyM41W4nIM3FvetHD
K/mq1SefNfTP1X2O8Swo6sVrp7ip7mIT3/HWfcLSjr895F4wwn+mrrLms62M297q
hRjklocbxvRTqsbQ3Sivz6C9rh0vhxZnkEZMBEQ9RtD7xhaoDHF5Fiz5PsE4B6ef
2mP5ArZ2oneHn7YjWRhWkROIZbaKiYotCJ1F/3R5kyRU9qm8zI1DmirNY52mZfla
VTEXrujRXKE1SO7zS6A5A9b7gKnDGv3hxq36A5bub3JA0p+0gtfjnQlWQJQhPoga
NYwxM1CdmMf0XWhdAfenIVm4qYh5N4jhsY7y0y65XDEg9481ESSvjlIgylEsqz2D
Fhh7arHngXoHI8c+Zc9iSvhJga9iNdbLs4pvjjs8Xi1SiuBP37TUKcAV/mAEPWyF
lkovY7fq4QauVxs6ccyfo552AAxbvqqFCFh4s3iaTJgN6XtJIxP4myCp8Bmd0QAj
EYo+VFhc0mdxNyS7Ps2oogoF23ctXQNLKsfxzBJ8SMTdqL3gZA+OHQwanQlMHqwX
oheEPPrK4sjCRst/L1egzEyJLwPwyHPRkRda7gm8LDsBuICGvnshApiinxHF4Z/Q
/8c5hF/bVf2ZL7g8G5AxhwEPGGrMpvFHYwHupMyx/FaMzdaB9Jxn8CUyI1uFvsA0
pkqbNMFliX4J+sJP9w5EEZnUC6CtIQ3Mx763ia5ggx8vt6aWQHxaQtrG3AJTCEsC
n7z/2NFhY7TPbhhqsjg8esrhaxube9MwGEK0oQ1pChchXSN0bVZwDCNXhjUeLd+A
4D+RySBZajdIotuEDQcTslaE+E7DG5/8AfOeRTkLkuJISHhwqGxQoLRLuA99Tq+s
A7spvE/6ShmicmnHV4fgIXNGrGC8V+kb6Rcbg/vjuemk3UOf7pxJ5FwrSImT2T2n
JdiyXjsA+6fBD0pifnZKRqNB+D8ocgoUajcx85rRgPCCuY8JItfZ56/lOf+xeDRr
6wREAU08Ij2mgJTcxvWBn8SVXxqkiy8C29uxedKDwKgEZorMz1h7MITeFPZByMOB
3HaEb3yod0/JF01AyTKq1mEYVFBIIUblZFim5eQTzX7BI8FLLyjaieX8qp49vgaf
o4fjw89FocTAB4wIyOFkFroPfYwKT1ikGh9PlqOKfEThhseyzLLIYjeUVvIFHJHb
pNLbOPhRQbtC+VAZ9gh8CFK6umArGIw3FOWe86OvyEAlIIeold0C6PJ1strGBYCR
ndfoSAexbk4hXJKwHEZL/nx8GnZqQlAqmsWdqYg4/v5HvUs1bXA565lqeHdA0LYi
clMlQBnpSSMpDovMhLX+zYLMF+ZyFEcELZlnxdpHy5SFTA2kyk8EldMFDXmFtomT
/AUuksENxzkWr3AfgCWYSzJ7LBcnynLJwKinQzPkIxFjNOFDYHclAdbjAI+1ledB
ozcPSBtAI6oPHm0RTUvV5zzyjUEGfUmqzFFgPFkuzlvJGQsS9wRy3gN0KTjVAKGd
pFdv9p2lqdaXQN1mhbFZ6nLATtLjjduCWa8/HKkajZUu/20yJDA+m0yzwalMECvo
dWARjJVUKM1nspr15yENdaUeukhU8LT0ZasUPm8QG6DWlr0qeic5q0WujIJ3KFFd
h99w3xTv9RDWPb2Ed6ai7EwOcns4lFDchM4xD3bpCCd349XKC7q1ZBNA6H6/nnRz
OzGtXSBIKANcIcb+WLp2BkugoiovjgHAYXZ9RrWehzypSjyIVh0q9HyMO7OTf06k
aNQBcGDVUJ/J6nykgBneq2DN1+6L40gBuWsZWEO1yhbtZvnuhFGGpbn5EVKMWdB9
GKSi3H6VtV/jXoQFNb+6ocX/fpFieOxG7O+RYMnaDSBTioXz0JOoN+SXbJoCxprU
Y8aVqoeYtxNNBchwsdkEYT5KFfQsmZHfulsF+5FD65GGiv8R1kDNaC4GmImFMmLd
1r86mqHF2OdZMo+/EiW0UOpUmkCTmLlb8tGhPKh9ju6AyvEEX4XCOshELJzoBVWF
e8WbrIByackrcFCgpmJNPo/oTEj6PrHQoDZ9n/MJAQue1nrEejGDMVFE3sl2VTpy
7N6F1wdEbWV9dfFPQydw+gX9LhpFy4OcAn2woBJ/psf2wsGc5Jfxdv2jBMhfU472
zdB9UnwErPjASPzNoMJgtvlDKDQabgr3vANfBL+bbY4zmF3yWXSIz/WtWg+8a7dV
nXrR0RKBecKdJE2lJwqAuUvTyMiDKt32ZJtW/l2iNMKcI6Pboe6nYZh4K6c/eRPw
UTdkJIpzJHGkUUFw6PYh8aVuGIPwMgcAEvFDas+LSRpQYjrW6HK3hS8+JX57yl5/
pH/WX++329LjERYm4IRlrfyZnFzZM2tx+gkpNMXn9XEKQTQIq6kQViLTxP3sxYmf
i+IR3j/gpoh94sFZLziFpy8ii5CU7vzNfImGbjZJVut4sl3NKB750omvKx2V7pGP
3cGA9+AIhCtRfrZ/9mK8YbzYR2M0wiQnjbj/0nK99RJnINPHX5aH1UdcHSBjdMY2
jB87BXreu0VJdtqe8LTs4WIvMionfJ7R2AG26WoNAP/KR+H29a8uP9bIRkO15xVF
YAPFWmLZBw1dQkpHR8RULHD7k4QCSorK7y0e9E26bMYSdW3iJd75s6lNNE9lqy8E
vT4ftOu/crYHwEV0b2bTdsFrDxrRm4v2PlOBFXwZuTM4vMlHIF6v6ETJGS6HyL8A
281cq6nQBzhQxI38EPbU1EYdytehbkX0RMUYZtps6hIJHA3ilJ3DtM1f6TsgIYbo
A8uVK1jmzL8ZY+C01O/i0j8atoWIYQh6KAOWES1Svx+JaIFf4UcDZWMjDu6uMVhT
busjTobg1EbzC0GnRnpCyxLaCfkqoyOiYqPRORjWc/X7IeFuS283Jd/lZg5P+AJn
djnwX+D/WnAVvW96I1z4JSJpMITBIXZ8woZkQvKkkCiH03/U2BSCQbx5YBPnT6fq
pMBdHBGhwZdPXs2nE4i646rePM/b5Q8QJE8PwCPuMDxrecSmPaYYLIUKd3+ve4Ab
BhMtialKLFYI3x2ntvxLp2HWXgvKBpADs2xuip4B0vNpHGNk+vb/lKhQasryFGEQ
yNsUlEKovxaYvBtYlq+vohzBFiKrmaxfY2z8D06LJkwnqamgWI3alpD5fOsaHTKy
FTdVqDCxnMb1Z2A77CkscGMQdKWttvamUhlysEkpminhVgU/ApzAliTS8U50VKy6
ebGE2HVaDeB3d/04Lf0h6XiWhKdXtBeG4HDKSY5hb4fHor60dusQpIKcXIpXfGJC
6CSnA6APqulTpvxuAL69ZtoB7XO+wPCNWl32YXEsuft2apPptuZJ42uERVBtwWSu
PBDX7jDv5L3fi/M0RhgbvLnstGe2svuBTuQiSMA2GyrmkjYp/FLxhnLQLw3p8WJ0
PmvdwvESDRjiwita90f3ZIzdb7hu6R5o1LNwCA4N6amdKvCSVPF+/DBfmfFChiOw
PgaYnBH6xGjpFzpM2XsrnlFaffau2cefG+eehruwmoPJY+tSwcI3xLB/1NuLMNyI
Tzmr5KJrNYKJww+ZhqV+HvAeDdNLATrpRz2e+JVmEus38h6WtWmnvFC5yiLwtZ/q
Vqz3t5YLSS9/8EDTMQT4DFFhPA2bsujluUBPZFjlQOaLMFhXlBvb9Pva1Vk+nJGR
2RYIgjv7SJKH8AIqUF9xFNQoQa949qZRmY2HlI34WMMhC160ELuUu+UGOHgi/ClU
PGXysh5E/6NAyyBzsCAHJd3KTe5RMekxgbtyg1IogmHVaKBJGe8mpwkwrO0kGH6o
4IclrtWXxKlnfahAZvDo4YqhjfO5JtgyisvuA9WLANb+ZMGOyJX/0KAO3CJyAqND
LrgbAb6uglQ+WUQ5UsMKurHeGQRJLy8qiSgJhyqDMcTCzNhp0nLPOUd19I6Zzuge
O1zJl/a9jlH7OjZOrTsz+jEP31XlyCXkMwzlqcSoIg25GBblGCC9t5dPErHOY9sQ
kqfIma+M2NQXaywubxMO9cGCllZEmc+UC0Rlpt6i1rPCTn9WHvDniDYjHvK91QYM
S/Xe/KQvISKoBbxjELWSKCOc3Z3MERqVUeHIuP/q85xDagwHuvpq8+rz39+1/LLr
M0FBjm4/8HFbHqCbmuQwzIZ1T1ym4JoJ51h/i58YVZ+zy2WPW2G0dn+vSURNdrK5
/TfYMBZdHwtpBJL2duAPIN+Z2/bdzDmDMdayU875AEwobP8nF8cdfmoWIjG+l+hZ
fDmz7Qd3MqmKis78QhU+VfGhG1gvWhSdODKGyyRLrdc99Fx/nDqh4hCkXOPdvH+g
xA1fYdcWwgYYspCr6RdIfPH4aRDqnDHuSR/rGzTeziamM028qfQZ68DaxY1jpron
i0BEXddae6FQbDGt6XNVJZ3pOovB8v65pfKrckf2xQ81tmuvdPuc3Orx+SMcKbJg
2nMQ1+GpZp0fan3YPAFVbtpv7H5z6UFi61abdoJPFfzL1wzKGiIueEUPGyG127d9
yRFNSRL+iKKx6zMWUKv6up9dxyShdiedhqmEtHVmmOh56SPB1BbymNAzbaR+IAho
TIM9UvWbvJzl5Zh3bYSvswM5x4vsCy2+S2Ho1kdn/HbM3gcUeO4rpJp/anBN/R9x
YEFLSDjyvUNNMmc+QmE0O1wvE9C6XuxqKkKTEaxl5ONvLu3lWxVuoDLY7dHGYSXC
sNFy38eumPYAvPhzIIPTCZ7MuOImHtbI3UfF6ldpoaAIgGvCS90XLozLwnArKEq0
GH7jrHKoxG9CZPPuVgTY8+7qSQY2KF1DIhpEv9OY5yQun7Q+a6a5Q5p4FMQ5SfIS
O2S1wee/64VLuN/OJ/JGDgwH6jGbr0hHiPfpj7PSZIOkeSDnw2VkCQqk2XWeW2cJ
IaTspLhyg52iDOdDYhAzlYc66oQzZFpAXZMIzr8UWDyfFPrZ/rI/tWDXyGjU0boF
Yidd0uk+h/LiR5Uk58l7mq5wSJf8SSIdYmdPBrQsRarbfKtdydiO1gb4nS5GDQeL
zvRVe+2xFKWRpZqpkJswZQnifiVgNIasatEuPojhm+UbyYKnvLssl+4unl2Fu41j
q4tnmrZFNLB0PhwUV/BcKvMfDILJsOywoV2bqtVSolVxZpODaMVxsAIvSbhSuiDL
YI5zTsVo67prefrm5VY82+5tDCKtV44LIZd3357n/x1DsQMxtXP9suPkpfWP575A
6QoDm9vdSAYzRk2I0dye8ovsbCA1T4X8rhUr7IsxKFWuKkaVbtm0Ib6dYLny6rkS
mfqDQoF7oXJOCPs0v4yZeI0zZKcrwVLHteJmdkM09Ec7lAz0yY7zqZV1v3idPZQq
a+NCoqthy8AA3DjE8JKLR6r3qNtKLmkygJLgKyt0S2OmeQogdGBRzRsFiVTjMlPe
AAv7CYffwg11+5hFCT0b+J9Y2c2lqAWqvogscwgc6WIGr/T1UrCfuAYIZ11MqGG7
6xUn8LFeni7/ZCdamSWGnbrMJQq6BX4iZBe8d4p2GinLnrpu0HIR4LTIVBB1V0v5
vtcMOvTJ8W++0Xu0YOU+Lw4CP0/8rnvkd0waHUkQa6aipqQYnpriKLpCoS1ftCRp
J7N7fuX9nNF1UKtFLIpfpluLpghg9jpDcdIZTEOx7Or8axHivWq8TAK4f+IOY2vL
WPXQ4/q/JwWw6mq+JPu8G4ZThBbsgtk7aTL3Un238bjueIg09Jj6NOfxUnHiFgpa
UyP1WcF06p9Sywfgg6HV+5RjtMFn6m2gSL0VeR0N90JV9sIwW4o/VwOVxpQfJLKT
o9snUEn1zdYM1zH3ab3RM66oJL5fBthYjtfNO02l5DikNH0KQd8kcRJxwLTLeOuv
GWHXfyEapNmdw+J2ROw0yaMPC/aG7u9FRCY0GoZLWP7F7jzag+NAmM6zCZwCAst1
zCv9koDeGMb6qN70zR9b4S3rVVsbvEPzA2T70iUYNcDE4+v1IZrAoezdgE+Xw5tw
URL4yJfEm6uplgzQpjf//Yv3xz9ue+MuIb54MVglxO4NxCm1biXWQ8t+RabL4gsV
n9t/saV/xwbEJWfoJpJrJtOUmMt1WPGhmRjPtYoC5shPeCFsUXibPC4gSSocrxQo
ZcuqpYx19EfTKaAyDAzzTTvG3WCm7KNDCfHlMqE/q3dTLzcip3nQkFTGJXYxQPG9
wBoh7Ytv+7QNEgGH/y3jEZ+dl+03H+SzRFlOmsbHVqdbd2s2KBDbMXWpoHR2pAcn
PAtsU2LNQvBE17sS/qfPtZGnSgpIr7SbqYUGqIf8gBlgzg5sonIC13kWl1ydkYhi
YhEigzi0pT5k5dXc72w17J94kV8cErFWJTWOllDN+YsUyiGIghskRvY3GhyFSASB
9TUg9VJrOw74TA2SK0rS9vnC1es3DFfsF9gdj1TpyKgms79DUyrkUiCUMsA+7VKO
m3XKnCSttll7FpMuSffpEijTog9SgmAPuJGIhYx32glzR0eW3WIgYBvm6RT5zpDr
9PtR09EiTMZ/ROMMYxiTSQeS97wdVVeTXEtkArTAfkRm5BgZa2aPpxp+jagZ49nG
WEZXHRGYYfkJC/+sg0GSf3NJWuZUO88xuFC2n0PQ4z7oB1FI8OVPBIK8HCgKZdd2
RAvh61RFqqv6noEJmXd5ellcRl3hsDinlUewNhZ4EHVDGeDSwOB3KYQb2PPriRA1
enyC4nRfK09JO8hO9FOq2hxEkL8hdsaI6vNITOl5HtbDxf/QOatWqCvsHoefL6Xa
9sS0Q418VVYeH1gn1YHT/U5ATOvEIMl8PEsSS8Ftv57GNdBkQCb0NekL8AklU8bR
QRMMbW+vVrphYY/huhMsIRUy2v0KpYxYKtIfZIP8TpPN3+7B09BlIcPoGGLkqsmw
v4Zn8ZGzLNfHTXbRvwX5qgDejiDLieZQOPJbHYjmZonXoj0FNpCxuObx2UiGw1C1
zSZHRNzkEs8LIKjNTfJyFdL9WfACkhRh51KQiEApiqpHxRaAsNr7E+A3QuCI9MHB
Ykf/qKgOYcu8rnIQPdPxdrxMISqdK8RgkcS8CsxRXCLDFivbNR7vwUiU3J08alwL
bf5wgIbMXG0u8wjDzBIPgfQ4KatZJbU7gcxTOkfd4Vxut7a3BKU8BI3LQSdmLm9/
DxxWcAAcuRCCUyqmuVQ68znRFjKWZt6xW3Ajcq3W3ZL0z50TLzO7wbCcx6o9+yfu
5gz1+kuO9uCOC67K5ocWjLLzBZsdW7vZTaNTWZosoUElaME7KtCJaAGAJCKI0y0H
6lh37a1Rpg2hjNvXMDzMcSCOTZh/+gUIEEwWajihXBXSYogd+qOMjOnhUzzHxVje
gfjA1SsBxPsT1pur24FNIdlgf+3xzZDTPVF2wmhx8Uj8cXDL5uUve0P+Rp/3p0LW
Jb5Pa3SyTSU5P3r6XBrLDwUtZpNJoBcT4HkLkPFchaLiCIYzQAFUqKp69j967nAe
j73qoPkx+1848wzFwtLEpAUe6P67TV9bXYKVC/6wFHuGPecL5CbtSjbyqzHAV3t2
3qy3zyI2apgphy5FpzGF72g6mT3CFy5N6fOKyS1X/Uj84+xdGmBLRLLA4mzKZiae
uBJmcqDoYVHFrsx3BD9EatRSgVoL9eRvGOTjA2QZuPt1zQCn/kDcGq0I/9ZjOFgX
WMs4lgWa9c/qQuJPJJZohRcGyF3z/etOBFcUGXC5AA7BA9My+Y/0xH7VEM49HjW3
1HFthC+WeCafT1CWef0xlr+0SfdwjzxE4LQqVwJHHxMCJNW+o6LJvcY6kTB+6At5
NQAXonj4oqvnL3nBRukgQetOCaQymnmtAbkIaMb+1PmkgG7hlq92g/wYKpgaMISu
Z7TGa3yDL7JkGksIMm4UDdCDL7mxYaYYXYjc1CWvq14vN3U5EmdH0GltaG7vnSm3
2SWLgL+HZrPjZ8Gi2EAz4byHNBWjs0tuDJ9RPMwMZL1Q0AXlqrv7L8BSUC5pLD3v
E4X8FnasFle2RfCGPlBJMoMYEGJPze784hniv+0d6ppuz0BwycgShLg50YVLwdT1
ApvD3+QIXwxnDNpgZ7fIrj4NuHWT3Q6h7dwokz2AReEIdxwasq1KlS4xKyeHSdij
JAOKv8rqsxIarr+M45X4UkMoiuXSd6/qysSFphRIy8Ym7WEfS5eNUULJvlo6tYy9
QVBdmpFZ70aTkX2qV0ggS8PqT6XZraTQJpQjiq+Is3LyuC3NhyiH2DnS6XSgt7oZ
e8YG+Vi4hIPc5h/dMavyExsnct415pEkweqCGI9iXza5X9pI1mbnJZM1f5PyOlSF
Ue7H128dTPL31JNUh5to/pIlp/GOTzvyWo1Q1SYdANkssifewS2G0HD4i3NOUXVb
wDpOqYCP6EWrzqWJ1re8LD/U6m5a6IrVqFrRIOVBndXnEUjacM18a6BbB7b5bbs1
nGU5Fa0ynuofzycqh4noPFXwDBvRr6hfd7elQ5M+pH91VQXUW1/Gfi9XSIL05UlO
pQWTyHLu9zZQftNvxJjteY3BSnZ+rkxRnG01YOLUaHQpXvx14w6CjOWAlbvQ2EgH
LzGfVH983N1pgjwS3hialcej3JR0u8zNJH9OzOIXvogWEJy0ClNvTNsZo8hyhBjF
ZmTa+f58dHuup2BIpT92R4/7+uYaMfT9Gwd1j1cPHIPWazKR5sGAMhJuoFrlq+OS
4vfmOAiKCi9XKXIrepgTtLjzB19ap0t6oclG3L/PGzXboYqUaIKpgqnV7YIGJjvk
F07j3hfIuU1yb/XsYl2HPVSRCXsQcNuxhYAIf0us3cC/Cpep+FoRzY8FKvdZ+5ny
fBGDCwAsxVJdFIGUeSebpbTdvu4XLwSSBPrXV5k5rq1YoB+iOeqKsK8MLsso7luw
0/y0bkb9QoIW79dE3s+woFFcCVrL24fgMymRAB1VOAw+M79wyZQVuUXKNUw7I1dg
EAWZYzqpCiRSa/OzqOIN19vb7j2xzw0SspXtM4kBAtEjhOnZKGbahJcBWxoxFsCV
r1iGDIyB1TeEO5Rge7NYOWw4hhQ0YjIowMCfNG/ZAUKcTPloRrVv91xTfAbUT7do
zy/RlHGRKGsxjBuBJMDW9w2MfnCpEBvmL5RU42xWV1u7J+sSGVANmBJFtlQWwqHt
BlXpzcy3oGbM1HgWXC6kbdBZU5FsGZp/K3TPmKgJLdueg8shhilAkEvZ8jCAmrtf
DDT2Xtkdlm37I8FhzZf6iLuJwcuzS3MCVshcHmoM9aBrFEbj+peI3sWuzkZIa5XC
x0QYNUqTbUb74l5vunAHBvoOwpuo0wMjRHqT92LctvAI7U1wIVJ/VICHh+OJrGrZ
bAcQb8WtJctsUa1IBA7gGipChO0CjSDlGrd+H4BCQB/RZIgghAMQBMQP6ld3hbXT
gDm6TxvneXUn0nyTYG5k87+Ds/EGQgcmJCNTRaLpgZqpzSoktT9vTT1zu0Ny0VTo
gvBzYk7jGXekggvx6Gbkdy0zFdkT4Rz24CijXoR6thROr8Q1ioQz68CAG0QkcY+B
sGqRTpS+dZ/1O1GqcY+K6TuhclU/dZkph39bFelhJ3DyJNt6AFLiOIDCK/9I7C+l
kxueKINSCBRFCmGouar3d2AYm8yvtjd0qyDW31Kjlt7n/DNR0+UCniWCTtPV3Agx
rOl8ar+kpoJ0YzpyTebmrhggGwBIAmqKdthf50li2lzN000gYfGaQXKlZGcMYsO9
968he719HGc3ynlQ8Mzd/O5JfxF8L7LXBe+QPJ/b81GGvlQedUOEFW3BU9PNTHWZ
k69xMicNfsBk4Q/PAxw/VUyjylV8i4am6ZFyUbKM5wCtzIKl6EL/tFqcj93WecSZ
/IaEz9KvYuQzg9OK4EBk+aGEscNQavUd4NRPuQjOShzlexO98qcqwBHadKwhb6tz
MHVGK8IKpBP0MwoctpknbnOmwTl3ABE2Zaz+hFDwyD5C3+TtJ0lfep8lEYwXe/xi
hHhiuZ2cO+EETvd78OygA/mTTQyXn0H1IZEE3/lnZMNeslheSICZstkZmLB/frJn
bKNSbb21YNc9MLPwcNhKRXS98ne0sKwyAqGd6OzvskPE4EOiZGVCtZhsBOM60ENk
zFX+LifRn7u0NwNlR763FBRmImQV/kP/XbCyCSELKzpYl4l1ymuMahYyyhx5DoG+
xNZHN9bkTsadNljfHPbyFw9KfyNAoPI0iEInHwEnKJad6zEMRhSlt1n+E4G8/1zi
uopvIGgR1RlbihFfzCd9U04pCcejAr4bs+S2TKm2SUWfAS2uadEsq48Z5GL5fWhm
aIM6LhHuh/q7vbEvVoGJaJNj55l2kiWKz94u3hdBG6B+e8ON5GzMVPHAkcx7ZV8t
c9f3wvLVcewzGErePmMO+Ul5QjDXKGFyK//oBCuJMVNUWyQt34zbgiDxRazAf3Lp
9OdLG3poZVcGkoW/1mLfshnBKp3b6sdsY58Hnf+icqPaSzLa3CE0V2O9lRp+ouBd
FASNc2QBC2aXKsedGeCk81RS1PrSLR9s2937ji9H9grXN8rl5TEY/rKWYJ2LZNMd
SOZgf8v9KSfMoFqn9JUGTaspexrUIpq+4pUhq0q0J8YffhjNWdl+GhXAVp0w/QZP
syy+c497rGBq9BE+7VFA0BdoIQecOw+5F28yttuXx86OPTSj5S6UwfsHZj1d3q9j
bN13ROxSv6vY7uvAdtgZzAXAVwnQ9TsItHLYHqfiCKB0/fMrrnA1RjUgbF7jZ9UB
W6UA9eQ5n7CIxrGWLWPqjtoJgSVcNWfW7p7eC9BSK/tx92hJd9Mg5K0xcobEKUaY
Cf0trGnwRWtm9u1T/DqVKE4QUNQTeRzsKSi13Qz6EKrBjrxj0Mdszv4eCjT9jWwi
7tlNT/nELdBT8PfBrA2l1ijvev8ezPLVUh0LR+G/Wiq2aSTpkCOJdZv5n02I+Pgv
7AfCLdBdcJo45OUClR//IXlgURxI4IfSoDIyhiNYWzPulT0wqbbiEYiyNJRipZSH
9VCaxp2eYkWLNF9uH8nJcvFER8N+7EkLlvI+um8qj+ljxFv26p2jpA1WQdY1qR5v
rHsYlrUCZzkh5eW7mRq+BVtlQ9Kp7koe67b59cyBzD5oFCWsbwgApFokEQtEnPlL
PG0F0eG2U9iikmAencnjU188+/nNnh5G3EqwgubS8Qy771OYjOk1AT3viOU4DXM9
QurqR91Yv+CO8aWGs2vLO0+Gx8m5BEFVNC1/FX/LS9esN7/2q8qVvWeNw/fOPpvd
kQ+fGUB27F1Brpd5C2Gb0jysKwVEQqha1KBBG2fxJhTWKDKfhHC8oiMUHcp/OrrM
ZPRWPR15R44lXg94IQUFybVMm06d3kSjaHY4BtxbW6jnEiOWJqcoMvTmKgTGcGNa
HJ092mrM1zt3kdxSGIS5VJyBOtzaIR759MeNEg7V0bYYQUiRspofT6wxDcHyrEqz
CxIGfbyLXQsTj3M7LRxLdhVElvf8w2c8NHK0NHpmm7mZmHQ2xm/Vf+hwZZkH/eU1
SwQZX3cR7DtHyu1jw1l7dHdxxBCBWclaPk1TvpyPKzPnb3HBMgKgLkQkr6dMnr8y
FI8spkTO4i1kXbA5NS7w/16QwtosTgDkiQqwX+NiiK5Awaqv2sjLHYD0XWPLYjSO
2Yoqr0iWPEYd8EvC3JTbDpXYya9n5xiC4e22PT/uD9glJJYDmfOJRwHro4dhQR6I
1G89v8hfPxWHZGEM/STzGgzUxjH3Um2r3WBqWEhGoJCxEICqLwLRxeP5CKZ8dIkC
ZoHq9ZI0Nb1NuGmxAD4i4e7V6DVBkDi+1cJNV9HXmnIMJLH0bK21urmas1nqwp8/
j/qr6S62m36rY9P4sI8eZPBLoZMT7HKcwgGb3D+QpHZ/5TdVoLJQ4FfUnznIERQ6
IQ/yelIYrrtFBhxImGKWUpO28vfjGY8kYpfghtJIjD5tgAgig1Y/bxi6aREMq6Fr
6ate/HnO/Jx6I5R6nojR0ess19A0ZV2sTtUgUMMSHDyGdLxgsSsvQKy4MNztMoXK
Qhv5J2r5jyJqAo2BmmpZRhb5E2f8vZ6v7MkE4gKjW1BugtzJnNEjbEABOLYb/OmE
wJyPhUrOGRkvddfiCPGyeEnneoJl9spfc6DVuHc72XihRYLHv0jeS0X4dalUQTUT
Mne0jAlQ8Uf/1GZDL+E5bBIkLp5rR17J9In3+zuIdx8dnvc1wbIj/mIuhm5SoXb9
LxT+1E+J6wlVCsMjPWfU35+arFDSjF7zGlmYxwIg+LuAV6xv2FqG5Keh2veIo3PW
H5U1IeK2chkwXh2FSRq3k/EXrzOxPbDzqKEZO2HpdAnsUHNXjmxk54ank89RLctH
+Yj3qF5cAriU6z5gZnYbrhu6NDq1krDj0ixq60ZLC0AvA9N5CMtvSjHa8zSzKtpu
UsSUSlaNRWixR0HGAh/WDWQNYhKqK/w8trl+Q9C2Xpc=
`protect end_protected