`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1952 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
K21MooLiMCXVPibvGUiGAfhs8h1SsxIP3jvJioBnllwccW1ZWPtmmt7QsOiCXEGK
08gQZsHAID72CbSrLPJi7gpInDHhHApviptmpJotLnhgX4kbWt3zi6bR5V5LA4rh
On9rvWrQd8+JDOahh4GNfMd+Vz84YGHKHGupcZtaYXuHIef5nW1YTcXZ/2OtMQ4J
T2w6pQTZ1xDV1OZruLAw53ZGYUyw9FPEEWqZV3KN4kWGGVtIm/7qaenUv53nY+c1
pki4TH+MQY1EnduV1K0JhFrehZXijchw4sVwLIa5Ctx4egTu8JFJ0jOEwVmDYZ1+
Ou8fi0UA+ilCXdBo0xnmWHfsU0nmn1wq3a/yLhgYwN/xXp0Xh/x+UkzbtQy5UiDd
VvmrPTofEZi73VH8HldyKa+ysDVybncaz1sYEBG65BhsV758/R8CS9Znl8qPgsyD
eBZ1U4pxgKgde13JOxrbmKdcHF0zv3LOQaVkH6OhonDmEu1Gksqb+9ZZlbV+oGwE
7GlVqIrunlM2o/3I3lli0oUpkmR2WFzr3LtU2/Tw5nrqpIRaTa03YwISGxKO10eX
GwGbCq58DJZgr8iEIiSUCPBMOULowjjXSQfO74NZNB+RR8rpFz59hGZUXFSoeybF
JdzYDlyqckpJmhsOWdjJ3jBXxPAdhPnEwWo9dkJLeRGEJt4p2MC3XPwQ4ElFfQBz
cMxePb4EePnjnBfw6C5pDjNajEQ3kfF2QWt86DzhSDy8E0Dch7DHpY+A5F1WP4kZ
NTH2i7pf2NuZwwGGUrugUCrZ8qUWjckgUAvEEOgqKy80Bpuf2TdK55YmU4o5ezpE
Sk0UmWSym2IPlSI7Oe2KY5siS7b53tRhQ6kWJL9zXJG0INEkM6w1rIA4AGycMXaS
ugZls0ansqTJ5JPQz40bt9liyGg8yA0i6V9D8CSfpF4uY7fV+b/iBhR4SX2dSowp
lA5p2eFwuSbDZk+P5wURcsaONd2XhCihMmWMSGzF2voa3Fty+lXE31tQ29Tag+bX
adhPX/f89h/2lHQLF5X2gy4843uJqZ4/Nnw1AQ2QVOE+i4oyiG4SzhC5IOE4hA1c
GNgmGNiRwSY03v8WeIakw5t2B2r2jS08sugznyqViQmKmeKbdGIaJXvS/RzwbGVD
6is2VpHC/YmCOyqUOIeQ9Zj/nken12UtJHU150VGWWI1b40wRTyLx/L2avTxpv0h
UmbK06fHYcXOMDDE2hqBIUMW0PJmxdm4Ct1oqm+6Kab5F6y9Fkp/etAWPQqfpDVY
UYNwgAkbU1OoETOAOF355FVxiVvDzPUf2Amr3uBBOaOip9w7rOsovhaCX+TmMT1O
rIFMADD+GjtehQzPjjAqLGauOaHUquCV+SXD9MqcS0ojGKV1roD/XQMi0BwZBnQJ
dYFiB26ev7ywjeRlPKsCzGbk12pWybGefID+ZHCdiXKpn/LRVr4+845YMeKbThPn
niHOguaW+is51Gy3ef2VoptDwXOpge39eZ2y3Wq7/g6bUAfDqNaIYmXZpI0brAoy
oOuW84J5CgqTVLtjSdrneJZ/Z6tbeHyDq3xwfq3OFgVtFJW1dqRHUde+eCe9tdgI
rBoWkJ2FV6UwK32hgayG5gtpOgK+rj3rzmMchItxKNm5XkPNV/BL2SXQVuuuPXcD
x2I8rwmMLMfwqqyc3QdP9Ojii0ukeB6dGBSONu9aXQHQ90ewlqIaSAVFZLtu/ptE
ESi0X5OnZOA/oiizoItqDFeR7s5iVbtOG+IFrUUOU8nKxBSOvac1wSnzV+wJSGa7
0ORp0oCjDiERyF9CU5PdEvOBWagOpI5rhUZuCms/1MUYhlZ9IkogmYgx3uQQF/p0
3d6aWpYu7+yUq4wmZF0Kbx1J+td3PGZWBj8ERo71u0T7Mrl6IyOjILPMsWV/vAbn
sDomq1E4pr5CMuMaauC9ldnTtaYAIozppkG2CGInMWxwrha3AQ5vw+RIDxw5hl6T
5SQmP4nQlTjTsLXXKgEzw6XJvDWq96U9XZbudtPuv8Ppuqt/12hssujRNaTVPaRg
BFWptLukb+cVA8+lGMFRmxamlOzTyIaS+6+s6W72oeKJ5HONQA3KI0YHfqJ32PqI
kf9yGjYGXkhMLCGGWz1rnx7IACxlWe0hzKtmsCUs/73s/u+RetIrV2Bmq6gxvl8R
63mM3nWV18hcQmRLaDRrCWkr//7lb82HuVS2uRW5hKkzyGAqpg4rxgvx66UG7Uz2
xk4Ph8vS7PKpUvqLuerJUXpuU5QlrEl1Osb9ytJsbuj6Kwg7bKRfJkWKB6t6x9ED
J6n7KaKgyMI2wkQSzKcV2kRsFe1o7i9pvA7AzKcmeReWYEUhhy+cQZ4da/eHOnQZ
512j5MkkltQ50y3e5T9NLsUfFEPVnT1UF4TrtiZevdPbt2xJahHzUoP24FthEC4j
5UyBcaNkzs8A0RLgn2HnqtrkCo+MyyXyZsFmN+OgEPY=
`protect end_protected