`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2992 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
wcmpwSk7Xh2DEFViwcIwocn+IsGqsYMDVY/nyA0zXDqKMAGlPiXBLpMDMJP7gi4D
fpTyVlnAuqQ8Hz6T9RzaH/1lCSG7Ml61WEuaUhsB1F8u5A66s4dwoQZM5i0Q1gWZ
DtD1/ngt7+BCNBETUMq7OdG8Ejl2J+Kd95I1u8hHXeERUQ0yUjH6K7Xs70S+8nPW
xIBwZUTCGLyfpxlR/MAJDuTeumxaC0fz0iaXUSB4IC3Mg6HF/Juc5jRUus9ABIzK
g/RJp/38XsBKZjSCxFdWhDOXCn2UKn/7gVVNOrJeIi4LLGJ8YVl5QQzjw3ZFrO31
n1EdHOPnKgoBjQZa7PgZ5fiNe4ZIAF9vT91Wzav097iBiYxx0WEzb2dL8Wl3QtXK
BG156v5a8o6uhRzGBow3leil7mYyz+CdVMQyNJ7hLjjhgGeSF3OLDF0psT5RniXq
/tonvKhYcONRJPtiF3EpEynkJcxnCbjsxdp15qvXvt0qDRt4YuyngOstekrPnhvO
9B9N9Y7VZKJvxmLVHhUcuLHTMO9jww24nh6dwaluaS6R3S4Aw1BjZ52qA2tcOEDo
d5c9t4F6/XQb5ZHaBWrPZ2pCxeOM9LG00MfD+br5DOUTUiZvyzFiQMEUsxg0AHUa
2AvVgUSJIOdGyfS74KDYkHlLi1RLnwxVGQzf0nVvMQQkY3WfmtGvTrmPRjas+YGQ
Tu/rzduB6At/GWMczgcFO5O1UGUiQ6ZgsbodnNCviT329OBd/9gP9jMitz1XHc+h
7HVAJHVsjF+4jf19LGeiE5cnb3T0ChLNDhL50tq7a0pP+uv7ov+QJRNOLAZ1goqu
ZsWz0jUHn5MnX3YflCCQjZWi2Og+VWttmo4MPg6t01HGnEhEC6PK6eg7JHbLhXWs
LJQxzfE/kYhYza8skqCE+JhnqRPgNcOKzhjZ6Mqv/JHr3XTqT/IZzDGKZXx20yUJ
1VrquIC6sVM4HfsY9LzL0MXXGED/I+swN7zdMQSzOH9uUMOYlaoeqwRurJaGA7i6
ST3L1QS3Li1vit8MgpmK1t1Qq7fjqw6FjzWLmYCu4bB7qRCUBcYjPIV0ocoERPmj
0p8PIBBqk/aQphxyv8PJEKV5uQZ1lh+d8qrqTVaXUjV9jZcvF4MLklK0Qncrba4a
9zACmNqJ/j3ftvdONpztrfCBOcT5I/cm8f5kTXeUv3EVEXMmE+OU6FneIjQlcBuI
WH36rxKK07RlZcOkotEM1jvRA5b0rUaCkSji7gRY1QHrAoSPoXGOhjG+zw0upMTv
EgkTJjsKSpUZqTi5MdcFG+LGnx4YgFTWm29KdJW90anJwJ0+LGary5CuTZJdlfe3
krTYeLbyRS2f2QCzM11LVCRvieaPGHk2+uldq4gw1BBTCgEvAKRzvOfgsr0yA+WD
FLU8IRgW25GfoJuckrWWcqtI9sda24AdPZfVRKgn6s0SaMqJN09aalcEV0qijGg+
AGtTD58Diw668Z2++PbYw2IQstK9j3uDnwPPizqnUA7NZ0bj06iRs7P+kKSA+oFe
zq5IApPZOXRitZ1JL148yvAg4Xaj0bYqg887f8OzAmOU/2uLLxukpK1gViu4g48x
mjC9VePTpxf2KVAje+ophk8g0vLmxTh0MeGPsBFN3NqZgb6hwATl4Vu0oV6xL8qu
OnDniE5RqeOjxVAc9uVdh/g3qg6eNgAu1zABzVN8LDsgplybtVLM5nI13EVvlw5S
St0jFMUFuNjjHn8vvZv+JE8HsXbfkYywL9sOiAcKGMWUB6kDwydFRRfXY9SJiC0f
nwnp3rDhTyITP+EAphlNe27TFKNvUlwS++tlD3weES9yzj2Q0T9N9yahtl1KrIHj
614tnzhqRKZsHrhfBLthyIa+FxBnC3gka4ns1Ln3nAERlhsQ08OGgJSWKGtI2RZK
PNt2GFYoRZpYc1uBQm4NPIwAKEr/P0ve6uBlEmqRbQ4CZiMGgsd1FQZvejBEcxtx
2jeXyu/N0iXIZ7YA5HGUoxgOcL0ZCNYkxXzjzIZWtkCqj7wYhP+6WHP2h+zuc3xy
Flk8HNhRY/8ODeHuHdSrudrH5zIt0bZSRIjlmMS+rlVmKi31Bl1PuuYmteKyNsG2
73uvgHV0tkVeN7MN4lfXeTLUhYJBqXrIGWSEWuHGf7HzolRfp1V5nDDZH5sOC+Te
XpALQyFfHCGtrpdg6vBOuyTYujBAYrjixuH+bO0qQIdw/a0NRBOCtRrReLPYv5xM
zXMKWlkCb+VamI9OOvRp8NRWGv93wuLZlR5SaFdXgLEgptK/kwAV1VtNELFAxSAv
TdcnjebFC8z9V6mGhBMRAjGs17hjiO02OIp4SUeD80LG/ENl1PQC06RgMACi+6FC
BSIvXkIhqPB/vTCkTGRNuuBapFi843Tczt7VOUgZB1o17RuB1tVY361yr0L+Wb2I
fsDDO9000kSdHZe3j9lgI92Dr8e7GFxXgzxgKevq3Ln9FDtynRPzKfY/XwdEoD1P
avTOUaYsZiWTuuPnJ6PRWd9HMe6TwvxYur8jWHoKXsPTGsO4enboMlaQABrdebCD
I42wd14r78paPNNqVhDAP/tguSB3IgQeRcDZnJzNVKlu64BVAZ4OERs84oaTxk0/
e7lNxwRGvVcAS22D/JDQfbV13wf+vjm8UhPs+jzSPCEQydw6tkQgVXTXx8mHSh8H
jHheUQ81Opr6u6lFdJYt0YW1m5zkBtsl8L6SJgbSA3674JvqOiqQK6q7D+pPtwkI
pVLoPp92t+gFNCb6bfSvU2dW0jSeTgmFcMQwZPMY44B3cbJSqYmNVu6o8SiwziFe
qa+WIDlTrIKGIEJ0GwgOdCYqYiKU1avvUSXin2tibQMoLabb5YAc2nAoEN5KFedv
ERKmpeJfUYSj+ITrJU4S3R/sSCTaAEK9Hs9QFw/3X76nnENXXRWyU1KeyvLqnBMs
Ot7YAn64gJXReFKqLUH6QnNehxcI4WqBpFDcok50IfUDL3ZCAkwX5ExT8jRwzWsb
rlpCyDyCaA6RzO4jqOFD+G5xhEXTXbEtGCAeceO13F+YAHR9QVpqsb+xeLlgyePT
q7A+zDrVeCIz4tm4r5qcWryuWIDADMR8K/f6rEWdv0WH+Awi0qIKFWLEYctBswju
XauRlW11b5Rm6pnPbRbcT+gue52/qoGbvOclfLbI4QK8/CO9R2YfGEBFUG7hbkbe
6RuJgu622ENyT6ouelUV6etIsWQHPJMtTSitCHrhcMYHw34BrIVxTnGCfDuIyVso
9224S57Nmkeh7kOPZBoV3YbD+2xwL0vITpANTtYln/Yfx0eHqM2YJiGnXspZVU4R
MtFlrKanwleCWQx36H4eoEiibBtUFoW4cwS9zJRy8ufSlwxij08Glq4BgDrjZjwQ
/+4elArRywOfk6ABVBlm5QLSFWg7/pnbEaJUkw5ReRjRtu208IlvDgTtMay4JK45
Chi3IYTMYRyiyTJ1KuVCk/e2xjtpT6iv1uK+UOWxZeRDmQ4XKgAio1cLxaQNqeD3
Ps0lgFf+l6SoSrvOnBc9FkPEedhU+yuuGrBbOwwrrbpdQqmfyzOTpX55xN51Wy0J
Kq8ltkLdNbK0kntovnI9F+dE8HQlrbQaXhunuPEtCar/tMIeT4U+51CMA4cl2kn1
h6idHrvlf+9VoVRt3QDWNtXcIAOMF5+L/Ce1pgxBU/eW/hoTlfpOvyln2zdf9nlw
LouetGGB0BlzAungtCW54mTbWQIG00Sdgwky0Eo+Bfq5psRHhbh0UrMyXcGo6rXB
sfftM/6SnhbjowJU72eBXSMIoQ363F1nZnTpkYyTtxQlu8G9FMR3p8zdF3Lmp9Sg
bPMjU03bp47+lExxBCDubg==
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2992 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
yLhC3vSw3ZQMJzW1WqPsUfaYirrQahlztuJ1FqPEh7xaBYOpUfb34BEyiveQYiZl
Q2Il7O1ewNoiD4cZk2y7QNXPFeDUDwj12gKShm9Awum996lorzcElTih61GhiH5R
4ZbpFIYHD+Uw8xbtmpyepD2BDOsP1RHXE9z0UksjnuGjvmYJpJIxNP6UB+eSrgme
gSF8alFKGPKPII+vj4/Es0qjmQQ9tnO/Z5oJe5uzM0A10otIlzQycvkM4pDHxLNd
RW5oOuEDUKJx27J7hH21a/EpAJYqg0xTrMW5kNRO7fZ2Yx5WQzfkPSOKi3cqOGNO
p8qJ6R84X6hhXu9KO2M0xm9vnd4uFT1MvXnvLAoDZHUOilSvdzBZ/3stIP9jQSaI
dKNcTVBtkCXQgghDrxqs77hkOS+APuCdHa+QRGvyzbCoKgJP1ZDmQ/BeGo15wOTk
rsiqLGZCYr+9YHHfFJULL00yKCWFDQjpZU5gorZLN7lqZiiJ0DIBJ6tm68wS658s
M/75BRA/lESniWEmv0XJlTAiDS5ERqletIZ1JqQbhiMtYoEX0fJG3JmEXpGJ8sbm
6Nhe81IvpmlDF4JFmNz77BZ9am1q2gl6DUutShKyaRF6jGdeIfh83+BECKEngh6k
Rnz5sza7i9qo45gYfDnVWBC8KmyrNkSQ6uUEiZ+U7dmJeDTmtwkFGroIE3ghkhfn
sooxWItvClP0rt9AwaqKI4kapDs8keboz7d2D1Pftmbi8vjbGO7UYhpqwzkDwLyI
IsNH4lx553F+dR3hilurGvy473U7mpjk14T9poDQF0d4jMsigRzGsyAAQi6ccSzS
fN6cz+XCzfYcRRvk+R7xjRh2nI4YuuVVh4593K/pAIG9nXuoHV4kAn4wgSKYDWnX
WbpLIdxWGlUIo/hZALa8GxWwkPxEVXroD+FWFCwFLheHdAMwfWgxGh7c80eN7nrs
z9TSaMxzDc5Fg7uG+zwvz2zteB7Ei/z3eDErUg5nGMwxzVLmP2IB82YD9/0vvQ9r
TZB2TVXnch/kI6G9kaXOgEHsMEqBQo8NaBpiztvZxny6+Q5NshCm+5IBQEruG+la
AWWseN+DrQdu0aRmN4Sd6jf72SeuWUb4gnuuWQEipZ7WAxW4Qv1L2+uxdHiH9Yua
fS3183PSwQIqNZ+0TGbBAvojh0PcmAAe4TEYIPyRpe640Q4MYeCjXdV+ZBI+Cze4
81cFjDVriR6aJVbaB1FXt1z4I8oAISFs8kMlYCwq5h73FwyeNYDbISdSne5QIXkH
KlbROoLsIUWycRUogSOa8yJgZdeN4KQJzBhf9lVsvrdiCuu3J6HCxTeUxxuo/59g
GDgiQZXwX/8JZCpST34so2H3hxJcqM4ttDBPcJ8W/0E9sswRfTbcj5UkHyJnxNMv
rt3IQjOyrac2B28DyWTCoEdTF/J1KBxzcStuOscEt2F+kt0qIgPLWtsiwbn9chJn
xj7UYVD131/kA0JpSG2jeDcE/O5cRRHQwhKTJiuviLYzD6+A8Q7cTO8dIYdOzLti
MwzrLG61bPomVylzZBeUZy564EdGG0iqS/pGjjMdf+hKoCosluqZ/asAEusW7cHK
N+tPTizGFvdQLVtqr5HWowukXarLzcpZ+1uygk6qCKcVl75KRWNVCEyXhWERX34M
f59nu4R1JO9O2Tp9EbWDC+SGvSrDYsVkAmjBcmXLr7pRNOSTclcCD1GeWzfv5twc
RkivyZ77miqQZklx0bWFMfyBBNY07gl9MUyHXmh45kW3JrXd2iofq4Hi7DMuoSHN
N3cyKXLNNY+zcwRTdpmGvybc4QYtN6Zkk7DYo8o3cCvYslAIevBuG4cZBVMb6x9d
GHMrIHYWrCrwfdBpahtk0FQ9c58JM2iVOzMdHe1RE4c+WQR1CXV4CJpt+WZ3oPVu
/Ka9yL0sv0rEoxB4auoLQtJdqGiDlmfyzVR2qY5EwOWaGq4OblW1JSx+aAfKFXzI
8tAxf2LDZ8IPD+6oz4uj8EVu3pIDoH7V144OBf0RMtkbWgf7UZ72zHuert4SI4WK
RLROX3WBP7FLk+IBKyg6wOZ1LQxmkgzTOmTDYSPQNyvWsOGhKAYHkJydINL+x/xc
y79eELipaxNjuv0ohGK+jD9dmNeb/K5SZuxoo9xlWnBxJMquasQS9YpG4lV/fL9i
V6h/xt46a4PN412shRtvQD+n223Oddzq8uUmnTY1gVYaDJn5SLOJ3Ox4evI28aM5
asBVPEzhFqN7TTsS2Ag8lKxbi5X4mVTyubdPWmqKExGnEGyVjWBOxM3LezL1QKZB
zd9vNbmsJu1U37BP+nyinpa625f4qNxjFWcxESMLpDlor8HY8jxKAs0ncr+BWOU0
37a7UlLbZIeiJRKZZmm9AxFrjPfrX5+QADESaKeYpr94vv6NHQsgmpMRSU6uAy0w
vhwELVzZgGE4QsDRkXcCId3o6XCnEk4IWslNFS7LGeR1aTw5P0oQBnfnC4Le/gz+
okneQRMZklam6RQeEKk/m137fkoH3HbsOpzYRcOmiCsTY0V1d2/rq0pn7+itlm8t
u6e0ms1+jMvSzCwhAyjqd5rm6dcIhhhcqOjSoAgewAhtDI3yxB3w0NCpxzgd//Nb
omHoUO3KuF0N8dmilkDzQyJ6zlP/z4ViiTZo+NoU5rm51C6SNPB0XsBgEnwZt0tt
lY6Y3OehbyuLxrSFyjcqbCm4/0JEwhRghWeduIrJ73HEz15aCUUEB/n6yQyuGGyf
y6LtRohmYDvxb1ZHCSUq9hZdh/4j7Q3m+Jds26K1v/tFv5cGOgMOhBLNJLvoyOMa
0rlI17/wN0Gkb6kuDkjnnN424k32S7MN0Qda9DpdxWWtKq6aub5jk07YSTI8GKzh
SAwIVyH3SPkxSPnkwEJDw0tmMymHkOgn3MWeFhaHC2t25dgIpS/oX88wwwOcZW3N
1ll8rKtTfQ/AGfrml37uEp0GKV7X+5EG2xdyr0nuT79nv57zxTuP7hvIiX+Sc741
z3kwU5VyC+0h3cBEuha1StGi38y6mHpBQWhkibL6R3DvAxhaod5h/qvFzqJepzC4
F8JqH2FMIX9nGtZcCdEcDpXJ2oG6QmfsxUIRirtE2C51TecQkfaWxijolbnkN8P1
d9CD2MDVdxUIsn/oqvmolkL5asePF+OVQk8pZKkl5KRk2Gn18cQOgACx6BaW1TX/
UHiGDq+fTsElPSkxZXR0TE2yhjMoBK9oTo/+Qtq03/GDiOpZJsvmJfrj2e3jWXOy
ssaQs95+Exvwymj9SnlzrVaA9lYW8HJmRGc260xYkXcytvYabR4MbD8rmC2qIAkz
4rwDIpS70kJ8lU67XuAGJHz7HU4qPO9IzbOZhw+LJKYmRdWj1duHaOtlo00CZvyw
aQl2vUN09kVJDnDsoxAzzmVvBGNchIL1+hr3Vo2ZRAMEqHqcfWjNYJw/4xua0Ly6
ZfDt8XS417i87emCS9c18Ko/SLJWCs3GDHzLWIN5vO5wvzFag8DAubokBGnFzp/+
3x9e869NbBXrMa7/ujDnmXfNgrR8Ngot5lBHIwGORO/BDx+1T5hMRUcgD8kmkPUt
9eInr29KFioivMkHnxx/t/M1OUIF1HhjxLO8N6u4jycSKQ1KKOS0+xB9EKQqydD8
nlsEx6pscWAeLiauS7w0K0x8ERjATy2pFrGkL0aj2rmp7/FReZiCRmjdcTisfMUz
rVq8o58OW6m/bTkv/YhrLIAsKz4aSwbq5Vf6Cyv/9fdiqdltFdShpU/V24K7yojj
eb1I+IX0FBEUeTl+tMd9D3Pu3YXiM4QDXYEOTxejTG0zeexeCduytOedOUDeRv+R
XYlWeKp2Gl16oHzBBbXHfg==
>>>>>>> main
`protect end_protected