`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9776 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
L2bRNdr1lLBT0eERw3vGlJHdB0ZItXhoSTS/Q4ms9sN+MknGU+HyxmMzr2PEd+8s
3TUzI0yaHJRZwXsFQe0VHI2enwhJ9IWefCGy9gArtML4C00IQePcdegS4iPQSXjf
lZLE3HqB5HeYIBmVrgio6LfOQsp5mRTFLAIhdE9HVer1X/v59VFJc9A9pCKOay3z
9s9zyYnkYGL9bME4UzeYoTIxDIJyJEGTFTB9tZEcuAt+ZZBFvO50YJ7pOgyPnNU0
FQk1kZ9Nuol66hpSS20YeqmDLR5osqWarWWJD+7BpmmTkutExMxiqt3lC5pvqHkM
A0vZd8S7JQHa0fxrrKnATqdz/AHZRy6pHNYlgtkZtCgRmmTvHOH0LbP4DhYqUUBx
0qber7obcMKVmCJNFgIJRs4Me4PC3u3FL4cCPsS6MAJQ1WQEDzi7P+CzsbRJAJVY
mmJBuFGrm0Zxu9CFC+x1wiRv0i5mqGev6PcjcE4V7sYigN3bGGlcEqFL083EFmgo
sBGfyhNiHod4LL4MHwsguYNiIv+wQGuK5miNr6LsZkloLKm1rjIs7M0ue203Twt8
2s9AD2txMzzV76T8aExRyvbAsmeoyunQVSzhUzLXIUTypzzwipTM088E+Ztxcsod
ZkzHQQFiI6rjLAts9w/QSZhmfQ8beMN1sQS72Y0rK638EAMMqGAbqYJmNoqKQuQm
NZ7WcY7ItxcPRVIzB5o7SKWeut3plVSEjHp5RpANtYyTK8sxeVGbnhjWHwh22jRu
ApgGCNYwP4pJB9K+aJsDCphQcpTZ2IK5QKelmzpoahIKrkQY9y9+/BZhSRX5Dqyr
oLnP+M1ShLgTC2Dgg2o+LS4pOKHqDOLmtg1ySDxpVm/+q1UtnlGjYExmjAq5D9dD
5QcyCuTpVMjg7YMjuh6ne95DrMHcUdvfk8YC/yQYl+61zzrIjPE+VyATlcfCYgdL
PEbOtTDaOAY+j67MPHzACTWbdfowm1ojFu2Ezu64jIy3OgaIuBUqQHVNqF08j79k
cppb4B8QA4wQrpQufseghEOWsOxZJpojqQLPoXqKYdN8gN9gxAJ6pAl0n2Pz6omf
gpfygaQ767LoMPmQ5jeR4VubBrneX75sZ8i94qd6ukPvv+sHe5wVn7djHfHGL808
sEKeeGLLdzt382TYHnyqn6uIqMyIl99W2sTihtElrcSrFHGcUVDK4mWKY+En19nE
e5SYmhLni9xqOisgs9Ql6qcKiHjco5+Fd53kAxkSyUJfusS/NfbArz5PmVHfa6kc
ANz/zrfJCnqdgut4M60lY/KntcoIXRnkZszcx5Zr3TiIxOxZbxyX1ihvjbIHZgvl
zdQRmTIAlf8fsLJsgeW7F2Q/88Z8yHLOkX++vtXe6WQOhU4F4VW3QLvl006+RgFB
aVn8pDvvXVsMPvCzryTv3qJx/+bcC2C+xYJVY6lPpqZMW6SYNO0PfZRNOKlPd1Hu
1NpD2vXJi3sVLLHWZwDGG1/q9o3POagOt46bn1DYdSmaWDnJo+GkKdfffMK1KVq+
fFz2Rinsje1z7iE4CV0wU8Gvu2AAHJ6xnlB2/EeVxo//SLV0YZv3SMi+ZWaVtqKa
f3ADg6WqG9DPV+FLm6Jrq5ccY6B9JKWNV6s6zClPzVZkXC4yS1W3jMBcZYsHk23Q
bMtW4q4qePnRRDwf3oee7E03ON20BQ/X6WkO/GBzPy3FMPAS+yR9x5SJxS+5+tPR
/6Z1vxHUwgSamdNBnQVF3DGVAPXT0DhazwlWpRcwgo8Rtr9CfAGtEbgR3S/RuDHK
Px9j6t/QWfkeY1IdA05FcUFpdbxPrsKO0pakqR7Qrnaq/A1f71ChOclQe/yShzhU
Jqy3s803ltpDHMmG05JcBot7K+4fLPLrISkPZmbmQ1HeCa6NftMfryDkMhCu0EZk
3nVL31E8lQnNBVC2BVLlFTF5bPW+tXs2ffDcR3589J30cj8znthHl29LjTaESdBE
MxMX2SVD8F+3Jyzaa9r2thp3WLSW8+NQfRj9IfUIQ+vqZGM+gyQhpmQkenTYO8iY
IdAnEW6z4/BjoFyngH5HXNDO7v2kxhMJtnH5Qnd4y4e7isN0aM6QKdNQtTAF8jd9
157b5kAtlJ3jrMV1gE2zVhMQYEwf6Qxg/l4T4120+dx+0lmmlmM7r4gNY5LRU2Vw
wC+lq0BUDR2wBr14qf0FysJjRAHFK2q0aExhwvlZB2KLG5iyKl3qbrJlmslo9Glv
exf4GYVS2foj7lXfozZCR5XxGxMpTVs70hdv3h+l6IJWeyfAPrN8DBRIuy6UBgjS
v8A32mTmX814MkDDmqKasVFGMagEaUGE0poeUFWV5PS5Iq8i1eE3ksqknl346UPi
I9vD15j5RwUZrZXgFOAWSzInIgGROVFnbRsfju+5i2eTzG028PclH7mHZKjhMxTZ
UeqDoUv/TxxrHq94PHJOMMtpYWkBajY8jSYTrp4DT/7BYfJmC0MkTVmWi8vt6jVr
pwayRcy8s4x6LuMTrxJyplj1Bt+Oi7pMoED61FNoASs8KSYsktNNyvmsCjSh8jID
HxmmeYxzbeXIt6rNOimiwSH5/Dchwfp9iTm04nkPTxI0WnGWM2I8XVNu7arArift
9kwMgfbU8m5hscmJiEqD6q9kElBoW7wmqbAYZTfosmvwgIvDOpmWrbvVQNs/t4ST
e3jjAYpAoPIdUFQLBofSQG1wQoHjqNDFHRNScZG25vXLPErlAheyT9gpuKcY+Fle
7b+IYZjbYzdN2EU0l+550z6GYMU5e1An6Hm2LLDLbrPOXI28DOhFGX7wuqYWi9Uz
r0V1+YnqTHo91FMRLxDgvXYgIoiXSTXPnQbD5TL/CQYTaBp5qpxNcs3Q8ZVJ+Vtt
K4kWdI3VxYvyAkM8P+hYYgB8B0Dd6J1lsQmleUU0ViTMhDiOX75ukMbansXOJE9k
dNZS8jaeKZ3HYI/lIxduzRKrOlL+dZ6tjCFqZm+kiZhzLFjbx4YFNL9Szo/Gv5ip
sd41qRWr59ve4IY0RkvnF/9F4H5V4LTkFWM55N7A7Y+eBGZhNomcUu7b0KpI1ePt
AdXlrNkwulKiPtL0+gok5ubtpKqXveNafhCclfZWWznLgbG1qS0FMuFtP+0NeBgl
Fk8gM8QS96bKvaOuJOSxDWGAkLxMBAcNcACYmYxs2hTRCaQ3/wQqLyAwQgaQv0UL
w7a9D7DwWOGm8WOOauGVKIu94dtHAwKm+o1OwfEQ8DgPc9Cm29p0zDLFx1wiz7b9
9czmeoqDYQRpc+KAwE9qrtTKIWBpb9rRNpML/AcrzJlSGba0YdcTkKTA6uqkrbxa
NfEiXLBncURChlfqXDNNqxRkqmNLRouL26oMBq9c5nIWW9rMJ3PJ1Hf1c5Vwt4gw
37nrLP+COtxO5NC16Tby+d2EZWD+Uz6MGLkS5NVhFWWLqeJxrCLu9otynSOijQBj
p1nnHPdpsFp76WL8Rvm6u+7rUEwyd91Jvd98Z121vHOhHYOauQ9dLfWNt9Lh9w3/
DITmiHFsnX34Fg3ELlw9sviCvZy4WuMR4wdLimR+8jMKnc2aQthmi0rwpVybcs45
PM2Bxg4rhOer/fb2UQa8LkZ53PBAmYt4BBrDbhXx94MHdKfoRz+3y+6N1YUwx4Dz
8mcQ/c/fgoTTBgDmd6qTJWAhyexZGmHSo7j9pyvF5m86x0Hkp0inJKZH3f2GisRS
nasD2bkEVxMzfVZCRcAceAvmXEr5xw4KpIv5Y/bzc7LfLUasXqNxmSBlZeHoeoOk
7HhSiJ06uRrxyoDjpk1xpcLnmFykLu1LIDoo9yr5Tix1LvpGegCuUzVc0ii/MI6P
ek9SlKsch+j4KYAj+exDkfubgMWjWNfehmjBh+YYtgZGKgWlC6dTS9sYuXssR3b9
aWWpUTqU6bhEaFVHw2Ofbo+z5BLFlbqV14rrB4qampgjlBOEbhWc19vbPigCIDml
6RFbcXWlxx2jUxiBaOhGn/B13YNonTk21qg3+1bsAx1ejRN4GRylpARlyS4P96/3
vn0E4qUSw/PNYI0QrlEPa7oYSdrv5Rboc4lqRRhl6cnLnb0chqxfOs+Owur46Yng
MqdR8kg0VXp3RXwJZzG4S1xcNJlv+rDhrHfwcH4Wx0eQxINlo3X9CDCkV4Vr09tT
DdwPNcTugYF64K4W+81GqgiSqQhUDcaJfpbO4VKFm9uav50WZpEgWJ3n9SIrnIrt
2ya5g+7D4UwjgwQuwpGwvgHA/A+bvY7LKfiyYMv2Xfvqd4Dz+AfM2v11TOC4RO07
pFTbeaqYyumCdlF0iLn+dItzjl0vZN8/ENDpgnui01sSuF0c6o2jnXgrYOJ0jNhB
xJz3PSxUjg/zpp1N+L0bQB3sA10km0UgfSsEwMPRZSEJIRlxxX+jccWmUmVjvut7
WqyLWD3hq0x8sMwkS1gBcNC0HoC7zrV5qavmjXHjuUodvgZn+jMhxNxotwCb04Jp
qPqLEDk/FgIrEE7mCsocSQssdBkyMtqV/MMeXNGZxzlo2IrlDV/ruqin9yenmDx2
Zd5vX5TsYbe4YXY/bPxBIZcABHNtq3o4+IyAYx2kKggeB8TmQLwd7qs8ehKmustd
shLgO4mmDLybz96QkWp73ZpgyaJ3rxjs82+xaLNVoZJ0D5Zc2SaEaq5xhjOgzHyo
gkb4DlzGDS62xFY7Ij7yjw4PxoBa74EX1bMlXvp4J52d6GfHqHoQEnIWl037hO1i
Lqy9SbazndJcSIr6lF+JQdh9LoZXlbefeJ1jxFPuTr7NXv1WKVNkiPvqJMcEifGc
EUY3uLXdGkTpp8geRToadfKgeZmzCVlYDW49S1lsle8fMB9Eejlu06c1qWrYnN12
j/ttvQgtH8B6nDwU4YeDLqyeXzt6532RqK3My4ab9V0MW7/fIxxwquIzkuBgC27Z
nM8mM53Z6Xpb5fVk5BcAmbkSQFlH5f7lSmS6wDMpQ8K1+4npef4mgsMX0cIAzHPq
3wRfCT4LBPtbq4asDHClQFzukU/Zfh6zHX+FNNGsUBJpplbunJLK3piWzsOlh3uC
ieu9/HKnJcy94YJmKSlDzkg/8DFEu0vsHYYZlaujIQCx9dHQyo3JYiCSJiLq5LL6
iD8XO05Kz3/A4vdmgE2P/LWrooOFzTyD9pS7g5zYiJrw6XMQJdZwoxBclYyIXi7Q
pFBjbXRlkqtcU4M3Oh6zXsb9Cv/gUbb1IFTo9h5Dune6CJ2ZT9S4Mqjryz1BYg9S
o6ir7VQZv4o+KuXsRt7qJAtuLRKxyXXMQaL9OSUagL+zJeCeqJs/7SDu6QKmDm8b
mvcQB0yghPjHkp8fmDZ/Khc7BPzTCpI4LUH5LmcV5HnR1aYFoClEcFHiR41W17l2
psEteMuur3oO9PpBCQifuFU4AfIr1za+sBUyWVu+VVJKQaZ3siYAWqEBt+/t7vSR
dtHfEPy24b6C84EYydMocxqcW+Ion816uwVwlJB02KCx7Kx+BhdczAkIOQrBotR8
Qtk2s1YFvzy/JeDxNETDJ9Tlnb/zEc1w9eOVn1L9KPiTdVMx1vTC7bxyJfuHro22
Ss3Jn2g1ANWy9+hiNoXR7QKT6JoEr2/kS3MEC5yIeGfDJlmR0CnKIkPgbzK87Y08
Q20TjEZlks+QOVa45aTNsPCrBftETDXyYpnl3Nj7ty8aI+OHxvwiJvooypQNKE5V
VowArjyKOCaPsYTa0NsAu+/OywnZcTx5jygmJc7Isj/r9rj5zVD7HjLz/ELiD7pF
P7kWcAQUZjA5rD1XtiRAZExfwMK9MUtohFv52N/hKWXnJzXuUenOz5DqjHsKFNSb
m4PQWrtAzrfojpdJouoklVvh3O4fJRFMX4VpeiVtAqYS6C3o3OEs/jFhn67DXqOv
6ihckxJ9bwuovmDYdJ4Trg4040sVMU3gS7ixJ998ObQJVEVSCMbmzvgviaFF82Pl
5So15rweNWraFnmBcErM6nUZZCw2eJySq9bFB14vBmfwPs2znOwwws+PlMyp4Dne
nBgxU3GIvs99Kn/zjgbZDZfPqZtrF+kmj6mvPwDFX8hb8Lf19GBvWu/27+OGjL55
GolG5wOeh6gQKp9zQh7pno3bO8c3xPgNTolIlN5+kwtX4+OtGsdR54c7ElHKoOZM
ILcggdzczz2xajhwnMUbjXEoOLcA11/0rfdnkzlTT4Q6VkRLBirn0bNuYyCT1SK9
rISkOBInu3fXo6PO1ZqaWuipmBqBWfXbJsSaVzVXmcioY80SSVR/boF3Y/lic3fi
WKLeTcd64w+YELNwVtjUjIgsmsjqylr1kPvO9ZBIGocymZT7FGjBJ9l+YXIZmJfx
IhRk0vyJN4u4pfFx7Pgu6Zl1MOnJaqWV5lXcfcuYtc2tkXxughQK5Bt7jQJYvP4K
JqzOX5mKC6ur82QazTbN98hwmxXKO5UZee+uHiotpqo7zrgYiKj8QGYpkgCi4pJs
S0GhijRsTrhYS2ZoTFFYl6Sk8nr6m/9M8oTjFVUV5Jw9xq3cZic7J1e5/H/l4skp
dwLnN+fzkPOgDXcj9hsT472E5yHzYQ7eBv3zJKSiyWKx9rM6mJW0KiaYDMGWSU2i
UgB4+GOiUH+bCbkE54CUyvj3GyzfPrd2CxoqYXLAKDDt0+GakTnj0cfvLKQvT1+R
LMU21xnGiraXS5ZYjaU6L5XrPOpk3QP4cT1srAfQx02RP1cAwMH6/l5DJiP3ahPD
uyk8H4kA48KpW7TkQAs6p/lHUKRRxgd/U4XhChJUHHujTW269CyFc16eIejyu9gu
GPCNDUlHlKxGbwq48yOTJeJZUovYCDLIz7KnCQoZdoa17I0TtXnGFj9U6YLUrHqh
CkXD/akKYqf61qFIkMf+KjZHkrC+006nsa1cfyTu21zmJj11qfF2U0z0+knLPWPU
QyRFoT01Wh8GE4vO/Uh/MoT8EiTNUCOZokS2STHf+LiH7NzjowQYU/ydtHFRdzPR
JQjktphQbZrSV4mEIrOk8MdvyOxb87AzAoPE44ApNq3gRXYyssZesn7zkk97Hl4f
p5PaECSizNXTCwoT/zFBrCN+j/e4XG3IszhAkX7XAKc1n80lloBqMhYZWV9USfL9
LPA0qMmXlqYxaY3Bp9GPTTq2nTqUfR1gj8RIItJsxMxwlYBZKxGdaYicfoOoeXih
gRGBRXhWiR4rfRQanFXaycbiry+TFNIa7I+oX9at5a0KkjHNj+W5bzTYjRKnm+zT
rj//ERWQwzTu4l2pAuCEFnsSKfb5XDZB8oWBfHmsnLWMNRmzKF539KhsCJIDe+S9
Em6BcL3qlgbRgfeiFOqkwb4YAMt/6dxZ/sQySrb0Fm8F+lp1FgAOMVLihA4COKvh
jYqmq3IU7bj3rsbMT3ELDM5h67GViPNIdK40my3WnzkjEA0EMh+2WbgpMgLpeiEA
0uWLtWZIfKFR83tMtnMuMUv15M8hVxgWzFDWypa3cY0YlGHIoVeClmMs8vwBZ2Q4
Ud5t658jTKxYyxyuCRm+g/N1447naFmUC4i68yjGVFBrCjyu1h46ARsvVo+TjhJv
dyZCIvuupkmtAMALHNT1d+yuIu53F9NnaETNUAfd5TxkwKLELvNx20/aKfJaSm+t
JS9ksKjN0FFemCkAyBdr9ChR0jhIxEXB/d9NTdMlZaYvisa5pcsduSAPG9Aut1Bm
H+BHFjhQsMygkqQgjAECOpZvQx96R9GlxQSjmbkTU4IALpV1ZRSTO2XXleLEyLkh
yD7ta0rkImA2Ybiy8QG/eBIqcno25LUYNH7OcNrj6k05dJV6jqFYOcV5JsS+E0sp
9njrCrE+rSc9PZGspfmQBlPjLG4XzaCMTmK94qoKqztYQ83N3+6NF6wRL6+2XPwQ
qjCZP6yjnczfKTY+pLJJqCOThNdh7UpbL5mbXZE5y9gUJ8ItHZQYe+Rc+fw2m1qG
W/r01xuV37heTzGFUnTD+9H/eIjifj7gbmuyVQmMqDwu+vCYKwYnVHn4+FEA+xCX
OD15eqPhrqehoilJBHlH/QVTrMxTzmS9z6PTlxUq1X6HMuq6pRqQ+GUkK4O7wITz
hbLZFG8BXuzywtgL/3D2uGDMt771fJW9rnOklB7inJ3dyRecedGYR9yikVFpGLia
J32+1sDI2Twuq0wo4FQmQQcEWBlRIjI31cOFtS5iCBR4CSn34NBlYm8lC7n8Wexd
N7K/Noe9lSGePSTXLYb1dPQGu2BNP6mn8PFxGd/e+u+dzKXdJM/j7z1/MG7dhFmz
sbAo8mQfzlqRvCG67eWF+c5tJJUH++NzxsPVAYm3tdlM1bj9B+FL5or0Pny7HEGw
GWiCyAAIR84HI3XJIbviVjEld4ERvmwssBpi13lmma7oapNovNikqXMbKn8x9BNk
q2/gTPni2q8j0murGWS45dpT7Bb/G326jgtndGFVWXQC0vPhXATzO7pnLh+16Bro
b3m4kP0Mr1BBR4ClDwzfNpCxPoh7c9Pv1hoGIokAYHld0T8z6qE1o0Qbl6OdRO/2
WgZlkWgyyH0eLUh+KRMhyldvRf6ZMVc+1vLeLTsMLIyOjrlk5YQbTlcTb+1MKtIo
zx1iip5mLapwxnSnZ2OnuPjQ0ead+kzIcHD4OVYYpWu08zxodmSMJD8Y5vhai9Pc
mosgns10NMh4Nvuyg0hr/sq975WkKGvwfZ575E6I8gBuFMUmanMrqnpz0FMAehi9
Qg6JLnC5ZMlfb1WPc08ZGZrk8dlJgXmnDLXOPtFrrldD8K/MmLkpj21RmVAKAO5g
qbFHpLJXgReajKbzslg0rv8QARhDDiOlZW3ua+8y8hBHNkNeiHoZij0+n7gFHSGu
aKfcUY0TpsGF2g7BsewPNv5xNn+8UxpqY4FHGYn9R3eo8+XPQkQ53KFTB0BEmgJi
7cBRgAelvMyBD9p3WX+ZY5huQ22QmPpWe9QgU2l0SmFkTZkNpLK3Tcs/gWY52Dox
hDTips7Ge1NXQtSwmrRgOScu4hooDIYljN7VhRhj93XeJhn2kNFKVy3h/irVOHVB
3nCBDwVQ1clft66CH0S3wFGERr9SL+s6FQ8D/Th5bh+jD2K/f1H6T8Zd5yIVZOpQ
7R7Cy6F0Z/IsNtOBQUYwlo4XYSZdyVwXSlV9P8XNQn5+6oh/5wzGB6iYqD2xCYcn
Mcj2Vm2kBhVorwz3n3xegu/AlQ3fp+9jxsXyRdEJMIsw/XpRkPUQdQICVm3KHL1h
6gm3IkOuvTIZXZFDMG9js0kehjY2oPohZjA15XeRLonXEZ3Onqo34XSIAaaykw9O
1Rh+KV166z1RPGOhIu/Qg3a4xO4ZAoRDaXNafU+FvSGendVXfr1ChNcCHcCa3WIq
lE3XcOmPwUWCuvrcAAtBWXzjMHl7nfHD3CWovLu/lT4LH5exV8ZI5qBOpLKrHFEo
se+8bjQcIaz2PIJxmed18XaoA3yblHcU17A+dUgEI2v3Sw2zS5luDdsQr+TsO9mE
v+V/qbhSL4feevcUOytjtq7ZaDcDsloBsB4mCOZQiiVYb/QUORAYNv1GRGgU+r3a
OLT0M2ysL0K9NLjI0Z7z5VV9SzsUuoOLQOSsHhgpSd+NMDwedRLBuTyLuvu9fQPt
f5T6Bc+5MkyEDr03j51uBPay3BScaitXoWcToLFQzMQVPsYcsbCPINcW5ZgcyD5a
St/ETpYm0UKpvFakfGVXhswAwT2Fq6hO1VRfeWFUHYF0yL3FsIXl1Gpa8uJGWU6C
DN0Rrim5wx+mFn4SrWNNgODIlq8L9uJbB+xvPrr6lkRpUt7N5qauq1JHKP2psWdm
/CnScrfGx51hvBRlhoyoLldOfOnmrx/olAnRlSmEQ9UEwQOobJeT98Li84pAgylj
0JulyQnAmd3BQgx9+RnZqt0JFwdtSj6vh62xqc5h637mWWhms66x71GxqyFCYmIG
eQFE1+1dcMEcauRk4niOFFChe+o/g9cbOZKa57iN/Oq+78iPgYyyPh1GKTrHGp+N
2oAN7k5waAcNycYws99C2oSJaJBNB2oUL7vmfj4wvt3PXK6Nhzs860BsZF20dvuJ
rORSukJ+j6TMwXA3dun5jUI63OJT/1qVK6+DxVp19/fvm8eyedvPTiBqgv6lozmH
pZKDftjMiZdf2i7e/UMglB2+3xm2R4FldGsUzRphyW3gFPRa4cRuhqlN1CnG+DMP
nkjSLxspzZWKyMn7LDvtjuxZrCe60+I9YVAu9bqxxrRjMeUm6I+X8wfW1k7wdAP/
d6AOLHpToL/+53dILC502tqOrefU0mvfwe1GZlVNPd/AQyoyAzmobydhaGrt1QCK
+O3IKRQleO6JKwd/k42GAoNghC1xyVi7m5/5PHcw4+XGZE9NrYmyhp1W5uqwV2Fp
Uo4AdjjJHl8P6ysyQXNRu6TXqMWGyNC6cJ40EjNkduQ1/VWeO3w8wBY4+Q+Zf6R7
P+Y+2iDO5u//gYpaRefKNlUjCgJBL8XTaEpqI+r77N8GuxutY3mjYhZmfAJGx1LK
TjGrb0M/GJI2DRbrfE1px78iLmbhAqLLD3YOXzz9H0St6ykFQKVCIpt7XAIHxx5e
N0oEHkWuZLsHO3lmtyuK/9nXVQAtVJg7Vb9FwtU3CTzCemX7Dr9lquZsCY0pop9n
72pkJ4DPBORaSkn2sQLfWZhfZCqHXNev2i0fSNRPjf+TeuWk+MaCYKTTcf+pB+Gp
apW8q3F252h/2fAYr5VHyRHiLP7OzmPCBCwmhvnWywlaw4vhkbyW5FcBhdPIO3Wc
bN/Pen0RIss1/CQstykO5qV8HN8mo00oNv5FoQmK6zzGJ1qG3lySj5HNvXVhYsPV
QDyleCEXWPTQGMLypFsoyeEDR4rsLknR8qEKxFQrZtu4dbAvnrjP3YtygUs1aPqB
/Qe9HbeD9SgL2rGEQEH9fZXjJHwyNhwVdVPpo4SYE/HThUgmlRVHJWjckWdZqA96
bnWsi/RW7Ig5MqTQCHdobdVesIOMiEuxWwXTRBxPpykbiXeWaPium6/DLBQGF9sH
04QHG7kSgZrRBQS7gy3Gsc1lEAYVZqfTmUgYS4alKIrbnpzkzuMiosfhlpr/IB4O
FXGsttqyDgE3dlSxY+UQOGF3MMNPwBkx7D+pQyvSddAU9sNcejhdSV/DS3dlqleh
xHKvcA4kduMVRXyc5bJceeZGdGdAhr3AOy62V0aXLi9LmpWkScKBr9qgqq7oo8/M
HVbI7Ry29hbrgrBae2mlT1GiiuIP16plmU3olzGJVZE9tUezUbDYSJfCtPhN+oQZ
cAxlT4V3auBZQzbf50h4NblIHSK7D8ZMdbmWnrins9Q9xh4e6wIf+r9n2ASbWZbG
H9iT2u1TzCldNtVLn6m5qn/Wl2thi79QhHVvxtF3PNSStjAJJz+yx9Xv7CT5AO41
8ksieOnfcCUEoLYe/qC7+QmP8VounmQIZ/2hjGrNsQxixh7xlgQYsO++KMdstdBH
V84/8Swu+tS5xXarDPCNzlgxe5q45GhirDskkE/7i4lgQnKymTYL4RA38ucBUACf
FepaCotvekBbeeN1PGw5YyLrYSeIf+vxGTyX5MxzNM982IoGQG5flyawZAow0tdM
GvsWXprPzaXs5fVxy7SKJEj2VrFLMKyq9Nl8m8BjumLrwGPv/df31UEodfS4EgPy
aUTx3MqfHmgfOjDDA4BQqo4/kPBVE+UpUfYBRAcN73sPivZ206CPgIA7JO32qDN5
3YVCJYdoavrsXWsuSyOwQuavY3XLoFBuYxQM3N+7BHNE8izjqskcppEaGzQwmPLk
1S8bTmb9xdN8o9gm1Wpl8Xlb2S8gEzyHFhT3Rbp+2vM3ugJnwZxoC5owMkMN+Pij
XLkU0lmqrIrk3ZJm5UlykBiLOk+EoLd92cQiHSs9V3dHrJvhhfFTWR6rqW3keBRi
e960V5cFdo5wMPGDoeH2gWFutfEfa5yBU6liU+u6vmwpHwcktqmDvzZAD8SLaPkR
mrsiEFdR0dyJypfxUEQ3y7rU6JkaBrL74t6tdPz08l5rdxE+0XZBAzdmI7ys46OZ
7mJUqoQzGUZEKstBeNc6uSPEqO2QewNNC6tCrBCF/dMsfZ0dlM5uOgSe8MricY+D
FL8m90YxJlqU7JBxZm7Z0QpdWVduq6zTJTw1tLwSID8gDKJikjB6iYL0y9xENteE
I+z1Adjt/k4Y40Fw6BhreF+1IxZhmCs/H1hUpWwhCSZo19Z3Kb6u0TPOKICtm9Fh
FjlyLbOubETLfySVFGc9zC0b121abUVYQ80WBOL4wf5S8Jn66CuaqZRYgPEs00t2
2jZk81V7xsUZKtYWBMw3tTgmQ0E2qBpSzbGBjrueLxQ49NgKQibaVZz8CLqQ5cOJ
FiVC0xFR8MQih00Oy8RGGokH8R8ZPmUtkZpuwqs6x7Sl0xW3kS2xdH6mdDttEA0B
N3djOiIBojt9A4wRDtNt9ephFq5MQqKbSws6qSn5mKWow1Ic+pyjOzcu/c1ZQ6s1
MEMfUuOlCnCViumZEBliWk8Q1gt7SpPKFsDg5GhhcKnK4GIXbesVq4y0MXJlEo4K
7j1qO37bQy+r6dxqvoeC4hlijj38WKuvlae5qOxNKK5xj99TxL3dOP2/g3HJUNka
UYwoHjz2vgXOmWbgLnJDm6L/NUJgqq/vbJP/Vh0/HV+Oto7TjqacIiA3uA9GveAn
Cb2AhHU5dz9a4viPio6AgI1/82XrHDLDb156inV0UxT3Ek7yvumDeTzzbjk5rgmO
60vgHXeOXsxXfn6KjtnixXURjxIrgai6uzpnSDrLvgRmz+whdRj7VtjWLXTsYblQ
JXGbsTP103tK4tPFyXFUTrgM+rQlrUllyJYFt5ukRIEAsIvLWKl5TQMdUeyLimxj
b12SaINR1sPjFXD7sxymHCn0z8PWflvgI4HdGZhI4rs=
`protect end_protected