`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8496 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRvSzIdqqwO5JLOHm2ufP7ErxMLNy/dY8s/nYNHSIBPNi
jBYFXhYUdNAO0R8/BBV2l3ATp4QF0HTZH1iwbZCSB2z1/VuiJ0k7MHGNN1OnDfLa
IP7R4cxTXoZMs3s2l/EVAwfrZineQL/+ny7cDtaWv4UAJbtBvwXAuSUePaYQqYp3
vL1GGbHe+Bmzo9r0R1F1aa+KtwvvvtX7ovg6AE/aIaJ1eA+gMRvGAGwoehjeAtMZ
Ppfc1U9WUZBIsgbt7aXKa7uZjzc498DKDBOpW3Ysnx9X0aRMWr/fa34Pp6Hhlegy
fZmR5ruPg/sKTBxh/RsaIJ7ePXHdf7/qsD7auhDlMBF87fAUZWRdu1GoMzVTayEa
l/aCdHmgqzeTuSBZdtipbykR4n5y167XdyT7nGGRTRBDfsdPCo0yjCM8Ru3TNo6C
jOi84+DwfoQBQztWjYA5a16PIzYrnOGMK5iiiJ1IDjXgBE3Rj7jNNRCN1dt+LmQV
kVRqsMc6snV5nrpkBk7qbp7l/cz4A7/NKadAuyMg1T4VVnkfVX1He5Abb0fp/iEE
A+N4qWrCeUeXpxNzqd9pSXpLAMwFnSTMMBQrKi6/1bCJCai1kR4/m3vbDanN/jcW
uUhy9tGdO0PvRD5rgQM16pwzEgKK30z3BqbpJGzpW9YN707dogw7uvPF/v7ee7+l
etvGlwJnjRs3oxx/hVtMTI5jQkxzd6Dp/y1dv9zKw56h5Qd3yqab4bObbPh6MwrD
ylttvu9Tvckg/bH4QN2QaENcmTfBFFBl9/pjKRrRkcx04qh7Qv50DCXjOA2ZZDYp
LPPwqgR1i0GZnpflKayPuGIiC2E8MXRxnCUGp9ouMWbuBHWOwkU/5jch1N+yuxi3
AiCN/XZV7bS8EB2fpyVjtQEDuw+y9vmKUow8VMTyv4jvsj2/J0slyC8LG0mIcePJ
50V2ag+DUo+CUhCWuyQy93GN/xrWV4y3fI5EFrX7cc0apTdmILtKf5rSHzek+ur3
gHqHDgX8Q1vXZz9dkJVoY7gnkZpZXImaHX05Nj+wWGOJKoikl17tEUlCkFy757eE
+Y5s5YOwidMDWlH3l+NgJcLF7735McowF9hKLMZ395hvtRsqStSPTU+1BbA76K0a
QdLyUJ154V5Z4cpy6H3juwXpU7bmBxZesf9f+yQ//7c/SB2AXbhfZWBcIhPuf+XL
w4qhwUYr6JMqi/NFKFnHWhq0lZUds6Ov+fmz2oWjO6eYz+gzMBHB9ImYb58qmKGt
E5e8BGi+4Sg+l1f6vVRFx5FFYH/Dfm9gNgzqs4G2rXqgyQ+0Wn/GzL5xMVtbl5eZ
bBy07Dj61ipy2iWvOg+ATdkptH/FHIwHCcc9AgSfAQv+BEKhve/qnhOxXVHaaF0g
oZbJhRWZUeVXji9NhalcPopMlxMjVAKwjw0BfzSoKGy17mK+uZXJPtQ4dCvyG4X1
iFVcDIwYKbn9L0jUSvJloxiLnYrJbm2RAsnNSOUkjdgiSrCAtMLLfZaLm8KDQ/LG
q3/D/kiO5M+1UgZqQ2mfqkS9Pk6satdQZRNCd7BueXmtU96TSdsRNJ5XTJYX2qpv
fo6ddCNIb2Y+7TNbKMSOS3L213+vSNgPFK/JrtDWAXEGiU84bt2z5LaQ3OitR47t
j0iH/Pgt7wp775HzzZsKIe7tEBsHAXhsBnwGhyV51TC5mH799lTYoAuq15WkQ3cE
8CxQn6Rw59TzAdOCt1su+yJhmMXnIH10+yEpp0I4DQgCj/kssf3cVkJ4CzhZtDDG
lzzGKcofPb1cqOcyxBj5gDIGhJoxPdfr+FJTsDanaVXhwBKBwxZZgYReY75hjCNR
ShxrnqwtM0OZCUJcnIcnDCkX9kXzoI9hhRRiHrzU95Pmdkuq0KvcJnuwy1Z43D1z
N2NHwdwOQ5KW302OhT+VXfLEY5PCpjOpDEXbojOB+Hd1lyOnm/qLl24NyIaHcXM5
7xrmpfsvQ8K4RBz3SR0aov7BnphACCzm4CKLUlFNMDwtUeuWNyrZjKQ+yyim/yus
Xx67WqquGB3Is8ZPWs5EdhWNUUubZUzMkS5I6yCPYRcWCoeM5fURyItiP0uu3I9Y
RBm/3at5GmVtLFPKXBZbImOU9xlOjtVeS1n5fO/sNhHrUy8hu13ifA2zrK+GRx9k
ajSt3INL86clZ1BxJY0/DWKIJq0pLNPBAuhrmQbJgKYVYhXLFm1kjh5UhZDGJ/zF
gFThyJrSUNi9+lgWVoh7sIXBs3X4tSOG3k/UL4WPSRqoyo4DWRmb1qo/2nbCTfC6
Ezq24kCgTpYqqjygA9eYpot1furcKfDCFdkTP7wcBd0DEv3VE6oNkoebS8EqtPz/
ksxPre+hFFPfkBxyFSPNAyO+wr3lkdx9c2AffTybdTPeqiiSCT8Ff57r5ctCwNgR
Wh2nArpUc7moxrQcMalkDiADcGfbsivNcOuihwA98YMYi7Yo4aQqN3D/7RYYVWbK
Qe0szd/VvPvigHinGy+bYAxDbC+C4q5ie7IRVgO2YqENTg23N2GJZkYqEqMmR3oR
PKUmBioohP76sQUEvxENyJZSwIHxECp6NVakyalSfTz0/tNflO7ynVwjTd/uUaLa
242Qn+N9KT9C1E1OZ4gFNlcM1VQbZeI59MIq/jcyEzV/pbkv73EgIHHRTCxTGJ/B
mEbxxFxGenKQe0k7dqS/8NYS/ZVtjSCzU1D/Cz28HnCbcHqgDvsVXpjqrEnh+ixR
85Cvgv294rpjjUxX/rsGeTw6HIJuQe0FhHrZk+8WC2/4AhACUBi5xychSpL5CDfa
vHS6VX6ahFEtR8aBhUGp9joMNpKfMyniAHxT31h6wZaCv8s6ppkJTaVkTOpS2aaC
37zUWmir54TP94+uKW+8yP8vk4OKOW71Udnu1zda6ZWleV3L47FX/J7ZeF76YzN8
JleJmwdjbz1m0ht7jrhxf0UhTQiUv0+4+TaCM76tPT5eaU+MYGihtXSCzUWYb8dr
ZBm2lvDiV1q9DrmNp6CmKWw4QWVSTVfp4hApEx9CZwncKAI4g6eLFxfXiwyVgnak
t8aWzWeWAXQL2lV2x/u7zJfKCEHxwgAINOCZcSFlH2cPg+Gzr2gYr2RWHLZQn0v7
85s32JDoh52x1AGYqiI/ghCY4cyAMlvJ8sfACiLVnOmMcULYWzlasAA/Y2ezzYYM
zqfLRtcno2tlDdFS7azuNk4cSmgzmunPfr18B3eHK0Jtdg1Z2W+HMiCHPwj2U8Zj
rDq4fKRJCfRymbnNG1Ydz2xOGxw44NJMn0fzKXXFkxmmP/43INLEgMlvVfRGszwk
SxNwLXE0BJjjWAlLmBhZQrNoq/+CbMLWkUrMU4rkAnRoSpdXZhccrHHBneDaffQ1
ucZw2skQSv6TpSXDQljf/YOb2H56YU4IUjHyBy1pQaKg1g38OsusNP3BHUoAI20n
68seK/cJ85RscHo2Mt0Hipaz8Wf+K892zlaS6C+UnLtXsRur7zG0m0QoSFuxl3FE
Q4QaxBaifYDfwpGuoCY+BEIhd00GZyhl5iXg7sxcyN2nCe6LmHZwt5b6P4sWfAIh
68lTw8H8irnIWMbtWKMatDTd8K2L8m1Z7PT7CtqmEeCv5wqdt2cUAwol8Od7GB7S
DvczOCujhixd5F33+85zLq/q49q2fgnNHzbCL+hm9/6iKVixwRJsmmYPnWbI8uwn
HxWvugV5P0ra1FwjTywS+Kg+WiKD93R7lT4x4SkjRfcLH4FYiTt+57iiY5D90wqg
RIyq0qxqKcW31c0oPn2uqHxFtgKqMyjtm3siU7hVlggF26GprRhM6+l0J+YheKsm
MRLD6T+FW9zAs3ptKG15QLN68dJ7BvRnDyBkXItxEpzo94MplpxafsNbfpSZE5mF
M6L6bMrpBDyAj3GCMppptiIxI5759ojjfLEBKjOH2ywagukwgJKz/pOKRHFVYmLo
++FpwEFJzzSDZVsIxF6e+kNETDuMmuTdkcg84OmdiYds6t2pckyGNfViIFEhWkVu
4TliY7XePEYM8sY0UMJW+oMSbgrwPwgzWkeVICkcpTbV7hhzChs2eiTlGSVn5rv3
sZTpKufXSVQ4BSc43bMep+erSbH8Zlzq1A6Jgxvx0Lz3ytG1HZjmwq45lK8SAxjr
Y5HT4xAX5rCawtD/a8GHMfpdjZCgMADA6C9C4OpCPH+x6weNEURg6hFR7KEGJsgR
/W0Gdi00AiTbUIc2CmLBKRWT7SNPc8/Db6HchUcxqw2nUGMfaCPQIsq89AhC8n5c
UBAD1V2snGjMy64m4cSjim+VTNYOjgGHWK4SUaM35oQVF2uQ0UPeG02iPsKO5B2L
xWKxNgRavF+7+yAG55kUFZ+gh0Qhzh8OmUqyUPgBIDlDwhI+1yj/Ck8K3J2wToKu
MJ0rYWCfQos3318Gnz0jv1HKvVhFvSJ0OyVo5EcvqzqZAb5M27s8lwNknsJTKoHM
sv1cOyzLFvt17wTIPIp8T1Sy6YmAExgHaLvRl+9VpU7B8gkh7hccawndBn5VASYi
nbiJcdyEZbApbUABCVgYr/tpovdLNStK3oASXTsSTfnUjwHVmKqJhbsF5K9DrR3o
VXVwpzONwPrDubfb2hKWgcDxbEcQbAsTYlc5nk40JzWjZBAQmLFfNGdEdD0Kbu3/
/ZjiNGxgApb7C2/DDAvzheyExvssEWfEiv1KsbHVu2iAbP6wrlLTUX4jHjcLVx1d
FcDWLy507z9dR1tDYWKt37E+5hwXr42hAY/Rr9cJWvdi4DnnwdNFd0sY30h7k8LQ
iS3WI4a6h8e+d6ZXEY5FcChdS0kNUuD2wLzMEvTt/U/ov5OBmGx2OmGpp+uVNBoX
CA1gfMEZoXUSjHYAwEL4o0dB2D0Le4etRP2TJnhLc/ZQxroJ7M/wXnR6IAAakSgI
Ts3QRk/V68bWJA7G+9tny3No3zmo2UisDNtK1ZLLQcsoivoaY34qBeWHi6DLIkD7
9DG3/9T8U7EjBKMWKIdFWCCaCPw7ScGHNROf5rj9O5xVW5dKI8jyZWUUIDDcyAWW
C8o1KWx5YhgXrKFUeYxTvkrTDlknB0Xkg1Z+diZ0CZylkleVSxAWvXrgMJ603h+O
51HEX1FNj6BITFT94IEiQcv6CJFVXrO1kxI5liVyu1eRqec63IR6QfhE7Valk39C
+aBosY3HrDILv5yS89arMI+EIY0J0fgDUpBQZP7KmQ2NtblvYPl7lxjz66HseiFq
Am64wo75yOUIJjum8ZLJc0twv5hQ8ugu+Mvz+KKehPTStUqpKJ3D/571KkifOcO1
XINfkEvS9bWVEiMKoifQfCiTzVfcEp1zIWLEWBg82y1QZIR+JcEBnSl7sn/7lmRL
mMc+9yEHzYxUom7Xw5ofc2nm8cemN2m5S8xkWywgHX5e3qW8LOynQaoqwBGT1Go5
P22HScgSHSdBkWnF29vRl1GiYEeJVbvi3LJXPgT4IsyjAqXPgpbhRHl6q8EnGSjQ
rWh3R2S81RGrkpaPZdQW66bOe1M8w7vbUmmyRt8zDJ2wovHX3OR4FS3ywE/K4iPw
DN0ArMXaxfB4TrOfKbjWL+azfBNSa/0XehG6T+was63FidQz2eYHJMP3nTKCua0S
g6DdYmssgaLPLq2LyXGJ0lxW5mtNsADr79lMgS0ZscUxlF26XhzT+Hh9jDCAGQQS
u8joUJvIcFd8nmDTpNWIozqG/G/TtRK22kxcU/CKltpIhg4VcgZBPKPtErtMihxu
yvRMAl+BiHNHkDtBhwtSI1+PE3GWOfI5rvPYnL7wCKoTCgJD/9sQ1tylCrbOl79O
a1FYucHonb9JjXjnYdvvK90FW+ssJr43T+WCjKpsAklLep1MorxZJA+UaAli+5/A
x5fCSGQ/y0+Oc+WKQW+/n+iRTuHAqVtBD9YviPCZFcW74TnIiRgJp6FbnJNbx94Z
UCfQoXM3aIYBxQTuMPWu/3hOZWnvK4XRqCFiHoqOvhWoIxqXEeU6H8PFl6D9SPTu
dioJ1qDN9yHoyA+pVg46Mp5ZvlbgpYADpK0nR6ERDRRY/G1OKG/TZitmiPCyL4cK
BRbVQGjobfMveX1blCQf68HJI60s9sM+ZCUzo9oGKIyXhfd2tvuUp6H+vfGW6LXP
P4qAUx6efjXW0XrBieOp+elRlMjdshhDOUFIJVTI1pLbkaxN+vMcrL2Dk6YubMGQ
+l2GmozO99WIG2C3GOlJdhhnF27qtZYbDVb/DUFeAQk+74txsuKXnILPdN0XM6U2
6snJeYC0WMF8cihIA4nu96IpFaUoIH8w4x6zbGRq6hYLpky6xTcRMPRF5N32BsTz
SWTDno5qaUoGbntrU3pz+YEuYDNMXkmICaInJ//E4NhI6wFEoFduG8omcNIdLZhn
uJDd3zBgYno8lemyV5Zhwv6rGO+Nc9PWu9KBXsTnGUL7BA4/6BXx3Ulqht1oXjDs
HegAkz8Xo7NWN7D6p6B8boGTuZi/fk4PK83dX/9/9f5rzO1SNR6f7L/y57CXlaeS
9jWwEIFmL4TDvxsjYZ/WVivFpPowxjR8ccD2GLWheiqFLsPb28XNpbY7X0cjp8Or
fex2OsFbKSuq3DbX8C0vxpab2EFzprasBLpDZKF3RKPSxhXo+IrUQ6rjo4cqM776
Sdobqp3ppRHsBTBbH5FkbfL3yiNg9te9dhbL2SUiIGgvyHd3Voks9MYgLxVGjRQ/
HWDBFBOFCBhGKmUlH1aIVYr53jAqs1YlSSP7mNKNFKKkhtSBVsJXUkOzhydepq96
Aims6j9N8T8G17wi1O+KCjBgeJ9qLk835RUmDVUG4YXn2/rAoDp4JPTRe2crsuK2
3K5HwMX8spIKMysKcMPKQHWpc95PpE5nKHrymSnoDq3k4B5adZHJFZvT0LcALCq+
zh5BtiCfOwhCdV3SfRlE8YWM6di4E2f9TgAb9b0OUw6hW8xxrZJYaGez3tkkArWt
jAmY7RRPVByQloM86glB2Ut2DM18z44J81NG080oA9AICbTYGQp0CZkOaMHGBF3e
lFVFIw/YFykV1rOYOLl3A4TKZg4BxistUL1+TQBer3JSt7MKEDXr9jufmufGVwb7
+qduobIP9dHCp0qagLgUHpKzrbzhY5C9otEWcNA8xpbvb6GSU88od3k8yEzubyG2
/5MLYTkitgBso05r6eJ6QrWVXaSZQVjTPIJIQZvjuF/0muKdGjaTiQs8STDL1DDx
crrKP9NfTH4ZNbd8GK2oAydWjuKekN1KFZS5uljSwTdPYH6C0FhFbpe0oIpd0ETv
3+4PmswRc3RUgAfymKEFFDe+F6ORukZt7C9q5bbNrBjc5xxfjAwjaFmJrsH/fQ9f
LgVXsiCRQF9Mfqp+y79+pDLIKX3MjCNCrF5NfiW8fYS9AnEYsjYoU8ugdZT5ygVH
wXZkaneaWd+xFqsV3O6HV2Qjpcb7q062QAjGsOt+TibdhAMdTjYHTpfb7LvSkcCC
fse61es5EFT94nZfKK1l9reKSvfxQ/x1F8EpK0fTqvsGoqxyf64U3wjdnPR9aiQz
z6QUyWj66ABLrkBGB/9D28ZeUNxElaayM04H8XeWR6fHNp5p0jCCcqHcSnx+Ur+o
xDUdp3WdwmilPIfOWMuJlmsesP5wQgwjvYbqH0CzcupWg0C0QUe3k9bxWzQWNzWO
2PbZ09QOz+hL7Ts6Sr+urqCmXDfDjf2EUlL19h1f92B1+pPvd7DANOSJMUXjhKsB
PNvK3b6Cn78EfMECRmYP5Fsqlf0tAqoFGJu9O0lqcZfjbR3+XmPeZ6/aUaEr9jwW
cklLTPicRrbTnpnQZJTWlBmmxZcACdGbVnenVmicPCJ8LvturU+0uJNYIy5vtisb
OLnLH6yF+ZzFIX/gs1BxqrYEJFz5THElIY70yxaIEWgY4XFMlRd9hoorJD+HzSo7
CiZWmmhjlJFWUNMuoA4DDKPMQGKJw1GcX/3ZVGQCdRXiOj/5t4tERcXtTu5V7v4R
uwOJmmYbXKbYOv9YZ47AYnskmWbq9jhuBmEhJbT4Ouqv4KZjATqgJyIa3RtzwT2H
EsyMxYmdKuXMay+XyCOc6Sse+FZTokVy4efUqfAgHYLwdTNVs28s/IVTWAF+vBRQ
IyDc6LBNFDJU0jyhSsNw0n6+DUBpOmcwyGD2eKUdTOCBqs3du2mpo3BF3L2XU7Vo
/cOuaENwx5noNyyGSr4Jtq5PnNJ0z1/qBSHD4eLdA+DjGiZkFZxw0SIQsUNEwzv0
67RmYkmBETJzOpl4YeOkMgpNVxqVPqSv+QwM6GXY48fvh6QzcyqlxXKIPGQGwhcw
3qyIBRSSpOoqJp4+Z9wxT3S+Pl4hfSDgxSJo0CI9LU2li2eyP4syl5bFXCQxpSxJ
NiOKO90+Uiv2BZ5+L50SBM/eHPPpTMFqvSTx6P1v06jtwJPwb+bpoloHFasdS0h9
68zI96xgwKAFtQoOyZIeCwyx3MeVEt+Lxw0ubt3o7hjQP3Ed0tx+BTqGsIqaIwVy
Bho1IiDtgUZwA50swZChcnEPJSmcZn5fLOAo1iX7B5CtQDmEuNXbxqV5bNMRG/PM
8FDRH1+Gh0RCVe9nRtTIcEzxPFjiiNagumPotyXnbRqPeXtV1CmFUpguyajn12hH
YgrotxFpoSjVDCgUSJJLwQJRRE1VJq37wyRyABzyOflp8u1manEgT90l8ZKeq1ED
kcoxkLSo2VHHUdyFDIGyJa/dB5BP2PWooNcL/4HtlJ16J5Br8g9N0DjbvAdhgvgS
9LLCa07gzY+vQQ0IrTkCGcr1/8LUE1T4qcnoz0u6kTby4DWxGT+Wqzzjh7IY2IHB
Wh15QvIs/XDtQnzZHVrxDkUrmBFRnDCvw495hUgo+pnvuX5vKhyrdVqk+Jhyafmz
ky3UNa4315gVJs1RaByin5g9jcSeL9jCixwOKGB32GMLC7Cb+RtGeeWv9b7tnM4V
1tU7e3OqCeydIlpfq+hFy6Eq2+foRPQr0EJaYLKruSQIL2vkiloGtz9c2Bq6YQoD
X5CYEE+3F7CI/dJFbwEvr+DBg832ujKzR6lJtvk6ldjOavYj+BhFlrXt+VToXEBg
pf9fkNg8vQxE2e1LEE/psGvP86ZnGOQwJJekeKU7rtH8cFZmHjusnAYhY/5BGHyB
uX4V3jJFkCSsR37e/4CWKpOLbuOZTwRO8Pj4ATIS5TKTdOfELRl4wLjvMEdg+DwW
XbpG37pq2AP9Le0jNtQP9yyjwFwarKyv6e/4lb/6odfqMDZqQXJ7deh2UCZVEBDX
Q3DHzNav0HQZ3yg03P1MZ8tcX4Ji1/jhK0JFVqBc05SyQTWH+19lHxvW59vbAXro
7WcUohX+jOfOaz64ijWCmAyVPaN0IdBKXK/a0EuC+iKMHhHUzcrJ5EWpVr1UEvCv
34uv6pgPw6mD/MmucQ/xfvoetqhZOhTIIAPl4P/nOXfn7qPIB+A5bc8TR25LTd7s
1grfVEwa5coPQjownX1qcvPb1czjK8fsVByhff7YYF6CzNgH5CfleETtNyftB8aK
aQa8k/7idN1KLOkIz9TzB9oe7KfU1KhR0IuoyXpK9sdbbe8huPk2OCzayGKD9BOf
wszzYfPmIhkYZPwwfRHp4tKYpOv1W0z57+6g+OiHULiTFUS9v1PtVd6AtpssJ+Dj
0ruSerVMnhkRJ8V9QjC3PphMZw2hGaIL+nd8+1yWaoT11Tn6Mh3e5hzQTvWPy1f/
17Ujd8AYtRHOt+FJQQLU6OFQAzG5mZQHI/K+lMr42SFJZOuD4snKaUnytG9DfWvw
jeKoCM2DTl8fDlcZg9MMZyKvsAIsoxTY9B4EjWouT4PEo2Irv/fZ6MUo0JAn5HHO
7l/ilBrLvdVTaqMJO/Epm+PoP2WlKK7oams6o9F6kgX7Cy6yDFHmiKSrgxW9uHyG
yGj56a93e82D/b191W0+0l6RGxYqmKqy673ZCFVZDa9GJ8DeKU7wTiP4SQGMNEr/
MYfD2cp7tlzGbboTupzXhXvKtT4MVPhRhv24CPC8vSCITYIpRSZTRI39kY7h1vH2
ir5UpzMaOYR97Q1WjQDrwmeRZQHff2AIePVQNRfecyn4xPzExNXC7MdYK6mLoN34
9fT3LrCt9eFBuqhdWTa1Q/JE7NLI59plIQIBy4tCznKJ58YU1rpbJmroq80YqAy/
D4MeZWcXym6c6rqHBaP8bJv6TQ6f10JiMuNk84AoipM+Hom4IKm8SVkIxFc2oESU
DX3ewOSn/eQZNa/oFI9hGtHYvrnlu4Jeb08+Iu3Uce34Xjy6787KPheA4H5Lf1sq
TgYowVl4GSVaAUdrudv/z70HHPJ/aq2q9xur0Cwl9wD3Ve/qavfozfxT3JfBcGNO
sBMxqk2TQZ7P2md5sLNSbNpIUNoa7Rtiuij3/KfC59N9VNe3Miqy0Lfe7BcT0uiy
wfIVaB1dT+tfiRI3/N6pyO8m4JCfVaLhe7cYE3Dc1pLRcROnQCOv7cEh17C8DYp8
kR/ZAG7dzan8PRkzAsTckpH3vL2f5fTeL8nTSNbJ7/l1mpUMxEdZC+tiU+4N5hJ3
0sXTMfWyb9srzuk5dpquY7jka/U+VGNZHkn8N7BnfyHVXYqOlhczDnFGWgaFXD85
PcPZIX66kwbW1wa/zKNis+MK/xFC4K6qSE+MUnnqFtnnGwuBAdBH6nIl3jmwqUIX
NvwyPgL4LLZMUVvHTKhW9cA7gMZDGzTI+tUBM3uZlQvibRYj3zideUu4TmZpqYct
lPpVWRRSpvk9AuKzna2LuqHpv7p2xLFVPup5JM30jbYdB/AaoRpr664TjB/uCZul
+AfCycF4AaCsEfh2h/oXH2dcE3MUnoW81Q21N7fEls2kNtGX/qIeJOrdJVxMa5mY
bqrzmhCSJNsNMEVGKYSvclz+6Y0aLC7yjR0NZLg3nYuLxa8sGOGkdJ0BA6NbYXT/
cdkUz/B5jUCM4KHJsmlCeWtpPQdRz74oGjEz1C9tJYlVYmKsBBhXkmP1JhxY37d8
gld6gAuHgPQVbADZuFfRWHqsawKXS27VCIM0KgOSKUvjxh9aYzGo0TTHikEubuIZ
4B+zOTTNHWSb+ry/rM2MuL1J9znBN/9SJWdWzTmb3vNPnYmXFXAjN1BVxIF/9NvD
INwoWDdYLGKEhhJGBVc+DcUzwROqxcxZQJQPK4vQfdl5Dt3hGvSDZFSf9S5eqI1d
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8496 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aXtofNDQzja9NaCJV9U+TSYIyCYjubxSSFgTHi6BMvfk
vMX+zY/oum85alqOnLzQzl52M+zSKzVtDoT9vopDmBJoM0DMjz+jgXFnQ1lfSRR0
4OknDEslfcbR/TnlyO/GleP7OkCqRuxkUVALpqKLhJAzEu4kJIa3/WVbBaRxZaQE
90jNkVdcUcgXSgiiM2/OIQzIgdQAzj6tj3HoSq4Bhik1Fta+DQuT6rZvj3xKyIUw
0PKx+lfqbez4EFbK4qls9VWl1g5jBIG66bFh9ufG6H1sWWzBNaiFi8H8UPiDheN/
PSWF1iOfSRXRUMxeuzEGFz0pUwnvxaGDaOm1e23lTHWskZ4pTii4nPBWCGuEgq1I
UoYl3PX+L+/fG/6NawuYg57wW7NFYAtJ66nfxDVohsN+UAZv+cQMnaklalVGWXnj
HmiXEA3gs7kmK4vk8gh1htq5Jo5oeWVBTX72ErhgaFfKYS3J0CC6/DYhrj9XxD4o
i9rFfXoQCKdO21BuDV1Yqr1qeYCj0nUuUf36/H6TflGUPQb3CvmubOYMf63fXFQX
7khf4qxuq3+FkY5J6d2okv+0PVd1U4pMt65mo6btbJeVuZO2EkeR8GXI85h5oq23
vgNSicmJcj+5GQf2FXqyANc3yJoUYmq+LMe3kpsiIWpG/WkJdsmSE4+XFCpSJJfQ
OLRzGNA/Zx1ejYzhCLc+OQo1rzwzoGNzKS5seIw8FWUD52hT5dZ1wXiG+8+DTFLB
Tl3SMbBNhHfEHlvf9Y7Qn/kuJn3U+bqUYQMy4LN/ByCISJ5kF0+RhtTRAG6Vlcno
/UwTeBFVQ8ZrH/OQH2GvX6HPmfHMFrvuQ/zFIZG91f1FltgnB6JqRRDwe7+HMLcY
InWWaJKoTqyMNE42/M2OLSDYhp2a797yPzZSQLNbPaoZO5vi79X5Ysbb0UqeiLEO
BaiTjbzmHKG+6gyGqqIa4yZHnaleeWf7DoCe3ZD74W6THWZBG3cekAc/XoDozPiW
POCHLwF7ljgldBkPRONlJoLVPMeq0dWXklYaxRxrvBwOH7ECL4jEQyAYZWMmySo/
3dk9C53XjJHBn9UUXOeXa8xpMKDywpZY7MuwRILu4bwuc77jDkdUcWzFt7RqCDgB
bOrfyMYoL4PhvqbloN5+rVPAA/znQFBHiLQxjo3hibD2AJoPgIfN6k6r2bdXqnaf
wGb+pMwkShVisj8fzyGpjkfAceKiE8UzdD1BeJ/tr/1Kla5ExMSMyN3r/y/lggP7
NN2wrel7LqLj2dbTQcQpnlHU3M0iTaswS7ySw2D9By6IdxonPOtsXOFbkY1RfMdo
/xCOSfOPPFE/yc8y7kgBMM/L0/5cF4nlovQG1svalOkq19b4FJ+brPxadUKgbjWJ
zCS4w05vVfbIRJKByastCf6FIgMXti49pJxvMqerRsghFxocC/JKqV8dtWKvbcAI
qpGlsASZhikSja5MVMdMkORjUvKZzFKgCskZrbwPeOqH3KDcAuopHjjOn4lUBZ2Q
8djdRiaQAmI3nyX4o3EJcSKyK9ZEDPG5wOKSOYqOtkIFluwkFiq60h6CuRJdnj1l
e9OaTkZRyODwqt+Ob9V2K/ODfAMmn3SGEtjn8fa+esRk4PXXAqrzXaQOFIbwCbjj
fAtcZMV+cZZtDGU0Okz8PhMC+NJ+eqQgvkzF9JnI7AauLwINXF5PEy+mtNxgqjuh
F9BN1ATFh74TUo5IbzihQUXeYPhWRc4h+ec3BZAvcAaSlURxTmyDCVj/9lMxnIH8
tdDtgwtHqUM5rgw1kvt/vBz/wWMEzyQE8+E70uGBWnkx/TyFJrae9X5DaJSmZzIM
5kkkKPW+YZwBYqKec1rIJnMAayiCh7h9zFCYGeI0Krq0ICycSuHi8vQ80aUqA2WY
zWYpDiAzu9kULERUwk/uD+pxq1qbp7swyrdaw/YGu9BLhtNzqDuAghtJ973X4PC0
hWSNc09BN9mIMHhxO4Az1G9IJTZKeTVFSa0hra2KyHQX8rJoXJ/y4Cm3uymWIKeD
BMS/Weh3VKRE+pS0a4AaOayNWZXrkVPi2oVMO4uX29NUhnMnfJ57VSgn5dplyhA6
GU/pDRcAL1qnQFPDldoHAoLrhqaMWdAZDfocaEsPbeLhDQI0pvUrbTIVl9LH26P5
nJq93t4MGYZsmByGV7OA7fRnocsjQzMYIilVu912BkOf8LUxH8eS/07/8OJD0MYa
GJGcj09luqsIlGALK9sAJjKEZRVITLlLz1iI7d+qdiTzIhfp1T/5f9zoLu0ddp+C
ZF7XsgSWA3k+m5jBVCX1dcisNKfFtewVO2pJF9j/yCh7aiNrrzYqUqmpT9HKNauq
MOubieZdlwQ+eHgS8B0j4xu0KGkVcTcY7b5Ll3jnCK/r7nzc8a6awvc9d7TC4LZ0
peRV8vltf1A4hVjzLM2Hxf8Y2EEU+0k5adWWK0821wuK3n98YzpWZhHTD7T3jhTB
ZkuDUOKs0zkOCfmzBHgE8VzXaOiwIPialqAL2oND1YtPUQXSORDmWM4/pwUNyzr1
49sm2rZqZNQ07wTlduQZX7zs0hcvVTMI3OicEwzjs8VZw+/lcUzljhv0OodKA1MX
EDs56chhzD1XdhMtXgtjrRzjlrbC6VqzM+iBKVmIHYdECrG2JvuLOaIQHpzFe8fG
viMJkXK4qn8SnMkiOle3gGaQmoNrSb8afUf0C0AEHeVAY6dpFiy4qdEwZHIDUBhd
OVYBGANlrmVwFIPgjjK4DoKzt7jsHueeVO4odMxMADimaXpmVc8a4MzWwAwThTxb
srQWbW9tsU7CQ7Lc+inP5HMMd06hmcDw2w23RFu3TW/hdB93PWn+wHii6hx4YtwA
m7gryoSWTx1dwZdwwTGMOkmZt70iMQmdLb9p3LZqkhL/jbLXuczimhP3Nol97a8N
BJmXDRopIEqVWAD0cWMko4Ld857KspiTUkFxTR4Oi4TbXY5Pb1MmE7AeiMDIHQLY
51xYo2UtaM93pfzGSxE1tqq3Wg30KXBE19jIh8L1RCZuVugTKrLBLCqmwL3OO96x
c0wP0UIaGOabKHMnJlo7VHo969BLiOoptWAu6c+993D64UvWf6Co8tnIS+ycspl/
p+QMggHQapW7/LR2PnUMB4PmweVtY4rHXoOoEU0tpvFi4RzCtKl+1utUQppBSkbm
G1O7QO131jQeJLHD3ETs9ZtsC2mFvYvas3Uf9ziyU1fc27mx3vFlXcsM+0aBAs56
v5/tDLJUQwTusCnkhguT8rozxIf1u/kw9hz48PiOteFHX5gmCB7lrDADOKqs6r4x
0NBJiY/hUVOdHYoru3JVvvHOMqI7JS2vFawIW4/481whxJUSPH0CjZh03v144zTO
rLedmkuZITP7RK5pjwGon8PgScE64dgeaoOsxG/whxuK0VdgXOkj6ss0AAlpNjvC
XYOPPJOaZLcBYnqUA45uaudt7gavrwJa+/Mz1WyssORK3dwvguJnHvVUwhOm3xGe
GpZ/4ASAZ5H2x988Ne78YlUn7U+q/8Xzr3Q0/P/ycdFiuXE3Yhb/KgwZrnT8KUGS
z3FTC1WVOTa6pmjJAZ67d8p4ncxAu6Amj06Xv4Mx7av25JPMHfPOz7yK4Gs8AcOx
wsOY+3Me17dl6v7PHSkHTcxgBgo7zavc/Bt/b5EG6TLBLPO7wIIAZl10EAyy7S09
ihG1NbieHmPByHV0hVaeIPCpfHOocJpAKZGjS9m5dBk/4RIcSToluZeCrrphd17m
TsMd5cmfydkSnx9W5G2vVhChMPwY7GuPvxYrJLcJ8XauLKXb/hyu92eDT28tStDW
EutBrPZsu4bPCUfx7GNEbJuLpGAL6USUDq55HhYJ4EUiLUZmILwHztW9KRsetCPr
GeKKKH5PFgDgHplRPmjhYmK68bXGH/duKwD3Y0Z1e9dm6AaWN8qpUgDt8vHO0wUn
NfNBsipohSz4SogN/UesDQcvdUavSljNkHbYhzPLbjfUC1YIRGmqKFQuAJjKYFfl
Ci4s3qGjXuQ4rZf5SwjVbA36II+RPtGED9sA8bTN+3MhPx/J5Cr1a5qMdKGgUzdu
nrRM9kbFXYewgDJUOa0ypyscgWdv0l1TcZKRP2Ull0tKmkjoITLQP4vY1Tb+jrov
aYol6yNn1eMQ/S1cwMDaSkHRPkObj5sJi4bqTj0KFcS9XazMXl+0t2rQjP2egHoP
mrr64cg1Y2RS95NyR+yMB1zMRZY8G3ZlSBNz6A17uRAZ/ddyZutWgj5sV4T6aup+
BeObhPeX3kLMtUI4TiM7IfZEsVjNeaaamHlMbQat7g3AN0UIX929gcbvnRQLh48V
pYlR4nyKrS48lKgkfDisNpJzggUKI2ifBObbgLiTi4fdyCgxNFkuUvYcsEMif4hG
tM5swdfuG9/7fN24gu8aHEWeXBTCCSZTqiHWTrmyys8wzi/WqCEqKOyh2HWULwyh
hWt67Jm9OQMMC83oKZrKRImMmqgJurVHVAv7uqiNXruTzH1CjLj83nXR+in6KU3T
i+l+CMRqBSgHiw2FtavVgfyPtk565BpxJZMhV7lq9vox3g8LacJweaAOVtTDQ+vf
TwMk6Ht3OYD2k9gRKbiwDTGCGeYTF6mbsrd/IKBBmcQzX/43Xlq3a+jNxR0ssu71
kqQ5c34wy1oyB12BURt12heHsP7szCCdtDUCo4fg2vdbfoFO1NfHNml1sxge/D/A
Og6M5grxcrgNwyUIFZdBAJG6nTm7vk1xxuG+k16jRoR1vNY6iXORxZXjhI3WVzUn
f/8AGSld+N5T9aKIE/Vby9V71HVhO5c4bQDhYUXsJNhnm2EHtuWhJ44IRV4FRAGv
GwIcEPFBrszgz7IUuVjlYVv903mMCXjKyMu433he14cTAigzmaOKWI3rNDD9eJqz
Yzp/pdB/OxIm4uSludi66J5VbR6c1fdBYc9/Tgq02auays3WfJfNBfj3YD2IlHX6
fIVPvwllvj4EFwU6bz29YTnpPjphw+YrkKEr1HhEcwI6hpNG25w5QmHPdHwCTtgP
3VH08D9+PUqbbqrvGpF/ErdvsU8MNtmLVoveTaJmuMltBd/yRH+rKydOYMUyXPQS
4vJGG4pMfA+i1oPlhQSrzvCY1cJYwebs56dW9w1jZQddwZzgpHRPjch4nBFAUq5q
RFHcpVm2G2Hv+T7fa7EUGYTWaoecJ+eYBfJ/9xXXGvI6gVJUqub0qrSyCZA2VsbP
lWVwb9E+23HUY5PiWA+Cp4VCTYe2hFtgGsK9HYEs7raXd1OHVtu1AUJaykrHJUYO
ib2zx3eoUOfx3FCIZOj26vsQufpStG2gmeY33hcyUthtzbFqoSp0xEDH0N9jSwjW
VCBUW3nFzvfbUDrZniM1vxANbThoZeDlXiexVBuWS5UsdT5s99fesu9g2dr1jSkS
Av9suSYs1nPffOIIvsq+tPddWtYNyhubaPZFvy2IM7EeEk2CQ0JetX0cr/p6xzcA
5xJG8PDwfGq6GuY1dnp9pldbizgjB5O3+pSZwIqxGf7mW5ZrSmi58cJWf19ZRPq/
wpVmCGFbYOxohn7DFrI842baEcSHo8Cy6i3VIposzOAJ7TfjjnJQxY7QzKHENeRI
nWXRQ4A2mHhIaVgRvN5r5/CBUvo9Ex+xhmxfa/H1s5JxugB+pjenGvUg0phDTE93
T+wQshgy+uyqJ8EDQLP8AgU1ME7rvkEw8ijbCVTI8qUirHtJwHsyL5Q7cGHhL30C
EbM2fWQ1MD/1jusaIhN4eJN3vVhhB8OAJOigWfNIKV1vfYkWbRDE5pFnD924Q4dv
wC2+BmLyyKKdMG8owTwqRni5+hVAhIhpuv4N1Q5pLwtTQJ9VjTSz77KZ/jA0lttq
qAHQuBuWkGiSb+8wFKh5fIAIGuT45Hhbm5nxt0YmMLl9O57p3sH1+kbuVVimP+zH
v+WJqA9S4ofIJ+KaMxTvU8SVe8jAFuLG62Yo6A3OxsOYYQCAGn8Lp3/6FjNxm2VI
OfDN/W0MpLxTHEYxRMQY3GYwJtwcLx81KjSA2DbW8VFuW1KQLr61Rkzz3jiWWEbA
OCxBjZOOQM94cjoQ6i3jAr6gnkwQRJvbYrGZTgn4Ol+9XmkNVUNW8sk9kBNgnIVU
cUFV0/MiU2JKvJy1JEEcUloL1VD5k+NMRhm9c0Dc3TPURkMG2VbBgNF2o0w62nYx
J72mjh6wVzk6wD3ToI6n7yRltOr+XJCv0oXJCJyY7EQ5LsTkJsfd7d5MD+qJCviu
GSOBlnbe2rjxE+tZgXrxXA+5GVjjp9aI19yU+ZxwJL3YIhfT1WH/LV0hTjybx9ER
AnK9EYzM0XyaCsK+K6fX6WUw34/2n3A5mV+oPO1XM0/bEVptflpZ1FXx1BlGRCWT
bKETAelQij2uwJxntj8bNlUfOAtml2GD5+j6vQ4VSyCzr0ajMOex+ddCsfNLUdg7
sBHUYnCC4tg8nYOA+mD/tlSc1g89J1rOUI2oBB6qVJmvvy+oRVAtthxhhXhMDU4H
nensbCYzKfI7mNhxN5E9qhmlSuWTTD3BOa/ESy4V3aGQhiZgPU40WeSCzpE4yWy/
vp4z3W/pkjylidTERk5SlVSeqxJzNYuRzgUcwQ1i90oOGRtINdDNNYEOE0eFBt3X
skymgYBrsyXtgA6T5OdUB+ta3gl8gAIEnch9wR3sSgZYzy8W7YhvhPV3gV5GSajN
1fVFHdnBVixsHA6jNNkt4ozaOcMAqnaz8SYT0StI1WjqZGPTwCjAz4N0oo/CfiVP
d/1DDlJ5BVyx5KHwD2SunjSqN2H9pmyt7Iwvo6ZiOIuJk87nNWxFhYzGQnVgke2s
zLsWyQlpO9y19Gnhpk95omCrD61Cr15ujcgEhhbUMQ1w2TDaSgcmFmcl0KE4YGjH
BXFZZ1LqewV+B6RYfLGIV0FaIs5D/5aIVcZybDDJ48LaLf7qGUYwZzOdJinss5I5
8sgIeOEZoeAL8fm/Zk9A+np6GQIysDl5rztCKdCzZuNyq7j/vGXWl6ud3TVuCDPs
uJa+dkZ5gi8b/JVBI7PXHJN6bx6ku1x1pR8NXBxjGKXCaSK28iN7XV4xJmlX+vQt
YKvSJSO5pcNCMPDj9s9XYHDYkH9ImDn0m2gcUzz0u5WBJ6avCS+rolHi6uldfOwa
JmlmU2iHemhRs9g7Qsr5vpaTmnKfcLAqfNjismOyUrEGqfjnDvn2G3gkkwkXUCfC
HpdsHmbWyqq2o5dy4XuFYNud4Gq9e+M/2V8voLZkmsrgkxKO4bUFgETtG59jOQB1
I9nw9rPnSiZRyLITa8BIvHYz8h68K/WDvthZSEr+hPF6xO8O5PJzcmKKTQ1YKKAP
064CJSMz/9288ZLIqrgX705kedLMdDm620O+8QeweePkeB/FbQ4kDDOarYm/ScIq
3h4PHlwnFzJI15AkoAc8WP8Ba+dXp6yFT/YLCe1hdd/+2SfcdWuK8iKmAOBOE4K0
OU12lBw7YUdP1ahSBoVcT/l+FKTOaWnjwv3o5Y9jmx4VtuCjzFK2lOSUxDOY2+1Y
XkDREumwsGDMxa8ZOfQSGdLoX/mS3wSCEz+JNk9yxToaHcrda/X1LWRJ+bAQjf4t
Ucd18ByV+03az4wsKuzSQUZCzU/bmv4F8RzpUMqggS8KUn/J/rYZ/qQcvlOPP/lF
Pqg1pAVgn5UnSQIM5Dhb9G9UqdeMyiDwrkj8x9R3l+8AuEdn+4BhNhWnKor2znS1
7W4GLNUbHRkS//hQ0hsbiboKFlnxtQaGpchsEdpBpmZjQp1RPC/qEay9Az7tciJf
W6otIUDRuDDvQCvDP7ItLTZxgzrjGRO9M6TPojuoed28mF3yzfCW+1O2nsdHaXH2
7USOjPb3NXO3M1MCFGht5Dg227uqCts9uyNzPC5t0KPMghKPvUOgJCJL0lKh/rax
x+BC3VgCkpjmXVEdsOPltNjwCY1hUOlNZObX6IUMQAFIlgwwda3dgkUZqiMPjtfE
KRiLGBpGtVg2ELQSXGU4CaJMT/v8D9opob5MKTGZ0sz+GY7kJeXGUTRZz2VjlKM4
vkS1qflXffc04IjmZBYleHeOYu6mcgrO0e42h3mZAAQamVmkkcIvr41KgrtOs14b
qz8nA04G1ps0JXUeq+AbbF9G4gcBVhj31b48BRgTJL+5Ez0ysbfqgRioSp3r8ihL
t392FKetlNpCzrR2Luw1uAlK64gtadevzMWd7Yh24GUjsl6HzH6M8TZAmzVnOATd
oX0q+fA89Gg46LIfitf1cHqxG/i4ulOpkp093MIQUAVfI1tGeyOe7EdOcJyHvKPt
jWOKP5TezEZ/rxhlbrxL6P0Yi37rTfRGqgbWgs/pp2YDkmzQU9cEPgc2M7c6jruV
6Ky94PPn4m0FXf0kqHnTPQw+u66RvE23PhO3VZpXShg3APIYz6MZSFKmv2OzvONX
efXkLntR7NT4kJCx8rhTmkm+uPsJxPTn8VdTLRhxw2lYo/qa3+5oWB35dv/l0C7H
tSXvEjBWEf/Zfx5bKQ2RALX/V2nQiYn8jn9QXeWCb/cCaTwSOrWYno/q6uJr7i6C
qFo8zrafncq/pjFmuwjxcBnrvNc0EyhtYMkn8NlRsJTTydN400rC7+8bBEOYT70J
muUq6/5gajV2ciDeg18OdtTbQ3UPcfLIJn78kZXXF5F4/x2LiMCLCT3ln40spuzZ
gDz1++fHq2zHuMevzMLPcr+iQzd12mgaVNMLkpGBX4M1WPdQe4ZKViKETYwoVsCL
C9lxd3MAqycaTRI70/nZdqh1c4JmM1PB0FW2wE9s3ivuVhmbS1llIgD+Uuo2WVis
D4P9E4RZeOEubwaZdRJSJD3AqbE9T+y9PPnEb0wwWCyCVyYscCnLMccZHI82PVb3
Io8L73F58KKMvbkp7zBbHHK49rnonTANzgrPHaciyBXKQ3MsGJJitKapCj9xRcbH
TrMHaD7ZQ9hJGrq7eV5T3n5gh3YuWACf6Hf5bkK45nh0lY3zE0/Guq2r4lAdpIbq
Tvdo7xAjWpo27ueq3I3thwYzQKPWnSKZGzKoVH2aXcpoDaf6C+28+pggjvZYY9BQ
l1VrfeqWjW7JDN1ZiQIuXQzPdJQQZ7ZbBT0FQQ2UnxekMt1vUGEiYQX6WUZcZb5a
/wCoHL7wkW5S/fwKx1vZTPlzGmabWC9zr+XKu6LMloYebY6oZXjoJBWrtv8YLM/y
85B9d2fEyoRgOnGtcxQ/1D4z3nh4bqNHuLTA2I7EkaTvUl03F7qRx1QrPKPSUp/8
f1lVZxkSLMl1oEnwNdc+5bZo3SJ9ZGDrpk9rZdQ1+DqIgvYqohgWPmRYviKnbSXy
P8bso7chfUyp1LvPMZ30t0fwiAL2Jj+WI3Ut9NRQ+ZgMk6+jqZHZc2qZcsBDIIr0
JJxbvOiVO5hEk6574IkGS5mFyf59NPw6On8lisU0fb5C8FVyAMQPVWD+9H+H0aeB
68DVfNpa3cCO8VSdbW5ZrtWvqVU4gdM0FtQdVM6dDRiJBUVqke8EbtJQc3ySn9M/
RODBWwW1x9CyT046+Z4qBQRg6hEmDZfH/Il0rg0MS4bB13vzc4EKWFe8OixgvZRa
IITngZBtTC/8rX4zDayHpivZfFiATRc0PDXEfuPrmD8tQPXsUJBkb7gtVZIfaL1A
o2+cRWH4nyee4CZ2dYEbOGweZXogdMT+/gUkec3YeR/SdP8ORlZ4xQbYLvTHd1ry
Tl5edDGJpOLsgFlVDwcrSkm9hGw19w6LC3NhxFTaaIeojnFSMy2iPdNEbYwnfT5E
feJCAYKebp4VlyqcXml5oliv7D4zySRfy0HKyt3mpOr/WfG0Zkc01L/mQNXr4U0I
IY+buA2kYUgMAU3bSJOAL+VN1A5G44KjzTqKyPcMBGbTkbwg5bnEcZIX7tNwll8X
hrBNrOou98WQjFzpMAB0U2Z5xZaTZFDjrIFIE+v/ZXGtO6LUP98eEAN7sFq3c+D7
IJwc/lAG6GOlmIER2B0EkDY8T8d5UM7K5sVgFZfwclIj3Mu4bRZwbbhVHbxSmNiZ
6HfehQth84xzpclX2GnQYn6lDd/oGbRzL/KZvbrLvXknWRC7r8nmmk62Hkg2Fj6R
rM0m7evxQoYzBo3DF/DHzb6RBBwuUeqAyLQRwoE5x5uP3RkrpbL7oobdmgoaXG3g
qSHBEwWbIVVMAg+HD2Y+owwU4rvzJk9HAzQAP8W27Ke1QzFNZS9lFSU8c+xvABg+
24NvoJzaecSVNRUHYxeoFmHPwuml8B25gmSu56a7LSg7fo/fdzmgXUPx7RffX7tL
zFuHWWmmsd580CXTT9dL06g0CSHfQMlZWxv/w2XKrLvup1iHP/ZkYQtf4cf89naZ
XJHv3GRnDfNJoL2zs7bqbmB9KJpn+TiRHZatZt/HlVfMs+jLR9i9vaxlN5+uPAAH
Euiw8+BTEKFCvshD80xeCNi1igMsVNY+PdrDIe37lRp4X3lz2tb6ObYUgBACWPgL
M5RLaZlLxzhVOyuRg780BbO/CfvRRVybw6sqpoiQjsAs8CRCfMWREidz2XyTwFge
U4F8PVYOXIZHDpfy7d4Zf9ec2nfhU2As3BNat2DWx25WVco56fVPKhX8gtM5nA9L
A3pztB4iYsXjdJ+kDVwHFJuSZeG3ysqGqgMZfkEXbp9rnJHFzZQIKRROhsocGgSj
b7o+gQWDw1nqIa2FPB3F+x1hXmNYuu1HMKLn3KMfEO0B+ISpSfPMEixmx4mm3zml
jRKpl6+E2zSgApfeqhgmBAL3PYMyTwQ8nhGJFvq72iuSzdxDEgyz5ROicv7/vMnA
zGH4CsUR/W5frvc3lOi/1Bt6jEGFkdW20P30DFG8E5lUDrbFxIix1Oo7vCfYu60C
yKTxYO4WOtt98qOMv2pPzmuCVty2gOsrRBE0MhYZm4GUYh4hrr0E5uKqAyueVRDw
hftRCAJbsd1StR4aqBu/LM55twv9fFi+NgFqAglFgFDyFFKMbxPBKm/w9OEkcNaP
VnJ3oewQ21Gq1EoY+MhITMhgUjb+9wtVL7KtKn/EjbyqIw4la7sJIRksa0RFNc/K
QYPwA372zbTQrgx9WW5VoOd9jJsOpmPZjGw6ZXqTiUMWCctWiKSFb4J5PxkcqnTz
q0fga8sL5ZZOtGzQVRvr5i6YARxlVYjV5bOYPBJZKSOhzNoKc1jQh//JDqAkhPNn
>>>>>>> main
`protect end_protected