`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2128 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ajdsGY4KSUwqrig3jFMVPxNrywouAmklN0v2ERB227uYv0X9XyYNwGTmx4tIoH/j
xNlx/b8OC5YZvO5vxNqB53BUsjpa70JOurKI7hl2fGFDy7Ld6uYaXb0k1cJlKtPO
bzYmuZCf4Slgd1/x5wTgnVbAHNZEHuz9Y+ajlZ4AvSZgy/CoBasRMx+mYVpMOm+S
/lfBLLKEO+MqB9Z0OAkPyf5nG9U+schnjvJZ7WFyPF3IIfHuJzHF2YI8UDeB6FPm
xBlMTT34VJYfZ/0nYOTO0LQ/s+zO52O8luf0a056P4bFC7mGd5P9gXU9UKoGqDWD
feQy2KZ+gPXEXpNfy03nBVFss2FqS4bfFQuKjiohJGiKm6zYbiLktVZTONGooKi+
c/ixGgt4i6ZBu6YaC6b5eiRglJ3SKU0QJApx5ca+ZGNBVfjFsQykbEy6+VUyZXNT
MartPhnI3tqHcVrwV5Mf2idW4vRaZqnTdhxHMEzkBvoDR5vtHX5imNnzbr80pVs+
G0IeepgvmshftE+iYueQQEGvWuLzrXYfA7tFw8lLh5y+4xEiEM6L8fwgPBbtixat
8gcdUOrvrZ2IPCv36kOFjqIfne0PgADqVSlzSdzDdEb9SAMlgvuuuPKmgDyTqKYj
D69pVy2tiqXofzZbjciIiiTAn93vbfs7+34jDfH3n26ohfZwhMbOo/+tqrndjIuQ
IkfEfFm5Jn/Du8pIs2Ix3xV7h0KDdILLicbheDeA2RK10EDRVrV4NtKAd9s4WLU4
WTu0Zt3IDO83SVNQirmitmjh5bNffKWdeEcVNT9Qlj/LpglFL8Xz03siQjpJaG4M
wrK500hFDvKxKrBzhVpW99OudFYxrAigB4ZSEAgMlZAyarHSYo8UWD4xFoQxILdK
Nn5O4eE8sShi7uixc+UqjMU8jjiY2PDwiGqoJpNvWp/Bc8wHjhiqPsGoXsNSroUp
/qQJJn5IOaFTelHcrxdrSBFX0iDr1vkDwles0iTl0zO6S9v6ssv3XjxlXnKpk7yq
Ncs098NlMs1/Zbr5LCBjxq/7SrNrMpQozNjOPUxiaGYADuNBroCPXN3tU+E/Zmu+
jaHsvDsrendwpNrEqq4YlK1EgCspvLdjGjxlpruXuJRMPZMBQgEBOhGM2WB1ZruA
ErWqwLDfXpYZ71fmWdvPMPZWRXSHkMmCMD0dO6ee4YJi2J3bUt6MxCTR0HTJmTH3
0QCRxGEr7rezpzZ1mdLXzg1eVYv+BNJfB7plAQYEeX8PDwArwsbFrIdVvKxfV1br
H1E90aXpdiSBEPO6wU8j680y2t2pScVjIfc5r1/JiyaWXTdU8qaUGZgCz18Ba38I
dYawcKnvwpZ02c5wwQbiuEhKUXBSDA3ZrUQ9RaHzQfr4eRmkF4iHyZ86+yQe1r+u
1lyd52oEC+K3Q7MCycRjJd4sNacJcCrVwV0xjpsFs/i0VQeTKpwoEazrM5Cfy9ir
R6M5rZ/uJitCTtUbhnmhfMJD0mXcWm8MowAZBASo22hn2CwnYNy0JF4MUiRygQ/U
heEaLyVMalqqLueAzrScAkHr92YdDDN8DjhHo7XkZrhlIkwzHJW2gaNlWK1L6rq9
l1XSipUDL1uzzJDoNHx1ECsqBZ1l1o7q8DGgcb41KpMWqfjRDP69HZUR5jDu1sqS
XCBq43gsvYMi2GAgDHsE3/kdxWAjF0UHlFA7NB+mPLGzxG73tarvVLTrJau/Tb2w
CEJuL64yu2/1sUjMRnYTzdLKFY+9T34iMhMbZoZnO6GTUO7fD+aCFgZceNnQ8ONK
pR+0eoYoX8AgO4Cb597w2pN5wh/UR0BOj95YZHc9UCFObx2SzggWfuoFtC7T2knl
yx9KufkeGrgcVI0wWhxWC3tQjVbCxfS6wSROZpuJMWIyICnHrMJzdllccPwQ2GRt
JBV6ZvyroAn8gJElUbAhgKguqHwCanmQd5zl09+fo7MPeYh5x1Jr1OS8AQ/1WRjL
btjBK0bA7XA+50D7K5I+wfoJML7B3ttZGln0d9Hw33O1VRf7X62Myde44awEx1HL
2jj2oHdcuvEa2oClupr3cRdJ3p4PkFdbYkNdjfH9scKEcdPssV2JOHvbQfkO0AVJ
UPlXQuQUXjpKdV5HN9wq/8jgH1pxKgeeIeBaYLTcsVQzKTm2y0D4P3TNJJ4NKPH4
PyFZUwpLnGYQWXBcK8bHSRCW2hVJ5FJ6GMZ7JuuUYrJu0J0lwt0uR6Tz59y8jUMS
MRY8Z6hoZ0BZO/A57o2WujGxA18PxkHuHWv//q2+0IYUcp3XTHTs6/nOUn6MlbBK
ybbEyuACbyMbnCcKnDakNW78BamQJC5kc0Vtyyptkhyii2QQTqEx0piKyKOfxifA
3/hPJ0SOYbSIIfrWad/2E3q6CDZObM9lssJiQOTvzmJJGe1cQxxMXNLXpL80rRwI
DN0HsZVOsU81J3savlmHqhYpY5kZJUB80lzZkDnyDJI+zt7MqWycX3ign1KSjlER
1tdMvaq+jOa2kFXWwyUNR6t9kGuSHd2WmFz8Ck+z1DHsyZM2rueQ9e656ZhpWlYJ
VERE8Xaqgfsnhaksq3V62ZKRj2RlLVsiYPPY39eAqD0jpygO7UwfVvkXe8fG3oOX
rHm13j8Ex5YK7iUwMhWvDPGvCKr2gV6ZQB6auLwfos6i0XCEEx5O4ZbbwZIw9ux4
wf6v4Q4tng4m+61/YXjABw==
`protect end_protected