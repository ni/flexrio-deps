`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
hVdJHWSfELCmA4ds+csnOQAALbB3ps7EiTSHEDd//nts1r+JQrRE4d3bDPRJpiX2
Sl8d+xAK9BIi4i+3ruAzYvB6kuD7r+gs02Jsvd/1kn7JYK4xBxCjtdDFjVHOTEl1
sSh1oNiYUwLuwR1yKfP+xBhqxD2Dv6pCKhH1NdGilpJQ6cvivGkSunAu0tzP76T0
4x1pB179E7uIeRplfHWX03KzEBF+eVtfgXVp2W1BGjfAe43y1pCvNYZOh1+TY62g
EgAFgbo7pAujZxZy/YSiZjUr2mGp7o83qMXyusx8+rQ41D3X6rxfuP0RiId2pOpC
6oq5Dfkx04a1dk4s8w8cVg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="Sm9DkM+kBxuxXCFA+l3fFkxuSWV4xqRc4Nn7Ji3ukao="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
m2emGBqRy4AuduN4dffN8194qYvc9UXRqiQc56IrQYMiIVQPyh59I8SYabcDdspI
7AFHnvKD5YaF6tQfxWm+mlcmMEk2Y//aUjxeiGGs+RkKgbHitJF/K7nqg1dmKvDg
a/GaBCq4Bqh0EehlN4ntP5HxM4qcvSfh5m/Coe3drc4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uG91daMWA1mGkhgP3oZKMYye3UAomMWgG80HuuXg2E0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
c9NqBF2D1wSep1rW7utzHsk2j40aow1MnrccxUTvKej2Q1cyeDDbgAml4eTSXI8z
QYgCADtWi7S8BeChdv4B2VxKcS7CMq/DaQrOy1MKTfQzfAlK0iubmlTkljLy0Rwd
Xim13c6uwpYSg2ONMAUgYaGs33Ur6k21Byxp9Yxm1Gaopls230u6SupdOaBDKWcD
ylbGY1zIS49RZJIPSkT5CkYkZRrsy/zB+TprtSR9eXiOK28SxBjLebOdxJ4urbzx
FqxgpGWLSCCrNpjCjPGZEM0EXodOv0/uzKWyBIgY3UNME7ew0UKG8lXDz20seff5
BL9d7hmtxHqJi/wKx8gEgrZROhZechxn9b02GErP3jrul7lsgDkMRAUiYkEHJAXK
zDJnv0mKBfXhOz5DYcPJeughR7XOO22h2hDhpbIXRGwqRKA274H3wgUQXfJLpFgG
JklRUj+iwaToyXe1ofetRT+Z6dvcsVbx42aGQbmtjRNT0Cr3p5uXP+JCzXAerVmS
xKhVKDqWYK3oUGqr2ieSawB+sKFmIwRsghTc2wDCEod4yIKU50kE+JLxawFb71wQ
e1iNwNb8A9slWNmnyk5g0h9GTB4/JZjjD20TqWKtcyd9okf0CSJWs/q8W7Niu6Ux
s+CIZRkVn5qK5QMcEInVfdpsy0HW+VWned60i8SltbCPdcRbXQM1kovKCIQfVjsk
KSNVtNi0jNpV+7RaXv6l/6ZZeh+RKaFh2txjzRzPt/ObXr8Q9PQCnTIpxBuhMzBy
a2l22MMKY01GNFnv6pjTwZ1xYfMyCVtpSmftvjJic/zthNlIfgAS7wwF/eYUXnYx
tpYXfTA0cIKTDRg0aONcDAIfkOV+Q1uL2SX3OnFgql0kTUsGohhdqAXkQh9iV4RN
JCdeocty0UI+ustYMI+hdYUQkFS0wWl7MJLjJrUKIQEKIqdltTkWWrEkCS2zxjBG
dE8E7hIpWgiu2/wFW8KCtipbiln11+EdiQHgLGuahiHX4pWk6Vk7n9W3yPeMEk62
4/ZnbK5YxlRYIopORfu9dhcu9JgDTjXHrfjQnrpAXGw60T3TG9yvmcTAPWy5ZJX2
IPae27XVaKp+RdafysmAJoNBBzDJdE7k/YpiYc17sUetSJrL9tDjMRLaGT4zrVCY
rUps4KAmNgGeOkEp5vqhLzupkw6DMqCwLJJCyR4U6+0wbcjNAu2Fv4Wg9oQ8KzKW
8D/61qVWs+FiJidsM2w1NamSWrTy/hYQT5qYExMSqW7gumS/e8/0i8r8XNEmemxV
xi3F1Ed/pbbmTvLYc3wfvHACmw+Y7be+XAiL7fnUlc9tcWta4ND8sNcpqsYb7+kv
SEz/JEy3uyP3v1cLtU5KvMMBYBnzNvjSaVgJ0b/rtA86gA/G2tjpA+85gFO12eNu
VWTDkCZNjtJXsXEQUXniRkfO1g1jLHsayIOQf4xz9x0nNu2gF+TeHAy1uN5VRSvL
yuYZL3Ptj4zMA+Kt4ZVpd4H7QyXM27FgjUB7LEPMJQL+8xHvm6CZzCmfjmJRsNIs
kVPeQ7gXQTrSIsQpgitibQ8lWWDigzkx/ePGN90h2zraSuXNWIDaJ3OYAJ+ygjwL
7QiOhPdDYVeuYkYjyUh2fq2Vpj00EPid4OAs3I28wUGFAES6xObwmvtqJ+0Dbm36
KvG7i7hVn9Iw8Ar/XfJj9cXmRK8S72Nt6GnkjHaGbUCIpsTsAUeROuo5NqYcDsdf
4nDzQR14VxgQLPhC1sJ9F4r2rr6hDIdEjADARvz8bI16jX8xRKM6T1xnnJGHwsM9
xYsbPeUdc6kQhueWcqhs8q68/DXLECGjU53d75WSzRH1f9qfNt+0ncAqtztognb0
1ECQBVE1Age/wcqqf/M/VHSA2f1GYrOc4JoXbaqV1Lsfg3Ib7+c/AiCq7Y5SkDMl
3RarnBN5klrDlQNwOI5z5wrLRvXr9I+K6FCqWqW7artuY8aOqoXQXwDjaWdpNMkz
iMEkTMYvhe5fWqePMpT/CafKEzYvM9EXyAfk7TYjZzzM0okbTio07LYRSqZHwkXC
TBN2o1o1/fDU3YSry0gac63SiMFhSGKuhFhyffKUYEdYtjq1idyoqsdwuXmjxKwi
8q3BJEVCEE4wuZeeHxT2sbNa0SIjPNWUoBQ4gQO1pQd4cD/GG8BHqLubpsUwebyA
WyBWEKaowUSRjNVGf1xM6NyjaArg6fMXdeFCjeNJ35FQCE05yg6HyCWsezrQc/gd
48kee9OgDp8QH4ta5QjWl8b7LNnr/K2NEad1u+d9c/LlSofC7TTDtLTdLPzw/S8K
xGXofNVDGlqed7OcVPVRgdyHiTR3/nksmjfZXHWNrwPfGGEY9WDQDcnkxy7oDYhP
wK8mKujUc133MiAW5tI7LWAzvq8VjV90ddChNRucuA+p0kk+spscUJgEk0VtBfhu
RcP3c8ksC7JO0HfG42Oq4qkijjSmRcfdpUBxQ+LdvFRObUhncsEvi5uwZ01em+lV
f0k/j730x5RU10kadW8S5cFvQ4ugx0ynDl7rEFQn/746uJ6w5P5A6jGD1/37JnCc
Gj6a1rkCHJb6cTid8qmbpy2SrYZ09t/jWX1VSpyDUVpNawRltUk/3jFRWCu8iICn
3KX+8dfze3QEx/gEqiTRL/fxQPp1FTh8us7fqz8csEMAt5NMBFyWn1ueV+Dqa+er
Hsg98pboMQgL+I6V2IR6xDGhmEY6GsbN0wf2vNm0srZbmwZR/XkeNhsb51VTO6Bv
8YhrGmcM1wyUhT1B9UBKmaSAMCSny6nNRKuHxX7eTf1lzCu+FQC76GLwjFCeYHms
n415jmhaRRWmTNC0NbHB4nHt9sYBm/xyeq9XqRX4W5ztJT2DDR2ZLvDWMZrx0HP0
ONvw546JUjh50L3Yd+Lli6MrKnHbLixTVSuGL8iiM6TL855NtbRoq7Vf3thLupzQ
DB5W1qcthLLbff9taNsxoP/IvhfJUk35Zc6jRu2QD30RQoMyEscrKmoxi2LgnWK+
/g8IekaqQE20lkYNexn5Od4DOAIAP0pfqWI89R98VyhJ9D1O8gp1gg+qLD5UjgRG
VhmI9dSI6qvA+sRVSMjTG3ZcVcg3yvJUMOqlaVKb5GMs3phEspE28fW6nAWf3XSJ
tJQJGCCpy0V1Xqfa6CnUO09PckD1e8rH0NtiWWhU4XOeUsEZ+c3mvbp7mKhwAwp4
LjF7/lw+BcC+LNldbjt34vGHLTZquUfnyNNxsGRm/FQQ7OkyS1aDit8tlgRaiq+c
cK4AyRKxPWmK0IbD0SpqHS1m/zlmuVn9m8LYyStvqZoS151Y6FDguLtroWNhhzR/
rDUtf192s4T76f6cfTU1fTVDgrMqJienEUjxTG17GpnCShuLo0bqVtt3edzb/XoL
et4IvsyvkG15Ff6g+MykB1CiuxzZMaQ41gPqN2IFJ1BcZYkuFq/lvt3L9Ru4jdHB
zz04ySQmKql8xcXuesKeZXMt7k3Lw2AqR+4382J1dNN6xVXBHmPz3MFWLzKTOeZK
RL4tVMfxe+IFI0jy6NzCcY9lwyjkvXNWyiF8hMem3mb+FKhwVE83mU8a1iiqEDse
vKq12f4RNp3ZwHgcAeILK1kcjvpgKE2xrzGy5G0bldQBkjHotpk0tGFEv24giLxb
XYPUVJxX3oSaee5x1dP2/Eau6Ml5ZYSOakfDq73lA6K9ANV7ypOM+5ho2i5iHvmr
+1QZ0wGfFe2U9Tj1R6k7iWzfwi8FOqFXHiXaYNd48WFOv/SetlNFMp5nWkHoXQr3
IPQHblhOoYlUln8QhCWGbmM/goJiz0r/jsZ0VbwFJJiZvMKWt2pX7pHOXCOoOzM6
PikQC5wKJPCpZVjOScRz/4lcSkVHHrtpnwtASk1MdQ+/P/gIgFpIMC5wW0fD0V9L
9ZfPjTaYvUnJBp4JYn6YMavbQQWBTXM1nC1kqweOVrW5BTsle2+c1iZrAD5+sko9
8Rn/STDTZlPzR9jqcoVJaLvgHeDRcChmfn6q+oIHkLn359fouCclrZ106OrWZxe5
T3xd7tll04EDnVHXrtGr0WH5VhsAmF5qXqSdmXahorUS7HQGkTFTifwcpqZ3120C
Apf/dhNlYqHRSMs/FcVkRmOQNC7c5cHt6lygYQ0Hg7ZV887CvVvf2jC82Q/bhP7p
/7SfSRUtaUojjiM8480qzSxnFoDvGluWBfPXWihdR78Mj8kIvMaWhM8qbz7MVjCn
Iy67OMk45kbYp4+sRF2UnK2w4SrZjRGCZ/S3/QmXFN6FZ4HeujcsiakzbqIW5FqI
O3UR32AqgX6SGAHoZKw/ylPYikYgerzO7CaHAqtvv+T1d8TMPbaxJ6pFLpeQcxe+
35D8z/R59ifcZn6JiH5cVWHl5GZzNXXFWAYvdVP90pmlYiJpBUd64w5MsvyT1CLx
74vlMsTJyuZ2KkkuIbcs6wMXefAJ6QNjl0u2v6q5tLO9lHIKjcNQBUmWuiGiEzSb
doG0Jl+nBo/QkHrwkKH0AtQ+awLJ7lWRsC5SSoKX1OxWLpBGOKGgg/4esbmKkvEW
j70pi8H2jX/eGQ1HbmKTBBrWH1iMZcu5NttLodaUjF/UNS0n6dnslaa8HD88e0yl
GMc8riMw769Cs+auFZmZvBV3mGkFHZ6lNy49+bEVsntTrZTHbsDF2P0bfAeck5DH
2EibPs9DeoUF652JJsHpny4N0K8xDQhC4lk9SbmvBPSSKY3LhpnXNKB0GwfmtKwI
i/LHFFcRvM5YvCLxmEm112V95YA96lm7U6zMGd6kc7yXYAzYDaPB74mJu4PY3w6e
i81V4cT1577RrT5nHgcdubaCbHJ0go+a064sNZxQzrT0XgxfHKJSqcT852SmAeTr
bOdaJET/MkyJvjdhYAY0B/xnY93RflRa//6jTQdqqo2V+H0RfSqhGZ+2dgHtDImy
GIfrW/o42gY2INL8vBTwsaT+DrmtPdaCi525pjAKt5+6Pu2qrjLKW3yby1GuaL4e
fJ1+Xi29wjyOOnWjw8yVHNWq0tV+jeDlQXPMblmooOM3j49QYQFUZtz1ettyJfyn
dvP3g7W/rthg3irsucDpDykhvjvWE+S+bZ/Ga9Hm6uXNObMRnF01/FPOQEMmRha5
nlm8hwycvzRY7AYkQSafE/jwjDZSkTYNS3oYxFelKBg0LKRKMyFa8siquq9Ck8TF
RPh7UudbiwRZfReiP4noTThI5JlLGyQC9C4Vg/tkP+TULvG4M1Yea2LcaOD/iNFQ
+NjDAkuoFYnviJH4gTEaLdmJbMdoLwU6aqbSUaayFSYbDqR798+Bi9njK9iU8Z75
Zny/L9HEoimit5jRlS3sUx21+XL5ExbP3TRVT2AvWiDP+yySnYnPDGbvcHYL3mtv
II9Tg7M7QmYJZAbQds1z+IsNZ/tmmdoj8y+srhvVu6XrCSdu7oPzhbSf1hwTd1SR
Oh5Hc09LHZIaFT7PbaY1ZY5rvbGYfzhRN7wEfeMZAG8BbpmkmxlOh7zutLtXIGC/
zxKRIvvUinm+NY9P1VFDbLAqUSsnMKsQD2y3rsN/2QXVsGWXZcabj0rimTHnzcj8
s66SJYXZ2FJ8S6bbu8RBb01pLpVwA5s1tIU3OrVm1GbYe2544FWzFZdK1DUlFWsN
4nB/l0pFryDLx7v38I9ToTk9ZF0FzQG5bhqvEqTEJ6E7RNzeWL1GSdqXvohXZQcc
a/MniSXVV9/3SaldpOuZI6PzCB4kT4EEUn/msQo5rz30hha8IO2FD3M8ICXLUhks
S8jkJD29B0+Cky1rfwLV6aHZakIYBv5Tk5QNtd4tt8K4s/Sc5MUQTkIV1aV+7Y2r
nw5JU58YSbnp8GC20/vpuBLM0XPQ4/F5VAt51+/13CByOpsu/kmfuyFmLFt63ABm
H8k32UEhQHGVF4XMdExL1o7vjThVzUyBghKM3eTVus3KccM02zXoFbuKw6ujXAR2
AKJJrQ3nlZ+Xuti7rm0PFsBtUJDYMAqRPlpPZtOnRUNJTZy4WIKC7WhcyeTYz0ny
wH/CUzbiKk2WLCDPEARRslGMAZMv/VQEJxU/u2Aagxh7z+eJVkmt9SeJiPchDxNU
Spqnqzo/OedmFs4y+dYReKkJxasIsee4Xp2pPcBvjDamMslnpQkxyGceaPJ608Xd
v736NrkEgqZMAGA5Dng5DSqur5AQOVLWeoprgE89L1XcgaIjt0bpbJfJ7RZzfM8b
dKNcCkGv6uUZ3ATMAMEd02/kb399mSTFCuMIJJ5s3QrnkZGGGSQELaVrwNayA+OI
6CWJL8D6M1RpsbOpYIHKe3/0OsIFxBluV85IjrfCn7+2pVxoky/br7T9iFXsmIlm
jcsgeUfs/XH1NMC5nEfdgv8hcmW/G41qclzzat035VWEMmgTT3XHxM6qfp43rGJb
yP0hdHacSgOWIbNFOn0tMajhsdm3SiO1XJZcpWiFsTYP+laCxUmTK1UCumockp81
HyIMH5ImPdmb/XvXvTyuxhSsROW2lOP0/2yJPzTOGI+DNBfRWhnfwVvWOncl8ngX
utKkt+rpjcvyMcH7z0tOK+2XDqC3YkvJaTtD9b8WdeB5v/mcVVlA7HbAH8ATr7Fg
WLBmy7FcZJLsY+tPs7o0mamcuEK4UlCmhp0pwx2ShPViE/AG6gj6/eiCjlItUfBr
Tnjz1veqU/Coa3gIrqdwkP0hz8tq5Jvf8mWd/05UnyX4kvcNqSwQZsk9HvQUjmAT
yOxCx4K0fIqCUdFIGaH3//piOV+UQcnJ/JW6BPxhPzfr9Y+hTl3jG7tTrMUm2kmY
qjW8CeThLl15hTcn0h1M9nyX8a0afZmV+0CR+yEAyx1e6lEhLqCQ4Z0RNQXsywBy
M7ecIkv6/EBsscG7Vu0QJKqPv1W73HdHFl2mZ/CqOAMS1aqnu7jPc679ulJkeQ8K
vR0dqp+sRWIwl1ViyCdB5nASFBszShmGAep3o9aFEl0fMGiAqy4737U2Uf3fzdhR
AIKUF10RW1U6o3ky4KIWP0TMZQXLsoE6c+7On75pixl57dUCZNLtI1uc7oHhTRfG
BEJhWNjt42DuD4JegUp90GjjeJPMAmEN4XiohEM/FVYpB/mqRYj3DqihLE0rbr/u
Pi5/v89k0+ChfZV93YefTiXcvNPOlrMl0Pnn6BtZUHpvR/e8nlkOK3+tThkdyAkg
AVyihw/Ly5elbZ5Hi/66N+NIKdAhalPkqllQaFQZrg/1qSvjKtijM+yGSxO+t671
fCciMn9JiaNLaTE7BAvJqlbcwKji5ASnTzuYoMJ73fEk1uZwHdJJfkPXYth8nHgC
c8164Z9qH335G2GKGbtyF6AfXRMRsaD8KpnKjT1SLVTExHVUBkck7KdX/0ZSXaNR
loUzhsuSPECkoLIxSSiV6v2MP0IgoRf5EoXq0TOZeMR5px9gkij8ej1v577om/D0
KJ/q2Z0+sr63ZtWKsNAUq97ofl2jo6MZDchs1d6hdH+za+bQpk0T8G+JqND2mZWl
IZw9KUy1GgyevR1hWj9F8tGCkA/qDSVSdL8i64cXYKQI3VGF6VLvwydoPVZnNYPV
9aQ/wzQlzuvjVGEugMmkj9tSyQvbvn+Igr7pV1nrvysxPKasMLjTPozncLPvSc4z
1FJkii+8DT/r1wRdd2EJmWAnO5rfhdDJ6KuOcWERTT+buEyuA5Ec7VPfLWtSNaVA
a4AwU4FFogLR7GrIjwp3IiTTqdlt56VA3UPoTBMkcwrGi8FEH+gDmWrvTo7rTeTy
cI9fGYQ8iLg+n/ucpYcCEbXC08MiknfI4m6kuh7Er15E42XmeQW8cNkQG+X5rVGR
O482D6SX92IG4h+T4ArENatVRol08ytJ4+xLCQrDM07J5rF0ZdrWydDhzrGXt7nV
2r2OSLUWf8P2jwGEp398ZpszMDWkawGg3QC1MUnbAYN/kn1TRE7uH4IQ34AosPro
7aBweV3Ay9baAdxiTzzcb6NdUzas3QqIGNVcLn7UjvLyHA2iRobK90SQRUXsgHJK
0hmXN0wdTnJbZ3ISD34WeKTATOpjJADbH8yJCJ/72X7AZrT3Ocq6jGr1NT62hiO5
8Vd3g4Ced9hubbK6Z39DHzaEJb7S960kRUJAUdRCiQqBpl5frTpVzWEQQeG6nXGz
pRYo8K6K5SNLc6OJlWqe/acA/8/K+lZT4/uK39xYlc8UcJfExze9CHle0f+t4ZHj
EPVjeDWG97T9qGSAcW+sJB2rNMI2RN/DbDznAlyqePZF6ASBWH7o/glFiMPwAO83
siC68s+cLDiFW3mqPEqQC2w0tkIbLNcTXtiRkotbZ2UAZKxf2ZHM4l+OZgghKZ71
unvGTZZZ7MrLBU6QFRx9rv3YOIHTJm3miCquOyxMaJdbNApf7BMsIQjT2a/MqLD/
ci0GJ1a+yW/rzFlZf1cHhAcWxgrZ4cPz95Ooq4ESfLTQ+5jdnFOdyk2PmCb6J55L
/E3LidFjf1sGj6H1p2oGOowTsgR3d12nwek4gxy/U885o2AYz8VBwQ5kqfnFF0j5
AiBz7s7DxtQpoQUNskB1GVl0dmSpknQctXyF3pYnRzZwzrMFwaeBQ7wdXCzCGbdt
7HBLESywN/yriLGaGTL+aX+Clr5zZtJuPcNY6BeqfoDBq+pmcPlCs98k5ztqF+ah
AhbuzY/q197kCqfj8g4sND0jieIQSq9YzlgVoMqUlgyKQspRbiXoAjyiB2jL1Jbs
oPUz6J6yxJsj0DpkbdBsa4y79Z2pyFhEr2/VoG+Ldc+nKIsUqJWWATxVzOjrG4nw
KxwRHiZAD67WSUI0t9rnsl9FNR31XT20lD/7aywKLeRuCQ4+R7uOmJubLohzanKQ
mzhF3H/DL4UOdkhbhL13l1DtU4ddep8/Ry0opQQVfSKqpX4gjLKEuietPotSaARF
J15Qy5tD947s6XoC6DK2Cs4NvsyFI60CcMjm4jJSnvMjlK1SKBFU2Vff5aHoMQqx
xVH2KRATPv0gckyyJpRaSG5hVLT4catWbXd1RUUHxwLMFp8S39qkKOhIcJXknwIM
xDm6O5cUW+30F9PnC189bHxXbDo+FNYRUMqxUYMkdGMgnTWcFAZEqjY2UKaFPiVQ
WkBOw08L8KyEf2bFCLYAlrxHbQiHzTivV6CvhUh5CQh0KDV8bScfONvoZLjCvSQK
E/xxT/tuuwwWViJmvZI6DMaUsTRvFGukXvZ7SLIldELDrI2Q8TOcFEJkT0vF+h8Y
Q2cVN2k+SV7SwGmrnyRuReCqa+yTOa4IbcYuJkpyJW6I+C/s7IJgyX6HMuQaWTr6
UXUWos4nQm5Z4Trh7T3OKeT6QgmElLuT+0mOwC1/VECLLXSbR7Ddj2GJkT2vRHTf
K9i1d81siRrtVmJOQr3q0II8JTiERoSWneQn6zuPuTr4AOqEKuX85alio7hUwgnI
cidBwLo6M+J1gCOXkQ+7J+sAKb0+9y1zg9rvlJEGMitNyiurR4hZ/+wWwj7GPZnC
E8e09FyFJAiMPYW6NVx/e8AIObo6IYmC8hyzoJsYe2gwQkQuQTDJNXBohVKtAXhA
wlyOZh+slVmRwT3tOYo7Gi0HozD8uv0PebwiX5bsLz1dpsuoOBXyXx7JsL7/o0TZ
cOPRCSGT8wl+AVtc/9MWDEhzDA9zt/UF4XKtxSkb0LjqPxRL9xHkOSfB/pSWfsTY
Gmzk2tFn4cGqcqncAo9A8FvqSmsSpoGJn08zIF8JPBqCEimaRG0UXxwevCTYOL3J
Oa/JCU0hWiT477tn+XNA3YqJ/CyjbraC7DRmu9lgLCrhhOvfO9vnzIw1sPyOFXC+
awSp6MHxeHYY4mHqq8kC0qfotI4UZBHAkrOxez2iTqQRyo86VwCThkkSp+yFGvKe
rnVhiAgm+da0KHlNVMeSR1fWJYwUeKJIhYuF4H0N2k7rLWu+OwkXmeNpT36uA6hX
GCzvI0WRjgXC1E5JDt7znp8OWK0rldKp9p6wHD/1hPzqGhp3okM+kH8KkWlfKlil
LvfvJMm2xe/+BqRpCvuRiHHec4mNMnHeuoeTZSAWpE3fSaDs/FPJAJxWEYiMv459
MF+ThFpwAjBHol5RgPDWxKKXBqYh9uqhorPPFp/mnKd00P3kjRY7Mb2UG24wW3Qu
hyVjWg/b3nJj/DG78w5iuMibK9L1he1BJ4pNaF375SquMF34IREN0f70nH9ywZe2
WYYRsAzv/E4j36TZlQsHhfO2pwxYvbvt8gxGTrM9X3saTEPbtyDgX5gWJHnsRbpc
Tf8qwLhTI8PofEhVJWN5mmVXWkr7F+tvPku8wh3eV8fewKJ4d7RH7FCvQAfQlk4F
5XKjDNkijrIA68N/BuZzfdQzAdRe0yw+gU1VNKWQOpoVMdYONSRz/ZZkae3zM3UB
SjHFHX8xXKO6py2cCYA/g2NB9e9ZMwd6dLNMtEiJzdCRlG+sWr82dUoL+Egh0Q4o
99yyHKdBNsadTAgrUfDGitd7gKIoWYidqCvvZgEunRM18TOLP5g7Ss2hX4HvZ8MH
9Qi96122mu8tOBg1ewlj4PClbG9z66oF7nKiEDCV1kg33i1XIUJbNy09Jh2NHV66
W/LI581bNmDthS6fjJ6s0BB5Ori9MdeKFNKEyjOI+V6hUaNycS67OhwtvyDi1TIM
vbICqEUJt03vTDUB8kHavFaTZQHzRhOc5OWC58kSOGSxnKRFX6uKO2H8WCLc7v/C
zyO4Jxk32mmm9NR2lELtr8H4YK/zkxzZ3Lc2ULXoms5ZodIsgCXKsxDXYXQ/ZZ2m
CP3L761s51PVFHMHgaec9FRLkmPjJPkCKjsgwZLVVeCQAovdJ9C1Hwz5h81E7Edu
w+h/gba5xnO4MUqnojbibP/MPJuimmfE3pAWHEOutHMUu0eO+9MRGcgxR38jygNH
7IveaUAOyABMvki0DJrdAYO9M+Z+SABLOTrtMozY2vxuMoNQX7wztH7JAA+ORSQa
w4ht5UniOXlS7lSqi3oyDmlhaSRKpR9QGs1x5TciCBubEBgU1BlcPgUAtWQRRlC8
lePVRKVmAl2OPvBnf8EgH7wry9hQjTgGFFKsl7bUykTlSNSd42RrInavMlihL+wF
d3V3Y1bPcbCzNYO991OnvbENVUS87obQmlnR6hVtrNvXSamfvcdOUHCf3kBcBWcP
LGnmFZ46yQXe8iNLd9r719FuOH0MaYeYrmHFLFuySCTA5iJntsZKZpBdkLD4FwKT
JSumkjB1lGrGRP1DZAQ4mVp0lvO/wBZrUUN7XduV7/CPMZUVF2qVMiiZQqZKXQJ+
U1Hu+047gRooaG1qwIKVq9NAWG16m5ouSjgeNGtuSS5kV3gOXwBKnwUkgojjA8dK
uimQaPlA6NapdedUBe52JaNGmKTV46LgGQwVkUTMfsN5ake5FhglVtSyz3OkVbKb
YLsXOBpBxEufTqu/2x73kOee8T+PNs3hSHhnFgrlsfs40zfOyL2o7I330dI4d/BI
a/FWiJ7ukpM8RMtbWRNgj+gTRkmi8YpyGVFy+ajuiyMCWc3NhxnhfQUH4Pj2V1gc
nfy3OfUFmPYITRWLmVHnkdysqdR8IwiDJIgjMBaj4SX5zqhSgc7cUWDpg5cZV4PK
u2zdhyHIH+X5ZGJLjv2mF37WwdLIwAtqBYNZnjjuIAomBxuSS8X5PESoSdjL1oD3
yu4sx5DFdaXMl7ElqbHOxwn9adROaGNC+KDKVdtjL2RXfKcP4wNMxxPuNun5BscF
bRcDKQA2vBUY94kbrysAzLYj0pYmpI6yFK3xaRKKbGfMpJW+9Qfx4BibEA8j/2VG
IoaoN6AsvQSwH71dKciCPQH3AJ2MQZRCldbMqBiSBJRCudj5mWMjV4eMA+Hi1WPM
OVOvNVtz8f71Hgl+VhexaWOuVTTCU+Ns31aVRIUY2peLJfxZJnWiGo+YReDw8gmo
emizUxC5RfFpZjbjRLkvs/Wjd0VNrbazFaFXdRqX7HXD8DYDVwuqu1tc2J1CYZsH
yrpBooKV7qm62j8snl3ULN7rw9XJcPuyL5rWJ/h/PU7G+KrXYKeJ8E3soWaoQzH6
cN2tOihUbMxUNjC8yCrcj1KOMX41ejrpzTf9lkSmxN1NIKxiGanma/G1KYkZrHO3
++EDFC1SRiddNQJLfx5fizgmNnZy15pcchY+oY9RYsTxb2tu2UyEYHRiokolpR1S
Hg6vUwMU32VAaikbHIrITcUtu3h8uWcRC9dOIwOP8cuwQzbBQ7u0ujr5EjZTcxTn
Do9SRVTBjQt8S2sJu8rH89Z2X9bKIlcYf0KwF9MYoa00ah+ffDnHYKRtdWOIfycf
5Y5tioQU9Whx+kEb85VU6+3O59hh0XaWngQyeFU+b6AhGfz1nDSIY6ZRpPKg5CaH
fKPRAobLUHzYR/AF3J6rM+8uguI6b2k1kDKPJppUjsyflGVej6GYLUwWApDVsevf
iduwRF1uqt23rgGG8ejhIT4lGwZg20QRvnbXofJ6H1YZ2eC1c1GrvLzrqpIFf+W5
Y1k8mp6RlfejLHacb+Fli/NFV5pffDPIZQ+Oz8sKveYPjN2aj/wFf35ESX+BmGlc
kqmVW0rq2HVpqsvo6OeQDstzzlLg0N+JgAbPDlUeM4wthRxchdAmgrY+hhYZwSAJ
SFzIeE//jk4Yu4bA0wwrblMr8cisEkMSp0bVlorbOOaKfBk8o6uBJQ/KZpMrQ4Qk
BgV3NoErI2/RL+NeRJrQQFXeDjLGF656Gv0lG7mTc/Dk0BbtpHCafuvp2mi+zl/u
iJLpwIOBFsK52Rsh7GM5bKiPdOepw9Ykkcl8JhqkEKwIAjl9l+rL79xTw9oASX0Y
U0867H0Vkg0FkoBUda9ENtMobzMOyYV7nTLq3+ujzvqnaPdymv9RbkmipIKRNbWo
ANkUFs+q2nrQOExlK+ZpHdwl1s5dVsV2Jx2zrecj4adFiYwRgMOCfo3hlEbYC+es
XcyKo9HhNMGNdagPvjA3NkyAmOdsX+RbQR9lh6dbBVoeV33Qqc8CJZC9a+ox18MA
SEOqkQLu+rjC4/eFJEx+bTg8S4Kr2l3ShcZLUPmpW9XrRQj012bePYhcyI5aKXkl
rVpl3HQx323/d4+cPcfruFjmcjNkVU4n264nA6wRBsEqGRtFSZZPNZ3I2l8A6Y7l
NHlVM2WCt/5rCfym2uBjQ15B4/TMVYk7arxAthhKXs5q4j4COxZxI6JU0s9n0lCV
whv/p1Y7MD39N+EDDB9mvOOuaoZ0ho1+gJ8EPExVGm0FiF0elkRZZfh1rKKSY3dM
9Xbzzx47dbFbV3N6IfpusiJ7eJzQDXoP+BZNBT2Z3DbbwYwKzFTTNvXNcM4ZQKV1
0j8VFzY9RmW8iOmsfDnjz7aOOSe7qxzPOfm1i/iTLOipWTzKu0IPQgzMTVebJPoh
ftcIvPA9mwTFR8u0VVtrlv3eqNXMnTHaMM6WPDMSlxmp2/0nwfCCkGcgBy0lAv51
LvdriZWF44gNJRFVB/ALBZppmKl73C+eS1LEwwmqPB+F3Loucu9AohOxGbXzX16w
rta6X4Xetr3JoYDoLhNszIfdY6nPkr59Q97opATXi6Op1jVGnvGuvzBqWM/lUw3j
ihMnwTxYC1rNu2iaQoG8qe56SO+8/2iVNpsG/Pl/6xWFwRcb5SN6Qxv740U07V8t
yJJd/tnmwvMVFBd0CzobKWgK7ZOnUxfzy2HJ459vj54WBM8d2X+rg3YKb/Nh0eBI
F1jE9mGlXkstbPsB3FrA1gaIcgEFPe+k58BC2NcAqbvDFKCd8v4MBUZLSvx6xFz1
dCuA6luXJHkAIXy7DS0CHtTgLMghiyxWVgV3dJ1FD1mOlJTOyCao1Z/3skxHlLFq
Y6oMCD4YWV1bpSoSxwq+H0pQZBwLWQAeCxcxarGDKwFNzdjOuW+MvNCMRoBsjbIb
/4XRZsZiz/65OBe+UArNQrOjbDkuWGpm6sUdpjv05+st/+5JcWD7DkafVXdvuedL
teJjBmdug1NbKMOAILMParQ4OMzuPxD/YfltJKGyvLHPfb0xiDkw6FFGMlMLPr+K
kzjTqNPFAj6RZzzt5vS3t5iYUiriNRiPQnjYhTQaBwq62h1pjRGKqQt4h8xM2Y0q
jmS7px8APVLO8wNj4Mpqkzep44eL7tx8HoJx1P7zGfJSnppEuo7uKOGBBtrH/2m7
mkAKuwlYHnbooSx0/mrLjT7gX79vxDE+nrb0JPWlMyX9Amh4ByLKk6B4nROoMPAL
1exTwWHvL4oM1wMfvWAVRnYDPNMwkEk73vz05Yhkl3kek+1HHLe4J/aPjcI8NHKU
DzlWf+eAsO16zPafqi5E+XuO2bR5gfodPMg8NjDX12SbsblrRRwBuj/eBBP4p6KP
6Yu7lswtPq5+woZRw86GBQp9dq2ekdJlqdAzVwK2nhW/jFuKDErfUCZLQ/zb5pOl
IcDgivIEdF3tWu1+c5Lcj6JSuJdb5NCRq83WRD4Q1KqILysk071uhzObQ7wUr90/
Omd1TLNxSMgF9bldPv45To2iuA376PXCMui7TbuEwS1z4Ipbr0a06qMy4R4ZtlOb
0HX/hZ15ky2u2Keue/NTfXQ5qNWcuPxPig6jKkxJlg0skfafPgu9HPrRcQ5Y1Jzz
rdptFAu4t1dmd8h0FNkI3wzjFNmNu/aUjGFAsvMRT/reE8iR9jNOb5jP9jbLlyr6
9fBs/9aBDTw0r5RDzArRZnNT5LGb0iV1wdwl/XJSlwGotf3QD7pEu0gCvZ/YqcDE
sZqYeSMReBj8DJWEfW/g3B5/3R1JrBzjieJAZrL0Yoep8CUcYwvM0uEBQJF4eQiH
z/kz+V5JlJ1lk2wRp7RvOWTujnrPRljVS7gqq8D4CpZQzX509G8YzWaF1GRy9MU9
JHLwlsSNO+Sr+m1v1rsFPIQQMX1CIN/0nxy6crXUP7Vygb9OzbtEds2pyAvrflch
zB4dyj0lJ3ld3FsSmHmR9/Vb4frB0CZpquIYaOkx8tyCMCYnMjFP6+bTEFUXtY0X
TSfljwSHh0mPofDRgI0o6z3TFdfBqPBlyK2yxhd8ztTUHHN/7G0QN3bpPMGoZ83y
x7kMs0c2s0e/n4Pb/nXr91lmB3W7CBeCxP9BXhDZG8BI8+sAoWnzf8rIf+xzDUBq
GWqd3FW3AE8Il1vlTvz3UccPPwS3lJMseocylcOWACcxaEz2ZpezjAjfaPfA0k7T
wYzBP7r6Y19lfGmuv0pGSrZbr0QNWCmwqOJ16aIeNLIwCeJaDnSL5wihTsiEgXs3
qX7wiMKKSTK5kdjrnxhZKulXAuEncpj1TKmDC5UjuRbRhbvNO6HyXV1X8Lo/FeAU
uftBOWeb90vyFGGXQEs/Xi+pj1CwKh4LlrU/mvKYsP8UJbbSNy8owkzByY1QCSOB
usbxmfSVlzSuSBXtKh1BSdOWGOrmnKboH1AucACktQJ/HzApNysOvCjf4k++7vMa
fisb71gCvxe9zEHjk1N0s+RlVKlYh5lrM0V6l0Eh3SfveF1lyUbWgtWArS8/K7w4
XvVkMA7nYfOE1NiwxX3yHEaBsUxADoh0wNjlCqPQMFpElcYkY4sU/2RQ+pDrgeMX
4lATZidqGx+NZGpIS5eXzEqfQFhIIEIXK5TYFMBfgEuv7ZJ/ycrF6uRg+NbPhkRE
onCtSsoa4zMaBtRE8VSu7PeIpz6k4N1szVmbh+SGEtSwL/iGImocx4xNsgvuPxOw
ubPsLCKvFsTz3l+sCb56v+eewlPFAq5eDUDYtYn06IWK3Kkf4VI/WgMb7SdROtRW
MQHlvDs4Cn2bXdjkdtVbf6AV+FZD88K+k9bpkV4E3a8RTCyA7pAXBT6in06DKFCA
wiZz9ITlM87NlnLOjfATPTVWcp+0gEhF0mdl4gB+Vh3QZrUIBZkWeQ62FFmCyjKy
hbYDSawHde08NXBCs6PWSS1aWrDNj8mcqoQsscdePQ01dEyukhAAuqUGpRN5+4Yh
ZgkKJUL8hQfc5rgijyrmTkzlUKoSsMuhirU5OIU6bNeWECRvMsb3Mpfqq0dRmp1d
KOPwXVG5h5KiqulD/GvDBxqjEaiYp4P3wVrUgO3Co4xSqcNl6H/HsAOJswJHuYmh
aspQ+W49ktBA5rYloAcZTtTeev2U8JJ9FJO9H4cP3BQNNFhCXgvd/OD39JPQQGG/
wxLvWY6fTob8UnkXLYa+LotdOAmacNUq6xG6Je2Ak9jwBAylaxiublMWPGAr2XCY
RhgXAAxX6j/G4DrYtb4AXb+FwdvZzYvb+LwZQq9a8j0ePb0GzgcMRkrQLfh4yBvL
3TQXTEgPDhSIsM+gzsMpKPdzaQGCI09GvRNSMqlGHy2/3IHYRbxwr5SgKj7QeNsq
rtRgqH24XuuGS9ojTPWFJtr6IBf0edHWIEotLTo1JHUcSZYVndhN28ngJMY/mDJM
bMQ4pybpknBy+TE3vWeCDmULe38WbROEgnHJOLbXxuvgfbArGS+PQszSrRu6Rm7+
okelsplBf4ItpY+in6r4GhNjWIpfSbnuIS5uFHs/k2ZTR/IkWYphk2N5jJlWYP5x
Lq9U9ElEQqgIFrfVHyX27Ue+vWpwKGgNU3wjccrdOYotWmlch+HpZI7If/CczaTe
0uhCeKO93uebPWbCmGTEhZnXp6Q9bDV20d67SzK8JjHgbTlG432hxYvfWpYDe589
TRBtkfGUleZ4YQK2gfwNDIhLw5qrckvdDcXhsZDO329FfjMasCyBYlwCUT3zo/pm
mJa8aMnjNBcX9mfrc+rFX+rgn9YVSBhWLt0CbWuKnIWuGcxW5uDzZLuwjUVI9k5Y
0mTFIpEJFI38xs2vN9Ao2Kd+YJDHX4nIrH4UQoevSDboIp6LaJ3kGLkJunfGV+IL
zA9U12wB1HgAqZLk1bl3fkMZzIwqq4pfJ95kH4FIFyj/nAeQkE7kpMybs06caLfx
835U1bkMbQhXFv2SzjJhRyLP5RBH79zJFsNiWxS0+e2b0T4FM3Ox0IydkKhSVQGl
Q9yR58E9JRsl/9QKauJo5WcbDm+W2uOporzgwfEQavfFGj9xzv0Ji6xlaeMDrNux
fYPbFfMVBNh6vKziBdS0vQ4b18MNpZXavfL5L3fkE61zaC7cSk1ebjkVd97gZxrn
eFpldvtn58KgGc5nm+YVxZF/y7C2YUk4Mof3wTgdBD0WH83DTpT+wV8lsPhkGM7B
10kLa1EiBJVLmZxrrUAB44U7zfIvdsAEUbOZA/aD5RwpnpUA++Q8V09VTH2dJa/l
vvdS/hVfgl6k0Q10WfIaOqFhwFO5bjiU06FgFJ3VTHoMrYWH8YIcAEynKP/9LkET
A2M8PSRFkvRLjH5Ku27Q7TGqSVnHuVR/i0Zsf/QNGELr5mjbZYO+YUHRlYBFBwIC
nZCK1vLrczjWNVyBx7AOTFMfaWIq6vCuINeR57VKUtvdWOIh9UKqA4urSRc9YNUy
IGJviVNIv0e0DxOdq7Q549fzV4PkMIdx4ISnMsxo0vUSh6LY1J1HcgEe94eJsH1o
RfmRKXAmtSHU/g7TTe45ym9UXjszazEYxOsYJ0yaa747j5oYa6cg6VYwAlUfjyJl
CIfovAFVzRs/3bIP3Rkn/9RDX7dABjeddu4gy/dloxhI4CeY/6tnp+uuOLEVUcr3
MVsIREb2jv59wQnwt4Xm4DERj6TDO9n35QUQ6fDCfZlLzohcGOUYUKO8oou/rEgF
ToUqJGNZ8lh9BKQFYIxEOBpzrJyToNKet2GD+UdggphzeglzNhrBRFpqzepS5cIr
bdaLBOKhiGZ+uCbKXu6AoaNW/caOh+/3qMFo7r9+ijeMP1hH8frU3OKPuHu/PKN1
CyM6jH60lBhOjK9gupHyWX8C8S4uuiRTCcUn57J+mRJo5qLLBRWh0AOWN58OkiYY
XLg+cq2DBl/zDPtcPf7gBbHipZqpGDtP46ZhWmN33kXXPkfmun/jV/kYNW57sleG
7lQ5789Zz/UUSpSbatNJ9r2VsYxkFKpO4fjgyPnOA0vxN4Sca4wj5tB6i4krCaKK
TpfR3LUK1rRSaMLdEvNzEx/WWRqX3m17cQ61g2wCmpnquWiBXqkxYxHhfGxnWEVB
BqrXay11uNFAEqYIeb8F5y7cR4K3kfTXOzhdK+1rV5LI5tfgQxdkcClsepxyrmnP
bI2qS4X5xXhsR2SJ5+rCX9NhRfDcw+Sqfap0uRW/D+IQo84xup1wypxrwl3JchsP
7dw5uXFJMoUGL65MKWx+TtBD9tzYJt2FuVWiEkFQjfEGlTNCvovZrHd3ttcWo/9M
NLpEOomvUiGQUz892DeErTdo+NwldYYxUTNfWGIkJyONHzCWq5M21iC9roqNhmSJ
YJdLPc28op+9cEAIrbWFnSSH6b5fihCXhNL704XcPCq+WXpjZaXGbPMcNkPdubXT
uJf5BcS2eNWgopq1Rt7OGhbxdS8NOYENtGQorf4vhipX9FoTajH7xBquMsZM4asZ
C+8/jeLcguiqLc9Lk08coRg03k4uUR5VcUI9GIgFqJ96/My4srHcJAvMSvYHiqB5
Ppea/OlYZknR354yvpFYjVuUUKGgZ01f9r36nKkSp1wV1PMBJzaGz9Z8iTNA18a6
ppbXLcH+etUk5ZBjDiAXt1eOCd31F+u7itZ9PUXnxyZWCAYFSemZMmEjGhWuNIDH
AbJhz5IlSFs51iju4asEZYFWIQf+u88MSCbVjFisBZ596MAdq+nnaepisTp+yuTx
hK7wMskSeKv2OsKri6ur9vo/dMxps6PcTqP/k94S9XfplrIQ1R+hVs6RwRil7igd
+hZu2OtrIsun146qyj1OS5zwOrQW9/aBLXWK0+E7cdXg7Ex80/jKbZ13GNba1i/A
gECe0CUDwgjleNcCndcLP9wJ72tyBsm028SFumXbfR4q1cs/dumHImmCLCH+VlZW
AHUnQHb+L5/dHYXa37mW8C8BEfs5D/cy0OZDHYVNGxWzO1dUuxt63mG44b9zkqpo
qgDwath3J6R1zhF/rJfvBUaHCSlakMHqMEuYC7wUKOAJZlQqxtTQ2vgJmRzwNidZ
sVpe1zS+DtAVyM4cmGeeFm8g4wxfY3CPQ5PtJAIhi/LQ1X6QCdOJg1XopseNT9IY
Q9YJXv+KmuL7T81csgXMK+TpZ6yxSXMxHZK4g833PT/qQHMLWvlA1uwzLuR0zNIN
2IEHg8kbRY0TRjl2I4VPk+5b4CNAZ/d2lNSfj2MlIK4C4dscfI2PhwTBDKHqeJE9
3y0rzCd9VbiW0isjIZzDByZtAsvtuKFGaL4lqPfRCu/5ED3qjWlwgjjL3j2xjGrB
XrX01owi+hw2YYXNs55eERGyp5HCM1vEjaHt9OPGxncHvqfQ+bWO4/j35IvrOZjR
HUuIAs4gDXkmWUy5VOPDEpDI8kfZglcxgQf4wz/4+EOf0+aFEMof8TM6uqDmFLeP
FZbe0Lo8hO90zTH0VUDCAxhUwC+uqfhx9BFjigfJbyT+dFpvgcA2QE81QqmnBcV9
lIjdPTVY+3fRV0mRqOzUOUuBOAQWKQ+Zj909uuwr65pKDBEFgLfZM5mGoT4/Hpj4
nLH110g1cfe7HaJG098yUfKHqKBcNdfkKfpQwGnByqE1ehKX6NyujbvxiCRMCu4b
24VN+qwrIXmJRqF/4gUTdtRLH+pSzOXTY0DRI8XLC47vBB1n3R+lQpbqj4qyd8tv
jkAF1CQawwAkiyIfLsXENPEDzaiHLV9wjnbNzsNbfckE8H2YhO9Ks1IrfrgmZP0G
54cchkRg6dYRA37BNiM0baJK494qOdO64mVXOTSbo2ZoSkUTAFj85hNLqeG0p3a9
hs+WIbye+rnCkPvF3libxEiALdpQ62B8v629qyymQKIxhNqQmlvuVkTKaTtEqgLw
SqMfJ9Lb0z9GblifU5V16p/eijPR5+LIiAlrNH789qIVvwsrBq3yzZhdKc9jVrjN
t/gjnkb29bgX/9K8qS5TReCyqiy0FK802+Y+QHAp38XaiESo1LJGzx4iMYPFghwi
+WrwRI7gNeB8e+C1oQK+p9nbO8qnbZyZE3I5jzPrhpL2TWiySuAdUT9+1IGyw6Cz
iS2O/YuzcMKLS2UyzAi5DuHxtkRucAPvrlRGuAfiHSkee+AHEa0ocIhYrE6fMOhg
ruSflT/tQUWM4Ep9T6lz1U84haiZma+13SnrqBY3Ywpw3iTKhfB56DqCDJA3Aga0
hWyCXvLJw7McEDynCyk3lz1kK3w5+zBmNJZDOZZdYKDcBoeCYRRI7h5W14w+36MM
fHktXyN3G/0JfvZ1vbriEVnMFqouRbN7ej4hdOv0aB2QZsBLOONJko9QkoA4pSWZ
QybZj73s1sgvnYIfHPP0Ir9uZJuNAG+Wq6SRBYuNWQX0pUAhqPDEbgf4pDIA7SZb
hBrEwB+ZkGiTu0LERapdScyl4rGgFZ9FWn60pWr5Y4LzDqyHPjVeF4M06cyqSJl5
UFNrPgCnCj4aCoAwkUwFzoTmHChR2+HDQLYKqVYhxUTLKFojv6ar/18AUHaPXjFf
HizwQdLBjK3FtVjDN1eO7959SfuZ4dFPzcHL63OR+qKikj32y00VdgixmIevG1mS
Bqv62W7Cn78oFzIYKRcyO+LwM9tqGg2YRQ9PSuExx4DguGtclMhAtbLBQjOk/oKv
Z9wMwGGETRq9NDTTkkA7eKbdCp+0dbEh7BbEgSBYBtgTP1zLwOwXBbC0DyKoW0nx
EM7qwlh5Cbp7DtWB+AI4ItTmVvc7sGZUyFipevFQA2124fjD3qQ1cNTtwxetmyWC
ZqRt0aERkbpHPmLwwvyhhg6EYWw9t/gHgh7zGxYERvzfaHt9Q8qg8UPU3jeHiV+7
k+iYY+8wmh8i4CrFgvKkTzCHOrki5RQj+VtkmjHTgWyMGDIxeR4yQ+BFcy75e8nm
XuvWbzi0C5xI3wUJwpXdjbc6ZuyMXl2jljJwKfOx2EOz3rieVDY16L6mHsjOoDJp
GFAM0eZh1A00wd3GTE9A7J6utikZFua1wfXq6iOu8g80plRW6paZPAXHgwbMN3Ki
MOvIZNCU3CJ4svTk5A/Gpa0FiWIkESuegT9O6Gw2Y5/2Vg9yTwoyhEu0OoAOT+l3
f3IQf2iF2W8MZlGVprPLGadPWABaLQJWQIFyKOoQ6NDBeKzs7GfK6nWwFlGgNUD0
6/cciWOCzxKkfXiPcjIkRm2A6qu0Cqqlg7QjsI5D+R/Yri718kiJTGtz3IOlK6Kt
QxJeQ8yahRWbm3BnIG1RNP8Q4/xmUKHtzn+VPDNXetvXQ1YTA/ZgeKjtRzftHREo
Inp0m11E+ON4ZTY9T6mNeT4eM/kQOV/qTItefRbQwr7ZGCh99TobagN5o7AYI+G1
+3huhKy8Cudlri+ESXiHeN7/K06/ClNCRjdZnKg0kjqIot7ZxiJ5xTCrkbbKhs3G
Csqcaws5RSfJ1t/gKbTiWap5gq62wrDgS0Mt6MuITN4GgWHanZPpv+yBp1IfrELs
91h3tDlT2TQ0iYKclU4ZvGvgK6CE1P0NXMKzhKOLBkXV5NA+d5se7xZbPXcdFZYC
rgROzFDSABkTuwdLBIlKspM5qs3AVIYyxOh49fqhx6NQ5hrzTenfd/DzQCaiFlQP
N30ZUydyMSMh5hthQrRObgeD4zOHss3GNyKT+kOC1qBH0ORaHr7rU2YsOV5BGIyW
mrjQD/ppEybLayfU+Z9BSWP8hkD29iQKNxqfdvYKs9ynla41Tzcna8nPSgo1HHd0
uTOeTZP/8hcf29YHDfNzRu7fXyzkXNY0UxpFjJZHetovy02nZRZnbdXyV5VyLfzf
8612FP3KfCL/2hOl0oY1GdH9wMPFk65feqX2Cal9Bzmq45RsOQTsR+LFQ6zXmSL5
2WBKOyLzYqN2RgOTqwN97QUJqu6tsOcLIYkNJmwT7ahZBQEsnCy0akx0LNJdkvkz
Fa9LLW5I3dLJIKnQ3wMqEMh5n7bX30asjjN7IB7U9GIIuCV3tz4AGzpdhcfMryWk
Sz6npsNxxjtsbcwj6zWVljTX+LqmccR9Zj+3DeyYzw3eJeL1uxXwZfC6bWKZ6SM2
pCkfz1GuD1xOHfrRZM7Uohx/40RFmaIPWGuiRgrcFtkdzuBVqNAmCKSVOrdWszXO
oPaIpbLd1b+uJiAvpf6brzlbh6e3+nFLs9PYNn90OsBpY8I4kAExOyK3Ss6rFiLt
gnrxQgqY0HOlL64oNH6/qFgv/liOkReE0VZj7uScO8qAWBdp/bag2YmOr2sW4SNI
sN+2pqG1lxz5hCskKOMKeGkEx2em0ij8EdMo/Hmw+OVyWjwfmyDgaWqx88AY9qEl
LAI5u0yxokl+sQMkb1zvgSzVY9vE2muoOgdolA2A3ibEj1k9UC69roFuDxU6ehAq
X9XIWSfKCm25OX/qElIov7rw7NyCZbL1q+cePAAIBC2hrQT2l1msN7iQwFIswgRD
nchKX4OosiXtZyeY/Sf9YsjcH4huy//hmbkVLuoxMME/E9ZYEwXQfDrv8tuAwzlq
mUduF1Zi6XKZTteSy4n7/mZo+PVS4CgeLbkMuO3ProtaIgD+u/qo7Ec7aty71XVc
qXIzS8tWZXijFfbQ1ZH+gDydmQ7NXABCifhtKmMxGSbqCCMdCkv9jgAkx7shMEmR
efUVDByuFp/jEvd5hYT2DhcmFRTvY0AuUHCrvLV5FJPnKKJxw1aXpHth9JDu5ErE
HVBfvGbRNp9pmyiOkhQBW+BTS+qGKrM04HkxePEJMrvtYFgpl1QAnvdPfm05DYk0
5SWCFR6LOEGtXoc1VxbzAFX4GE8GMyR8q18fBN8A+oR+wHfkCV4lAbjxeTYD49bU
Eh2US58NkAozkwjiPdZyIfxaXSrHmVNKhfZontAAYSF7faCPlbkdfk39YoTBEEvJ
W+exNgiJRSdxL+znk7PjrqK7FHEnF/ev6jIIk0ET47PBKUtexIzVSI8UOFzkr0D+
Dd7KZB4lx+6s3zFDuvZjXihq0LwijlLiOaTJqGTA0ZGVvjRV2aJH++GorzjOx2HO
vMd5Qk62Q/srUkmBByPhBX3omWfzHX7EwLtSezykNeDfCi593SzTPnoyfCqX0rVL
jzU2g3QQfDr+cuEbw52UnGLwIgR8IJFqik9kbAd5hG4BWq4sn5XDTygWm1sQ6CuR
GhT6Vlef5XyGWVkQmFuUgF2QSPwEV4zOe2LD5KaqwWArnVV+jIk3tHJW7I/oyBOK
5odc6P9KNCMgo54fmr+cvmxVfSVWc9eIqZRpHg8G0lkrMjv3FLMdpINYsY/3OYyS
wZLPD/dUppbOeJAz0JOOp2DgeEfsiOIgcCaCEkeRMKSHKlIi/esWe5dF7maHc8yS
cNa7Zjl3CIbCWIHalVexa/pSh4SF592AakbbZqtdFVkc5uLquKeaSULMOS04Ud3V
D8XLZ6HFhNxqgLE7CzLUx2hYHgGhum+DEP7+XBbeSj0Z4TxDvkPzWTVQ3QZCTRR1
OaYD5rk9cY4e4lPBTl23dYRFjHQh7IdlJdKrHlpHOhz+9Y0Ee3+O0buxZWI8lMGA
Fn6tcvaW9zURv7w5Aj1Bd1pZGjjGb1JUQCL+j5CJ+rJ2HaCH6hn0LWUQhDl+/IFS
Z6Yv2Zja50mKvTrUH3AnvQcKlGF/POqY6j3DnyRWe0lKrSqW+3UsW3On8VXfl9IA
pXjqg0fIecPu66iYhGf8+8OTlNozI/lr+LOsioCUUoWfX7Z6KlP1YBzT6V7VvguA
e21KN34gdwi8iB1QCmQSEIuvOi3LEdqq5YbU1X8IWebICdp5Qu/1Ptq4MR00Gl48
JLfyLn5yuJbSZPQlujZuRS6YdFxnmKcumap9bcgPxAvomJkwqw8tISh1vBkm/y2Q
ndm83WD6MqXyFrF68xUkRRvqRBQ/PxLAsp7646xIOllLPvglNUdDHi1x6Tth914M
5mZs9mhB0BRBLfs3aL7c0UTcFw7j38UXNqPUoSFkqU1yyv02xCdW4Ie8KGJQgNBI
hXc315BzBNEnp621w3du6f6acxkKaDvxnMIo7gI1NQjZCdOgfYvjrrFBYkSDxzbK
GxOSrBZKO27M5526A2fnx9pxFrVXGzXiHsCuppvipk0/5IBq53x6zBEGjupoE4kS
dkMOvQop3AyTMPS+RDvmq7L0oR6Lw00FoOmfdQparsdxKUQWAex1tMYwlVPBkSeG
pwGwxMAUtkcrk/xDCVHgR6qeyZaOYovNyJArWdpv1AuTn+Tn2Eco3hwR/sH8Fj+E
zlZAD4BXqH2VdHkC/WaIoc8327w7nrtLJvn0GhJ9S1n56qR0b3VSdijHylRyYboS
dIdYE/b661aZp/Pr1w3sTKSpBdFiyBmoxhaGMJTBp15bZUS74SOXDOqUdEQEH7l2
IFNXdV9u9v9iGfyn8sPdRpzHRg3o0rgMpP7sjkGYSegs7Q2NTkTDVjPJji8UEl+R
FDqW1DjxiWyjYnKG90iexNaqdFOjP4k2C0z7qEsZGtvxhHtilOMZE9jPc3rEfkWo
5UXDjH8nEiLCcLQuczHpT/KKEDV06IuR3SFOvVtB5DRjecKQ+Da23JpBJQL0d8gJ
OLdUDZuHGmbfrTmmUWDCaUM0SMD0A3idM9cmGvjcYrELA601X/FluCAzYUVKj1Vh
ZwVMBqI1WNlQNPaRJhjG3UwbyuEAzjUSY1OIU4uELgVcWPqlt3ZEpdEXSVGlbAMR
IrgpNU9HqLvE8naY9xCODQrHhku5RP5bnJwbsdgtf99q2y2bbwx9QSL+87EcZOEf
ljbhYL9GU60eeFgSOj1G+Go6d51AGGDP/S4x9XUSt3piHU1dgdvcPhAE52v+IlvX
6BGvlg47UHAqr6+i6/aDLN6+gLpY5p920QnIEc5V/g6ZST1qw8wpWq/DEwHxs+WO
vZqrr3b9x1H2D+g6B+2toP9Hqioe9X3uQA/VJEdG3A/AoDcyda2Z94CjPQvvAYns
nAiKsepfykgYZv1PT8JWbjBW/Lw/XhP+BVd78NYA7SROYraIKkImW1KTTJnKFYd9
LOqrwuYv3q48uxvXBc67ipA6aZC2GEugTJPCHeXqvxcr56cegSypvmE0PQXaEtIT
dOGDgMnHsk+Ssywh810f+Ct1mamTTWlseNEFZCfvUW59Qz+9svT4EyTrBM9z1pcH
gfeWC+isVdzAv7wEMPfDBO8Z2dti1eCBQzlty6oFG0XWVz64PyoYoLbols4sXtZn
IOqZYIQv4cVzHH6A/SVez94sHnCHhzFdntbRTOl0MQy50naXEuzE5VCXLamdAwiY
Di92/3iGc2oJUyl8qU2Tgy1ltA1mr+Hk/wvouEmK0ypf8j/5gEQOfsI9Wpo82z6/
WaA6ztY3wpOwLcH5gVo+JGbl2RcVOqe0xM/40yHRNxZLudGdsSgi/+sm8r8jDJFZ
ITIMXogVYoml0aZtYd2US0HTPTR5aLos8rmBWPCN/GjsJHqUBqHZVTT0g9O3iJwe
0lVMNSrpBsEkxyC7kaXluXJsffOO+LaEOgqiK4bPFlW/A7dmFmX7TN7co7hihCgy
RWbMABCU6fLyAiSQjE1bHRPUv6UsX9nnkScARE2m/cn57QsQhUVRGpyJxXHOvk+J
shTWQPJrBnDqvhuiImbo+jL/8oup2tDD8v30pt8+f2LyvB3dxAz4t83shYecTuWP
oIEAjI2w4ngCIfcyg67tJws7DSWGvGpC151wDSq7Fe6V6v1siGsKA0qSm6eHZhhE
NgILrkSEyXdsbL+l7pIbiWKn088RiVuxmCholddYX3z97RlvlAX641H92fHr1t93
4x+YY/Le7rNJAp4xZEj3VHEewZA5Snz4Lyo31BM2EUGN7Iht0NedEepn3HOKoCbC
JCTEb/0ACubdj0wxriBzo6z+OD0CI5JjX6zwzNOfSEGdpM4s0gJ3vcpPrPTq+acH
ITv7XGqziyP4s0KhS2SKBhh3ASs4TbvebvwtNY/oWJnH+/348jKYG2Uz1GPKZYcG
8GcSnTPGmEoENZYmKPg3T5iR015h2rUeCIO9ZQkkjfuZu8I1Sjf0zR1umL/qGLzB
w0IwT4jxOiFbGzt8Sx9q9E6EpYdoalBMgHx6g0sNpakEa05ADq4va6Idc4svtq2L
33wbMvATAFXHjR8jl3voEW7uugd9muOwSO9gAsKkzWhX5J0ucbGngEFbw5dfMVI3
ZrL/EQCNW8qcM34N7zxNLrJq6SJScLzu26yGofLjMnPYQcynv7hwkEy+uo9nfm63
59ApOmXsDFSDQR09jJqay5FJv5STtfrRFmjqVpucOkQaO1ghKS0pyufaOSZQU9eM
74sEkOCp4NOdvmYbjAzc0kOCsX6IOrqZceT9TVc4Q+akgWLYdwGvZ3fSKaS/+T1S
zS6qhy+C4BhzFk55zhOVuxyN4CjKCAGsP12DQEfZgEUTLc3gnDA+QdE0AGbv2QNI
zYhHWPkU/9i+po9pA9hMU13aWp/F7dbcShpb/nx9rsbJgmr4cV8VnVFxbXpCxmTu
hvMbeemSJmnfHnyXWCYk16m9h3DLoMjA7dkzCIwlk1LebNK132NpfUcMG5OTKZJ6
5vCkLboLyBdXVsJlcDYouPbzhHjSVqNDM2i9cfFuCx+1QtMN32cGMOVU/9EsqLI+
NA5JCpQNBMiRynYKXc4RXGixh0+3sWOXalPPlDtdIBMISCtgPqvy/H9UkCebudhH
6mH/ddLGsmdC84oCDiQk2LA8KZmldCZ38Wy1gFZy2gIGRrxDh1LiaAS+EMpVfqSO
MlBjEvK6iHOOMt4vkPTxd1FJ6U34XZQoFyoyEYTqD9Qg0qh0QmN7TmRWFu6sNDy+
L2NSGsrW29byrlCA8XnDrTB0gZBvZ2IRtRxE+BlueDnHdDwYfgIJDJQrFDe9ErtP
AmoZmTYL/K+f7/rjlxpHbVzwse0U3CyEu6OD2cZSpHJQ3Si5FDugIAtXnSsTTeG+
iqlHz8D6T3V8OvFxZZ1bH0qPjNmexAnnZrOmoVowKqjkjBO95B4dgZqzIXE30SZz
DnMbKkYcqjD7k1OSc4Na6NCqrEfH88sWUNYScUOpmAarw2GJ/x4IRfvLlEIqR90d
kDkoTbXB31JHstIPS6P6PRR3NV1hdey40Uxf2fgH1OwcAwlH29JZvhIZ+Q07u7Ds
H6HCEqxWy6R9Rb5HO9s0NPOIvBZgPEzvZYVbfP1HHAk/HHLqA4seWxk0OUyQzZ6Q
b5gH0JsOoemhfXfndwUeS3Trmc2WQjWis05/pXlyR6lFfcL3Ln0hUVONcDGan+wQ
8xwaQONBc4a7fMfswyzN2ZHLfzdBfHAkzHZp8spXOG9uoWXzvBL2NmBnZ2IXj+pC
BOAgtMokbVSG9a+8f0Lie1cvRWBhBvfDy6YQQ5UdZMCMshIUkei0xV8b7eGDmXsu
e5b86F1VSkArKmBZi3w1GJGoFTTUiyXgR4e7ckBo+lhHqlMhb0I0I3BlZkNeEo98
plt8C/p8Jtxnv924T2/EeZd/hLxS8J9dH8F5LCnDMIH4guf4Jrn4xIqKT9Jqw+j6
BrRNobWJGa9iq1VowYTMBGGr3oCOGZ032JXpYe08kKYThSeMc4Edo80keZLqj5ng
gKy8W+OPK2quRWgYEDMitxzHDlLtU1ccGc1d/ttTqpjm08iEs0QZIS8qLJ/rJAIL
4CzRQ3HgT0AWskq2FvhdqRPh/S+EHGNBhi50P7ahKQLOmHkepO+KgnizUswvFxa0
LCVyGgocayIqWzfVlIDzvP9m5urWmzwbsgqqIF6ERf9fK4vskIpXk4qOkC++xYNz
3+wH21/L5aa52cuKf0HI4MHxq7YRmFgaUcu6spdo8Ve6m6qOWqVMJXZ58CAe5R8V
AO049vrJ/3JGrFv0WTRX9cGTk3dUjiCVeoL+w/XkVVtDml0sll9b6s1PzVjQrWIn
OnrTguKqpdxn09HuaA8mACmY/cWks6tqpgwwM7HZZObhBFTQQ5r5YA1axwTD68G+
a/TOKZ8+2+Ra6TDZK3IM8IFyAJDD0Y7M90LPuq8SGgcDZfMnpokAvSB9AfYLok6D
yUYuf79+ONtpNx/DucomBCyOPjR4GZ4VqIK2mREI5Q+WfKiQuVg/XjKgjnf5bQkq
zxH/5TI3XchbKq7heS1B5rkXquAxUfphg9YyiS33f5OTuz4UrpBUoSj+yGArqUro
U8ITZdy6DDNPocQIHUF9A0n0uMyFXf4awXHlKyYYVwW00bXmUNJE5vz+WkvAtqz/
pUj5Bs+lizQNv0SJWroBXFNVuLTrMLSB0LbybjnRMscZfjPjaa9xgEHMpz33Wal5
qQC0rlcBZuetZxka8U1cQJbtMg2o2zEY2CV6O0Pa7nF9bZaKOjX5+xJL7wNX/PfB
sjr5ASIa18PYcJ2fzYWqEcumtrq48IUBSdXNygR6XlEz50/MpEGM9944b6Gj6YUl
P3oWJWBxhhGgTlUXaPkcT06vNQr8WipEp19tacBXlDqFphYyVEGzCMI/3NjqIjxo
3XWlgGrvuNHQWx5IqJAEOFSKB1hVWnwaLhennwc5MJts7xOvPatNOC+y6n/MoXrm
O8ReJg/+DdqRAWDK++P2wM+TCatRuYfh13lHlK2snzwRYPL7iS5yHj5ZY4z9n5EH
dP3xeFBsoIqvevrnrYM0k4FctTVGyuVVF0v5As56hjT2biYm7zYwW34wkWPzXQt6
Bvmk/TsAQtqVsW6zI2g+fmJPn/OyRghdDmGP374wnRH8WVG8JQjZNm/A1iWLhMoX
/YYoYqjF7k5DjRDPK5kGQpe6EnjUetB3vXLkNDpb7yrHi141tKAg+wUhzSeo911x
sJeYWjjzqJCZmqHCpu9+xQm0lvcVGrirU290fT1ou2EqDxl0hTQFgUqK648H5vze
5scRsRifAf+NzzcS3Ehz4KswZVjmaYd+0xvjZWIku16RTyC7VQ6qh15H+ZMVWajo
UGoBNyMbW7jfj9Dsx0/iFs1xH4ed/u8CSqH9/LAsxblFNzm/MDKiyJ/9h5morBlQ
2aHMwqoboQ/He5PvC3Zpi7F0mhfzcPS0RhuOkThh4p9YCwa9hcci4zRnP7AaM6tz
JvFNkSxky4WTyI9SaM5wjUvk6uXL82y59mNnaGf9E5Gdbq8FD2Mk1bKeknR7YSrl
eNfEYkEhyCL0jtxVLje3qeeVVHASaKHedzyVnkWybZ/LyF3IaRhvRozSzdm2q1Zo
2jPVa0Eq00T1PDI2NmSll+4kS1OyyChq7IH2IAh2qQcWIA/CVYxcg9s3SR+5GGm7
fDPZbxTAUR/w7/BJruNbWPTP+wbe8dqHLEO74EV2hv24TazAYl7t2nBoXnmwMs/o
Ajv2Uksw3oXZT7MGhleUGszAvXZEXmMTT8PkbK1x2OYd+DmriTiv3YNsg2Im1225
U2IEPeiS2tvRMXlLJJPYuVlobraCppAZaRLo/s+JBuhDMIE03TxF7nC8pXhyCKVv
0g1peDK64kUgQnxkqCkbpBy7y/GYYutok55/5q3LN29MHPFDxPS8PcjRCIOAL4xH
RA+kBBcEMOYUl9bI/g9ayPhyJQYQaqLhvj+9Fwwow1DDv3M3Wuh+wkCy5UUkmIlm
WSTMHeWxrb+21X32e1zQdoLn/mN6jLMYsTLrt08LepvN5Z278mPvtXIJLWyPryzQ
Tll5RaCX7i5X3ils0Dgn5HONWTE9zkkBcqjotjBL4LtdMTbcnZT0mLjutX8AkMq/
MRsk6aTKO5nYriWSlKwRzyjkior9KRmmn278dJqCsEQr7wtPflUI8YXH+y2nLL+W
mZEtRd9rO7Kc3xGnTHXaEJ+a7j97TeMe9HH+OxkXWytljv/TuRLWXqygwvMPyzmr
nq/heg7+N/M+1s2EWzdssP5p668pdsjp5YeNZoyoleH+6M4f6nrMZ/kSwdkXUtoB
76m1pGAklCuENjjtunUIXomYhXOi4IOY+u9IijrMQQukS2VO/Trv4f1Qf+k5gROi
q2lb+sYP0A3qmrRiY+tJOboLiUIClD2bGYZn2NVEZAICqT5R4rKa4t7PWP0IoaWI
yEMufBduLd9xerP3Nvljx0s8WmD/iSMFowyHkrxW4okK5GqgdVwppwuauqdFlrnF
SDIMLGLR5E+esdIr73hSXvrduvn29sjI5EL6gjUZrOoSGXQLQI1c86+wU0A6TioQ
SBZomQokadUHMRdax4rfb8AmRvCEVEh0qkW0Mo9JtqLOFAzag3j6DKRHPykm/Kli
iu7PoPCoP37/z3gKZjpEkxDj0jxNo1bsdXV8a/07XD3wEkhT13nGdVHSAgy6Ol6p
7nezjmyQPxkGvX9489b1Y/wjJiN5rxyYaBpR6HgWedVMCyyrN84j4nyxpB6YEDZY
0M0WhnkF65QCAnxA7GPPXdXVRKaPZEyFHKYTEFiJUkC2eiKGpgARZli9mdQ3Kfyr
vR+siNax1cA5gq+li9oZe/Hlesc5Tysh4lusFcUEi2qdROsh+Wf5UmueiNMKIB+y
g1sMjWPo51OWwfH9cb+eWKN8riApJgBVerXKqaeZbWaezJMPa2f37BBcwQE4fyct
7tq1scsx8bFQfmq0o+vj3RnjbIl6R9Nh7zzqPbg9x7/ADiWSaZtoN1LgZENHXZaL
Ig1uS4pyKldWXxtmVC5PEbquXmY5E5O7zlGG9R0pCZZgQ317Cz2lfikieaPhQsfr
embeH+1WA+v4Iw2zwzQDutM3CS1W/7SmZHyxym0XdiDdvQ/kW9lX7YALmIlE4uSp
QlUwf0y2WP44D78H41dGG+AiEWxzfsbh2U+P9zC3KP79UNb8IkI+UojQZoCDCi9n
/TucDARSNswsC0HNGSjJuU+/45AZzLzVh/vC4O0ZUQHMZV3NYmpRXhxR+sJ1A+cF
C/MY6cJhWGwWuJG2W6m1rwg0QfSMr9+FLea0wNRgtr7nFB5CvUPDC8iOHYWxahTA
lgmJsmTBWldop5IcJkKQ8WAidgZrTAeMISejatjjU4BZSfIDo8Ltg5swqEeUjvj+
kBGn42O56XJ7WCBJK8PMPqT1HhAFcli+4WyIBcgRdw2PLCqlFPFiBXnePdSY4Cgu
sVtRXBtd9Gd+benhnhKWBNLjWKYFA7ey9BlVb4+DF6T6QKj0TsUJWF9sDn6rN+fu
Cs2NvDQs5Nn3vn/rXpYFms4D7SGX10WB4yEMmDexuIai8NnWmGAc/zzQudHD2TfO
mmotB3KmeHE5dfurbIZeAfsR3GN1zbIaNh6AsdwlnuD9xZz5Sa2IJYn7NTwd+c6G
4gd9nKDUKqhn64dIM5hi98irW7EtLqkmcC49p4/3GIL2jCKz+Dn+0I7iX7GuC3kA
js541jtLM3yyQATIdlUJEbNmXPrhepn3VqAu953o0Vyj4k49DZp5K79el8WN3zMf
O6ErDH3HZYh9vRKOvl9ajLPzPvkwxcx1dztMCWDHQbkNjydVt+7hqxgoKBKU+RZt
KECt5n1F8oZ0IFqipa6ltm7u6kpUyn7ylccKJwlBH8rNzfJdYv8dhykpJR6F78dO
ncsDfmYWs8IuomJnEITnlmTpsI3GCmxsgtLDXYMGb5fThnzgq+o+Si3Im82GO4Ot
tCUw1M5uKZu1ec9f8kzm6U1pQQ3N9CkWRXEW4hQ+OosrUdFmqUdG+PoGpcnhutKH
3faZ6SSdsMv4/v3QQvlD0v65dByExLovzj1ZNAvSmPL7ZXcNGutfkYUPEZeIgJlH
UzQleCbsLHt3w0KKXuHy7Iak2Gf4nvG5QdijgRAB/yTtn3xPX33hAkzWL/7+rhOZ
XHlLzD2Xohi5OC0/U4TQlSKAE334FUvOFZLAJidLcrVBQyn6MVRGo/itWZm2X84I
73szxcaFcK8VSgjLq8rxP7Ygaf2GsBGPgOLwxS1Xj/dcVLUOaRHQFB1OBYl9eZSy
wNUC+qXLhcZGT7IW4ngHJq1u8crr5DMLoDm956uOFkXWw09aTLo39odoeC1f9kSX
v57wrSdn9O9Cfy39coDaSKF8LLiqc8eQtOTRw3G0hplxTJUCJOzcgM0ypUozfL7U
SeKPsy8yFMUA/ovj8BzgiGZRw4e0qpQtmB4g4oqK7hu41kHJO143nODFaDOonQxN
t0yr5KSaahKPynFmthddG3jr/Gi3hbXYxxNtr26SHNEn9KF+ahIkB35RuWyfjbkH
5LttWKs1jmura+k2a9qE3UO0qPYuSqwrkvKl/uvMfXN3lfnMsouOF48yl7Jq+Fe5
KDeuYxPgz+mfdiBpOk/Yc68UcNAedtR/6Hyg8HwKbzK3192+WLhzAoZWQdu60X+S
dh/GCLMvrRqE0oQxPQbF15narmPfD6A38Dpmv0YBvlBw1CzWXmM0AlMM/S+WvSLP
kWo45hdc3waIVVR5IKmx9D6q0aeSK7RIYvtd5+/wtgbIDcQQUium6oL8V36K7zrO
QG0PUH0Se4w4rNmCLO/nTr+6Me2CB3ZZ+fz+kAuPd+YsCdNYt+Y7xwoFk/Ad1XuD
1s2WwlMfD2ExPx7W9/M5mbL1y73XmMpTaJo8jjA3UUlqtrK/HnJFLej+dC7ZwoLa
ckQKEPQARhYcZEW0TvZYxdKX+q/zUxCjkd0IaHaUkfqGsRHn3mWdDg11ZwJuy3lb
ZhNf9jQi7rtHLJa1Z9LVUjV51D28Qdvv8fpt0dpaZF/Q8660HOos48gGXjp3VksH
uldSPWEdTAbn8Mv2i7W8vT5U706hkf0U/LYa+uI0wm1U6ROFRqBRmW0VRu+770H6
+MTMKnzKhiCQnKvO7eqe85PzNX3cEQpakMPg6G5nwWcE61Iiu5V4BbDsJN2xTSnR
O++Ftby1T/Gf0mVm9XJV461aFcTJ5ejhXRF5Qj4UwidXYZzHRPwRmApG85w3tfws
VvThGKq5YUsrLXc84eIETJUoFnK1GZ2Npnfbn3C/OaCZfBjF8zsWuKGdHMQpzcr7
yxJ7SX+UVymqbCf7wMSVZMSTwsn404ABOhvHYYXatlSAzti4KMx9h6CtgUewv85/
V4wP8qGpnO+XnYJxJ8L3nRl+JTmORtzQVla3XRw+V53rycKciIE2rLwmUZqiYh+7
gJP5NwHP3LRsIOWHbpCpUQa1d8E+i7vooP2KcFW+Gl85CIbJm7C+h0JpyKkad8Zv
w7c4cQpqXabju9wILEilHczM2iyGBRLprJjfCc0/MSj87Oy8K8doznE4TFCu7jjW
ioNzcKHrQfXHsKpKGTQ4kjkTH8LZ/Cu/+ueupqovUkmNpoxnrgmdbueE0/RaVtA5
uf4J8WeM1WLLg0VHa6+UV5kZoDJzD1F6L3JAnQVWSMD6jpUN3glmA8aG7lA+Xv3S
I5rdlmXt4R75qpvlUD3Z5OPlx3+Hvi1CV3Cr2agMtwDjznM7Dxo+MMmZ6t/gCFbm
889/j4VaE7cUhRKCL/FbXfNroxnDE6KxYhfLeSc0flmb2/u9iYLgt6hrq+4dcFbN
NBXFaoixJIZ/vZRJWw/WgHFj4v7DuJ0y9f5eZWaOZrMPKBmtIb1HtUlZHj6VbJT8
FR4Ip7cQpntlvsEENVGEJxrDWQGBBhpZn+kj2UepDJl7gct25nSRe1dLgJrwZy1u
31BfO7Q7MFpTdC9GV6Q1k4mI9QWF8x3OewYvsRfawalj4ewb4kMbSVFK8DQlSgA2
i0mwchz27WWypn/iZH3XmKbCfLyIclVDaLsSC7tAn1krjvp1lLaZhFprZ1b9jn/P
9QNhckMTlZxzivdYDam6d+m5jUk5Ju2aGp4Ffq9wUsUaQ/Bx4rzfPLFWm0QQFNOo
I6kMSA52XZ0lG2o3DhZtTiHswYd78woObOU77f4a7NbZSUOY/icd/pmagjKOSfps
Tf82Y8Eqm7tJBBW0hGrToHNwWXgkZ5ok7J0+qdIe66fj8uQuhGNo+Zg6FvC8iXTm
f/CzxG7IL2crq6RGN0601DYC6alrj6d3wLOgN+NgyYj5gkyPqg9Az6KEtub2juXg
Fpu/nMGC9nS0epy3d+OvLTvFYQ6EEFSVa/1jrKT9Sgl5U4q8FxRkuxxMGk6ynojZ
iLgwta5iS6h9hbl0QOnEZ0dkxaPU5XgAcTGay6FA70N5Mk5+f2iwDWZaO3xe1o9U
GdFpd8WuxSv/AvQrVDY8EM9BS8NgrmoBQ/JZe5JrL9Ni994/LcPl8uayVHz+yIGU
5SyoSKAc2X3jVR1mDDF/NxKVFeYHqSPnzoUD/sOOwJw96iAhHaOHaMbYmtz9lht4
syyS8iKSjW4r14i8ArSZMl84akE6ibZDB2ga3DcfUIhJRGqZfCLRYmgpHbYhQsQq
gbpcmtkhEhQy4cUHN0LHb2pDhSHfWhzX+2HjqamcA1HYAH/A5x4F36/wl+TuAVaj
DDT+p4G4wB9laFb1JZrMxCNWl9ohnKa8iRoIhwUbiBwqj3PMp+AbcpKGdynJOEQk
1Fktt3KPlG3cpIvi2n9tup6FxZtyMV0a7R5gGKuwZJuMtqZM9RP6nU19TL482NKn
6VdACXQg0by7LlfHqvQysiM6pcdR5ZK/Z8BGsi/e1y2jYe1qj+OR0FMuAnNzm0SU
Cy4S9x1R3P9p5OxEIxtApmFzSWgkwwKVgo8nPe8QSfhQvOPnufvuDvfA1+g5hiI+
HtbfiOhXl+yZkYwuMA0Ugj4xAM2AhmI5vh4kPmPJN2q8p52cs7SQtE9hmj/vlHef
6JAw37i36M4adnmyeqgjPnU6ulq2VxG1quVsenQ63nLnB/ujyaO0FqvrtmjviiQC
Ch2MCc3+esyiEFHin2e+EAB7coJG+/nAjmxCXKpZr6dMZVgyr4FDFVylXZ1GOHbR
BWW7bURvXpUWhTIy0OurXrOJK6bKH0GK1xWfhsovyfGqM/mqRi/r7k7k1O/h8gRb
TTYA/QsFkgywoSYdz5J6kVnRCVjV/BTR9fTIXnU1U3upfHp3ZvVWzY3csBIGJmq3
DiAGUvszg20OPteEvwz+TdY+Uj2+c4YGlve1kRjDY9MXJ6nk+2YArnTVqLheyR1U
zzyjBnpl0jBNprzd1VhvBCqxaCj5JjVMMLKraMGEvSbF48WE3Bpkd0hz5Qkn79yX
kfVlurWCUMoObugVbPeQlIysiolCns+28k7HKDCo3JwsQO98a668udMOX2gexzBT
3YxgZGMMq+AomSClcKkZ66VXOc3n4vFu3FPSP2MVdnZlm2rLJOldftvYIQp9tqFc
c+w2NuBA0sIXM65vwulbUF7bMBpoqWK7cgxX7qEqGV3W/ihqGRKjFrzxMDWixiIJ
rm7vZk+3/Exld2nFJvGTLvfGuil4V4IRBjqI15LdDvc7HtFBH5k80cAtxbUG3VU6
8pcfKvi6RgS6Ec6nxl5Ya8rvCcF+70FA74IBoWOUyhUv5qvYvyTUjbiqJ7AgJ0rS
+SSq5odqMLZ+J/xDxlmRiodERsuf46DJwBGM6BgvquSmtry6N2a/J6PkHuBsI+7A
+1t3WOjWMD6zUya5ZstPBUWVrgZAbdxn07ydm7K+qJWkBfHM/aIAPaOxXldIhAJ2
DawActEW6880rUT4nKH5rvLe/Ut6Ijw1eWPsBUG3UIELDxtz73sbWFGLM+ibPuCJ
oJaPzELbiEgj7jnxybS5yl0M/NdlZHb5n7P0uKbFcfw5rUyYfoEOLA9nI1qtMK/G
ByOoLjZsOju7DFVlWi33Le7tNBwFKHMNFz5yxPchwn1ST41v3VzPAiExqgi9JcZ+
t0DKro0TER/SX4o+ZXQn6Y4Jgsr7+6IJnRuZTe3DsB6dwXXKHBYsx5C5sFsAk0oj
LF+Q0IEMnOS1Zsa8ezJb/RTzclqbwMvQeGeTsCvzR6wBrE4dHbwmV2t7AaNFTgjb
Qa8o6HxcyY5Iykes/XKhL99d3/E7mh967agojCcCgcWsSRSULsfVul30md4dvrNr
UX5bW8idYgPs5/TEoJ0r/CMB0YmUP+0JsUjBZ9bnekQ7YvIpoiR5OAj+KSrv5c4S
luS6DDTGW9yGqTWEjjaDPcGhMeNmM4JrnF88FpUXEmJOd0kZnrobVpggOj1I1D6m
qD0pC9Hmo7LRHZuSd7FzKo3Js6TsqKc+eiN7kFGm+KwodWs61/ziOWFxy9c/5stb
m/24wHNgRsr7Isj0aZdYpEYQmw7OMstL743QmFXXs0uFan7iZzA0MJ68vJ2M40xM
6FAWGQagcVowRkEBlWlYbQYy3iZx3TVojFEoQT0pmQJzv5tj3Ka3zseSnDcbpKTv
RnjDFvkpwbSRhUgAtGqdFed3TDhQvT2+QsmUxR09gT/cFQGuPBS7JoVHu7q20Mxi
8snjjZPBsxy75C5pGbDkiAxCfHRKjUMnJRaoMyUiUThDxF8B93XVcn9qFpNY8bns
/pRIyaoOE4EHwpr07fJ3nxjfwJuru873rcwy5bpaHSUmT8qN9TrNVotdKZzLq/xw
pUbjFzV5ktke72v1aaIIYedoHPLoSPwNJ/pJSg34yNSmLufu4Rg1DYK13RdcMxc1
5lJN8KxrLFVtoqrMFMk1ykHh3ohNkXPf7KcvUSdLuK6F/ScfFPPFIJMkeXzxrmL2
9ADA2ocGtA/kwAajlqnMaeDX0Z1yo5bohfZrsT19DU/8uhjVNueDAxtT048PZh47
My6STqJUpMo1VFOlCIzUY6BJhPtrC++YuKk0gOY0E4zcsGCEDVj3i8ceJvWYUkc9
snSby2oVYuWlMaQRiG3b77+EVMmOgeThvAtjLRPb5wHT4BCQHOhbBB0S6XGU8zp4
7HWU5rhA0Z/3SdUZ6I1yJ1DSC/QiQ3NuJfN9OSy/MG+Obua6MPcuuGdrSBaOAXUX
fdI4l3ZHbxAePBGNXTBCdzr6iwANRtOdC6QEKbHGA1kA6/+8MuZ0CCGZsXQhj04o
6i1DpoXIsn5QvGxiZEXCHQqanjqQusDQjysmQnaUMm1Y57XTkf9/D3/whHFh/82T
zSfBpvY7LKqkyaPd6wWkCRkDtr7XMh8tslbGs+Rh0dTIjkNtNJtnVRoOSFlinqey
Yi9nvfigg+nd7UEkg2hCtLXYl7BQz7ZYXS32XUaer6a1R2pECFFnT2Fj5ZxWok68
UqtKFzRm/P8p8e5cawtEd3HzNvZpibICQDNjQOkhHHt5EnoBkP1nDX1KjPbKypbD
y+S/xGZW0HJIKAMBimO4AgLejBRLdxkRwx3w0iTqn3pO8LifobplT3UPedRtt0hi
/y1PsyQi7tJU1aVop8bC76NDQjth41qAnQyls3L88MYb01b8t04fYL070LBQEqhL
yiWCvw0F/RFJ1qM1zF5XpqZ2XC86imHA1AHvjiVcc9cJLMEaqvEvwIiS2KPftDM4
pKJDW55T6bGlyd6X4mN1L9kfxkZVfqcdW/4gq5Mtd4l/nXZkb52X8jRtvdrPxB6P
Z5uifGepBOFSdJP49qRihD95AhV8uHUU2X88REkG255NtpJaO8D0jC/CBe5Yh18O
AOzioAKM8BUSuCvkgN/j6rBIbR3i4VFOmVehphRXAeTKC6D1ktoP1O6YCortM420
7ebM+hYc0rn7XaGYG0t4bo4nNFPujXl/bNkzXGS7WlYzu/JZXshbaUNZBLvOeybR
ua4ojs5/W8ur6WGGLx5nazcow3UKaOD9FXo+8MiPONPWQgRJjQTPou4LblFG4ge2
U5KXSDVWxdWZx4HPKc2qspXjg43R76EP3NbHM/FU60e0erDj4DbGPbTbphvIBWZd
4LiMvcAqvMPe/3qPG/I/k148UPqZBG4yYGCGwCQ94Sa2LQGQrx8xkYNHnRumJH95
rXs6LC9hWop9Y5VI8My/5smD5sEGdsC9Wjih/tLgkR3QHOMVaKlSGKQYkcNZN533
Up9RsBRNYYj+MorJuRkVEle88fPKg53e10rD66M9x3T+RITM5ZLTHNcR2APRHoV0
ZOR5iKQnpk59QvtvxW3Hkj54DM6mMb4gGYQZazH2VjAyFxjA81VpA7qPqydYRF5I
jwhQw9M3VeJIbRPGYOBefHnBbH+ffgr/Dhed9yS3rCDJmWLZf8IoaHHw2AmDCFil
81l6gaTF0yugMpbgmHbdp+PrVJftioXkv8D8S+IbYTKxkDrdc9EfKlse2BmDv6Ph
NXpEsPGvCwIkGkeRaQlbnrmot6wmn3NiPKHmN44LoXb293wUiOPrRnZj7xZm8PoO
SIH8xWB/Tpo7m9ofYOjHSxAyoAlEUc48pKU6AANDM2P14isDswXRv43U02bPzqyi
8r0LqV8p5yybhXZeB4mZQQvadehEVUovfUkOIVga7PqzvPFFVxCRSlX0uKPSqg9t
iLGSEnB6hLjs2gIQ/E3Wf0MlS2cwGFqiSiWe3GA61oQ/xu4rHGm/zsXN86MimQEi
zywwMlqdmw9sG6U2l48vkVSUyXW30HhtXNnDgz3weNEMdZflwyjAZ6zti4Hc0A70
lGCFBWcob1LnsjzAy3O2OxW0yO46DLyVLUbzNoIA5eAMcCyHhbhzkYXrTJawgO4M
UkGzdER6wMqgUKFhtGluNTNtkOx16BtYHct1+v5ZI8l4rYpiMCZInJ18q6mPsvZE
0BY1q3/ChGuxzrLyWB9xcsWFR0rB7GsVh3+gY5bm6PWWk9Zk+8b4ZxXXBnvfpAFJ
jNqHOclI4lKUA1HvDNJKf4PCXLad1ZvtrepZjF1gNiG97RXc4GLpAk3DgtnSd4ns
hFXbub1ud2Dc2RViU0bezVOOpN7RfYKCZMMoB8Q3t0RkQEhK63SCVpCtjRo8f0gl
zbibn25aZVO+V+sPuasO31vt15ySfOUARTgNp/iVhk5VoZA7LtADUtL7uHWRAkQi
ZOp+LqWO7GRQ/M5haP5xgCxTr9QaKWOh4gxOjboR5JYmPvIqbbAG9hFap29dQEDG
5yG9bnj+szS/X3vuXrHZ5DIe09/N2X7LPT2A9uDATMQR8sL9KlyD2Ghh/BW2zexN
QoAGET1oXPn8tmBsdt81Pb11gZlL/HoujKTDI8m5ikvgsw3uTcgFqwUtfsk3IyPm
CbNsEFgz6iWQSBwR5nQCZIF0ntFuokbwjtqobi2d50rikGFdVMqxDqTg/kyp/GPw
rZtV+u1z7yKD2jXywgFMfLc39Lhyz98Ntk+qp/X15BNqXNF4pBI3+DV6NzPoNI34
b4tHFAYMeDnErMH98pLvvnpeW5x8UkQEWIbZMeDAEuT35G3GoezvDZXxdCegvezo
EqZafk6sqJM3X9I/bknPEmUH9thj+4qlkFIGdlVGA7Kps6opDhbpUBKo7Eqygxty
9uwM/W8Kg21JPYUkvaaqDtLIle6eh0lLUY8V2OYW53u4s8KOHA2UgAUSN7kdOLgo
P5dwZJyo62eFjvAY/dWcKZ3E2ddonZwbQNOvLtUQ6RRktvCZfAM5E2Y1cKLcWcES
KtbYeXV/2LAHMHF+3DYwIu8o19+c6hpP9nNXyxlIjaJMwQb2tE6ET0mIOJ2Aut3t
l58spuezIPBmqnNVV+Qxm+hYbOMtc9y1SoTM4iVHS4eAUgDnw/X55wcBoLh/9ctH
DBK8izxDtUpDrb6yGNDW5C7zbDUmzFW1CjyQ9hmHgG4XOqGkSSeWQH5fkt81eMVj
/J5CSyX1R6b7ZEaGc5x8/Axp1TrKPUIKHrqtpQNvfGfbRaGr6z1moY0JEQM18DhN
lqjloQaw37mK1W8S50rmu+mrgH2xiNsRzch+Ta0FOuvzFqGfIWVBrUwZRBUVtg+b
bP2hsJXPfMdT0Pi8omXjb3cmICr+feCgrz23+pLLVsxhhGV9W2NIVwDAYUMO6mgC
iG88Sb1zpiwx7tW7MbZn/ny3d0I267ooLcN3ta46h2qtX9A2z02z7IA2eRPKXRQ7
o6sFKMjcUEVPc2GQEjPmSCb6ellYYaecivTmDlY0R1pnkvPeHKq0MeG04ln51AIh
sFE38DLZX1QpwJ8UmLlM+QKkzn2k3I0jv7ItFFEk1lVzJq2KAYQjhyAPOGmUKwKA
7+d0O00kmKdfn0r/FlSYs1+6oqw9ZLAuA7xBgrb677oypNURCEPIV65Sy149uMTf
PHJtSZwhy/Lm4DFNBgxV7mRxMeda/dBoFqAJ7nwy8AYndTfkJAF4zL/E80c+BFhD
Qca+HKvui2IVJqpt8uLROCkvkS7CcjbFyrcsU3jypsbHQB+4iCIt4F3+go6Jqy/d
mexA6b87UqczyHWTS2wjvOPB4ZucvUclLp3vSCPrIGCQ8GtMHLiM9fQ0Rfxaqi8v
X1KYoZN8DmPS7L9bIO73NaRtp/kP2EkA/NQrli78sGIzYohMbvTnyi2iF1Xm7vgp
EJDWPr5yrMl95qYBTpxtjAVfqGGV/Ay+wdFpQ0DaEg7YvyzMaaSxzkEjQFwWv5nn
44edQ4UCiSPuszij8I6hCpO8iBZWbybORWo52UGcWBYQvhwHuJFm7NPsenGKYM5P
j1dn/WE1udrUSfSPynRxiXVLPH1AsGyYULe7te7fGuiF58dqMi+liwojQbZSNlyN
1ojV2O+7FBL0BesojPzbZ2iESZlvkih9r+1gqB53xIvHXy0pNRCYXGz26eRsGgZY
80BKH5GbWZFv1eOXdqKD1Ioz8qSvv+E2/uxgsuWyMHUGV8br/g+sGvjVQDOnzAxF
mRIWEG/jf/AvD72xm7+0BE1GXtr8hoUaPnIa0g9xWolUDQDrYb75Z6ptNonIlEFU
N7m9OSvyzLTd8YnwFU2YKmtQga71FCtXeRLE3uzJx2//+KZCjQBjY38XNhyVZtTZ
c81pw7tbq6t1Lry1jr/aryXuYo+eMcpnhettektVBODl/3xFW9AUrXd6AL1194+M
onUNSbpwZDX4rWOp+Azlph7oUvFA43z1SGMRSSo+a221S2CJQnpMp9sfwIC3Ls46
xqYO3PElasZFesZBw4cxB+Jkiv/N1rhWSZKilgrqJQEhfPgwMZ3PXm6r/tDsnYWU
+2EIueCtMijp1jXoxHpYgOSEwbelhzHKTEoLT0AqY+nJwP98k3FSZ1wsIEqxdcLr
Zwmz3HEHoTWWk6GFw+AEzNgTjzQXCQGKxR8NZ9+3xpkLD+jJV0mfnVuSvwp/CcTQ
1t1DzCMcwJ2YhFlRdmSlzzAYstDY+yWATKpg2GKFhffd8E/z7dqwRG/BVpu9cuT0
kyGueKaXHaIKYb9lGoohAMRKWxjxGdCY/Ez/ig/ohXnNGxhgG2c8l9JmqNgYmFRv
MV+7IUW4WvncF9MR19bbdtKabi83PcCMDUR1G8M4aRjtTQ0+I+I0f1UGtAPO+Iex
8mKY7rjzZJqyj4Y6gnasRzCXZIElbHVPn8312Xb+aKSfeLAnC7okth0wTfi6Re1R
4Dmi9GdmRdpvLPmLAGJumpTPRv23jnyLQ4Og9IPYRaW1E1LuJd4o+HyciUCY8Rbp
NyyyCt2mq+Td/tmjciLFR+1O2Ds0jyO14/VPzG6W3TpZhgPQP1JnQ0r2tnPXb5wA
tYl7h3836zIedIkgwpEO2WmLiLxhnwRUF17q1wCnQQkhMnnWocIoHucjrJVPapiv
zjVPdlz7v0CEwcudE4JjIPCs+4Wi2PQcb89qNjeaaU+LARkluzOx87YMaNNyVN0j
6A3Ma5oyYVxqm2tnT4Gdd8/qcqktX4duqzhB0uup1UNE9bIqxgD2V8RimS3g4iN2
XLbkxpJk9ptZsL/W8/WVmSrd4Fbn3OwgCIBdSd4mShitiwBE6hHmn4Ao3ljtQh6H
vxT5fIwYj1BS3VobN3l7B7YnR8GbHXXlZAYRvq4+O0szRRhcRoNJYuAkIjNq1+/c
FhXugXek3zIZ6h30M94SL4KkSnzxpvOywPmX+3dJSAfNfiXSGo2qz1M01hRVf9Or
8B2uX2yU6denN4QcXtCrIkKfavMiFrHRGojCaNalxjNDGFCcfwlhKIo/zNiQqNN8
K9WgHmnhNiEFftzP3BsUyrwiYDYhTgBREuUekGd/XTFyqVeerq00Y7Ijjz0gQGTd
0mcLnVVLrlyY/qeELzbVTTZs9ptU7eeBBNzrg+zJhZ0nU0hb9UxiYPpDVx3tquOB
4XW8gIELj9JJTKPVGDvQa5qj6nTMZa3qGrCdVLgqLWE7vXedBDa+hW1EWGRSXojM
WAWeS1ePF/Uonl8h4v/Q7LwT7ZyWXXwRzuDeD3Kq4EfKVceQkp13pyx4TrfbGvUn
3LsNyZZDpt/o85cBRjIBg1glknNM2g8mNhCSgMtvYyKV8KRYToTs/LLL2wwf4Kx/
0ZaLhapjg5aGZrq4OioflyEe1VOLPFyX6KOnXDmqArIw2e8AL+ZESL18oQ7QQ99t
HnVSkPBEzHmQUIdt4e41rAnncOF9dEkjn5pAp3kjWIcaSmfk64ZIYA6FhUtEZgVD
Ak5Sfl2gxLnBru2WMsmyq4lp9hVaoi2fZKRKXO/8DGr9HFkldeZE7TI9psJTDz2S
DbGyncCMSbnE2mWMTwnj1VtKIuesNYOXTIQ9NyaxBMau9dXiWSVCGuhjNxsKPAQK
SbfhJe5VUoRnZlCNgw/CPTvliDGBi7s4wI+Mc4z/AATXE4/vvYeWYdxeP0HQkxKq
vDWz3A/et7nnS1C9ntLbCaN65ja/OnI7Daj13o7ui6+Ld/Wp/8Bs7556W1Nol/Gg
EYoponWChVNoG+Xww0EAn6Lywwe7RoUL++sQ7XAwqhHU8+bo3qY6ISDljN70exh4
hljXGR4Ihi32J+3Td8oNfIHnPjkx1mYLqTJu/mIt0ZIJb5O30DZhgNWO9aaaCek8
58V+HiwkLA16+MNHXPnCJhbp5eQVSP+3E3l7jbYlKlC6zGpkQL1ZjQK/RNq9MLzu
PzVhTsQA/6nzbod1k/0weShsUR3V3ce8O9i0v3w3pE1AqAmBJOZoGM4ePLlAttNi
Zjdfk6Pti1SAmbbAZWhjQWeTA6iu+pxawgWiMGvdCcex0pRniiNIihUM0R7y7zNy
LWtMR8zVY5MQW56UeIWShr9xK1G2avjxmFckck3HQ6gsSWqCMfmMD7R8gMRTttmk
2C6+4vDdG4915Wyr6f9PAXwXpQIkcBWm0aQl/4TUNrUkFmmc7dNAg2yyHWElQd7k
ZZWwtoKkvxHUKYvLbCjWH2kluYQ8PsloIsy9qWLLlKcsiRAnB6nFO39wZ7+DQ+jf
N74VdQRWVgVgTQmnUv4AzpIqF1oIi2MIZd8reu+H5g/8PmvBt56Xt2dNp+SFMaOj
KvPpoqZVd/40hiKvAaQeg6rCOhWl4Bw25juSXL5GbwE6gS1a2UaXXx2fNHy8pYqg
uITyWMycjz1gWs5Na8FpQaR5DMfQlnmAWUjxjvqZVXLASZtadQYqqY9iBHHkuKie
IqNLpENHQAQj8UGuBxtQWpLPFNXVlHygt2Kyl1AS5r2LfawzKV/tI8sm0mxvUbXG
qhj14C9LgMHDlEn9JVp+XW4p+8lEzh1ePT6xXbfAUuC60N9NJ+tWJp0sgHVOOMDX
Ccj+w0ZKrysQqI14x7C6wBCFBdIjRTBa4IEglidqmx3hHn8Hp9YNvVmhownLhffM
MYqRWdKIXU5cfMC95BypgpFmmJ0DO0MYgaEGnG4xogWJSMsQFUv+s5c2VPOeGryl
Gi8xWTGYJx1QKQdOtvzKGjg5yZU8AplWdnNVUlLHJTuVyuJbbJpHwbNVp2mSI+5B
v7G111l//Q0/naafAI8YtV/iaIjQ+b7WQApDOQ270E5cFHnUIzIRYaupLMwkW2NC
n3Y+SA01EXtv0g2JtSWpY+r91TaRhVYq8skXqx/pcsDtjnVIIrxkDbqOrrqj0tKu
w/zG8MdF+d4LWGeKTApSS2uWQ/qy86NDusfObEqS7Peft9Q099UZWsXSzpHTAKTF
jnQRRYqfSj/KgRNo3CRs0jI50naWRM6qwBPr5FkfSKddC+YEtul33HdDA3WPeR4b
ewbMsIwxUluP8SK9rVy7J9TJjoG6nvemm/yZWf3QF7U7UCY0Di0jMLSnBydw84lP
kZEEf7lToT21xMZAlnoT2Tx+bVrXuVYSc0g63pqy2aAm4bXA9toN5oMOA6ItqaQm
yhBL4pSBXPiWGSBENH9lcU6OwQWIJUXR2eC3a/40qz69QpQr2wpP8XqGJFpaA3aM
XZjTicvj8LiUJ3DUvuYoJc/k0lkWIfe0hzn8X781yV+yQzP/lXi4QGj+OG1TyE9I
uK/rE/u+A0aJS9rcY2Rbe5vbCHacp8EKyolIp19H20vIQCoycgH6w3/iua/UnL5V
mX2KphvU9kEW3HkSETkibVPBkSLi0zScoowKI980mcMgdmrEzlq6gtJmBXjNW8Pp
OmqKRIkTADPI2EvazLXvZshKPpkUJNUBXumFRyLMLr/9TNl7+mRUFw+ZmGWMUFvu
QfmiJ7xnba1iA3HEhq7o1UhROXZUMQd9KqfWOeZwoLphOZYu5bohTmmJQEi6EBZ7
VwiwODBddlmTqcClzP7Rk6HIroZsZ4R8BDfhk7md0rVF9Ec2mSBGlLfZgQzILxz5
Ux42xVifRJcT8FcE3HH2N7zjmyAYbsV9J/OhQaa3wnoQ154gyXw5jTTmKzAV8CPU
Hm5WHY0TYx7KuZh+WQSltT8m1ZpSzW+Gcqf3AG9geYY8oKGfKUohaN0e8p7GSdd0
8ZkPh5qEU2nLJ0zaLn0gZ1NxF6K4Ut1Dig7rsgIB0vyjf8Tok8IKwJYdTpsofhlp
+yBjpx3guFAoNjFDfOXMuK6fmKt4UfQ4TzedPSNm5X5Xbuvt3OPHPibeLv8pJHLH
5/3BflNyJTdiGWrhdDfQ1+iij8tNDvtro2PzRxkKHSSayuJTdApnCh3xxQIOSoeX
YSs0HtSv109TXc2H216uD8jFkzz7QSsA7sQysOtbpMvJgTlqWQLpo9pYHkmshUgN
Xlvjn4Dbrq4bl2tf1llAdal0DVp7RVHOxzySPoUwfpOoc9AevEuH/lDbAb4F9rbP
DviQCQ2Fy8yImhQm50TXyihskgLUWYmuHArSxliS/TKcx+oui76gT/GPxPQl0D0i
lQwStM9HExbosq4n4VTt0jpoCSuJmYbSzJ+2LymkiE1nuGIUrkYKOStqiO8yJtp8
QBEOeXqvQp1YYTucJPsqhsWXO7X96ZB7wbXJOpRxIlX2RRVMzHuNR2QW0j6bixoi
ob8fdalbOTtCWHjcket7HrQ7KLyhSGyOg4AmaC61vQ+2JcHOBYGGp6I5DEo4Y1Zi
BS93B5eBjYc4+7knjfx4XxFTXO7pG5acKo5mSdybUNlB97nLxRyFHjNpBYauuvZ0
l4epukN2gb6Fn5FcbCnRQo8P+24p9LZdSfGNquGGYFd+bSjBqY+eRDNcqdFkJGFx
JgTuBkNUObmhcgYjg42/8Pb6VArAsn8AbB+QjspFxvR3Bu4ZyhCVTjTTAerxdvkh
XY04dVfitgveIpct0sucvR1KWf8TNEk8OrNke8Kuv7i8psaHX33ZObQZBo3ghJwM
tCbfeb39EYXYxFrqc6vnxypRugxXPmjyE0DR6S/HqHW8aMNQO99FUrBfKTwntBNG
JAgPL86oOYLhC4H0d2/1mak5g9ha2ubpseYqI8xda3VyFptt8EfMX17P6Tu0Rntg
NELL1ixrQpbhrKGdm2Haxuj0qRNyiJDuDwNq1JYSXP1jjmV1k9TcWk2zafR14GsG
bukhb3seUu6POgRMRdTPp6MeUohk1QDJZNdndde4cIVTjKx/Kk3nvhQuS0h3ppqM
91jViQGSvnoAgJxxkuok/4SXncuKMSbq2hOdEtj8jTn7R+yW4lrhFEKIP7jz91Se
BAOvRJ8arOyBf/ziev3hzOfe8MIZd4k2wrrpw5IcPC0lLvfAwgwyCnoeda6SaoFw
wabCs5QdJZl3eyS0b2nnYvjS+fAir3apXZHeY3eWcxrag085Xzoptwob2Wr+y7c/
+NRdwTxPdB5WxpMoYnu+1PpluVVECKrS02XboABae7TiXWAkfMKhZ067EeABiqPo
pk11rO3rX6ERQ5LuDmXyCBBEA/K7ifjOGqjx2xHUOPZy/2f3KSuWyAzUYEYljw4P
5fECj39K5eMNOvcUjacnojGmq6BxP9aVqnHH5LvbnEsnOzf0NszvrSGrKnsCVZUN
JPALAdRjDdU61ZCicnwxSSm6YqPxW2uGfQS0Pq1jPKKdeMadnSxCA//jdF5/b3hL
ZGsYY6A3niAMu2XX42/+pJ9WLx3YmX+MbTwHbmwKbeBYrZXbxYNJA31L6UXeTZA3
3rRPiod+D86INiS200wFN+kTuBhfaz3ynlgjsuEM0l9uUVrfIlqP5Ax/Xsk1tQ8v
nxRPJh3V6wuMqXCTehqE5O9ikiUfaHukE/8z7UdPsiMEsz0ZK3BpuRFOlnN5X5vj
FzomTHwIkCeb8zofXrZj8rX8kS/f/aRKiMVsy5vMZlPj0n67bpQE7GWQiUQPBgEl
rkRuOtexIRpucihqLi6Tdh22kDHWFn0mqiHBCWzkdMpuXcjskRtoX8jUe3GNgWTR
61FRx4TUH/fYFdsI3ubvvVfQBpo3wXAx1sKzK0pthFieBB5H/2Lbld7jVH9SRe1A
fmCxJE0zieNr5bE8B1tDp3ZQCRtnoF1upMn8A2IMXyJcx44xvDmi7acdYDgaR5yX
k9Uo70gmvgaLMjrKXssIElT6ww0hXawAEAEZAGFAcAJ6jM+KczyWdzlfZCjRDwzh
e7Yt0zFV8+IOmqk/cqX4BmMX+KmSFjS/yUSG2/Rx9yGGPiGsRDCjm0deyD0wGwFb
tvfc2nIVD5NzjMWx1alwjRAzqoB/cbh1egf6ReJI7/hd2a4f6Tlaao3wKk+8d+XN
X0fe5WgKZ9tUhsIxp+UfKUhwscyPJfBknuW+CjusfdLg0bxq5/io0F/yIHV+V5uJ
GkFrWzNcRK5UiHTZAdjyr1qeFkocwvkASWJ9y65UFicJs67PNDMc+5+/UyFociWt
cWgJpcW4t7pL5R+deNbJUTBgLLBCcJ6gJ2lEOukr7tkMl9qtcV3CX0ehwmG5Nte8
TBE5f8ANzExUFnN5yMlYCBdBRWnOW3pJsf089BHGc8pzPiNjtP+NRmotmKu0DgAW
XQgl6udQ908er9VzZYfyLUJDr2BUYNAn/SEZFpH5fV1Bxb33js6+f0Es6nYsU7tv
bk9UL9AAVzZ+BHEJyBja+7GI2M4Y81PUfl8EEe/Ik5tdCh0Ol9g//FYfA4QHJHIf
oXUdFtAFgcb5Y5tUXExr8iQtFVWFRV+yNesVtb/sHusMrA7ZdeqrwyLADB1n8OOi
nxfYbE9w2JKlcl2wB0MhrSAqk5LNiKa8ME2yzn+VxhbCMTF0lXZnGnSZCYBZXWxD
O1kEdbyIjPBafUQl6gSh59hgP+c+Zub6JJ2FO93y5XCk7m1rl0q3FSHevAsYzJnc
ADCqpAycf5+9C0NTqpW7dNYj/eXz0pSJg7S33Mxk4k5W42RbY+oVdzyvGdqiuuLO
NTcumKYMieNs76V+0YaDAhCzdvm940Njk/NyjcZXOUG2XeDw8+Cfcy/y2IWiReeG
2Qak9sKACKpDc72atskSOoLrdTzTtw2xTgd4aOx7YYrTC2w/L4p7W9m0070jVOb4
IR++18OQngjuH9HiKqN9YqMMA4k6mP3eXwtRtAVg8OhZEw5QUnftq3Rjyxp1eR5W
lsesrIYdyqKlpKjwHlyvae9TuOx4fsfHTArx+L1a8jSluIfKJ7+lQ77pm9SPn3t1
gYFf5f8XpYbWoFQRxdtibHC6ASWwHu1QIGzJOCJRWNooJp1EWY+tRVZaf+y/J0sZ
C6hsYWgESqwc0zaqvj6b7DXY1AcnRBbKqundB8Ol+kE09dOF9fnRRkw8oM+OeAUB
alAE8T3GZJ+CsBfQ61u2X/cKI996ZXOaC0f0tEODVhTQ6yVtL5rwn81owOHD/0nt
9Kwv5gk/yplKWndtRFLduBn0QPrQ6gLGw58cyWmQpbftXjkdULAXeCTfRFxgtGtk
xDwdXH/G1E1m14uhK5bsWsE+wzWIwLxONDrgrdfQ5feIjsLYU+Or1hDgr3txZInG
rbKpACPuP5Sh12XeGk5rHKSXzkpr1mF596fqMWIA/ZukBbS1pzIWuBJpOENgwyE0
v3BvskXJT/ElVZQY7WBig47/w1YUpCrEWvnXPksRvbbmGlUQoLmO0OgJ4hfSNji/
BbYLnxRTPJPSzHOcfeetrUNMgw0FNx0L6NXR+NlFWTpNHzPx0tVzGqfSEZpvmdch
xoZekqGvXRMPc9kGGoDc95oTNlGHQMhXr2hyi0cdCyv5Q8EjEhT/HubZrAJIkyys
8VhKUgyu5HTyx9f55KnKAKoBJCvWUFTzMXpJUkFnluVuAzLnUuqSLlDriDeOjgmf
v8fZPoh0VLKijQiiNV6BFMTSBkEePArf3frfpRlZOUqp7/VsNkITGD5oVORjv6WS
0A7dpQBA3hvKLe1+f15kjhH/yYW8FgzmtCIyYjvUvVJtLUk01Kn3rRxBB/LL1whT
mVD6CLGutmQR2Wse5nCvNGhZBEdyKXk2dP5SqTC39GQSUHa07CzvxUnoEXzBH8ak
Iy862LvwNIXWhP4Ou+pxpUX0ZElKAbyCBMVzjj2AE90iV9UBvax7H5GIDgXDbjIN
z/jDkbygnQTgzrfh0bDcucNHTEcGEtPPwDK7J2n/saoY4qRxjuOB7a47MwmZ7jrK
kOeA2Si28fmLkM+/GlvdGwsKGSoRly72CUiS2+PIWx2XQPnm9m1dYabSgniOUGM0
fn8B1s/x7W/Ag9az/aGhPEoW9Y4FpIXdkLWMD8PpEssACXNzYvLJTL5LX0h62PUT
3abQqRmt4U+48Y/x37gbaz6zn+MYjjaGYnZIq6wN8XBLDlOkT6ezT2c/CqtHgcPb
qEO6LxgB66NCYCHeQaMrb+NzWPV9cTAdT7TGC02kiiB5bTlTUCLSxy+srXhAQhjr
+JN0jkfjZE4ONDO07PwgGZsqrVWDZrcQ47YP+JPhPKp0THtNa8PSR+4rPuN09a6K
+xxBiVzDQ6lQa2WmhdAZjcO7sptR77vi101pyO4p8agaWa8akwCrBKM4k9FhqfV8
mtohDAt+DOnxRlUR6lT8ULXYW+njvH5xbUiMXA0VuVnHygfDp5AlBgTFosBB6G+a
jPLLg8OK6cTDAxQCCEcKuYu72+fpvHfNSoDnTpOgcmFrvQ62Ch5Hp24T6pwG+4eU
7q0aBAmWpiMijHE0Uogkc2muax1gQ3RZ7MWlXlqGkjOHheS177lOV2aIGYyAKRbS
+9GCSrCkK2VpM95tkJU71xeIyfFIrTqR6MuXBRaem/DLrc+qgoStoKND9+JPUkmi
DW0xkzfBS2GddCgS4WJwcUhQStmKm7/2wvbgmduET8QlDCrBn8ygubrDWrn7+tFE
tB2OteGGVjxJq/PfmjjSCUbwwk+b+Wn4IxmNFOOw9hRXdJtUh3RdGH+L0xySxnWb
KZoGzV2H9/BBcjrpgwmL9i8QHQFGCX/LuqNCS4guM56hEsjR8osvkMJejH5VUWC3
6/simQLQ6I2AdrbKmUk5A3HqK12U8mW5OQ1OJsO3I7yhGrIlnhFMWmlQq+ffUcdT
NvII0Xc0aT/t0t8NZW8n+Jv0q+vyb7PopMRbSiMHA2CU05yab5ADBcYJuNIVVpMl
bIsrQny57LuD44tfazPv377eIAeLAbRasmpOrIQHNQder1T36N4agsK5AO0+BCEm
qWUiQ0nBtIX5V60WImlvLxVTo7+k6Df7y5cg89Tj2lSgZuNgsb+YVUm7JCiON/8K
ep5SXpsRdJKAidkOnzE8Y0Z+NoGARUgtZfMY8v6thV5unIf307sCnUgo5ihKITuH
/Scz1vHq1iG3O93PEm7azO2GR4WFrNEXnqEXCbzP5YONm95kHEr6i/DpqgWbTlph
CK2GsgQSrEmrLCe4HsheEU76qOUte+07UDFgspmxwJX7dqY2bXOO7brI5spZwIsM
bPF/3a5x13uE+XJcI/zvY+SBOn25z/Pf2LC2KGHOB1zK7nkY/+m5GPIO/h6CgrgQ
vaKm1E75wnIZkLK9r8/6wBdZ1l4ZH1P9Q0avILWtt4dpua+RHLIRAp6IZ6NKq8kM
d+XIURbdP9dGAO4N1TX+SyF3n/+elePxYPhvcp/MrDmUdymJWIqaxdQIRUHWp8RO
CobUEWvCV7vZPY0lroey6vR+sSBYRjAgnyMNm0dF/Bush0Ia0+LYs/iqCwFgAuLg
Z/gNJ+gCV7z1PGz6n6VAK0wXLmSymLKuUk/1QZvbJKoVD+hMXwCp854DZvbZnPiH
Nb7ahudyAHXo/tT0eewtacql37EWLCwBuJnBj8Ce61L69d37fg7zq2+k55pTwWr2
vHCLeR6q0M9rV75sOkN/7Y7zIKDY56x1un/ikWsrsZWVAKDq1GWIwFJs26Hgntrh
EpjZR5fTV5RpS24cB7aRXeDyn2YYdubUyZqX9mft0kmIOjjJEOe/9rlb3LuCM1P0
cgW8/0nIY0ZxHIgMDs8Y2Py2tIHMCV0QjyBvSm3uP7kPXwayYAkbGESg4kUrFdpJ
IfP11YjNHH58/EGxgU5WgOJp3GY2GIj3vU3vgasHsiUrNQEeGyhI22n6j1HCKVj4
yoOFxz3vsV8wK/wNGUJ8uQSkKWp2iP2h/InN7jClNT52481AYS486k8Ccbm8xzYW
HG79c9264XUYOa8NA4pYV7SlgGQ3aOOUo/Gf6HgYf3nJfXzSQ6LvgvyFtjgnTrRZ
9o4N1874l68TJj0GnrszGPVSx76xKaGXWeINYsRmeZYNOjRfGAYFh5hfH6ulh7cw
3mUP9QNGcVaJOL2IzF+ZTLG7dW+GRVHLZKcNUOeC58Z86sejdfK/38NM10oIY05l
fpsdJXOgMdzZ2vagKlrgUGXeKsih33b5H3qf2h6O59bmv3010o4rCPk+YgHXbSir
VfZ3NAuEEWjzUTstUSSEAi2HunNA5/Ud4ntRM4Sh/mWqucN7Co3ubBDQ04sGjwt6
JB3DysvNGhDSbyoepKVZkLD5qRV5yovMFoBkat///skJAw+1yjV1IwaRKsvMhEng
hNWWLId1gN5w2BBsJL0GC5gLRoJ7l0Z0r2WzDJkwemJi3dJq+8lky99Ut4y2LtU3
vngi/4cQy/KYgC0ihIiLvLkNCKNlmLRt3mpMzAkeMrvNP7S2hFXmTHS+uzDkz4AS
opv2ShplTQ9H+NGfLzH6iGLmld0Z2dZU2nvzfXLPoOPkwynNPgR+0Oc1dawZmnwd
Y/+ZxeU5t0AS78rpZuomsr5dIouPXwrXkeF9Dua20vp5Yk0PaHFNwg8Q9Oejjsfy
gsJL9FXa8KKSlvgurbrHV1jrGFmKFlBwWz5c250802GQp/Ipa1Rga5f0Vj8Stf98
qTPG7DRFv46eRDWdfLIREzxkZTC7kySG5WXzAEX1kILuhN394azxN6KUs4+X8se/
HjpAvbiCfT4//UkT2WHBkN6cpH9gY5t7aQSvANIOgzHD2CDwBvXrYsIfr9xy/Ue4
EWh8JhXo/G2cfP2zj7LHxqNMesTqpiRIv2FKMWR/t4WlaS94xuyOBwCWuCdKcT+9
EMtNACkvq44wDb4cG8SDjYsn6eRwJRxzJI9B8/GCb44FbGiO3Er8neRF6aFyP/Pm
l/rBnXzI5ev0v0ep+dfz9u1Hxto8hGSZDtUhuKomu6jak2aJrnCBF1ycRkX93FEk
37IBJsEzXy5d4PSqYFVneLxRQ+kcocqeVdyBfdZAYNeDKtRN9idNWSbfWwKNcMoS
h4O7AG4I7UAnY1ZNT8K9tcsmf+A6j77IqH9Er1JXp+vYBSuXEsEhqCwoz8PwDrJs
eqLDAFS/kp9ZFO1oOpVmwqWlyD1PqPz+99vDrTVZEFNXBzOnjYCaKw3CERiVRwLZ
hgcCDelA6dH6H+tL4QBo91F+tqgzW8LNMVbOdC/3D1Sq1yYwremEjM35zTepd4oE
5nb4C20U1tI4VfhIKhP5dScXPsriY8T66oY78055tOcj+zZeJ7Nx+X8JYHux+cnC
j9cFRQvIkid+ccBlIR9hPQwFFF9iwIm/TpJ0Vqhx0T7G91AuAWBbxVQyfu864Q7z
qjCOoEhQdCoAP34ddr8MkLRNVdL91KKtlhclPz+EdRHS1zESYqU2L4un1LzR+sU/
+5FaPMXhzFds7fOB5HAATRAPbbwW/6qmzWJ6ku9/nJpOHn9Qa3IzCe55Tt8UONHO
JXvZb8ZFOSXVPZKvyswWzKgr5zmSEioLfIDcjhEhbnrcI8yoPGwhbXDIpbTCH5zY
HTWPARC29M+RDptRL/kKymJX17pnDCYebMY+QjMy5YPMOdF/5tX431A/YLJxBvbV
Hh5j4sXYPiWu7GpypeiAdgp/JYN7i1nJYZLrId2S3gqIiWYzzwGmtPIj+qlFc6u3
nMvU/u5VRGDv+evagWME8IBNFIQOmMR+ktO0Kw4ids7KNZYfVmolwTrpZroUk55d
Lx8DHA7iC6Nk9hbDzhkNVyO1rGSDDClNhbVN/wotgm/ynyKH/9Y3KyP9bcRNGyZi
VW4SBx0lG38cUX0CgmloD9pRfNh3uA7BZrBuUqFJJ/gK7VJFelKBxVn6cM1FGY+t
lnS9VrxLS+VdwGgJL29zsLRZ2L2b55nGybA4OW/4wQGXTFWrc/9cdzmhl26b9nXN
TRfDKz7GLi7pAzTCfWdjymzZ0n50IaSHQ9cVJQZhWtMT/TCB7a27+Nu2iNiBHz8Z
MbP0c8H8i25o6GrBCBtwd2bLnErm5E4JH2JNf+mZYyhGZBGHQfPEDLrf8BYGB6kJ
zQ/A1ivmC8Y9lIkVhn1OXICqm0dh7V1eKrNJuPzGWq7MKdfjosXIP5QJStCemj/4
ziUx+vjUfoopCN4tMv8gUErlsLXjUUAHCrhr8yYIu/W3JuLmZapXd3VlStVDWGKY
Jj54DsHeIo75os7laxf5JV2BYmTYoFlMgQm63z5UkzPVpuGVHOgChvYfaYm7PS1F
MBx+hvxth2m7kfAdDK3kGXoCAg41/cGa1AQwgWxGINT6oDX0s/IENoR+0DnRNgyg
LgRp8dss0xGmSV949Sl30JAQELhzYaY8BRhG4ZzrRPQMbWPwwDoXAHpCUVyAhitd
WV9fBPZESrGRJATXrrjKXAg2cvh162V7aymLUeZlPGGsRvVhXn0DIUYEgVtdFB+f
UlRJtz3KDOemE/ErgvOT/YWdbX0HsJlbR8BqgYF+VWjeCh0gyRvfXloskeXE/zmb
UzZ6P58GKca/+KdSF/tt6MIBE511+86lWIUhLw5Ypd7AfgEa4mmhY+ey/eiZmHWS
JAqVGAU3FkxhXe0hqYo3rgk/ZRuZrv+tpBalDhowfC2u9RI9Alshf8U7G4E3o3uN
dpfBiBVvPwOsz81ulH8pvUu4c15m8YYgHJbGohefoHve4z6Jqc04xJexZJUOFd7k
ZaHTXXdAbR3pCGjJl3ClCijCk2MaWTC1i5wvZ867uFfBmj2k1WJm6SxCm83mFFk2
7t/ovx2BddJf8grM7uFbPjEz0dKwAn1Hm9lUR9YthIWdeq+A5UK9dbRqPt9nXaqO
RQSUJ9n9IysGc9PEtnPJX7YU1+dTt/42oL8xa0lxy+RtZ9/3KKq82PYsXiVepm0V
EJZhhaUogzI6kTg68R+ex/7a/RABFXp/+xP7C1pB5qn1TIoXuAbQuTaJCe/VWol2
zhq7ANgCKrr4hHmMkaXnm/J6XGYlmtwnLm+pWqzAsdz5+6Ja2u1/Q/8zAOCnPcah
dtEprnOgRPNE8vX8VdY80puwwMhk/FDS5oQyaFTde2sMC1/fhdnuf8eztby2+Foa
tAfi83qEA9rm1uFy6/60/b2oO5/u+qAAzRyPwxMlZLebzvJCQ8llNlJmiH5YG50B
6aQaY+5EGuBx6nOW8ENQCCM4bav7apmQjXKMh1qRRerVGYVSmLobsypuDwMKPwHg
z/NCSjwOhFEAUBjafIaIuIfi4Z/GBwWtJ6NZNQAnlwPk8yhorTGW1Omdf7kAkzNg
SZ9RLJsogzi3EdKtlUzPKeeJmJV3EtHHCTeFtYQINJWS5Y/9v5TW2du09gcwhMo7
tXLI6gHMfXaVKtlpwHnYLoxWaxvxa1ubi6D/OryUiFH+c/gdw3qJLmFJsk29eZF/
k6kr5Bl0xc4NInMrlrKAy86fSn4DT+Z+OUfPfQikeGPoLSkJM9thZAFqMCM9IGkL
72vwXI2i6QxfPIC6Hak3rt5B8XkHqFyS1+WYccGa0Yy00WiG2LnCjLIAFyvM6AC+
mabUXwKMK9BvjGIzZNqZiVjkX3mvjAssgXCY7jnRqm3p98/TtRKlAuMIjvlEt5Vz
uNFPA7/ApdGDli8gznpKCv/qH8nvWYvWvXIOKmVULNl9VfwvZzE1AXy/7qdW+azi
/u4MkyikRbdA+yoKdMr5shMlGI/DksImqKJVTMVCohy6yv0PfaTMRMryr0FbndFA
OjK776UKeKTLBRLtmUrZOnfWDDriYN0VtAcX/i4W8V62Elvz1lNltrDZm730VvNt
WEQSAlg+E/4I4IrnSBAPpD0YGZX0fkqfRs5b5ot+86vbOoowj/pIm5upmHcdDuKY
i+luCGO338pjMNCnLg9UwKMESaXi1ZjK8bindQnJNDkRH/oVIrpjskfaCLr5vZfJ
/HGDrYmdalohpKZnKIit9UnzhBvJHhv2Y/BmBKwmlbRc4di+lFavvarUOLkO/GMN
tAVLlkOyUcR9oqAroKmfEdjIXDTcxjjU/wCwLF9VdtSozEULjY7Cgbs3E3wxZ70A
JjwLaiF3GpWRLYSlMEcuMTXy1D4VcEXf5oqYDP4SX/ixFO4CBfufXpBNtL1kH0Ml
fTv4qAglTwFeooZ0Xnkt576e4gD3NPSrZPQ3QK0y7q42tA7NlLulsj2QuVy5ZO7k
UNk7UDwXlSbwk9/04SL3VNQq+JoDNz9XQaGZ8cd41s85g8XQEQUXjE04TxdpoF2p
7Cl5kHKLYehoaTIBtBgFblLjc9VjEiON30yCywqLdDtJPyJm3vPv2Nuavc34qaJj
NodtoGjTyIKmUvo3rXsG8bG6o6MFIZBrp+xd85EwFi1yxC245BdSqIAAjXlRe39F
H3HPWlO35jvV7GFnOwEGhXaTBgG75RfjXvqd0L+rwlwcarUYWJbwRyk8l3sAjIv8
h3u/9hH0ttVxQUTcgSd5HceAJnUyYSv+ykbjlp6Z/r0gdeo0Pw0lWRBT4Tk9F4R5
7FXmdd0d9nkQaFpEeMZrruaO2ml5qSzZm6sMCow7w87mrtHFrWLke5U3MLRNeO5v
Qlk1FhiJEYhLj2S3ttFKJVMj2U/vCjF4RCHD3pgxn4B5M+6/g4CNSvDcxcw9YtRy
nibp6N8ufxmHMLqa0Uqa/m2p8a7qO08m39JQtXgkxIyP3wqOyTQfzzV5Gu+NekUY
kprWhpe3HL2mF6YEHN9aepT2QmXDbLgTfA2E7WMjzwqm5Chi8wBCEzQ1AcsyIsC1
v6xu88boCYWt5gFFHk1OkD2YEldlGAQPhPyDC9IptLLeCMz+P6vN0hMloIVDYOnJ
XOcNOYpqei4QnNIWUKyHrgd0iOS94XaJNZhZ5tUnxnVXTVhCltjr4Lw4GfBxe1ST
zVgqaGYsknMMknXY4JD/JYFgXG3WsvjhVrKMbaKIDy/6MIp/+thliqCtcpIlI6wr
zx/w0RBm4/JHvRH3dQFuc9U7Z+T2QIl7MUYk9VwLyl3my04KfJasTqIKDGavdK1w
YbEVsTKD+E6Z84lJfH8pws/CmZzjC3DwKOEOTjFZfMgRss9Rvwa1jw/DcwIW2jIH
etHuRlfhNA+wvKNsjCFXnJyIE1843rRdFnz6tGCsCCu8shiZe0mo2QZ0yY4XL7Cu
GrcH7jDb60NG6wagnl2xrtE6k9ThLdNldTifYJLquf0hBOXok7toUBAkZyOTCo19
xEoSJfsU5y8sdoizQQU3TKvmYd9DwRzHc7z18n4OoXaBn+TG7TsqArS7M1Ua76dV
kGf79oCkZhe6GPpfEWfTUQBbK2xT4aJ88o94I9Rz7Bl+GWSsygzsGKC4HThCpz1q
fa22zjmihmr1Y4RkrebOPIf/wG+fb1Rq2s0TpEpDl7QJ5tKMGBK5FT0gepLYth/Q
Kq6G3IjhVQ5z19x8kofvtyUz9qJjF1wOF7iKo2gJJ5318rMhUGeTQjHVdVTUPqX4
19bh4RU8+f81p8iCL8HPY5CtPodAeMJfmQi2KrxZOXqoDjnjZLi5OCn3hRNqPePU
RJmRyc1t3YWXGaFfkNXnCo+x+6Vph6ccVnhOJFacGnECZVTMdBkrBbBIYNoaI5my
8ylyyY08VvO0qeDsKDnWPKPcymgH3jVMpmWLKaevwKTPJ11MZfLda9wHAK5BIpdP
WFEx0ZW+0W5cIeUjp+HbH7O69mWUeBg3xkGTM1nb/Fc9b1B5YywYJJsdyP09II3F
t3hjz4FJkfcyPYNl1xfofVj1HFGpEH+SLgxo0BYxKLmQtZiFPoXMQ+XNb9SCVBQv
WzhsDmB2K4Cpb/ythRPUJNSy4p9/pcdpbS81Hu7T6uDpAewicBaomgGOnKD4fNqU
qArucZT1cOV84nBTecgfoZuWhPCv1J3U9KvWYI7xsjnu4hXQD4GBu5gbZZqNylDU
YQMYmCTzDkG6Am0xWbgoujLs3gKNlgyW55rdrKxBrP5WKEt8aEPTvi9RmIOqhZrr
aVq7ZZ2+HEERSDLbLjJjj98ULpzIV3WQOohgzrVdzbz3Hq2QW6kitQ2AgVV2N8oR
mhTEFsgcYdRt3/yxrJVX1Fz7KdUu0gcBcySJl9S04NC+jXC6tkh10LGT771MNCUb
e+vDAI1sLauIn8foAsUgvOUfe9iMu6g1Z+J1yiMF6yxBLdX5dNNXtHCQAo9MyevA
AAvZkuXAhu4ORT0TVrykietadlUxio9+tPp+Ek4nTBPm+Nd8lJPNpzpCC0CKhwkx
9Nf9AZ35V8GIUpKRxEvJs0Td15hwrgUYT7lPNCprUJl9lj1fek7s3co2bsyAZoPq
TZfVdfo/UADsz4rLjRr8xCt/NbdnrNS6mDAGseAr0KjHl9tT78WiRxFP3Oz6wzmm
hp179VWpbm3CJ95H+m5vomzGw0gxxVz1jkzzmBWimwKGDXpU+ORJnF5Gg7eB/Ti/
E9RRmLCieCar7QQ9e2TcWxZiRXoHF5Kr3Zh6RBSD1C/clo7hfGWGxCCxoEnMAVse
Z+3iZS4O5wpaIvKGJWECNKoyF/55WSOTeU91DDNFky9p/DoVa2c8W7iQBdrs/zBh
muIchtXkQbqZDdbl9u8epaAiVZU/D0TlZbjgk32h5qxmgxPJlnEUa/D0BsYiAoX6
GXag9dW1zBV7GKIpF9qz4xnvOy9m1WQA7k66480GjyrxH4uDHCsq5TmZ3q71ehnX
L9uw54OrtFxtqrOBiZV4spoWLfoZiVRgyb3XPSuT4Rafc3K7+5rvZ758j8sOPVGM
wVYV7HdNmYV0wvkIfnJTcnvJiZYC5Pe7ew6mokoFicxU+2Q5ZDQo9ICpykTP4nUW
zq3kpAa1v2wiFOL2G0t52aKI0IGP2gEOQ8R4hlNcJQ1eRva5nkO6IDy65qAtPIvH
CyVib1F5tArJyZUMRHPNRRQDTvvLpCk5bj1PpxNpq9uOzUhurnCzk00y8AfThu7/
8YrVx2n/iaE8eM2PXe4WoskDNHjxc05yeTVFAUTVbHLWPxBAiGn6+R2c1V4kZkXn
gyINlhO9FiomhMuLwNVcLdsla02j/oV4FDwc8gaJoA0SVlaTWGfiIa8f0VrUlh9U
8QsdTZSZNNCiSHi5QtlGJBOSY65seaq48ZgKs2yecRkj1aobb806WY0XMQZb3txc
8FB0XXkfeFIjy8a8mO7JzAMRuRnuqakfCUPozN7/WDy+5nwjMaN7ZS2blde71vGS
el5fsU8kWplzXCMdV2HS3U+w0PB2lDObtG9M7egCaMBI/o2Lw6ltGkwcBloh8fyq
Z93K/xCuKErh5Xr59Wlvpy2sLL/t4kHg/i0mQXVcJZiz2hphIIDob4OqKriWREwf
PDZNHwWU2b1Aha/Qjlnyjpw7Ws4IBHj2v+1qnlDYb6aM9xnGhp1jagSm9UQEb2Gx
EwGmH9S4mZ4vPCUyAhUNX1FS3B0BRpwE/oooThFxnQTxKhAgPMLiwjEO1EI92noy
Uvb4mOPYHmU9Xhmw5V60+DHzQ1aQs3JmmrQgx7LrrYs0xsWxmcZ+4SyOwr8HGSqC
zGPDTmvrorgyWPHhL2EhEY++G6b63ar+RnXn2m7gFEj48R6aoxVoFpva1WVCJk25
5qpc492dHcZ2JNM7+uPLlLibWkWSnpmRlBgtXqPiXkoBBglsYuPL7CA3AuYbjvNo
o1+zc5BS6YUtESodCyoW+2Px7CN3jm4wS9LKsiShzzwV7NtGcdGsOzwITxwngWvu
V0XEOl9/eUkNh6q92nSuilQQ7SOj2DuYayyS7YwDd1UR6IG8NuRB0+2KELHsG/8v
ZAJbgg7Y46OkiLvmcUUI9jVXoKyM8oK4PUGNlWUYoN6zd1IGn/N747+nCoU622Ul
kgM5aPX1bGzSN4kremPAf+EJJ4ON/EEtYPiruMXubm9EKZ7zTa7Rz2OyvaZGkR+2
XSUNjddYLCXYRFJ2DpffuxYWP8Qc5Ezyy7zOKifEVwGtRJbsYA1G90BR61dVNUS4
lrMHZC8hriYPMirErO8+WGRXCnOcA9+cqFEhLjiwMX1QXIIZNWKRTjqaNe08W5Bb
gww3+vE3drf28Vt4ju27J6QRWJov63w4Z/MCS28UZegW16mJ6tnsVbvMzd8Wg+CF
XJfjQb8KTIvAANUeFr3wGpG/Fi0UuyrswYw1P9ax+PhnsYeuk8KWm/wJMoHeaYnu
apbtl8ZAxGzx4pxSDJ9vMGEJs52u8IyFnG4pQkV7yRHGOCvo/vQL+HuqgrL530FS
rPMq5mQJX7NfjjlTjUyafP6w99RhYJMVbHG4UakGZQjyuzO1WhLtmIIHnkldNu4e
9M4zC/uDDuQjk5EdYE99z7Iup6721n7vNDLntptdLBzEDM+wxczAzTFEYJcTdI1H
khBro37c6nYv9VQb4CG5Bx4gkLcCVxsxVUOTDTza7WOE+KOlPewGnhgD6vjYjcdG
zn45frr8rDOrC1iaSRZfszpMJIcUwpmdem49kIcUzroenZu7F1do9SCSHq0wilo4
oU6PwRai7xck7VeJ2T82xgFf11I4MsiqbCj1OLiWEK/qDpeUROQDyrY6CEFwSye8
P4N1VFDhjJH08LJ+ar1iIFQm1+K9MnvSjHKy//G757Vzp0XdB3keWVZAG5TZpmxa
nD5/Tqjkn3h8rCM4MPH/bGK7bveMiPg428bVadzDxFS6LDxpSUwv5YuksxxiGsXo
665YHU1BGqCUgloYBVr0LbF30Z1xjuonMH2x3xAZ01Aj55EFRi+9aKab76FozvNw
Dzi9S0oReejaZiHwW+/WRU+czijbpdFX5Yz2XvZIoDn5BSlOMvuVSrNtxgwKa3JX
KcTgQzUDzmJNOME5A0sodgQ9ItJPIBKxNpnvOL1QkSIDQGEiwVFpYvAXL+zFPS7t
RZlFHLwh5N0/T3LNC3Ko8WYwD0Bj/LTEvzdM9gvDm36iu14KLWbJBLFNOv5dkSwW
C2WVRIcYVQyXqKuT48uzTLOmnECufqkaP8JmExdwuXwbMl3EI2DARBCsI6aLEomh
w2wXONcG+yaPO+w+5/Syze2SKQ84KvWUBFBuCg6+ycmtpUFK2IlnFybJQKzQLopi
/DA1la+fTwUuJwRGm8ASrHCGHkXNhEtMi8WaCUeqbpvRNH83aYirL/pNn6VAP6Au
GoYlTU6/MVkTcuqWuXiaUXkktgl+VEdUoHRxxiMiDWQmqzZNK3UkNkXM7tNiXhfe
u+xUWb9PNmRVT18t2LM6NceuotQR3lYBzwpdxy3j6vk6yXHU4hRC8Uu7ucc8IXcm
suymI2UnGWWuc1oNczEmjLRWWQURpC68mXe8G/NB7zfbspyeHmdpTvlcV7hw5FwJ
dTy7T7i+YxG3yOLCR2ZUOu86PbdKK3Xzmuxh6EyI1zZdSxJHq9m51ASI32b6Q43a
vPDpd3bpe+NaqEBeDJtz9ONYl/RR6T+63IdqTp8iG9CqkFRwlDCvFQ/8NQm2EU7L
Bq3JaR9/XTnaYFCoAIol+Mp0bgq8cAff1DVfy6vd3GWDqppLLasSUhdnlNin75ku
7eYgBt15T/MNuYhPhLL/W2z/CnF7+CUh8WZXbZBU7WOoJBaQ6gKWCIjrjzY6+/+C
L/LyQ3QKbNtTHBRpAl6Od7bCxggkan8TajvaBqOxOGoQzlBeuqVqBo+03pgN7yK7
oPBXzFrAjuZPLsUrfTZCif9YX2Arky9THuHmB9Zu6EN2diBlJs5PqwYIoCjdfob5
mUkyOItq6x+y2blhXTQBo8T7i0lz2aY9hukIWHrPQLbX7UxnpWe7ct7+l5oSUOF0
8FyVu2/vWpwh8/KMiIGioJ0rP14dpce6kI6fKTiGH84GQWwgSE6zdsxRJMKNsb+Q
hzNcjyDF06I8QaIuL0wIjItIqZHeKzDVir8Y2fbPgwVgImpj6ld01SNypitHxRpV
8BiTzYsPupEH8U+5FeZl2G0wHWVo9fR6bWbMxtq4L6EcbztE2mo/6S8IuMpzNfOE
hmbb6uEy8vOMP6gGtNjto73uMKx+2ZB/X2KRV+NEQ4FDkP6BnpEaa5i6o4TawawT
/sLBiHevhHMFjDfEaKe6NHN6ZlcPeUe9nZWZA1WD7UlnNOPR0sPIwGlpbIMW8fWB
x25uu2q5JMD1pygPTG9BCe9ynlqY/LDfx8+l8dEUv7aZ3bDxW/otfpBgqkSZmZZ6
Pna91QTy1dR+Gkfjrfz/QXrRwdF/FZJBiWZfzpeStvqXKr3WGWmS2IB1SNvLGzd6
14eQ3AgL9pzCezSlT0kC9/giQhnZmQx74BI2GvxIP87ADLrrqKRIPtX+/tQIKQ+L
1Z/vEw2rKy+QLCAL6G2aYBQw6GUGjk47PI8qHdHt3DEYb9adCPnKHiiQ2MB1cPN0
tYB2s3N4c87LcQd9A/iHI5HWLCpP6Xp/deaIgM2SE954Erqom2xs+CnjqSayf72Y
g7FQo+ZhoPDDNi0daSZdVQKbljjdkvke5thlbFyV8aaL4f90OpkGiIdfvmTYYMvC
fRjdbOvRXST2l6GkeNXVln1sRINs3GcfcJ15Yb1kDOK4LP6pbsV0MulFdsRpiYXG
vEp6Zo6QftJG09xJrc/Syggl0veuByrloWdLGqNxUKi8zu1G9M/OO+mv0aj2v1WB
OBNUAZ+5xOpuhPkkOWdEwQ6MPefJXrVtMXcXZl3ZRyCj+fVJxB2QMmpMgLKwdT4P
OPseNK+vtNwqwvF39fFeuYEpuy87rFXP9yhvQ6J6xdxmjlh6OxCmKJ8Utk+rQNID
SZwYDeKr1bHNrRuqebjFrixmiXmxA+1nZvdr3X6wZldRHIDzmuHkl1mjBCN0zASF
AsuaYBJ8kzVMnLVTW8284lPTYIz8NE5Oom7+Cfhhym5jgMnq1bJNdxdKBhJsST0P
PzO9Cr16SIYmoHSg4jk4H0d/gXhw9Y03K7XPIw+/EvBipmEh0yAdnym0LXGR9bOO
i/gH1DpJoDesjGh4BIFdDuN2HSMR8wI0ACaS8E8XqReEgk6HVWAR3gra1QX1pa//
MQWkfL0hHnCh63O70GYK+tNKfMPA8qxHnlTkm7XZws8NDjtMIT5Wk9hjSct5x241
9cFvZFPNRvwlsG8TBXlSgV+aByaRPi/qQr65fkcKtPeJu6YzUmnOidKvc9yCL1dl
fP3wevq9KHVzddaHi2NuoHFlPMXvQLaW3e2Sq6nNQerlcuyVoYOMDeZzfhksqCr+
5lTqY1h9UIFpO7GDK7JeKQIG1FGJv91oFpV/TXT5+Hy77xgQL3haK2HjspI9m1EJ
4HjjkTOWn9EuhvLu0PutPWJkJu5u1JlKbpTdVaBK1EG1BPRcNAiAZ9NY3R9pTpn3
N6XlK7nIyKYpbX9IcQBOpRISQxwOzeGwX5okhFh7NeshKcfzHp+H7Mm6aLmDH2IW
vjvDAzOB3C0xFeCOPtNVlJS5J5fVg1zKBL6GkQLcQ6gCuMdBVeXFiFBuh6Has3Dx
0QweUllgN/79G9ZdpsaSkeqicXMFiQiR+5gaKl11RlkBEjuKnMWi0l9Xauw4BhDP
jlsYelRxSEQVKj1ilLIdmgz8b3A8RtlZWMTPBBITs6ddphci1B+JIvVtrkcuIpu5
togHdpvmqsUZ3k3qDbjkbK5am8+BbXneTs645/iGXXr19YwwJGacpI4BHHpFrEWc
dMhc5GD+hQs3ZWGm91kURsLi3LJbwx41/YJ60WyoyGPHCmCqQ7Fl5p3fHsTO1EVW
nfye/glDDYfIx8Aq/OU13a4kagOQo7RaJwKSi46CvcGHaAAElI3I28JOGbacmd5G
ENipk3WI1ovUWaGaJJoVda4uiWNQAPRtreZdDPHvwPpTAnBkSOc6IrDXxf/0oEQ1
+XprCNgtg6oZXdWc6D5mKYooENp1cyj7DxCarqACEeX/PJ5qRVWoaEk67UcJ7r9+
BKy3XSAw6dsPT0T5Nz6uoRS/nRBw8Ryi1qgOaHHAyAaSN6tau1oGRXe0G+rwittV
wv5XXJ7jPrNtiZEFsAg+pfBMxVqfhUlNVUAsdwii5wNWnLkit7FSl1ikmvnrJ6vL
FJzMzzbW9Woy9xC6mwoI7Kx/Oa25iW8N6fYuvcZN8EHcXowHUEokBDRryNqx0cn+
47+hfc7BR8O9CAP8fOKICH78AneBamuIIPxP2ilOg7+Ks9yjnPk4Y2HZwf7Tb5w1
xxNUokeGN8Pjo0OUHARM3dqapvln671Ttn7VaAieU+rjmKEqQ9cTMR6CE3sTnilF
jBTgjxxFXvdzNwN/dI1PW2njG7LKlehI2dQEFitCAQKLQDplyv3dNo9uWKW23FOL
nqhy0vsBm7aHJjzpf7gGcwcAWcqsBwiRFXcROEPT7aq98ixZ5kZylAclpsh8M7m2
XIwb/scwfbTG0fY2QOaAXwfynvlfG29wDwQOkuchCKolT3yOfyVbREpFLoH8po55
vZiIWLlhYR8lggM1OslVObwOhpXWxMyJ9aGQckvWLkSmkT3TiqAnu/xKIv2g2ZKG
Xkke1dV7qzdek2fx1MJ+ZXrf6yB4sUCSCalwaUPtLIoOOijYtJAS4AsvZ0kf/4tm
zoGnqwCZRQLOEzaaERRf50t51i52+QKQgEdmF4dXFf6m6rn/C1LM6IHggdJJU1BK
dyFbhUKBYFGNzEorhVU2W9Evo4+WTq4wwItL927xCHZnC4NymktmKIPqHiDd0Axu
FM2YZjDtL6MuWZ4ROSWaxS9cEQZP9z57iuJ0IOcwS57hRDGskgDEWoH2ccfaD067
07D1bKjdmPqlowhq6d+uwx2RSAoncSfLJ7A6S4tgWpawzOKQYJwUSN/PEsIRZh0s
7gcPAvq3D5AQZv1GE0VqAQmQOmxmImnjOg97uzL7/7Xg2iAGYE5Fiy6lBgb7Bxsq
rENwweb1+pMbWNu/idr7daRLDlsIIvSCUWbC9G2k9IZlro/5oZVzTpJ4HX1B2kGf
3Tq5ArjES7zrq8z8jkoqHKo6qyl8P/n72OuD67Y9qpR+X8JVIGnt1Ws81Gk/61Ub
6pmIT0b49VItRa9lPq18SwNeDUZIC3l4xMkdKSf7zxOqzS0XBG1FEozHB3sY54gt
qLSpWy86ftYbD9HAUU1IDmMIICkd9BMUYoOzsodDPUPEiZJ3bc46K3Hiuax4U0oJ
5jSxJT12GwofxpkE9Q7od7LJHvTwiyrVYRUmjhwU/n+wlHh5UiAFep2tzTX5UEGy
DJq8V8T1jZ736tquzxQpxaG3gnsi4j1k9GmQfRjTdz7D/BdEvgsQEGm5UtaJFbP8
9Byhs9v7V+BBo+EBwjMxoMEf6EvkIOiWw24tMAEKRQ22rHPmWBeBYaTcBGLgHI9X
059wNO/Gqsao2WYjZz05chMsElssAatry+xB9WI57XwJ8nKQeVtFIdyJ2DPAoczS
Q+EgxG3OfkQU4hxgFEdH6vwE79USCsoemauqaCJloO/cDkq46vSSTqoATKUPVN4U
YhmH0fYyfEjOJr5mRmlG9fPAo54NECl7tgZvymu5+6h9VFT2tPgzdaPnHa5x205C
uAZcpmI4P3OvIpw8kKgdXxEsj7yq1LSSWKirUdZ9+SiLJrGP7DkAp8ozwbBanacT
gYd7nNMh7E1ynCTInwBldM7SVM+8KO1J4gOyGIHVkiMZXpcRl/xFLPC4+dxtBDN/
tHde+ybdHfJp0LGUBukSOL6M55j2yweuKW0iLT7JuMc0iW3UMUhvdk1/2OJL0qfL
nEPbqH+I7MFr1Xh6hU4Vcl05OW1Qi6dx/v0eaiq1dSBhp+yx8df+d4TA6lt+9yeU
lsfFgIOZcp9ljT0iIEPABXkDF5zitqNuM/4HBX5GrcJItbSWZ5XILmyD+9P3oumH
7H3wpUHjZY/XTlbwZA7N4ZOnrVMAECI+kazI3E2th5Sd07mH98EDyVSC3scv7sQJ
oTHbqQq7V2iSqJKra1SiS5at8t8rXXfMbLiKzYMzTlkAaUz3+ghE0iqOPBGgxl/B
lHHLCNXMDqX45lI9NJuZIlHTY+J6RYUdUPeAmROEknQp666Ke0NheOq92Y+do87x
BlH4ogkog0Ufq1g57irmvi9JNmI1sCOirZgtA/WgzhHAkzIj563ph/hw6ru+Un2n
R2DrAGEK98tDGbnRNUT00rw5FknB+/JcTOm9ej0oNhgpzwJ00LvGvgWvmTJSClI4
5cilZJaUX/Fgq5YIaE8Non0bwnSfMlrUY3qxOhhWkYPsBagtJrHu1qwtnfM6FAZ4
d3JgJOTj9FkZVTpf5zXn3BIiREX3MTCJC0QSyMWVOZ9x9apt+ZUldkgyh6Jj/uKj
t4cPoTNA0MbmiJSsGViSfmbZWD4mAoOUrmZEgOJYHGJI90VioihGBc4vtNJmxR5c
nnbvgk5pB6sK0Ny3aTC/rQ4VByioZxUgZToY6lFWiQLwks6pYythrQpirBTXcc/v
Bu6yIHrrN2uMEtUfZnw8r1qIFLdiCRP8fqxBzsYwXWqFy3LhmxCzRSKWv/+U5LXy
qQ/2obeSbfLgODtxCab0OfFV1BhayHHH7fzruSwxZ+SWfflQqXpF609VsY8Nkwz9
rp5de+TajkqDftJ6aFbAejBfuhJZtfHZPc2PCR3doYS9TwjgEgjA9lepgTC/WvUY
o62ZCbr0x1g0JZzr9ArOxgQEBcAWhWpJ+qNASsNF7pUzD1k0Jc0uaIU9Xn1m1PNt
xxMIRqeQCfgsooaHvJy/lj37h/ZxPch3rBOSo9ZOLTmbw4eSYupQH14ZKdhxoUHt
aT9fo1js6E5K3UBOTl+XvikljiOES1TGwD0l4vYQjVRqX+0F2+UpmBPQhNbht95R
6Jlpz41WEsoN2vnMGPApL8F4HzHwM8eiD6TdGW08zNvZegX+4UnZH5cslhMqzA/g
TEhjeta7idqOkPb1GtE5HwQE8anSg+l8QRpTeyMqn6RA/ti7n0blGjafzWZvyt1y
MJxHls1pmM8fs+LVeaI+MDQm50jit3B2JRCeSzDdYcsnvnm8I2kU9qakPuD0ohuf
vcglG9EUCTQTMxymawBkIu3HU0kfY352I1vZ0HstcPBzXmtcqyobeFujRBkTLX0r
Sjk7d6rA41jUbCSv4Xe5Es4iwaQjIfSbdiLlCZCrju9NzIw8qru8x7+MpHwzbSTq
yxaYWcwtLBhIDd96Td2NL6vcuxuArPWS1InewIxRYBGitj1dJedmW8nzT6YQTmfj
4ATTi8aOA+64S1NLYCjUGDWADqt49ZcFkE68NKfux1mc8BlWFe2asySNAmP0WVqx
KrgPukTbRUsDdzyHHtFASA5EJeJ3KptE8uLWoC2zPmGFALdSUH3JD3qTKrbSsQTJ
N+ZCcruhBXodKlS9KRNnQ+7A0nPlzNlz8XJTsGietO4m3pHFtbzMqYJOlKVPgPK+
TlBJ1YeO0cMbQIZJrxlklcFCZosihN0la4pHuhOueyoGwNnpo8MGerDoxet+LpEa
NxRo085kvPI0yzfKcl4o7m8VTeH53TWOnXS9cIAjMfR8ZXhjYWc4BcW0RKnn6ekS
TT0S4yILGKoOGN9Azvi+PEcbwjA0MRa6QivyzYu66QmNj3+6pKUz/HnrFnjGR2yx
jDWsOvPfc6w41PiWU+fJiH/nqRE5NjCEd4hBh8RAiJTFjB/7HkWfrz6zdK7kAx6T
rFY1SB0Pjghud9OJVczkXAjpxf1AhsEKtytSipiCaERqjylnZNi1XctaBzu8sV7t
E1cW2qZ98cOTDfTpIn8SRSmUVt02PQ3iLI10Hz+nyMbCo0WAE03l54fHiF5Bs715
ZovORNRgf2WPgAancWuFdUc5QmScw5nnNmiTZUBLCih/dzgBKTiKJkdzpCxFXtia
yyP+iZqzAq55g1/fdcJwU7PWradlQD8H9q9nEtgHXziHs/EYYJm4QvJLBwgzTCk8
pAzyJR5JHGnySfUR0/IlaQmi6DhzdBAZnPMHU3RZVx7KXEWfYAzh2yUBwdLCX0ce
nK9BVPl3MHPBf48q7hxNh2hSZzuY2PeAIo3Qo2tNh9cipiDi1wp5Zl39ZWSWPQDb
6bB1em3uRcporAq7VavHu6svFtWscgn+DFz1q+oen73GuWrYJdG3Zynw84UjqvY1
dEEZ9XJbOLMapTyLcrMa3FRqtVnJKEzKIG/l51+e9rAionMRYiGbLFUrE9MqvXuG
f/OuprNIiTZ0JorpF8NBiz0ggwtE8G28FJbXDDPs5Kju/uQjVIc0KVm9bhDXTZsN
Qlh/8cTc4eBI7tL+lA9U3rCgrdx3XGSGrbofp0jsGcznq7sSti5Yx7nayaKnJyh9
ufhKwROHvYbnej8J9kOxEImQPzcDoPMbsKFs7lDqKJ3jrtAW3K/m7wx4ytpqm0Ex
n30tNYV4dJmCHJaWaxRIeuFnCQsbIEeD+4RpLmy+cd8EDGMbjTLg1dEhTMdPZCmb
EwdS9yLAUa9wTwfdl9UP7EwUDhooWXugKBZACjNxEJsWucgwCNNPpW/adbSRsJLl
RwPJ2BVaOzVRo0DR0eUustsnLqAr5DnqqVp57tHT4bNoouYUsMe3lRGFPurLEwgg
bUMsk1V9HO+p9Rd5WMC5jx9Pg5GpZ/nBKyDIIR7TwP8CC8BFPWbzieGhMq/mD65C
sX1NjIK9CHHO8cGYzw9IzwIuSyNkQadb1DqOfA8P8mwT/JxRDMoEFHXzpVUfKydB
vDCYPdDMwYMmWJHMNbCK9YzX/GayU4fJaZ3HtndW3KVmkuoNgGcgZ8w40mI7w5sd
eVuyAnWkCApu6aCYEKAMXuPRYWqjvWXsXjTwLUTrmabB7QqXBJWNwiLb03YZfbHB
zYhwg4fYZ4OiHy1KHOEUrDwYt4FZ5caEYQpQjq3BgG06cW7J0f5aq/XX/OmDrx9Y
2tOIRslBFi63uq9GL85yeroUD3CP14dRrmilxt4iOfGMdoMBYmd7aZBLyn44x39Z
ydxFn0JxPosLEfzN8iH0NZFJ6BXRhuw/1OpdHzQhkMNDjLModHO82ooKBcwydO25
rp/QIVIfBDRoeJ3F9Oz8vg==
`protect end_protected