`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4320 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTAYHkqCG+zxoaJdVRpY7F9msVL/YCMoGx023t3FwXRtR
O027Tp7/W6O/0lwwLMcG/3jC8DkGVpcf6PilS7yJbjTOtwz2SQy2tA3nK0b2YF9V
yRfxMZ9DFli/pii1c0CTTcv9CR3z7TkyRtKFWw+ZYipb7uxPs4WhVH65XAEMnd06
S9apLYwmyt1BTFlTyFukx4/8fKVUXVoqMN67a50KF1qsJAFSbtAfxGtx8i1DKSkF
uBsq7k70t8UMjGEQfj5xpvp0fuCIdR3MwFBZpCYJAeljpbSqwN+nQgmeQticKpGH
FtXXMkOWSJPL/cgYhaOeL1g56cbxs7Jvn367R2EzRQ2GqhlKV8mdzAf++uXoopWb
1po32gU88AHXtsRQyPT+BAQCoMrA15Xb5ffl0qKaWwnQ1WrAuSaArG0tgcM2FDjW
m5XMFKdigB+RffJV6LpqN/xnG8vKO6F6a2XN4k2AXbepv0IFRa7IJTx/W5NWPJGz
9ZfPc+HFmEOJdCiUxWnWlhqWC+q6NYF5wyJAcY09FrJiNT/dqDdfqFNRpmU8dols
DULcWDmFvjioaZM/e8+s/iDBTSuoyhPoGpx7REbr/2jnhFMcI0GBCcAkkC6fFxJu
TAYWhwLLVC2/+4No9ISI+BgDLrLQ6sZi8iONlcYRYKn3fy4iASMVh+TyDjT7NUk7
SoSkak1vnEFLNfO5HHu9UkwHgObc7itIUoW7YcJxr3bTSAK7WAOfCa9/79/XJeiP
TqXzqhSZos3hQcC0t+g3bnWc44xRkNCe45H1lPhcbyrYTxczgWzzrmKqyd5q8JV/
JpSCmLDxWVE531s/rtEJGyMLuqR9SVaw/RSqNgkyg4srsZQsj9uTTttqcDXeRnvL
xcEFWlcNJ0Wc8MAJDJwrnfUFwE2YJY7A+G8csJ80Vh5YKEGY7lXHr0EbbVdSIWCM
86BaqUnLFYi0uVX5OiS6upTsWSyP52IMPsfcDawrE7iGPbhYRHnjCA2iHEEGTUpk
Sp1PjzUSvRDqXzuoCnrveXc4y9yvAIaAHkaw2yqTgzMJ4AxIgDyL0SO4DxL/oo1E
a6xlPN7tMmfyRKp2gO8wJMNMxQANLfV7ve62xARDiwzj+hUPewzs7zinkIV5LVsY
Yu5Rsj2bux1fTglBwKmRSYQbV5qgsJfucGnigho4Zn/5l+2ERgqWIKN30JPnPBVs
38PKK/zkk/z17FptrrqBffwR/OQwu7L56ZQ216BBj8z46Vso1jVi1f3kprwcYB0X
w/USbQUU6dfOhHjYd6u3NhDD7Ryn0pVEGGmMZOHV4L2HTQG6k9JrFLvQxgP6wBBA
AnKo2ZKLmNWLYc/H6VwhCo+TBudQPZCYtS0HFYomjXp5Dhz4pF+JFYkC3eZWp4+b
lsA9aynmy3aT491Y4galoK3F/l77XOsJ3aDAQbCVoU9oBsJwIJfVAbXLOK7/EZ+V
ajFxloCkDQVW+8BEtRK1f+WcrXN44olhc/AONaWFPOjFctrYUqRhSsE+ccXiI4Yt
igXG0K7HUJYx0qKhn3ES8geeIdDgmG/Q3CXLh7Jj/Lqk5Sny9EiXjr765NjOoOtr
ZAYj6BU10lPTVL3T/dci55MuG+xCZ4QqGtauYCMflMvsSnmpkN11qpJkeQ8phcwO
I40tHyU+Nxjg0ZZQ68BN4PbqjzcaLduO/2cBVtNw8yAenu7Vey7bpZ/4Oo/FiDcG
iY9EOWX8Vv2HgrydMVcmuFz7TsKmxMf57fatkiS4M/flYDDEzZhebQ/6XFwBvJ3r
cpB9lG5dO7Au+IBBx05DsQ9vtDjGWvtmE/iqGCgvON8xntWu47Pa0X3rkx6QUBi6
ODDxN7GcThCV0Xhwxi5ilRJw0sVGhPPzJxEaR+MMBll4qKUVKgvEVtd4NVWB/jGS
8bCp1vy+SQxkVhiKWaoai1dUYgAju1GJKOeqOShWDw8DXJVzN86Ny/okxCxdLlda
xuUrycJxe4Nom8GgFFAv7CkcQ3PIG6k3+1cO0iM/VL0U38gpepoAlp845RHBnKEK
7qqD/LQmw0I4tY3VnvAg+aBUFKdFN8MtD6emkRjYx2M7M1ckkvZ/WnaOiox/r2O8
6VGvEVjkZ7CittHCADZpj7/NQqVffXRvM7WxRsWm7LwH0iPrRBHqklU/y2J3VNBj
uboarRKTAyt72slmlnJRfWUeEWqqtobITH/5wD7VcXa5ZcVWUCoWGVS6CBsbGYI8
19PaKWckDG++7toMdO9w4ISV4p1hAExT6beeFbgEqEpTLV7ZwegySDkzaqjENoNi
YoMBU5EcMMdRYgGpOJ4rzPx71OI4Jw7AWOCHPbCl53X593Ipti0tDpFXe81aBIS4
2zdWcPUANZeaqZto2kolZTdwYCcxugO4Q9aYwMcKjuvFuiQ2+u1kLSD5awsj0vyz
UczQKq0yB5IXRcAxph4ePYPqYIpFaO6XpSuL3XFt/pnwQFOVhLzP7dpWSRyIXwu+
OpCPGOnS4OJPyy6NFjYx9HJIdOSlAe1STmtHfVFEEFzl4F/quShF+Kjt+Sd3SNGW
asAYH19yzjWrv3WcvR+1dKhcwSm0+fd9SPs2AUhNM0CjeaAMYb+I9N7NjHmj1I3U
8TDSuRVleme/sVtA0bg9DVaL8Qr1OEL4HTo2jK/7BU8+piA7inRlfTnpOLsib+E2
ZD0/pQIe8EX1mDG1VeEAgegL+BCSDL2W3AFwuPZBN4uU26Pptkd/tbn3qMUEbMvI
+bPqupPJw43/a0fR7azhZyf6UXpaz2vqOOZKSVCekXqUZ7IGyTh75fQBE6kpuYsM
BZNDSMwb7n526X5KMjH55e5dIZ/hvGNIPnEXUyX9w6due01t4IjdJixjjEldyXGd
mi7f6cgdjvJ3rZDcWOb5+GZiX7dePoxM0HUr7LfDK6V0FPmXdp2zg2IQ4bG72Yej
WfeZfSp0sKfQ2ymreN8qimGazjpCLsduI5GddbBvWfDfAU83SIFOo04QJLcNb8SH
m7GfK9vjxMQdf4oZw1Mlf6P50u/z0jhpU+FximuFurU/pupIhKhNxmYoAgvRaFTn
fYozWtL48uKw92sTUmio0KvRB4nlzudfrQiaK5Ezx0bsigfbakENiqh/DzmOy8nZ
SCj2G8VjNNzPnPuIMo2cJgwyU0DO+MdwhisN8MCXhAqpCtz3dPVdZmaGJwYXMBGu
dzmTaUKhbMvwM5qo/wc2nmYvw7QefRh9MXGL4Mq9bUJBDuXG628/VJny8AfO+nSq
5fnvaeL5W/kzOrRnGiJrUwwFGjuvCJLUcN2FLss0SMd8dbBkL/SglXL1meAWNRsL
sHni5AjRkFyCqjjjFJxyJpEczK25HZ/ctgHOpwZP5vsqtDjNYheFTdHey7QxemIt
GcrKAecRmVTigCuN/aRGfsuFSN/xfukY4imhfOum3BJYA3nlhK8GsVHIMAZQCKly
cFV4nuoeuM8DvbG7RSkBZqkpcdbg194xBXdaTgaSZFeuNyyZ+PJcOIlD/ntkc51Q
20Y8HvIwv4wn5iakGsqYSdo4eOeRJkGRFQkuaSHbHGj2QCdhzzU2fzhR0NVMf3kV
ReWrfFMkc9j8TXcEr6pQqQ3HRgCKsMFYxvpVJuB3ktu+hYqTogZXcXZRLLRHWkCy
o3sAz9jCztTZ+lMrYgVnPXa0y2VZoCCZHtq9NURGsAbi+GoRnAqfcTJ6NKH9MgEw
ogvRVsWKkb90tdsV8MjpVWVdsNfhLAVhVfFukQiJDuAV5ZpasWWJsDwDi9voRE3d
UoKYON2wqHBM8uWuoMkf8a9qLJIgu03/ulH/AONlYdey6QUGLLy0M2UW7FouFOf5
mkirU52Shr4qccyJ/CAkNsw6Ybl73DuwydFJRnGV09Qlt9CXaZxl84ZvrpJdrx6G
fNQFIQ5lX/BLpYEWU/eaalrf7GG1xdDkDYwfH0/+cJa4lSV9s9KBcaVXzwOCM6Sp
2UIE4DxlafDflKhtT4b31YtoUWPIUAROySxM7Nd3v1988PBDnXHJt+RtdUcDWdJf
ju+KvvuQx+ye2rBndMYV6g/TVEVnjDZJY4ixTYimWW5OZyLGUxcot2uq8Md1B/2Q
7OaVdWpRYAo7a+5E1y/xV+tyRogk3mCYUXKlSwGSRJ69xjMk+76OPk3nDuqJmphz
bE5zCrgDuAmQjFUT2+IwX57RfTy6Kzqbki6K3WWEuiWjOJ5dqUzdl3it74kBAB3P
74HhbVRMv0qlq22EqWh8Scs7dEhVVCIUsi0Iu5Me28fjLeh/TGp6v0erVtahk/SE
X0wrM0sh/TbqkiP8lOzwmALTjt4McusPE3kT1PqFUwA5ptjQo0QJvF96W9H6r5Kc
8YB8HbmhMUSTZ/ZHOa+tktrExdLMetbIoJwBC3+5HnUEQzDCmGfaKwRn/9W0fkbJ
UkREE2FuTlzFnEbSkJAsIvMzuyajIUksBrNGI8VeKCphbw4UY7moKXs7Qj81tr6f
VZL84swu5ccfL9TF+YdrC95qwG5mriH4DTXREoroy3ZBw3x6RMib81t6Yv+a/Fon
rZyOmStlVFLr6Lerv1s7p/O5lS7wIT14VWqAwYl77JH22M3PZT7pYmCiYcPszr7q
ukI9dXssfvmYCUo66gRpJo/ROzv1FvtMxpkizrkNryMBbp7oQl5+B4vj3nODlNqg
pgtgBVgFUioKlKbjfO+HYeCGKuBhJL9W/W5POix8UrwIFMlijZk53cqOJjIythrJ
8/4JUW0Taw2myD3Lm7YMr0JZACAbVukL4bDwuiSKOUYJ5c7kewlb/MoHw3Q/sUv8
LtJd1GxVIloFEpb3j6LjimgdfRp+l5N2gXzAn667SSpNkx/6xdOHx/yNd9FKTWmV
WKNRA/jPWfGFCH8rMwMUMSoNtop/q3MskMPo5I7GstCkRTv7i6E3UIzHFNOc/79z
L9618he/NHTVDMh3gJif/PXiuq+uGqYJG/1UQZeLEHuK4MbLf+Fgfq7u50062Z6A
PS9IXAtTyYfbwbTUI/TAcWu0Jk7bmpKMMrZp7M46nEsGvNeomctpLEZ8y8EOcuTo
VTLkcOoxQOjLEsZb2ZBEG8MBPngDJuTWfjhsfqjR5b/RfiAo5c3xVZBbdvJWn0mw
uCwo2xTFcDp7Il3fWop39T6vtHehC4dL996htL4YZ16RochU6J7ioi3/9CEELa2s
bOqOBUzRnI9rwZi2wltT6MKmKbm1RHshpL0ytlZXuntZ0zfC9LkKMGBUAOCe0l2j
BkJFGIp2168GRI2Ee1mVFFnKTP4jted0WkaUtb6pzHYrDo2M54e11NI5CqT766nw
cVc1wD50a7pCB42KGoUBpr5PppdnBv6lYPHvNnKu9LEeyONnv5+CQzWAnLMyd2f6
h4H+9kvI5vpVwTxIQZDUC+60RZJTpQ5mD6GU6rwbv7LNcCxH41RFjieq1y2FmFOG
idse4atQpvG11//YtNYGtBKOyEpMY8QRrEQ5afOWCy7qUgGp3u2RE3tB/ylzz3HY
VTeH61QpfJy22AICb/QhdkccJ4bnwtOI/Wqy0pvL7wXD7H6oO3dc/2UcYDt3n6c4
mHzKWhfCEGVgSnWXTty4hTb+UVzvGWahYmrpzW6D1/lW6aH+aC27/NOnKn2eTK7j
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4320 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
lmOQgIOM5jiJrGbWpsW/8vW1JpbRiFgVbGCdXf//r0/3gW67VDte3ft/qgIEdOtl
jMtvJPzkWK/l/ragtlhlWpp8WWennwbYK6jp1ZV40kBYshQGi8eI13zsKswuGClL
VXFWZSMwmnt3TsYSQt35DSzYziljvefpU+lWeCrcrShcM7d6BOpNuMelgT9CvOaL
POlZ7ZO9gBBrClo0neTBES/Yf9lQVAZtKa5Wp9fi1913Atmg+MjWmRz9Os1ROmcb
RdNAsRNsutfJQpNRWHVHeNm9mKu5FB+DYyrIzPQIaEZ/2+dzpW5oOwffAviq3HnI
InsBTeHFrk53wirftcWwt+bnAc2HGzirTCI69QcnRnJbFoUbU6rhZETTRT5m5jsf
Y8UFbRP9CFromWTI6HP2fBHU1juiyt1pkqALjUGC7qgJLWpVurGH2CZ3kQxJcX4T
rWh+pC4tAS5oIiusayXvsdWnn3kqcDElgQYYBe1oxe+ipbbZIW/RKVF1annnMpZm
3EJCf87Dh8iz9Ye9skCVwK9sfSkZswDz4oOr57axMjLQR2VD2ZpT/RJykc8QDnP1
6r25uxMd3jtQhi4XYW48wyTPkSP0W2Jj1YBkjeRP2E5c3o81AICH57cPWwinPIGe
SbHyFvHi5WNitoC0BSlj1tykmiYQDjM7csA8J1UreuOCOn7EC+iZrQRscHaJBMG2
vemzNqCw3+xFe5Z2HwaLO/TZkGvlfmSvL2pA3fF04x4CC4t3QlDw2MxlBL34qLeo
SqTOvz1joCzodXBuJN1f69ufCms4aWW8mvDSIM7KafJvaIzWI0JlajljOpCYqphL
atemWQOndq1GL41tTKDu0O2I9nQxyfo2LxDBEyIHVv7TdlfrdHIP9Kqdxz1ejbWU
d7+Zzm7JtsPlcpw8dRvUbl+nC0UMvKgd0lAAoqvFwvaidDYGKHsZy2TAErF1e2FC
BZwP/uQ3qeekoWFKg75tm7wKSjbhe/AdNAjgkXksLGpP1c1L509USrJPg3xmqdHH
e8E0MiW3qWyohIZfgMaTIzd7ebw9cB9ZY1EyNDIoazwUriuUNtdMmijjlAEyBIF+
+OqtNgHEEt1jSeV72gE8gb0iWIyAEcPDhmkv2950Z9ZOo8I9/F2/AyScHSYpV3wl
8lC5lKLxvU6zu9e4TzCNnrdXx1lcRae0igXdP3NhivH5VWwC7R1+aSzSfoQPinAX
OWIhilc7eFAhEmy+1ZfpZfFloIRrSOsjresKy7uIW2N+ofFezkX9qEZBf9ujKTWo
Zy4lf+uSERFvITA3vToGjzF6vXwUjAkh/Jw/lmtnx50xMDdl9cM3ISC8QdDZ97J9
WQ/cGiZ4wr0HilxYBGH5Jez0K5TqwnTC75mvGnW6V80k9ipNNYLKHEjS0cWo3KP6
5OOM5TvbVKXe77Fva6+7IxdeKRF5jDS9+kPAh1CZQ/4hypxSI6d4Pg5UA4oexZqd
wohxlkn8D608KYeOHGSulz0yJCLY9YJ33d1AXB8Tvf1gdKQp5qkjx813G8lWT528
5NU4/YMZeI3burycVc6l7Q/URWvvIjisPrWzYnxi6QxJkjhf6QM1TXYinkT7IHHX
e854xtpNxUQ/VZt8FAhQ6mDNbslbiDwZnawF9qWu9Ijazr5b4T3XHe9VIIjOYlu3
faoa/vkzwMllsSoQ4ZEwAeo7/jdQli8h9OChPvdhs/jc0q/fDHfiqrCdpK1+lAzP
ZZn9gpBvjVJq0xImrljAgfZ4HGl4y7Gx9qE9Ppzc7PN0Q8LAOhNkxxZYPwIURvKm
wdRxZMkGXy30/BaKufwVhkoUb64ufkIvu8hqnk7FeJW0ucMMSNL1ZXCPz1AAJofU
okNUoYxWF1TuPX+DRgi4rwqXT9iq+8/ooNrh91Z8cIL3MF0WKhVX7lZD0sM0UQTj
JKogw01EjDk1Im/lyr5OIbbn6FgoD41hRKhRvzsxLueIZxh6Y6DpbQQaITFRT8qW
vu4WuIplOQh6yfUBApWs34fpKOdcYOWZRDZxe984V6imKBZOB6yHDI7IQcleQbY/
hIHxCtTNaJibDZ6qfAmDV5fSS4Z/10lUVp5eoZkK1qLwlgcGNTvsHCNd0n9Y34kG
vF1suQX3S+oB6ToBLSsLaLeSmP7W/sB37P59P6qBgvFHvNeJJZJVhwbcZsn+aHzM
Ja6Ts0p6sAkJtEjLVS0Hk5Vm8/nOHOjEE/HzJ1nxAnnhyfd/VOY8eaSDRLRQwz6Q
rWujQTuzFd7XA3UdZkJ9vJPYiZjCEptrKe69ZSNdZB4xCBhwdyJwvYO9/pg0Lgj7
TLL0/fQzecMVxyAH497ZRBpQxunlx5mzHyJ26VMHIzo5cnsgfUMYPLJ94wextPlR
1RW2EbudkWx6Jdxm2CTuql+d+iDGqdWsATIP7153LHPoRHhd8aRc0Mpe5FUkeCpU
SGLID5zxQ5EgFHPeAqiG148YESz9KQtSvtgFTgHCfjCapViJYpL7bqtKBlY8DRsZ
sbeIRxC8lcI0MsugP8Rhr+6Bni1qvr7uLKdZLYlmKxAPfBDyc6dfMHYMiwjtPt6v
Vvu3ywohS1pQ2sXP/0Z554HKl+lMwFKa43dGSr51UQA0sgSovdOvJvUQpdiJfGD3
80pGBHFU8YWGQPDi9lCYiWRoWDCLTbLNOiSLwp9TEkrEyqMSAtda6aBCAFsa60B7
c2WzOWyPWHWoEq1e7HQfcPFa6uoR/3sQMnra2nH3KCXocjsrnl1N51pnDA1Hd1wq
vlbUzoPhL8c39PenaubI9XUfU85901Siyi1poG2omyxjUKyv7fk/20o8c9hPvHoR
QKO/I1Iwn47mCSdqb206OgKovuQyew8YacTpRDclqvuTL9TrbEvhI6UGkM9ni+42
4DdDuR/GLGeyDFN2dltVbVjVu6TBhw2klE3eQkuBKnzP7Tb8wwfDiCUZ+7th+NGm
loWn4kSmrXQ9iDlTLhmkG8ar6BtQ6MuR3/J/K82e9f+2zN9PECh/dO7Oj/jPNDHX
D2/pAqV9Otmc7uz8QdijJP4CoGzoJg2LQ/V97UBCEEDAz5lnYRaeBu6hG68+UGny
c7T3idFa4JjzdjTiVrGEBqyVj0brVm+4QcbLt8csj0TGp//pIiXGTSN5cqt1nKDG
EpWBiJR9r/ckJzqy3cGVRQZMH3Z7FdfL+vSbjK648E3awZa2i9pCUZ29tuI9lYMg
7I0UFKBvAojAIP6+vHWxwnIYP5fVNDxLzqOUW2hercdLLoBvlF5BY3m0Mqb9n2Qd
mKCapYEYd7ufRaQWenlB9vwY15v7qXVLJCRHfwfvcOuvfEgDEnQNVWNzP/dgpDIr
YGWFPFymLg0C8B9c1sRCDTVPilp/O8l/dwVOs7c0XNYGc7hgJamfe9Qt0vee7cvP
zgFcnt5G7DEA8gSUDGFmbm38ii/xJ/IzPXCEIqqVAnsXosu1rDKh9WYqbfB70qr5
ozzjZW3Pt2njxtuzXG06LhzvjsGfDo2folka1CFKZfRUAzA03XnwUsyxRBmGhuZ+
7Zy3cbn3BZgU/YYMSC1R8GlaDgPOoRE1JtoM1cRPuBgE+Mk2hxF+vtKoNATmLtCb
i5N5YGGdv5gPTEzz1tUs33VG/Cg+4OKCo0dOjw2EjDhamJkR+jX5Y/tmlc8QKPF9
34SBIUkpMhP2MIWjGvNEbxyibbjavpQW9ITmDy1UwMATmfFDZEGJWxXXAn0XdX12
RRHdrudT8odOZV9P4zcmgkNX/YM89nwtIE4B1rk6BSQSHzgJMenBxFLRCZDLWVa5
iwXsaDwYtDrvgoUWdRk2SjdoWACDRA556yExLclZUNX+CxhdnR8HQLAUoItiNExo
V8CaDyUBm+9NsHT9grcLoRF4ShtPCcOe8K1kNPqDYIJbpz1E+TYjWm8N4GScOlTP
1zbwNBsYsx187K4jKQQvDs0aZWc1sSfB2CIQ7bx3u802OrhE1jorOavJmmzOkZmy
lrWv930zWM6ANEcgJ6wJa2QIChJ2Naasy2vhSZLN7oRMyrXXWJpbcqnF1sbr+Oi/
BzjB5thYbz04AzZYsuNP8/Ks+XZPgh5Yw4gciMoD4XQoCEr/anRpO0ytM6B6oYT2
kK9Tb97smxYEuD9zR5ghfS/XStZwrkeGVsdov67JQ27i1S00GKKWNGWZVmYrgF/I
tm3YUrx53FA/wVggqo7/LafyAKbT7Sf0F7i4RyQ5N8NuQHDeVgVFJaJR91ADt6Vw
sWQhyeh0r/XCS7iWpoTOoKdiUqt2/w0jSFJtyI/RhXzJdlR3fYuP3gx4nfqfz8sf
TFQ7JhVn8q6WqyW5DVniopMeDzqdZ6/6FeNq9dwSHBMkl6cdbGbYpKS1rYlfu6MR
FFNLX8cRCsLp5w311oVsXNL5rLZ+bZTE5zVAsQn0KPH2UVgeMwzOdikjpmwgSApg
PJivYDcEwK8GznD5lk8hfxC32ga1m7kFiXxUUV2lozrG68bvLJRBJSQQpwEmVFw7
b1cqN4hZSZ+2aPSE5egYtMxalWBWqTCoGjWrvc8wfE7ZsDHAkZgvs3/Yug88NM87
2cxof9Avm76Ux51Yzp6pm7/v8wNf8VYkerWFu61Uo8eosuAhsr8rY3pZs2xomHL2
+bVfH6UUEGSNOK8ExypeJhwsaij+GsQ+RPmX+i7wUpYyyII5ojw9UYZ5w/dyVaSv
ixOhJnaevybbhg+xfe1uKQ9JFX2mR2zmJjH3Ihff8oGBgXIozwlJ9xBpPRtP+awM
naCVKqjjYpKJKV3jc0X9fcxU+YAWwV8yshjIN3loFej7MivwzVTFOBQ0jXJ2Yvbn
P5xPBSnIzUXyiaBj7+qZD7i/20fd2Cv/iqXo2om0u8tKmobGLy4rl5Ntp4DSUM2S
Z3oLAFRqSjTc5ICmWOatHLIq3AL2uwaLHYYCwNjWFM86sbjdSDlu89XQc4g2JNON
GVG2J5+AMW030jCorhrah/IW3UizYLesXD2ZLplm/mGnMqrQDLymtsxzFIr7N6kx
p0+z5QcxZzgBSAjvUKd3dGnFMcu5yp13tIbeDLCCJYWeqeUMxXKcKRtgXFDad5Mc
nliS/o8v4icn1z2tGeyJJoLmA9+sKXw8oqNXh+D9mdJ+vZ6NdDC7ZIyo/aPIjmBS
MEL+aMqYH1xxiHdncrSRhQh8kBCNHzY6gGxcL+lzxI169Hv84xmIOzoHf69MoWYA
T+w+hdV6PTkXVNtxYiUZ42GGhLS8HPBJi5WzRzBFqtO9b6TgYoFAh9TSd++rOtTa
lM0fefv8yFSZqbxDEl9daTcb1Y7WQeXUuv9eH+XpOsuFOiirddGD8N151duMTEGA
UG0v/h+8nYuQSPSKolXFdLxBEkOP9Yw9wi7NxTD56ZYYMvcEqy7Sy7G6A4Wtg8i2
ObflY/scsLW/SrDSBJSF1PZPy6kb+Pgn4THa5FMJKz+zfEFxfoJOWpLWbgdUDz4n
hv6oiM7X26kqnBVbnhm4WZO9fBcMVOmbrrDx5OavwvLfydkBumfn4cLWvq0uMLE8
6QqImBiH0Ib00gbGhgaaCZrgKcyv1pUZgkQDoXE1/47XerWGwLJ/ycApw25Fygu2
tGQArfww8E1Mbpm8+pzUuKc6luYCN79+V4mMTguCqK9lNun3AoUcmPqZWWhN9Z26
>>>>>>> main
`protect end_protected