`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6288 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
iOS4T16637ogvUHHJHvO1GKLK26X4c+6W4EdvCFx3cNf+Ra1rB2ggTfjom6Bl63k
tPRs9tyf4e7mMk2vZ2ne6hkPuQed120MvWx90eN8OXTmSOT/zCXO+Btd2XigrhKv
a7lwnYFhEkQ35sJDZ+m2LJWqe34VlAu/0VQdYSA6HNa/nsN2cAs/sujSxo7SiMfM
U4HiMgdad4R4JgxVOaPUiXkTLLuP7P9EgzWIf1/pJ2S43xHmYZfsPn64O4QQy1OZ
fN0eFqe8HQ/kfWUYQen0gjJ1361zikSvBD7Ez05LjbI8TzrV/yZoIWXUOEgUHhg4
XkgkQhSTPyjOzDLWARfBc+tfbgnEBBnGWbM70TSU4xH62djOO3NtYhzgOvZ8pPu7
mg5z0WQzVljfX1TguHyhnglEMOyoHBLwGBnrBXPCWF70S/K3cWI2/ysnxvQ/i222
TP60cmHcxoFgKWzDjbIfkQJ2l2FB9VddF7LuQhvZuWhwU+rLji4EmquRLWa54H56
LO7YWVwjtxm9CyeYpCNUBrrf6mcGxNuWgUaz8CaRUoz8fW1ZCBkePLJo9TRYugcF
vI24U+RqIbKqhXoaSVrIicokcVbK/LK5ZsWuqybkJV4Wo7v13ypuScwUSMKcjBD+
ZyHzWylSMgYP7JLzZZ9wh8uH2hrPfhw3+zpoduaIJIsPdg7IKrAUo63YDedhhZjj
8BqMiIkMalIs9jAGxbMPTNx+Q81Uyn/Sp1g59yZIOrtLR0276nODIV0nitd5V2s6
GoFKAHhswytYcMQQMsU+33Xk6yvHhgGWBb5NFytnFkW/sHqe6Y1B395qvoguWyjs
DVBcIKITsfPfepOw90MzNmBI0udJBig77MsSN1Q6mVLCymYbd8Eq9q97oSm0luLj
hgaDPhahMMFY36dYLdu55TOTI7AJpHkmdDYTu6mvYvKB5ojGUXDnxO9Wr7W8VAkd
sEnhlvFkss7swO2kXpxcijI8RsR48bV6TVeqrLrVqv9DqrgR78N26JEhY/KLPct7
XrugPapteMuJbjFLgI2rAELkdsvAtEjFgi6UFzuqlhaO+F3jEatAIYwCUcy4n9sK
ZNRM21wLYAT259Nz6uPo0yRwd+T4liKDN6FRelsuuIHEG3dDNPnOcxhQvhMFMkom
dSPM2kD6bJ2Thz5vHqz+cJ4ahDCSECitc8sRHNi7BDieCxo2ZELiiUVTqR3pemIG
FuQFmbg4KJyfQGlFXh2aJ4lcXvVHCIgcKdLAhmMY8T99v4joFhmtGbcN8HDgDj4u
nTX2YGVGI3ysjpuQjbNchix31jy1kE2l0ndmJTUocyX/cmSTzcg/Py//iVjM3lcR
aFyOY3S8YSmZy3UZV7wI7jD3N/I5EqWbDOWPrw2HuBLddpoeHawjanRh+umelfi1
yjNq48DQ8S4or7IG7T0vBSpbSqWGrSctcsROOdvvNxbFMcmwZANrquwiWyhn6a6O
Wnh+IqOhYXyIilxhGlUH+S5Sy5k88SWDkw35g/EVFui2HS/WFCvniQgJf5D/Uh8T
nLzmrsAyQI2McybDHvSdUeW7mDSmw2n6GlX1RABQeNM8XGQbYIj/xoDG9Oz5gqCT
JZl8mjkxN5oxOPz/gBAM5F+4YQQfxlT4hTaPD3MFannblEA7kEB4F4vpgoVkr5yv
Q3e5p3mVdqkOA6dVvyvSHRvBM1zS9wmbN3r5NfbCIjYC6fMBzJG+c7zxONlUZDRF
SQKmjcBpAJUF3d4F7sBOZHlknn74WSVPRg0GBlJkLorzDfZiHAM8gavd/wewn3lo
sUj2bC1kWnElVQLBzFNGkXFtUY6jCfxotWHf9dB2kDwYoZHfEudtbk4hr7jGLTYl
KLk6cwQEG/7pohh7TBJnopIRn8/u4JoPJ6JYj3+WbETj4Gk9l4z24zQEGQ79/SjF
21L6505jiu7px3Os961GlbiwTVzsTxbLPXl2oZlqRG5nIZh62wQNdeiBtgMFWUkY
/36mxPID/22FRBvBssDpNE8thPh9i7LEkGHwjpVMhpL9/lMeb/v6t586sNrUIQ6/
1yT1EqBZkJCqa8hw35/MIAa5NIkoHYTk1u960qXZ/GeV6VFHRlGdsODDcQabeRs2
Zwu1tV8kjyRVzCSCegqhHor2AFOm0a+cjrCJedUoGk2azSJInBGz3THrULiy/H1H
bxveq3upfE++1M776k7FPFcIm30CqaopzobxGpEn7Ka9znZ/nKhIlYzl9AHA8gtP
3enNlbxaxSGVGojoZdjWea2HnykQd0lr0BVCvGmwtsROZo1rHsQCDik5S8/FCDtt
ce8LYgdA4RwbKcC/Ep1Itc0TYXwRt14xtkOHZG4+KbgIlQMa0DKyNlh13+OE2Hv7
2Hwl+aHGTsjykNXUwVJ3OkW4bAdaUIO00pRIdRQ7UZ2IVixuvtMnjun858rR54Nt
OIoQ6lp1KNM+7XgAJFz+pImXHdZ92aHdYQcJVJBOhG8B1oejrDsQbDna1csDoY62
UJlOg5Yp6y/iaAt3olV2khE3W4Oto80s83zq5j4mFpsBiiYI0by8pz23tLiUj68h
rgdwxBhOEN55wSfY6dhoSd/bMXwxRn+cAH3p5Nm6bTWLJNLh5rMqAqiWvuuaD2ps
ezzIyX70lJP6LqwAE71FC+wwnShI1uckNOHql1SqeR81zspW8tViy+V/4FnSTJSl
z8GnoFXcZ8rH7HbRuWxZpWQIsv1aytpnJ8UdAKlYsrJxkCIfqWqf23U/77XSlJDC
nUI+BBXZEcRAs/CqDnXlYtnLBAJrNO6Q2gFXWXuwTqC4jtfKPheyt31DuHSegmnZ
nZM8lfMiw3rD/yZXJ28xUaTR1NxFJylfABOZ7wCxy9BdtRaMAd4UAUwEWc0xx1nY
mfZkTgTZRAYaKI8PE5Fiqo3mZMSobz1o24iXk00qsvnpNnkS4AvidmqyRYhLyE5u
l07QJipZG5Y7DuntpkCpe5bPUrF5r/fOa93k61YAXGSgqD5xglTCDfnqDEVxlDYa
3Edss5oV7qEyKfNAjIfdVQaJCIkG78VT1WuU4w76TVamu4CEKYPOt0UHTC3M5B4u
34BrWZcHb/XmObS/IXNMALJvrj9WJq1ZHFElRklvElreGbJXK+P0EXiWuQJzvLp8
uGBLazrfrJvwlxHYDoy3BhyY4TakpBrAhvXTKzSViMUHk7SX6ZSllieSNJSItk3b
RNNIDD7T52dT+eFou5pE3vXZndr8jG3WOe+aM413Iqkoh8KcmIVrqxjJstrhzen8
wRPULTH3fSqQiGogcp1zpDzFo8gYVnoNHaupS5YJ8Hk+H6Ig6g1hkHacs+XA9Ptu
PzYpA545eAIbQhSzd4co23a7C/1aVMy1mzYmTdIYMWcLFSYpvEe9Qz7Th1OAtm7W
473NPbocAklxoa+cPD/9FrYZY5Uu0L2uhOWCOSezbTYaD+tW7d7ODZiulun0Rfn2
e2LQ661kscRiPcgmKexOlQfBkieXQ1LjpWpWOr/GDDAPc/A/vUk/xQPlCnG0RO2e
P+NURxDc6sVZMRH1b4WxQopccwyyUKCFSmyOYybMtUwMTMyxXtZJckpHjsuYxpqh
xni7NTHXnbY/t0V2uKdYxtqMphHHq71yJcDuusihL8cXChbE1odXivhj/KQwfN2N
lcU+bM9NGcPhlWETWCeau03yZdzfbE7/JnJglRcUlDdtUS/MU5a+YX+IANEm5OOP
6eG9SJEhzaNwPrMYkSNfJlBkDovGydUPizMZiWnYC3jp3q8ixzjEHmQs4D+j3kN2
SLk9WmuEMZxBsGAGuVifAuM2c8gScetYo/wVdKdyutEbSLQimwl/dqTBqleOUL2r
4/ziXYEMSnj0tV29xEmInDF4Aob+13TaEy5lfNN0Jt2JH6L+IjiP2TdDcTCE9fPD
XeauyP/MBBD42FWlV/SxWzNncOvIBpqh/E9yzBHR/il23te30wGalow6fk0+s9Fd
ux7i9zqPHXTvz5IY0BjAOaTkfqlgh7/7D7a5yk4uVYK1RXlhv7Xr1pw1KeDOBZvO
bgAEqqbeVsej3vyiy9R7JToLgiozeBhfRQ/rVamBw+yCnG+quaTpnmeL/tSVb0Mk
k5bPHdMWylFthDmdx430S07zk8omdUjYvEBcpm24hiVARJ9gQfV4Vxhfd2VqKGtS
DR1ULzPQwcUBgVi43darQpt+jrDntywKC/dGWj8FDAOI79fcgbasXmg6SW8ZB2UF
p4/rt5fGjGg/KIG3iWkwgYgV6F1+SvFSb9SJb0Fi/Z7nNZCkwY3WhRMvVLOyj05N
iYPexNBBHVe0BkE9YXbh1/uXZ2xzB1jyjypkHkRcbUIB3NjYGiWnfAIdJjDr7kvR
457zWupCqKu2zuAkiZIGrEyIYz8sf/VfRU/3DaHRwZprnIbg2Tt97/gnlH68yTtF
L02i+KOfz7QPKO9hhJr6jPo6w6IdxUI3Omm+Vy1Di2z3j/V7h2KVHMy+lS2lrzDQ
3VddOk7EIi94yxFSjag6mfx3KsINp66YHHEGU9qUQQqiDujrPmic2kDq1uMCsL/v
4bsTxlRzNztyaE1JHMM+6VPjg5nci+pbwFuS+R8CBNEANCeULYFLbA9GUFj/KNv0
giEcb/Ao0nNOWjvJ9ozEEndabmyFt+FDZP5s7Jd0t4OAV8GrNl0VtbqirWLy5JNi
LM9sKLG6EHUs0olSMJt1HxNsb+yb2mG1PQQZxonAwTAOEddv3A2M4KDEwHZR6Sf2
KQmnQqEZXInxMEeZzJgf/59KwWpBbJFaKL8Vj1MhVTctSWTpEoHiB/rUn4KS35bO
TQusvBmc2wHISJWliEpqzG1GgMFs5MrVTbBucrpCNSSbSjL8XSqkQij/qmF/CWzn
PjHrK8JUxXf82E/Q/ZD0SSATxTB15AGb4uowecSwZif2ss8cMPnza1xrmHV5kqYD
iijJvTv/xKdpgB+2BrxPATlmBLYwy/8gKduud/d69x3Z1B+0zvFfwSN0mnefSGfF
9zYP+mGHZ+FEA1HrNgX+Qsyi+hoXgchy6hXefxBgx2ow5VQTYP/7o9E3o8FmURvR
YAViWuNe+HjV4AriOy0btjRQH6q6bQNrmF2v3GlHP/HCKgMnS4VWx20IGKBzemqk
LfuDYFyMBOlWnmeMT/B7xqVGybtZ0FAQjmNgqJFc16g6rcdOwQ1n30HoSPaIfHka
e4usI8RrnQ2K3zQYZPSIm/SYID9i5D6y1ax0ooGwJNMQlXP6FSBwtO5z3igjuo5w
gTWJPBlXXemm/OWQaS6eueLOPcKcUZlxeDqqRGtiAmPctyYcLBVQGNtiS2kwL9Qb
Mdh+OwJYdpOMhyj1O/O/xN+ACgwW3YFceNXSaRRbyIkU14rgqOFp99eTU9U4+Kpz
bB7DTtEJ6M4dEEAcAqzCaZ33j2dJDad5fB4b7Q8MYeaT2xNZv+YKI2HvOVErGyra
Tyg4VCGKyO+XsRTRezwpBTvwuZVfJ7nQJwBSIktIcqMKQ8bGnrioQBgJYoEtdRus
Mo8P20dm6bRwcxVNZYO2EllIjAGt+gMI5v3/6KDma57Q9JZkeU7eLA9Z/lXkSDri
trnV+CkbII084nfSnP8NHpGESY2sA7klEefx4MPduokcpyw1WJm5sstAyPBKZf0h
mExxv3Zelqo4XzE3n6h93ew9AQAy8HbNWez/0DVLrvQznVo5UTbvgDSounG5Q0AV
5/DdwoeiWpByZMMXS+iwSA/CxhRDU0Fxxp+AaHR6QgSkEdizC9zHR57ocZoNFZN9
hebM/U9gRxWqOQmd3Ian2Kg1Rth7W/QngJLEMCmDYpWvGGSnl7XvDNuwhFW6z2ZJ
MKIg/bfQzlm+5Fe77KlXM/vp4oQqMNMyGP3fKBoS2JGEZPFkRzIojfOdl0UuFQSQ
sFbmbMaED2WhdHijHU+oUouolcPed8LqjgzF860zjYY3t1EResxM0nwlVNMIWVtn
0PwNnt9+mITjEjHaZNJ8irnFyNYrWKI6Hg7cXtj8R2mve99Kf3P8k11zQczl6Sdp
+npp0KJOrW4w/NZpXyxQHud6oQdHVF3eP7JZpyGZhltOxR3I3mnEFDv7DYkDFqeA
u2cUHMH6VqXNTF5xq2Ta2tEDRjqx8IaCUf0Apjaz1YnMMWfTrXUjFzSBhusM+4Zm
XD+nO0jvpk/LJ9optMZKG7vOKMNmTKU6y7YKj+2u48aUWK0R6SYJsgld/6cPowbs
x8PgJfRDnu2dcS0t+8CWUBMWFaObgvRH9gLiAFsJlY6SjKNxni/W0GG2HiFjOlfU
Ni8EAX33Wf/LdiPCCR7ra58BXOCCNf60PsKTss4AOFuVN+imPEK6VMvbhnSrGrQK
9tI4KCRLeNWtgxJ9dxhhh0zIa1Qf/4Tekjk+nLK4/gocdy7XXODCF9X/XGYXbJ26
bjaaeogfmic7uTi/E1N7i4B0F1/iz7s++JIB9KcoA0jEeYADVtpoiFjWBOthi87s
NmVecW3BAkdvlpv9twku8GfyeLZtR1W+UUmXPbKjNWxwuR+74j/B1BZTZ4ZUGaN+
ugDeaPUVXlDewWms9eCFTsntJnRGvosi6v8mpkafFt8tfNxAGVo2nrcXMR8whvCC
8BYeHoupdxb7kOL8fTtx2K6+wNFxFQ/VWn2oVLMEvZIyxA+8nmPR3Docpw2yQ7xU
gQxJyk/Sng2l7vghzRj5uLIB3/qdVsUfQgLFLgtN73sm+p3WVmqvDWVjp5oNRWlj
qL17phPLaPGlpqYZmRSGXs6e65qCQyEeSm+Uoel+feR6MYTgjJXfEwRFX615lPMa
5eCEidmW44JiegiqPyTRWCb7no0OqOBt9J5C+Tx+fu5tnz46RGPW8FRXe84I4ARZ
B9ZozdjbieuJv5GLtcLN/dvVWR2SP5eTEAnuNWYxllZ/i7W+lvaCUmer7NlZl16s
ejr2tl/AnSXgHklQsEYjs/F7cvT1YNjawVi97VeScUmlAXjiS3K3zQ34KpRdQ5jV
umEI3N5B5byndvdXvtHjdRr36fZB1mFbshPOWv7e4VonY1Xie9B48ZzvfxGMfEdb
bNtzCJw9IK7VvvTbAmHUSC1NSDem2Qo6uQ9FKheRh4TnXxO4fht2y/y7uj60iy3p
gy9XoY13uY3gnfI+EoJYOVtFVCScDLXQvP+iBzGkbyCi5qp9LCA15epA7zDkN99L
nQU/ERiGSWIiFzs66jL/b7HU7BzjFd20yBpdaDzvYjRtbe9ki0o9UkFOPPaB9xxr
ZwBIOEzuz6Hw2wlhUzcNGMY5ZrMwZya+sTRrL+ZMVSMkV1/1KCB1jAwq8U8GDZbo
lF5GqwuiV82M+OOpkBL0ggTO4+E0vVM4xdvAteyd7YgjJatg+55xgUXu9nd0vuzk
6dp4RCPBzK2T8peo9nzrEFk5B8CMKjVlTFwMSLExbTNuTEG01bBbbf+BGAnOwSKD
L33d2qGzK4SSeORruylMr9pCSdWCb2QLP6R4lkdl/6I6ObxxlfucMSfPqWdfCYxU
cKYDbHdkzcj5WvmcnqByjWNV0LlaaxWXnQ3cG7Ze7WMoikZrmXh2HjCQkQ/2zkLe
xQxrbLI1cNYGvMkfKn/OXghtYvHreneb3Th/vpEOL4wA7zIgErAyupvy5T5IYYZb
NlpXDpa3cVxk8U2x6A8wbkP3wIwc2IcDxh+BsjvHfbwFz8lchmfJiGCkG/EBEgC8
qiqM0DTAhSUn4/fR+wnYHMEOSF2dD8TiaGYe27jHC5QKsQSWJ/qzNNedYa+s0Ejj
s47ceSMW1fEf4jp9gm3QQYJAxsEDGzHeBn/qXQCLnrjlqvPoEgBKOpTjpqX6s7qr
4ZnBygdbxo96fe/EPTX70KSmktRjTvLg0RVda0iwfubqHAZlaluB/qrm9ZkARptR
RuAkMm7QL/mc2D2Bx1tc0OSFZm41lmisJjG6QaokmTfBBKgEqrNDT2+3KQ2QKnnn
In0y0hL/vcn7EYlTSryTnItL82WEOwwTbxaqrreILfM9ilQn+xDDTTJ8NQSNbnbf
JknsG/4Hh/iM6LdYo7EKp4bPNR0QFsoNXFbPfEt6xZlp2KI5dSCuyR61VaWhS60g
sWwV2rlYpKhe3DeoW0ExHcMFTY8oHFHQT/nwnedbSJPI7fvNdEPuW0Xz6hSffxfu
jrKbCGkCHBDhyJQvveeKrSFgXu5NKr72p3LeDiOnhqv99Bvax1oZzy5TkS1xH5z9
+/BcrNRW22vpwcznMau47QWY4brHdoRb5wszkig2zTt48drRwNLiWcFk4L+7p1lO
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6288 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
vWaiee8LnCgatAmbQJm76O1I4IXSyRJhY1P+pBoI4QvgDqW9kg0aVe/0uIOYKuWf
OIsFpqZz+smuFUViTZ7DBMj+ZI1i1VFtcL26ejajoAQPOvfyUJVPBMDve/UqFMmI
IiKKMi7EX5SIgOCs2E9NeQIFv8wsMjfT6eunGFsYL3syHSvwtYNlqt0q26AA2aSz
DhX0PCkPbhK/TJuVGEFnLa6lfqbdjbyVFCGzfgZAzP/8geNZriQfhKB8cyWMkugz
GrVp67Evtd697poWfI6+1XJ44N5flzB5CM5F6gEiU0Q9+pH/1Wejj06cp9TLYsBT
c0+JJgUx6C0IdUY/FQM88/vpIDPrOaYCin919sTitbH0yNSXZF1Q6DXy36nxx38c
QSEcWbrxy1zCjZfpeyLLaTy43f5xPhDvnAOzbpgmeb9WKff4nfoVznwLKSIHXqCd
IcJVMhbjEFgFWMmyR5mIV3X1vADT3TFkJhbFEFODxuoZ8/kJEjMrXOxxRwFVLQwj
W+UsNnfX2r+gJ5UrylyIp/olVX/Co/9nqmUQXlBjz/xSXSqA9RB3LwT+NmuIBgf0
NPjXWLaXLwqQa5J7Q1yaahPXLmfycS61uY5fw01bXO/oUKTPwPjClyHxtESBpSob
jtS3DUzEMiwvIDL57WfERlQ7URoIfgMEyaaayKGpJEVWqvvROx3nr5mSSbo5vOkm
+rgoF/BmdJbsNd+mTQQ8HWDE+NAfm0fAq4u++7FNeSNq9xk3FBBPZJlNsyr4jsTg
A2PWRN0wJQl5EuxyzeSEP5/zSA8L+WU/TevrXx4izdWhXhyRLARtM7UlDyHAkNt2
ftbgMkHS8UlcW15gAlAHMWiQcCI3dy9KqRwTKMCGvZGJcgjSdzo79PHXJj1EK/ne
A/R3z+/4hW883LD7JuEF2nTT2WADBGhK6bjbwz7Op1RKwePgBRdPAnIOhc3d8+P9
eFa4VhhbyCdriWHivhmhLNPw9LPM0pjZPHoqLRKOWBgg2NFqPoKtU6nIqAeb+T0u
7oSRXx911PoqaP9FcBDPiv98jJyrPbiI/qS1mtJO0uAxRyhmbvRqqlTi2geOjdVZ
RHJ09TnaXYj/MpACi2eUgHWLlWT+GvFnGUXcRINCSEKtKgapIqRCzYtXVImSfVOo
TOXoF4ojQ0syV71akMrYNwGe6J3fxsGuqJPgeIbnjikkUKqqGvdJvuL1SNS/2xW3
UKoRHpOWG+i7QGMYOacctHScxrjN7e+7P8P1ZwbaR4iMBzlpnm7yz94LKBD7Q561
WHhM32lfXaQOWNIzOvmiNxUDmOjXHJt9wQtCkGIFxuhgJckkjwLswq5Z7GdKdgHd
JFWJxfjZLv17IO/6BLKxkLMDkBmjJrG/31l673VT8ONGjzUf6l5InZKJBK9LzlLa
Bo4U+NG6DOKpzMhher382WPd7GCs6USyFnYfNMAtVTltUeUDeW3gHdho9xw45pwW
fSZL3UeMcS/Mym2fIDiXZjkGVEq2a34UFev9GlQY62tXcxjUPrxinMTNVC+tqbYC
KH6fywIdP4cL7eGBHDwoKvydthQnf7wpi5zjTv+Gxn5mz238ExBbk1AfKZ3eZoYX
UmnElVRNVfjkhIE5clizUMlTZT/FyqVQsPHomTp+gWQi+jgThreRgZHKB7lF/sWt
5g/x5FxiwuC8lugefegQYSqsnJ36KvXWwSOZg/tv7W9dTxqX3AlmA9JaPnNVKZpi
YjpoHm5CjBLUfjPNnS29QkmxGufhWn0p7rX1koUqVqlC9qPhNwjaDAzizdZOAIpG
wbECWvwJy01O5b7vG18KXdGOVdeFM3ip9yyrlhQxN4KcBL/mI33utafEzwnlxAS3
SNmB+LYJNF9GZnZMdLGzRhz3bTIE2chLaL2FIF9QtEgNXJMRJEi7xJ/coiIyJiaK
n9MeY0Q8w+tzANQQ49HyR2rMuNyuDEvoYJsLwBOSM2fWm/M18WMLR6t2bNTnlynp
Dwk8GL6ur+u4pZiviRDCCRF1LgZmYy3sVM0UkyuL2BjKOhhYu49s3jCeiZypqu6i
r3l+N0iWPGKFeHQ+sFjIdEAfHh3MMx9BhofmnBjno7VIJ/cS4cumyNRNc7EW/6SD
5OjrbPoZVpHTN74pHkk6aEOg0XPEVPH4hoP5q47kiyDtONobU72HOukMsjn/Dgr1
Bi5RV4Yop4qsutFVnur0iiTQ2zbqMWTrY9H50SubVTYHeLovsKnCU1VylBmhxoGH
Y8uUzocMHrmwo96XeoZDOFVIzJw8ON25yDEqmJrYtdcFHEsjoMlES8tGaFPWB0QW
abVX8AKwZNZ8hhLGWU5ctuRitAPRliidiS9PTuggRwe8+7TTV7DaAdMDCFj+4SmC
mL5t9t1npRtIsulyEJ1uAZ9qUNNUTVELZRNbnTm1WP66xWbhxm5f6EwFhdaWF3sQ
XOVwzbh2diN0OV019GyURIrR+8NjJKItjzY23gyAA0XhbSLuxMlIvoQKu2cLkTIm
iehicWbdWQUCTijGkWzH1oYKoqom8XhvnxnWhlVGACJRn0MlCwjvEScENLntAI+n
RMe8S9YKCsZYxYR/hsm8AJi5gOOwNvj7Vjh8S5KdntKjZala98SczfPBHNH/UPRt
kVP39RvWGwNkVz7uQSHBVt6wsuwW5I+fXSpoucuSt1S7WERTNjd9y6LqBove/0W7
oB62lVkjKnpGvvCYHWivzqwrxYsApEJFcqlNsPTvC5SbW+UIKiSTPuKc/PRX+Z8m
1BZ60Tz9x7pHUJA7p1muVNvd+uHGdrc6bSD0DIvA4YPbixIMMIFuVmAxLmeqCbd3
Vq1p+Lm0+bfbSE+C3JxH9IeFrUcukJbmogPi+vQME6p5QuZ55pXqTIwOnnTxTInU
SVDI4+a2GHQWHoZNUht6DB6+Tv0SD7slR0ZLWYe8V6A6+uQdzJvnfACHvKiY+nV+
xLIfbXtCCoE2STFq8MoUgDtNKVaysaVrw6yZhlut6U0moh9YLxL6SEJ6imoInyyC
p4J+TLqB3NAlhkzACiumn4LIBA/5JsdJHmof1sVV4fskj0RwJ759/NDiBiA2Hwyz
9T2rPpdbGV18afcgwtzB73OeEaZnQeqDBdrgxJxnS6Fxy1Ci3VqsOaEeCpJ16MDJ
mqmRNAuPHYs3A/GW/pv409hKGCmimn5F75FMOofdPoEAyaMofsR0yTZqLg6wonPI
/Hr8+ONWSD+SH2R+CcwG8zY53G4FI2lk7vXi/i/XbbRU4nt4xwjA0ryivSC/Ouqc
Xhsl5sXiIfQLZls+JVCC5B7hqm5GiR6HR+nswvVx8ThkDr+cVZ5OjfnnQLhcWBMJ
tfKi4kfbnmFrj76pptLRHo4jxLhigQ22dRHca1sKPfHYV1+oLQFri6/AmwBOX7df
tsefhfaMU5U2Zv9KAIV5Gtwc7zNkCpAz/QeUfdcEpbZ5LZMYcS5BF5e/Ob6EOoAm
AMj+AlqjGMbqbW9mVFDRQ/idQeH5cDM3As3RCrdDtZFQ3lj/UW5W5pjjU8a+iSXD
x58ZPu2yV1qqkl57LGhXmaezav8aASwR+gs86xSI9DAaeT4PReD3F0YesV2sxXEO
4Q+f9/uxkOkV4Od+Mn347sxVpP8qQXcqqCsEWeF12l2dvztjHXoczh5WJnKvZaYF
D2eVMjmXSQCgQopvC1DckzxQZY5KhWGPwdNxCYBOaUWOUHrZwafOP7HZ6Jnj3CvD
eGBxnxxselbzwZB/S+l9AN2nYzQvhk5sIXL4jAZhtsBOArE5jCl7ZPW569k2hQa8
TlycFE9S620pfNtlR8hN10ulhaWBOpJAVvxPsF7RRUQTO/i9GwOPO79iQXZaJAYl
iP4GZ56vAu/GgcDI3QrPQx+WTWc0fDyP4r5SNWHMOl2zf8mBPo+mGnjIefzNc6aD
sc+V0vc8DG245oi7+Kkmcei/0hUkuAfzwBBFyLmnp9heMbytO40VDbxaHioo7sum
L12Slrc74iH3bObm+fzRjVUSH4QFEbja9KUGW3C0KvZKE/7uBJib8y4p+9JEv3yz
lT/Et8UyjBVo5x6wy9A1LnkB+vwbc6+iaSanRyWY7f4Blhy5SwIepJJaLAhkHs+H
+fwmfWK7FgX2u7uN3MyWVp99WFFjWgNT5BHdZ6yA5npCJ6s3WtIOpbx4p/NI1Ssk
EiyAEPxYXgjy/7SzWNFsEdpEN1LheviBI7KVFCG6bAAGFRTYs2qzt5RuN46T3A0r
IOO+H6eZJFAuwhDodk+UdVuXStx9CkHshx8J769hGMDyz+gfjmHhMmR7KXBxkDLO
KKzvD3q+u3st1F3WJDKAcVRSbGZj52gqfArTUy+lv4LxmdSF9/TodMRo1MP3VJ0I
2x8/3kB2ZZo6Bc4PAnV9MbGzRNg4aFcYt+SQn5q2LRDfa+Y4a/U5wt9B1pTVQvVm
shJkW182nC4F70eyPWve+QWz2zR3I510ac3Cc+zDvDXyUFkhG0M0VRGjV4CcSi7q
Ws/i1Hy3Oi2sj+rLObLgikh4eiRu+uhxU7PT94ilSW0A4fTAV4ewniv+AcDBVsuR
o+aDpjvgauK0DTRALKg26YzCrsT9Ufm75nDHWOLfGSPQ6JBSr4OEy6gvEQPdR9Zs
3jhidSOPNvRnXBlQ0hv6TOINgbn8BJ280jWg+1HE19RI70XcT72NrsNd5urKJRNk
djmmUWDWTMerDZwRDlUGVCMlwogKAYTL9lYux0U+GY6tgRpYqAU60pZxe0bHX1dy
lA4JGrT0qGH0m/iBSUp5eTri2QC3YJZHMg5/6/lHPbWiTia6sG/jVxhG+y92pVIC
2HQA35cyhxP1Jp6YJcto6bWS9JhO2wUExDha2KYfEzddUa9WtHrl73+7QIIpyfuj
x0WOBZhY0+l6W91tvajUSWzmBD9irHqrFyi9seCVogw/PY3mcCUmAy9w7GizSQdf
hDw3qrGzk73dDBHuihlbzCdSCuBGeslEmx66ZYOQTyUGLrIM9I0BcYwn1CXgCsiG
v9ggKszDFu0p69GTlGYZfbAcjOC6P30GWzN1mikQI+GlrdkRLkkiOS61/MNVHDDI
Nt/bxbC6GcGfHuJpLh5XbJ/vsfyxIjh90v1q3xn+W2WDDAu3UAjVMeeefXaKsNgv
1EFEPSn3kMAj0+E2O7Ik2gGCNMJ01G2FGpfFNWP86+O2WA4Z1tiLfUPXToLWmrSh
wWH8Fu4NaHHeBekC0FfeKfOeCmHD8S33/y63ic1TIPDJMvXnlTK0d/TzCWNxKyqd
4ySzNxEek6jjCtAlYTphKVBHRJ4BAE+kUowiuoNHiWPVzKSBoCA97+NRA4kI0rE2
ZWRxNf2Ttqi8h4bd+pxrQM/OK0uviZCqGQAT3mANzTzFvtoFuwA629afOrWhskh3
7UC0E64tjX/H6ByDGFOZEszhKllrj3BcOhr+jdcC+7Ra050cnOcdoBtzfMkvURLO
bptPULhIxUyuA2xqqkGWmI4gjkQIizBOqbcmam/IsonmZMRSTAC+1uzIcAnQWH2M
vWghFO0YeY47HVhENtmkeOXATc95VvgiACqGG6xlFGVMUzZk73n00IausxPqrVrP
AZFnYBAoxDDHr3PQRt9Q9OD3bdNBDRPS5UMpuTbXxSz2EjNr9/G8rlwlkE34ZPXk
A3Xou0wJpRVbY8vY0nhh6s0QhYtm+ehWusd25OiQicgN3mal8kOSSCfwQuefOgHV
eNPmUIFoGOpDU5Bs0ED81bfTopeXOtC0K4C3PUf6u+eQPpaRppO9G7t+IArgkF1p
gIKOyJ7h7lUhei1w6iq1MZnk2TABGGgEn/+GoW2aygZZWeyVa00118YXPaxmTjs4
4lkQDTkrlSh3vfxrtvRIweC5x8Dv1bn7VCIPar8vLO3mE7w1/L3YgT8vhFLrM8FI
CmpR1KLRteF1JCVACaX0r/jO+26mGJPuOoApMuHgc4RgMUCPZD4GaXW08oR1ZC0o
e1wWubBhFKjZFMExRirh5Rjylme05RQNbTZJeb/Oki1CRjnAB+3go3Yy3v1sJR0i
soQhKSKdsOVHOyqiKZB8Brvx+yN4S+sDpgSbIc8KQPKC+bSjKESpGMexSDjRMksQ
wC9DXiEjevnO5HV3qsmiqGt8HTtap9NM24v9M9RByrZUx9Z+2cYwiu51ajJSSlUR
BO2qTpXiQ+J1O2+F/tK/r8Jm+ynr/uyJzwuu2KIz4USXIIYSPrAFWgfKHFA9w6Fs
irWqENP1AXe35/COllUTcXfMxsVs8z65S6e0OyBJ12S3+wyOYG6kEfj1i1/HC2it
65nC3osEAeXV5XzOLIUAbhky7Omybtt5KH1/e9qk0liVU1ocJmrx/TSvoD2cIlYn
0j9XNu8C+MTdsZs0dT8BkVcjYHSPMpklnGe7bvG+WQCR98WKGhnccpBkrcrhrWCV
2ayOZlDkexHSGk/Z5c9lyUwCsFgy3mCEzvV0oz4Fg8HKD27aikuuxlxog6ryxIIB
pzc0WnKvas87ZljfdX/DYNNSmk2pQ7Gd9nf6+MJZaIBM1nyVgWiZbiySdYCHtoBY
cDIf6EkqE0xVYcrA3drdM+SmqSgPZMvAaj9jZg0BsyD6GzvE3fUaUCVnII35QuhZ
OJ1su56Htm/SFIU9LkfqeqLVCr+fpI59EWcy3ttmjz6jGl1UWON7DIIMzm/K2b6w
16Pytmen+3Ji2JZqk0tWmmGJMfD0VZGypFKekTW3kox3gD2WrywmW7olhEtHFduG
Y476Ahm1G8XmnYUaTaAWpDcUBi+ZBzgp65GJJ0W5ixgcvHDNOHTMcixApUE0UAhJ
TkMMQdXpfgiiowLji7ZUXRobroP9Jo8f9ZuRzdJy3mGw2sdmUvCcYzH7KoHE2xtN
a8usWDqP5TIF5t5tR6RwE6/y3b7pOjo4MWnSqs/HGzckX6gvjyQ5ygJP29M35R/E
7mWbj7iSzVtzwy23rS+g07LFppNcuSMOqBBZTdmyNHwO2c7xfuVBhvAtK/La6SQ8
0hBVq/s/myPhcdLNpDMbKSAU0jov7MpIDqERsAI6ALEWTUqtBUKEtJ6/79phzy0R
sO440yYEgw2Du1qPUYLNFgpS9nkI2CZjbK0muX8oHLLeZo884W498Ek6EIXqITIE
NvZhuXVvHqnL2ihdQjqPfOCcwJURLstEZ2BzA+faHeXpS8KCxAkFpVDcYKCUHHM5
bFxobTp+eusqWkO3uuKgwbXgNq1lr9swYCl0FnnDv7zoV+wAduiJYfJd+gkZQn8n
ZMhi36GzoQrAgkntnM0Tw/SSsknv+OxJM+kavm1eVoehZ5QsgvrifJBSsOnNa6fK
o1qays2Z5Mp3AixYJwiN7qWZsq3ir/jKIZCkFUCm50Okpq6/01PAg43mgT9AljrV
0Y3/r1xfSslqofMOF87mSyPy/ZVUW5FTRPj+G09hwYpFMaVmzL3c7mmFH9IRghi3
NrUcWhB30GyIt9A0GIMunY6dTHSiMTjik3F3wi//whFGN69UmgAtvHWUgEQ+ugit
pss+5Py4nMTzcUNBzW9z2YBbMiE6joBWw2G3h/xtWubGWAOTCQk+v4HW1p3LpTO4
eD6rWgxJhr6uGUUsrt3+f2xp8dXyySgGUT9f50WZWSa+tuCPoDsCvr6TJ5fxz9kr
HYeRfEEFukFLGYzCcz5W4JNUT/4mD4Ed8xQaZbVjrO+ZxKdY+9movIrywBtk4g1G
WdWg6/csvyJF/Iv/nHsTzsQxEIZc5eBJzqNBfI3/fWAzMLejGC4aKF5GNSeLOxoS
UXBGSKEH9fwZS1iM7ilLyztZzV6wnKXachV34qR+xbSHAMxAB6PBMK/yWJLk1KJo
HavuMGEPo+7e6xP8lr6/mhVxkbWcQ1BhGg0LGR37Vo5qMjA0UxfuJT0Q0OJo84Iu
aczMRAttIbbcTqQpwsoT3Yk2pmMH6brPefNwV0ehZ0KQL7OhPyl1gR2Qaxo4hLsf
8j0ubr0PQTS5jV4uydzXPfi2VrckYIdyZ3eN/SGv2l46waBXH3lXa4XfjKt8Ja+Q
SuZ3k02uf7RR0/uJ3K8GSamIpyS1IkyO78egkR+HB03CI4tlKvDj2MJ8DchLYq2Z
tFyO6euhmevnOeY6Rw5HCpUvI/nsHE58JNp0RGvS2pqRAXQ6BsN21/X1cjW8MUXg
tYFaFuS3+FrhNbcCCITFN/zvZ4psJl/8cihu6kr5AQNUWSBRo2q3rdOshtqEVjJL
F9OzmM+j158L54L7p2cVP79D7FhNNrckoYZ6nMIHP9CaATx5YPk5A1DmJLZsgc7J
>>>>>>> main
`protect end_protected