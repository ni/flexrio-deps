`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 19632 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
dnVBOIGMhMFpJZXzCENQ2A8y7kPmzdhNwn+NPv8A3dfzBFeHO6nsFIPrvipKsU4P
FoovXGs9OMW5vauraPvfuLt/4VC2Usm90RYbEmbtKGYemPQxXHoA92tzweKvjUig
NvUf/JqySxCiPvHvoAuFvoinzQfWFQtMurPvjwNzfugfsVRtG6kzV5t4m9WJ7geT
l20UxUMFCAKs1bv1Iz6Kw5VJh9BpVNcizZHKAsmQ7X98COwn1uSpSpP+V0dSBN32
iqmayi2UH2c+0FJMyrssi9pzgXBkkyU+KmzFG+21nHYT4VZeY1FKMkGNCK5SYUXJ
XT+TmGy/0v/cILfLnCQqUdBgRp0HLjpKNEkcPQIbQ/rvkNw8NB5IWA/ed7Rjtbi9
HjXedKav0dnJyCtwQzGCILbyVd6ONgf0vPNJ20RbBPFCHQpuZTxL7EbNQn6N1M3d
X+sQERAxvJm+j7Xl1vHlFk2BMl1tTNKOkS9blb9bQw8jGaalQSyz97jptnMvqRie
Kw1O9OgAB7Xp7Vg8TCi5A9oPOZF6/twUHXXpTdAGqlwfGQ22q4M4AuLAbayK896N
7qCTBexIUz1Tj4ZglPbJwItNRGeBh65R8I1l+VmbBnDfFih501r8oOFH5+/bmWax
OJ21qzymsV/5YLHfUWW3JbTeCM/w46t0jwvnaBJQk/2wkJG7OoajS7MkMl0HxZyP
N9ani+GJA72wEDhEERKVQTBk+7FdxGcw4gDh1wRzySyRIvBOm/enq+TW6fh9VfC3
yAe+zde4Tk+/lb3IvvlTEc9WtZwNth6Sdlxrn9PmoGCppSmb70jY5IdJvDtih63+
14CKYbOOrkzoLCxU6GguBRf4ki/zFSdRUG6H/AmG6k+Tl55nPf6xVhxNIuHzFfeF
R+692KClVDAAEh0T/Xr3m+kyTtI43nTIF4FHZgvFaXCMRM6Fhx7L4Mk8Pj+faWBK
bZvbhFngsB3ITnwKWOSZNvhmMBn2C+1uqqanACyNjS6WKO3X/92lo3P+A34+LdTR
OLsw/xaZEvXO6ryjwJbc4/2nQtojL1WCl/THX/2XCCSwGo0vb3uDnouAL0uC2LAa
cKCYcZQd3DCG0/yoZVV1MB1Yze+gMVlJkx/Rn1suIoeADX5eanlMKy3501m5SQmH
sgwWsRS4iorsuAhNh/Y7XIHKpE0T428yria69iTqcF9nHnlop9fDhWN6usJgb2oG
w06erIpiiL2wBAJ+DrUgxwJ2Qgccm19Wy4IdHrQYmu7dL3oXsjeSq4K8lj77QCYb
0cqut6KwK8Tw3bn0kivqHBJPu0UK8mANIX/Cl4gHo6PEh808duy9fo4XEwBCuHqg
iYfnoTvhX1wYGIZIOE858W7uSIULCKtms1rn8LCSkBcyiv7xopHLHTnjHi66fuwt
6nOQ0o8KPLzjjSn3xncVGzkCkbspSgsI6XK4G5MB/Gr9wCxg8VCkWYBRhtrLXv4a
xpbLa992uRahD5VxbDoNCLHsE0lwOYXfurdOr+Cprv3Sga8okotcmirrOZsxcDmK
REyYSgjXtdU+DMQK+OcmlyS+bOTe+IHZJsW8I+TLJwlycYzGQIDMqAV9TljuVeWg
qu+P65eaqSYnOLqOr9yulK0sbT89PChkfH4tiykczJnZYqn982yncvDchLJPdvj3
LPB+v61WfrJvSw1jUf1BBpwglyHIXr6jmvMI4Bk7ijL3gkdmi1wO6vVZ+FXtzpIV
w570TRBjGDFqookZ4/k3UzAvN66zySkFE9R1a6UU4PscyHipzz3kLKJiMTOKW/6/
t4DOqYrSc0yWXIksFKCThBbOzDsZfrDyi2NASOpczzyIbX4yrv6OFbF/LCAyVp1S
rfH03QGlxALThCSWgFeAG3sF5NGrLLMg8wOyz/cofd4vOAu+c+aOYQeHn5/iF8lv
jooUGQYPF4OTpUI4nPjbbAzueIczBAD+csBhAI6brhBPbcLRXj4Z2Lzx1KZiq7Sm
JVf7AvFDh2fj4hHazpH5EFHKBP/8bzI8ajW8j63WeLy5ne5V0kKhtYryLAx8zjfO
clXlukr8gY6iuf2KjxvU1FeWt/2BoJ7W93BrWRWVsHaOHVVTyGTMyqU3OglJhPO8
/TBBg8y9Pj4sweW8O5blah0epBDvB3iktX3o2dzbr02fyzqnYBy7jXkpV7/TUklr
zq6hCh7myGFyCNMnzyxZhW/3MUkoYdcP5cWitXQv3dVSghD3+rXzlP3suMHm8w4t
JA3/hYHoZNIuZW5HqSiOAi+ER4Ejrt82W2kDIROvqnyhz4n4T2TFp5MUYGLT+O77
prXBvzblXIcAmIzw1hmpxsMV2TpjO92lYe0KiE/q3yR3ATEpywvUEBfn3eGAiEnB
UNK+LG33S2OjHIOYEASpzqKqCecd+ZgSHsG20uBjxHeBfP31SnCjSXYgsbwtieK+
QcT8hZgECQX02d3Iw2N25gRTVIa8Km8fBWQKBs5NpZ6IszEraxNR3T301R1jtDv/
A/lU+Ki1mAg+GbEfBIC8pg/r6HFmUX+KdibBpX+fJEgbo8KoGv8X4d/tCZliJApk
Jsc2O+SdnMS0FNy04CxN38ytgme02z+k/BKX7+8kT6VsV5y+l4Nh6+d6xJjxqXMO
Pyji1+QL3H5KNKY5xGQkUUfcbZvIJkejc4HudmF1FV6hc2z8L6AUgVaSH1vYgB0K
thjhKNtMNNBMDULeCDYP5EmCzv2J3+cr3Qsw9xsHNaQE4HMkpQ4O3XRrHM1WFuB6
zuicOSuIU3e/P1g4Ksjtv+ROOcWZQB+l8fTcgzyoHnu0sAdcLq7AGb2rB1eZhzWV
po1zAf+BkDWQOuzbZzmtn7BlVbbCjoWWFduaoiYrVuCwSLCdxlUSuWlMorT5sSA/
PBg4xqA4+3pn6SNsRrt2FRXykNFeVIQburx2h9GfkV88gRy/Gx9fRo3XgJMKggk/
7UXAEcaVgB1q6U9eqIBUHVLpH1F9OTKoy5wuVmrSm6h24P86X5W23lNSUZolKptV
3dE4KctTpxwJF/Ccv/+aZQlm1Zmmlh0eRaClIc0UU7LSXwXhayAT34xnZ8t9mHxC
HZrWZGwQMslrEQ1qs4iC2PZnk5ymZGAIBB4ycTg/E0AtzVjSKSGFCb9WqPqYW4ny
6nYb8L8PV6Afk6IbagVFck2+h7wljoHhYsHF/d1My6/tcaTKzjyy5HQEgEchTcCd
VfmGH9YiT/9l2zAfmIV+Utw8SQLoaVnRm0+9RaX9hNYyCMqrXNiBZQa4IChdcYeY
+LmN4I6h5SQk0mNBXp6eoUZfkOyuQJNKMEiTv4aX1ii6j8V3QPjhO4+KJzirt/LV
OqlBvkrzamXHy1eOiI/E3vN8Jpj/LaK/EpuTHMws7UTcsIQA4Vyy+HiFNlMnxtdR
kr+zYS4yxZXFoYMwnCBYe1VJYDJddkttwoQ7qodqxd+OFS2EbzHR4g21W5WMOyeT
65x7p4bH9T2OE1kkpBncrykJ3Adf0szHkUwfOCtd9+zR7CkvWbDovo5wGgseqUNN
t4cO+QfDasDiS+BIs6FRYmyoGrZNgLOlJ2uVQcrwWyFc/RvIUHiZVe5Q5uW870VN
V+ivaWMFjkExfnaoI0EsL8UglSgaAPa1IBxShLFq+fFeo6YwZYNm58iGonYbvKHC
Qqxi8VK+344lTvvmpgtr1EIZQ+i9WKuVwi8qBTIUhMSqBVK81VQxNMfXHPScNaGb
m1M6Pj94JZnA7rCuCRqpoBjBoE1Nx7WVyJpxuFTmUNdFjbBg3hiEevqW7IjuJuh/
MsU32JLuBt7H9SI6y0nobp92duC848eRHxN4N9evyT0Meyoot3lZw/0xl9eAArdu
614kRLE8Xt4NA9h3jgRUh05TbWd3gW/lUnjnqEIx3p3TYkLP/UdFr7+JxlLHmnnH
YwOwlRq+icZnDKijs5kuav4mkK7+xr4Gl+c318XqnrNIFvN0R8UfWpvl7kToToA+
sOtvNVum0dRlUKCQ/3wzlLkxokf83Ydkl5ODCbNWCOeUpEFennru0Tg+AkIhEum+
2u3ggw3rjtwue29lk/0dDWbOzSEIATPFSvZRgSLcY2CuDVreM5V7vxXSOy4gqgsW
82KsNTT3aRNz+SnpRpP/fvi4uZImLrfidLsSfVTYigO8+Fol5xaHTb5EtLPj6nXM
awVv0+b4v1UxeM2LilScP+iRC2cKL5b06Fv7TQNA9vexNd6gEYAPUVO+lb4I1zNZ
T0EoWZvqUwO9C9KdcDH2N5DlY4W4Z8HN9oYQbKMu3AODjp5DhrdagvIo3bS1l1zH
fNKZu8XLfkkFwRw2gjhalDW3PP/Ft7HPcdpZ15fulwGzugtcruSM89ZvorZurqtL
fwcFIsiCZDWIyCSDYpQYqNDyX4tcis1GaHcf1rbPvBlXGabxOvAE8EKJbQNylMD3
KQ2R+ZNQ7V2LCOGrvaCEndxbnrZX8DfMKfKQONhHb2XxOb9HWgi/d2Z/nBFR7oJn
SfTB+SE4qA7xlnpwOw+jMwHz5fQcWe6DYiOxWhMT4gdkE6nipvxB47IT24jzI4uY
Gji1YJ9LW1FpcmYeB17ZhTDPEo+u9OzwH4oqLxtRSNkuI2gQeD4gKeGT4R/770hF
Ew8JDo57uw1xYqDtIO0Tk6hLQkctPqDDpjjI42RA9t1E6wS89cG8Zl9jAlQ0U59n
NbtdF91ml7mWYzP+xHp+VYL/TRl9ABFF4R9NXDOMUSqeLy0FrPu7af7sg5bnEWLT
e39Zmk1BN97hPU8H+nK3LggSFPh1cdIjKPoL+68uMAz8C/PI+dMw2PdsH0v4LFio
1fMt/4Wp6OfAzvbPfqX6TqnKld8ba7unZQ6wgM6XQwWWq0o7cLmS7Z7pbEv9sUob
ab0RIyrjLmyZCLcQsf4xG2X3pmCLnGvE0XYNM7ORtVll0744C8F5dUe0OtIoqMG0
eM/xXb50Gtzaxbj9iL2RZOMOwjbBq5LiHqLMKBxZS2/bDrb+r0PjX3fQF1usdi30
hsz+9YvhOpgnZCvnN5Dkaq0LQua8PNUgs15zdUx4nWhzI8ZBkq3h/RPEGHaaktWF
4kh69sgq2LluUdN6fEA46LGexWcQdk5l5ABmMJHw8f7KBj/oo8l+dhlzpaXHpX+J
gMbtc/Rg4cagep9/4MQIwHhGHp8HDVJXXNHvD8ePz0olcX7SqizZH38UKU1tmU7C
5gge6VN1lbIV9d23JIklRed2DjCizuNKDQ9iiKF8OAaT8/od35cNpxzyeFeC2SVv
JhEYf+aGzk6TJhtCBkWiicCWozvTCawCZMPkxk+emD5nHtcF6kBYtM711wNb9rDz
ghC33t0GwbyG2Cc5RwjnqyDZ9fw6g+Egb524kF2eYtYajfaN79OINzmXyeUvvXEK
RfdJxQQzEf4oQVQYF34U1lQlXrL8J0YQuW0Tg4mugqA+MfbCve0ti++SC6h1zmAL
9DP2wZzs3357JPZcY3pSfmPf0B/v5/HOZiFOLaIxL6PuWbBtDhqe8b2uhkA+IGTr
agHdSCKJyiWBhwsB20FEjofd+ySji39xyn1v3w84XUErS5hqXiUpfVzheP9xxQej
KUxZ5/OpzLOd5G6U6ef7mfoQ4TQH1ptZoJDhijOOzpxNTD9bp5FkWzqi6jJ3mOll
GUDX8Ff+8kVey3bs7RpKoYrnMfzipp9ki9waqEIgiLBtM9q96Zt3kefMx54uhaL7
APbQthV8/MQnf/S+nwBfzzcQw+pQvU0++5GDWVUqejW1YxdAXtADWUIg5E910P42
WI1xvRj6uK+pIT5AqDDeaDx6EUrNT44XYB35elDgtetanrdieuHdpWiHwPk5P3yi
jHHpcP3dqGQihuNuGgvEHK4fFsvHO65VYnEVkGNYplOtyc9qVyWosgxNpewJNscb
2z0IJsp12jL+KBBASFHGSDtKSx9F3tVhO28TzzIyFV5KX/tNHmUIGu49cMLyfh+p
oeHJ04+6HEYBnbVDj+SHW39xRMKPSeI8SuT1osXd76bysxeWIpD0CtR2z/ksjrJp
JrIdwbeotGtR2F7wRp+peaWHG0ar8uGacy6C5mo9zRleCs0reMa6dqS4Wz7nyx27
ElSs/gFyfljmA3VzAxVRgU/kVGatiadl8xFlmcp20C+DNOyauxAVPSjepW8YhULc
n4XApuCPquAK35P+O+dqFWe+V+znum5g2LdIumt+vk82AMRtZoAaKB+ZUT0IjJjt
3RNuAvLOmT9FNW8XtXAkY+6mKmOfrzsClApjrXuTpzNXFdYJQpexpCR08DnndFAb
Bz6FVW8MzCdHPnhVedUGDKMFarJviOp0tlgiFYAwvZRv9BgvhWqA/kA1bgRMVQyJ
5N1tl2UVONvcn0nuHCWuB62YyKDxpCFED30ehPXQJVVM45oo0YGFYfHhZ9NwEs4s
5cZVHAkqrImsAAgwSS1mEtljjQdaB72w75kBe5G2TXqMj0awrUIA9KBjPkvZbBtD
0Xb1wEI3C5nVnn0OfWYIsc2PujLHyYHjDN/MMM0BtYC28hwGf4RNZnbGheipfTOe
w/guCJFvByxDMD10ix6wfx3R6lC3h/9vqfivcf+OD9G5/yJpVdKG6cLw5+vA8B4f
h04QUBVX3kFS8F4L2nfkT1f546zrcEhGrTBoYK6pVFNXS8VIuK53wUBzM1rrBWY/
IOhO2TIqV9A+YyDfsck0oPFJutJIClirTn1h8Y6/NSIsQHHqLmmTH6BDIjn7VruX
865Ny/jE74nWsksPGU6oNXDFsj8U2uuW1G5553tPzXHtANlTZMp37nAoaTPT6gFu
XZ21neVgn57RjJHO9x6tIm/XrU1Im7uNQ9H8KsH+FlD8sbmvWCwyj9SYC0UQOM/G
gKKfGro2Et2HknFSM9Z0J9Fm6+MrINWFs1UOm+rX5RpxEyVri3vfBZUMzyy4fBZ9
nSdTBZ28+1OyKT+2ngifwrUc+gTTDu/WF5RbzHMckbzV715K3MANlFPmI7TuhOg1
2gXOh+5Ngyw01IbKxfAna1sa3tg8XJiPTooJRxFcFVvhDpoPDNoXcO8K0HBIs37a
VpkML4tZf3KXmQWvDHzMvX8c0TZUymboVNrcX3KCiSF2nhtsJGgI1xUSMMIRRho3
WqnQrA6asEYBG+JJ7gwB7hENywK7Rlmt5u1jpfUtckLBCcW5ZnfrrjrC0BJefU7b
vL3VckkNsg17sOUDHyjDGzGYbtkzN/wp6vEb8W8/2Rju2x4kKMyrMt5qlaeQqWhy
lKSn7RMaHxybhAPVJ88/iSCFjYyvgAr3GL7zHWely1wyDdxShMLZ5lMJbJtdOIcm
rHir4/cmMJzC+lex1PughzMecl0XlKp35YFZRefeZWdIAImmSFSOnyZXCqVduREg
qV9KPNNLOVLa3dhALR33moF7B1yDdq8xusBWIqDQNN/ZXjb0wXI1+Py7knP3N6Yh
E5m/H4oN6Ot/ZlKT8y5tk0cl6G+qQ8iRr/misOflFxjDXGIP+YecJgmPmNY25XUM
OQ+GXI1yNQP+1ls/hMPqLPdxO8V2FET5YJAt0XyZgtT4HWUe9cp8ScmZWJ8WvV3T
/l4uisZhvpJTJBhuftWEo1KGd2tJwgje/OI80IMEd7s2kToT6HWCtWAmAGTR677X
hqhZy2GZR6+ZDlJPFBDm61h+3HgZBkdKwJrU/7wXEa6S3HxHY+ro7frASqO2x0+c
MHeSjmv4IS6j7gFTxVd9yaX/P0VlpJGhy7TgzWJSw1BTkY0xqndUx2kyjfhd7RJ/
O6ViW2OXJr8RJJetOlOjAR/dwg0k91+4j2h5/uXWxoya+M9JpWrtMovO5jc7paYx
ugjMBrLjy8dylJ+Ms8oCk573/ofGsIBYocVxnpIsf3CAtE68F18WndqWj+nfUpR/
iTkQinCEXvgXddYpEEBYiVqqm6WbLGjF08qcmIJkedzGdoEeatNYLsazCEL6F6G1
Mx3bIwI0j1X8ZeODeZNpKMXPO+AzU5i3cunpvrahoTN6y+NxvJVYftE1hmrZ3rOH
vgAKRXsBY41zfXNmajeCl0wg8IKZpKmH+35w2FeuowhyxxQsSPwJOAHeNP9J56dm
NgJM6zCXydAYOiRlLyNReCKKDKIxUr0HhN5n9vqu8c+nuvZLATKi+H3w2gNOOSCU
ak2r/yU78NlVSJfF1xZeT4RL3KDGsnyIS8iDPQMnMYnNmcvBOrxxrUhzB6KJJ3Yl
l8lyCFrGx86hQgG1CmfCK77IBPaqiaPC5lGO3pErFaqybn58DS1RNtjtbbbatkRs
/oP2ivwIhVVY+HlHLRx/h/pxr/oBfNKpYbyu1XmIYcRABCmbbHCdoj9oWnCGwZZt
6tye/klHXjPFo1qbH3yWY/CLEDrGCDN3VvGsIdkq+wzaPsAu3b5SPnyDuWA+7I35
0jWsHRnaebMNpFx6NjIHZUeSnreelzp+gPCVm+qAcqBUk//tFQwyHUa1eZBGzuiO
dM+GwHEbSgYhBa7Liqi2SWJ4o27MQUG3dHwv9C7PdWlBJCxt5DwvAVyy9MldquD/
atsGjYcK9JjPCz8FrAmW8z8dXMreYlsEv9EuYqGRgY5XAdW+x6eWhG3GF2qaXU+J
EUmPLU7H32bvmYIJvu+3U9NnWy2GrM7BHH3Ab9pl4YpFb7M3m1vHIp9ekO+BA2xd
XWdx7Wx6DK/Oo35fY7aaaz43dE4wM6hmp2TdgbcyXrYw8deWINMjXySxCDuwi36J
HydHR6Y9RasWaqcISrXS/avExuazy+OMb8U/F41Fk/fcI6xAH1yOWZuvxZUIyHxn
Ln93A46q6FjNe4xYwQ44aSZUP+T/mKT2uFs1X7kIRlTKtqSG5Z+vFocZP30WTd6G
GQ2cLRh2WUMaJAk1NJi2/OEtuKj60iGKXbVQqfAIopHxG3nREPN37jRX9Qqdvi/6
qV5aepQ4EH6tXKW6sfaKnRFL4MI94Z14WY0I8ptnPZRg+Q21HYW4k1w0OM/dQ272
OVvu2Kusb31RiCzCNpqV3kCUDFTE1OVfGDwrL7UT6tgitiX6ENHMBFqct+eMQep8
FkVvHt2UPa1dsCT4ojhFMUZAgH4LjQQS+1aXlKwbpxxOQNgJhvmtjQTqlOGo3pJL
4I7NUPhqB/kb0d8/yEbyUz6jyrBE0TLrK/m0sGJSYQgWpGIRJ/Hn12Y7dff4fXle
ohZQxu4P3kXljJKHaRmZH0XQrDOh9tXdYhsuocdOdOc+/jjikDX11PoV+LMYGZ6w
mijOKnH5ocMXXEJgCjUa6Z5ekFSiDTRGZzO8FSRmdXwxACUzq9ehcDo+iq1ZBoVx
f4HRmYj3odO1+NWwFMjuVvWK6faE6V7fZUZ3lTf4lZatg0xJDYewQ9tNUlr54h4k
jqDm/Iyg8u3ZhVO4u4x0sZkXsxKGdK6j3uvixeQL+SujWztQBAauZ3ks+RvyLxUr
SRwuLDy0qXUtQ2jQ0QKuDowdU8qkFaUIKE0QHdbFMLjpp64dl6IR4Nc0EgaBFVCm
ylqsq6xH90t0zj0KA45lwnEIkz59UgwY54t3nnMmQJRKNvSsVZcAzv+nsCCWft5P
RJDHnJYGrb6G+UGS72H4B+ZFxri2367/3xemGgr0TysiDDrIIG86dOycLpUlYVPM
Rs6AytPWaymxIdHWv8R90gG3Qr+o0GDB6trn9Pn+ZsnD8mfrepUas9owAjbWcLe0
eiLwa4v0PVYHP7Qna+Faw8n5kaYBMBD9Usv2GE88oFv9Gl3S09DeFZi0BsiWSTfY
vMVPk3uKe30NPxVbS00JCtgHZtu+h1WDbT+X0HkK3VQ9eGM+VldWfFfHymXZJHpz
t1wJ4R3y1uzHMym2xSwHrQT9AmdYriUzXl1sp9+HwU0NSJL3GzUOKSGg7EtWceJy
LH7Cxw1bKSceMy181hdDCVF1aZ/Hb/Hwc0+NJjRcCbOkUJ/k8HH+vHV/HK1kjci2
kTmjAgYjRfyLp+CM5L+/PivZdlXn1+GHrV43R+Sb23ugLD8x3pbFgT5+TIBwpAa7
jMIII8xz+gOkMsVeLaUKwjbyFql4NIcMVJLznfLHNk+XODgknoUOa/7dElwi5Px/
qavZ9mJu3cQKJudvzKGR3WJgLwVxEyBqVfkI+VTVcfMoHGZVJiVLGL93R/x6LK1u
gR89UBRPtN3DnYqB3fmZk4BGQrvXtv7bg5hqDXb/FP0u8oGweHcDJLPhU/vIURdg
rRG7ILgNADX0jMViLbf857GW2HC89pvkdtkGOYqic+mpPawc8t4JVE/P2DzbU/7E
Os5MVPzVXdKsWGDCDLU+QWJO+OaJZ+qR/SSn3oDx2x4m2Pi9YTZzA8rZ0kP1OEy1
bu1mQA5Sp9i/sf11ztpwE5J0yVfcLmw2wAk/FLmYyt9rFOnv5Jt2G6M+Js0Ap7O8
85HarQw18ejT8GUSyDbzf+m1LOTgi7ajjQdu6NP0fBnbJyNWHyRjBWvy/Yapoco9
25dFCFQdi8CDUSbq5HwaPhC/tsHN+YJVt++pXjl8EpBwS/sPAn/NKvlX4lQp5hY0
oSBl44sG/bHvpN9v0qyHjepkGMzwKqgCQheUo35nvN0fyDZnxME/RMGuAtRiwDHW
+Dtk8kt3ba7ciC8qgKyN4fS0AMnLarwEtqraksN89g6ojeY72aCG7XcAuRIXkUvL
Gjo0PZPoC4sOgNX+xiZ900+FeEqLLscLIgk57QS7gnZHL3JMQDbyOcAIRZid7Loo
mz+pagl+NKPMGfh5WfFp7FLEvETjGSpf/YxjUJkYY8Sm7QMgUdX9fr236YxEXgYU
CfvYZWrpER9+yd2N1MXT9Ym3Q5lr1VYZ1HB25RQH/WX5Xxi+wr50GLgMHuQJj7Lb
5lx+lOGGIC7UTI9HYyQGL4GGTJQFzevdiKXKiyghWCpVR6mU7kJtgka1FhR9eygL
3v0/YykQycGoOzD8RmBitNBwXKUD0xDyxuFJD8MKRmcPaPixnCKiUHs13IUhHkI9
omv9MPGFo6XTYiu+uE9K1DSMgYsqWE4/J0YHM163mLAULIL6lHs0FyZ/KfCXuto0
w0gklRG6gL/TW6ggYWpFM3zhr6qSkGdxoyWHyWa7xcold35CwTRxfpZpzYoA6j86
d3/wUB4+W9QIQ67cQA3b4McPXAzIB7lt3mNN2qHwlY3qQXGRwp4m1rL7BSrryxE7
VICAybu9EhMC8qd9f1aIuH1k4CO5xyBdeRS7BEft/SAU7Uy0IvItKhvX2qix66VQ
ZdqYV5Ngi1Klx4d3KXfe0bSkYvmmM7Fidlqyt9ncX26+Z+iLq2XDJcXL2XqiI4kt
2eH8jLaLOxgMSd8HALBXFcVKfUCC+MEbvjLKK4l3uUf1yS0QYFZ5j7rXqjcb7AqR
zFa3BPN2NdbPiMUcZfyHxcmQ/zOEptx4SjzYWJhXI6M9nhhDMhccIs14Gydfwc9C
tuHdQ5RU9R/wRujyDv1QDWn0bLGKm2qx2Xm8RjivyhrNxfPgIUr0OMjIyQIUpCD4
3Dwwe7EaiM6dkgzxwAt/73h5o2+fjurrH/LPZHEl4/ATRwluFikbZm8saHMa1pc1
LMpMw6WpEgbMOACW8N+1QedRbRhXtp/JZ9qXhn2k4LR7PijfWBcHwXDGGfeCUBIM
NnODieR5+fhRgLPnNvqSndKIXRj6dPT9kPEC8EhJTJLXtgBQECiXjMrSakh3b8gr
wYWDXeCeh1Sg/5S2ILR/jtKcWZrr6k/PQOMNyT/dOkY1ULcguhNlRcYvYTkvoygq
VoVihCFn9+O0hhXaF0Bhf+cnQAV2UfgzSY2bRMcIdXCpIzV1fhbBBFDfESROmlHW
aE9nDzo3jWKIsMzAp1zCtG2erBjywnT0DXC6x/TSQrMBEZxa3gJx4WDrzUPE1BDq
N9VWZw8AbqNt6RWfsyofKgedtJ9seJZ9SU8RNCd9bPpWcv4F7KxA8WW0EENtZN1z
4mlBQLC4mJSK9MfAuEX0D1tEcNEyV5bgF4scER3cVLQy8scpkUY9cKYQ30j9eIaD
Z8CLkTKh4lPckjnnSZiTu2E0n4/2MPUdKSGFepwXwMLJDuXiARKwd1uZYRtH47J8
orB7mKYouBu48ClaByAQ/b+oPlJQbrBZAYwcwlwiXMWFX15bPAXZ5P4AWt2TiLU2
/eVujvag1VdmPiGysfWkSGSIs7EXI4HHRN3a3yLXTefd7fBAPGlMUuRC6Mv0RO8V
rKHlKMvwKGjSBIf3tf9IQxo/nJLw3pLWfc/XFAP0Us9IkBO5tBVAp53UquQJkNC+
lcjgMH4mEgEsfCpxtjvwMLnQihUG76JWxc0rY7qLveRoTGrRH+zlYHNO6LohJcAT
QAIPvPsxVV7MGPgHD7IGDg0BiWu4MuLCEfv+55Wk1MSitGgozyFNMQnwKrxepuBS
aPxDUfDGwIU/mtAww7XulofJ4tvuXUljqOXwuALSaIhuJOUePbKGLCBQlRhqPMWZ
thpLdOnBlErEtAZ44pG7Ll7ISWrXgJIHKCKmppxMtsVPESt1G6CZuhwD6QFH2J/X
zti8iRtRT4cSB+9yX+PL1fzmg8mQyy6Rl7x9rb9Kra5xUGn/mAW5JaS3vnvqqaRJ
y9q5ovvCxKla31VzVG7N596M0cG7TErYACdMYz2s2RfjNW4o1wV6nsa5Qj4p6V0g
IOT/y5kLSqSTBeYd6XvOn0SaFxXL8e05e1VildMH4zsjjyCJQHRsvFzaEzH2N22K
3vvoll8z4ctrQdf/lPziXTADFmMLDcuwUkXVfHI0mxlfz3jxQ8hi9G8MxbMKyoto
yXRjk3AMnuSB76zyGvw8MSUkL1gchFbMM6H5ackvcmGURut7tpykjb4P2rAtdHRH
52oxMGygqvLn3lRUdNm2Za3NC91qWS5kGCXLd/l1tvG8GyhyaZpIS2HSTBCPP98E
kDqm9nxkSftpzCCnZwQmiL6pE9nauP4gGFZh/Ykrp5aTxbKmMz+sUWUf1nVUW2vM
+lT8oDbD8pnbHNDvFiTE/ThQvi8kuQFujiaT60pFUImlgPUe/CcHFakNOpOjXeOA
0Tpo7YE7cALUFfP8gFUSLjWjbVfQbfH3GH1PIjyzuYarec9mWe+K2/AIGXn6Se2N
LleACxRzcW+2sTc0COvP10LIMFEWj6mgoSr2Su/cAGJuw5usC/i459FTs3uZx2Pc
/dftRqu/VljsC/xWDU0P+1+/mYI1eFX1/ZpPP63hu66FlaAzKJIN8ncU4dXI3HLv
cP3EPatHG/ZXANRA1dBko5uoTJqsIni7YzyaRcYLqsa6zwo1NpVo7Rf+eOB9I0GD
uG7xBjgO7CiqnVttoRTC0zKXbTNE2b5rsT5670kNXdoh12Dy9AsApojtr16pHXeG
8elooKsHoyaIHhNAf+5zMdDWQUz4lrXH50huQxguupRFrrhahVHC/aM6hFmhf4+W
N/onCwkiMd19EBQ2WjC8Ao/FZONkn5UgRCca21Xr5sB8gZHvK0qVcy3kdh8acBr8
XKVOBzazaRkmS2SKecaxrPmLY8Q2zuTv/6PuMk6IkTTQ4Q+FgmzEvE1txjOKsaqA
fjiWMiBxzrZblDQ5OAlgbmChEXxFj915rkOk5jJzu4vf6q8BnkwpEWMAwXVuD4V1
lVMUaui3Xz3cyXSgIL8zvYnJEcaLbC3JajQvOZ+eg7u6DqpWWCftkwDz+W6ICJTa
NvH1XCSLO8OR36pq5Yq8wQxNGyjGRiSq+LIhrtqU0KHadkURMx/sRp5MWAVpglyg
Tc7MXhAMqvOw8fyxP8wi6oHIz7kULSlvP2Rv5CtRZdx0BZh6xPtH2vDJyBwd1R5M
YiPYnfqXecea8PhkIxuxVgxWYsWk9va4Ei82ioqdNW4q2TSbyIkkIk9+hGv9Cf3g
QwdpNS0aF23vqBGyH43zijs3nXt+hMQaulEnamEf8Zn8eEFtbV6Ja3GilZs815pF
q9rElCRga03aB507Qeu3Kb1vMiVp2kYKWadid/E0iLc6tphQa81ZmBKEJGYz8cdQ
MBr1+jrwC93o1IUiIG9APlu2VPU3geq554DeN+Z6uDAZyoHGRdv0wQNBdWAIc0Hj
7r7T7JDrr7PtygRZHWXmt2T/E3RSiWeVKzTxeR7Z4P492SMR/tNpNdV49vxwYxzR
6k2Y1IWSAsAr5NGyxGM/pnPTnFN0dJs8x02eU2lh0yWsgkdc22820dlV7yIQOt0j
w7AaSXZeUoJwa3mflBLLOkXWIyHf8rSgMp5sakBOLOXedDdMYv8PAICflpCvzI9N
R6y0sWGgSjhxNrt8PjRohtX9ikc1Ryh2TqrLO+fE6gG8frGV3U64zoj3fn75x7ni
vguef/hh+7Pg0daL/d+Mkr12xDYViEwq3ylMU5Y5b6iWJJmXQskoUc/YsQMVaMqS
zB8sKxNwbbL8sga0wjik0z6M7N7r0xp/7JOq0yXIG0LajJtZUsXCPoGv4RPO8M+G
DQ50ZQ87aratQNrbzIWQPH5YhPKg49gyfftzX+3Q8JO02iUG0/Gy71MssO5IKa5I
iazZOy/7QW8RVb8NLLsRgJhs4fPoyP4oCQrC/KV7eAeCBS/0GN8uEoyuYBHvI8uN
T/3boI2mfeTpiFzCJmMOkk07lfb140PeaRehl0TjX0Xsu0xCdMDzDwpLZoxv8kJw
aploAzYuskuZpRRYuvl2F8nNdvNJ/kqbZiy9WgKJFNnu8TzCH7AoV9EqPfsTmvvg
e98bDh08vYuoOyfdzrKmoUT33u+tPVH0RNQE0E6nBJD0x2hREP0aQP67EHbmldup
0Fguwamce7U4Vkfu8im1JbGoZbcOet9C13ByZjemPL3OqQlixBq2Q4dSqEheZsuC
G6Pnc92TVplL9cQeBD9bXdGpYAUOlRqXGrfeK7b7bdLMTimroEWCxoHnscoy7eSb
oyDlU7RwvsqJKqPRXgdo9kZ0itsW1Mc6FbptdQtS6dExhJquh5QPbY9H9P30vbeW
B1ufaBxG+WpRUqljykxColaiFHYaI88nLxue2pps12xGDFG6xh9nED/jYiwXjJUA
7DBKrHgvd9NuEungl9VDsyN2JB20P0fFDFC0yjlI3M4dtFcq4m/FbnwiFW3ABBI6
4jC2l29gCg2XdhRJq3jJwcNMfZllTbBDthyblgr2BPJ5ASwiTjF4z2iPnh0SBu0U
K6dxKFzI473lhBUIN0bNW72MjW9k7BWPVmDLkmonQkdLOm6ojaJnDUfBH0pjTBPw
Zb0suGNmv+hezzIfj+XygFI7j/l2t4gVaTtv72ndvmq13szQYmmAyxIcSR/wBacB
mXQXK25fHrorVWjMah6E2CYkxbBH5Jmfp8aWtQgZXyeIdqvkskxx/ckzKah3blCs
ZqVosh7H2kA/MpFAw31hNAf9HsDrxZdYIi6KhQYN97t1SYd+YI/1t4ifpwSY0n7n
AnAtkKRBhDaI13i7aqi1VlZzueizc0kSwQXXbk8avDJyI0h2JEu5Io2YEZEHSvcf
G1wAlLXKDEjtyxz/Ft3uBzJZOvvBLKQqd5GUXwKCMMJvBwCI5zne3kcj+3p6Uhr/
TmP3lwwGojkLfktR7wJKdnOxR39nQVPZ+l5B3Q0pj/iZhkUmeU+oirYzldQzd1Qv
UEBAv5chbiViTEG9WpKKdJUhyM8OHWg8h8egZj3+TU7luCZ6u5RjvEZab7F92OAu
iNv4DreRakrQHa6X9Keao4T4VEl322i6mAwS9hBE4LhRDIBfnfACVA3p/wg0wihU
diREuYPFoy5TWuuvH/SYdtan0uzsayx4VDF8m79KQT1JV2pSGL9snnqTcHsvKFzi
Sdq2geV00f6dpofA6VRbI8forzWAhSFl7GSR9BPcjlBGU52/2Bqs23AmO26mCPYz
nRonBI9GMac5cQCzZvXzSzVmikWm33pkfnvRBEs+vWK8qoTxRMh+vkrzf+iSSjnF
hdkdArxWNYPd5fOPO2Vu7Ym8xvSEEdd7hPDAcLgioH3anPgR80DrziaNuc61chpv
6/GXuU9MOe368ksSP2nyo5ik0ON8h+lmXK4cIt+scymM3gCwWyVV/IFC8sgX4kon
PhdHsNUlLuBnAiv1L6zWIUTtbLhMhLuFMuRsKqtX41t9n4QQwzX5hXmgaBb8XjY0
Gi7FPPelDWPsglNsfFo9+BPQJSdaeuey08ihNb4LCTswJElVIhcOTeIHazEEPSeE
ZdB+By5aBDoU9trHijhk544WjTf2jCayaN78oGuJNNTDd1Fhoxk9zoXJpIrBF2mz
UzlMuVYrg7pLmqMh7Mig3rbitf26f5IgEppH1Gi7anLY/bTtnIAR5TqGmmrAvaXj
vA/TP9d8ZjKW7R0TuK6SoCAQHp1EyPBFz2rDeestufLFTyteaL6qXh4gH/lRd/LP
mAs0rzPke9P17JqjSAKqxmHK7HcNk3ZnK2mswEdh4oMaNBIbe0K/BQbXvrg0sIIW
HMILaS4yUlNZExu2kripET2bJUcra2ha9U3KiNc872MV1k8BdpI3//Onb3JJEpd7
DKHB4OIiyv8rScJbx150uVb9c0DT4zmI02i9NijXsKdxqDDgRmjfejS1ZNTc0JlJ
DMDbrEHGH14XJ2/mzvtd5ZrtoYMjbSV7MPvyQTi9Frv/YQDpOjKhr/iTqJTPlHVl
vTO4Rd2Abd/8z4SJQu1+UId+KDWitBsVGDAhKtMyErHGBcDfQM7WPtFYg2oWIRva
dH/K5edX+hlSGelqDMsoKlNWg9X7VMnJFVzws9ZkSIH/J2pMT9Qyj4iE0EzCsEfM
oig2z3tIDwWyEOgQux/qn8AmD51xA3bKJyY20FN6mDhJX/ci2VQK50kt+Jtyv6tH
88Oy32/fqOlU2DREkcPePw/ce9BzUR/YaWfvfo/5h4CSSeklJfLYprTGL173CQdr
PQrPLjxKC1Tzq8m9gIAFpSoRNqI/vZfBaLDpnCjUDwHQ2ow2eqkHhulyxrlzDxXN
KgXSlpro22SK+/LIejsoT/NuFlFKnPWLkJt4MsTSpeXWB+6m+BJSa4IpT4g+hl7G
Lss90sXWaO5KS3STAW7OWEH2tzGI4NKlwFTxXBSD8I4kZ5/Cs/7h3wOl5edgOdUy
e7yejoMrFbm5BpZ3q8HkGz33Yz2pi2NIBL/4WoWUHqsaSbpknMtMs5pA+9Cj8Iso
F99SHiWQSLL0dar52RT0FgBLhvNkgGBzeGNBJWiP94tCpoetARJkO4lAubxlAPUq
vJNNXFVQSniRf5+SwAF1dy0yKTBiSxa6ZI/BlJXrAlGSfL7jBJ8dKGAxPRRmIHpB
IReExT1IzFpicvEnUcntQ3IDyYmcuFpU2MWNRBQ27US9bjN7M4D+Vsja2MN2khal
NQuzn6Y3PYTSYreKdDwx9zd+dI2gI8bREsj0tiu8HOOqopmXBhloh1aUBQInDiaF
3YYixRVQu8bWmWKONqKaZO6VjgO+Qrx6+VoAr0h7TtXbOWYtYU+sXtzrPmMcprof
rOIu4uhfLB57Ne/ka/hCJr9/8FshIjw8cZkRyEHyAwL7ocE/4zaN5UYKyoWtZvvy
+dij0Z1+oZ3jecvmgAPhWSPzjyIu3C/fmvkYa2CzokWgvasOb/yfelFDocYQqU5i
32Ci/80H1NOo032fNnLprUQdK6/spSy+OC4pfHYnpldLTMoh0hz7dm44njM4daS+
ZVWHgtzNsHRXxov6XjxeaQ+E1u7C5zC46kTBw8woBffzuYX4PwJuQ2I/UQy4Zdfw
05dXJlUv11B7zspdsNEIWAjadorvcxkEFx/Yw6mUAiPm7khsTW2/v6FedY0OfVEu
kdZiiZlIVzC1Bm4Ws2NoG1GzsTnHcSHHLk54FCkJ58sfNyzfm2OeO5wp7BgN5Go/
GlyngBaK+xq/B3OBm0pbordPUtBG+gF1+hIiD6uwdsZAFR+dhxfqDUyC3XBG1+HL
hik73BuK9BWKL/5gslhkPviK1Hp7Gb3d7K2+ZrBQcB9KXnD9eHxohuVCOJnMmZrM
8BELR3ESepAHCv27xbqaFIHVzC4ABKFEKxblLWaFT5JqOPlsT5lhwjEejMB6/jZy
4YtwPhWOBstMBRIrgmAkFxyjuylI4J6Ec/NfJYNiM0o3OrzLCsjmpEjKlR66Z+TH
YEJStnW5o8J4wiMSkPb41vqHTt5saJyY/+kwP2BrQyKaFIMkHoeddDICb5qRfOx9
JWEPtDQEx+4Pf8xoXfzF4jS1DGKyqmd6pgQWHpE8WOKxVuK0Ew/01R0kLuUSorwQ
rnHkSnzRfHVQBedP4pBN2B5Ed5MSBtnJhFqGp+qXhWmqGeHvY6wCfuzdzBWEj4GF
xZyFrJIhDFAqQ6E6Pilbg/aTLbtGyaf+qZo5eLoVJqGA0MPxl1kESQMzEaQpjkHu
YhTsNOJNbx1JMQadHWzJad4EkhmKcK3iP3lJkV/962at+7KqS+vlRfF2idEh562f
RfJjgxZ98Lid+11nK6WQ0ctEStN1orUUb3CENMd9weKHCi2Jry54Gscmb8dPGZn4
yyEk2d3WAXOjZWaaYuzc7VvezBH1/Dk2xp39498m5y50n5T/Znmu2amHUsRj+CvG
egx17xdPIZO3aBKddkcAAFJjWd121UrCYGPXeqSkoobvDNS0PYq1lUO0c0rdz+OM
Am2HEU0ydWlLd0gYIK4p/9sVOvUbJj92e7dzuGtlk7PUI3bPNGKMDu5a/VvrTJmh
kpHETIWZugGIj55aX8qjIcAgyHyvzNaTiv5uNTlx/3XVRXCccVgaCzBZQ2mg4/cA
GSEFMaOodWvgWfrtVBeaxXRZIRNuUeQZkaWpF1gl/HiV93uTa6W3KPjHebSpSPbt
X2WSVzlmE7v/cTO0vndecxRRc2GPaBoZEe02wfI7fpcB4mbEWoEzScIekt8IHhC9
YUHhBl780uxxwCBqzSBUmfSDvwLSmTQYr9SK3JHKLcauxOHcRg+WRjo7zxasxOXd
eQXqnOMg7n77ae5AxH8G/56cDplr0+7JvgGYb+87k0nXfbhjgk5wHK+klkb3yLmP
iBEN50voRCcN8TueeRpL5jqRNEAQ5IjgP1F65eHlvb3QgO9oNZfH7TEAaAOQR3Ei
HjktFsFFeS/O8tWq/6j1tuSk/CoGP4VfQT6KrE2aIKjUL2MHvQedxfpXYcxGb+GC
jCrRL8fZbvnDYHZoPa/U4LLrnafEVECAjkOW5AcAngLT3Lsw+Jz2Ani7ZaBxIFWS
koB+HtHiAikagmaeLSEwO1wSOGG3LHcjmjjhY52ZUb1X8r761xatNssvyPQ/xq4V
8+fEzmlvNUj8qR3xZIwtBXwtAJHhbO0jhM8D99Bb62hf0g0ugYhRnn+NrT9DpYJn
RmVs4J9OPYNnay54Z7yqXHoHtZqZwDu7xRUFPl16ZwlIrC3FyO9VDIZXGDFcHHIJ
+liVRwQRrBaRIyLYTj5iAfYt2tpN83iH1DMOiwcqasBNqsPbd/K+L1dESESMI3GX
Es+NcSFOsrcaqPeJ76mSZEcBF0pDiHzmna8KXMxJyxnS2vAVB19Xh4RTEIBBydCC
zrJeFJgQpc0bdR+F14ZEZgqQ8c+RUmIypQfmGYj7TuWY3N66AMJ9rqvBSx5XBuD8
8Pr8oLWjSqhvzNWNmyMIGCV9CQqzgbPfWwQI3+CjGYgKZwqwqrnIqzEp8ospy5w5
VrukG8EaHX67COY/F7GGqDuaX6oLqIfOE2H3BdBoieDHTNjc2ObH08XeEmyYbEVv
7Jn+mQWa4ZYIDom8d8IDNz1whU2EuK2jzbdGHXelczuMznqQkv/9cSv+I9XDYyxX
+1ZiIyef+I3CVIRe4DJhXmsSDKql6Z1AFdQDyDswWpb+Qg9jOp230Z7zz5McZurE
YlHBL5XU5wDykPDmBPC0kXwIEeBZTm2CEMh7uiopCUnssjprg9jD38iNArQdLYR9
rlcrcI71UJ9cAI5sYcxL2k17nhWtvD28fDjbIFIg/1XZ5neiUd2irZAtB/e1HrH2
KxqlDByXDJoH/numJukYZT7zcLuihF+Kx8z40hPwfmjhHXqIEdF8r+QYD2wmpgJs
30C7hamMTXJl29PN0U8KvkDT3xYbJqFakdXW49+kb7CNckHIX0SlmZRv1OMAcR4y
G92TXhWUzQ6UiKLyGr38QH3sQTFtbw2ZPKABbSqRw95V7+d3TsXEMqutuccPX2Z5
ij2nHpTg/RDQ1mfhjmOOiuq1fYfw1Ck649hVp3/pZf0LVDn8CGMgDvppq+QS2s+j
besHZJxvJObDWlTwbl9FBPPNHtR0edtqAacJvFvDiqTHynTm61cz5pGc/FQEwmi2
PZWxhN2uAtrgTZTmWb70h6UL9hALM+L3wXIonWt80JnsHOxiULm7bAWoNud5APX+
NGBbSao23uBFdX9Ftpfig8S97GEnyE5wX8zrRFIKv+mvbHgSpmbSl+rW45XLbCXc
sHpeD96B+fypSwmFl1SnIR6/Pb25TrFWwcSeG/+mu6lzv3pFa02+H2zc4OTiiWvK
q5jnq6aBysAwnsJ3B8V/8VfxqHZiAHT4nD7CPF5tzpilSbCQyQfNozqLOWmXV3+O
ELS9R4Sruc5AYfhAmfOLEnzakPaDq27Dkt+W8eJdPSeW2VK7WLZZWMwe495zy3Zv
9jOq1AIn4AyO3fAGdtPyo+9QjfAuXuEOXhxiv3xdmXKgvG8lvafMuH7RAw8NNA39
M4WlBsQV5ADDszme9gUXY93z5XCDSyd2ptiTXCRwl1uw2pYXRyzvOmS7GuRL6fDH
UW363QXKVejGAoSgVxzldr252qRK5f8Ff1aiSVN8N7aknTy10aNytAlYwYN/yyFr
Q29SvFjOsGDBB05DdQshM7+e1DaLntRFaEHIfe4HuFWUmWAnH7YK8Dc48sqOStqq
nqm/KBYKarEzhmu3KjFs+FAEmIHtTYAYmXTZF9mwlfbhJxy/2YhXGAXWMNdJTQ51
OYKZbWMFZq9NnygEbOlYf9YtaFAAPW/Nyyec5uUnpiW1DdkSNeXXQfkXMI7mnApY
3Euo3fdLSD+z1ZpN2X96N04ed+SK4LMCqjsxqQwTuKjpYFWRPbJsf4L8c5z0GSrN
pc0lsQ55d3Ac1VV5P2nDLMm2Js7XIE8hh+gnvTPWDeGtxJUpg5QZ6TuwygiEPYuZ
6pmqXK9Nv1OdaocQwwyXDHBpnREtQSEqJjreJ/BcZbX1TAKEwmN22dtoJ9IzaZ+P
MRCgrW7AgdvE6CCR8NXOuCw8N0yP0BBocCxB20O6iIxDlmEe30y0n4zkZrwT8kdR
l9tJDbdXQTNFHodNop2BzbnSgJodu5EDZvqT6tyYC+wI0T9PuWzymQeChkpxZrpi
3fXnoADO5drmJNfysUdFdqqcVPML2szFv6yJXLqRfH7EHKZN8nKVzhK65TB0bVCf
t2NRZs/AXntrG9WewBwLh6HkheutodcRyM/clUoKOW58RNcEihU7uJe3wI0Q5nKz
raj2+icpvghAxKRvGSkFEcZAOxl3LkzpevH//Mz/MX7awxXgDHbUQd1r63iE9YEt
csLMVMuntLNWF11qJU82GNBo8VMZ/hox4Ps3k2kHqXEHQ1/zcW3nXqsGBKi3V8e9
JIn4lvTz6peiRiGdUsNBpGOw5YPP/FWV/dlvvh38Qj+Zx0b6oFN7SSLrda5sE0Z/
uTkgWAcRFSeSKA1mlmS87hA74NzMAIo7dKlp+kbPoYdRz/kUADzfdZLkB4TVQkUM
fN1i5p/c3+4NbirzkIYTRFxiuJjGtyC2IeCXhZPTHC6/SEasBG5U4PwLMkdcGT3s
pXM9+20/poHcMZGt83OWKqayJHFWVuAHOitjeakiHnL2NG8stWerGlEoSaaFNlfx
DQsTN6qZioioL/+B/J0f4OtLFeMuVN2K9PLrq8GgxozXPCGt9LyMN80a2K8vRRft
mayqdTt63ILzsgQAQcXmGwNmiuP6QkGG2vsGxffHZ8xcTC6ZmyHNe9+UhaNRuplv
TSx4Cte4598OAuirXXujl1CZku63Fb0NReFXf4BiR3CmKeJv+2caLgszbPCNAp+e
8kvkG+aWnidm//TrT2lXRb1wfxUQFfYrRDe9HaJLRPSj7DjTf4zLP4lbQ3Mq0KiY
ZRRFMP7/9u0WuOef8e0XaMqVpaICkGaQCVG1NZMAFu+h/2sCvyi0yyG/hBWlNaxr
JXPSBAKQu93WILiHBJIOjq0GGK81+qeMQ/+OrGCTeky/iUIJ/tMjWcn6uFlAxJ90
X0KK09B7f+eESLzv+DkckDZ9YT3iJ66jJ1YfIBH2h6/pZx3RQ3erDsIlf1paYKN5
kcPCtZ9YGSgBkuGm8x4YyU8i6LhTOhLbxstyJv9Yp5uXBJ1N0i6/J7eqQoitSZfX
7TBI1C8MPdRt8y1+ZDriX2ruhbu9bPmStBv5P94yHKNpdHbSLCoTRJewRZn3fnH/
ZXXnbvbnEBsTGTbQM98CuMkodc2585oRqOyv8Qrd9cynsteQorFoMBgLYFuEu83r
sybk25LSvSjR/8fuUXETIJbvnfqhunQWeESvQCgzOGjzIEGptMoSrsKLst/2qWcw
k5IgZWkep2Z5hCbkc7kfeoJb38g9R3M0UGwlTFws7MDtLB3IZQkwsek1bmK/I24Q
9Se/4QnjrH2bXpJnlHYyrtoTVbd4K7DpokJyS3Xiq0z5pITgw4Fws9GE9tZV5JB9
B51t66QSk+GGyj5maPwZ7KftotOcxXH7pRwynrESXmkzSCkO1Cg74t2NeA+W65Wo
8DpnezyBmpK8KIiumXrKv8z2VKNeIJykaxO2OfsmDHs0arEdUY9Nsl527opSbvhX
6JVjs60liMIwIh+2Adze5me6eudoswCvQopqVPWK84PI2vNdVmd7xIuQcQtjXg49
rv49B3GXmspTO0MyTv2cjt4nmRa4v6MniwFWncCIvbsW9Kg2eEOxHhV46VZNwiwm
LTGjlfCikwubGR979Ujfm6uu8R35tvwLrTMzdBNcvPjqlr4Ca96JAMJTbZT3LUDt
XH3Ye2FXHeSUb01cPB2NK897+WOs/Lv+EaFSUTJrANB2Mc/exbUvJIJxTZP2n44i
v8lZWpsB7vQU12k594AHkEVKuHj7MqJvO6YczzboF+Nnl3koWjOFKG/ASO7TPzoM
sTkK/qOmka57IdWBMQeoDrhnHrDqU/mzGdNhmZvSNSoZvPuDUvPL28Dz6VNBEX5n
o8EyGqiEdmvYxFp1L+Us3D8quAsklqyinay/r/b37xiZjKrK9Bqy1OLX7OyPmPEf
B4Zdd38ka5fpc7muhViBh6HyItLQzqbauuJJrin9smbqTnDm2krUjkI1RdGiPh+N
W/S9VVulpxason6C4pU8BFa9rlCcgp/1YV47IuCXEYliZDKsvVr4UKtWTShBCq3J
308zAaEPexAEsO9e2KENCa/hA0U47W3KKCSqJntQVwAnv+7dW/76BlrjdAbXdL6N
lJjeVnVfFOQHgG4AwDsnkQ1/D2XrVTU7cprmuDQmO3KZkCIDQNh/RyWLeq4usdgQ
Oq3w4ZWd8Zeshs9G8QyZoG7D8KcAVnBtoAszyLgLu4jzf/Mt/9V4A8aOHbZyvTRg
HyrxLACcufig9sTx7mDCw5TZcnaVM41FbBnLLFLmQLShhHOtyqV0BpO7xSwU6aCR
vEUfCfHnffZenS2eJbvSl3DBjfRUNMvgVrL75Tznp1yOLaPy8e37VwAQtwue16gX
CmSzDd7P5jgsrcVUCYC/FgcOODw5+unYOU9X4dCybyGPtYFieVYpVkYgtaBhkI5A
6CUl9peN4VFPiTUzJVKyeIRiTG4jWKaLn5AcuqmllK3wmWNG/XJsTecCHlpfrJs8
8e/Q/2NOAW9Nd0OERmZr+0J6xjj/ApMsvNsWUryu9lh1cAOB3LbsZ4IKel+bsFya
ZZFhLveEUUCdhxYwcrHrzusvzCupP0nmLmSLwz3kPCn/cx4s/e2ajaDnyZfGoDLZ
nsSyxNiWwsLyonL5St5gpsnVeAnPUtN7Q/9EkxJuKaYGKz3LREaCX9NO72l84DdB
tSvdxVdY+pNyK0R+ecIdD6ToCbmtn/ntyETj6FkchW5+tmoQkHPhQ689BmCXlAZL
n8rD+C704pYOvlyg1w6EQxApM1Zxy4pQqoZzb+BmWll1ZHte78akuFjO+rtxpUcJ
HMLr/zO9+pbxBRz9Jt54pSINxJEAXGftLfK/CUGqWtyoEugSinc6Mgl+PXjmHRwM
AgNrd7OmOQYneooChng9q09RQNnsXP5SOx85e/2yOW4P+ZMu3fp0YpXHfFlrS53S
d0b9DKHaJYDujc2osRuv/J13Fj5EDOooOCD19lZ/agaJ7+D999atV832/7KNKKa1
L5BLQQaseprHk809MuH5an7RRWWSFdIN+uAZoHOq9lgXLPv0SblNn5CaNIIERTaY
JNfmklrUXqMOoQg32TS8yD+/+yo27OBuKeRIixmOtjID0sj/r8YK6Mx0OxZc4cqi
i9dKOQIqb4n4YpF1XVBXft3sJnQQK5gHmOJEB21PHFp3cGJkCantTIEYEIB/PWZG
qU5NLAnCs3bVgh49q2zKDegI/wIeDLt1NpMIRsGV61x52rZrn0Ugd++PPZucxjLL
s65ebCtehGc8Wvdu8GsQR1pr9mU5UI8VIr9Hogj3rxLi3g6laKnwmxhZ6Rc0QQ5y
J9f3rhTHUqaMKSIef+it2zTgBVyoAmFyydAVD0N6/xFenxIZBmd2jifZL4i9/vIg
IyZD8LiPugotU6w5SklJMvzIRB51wnYFW6AgPUVOZAZTnwoHEpRs5Sk+0T6Zqrtv
wwa24rLRBZFlgg0o7JWK4fq28nVPa4sN2aUk4cS5ox3IrFojUB7HUIrJY2kvygfV
WA3hVcoMektsxrCGin9vDcRcfn0UEnx7vZ6H970e/yEuSkaffXlP3CsPvif2ZH9R
+AvXcAmZG7mfhLlbQlnzT9i/DuLFhunt8dk76ku2pAIwLVIvUViGszpycr7IpElG
GbWs8mCkZee9k8vKjYgUk4PNBZ83UgrOuXEaYtYF+PBQ0Sum4zwGFkNBcOsPUNp5
5dQNf1uuMFqxRkcMeFLiLcdUj83gfvULTyzy59IsLseZoXr/lkzQenKxBF2zHAmY
aMinoCg4r6yVgPGoe6wpGLV5Le97gqS75bqQssOTTonC0bMewis6bsYs1rrK8mI1
zFmRMmKiNHt64DgCGzQPDlAhe2N8cfhyAp4+u9mgMljxsLFjqytIvOgIuGMJPxRP
+lhdj0bYH65OZO51oNnQsLGKNgSx/7Am08NnFuhT/DPe69Zrv/Fi1ATH+aASXCrn
AA3oicqsy0rdbmVjnBV3Ok0OvthhnjrHzPaRPL4vMYEQ7DumJrKgl4039tin4Ebi
JG38BT/gEsqT2WSgIRBHeejZBiJsg8ZhfmZ1uDfaNqt5hwD/nbzd1YFQO8BdgvJq
KvYqlhbJTNuSjRMzldjcGcaf8UDyIY1gYZHlWrupSYPqqMLb+HbkBsyvLCnMiRwe
pfdGF611lN0N0DuaHVsRuxS59Oq8jAcpO6LRyiYG7bWb3vRaS3hZiBtUzHDuFaQB
gLqVZEP4ul5vnH18S8TqZVfA7fCRm3w/hxsDJjTd5jBNuqxeswbR7OXWkNIgFNtb
QxpklEWQIXEj9xjo7fppjOpmnxq1o6aeo0eDaEQyPwoT3g0lufDl0cTR0pE++i/p
4dHaM5YA8m6OYNXz1HCgppiNvFZOHxXWu34xeSDwzuNKkeyYvbfwRu2z8IqKb9FG
YI9r7pdOgMofwDapRgCyvFaRbBo10atzmU10KcPgaSHUGqKqAMpUVfSw+4tjHcx9
httnQdKq3M7E7k7oTzTkgEnvD0Jrdwd/6KTeiV2R79tNMIzPbccBK63dm71iRFdB
60KTI/SZbZeEsqZPUFaym2p7weE9FVqb7Df/fR+shR9wYzknDNmPyIRIzc3ZuDBE
ufGcZvOCJVcyMpaudZug5uWXY0w4R19A9c5f5FYescag6113Afi/TFNzMY+0kf9U
sQ4Wa+uNtHGLf7UfxkoV1MRQvXiSnaYNJEd8i+zsqCYQPc0/L9N2ERihhftBewpt
s8MvVYef7OjzNlbmMMKdRfhZw7LADap85LCvwRUNDXs0exsOcTiP8yJaK8r+bw02
`protect end_protected