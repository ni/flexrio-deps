`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4320 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
L2bRNdr1lLBT0eERw3vGlH/OslS2312AA6uFwd05okOofOvxgzpfeaHq8GTq/3kT
zsy6FXxCoPfr7yyceoHbslAb5aexxIXcnxMi/riokgQS05CmCDu16ZG0zaeYnRlE
yc9Xy/tn5n6g8M59bUnC5FEowqwmn4d6O66nkE4MXTT7hTb+mZaCypm5IrD3aF+Y
B157Raurc7WpKAyhkbb8jfFvdJW4pczrYwkwNd6pyf2J+Nh2cDXmqasq8A9hYQ+l
cei1nxwq/GvnGtr6Be4iF72g7Zea6SRGWrBQof/mLDqpF4D9T0P6TBkm9TFfNXJN
upqRvzbf11j1/wTr8xiPKruLzSUPpCPQL2h8kvFWPc99/4zW8FZywSvlRpav2nfX
7F5tV1T4ooYi7LMyzTUKisNJ096b9oYx7/b8ZqJvMmjTt7PrwC0/wC9b++ASet+J
rb/kDxVqaIxJqA3iTRyfSG6sOWVmP5faY1Ye2An8u8go/Axk6PPpAbqvLhsstlNH
yvK8M2YxMtYQ/7Y4aEWbGOqfhbqoPBAmUQSCVNVmfhoQ1S8Ict1/Okfo+Vx4bTQx
9+i+mmr+3tK62Kz9q3fKIdLGS3guqt7q2gLYiwCtQwGn5dsIBO+Zr6CO6v8C9oBC
wrdIkQor22mh+nx1974sY+VkVclH4+PeNCY7XFLRWnVcA9fOh0XwmyxGOhu7W9J1
J0vEk4sF4LURdC9VVkJOhWUoVnX2bsou3MXXdI9qmRGgls6UH8xOeH6YLFczZkLg
/M/nzJLB5d1n69agz3IrLqKMDKj91aBUz59sbNN1pwUSieC8VhJ8/UpNCqfYRaq7
ITrGX/FRdAvDMDH6mzcCnSq4nJYhSRGppgYT5yeJC7zNdJf04Icd9oDdVzfl3AUc
wlfnKq47j9qNj7mkSe+zupP4q24Fdn6yMzxfkS4omudNBF+UqrcRjMmM3OayoCD8
0G6oRJZqGx/LsID0XW+gwBRBGQZRPUqrp/0hnhTYMKwaihAfWZgjD0TCHG/GZLzl
pkZ/rzp4FaNBY6qv5Pt5gtwbnfp9npUbS+wuBkmP+3DxRYJtroqY6VdMs0CT+z2S
h8tNk2ZIsjFkctN6VtDr0nGqPu+f8t2Ud+cXhy9D50BdZw50RD+vCSrLXJGIhAVR
cHFUH8WW8PSzOv/5s4QFjFhPDY1+IYHoawrAUTYJFhkcY3bUnJg5A8VqzbxVVKjW
SjJopQL9PhM9x4P81VaeU8CbaEljgWlkjkp+rM94oH/ZGyamx9yK5vsqvqwl90u+
TMtY8tW3aq5qfeDGgA31vdcCc0NwFN+D63TiZn53GGtJ7BKhLYidD+V5orNvrK7M
7WDqEDYo83tdbH7dr+8BQmAHAF101zL3/dFXdsELX+K10dhIXBsWwFPTESRL2SyX
7+EtLY4A2nvigwK3pcX4xMuwy03XQ0a5t3tCgeHIiMkp5lhr2tcGSN65TzlbLa15
C140Oqz0/ciRt1oVTh1SBxRSQ5f3fEQUzlh0rkCQ7Eli5lhZ221OiKcUSwclAUls
UUBYTYUDcMHpH/Ihh2FbISCVaZd87KwbEFHLfJtCvWym8OIw0kdHuHqPmpsd+XGw
TsgPFwBcvMQJl+gwxxsv1sBCHAvGT//bbsmbkhL4fgJU8LS9x1Wfc+ri0mrJ1wt6
WaM7C2S393DGvjWNwwQTSfMm0n95GDH/mcJwCpBXG943x1NRuOKjueP7RuPtboO7
kubbsPVF6nhdqUYau3V1GseB9vnpGy+IwELSluhHd9coHNkiGDmahrb/4+d7OM28
oaO9rXQN/txOuO0F+FrBCQRcLuZG8mvPEKCYJscEMLIxzqEodAAFIOPlPvm7ZmfE
LvBxid7EV4z87SseIuVYH1mp40ntkseeV7ZcA1Ys9objtAue5yKd4mR/NR6ab6XE
aJdcv6udnNzjfyDNxKCNrmSYq+/gaSFdX/PZ76/yVruKMhzOQ1uyht/hcqNOI7i4
kGI3HAC8aUBLBAyssiRMKImvVzHxbaSluBLTN3WAZSjQp9SatwFi94jU4+ikC+H+
16Kj2uNg8KHCS01/2do030bJethQPFNJ2h6+9ifcZW2CLMpuNydnhTBh6K3SgpOl
H6+dBit/+JC/QLPwMSHT3ednUeXr/6slGP04M5ZTN5oE78ks1L66pyq/7KWfyjaY
NPUQuTXNSH905WCIJZvTlPoUP5l3Ce66bb0lVU2grUoW9xrT17wpVWFGYxXrlNQ5
xjzlKUmH9KfD2arV1jmR84EJJ6FqK2iyHCqs49NyJWsipnEd2fpbzGlf3UjOpVrJ
jadZKaRD7ZcEGJl2iWaTNj05Ds2OF8+w3AElZN58kEY5r4HkAcg45gQqax/Bvlej
HWrVPfjN99Y2H4k1I7/C3uFjNqQfH/9phMUH1MUAS4WlS+khJtfl8yurJ7WhYeNY
bulkIRVhVHe/dCnn6EnIyGfC7TpHPHqEeOg5sE1QL3owV8Caq1UdYR6Cv4V/Cwxw
/lVgOGkHcz3fz5OtKeMITnNGfvTo7qhroHsD5op+B/mRZ/+bFmvmAKJ5TuAejtr6
eivwvupbHM/MZm65Iac2uzzmhlze0Dfb0R0qzZR5m7s2Caz4KpMLfa9W7WbXXh5e
hTA3m68daV6cTLGG6MNCmKk+/SfwTE1ZNV/Jc08Q9/lxnRELjf1uKLowbRPyaZxR
cNT94z2d3ZEnZmCR5XAx3+PiIYwbzdWcecmrKj56E6A+76tOFIH9t3CfF1OXMUhy
a4WD3TIeBPE+aHdo6wNOzizxPoq4KiCTpIYdMMQBEFD+XSHAfC+ipeeCPWv/1S9p
HTIP7Gx1xI6dn+acGug/TrX8fQqa+N0Vhs9fK80lECU9JbFPeo8pRSBcBY9KRVSF
qpy5+3mluR9AsQVRvI4VYR8j5jIufKCXvn4ExMrdkIptqMSZOMVB06e5p2eDmIRL
8SrYkYSsp99vxmjFeZG0BpFOUoAinNWkeC9N3grr9nas0vNqJcQBKQ/yFiBX6rE/
TslvfAQhuhiAnuvLJ20dAhbJ/jv/sGVKZX5mLrCCBf2k90RfCSbsxvJc+YfTCl9j
xd/K0qyHbNr30RqqdU4bIyUVVEhdR6QrDLbyttNmCI/m9jyOEN2JL4BYp9B0TqNn
Fft5xf2PGbpOIOswDv4CztGhtL+g4eDDwrAadYZeyeZU3dI+Op3QBLXSVyUXjTWo
PUS9fH2ioUwM1593oZliJAiTjEO6G6cGG4zb4ikLNbZwV5LpA0guM4UdZ1ecktxb
mIke9j2VF0huRuolpFl7zUsKN6H3mXDuP1bQlmAD8KV7GbfVxHEvwd/sjFAGekh8
oZhD/OcBIHYgA4+oovGT33DDi9OeVfpeIXX7d8VswYGZnbDVgm5Gy/TOGST4mCMG
+/vZhSmXxP9o8medo/oL7w7PX/bcb3tWlvye/uzVvGW5XNDsXcEA0JOYPCFwjxp9
YfoV5DQ8hI2lqSOJwdReUCadEE8NCEDVVsoAGxuHfV4PLEjd0NXllXq9E5qjwoAa
AEC6LPUR0aD1i2wqPlUsrbhJqtAGq424GzkRFLtLas3BRN9x/TGkY3LKQyGh3TgM
RYv38lFBDu/VqwFyxU9hCX6qkZ0kiMdVNbS6PTfNs8fJ80uwx8j79KZN8rrfg/dn
LMCIZV51BzvLTMMhzNIrDNtu/O6SBqEM7VMrK7GBBFZD/x9trLVsREjNxlK9nTuC
9oHqUcDAhlrEJanXbTsfJVL3LHz8DDMlxriwbOhSweb8X8o8zXO6Iz4RGQluIVfs
CM6cxv/EQq0J9nlWVFk5WwiG9fQk3k+TafZ/KPqr72AN7c1VBu/EYBM+oDb6+GlF
s4g9Ul46F+XLOpFjxjfAHfcUTeWdyGk89vQiqkh8Y+b095OGNeTHZiWxRPEwpyZo
fbDmg87C7j93RC8qQR3KfPiQeaEnbAYWgo0C7c0zY/xcoq606sn5MMstSsHEMjdx
YQTEmf1GkCLwlT1+MXC/XfgqAawY49VkOFA1gj/uoTw06bxRzeL/H+pXxILU95g4
lRI4vkZJpiE8lstcgU4QjIwNlHDnNcRqrD5dqxNikhwDXlDGBTmA+nZb+No2gyv2
0pLIDNuebZljXM5MJJhCt2VdKetGMiNK6wiDSyjDSXqANQGjszc0gNbslbBb0/6A
jZqioJKYaeRkF+C4CFQAVQpCBPfbeKsB/17lSVNHxoqvEqaYLjqlQk50F+18aPxd
BkgLtF10eX/wJr6oy1Wtk7yESfDdadDDeDubWmAP2YntqaoxtZe8vXHukHGixDji
lfd+O2Xhsm7eN/zBbVeYIiT8s7+5lW+7hMbQT5EuEte+j0XA6gCzkw5zhKQgcRHf
e+SYUdK7wM0WMiDZQ5uJgqOUgFkx/ixAWXGGW27XWH+z8lZjxKynrBCG1cTqxdkb
Hpvcq6VKbZAIBCzj8Psfjz+ygolBysNwpVIJBXE6g1/rE/hRu/Ka0/Og5TFok/Q0
UvPprc6thwcvX7rhmwZeXcvoAuoxIBHlM9xm1yST2cBqSfkogyDZ6n8MyW/4teCv
CbIIKzEGpYAIaOuTar9bKeqk3xn1HhZzE8c4BZSWL8ekbwtBdbdDkDqT2/wyAcbx
jIK/BSQw+B/xqnuRuqcq2tOb5lfoQnyKt+ReuBg5oojd+MAUQ+l9YGQugvLyj3CW
bR85x8lilix6BLjd/EMIQlivypr+GPvX1O1xdQE5l53O3N6uT1vySTBzXYECrvv9
Iz79IH+bCSGvNam+4cy7whi2Kfzbn3fKpDyA2lNqYGbN2mNwheXc3lYwW50sQTfB
JRDVwVY8QRRugRID09aesyw0NP6CegnKYNI724U8UwUKbS1n74mvvOKC5hcM3NGf
Rx1Zb35wJnbOjwE7cSBZ08ITCkvgQjqqHDST6F/hHceSuKCuGFstYNNQ/uuvacgs
1n1XPCuhVMagCuooT1JkbWw5kmdW2rh4gdfgwdLL70gbyyRxYr2YOY87cD1usgbj
WsJXApyO0drsInD9SwOF5zeXz2cRQGPSZLdhaKFQSjRgTb5RPUjRNKgjXBuocUkj
Z1VksJXnSRYB0PrsCnOpM3AHCePO7XY1BHfaw9cO3aFOYFn0kyld54V1um+ipMYU
UpzNGFq5/z0C3hzOkpTqUTMX8R1TZjfijH6wnHIoSDihiiJ3RDyF+x02NrXhgM7p
ybJhd8UQ9n4LRXYadGCc1eVCAOupazPHZwNpcujilG0XlTR4/1w2hhTyLAvgCdIk
oomI7spSFx/I/+YjOZLFgaR+989PJaVCytwyaTQDMdCqDBq0FQMhqHhJVS2JnMQb
Rg5DzPi+JSvvb00+fD9VlCf0j0vFw8FjatIyQObEwsB8iCiSODZGMX7q5+0OD26H
3T4DqXSX2Vp7zdOnFncGNZSvwdmmi1VYlLWYZgJJFdAiARF7HCuXjHO4NZaWZ0ii
QQr2xO4930QImY1aoWYmSqOqYNMIvvincQOGY3Ks0oDFHc9aGbJGRzdYcZfo0OTE
zmKTeacASCKP2Id3wRJlDbeiOdGhkfj+D94wXMyOeJJ028cD4nveey36KKKC7oAy
WUBIgWyT5HHx9ANCC5lqtqGevRibqlPq+5Kv1B6BUm6LLuBLIj2kUj/FMAWK8uK7
`protect end_protected