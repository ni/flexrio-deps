`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11040 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIbmtDsHrDP4hDy/xrzKHF190yQcy43hTtXCBsCYQohkUN
ubueGbxLkxiMi9s5/yxF0SwSh/5+DCYAGPYEUF1sY1yTWkyzB73uDoPjYsnTzPuS
146sX080+/QkbSw8EDwMkVFEP4vMbHZTYydt6U73/+dvQMawxzM2/gmguJg0pQmw
qVnG5LggLK/vGF1RntqQoXeODLsosAH0SGHTkVnFodDETAzAbeJmCa/agSRAa5if
XGJnfb1jTmnzhUYj5HXJl2EvfWMiF4v3lReKe9qdnSk/KMs1aeeDvn8UEh4juumV
cEAil9DuFw+VGh8P8Ra0qdqmuLVtJ3KNThf+9s7lHbYDbweh5E/IHYNaZaSlUwoR
dLrZ3I1kA+Czu6iwExfagevJcMAiUag0KaaBPVoT/I8GYYF95dNrCo7uJKOSNcAQ
xqA7Pia6u8c3xPtNzYyLB8G8lEIToT6TJrX4rvAVtbaT2dQqbyrPV9bXHTYk7R70
dKvKn0hsqbQisMIlK3OITHkPYI8P1TYZAHpF97phvWsT4gd1TLP0sGLFx65vdt8x
3UIZxGQvOFizChKuRqg63j2qrxXDJH1x9WhIGyq3rdQizOw/DSOKVkBVdlAMOYw7
nmHuuxjHDD9tDBvx/P0NcBfOnw07C/OnxdMyXpvwYMHgGLOOmRvChFVnY2pSSK9C
AtvQxKyjOhUa8NAOYAAYf9p2kotGQpJBSKyQkvM+rQOi4tfyqm7Mfzp8B4PJqtmU
HUqyWfTzpGAyDaR4wH+BPP+kusm18tEsR/mP+sfT9wwO5tqSJ7JOWth5FMtgA2Ns
knV3Yupt0vOqf5/yMjm1KGKQ2ukRkKpZu9Gr7N9IxzV3Si69fCqRIbiAFKnWYDZ4
iQDcfVKEvYoGvzMZ4NMG2m7IvBQcmfNm9n7MUqyIIACSVXhPUHtMf0I6mKlLoX3P
doptcRICsboi1Gd7a1jpQJoRkIomHE1er1RhEPdNqlQ94730onon1Do0sTADh6PL
r9urb1vgIooWfNiRlntv7w3WTk3ffRD43cpO8C0E/XkgIMVTnq/UuwKQslBmgjV5
wJfmFGtedHwlHzWGpEf4Ls1FbQmT/yz6Uuqq657SC7p5WTkLV5QF9b9uBynqHeUf
o5TjL2W5duA2yaTtIIwAxl2NPgvlDkNO3mG4FzXEZBPjG+Moe0J4H8tC3C/MxFSx
+mpnozQix49Rg6GfzFJ+RA796jq7ZsBYONUHP/kQCCoTOV+FA3wCPGzjE+enE+AR
yGSU3ka+njU6OHUD3JrjvKvNc3y5SXxdrhBP5eVID5ozO4VRkARISg1Z4aEBB8kw
z0CX6bfSIpY+Q2VDMyqAURc7BgZvuy6Q7kXSb/rC8Zfx/Gwb1F9pauZ+GGxho6pQ
Ajb+Oade3khTcT5/cgPLDz/GLGlamj3SRAJptHDr6rCtuTO2YWQ2o0QE8geItzug
7J9N1myGwWhH9/cv/+tKDY3oo+mtBZkfus3SOYZzDaHQjP8SgxCqh49qhHuQgSLt
JXCQFNZdVayCzyQqcsaKRjFtHIbO5QT9+M340n9s0Jv0L9vHTqz7n9mYCCjVkyVG
VKGe6kVT3Kh+h2x95f+NV4mAkTsRGojayJcsNKlaTwZZkWA03aIDFgp/KkK9HjLf
Fnr0S5gYivJRFL30zcsJCO4+/rVNdHDYel0qhbsSFVVeVUZnhqNVXtM4/KxgpzBF
oebNOs8KYk95WC9nAwvkiwEFhXnXA3FtxlM8CoeLfxSbpLx76tsTGNS64wzPfr1K
YeSKHJDTgTxlF5v0GqXeLe8AQAZvVVVsYwI5QOUbd8HPWmB7ezfQTn2XPlIt0foI
Jybmponj43U35hQCq9168PHPHTTNdiHP7a8zljUZzIPTdwfIZEbwUoXKYBZsnC0K
KeyK9y8MQUAetnBNDGwL7uHHVIbMqdYwCAd3wZgHPdkiW3YIJAgIKivBn6ZWKinj
a68neItnmC/hwrwwXvcSA7vaGvBYSYvsdO3pB3tOva3ICSF1bAvpXtZJqvsa/cUU
vxHUj6holCpBtvKaHq07Q9+ulKcoEDEhGHOSbjz6d1UhFii6nofnFlZOlfCpDP0E
7lbILhtm8lJsDraF/xCEpO/zvIcx04qhOHOllTwbJxTWQavVZpPWK3pU/h7vnqMX
TsV8VqXLtO0bNrTgxjl2uGiRTtXaxLnW6OQchAQyXo/P+vEmWFI8NA29MOIXsIq3
8Z0DSYDBJiXCkqS+zkPcD637Xu12eH5xDip8HBgjvPUElAI4xOzowSLb74Qa3HyH
P5vHTIcBNUoabZEWAD2OUU2HAf3FaMMVz6Oyf8NvJN3LEPEPlBWKVu52Veeky+tB
Lb7uOLAT8QWrm0zGlV5+0dtfkBrT7P31Ne7NImpjMl6ypH6KL+S66dJpwDulxlNM
CRBZ5wvxUX0uJJjhfdSeghT7DcgRClX0w+rXGpi4zMaoH0/EooC/oRmeNxF15Dp/
dJHaeCKoCVivPwq2V1humicpnusDBJW4BeoU+zKtdq+OCluBkuyICAfBYOB16jKO
EfkXx2HewnoB1mGzNC4rpa1/ShtG+g8rcz9MRP4V0zbyl4EriZtAqaL3hPgwn3gj
RXb//oMXxM3pCzL0yjwh9c/yAT2nyaMIk7gQs+vZFaGFPEp+9kGmCIPVMD3oo3Co
2Fd7x6/raD45z+rid/FVtJL7pNYa82JxEDaqU9MVW2bfFwQ3XKOTE8qKNH26H2i4
iQGjW0CAkxt+Gky5jB6C7d5HjzqY+abpqoNN3zffJ2IQ1KUY/LVa14i48pU2U8KL
aMoEgLjRkwsA81qk1+h1OFWIP6K+JLVumt5JI0hwRwOxL9xBQqkyfUOzGKqlFutm
Uf/GRMfOjY4z36aMKpf6fbK/YOPpGFwWvbGzTLh6dNQavaOvktgkKnl53szwXS4F
0VISMNVuXZOxIjUVJm7QrkHV3OzlH0G7PF3fG+1xL8Ox93uZ+fQCOYYOgI0rbJQp
/ACGNgPTRuRC755ayuc1HygZKtpHMCvcg9mD4jDO6KR5GmzdqL7xLS3k6PuBVxWN
Cgya7PU9Sy4Qj96MIcmbvtCXv+61D9TvYNfsHbJdv1E6FlomXZD4THBQpoCVlrTL
ITh2vcf8Q7lB7uBeG6uVVrgsgry6RvI+dCb/4HmlO/Z6Z1cKGyy4/pzprPjw1mjc
4sEgdOEhzJ6nbL3uMZ0HYoNNJwwFCRFyEBRH7iYo5vBcP4qI6PDMhiUduw+u7uuC
cP4azDVtUCTuMTbGYW6jr2kBgT9YWw/IQ9vGWbAB7u/My8Btmuns6bsoptAc+7kU
QTWKveCFwjFcGMtZ22Qhy7+8pbHVZeHRhA6RgR/tuXUadIpQ9myS1G80lJIU0gQW
AVvmAy2yiCADKyDBedxm14CLpAllNKYtxyDXNnXpqyqeJ2Jxf85RyNpP/jJB0Sl7
weJHq4DLOWN7+MsAbut6W7QOQJ4Mf3/lntK8UJDFNGtlyw5sSfyaVI9G8alOQ9Sb
t2fsG/tg6euNejhxMXPa6wEe5sKcrV5ype7Tvl4Q2vfKwx7pQzCE15L6hpplOAGK
yDKrFe8k4W95uMXE5/Tsnuzkd1vVVpnyhcM9w5Xk877prKg4WZDJFOsFvE53gp2V
sCker11He4S8WSU00ByK+tM2cNeaWDRE4DcUcZyn6jNLVo827W9slYmHLsSVMGFw
x1PtoywFa9DVF5BYquNGeBntdGe8xZD/tMfwxfEgIIL3eziKa6QviNyfZ4Xg/y9J
u00UPx3Umrgi12w1rWHiwfaGNq8cnhRchFzlS2oZojBSEeSkEcVv1/kMSSk8uyq1
2Fom2Ax1bENA7dtqrFN4Gq87RJMzayRej9wY1dj/SjFTYzmLI6Je4Hx63qSyPSRL
1tuvdj029aqKVbcusEgOUrE8dLZADWM++zvJ8Ta/qam10/xFTuPNjs5FGuNAP5Lc
O/uje6UWErahct9C/brebIHnHxiMp5y/DEFv2nIZOjI3km+ephjP/BiKROj+SIk9
Onf4up6+6SXx667u3qnL9YtnjA/NCDH78w0dZf4Vp4kYGB8KIzPStEix7vAXsbU4
qc3woR/f+s+BT83V4zn5WVVHdYFq24ZKMAOTQe9XegRAvrOzlIdnX24uPpY3DYeX
bwfHoMsnehjFYdNg2Vn4Qh9h5dy7Jw3HbW61mlp2+9yapgqm9DWwdKViZOPQ4olM
jpycj+OqUC+DbRnpW+hVr+RPLGvi1KKlWmnxscdY85G4V18F3gsrCaBFGAmTFpSc
B3aiw0vynuIOQS2gZeVi3dahC1V1XJqlA9GPAIUcY7ATO8hHb2PAfl2E5YYfcVDH
vLp8f9kTNtL/FNZQfYJ2IHqso/dzk8DkJk+7pxc0E54EFDIAolyYEAGke1GcGRpP
wv+2JJNSaobi29seB4cP87jD1AqN93SUdUucqk2qYGaiqW0InVBHk/CwLH84niJc
aU4p0T5HN3hGGsm8yBnnACJfSw9iv8ovQqEoG0aaFAqgyvU2m8PNklBnJ2FOefVW
GWKtpD6FoGRKz2WUBzCPQWtDtsotvSiRM+BjKZGsG45d/167uD7YCFcY/Xv4HCJT
TSSEna33tUaUo4cwh8QdVqjUBaHK8gW/WhLxmgMFQHUK/Rqb/D583MGCakR5mF1T
E8+XY+2utUAEl55rTTjXjfJKVue1DkvCmyt2YihYKKwHic1D68Huykeu2pLoVzfH
/K5vunhSxE25n34LXS9tog+sSdZrLpXas0d+BJyaj3ztca7bt28Dds+R8SQhbbWU
j0Auu0nMHJkVn9LH8YB6pVM38LTuYb/z8zHpHg8Gn6YplkuR13P3cWq9O3E9qS4U
PtT17eShE99HGPQP90RztP9sQbMS2kyt/U3kfdwEFA6eiraXneWxV43dlfXI5AS/
WvvnWSZPhq7ts9CjnpxGmcE4IcRFFHr0zZ1/y07ijGNoIMhU5pQzUS2/KmzORE9T
xNPuXsXadDB9FW+fmMh3/6gJETKzHqXKmuSFj+hk0OtQr8ArsIFXck5+v4ix1d8/
zpyA87gNARtYIEk1NXVpm5xGBqGH3WwlMFSb90rWw0E+PHpY0gSTfQ9ah+U7WozK
NLeh8VpG5yp0SgNieBrU3sox6hd/U36KXEppe8TlzjcR9m/QzrfOR8ZSGGEqo/R3
U0oPDOptCj1mG0C8Jb2wahwqmz0/2J2yRR0pxRv/9kM3p0qfzF/f60JZDf4DVEyd
wi7JNM5R6n3X9xULef5EEcMDB++AWWGhEtc1aV26Zty+oEdcvfNg6icVCKOOKpLW
9MJUtI0NzH+ucv0Hjj75lNhJzELDRVge7bVsyaoq4k09mwKA+oo7iJpJjAuwxZ8o
4U0kTHIGppksLdS1P3Ow7V1YalTS0ezRtEvRytP0WzSKAZbgxW9sAIVW0SlVvPTK
jJC6l0JGiG3wX7213mrmq2B8ZZ5SXZ0mxpkWY1id+XxmliIQwmtJ4Yz9eGsjtzvK
s2lYyG/R2HX5SktIu09+MqSq2Bcw6ytBz2VcKovAXFbvupVBz72TLQyazGRVMFUK
G3GVbSu6xIqE6ox64AtY0DqUjlgO1a6rIdo0LCFwygi2qWcN6kqBfgXKObdzfvkk
gYRtX1nIvwsQc58E1l3r9dWpinDwu6Q429tYRPuE71GUN2gPXf3/V8pX8llNbgiO
0bRSz/yjSOtXqDLcv3utX+N0kXyPXjafX3CY3KgXOaB3Ecy4LaDJyp1JP815r8cF
XvsHeyW0MSVNs1DrlEcNGWE+kURJfw8No7O/siWDjjkuo4C1fB8hyi7jDAxjtTzV
QASwgWU2jW88rhUZDFkLD3Rl2h+jD4eJYS39+lSK8nNe2Y7Crsl04TZL1FbZPmZl
QHIcMyBLU0KyDEelXZXVAFjewRCfybEwxwtGq5+QrDvMKRluVtVWCI7klt5C8qGY
oIgPt2bUQJcH6wodT3192dSaL60dVgyrLUQDwQp/bs6U1dB/EUm4GYl8YN6Z77DI
0O/zJCGV7HRQF3nt9PTR+7fXG6N6S3UOEgvfgMJblJj7syh9NfIXPzF2ZpU4m7lB
kZUHczZgwaJL2C2huSOBhlYIh4fsVf0jyVStp9l9m2h8It5+rgc/Ibb1to/UhuCU
nKJh5O1XKQDzG8hDqhMz05PbFMG5j0bK0pDoB8v7Lv80wf8DyKw80IdlZaaDw3HS
h7a7AVwtfzrFmJUspsICaKMd2YXSxa6zEpq+iGIFkY7Lyz4cF2KYl1skbua2nFsY
uqce1jhzDi/UYOW6uwwe5iBqG2b+KZ8IfhY7OdkFsPUBGl/WcKTGHV9hrTEdORaZ
3CkZSHtuDWckEdgjYJBP+OFASpQnm4ze6xsy9BrIhlnl2FfIbb0b5rY9sm8Bw5Yn
/8A6GRUpxY0cN4z/f0onIM3SauUH4o8FzMESEB8TM9FyQeMBOlIc/bOHv1R8Zty9
248D5kBOCfSwQxoKo34b9TZK0CPL0MgHQPL3qfJnuicFthY2bshMmhXmm/q60Lhh
U20H9mePeiu5iN8kck7UxobqZMwn3tlhmVPUBfqh/J/VZNhYNFGzprMcShHF13UG
lcbbYsQFZ0OSyZ6Ilypwzdju8S+lfUP1bE23oZp2gPv90OsOfbFuI85tez3+ZTdV
J3kJNmj3wf07YU3bZTxDZZN5irpYjXA02d/3EPNGn6FTJzPRxBPo4688iFcximKf
n+MELJj2roSi0tJh3gThzHTMRDk6tFsdiXjbXL8tlVVb/+qm7e918HdY8x+hlWyl
8JDzK4yuONh2qjma0YAKpnY8Cevxw0DZN6E1ul0yOifFAe2wjIdeC+uJwvRiVe2H
WYE773kvoQZPQInQRuJM6aWomzCXa3d/9itW4YrHswbOvFzYDqYrC2yJkMIzviYg
lFoWi68FYk5Mj9BF004q8JoRfrehnk2Nmlq/C9of1oDzKD20vK7WTzPa6sHbNtiq
aTDc6FNwVPTEsjTEStA+GYpntGiwYgtzq0vvD93YtX2AOVwhwgZT4q6uWwa/9SsA
2VSebgzqgCn4cnQ0t3Z+wo9XftTU8Ww8PitPfidxfmYkS9HTVP6ElBVox8IWPsBQ
OkYsfr1+YGVT+/6O5pgAvdKKjomd5nzaDqcLycJXXDqK+X3ppJqp1UdgKnX4rb5K
n+OgGIdrXcd6X9CPthPyCzs83ESOaT2rfyd/1jqbVCxEHf3vinxQAtZK9Oi9KnyZ
LxKxrsJza/IpFR3QuPB64D9t+qNMfEXa5/bsot/tcffAXJFbYwo3Hr4Vd1dqtqNw
MWsDylEL8PPEZyRcMqvgfYsisJ84v4Zk1JZhqXQJiz6FK9GkI3ZjeRYBf/Oe5hlq
hxIEi7dzwvXKtJg072BW1ytV9jK4fe4u8sgmO2sLl1oJPls03trdxjjW6DnwCnXt
KZHuROlRbpw3kIujgOfhOWTAzxMsFUTjYdAwlo8qEEHKf5oWNOMfzDbcS9ZhJugQ
ZcPE9RsuVI0P4kj7r6LtFOCrnfbhcqpb7npy51FWdFANXddl9w1HeWeEcr7OBzEt
LF+zlivrpPg7X1gIiGef++u9b7lsh8L32x51Uis8/tXwU7jrRwMSt3emGKEnPvei
MJWFD4dcfAXDtEuyGyEXZCml9NcCdOxyyZ5AVIIsy0Oc/f4dipptcxVlP6x+dtc+
FDoAq+a2kKIR53AngQvzgbpOwHpUWH8w9HbNSwfCqJurykM80oh94ZM75MfnbGJb
cJClViH7sEmW5y30kt3kvzxyQATUNhn/hJYqfn93GmUa/6wwjQx36kLvXV3Yj3md
yl1+gfgnwubFJvxBwINYzyFls6i+7iC9XuXFxY39YYsUPEOrOChXasi08o+jEsbU
Ci6QNvbFgaBJUlMf/NwfWiVdMbo2RmZUGiTfO1pbUmyTXDnI2+hk2ik9CCQp0g/M
8q+51iAONCCKc0mNY05KgaTmEH2SaL0OF4EQt9nLbjr/PHipDOdH7zk8qdWjk8Aj
6NCZ6Z48jG5nJWUAzIuiFuc6UcHsYGHnVVz+H8Zbrph+DXqJj6jEXHsTVQ+XTA5x
DxvLnbcNbb3/5aDibMR70fja76rCRU/U6RRQE+O1WUr0x1HOC+5xkuuVHSsLDh3r
RKczGfia+ZkOW4EOiC6YJuif1gSaWWbeiMzv/SxSn+4U8MTcpqpyczgC9j7wL7Hm
Hk1G/ZR4fZc3k7B4ZgrfOXYp1ee2IKSERJon1p+Udm2YySTA9gKZoY0rk8byf902
Ek21GPDthTAYfWT6v3b0g9JoRg9C9zSI+AWhGfKb9cmB7KAPjC6mdq5otrt9Bs0I
UGa35KdDIpN+qpO1Ezj3prQK3GyIaPylG96VjAPtv9OpMTAgLJx2EFEZKgOnYXVB
m3fJBtTLa69isjevO8jNLkZsH3Jn0mBQ3aFglR5v7jJRrqITKjnuVD6If2rFP67D
paNS8iHbL0SJ51MC+TUFniOgfn+Gskq0LZvXLdiy+LY9+Om1rkY7F01S3V8ZXFv0
vxc79bHlv/HVmVwrZmtOVLicjiZqC2vOMt5asBbu+wVfYcrsHnYuy3ZCqUMhIE9g
f9lIKYGp6M6tEJzwFrEkHqCtpdkK7xBQcdqeShME2R73hNb/ekQCCWcmIDGJEViN
PTy8S7x0E1xnb0cD1wQfhKlGYb13o4GDzIl0smjgK1aPniMo0LZ5GLFJVJxrOKQS
Hzf2hH63R0+fekBgxBPMUBVFE7SWVUFOobZSbdD3MmpYLY4MEP3Lb6BtHbEKXuxi
I1lSeFeSpqXdd+8G/d8l0OrWPAcDRfoTMTyhZe7L3mLgYjQZ6kWEPO8O3mXxi95R
/CzsO/EuJW9kvp8Vyjq44qxk2FPZ7ZXGiknorFxxY4l9O1cylnIXxdmCrRlOUEu1
1rrxg1zDhRtOIFOyKk1xJ8iSySpqtVc9WrCMulwB5Yr/YDERgPbTupzmUgPssEcz
ZJd2fKKOZ2N5/4XrN8D7MQdh0di3XK5Gm2Q8ZT5Za2b2xCTv6KKYDeULxR03LbS4
NcL0FTusTBGCZbTtapOm9c/ff6UC+/4G7kTsUAOxv/MkBHCVhrAifj+j7V2ur4eQ
ErqtMDiFlqhbGmOT2ul0aTyz8DPvtjTMPtWkTW6j71j+SPDeRB/ejUYtsF3pG35F
zxUPhurLNiplBEmdu8EMwNEo4qVffrTIGhU5MsZvoLYWgWMyNtEFZZgozXaP5cpa
2NVQeB72pPbtPn27fbMLrIAYqgRIOPGEnusEr5FZlMYRmM4RkuKGX/ai5/cMAUw6
tOJYNJ2gGTka63V5vvyHYYPGelgz26D4agrDp1m/EDni898FuAWEDCK8nESt+FDU
QjSDSNj4TwSIqx1q4Irr5HcVblNy3q10+4CLdDmbbQ008vZW01VadWeedWrSFaU+
JK7B9K8rdks1PD7eJw26oH9I8f9SVDAGo1MT0+nbpmmjT6QUd0EXWCygDeS9Uffh
tTGPSb6saOL67PomH69wf7xDUMJa9Se3IGkDysevfTYArMZmW+sS+9r9bxhjtYv2
yFXYtnYsZa35uvyzpTeFpad/kmIoWO0yoDT1vfj2LEBF744KfGaF0QOOeZXHrB6S
GQf3M95NnqnVcvIeBWllWjLSJKNDXRCZeDN0vTXsN9zzdG/heyjW8vlfkfgMzuiB
bOScq69w7S5pCVmOgo5tAa0iLwoWA0OU6xy2mer6ZLHgrvxlaXy1jd1Dbr/r4WSK
4gnBeT4+Y+65kx7OszSFrK9Yg4gwAu/RK+/pV4yodAPlJoQSNuUqFQcwQGfb8Jwr
PTYO5Cm0PupdXCP7KLkeExldnsALQx8uLxMmUMDj5/EQkN39f+xrUyjAqLvLiA5/
rEBcGFhp3UqcEf/VsMp3PpPtYoNwEaEAwSApxRhO7qrjdNW3aFZjbAWJFpgWMaiV
8h4u7PlqQbav+0PLkVJIhJWcbayuDI1QqIRQanrIachmt7kgeuXLQE+OAPKGC22B
qSiCJVP7x4kpHlv1Yh4+TWL1bQHbfxL2IG55DKmT1FU7Mzi4gFzbM3Sh74DoNymy
g6Oxg97TrLVWQvZS4DAdDwM7OHnr86R3RjBB2OR9efG2okwcEvkTJJ339t/RSg+e
HGv1l8sSVobNBAKCBQg8GFf0hKJlR26F6TY/oG/OBXz/pwKsCFudVQEWdLOkY4EZ
Icx1gJlXdHT/CqFOpbRHDKekhHB598zihDU2jxdZOBcbFhLQRfnwxZOYrrZVuQGP
b/PUM62JmRwPpymeuDM87LlAT1kxTdxb25SLbAxl9DNKZa06sze9CjD0874GeboZ
E9e8tunqo3ZpG9Ow6MTDNx77c44HH6d/hwbOFJuuKepDhBLlOIvRbw71OL9RTktb
7knYNT61f4gbzvQf2F7ZUuKiakLd9lxqYe1n96wbeSFgYbPcNfrT7JfYlqslqAWO
F7EtmXyaaD2MI4pqlZqA94liFACtfvBE2iUQ/A+Sw5T/w37BOM9tR4ArrJswsRKH
VTWSBollxN2ohZRkmZAeMKYKeGi+7L0FtNHcNH6KCTyF8aXQA5ALjxXtmKj+LE3T
3+FIA0NVdVJaHo2BLjRQONFrbIuDa/AL+U439gj+X2vgbRQ67K6plhN5fYZqDvW5
0TrfMwRkjhDqh6B5OJoMSp4DkQoQM8Sky3vghbYl1H3BPkyL8eGTJHBpJmpDQa0f
2kUhTapzzAA+AU5Rywjo0l6SkRM5Rqm9mrgcl8RZJ6tP4Rv8pjvGziZTyg7G5AVl
+MmuAKI6vhxhIiSEeQjBK344qdhVdDIK2zEx+TWMqexfm+0j22zZHcMOygRJ60tN
7S9Y6hsZdVK+TKmqua+CoDX1bRWVZTXaiJfxd1J+MSVYi273FFxrW+nn53SHHD7/
puqHaw9fyNIisq+4pT8tN4y7Qs30Kv6UMSFkORyYY7ffFDBQPsklTIhIfWeojSWp
8EleALvEbLO5r2YQws7ygpm3rlsnkzz9hZITqyTqOGfvW5nkD+ZrPBKOtydAOSOE
bx/9I6HQ7Kd6MOUY7SLFWEfHmK+ZWchofWQe7huncU4EfHaNr/m8c5RQr3zjMYsE
1MbB/J2t8QCWBoYoVHlJxfO7Zw1E0KjfrtVD/rtWcXqHpgniE4uXH9rvNFf231+h
b+cCqmmOWqtKCsIP5RbGiis8kCJFW6rCRnFYj1p5w/2JA6BJZ3/Xtm4+D6arhmK/
Pjr2ou/BjZ+PoR+hOGLkeVpd8u29x7rHO6p0L2gwEs2PPlOAPNNx8TXjTrLmjA2J
0+aeLSiNweFOor7ryeFJZMiUGRmDVFPoid915LpemQrErrPbvF1wGIke2yEaQOSj
EzIw/Mu0R3eKyVh3fRbWAWXBm/FiBPCC7mjnVtkL0MrtR2CxTBcN7gQ54RTI3mc/
CDeF6hsFNsQR3l5VQ5Hj2DyjF1n2b471QpcCIn6diPQ4ZsxbkSABYVPLZkwFA2Us
Jt2iOT2LfUBtUlA7HB7joFh54xIqZdGx6EiHicLAasJ45j+EfhpZdDS0uARWUH4z
AA8oQVRrFJc3cez/wz5lq+P4zCU956r2RmBhgL6XYzyonHjHGGYrAh8FiDqNfs8S
9pv9DpgFqCcIRrbjl/VEAM5+Lbz12tteG4bBkmFP5nJzMjdn5r7tapEYTk+N/xTZ
4TGj7mVNUjAckiDT0GK5pduPj2ih6bzqufPmdGK9d6Hy/KpbqLFWVARSH8D38ZSV
VG/OL5Dyupg8/6mp04dkrWkEoXcT+KliIxaxFe4k2x/hbdXv5ey4bNwajIT5CY01
8AqyQHpT1A77FPS3JcMBZQTXRHG1YCMOtXrc7pb2zecJfGwe7zdb0RGqL8uViDVN
mmtQZAjZgCyNCEL+EFSEKE3uYrsJYQjbBakUmQP6HtFM9ymiIMQLzOYX1Q7+3IyV
3NeAmClAm+mji9sRGDe1Bl2wU884OT0GU2DbyxWOtnHORul4Ox0QlP1Reg21/cRC
9iHR8/oexYXVrT/70EONIPQQ7pd689nn2WynoJhosR9rHmVDjfSkZDRCYq78saAf
QRCXcyAtfTBh+/8u9GmxYhIbGRhQNv/LQ+9549PIx0abzIlpK38GA5ahYWvkfcY/
kxBB0k7oEHIZEEgspI6R32G4zoRWJhsH9GhONtgGPVbRlZ9X3ZNlVKDxLOASZZC0
C3HRM9pBKl/MqcrsiKFoDZHtNnlFiqIx2YbXD6N2EW2n7PCMo8RCLFcvBdRtWbiD
7P6cXyEGLt8ZvJBg2ISDTaBhBFWDzzpylfjvtjhDe53f+ExF1qW6xxONxLJGhx54
QrDitkr8IcyD7P/gYd4EkzOPv1NwqtKs8C0kxW0aI0eZO1p7eeG7Nn+CRBCm6fsc
8JKt3/y2xO5HExAN/Gy2DBVrNWBX/7PvPxYcND38jnEGPWLYBbRCaesn1v7Gx0zy
cGued4xKwblF0YR0hvon73f/ORMXoImEZiJ7GAVrEYQBtxcfQMX/70MJr6uV5TT0
WgdngOrWYsjJ4USDQRqDKVovBbsDEE/ie4u5zKL0i2ge5PSYC++Zzej7l7Ybf6XZ
I3ng1/WI98I9vC2qB0omploaopyIjcb76yQjljtJmZtg7KW5dB8O3iSlfrWz6vi9
O1OStfcvx0XeuH6jhcK93qYZOwXUEeYqyePDpEUCDOu33pTgTwrog82yUUK5dNCZ
grgpumSyTTbrff9tk4IaIhXBdaGrHaYX67IggEQH7gHAXVkdbaWdS20yR4clG5xI
II9O5YZlQZf3LOHn9FT/pvqdL6u4U5pZdEiLT25OYOz4qeUk+j71IQRtavEY+D4L
2Kp7NFLQLtHZRlZ4aAUNb+iQVjlVD+DGGXwyjjd+Zu0s+DrXJKKzg4fvhdeDncaZ
nWGJiAmYQc9xOqJDjMLxEUcYd5T1LXa/wbrwAgy+fXpQALS+Vbszp2QywAZj4IfX
uVpI7cYWjL6YBBAwxvjlaU1lSN+UJuHYdtzFSKjXhgl79cjIWUp+cMhxeFzo3yY2
+8svzhG8m2fXw3C6z5Kz8xytXRrjp6g/KjshOXuVzv8XPKRreeVB0KJm4fXvZmbg
cnRbNya2nNvgODegj7ur4OJl3penqGpOdECshPEAVI311L5CfUyDoWHEnki/eJW2
wWymiiRbpecDWWhayojsjbOORAsvp0w7smbebd+AbjM8zgLjbRmIxxi9gNpz/7cd
mWaDNB7czuDjblncI0mJezD3oMV28z5UJY6cqMv58rPvOJvUmk3e58efioNYc1+x
ztHBeY2CLwlBctHRWTj8qJOpF244a8en8dvmD5JpR0KefohDAUHn8SxcCHQrChfG
ok+0LOol9DMJD2LFkosiB9pzpJ2n0P/YNpS6lPjz3m/ueA8DZQHk/t8iUGnoSEY3
SXbcqe6IOOwicPJLeizAiV2BOppnJgDGo4z0xMWShjlPNtkEuGQxJxnJpCBIIr8u
SpZ1OLMTJ0C4RgxyRw5iocQm3AMDYjT2+C2Zsf8wwSJWkarntjuGnEk09sYVwX7n
w7Q7XRI6VjfQAtb97cQRCOzsOeIIljhFCtIrBfuR60MypfWIdYgqodwsLv67TBEY
dXDercyNYrokKOb2jHhuM0p6BV6X9oB29bz9QFHWBJutcjbBrZ83OwAh6XoTbXSQ
UR1TvXDG0wmG3pAUyjDKMW3PEH/WKkHKsw6NSS8ylBP6diPFHRCGqGpP/AejUkCq
ib6KJC/zAIvDdnQUd8QAcwDiIO4XuePVrPeFw+5GoSfJUKDtxK2/97FigY1pSBaL
D4SgJoLcf3/EPk/F4MYTAldIoEnlphHVBcSRnZzE9bpeO2E4NjcAmNj9NYlDWa4I
nAqsr1U2RMtHNJEjNaOG2+Co2xuw+wmuAyqYEt+tXEftcuHNZ/TlN8FvisxYsFzv
YGG2j2OrtByrG7RCkwTRgU3xd4CHMsnf4S+1Pqk8/m0DpEQGbUrK3ZzJaCd1qREg
CsKDAjtLCPNdI8WjWFzPaPyu9ajbX7V513/b4mxmhJWfUzlaaCoPRh18QDNRTzxz
jXqEIgREvB+hHLAZ7P5fZiYqsAlEt/40hJjyBkHAIivuIuIrLrxNTUCc3jBlVHec
mLxXb8fPQ6NtvIlIH/ua28Iv67jDHXKN4U2+MnvcCzrvnHvbZ8fgFBvN20JdxU8V
VWgvV4k0Qv5AXRR7bwXgfrgoEmsf2xKxhLwXGQT3eu8JKAZbMrQcvD+ShcXLeb8i
dTndltsnlVGWT3SoCz3dPwU5OHrJIwl3DtSOrNORy+0xc8Tv4+AoM4fTF8W94r+C
OREBETjHYOUBeH5F/Y8pQOzmCDCOhsCxCi+SHyMKgZmwLWP/JHBA86SEX2wP6ptZ
gq60TgFFwKg+CNRfmStIf0qxJEe0YBVNn3i1PjYq9PbLthvfo49Sq9PB+6RkjB+R
7h2VAjbOQ5vHpaLkG8A0egn3boTOYhuOXv73KQd0YQId2K0pJdekBl9Sk4G2cFIr
n3FtjWVEqGP4bjjEaSYtQ2M+E0knKhEFc4pSbJVI4d5OrxJ7Qcu8q1RtIjvBGJzc
8H33A85wFu+9ZSGEd2iiyO07j9yeaIfxCobxeBUTzr+f7utVuUL2A25Wdz31Mipj
`protect end_protected