`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 57664 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
W6MqvulZH+WIzeIjX6w8v4Tm9mPnc9jZ97Puaqdp1jzycIrV9vWUM+UHxqWGvlAZ
7iQiTsLrnByuACehuJjdruD/gkTPGBDJQ0xbDsLre76iWdhoAUUBHUoNAax7xzvr
nm3mpnUSVfHpwr9K2RDEWbIX2Z/9TtcLM7KIlCbm099Iv0mi9DHt8MkPSd09BMFP
djue07NfSvZc66BGY6u3bTGKJc+6tiVj0dn7cb8prE4kdK6u0LvrsgsFZSkatpsC
4veYyywlaHcVeYxVCB1/YfHKbbRe56oyA2nb9l16FPNcWo5adVTP301j/dGJA+Ws
edCuSE/XsI1Oul0WFy+6iuQ1tdBN7+NKVe1MmFocD1eAmjWZZj4iEr9IGeCu40Dq
ydItkglTJkyryCY01EARtRQcM0oCJz9fs68mgYC3D2IqpECJnG0la4oGURNxoj4i
I4mF63MTGgZu8LQnKuF0djdkJGqbYQi2dRSkfKwcqQUYliyQ+e+Qgk9SiCPNx9jR
F94NwTpXZeEHMpKQNCUdSag3QtD0i/pu9laKXRnCZfxIcLsvrohRGajF0o07TO78
rFMQF2NA9ANjlpPZQFOodfchRAODRROTfqbu6u+MVa//3s48wJxw0LMgKgduZPpv
LS+983csbdXUoha8WiXkyM8bynuZgZzAyLwlmTKiKkuX30GOFxFIZnvXf2y+9zO4
coSH0/56vHQl3Sg3QXqkJa6Sp7aUhXKckM8yoUJySRAh5qrGM0Vwbmrh2QEu4YaY
zuNx/JvmWDnUE5d0hlJinEeOzWXyv08UtsdRQ7PJXIqFf0/6eGBpVhDlgWSN4Ezd
IJz0md6yWs6q5ZfzQbMi8T/m88JWQ2pG9GUXY56VU4EyWH8b9eDOTx0dsF/U+cDh
vtAvE7UQKWcgw6V52qJ5o92zNAyQMaQ1POKbqLJhUNsnGfyZ11u9vN/3twVNOTnb
l31l2bgbYmK48OiNmdAf7yoAPXeCrgXtDGkO79JKhAbf4nR9EpTMvcKltTwtBmnD
+3zrwE0xTrja4FFFGbDO4zesm2ZdIHZzocKY9P3z+uIW9bBVdB/dWxCqXLrI4pbC
QElBVKmJH3SS2MVqpWwbyJq4fD4hVGESzkJ+IY3HPLtsTZ0+rgl65F1sKSTnUYWC
cKKveyZEyxSW1m1vxtAQVAS/932Md+y2Ss4a4vpldte+6MR43LG7eaC5DpsEF3iC
AstIoS/Dbpan+SsW+1QE/46vpFptM4Yh0rJAIfl29St8C3MBo5dOrXJAHETGPuzt
LfKOKg5NPAM3NTAGh4xCMAZbNOyOMnfXp7Do+xmveMgIz+YvyBpGeTXHWdUPu0IB
IzKYgrURSNSVhXpYuWFUDm3FfT8IzHivWbNYlBdf5QdD4oCq92c7Ai+b4lnWI81B
cKFI05NQT/MRQnW4L4NoWbiVPLuTHLy6rgeBt95/PAzP2BKZ+NAak/7Vt9NBcRPT
wHgWcQRX3jRAolkyZ+nSRyppwK9La0qC+353cIRrmSywr82lifUV9OLXXm4f9Vby
yJiHggTS5+YcKl7QB8FFGWqGp1HqPZoBwNcaJMthU6wvpKfB0iVxGB2YNBFulJX+
/qE9j1kPZfT1+IqgHxrEVycZ0vgKmkPPxurbrxUR/EFtr+OuZfsn8Den/NDjLEC5
1dX/7rvb05E0EiLf7moKeN2ETZvwwnas9CdXCG0P7GGMTpRCL/S13nDZg8u2QISE
7w6MGH/lMlBpvTrpCsa5H4XfGO5fMxfvRi+CDNvH63cMFCPK2O1yC8ly7u3yf9e7
KHJIhwcte2hV014wzTyZdjHD+Kt3goYbh04s9TocS/Xjn2Gf9abJni/QDPVC21SZ
Cqv80gusY8dNJEtq9Hm7LGdYPcfGuPir/YG0ldnCIWK4ENgIuipMF06WRBeIB7kS
gDSfyyS3IG47hSyuOAilG0B3n+bd15uztxeZ/DnJJpu87p3/0+d7Bs0mG4/h5Ob/
M6zFHsmyt+N4tOwMQy5uapteet78Cak13AkuUik+Xq0P3Nzou3UjSaBh7wAbTyOs
5ESR5tZkAKVRYLxD+Al7/gTBEpx/nuJINZOX3fFAbcTNfcDVZGAq+wjn7BTwAsJ/
ZUt12e/9v6E8SqidoIdVO1BjPflsE2xjddqXKH+JNWQnlhdaADboh0tDl7xnE6Z0
dHhJWthIKFJL4MQBGt/It1v11oRruSPiORDR3PrfQaB+0WpH3sPkmZJLlWSvVwRe
3AAqJIz+nGPoC76Bc/X57RlMUEcIoNJKm0g9g4YUwwLaDuc7QuoVljyCn2AesHgM
KPn+uOdHIeLBaIOwkB93LlvFmUOrzzOLubE9BfMkEOsu6Iz9F7MZnT68MIeo7yAD
YT88WiupRjYx4S/745yYe49Ff97OUP8ZjmIeIQcFbF3hD2QgBiPUz/DPiouXUIhB
7G7gjqyOdbjY0a8x5dPVbaxwJrU1At/JIilzxs55JlPQJyjGjXY+y3eOaPdtXjwx
bn3Oupf/0CHNMB4IAxu8vE376dok03gfT92/gsFEOK1yCLzmg9ipWAmS6VvR72uh
kZ8os8khdHZl8JnXQ6ls+HEnj8N2eWp9zqIqygG+5ah2CsOgD6f081PVxtLJZ5uw
EtzbNP0MnSwk7p8WOPjrTGbicMIlKX3aOAoUMls91/OcEfj7Dtmx4eSnP2HB92zc
qSPEjpa2tl5tndBAFC+79IFjmE5T17kbsuaJY7r0t4OJTAPeN3axLOz/yTF3A8sF
zLkHKBaHC15OWrlaGxvHNwEzVCRPf7uUAZOoWK9AbUhHoRwqxpe3dUZeEbeeIe6i
Gm0GdnFY/7MU20WjiUw+Iw+Mo7VhvViqwDXYLCvp6fNfCw5H4SS2G4U9lnpLrtoE
i8ScTrIG15cy05E5EU2HSIzuu2p9D9jBqSf10fpNNxYEiQUIh2nfcw2z9uzvTTfY
YGnU1vijo+8JaKjGgMEoRcd4lmsyIaKScr2veSeDAEtb21qIG8v5RRDhwcM25I/j
RW7Y+Qc+SK/MATdloUkWWXO9C5QBiPhnwo35ZkpGe2mooarlAYoaYr98uY4Sc43H
KChluXCTwn117kIRYD9wSBsjUhOb6P16or0e+PI89AWQHSANaeDfBlCksRa/5xo3
4LF0DUGiR/HXzVel8hTp3Cnrrp5seUy8xjvZ0DA8Z40BWgabJ0a+8vYRedoq2dd3
fIjmq3XffAyB1FxpfpJdLO0OP4IR0gk7/JJPK8DGvBAe8/Ao8iptZQg63+nxKa1s
UoFVd1+jMZW1+ybWXW7nXdJPZHmmPE0E52zL8gfpJ56tSVCMWq+3rZUxMWLjFkfM
ym93BsSCQOKwy3+wa7s9JUT5gz989vOZaLIux6Q8FqDfBwymA3sdUAX/J3AIpK83
ILkJ0ppHJBAGLCpCvbRo91+xH5phy9BDzwEtZ8YaDaOG7cbeDkvTvg4S428cYEsa
EQy5tRSI+ckUm2RTAqVIIxZYS6Tvi+a6O8j0xXo4rpTOEvmR79igAxT6NvVbl0IW
YVAxMtV8mF2OhfPdMdzsgwkMnZ2wha+TXYriPOgDtLye31Hpi3fmVusyEk7cQaoh
M7FD6c4nwLgiSr+5J+ThcycWNp736jDXNTtOfuZO/tHW2PijAHPyPCf4yrdgAp/4
ZJ/ZLWPYkghYsatXyczKpIIpFL3mkBzBC4jM29Zp6aZzgCS70E/xvq3QvdMOcFf8
lu3yDvhBJjB4Zz1IJq3mKAyrn3XYzBqbidDXSnyF21tJH7xLuZcvxTogyNxQA0Xi
i2omBaMqElXo2fZjp78MFTzMOPZA8CUEwgUWI9YycLKwj9fZolRakQ8FYWhE+AfL
2n/7f4clgVbpSG1APqARazFKnFKXgbyDbfdSl/4PvRTcH3hLRefQJ0/WfwC3LCmL
sNUz2LhNFcaIfmmMFcWQ1Ht5lM4/lu0PoMOIXCgWpTM/yjqQSJmhDPIUCkPyOnEG
TvlgCZtpnO2D1wNgpGOwDlAEcfnoXHFpkXmZfkfBWYLNh1AQ4Jz0xc2GK3WQcsk9
vBSqS1IcniKw7bnsqiz2+rJuauWfvpjuguetWAO78Kxc32mSnLZcWPnIILTjC8Yu
K4NS8+IEml47gfcU3U9uhtWVnTn75haR+/9dI7NxQybtML+lQQD93MIXG1mCCCid
sksvYj21AtOdq1CB8LJbBxf5KQDx9KTfuTZgZU3bcbExlWPWbEtyxkwG6aXVIpvu
VMw8KsxFQCsXltVGAjBrC3sgQyIjBBBFVQ3wt/3/seUAruC9KsRr3ShWWkmdSYpM
VYjC6QdtcmU8MN9ZWeIantbuNZum01aPXQB3o6ebnasoad/Uceex9aaMfitVFz3a
BYmB2pOCKuh63JidKypXyGNi1YZ76WTVckvjKvNbx3YAIscttY6YTDyAKKABHwZe
N1acg07fJcJ42XX1jbKr78EoJuId5tj+F4eZGLxbc//QtjBr/NcS996x3F9KtFqP
VQ5U9qb0RUvfFe4yS+4WlrxR0N3V41HwdQxlqIfwbJFwxXocyvvtvat3PTY0DMDU
ZAcG2WpIaRh+bPRHb62GZwVLmQhJQnmSRbPjfhfDo0aR3bQj5YKQayU8DBSJsPt4
0DR6/52D5K2udamXtaA5ZB9ZnsAvtjpFBCUNNzSlSP+UvLPzKt1WqiaTc/ulK8FU
MMmWmDI+wHnNiooYTGQkkz/vd8Y89rp1cCWQd5BZFulGXuiHDh/+MG0eEdSowz5l
6spYuugRDiTLAG0N7bw+X3wBE8ZJioOULoa3CUbRFpvWzmC5FTCe1l4qCb273tBB
qZFQam/mphWuGJwMBuKNffoMRIr+h1cqJaVFvBnyusYa0mYutspJL6Dg/SpxTzku
NAiCzs8R5EPlpQc407Fl8LKXdScZzHfgise54lqLX1aRLXRoIQXIxSfhy4dm1Vpq
kbuhGGeECNKDTjpMu9gdvY95M1UuJuJV+ZThL6LwJOCPzOsGsgb5g1BzLRA1HpVr
bzInN/p7yhQywCBTY/7d4j99PixobW5Mf138dbbH3IVk2EGqE94zIAOxf2cJCfwC
vCEI50lu8LUL6t6Jujqb/8uGJJgwyn034eKd9EnAzHh9P+qc0AEmLSdSk5SCnyCq
u+XPA8OGMqvbLEfSnWTlpkXpaTcUP3Ir0RQzHsbNl/XjsHZ07Jw/92yd4HkyehDz
MzB2l2zTw+e9XoQ7FiGj13DgrECMjL+f//v930Mmq1t9/D8eGcnxAJyrE9ESQpTN
NR9aJb3R0T/fESLZwhLf2VmU9qMxu8/wi0Ix58YL3aKuK4PjYjDQjrmf4VQEIPpd
PLtauPDC/7s4NryxgEjKNI3rR/mUIr8WErG1/INK8d6JWYCPX1cgHziDlfJWUhTz
v+Yky1uPCYaxXHPIZWWtpMQQQ90MRy+cJHV0HoGbfuZD+ASiGTRFQyBkE3CJzp6G
z9A39w9fVV3tbNuyZVo8+31XMZFbb+CpZ/oa773isfEy9RsRHMSp+1LGPWTe9HbL
rjb5tMyNqjVa2e4BLsySmq6gUSSUnNEyzj2ZOlfHIRUjn9yJZV2SWobzt2TxTFyl
QR75D9oFqu24zzoot4qPXfUcv/6VuDb8uMCfyTy8UkotiLqeggYKWmsMnpuaUfOo
c1OXS8nvJAR/rKUgKq7d2jaQ3WYoR1l0rmT+VW48KLwFQRMpEud5xTauJChAHGiI
BERfkmlyPvWKX8dp6r4zExaU/bzkpWQoLRpVxK5IRs61mFScU1EQYuQ048oT2Wq/
ulGFVBsKP4gZl2GwRXl9cJgWzdPVwhF5KBvot79pf6W2mYY0AvmkKzN3AUjSMnS5
cvWTZbRqtypGix/xiM95dr0I5rYUZJ4rY0icZUHhkPkIQ9Yu86A1q5bYvcD9sp/4
9VIZkZErz23qvdEID+pMyGHxVx2fhnlEHuQVoI5dLrwZs3WWWlLenE6fB/J1a0r2
DM/QS2zo9EKxy76wA3aR16oSQVxpnVQRGO1A6+ZIOcjT44xvRMj/0jlkxZj9H9cF
g/I26LSqDZGzeXyBffFpcObZ9Jy0pTM9TJxso3e8RdyJnJfS5hst+GqsoLaP1jeb
/ip5hPfTThP8KZQVV04l4PJyfofcR5VUPSiLXV88ExoRcz6O4KS18rHO4ZjqZUbG
KOe30wUxNgA/Yxv5A4z2W/Bjrwpx6AbAl7euhPWFHM5rOJw52EaHmYWqTf5lCeLh
Dj4+juXBayP9B+P1+xmZbJ/jhG2svEDL/kvMjNBXAIP26DJQMte9cwbBdn7LDDy1
F3HAyAetG5HEUBoDXyj6jc81g6gzu5HPKAo+forOnB5AbZTHayrxDleFEzbHxOr5
F+Z9kuo3U1bmgsvUuucYEvRAVFnDz9/WSJMX89kSPJ4H0cSk8erCz+iTzTXMG0iS
6SqihG5qwXwPeR1vKb9sxTN+490ZeYomy0Ha6UtrC/wtRUcITNk/VOjthoRf1U/S
nOzbSkLb4pmeaLQrw5CW8hcZbfkkf/HjXTbJoAgiX1ijHQUhxDDn1PFafip3hldN
+OwhpcKSRYsYe9NTRnaqqoiiSuYjPTIIq75kOH/HaC5PKrk8y9M+MHMsgSG/zsbg
BmA5uDhi2dPc9Y3bmq3WNeiBqXzbwW5oI8c2cVTJeVCQItIdh37kWAL8BDgyQHlB
19b3PxYw0aLdSLEbB/GfPb+LrjUCFZuUlc1mf2JzGs1Ws5+9FwEiuSJZZI0QHpym
DXnDxgJE9sV0pyBSPMkfp4kHYgaIuip7LAXsNC6zfN2JAFK8P2bgUVTV1lCFHvVS
eQR8YoGH0AO+fPkCNAEybMrtm11YI3k2KD6rKGzZmr3Mqu5WdeIGVhkBITFVE026
9a6ghXeVjn0wGGac3KxmXRYmkwBGd7CU4EUNKBZCKqrmuXpKPmFZ2vWMQ2ovXjaf
lw4P+YcTlT2HKTNp1iHp/S41kWHevg27Fs3uNAmiytHe4OXHeZYeWKMrItwho1lR
BUA4yCmo3BEnOXXPOIyZBbk4X/LSZH3EtnSV76pK+J5MqaxF2X/OOTmf5wiEHgYw
SYaw427oBgOJn/sRyAP1sXOGjLWBi6MK5kjb66keZ0cJPwSnUTNNvBule1G8QAng
vQcxBg3X6eIl628Wns6eHBOU6v22twpGaSzJFSDm9p7tJI2MDcnO+XL9Ev1wFQTn
qmsJFqMUGHZceatFaq1qvktflgVnyswbkbv4xZm8rKKPlDvIS9ZwnzJDgIZmzBQy
SBfmEN72A6GQcVFwHkxGZjpFzUPJlvyH/K5GbrLgRqkKIz1wjKz+zsjXwDVEv059
CO6s31Jpp4O+cBEP9DdSZY3WS1vHWuBG6A8WjtUw3DGTrxjscsU52dr+VdSU7BtV
5sWyEiKHeM5/k7yqa895P0UASeuoQjJOFeRfKq7pHrRTWxpCggHQ7On6F4bTelQO
EbpSdDwwb3MayOql/SgrTTubV1dPhnxUHbm9zVgKI8bLmWDnJuuPoKODyvy89Vg9
ZQX6sUWIUYVj29MyJ6KoJb3VbBJc7nTLZ0Q+ykuCsNFuIVeLrfT0YJb/IDLZRVUV
UEu06qfoTbXETUrDp6kKMSc9+ysSpoOzR+YjNvH7zfFddisF2c0nOyJiS2rCN6ky
MZrhHN7xB7QLHl9/b1Q2bLE9qf+8bbtzhFKYOBdDCLuCZDMQVRpSwIVt6Dc1sktE
sjviX0TelGmDBL/eu0HOne3gp0JvalGD4BY1KE+Q7k0ewi2HWv373H9RnVHXK6vK
wNbIYNL5zCPxrlAseGfD4+4a/z8j2qvcWtR7CvEme0LuMv1xsCpEt3X4TQH06noa
PeTw1B+4sGxYJ13QEr2+26pqBtL/b52M2xr2cy6sTC4bv3Rl+Vget0+aO/3qJqYE
FSwFzWZAXNAPl+pGDQjTHISUsfnzCaSvV3ESSIQ9ccgScVfohp8Yj0rllIc+5K+o
0j804ZWzZdlZxf7npUfYrBP0K5bwspBpwqDz91iR2/UlXc1Zm0zal72YFNjzWmUm
HKJpk+xkBHCjPztjgJwOHYukJOCny99DpJG1dlCNcYKFAdAVMJF6JXwP9GgB82e4
4FHriEDIbJQwhmg/Zv+hjv/wl7MScmmaAVr+nCaylN8oXElFGr7lFrQNCyN5TY3R
gXLgQNpKi45lPchnMaQI6Y2hsKfFk/UQbEEwa9QhnQF1+K2EV6UVzbDXRde2N8EL
Qcoe2oWjN9VKqTS0LI0tUkbY0ocP2W7G/Lg6IcAHvZbrO/FQrmZn6U8EepJ3rVql
1bVfHyXFzbl99Apkf9T7z/q6Bxhz1SF/zLhehDCVFLekL2zoarna0GEFB5uCSqFG
zqYqN5wNjIVBbCegKbCEaYQQMJfx5X8CK9UcjkHU6/iZYn2rPuEQ3CFz3R6Oa7W7
4ApCVZctLZHlr3HqGFmIcZboXWVskE8An+6AUxLWRc4nK2clV85jeaJKGWofRJNj
nXkuZFGx2WF1dmgm7+89nHJQHTTvZJoAwj76cJywgsLs2GnJd0pfJSodweCB0Z/V
qzXk6ivfeRqRooXrU7kckvX0HPNKj3AkmbK9/gOyCBi3oFU+p+ecc8vD1gpX40QE
cuHudf4MoATsTNAi1KcSZQwqsDez0y9AkdCawI7Lf3pdZjO6YyAmeePOsMZy5zLq
wnhr0TvJrMEW3Baf31b3HLKbdyLDgNq0FGkjbVUIPyO6wRaVqA//gtAGLop2RS+4
XD+aJLWhtyY6BX5Ad/LMulQi/bY01b24vzLr+MdvYOmmi1kioS12z1DoABMt5blA
+Zu33/Pyvd9RcgFX3JFZXCWvkhf+y0cOMEHnZHwqgXv6ZaysfsZPW5pRE2HSfYHH
TFTt8bPRfTDhydb3pLn4tNIachgRie2A/W5BdeJO/NTZUZN/n6DSXjYKGlOwp2i9
oxsyzomUtrECmZ8LqOkE3ZuZIgRNtq+kz89N5DmqEvOJmYMIN6ZaxSm2GKzny/wB
PxqxOOorZJK2m2Z5cViWhb9pCZS8D4NUkcPcHRLJe0aTXmZS5iJvMCOAZ5A1Uz/h
O1OiMoNmRMRPh4My5Hs22413ZQupw3C0nrtuXe0jSvcq4VoZuQo1abD8R2oGMm6R
o3GjLPCZ6zUQ458AMkQd7UzxZpT1PRLxc8di+gU0ZGsclyDWR4mzAHhPkdkF6SrW
QpXXtkHNkdJjdIH5cYjcaFrAutBkvJ2VK4AJEc9S1qc5KbQf/dyANAJ4S4AVw3lJ
ei3Au3s4NX3kSGK+rRs8Y7aCOt94847bfUsz0wtgsRoH9hreQ91REQunzp4V8viW
g918o6UrE1LnnnEOcYqwlq1RGs5deYzo4u9ntdducW317cIe+mOdmltq9Emya6db
H5n96cLJaTJ7UF/selzROFLSRZqQ3Bt7CReSqjM1SIH4jnWF4SXfbHQq33E7lcAI
8nd77wcOK8FhWM+HDdtgybSwBd4gh+RQ+gEESXWzHXmKUw5AiQGUmZMMMWjqSL7e
HzzXpJApijzPeGBqTXI5KYVFKW3SGdY3XCwtYJZFUpqaxxV6UnqHP8/tIiU+TyZt
9ok7x7tTS/1GwFTwahZwmGn5mktQgczg4811re4dnUn58IgEtlPvRnF0GL/vzA+y
1UPYOYoer7uJfRrvxRqR8PmjkXv1R4kndAsfkVXll+AqQiBf23zB31vhSxS97Aan
xISLTwTKbiXFqHMBW+RtQLlg/rrGKOcr66I3zgONGJVykMApgJnUnmWT2pRfUw5T
FcBM7B3aG3wyI6PK8cHoohKEBdtehQZ9X6dLhx/j2FBV5n9wRoVEbh2VqKPro/rB
Ba9s9VE40/X0Ek0TBdJs3dqa4BKiRUh2z4sodXy4+2LcYXyqRkJe/o+mxp90gu30
ukC63ESXWTkMy7LO6/GxH94gwkykkQnK4pfBEuzhVso4/FmxVUFbQPug1npC5xiW
qWyCqnFzBkslYtJ4LRMcsKqWpt+fIi56wOiqhPde3ja412+t/2KraxN4HAqAZloc
eAVorMBBQlytp656ZRVUkqL9fYSyYoER4jLGxkTfHE3uhELKmgrBReA44NIsEQJW
Q9k08wJN1n0PkcFQFFioR5WCl9ojnDSHMJmQmK2ipKqZLEsptVb9RlXvTo8da4nS
8UuTzbiR46a7X+gOtpXXxZILMKWAeIsjps231SUEiPvwAZxTuDUYCxfJht5CHAS9
lvWd0l12HlBVwKmFvy4il6J8v073Unzb/xMJnJvybZhIOm4RvFWi09O/pQkgx8nn
sDhh9z3SfxTHSZLtLVjlWS2fPhXUHAIok/V17HQY373crZmLkSwOuw1oBTXDPl3a
W3+SMvYOvSx16wcs+5asmWWSEMqWtOR8b3qc1OiLsHN6kHLJ211nBuFe7eJ5lYOf
tEq02OmBfIY7X/wfRp3BDQvzz6SOlzphZrtCximwqD//LELVm5dg9IFaXn9iP5v1
eSq/cFYVAQh9sNNkCb1BTn91EM8AUEkGcmuBngeTK7fIamxIVu++dno9+KSKW/AE
YXYG4U5/ngY2tbZ2hjLslMCYka1jChijIIgQCa7pCzf+okKSDF8v/F2TlbjXLKIZ
imFDJp0VDk9ZEBmH3VgNksD1zgYs23FKSD/ZO/MkMxVzC8FJdo7ByZcjNfM+hbAp
BUgz2CL7MW/5vcoCdEUbO6Qret6GGbf8q4zS6300rHFIOkPm5kF43d03I6LB31fH
VN52yYkK0TZMuKnFqYAfsVs0XAqWZpxuJMKCQ8kVjtUguXUpr0LiMK8F0b5wtWNU
nRkceR6BQ4VkDBlbC5+rOtRV9Egd67HfvV1az9vZB7Fe0nkTGBydgMw9nF67LPYr
cP0fYbmF4wsL6cnKTyreyJUX1fx0Ri8gEFWP1ID7EQiMP4WHdWPk+Hpdf38JfWXy
4KcyXWSc2Fkze6PjQjIgWTZd7wwuv+uW+MeCdwrM1cxuactosTRr5jo9B46hkZ4R
gZDg/WD2sNwIRjacM4YlfB1Ndp6qrQIgVJc0gn0c4jshs3Y1JdaDHXsjdETgcSyL
uwiOGR1AdR/z1O9TILgQEzFc14F/1pJ2/2d3noUg77I6ZAr12J5fjnyhPIUJRTKq
4q1BwVIyyR3LN7mgau15njvPjOD1X9IUq77BFOjcGn8a335Zcbe+v3OVdINFxREf
iK2UogRoN1z/za1dhLiuOunQeUkqXDpDZU8gpDv2Pk46Rzm2eUFPsZzHNueVCtis
4RiEmsixA/Keoyn9uh+KjRM7TMSx0ep7OFy+neEZ0F+HCVATU2dY4iV+cWrhtb5A
1+Tl0zdFtOr6xdRWfdZMJRKX8m43GKivI5y3M3lCOt6+EWOSJxR68KVR+rmcbHBv
H9NCn02NdCA9d0ae1PCDCpoUJZczMAmwgBYjSLc/106xP4qYwAD5qipevIoScHls
FLMWaks1lGF0VjEyH+ZOaiC4odDh7QC9nb0++GT+N6F5Od+rBbMgRmU8GN7Fc9Hc
etmTvNI/SHtLbJxqwZRphZkJAjs/uLfa46Dnbf8bq1ClfhXsVspQiomzX/PkDPSz
Tpt/GZQhplON280Yt9czdhwZiuoiOOYmOV2nq33lz1YGVe1/3JCHlnZ0WSXxQbxg
Az5LCdtm5tfu6+S8JM7AzVYda8nsdv6jtY5Gl8Fwnnkv0IMFNxXXATjusQEQnLfZ
5KRKWe3ylwuSpc5WlTXmR7Td9IZgnReXSY9o0g4YcMonbmmn/DAJmEM1dxkebo7S
04LBkIGGe1GA2votoCM5Qs0Nc4YypBpqATS5kOZmn4fKh/C8uSeo70Jx/lghcM7M
w49XHSpysi8u37KPXq7Lhwj5EhDrTiKu3AhWOIhqpzEcKgRSX8T6DAPGYiJb4uck
Ng0nM9RxAkePDQOjwqXDC2diNOkTRyJaghFrJNJQsCq0eWwzeJ7Al31owOeykGWN
ihTLiuygAZ3ZEhWo0Nf/BjOoXmD4aSLTXgICxdm5WqtAPoAGR6jo88FS6LkjkHlB
fYalLgxELVRvC8htwNWAXyYLVE15mjgT/rsRYiPhNxhzsUq7ylLxy/pEtfGfgAKa
mHH98sIg3q4Mu0+QKyenrOr/JfZsDpEbGDPisAIMs5Sx2py9HSZ0SMmTap08uElC
PJArNYhTJWg6JW3bz2Pauf+mI03ddE0BlO/2wTJz2SFMJoEr7RLSrQWQsXAqnrS8
ulqMEu+F5x5YvkrDd5WIzZoxOjIYY+apxC/zGeHk9OlkwWfoAFZnb5/6bnS+vMvS
eJGH3+eSbmBUhN6AgyRKYodWnMzyDoQ0/wNsFB+jBJEyhDYD+bhRmQ1J7nt4xzCa
mnDfPtYOuXgIgtdmPye9g1/2CmGSF9txo5RAbjUonDLwtSKcsGfhNofy1ngBoDA5
40vOMC4/Zd2aJIB5aSPvNISFacYf6unm54F7v5W2J94AEfmkg8bKsbxt4r/+tkwf
maZiJ66zB/75itZXTkDM1xh44Yl+UuOkIsclXCjtJ50MntCd+TtS8nVorNNgLavJ
UpjGii1ILkVOtXkE6kSqe0/jeupXvgQ5AuLc9dNoNfYeJ7Mhg5JfQ0hI+u/nlTxi
WCDT5THaIpdhe4WmrrGwy5Bkq1OfgTubkkTZlbEyNE7ye9/dh98dYBRkAcOgYQEe
oFcQT1t9kAFMtzTwBq/k8MVMo8h51F28nkKo3dXBgrY7Bc7EgOsQoOZhPWN6dQTc
JV77YjZFFFFPHi8tn4yVpLn2zsZLk3eE+olQmXxHO0BW6NVliqbakk/vWCyAHwC1
cI0YlgZloEuAkmF5VzaXWl1AJUSso5Gz7wugl+JKbXKDLEdv9vLTDdLPSEiJ+dKP
KukzxDef7AecYksYo7IlBtlFYudst5tOARcWSRV7IYDxsvgZlv0ktNOS/eqOhbKQ
adO/gYkU48QAVHVFmcpMP4pxKCrL5rKGtXzS0zN913dfIqgG/MIsTcDs0vcArlSW
tCOeWL/fJXjhVx5UnOK+oTn7sIJIA8qvphmUiIZhaZ+8eyCWsySoZk6dffrALMlX
Do4CQkxXPZKzdEBxSuMKm1hQA4k2fnwzSAl5UphXwGUG3yZLi8+2EAoEKQoz0GBn
ASzjI8BjW6DvDICYOyXdEqzEafQj4fM3v/m0pSBrU+WwThAJSjU2BPrPPfcNhfsj
4rA+WwSa8xvH6VdnVJKlu9eSgY0i5Sg/QPrb/oNR32pcfVkuwHafn4QtZzWXFdvE
MAqXkfuy51CtBpIRu0J87QCxyFZMu/bDH2HhvZ9CpXtE5sPIL4uwtfi6sQd83/r6
gntuedP6pCXgBs1CU3ASBEkM2nVG5W1LLlHNFuoKu8DYAL3U4T5gLbRN7/Agcwp6
J+8X0YPU+10eyx0T+4VoSZSmXfysOKDxxurk9jGYJuSN20Tr4/kO719X8V51pLhT
JP5I7wbv2SN1moZLqrj26I46CQ+VU+uPpL16oeIUwaLQjaPhufXbGfyQLJW+vg1Z
xqulZsZRZOglFS12mcUKpjHzfXPTUsTEiLbvWQrlCdQNU8UNrtGD4jEUCOqvJM9x
ax0Xcn8VAgdToCIiQn97YMdY509h+4KzUmhmZfdTBpxfA+rD8/rTT8SIFup2Wf7h
cVs5Om7jLKUeu79KCTTqcPrzt2Fiq6xfB20c86H6iCVPdkScyZesFTI/0OQ5gJAd
D3F9Hk+eWL4HS1BuKhy5L0zcNdNEu2lpIASjJkIuYXEXvVxDT3wssNm9xObW5xpQ
qTSl0j7kImwQV3/dA6syVU9m71EDVmRFccpeYK/XYRlvH3l3a0/7dRahXm2Nride
rmqV5tHGOu44dVz9EIIpOAzcMI4TdtcWqGFfdDMg/VFU9Z9lUvDnVsKlRTqFsq3j
HJLp4WObWSBTwPP0CQv3S1isWH8aFwqpUGpAswnNke/rGGGYUwCNM4GBhpElctNA
4yM7OPAklWWmJWHG+Vd2rLKw4brFzqRX1fOu6MEhGiaB4gEncDBVvKI85TDH6Y49
zglzZ8rlsL7zrS1qpvOLp6b0NoP4mrbnBweMlt7lB4NDJjDC6o0QfrIyX8OwUJER
sKwJp1B1tNc5JQRnNm17FV/B/xcZAwQe04Zo/czna9cEbvdGI/PLZKDPqNl9U5jT
Z0/ZENdpB/AXVLsvJWRdZel2k/QO08pXYS+MTX2ZG7ZkRGisnsNeeznLzKU6J4Cp
C6nZZ2ASPF6V+xiJE+c3tPHJc77iaFSqjBglc5+b2zrNgL8MMQknPB19zD13fXHZ
y21FTWfAayHyoiwK1IT76d1B+KmbmE1b5PtsiB6ZeA7srDKAA4SqpV/CyaZR8uwd
DCpFlNqyWcv6MJ6K7xf2JZVIZ/A8RVNj2spUnDrNg03DMba99VKPqKTT5ilS7Sl8
qAlSdxH+ZQqO++AxymqhfK0KbRGK+OGk8SBpGNHAUVGevv/1Mlp6t27bX8WSnmfY
txfpRNbkwnVwdovKULD6Sb8B6K8Idw4PyQcpIqZ1eBmyF6PgQLTE/ADcwOnG0/RC
YLnYdtUA+LW9qohhCVpgQy1otw+xgInmM/Qa186iBsJZ+VVo5IuBFgu3nYOtivlS
LXPMGHClXhCG70Z0dgcdnDjaywC0ViLEjmosR418Qu0yAUyA3vyHv+uRy0P1UkzA
nFuSiSkfznkW/MVVwaiGyjojIiyd7+mwCCIOW/n4Y5bcj0WF9Lol92EFCWb9CDlJ
A67dMoy8Cu0HBPmtJtU60+MPP26Q67IYvyHW65+fhRFEhXJhHRyeS/24FVjSnbLJ
0tuRbzfAF65sIctY1q0b/GZv1M0yFQ1xuxwHi1pKUqwYAGkPvsMc+KXycmHsxjvm
etQrlQslSMP6tLceaubeDlSvgX72JgE2H8jvQ3Yt2fPkoAtxirZHd4pK9+nwYYKj
3nq7oNLC6Fc1gcAN1f0EwgbU1JHRZl32sCJEzm6VyGwqnsMgbAWIKFgbqredHq8l
1Jcyxmu44En2AIfRNTfMZYJbbqUDJs/XRfSUQ/b3eL6Ba2aX9J/sH3pgYEJMw5F6
GPNoYa9SuNPGKed8xdGeB9eFBy03oXV0yoTDoQRwy07MoWeycFSas3FSDQjgvFmt
3TkutWtHmPyV5eNRY9d4d3eJ7NExxne7OswQ+NUYU/aQa/dec3My3tmm+KhpKV1B
xdVa0F9VGF/bbqHhXf6dShHXs2dxCME4wQMCKP2n/fOUZpY+owoopUbu/oALP+ep
IYgnb7MumJMkBdCtxXu0Wug6mghts2u/cNvNkGbmjy6+r6IJF8nn3qG2cmRoA3//
h3i+SaB3t1SJEniQTGBRrzNueh3gxrrjz2wMPUHJoHyNY1BrFZmqQxe2RDb4Jo3y
nvYjeuA4y0mSMSXC3hQdKZGINpFpnr3PD0nVIdT+jJ9Rz8HEX54Bl3bHTq82OHS3
qDvtgSIj8yeUGoBrmScfvMzZ50LFmbTu7tiX3rtWEPPjwwxU0/yi5RrROuRZC6Ty
dOFtFC2Ub9PxgujaXFaAzfRkewEN/XoX+3DNC0eazzWJu9yX76WlC1dU58zwKa5F
ZsD/TK258o/H+mD01q7z+O3aq59cZ3g2u0UTxbVKoGaltvHFB652P/eYwIie9xa0
7T05SQTQ9sdxZwPz84V/FLFYniaU6yUordl5chBiR3riYaoifVQGPFv87dbkPbXo
BAGMT1r68MT1HGc0V1LdSZRUgx/O0upSRc04hv/6Z/uXe9iLKzUH0YhpTA8qpiTo
pv6losoYQDRC4RvfAeT6ZpwQA3BKFUMmBC4GheiRBrtcpYbKK18V9gR5fjpR6daS
4rnmK7bsrCQYrj5J6zU2bi2FxdvULXBBt4GjUvk2iFq6ZRtiSBTpBMYWZo2SuEnJ
aGSf6+IzKKlwWrZHsYmuSQFfWAVHdpldJMzGAr7CCAsARTZyjhj/BHiARNpR8vmV
/3Vsw3QEgRLe8g3ofg5a/ylgNpkd5N96IejFEIG4PsiV8O8uAQH8jinkS4a/SVfd
mBgeRU15Dci/dB7vfneqcOahwHNZb0dgqYV4+qRMHJdx6u6TIK9LoG2xPjZyI3aF
9Xb3pkBaKZWyk2N27C5yr6LZNrJmTN4aQlmZZFHE6bHqumM9BfGMpR73uMat2F6W
zPapSCUH1+4NsZSgjQ5kuaiRgPFLLZHtmYEnh5G90Tj3BEa3Zxm9fC6062VD2epq
iUU7kh41U2tvBfDYMntXq1oK1Es4SJfx1t76XM9EdiegySHtVkXGqjynBEyDW69Y
DAT/uussLrCqRl/VhXVdetMhA1vxyMz27wEh+iIh4qzDMHNqtLaigMBIPz22ygq0
tv1Sm4K72mXp3AZXRQ1mM1irZr0CaGFKWO1HhS53n4hPfgfsIo0iTefWKrLxugzs
Xyb05QWr9ZHWN0GP9zu3KrQs8WHTfiEdtQvIMNwuJrzIx5UPDhrCpYVLh2pvdNeD
3wCRyZ2QQ4GPvhMEusGRR0b8yfhU30yQk50/WILPJWZ6+jud/WfusY6uVt+/4F4k
JHplqUua/QIjZ4JR0U4/ZzAeIUbn1Lb/M2xfja14tTYYgNrd/NWJA3k0UFApOIh4
EnnLIlwa7r3y+DgRWCJyZC3Fw3p19/YsXCYRYhyxMGWkcea37c2RPpQKcdX+gjVs
aoqsYDEzgkWaKvbC2t82936NbhRrkyaTFAlBPCIN/bjrkfgHyoQXmEnnm+Kvl6ka
f8EQsoZUbS7Q78tbLLK4cCZQy6POYbS2JDazDaUCOOt+J00pYmsL51c8d9zlcPsr
q60g2S5QvbQlRJQkAfwvqmhnlGdRtcqT7BiStgh1tb3HN5RK1N41qPygd4ioFuiE
4Is1RGw6RWg1MAtHI9rz9FnnoGdRJuURKid1R6YMWgwbTIndq3MuHPhQXw8pnj3d
CjxWtRlc/fyoEyTfV7lM/z3vwf+1KkV30eb1dSP5qHdEDp+E2T5ZNCXWNrSiztru
efs85RAjOL4sVd2ptKV60eRul8cj5N3BI2iu/+VG9a5weSTMtO2wNg11GqUPWH5i
mSuC1MtAcEdI2BsscyprOBnaIqz1nJy9xEsR1FU5EuKoZEn/AkInMoVTDkPuGx1L
Lpz0xlDhgREtbMmjoA3UHKdN7PaOiEVxVetGzGPFOpnIjTh7lXOY7mOOUKZF/Lmb
zgrZZ27msmIYfr2FnvqxytOttOdxHZCu9cdEx6lEJPykuBZNG47zCDGNMmYtvmLH
I1T76E8Cl2JPIve3nAKghhmT2N6YfGhIq8A5CHb0XQqWTuv1Njqhu8r3afvaGYC+
tMopciBZTDLCvg97FnwLydSBYPJZJJZF/qbmnk5G7hdMwj2D5lijs2ckdXrNP6zm
+me8FjdOWb4DJFeN+dT2sUaC7uQOGfPjWkd/PB+zjVLRMXWAxnX2UKHHkfgS8mxH
7PL9OV9KUDVOB+ExoDggWq8Db/IM4dyx6TQM3v2n6fjQfPVGtYnCwQWZkGL3sy8X
Fmzp0VKkImxcZ2yEFK0Ezit2sFT35c9zEzeXEjvAXKMSg22YJkzRGfni/qHgKd/I
5phS52tTsR5+y8hJMl6Vzj34ZOmXqZjZtcKVciNaWhODhrz0RD8RGlOkHN8gnUmn
ED0NyM9CBx7r4OhL8qwgrL6hCOhRr2h+R8DxOu8u9mRhn9oPFRJ8OyDhGf0SqGtM
YEFAitqYH/mN0rMnxvI7EJFObcur/h4WOWxiXb7m22WgPrsG52jo7NhqGKOGRvRV
sVHJwyYB5BG9VhZ63NoNUzQxFYNIoM1fvmYRnxvaalqKKIR6zgRGKuGhkJ+ngGdz
BGSbB2A4HmmMYepdwGWPUQMnylNNDWp3D9NwClci+98VmUTU8BPIVZyHOF88Gxc8
fcXgHTC45vDswvwA/WhBwFjy+X9efItoY4tGyEGUSky7HDP3G47iNNMwPx1fJVEK
Ob2ASpOZ5roSsC85+NGS9imez9Wr/ZLrWZPuJsjQ7eak/w4bYb+OS8fr9Myge2sY
Xx5DWtUMcSJJNaf95Mu47urbcBlyskSNGE6Sw/yNfLo77hTh2zlB6Covqc1q6chT
qAWHtSt7y0lsyZ6UMpTgR6voAAYe4SpMOIamHfhzhPD1FavjMYNXBkx6T0RvCcnp
EEIEQMGfXADw2Gb8eoV+LkmHbjsqlFfPKjqBEiucoE14sG2RIKxldSNrLiIXyjUy
tU8szkICYZRqXuGvbeURLGULNbMqgtas4Kis5T3AbmY0Q92xDQD0V52qyGErB0Ke
jeQTUVvSmgb2E+oJ2+us/lb9Rbf/K+iqfxYT0iMAdv7OS3EvxHYGS9PmYDXdSoSV
wtJHlt09TK4OXJUEKYRoXJQfXrvRO2oIXecXwLZGcMehmxpH89eL5HCCe/Adbkt9
KKebVtLrea6ZCTAK5xii0uJ23hjcJHuYc6G+lOPq4NfIPWX3EUnyI1EMKaaw67R0
c4pIQX7YUztjtZYXWtHKTQ5fFMIkg+IVwSVRIlK3nsyzfes9LEms09ofdfdqNMiy
m2j2eBwh5Fii5dF49eGxFUPVH9l8x2c8bzTeCOKMYjLTxqH/nH7ZzpfC3EuUxRe7
g5K2LNucXLMy43ccMa2skGREH/9UO0ovmjO0gfbjHYUCWrsLkz0YtZbGaQYWW7sD
5xNiAL1fLBHXBXQgnEyzzMj5B6FVupDLf0sRWll7criOHhnrvbiT5FCi+WeDTOXC
H3V6mWagphVQhCxSF6NkU+6vyxiKG1v2qsI4Zp96Pzm52wfIxHJ4a48s+Epk/LvH
OVEwzlPOnCzeED4l3vRVfQq9LT7GDlR4/5OZ+yngNWTf3k3wK071erFvsOpX5D0q
+ueOK131mcFrI+89O49HROGSLSP9W+EwwmWFj9/iRm47O/UALA787c40MruP/auy
bCfhx1GAQXzBB8VMqRtSt9K3Zr3LEo9SVw4pJG7b0WWcZFJo/BljSKkJoK4XZhDp
tKKa/0T8IDzCGj9qh86+dRt01aMdK5Trg5WGVrWypQINjZ7XE6z2WKsT6YX2FLCq
eaiQxKL3i53Kzr/fCcJzxuv72nC5HX/m48UZA46t6EmaakSK36SftW8g0vKFjvr/
V3colg8DZ2auTkkAfIw31LQetcQ+fh3iWZG0JTreobvc94NKv1YCVEngvihDfMsC
uL8i3kS0Xu473UQS56CkRDvqYnm8XUJR2UhuOgsKvPdYqXT66WjL6SCpaPXQ1Zcp
gf9ws/x5oi7ihIaAlWtsofYCslycLTekGENbH8szJ0TMG21Ss2WILHpz6br/zEmi
6ZqrVxmZWkO8FNaRrZKOBZ4ynJxklvL3ZGeu6y19w0mfiphIJovYnV8mlDQZNtTn
gMfGrBVQpsE7MDhYJjQ7veJwOsNhuJ1txeahM5+86QfQgPKsA3giG8ZOIyS1QYgp
i1SyGCZGjjbJTQMiShjUnWlrhid5VuerRBRlCFtq0aaN3y7U2q0C1LyiiWCNW3BD
BHposdoQrt4KCRYDi4jK8Aavdqyx8e4Jj1WX/kijBYgZAIaCTxmSBpJBqzpdufo8
aa/pcTQbQfkT4GVTvQSVAiQhW+HCe/9uwB0jAPl8VTvyj7xomiFVmH2YkhafHAzZ
rYGORN+13XCUfYRZVDZr98c3/ILjiItBSczYCCGuAb6nHDLiTdqElb8V8BYEcXs6
UmF37/gJ73xhIBj51j3Jw4BTsghrEX0S6vtXR0ogYB0sRzhQ5BY7U1THVxFUogfU
Xg2X96nuI21bExPZ/aVi0JooNTDODGepGtezJQdTKBTsP5wQ8L8nMbfrlYLjvgbF
baJEs4SnUUuQkT14/W5muSYY6o+J/6mJMnUVC4oybo8SXDdf/hs6+fZTmq57JgNa
odTd7W7rMYp/N5nsHd6S7KELr7mnvOyDlBXlfX0bXajZNBjojL5Yneo1nHSxnKd+
ILcr4C/JHz5GDWbiQkdgv+4FYZXecrDKHdFhl25AawVzVLw+JGxh8T+CCBDHsEHP
C8qSLiveCmrC8eCag5/QJaIPmHccYFR7tvJinwGFeyyq9pGKkP/5l7vvu6fwmvt0
3CrZ9lzL6R8/xbQRYXn61R9lqO4JXNr2gIAGD2uerC5zuDY0QEy7WtMBmEO+KfqL
bxGhqPdtj9fMcYK+ctLOvjU4krZFZmHHNUCqUoM2uE/PEBZVix/+X5X6OTJ/YbYN
r8js7bj2Zr2Tot0p9JNKEl3nAhKkiwf2HurgI/y4+ez9JsbGkYZxrTyX9SRhckCA
ZWdzzVHGnqiTFrbr7Xaa7qZEu8AxR8o21+MHdUOHrhqvoGynjtegguPhaZ9w1gD9
m0TGpgBqSiAZk55fiJ+5cVmjjjT9ebo3yx5LzPKQXPA/3VgKmHHq/pIR2OhxXQ1/
QIOuo00hK3MU8/ShBWN9WJLRfvAsVPeQYfpBdaSKgUyGYkKuGfjBBvtC4cSGnDUk
AxlUb4E+Oq4dYy+RLot7F3RK6IbT/qdpwOIv7HqIrH6+rHpKtBJZUWcc+U4Cet4j
pn3n1ISz1Tj/si8ZootGugbE+fPL/WzWyzYM6F6L7Wl7ifysq/Cc9BReT04iH4J7
WF8YZyiYScbIfKBtNuWq4Vw4isWDdz1NFSGIr3S7uOuS47iJLSz9t24Mc5b4MvWn
ymcUyTpcbIsZuE60bnO+iQJmL+IMpoq5MStLzKPwvtYczmzRU9GnS2PAINV3KCAX
0jcT7u4R8/BZF18tY+3Hsms2FbDKkYfoefl3GDAIsLQKRa1BAaXDpZse2GZGWxJb
ioVQayXdrzCtHRLWN4kOPIsoti4Cs3JY4CzsukTIBFTvQR7/ln+eejQP+gqUUfo8
FE14PzfBDPNa3b0NSOS76izHUvZDq0tLTU22I0JN3iymPh3en5j4RtEECEsMIqda
sTJJxaTDFRmnRsOgS9conzASqg35gYRSqdwOwAVxiDMJxvHGgbcfCvbD0djoNz4E
lBAxCWx3qdGVu05MS8MUbEb7qncRyDGuPmJgfcjWlVMe1a029p3K1MGaXpOZ9zA4
qUH4aeayebG6v2IJn7zk32y+JK1c4jiWyvzVPTm+8wsLLGwYrnadNzYnSqi0HYT3
brAW4YUTb1FyoBUCnP9iIaRSchy18uYPPZneCaFn6uJSm542Rvq22fGXiXqIQGEE
crKB1DFNKChlQWvrN57RbJiQnasOVEqTm1ZxUrqKJ+x1wra7gBbkMDVPqcqWJsNq
3r23v+nsSaz+Rk7MRnEax/h4cyO2b4OoT6brtn20dy6pM+iEUprvlzxLSOlGAhxW
zXhY49xHuESIhj1qp1i6x0R5ojD/xbzLCigYPfIoE1b1Hfi43i7mjIhqgthAsxwN
t9/inP2ksU9sO5ylfCHegz2I15xQXqMtaEVdZ9oyQQJz9bXk2HryseAWsUu+bSW8
KSbR2b7AJQ19eCz0B0I3PYgi65gSuhGrO7+rqVhNDYsvbsmPKqZ8Ii2fz7lNcdyb
8N/7/iW94xNqjNnKHA/I2VbSOTokUz2KVOwSQctjWaRan0O1BaDn93aOfaIg9rpZ
jl/2+OyKUVUT07D5DBh+F29rUltkrFoo9DJG3+TV6Jeo2KVDPiYkMd6UXTH/7eWV
63kUk8SuUmdoUUfQunqnOXdR4CJCc1HAny8p0c8jdw7hOmJUGxpkc2JGKIObtfyI
Liihgf+OAKP1vMc+g4oMs3xNjMUK6HOxWcMCjvEO+7a6mUgWqrYfRu4nO+Kpk8eg
ihul474R94zR1JIT4pFwIsDsmRj1p1a/d0uLVg+IADLARPkV2soEiXTPvj5dKqfM
mz2nKRPzU8njlhsALZ5q6KRnRFGnltkngMXze9s/hJ8IOqnUzR23yZv9m5yru8ke
Vcw78m1HYxeKRfbd5gyu6u6ee1OII93RsTr2+kBOQ0Q9zc1lwCWUN+/QuNvXIgUG
fMRxOWbDEQl1L/ZCZloNbHdqP/4/nY1cGFWB3h13BtBrG/jZzaIXTjHObB7eHW+q
Zbhh3dK7ryRsPRTbQ1dl7IVIh3C3TdXoVLcII0iSN86e2iVEMnI6LnhPRipwimk5
bGcqcKD9GWR7SbY3rTcZieAlm3J5ROC+Uohlqs91zC1L28Hwuxg6KHUaq8RgT4dV
rzTHBRavCFLChMTuYbXiOsgkMZjjaT47cwZ/FhHzJLR060SUDSitFegk0HEnCeII
Gw66N1nijY6aLE68Tg8j2WbPF638oPUQdfwUmhi5K/vUG2JK1Exz0TOblPO8mkda
weO0N3IhFk5PVNRJfnoz7mHIcAlJmpDeaNbGO88tuqNuVMUCtXC9qL+PW4AqpVzU
rFm9D09PhXpLjiiR5jAw9FYYiC9rmUkx2Oeido4dXUX54HoK0UUqYCMnqFGrfvHI
d6GS/X0oTjCJkd0Pt2hJ+qdap52V6SrqGKtF0YGguKZ6EYQ4d74GB2n1XVyM1O1s
iaUssYMb5p3nsQliRpvrCUEaVqJ4QcUO0Bb7Dm3F6Yt67/Dd+C9C3gsnLomi1A57
EfNyqRiSVavFFf93zcvwWYO2g9au7PkofLrFhx8b+LhjL6vYEkHwtKo1NfDyd/xM
/Vs7tGuj6OURUfEooyRYN4yVFP0uuKgSPUATBkJPzhGCKADECSoBLPqRxMLQKDSi
h2XUZHztCmK4nwyxoV+UHTZvti+X1lXTYPW5MO2twC7uDZwdpUe4zpuArk6gL8Qu
Xpg8oeBtBy3KaPlYe7x9dVnkQTsHt40D0fXRhTffj7hr27zCo7RhRtgL90EqAuzF
/jN9PA0Qdcsc5clZDOJy12D8LcLGaJgr3rvaG3Pt85WHBUCFmoRejsFkKtEtDXgS
uap0obu73haOrkEt9f7VfTUiJlGdv+HkmVlGTmPK3tIzr5pQDqdCxy8tzw8yDLOn
3iDTWRZjiTmfNoB41xzbfeUsvBPmW6RuPFvnnH80WpOYuwLJIb4Jm/SLKcnJX0MS
pDaeYCoS1vNycaah3SYEjCaY7oAbAyYMCiMY1m1NFHYIUto76tCkJgf6UPpD77C/
cIXD6xtYBjY6tCR4PJnTQpQPMS8djPE9qDklBjXbSF0Vz0tj4dnjdQAqguRMchIw
QGkySquZ7TuTVFt5vLLdjLcAqXEQ/oyWclaWsy/yLdQJHzwTjy1dEPOytGrsh8RT
vYHqpR2xYoUmzL1PpQARjVimzt0uTK01sUKh5MI+8o7nent3J9DwhWJG494d8QzU
ONepg/JDEfIR9mawmKP5k/Cl154pvCC6iHOqsicqPZuWIquO03HB5m44SjFd1IkR
iyGCCQdUQAXaegXNapTlVIUqid8/qvo0L/Z1Y8agcQpXyI2956E9/gCJ8+K7Lvz7
rOfnw4KvASJGlvJ3uuMoVvXz4mA53l/bI1eFC8wYe6LGJi5XJ3GWMFEQ65Oksk3N
6h+nJUAude+nZwNGew2p+JJ9sXWeburwXGUkAfmQNonWShkuZppJ36i7ueTCTsFd
nGmopVh0Hbrdk2rNpvAa/T51Lemdd0AyC4bKtJLSqupi9tlVDnLk0D2pryk2Q3et
jtJOadZT9CGgPGnXm0VKW+/HwrVeNhQ8GzTQOoPg/ZW/H9hACO9Du/q6I2Voh45Q
svbGAZ8XY7BopzR8SwgK67Kv6VA2Y4oDXJ9fJy35mMi9fsrMDy/Enh7QWY43Z7RT
TwyVZ8dTovH240wGo9UqkV/zGTiJVSvEE67BQWnaYy3P87PESANVyPbRo82grMc9
Tshe3MMrYEdvihrW5yHp4fK4WpYRSB5tYf9nUNRwpoIIDxZdaWOD7ofi6eGvJ6Un
POXpMOqEFbnX03InDXSWS2ST1pbpCqKYfPt1VYwj4GcvhepbioZIUhyaII84T1Gb
iuIonTN0BSrfiNzz+A8KwJQsgxn3zPigB2Tsh/QoECEz9RXUuE28FJxQuirhktky
ZXAnUxyLM4NiEmfIPpcsNvcotDJOXdmdw9BF3Rv0hFmIaBmre7Y5oXFVopoiN3ti
59DOBlo6LWYX8LRlZDFkzkAEPIv6kYkFHtS7WEh+1ntDcC4d+onMc1Yqzimfv3jY
MC/6PSf8ds45S/nS8ihNLJXC6KZr1tEA5s5Ako6dm6AXsCXezyQscnFTOudOt9th
eFVXUAZ4i2Cr6aAsw82xtSgcoaIMc7VRzov1ND0qJXs3awqkogh3EJNn2rANANvc
lVIstyaQ2j3AdQnU0AO4mj8RIQ8qvJQMzTl/NBoQEl+9VaoaEZM+i3yJXB1PCXiy
S/yV4xg8RbeNlM/5Eoe4QJtgpiz3hDGJYUHu7qbe6am3Qq6FhRX4J6IoCqBjkusT
smEED3mwzo8crSxIQriH+WXged9TMTnpy8CsOntT5B4fL4/tWCgwHQn6b+binBdJ
jgdGojEcTme3zsWZUSBRglj2bDEegcvatlvmMBFVdxZ61XBEjd/9NxY/Wljqu6gm
36mdomYL7TEsktoan0yFRiIu1fVkZv2D7nWK4IuvGzznBNuqp2cJTj10T8c4bu/W
sTFy/zellxmIp8ugHlk2VFZTv8AMF73W/k09i2BJjA9ZdCxLXDZ1zdI5U7emzJKd
mxBGamGx7qtsYaVYb1Cf8dlSm4J+hsk71MjfrxvqSCOoAZYHACf/8MlnoN2+6Muw
9azQgHx63+wh9ss1HvtMuYsGehQ0fp3gIvJggb1AWf8r7FTlpswXIZLAaG+bJp3T
TiTvieGfStA8GnqX66rbYzsiZ4IE0uBLRKuKy80DSfGDec+Pws8vxlHo7VNz3TUv
xTgcQNb/39o+WcdQRMxGM3H4C7E2JFcDu2ZyP7cqw0zMk5vlJHlM5zxXMNK6LyFy
NhrVtqprUAmqsAZ4O4yfEyMr7FlrJVEdvZBvyOpbZY4D4HtMAcGpu48vlpI9zcHu
wJacKPJwfNUMNeVVVRO73xdSXYpBwG4CSDphPs/efjUi5UsNrxGwwuI1k+5uBRdE
4xKkDU6LXZey6MJbMDze5+4E6FFVvi0deiBXZfP2uIIUrraNk2LytJu7ibJf/rex
j0S01atBBKguUNvvqG953iOK8D+SbegeWGLo9otq3bSEaeuU0YLqwegEIs0YJsrO
EJ66llaHMYTZeA32dxfDswDS4E1a3QgYAS25sUK6U3lHqr5kHIMVnAWljGi0ZSaF
K7fxyYnho17Sgjq8RshhMipHAvUyx+0QilJqRJDulIwNKxATn4L/5U1UhgBpSwAw
LjHOaL1rMhu3cQoHxb/UsYZIfA4UsP2Iv6yGovEP73QTWdjeO4JAJGTW4rCRg6t2
4M2ih4PVyXmKCdjz0K4e/z+euT/MVn5j/QXD3KViOBDlK1iDiYaeuqM/MsxK4AhB
PA7MgD3xe+h3z47QdEuegojaBdexKdisae1DTt7UmIbU8kmHxTZ96eZiKX1p2f9i
8cFxCEa8kaCh05fhDFTqyuNsouYI3qykJ9Vu5JLi6nPliSrBx+Wwat2zAKePEvj9
gPl3U89Ijrdyfibye0FvSiMt6dPqqiFBztNzWWxPtFewn2nrj/ZwLfNkFg6Z9LV1
Wt+av2eGo3+/EXOzC8IiVj8S/al3ifPz/mEDgEZLdrpthmWPPQXt+Jqp8ZBwpPFg
vz5dS6+wiVIy5Ww235yoIImhNBRSCDehoVLbmCqakcoCHEmI9YFT70A8sok7xWxS
2bH7rzZtSOjJdD+indrTi/N75j+8ve2mkTAXA0twL7boABm+8NUXT3lYkCKtp2/C
AS0vbn7Un2Y7/BUbK6JC5bMgX43SIaYFOAOgiQFc5p8DrFFMN6/2v1YwVmRQTERj
c5k4LXnOz6xNqk/5L0GB+LRc1Q5plp252qskWMXO0hoXbHSOOeq22xR5TK8lKHj8
oACPUrJvSD2IdtAi2DMl7ZKr0yMkOpQIeWwWOcbpbSIRGyxCRM5vFqUjl59zUNJC
EnfDsehLIXH5CnTE3X5ioklYLMKLh/A+DBpQcjHOEyQP3FIeEy1F6jJDf0OFEhHz
xV2RSUQ24ldi3pBmOsBhM1dQp06phK1uCHxRowbSyfMyudm62Qf98D3RbYZ5eB5B
XE/GCALKjGhUt+ysF/SBwryoq0hEFiSL3tpZaFakarsYOzdRtXg/Se+Kv40UBm4I
U5oUuTElOH0ZOPyc4It6LIGKF13GUgiSRPSnn52ElrHqgCRIIxvDVg+NEJ6ZWJ8G
Ae1U3ST4nNUirqLYfI/M37+iHwkSp+kloULkhiMb46oLxdE+LXTR3jq3uFZn0RAC
olUoHUPuPm0xdq8O2z/pFPGSCezbdvM9w5r5N0AJgSwKpzdOBg0l6bIJsQzJWCuk
YtcVGpx+xTIialRfy29IRkIByabnYc6OIjVr3BZuMPRj+vmREG1cp8Ek7r7IQ6Dm
Pte0kaHrWdd1ruQM1v7W3IcLX+W/EVXzhs3rEoWaUdNqqiHVe9qajL0ApefiEz+l
cL8k3zLFjaR4YXnog9IgseprmyuJW8dnPPm7k2dobKikUI/HMY6+5nEqp1gsARV1
z5GnmLJZIN9rqEbQZYiKU6jABLO4IJFaYoiafzCCF1CJ4Xg74FKKCs7KbPiuNYgd
1qI0PIJmJd4GdT9btUzbzL8Y8Bfd4OL7AVHXxlZwLAxoXQWM7SkIAVWuMJo6TZq2
Kpq7dtCsD/dqYamDbDwL3RQ9S45w0TvUsUxUqr8anNWsrVOgp995i0Gag1Hif0Tq
X+qYpx6R6NuBFeSYcC+dEEZcy/hQJcCDqlX6Z4EFvlqx67rdsvWBVr02njL1/IW8
81rnyMD3Yor2lq7JsSu7UcgczMlnicMQiD9tG4mKgFHEU/cTrVXoDSF3OiWt/pwS
r3AplRzxv0h67/jYFSyMLB3k+0RdTyiQG5dNVLvQaeZqk4u9RWN/tCNpxBt4yh3g
HGR4BxCz0sdsUwmuSWUJ7YIxMw3aDTMz98eCSBIJEN5cwm076rZccY8cr9H5QHcE
qzGC+08NgxrYk+hjceyQiRmSPkxiWuV8xPOHYlYdaQIM7aZ9NGqvL/c0H4r2/AGq
dckgZMuopJ/XoeI13/Nn5jQ8qv6RIs5RULiD+WR92OcDSIjNWBn6PE8yGbBJogqr
FXa+fr19lGKntxYny6Jk3ZTsu5ejSGIkus8oWDZ9lbQpcfK9ajbXUoVy5O7/jU7d
IA6sSoEYS/hX+5WjPJcgAYgapLmtOdcrpMpEuwExlTfxKp/WpZS5eMcAp9wXA0k3
KnYClgLHuADIWhsvtvG9VyQDWzdc9qzrT6vOW0Ed2aGZOdKMyzKdKsK6w4UweTnz
VfaQMoVcu8x3oQjI/fXeEnWjRyqThQmu34u0JlamdDyLP0zvkFV6L3Y4P78kOkDo
QoN/ypJ5abFXDESRDqUFuNDzq3kbrt29l/9TnJotvg1vWSyd+Zt9a26UIqhxZWZ3
sMC15VZl/mGu8B8wif10q9ti0CMnl1Jc1dG6g0YHuyLajTvokvcT7X7e3Lx6Yycm
Qh+bykyUcrkLa1ePxZiw3mirkwLWlMmAFXKkN0Y+1VEBHnx3pdcAtRQtUwg/QndX
L9MYEunM1HFixLQv43JsZVvR8Tyk3n32/S0Kz1WEQ8uKXv00EB+B3yU4HQVb8FlJ
GhFi5nHs8tpwnY5Esq0Q8JWg7gvqfeZBzfdJcfm7mZ7a/K7JqzSkiMU5kpJKEwWC
3T8wouhl/LNk+PIDu5Ve9Xg6TKnKJ8jLtl/9+1VLjpWGimuiasv/3K9yoYhIdfLJ
oMOPqWFUvV+1PkmiixuuO/Tlg/1d87FkkpfgQazBhKXzi24nP/TSIQjbgC+tD+X/
CHufQosghEozquLvvrxMVAxzrYnGjUEy3e4PqxfqNRyeebATEpZhRIrR3xkBq2eH
80CyitlID58PwNmNOucQDyrKBrc1Ej52bFDdlUIjNNSmD6N9r7a0ciLb/Tl36DCp
5UnChVng+utOpPpSREaxP3NBdLdmm26M6jnPjeHTJGhWtuihnLcTxm8cVDJUstq6
2sOOsx8IBYU7mAY5Bi1ig7F+pSQIbq7ZAb+y+4lwpzFFN5+ieHGiqJ0m1DJ+a3Nm
X2PNItNiBIZq7V7/oeQJLEhjIemu7jSFvoOr7zxFLo28QY6jnpNdaKZxp0yntfUx
hkONo2/b++z5Uy9HWtK4Mubr0GKOcGdTJ5XK+qImFShNxODoUOiE7/0+LGwSisTL
sJ1AQoOlV5/J77GRGgCeyn1V3FJWFze+EVG3/FnrIUsYWF4fll522EXY0prdFI5w
M3EiWfAYXaiaFirnXXidZVTeiY4D3V77Ry3Nlmj5CV0Zwi9cFxm2QwTijWokZvge
1MuDZtBqGOtBp0raAEZIwinh+f0HeMuMKo7pCQ6U3vNBdWUYAY5MvOOIrU+jJIqa
zIOj0fGJg5OzaXavKs12Ohl1kAHbo0uTxlDN8Vtqx1tLQD9seq7KmtO2fiU4U5Bu
mEsRBFPiZx7GA94Cw3LtvHFhab8rSFZDsOWrNdSoUia5xYdISYWPS0wPhnrEio9L
ApPnEzlb0HT0YhZSutE94DxcQWZ2EUTnoBi6EsTl3UbYCPAJrnrCE2YUgWEEaI60
w/GcF1FH7WDillB7sVueAc6zPI6ZrSevR5xfGgET2b5xaXKxzqSExrYYbPjS+ao9
tyHK0y2zf7Vo6b4W7R++iy1Nay50TJL2LZIFt49wIjeptlzGPlPUc1tDFySUuT4B
YjeDdw8cR+dGJYG03SC2rLzi9xzjJAErVT4XEyOuLr05h7uNenZZz8olTmRL0s1R
PkWT/yXcjtl1NTuPjHi7cJeJAnSiHYHTn7yV4yVHScdYicTabRHDVRn0aUbVWK7i
Doq6QpzarU+s8u+OuHxki88bvfFzUgMGJBHi8FeI1Gy7Urzaw7EORTijCh4c/Apj
ND21R36qZelNn7e/fWU+smXCKCZSR0RZtFVM12vVaqZDLq1aDaXqoZw+d52frcXL
yZHX3SWUQFpE/1G1joF/i/eH8jkUAGvEz9/AZbX2NayjWIipSpAoXy3dFJOdZBMX
yNcG1ZAQqu1HGMUmKN1V8wSnLNfTLq05AScZhuQc6LPEsABd+wzdcN4JXxZrnG0N
MysGQjUwjHgD4x/bmncmlPWv3EBVntZVQR1HaZ+E//+KjSQOPSuDfLNd/+uqvuhS
4/XYF82rcsV/fXRafa/h4spOd/Tu/MsFTtLdfm6J8nM73pWwLeWd2l0NqdjSDKdl
uimZsUJyp5rYj5HMx6Ho2fmHcWgFBqe7PeMMHauVpxMn+0T838h5EMcUlS3AGA/H
QgwHUEJGdbn69GEv/iVyU4x+6cTZcABRdmyDuklMXqnsTUpmiXyl5Yt+EPCaJfLo
Dm59l8ZGwy8AERLUcC42DraqXqDHAyJeIIuRd888GrcJluZOKmx0dq17tVHwaA16
+lUffE/0h23XqeTdFvvqwJNGom5OQ1fy6ZbZa1D6YXw9TpgRvLDmZLiQunbHdtCj
L28m9XW+x2kLHeXST8xNJHOYmF/GtalNJ0luaJ47lGCKMySwaGsY2qWI6Y32ClnF
iNyNtQh9CR8y0qqj8i44DB3taZeAR+Wb0IT5tb645mmZwegBB2ZpoqQjIwIvIfjT
uMMym/l7cnPD4kJej1YJC03rZBOyJwsvCPrEOchcONfrCyMKHYXag6XNuHp21F7Z
cz17bTphpqkY1eion904U7Z3URH4pnkWFW0ynCshQDfeDE5QU7r4Fyr81RqKVwDa
b+DmM3B3iBVUHugaHQPbm1aXEGevOd9Lu+A8qABmT3YrbqCbUXmqyBpp0ZTe7C0a
E9OsAHRIY45r3qoXxkM/jIOR73hRcMHzg25stfy282FTk5ZZMHqrPEbVtAbp5h3H
5MMCSCxRFvZK79uPO4MLf8OkGRujHioZ2j/a0j8yRzHTpa0Xu9D2CaKCDWoaNpWq
YRLzcgRULnWMhx7MSmUyqbydrM7kakDXJbDaNNhZPxaAfZWVLloB2ReOKlurJsQW
HnbhJAvQYi2LPmdJIYrAN/hBd1PHxjswMsueHVvHLZNbyPlIoteEIyUg3IPf6bDw
EbqMOpYKufys7za3ubgCv9Dz4c8SH+dn5Yfxago8h4/WAq15tannRgR1Kf5vBUBs
2PDI9dSg3v1rYWAGpKWIkTM45XbShHu3LCcsCJPOb1XcmuwTb28W5isXShNyxnuD
22SMbrUuyDMq3QYVCFD+O4Z2K3ak8r3vXYCIAhIbE5nWTrYyN0odbUbtQNHQsz04
fOHVkk4jNgjwxGFHaBkw/cmSALVDhLha9Cc1PKk7FaIDYxmT6Ffgj0i7z7uCca2x
Dy4ZBTrw1VMlM2RcALbtI31pmcMo0pyUT7yMIo6hXSa8fqWFGj8QiFp8ldWRkOoz
N35wnQfNT1/Xt6iropCgWSJ/qS9yUwA3X9ktiDfdIkcfNvPZZV+ub2N8I597THre
A2kPp/ssM70VHGpNn8lTxsYXOMqfVakNzP+E9nAH8czVV4h0tWKyAncgriUnCIvi
kjh0aebtRR4sjeGgGxCS8RtXjHiXwQ7OoWB72OAwMUj0XpeRaQEjWO3WGfGfOd+a
EHAhGZ7l5nuZ546UQyrH32vKGQDCaE9lgubL1Vpj44T644l3obp60XqhNuB4jkSs
m3/8brGuOWzkXP6RVh3Eu4XQ4FVQL3rqbOFmrNddDfwsZHkK8TjvfpgVa5/bi+ak
nP3RN1qBmuRmU09GRSqPUO21ifFUKjYymsuABfjnQdb6tctdApf3IGX5XenpOXcA
A/DJ69Eho42OBmRtrfnJzwpygKP1HkjePGEUoXQj75uJNQdTSmUkzQ+qsrCG3/q1
4x2I+SeCYhlPAWK1N4siousbESqntsa/1S1Wsa3uQrWpnVZ+bMDSZRoeLkr3w5R/
rPSHvM/6Djc34rJO63nCLSp85Zx+r8IPOdg7JTpql4sCkDmVkN6wi/WYcOoTNY6j
YUZ/ByIaBzRHZXpHAOyyvCShVVq4O49G46ZTK4L/6OznkTHdmitmKmeSkYAbdLo4
NOvZCCky70CETm6wvPJb7S7WjUjsPPR9fCXD9TRpD2SWy8PNiuYuyvIq20tv0lZC
NN3bUIAxukdT/DqEe7eM/5920IaXUOprpErOJI9qmXYS68qFLW5quyuTQStCJhT0
qN3fXGv1Bd2fZ7wRcesfbdIEuOZ6OS/8cDUFRsnqibG3awUxsta53MGfWOPhdjQB
yPaLS92QNGan5rLHl/ODuxIAhvi/1VG8b9A/pXmntDtqkBXiOZLlUri1DPnbVq/F
qIeyT7OvoeHmzZRWcBLVpNlHCDYjoXl9TCr8DcKp2+e3xOCsZV20wmruLWoXVIJk
s9bsijXn3utDMSMkHNwpMacU1zd0BwnZkpKkpngBZ2S7NrqWXJVuEkfenBzaRQe1
4y03reLO12aZDT04Ckd50QDF6W6S/88po1pPwhjBerVokcPHDmPF0mWFUYRIRLbm
7pEeV3+eZFFHgShtwNpFLsMVGGbvpVn4hNWk7eohXYNPmMiCdMF67UrF+Yx8fWZd
1Wjsp8Nm4OsgNzg0bwHUvTTioo3sMNAY/aP/nPx69tpUHIR5n1SwMtSXWLEjK4wh
8zscT75lqa2ItO6nH9q7iJDMrLialUmpe4wRNyaTRy2VDMCLIaNMiYGfAEQYNyxY
pKYwnJfD92R6kmgPJ6Zu43a+pvrnQP3o3RrHwWmflUiyNRai+vfQLeuCR2YIa+qi
7jN72hLwkE5yrdVyo4+CnSIV3XxzoZ+J1eRVKAbp4/EuS8j9IIErvzwy6PPYwzKp
bb1h1Rln1Lb8ENRDfd7NwjY6O/8Fe4lmiMlfOOGwIm6KA5vEd9uVUzBhs+vHExAh
0d/AP+HpcN0bqalfsj+Wv8pIC/fRRhbUp9LoxRdQMKSoRMrrUNIRWePPHT3vtKx5
OZHB17+CnSIfd0z9VuOWKdfNj8TKVuTGFAPcEAg5yUieF0md9vlUA8hsBZXNsWtI
3WIbOQYpBBIMNTohCl/IoZmEAvVBC4lVzoNZ18Iy80e4N+B6CGmB0g8ileYC3yyx
KIG1atk7xTEhO9WozJONXYE0q0Qy5ahuRsne3Ry+D9GqQy1UGMOzWBuDLsAifRAT
w+9cvLJ5c5Tl+q6M0ap5Af+ZW4YL9vSoM3qbeGARl0BEubRKCISLhc1g/CeiRU+8
lvHEHOFLwDPKdNjDIXx5YR+pRojUVsbkYVd0TgWeA7RIkj8/NzX+q7gvwOoaW/uU
gEMH2DIPDNbNPNzEzQ6E6QI2KqxLe8ly/clgh1jn/O5N/LWGSvN/+XGEosAL5lWc
R4JeXddpvMLnO1VjusYAHUOcCe9wquPTOi6Vw9XQtwA58+YLIMxmbQxFPgGTbz4G
ab0udM/fIfwUcQZaV7DbBmQ1s5H+gF+8T/4gjO3fk3KWQyXWIUjYATcMzijSQ3ew
3ghS/wx7m+md035Vwd0dv87KaOaORblu2c46sLGJsAvVM+LQV7rukxB3EUdb+T8F
RLbS2y6zRSYgOXFRK1SGrRbKvJqMy858S6fImHiU0iViLmEK509/sNvQHlxJTojp
xZ6mHHTWn66b88cgU/RcexY/9vHI9Nc2MLSH7HV2nKlKmJtlB0+7dcpfSvwHUuaT
je/Fyi7Q+Ybnv/FFXY006ox3pSDtwnXUzacgbZq/ukxlqTFVG32b9BJg6CrmEJL/
nh9IlGs8uoY5EOlxds+3kkbCSlKCyEomjfauHBm/TTbmt99DY88O1BTUjHrtjcyH
/dhoDHkCO+KL/Er6bCNarkEUFQHr0QIC+bN1EZrKSprEkUo36lCxSMFiH8QEoMMJ
11l9e/yRgEom8y1uyTqRIkbMPow5q6vOblviOb/2jQpri90PkSrrAmc/h+W12wl6
aoiZ8k5MCLoC6DMvG4wcf0dV5sLfJ/n+RqXSV2LMh/PHcjh+Vy5griANqFZSYpcz
5ipxdJn/SASzK1sLFNJf/+LE9Y8IGJWTrVUAkkz88ciwU+9BPL+Ut4QU4dSa+bvq
f3s3bi9jgPXBT8gYpwOCO+f7mNRcqLCOyixAIzzC/SFpsF2x6v4iSTwEaRDGZ8dy
XKh9VXG/DhRJwZlQBq4ueKGqRt+Imh0eF7JHDfh7qb0ak3YaLn9Ha+hUMMKInvn5
NAjnGgkmsQzhzlgIporwzKLJL5SQBMNi3bqqpb/gOGiJ0r42LhwzH9fYnz0Nib8m
E7szmfVT21wIkj/R4WTtcj+sfgspIypy8OdA9DRF/mR0kwR6IcgAz7z5C5IN4OSi
uhJSQhTkl6BUHOJlNcZ4ZzHyJPgTDjf1aEWxD7THd8miyeMndZO6f01cOSBGbAc6
1z0mT7Ubpct9XqilCwRRFh/QbE5/9cMOKpVF47L1/nZNZcPNEEoJ3jj+L8408A9V
fN4lBLoJGmBjUAIaIVxTkjyUBflR4Emvv4pexP8vSk229CryCWi+hhG6ZJ9hS/mF
yJ24TzN8WucZrPYLovKUXxlvmlNqzEKRqac5u0Tw/mlCv+l2mill1IpB+WmTLCqn
CAlECkPb+azjpD0KOxQxsuYBBszFTuh5815LWdGtOho398aX7kAb3tnwTxVL9Jog
ChsrcIi2pbudU3UUes4+8wfk346d8A12S0Ak+p10yc61+B8Z5pxlmmkvO5uixkoA
Dc0uFKwB/e8QDR8sUyaHck2rxUTokqCDTCFYyIN15D1HZbDvraJIq+PArmv8yzr5
muclrjeW6rpXJQbXD+8HCoYllYUsd7qWCfLY5G6WMjDfNNQqWCxFFnUPal9bob5Q
U9SGMRmWM/EYmK1zRoHUcKgYnin4chYSzjVjsmlBgb+usfZtSQ8HsSn/nd3gm3aK
ZL+vR/MeeOUDTupaJT/Az/vdhOu1LhepFawak3IFdUdQII96TLRYGQmyQs0neW9a
GlFly1Y1meNbJRDXl0gybhtGbMOEXKUk/IfM3hqAItjA10tLdptJb9acILufcMbk
OZ6eEjdrAjz65ZpDPk89/1rqcGbsKVA65qWdd0XbsXpdtG6pEC6/SFG6gr7BSa0S
EsHRcFVMroXmqBoYGLQXinpuZamsoxy1RDZfTryx1T4lH75FyEpW+oqJn9Ly9+Cy
bXYXIWsYGthu1FKpO9j5hI8sJ9B8dp9hybYG5++js2nIoUQn4Z27xfFN+N/TQKPO
29yiGBR8qWe4ykPgTftOyjF+3gdEmvjAzNWezUgnBA/LXnA2CUppHL1xPcCIq1zB
MQ8mwoedyQDSnuB/OcK/nFC09R85KsPJPaVrh975GrwyXSGcPpMqNK9Zc/eebYB5
QyCxK47dbA3QwUclXTZDVtgpxZnP73C3ZEL6ds9mkLuN25x/cYZOe+eXy1AbvNfF
RD1sOus3R9tEVYdRS27Z9PKW8nvfEsXlzODLwovO3j+U2e1iXFkVyYrenG3Am76x
c9Tju4NR6alVqW5K+xkdhXkYgjSI0Ow4FLmCqlSSrbUjIXokpDcug3DjcDjIME6H
y98lohmyRiqHMHzU3gvc4ZTAO90+Ut/KsWpDCyR3lQ688Cm4y8RgiIDw42PbZZWt
7oeUtZjkroExu5Zncs88XQ0BJNYnpgbJX2QoB+f8L1YY4KKD3F2GkpZqgB8UGqjH
8J+OFVtZjq8LKg00TzaoONRuBSHdpviMNcM4Z+MR7DpfzcVDc6e+qCleOvPu9KFU
LPLCmDe8aYhrJLDiLMCaukQnYR8U2j9D/snDdfad11egwVYWMTY0nsebWBU7LqET
dXAotIc427oZp3UjzuF1afzkVvcVZCa7UIN1myGJd/A14U9GNRd6lf033NAp0Waq
XZjZgpH1/U9IFSCyyfaacD9+/cpiLY/lkdQB7QHpU6Oh82Bu6hfQF0DATZViOL1W
lW7B99xN60NyX1bV6SjXjcdNhU+V0pWrTbVg0KIcFUWGx9ujATCBfJnE0le7MemH
bDYl9kkrHV+0HQmNZrfz5UGfawDYJeJuEY+D68YteWDYyprHLykkJn2ibeMNWp9M
2+C0KL+YnVnzHXJP0cmY0q3Em+/uQEXTeVuZjNU/Gu5F15gqLQcwCNyJbCRb5kgx
XXLDlKVI4AggOj6ZKGapfsQ4ftkU9szCTwfOgHea4oWGKIvPegW4lJ3xj2U6JrU9
6ZOaU9wkxkFrB3S3H3lvzYEjK1O7bQAPHuxKjoEeDSh0uEfUOxX/mGqkxJKySrBL
WJbPs82ukqzzJaU0+bh/utCVlcuA1OlCD9RGILnkSZcvXyO1yryKOiu3QTdFDFHU
CPw9804vYR6uZGosVzhY6a/ptvC3d3LLTFX55ivfoxCOkzTMiCsl0+exoL5oVMB2
R941h+4RvWh47sSgROXpMSIzzca9+ORHB/NqGytxW28UvfM2ckwEZ5NulM2uJk5v
u939A/9Cn8TZa1XJcGLSd1iwGhP1A/tqxdH5zVVDXICDT2vrFGdA1rMALnWyp/Es
fQK9diHkt6Ty8LDMk+uP+6TM4Xze8Z9NUh04bSnchvrMkybAG5CjAVQyxkl5Th4S
r9dk2b5fP8FgqtzTo7Cg/oH/wMHn4uX7iLj6dRJuGmNn61rjvgP33ftsvk/WOXOC
8uMfqlAv0ILqM2hxOaBV08w8U1gJzMpHyBB1xc2d6u5IoFzvoLi7tOq7SGDNNa61
6eArrORUPa4s/7Im0BnZ/RdTEXjXE40Q3kawnC2lRz6F+Mj8Qi9tYKNwGRhhuMHQ
HJJC7uAFK1YHNK1JTpG1iyCc2Vz4T4puWKhEku88mxPjZR7kj2VZ6dBgaxx81MTQ
j5AX9gMq20TjM4Hy/QHY+6omyOEyNPbeNGEki1kT9PKrVtKuFHwK4l7JooR2+EXp
2A+6xWVZED0mEBKo1iM/mkTMoHl9l5YXBMImZJwIYw3WFODnTXoHv+cPoD4hvUke
YNppYZOlXfrFNSR33e0+Vsp+qPxeD1qNZmYpLMQ/sTyt6Om7A++LxCCKoF+JFmjU
uffWbjMhmsi+vbO2WCHoDxqBaIJaf36zc4CTgITPV92aXelfSWTx0MMhQ2nuUg8U
yTxIofxq+/DrrayuyUYuemk/cnzjW5bUeC3ggYUEWwFWuaX2hI84ybb2VN4Uknjn
+H3swLc0qDkWBXc90bZenvPgLcrgk+3o3oGypp1ReBJw3eAV+WTRRwtDjoInkQ1c
YJzxNmEEwYij94B3VWDKGzwhuNh3BOicVBiCLS9NZ760xwYL6ICvAt+Wt/NfrGAc
aCRXyNsai6z8mc5zlsavNMjTTV9dnMAn6cBz/zwkP1L77e9oxZDl+x+yAfhdV5H4
hOgSBq07k4eB8Hvl17KlDrqECvv4A24ndHdtPWwq3wCyaP1110gQuHvHURxYMb9s
gpsbgKBmSdx8QD/zko+3/qAwIiW0+VWTFShI5ZhKRD+b9MeJ0JLC6/ieAgZbxTci
OlB6qHVZdauKr5/YC+wIofCsE8lEflw1ViqTQrCYlRavU3GQGstU3DnxnA73JhiX
HE4vDO5YGrP6Es4tBNbTdwpONtQ1M9L8FzJDoQcrgJFc+sRL2uSZTKafWVwKm6gG
OGww6tjCN3RGoyKc+4XQY4mohKEePTRBlDSPk1SoxRSCp6H/ACaw5ep88Iet9IwE
wsX8kZb4WSIHzH8dt50k8XTsFl6dlgvJNGGKAy52eMXO2/VjO2772yA+C91DNj1z
J5dAcbAcpJtsHqmGLLOq2OJsxowPFyGqDQfoKFfkExN/JcVxqEEhaHMBkgmukC0U
CvbEN7d9n83c9CoQJeBPdnJRndYS0t9w2aOZtdJgRtThPuTLsDSAmAZ/1pKX2dxN
NB/lnduoUd8/ooXURPsFgNMHu2UM9wA8l5xhuU9U4acQQmhGw2Cgj1x6K43dhuEC
SqVtpkLy9M3VUKCL04yZE0MU6CtoLCepCZWJpqLQmHCT5GaAg2DtqLRoN+IDugqE
iDTkDkdutDlyoug5FVs3dJOFaNXsn9CtVRilqtzcfvRgaKHP7qWVPjVRVf8z8PyA
mL4XOEBoJUPLMoxfBoqkH3uXqv98Z8DYuyzNrwkW+sOqh/E0UlWnkd4JY71gCDu2
MMxkmPSIRv6p3Ou1TwGU0BZ2uPeJZhDABkJ1RrX1tl7KtCPDqd2kOqgi8Vltk3QT
Ohf65ItaUCyhwgY/WBJEUoks0hC0jMIEhRwPI1iKAayNXo8lYA2BO+p9Uo6D/3ou
8ZvYJtYAAgi/zkNnbItFAxaE59uGFpu1VkvMxzbgOA5F4kueoimYAn6gKZikk8ek
lAB2SsAme6cjZYB4tNcqtW5259ir/vuPb1Ods0uw/M4OutBEj0f0JJa1/UzV6FWx
RdqkLbAWEg9oPKwRXtf3sJJ21XhwGY2BWZudUBa5WlIjoTci94xQrOTkpdmBkwlA
4envmoSx347o5H+M8gUe6k8+VKQsuCIuJTbU/LZL4RZLptBwE9HNwlhJ1dcWH4aS
37BZ4ThMjOROiAZYDJnxwtvmFlhiIwkuWSGRckt8C0eXxTW6n19s3cLvLMn9UZDV
U2WvUWfh0Jz0C009zIWfWqER67nWCYpbgpJJKI2KMIDVOVzhdpkETIrlzJbsl7jC
Ta+mWQxBkgCaDi4zdSypg3ogqXaHQVf5bqHY4fy0q4/RMR/7GAk+6Qp+AKNB8Wbt
PeemzLqPTBL63xOdv8FmHvk+9Zu+TNKGHzZFGpF3tfct9M4JeudKgMBzk2/qYspl
dBHaFt/zWsYUjC7ybgLmL7XSZsDZuhTL3EUbd1Ecq6FDUE81qy5U+3owufwkR+GZ
sPi8YItbOP1ew1TEAGTJ4QiHxzmpqqyhKYpToHOHSRRemkhPOsrwLrQyu6AkFXpI
7/SHxCVd9K0fTL0HEsXHKilxkF73y0DQJ03MV7iQ+FguaSuwq5T5P3NN4edvA3ID
tO8c4unxgr3ZRwCXOlRoyvbOYx8Mdtdkr2PLogA2HvJGfz0vjgyCTgPmtdeBF09I
WZPabskvKbP7HE6c6c5+Gz1l13D/Xdog2B4uvRQv2+ukgo2lTA1smLnTgZwMi49Y
fLClFhVaK8tVv8Yym6DQVuWDV3sjWMU9/89GcXRMeR4p6+32nVMioeBArIR+IQII
oI5zEybCsK3bRRkDH6lny1seZ+67Vhlahh/bEOcgZwcISJwKn3JH6t/nA0UJ9jVN
ahT6zqkhKs+PJq/SdDUMN2M+pXyjjJGBBO6oHJN+jPAIYPwbvabD6nTETU4qIVNh
8WJ+RJZd6kcYaqJGFn9NTyzRP4kK2SO4fP/+VPe1Ek7hXwwekExexIHHXYoU1fat
ZzAmC7gJ+e5yOls2Eo4xDhDw5GZ6jdY7bbAYBDMfzpJFqaJtCD1mC9BzC8UqyXb0
7Lj2SOMCi8+xcLk5xUDJkJUipxLzHVdxRT82buy9xzwFzDmPCMMbZFhvo0a0kab2
qNgjrNXihFvEJUpY7NZM1PU7S+66aUNhwaCoKUMT0cPJydWpkZ9kYGrHwGNucqFp
O9osxUeKLV7JvzTJyYd/hEw4fzmcHTLkf8S/SkX9dp+ZVN9QJ1toxjLIo6/tZLee
LynU+G4XRyWBqYivcEZj2gO7Sk1ETQQ4zldGhhbSRPrIflOkcQUgMiNOfGwwhUK8
RgHrmNNnzEnPXt7GgSg7KYaGgpL/+d04nSUZzJmD0nwUAD+ycb84gEN4o9P6FPP2
dDGYGupjWWpLkalinn4HDULTKMz/e+R/hhi3LblPj/JFX3LXhbVN0wh9OwF3E6Z8
oMu/3G/AeEMZn/fObzRB9czG3gk3cfflSxr9Jf0a5qBI/8qtuoYUB6PhOvJkZqYX
grvXqeJLvQHe4brAYd/0FXZ9CmV18rNmVOupO0DeCZgrKQZODNWCpJRRIVcMkisQ
VZAyHo7FN3FjlIN/alEzVR8JwV1BGm4LJl2P+F2HND+mB1un/T9cSbXg1xLQn2O8
zky3BNeq4ZzOmH7ta+Fkfynikb0sYkjodB6hrVcOQnXxCIwDBoJ/GYE5n6Qc4BK9
tBPmd+YB75zvaZS9m2au2m+kfb7VUUA6P7jZNU4l8iccFNVfEGI/KnqLRIILuIvt
TJyXXmvWklD1tCf90jGW1RwV3fD4NP5uDm+LkUCyLBcaTha92M0AtbSojgty0GYv
6Z9YWL3FnQ/cFLS2t1NdqvCkwSC12WXPEK6jWsdqwJRP2UMaSnEuRL9fHn68nVDb
8hdDJtjTB29nXEVI4JSmF+urIcu9YQAf2Vzmrc2y1Za4PikShOxMTGjVRuQ2cX3a
NIKB6vMemXB1A8FSW4v8CPQv+D0MjMM/pa6lptfufYV714TB6ZnCdLRTXDmxzgMp
zdxY9I1HrGNqAdfpAQcnOs0wclYs/gsPvCui5nrC9wtsraqglxVNQKE6+lObmR1x
3tGEZJKV+WKeuXIqauX2AYjozcVZmnUFAjGnpaNd4oW9EzvLbD3qCYgWr8+wdiSf
Pg1wEwcbQPaErRlmsdZYSGvwM3LIiOFxUJMSVRhASC2+kpHOGHF0hED1NaMf/65U
IumrvZo3Gim4hCI3ohC+jxyG58sKSRMJuCZky5PA6oe+HTZJomk/KUGOH/3gJSHs
9JjPM4ow13xYC3nVyRGBXLYc5sMrBZqpngMew7YZIa1e9piPN7oea/5PzsacleJ2
0jGYh7tEEYXXNL9FdwWsdbRPGWIOVADQlgNTGdSNxaebYTdFXR1WCEujSdx+8kbB
TVQi8LFpcBRxLxHSORQ8PTjgZedYwYJWkAeyjdnq4K3viw7hxaiksFSc5D+udcmb
ufBcyThkqr4qSJtbeET9pHBD+vKcD2J3yy73da4W6HIOGNHIsrnKzhHr3VIfcTuM
dd0No+LgxibWC3bI2pMSv/0quH28Crrug4K4jYeetLey/kRzf9BCj3ddycniIIKM
4S/veHqugfIm3RVUq4bST6sGNCQvlDYW3Gy66N2xCv3jydpE8f1H4DT43wgYZuMT
En4bHo2goGMLCp8FkLF/cJREmGo5wtIP8iMMOBq75f3R9mJp54HFLj6hAg3zSm/I
9tFT0WT6sqNnh4QgEjQI/KFc1osDcwTacBE5qK7K6REV1qxS2oWGCEmFKBqePZxj
9RH/Rp1lsP1SDNmyYOEZK5+u61k4Tldu1Lou6lejqX41hiaLtqrCSNbsrlz35UZ6
cEZVuEYEIRwvucnfYNUTpJKDUHjvLBuQ0M+1Z88f90nW2u8Hprwc6HkeCgLhGC8B
wPxksCIRI1oIamwvLtRcC8YRbVc6X6fVutwJi5/DPOHQBbdCUDj+hdyKaUEFbTao
KRWOyhCVzco5z6Cx23a8GdZl5hRNOuHAyFh3J5WmIqeJWn1RS/qkDaaCAru3gBZk
skEVuefFT2M3v+Cu/T446ATcdiz756WqqJbQuQVOBLERPIYjJ6P7Oz2a80sWT9WM
2YPzRZQORFB0t5fxTWikK4INaA20mlFbsXMoN/+M+HY3IfTiyEP026POk6ZP8pv8
aLudN91QjNTMZzjqEoIWn90vJDUcSSNLMDbThOHRMB1MkSFE0iL0pZDtCy/wP9FN
OOuRTxlIuZ/m3wxWh9l7NAPgWPKSJv3pxBiMtxbz9YjNAitioFpvGB94b5ISix9A
ItelYIGp5k/NQ3I61ujEZfSZiDyes2at3AGG1N5kCQbzEYZ5gB/jYoQhW1rvSL18
PO3rTUZWXXCckIXpo3yvXTdy35yKUKw2FaeBIJwugQFHnmj1wX47C+q7XKTha3aP
6/XHz1ESK1i9vrZGph0rGs5mCBqlLrN+k0i8Srl11r3AQST+Fm0TSuYG95sKDskT
teJpIUqTt+lYWjDnq72AZUviPq1BhsxJzQkh5W78kpydV9PPTIJm8la+ss18ODYV
7EVBQeEYuhLbNlGwnU3qQhtsn37AxK3g/RPitRDjvZQ2Dh5bQF1RzqAr9ymP19lE
nM9QRUrKeqwbgkk9rkHDjcDZxeQrAMATYOo+chstRGRKddLT41KB+Kd8vCq24osQ
pYEcENoog4+kyukWW6D2YAIF97cNyh/iap+FmZ8z8X1MmvQUD2gRCuDu08Jb+Lax
GRQ47vMVBLuYygL0a7D/N9nQFwEV2OchoA5Hj4Sn9JaQQaebUiHWDqpf0FQxoTKX
G7qLd7F5yYO2X7SjGsrjjQBSaaDtCfa/tteS8B4jNs/hFgQeXRXfvACrAxRmLass
+uc0gwwSFcC5zFHZXH0V/5HKYJqSNW2mDfxPNvPM/el/ykN9/FD3l3BNbeiWP279
K+um4ELd2UA/NI5TL1jgQqyhID0Lo6SQu8sKNqJyaDtopq5TckUoU0kcWxm7xXnf
v1xljlUevGpEbVIgr+mtWVWHXEm5E5I8lsqZEX/sOMb7WyWiBdohJry451PFALMI
fIePbOO7GMW6Lp2OyywuZZSt1LBGRcI2tVRhH5YBwFb+zfKAdUdSZXdEhOySmKw/
MYQ5oI/jkG9sG+ndOWsK78KjO2UHUI5pXqLsfwO9EeGDB9XsaTlUFdKgNNJUD0I/
KUJXork/HeSq5yq20/KbT2+g15RN0Scr4Aq6nfvOcDi75Sb2QROUEUdSkSIZvRNG
E2CCaoczxcVDGctuZ/8huKaiwsBThHrRjB1wTlFaCShmU3740XG//xzx2t5I+Yiu
MemEf0/Az5OCEcjU3sFwGFnsqhMvOpSXpTBuLxCLOGLCzkptRLQS87uUiKFnlZS2
gHd4qQX0Iv7/vbELUlGYFh13piwKdnWs4T03HOrEW+dN6L49SlDl2b3HuFzUVqKg
ty62AG9YzV7vSk1PoOUwDkmNPMc2PZ5fMSmbvahGwV7+AsSQZBBQnkM7lGbHpScD
Eyvozq5UeDfdr9OM4e0Jhe7dyn+kyp77xEofXHFUTqB1E5Ahd8HgIaietDsjR+j8
Bs4qF3PQmExfFV+oHJArsY7CVyEHUx8RcjN6ZoIZRtOaEGBgwZRr1KzNgAgsusVQ
0nwtOIgr3FtKLG4OKljF/aByQV+OMuzt7BIZmE4jhOVaA5+JE/slMqkBh73e/CUK
WufKYOjw5cqkegO/NZWkRBKOwpjeRdpnj7ih7Lj4FRYHfrVDChME6WYJxiX/HYOn
6J7ZUBrMDuDXK9tZEV8srZxYmlJeWmVlKLfxVifq6Um+akbgm5k2/P90SAiePcZr
++qSlWblRTgX6hwL5ChgysU6b3mSmh0TDyI3RxlgCOjSrKEHP/5QdGEZd497anWY
JG8WdHR87rjYHe8qO4zbp95wQgF3Y8BfV8dDcPB6thgT8UTMNZolWYO9yfMgA9Cx
ImaHgHqGTi859Zq5+k/0dgzB+qK5zGkLic9agkctNRztmfOuPDsxOUH3rFndIZQ4
Hmx2CG4BOdJBQgF8gvQpirBwifkya0GSxfuwT5+0zFbq0qJ5TVthuFm02m/yjBxh
vc7i8PCLd5vPVvS6DrbeYBFtNT/UWRtggdjQzluD6DK3uWW+pSNtFXl7lqLziBab
eu8J4qFYkwGQg9HsVtkiKaHSJ80SNKXXTBt8JUR7JBeMs+GLd/x97tctvuiSFJj9
T89wH3x2xazysIyTAuUZUwcyjFK9k+kOVsEj4CuBvhlY3ShaAkCxMI7D5+XFnNyf
EEpjFb5TQK5kpygCo1Bse+j1Y9b0ifbaqTBI3O/CEmhaBERiiqTMBLvGCoPuNMOg
WxM/qccfMVGJrWPyrhjXVo39z/ojdYpitkWS2Ps4pq8EJ4aJvxUIjKFD6w9Ctkfk
NsB+2vElA1WDYrIhY8g9XFEkKTwjXvnPJYZAqPNJI0YKYZXC56bzGF3++IRKg/rR
uHv387jz1waiAE3XIuSDYQXbEb5itDNtBmqjAEPjkLrhiosIe8dPRVj+XOFfdP0z
tW2kln7fjENvhRlnCOmJXCsCNfio44mPBdvL5nskKX6wKjFCQCmIl1U14hTvmpJ/
vEik1spAchrKuG/blrL1e8CC3USyBMpyXWTSxfXFPGJAu5xPufzQ2YfxcixCq68Y
MMKPtf5PKieDv0MO5R5K+2E66yaZlkGC3c4JCXTarq6VVr+j42QA1VvByYUbMyjg
K0JaYU7XTwVCdRU9HuhNtyRIHH2xF10DlqC/ZCqsk/wjvEHG7Q4KElKFIStUFoni
4Z0V3b/6u9J/dbwjtjeqNyELx7xZiXdWMeN81yhELHVNs5fv0hSLU+8sqlgDafGs
S1txWZ/FEbzadIK+htHrl4KfKqMa0gegXky76W+CtalM5tzIi6DZ8entB5idECJq
72SfkXD3LEnU8rvwVhA36YakbamZ3n2Ol5mnohq4IxVKEScsgfj0MrtWsZxNIf/P
WzPPBIuVgp2rR17qv3M+1+BA1eO1EtBgsfjUA5vkfonqwbgETRjgwDcBzo/gvDaS
Pvuk4VS237i2J8/32/YO0FntDwwpk8guy5RJvyJWXW76wnczx6M9qOXrIKmxC5JB
KElJSVO8HZNUGuXBrLlIyTlY6j/VKXnRe03vqiPqaS8Oq5yNCMMNNzpp6uQbDyHK
Zz2mHXVG29fUHde8UvdQ40wZ98Y6VD7fn3eeCXoH++PtQDPgm62G6sRbGZO/R2Wc
bRTwaeYZrJ9XpXRYn30tYviiwbnQBK8u/wh9VMLSoUUzPqidvhpnfugY3kzx9W9x
RHe+jzjYvtW7jkVK4RtLrPn7gHE0xg3LLyBw22aynOrRGQljMr0UY7YmqAERS4JW
efh76l2QrWRaHcJO5luT5B9ZsfLoTR/Vgbgg3LBHjoyaCoentLWRUiOPAzqFody9
THZ1CVcp3Ceh96Uyk6Hk655nLRXsUQwaAz9HKLNdmLuYNKwNAuIrCmcIGLhiy1mW
2qJlqjfCzjDC3W8ON+3J7HibskAccEsJ234tHFAxcvn4dpVaEiNZ7pZS062ztJNC
xEW0s4nAN2zMl0OiF77+rLLX2eR8/mgnfHdZicxzIwkb7Zq+gqLq70SWHM8naCcN
4VB2v3ukx51xmTdNalqgRkNxmS0Iusoy0Xg4/OKNIovjg9X3LKsqGHILlsutTJUG
dbnRnNM/Uyo8OegTsCrj5sAaYaJ7LdassNbBVkSI5waLRKiaP29ZdFfzpnZRo763
84lbg84Bg6nBGBVyuD2FtH/MZg8E7VXzXwW6zB6eqDhyaECLi0TaTGtRH289lNE3
f8q1P4MR7+Yw65aB9ypAlISDlW9/z844BSSDD5Oo0Ma/3oV0th+S9yp+1iywxOCH
yMo1LmjGpjpXTZowtfcE+UkFMJQ+qhKCxzYOv1P6S/NJ/HnvCiA+nSS4fHIYMFMM
Hilkwq0feDKrBg0p7wuhR0nnuBEeaPMyrWZmRIglY0D4zoGg3T/fd4iU37nyospu
GPxWqaUQ8LqVdCz+0XP43ITnefMOscpt5k73w83BM6evyNg0efW6v6CvF++U8Pnt
gRla+g/FYClwvmBikmZIKmWakgUOmn/pfNKW6n8aMllKxCKWKT/YCPa1w4pOG6jT
kQJOMJ6Jb7lmDa2R2tDH66Rxvs/Vi4snjDG1sr260pCuAfYEKz8O1Iiecv8zFqxX
YzGbsrtNluHRgsPm5lt8axRUunrWLnyXWT4DKiL6cYVU2cD4Qm86dKgELjY3GcO9
GN7r2wr8rnDPvB+Ei06va7feaf2UNtNE+F3Oc1vwIO5r2fJwMEgweBNP6i3gn8+F
pM2hEgPeByk2RFI5L2G5Tb60yCKSlNUFifpP9N3SFocvfUpIzGMNw/jDbFhyrakD
GsXJ5Nmpp8Z2MzX0dcvkYviK0od+LqxqEaaIfItz2Xa8o4h0X9AsexqBvVO24d0N
idczaZr/D+LxD0/950Tx0fhpOY9SL48nTyX/niOX+Wb5smcDR/ZAMJYKhIXxkfgp
bS3aLCS48yJar8ELDtuc40aBRPQQERKJI4WXorqXc5zoqwwwhOp3K2olnyERYuKt
6XZPKrYd8VGdgq3Fj5kb7QG9IlEb3pMDWgDescLjCLCYVS/myen7AtWYKAn2EJ/D
p5JjHpkXaaF3J+4SDvd7nwDay13S7GFX+P/yw8J8R8Q1Fq+uYdn2eiG9BcK7nnt3
gad1wriaWlBfwkWhh5o8PVxggXu2f3vqbQaqxOQgNsjefm0+gZQ4OMlVIPfb3q7F
B21CYKV2hJMpaYeivQ3iwX8/KhBArsZlKg1wSR/kdc3o48ZPlfbJTd4asPKKUg+0
7PBPvZVoXggLdwch5lK8PKFscs7DGXsBauhu4gjsFDT3JTSEceS6eAJ39p6rJl2B
wG7sWlbhFt+FVudKulWyTtsa6TcfKdrg2vXhkWqS9dykqWpFbp3sgVv7I38muw8o
gGoZmPwEZ9QisyRsSkZnQwxVGbEqmMbnJWl1EPLmZKyup/WXXqURbtB4S0ktTI0a
4TDf+DvCwcknB5fkgrO136CGdxXdAAoSJNJwxzQ7HTxJtqAYnd6lsi99X4GLkeA2
6Ozf/eLHz3VclCxIQGOEuB9zi6JhVHzvOWsVFvFhpw3TZkmhP/2OJqr5vy75bR6I
X0NFmmGup/uHgEULCfa871yk0LILolTwYsFQ0CNqrg4Opmig6fNvgOAJ/PNMWhX1
Gv5tcYnEuG7SPk29ZmTq3ffWX2yFbWx90ONH2GyT2g8+fA/keM6zSSdBMtlWI8BU
XJ/HR5Kc13eZNXUEqeVibbxLynwaACVs93Wf3MiTNLdQEoV7K3tiUyGwPtKIW/FC
1cwKHJKy9w7zOfbdHseWJ734F2wn0fqVp9vU8qIvFgKqWBEbApcR976JxooU8QuI
y38vZZ6tAZkuPQOdfSKO/0Y/akgExVIPXPjqn1XAR58ORTz+qyQ9JenrU1OEkEHK
HRTdu5fQx3ApfefRqPE3veIbvQYF6agdBvJ4RZpPtWIkNDgEB09N/hdngjkoIrkP
S/0sti0ATczDmFv5YVhc169vQEcjQrzgLd6azlbcS6RJOBZhMZLgcPbmPIdBp68a
09/ZHONK4R5+zLcG2tGYFmiAsVvhOZQatQrCYqHprfwcJxyAkMNUIpmHcpxHRi4V
GkiRYlNO0Ub85yNMwMhCZh2Yt+od+Bn1e9gLDVeKVOJeSp21ewkxM8WSfjCyZqN3
WMdJ/ZQk7RqMYt1A0003VLhyrG4ztil+lkGlHE7mUodJIpDJzRKyjOQF2sw3CIDm
rCWLoERU/d4fomHahWFdSvFpG/U9OMOL/Lp4h7QCZAZ7R0vmpf667XOyztI+a3RO
hX6PBPmU8CYDjsA+8Vl6hvMYlJT5LzJMGhXcOPr1sVCM7xiS7OAXcwE7HL5pA/+T
bOCl9Cfg6qtIDJY3xH1rAg7/y53FY/bDoAXjIj3TnnPrgd1EYb843kM6pvtfZQli
uVYRvUK1OEsrQhyalUDfJCjp44hMrbpoGGIafNXJmTmywYivGajclEViUPehCdnV
Rxby3FoNXCccCCfE+xwdvJ24HJ8pFgwvJ1wf+hcGvXARQ0X9kD2U7vbyKJu4hJKZ
vRHEV5zn6P3JluNUrhX+6eXmoEA413azmQ/yAVIQmTnNUojvKwTziFPZsKPogOOT
2wqTKIOe18tBQvBGoBS8U2pkom9DHd/+/5ZS9N9U5nvlQVlhiNRJsL/5gH7yIrPQ
HSCVJFeKje0Yo8CRr/5AzkJyrPgvCGC0QW1viYyxEsO80vFZNMQWvBDbvaVNbu0s
mir/qm0GauOePtTIgVHL/cEsjodsTv0OfOl+Nma1z04gSh3cSrlchDo7SUmNMBRM
UnHm01KK2CjLF2eXr27r4O2eRy7f88LUjl4RihyaOGJQBUEEo7WeO8yR/mGvgNoQ
QPrg1sVBIcysE5cyYNM3K7SvjfdzrySAMG3p30h6qgoj4Pd6xk39omjaqq75ENqn
Lu3m3IDBcprQ5q9LwJHy0AJrLEGptoIQpskcNBIh7x7/ZpAqzpmDTCM3kXcPD71d
sBjiG9+DwWMswhSXdmQs/Ne76gdvwNNKfnqSJiXDhtAkLa3ziUKBh9qWJ992FCbz
Jy2wCA7puXqcuNsnBHg/U7tWbVYSvc0iNxIDPmteddEJXs+iewzODMuzKwCydwQx
3gvY0Ans5nXcJ7Ufh52yMAnZihGILd3KHw1eV2CdXEk3M9ChvfJOqmoTaTSPRncQ
Zmrdc74DLsmdGRv5+6CV4jDsxrg7lnrLRwRULWJaKaUB1/b5sImZG9bKnq3JnOo+
9z9teCzxZafUJinQcqKEzJoFr715AJmstS3m7UXxCrJXfTByzGurYewc3GnoLgi2
pUonLntPBnEjx8lLJ8NcUmxRer1wO12q1wUHO+Wrz6ervSCQjG6nk8g8HmExScSX
2Jz7tVVxMbzqvQA8mWbP/HLZ0bCWoZW6E2slUrNXxnJ5UKZMXF2GuleNgkY2VFuF
ZJAtjp2cE8YyhhEpnl5sRA3AVxOAwPSMElEvj/YL0ENBYe5XxlYXFFYFSZ68IX2x
/3e+j4nzOBXVIrKY1zGkt/u3tZAYLjThcap/T47wQrQ2cfp4XVLaZpsIkKZV5/Qc
ZohK5YOEIwkOueULj7wf14cYdClz3lv2zOPMVhPu2RKWcvQ5ZFobcyFZ0Lg2Or4R
OPlxzcoBLgfKWAKc/Xh2hBgX/VA8YYl7t8yCgAkvl3BfG0tQGMuoAOg37na10s1s
xEbsCvm/2wlVC0xMaNRdc+e2jfe+scz0H7upXCncUhYG+n4V57fwH2VjbKOM8di0
MH9PiD/GtgipJ8rlt72xNcfS2NG3imwTkssePG+Xl8zvoyy5fSvxi7dyM+0ZOUzg
nIzpMlSHRQEQgqNhgSdW7RJqabzQpdOTeloG5cc+y2xd0rJt5Q3GiK5SLiU/lL/q
ZbpVHcVD3DEJqllw6qOgoT7LrQamkP1ehvBGVf54AdyysFzdhBlwS5rhjgMg/KUY
yv2j3L5NPfO0AsrJHTIYAIW23lEw5oQeTxkH23/fQBYHlWU5i8mWg7i8Yb0+LITP
sAyKlj37sQaRb/zRaHK6r8H2dIM7VtRlmp4zqzU2ovbTUo0YeoVuctjGX4sVe5T+
JZea5rMcSXqlsBLHyglcGGIgBA5BrrTqvDztWCLV+1OFE/D23bSW3PVMI1Bf+wLF
9mPLFnb1FwzaiIQlgwHlzJGLTFt0/zmE4olhFJMlQFsRyl4cC7TIHiBanYVCz2ZE
IqBmHYgzEeaOJg+ID4s4dLUKO0qRYnmJ1UuDU0yCQhvTDVdOnNeNlZxxhUHASjXx
nb1uijAV2kRsXvJKxLCaQW92wLkKPXBXAbT9s7ug0ag6WUQ7zF0K3cnYjP0q3jm8
mi4qtQn6UZObUY9+hXH5BwZnlXeTEU/TWGlPuE9dBAT7uwgtxhgobd/+y6fVsDyS
KYhokn/krDymjToh9uCK1CUnbA7TWkkNYYVGU5m9um2DcnqwM+mEJm2AFaUUzPJh
UgU3qzL2afbfHl+Odo4q8svoR9u47FtWtYSfr4FM447qAgZBAXSUEDAz8xHEHjL/
ecEaggE8sWpcGxdfMcgblBEbzOF62twRqBCIRXF2qUDOhqbOHRVxx/15upuxZt58
pAfxTw84OW105hBMRTWWC4eh+nl7TJdqRWMlll4KAVZk+wuFuSx9dDkNfrCBrDkL
PdR7ZQSX4KPEmjwEa6LYT44jA7X9wazBTIB/zIL1V1gFhZG0m1bh9iPPpTbs5jW8
cGD/WqeBrWGqUeBEay/u4mETdMimbWVYjTp8uyUer6FpqZHK2T++EZ4qUf8rXl4K
XjTuvzGWuJltBu5lmmbnC9rhtekgOlfUP704PuEG6wZHi2z7WpH+gkyz06wDjGTw
UFIo6nuckEWw8e2HmTreDHiArvpz399z2mlSVE1lvSfU+Iw+d81TdVjljuOdC/eK
FAfShUe0pNg38WT/Ve+BgtIG3zeJtycablHDYGgr4w2QuaePUOv9lO/2IceiYq+g
u7uvhp9nXRHNTnqsRG2OFwfTT0U9rl2cSyyVtIcHPHBnlrLMovM3OD76jcHm6esi
kdOM6TkU8G8TfTgobpOM4FXiimnIkvanZx1nV4oMGBTNvr5gCeyyrlYUQupzvgI7
qj6FPJAvEwz2WkoJjElyVUao/6MfoG7+q4Vl/oBDGBkyPZf9vNKUiGV2iUj1d6ib
Umlw9urBlnWjchnAUmrMS31kCsUyu/vLg3FT54dtgnFyuMCh3ifJfCcHMRY7lJ2z
GnMtjTL2CCtKr68iRdwvDTAZRe6CO7fFP0TBf/HlH8My3/lH8RTMtyOJq2G8lu3l
hck5K+sF0kWFjR+ibQdjpzf/3f5mUpShS6iJaXlDe9rCb/qFlLQtQeWYCwA68Qlc
MD5iQx1Mqs7J2Gj8PWSHXhZQYCF65lnk3kv5daCS1BI036D1WcRiiFLWQ+JnKVIa
PPqhZ36TUU0+tMTKsZhd5mBikOttjZ21JvNoqXh65nMDs7b9TKnVtRob4XAnMyAJ
0ATYS1PYyOflTqNaNDSxymBh/WUUDLcLeOCME5E19wM2DLSkya3QEC0Bv+WFjwHw
2kF+7CTCYE5mBQmESjBPQUcjQleg+r+kyiBDuR/gIbRgAwTopVATF9Ycw5dFk2BY
QpATetkXe/VUh2MyrvVx6pZsraZjXJEXs953WCMp3Go0iNIH8KqVAwIxHTLuqAh8
CbnbCJINvUEC5cMw6i4Z8c9CVdjTahMWsl9iE5WuWj+esAZhlhHt8Z57EPYwa8LD
5lbveRJkA5UjO6wkUTxqHntnoowMriyB/U2H/n72XD+uHapRVDdXOcRWE9jEtR/Z
G3VfLZX5c8S7vBIiVl6BAcluG5mWTkNhsQBins4Dds4rC98Ivl+FeJDghkJMAZnF
GkeSWUR0dXEwBpZ3V2fh6qujJh4FSY0BGE9LULjOJOQxyGtohilPyHN60A4wwj+H
rudPtVB5RTSS+5j0DWNtej9Wn5D/1kPDJJCln4LPLtUNGGBy7Mjee1nQEY1WoDO1
ccVYTvspluvAG78ujWuASeCVdKIw800qXXAqdh+Pwme0WQIf+5QGdF0h7JJzg4SJ
mYjNgttFjKNjfAZjZEADldm6HSAa5S7V0J14ysp0MTnyEQYUU02e7GTJi34plnvq
xLo98t8bCsafvsJ02Wyx3S25ofIkhbkt86PmQqhzA3cfV0/kdbW424ikNfI7fPSt
njrVyoYon6+cb9GXaQJhS4XkbyYb517yGUCpkQh99y7sc7Q5tAZobPHFm9edu9Hc
MDmz/EoaEM4sJqVLoZ0FHtaORemlB8k/0U4o18rG1XP8zcOkLdAXwDcuE1Q+4IVH
bla3/lf9e0bfSNWH3k70ITFi9XSj35nsLAGuATdcMLeWMnpIBp5cq00PGbaY2enl
CrUXrtaTGKRpx/VCkCPXBeYfSwkgGQfL2qb6m0f+f+ooervwRwXWLdL9T0HV6Dqw
xjArvm2bM3SZun2MJ1h42nUXDCFGwdjVWOlhGy1VI9xont+1Xmoc9abwg19VR5dD
eq40wlA1ViJWJ9t509g6RU5BTwq6Idjnm4afltDL24W76/GqvnFr4nDrlHfRVoya
7Dfv4vsJPQ6fRl9gqhRiIe2I54yuNHOTKZo8zqK+vj91KfTvOfi/NlmdaS3JIEfC
ipQRHhBOJVbJKq8VvoFzoOId1xIn8bck4CiU6Tf/PF+Rg+6d7vGvdyNWeRo79PhY
dfqB7njhn9b++iSojI6OahbZvQ6y3F7iWEHtbABfSOPek1ezQwtNLcC5IdtQKB6p
QEzp01acchz0h1os33i9ON1pAGGxXWO4PoUl5UP7QTShaFgT9XXZhji62HgJrPsl
nuFy+0gwd7G6zLV28Kuu9b3c+0c4zREvNd5TzcGdaY2m/g3+Rnw+gExWOmTBn2kI
ue0qTSWkHQMZcUt/rW4jhHRI5FeY/KxRtCSLqtUdwBQzeL3LDvgIktskL0LkZHeu
dPrCue5zmbFHCCXG5TKSln/vsPKJ0inrR8G/B5DSN/2IlF5A/mcKutwRG803CgiV
Q7Ft17aAxAvWVSMIUhoEFHBVfTUKh9uwC1tG6cvXIf+PqrwstGoaU5OSwOhKrC0/
4QHSYAFjpbT5oiBv9xWQqNADRmvRDP3INT10ulBnebGGsHTTM1bXJl/X+z9REJN3
DTY7LhXFmiD4jRWujIl2Phlp5yiNYE7JeX9LgHB/GcXmrY8LfUkACGxqp38laN40
R1RX6069DBNaCFBiyYL9xWEF3U4Ru3NbK3enANlNYNHqvcjAW/xJNZm0iizDFRXB
5ZhTyctGpdJ8qcV2vf53HxkfmEA0Ho87YC4g11CnI+z9JwcxxmS0CTzh+IeJcFMf
BEQQ2w2LQMSb+ma84Zg86AB8+nf2ZVD9HjTCKZfXYFLyIxyhSR+lf+YH3rN8f8S3
zRdD5bIj7B5gZpJMTIfhh/UGQuPwRHDSRwoIhV77EdTj3HFKcLM/X1WpESVHGfW0
zzeXXUTFjvbQ0zHRUGx/F2tjEuTqNjrMQI7LabBhr4spKgo8/A70I0g4prn3yd/+
fyKfW9gfpYB4ukwcc4J/ivnePXv4piN2OzsfX8obJhBftSYmKsEB0M6Py/30t9oY
fCP5c4vOttQybITYWSqybwbbuMrYHAa1dPzBgsQ0HbKXUJV/U+11z5uNLO1zjI6u
CHGSH2WLLzmX5/6+phHjBdCmVQGC52MU8nTWa+dEsyNcfSoaqp36va7nWodmwN/u
FUI4PSUi2QxThE+4AG+uWe5jb4sTPWnWcMyQYANsbB3+hWWvBkGfySOsLdItQQYw
uVrJmLB5G+0JkRx6M/xlgXOWFlKEb7vgdBwf5K0J0LPfGx9mULp4GfCvKz1RtVfh
9Z4//YadYQXLv/+NMinsm8fSHd1z+7cwtqJ6gemy++gbMfech2YmD1RIbrWllk/X
gR/AspFLPA3tUG4ah5POdZAKSGdrZ+T4mnJRV1aeE+2ncBz0IyPu/Inpxws5rJ/4
vaIgGPQBSfTfj4Ck30pQztbjGQHrcC6TrtrOLQBj5z+x3jaF5zagAPjQ2vaR+2tS
lL6TVixOZU2A426e1ECLAHIiek3ZQFxmFWa+cwfMgFb9y5+X9g6Tu4rvoTOH7+hw
nRVdzwrxm9OIbY2aWEp0AZSexenQHF/nD9RarAG5QesW/tMXVPoER6B5SGj9iYiM
H3vHMtQa/2FMuxhxte/aQN2q0m4GrAzy4LgzkXBdzV/rZZpdWtWAzf48JpPR8ogf
3BKchzzR8RNuSryc2U8+whEItFUjM6qIrpQeEsu/w6aQbDF5fWWMrsQ8c5ASppL3
oNB5ipIXqRcVPfrwIdh8NPkUqhKiQ4k92nEYsEhQh3K1Ohfd/+fkSaoKVzEQnqH6
hoe2IdFk3abeC7uc7tQerieTqEJMBU7xcdneyoilMReGHUbWsyDqon9cXUKOg5Sy
M3T7YibP2HRXgXtLo94/VwzC8m2z1WraTUbqy++Z1FS7npUnT2+aZWtaAvtNOT6e
xdSo0CMOdDdF3Qy4q9zOlYVJ+z7wdelWoWbUT31Ml9PzwPwSatue7U+cpxkKvFCy
M1dDjo7Y92ihS41nYdCDAlhoJVGe5eU1yg6ber61yHHYBELrr345HaJmtBd9iOus
6N/NXrsTGN3DL5PN4AWkjC9t6Hmy+j6kaTWGA95LJjT/QfIutGMNXTtuZaVLRdb6
dXhyNSjpLdmd5OfsE3WfEudI4xy8a6qsW7xl4GAV/DOl7DZJ40K7elvG2hGgOWrA
K9Qk5AHQ0etTwDOVmXTVAUah497TR2ZINmw5mcjamBJcUNwuuSBrJmWoPxvAaiIR
mwZMKALA7xgKYL0klvHFvEkqA9izRNuSwUqav9CpkZU3pWP9RadCRgjOpo0t9elc
ibL3oDrqZrl532eTTQ/BYcPWLWR1CMnP9dvHuQgg7eOozbux9UfPBDQxgEik6h1J
+6EqhK7NNMPJr6q3ls4z4VkfOgTA2nPFHdxwJabKLWzF0qIG8FU324yf2lWo0Rdh
wA34EljPQAkNsfKELBYPdWlrKdjt/iexveXb/2pP1caQt72lyAhjtQV24hFbiCGx
Q7cWu6iHUBMZaHP/S9web0ZZy7+KFQK7iyqnbpWyIQDuSXqXsX6y0YjKhOieRdY9
d7TeSuCy/Dxh6jVLCu2lkoQdVrIWUmHoCsOAmN0ZL2yDWyL0zQpEo1ANX08srdM+
L3arqxWgXTrj4qeAV/089jKrLwhJsFFMmdpRKdukJgh7VQV5+SvmRz7RFq5vot/H
LQ81AqpTu3KJu5chrokb2Yu0dfvuYifgQHgUv/vP1Ke/DjLmsQq2d5Ve72xBGqnh
jyyha1UR7UYsE3ak13k2EfNnVHPDXgj24cX8+Om1JQJq0eJl66Nc4LOJJq4MgS6S
vEfsfDipxWNKwNsdSe1j6CUY70wMjxGbeMuiB3cVrQ9VWWjPv8AEEOfSYNP4x5T/
EhzgfRJxQxZi1DbK1r4GWOu6WiQqKyXi+czMrdsXpvv62KXphTac6s20Z9xVGW3I
d1oE2a+kCPGbUfRe0IynzjQcF48sMyDSQflfSwiRDoyTPqPVyHkuorqRQYbqcuXn
CG2aB+0iINHVv7ZKo2dJUD8vwxv9acYMdhoNyntgRXL2EBKJNVvWkvNaCr0EOVVj
2EBkv78NHMfNh1pemdA2oZoho8oXE32pLH0Yj08ihqtT2B3DyfPndtAFPJeUXKyX
DG5iFiTVVUMVfB+nWLiYPdMM1cTNUHgsNbl7G0vx00Nvn4n3sCxOI3JsrxlP4B2r
FgmaxzWmW0/GmHVKqeOg6v4GPBDi8hCopU3k69vKy7Qrc7jitF9EoRa+Nb7JupR3
+RauKjdokPKfovYdLTrdOiqOH66tJ5FIfCXLJSBKpaLsqt28pYZxDYYs0Gfkte7X
W8RPDih76dSFJnt2+jEclYS7NTdhBi7p+kd86UUEAN6tRM/+ieAVd0sH3ZbUwssQ
YHYWzQ1ZKQK8JXtg90cf+AsmQF+fq9a+NmZ9eTKsq0++0LCdjTgNHm9WXjLAIjGM
c0tKOm66IYpPUZ6L7Oh9zx0b7pUKULHyXUk+AOr9ok4qvV6h9oWAvw1NTm/XVKkv
xWDHe+e5klv0Bxu4K1ZUN6tsanc/GzJdEValpG7p2OiB9syONZehLrWxEOsTqJm+
cPRFg3hJYc9icv6zMeg4krXZcy38R9sNYFHbeg9LtnThJilHnEX2GTtxCQKjrt2S
0uFD6VLqRuPi3+sPTwSJMiiAcEkQRb7CHkCcXEyCqQm/jz9Wd1KsSAO9fDsGbBqG
3NMAZx4C5tSPLAMOqF3rA8rlIhpIIUHVNkpCP2sTwfyJcKyQK5pbWGclMYtVy36U
kRJMMoGbhMuNJTG+v02a6Wn6DbjZM28bGJs2cKQsgHEBWQJFjtEyLpk1Fgcv2Ja5
7NiAieJ5faeJWmW+lZjMEvM1PBH+IuNxXKv/vdBpEZLOsoA+wvHASzKU+vQ33OMN
alofrRUAaMCDokg1kcr1t5C5cmjpLzbMzhzi+5HCECiasnK92u9fX+yNgPGqUEot
3FnKaR895RZ/sVGtdF0g/57hlyOE1fJEl1jeVogojY+YLWRNLpbJXZPnBrWIwdMl
bQt+SeSAhAaPlfrCLwGCWRvGSHeQayMoe4dbTpYXO8r95wLiKoqeFI4Ycd6JSFcW
5tbnxOTXUBnRNkm9yWszsAonWgNZtAI9bZ5xkD1ql8p3Z9wZSR7srsSXtjP6JFZY
Ckz0y6rWr51W5XqLwl9La+n/6U/31vHyj9ySy0eFOiBg815dOE0NWnWz4ZMx47Cp
qZunWpDRxiFCo5UJljpR8sUn13a20pe20QndyoXwju5Av7tdhtrl+moiA6trXwj3
kZn/T7S8bPckcIgpGYufAaYJ59yUQXCgVwPoq8aFNdoNcaAezpGh44NZpD5YLeqq
uI+3/lbIuYFs2018gFDX+lEW0MY+k+drzUTuhwDR4TZM1DHX+Ot/v8lDgrR1qnvZ
1J0wc5Bwg1qJRkPMnqyaylS0S6iztO+W+PNdrQQlIgskfkzEOZM7XHSJlyITRSb3
G5kMEefuNzH7sHUkHHD3VIQSUzi4xt1rPVGRsIkdvdHSAXFmq4+E2+gioDtEfrsI
a7u9HIPkEXHfvF6+7F2KCpN8mlv1WwkGuKOmy1OWTey1siK+q2/TtRKsJNc1Jj2W
7oYb4ND4RCCzeDZKGioKDOjLSQRLdAqiW73+ef1P5IeVnAhgdsw3mG8QApQssFRX
YI14C2go7P7nmya92417oOh+xvjNUDB8idfniRXVahlBSlELrSvTzDwspS1aQyYn
FfiX34QOPOvFmhC0MacKBQEqXe0k2YlqwSqUthEcSLGpnT+NocCwJgAPzAJwdL+2
gr82O/xDAwSDmj8rKbRvC84TLCosBlUeTq9WtJD4NuVIL2qreUUNwkvyQihBOOYQ
xabT8Oqxh4v0/72O+bm6cfURxcaW0RC0CjAZFoiaYze3lqfzvh7SnZ+RxIm6xBMq
9vJsdxHMsEGiUuQQMv3z+UFq7udwp4736eZ6WpMUrjNnfwIK1QpYK/KXZpatNlKa
3ywUzRsFpmfshLmE3XxgwwJQAhzeo1mk2w577oZOKTbCvYgC6zJC0PpQgJ723VIE
x6nO7DYo/dkpm/ztZIJYwarLQugZQNhS1GXOuE5I9NqyA3IsUQ0Mcg+jy6K4Q5N1
eRe30eIli9sbRgCiqiazYpBaPIhX69tUUR5PuOFsg4fy470L6Ad+hIShJunW2J/3
9btkF1cz1kOagConL+bXTXOpODJcL1hVC76f6FEgXgFmdAX3YWStcGyMF1/fMAR1
Qo1aWIqaCHOj5WQ2n3sPoR2T3NsN0AgUYElsGW8xWnxmQbGMFKVm2M0heX7zErJC
li8I3P/vKQTFMnFjQwwKQuWrppV5fA3Qe4CzmdEwdWDQqGzzGjMu7X8MmdBgDeAy
HhcTvSO3Vk9ZfztPRWhpGbS+ekWkG9iuDP7jh95h6oi6TuD4SmIuw78Id+brrWmg
DeOH44PoW8nTREFg/R0MseAWDJX2PMgJmr39uBxqvGKozD/008BLd7pwrqkiV8SQ
QvBzECln4yWcNZmqigiCz/uIB9rbQPoFLyZ8b1Du4BJ/8mWzsMg5exPCFm3cefFk
60ESnW26w2aNp9ilxNfZhVPID09IW8olj21A+fRzlOEz1dgh7FS6hKHlhOzqrGQU
OFu6khx/x4NrOWX3xUa22v5m1yS7O5sstYGDKmKIdFrUJCTdlbKDTbl5PZO9tab4
5eLqZf6HY8V96YG4bjLUAqGq22WqVPFF349rUahFw2JKQQK+JKRvbRfbaJbpUQcw
WlLO3WSlrTTm3cBIh0cfByWLqr0iUSpH+k84X0A2n6BVFzQdzal+znP2+lZriVyw
hUr0DrMcrygKbfXTxrLaPKwiD5kf/Ymz14k1g60nqU8io2YcLjBoPd/0A9GoScSx
yqEDlKy7CgtLlDfmdAk6xJgHjcFThWVIRwQTXndi7QkSjQKD0dmw7IrmZvKzV+rK
fyJj/C6uhwkE+tMMQa8CBGVQeELZvmrLilP6TSfGgWBvZFZItCx9pDpTAZTW4+yN
/WyId3+lfAuB3WSotVdzRNjNnBbkDjpxyOGtqlvp2KKk8pBMJIAGFjCvFkIj1KK1
kWayiCnaArvXxIqiNbJ08bwKOKMka/aqoqYGI+xOO4IuZOY0LUmyguV0xlb4fLrK
oruW+cEmFx5KP7NAAI1ZlxAgyPI5V6uPAj+qhsEQgl24zgwjYR7WbUqJwanm3Scn
QtnrllFZodE2DCpbJoUKhxltKAu6N+IxjtBcZCjbh7Fgg+Q0pzaY6zQyGl3y88sy
EL7FhbKFermiyyAyYUsqbnGEpefs04coCYo533jcUD3aOQqr/zw84IkTwMdTcj2/
MDgjbBzuLZpmm2ePcTXWzQ3hOhNZ5gjyH3UAzWFD2XTPJ0Z3LTCm0TsfKRe705rI
Ka5ABVRuCyoRlONdZaLvGm15nknYYpH/AI1P5ozsiqIZhXh0uadxdbV4QOkEZWI5
MFfEDKwwYCPo87fdL0TjlyCdl9DSVDZAbuiW0kIUMEshbGNrvzTOr48DknjquFfa
Kk1UvLEC8s58epa7Z9AA4tsrecHrGxlWUlxS4FJb79SJWh/5DrdPv0WSkDRfMlXA
CCc2SWZE+kta1JUdg8INvhxfwIVF8bRhS90UpYu12aj+u05GLKs1yDctMmF7Qgk/
yC4OHAkBD9qwocdJz6RuIIbcqtdGPLCS2v8MjMf7zrwnLWvRvQH7bxBwdcr2KRvM
tL+u7RUhlDtpD9vilbPGSTtRRz29nDAKTT8PqCmDxqBso5u72G5SUdtwzmQVdX67
0S9EXSrVIsHHn2aG9tbenzTvgWOsxkSZZ4EbAG55h18VHD396ETc4uCqQs3arxAX
R7+QwmyREBL/S9scRemGP+sFSV8Ddo5GMMUVfHyqK82PPcDiMO6p/WrFaOr7lW/W
p1cGK2QzGwIb26IWQ/XFs6vcHSTUubwg/tQDum+ZI2AtWlctoVr+IM24xqmeuZif
JCjkpEHjrTo1HcSYvyJ9VA7hXd9CvGP9traofnBamamskKIKuI1VjehNyiCuBPel
+sqmXgIcaJ9Rbi9zmNFFnQsy2oRcsO4Kmqz0TfVgTILnrE5SH0r3KdcMj3a66gKI
QeNVcz5KL7c9HGXezT0gV3fTxHlrVKlLLtArTi7NR+vR4ZkG/VTNNenpgwe5NXqV
ww/5BJ4qQfEfSSC789365UN0WTLGjbzEsk/u+TM10owA7FzCb05bArAtMHaMLG2A
9CW9oI5uyvIASEQ87w5A3mwfbfvZgHPif6zeK4qmYs9R77NS8eMXeitzAerRwVHa
drFNEYa4s++TFPXgwPgemEeFsALGMc/ATNOXMUv36keG3PjN6mK2BZDOp8c0SRJK
4nf0yjUm59WrrRr2CjnMO71YQ4wfU6SSSxW5T/oeqrSU7IbCIHyUWO1fhBTbz/re
Q0+RH4wtkwtzJNWU/CcOWn7/rg7e4TqSVFK3PXJx5z2ssYVziHH3kGVyTRIi1ZE5
K1BryEivx/zO/b5GZbnbW2TpRpifP1MOaxR441Z2Z5H83V+iFmW3bNvZnaOpXGEm
/F885fczfcD2TmyKNISQ5w2wBC4YV13MZtCkt1XVF1PI0Kntg287cdMrqdzgiRvF
zmvBnLP2qSyD2kF5i5I6YnA46Z/aTn9HXz3N8bLKHOu6tGwWyqHWyBSw4i5UoD36
Q/V0iwZiseEyOppuLCXKObmiMl65kgufCttOGxesHlnLPv9LzYijkXwDRXBlZ04q
odgw1m98KHPEDFxPph3PPrzk+djsUwKoAsNq4V/BnfSX6JArESdSZIuZJIIaL+KZ
SGNJQp9/CS3O0Ya+7dILevJgCCIe4yOoBUxNCpNsM02lfnSXZ0xYFQpV+FQLLnCN
c4aCGuAr8r5s/FXVhGtCtihbqZHO2G0gBXOGlQJ07Q3XiTU1hVXj7nCjqzb3INvr
8WdQPXjgzYfG3a0N/unLXM5LrC9dXG99U9O1XroPCWIPq27c/mgvIGploTOc058s
Nz7CW8pArgJvknSX1QRDhjS7H8uE2ZK3oDDdgn1bxBrrLcJaibcGDLxYffUo0R2H
zAvLNyenKp4JwmvEdxoQQ3x5sNW7NmUuVhYrbow/oNlsrD410DO4XMFsRRLGDkjg
O7wvc6XU34vWAx6npzfDZq8QvVxFCHNgQAPBhX9ChJu0+yFGIizRO/pKxkO+uhFD
qImWQR8W5TNJldXb46ANrUe0vl7CharPdPTWrsVnJu0SVbdgNEYebOnDMqyu/C1r
Ia6utGfyhHa1R4JKLUSL0pEcJYNznZUFVdJTxXuNznyfr7C0D1y52nCaMWXpsbVT
TNb2Eb+QRg3RO/dcLyyRpj93eTsKFTBRkTigmUa5GLnElFnVpLMx7CoMCVQt7MZx
ppUrlx9Mi3LPWVoiZiS9v0c57SHy+0UJhWm8uyShtmoo5iSCfsTqIHqr3ipOneBe
P7+PzlFZe9DmvaZaCYCTrcnhXvfQjc4LgCKx5TTCiMTCnnbz9JtT8FxG44xdSnxU
QbW3xInkNN1e9BvHgrQszC+llRGJ8i6Le5OHdGSX29JVbYrdH0dDtT6ev3y8iGew
p3e6TDlwvVtTOgKjuXPVg7pioUj/UGbTdqfm1MCFCjPVrXUVJ73qci2zAQPHXO0B
4tQCbP1Vq89m2h5xlvpnMTgr8Ugr4l4dEcRYp8VtNRWVr5UTyexnm7tDq8wUFCHB
P8djw7wMBsi3iiJu1GpJvTvwIaVSprI+n8ZEoU4/3rmnbs6y5uQxUINWYdEZY55O
td56fb0F1Mwxr+DED68d2j29/FBloq4CRqUsryvIFgAoqcLR5tGGWQTLftBbLmgJ
8TrNpLOwerBSDBPG9vc6X2IEsz0/Uyp9vOIOX7RA5PSXjSByV+hg4hQAuQMWa1gx
lorBj8CCU72SPXUAk8PEZw9x1lwF4zN48FsVFiPa3AiC55aNOm1UQiOjC+Hr/w1f
ThcGhr7fpLwjOhD9OzGuf8ec9dcqrdDUUPSq1rCJ+7B2KEWFh69cIJCqwy0PmrLQ
2ZEn7wqek8kZmauyZlaeurpNz6dg1UgD0Rr77ust6j8OnChjmkSArsJfyGZf8v2I
L3c/94dTCaUFiRf48o1PG48I5EcaggGA4rPslOq/6gVb574ZI0AtS0Pce3oG7IUF
GHPYqPZL5xL/rW0G4/JG+LV6Ea0C6YnwCIxKzd/hITY2pDXpnff3dtXseR35NT7K
G880FANsLJaEQXOPI1y/uv2Yhwne+kyUjPcNe7+cOXK2VmiZg0olDNgPC3/XEAcB
p6ALIVEK3r+GBD/DLvqPaMJkZKYesnVWrJ8n/0jeNPyEItCSmsA5aITwh7NA9IrV
2gpwRd+LJJ4VWCCjniFxbWJzwbWTx7Yxl/0VK/Nz77mn7cE7GiGJ0dqWfsOMKqIe
SHUcDt/o63MCGTHIMEhMbuKuO1bVyZz88s0a71k1I49nTiPV86YpvVFE4FXZ1DO7
t0WhYceufTSj/3rQrG6zbaw8xfkbA9hxi8P6/qqNKbRiSlpJJK293MRnK4qMC/Zw
e8n9GuYsJX60C1aNXJUwx5xrbAVCJQxzpEwKWMWcR/6yEI07AJXRNtCo0UnWNaoU
uzpq/e75N0tVs7mlTMwp1bXqIPS6wPJdccFohDpn+y1AnuSgs2F0c3+57oi2fDNE
e/Sq+ECslnNWJk7mVMCHjq6hYitWGADSH0rHlzPrTTTiehmGvzNtNc4PNdAfnuBx
jKDUgTWROu4HHnhcjKY1V+IH2w6tDESULXiJjVGe+zTAE7GD2f/L8qeo/uXRZjSy
YYx3f7BgO5ohVTtNl9KXb0tHsBQk5hKl0O5/YH/Vpy7UCrT7pMopveG/UcJgwn76
B2S3mcWV0XrEs1oiFV39nKbb4A/0wuiFdb5pfqr7vkQTg1IadAFz8XE2ZZXT2kc+
xdcYf/hSj/I7SsIU0xTDKuT/P1CFPx9Quy7dLVWUGErutkzh/eWxiE+x/E5/BKJE
hwGbTfZKk6djhYO4yH3v6bnTtv1pfa8lgs5/DBhnjoa0OfAqSDbQZVCswMGAZ0TW
8nfhIxo20Y0s5n0f20kIc88BNeNAksagpUrQuUtaYD5N74nDbTBN/92QTEIKyn9B
rN7AfNtLUSNDjPzhdd7uXU6L10P6AWva3MqAnZnaO+dpBapKsGKP3K2o86pWoMFP
Tk/ng6vV5OXhygs2MDzetOxU6ozpOt5OdVwsIuPZ4iFf4HjHSTS7nXxtndMSv75N
ecXbjnl56I0jcUaXj/kYirKWBqgGpWTtjD6/VLtLc8097MmrvTpJ8SwgwiSwwJCF
9D4z4+P7LrxjpWnyyjQk/xYHsXW9kS0T1QeSnsQiDkVFvgPLR+bkBj81OKszmu0x
6UMkbFJcT5Kn2Z5OuX1dwSqrlbtYDx1PDpQV5StEhGuvjBuOuU784ExMV7Hir+Hh
PUhfPjRECL0dtadnTTVtsLhUU79Nb3t+WrITMaZmtTaqaDiOjHU281E9IzkJJAg/
lnjyYEab4SW5F/ht6g9kXAtx5JaZPzJCEWsn9/oD9sBB9qGi/Zp6e0EEhkCS1kWF
iL23AEvpBRtWa3W+m4MahZwHIzmoLQZJhzBbkvZq8JqMSQVHNhpv3+avk76EkkOB
fDn3kzoQ9Ps/UHhuft8b05UpUcEKG2sVzyUl+EnuC4RFM1n0CwjAVqPC5JOzQbTl
CQldC1sw4wxJ+pQv71p0ehhT5YW+/FNwyUpyaDJJdnXsc9EDl9Q0m6rXq0Z58iuG
IkRGfqiNm9HNd7eHCJe+t7VTKmgP/gcqi896ACkA5wXtWuPpPEf1AhRd5H1HhmA/
M6cAq1tQG4sqclilw04cr+M6Yvk4LWhA4fre7WKck8+uUVB9xA0gW6Kr34StHH+K
KlnUEV/GrOsyuDiSaw9cOX8W1lK4Cu3MKnSo+/YbK1SlRi+Pk6TsaQjWI3d4AUmj
1DZaV6eX256psW+IfhP8bDjJZLBo5RX6b+cJrDcpMzAu5srWfg4edmPAi6zEoN5s
U2iL6aQfEmKf/g6nN8gAWVYP+iDNcujdwGRqKI38xMTaBI7Eb10rPyrlQdXDuhoY
QMAfwvdHKRDMSsbuyPYwvqI6MDGLtcBtpNp8A6QyIbI/Aqo52oqZqLJdn4TGv/zL
/fTR8t6+ue8MlRHU5q+g0p8ViXAloaSGQ2S3NHcbTRjAGAKHsXUy6aJE7h52d4oi
tEGr6JL/MZizUQycQyNuqPYYy1PewpnR/h1jMz3SvGZV0LSBBJCXTL5EpgRx8uYT
41igfEx1fyWR/CNmJ7QGxvITnevVZFLYKhZWKaAoyIf5vfJpwjQzyf41mnBLd4vR
NS159E8pcFp0Z+JAKnVvFheEU7JYHmarBR2RyqDbTZkSOkionIn6Lf0tkFtvXaf7
2crU5xR57irhh3Prl2uOHxKhy6MFANU8vKOC6oNPLGDOWer4EWv3OaOIwFlqu4g/
dRu2yMoUJKvBvbxhqnH0tIrw6B/tozhF8clZ/U+YUbpi0gvFPItVvHxuvV24ae02
0YdFD0qz8OfzWcS2YuRvRhErQ1OVp1Kel23XQyrMr8fe8ztkNe2kQvvWtP9qZBDX
qVZz+Iv/VNcyrwxWZnBxwY5HF0yHFm4fLmgkImn95lDF2OECHXc3NT7nWFUgBlJj
5k7Z/caW0MjRJGZmELoDKpR6LRIhBHJmT1QW/+SdBYHvrltj2DicTy+cWGPEaiZN
/EI8gddLFmURA+uFP56O/NArdh7qz2t2yPtNpwasQf2rZAkg23AWceSOPu7BX5c3
kmv4UarzAn2hBeYm96vzx8MeroDhrfjb67nLlAqN+LHCmbIoMhv4n9Ii/x+uGY4Z
3tYhZ+xF9WlAMRByNonBFbSFZ1hJDMhO8XztJmWFeo6uBpNPI3ig0HJOIPSxK1t9
iVPmC5sGHAmh7JiczKjUq10WPgHwT3SSv3uBDzRbXeIgvHQzrzQmo9ttsj2rdpbk
e7l9+0KDsV50Vq371FNmiwKIDOs1p8BjQZp5IkFGuHOb76o+M3EN/7xGzg8Df1Z0
DqfRBIIu/dYnH7R3X425Kp4Rdc5xpD7Son8XYgn1W2eDAE6FOWEx+FBYYdnwWMfX
nRbzjeevY3zY3lsT/uvp3WWPV1R1HOljC4Z6XOMSO5cYAwszZUWYRTGn1mQj9h/x
v5kT7qI8/igtcheBr7aT8a9IqTetDg4p/efTm5uUh18oxe5IaH1dAHl8xo47XVfP
oDDT/vFUlHj6uXjzW0biqef5jFEQAefwqDp0ZJ1x6Pc3lQzAuCxOEFgMI2layCvf
EjzMlCIIiOlF+kPur7d+DnthnOpPchy4UT2Sg7tvD9PZJFJhcdxd+zKNmssswccY
7RLz9ljZYgo4y+wAAFEkJNKed6QXi9sN7C8MCZymyqI5M2aywnUxhZGxahlziK0G
kCGqWwYX9z3L71Kz/e4cuR42HLAks63yGjEJEMRCD7I1VeF/1dDiBwbOlnud24p5
SZKKmHpELGDKNk88ARpqC+xDQc3Hg8xumHbn1woU/x/J4LyhlQQ0PT/bDtdGgTne
GVKzZzXoMiAu1w+vYcP8yMNx/7iDjExp0y+V/JrmGE41czkt1eo9wlgm/PNb4331
TDGrtO3B9cEgnOaABswksw7o4yXlmilSrd1RlrmbnJOrsu5ZrU/zg4ZW3m26eYgK
NYf8SDmawQErUjPwNJQxAYcHmVzerzwJraWAV6y+xL2dtwT4bz4/0Py4L8rlCcpH
sPCRF+7vxyQQST+hpEkGQyqVXhZZbIfqGwovJKg8dFWE6DSr+KMcDxhdAetPURJA
A61FFIL/rnF2kW/A/nTzExX6UUBrq1xi7Pt51e42EZWJzNe4JDNEQpqTYPBnEOX7
GdbdR5LWCPSvuZbcLJL5pc6cIv7/8+uhXFZGGDtJNrkMriquHKwgW2lDSV7TDwd7
9Pv+adWXQf+10uy+XmN/ei9n9j0aipAd7jwxG2ONzSCxyF0oZGHUSNNHMAvxdhAz
yfeU3YXXDp1i3dhpzJXvo14dqzDvJLzYUpqVZKQVfVt/ECkMIs6IfqTdwU0IgQbv
WovPY0yn4AFymuu5JPKZjPbJlAXxGRdjriRvpmff96/B3fCCU8wAkWT1i5fm7scP
c52SLotVtkOcEhfYoNnzD4se3dTLHirCaDaZ2uwnQ6ZSj+3ZbtNAkCxJUrUOwll8
eNcZQGOFWdsG3dgBrYQ6iiyxXfvwORRDpP1npkEnud8usDIaLpkmtHSkDZ8AxrL8
mKZlTPbCuZcZ9388LIFkP6kGPbVxPj79PoeOypL8zAMNRSFLpZI1Pnd58I7XY+DU
+9wZVt++6UtmSvo16THKgA9bLlKmRkOWEHc34bF83UcrU61r0rbRSEytTRoiCrt7
mmh02GJaj/AxiOIOBHmznV9Ta9uLjXOxMI1WfbJINC2VsdxcpT9YIZIOoM7xoM8b
sREcY/xC/m6KuztkUw7FNUYZzYQaBiFO7suyeXBwkI+o2YP0lDyn9hhCNLU8/0W3
xYDsSr+jlLB40zOahG6KJaiocZcOAooKAjXkqOOLRKCBL/anM85BN9a7M+ER4r9C
cJb3yGahL/uvH9ernHjNt276Xr9N9I7P++Z4NXlfVqauiX5c9tkb5IATOFvGwdjD
GPxySe5pqhsnu8B09w4wHetscHf5X6qxPDQ9hMMQFowQN3HIoGD3D7hprFNefCbW
Yx+L/ixfkvFFp/AaQLpVrulojrnJnw5CTwNm+/oqGSeSh5L+toyTc+2po33ppL9n
7DJ5bTVOR4Ps2GXLq2oL8wEeQ3K6GAN0TIL8uLPu2Zogx8eVbcc+0pP3i+mH6auI
ZQB3lVF4vWyWkXDjbt37zIQhQj5tPjeI1B06aBoru1jcX7v2WRgIVtYNlORYirrF
thA/mEj2wHIGSUSopo1STfmknT8XRlZ7vw5op/wZWfMjELnwGZiXupshFj39e7oO
ldloPjE5AlyM4yJuE5iYTQjWEM1hYUutEyPq3t2NxvnJDNr+8LNt+hGj08I5IvLF
2pp297gC3YQ5O9grnN8mxrW8aXtr9WZIF/7IiY3AtjXokVAI57oJapWkmngYBM3c
NUUrpwWXJ1SMVSIilbjVqwc+w4P7OWhIH2Z+zBbLIVOWhXz9CIfHGDVWMct/64rj
oGtq3KZ392ftvTkSy7D65deo5D5tSj3N5ON6PGVOrkpkeMUgfaRLDgtnunjuiQq2
JWV+fEJGLupwH264opcLCC/TOTdfbkhlm62EJUXM1QqKGB5P1kKns3WOUBZ9aBN9
CkY7l3o6UWwDnZedBj6N/y5GQ92TcKXaMz/7nFMFnX7ls7YZ0WZugZUVXEcOLqBw
4OZ6wXHD/zsv0TH8SJRVFuzKfjuSZeWZSac8LN1wCY9QbYmOhChFa2IRQoL5gYEB
E26atGNPD8XuD2bpgrD7e5EZ7uzh2l0ka88C00BfPQ6UDJF2FeenLeXihAriAe9P
Jx3QuHdJSPIPFI0mb7B5xNzliiO3FNLxfguCMUAMiWHFgctEfzny6AJP774eVKK+
QVfjCseS1duol7ck79QTaKlgnHnigIzLAG2rpqxcH07LEQaIwaP2Z8aCGUrwAskP
et7z3ITI81ykN1poioi8rlsdwbkZkm7rRBNeuZF3eFqRzSBFbHONPTyi80rOIsuJ
qDDBH4NreL1qF1wCXQqp9IJZi8xoxWme9ppAIcGwFrh6ZL+9UzsE2Gq4vRp4IHkm
iYvXmNtJRLzzKFKIXwsZUXCIHX0fFMdCI6Qsek4Rk1gmegKQPDey60kzWKPTrR3Q
jCj4K+k1QAHG+melWCWSIOC0u611tl1AsJxj/YDTAXzR+ulNdjjmjndG0eoHigCF
RYh42eyZzoMn2hvYvbzGt5nI8USN9BlzOPrWmcxxWZ4jmwynHuzB4aTM1eQ8LWSv
q6cgYFVPn1GtjgxTDfCPxrZsjvXh9DbyUPJRxLtrlXXLcL2WJtAUu3QpfBNOGQS8
Hn9V4e6K3vAg0szucP7jxzDoGgqtdHwcY03M+db7QBe77KkgXvYH+KEvEoNdLexX
6ZgoAs2Z7V7xinEkj3zKQMrEYRif09hYkY/Pp66lrNaY3/zF2KPj+Iw81T6UtU69
XWpTTb+hSV9CgOwPLyQeLDLAcHpk7HG/NVh/yoaIFCvQOKZEZhXmNkK9ZKG+N5b4
tMDvAkpk5CzgXyf8LqinZPWTfWe/UVUYHbDTFpeYBsMUPahz/J4mdVaQ+3gy8LID
EQRlXP3BjC5gh6dJXmu2Mr7q3ti6kJD8AKXe2+rfu20lrb+SQ8tdwkFbCQGJpizI
QiIFVFq8dMOb7CXNtYbuPLWVCjaDuQLPRrz4aGmnThekYHd8EmFTstjpFWDaEXFp
mvREpeRjtUidkMG4ruOTNybJMa1OVj1/2cjtcddJIYDXaDghGT0xCw1Uim6h8lko
Rsm7YioTm0URip4noNPSfr8Cg7zRp4+qnhhYJI9z00BVi/5tcGCgcE8Ib5d8J6cV
NOCH4E3Ybum0uqAF3Rdx+IF8fHf7T4PA+ftvA/QGGxlXXTC4HKqMcAbDpLGhquH2
dumkh2cmKfaliVeKClgDrRESOOYA0gYjFikQR5kcYe6ZErYnyo1cV4uES5boZeQX
beD1AuC8aLrC/w61HKHi3E1b3GZ4cDLk/rDXMs8RS8mTXQ1IP8R2DcM6HG0hQi0L
w/HP2E7MzJfzubOZaf9Nst2Y9Hs4avIXZTO8Um9pjJqc2+t9Lq+fvjuzdnAeFPjC
26DBpNc+BxlTbedf/TbOF5fJGFXi1Yf8Yy433wEsL5DWRsxm9caLePZvwuVzINho
C9vjTotvj6o0kJ1E3vctAJajPJAA3TSr0hTtWU2exMbtt9S6JePt2sDB/Hs+ykiL
TJfnIvbfs4rN8ibdHPDYRyp9d2KK90Nc0Ls6+xBAK3iBltLDaitq1SaS+FG+mXH6
1e3H0JSgNZm7NOGBBA6Ad9W87febYR0OZIzIHcSm0VDE2j5ruqtQouycwNak2kua
yAW70jmJEIfLjyRThk/MpHdaxld5YDUcPTubnFVYjmMM1uepy7QcLrx68d8kkA1l
yPcotg0RpXkgnMMs8b87jfwc3mTubKmX2TSAJevxsZIoNLFDoMGaSHdGiFRe0sxz
IG0uQ0IEhxQK0vd+MZvopZ2fTMnP6Q4WutxRCiKU3O3cZdGJBykNsIDt/dX6EGx9
GK1FWK3gaZ1eCDETpBne+qUGvsngPami+ewspozGwhf47emYs6rOVUUTgXazjZ1a
6bLeTYw0LkqIPPceOQFVQTvva48FbHUZPm+OlkeoMxtSdYbeMmia9ecJultGzwUO
tSPI90ttACFDhV1GsYQylcj6bnzCENUskw+52ETXVJXnmb8ODC0Ib2CX7Ai+w7cq
L7L9Bo0yqs5ZyV0iwFvOmYhQvQPzBR+FimiyY9BxM5d6T1mPWlGyfg/GCSnbO8fJ
berr0pQDMl7L95SGiaYPN352Ya6plQXhU0k34uAe5/LCVoVo/pYhcxYVfBMjrWVz
ktD4sU4llL5epEmfIAhtYv7Ld+vKQcmC+uex424c5py7C+k+me8vvSwJ3jxLEaOh
4031RrCgoICJgktZnthF291u65S+Wrz0CYwWHACGQ0z09dP00FZ8/wf1imMNS7Xu
fReW2ldIP1JTkf3Dnb+r4tjTfyb3Tb26ErLfZ5L+GNWN9bPCjaMXywoU2lkMdJlB
tCqGeC4vdBGNwPnp1Y/wG2XtlHuwfJt92s8LJITQNaTiWEe41EnikQa0l2D25vrK
PsvtuIGjVmySktnoAkUEHhzrpll4gcWswsWOMJuZddUIF4zeeeGdGerk1HoZcnPo
EZlQHvJ2FfrEz5b2+APxkvEbuGoHBaYXXHIRDuGiyWSQrVIt/wW4Snpat5vmeJxI
m1ro1uW8LOhBefZM8LUFKpxQoJS6iRXr+6ZiOz5ayDDUKzzQI+HNCStTCVodJVls
TfgkloA3Jcx9zYC/yeA/8nDh7VPLduNlCnnA5XzQwOgcHlmnf9aXawjf5xDOzIsv
hA8e/k2gSUr0S4dCRPFNcTYX68sH+4tPIwLAzsdFgr15Vrc5lwP05ex1T0MpaR87
jvZ8QVmcZiG4TYRYv1L8lTPNjdS/OGG22I3xcz4uS8zpiATf10RLJv8T4MI6Tdqc
3KVpcpM7gmpp5acxfeh/SA259UjBKTVaewvG4FkDBaSlmYMh2ylYnhpkHSOfuKHE
DemRkZ6xzpL9gG9Mr4Tm8KAXKyEjOu7sII5hL/shF4B/EOh2BFDWYpavNDyMKgJC
gQMGxknMGYKIQNO9jLheQhAZXrHUiW98ro8J/HMC1NIA/KVedqzjGMUxsm5YqKod
9jHEnncDvScwsbHhNaQTzHoJZiB01AdoiEBnA07ycwjb8L8B7zT23XmVz09oo8cT
NeZsv/1/tfswV3JjcESpxXtkiKHZJR4VggxTH23yrKANGlwZqOZdOAGx3CZ9BsGq
g7WR8KxYtoQi7eu4nsvkJil3uLpsOopUOK16xbVe2re5QsjAAWpwQK4/Q5m/eBWz
lVFBBqZAgTnLlkZbuLdMMYHCrZPgJT6J+QHe6rPsoU+We4WsGRySpNqEpIQv4cW/
/E00xE3oY9TeL4cXkhX+ImtBOFfA5c6uL15ujQvpQw7v3ijAGwkOnfc3AvAGQ+ya
gMwN0wRmWFkl/Er2T7IHFQE8PldJHSglOjExVHSwXREdNyhfjFZkI1plAmD2U8Dq
0j1q5fTbbG+81+6BBQ200fT1y1h5Q3ry7X48vriai8TOXP425cFXickLaiczxKlO
d4noo1DZSiPcbZUWgXhvwTlDv5v4METEQZ6/JwZbyid8ugNLat3frqAL3jhUd20z
PkK7vNeHydtKnTlDjq7ASwG4eBHwSjmH9JPBtxdGuoLq3V5O8OtFAohgD8JIwPES
mttoxJ2lPHIfnd7RMlapR1Hpm83/M00TyK8D/xwN3ldmQRfC5xSVjRDBDqtIrPrf
NEo3KbmUafBmHwrZyctuLUFLdToiZI7OipWhDX//ytINd9mYKIjPEZ8ty7ZB3Xl3
N8wVoSUxWzTbxkrGC+VcU9w6hV7SCCd/0HqAe0ntsZnP0JYjHn3cG1QUFLGavZPu
7vd3y8x0+THX5uofxPnkBVus29wubepzQ9unvqZ0E8TPc/Vvp2AqSdTVTAr9SuBb
G90z1/R86/Q5cVJOJKIcm8VddAFM/EwSHOVSiSbDQ3EzwDIlJIAje1dfyOb9xoRj
gqj560Bu6tr1Dg9WQqRIqQvEC2q9l+wijxET6RKIlt19l0LeU1kWPf1HwSGP8vZw
kme+dAu1Z9jQY/oQhX+wA/zvgZOryWdPN+MJH9sg5xOGPoukQ7X8B//LLNTdJ/oJ
IXQBq7z6Vx6M4pjtJpAMvG9z32UK8AsJ/LYZ8XJ9GB4sfItat1u6FWqPNGo861Fd
RYBWtJrWyLM7Io1uzxZmpea8dBe2fcDl7jKGrAG7kd3FYnmWzY9ysaE0AqsnbzHG
+WBT2UReastT8VX0NbC/ljoSCBdWbJP+8Ak3kaF0jYilVSNK71avs71YmcNiya8j
vjvm5GxcYwOrBSAzfXuXO0shUUbbVr5oGxehhmYo6+7rIf6V7OItd5z1KVZneI+o
9TMKEpXZcDcUB03KSEb9DlSbnkumqNlIVeISlR+V45IzUgbuwKuulcNcQBnApMwn
amEU/+/YMJ/igPKVvVb+lgZl1xz8KzrV/eNooVOsoLDZTV8b91wZBxXTUA+xCmvU
AEfZ9clqCS/Wmqc0PHjGrk5Xnm7vMIpCG4uVHLDC934AwrxmoQ5SNBe+U8+VhW6Q
WRFAJ+v/UXjBf2q6AgWxlpXtCCOJ868Nl4KeVIRj4L/OM4HrSHqNPikmaBu5FkPs
toZgYYPVOGH1NWA28frS/yQQ12U60GYyMezAdJCX/YpZ0ms7n6nT0Scs+RuzrIrF
VaA2LTB3ZUe1bDniIIUjlIYPgq8Q2cEbkdI8Xr1x3DLClCtLqexfZCIyLUpV3DO2
tIIXkLi7pFjOSE4N+vaXq5SKooMa2YfI5b7jpRgHcFUdt9O7jKVe5dPSz9aPqydl
t3FIxLIkUVlVQnDEud62fYu/X1R13MQ71qowxbR1z16ciu+dvOsOnScwfeLeBjY2
tl8Mh1jvuaLMzoRooFnC5FeLAOI+73tHtbpExUGHAEVENWMcB7pB+AB4ie72tQLK
cb+9k8Snx9WUQLnYfVC2eukUDejNVIL3diMQaF4dED+52PmkG2t6r+BdJ101Mh91
wwQ1Y1ez/cqOUMMSwA+okLmnakg3Y/UjmEzb0vFFUyOew4qj6hqBX+ylTsSudGFq
/PiXvoY2ovhaxv6JfN2gx8QrgutFoM4BAhauHgsizsTa3Fh3f6VbEDXmIOqDN3D3
ST5y21MBJyiiMUeTDjTD54WnmeR+57VxYZPH7e8PqXzvCNUNk/0bKJIrem+4Goq9
53pedPTgCxMddaXkL9Y0CuEM4m6yoO670QtHPoQjcgc1UVz594zjj5+tHQuV+olu
qq4L9XV3mEieSk/mZq5uGWCmt4/g6++7PEYp1D/L1LBkSFlEX5n/J4cz8Xy90qK4
JqvfJcxXM9JfNH6tLo1h3iyuAjHoh46+wdVIuffFSztQuw80nFOVGg7NjYKEAute
yvOlAJtELnXkkmgrmzjni5QmSuFlMIcWcnlrG8LNaj8m5rn3O5mkDzbiSdns4v4p
//45CnG/8IM11vUspzu1hq5rcbEjinb3UVugGZQzY4KxP1mAd2eSxg4UyRoBUY6e
IBM6BBInc1n4BWQX8k+k4GJldzlaeB3gIEbebn9gLfk3iAGtcA/DD6x/XEasS681
qH+1nRhxL8xmLP9dUaiqql+sFikKJI84apCLd8xp7F6HxOwSl5D9mxra6N4QpIc+
9jslekEOFTs1vC7mGu3q5sPfLRr4UhndB4lf8pCF6IbhEgvQzqYpkp7dIrbXrbhS
LEJQYn1zSPlvPLm5VUOyqMhzeslq2T3LkjMcuu84BK0ZUvhfiC6ncO3Y2ncDgJy/
NP/5L6gO4WJjcWZ9lhTLVt8KRSLSCwwGrprWyyXJID+7dZCIBOVIPnU5wdsoGt3H
nC2Pn7A/LNrLnCV0hrOyujKCgl8CJNUrbrrRak0xav5T64u5SXisZR3waa+4vUNY
S+6vqrDAVa8xCzsB0to4lncuoQbAYjP7YnSSxpiZ5Y8Q1nNgHu+FY6nmc6w8i78u
mEof+AqQhg7Cmvk76WtEBm1B3IWcjurkInmlF/BTyJHSH33fJn8/mw+uxrvAp6ug
d6zrY7xxiVyOglPu22phY7tmQee3QayR/qqyQ+SPr77t6yBCFN0Z3vj1O33bhiQh
spsVJHI72311otPL1NUZzGR0m+Eu+uBQaM2H8P0wYL32ProwAq6XgzDJk70svL8s
BRg7wRAFKB+kDpC9Dr2SMIpJ6WSpwFrLceiOBMMYlR1M+VZ0/IrNEUZKGS0U9fUc
w+kubeQyyxKxpX59s3XfU1ykpx3halo6WgHiDyKm2yBWWIbuOHvO3fO8a4m2EH45
5tXucmHprsuvLtcONvUvul7cwhKnVB32kp1aAjdW8XxRInHRe2D4K2PMuQJ2aoJ+
HiEV6h/0fJfnVgB+V55sHyTSW4MI/AoEi7AfQq9f/H9bS3rS+rzvxT3tkBrEK+IB
TShizklSAxE90L/nAodvr7SoKR6cPbjexkh/L7YXbRgvoZmVO6J1VXcpJA/USiSd
MS/PezabIXiHaOpAqFK/kVy15Q3UlKY6+bUCvmUwggqFW6/6w6Wr5pG/n7TXjOTQ
htLd7UNb9CUvTJL1f/2FNYw/wkpM3hwOmeyvDklhd7P/bYAbMpp+m31/SEshGPs2
t25tUqf9TwV+ryB2vybLbLmxfQF45I2DOWo53+YelvOPhddAbYEaibe6h1zafWvS
Mm+jg7nHvC2AoXD/G8u7Sz6cww4IHLR3hvLqytaO6NkrzPCeWAJc65X5+LqYsGxb
YAnpMc4aF5dgj4ni8Wfu/7voVrDXc8v8Z4CAnnuXze6GfGdG7U610Sn0iEJlikYa
womYDRyuuLAFguIZVdFjjaQJwGVbJZrbLi4/C5b2IL/99TqwimQRDRsgX3XsA2cK
HIx+RtHtn8M1ePZrbDaTLlhBN+R6K1N/p7slzdCFIlIVf+PSlIzgml/+qluhdXDF
+sPxwzaRqTb7oFHJ+oU+p/gZ6rzvxb+pDon8rQjCcaB28ykrI/BmQmR5imfUJopS
NbPrkwvg1opjWEqNqK8j3D/5pTDuyY4HCZKHXhqst5U63XtSCS9ZkuFXVkKBINVV
VwA9So1/WtDOnQ/rYm+90+APeuuT2/E6GEnujmozUtSd6yvwqBdzPsZb3OGJrGzw
bCpQkf7DeWDoo8Pz+hc2kdULL3Plidnm7uXSY7cnyAApuMqx3uOPpm94jfArIQZy
l6fInBxHxEEG6BmpZc0aom9hcwquqKNF1FxsYSrOTDh3z3Xj5CkB/TvzKX/64qCo
jsA4Q3LaHBUHB+L6SHgXFi4zWiZ4duQOz8vYZgqSBHGzCysvqiOy3+PCCP/8dnVb
VqZfroRTRkjfUomicIWGXfCDqlVFk4XNGPIU+9+UR9tRcAE9Z+mjt8onc5P9A/WH
O2/XBJcqbeo7EXBWTpT7bMqXZIg1fdhCS0AiAi/qD+YtBwieZHgANkTYUSMkIdnj
rERFSqrBOczyz7QV2UO2TfJY4KD0FVwarfc0TQy8I0XG66IW7Kr1qv28n3/OPmjj
KHYkS43GTn7b8KakPy3prJlW5fQ9+Qc+W/AXySsZJGOh+FQp7UzGVDwwSc+UO4Vb
WJ4N5yUXOzQSzne8UFa9MSZmfXyb+9rpaWWwCGdGQ7tNc3N2O9vGau4eOr602rKI
XievT+OXLKYNqJIJqvkdE9GuTS6hexdeF7Hnjr5ZYVSXoVh3eskOtd251qK6uQYI
lSeD/kpwDqt0Jnl4cjrhjJPud7hl/k4dc9p8tLy91AL8+hL4ZV9G6syOVgt5e5pe
PX6HUnGD9CxnjBkaCXSFM0QJZCbMUX+ieX6ndVh9wNz9djUJq6aphcLuuDDS9FYm
0p8QIkGvMafIYCFCQrYPc5DK6i9xNyqz9iEjkQOEKFN/UwUIi4gcT3XUFPLT8sre
AiAsFtdO/8vDzLp8Tmd93tAYGXSuNvwVMTLZK98S7uGFNq9Ov+6jgifZvyllEA2R
7C1XTyxFnleC9QwHIPVizHU+3oX5U+2pRCbdlKzy00hK8qm1zTm1WYJqAgr581Nw
LvwzXjr3I5gcDFBux0RPYsP+fqEAAM4j1aOHJBAbzM7XI47zyUAp2fRR57Mr8WNL
IvRWVlW8rBDrpjNlJpMG3d6kObyIR0dWPOVvBS4t5uJTx/4sZX/dRFj1LBVWpqxl
S2kYvEH00UllXJdBgiOQtfJmiXTfuEtQ33nFSFNWYfjWZnDrg0V20NHZOibf7S+w
jMyEfXtL2kx9yEaTldnPfpV9zmZLZN6+Fwsru76mVMDCncJ9KQZEk/36k6Bn/9QS
j9nrHSVm/t5d8UeqLL7lJCNB+7nCrnMXaazxTH0JP/AoliL1h6+Or5oxU6NY00aC
uAp9gXiBRqNWxrKeLRzjOiqTk0+4s989YRqjNGdrEEhv89xf3Jf8/MSCZDcL+SSa
u9L0FTBYsk+OxKW5MSIQHfge+I5QbdG8vRl+FsK/5K/65BCId32PqLgkifACL3U2
bVZ7fsZxUFP7l7ZKEwJgjNQPRS850wUJo3r0vH1nFv+Y/dqfaBBoI8MqKmStCmJP
mInorZhivBJqibspBvnwoUQZ52tkZ1It3Yb7jeZpNTQ1WiCDUKZ5UdB3q/J4JpAk
VdLtYsEDc+ZpyWe0nLkim502LmiYwnNZP8mLYOi+TywE1nkRHPN1VZmpkzwZcB87
r6+DS4PN4e0j42yfG6SdIIafCggSWelXj0POUT0C6nWi18dp0+jjW3xtb3uj64As
xCc0Bb8kvjtuxaQaW18kRs/wKAiroarZDe8p61sXKNqpuS1/qpAYN8it5XGfXYTN
3qOZ4CsaUikPALteNnNyPlwz1PbGEX+mBUw1hi6O1m966PRD191gP1GUaFEjfilq
+YdgfIH1jrzj18yWWrExiPpjawMJIugwIzuQTEKdbmvEn37IbJYVu+I4RhR/Dq/n
qG6772YZwpSycxNKCY1Xif3xAvnWD7HEdNJrADdnIoyHyCx4sY7TsfxgNls+nDzT
sRrcBTTT4vgX7IppcTx3IL6zYeucAJaItZF2Ul75gCC6IHGJLJxsElcePTl7Rhah
P5PvWdBDBbggmqVHLc2aGGIi/kscospeeFiL9AW+a3cl0vz7Ra1aYyCkOF0qJj0W
9+lkqahG75i4HsOnXN3DCQyPJvuu9w/eqndvIM31Zg/ac3b3BYe+Ej4eFSv8avE4
m7/M3oLYUrWAxoqIyxiZ88a0ZbnQ3adsK7+HQmb6zM7dD0ef8GFJZ4xZQI/24sNr
IPHWt367ejY+99jd8u4nhzO0yl7A+Jea8vKVqKMczHdRnyc1hnK79gazzn947QPU
HK87r86aba8wrINF0nkcAtfCIx9wSNarkgYTivUgCDtCpDPl9qo+GD+wwOrOZzz5
q4hIYMk2SXvW3HJXzx7Bcnzk+HoM1DV7zjFVPbY9KRo3QV7j9saTirgSQWWcJ50N
2PNuxmc/+7AS692dA2h55E0gZD38wgPTOv64VXBTQPVby61poID421zOqzAymH+d
K9CoGZxroApk1vzXewhkp7L2UPZ8HiTpJppxyjYBkSWMfOW4VRf2pUgKWK54Itta
1pUWZoxghoYlKTQ0KCzOn8pQkNWM/qrZ3cyrEH+8jlE1g4PWE+YL/dAX/CF1F0OY
DyJkvdlDHA4Q+ZiT7+tb+DY8JTetmeXMAX+7X4CvV2RkyaRXV6/0TdStUUHt5Sci
TM7zYoP7q/kYfKlsEekS++Qa9BWJQxxhQ+JrIpX20DytqOBJr4JBEbte0j1c5mir
RS/E7mhMOJ01vx784dHOZEm6VPbo+PGcL8j9hzo0D6rzLmyq+JqTCZumcL/s4WrI
K3HrBoFpheGeOqlftUV+dWJ1bKcwJBCe6DIg4ujdWwJAUctvXiCmOOPne812MNb1
oTTVwKHapZ+7Cch8TrAOqisqM7Oh0MbfMUjvjxUXGBE6CfDxDp6vXa9j66o3s2ck
DycJE+MSli+KzvP2uRKmLkW4YDpb+fiI2j4kO9LpCPhNG+UUyN7Dh5Wc37RCJSex
Kxo8qEVBy2swZk3fClPCwwiGX0xCI/HEKDN4FrHKPvxjEFTO/LcaxUt65eYrUnFC
3TbqBoeKD3tgoteOEecv7xiHn7sip5tu0pgqzRSHp0/gRLvY4BkgqvUSDBoKQLPk
mbDemD4ayPj7+ITz8eWq0MnLv7JHkPw2hrgRCuII2oxYKLwt1KJcn9C6V4ST6av8
L9mO+vYUiF3qzKxF/uIjEO1FJ7ewvr4U+n2I+4AwCM9Fyb8HUYlTCg4k2WkyVxZp
4N6PwixRLC00GAXmqAiRbeF88vHJZ3sQuLMYTyLgB2O+6U4PFUjiiadhglGiUOEJ
3zn44E37rh0xqFwrw3qRFaygsqPFOk9O7iQ/sYBzUBfKTal6gJZ4lYiFqFAq+zPE
9LE98ClnPbDgIPkMNRusqYb50ddHgdKoIR3I5imB94ijmpUGwyiux+hmLhoUQ6Dw
e4fAKvH5mW/QC38hZE8XEr3YvDM5zYOHcGOJZWuk6OJ6gMfG+Iq9BVXqc1fVK0LD
6GYPnqlGvnbTGyJa8BfeAHVbCP7KQUs1yN4aiJ4VyD0BP37W9TrOYfTn6aoVCKZT
pURuZhi6AmDovhwIfkgqkY7y1iHVi5h+F2YWz1PNmzG/OznYtlW3kZ8y/xjF6nIt
SpK5+TyoMuXoy+Bssoensc5KgkkE0pUYOIsGlQ/i3fHdx8PXCNEUpXL1mxyqSxzE
g95ahnJQ3nGyJZhzohpAfNjRoaoLPTgkVkl0fYUAs9PPqLEPofWiFWXg+TwlUHjM
2wYnukOJ3crsV10ZFs3HUS5yYOgGbBrVpYRVsRRdgoci84BdEBSqfToEuQB1eZ4E
e8ZGt6ztUz6NggplWjYuiKI/UsieybWEIibYHr8MCjmE8uldMJkgBAWdNzZA7lr0
0OQZVZmw5WN7q+0g7Ivcyr4qff35y1yxr3fSqNIXyKuEWsJGLz24Fp8DdhqBV0v+
zxc2cidSiH8PaAcG6LCK+9ilMHDQocJKOLuFMYtpaGMIRpOEUDDMbfppieLRI5pQ
LIhhOMg271oCwgUvF/DtE571vLtTT27Fm4ViF8dhj7GQAPbKxVJYnKE4ZwNNyfdR
hV0OOHHhsfWCuMdeDzYWKjlXaBeYavkkxwjNmYLp7Q46G/GqLy12y3sc7NNiqdxF
sv7yVixoBuNN9tZtR34sKuTsuKfCqyofT0qNaALmVXJA2K+m9Xi7vFTvzK0vpRCZ
JZUZgSyo2jxS0wPmUXtAn8hyNXHs45LEOoa6XB+kvzEb6VgLUZH/GLNDUSjQ33CT
hXCYYlPjswW8gD3AAyiBGUMeaiWG/HRHxPv03wg+4zTpTCQ7UzJ2iD7tu0h3PimU
ZGE+b3FWoDfuObTZsakLbR/9SDuH/xYi+5Y53Fmxe7stuiiGWg6PMEguxmDXKmKX
0ZAwZOKScnGLWf/3+LnDllI+8Wc8ldq3JWpEbdV9w3VxzUSr3Y2guTK4hz9sDQ5W
VM/qlYDFdBtH//u3EgCsn6UsjVnG6niuCCXFO3i9aIell4G8rlZ5xhMscPL5YeAc
mQazzlSoLllj+sP3vb8jIFRRam/I1nNzYUAg/MpvkctLzr+jsvNesnos0Y9n36Sa
XrOl5UqagDjJ4z0WBs9vb8OyBRzOIyFDnvYCCyAWjy37R3Ydfuc30KCHPTQ+SLQI
JzT1GqX6KIsEi1n59F+ZkGSdIWMbArR7gqrIj/FqcgGlO9ZxRApkYfSo94PFZijb
dqQIfyK5Mkjk+fhrrTWP+rY8vhzIkBVRwcRUAvvcxXG4LV8JLOHlIhaIlay/ZBqY
WNA4qFxVMJ2PfKEJprcqOoNSlRhXMjLYf+J+MuW1zyx3HJWDm6rkBLU7R2HoC3E3
t6jZ9GMUcHsAsyFZKGdvmb1G70lQFW7tompNDmaG/8Fe12ye/ViGKOVGWWf8UCeb
J9MQz0CUQoRwo+tp/kMRupqyeYQkgMQIYZ+BgMRJAs9iAEGech9L9sK1u8fGHSps
kSXXg9/pUTkazhwB8B6jYVRge9H98bp5fovPSgUrvSzprxng7r/LsOD8XLmdycQ2
qeQT3nDE270JNqDdhxeo/3iIb77Djd1lLKRvJxrwPrzrkrsDT/5uQaDr7TFs56z0
G7pP+TxhhhCw70hhl29I7fa01fC+xINpbUhmTD58VYWsKGqAPAIuHvYKl89PtCZi
RP8slucIbe2TOYxjqb7nhVTUGNT/x5g47meUa3LP7l2Qg0JKz2/yjgBRaA+7alge
WDqwoKcsB58DUSQ9+qNLuw==
`protect end_protected