`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
j9eMmSPGcKCWAR9PvkqZ1R001FU8QKTyJzFqNLn+qur6INyYDE1AI8LWcxAzfnTc
IpZG7ua3uuk5/kQKKQx8ZIPLfmv6H3t3eWjki8YIAtY/d5E7Gq8Z5mNxMYRzGGTg
TCMm6oOrOTVYlCXHE0X9AW696Z7UGfWirVibl8hs19hrFdeZKGiGht4r09vHR+Gl
FQQmSObM5aSK5wu5KOrK5ZUKGHyBhjnIQO5NnittDjOwxV/57nHVg0pdG6JUqyvm
tEgmCY36RCMRGWN7sekPtNHjqpZkmYrVX1T9QF3h73+8ZekZYd2xY2hpHHGYYeWA
t3+Fmb/6NUmoP8+Pt2hI6g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="wX+NBVcG/A5ruHK3pkDqG8ZVPdOz9TJPJ5saXZYSeQ4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
j/hqWUoxjK88VtH4QmjIrexFOSwtsLKOZ/LCP4cmrqgzmR/e71apdtoL+o8nlfy6
eZxDZMmrZmJGoazz2oK6kz7xJU85UCwNc4cxAsVxNdCP19vZxph/nCYZQ9lUFkLH
uLBkOeFP15CD3jG5/dp945fHP13J9SzB/L9PWvDC/gY=
`protect rights_digest_method = "sha256"
`protect end_toolblock="sqDZkaglKf+bDjC7VKm3lOELrT2Jlynh4UhPg2J0Q70="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 27696 )
`protect data_block
f9kZDbPp4NLiAOFOgATj9W35i3s4a7wbt9jeHjHVcJxMoXY8rb8laqS5bNUhXGW/
MOc7UNc1VwolqhkS7G27SLamkGClZZtXSbRcN1N+5kYdRMAqEGt4OHQHIKzxxfMM
am5VnrC5dYupkSoW9hEBkE9xNIzdEPQIb5M1hQWWHoxKj63M6OxQLFcx/7fxPFdL
V2YMgsR3CWO9wATV/LXYJse1NN8TToPt3qrjP1sMOA3aImp4YO3pRBr7HfdwjaZT
ed1LgfWd/itwl0FNxJRXemDycLG+MyJzcnHjWuKD0t14kixiFS6YnE3vWi1hBM7z
0WbcCROTcKyH7nqr95mIWw5qHhL7lrKv0cQ4j0lkpyAWur55OuXzpjfUfufUEnEa
JdvB2Tf0/ILjmBDVDKo8h4Df1mb6jKBqEbTuakTVeFIcdbQ+TneTKeV90Sf/d+xH
i/BFkXdOAjZDmHJVbIkxaYeuO4dfL+WuUKXeXD1sNmyMAqmfNpl6MCnRcdaS7XdS
3ywGfMvVRLpRi5QsxYDWREDR2Cq1ebHCQ8oJszURNAjeH2JyYTUGaGG3EZr+dink
sp61JG0xBx6ciRkVqeHL4bbR6jIO6/3JrG4sM5DuiRJGq3RaQn23JLJ2ZOUJAPXj
JCwtjsdTVJ6LFnGu2Alg7AZc31Ih7Ng8z+lXeaLRse1/TCAh3BdmBeE8sYyRhc7/
FEKM3RgZYf3AdrwAiaPS3CsWJQ3rxZdLdPPMHHcfX+G9fnW0+bbAm+fET8GxuhWL
R74CcWg3762OFb3xQ3MJuq4f5po/qthdG1ds+AgoZPqC8JqJEiWhO3r1BqhSQeXU
gKEeJ5lpNYOOdc1HoLdNbvwekFFUEa2gfozi2vL1wcbVW3G15zHpHbHmWCoU3rk8
t8MSd8qr50jEdihR3tsoOhWv/wmFXca14zh5dxgYpGnv3Dw2FMLQEyXinWpPluuJ
pGGA8Bnkrf5Pa9xVVptwwtNKAH2K/wmvjhokgr1vUDFPmuewdwnnwyov/ysqs2U+
uLYy3REUx4AnUurQgLjBrKCM3Y0A97Ds2dH08zqerNaVXa6eGwljyr07XErF87bA
hbZSKGC2dGQ4CgzfzJ4knnpnPfkk0MtqRZ4SBUt6U6y8j5l8mVQth3dTgcpGDFn6
WJx6AwspLCPQbIOIxQ0MTpgARfvmxYIvMHWr/eZxB5mnD7s3y/aVY3RFoFFocqvH
9Gp95LT0fse050+NTa6uvJl1S78gytCbtOGGHG7IQHxfwDILZPjuzPZw8mdSrr/0
2Cf6k2lB/y4u6oWjGoTaKkQEiaeShWfzqigeM+uUbU/m6GreC+KxtOHmEFrAP0DO
/llnWnqU314qHsUXuryk1Tbxvcep/YJNRhS5k/CuBtkCT6iJGfMbn6Ianq6GxE2g
nkFwsNdlEeFyRnE4QmBFU7hxgqNX7rIqTuWQNhuKCBF4iWv3Rhg8967ZuED6pYLu
y5+0RZ1zU+aLdiJ1pLseSvmECK59yKrFS/V6dqrkfGEt/fBdv5ZzH8gv55Lt+zsH
XOhpd/VmYfaWuGb/pN6GujHNpkNbxXobuh9nTnhiHhSsisBfWnPtBi9w1HxF+2Os
O+EvtY7T6KqzOfjkjNt7k1+jQbm+PfI4+aMthVVpVJK/+CVbUPNB/bH7Ge16RSxu
dYS5H7EhzNRhfLXDto/l5t3Dz63BPK//84yVsG5yfuYHA5nBX6rHwvJPIHtcZOYg
5GM7Ux7SAXxbBuxWR3k1Hp0GMgXC+23zFw6Kb6gWYatfHsYpzQNt/PCljEtB9fSs
Qn8wdoPFeeIjyEpkDN8jAT56Eu59/uZnwFe0G0/gg6cSVTV8SNBdhAEYHqx3U8e/
jS1DrMeMTOCsx0zf0dF0r56sCiw0ptK/kLGXgKBFwEwKBZcKfwTWBJ4jva/MlDnJ
Ms6CJU47OnW6JBC8Mk3PgJMkiLbMf1C7rvkPCfhzWjAPamQAwmQAdefBalAKPwDg
i5IptkzrTvbVX3tqOW6nf6MFW6Bw2eZzUyKl4JgWEbtW2301UW5WnaIVgBlDPrFM
hirTpiOPALP5q3opX7N7fTQKq7DVT9cLPbpmKs8Np1SV+9PoilDH7uteR8pA7r/X
+nAAOxJQElTUtikqHIBY706a8HwXnV+Jj5uLjBvhqBMhKpuhAz36kdXZdoKXx7DW
YCaDAy6Ep5fmEcwr/uUsm8k1xh/7ShMZqKHGK9d2OEt/oqJ0ji23dUdwGiKQvkLW
t8LdBMJ6Ae0CUL4ip0Mch2mp8HRo0Thg6xgWKve3KwUUzYev8vr2GjazTj2340bP
eMfMaJvz+0YhFvkfOYsycsojgS0H34M5a+0diHz7jTuxhSUr/7Hdyb8kGbwr0dge
I4+1FIDedhkL36ISAUXQd8Je4GXGPST0tpQ1tUceGs/gonaIxZQ6wP9UuDPw4kTe
Ai3QwuBP0yT8s5tNUdY6F1/KYCgGcd+LGyWTCy2H8RBYFGaI6KdxQHVEQKG96mDL
XbYHrrOM2qf1OlvGBc+gENoXW3wC3BrTfBB8MbK9bhh1T72lPXOaOoL0ik9orGDH
YxpvRWNPYqQFAKf4Ni0yxInm4O9knq1wHpuS08JWpyYZqtLheWc/IrCCwpjICAv6
owePSQp+mjeaxTgH9l/YUEGfCbyjmN07vMpkTC/L8X7cdJhzxwR439mvFeST3fMZ
iGO0vUnZ75IVZnSVgEy+dGNWn+pVVnsndlDQFbQj9NVvF3XJR9bmxBz1plMZhG+J
ApNIFYvFq/zvMB0WpITURePRvgM4Riwzwj/JG8rZM31MIXE8r7UaaZERBY4YXrxY
TM4oVZ3W1yJc2X0RMjnJpzUdTyk0r3pMZMpdS+wRrZrnnv796y9W0FQLgsPQAGC8
T+RZjmj3WSDwVR09PTsx+GNSKJuJFOH/LB6j6HOuvx2maU/ZH7BDxi6zCfN0pTEk
dZ6t3zb5WZ34Bi9kFy5eQsou/uqPc2I7jrWShATeZucJa6E7LlmvilPsQe1EGnuv
P7rpfFV1CDMHpoFPb5rmG6rcRZp5JRIKrJQCuuMIKoSoDohQ3hDf9JGLCPBOs+lp
nwSFW3vi0mpUByO5kpNxx4lkBLUVlbq9UH6qVJ0fYEcB34Cj0di0YEJuoBnjhq4Q
vtASnYClA+23f1UIQNfkA1FvXdW8Iy7alY7BdS7tLChg1lulQi2rAG24gMK7f8hm
hv7Veo7NPIhv1bW373r/6hDEeLVXEoBiEMLqckOBoQ/ztrC+5DpbwxCXRGOj0+Bo
skIZUk/6RARASgH7QZGFIa1MW02SEWMQnoTqDyiPI84ryP3MC6kasuIsfVv8c1A3
JjVVgIq0RpfpK4ExUfYyVc62OrtYJSyl58onxfN3lr7vHGEEXpTWp/lb9Tfze6a0
ImRDGAvRTI3oN4sOpvEJm1Ud6c6NVu52FgSrx1PzN2k+jEpWBKT7dZp2WDawJN+U
Je6SZe8em6NbWt2sxFyznFWftCot4y8DQ1gfOFppFixY6+rsgP/EET3wDFCSFScu
BFf99udLb5la+5fD2xW3mbdRC07b/s+Netvqa6CThFwHDt2lt1yB+uz26sHejUvp
5WcM2fyKCNRc8Kv19fdbV9QkOv4NcZrD+hlYFEBSp6wsgIcXYKc2e67Gx269q9w/
zfIzYUD/Czufj3atSD+6ncYyHtRG4/Sn/pHLlbpQ4sBdF9/dijGBkVs2NBvh7Lge
l/XsP4SpDNa7j9hzxGMMkcX+JuDoKFCbx1PUvHw5jAUCsCmJ0EeALKasL6VQQtre
Iukc1kWSnD37tpgwXJdpzVh9GFrsO5/T2OlqNJcSxYgYwUeFmyvaR4dzPxGoTmvu
wZEiVNuA2Qb0ISrYnOXQsCqxtJQEsgPPCnDbsZ+hloob3sYbO1p4XSzh9V75JN5Q
TmrY0fTOCrG7SGtaCRWcFW3VFf+Jn0uApRynRsSnbs4rIbYRSro7+EAzlKcnJiei
SWmdImBhLhDYPXmtvNFQM8Re69MftFG801L0rot3wLFL2P/khTKhAtb3fBEYpjLh
2IXc7h7jzpCQ6uyRTw+1b/0DeSUTFlJ8qqyroShcD4C+bn9qCTVhPG+njcnhOZls
jtPMZPxJWw1tPVgMFeK71F9pPNCzYqCArbFu6J/lTWem7CAPQqXeMIO35XUAKmQ4
TwJ5BuEa1B2+CQ/id2yhU1bfRAU6fz3Yfr2z28nU4msyK9fdvvrdrQgLMB9gLjTp
znuib9z9JnkJpMAXSNyrpFf5w7gi+i2CjtXVP54gOuc0rzqCc5DE5Xpg4geakmIr
4ld0bryzGCZw/NeJ8Vjspo3x4c5UyxvKyiNDgNHj/9IZOiXy4LFkRvzaqKkDjA96
9UZBmbK9ShCHflu4gRDRAoJmbPxamPNOOe0fBE9W56/B/FH7Lrt4/tb4ZiMWZEvf
lbduaZehMeCvwf27Dy4WbS4vPP1vrymY9LG0Csfp8V35NMwh2x2v2C0fDeGK2cjv
E7P0PovEnkkN/Fgtz7/+4EL97LUPwRyk1krO4247tzUUoWu5DPGC+C9Q3Ue59E4T
AMiwDNDsMLhsl4ER2NmE8MrtqjOlbV9GCuEhG8/ZLwLMUnSrxGkylcjIr4qqgRdg
G2zG0Bxl9dLCl3ecfQnF+GMI/NGEr+6VF9IbkZNGUOtCVuAV+7gr/EEDkJFqr6Dt
BJSfY4ujv9x7fCA3eqEcGxOnDnTBEBW1zCBWRTgcU/MJ/opJ7vvZG72ha1IdqHRM
fU+fUdBTUoR0RiMBXCp5zp1aanpqE5COMnmHwKIW3hfzydWX5Dk/HF2vhMGo6NgW
E1TGK5TkJxHexZmShMvuK4nIs1dbPj6nv36+Qtb9S/W8O16psSh5xecEaePj7GCv
Qt9b5YdN+WIIwhqpT7I52kr/dG1a+L8ADDayKfoA0Tkcu3BFxUt2xL4q+MEzfoo0
vHkCsfjp51fgOdFjcEJLqRlgduuu8bt8l6G/tgvFnCKWp2Ur3KPkAE3XBPDihdat
z2C4fmYRZ8sTzpB1SwaAWXkfGlvoEBQM/m2btKoBq5wOTOxeccBnQe/nnD304t4T
8O1nnRYQIZUsRK9Azl2p6Gg1kKtyqYOwgATvl3piupXbw/Z6YqxLr6BZS+jr+Z8+
bptkxQzQQJZ2mtUKdeugt+nR9HhE9nE2WcEJMzvpG1nswDIU5RsZqDdzXjoYYsUm
T6ciepy6mdheRn4eJ6iQKtl550Swqb34A/7BHjM97lNv53F86k71EsnA0tP1pn7S
Yvj2cf1Dm3Md7qpCDVeznV+2Wb3eSXuzGwpvU1t2LSBIyTd4MrO7QHehMoRjLtSu
vKTi0hFY3rdMK2H3sGPMA1gHurgL17vrNWtYXgXF/waKnEKJCfCtndPhs5VLd/TG
jzPJ6D3MdT5KUED4I+Hmeyt7URckU6EFNK2TAuPbsgXWZHKTMnCqzm6o3M3KRmB3
vYVbabssTasR6P3q/MT46oJp0p/hCKMQiEwR+V92v3VHrqikvfjB1k2ugqBNnT+s
IUhJxLMAK6khtKdHGaBPO9jOEXmOXhgIh2tDFYaO80htoWLhbMupa5znHQS3S0WE
ksaXS0E2XKkEeUPzQVKQkT3KLRWElKOw/HQH3UAyV9w7VLSbOrojGzHc0paQAqsY
/UqGm/GR8VXK1SlwvogFMrtriBooHGVibJ9C2Mh0VWnhWRdYPMDt7JzbclSU0v2O
zFjXeolaE7miRZcSIiCJFN/rR2vlIZPcUxqLXdcne8uGCgoFqvNkTClN7CyzFAHA
Fp4JHKGEWQllwczlKTH9WTzlFDs5HmA4XT/L7BNDGX0jsIHooXa6RfmfKmFWMe39
Qp1PSfuPFsbzl9Ru0PUFxSh/8wt7jaGrlmff1tOoQEnEZ8AqEA+x1yi/tpwRqAvo
uHDwVuNmF9bi6wiPJqlWtbZ5NBU0ZEHnTUtHdMRkn1zSzCZfYI0m+3Jkl14fQXhl
TQWcFmfih8I/JDbYVbu2o/pFHwRsmex6IDtnpk6BF+uIcVo0e0XM8ckv6I1gCnJl
CK2/WvtP8U0H1ldcYl1nvcg+2vI2gACuUOKGOMpH0X8fQOglPIHPiGXibk7oyRuN
j08+VW2chnPx/65Pi2WLQDUQ21z+vQ4edH8y8v7sTrUJ1LeysLDiOmcmrISX40la
kNZuS844Ivs5YL98Zat9MZlE8yapzz3Vkxb3g0ND1NKQGCCRwXXNzQruXn0gDZWU
VGAYuNQnsnc2pZxF8lhbt1H9Rz++Oj9/7OjxtmOb7YfF5wi4r/8SMLMaNgXwFIjN
Z1nd08sAo6a44dyz2j0vrrib7drEhVJcwCvARkQHnAWGed2csVqxrkSVcBpwXPb6
cK4aPGv8pvbpdIsKrw+C9Zpm0Byrdufz/K63wkO0XAKxL8K11V/KFkVA7MHKtFtB
705bNFlBA1lzl2BgGXV1fZq4L2FdlusyRCV4xlh6sLll5wYUZBvrfK8h7SusrLfF
qilhPUrFmFr3fRs7ZNkocVdvn/gJIYIyFOLtprtDhfjmIlJIAkKyNcTRBzh8rGHV
yTLZ9IjUMzOKU5fy5WoN/Xdl0Vz8Ygz9K7t0cFMeD8qXXKuLRnj7SHo7zKGC4rm3
j+0U540t1ieqyGgkfdrw69yJiOOibahligkx8G/wVYfDGcsQzVj6w/Sqx10za+BT
Brlvu9/dhebQTlOQ7VapCvqtSMo6MhLC3CgbcpJShJAFb0gW7c64/Q9RDiLdwb70
Nlfpb+BzfAHFB0dd1OQ7okrKcyMqfOikVGN9u/bTm705fy99MT79x1ZPxBKGXpyQ
7l5x4tAZIAc9Vel5hOhQIwXyyGWJxUmA2uag3h602uyXokXiJrxVx4cIdh9vEZLb
L4jEZWMhgY83d8rsPjLr+haOVmeAKWtm8bXm44VrFjKo5w0pKz4twpZJ7nwBihWi
zlbtS5eQirPmwZSsQKBN7NleOY9K6qLTpaWF75AJbuEuQpgQKDZx9bk7OKR7WWfw
jlDLsPFHhdST30yObUYirXcv8LhSYIbZWAf4w4Yxnuoa7/UOh+ow8rRkfoQco/Bz
/mNoym493vbRVux9M2brE1yaoaqhWFVxKtkpa0yhCGcROCGSBEiRRZiobxHoPl9s
UDSQmTo8qprhTfeURAM8Y5laXmONu4j0ZEqkUQLFBLjenrjkZoW8JRe/xG3+aLNO
v24zv3DBlCxNYbetfSQ6xkHizGMpX+z99yhyP5BTaFjq5uWVD0Rf+y1I1eW6DVEm
G4dLJFX17/IdnCK17ZjVIo2ZRNupHS9cFg4efwlmOYSOmarsr23hr4pqlLC/5pLm
zWER5h2kf9Xzy1KhrhAvgACMcqkBPRgxhPQDOjceaNQMPiBQJN1TycrP9MtW+o+Y
GJ2wgp5NRJxuyEhE36wESlwZbGRni56GQyrbruRpt94xY9MPV8ciQdr0xxwjW2At
MKjFhFY7HcAO9X2efFEPTQZjDkj4Q1+XsKpI46+QkdbGFfz09Q3QMmkeDLCiJ9yB
GY3ez6M1qmhrbPgJEEuISjFHu6OtrqRgYyJYFD5VsX4CaSGcTH8hJurGoYpVZuIM
gIfjoNTNGkTFcIH1T+k7LX0jhwugecnVw9zMNfFcoMJ2oxfPS6PE7qhYPfNhPt35
6xiEqr+y2tiSFWj62gfXzJxOjmOrmWxORYWpewmnJbE1D4b+H38YUwI6xRRqyQqr
hpMa6RkXm50bjincaySBs7JMXL5P9bxaBylIvRmBKcA6sUsoLaLzuYh/UNBBl5nW
cSWjABlIZtH7o+n9KtRmYk21UQtykA2/uumtWyufinBoX3YOv+t24LRwh8YOoRR0
iIiT+h6Mwg1CYGZLjmcUwAvxFaQ5NlQXgeCULqIalO6rfnqDJE3WCtaoxAyxfbj3
EhvKKT+AzPLn4VobKgsuswvneUExZm7svtvUB3ICidFQqSAA/ZNnJ+Ayaf5uJ6eM
hkJ0Lb2rCojEWWFZYT9iB3y+HEukl1A1i6q26YnWfp1I4Eqgm8KM6fjqd1PMG5f7
g3y4mAENGYZMmw4K5TzAKFOiGvDbCvhVau3qENkef29bYUGkXWlUJtRG786NmGd+
BrOufcjQGa+JicXWDVc2F1aSlItNyfjKKuKhzyp1B9kk1+TLHtB3MXTzy9pmhMPO
GGWYsflAiSEIl4U7RVPzWiGPNvPp6Ly2KB76FAJtv+gTq/87I10li4Da9zcQDF8n
ufCQmkFRfk9PGAXJKaygDKPi/6yCgYFJI6tJb3huL8HxnaoMHxx36B/Gzs6NF+Ai
9K7S8N6+0I2ffQh40GV3uKHQrAr0a2jl/f3/9INum70E8PqUTwNp80xtqO0+yQT1
qOO6YnbBD073VxEEOVWiTVcFR1mXa8XM4XuQcq1yizQqCFQ0xpWTOI1HNMNelKzX
qVy7EDNBqpcJO0eYpPX/30Q2CGfQ19NjJjegQdLyULiNgPUUcJbAHaedbj3lhBtf
80xYuG8z+88xtz7AvN0yb7UrZQ92jZXUxtstt/uCAXfVFtIh1F+OroO0mqByrGyC
sKqmdZlejmoYmC1TlrzOMKaGfcVhcxkvwSzT0P9a4sPhUXIHHmGqcRsSMxqcRyfW
FnVfhjgON947KcpA5rxaE2SYh4DuyfTkzHkQRkPcxDq9kJuGkZOvrfWsC2OQnsgc
hYkC4ajT+H+L88K80RyNgxCI0vs1e6f6O55/tWqZ5hXCv3cHTJ4aDHWkuk09gfqf
Wwz7mSy3nJ75RpMdlAp1ezGWivcFkPPZS2/qa0CO45s5mp38GbeckOtoAh6Jbufv
FCzXLZKsVnQkGLJS9Z9h9HR5xA+cuzvwqsFupRxgCqGHPpQokkMLwTjU98NyxNc+
TaOL+nNpuryC4Pke8F3DlYyUhyNNEFMf7BWFK82zgm4tPOJOd/wM7Fmhar7KosM9
HeLBDmAkoNMSfk3HFlwdKV0lqzXOZ4N4JJhUZgdiMxwnBJMts1+Ytimih8rzfFpl
XZ8QMpVNlsGemYHaw8Cv6ed0l2a8yNw+9CT2+rrAYaoQc5lBXBYahuW5JveEdgAD
68idwK+GX1Y8ydnh0o9/OdSx5ZQnDLzpz6stmyPvVNMJxI//+EVd6hU0RNwebcUA
V21qAEdS2SJR5Nig932C8+dYaFi4E3deAsNmqF+gX4l4KBXb54X+u1Xl7o8j7IJd
G0OPd0OZwoiVFKTZQU+mA50oFIQufXW21cA2RcZWaQ2q/fu9u+bR87dCXIYAAqCu
Q4a2+7/Csp9+L4jSI/isvf0KgM0FQ8+QuzNyELtIa/20G6aPCByFYLm5estyp8zx
+c26VErdnmZPPpmPP9rrHOnwBvpsEMaHXJvO+AkL7MWCVtgC/gZatXJyOAYc7Kdb
3lJnNGRkln0UkGa2qE8NFYXqSTwB3jYlRApEQYyM/Lf9mejFeMW8cYFaVnJ5rxo5
t3kMbKaeKJrFkri3QWnIZZs0PvqAqpUcDjRWSnO7AQb9o99bDHl0/u1E7pBcaZCl
tgfaio7R1RlpNCGyVHfyIFVl0GvgFoG6i/Zs22xhyFyRBQ4wag1vCQyBERwekJ1m
G1/AqbSwCxHLApn7MQk0uECCf9Qy5Q/hBWPokbQNX4Z89KuTSsakAr7meI5fd3I4
SsQJgFKRi1svBS+j3rYvXMbkZPiIEBLN59HaYrhDTM0Dv1lu7+PRgdzZBi3FiJCU
hDb4oXjpIKwyDYwCa0B3gubYM7dETqgxv2en/qb28wEOCt4EPlNjCY+iTktRWiNx
9eF+JQaLXVcNbJz3+SlIPsKO/8qWnvOktSn5yO50qEmdj68cUBaAUghF2H3Z3xFS
oWXXpDbFCyJbobsrGo+zh3aMBruh3wPE7wNKjAxu2+YBDfuojWFRCYyZbh7SIcKH
i4W2HfHl3xnbIhijNO9RGR3xsAvn64T+98l9+4XtsbfpSRPNPYoq6U8+boo7q6om
+D/XBqY+Mza/wfAxRal8fxeIO9OOS3PDId75y6BlRNxHxLs6R9N0KJM5MLEBTls/
VECXEahRmmnqsgatZxfJm7GZ4cTJ/saTG+54+3Ttt5V7bGe5FbNgxD1Z4uUiNzGO
I8jvhkxlPzu4EZ9pMKE2AYh8qZZsG+7yqvwprYysuvku80awQPF6zMXvLCiUvz+e
sshr3QSwKGmzA7GHqlzlzrm33UXUi5N5ZkAE3mtGI5ZNXGrEOb5SWFstaTjxXI79
vnJ1/kwSdkg/uQjcBd/y6f/8/bZF80OP7sqwoz1kDph2jGyA5n9kEJckY0Mzs/QY
BAz+biSgUsWJ4Mdact/P6R6b55MEU1wolgs+2qgoP4W+y8BB3kEkmuFpwTbYm5ND
Bh8e6wWZmVYC7owEg2Ry0EZAO5YobMsiwUOPCWOv8WPdqi9WhEKmnunhQ7p2k8+0
WEgw6ZRAKy6vOjAodG6ou3SXRMK6LJY3U/R4aWCsOYQYS2czvlMULMucq6zWQF8P
1kc9xR1xiWGJUlvb/eReWThw6fdXrjJg0+WJCf44b7s4QvlWYo1ZGQBh+IKr90bc
B9vtWe1NRO8DnLt36I6UwN1DxiktJyuDceUMyP0p+ShwHY4Oc9zcLRv+eK8Y2No5
ke69ulqftTI3dfV9OhRW8LosIFjM1b7OOVCn4iCywzpVsAhkYDd6lMu+jkmROqen
nzVD+W/KdXzs9WaKedb5MV7RWTHU8lc6WX5q9hnWDxddsILZAElkxzZS8CZTAr7k
xD8mkzWEt8HiNLbDvLl1l4CrPwdNdO0zgo8v/wLaFGYLM64KLoj8hOJgOwMxVceh
u/fDDpveg+Wk+GrPhPngIRe4MqpqBHyMuHKzFyKm+JB0WtwpFTkff2/KOGGxfcCV
su5Db0sDR/c6xykOMfVfy1JiutsD7GXpK0R4Yyr1rVkNaaUXAiSwTo6eAPUBLemd
Lid5sKyolqLlErvbZckA/A/mxJp3tdmXu5rqNGupeyg6jzzAoSSBcZXJPnL10Mve
ToKhU9H6MnHb+KGzGQd/WVj6TYJyMPKDsjrsoMdc8rRWS33s3OYxWmCOGbYif311
nYW1OqalhP9ebEBEhzE25lcooSQ27r0J004dwyVUXiul+KpZQJuHUzt1hMOr2D/+
cpz5tGM45jclhLrymOkLnbtx3WqY/k2v7QpcdymcVw1iMz5az49LdkRXJ2Sg8Rmd
cq0lkLTIiQ9sigtClcgedtOvwEsO8tA+thU086hJqO4adxO0gr3nRk3ZJ7/pJYgP
8XU5LZ3IajOa4EMhs3cYwbDSC+p3AfVBtEXe5vsdYVMSq7N+puQEN21a1Ebwg8NI
JC4+CBJxziVhj7+KMYuArryGMiWQStlBdUGERvYdUZxzWaIsx9f/f+u0j1JiHcyV
ry9AmkuK0+FrJ2L77ELfdvNSxqnXadMqLkXE9QrFP9X7AEvEnEvSe9US8wJg1+2/
lMGlFQHLSKb57Ez+OmkfsxAKrJlBLcoiebRKq8BtdlgTjJQ/wcU3DGJNQB/MNYqs
XnhejsLoI/73gjybFTPc0iMJgxV/PqliHZuOm2NaZI3UJERBYWFw1krnyWVpgcpl
7T/saLi5p+9qmaN4VlYy8XWmpta5anB2dTM6A/SXLfC0oR0l+UB8To5SUQQ8WFBb
kplZJZLMgFB3QU7Z3gYDrIZ6t6Ak9vqT2BmSOAS+gnTy4vqgpeveN47AjE7HbViU
EJLfbxMH5CbaM+x98stKbKlfS2IeW43BqXtMc9dDWXAL2fvMHtK2CaFwLNEbyIOh
1Pisq1xRjiW6wHY007+xMneZnTN64YYRYtYuoJLr+MJuqb2xTYhyksoSJHuXq/ms
mJ3m25L+jZqDnY0CGGzADGyhV73ICWrYCKbxuYN/i8/zVy1LRPX6C6Xxs5+qLn3I
Jx175sJzGFAh2J5OmAB4KzZdskfLAiUX1eFlN8d7QCK4CYqw46Tet0p3VrQUlEYz
5y6aZ8zvx6e5CgkW/13UwfxVN6B841mBViSRxIbYG2O9PCzJGvensQ2ifQeyyLQU
o8GVuTOWPCzHG0AaZTanEMZvMVMriz4VEvWM+hHU7yr47MCOCfFysZS2IFgBBx33
Ge4uNviFznICjTBGsHllCjELyZFpZe/QvHKmPlxbiVzEP576/dR7KNZVAhyQ/Y5v
v/prsmztxsziQ9XfWuP9A7AtvNSzrfb+jBzZPN/SB0yLWpCNBt7LHrJFiO7uEyqq
13Msu8ygjuH3iytSoOFqmBAxJ+Cj9oZKepxSU5L5zlh/5TAV7JcxtHAOs0GOhGLm
o+WlsTvyB8Ap6QtY4Tgn6TpoE0XaXHfRq/us4E8w5A3nMR4e1LQ8IqGDggstM8xO
HrE0ki1Tfa2bcwe+QGxsh0MbZHPdSACHvjrPOk4gnuxJ6RLjY5QfukYvRGiwpN2M
beQcbHyWKI9csB7n2zS3kxkNQ6HHQ00dQSLsKpf8eiufhrDyT+FJuiYZJcPsHdFe
LyrarMZtqV6+ldtDsCCFxwyy4W/R80W2bindftAC2iye7mrD/ZOA1R026eBWNatU
w/iEzcQEsyV1XhUrNZD+f60vvuPX9OjDo23CAbgkwjl3k8Y37QVJqH6NdPnTBSRD
KS5Ujqu0YlnzyBvVeAZ7h4GoXcZ8pZobc0N7pceU+vWVeHjolxPWASWGt3fotWdC
0BR4EzcxSFNiVMPzQyTn2+21IFKN8p3y8koy4eiHnHxhH5dAuOVWjGa6LM8wTOg/
47koauunFYKB4I5gjtAVyKNjmSnzsmcmwy0/N7Abx08O2i/0Bue7GnCliKF/FO7p
2r78R+H/L+gvno9kPqMo+SUC2rBDvDXn6d9S/8OT245a++zFQXqtCIfEreEteV9g
2uVbOwu0gMc98oeP0ogy3ZidOYnOs5Fe6NL9a++KSpvVXT2RTL/wzW8+hMI0MxV6
yuQT8HCJq1K3IGe8T2Tk8l5yw9pSyf5DXN4ld0pFE5ZrlbvZZ9TXyz7MfC6GSNiq
Hdm0UieIe1Jy8HONhSjRve1+szx8nnWARb0QmFwhH6GgMdlZxMm+/KFBiD2ZQy8O
jU48yNhvNdwa7iM4f/SozRLMgrYenlFoNEpK6ps9QB4g9M2CGKmF4UOH6VsU3M/4
K5mS5jF6djLpESizVMQ7TY4ymWz+bcPHJiaDwuNJ73vFvc1n0hEqma7nFOGCVaJq
kzgEDdqOpiGM4tndEpCoNxyBOCUtwct2jmQZ+kEKlnMMfVvparME/02K705RGf4+
L5YqTHU73FnpAq3pcU1sV3Ox13hrKaMdwq+NBqft/cTTkt0Hg2lhSZUYwmTDAk0r
PsHPeL4qY/7GnAgP4Z8iagDLYfZKx8hvTmuI/9+vafWLzw+ljAqPxkNBFW2mexpC
yx7ZzHJhUU2Usy2/TwkpYQrYGL4by1Rsa+bnM6/FNDsu3nUOHwyDe8RHGGRFxUZd
cSGc2movERyqq2uFv1bucQNrp4W8JFS7KnKrr2Q+5eS2D60wwBIgVqutZfD1Qo2q
O/6wT66lCtAnmFW1INgiU5BXugJ+UyZFm49ZqkBsF4zK6t4EaQBMqU/dxaRBLxAf
8idoiiZHFDAShAfiOO77hmu1Ubnow+qbZVbPjI9L8CXMlf/BPJtiQDm94q55WhhT
ZsUpJK9zt2R/i432WRtPCx9OZcM1CDz2rg8IzgUR1SYV860s4UMQ993w/IbczBUP
hNfoUx9wAyq+W5ZHEFAmCmpLo4qErnoZS+JaNFZHqyLlXxz60tRKGwOjUrh6Lokx
edgqG9jZfoPtQYQ800C49LeYo2V9PxqXFD6kZHQcUVSCEs/gMR/D9MTGSjmePq/c
6BNylgkqAkeqIpiIjEccShJCEm3JHPWLJ+3UOOBTSoiVoNj/hy5Dr7ezyCubEYJV
ClCtJjA39cjTfbESYzOxGL8TDEeK5DcuiyYs01UMQsd9WoEpR+TLdqXcpczN0Ek/
ZKljiXCFzsDtSHDd/T/6zQvuRrhdHCY3G6wwQQxtF2Y7w96FW+4VLHqB/Qhpl3AU
ZgWfzJAv0IgkLFu4KPbcXAJY6XQX8+qMJbB9ad5RVNn3ZuQl6MsoYHGy4PmNOPKY
Lzjj/z4Sse+LBEHU5xA3excW5Ej4VTiyoPNE3xAwRfYHasTaaqwHahI9gYPhb/hd
Hta0CNbiVOWGc1xvbwPNl4770yiTnF3BxBhwBzLdJfE+xViFMWc1Lv77iWVU/7FX
Y8EY8cvzpqfSbYnBmu7+hM2EzdjYpVTNjr0etpCCB3T+u5grwA3lwtKPm8/2ldZQ
bpjJSsKHaRRBh3l2YDV+11FmtIHR3pgn/QtqQqEvkc30eAIuBb/0408PSFhqmafy
1IpRTrTMbqiX3QyeHrKwoh8w5e/+n2+yamRhCElrA6sGcQwd3ns+i3SgnRlERf/1
1wb//1m/lf8DNp2qSbg52EbbANlLHq+qs+NsZJ3vf71dp1Lh9JA7Ngtql8dz9rTN
BSR4BwYuNxVPXos0uJ/OngDXkkEiKCUzLt3EqSUodWWK576PYbsPKhlJjnE8M/7b
5PpMH0mnn/Unq+NX9M7XgUf1I8iRSuo+U3sTxFzlljBxv0QFm55PVodJXwDs/CyD
1OvcAR11UyBiqilM3PNFF9E5ZlKF+g0OGOo2k4RBwvUu8WKuUKfGlGe8pt+g3eGg
OAjpjG5Jw0jkusYWiXtq7YpawEGnvPha2isa56uZexAc4d55YNhXVYzGjpcOi/jk
Yw0/S70K/ZXa8XLQU5sdoNczyvJzQaKnc1rf+TPsOK5YMRczBNq93VnQjpLwDlzL
jjdZSTMrj/gAbcMY1X+6YNZvElBMrwNDaDwE7CbghL8SIwcEj3NxouZUtBw6PGfj
JmipWMruQq6UPCU4iQu1a1d0ouaTeH76ODM4I3pzpeR6ddT9yv7Licqtd79JvmaV
mh9LvumddDL405UnyInLz67nQvmy9AleEQfO+I+vzTgU2+hlABflwE0pfHuEAME2
ABds7enM3xlsTf8KjYYMud46wnd6eudz2C6NrFw/OPI3Iu1+pG4oIgU0/bXasEpj
+nmjYCgRAT5Js/YpdPlsq2xVRuOgueSdYeRGHk2C/ZdC4b7NBAelv6JDDjtdpBqR
bJqTjiXsjZSQpVJSTCxQUvdJJXSAvBkYsBZvy5f8CFV5lGcfEG9LQ/TyfCR/mPLs
nMxXTHtEmEuFR2gewiDI91Yx8sBWuZsGhG7xcEjTdVWa9hD6ZZabQ4pavIzef5Pe
vwofe4YsDN1S4vLt9JPBJorg0LXU2J0Q0dQSEZo6xVFiA93/o4x0bhVcPISM8Wqm
ei+/iNKkKmWFDLg4JfJGzPhCeqYTd7CbTplgoSjgyePIrQQE3uuAu2pHcPAR3m7K
WFx9xLx43wxw+swZOC/lZaoCTS9EYLlfUgHR4vzwEAqoHjtEl0KrR1nFgEXV5v9z
XWEVOkYcfzkRG7NVCgjgzkjAot3Z1M2DoyTnIf+6XfkBATl9THQJdDGf27tHyZ6A
rys6PC3t6pILXEBwZwhs4yeSmX7H9aFy6akjHDL8pcmXTQL2MgkPbG/slGhnfTdp
bWuLgRt1AtFTLYtRpZBXLI9u9mrZ3W3w9E9rqAMHJz57uo2VxfuRYqESJ/yKCZZj
30pLErDS75qPX8Ar/Un77eJQbLQD/guJeMMclI4xe1q0P2uUfsHXvzWmHkK7fBH0
QtIVwCvp53aJszXZWXiIBgN4gmht3VyxFoItdk12K3FnDqSj+wr3rUECECnS0UGd
0jxCoiH4ohJaMph4yllkD8SOmVF+RkfLXEATpecaYMGyTfj89aetRpSjwnwPii2G
3gzYdSLoaTwfHK+J9UD2K+mrsCjINVwfKVvImf5znsmCk4a/oIgKq6GasRBjTX14
w6x+FWDX4RZX3cs5r+RniZDZz0RwumtjaNdm2dWVH/8RgISAPVbnwq8vRZnDxOkP
OXB8HhVX5IajNq/jfUaeQUdoMVB4wL9ItHdtCvCzPjP7FAYd0vq0PGbbHiM24akK
kqJZ+gy7k7yrNkZNiFCySup4i/r9vmdr98AiTOjZDBmVAF0DVURJ8V9V4riVZPhp
WfpaH2AasPd8j06m81EuWcKzs1eEWPIDnpovAtRZL2DRhqLZdKmrphSFfCbtbMjM
GHpkZ4PEUx0grVAyZcGPbNtoBXzxoDRoftH8Lfad2rnTCju6vvhRKdfZD7VHss7y
v8knOlbjjn/adXu9Nto5b76pxzRGWZHKwoLLCsaNRs2I6eh6M/9oTohJIfd91ak0
5x6Tg2YYNK2vqC+qVrle5NaoWZxVza7vpvUpkTVx+phvNhTT+w3Lay7tw+SHPym8
ALGj36xOc9utNTjVkLMyPa2BVZ6nPLTQWKA2v+KY5HBo/g1SHBuWNI+GhNCq4Xw3
dn4OJp2Ufr9EOSCOteE0zXGf/WFB7mm41YU0MOJzZoV8MvezU9Gx7h3lF7oS+pAG
tGv0JrNbSwFsOCc1Nzs39yHaS5p4idMVRJKMeIl+wurJpyM07bJZDA7ZR9Zz+PPI
Rt4ulKJz8zmi+PIR3pcAXYlOY5R789iHGCpG/V9J5lGhrLtVwGfIojDMBdcHqZxs
2gqeMQGBzeY0ciJ7RVeq9XSM5brzjubV2COK169SYM4vEocKGyedVwBa6w2/ypkk
ztdhK8UDNeAfZr+9tSevDYWIOu35q/28EfKtDSg5D63i4nT5/lQMfRAVFfr3dsZy
RlDthF+6SmmescY9lvMPpQtsbxUx9fI8yEw3qr0Qd6hTOrwHBV5wHwFKlzldrhx2
ysTpqzNf6OJuxr2kNZqCGK3LhFj1CiMFRTu27LfVmt/04FR/kz8TohGS3Otn2rrs
0I54cL1LhaonIN5y0Of+oW75++Fy6yV5K/Z7ixEVEh9HOuTuiMN9e9EBSFTxceWC
0A7hk8AqDBCdodo6IkuPiOYvwZ2v2UuvNTYJHSRP3ddk8PTqgJBY7/iYGYmo53C4
yhxba9xc3ZeZmw5HA2Y5MlJjTjXG4Lepxsdm4HfuT/sMR2egOFVJQLGfk/yxjECO
N99tSyuJyTWShBrgJ65NJrU3zXBVAIHdIM4RTfD/oLHQgFBTqYs3atou/uGtmxjq
UmowFRR3Z7uS14FoDOrvondUIK+NMCdT9SBZzrt//T0lAS2VFaG/XtI3nvflbIFj
WHMNvKfDaNI8U3De2DXEWVMJYb4m5kaWawMuBpeulzOKdXH29ZAbpFJ5CID+25W3
KeiysvuCjVGlKZ3u5ZUEB0tahqhrpYKpLiVpHe920yEG//+O84Zr1gRpJEluqbbL
vVSgt0mK+WGi/d+OCadjSuzvlI7NVjPP8qMiSFglMimSwpCXOGUwTFczeJJ3sfES
GoLhLZerqJX1ghLfL2hE0h96ZboYndiF23A8wOe/fjTocWWZ+AUNzO0CGv3OUOAM
oz9Bi8x7gDDpPgW31Rn58uiK433h5PN8pYoKHBmkpfD/uELrGw7CWO4oWCQPRHzp
upZzwb+hUNi47R0IITjy/Ad/UGkPDL58uU4btuyDwEQnSkYKjfkMHkTQiGsXk2SW
yigdObWQB8C3uxPqmj6hIh90ZFqpxoit7jm2snA4agJu98wGkkf4AqSQTXuG1RMW
tsgKrXGdMfIsX7m527tonoQpQ3pd0nln6vww6R6I4qt1cCGKYBpXpQOj3gyXv9xD
2XtgCmPM9Uga2JA/i+YZAw4dYUaJQZRMKAxhqDhvbmUW/PjpMa/23ckYfMj/PivP
hY3daNMYS/Sil//7k9fklfskKmPiuUNpEmRhp+WyvqLAI0sYsD98kS+eZKEb2z2q
fcOD2ptM5hTyvwHPzN23uAefTC+o2zxcPeZ9YqvL6HBRGyFV8JvKeiUYEHQ5EtYW
kc0YpduDfIeXpjLoDeAyqarzRuKpJ6WzFvBxWhynG59FYt9eQLY/4Jy2wI1adRlD
YTSeGu89JohcLyVcJ0vgpFWK44PaWIwWC+E6eALYms0bS6BDCB/X5hC8fjxtRp9M
4mHOqZsDvkygSmFwGY4zW5yuEgqoDGe58F/e5fGpYzT6nXOR5XVQpNA16vPaKKWk
II4BbM1a8QVDaoC8GMla5wlJVq0/TvSF/7yImRBUu45zlEUVey5GNR2oGHwxnMxv
6IuwYnyz7WuGiVEwfpvJ3KEheS3lVj9vfGhxAS7jc1Ht2FEolTKklEk2IxjD04Iw
5XOIruGewUSoILFyUHMMTmxuoIjdVHLGRfkfm0lWrqbkM00r8r8tgOQfe4AuzbM6
dLC6XRmmAU+tDRu0zzlYH08Tm0PFvLFcjnSdGOSGQDg/9NR2Q/Cd9/4hrMl+DlW5
UWZRmqO0DVZNlW7rRktrHDi54sg+LlA5iYLSPSEYBUHKyS7SRAT2WFCKxSahW3Yt
5WgXAmCXa5uAJXjrYJu/JAtbYsIP2cRLlF5AWjaXHJXcBZUWiP7OHEZ6ciFjTEqQ
bwX5IewgL/k9BI+o4StZu5MjIjuTp4UT/YygOzhGGpMPO9NUPdsosJwKNAUAy3Di
A4zoC+e7aPHxO23O45YVOWxqcERmvPuGTatzKHJwekLl3YbAVz//t8IcW/YSEmef
cTUn6hXJJIDxOMMT8RI0zXmsUI+4XKWyuC64hzCHsJtcICm4BFZBD+sorOZqTMSD
+5saQsBi2GizMkLph39hnkgdUWkEMkTgnU9G4lSxLOvBHnTnJNkMeD+0j21deNrr
0imu3C8CBrBeKNEYcpd6MEKzqqwEdLTLvptPlDp944EIyV+/8o2zpY9apbDZubZO
LkRuRWZw9dB5rX9wTUDpjTDrSyfirTJ/wxuYNbVKqmHXZ0mwjTHifd7ISKa3Apvc
wF7/g+8bce/0pszEEhrF3q2b2yFWl0QnxBw/jmPZyUZ0flxlPgBuVYONREw5rFJp
Nc0BOxEQK+9Ds8m3ks4q1wXScjQo3CjNyOSdYerUolsd23MuWbWXRa8hYoaCEc6c
ZDVgEoAgaaZYAiMqoze+IA8Kd9DegJr+liVC1rbKSaph431zV6EPFmZTRgBctyrB
pjwb9Z8+AdOa7aFL01Dxs9vdC5i231RBUWknA3lUNE1XytKOj1mX+7zybPbFcBQB
qRbjZ6l8oJCCL/coA/YMUtGgvWB9JdfzXaj0iVOSNKkSDQNvaqJQjSvMKEH5vid7
LB+O0gMbD2lDDgcAkaOLq/steCWmmIRM9A5h+YKBnjwWRs51SvBQND24IaiO3XFv
rbWuTj+mPKeoX25LrMz69pAR+oBryFhLOZ8TlpjlJ8VIc3ocm2gT5SV2qcJaQT0h
4/cs6zA5WQ9PYwOzNkgvaT7ZvGJGdUur+VRHLcm0nclhCKl3vj51gawSt/Rq85L8
ZzIXxl4qtqp1GONJSQLXujMK9EhyzfG0ts02YaJDVea9Y1h/50QpwJALo6CUm6j6
6JICDEASxAdEDufD1fiXZyAgcHL+HM/utfGow/caj4yz6zbxBmnwZx4hhHnbDXKE
PHZTFB3MhZkH1hksNTas97rdWxgV6YHYx/3rVvVbCtC9UmDVEvHKacEcZBaWwTQh
FGbdRkHga8Y19W1dttT1O8XYMpeyCUKuvsVFOXDlG3Qt9Gn7hSomjuSsU5Jb8AR6
8TKc+6JN16GrOudD07cphcdgWZtWU7AL48WlExREJeAr8X2cDQNAwRSb5ti5ggSL
vOn96cqIFQwcVdHohxFrANUJM/KkjVws2C3MAexHnEdnK8d203PpgzjuWd4l1vxP
TOdugkIPSkO4Hi454irENKJG5poKTCgkKPvBkQhjl4RkNgBC+9uRkeB6eBAtXVdw
EYN8lVuZLZjzsXtVeq/vKH6CkofdaEECS3MncdxHlhbpEUngXH15ivUDbVYdKrdF
NdIXmKfa/ldev0FqN9BodROe7aKUiZb0p6KIQqy+NiYMxNtPXpLoRdYUUropCVfP
wmxp4WHwmB6IuDMp++i7t7YZ7kGrawzw1jWLs8sgM0gBYSo5JecENwce16mc+Fd5
cjFu3nWK+szt25vKTpE3Mf/84M/ETnUfNq+uUhbX8wAAN4DfMxbHyJyxZnWUCh36
8y+oX81OzRrFIshD5BBowv5oQrPVi1wb/m1A6unfCsv23w27c5JmPPpMjqeYQpdD
CWYbE4KZYKhu9QvTlDtx0sWezqAZthYjr7idhvlAoTQQGOwicT8FDVjOTt/Otxye
CBKYJUXobDEfdab6T+xWeRY195rcUHlTzmRHuGTKuHw853dVMaX/r/8mF+FrimZR
eaxe1bKZAxu+JqpFMLLVafnMd50TFFjQ+4gJb1C39U8/R4gp6I3aVMS3KyQ/UhU8
vTY6BCzB4ghUUU240D8trUjep0dn6cnF1yxPOFuku+XnLKgbVo+bmHxAG4Y1Blqo
TkEJ1GFqwLhY+HnUxb5Etdow+Y7iRmWQQ/BO1xqX8Tluv3lWt10lGa9dvlb0Mphd
A7WmLp1RUYgSrQ9RwfhluquTVd7QG7oRc7JI+hWJbAflHIWwZf0FusSieg1hyKS6
/ROv39NLJGfON3I1ytNjlE9UJCWXNuDacyO9fMtj/DqYDS8pUshrz7D1p+Nexf2w
MjrsvwTkPci/V78TPANgye9wFQ4ExSh/7AFBsBGm3y44QNoHix+hznCb0BS4wFUu
YGmhlSmevZf5noanV7EhaAghdEGRPfo9G37D4459wlnQ9LETjam87ajNvvl3euWW
bROK4GPRA/pMAgZ38agVAo8SUgLpensHUfZFVhx8EUr3IzjDFU/TV30QnSZEeFkB
hcSCLBPZS94juSQQfSPZ4E3uLzf+QNDVLtEu8wdB7FU587HPBjsz/ErY6j1ELbs4
OZ1OTG0x7NFf0lDnUD6m7lYyLxK5X4yh1RowsGgg+xlBZ3via1UN5BtiClALcRRp
p8ZSAxoGPHMFZUMCvbsUDB+fZpTrJXUi/S+9PtgfmdmX8qHr0JK5XJmfDEPHZVJd
v6CgEgMV+rehMIw7lhG/pQNRB5Is1FJoAJ3HJGff7370cD6RVHRfYreu1Dz5gZ/2
TeZVoPwV/JVTYzQkfqKeD5yapMCcGdffk6JCZH/nRUe5wC3GxGAaRh7ScnXdsrXA
3EQUdiPMTIpbD14sFKQ6DFrnUAjqryhHbcZu+ruYPTvtX6vxVMS3Ao1VgFVi4RgE
llCQDJ0tsm5GODvC5OWHr9wA+CX0wE8mG5VKhFWJ9e3gNpM48H7D8HpGqWkBP88W
NU1J4mH1s25+5xtSHISQfP62XTpR3FNhDZ1SSYOljj93J118gsEPjb8egd2MaATl
izmuDxUE3QkjYFIwAG6B5jqwglglUh9h32OavDNcBhzBiugBPdZVAzpB0bSgMTGM
Q4QXzfZdG6KjL1PhwJjV50nY691BAnD7pEfIMkOWegXyZahlSxijp0O7Fipmgfne
bc12un46VAeLdJeDv2SvurmC1HjKp2jczFSmFfxeMB7JWMm4D3I0R9RHUwWnKHn6
NwjRYEcgC3Sx3SNr/281HaWG1CRsI8/wqKxgUvQMVUQ14yN9wXlLD8mmcWenV3xK
3b+VIZ4IBi1PD+2XVVH35ZgXKxlfWzcZrpdIf9c2SPKDSz9U8KV1Eq476KGn/Ug4
p9uE2g1pznVZ/0R+rqX5zO+Kj9TUxTKAoTkMjsBUJGK4YopQuhFK/Reu4nZ+5WPi
UIqXqIuFoLkHgn0Ije+5kwJ7OgHkcOwt5gwcYoHj6z0uoF0TjpR2gVgQH+3+u50E
sFRPGNXbM/WlB/EyUSbDR5UHyouundhl1eA1XyKkYm7PtmOsTQpfwLBWMrnFGOnx
YxTMthzt1VzdLgFzbiuXgsdnvXO/bJrvXfiz55FOUkyvQLIDHVLnL/JPgMTjvNQE
HXPOLh5sZTBOvE8FgIBw2SzyRnjyo+Anf2UwT9B6Jt0bStXvSVcFByYFlX2kSK14
Y3KGwBy2GXBPUkRr5qrs2MQBbYkpYM7admmWb3txFe+Qu/qzR7Xa0zDNoPeLKU1r
3kiXjFS7rUv4Tq+3g5E2Xb8/V5vx6dA3x71Dkcb9+Ze1bF0kXF9pf4+yIOBa4ECl
Up9uWZahE+nWkMz7KS8y0pJ38kKz2fMk370GaIJNs7D5VobCgLKJf73iL4Zgk3/k
6SDde7zoHlIu9JqlWFZZXUEx1U4OHKe/zwRqgcgg6MrK64o6b8esecNHUs0H3+/M
utvkJLJvX+p2OHM0vTKlQ14XRcLPbZ0CHQvt10DMMB17Ehh3YEWnANl/V8jivEls
VUGZq4iTCcGe4Q5qybNXFijjrnnrMvZmtu0ZYkn8ch7ijKtKTzRlAiV3+1eOLkM2
sKSn2qDgRxZVHVEz1cjGy4g6A1ig7Qsa7KY1Va+FFJRBBZ0p6Qe0VS6E3d63slQG
M59DvFAvZbYcYojveFeO8P8Y9U5nfkjH4JJlny032gMR3DtHwdKLfela7Nw22jFy
w+X9VBZhwMbw3fDHYkbnQkyWZ9dg5VlqUEJZjGBChDTHVKh0AGF/+MKVD3GsEKY2
YTJh1wE/bx3di5YCq7LCFH4qmQN2wwKZQAY22ERyTqlPOx/3km8GzYPxcb5vXsgt
cfACMmbwoFsTgdpnqwXBy1dlZ0Zwsv0ByTI6FdiIE9m93TSod7m8Hrlo/wVIPmM7
7aUNgeJVnu70pj+SUysyJTzxsCr9u6ogx7MWXY6Vy2kqFHgsWBrIKHBDBN6j4Taj
ueDgovpwckKFrpOTZD2tiVZsM/4ysiPtWa77mrGtpWC/qDpMJU5/cshhujMzA7o/
yrCF97U+dmOlcjerqEUivAP5XG3F86+WYlMUKg5I3B5LD94FkWIGUpN1H9V+jOvp
tuGsBKCcXmPHGq4Xe0pCCEbHlFXlqoKQd724PIdpt8hJztG+e+2oz7vraDN/RMvq
4tNowcplockxJFiOkXC6PkWaUjxQLK9/z1dRrjdeu3jxdSHecwiHM1QappycfRCE
6XEmJ0TmyvyCT8c/kwcduemO0JlH4FFxmN1EKnu8sLWSySIahRFEiXvi3JW4ci3x
kBlhcULB9R9yMBQHJAxTZCDMwSs4YyFeQoCcFpoTnlU9K0t0vRV+VLkGxIQHU8zW
ewYNsBMYG/Og5L8LNwuwwq6MguDCGPh98XUpJf2xtrtLqmxCbTYlhv9Jmj3oSlNi
NaNe0G8YhJZEr2eXZn2Tz9bFLW4JTw1+44Rg8BB+H34tNytx/mPJ3tCrS+DYBqPy
tItRETgvfq50zFpKgpxmCP0JPPw5v4ZPwTPelnu6IUf54Lfhn8Z9rE6JujiabxRV
Vsu/kG4JTYv9XueKRrU1IS+W56cz1NmovnOlxnCdpUGpfn24+bOMmu4Fwe8iAkQp
R0rSfBOKJCxsUNpAaLpibEBgfqkS7awlj//k3tJ1c0ng3fNMzdEDAY3EsWWEv2TO
U5gW+OhhEGrE7qJ1ShbfbdMn3+gGrDsvCYmr4QimRwyZdECvBVe4zbOsfcbGpFNP
erdLTvPchrjgLT7auUvwdI2SgMjzHBuy/QrHIlBdOTfKrw7oN29jxs0gAt1FL+mS
in6oHy4C0xnR/sAfmTxJx/vxZceLObOQkePVNqq7pgx8n0cEzKIt0qA5EeH76adF
EebjmCyCZT58huwI31naZmQwDJ3/NDEUUQfLyvkESL4lT7wg20jdck7zWdFQriMt
aX5xO9d4aIqU/X8uUInPQDSSkI81BBhcHVVs79WtNX25rnqZQaXxyghuRGtlyM3O
bESmc6sI0MGGkaJQoQkt/3Yj35hA0KDtUHRMMpXIJ5VQMxnCC0eBi50MJkfjLb/o
dHRRpI7zfzPlUd/x/ers+gw3V77MSk+khU5ruH89XbONtQvog5jakG90+pKrsU4s
O4tEiAhuv87Gyti8dlNgBKJjUyQJU6MZNiBkhssYY9s4fjnJBjBa6punCVVwXDVS
EYD9Xuxaiw2zazKHJlkTby1pnzy2yOQ/6Vm13/dvQh10AO5qAUEvttixIYTbG8c0
Ye9TEEFkkYkrPgQCOv89o9mYlQG2UvcjW4ObKt9wGcxyGEFY8oewIxRnz2rZk8ty
gyuEUzlEEDOmORZ3awAaYOE9UaW3MPRWyVLUlSx/O+ZD4M7gkGz4vCggC+FgoNJl
ZfHpGke6uSQpvII34Be+fUNXd8ojX6EyzDcT/uPZ1DXNnxChk2Jv2ZjJaZw+7Xmr
mZLFN7odI2zNQXDbG4W9teudEPiwbFvZG1H6o45MwKwosElene3NkHEVA21QrCNh
bBznMK8YVFoD7tL4Vl6SdQsqOrqHgz2/yDmWiCeHIBtc/6dxZgXrBRqAd5Ko7eD0
ohDicyiFc8d1NW6LmrieH3w7tguKi3lDVwYDCvzhU3HK6G8znr9riqrFtEp1agyq
r2yNPrqblVLxDnM8qEQZT6h359cAj3O3T8swZvK1lq6W/8mjf0BqBIBmhoVM2m0D
rhphZQ5mChzIcp6QuahGfky7frOfiST1RsHm8S9Sy/yLqHt3ijmRBNG/zGdokjhY
cwcqNS9pJyD+f0PhQE5KH8DiXDh9cWGuhIsjodvgnKryDnJSYBPRa7LMR8O47IBl
ZxzLr+sdeTD4jRX3bxCnzX/NKvun7cqle1XlMSwH3RYPtaYwBgJtHkxb8WlC9yQx
QNUj4Bb+PKW9ENPE+lhv3lIFaS6i6J97A/wWa1xNjbGhUZZlwLt3w40IyojYPNAs
5gySBULjbmmU56RasY9988f8oOHDrr9Q7soejC++JakfF/CVoKsulmGhHGD/I9Jb
JS3CDf6jS8HJNsUerCy8il8vx/+JuZJBMoHIsVlW4KPLhVTD8xRmDFh+4xtpDOF8
7iLCS4PhEjkSxR7sDipEZkyG2c1n5wuRRXm4RXpo+eHNVMwxVCGKZE0Eo00hzUvi
sgKF3srxyIYovx8g7QtKwaU7N41/8cVKC8U/UHFWC63r3e5cCcJgRltEgUXY4RXz
L5JDQTIASHovd971ZFuuwJ4MumcIlkEnaUS2QkHBzFnuHagzV+ZXUaqle8z3MsX9
ANcdxTGZ/jwPGWDsofPaMkXogQSWf/e+f8esuJr6R+txChFCu4PNGd/im/PctBxb
6hKpadE06a8MKZ9RSqcMcseYML+1N3bW7TY1rNnYQsNmKldqr0VRAMpnvIMmpCqh
j7JxJAoUMkYJVOkEemOybGLE7sgryM1ByQ+6OozozNHUscsCMdc/Ky1xL1o1OHOB
u/NoTOwIzPD5XbF1+9sD58mwCvXHX/HuCvRb7bN2heH/lZxvS0B01nXW2e4BqNRA
vnqvPOzDHRyjUuhYEhNw0lYISyKLRbjOr11fCytKDEilfHjlHD0ztbYxVNZ7RjmK
nLnHYdGhzVGqbvkQkmwwNIKbXaMhLGcFhHlgasklsIZc4zm/G4weVQ4MwDY/q9UU
QVAbsRgeD0ZBMTKBgFCdvrUwDI+RFxyPHkY67HdM40V5qdVBmluWwzZH0PdlnUib
Hhe09keFqYBeA9F34XpyMwWE+XXadxyBfUx3p1AMNNK6KJl4r8/WACGlNgLBr0/S
3V09Vta7ydqXscNVKbW87UC42g3IpXvIH0owz8n+D5UFVgTRkNVOYIuDpAhefD4J
yImBn6ero/9xB5V4s0/F803wUayFZ3GhnPRZSidgMhWD1BEmbeAAg2pmBw367h4d
or43L7w+Ja2AAtnwlv+ISbcGFHk9VJIdEqlvSy5IuiYM0xLt00o7x1CcH1A3X006
zszRbmL2yxehawI7OgMkeIzDKbouf0Hk0DR/dQizQyITXXa15H7CN6ML/jzxlwTW
RAPhF2LqhdapJBLTbhuuGzcrxWO/Uy7J1CTOr+WXqQMSvgnapwMLqb2o2NNct9qG
Vm1NWDzScInOSRiHCFyevn0rqTFVFJk/vXkv2ICH0PRQyyhBOcSC5DpGHfuG3m0a
Clrky2YnUFokD3wZBFYrTMEoOJuD7uVJI7IVnEfna/HjQLEr7r+LBYIW+0xCLGgb
+aNFYp0YEcsASGe9KHIy1Kn//uGjWMqHHYoNCeZhZjeybLqJObVi08wkY5xXE1cc
U0TFaaZ2rgk07wUtLcpY7RdteFl7y+1IWHL9MvriV3VoHJnG82wAL63MX652FXRs
bImJZU3SIznXB4tdEGNUXXoSOQEyZ/0m6/EXEsqcL7C11Tx3VYkm/7x1W7iCDcLM
L7QYYqNMQOUe+NyuVNs4Zcs+DxqRsCB3A3eW90bXVgo6h2xBZ20I6Xn987klwqz1
vt/de1PIq26iF6xtSmSEzr+WtGYgHIZhkWf1Lz3HJw9gnnQQin8utIpWjXS9n5+K
3lcAhpzQUcKJwWII19oQ/IqQnr/KL7N2CPCo6ktIwQjvsmMys5SN3IgEqiac401H
m0pIJZxxsN/gwiLI43nFPUWYeeN1p3Bxz/+xyxzauMrYCEl09T2cdiP7rSJdfirt
3FzRoSagzhRHH/pPIj2m+DDFvWlsjZCnCjtBcXmxlaILPg7NPHWjBQ8Rg6Q3CQnx
Tu4S4LGBn/yQofqMRYEgupNud/wSh5t4fnx8isGGJANRCof2itxDnjOZ7Ei6Vrse
9YVP95z5QQ9BAQwRGhOySwHsSobTdILq3snKL16+GpmmJdqLv5umK4b1tExrgcCk
+GEg5zJE3Iv8/039F9OkW/ExH0BCixB5sS0hvHRnGkkNHIYp1mIJBiqzjNWe8Z3h
IMTo0a1rwgto+IlZayki1uSOCoyiJzC62y2cmF9uIDj/gQo7JoYmm6zTGBMGGJF7
i2AzyJeSaFUmWLorAebL3NBNZt+gj/tjJ0BS5neClN7SjqUV6917hPma1TF84O6M
rbpuaP2xL2t3yh9Z2VQ5hKZSJo1AzRbedE7Q6lX5TMu8FT5/qY+Cn7zVApak3AnU
6JhSkV79xAew8oxDoBq6k4B4CnegeYkxEpErwuKN0S0B5o9bhnzXQrKIji9cRJrP
iEg/paP4NevG+XxEys48SHOVQCG0zOYXe7MJJ/ttgDB+cfHA0PWQEv+FpYWk4O9Z
X6Cb8TDFNs42fJo8YOSup/FtY6b3ws3qD1mPu2YCvb56SI8LsP+1SpBBU1iMoc+T
xro1x9mggIzFC2U+9b6tlxg3BzzBn48ZsmzGIJgk+Nih9rnKdGBHvKlaqpIQOxUW
4D3NRQ+tmvO5/U6scM7QKd8xB9ZzM84qz8O0NFIcP1QMHl1lNuhU7N3PuSQXIQBo
hckIfbxuuv/NLnCJsmIdXBGLL7T9pExoHEfA5DRjfx3ZUvOml6hlXKZALS8YBkbA
VqHCR+fjKmx24mk8Cz6SEw418DBjZxuiPsKJ8Bho/yF0GlPJmA5W4zx+TiLN3Jlk
vG0QbdBmjbM1FLEvlmrv0WZUXNxvvFnKe6gLL9wj2ekFOCm4PT0BSZ9oAxBweNQn
LrHIZeY1WF+BZORmndfKu7OaiaV8DjJ13vG4xvUh4HmFPv5/xrUCnplXlYvKRAbA
DVWSvA9wTW0+1Qm7HJjmMSO6NsFy6fRdYDWmUEsoYd2GPH1RqpwZZnYlptrPXTp7
eoqUB3bp4LT9B3Fc206u2GT2L0vjf5bEIqif0FbCudPftX2cCXMy/YuaNxLj7w30
FLXxS+i4GsfU9b8pnuFZku+4EMssVjEQQXa/C/J5e8t9ThNx9VJ4lOHM2nXLrwyw
Fq4PYiF5jgg7LPfLL5Fmr08GBTvZ6yotGktpM0nrPg81uX8vF4iEF9IoubW9L+9/
oY1YrIAJPQucQv0ibgxZ02l+feYYWCLyhgtu0mP1E2tVU90ykI7mJQ3IVABnIaXY
wJhHPcMTJ2xfY5an+tKgwRLVL5+EABsYdLDIavQmRbbKLcsd/iLps2E19MzR00gY
dnTUdhGGXYU0mwny4sHgwLyQMjBQuiCxQc6S89+IcP+lDll7rrnRenX5d01B+Sup
4zjc3EYfQ22+B3sUDcwPnSrLUoey+12WH/Nc/MPlc/Ekj1YT8qyjd78EejvpNBn2
1KBPkRTNojH0IgSjInYYN/ONZ/THvNe5SQe0HUda7oPMxXwyCmL/g8H8WH01/R/0
aMdBm3bMADZUCBEsK7IKoXTASxH+T0wZxcbKMJsXMQzv+a8TPP2uxkVETnFwhFsm
4TRVMN3oTG0VD26tfxzbowOK3PH/xPNzYeuuBkJeKGdeGtLydLYNbJ1+ikidVlvb
uqkst1PMjMddxa7l/vb15Xfsn5Rv/TKzPODZl2RjE2SrjbM8Y76ttK9pScZY4XiM
a4sOscqVIv6mKauH/29Bt+4fraVVhKVCRBcvIxhfAcShPBQjsDByT20gjeD5HcB1
Y+FDLmWHo5xPKpk7sCyEuQKV3wFW0AQT/B6hnBvLWk2xSlT/nXp1ts6j+8hqLL4v
UcGz5Uuq4RqVzbPu+R5qUGNAGud/pkimA5qS84DyEGYPzoZ4+Ni90Ce7HxbXwmHg
w+iEdNTRrd+75/n5FyGpsHh/ibbVgKHQJ+Go7hLMrceyjSzToL0DmQbKGoY5GHth
Z275DiKs6U3ZT3Ioiwz+OypCMIPnzB+6t9ArxabM4WMr/8DtYW7D7NmQ400gvz70
2m+drs5JwNtJQwt8jeYh4JEQ1xFWZ8WtAflwg0yaQgwdLXnOcQkutXZ2gzSNGHuB
Jx8AdgTpNekrhighmmB8YHUZnYjAVuMKImmrsUlteCfA1Ix8Or0onp8AZpxTyF+K
kUpRYDlJ3JWhhEsk5NVfw1nzIrt9Eku5Sj/aFJnE7Crix4I9TEhyUbr3zTlPJyCE
U4BotgLPUYnOnWJ7i+2grQqyYDiCpICsw7zr+jQpB4p8d4lSuB1hJB95zbv//pp7
wrKyeMkjEmU5HfMcNmg/JleNhYhPJaIgE1UJHcCqp/LlhBHvSJ/BDTLv23K0UmEw
alDs0PsaQaBdgtMtZPWjl1Wki1ZlS0M5uKOXeD+8eivC2FfKDVqDnRnvxdtYa2gF
exIBiXz3IwBh9FsQ5BbLbVE5gd9dXM1UaEDWDOqf7TW1jDyc0f+oIJp4eGRxkljZ
aB5+Z/XI3umuo0VZZYCxaXRoYjAR7nK8XQWeohyhinZzRy8A59nqf+e7wJXZOHL8
tymEmUWRwqmbrjZ7NIGR2ad9LAepHwUjFCvcZjxRCzsBD/GzGDBTp5+Lh9thE8Ci
48nVEeSXQxpuePS/KidUpKqwsPSVq2Nj1YDNndlD+54JBCFmE4dVG2f7kf6qxyIL
kFCCF9FhsRFNiSGDrdspjZ59s59bbNOZDypkvpIDRRRkIZLGpf06KvN3UXgMa0UO
GklXYoI+CqzGrjccfnS7ndzdLHvowLX2b5JlnfYzGvVl/6MSZLrSDZPG+gHLjLOC
IFM+IjnOUlXV9MiJtNEteaRJjZHbtBZsvCcpr57S9CafdVoRUo3lPi1nvY/uJIx9
UzuBi5vyakZyoVDNHDdKhP7Wl/eXPDmE4Mj0exu6y/ms3aUKYSoo25Dc5R/AXniU
BF4Qt9A3UYQhwmDfz5f728rU0RWuqavORARNZi4X/b5mUcW1pO/KNbfVbDkvai9I
jZznXT54cv/a7NFEXXWzmRtF3pyGeZ42Z7/2JdoekpnJJY89yHoA8/qJOKylasQB
Gz3GEK2IIUCc0D+L99HdnJAOVNVue3I9nSiggtRv9FqBMeY3jhP+kaX6ofCYaR3T
Ehh10vymAXFs9j8xPRUlrlJlacPeGLZ1Dv6QNX9w0SYK0RxQ31QdiFLwtKzUPef9
fMh2hPjf94Vl4oRQZG3K282TAwik2SJo8b82WR3/QpJeBSxuVeTI3dq3m0UQMamQ
7fMzEMCAySF443XI0HUgX3S3/4Wkq9hdJVwdjslUan0d82furQMy+6mBXODbAvgt
brsO/Xcz7UDhW5GXQDAIoWAzLOO6ZOSNPDoxw6U9o2/JeOUf+PXz0iLimosuS/Q0
2adH3QLXJHa1v3eyhQkeGYJJstf4h9EXUHDoZ45xDgqgZO8aYZLEbi+xM4xaFjgt
U/YYAw208M//oqfFeF0oPfLQ3K+eDxARm4bxqZjVWMRcvdtMH/UAVAg1vK6zHhWL
sQZN94PQZmfGrdJBfVAynTps43VzJU/5rpkk7uFI0Kn92uhbDpStYYLQ/kB5HoJ0
FXE3tsvhjUp6kFPZgVPUwj918ADDqX/eJ3Wn/xeknP89ygDLOMYx4b6HyfYhqsUF
AUO+J+eLs0AHinOkIwp/1UtocScTJ/2RUXmFXTkIBJ1q5pgyCqKgA3lT3ak0qYRt
F/5+hmu9vKr+EtznIzRxf6NRLrGoks2e1M9oGuGwr1aaDlhxNAx0cCTGJxnxvt4R
4hbgyX0NoasPkHW4BXY6+1BfCVWuC4fe18l+skiXqDPMC9bldYGRB97jNf5N84w7
0jiaM5uzj1R9U+e/YoxlplKhz9IwqHyOJLjyIGiYoNUCsepMF9+TJD6zsH2SuKZm
fI85OQ0zIVZviu9Ga2bjyX7Z/IWMBo7XUwCCs7xpocdbkrlEn8CnGLIZpd0Z41Vw
0xJ0EjdOh3Lj8jRtV3pOteZ/dQC3uCxgSifIL92t1AHurNPHu10q/zan+gnb6jkC
GVtNH4H42U3qNbjqSLaaeCGUr/qpCBFZus52/IrqtvTPqsHx+fsMo1IY610eELjS
7fweY5hIDoRhrjhgnFdCBFaLKU4s5wGLWJ8fcTu7KwofkYHYGCH5AvOs7s0ZWSeQ
AWVxZu4SCUv5xG7yr8tcevcXDbeWvs6RlbOLhVkdGSFeRUpW4HgbllK9evYRzn4p
TS62phhcqPD8lJRBrmPvZpaIQInYhxe2oqD+K/Q7WZ2ibjSjry2GFPOHoJnr9ByN
C7omvWUQDSqYJEb0OgOkJ8xx9VJf+PQG05OVlF8NtQATSCBeKdVZZZ7TSp4ig/b9
0RhHC+y2xmhzTjWLYlALGtf4TIMu91+rhcR0hOTznSRJQpoz4iWaGdCPPR9n9OYB
M6i+O6Cf/diagZhQ0rwKBNJkMKaBcGnqbCnSa9X7cuLRQZHynaOCMaMFy8WWD5Xf
2EulFbaNh4X+ORQJtOvIi842IRJW1QsSmHVzhMtYODSP7ieWU1uGFPg5bP6c78jl
CXodLV8MZZosTd/wL1fDTVZsxHZr+hXaMGbiKt7uycyX6ATH/AYPaQTnAgwbgyeU
Ki7QBJonEU1NDZayOAE+aqYn0FJ/6EY7zhMDpWw94ukG+eiJuNdwvEQE5SVFZLrp
tqJGWCq0fD2Dv44q+w1yF3X1Pwu3FNg9h56lulWlAKwXMqZGWkAYn5INE9mhXgJu
1xOw0zlxMle3irix2BxpXbrDSrp0AEFJKfXdDjcd1hGB8EhryOKY+lBBUWtdF64Q
Zo87k4WWEV3vwSMJ0O+kk0vbI1sXZ41Kx5thXX53pnRkagHXXB+Os+mGZgamMVhs
YnryplHRXGB46iCeN3liDSRHI3x6nYxfLXlY6YGcQhvZyDdNtyAq7lpoQkYqRCvg
myCHAfyHU+8hXmhgLfwRN47hApdQyhbq3JfIy2bF9O7MxfKFbvIIz9uWuVgK6cx5
FHz7q5vvC20mvckdnsIP4Y7RIJ0qrdqnHQmJBrhvPeFS5hMlp7Y003vw/q43gYUZ
1kQf0NK2iznZcrxyym3TyBIwzY+zxBqd9mWXvRnLcRIMoXqjtj+koHFCSAkf6aLD
/2FvvAqFDSOJtnL/Bsdo6zpfMb8N383NqzC2eyqQOx/lbFmQLCemnVh5OJIf8wXo
xtYLaBUmOvcfDsCD3uNVLfmduYF5uNTrKMR0YfxqUtSFlacmwDFDUO7/Xpjaa5Xi
TFBeoWUnf7y7w6uA3Ni7fje16f+/DFKpMc3W09+T155pSP7cUrpGGRs1R2oUsLHD
C1tqpWZznstnUH+v49i3lgx+Bi3i3yIQLOLT0O5CODytt7+4uxQCIfc/JtSvJXEI
KMhuxFKottLANUQiyAfy4JdCLvKXJMSVAQyfGytzTmKzD9AOkHwhQUx/QQNIayOi
SIzLUqnuC4XV4aqGMBD3g2K82mxw5gyR8vHNzL4lzKIeeuyfBFb06AFUe0SBSgld
bxQ9I2TYXtUueL1ldRqvSnqkA7WHpwkNhb0TDiWnkoiu3Y6do4StajJ2X258xdmv
QHMPz+fxtF4MDIRf2dNQjhVM8q5Q/ePkWddTtp2QQHuxV2zYpxgl5M1qN2sE9NYt
Zh73ED19eFcQsWkSH/nP3BkyI3Tot1ebRk3kwbLsiMaP2o4M4isHWUWyd4AHzy2n
wFwy0kVMppPJDhNtf4b0nZIn7eYnRyAJOr7vgCqUhzBR6Mpa1b0Q3CKZ3ElNlITe
sqigLt9H7BGFlcDuRq1uGPHzobPzsJUCMGXXn53qk4hJPMb4wsqImtU6QI1lu59q
yh0JeWd2yhubSuS/IJXZSme2NvvtYO2N8ajVRvc6/UYGnrPD1xcV8H9GaBItEvva
Ab8CnnLJeDk66F9njvwVO6lAcyuxTcQWpmxbBZ4JsVmoPCRDiK2KA6kLwIhhY1ia
HlJxLhJcTxvOF3ewZWkStQCjnpKq3mi8SJcsNYNVffCC0KxULJfZx+qUpK+oEEPi
IwvDCxh4FQHTpNkjQ2tdJe0hGSGzi1BzSD+Hc7X3M64Xnr+mkZtC0CS8koSliIcH
w+yc0di820ouGwVeEGUkd6hXsfgV8B62h8T+4LKUYprfldMBx8ombfcqq4i/V0tm
JSs9nyQUihDUQcXin5uStC3pTf5wsnFhk+weE+qBs/8pawrgX1OMe/h5kEALtSuh
lKgXeG5S3TP1LyD4CHJcjzxGYUGFm2Pydrqpa8myTrvDjHCZ2rXA0UucfxjMgS1I
I19ziY5lYz2IGgpZUlhwUqjTMKsjj+wNnqfH6STTTdRLW+R20ZIrAvUuNqxvZ6ca
x7UU9sK6/GZ4gU2ol4mXTlOh4xon7KnlsKzj1VjutMktP7BVLlHNgM4yyqohYvvm
GWOXMK3YT0+hv9jEiJcwGHatN9hb/rFLN4lSN3IHZOQzF6MshfBnl+3XWk0pVZu+
bl084TXmQVT9b9k1xgCSxlq8R2TChw3vhp2M6HNPKtXByjf34ickv9U8PbonCwo1
yEnDAXvf+q4R6s/3dlcV/2KhkchWrK6WL7GC/tVAD3GqeIbneEqC8Kg7ZVh73r7a
YU2fZNLBpteJ0mLHrVU/URMxGD/oj0xH9Jo1IgQoQhTCYAtsJcUhD7YfSlOFKhX1
4w82ETmcQyMAEdjUM3XytPGbxi/NPEOOA+cH9GE1U3ro/OTeMwUd/Tx3qoYjdr91
AZ2dFIYDQq8mImLXpY/uMJD8vIVo7ebc7I+U9GdX6RfNdaAEScWnA2v6H6XZTo+z
BS9G1OUc4C25DKP3/duzbphu72WpKOCxRYCw2mrq0o7asf58emgiMfP7mwx6O7ya
7qbZPdcZT+uwRphLSYX7phYD0YrUTqaDgDmP0n8yn8OIDwmBmWyytuswpwW8NqI5
ch4bcJapTN2kP1H7JLBVgDYPc4JN0F3QY5Nth7X+05HY4hNXiptTTKjXegI6PEuW
UfRQpi4neLmvDOWdMcWdGk70PVmvpGbk3hZqBvZvrMxG2ceakYxhiZ5Wvxztc9lz
jKQZfN7CdBd5cF/kLjbjw6bzMTc2wiiaVA59Zsve0wV0SbYRW+i0byuVKnTR+syl
dtQCp2GHNvt4V8i/m/UV0NZqw8kY55qZtKwKzZ5oPk1ooCjvlAlKv2c6FSf8JT/6
1Y3rHR0+HTOnYUDL9k+TWV9QbZhmxwAIOC6o+mv5l2L1xXXsw7bB9TKPuTH9L4T5
QW0CCR2/xouIaed7hklq7iikYI1/xeCTvhWZVWK1NUSLVKWs5DdoOBql9/RwGtTF
n9fXxQTaeD/lXuwh3AVBKiDvFf+ScU6LitxgMfXQBCfBw0Hy2cMwQTS+9QSKj/Cv
m7FlZ+tMTw21iao+nfS8i+kfSTxEnpfhwZhSCSXYt26YJcd5l02WhqjaygSYW9mV
YTrAWGdFnLEO109HY+QFW+18UH/mXHVdzud1f47AMT/bHGAXS5VjMDvfDszb3sH0
1zYDMBp1haCgzAS1lY8VfV5edkvaR31oVWAYEqHB7MMePkCyFmZn9PPWUVtA3ZYS
5g8umFQK/OKCoTz9a6WIjqJM5CnWpbYrQrWxVNcp9xTpjZdtJcxvLbHm2un/V2DD
sLAbUuHiig8Ofzr0Mm2Mt6cPoBUxmvkku7dBH9aep8uSft2AbJey8orJbTAYUVFc
vTU2FfE1b3ufq4FrfSOnw8UsXY+77TdgKQKrnucTORLq2wNSS3SXyk2Dajk4vPNd
9DUDNTYR5rIH3IAEVJbtz4yZcbVN2Bly4eKRgovILN1ONKCP6AxKer/FOG2bkS2G
T7LxBNTC/m1Nx7La9+NK54Td089Ir3DuC53YBTbr2DIYlkU7vnp0PTgWiuYbjRzy
RK3w5UoedD5+67OEe1JGAjzTQU012Cffo4EetMnh9IwtoL9HYAgKmEVUEhSJrlBD
Jj0bPzQSoz3PtavPWVPrdljHRCOAHB1Jd5PqgyPHQc1hNGK9D9KOOllI22//nwGG
7ZfoLLm+/Vk2YduMjjk/HW53N9Bjyu+fcK1o2RpRxcsbyUNp+TmJg+RyunN6OoIo
x0X91locBhkxOTLEO5M0SWyR9S9sR/TxGtzehQLBhvcQJUqPpAmwm/eNWk3y10n8
qbXnM2B8/Rb2kTOZl8wkvi0pxq1ZaBjLZX1QWP0NNa0zZaj+hqptfgIUfBAT9XV5
gNWuS8CWx35Lqc7e9BPxUJL0+UkS/IEGqIWGH+ifgxv6+5ZruMNo5ll+xC0G9YPb
8KrpMZmdFnlOKG7HY8b5FPAC5KkvfC1O+Gf96+nTjWxalvg4RnBtbDfI+HEfvDe+
Izfx4ka2U8HeBveL93TURvGhp9ZdtSfAiye7NN2obE3RkDDZ9tT22fVAbL8DOH6o
tfRN6c4Ej/MT4WSeg2smKTT7kADKRw/nWamFkMRttgTI+caKnB/chBrkpG/VhmIr
jAjxAKMzQ26ohjsXf+plvLlaip2bMqpuDFdqbBCj4iTneIX9sTdjlNMWz3x93tAm
D+P+YBTaBABdukcOlbp1IPebjaQqYP6Q5t0t+1YwrGh7mZZ7HoFVbVoZ2C2z7qLW
JhSwbZ9BKKQ44lQ6nz0l2rRE4uxq0w20pUipUAAl8G3i4sFbHk7PB0r5dGyaRTdC
BS1SWoHDKU+73R/LmjiN0VytL1tikwpGN/Ll4GAJnUJtNZ6RppRVHWqMEZr4RmG/
j1ZgeIY/2z9PvVr+qJqJF8UE8u/QaFiEjM8qB+QxhxKiY1yXDRyhAErTi9rIh0Z/
O/GpElc6OVeEnczMV8mdWWfDKS2Zga5Gnovxr8pKdzoJ9zmSaxiadzugXBFqGctU
2O5/yRPRoGW6WKsyXR+PVwKGcIL7ZfI39GSLw5cUMmVXOwKZyCTFpeeeoCAKg9vx
t9nNm8ZK4L+VOqILnrwggZbJoueSEIgnDDohTcilO/ZCoDvG4jrjhBL+k+OgsATT
lUZh+7tXAsASAHXeH7ryoI7dm7EqUXTLw2TR9nPiL/VC1ayPmdqazHfPEuXjnNz/
WJ+fCPTD+OGZ56a4o1LNn70ByJ5nrL9mXzjk7xDKf1Ln+xdD9eDiWfkO1/Y7EMXW
YT3xZ3fFD8k37/GV/R0z9B7diWSCDE3H60s0QEe9JAqUC8bCW6RKzLfeX0wJR9Ah
0lzbVJAe0p0xJM7zq2tmKh++Zde6o8GiA4QtVf8aeL5docNa252+Ylj46vx8gw5E
zomVw3zbf8L6ulM9APiFxpLmLo+cu9YIoMYJOeAWnsONdCGvgEWwY9jdwTS7okSw
qHelvVMvuMZHRUlpoCSqReAac+ZkyVGvycg6wJwftUIkx8wg/GrXXmE/7E4lnU9l
MrmgPpL1IJeGH5JjSRNd/fPYSlNpoweR7xfk79bD4WMdFIG3AQFegiZ93TzZKLfT
AZ0lxYuSEzAMCFqqa/aLyR0J0eL1OIlXO95+fTMcGckUkLmSXmFeumg3g5GlQFQg
WfWNLP0uCSQ4XM8ah9Wfrrf8lzjd8YaGHjwh7HmkFv+Zd7LboX9YioAzmPGfe+T9
0mW1IEeUamnOLgAfzv7KeRs6kEXNBveHgVeYP3VtdX6dWs4dgk0qY7C3vCHoN+mf
hF47r8WJeGGDxJZ4vSj2A7AlfVxT9F4g1VyUDc1iHjG/Uudl0VojzFtia8NGo9u1
5tY1PY5lZIuM4bbqX8A6K85aUP5/sWw1tEkiS6zE+tUAMMXvbiq7oegKIhtrYm7h
vAIGHF+qIKGa2pVNvTgaKXetRZ3n8lzIb/fYl7ghEOk9KfN/lP2UDYj1V/SX0IGx
3q92+6bbJVjsOkoMdX2Yo+Av/1cy+AdpHqyOQzh2fC9keFV11WBplsf67JluABEb
vILGfQWcxNl1+cRGyDE+q7h94aAjHu2V1JAkka+tSpAlO3Xcz60IzJ8hJNr3lqnk
+jBtLQKVldLhrCtVVDRxacVcGbwbV3DFwkYua4uAahZ1+2ZZBYaHj9Kyf8VKPngd
+RoAXJwcl6bUMIho7mvYOhjkh8TqkQP1lqK84lPc13tWeQVI4wEGn4cJ45kdvJAP
8HYhM+4dl3TwFDCUvbWtOSeJ7UxQxBD2KiW6/u91sbw7xmIdDFEJTF4x/k7Tf2FN
70jKCqAL+PaIC2RKbVSfcPF+oBJ0donW0RmazpDKNjCbHUie4VFGxlaFL9WIHGKW
LD6yO91oNphC50rSnIMNOfp+fk4J4Vmzvnzx+VbeRs3QTpvn1Xd8HP/ycW1W6oBe
2c5R5gdobNppBA6sWkm58Fm2I6dh4CFjgBneRi+HC8kFNhgAPotxKJdKC0z/IyWe
tH8oYcncGx2WO2EraIH8eQMtWT2sFbW52+nu3T903s/KUFZypgvP6g20RnzqzmBm
cjnHEHGpoVokoRhCec0YMQlLrbwlaRenEa6dKL2OahBAMHFjmtgHLU7zPrbK34g5
E+sK/XEBL2kUjf2G+n7AYvFzauFoKcVu+dkxLzM+jee+71A3p/tHLmbqBxBYix6C
xyiEPz7oKQq1YzphgtqQOBIgSzPU1EvvFJYG8dBeoMfkLa7bV9kIKb+0CHiGIG/9
`protect end_protected