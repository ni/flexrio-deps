`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 17440 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpB/YeH6Nb8mC/T0P7RFHOeGxk9fePrEw22QOUhOTObw+
wNOmCgbYXHkq4AOEDAGRuWmNpZSZ6NDNWeF+9uQGiRoroDX4qe3LNa+wzcddVt/Y
V/H0Wg5ldvaNOrIF+lAOYF6BOwguTNssh8ZCtuxdYGuYuJeMeX49c0u1dA7Ze60d
O2qxvWASzNSD4uZqzvHcQMfgpqgbxcig9E5skDqv7vzsP+U1L/5ZYDF6jNwaf79e
HfLLCDY6enHchrCBNCjwk3k8ke71WgR4I2ncR2E5g51BKD9SrImob7kwKxEpxgKw
0uPPoj7ZFldu1BkusE43pb6Vm4nTj14oqXmy2dbM3YX5KpC0VIHjXX8T94WeITyO
w7F5Cu7rHq4jSidhDZJLTW/7SxJFvs7JFmiV71r/u3AtVQWVQWPzj1qMNU6xQJS7
9k/cGJZHbxWO5Vw8wm3LBoh1T9YzgfAK471RWQOgO9npjchRh0vaNb8rmBHW0JNm
N/c82DMgfJ/+e0n0a5KT3Y37Ihjw+RyxALBI2WVqxbB98D7DVrYyEhgXRtpz9aTR
Wd2qbY0U8F+GkLcRR25CUx9XZGvpBWjviEvYMhkam6UR/ACADvuP9pH8Us/Ys74H
ag6FEPvBnIL3X873fW+uZDUYfUu8XCc8Qf+fCHWY7WmZFdASCRuClGmvBtDndACW
thTHkbYgmCGVB7WNbjikca/Yv/LqpJX+QvBN6w9yF5e7nO+/Sb8FT+OaTkGfx9zR
hETsPp/L+0jQKgVIcFiNdBCF2ONgDV0nCZTRiNlKc1iQnibsyOgplWrzOwW8Ok4o
vUWiprFpdRQuW3ekwvybxo/v/rlM/zzydjhy7rRQu6j3IULlCc7IWljUt2+/xcTj
eVfotBX0WKBCDyBlyPLAhbXLeMb4dKDxfalFIiZzEEjRGmDqU4G0qzUur+W8zUuw
9Tth3/mpxhXs4FgKU6888uHDTiptkvGqodtBx/nPFcpnUoliTUhDu079E2rfj2qL
aN/KuAV8QuKsyG+WSu5tpqry0CE5ZFkepvuj6yeW0aMvdZdAwkUtZSetPr7LurEr
tSXCf79xATdLzV7FmkfJYISYDR5WuC7ppnCXTryKt710f1kE1hb5jJ8177Tvbcqs
XteTpL5c4PmsjPeEVw7HXrbzY3gZGOFfFoyqkO43rfsIhfTGpcV/Il0us9Tw6p7V
P4RihAuDLqPvq9fjsLK7C1LzUGY+fGgJLlx2oA7sZVXXfo4fJ7VScdQtQJpNznAM
Gan1ztkYJG9Vvi9qQ0kx0Y4zXJzryhgvGQhljD7xfM82mLiJTxV/iU9lBs5eISYk
29KY9YVAJGiNoIToNz+cZwdX1gUCW7IqwH5kF57Si2GDS1XGB4F8NcMg+oBpVQi5
YFqa33PgCsMQTEBf5LZkEm8zBwnQ4ZaSYEq6FdN1Vit+Jo8HDUxvBaDTYsxV9aLr
tIB6DOTEtQ0Te6sNrgzGrpDs1Ho95l4Mfe2yfigk1+mpbT5i+uwwi6r1YoZ04fuF
WsHbGVUwLsdQic/q2kuLSqcKvirmvxEXNvYLHSfqiODT22+6phCID1U6SXw0SF8+
ROkcQIgyE2i2WSMTCuRHzsYN9byh6XMjl9HXOMjp+F8Ce3QejtlAnR2zX1WF8aFW
u2ZeVjo/FQSd+2qcnNN1CTPDWEx9jzECH49Opvgb97L3BJYhKXPBhLezrWvjncQf
v9o2yoeAJMSCpTbzBhiH1uaEH+rVy1hMuKq09lHBXI623X4vGTrolgQq/DISGWzQ
btWx+b7R1M/6jy8Yav5N84kuTKEKpum5wYIgUKHJt8HpPtxeotlynBxQqXu4SZXK
44l0f4E038nBpUpUQdoT+dwSne+iaQxNq6xiftvNxVCb0YF/g9rLtZ3/0qNZ6lKU
Bf8Hrfus+Vlm8tlJdHpBHTU4L070mKzdjOFBXvabw7hLE0MJu5FbdEcxxMyjjPb/
/ajQ6dA3awpGLlKJQ0kEkIgrrWqJ6LMdq30vDxxwv1HDCaJ6TaeX2Rvx1rAE5A+b
+WYQ4IglT6G3JPuUJ3uVLaTVkyOovMlzGS74VeeOXnaQ4hhfxLTurcVFAK+lfM75
BPI01o7a4B3kZNHwSKx2aXU6IKs+zhsh7/SQs50sLAQGOel/gXc7mydGQN4uPKBn
xj4ZtiBf7/F1cn8Q+sZ4AfS5kZF+rNCp4cPzvVAgCjb3wMcGi1pcWqrSshUjQNR7
kUWlgv49mIWC4rvG5DbrO+5UBHSPoogrdai4zs+ppSbzsKe8OF5q+1+OGqn5sUH1
MY4EOtikFXvWGObCoBioyodH0tY1/pbySYgUMSGogvldd7Bs1s9jxqfKTHyUoPHr
5THahGiwbRoBAFdkdCp6mmt/VgWq3+UMo8i0HPIn8NiDRrxCw4s1SWbY9d1OtkdP
jaLGNQYoLiLdPCYenEvksRzSGUwDnFLhxPvtQHGyPcKCAQmrUEeTDaTHtBZXf4Zh
gZGja57J6rr5miwa9YZztFnoa3vKtfbdn4XhIJbXl6Ej2Upf+NtHod3nVs/0Y6LM
Chj237UnhwzAr8EhNS3WW3lTtHhV7LGJ4e3nH62gGCc9SYKthXQHudJuuL6AjxQe
BNXW9I0pdVDKHHUykUEnRKGNxVXGe8SaSh3b7HdTNYALX4/JOY14kyh92FSPngVN
eSLVCkdw5XLH35OVGMGs+DNT5Jj9NbZy5d+1Rhdoin+nsfOtlZ1T5PLUK9Jfsh01
usELAHXJnpBhcbP495+cMMirxBZq0ZmCHP5j77j2bqHQZi1Pyz357rNvzATHb0up
l41suv+Vw358tfrtKcpADNUKF9PAYqA97zEwvnHEIKyfTkL20oNjO2kfesD+CS4N
DxQaOhPXj2OpCbr2qxbbEku3R1fJ8WmV6bxP/SVJZjFES+3/Xf8Y9regX6ZQesKr
WZyJ4XinwK4CEEDt9E/OcNGTd5mXnucVgW61k3LXE+00HIxISF39fW49akVkmmX4
TpYxeZ4ZzDYtcauOKhXFhLdGLx0Y9kVPJvo4TuXDriH9X7kZcfOTbDIkLvIaKKbY
p0QET0xSr009L0HwDffStB5nILJoDtz8DM9oln8/R21o07OJtPsHmX8f1D/FpiKb
ZXSpCHTeN2OX8n+w9xj+eKx5FCK7FVMhXfB3EhJ+fylVTqdBc+r1NlUljvCdYoda
vxYvqxdLEQLdjjW8lklAt34ezGeb1IN4zMYIzl4O3npYTkVqWmgwStjsJQjhaWUv
dnFhdQuthD3ZdRTDVmhI3yIMtLKkDtIVNKkos6DIliNtFB/wxb6XhL232NN0+5Lg
8vJkPFb2fhd0IjXJpyFkvBCV2fYPvjSeAxNgWNs5vY4SWV6cXCrhMwJQY5FdCbIO
DuOI2CF/TmzGSYrFQLwQlN5yt8Th5xcHrCaIAKAWK7NAhC71M4Jg/G2gtPxDsH8d
NZ2BXLGyuoj59fY5G1Tfk64p28SY79PiyTqRV8Bj87i6L2Y98B8T+hIlG0UJslYZ
vEy/tCoqsZMaMTTHhUjqMecb/yWOgJ3hSv+cKXmMmBE4yC4wrxawJeVJ95EAUkZB
vjj0HAJkh2QMN5L8LyrHoKvA4VAuaumLPfvPvoiUHcL0XCvUeGkOzQRbg6J7TkLg
i0xoZSkWxmDTAjj8w7U3JrZDc0GnquEcNOHPQii+qD8mEnnSn89Nts56OtBlhN0T
8eWM6+dP2cK4sjv1IWdm8hOuwBlfSK8x+vHSTyZFvv4rtw/HcLroBFPGOZxUxdKH
XBV9uoV2rMGlgGy0NlZOvnlELson0OtVHKEZmpWuIBSSnEBt74l72y6W1It8ifqx
PsoK+9Hr30HqMDi7adk2CSpb//Hj7e3XgxYWjyPtSyECz7LUYX3OHja3TsegfGNT
h6fiHJkKDIwK6BsB65PZKddWD3YhoeQTQbz276MgnrYJJNvM0UVleYXZCDVe+AhU
Q2aEAENJsTqv3UDcdYzbekzvWZeUvVNgfNPc2lqJvGPDj6vXLqNLk2jVGG8MAXGq
s2okzob3kvB3O+XDOdRksHp7v1Eu7bzVp/4vUTP/UrySasfNiPef0FPB85c/lrWs
bMIP5n3v5PRXbZ3sD4UXZIBIcvOacGfGpmK7hJJcvsAPPcCBhlrXZld8ZKgVyny/
62x0QoPB4G02CCf/rguKAi4P9QGeCmcMT5UAdcY7VRlgGS82hbKku4uXmShkfQ0U
eYB+tI93HBD/p1/pXYjsT5nYtnslGRhKmTaVO/CU2cnPjxgx8/MYRbyDUsuOG6hj
aWWz+JHYA8ihhBzJpuiu27qH/bmiwc+uQWov9TnmVKgTMTRYi6adg0OGquXWE7O0
omXJQBmk1odQgOdmhPoTxdhcm1i8DkGncCikGQc3BTRK05yCPc53N4S5o+XP3uRC
6wMbdYWfdybKOR3lAhphVD23kB8Tn3yiAPqL2ZH7F/+zurC0ZyXuV/qMPRYPaOCf
gsKJCFFcXv167203DaABV+6ymADpDpoWDqnMSLy5ooPHcIbb29JmGnFkCE7HGb/B
WXBMXK999pJZ6iZTqBAHxx2dzjKWd6RKRpUUK6zky4ryZ4KIHotZBFJMMKjxgP33
XC6CuCi/K5dye0BdDeYPygfMUlv/bRmTVkNrkpGUHBBeKWEfKrJH0fl2bFQtM85h
3LNk3VTXQOF+Gtl34wo2usk0Tqtt92Hbuo23R55HVdlK0jAnNAfvGmKcNDJ/csrX
tWHZQx+3Qe5Kw2HFTzoXPLvKzSCjiBQFdXKINdQvPB9uh4OGL/hHLtSMfDc7sORk
GzVpDAuGrdHIygcAhZwNlrwT9Q+Kz7+DiiD84LLYiPEE6Br8YBnx9pGX4fRIXowb
D5+/I8225NDVcMh8AlDeTBEmA1G78hok6qWq97sHxfyQfUfR7I0P1V/nWpkXVNtq
Ufa2HBN6CgkDXJSybmHsLQyaH5fRdpe31exLgV4lQEb0KpFeJY0qgSu8jeBhNs+A
PzxNz2pSYNUTDKROAmH4/cHXTJa+IxRLUNYRGNKSkX7zsFKOHW28xz0M8Hm5O9lV
MuOPZxosD6Co2SgcRXbF+wH7hb9YEaP2SJC0Zg1A2SrIj3eFZh0BF9Xl9H9hZdVF
2ERK1fJQkjxpXtBaplFeZM6D7sqXme6FaUiB/BQGCRC83Wr1mOBHfV61cb3HYfQn
xdvKv5m2qnWNje/jcaE+cVLEt9ZOqTox+j8DzfrZIo+l0MIS+9UxNPjPe0KysUGa
fZXSZ1qq6TKCFALl1/2RcP4n5+F5z5CJ1F5VxaEbpg6kg+jPhVzW67lBOO0CPF6k
qnaBlbUBq4o4CDoYCOvDwLh+zsMSU14FgJ394EIuAQKAeUkaeC7Tx3PrEHi+oN8e
9bSssXz9O3FVf/2jtmMM2EKaoIptRZ8pt2YAtPeRsrN/PfV3IlgOlE6VsAWgbbPF
5357j18DHg/Ke4dsC13BiwYLYiMqGbr3myEwcqD8Ddhtq/IA5v0yPWF3U0lc9hOL
tYDmcxzjf2yvu9F1cnX42tT5fzMANfHFwZEPxJxIoNEhkzqFG9xWxZAV4qhy1PVs
182yaoVmkhG+56SXrYDIz98EuxnScrKTT6sOaQyrwLOinexewGmXX8L4fymq3B3w
qdk6Vw8l31S5doxFXt/Xoh1MFeILdfa60wFC1nRwP0Q3owWp8CjJjVaBqVKAvBuc
pR4WhWHLO1t0PoAdOmEY3dfq2lVgPMaucklqqe86StTYeYiSfyKYAC0C/w6tgtFy
+8UjI5ZK+Rz10Bitv0hJDQtRXyewtsb28x89D9PEyTGnBSBPfhua9Ou4fm6zzxPY
yuGh2GQFsH/irM4tBGXGSdIB0HEklA+smvzzeyxKOy3npxMIAFBrQEOU8KEZXltN
kc6+WETBdApz4LWfY1biVjKQz8rOCZbA58RnnE0lcMhunz650aurSQ111GKRROAc
9DkeFn6DSVX6jFcMAKMN0shoXVgeNM36u9amnT+ZoZxt1ko7Mo1CjGZfHkx2GfPJ
+zQWd0hdP50d3d1nfOHpG8QkjpDGVgtHnKzl1YIiPgpO46OTgt0RzIyBGR+gWLKv
90fHeVflI57snJHggMP25PJd1uxJo2MTM8MghbjoK3CIZg72vHN5dthKzfwpgBXU
TuoBszCvywE76HYCm7Dd2Kf1GU/a+RSufKokRWkL93MUOzSL7e3shaImyBc9JywE
kgURk6U2DL2UNkTsg8rj5r3p8t4JwCO7Tq9HkCxWqs9N2Ro//SkmITenBWHJAupY
1rK1oJhl7VgafJ9hHN0MehtNtC1E21pK5U/Kgwqksj26kuNBfuINjYQ0Uzms4Kmr
D+IufnS/JP0E93kdmAU8X9fEd3dk850DqqyhFWg356RJhXLKo87/HISy5k5PxbvU
RSZES+bcXp1P5uTidHeJjunNHqrEmJeXg+CP0adT+L0LGXGRkw9dNIA3b7Hjkmgh
yxJDZYPyD4CS6Kn63p06bFY0FmQNm0NLaluIsfqQetiuqSe4RKshzzw+S8+XuBAb
rUFgfv0O0x22IfMP1Yv7da9DBN93487hm0eNMsjh3Q3VEuBpa1WnrY1+xvEzDGM9
6iZi5iM75XqnVESmBp2mp32grLrXS3AjZ7ApO7InwIpXruQKxIhdHEEZ4A2Hocco
9F0y3oTyOjTLzPTPxBPMJus8SHx8v+8p+8UCTC7aQkhGmTOzWOxtjeAwMKPkEL9N
2eeMPoN57Aid4KuJ0JbGqvevyx/K5PiU+NmPO4wRd5OYu6ItqXAV7jrr92i8Rp6D
4t8ub4coUhdofeSL3NOHAp2VCVde1DqZY2lPYN1Usj4VfdIMvVxcxKqX9JZh6lC9
TC1E05OFsQs4UczvjLHfxrXz1mUD3Q4VB+oENgH7AVKao5lPYbxqdpyqZAvy4kja
c0q2sDByu+4ht4N8GLV29FDrlq++G1c1hZbJo+ZhFOfj2agt9cV5jieSq8r1k91Q
rWwslrJqOUmLCQppa3+VYAGpCqAMFfINURIx5ub4ydR6uCbkwOJu/7vWoEEy4W9h
pCxzlc2xfJKq1gFkMkrCnkUqbdrRj1urITMW/k6gD09tJByBLQBkt3W8l7OjDrnt
mj5WIfieSwcPO6BmBK7hHWA/2x/ez3oz4TEEdtksop7b9edoh6YUa30asba9nESB
TWEIDiaYHc75wiVR2jH2cR4xyWeNH5PT2xOVM67S+Xphn34Q5dTwBLpxpbf7378o
PeGomQ3SB6gtjxTaYaEQbZcdJMzsbtWSDnwLxRXFDtMGtbN7gB0GDqa9U95+051U
2HCnEZGB5gRmulEHjU7fleoA2wpIgk1mQ1kVVFz9iecxwGA1v4L/CsTkwuzhCMDw
aK7xURNKL7bHPsNykXRGiUxJ7UPtwdLxoftHMcJIV7N0rDaXd+pcmCgETMlH0ZEq
GCvlEi2+EHuGjB3DHzEPhr9nS8re28PCnarbo4rcH1jPm6DZziSZxAHaVpZFu78L
5ANvrojl3izD3UPfH38VwBAJUETp50aY4S0B31iyO4AmwvYCOFhX5NDtt4IQarnA
+T5iEg23MlKyXIu1oyhmYCL6/IyH4xpIAbk/pBkwQ3hhy5QMkURCF3869BPIZmfR
9aoqCwabGoXAGCt4ZbwlF8wsLO1Fwm14ke7Khjd12DedVIFF7De0n5goun3//g8a
088ixFftOngjBtD4xUu3TYAoD8kAKzcavqTnot9zqqC8+ElJHAHxlfZFiabZacLc
vifXOx9LH3gOP3YgCMG49C8zcbDKTg+LywH0ch8zcXk+OSTITgRgVCh9//gRgdwH
f7mqOwyD9IcujDHCnu5uqK/IyJL+vA24NVucT3AOic3+XZwRnBDpZiyrEP9zFXGH
Qb6EGJm1IgpamsZxGe64N63I3QB+5r0hm3PZ5mr7MNE3YbS1nUNaRYvl2aa2uKGq
AYGSOF4AgYQ7wvAHmeXYMnUFkYV+6+qkfjtoNsyd2plE+6b5TW9vq8kw4Q6wUHWw
4HUDexDFSvvYBHE03K2QP1ELbWJfsBhZpM9WuyKYgG8IG7MJ8fnP5N6wTaoSYUtF
nEQJzxYJTsMKn7x9bIKkBPvTdz0/Pg3al6TEwli7TmQ7NjecPaBqjn52aOrh+AEB
18MJkBxFtMPbFQfpPeZae+i22pVjf4iI2+ceiIdJGypC33fXrmeNzPhW4Tn5FLzR
mS571fLuz/ZZV52A8+zetMwKs35yRms4l212CvVRpVTDv8OWv+8o1QtPN24+b3tP
ZYLpjxFY7m1/0gtDfo0xGS2qm+fnpdKAGs5KbyrsBsOlUG0UHEBnK30tNFCqdW4u
GQ4Xxwa7SVNa6GpmvJBzNnfGm/AFl3djQ5gYKvXIy/wCHqpwskKq4cvKa+N0Ypay
N/ZHEGDoJ0tq3bMe+gg0pWvycBBVknlHywqWXOO5jnna1hiexcFc4Ry1wl4JK40z
SZzAzSMzGo1ErB+pC6OMmJ8ucKfp4yUEMAjjflsgjNbHU0aDU3+0zdrjhz/Vmb2e
Rs+8ri18qSGh+pRqIHoYXVU/m4BADMIjy6flIyw/Iqyf5ZqISzoImIygy5VUtP8k
R7k/ojOCKbtJeEbOIC+LuV+/FFxGCOCqTyqG1r+4oLPbC5D5iOhPQGsszsBnVhd6
vTigVboT5AoFpHPM4xs2WQWiamPS3RvglRa2G2mv2l1qFkDvynYstKp1eHtxi33f
XJryQjj69w3lpYkwdxK2WpGdqD/a6ShYzDpvbnvyUdwJGZcxtwe2ZyHJ9QOltBnD
tY23ZGZsmB2SaaE4ig/904nPATHkuki3vDzenmm1F9UXKMjFJx3sn/oLgELGbGbE
cKVOtbvhMTUkpgAT4xSJK50yr/vswxouKXUrvfZwFVE+VHbIT6sWwpIJ+XtnRMAV
kKh087otg60ihCnhwWBLu2AO0QqP0PlGheyWRqcsrXklvsW2wNYl73Vyje/hE8S9
pRkTOrRdl7wR7iv71vNHltvi6mCcrPW2STxp1kGiWABQqMbHgerPYAIsqAMLQyu7
NgTp4dxe6EVTBH1qsBQf2wNGNoD/oydMUQQNlGGZx3WVmMJT/+87TsqJ8GXGY6na
MO0VVG/LteFjUsOEaSYF7X8T2KM/mgWr+A9fnK+D6uE77duyYHw1D4tzuFfmdDTg
mUHN0HJxs+X+BpOsLS7tM8XsW5Ueb7TvbZlYYpSq2ylMsMCB7v6zSjE4D+og65xF
7YlN9Br1lnBFb5Z4Q/dadw6NaMb56keCmFedXuQZTWOdH9AOlKmKck1egJvI3jYQ
vBGfwWlSoYQMAR3jtDe5idzxVRCEPKmGRUafAN4tvHpeqXx2QNUPaaGbAC2MNrX6
DR6ikvXXLW8Wm81niIuS4gVBL6mSzCbAOS/Jgix+uB5oA7Mglc34Y0RJaC7TIvOe
mMaPwONpKqvPK3P8mYfpkb5LskRw6EbPpZuWadYLmCIXoSjT4BHAkOi0lOjKUW30
0QJkEeTH24tAH4uvHXsde61lP7WwF/wpV4zprh6o9nd8ng7aj2FLp8tIboVryanx
XCc1jHQa296/pVt8BwUBUY4wpNv+w/GjN1yN3mEBE48wF2aCAbm+b+ZdvVtLhp52
b3R48Sx+xSkG7ixj4uOG2MUXFNnGyF27HS5Q78I/6NNcrGXWg8jN6N6V8JzE0QGq
jupHJLSY0hTwDTxFGQr2Bu1nueBP7RmSCwy+0Buiy8Sz1ruB1+Y+973gjY923I+z
dbPRvAD/xiD9xJupImvVEbO48XrSnk3NQmGdgULp/Qqn7PcNNyWh5im8YQO/7pN/
W8dYpHDoMWM42oNNWH4I7yV2yCbjFX/+f40LWXJsntoY7JBgHae7/6lyqKm9mQza
cy4Sx4rcpgGJW/Ys+PmtixiSwOY3fHWdevw7MayFFYxiZw80IYoEfwWlvu2LFhi7
UWVBx5Lr0Rz6XnryUZ2r2pw51R2CReDXiZfFz8qceqYxpOKhdnYOaeX/47dz6VOC
6W73FTYXvAS9oXbYCskhNFq0QstENMEt7UQqNGvRjIuw38TJManH5/+Wa2l88NkO
SxfRB2zKXk3zQhQWrDKdGjHURcL/Sx0+tKuHTbGAV3p7DXkhwNZRKNfHHe2RG3BW
pOE4UpMnxj6t/neR3xGX2nAWxS7fYPnXWs2pOxMdupheqj7VitkrJEYH4FGCCpd6
fsEMQzThf9S3Vf7RGeIKA+gMl0WQNeFNY8xbvcjsNf3PfgkVuLUSV6YJ8LgOeMny
A/zMR81HRzp3zZFCWhjjdc40PsCcvpHCLWj9Rew+wRYS/yLoj1UAbtjSe1iSqCYq
IDqF1WtIJJ3PPgRDWWJIA54ZNkLJyf8EtPj77XaniXkTXYsGyHGjUD4fWRzarcf5
i0WYr9zwxjhNOW7Mfi0gVyvGsxBP15IKpTxaXqBGsmVndrrJ3MGNKuyixUqacNc2
oqq8vFkXXWboZiMo9F/lQcNKYDlmrw0a0z0I+PBkLjQ2ztqNXnDR7e6LSbe1pq3k
5adTOreTw6gBq/vZIE2Vrw8zVLzLU1AfIAXkcjTUVjEI7AIux6OlSUpY+vZeV6Vr
Ej/p0D5ijpc1Cwhhz0bRfz6F3rv/9Bz9o4eHRW6x3wERQgMMuJnpPaZ0pvLhWUX1
BkMjCHjjff9iynP7mVwW9dKAOhuKxGig0eS5OjTqA9aWw8V7ETC5K8ytHs9nvBeb
8boWFgOSrXp75Pq4wi4p2iJs/GRKB+SEpnhqxQp0anBU+nTNugQs1rejJeVHAsuJ
LbrFKQD2fLdKo4AcJtae4RxysCYhomLt3D8VZx6olmNg+fWsaElqqO5rNe0uMLo2
vXSCWtLxka3UuZa3ZM6jDDmqDHnT3WbYE8FgxTO+x6cLVqBcO2EUrOx85f8MGcVy
7nyFpIH8u+q1I9nOG2/ljhtmBctZU96oUi+DAyl9xMCyJrLcGtwKAhsxy0lBOFbR
gXLJvly1blkLL4FhelfKHs9UG42W3Ay8N4b9eTl8ZNBRVX6W9eOPAlgr4ltz7bpU
Yrkn6N8Wj3WtajWdlCtwdJaVxdluRkKQMgE/aNUlcwwfGS6SNPjgaIk/Nuz7rIlj
+pWqrO2laQpSeyaBCRhtRfSxHmcyvgJdk+69UIuFy/HCxiM598aOAljnMORaF8R1
3NOuTMTfc6MfCpz53eL06Tq8WjTFjtiQGPyHWZo1tGZm6iWRzoQ3yx0wW8xDbR4I
UZK7stDFgvOwSc8Wv7QWpVc9ETt+fyucQkSRw2/VTIVpBMolKKcXPrt0VPQnL/v+
Bi9DONL4o8vHzxmUmnsJVMnXDCPaItXoJs5IM1MIsKU9CfDzjuntsPrnl2xjqk0G
3K3IJjsm/MWKKeeDHuKsCdNKPxuTYsWPMvAU+ueel+oyIXkgU+JzW2T0w7eFZm/h
qdQNGBbLWt2PqJCpt4A2VlVGBfvaVLEqNBvokPvhWEON6Yi4OlNnZKwtpRut3KiC
iEVOXACobpK/QHqAVrJlOHAOlbzMIGHPYCEckxheTbxgOP4uByVGlM0poSD0HUDr
WVdx7A8VSwD+VlayVzFHyAfxt+QvccQYJodMiD6xtklQoexVDMCIbpft8G40BjHY
4V+mVqRrDRR0eK06bmOxGBc4PnWcankMbc7nhh61dsvFRt1bC6ngjyQSWyZaxn2T
enQyOkMPDRVxC7KtJi3y0dCL4EaTFyCGCKm0JYM3s5lHiMilycU+LpbFLgo6N1vb
hLNGVBxvsVNmpGdc0O0XJ6kcjxdkRAG0uxBwqSanYHL6Wbm5hjYrxeqIh0Rmstt4
goirvVrL4/D8IZUckuiQJc8hC3e7s3E9A2p6mOimfjI30LBJZlHYZOuxE9/3masa
Kuk1NM1QAx8pp/cFBpENYc2KiX28s8Hghh/2f2SBUWvj0vYq2Ds90yDP7wzF3BmE
OgbSwSX20prJWu8vXy1wb30kX9mR28fUJTFGPMCzx/RAj/hb+yeKiKi3ah+ScMD9
ocKk9x29n/M2r5LbMINX1P1ZGjE+8m802L36xV2EU7wgLy6uQtxhjESspZl3Qu6I
A+uyjcO/I3CtVGNM8gEwy6gIhq+S5RZbrU7n9VQim85WYIqsi4lLc554y8CCyMz4
k1TNhYAwNJSBxtWBP5vE0Maban2NE6uA6oUPrrZ3ty/LJF7ilGWREdISXHNH3A98
bO3JFqbdmB+0HEKuAxVzOm5SLMxaJTGHJ6yUvbaHPprZ7vYGzexRAScLBFUhmT0J
jD3aE6gFiY7/mkOksl9b4WoRlHoZIViAZncoBo4QQ2gctl3HGgt9AyCOR79Ahtfe
QPnDO0zBHW7/d+LwLMMnjR1j/id6aaOa+PIz4AYoOWDeXs/XTmhpku+SrWoPxNaI
itmdlhyYhk8lHNJYjNJpAIrqKyfripCf8xhNTOXa8+7MqnBOjJj7ZEYGb2OjVvQ0
krHO9ZtUquoSZEtrJ3qm8/bQJw+bvjOFPyPR7AY/eJM9CCBjvYV4HrIBba8vBBu/
3l+pYxPUby+iF/Yhcl+2iEqzdhr6zEofuACb1gHxoLg6pUMJXJYf9uhwkx+Tj4cx
4by9+weBngiaSd/Irp2SLS9XVQJ61DMjlHMVxqOgTnRjDdiDTmrFeIb3BCk/1iXz
rYJ2Lhjzw5XweiTFo8hWXJLiP2RgtDzMFzE1UKbT1RjVbFNaNbTkWYC0ygNV93Mh
cZNPxJz+W36R4COd5vBHll8hfQ8/LF7VHJQXMs0lWxBUpZl4yqFEchAMIqf/XcJu
RX9eap6biJBl1+D4RoWE8sXbvXqtdlLC7YNzU5AG+edvYqkaSceKBr8243J0oW1i
6O7EvuV0F+Zgkox0TafCzYQumhvZg31Zz4y9KlR+6PqWfEoiwYPTFqDs4r8zcofu
3b+AgXbM7+OMDmFlsX2o+RLibOOEvmntLBMMzh906YWEKr+fmBNaklvmOkv9xTw6
NcgWkqWZ5931LimdEBIufRBgbTzDECQb1fsCO9xgXbiMJGY3p3alTOB8GhQbtBfN
a2eJjONIZbgQzN/N3Td1oROSgsozmWX0DXS4nw50hJcqrd2+U1wBDmgdzj1GujuC
VQMOXSS4lbwiFN7T9NmBo+qNcEjh/MY3y5Gi7XUdeL9c6eOc8VSL/WYIGtCVqqT5
wx5xAa6gnVX3Qp2jXPc7wm2anC9hkrQ26Z15XuGTrtZPfy0NkQ8qbFn6K9D4qBnG
ItYOs4y68a5s4otV4Viz71T1HRJdsojXzLn9n6OKhJKjczJrLUeA/pYfKsJdLya0
iTHNXD43lEzg+kb6mAoIF7OkT8vWELWB28LhCiw4AhwouwaDZPEIikKTTcfbNm+L
8ESKRLMnjrf6i3m0DEBEiNnH2w58J4ZG9tYMB/94xEB5SSnjs7tZb9H/rtShtLzW
nPsNEWakOfsMSvLON2o0oE922kw7pQkeIlm0501X4OF7W6IGRH/XFMiLIRf2SOWK
4qTVXERi56jiqepaBg9LlQ62wxe8FZ+B6fnWk59GbQQwSnCVCKjP2pws/+0o47oq
iDBOW9DfqWLyCxF4nV08iU9oDvldAW4+qYLFh9K2dc2QmzWzv2RCijf6wr+CM93T
eN4HVcPkBaIJJv+PlLehUgu0czQCRzhGWd7w9DG+NXj0Jeg/1FywIHYjaloLSw98
Ql48jkiQKizNpZcTkZIHxGuqtoNWnx0YgzY0tVNkNIQxa646LbxfVr8UCDmSw3Rw
4HgozYdYssgBr72ycU6ly7MZyHTN0QkwAPBOwt9CF7d3Ht8xtbKehssGFilNTBBP
1s+BGihOHvbDOs+nOAlY1+mq59GKzMNiTfLcxVnRIhb0A7sV/W0pJSusJTMX68Za
CHedlxZ0B/UqsuavQWcFRFoGzH07lkOoaib1BqTqlz5MvmKRS3uqiWwRRgM7LpWu
uvTXd6e4mF9IO5Dynf8lXHsHBUdT9jpul569YUxYj5UoUfeC46O0+PWFV9LfA78s
RcxGkSc6dM/2OVt2DbJVgA4KS95Zy623Dkvn8T0/+z+rUk2Ax9cgfJGWZfFETP+D
+RQ4tyvhPfSooTycKWamfcpBTFJ598aDkubQ57TWcasS6YRvfq1Ga+GkZjMQaH0h
jlMzx64xLGDy8mu2zIRHpC/K5zDZ8qbCIodc/IrOYVK+89eUGpfn7SJcXM3CPNQL
Zpej5FUwb6eyjO7HJO7E2SGzKgIFV/vdbadhZRQYExl8kHFj6HAjy6fMUGqoUFhC
Bl4PmUFGNEhvPpHM8WGnXjbIUW8AV/kO2wwGiNkuZoVGokpg9tR0kCVs2Ux+t9Ew
F61dVmfctbPqTLwmtjwawxFpPZIaVw+pcg3y9ruW5Ck6SpFtTuTDwsODObsU3tV6
nrBcPxOVTRvupFZ+SADEJqamAVYoiz4B+IvpWihQQpmSyPLUyM19G2KQEvSXhAVX
kqCIgMga3S3F9oXB3loEwBhPE99G27MAYdRS8Ia8XvdqStbDt3H2bb+j0M385CAN
jms05maTxgtc5DpS1duPkCIqeogEfAWpw6Db1w9iwSIxhyYuNezMaVw8db+V7W2Q
G2yiYLmwK0N69EQfUZN/3wEvhYAR8CAtX3X09rRszJWEWwz7S+rYC5pampE2zgiS
zkUoyyY+mcHeju5TViz7IbCVZJN/H2UlVRc9jspyrLx6fWO/n5ZODwj3j60yQ+ZV
ge2s9wTauPJ6b4PeqNU3HdoKcIeTHlK3pQwYMLl1Wbq1hX64vJtowkotrP1vY8A6
C+JvWKXe+/m/H23/Xg2HujoFx6Vh1C2qGXmjbvVToyLFkaWN2goXeuIVrr+QOlKI
aD98XpoNhFa+xDth6jJoOOIOVzYN/v2zCufTF5zUt99FYbNe0wV/LT9mNMqSNSR2
GkNNwvnwEFn9W7cj0lzxM9oW0/JKXPAZ5eMQRy/asbvM0UNqpPFIHiwbeDSfk5gm
RnvvdCUaN0mMwH46tZuS1DwP+25yCIi5ggdizyhMCe/4XQw06G648y+6TBRSHJ4m
B5VbF052xZu6FRMksAP1mAKdZIwvUcBeYiRvgUuD3HP9O8dzyEUWKvwA1KD6EFC6
uLf64WV5JqaCKajAGLnQvXgJ+zH3OeZ0pBayPt2a/93fiVEPctyzBlocqf92QN0n
1Wq6O0SezzbYhaFFzd2wE+pqj8jUUs5gsrSqts6rjExb70cGLat28KmC4jAZUPjL
U2+FksuVLwASqDUDCeD1wZAXrHv2h9jDzK4IthQLVPlh3Ece+CPl63iwenz+xC8Y
I+htfmjTzBS6i31zzyj9wFkgnn+oIqkhq4hbJoy9v4Ztu+VGdY+Nm0bl3fCDbpLk
rhhPl3gnS+XYImsygduuoQpDCGiXS+6Nn1pkGC5a+Oap35+pkMAkd3Vb7WGu81W2
IHubnCHKJCdMaHWhgLyLNnDsUZYDpvLQnPYFabqa415Z+DO2Zg2vvsMQ/4/S32/C
JW+dBRN1o+PS1QxvS09zn5dOtA3DSe1CRYLKapTwAyVxe+fq2ITLxpLoWEQFUZAl
UONs5zsWVRnBj/o5tRjvykOCxvFe8zJ+aDG3aWGJ9WCuXKs55ezHm73qoHZUryyX
A3zfZnlTagmaLdvvkkUeGPmZM4SYoPrlIbnw2j7rmtl3qWlBa7MQ9Znv4siJLzUv
AwjRx925X/3r5zcRiTr9xHg8rMHi1zqe4d2VLnTz4Athnpu89Cq+wREy4mI9MJmT
/nLM21MTDQhWA6vWjM8edELSx0TEbCMqRLawrQwmHPMc31DJU8nDn9ahyLCeFKrm
EJsM0ukw/YgHaUxkiIR/oAMLK0RwmR5WrFY7PAnvFP/47jE+lr5PBt8hJx3QjKX7
J0Uyyxn0N87XX7QVIRuDePJXwVO650VvrKX421yql1MCBtAo0rdM2n+a5PiFSIAG
40dCEV5+1zHAGUvGqUbXeC38Z4062xVD+6YyXo57Hv3cG/P7yyT2A3gRJmk2f0vk
gMHUYKsH9IvT1EIiCXfDxgfci+PoaJwRzEtCpb8Xtax6cYJaorqoSrSPw0pOdiXT
yCKNqMipUTVepkdhjR0qVfk0Y6Wgt/IP0oE4prbOiYeuC2WAizWERlT50gJW33TZ
7YGj8otl/AlqmBInlWHWWKbLFw0t7Gho5Jyd/7fDo5fZ+a3hdIZE0WyEo+J2mqN+
e2kHoYiWYE6JhQwPGcBZxCupYNKkU3F+Dctx/y9QdWeGF3rI2N0gS+1IbYuLF3AM
t/j/486yXH1r0LT/x/h4jHLwx3+JbO/w9/SAh0gth/a+8g0a3KSCmw+nCTAfVoPD
aiZq5A3GNvSHDuYiIEMI3tVNFiYAtSDfA1DN2GH7cmNz1GSjhBR7oMroSC7vQsHn
f6d2SYjqr06gPo6IxkQQgkNc4He2XG8GIAjJ6SPk/svT6iCWN+dI2aFTowsZ3MIE
aoBMlxPIAV9kYi+bo0tOvnLsNAEmIfvB6ceGX0LxeGenlI8AdGZBk0DUABRINWgy
YibLHHlWtyIqUzpBPuPKkKigTUdElWm3e4xTeZp25XDHi4yZ0pTEpkuRHDm+j+rH
CWGgbjjHcSMDxno0M+t55ToVN7V5AoXwH9UfEiwVFIsx3p6WC9AmiJScCvzgCxMO
tVr+xqvc2bWvhx+eh+NMaGXoPirZKH3dawQURUIW/g3Haq5cvmfy0RegJbKuE3tP
AOUhiGi/HFMOREQZLZ9KzBP3ybHnVIoIga4H6eWAPCAGWqgINKAuNCaKjaOL4iWL
/GpCN3IRhuyQxrR18k8LeynmBB71tkyd9KbES1YUF6MHnYrxr3c6bx0Ea7LNLF3R
0Qv+SRYyxKwZvzA6BnyhoUpr8HqknB/wOIaH21TlM+W6fpViEKjZ7vjmIBOYxx82
gDodGNBeh/OntXZ6vl5iX7Vl/8GvL/ssuoDeBDXThzs5iNeZwmhmip7Pu1ZSXue6
L0b9wScZfjad6zs9omgT+cTONNuCOzfV8uPEfqsKHKm3aps3b0q39iPS9Ndi4uxV
RIVt3PoBcBNe328XMt5r+3qOZi/BV53hm2VfXj3/ckStFcRiS64ytez9YC9DXcf0
5wPxQHcOUZ2zQp1PUvURemUoDmWHgZGdE4LrNGXSsCEcVMMwkdxA8j4OsDpF/GBe
zfJ+IkswH7LJKYwGBAeOHffOLSDHqzOzdkrMM7VBHgzgkpGkH6gVmTfa1x82IChR
7HUmjl3qnqYYWQ5xgmXKlzCZMjJIcB3th3HPV3KLV/+hLmpTvYx105ar5AZkE405
X8DjGk7d0b2NI4qvHKrHdYZdMGfhFF/Lg3JmMMorhBPaRy0QyRorbRF+PtqdgYKF
9eri26g7ymmam1iearFulP0rnnYKB0Jz05mBVQUrsP/4WAbHjTM/1GHYqdl9alui
4ZZHyfI0J9VjwOYSEv9xxXlZN1HHHW+ctG06MPI0Mkyp3NRy+isdl1noxO530PqA
5bzexC31B6jfXF3RIv2YHrxfuB4mmYZVgpRJwOtHspmKOipoe5Kb41eXxoMQh1Vm
Ue2wMgIbpvkCx+P8QhRL8OrBmbo5MYImhoFWlCk5fqlu2Pg7wfuwSP+nIzmkGT6b
oAUTkAd9xkTiBVEQlL+5y9E5l1rXQOoNTafVFr9NyIrelnQLi0EFcAgUa1bGkxEd
4nJ5TYfjjTaDt0l1zf4kldvTVIpCexKKxshysYKoZJvm7qUEu1L+shdGTxUE0gej
035wkwwy8Q5kz42njwE8kuD3N7kw/5EYKXjV6aMPwp92C+BsoTP8gd/DjpOCXIfM
DMABSS1Mrs2Tlsua0redYvXchv9oeJ13UJ2PRrS+hya2g88KU5UWcb4225jT+Idc
uz3TNlbJp5oo3p3BQc9HP2mRJ5LrN7SFwDajN4a2gnI+F5xHmqzkyeGsX1JAM83C
6aJA8PFjoIbSMGEX0z8Ymqee4ONQDK12M9ejSKxxCocnAQt8a1/A7Br6d3yAT2EU
3+mrVkBpLIM9BN0h44BFwkf7RmgL+mrz1LtFJ8BDjeWrKTw0kZNNI7ei68EhpXG0
GKtzxCLD0GXVWU95CT40uHhAWalM9u3X081HifZqp3MAwKyBX+J6Ig/YqPC1zs4Y
6j8fs13rle6qlKYqrsRuV9+bzzZmRv1QTaBddAfXk4Wcfj1qp2Ov6BOTrFosXPFA
B0hg9XoxRzp9v4NqA3vwORCAjHthIEgULL3b3K20QXWKTL/nTYu9pz8/e/U9k1vw
xjLxx2cF9UonZQmDzcyJQhZKd5+oSvzoWqDHU8y7/oNa4d2iqXjJFKLZSow8EM9u
HdgliHO2b1hqUZWNaHxxa+nJZ8yX75DnkJ4J1lQJp3txMQxc2vRTO1e48sDBRQpW
8yVEI02Dh6FCq93EMcJvDF/HCmzqYpCPsrQ0xAoACqX5azM/2XHP/1X0XtlDzUHJ
2BQLTjuiMtwFWlt9rFtc1nPAigfV02YYnXSxmEXBbWSjlrNirVqADdY910HsF02G
KMdrgmVBY0aHmLuhF3qpPkf/OVWS5jUegOgnaHfWA9cYH1DPaP2NXHjl9eTVnZCl
qWNfQxxUlwo1cRDV6WhxD05ES50a+gFpkzjSKabxIe8Ppbzv/7VnBCNiDNsmY/7w
9moABnC4CDrdYyGtkWNZ0WM4D3celOPRt1FUNm0shhwtqULtw4HShzu6XSHh9Mo9
d5slh0NbEvJoxHF7nmgGmRj29hbtO1OPXBKUPccKasMZt1ivEvhRNPOBgFz/Tala
npNAfCGFhZlknzfgrWz6gDZ8M9tOl/ks3n0gD/wXmXuAySisOce0fU3Dn1i0yArH
xTcFQDDn5FbHsSfzoEZnGRA3WsX69v/rIdZL1mtoHFBaVk9OYqBXRXDdyCMb9OHR
M9326oD6sLGWRGJiP/aI+xZi+UcQwe8ZTZslzw8qTDvitFVepaF0Jp494R3O24vJ
BS0IMSkCCX2oupNLtCuIRlG/+kCgSgg9xkqSI29pNa1xLayVGQ57GLhTwxVzLMKT
JIflo7cP+9RQsfT4o1cY9dm/2qtDPH7knXuaz7HXmx5epu+OKNYlJGmogBBmolLd
M49lJIoLoroIonmB2KCxQijREHZNpcEzp4Jt6m2eVuqb7giEPOXouDAj+uAx/0tF
+9ePpZCkoaebVqa+Mj8AoxhNyZ+bm3PZC63sKpoM9OHQcj/CIZjmRkG7doKIh5Wd
mAWYYHbuwPicIg0RjWQgc46GOfEkvqpsvvtuBLDC0sgmaZh3ku1OPxSTz5LkPwwa
DT51LiMSVRswXTJqY07t9qvzcJv6p/ZOZOpjJAigPiwiMmpvJhANCGeSI4NxWUnh
Nx/I4+g1ogJeoIaMEwKe0V30hDw7YXeWG4TIYOTxzWrii1rBpDvmbydXmeD8L8lu
P6JsTrq6nX8PROmic7YCe5ybRYiQBbAZAKLYm6/wLHv4C3cQdxMV6qJ95UP62+7b
NsrNkzzTZ7vuGiBw51FavwDvjQ+odF/Xjf95Wxd+cleIK4/RZPxoULUSW47CFxCf
xap2mkmz+MOPKIROTLcF3tTviO/78aJhppELGdlwYq/baGf3s/oNCSRr71BaTeqk
tOGyrJ1NsOrnNy57hZ8TM1AcFCZMdoEe7kkKBuJ+HJvXxi/XzkReLBsxmbguP96G
YD+jnz7s+JgRSlJadInX2JzOtiFxwPZWpp0KAny82A6QJDqSpy46HKwYWxYzvbxh
C1NNYQamLpsGbnSOjMpkruVQsbWwQb4SiGFD50LNUfx485VuozPsVHHWolZye2kx
6d/mUN7i+YR5nL+jlqegPW2zLFvJxTwZzhH1svUNTYkGnxVdsGaPRe7Iyos+h4o9
e2Ze3X4XFx0WCG0RRhslkbOKArg4un1sIGJnRfSOvdj9BoDlI42esGVE+frj3ERl
rcbCQqTzX/rcQThmnxfvJ75IB0JFWRUFihzMrI2mNKExC9j68rzCoJj6/ypApv6w
wppn3pT5L9tstMsPTYQXjY3Pb3VVECxdTuW0bIodfohd/owjrCYN8X96tgoOzU5e
d/wCqFOA2M0XFx2fonGLYDxDvHe7m2fenonqlK1pT6oRqXCSsjNyl69HFjEUMcmw
nPVEzlk6hXOPK59JbcoGdSbzN+3gUJDl9JClT9kKcXEXJvPIchZoYijUEYWx3rto
goXFyUyr89pShc3484ZT4ismZnc2+3hBuyL0tYeUyVv/RSMHMm9T+eSfDzXOtoBI
VuwRf3cdWVqAgVGMWOKZTrOsbt8kVqg1jQ+YCJZyzBC5J8HHhEYwMqZdl5sAG3H7
3Aze2f4BaFEvj+hecER2pjoZKVx7fuZbkt4JxmdeoPq42bxe/pbuNvLAdHuqfBQu
PxLTK1ZlqWsinxB7M3U5OOeXSNMRa1WW1PxtDYMIE/boFVHXPiJaehbTLKCEtPqs
5RWBf3BbnlhQsed/dwoYh2QAYbkIpT/uXMUmIkzjDbXk3YwodTTYuUr5NgsDaIK9
S8G61Kk4tAOhTD7+0nlT9oh+OKNWdjseW/aykQ3T79oijlSIHc/PobZR9PhHCN2A
59HIWyDwrp/eOP1E8cqtDikhEFCWagLu6qXCTIu1kyorWCoufdAYUzcsrVKepJse
cP4uMLm5m/nX57cpp+DAbfnQdcp8cWqvrX96WMuPBe23/v3kghj69yY/fN68Vegq
YgTN2uuIG7zg6uMCvnDhWTz3BxiPE7zlp2M0K6ot0wumsZnu6QVFcZHxBXk7JK5d
yFspHPRK4p+xlP+Ps5ufC1giO4iLZShNquRis2Y0gucBvQ2WhA8nNvbqprbTnY1F
GLbdiTMlmv6iwWXNn0oW2GeAXAPBvgemtx+79F9UlcymQjPDWTK4M3BxHGJ/Xzml
dFLLPFNEpmc3VyKq1pPFLuOHDEmpJBJB+OyCu6+7a4DGfoQH0LH9nl2WR3mcVOM2
SNy9qudj0yVhSTYlSEGy434H3r+ypiYezI9nOm3BQVYVU+047cTKll3nFN1mGYtS
GufIheLX62MumDyEc86RXCvKHwFEVyPBcWTw616tLYXTpQqaBKWM70FMQjHq5Q32
e13iBTihIap254UgqdZCJKEzk8X5IAWhzZfzEq6Jw2sfENRZbzYd1/DEXFj0I9hp
V6D5YtQRjZj5H62L1PU+pnM9Xos4TtNyvJg+S3bD+zmLkk2/nPPMHor9O2K0C1us
1EpBkWnMX7i+sNcPB8uveLNFmoBbphpf5gSggeE8bRF0VT6Gt1DnUyBuVMZwKACj
KK/Z/hg3oytjS/Ois2FPxgmCvcfgx2TRwIga22O8BUAEu0tNHp/kocdoPndBZjyo
9L/F6eDa1ba+8fKbJqOrR4Daw1L6sX6qdD8CY1BJCaO8Gm3Zzu9emkiwA+rAbJN5
Ne8tvbvVbNZy4Tnxc3D76y+nNJ5/7/ZCmRzcYYE95stzf9sikOoksL6jo5/4syBx
Nk/WUDPSxEdPKOyb2kYtnCAkeCa/CGhDL+aQbqRoexhVJfDl3SCQHbQ5QxQqxLAP
83XoF2r9n1PF+c9lmtlf8nBp2bTME5c/KTeUu6xftWENnUeyXGin9/NUYiBb1jnZ
YFzX6yVFTUNbJYRuf+/tkTX97q4bLSm9W31orLGNLiww31wefW62DfKqDxsGATgA
KjxlCd7k6XB69tQlUqVx5QlagXChZSLf40X0LKppW/ZstI+GJadULLNc+mP/KMrh
VwH9Pr26msADabzEYazTzPkcspGcO+QSCsHVLMxDDBLoOcdIymBRI7DAP+gH4M02
yD5uITBwuMsetnTdhfjHFf/ry6zEAev2KL1YBQPORf1eSUEw4lpiBEkNE+sRnvpI
E1YqJLqYfB6zQKVO2u5ec/EX2PrHQc/J6Hj6eIt43g22xH0QGUd6fv86zt74cDOi
FNs9i6xzhSopMi+4IckNAA085GLprOVkz0MO0ZcVcg6tWq2P/ugdg2Vl9Z7wAWqF
Rc2bb1e9NB9DtowRimeQiv8fN9m17YSbmD/jyeigW52EDoamhwNAHt8VvHyyupuE
SxjPmGLF3lVNolDdfd0BgK0tiPGvThBPlOXN7lUB4R3jmhnGnA/cu63tn8sVYPKT
dozhM3uu6bYwywgL5UiCTzFZsZm3ikePtDXdBYcvGsk1tDPfaEuIoqnKGRyCo8GR
aHtVFVFxV0a0kjv8V//j/SE9aNemTp7+lsh+DkeTRlF7K4AYTUDTWXl99BaGeW3G
Wd/AJk+pzFgsows9mQz/gWecDyXA/HVKui1kC/hZ/6ugQYVo4l5Gl8HcHuD/NKCy
QItGj+ICCaniPdm6EXaVSpaHMblQpV1gUvyIAD9YU2GtEjh9JblOuprJfBeuVzHE
zATuC5bd62zNkS/7+zsp3BiwbvYgceCJ9UUTl8yQ7CbCXNu8C/3J6+E7ZXPstHqJ
qJh+W3hD+IlgFtLyElT5JSBdVinbhYtBU8YnC4UbJvOgFWa1k9nlRY1xKQPSGPvB
Ac/esmLIrSLlsMIfJu+vtTU+O7m7x3PWmCQqHb5c6SKm/O9ylqWeeXHQwF4esQ6C
FIAiGdXX64jYcdl3Z9xTKAAfnw5z6Xrwe0OA7tnywxmCieaOXQd/KGUzbP508ZEV
iegxSkkdyfv1PUe8x9DxXQCy9LMnpKPde/7Lmk/WpK3lRl/8hD5n+78SxWfOAW+U
xctvGVTWccWd/vAOUWZpcqWXuVS75OK9ccMAy6QFegdC58/gxQNhiQMcfqFtWmbk
z/0TMGvkooZKqEWbTPhsKgdv1BQWGFkSwbDu82O42w1u4S8lW66e7l9X8IiqwUvN
Z3h+EiVQGCORqyb67aZPHSAXYdDZ+81Q7xeqR7ooLcTZlPeATVgSHWKw7CIlL8uh
IJRFMQVW0im90+FHUITJt0mQBP7s8vTFYqAIzOA3slZDg/l1NNGMAWlzBlXVro7s
B3s1oU/wjOUnBmrHRYoQBFoEHcCQiCVXBf6+sG5o1jB/AkSqC5nrbJC/mVMwh4tI
Pp1VYxdnJunFz+ZPS84ENw8pE56/JEjdPil67vDDb5tgoGmfRDmis8PkZ6zr1hXT
hNwc3iYb2eoBhkZqYb63ZORqSw+j4JYdW1krz7EgL4HzQw9eetWWW1llyO8y5ISJ
t4oP2MMNBRMVfc6QLPFhQxqZQYc37bUb3nTNR962WB7ENeN12ilbkw75Hc1e2OCm
58CLMgpx3AxTiYc7HCWXqw==
`protect end_protected