`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6288 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
YKazAXTwZvVeXonKKI9l+/wvqHQ+TFtxpoxllDMI7RfTN5cHkZ/YOPJPerJreCmX
eHHCHA8t+lqyawBg8vyODqhPWYn1Yq8E06mHwXc86Wf7AQVaz3hlPlEGbHuEFbaL
Lb6q1drgYMJa5q/usA1zTfRgDLhJTpfreuhyov3RRke1RTd7TMu6zFefKF/n32gv
fI2LGvcOkiynj8ukodohCf8eCBQeJq+qddFSXbTW2veWoKe3Teb8R754oNpxNzrN
J1Tv0j7Mt/Lg52nbNfXjZKywXsCaluMTzXQJHCctnf+6oW25SKh3Do2qm5tj8hbA
Zliwn7ND4B6HmtQZ39pQycb2p2s/xw1BcjV+7YXUGEeWuoHlHU6RBUXBWI/9J5QY
8qlacIwt8dRC9EifB8xd5y3fptFP3zuLZCNgYsPGML3NCQt1y5ncGHShgcb+FfQc
JDRKRZZun1aZx0B5q/jvuf0EDTyiKF1h0IfVP1r+r+NMeI8J7HOjXVwX/LELB3fx
026yV6epbATPMRlIeRpxdGO3z05biKIbYL6ik0PQSq+h4dHS5yfjpFgFg1mJIo1w
hDXr9uvlyQXvffdp3bnfoR8Sy4S948OiyEo8ui6wbBoqbv2J9tna5l5OeE31/LGh
nDYLHBOSJGwjD9XAQDL/rQkoCltFp4aTE1KcUb0TT5hz1KGZ85+k4+iP9c8pp3JN
g/hUZxK+2OwA/Qvyvs11GUBGtOIePOxIdqcccYqszzYk66EpSV6e1yJd4Qafmskh
w4baflO4jHvSZAyR2kA39GYvYNzwojIgLhP4Nnays5OhxXWbctC4+bjb4luFIbvv
uS0FN2AOWcgE7cR2YUwnneKRkCIChzBOYzcyR7iDrXxWgWkY75Q24B1R26fz+ZoN
4fkbUKmAmAaUtH3U6/kkEt9Y4ni6TM/ydiYYnHmt2ShASBuuG2YgDaD98YitdKe3
mM6T+04LQyunOZjYCFtBXuZG6Qv+P/LKa+5Aec4DNZktZP2+pGTdV28X/N7hDqlK
tvlRzD4yMhjNlPscaw41MIY/6sFEDrc0GoakyVCvktvOIwcehPMNiE8IL9yt/pRY
uiq0bOd30BWIwsBMIa+Jpc2ESyuRXPiFpbgawZal2/jXNeiVAW9zBpiYATW/uz+2
5m7mJnhFmUplSMcgTDV/1inbN1Qu2N1MR2CV+R8vnF+54V6m8mrfxqUyhYrFtJg0
M9TWhH83xmxsb3jivpaNm/YFramlk7fODsKlFwwFRD4L95sRxwgSq2DrI62mQGa4
IovI0/6n6MhrTAus/OFb37+SCJnh/dxa/EqnrrguVE921uztnSl1dzKmyp7VK/vd
/Ph68wU89ezGHXbzeN9fGFdA9OcQzNn9/wE29k75GORAoLjg/dOHly334fdT6kYR
V0U7I7lYB03/W7YFIc+8M4gTR3rK6vtjiX+0gSgpl8wvXc+d0gtnAlVvNY7BqNhA
nBlliXDswOIFg2Zcl7uFVRY6ZNmI7majviUlHZ3zxXW9VRBrJ36/79oJO1wQscPY
uslC8ydpLADVy9NX053n5cn26H9Mps1mHbgGby7dZzLpqIuL3XDFPzATtn13Y2rO
IuMk46mIULG9hdMLROSjWD9pdwh5S/67DnwEMOeaS3yC4FxOu3yFsNUR48KgCGip
+4BqmxuTbe3xJFGM2p+4kuo3ZipyJtJy9eoHc8sOo8G7+fDkSnNnuGSfVwIPXWIt
dcH18/E964xNhUC3/W94uyrgrRyIEdfk/Ak1XRRUEBfRC/Ei0qE3FiCtJnPCq7BK
MkYTlpA5XXJcC+EH3GNGmqirVqH+Su251RLRoQ8fmepnv3f6f6tWup5hwoXgfK0+
0G4uCAK8WIL4MPoVeejF95CrA6+7e3T+pLBN5kx3oI4NmR8dIdIAAL5uv2Ip6S7V
3zqK7zDpm/xwKkRSpZx7zAo81LSDBBHrwEerzNFScxUwYKgy5rAFp1Nowy+p8Wrb
zlyKT/6onOvFlJFV5HWxb4EsMwx/03kMNZ0p9JpNqCzcjFOd4n2JW71VrPOhbLZt
onMfu4ZP3zGM8N120BIOGNWMss+6Fivt6ViJYoLkkE+jn4qsPSNIGOtvwMXAErqu
xmWzTVf5egK8/ALmusl02R8rXOhG/1Kkqo4nH3TSid9vnffkf/51FzPggiBaFA2I
fcTsAMJcRdCpUWdBv7Z99SovzK9KPtJDgCS5iOnLX97F1dxP6qpU0ai4UEOciKwK
GJ1GxqcM7HwLVOTODh/y6lZ+xrck4vQOPUVww4WJpvJ0APkJD5Z6R7gZltloDSwv
LlWT8hYZRr7PF7OzIs2Vae0NPhOq0XCcE1Sf5kT2t3nPScSinMdzhkNbi1cuWwNH
SvVTHm3JkY2Ts+OiqpdXV4v5CEBbOpO7hwOpCSFF5DlpD1gkc5TrIaqDnkwx2BmZ
kcwX5LBn4QF5HXJ3pJuHklORpS0TTNLkLjTNUnsPnlJDnFG5CDpkYJd4WqQ7iRdv
qPE1/YJCOnILPkC0HRpx9AfHba0lGNIJPlTd0/m3IonttWHXyOYE91EHOoYKNnT9
d0YCtOL5MwLDJX/I8SCZvhBcEWH/krDRQDwCNlwHxtd/4CiaDZgr8JQjGYCiEC9K
oARS/JUNwFX3hbJD56jdv/MPkPk4+l6hdZ2suilAjeMm8BpTeNDgbYmeK3v7KN0v
Y0wqrKd0UTBxS/jQQx9+x+DJOy7Ros28JCu2yMsSE8QEpbT0RYBn3eT6AW1bSQVj
TRHgScgZC7f3yqU248UX7t1KacCgQuuwR5DgIfzU0lPj6XlelDko4UG50zbwiukX
mbtFrBvgXmnrGjaPc1AQ9VZviccHVYFrVKgdd5QUviqeJyPQEnNhiUE5bBibJHVB
y2Ea5fMciQWlTx0enj2gtymVK+yOQUCsDR8BI0D3RZ0uEIxjXKEXn+WuweVBgclj
qb8RvbZIO2hqGhwXmlN/r7V1tALasp4d9sR4nS1SdQadbbhZzDBaD+iPayOyZPKu
M0yw9S96+lX5AEzhMPLyhtJt0s6I+IvPQbInqHbRPDA+k8g9yZ3uZxJ5h6nU3R+T
MZUmhgNooszBcxiEeBOIIRzkMQwaK3IFlQcfqdhjpW6C3567KqzKIBQqVnBe1uBp
v3BiUcv5gkiJZxO4kzM3RmlCt5jypTIxsYvsK6Z06zHhWBJ/F7INNPRniWxkzG0h
Fbp9EbGvW4zxFui1V9S/aUMtm1+v/WszfBymRt/e8ErRDLmwAsKIHGoWr1zA0pZA
KPWgywFRggFyyKzYqkRLPIO9148a7Tdfdla/Oy94PLn0eu5PtTxhHC6j4SdRBMGc
aw99dOUjJnFROQgqIc9ys0zoejK/D6Ldme4J9abFZWixxuJfVi70cOxCGDmKNJ7E
1a8qUPkDmdpMXu/kRjrjx0MtXEwjtJYy/ZxDoFCVAEVzmufP2Vn1qW2DWie59J6Q
T5kUcvQiFSIsAUTV9x606ekWY7ULJlanUdxw7uFj7TbwHOgBVeKjDki4cLtKU6kc
qeNL3t6zJsomcxgly7CgNU4e3frBX5XxaZOb2vTa24EIhnwjl1oEP7QtxKOW3pBJ
b/kaeKz4RsDph2XmC/WHW2C6OceeacqcX9V3GXyVa1/JhbDlbLoFvRoCyPoWvLXI
s8MdDpVt52CQCqT95K9KihHmyQqRdluQJyUdfv95sAVXLI7Gpk57W0KYWGha1pqQ
/OhXNHvzSSdB6hK13WmN5S0o+VbWpUrz76ZGpRsGulCPG6H4VriTfTLKlSuE8bJ2
HoueIFTNxMC7f1F3jEAuCms+X6HBSXVAnG84HDRmR0j/xtsSdysxTtZ4NIoiQ8Pn
aD6p7Xr2kbhIyiNblv8Xu2wXwjKr2m6cFgjyYy+6CyvIXKh34XekLWUt6qydcfKm
xrrI5jnBxuJmA24HKTdi3dHKNSfNN1HqGJFhSM0y2M1ksV8J2sdPmG9HOTwE3ZkC
Ue089DBhiAqUqikyhq5DqOQxGYOcsK9v8G0FpCmSZu5aTHjoY06wOXw2uDlYESTs
ylFErtuW+nl8me8aN49K1rA5+7iYAyFP/mTSWsBgzffmcJuHiWRYs7msMBM6RD/p
gvu8anehtUziC6oycY6pqQM0ws9eiyZXiCdZaksQ/ud8v15yL6vVJV6wk3VR0dKT
H2vFbsmjPDkG8mdqcc5N/HJohOhGU4Qjgc1348uXyYwprfc1e63saNlCAnE3LbtZ
avOCGwlPtFgRDcK7qNrCnKiZx9LkA1v5kn+zkAJXw6aqcCZlhSJmv3UbARdpcUT3
O1LN606cPVEC8pGc2KLzFaUUAg96iCeiA0rTQ1nQs+GKkYyyUbrPen59a3g2I8bq
kA2ZHPS1lbWW+opdA/+WVeq5b6tSnFwye02sGeXb+LziSQlt9A4KtdxTkgO9yqXQ
sRuc+alQ2U4Kfm+WT6XloX/MEAlR1xoQEE8MXq+wGAv1SqBHuX9JgA16+q6/Y4+S
lEcr1wGBCEt8b+zrAy1/+mlFSEZfkfJodVEOWMfjc3XSIWv8OHGysRKWRAfZzXLw
7TRoNjCdoo1lLrBIzCOs/08nYRcOdGDYHMIjWjjyO2f4HJ51XvTEVyTNMx0945CG
wcZAdElVfr6SISW5C7Jol0BuCVuWDN4Wondy5gNgwawAS38eLDlXh0LV7iSwGz4q
K0fJ2ZBLto/nE57Q5Ggt1gEzl8qUqxaQsfBIgzGSk2dhjOvsTXUW5lK5iITXOo/0
7+mXu/6E7oVo5MQNaAhfZbOjnTam252oC93yN1gK1PnDIn9JwQA7j5a0GsNPHuAO
WO0kZeY0nr5cQLbtl5LBD9rW3OGyD3IrYZkiPspSnGaekaiW4X2RR57yQ+FAJK2s
7g/qbCHzXwG+Zs3NkBMV+5nrkY3AnclR0EB57BWBz8sgBdQL+gs+I46jQ4BBv3wP
V8mymehv/BYR1bWwPigtEXcPs4Dpad7FSLzqbEpzeBYOCfEK+yTiH7JlkromsASB
NbhWWyCqs+nfAVuKSZfbqY++2Kf85SpzRSlxuKp3M9o8RvN8V64ZnRnicFeGgrN7
1MAq8G12mUvnmokpTiaygp7fNo8NHxfVewShQ6vPAxASsz4N+Mz17oxhtFSZbcwZ
ATxbH6RYPy6hNnz5rS0LXoNjW9bwP3kNFPbzEsnZhf2RfmuMn3exZge8OYOlhFou
0EaZe5OdZxp8b53394xsdGe06mhihvyKQ+c/rKRvS1V033RJiiS4YVJ7td9zc8zs
hpZqT1iKCahc+gTo4iOzs2BEpZkpryl0gAF5gqzW1Mh6eh9nFcXR7jeXTkxDo7Wp
FUhntebsH85xARadjppUkBqLiatCE5KvgvgYmIShIZSjmj7B+sMj9Eo5hr3Nn9La
/px1RYos+yU9K4CxDPhEApbXeAcd+swUiMC4UU1wF5rhed/gDgu9nb/ofHXL3G/Q
lYCdrwIlLUB0tf113LlKvAtLa9ZqwBmUblR1PzV4/OsVbv5nk3xKKI6p6nq3boTo
wjXMJ9qeQhiUgNeOZ6TSuISpacP0NJHrX2NteXrnRBuwFwuPlNfI2d8DLSfi59ig
35gI5Ho3zyvuOr29dfteBCXay0WHBzzROHX3zm8eboL0DKz1RVFFDfppumvldUoC
P28UBq8pLn0/uDQ8oKEH1Ta5NnJsVU8+YiughOHdNIHDhEtCXQsfJgPzT5CnhOcA
9GtBqda+7GdADyj42n1vodoHb6CYXJ6wrUS4aRMk3ujTtTCpCrUZwl/uZOixpZMO
S0nIgjNkKnvfYnYRt0XzBfXg7F5uRN/dQ/nOm08ET6V9Mo4Su/ILjsQKEhONxif4
KAaoiLqtrxu9g/BJN7F6cTbKR+B03NYe2sjBg91c2zLQvLsQSjxOB63nOisvsuNh
OZoXrGjYFRKiGz8+D8QPi0gM8wMPtBDCbEWoibxwYohwepti/KqiBn8Yg/PoOUrj
cnYcIsC1IBiLzsYON0MnmkrlDGFLPR+q544qF74MmnJpn2WRtX5oxOrCMQXygfLl
vdBlnlY/K1zMraixsPsOwbsvpo+M6zM36Uvdb21wg1b7M7hvnWPdJ0XOmexebEXE
mOWJ+++GJKOGbYwNg+4k1kNKrVx6nz2mdQpf4saOCINuHbHM3S8ReSZDKYPsSQFO
fr/LWnFm5PQ0b2xlh7NVkp9XEJz926k8x3JCUmTNKes/BIo/cNqelbg0iXtVTxEd
er6zgvDGoCLtCKdkHK3Hjz3w8jhmUtTFnD7R5RJuc46VRTh/H5iS+VtfEqQnnB7E
5i1sZjLs1ZczaAtn/6HpUgNN87aMUe4njJNTzEuJrH7kzdQseMtrHsrZlFDoUY01
PU7l3/aMW/bY/V1lCnIXQUrYpPXsei3M8s7dq1Sdh6+NwXZ68yVdchcqeGDybuWH
Sw7X4IFgkgr1f9zR+DvOjEkNMn8K5penypznvsPtVZb6J7r3/5FB/Q7vI58NLBC/
Pm3oyuwGMZAmDyTv5XJwWHMsRz0tyJo7Ykbqgt4jj9AIVYxd7ZIEoQIPt4UQXRLt
TlBchhizuKoywaF/+lxt4gX2tyAMkvgORu/2tPwCS3WEBABilAVUZz8qiO6vrFeF
fSh5eJbm/lFIcZ4QZttcMhF5AwE+cYU/kYnhuX2LjOvrCKuatD1zn5i3a3BAe7jc
SthWrclGYAnQ3D0sNW+6kK1txKV26laeNH7CVssiTwSqn5Li/A19WX/4aKxc7/sM
z4EY1upKzz6miU/6GQ/9yYgOiIqaPUXWU+sn7LwLTh74Cg7RIyRR8x6aeYsjRu/D
7lDXPuoYykER0iB35RMOPtRGKF9PyndEko8ldOqtFEKt9CYv0pcoiBYVfUW85kY2
zYqKkcYSeH2KYeJuE8OXAheHUTHqd1yb9ZWA483WG7fgk94z8fvOOIiD+g4Ho0gI
4c/oeMFR974cclCFy9MVoBQGR1ymN/LZ3yxWMwg5sMhOz3p4UW5FlUcuulWBDMyP
EKUDaCsYq7dYkZfSP/YKuSIhR8czCrcHQ3Xq0EofuXrtjV2gifNyRS/jV/mr/4Ou
BZbdexkSajaW6WfT/ksn/ynTl82xkp7hCJdFRSd6IUjtbsBgGSvzuRwEvhSOI/SH
B1Mjs1O3WjMg//cSUG4OTovlryUz0blF0EcjfP8xQYeSTsevKSf/lseBoN6HPuqY
jdAoQZpHAfpQw8c9uvlkr/kegTzxJZGZe82CUoP8jr0rjkAX41XU57+VQIMCAU0X
p/VqDqNEE9IsI7q9oJYH8B6xVm6E4gtPhG8PhYtyXj8vC8bzfXy866r/yEady9eo
nFQm33ho7Qe6JxNFtvvDRN7DcFLvO85vLRLfdNcsFzB99obaXhu+9hAvI3cy3Jz5
XNV7GOr3tJMG5AOJo54fDNlKz2KIqigCVqsSugS56DnLtXLcM3qHPEBxPhB8BOZ5
ELvW/DinSqRWyr0rejYAdsAa6uEbVFdt3O1SjUNiPD5SAhs4mN868lTOCiZ57lKu
/Qw2hXhtmvBsoitMdjG9jaFJQ3RLAHCzcQD/NPvnyKK+IYRsNQ06z+UvAwz5FrMG
8w2dyesJkh760GefUEZP9TX7hpHDX0+RD17LeoyEK15IvaOSSxaiM21gNPL4GBhm
66BYyWoL6fJlDgUTxq9EmV4aG9Jdde/nvEprmZwVPf+Cqksaj17qkttoJJxT09DK
liXJ3oWFKvlFN2ouAx8VSjIzPRvEPP0tcdc/4lp7jW1yGVFZA8NbKudYiFr4bJjy
KcjXEL4Qi44v1PjVsZxWa6alP275kk+pus+LWEWe7pvLApngnKtD7hR8Pdfo4lFn
+U0tM80dtO5HoZjDXMqOaEnRfG9Dd7sDTwyfoUwQdnkW9QBc8YI7MhB7HBkNHxEH
MWX5pmXQqcVVtbmHaHpMQ14ebmK1N+fPyzJ3CP44zRFGsZdTgzlKXMAdNoliv+Ll
ZkQ9n5LgH5KCUcxniwsjv9q2VbcOmgorIr4A2UvUVixtL/rGADKl/QMmMeI8GknM
Y4G4TRNrlwgml4PWkM9jCv11J6m+Sv7K5xHkLV6TJrr2aRvOBBZu8OHojAO0lDBC
7HY1Nr8gOyYjlGru3uBk7U8IntcFhs+MF3bP/C/CeNAKHEdYZNYfNff/2WbDf4ke
YdRGvjiPy4LlxFKN5iAdF8X8OQXSnCU2J9VNsqR61AhUKsSjrYbkc3BJwfC2o2vh
0WJIGcWXfr77fh/V3xh4mRv4U6gs6sQXofzT/mr1QqQUXYcTK57ESgI/j856GzOb
`protect end_protected