`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7152 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpCy7VfzPucQWBxxbAs+GRaiXDTVGuZKhxkqAyHRyMusY
fIwGNsEUSZTW9qszjibKIEHoAYUpqUr02PxvykIgs/813J3KpThopa050aTinE+T
apsNih4qU1sFzo6RzBmBB6eG4BhHjGDyBUTjYdP3eCyr/yql5sdenuVaOrxE7YJB
9bN+ao/up7K+eSa/ecjqiHF9Io0m0cS/ffSlR+7kgLNUFB7b1VsHuRMYZVFM3PtP
6LSJ+qUQunCdrFllPOnyxH5ZQFHbTAZZAMigMJkTomhp+kpeHMQNbmCqQvp1S8jw
IttDlm0KucnlG7q+TjXDd7N/Wen8AfZywPjQQbBXb3UKNwXdP3PxcDYzPstjH+gP
R9b6PFSXnYSglcobt+PSGAdogjFgMKfu9LiVTBXU6rbou+01mBCak+XSp2i/QqCh
CyucK0vfVVQany2LCVOWOw8Ml1+OMIvCdafoUemkXJIBP2ucv3sboThaDJMMYUmp
REz7f0C98PHKqmiidApXz+VFHJxQeVf1gyvpo3EhNBVJG8nPt4Eyp9Iv5rM2CReb
Hd05S1WBAJ3BALrov66Qxj5U3hqESloSvVO0Ml83aXbk0EP2jBjcj1LKOnQBgs93
iFgF+5PS+auv/GpNy3hK54pLsVnXlSLOsnT+5sfn+jG+UD8nyZHyCXgcBEd23Rs9
C37plSowUGm+5Cp5nPUEDNr2MO293l5webM3e7pEqP38uZ/F3XhhHp6ZwEN+8E0H
KS2P6VdNXu6ACXSoD6a+ZUcCOP+EX0bx2zxKr7bE4u+KCwlK3ZIQ4rCsnNUJkl/z
+wqHhAQ121O7pgw+hKLZEZ0MpzyeBwaAtJwAjHZ+JmWMKLEsq5PIwU3uqSV1cASG
K2JL+1iLak+OhIts3XepeHEIyBpiZAcM3joGe+UCuuIiqOgiwIPj09zuvzIjG67e
rfAxDD8IJSOfAPvWT62x6Eq6fZW81Ww8+NzWCnsus9uXtrW0Yh981mTcII9dbOEi
5zy5fk6sNkfvgcvewDevR7pDMfz4sZuAoMh87HxXhAM3cczqTIk5PpnZO4lyCgA4
PRhDL5SrhLDOQY5UUTO0xEeV57ZLyIxyrL0uaWJZfVzHvSYFojKAB0oZOpMKoSdL
MRTADm34wb//h3YtYA17wmBBf+SXBO93NHPu54GPg+T3YEDssKALG4yKc4jXXe9D
simtzhqldh/HHJwWyC11v03ZWCm61Ab4eidzfMRT8Hq2fut4BqByUA6Efagpp9tV
aZ4IQkskWEtSOKzzN9DRJlWumoVmzruD26/ECRoeI9ofmipsf3qvq+Hs+4SKe3ts
Xvk07IAluDhXArnfoGcblAu2f4wkIJGsX2wJdFb/P35eKdU0XvXwO/YkmmzTO2tA
rnWJyPJNfR4Q22+bQATyix8dOetICfkCquIdhOjWJPbScVJ75gfopHEyyj258vwN
H8sbqeGMeuu4/GPJuUCAjFWs96VKKvDzJ3AFd8vObQOHgMbzI6cm0cRHMPWefwcL
78vgBe+4oiFDd9inoNtvYHiUi5RHgB6OOpAqcCY0372GQc3mDa4hGdYwci4Y3usA
+tpq0K8ZMyibqL5VwheCbwHbbFe0XDBCbb87+/TbQciKCLn/G7kYW26+8nn0YR6P
HoFDPydH71Qe1k9KfVTKAHHWp0jZYrBTRS+ULoHxMUvQiICBVJjWLlG9B5eior6I
cbD7MNUNMH4mPTD3dwlDBBhJ8PHRKF+q2pIAko7KMJTGzC+3RVNIHcKfGhagjirF
0ogfgEyLh1ZSddABgFG7L1kM1ea1c9oIDGtq/audY0/ZRfNQDo9sBq8LMsOPDzCq
R6j3mYVJK0NdivwAkPqDC++LiQMjzayctfO0D2x/6RIX5MBjADQGkBbnzEVkVtMz
O+uHkU5OufCSNWer2O1nF/C19APK6zBOujTnPXLIo3l6C0uhH+nzHYrO5RhXNCRl
SH5yNWuO2hIadq1vq77yfwizOdoX+ugDMacLgUsg2bUS5rLC9jPjJdQfLKdjmgeS
507ikEkBw+5yXFowmx03QydnnppaVVHH+tvcXzg0tZVozRpGlP0bSQPSAOyB+ixG
n540JlSGsmshSD3UTjcM4ZMuIBeOjYPp3t+Ps9LsrLY1XuRVRbaTEVQypLH2S7oZ
W5567udribPLt1jf0a3oo3Raw5rZkYMHmeDY8THE91nau4Q0oM4sLuPaOFSMks2n
/xvrxyld18doxubf72YjyMBj+j2UYLFymIAM35zjTeDsSgJyH4o/h1Mxg1XAugkm
D67BrFrT28klKuO4odkDke6iKEPVV0yVUcurVUZVVAXtYuF+hl82BkShn/VuZtrE
EqauLbcrwjm/gO1T3KMJTkVVIPN+vu9jUGy671an4Ep3r8c7uoQLzjpdni2qziec
rMmeHZQp8FjSbZZ/npawCntzsIxHvu9kAHHYKbieyVUTQlr8bv8e/SLbhtTIt28f
qL1wB0+zhNkchkjN4TexyJgNAab86Xv9QXc7O2c7Lb5aRCbUiARohfgQS8BlKE9S
VZ3z+sC/wpkntDQ3ZclGG4i9GL5ZuchGOxw9SfwyvEqSy+JtWc3kETPoEAPwWzun
Rqpl3B2/dEYn4IpuFs6ICG1nlsa8dEgf7cUKbI1pK/umvpXzaZHQtYZ67QVVlR62
aebqNdJQ9enKwQMKrVCT+G9J/QK1VJ9pPbi7Ylc+Q5h3AvjKCcg3Ch8PS5yHpjqy
KAjZ80Q3sQ8H1tf2EmuMmPbZzD3/W0p9MKXHWhsbEA1HT+IuOXFcVK6y4V+Eijo5
AQHkis02qn+Nfp1gxplf8JFwccE3/TZAfblBNpEMtFgdhAzi4TFZAYC41f2sLtwt
WaXXvRNPh0mFEeVy74zbJgEeDHUdaDWuC7tZE51DnRM+vCTYZFprKkimt9Rvl1gw
grvPJin2YZKNyVko0kmLMDbY9MpeGbU0slOlTJ4ZHmlCSCqIRwVUpyD7Cvne0ny0
kYCI5z884mpHPn+PN9xEGROUoUHZEd1ZnpXnuAaA6jw0eVbFOinw7J0tkX4W1Ct4
tHn76SakkAt6ou73p35CdhMHtspVhyqIMOAyId/ybtxP5O1KmzAUtgq+RvWTaTJV
ieeKpyJCkvgCKpJi9F0jHKscfSljNXZZGxVaLCBOztfO/eYDzWjhM1Jl8Hxl4bU4
DhKa+mIOh0lcpMJBJUJOHGeeptF6OFu1I2cevi8FFG6/cbwEWwkywC/w/Ue20dxk
ciJnxTozgtgQ37OOw27agTAHjLRGZ06yy3egtQhpsZh/yZYUWrx3C/16UGlKJuUC
DgZL4cWbr/+sSwaDnXK6oCklouIRX444i361u7SnaKnLJvwtQ+vuCHQqNqDogwAp
A2ZDUDYT+OQvq+uxZ2tHern62d/tRN/DtfeuaeIj/tHXk1Au8CqqREwPPX5+X4KH
0fC/Rpa4E1o/yYqftbnrXx7tiRoohBRLk40ISlH3YfXrOfekZNDm3dEBsx+YAMNk
LgjAHblIUb8zZ1u5Dex2kaEY8iuMXyGUJsXh4LYd9hD8Rf2ujBBE/IHFDDjbImYi
H5abJKx39n6yqddRsR5TpW4iKSad6pySKUOmejOzZKAn58PDkubaPG7GiMFT44HE
pBBBVIo2rlveBYqMXb7RFwgbvUo2sO7Ac9wppcGq4g0ncRfXWRi2D8t9uvHDYsjC
IgmIfYctiJdFaBeN9NWdz1YSOMcwfG+bgvcJzXcLGsi6ApQ0PRorY1YheirLkq61
TNdFtHBw8SUzS6JXrIMRYR6ut0snn98BMnre0VL0jcYZkMQ9uHs3Cb9wv6wlsRUL
phkCKI8g2fEJZrRKQ4E4qPue1uzA8jOYTouasa6iTzYfsJTqYofPKtt1UqU//JlU
MAyuylK2M3eg0i9twKBb91Lb7UNv2Td2fNyqs2jq6KqD/ZEmdE7cD2hWxWJFIFP2
pgtNFOYgdavY9o65gxkHMPUtfxozs2CGCeIKpKoGV8e217v8soycd4RZD2/+XL18
xuWJxgIH3Miw+PP3KfnkEQrMKh9C+/8XYzP5YcyH24pMZx4sYjBRQH00sm3ct6b5
6963aKvhWkAInIrq+l/EmwbifQAXYcZFhjfoG+HYfGZukFLSWj8anKL3rJ/NdWJn
lqeqgqy1ajAaFe8+PYRCOXTG8KCUM6elldjNpy1P2HQ4PTR42VM6+CB97GWWQD2B
t6oW+8m0ZD1VYIZU9Lq1+UjQF6693T82LucKJk2C2DX9MB8fhNm/eupW0cZNGDyY
56b8tvzBAoGhNm9ZQac93M52d82XpT2EEjZ0XDmUEIWee8uT/A1dCgSvl7zm+EtI
Voa2mpzkJEOUb0vkOxsDLodpn/82OhSdNAz1V0wyHLs/pkOajqq3jaLxbSMO96wA
NHPcrXXE9ikgBO9Lq7hCw7aFR00kK9jkZ3g4S4Z6NuP0wSTGhsr02JhvtnlWf4eb
2SXShHFwQu6FIm+6XyvAOSqiRgMIghxQhM6LG+wGFz0a6/qAX54NBoHVTXdEJXbD
yim89P24rfW+i6TExfFWinYeJm3vWzXbOWbUEYpf7aQ9nBvsJYDdOtpe+lvWv1rp
MvC7+eLSMzwfP6doPgpLPK4dvvrW33hMRBAxifUlW845U/WEQ3sDtowiBpt/g2J1
9KDNJvlLnz+8qiXadKQwcLQSO/ZtlZCjtpRz8ajOld+UEcncb09wIBd8T9hRzFGG
YXcNTvEVRvvbgxLoq3QaNCzCXoiVCDmRaqZFHINMG3RAEJ8RKB9hybRy8qdvnAZ3
alGMvK3x1bcronFQPpYnhXCG7t3VbCWT5WDYrs8e5VLL3XWkM0vFKx5nkjATiaIP
vnXb7epbxa3MhlpgP4RoNCduAtZ+8Sen5JAhVYaluMalDey6bnkjaSU+opuMR2vf
z9e11XKWUehYdw/J4msJwGuAE9Cimo1veF6FtzNLmm+UwAPtq7Xtf2Qh7danVNEo
DuFs4DNdMuFRtgJrcAX8Dtl4PkHKI25ITFKKBjQShQieDxBjbXEUdDBSob567gpl
V8WCH8MLn9vf4H6wcBQCoLE9cax9jj6r9uK5vwzYAHeDuGHV2iQPgrGq+APo+aJC
cs+XlZywYg4RzuXCaBtTGIKOdhpHof/kcIN18fPXBrheLk9lLebZDIYiMLkI6OnS
HjEEJ/RHUWB12fdbKTADtbGDdfRTTbs0H8sTFtSVol5+paSXkmYUxD14j/xV7ABh
qTFRVQqeL3PgPpyTNjU8JmDZoQ3t2GmoPT7Ri+UJ0fz4CrCzQyappsau+QKCDWpG
c5phkLYZzbU+w/jBxSAgRLGCWQK+b1PkqGm9GdXXH6EyaJkZqGnCu4g8CgopXwZc
1Q1C9s4hNpB/L19YOAi9ApEsDM/qZU8TtxmJensY1ZmY/RK5w4TP5/82MhBvzVd9
UoyJd7C9wt95xOpBbTKueJXzppAfoVUvAMGF6tX8EGEKaEHx8f5nh3epXzA/KKf1
NoHKhnddvL3ABDpLWqu+ZAmwll0zTQzdN54zAxG1/2gJxtheRMKPUw6tONIxA+ot
sB1aaDpzmDNEcjxH1/rAUJCwGsURWxBUzif4KFhqRWHc+ULto5H07X0ZvJCf0JM8
4CR+SX/QOgJOHSKW0H6UkDucCVBPBZDa6A4LyLm0BcCItXANJ4sjxXknY/mHcWAq
73/fN8T5FVx3/0noXNfFVkLpsjXdMreWUaygF9ct+1M55YIBvd8beG81vwKE7Uvb
5IPMbe3+dq+BkaQJf1k+H+biOmOPDIUdRuFC6wrOtKNw+BoC+bnSyrKV0eG4xxss
3Bl7gz2mB+/keya5v2B61i9lXqWjBhN88PmKTm8hV9D0kZegSsez6xFz+ezEwXX+
gBvp8h7sYlsKHlIfbIZWgxsFpGVDXk6wxU6+p+VAhKCJncDO8bEgxbGtXB/wTsq/
+LC1kYbXDdmqZPyCxoaHt9uxjNSNN6929sMuLza1/8rXnx5ioRuoD9R6Jhj6lVHG
eP/4mV+D1kexbyZ+iqnQ1Htl6I6GjPLlAyotxKR6qNZsru8T3sIgNb9rsIJIQ7Ww
tyeMlVke9RjYMcPKVq6D1BDqBwdVC5wpio/q5vfvtW3VVblj9EPCsfdOVOLYyGQo
KpWFuy0hHQCr/5JxHMQ3SGM8CZUnp8l/vXClOOJxmgF8OPvLDoIYoQR4asfXYsSn
QWxG0Rq0lJZi7tfE4Ef26aA3uB4A0N6JdDDYTg1/obS/qUpsR2rRIp4xsVQcWO4f
piRijTuKQFepX+Fbx/+mpVu3hiFRJWCialMOBHwurcNibKiDXcHV0kCRHNDbYx6/
J7+x4btOiXaOql8hwQ9B4WaGziG0cTdWlvxoIpI3XNCpZEIC15gsa539SoZqagsy
1XrR43gDSSav9ZJcuHcGFGw2Tn/XpMCdmOk+CrgnJVaIFjfxQcVsGzm8H3G2fUNj
sX5Zh5lpCVX5rd2g13FkVF3P0HP2pRbpEcEYg8+78TLUSMBSmmgH7TsL4bMvcXnd
x7O5o5EQxt1i/vzCmGsZD0QbkM1Hz7eeeWQPIpyTSGmo5RY3rod4O4uIP/8E/Er4
3uE+OyVjN2Di7kf0TIM8ECAaAK6cBeMV7Gf/W5N/cD74Jd1QkoqRqFv8yhbxnbLO
MjMK6cpseDz6Awj6rdY4CUEJQyzXiqxBfLy1zVb7EUxRD/NUm5hmfn4DG3Oar/Dn
7ObLENGbB5920IPqsPo9ZtkBhLqLK4qhcx2PrXarGsC6bAlBhgUT+AEnfXMHsRXP
3slI2MpROMDRj5BNQeKrjGwHh76pmAmMFb9HJxQc80EALCxZVruKALWuvL/Szq/h
UpXu3Xj96Iy+LGPb3ANtHjz1PKJLFW5+1U1b77sS5UBUXNPZKwFflv5xHucWSf5a
3r/DSk5oW5BXMDi1FJEoio1kSoS79JSODC7kYDzJuCZo2TB3RzgbKKXtQBBy0C0J
2sZVfZjrLqSsaBH2a8tnKqI8jFfhGNL/J2NnbjTz/VmJ/X9rijLMjGi5CDhJMndk
1kcn658MFJQaR/qB+DOEETHWdM5O7dYkKU2qbWamMWfWsELHxWu3B/Kjl5GKjcmk
tZ+QvTsWbw/vGzsmUmksfAx1FCCcaY0/kr+MVa7UBSrjsrJ4D2HuQ9UZj/6GA1uS
RpI0IW7jmjpkw4rxrRGfvTpGp0wsXE981EGy8sCtBlbf1ifpOw/jJdjhCMFgWgeK
oBxIr1B0SpWH7G9Ls5VrSPlYxm4p9Uc0wWRsXDWlr8V5W3MkxSlx+1aLtwsjWEye
o8xLSypiAdHLv4+oC0rUU6Om/EtoqmQe62dFusP2896El5+8HneW5B0GnWEVYc5/
oxv5hrofgvReF6RrosMe6b36JkTVqiSNN2EoODyOznwq41xZNafukOppWbpQKT9Y
XD+grxT2FosiD+QAl3SfFXNW4orfila1Rm/AMdlH6fbImLZdOP+1NFXaNwmf/g9Z
ASEMOGFta/iOS6ehbqb2CCDEXBZnEBxsLlEtJ8dBi96inJaFKRq3z9VH5UHC+4au
eeJiU0r7ddLUEXcs036i+Y2Dtyt4zJX+ruGd9BQ4bS1bWw4cgQ1XndcNV7NJhy60
eXZpozTZlaVQqfSqxHsHLqWDXcd69p0iR3UTfwfmQhhCuFeN8Fbv7k5TutPI7+Ap
H6/4E5uAYTs3xaHZyMjJnz/aulgDf7wz09x8ZyBn8IJGnGGGd2CvLcJq/ZwjcuQT
wkEZtAYuFw4WDiqgr6vg7Ve6HlTaeFi89RjZf8kmbB24JtBDsmR6iJoM3QpdxgO6
3Lpb6ScuqnI1Gk60jK7M3ceA7AjdSAZ9jeGtrNaQFjL4cqqNRECN1KQQNUa/TTM+
hRTArQ+Nn+mGDmEGDORb3tPcWn0h9aqR7IVSM/sM0jAeA3Lz3/Nf4P4ML9Oqjjt4
0sHaSRBUsU4J7KwnHPngoImEns32zBsWk5dxLPh4FRU75ATWrIvnLAYFKYp8EOSH
G41UzyzUln0jAgnXivOtr+S9bdysVfNIrqXezS3WasVj0cDSOu/s2vsKJxK3DlKV
7Pm7aYIGCv3G/C1WF1gUj3hCun/D82aKwLZ1OtP5x5koAUKOgyB4uUzvr6uT2d11
Zsx7oD3tiylM47+BzHwBOQiz04oaUCmGMuHWVAHHnUS3dDDQn6kRvMhByotabUe3
U0RaZ3vsdpXIDBhHMY8peTOIcdyzLNXD3v4I3eBFbWmu2GCGn/CONC2hUNixoyLw
t6eW5H+wSpETz1EFNfg3gO+Zl8FiCIo5wWik5qPHNZGFFS75Ql0N+ZP2/5qWZdh2
pmtzQR/V70hgL0l/E625n9bd5qEaKaD3MZArdrTZW3prFQ5qlq7ywsFhhLCsAmuL
CcV0ZDBEdcJgHNUcKfHDodQYA9TEnlxe0S4kkgyn+xWySfU7yOd8nHBLRb/ajWH3
iDnvssRB0dOqSg5WzWI+gKikhxPUz9Y1cdIA5b/7Ct2JH1NB70gNMHzxUEaHcPCk
xQ/dhuqgZW2pmQ+bIVZXZLmYPhHsECfGIVjgSOWwF0y86F7VHguA+5P0equ1RxCh
f9JWNPccHeVk9jx34I2aOaSDdmtYrSNqnicsfEl4dU/Ms2AwcWOc5cAR2+oVMcwI
L5f50LzROsr0uYV5GKzpGAkB/BmnBlvEkeDmmIBuM2GvcvATTeHFj+p0+J0HNtTA
G0YLogoZUJc1jEkRA/o3Elvd2Y+ECvOEItY2Eb6VWzThFFFU9Mn1bOu7zRHwPtxQ
A+ZT4WPBGUbHw3z7VPySLWjp1zP/1zaaxQCJeiLLSl/npuRh8josqfuBDExQtMzA
mkQbPXQe+XHsSunYlChct4FK1NmsryLs0Bcsku7nSAwkDz9ZTmfifXEJRORR6SJZ
dZ7i2ONhG7E3GoTYb1PiTtEoLr994ZIU6FnYZlrfjDswY4EJvugL2ESyPQ0UoGF5
t+cu+62wbnSKMUud23KSb7hCQoCd6PpY4u0bIYRpLil8Bi8F4KUPb2NxMIHH18PB
uyhwDgdYNrbk5w4hQtb11T+kL60jeQrIx8mYUgys7xdccMMd5Xkixb5gSAJSxrU7
tkGHdLsGOVCFkTp7g6Gh0jxF5DK+byFQ6n/il/0J8NDJT4c5meWNegONNuJ7w413
vN1mJCLcLnMwIsXpqDxkaOno+PZ9pybFZbGcT+arf3UHufFAzZLwsypbHJY9JUpG
7oy2/qQrvc1QgSQgks/QtCKdGHbbIaUIL+DVX93wtk/zlYklxhxX+tCy0MrMZxj7
/EiJ717fSba4iBeiUcZU/HSm3LXLXRFZtUfTjfteT/R0p2PbkosLpLozsejcZuFu
ZPXAQWK8L8JYtZ1ezByMwpqGd7XFGuSW2IjLKlen629t6/ejjlE6N0YtmIhejwY3
`protect end_protected