`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8672 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aeX9seC9V7j98AHI2NaHVkyQ1n9y8bgh0Zm4AI2U9pG2
VYFuv//lNIjVvWyOfI5LCMXMJJ3JxC5s9hV0cXHsHbHgKagdCPg1rGpDH5MTJKFq
VXSUCMQmvt5rvrcZHzWI4JFY6V+l+w+mynKPUWHbFq6ogT34YGwoaBcrMh5ykSQG
G/ufrWzDzRFYoWvG0cOFg+pIRuimngoxEMzWh2BLKwn8hJ68KbLSstvO+MGE3GmL
0WhyfSMu+H6JPfA8eaexp8IxvCkVRCl4ZIkpwldRA2UDY6l0xyDJmPFep19s6xLr
zov3HhoooP/XqSncMKl1aFTV05Z+YnDRkL+dKzjVFaIkPlezsnktZ93mCIx2Ct68
I/iz56afYUdRq4liPNY3aj7qD61luG4AsN11x7GSrWXUvcrJdBNI4mbCYKs8U5ok
tNS3YE8aQiWybfic2QBQBe1trlsf1/eeS8NGWyDB1F98Xb0j+yIbqUF9RPuW3HUx
Jc0CcHYdxH3JBBwBz1KLlpvd63tnX81UYbRB/0BoYWb3YFEMsnyLbkFBct9p3yrv
+LZCY1/ljc/BXLEMOp+Xvmc4piF74Rh98SguyEgr/rm+KQIGf3HxCIjy5qvyM0Zz
q+nCJ6SsJM+0oVpEerfBKwWWPzWddq0EFBDx1R1AXXmfPhYF55TzBjNJzGmrtmA3
SZh9MlUwI6zwqwRC2q4Tf9jvPAb3pkQy9qmRZCaZB0nJCLYs73vOXa+TBdUklFXu
euq8RH4Lzg+L1ZpPQvdz/8GOaK8HDw34fuuycaKgl99vdaMb2IHghuPhjJi97o5D
mnRwDSXFW8v1Mfv9j++q1VhYFR1xu3P3IuhM/+e3LEfKu4Xttbb+J1EhTM258HDp
9txT2BqhhSfMRKzYRwc6hZ7UnL1bkF+ApQFXsl7S83L8zwvFGT0FdAUwpL3OI6Fy
h4t15eoeSqmTrOj86PwohV1i+bO8VeaYAGaqDMrKu04jDO3a4sQxPvjqHNZiIsVe
mIVwB2uY+ObAoWqOxN8UDbWuB/vws+7tEvqBO4xtETz9DIj0g5XwKv+rxX+ng3q0
nIgW4jl5uCF5Tusz5bWgTevZKQV/3qftfZfAB5QnDXk2mV9d42o9rwYQMBMEzMYa
QNq0gyGBkmB4N5UUc99hX86Gxks8sCCLd9AALGoIEP3nrQIPYHsY6/iXfKLqMnBh
y52JVdGDuEzHsVHwQBRhTaYqqHgMuVLAilBaEp/nyhH+LlpZb6NqAfTVIfIgQvhh
B0KefoOkBiVArwHvVIaA8x/4z/rkGfaG7K1DnpK2VG8vraQvNHR/EGk1EKjzcx4l
q1K69zpjd82QAu7imMw8UFvJtWHyew1E0DVi7dapCTGi0ly/dJkNcAQM6l/K6llF
B/NPK9bPHzxQwc3MMZitePIta6sBNyzqhjCtQqHl7TmuTce8YpwkTEahKv4EamEZ
LvAwaH2supzQ85j95bU2QRmq9LFYC7NefiHZMRH/DL6K3Ty9RmmDsnF9tTc444C5
wi2iXIXbhgztef+z6g+decjTeEtDpZ2oBqYyT/hpNxgCPk4yCVw5J7A1L40PK8tx
Vj2FFZvfic82pi42oggqgVl7nqOuj1fTNSbydFlYVFiL8CboKQTAb9yilCAbH8QW
NqJcDEQy/kRCN/weyCoiYxDXGnnhJPn0y4dmFBDUW+rMTInJ4YcmVMb4vuVWclFP
VUGg8caPtuLN8neE6zVT6OFYsBAKwc/Ar25sKE1gR8xHBLzfx12KrVjKV3KfonZ1
3OLMIr4IQOOMPgRfrCDTtyZF8XwD2fk++zsO6H+KbmrE3GSfl2jDBSZZGCc8Z32w
yks72BzKifJRe1SWB1LLL8Ec9IRzariCu0jXVs/G1odNQh9/DaAOmsw9FOUraey7
v2/0wKylKnZgRozaEDK98g/tEKXDqgCJhdDOyrv4ZxkX5KaqS+0YoddoGSpPi3uP
lt2FS8xpZGgw3zNUK+SZG/0NOIib9P4h/OmiMKuevqXsaEYp0TTy1IWMAJ/OWflz
VW/6FPZ/h3PeXYNSRw8pi7QAdoIYZmNAXKSrP7L/Oh8juHCU3SI+c+IM1/NVZr3+
0bPzSvkd/8jPUDeeREZO28JceiIs5NKjbKUthFhf5eZGTNhDOB7NZlswiYhGMsn/
relIbziZSMmYCzpqIe9tdPAH11aJcC1m4gbHuSc9dVYqouFIcDAvpxLHtx37aUJm
V1yYAHj0qfTBSmCEIWH/j+FjSpxJ8vey6C2+Jgh/Pxnm3/m3AR6HoevcEwqYOZaD
wvP4UpGE6TjPB1T4puMtuAsvGBHbVqQ1SqE5wNKyG5bdZUexBEKtXS74HRwWV+bA
bg2GEN+/qsUQ6QfBmqPvGTIcAa6vepKLUCghy+ns7XS9e8reTEPChsLMt+WGDpb6
Z24Rou+FGyvHmv/8jhsKI4Dq2FXY33nM/4ThGAAbVFwaJC1Qjjt9c6Qbd9tdcPTh
SzNvnrfFAF2xXwC1cTiXkyTUBxseXzGjQIPKUVR+p6ADShWlwKBtfFeA2Fs4wXIn
MR7AiR1T/oFkyy7uWgssHpvV90mCbCoW+5XKprfPkMs2gDukKhwWbU9+wZmiYFl7
T9ySro3DRU6uGQSDl7dzq1Vl5QFyTjvzQ+FyMrRBeCkytq8JsMHUNV+XFXdFNcdm
tTipZ+hjDxId2v3myXVnHvCjvs/sol3ae5qVmwcCKLo35qZnodBbv/lbK0gMNOSR
P6ce5qbqabtmBR/W+VAVYPGbBUzu90+w2YCePnElkDA5J3Y8R67j7jkheLVctnC8
oV8wNwYrCTmmN49RS4jD3A61aAnhzwMSATV5cDE1Huv1mdu8mrzt7hpObo4aP1s1
015rK1MI9PQJh36ScJlcKAC6lN2J1JwcQR8mWjFu9hhlMofaPCpl+ecdIii+rMfA
GskDoe+2vKA3KHx2XRGcraWSw4u3q5wkSlBKjoqja679cCaVQ63zKmoqfZfyhWAu
wfLoKi/hFnXbFMUBdkzGyleRAscp5lxbYSg1DGX4cxobvZCDu4sQ3fVsoi1MOgUN
9/MhyyhBjS0qxBKIkj8HAwv5dbXZAhXSzrnsIcMCM+LYtDcgf3lmMHBFmw/RR5GF
Icd3XeQvkcCX7Q2lQsSpIj5zxGN7BTUJn6XIwtyZnkQLpkutPhNuj3y7NNFkzBYr
cDM7qwm0c7e6bFyDadJ4okWsVPh6m0C6ie1AeyC3CmFLLNsKwAXSFHxc1iCdOi75
YapLIGQP3kUsyLshCG9UfpKKzMGPPSWf/ULeCC2wCFVmFwsA2dHGTbestOIBMu9v
v8NZG2l9hxK0j0+y2P//mcJCNjq7o3xlJapFRac6JYxyYmlbAaKzJJmkiYj0z0Zv
4BleJ8NqUm6tYiI0jym/uR9gdogrp9JSlTq3PNn3ynRx068VUjhGLIsZjj9pCdcR
MdYKdkGH2MpPWFPnFdcYUjx9l/R6al8kddH146fvSe0MYdEhHO2B4eurj3W/JnqS
yTvDXvkq0U3zbA1KhBJTpbrdIabmL0d+7y0RrLY2bG6hCCpn5w67Z0RcUuKWC1FL
9bg8UXKWoAW8pCZS2zsI3kFxf2Y5hkAQx/2/s8LZ/ahCygmTsK+XiAOu6wTgfi+G
pQs3hQQ5GwhxcKOsDwrEsuJ+3kiFxKiIYhZOgORTb0HMgGKNhn/TUKwyHSdZQHd7
GXWdiDjSI9gnMUz0R5VQ/QYaqp903R17mr7NC0vza1fzNOpX7tCtDtflp6h5IvX3
wxqFRBtfOzV98GyTw2q8m1AiofRMDvnwqDIW0GJ7OSdjYpS0JK2bDMjNEKHA8Oiq
IDccaofsPm1grlJwd5q+HW5nwZtXm0opi0kjDpp8tPL4Q6SRvrDGv5IiO0jWYdr7
2C5ecXeD1ZZRZkJ1oZYB9N3Xv/HRPAYL1TQzBcSe/NEfYy6cgc3TnovFCr7qZv6n
z5+E85NF9LQTGPqfzn95hF/jsXQ5UHOHS4RttC0+CeWZVdqfoAjajMC5r2hwR8EX
lK5vmwbm+vFB6IwjF+2JbD4SbuBN/JjiFVhGYPRLjHviX440t7mgrScTZWeUBeKc
fmLOMxEUt5n8RGqfRqBl2n/4zrpF+yI/YZjcYJX91jDh5tw1Y6cKcl/Anzu2t+eN
AGgjd08krflsWciMbzfRkmlUmfak9aZ4RdbPaoGunMcq4rcGa+0659tdegRoPKDG
XUsoSnSj5Wl45as9zSGJViHCILV/fqVUNEUTeXfNQoF3Dk6GLSNHRTZ5MCjZONFX
pXihgIQ7LSfuHPSsG5JxghWcSyTlFI9a9CbYPFw73C/pOXcR/uo/6+N52ZyZ6bs6
s4YLuqlFi2PbJo1RC61RqcdnBjk8mreU53GFqP6FuDdLWSvE1H+lJJgov+DDxElO
HRSG7EEHGVuPkRatnI46Z8aL3bJ9M/b+uX1jWka1NZXkmlxbTRVlBVuOyq3Bcfri
bcI4RXrG7V5L0fJvm2JUtHLYSmfEOMBSMuyu0KN4pcnOwb+Kip57lic28SsmYUv/
4epqxMlKf1hmMBmyiO/U5w/xKEpLZDj28lImQC4mi5R3wD7rboeL3pqYGPUkEXn6
T0bmcWpz0kaxNNXWFXeeYJEEC+d6rC2fhhvv8RbXNX0YFnjBtKLM4RnD3zQwWePp
Ls+mfoSX8AGVMBma4kEqRwfBmZXq60s4BDP2o3QkihJZxTbtYjSKZrTEf5vlPo7c
t0TEIl2UAoMgMy06ql2BJ0Rt1E1IgwWdW1eoJ6i+W47ALFRRrOCAuWqvZvZjNaS3
F4E0+dmOHaFz8KJZ+5keoPzqvt5+dzlJ49JJ86xmfX8evWzemE13jy3uIlueXcHY
ZKFjDlj9xG2zFKesDLk7Pm1F1u52nrBFb3Pe42XUxbEP+nUXpK0GYOBLjIvmFOAY
LSNbQAfiZ/Bm982OkUXkRYpxF+S/+o89ab0PqnlgOtg2NipQU4ocfhsjf1tl0OxH
Toe2LfdqocVW7wGuAx1C62y9ZbvDIxGAMoy0sNF5jcwhiSHt2KsuWAKyFtuAUkGb
drntBfV7QadMV3exLXO9fiRbR14dZgWj/0c0KkfiUtqvdLGjHAk4tACszMsKDKhE
JEcYOrKOHzIdeLJGxGyUvo8KbN3Ryeg1WtpeNIVLgnxQTqnUJM1FwlFlFaAh9PPo
et7/IB45atvCVH8z+HnNEmk9atF42GUfuzAxKjp812f1ZARUe3SBGRv/DEm+CPQO
j2IF2T/OcagWAwbrLv7OFOQXcE6eYrmAcOr3MRKSlm4d308L+mgExY5HlzU0mOfO
Mfj0dtrU7aXP8enPvXTFtZf3eTBHaWnhBYZy71rtVlMN+7fWc6BzpkFzUARTdrck
Nm7q78S8wxQk7cMmCuSqqT2VAqT1E3c75GyKnrVDVZk9iWBfmY7FFcCiLGVAeJdC
sems6ZG1IsLRwJegFNkIzKXXltJyJ3ar8W33qJLIwL//bBhP1bO0MwmUhHeLhiDv
Y85M+l+609qRdxjfKz+3nd0Qs+NW9XXW2IKP7txSivrp52Lk4pBJFYucuwCf1MOL
g7mi5P+wxKaiPLOK1P6qJ01tPogzuQebow8D9UIzo+5JySfE5/xZnspHQ795hJPR
IePEC0HW7MY4UBWfHibiq9NliEiOI2Mxw8kPAX0GZLinALy8IyqFNxC6W2AB1Vtp
caYOyKX4NqdaLEA26k+2Ed4t360R9cBIpYKNjq4nR4OdwpULh6+DKv08eY6XoNIV
o/Ve6qnzuvrSI/sbM1kXkq1l7se6pr1k65NS9sfCH6Q1+vsJDM/Tz/LCfuYQ/zmF
PUXRJwRvB83uGU+cEGH01ZGxJ3f/9vtWL3kRMVweyzbTfMsEhklUINg9YXHYaK/P
qzCNsAd8IBhJB+JhlFXTJI+hjmzxdCJKFqZTbWN2501rsWYuaadkmyuRTAHbNbnh
91NdaFeIfq31h9foD3yR3DMb7GsCdITGSkEXYgmj+2OsmzsxESqCghztyV5HVQZD
Z6ZoiwDlqLwtfiAkP4DoqhoL55BtHh/eBppFi03PgksSRLvRexEi7mxP8kN4yt3g
Ha+iyGhr5qdU3h/br8LGZyGWC3wJgCE6BcwZoqWP2yKWwyOw18DfIjewCA+YVcjv
EMdMeT8pvTnJUxbg7jsVI4IOSdAZU2znEkC0v54RExezN4d+1krK4E8takaed1Oa
kkgB3QDskjC3lN2O7ZNDINmfk2nx7Qq2PfS9w9QUMvbccXc0QqwaZGZPgTP5DzXF
6OrUe4IaxlmjuXTwlyy8Fx53HRAwd2JjC44s55qYakrTkRO8Riq1VnuBaVbalZ5N
IqjLsaDQP68oscE54O0OKfaHw3+Cy6ZuTuZmOXUJ5N7YynDZqA2UQeZLDJmqAR1r
9j1lXhDCGLbpS1v4tr74Qh2jmg4dHet1q/Nl+cecbHmSnJvB75Scz4es4juE9HX9
6yA7f8ri5RYX6R+um/XCQeUkK9D+i9nrhX0kkV0+d+DYoedAPk2XOAuZ5j51098/
JelBXz2DzsXkLm/KH2GZNj3zUzg90edFZqelI7WNic6RRDaeoRvaKY5Bt+3IVEqD
9TmmoEJzk9ZiCvjxiZ+iY/+OlylQXnrzyDQW4zqlCpl/5zJgJk8ovfnQmzibzbj9
W5yRVSDT6SV2Z0LkmYob6YQ9yOPtGTafag20HjllCk9rliTLxDStz7rF0tzmoRcz
VMuNp6ixC2VPEj+gGbeNaOQXQCnxRrbRuns6jMtTIf766mmonhqI7B2DUl/3RDGA
jPDHJmcFevLn24dnf/T39xE2O8vw4GO3KwV+9ej6zI15ZYLSlgbhTDFmzz2H2m72
b0Z7ys0mRp6kIpf+S9WoQPvOCWd7MET1ixOaFiLCt9bPgHdqyfLpUIfWYBRPji96
Nv3d1YBIdi7eYPdQDb2QUtAESbpxZ6xbS/4H7ttWZU/agzUWDC2FBJSfNml9+llM
xPv3PsKaYbGEKLAg6+exem/sXGoAPfx5e+yatD/bkh9eQKc+OboCKBAcbBE7Euhr
KXcFbAfYSehMJ2/sd1J/2H5hvIzlrwN4ZK8//ndyKc4oeA3YJJrqiMfbSbyOJLP2
JwrwoJNozU9JbF3zwED5AToMZH4ESqnGF4/4G+zp/Ay9HWNoXBl+SA5/aSfE4VWz
p/91Ic/k0UogzsX6JawJI772PhZYmkg9pz3JKtHVMTgTC8s8H6UUeryfrq6q9AJp
UIRv027HbWEfc4sWqzrygwA3/345TXHmSpuDXzs4KNrdlmjNoOcQPI3W10zqNPJG
DryMbakw6IHGNWgcPDxwLd/4awn6SAWMmbb/zEFkP4wcTH7S7dOY8dAVOtdsenXt
BwAFeZhZcfj52xNsYAINBv98bnkjkd1baCnZ6F6rPGTET0hKEdWpdvvJojOFrsHs
2Q5uaX0FxK6J+0dVmcg7tNGDq1sQoRFNqB90Jcb7t5gy0cExGJYw8wv/rq2ywGEU
0iUnhtVs/8mliBJyYfBg9DEvUQk1MfHbX4gGEyNpqxIK3mLI8EehT8ABd9/U5BkB
8AiBP5Jgo7o3sWN4iys8Mmb+xcaD1tpuQNC9hd0sIiDQwZIYGmApsDME1hmBAjFQ
JvTjSkRGiUpES7Hcq+4T1UuvxOTrSubAHWf0v/WiICzMJ3ExrHcyR731JbdH1Dhu
4dZOIDXSkUFvoJc5gjNG0no7+HdBcBmerGK6MEzhCEW3g+i6mt5aYC1wntQfLmMS
25PYcwKZOBOyzv+HzlbFlYitVz8BShBYKlMWNWNXbYYvEWImhe4HWoU2kqhOk15r
N3mXbLUUkg6nHGzP5tb0iNw/reHiTtW70u80iHRO3jwq/ruT9nj0CuOuWljxzn/u
vnPiKNlqn49+ZdgNJ0H+Kt5qFMmcBmt542mIN3ar+uEd/9GmHM5C9IY24vWJ0Isl
Gia59Nf0cJ95ycwRUvw6NPXN4KQY5dEb/9r2YVi2TwFJpC4kcUf3QbuIS+uz3QlV
M3rkpLQMhY6L+jYNv2sMhWsBwQiKfmhz4D1CbaBltJ1tBBA2FNW4QnPk/8881+Gj
a8Li8HASWuPlK6V6lAl75k/EQXrrDQ/x5Hhvk7De2rmUhv7OzRK/H5YAvsqMvmc6
Elrc3tFeluBthwmudy1kIwyFcGvXX6XLznXOZZUPre4gZNAVzcgAM9cyesBaUaeW
nwoMe7/hsIGm0I9PcTJr0pJNfyF9sGN+7YGOCGGhuRGzXSEHpZ0bInTNtGYTgqmc
YNwe9RxnKVer4BvWBge5ZE3Nr5GrdiH3yAvuPXMGSKmXAWP3O3pEuk7RIapjVKkq
S9DWwIqMfqdKPxX8dSEBtwkYihI8q6Xhit2kRZ91zM1ohSwYf8z/GGs7Qt4D1pRK
eyfZcHBozb9G2/FaNERhVSOeBtR/tiL0cCow2vFiDu3CMkyKIO2laLJJ9n3/oupl
3Omr19HUVERaoXnkFYmap/MAy6o0WKGRCbGAf+QkN6WNTNtE+8MfZZpWIRD7vt+A
wWrbbLGR/lzVb6PpIoN/uizDHQAyXt5VavWtpcT33T3BeNpOd/e3iHYz1CjEOJ8N
RliNAW24CnQlA9f2VJ7/pJSZ+l9uHbvKEhyDfwQchXj5mGUBrQoSUNo82CZTYfui
oI1ovh3mebzWI7VeRpqLHZ3dEyLy2BEfcICMNVFkL2CLJmqD/kEEpi/yC4ltXmX9
8UoLzcOm8X5p+Oxf0fJTopJEx5/saGdxL0522bL8W2BtkDiWLi9i8e1a4FSLbZsY
fK8lvrMdlYTI0g2sCuLfKwDl3dLG13lu120hXSsUEK5fNLfwLg327OJ6cmxDyUkB
4kSVKK49j8Uq9OKXzwWrXsPK3JxVjv2/qikxSdULQ36iRjaYfv4pw1tz7qc2PupR
iwDCJnDLSXAIhnWdPl3ulLB3phx72sR9okqK0ElVhZ+X8yfCkHY/EJRF7IzdDLa4
EYUzZG71vOxh3xxQzwvPf27LbSobB4Se1egfZonDhucaoq3372Lx1wbH3shrpTEr
gHzuOgGfMtIzUu5xDFL8wzDoXZStbsbGCalTYysxtzwLCZPaTAYAfH2RUlX4PVMr
z1d6X7DtK2oboS6kewkk9zMYVhkLHa63n2OZogNRN10qiUTbeMmIYi/VfJERc9wY
6A5jI3/fK3FaP3w+bRqA8FowMsH7bvGhCOt5LrMN1AWzij2tx292VA/fv5yS/mDb
pFGtI38RHw4x3LC5iLVfQJtj1mrFtdqcarAo6GW5cZmLucb+nqAGU4nVdOFmYu3/
ECdFx3NpeGk1Xf9AccQVte0so4LNniaTKns7Wy1zBNRrxgBqa9tE+Yv8eFrE5Kzs
NtUmXLQKplI1248hbkDZK3MMNRPqpd8z+XAj3xzNY6hdg7wkulB0SpUkRkomVrcA
p/Fp791PdP/3MXM5xXA7puwmCD9/MxEwFK902yCQrqeBkp9PK8EIwhroWy30ko9z
apO1TY5Sgx006uULbqYyIxe2bfGHcVdNScQaRIXgq/Uq9hYhm7o7JFcBEkXgd5Bw
VNhVsZioN92U0QrZL+tr4aGY8wijTMMH4qWLTj+98NZQQj+nsCZfmcq/F0mUZqp0
proIpkY/oITFi4ofjUf8MJN6SuyH/6L04GaOZsflwRWpxNI6llK6tufDIXpvQb26
FAIIWwFi8RFIHcttZV1TH4sRsreMAvfcM85G+O5K84It3omqEUbzYr/KI9u+fBnN
IytYfn9wmXoBZE1m0lT8OOQ141IbpraSJZLp2E48AmITvh2hWRNJdt0em0zCSmvi
cJ+YSW4YPF5F9sQSwmA90NiL47jfFIIzA9f9fuVit7Os3idEc0m/SXGspWIoIGKM
BVgtu/yrDqa7zXUFTxLOCu3qiVpLX5HHuCX1/T1d39vlrYZWKyLic+QpYBdskqhM
s5hatL5bsrQ5w2paY7VcqesHHZwKoZE/mpRNSHyeB4KyUxwby4Z4kv8aFg/JzCLo
dJQvjqVvKchbgCLS4oL9DXKSXcgtj7qx7ltBqCF2+uLeZv+6mTTf9xU8msEse0nk
Ke/aH609IBwiZxJLPjYJYx9OgahVBHY0w8DCGE32ENx96+me4SHbconpUUSPgTKK
FqMhc7blgaN40n+3NkQ9Q6/HRhEUSS1j4zPm+EgpSKaCVew6JZpc/FYDf919mz6C
EgEQKOMGK5VAvpV1DqFj7CU+4z3JM/dtPbm1ib0hiCWin5Jfjnt4xj4UPLJ9YdcC
LYlVMRYUJDXOxMUxYe1JlOc5FTw5TVSBSFza/FuB8Juowg/kAC5RcIKeRDowF5d0
D+qA2W8nds6E8QMfU6/JxZ6pOeS4dtfN0Qti6iMF0KBuypzFsjg208RhUIZKbFAE
Gc1Mz0BgkFSQIm6+GLPq+XLoQ6CMMJ/IXwZqaPb+d3nGrrN7bi0ajYNgG1xfg+tL
649SpxexMerYjE3DZzDmqtIGZ306kUqvxnHEcPzTs2RN+x/zOiBEflFwNMCIQie4
Qslzm/0VwK6NNXJkA4vYoIqyaGnINVLRORwQgruNB3f7yU+46QNJicH+YrfD2mhm
jLMbxNBiqjyGaWRoKdECRWnfwKzVSeRqf8bCoCjmtPSIzH5aE/Kchd6VSyy1xzO0
CulvIMPkK0zHrs/6USluJvTSqP6vptHteuQ4MsA9IbG8y3Rv/EGGnkAhVFXX/+dI
HQc+K7ZMUjZUmpp1fO11CQtS9ZknarEvo0avbGJOf63eTAU1OwDKGEDsfuZ+BSTr
A5N8WDZmIEQmmUptqmGL1Dh4+23ae6ZhjohqfKQuP2oIXuuH0qRHRVmyCCDU61E9
FQJaLpZ8ItvnuejoFdighATYs/5FmCN1GmFgHzYG/qAAhqrp8c3AlHwnxE2KYTql
FW5GV5+fP6qoJT/QnU3wXgsRlgp+ml9HPf3Xb9z6/tjzhot/aAjLtHbKs9cv8TQC
KNIBnYgGeojQrnxV2B5mybCgXi/p7rvYT2YN+Mcc6Q06MpQvRMBzKpWZL46iDNJh
QNPD7v5dvi1EKc8XdS263Mp6/xlDfkFNVMECC+N+ZV+06+guMRc5Co26uUYykY/8
HTpoa23hhMI/ZZwp8Lz/dghufeuSo3I2++bFuxXwYSZXOoAJdLQQKzBtMmp0Wsb2
Bx5298rZ091FIzj2KrRWKtABq6KuOILhHpY0lPNEk9TEV9NvqQqFdK0z7LiggTHx
bfhf8TQEdjig8wX4wEd6FBXjJiuml3e2SuWMGpXqBg/Bs+AFGR4a590sr+o3BKiq
/uE/8PR7Se5eXPKwgL0GKtgBTpxp5ZLW9MURw15pYTba4+lGKSIaJaVFboNLETVj
NqNgdbS9pvhRnv1IdEiXpIs32hghnC/IP8IMNswZ/D/yf+RrP+mRpdu4vUCNw0zq
jYHVLExLCeHvylJS62IimdrgOvsA45Q+gCu72JnI5Gc=
`protect end_protected