`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 33072 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
Oc4fq76CzL4QYVrEyjSlCFKNcw6lLYIiXu7QrzAoowSp6CQJouNkj/O/OsYpEfft
INZAzpCqRzrhTJk0TwMsYVKg/EW9nIZ0qB/MAtugbiuii4mhuFTmNgovC6QQWPvT
v12Y30w61ULISCxLWmqsRnC/K2VgEA3+vH6kpgdsqToMnC4XAFFQmkeDra52KNbS
1FJjrU5gQposqv1YldtTQDW9/FgU03iwHmPxJmCVfD0ZJIvGHXl9lGDSy86FfJ7x
apy0l00Bw38I+B3T1ZpmT6SBh2uK5x930dNg3LtXNvcUF0Ekhd4ZrYqcN+8v4o24
2h/vSKbcLVSu6DilX20o+yzFEzAlPMpk1/8SbiwXwLVU8eTRoRWrmFNqFC0PA13b
TlURZA66YQ1yC5DL3CNftADXsaLNURh27P5GG9qID2pBtCTuDIJiy4SalHYfLZWF
U3Ac6oz+RYaq9U7P3YCWJlTfOrqM4O4ivxVQbtQYsqW21MvIPNdrMTRJE2ixDdhW
XGH9Mmo8CFEdEJUf4fst+zXZzsyDNcvCZ/Zm/4B5E+OFEfpS6x5tzbp7sAkkjNFn
gER7Gwucec8u6zA7K/ItpX/UDvdJfFtYQhdiPGQoItKWY5sb0U4YQcEpCpTUCpbq
xbo3bzbvmJKoMOwz+JOufTi+rG24EhzY1yFBRlazO3Dr/IahudIMMT4h5ceDH7nl
Wi8eelzIG2z8AH7etO5Iszr7fDgGAecQruqHd6Jbe7rE8wv+IaIy/je1wvQpJDEh
DAGSTlU7t6B2F/LjeF1E1NWud3Ivg8qaXQu3/mjshQLOcm1GhaysoknESeUUwUJE
bjGFABhNita3V2mG2s6Nm3r+Hm0y8gkMk0qbCj9hEP/YQ63umJVxdlIHXZV+ONK5
00IRCufy/E12EVcjZWdnLPMXH9O9EmzIj8EOUSXmbF1F6bwZSGdM339wBLI1T/d7
O4Ut123TqtoAJnPmjfype3SptPQUlTsVeN8WyF/b5QzAcRYfi3iejgGr1NRImeY/
/1xx81NSb6k805idC5UL7I3SkonNlbCRV7/fZYEQ8uh/SxDxGnncZakf+6AbGh2Q
mzWqgxm0ymjRpqCHXnWUXtoT6S6ucakbJRNL2U0t6x7JB/Qdc1D+HS6pOm5c0Czc
xJM4iLfrizQfbbLNLR1SNYwGgpOz91DwAJt/rwnFSWr6zM5SbNd/S8saQyxLjOIf
f6S0EMxORtoVBAtC4MLSfRxt/aSr1/k5XbmYIT5zynGLohvGp3L7AGGIFtTAcLCQ
lUjVbfTytB2xbSNjs2Mqolipr0pMYZZtLRbfB1pj5TIBLGG93p0NeNwfZBNXpxKh
O2qYwknOHIODSyjAbigK50BuYveCnht20FzPdgF+TD55MYHQbjv+GLLAB1Y7jJO5
/+pL7zAxsZMyCNKQ3ok6wu9OowxgVPwZOjx1vmp6qBZF2kI7lcl7v0wgNLGwP948
K2wGKi+HH60hDwLcg32HHqMpuCy+EongQDdrqX+tpJaS1MgZTEpk4nHcmf678Ihy
fbddVgJc78AjIArfI+KakaflkIyhhqlepmqir2r+wHEUHWFISkxJjMl1PUAGTNf9
7vwUzSJOK1xuMxfzsfHqxhlTNYhekyUQzGipYV+J4K9M7+6VPDiXFZczRyS233kt
BB1YxVZyzl/rLiPnckAj7EPASJiKz2kLpshC74LLrrf17/BcHGSGXmMlsFsdv0Do
Dy8dyLXESby8Bq3w/3hl69VOB3cHuaOH2FY/VRP8DN/15zmHrTloFkZwfEDjbFRN
cSk2ysL8utsGeTRtr8TWBgSI3oiUT90sn+veaJvL39vYueUi953Kv606rdvOK222
MXeRIwk2PINve+lb2+/8DFLHuVtpzyomC8lVSUiYYTQHFwIz8GVS4SRgMhuZPX7H
ETWVjzqrVXjiubfTV3y5WWTlvkTZkICYff6nFeznkkTCJ6zp0q1ioGnVFvu6Lwcs
WeIFoecknG/Q0QherbGEpiSpEzITCaj8mzAtETd1C6NHX3g9dsdWmNytgf82vHs3
6mjQLgLHrR256NcxIeg1+UVlr6CooKv+UmlcYbo3Y9M1PCH51RswzkEJkFn5o0oN
3XmeJMpk6GpErdnMc7By0lD0ZCZDVpoy+DjavPAXPOgDeMIRgWNIms6NovRBWNh9
mHnKC7f1vuFbgROcNAzowYseUKrtUaZkgaBZFPLQOwMAmHxN0y6NvzxybyukNMUc
bwRqbRUCT7wuAcebwcp5rjiE2vkOR5k+71pu9AILTy7C8ZH+B9Xx7SHdi2QDsjBE
QU8oCHXtY+nLf6CX9+n6eXF6CFAfX8QCQ6Igcyxm4M2Gsv9XJnwpNzc/CRL0zyro
Rjo9hLRmgeMyzhQ77BbX8aMbcYEDKTdL6bP0b/TX+LeRxd/uc7u8oU5rWtOBby8E
qbJkFnV7/z9Hh9Bf9gtwH1X6a4ibpLgw1/9UrKteBoYrOHpXFyg656GaGRkKrZIe
MbaxVtSaza0Y4uue105E3MTLnD5PwesXUY9/HYB86Yw/mPG6rtlD4vtIMd0kkGJh
hrYcfgkLLho1g5TSECllmA82XS5yKqGciKoHN0h0cwBS3QRzKennWMdF88uTbYcD
RqHego5icksZma7i2yVc8GS+kq15OSWRwm+bvz6xzso7QyILNlKsEj4Ad4ebG5Nn
QaumhsAM0Co50MfG8vabgrbG4m6HgnuL+pP/5AUC57FqUsgCMO5XuAEQUM64BvBo
Z8Lwq4fFlcl07NTRtvEkDLHIXR7aqmAkZUOiD49LqPsiBUeC6U9CAOc5PaqcEHz5
k+OMBAWEefs8/YIUMbabT7/SypxKfbR6JwbPlxSUs8zX2uuQDhh1e+GtigDO5Nhv
BkK8KFmzIrBlkisOIjopd46YFt5X8z/+RmjqBSA37YhmMTfk/7V0hJk8mwpvrrQ4
IWDzsFpr//GBSVzKAdbkdvBVJq1zxm9pjalBLFBZSCY5urO4y+olH2n2b7gf1DgX
jBgxx4mHMb+Fn42xn+rodXrmKzmtuI7KnA6XOnlLVUNOfqq5yZ0ctq4Rym/QuNWT
NBaG0D7S6ouXfmRFZ1xWGsBKvilzC+/mblpIfh7ZBd5RFrBawfTt8+JwGuACryJP
UipoALPKvt16afPbr18z91MJ3JxDxWBCnPbsOrWpO1yVBdxddae5cEggBED0wjy8
uh7kqO0LcnUfb+PICDgmRWy40bFdge1GeHpmMPgrvxdyaCgDfFagQpOG7fR9YBnC
Su+WpBMjfWj7xm+jV3Xcx3QkWqJGqJ1rmo691PXGYiZCZDobhOHPhZ1iqH0XA2TU
bpGGF1s5RtipDpmKynvdFvwaVT9QZMn8OyUsgO+DUZ8gp3Th9o3E8nzCvnvOPXmz
CzhMs3bEhK6zR5zfR0v1NggDuC9+D+PmWBktA2sWSJI/VKUATLbfNQG3qLS2jNXs
Cho1XZLtXkqP0g+OGmI2fswREdtQU/8vY5Sq9zXjOdYc3O70GxOWDh5geBcclhlG
/wYX9oTvUexrbrBDPjDTKq8XLDr7wFIMAddvrW1y4YgwRqAK8VsB98jwzDiYmPWt
KcddV7JIyS5mEQlI+V2gOSFYirq6FVawvOS4HFHq+F9vdqlBLUoejYWslmNjsT+0
cGn6Zw7jyO2AH4Uyk7EoiXXqoLMcT5A59OGreSeYsnd/WsOQpQiUnUAKfLBv0L76
m2nNAZoGeIEZdg9Eefnlgni6ya/BfFnBlnXELDLSuTq1A9/L49a2NPGtPkFr/Pea
UjCssu7+9GbLN6kSAGl5ct9LeWARV7/n/0AlkB1CUetJKHkM2Hml7nZXtx51hIyh
rGnaCNbcjndOMBcO8F1s/xyiF6LmyVat0ME5jxJYt4wXnLD3I5ZmOM5ytedISwbk
7/10p1DV0he+pindeD0hJqMpzZ4wxXyyejyr2X3L7g0xoecAIR532f7Owcm3fXx1
3LWwwztKwgJjgf/fiP42qO78Mm7X5AWQFUvpJPGdIOrLneZsm6btu3H9uHVdC+b7
ZHjAWGP5Kprli/rW9TcJjFJNk2/51qBs0mhxRhi6YjjghwaTGiO16qdk4TdaP2MG
Ec/h2ntuHBn/nbCuQQKhTBHZ84+1IvyyPM8YGSPuZXEY29x8pIzSiAg9NXJFibcZ
nCrQEuoHuN5LgG0UdLXQ3he2337M2PI4yUzMpNIwpaDlhqDgVy2ie0QceqFiVweg
W9gCS6mNJzZPCMFseRkztWPShB0ZHllEWgmgortkVP80E2wGGkUdNjXzvQ6qRsrH
cJC8jFrUuRDSLrXU+FzjciUhrJkg03+yqOacSEBaxusS6BTNErRKCAwp/ZL6sBSJ
VmRmqddyb8ozC33WjRvMq8uzkYjk1S5iTJwAMGt4+Zbq3wQXHjKy5bVlt7jvlWq+
Sucypm9qSV9hTGQf3dgiQNloLd8XlH/pxwWSYgx9+Sat/3W6JVzX8WE6IdLB5luq
wSNBoqjrxDKO9qoXP4LWjpmcXltHyw86w3Og4Y99SlzP9sHnak2tKOwGvSFdwd4g
22MOB6J7k3UkqFkcQJYqkLwsM0Dmfqg2hDgfo0QNyvZhaxb2QVa7Qo7nXuxq5rWl
RIrs6tYoc6pldtt63eixt8jQve0i/yoYA5S/IfOmPmorxNaUkQ9hZZgptZaI2hMb
Z9vsB8wfqUHPuUxLeR5RndCrqZkH5xiIoDGoQ2+YxRMHVOJb1SR9CKD8WMUtdIms
26oukAlUAJetzJN2fEzlG3Un70VPmb81dUJufueJXE4eG+g4J4Da8Au0fKW2fa4R
CdfUdJBYNEhlzigA5cGyGNEj91MFP8S9YbP+S6uGlU96Ayi7T1ClCR+R3ewX0ADM
B969MraD2sRgnJGQ/otIFhTwHzdPe62GM5QcdsCfZniZp1zjnL2FsyrRRof+khd9
0BeKXETERFkY4b6nhga3svjGfBoOysUXRJRjj1oSTk2XwHHtBVdX0bvBVplEXgyH
imGEsUPJ5iKQrB5MOksiYtC3tV/7a0Qnb7uFuxYjwYTnIFgfck5WWNBhfOl6HWd9
yzqV9QLnF6eWDUZ2AWncqHDefagqbBihwIAeKLqahULj93pb2UG+O22Fz9XidMAd
phneTQ80cOodHFB6cyZspgppcmNiB4dARDccyxcX8Gb1TrHChvgG3uD3DY/kX0X/
6H7nthSqL1/Qtbm8HijdHUewtAt7OySq6PkZEclRBk50PXIWqwL3WdDnbZ03AS4R
MyNzjc+nkyhyP/T56lYVDTJ+Mh8eEmlECGP5HtqeeNM5w/tMFzyjVku6TRT8n2hr
W+EoIVtULfdRd+xYwUzqPa1Juycu3QmHhbM4ORZat8ptc/kGglNhu436qbZNMjKl
aQnCW301wUcrkynAOOjF4RWTJKL9XhZnzU7DyYTu66xLJwdxV5KuISS9sKllYVcJ
UNiKiKmbiTtNp5OVqjaTe1RYz/iOqn9ETsufgD+oCeCBYS/EE08MWWiaMBGomDy/
SbfUCJXrCqPoamJ6zlMMK9rB0cIv8r5RcKa6l8aDbMBUr6mNOO7evdr0xB8z9765
xp5m08EC0xkXJVcfGIxFUQNsld1qAR+m1pp1n30wpP+sMfnQMhcTa66bqVwARo8a
4JxbNrjDlvtqBMArY3LEgN7tEf8lDhWQ7XeGDnJ4/pI6FY9w0tSMp3n+J6/GyMTW
xNwJgmqTGSLL1dlX91Ifjc3cILckRgBuPckwGkJTJldUNqLD+sN9w58Taskl8gFa
c21KnsPLGB3pGPt54N5a7drXAPwR1NyqqG/AJSLXiYyH/jtdvZop/DziQoeGldMo
/dccdM8KqU4Q+U0Kop6JjroCkwToAdFfCifbVs/BR5zrD0RlKeNzRDmytczK5Uf+
vN3c9ZmfEJysSU5DcGoMoqW7nEUOA0sZh0tyFcJ5OXQBs0bIiYO/apK5IlgyzfFf
qyydVhg/ELdcMtxwPbxLbmpJSrJVttZWTDFq3cmxpCAx7vgN/ZPG5FP6mdgI321w
DfKCNLNUYgXFHkVO5yJxOQkwLVFttkGWnFmaMjgFhSVcwN5FCQvbljaoHvjutKhP
MU/rI8hgviFInBErr9kP1YkexM2Bmd+apAz+q2y01+xmei0WmJEPMQiHwBRtsx9q
G72v86nAwtFWeDQ/Iwz03wIrbquTG65vP2tWEhNakC3M+JxyJPxWGyyUL/is0LEp
pWTwUmPWWjSRhXMAgkz9mGxba64yRIfWGTS44juHcHqRwSIjZm2QPrk08i9KGHoB
4hU7QruImpJ75UWm5NLk0CRU9IfDJHb/7QhIaLHfwkN+OYtPwb9z9L+ocJ+8o/SJ
AjBKhcYoCYd6qZRJoqc/jvWSUQgODRm0Dy/0yXi7lFHw2drNlOqDqdW8Zz9gu2FU
0hPDpNUmDi3Cbb3VZcNT4suhdoPT1VQ3Oga/591bnR8fIMglNTVzt6KBUlLxfU+4
vdmiKyPBKK8Hy5FhW9Ppk8wN6Tw7a9MjwvPPc4u7aeCQ+PCLvhfer/qJZkA3TTks
wwK8zxMdWYNiYsybSnl7h9aJyIYn9lmuRdmJkHHiBQlzraU8K782HHwOEDAK4Iks
IotDN9yWMFgQUti9oHDc6QzsXqXUMw6S7rQsf+O6xi6QuWCmYGWadhpszMjBa96s
ZYv/SxbpIZPG7oKvisEz59dRdKrsdUvXNTWncJvj347kPdBoURiA1XZhVBP09REA
Labbm9mOVYVAFhJrq5W0ATVCqB1FxrclYZFP97ddOZ/CuAZ8OE/sEPBjWtOma+FO
N3Fk55q+wotTKxUrMlRc+EAUxTWzuX9L8ukVlm7zekkLXsO8Qe9HFZN9CQCXM4P3
Fmke4lDJczvA9rX3i0eBsV7O6U61FW7Usn5w1pBsdrmuCfjzM8n7a4Ya/2HmkSmC
f+iKPrXcqr8HiiAxr8ivdk+WAbgadYPhqgrWLjW+4z8/bEHtIrNwsnTXNzUXWa/b
4id0MnRZrmv54bMn65q7U3B/n0Y+fjEo1vf0tLIqOynv7bMGgPAQAQHYtuhJ4bQ0
7l3RLc7gPWNeqIyu3YhqwOVDZ9AdjVaTkhATW1Vi+Es6qOGF0n+6Yd1sdRuC5+Dn
jdO9764/abZXV6XLUlDGqNQBevXufA5723uFmY9lslWM3GtP7GoLiUCrCBqSookN
oo9WgPqDpvC05d2U0CNnMi3JLMtzx9TOVJyqAOeZD+UZlvG1fhA6fLOYhFXnlYG+
zpkErXFvrQtYDXygAV8dhqAIMthi3bShJVi1v/s1E6M1FZMpDnscPYKe5PN4nSBq
gMrBEZWwj2ITEDjL9AbsmczMOIQlu3pJgl/DLDLeFXwR+W0l3He1DUUNcuIYzRd0
ZXYdZDsq7PpcPvjkTVLCK7XR5XrU0o3iYZ1kcL97rfTc4/FnzAV6U8XbIQE3y0/B
AvM/XgpERMJlXvBNkOq0FPIGuQNgsYdJ+/REHVMnGdfxHEuygKg8fgapLTftcvHR
F8pN1Ms2ad95F84XgnqNsUcjcf9APlZ54dTbSuYg7O+qHQd0s8YyXo/esVlaSxYD
0A7wSq39N2/W4cDgN8lQCs8bSRh9oYCXZdRa2RNzWLyJRoFwZZuzvCByUClv6Mm6
tiEAbX8vK2IK5NazlfedQfgDX5o1+ong4GSRvBV/Fe3nSPqu6RFT7KshgSVNk5UA
o7/k6MnY7c45R+NLQmYBJBQZN0ZxUJmUHvoJbrGcfrtgCNQXtqKoXg9LIIWC/oRu
sr2rgtTvAK4lpMGZMNMWnmhpHC8z6tPqCZ3I7S4jnxbsG07QlwHxYEdndHfSfIH5
Fxa2EUnTppV4GqE3gX0T7h4VHizmsGAtDDV3+MY6knV++MeRHEU3x4SlteR1BsmN
koMpmtC+LphirX55IWwhBRnCvUfN+VS7V6/jE6F6+18E+jYUtIfVzvRKJRvTsYI1
YF7NFuxeR5IRzYtsA8vzgQ+8H+y6D1sc4e1OOWkU+hiHxmt5mi3uNFWmrWSx31/r
HfZOCo8wXoVzt4o1Nsf5IKLrd/BRFECGk/Kl6vM7mh1/56mHDjgsNObDAR6XiqzW
1KH2w2FErrb2wJJ/Bq4g/X5TQ4JXjLIZ3U//77CnrlVlrS4woGb5LQGInX/VrO2P
V/3XSfuC4VKw7cMM58hBRjC8YuuU0xWASPimb61mFQMsAX2fXrhu98VDvVq4xFZj
aiJvkn8gWiLMXP0q9quz1Q1rxPgs8uJs6M1CkJn70tXszM5OuMfd7sG2VwhBchd6
zpnTmsqWVYij3+7dYpcoqtNXixc5MCFevmSWzNE3usJEM0G/8vA0iATRm/Y18kQw
B/xZEdNKwfyHzrp5sQCJMOIhRDHZ3JTfoMKEhLB4Zpd5zWO4dUd7c0+l5SqhVW7D
6mqwO/AX2LelPalLCruv2r1axF10SaQBC6P1mCMJOhZOccbSr70SwX7hVbO5scqq
e+9Ktr8uttZNAroqKndKsnGrHshlf+hnxKcJyNzxHMPYqixCo3IWMwFHrHUkIbRS
KZkF/d4fka8thC7SESKl1nhdfrUiRZbaDl+1LcvacKSrFWljT71fg/pp9ExY/WAc
5KB8KBRYs5HKAy6EU59zvhEnH+PKQurOXphVjUcVFPoEoNjDDWJAbuuHj9vwD5J6
r7vPh58zfQZ+gUhkCLlZcKjPAV5FtgnSqiJgsQxQDnUgGrOt4QPmUKXGagZzz3i+
roUU+fmapohMC/Jkuzu8X5h4T8bOb3P5LefaLaBVib5nOjpMxcticHLExyXBxXBG
B1c8VO81kQ5PQSLVMwXyDSbPbbcSjDdk3bKCFvKFlUyMMrZw0owT5TMgj5Sx60l4
UyP0PkGkk94IhW7Qx4acqTjoHxEIG6WsQdUoNLHk3OXA/r7ZBSVIoOovqkq7h4IX
0ogN+izEd2T0V3ReU7zITQZiT0CPfEKoK/aPGUwrir0kPViauunVXyuwYzMzrdHZ
DPTRmNlp2stCXltQ5mvBwNoc80z1Ci7uC2PZCc5fvd8D/7hHyh5FPFNyEBacLXTk
w+EXMLBurunEoyf5EOn5QaKQAWRCnljPpQngbmk5hnY0l0K57xfqxYlgrRYO3FFy
xnkN1YRj9fxNTP1Yj/HfmgLnR59MWMaVtUASnJFt0RAbEdDWPal8Hc/87qjJh6PB
9Je6/ztp+HkLwkp3R7GahFk8X3bshr3VRlTXY7/umhHJ5mj571BU+bTl10v5L5R4
RCFpua4sDgGEWgP3MjdNq1riL3D8b3dsCrOOghOYMTaWOOnuYbV+75Bo1MugcOkU
htRWOMaJe23wWpef9JjJSjWmhuLENSsOIJOyxC2IbvWb7urBmCMWbbkHEHxEhT/m
t560OZgLnm2V0zqcjow6I5OP7fS9Wi8psEglGwshgyi4Nw77wjhMGDlZi5cj3QtH
b6z3OlF1e28zmVYU87wtixVcGvmsVFnGi50z8Gut/84h7LaROEcLKzz4KGqynvTt
3bqf3l7gK419inso89rJ8uSSDggeeV9B4Mo7FvNmxxg4hX9jzDLxmzGAL7rKz8c8
Ku8RTd3B3g6AfwJjK4s5LIgErXv4gMIc5Sdu253uNo1F74CfmbH4dK5djvhPnrYq
XhoVc03zOSBi0A5RAd43NF2emLpjQQEAYjkeEodXXerLNmJGAnzjJemtFmbpUNqS
MIQiGrrlzdVbrq1kimkmiryIFbxM34Wy6IT+rCN4/1bmb6+dyev7uMujqO9e8T7f
hwNmkJJrgtwrIdeeqWhlDlORUJ/ePqhyUHAW/2cPY3Fb3GeX1BG/glPKtbx8mBzA
kmGT4XkLLQWBj785acBpDeSS8p/CypZcjE/wd93I6eZxa0SDU7shS9S0saaqoKNx
hxPBd+AaKocDAf/Ie0RdmZdAZDkGDWmXobB73x2PQfg0hjneVF3GOPyPLHYeu1Sh
BOH36Yp4GykeY5mRInlBLVIMJJWzB+iHm0vlnSeDmkcNOAc3W3nh3/ctjpXOk77H
m6JA3xs980X/mD6QfWuerpz4MyhIzA4BsOn50fGAwxtCuIG4JUgGZj8uLw71fTnM
tQnqqiP/EoA32Dmrzd4m9ClHeyRn1w0A0cNWyLf9KQYeGpdk/MD+BEyC4fYTmub8
THwlt0zC5Jje9oA+aF9DepIwrSZBVtK+CvuA5y2juEwIEN6GLzeT7WOOqk3X7iXp
o3jPWL1Klb6KkE/Eu9FBEi0hT0ouAJPSjLS3m0u1X1sGAaPtSApCnVVckBjpsg9w
CB8ClWHejCYAB77t4nz8cMdKbeAWluc/x/RaL7YpvBRr7+eFD16L4FmQh4AHASw/
0fSxbMf+vONDGxU3/i379bT/QoyiPU15zDi8ZDn+9SZaTEcw6NRlIz/GI7+TgC1J
godDLdy4aKF2GT61opD0M0BrtkwMNVzSrNUWCpNYwL9WwPp6EGJL2VX0PEe8Txxn
lCONSqJbbHqAiUnONxDE+zfkbS1DkKT5LjPYMgGtTaSTzXpoHicxm34PCEJGwPx0
PxjBPh1aL2qpDi7DQPb9ns+IJluwwNK00Tb/5TVzUfaQVSg0Zd6G6G7Dj9Souw9g
dnqd5QmKewI0h9vy9flBY5m0RzlNTCkGtwSvv/Lt6iuKYRYSHvQUh4wlMcylRO00
E1AQTvT+JPRC+tu77RYIA65k5axbn+ph2gTs0QbX3w8aiycmDHmhkpcvyvndCglA
mn5xRYb7V6hUyTRuGLE3rW2z1hhmXp5C/p7mHT139keQ5RxFlwryv3vzxydbLogD
xyuV8LCVUrgZuBeUwFbi2QJSAIYAkmiOEJh4fXVbCsM4umGnHwG+E8iwORn7dY4w
yJ3NkMtW7JZ/BfW9GQ6P0UpzjueEVJQdPu1sTeONvgkM/tErxYZUF56bhl5T7pRp
sXt6ErYEo2jhkTK0rK32zHWlJ/m4TB6/zEXMrpha0FRMySgKmi4fmKHTsovYT8Qz
4OoL6WIun4zlxBQ26V7SY4++JDesYF2ZFSSBqG5q1yzEudXmABaND8H5G88I7sOo
TrhYfh6aEdmldXM9cXRiJ25+yYhTf/b4Vj332jbvEMojwRjIiTZJmpBqJOV1E1c2
cROYz3Jrm5x4plTDjxZz5lBp+kBNP0XujKYbNp3iBO3oC1/1XMou4R4itGfm48w8
GbGAjunLxs6xzTIsQr8PgvemPNLghULd65s/uGG96vYo7pfrxcRQVaH+GRbPA570
K3SPWd66AchLiasBljbl8DkrQKm/SxgukR/Fn+3j2If6uZfilzDDnLkGSzkUPpD3
Aj4Vxwpf8dJKMi5zXJNs4OLtW1he+ZqZDBSrzpf2F4ZyjRZNK1LnjfkbmxI1uyKZ
CjdvC8VaXXh7/88rHIWRQNuMEg3QOmAQzauFQ31ETCiYhRaXtpPh/54AQ7HBHN48
rr2LGU+emFEA1/uNZjtHFOMVrVrG0XpMo+Ys1Dn1xe3fEXvCI5M7SLG8/N7VkpsT
fvx5OKVfy7bEY+4JMX+wwgPvSXt2ih28bXNsTuFkJUid8dpYjPnTtEfJWvfPAQtl
FjZ7jJfA8LX4vcC0fgyzSl7J0rL/H8H2FEwintGWzsVoekHS3W04ERCcoydrTLDA
2FxPpnzTBoW/bscOW0qzseksAO2jxuXkBYq4gaFZNo3lf9JLZdWkV4Yx1ns5wMfH
uTreYRZ8OTXSleyNGkSaygk+Qzgc53T4ufFDD1fpHDrKw9GlaJ03q6LA4XpmJFXf
d9Z8+EjqKulOP3zZbQy4BbKLkxHtNSPwD0hO6knmZa/nAnZTRoiI3AK4+KlU08VG
T1ffYiXfhLaqEVGXyUTH8rjbrlLn0Ay2DD4N+LwDSgZcGycQHjUotuOxImOgvVLf
6XmCWK6D7rYLRtsYBmwXRLw1U7T5KYkcqHSqSBGAG1g6l/cLF6O1P8GVidjNU26n
LpRxSTpuz4BJsNU6dpywwDrS4VYn1bNTfwNNIj5Yfmnr3clJUgPWIPUn5pgZ1Yr6
mvnIRvCm0S2k/NpK7o2/RvyEH7b10UuuDnSsOmNIR7B1on3hZxZ7j4eLdLLUXujS
03TPxVlgAfQayCyPQuemEEY3g+As8/d8SHWykht7Pgr9t3XTnb0+Laszbw0LhrBx
OP3vGUn8ID9NWYUyUD+yqONLGy7Dg5EkpuQXizJk7goNS2qp0GUPToKfVh072GAJ
SNaispzog0NRvN0R2GqOzHDQUgSvA9CbaIQ5zNDAFwzDz6H8cScsja3u817rTFWU
Izzy+XY3D9YkK/LVN9aLtOvFb/cj6BG134tSGfEkUs+V+EMAzZja4R/0TFJLZMog
70niL6rPU4JnVC5DRee0eFTBanO5XB3kOGmreAb2wfiNRNbVY2wsTlrZ180lmFlP
YSowGnZUpuyyRUa/p4UfC4zLhe+hDPlSpSgP7MoOLiEP8JvkJF+r1mrJ7LX0N6n6
CH1FC/TKW/K0lb8uAXOn67Gan1JsxqG4dHTHj0M3WQFSv+a2C+gCUzGgdh86yiZO
JIMAiSYpvfsUZeDR1+08dSnXCpgj0R/0Pc3SnyTPbqh9j19BmmHzFXLYU/XPr1rV
7eKBhu9aUlku2vrOx51OPVx4eNJBwplO8pPuIL0BV21cPG6iVcLReg3eFjsMJvPW
P6PxVF9GUeYvI18vOgTIvCFcdJb8cZqxW/8oCnJurDSxXCWSKs6etOXHJyXaJHPS
76seCguqxHZ2K9p0D4+Dn1qXf2YfwRMya0k+eDgtStW5HhDS51n82mMXifYYku1e
xVcQDMON4UVn+iMzL+GNwEfo+BxmrkM+Svb2Nd/eGKBkJxAdcl5HVW22BCvaocqU
89s3RVxhvNgTMu9NKHLMTCr5DXMXfS+QXTNavU81D5hLT9e1B6wJx8iRBLyyWysl
MHmViiOT++dGdwT1SsGLVu6yWqRI+c4jHolhSnCHdXQFMUpsKCEhh3kmWIpOCJlj
A58k5d0qOpV9HTMwSL0wNn4dAw60aQuDc457Nl/DDQS138maEHRZ2geOCA/SvcEA
y3P06sml34j91RE399tSjQ/ehKbi8IVPlqDXw+LW8h7k3u5dnhba7ZhprF4hh7vu
C3QN82DBibMxeM7rdU7e82EMZgbUDqVyAOJT7XvCRtKwz57efeL3Q/JwCI4gMC8I
7vmTCuFqSGBeZuqzwZ6hnXuXWB8T/63MabAIa7SxRavx0wxS0Od+UmhzFWB7dnN0
QbnKqEqDJj2hHyhMF8GxjN62y2xvG88xUdhcm8rZWxVMVrNwM7bfuDq65K391JV8
q9AApzYVpdQ8XrKpAW8lHttcJKYrs1gqZtwJESnDd7EL/rGOmFwGarNWKYVOmprz
H7TjICPw0PFJxTK+5OTi14HRhm/lGx0cHBjRpiKbv6HslvaH36973w9Pr186ke5j
A3i4GHElzkNGj0NajV6ZyNuzFtQRpPNDcQYml/zncuYmpC+WdIm9NUJxzuMz3cGc
mpIqelTEZB05qOpdhh1yAxGxBBIb9DXDyet7n9EVywUbQzUIDCoQyiH4sPWbfaZc
EMLiAUOcytWqU9wNpia7HfUsUNzdFpoemFdGMh/btbQ2T8e+4sBJo+raVQUJ31YE
Olj5c+CTNKe41DHeSzPsyQUCTF1UNGLZtyKldumiz1qGeRm52hLT/ugs7cTN1QTy
plEmOi+yI3rFPGjSIcun01R/qx1XiRgIE8h3GPuDGG18z4ILah2g4ne/RCmCl24P
5ngA8HgcP4N2CHs2Y/1mEflb57U2jZQZCTYmC8fVnkWMdGO+fE+j7eyyLsWF4VTO
9gVlBRKBHLPG+3Ien44T/cW2Nhth4UmYrFQvIoaHjqvkotH3l6ifwppvpFA9uPJa
7O8YwsDuGBD0216XQXHXGh4cqOKnuzYlXPyIL9BPSWyEZKIdIPaZZ22+lFV6xb7a
f5CupTAkHWxEzxqjtKnadkD4XBLZVzUoccZlGolkrjT2vOO4LmqDJwC0Kc5327K9
LTfSeZiWAajhwFHQll5amsRN4xcoc6YS74yVxQrGy+F/e6STvgmRs55XXKxSnJxp
QcPlFqId4Sw85d1RTVsd2ULwoBC+zNQpF1PkFb8vWKARLayASEjEK0dpEj0Rgbcc
NzPosADf2YoT8dAIBUxtP6NxAnOlB1hsMzhL8mntGT8h/ChVLZquIYuE2CrvpH4d
6vUNJWkmc+PMMK3LMckwv0KqAPbauzbQFwH8gu6g6YmYijg/APzle7R6WSUs7VBI
T859QISFOqdCFs9DxkmnyrJitlNmgo4xwHkSxVEiBLY3dxgkpb3u8yJZx7Ibgwwk
426DzoWfmQlcxUIM8EFwB5wBiYPg0DgSg18WmlKRSGGcAX5slJjziPOLUD01k9Hp
Rz4PVpoibGJ5IwAhUgca+FdQy0jpbWk1nYXOTzdTo41SFxuzL5KqV8rOU1yTNQ2H
6197GN7pFsftMjb7abTKc/Emd2rOT/VzqjQdqe+wv5KtNJe2cu6Nujr8KgDfGcMI
042MipBo7CX1Jlft3o2VsY6uPQFAyaottD+PTKGVvrl2SCm5BqtYIEQt4viGxzRl
+x75dKTbfGVHd8PB8p3126tmzqi6lx/F5wiGzaueg68ZPbdlYphmW3hfjETbUuQu
exegllCkltPXDtswncY0SEuLRBHXfjnW+qb5fRuMBmdTCygaDXk4GApON2Z66nuj
KqzUdpABFWDPOhChhdZ2cuQT3Ce5c2YuY0vZ+TFkp8TqMQY/L4EVjuB1Y8lid8h7
mfN8C6p6Tc5Q6Qtj+ynZ1PuRQe1ccgm9WHh/jYBfGY+FsCvXerIc5GTL3mk2YCkl
EzeLyqIN49eYlHTnsnfoBUi+H17B+VnHcdfa0pUCyG0Y+znUPbjCbQLyMAheBvBc
G7cKWLr0IrPPC8i81GFMwdcv/PjjAq+J2PckFaXkLcW+KzhTskdVw2sql79IpzH6
EvHPGLrfxOzXAF63hYjypPl4/Mrt/T4TQ+y3sKvzXzdbs2kiEfgphgtVH6AkMYt0
YDTCuD0JVDAs6+uzjQbOBtKXB4omVfmyMxaokGk4CAGbCjiapXlpZ8l8/2fuWZUB
IaTq46iiORagllMNOn7j+JANN5yAsJ+fwKdl9SvUqUOK7RRo+YcA9zhCSio13EFX
rk8A4a9WNH/8oJ8c/bXatSwmXTjN9brrC7bgGs8trdOjMgnX6aNY+HdO06a2xyk8
+2g7EHS19Z9Z3QO2Xl3dFrxn7+F8YdlRf6Z8FxeCK4zw2hRupwzaf9VF8yYfiqJH
y8HNHS8S/YiXMdExg1rzKbzKDZrpKKI0xOTNXboygzy2ntETss5rtwbffJoR5DLQ
FVGq0PBkL5uEdGGr97fW1s/GnXw/AkozszzM7RBixseo2Sm5+6Q1/f/6geHpKWI+
3qkCEX/ufN4VNMS11MRglOgN43zB2fBLbTIrTExUQZbU1Jt6qz5dSfpsxGfFO8kS
alzdev17mbBreLaXa8ekLtTuFvZNXOk9WVA0kl3TvmEGdpcAGJYMx6BoSiTOUeCN
s+g1yC/JqFzn9w+gk46ogwIiMlHKHGt7y3ce0rLKyEsGnFViIImO76xY14ASlmyA
7XzF4WT5VEoIo5DS/NsiTjJHk38yDDJh3IB7As8YommjuIc6yGRgQcntvBhnZ5ND
pRhxtAPA1/NI5eBi74m8rqTex3Jy8oWQ1cQg+/M23czBgDJL40abxrGkh7rKbRUI
GRI5iKmhFqF7BYuCuUNQJ7TYsPSh9slVuzGmvIOpc/6DoJGw0DSMsF/MykeNeSp2
5JpxCBqgMtYnWmigDIX/5FOhWOyaDRM0+Qxh2SpQQ8vOxW4/eLXHP/2xOSv1TFNz
2DxdwckvJJ+lTmTy2iSzj88BKHbXh25VWDblduR4imvsnP/dO4c1pjxCMoDvcQvj
DiiVApKijYYFYSJNxGt49+4TReZ1OIoxfi3c8+R1X70SLKKa5Bzbs1+HG/IZJDX5
LDvSD40ejtC1h9d46vjBcWSjTIGylgLbxf1BteO/vhXVqPoyjbLQQDpe9TAfaVxg
i50OJxE2ImFFOELCOERyk+4UGLz6LR+rJMiFM2vy0WKMRM3tq3SbbWPATgj7Jn7l
6wauUuKua7+FybI2lT+bsq8tYN6eLiDZ4ajVY8p15nL5vV28FhohxShKxiHqAYKg
cClBY2/fK3OBY4sledtuwuScrOy0x+P2hMhK8Wg4uSkSDesOCKa+/EdCqzpkwcJG
BBoFDJr7/v+sEt01JOXyGqmNRzQWROyrhvo4T4HnCMyrkoBi7KgEC/WycSHpIYEC
wvJAMuCRBeNbQAJL7Y95A17FL+luXBYJwXBTBecQD7Sl89TbMM8uPMYZgQgxQZT3
rUkgyhvxVTPuDV2MqEzzcO+1l0LaAvo8ZRVP4vY5WW13RXe1/SrAoO8o6VVTjzxS
K/JHqHrSWN5MXmgHpxSKy9Z4vZE9cy18XBU/1dV8oX99xC4zNzQ5h12ObCbRT02J
yZtB1Wl+Le++0D98VVZAZ6j0fW/zUZ1BwWFa0ZGEC0KlCqzd0yy7D7y1EQ2yBs5T
JikGHU6u5WIHOOqSafUPmW2Wpzf3Oxy9ZxqqCtPoXpHxvuhOvrmlCRqCOCYDJE1l
4scvaHp1LSUvvQOr3R4TGc9Dz+8AIP8TNoeExxfr95CeXyG3evb/wma1JLf2kMlV
ba4MVGPxD6zK+fHfKKTuE60/aS1hNIDRBZCL4IRzPb8J7l2w3cR132ancxT6W1F4
fd1BPW3gabggeBUWSh0oYZkpfQn8rUdlGpqCvO9Z0bmsuKzHGqC0OX6SkU8JVU4N
O10Vr5k9Ng68WhvBNxcNgBSIFwutjMU93wvpkrh6hivRXyOTY6TSp/DYE6BYFeFz
Fs3J5qicL9On00dtlnMLrx140iQiCOnOBB8908lJ3noC6Lri9ExSCKVuSuhRBBCF
5F1aAtMz98rgl75Ace5hLb8nNwMAHpJoZe9p2huCu2yK3zLe8arONXmJItrUki1k
6Nq/SyOyCgfAPHMjUwj7/VCg+1CM3x+RWYvZAlbfrSAg+GGhwD40UauPvvJ6AuYW
yDBDJE9EumEUnwMyey1uKpO4nEU1EPiAQutDfZJU/h/yBbXhpOkpI/i5RH2uQHIV
yf3mNDutSPyjKst0FAk2IJGTZJgIWXUuCJtdShGLTHRCDc2yDjMg455VXxQ8Upuy
+kR/C2RyDWmQYDTs08uCsDZ3TN8cobko7H2ukch2q9myv94BJ4gKiOriO2l7aUCu
YoDjT1msitOFaqDGhNqN/zrAwJwzR6xuEFZN3qMFFkB/J3EwI+02WeGZX9pfOhrl
9ZJq69cgYgbnE6EGk52S3hH+/+gZ8NuyROfDncIvIzH0bqkpI3iznhSQ2XBEUGyP
JcHMfir9j8h7qTm6zhpRbSgwYARg+TfCXTZbOwEjQt08cgjnbrFex8IJbFaL/g5Z
MkM5HeSYfiU74d2crRrm09LSKqzQu+6eOcwvM+hbToj7IeH7zMxegRm7KphK3hfe
602x34iI2UvNaH9Kk4BiPP4Mft49CPYufSU5gbJwcMPqDYnwyuQ2e5C+uYyLOdVj
Quk4xmzL0BcPJvqv3X38z2Trit7BTrk1RaJJQ2MAkF9RVqUNgloROOYPdEJ+IhYg
yK7bUUEaLrFH9VaNcHs7rl1/k9YqgVmROsceiEgJZ59OeGKnUNx+KNs66DDJ7vhm
LlxAfJNvaQyRo7cZ6wn795nOVagPlJWrnB45jIAuBTn8t1G3reBOx9qr8HRsT/Ye
JFUL8pMrxZgC03IG1UxWtLWTRn4EN623ptlzA++0vqIU0gXXgdEhjNasnCtZlGNl
BJNImGTLx76QO3nUxqP5uFeJAS6tSWX/Vr87MYPchvG4H6nbXpBIaNPEgNcvO2oM
JwZQpsbgwDwJfO12Y1GhQ244TDLFciue/D40QxPGGjsP1kXTeef1Qn9f4KdsJkSY
rd5c0FmKFLYIfSYvnX7zD3nCopCizuoNZgGUlmq0qKqN3kLZF1x/Uq4eEQ8qNdGC
0/xYdC6v2JRk+TDzqc6fk/Rzl97se9q+eGT+mILtjfM1z+xWPPGXYPURvoOdMfD8
uPKp3qhqmHhtTqWqj16eRMqRMq7uCSyGgFmAC6PzCaJMtIPB7f9vBrg7Wc6pi957
gRiWKYQi0cUk6q8dQqeF6NN6YGci8Mmzjq51vlbz6y5zCxbaCWiufonKKQCIASQC
GSoY1xINh1kAPfOMgMTjWhYVu9LjCsecDVocEvAwkkx//kYDIAYRFrcPGcd6OFJo
vpwWQoau34PvcOhpk2WpB14WO9aMk65XuFYBzaRkXTx7knh+yQFHtuhacueHAZ8s
8vJDoL3ZJ0WMIK8YYsSwg6GQAdLqkihHPPB+sdmkkVCXWXoNsbNqMXISVEXw6ySE
g4nXQnX42Rusa8DnRkTTEworEe4QnZJ3qLtv/IRL/KPsSdhPYeDZ56M7KIZQtT3t
dKC47fjn5Ds4ONxTGGI2ISswjPd+aPZmSLAnrKG1LryM0G+lDZb7F7lDXCZz3C6d
oFfOsgnf+oSxNSwSAMcuu66WcB3/ifUZ37NpTEX3apYp7QnWw9Yxmq7CA66a0aTT
YL+HIv/ZvmIyTeOyhPWJbF6iBrWdUicOnb9Rb5tdtNwVcVXwogBHY3ZSmXAzI6/P
f6vqUAn1po+5/2jP7YJeRkIMLVXkb80hDpWfT0wYSDp8mTETn1JADj0nxa3iSSIz
h2avaOFMuXK4VQrcK4F49/UySBMQPSNnL/nf4UekYBgSgxcglNrcZls29yWSF9uT
HnA5ci6CPSkG5t8D2cnpoxcc2sg4ttp2hCV7LJxg6iLkxo8DVzjz33+k9I7LLWKE
sZChk0omPeOl43UlztnKpHQsjOFZooSkHT4HqGcpRnd60BXCS860iefxDw8JZ2pv
3XxYsXMVXMvPNQvrMz6uPPw1uQpYPiEp2qQ+K9xYkC+XGpMHvd+QngvrgkR5PwlM
iQjzFwz8N7oxzyU4dgrkrjCIXaSR/iR6CHMmBHBsp8ti+06SpXI/fNYp4rz6cSUa
5slinkNVpWLWaMFzCsPHpfsJUa+FDGeNWC/aVkDl6RIlcB0iszabJ5xa00MzCajM
w2WTuV6W8WvcZ+jAw2EIsml/6OBkYRun2FJOUn0pZ3chCB7gvCsu4SQLN8z/2DoS
q7p9mk19ie8syk0vaWNoIGTdS0sWUYe7E+pR9pQ4DYa7wtIzdSUtujEWOolwzFOB
Qyx5YTplTIc2qD6jl6H1tXpJoSiKQrUXdR1pduh07YWyCV/e3GqlpCHiY+O1BIm1
2F5QK1G3mV4PcYNvwAsi2y+EahfTBZhL/VnX4b/Mn3I5lcDj3AwD21zLdDHxAgOo
7Xbto3ocD6t4u+5vhonOZ8JnKxuG+lN4XPk3z0bPj28H4uJM33rWVALiEzSMRT2m
Bx9Q4CYNOfwnfcEQ6r+0WaBuk2TtLRPpQlbu3GJ17RfEW37vijqGYFmvVD/t8lT6
HHiSoyYCxtOsCw2jpWC47WQhyJfKkf3zmapsX0ldZESClQtQN5xy39Q8t5V3r1BD
rCUKS//z9LcNZLKKN8+KGH5f77cawzJ38hMbJ7m2Jf+fy6xUghaTWp3HwoZNVJ46
tBCEDNgvrdaN/CIXchDg0KlfUFvHI/HpO+qUduYYmcXlG+iKB+9ot0/5Bb+vR/nV
X9ihehD7XrVC01xgYXXQUczbHrH/CVcZCPeKykY67DaSmtMHf0qFVwLHndFJshxb
j7PEEfh9Tx7zBlNaJllBa0T/IzJ1QUU4xvM0XsFZ833j+WCsdFIgyuzEO/uNmTBp
9x6/KDL3uHYqjVRcxPGNr4MuYIm2MUHkTY4fUABHRtPg14qxuygpUEGBVMoPuO7K
H0uDKQJ8wzb5U6G7YkeD0ahvPzxPQerWUNjmh/bT0MKPk1izrF998zpursu/ryuH
gPjhZLqqNDbigb6e/ut9QGDp6xWT3ME8RWWHfixWpgc8OhbUX7TmrB/TDfVMlHFw
nA141x0X2PIMBQSqcNFw+K/K0k0LeQxhu66QeDtrFZPfQTxePwA4qx/wXahkLRQm
oM8Tk8T/gpahpb6aN32rJO4gXhEh/FaPKmbiu1X6x8fzXLv8+fY3nn+/eDYePhGC
wRq5Ug+jWi7AbvGlbXsLnG8qy6tgxIVAw3NYd4/SkPIoc23WWJdlH9oMiTQ0py9y
XVq+46GEj3pc9OEbmkeO/AiiPzaFoBLeB0ZReMxO3MYs2jJaBLuLI1pXP5zJsVYk
EmBMwCpq2YwMaTlCAT7e8XIgDET6Rdf96zxVEqgnBOnrtPM3NHB+0dUxxRMbKF2o
nZRRpaU0xd3Q85U4i9dAJqMp4RR6omRFOUHiuipiSUXxm6MB4jLoFI/LKvv+gH3V
1evMdTlly3MUrzAj7DV7zCPbv/9ofxyb0K05B7/zyjaZ/++pUBLe6wAMtRm6f4RO
niyZrHzqun3d6qoyDYQFZZuE1csQhQjsx/VNnrsCzm+aHgLQy660lpYMO3MFRVsS
AWseRRFrt6jPeNw1yyBGGY1nyDVUFOi81+mHRWJvNVeUuYtSPuk5hgE7TX8PuVUU
KSYCTJSBkjAU1uj2fVU4BkcequtvrQAq09WF9wlPpjGo0bjB+F8JhBXoxls1J6LA
dUPcWoZzG9e/hdUGQpZgxJxzUBencR26aRONQEAzU1wgxLNQRVu6gp0nd7cePcTV
9Ew4clURZr5egNHz058Lio70oaWrh9XYQh3oyaQqv7JRnPXvt3gfnir42GDm2dJr
7cW+OoIq1a6qyKelJ34bxkt/H6V79dWXM5xyfFWQLifMtUk62vyB3CnjVjTORs3R
rdR0x7kKZrUvjC2DLYs8WZNICtD3m2vuKuFSl0gk/0tL1YPY1etv2Q8O8rbx+PE4
6tHy3i8B/xc+84G4UCFWOuZQ4z5l9jCXMDNE30fs3lgj+xx82wxhkh5IFx3VSh1I
JH5fz029B0dKvIES4DIg92vs6/RUGEAFJOYXn7OOqCic8LlWTCcv50UiHAwdwS06
pbV5syiE8P/rvztc6KAfuMBCQmXR//kN4vWDRNOr/YuKye6mzQqOKQc4PmrqkD9L
vbNYRnwGXs4r8U+5EbAD4GG/7lc54ECoVOMYrWRqum8RN8FuK3Sxtxax7yqn9Ae9
9KhAP8dCHFVxNsg+HVt+y+8I6LOHfFFepvWqKnOaA6U7MLsg/4uY+6Ca/hPYNAl6
K6HGAwj1j2ta2g2xruPZoszvWc1umjY2WBddZ+hdAPG9mXMjtJuRPkjgdHrD4eKt
u9iZTAiQkIkV1GSVMkxwTuL5N/QlAVpILqJWogkm+5FSurF6rLBL1jlB9CkRFxWP
r6tEJNxhpVdfe1SP342P9Cz+Cwrzd28oaW0kL/H06WqvONWBKKDfGbFuAMKdgvO0
kSykIEaDUpLSmD5GEk3XA7hv6vT9JIUiEGuNd9TwJ6n2le6iSkdj8Zt7DyhH8D+i
cySxspVpexoxMDsVtpCuTwd8S0g0qVAKV82zqxLDNO/SUyGmwpQNlhoZo5rT/2up
IWY2sHJCNYsi04kAJIe/oc1wWTDgev2xRqK7vnDIEm5mTuEviPPXmRO0Hh+xwESC
vPAKq69b4vRl7nR0IWb3VzlYlESB0BLhcIXty28Xga71i0Q6kxo0+gp0VBZo9581
0IAeAcfwojfajJSFDyGalVd0CFwU6LNM4B4SBhNfatf2kLjDRFvNpBjxq3OTn4Yu
1jWY57kPIR13rCdx/n4Sqrg1PeX8lXnDJWLVJN28NlIGI2MPSX4Wy8Qv7Ow+kKVK
LiXoGQz6rv8TgPflI7s2lto7hkc/TAEz6VoKUKE5W8u0Nx2og6BWHQJOlDlcgKzg
1+QUGMkQAqgUsvEklxkTX8q1nxmf7arI1gMCYcByIkHvhVen8/TLZLo7oFxmfSYe
txiE4G1Fj3/UUjS+XNlH0MQscSRhh9PTGsdbEXYEIYwraPEclCIh2Dyt9hWJgom1
XhWLcdAp22cXkEsAqJGsY1Eor4rBZtQp3DudhoYhvhqwPtTswohxAwWUAPnN9+z8
zyZHGXkI4Xaa6lFlhWLkW9CsAtq0TLoyiNwcsGSjySA02Q40BrQWW8VFg9JSD4/Z
xQ5JTaKsVdyUJt4JKPi5m4P466vYfXCkKHGJc1JsRXW5flOZ2FDPOejhNz7HqDYG
S97hUou/zw3P7euoL1wINOaxhCWh3pMgJ3lEGrtAnUkBJ79KYshUP9XSD00SwO3C
xptkgeOK/oA2hN4qsBEz+JcnMo0UbbZ1WhS7iQmqBSau7tY4ifSoH6Jf3DagE4FY
u2xx2cHi0MSweXNtQ386p7UcRn7NAQXVE7CWUJE+VqtLfq25wBOIauH3JRd/N5Sd
pBqJRwx21UUFsmfEM+dZLWlTsNRZ7NdoDqw3O7+ibGVmIGt8aeFs9srDg1d9vg/K
SJA3B9Um2Hlky2MmNcQdyMbxKvoWr1L3g06ogswNjbd53BESNeHo6UZUR1k5Bc2m
AAYmkIRdrxnL/l46qZzk9XATnritReWJFm8+ttqreNC0dyUsglSxTx0Vf6VCGP/5
FNFMrHaYsVv4VRe0EWpJ5uLxAAGFgty/+G4JyX8vk3tm7bAM1rZ5RCytMg3Rw00y
NQON40vw7WvANAXflvGwCMcpQTsfab5AxiMIXxVbxDV8jXkFz5h3cSbjkm1NWL/Q
kEoBMl+l38kKKYDZU9FTgHIOkTgEE7M46s4gtrd14Hjgbl43kxiZJGnXnXleB1io
lqpzB/d+/b0SIhqUXbs75j047xA6d9mz1EEljcXl2F348vQ4Zz+YeI6IZU3UCTpx
3gPwP2iE+ReoQAygB9nzFf/Sk7fk56hIrWdJwRfYHhTwm6Hblx6zzbnnwA2ROAAo
23msUQLQMjQfashUbKZtY67y5rwApdmEV7eKCJA1k5xWmEsrUDhfh4/nrTNDOZ69
Hcax0WR68SyEVWquSbacdBtGILHWx376kLfuxYz9hiCdEaTCUwiu6/G0kbzWmAnq
DO1uQcHrkYdSq6Ii5cRGP+6nYjAmKC37vLhXQD3Rq0An2iPFDdXJJ0RIujBHwJUt
3jBjoGeXPjJd1LrX4DzUzkVE+/RYzOalfH2Vx0KkazNb+U5epYTwlFxRr6NbYw/k
NYM4chQZ4+8/X8kiJ9zNYFO9MJZR5TrxBU4FHQxpPFCaKQwcS16y7h+D9Vm+epzI
3i56n4Cx/R7cnSWW/arQjsqzIgVOZRV9xXQzAv/fT2UqqAQOLQRiODSjFDg5waHC
Uys4Gkawa7wD2TSFLUesf1CY54kKOtwsNFcyGQNwelJQP1RD8Jh4VQEPq6xlapXX
njEh8n0Hf8i1F8+uJcIPGSnFe36pZsPLX3bD2eD3l96g86oRDt03gdZe8Z5zHCZC
I4Tl7gUfl2wDrD1hVqaf/WF+6IemV/Q3Laldq0eYAP2+kBT78LYryGZ4GIV2t8ge
EIRninqV/06Dx69mcwU68Cn9sHcAVGXoFYNOWu52LJOhsaYFEZTv90SX71m4FMy8
Ob7AIMfcCx6VVqBYuzypBq8bSCNgug11yFaO6HL3BiiIMl0qmg+TBM0mrdo3MxT7
57z0RMCuXr9YcGn1i1dZiRe1MYhKXQS9bHuKHILdP7vszF8oly0CtFNW9s4qBh7b
SF/UmheTxiNQZ838OwTE0utz1+jMB74CP9gaumLRO2z+JFpqs8XQ3GeTa8sj86/5
w1/yNRokvMSSzsNWqCONOuNurxVoI8h5l4ZTXHwDEfW/+z1O3i7yGAugzyoGbfZs
uSqSybZZZyDCDuGyhiUAt0+pCXT3bF1vQVdcSCDQ7wxpuk9wka5tTqEwpA8Qh3LT
XUbMCgK416I3fwEpAHnxVDtf07/BBklAKVGxspyn4ll8/JV+9vpj5gIWG+Vzaz5p
BeHKhStr+IhRoJexdVXa7+alUOTLSqtkjculA7brjsF0lpqqM4lHJvApQZR0gnNc
DyrycFlfuVrSfHpyOTbajdxwMWWsobpOGmX9zs4iIxf4K+seT0QoXksAoVqCyjsb
9oTbAMezyMEcSENTzG9k3zMCQNhudA8REDIUQvLaIbWymw0Ja6ek9I7Ee1lw41Wj
tW5jyh3BqxW/20fGLi97R4nFJADaarqccQQ1Na02GrFAFzLE8WjK1AJ2a893+N2V
mmcZYku+WYRVO4Vkog0pRgfZGHdCdftzxhAcTeJaAW3dyaZex0m+NMJdzrYwUyIz
KMPN/FYtrroHkCsdWhWjOScVXwigF/FTVqIkJuixxapV1GeK/A5QLw/5OXj14wYT
LGkuObevqRAWZHKl7LkZAEe9JnWXv1IYe9f3eQHlZ7/g6jIArNqmvWIa/bL3KA+E
8+knEvp88YVuKbd9MmvT7y333BzKfiJU2DCCNelWlVsjxR1wLBwDH2rEgzMJ6lQ7
tR+R/ECZ9N2wEvZ7D4G4pZMFaw2C4jnMIO+sfAMh62zgn2MCCdCobRV7Ky2AjAZj
zQ3/MVCG93H9me8S8VHuBi9XxmLnwZ+yqCwqQnFyWHcN2X3sdfg3nmnquXPOJ8YO
ZhbYmoZGTP0hUsuDcYgZsInE/ubc5clKRu7T6gVflvoTrd/EUhGPP21Mx1jTNN3H
11bqWzG8X1MAiTplq2ACe+Qv15jSc6T3oueVexE15Hagq6M3oCdEmUNc/vnIS/Gp
VNeAA5xVfPps9faUvh6o3khBb+wAnnrPfZ78AEdP/blU3w2TrGo5EfgAOvvS+k0b
nNaVSq4T2Z6nmltbnhWYfDIVh7q1PfU6Dt3Hi15EYwWJ628abwfa5z9dqNU29k2G
g9G64+VKiXcU057y/5JaHJcnhlp3sbuS1xsw/8b4yIS9cvTfWrFYScqAOOuP56Nh
3coSJW85aagecRiIBlwCCBKs492frrbzx5fGaEx343v8U6Hk2J92ejuuxbG3B7/J
sDA9zNHwH+ZUkuuesBgvNWcGcjNrdETWXn+T71b1PCEv/Cm7Pcm0SdZ4cxj6x9/3
gZqvbbXWw5rBtQw3IMI1VDSCBOs8A4S7hGSoyfRRRDa7VHv2xcUj/mZjwurz6CR4
SphAu2fssJVNpSypCTMgJtCfvZU6FTh8+kVDdBE9pyygHelhwdTuzru5VSVwfkSO
d2/EPIdIQOm3jhRI2ZgOShzBJ4j2KP1bWWs9LVM547Oad18jJVpsjaDl5Wj8C315
Kc4gg4nJCxcKtZsD6jqgKKa9UMo3qFu4byTTNwQguyrK+iiGbp1UzE9i5QhVzyKu
pWDlHWZiFnAOGrbzF3oR1dOp0gg8ecZRmUFokkYsFUOcikuEDm4vdpVjekGfmHp5
UCgEWWQF6AG1GMXDX9kr2ZDBq2Judr77EgNGuULDj8VMDZ3U/usjckUCexx2l5k7
T49IE4WuLqsYvscAnTGaQ8bcjva1f9D71yC7OmdRiIZSTT2pVvIqcokalPqYMWV5
dJZ2Li8QKeybjq/DYbZMHvActcJ31zDMKGnetM9XMxLx8UdFVnXvZrzlAFYEWEny
L6H1BshIOVYu6rOa6WbkBLlU7kyUycbwdbMIGWqus3M17OrVRJ5t36paxucOvVn9
rUCzZFa3VQ5DYNn2EHwwvIXR5mQGoJE3KQz/3uMlKPgKCz9z5NGqxQBsRLZLO6e/
FhOIZvvQh54DePintw2iI61qac3Iq9mJodpHYA8yOXFyLc4s9cdXwkPsyJZ+TJQb
eLlF4mOUAE0cS4pt+0j50umJEmhC7XSkzEdKE1cIBASwofQrOcE3+kOUX1DGz09u
viOicXPwwzN5N+vp4AbBmbYY76OwJRdCQUS5kDwnuzZLEbv6I+fO/KHUFchIVuho
5MHMpxYgrjg5TC8jEV92+Ygy6opNBPAfQ+ItkxcHwUoP8xUk+C3VFu9OHI6iis7q
rI9W8ct2RBKZAo9ctdbx/YlZre7w79Q1RR8nzpI4+hxJspBO04KKQ2iyVtcZhaYY
ee2H7B50GNR6zvq0oRo3ZDiDmp96pBgtlq4h/cs3pZjZ/BxKoxechl1CjMX/pR5a
MewGSUOSnwCt61Y3IOG+jOcUAubGUD7kLwfCtVKW/UuJtSxkBVjId/zYseoy02+H
6sXYlwWLFQj+a1CbKaqSH4de20Yr/2XJqd70k0vDspAfEw4bwXkrk/41pYTF8PF/
zWH9DVPBc7l5R+L1FZ3YhiER10fyo10lyDWayWVTeioLFosM4Ts+mYfn1jLbn8V7
qd8vgarUvlAdYtrwqHngGNmgvbNEj+OV4FMWYyBnYYDxslfsonxUXMjvY/IoTdsI
Y3SjEM5jnOo4ta07F29HgEMKAkL5Yz4S/h5bsrUrpnHLrG0U7CtfXfUngI45LgGA
1fOC6xVVW8aQXw1QooxtFrgnEc9kHbeeM+kAm1s+9qJ/uIeavSYMzcnswit8VGll
wtySn84CJ0l6Bbi/3yPQFbAw+Ah0GnxP4Dwmpamxpz2vMSqHoiKXW1ZFPZ4mpPg9
+FOiTdin0eTtdeWZ0MacXkTAEcmV/uBSB7Qn0bPyge6Ine2FrUuj+R2pQBSN3GJf
R6dPHaBrAObG0nxiKWOZ8rcf8MOHz1gOL4+92mteF0E6YfGyNu6edoD+Za2y1Zfn
Tk8RIjws067duuImm6IAjIXkwxsmyYG5sy35YM9WqWPTMWliusybWFPAO8iZ90Kl
0v+ujBiH072q0orL++gnHl+tbRXXzN8ssdv6OgIuIwhaAj3AuC3xlsLaQWy05+be
ziOdc+4A8vM0uv2+FC/DfEApG1CbEGyifdbx+SBOaclPbw2RXzolxFKhOws3hvYW
5ToeB6CfQDnxCFdBknzWLnO3y+kxhVN4ZBTY4f0jAGwzLjtL7DhXeC7UFhCYNuDt
8hPbEyr278jcBDyQZ1ukx4ya1SdUs+ZB//I9YWolVd88X1/nROTLGYsXgnAYPj5v
DrXMlmHQvHbcZn0pjQ6osO8xR3OIv9uRkaNIgBAMOi77kLF5NjKszuL9AtB2mtQb
OJ558xQJqRmY94dGIpp2CfjaxjQAmHgzuEvZl1CeMl8SEpVPzjAmBK3iP8R//8my
MvvF0VF38POl8jcRnak5zy74cGXWjNafSgKsNYKODn9TTJBYaeZJDBEGdVrGM0vB
0BENWczAp6y76tqAVorEEbHFigFIbnDbSisI7fRAqM2cZpCU8mQu7s9+VtwbEpLU
4vitM2DuJ8ZYebLkbG3QuHSGkG062j7luqdOcn1g1Bzqx3kLs8v7sGWBphI8ubr0
YEUenrSf2UzaaAY3M8yoSwoeHVzERJnM1aNv98pRHrc9zeNIo6qwqOjxhLFutKXW
5mQLRJWE7pbTIGx9nSkadvvhS5LZ61xuXKTYrB8WSnk9w76CfZdc7rWMhc/YZkZj
y8vhDYf6x1WLlUOlcGmGYI+msQfnPSQBDFTclXyykkxbCr3FL9WyRxa6UAHEbw2I
A4C1pMCQVK4e65Zz+P4Xcji88PCef2HyMApIiJ238JtQ7Jw7bV7UG3xgrga2vMrk
JZ+SfxCTqDs2LxXUSei0qBsu6Pcgqc5cmoGMuPSqW9FPXjPFFIiB6ZLnOAFjYtWE
yM8sRJIQ0OPXOP+KF3Zye8r6R1nZJZMmAel6NgTL72pzi+lctWtt3Jm4gXBMbEgK
u3cod/Cx3m6FOhDWCH6HErzEhYsHeU4zt9xKkdny91SMi+iRlPZSGJg+mo8aUJnG
0wj8d5uzUmhYCk96YCbboj1AzyTVQXKplm3ofsfYfIoiS+ja/uCMO05lYIjOAc7Q
vp+Hp72OSwi7IefSOV6LgPa/3TS8WUG4tvEKNsqFCPZ0533fNhiBvhAUMrTnCXH2
fjEtdNXOdQYP5KuL60ZvxwyH4YXsu/um6XGxBLRgjZuWf0ZD/LQguCQudL/mspJ8
67DPza+8DUoUbh64bsnOrKh8L+tD+YXTxUcksl3HM4ouV/W5Roi/Kh/lWBHCobA2
TODibr1hn24A9U6RvM8yq/aI2ySR1aHCT/HpcZtqjXZsS5sEFDyzAtkAu2JPoKMZ
JB1ReB0k+VaNBwUl8ZisUgEl7CqVUSRbQs2HFEjHVmd4xkChxynJ5f2dVVlsnOYr
JMSTAQAJbqdum8pRkoUbzAIP21CUTZPcXDqiPSfUMzUOURnQbIUTJKrjGYUuuRqI
7ayVq8yPjbf80migHeYmJfcX2mBeVNQIJKP/X1ghhAJftJd4wQ5a2jeDUJwpb19U
LHEp7xmmM2FgbdmyfPZKABdLWuWXTAJL74Vty6AbGlmcqztikKhViux5g2GES5ZM
QEsN0qP0N7wNJsDMz7h2ntGKt6MFrmULsRQsw0EoMELIE7Flrzu0cdeaJDfRTu/k
w90OmNf7zH8Kqb2JIYB8waCAbpPXUBEisfeebM0YZ1O542Yd/RD1IgLkUz+H8atl
SNVt6lUamtThJ2U4uALgMA5Ng8Hm1vMztyjkdHPzGcVMzADxg0HR9o0N2903W3dY
w0UdcBfFmtbM8ViPFM7O2DhML21j8c2TGhNzbbAEhMH4u5PMH7GStf2OGQhV7Em5
ZrlyW1yXxEXjjJnuPhjwdZ9HLJXCHhpI1okgCzgRZRmM4jCX1MFkPP4DgI5bxWyL
ESnQn0z5bSZhgTAkdU64iSLiIbaFQKEDGMR0PBYTRbku6hjeCsPt+6HxuB0HKpCg
jEQLlDf0G19uEU/bHuyh5WbXE3BzEeD5Q0Ug4yCustbR9fdLfdZAV9tfRzeU2/Rl
2LC5r3E3PKlkxFXl9uJUgKkGw9n8joJV5NL4MOJvDEpAbvw2zJK9blcvhUpCaz2a
GAOpzRyj6Dc/bFrjiDZXJtF2h8Vz8U7670OLgAJf1O0HDHYmPuZepjFoOjrGM9J5
sUz/2J+kMa2SjalMw2iYncj57dHN3LsQAfmzSF/Rk1sjRvbh/pdmvmGE61+l1Bwa
sa3SIGRW6wj6rIX65FQqBOFU3ctRgl2M3eZ+6LayWxXLrZCvN1sMVQmX2yKMG9Tr
SVuvTkBd1+ZtgW5gxITgQIbOpg24cTcWDWn16WC5wlh+ITxNIcS4DhBrTAdmOYln
78+K8bXeS38InlLQvxXau4AKYOAk3Cz1ODlBtpwkh92eO0jX4ofn03rG1+LLoRAV
aKqaeCN0nZxirGff0tiMBceRMODVkTkCU/NzVRKiAmalKNecBGvN6jFQutYxPTdV
X8zppHTXvpyoQMJYxTzQkU1Hnp4yskyHYTvgWvuoOuHjg1kEQI1JpOeqEtftqRfy
FVXJaIu29DDWU447aciC5BSwbmtmJWsbgkz7E+QYvmI+TG95W68OOfztvKJY9MqZ
7LDweBaUPsDXJ6jx0BtHzmu9oWEF8JtixJRDsMf7oq3aAihYRaxxCWN6uDKhVloZ
S4Dm5s6BOFTEX6DbzDKXHn6EEGvyH22a/vu990AHyWj2GAUgqLOq8XGdBb/bo4bA
01QRncCWStQh1ni3fBYh03fMdacTKi30KCqV0RWPYd3ZGa5D42YCMTrywKPFoPLq
7F+0Z/ruQrF6iA9xLU9FmDceGXOan1qJlQiDe2rGUoN3Mt4PDGrpCvy6mzcZ0NVt
ZDOzAfF+7JKuFggBaIQ9/8/4JDpWPm26S+NxqTv6yi/t5C+JcCNhK+52uug3/IjH
Wcr8HmlYItya4S0XTuweBR4mmOz6qiGftwE+nYhRyhwVXVZBSPtJqwM2Vqa9XbIl
FjlUTNHVXVtX51tB7VhYQLk3syiQRhNLvOytKjBbbQybUZHi1HOFGCQNSRuCrw1T
1aAs0hXOSbCndzMUICc+lDnttktDIjG+B5urq6a3MHqblO1Lnkux/aiNYuwzytYz
sykjzVH7M+46XG9VN2AUeOUl/4xBLGGACh20lTEPY2a8jF2XF+CE7COHzDyuauoK
z8+brGhdkEif/ivnxA2ARx0Bg+0VnOwQMngAxYNfLPP3EqOiMDnhbgfFDSKKkrvx
rT+ACCHVVGW19TFLN42O01QNiDAVsvc7G2BbgDIj8WP93seiNZMjch7FZqZmQfJR
36kKyDpcvmXO5W1OfapI6URq62pQsbjGN7ct96T6VjPui7VyaYrpC1JczZQkiyzR
1Cu3E1dClRVF9lHkBsSJQUph2igtcKTz2otAZjzwfCr48X4V/HEkgP9stC2kpt2q
OKBROQ2VtnqArm7ZoqSR+nLmPFKrEHINbh+c2uBOorkfCUDih60vvwGu/7Pc/oxW
EE5JOGhL2STvpJwEjuMvYf/8ui4nLCIzp1D915WCu3KIaL6LHPN/EGrfKMFBU1Xv
Jr2CNTbl3SBFGjR9pIc4EUUVgyE30o4U0A6DY3IzJY4C2MNtS4uPJPof/jR63SnU
AHvlFlRLtL9k+oh8dazeXFf9B5hyHijK8EVxiLJY6eZ07CdFljy3WII8GQUsG3+G
zsjmzth0dXwvu+9LzxrscxEmnPHQA3mz1LsKsDRd2rYMnLf3EFrb9qURi9PLIFI/
CnACHt8IAuObNEjIH/0K/eu+qeHWkD4tx4INs8mffXztHlfUxmv3X6VWGoWNwMda
EMppLElwN6QYYm2J17ZSo0OiSDi//jCtbt8Sb8haYRE+iz7zyTqtuUhizZxNFbto
ZpmYaZaH4sbE8RbWivh0cvWXd4SanGZ+phcpQY4JnOEbaqICLCb8d0pG6/je9TZc
X/5GlfzJzMeemK1E6fF0OTOa6lPOtTMeR2Mg9N9600OO46cBWCk39mxhOHP1jY9J
RS9OJQ3bLfqWAiNbqHSpCDozM9whlAkPCXs2wjZMmH1r3fiAQR0wxoFAOaDQ37v+
Fm8UmHkj4m/zutxD277nCXU0HDnuLE6OY2NHZGp/SdGzPoM74twjNMxOuwIKGtAv
/KW2BtED8AmJ+EVHzPeW1fttFC2CE2VdZ1twjY3RsF/NRKzf492DFpEwt78YNFU3
9ZVfrUK+NTz63K0mcUqzaR1fYSKtZ7NH1J5lPCkWRCtbo8iNkckrIbLvAHohdxGx
d/228uwe8cpRAy9oRr3nhkP0gW8s4y6XqJlGJQOVMdXZzxqMJneXKXVlmQueP1T+
D3eTsnBMaqWE/kYmuZM2ZAhBZmCHKxAutnU91hG00U3H5+sdiS1tpu3PQSy6Vrv0
Nr1HS/zD5l03ujDgy7mDp4XmpbtPFvMsgmu1QFU0QOzVSCtqkLl+fOjIc+V66hGh
0QsBe8cTfxiekTO5EeHv8tH0PJ4DSHs1ACeEK7OqJTlZ+DL8NGDuMQcM9Slukjwg
afnfgZLC/R3eD0iu2J7HMF1UUvTdHLSOW3KR8RogcX2jCH+LnWIsPkYl6zS+cTrB
sqHSwVtEcnNIfd3bRG9ciPs9cCMxGW60miokE7W9ymkadfzW5eL6WwSaETR9lzbE
sDo65WXVEYEu5FLcoKz9urNNhl4YwP6RSzVMncHdkwQwhB4gFiqbZlVmEf4B6b1T
0zrYuU1gcKUnspc5Ia6kKiKEmZuCqR4b0E2xgImbJDz3ADrk4gb+jZzdDQvJlimP
yl86WSFIo6b0szeXJyUyjqIJ2gsUGRp/ihpF57BwqJk0Am0Eq/5LgMmIoINgddMa
NwY5k5soH+gAsp71hybsVeNGAhbi95Cq9hSHBDHAlaD+SFmShMMP60cqwvwYcXzh
6tQcmX5mmHfrok1Gw3fp84Bsr0v2G/wZ7dhMRPK92+ZpvQB7iMooil46wyLKWvGe
RgZ6Ae0xmhYBdBi8quFZm1+GGHmaDj+4Z7L0l+ulh/X61f9PhJqETqtoZ+LBspMe
wdHwzp5wjbuSzqszf2ClvioWGoxzAmUu9+07IZkTXxNNRhNiPb0d1mDO2mLQsDsu
ulVgFfq7mX/qhpnHLBRokA0dHTmo85npYRPt8QltjKz2P+gLjYT9oTf/48YAoO7j
J+9momqwOPqvOAfidg68IFHW5wHaiBwAvkHRg9P74BdM1xIRoGnp1kQsLoE0g6xd
MJs0Ldg6WQNiWBtoydp2Spk7Dx2o6qO1CgV3Z/iWNbTv2NebJST2vYgum1+MZ7MP
c4OjuTPdJqN8mHqC5L6mylxkY68xwdmTzieCrcKPYN+RVYA0YIM64bHeFjF6pgJX
7qNHpyhDuAr/y/owYwSI1gjOjL0gGdtOIw/u16rRe1NhFQjsCxOg84btpctMvokS
zi1z6YyANKOrhixTxhXGjRioMNum8NQPe6SAJB6MhaYvK9lorq+M2Grla/BF7Vgn
YBW4vZEfwUpA4m48A3AYTZi+KptpjtwtmlUe8IGXbsjL8RgdRj+fuI7wLbRtvBTR
KP/71/5lBUs1tWn4Q18LovNdopnsISB2WjDMRwxNvDhbM9sdRmM5VgtUgmHePsbL
chbhLSdFYT1Y59prxN20ukZq28lLmGZ9d6UkrzxFrKAFyj4df2zznnc/bAEnzueY
qkL3hXxfZJ00NkbolcPDrWJeAjd2+3rhasP3tyyKMnFdGZszXINM7fGo5Zhe3P/E
SUFQJK8mWjKM7NIekHWeHHdjSHU9abLyjnQ9lN3wsfILiw/p5SImMOvrzEaueLIj
y/Lr+ArwQhgIigXS8mcZzOLNjo06IC9ho+VtIoXpLvfuunImjzEExS5CHNXAHQ7B
RwPXt39SFqUmLDywk5yd8W7wrxYEwxf3xXN3i8CGcmEKPfTrJFTtJ0+yDxd/SNb4
GcqzuEfeE4lFDrlqRXAqYiW1Tcc1ExpvBR+vWCMKnRoWRvCzbUe04VLRnlE6/y/n
lZNuJdBqrI6g46QN3jIwGcVCqX5xtKFrbGckR42VNuW5Ehdwgx1XTrtTONP75+Pm
k5DGnuxIu1wAv7ZrhEerBcSINNHPZBfDc0a9sa82UgqBne85Ty1Gp4y+TmCFKg7J
vQqLwGCIkYk7eYo9VLD0ACsOxaRr8v3JRdmfC6CUT8wx2SfOnMhfmPdOem9Hl4OF
e8gPbqh7z62EpSrN40YFEzt+ESmxlXhBQjA3wx5KbMks851AaJ5zx1546uMKe9Kt
UwiwXvbx87BdpZYifap/um/kAaiAqT8IkmaC3/YZRVKg7+9ezPmWtIZdqJ0seAIB
GFDLxBmy0ArT4rIPBNrAP4vHuVe3ULJq4d6JZAi9SyTr9eedRBmZFoaEdPsky8Cy
gIaBk5Ukl0vxIGLsa0fn6aQh5YrsIGNMvq8ibXK/pmybXvt4NBq3noI/i4swrg8O
dS5HJridvneNw3sY5DF4DSzhDXIq0/wxnbFEiMQy0AyGCM9oR760oy2Y+4PKkR2L
1QOLbbEzJ+nBEqtv+HBSNsAaCrNn0v7IlWjeNRL6QTZvfEDr2dSPSzToEQUywXxG
bvHzey0e6JPaHSdQdb0CJmKzT3wg0nZykHelGJKqMmN9NI2QukGwGPaBFFX2ebrK
74iHOp5664tegpz7y8c56eg1diDs93ox6cvbHelsbO/9d2UzRuaJEhTzmQaijju6
zPyD0m/X9kDqoAF1QpBkcE/fsrkZZ+mtM9rHdGRYngYcbFruNQZ+u108hNry6Yb5
++92dkZ+o2exAY+OscYhGJdsSZmPr5LXobO0wdD3yC97pgW2bXLfDfktravFRIZ/
UkzoP3MyLdlDw21h8AR7QVLazbdQ7f3MLM0eCQEjafGrR5H3NQDLogeUqmDsviKj
S/P1A8ZrogoByozJ+4bRh8FqZFzH1OzlYhZcMuOPrTNRdMsKB2fIJ2JbMA3IlJ4i
+uNXmy8fwKGeew9qoHJBdczpnrBhZo6h8lLPPqOL3Kl8U9Wpd8+QHzM2l3+rVYHZ
pfCuIK9DEFmE+ycKveQHat9dmeSiVkBjcVrIYu8Cf2ddjwQQCR8Jq+i1o0G0damz
xZNaTlgvtn4yIpnqdikSgB7spNLf99kFPF1ThB1+bwGrvIVJI3UJn2zAxFrb+Pso
ExvOXv8btObIxFnW1uRITc/Q8gPxKcRo0yqd3g5TbeMrXxUJojckTkMCUqOf3R6f
BTLNm7cZbSTZZHB/q5ePPOSkGu0X0pxnYPfDUxVfeGd1/HN2SHXRaRcQa0BYW6ua
jmHSV3QKY4N+gD4n2yaNPKylgr7uRV3j5TIjFthS5Z5ZDvveULLV4c9QoTMV/xY1
2MZDh3xeNGC5hFHWw4/dWcXtRdSeIp5u60ng0/44u1FCnwTKZ2DXPRUpBXhtjPvl
/aovhwInT9TaxEJYjZN9K9E27OWJASvEz5k6gjvzEQpX1XPPnGce9Pn5O9fRN5QC
Aw2twKKqfyvJwE2A8pPetGS7UlAPhvmy1+gSlmG9mIG2Bzpef8v6JkzUTInl6dNS
sDZF3D4/hEkRdbAkTkV0jk3cyVrd4ijCZLavIIgW/0vEqSuRwC1yJgGCEpygvp0w
Ptt5JZxSeIos5lKhrQhfEMOH8IPz5440DVOHZFHjSkw+pk8cT39qBm601UPUSt7m
9u2J1EdTiz6i99i3YJBx967RY+Tfe4+W/d317nsdcl5HWIsppG93JhH/t9tL4pfl
9eBcoBpYefLSBWqkl99pDAZToEwabCAPl7ay1nUIJep//PKzQjja4NOC2pq6/Zaz
ZyHrmeGtJq7NYnXQlAPBZo7Af5h5nMdzZF97Wsu5B9kFod9PN+NUnmiwF2vHL3/3
q9gyKrJW7IjDMT3ozqZaOXoRrz/Q1eJgkxfArPqsAL2qIt5Yu53467gvvwVYXzKP
FR/zfoCV1i6MD0nVk5aoKWkTllFmqXJfFhWy7irfmyRLSj8373TDCn0vvG74Onf7
hbWDMYGgo6qeDFINxZHrU/oaH0yu7bEi1rHfpW8aFiLABu/U2IyhckMpFGM9Lcx+
PR9MjNmSrl5xjPnCyQ1I5aGNbPs+FtnPDbclnAk8Qv/d5dEUzMhgSCYeRpxDBpsj
Pcr/ntmRW9mBoUaU4SSLvsp3HVJ5UX8ustFEhiDypzJiArcRHNcsPJ4452eEc+aW
h4EfpkAZEqa2ZYw6/L6U2GOplX2UUHBwJqAvINSSs/S4Xfh3bMSoxkb8E5Ro5ZSd
8ZRRINuEhFeOZaws06dVK7ui1OB6fkJX6JsfJTp3cjQXeYC+goUoU4JNOkLbeoDO
wbOGGTK7XY54UqN618OpkPmwBAgcnnbE2dfT1C+DhK1Ns+7s+67edspCWFspYVDT
a+Ex64kspOV7HYwUPvW27Ijwm5L/Zllep3Tbe5Cc5qmoNvYVCNEBM1gVVBTQJwtZ
4qmTI3y8M943k3/FSKwz1K9NeKhe4l8uqUdfKAjzD5FS1aWse+UG6NEM6F4xG2Aj
riTVZOh89aY5yLPpSEy/Rw7YOZcgx1Hz3aXW2rWFNO6pFSj4Sp/znYF7oNdBthUL
yYJChf6MAiP+Z97D/EM/+/w1IHqutQ41loaVo0J6TomJBW6UftxiyeMTnxj3porW
rtdvBQ6UEznag+1PXTdJeMTJo26pnFb9WJq/KpkQfVP0gEK85+IKI7xZDk335u6p
RdtFg60zdV0GFgGeShkelXdryAELrrDhOUDS/nYBZytkB+xKbPaFVQmlgNPqDuZ6
uZqCKG5pvUj/Y4gWzEVqQiBDv827rxJ0Z8PqQ2rgil13/PIwv6tP4Px6lXtAUaV+
tuJpD5qv+t1GcKh3toOzQ96+2D7LlWZ5Ase+PO7I41PrzdzoM2fx38JgriHcbXFJ
4qdPdKfJWD9ZKZ0aQYTJ1tbh9Ku/YXXEFLxPEuCqxqHbDyMMAjQECcTrwVb2ZjWw
UXN7j3dUmh0eGeCMs+prfvtMO+3m4a7WJPlpog9avF+bkNOINDcQqx5wVY8cxz+r
iNASfehKXFDpLm/1WgwmQgho1u/YyNp/kkIrENKB8rJRccFowxcyx6VAVCY8xlVO
H6F89WGFZIpjMznr+QCWZC02xJf9q8NEFI7JZQyYXO1AbObf23UEfSv0K5D2vUY6
Fvp+RTmrQaI/zsfbXzELPBuJeuiNNGE4tk8jjw3i5aRa02PjdtdUMS7g0jeFzLVp
qqEEMx8IbUD9/K0b79LasrfeI7LzbRKq5CeMaixII2LXNoH0AlGia4HXgWoIcuqE
OjQlT24yfI+6I6Ng8r+WAd1H+9SZg+3XMJmaF3QfA66YdyyTjTWYCUFXb3cZAWdP
x8BMCJ/Ik/FZhoRC4f1mjC4dIYjpM4xjTpVyRY5oXxYKX0zKgwOPEU7YWB4aIqqQ
0oikrf7VozTZMkmw9Yyk7RYVI8l8eWHnMpWX49tEJHaPf4e6Og4ctG0okyPdohl/
wng2Uz2IRxcNKYpsemuW/KX0v6csINTnPsxcczRntHFKCvQxcIGB9pvvdEr+DztU
Ji4rJkk5YYDB0IJQxrPvZs75lie86Jf+R9xNxGZvIttfBwgW0HFJ1K1SXVGnhSan
71PAbgNz+f1pCFxMD+WaNsdiEPRWlwQKz8BLODr6PAQ+VDFHkIXUd5OxIsTxR/z/
QiJssFCWxxtW0KsxGJWYsHkdFAul3xX5uvIXnYYbHw7D5REoxmnVjsNE0RwTIDQa
+PXMKNce+sXRBSE5wkRSFdEXM8zNsSEdB8VQmFZUuO4tr38AqdPvzquY3yVSOmf8
BX3LTtMThkMvfQtGRh7jD1WvJ5b+yiOUdDIUwUCGbooFPbqleJuJBZ2Hxq6i2jRW
fcaYG+iY/lh7otmQRAUtQAd72cUJH7C4BtiUiV2jwkL+rD4oTeqI//ddXz94VYeL
rkUonLMDaRieHQA5oilyHRRXQ2oCHUJgCCu/E/Z4ZxbHI097jTU+ilo8jFTGUNfN
pftWsFJ4eU6JsCi0+SjfdfHAY3y/9Bz5zF86LqNDNU2dXhpHP0lF7mKsSvpwy0lU
ih3y0FEYYkBQRpH3jteKZe4xDoHzrHgQV9EuPdehyqjR166OAzXomut/jeM4sbKv
fCTGB4pzDuRcXnCkD2lkxlv+KwUK7Ye7IEj58VJqsryU4zenTxgh9n7fz8BevXKc
OgWw/FgvPCnAp5N0YWxVQ9n+8XjwUoq7g1UogO+CVNUd4Uj+VZj8ED1ymQIPlX1z
9Qbijrb/LsBc+H/sj+09SDJPSOA8OQMUnaoGcNsXIfHEU5FXMIbxKJcGckI+e/Wa
hcgEwZG0BhBRFaLI+zo5BAmba2LSz5h3YkgH+kwL28cnIwDxrsqOpjnUUddLj4I0
MNdqKo7qEbE3Mr1q17yYdfOY7Ay5sQhd/RBmNzKsIAwV8G5wd6Y8Gm68s7UVXuER
1/zJuq86WeA4GrulWCpyQ7Kq5XYK8p2dx2c/GRTKteiIhk5oLPS/Y8Qg9OeAtuL4
NeWLsBepewHKQop7fqiVcEkDoAgirn1cJZbMgWCCYHcngKbalxhnIX7nL+AAciLs
XcBgi1QzmpTFaGobZgsbUIhodB0GPeXgXh/mm+lncfjUmsI83Jer668ILe1McxC8
idFat8wlxyER7+EXi3YF+n3j0fU7i/KHbZUcprW1EZJlQRS0MGTpImPEJXyYgZZp
ZZ8XmTZM3pawhLyFVqt7fkHYTMCMFZTcQAK1VlE5I2pFK3kYUurYIzdM4VYps8Sx
r+IXjCXMcRopHDND/sVQmWr9dp4B4fcyYsb7/8zkrtVywmNSA7E7CI1tNy687kul
+UadJ+6Q07Hb4aQnyii2MXn9oxkRFMxxpya3te0xiDEcyp6uQhN8MApnVl9n6faC
LMiAOo3MBnVNe9aN25brnilbHmfaFj77f66KNG31i6ISsfZ32KZNWjlbmx0YogUe
9ow8Vd5l94Cmez1Wdcxm1klpgZHmsSDrKkct0eQpjIDSOW8V4dMycyOMaf/WHDLu
udV/BteJDczttTaznQYqcW1L/rdxt+7PR7AvL+gQnFXfbbNZs6ho2teucym/rVuY
j5XSw6+0tLFaMJGZWssEyQHNlrvlrVmUw3smAPlmOGzLrecg026VbCDiCdEPssLd
XW1ML20MRfe8nJRbNqrYqTvdx8cTpQuUnzjR3b2XnkXwYJbg281cHNBPz3wcsjig
Fu4jiz7UH6IUOIhXNjx0ErtHoHPms70od3hBeNCYQqHSl/0YSLrILdF4gY7r/J1+
lrjCGA/5A/MxhT6UOqKsoW4X+Czr1m6Ei+Mc4y4sXBJRA0UlzRfyPADfhC9QSOnF
ICrQ1/vjomjNnDl491QNSkYATQam1Rx3godAGq/A/tItjst+GGbn2AApj/PbNF8V
RhAVVj6SK/nfYyPiWOBj5J64ibkx1JWSWBoBkNsaVSkXMcuGJkLN+ewNyr61URwT
zUFfJqu1R1kTxYgQMiIVrkU4a1kT51/71DRg7UQ0EQABqNW2SCPDrAERm1CjTUaS
Z8DQDZENC2SJYVPCY/ypdEb3HQfIwiiHT80gAbybjF7JerHZpVbxyLv/HKGtBMxV
7i/xr0ONk2A5R/ut/d3jkfhCCfTuVvZZE9TboDEnlNSUv/fJ0QYwXPRDhyixU84X
Lkym6JyM4weF41grGuzJaFD9RCCZ+K2tE34QGCXFnlNFPL5x1oywEi0JRu+xXlOz
WBGkRfm9IT51FYtfo7pZd5OfELv5ngN8UDxnFrzDOKC38dAes+1FEop25vlecIL2
m7iBJ0UoegzuOGk3l5R4YkX7C1zSi//rxkfVtZLe89ghF7K0BcH5XPyxr+nef5Xm
dC3wmFbmZMh1TXJJvqWr74ySBVkyDURTe163dPkIQnybY3Ow9hO5PAgQaMAqINpp
5YYDa+2M18nhTkO6BMgQc52Cg/J9F5f6CRDR7bC6tpHzZWP08Z0N6dGTtUk4Vjrw
EiJtTz/bTkNeMfePvUQSiPfnDGyyZks151bs+mdZOt33wlQrH5baMrjiw70iG04n
I+qcLRl1HWRZ/z1X1hb45+lyquuiBbXHJcHW5ZkLP/Cr1WoPfMD9Vpp1Z9A71JwY
OPQgVG3Z3xtKid7/bH0boPHedZwAw39ZJ9h3FgjwrMuJl3E6WGxaRq+Rn84hrbk9
TZ3UGukGDgLUkiqkR+oaWA2C+PaE5v2I0V29FzratZ34myxzveUSv7DTmHgqy+fD
eZjnJudNiG475YxtzPyhPWUCp+QCSYRt/gVi1B4UpGM0/t1DCRy3SwaQ4xKDg6xE
e+gxUEwPHflv8MDWJ5PYBeYD0PQhDPGIujAZkZHLtgd2CfL5fL9X1mMDQruKFKdz
1Y8ZmZ0QpwreVzOnvps1a4bO9kIxOoOlat2qtb/iVQUXdmQcjPXaa6LOKqywhM2D
0L6vspch6I3SwgmpItY3AYTcBIa0XTF0kB8Wi7Yqr2swDC2FzhJWDYIUTK+HmGin
GSlL05Bmr7dM/rfSojkxKcMAuXPJ3Wn6YrKFXqyg4O8Pz8ZMQZ4VgMc3We2vDNCX
tnL3tp54AzsJReYA77C02LJHDS36WjvOCwO0XOe9U4TinYndyvvNnXQ090g+qtpi
91NoUeK+6uK5fOYY7lHp09THgMkfvuEcLuq7U5DLw9HXA6CnsPOl1b7uBdhNnjCs
xqabneRr92UF5tRPFTs0bBSQU/vbEp6341uRjkjVOsXzyqLzpeZfwjkXFm7KsWU1
bk9qjNbjzuyZTLfRf6W93VPmXh+WjxuxY2mhVDhlHLCZqNLZFdh/YKZ1mJnCGPEH
JGXyzK/gZ4l/C6gfTtE9q75QgxH6KD1BY6QBjCvaaCQtbS5zd2bZ/tsIVInX0fVm
njW0yFVho6f4xpcm0dj+F1IcmNUXz6Xgy7A9BpIn6OwE3AVfmKjUAQ4Qb4WwImQY
SZ6+goLlw/xcnbqUW7nCjiFiBrWg9werdBCQnCwS695Bezb+99P/FobP3d4URWOn
s2Z/tUTLpTlMNAUOyO9fbWbxLnu/GAJkLqxZvJnGk/7MKFJTOHdt9LUQHyOiRcRy
ihdMx82WLsFiW0AdqGrvZuBZE/1uTxdLTk3cozEdbPUTfONqckCsT8pbV/VM4nML
ovgorguh3wto0PJ4Zp7vGDEx+DtDwtT1tBMni2bxOQVXGzsN/APjqNniBihzzGos
yIlHVSCn24h8zGnLET+JxI110jcQPnuF00OGvsQ/s5o3XpcCCyaSEEnXddHdFykk
3tr2RwA8uMdFftu1Js2e+xaEfyA5p8gFLgMJEeOPLjlgSaOFLBlYKvez6P6KYi5u
cw/bL6y4h2KrtK4Defsv0qGtdD02bk8syHis2866zd8COKKoU9MIdJGKFU/1iLXH
qrxsZ3iXN+0SIFJ8Sa/bj4aohHv1ONCCjS0PrK6HvJDPnoqxlQIPRsUwymbWmaCA
PeESn6Ek4rkGppv5RZH17Hy53hTVNT/Od93lMWIA503irKlN75ZOnacJmShbkZ7A
Lrjso1Qj6rtnteIDnwgiK4kaSUbCdh/H5HnuAU+A+TkypZSnmMj7px0y4nnps147
GpJ8YZkdVQ1QJ9hHKxeHf5x+rZSKyyMvIjiJeB5UCCaASLJZ+KiHq2NkSvwqZcWg
xgDhkiYzIZrW2dxCv+oCUqiBhQkVXMZhvpgbJFZ2hpPdT9vKTYAIon0li6yA8gFB
P4StiF6B9kpZdyg/NAoeEgC08vb13ddotBxhwmGziDuKL91+M8oVB27HV9QOWmOx
aGBw9hS0IfD4mti1um+5+0VvxB6pL8BEmsIoYKTvxNO29EuY6ao3EatfDHCQATdI
iobNkX+IZqK1vtjmHrwKXBImVMgkjj3R4x0mmJxx9wmY9+qSW0H3V8bL/P4c4cbp
LpzmDO57xY2XiUKO2ys8/UUx+w7+Gqa+f2jfez/UpNxOyuqcFSySb9QAo129SFAm
xnMZ7S6chSigJtzRqIABySRZQ1HLU5FF6H8PtXr9bWQ1vZcd9D9wUwz5RwlwlmxY
hXCuU06gDfMpzLy3aASECga7Kop/8Lfhtpl7xCRQFUC2/voKW27fx1ilBxHyfBfY
gTMhSe6fZYcP9uKfG/2d1qhVtH9UJn+jJech8lmUiwHGpTvZBS+14wRxuGWrUnQG
I9UzfdHE/TFqgSaYEEmnWpuRlzlRwWXVsqQ39CrUxmE52Nbsy1AhpUrxdNV511ta
R9uWmUFPVXleN4gpnv0cJpl6VPBsQZ2zu+glqiBMHG70AUeuj/JbHYbP7PH0XZy7
UPL3bjdexYpJDqjcwpvPK6foVOAeaOkS9iiRj/yC5N++hFnzzvBdrnUz3Fs3XhrJ
/gdRi7nc7LXeAUGSMKjz9H96AxsyPk55QtcBD0yDVeR9TXdfhB+f4+MyEwyWfky9
EUfuz9itAEDd/iMU1TKC+8ZWWJa9C6zVdJv6jl832F0uMTYsD5dcWnZFfZYiSyxV
vU8/vB3IS3Oc+DR3lgttyjcdPn5K6PxGsaU3/yd5mldukJE4cOHM3JEfxeR2VTLs
jnIv4it+JNf7ykw1g9fT0c74IC/dfUMshDRR36UGTz/BJWiOLHqMQGVIGAd/xCsL
/MaaSRz8/fABsb7S1u9fyBKFpegmOUiKKY56RKIcZemM9UvQ2HCcdiiK179Uhe8a
7gUIE8I9LKPl+A0rv0vfW5evc01gYkJR1hlurEm6FtIGFocpiYM6qWh6VNw+Rj7t
HonKtmuQERiKDND5Q2NsXx+lYYGTng9PJFc34da91J627eo2BsXI7oaLiFiGTW3u
MNo1AERWzGYug0Jl8fMbsG90ljAYnRHkTtxfbwNCiK3cWQQwjqu7GxPVLb/o1Y0O
qelFPBH6KeR9AQqklu+IQMuq/7Am1NIkYM+UhnDdLZKpxLw4FPQrVTbLjGyz5hFw
YNVqZAhB7Kb2DtlO0JnHHBD9QURMDfF+Wzmp2wioQwa49qqLn8d5w5feMeTDvdox
QNdDL1OSpSHJPtLTDTpUn/Ry/eARLM7IBsIHHGj25tkfJ7ESAODSpTIi9ZMBlx7H
O5T196xaEY1UVI3vxVAvDiFqV2bgkGIMWI7lB7CQyys5DvNwJuqQ4LSK9HftzA7i
pno+NbfYwsHKxssxOVFmgbuGtT7b9dyfDudgh+oLP47S9KZfsPoPUZbL3lgHYH9H
Dl43Nbp7LASR7y03ypfzYYbkif7JpvcyQ1esGe35QAc4Jx9Wjm5ezWLaLZdg3rwy
G0x0m5ktASU/JCEu7YP1al60ZEK6AtB4VC+2yN6h+9dGtcC9RS20hA5kGok5wREx
rAMw8Mw+/wTDKmNj6zTk2S717KBDfjofKyv2bU9q6/hj8w9oARJi2nLrBqo2prmB
aNTQtDZmaViCG4J+oAVP6MdZW8VQlv2xricYR0lWsGYAxygdQ9XILt7q5iEXkNF0
0lSB2C0mLVnnI/eljUKdt4P1xGaV83/Hp7t/HLcYD/OEVjP4s4iU9NUrzni9sHH8
q4erw/W92yV+G3f9ElDaQYBdEYWzGjpbYcXK8nvQKsRxvf/3JuKt3wjncLD23Lg6
Flny37UHP78gKETInjrUa5RRvO+Bcig76jJDtZx23H2yfu0D90qANPPGbwenZ4+w
45PZEC2WxSK7HQ8Zd7bkERHn/NH0YTdsMc4fV1R2+eqTK/oFNHmrQecw6XYo1IJT
tuw5TlZh8LNPkKibBKbmONHTj+8obj9KoHqxtRto6cFc+CMvAsLWu1Oiax6yiqKI
OtuMzCrI3KX0MBZm84pyaiV4AUla8BicjJaIpbn5/o3ayX0s94jjpsiNGOIY9eu2
Oql8u65GRtAM6SecWl6ax3CS/kx60rDl4giDbTCugpx5maVwrcRL2ZGHL5S7W+aF
YVaThStXU7a/EK6iZWqgLOrCvz7piAzmfkEhrVIVfWZWMv0QKUyX1qiAoMTSRo0I
OfubUntaWyPHrBjDMiQnSzO//QcTC4DBinmFxzwTxgiAeHrxt+oYC1oJbkJ0J7h7
W/kA7zKZMtp0evYDelAV+RPu2vIMk5nGLbJkakosUiHDhy0ErJk8QAjqCq/hYNTb
cbOb8sZ0ZujX2HJUglUTJguUgHKcGPeVsMGH0keOdXmV0nwdmtoCb0lsjyrgy6j0
br/uoIc8W8Yj8IDm05eE9X8OXgagO1uf+dbYj3EzDirSmbIfKpE26T9V7BY6vfy0
TsUZMs/x3Xg+S8TVHq1Lviohy5QUXbrC7nSfUIe66EVu1XUhVl39/eOo9Qk7fr1T
1Pm+yjFrgx+LnNmN0uGpwryzRfvwotlC+V7YXK4gC8GZx5cqGQyLcbEXp2JIYTNs
HmmYM20G8A9ZHIuXFHjFxrUG7yLXoalbylajslXrEZxOReY+IdFRgdgdwysViJk8
UmsWpFYm/JOaA6634oulpchyFe9FmuTtIgYK1ZV1X+idHmyScm+MLzscdI9fnPX1
oLv+/0+Ola2Zn8SwQmqSxcbBm/AjiBQKl+fr/teImoTj9cSSGpJYd+YiuPNgAEmS
9gea/D+t9I3xMNXLu+AZNuNRULjEW8c6ahH+lcb57vZkKSBL70fkOsmfAlUSdY/b
NdnIcZVF2kGdpxU2+qP5aLA9veF7s9ur3FFI+umtZBPGLCqxHFduI8j36TkVtxif
O5aXypxZlMTlmWlhc/F5Ur9YsNdOJ4H4y6HWV+HDC2iRP6yoY6ZzQHRSfc6mo5Hd
CxAv8H8oZOkTTLKJQ9bKR+WxRRyEk0qPRIZefGowfTpHuUfTgcFNFbnmZZCTGQK3
/f5gYlpdPuX9zGgnOiTDWq0IVvUm50Oi/G+bi7MfUec9d4ZrrMlYovhbpuPdbUkv
rAxpoLhPvhhT07knwEnc8amUBbKDX7TOESzcUeORALaLENrU7uWgHq6NbtuoK4NA
kZCh3lad/L3VZjPhQUSew2sxbVJC/vvRfPWS53zYQ9LHPMlEl/XIXbs7Jakd1Dum
bV9u8vpPA0AT1xmi/S8xd20LQADLaFor6e+dQ7J4LHMxcpkHU0MOQ4pc/1jKRK8X
urSDF1AQgIID4STMXmvtyIGdNz3Nar3t6UPPdXS/4ufEiTiRAIQZog9rkW1Hlks4
3HbyCEyb9kQ6d9tnP7l4iLeWn67jzsP5VQOgfvCRx/8QDWo01ZFmiAKaG+Ny8AB2
hbMuTvAbnKS27qkAMO5w4StU5IutfXztjqt34Qc6yehp3qqZL4NnUiop5xNv2zTI
gXEyVpdV/ljfuQoWheR6+3ottXGK+jmeebUpzZWbMic4m2unqmxpW8sAPobCenMv
i9q2DIoa3BCkvihMbDTlU2LdkrXVrxTgKIo0E11kzw+Z2c2OP/xDCvJeAmJSC7CL
`protect end_protected