`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 45040 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
0ivLeOT4zMq5S+D+IkEISP6ghVrxgZ2wRM7mZFGMs28OKNzh8wzSofPquIRF7Z3e
6jofza2dGmf4j0CDWIKkcpDb7YdlRCYjLml2mpuZNFOI655tEIn4DNhIO82rylHE
9bhM2VzxWC3Fu/59ojXYezeI2XQJwUjAI8/6YBXef3TPCswzpebU3obMG8/taBUt
DsGKBHcRQXcT80FYk7u3+RiVbswviaSQQE4nhKNVA8dsUN4vOCAcYa7C6qkz+XYv
YFcLtt5AjyYpWUdUCPdGnOb8kcKDt7u6WVhuuXebNLwoR7ozydQWsg3Oxw3U+e8d
pBAXDS9YPTg2QlMx8cLMupGfs7RN+3oBA9jXXSmgYmGkupURw47edN1eKU3RHQw6
iOeFtXygvKNdiLYP+7dpbSJsZn+AwqhgAirrTwviTIJuozruXKpM6wYnCvp9pt05
Vsk5aKR+lvuYv3GJPSPvjq3DD5zICgo6680IT6hcLjIdR4Ws8Y7qsbR0+x9RT8FY
nxkHi/jJFEnYWtqZNQitwpmGkbQL0MFecGefLfFd4vSEDLY1X9MhrlBV0FN83Jjq
7smY0szf4j9vAPwEMHprT5+5hcaRSXQQnmGGlor6sClgLvlSnpOJX5wriJV/5Fva
asTcm5BFBHo8rPCNSoaaCjGIzB7emHzHpaMWt6qnUDFsYHH7/84r6JBWDgvSEE9i
ykn7GiJu5W+x8MAWJJULE7xFNMtOK9+QNTG0CoRFijhK2NwINRoQzhp1rgjOENZn
Dwb72pifAqotNmEDYJWBywokzQ0q/+B8dDDW534DFybCBdMurfR8AieC3rvJxzsH
FcfGv8cc13rcP3nrw2MrZ9awrkZ4ukeT9+eWEp3x/iCiEPKxkcHxw1btR12K8Nf1
rvBlJyY7+/HbWhiXHdcW+oDDuMDJ9zrB9UxdDtR1NXuQJGPtwxTh2tjsg4vxJq/G
VSzYiyIhACIg3cCskmkyUnCaUe35KcZIxSZ+7oLEzR+iKALuwQCTD6E9C9dU7QR3
AMlDuVdku7c/rGbfAQ1oZQgcSOrkwoT00ZZTLOe0lk4WmPD5DlwAjL+1IKco8UYL
jcVivMFJU/2tiumPOwKyV7p1J0c9PtYstxLtxo8plhPs5CVHlGycaBhjSkxvvIfC
0svdWWt3SioR23RQf/HZ/QzI6Bny8AhIH5UOHjpgK0WPl1Qm/iBz7sZPlDtitnDd
yb6eGvgag7+C5aRC3z+35/EErOzd3rFjXSWJkzv4DUiIbdqxyN8KFfNn45J4QAOX
NKVaHE6PRjHlKrK3Ppya8FbFrER9lOMvJko0Tw2W7LhOtC+bij9aqEW6feF6ThRZ
8mg/CrIBlAK8rgAMOuj23v3C5EfLGQ32kc1Kn3RqXpcSSgnMHGYH4bOAUyWWtHbo
eXqnaHT5t+MgCUN9osQPeAwTHaC7mHxNuOA1KiZmnsWxkIC/SdgSxNGM67DwEMVZ
3EEIlQUBgP/TtfJ+qRtiQWZ3fNSavXH9nvteGcP9qYANZB3n36gMMUxEUU13YT+4
D2TW9NSp1b544KSG5fKO00irK30r1AyNveepOFNraZ36JuUVVWDNOaovDZol2nti
HAcQ9kHuVElBMiCGlCOC7FgIn8B/koCNfhO1iw+XUJltzfG2u+nT0jJrGR2WH/5x
LMSUEo5FzeuYAxi+SO0ZoWRDCukmJdrSf75mJjwV6EPuDIg8VTqSJkbpCqtPeaar
/CWlixZyLcKNginrfK6XyXTrIzEKo7vDuSqbFm0/skr47Wn/2T61IUyBeiU9c1TE
9JDRwZ5pwtxEoszqOJYrXo3H7aVAlh1Ri+YyOmPkZ7BH7ZWw9XM64dTkrlcv0tRa
CYwa5OigD2M/COetx678Ks78t92bvUNsXDlEoOjsCZ+A+Ow1Y3JPu+S2MaP8idT5
TpPeOqsCsGBCH8IhPq29J/TOInbTwhJjzwV4Fujg+mIwAzsXiyskXon3ESm49ItT
1e7CQ6OM6Y/4VvyTl+D31GWIvhbcoCBb0XyF5kCIxM51tUUtORnFC+1hNtYijGUS
6ukVAq7kKkfVhmG2t+8p7Cnc3ACuMQdvMQumNE6pV/qx0R5kmo6Rj3Psmdz1Y1M1
TNvj/iKX1DOFbxxhXJh+AhkGkzhV8nxWk4QNK/WtKZJC67v7N6aSLEAhbYiu+Vln
PF7x6vqaPgmdXAJXA3fnYyMhDpXfatZKqpSd1n1WseVC57Itdl7FCNb1fohW6ANp
MvKli34gqXaY8vj/MkR7nDZJE5HyQ1aBXAskub16Kvp7f80YOAZHvUhcT6dm6sBz
qhLScxKppvgmr8bUOBnThhlsoSwR/4wt1CZkmbLI1nvGliqBGK84wNOSOpTF/ebz
PHLoupv9NU1OoQswEEXlmGEzPVgUypsYA1mRSs7Bh617edSNzOiwIfnw/j0sS4rH
+qawlqkgbg4n1BnSRHKBLw98lYVFoATRMoOGpWBTWu2uS4NR8dgfzyUrsWnZEbRK
eAIdErTpTyipo6W4szY6v4bDDx7W/GkVc8OhmSyHurXCoZj3pDbHaESe9T5QZLjz
h65UcQj7LJAFiNJ9atmPYbkQBnzx4vz/nETa0mOH4MSf1GIbzsFFdXbOqoLrhrc7
dgY3X2WegL3tQ0B1njstYK0VtN+3gTr9qJSNiz8AodiwX8xqhWvZ7hq+fWnM6kNq
k1c4JckezDiqF6lhaZhgz5GqIZ2/ovoTQQWBFe5deor9G4PVoz6SbTX4X/t9JzEK
ui5yScJjY0vj0u6kpiAQj0qt8a9dNQ8/sQWHGI+4nO4vPh+75h79524CPxbS6a8b
zXBF2DRbhVOCIyK23Nz2W7XuTpP0LP8rPTYAz2fHETdnVSDI5VBtu9IRBl5itECy
V3x/FvOPq6wxhbyhc3L9sDUrNFaWXfGNz8wmXi9H6x7GuXRrMUk2nOIJ+Q1uU5yF
uWUTbkvTkB5eF4M4wE4rvuRZPbt3q1xHa/F+f62KBFHQ7KQLnFZYRa2SLsx/M9/c
qVXIpduoc6s/nHMfDI0HadWKB4nsT6S8NoIjkzAmXhMVXLu8lCWrO0TqQWRCiKbl
o4dtTprnOYSy4pra2gv2mii9j1FkBY0FpBGuofJzdcUso2B7WnpfjGCiYuXAh+0i
CorKD5fYMLz0zwHg0njQU3f5dldYH4DNdYf0YKMWupZGd3ePaulSw8FRYBssbY87
pcVbUgbE7rv1v33JrCqS/lgPPXSkIweRX/A4Wf369OV66WUu4aoAdjWdL0/0I8+q
gWStQFxXY31WPLBo6zcFitY9ALSNs9ji1VquunYgOUy8tpMBGAzJJqgjVUZhvq6v
Nb0pvP77F9hZGr5j3uDfLgRXI/xXWKJQSGDSrynyFr8+4sG4enibU0yCrvJ+IB81
TQx5IuE+/kD4VC+8gA72l2DEo8rUCoqKr7hxv3CZWWNVA6m+GlERUSTKzQzcjkpE
L5yX80AVXqFNDi+bjd1YszpfoHzXtamYhH81afYBKFdmXPoz1im0czeybHrmoUdD
yE0OfeGHacyERas/WX1WeozDql/PutreXxnRLtIrldWqAwP0jvHJe+NHx5Q2M0n2
BGF4sS6/dDqYNm7F70uZIio/nZn6dL7Hdxa7XuXz5//piW7CDjuf1N7AuPLtkvNt
PpyFCBCU5g/nqW+ZjQndio4zoq2AORSx0Dxcz63rXKVxcENVEG1rk9gZnorjTgif
SqBX35fQ/D/d07THrWhD5OhPB039u16Y1K56LAgUS3qfhtjp2XfhbqkJyMF6ITA0
zAM6Pg46EgLXltuAnQCk1RKsGfiYFVTWl855ZEjCAXsCIdVn60WC+4Kevz2sO76z
Utmp218gWf+YaAOIDDFRP/UQU1kQrxrdLEP0S3hhDc9MSq03vCX+GOZY0n8i6fpj
K7WaGzxyl4d3AdUZb24JOGk5ATshF1RoJPXhiemuGkDjxecHIS3qeA9Pfi7mJWEB
6FflX878+yLbSzRI0pTvIrZZf16gLTEXDbAF+53zSfDnhugI3gcRdAvzaN5UBxFd
+/cnTNJr622bK0r6V9QVL/SYclwEiM4XfIHva1OY2TmxDJo3JtkoflqKCyvKlosC
YdQuKx/nuQUpcakF6G6DFcrZvIeJznt2HNufMkYFVnZYvEHSedGeWSqj7MpOaPRl
n2UvSPVqpXrMrJeR4flLAm6vQHBK1bS2vcrirbucVEAcluoZiJwzCwBGE8uDNybC
MR3WlBYGRoh2ItzLjSpglkTMFuelxdkI1RATYy3sKcO8RHYN3aW0VHKbdecNsrnx
lRiz+MKetoTTBcbar1KxCAdF2K5bxizOngePXBKMeTJxdUBzGegLJwAKJg3AusCu
RnEy/ap3sJfTEawdpzszTxzhHF4qf6ESBqmuaejYylhzf5OvhdLVUFF9paDHLUKJ
syOT6BLtugCPneaI4TpN9KhgfgfQXkVyaYJcON2Kv8kAUf0pO4EZqtQVz4OZVzyF
+332eb+MOftpAcXvNAz3Rs5ae8UCe6Y2r/dovy1wN+HN0nE7X42Zjes6JT9eYtK5
9k1ad/4lxJiCJvtKFGkQiTG0eQVm3Vy33MJ1cBGmRNak1CJsN21tQ2bOYJjZ6FYZ
WBYinUJ4ybZDzKZ/ntg8Hy2D++JGpmJRwOxCTy3ZianJgiYI8Cccphdgpabfz8Fr
ztuWcVICQs4hCZ3mP3g27hrHwoKX/D6njtrGby6T9DC+iGbDhOpgsd2JBj3G3t2T
W1e8nWgXl22SgNaxpsGkK2SvkS/qW9L3bCNnpxjagjxTQ9VxLfjBhjgU0ZhPWQZr
kTYtbUKrKsz89zqtAK714Bk0M+ixuOPsXbqCiFIvN7ihtRkqzm9udGzW6/bt3pQD
wzeqb4mJ2lzd2Sc0sz/o88Qt5umlQ28n1G+ya91Z3vtVR/E3vrirDZ6grhEQiJ01
EP/5VKJ2kSxrDfQ09VM+X+l9l8EB85KgTGDtsmK7kbqgYmGylMV7u79JVS8U5jim
AKZ+dCO/ICVdo9LdLYm9BoqNs46Y6Rqk2CBlg0p5vsl60faF6Yk7B9N9Ns2St17Z
3tO4QlRg1vKOQH8xZQKS2juFoJE0p8oqehOzjyvZC6xq9f2+ZEI6MRar/n5jHsbe
ZV9aql4lacguhuefJeOHPNuHkPjKqmzq5nZCQ1A4xgaJKv3g+oWPF1ZhmThKorLY
KIRKGKybTPn2PXlJK2ZxSgEwEbzrIM/9wVbI/ARSuyTMXkhvYA+90DWA4YnWlS75
CbAMo+T62D429AeGAuumgjSntyE8WYk2FJHsWk2SdSgZztpReO9wrMCjsDov3Dd9
Co9YBug1S3wgvuO8VPHjq5IOwlkzpV2jtPWiSNoWz6pF+9Ni555/modWkAR94EXY
q/jA1x/mWuc04iH+48Vppls37s7dS/XrRc6PSkKw/PQFyx4nZOevE7GXXQ+Vob/M
0TTYSu5Sa67OwrL579sUrqTBe8WzlOX/+ADNr5eXHRxky6QGPZssFnnjqYU94Uo9
+5IxcIsHpH+rDmdNMdSr+OAPZf1StI1i4T5cn7cI57XmzGFjWcdQb1auFLPbY18a
qOkATxtclvE2BVGXkdGOkj9esaJt35MuqSKpR8ILEi2JGj4h5fJzCCgXK+VhRVgn
fZESUx7a4tYtQrTYYjp0qyICOYwDfqTDmOtOkHFwx2q4xn39WhIuMsI8pH8pkrx3
UiCoMacIRk0PIzZhRBnBlMb6ZRoBlEXdbnU95rkvzvVtAw+5VZnRahZwQf8TMTpz
88zAkL8c3YZt9/TFcSHjB5gSVS9STkxK8AJS/3Rs7OOsbuGUaijBHk1jaFA9jlju
QY3FtVOfjjS+SWLE3sYb+A+xuHXCBb3VM6qNibFan5XWuTk0k9v3p2KS8kAYztuq
RtfSye2DtktSH/3DIIdHr70vCpbVtmfzYeS9cDTZPCU90qPb7CacPG/DO/50WB5Z
/9Wp8VY9PXxR4GIlUQXhaWDfnzHZzGkuXpVwjZfcXsHZjL9KgwdasTsIcwvR8hy3
JGNutlVS1TJ6vBcZKmch7CSdc0fsN/+HDY2DxTTAnpUoT5jQu+BeOUqfCWW/WbZI
Yc6ze0JtfFcpsS2yA8b3eutwzoGqZnizk0fA/gKGH/FpIHkOv2lRiVACsCLKvuLk
5cuIbMHmngINKMKzeaLjZdOlWzdiXgMeaPZjnlzfgT5mgUs+7vLlH5ojXEwXU2bA
Umd+YLYQVwptW5A5O1Kz0DpyBC6IalE97bZRjpI7jXu1T7vHwoj1L8vXtsavckf+
pirmFhX+3agAFmZs6a8RSAggbdL1IXdR0W56viJe2Uyzp+DV+BXEccdQyEDVWEsr
eHf2/lpXNWadQde7Sik3YHrgaGiqmTOt26OBAROshyxIwWajUfDEbDQFiIdi576o
WMzyjlY6G7kWaeDFBEHFknTz1E0SFwyNThaEhKjA9We1mtopvsjPP2FzhtLapSRs
03DlxeXc/ZWV9iPLnCLJNxVGO7wDj+qDpmOLAyjmBwUDILhPUrQYzedXcNKoq0U2
oqlbWW/9oKnYbd2YWzamHISGG5LPrn0ybSp8qxmucB7lVfzSlv1grpbCTswEDiW5
ijVQ4hL4Fz8aeiKTKnGvPheWUWMd5kFqrSlr9oFVUTTsLu4F/m3ePvRQNDKJVhFA
Y7TSx7MEuYUKPA96NVajN1EmlMU8ZTlOQVGEHjE/8dtuU2S6/mln79MqYz5dBI5Y
ednDgA9V19d8+9uZJAwnfn2ztdhQQXQd+XBqAs0YCq8Hxy1TlCYmJdf5h8AsoFuH
srE3+ipKFoX76uVKW3oyWiWo+lpd7fcRBlvh/e+ARCehkCrxfXcUwZRoMsmaHNIw
/Wpk6lr173AQkwSuJ0ks1H+FVeXa12uVjrCTRcBDSOHVmJEJuTXsYm3MC7eM3JRX
ziSII4pV03O8D/eB9gnuINU+K02lB+Z9eiAUYHAHTw3n0q8Ir6h7EG2SVdMD3fUQ
sYlicbwHVchcebu9OJTTG/w3FoVQedHDRfCWRutPsNq9MVfWiDqDWfvH5DwRNJaA
pqJ6wiQEJf/WKKOVxvUJW+t0XK/Z3pelneTv8GXSkTR67JHw7av2E24I9TlLY7f/
1ZHrdBx50VrUDKHXwir/ve4ooUvitNJuzTqtgbXxDmrCubZ/FA9OziNu7AnMZ8e0
KtwsCc4P1wRCajgYuNc4wZlp2H9iJdgrA9UsOgoe/u4dsVyRwRpKT2JVLEu+bPgJ
hIHXVOmLK3fHHp33MjpdvvY2dNVgJSBeedT/FhvgSxMyg6IBpbkL/SkaPC152F7v
wpnR+tCktXmT4lwqTicO6SmFeGCwVAW7I+xy3BGUtNTNOk7YkIlyhiWMsmE59TXK
kq2ks3Rzumh0e1f3CWadi+qyayyHBaoby9hM7EQDvN9w1sXzSHAN9TnjVIm9uQRm
sNU5DK7kTpJpRuQLFuYEo99uHT8nbzIT9SVXVrvsivA+EQg3ivSCL+9fVsDEYLa9
I68i0iwnB/u8zbmibCM6gzyXhNM33MWg+q+I8yL+SgC9WV7TfCZ6MTFw7Wbfr4Oi
0fMbHKNlBIFuQRQAgBPibeOC97CpkjP/uwkWD/CCjSy18qumLYMw6Zc5xEhFSx4q
y+gWn9p/o0qAjR22Dr/mHFcy+eJ/ed5PE0ApTFwKohBqrdK/10ZOVFhtXf4XXssM
qlBY2f4WjsAbuX5PJ5T4A1OgjBsjwHbs/Be27xhfCQSR0DvIg6IofbCYVxTabcUV
Mo79x3crGvupn680mYsU9oPDZOpycNGw81YvHgBfuH+Py2J7cq1PdnOEOlgISOl2
yZGHAn1bECEFeqHIAY2Bql+G6mSwhYIXNwyx1/bMqSkiamxBtXwWGpx1i9FTvsty
YYgR/87IoJmgX94O/AFTRJ1pfvKnIjrDdb+jVVabvSLLsW2YkNSo9oatjwaABFj+
GzbaCV3YNQdetDOeSH+sBqH+USXCX/iDLOWf3N5ozO6QHC4DSceqdwVlv0R7YCh9
kgnyIfkdhwbr8he0OYhG4yFcPvoB5azyB3ddRRLXSgnUTZzfTm5IXAwMLLzxy0q5
Q2yWhRKSkBL+he18v0GPY6u4fIVaSm4Aln27BSv6KhyNDhhXaFByTqhIkXJSgNgr
6m5mL/n7kzv4E5MydclDVv5emmmWNxhS7sWIhlXBCXsN3oTxV/nI4flLUc/kEcaA
OHv3uHTWtw/Az1THq0aYxQp5ln8hGhw5oJuacVSLJzBHTFWpKzlHBp4M91fTYQe4
LMeGvWYJRuLgPRMEtCvtcO7+UkueO4uiDhw2FipJ/htTanUG5O/IWhjC6GtILfaf
qDFQiFswW8Fm2IoL4AcrHnu/8qk8mmsBR7V8U4s//srVLTGCP7ghoq1Pa6YKIVcx
7rPMIMEcRkBtdN55IQAK1lg3zZ0buekTEG48smWD19kH6zSYhZ2R6GFNN9TVkufP
ClYGA3Y5FyKb4ogg6wZJEfgDQFJKuC4MO8hZsHV/PgYWc1syJlJ3ZIEQpwp3Njmt
392Byw6OouurxThhXpOSUPo92UY0ZMgdEbC/uWrulWr8Ey7DFLRiABkwpmZ23zeU
oRf5Xv/26FfuyqS1cNPFRG5Aw4V30Xjv1qkUpK9zPYEDOpPqjJRx4cJA0TZt/uUa
GSWb3oszRE5FLASGnOQ5i0PSSIh0j2Iwx6bg1OZAKQQPAp8gO4erHI6sYnFo370w
vHcbqj+N8oXK9OOHnt2sPjtqqY0BBIYR6kvUrMAqPvL6r3S9E+KmPSrTbS+1Wy3Y
Qhr14ICKo51kaDGy8bEflFW7C6bbkJENxDDZpWctnkIVfmhYHZaMgEgRdIlYnWIV
JJDhWEzE846Xm8W7hd1zn2cPNFFsDebc8I06DWQUlK/gwpDih7smn9mt16Guf3q3
hXJlCLoV49I2KSSMSGsEqP/KVz6AFAjP3Xr1ytttCku6EWCqIKg00sGekLVnjv4G
asqJC4OORK8sYwBvZMK1F5v56awCIF0kqbuWggFYT89NU7flj1Hg2CbSCX4NVIsY
9P/LSQqKLm24yD6qrMVp4lBv5AO/79n94I06nKrelwdd+AtAnUfL6pw6JbD5JNGL
F5Z9MIHvN5UBFoewP53Yy0XFy6InaDRUfETIRB9UZ3M8tGbZMGrf5bzP6s5AiUbE
/dBSsXx83v86j1RcY8/MDuZVD5X52rRVRa/fIhnrQSxivFDnce7xnw6dmI01hAtj
+DOKyIlMQe/H33IhXZes9kc9sOFN+ql+t4BzYNkQKhwpQeOIuqC51Ecoim0szyRW
7efeaqM1oVFUVgj1MUN2T7B8PQcYI0uuzPHA1MMPDjNkkqpcaV2ieXH18msRv0qJ
BCdvUR9d8vISYdzbAu/RcM3ZmKc+M1Lynuy2lcz01Laduhyltr39cGs65t9DxT/O
nGTN9GRYC3gqjYdHngWn5+//B+ZYCNKhL4QtN8FSqD2e4B6+fdP0BtWFVQiaOxMh
PhE0aHorpGgPtufGSvfNQ8vlPtPpxSUlBIKk9zZq6TMfAeIJhyHHQ73Bpb/oyMpB
ftvPcWeuMVfY5IKLFvNJ0j48/CN+EyEQvbGZbjI7LdTP4pie9WVIyPgXXF++Mbd8
Q8piyiY0T4g21gtI+bsmQZleSpUI5m+GDTPKlgkPtFWRq0EUNAwH0Amzjkz5Zcl7
DhNfwb+vL7GAWnSi3ctfojFcstJE40yBmVs3F60YazIKu+sjlvGXUQFX1lS/Cn0g
IMPhjFwEKr/QaK/om4Pm659VkDCc2beId3ANJZMTP8BhlVkR4HF1GnmsfiQlmaXR
0BiUGN07NnywNOaK3qGcrNBlWg+BIhpCjXIYk2RyQSz3J9eJuG9sJsRTG8Hdiway
KoVv5pwCg6Bg1zKJrgJqB7w5akXuHO8UCAczDuU4v1GP+71UvgZWmbNb+TZBjjUT
vvxWZ5tJdvXSJ5Ag9YD8gVofnOJJZENvAlhEX4Xf78+ESdRjDDOQggZ+Ve1CSo5n
dFXGPbrB/IQb1kVHHJ4ezrSoRy5yPK1JY6W5zrVnriF6FjbBXefMutuga/9NPAfU
yFMTAz5ege/RIkGSKmXmNXmLnghrMR9SEPpBji9+2FOO/J5SAFHENGSV89MI2b85
jhjSx1GiTBWTRDz/N0uz3Tnqx61tQ5ScbImw+fA/SfK0dNRhY74tTjKyVs3JcSRL
pi99UVu3ywROKNS0+bHZ7/u6eXgCPUsp9XXdjsz0qQDD/7C/V72EG0Uys1/FxgIe
DktAvqsQbnskppyY+J+W3G1yHELj4hcOxK4bkKarKKEKWqC7ugqhUlW2PDZ9mHOF
jhwryQ6bplY6SC3bqgf3PH2807eVCT6bzrHKQSyyi90+iH79eyWQkJ8blHAzIsoz
oGvbmJZ8pwyNp76k/K1ApSCjPHZTAGDpwN7O70FlEiGD1W7EEkDnmx9ChqID/z1l
6tgHa9DyvsK6WkUUKbGoCICvwhSSxBiV0jzD1V4hIe4eHMTl2+VoFrkPjuE5Aw6J
zO5wNQEHXpArnJa5dnbZx/p2OxUXdTmdvgnk4dCSIqaB20u3KPclDshwmEpJT61D
U3+MJqEElFY9PDoSeYv2MaCn7Nmtga2ht0EjSMg485RutOoo4pWsBQqwD7Uo/T/6
iaYLb/xlIKeVABMGoELxzaz1lW06jX4H1/oliya6o69OEG5M01452LH53uYVntv8
2EAnzcNJQrivDPsl55bhWIC4x35CebI9pprd1Be/HrrJkcNVPk9D2NOqhAz73y9U
FMoxPmPV7QUw80C/ibnxjsn56Iv69L7xn2Hwv4Ckcc1t3SlAwWFgsfdFngWWeVEO
lhGxHVABtVvspCQhTJ0F/YUXQBQiw/I6AzxvOSEiFuQbjGAIv2x5lXjsXkC3csHs
OjFX9LeUgMZHRUExPxqTM2szBfDNjg3G8p0/5QCyF4CVJpSM55tkbg5vlpF8zCTB
RiToOZKt+R1t54CuKKmOjd7SYklQMNFluCxNAEOYnU3jtLVE4bDH35sr3RAj1wSq
BTFAiBWmfPkfhFD4y5SZdUF7sQEpiyyE/7d4CWkoaqvRkAaFBcLz4DhTDyjsILFe
QMgikuEJIl9aN1kQ66lD74D5CK4toe3Ocew0Wpy3TVOfboZOHWKRy9WcYLojEbnS
TeMfy+Y3+VE2FaVtNJnoxXnRZk8cCt6Fm1Qg3VojGqNBfvpyXgBd9I7ChLX1WBx/
Bb460FBpBtm4s9UJzxWaCqAlTpRGS6atzbw0hEh7BFf+cdZW7CxK/OsiZvL/T9im
KhCL63vy8jvOJvw2n2TFAFu28QlXEOQdo3ZcauQkQqZXgkFiTVmT58MTOxr0DOV/
wXiNrb0qsbe0e4SnhsE3+T4LnxCxhwYQO1tk7joVKBwiB/w9T/4DlRF4bqrxNc/n
wAGI2agZWe5vstbwBim3cmqKhKd6vcNPkHvW88ga+gAP5QMQvuSVYL66MXgd9VcR
exC/3U2/hZWgph7PZwvtYmooikuXqfTz/0EIID3M6BDn7hRDlgRhZHdcFYGbBLqE
vH9+c35dX3wWmi1xpCuWLfXci7ZOaN/SX2X3dQ5sQ/UrYWcRxZC1M6Q8Ul/MQoGq
G+bOSvDd18OYlI2Qr4VJB8DFErOs8wE1Yrbhq5NxhyAgkWDmCm4TT/kz6r2YTnnP
/4IyLUgfxZ4R+nRffOrOB4QX6n8WyO7OHKn7lMI5bMBWtKkOFLaxhmvPdFUBikKe
IEM9q1eXV9S7EAWC6Df1neKZLZraPWbQHdR2D1vfnmIfwSQYVWX+xa/1t9wruZeK
UpKlnY8YsEy01lGmCcw//V7HK+2E9sS02w0Sm7p9harVcka5snnqKO90FvHJdtvf
fUcomEwTfNNzJCb+cb3EhyJQm56ET9jXerX79v3Wb5N39mT2Tps9LB5ZJwc1NA3v
VFUwAHU6Miu8APcg8idXkXuSAo0TxLQMwk79C0g42H5hp43Tgzkvzp4j9G6g9fdj
Fh1Hx6WxrmRdQnnE1gTrrtFBAJMB42kbvKT3evClzDd4DeXzyyATyJrnco+gt3Bz
ItZRfmzeCYmfc+bvUsFDpfpASNaSzskWeB/dcknMO4Xf+9UP9Kp8cpK/BVJdyD0g
G+zRnGd5wPCRW0otGsHVhacpQMgVyFPKHhBQnYcP+ohfIJSt+Ilm1QOo5STJnGkl
C76BRAM7YPFo0EUtpPVJC3xMfzXd/nM/q2ykHFzuUO0R27X8vWmoWHp36rfSXsho
kUhQ9Eiqzi9kPnjUvMQlnfTELunHIxqgkyoBf7sODxg+hEJOI9FRbom9ebtWDAkD
RvVpyN7eKNF/DbQVgXV2V7PCLCCDegc+1qBABUNTfNqTKGx2VnEiWps0Yi0U9fOs
kbwMu8qHpbK+tltmPPVTs6MS3M1RW+nYnakf5Ys7Dnue8L1bjlwzuNgsO8U/enAS
J2oAqFg+QO9Dy042bVwsA6MvWihKCOpC7Y+Lyyat/6/9AVTJIoHlK+sD6aeCzceW
Fv0+DGBsnsmQHJFvHq65dgZaFze0AGYvrcm4omqe6y4uLouecWryrApi+8dEbIXG
lO85tL+M8FZZ6AL2OQXLmRntPMt0qG024NlMYYpWpf6fVv5EGvQGN6VS7vxopiHN
sn7NgA0rXaA+KKyYmDRZzLt8VyeO6JwN2dwp0RsHBLxhkeVP4RFw1mpjXqXV+R6I
rw488SWKFu1Vja6TWYJ0xhLPBZ/rzZkaQpZME5oPsW96hBnMQcNomo7EM6i/Upva
abTbLi+xPcvHlNGLpS5aPafSE0T27ksYk80M9TRWJdFrebDGjb/xis3NrY8BAhkc
pD0hiiLva3Bc6LOil44fQm+YZoLd80/EFjRO932NhsnKj6BWfSQiyt9SRYxiEKgV
SzLqt/+kDC4k0tFwXNRgQXAnAO3NyUXetBHo2TQ2aH2PLfNmwyqp9fmuLAJJP3WZ
LQ5WuAy+XZIkMXO3PvI7RnLHDYlRSaPOjgU2MQtPBeSFYCRfdaKCNO3q58oP1rxp
CDPd4BZbZMXHUbtefnNwJS4N5LPvDnThZd2Nem5DXNNljt/2msW6oCvRS6m+bRsw
DcEPQP/myaW+Mdt2WPDBVyK6ZnCgaKTaHs22P5B6LfGt+qZIbfgHRngBOXaX8L8w
EBOrk80nZMfucpLk26rWF94NxTGEzZJ3mIp6VGz4zUMMntRH+81inW1KDttm5SvI
5Do9MFf+XNpoKrIfW+5VGYCHl71X1KpqI5sXeONBw9lmuhMLQ9NXwoH5j5mhZNfe
uITinqAynIEylmE+35KYeNNkDKUuMJiD+S2p7G5ZQXIkICz4EqvTKosO2BhFH1MG
00vOUgoviSHCDlf4KZ9RbHaISei3U13rBWRDuDo8+2vGEOIFCHBRVTx1/FPqGFHd
BmUcth3OiWLQuAGvuSiYH01HILxF0nVz9OwhB2aHYe33HYdr0gMG6vAeM/eaTtPf
ndX4dXp4eCs6BbL5z126IDWI73p43mARVN+YFZFPb2+CD21fbKOMKOypd6hKHW7O
98R1e9ftZsn14ZEEUVQoqUGu3ifixxrESBxpeHts1qUsNAThVwLCLOSqwphPBbcA
JL/0VXZ+N0YQ9/SCnJfnbHaLdu0fZXWD0IjEV6UTHYynLmwa38gdxKD8nyCMwkMb
bsbVStvoV5kwdqgYFwiWzFJfEaMCSAHf5ng9XBYcn2RxH6U0sPprD1ya/+SSvMrK
2quvSONdUOYskivNVuK0axN60N19D5QTabeivylQAOqLztNODA6C0fufR8Q9LyKh
LM0PS8S0HxWrh8ex3op3Sqk0jNmDYrTKLBBOYbja09fWzo95LLgENuNYaHPXAkk3
Tpda2PQb7de061l6zSGN7KJJoJkimuyHMlzD8O4r4TyuiUq3PlePfs7OHrZf6lBW
ep7xHZ5e7qkRF1oufZ7bBOjLu0v4NBeSJLfQTS6PSA6w6a0js8OGT51KH3/rGytI
Yx8qICzVIvx5RsGbgcuEtG9UZDlOz6hsovxWFH7EUTlDkW872fNPSzYTHp5onCmD
YRIMxmvk5ACH1fYFr75pHeI1VdQHAV+2naDlmUIJrhm8y6tMacmqgVHotv82ZiFM
egkRxcNEIhI8iUbvqM9qtE1UY4GcWxZ1TEzl2asKeXLd/onLwMDg/tODIlg5z+Ea
udOaR9Y2uM1EnLhM+RbRjh45ttgs6l/BC5+4aHS9quKRhbTRoYVidw7O59QttJhd
h2dT/a5gXBJrVOBSoOwjbUsZN65eBfWtUuxXQRA5Y/G8/6zi2MDOd5uxBcb7n4ks
ZlJOuNwEj4MU0SiX9DhIY6hEXSth8BOYhjfMuGEF4ehESGBhhJmzCXPw2KbDSkSY
msXiQtoaWz/C4oD+CVVtgJN4dMrC9QsI+hSSAaCWu/9wabXOkTCxhr7v607FuprL
PG5eYNyWCgWQ9GxmRCkSiqjJgm6q3nGIIKecYY8xoRLo09jeGVnQjdpeG6DoaUof
H0Ibf+vVnNUO6sVNOiceklYli7ktxyG/2achlkYFK244NkJ3metBsumwx+seJ5XH
QkUlIu6Eb5kPu9cnbwmCT8ghMMnEdDVpP3RG1ptTfpzcc4zJsEfM4OfQBwridSxu
GIFBXvHlp6IUuq9SDfeM260ly4JBYjNZISlgTLji5g6l/D1U6kuWoHAhuSCPmskI
1W/GWAF8LcqAkGJi0HJ7fAFIAb/6kjVOXrflNzfPk2mie77CwMWlBVaoKA+bgK3t
a9K7x5LhE6EMPBeMoPowU53pm0aokzoD9nTZA1roDw1eejcNcfzKjE8qtnmZwx/T
SXzc5PCSK0crNn73ZkJZwuMyAIMy0ihzeR4bxh3Apbx1AEOAZR78mXtdHMa7b0NZ
4o4AQnPysCx/MegcvMeQnen/Hs0Rip6jHePOIC3q5RjPfPfvwdZuPloM/kq6o81/
NVdYh6LvF3xmdol6AdjHG2A+4NkvHhQcc1iU3Uvx7s4b3S6IQ82KhHUeQ//ywAjf
9/ekoDRaD1RloewV3El7c3WkY1PIANyMyrPBZbWLFTYR7gs5cus9T86SSuWMs7gx
yzdKZVJvTQzotx5gioITI7YsuTua5SOCtI79Xd8DNmcyHzI3l+DSPmUpMDwTX9Rx
z0+3sCN80xvdFAlc7fOh6QwxnbwSpLwzfKZuIjo8PTpMJuJ0SDCiTWhk8nUDboDV
o3qgmRJeUP8WX/s+6qT9m+WA20tzdsxyTzalujYXwdrIAGaJVKlY9VqtN5l/SxI2
4dr5B8zM+GiUeIg4SX93sXPpGwuj0pXdxDkcM5OLYQcR+gv5Ae3fIXvakwnBdoyn
o6nhE4luzxrc4vEV06kOX+/jt5EnQ+kwaYV6Pj1kKvWBJBBtXw6hjZxnBdrmrY/V
5o8wnRB3bbwYkMvPXiASJnB7hKbXY5unTnnJb8S4kbYUNmgLo8eMN/mouCEV/YlA
VOYvWC9ZXXMSaXlTztNEFOxi3tUEu8oo3XQv1BEILcy3X7Rbm78FRM8APLJw6+P6
ohNb+jHlaECOl1RDHr8a6JTh3KeFUuu64ZD8E6Opm/1vqGulYJIUyRQeyzdkb3mt
X9FOE7L04kJhnc7tDgB2JR/paQaER/71m83cXYV8yEdiV6S31opxZmlzTZQMN+bo
Antl4oxpN9XD++Hf1QGXKREBMaSYgOKo4KlfDNCuqSkWobv3tJDkqAKdC9Uw6ao4
V1ONcgemCCbDUJwBg61efKGpE/T+pUVXgcg5KJ1suqWpwX4BVAFeEewDT6laT7jz
uAdx0psQfH8fYjuMLi80wFNZTigDyvKNJ30a8ZrQHHBuV7fYWE9/vk7Kv2GKXdMi
i22W2XCpXyW88lmdKPBxmYnwFdWJ6daWpTtywiIy09P3D5IqMhmW1uE45mlB3z1P
QFIQiQxSZZa5jpxx0ZZRaQYw8+XjDAb9QNuaJz+ce5JuNeY70ZPOqfel6LNomBG4
hU+OmknRyogOrJrn0uBGgRCoBFOA5kICIU5qkQAZFn6KBCGXNNInIDbfC/wfjefQ
gKLtTGQySRoTB5/MuMoJJ8PcQcgkcXzUCq43aTuv+RtlprKkcFRRjR9VD1D7BULk
xsXk3r5PIw8VWFKxvEqcR1CA5Pxj42ehb1RD7P2383PDGjJyhsqq+izZYzNpFjgK
UJIGTeCelJrFQ/2ZM9ZufSoi2W6RIkgL+cGJUH+kS2LfPrd/tDFKq4XhtJr+W1+R
EP8TZIr5MerfoO/5Qb5Ezb/+c9AkLEcUY+kMBwgP3eT2RMM8uPWRnSO1GZ0ki2bM
zIcuXtmmEhAVn7vhQGiJ3pnq/8wA+4bPdkgIehw5i8o+GVVnqJJfniwJm1YkAPyO
5tpKEv4e0UFfQZ2UTbzV5pkppnyx0thI8qFex+I1V23Nl0CeiuYwP/l2vytH5p99
FMvsqlzG2wMtAXFO5FaQfnh2zW7D00iAtzyZiW2+vv5CZ8c+1AvLhoDvAg3r8HW3
QjJnwBw21t+FH8ExI6S73Iy4kLJ4ukvFjg3yeEAlGOW6Prh9O8YndqmYlQRHSbki
rBEQk0wU6ldg29UOq/mY1H7NquDNjH1Hx1gye+kvbZ6e6x9V9TnCMfZV7CQKku4m
WakSOTYXunYFnrOr7ldrsEXC5TRfU33SAD8Uy9FEgHag34yRQQ3VGiUgB92u9EyQ
tALyT5rhnnHY4Kmd9Pr2k8LjP5/BwGUUrIppoIxTbD8VNeMp+eHstU7MSR7++Ub6
rbpJYPXeJDTf3GGQTkH7cnAE2X8Dsh/dA+VIK5L1x22Z4ssgpTaTbc21/6TNPCZF
0RTgnyBg2aWl602Zw0ardtEd4DsztumDw9cZ6CdDDrbsEFgKnVA1GhwqbxK53yyC
wEIHLW5+d+/yvTfEu0U8n1YiTmwdk4JlchsHO1yhaF6Ml5Eq4B9cAFZkVM1vs/qm
9ReMLgC+QUUUIzJyUxq95npNP9BypGmVFJVhd61/pvBJFYrPWnM4+biAGP8cTbVF
NCsCQyw/ewQWJw4E17wtXXnLK1FRuRDyANPRbIBW4WEVnv4VkEAiqB1mU4w7boOY
p5qP0rJdkbaFAKjNtbmVP8d777ipLO//tPv1DUx02afRDEAJSSP508yU9PFh5jn+
KUdvJW3LlfixtqlsmtnM5pqHrHn3rj4Dp40OwwS3FtGXtwHV/a7MP4MpjdWKV4hu
wYwKOJWLREbOkfrYbJ0XNSf1oydNbd8v8Q4gkemRDpz/ZfICYzGH2boL20bgFoB2
a5d7OPRZPtnf+NZwHpD/5gGQDEdfG0gEjhPoQfvevT5zbLsOv42Lajy807tSGnVW
YsE+1Z5VQ9P1sPviL/IHCQosgXiMOmga8FgDJGfBbUEVyRXA1hXE76k2tzfTddHL
9pxftZiVieAwWqPupdqSX3YBAp0o3d5AfIAqzgXjC+875wppMvtngcUxtLDVNiix
1NgGXx95sqLo5TfnSoUWgo/cWnnT7LVMNaUYdBbIYlTRV9+dptSrU3NoX8l3BsET
w89ndae0kouDYZG9HCz+LAzC5aHJoLCtKdETkX15vzi97VPC5VgSaP4cyiB62QOM
bcZAJb7pND7ipYfkXA6a/fWysgxJ/I24YnVZbfEJbdaTT+Wxr3wJKDtOr2SBmiHR
t410t6zAB0p9jYzBbs0IHu6Nu+h5JG851+C91ePAEvUmeY/mHM4bwrpLKJjANaV/
LgOB4A1L2+WRPy1Ygd1wMGw60OvHlPwtnvlahJ1EyRshkJ9vZfWwENeDi05BV7ZA
MdAVC/zUzT1ox2RrR2MNC5b0ZcgqF20imjZifn6ztu0FTKURaXqlpzDcwOjHxfas
//BRY/RktFbbpeke03xn7zvk3LF7hA/OIVgPupdgitR1cCo18X3xgGk2D8jNTFNq
nuc2Fddm9o2dNQ1chbzRO01HtlLnW+63dPLFTDG6JfyPPVvRQ0P69nkEfzuCagxw
R/jgsaKAisCMoRA0v/zOEZdb9HOlK5mbgbcyJKMr2q/A3gwIo2+a+qOp1qXnFFzo
UONa1TZJIoXBBE/Qn7jEfBptwDDag/dUdlz7CpSE4+H5dP19brOEGpj4wFn3DARI
Mhr+7JFDU43i9NhieZB7weCxv7MFiQrj1AbcuHlI4kPQwvsemr0wHA9H7xjJAey2
xTBbu6Z8dcSi902qZtt2MFEW1YiDFYN2c7vVXvXAx1DJlhtMbyDjKBmM3DauvDIE
01wSwN6mnH25AMzVQ/RpSIYiLAEzCiebMhYJ0xHA4LYb9N7awYzF1nkubp/bsja/
n7Sd57K/ECfrV87mFYjncgygxrYDOX3ckJMd5tOHugthXNfzVOneZI+I86ARa29d
EjkWyvShnoH164XFDCkx3CjGsYUubTEcqVSz24GNq1JGmhRmt4w0aUfLZ9N972Un
Lcdtdq1QfEyMY110wo/nLeP7YV6yV5gaJLBZwLL8k2+N/cGcmlVbC0wDUigboObO
oeEYCh5Ko8QENfPKWlNr2J9rTUMP6+A843dOkEvw8HI9Q5MOuIZcqFjCu9AB0+fG
CZnyHbag8PtScbZUhCyZRorzzNX4sFeLyEZy3I1f47sUZLu3wk6e+6kEtylgqyCX
WngiFApQ6bwb2RIqEnfQNNb0nEdnoh6W8Zn6+g/tTyuu1JIUP+Ghh/aBd4NpmiR0
TpRK4VY/AqzvR1hkVlPp9/PdXJetMF0FTHXzjdgSojl5OJE91wsoCj189yO6Ysw6
mM/A3gwVzoIVZG3G0HSDznMS4enT169y+WpVRbiKzWZaWrcF7Zw4u5XpXq20Xv6t
eFnAkYHhGjd5wTatL0fzUIRnNeLQFboH5MB0syQdmXZobTUoZYfyyQ8GP5lYTofE
flsSMhWTbaRai+gwZGoJwa61aBFvF/CHzVexUPrqujxPGKguybQJ5d6OEfBW6fWO
95SAyqTQ8KLOHMGTagt3rvHmnOF6pbbSTYA0CYw+KhCfMTZ79aZ+kDarxmwoJ2c+
IiyjMwHKs3gmHwEf31Da/jtPRJN9K5BFH8Yo8QcZHWCN1+iFvSuZVCzMeX5s/0mj
FUiCBDdGJvf/ftQu3XQo6OcVoeVurxUYKiYospoj6JAHoOg5eYr6UImRtJHb5YA8
lhd/safPzcz1i19GaO9GjDSD/RcGo1K2WfWgzYYX1IxB3pJ4De/qsjkSTK79JZVs
/VFbVgGQQrE/9VKE3r68CjsAnHg84+sLRoNOELQBEjRkUeM/4YkXuD2/5qndIjue
D7qcAYDhCipWdPmW9UN4iLoldjCjcQJpyaLNFOgXXDc3oVgi1mWZ710tmjQSyhhv
GkYJyihFIltIcSPHOpYV9vJJy2A/5++LZY6AU2s+i6yIfJCZbimRPTO/zrm9zYlm
U/JLMvuvXrFa1CMdsCJCLt/Uyuh2nVBwvdBQDkDZMQNuPnfrxBOaNjSUCisHdPgM
AZdBxPpoTWuJxVm9vDvM8movnRPbSX5koceczhnxjab4Lz8XfEft6moIJWnYWRhO
ew1TFUjRVvFmahOKjrsm00H80ZVU9QU1P9Emw59hC5YKfXvIlVqeaoL0wlY8Cos2
hK2JeoJx3EXxM6u+73UrBbQKNqJTVbarLOO5atZ1zEeHfOU7QjiT0BFCrBRvDJ0c
DlreanieZA1HIi2EMrGydzrgfGFlwv6ILeP+uSt+mCBJlULSOmo5kUdt9KqnjDDc
QsFBnIWYWmCyVrxjezBdGgue/Ph9jnf9oXdD0huMY6Sbz63GaBSszun+HjeILK1k
B3jemEE9utgIPreXYvWTjNoERRlNIi8CvLECoOQBOz4mkVecaR7+UWbIWVbc8hVc
ACl9xNRa4xKspj/TmM/+iwMCRemVj9wpANO1WLrmgMKbP9//H54XSXLwnPR6xK4a
gIXoskBcGuKof2YIp9gkL7rmKl9dODnETGQgAMtfVgT6yQrZSVgBkYv/m4OR5cyp
hi+JMtRhQ0D8SyIMCi+hQhdDxI+a7ioMqnyo7MZ85JCqWfECHYPWG+p2DFJGsA8q
YbYljlohr8UNjJODEeCPQYpruZy1mOlVuLpKsWCX0sfTpi83oHZqXHVc2cG+OXqd
MbLxPLok7AOpIWlbkfd7IiGICLKmYzWWqONAYGijbFMRKaJtVspW+rJheZbSi0Qu
k4ob8MF7unulbUdRwTfsKrPZ1oIgioxZohh3/+CYYSmPcIgYd2S4M4Q1kLVSDlYa
Dq4AoLAETSO0TeAqa53rIhCqqWWd1P6G/2CORqnypsgr7II9SvfeY7+L8NVfRmG3
NlIvlKmhazQh1AnUWQY4vxbN3RKSYSN897cnZkqyB5E4Iw0+xmHJMRujNKhSR3v7
lG2DMpAPp706AJDClrK8/5nySW0ZWk2df3U/7yh/JIhanYZxl6+BOg+1SDHHCJXw
61bE5JZ+h0YUkN1ZNdrD5keXkmx8V5gPfAE/iASFp3aluz04aQ8jlRqoS+dy45iG
CUYt4A32uE/2ARHkSAQoR2EhcRRLdRk5sAvfBvRnB3gpJiLD9qu0q3Rm2TfzTggj
seQgXG9RtPR9FTdf6jp5CuxvvflbfxNwnrRJPKRjjL88SfGojeUOeUszITYEFNxp
7XHgQQaTRF/LsaXjhtIcOGmzsAU/2YsZCaHL4gVYLD/7IVT6Rcqoi8z8uddRDGiW
9BwB7uzSBA/EAFfjtEr2O35agMqzYO5/cTr1wtN4RtG1TVtaD2IqGShZfJIwbRVp
sMjRlCnXg7aWrX0ogrPIjDG4d/ooiurejwrGWtMqUTjVW1pMSYzRjpAnabYpNx4M
57krTiVkKu++aHxE4qLfvge8PjOAUJOfVZszb1MZPy5nI5z+J/FD/0T3/zA7qN98
eHB7u1W4o8g2cH+9Lv2ixiYarNFyXZNvcY3hPjrbEt58MS7TuVZsHSFiQbBfjNUr
R4FqgR1eFSK/qarsSdvXtxGLe+O8p13R+ijs6/J142Bdd8VjOhS8pEZyxPuztGH1
dRZ35mCVWFP4LgOYxbt8x6GhDdx+HMHDAH7XJqb0ao0HGaHMx9Kc9Jty86dhv+B6
Nh+BdTtrOQGJL6/7Rk1MU0oY1dwpT5uBm/UuEAjSxy9Ojtlt7lVsHX2LEz04cdW1
BQHQX4B1sKPnsLm6BjIwmAlxsztQ17xA0ldHh1DcEcH9Q7ezkZPxxsF0CK1dXZAE
thDHooKJrpKXEkNsatF/tUSjw6LvpkpHimyTC3KQ4smmk5L4AxBeayUQe07pYCPD
rpwxX8O8Mb6IPHuvVZBrRHKzUQy2HK+oPtqQiJW6ASqWAVURzM/UHGocUlZ4xTVG
wl2zQzUyIBy0NleChMbJbummnpRB+jLWCxvgx8nFv02BoVkeUFVGqWwBHItaigX8
UhO0VYDz34K9Tnj4kUqln31ztPZfPJY65X8K1W46jE7fcfb6YMfeVTvj+kHLdA0k
BJUzdVRiJNKkudN7xatwbGCpZS8FO/rK47l1XFS06HpVu5sFuztx8r49YexNvsg5
LEQofmycW3bRb9sfEt859HGbbN3WDPmb1jIJqx2lhy0Xdpq/6F/3EXRhg7rHLUgI
OxA128HTpzIe+ARIh7ORZl2Wb61pPZgtBV4ULtJul3MV5NYosGweYq5oCRM3j3Ba
kIcxONSESpfRxM0anhe2B1by/fu8AHxg/qxTZEuVIMq/zbKViJvVHboGaOweIWIT
2EJRoKvrHa9Hfsw8u3uao2Gu8au47FDuHHfsRmwObngbaCiufZlVV+1wwkVtvo14
O0rgqnLRPQtODEnyKiDGp9odOFEEnVBWS3eAXdotHwBL2K+yyxf59/uOgTjFHjsr
UwZtLnLiJTpo28fo3JL2d4j7IuQSum2fVHNMgaUCQalGlQQ0KUw536Q/IJ1xiv5z
S4/uH9pnfkcz7Zm5z6gSlbJhEc5BbCVXwa8Js7Iw0rW1ulPUv0AcS8yQUFRjrXin
RHgE7mKGxYTvpP6kbyp9WIz11ZSxeMf8wnC3sp3eYLIKlprqck1V+Q0A73t59oAY
ksqaed9DlRaTmQCZi/CgyGvuLJmFJWNbGcPPxpqgPmoJXEVddqE4tgKaEgZ4GXl7
RA1a1B5uUOh8G3n3hVa3SRiEuCjs53F/M4/U3mCanrGIAwurwol7xx9zANoq+3nI
ELfOSeuo8GKvxySwptjJH29JtYx9QUgmsKQZ4exVP+ulkdsVD2/bLeSfn0fE01wB
C+A9F3HeF/gvlqnArJHRL95ibKsq/tmFsSQLXFOWPq52J51gtwsS9oa44wFd2Fu1
pqs8YI/ZT+R746+tuUTI5kSeTc5hl7Yr1A7GGTZy3AoD+bKO+JNflcOWAIjY84Av
DsBk0ANSMwFr1Zc4sSloQapEsqgPilnZE6TUgfatfzU2qNKQa43MV1LB+h47IU9N
FayWyKJOZKZnT+SwtrEYnUfUJyKKxgKkRi9hb5zlnP9WIjPI5fo/+mWtxTYso5G3
4/aI6KrNa0P7+8lEMDx/HSGvHOQBDCtKCbqeA200DSgLQg6wcr2zx8sqQ5IHKp9D
2RO7t2X+H2oHnPFiGm+2+tWsMF+4i1UDmWA2AaR/CzpP5+bCpr67963iuQfnaeca
5MsvIuS+WYzQi8PfgTJTC+OOuv93gq27yI1HXeH4Mfodqy4qbkJahN23/DKIjwWv
0AoA+One2XV7lkw58zoFDjMtAt4XbvnY862XPaLoloWbXVVJnTQVysld3lZRfKlM
nbu/pqcvBTCNUuM2/IdbS8XxgheyYWaIM/fefg1lkSXz0HSvEY/kyTZp/j17exjE
BLPyiTtxrYliSWVq66AczFa3bZw+srSeTbrnkHJZ90XOfBDTv4/YsbEViDPAKmXh
veh99VL4K0suX/Zm/itL9lLXid0/GNdR67z2RP46llrcrD0Tm04kHra0TBawHYiK
iokBdG6BJqH8xhTdB4lBX/OskIu2QfzRm7UUaCLZr5Ge36qSLzPXoEI0W0A0qMC6
7uztaJ2IRLj7wFbvlSgebieKHCarwIWnI8ztLpuEbr1f9hmfWk6OgIIvl0ljeMjZ
wfMvFIvcEOdCgOAcqFGAla9ZJZyWDY6x3su98KohsCNjF7hAUYf+mhr0GZ9/6Yst
bvfJPwpC0AvqaMqIJFIa2If0jJBcFOaLZ7Sx8zDI9RKxaT33pKViXNIoKpLx1os3
Z0OaPnWmdukAqLUveVoNoo3YQthbDuqmKlc/RaMitek6WDxEIQQruDqP6gsGOS66
fFjdYmqGorPsRIBHGeihZkN9JKX43Ue7FYBYSMbdPnQfGhLEyCzlGxIib4ikXtYS
2F/GzUWAhF2KydUn/tzA1tUn04tNHAFEIkCechORSLDiUtN+iPC95WTsS+5zxX8t
F0h7uavXxG2bG5w+GveKU7h8xA0uGzm2/Lj1ty+2dR2iMbnBrUDNNy5u1fRJ9oSz
7+/Xq202/rfOZnT/3HyXJCumYVKmnOMiyTigOZ0u2nptUgjvep/XdaQkYUc3cLQ2
CpFXmO7LxRgnzAmaiN/4tVnphSpRVIHSuI2+NlrSEnex1OOcnDZQa3E4BQoGhsu3
NaMSJfZxBU9hcOVT4HiTHvEU0rlKCQmVkm1S9UuKZVg+vsWC4DXbb/E/5xYbdGrg
hherF3xEaNcZj+Lx0mZlwiHJqnQq3cb0R4F3bK5TjUA5QvgiFmavAhObE5jLXy8z
R5Nk/HAnib+9u8ztWWGKmdX2O0ChG7uINMyCO2BmD+tIjKQEHhdDmZejCm85KZ3l
5KYU7pfHQ7qngzgBQgWqX/j2imx4YgF+Iqx8YtQMYg30Mji48h01dq8s08QcO+aT
JMPjnUgmrjRw3KMCLE57T3+TCRMUPLda+G+VnCvclt47GhDDrScmMTVbbE+4GkL/
+sc08o7XrZai74OWwkaR8qc2MXKUPLjiGerZZDIGjffj/bD1dJ5O5b0AQ7+Hj0Of
G0sprdyIawMdUwJYbYiYUoxhdV4QW6cwlrz6OclCofZ6TqSNQdhGAEYT2/lYrUsJ
GN4L+0PIfNetj6PUWo9ESDyfkURIUXGZqhMOaihe2yphVNfK8eU0N3h6Q46hMXRa
N/y8O4SoXaqY3rIm8drp8KJYcggHddPNguK7pFHYH4JphE925Jvq4qGAqRwJXCkF
x86lzZ3Jxuiy2etevAEwL0icHcDpZ1ZYY50mEl6Sba6wTNQlliC8RmrS/UwrDD7N
gDyAdtJGSsimMbJUhiRpoqdQsiyxNDMz00LP/zOX85JWA6dWwiEOZR/3sxtch6zV
314Ykp96+z1LPjFH2vKGx8N8WTyrsJY9bFIm4R3XZhlJjTtqerstwJhhuNItoDd7
layZl43/HQpM9WVdguD+uh3WhzRzua3R/fLco3UYGsWfV1Pd8BZdF/EjO2OxnhFu
7XHbHlbtO2gVXTXGvVYfk9JA6lD7N/V0myoSK8q64m/uKfnveWFa2MTjX4KQCTeB
PI/YJh9cNB+MslCnn0jjwxfy0pJ6VqMBxeYjMK05gquPghovX487aQUdX65zPuQz
LzImzCfi/7/DzavGOKlJTxmgGrPUixCzGHKF/Ot+nagCVkSJIYHTvhol/ABPdzle
/2/pebWI1zp5Zo9h7wGHE9I2whMc88/rJfuO4tGH5v4BFFhgskYUlafxyQn4YK/b
yWLKKhN9OGmyu90cCqbCxlf8npY5F+7DQDPpQpR4YoTFqJsKk6oNCeYSPOcYdXO7
pyU5ePKDjWwUrKlYFmLaK/D4fV1iV7VrAfV/hnon0o/n625r7I3vbna3GZIrgTya
rj+KhbRJKhBRflAcB+Y8F1PlCtZKKyklY0oJTWiyLegg5m4nTCNWf0Rs3Qc9kQGe
1LhPr2ZGyALG6NmI044ufZEhLA1qmHfd867qzICBPewRahxXyS3A0+fTbTn4SF7M
/RbcSJ8cz63MKkom6kgoPqZgBx6tirTLQH8CKsdnZvNJ38q5GgbJueVxDQh7TGFA
y7PtLkrYnM1GbWZlaT3M5c386ih/KDdcnsZh29n4ee2PU/hY1pTEYyjRlNCTdXZ/
/SnQRXpIbYW3IE4Cb7Gz54Wm1lw2Q0/MLzINODfsH/Nqiqou1fx0TGIGebUekLbQ
Xw13y+7HrskWhOOFXGmOc7QHffwyOxw0c4ZxtKaEQB/QmYFTbTfBqvpzfg+R1Z1e
kfQOGsp44naYiqmlFEoNKEBnHrr0fqFKTUGnfBGJLwvB7ZqTc0SYkQWx8M2bNjpG
UEj+Wvf7d8yZanbEzkQcA3FqVbZWyk/Spg7Ojb2XlkIMG2JFLMKZF/flWSXJ4Zp4
m9MwoE98knpjMFgcTAczbtofKQyGrTAkAbEh/479tzYMBWpHuQWK9kxN6V/0itfD
AYU8/1RcYHx6qdZn5SYzM43YZDgoL2GrwSAfyVF7sXBbk44TLSHOdBZjXGAfgntw
T3oQvHvcwJdCgdF4IEwW5h1zsCiv/24t4NadKp6+ZUVxRc7B8JVLz7ZEzYec0KHG
PlAKEZ1p6j8eyfHtgpxWeK/UhD52sxHR7+33XmYmJfpP/YB/vAk5cJiMrD3doldR
7NFCorAisBaiDjGsVQvIPZTldbI0QRlloUafCohspRuyk/tmnnL4LhZbmrxwmquX
MHvydFj4apOy25+wauxpxrLyOvSjGBe/Eik3rvEURhOOcXVHeF++2vYzs7ccfy0L
CAEaCfg3TuVbZbf5s9kyYfq8+6BbzPgat67vaImA3Tnd2XIvV1y1jq9cv0S1P+3r
dYbPl0HYmVA/UQnId6cgVhPOpt8ob13/1t1+5RxGYYeXN8Pw0+7IsFtd3DD9Uott
K5Z22f+6ORyfj+cKyA/D1HICp+n4gKSzPWcYnrymZM0bFC1DF8D6WhMw3K6QzLNX
Vk49M9uxz4phZ96hJEQ7FSpwYFaE+UBVweBQHCC5YCio6lkBRw0uvCCATfXyC1Hl
23nE9npzSXVnKZx7NpbHAKN0qMRB/bv51yOyO1FCaVU+2KR9JiCbTezc0aB26jcz
GitCJM914j2ch0Emy6nIbXSg/zebGVmroCEbOlAb0ASBJpbN4wT7Bj8FfUzz/Lad
FeifzlpUeuwwvioYpNZ+wxTA7t8A04XFCgNbB9whEW/JMG4rJr4goDAVNzTVUe+c
AGe0COoB6QvGZTkkPjib8XWQuFNsunfquWKWPPp1PMz6P3lcxM1bxzeZ1Hd2B05E
EhP+t63npxwBm9c2jQR0B+4nlsJ4bpizPT0ovvdjRq6KMorLABsqwjmPYjgUNC1j
E2JsHafGRc1IpgkykFdBJqRFrFrmpzE/gxxamh6OBPrkpPsedXz2/vLbvN8+G5HL
GRd6jzkkfP0dDP4bV3NisG78cyG5C1sKPRKfQ5QlOYgDYf380w5MXv/P10RKeifF
cqxI0F9rNeK83Q4PYZ5fD5XW2Z0KHH1x/jW1EeKNki7WzY2rIkWMktmdygxOgCdm
C64yvV0gwJQ/ezx7rG+HK94AEQE07w8VTDYIMMoft9JC+ee4JHVAOEPqa6HckS41
dVbr1JbfO4aJ0i9IgrsJUex80sfC4t6ckaGArA7ntGDrbxMktk+14LtwmCIpHm4V
kPXUY5Oi5fJ0fs93Aukw4cpLt2iQBVwwgFTmaqZwdGt5l3U64Zkmq/kR0+yjgFRN
KZ9bAl5b1K6nKlYW2dWIapKHleQFYZ+ezjnsf9ZtzoViO/7CphIAEIYQda4W7y5s
NUc/RnzJrDkWJbiuYnGqkGYb+0QKYYDr2qHX6ADEBOugzMkdn9vOJMXjHZqSPb5p
D0oqYGf8PkedOp4oJtNue4FhHOAITgs/hzB6pxnn5Jk12WJWXgxNSaxrkKuPEh8r
4xkwxsHFjROuqhHPRg5m/32+ejxEj6ywM66pIy6nSjyoSq9mgdEmwh/j56b9zgon
ryihGfSE++tbCc1LJfnhJMwBPEmf6lO6/wiT5fQ6ffYdChMIlUk36GQv8QUdNvHk
8QNW3v5yBbaPmj46hcu2FCtAlQY8eaGKVuJRRkdRouhTaAR3meM+ugScDRLecWpK
w5cfOYGe5uQYzatZ6w7owQcix4gPsLHX4xYwmUJfvxt5E4txtjl5G2y2LNOlbLHL
CX7j/qqBrfc87QsZdbYqgW5/BH1wS6rQh3ojrQ8vYov3zrXyOJtrV/aC5TOY7C5i
RzK3QHWCr1zPM8YEQtL+djb48GOD9DUpaNLrRToZWaxCZFun/eNeZyGSdQp4qzm7
ztHqKM0/6JZH3xQf/L+bxV5BgWbUVhDkMtAb87/FPDRdRINHnvmSF2M1diZ57MO8
4rRTJud/5FWfPjqQH2fDLGJysQK8Ft4XncLIB64V5HPkzNMleAlt/YzKJ7GWo9eF
2inm0sp/Nz7JVOKj2hL9Fige2Z/H1g2YSeWYQKkennw/QuEpYVuHM2rPHd2bny8Y
MHw9lq4/kseP9uT6ZSEBbHshdTK5W2bUgZQiDBtPvMz6JYwauEqliNTMuBgCxvzq
wJADHXvYVgnpy5UBykeklW7xUG4Ua+AlqboRwj8Ny/jqt2e5M8767g+PXEnrB57C
QRekpzcIxV1crqGMJuy/1Tu4mZe8wD4pn1VnxBG7Uhc28t6ycidI5t23ZnXcCvyU
zezDXIzPXjdknEgypFiHgCRQtoRwiiXd0Rk7zozFSHSldPyl90KVGYatCV4BTBgR
DSWs28xrbTAnZk5neYgC8zFQrr/Pg8/ip282AfKJav8opm9imocFnfsPO1LZ75eP
JC5/9X3vb/Pfrb7IIyhvV3Jp2JFJbHsxDQrRUrTwizJ7pWfUaNF2UD6olxqXDWOp
7oTrHtCExaQHxqnT55MJ5SMhvQWukic+6tU5/jDQXi56fZTZW43ApdgsiJ5zIxWT
yije+0tLehPNVQMirk5u1Ecdr1CHbvS77d/4j3edAXryeTD073wjL1UEaEVsEZzM
gOt74Uxtovndf0xF/kAakC0IJn8uApbrT/DLumPsxzvn5Sat92G9/Q5QF6GJfwgl
a1Tko9TYl7qcTzxk27N5aZj93fXZZ5qQBfN/HqdGEkThR/VWaCCPLcCInneBiE/V
MdoUsE95ZVNF5izWc7Tav5bqAAl0+G0PbC5c11eUVLCuv/H/NnvQBY6HtFtsrL6z
FxvAkn/WVRAhYCPUxCZvD6mJrYYqjJaSB2Onz5RyBmF8492F2WxUYZLcGq11rT73
pEB6f7OvfjjcfCMP6JoMAGrqL49F7NdMbTlu9j1bcZ8d0KMqZAFG8hNuiZjywSkd
tD5NbSxUw1A5KcecHwtpBEbjCCGtdgq+OUWrILz0algId4B1PXyI72da7E80Tj/w
C0DohM1Anx9TH0EKiVZfxcfRdWh9mPdHwFdiEphszqjTmLiNEXhnzey4M/Qmq1+k
eNLmoxIKpfmfuKCzGh9TOKdxHhdZoxUma1d3tSxSmU4GvYk1XKZapDXgqUZ3Yluh
GiTyM2to6GpRWC7eQnIHjMHgqmuAqZXmhSdQTWPfk6dW7iE72xREUEV93Uu1oiKy
5+FOxJ3IEjeivnDCJb44Ca7/9KmDoE21tMQiIBNlALAy5PEX1bbpkRl1y0r9srFL
A2LdUaDWuvkhzJSWFyteYcOTu05MWNei15vaFy9NWirg5DnqNcZJh5Vg8+jdfxWz
GcWcchG3WGlnX6WKIMxwtqU5PO1fYBaLITprqyLd3PXQh7FrdNmLz2bDEz6ZpRre
zpBVWcw8vm34M2XhNFZPjdGkffs6myOh+J08oLLo9XLuFeRl9alnfb/9YK96OQeQ
zLd7SV8jZGKaecZUsg73Wu82FEhZ5EP7o6yRHEtUHvtOl8ah/8C7b7CwfmyxAVot
aZ1PwZ0FvEQY1KFfNnXuWsu5E84pnp/92/V/QnKtAKJZPuc5IdR26oGra5ji8mZr
Zls5GJ2P4d+Dr86xK5r52RI/5n/v7xQhAY87LXz5TZy7vqhWRBvTvLDVuM5emIWk
BhgZl0H16NCPm5RWWfwOWIKwuvZyTGALqlmOoyBt5TydQgARvs2z2RJKO94StTbv
kdbp+Xd4/bxbKL6eyU/osZGarZxYLBsW+iPOz790H2DBSvrYHK722GTrex/CoBNu
CNNF9hHoImuPKDSQGomy/54+r/mpPNGbH8a9clUo5nlil919RlGQdASE11UMbQwd
Z2Cd+hciJUrFo9BvqKLdKjILEzwo3nnW2KLDu2RLOMoiVjIJUrLE7BBkiDSu2OlL
7YvLRhazhuz8f+TvFxyRPNfZ2Ibtl4xMZqOHuGdunLjC3GMMGWc89oxu/xOFghnd
KvkkTxZKx4taAptH4kn/PMDMwBDMBexu9rugUWYdm9nKtHlUnZvelC/52DBSNo+x
EzuMAFzAaFY2SBU9hzjwLsG7vWUINzO7pdY+SOlpq9k6901sn8TWBbwqgMHtj52M
SdnAaQ1ICJ91AHwVLFUiSVTQSYJfiNyDuAx0y7kY3RxgVjs7rNm4ymLaEmY28Uwm
y7eoMx1/jQYnYw+BmOT2ADq+ybMFVZPbYIuJIdV1yerMs+AXqR1G/0TCnRJ3Ieyz
B1Srw703sVOyyvlLFMNhhLcpR23ZQsrQwSoUzO4CBk4RgEGYitMoIRcKegtFKDBZ
AUI1nIp1mkwwBrrsKibqAzlj2KnAIgV5tf3W5QLrmE+2NRs9pwJgoOaO8szytpvV
7CpzYE8aoO3AgKh7OP1/b9L2QoUmIw2bZk8Q2pqjkMyJuvEwKKSZQXK3m05PSkDJ
jEgfd8tM/jf7lXBjinfgu+09+4xBkBfb37DlyutwMacNoLqJ2WewazDseMS3QvBu
X4FYYfPW5GLg3shTASu6QslDhQwopHYea6DUeMNvsNatHTRTKdKGGc0EqklNk4GE
BIhxc9nkjCKEMR34fJg7hR+a/LACwtCuXGwdNLPYKwm2DwgeOMcGOqAXGSCbaSBA
hEFb8Eu7yitWDv4pj0H8o3jMwICgCcnrlHSBs1UZs4fpMWsq8yUe/BFybtosV26R
PsKPDNrW5QxsDD2lxsyjEjlrQWQT0Uvkj59WcJNs1DqqyzmCsrVeBU6xk3/atdZs
vKZzt084LDPR0hn/nlEt9TdkFlgoOFOz4iHRwYH0tUSKq7V1t1wB3sJTdEuLzjAa
dN29/d+58hhM9Ull6kFcKbZVVdx9xsOcxI5KeokIj8htIFkilTV63TIt560lLdRp
Pitcxc34ELKt454h9+q7XAYqFE6zOP+EzzcbW6hOVks3J9ImDnI9ye3ukJsickrQ
ju/9IdX4TMiOTaiI5RHskLJwMCs4NRVBpTC8mPAmrRgVS3qLgdop0AFAyFc5BRYH
KuqL2us3HwX+g/WIF0b9zdeKaltAyx6XdYkQpLlch7OxhJMp/hvkIp7PEQOADK+y
2mowYHEG8VKH18c0NfIAVC3pUmszDFsXH8KHUEOuUCzL7EWdR9WxjL0rkIXg1CIy
OaHa99UQcuJk/ykf7Q64ULvLmWPcVJ2MqS/i+NOZwyGRlfhwI0LwlETHiFI6zX9+
J3cieFmB5oXfagPIG6Sqw8eiBX2Szk40Pm8KqqN/0+d2m+gpwzmv2+osRn0bCb7P
N97eyliIqOewJUYYfv0jHuGeIB/Sk4MfK7SVmO8Me0gHQGie+GyHgdNU56O1ZeA6
FlcsL1RWSsLf6UIEWQOaSweYbjbO0VjQLGZM2V9z6h1j4BxKesJRYcuFaS9WBh5B
h+akEgPbm/ggwcum0c0vjAfTQ5Y4YkUNTnWmEUo43Odk9Ag/CNFwvyMkAmo6JY7U
wyYJKws+0SyzQKkYOjqbbwFirapDhssOPin9iAioExslaJxmWmLwY3+ZcVSRDRhB
FzFnihyiNqX+JXk8SisOdM25a40dhTyG1QIGbUndld0xyGPA3QJFOmeu9VraKOMl
EKLyYTfydsRBz8jyo6xrzGQGxMAUllsA4bLT7b+ItQRzIwjdj4ePj/dfx7LFo/ek
wDVjdoUChmj03IhEjcvcNFCWACTT5nfahcTLTYP3EOXOrrBI8PwqDLu83tlTbY1i
dxmJt3fJ34OWfPxQDKnzbagX4TkVTNOWcIkqiojImFeMkioULwXKUdgmIptE6PIX
Ji+SdzhzhQ4Ila9q2O6KS9yNvvV/5XefbnvE9xYt8N28/cpdt4xuPjgVuijrJ31N
Sd+yzqzajBoxaVP8SGyocaivb4OVcLX1cIHai4LqSWaU3QASquhIscaYnR7Lu8RH
D946jLFtrRCv3QxR9cq2XemHEgN+rBDhx0goJtK3btEkkztL5jMqbm+HgGR/PFEK
nGSMCaArnlMDbUDmrZw3vmxUwy/SquoM9F52dXQGnOpS6b5XOqRPdv1Hj+/et2B4
J8VLRySFYLzlEWwacjJAeqkbXU+Wg46A0pop1c0EU6RwIRHTMlC9ZHgu/65GuGmz
BHbZ5i6J7jef88RKRGbqwq2WLlCpFkRPNAUDtG9QvBmc0HxMjUmeGiwi0wGsP4Py
2qtaCHrz57NuNJdkldpm9R+8zY8pBZK5tP+x6qy8r+OhH1aJo9mPyRkfXWeB2SA2
29xBMnL6QBY8A1SdXDfpuEvcRxmpl5fBQDCoMUUixlpKUE/J9FtyXZNUyXjbPZg2
OVK9cZktc9+p6d8zU6Xw9A4w/rksvetkAXI/tCn9sTaseMTwg0BLp4MDuVFvuwGZ
YsDzd7wYj9dj6Z2bvGmAeTXogfLy7TJ2a31JygHYne8HtB5OH7UJVQZYCOd3zT54
RrdID68LMBJLODxIoGSsApjV6MTYS0Ys83MHejfi3OLdcpUMwPo9QAGcNXOOFKiT
ihIWaBj7PXeGSZz3pGzqqhj/OD8ueUczLyodlS4rvXzjLibQdwDcrUHLFn62L42G
7qtKRcG0cU+OY9+q1WznpogkFsuoOraEwZlzU78fonLlYd/ZVNcUogGoch8Pu0Si
osOzZdvlK/uC+SufI+Fq1Y+HHJ73MZO2JDrb0xbJB2PjmcMMFLWQLUqhfukywM54
dSVV0ElEe7HILX2mxW67N1oXP6z4Bb+p6diehDz8wzjO74pUwU5ssmluh+lctBni
2DkCkxL3LcxeWTBpkQJWtU/YzXQtgI7TKyMIFNyL6mnKgTASHfpN0EWodjadGeb9
TuYq15CZeRV5jsvftpOLdjn4dJ7kE4QcU0QT9JSI7bfGtF4ObWKNQFN9IH6SEIyC
GTqDO3lHqPNKTFM5SFtNtDXeAsk0w1VWZcNu6Wku/lunHn53nKwAx5Gm2BxccF73
h9xdGJPVN9eW0KQCvILid9f58P6keO4QpLHNtQtfo5oqav2gQoHClczvnO6FBW64
hlhOOiyluASrdZoCLh9pMpM2TT1YG4gKLGpNZit/Y3XhRkSuOu0TSoBMdZk7k1xC
aNRGjT1u2qvZbMg0x+aV61jB9paR1xqTclPrVBsdxQXyszzxhO5x3ph0OyjkVe3d
EflGoHjGiJYELz8q4JhOuL1JEKfkx0A0Z6A44QzfSOBhL/d83rdoDS0nwHi+A60x
FfkgWrLekqkX232AZ3eAJj2I+wiY07HZaA2HmiDHD+Pm1kGHnS8QQWMtIBTxOdJj
h44H/A/v0dgfM8JECkp9GCODpxcqU0hiY0q2El5D4gr1PW6Y1MfQQaHJ9XIroef6
FMm7ZMqiSBMR6Ar+SfBC7yZs6wH5b5EQIPo5Blrp8MjtAkwkMgnr1KC7DyB1U2pS
Sjb1SF3G0LwC0mU76wmvUWh4jpycCZ9RtcvPVuBpcMQQswLy5gcuAh0HPXMd/45f
VZbEjUIqUq9Prz/RGRxAKFiV0WHqPDJFqvnmx1hhL3hHtTFPp3Qr6ZoeThrTqeqC
610AZtLDO0l6SSIZ26oDga52bLdrr/IMWON0Ln9yXsCAvgSADPDK+n9U2WeREaRN
O09ET53CwcNuKFbzy/qhLHHnsMcWDx/Vvf1o5LXvm63qKdyreUyqJiUu/y96QS1O
B6s0sHnPkQl90Svd/fqX+aqXLqZYvxgWWiTbv0A5FCH3lXwO6GOvhEGvor1fiQkJ
A+OlCWxTudgPMHE/mmidlH6oHAIHam4lChaR42gvWy8tKZse+sCJYHJSec+yDnSB
laBtVSRPe9VsZg+v9nBwOsFejNH8EMFMBk7zacCqca6duhBY9SfMBIccEFlUpBJp
hbZa5Ly06wVQLliI9FWj1rX4FkXSVLBJJw7G7RnXnqWzWAm1qpcTLKuwdhRO2HCH
zzWfc+R1pvHzhxQ5tKas9SlGml5RRdwwA/6vw3QJkSQM5+uKt1uV035kX/a4LY87
ab5gQArdy9gfzpS9z4VEPVk+ZaWnG7bg6FiIuaEq6o72VjRhO+ddzMEXLPGN1RVP
1ws/hScZlVJlhqx21tmgupfEHIByLis4Dv9fj7A+mAd0oe9NSisE5e1YkL24qet3
H2v16HUrPqh/Inmrl7g+jaNmBaebbzoQFokFtU3IUxqfBI1rHd/9/swtY1aciJeJ
kYACwadQx95fntftv1RR1ho3Ugl23RLAnNZEjBdp9mpoZfl9xh5HZHKo0cYCPVju
5RfTHnzTR7TMIhm/SS6xibH/3t3Tn9ul1eUbnU/KpFUDULWgrNaidxd7+4kNRi8G
JoVqtc/Yh0smURL6Te73SKVXeOwwqXD8v+5w1xTYprnrDH2OFBIa/JFAJAgBDnVD
iZqNlEA5GLlnmRXWpQAmcMhTiYNRCaTQlSvqS2wjdzd/vDC3vAYuqtaHqO83lssl
Arb7heZSr0fJQCJY2BLE/AVdvZ5hogDPWb8mhyms7Df3OzlUWPIvj13CNXiCGhVj
u7XIh6N8KemJExY7iryKGPzT4zG7P6o37IFs8xmkelQv+HHbKJV/kNToQZ+uGF7H
8QPADCPagK5bz1c9SAsB9aufyAXAy44Hss/+y4gl5JKXvcVK/LqpWS3JtecZxizF
eyJeazMgsjDadUKjFZQrBZrKhOP+IF2Mb6Uy6ZAlQb8ASSskyHTCuj4MDPfrEi6U
6x/4jiyyhpFAV0qJ4mvyFG4IRnVvkeb3R6+/IPcR7syok9o3m7reteFfMajNHpcA
CIP0L29bb5CCGH3HdV5r0Hi3dC7QImAALAvFda7zotUmhO7/b70O4EMm6U1bkip1
MmPWSpKVNjYhU4nYJSLlx56m9ziWGOcEkc2qAIxzhq4rUByY5NN8wov5HBZV+YGo
kFHcjCAuoNg14TBn+V6CWn3o/7MsCRUWY3BnjZeGr7apHzYtVWFwjERXWEv3k/WQ
V8W2EDLTdMR3mzRmh6Qec+hsDcU8KZbsgxJaSuz713xZ2kL7DVOeRLPr1GPZzJaV
4vghg6/ZT4Y8VTGc7VNREe+nzATWkZB+fPfxsoGwg/0u/46EiWcX+WDbEOoIm2DN
mZi/d3sFvKDL7Y/gtKjssOkjfk+c1hQptjRtS1fRsFNwlJS8G2KkABaEb1ZEUcV1
JvwqQeEY8OO4cLPSfV7IpASWQdipf9AD4x2wgC5hfVtyW9QCeoulckOGtByE9IKz
mfN8iaoouGxwByuF7Lau+1DXMwz3MMwiGCHQ772r7tInKusspLUgccTqIoko0nu5
ktDkAs5ahJTPKBpfLl8sj2FFbZpwW48EuNUJbA1lc7MyKEUnM130UeC7pNPaypMP
rBfGjxfefjC0SZRXm97SjqoZBQ8RLe31cMXc6qYzPxmZehZiiIkIL2yXfCYC/RtY
uaqUOi+0yvXDpVJwdRmj+doy/80y0q86SDxeDw+coPKUis50QzON3gpS6sJEcI2D
9t6aR4g+hw33u6VdcAy/gIq4b1WE6rStxmwb+ZjYZB83bm8sFvVEJDOoOGE18vrh
6N1v5WIHfafACNWdkKI6FEgInuJVLQ8fID1GQgIUf0H3APZ4rwFjQWIrnteJZYNW
kREPCY7YoSX6iIHuIofQCju7qtnG3MYBAlXsgWGHDLRa/QFaEOjW7agIwjq1/LFu
JXiCuvXGoqrEwf6RY3G8pxWmPV0/sT8RSBB3uHR8e6Lu+vgdgpRJRIxe/JNmLWat
27RxrueGw43j/phJDAwbfjZX0QGQjdPiIEo4tYe8MKn/ustywcS2QvtKCsf2Q/q8
XnrEPPHKsoaP7FXWGVAHo+ECwH1laMJJCruhC+uhiFxt0pP58I9O+keNDTFOWEPE
ithxV/AiZ6CqOuPSE5U+lf3FvUdd+r6EXExjXug4NTQPqdR3X4lqYebkoqk5YVZO
K71oFFyQWKV1DPiRloZ53SUUoI1sEsdN+mVVlu1WZb6YPZhdPASo/ANcw7ZXhaWt
/ViI8bSuscq9J8Tf8OXs6SXXov63leFfh8vk+F5Wlb/lcb9F39fV6bIu4qluOtgx
Ew9xMRkFi6VUSrQ/tc+Ie1KKuyiqhwUW4IvM09CPqn9j3nJ/3Fiuf8qlBxj5hIqR
xQ6vY3Q4FN4yTGTkjyUA1L5HCg09ZC61MEBby1ic0uikxqjmMxRJxiPDaaBnxZ+8
PpBT1mQu21RZzoJbyb/gfWHomCQDsjA81FTJI/mN35ojuTeL+3MnBJO1Jq8lyT8q
N0kRi2dyfNKUGFRtB/oxEEk0WovvJL6chCmgFcNffjLGVG1cbOHlrAyi10vvdssf
b6XLsFikaRBiI09INhQY6LIH3JUQfgltx2WfXoUTx6RXEhmBbeevdaP+MjlxtXIv
+dAvxnB0MgCJ6tbsektXTPOgLq59SeeoLMnTX0ignKj3jaAyIvAfdOV3SKk9lemj
UalWOnS/2DcZwv7Z/jNaDaElct39l+S4ektzPRe6YpPAnSLqwJxX5kxTZ83TNC9x
mL/4SmPGxfY0MYJ3TZOZCA9l8UN7q777X4bTsKQu6XSsUOHMAcLbkmWcBpBJyUTS
hUAC8A1fh3epVdizcQxIQjd1D2XIjvC548pfAfHvav1pPq0WfkYzTypmA6yVdbVM
axNKzFG48JnDv/cSNrjzFbWAm5z3FRHelNxN0mCO8/uuCFIv9aEe4xEOFqdk1bbg
wxnL/SRbCNFezdO/8vzTKSiSH+81VEQUWwzpP4EaePt7WHYOs7pIEkQ4MvzVcxki
hMlWrp+geg9STDLjuVYrP9CyJcSofHx3PDFP9zQDLJ5ufC5ldlWIv+EWPnnCRGbi
JpICiF26u8ge+GATBphWwIGw/v7fZ3F5mkfTspX80aMtKCXVjht/I2CNUCMt2UM8
XuIu+N7jAPCo+uUEXDrHAW4XYwHjz5p8+qrb8bys/Hgc5zI/aIeN+OC4N4WCvs5R
s/DNSIh36CqpNcPoTyWRAKoTmMTN+TIAT1338QroBuoMtDzL0LlvxxQoUzvbeJ8/
mPZp6CXOhBFSU48lCOVkxqgVjsPSclItM3bw8L32E47ZvonXoizEcGn0DjyxaVG7
2IvrTUAEh5aYPIWl2fG/m3zR2aKqw8fcNVDpnsL201NYwl8+lKmI8qpOKkV/A9gy
CI5eI477ntVGvg7MdGMgjmaVbyMHThohdGqNRRxGe9BFsE4lbO5XHqiNKgXZowbI
jXcu4kCzHUEC4NbJXc21gneEXqXHR6nkILZD4FkBtTVNm2Kd3uUytsuZLEM2Qsv/
yawe8Z9jfzZQ1R4m2AczGZhuadeZSmlfZG4CH9hK0BLBJuZCnheTHkd3ZaZBbNIv
seNwRlfvJ38dhbgtEsRcoJX9CFQ8Yr5PtTQQ7lXAaTHJxYvrTREZ28FkJrogYTpS
qca3mCGcU8VjpX+NuPs1zciOmtHVZC1Al+8SF0EhDj0g5otXHnyBOeg3CYiVIxDd
HfKfpWbHSLJTSKILGPdS5gcrkG5QPVPZwItgU0W9C6I87ICYNvtS66QAeR/NovTe
cye2f6SfKJT6X2Mu0sulH14TEMidinlPaqTV95vHSC0aNrW/39Hv0SyMysoCtLDF
zy/nZYrllpRvL7EiVvpe5uCtEgpNRBAEaAtn2i1OgnCLE+03Fe/C3riMCDNvF/4L
nPCTxn2rFWPQgC3zZI/otizh8Dh8LNmM1g8gOL6Xm3FN/PZTx2vg+xE/+qFk0yG8
wDXu9udK13ENlkxeQ6iFkkSBVXH4dyn9UdtbWR0j5WQxha2da/dUlTkc7YATc5fC
O0NjpGdVCpqjXClnCVixKi70zJ2qOMUyYbHo/xkVeQAV26v36ng2bSUzxXyHZwml
9IfjisXjK+4cXtVoIPnj2dP+FQWAwoQY5P712xNbLgIWlqq517pVmroes8GjxWvj
Q1+hJRbxZ6gCf0cHGJptmoyRCd4e7lSChEjkgxm45lAgEOrnedCUu9Or8XJqj9Kg
sW7Zrd2PJSyv/nUW8xXmv8+6DGPlcfk73jtuCNJCB7YfKEsKGLNIATexmgS+E6xA
y9XuxT5gIrdVFhO+wILv1N2xvgGcVMdswbD95mjHJofsi3kOBMqKHHf0zOnVciVo
HoJhPiFArXdq+GLfEkzLR1wyWhVHHFY+aDo45ZjPiJtHpZFzSmruceOx7GWAMDiy
BGbFZgz2iFZHr5f5R62QvDfu8aWKra37qjJmnKK+dRpx6i11vLO1sKBjlCul0eWa
YH30a38u5XCJ9U5wILP6w7KGFijOM0PhLRrpo9nTiK97UnHvws9PELE+nt3hmK/2
sGYTO/SDMmJTvxOQOSv4tkcTC4b8OmwRqXsSX6mA3lpI69w8ziR/XdVKzHSBPvAA
A+uXf8WIDxgcaJLfoiqRjIAmdJnUgxWt2hSmYOmmbF66XtOGqORWYy766ixK25Fs
b0HZJ5LGErLUgTuIP+Yf3sfT+uIux6FX+twQZbV/sZz6WH7DoZbCndoGRFBoGZkX
oAvUYDMptgJpr+Z5BjApif3OghSZTG+bQlmJj2w7uygpTboYM+xjtnInNCxXT5Sw
5qAtxBXyM6z4lENRjWoI/ZVkM5EhLFE2a9SNSPhrVtmGJ5e3nwBikG7HHgj+qlw9
zJpCBorezx5ktaToD8Pr/gt9siOMTgGQ87JYU5rFaBT5o7RV0TmpeYxsaKGBbGix
fF1g+4+7TGZmSUmslCcWhIc9C795MdedAgVnmhvJogHrh3hAUp47CheOnkulG1Ye
/dli4BII9BOFOrHImW/JSojxoE+0HA2mjph921+5IjH+fgu09nRki4uS/E9rhOGS
vAw+9JnUmfiYKjM6zdHyBZqWm2YZXvu51xf6Ox6ZX52qXSmGr09H1yF1DfzFNCP6
7MY7L1OKmcrRJBJloE7hlND9xOaMK+8vuCAuDXhSQojv4viQP40FsJYp9CxTnaPf
QG1hOxj080mFNm1PgJvjcOAsL6nOjvrGQchkKeUSeZMw3KTQu2dEkZf7tutVnR2J
1Xc9fuK8ImwQZgRjGWHcADkb+x16sjaNY8e5jShk8514BWyMD7fEPYuBsTQOLtWf
QjKsKNsQGDV1nKj42TsZsXlKy7HvWhddZF+tPn1Dt0sVr3R/Po4Q5bnKvSfj54S5
at0PDgPriwyAzuqymt8OZPupD6LkdWKlIvv1nAE26ONODZeuDgj9sz64b5rPmwDE
LXMIDgJJqUfVOXv2BI13rOAvmseGRz79FQuZIobCLoEMwWr4KuNFLyE/2rdndDPO
lLpJmmooCbDCvehJ7ZTu3IQc683j3Q3B4MjP9WWkFWhzR6382JjNr3T94lEAfn23
nyp71Vc0AiIfULsLCTeoH+Mx16oOn5P3TyiFRZQM7iIdsykwwxJO7qohbPzqKTK4
I5jbt74rUFB3p1PoLel3NViEYjUpudA5KMwUdkE1JDu7QQ2qemc7eRhllv9psw9V
wEEFGzmOWsUKHI5hAYFOOXJKg7djV8sa9hac5IbU66wcAVFxIEK5/qm+UL5cCEAe
LYSm3algyl2U9GkOxJusYQ9VaZ/Q8+IFIpoXqwNcWCP+MPCEke2Msf+8GM2hi5eT
2hCl9cqr+8TfjSUDbeIFXLt7LfX5A4fOlniWR6q1Pc28pdjNuzYfWQ2rbPN/Ttsv
AZKzDEmBYncXqiBmVUAsqqry/RkKJwaC7IQ6w571GyluLks1KO4wqMI02hniT9Jn
Xj66r6O0mKRG6ci420JKu691M02YvM1eo1rVzpl+oidxTtLZKKdmQ8YRqtSBfj/j
gl9fNVjVV0y9txPSugaJxhfLVwzdbBtDGjeFs9un1PHCBuKgJuKK/k26RhrwQV8y
QS+QvAePE37yo539Wg4dTL+aPBKJziE3bt6SeHiemRyQnaSk06I7ws/MbZSHxEHb
8PiJLXZEbJm6zyTnmksOXcRf5hYdTbI2JSS32q5O6r82qz+ZjbQYcQyZRuWX69hg
jhccjXsjvF6GZ/e2orvXwqlie8J+Mq5aHQcRZa2ywScF3aaD2bjj4rc87A0LU/uj
3fswLmciPsgiTdsEAjZKKHL0jTdzR0cgLI+pVaCuuSE/ZAsujYhjymhONecsGhq5
MHkvNHhEeKavcjvgJsQfzgY9i4B6jJegykT31lj9pflPlQqLtiBB3BKi9rv0hY63
32F5f+roG9DPEcBnqWRLCs76kOJK6V08QNcjS1sr/svOnkY+MgUqmDdQ/s81SbO5
qTNrweaJk7tUN5X4DcioKjFTzloIpMtPnb3bGZgLzbHMGub1L4oHfYWSS64XheZX
/Ep7xAhljAetOn+UHKRTVgQO+S8jl4JAWnkNroAWYJpmoFzR4IsE4ntP/OBrzqfu
ICvRt11/96zEXn+0+h/XK2J3mr9p/L3dn9wm16NdeQsaGmZeSZ5eQ/lX6ejc1d45
RqqoXva1gbHXtyH16EM2LCAAYhmMfbrQLKYasiYK5XblTo8gxWB2MjzoA7KxNtEx
L8UiZgkYEqMLcZMfmyGDPDv65LxavUEKeDzcdwamL3pZjKWzsiW80+9W9upp18b9
iS6psfb87KjgePaAt4LmgyIytEifEWuEKMj67qKRHtTt5mq6csJKcKrIrCiNGrFb
nz1FKpiZkrcZcvnXDv5WvF/ffwhjqB1iKxtFQY2Rn8OHvtvsjCcLaQ+Gi9kMqeeE
vc/qkJWWbqdmSK/KQmeNk+6+FEkMrtr6ZIVdRG57nEPulatN4Dhi+SPVvgs2v+kU
uXXCp1YGAZFS7FNhuedPdXnGxH2MdTnhhwtDlJoEvb974ZXEwVGUju82Jzu2jdFW
tV1fM7LBtmlmBYFsPhE3w7NGuAcPRLkpcSIdlGU+Gb0CtWnJfwTZNq3Mbm/5QW0Y
1LEw/ackINP0iAoUZ1n/j1BVAaYX0N2+Z90SlJfZvnPCOtrlvIjJJiaiir+FHaC3
QStu5ubCgFdmVkiy4jSghGVDZ0Gj8GPtrevE4w1VBD1UrpbyoGu7You8SAkxusQQ
oAjXM1DA0PGRc5mT6wge+5bFz3+IAc4FZ3BmcIWTm9ZjxxgQVYwqVYt5SHzRlsB3
4CS9ZNUC19grZ2KRMLb2rQ3S2RflWiYZZf8mcro3NT4Tt1jQaVQPZs1WJ4LfYNrB
+wkPBo+4EGVG35bFEB9d46+BBxUiye3ZQS4GnaE03OzNMbnzEEwN2dawvMf6QQRh
8z3cArlnFWwSTMwhkUUUj7+1nY/ksvvlkrU9d0uGPB4s3M1egl05sv8ZwicBJt7T
cPbjxovqeruW5vItMdnWc29aAkhUtscqJNlJyounjESDVVW1o5eiM+cCvY8lhOt9
zQvujkMuvRLV7qyw5O8fW8GUQC5Ulr8yzJy7SaZZcrrU76wxgtVXUfu1A7CDO/2R
aFbmm4cJBaq2Sz4564DJWfho//smyBKPWIO+t50amEPwdbup15iEiHjyWvjC9Njf
RoresK0GdDURCyXa4bZwa1KAExf6WxqfwusjNtD5tAfJEGTqb5gQm7Ba0RbIsmZY
WHewi7t0PwxilETvG6tqEqOVPlgCpXTm03FkqYbDIf21stdm+SEFIdNUhCeOMb8p
t3wD3eEmYM1lA0Bk5ZZeaklhS0coY00U/+Ww8+TK2uXndH4dhueyl9epBLtNoFiK
tPRbIX8Bv1s7/T3XIFQy73uq4cV/9Et1m9jT3KJvb86TJRxuV//wZjftJclpOBNu
qRbfd0xMkIEaPwlPfx2q08mpaeK8gKlJwHa5xZR1OOlJPOfVtBscIHe67Ln4cayo
5eGGpMNRINfCKPVVT3Frw6doeTRA4OfOkad1OdqXg0BTNOOe5hLjish+UyYkyH6f
F41DgSfl4GkhQ22DFPjBATvb6d0w1W9rNrcHpkeJrTooht5hoXfhgKcMagr5W5cR
X3wLyra5hR0K01EjBkwL6OCQr+XP6rkvXoZ3NdqJNZpa2s2QlmqB19NQ9OCm+1l1
WSH7Xw1ui+36tJahZTg3OvALAf/rd6MQYxiVTcacVggG2+9MqdgCv5Fyx+ZX03k2
qk5wDLo8hK2DpRHaKZ5XI+6lOTNO8L2B5MkmQcYIQJH4MgJd3ep1VH10obZ/i/IM
eKu06teG5dBROWf7OoaT2B3k+0L3RS5+cDH8hwVJ1YlEublL+pV2pcMRrraEkB5K
4ma5M+hY8PgduamYCrFs4Vnb3CFJTKhhPnmV6ZkKrPiq0nPOrFTNwalia1hirlaF
5PPaihT0K8LXOSlLAG8JUiWKO0hIHkXSdcwwvxLNi1VLsXCb55QdX99WkmV/A7Tq
/QrQWQXya2hiKYoRmK2u0BrGrLfIRVkGeLO0uGjIEpeFv0SbrGc6UGVK4mTNHQQy
qJzfvDSvo+Z2eTaoS7QfMet2YYNqBQk07AA1qt8vY9fi6pMhmft2g1kJDzd/FKrm
e701/JzSP/0Tyj0ZjBp4q05jRp5wTgIbpBGHoBWobqIwzIigZB6lHq0y9/FELkwe
UjUpXwgTpM/7mUoVcovnTApiClW8AzZqNtXEyg6+/ng24F8JLh0oU/FjM2xc0Rrf
VAm4fX79b2iW/pYKBJqFqUPwPjoFP7vaFHIlDy0mSwHYHh47Sx/gBmSCg4ZCkUz9
g628AslnCMqhurkX70sPtY7w+PIgJgmvhRuSYQ4Z/oasmlJNjWajj8JKchJnocrG
X88WuatGgEWMFYtl8jQ/tHwCHHI64PueprcDplXRLxp1RfkF7Vl+G9bxp3NqXIaK
hIsobRE+br4pC1BP4Y0uuCIgjWN2F9vUE08JymdutfrumwczHQmkD4rpNg7mDA/C
d7yqwh5J7wrh32tjNxPGZKeHbLjzml5LQQMbGKgVq0aEmk7cyzgFniszHmwUIZLU
FQmlhU64LDYcHQtfMafN05kDorwpFXrkJCpztqNDUdEM8BEaUiMf7QXeJXfc/rmN
sv30BGamUA0pFIlq9iVZasqAa5zmOyG7CsiHI0fQu2c0pXrLu85lD4i1ehTDdylc
9GCOiQ+UH57Q/3pdiPGjDz40tBaiLbHmK00n1xxt7im1JEotsbvUjDog/zxLzaJw
2NO1uytxscvBKR77sUmxKOX4W6O8JeaMgbU4H72FoZDmcDL1E4HdeflBTYgotxzv
SA0BCE3Ktd8qjk0OcjOM7sHK4rlmHC0v5Ax/9SwfUimWcazNj74/jqCGymbn9Jsq
NPmP2kRkEVC3n+ZonfyoGFa0X/Qw10TxO3MHCtlP95GFZj9QHFLjgnXmLfVWBG1J
S/uMUuyi7TKKWZ4LN3auyHFpEffNbAGg4aS0hjwOAUkFt+nEyEHa9gpV10btDxKo
pO4+GPahcWPtAHLvYtNstTNtDc4gnrtN8Ue7sj3WA5+RXsVRkJZZ1zlxfu3RHfG0
iAkB9xVshTtGjCvgSJ/G/3DdefeAYX/qgrPSPcz9VyPDxI5aBgBeY++gIYwMG/VP
Kg9Jn8/vQpBv/jMrlYB2NFUArck9e7Wm3BAkX88wXcexCmK6O5UpibHWhGDgB93i
phhFoH/nYWG8UCsYlODmxZ1u27xJ+VzuTcIryZMOZgQdijK7V5hl+RyGSDgJdCtY
6+UA5CoK2P6k1mIt7LHlJPLiKPmfj9BJEXaq2VG2xs4shywfFQSyVnNE8+il90Tt
ma+UmrkriT1eiu3aEOgk3GmLBL4NKbr1wdqbpJeUGNRfPQMyHRlEHoJBYapJKehl
Vnm6owhftfY6L6mcxFcmeSGnVCiZoWdXguV9mDK2v1qFyY+t8XyPWQpGukijrd/z
FWEocCpr14iejqzMdXTvlwaM3a8U9MmYWsv2MeBjQlybQWzo91kMPl9zLEsijDk9
noPY3TB3Y7zKnF7vu69Zd4d0azpMsrHztLnb1jr8ydwTXZ1IkTtzkZ3caLmkxR3f
yeNEgcNYL9lfj9ZnaCwnM2kNStte1pZNHKLRfTrcZQXEDj94FX4RxUUAYVLEfy3I
/GHto8MN7EyVBsvsh3+82Uy3Q8WEsBaZvkh2JZjtfL0iNXzKIdo0UoO600NBPi3S
BDgD1z20zqDkDoIy360EzRfRYYnBNqkeVdBGh2tZgS8Z4c6pIqmoSfkPe6EAuO4l
clMyOlOP8thz9N/0s/NIge1xCWNpx30h2NJawkqH+rRHONSX37+9TGGJkbU8WtJy
uqWSf/ooQcDd8E75B/lpJX6kzJ0OV6/i0eJw3NJVScryELCUioo4Q51yRqX7hh6A
Q8HNXJGwiQsbYiBz/p17D/5caiUdt8Q87xlcokKzsp1cJQVXjcHEcD6KSF/hWnEM
Kzwl8nzbuLC/FCzC+bA38TaP9T+U70QA2fncIAqOezhlmfntM2jSglcT104kMcud
CtC3IJgSBmuty4QZgKR+nqZDOAxYzVPuGIIuIvWhX4425IKA41KtRJXipwqYgY/k
Y6wyuTuXxiQvdUvMuK14wm8erXv1hWTdvwY/UjPLU3jeETlMS4DmufII8yHS/Yxu
TniwP/q4hJRsXxx2svtt5Y3iHnOQ+iVjNg16WCvABVuHo0S3Oqyqoe9SFqyoTKSL
oImFswontzbvZpxtM3OkRjlbFYeQAzndZ+7pGrnMVFF4bYDNFFAPA4DeMYiZxC/5
cYI7qHBfxxNfhBsB8//VJp0iBbaxg1qZMwLZhY4GXFY7F2Z2FdLtkVBfipUQWjH6
UwD6Az/N/AjwKACwqCEnD6YMiruzfvp/lPq6/XmTZHzndHLEGSfeFoYmrF5723aa
ORNCMIxS11AEQGL7k73Dxc4L6iY13QQEsiG+dzJu4Gj2Yzrx1TrmQysM3TS8PjuX
rjrR0kwLmvNt5+94O99q24RJUoYVtj+s3CXqVfjpOcU2yjq4fhAtJxvYe8twhhd7
Vbfi2vglj6VczG918JgOEsxyJFIaXx25huY5DU2V/oVYrP8NSa84aVRraY6QQTAA
DcymOkjrEEYkGz3hILwZJjZviqBZIV3r6TGvHjXl/7S3pY7pvtBZSroholk4A7Df
TQDMH/U8P/Of1M1nE4ykTPBLbHA+oAmvCKgxzsW+C4HGUYlA1HdcSptnXXd/MErg
tXsRrA1NTnrwkxQ9kb5JsRaE/1+IWjw0/cx91QF4MqQxtT/DZgAdL4x3yruaVcmk
WRG+QrGg1a9zeQs1kcijqcEf6hlVPDkTOmXGcOqRHLfu04a7J0wxE/VTNPXj2W7k
avGt2t5gUl0RyNwatEcpn8CS92y1t9IcWEx5Ovs3rUlWW2CvVS81MRyCzrmLobz7
GvVnY/L1uYhTimfhmeFAim6c50SnF57NNyeXx8Z0ISJDe2swxGtTCtLVxzf6x6db
vkxbiyfVAewfIRW+RsQuIa6nytso2jABSJJudJ9eCPaG8EYe+p+RJoCUsErgyw7p
zgxv0UMwjbJ8s3c1RsHg46PRx/01Rr0n+eyGx3q6ThYsfwYcdqIwCw2wJVLl+zD/
UWwjpR7/RE5EZXhVyxBpq5FjnudeybnRJQBfcGbKVPX0jOGwy+WuCTJ/o6Eo6gX5
OfIg5s5Z9Ik7hFY6VvYkt1Qqy1yLncVNnLKhLqEzaX59/AcmgrLs4QPy5P3PSHxf
JXapGxwgRiSdI9MvTFYZvS1SXHqE97lxtB19i+2EzXCfwb02jn5WmgdmKTy0xpj1
wZJKXoSYUjSqQ0HC1QHFQZHpiFhSnmWME3g8ic9+kJ7cFofA+UAmT/0EWoiwtuxl
wyXm1Fk47lO0DjviduRQ639FEzvbzRq/WHIm6q3MWukYXRXVwbB2glAENRF/1XuB
IYKWBCZFDr+/JERCcoUF9HN2e93UYdKzRNlaidlS2CxZfv08ss0hdJvdQd3r+S28
p4d6HvrhWWdqObPvDterI9ARx3srsPeCfbu/STUPodNv56pKdwKDEDiqgLeia1bm
t7BauAR8+ZTpInFAVIHekSqQt65dGFwFkKyHQEuZ1MCdEjG0QoqgQsT/D4eOgZLl
8r6jjb8Nns84CnjYvWyLifCRzDSBEW1TUuZs0ztzS8KjN2fqQzVp1yahluOP4jsG
gjY1upQ0Hwn6VbuAcH7EUiYDHxodLdxPLBrxafIZiktZaqiWrwrILLYaHb5DgGIc
BfR4yrlnDn9cEWukFRVfeXyizOGSfNdX9Bj00tuUsN/TuO1vF2Mho+zZ0HgICH9b
0dVOMRvlKEUk5hqq4RIR8SLC+gbHDA+zi+Xrz6r5prGiYDjYGRaAH384hseORu12
iR+b6MbN28PsXafbHL4fcVTvX6Pu5FWZ8l/bgifF1WpTDfffvHJW8vSUje+XxRzH
DYMTu/lfSBeyrheFAkURfsoq/RCtPgXbNQMpKJXAUdwrKhvcvKe3frNcV4M39HbT
NM3yFFVYaLc697jQO2rUdHRuY+BawVoV6dpOr/Hd7TvWv/amJJQbK07LBImZD/BR
1QQR8lBMvqMWleTY/PMTi5YAJUqGw1G9pN/9PVj0g57OYXGsoNhx+DaJpjGciPPp
+HTjQSHWIOtgzBOTmQbz8eZpmNX2TbjD03byt++lcgnGsubKzVLVlXotELQLZVtq
JJkF6ElRLp9vzP01Ago+F0Bs8hZrSTp++0aLCL+4o3RgCxpNCQkIYmLwg7TBMrao
mQO8tOEonQpqpWTM1lqGpw0kBdYLc4grztCe8rZAs02cS/LSN6RqOrfdDoEy5Ya5
stFbVK3Nt7Ver44kdfjqFf9+NRTgIKOY/QDUuq5Vm2cS0FSJSP21nDHG/YaEB86V
y8Qej/GiP6xJpTomwy3g2ptsJLAzHn3Aecb/EA7oiG4P2ARo9jKRpM5d4WthUqE3
LJwSIBIrRlpzi+RL6NbWxIlpJ+S+FiJK7zq6qY9dQKrueuSh2I/VRt8y5+3Wcqo0
KJIeNo7+7yM4B04nO/u8P6tqBCNo8DZiyfwFVoE2pNHWYr+4t98eHhR6TeWL6obw
UHZQI7Vk54g3xReZ/6YtKti0DH0J3aZErO0mt/Qg7Q38t4ESmhGQmHbtaaEst7u4
ZfGEeSRHD/f8/mq5OjjTb4gA9Mhz3v0MGevufrAfHhTO+xyOW6BTlqyuQALWs7rs
8quMirlh8OOOXjwVgdV0DUc/GaQf+QTbLEgnFEvE/AjJAg+l60bkgDwGeJNArXqI
RJmBoMd5LtdTW4rYmMZtwBfEG9RQLqY0gNO9FdLkRCXdYSmjBP7hgXJZigGmsJXO
1rQcPD5XQj7B7LQE9OX9HivUkUUUoc/BchXDTQtdf2qSjLfHFHgTE+h2f9RmHQ1d
JDa2AsqunNK2TGE7isck1Cf92Jbcfe5O4ZPpMioQBMRxnvRJbQpa7Vc7fz6C0bQd
H1iiu3oMQ3ASqAamqTTdIshw8cHqyWVgBwRwpEnS938N3J7Y0BJOrvrZgfEsDDe2
rupMC2P6eaiAD5YULI7k5yoo8QDCVZQE84GjFjmIhAaSgbB0VHACZvQqZ1KuhOW8
yU5WHlVBncXT/9ojA1cEa/jNgrZVmDMMtD+tNukbEtfNXSxT9/pH/sjIUiDYQ5uy
AlcZXLOIVEIB5Cv8iyn+8IoU0uKGHscUOZCDEydMLOtzkz1FY+j/wAnaL0D7YKor
W+qIYMwMa4mWfRnBAkCagGxFTFFAchodeEz+x4IX0AYtiUQH76KmUtH2HG26Fdpe
SxDZo84DtX79D9qpttJvE76w5QUzztDjRRObMQxfg8v0vmQJSyjZPa5UL0egqMi3
j9i7TZSMuOJkeLwwwpsZsi8gCenyrkq3kvrQOpwJY5xty8T9g32H7xD8WF7FTn83
ep5a1u7AZK3h8v91S9jPuHm1DyAB9Gy/9+OXaKRiNt1x7rBc7cqG0VUGwr1BgYzG
kAIHXrN36Iw418y3zJVKZSFlDgGuxUDe0NWboNRE3doHR8mESkKH0FP3oJoA8wS6
KKekt3mmKQqnKZutJpJAhnxBSofoUvj+clBC6YMzdceBTkQrLu8B2Lco5ppc8fI/
ka0l3J5D3F0l60vVCG6DirdBpr/WNtxv2DVj/2Tdxx5jpCqMzSbTfJuVlkzC9dv7
HF0S1GtC0wmdfjA5w/6Ivs3vvJ4I4dfwxMF9/XgZZUcluEQQE9zhoEbo/JUWcw2U
NIkShNb7X+4qJ/9gYfjZRlq2otGw/2RKhKuPnzlkFtvVZ0y54KabyvtrhaZD9EFt
XTsZi77xm2QRf0N7zj8hSqgG72BJxm/Ma3ks5HuFwxmv26CGQco3r11+WDQVpmcS
Yl7a1TRA9NyrrE1pZ8UySx/nxJvD9zoNm4zJZkyw+euoGYdIRqKgYyt+tLJb+MLl
WOrfYxBSF4tkx9Nz06qRc7MdfTYbQlDnWVXCKF5BHNe4OoKAC32BSK8hJDZEzKDV
Y/uZ0pukIyqOsKRqReN1kIZWCMU8Ave8uHtlkG4XNjA/XB0afcSR+sFuykUF6hnr
OYMWquIv8NOo4zUCUcsKwd6YUxw6EIaJqNNBpLj3nz97HimFQjj6TJk4yZOtKdEU
MTTbQf7zb9iNA0NQUnHCvHhdts7PEsrADee5d4DaZTCsYOlehvVwGXQP7eMq9cG8
30VUjOOm0RasR85FYfZdDfLdT9mMYhCV/kt9d9L9CbXOlz46Lhiz8H4ei3sFU9R7
j65t5EJNLtLdqd/barnuHq1H8+7pHTctD7I5IFnkzWnZuYf1oAzu0fkzfZ+M5KlP
LaQLmpVpuku/3EoGUHaNKb6UeXhFLWBohHFaPAphRhrJ94s8aIL/mZ+o+I3fAhFf
VpLnZXi1/fPp1cySIFUqx9OILfd9bY7cY3r0KNxZ0MvZ8iwBVXBq1PKt48wA8g05
fHvVK2JrNH9BVpTaOqCN02gExnkOVviNyU4JGhJh8t/zO/BFMVXoDHWFzCHi4kXC
uAMrJ/1f5qbeyGSK4qBQ8GLqn/YYfTt1o/fQWFaQ27rRRX8qN7LFcBP+bOAwa34G
VDhybjf8xXM4RfnE+vfgKGMcdLPITFtgw1Sg1BSE8xIw5gPkXatvEywNTdSkUyOd
sni6b2mXt+TJdNQdVIH0R5j6zZ8A1YG8g3VWJ5YDxSbBYdl+1wraqDx2d/RgE6mU
+x9yr6yQ+gi7efh1qgEEl6KFQOXJ02RzNuUwXn+1rsnt+SNfMLOHaw3K2mKyqKvB
cPk1cP/i9isxRUlVN/FWaCAPMqappn2Y7mQ7khyfvlaqIAUCsRra2Yp+34mAyWVV
wgsfHRMZdomTPMi4cmGzg6UXqy2cBEO5ym8y4zrAW1VCKRWosK30NWAvb8Ea4w2j
xXA/GsGOXgzBUu21ockw9ryMdq5SWyNqjDULPkP7XV82Som0NXch3uCJcQfGhdoa
ISP8I+ZMIlAzyQd5860jOGOWoFzBLKLCFvDcm+uTaNSNz8XSykUAvgFibLrDLcHo
Jg3+VhuTyfhiOzK7k1Ma3ONBILRHSvxzNMJMA9swQjwb3atO6mw5xl2yPSqik15u
riyFzUCSMiaQVY9N1JniF5VtaH1CDOuS1nxMLk1N6HZD1Qs1D2bkxSYIjP829BTE
21LpAsdGgewCI9G2blJZ2Kr6NuO2XpVJRWpgvOWTYn/N7tPq20DgbENGVHqP2YvM
ZHaaKDM/gAgzdk02mDdPDuseyYiJB6MxLG/bs/ns4R5KvyTIxizyvie1FjuEBC6R
+nyoWHXkRzvwGTHXnMVSrFiZ6FwjPBku1Ah+QrjiXWL9EcE2EcZGeL7HvxdsreVg
tKUOJqWcOicjzT8oJEOsVdCfP5OQxUicJFjuZ6bOvX5osE4UgrW/5OQZlC3qwevk
q1zjvgZ3mZUQ8O6aecBfu6aZcTLk5SuiJ2+hPAHQO0O0fZge0eaC7bHGPzRshrR/
cSTuV2eojpw1MBDVeSeK2xQI0+YsNS9KmQ3F5Zo1UiRRuugHEPilaWT9kBwBs0aV
AaffFO/nMm1iejykxEmoAGOevt1cpJ173N6jZe+G9jsxu9sISPPs2r8+Q7JBC0eA
IXctMvbrSdwPKjua0iYAQhPWbLE7b1kLcyL3r1LPU7JrAL9om8An+9XSy8OipdZH
O6OAOUEcaAaMXrYy4xDqxuzvlMrJVAR1xb5YQNNmD3hUvqMrfvwQO4YGMLg9iACv
TregzoQ70F7avBCzFwwwDsmphHyVx5pTps6I8/sxUJid+rlnyuifCrEdjaCVdF4d
1DIh5qGZZBEwpJqzEhDYLKrJWTwOIc784KHykH+A2o3GdwiJlzQHGiMCPNUrIdxT
R8C8cGbnRKmT2whN2kfxIn5aH8gfblZIxwlL29we52UsnfuixNRMv03dL7O9hF5s
McYspTDH0tVbKf8cPFYHMWQdPB7CHdb3nb//u+fZYDB2KGhLrFxsor/GmPPUE/pc
ZxX5ClWhahFWOrY+4aO4zNp3PGa49nbim5oczFPTxKF0PtW+WUYNGqE1m9xxZ/+n
ntSh9NJDR+KRwooBQGz0WPekSApluzQWHVkxB3bduHDZkBVA+xjq50hqA0blXdJt
M2F3x2YaphppyH+o1AGeJZqn8wW0MR7nDCtN2yzkHt5bCanB8/6ItdMRIP62owv9
cxT0esLsUqn4QAT02HM4qnarlEQsuxV4wpPZweHRamF58FE1HMxbbdu6qH3jYY3c
BZvVhd3ujgCBAqOXLP4WcJ6Eqgl4eP7gqmlHWGgNuSYFijwCGzL4fE14ZGif15Ck
av7xiv8kImcQvbjhli6829HBTRuORNPMDSHjnk/ZvNBsqebttd4pNE+Q/mjKzv9G
znpgVUSjJGTBVHpql4OeNTSYkIlhtxMSv+iMNUFiqY/iOLlba0DVUBa0vqjZe30J
tLWa7UKRB3X8KGfRqJ9pOTN6qNLln1+oemdkBgI6UFXXPVx1Pz5urwR95TLgl4Uj
7XLvOkUxNyeeh+KqbuOyLumybvlapqPxoX4hqMfITpukZtoEomVERAtSmWS61Bi/
FbxPE2jHRKcgZmlwUOyCPN0wpVutMFgppYVp0/nPHK5/MrGh5mzcpDIq1oJFhVtT
WHVo1/lHmEI4wcuGY7W9IgnK50jz+qI3S1SjzmzrpLCTeMOUsidXpQ3WxbxJa3di
3VqKcYtxhOqJAxubDqFo1LTEkOOU8usifFw5JHKlzMNox6DWFi/KlPAGs27cHjGY
q1OaGJUQTnrE3/nw4JPXDckp6mB2R/a/sceCnW7p5HBPcl8n7n/NkYKUiEIpxC30
qM7lbVlIY7J3kxBZw8lvgnPvUStqF3cOosfXl+ojwURwoO6J0LhK8/vWG4zslozY
Rhwnn+cenC4sGXuoPPjeh/ZusiB6oLvaHQoMXLNwg59IlPtv1p/rdXaxPEyI3EjO
1jsqPz8i7bHinsfBujGB3au9YEnBqY999pWY3YVQxuhGD7E4Re9Z5uDvB7xkE8+a
fCZJ4J+6CrOgaijhvaLLa/vIcz6QgvrvndS6pUVmCodV1PFbm+z3NZB/a+AWH9dc
U+OoTig6RdBc5sfWburO8RDzqIc5qe9gjE8C3cdYuoH3N0pqlYMaGXVHm7eBcTYH
pWminF+9W/SYwQ6H1I8f0EVdX+iOstg3SAqbMnc8ZXCMxkGRI8GG9O2WlhTpQuKD
vRHS3dDWLO2TW6gdz8Nxl0HnX9oAru7AS3AEKyPAkZKLgIX6p966Ms0RfS790M4w
l8F98vEoQXeBtSaAW4bXMNOZsB5mcTPyu044VanmRHDJ5v2TWnJdjVGPiA7sT9EA
JtAL1ZKbnNAmu06rgB6iEDbtcMjly5Eo0lgnSZZLkunJk+4V1JsJN0lY6b2yp5Hq
FMB/m1Xtw6OqnvYZSXiP56OY7oifhyhTFgSQ6c1mhZiX2rtTC5z6uxbnMUX3j5Cc
0dcKwd/07CizIBDzQNpS6pvqEhhubgzSh6TdrNFeN94w19UsnBEXgqLS8w7hXvrJ
J1wPtAghdOHgRp3IVxFnpmVE0GBlPoULrtu5y7RlaHEBHE87aDLsksxlSP0LV/RR
3Evg4N8HX2TE//BKS9nFViM0eUOP4dzn9QFW1NxCnKHMrXJnFjttzhyVChQ5d/m5
o3FB7OiRNoowp+cVO7uyqpPb0KqNI7PP1tr20fMZhL8Ku0V7gLdJDM/vMIKnjGO5
fn9sByx7ld1BMRcq5UifxK29olrnTFBxL86bHHpqGXh9ZGrUAMBMSIVwZloY5luO
IQDYKcVdrteVIR+KUE+U3WszOxpmwuv2jHFSinV0ga/QFGGULg+cqHZu1MXKA0pE
/73DLTLLOpWqPEWLjz8LsT5OyxJzZs110zD8n/g9StgOoW3PTmEPEu4vFrtcFgV/
NBLTOS89sBcdyf6Aj533pSJqa8mCrTLsSi/ZirFhuvkEC1zvhK0PVKBecf45kTb9
gvd7QPHe+80EMK498Q8ZoAKqrdRUbxZ3x6fW5r1ic6PWoFZtAxD8GcuppWZIAtsT
rOaDYEUPLyxMp0HUHceglW2yG1ODp0+7EhUMGiNL+PM01c1phlX4oQebSbetc/UX
7JCi9G1SBSNSb6elI795jyh1k4jkJ8Bxyi8xrWP6OuLkgSJNGNwqqtT8v4g5FIq9
i8fj3WuP8L+1f0lZemhkk4anRkizfejgb40ehkjSrG6nKlZyBzyLfMXruKgMwgft
ncbSM4D57NbHmx1B/R8LbMf+kxt66rMmYzr8WafFVOGmoJcYf6pSv4VjfZdudany
c+MwNxQx0aNQ4QkRg0ZPycXG3CPfkWp16a3iUjVjc9jd8GDy4V1KmjwJsChffZ+V
7crz8rNrnCP1BaKRNtpeeGKKVHlqrjDyPmkT5MhrTE2AMGFArtkMBlxcgCea9E4j
Y9UwnrVaazNTjOZ8XkmNS1mCbqnWO2wX/QhXMuv5nsoewDERVioFg47H3TrxmzP6
q95+OSL4SeQXYdSsww9qc8qAzagosJlOBkENzI+sSWWcUijgH3AXpP3jaz6h+4r9
7mIA84aTRLVN5O4aEoFhEPoNi973hnAtrj7phcw8uQcWz8VZUCqX28QZCahIj2W1
PYMowMKsrdu7nJBVeYkByfbQE5cMh8PsIonO9tlv+Bt1RgYnLFymucM4NW6J1Rsf
lHT6XCjKNu242sZvwjjhurb+dDXAYFgPUvHllyjG2SzQtDUhw0XL0LpDRuaq+4y+
V3UnUoDEI0ck4reca1jFhWIR7Klq9ZoiCWtPe9r7bGw9ZR5VAylpBn+RQd0d70YG
JqOdLcS6RHWr4oTFvVxHsHc25rT9gdVoZph0FrUdkwWpm1ADctUvHYem00eIAY2G
Em9KZKZL8DsQJjsjlDDicZorIbZ/2flbGIj/y2XWGc/TN7YufMk+xOPO87aSOUM2
PMKz3Z4Ts8z0XmMI6jEHcA4VLpzWdOLG5zdbz9HI42NJ0guWnux5S/EKD1viohfo
IGJ+pNUM5pI0+dFhZ+KND/parrkRuTv+RjxwWZgBcm3y2o+XOZYqT+DpTqRsKgo2
0/PoJIlFOMTkjEWWEH9GHrsaJpi6zNq1+w3YcYirfMnrl/mG65ABufPGlb4LBzfs
kzk274wrdof02yvmKhx5IkeKX5na735c0FXmxWJeFjm0VtXZaq9JkdYzjDPzBaUY
w02wLaJiOslqjDE12nNXiu1UMQQtS2HxCE1pXlAT7hcp3ShBurndMufvHPJGxcfS
agBhLxnFo0w9YnG1kaJZbhzmYllazYqmnU7+rSRXX8cnjcgHECZ/wYVuh0JtoN15
9P0vJoKSJuwdVygGzmx4YubFJzNXXkSp7o//akFdWrWxlapWuUreburVG9fL3a7C
kQQbkAeGgEvIUweW55Eh73EOANSpblsciDm8dFNzxtc0lXVGJggrIbxxzOJX1e8r
YTHa9GCMO53ufvIF6669r3W6wEdNyxXJr0XsitTNjyt5rb3bT7zmr5HzKQnYGNnz
8LX7UWFlEzYj6hpO0fFQZ2Rujw3W7NcFI4/vbuAsgGNbOKeTQujricqSHJLbaNlz
yX+pvfuhTxidJKmv7EPBbdOpgxwxKhH0fLMCO9Hxfp3cMSWcmplmZQo4nGfUIjCP
qvjUqN2CLVPDtwVFVvQW34h82Hbl8xTAOJANSQ4M4oO0gybp5w6HdqE8tavrNe4t
gYYiH56aX5iF6qhCDohbbL4xRfQrso9Cw25oVD1YYrlU5oz9lksIGCHMz0vYgr2X
fKzrGmTovzQSnylTf5i2hV5Xs/wm6bryRCPnxTtTo9u5Q1nhWhLhm5HRgRjlZX0S
7FcwgSgmhkLfulo93jKiuxwtcy4WY557pz+FVSZoxilSj/p7htD4LixF9usb3SYF
wCcfS0GazhxunN8usWGi37/YsBYjgWVdAXzaviEQdP1B7gP1FhkT6G+YyO02T+od
O45yrFaWQwxWJXyahonUYCjMqgNPJtcokOY0EZ3/jl/Rgs5kHvEvHE3yjJ+PBZ5X
m0ExIqyZCiC6Btr/EfcWtkYGjuBnjaU6oBSexskU3TuUfCTro8AI7tAl5N0yi7/0
A4g7FsZFH6ppjxBKxi2MkrvIdjMiF+HyrBrXoJptmfbu2RQRNPzrGJidTVPBKdQD
gOZB6Vw9JzUg+rdJGsc94vCqQQ76lOtAqOtwZ7UdqB8ArwfsdliO5m5cfkWA91iw
5BLUtJ8o1K6gJm1okE8e/lVVAt1qq+HKu0csuMlJAXtz8nmo5TXFOym9cOS3z12s
olsZ33XPRx9rmV4DXM4EgStfzlTQrr2Z3uCKdiF2zl23bm669rF8TYoqmb+nECWU
34X37I1zTo62uKrhlA/63DN33uq8Sxu7zywJpmRtQH8GY3fdY/m2ZxhB2OOty2Vp
6Y+QRb8Y6WO/EoJrjZG1Q17fXfx6odg+ADrbN9iQKFOy9N8hcVIhOKat9cknan5/
ahOthT7PKHPSVp0DgXGyYklkujuClwhISLyBWpgtBKKs9pd5kytb+rpbodWU4Z5r
+HRAJouorapr+p/Ya7pqE+FmryFrH0HzbJ6N89t5ediAp7I31DOFNIIsUqRLpuQp
uOfOKsHWvESTl8lC84djNUSD3R2UFNIxzFQJvcSBF6c1nX7yAKGMV6UNX9wKiAX3
EZv9d3zQa7vY/nx2dmZgJmEUxBdcSWm0/jXjTxO7LAf5S7OjkR+Npi6XLtIQVn7K
Lj+vPNeS2g+Bl3PC5hSJ5trsPThT8XdtlnE3PYYl+E3U49siYq6PImEzixoyKb5U
UcMOedHpmvJa6m2linxWVzfqDORFLME1twr1Q3KzNt/G692gncoYm/zLwsmyzF8F
PHwWCkcWD7wBcw8x7CQY7IrugBq6liuw6hr75x6cNfhpYZCBRNXb53yVSvntljwE
GaY4bkj9aBPU/oROYmPZ8cD9h6ScxvWRrpiv+ChyrZ9JcgPY6V+gD1uxDGt9AxLd
t6vZir0XeDq11FNBwERdeQnBD0nDSLFAIS0wtAjxxk5oJwIAU80YjqIpC8kLOcsf
QxShtwt75mATeK6B1/XhvfTsjQvRiFd1MV6eQLmc/0qFv3crT84TV3o9Mx46clUX
8JoHR7uyx57tDbjEqQ8sgbObV4yDm909hNtPAsMD8sF0hUtJtAL71lb2pxkQjbGo
D2H8rt+JXhoAPDB6Rzb6/d99BHwkKla9EJeL/wZRhzeLMLB0at4JjWMHrbD66kx6
+C1eNe4ixLmNyHmr05uW3k7wTOWEExQ1sSnQDrgynXZ+gZoUa7esZuZmnXNdu3l+
maHQtr8cGJFiPSvzrxiAZyPUs89Ev1v9WL+MSbRp7c5aMHSAxn+tQbTdTKrtbVhL
BOxOTUOUz04ZWSEeXS7qyZGSm3X9khoT8J8DhwxQPmOm1LLFKO1/lL7HAj+u4lh4
IkgdDE5WqPqm5hNDqBkwbUmH4SOfRkazbrkfRghBXzTjhKH2bjvZeyePrxpr7WbZ
FawlQiAtpSOl4KAyXwfKExGxfG7WsvWNVyajskuGvwxjjoVp2kbxDd0apY6Zr8Ay
dFQOnDSdFbk73X0npd0x74QNnW3ZH189N0Zu8y1pYyQnzE0H1EhBpOSaOY03N8v5
UtTpRpztKPhyRfQIrEvvfhatwf+LaQYxAvd6bhC9b330ne3eQq7qooA0LUFzhhB8
7AnLW6nYeVefvA+FwYI1FqzvlPP8enHS792tNhfbmMdzQ7nezcQwy9GPYUrRu3Su
Hm+SQMbZzWaoO2PDYDmR2aN4Xf6uU2nlK3MCgf7PTUnX1ty8bjlvlCsz2doKTr/l
Bi/b/A5oEt4dMvU++3PG5eSCxJ1WreirtHML596YSFLm5+OrtH9v6wH+o3YmwjGP
NWeIezobrz7aTyxAPgiyl39r5xW00CKDW9zUHgiHCUY50WQoGrupWkAksk/52fiB
GZqagzorfjtCcZf9/tfpUiiZgqOkQlILI6OqTciP/jq5hy4xOK5zJ1Wq4BF18qFh
9p3aqkTsVl3lXQRl6/VVe5wJmm1FKiXVUGqtstPyVAmd2y9Zyayox7DRmrMZCakA
OMiE5w/ltspGaiDYHI409OamrAYUB4ugK9F3h2NeT4fq+T6bCunGs8XJQN65qi0X
9sz3+3hO1h1ORlOwyRYrDANPIF5+oEGT4B7AhhfKLVXMok9ZuH/tEEne4VFcHH4g
VARkfFOWuaHfI36lW1YIgUBRRSIk1pduFcbNMxdgtLTIQKbgGTCti96X6gz5jrOA
H06fRsosE0cg6vT+WsvShc1VizKYrBUnN07KDssMCpiFOAacHN1JQ7gGOksOAdvX
tAPQiewxTYsiT35FdMX8wUN5kigkVN7FyvKp19VrXPPI7T8HeYbQtjwnh9T7AViY
P5qBWNFsrUAdVqMIos7iPgCS1V9gDQiNr/tokt5BbXmiLGuZjju4vn3JLOMivR3b
IJphMvQzFFVeme2D8q0EJ/qucwg9XlfVmLCkngLbc4w+e3p4HdtX/GQWyqlmZfkO
0+qACouEGTADYtTlpT/N29+s7t5kXPjPyGIWU8Y1q0BNKUzO+edYazSZUwoyPuvv
Mk8QboT8r8RjiwoGMX1LlP/4svvAiN2sg7rWA534iNo9Y5FRpBkHb4UGWGnN2PHX
/173csEtbV8JDa0e2erZSgcgksDBG19wG7Se63cLdVk9Z0MUgNDVbJPYju6XuDvu
aHiCrZJLpB8Y0BFYmbsRQBm0AI5DsT/xC1pYcUt3CquJKvjQGYrmQo177YbK/pZb
gZY5sqKvxs1K1c1pI2KTg3kVdWOF0rj/fwsDSvAx7D07PmQigXkQxh8MZV39a5tz
mvizPstluWOqDV58mnsn0RdzXMae/pzgA4JwYnjIDGmvbpBsOg4+1/wJXiRxjcXZ
mdH2R6y919kNh9EeVN/50cM3zHwew3/4BD+P2s0QpX6cdSXNZeg3OFNtTkNBH1XB
wgWtqvosfXujMNmjPpYg3nJyKG1QdwSonLt1+wOoX3oRQ97x3PjCIDrXmhiojaNB
KB3VfTJ7KhNoWrMUVfKirdcv3401hLCAVP1euti8E/tRNJb11QEHeX83ojWMZceZ
ITZgA2RsIQgM1jwZ/Mui9Y6bFvTckKd33SlN+hlOF6JIU+GgoD36x3DE56XD28++
s6VfBYw2U/JKeRzXUkuJwbXtsGFGQGKP5dPePJY9F5jM3MIeoRZrogau9qzJJcuE
L0bRBE1HiEEIvqaB/66xp695+4+Jx/jGJR0ssRn5UUU3a+bWbmx39rfxAjvKgbCU
kqw19vH96MUVDpr6HfN81/HaQyj5IxFgmGcne7sS6jGoGX095ajK1hrz9ZWQFLy9
m/Bs8ZFEJbNrypp0i6vJJKpQVgKfgKqtdDwa4D0daPP6au3WHLo6MVHco8o34e6V
OedhUn36AwdvmwPFPdgBaGBVJg0h50aAHxn0ceaONiiN8Bupm73wjM4yONYINT+l
ZAYuQnlLbgfQmq7sN+veUNe2oVN8ijv05Y6DT+GvhFrfgT/CC0k6G6rizf8RPX9/
Hc8umoxJt34FK+pdGJvX4u5nUFqq63m0pf6FKeWoUNrl9FAcd+Vh3sW+FkPs4u/D
aoTOzol4SCvWEEk7Rgl2GD17c7SgEPo8gMHmOMLMvlRU6ARJI4zH76A+GEMz09rY
jn4bS7WUafXsNYKNXpIpURdCkO1dKK0Abax18eO/hm0coAuqGRnFPVkWQATGpCzy
R052QqzP0uZjk8jpvLeG+rQRfbD4+CJuJOnleXdng79OIjC7rbz/0KmrU5WW8HEZ
HqWvfMGmKHqW46bQwdplJl95bcVWd9rSKaD5GQtN/QP1XQJGCsOVUE0kUaJMiAxl
iX1zGvedDeYi5WgEORwvmaKGwOLIm8uKmwBqfckFrJPvzqUFQEUg1ibgrTSOKsnf
pNcWYxA5wtL2UyammlcuOkB9aGKIutmF5eEmABIwTJnd/pN3gV9v44duzC7vYp7U
Oapuj46p1QeOSgc+kuLOUI+LNHdcpiFxT4FObLIiwgBHzLdCjXvMt/i8NCSg0his
s/pQ6zDO1jXkIlyZPV9wK4U+eoPzumCX1GvkP//GykKPHP57Ltogalz1IblPR4jR
DoVRvPPjQRnXUSSYCDZwaeRnE7Irgd+fm/YDemOH1PKqAQDhQOqBYHXlKgiS5gRt
tymfyUfGgrcpaitw/ft8nPl6J4p9sP5lHA3aG2AJGX6Aq6EaTOZPsW0DmNnyP9/Z
I++ypa7vgGHwi4pHXhK0UJKhlBm+ruO8SFTawyY1rKjNV8HJL2/OajSRsDdKfxwL
D+Qb3WgUm1IdfD0/NCRpm6njGXj6y4HGOtoujSmaQpXojei4zbGp53MOFWVgdJ38
ek5JGIhxIaCeiq3euxFQN1jSe5lKq3f3C9JH38t83Fa4pzXI0i2Dz+/27/jxXQwK
ukHCr6E/zMWpfDpAsgNEgvdrdxRj7rkMtbDjgTfVhTF18FEeEdHneSU9L/FjQfUZ
ZYG+2rdbNr52VQyscVPLk8OGZznvBlxLGfplghpZQSZN0i3+i2EzfujBp9ekTx1G
Ci2+T4VnfO96stBUK2zeXS+a8QMn5kDZYHtyPcvbbTCAd8fLxwn2Lu/T3+Yo4u3I
IX6TVK7KVQuqEJ8i9nwasKZpFuw1KdWJlEMIb4qEUclV/OGWDghFOXNlAqLl6K2a
CMM9lx7zebYP0JbJVMGuo75jAlLZhjB7/TfBX7NYRaPlWAfYHAQoFQRijfr0dQYk
vYg2YIoY0JtWcBtaOIXbRcnJTFjTdzRps/QNofekuOjUYIzR6cJ7oVjjRoVKC1mr
v0XBr6ZBeVuBblmeXZCyPG3OGd3CCbv+M1MjgI/x63sOmle1AWtWdVocHvWJ/FF0
y5cQPAzqCC+Ysm7kCiFV0ToJ5uMbY3MP7AgSIr60cAvinuKc+HM0KxjQuQRWOvvo
wclV7G/87nyBT0bpKs3TveCOqaxgEZKnpYhH9SryBtjGkprMQNBXa+RFIK10mzTp
cP/QqIF+srwKxzOr2tj2f8NUp5AQCt0vB2+oOYmkhG2vVv4DigHSjHHccF8MI6b2
qhKRfQkQ2QuQL57yaafDIBQqADjxzQEvR4JTzYbRv+9zDfeE1tI0HuSNfslpa9MI
qrFrALHd+dMCrm+32/SKHdpJNbO+Wmp4KyjFRWcqmfN+hDlNJabndVIoaOjEfNyJ
TkiW/6g/C8wRak3iP5V0dtsd+aBKNVPSRW63mtagdY/Xw7cAODa2zFi8tZZIT1Mg
jLmSAVhHQy4q7D1hOPP8Vbqt3lky0AQTR2L2FOKn2ZS/110+ltomnlXF+RLNCIvk
7gTUJvesYtCiR66sX74kHTrBYl21DkM79P1F3oqNln1yml8Ob55DbOg32qgN/TZG
H3aeprmKB3fETPKJxI6BpdXADov6oR/97SVRbGuZErE6FpVALsTMHhX/N63Q5d0P
9ARxIlnL6Etj6mx+M8W2WwEe890HCbl9IwP+AVIkVb0upcz+e0ngg6JViMdpdvEf
T7jSFHGw85VZ1zzB4yo37dWMlLDYARqkWSgiYXBueGR00lr+lJ8qB1z8SyU9eSiT
DPIKVa5T5b+akLKY9TcmfhNZCMdnL66V5/qW4G3XOyPHobWNfUs9CxArr+/VUWiq
HVFu920XgSInNQbLq52n6XceNlAD7CdIPXVxjgmID768UMGd63W92KYLUrK/F11E
2N00TA3WkM813NaG9/zzitZe3GsDUoanXxSxU6ItVo2fLUDZB3NHFXhUGJdJx44J
ODtsvN7H/wiqogBIWVIeAU0z2zp3BWH6C6rZ640bnFIhwU+3qOVfh99rQVi0CPSw
sHV5c9rTrYG74zVGcdW8LsXycgXCDWS67nV/ahykeNX9zK8hpAMKdrm/XRbEv8b/
Y1cWuui/qDe2Jsk7Xjm1ZwsRoYejpIZAz0hCbqTdwJiyPddtBkLKX+Puegjx9GuU
hJN39XcADG7WMCkaq8PXLbsJD7kYCN//ABx3YLSMV0AGjX1qK/oUiUcWpz/yfMer
CYd/LtEAcITHy+cuHPo4WEjjoRIgBirzNYEHJXVX2xnh6+coY9LDQ/n8M/NYtZ/g
1DZFROqw5BL6XbyhPBT1aDo82WuvIgTJWWDU3dVtNCqASureE7jhysVFgEKWCwgl
NsYJ2Ai8m33BnsfJeLfuraUwbyGGlSJhFTxC1SKSn1cGioXPXKQJ/QD3hGb8YXAZ
S5oWUSX+Z2byU2IiIi53HsmzUQbUqWztInJFY6IEa1dNpvRV7Y2jbj8XRdHmLEdW
GAU6lenHh6LeOntQOd0K0omF/xnQ4R5V3xmVHY9O2sTh9nR+0mGPt7QBc/cORecO
BSsSK2DjEeoGTpRA/BwQt9FaMDjQiubyiTRex0ebJijG7ukB1UFu3xBT6IrOvC83
JFy8wMr4XS6c3eE5HnMzveNQ3gT5+3K33MCmKJ9qp11t7PS23b7lAw4naqWojURo
fR1ira4++rXAK9gDc1WcgQ==
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 45040 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
4NAZGBPmQSC1EoH0Jm8NyFq7LL+I6XKWaSZYzH2Uo/uRl+mJwOGFU2bwyR/UQ7dZ
SPJ5XMUayyWPO3HKo1oVMtbquxI7WowsLxWi6wKnoVbPQOyYfg7SZ0IUiswTBg9s
KDBtRPwzE/UtBhTT7IyC7TZruXG81/AiFxvauxJCNE71WY7CC2SL/UekUcLLO6MX
rNZkX2gpNGmqxcsexeLur3asWZJDvuv+/1Vhiu73v87PpT7YU0RKsK1WkRdO5P38
HEdEOgf89lWtVOv4zzz8jdZ7A7dlhipS1HNQjKGICSc5ZfoLVZeK6sTchJJE1sBr
g6lZT4BtSogXSHQmJOUaj/V2BFOx25bi6mbG3McCk1oY0kMP7sBYd+/mCOpK24Fb
Jg9hEy/M4J2xfxCFpr5XWSRbM5cewuGE0Mxc/U30BpvwHAgv44Ot71ZbuJ6eJ1jh
QakRpGYCEnyEyFRI8GV7NjyDyUVRLlk1BjUJ+/MVD3ebl8ercj9JrNrDedP0H8MT
HFQWUKtBSgx9O5f19evTVgGYu9wkrkHoxvyrlXKxlut/D50Ame5oTPoD0GDvU11a
7hGxOuZ8hazQyGmM6jI4Ku/s8+ValGfF5aMdkuYJs21J4yimAMoRIFjiv75l8ode
kMTlVscUaye1vOKx7nwmwJ4WcAr/7XCquqXgfJ31YHP0u3hm5ae7QMtFLNs5H0bZ
rCmGDUOgzPPgIRH79GxZ0eeBoGvcpDRIB7tTrNRN8bJBMKbS8kNrEUVw6LSJXZnN
1PALQSzkKPxNZqHGyfHLeOxPHzYir4wE6WKG8hZkgkUopnRBmiblknk31vFL9mjj
qecdF0/hc9kWtGKAbjH71uefxOY/oL1qwMegeSGdjY9F9TTASZ0+C1Ct4WicNLJX
ZE5x/kDZhVFKG2KnD0XG2g3zVT77inZdhExK+A7WbPyDt0DhKrLZ5EcWv8sbDi4v
e0PIp1w8h4TwYtTAARtwJrW0nI960yuPvvd077rj56jeOerEUmQHwd448966kRqG
5fKKNg0qiNS7Lr8afb6dZ7THPTsq4utiaLA7tcA0uvHXpuw29m1rP4YAZHVs1Kz6
s0JasWvz3x4j7Lk6Xdni/sYr7eo/A//tGNTDOdXnHbI8ACQ/icgyVU7MZwNQ8bvS
9zZLLbDbaOHIA0h8u1Rfq3FYDrUSbGI4xXLBkeiQg2BYOXq60v3L6BViFWs1lpr+
QpZV4TnCjzvO2hd0VaX1Y1rlT7malEBwTA43RKUPq5wIDB9iIwCAtduvgx8rmnhL
iNmJFi5Gxgv/+PnTlQNfFznqvefx4XGJckyC/NxzXZlQa5DiZnc8dbz/NKa1Ud0n
66bVG7mgJQIcxCaZH8lb5DxIZtpWGNjXy0SEWktrKBiOXS7uVGGndMsHp3+HtgDT
RNo+aOZgELWse7EVf6mgF+2cKxdl3Ovq/Kgh373CkVPBtJyLl/s5xSxUzmVoCiEJ
vAUTbBg19bS6YuwTmQ8Wu7hqQOtrzK3i17bNJd+WfAgM71NEL1ZENJr+DvehFtlQ
inLMe4fwpEzjpVMXSm53tM0fdoYjhlOtkC7Hku8jUkbDPUvBT0bWLakXdfzgT/OO
fr18V/i0Wve4gOGSmYPxC9aeJ5+noDeYgIAMhwmdxSmdSs3mp08BNfkgqiiYNDqy
DP4k0jXiDI0iS+HcKXJYIuDbIldhE+vnpEyqVFigSU0ICloJsZyyAoEzgIi/bHw5
J4fD4aww68vJBBThZF5hkzg7kLoGHA9F0PMRJCGziqCYwfHIJxasAjM5N3kY50v/
KE6WTlfa0M2rYniRfkLR0Swk4yZU9FWWXhUM61l64XT5y/g3lxdNFvU7eb7lgGtv
M/33poP1uJQCJOl4JUP9dyhF36zhSa0twIF9qtIE+kQHf98kW/LHH2xVPCUgottV
dXImr1ZufSCrLEqtGYjqRJnOJJpzrRuJ8wlGNGuDdQtWB/bB7Eu2t+ST0+VJMOBs
n2p2xpnDCG4oujc8QbNaxbcIFeFGiiocgwOQNSGcIh3DuJSkRf7Ny6nBlQbCQnzL
paTD2PeiIOQllZ4NaFKKKpk0xt1FsP2m8zvbfcMG52xJQz81XgH7Dx0z0lOjHt9p
3r5Lio/f2Q2YRXQZWOxMvrdBfBSr8w1G6jRBacSTVq9lnP/WPf9uYDe5sRLUNESg
9yUiwtvGZ3NTcZjqfLy7mFgWQu/EgFJW+Yc4vtfG99j2iy0p+WJli5TNusWLn/4h
Ehcu66avH4ur8BqvNgYCuLhJxmKCtNEi2H5W873ArZmvOWebqIe9nK0exf+5s3RM
kYxBoDPyiwx5JCnNgxDU0A1ZPmPt6VyFcd+Ioh/cZO1HIBW5/JkCOFBGGTTG3w88
37frUGw4lfj3jKFKvbEOcDUIZVOZtIrTR1bMhWYuu4Xwpd17VghSLmvP/kHOq5Ac
yGUfBxTV0TUBf5/2xsneOVeP2ZVF5EXzNXxBlibWVmTdEHO6P4tknoY9KOF3LDfs
Z+dgTWlgK6HwiGiqVmCnLaTxsJpBg81MX/v3VdPB7QNGgVzwFnq5EjMMpBrrpVm1
oVhKDKlVxIQyKn9f9b+OEfTP2tVUJLPx8JB+EdQ4bMRyO2kVkjEoSw6rR/DULhti
Kt56Gt8QaNH1DAVe0p8uadWXiAMnIzekSWm/UsynfwZ6kXf/fTauwWKIK3GBpcbk
1xcyilKHCLhPv0Xy8bkAdwNEeFsRt6ihQy2M2ujVz5B0kAYnCmCaXhRpCfD/Gm/c
bbfH2R3oBnRYeXy3nGhSeJeoAeLGUgB+ekRXn6z44TsFcSHVFgqOO+wEseb02ZUe
ZJMI/WIwM5u986FdbVh5d1m/ei1qkSM6VZlrvY37A1zegBx5qhf4wZQaWqqLHfJw
gTAFvShQPWw6iqYSZL0fZJbx7BPdk4aIhPu+W7uZPp8Ne45jl5jdj3xXPuA5Pnq5
MyfUZfmzfWXj4MCPAA789lVDhO/G/zzunWPbHw5RnWNLdeT8Dh6bZXUtHbmkg0i9
ZGDjNUcEXye4pMOdSBorxIDsa/LNRV1YRAcY67wqkDjCf0ShRB9nFYoR+5iBT8os
4eDcfrSciNF0B7ByfTSUnmuOhoaHUvZJRY+47RAaxTgWfCulkaqiH7AkKkDb8uZD
gDsMJsAhrnlzostf8qSUkmDwQSeHYGIFXL2VzdH9B3QopGwsPZIPAGyrw+ceyC73
62jP123tMEb2qm3J6xUtoZR7vnO6GMXp2mFiCX9jR47vgwfz9LK0OIPls5eAnEvm
kCgWQilx6POWKawuow8QbNgLgWzPwkYHnkAchapvxou4SxjM212nyh4imHxEtA1J
YmLxXeX40jQV1AatW2AOu2Q+AhQT9Scwg7pkv0hxaoHqgNQ4+pGZ7mIEOO3NKUzc
2cwy1ztI5BR5CXwghPaVus5IZEWwfxjs/6c4mGHdPPtBTn1MHbgUMLsppqJvJjZD
rFaLaVB1OUwyHVACm0Ik8+GaRzr8HI6OkceOmvLt9CB8UAbf0KAwAOgqmXrrqkcP
Gjv7risbfsWFJGJFKH1yDcq3bPyaKz+PuI6PabPm23ezivA+prxPYU7E6aQ91u0g
VMv5GPjFrkuK4saGFODc1zpgAkvLtTuiMdc5YNUaHbufkWZTqAbRDKQq7pSamudz
+5nY0RRBpYBKklDD6mHFIHEFoBdntIxhydK4gTxRJAWB9E2pn0Ac0DQTFeZ30HQv
8DhKZjd7itujfs8ETtUlUPLPH3+jIy0xPktspiuAb5lJNkAtNam7TE2foXn9nS27
729BYoMfgRvuNuoa+zhegicFjxzqhhyzgktr6KwBKQlRnUQCks2Wtk3QP48piUFL
GT6jit5InCxxECTMtwpNEt1eW2DS0oVlIfrBD8Gn1BeTISV/8tlhjxfqsDgtyVRE
/Rx6ePYkv+885I15AbLTba6Sxj9z1ndMbApRUBnzse6JZuOUak1MFIEknAo6ZBPu
3zB+nGcjq3oRN9iLYj1hBTCnyEB4OlASzJFyCdtUXN0Dii5oI74hW6JVegW+DOx/
TVb6QW2IloyKQJT4RTdUCr2SFotxSdi94j4YXVi10VUvLdbp02QISsqS99qQjp1E
B6XKZje4S2Hk2bEHJDBGvuaRjzwucURmiDfNPlC0OWJ5++5U93HrI43rgkWg2Lmy
S4NHsAmnAM1Y+N7ail/8lZm46HGfv+02p8zMGX/YcoBoBixiSTUEeQocjWcPn7dn
Ccx1m+G2bfKWhvu6VbbKH4rVILLTG9l3kZ/sRvan/ZN8dpj+8oJqYHAgEOUSg8xJ
K03tW0z68xPDHZsMe/CLplN6+ahbtXDAtv0opZjfegqfqHkO41rtzLTHb2tEEXpj
iISw4vuKhIvHFT8AQ7qkoxDZxnKJidtOTXr8YIhseTI2VOq96YRF3UzZERAPsHlE
9/H7oSlW5dkoIYm/gAJ0+gHlCVl0vwQ3C4205/fuqi02T5OOzjQlwI2PxEOQPmMQ
ZbN4iKKx6uDw97dwUpWUVxBoJ2Oiv1jNqQzM34VgjdAYPv/ApFd6cxsIP8GNrPKN
K2UTJ+duKBI7sZymo1opMYYqiXBGLuOqkZuOLS648mG9xr9W7COdjJ49VvrQEFX7
g7JgqsfSJLUlgbPuKhP7ceVDsfuA5E5IRQpghIcb2VuMa3+o8Atu7vPEpWd5+hDg
LWDHf0wYnazjB52Ryst92WYmRIoVc7b6cbObXMwGsB+1Z8DizHAYd3NuvOiaY7kz
1doKm2I9Qb3Z5ntMw4hkoNKOqavd0zSgeiN3mq4Uxi9wPT9MZFT51kpkNQrHY0t7
GtjS54t2Ct/dPdhrPmqSvvruYPpruiNY5BlZhHYsiHkCG3+l0dJaetpWoWzzAnhk
emAZcmvmD+oXYBob0aPJg8wtMDA+BgYw8ceMDwog00rKMqsLFbHb90/V1ou1M378
+NJi6gYzrs6tP5uRgnNwlffpbBjOHc+bEKSKo8M783QZ+GHrXVwZxsftsQ7OxR+4
2rPZ2+w3mQzGCqmsNJLTe5ctc5lITUSHCCSxLqo3f/sQl4QCHnt3TGWHX+RJoS5s
ka/PgY8b505TY7dTYKUN9BKb41LCDZLPhaBArWa61lRrOpnVIfDioJ8k6vteno9x
5R42i39rWaAADtaVg/qyLaOUK2cZqb32cZRalIUnQrsOwU2xqvBIFOX0/Nh4UH/K
dlxwbqDIRbNjztOVu/KwgJOYwEpHaJ99Q8AFhpgpnGuoCNRNy+gxg4kHm4VJ5ZN+
8vQHiqQCcF65dxIbJsfPlBtHPtOmF+IRsiuaN4dAH0uUtRBX3iqUVvXdx3rpSszf
vOa5jJwTz9dfo3x1oy1KB1IqIU/cpMSqMNeavA7NVF2rjDsq9uHjUzShd79i5HGa
DbkWw+B9s4fSzCXnnRu6t2I2UULqFt6PxH3GVAYItbQkVT/Th06LCr6JYtJiuHzX
f+uCL66B64/EbLA0I72vuOFYlp97lra3pVgfWi2HxrNWT9XEARXYsCWm8XS6aUDc
KpI1JMIRYudq/LJuZU5QSvSv79nkZRlXFbEOih7OU1CeFLMnDdBP/7cl5SrttPR9
UtHJkA8gQcS6YLe3THJ/jn3QivnaApizyXLhUR1GaZCNurX16m8BIVe6Ity6P/nJ
H8mCTZ74ZjniQAuQdlAz3lDLpVajbRpMglX4e24m6LBBJZwdm3ulZbizhnfEklwF
ezPN6mM00xVjAcgX41xZvJggh38+q6qIVy2LG0JH3C6cJA4rdY3pfgxDQpvvkXX9
/yvWRfP2qzhGO/9yKSAoKJ2HUG5nj7X8SRQMKBFtNNFVhqxMUcPvHqcwAuizn8kM
iDV3XsuaX27pA++m7u6mY4WEsJAkEb28YS1ZIgeE8+UI/VpwuqBmhJjtgDIWD669
Hp1KEarc+PNygEp0hSvKetVaY7X626dMfgkHrikTLyHDChzI4WATqQKJdi7+trDY
O/P+Kr6Jso6yh/sNZhBYRLAGt7fhwIoOqtEfIzD/KIm1qc5ahGIGFM1deRIWxk3w
pNFjR5uhpW5DeTKyPLKTWSierTlfjbgBbqrhJaRYpeAOnNmuf3dZNDn/OvNpqqSe
aMxH7Zpn0EtiYfM/utxuVDJZlO8wd8a5LUGj0MMnzQLxT2e8/BscVSvlxdmd7WYd
LZHHGKrsiTyrrrlB/EK8hMIUM1rMwaE/NKFq2+AU/fDxCZY1JP0kcovoi9DJpjGf
yrhuzC/5COxAY5PAjA60hp/EqwQQxrV3+zegv+a3jlJRk3CIZUhbyabQfmelqmpz
KlASd9pzA4QFF/hT0WvpMbBgfxglWJMEs+2ZViRvfVMVVEjqBlIp/IX8iHBYc6C+
J/Dr2UzMq1GrkHlHhV/GVvGBYnZ4/EaH0ufIl09oeEuKviK8QWiF0kuaPBOcr4nK
EzQ4KIeO2oQ0D2uQ5vTQQ83EaTr8iZG7C/6PNKK5efc2UXDaZ5W5nrDaAlAePrwC
KDNc2W0iaCAdfbLON9Q2X7mPiggsj/Mv9P/ATuX+BszeQ4APVCgqm5Imc7IAuYPg
AnUD88qw/9Vrx698EPxz9WcHk1Tco53HfBJ7zHTPW0IpR5IX43jU1HDHRDTkTJRD
MLyD9r6ienvwKEV4ERiK+oLRPJ78fX1gvCg7f76FGYFuvBA7DRnuuwZ77B9agJy8
Ml6ucEd7LunQZe+SwJ1pIIJIGW8+y5GKQ0gOeSgfXqjlHI5QIdPy+wC/ph7PDTsV
hguxsC5m1ZQmjigTA+eb0Pu4jLxVYgqwI1sSzCcNFvpqRmUsrGw/Ya5Z9AQ1iUl+
J0b/RrOidPqenOW0paG7e4RA8dp4xGmIYcDmbApSt+u79k4OO3jaIuvhi6YnWc75
PJ4EHO2AmRUFl2ccvOtvxkjkij7smpLjJESPzNNfcMEPxT6H+8CORXDuW7+dwE3L
iyzQlpOMYaEYV0jXbsds6x6PnVKdhQe6/+nFdMiqFniJvoapLR9AlcHW5Tn0I0OU
5+sd+cFPtT+x9nqDw0kEbdDA/azOvDlK9YZCsbdWM3KV+mQP3TekTXOx48VVmT4S
TyiUBDkRBBLZpKPcjsANdaDirYIJhCh0RxZ8SNGZHzOShGoGn3H/I8TA2E8ZjV5f
c+ydo02SqoXek3kAsmfzcVBOvYWc0ILuHvzOtvaehOU2eq6wF4ecaj4B/UJdOHRZ
g3Nkj5mLC1bxwyAB84KT5pDdMI0MS1QhyU1EK8Ztol5n5DWyjq4/w39gxMd0fVIy
BVMEr50wmhCGA3511tJERXKedM6N6GLv/UXzdYleQev/mJiUj74BTd8mLg1olC1A
kDF1VLfRncCYnz+2futK19x1yxqelMofATLBiM7NSMUcL/NmSnRGX2YeZ5ihTQiC
F6BWb02VlDfT04v1SJIBHY7NyBX8LmC0uaTSrHWt9sTNEYtxkcROKeQcYk9AZxxh
r2PrOkc2CbTML7nFTUbRHk/Lx9t56cMFRHogpnUMjVudEFtEtaC2lgh1uRha/o3s
G3L9jLMa9+qMpGpwYBd+vVJv0hSJwTwfX0OfBlxpQknstRn2qFR5kbQSAKO8tDxd
II5w3hSkFTUE1ioAZzUptJxY9uGOr3EANUMZ5Of2Og/2pPENyIpy1SfJEVQJX3sm
4FJkPsSRoVgBUzwi9ND8PNNuUZhYsNjLnPCOITB9brfXbSATXOK4UExfXm6uX4pY
9rmBjUqtPM/fmPKLDz7WKU54EBSe4ce+UQmXJQqu+lxAbpYkucfr5SMOyjcOYkmN
aThrsGULKr7s34tqvWdnfDD/89zWseb+Jd4dZ4JOWJM0rMwJ/CGRyBfGHS0dSo6X
E+n4IN+HsnMVFNuClYfkFZTObMDKXo95tN1rwyowvnnnbuAVgX0vp/athyoltS/5
RGY3LPEk79UiYMZnyBjwmQiWgXPMxSytxSbnR6kGzj/p1Ywq53N4t1QxVRXrAHtQ
Rwp/VGTNKMJomvzNIo4E1C1t0Yagex97/yNO+r+FX4DlcZT0+5PmHumHjYjDK/Z9
+/lnf3h8sn0mvFSDxw/51H6bJKo/BXNLk8UTjYu2GDb0/w+vlYMm10JXC4ybwlWJ
yCDILzpMARUcLI6mnMk+MCnlI9DdaAksvw+dT+5pBIfS+QYSnqOr7GU1Kt/ALrBC
jHb282nrUdAa3Ep3AbFEEkZWTS2E1V++PieSTc1hjZoU9dNa+af5NgrS3TONOXNO
5hNNUpP+dbuNFGO+Ka4sDyyg9KKPp8obeQerpqRHQPRe2Dwr2eYHbVs/2uZ0j142
ij3AHcdXXXUqSO9B7hkPlhu94LmgvtQx4YTNqNjm/srtQ9/0Ltv70M/KgjKMRh4R
RqTTPIJ2+GfHmXTwkNKRA7ZoHoscw7liFcrDQCrJwOfvXYi8eT2Ldz+IIwyjmoUb
fkbX5liG66TpxTtUmHF7ajF6bwO9uLGcxYrw3iZEtzifnlPZuysHXslProiCJ8uk
ZW85Y5BVFwZ2gxSI0AsDw9pqpc1vu6ovcsesPfcmmaOe6S+EQs49XO0vHfCjHti/
DzNT9zsOk0HKWTWj6kRtDFHZ3FDGqkr6FuiADRC+fwoKWypvYax8Y69qI+k74l+p
A+rDZPaeIv/9aOrxmz1eP02W25OEbcagEw8Prrb2w7gZIIk8EpsShph6GT02jEM2
SZ4QuUZ2sZEdiGmTwJS6rCAiFrIrHFs0nCp1Dnta4Os/crnBiTgchp/f84USNmvF
qbGx4HKQA6vcUS3kxlZVeHzbVhjo8GeH4WONnLTS/eyzl/eJNTSsJ5DkZT+YMtxu
STClevxLRotKp4XBz8FUMmr0hMKZPn+PaYbd7WUppe5bf1okoBdSHVSXu6nriHFF
ARRkeZRyTBJ9c/xAsh6d1F15IYdZGvpA+r7MBAHSjRv/gcAf/fCABZdz5eoON2dS
x5RUoKNcq9QhtWDgI7MAN6rIp3N0+BwjjZ7NmaDw3OgP5ULJnXbHt/pkMXW3zxG+
4JDLTKFggVM/3hiiH9V56ewRmN6GprkzkpTRtF1mwqjKMFHlgWAM2hNth3jmFOHU
O9OYvOx9n+S2984/opEfC0B8VxhaUzlvFtAnYah3qs1dHi+hGS2sOKci2P0VH8Cg
wfEzpB+aPX8a6+3qNg6fFijEU7cwPesjQvZQqyw847opV53b0mgKwOND69318T+X
5O6tppviU4wNYT0UZcUxPiNrJjJkSQLdu8HyhNjTVOTmBucflOvhAgT13rErgG7r
xwBrQAc9GrK/7pFLyfOAn6Bk60NBD5KxKo85Xxsks8/BlgwhIR2BWaiHL7JsX3J+
C85byNU27SknPmleRZEGH2EF74fBlx+jxfOP0blw71n6axNJpPdRW79o9PbftxoF
uqANoofp5yAaQ16XGIxEMizBkh210zASLo0vcxN56LUqkAfqF8WqAIfnaF25rnf8
hOXq2ytr6x0qwHfXYp+tH2PUE+ayq31vhKjC5I3OeF1qabczsKX2Ch/OEWwok+H8
Lso5h0CUCeUHN0eoakFRAd49D2saaR3LDjUXO7gWW7itF3PbO5AwMFdjkMzM/eH0
TClVZ5lLqI/KWFl/0YAwJ15BLL++siMG6sQvBD/QmgYak+RWLLOvKghAGfmNApmG
HL2yTzWjzuZmFIa9bYeuASraoB9gnWGdlEs06kG67tCDFHzSJq4C0YSbyzVafSrV
VQt8XefLeAEamtUAL6DNCnklE9PzYjSQ6gs97Tto8Jvm01YPVOf/2982adHZwg5j
7BLHUdqiCQJYlhrgm2iiS0a2jcsAOiUXydy3UlZa+5fleSkf1h0IRH4+0THU5drC
qS1kL4X1ST2vDSQSIx0m5XY9GtV02avU+h8DTSw+n5mySydouLbgSQ1BhaGWLNCs
/bV8OBj4YQ0XCWu/TfP3mwtdzo3241iRZJ508L8VLWJ6Teix9KtJQIqPNr3TUsxX
wSv757YKQG0CzjByazjVD3Y5U5GZDqJ7Q4+aURsJ+82831VYpe9o3fy4HFPDRusS
K5epRJmowbPi1rsEAi7vfnuqya0g27g314DwnOb3GIZW8RtF4UslN561zncONxm/
0DdtRD/Y9Bkiu3E/kuWDuj1cqGl6/j+ZpZ7pJJKGIHV5g4dLe+H94BFz0w3XIxlM
Bh+PV0EkXQcmSyPGgRLsA7dMb9Hg8K0JLXjL78QVbLWsc7SI+Vu9SuaoyNKfiuh3
t8RLwbo8giBX+1duFFKG6QwVKGsr5V48j0eNx9RASWWKBFKkXWZIF94DfuLrlxBW
sCcsaNCwMG+kn1Q1U2zCIskH0rTAPU5s2dzohzUpvdLDvnPB+s+L9zSpvyrB3p3n
e/JMKwqQuC0JPog1Enm1TAYr3te/qqulXPT6HBoOtvBICgySt1jlktg/RWMoxQSt
3HRZO8Ukab9alsPe095hgSRpLXPPpr+0UGrcS/oRwvOgkq49bFA/HK9lHHtyOX0N
KLX/oSxDWJLkmrVdmdUPwwYgLXKnBwepGTqCPTy5P9D1vhMOJpAhslrvnCHVWG5U
jeBX+e2HHFmkoTMUbF1HBevbmOlca0Rgw3rhPqgccjBU3So8yAL1J471U0NEHJ7Y
zH8sPRd8gPmHyQh6KKdXKMkPscVSeOd3z702DPpdem+u9K2rli+1BoYLkGZMKdk7
VrcUphmLi0XgtpW6YGLTbiQTC+gZoCGG/67qNT55mD2+fBHmm7SCk0nHr2J1SDnD
X+WRMDV2GvJFdU4nqU2rit0hhbIa5VCgIjOjX58wWCvL1HvRBw2SzRPCrsLy9P++
tvVsJgq2+6cgOo+9T2kRgExWQT3V4u9BGQ7ps/jZE6sBcuTaNrRV4f/uxOeNSyJA
FIsHAGhRZ4VMyZ3zYk4fS5ZLeUphABO5BBfoN3WHjtaINHRE+iOQdHpLE9A0wE9h
BC5LRlvUaOtUA7TAfQcXemCKhrSoMHqm+PEL1ENH7N4ZL4x2CAjZaUil9qnOp814
sh17rNPC7FCcG433z1+0mWYyo1+7qZr0K4wr+vES1uGhaBeIHTXI5e6OkoOk3atY
oDuFnaPFZN+SFtS/Fgjmj2j+e3oOUBDtJu1L/ipa1xg76qpY3jVxzArX3ULwNPUf
zrc9tccmHJPEJ+4qxxH0i4Y9FyYt8Qf5Y+H4d4gV03Pc5ErJ//7Fx2pFxgGaJ1Ad
sp34j0UV2dww2HfYKopPRI0hAJDox9EzgpwXZWY4ouu5BGkiZPz/KLqcfDb8lVMk
O1GUToEURNDOqIZ4jouWIixtsbe7+FZlXnsrxKeZCxhKrukfiEjFvd0QoxzRsTlY
Ztwmasae6I4mmysDoBYS5UyjDeMD6ZZx+dO+sD7MSDm67yDylvq37VUqaUjN8DQr
MaWxR9HR0647Z6nupSUVpMXuxWS1Dgxm6sKwbdXallBndY0Fiei8xhlbHh0Yi79c
UC/GA1aPKeh4suBX0g+gy3Xj8G3qPNx1vUedH4UaJ2S1eB3lTNIlhMs2Tleqlob9
YttHb1PsiVmKWB6yjL+/wwI6IhPW6HBhydVQfOxLNkSSY6PO03QFBLkxDA50bPpj
Jb9BcIR0wlljPTrYYQonP9vRHQQkhDjwS2goV/LmPF4Btkj93QxFfp5CR68BB67r
gny178Msmmvcf70QAph1p5lAfcW5Mo8CrrGApZ8XV8r25GHEbDtLoZxP2rtafdOZ
pNkxmu7+W8kDFIQ59cMsYq4Z3yI+ZBMCx3wmfOdty9tngAGKldoMrA+OkP1CsWIJ
Y3V88PAToNFQSB0FJ4LUiChSoR+ljdgMIj+yi3ojNyR4TtQhwUShvR4s1+/qNkG4
RqeAgJEaATZGq8vndAQa69cqnOm1aewaqPP3Awtc9d5+jzKU6JTcGLWzXxCCqB/2
fZJlO6DZJbeLcWeMRnBg4oKqYrGojj0UUIVQxOrX9EqEqISKfrbo+F3t6adMTYMZ
GGGBw6n9lENGtZLstp0+9h87Y/7IGZzW92ZOHU6RticTyZIo3C5vNgqRRH+g9sp5
lcMS3sPRJc8xjAdWt3B/t2U6/ps8GjMLtKmWGEDXjGbX08uAZEOY3i4s9iR1N9/J
iV21aRx3fYSgkv53HmpJALicSvs9VPlKblTYmvSsTu1l0MCgCbGlrYwXrUGgEOwu
MmiBHy7eZkqlRpEr63lMsEkC+GaolonC9m5cNF8GFjQBG+YV9P/vLZaoqfi7ppPw
3ccgdNHFmrAZdXenkaYAmhWSwYT3q48L0W7yps0lWH+B32zmaErNLNRDZbI6ZFxw
caVbCgY71Ysq8k+f3jmmqW42G6JgVxAsTgPArmVc/h+DQ2MvBCO2D9T0H7p0GwcH
of1xwxnwfM87X9rLxKh13rISoWE5cpHt520Dnn2LJXj18Z6Xp9jRSqRCEtvfZyCI
elb0bsU0u++SILK5fskDoZg3r6ZtOyzuvE0Sq0Lbl2j6qGoi164RKPRlOcaozDcM
PaIXX+KEnOu+moZ1ZBs+FHW7Zypz/shCgFz0L+FRTntgVJPg2rQhcHO5RQadfXED
CACakQDpXN/Gu+folFRKZ2yqyUiohKlYnF18NN8Hix+dgYKmXrAQVB60C5YccZtm
3GsCu6CohVdIm+HRqxQtZ+Zdq9906nzFHGfnDOt7jnhknMx1tcvzBWNxeyEm8LLk
s8jsdRj6MT5n6Tt+5q4C69JlwS9nH+WI6hwqQRG+bxY7fXUcn+RWgXCKKM8G2GQr
T6x0I0od3d7Im8hXXDIXvIyX2P8x5HIFNpPLNrOmZUA4JbIYRB41KowlZatgHaUx
ssOgwwUFr5QFdUEjNmhuAtXeVWVb1jcD7jwGvR2piPAq3SnvpVMwO/MvSB37Q3uY
WsY3bnnSBUi0zhLyO46ZSr5pGKLuO8cjAyAZQl8VrAbUD1HXRKBxjRo3JoAplavq
dDSsaiu6/erJvVXP3HSaQKaj/MS3og4h1g5gYGOJ6G2BNK0xL1h/O7eyZldxNCnh
vA3QF62oCcOqulkcMaPjXI3XyUuPdXLWGi4rREMzr4csRIwiqVKDRI7sdAl/E206
+14Hl2XN9itx7YrI7VHbo4m4NNAfE77GxtGq16pKfGyFkEmiY+eup7hGYB+BLxlH
2Osq5AGA3r1fMk7sd/MMt4tJnfXwjfQU55f1BLYGjpHN8U5H+aCZ4s0mxyqaHjFM
e1IXyQ9SujANnFWgxeRjFEHfsuI8nNg4OXVjxvP9Y2GxRS5RBR6Ei+Ue0z+QcbzH
1qW5skz75EIJxFpqudWHnRKigSLTtjdBtmsAIwZsKlNrhcmk+Q1pIGdWo4M48YKv
jtBgzcqB5UjdrFAVKfbx/FN5QiI1JwPvBa1sD0Bf82dWmEd5UBEkrbFAEN9NeWYO
WIyzp54Okh1L351xiZrPQ62ybJSxrRpcyN5lyAYEDxD6mCRaekp4ODaEITGraPJm
+TomFSYe6OgGqVVwp7JKzwRm+Z51Y6ZHPgu2+nwto4X9XUoOLOFSo9cIc6LOjdOn
DOFF0cOxBHL6Zrb5FBn3H5zUTDowC1vX54JExH0WG48ovDTyMclPFjttyJFxeoeb
VSIIdnr1q9fjnEBTNQRuEkdcSOgaLrxWCgq44CPCO3TwmZ0ZwGIOak1O3d4yXx0p
PUeoyDcSfoQDkUNCdwD9EPKTAQk6QCvKEQ25Zdiy8x5LtuJzrWw/iYuU+MPRwGrw
g9KtGCKAnVwJIRzw2r6hJrza6lOtHrpbbU/+czflJqjZAaNAcnj5O2DKELN9m7tJ
8cVOfGGYNttL+dxKIkgWygPSQwaPq9IdMUV6S+e5GrwJahfTtBcxo1a0p8MxJaJB
wr9HYTEz+TKmXHqx7o3kmDBPmqlW5S9d8FCaMdNYh3UfPhOwzaMrPbyZZQkbr4T3
bAtiiqPHNxtik/fWDML5DizCrZ+oKKo/dnqez2ooSqeEbDhtXJuMThCODnlMXfoN
IvnwOnCUJzCUGudocRyOzK1pv6TAHRTw0W/89jXXQ7XnC2RZxPWgxtwQ08sAWtBO
5KGfEYV94g7SVEUO4vXZhZ/kocfHtNius3EitBJ/+ItsMhTUzygeAE+rE0FNHorE
C3HeBrbh7hLgY4cxmu0bU91Dr9u8Q2oVnsnGSV9Qo9a+wbR6MYWtSLkKN91V86t5
urOXEoYQO3fuTTHGi3UbBwdrDCkZcTfQUWUqpV42cmYSwXuhKx2pQXlwaJCXe4ee
C6b9yvHKYWWrYLKBJv+wZG5wm+5kRND287EDx6BFzXV9V2Hv+isP1vRBwhqZHMTc
MbYXIcXd4k+RNi5Vr3UQijhXrvOc4ENsU1L2stSop8LH4pKCkmbzFJQKZ3UlAZ9C
cHQ+sVf9cWf7jwPIcAAJtboUsYp6I7KaeRgxLHNXKrmfW8A9IvDXVHTMqADWYSYt
hkR7N6Za30tTFceQz6coHZAZ7it+ED0GYn/f8jKzmk2J0utkZaMxAozLdCbWZzJD
9qqZXE+CN40WWUb6CpfOfJm/ikfc3DMM7e1RRQo7ovU+Al6bTOAO0dOfHEjuini7
R8biYHYNPtnTsie+4arIIOTVnCpaJpVRjP6y9+/AjXtcTqjSARb+xEQTcVFja1AL
CPMePZb5mZB1jMDxh1acw2wfS3uLinH0b6wM2MWYNjDp5RQPjE2+nSD8qptJC1Qp
6OVyAzzt5eXKjOIgOH5P/4pjZ/oX2zzm2c9V5/CiFx+8wqGx1svSDhZTV5I5Hqof
RUPh9BiQ8KmaG3tOKaZqmk5uR2tPjN2/g3n/B7BzqDZhmrG//tbdbxsfDBs7Uagh
k9xZapvcN7d+/R598gZOkmxD2GUCcB6J/n6q06NUT/L4Mc96CpO7PDpwwWPn4xpV
xqhBucqSeL9CLDAT/HqpGOLxcElCdyTWUugSoQYReLtECxSdpjGkVbPFH0WyUnNi
3nbTSQ+lRfIjMoNHWQ7L/Xqqe4ONyJC9CfxdSA5g5+EeFVkQYB8/UY5UGDa/kGbP
y7jw1Y9ybWcMliKiG7O59BIO4d9juq25yD/Ge4fjb9hI8376t0/xxHBKR37r/tPq
9PqmEslNnz8Fjvruy2TH3yyOkAXc8E8SP2VABqMveWpPTFvKwLTcsGvXBrIpWXwt
PACb5YFF4UslUaE4Ta2W4oe2n4rpCPNEAQxTMiLh0J7qXuylGaI4wlicWDCrAFAI
AWe9dmkvXTSIxXs/z5G0TMmIvV42hX5NskrZPQsjvqo4nLnNPf1QQq/S4Jd3rB6x
gvQO+nM1STIffFcKaspA/oLUlsJTEcQCzAIFw6nsYTz7GGYXe9BJe+eCgy/iA+SY
cRo1dteq+AshXi8+4balP2pSycX0Qmt0+Ds1IZ7rxUelWKl3FHdpDwgPLKjlVq7c
T3cgGQ9wi8NJlxMbEX4Sg4UQO/i58e9ydtRvYI/CgODAPXKmEfv6RamLR8yncFst
o7KV0uW1wvSoDp9dGBGFlXcnHA+1z0OVg2INMfulLjbuo8xKNKfcdoh21m+JiVWI
jq1GGloxXiTsKKlMbHG+Ai54JrX4oJ1d7vE8LMwoXdS2ByyPw7HnNMSsitCdan+9
FB5U5nBnqBpajxk1rQ57iVwwK6oZBpB1s4vt6EjeDTExu37rDzHFvWdoOVDMn99S
R9vxzohQwYx21Mi/ovS99KBowOEI+jmoBY3dPGn/6VKu32v1OiYhFNncicQneazA
GedsCtp5tXfzSW6CrNsSb3pRVwITX9PtelOi8Zfix1UIWSTTRztmy6LKOoqz8jgn
nbr6ltqG8wBpCQH5ZMmc8M7PKvDHHdjS/01gZSAuXHAol6B1O1HeIjFBuF8/URBR
eAXzaqT3KnqyFNpFgdCkQpsUvRgdTShfZytA+xXz3PlQl51UKqooiv3phmS0VaOn
ZeS+bXbTtSDxoBYOf1H7sfs5ElkRSd5V58So2L2ct3K/GKkMzPG7ABynWfyyejvm
g0WdOz7uCbtEVh+KUUl9KYHvW7enIt92psyF1U+JfyUfTntdJz5ZuO2pnGtWPb9D
C5aTaNxSCrmXI4RPXJxe0sB33VGg75jM4ZD4jG1w5O82JP4KBtJiMvielo2TE9DM
OQixiKLipVL+pXgtXzwP43LI0qawjuGjRIQuS9kpD+Kui1q6Y6eJFyMA8qdS/uGm
B/8wA3RjY9dZ7T7fPBgedVlmMyXxwggxBV7cv2UmCjPYYErzx0FpVOCED+ilWxGz
n4Hi9sBARJdv5/IY/HNpkQAwHJADWu3r1Y7E2meDD1v+e8bG+w8ia6XLGHvtFz+U
nBLQ6MTu1sPx3mbLw28Ujgf6Fw4jmDT1sZ2JQqHY6g6vVlCjz1RxUBhYZO5BKmH1
BDMGbOP4at0JcLsYcA7wnNetcF3xW5yNG6jamjEDWvH5UiJQYlr2QeXTHWNRFm8I
/dkN23h7l4TSdBphpcqBcXpV9WdIl0YK6j8CYi3qmNxcauLps40lBwViKZWpwwX4
u+iVPXwUq+SYhmCXOcHNiC5o6HS4uYyFc5uuvBhnJTV9W/UmMf9TjJbW/081mgu3
6pBkkeXV2YTH9X7M7f2+bJ1pmacgrLVzkXYtK3sTkjV14kRRsrfBXF/oC4p6w6B7
mEF2Gw290BS+IsM+2WyOQP1ZhDX/jWbYQVCFG3WXS7YSUUhOBunFcNUBRYT8uR2g
PMnFS2ojGodTcoXe87559+Y9/itSs+3PdNx1kVTAx5PtljQGKNF7hy2pArE4FiQI
3v2TksB/vAiySqZ/i+khUXcLOusr9m4ugtKpv575UuPahdoI4F+wjbKsUM6pD0pG
hAwzpRZ6AZP2jEMN3OY8mwr9apSVnRtclJdoKcEVdFQJMWd0lv/S6S5CdJtzOSqJ
Fc5a8B8X4lLz2YU3jw9kvr9beU/2FKzJxJStqj+5RTpHvqJCPmU5C6iP/aGGtey+
6On9lhKsM5pl9vc9q347k0aTCPCeOO+yDPGD+D4OiKopttoWCBiYlxYU2zICKDeK
RElc9FHiyQjd5oPIfao3mN0bRBuO24r5ZLR8NW5R618zZ4DHNVyD6dDk3N7d/WWj
Flj3xHyFU1Gcl7z355n4wAUrBjSDtgEMSmK3LqldIhpVVZcjKySlZ1HMb39VlNTD
EjbIX/CV5GZYzUrbxZndXOLMPtYGrRlaFhHCDqO4IEChcolacK52OQ4mU7zu+OJt
FFEWK196bZZC6kXiQrBm5vHkF3TeNYMgjEFSdh9j8ZzFSdNA9S2nkud4tj00D2KM
fpES7A2ZmztEaJo79hgQrAR3n/Vy6HDmpfzS+M5pabYfJnVKilXWTZZN/K0+8AR1
w+KAsJYpz5s25RbfPAMO/InOqjklKIDbu5eHUcTrHhiOuPitTvkOHwdujijzDQDo
zJmxHNdRi8KuhpISzn2Sn5V0FL+v4Ndae4w2HksKTR/0bZWFEd47SvoglQ9nQy25
vkhB+Lob82hEFJW78/OAnKQnqLKGS0aQSeIMvLYXcA4Lfk16Q0Ziq1ro7TFSjo6B
Unpc5iYS4wrPBxm+mnpWcJUZ0i5VpobS76ujBQ7DfkZVerZAGuGU8JNQpozAySzg
9nsTxMcA3y78HKE9GnJ/YSLItpBc8psmm4HZPUkQ+FbD9KT7GvBR+JCZQX+l34oF
5Nn/ATQiDEuxiInJ4oyhFnF3q7k7s4ZubTc2zpW7vBN9HCSmbI42eThKYJ/Aui7U
nsm3zD2Ht+0dgfU7PZxJEXETa+0gMKAjABG2oibCrzp59dfWie8k7wcpgKwgu9A3
EE4d6yA00eY+qH+IYpuoXJvzFdYhVyfwQrIi2tOBaLKYfPmmglj+NzX4e9sxjfcU
N5vOqKz4OAMP5voo5SB+UWuG0zF3MWhLNgMBUjDc1R0wNYeegXXBZcydhZ1GGkl5
o3+ykCozDSjwUM2EA+/rg3Mb7+cni+IP4+xAE2raA/4+Z7OHledxUQpfxzLozCau
i3iG3YU5M7II2JR0UWl5ZlCq8Nh/QL7AbV+W5ELI51Nx1V7G87cRQoWEHGHZU9RR
8cC05qB8jsg/BlBgFo/vU1EuaRTh7jRIMyCl+1+0R64dckl0o/PFxqoHDBiB0RnC
kik7+gcBXVLP57HznXDRsaO9+uFiwRe5OETurFPWdnbsE5sALGybyx9zSQ3y6Kp1
eMY4hSNTK+PyMt1UPNLvTf//ri7kjzAjKlZ74hm3ezrsHrfOkOIEKkBCfF1zrU0C
cC0ob1IHKbNkSI+9kpiILGrkGg8sSBCzjF53Ydtrs7CDMDhGTCG8elmyZtrU4BPl
EJwCpVuppQ1/vJJryo3/5SQW0SZxITKJffO9rK6jvXYWQVLM3tqYnZiBywIhhsHK
tSRbP7aXd9Zv8QFKcLhtAlWhbb3jNTB69n3OOOzFWH+VwXSt/1OH7stUIfyxFKj3
vm9dXoC2N7S5eR3ZCcsKx7rWSI7a3ugbI9jeE4yH+2KxImdxfLjWdzqkKdc6jpRr
/i2JAc7gsJotgc9VfNiphJLEDJbiEJ6Un77fqgsGp981+LmFGZh6Y6x0S540vBn7
L6pFLHCVA+x5VM7GU00vfawgmgKSRyn/OTuUZHIunR8Z65CbOGD0fdfsY+gDAksA
iWkAJhA2SeIleShymnLt2jDHjvyHsjaw+g7cD0tIV0eNeCPXCwKD4MY5WQy8eXNk
Wyi4bne/3bZVNKStdnFVoYw376UQrwJwlafztmxIJoJCKIZ0JWUwDaypjoGraGL/
Uk8HdY/jGcxjzRUafB8SCgbkAMX7lNbA9pNldMzEsHfYVM0yoQQ+Yyt0Yx4kFw17
ih28HeSTV5/So462Psgm1TU3bQhBM7RYF8lc1rVj8Bf/ShhZpz0N0VFa5vOy8iMQ
/JsVky6lSvnZYwQxJaVUMoZDtfe/yYHYL8sJ1Pz+RF+UeNgyotOPNNuSPq6trZi/
tPvXCZE1WidlowfIPzLBB93iDQaI1yHJ9kLKfDpLdT+izQc4c7r+a98vdWG9rcgw
014qYNW45e28TOCAJ+xpKsC9TXwpkCKsreJbxLPf7bMWHwE9iiuo6J5gCASSul03
JfW6KwuMBF0qqc3FriCySJTJbVoZnPK4B0a9RqIbeqHS2oOMTXHpc2BfL4giLYFk
7X8pufcMdCCjkZumBA126hx04A8w6PP7sqktIqxsc5fhDRLeI7I3lVZkQ4uCXEL7
18rZl98Qgagq62G2kzClFNtDKBcs7Blf0l5lMnu4Ez6DCN7wRCe9v4NXTVcKtuoT
Lkm4pAqkvJnB0molOJbrkv9Ai3z+19j2qgDDUP85InwbsfvIDmRY2SUGbZF7fvjO
3wNycily0S8DMPsvocJBgN9G2SYSFhrSe/Low5uj5SKnDHVHonD+muPtHjfSuTVA
ttp2P0RC0mVxNEu1aLDmfb4wz3w5C0y/J3jTG58fX9qrty9OOqkMe6TJypHYs0PK
FPOLfSLh966rvE6VrUhVlVipalKvwuFbuRt6JE/K4gYqKaIoczw2DRQPzIOl2R2q
4NFgNCyNSxhcF5HehoO2zgVlz1GxGfcS5XPkqWln1UudMD+yaupE87b+IdIEPB2I
pLx/KFkzOwoN0oVv70zW6ytwjb6dkzpV2S3WNVr5m0c2yK4JYlRQ2onSOnKzshvk
q4CPCiRmGNsgpmt1q64AnjXgQfsQm/qB6no2vTD736ntCYJJmv8M+3FFeVMGd5Gb
Qm9GUNv4TH4caRSGSJBtIwPri/zcZWBAXXCL2fzcAEAvcjvIAxHIbiKJJgU4KHOr
I/SNj+oXbRF+wE7Mek+Jxv2npTzWvxNHvucbTmk1GUd3pxpeKgruPyxYGMCFJxqM
Q+8jbpKJyluSrMUkTpNg0Xw5GA57r3K0F9Q13TWUZsXIF9gYy71Ig8UVYLu6hym5
yigGyFO5Azpw/bqhrC5akIphjpcXc8k1JIS3zpS99yfLi1GwcPVI8hxJJr2svvmG
RheWPjqYyoE64sTf/L9whqIRQ2ErST1a7alrkMzaSYPGyNEvanrXRQNWvxN/Ej6J
c500NRCDfYxI2yC689Sm3GuCZHRruyxm6JEKeko4vuTMoCn++Ow2DYOEv4sBn5ah
jMk4PvP9pnJQAtidoKiN0/W34y9KEibYebcXDaXoMoQ/lTnDJ6XgglGk+VDwR+p/
1R8WGKcSoxOx+4fXZuNTiydAjqUy0/o1IgDsr+fWIQ0k3DVbxeTf8DJ0UTSXTL3O
nKrZFv8PzdQ6hNcdtM+OrV+JwGen8VBpt/HRH/EKP58McV/M1klRDE69GINRRKub
11z8YC/fzkLazQ/0WJGtAtU4L2zeauAS/8+/P1rDSBaFcVua01JY99C0MmfGI/Vs
RH+MNxo09LKPqgvCOwIY0vFSrM6zMw75YHCE0HiVXOR3OqI4y+JKE3gbKc4L6r0R
SIBksIQRLUl9YPRDkynHKRe2NwZS+8LQGgbRZFP9JlNROekrpYoQjOOceNvqPPSN
slFhQkYVCtVF0LMQb4bTYJohavnBp569UYlIIaV4UBMOMVAP6rHJSQ6tyRLbKmBY
iRGKsUc2nK42Bp3HXm/oc5Ax8kPgT16ty+Ov3bac61XhV2+Q1jJq6c8DHH/hPKEw
CfGP1GV+Q83VXCVaw0BOSibxyyQ5g9Sjmj3YVlfijFkIzMeVXSYgXcE7qZI+oiw6
SFmRvQ+JohL2yT+0CZ4oMjlAlmQw0S97kuRkbmdbt+c/A1T1gMZ+DdrrdoZgD3xw
gBbiFRDa4tSKcp+iGDZ3Ip54jZrsG71A0CJ5e3gXg83NR++qjfb9pGkLFHORolPq
rGy/LhyR3Dal9utASZ4N/Gv9H2be8CnELjrI13J7LysVxgIPIbeILzsgym6g7CZ3
uLiJUINGcYNkrS21mA/GjVdxRs5sLVwiAKd8LnDsnV9a06wzJvJAp+wLZ/qxLH8z
H62+612yWYa0qDplk3h2k1ZeyL8Ny7xByD4e+mNb5hDErNrbo7sfcTIB3RjK+a3a
pVazRjwAXZuNokZD8u4PiiN69aNnBknQktO9RIpV+Rd4cHcCoNG6g5yCC5CtjdM7
6mHtpSMQrpH0AjkOYukyBe5meT/F803fD3wQ1bMhfXPsBRWIw21bjHZ+wOBSxJZm
544wjmA/Zea0mGhwuxNF6RL0iaWmCu33n8d3NnrzPs+wlrN8nR0ClVW6QOQdPo67
FvNFAukzjjyva8LaHipBD0/HQjNjQoKSx8QggWvK/eyiTh0/ctkP3J27wH7Xw2rg
SpwYBq0UTElm3hQIQ2hIz6AvYCJoKghw4x1mGxx3UFjemP4RtYfeqNJDuCbj94mc
rEz/q4JjjTTjiwlh+JU9Ys5k68bSzTMfghYUSpI7VN/Y3JNPShZrVezKxChfWSmP
7soK0KZxPvxHpfyW+cef6g6R1xleZeNVFp6KIck7JeHNzMptYF4+3EiW2XJJq2Wq
vncJWRQrK6Y9EcmQZ+OSXmFgJF4tLqLPL0sN/5UTp715CU4pK8bvdLWYdGa4ZHVP
A6mLmlkEIzcAFZrSpgMNGCD/e9EaqkM1RsFj5T/h/F1XhpipbvQTV3xPVgxChpU4
zTwQqh1gAqljnmRc4/Klts+64LRCYDyp/+afedxloAOBvY2WLrZD1rqanYrTkqDz
BvYxq2zSbs1Mv1ncOF7x0hJ/4JhjZjCcjiIxhEFPh6QKGLwgJfCK/MRE60fzxXAY
E3COQSeza5A8s9zI/dvfRiLPCRlRqeBqCekNdFmOhxZbH6aYL04R7wz7MovafgKV
0d0M3vuYvq7a2W7pF/z5ayeerUflAC+xbCGBxWL1kckSgUIUxYm69nM4gE+u+2bM
a0tUYkZJqGIXcpJ5hGYDeyJF2ofzjPc/k9bGgwZPHVCxTUWomaPFAH3SAmZ7+eVg
cWJo10Tudk4wuyeMCJ6w+cDQgLgYg3iZKuCi1bYSmTc8liAjrgJ4Vv5JcBwNWkja
qMA+RBsuGs8974xFa21iQRbYR7XavGpYQAXsJIfJfIjMjyNueiHeIcdO4PMBFfhq
EMveSMkjLjHD2aQFnjsflFyyvDF6GFrkLwvclw25Nee2LIG8e4E+wustBwFlvGnp
IcvQ57NYqRJ33LU48932XhGI7wO9dl3uZUHwmOFcRrVjdx+hNxJkGHseL/sPHmIE
LFe0rAXDT5qbpAAeutIUoeS8GCuS8J8U+j7JKCjK16HAf27ciVb+8MHPggP0Kavr
bsxiLnmoWYyBIImpQvCLjNsUAs25DdtHms+TL0DWQ7f2CCVW5jy0u8t+YnXZMQtN
eR8eylK+pUcola2zAyJMj6A0TVj+z5ZTt0R54nFxbh2TBunB8moCSMzw3LEAb7dy
7Z+M0XYcFWSKOxEmtS8Zmjk9rqDLlAUWvXAseCDBv9zEmY+EG5Z+MdevlK+uq09k
ddrwyfmxC4ZkyRuibU4Kmj3CW4zseBeThxJ4N+DDq9GO+tzst0EK1HcMBw1dIA3e
QZbQ7VCijzGKIZkK+2TbfQY7GUs5vLUWjtfDHtlR9RnXmkUmntyWjfJmSE+UTUSm
mfh9TPk/3v8bT7qtVrt3UWfIf2Ct3mgWKiEQGo7daJHxmQDC6lSklHm/SAMYMYNk
rkFvDa6AtDq6nRlWOf9U4o1JNqPBAhalj1NMKrIlv1UBFnjYdY+UZO8J8rlldBwP
arXFY3Wq2JA+P/Hb0NzOxFW+lWb/NY8ZuFWLRCIuInXf+88ylIoefgmZI1gOhnDT
/hOXI4doumRrcCjjtqVuK82FYb6e5n/JpelubydYvtZnd0zbPOH+BtnAknOzpzKS
3mwjGpxqgcDRur5oeUgDrVo2sdkVqoIP06Vu5c7VB+KtlVgwojRlTn0+Mjq/4JAd
UsV/5L1waOovSCeIjoTwuaF/IylEw8oQbZfoVtpvVAFktNDY/9T4tn8L3KyCLiIH
+8ChLVBH2ZezYx3yL3dSNX9AY/biBBdc8aLEkDVnKjtb+dGgUcNoL1R/gRaxbxZk
FG2RUaHTCXEvbrQKfeDka4UJBVJjg6tEO/gQUUvtPzCJcSgy/tzNPTOl501GxN7j
uxw9ZaZrGcIIkjFT1ajCl1MrUDWjoTnrQGhImQIpvovEywroJeBnfelFXK9lJFDP
tUvk4qA1LmfXXnCCbqyhueLiDtYujNOjxo4Mpow5INGXNBIjRbToGS3a4G+M6mW+
5NP5ed7y0UPx9tm0iIOT6c6aDDTsPC1JoG2N9/g69FM5TnOmdjHXwrkk4aFPHcNb
bsQv/fcOplnv8FBEWOW/Agaz4xIars8GbgsjY4Ov00+u6il4ffMTNPXdJZfAVU/7
YpIko/monVAufV3iiGwc8x9QkxET9MTuf5ON7kn4Nq+NOWLAdzS2UhAOXBpdAHXu
iSzmbe6wDvAsHcPzJUICcObg93JqJ8DpZTcIRAwuAzZOkYnP3p3tL7dFCtxJg2xY
4mqKUj4/qcn66p/JhY1TX9EtdbMOmVxT/p0PdViBXDcCTlLj6xSujo/R9tq9L9eb
/oG+uxSF2g/wn4GdFnG0u1KonRYkyfFQPjNfvqt/0sLicfaJhhXKhZi0cI6+Lfgz
AFnicHVkrDN9Nk2f9+5JBwVExDIZ9rKw6/maNaIe9ihUXnEhQ7kOS0Eq+Qy/m1kL
ZCe70UtV4aDnOYVKLabMqYmoiSccIYXDFBEeuiswsu2AB5oE1TGgnKQEBXmbx9lu
98hgVn6dTN4IBoxDNvfSv/9o9bWeUSzR+hql1p/7juwc6C3N73sdZ9GESIBInpW3
uUzyllvcUYJpENX5VRtpx1dgK5tHGxEG+3hi8MBZ8QW/vyQJsIEyXdVWBFpf72OQ
vsaJlF4NVCteXTYVbTUe8FGMT/3eUH00ylNVsHrfbJtorZmpmpMd7gj54mP1Sv/V
7SUxBwp1KjHr201YFSaPRPWnszHhJkDY4TLcJYVQlv3yulgJAnF9mvWzrL8gRb+C
h8K7YD+hZwH4ron+XZhm6cL9K6j/9h3P1c0+lFtXFfdxYSfXJG2W04oOTt5fCLoK
ova1FUqDrPNg/9Nw3yRIo30Ehe/Ev0hxbZaO9LLXFvNdFNFomyCHmusUYO3nOPWX
w4O4kd584MHtWcMhPPe5ozoLUBrfY/Y35u0PL1r7idzkTx1tehnyEy2A2Q09p3/3
T/34Gpj8nkoLgwcG+uXIrTK5xECB1XU9TsvZLQe5a+5yHMvrhIBiKZpW6zehzkaC
g6hYbHr2ivtd0Q3tqdtip28WobZF/gZcRdzQ7E0pSlhMXbwybvZmkrhKr/p8j12Y
YtmPa9WZQPWHwuZsCjZebYTDQ7uV47bTxQOurTign/a4KukhpC6xhgJZkuT4ldDh
Twu8CV+HuWl8aj6rmljdUMiE2VIPuiuo+5FIOY88e6/ovN5hG2GxA4ElrRh61sQQ
GoIosveF82E94pi9J3uumtanHklwm/vjHkSdKz+DQgTkXwo2rsNyqAhc1XZcfiJI
1NnkeHEjQYZrKz1SANzYOwLp4NjtFMrmk08kMWGV7XHV/G6468omfSjJnF5ranpk
ssFIsCTDYVoMDTcj9s7AJYpyrWlHmZwGBL1rYex86Zc/YZoQa2XqmCIlDNn7OE5e
obEP80Z5kBQeKZ7b5rU8L3Uy0BQDHDyhjJyx2nKdyPR5fDnsEKX+3/sPJembPjMZ
K1PydijgXRqNJNKdaajK7mQAL/JO/niACWz9QaD8WQrzTCtohjqqqE2Izf+fr3Uy
oWMhFHMtpfV4bUzBjLiEO470KzVw9g6xs5+WH9A6VEsl0WM0k5xUKxoK8EB/5wzI
PCNw7TnH593+0K+1b3bUwggG+UnpYw+K+XV/J3k7sFAfR5VMuud+3PAnYBb4X3wz
LnXNZhZIUK0EFWQ6IooxEYPILmtdYgx8hWcUkdyCQvx9Da4UvJlJzMMxiV9Smyvl
w2T2apEYT64zB4klQHubvJRLt6+UHoUEu52/moDb1cuCxpWDLCgEuiR9F0l4muOr
f9GcWuQlLxfBGulvAyvARtocPmDA9H2wL1JEGeerd6obRTl8bi2S5rBRVPlp/Fkb
ebis+w4Ta/tJUB85VWlPrYHlHSK4JeLpKlPcZIqa8QATaHnnV5mViQuX8ttZEz/j
4j0q5nad6uNRlJBQfkCteqb6SMiKPMYcx9tPusPx7OWyZa8bCZTs3FB0wrl+6TfA
xVm4CWlS7hlqvTMH2KEepSVK68O7T30HmtaaCSWdDHJ8KaUGfZhXNreQZ+3R3CJP
Ju6w9LMQm6VgFWM2l5EddFW3kUc7pkQBK9Mq1YlwQlouoCIstEvMUE17pqwEnKJy
qFkF8/7gVkoXaMfjYw2MXs3HtOlum8Xa9cPPCtnqi/pWtCF0sQIhH9zlHGa4a5jS
pxsuVS6seRYgk3N+gdSf4E2gyJvKdGzhjdwAMFqqoa7q1OAp7jRY2YNxupPmFJL7
ISMQrvFf1fqyN0e7KE2kBvw2fTg0BNrfAnMgb47fu5YgoDQH1A7PqcSc3tPrkIay
abMzQhZc1TcxTcPk0wBSvp+fILCdvLUrevzVlRnxQEBYnR3v1FDwoM3aFrof9Ksy
laE7BGtkLjOLwwawj7OHebysLFpjRrAMjwHeKp26q74DE8nWZAvO4pX3d5Nzr1OI
p6SlwYLkt5XqXGk5dW3yBYlK55mW+PrOt0iKSEMykrlk2st1lcyQn1adLuMUm6sI
51nPRFPyds50l68u0bTh7+ZKe1SV4693kHPleCo07ow9hLJnX4rMRBafme47XRoq
KlbdiLEAXgA5ejWCabDcWyC3W0pCp5pcygoEFZfTXcPOmn+2PzbkGM+//ARGD/Hp
m5Z1l8ek81VdbLHf+iDdt0y0Mlv9IkdhLb011kYxz1051ZU8FSl5mJhXrCR22VJy
E7/mxdDazabuQc56UXjRA8hKK6F9trCeAlY93FE3q/0NxQ+3MkPHHyqAz4PsvZ96
GcXs4PJgxd0kSVZ0/Bb4BHXkCvqWr+qK2qg/MUkYemAy5hqIJKlUHGuIWmwaPcNj
oMCc7Qu0eYhaKCrL8x8r+MI+YBcS3/UHQGDVdE3Rd7/gev3o+ASNbx8wuztiN699
AHDCEzmzFMNNStUHyIstw4irgga46P2J/BiVB4rpA/R0oyHyXnVhHhmbTuLdSxa4
RJA9kzkgDKXPHMw59OJb9qkkatWv2mVf0hbZ4VUIphz2mGg8jQ8V7+oMDPM8S5yh
tnu2ZwsT2DLvdfr6VdWxzUxp77YpfHvVwX7XZqnlJMjgZbLbdu0aJOcNuhu22HZf
SctC/1US42v9OgVzA33aUAP/6oUtsDpjNGqy2xFqLSBbwX6MM8sO/5m2IY2a3kbQ
gRvYW70Jdf9AClNrmiaoZilvKYm20rJn/XB+PY5ZX4AmcfENrvfnbMnyHsz5wwY5
vP6H4V34sYFC/4IJSkPXTf0fx2a3toMltv3wD73R9JA/tOdCB0aMKYKMb/20nME1
q7SFwLZ6bRdmf68o01fsXaqtg0wN/ls+F1jQchmlr6KuNyX8jUWm9hRkfv4TDOZ1
9HcWJkscMI7u+JleIL+8xQVpkYVPcdPLYCA8RQx6Nuwy3Iy4SN1H/YCOILnrFTdp
b4Ak+Merw0Hr3Glwq64WhYQqnIQYEBPBezf/9aRZ2Hu8W8iGdvYx1ye9FfhyhhF9
GUP8wOGEQ9OGbPia5ulbWjyyLUh200qGJAZHhl0DEk6VTNoM7D5w5Ahg5JCblrj3
DZU5A3nsxC315O/A3sbfUPnbqNl/o8DIxMf3LfxyylYTrbMCVPNNjycoTQMGFopo
1V/Kn7LK6gPEdalq7HDQSGRVUROOLststJut9OnjqwK+Jifd9C8MRKa1JZCBjAR5
uNO7GPWmLyMdOrRfFc8yq0O7Sh2JgpoL7wEv+ITYLvL4X1yzevAknH1J1Kh8g5EE
UBIAgyxXylcY3RVIUUldZpdZnxPgttJR6NEMkcWVW6a5YalrNExKp8o+Ve6Ze5M4
MWOAgeygNzSmDdakLefa9BdNKeeBVLTRL+xyQzQBsZiJ9olyTNiTHzCeDY+sFmSt
7Waq8ltqfgBlfasvzUqCb7b4vS1G/+UaYs/kATaXwJZ4Ax2DfxUwBCiPlzIxjNzN
/Zcc8xzkGQpamNjjvC5s0ExCkJOjTJRKid3xcH5ebcXdxp4fzJrWoHFuKhMK1xAP
CUkY4OD7upwLyFsyULwjYLm5R6APoYlXGAjNceeJ0doraQXdL/EV4Rl+W8e4893L
Y2WI9/JDbvpYZe5mLRwhJ5r4p4rFMjVvIRNodptSAptVmH9K5LFMUerXzrgnVYJz
JbrHxFxLzzy3iCrPtTQ6UnirTwoFgPEfqLR9cK1mJldsXolv3WCEuxu35qjykiDq
3CEQV0zWxni/0grNW4X/65ANNOOjbQtjkuBJzjYf1SIa03loYk1jtl+ShShgTeUx
OrLLBb0uCrX23kBQ+TQbPUvYUsrMmE69SnuUQwrFsq04DW4OSiKPwUKDdvxlvAMb
eJtLqRz3ey85OhmNhvUmx1WRQMJ8MWySXE5qm8aGb4qHdn5XGKZXT99e/Ofyxtxb
g75UOSmxNMkglzdAzHzE9NeK67heYwU2pDlr2bgMHVo8M3ndvJO7WYHdPNRPh33C
6+0u0urD6A26ix2zCupWVTXo/paUUUhgsteMb45Y1ZJC0Pv/asHGDHCAe+TfP86u
wcUD2724MDYCNkCQIzF1kKhwH9ooUMnQGapLWkJ+5gHD367Jp/vItU373TVbyqbp
aqOIifuiqsJd45aqfsKaYLox3IV1liHecN/uwJxWlssA0olvZfO0SoAWcKB+KYVG
tjInOw+PPYB9vDGIm7tWntpD4WBRzLuOlkLPKxph4STKjN1+Hth7E2EsrfgqJbTT
TzzbrYJB3hcLCxYLsbCF7OyIeIQCuXlrEvglQHO/L+vDz3kcJeu7RWpBtgyViPAU
jqlS4YUFbQkVIRXPtKFdwwSQVIdJkg7Jb1l6TFcrisGI/lPp/pc3mAfo5CpiGrzt
MHrw+OdVV9YbM2uaeyy7zYs8CGjnsXLLZdahhbpn1oc2+CxPUGWlC2QRoxYHyc3E
TIV9cpjp3p3sWfw1ZfabnQJfTNxCy9vUlbotSasBhNw4zOcgmoiwrkdl0uA87PQd
d4py2VfvOaOHPHE7rCIX8UtEhqvjErFYDAWBtEH3ZxvCZRfv+nw0dckocr1cYff6
KG292uw7gqXrznyKTZAov8pn/5JfHmbtrR/t27XI57l0bcg2rKzxu1FlPNNjn0dr
nzyCD31cN6olC5fp4nrVFuVD2swVRBQISBpF8V+POkjTOqJSwkr5sYIb+wpCeJgA
BaoW49Cg61bVjG0hgugxmUGTM0LfJhBRrfOd33YODZhPjnneVTsFFhNJyYquJJaX
I8Iyk7PDkNdnasi3NEaOjBuUkwZpRXdJESM2+6TiGAggN86s/XC9uZ9R/Ha7onT+
UsuSF+U/X0eA5mymrsEKHPjoNJBMyQNiWtAxCTtVfj6meZiuM1+jdseeK8JQOCdr
AZ2R3f2fFA4epDgVvdibzhkGKobho4PJUM1y4iyHmcK1GctaubWhOUBR4zAm+fm8
Ngru1YPEoRM10bW85yHvomyT/3OEAqrRAjUQ174NdWMRWnVXEmvoQVv0X/byxA+N
Gi7+eCNYLO408v5A77vgKYGDzN0pTKbrqFXdxQaCQ4Fg9nNe718TmLzCvQQEcuNI
ChcsTSBZZ403IMyVAccWzx6BpKvu0GzBEhAbhe8hMEKtTc/Yd2aiTxGb2pxvAcI3
/nTHLGltucAzOa/OMmjq2Xe0JVvdMoThX745LRJxxVOP6eTczg3v2mzUE+ikBkX0
WidVzcHReEhec0JlKQdVoKUGUTbIoWWZQR64GQ3V4oFRTSTNnxYYxd1HDdaN3beT
xfXzDJWf6p5n5+FAfWlodjSE07gE8LZ9eBGtgj5Ncy7dM5N6dSz4HdGt2zFzny3k
hgdxTF/1MciyrLMYYlOC8O/1jTHqVNHk8PiuI0KQUwtfXGVnqSpMOC76mzKDMfKw
zEFIg4dffxC2+/JqoVVbZOXOYAot45QhZeEWUcnA2D3Pl7pvHikb/L11gBK4ZL5I
Ft2A3ZJWQqlyVE4ZUDP3vhvSj7WpnCDqKQBf099foODgqi8V6FE2YQGVeqSbWsG7
GgPpboH+2sIldjqL02LPYw2zDfJMd+jtuqBUXIrDkrnpVClztVJKKSb/7HQoPDNB
62EM9wflXmhh4I85aSN2zCEeWt3KCHY7qt+Ntfjgj3WC+ledO0ruqgVPteCP+BWz
HeRNAhphNf8QNEu+hI82IEy2RkgXGfZ//QuOvEJAl4XaqpUMBaXckObd67Zmn1Pw
z4xLSnt1qiT8RpwO9cTyRGE5FYJuSzUqvN0UKWrVeXm5ci/5O7cPNVgq04qrCniV
OeT98GTIIMZUo1daVA1kKgGVKzG0w/JAImHeoQmppI0XakS4YgOGkrDGc6y2D/2+
3v9ZMQw5/RbQ4RFsJ7L7tX1Z8H4A1BFVyf2xqg/cxle55+gdjummNRnUYfXhzzVV
amy9YWtvD0HjcYeqPFGZd+OYMxO+PNIFNklk68cehdlveHgokclCvgZSSqUZXND8
eVIVmbwYKGP0mybgVjVk18TuWHwNT/3iUc5rzb9UT/qha1B1tfuL7NZn6zM6+mgx
MtQoOkJC1CIehvVXptUCWbxGGBsQ7E9Os6HqIBk4TY6C3dq7Kre2CFLJcTDiVtpJ
UqOAL6/+gQWyrjwBM4xmWKIJ6jxVnZIBoReds3k4T6Z2QQ+zvsXxUZ2MfyPYEeKg
M5BtSV+yXui6TMZwYYLUEKGoiyMamrhBaZgnfYWvnJuWpws18YiM+5U6bAIBRVfI
3gAX7o3lQnVbpYlxKHdkQWe0tj4BzbuHT6jT2sATOoThIy81Y0ugLvK/BqlPDuJz
iNTwEDXTWeW0OTkIOwGFkaRT4ALFOf63nf/MOW6aX6uD+W6JVriXiqveqKgotJfH
bKWXPI+gKUCE/JToOfrHELUNsN5Z924Rf3Qzzul1LcJB/378/++rbAk0hePADhRx
ZHX7lOq8UPnxEmjtGCNhSxBjv7pXMAQX545DA/xWGnTQ6IS4Kzq1ZqoSLLvabmqt
wR7u8AmSEuId2oIKvng1Bs4PxdtvEO+4Vs6dq3/ay+mmkiBgNvBRI6I9iqpdBZt6
QtKLoEHr9CASVR2Jqse1ILWDv5FIBUIcbpjdJxSCPfWs/bmmTqw3/DccebJk/R7Z
5YhU8ksYDcv7gXvv+wRhL/INtCAj7A2VUVFToerhfhiO7G81dadlVUNw5QxqFSN2
nKXBuTmSEyx0PR1HilqRtF8I9z1uvieEL/UU6rPSkkW4q+LxsQljB2BAZc3GcfyA
hLuE4+NM7eJ3GRxfKEStPPs7li7WhYObGj1ctcjn5Yca07v1Y5Z1vA4cNyBnjGoL
WQaOkjd2F9XPAKopjzmMDq40CR5c6xgBW5QcE/2bYDVKu9IPQHesdejoRa+yAcht
9kSAWTFXc6hkBNUfLLEHmx3f4ldSrybeLlsBUgX2y/2Ea66wqxZpKBv1pSmSgp00
SUY+W0z1bFi9zrD7khtPzHHJIW63USJyyEhNgosPc3sr8rlU+0KJXqzOYHb1dxYH
tQg/3dP8+9j8NQUPS/yrU7TBzpuMmsG/jGYwhIADEKdzNyCmxzRlq3tB6rxpTX6O
WKgmx/xrcJJza0ltmzlpDO3kDrKGXxtv97bURacJSXW2r2Xa/biOAtTIUmH6nm+p
inv37DJr8HZoeMTwGSpL6LS9PtJqruNH1mZPffVWsnQN1r6hLzEj+PbXwWv1RPU2
uTfdWlnYYn5+V4OmzCgsEYPZuhAgd6CZ3DdG8gEWxImNu0LK6NMwZbSrJaEzY3hN
LrMSMur5Jo4LN1gWVRb5yH5lIbrRHlZaqa6JudTC6U9yz+cew3LCv5FxX+VlP4zx
kDyjaea+eZNMjrgWRT4UO4Qr3fCsIg04lHhWmA1kD81aDzJ31RxRGGxBp0FNoRTQ
BPtUojPhFc/J6VXjtCoarKMS3GF14P7MdzBJSJfK2M/+NL42yq2DOMahR/hgvMoo
0TA1T/B9ZBWsMC00qWccHoyCOMI81+Lj0suodS06uWTD5j3xqS4D2D5W7HC2x8wx
4+dU2FO5QWt101uoaRuqxomPAW98m1sroljYSaiEbuqmvQb4im4uJpRrxN8hYJk6
upwlQuVHNscM0m38u09uSnDpVT7PAVAysgUSCl4pzVAPyTZr4QjAgk0jbnCBhNHl
QZCAViRt1bWBoWb5GuNzFYXA7gx8nw//wLK3KcfGar6WPgIqJ+2EVQZYtgcXtW+C
RPROlwMdCOrqevTqZHq6G/OeBCqj6z3eZum3WcphXjlw84YeDHyAVyX7BwwprQuz
u62Jle0enYh4sPImRf8K76hSrYnyi0OernqQsOlax18DDyUm7YxEcGGefqvkQmpA
n9T81WEe2GhoPLTkqa5C4wdvKQU8nc0n90zwvudGaSHz4u4KGR9jeGCls4jc1aPR
gMm4il+rF86HtokolM0rt/n3DPvrFhe8ybyp9FsXpuTCmqops49Mn6Kwfu2ghWZU
xPZyVQKpsfyncZSz7m0yUIPJUMs08sEY1DfB5btvNv3EehMXjDhWKJHlSrMTpM3z
7vsw+Hr9PZlBILG2YTYrvwe82Do1fXaissXa3vRN+gDwCX15aIn/JFkUry4MDplv
LWbruBWesN6l4UiRtx8+Q+HTwWR7Ko1CpjI9xads/zeH+zkHtU3ICyB6rbR0ODHw
KVz5QinbR31J0i4BO8FtysB2zV8Uv8fzktj3fEXCEqIn2HG8WgPGgH9Lsxxd0TAh
eChhs7CfygwJ8zZQDAHrfqqeKO8Zt25cudAEqagZfSz0PYceCziSHS2el2ftGgFs
bdpX+zrytqFyR6aKO7M7BqtrtfjMZeuxHmeLDLPAefcbjjPRPKPuxa0nNFKUZbKl
tcZ71PwQVYb1bthTSpzVSYscxBw3jUE4iKS8OlQ03S0/0HIQdMX65H5H1Oz4FHuJ
StK207dJ/5FfMxLmhtdla1GL86zt8GcfzaFMrBkDUjCnjTnamwOBhI/tClPWBu63
br1SzI8cnPp4bJAcNh/qjeqUW3mRS8yIMTrn0UoRJ71mv/ATw64uxRIepE7AnM9j
RpqXGHDDRdapsn2lhm9MBhcT/QC91lJg+EXbhDspGiEn/iYgj5W+n5WSdICZ6MgS
y3D7skrkPv7j7AgoMNoWPzN970aOaj+RQimECKRClteLe3tMkpZudxsyvaJV7+Da
jRh2bkgtF3FcRUnBz5FraKZ7O9K8bHpkEo0K3BHjVuoPvlL5KblLbaimapbdHQRG
cS1Vc1lliusB+4u0c/X4/amG0VfdvwIxn1kAeFI8WPhebPOSQ3kCfLQoVg/jwppQ
CqTdRA76mNf085DT/yCzGGC+rgdJLMN+FhMfmZbvY7yYc6/h4XXhL8l5b4r93QXd
Fr2D3SNZ628CTEl7SuveXtrCwTbfdkyvRtCqNQ9/+zA2f3eXUQ6u4aFDSf79MuDj
2TCqLsqteIsiU6KheLkMO8DVjT//TK4yCNRXkUASrKS317d368z6nCFQ2vqPMB4I
gXDIVeXg2bY/Ob9uQSaMeUWM+3+Q+Z4/Y7nXhuzgmqXmiDWOb34OBigIQZ3kCZxI
GukYbsw8HQ8E0RPpAVj5B5GeHnLNbToSfotsX7GWWKrsyFIuRIkC09XC29fnEtyn
JHlNN0+STrsBzlIW65mLRg1zl9J1UxSNhtuSRh7Vcrb5lo2ir2ffHDNl1GnUHUjK
nbLaJcA2ZVOOH5m0pD86o3BhmCn317jEHizsBn6qGQfN3KCxX48o78+VbhDyQdoI
d1fxXcQFLvxrLz0gqfeL+h5zkwsppKtD5q+OBmvBI50cEsGA5t8Un+OMDeX6TvG1
8NuVphITzZ+o3hSEG+5hMNRAjR6H8OkyazbiBkUQM1gJuB/x2vLoCgG5DE/8ejvI
uMbM4vbZQ7IYE6AI1N6hh0kgIpbaduYarDhtMGnnuCAHtz1pJU5RWlPh8EbVvnU0
+XaVTPH4/tDJ7Gz6iIUKKLLb6aQI665Niq5Bp6ekmzxtVjKBaITAf4ZCtOup8p1X
uH/VnM2rkERdK6h6iiB731JuDCeJqQ+xVKRYD8FuEUEjjoowbXPvNR/cuqzMh7R5
DqmMy9aC/ZloL/x7+K87mZkVgNc4K52I+aFjRXWwoUF4ivSh/G0Xx9+zY8PMTQmC
jEbig5Lg3Dl+6tjzWTEO3UXyWdQYmSfPcbJlDGxChfpRf5D9LF+u4EJ6GVmSLZFF
3xtJgVOwf/ZFG7UEibtrSu9B9zKX5cw+SwBwD86DHIOT55SCnoo4Yw8mjtrRlB3+
O0XIGut0Bfj8f0mpxpRiy6UGLcryAUpGsV3yEOxMQbZteUpmXbTmIxrA2BElo4/R
0l8DiYFKyixq8eofPCMur2m+K9ItHfiMBYUyL2Isr5o2nl+wB3gjqkEfRqtCkC0S
2XreRCpNF/NPpiEI69xeQ+7SVNjS+oNuZD7eCW6UUSs2QpD2/YQmEvaHgyGWmcic
yDNIZ/PTBHiEQEEi7V9CmGWqByUUl0fEumB29dj5lSoefkVcChv643O9gYUgmuwz
AZSDfpfHgmeRma6kMaPLEWctw7plKiSGdm7LzDuhj4SELCoq2GouLUOWwYLtuDiM
PeF1LKXfL/SUUmXVFjcq/LhpomI3eu894Y6lBrPEJjHQdGZvr6Z10cP9yy/Nj36f
SNd5wvIH4ZB8v995zftx6nzgWOL9AWymgdrCaT03aD0MJHIV38Q7KEzND8XeLQBl
V+4NyD+Htm8q7pia8rTxgn+5RAIqSnFVIAPKl8WRuE6tJzd6Y+UT4n3kay1H8iCt
i8HPCluNv42xTszOkLX+t1pl5qjU0N0wSc8iY7xOLNg1wL23eFo3qE9biiJHr2AY
SI6rl0rkdIAXLItOBRC/1r4wHayTLaX9pM973Oi/UT6+qE29JTbeR+AuRJbptxy1
/DxJaapf4vPIO3vP3m2e0Bp38gi3gR2OGcJpP2NYB09iBpFoi+CO62xznap5FE5D
mielZuN/L4N5uTjw4ZL+FRCEhuWYFib/bP36M+EkJd9xLJ0N2Pk5JreJamVstP2U
Jlr3ykRjPcChn0r8GQCWQ10uz3Tz029PumU5+zwrup1sZt5dh8h13iTVryeY3Pz/
G1lT3tUIMR+DFfHaWYkRccVmslFMNT2WUM9V+nBHL+V7XVl9pM6e3NvpPgslmZvm
M7CFdi66ikRNkufIeoigajiBINma2saXomk2wicPtpUbxDZpd958ty3xFuve7dYT
7Cbdkk/pxpfJ+IlKY39607b5zO3Ni7ibS+gUR/hkSV3gZMaFNPSiTIRv1fQ1jQXF
T+OVp3GfNcnKJanklDYujPLwf2onwHfO6B/AF4L136n8jd38nUHNnd0zJKijFCZY
ciHYL0P4wcRy7H+4XmnGjTBv62Wf4qMbfTU1l7wF2Fci7QLxnJdejS93elRbouYi
u0yVVLQEOS7KE1cnx2E3EgF1Yi8+0twKhoD1k6cKG+BR1rlLDRtcjYtL3RARhIa0
2DGVHWKI01AWLMk4AVL6Z612boKmJD0r115xJHJycHCsKq9cHh3uQaghdC/V9aqO
mLN774vnYhrroGOZ0nOk/0y7TIPaSke4lVaMY5U67d+9qVyYD8twXDTrBAQUs80Z
oFY6gnFUcHFgThWHbtDKvMQ98RK4KejNfBRR3x5yhXAQlCwF8PaCeorlxtT3qlb7
mmlyERarCHIFy/qHOP68TuHIb0tFGyJok/qlv5hZXZc2eOJ5fh9lrxSN6ZnG94Ry
K2SKXngk6Hn1XR3kIyr4fyUt9p2wMaGI9uDjjbQaeGLFI1n5t0OM8Cebca6eMb3h
Q2p0h5elt7rWvXKsJp7nH6RHUkNdVuWggdgxYSYIUqyHrOVg/Re556HhOM1jgM2j
O6OlvxprVUEoaPzXzAhKv9tzG0GJN3nDCZQJTGZK0GBuJhVLzFK4evKYXSKOT37s
FqMEIWrb2knFewT1I/l5ostn1HM0t5ukmfPTWWG65M2RG6OSbjGZcmPRaaqkZUbv
X9l9S9rrYa7IwWGYrGAwRPsY5Pz/XZTmz6gMcEbo4F1x3Y4zlNusH/YuZh5VJGN3
B1iK/tz0REYWSQ0wtZxBgXFaLNlCHo5tlGBLO82T4so7jNTlzpuwyVX/vsDWr6eX
GdXozB4P2M94UX5D1S8B4dhonXOmiKT0eWmWMn8XhT6QRSVNFDL2C8ly9HX4BeWg
DuihR1aoxHvrhvC6lbJRe9fzjDuLlo+UpV1vfdfAlPt/bw3KC9W4xvSFbTRJdZEs
rxP8GHaimaEpbwJI0N+CL8YKA8a9Ytm6jY2MPo1HfxDaVD35hDF+dCZd88eX++sm
6q8TrFFIYMGipaVa7/XRj+vAzwVEZKQN7F4dIws0NiFA6+azbhtdo0qLfjiurjMO
QqhMKdZQmPIfzcqDuJhMHygFSjnhrqeJXsvWPv1b7R+cW+buYyzogmMV8fP9VyTP
yySS/qTYs2P/e/g0a2yrCfYt6rjZSVeKDN4ovHkLb93PpNAidxZB0aFL9fK8SPwj
nC6BV8s2Tp14hbBtU1TpLLn3t49laSFodTnrqGUp7ohwgV9u+ovDz0klopY/Nfm3
D/+mrC0G8PntpRMaPsmVripa2bizRlxq4Sf5W4PHckC7/jvMUoKiGCFQo8/4Stqj
MbhJ5HWAx0BKt/ADxCXIRzMJK40wJp2yt2+R4D03jzCmpka8cAbEieBgXHiJQrZC
X7KEFtJEtFbv+zkRRucA68vtGiDgouVQhDmcvU1ubKZLHMdTUYqjalVd72DnMUqe
Qp4TZRT2oYKilNhn+Mb7CpWq8MZt8rTkgQADu+RQe8nVqLGRbvccQhzgKIZaUXBU
DTEHAnmpbmtgjOZCeVJSJy4rRXeJb9lb2bOju+AwCsKX22BBhLkoe7zTR40f0Adm
BCttijPJhfsWNZ33y0i8g6Rq4M1WvRkkSawR8f+Cfg9liemFdg3jqa71od0ZErwt
6Gj1s9/VmrKWHQ4gyFbQ+F2+n/To/fNv/R4fmyk9LMRNs2hLe+m+xOTiG+kBan2D
Sk9v2+kZmI74Kw+XGDr9fDwDvx/nMezKqRjwdv5r/7pYiOFAiAH1/wHItUEiwtsQ
uXJmowIsVMaz5qWIG1KkNrK0C8cZYZB82vqz9+4J/hBWD08jrWUz7GqtZ5HHiCRV
vdjHDB7VHPcRxd9t4zpTadscRqHVtGjKRTG07rpuJp2BIc6bTbAq9d+LBj2h3rlc
cKgFzstQ7ingV110p0nKW4q/u89z9NajFlDZuhBSTx9zCI3nviJt0tnknHHmW27w
B1Z1+5QXQ77nNDLLqafOYjGIqe6gUeeMkajiZR5ghrdzyhAOLrYn9IOmLudLdcWd
EaJIPlYP/e+6Xp6ycj2O84qz0qAQhyUhGxiFkmukJiDTS3FbO5fWCyEeG9mThTrT
Pd0bkG2D5GhpoUBus/jz5nm5U8qUKVgmAgG+1QGtaD26WGh37hRyW/q+L8+2FRgB
31hhCb8W9T2GexLEN+anXpZYPtvl2emLE22R3pGdJPD0lI0LEAiA3HbhL4CQPJ1o
5bm4ijMeA1Dz1oHeClgW9Ztkcs0aPNUHwrvT3uhnAzUojzqaTYrlBtfg9T2Xp7II
2/ssQUaYvX6Hfvuv9heIC4ZaoZcKqlYvrBJYvhpNR00xHZ1O7yjcwibZD6LPQ/5B
hVnA2sFvAx+IjFaFHEixL6XohZY7J3WB0HmTaVzK5pnZtS+Uhf52xebNAL4QWb0e
NxS3CdH13FzWLc69u3pi9hLqGfjuAGAR+/ocHASfxY6SNAZ4CTT2IPxxiW9OQaPF
+gjk/DoaUKidvORiNpbvb5heUmVgA1k/gHrfjwVam0VxGpFXXRFdqIaTIkoHwM3L
ZETWliq7ZQxiPUt/VyTgPB7s8MZR5JL+fZ3GtZgBHKf8gIKi5e/DJkA1ApkRwRA/
wQgtVDqdoF7hjmfnff5afX8tlPpkeLg05Be/c7ySNvgIt77NoMoyNq/wpcNGd6Oi
OdK+Foa0NuEV/1sy3KrIOgLg28FCZxp3eCeHldwdXWvyKEDKpjgtJkS+0lJs/Zs+
WmhtQpYKc/Vqg4C6oUdF68uk8kjYEZDpvTXkGbZR4MKrp9GVOXvLS6E/G2PMQ4Cb
ZDvXjzArCPEM41EoqLBDWyJayOl88tGBHTtDxiaey8QXbA7xhS2MFdpWCCZMuyGy
ZOz+DwPB1F+iZz1Ifxt1OVN0onqc0XE2LRGHdHGoNGAMdKiHGLJYwnkGtwQN1yGN
VVb5GDCrQBwDlvbE2TBdvuwPX2LKHwUNj9cX87VQ6CQlG8dRnh3D0rHGgQunMt5e
u/B6BCrrIVq/K/MSeTCQlU1Vo++E9P2UrEBLvimR38AHWvxwdj27zYiifeK9kULC
Gc8C9kTZPidYRCvCWTmtTXMP+0YH0EsPC3LAZP2TdAmSVc4HVnlxrCZTjkGcOu7c
3tm6V+4tHvdpztODw7SilO4Y5Y0zAaH8bGSFeYGjQWhzGfv4bbrUIVYJSm/S4bt2
W/V01E5XczwWDLsnuV2GKn3DUpPDha3/LPkL0vNvoWwrTsUMsIXE7IbCndwEtESl
ZItqbsQitdyEoRs0YM1hLig0gU1CbX1y6pds+2dWKBMoQIGA++6BeXexPi/i4LjD
HQJnapDaR9irDZ+XpHSlkdum0tytkD8te3DLTP03vwRlh0fK9bh6QBihce04+/WN
6HjTRW98ehPCPl1l/RXDnfYsFwTK4EyT7s+hwGWquK5vkh/N3jJefQJ9UMh89rJP
7VS7uC4jBx2BErTW8KsOB1gL73qMvFk7YbQSgMNtolBw+y14q9iT2N5I8lnDJPuq
cUEuh7Lh87NcqAgDQB9Ai05VLVXLp/rZp0fIWbT9bkp1tSjIHlji14w4O/F4CASU
5ThSbHeXPll6eoctk/o2gy8VlddEmahAal2M0WRSBGgIU85OoaWrDcFUkLJUdLc6
S9y5fqpfruIBCrVIAzU294ARthrlO/mWEfVxlmQwzwU1Nrj9YyXrlZ8eTdFhKNFX
oRPHglLwAXqWClgUExF6nbn6YmcPg6scklF8NnI8MzVkw56otxYL3Mm7aPMDN3UC
KUTVfB+Sn0E1Jj93C1x85E4KMLUrAZgSNnh5vriRPAwCIbJtfAWRJhoBT6AfZksU
1cpR3ANK5vTf2KwgsgvWDz6WFuStNe4OcNlw4NTX9+eVMcXIWt0/sWifsYV1O80s
0/h8ZBigyIxG34hIeQt6PoT8PnFCYMz3LgQFzBBfJgmEQrnCITDEnnoNxdZKkBJA
rgsp9pJV3xa3lRe9upPoVlGAGmiiM6jcotr1naQZazNI6aPVxyiP6L/5DhguBuyJ
Ipk/YkUXMCcEZZP6s8URldPOKf+ZN3AWcNh+D/Zg1LdRWTJewP4VMA82nZq7vppr
N5eWaxQveOt4vQHHqGxsY/qZSHTOinq7TPsrdYhLvd6PXsV1fK3C79ZeO4HkxeyN
YaN41JC4snoAptkVuljVyWBuOlKHKz4hj2pq+xz5dwVW6A4X/eX4q4Cvi8JBNAQR
pMS0nRe/p27zge4L54EEXYWx9HLFr68PMR3Y0xMAOeYRy+PVBhrHah/ghR94fVX3
iZvXCuaQw9r6KtEyXKUAdCBy2UgKf9lE0Sdv/GIRRQ2O+ojCQctf4J8xkw2GbJbE
rPfMvuP8nyF/MDKB6dDOOv6KrVw1gnUPkpC1Dv0jWS5ANTaeXFmu9186adgnUS9m
x0YGiqBzt0ifZby9FsMMKI+6If1EvI4BTePOZfOT8GFPLFGBqydtrNntTO49kz7X
Azu5pBD+r0aJi31ondOOq6YXshrJWkZ0PSuSBLDPsHwV/EBg3/KgPo2OPNGHMb5U
bXh59eDRQpLTyxAIFvzIbZmNRHSLg1uHynVI7CRPPcLWAIF5ST7sTCceq6uhvuBK
16Rdtc1Bu7xfR11m+SD4qzVaQmDM9Xv13rZkNFXqsdMfNISf5FRYbFtA1TNIL0Yh
x57oyrua7mEfq/iSXIjd89ZRMMCMAqBN5rEX1S6K7kosanmy6gvyCacrXf6YqIPc
wtJrMkpnFJWNlML1Ew6xmsNSg1RMtT7qJ42bHReraDgeU+gZWGBmhoLLY+RA02Nt
hPzOgbko6kWcsEe9jbdXkeqsOnUk2/c5QYWDJO9ux9XUG2FGAYe7X8NY8lFlJGRH
kHONKJCksF6rGUYd1Mw2HBUDc0vHk9LOIksnPYnxggf3k3m+E30bb72iJ46SJnfP
F/1qspnMqCHpr+1aeW0N09UQakJBQEk58niE9MGexWVC9rDq4wV9N3Gf2Rp5z0ES
1t0SWQRf+OLP4/jjs7fObk7PSIy4ItZvV6KPuOTMlBkRV/ehKU1cnaJx++3/nZ78
SsRHywr2WzsvEXk1yHZ8VNdCjPDldzyCBQuyfEbA5mXiHw2n7DcGyxBY+FED6cD4
v6UjrTkmCB7h/0s/7isfmAuiWOaq9IjeFVwLnYAJp0KjwlFpCLfZUBqet20iMaMV
oxv6Xvrj4bPTmUE6Ch1FKaO2ZqnWE0Veomvak4M1u9zT1LcV5Buoz9tZ4jYci33k
d2QOEeqdKLBDZ7sKU04IrPP6EEwiX5iBTQpwWGbsDQIiBmXhlHHcoMLi9gwnN4hV
JB2nz0gWEYhnun1cNZVg0ir1FjTqDlHEXDXv5ik24p/AIIJ4m2Nj+ygraDkjAGK4
XfVmVdBwcHTUnerebWTPuwOlPjSu1fy4pXU2aQXGdaIRXrEoZaDdLg/cr62LaxN2
8RDF39C39ezY4G7ob7SQcUG8oWsXA/x5ZZg/tATclr1M+fCDELOf8RX93F9LIvBI
gOWGNHhfI2B0h13E1pUij3Ss4+wQ8LTklFjXh3UoTq8rCgNSAoqky0m687mrm5PH
JxV1WxxE1uXKw/00ymdk13iUW2RuDBgrClaXtd36wmlx0BVsENwB0UFVJFLCizGM
nIShpHEJrnVMahXC1/MuVSeXfwx2tnmR6Sxiw8xIildq9UJcXWmsv8ushzYYMWom
i9tqRL9pSsO6Y3wJFWttcmFmYPF671jrhdVEKqMDFgIKcaNnTIBlXs7hWDq5gtFH
4dI2/hM78gcaLYYvH84PPIG+q0qKvDIIpymrwcMaxuXquyfAX23wWWkUV5ssD0Xd
vofD8BDfFjIu3c0NNfgP80261Mvux0Eyif3YNCia0BQ7Qo1FaF9sVjlCzPA8MzUm
snVGVwMqGT7qQ0AdyFTpx8IRc7pHqYnnWFUMmmlBdhp7ffdBu2hD7qNNLRuomZ8c
97HOo064GdFkrok7jEXxqcqEDVwGinjjyEZaiLg2D66hMuKsmgh3RDfXhD8pgNhv
UT4pO0DWqRfSomn2lqO3mfzlDj8VnAMPr6eccsI+zAtdZj5nWLgGECBr5jBfV7tG
53cY5czNlPaGEjxim9jy9THEaF4yBem7lMtWA7rH6P1VAiagFqxKps5fMkAYMmKe
rbrqlLBlx6f99npvd0UDieZ55WxZaK1s13K+B93OwDHhgiJOhCs306nfRMLLjvnm
cXfxta3AWAU51cUCfvHfiseInCfdHipuKg9ofCkwTbp69my+kQpdEKOGG7fGODsI
Sd82fgiTU1JOxjMawIeKN0tYeNt8UZSI4JWiB3LZsVLv0VJ3hG6ZBaRkOAHtpVU4
7HCMleOphqLTyrWOf9tkSXs5IeApL770eMuWV5VF0c0hFuYkzpT6xMV9mIxRMAiS
2GvlEu7Achsh328WPUNRzanq+XvPrjt54oznLhqM61npZMkCdXW1xiVMC/1tuN3b
pIZbnI/pECrKUaGPM0JOQzR+cpS/ZGThF2N8BxWl4oqNjS1nyRpF6NkLNmU0gJm0
7jlHzWR66RH+FVNAf7BtdVNWfxEWickLH4Pl/CpYV9yR7Sx6hKdsFwOC11QbOnjh
vFktINwJLVQB/vcx6dBDNYuNUHuLWKSlyEOlcralNdnBcmaJ/zt2IgxHuDO07Qst
lcmSvrT5N+CoN5/88qeb0VVPH4N/Q2fOlu22zmwlRqXuRxvtRibZqwBSAfTMlQWA
mj0aKlr7U3PL+vsjMehtHdxv06sFJL/X5UYzDG1+Ta6IAESrdLNgIlqWbhUCMKjF
KG+XzQfAdCHV//5r1rfXaxlBo6cmRj3LHBCYSu8s0nccb0Kqui31u1oNtbI0cS4h
e5fb8EUljjAzWBWHTRj5yEOsNqYFUse8ISSPAZmYKG1ydRkGl3LfVuMAZPYJbwed
dy5rXfX9DZpRUTNcEwTVYYnAYrjf6qNIt0MQIFWsR1fB2heuF2A8gWkPg7zHR/zA
MkugV81zYT2EGOGjak2nzy1YjM/105CcVYE49upGr9BkyUIdeWWXciDuywa1T4hr
aopFvdiZORZe88aCwQLmLrS2s7/e3ysX8z78CYX4F1OmD3FCoIzWQD7svVa5oSP4
JVf/rxR/ZBVec44NbXKTsMDI3Np4LRiBtX45g9NAmzka01HxSZLStCdvSGxmKu95
d37Ky/nZQAAnroooi3CZcEjfiObJf0XENcmGALzg1E/eLCeyhTG66K2Se7gDc7Tl
6CDRrhTQajeNovdmskD3fkc+QTdWMQ0KoKjdbMLQKOjWC8wm7HGoHtE+aGgcdgCB
NDIjgUt4n3CiVEkix9qKZr+bCu1hD3ValAHDjnchIKGNy4S2Qz8mdMZcLki+kira
rMKHXvxqBbsYJTwdukHuxuD4rgwVer16UuPmwIv7WzZvSC7gRMTVvY8PQzPBZS6q
t0b4o2eq1xQAdsD1LwD77uBI6yPplfeVh8NmE3x0kNPI6HVt3tjP9swwxhqq4G89
5DmMKifNiAhFZKckep4bVg0HkKUPO3vM6y9dnZVAPbv/CpuHSi2EUxP97dqa0qkk
eIGobl+NNgY9GC3bejt9VkEb/wfdTwspGLOFcwHSlJSHlhySsvCOpsJ+POu9fIfM
h7WiXZ6k2W11tKmfnitK6496mmdbHegBYcumcrzzyi3QcU+9VF5GSu1zpP/zjBeW
3dvBtqTMLWzamjJ4csqASNQfNCnAFOsvWtGyCQtkRtUV0Sqr7AMKmMnBr8Y7NWic
6KmDeWsN+aQWGASgBbRO7gGYLAbTl0UgPq4TCD2EZT/eBZ15pNZQeYqoJ1AWLLrJ
lMIHdJwU1xHB51kO7h0YUTui8u+rE0FodR5sNlholv1oP1flBhKly8GqP4wVit/Z
Zz7guDHZ+vQ47qjHTVoJGuCcRmmkqDA6KVKMLh9K8/GUolfK2CWw7VOHDVuYTLHl
nh1fUYjEM7cexquZfwskE9ZTBMWa9AsvCMr3KrQ8OGAkcD/upQV4z4udYFuJVd1f
EgpdfY6PCV3+fJrf3qYl8dve3ddwmG+dfIl3tDI/f5n0Uy75goym45MYrSAXpCpS
em+3p3zoAxJltAVoqULU9vtZ8xjuEqiUZ719HGwRzxgQyPLHXau1zH45HQ3MFrC9
ulRstuiTnUOgLYyb6yeMMFyh79FRur4pPL6Os6CxpJUwnpjpphfZsOc5YrmWnUnU
I5f9RvX/VhWQu6/ETJCWJeCxTFrTLtRUJr72zsp2Nqa3hFjph9eeLjDybIzxP2PU
Z5JJ0isw+HMVC6ZSXUJBnn+2Agu5q0aeYi1wWW66tj2G0ipPDF6ni7L3TW5Y6xad
DfEzmf8Zi6WglYDt+B+/QMKf3ECRA8ttv0U42SvdumCacrO9o09wtWCZFVcy9Ju/
K1xAVUpCBT5busuQCEtt1vb5tlulfZikDGnaWTppgps8tL1B7KgseYd2VoQFyN1M
4w6D5shewfag2kqRCBifD6eRXsLMr/glh4Cb2WbqDptzTUwYJq/pGnVgaGWhTq1C
H8aBk/fSVlDIA0HD0LzjAvldKaXoM1MXzD1GwcqN5IysEeSaShDQXMUp0aPbaXYa
jiA70rjFzogIERQny8ry4OP8ffWWr4DXDXq+qyDfgSIT5sEU098NkvGt4xI+qo0K
wplow4bi9+Gzjce0x/RN9DZECe9UZt404muWtAeYRslSXCGxnKSB0txQEqKXUR9R
hfJeKTnSwg3H6SwM0ooN7wawJ29Ng1McPnf+ifXxEL74QVSL+S3GJbs6BQLCrQtm
1MDNWyg9XNy4O70g7iSZZEH5rpb6fE1XrTxUrdVenqumTfRCU1y6NbP9x/crcl9P
IOJ1A0tkuO0s7M8KdQk4skkR3kZlTlgKtgwooe4Xe7uyDY8ubdsegEh5pTnipvOT
5QFfHqj43E/wyFpovf1txrbNnXPERWIkNW8W/k2k+b7Yi7qqKMjwoj0OkvjWQJ3f
wNNkMG3X4CsGwYLA93Cmf/RNmIEfXs4kEvfxjJwNrEzjEa0DMPnymou36anygaYI
JVW1u2VnNh/n3WbJBWK695nQeaNihcLylEm7KgC6LFInXCspu5wznupWRUsTNG1w
fhSjLVVnC7dMXtNdfCHomDcwsPLhQiFRx1s5R42v2qkfudT+XJU29riWnshWzPNv
0xYGvhsYAjfr4kr+7f/ovxrNmGKdXGMiZIbzKPk50GCVLPXpjRwd/XrR8A06lY+Y
Xqxt8FmTnY5THXR9FyUoVyhhGnUb4ud+2tlp46Vhbq56jxnHkxBtaiZ1khFnjP+3
ZIc7lNJEtyPnW7PzzYbjxAgsuKKKRLQMBiVVKPiR6r+tU4axBeFGBiPDoXbolFuW
YztE375OuhHA+UQ7juBpOPv78cHGPLk4McoVGDf0KFkLE7KMUKCNTsPfO0nNHmMf
q+51UJn9Q5l2DKMH1PTkqk5nPUM935mANlE6cTQFv1Wj+sN7vWpEhp8sVpcgx9Li
/QTrJVmRsajHNk/IZvMD1WCbwziwqxBQst8sBa+xhvdYfabeJOwguOYNVdJh9vf6
O9eS+jLB91JVY10PgcCC9qTvlmND7+j2VM/wCoS7O3e7f7ykxq6J6Ub8cdq5v4ws
n9/gfY1S2wDy4q3l6cN8ALPtDivD5I/pXyVaeu1fSLNXWKCWJH3/nFlKsC4HEgP7
ylfJXeSXDciIS6e2B83tIBjFcn3/Bkr+cIgv5tu+fmEZvfYx2QXQemu/7VbhjGS3
FnXfQjgJfu01V66eQ/uiPaynkdrna6gutrHRKRQhiOK5lkbY2ctCghdblqP8vAoH
nGmamwzx4zxcqdg9nTDXrVhPbNQ9FlR2LsaFmpcDYKo79HMm8QDfIUn85Pdi+GEd
yWFaV0/HSdypYT6nIYvYESUouSxPNt68T9omgvbW4U5a/IGf5/2F7SdtTXObWoqn
keHMyraw9XLWBOqiH+JuQISo5vecA7J19BG85DWMsSlVUPGmtacgQAi/0dUvUyD+
ny8aHNq43S5ClU/F1oVAcA9e+pZtxSstFNJuEBP5OkfblyqiBx5bHX9h1xsMy9Pp
kMShq1sHm10cVAs6hARAQgKCkl0Bm8kwvRLLXjyC8GN/e9yui2fhixGOMognGGrH
a65hMxnAxTxME8Ih8UI1v46MSjGQbwXK9DeM28ND01qUuEmQ7vvC9A4quIe+PHTn
rcQZgMM2gdP+cFUZoXRNJE1+4f/vxD402DDnoSR+ogLnD5Bfl73i+1m2Mpj86ZTH
i67pHpl9M+E9hgSQkHeeQ32/ye2Q3ZJLUxEce+9yxUtzEkg0rI0Lkbt2ZUmOPLLF
VVRvTHCQaYc+QAUUAuAuo/JnDeYpep69N9Y8FiXq4Ds1dbzWBD1/vPgJ728d/54E
hvjWdaxphZotQVQnVaZEqF4C/6YmZ8bOnmRGM17PXKzd+N1WHbpICd30AS/B/ylk
FcXJC6s1V9peuJcdHxLo1zq6BdSFhk1c0kGCFt9A9UOV0CHn7xIARRq7mVgqYNsR
4GKV0a7GnPH2LmOO+MKP8ORlAH3qZ20P8AQXqUePL/9STO2PNAcYiMLC13qG893M
zeg9q+4xSD3+IOP6t00R6suinOWa23zDrBriHjZXVag99byTO7tXjXwrw/v5t3Ju
no+0SdXSX0l8SCzNzMLRPqMIm6uCbwNzt7kyRCn9o/KVZGbjs3Jy2A32+sQYLAn1
NZghEHCbWbd1+hAICLPi6BXPjhQ0c8ho1eP/2yRrhxke2PNfxsCHm/IY3hwifZCd
ZzzePN+PqnHCvZPQ7bvH22JhSz/+FAlk55cvfFyqGrC79w7+EmJWn+LYTm1jrs6D
QaBGjexJYbQZrPBtOseV3VeX5n4/ZkHIGP+3Hdjsfhi2xPYTnwJD8lPYmfpS9NM+
AoJueScZZn+ZYOKFe8Qsw/DImuLr8dqLd2EqKTFyBy0J5cW3/RGE8akx/TYex0TN
riOvr5fH2ih5ZkOEbIlURK3YrtPBv9J5j8ohouiiuUUbz3hKYcZa+r8LNDY+T20H
ZcHa38JJKQuthkaoMtJBH6rpibFxmSE5jvQnTm20LQf6f8w0aaWV4gKk4hTBiDhq
+mOeumQxoiH1/60Jjb1jWCJbRvpfnM9XTNOKS435WaVJFlm1mlqDrCCUHZNo+MqU
PEY74OStiIUjqoiWOPGsZUCwWetpKj8m0N1MbpnHaHD/N2IltObOF9kP54/sLdS9
BR3Kg6EEat86SwaAbwM/5UIEKiHPQdv0c1XYlUyfOM3m8XJXJgRnIJKyDJxFJD21
wEOBaDRuxJABm/n2NUCMj6cO/xrW8o/m0Ii+Qtakwy2lzQGm1FdDATHS20E9HVxo
h6WhBLG0SN2a2ws2kyf4CXQZkjaLamTJBxjNBv8ymxwiD12t1sjyKWOnEtHR9vmb
6uD2cz7n1gzHrf14LXGy5EUco9synKYQqJIq51FVrqg/NeaJhoL/dDMSpWkgYgMJ
HKzIR5ZtoHnIzTvqB0JrKUM3SLs7mWwI4XCf9y1nK5ma64+SbEEp4m6pLj1vsV4/
ASIaa6d3d+Rw8UgU/y8XhmAIRZULnOm6NcnIybWg2prJceO4zJ7+YLPfRpsWZhIW
vZE2a+tP0p+Hi0ColI6PKkRAquPYbJhEkXTUV1dFH5diaLoUj0sCYw421lbb15LZ
No2HQ+vJMAHRExE+LL+6lZ7FdVdy0GGF97b6d2THGd/G9vcE22Q2yQED4xKYyWBt
Hp/KV8ZH/mrIMwfxIRsgVUTb7T/q3t61rantsOb2R7cp4wMpmvUydPMqHs55vn34
Euy8rKfkLC6EN9G6EniTeBLGyq4UX5cxuesG9tBfbCeHga/jjGFpXM1mxwI1gG32
qvw+kOG2neBFkmGxhUkdkXPMQIh9mPGanHcx1Lg7JjVKnJisAXMjOF810J3ifUOv
3fScV2YMp7a4x84FI/M3GFWy0tPI1SeBF9avtWx6XlCKs/xrPe3MKuZ3Z4WtBgI1
0PRfwTbNdy8guLvPCAvaxS6vGWeEupE08pTbYxscZ2L6NcCFJYF+c5Kw50E+YUNN
Si5se+qCEeQMy9qRRqvAV4BPoBTytMx1319hHd4JGycwTgdGLeGQBN40hIykDQ4E
7G/F7YoxlDSeZlz+qKmxgLOIAnOFzf47RhRxLSEBIG53DuBv8kXCUy9OGU7Q8IY1
LddOVOb1ry27DD49Q4KR9/tmkOdMtpqyncTBthUzkxjbXx+7S6c6Dhk7icF1qu3g
ez7Jj2BQZ/cdDngeYNdher48cGguObp5AszlUzvZGDWgED4JVIyKdajUytJsszGj
HLXC32Lsjj0xYD2i8UYKLhHu5kW74f6lm7oM+xYtVvQpE3jxFE8HpezwuAwId6zA
3ReM3Wo0rsWTuJwawiqBLlAm3zurpx2XdC/vZywWy21va3+8Rnxuq75tGXHtbfb3
++Oh2pm9kp2nMBB91IiMNMkkL4/YnvZQFohnSmlplhzTzD80mjCeaLltYhSkqYpt
2FW6HHF+zX4sEDyWA0ILMte/RbZTByEt5EKPd02QC4hQBIRAjDGZ3JfslfndPbNr
QKV0e4Ruev/Dot/rT78ZWhaY1KxB4bHuW7dBqaHn0/Pf4AAAazrUuWJO1HlTAU/P
Bk7kazEvliGN3NAnp5yIkMsav3ezYcG1dNkxt4YYrKzVnnsF1O6yZs7zBB3rWIwG
4/kpOG7ciTkXiIZ5NV4HXQFPtY7xZrdZPssmqUYEJLC8B+23oMrKil722o8Miqw7
b13EQ3aP9lb7xQ53UvtC5ml2yOtkp/faDKoJfBTADT72cZsOBwMc8xwNw2QWKlrm
uIhLVVbBtN4gJqve1Q85I2We+DXMPdP8nlEW/aeQ1Z7jc1JeI2mFAvRI2YTnkF4+
AH2wP54m+A88WtFA+F40FSNtTOXNannX8Sr4NJVwtSP0FQ/g4aTLElogjRUXwe9b
IP9uhw9qK09jfYCZ4CzSi3B3yY+qMkJkPPpwzc10CYsmma9kt2VhSGGB50xw83+B
n4qFi5SQBJCM2RcW18szWebtaqOB2FJDkzJmDJi58zGLaVtHzmhT4dvF1pUdHNZ+
TDZjMbpEaXK4Q80bCkn81U2g2QI74UTippsI8EnhNgqFTYQVc79SwKIQTs++QHz2
b96GFTZWtCpv6bVQG9d5OmOaQtE9+k4VhBGcTRrsuDtesx51F4T4HhvyjbvWjyoE
lkfUdv61GvZgqEZNIDXLg1umbhsau9jwtNNg3kIfc9oaB4VM1+Gt+KdV0TgK4fPb
LLHJJrehNkvrykAZ24n+snvspwVDH+b+fTl8rkiiv18thRkOnLIf/adw5Tcer742
u9qQ8unFAqQiqOcvU880zV6PmFExNYRVQa0EI2SsfVvPBCSc4TgVEIuhooapIM9W
o1Efgrc5koCdofl0UxIqNBx9YGjHlB3TzqDGcyFQru8tmuYWzoZosb3I5g3MBvTq
jUOBnB/P7L8aKIoiiF8ilH31G30Ct50r/ORUi1r1pef2jk4sjEPb630Cfn5GhRqO
m2PTkE0o4NJQbKmtG5NF7Pr1vHetJMIH3usOIR45zdg/GqCZtwyg1Pp8YRgHNvEi
246/wlBM7s0McSj4hTUujqekyK60lf0Q4ssNnCA52NuVNmvu7wOxxtqNusujWebD
UMkKqrhG81tsQ/AgzBEe7x6mBuDR0EVUVmCIKO3KF1U3IreGbVsbj3SmuLuIKsGj
UU9h041z+LLkPCvNDnhQAlg9UrRq2WA3aeY1tRfb8K6TI+aHyROCLAiSShFQFyLP
cGMyXu+vfF5I82tfXNgJUOv41n/EpbIdNdKSiIORoOryNz0LjwPNo3H1nJ43Jacm
LfzctsUxTWNBTUfp9q435C8O1d5fMI4fiNLL1USM+rjXfhkUKZ9+71+stBfHOtIm
UB1SmV022tflqDmNk7URI4GPGVoSy8CI1s4mArxnwnpjT85HtcQb8RgfbGbK12jF
YwEaJgxzIfCCqbJVYilFBAjWEeFBwWfegLPE1RAjqjHAIVym7eLS8Z+fzB96caY4
3l2sHYVNM2P/b9wf3Id7U76U90gQkjO9ZwRiHot/Xl8RR2MqjlZFsi/I/89N+V1s
47R6sc4sl7IdBFwhk6LFB+LqSdjGGus8ivN3ydQbfYJs91+lyxFkDJIvlwXOKBMh
1YC5WVNAuBGNlgx/DvZ3Efv0KGw2P6hAg8SDytW9E1SX6sqzBRzPNbH7uqVwXRv5
TAVV90HHdqgpuNWaIPHgo/znbZD2xOjVJZ9SqAZb/3lne09WZiKXBMm30C7RHyih
sCMgEFarZTTvZ4WOnmip/b/csnJo7iWlR6YLAHuMDfWd4kFejQaGW+dhHkpeyqHB
cT/Y6zKmLKGo5vuWXOC/3/qFkecFvoOfQqcu/KF/abX4OMnURyVi8AAY99MDcWCQ
ak8fGzJtkXLf/bxUPkelMejMqgRT30VBoRDkG0OOqL4OTnbcqflI3Mees/73QCzx
ncrwx/pSavx5MqcZ4ClGmY4hz1cG7nPn8+XSvJzN/Kz0OrKvf/ETXTM3Fne+AnJG
k3YzNGhX5zQlkLpZvhr8OaNP/0A/r8gm2bFvEVwbW+kmGBoOYe3QJg275TY85Hns
CG15mwJ2cIoK5ji33AFtK1zTcaLmsLsFTh5rV1tUUmLREGSWkQJrU4+Bk6M7fRGi
wYru0IJie6pTJt1xo21un/RvsJfEC5p4APqKzGFel4bFOGMZ2S+XowgGgrzFCIcq
AoC13wITWB+pHhgUtYYWo9x6kPZWtWdf3BlmPrQrsxWxcpwwbg8VUUkwHp0sZ5FO
vJtRqspGFHqS46XpYPrXKL7LAza2m68O6I/J5Kr/g8VOgq5JLbGJpm6wwbMCcQa7
iGTTJQ6iEHia6zcnEz7gcqr4BCF5qvj39BDPOZKqhFTU1wpCqaXL+35RsUMnHCBl
T8UbJ5S9kpdMdf7OaFv8U3GEXHa498pnFvlTL9h6CiFCsufJsrDZDxqEs1r6HRM1
yjX0BPpsNvHe5g2LuPw34+hYGI+KkTWIC+DMt2opEGc16ZbkCulUdQ39O0BpL8+e
iKzwQ/CVFgmZ9JI7HVo1fKEveLU4y8CMtCPwUQllBG+yusWVXhTrky4QHlQl3Xk+
DVKUjenNPBtW19VEOKAWyTl1KFAOztNHEwOjU8VSmHcbqzyXv/HMlHQ5ZWwPAXcB
59D5b8nhUBHK2c3IgujHWIlKrmLKPj3NB7meNNIjgagVSXbJLkCO5aL9wspdVySI
etvETzdUnfZ+KUPznz2eIs3OrSKakFdXKgmrI0bp5ZxseGeMzNRYPdCoULDmTXBo
NcHNqkdZ2ykL7Bt8lxR5Z1ipyv7JhoTxJ09b3NFpg3tBrmbTPYHD20hWGyLW/Hsa
tstoj0G/sOHKXRrQsqmaf0cVlhAYh+rn2IPO6LgHKxcVTJnp6vKyy6WVGOXUBGd1
p6XFedi5XQrBZsU2WGE07pw2FpKa78c6v8kUB475wKeNz/odAZ9KusxEKgu/AZzt
iYMJlvgkKDPUufLaJgZ/8O8hdu7UwsIK0VVKzPIIUKlpHPD2C/vwWsmVLZgYEhzr
xU4H6WoLEmAyOvjFrlBT+yXXdXe5V7hnDl+nuV+ujZ++n4PiN7NN7uwACyEpRkA6
Wr90Qf/7C8qJ2tHZlOvaA4qLrZ9JVXokNL3+U7HqeFyNCgutPW1H45GYnzk6fxdF
nD8BRVSNZPwVzi+HPNjBHMH/wkDwGICXWI4XKfnuvd//tQQRxOESCHsaqSa5dau9
Tc8vSItXl0kdv3nIdAc3U/eAQcn5aztFAnMgNjD/YZJ0JB/XZuQWiiEuaYIk4rzQ
7xjnhteBIHrzD3RCtq9UkydhLFwIMsVFNnETFjB8wxyDbRyQJFsuCdf/XWaoMdUy
Q/go7Rkc346uZZUxX1SEJ2HWWFuUCUsAda9rlT3BUtdQRnc/a0k0Mt38rkrWVeeR
u0I4qG8XHl3zzvYNB1mBecsRqsajI7SJiu/dQgbM1STMaTnWAVHDUMpj7BUEoVIN
k6S9Iu+bdXa19SWbYO6vrKfbLIBOZCeFwvtvhz+yYaPW6FcpjMtu8TvOPbSV/YJ4
Y6SWZY4aP++GhOzE5ih8eyg1rdYGMh56NruSaN0K8pgOTJN31y+ovLkNl7apYnRa
+3HQpXKIWX3+0U7ii9VujHCsSjjhSYkba6SNriu6i6xm4fS/18Fk6qrz+0ikbjBt
qzTOQOF+iP1b0vBWdalqLMruiBekGwGCni6z4tJEZXkXjQ/SYeyu0tEBGy0E97br
14sALysR5xvExSAVAwE/XpYE0B1c2AZJa07cU7yEPLeXYa3WcvWyBtDipWKPEaXC
L4XJeW9weCqLt3JYygt9rW4C2gyM507Xu8OLxU1uXLeQV9jRwvShcOWwV1ZsG9YE
xPR2ecXrDk3CEp/dwsxCU9PrNq9/np4u3fz+haDIweKSt84Yo5qyEy8hsTi2sIRc
s2xEQZLTmCiI9dYi4z1knODhkjpFjIiicgRQ9OaNEX8jJ/Q6LSaBUBxzttBxmcOK
dQraL1te6j4zsCfXPL8FLD/Ap6YReYaR039GUvjxZ2m+0hIWokuqmUvJTPjgpIlA
Ah/5ccKWT1rnCbaDILd95ztqWapA0IdouDwBJtYZHTziwEyGSZ4JnFJB7f3slt+o
h63i8etuNb1HjbNA9X9O7Y0AYxvpYZ6yWGi7Vb4Yanw/a1QTQaFEyE3K40y+WyVE
kQf7nMdTWf/R9TBMmSLu6QUtIbKzkgfhWCxf4m6sR1ovgyB0xKNlT3jmSFQ/2xQP
g0oqaQWZ62J83UvB2QXFhI890FGrJ8X3NI8wUForLBQanTSQ8iRYnKoiVpEbwS79
jQWmN/NdGCPF6jkBXJtgVGS+vDtljCpFQkoHygAX66MdVFs2g6XvWFWqk9K+8EB/
ABKskbeXf8XxUeW9blLECGKe/ryaw1WnN1hUbh2SiL6l4Qy52b4J1AujmuzYydJn
IHogk6bqatpljA+3phV4mP+YGuJJmB8KXh0MLPwlDS/VplqxUAx9LJJ3KkQdD42G
aAJDNI554ABLm0bKZO+TM6kpc6s8S/3R9PXHcMbOFxaoyRgjfWoRpOPCa222md8W
kcPi4LpHyQnnmAXoJxtjm7eKDQo7CZ49q4F37zNk8EHS9Nund1+3PcvIQySRoSW3
rGV9VHbZew3AZRAxc/jD42RPV62gWFqYbWnBWVnDFZc2NT9sLsscHkpRb2kK94YZ
eEH/oL10wTjNHDEB+hUkEulMbdf8F5G/DxP2LbpBiBTVVcZYm2ZwtJgvVl1J+ZMY
i6d3v/6iVvV1DbZTilliqfCY9UHn8kCKMfrNZO5lbJ0CPQgtwfazDTeu6LQqdxSG
N6/BshgpV56j/BUcnZX9wUY51hwSkvprsjqiJ5EwKapQzRduakNYfth+7gBx1Fff
3h5G3RrUxsLrb/t+P2Znhp0tlMhflMdURsDNX2Dhsa4ClNEyqws0RM1IjLR3ljR7
iF97NQLWja+CuHxcfSy94EoFo30qrRLsQIMntxJ0TDVJZVBtTiK/z6TbzIP7hPt8
psdopkA/+2o+i2bV2NqY2JPNpHKa5GSexSftvUp2iomWwMr+rutL4KCL6c+wcHMG
GHla0RMNrpFV76Gj3smyHqbSG+X8QEjUB+gtnHRMQaMZ/gOEwkthXfUQDzo990nZ
jvTjUH6bMrNXypESxAPrrM5nwmOj5s32STySv7nBxbNyo6aN66RmxMhryudwnDuT
xSHOGD8YTkRx4xM0+3MPHMnuOhS9OmC/wru44By/CtER7aGHyXvVqe3KqFbBTC+k
/d4yoxJOQ2Jjegk4kJB9wXPIQk3SxghVscMFKY/Nxiyap3f+p4zCgxcFHt75JOeb
cBgfZtDWGru5SidL+CjvTwjS7L2ewwXPZttlRSiGpWCiSVc38+qfbrnmKesdKTyv
vwXrmzgWCxxjXdP00dw1rERRtj7IRcRsxdp2T1PDuVV7qnJP7nTWvitAyqoX6YOc
SytA1BAS7mUnk4tQboet3VrIJ9XRZooOHQNnJ7ldHCp5thu6PhLnEM14ifL6ABOw
eujIyt2CF5LjAzxH6kwn7rbBZ1iwvl3NZcLfDy+lNO5Tw8f1/KAADPx10To0itDs
C2RyWCaHejlPTC1LAch8JQeASocB5rYVsvw7YqwbQ1FaFs54rgNM0Ng3d2F1dfKS
eTJFO+pAHROeB40dnCKcR8pwufW32Jf7UAeh/yKXKeFi6fTKliyTBX8mVctRpyc+
gA6mzZnARkkKx5xvHF7PXDG7iDiFpazieS8pIbqTbzIctb1BHhnWAKUtcggEoEeM
XlUODpBlnj3tROVOaeUzPXgAQFiUG/WXccE5qqO6T2ZN3UjkszIWL6QC3akF7u5x
ejUdrwqLvsXFQewl5o+tzFKcmAzvCuhELih/QYWMbiemmOjfu2AFiMvyUhSHF3uU
IEM+PIgObpeV28f+KQhF8Eru0vq+X2pPuF7toxWEO5zyABCOcLoM2ggY2/797ToB
RP3T8eJjWvtlZOVV9VgqvjW1hytKlMVd/44Ezirp9YSlyblkbqIxa1pLLimZZtIq
O3rK0+zOQWVEFK/rsLAT8uNr5YbDaGN1U+BmuijQLHA1AZvPJe3kNozygU1V3zs6
i70CK95nmYiTkGC/1OWFg2N5uIwfysuG8frE8dN4IPdcjWP2sk1qrOEWa/UX8RUj
CXuxouZ/uuq78UwPxSpWP9nN25E4qvBLtrTi2WiLnJU55YXjui1Xs7HZvI+wcmQK
35tVMpdYpWnKDgqQFdHNUcMpdVqtMrPBL49nrr9uXAvt4auYphAvJwm9sThfEHV9
gfGCvucvRtDImq3ksAtEfNI4WJT+77YUiWtKI4G9TM7pw9yuNqC1+b/dqwU12Gdz
NWRKGpO7HYAYqrWJUCSuaKKMDmJnweGn+e9clAD3XUEH8NdLlS6v2AFlxMbc+vjU
f9RgFTWBXLUOfKxTDUjiMqXDU5WsEDYMJv+lKs1sQLbaz+9pOmD1NFPzWZyRBX/Q
GFo8P2h5LP9oh9Imb+drBOTfewIa1xO1ZEOdH0CLUsIw1v+ZFEV3/K9ACSzKe/lW
+l0dc3/46SoxoKQj6Bi6Sk+d60gIDiVR7g8WRlJWSeVWlJrNszJnoYkibPeaN5/A
J8v0fnTxlAcAzMRVwcWgzHUWaIK30vuN978WFljjelk7AzSvfsGYrHOpWpc47VDs
v+Yxjkf1ikyHEo4JIo4BNA6lwdz0GjLRX2VjbaCvhmZKRmtHeft1vAIrCeBRVDwQ
Mf1uCh1EmN1eabJjyA9aUX0BBHCQYZ0AtU/o0QxwlvP6bFvnvMPTrF/VjOTl9jZ7
J6rejbLXGbmLadL8BC5tWrGQtqyCJMzG4RE/xU8M8jrydmHMlLPL4i0pDrZtmREe
NvoiHle2MbC7AQEzIOFyHpBTYq0ZO3LxS06aIHdEU7UYEiZgILwgtIMLc/F1iEPW
pckX1tjmih5BHIhHLOFMe+vfu2tyZziyxxtpMq0x/JYhw0XIJCPvXwLu9lBWcvBG
mm/cTK6hzzkWjkRuDUqlViSgBXSVfn+wFl1ozyFsqoGbubNh7M1vCdLFrpgd7eSd
xf3fNTajtBbjb6CzgfCMzgz6d/OfuGkQQHQvjQ2eSh7Njjkc2+R5yTz4IRa+bn2I
uPcGsXYGdyGlEYUZ0R8Y+etry0bkpg6XKVfIMp3uS4d+WVf5BRZY136oyu1I1rXa
aQWv3FM+nC/Zl2wU0+5yUZma1rbP4hhQDVu/77HPaYGBtY8rvkjFI8icgXLPYDYc
5YpVQilCYpUS3AAUyxS9KY0zGtmgraY31sAJgXlC1VHLK7R/do2//as/u6pXp/x0
R5B5yrmc0msNeVrV5B2UpoVTp6z6iQ+pHn03yvwgYtVP3Z5vx/IZLePHOwXOjBsv
f4wmx8Rmnjvn/BqPTsmYiviX/8EVZC95ocO7P0Z6R1vwaA8EXYtFSq7JlhkLxa9/
v4h7o8iXsWdmt8vo8WbU/s28t+sv8j9GLdLNgIuQcZy2Ub35p/x99uuxWHq35nTd
KWsFWKsgukIjp279Cy+4ITs1H+bb+ORGEjkSWRyZfAu0cYV6mSEh1/b//rUThkpx
uBYCxUL+sMh64x0VdUG3WJ/dCFQUrL1EZRImW9WolX2lpyhN5v/Cl3vOwHbd4cQV
5wGAyE0J/yJsHZUoA/narcPeSaSLfWKUVoSy+uK/brKsL+o7aHNSDedgamGpxIN5
YeyJy8FXLq3O5uOs7OB0saE/luLdVSB3Cc/WvLzQDxu3WukwXxM6ejPJXBYuSlwh
0o5cZiDalTFiIBhY1PdCpoiwvP67/BUd6XN26fr7CXJUIVzq+3GDLoG6UCpWcpP7
mGOZkcs7zSp3yLU2PC+ShqJqGKPOD1aF9mGtLJ0vuRafshdswxi7torN1hNKBlHc
r3Rfvry2iKbLFlkAmvB+/bdbjCIXox4qyLa4nsMMLO/dcL6+ST9nrI700DRgHsbR
dcus27fCRQ3DRp7sO72Cs58r85MDFyEjkVdC17psz15qKuWtl2KysB9YRNjPePJZ
+/QbHsLYeCxx700M8jpyHvqLScpLzHr3jMPSSBZ5kLfYS3LDU3rb/+sUfUnio3Zl
0tlcLUcy9dgUdiOzBhR9nG631t3DKO4Ib17/eir9FzkCI+PpGuCW5c0Q3Ks5k+gT
OcQBwd1+xjP0T4gOPaZVJO0U8zk+ULrX7+WZPNFYoPZL8KZovLAEnUN3kEwIYfZM
JhA3gWF56QWSmQjQjYP2uky2n6vvMQlFT4feLkH9YbOtfOYaXeVmpwCMWZsp/nPi
wcmlfNi+2PFSvk5wF5WIxoGHv0SIqfgIgfyBr5/UDTxu36Edw5SIWTfvs+ykN43c
AWqPSyMVhP1RqCgLjUyqC3O4TwQ3qR39e9nBQGvduvwAbD7P8yrcctfXiUg/WxwC
mc7S5MAGCyGR54Iu5fcwJD+hoO1H0ShbAziQT805VwYkYYMRVfFh8U4ZxCnIQqvg
U1GL0Ywx/pl9jq7+tQp1BHxS8CSxAvVcYYpnGJASKD/qOjcZu0GCl2uhrSPWvyXF
0PBMnWOs4gvjjuFs3gNWoigN0xJy3boARLQloainPgZ3f52engkBc/5vU7TRNLGQ
pq5Dv2ZJKzB749CA/0ipcmekptMd42z9ySWmGL0L0Z7huJsJyPPLHPWGasKaNprK
Rmhx3vMT38xrrgTPmlVkXZU4O+Irq40ZFAZgIVT+iUkC+p7Hn9l4YA7m3ZT5ax6j
zNHzVBpR7WhdExBkJE0Vvt273IwRHe+SrQlc1Qz2TnAo2iylhHUz9A1cbf9lm5aV
wfQQZj0SZgw+7GipV62sxfdCHKyl2C3E4XfCENdfdhgI0jWX/UouVXiUZSl58da4
bmCxuQVVG8hLaDfjS0yCMCzKE8/9dXSfhi3Akdz4T195c9UcdZ1iCGFKp3NFPJC0
FBVcqykTlM9mCDAW405chDx8dD0f33xwe5UNV0aE0E+Pg9blVv19WEpZUX/BCFL5
JIZAZrtZcQsXCNKOCeriiOekbcqheOVvULeoc/J1dAV5p9fiiCSnL/nVQNldLmxW
4wVr7dOSaMhqpyKsW0wq+g12BfrPrk1hPxiIjaHkgZYcYO3BjFT+wb4T851WTF1o
cdwNeh8uQdNmqykTP7eKiZvylVHjYDy1zudS0OAqPPSvp6Y4K2lRRRZjo54Y3mNl
R93qT10Zszc1fk6W/3lKKQK296wdnDnOgfGUBxWhUQNcPNFOOJsp2U6IpGlwRD7C
8P7YJvlwPhSKfEqPY8g8yNnD9PYXq0zbtnjB/r9IdAi65Dqxx7NQwFuC0IMv8jOq
VTSvKODsdL8cbQ1GBzEwCFOhuoSkTA+knmIBNMUc2SuiGG8y/uSNpyDFlLa+XRYC
DTv3xVb5I+Z4pqHlcGwlUUOL+JQpEVOvay5hBkqbFOLtzosNfnSZk8ukk7q02SxO
ZK5eXJcTNNJu6019qOJwzMwJ76kco9KbA6pIwv+esOKo7GY3NL0gGYowZJ5MFJo9
P4AqmiFDIvJxWM4pKo1u0aVXpNEoQ6x64TbKpBp4g5DMom0MvdWVlVmR3/dLMpMy
PnYf9VAighR2Yhd5Fw3+ycG0WpRTAfKKk8hUatprSA458tznO2Y9P664pyaSIHs8
+fdg9Y0t+lfXOBZzW/qX1oiKnhLsTF9+i568s+ax2IMr6JVv8RDaHeX+0XAzS/xZ
/SgSY+HzFIBa048pvLCFBNdlrlO+OO5tbeXZ+RPf/kMOp0cIktVQQwjfpssMrAPG
LrxrZbSV/R9R/VuSAGRUWMIDwQr7p2XK+h2EqoQLtTQkB5mTvLOBl20r5LMcECnc
bgZe8EJS+U+ZXlMfhNzKQ1IKvYoG4n0iKWphyzM8Edz0EYIJWN3DJys+VKi6S+p7
r2uS+x3DBqBboueUp/D04LYgjmxXP7zPsdMwQ2JcyofPpvm1HxCZbxuZUFAZNKnp
oGMk9YmNTcg0lVl0AviuuIGJzCPmpKTBK5ZzWu/vSi1uOxgoTFFjlzZ9s13N9vqt
g3Rhix1q45avkEb5RU9i+eLEkc+6r7pEEqVczwdAYIjGCOPghUCNzt4iVm9rA5Yd
k9xDVFhV/89yByqdCNURHaSfZWnZT/MtSRnN7qofRd9F6uoOcyXjowYFqXBEzXsD
GUJ16bHiKOjdNA4tjxHsAJylsjIRu3opsOfFVVE1xK6U+iF5FJPGbGH/qAq0C0HA
alNedEJlpUUswcrJcuPsuqXu13lBsnbyTDof3DDvqPs1ZzCC4ImUpuvCqDT+sq4q
NHpZplM43HgVtbdLjirvi973IRV77qBIcqzRfmMNoAwVGYVWxkIamEb6bLMzRu8S
5PkzVxGGPMbd2jL/9APSHbGl0LuMqwHY1TkcxKkrBm/ucIcMWDAs0PxiNETnKkn6
Q/3Qa8WOYXrubKlV1rxSBuwV2+Qgvx3jYLn5cy8QOr+oj9pLqKBT6+XzEF2/86V8
uxAofWoqKYhdfFpX/4OZDvU7HlK5IB0D9jaTwrQoPp9HbpTAZa9OXJrJY7U0LyG4
LFfffVpnmmFNFpIfunaUtOpi+ntcabc/KE2A66OvOhcUrJEoWVgH+O8VZD+lkrI5
dElTQRjuzlVT8Js7+hrGhQR+i8+yxPvA7aUC9fG5D1a+dvIJ+pJFmsUAa5bb/TGa
zknjox2v2W9Ss5ndCM9QUYCVE6nRvFtglA8ul5B79OMA/dZrsAzPzMfJhzoukCuR
CXM0Z7Z9mYvxRFhanpiavnY8W8OqI+aDmCLR7VXdR21f/TkjXf+rxBOW5IL53Gvb
ujlmNTBck8Ipv2FPLEpr+D6GONQDyDOtWotE2TvYtUayIojjJGTEHfCb5FCFLJfx
QzyFhFZ2MU+dlwA28UfAe9xBVRVOZJErf7HC32HaWZuKl2FdjaYFA789HGJ28LM8
LD9ixf9UzJs8azTA0fE+IAmozFZSH6wlB/HPobOtlnM7Fw/OFJucdSVGyuwKJti3
8j9+Yt8KmoKMJstEM/SrzowcZA9xjXrdi9078hvk3dthEqa2I45vXTdDLEY27FlC
itGiEMBvwtlZJaveNzOWz98kRdfkK7jc9HNGZyIM01fvk5lHH9c3y4YBHzfxpyFY
ey3Z3gGEYZcf+U9XZvQjGfGPyemN9TKSRr3/pkVEtaGvjftrakYf8C4o7kTmCx8L
+yGjKVboJGRDlILRoUZlYZ5i+7U/Y1wCI86PI2xIyDSXy9VtLGfkDh32f3NSwCgj
9KFKdUp7O4/Xy66yKZaFHccAlNyBb8Y3hEXVfT6CxwRrpX29wvnRbghBPEpn6oLW
b1gHHtomCZGvz0C4fwrfh+H7Cb4Dvjc3eFxNJOX35+Kl8opVJOeifHJSGB59/0qG
KXQZuFBhzK9AOh8BUddZaM/vfK+V8bUXv7uehkARSVQyX6oKnzg6230HF1bNkQt2
nSjxAIif4UlGuGGMwJBzcxK7VstsVtATyw6Y3pZW33kxhs1JGuCvURJ/FuANTwzc
wTcBPTjIP7EKEGaihLxBYuV58WF1xRvIZ/6KVY3aapyJA40RX6pTq5UP7jfVzFAa
4pl4MrnN2X0OGTDie2NajzZxEcYjeGqDXHZVzpbfjcw+xGRpZEPJshJiMueV/dkx
+shHnPgi8qD7AuJXP8satmoH1DwDgctK5UCKzhGVz4HRRYcGtOgCnkeiUPZHpKAi
aGEW4W7Xz++8bkEKExMnU+/oNQyz8KU7quqIf7B/81Kv8XgtsVLsIzJfId8m0wtN
o+8FpGzXhROwXQmX0CVrozsNGoOc1sNleixyXv+OG5ZByRjZUv+ebzDkoNF+JtqI
0eUscOgQHQGpxNo8jzjRBf12x5aPIe6gGLGQ5G/OQa0a+lIzyAlVnOIdsGfgCsLK
BxG70mHUdrReyaKdRWcBhNDJ1DTba4wPNcFd1iPI6RewDIV+xKIqoC+suZSWN8f2
WiBTNd2wmywc1gOo3fciSNRkmTUs1oYnYurf/mTlHuJGTiyyRxps8esI+B82/av5
Uirb4e7aGYyzj1grt69tHkk7Xoh32SyupXneAiUsr1W8l0YnsKKzqQbE/8f4LkTK
2v3Zosw35QVv82TPwLw0KTlrUM6+6Wleyn0UDgY/61r5mXqaymsOT9SfdTf/D7Kd
1Wxa0DSfpl0z7av1SQZloOHJOhD4vn9oznd/v7fVSE0y+KsFsZf0VDfIeCDnglfL
y2BsetDBYBaBvGg16uEfw3o+M3NWgO5+ZFPXt7OBSgslNbQNXzShgp0uWdP4iZJL
gOApdDHsZL0dgtjvJ1ureZ8CQ2yB139Sm3Hmuk1lyH5ipqmnJEsnnj8Lr1GwfSaA
hvqlmLMcisFwxgFZfOSwkcxZdERF0vAX6iVkD2Dhn8HhFRLwXSBqyZcBrygtLkkn
EEbBZvS0UKhLpLqk7joLdxchuiBm+dizcyMmXrj0vEr1XxLg+EaGP3aJ+QsYfcSG
4DEKtK+Gpk5peS1zpIsAbn7ZQ/dqbWg9UMszd3VCkaqDROkLa5c1IImELSOwCveE
72Md+deGP8BkDNkG7IFAkdHvmVmYcXEJrIrXbZ2CLKVGSoEM3ktdbUdwdL0Vpd2P
nuVDts7+i/VnY0eN2Zycd0t40Xo6cW4+RanSR1NcDOBR43d9+MWzRcVyd099MBMS
I1GprxKzF5TaOT8mrxKlD3xItlbXHBH0jkqkj8O7Vt5yDB/L2j6KGKbxh5yBSKUH
zMLKGmB2UeqzePd+DZhEqqSY6gJZKVUznl7ktqmsx+2z6BWmFPtDoPST+wVXgP1B
B0bh04Op7v5s9YjO3i2nwyDPQmZztkv4ip2Tccd833/h/nsHbJWYkr2nWZ4A9+iW
y2S00SKD/Xjw6s9dXZsZUnJVa35cwagAexN0csdBRwLLYR/nqSXvGSV5CXVQVyB3
cpgeCVFE7S79kMwtrXW4suKqiamym5BUeBlop4jMeF8ZlgW9glnPBzzsUMiyuhMC
U7yUHcR5KYKZLOoMca3hVUXauleRWDz8C9dkOFArnk9kbJkGI4Q4I270J1QMcX0Y
JVqHc/wk3o/DgOlAhZbME257yz4NgbSH+pkJ5sFIjr+BpE4VKnR1OBpdM9ICFf8K
df53Nqh1iPxHAH5v2JG5secsKQbX28U2yb4BXBxjc8ZXBaCOqmfRiofXZ5Y265n9
vPmocfXbL/pnyaS3yjuVRA==
>>>>>>> main
`protect end_protected