`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
gMcHP74wBZczB0bB0IzoP2xg5wC5NPjD/GsvSQ6VQgzYAsanETMwwsWi4yhFtJwv
5kY07u0WerSDf8woJ0stqW5xF501W3JLIS8KMiCOd55RHBOnavjYiaaLeu7oUCmB
TtTS1R4sO325rP2zOn9YwRbyyS5Ljn+PzFZZUmkt5xMca3p5NGqKtZW2dV6Babni
5HlLuF20Au601B75m2nv+ZRoGSrpkNElxoTibONmX8gBflpIVE7BehhHwaKSucEF
pp4QQ5zZAZjEC6aplZepouGVggAulz5AahlX5bf4opOVlB1J7IrgyjENtw6ysQ/q
DzybQ+ipztSXBGhmcCVU3A==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="jAI3OJE9Sh00Sic4PtM/KZ4WjwT98XM8AMZrZsQkxWQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hyw9IrFLPQsjvXplweG8O0lkaSLBN9Ijv4B5VdTRt6ipKJT9Kzsb5LxCKvkQyF9n
sGPOd5i74hRHnkHfYISGkfxGJCa55ieOyFShOsqTKRLxclm4oja9vTIey6yFm1BZ
54IDCG9h3PqfDiTD847UCSMRvFssyycwv+BRHQMQlFs=
`protect rights_digest_method = "sha256"
`protect end_toolblock="BnLuc3jxknmZOyxfJK70E5kp9u9O8IQ8cgkXv26kHA8="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
xABArkLxBOK6xG+7CdOOiGu0zbCbHMrEntFfAZEE/xRFxZaAZl1QLkuFI77OC2KL
XxG/mrHJzO3taVHgwRXNLDdc8ePbxbAiQfzV3NJLBO+gsBjmIymaCa480cPNpHLx
MvpLmpyOzKTdfClpwlkWJ8+IJ6BQSkacbcHTXlH4teS/Q2LveSMlvuYXreo+IDPd
9ajHzomHEg7WhvAhpoV5DeUNMvVIsEyX97iSN+sSuAkCfeUoHaXm/OAZ1qqvq3P1
PHNulZoIYoiTSY4qmRIWWiNiGSkPAeBdmPMMlpfb4QG+QbuqZgqE/Riv5SisxYGl
ThjTpC8f5czwQVKE5lKnwDFUjOJyOlTHu0L1LGkiX9w+2jPIywtSibWql4qJ39KR
A6smF6L0ttvxyAMUfhr2MkNIHsz1OQArcSeq2Lvv02s3/RqpFKLxCNIf6HdqUfdE
eKbbWOIojnHKXlNHhL2P3V3OKfLvu6I5HLDc1mEZlFZ8NAA7mpjYzueb6xGV5TLi
7QiV3kEIs7KP7z29R85cev/y4N2dMIMnqyxKlFhB36ktIgmyF/zWfMEN7L4e5WQ0
hmek1vRzTLNABag5xBd6r9reVLU1qgo5csmLrKF+BWer7CDSnT6cLnpxE1zRmaey
GdE0YGojUk2tG50eQn44bO9GdKWgVSPJnYstbUpRe8z4w2hNY+6IMMQbQ1l+ChS2
+M/JGonR3w2It8THLuxr8I/2bWCu/d51xOilpkrZWXH/deFT852JNWJli0I4F39p
8aYzBM4jOiC3UVPER6ahQuqKDdN28w4wvB/3l+2/MghCNUsF+fI7iADTuduboE4/
wkCdkzXa+GkMSVqxslf/TJWH36JCYmHNaTvPBlasAcxoo+qZl4sIS8g5ASSI+opj
kzsI4JuO4x79LFtPsXmyuIJOWRbGFAywMmM+Uf5LYcVziPXIi5okdAB6S6AN30P8
3vqshibsIhbAn2N/R9vjSCcZdIbRtXHKaIL5SNDDWYo+WxF9Txu8GPS7DMd7W72T
ZJ8VMSw1XeEz3cRJld8xLbLG9dCRW0qPMW80A2oSYUuu2CPNbeKSFzFqXLNJSMs/
mbT8LcWUzxKMN8kPSmpHbKVFkSWCdcBZWsfCNRKDKUltAVaMQZnAUs7OAHz/dXGS
zqyitf7O1MNPRqtMKml8UFxJ39KO/xh96wXMYXZMk6hohZoqObPx779mEkEBrhcL
9LF6ryH9KU1Jh54v/jLXNAmYUv0sBqNhnUeCYAI+XGHWhBdwQ/XRVEnelmz7yLIT
HH3cTY3ex9qG/cUPd8Y3u8vOePrGNjHjBQ5iR+fHsfFzzMCZw2l3vwY9pXQwPByE
AE0oKi1JlTN+Ugtn3+DaxGhmkWEoxmGuV9R6+Wz7T+KLT/bpIVQh93dVKPvFAmrE
8TWq/CsSjevgYaQB7nzwy+X5uYlzQO+AuM3UJg6Xac8xhlTlUsM1+1yw3RDbJboJ
Zs/XPcyMf9ByE26RbbjS8r/QCavE6Gf14eHF8iw6Eo7OTG5MvyZECwqY4ZLBXMvl
vOlBomIGz6B16/f1aiIEWbfxc+tjbTRyd8M8ZaPLvbBAbMCaoBWEBbh08bD/b5QG
dauruOBwel1r9yZPC/jN+hWArsA6vVx0D5Ux5FhLsw5RgPU3QjKgIWPzRUYjRJuM
ZS3XMlCGJFSD/Ftg4h03vIYBYOunpuBPvek4Cub2PbAGvGbY8+PX+z3X9YEjlwhf
DGrQBL3T83606vjkweuT5jwH3WNLNIVG3/svbfinmC/YFeJGzfGxtNZjqcOxzIXp
+1bVAH7TP+FZgA+YuaFdijXAYp8o3iKR+Q52W2XSrg4lPZB1yJbT+ixcY+3HZp9N
2qxhEjQqy8pCYxDRCRfJP0FBO4v3eqHAlJ2DqCq2gLSdx2q1lVPpvm+esRMa9OJy
+90eqznKKHGfsv3G6u+WDOumwZsGjmUcsAFk11figuCK0/hI/70YsHdjmi+Taqk4
viWJHEeH3/hKmgB2bZQtBqfs10xiDedteUCeohxokmUpYl13UJsg6rCBIq7wUDk/
+IkhM845il0d9EgpupufaYCIFzesn10yPUCbjIgYMaM8SXfXcNsxJEtEY08d0Pso
0fuQ3rDVR7HnUbBTv2PVYjKPJzgrknN66yphVI9M2B9mmqywyIcCjG/s3ICacR7H
GhSP628686SdorvTd+yQgo0Sz7CalZaNJ4sbrIihqbw9ZCa9mrR1NYMoDvsEo9Bq
4mjjXC42uoN9CQNjpItJkHvxwGlktTC56z2SYWaili0=
`protect end_protected