`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
wSlRvGACZeltNrdyZhP4eWHc3u0NosY88S/neykwPHS0N9EUB07m1oUnFcnfuB81
iWsnbcqZui9Un37u7DZwvFyUcUSZtA+OcGP/jvb1mZ7f8guGjLglIb/fl18zePO4
Im2qjsGiYHlSnhxG0phkGIao2bALf+9R/s1OZI9N60Nn/cqjmUqRDGaKDNiUSVx/
7oAsiNCyrvsoDAAR34p4ZPfV60Xv96wCO6JSLu2JxnJ1oxP6UMnbeyYuv53B1n9R
uQF+Nv3K4UkruAjl2TViIIwq0Zonq62+shyExKCaAaqzzNEDJxIPzXDbRMO21BJv
rlGh6mcMlgHcismgcj0pYX9y0KwDR3VWTP4O5IoCJ4vbJ7e+Zlf9Q2+qaWKwv043
DK4IOmUK5BJ95LqJoi7O89kn/dUKtheTuwv5OUyIC3c+7/1mk1a7e6NZgWSa0qIp
2A1aD3bUNza2Kpoe75Q9gJgR3H4du/lcM8RzJhZeSqaj4zJDmy+0rVcspNMovRC7
0pkUPJFPKRMqMnfLS7iE6qeIGHJvsqCXTi3pIsYVj9q5ALF4WnswCHQdV1iaXdx1
lg9Vg9G60tsyEGAhfWNAqMwQ89pkS5sA2HB0BMGJEIqkt1zCCPNnkhkOrCRB0eM4
1Ocho3Sj94WVVk0PtcBEp8y35NPQsaEd8iv6rZ0WjMFnrPqtlf+QHZaigAkR4kZf
S2VvtgoQTb81C7P6Kky02NVh9GEwHyknD9eTfN6tlX+5YY7sPFUw11NPF1reYIxV
VPYCerZIV1iKYg7IK5oZcIBOqwdVEDIfMTCeijywq8Bx3kJi88FLbElWoy+NESoT
RZ9Hz5E9Niy038HGxV7YHNuPJulGf2wd1nqXGtv4CnMvooEcMN1THhU9YWO8FVn2
OmpzonQorW1Rz87SWJwjw51DZQ79Dnc90XN8nx4yPhfNrXcUbS1IjxTt6ASSXlas
UOf2qOKGPKlXD/ZHwSSipBrVQoRhyA4xivFyfZA+u7jbG9Lq6qY77DK6PBYystG2
6ig7vVuln8xELqjZtP6aFsR8d8CMGaD4pJjWTGSjCe0n3SNWMCI9qA5wwKvbWeAv
iIcmLrYxGTx0Wpc7FeaJzunYGlGNQJQ0EQ5G2i/3QUTJfJsN2LBzAt6VRZjKhCtD
3MIOZRD97KaIvtm7c4c22Jd5+cnC1NANXQwNQrDZb5TqY9rf/Yat46zKiH9qEZmU
8/gqmxeP4h4tloastC3ffMcLmvsWtl7uAHBfFiybvuVwMMd8oB61bk32t/3k3kxr
PCPSa98jCQkFh4dBS+QZ3MyLR+cGl68gOm/ygqYd7jHw/fG4cGDwDi4/ZXOorj/w
+CCEnnFvPO0VDhnjAUXqDxfAJXKDLZdA0uq1/hWL6Vwjavs96d1XPQCUjRV94REh
b8oJ8HRYAXE9W9OEQTz4PSYtrPqY1gtnYm6Vu5VhzvmNqT3QRENBpwr/uC1RyX2z
ufwkZc1KSKA3J3agtIlTimaPLe/myEEoYiamfMu0nckv/bXdjMdmUoAcrW6N3JE7
VZhL1XZVDrKjqH6bDiv0FNKDSfuXdNY6fI6YEWzKm4loJC5wX4WVXeC5KRqpxxnw
v3AnC2dPkeOoidoxqFYc4YIU8M1fANuL1zkv5lS9TlJbsK6ed+SLqXfNzrLvHy5Q
SjNSvruMnKVlGZ4eSFCXBvrDyoMjXBLyb2iPMsOZqvPM2nJbG8edSo+BZu7AqoU5
a9It91FhDw/6cyN2Go5f1udFXMM2oaddGVoTeULtefz7oLuTtd1tHfK4+92BfDRg
KT0sQ9Xk5UNFAHLrME/+w97nl0eehnf87rYHsNiGFNcyunGYqKHgCG56E3vhe4rl
nFqau5qyLJLnzmp2hgFLjwlXSve9hc8N+0SqcOG5yn5H9uO9riL+b9kcdItsi3sX
pckvoe7uKX4LtHzPQGPt9ThpH8ptp97wyNpeVJfMhqEpkGOkVNJtC+tltRfICj/2
4UbNSjITlcZYJJCJiNfPyAO6RvGLBSpD21kbuIUzwvJAlPbR8PGExBt6DPwcpf2G
+zo2tzLo+qVmbtjEyYAnWM8fnmxB37x6NFCSIjPyVRemplA5k823IxOgV0wOZdxJ
4Qiw4iRkktEs5vT8ezeGL56hf+dNuYjCHjFFr2SIXqweMxLjPLSYmWEUT2UB9yTh
wPQO6GROHcp+Q/e5ADaBILtXgXPKCBwKB3aUG+5cJLnKcRB9SHrQagA+X7SV+rug
LiB13KUT1G66WEL3qf/jG6mOLzPja44VUImvuENiV/tAPVodbFsV/PCLClonDyu9
YGBhypf0ermKl6mkCo1bNSr3gGAO5/WnN2LMHCswa8mn8slTpJCj2G1q9HZW2qC7
VR63VqGMRu2K4cDFYMJk+zRurgV8sFNdnnt+J/um/9MzFuXvIWu8LyvghqVtoqeW
NEh6Fmf2tMbN5vAyl6TN5btGSbvU78e8eWQwrcg5hBuqod6LFg5cRer3gIUHjFhG
bLfkBwmYO+8snV9V041LPiXO5P2rIu5SE6QggeK9nSOronNB701isy5UPE9daOb5
82A8EutnUVCfolFO8X2WasCxOxXyy/C5BlXqna3TPm1jda4FnOxGB94DyI1l7cZ1
BEFrhOTi7svd4uBxKtMIgaBAjfj2aAHIH2yyhS+Cbbf1+uCwDV4Bd9X5oC7LTUPt
QWlOUZpumXzjQxEUZknTGQSnGIKUId9OpjN0E9T3gkfSAYTd+QLIJHgSVIx0c+MX
HV59OmLtJpRsTrCxCupHWBRHuJynEud827bRtiTvBAaJmkkHso0QhoMXc5lXodqP
yL/FdXSDzBXW9xtgCrpSbI4bMUxti0FNUHg1IOfltObVToc9KwrPgSUzrsnGgaxe
1Ky82olzU7nmqf270mId2j7wn9rVjXzO6VLyfRBCXpMV1grLv+0+BjhsCf/lfvvW
/zSWdm97UUmye9zK41pYc3BSyV71R+V3AfcG488HNTrrpjpYp0SzpNl3c+DsZsJH
ghAdlCWmUC5gEKHFK8eltSlDtfhdI0oeBQfhxJos6B5zphomjDOHqY+8a40CZLM6
6JLw14+gPstiHQPbQX/gLTUaASgKnW19rvOHllxzz99JupiUUPtZd7GpRKK46Z8x
2mikUs9Ft8byeADb8dOyJjcaBjFufsaIqLr842qDK7NI5Fk38rsT86TcfdyZWAws
irFj0fvFsabdXl4zB3ZGKv/ixPkYSlDkge550GOmy8deY6WhUnrimulRyPP0Wiil
9+CjhXr62RrASyZGMaNaxqaD4nlpZogHiJFVxuZbhxnDY4jB8aLreb65ypDVc3Fe
NDfJ1O65mFQ+/eoT03KEAXMtoAJFlZAHqY2k1Ag3V2+Joie9MDNJ8XoqdYhH9qSg
gSOKJzNdBv1h5w6BAMPWT9ehyzSrGsRL305UFkk7IoIhwd5sV1y4slhoMrsBkIxO
8X0jHRzK1OFJWcSp+i4znM2FZf3dkldcCUJouYXbkVy26u01G3bxRqjanCP86C9D
zUOKM0Urdpy7t+/rf6l8FIaxSvHnQxs3Znlg0/qTveFYnNNClOu+aqU+nI9MX4Kk
fHv1EU32SLQb1K2zrXWGiCaV1osdVwLkgtJ3QqGgtx9TJ4Qxvy1bCJIhjvgZUNAy
kZXy+0G1oTCIzc/UtXa55CYf4LV7Um09KQOKqK4bBUSv9QwHlh+vOmNeRvx0ibW+
VJEt3pED32nC85Y9nRtG/A6bL0OkOPGDomXXOBM0KXeUzQtP2WYHENtv0C1MFKhR
zoi4Xgq1JcDVBu4Aj46A5kqsei1yDeofoHNPr/aoJTYMKiiUODLTTGDmT2wrQ16i
o9j5tDY/CqDs6fGbQJVNB91bniJ7+jb5yyn9sTaZZdGOiDQXvcGLl0quCYCmk4GQ
KWFxxxmSs7xoqJJSQMJsepJR3BHvU5wTEYZC3yHC9wuz3S8f1kKUPGXnPRUCbzPA
qvqWSQDt3zIBvSwEphMRs5HcKhqY3Bg1n+gAnIgIRImifJmZyb+BU4AW9KU4K6Hx
bVlGTmEz4cBQ/lhtEwsUnAgzG2WdwTCBl9y5mYS/PzOssnfg9VzxRDbNFmXRbaLi
/QONYkINmOqa9nUs5raNrO93FkETIiMjTYg7/Sviawspud3eSNWp9KqgY+1rgtYS
ciO5cb3ehppFHQHXHT7jKPJOBe24Qyp+GfOzj4ryqDDAXcb0lfRKPYK69kGOQtfC
sCH9b44HlO/txF7S8C1S+skwlM75l4R13O7iBDvT7v5RL+KATcjgDHe1RdzNl/jd
HvMKlEezScu/yxvrOwAKiMzuofRpQwNMfPyZ82oLqhSz1icOKjwm5sJYpfErgJ66
Elc++Wg14T8WySwoJmxE4TPIXloMJgtnnVYV0pELdQL4GU/Jrj5m9ioh2B3Raukh
S8SIfG4EUaqrn81K1G7/vEZO1yOOvrQqxNkDZlqk+we+jdComO1V1f5MPo7x0FI7
aHyVX5i+FxsEUTc/L8um6MKha9lnCb4WW6tzYYepzBtg1P4xHi640OK7MYwZ8vc0
i2972NGG8YzojBULv6AgHLmmQRN7neyYF6PNl5W9CpJcCvoYFyA774/auTtm1oKR
uX4Keoa3OqpkDtcp2BEpcwgWquwvB+cdM3JacozMglv+keu+roI8VRQIhKs6Ijjt
LtJaP1+NSMrGqI+qfT6//+fTlY5nwLPPwT9lc+7pcpFibk8xDhNSPIGGiTm/fuMZ
grSA1Pa4/OUJvvj1yI6YWF2kfhtqszZpbas2GG9+4jZ4nH3IHkOrN3IVH+63ZCcu
8TQwDqxoml4prS4zIV5mfU1gz4hHUBVS8V0qcFF/GLCKo5N4HqQlPfJnv+obIi7O
az1L0xobb29HsWGq6N/F/ekJ/1Ih4w0l4H0rAJ/cKIWvZFosfrsO77B6syXSs7JU
OOr/VghXMr51yxGm2j9OGOPcd4Gns1VgNncO2yNBdMJ0WwoAwUeXfT0nivXO000y
Q2zOFa0MpYgaDt2OSOL8nfYBuKF79aKJ6NF/iynwNPReSKMio3yT+SGazYlZ4Fim
62/rX5De3xmVhzmon776kIqyg18IfFlUCFs3VnSWalkbXblDTdxxF4VM/xZRFX9I
i2fzMQZ31qgPHbcJ6VOWpHrKVBF2Ht/qjc+BpNU7xZMGA5WYnylkiPzxX8nhsQsM
UBBgbQPOBaSbrwjQ63YYEg8wrj3ObP20ov7tXloiV7NDbgixXBZCPHU36Aa561pN
80k0EvkEFcr/HMB2+OG9JqQnuXe9rqi1mVFzmaU+6DBhJHcHU3vEZaN7RsgC/m96
htlYunTd/Vv8OZePVvbOrHdW3cumox2b6NR9/78pgRvKfxi0+ByBJbq6GqrCDXmi
g6HuOYl3d0YwhC3y2xoBxNh/AvReQeyv2MZvJfbGoS77EVjgDjFG6/I1q2txnT3y
DFAKS59iQsxIBAVvK+CiZCY17+3ATzKZLZqQCSh3UQaCrBs2E/5z8wiAX+fkVMj9
NaqxB14xosWccMOzFCx1FZlNCbcm9UfdE4sT7HIYxbWOzdRjNHEg903SBliyhsWe
GEDpdX0WCETwZMrNADuVC+R6BkqwLigksiyCueVuRpuOF9hLZ1zXFRhRupc1/iSy
NmyvVc7BRgbCG9kfWr1+QSRQGcZICJO/+PU1x1k5J3QsIRgc22VtAhEVNVdESy0T
H7zv8fu88PTeWh3qG0iWbG+869+f8ja2ycQC4B8ce9epJ3s4PFRa/vya9G6jjwG2
AQTyzdxndFDzoKG6OwYXoKs8YREl6KAkrKjWSIdnxEmW7qJN3e89eQBUhaofcbJC
cbAAu9Cl2GqEufWjmUTUm7XGeE9y69qizPbrBeC8HRFqSxFTBtxA1T/Qe8zV/klo
ol4OtC5di1may1RJKhxA+nFoN8e6gf7razxdMbHZrG++HyQqSYe/lubtpHo2tVvd
z0c0VAPyco9Oxe7LSCy6Qm6wTnAaw2bh7oJAN+yNOSv/75Um5cZZvg4rk8q1ciQk
LzXJPRo1KVhcvj+Tg8gDp50X5aD+mQoSnFbnlrBgS9VOOmQG0+knUPmj5VZ2j/Wm
94F1yZ3EL2g/axM2CZTAF226GxDqtObGw96cAno8vcuEDDsT8PzRTpQxf9+NkmF6
99E+Lv0u3Xu88pkgo6cZrtWfB8iMKf7s2O6pHr0xiLwBK7CSiXybtapB6kOfGap9
8kY96dQ+b4mN1nY+wJ13uRj/GFEbyu/8IrF3+xn+pALKryR5mVNogvTnhrdqRdF1
qfILUGmGtOK73iQ4YE1h9pWEA5hYeLIU9EdP2Yv7gLT/X44U6OTkP7qnAKI18OzC
SGkkL4P/PAPtM4Dk26N8lRRtAF157913oOCPeDQiyfrIWEB2066su82AhOmP6ju+
/Adndt7pHKAtA6R/BihQOkErHEr/Ob2Yv7LBqNN4xuIBoDChrp15EO3REvXM5Onf
vilDQff/wSZncDMJXvqZGlL/17rzC2zIMxxZ6f6/58k6yvJfCoeKrf0oiL5nq2O2
R9t4l4hw0OCMm93sX60YbYga/YgTWbdtzYOWFGHq8i5s2rszo78quT790ZSVNSwS
k+zCYrTuWUQmUeoeyrMjJMPgitBpmgWGGvFGF0xu1h1PBPu12oFYV47UZASmUzdN
SrVJe3tW/7J3cbJ9iTZgNtYFfguhZ2DUt5AoPSlbJiMOEufcaUotUVyDcmrWA4B8
qotvSfFyBbLWICdAGN7ZJAIRWF1muCDDTnrrcKXhvU8sK2x5/A8yo1tlIttlU3mK
jhWi8aQwVWw9mYDwQR7iURVAi1500VOgfQSw4UmOiy6GXO2soUQMQxx1+mJHC6kr
+vMQJK9Yy/Xo9CQm3EWO8wDqc9DzJX237sOKPQiBiq4An0eZ2I1p9zM6D3fyu7hL
zwyeBccBJMkgOA97LgGMveI1xXJZ1wIrQlulHuuhfcP0n/+1OE3CRPAAt5IIAtF2
pj4RddqiCrOxplkX7GAbFgW7SWuo6lyoWJtFxHHWy8SWx+NA0swGXgeCyRFIXW55
BMWyJi/5ypAaPPVci8MJygoUcNqOC5h9IXX9yHW+ZPv8IIlystUTiq3MX2sjkctZ
oTvc3ro8bHocqJ5twdyBvBrxGIX0wlYeMa6pbehFUuhxJDHAMSSIrYl7NiggNxDV
mTL6vHhyLaUCXUcxS+zYaaES5f1Gq27n8ybdsnDLJISOm/sDAet+YRetaVMcWUTq
zSwywwCcQ9HOO0CDXJQ9a9OLPbIknA40z9+VMMpQPEk3rCDqXN1xQwORmaYz2u6T
WV5XlqYZOjF2f7+KPjBlzdPMHP/Wb1t+eUn3L5yYHjMFVyx34ZIrsEJsE34dsZpy
28+EgQHA66eGwW37FJDX7YiPns+uwNCXWkmZdBx+nbpDjIWuZlwEsAubf/og+w0k
1QCcatVWI6xdYNHcVDP+2MSkFLe2EXmg5XWEMlYHr65XFNHWzoXu5Cm8I86+RTvh
rj7Gfh1EXI1LtSczGvYfcJmoBeBDmUO6FP2BQxoRsWNaVDOuLRQ7u80v0ZCk+fPR
JoJsef9aYZ/Bz49bPEl7zHL/jbLTM7cwexcjXLnIwhN7L4JjqOJKXWUxH+bzzALl
nrYrW8ibCzJjhNzLZA5XKWgVqYwjnoz1MauGlPNL77K8kPHuWF7RI6Sz7uVMIUkG
n8hsdKlT7Dn6ltqjjG0Xb6PdwdsYKvzCYILL0TexfzPPWD4Uw7T96JtiGSPqoIIA
avCxQbS2BsJ95Bm7T5AZKLu6ijinrXL5BS9wHpaPRYEzjUmIZF27+q0bd+YBAU3q
UfM+k0TTwGWwe9fbQXBxZ1OZMTy9LDaBgpXgKAlb26AqrkjCOCsQEQhbMq4+/KgC
zNwu2XlRN0QZNIHxGlMl/9p1ydqNwa52zxzduc/52v84cRt8Z2vGOFE4H2NEi8Va
6rUzTSptvJjHf5bbfQVRBoT5Xapa1EIEkPyQGyoLJmjJ1ryEUWHfXrqaAC8oAFPs
LDOocMnWq7YvPf6yCSCgbo28RfvhRCjkAGSohGGZm91CMk8Oa/zDUrI66Mtt6RYn
MRbvlHA7UACFcFqxy0Yo3tBEtFkR4TMoB95UAkP1YEedCW05wbttuIUeGb8ttZ3K
xm3L5ZunJf6xR488wcfLD1XqBJz01SrkAYbmif80fZww0VSS2FKSp8QlbXyQ9OYf
o8M6At0TIyAwUy5hVyiyGOkEXRhn9aX8/dqBvxmVqPsk7MV9Apm+WAgCqCVKpoOa
grHctUAX4K6TQAlcYPe+xhGK0gGmEetWjV8lIIrG/PZwBiJct9Yn7LlMbNuGkRVw
//tQn0kUjqy+bNISkwgrCGj6RtUufIZvJ7OGlhn0/ijy109lS9gZbISLB/PMb/uE
ombz3HusbZ6YM3QaWKNcQ0mpGwMBJMPj+HtT6S2MPZC7REXveyTUYVSKYwdyKzIb
lUuauo3PmT+Z3FJdTkyU7j60WSwZnNJgim4KNOI6S5b0Jl9Um+oL4fmyim5NVLCP
D8Xtgnj7YNgwWjLYbPJfzBKB7QfWkrAQpapAO1xWP/zvFYbJ0QvYAZCl4I8tzp9v
G/sVGdXI0G2vKoTmDBCuFXddKoKIyzbDWPVeHSdUPoxoDD00Kguo9y+1qPqP8+va
T2yOhWCle5Q5vLh+1TIWyPw9CbyXL88+8giNAuTkCXQuOJEqBgXDC2wq3Hp5AsdQ
OKCz8TuXg/QAvxzruXkoEdN9jhBuxyy9xiAecd1Iw10mC8BWz7Oq4XR74GxxPzLV
MHxCwXgHa97mqarwYrHUntR1f+w2IjqcJgrZJTxfZTWzpKAcdxmOs6yMi0zAzLLv
DE+pAPHYdIiDKqbOSEe8bpWfrocUvfJYEh8KCwJSrQ/Z/W4fqQxmMmqGPKFLr3Ga
s9otayZEH8cyczhG3x7lJJz7NxclpktOjQptrYaA9gcyGNkPBRIjmRbfK43S16vU
vuwIa7OnUo9Yrv4xEH9lq4UaUbcA7SctyPy8YPHaDI5Hd3anovQxkfTkPRUPlVHH
lC+zMpZWueX7TECtt+nETgtclRXtOxwYeIl8NIbs+r+CPD7Aqrjr00iOYBRL6CZV
JeXcMs5mM5W52+PstGism6mYZGuh90RSAuLKFt0Np3oWWczAiieXsqWfXBYkb0ZV
Q+gM/qginwaBOEMMIOtxg5ZPqogxJjhSDvHlyirneUQHEULH91Zlh+OoLYXmipoi
U/vVEoiF4WcOmCgTIrmi8DS1MQM0UqCChJwQ2Hwdx907PxO5cY5XU36cF95y8BzN
JtIo2RoWavvONw67w0Eu4mGnQnzYueevLb+E+F1bIrogPHKoe6SeBKI/+w5J3BN2
BEDt2bRW5MvrVi6tgoOytXDOn/nuzjif5TtQb8RfJyYBX0gpvGHpdoQXn/r8nob/
aYR/z9GZ83I5IG4mI4Mj0Fs0ORpwl9SiXzzPG8G5OAj3FFt2TVm3zzjamgKdOter
a1VAG6Ch0d1pNpwRDHZrb8zV7/uN9dRf2/UPp77ZJjgstxjCvmjfjXAXzs/njCHi
sCyQo2dMIR4Y0zYen974+BPgO7k2QGWKa5cqoFFtrSVvwV7QBQ2wCtTCy1/w1BeA
HcKKV7gsAAdwu0COJyT8A4QqMFrk7gaDsRXtRv4EwGaqTZTdF7kSrE+CpGADJjZF
aKkdXyvWr16DBBBxGUTZd8oYO420osI2VYz4Um8m/eEZ19j0nqbmHRELoAoE9jKj
J16WQ6TiWDGD3fi0//9RmcQVjmygigDA5XdSM4OhkYx9RygQn8iBIwK0XNenr7Q4
YyJxwaEPu9ArWltSfo8OcFD7NVrqmjzFZgQ+1X/jWKuzp3aZIDygNcX5dcqkMJSM
uDUfgCJSGBKLZ2XbaRnxVW1Pja67sQlmvjRd3Oyqv9rfvBrUFuc/eoH2f3iqoIwH
NHSdibxJSXwr/HcJhhqfh1L5s/AH0i+aH0s5HBa2sieU1LlZTneHOIUiUVi1HRJE
W+VC/skTkPztm+LJWVh+6n9fSsozsZWUoeMbHkLDd8KXdS1qLQuPvsQwFoCOpPsk
zKpomziuTWW06Wf6rZH7MmZGJjUn8mkuvjvlu6HGUki5Zi45kwoOnwA2e83hNWEZ
e5FAJO8Kebz7NZH17FEb5ZBYGZJx731I7uguE8sNq/cWzepCY8E1qYwaKifUBnRj
04zTa3AysnAvfWg9QeN3SYxfZICczrS9HPDexW4llTivwK2TxfS0tCKcFe49daxC
K0MIsFbQwf/sahhSjDRzDKf5AXHuVWygR7AaadaWEFeFJtvNTAqH4Q45i0n76RXK
v6BY1JxiAfx1WYym1vRYSlqcFlbyuEaBcdxzVihgtr2OUndKE6mWotopS7/ajKcR
5YspeD/EVp5aLUq792ETCEp8cc1w7a2ljXM4z+20oM1F/DxVZ83jyWxo5tTSOrql
ovG991GdhnJxJBFmKA6DdN2E2UswpAjuF5IFMSgzJ32H9+KWKGIHG/MjU5tWqDJW
WEBn/K2LSvPuR7cnIdygFk4b9i3jemkogl2oNdd0wQ7Au+rY/wnvK/o8EsPvjl1G
3e02fMkqETE3ES3M/Yho2/4r/2aNfNhfRLQ/iVd7nFsKnRlnyKxW4WNaQ/KVMJRc
VcQqbhZNic6tNQbLQO+n7viQ3wpV5KoMvO12kyBe4tRV2xoYWjAqxKZQKCQwTdBB
CYB8/CfMbL/pmaM5qH+r59fFJFNBfJjHWVswn2HIydhiEkXhTDa7R6qnYxB2aW3F
9iKZ+aX+shzkt3IeZjmariZjsLbtNdtMOn26hZxSxdjbaD98x4oQJk0orXlv2G37
wh4DS1zscz5CqJ+/QdbhOoipynSCNXWFERIivAsYVi3zG7WWUm198OBb+4Chl+P/
/oT4JaOZy57lw9ixcSIAa0azVkZcet8xUYkSWB3HGSRZ2hSDSPMYnJt9uVdIAhUa
KwCotgY+9orrxmtStZs3iLsy4iGw6ERZXoIqWLwBc+AqdVCGlNhOL26i1Qs6osS+
c7ysyRd2yY8O+q/501DRDeGR20RKL6njMZqkKoATNQNGWAhpGD/0YIXOedVqrE0H
Lt0rHaqilQ+ZGR4LT/cFQw6PrXqKfczB0F3qxkWocuuO3s8PUSCJfU0pbizIsx9p
5dx2pCfBo8+zDyWbV2Bszth5d0j7wt7fVlPZiTpiFoRPZKebLNMK41bTIeqE0ZEI
qenmD+K1uG6xfQlOWXmZj/dDAsVwV/cpNT8wDw9L9nXfahUC+0FbKNPKIgCwNaRQ
yg0XwQvfuzYf3U4tpt2Vb53iCHmux13ai5Nt9zSuVk6M+GEsrBuoDb77830cfVYK
KAsWCPYC04DSbkTTGqwhd3fXytFvsjWKbLV9ZpDWvLpnhweJ1a4jAzzQlU8jmsuj
HLbgk5XZVddd5Ca48gzKViwX36LEaGGqEgh79aM3ZyG4/YMcso/YFi4WKL7+EaWN
dS409D9oHWc56gUkXuC13IqWv6WPrk504TRIt+gWnwcorynt/9Uyv5DhPUwNfbrP
v5vdnE5ZmzUuHxsFLYJk6JMZ3vGEIpv13Fs5/bqZDhYbcsiBby/fuUDEKvnAzzkf
XxcGGaqnD9/TXGv0kkgM87RE2qL2RkizV4PyedlsFCN++WyvTqbESUK+vF+SvesP
gwYwx+RatPiOSxxnr98sH6xq52IENsUVp/tozILUm69708d9rsRWBQpMS6mJU1Qn
+xrkBP6vzi4wTymcG8r5c6gb7uax8d7QQnsCiT+mtui1V6l6dRcQVbiBRJRGvxrQ
8IzUYAJx5v2KnLCRfIQxz86zzTM41VlJ/nfYKUKV9gdHKUMR8sToZoyAEwFwNTxo
67hKdkmLzxqbJFTg6Wj7nVykgc1cqy8H7cHigS85iRxD59AsCvaBawfIxSgWIzdk
/xwjesJAfSvtbUy+EOtODycTGfvNa/arQYM3qxh8U8eiFHuHFiBQJtvBFmcSeNWj
eTGFdVff6/+rDvgZnV3cNEvD+baHtCOGzZ0c3JxZiumNq1qKrrzvAFycRcoQ4Ffm
SHo9JGsbU9wTWFh+clmEHwcMSaQxZMQevCRbRTQYf/f2zHK+tcAUQYRATsyk+h3L
DdfWf7DPL/ZsK41M2N/l7pMDJAEG+ddChAJBVGh3aQO3N71kvtKVwT9e7qbkm7gb
gUNkyyqKociqKf45w4yBiJJWcFR3WaKYIBKCzBhschI4UUTAVf1LJXH3sP0Jx7xF
bysoPYdXiIkW766UIMElXHp5Y+Fl7YmbBDC4RXuESbZA9PEIAEpCDBNvNzRwCR37
TtNsmm1yT53rIeSgrORxHQMRHllADtOV7p4KWi3Vn0JILR4CkRgbfJqCCs4tqI+Z
6we/NNd6kT1pnbkzbFV9TWLFQfVyzrFn7Ol+146fPFbKaZzMIsKmTk/fwdvTJs2n
2UYnKQMPpBWNYB/5usyy+L1zvYgG7xKTZs4WvNiE8gnIj/qJA0p2sqyQr7jDTLFm
IMm7a/llG0x+t1E3xhJxj8F+QJ5/il7S/KcT4rfsCbtPKYpv/EsoEZ9H+BW54IFu
tg7kD66MwFUsLQ7bPlxE1LSxTIa7FsBcLk30fiAHoYVtq/LGroxaeDl5H4lAKSt2
xrhR397oBxa7XmItSKzyBeVnr9av8MBOrckDeXqrck1i1OPnGIXdmwZcQBy3UkxR
OPiW0obflfAUlVWBoF1FZv2zHSYpFg3QT/3wadsJUBw6hMy+7t0kIAS80zfXsHLL
/7wSJfVgbPFbLXLtIB7jHAEfl7J7gkl7IReScemcc4jn9pYrTHcCX0FLgRmJy7Tj
Jh6wGf/xyCQg7abK5BFuQZWZxjWUVaEZpkPVjwwKqs+4Flwb0tKKc0FripEo5XW2
3wQshyNisisD3T4muGEJqLaMkQWzCKM8RfEaqfoawLTFd5ziU9fjOzuEnajGFUxs
Hr0ed2aN7s4pADH7bPuE801wRoNdkPlnmWdBGXccBh5xTaDNZwnf0IdRWKXpBtn1
Q5eodk7ciqUYDTp9y0rgtw6V5ogt09o8cISzgi4mP4Oeq8o65pszmFzE1zozSE0I
oGS9ZMbxWxNMxf017mfCY6Noe1e/Rk3JcdOMlfYCSvXUANBAUbgMw9TYuoqojLpo
TmXbPpXhoqmZvF3HackujebIz+PaqAjVE2Ra79h+3CqjMPqfjIdQpDFOknvQq2W3
GsuRV6pptKSJFGHV73eQW0+m1ym/ooMANT0GStwLDgIryi1OuYLjdCveUiIY8FoE
NVuazcihgI5n0Z7tqPSpZMMPVeN9bpmriuCGwujAD50z5sJcFM5iOeT8t1ndeLBg
h83fqa+uCR5Q6AYguPMfUUR+gg7Dv2yy2Plt/495sfnFbW5o3IhEIdHDqqDL1Bok
42h1ElEFoUcRnPDU6AaTXIDpBuPtjKJjDXWWkaOSJ1z7RlKCakLSAoIq9Y00ih+Q
jzHMqNoCJf4fkilJ2EJQzCQw4zeb8rsIMCD/8gLu6Rp8Gi1Duw++nbirtqWr7NdP
6WNwoeeyI0IL6kqDittHCGGrCZX3b+h0ZJ0vG4dNd6vM7311ieesoMWQa+ghMl2d
/YWX82ZFYNby/Yg2+OcB5E1xLKi5H97OU4pt01RvrBDsuPWIM11mCfS39+vYEdYy
SU7cUSvpZfCeiO9OBJFkVm+Iy9pdiVV/TkRz8Gk1cUmNwCXyodwCezzK59/erlQL
7BtBd1Zlb2QMzeUVdQs0q2wUIzxUVDR8FrvDcNskWxfEygdKFOpTtnardMxdpx98
K/rKmnuxDPHEipWzfB8nyfJEmErH3j8L4sG5+9+0qVEQJycYlYNaWIOPItwxhVJc
iE9GsWyxoNjkDFLLyMxxY0J0n9TXnDhsM7NHm09PR9Le68hSiAV1t0sDpH0Vx9ru
IggLPbOaB4Wd/rVw4pJBw+I9Z8+tMFi+4xNxo/PKjliaswynUIl8YcsWzuwZJKei
LvjJ/tnq4rrOFy6uZIgvbmS/t71XihrF7exZc6xQUSgbyUN+Hn3iRNbzR622Tw48
qQ7fhZBwGdM3rqHmTtoNxLSwo45LmeajnfBJ1sskVELSVxnJKmoKQvqUUilAQEtj
fqG9GUXzeSQTL/RYGaqv6GT+OX+SGTFgTxRU9ry9TKH71h/yTGG+lMnYZnmv5sSI
ZElbpQ671YJ3xe2dCpDtaX8LVsx2SCZlEFwKEJSrQjRbMFzaBzU9IZmLjqUcAvjB
wrZwccZA5M874GfUzwy3mXB+ehj6d0Jloodfxfngg7wguHZglgKcBapcKl928hlu
4JNeNMtWZYtdROE1A02HX0CVUCHoUSomIU+4JpXfnPXEzUyZELUfkQ9PK7cR+FMr
BwMsmPgWytEwFjGpNCHwHtlPo9+vnlStJYghFphlxiWNrMP/TYoXOkmXzX9J89Hr
NZJY/ZeSN6RsJ3ojS5cbfv51iI1XJwmJEx3CZ151S13pxMxuHtXAH2791ULFtcur
f59GOcPdWDE9oKAmM8y5X/O2iRp5cvO4i9qFntvzEvVGrcC4ljIVyJJS78coGkhH
2mh1RyVokYiSX0mUqJoToW+ryobO6KgZ0abfitco101tL13GmXA8mv1CkYiPX/zu
X6va7tIyUiZMvZFMrpybLY9jjKOF2C2iIciJFiwokMvVUcejYvOfJylRLFxk0EW3
hgg3jUlaUXNurrxTUWTEk3rq1JDC7DXSKi0yBdgS7A7sFVNT7CnP53ucAg1RGTa/
YhvDMFiogqJNJxjtNWQO3ik4RUUmXJfag+f3AJciXMySamkZFZvvMxu/PODHLJdN
vXQl6IuWbip9AobIKY4D9s9FRpcb1zgnShqL7sLc21DlUjr2/C8GwUbnExw0ztjE
MHVRzgvouI3aK7lzVTtnYuTijgqXBwA0AaRuK59EGx2HuxzCVCarDGGUvmq3Rsuc
O1kpX+ZuVXj7xFAqiiq0O9AiIUgizKQMIig0iD10mvj/RjyHHURVxStA5LX+eSZ3
ZTtZN2zOr+mVP9Gh1HSZ0ewpm6bYdOZ0gFCBcxNmVuBhpsHNjQrMYNuH7dprNil1
OxQ/4L7jhGB9PF9/PyVp1mwog3jBVUhoGOMywAFNx5P74cpmrwgf/H2gskFFRUXY
+Gq56MEA5fPDZOgVxnEsMjVs0N/clv3nhyhCiQqE8Qc10tYo4mRG1Zqz7Z5oPT2j
k47UIYIpbTauP48io6qKemAsEWG1+zHwbjPnXJhNx+z6SfR876dHOhyXAxysxY+R
BWX6kY0Ffv8QV3ibchaLnT3DzFh4eMa4LAC5kg5e1PquBsDaEhRwBfmUkDlXOWrv
mhpUpYavQre64eZK/Xugy2wbHgzJ3UZ40IIbtqjZyuEgyDGyTfNyAPS/VctbSg1d
6Vj2kaCYwhJ68cjFohxX8F4TyCiC3Df/VEmSrijozVzpyEaS9E4u6SF5QKWoM3Gp
Ar+lwfyPFqDtfl2aAJRQh+xI5NDT+9w3zLgaze7JSQez4SpfyxDlxOvyYqlptsw9
yNAaz3ytn5Z0nKz5OPJB9zU8heYEEeh5M3PNXXjqcabCO21/LRoTIptP69I793DL
gTHlUy5ZgZIBRLPUs1/bUWpTrpDB0dojQocfwL4kDnxQVE/iC0hHGoNoh3+lbSf1
vbf3c6+UsPIAf+MBIk+8ZoLL1sSEINT/nZkzi/h4TM1d2MIDrzWmrvh9zizS0BYs
5t1No/dwRU3qQ8V5gK7FA1vz5U+LAcJKFF1rr4ThFAVE5kAy6HVH8KNQuA+ZjxlT
kDt/fTof8jT2EXwGvsdFKUQhpboEuEcKQXWAwQQ8LalvscHXIB92kF8OG9cCWBbE
SPywFKN0b1EMauAmhhVXTHsFNJ5kx0LMKRJw82VWSVWfjt5INtP8VdGUaWZTA9mY
oACYgxN/xzoxjHsbHGA7vDnoHB6OxY7x1fArYjlx/UidVgsaoUCereg6oryu4ZyH
30XVC1nf/LrgPcyoxgZQmicRS5dPjzwvzx0Hy+mMCCaTJdLmp2yNkyaz164sIUyo
vo8Lb8ZaNpmdyBuc9rhxgjPqrQTA0F0eCea9Midh92h2BdP0R7sXOu56JTC1Y+LX
tYM+JMFiUQX8jPwDkxStWlgdTdBrQOGocRwRY97+VuPygGqPS2JfCSnaDicCYKuq
5zP2MuXBN5b7yS7BWNoa6Q+hZjvyNwduryWpcOqQCT2xiBq6hdquO4UIbgHS3sDQ
qXLzmpZr6GYKF5STFXF6zuyxka7pNHUNioKT5UkBpJnP+5N6SVOC4EP/6zBaXq2I
2PIfTsiAJon7PuZnuTKmZ2svnGWTkXVwIXs+beQzDj/VJvp/S8svBkdNNwxiy3Fr
vqcpEiFq7tN5W9OdKpjuICc8Tz3MJNB/vfn4EFAT3Y+P4osqUvGPvgC3TujQ7rUR
Z1P9a6S2gPUxe25e0LPYJ5tO8/Z8wc3I7HJiGTs3xBxoLsgG9tiyimFYGPQhbqkM
3QRX4o5U79sVbC5qf2olwey7jT4ERYQfSEFv232gykL3td0IRq/g9N0CLsOYe1zJ
lg3MQGRpDEQ5oazt22dlFuwLcSbto2Wi2Byo3UdJxRsPEqHFIx+vC4LiCSrXPFqq
eWZzcnFJuAMNhd2Wq3jmD5mA1RaB3kks3Syj3Ia+nsjoWEHjVdHAtma7n8mJCbOm
MKbrrOo3IqsPc134NrSUzCMsE8pd4wNPmx2v0yIH1VC310rwMDest8pHHqK8Tb4i
wk5P0s0Lh/AEO8PybvjT4yM85v4I77f5arnnLnzT7xAfQqA2i+0T/AkyCrJyxngd
U3iNOz4O6IhDYTQeRFQz8GFPBVOAlHzechOxgy204CZ8gwKavAS3nJJ/18CLuRe4
VzP/m8cIsOzlMtDOOyYAQ0r8RX4/8zA+Euzp40JKJmti8B7/hg9jLdREG9jP9V4N
etQao8uvhJ0b3MPlbJj7OPteARO3Mq/LPYrIjVAUkqpx9oEKnQQWGdvdtt50Wnpk
H1ZPNXt89/FcuJbxQGpc15GgbZ4QJpC1JbrHyQsD3DBPeR7gr/ApEl57wtw/QtVg
T/vLUPfZABE0vlEJh6m8IKBnoMvZ/0abnX04qgI71QLyXqzMr3akaqLDTe03n8EN
nP3XXChgDu6hufgKnqPgoeVME/2rUZQCWw6xgkyfIL2Xk5OTUFBdkfoqFjh4RiAs
Ornw3w4heIJmVpGZG8lixhPkby6M9fVWwIBXrtquPQkPtYz2D/wN3LWb9rEg4kHW
oXpErSclYSpfqJVvk6Y02Pel71w/fv3U775dee+rgc9hdNTLG7eswchD/efWQLIH
1+ffxehHmFFL/nyGIlfdl+z4xz8ehmWpGgMbhAPNHZ02zW6mabxbQl3w/FA5nkXM
nuSkcraBjShTa43BjeWy2POoRbQ7oZI3giwA2cit5rMPJ0EJgtjmg/jLSu6/nQnf
RogfMoZApbybzNUv4rHd9YcyWv6AEy98q4UdCdAi6tfksE3+AOkPKlXNFdy3C4ss
OuyVfPca6NCwinmzevuKwmm+n1fda3MdmIw7tRnbGaR3WjI1idVCf0OXGvcujSfq
SJJhYlXq+G+MOm+uR+N+asfekBQU7ffzwHzMSkd2ZkyXzfhP70eTuOrmVbFvL2Dp
+YFZ7/1msX/ebX9eznK9MEhmm1AuThErUzXDWTGqMkMUrGGTDm+9Id5I72pb+7iq
DnrI4+5uh6rv/MbBiFQoR2LrA7d7bTu63EX4jL4gEP8+eUt1i5HohxsDpuLN1Rzb
EorKSRC5xWrnYGnIm6e5zqSbudndb64iqXWsR+QqX2/3wQ3er22HEeda+hPQWU2I
UZ1Gdxc2mxXthBb/UWduadfsKqY1zMGn3uEUS6bVGRVLKJdFhMvKB6RvlierZsaF
Klp4Ua8Km7ciE6aSKC/bCgCbS+obIbBHAPxiOVe5O2NeS2+qbfV9t/jmBpy/uq/M
vNnOWcHp0PrtTFxd62WcFyp9kvL+C7Wfi6hKUZKw1qKUzKJp0C3bK11F0Y74P57Z
RsowSFYH1O/ido1fZ6dBmYLZdGC/RGn9WuO4i5HWvcMzKAi5fgDyvinmw2sI4y4V
uiP5CtVms00nh6sO/xGvWwMgdemk678dor7KsPzGFgyOFXRTf4CP13KWY2SNkQDh
KvKPcsIuz6qExdxi5C38vfIghvc8JAVF0JmjZ/vHex3dPONOzjQO2o7aKZYEGkdv
aFs/7ST3z6vpcuK9ln7qkafRhYXM2dk5judKj8wohZ1QIh+kfmlN8v+wvhisd62a
T1AKuNe5MMT01hh9k9KoNxiVGZSc85feYD9NpdeV2+xQTPOZIsaBMBLiCt1S2upj
5vnP/C7FU/TQkuCX71zVMzbJRl1d5i6IeDS9WFoYcIK4/TEtKykTJq6kL0cLCV8m
DkMpPd2mKfNI7JtWt86SGITKdK7boV3xVpji2f3gbsEt/52Q0pw+yIn0rXKlN4sC
FoEn1xDA8cGUcKSW7jolMEH4JnuXMGveDaI9NFvhAfE9ZlU/yGhNcdY9PHDwMxzp
PMa+Inc2po3eogaAxqP0Rs3p79BcVuaO1rP2tIBwQTm1h6PnOqoT9YZeCMSs4cSO
zM9SYs5V/BFojiEC5E8ciumIn+CzrDD8FV82HY0yutOn3t5HF3Wuv73Z/0vp8/Xd
JxYa59WCw+tMY1o/vOtedBiSfvqJIj8H4JIbheqzTm2Nbx1fTgEJmOmkTcaD4CNh
/qcQ+WrQSxC9PNyj1W+6qZJYlM93UdBKei0NDKdQ4gDdQo0b9HGqF3iAfjLCDhq3
a8V5fT03cqX5wLGnu2xibHYPOyJvXRwqNqy408h1KkxVXaz+VXWUdt5rWkPtCKmJ
fKKI3tlIyv5rvq4HajPPgAql5d6ezTlqz9DIGH09V2vPGOYAaRSExLfyAtATCOib
OY6sQx0KTpwbJQeRN4E9/JQsp/805N1eq1EBxCkTQjDn4CisBRhHnzToxZn4zlZq
PjFvk7+8CpYMF+5UEpt8rX1JUKgru9ImwzIKXKVDvJ1jQECcUo8A9jWzeA4Liev4
pVR1bVBzgQClI+CqMHng1YoKkdqE2VXH5ibSnfFQOvrVX+DYmP/ue+RTOpKXpk2u
cmQ7GuG0Z3z24fqxTA+oHAJKKKU1f8412GgTzIfeaGsgWrL4QcUXzMvHdwzbCfXh
W8YT8ZTPVdrWXzfKdUPF1TRuLZUWZbKqmxkS4SA7EjexNarzA1QBn4MmVUd0Yqve
PyJd8oA8bJI3SDiR+IJYBzaLQjX/eZ1F9s+7/6K05Iqu75XBuCCqQYT4wDffxL13
1KZB9pWIGmWCTSnio3zkXehbcFIWmayaCVvRwReRoq9mmx9mFajuqlMBOeh0jjkK
mXzPmX2ecIQoQKuQPrMGoTLcKH80bvhRooSuHxqibivw52TLYebY/p27znIrTm+O
eP8Z1k1zPSDq7oWfN8sNVRSiIGMLt3oG3zBIoK1bTr0bGxruDERDkbQY31rYlfHp
F9Y0CtnfSNqGx+T4lTGhXbwiaiw023Oz5+uyOSnjjfq22kaU26yX9/5h6mmR/SEh
Sfm5v9gBmEDqjhUEwT6KMeHOqzcVUayFkXO+F1o7cGuNJrA6R0O3loCVEsPAjI5N
vBPIg64dG23PjQ0r5lArEOIJXjRb4kCdDmFZb4gS/Pks8AHWOtHXYftOvoBCQk5C
/RsijzQSyeaDPiEJkXDVCxChG+5eFPDzpFVj2ISQsX0JtJGNwkeEF5mt/o1q2HEK
2mLwceA99v2ccsGbiVrfwI3Q5iqri/NNuQ4TJKyoXHUH2m031W6LTbeNzXwXxzqv
o8M+MTe8ui+NM8RJuBxr2w1nIVxQ+9W5VWjN8COg1HuWhtFdHmyhC9oJt1SifOVA
dX70mOdHWJTuGaMEOlUCa4urwyBVDZ6azUngm87qe9gqRkrukg4SocDuIGSBihWp
mnoWh6qxS0k/M4AfCEzGZDIFW4OVyA31PWurJHU7rL7NoHjzQvnmsYZGEHrUx+ov
dRursqahhm1ZyJwcGOHGfLws/saksXKuOwdlGUDiWxCMj4LZ+cYib3AjXByEHiAg
Fzi+ccOdShnNC1Jj1YTrEknA79W+CfLG4SnjK/KAWWfYY/ahXxi0BidfYQr0364L
JeC3Jg3pWzg+zE2DGKYnlkejIPBl6rzpgK/e39zdV4Ltu7pwUUpDT52JXAkASxvE
5CsbwRPVmNsoJ/pRZ61wRxEVzmib5FybPCOWRnU8Y8NUv95Ru+Gz27xE7oLV0gnE
IAWlVHQei4ateAtpNpniLGAOzmwkh7nlMraI5G+5IldSjzaevz+5KzIymdsrWe6Y
D76o74uLh8AMX1vmBmnnNmEniIIKhRbuWbrG61gd32dxDcD/0iSR9BfeIvh7UUDY
d2XVuZ8lPojy8J1UEDz7gJLZVymFsPjLux/1uvxuhHKlk3E+Z4MO7m0FRFSpHsL1
wbJuzYMKsTgmm3DKP7V0+zl/of9mYhrF0GbBBSkUhTtd78D2t0E9oQJtSa3akMW0
Q+/108pEEAQ25vDlz/r4SvX3XceTlOnzSnAj2zdSKbhz944NB0Mamg6YShNy3h9C
bdMmxnMqJppUlnMxtH96Wt5PRl0lqG3y+vSU8PfbIljM/76jbDgSjszffIyHx5Iw
E9Vx4D6hFlnP7S7bFMsxTmk+xhbGw/d8ZikatvbTbqC7p2r2ikAg1Nqcgttf/ySI
oXO1+XMMZIiff0ObiPmecLdVz8VYAb7mgUUamxJVi3oZ0Mz5ikSRU8z1jqfQnCWI
4HRePlFDZiLpOacNp3hUWo2gwed3uwQuK2w78PSxDBWgBAyz2d8neP3yyMLZoiIw
yobyIs+vc29ypuTn3qnttsnHkFFiLIxiEVOwbZglPUfP+x3S16EutPoKQVmtsK5r
xsXGOD7etHjccBO5KsAquylyGy7QCLsdCldIGheOkUFBREPQix34ycZgnRwFo4kA
DSxpdeSQ78d39ic8iREa21UiXNXec4GcjtqTqKjCccqT51ESYajIiDlYRXEQ2FtB
vQlOJGu5agUMsxYeKn9LZ8QvQpknypE+GXpanAdFUB/3tWtbKopo0Cg9Auz5cnSd
slOe91ygBBBUpv8t6W+WmjrqvoCgrYmRiXGE7Xt3iAM+HoummAshhMej6fA+TqM/
JiAswqcuHNL7vHEAn8e9VJKDgJowhNloHv4SfkIfZIFXrYYUAgOeD/gZqijZ1ZZF
vWkWxVpk9PH0qK46jTc0EyIK4zxwNS1oz4K0TZ9X9C/ipxAkqofZsqZIOh2u3fHg
GEPYhUYX5PWcEN0kl1pPugzwVOqEJLFo7oO03R9e4vfNtRB8UmXsATrsngBxDGmk
/I5qLpmcGBjynnsbQXwAgP4ZP8D7vZ5FPYjcWvP6TTnZQdWTh40JXANLpT7PjzSH
eN0KIppAjp0Pu/JKKtqa4cQUKf+H0U/lovcOZ96VPSxwb21jqhZVTbWpGV6XxiSK
Pre8JRJXAHIW67OhgVyUAmTnuIwPDjv9e6Y95TbpUeGANmgd5tDp3EBhJ8O11CGm
2rVVJXyJJ+yi8iD2djcfIkh0DyvmaFi7gH9oU8EEAJK69NK8bg81A7dozJ34R0ac
j3wPdS0Q87iRhVFAdx70wa4lCAlNo8bF8bk20gakAOcQgsJp+luvRH603FLqtzVV
WDi8BDqKavxJFwGBr2AXKbRa5Vryq2qO1jRUs17BOvkdHtauDL2RQSgRzo29VvGt
sI3pkDXPQgHFg20Hzefj2iD2myrEzjoNIgxFYuOdXYol1Phx2xjS97A33lO7DXTW
KA73VodDUfn/PHaMBAQ4HH7YAvgzj6fTWTBzXxIOY9uLx7Q+oGHfF2odrjEnlZv5
5lHYhqH+kXqPPC/l5T6rW4KY2hQD2xnPZ+Y+46snkl24HHbOyUZupm1B4cmUNBSa
8WVkKGrxy0pF4Bk7weycFEE3yQ3ii99QPKrOIIqcnRzB0LsrQHCd+CLTZgPPMBpn
kSSdMQWLmiewfQOQc/sh42L2LidTpcRBHTW98eIHd7rtG0fLIXdn1MIGT+VxOLEd
cWCOTfflH65EBI8ICq9HSEp0VJcJet3DBC9HECHyt17NCLmKoFyHbAXvHeX/Uaca
PVsIMRkkzPDXe1fqhHyMdJ2jxa84fxYKhot2aoTCEMh4tJMCDM4Z/ppzgNImOmS/
TKq69lT8/8ld57tzhBjTMykJEujCVXolU28V7Qva/PDpnHwuvkfyM0UB9UTAwbWX
Bkh32oEzbIszJDqVjnrhPHJaLhPFmWN28t34xHMWSKB0is3y80v3ZwkC94a8zePc
mzrm1EbqFFyvsvWaEXpVaNTXW6qKUN0IU86g6/lVkPlFfy5Bv1X/C9n8rLzwCOP0
UYIS6cqQxH5o+p1e/EdYK9NQymHkKb33aD8nTTTU1GBFZrioo4mhT9jzL68ZYloS
kbXFUfguxMQWMBq52slaIwXwq6ZKR9RBMtfvftoma4Y2P2aZVHFxC2i783dJH/bp
S4XQKxhBen5aqybdmZieiGG5kZ6ysA1HhV6vSAoAI9iwYPe+1eJPjcqahhQR7pCX
xOjSSMsAHy3sq6FtY+mZwhn0/C9S4j55MdgizbdgnUPnse97N2mkgUWw6QYJ14IU
9uE8Z4oUCqw8U2VpS3h7qWMt6HLdIFzxL+6Ch0ZjKwaiBUoYFITPJEBzXezGm23J
cHCB1XpUFMs0dq9fZVWPg4VrN5yCCNQjSEnKTPfMUDd4p1xWgT7EegVt5cscGEvc
2P3Vz4mcfImAvWTh7cixgElU2dQbicVGZcOYqj+4kDTzcHP1ESKdHjlSX98DBR6k
XWy/AzsrvT7QC8oy/Wvo2BjhwkVKs6P+OK4zgml4dPBHNLfPtNLJFL3i31dO+B7w
+aGdDZSlSH9F/kHBeFlqnqolxU2bgHq2n9N3flIk06cCTnfDQ5fJGttZ6ejCzYsS
/HH0RnBVDcMFsxSsxuzptJ40Fv8qyrRWUazWVG0HdWqjjk9hNjbO+RzsUX6J3l0h
b4XX8wQclpnfWQVcH9IQCyvLrdS2p/RyfXF5Ti5A791+/dee2Lc+quPHBoWvic/k
se4yVQaDTeHbNBmgDGYvTI26nZS9WKdj8infRSC91syuGCICaOmwluvEmzZiWF06
4oFHPk7flRJ45USR9cxcVe75Ee1yunC1B1pWAOR8+Slw0NLuzwfY9Gm52I6KoUfH
r9LSrV1ADeQtfxTXGOeG/RUjbm2WO5swdZAxLZuhcRtvFc1263FX8FmgaYuDus9m
NRhT1h1ixnvNCBR9k2g+BW2zapJr8zc36Fub8XgpKivmGseCcSKQ2qIYIcWAeF5C
hHEUBhwVRUyb0UBw1kH9yB87OSZb6YLTcLzQqEVV4HTNdapVNXeUgVFIGTI4Y3DL
/tl566XP93thoMi3FZ8BgRziYOk7VXNXAg3yalkzA6UMH8/5Outvr1fJTJzXtURP
/qJg4XQrgI4T1UjAgiVcAwydMd+W2q+ZDPcAiVyOWR35Fr5TnjHE9GowNItuaZdD
2cmQDJcLbmPacylJRHVQXqrObvVCkCoPE7u7mIvAuVBsD+uHZur6joVScGgeBz7z
0qe3tcxLpGCGEQ7V2EOpRRXE3dJjf7sHSm/lyJQJhH8YeVh5Ri0WCc2AI1OT/SQ5
yMkLIDwEffnghedzV1L9OIpE+YoQ8mHXelC9UrQLPI20VkkP8t3xRb7FOkQZHsPZ
pSBRfDydJ61mr98Yc+hJb4vLqs9QGph/w+aEhnFl1/WjTVntmzPBJIV1EraRabco
YYP81hNnxuJgEteE7c12Ov8czeh8CEGDZLO3Hy7UWatCbBBmr6QtAN3fqfs0tx//
W7NvqWQgq2IFhF4yV0bykBbGtLgLO8fjDsNz96OJHhzWsGLrxZxLYrrWTUf8FfTd
QjQrVnkZozLq0Iabdrw9lz17ZtrDJu+4O0A+8f7jNMLJXQkKrxGET1dmwAogjR2x
XEDkeMv259Pk7hUu62sl67466tzqRcGfSy1bnwP+V+RWpDY/WuOKz6G/3aoTXknZ
DZw3ElZPuCSrA/rGl2lDBqGoi4IgHA5J/A31NQZgHdY68Ld5cvWiskqpuZXDwmSv
AXMuKY1EVPYO7VFOrAW6HZzEcktaxt9KeFqTcbrlX8ihPqG7yla0p3uqoJsATVrV
kYlfj5xNMndcarK96HHteyTvzrBq9WE5CGnpNZ6bUHGSK0kYKIgE2YrVLVnnplN5
XpjzzSIHcn7IhnaA6eqTIYlIKBYe9FqEi9Qro/nZRjaYUbW/AyOT6BB97D/n2r7N
XgM/VwmZ3eDXW/j2GsHTu0ZqJsESYsjDJq3eEddvzyrJSQy1hbg56g6lZ4Zq/9k4
t5+qz6JNCeSmnP/Ji1VbzGTXZN1f2Bc2QVotzv28H74VPFrY83EbdeN4x1KCTuwH
hNey8BGLJuBaixMvEOnQHPKuaDtbeE+beNqG/ifql7IotlGju1tqcr3oxZPpaukp
9ZYYyQ2DS3BnSk/30THcE+SXJ4dcpqR/wGOep+O11n99uP4yNqMh+OXiue4J+auP
ULpbHIYYNxSjIK3K8ViAShsUs1A7CD9Zz6FBQXR4LjEdjERKlF7fs5TWiFdkgCHQ
V++fjqAxwNzNmRPfNA6/0N7xe2giroxkZfBu2mAW/46cI1ADuH6m8AX+jF88pbyj
JW5skHr1SgH3WQV2OtSl+BGNsKfpC+y5wvcLuEzz7R84/cg5L/WiHzgx2gYwu5tX
/qxFPyWYrtd/tq2MHfbW98hCDmUErz+IJl/Fh9CC9KCWJ6Wl4QdC8UuBix1Y/Ba3
4TmjGArv6SS0ogGgB3pqOogrfF7Vkg+YM6PADjWx6PrTmrGy4O3uBXH+QC0vtbSG
FvEMph/tvI062Jv3Iml4ugHzG9edmCkUHGomyEMHgOoVzCD1w//jFmDcc/iv6S/d
nxMbC7kApgmFND9Nlxmitd+cPtZNlCLcF7EUCVhSIVT+ajOrwvmEFv9pm7Nb7JNO
AYark+qK92bYrFguO8l7ImD/oq4Xepdi1HM0IEopL+3RpVDFAWXZ1Z/Ah9IWB8Xb
TUaQ+zz/eOA0yJIROpW6wX6FhKaINWpq3+mVyVO6pDHkbaZcg2tXFP0zCKOCFay9
7CV/RMMcCrraZoZXb114SykSM33iAhio29rJt0It3rUH5K1yGbsaHjiWB63uJxyw
hpwc7uMpbqL/07JQt7PmyG4mzkB44wdeQ5suq3BEYUscC7RsNv9mnfcaa4Uix3/s
PAwbaImWOYsoV/XitpLuIMUOij1G5b62aJWpTv0GuNWMh81giwkqlhj9w2lBQu6f
Y6ufqmaThqRkA2Th/57pJjRhYUquCDVsJQmkjnwqHRd+5Fu3FPSGomCSgd3NFcA7
hqlNj5oR5muOU4ubeTYD1rykccyRn1N5LsgPrD442xmisMtGlkFJ6lOoNp7w5B2e
Y4/uQ5ldUTSAgJ/sjAByZrd9151F7q9M+nMoN7WM+fqzpxNTQBh92b2vAOXJy7yY
xPbIVZ2IbrSDLT/nlVjFQ2ds9OgrNdGBxvyQoQJu82HI6c4X6Q2NIpkIJtYB5lBJ
CLAwrtZdhGagbxTs/w5NjrfnTYiKTtQewTR5Jy9wLzGlT8/m8Q82Wjix01wLWE08
/x6Kxy6szFOeyM3xot4/C7qwRqZeNkHaqzsGXkmI4k8ksIdo8jMpMlY9ht2qTnCl
gaJwz4u89R78SNs6Ow0UKoe4b8tU+e1fNpANI4vyBuIn+A4SO73yrutjIZMT3+5r
gUvDyAut/9kVXUxk+qh9AeeV7A+Pkx+vESdnLOuXrmgWzGoF81La3kNTW3wOCCdV
KeVaTfKFfYbnh3vY2Y+bJIGQBT59J2thHCHXjnp9+IOGtES9lVCHdCiB8539IVWx
iSONOh424/zRWgMZ1GCbxEIguWmUIzGIXEX2H6gmwFygMyMkCFcovHxgJxypN3XH
iXa1cOnyKaQo6llxbW8CM08AdqogTqBrtosZ0NL4O0KzjH/JN7dqiu+cRQXl4Df+
O0JyjGY4LW7XlX5nMu1Mw1XFegP2cy+rd/UkYOv4tEsLn2IYv1IXNe6jZIvH9xlJ
ecSD2AcTeDqufWLOLDkgGai8JoL6e3OKrrTK/KXT7fRCRVyia5axHQo5YoMklDZQ
fDp5//vN8bfykYJWPQlXBiu1xDe6aHauabD+hntfOZdwBFA7TsesyhMWBf6Jf3Kr
s8AXSK/LRJ0ZMWfWBJ8lsytOvVv8L+UIYCpYht07HJd/qdTRC0DR2GWDEihR5m9z
0sqAkKXZq/EAZOF7Eoa8zxoReUw23hBvr57hYC1mgFgD5Fza/ZeWYqVT0eltJvi/
S26XoERUhlW9niBHDlVmRLShUD6Gf5tKJxi7yv15EKITpllHiCCGHs27uvBHc702
8flkqh6X2/f5ZJnmxiEqZCVxni9hfPk3YNzdzeLJVsm5qABnLJSsEJIaTxEIzw2f
kq42eFyVl+C8vvx6U9ZcRQAB/E9YyYHp0iFz4qcnhU2yO1ud8b/USWyXZugBErVQ
j0vx7Pf7pcIO8PLO/bXjXToC1/TQE/svTTr00Km2jTzcSG/Lto1EG9FK7BbY2IQX
C0tKJ/SIXh5m88qRlUdVdlccoqSTn0cr2tdn9aF1pBGZMOiqlDR81cduh4TFgKv6
6DjIOmxyPnztPByhQdC0uUDq4U8IcRhIwXk//TKxkS0Jtk4oGO4BwdarIgoy9POo
5t11/3SIwZktLznqSTYxX24p0kq0aYrXuN0zgTu+g3fHq+jNBWuWYvCBccjrHY2l
MF3vBG2aux1xVBTlQzfwRV/xJvAwSnOPHOi+JPz8LYKpv4I7rOwdkd2sqARPRvDT
OY9Icjyn8CZC9+2IwScpPt+DZFDqxVk3jsdohHBdLmhJBoHWt6Wr9anBoG0EYuRO
CC65HeJr0opwqUDytjKdFLRdRZ8V3IBIxU4MCba1HJZ7MfwIMN4cRtdRvfx2kKTA
KVKWC898mCtypL2ntgPKa45csHRoyQ3IabyhDh7JQC6rWu7k7eaCWwLESXKLs8ML
Z1TB73UvE/4cngqwGKemD7DJr+bZftKR/XwYT/KbF7fpH4WCHNYNlSA/Qdfr8qDQ
MzoZnwoXggiAO/aUMdVbGfvtIyrYwv87U8ddiPwkU1cCQ5g2J/hNGdAWuvi0nrvm
jZOxTeeH8IeZzMSbKGlRcaKY46+v/ZerD/uhUzFUoi9qY7MlCImUM8afwjNLfBd2
9vHW8Eu0+6edu7Cn/X1eOtP1Csxv4BC6ASBv+kDKz1GWyBjeqcDXqhYWTwIuyORd
U/WwRn7VqvsbyoImJyrh8FKnd6/S70I4DoT/ZAu1VONfg9rQFt31XTg1vNynuQSa
sy+6dmW0TaqfJXjEmiZvDC/3Ar8uKYLasqk3m5qYf26hFNME5CYggNSoNCZ44pra
AFeXl5kztnWNvrbbCs01BvW0Y38NzoBSRp2omEJE6HDeAz+7L3gUiybSzxq7J6iK
aMzHEbSHXNmuxdkccVBATW52fzvEpUVGzLRfptePcR38ysEGz+gv22HurccY94qY
NvBlfWKfbXGDgPrn5PjkU4HlKUJ26IMdggvCWMA2lgXoxcPwgUmx3yicCLRC2RjN
8wcbloTHHInGvQ/xfF1jJiHpS9/JLFcal8RCvAFy4IaoouZIcM9wCA18noxbIGko
FGK3s6/Iy9qQNpNnfZhvt8McU5TK5AxCpy+rHN4vcoB+j+yblEq1nvEz4fES1+mA
chVur2X4JH5v5k1GNN2MRGxiGMMUrrbfDUw1I/NsLk6FRYxljRFLjydij2LJP0Jx
0a15v/ysy8h68ic8Y+DWzM/PnAd8QBdzciONUP8J8C523hNBvbEvgsS/x3oRNgSt
G7W17qFxuSFRk+Fqe8RsgfbnNRsxqd0Efv/aO8KAOvSKQnBJtEz8DozeUee4yFZk
BQfX6vofrO5J2Iyju4Bh5ZMnd14U5fQPa3CSDE2TV7pKTBnS6tT39LkbpBsgZ8IT
y2LtLiYYCLVQ6tsVFogUBf9KGvv7SE/XiNSSIAtRG1CoH+hLupddlJSSYAwfnPk2
DOl7+b0PqtBelkYxbZd7LZ0uDDtg8A1+W8MT+6qV9uzgwZrxzv8moBzI1ZWikpCS
bI1omK6lPv2dH9Z0dhR/hXe1M2w9Wa8+FWGhA002boWl/AgYfljG10hW1MVZhpl7
zWVUz1/k3XT9XrHeVXf4iCvS5Jd/h3LSkf6Shx2ctJrJ6ej05A+aypr5z9pASDkd
7j2121MMcmiDJZMIDvqepuuvGavVcem0Tcz2WCIXzOcfH1k3X+W4WVaNcsqI6Ftg
r1p7vkvf0qptha0kFeYC5Wrn3Jb/2VutX/rqwCRci440bkf8edSqxay48MYOHTEY
asXRDSQpJXqFg92qEnG/pwkBZMXVNETk16qbkG0dfKaRaPzsQN0QESbIVkSEJFiQ
PViBxxhsOZG0Sr/JQ4Ndmllpl0sj/Bb9FS7h3OXumyXL2Untm9KYzHafAFm7FEhm
rWDwpvijXpxQdv9s9HTozcHE+UdCUU7hyZKelsUw0RLUmH3g6lAplonOTeo5Vd+C
ZSSQVWZtl0fPHcGGzs2yrO0LyG0uAMP6/NcAO0LXzwXoog1MWcbIwP/qSBb+xTG2
cLb9nvUNDh7/FTIJdvApknJ6P6z35smAbGJGDUiPz6/C+aW+5w4LBZlG6axd6cqQ
BAlVFr6fx818xaB2IF4a8kaCL9UFyLvqRNUC5LGQUpk83MfSb//OIKClG3S5R2ui
iA8qsj6rVZxcAjJvAYIXurRGbqLZNyy4DV7vUS03jd1shjkaSU8eVwBfvLGAkG8U
pW3DGcKiJJKRCcqafmCc37+NzbSbu8ouruNnUU0nAil7KyECFbhluoUKGYxfQE+A
xUQrn7ry4oy52VuQlKHF0UrE4mmpC6f/ir5at3k9zwL2STN18Btyw1Yb2mTYiRgc
7sp6N+EuAzq14EnyQRkbyymIDma4DYjYnJYQRqTPyPswUhdS5JL0ljgQLIacfEqS
O62aoYLpyEhLvRYRPsjE6ieJPiiqfsD40w7EPGw1ZU4zvaKoOPhFqZTR6fMdEI1d
lb4iHleNh1ArKsDnsOeShinXYUxHW4slfMu7fnYSHoinrHQfiMZ+vggFxM0CRfM7
V2sAknQDoQwnyZ+I7JfiJiGugrKF9k4pjev/lJA1ewkbEFXVG/uex6n6WjAp9kYB
1sgUqIZtacSsbQJgcGxJcGoU3ySJhnuKGzzB4c7yZtbKWeb1+iGrL00hkc31tjtc
UnOoKKuSjmbDibIVB1AWIsxMyCOpjbmvWivDYNGxrKvRm9DJJzUu6BZAzQrQHcZR
r/HgZXfSFocJgTcLiKW3by9CN0fQhYZcc1EKsfej0FPYQ+2iBJJce/cShzU+oMU1
nfRxAav0dlQCatoWPhxYg4+JyV21jT8aDuffQ+enl3E4GheKciCKTqMoR3VLvs/S
2fxMdLJbbL6ac2x0IcdT30zjGdhlnej8RU7W+7DwFHZZvP3YMZBtUZFMXXYjMUT4
8y8t3k+nT5gWu77XvFq7a09EliN9zPY+mvY+o3D4ICwr02+n535CIpShSTyk4/G8
QHcBE1uURuGZdqSwDtUkKm46ESCfXoMPJIu2Leg9TCqpztyn2/qfM4ehG17YwRmD
BK4SENWsb9Ira4YNZJUf5CovKr4iHy8yFHnTCdqmW6egRl7HBqUDJnMBE4oAtXN/
fc2/j7JfTiDt1lpSj8Q5n1G0D/XxYr6LpFhoGMR0zNcVPuSapUqIFHHqZlP1kXVv
Cwk3/1g28ZlWbCsFKhuFYOY2q+wPnUiDLMx4c6qX5Gkomndmh9Voyrxy/qJYjSaf
cyAOcZ5Hs/I4hGjYrlJymeUxtaJqsvsYTX4rVDS1avftnDwwh9GkpG/EO4LUcoX8
dlj3vQfk5ZLHK7yTnSAb3UaJvaoxtcnwZ+oshrX+c8ByIvkgpJSFcZz6dvH8YgB0
EvAluBXRkTZs/Nz2owT7WMqcJ6Ap00oVLz9Hp4MAtqabKlJ4+atelrHUCQ/i5f14
oBA8CDBs4bcm0BJWTctoeBDDQ7KdmyJYv3OQi/EIU+RXH3+12g+8w1FGlCD10tCd
nUK0YUzWeHmO5c2kHgWS29YXAZ+lx/reJTFiZ1HSTP/sDud36KwdSU4v8C9Xdmpb
SVIkuBwg2/GwXS8C/JlSV8qp3M8NbUPlvFkj5A/bBOmQwDjtYkjYAdTv7/oxeMhA
7SRhRc3giPFB5CBlZ9MixjdA/h+XDadM8PSFXe9Ps6X+IO+FF1/3pPKh+6hiSwGN
6c6XKuHSWIhC2Uw2ksDXt3c6MYppXtxFpzlK1N2T+uG9ZoshkccOUNyHgPxkQOwJ
dKdgY/MlxiA9r001JYVPU3EqE9FMxTUFkqAf9TImcun5ZZup4TAiLN8PdTVlAgvZ
K4kiaIxWs2rbg0j+zo1N5gBPUkgD5x5KF3T7aEqKdexem6roC/ZYsOFqfeo/n6Is
evbc96uNSlYKHcJyW5uyxNsfKfikO+UxDUnEmEqdZ8FrTzncQ+GzYZ1kHiklBSmt
56V6/BO2wt8A9b9LxmQKcxHOCzyOfWmmF7m2fQ7EsrJvifMpTgdzPA6B93lhzSfa
G/tCmKe2UqP7jC+J8+5MW5bWy/HeDrtaj5LzHGw7he3g/P49bFrEepR0pBiPdQZI
KAX9vv4nEfhSXNMQfwWQ4PIYITlBmJpY/8pPJ66FURlkXW0OYuaLEbPJBWdKqNG6
yY1it59ADFfwaLqH2ntVfg38aFPkRQgWZG48VqLkANGt3lpac3MKf+Gt7le7N037
NzqIXLNL3p0qztXVWvWFwHG7x2KtpYHOTbhR7LfYxJyeQQfkI1Lp1dxukXZ+ebPe
QBm8VS58dkYlCp+6lriDWHzlZHw+GnsXAttEmBUSZLhKPpjw2+ftIxjX/FsTl+xK
sMMf3KoJHJapZWRsId4K+1aqpr8lkt1GuSMKh/rVzPDmizwWZPYDSUsx79Oeyauj
8FpJ/MSfng4x7M0VpwJ3RTBZ5N82TriLbxyD9QNlb7cbQer40PuphIGf8eupju5E
3Yaeuen/akEaD1/Nv7L32KusZFlFHdHvmnCmanOQeHGtEHzdrxudx6Iwo6bozsvq
wKUi5pcFoSSIxCc3YXmUDi23odMA3Gx/EyaBpLfIkS1rIZmlVlPNSrgkn+8JDSIX
+oXpw/bs5/8rtohfQFunyazop8ruOOFc0MsEpsrAmAnEGlR8bQNVwrRlziKF+YaU
VD0Uwsqg3zkEFXJuDacUK135cJekupuZPPE7rFgWqhRPJf5ezVBFgIOjmw2h2jHA
JqORaP643F5nmpDn7Ul4oSUr5+SzF88ocyB0tDMLOfloL/M6xksmlX3OlhBe8evR
c+41BxVg17CgRtEntQmDGgZ6+RktM5b/CjXqwoYQGcZTnwNdv1WstLXQtywoP79K
SmTrtEfijKHuuWoXfkc43FKfOaTPNqwLvtwWgAVOtPSWsARJkvYd3gzGfbKDxjaE
WQZBxLi6Ph7hNpC1bwymYa1tC+7PN52AUx4RKLu+kHWWYV151/eG/c7Vom/74fMn
WkeBxkpQRJAlbBWKLd+sWDffB4XEE7h4GSrmjceo8QZLSEEV/EuI1pibrSgO6uFu
fP3YBw2XfGN5Cr9PIdVCmc4gCsnTG5Zx4nSJMW52ASRdLa5mOLiTqPo8tvozdNil
imtIEBef3G/hcp78oiVWaEKro7DFL3gF3jyarLOc2ZtrEMih3QjrIbrgnLQ32uuW
ejS9RUvMNSvEEPk7LgHsiw4Mb7AVn0GatEkF/c9ezPs7wNB2QXNnwG/5zwtOIoBl
CAr9NHzdiHoIZos8MgSpT00+/7yaFWdD22gYuE5LBeeoVmxEJ8q/0mD5hLcZI6yF
D6tYoRCp/M6JUv9lvLu2S2e02znT07kNZc0Xlj6obstfu0u1VT5uiqt2elU90GQ4
UjhU8pg8bgYZu3wb2NpNQ+CdOYi51I1tO9aioM2r8QRdAk6MxXhSy43lbB53T1UX
83H4YpEf7cHkAuPOGj/rsnjzuZ9u+CVBgqdVWFrBRnXgTLNeBLoXEaAluPnhG3oj
k0o0h9REHoE7p2A56YLZVKolD0E3KeqYO/j3nrgpYhLA+kkUCCMikUcCGoRnVLRm
biXu17K5HE824x8u9Z7npmN/Z92RTOOt4msk6Er4mhlu3L4RMXXhwgM2EGzAqcOu
1xT6pc+HF9Ok8SiRdwerRskeWTc8Ys7FfpWsSssKDDzG8KUAaODQsgDqdjf4+jyx
IR96ttoKZ4uBZi9JanSGxG9/IXlWMKPkjGGqWhR8FGVQTnguU8uyZaH7WUFPO0Eo
DykchmkbP+ss8vXQT+AUSa95/NiJ7Y+GkrPqwPOomY7f6hRb966VYt+5GsZZzwaD
RSSN4Kr7rTDI0LzQSLtAMcar5OZ81mY2qoxsowJ14SRfroPCRtovmMyKMM87NV2L
1RqLG/1mjtWpEwhPLzLHghp3ZiJxSHqYuGNqEtBVquTJX2YWwHXPtwK7aF/T2jK0
p9kA1CsjlwBUSiV8ubh8VDQSxR3OJ0trJd8I2gWKJwKOWhkoyhBkbeVZzgjpmrZf
kjMcTJjQJoNZOXmP70RB3axQwt+5hdSxmAFDzbU8OJz7jHEhNIGgAAimS/o/9XYg
An1gTxDMxuDZmNOXdRZTq8Ply+bSjeMHlx1o7Z7nHtyQFZFVuCRmB8DvA9o1eBJO
0hP5cM0eHfR0fSPhfpNAncxagtKlIyauiBSX20Zt99qLtKxODAu4HwmQuDQ/Biv2
CySaigsygjYT9ElG1mOTZiloGNt8h1YF9o5JGU1S2ahLtlRFbJlV4gWd5cL/F/Oo
kQe4ulpn1TDOvOumfukyhoPTIzNFRLGfN0Sf/xGM+iU/0wUzmE2qUiScXoogEto7
migBDlYYICUxWA0iggiKa/hvXDZ1jASWJmT9eM7x2ZqcRIb4LzrauLDbecltlkTX
RHnh2avoREke8fzha1SjdPewC/2aBSbRx1jemGyer0Rk4vKkrFu1wAJhQHorpg7e
zjS8x0yQusqwjZLDl+QcCgeAsUW7b2sy8y9I5NLPQM+Y/ocJ71RFN32hjKOo49Ja
gtY+heb+y1TDk4Cg/W/6xVQtpgVXxyTnO16ggF1vhzmJEVHZvmhb5wlAHGCufS1N
6A56L1Nwj4smyL5EGpRmrdkHVnVI80hFR86PMCr0H2hQ1oD0nb56Cdx65OJCE9zF
gO4MIEmD8ko6cEK6Bh5Y6HP+CbHMrps/6qxrfWi9yF40SxzCHpyaMhOScZoM0s3g
cp5E69lJTXcy4XFAm6jubc7QARDVCxA4ugUiI8NLzWplKIpIZ8DCnz6yOd8UzNkl
z3Kao5XK7wIxXvwevB4CJClQFswMspnfEfTA+J7U2DlDvLDviJoFEslDO8uORohk
uN6jE9cG9ZB6cMUHUX4LpWNTjQvRjFRfVXtIG9DiSOK8mjUocL5LWE7vvKJXn9IT
LkyTEOPSHuvWnj4Km8UV/Q5i/4l58aXLg12o3UvDGwGeT07or6FFIMXok6gE3M1E
mB6GNE7YNlniUrYya3RCH0UoNO8N+O61YYewJ6KfNVA6Org/bIHP/UADZIQfoEAF
vCBa3vo4f5n+EywVgGGU+dFGeaVbaj1kGQJMPLktcTSgwD4Zp43+siu6oyerLVKs
rHglqfGmnyRxDw+Fo90Sxgviycv2xLh5+y5x2YEpHyaOq+0H8ZnA+pKPjw7qOJ/u
F0RW86rUEG0oz2Ba4oac0x166OJyOV6js29ZrpWAfifwhmQUKO9QMKWVQTbMv+2D
vtDcbO2ycNbuw38mzcCFaGEVDbuE5QbLxreEN1yuof255N5oKhilOS2hJ7DHiIMb
qKleUx7HpSme7fO7h+6Kbw4WbmLqckFUPUeK6rrTAzFfaFWxB4mXBDvibjktHWWN
N4mDSee0dhqwiAnUgHjbNRTZIrSccEyb0HupXS+ntW8J/Ug8Wlf5CA8vmG6JPW71
Xtz0Emfj6P9IaXTc35ARByqm8xZvQZKIxfuryP1/HT19KtrV8h1d/rLXsBxQU3GG
Rf6BuPs7b5NOD5YbTZrMtxCZUSc9kAA3ap25HMqbp7eCU0cj4KixqCWITjC2HJKf
YyrNTZpXyPWflsK8jsUJmKQsiqaFTxuPkBBVlYkCF6khscK3Gq/P6APqHpZRnLtQ
z6WijyUsrfHVhehKnhB18Hlc8u/QlcFpdwzN4qkAwoO/B9ZVX8zgMEX951TJvPO+
nDbWTnyFDbPGGhEm4OkB+4KJ4xVmTDixKb3qkYAKM4jh63Hh4pSngxWHsBJ5Iu5o
ZlbQNe4Pr6lkMLu8Rt55BpR8jTWSQA1Z03m5BRgQMI9Bb9SjKKQ4bV9oQjLeeLsD
nCeCPOm67SjtqpfY1QDfvkKj0XINNWA+JfhZ+lGBBGk8JpSvWkLdMMy3E+AyGkJf
jtQzxpowhQEFRY/Yl7eqeShfRT962YaHADM9ID0oIMK3varCeQ2ZeP8o2SO4w3gO
196ZQ7QbP2hWwFAX0hfXR2kWBUvgA/ktFMMm1SK4kKsZddlXY74yHaFu05uzcqEH
V/JEIFdeKRkzZjtHCMc0OUACmndfCKf2dEfj+LDeuzJGXNtUYF8CZQ+K7cqzWUp1
Kj5wdU7TgMbqids+dNx2KSYoPePoWsBlv1UyvNF35fdlr//ypYz2pZJB0Zko3E/2
/IxwgDeONXM/q5W6eZvQi+0X6vMFIpeRmWGBITDOQwZjjuVUCdgypZ8XPFxIbJ/g
VsDOk7K8+50MFUo2KcVSLJFB/KUBsNPKf3ntOPTMB/HmHrptGdrvkWTxw3upp/ZC
pevFND6D4jKdG6zOLYBDcv+3YsDJNmorkigc01aF7mYawaPv6Ad+Yl+W//MbFV1c
w6QmHaIpecGZd0vu0s8ezMEeUrrLiJ83+i2GQmHjOl9HVjHdznAQsLWlZr5H4Qs/
HayZ9eAnLqJ+8ADxUDvyr+ZOhrWnRh9NpMxIDArJfP0STCMD1yX3arIabrX+r3wY
QQZRQfA8/t4vdSO7tigZs9tIdhBUxh269f5Ppdc4IlIvOgTdzWXt92T0rwIkoQCa
NRSquSOCUE1Dwiza8uQKsVCXysjgwva4yK9pWT9OTNh1iTHZSmEnPnptBEApZk3D
cRg5/tcOw53+4s6alnEK5iOCvH7VT9zZp/AFKFeNwhNTfRWiJ/HGlU1C+2LstXWh
01KG9A4jRuEk3Y5lTR/lysE3N5KpG3aF1N65ivHgU0gi5iW5idSdG3lHuifhioWa
ZpVZbYZC+eEBzR8f8yQ8rVVwpo+npVkPrnD37fMb625Fo1Gt6ZaimxNKorGECZSf
Q8p3rI0wALvxLWtmJUK4dbQPgpm+DTGDz0EDa5AjCoSRxQL6wADNRAeyAWCyyrJ9
VximpAGD5B0Dd1hGAnhO44ZQEaXH7gvyqUEM5g9ot7BlJ13DWIqX+Q7U5IUh+ooo
7pLyPf1m5G8q/uoSPlFexwL47/gKk+NeMVHcOChQiAgYd2vcmv0RgmlpaM7D5rqI
pGaQbWvtwQ3xk/NQERmj4oLmtLxEKH5Ei+XtodtE2k6baZLxejctdn26H+hDoD1X
20JqpIHzrppaTfWBaFY/F0IcyoPO4Lr7qLjQIz9ypWU84x537eJslnaiZtLJ+qfx
1e8qZBvxrSAPNr2/MZhh5HJkK3oiLZsQEctYHmCUDCUR2rR0LAQAbhk7ohQuOmkl
WT6IoLvUGNpYYtzswsiinZzR9mJUHF7UqQxXy3KGtdDwPXa5MkyBvjOOve7/7M9h
5GMuXhrn4gNxiEvIl/u5UTxowCmwYqPT3Vt6AoFEibi13h/pb3xF0yOiox1OeMB8
ukbUWDqV/c+TeEePLEGZsEOySAarYQX6YUfA4jC3XDTyxf06sY/oTGF3/4zWPqoZ
AY1yyJ2UTLHmnl/L/ZWcpfrLHgb6WeTyD5nSY7rI4skSz4b9U8ntmGi0RDVHiVv6
5qGiGc8VOEAwn6wFszgORbjcpt19F0hGROEj14u4fSGCiyczKo5WsAWsGGQ5cMfO
EnWuergGCj012LxvxmRlM6rAX1BdOwpQrrNaX12ami/+OONvwB0n0is0z18116fQ
b63me8qdVbQVoO1xViw74CNdnkpbm6h5xs9rrUqikZzEliujmqWmqwiqb+s3qUGR
sTIPSZIG9rzMG1mr0asXOU2c0uuROS4HmLzoKDM2kcOgCvMuyF8AdWnw5kznQIjw
IQegcPWJe4S+pcBSq89ATKiead+UL3Ng/K0OXqp6q1q5K6L0OUgULNdVj72N/mxT
cVl7+McDWyD3ArjcQyTe2Sb2srKOX/XYbL2Bi6bfHNp1X6DzwtIehZhwmXad+ILi
Um7PMHxadtU2+p7nSa5bcM2CHQGPzvsylOMCwpDzv8dyhxMb31RnTkyfVQA46Ht9
rGAxY6bK9H9Dm8ws7MQDzj2B5iYjp7W82SngAodRdL7LxdD4XsIt5sF5Sv8/zvYS
AVoFH+zx6TsQ/7xrMxiFx4/OVDaEnc2VsHlG94ZUbE+qrJNEzuMitnJLpO5nuAbH
kFaABoTMIE9LLzEVv6MVmnO1z3PfTEdC4+DaWYDp66CFUK2sjf6zWLD8kO5VP/qw
Hodz0Uq8hf/dT26fnq4nmbvkx34k3A2Z4MwVhGhlWs+IQ7EiOVk3ZfeJt6CWN/C4
qdHynJDwlTOBxdKW4bBL7DfJ/3W2HmIKzC/hsc8bFFHtEm+dn8JogNnGaow64EHE
SuzmBHbR+tOtOhdaT2XmS+fkDFCGkE3woGHqWWTOsg5nPVloLCzPA8lFKqt43yAr
UJ8WiyNV3FGnNPQbvAv+9Q+xI5SW6dYtmhBCvUaB2eyuhTR0QatQfArlZJ7yV1bs
DoqWrHbbrTWddPPiSYFgNTteN73NBXIlmMeIBxEOe34Elf8M+GnDY4ZEmzVeSYCP
VXrwAZWDDf8yf6eMgpyIjhW6YeoZ91nLghnCv32nOkcZPzufzrJkLQ+UEHnTnOJQ
jIuuBCHyMnvanzjBLjXQaeOWsfSmcVZuH3JA1TnbaGOVwyYjedXw9Fpe47DHSrhv
GeuW5zGfFVVeHMjh8lCz02mWiOnmAiP+YsoHVCvVijY6fER/HJqBvx8RW38uHend
Dqiyh7KhGSoXIj+8gzl4FjU2PTXg3Dq0260P7CZmS0zICmYiokOY6Fd07W8PuTe8
k+WidjZ0a/uEvYn/to0a6CYaycVZ0GuqNaulh9rcvtNZEINTf4C1EA/2wCX8vvPQ
D+LO+0qT2bxAVsTWi2NKnxMpwPvQiXriZLT0MiGaugSwf0dbXoApXHzvNOyIUE+b
fAyXvCf5CU1/f7GM1yBc1mMBW00hQ4DQbHJ96c1IhPUSUXMV/+WGSx9dnq1+rxT2
fx3XsFf4H05AleWhgDhUNTt8jAvizNMVL3Fvg57MyYvi3a1c+UTYc6Ld0H1P5bmR
i2c7ML57x8688qg6zBFsOtl0ZAEPxkJXkF1EibYyf/0fV417ZgBLcQW6F3zCn2LV
ruZxWrmfWJr5iFN+bB1k3vAobQx2+Abeb2v8qBVycZsZmM0gG9r2fY1WbfF4bXT+
qZGnVw9r6cOVL4wWgTRp+o3e2PUlX9psRhnNprr4UloRwMCNoa2wBzx6yCVX8nn3
65XNb3Wf3BThbEMfMv+o9VCFm1Qqb58VZzdmHylI6XoxMaxAIvkPQ1jKbRISU307
zblbHRyxRU7AQZ8uIGudLgDgkcrxrT1GEOPCOb9RfSKYl+cxf9nOGPSnc+As09gT
auoIsoRdKmV7zd/1dSHLM5DVp+GF/Yi+K7TuD4zWrVG0uj6ybtpRny1/+JCpoIrG
szYL8HWMakuaeW/E2LIAnaqq+zRM5cpzN9iNwwR/KpNCzJPV+J6K++0hPoyqT9xx
SD3b48dQYT25h3s3U39rvsWpm/bIy2RZV6ao/fQVyVpUQkoLbPmYFGjYLDFcw/dv
g+Sr/GkqYROvScez1pktQsJu5a4gKY1qhUj98rIAyAAbzbr0fb/K2YwNGngx3V11
dwA4fLBqAdynpiiYWu8DBrPnkMaiIn8hcE1aP4lvEKxXox29VXch1A/vKMISRwNQ
IDpjtwhxJ8oqBc8G8QP0fWr8FOPclsK3pVNuW8ZYJAT8hRO0D37dzopHErKXh9a0
wwGxoF13VuJPRE2aVDGk+0aCoHl35MQGJ1fU1Er/JPfVY++CIGMBip4czYEN1ION
0g/SQz2qrp5I0p0EXIL0C1fQ45dze+z8vn+0/DUKt6alWB6OHeRlc+G4cwh81SCW
n3tr7Ck+ubdEeqg3zUUaNo7kRVwP7vpG/a8M28pvnSPC/ADaCRdgi7h/jUIUuFwy
dSQvpZRn9L78IkIqlf5HlyOZH0WuVBUUmF2pfQa2UX1AOt4ltaGAIAS8BpFZ84wz
6r4bSF3g4iMSi4bjz+ItQLw+zCW9ddVPu/tyET2VubaGJOI6V5aAptdLVNd58QFj
gdZGihkmApvR1sYUZps26qGC96WSU4MhKcAq2HMbvYH1iqQlPoCXa6ID/LtgYj0y
iaf1zcxl+KFLy5zLvuLPSVQJ5D/h1GLOAxuvC694yi3thAacLopWKrIi4AWoY/fB
KMP6tFWkYhgTBUUEBnq00GP7yARzxDXqNJmXvb44JBe3VIHqar3mToekAhWiijqE
aFyykp4oJgdz4N1XWStR28xSI9XlhX1UdK5Qx+DPFJDEXBoiRP4dXc0nEFoLWLDI
SmW1kMqsnRuV4XT2qTZdkBoQ/LLN77vd9QcDgJg5rDEJaGOUZSbFREsopJh4D316
ium5KivpSRU/efGYrX+BCtctGwy5ByndGhRl3DNBxRLTxZtjqI1Mz9dHkj4k6Umv
6ehgO3eOJER/Oln+BgZ6PzECybWoafdM8+1M/a+XHuXA7veOVy3DRe0Ia20CE/2o
5W3O+8QaX3swG9KOzQUGvNJFBJCvqUs1cWthN2Gt5Z79oYE4adRj7HX9PiPfmdc1
I0hJioGdVqN1zuDCiJ5ShADQXNGbO3GF70V3+gwTBQe1MampqdCMstpEJ9sM3Psf
C3OoI0i0+WyDK4UWkKZ8SNroP2rl4z6DSJiBlWcUCHfsYX2sD1wA8nJ0qwo5LFET
SiKetcL6AhI0JreFjzkLHFedL+oi9DuTAEwCT+eOoKBvbRdezfPAaO3bItxt50Ji
+bFSPrBXcvi3/I0mkd3snGv6jQxqo9vcxHgzJt7rcRfUql7N0pKMpGfD9SwE8tgd
slq9cOqEDIzriAr8xYErVMtP81M3MoG9p69o5f0WXbXAxuBD2i9lXa8FYtQ71j9B
uKDywa+XK3ReRv13mj/3KrSeW7I94XEcZs7xoU61UAWiJ91CpPnFNI52tYUcpXzB
E6sdoL5vrBBHlqzRubr6H5vg/oZRScJnbRs8hBTcuvACfYV2RUeOBZlaXNPbuMhb
KIR+Rd4zzqSzBOrLdpI5oDguUtdnRF5hkVZoPZRLZbS4+hITy0wDHycrzwJJYuFy
353M6ZDcx0uzMBfubjvZiq/DXR8bJvB5SNtF+g5MDvDD/9thrUAj5wmxjzA6GFhm
ltIGUTrgs1VgSviyGk1Q020wJSdE0RbfzyheQYT6gfH6V/duuGrrr8GhKk0aXrw5
F9uLeRVeAsxJG70cvaGV5EYga33DDPeas1mzF9FQcEMIhl+PN24JdulK4eogRrbq
TXQve39j/MsJ5dz8ZY+UQO33IJZV1J6wIUlOCSgdOE4Ona/+DMzZFqX/2KjmUjW6
AxdRaLRdO1Mua50LdaBz+ABtDjkxsmrnSgyRL+SlTbqcKyf5Rv2AvTo60OvBzSgP
eE6gwrptZAJWQolb1heTb+XBtVw01JMHavvmpx/likK4OpVBrT6SCHUBEUfL4aW0
/UA/LpOFXlRdgg9UKmg7/TK+EhchjeVvKp5iy4U6OaZ4CZ5Iei9PAgKW6exNkgKO
lpEQBp80yvXYLcUZpk+BND0cEaBzO6H7dYrkZrb94pJYPRgPFy5v28WH6K4TOWNc
jlquGmJhWFyMdLMxNetelIFsPfoBOTrQpmhu3cdnCG13feLAM/D0QG8SZVIW+TF/
ScoUlOrMNeZjOK09kUCsU+wik7gyk9Mlq/65HFaDij7RMztP40pLZM1kEiKcvt3n
bwFF/thUoRIuNKtzwCgltLEfEWOGLsFQAZnd7dnKPqogIufHATS3h7uuZI8Sosb/
3/VYvskwSxEjAVrdc7xfQos/LQioNccOvLhvgd9ydvF8PmJRx5fUonaqzIh7Jt5+
uIm4QZcahM3ggX0DGk0eo7uYNt/EtSyy5QKyTFOWchVxJBqL91jUW9vJDt3SEy/r
x9jt0TvNzVe79OOg+Iwi+NQwLhXvIzndePr2/4BRu4Vm0PaKT+BOTWaagqhgrmH1
VZnvNdv1P4Nf39j7i19Ztl27TXljiueRVJnxl25eZGgAWV2iI82KArCUHjGwDMCM
nDD9S2174pPV0Nc/B4BIHTPxe9ARSDVMxKQR/4u9B7O797gRVR5KW5fK4xDvkNd8
cA8ff4khMtLtSxTA0a3iSslzZy4VWA3qE4XNqdati+EJj/5K3Et3uhEIqHu2BcW9
ri3i+CULyIJBuqmEWCib2gUe1IVzrMUqeTJNKtSummaHT6bwpC3S0UHkBY8FGX74
0M5gwGuDsDcy1BEIFFknUkb/JpR+BKLIv87nfgFaxlu/QtHnMP4Vezr5r9IsOAq2
QbTrWRICvHPrkeQVQZb4AQKcRijDZo6fTsiNXcjOyp+Opi/NIc99GIkF5hbgdYQy
HfgdgYXs9i8Qi47rEU15JY9CHOMVlzYKB5/DIoJQOimOu1cnp6Up7eBq9O3GYfiu
sU19PpiZohpKRy1BD6fyptUZzp2dJIP5JZCFKSyeos5dQGdrIP42jOB/1FBKktSq
lswNKwLf+fUwJRMwi16gkgEPduTVRKzohVxkO4w0mHBL6zt9Tv1Q0zpcoGcXs9+e
7bBvfe0eYG8rn9JIsR/0iph/x06FM9DVAmSyFu6gGw+BaXKiBKIdVLmqzQH+g9yO
Ck4BLTS/FWvacRQt3eSN9L7RAXeyKJO0G4SbXcPqTP1IbTKiY9NnSGTimjLIJx90
anP2LFPMbqnpKppKZFqTcwbk0jA7RqagD0J8Hl/1dxq0ohGtpFKPOsDg8EoWDmll
/xtSBxfjT+QFoedK+TFyIYNBFvC3apVUEDyuWl1Mgxk4CmtclhC6Rm6hgR0eThuO
98PjIJm8wkfelL3bvXhkjBpkBru7c/GIKN5Fha9mg+f8yVIVjtisbVc9XDhNcaUT
gvdEmFJyyF/cGeNECCHrLB3c43YDPCa5Xrw1g+lkzYinINttScZ5AAAXJbJ8skm2
Tp2Zx96e+KvPxz6gbu28KvlykIwzy2R0XyYdxWe+7pkX2f6vzlur2ZB3fFC22kIl
Wg5MI4gooeBpkT0O2yiYsYGcOs78m3g+7iHFGwElaNbEq0JKyRf4n0HV5op77Iga
hy2oL36he5UiDc4ZOdC3qdKBJFccQ1wrphmL8fuXitZxfGJitdZnd/J1lq9Zs2/P
XqONW0GcODin2fYwRb+lkFIQsRG4sbrdgQOtghWeAn1yAsqCKbacOoekBieRVCDs
mcV4SDpwMXpbnGBLBS9ilJs0qiyqbfHfnN3rHV560squdFk9Vdx0KEpkPUy+R0Jv
cDOqhYegkz+48ESyY0smvUAoqN8YcLmlfWPyeixwuYZC3X7+VVfhGM8QWGHnQwRz
qYN3Pnq/aEjJQHY7ojFe6X+Wkf9bLpfi8YLhEwt7kWUd14/ZzZd+sJuP446gf3vR
apLd6xaC99CGP71TSnzliAvIRHgNc/6ZaD1LttofwnOvngMzQNgFK2fGmRTzy2sZ
uEVYT2sWoa2KttDI5wmDzdFG6GhNeDBXli9TTBlD1sxXlWFv8k+eIGY1Zqr2szDr
e1omIHiWdCSd9ckF9Jhp0/8pYd0NqmRDFsfzFKhgP9tHy8DnJa/G7vNJHfqzUiEx
AuXGDWBvcKH8qb6R8rE0rcLOaEJxbVhaJivAfAjGJfv3BxGehpUi7BFXbDzoV3Y1
7eWQmyvwQkk9mzPpCHkMeYGJ0LzAo3jUw/Dn4lxWhnWiuRoQsOMwWGD9lQtXLI6j
m21iSs7KVn3b6vtDSVvx8ApLy1ktuk/xF/L+mjAz1iNuT4NUpbhvy7q7Wxdf5eZI
kDSVxZBILpG1l9XT+F+ds/56DR4I2VJU0kfBu09TahpTgdP1lEbViku1gdrEFbAj
Fhsva//2IZNw6PNibvcLh8fz8PODkHTm1wakHHCBiIGAlxtWGrcH0pWtccSmJ+86
YBVRLWDI5V5WkJLFj4TV/Ev0/XASoNiKwjGtNQbpGdFDBjR4mTO/nPe6SicoRIk0
BxQ2rS6IrIFYoAM2ORRgdUO4nn5VMnoJ3wvQ8YHoBQxgq2tNaRy7qWgJq+V6mUBm
6x9kL3r0WGedE1G67KSCq9jlfowtEaWl+gA/5Y5HVPwQm42WU4CyE+1wR8Vl0rLM
sOJ+MW/MNsGW5PJrBam3++d75B+WnxjAYAm9AqhumP/9RaW74JBQtGRE/igmo1pp
1qSd9t9zsnx+fDrZ888TfOd/D8Ww8mT2DKAIL3ju7WpvHVA76fE5sXaM7sywDD64
AKxdAWVCarqyEAGn2ro15CGvpBXKZ8TisMP290/ck6fPNsyJDVuN+B4deSwnNS8g
KydSi916AFIkzbZdx/74JYB3pz589geAdRyJpbVmlX8KYUxTKMUM2IA2U7UUdBQe
IscVvt30qaM4YhzWd1W58+JRmlGoQlExgzuNT7AvSI4vQ4NMOzoExpuUzUnUpxHk
J12Qyggzux5RV5BbSb70v5gSbk7uM/q2qtTaXFbCevYN2KxV2keY4nvLjUG1aDmB
iNzKRUxjhUJ1/a9Ypt5tDCDBQI5VPe+sfl4HQV06P1Me0awxGNN75g8KiF6xNILD
v5ANSHAbCeGywuMqSCNlsktX0aav1JQd43biN9wV2HCLc5imh+6VWwFY5ry1ly7s
n3fZEmPoqTyQpAE6JgfADsYTRdWIzSXRN6Q5l1BXgE3+QxEMCisiv2I7ereMTxpK
MgZ+PYo7vtd5W0hWRi/crJ74gTIqExVoFwHFcROQf2TDH+lYXZ6HFJ3muJ5EhwUv
jTvEFW306NNbPQ+WUBYFyIP+dAWZsD/pknWRDsQ2HbEWhiEqRzT8ALCP59vrGihm
ifg1mMHtxV0PN514Wyg/u7Qjw3lWOkhoUXJYAWkiUuaNdEcuJP6FaUh0oSEojDpb
a3BisF2a8aYz/7KaSDNzlQZpb3vd+nF+e9LqXfQrmveQd5p5LrKyDTgQkF5UUDUd
97CEpUHi9lRGNQ16ZG2rcnpgEX9c7A/rY0oom2nBCdb9L+PJVsygCH35s3SQjjNn
mRnE3/1DfD2mOfyklOD27x/j8IV2Zm/w4WeS2olic6k2+/uFvI/BWEcLYiib52/I
7pLqch96I8b+Lx3rUdKDCpbYqlacrgZnRiK8lNzhgu+lO6EP9y3oUpo95kb1kjNA
a9H5HvNA/nEpt7X1AR/dwQgXmOZMoDZpFC+9zrqqzHiG0CZhU1Wz+VRezGLwRW5j
OXcAslbGOm3AXTvC7QnBRlXVEmqhwXi5HSrHxJRsq+aOaB1b3UR1HQW23NYG81nU
4QFDfJjK8MxxFALY5gy1ItUhCNbpLTPgcLp3kDgDZtScGQY/ubkOuI91FKlVw0rv
nRY2l/A/JFJkDTEOBei6NRYI3wv1PygZm4rachX6x1zgI82wpAr4FyeBwryFfB9c
9xiWUx0MzqNuet+JnhHraFXtT3zwu1tyM4ej48WU0NtAIHuNFu+5NF7Wr3blZtd9
RUqc2rg6PFMu7MtqSDFxWDmlGY9RRzppIb0rCzSpJibF8UVYB2zv1OOEVk3brvUA
Tq3Dp+G00X7eRua9/yc/aqAF0aJ59C9li2m1OeOAIWLhMOSKqfWyKRqtR5+scwhq
Rh0AoYj+nnG+rS1uMKtxG7I8zthY34bpb+8npJ2yXxcv6MlbiTBw8JNMotUUoicj
0RrR6+56dBUIpRcfgTHP2P7SCWOiom4Ksm2stP0GbuU0vjZtU0URKnSKZZy32AQv
PwuSG5rmCLb2ovyM+SKdToeIcAMj+vCZCZJAzIIYfTSOqBUIZWx+CbrVmmrfJGcs
nGolBX7B8ydkMkbFxVwMjIN8JcCp5Nv4EhuYg5bZCvRqdofdGUONbZhuJCu87vnk
HJ1XpLDDUnBC5eC5NZ06eeh5eSsMVvohA0QdmTZvWmtDwHN7YoI8fP20jUUkef7m
xywK33yVXDsbn1kF2e1Q9PDKRYKFG+j7ryFKuRnKi9RbPOAjssy8+27+j8X13NY5
Dq7UBSHsa0UogN5n8fJgyVAqHuSrGPEijqRbKuYlBbmINVVBDRsUA7bBAKJtpK2Y
JFo5hQuEGfnHNPnU+ByW51OTCjIbISfuZY7QOpUTFS6TfXz2PoYDAZOmLGso7PXB
pxX7B8reDSTj85nfooHsr9K0v5raX/8WD76ERlwTlR7msxCivM1/bYNI01YV3gec
ClgGD1hieOJFmBYSMvR4lyYbmzt9e5eqjaRj1lG7Ij93YQuf0rnm76n5yub/5ZAn
eR9kec5FIX6FTnUECT9AMU3YMjsL1phzN7Jykc9Jv2Gs62bBOirxrZY3ckp5C3uZ
kXtfD0xcXWxjzVD2y9TYdhLprszMS34RB9KhAbks3SMqwrb67/oCeqitMSjDXRAo
0CudpK3N6JJifk9ge+kE8pRmmjGrHQVwOTWiHo0ixzpjjUZaurZgvfXiij6VQOFe
aPbLXEKLdLprT2mbDhc9zFRQT4OYHj1Hc/DWWO2KQlPsROwqjyxQs3hXNrf2/419
E9zjd2MkBYAiN7+H/pbZna02Ijgl9LUclZn8gN3WC/UKK/16awzu2M8rhmAlogew
TGIQ8WQ1TqP8TB+TAvj3C1CUcDPOBPNLBrCfGZSbSul4vTryGGUmKTCRR2xUxwFo
Gey4vptjaaK/tf5ITPHSDAe0lYkgdVtDSU+nz8Jqns5BSd9NZVbetQXK/i8BkXcy
hgrywoPX7VaCNZNesSXdW3/UbusoyqTtW7pGcxzCOLUmACvotEeBWPZT5mbFIERx
HVZddUZnBLO2Sa+rcBTzRaWZ3VFVB8uYB1mT3BGZ+y0vBg2HNPsw7MSmG0fn26oN
tZ7T+jTkwfmhka31UaDxDoGJ0PGvSwHM9YT6Jjkroa8v2q5FW127xc8tj4Hzdq96
VHXXpxoR6/MbY3IQqQvA98eXsJi4A8lR7FFcMImaDLaqnEktmWdTuKRkDKLYzS6/
5hHTjxBSSbv3k/yqV3E/huC6HNsstDvrh6THhIAqzsoNHUewrWTJR8sBszpo9pGw
jAq+DPshkd5YUfgor5LSgJVSursHtVAyO0W4Ui7nWJ5d3PdMFUszl7aBGyv/clfe
ZH8vafNtkjv6nq8rZrjCfoSMMrL3VFxwdsGdCbOug58AH+DE2Llbk42ifolKjGfD
PHqrKzdTd8mvyMRvznAPqGUe40IBrvSi2L2oyE5RAKPKNP+NZwCZCRV1yL6IP04m
7SLayxJ+3Qj3pbGwoeAMwC/ZwTDpZUt7DXK6DDIFXn1MWBG3qn1/fsPRbnT1Z2kA
rO11LGcCuGyaOJz48FIv55T7Hy5nch7eP865BBQ7n4NLfY28F8J08b9b0aQCGKdz
qjKOuyE6mEyRZTOAtWdhKyO1AFVfXt06EMP4+NYdOxgw+0Ne5O21thxU6RqNYPAd
Oxv3QKJgPUv6x0xWyT2hZ5oLmu0Mf25MNQDPbxEJoEHAYNHZv9pB/O8TnKmH2FkD
FrOxhqy5htimZXiO4QAzdlYkt4z5SmA0m69F4l09InNCZcqrCvUjenxDfNrkKwgR
tSoXWGYjEMtGGceeXItHocvXjtHDwBZY9PRmQGLohLQQCpO8XB0HpF/Wtf2l/vCp
lEBErb0l55A2ZrwcTef45anncAezt4BhFjnokx7mw+2NUEnbPp6Eksv6GhQ9UF8K
Nx/k90Nrp9J2VUESrAfq8cdFYhnUGrZfezL5ZKCKEUIvX2mEHvSbL5F0zTFH++IS
5gBTzAeFjoe2ANhGWbmJkTiqK1hKxeXa1DhyW0OR/jvCmndUKbdwZSbb9IswdUIr
d+LUtvWx3tK2/UwcoBrAZNZkDMxdwtpLQHr3sleNSWLN4v43w2SkMYeLxQfFPhkf
`protect end_protected