`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7824 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/Qj5HR5BeHpcN46a4J6Nr23waMN/8tpERdkBop5h73Fg
Lp5pL6FR5EO1michUKN79Q63D2N+Mh3rYKu6aaX0IktdJVz6U2ycLP2E9+YvJvPa
NX6Z546bB8yeSfW8xPtGCAmupuXg2jKpRgoEaAxVD6jr4FVsZRxPWoLLG1okZq8T
sKakOGKTLrWaXpLU46MRPzuR8AWel/WefjsND5/hFdoIICIMmJOQXWXhxDjBmYyu
mBp722BbN/tOujUbDACvFpzQWTyFNAZFuT/ehgADBE2pS5ChhTFhF0izFF6QPIBE
JYCnueBA9CEED6d0znb0ygyOUQetCoYM7Pirzx07XRcgswB6i3HOvqS2qwtAXQ2S
9k8HrXC45Y4erUdb41aTlkO8NjkqrZz6hiBXU+fm8mA9iIdZaxhsxIRrZyYkXnm4
5rgYIUltJiry92+EECrjY/wWudW4saKHIWHk4M/K98FkBIsx1I7KbgSX2jEDm/SS
4zvG+G8ahcInWFiFOTrXZfs/mmFGu/iYHrguVfST61tifzBpvJlPu84afB1zsSY7
UhaEKAQ7uDDMmNxz0G6X1+QaRUjDDlFQQXDHRD3RWViNcN95QjmWP+Vj6k/iWnKQ
BFTe/5ir5khTkU5AFoMxHprTv1121rdeDpZbBBOVHYFblZ5eJJio9zDOJnZjApAZ
qlOF5wquNnigEX+s/rjIsCVH6BxYaxFhd5RVWgFbdLEjhLfyDigY/W1UOC+9i6BA
JffdGG2FzxoFcpQyEoItBhNYaXsbmoOeIE4s64m//Af1QttuBwL4RjaYOStEIwF7
TgN+Z0bUPt5AgEOZ2x02FKTNmsEEQwPKy2IQ0c1jElb9eeWb/R3OZBZ1i2skHFYU
NNwhUi5SRntQ34EFUrNr8rjW3WYWgnDZg4ce19lOif2bmNfPq1n5VJDl9FWMnefA
dgHSEA1H5rklfFlUeAu8w+5ZBfqFX8pBCzMyyJIuTbPUOT4GBhqi9SgketSO9NBe
TWL0rJYkN9pHXKwCKm5NHNpjnyB7v0LqZr3BOAmARYLoh/O6Dk+J+bdJ5j5efgQ1
/t1Snfry1CGA8wtTXRXsS/4E9srmRQOBxscaM94wKSB3ZJZzLObwKyVG2ex3Gb86
N9GwCBEzbW+FD7W8EUrc7HWKJvpof9whqIf4Xw2EPFmbgFewtt0NzATvQdEmtTTj
cb9NK21NNE4IHkVZ4acFTp9BU1ZzMoN5df6yXnKWQ6h0QJ+JyGeQ6wpV+BKAwMKq
REgi99xH6scKmPELeDIe/ByDj2zZrEQknuzMFDDidH8DtXJWIIXntONp+GCpQ0pa
7ls5PfEBh7E0V8+I+TI5kuEerexoP/5W4LxZ+h845zNURzT52kAcpA6xBV+XLFMo
ScJzDjsTZyH/Haecv9te0kGSd8h3N1iNS/murxx3FcWdpNysfapYFrdNHnSWoxJh
hjHL1GntSqaS0zHzbjuKLxY3eamV5rP8tzR/yBj1zdbhYICw9/fLFQyqDF040NC9
9BTLr32ocrPPr/2JcrUIvjIkd5xzYb9qwFAHKUTORErbagPzE/dReQRUUYUHPYWF
wxIZbTRaf8jIKnAh8rbabvqB1PiVFgcGbxP9wxzyQSv91EIijcoaHaXkyWziHqDb
eMVxg7C//DU7MGjcPURmhBm55bbeQtvhrHPoTcXp8HquoQrd0IXvSnsjMwxhCrKF
86YZCaXgVufxaQiK+p7k6DP9ROhbsXahgoY4ECMDHlAdBH/XSOTPs4msqJzY6BzK
sUUahztnFI6KoBlT+JpKtkieDSrIsGRHqo2DB8Y/0ZC+z424xdmD6UMl/sStfIQu
SNC13P4bGm1K5Xd5RSuI6SNFL75YbZg8ccEH4HKWkgPfVeAO4ASQ/85nEE1uuRJ8
gU7GQSojGBr3b9ep5drj+cvk9PYdGdVBUoG3Zexz2Q4gxiIY3KfedEPOpB3i5eEw
d+ymGn6nIYgUpaIkz2zNWLn+IfXJdo7QttAVcK2tKx4ykGAUjx93vjtKi6rM0P79
yL/Ts6nn4sgPOhCUnLggFfWvsHjHFAAA1tvyGal8EpLcUE0GoaqLK/u3MhNZ+GVr
7v2S/8ZT0gVwLOoYC3aFYHHE6nhqg/DriqKk1NOvaRQ0RpPU/v9jI6Y77aXq06P9
DOxCwsTShfXliFE4l721SqNV5j4+RdAcJLUMBKzGuvApe9ezFTjP1qxI8R70fDvu
XcdvnremWMRgiFMlVMfMj1NFjEHx7yOsz3RABx6PmwPhJMB6BbABw+0ar7Lnkvij
w5ileV7b2iaMlMR7WBZEL+uu6ZXc8JFGUDwR76H7iFsddHmD9oj3jvoVGJqBFRBD
X5kXBXv/VCmS0Gl6jpKCL+fX2m/QShN3dl8XBmKmrjdL5iCcL1grTNDxev+YAfQF
KG7ZV24ijZszOtyew0tCIyvPjNzei5RIUIbbBjf2lu4XQoIOitJSY+oNb47Plbs6
refBpZEF/fnqitaRl5nan9lukY7KyTQeB2t4nwjRSPr3jqCNDbaSHAYPU5m0/NtV
KfVHJ5dMnNBc4vCibvbtNs6zIFLngRFHdcsThQAZ0ZOBXWLruHLifp21v9JF08Jj
T9CC4LSOHF+uah/VZnq8ZXVuIPYTVTYgr+7RKrO4znBdmdeKk3CA+hPd3WzfT6Li
E+kbOXMZqUJdrIaRxCpKLcdIFIVmE7ox+pGhpNPE3mGkuY6tpg/Bi+XW9axUKDgj
yQP+8lXKjCCX7fdTGImW9Eb6/pa2PhsHw7vhyqYwRKk7aY+x2JSo3XHTbTqjN0zI
ESy6ZYFIuojfQ7QRKWUaeckJc4CSgWVuX5GNaojByke9YZINEJg0Et7y+uHiKHlT
KQVXzY9X6xJVOXu761jYLBIqD3lwIXTz3M2sl8waCAcCyEiMLuHkotqXyymhNPda
DQXot3oKpgEEDjRKmGJBR0u+C2I8hzB3rnNki8iyOVqdXF5As4m5yji1M4TiRJfZ
4/ezDLM4oUzYasFMVXUSs4J78JX0xLbY/zkwce4RyNvxFDUPVVwtRLM+EdGQEvfp
HN71l+RwKuGb87Gg4DSkFSu3D/uQ6A9QqrFT/U367qtyg5Tsro9eGtalGlj31Kac
d0Koh0dXm+5OLJlRMM55VsRIyiX31dK7PrAjRRKJaj2kAWCA9G2RLnjAzEqj1lOU
juNvSFnDj1+QsARNYTRLVTwLO+qi1jT1MDXdaxsyw2l2Op6KStwdzVLwpmNtIiNs
2IVwY6oL3qANjIWkwjz7sxcTuF6V+vU6eXwlTjRDY2zgwjPholvgmKGExIiM4Knp
p9q3fFxwmNR35+8Es8OpAJUtuA9GLVdNQ3Yn7dGGAJD9kDBW/MXF8D4TzmtEs42O
b2WwZriJG7z4TY5fCVZ49ZemSslsDBOS2kx0+50nJsMfr5MT+ZbKdJTZc8lu5E1C
QqiEAdxt9MqV8j2kmpfOQpl5av3ASl6Fd/TpK01ZJwb+13SRRU4egVYW+eHnn7MW
ghYtxMOCEhW/vngFZpDWgU/DhT9A66DI2njbmKgZUP1BbG4EvNzPMXQtfq6dVR7a
OPkMxm8qrTHqDyKoB2EPOjsfW7fAgdssTIVgxMyjnQYg/5/AX1Bvul8cZtqeqy1T
CYBrcb3FU/vNLTPeQVuxE5RjhrUZ4ayupW/uOG4h9bgZj9SHko2xfu8rjdS7NPVh
wmRr3AUAQGQlq13HVjj9z5mktlSeNHg+AJgL0nBB5NizCAdOXpqCzFhf54ejX92Q
zpQAVI8xmAHieBJhbpVUTP3JdsQcCcBBIx4NzH/FFaorKvDnxZHm/FGZ84KvURJo
KReRwsd7D1UdI0kzNqM5Az+nWiaNDnFO2y1hx6Iu1DFlTOlCZJ5jExaavOzfV5Cm
j/Sj+bSJcKvCQmUwBRNohqREZeSo2dI/fDriuD9OZPSOpGq6vGBXyqY4xnurOnlw
6ZpQ+DBRmLwVFx7fmhcWzRsqYXEzTzl1P7RgEPsasFk7ZFGf6GuTesLErMPtCmnF
qkvb/M/4qi/WzdrEpoNJjGiTyHc7D2uJrPf5/K+a4McZpujJxdqFVRGnslkV40qw
jVpB5tx5lLzyKgqxyd21SAavq7WyfaHOyYrvBZdIzZp98L9V8gF6mBoyIgcfp+jZ
IMEpBKftVt67CVtRmG9esxIYjtl5bizhts7wvUf1EJdL/LtvaSlYE6ilITfF8wLx
JDzL6PM5cvpoox/pXLhSFqmvo5dHn7yb5AhVr9pLA0nhLUjepcGf9umP1gjP4NMs
jeYFsFeIhM0e72EgCt8THT7BA3/h1Vd11CZRtUNbRzsI/vUFDIi6sSzFEVKOPNCL
+rv5eeoSIgIQETH2u0e4n6ayn2s1yZKgC8Hqm3O9hK1JSEu/Fd+fKKj8vuGlFnkT
LZQtsACq5omu5XXOSnIP56rVEjHILGfEjw72n5rFCILWS75JxJf0vXD5+1q1iswF
xWCCjxw1NJoYxhT2NmplXJlNK0yt/SwXuSGk4NeoaxJjJ1sWD08a7GWpm3kB/p/E
iIXYXwX1dTrXlNcgJ5I32EefjLlqTH6aAgcYAFAeLEM9uELHXs2fEQ0jPtwVaI/H
ydKeaevLwoG2MgKywikvHUMq1vUuT5dDWIIkag8oZnEqzgOu/o18kX0YLUQiGoLG
awmE30zJIKIu/KwSkVNhnia5l9WRSmznx+5DWezzdsFocEWIgkpm4L4w1EgcpC7C
WtSlYBTNNdQM4p1nYhQfMb4biCP0+/0loe59IASvlqggbHzQcLodwhpcRNbtBzoI
gD/WXg8pAi3sHt4UEz3pPaOQ8c1eRk8FQYWVU9fxPvkAO342UTAwPAU5rGnrFp/K
YHkdD5/Xoko6449nw9rUxAX0TocONnk63xWaisOA7b08ABmeILf8LQA2wtTrZ6Cy
K4jWxdHwuXPEZREI8Yv2nYRYHkqSGTO1VkK8WKqaq4rqLgmWh0+cR3Dcjf+Jmvoe
g7CwvEySxyYqreP6E28ppkVc3BQq6ytg5lUyAJo6hq3dHvTms+GZDDvGZQsfMyqq
CTNbt+Q34mn4WbKE7KAxiO0dpl4ILPxxSESwCW+QIfdSl67YppYhsFbmV/zgpt+x
zrtP0Tuy+Jxb/isSXyP8+cuanuydMZvDImI4vd89m/l8/yudV4bSkspF987BGict
/jAoij2TNAk8XpFzUYbWvjhpBqtM8Iqlairr7PGsBYZKuJOVPaq7lk1WC6DJJLCo
YeNtedSUNFdNqqyhrXuDAN3vppQEtbOXC4DIIvwJrL5Lk+k1FeVawLEu7tS7ukUa
GaqrJkIIzOd8chgaLoS5xrOqJ2jabd0p4Jp0CRtY5hRY2LxUnwFxb/UMuyaFUoVT
Dn73THsGNn1PSUUNdhK7bd9SlOqxLkkS+e7x4Z+Y9MLRC1ZG6Eo6GCTWFU7uIgHq
XwHs5tF57kri/+yJPbVdR9UKLAQ5SIuFgquzU4JqQdpQ8Jk3dPl3blRkVZf3s8Zh
mFIJc7oW1qV6JgZi1BNcimpgg0ZShgvx/M2dz4sUhVat7UDwBWSp5AlvlIaY91gM
4O89jpY75jl8bwCsXOiMr6ACMOhfA1UFa6jTmYWcwQUgL4XNbzbmLhyTqmHFbffl
KrG8UDb7MUDlUA6BmoYQb54MYJjUj0buVTY6OeL+Pfmni0RKJXMgoMjoi+JthWnU
rSaDzLNs0/hqjghVK5ccIhGIaKNO8yjE/u+jM2TsQmwCCMPdOZrg/dXA+QXFgnfl
UMrGCcn/9755u1/W7VbGPAWE4nApuyrcsbkvFSEhaB1ULFEZYWvSVroJJFaEl/7P
i+OhStomqVmt6VC7WRmVvwV+iVzSljp5hK1Ni37OVf7mSa+X82oSGBOAWo3+BEFM
I45PuQwL8nL5OsBN4CviC9h1vck8RSgx5C8uMLILdL3PV14YDLXxcKMuFnM6C3P0
z1Gy5pymT3MZGIJc0LnUg7RUGrW4iYUtoKfceWKfm36mjdAX4VlEUWQcqV2J4Gof
XDf8CvaJVmJX+ytF/z7cW9yl1LXu1q2cOntl5O+or2tUCpj40PlByXczFUb2g0wP
fXfUo0m6mKfxfxlRBUqvFjjWUrob91fWLjt/C0HWXzfYLieHceEIkDLy3Q7gj1Jy
FrWbHlJNFkYFh2nKW9fN2/9OB2O45tZ3/0cLlvWJ2gd5F8mxTahwRuCl6FtNWI15
1936UA5g5aCCY7+g1zmpoa+peQbhxKOlQnZ2MqNvuuKwX/aTtJilrZIP638k3MXs
rEUkwaiJhxSFBHY/mR3i7JVcWbql8Qm2f7IMRKZ4XMkiazDPwVR3RRcr0p7Kn0Fk
OkfGhSrE8mesJVhaq7ViffYD1y/Bu5X49lbQqBM3TcaEFS9LdxStrd6Gyq+1Ow7o
nV2FAAbZ3RQBgaKLyFMr0F8F3GccTgEq/WNIm3Oif0+dwMSxty8Nt3BjpTDYwRsE
gKL9N+u6NxK/tjJpEkVXR5Z6ptG3WHupoLMUf5avN0c0zAcX2iEu+iCuF2/qM3CP
Nbgnt1RoMOpILCLpvFTvwFu5FDskRz0uNQAL8dDwCmkriXLDiF7/xjNT772Qao4/
LmJzokqA7C8lnyy5KuNIC3dNFgtJHL4Gj+Y3bjoofvw1M4aBl32Cs0lzifKeyYgp
PBafNbRZIyrFpuKpf0TMSOioSAt2MBKBjGjmMF7Qqaw0WWq9tWJSmkuxyBcTn/hi
hbWFQzFkLWdNhoHtts0kNUrsEip5L2F4tFy7k015jXQgyHf3mx5BojObjn6RiuZl
rJbQts/5TAzqRKSIleMbs6X2p1LCvgh9WHzW9xIl3ya4s3Z9ExZs30qgmAOg3TX2
IkwN8xTXaNzmNz0s/o/0Uk5OB1J6jga0ocj7OrlF8LqYQ3HQo7nNuB5/cRb+Wyop
I9A3M0bYhrTl1Ao5cYEvwd0Ho4E0WrxGVq5z3aioEFxdMCEcbFYx9UEBXHTZPK43
GGcVB2969u5t6Ywd1Sk1tPqmF2e31dPKgrMLMAhG/5sXl3+jHGAv1NSPHMYoHR2R
XuIdNZ53ZF45QSeGTTJ9HBYU/TE2XhzynW28u2LUxwIqER0Kehbup2dvpXaHcFBt
/Pj6Y2SmDIZE8cHzpSVWp3oP7UZNgw5i/06FS2A1vxB45wfl9IWkxn8mOh1wUiMm
djJtpkL4bm6bsaTKIrEyIMOhF3NyQLkS8APGCBo9scGzEJ8LR7ishV/5gorMO6HS
E5+8SX8jai4NKaYVC/mutJffPuULQ8dgyxQodjWdfj0K5GAXIZoLQ+zd/roh4AfH
2yNkDY4TeZeWhg5cscTOHCnD0Pbvg5r4BWPpLh0pl/rfmhFjr9fuyjgaZWb81li0
X8P/bSSUJRpxH8LknZANJIFIjVgkMTfoc2Sdghi9f5CsYewvsabx2mijem+fMA7V
UuCBipWqs69EX/fmANA4qbBG9PaUNG22FUwdP1hEkBTX8wphv+nmu22+iN7iHrut
sgbTcKdIvt1wNZrkHfFg/9hx++i6Hdi2mwTUpPS19asGOHKOWEFumJKxx/f4VC1i
AOs2fT1iGEjKvMXe9L9+YN7hHC64wdxPyH0v2uzDbRu+hqf0jqc9haBzgqf5fQcU
Rtw8ikzJn4RPzRBTIWpXlGAnh7OSInCutSyQeBEtMrQ/L9S4hjPuS1ZpeOU6vj5U
+aV5OatLxM+j0fJbND3fYTgjitBmEc+LnxOJ1LhGaygp49bXdp3gW5BsQaTIXGWp
XLoHWuqyZHjkFYDjGEx+OLV7rwA8crBvjSKhDCE/NIEkMGY0c0FdGP+AmgQRfJh4
46dLTp75UEnL8yT0v00Sfv0bVRGsGA1H5PSX7nlifuERWpKoYOBx0oVbPrb8UqGQ
KaC3uFA3Bu99IRKcLL3CJvacnjtncVCHlxlL87ZVfh/t0DGIYqmtUcbDW5rE+oCB
WIHrqUWppxdZgo2yqhJrx+i9kit9CgSt0jww/sZVHtL/VOXBCBABYvSwpFO4GFIC
TucA/DkN9q4IChle7D/5nzf+ASWUqh18PMJKVkhpY1WwuWla9jA4fEPnf/HEwlgo
nTFuljPJVbWAIbBQcCy081lecsAFyVEG2ucTjsNjNcsLbTAUcYKhhbwcIE3mHZEg
U5CXOgUVu+4JlvUrIlUKSuvlFs18WlSEoK+AomHsBF5EoG6kz2EbLIJGtTIvR6UF
CiZ+jNhU3/QQcLGUEXF0HBeQQmHba8Gc8lLRpCArofWeltJeep7i70UwI5Dbr068
NpkfQLAG4goHztaor2IEpZ4TWqNqjT+uRSWahFLXXEi3Dv4Qqa3xTKEpULyKQyiy
KWRaB304vNr9HmjekLmcpexje7FyWFH62RQcDYAQBjjEfAWumHmA7Z08jtHytxvQ
ALG1Zj7SsnbG2Le05Yk2/j/JUh3QjSmNFoQbOVOW3lD6FH1uTHhphPXm8YqdaBVH
9KGVb8g13zBSwHWZ9QOyOsJOvsV+SIt08mzbUos4L4Gh5I+hoDVCGhKLIVa2x8pu
J4go4vE4RhiqrJzJc+3D9e8kV3xcI003Y/tBifEEIhHzRM4wQzm/uFMHfs5C9p2U
Y2xR2VGam/4d3kSLHNGh6MXjNAsYa4Tpwpgq6QWHCuzMTfc1mX/4WzcThxK0wgTm
MlKANrxaOu1w+h4MXxHcz+z0fcrGthAnGqnhoaT3Lu/V6CpDUHP/If+fNfJQMgya
x9vJjZT9+ZeIq+/83LyDcmRe5twXRjMf1h/SJDJlr/cqAm899bD7Dyh7yccvuG2T
k6cnF90whCCCMHtudqzH1Xv0o7IE3c+gmT8512iRIXupLkHfDKjPVab5LkS9EsuP
6k+3JtKNXGAWaXEiYpEyAmY5oP2SB+i6HFRHkTfLFH6x1sXK14LldRKEJYfOrIqz
lUZazD7AO+hwH0ze9/TBEQ74v93vRzf/khXn5tclCnzS77A205LC0UJRY1FP0myx
8OkWpY7wUwYlKjdIjKfv7BFGXDXvVFlqXsLrMntIazyGkwcs8R72Wf/N9Rcsa/p4
aL0c+fQCLEhITa+XqKoVz5mc2oLGO6LqfF+VRKL2tM3ksenjTmjuN8UQq4wz3rpJ
5Sx3P2u4smG5rz67AAUFFPRD7VCOEx/CqGdmgFCjcgnW3F9AwskvoFpW0/IUh2Jq
QWqBx7LX4SNXdFFKSPi3kRUD6XxbwMuOja8uQ2uXBYSgb8+H/oDIGo4gW2vAUQxK
gUW9psOub4LgyWDWj2qqT/Wq5nxj7JrcA9F6tihD8uzQetWOihOE3dYg3CGr068d
DEBE1S2hlhpR0Hbm86EV5VNDF0JqNxmjxDA7AjK8pMHUAl3f4vUlMYpDHQH0ILDW
OZSZqSghS6nFLUIk/R41G0G6Tkb3cA8AlOeM4B7MefV3nqRWOxoVEPNPjXRxNX35
NC4LgumT+FNVi4RZRgn7TkOXonnzFptR8DTFVbvvzenOQsXAD6+Bw+r6JA2d2tDJ
9KQDBrfAZ/KTnHQp3K1q69ENX1XJcxbCJYHFpMvRwhyoqj20iUb5Xe0KJbqxlZGH
wQFXIzjfeHy92Me1RFlm2B6utM1KVtQj0GJ0vdU2cf4FO9uufDgYAPD19luRKWfV
FsSyg2OvfnJr6hk2MPKtJQm/1h4esafjhdtPIspCd0uWh4Hl1gHfLHxmJjtg0KP2
LZ+t/b30k3s+4Q0Ie0aglXAGK8BFzeEOGGPgtyUfMfsIwOESNLMYRU/fJIlUzDnS
sershxLOTs9WGPolroK3CsIf7w9c/uwP9UK6WwecfJTozEOr0iw1SE+sA3xkKznq
YFdgQjflFgSFvowuvrGjkuhNCHUalOint1u6PDdfuSfTritioQmcQNHXZvAGwg4E
aLHaGDLENgvFfaOy+jSFqez//qtRho0h6AbVJW3D1Vaha2jcFTsZ1AOypZzd51Ps
6fLnsph62UGvYgp/6aBBkING2+Bihd2wn5i8WFT9Vf3cWaDn/IuTegxOet2v7PUL
zyOX12CyzGh3bSS0h3HTG/1FmBvSifJHmJ9W2yOJaPXwyVj8CLuDO74qIxDQ7IsR
nNDYEgDLR1R+485ZuqWSO5hnGUoMyao6nHP9OfOf5imUh8PKWWw7ZAuVsnivWU7P
930IyUEV43Qlq5hzeUiyiqu4GI76qlbhR5Ks19xmbF6I7Le7lZrk2oZsnKn+D11v
O2cWzeV0VALtFSCXNyhMEizhQl5KLf5di0RoUQKlieIXOdQXG0x5PZEQSv+CSuJB
vOV9vq7Rhc8GEC3l/k154Xm9n8Q84+yd68a6n0AeP9FNNozALq18AD+1D3NiScl5
`protect end_protected