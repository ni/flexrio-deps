`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 26864 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10GXbr/0ybS3CmweZF54Xqu0csJkoL9LlEdwK1Q0L56ji
hDPhTsmTmqytC1wTx24RTT5gVTa0EhmGDqo27NyPYyp0TWIY6O8IgI12NOa2qcSp
ao4qTnFyjO44V9OCEBocppPJev0IF/n+XbpJAY84cpGBOvM0Rs5+dwgF587ZMTPC
dAzenVwKtz56c5XyQRVrgGfos8oxjOEbu60UZYXti6GYf2nnpsOlwEsyjcp6CQkB
uKmFODs4Tg0xGpw56QGDE4sfBOZ2fxniArb70n0unfBmjyulS3FJlCmPV5TABLIt
/STU7s/fUZPFkrPK80xWBZZESU5On2vxkka5jBwjb0LoM5BZCQNqVqRVqAUJSvjb
lftCHRM7aWkDAKwUcWdMbm1WoWHkACrvX/HBHjvabRbjylztvzBM0CiDmluZawgW
iYjSMWFB8gJhP6P2A034QqRoowFtm1gawM4K+W6AcWqHTdY7c+E7Pp7p2nxB+G7A
2Wz63ryDA+VqZNcq7q+UVagTpKvL13t02WU+yEsvRTBAeb4lMKpQ9uKl+hBIHtQU
a4L+YOmVb39QnxCVu/OCAEGVstDpU2npl7ZE7MrreE/vXlJrSh8nfR9Oo/QXbYD5
lu25l8iat1/LjD10lvOJu/yFYUe2g0A+yYkefbJYI2f/1JTPUTSxWzlH3+eHjC56
UJvHzBprRSRGckPQPMC5AGwcKc1EFhGK5/VKXyez19ldBvSXjy3JcMMiUQb+Pv/0
10SUaIOwuPrqMcllTwqNGiklLqq+C7c9MH99f1ZNUHQI57lpfZisxqWn3+WPCeJV
xT12/bNU711paIQZpdqfIC+A6YenLi4ED6eAFOXTgSgyVapOPUErCliUI5Q+aXSy
eM0ZO3p5e6nGFSk3EEGOBxBQM5PMxHONxeabvwE4vNVe/4ottRh4P1b5/oI10J6a
djqcPlTLyetVDGKD6qpUp1SItG2gILfzg4XoN1uEfbN38GS4dLDhkv3F/B4EbAM6
Z0++GwFhVox0aIky8JVlOBuhmkF69UQIy+zq0wNP7oJ+XyCyr6AOvoA3hepFaKl+
Lo8JbQY/uEdM9eW5+o3W0xGgAXy9nYWmtLMJoRafa2xS4e3o+imfIOzB0zTeOYRU
fdkBcYKXgNjN1UV64eDKOkp38nlZSeCmehxCwenCAjRIRT1NbsQiGPcb19405UKR
nslqeRoIcFgy+JYvUiExPOCKPQ4P1R5/rHymxwSGF95dHZYYPChEpW39r1IHU/Nc
tfFXyANufICuEIOApRmp+peAgqUM1DtpHAAgQ4rm0f8xqTcPp9MvP5kOSiZYtr24
mESeVVeEEWaohba+xRj8ukRExMH5/rPC+9xeg0b35upfCo+8w4U6TjV8m6wIS5JP
sNpnkG9EKzmF1c4vCIiiIJnEBmnQF0XVYJTQ5ysyB89AFa566WaFDR6Bs4I4KDxl
7Wsqnn8Oj1kNpnCdziJWji5Ad/fnCJ4np/uZbWnZ2WcgaIBbiBVTbXo+gE5YYN2D
fXSdO1YOTOhBRS9YyTd0NzGAT7txsoOTyrmNe1MoH8M6PIKNwPViGL6HP26tY3Bz
NelsMrjtGOTaOWvm5Hk2yF17pzs+Iedyez9j9EIri2kDSXuwUCgljiM5JJNp7nKg
G/Fqd2SU9DohVEBtOQDKezpB7XPOivtcPghmdD1Oo94fdgF9tIRb/7gGqoga112i
WCFUQ82nS1T6Pt/jfvw6GqlNtKtzIqYDShEFuF0Zc5j74+SBIa1GIuICPakG3D4J
Aj1zZWRQdngt6SdMsW5hzo6vwsVPxJNZhVGwSk8k4Zv8SYxQmSEuHkJXwpKWhzKO
o2sKPzXi5De3Ymtww2j9jRuR9E0cLqa9sKW2A49nN9ZLKqehZAA8sr1q/66o8pGI
kkBjrsbtDpXURjIikaF2toIP2A6mJWYjrm/FR7O5cZKwH2Djpi2fIGQO5fgq1RUN
9djUqPa8/ejY9OmHZeE2ngmFoJZVHq8CaxSC5YnkflX7q1KBmlEzzmSrbXeNir10
CwtOV9/70atrV30UhaC6JahSdTwAgIJBxp/3jB9ZWJtgQQZDFjL8K6IaTLAlYksY
JjO42oBfCf8PRIeAH6dtL/yQw47htt5hqLX/qRXLSBpcAUDWgN6mOaK/b7rQpILC
XmWIwV3sSnlXvS7QvabOlv8MYFzWjhPugOWXLdZk/aTBamtMNcfMDF9qiOhhhqH6
urCpyUSbWgouqVWk3+Lr3O8ZAEScDrasqGT+UtEHy00TW5koLcZKo4XwWktulyuF
Ae1Jyklw2HOwARXm2f/V6rv4ekE8P62EypLIFRDrR+VFiRFUBByzThfBlBPNwe7x
pG0qOcbRExGyiHo3NVBNVpfDdouGfAUs6NhP1L3JV/wlz4CIeEdbT8AstECYiqHy
2iNtuoZ+tGe+ETa/HRl6Fm1+t8vi/6FiGMWEjXUM9QSWIId8B0y86aELyFAmo9Wz
PimqOfOjipbi5QkPw/vc0L8BWT7IcbWODeEcWX5EeBvbbXnaXnOUgbjmXRW4L9AM
25bCzKVQ+wiMT1g0KiX/B/aU7Sc9hB7jEJonzmFop42o408s0qADw3AKdEUYuFcm
s464spzpNm7VYwt3S5rQzkXOiq/P6XnDlAS0St+4QOJDQBfpim3H2b8Mn6bqDiOz
EcUIq7wPeV/IuL7d2q6uC6qn2MgDgDbbVEVAiQCicpAvAMnLbV6CdGQQN3Qebuzx
KtefGdDCWTR6j+23jes9FbRTKUhERJyEcdVDim6v4vAn2assy+b0WIuF3KUCAbnK
oWfio81Z2NjRwYwRAl8tQeSGgL7Ylp4jKuw4Dv7ky/7LTnHJ0FnPTlijxD4NfeHn
RKZvkSszD4UakjdOBsBLCPKqFVEadP/Ujpd85wOZL1t0Vzoca6fhlVrB8g8g8jjb
prAhv71NqW5Zj1grhEH4dBUiyiGSs4LC0pLcmIcPZ/ocfm6BW0XhfaySGuduGMZ1
Ar8BJRsjdV0Ys6p/g+WrGacvJuQ7VQFBivlZRh1jvA3k1N7vy9g6/jrHaiurG94+
ZmN6ei+AOU3R2S5V0Ux8/ZAaFWbCQ9xkc3c1TU57OE5IjBP85cRF1M6HNBA3m0OY
eifToqAQc5dKWMMfw65KNkegxyeYaD1tZSLahDarUp654HdvXsqF+HhimMWR9Bum
QRLA54Yj2VTaES/o9LgVBp1wM3i4i0sFAv4o+tnaFaDzYC/sh7MRNErUm1k1gyut
43f2Hjhh9RxIfV9DbFuDxy1A6A9WgVlY6urJDCsdWmUj78ZoxCRSQ/0zsSu1WVqx
+JxdBtslIWKaP8k9hCu+H6SgV4GRjp9/gA/39IIwDelHZADfuBFFZk/W5TGsO39R
V1jTuMe8JC12t7v26P2YUqXurmLpLFScS4M2iaGHpz321b9b53bCqTB7K50TjAo7
hIx9ZDjnJWJninrApn7kw5RUAdKBASbwB6uv3QfD227T9tiFkLJlKuSkQEUvaN3O
/z6HLb4wElWbT0cQCKWy9EQ6PuZFNavCWS0bBaiiC43uDVAaVot5rce/gNGorD+U
RAWcMDBbWUrg/flpHu0I9zHMo7eOyQxwrTZi5vMfvpzS8YHVhAOJeyGOzcDivnjG
rLRyB0mLGBsmfKiu3SCisu+PT4Zek9PnEraivA0CnDGpO6caaesd5069oYwQ69zE
Dr6mZlThvz/peGcQmGay39/MUJdVUKueRL90fyFYNIHN5afQdJQPSUSA57TeSEiI
mJOVbFsNwWaEwrGr4iTha/w8CgiPuaXSPG3z1XQslhTI7pknpSeJbNCDUBbulAYL
hDxtUHvUGEUffGYyCnIA5TdCNEiS+7QyOxOY5jX61TrDjcx4f9bYDik8ilw09CE0
7CbzCNtqo4FCXEr9pd73npUIt2iOed7BlQC+ze4gdTjqkFW0S/nnSXxXauCSE+Z9
D/Cn89ohu75gctZWbXX3Z8dLR5egVWz4ZIipP23/jzpOmY6CxWA7pphZCmsXGOF8
06q3vL8qwzvnFxEM6iw4Wl4wybr/+lkZO8ZlUE15dkszBrsEc+6Ym9d+GYLcrrDU
g42zZ1L8a0LlTW2VcHLkQWEzoNuoWQ2OzLakso86V2bpgCZIb8g65wEdt39FcMtt
topZRRSOM+Q/X2wqQ+NV0U+L06LBTJLQyjqkpaUsnmP8GKDKkIdC1B/mI8/BELFQ
KeAy8eY3M+BhPi/Lbj/cfDISYMQpmSZd3RW6QA39vZYTfsPK2h3PIEvo5FrpRwy+
7+i2+bYiod8eHqTtGlobnUiXvMZznLREX4SUCCyiBYCzQFJY8GDzrRbFhXo86Y3q
Mz4iJTJJwMElMSjq59DvTCnBYaNPxox0HKpJSmxnX3EobbHWxYhARiyV+3F3k5TS
2FL07hp9SOY+ppZLlAHzDBuxSVo3kO4OzRNQqqWfZGLWHid7+AiBEROqCWfyjnoh
YGNokiLElFmM7ybp8cJ6kS8x154Tc2bYIRRpO9B9L+DFkfEikqhLTSu4uLIRCyvM
cJagYG9yVqulfWEYiT+oEDj9O0U390a/HMuJNDs+5QA93neIev/PP8trMFo/5g3w
z9/o+ao1HoMX48bQrweHk3fXRpjjqxepZ3oQgL957eI/p7FapIP0dd0LBDjcv2w8
hMqLKnRnHewsyxwXyxizFUyZmZppa7zbI5TPcoUPzpyXKH0Hk1E/mD/gmrAW+A8C
n884ar8rbgLlHsqe1/ofM7wffxLscZdpvOFhuUBlZF3+72Qysur7ITVZCSLg1pI2
MMgeO5Eq2I/0RZVPZRP7SPW7aTPNE5zqW+sfZ6rvjFQG1WbEkC+kusLXLSVyg+Ev
4yXMpwUsbv6md3acVkSZzLVc82PrhLd1Y2tILDovunWsxhowZ+3BpqKKKAO9t7+T
pxQ8YJXvpeIuZhBUHhFySYhqBiRbqv5SvJKK7bGKtu7XIdMIoJ/Ga8CD9QcXQ9yJ
FbybK+1CZJtLGqQvtqUoAh2qK8vtTQ+pN0szBFwsI6rH3Esb+xj/S3HdWYdyJfyU
B/URIewq9y31UT5Kduyr/BYoOzoU1uCsrPIXut4vJ6IEjhrkh+4S1hytCV1cqsHQ
J0kCcInpEIS9+DU5tniYa4QUH6iHgBqpeFyO6LIAiMoOi6sq+BDxFTrOmWVjC29t
AEsa1sprsFy3jxgpJk5CGkYPZrM1qOwLA9orxAzD33X3JJkwwAT7/Xwn7+DOOPL1
+nBG3N9ecWc6y6BuuH4N1P5JxplpCYppSTKQhWYE8V+ikcxqCyLMsE2hMysG0Uxm
VbUxqwEnQ/S57j5p1WFGnKhcrCK4jEZgW8diKfUb18b8Qyk1xXZF8kQZ4tuwxu32
7q3qB+6unutT9V+2Xj9HvuWcgbXkcwQsUVdEq0PrtQ6s7jw3N8OMc4tMPBNK4Llr
PukINV32Xg/IS900KKp081mwJRXCJGlpuEief6W2t+gxkcycPyoknjYftz4LBAhy
B7y4ehlJHGsZE9YFdiYwzqq3mpP3RmHJJg3+ioeykDuw37ZjjKVaiKY+vGBWmdGm
Rciep/1I3RfOZbuQ4sR1WOAfQ89kzvOBkdthinFhumQ8Pq3OSGe521ggE88kCe23
Jg8I0kKQB5A1T2yFKGyJyafv1MyEZgYD/zJwSMh3/yRt8jihzyGKEE/ibmCM62vv
Qz52VRyFeR8GdIRqRg3Uw3Cd115ubdy0mpQFTr3ZviRJGOc7mBnyx51iBNoECT9v
U6wsk9W7IQmc14Z+QLhtfUO4Rbv6Ap8wGmRKnnLuy9nZ5/QLkimO16+NhjIs4Kd7
5t3LgrPvi/B6mf5iHuXuuUqUOwSsP1d6DT532vkzPuNuXhxB6Bv6nlPKfRDTGues
E+U0gHad9Yu2z+Cuy29/mOy2t3n+5oq1hd3TnUjq/Eb8pZDdt+ie3v7VNqiH4Ud/
mCpXu3fadsRzH589W9SaFagp7x9UPo7S4sDqcYmW7yjZXFytFoyuV+qNYTWBqhAE
DkiSrRHDQdAP2/GkUwcErtOZS3coPoLUgu/G05YJ56DaGk8J4C6pzD2HhZLi3+q6
CiLKxiK9vu+/ofwN5MzaysYinrofzqwyBz2gXmb0aq/RgcD8nLei+sorGiygCUX7
+PC10YO54TQVjGFdtsxA2lu+15Gej4SOv4r0k23FbfMaIc5hf+Y8YV5F+J+I/4b0
mzOiELaIE/BwRntm0pyCCCj5ybqSnkuT+EAyuw5LroKzqEtO9SnLl/GeVMNqawKs
AfnKJC/DP7iCXsMIeBn1ZPdfcKO1zF/v6oZX5bE3Ur+R1rRDsbr2k2zDwfUjaAb/
1y2bT/XZbSbiTuKHwA/PaBI4IaZExASvN69LbLFyXkCfwsSRhAsdIYVz4qQIZHHl
YU9HYThWUggOJoNW5sZb+B41n75eoIj0OhZk/RuT7PRBJsjUZlEcCBS+lt/VcUlu
AM/rw8klicH901WDcV1BnnQPt+ppUyx5+mJYsh/TKr5OU6SJ/3e1ExzIGJxM9GZJ
BXucNQ/gvBLEJLz3at4Y+nFZA9AobxpjI9yWRIjPkGw5mJj0CF03NKrTbJ/DMKx8
MQfWli6wEgoN1FYhbgjTJwH+7V836XPI2aECnVlKjc4OUTOYeu6m/FJ+H7y9NLBN
YEcV9j487ohlVikF/eRMLDFiTX4FUYyvOX7YdbMqMZpSTBLawH8pz5xeOqQkqBy7
pAPCV2YuZdZfINq9Hy2kKjVrVBGfe8+4HdO6gyrVCAoHyKZaT1QpnrGBaGv8HTBG
6sUBMW/VGozw6dHyod1oRXS4RvHmuYnujWPM0GXbiIX7IIn6CuCBx4DO88+eH/Ax
On3H2pmtqvs1fkjWL4I+EMgmZnZ/C7X5BcQ4F4y/AvdHOEhW0g5E9aWqKjaO+eDu
JsfU137tOqKuc0HMaagBoQOpaE6t2mwyvjcre16bCGtldXGcWoaJ6Ywcu0iACpzO
AzCCGNRbSpXZkHFV9sbBY7VYvPr6xW0e/oQUdAtfdikoU8YkkLdUTPttzmwcw8zF
l2PruWjOYQmowxKGvshzS8h9OoZwzq6poqJMi4PJs7c4dfrWRzFyWMTfrtWWm4+l
PUv6W6WrZJI0t/qi+W0V2tvRJGBnM2RhUFgJNpKKxOf2PnVPTRyFACZMiYoU/i+i
nSEd3wKGc0rDOP+ZlWEjB+mDMeO2Z61IMkwFvtvtwDj24VQ3RQhrL7gztipFyv09
KjIfKKGVPW4npbdS3tpIiUKAMi6HFXf1qO8+Dc2HJjY8BC8qSb0/+KIGLBMce3eZ
02rVd/pm7KbpvgWGNcR2JVlcPm3yLl3uZYiUhbIcInuxPGkqDpRV/aSUNSxz7U0t
ng02H0ka6gHHDuttp6wdRH4myjwOjku3z2mWmI2KihAnNTlgY2tmj911cNs6ow3X
y+1U8O4snxFFdPv+5PZymkzm44/ykQcClMmSz/LFb6+N+OpMnJ+qAfVypB2I8Hvr
DN8Xy2Oyjt8S+Bn/fObkBJnoyHK+L8+O2vNrztB8DN9B94r0DFvQIpm1GTvG0QNX
gzK4mewO3w24Lr3ombbJWBMOD0r6ylprtt9YGXoS7v7sL02qselwolozRgOHeKzW
f3+b5nkjrvRYR2XxIGWNS5BlRTpgeEcbPBmF2+VJ8T0z9B+gfEoNa5VTMkIiiDvz
tTb+sKQm+G/SLuFts6Uei9JUOgPeKbqxk/r7RkaTQ+yDz03yp37S6rWtTFVs99g/
qP7YHfHZt1h4NqrRLFOe+oDHOUnIhFiRjDJOaQtiuUjgpq+NXvyoVsuYz0Icb1pt
XrjLXOsXe4ZZTXkHdwQhhj5PyF5FR4p+ra+7QwnmIHcubys/FGgTR1dlrICs2C2h
6iwszP4LEz4fp31+2F3kKFiUNAA7950pYq57RX9CuyPznUgf/zn32ja71na4+hhR
L4So4g6YSqKfWk/jT2Khh7ukOgsecQf/AAmQzrXDUscdKz7jEqVNP5XcJaDjjvQB
Fw6xbyFStkkJohZPfZRw580BnAMdJ7oeFNJf3AshILHGvnsTRvVv9T7CHeRvKAlb
SqqYczQ4Ce+lps8Xg5aSf/cHvh8llewW5v7GwxYKFZJxPpzjBKCfW7rEHgeDlguc
pusF0miGqSqkD0F3krL6bZK5aq1+TOtG2iopezKSwrgwqu60mY9c1KnZBtplUWuH
1sTMKmBO2Z8+poU+V9kFHFJ0HSFKsRYyUFB6m6r7TERC57jvti0PxcIg4oFFD/8B
l2J1o5IDCfFiPwsv2KCrksIzr2lzhZpKeAlFWsYI8Lmz3+R/rF/6dUr9qwaq3Gxg
R6yxhkXqToxEM87NCn0Dh8XeA7QhEZmi3k/LG+3IdZPgi2I+us+psRg7f7eNnyJb
fvrzOfjT/LnGvUeupNSE2IS3cGqRNvpFobZVYQf69shMA1909oOfCq4C0jm8me/O
n5PnhuZzwn+8GU+Bl72ubfxU8VMTwZv0ogG83acQAkOt264rmiSp3/gXwUYjHQry
5y7dT6H+s7xjRJENe2WNRU1eWvq4uNcutxYZeytMBwMQYo74cHDLCPiXNNgD7ApR
mq4mYGWSmcETdj0Qe+Zmf2ZD1FESFS7kq8ycdQjWdSKMnEp/X9I5DSkv+oaywJwn
uy1wpFwsvvRYDmu8vwj1xSUsVyLa4vZgQltk9oqlxv1w2Y8xOE3pDxwgDZG8Ng37
0d6a0uNNq62TE/fz1pi8aPNkdd1hEoPnftl34TVR2ku4mcyxlalBHGzjcB4ijkVW
ueMppnFBYjeF/klBRSndd1wVAuvU9YVc1IRnrYedxtqwPBdI4M12VP2/pUj4/tIo
5Xtu66BWPP7emj/t4Bf0epU//fhs6mB0A174Lcl0HUCDvdfkWHewhTW5ZqXywsrP
+1K7zgeomTtItDAkzJ9C2SH3RU4jDu8s4Xhh/phZ+xd9LSPNKFEKFi0y8YncRFa0
DYTrtRAORuK8JJQ1ULpQI+TNzDY0FvXL2vKnhq8obb9r13jeGAyOgL7dpzMwZvzI
p227B4afZqAG6NfoX/6zMLXnVxRxzkyXEeR78UWSl8GXZE82ghVQREOF/0JUoc08
T/1BNtA+joFMWLxCP1GxSQEDDT6+FQ5qkm4N9bxxeUazNg6sRbyiXDHPpdvhmVVQ
FNrARQN7wU4DzdCtePWXCOVBJ9u05uhYrNbWDJ11kso/E0vFc943FUT1khk6+gXk
39t1Dj5b+M4k8+UtYdf+/TI1XxnEEZf67IaO8j1nCtC6FIe7YWBvrpTwFM9pj2zz
AIZu+ECVDuM/U2Eej6hgG7xd7U0W/dZ1cjAozJI09poMSAXLjc1IsYkfydrFAIEO
ttgBnnuOUzMauHFlILMx7hjO08dpmngVI7ryZbE9uaRth0Ajv/KcjBPcL62ksDGr
4EAUbmKtADx4CWZsDmN8OA/uLs/O7TsZ3D1ZSqAtAeSpA9FFd1JZyaU3F8pe6/Fm
pv8p+gEjmRxoFhSUkZ1BCtPaU4vMWsgFv+XK1I4zWISQJ/17UemxXaPGgekx1aOu
C5qsUyFHFZ2rHsY22ozpJN0AUp7FYrCyMGfYsvg4CClXzu05MVaZabwPG/Pxauqv
OX/kusZ/Hdu3zP6p+TEQZf5MMizpy4TRDiTERQ7aUxSWNYTgzk62eK38EXnOxGbX
M0/RHega5tcDfwPnVF65JzWsOId2fFj1TpuOHc0yQ9WjFTEzXcRGlovM/CIBiVfz
Ucg2LvXwlre2aueq93zMqsgktiima4vWYusCwidFJtnrENJgLozJ8GNvzdxJuAYS
OWN/yzHfQI3U+1V8Zxduh2P5Jju/ZqzR+uiGEVNve/EsmLmMTyg7GpUIKbNHXBMw
BR0xErrFlYs8/bTQWr02WoWx6Lv0hLsuE7Tp5zWppp0KYP7Ba/T2fk5KD7FEQqSM
WottBGFWsMjYuFsMaSZsD6WChMSPSa5I9pIcT6VFS2JbzF8Bw0KMAci3sX7VT3AX
aojhB5QvtehExHd6TWvbiiY7kYuczpnqh9Eu0INXkOqmmcoNo1UfErYTcSCNWYoY
jl97u12o4VZW9rQVOiApUSO/56ImFQEbJSke/iQchXvHfmLBU0WF2OXVPhk1ilNM
2RRgaZxN5xDzrZsjSV0YtjMiuLsrDjBSBIc1aQLgyeffAFQqcQ2VYNJqFC7cZTB5
kGIrHNyWIABsMSlzkHlkjyNaRhje3rp2z1IGufHiAsWhm0UIfwTBJrkeVG9wTU2o
re0asiFUEdSDO58bTZ1+Wyo3O/C1P33rSMrQsol7kjFWJtb+dcmiRWrthxIsWW6r
irCibSv/cjWogFdhZOJ60/XHiYJKGxxmB5+BRVsTniVT54iQ0oGC9dd/9ZWh2qsN
0OYIXLrfdZAXk08A7xDAG+i6gbTpqBeopmt7vaA0x1i0amIXJfJFyOdtkrrYLryI
bShBKaoD1/VdX+vktWWnKiW5AjlQFcGn3uUn5bCgZA7bO6IMB8FzyNRH293I1AIT
M30YR+DhtsL5HKkdxcXhfOnlsUov4JqXAaUW88iSF1jUeSxirGH3ecEW2fU4AaAY
7oeymKcjTb9BYca0y3HWjhxRyvpmMrBRMU5XEsx3aM92tAgIgC56ypFFSh93Q92n
2E3ceeqmvw5gwTAiDuV93xh0/wylUE48PfiYK5R3LZo99BLFBovsqgvjs4DQk/hW
v1Xd1xCzjNaoCp/mlIFc8eKajyK+GT7YeUgm5J4KxNgJcMIOlGUO0B+wbqqi9dVd
jPwYxH/Kke+hbfk3LewllKB/sdPVkgVRJ0Y6Tk+sG4+MiCh/8u5f4fpq8bhGfJK6
1uaZxd8xYsAVRZ0VKXHvT9o/PlQJ3cxZK1/KA+zUKg+EgYx9apGDYygUAJ/GgJxx
hivuhssrJlsnozUFmYpCRYL1qa1bRnYT6w08YqS5VNlynyTnuB2X9AKvpyeZusQA
gOReBTT4dPqMxZoxUedTL4iBnQypYb8QTQRBNOFr75MK39brKhR2lAxPkG2MdmWG
dobyBn5FqfWP24FZ+3EjqASMQByat6RIyd+lyCMN3IjoMNrfC/TM2Oc1b+hTyJ+i
hdfMLprWAIEBNma2nwlvttzigTOL5byR7kaJsJA867kr8M1096T5Nu4kMXZ1rb87
rV3FyZP0FNfZ6oNOKq1GXjOiBspWGvgO5XmLKMCkL2CZd2eqIKuZb6aF6ZZBlvTc
blU34W1WfAfIV8CV4no3vMMhFBStldQ1OhujaR0bNEBBo0Kbu1ndYarKzVmesgp/
jKcx9Z5vTGLfwsMFDmNjjq8+Y6m7KCC6TNyQDdxuum/iQiDvf35jHexy4pXTwhk6
za/Nh7lnST3cUqpYrzxL/UhIMEm9tZCAgULwv+h13x+YjX+rrUDI8OZnjNn4NGVk
mVI88HJstaRNbOWUfnObaQtKx1IrRc6OynLVsecYcW0eXKgMLjbV4b3m5I6u7Hh2
g5yAn+0Qyv6VhrZelHFM/ltBVivFBvXum17QtsBndZUnD/mbMj8DKaSKSc0hbiev
HgSHR2tHuBYi73tZ9JB5APXlPg7bSI2xLaDipvubC6Lw6N8acftBBLW9t7tsueup
k255lLajU2KPxy4TaG4WQSD2ye9UDZP6osmDQH6lKS1bSSs3gHY6avIoTd2iXYa7
2gtyN1xk0IkalUg8BCo4shR8EpmJzSF1tQd7p+IqZh7kureAf5ghhzTckzjQwsvf
JAF/bC/cp48nAq8u0ucpESd9s82ND9JAeFZ0x5mD3Lh21LZSOFc/KcHh7ZSCzUl4
3KpY2Minf4T4Xi1eJtgDbr9cS0b7w7b2C9SGpOsd0vDgt8KdPUSNpTzovgS7yMBZ
7KveVb56oKVzMW83/Hp8B1RFHXOgvqC/dchcVMlvwMAo9OcqWqUHCasbwxolgOdx
l8n1Tc8OjAHF5Nmhp6DBcJTBrgnNwxPuy/88760bVJWrw4GV/SybFUBtgkAWOH2/
9vfoYvG0kwIULgrZ5hOcEuTgZRDIu3+3v7GHVpi2ylI1WZV0qOfDfZw9VWkO04FW
rQg4GHF1Bl1wGxYBQ+bZxK+tFMPzdp/QFgYCkbVoPY5ASGBUrEMCrVMJOtREkt5q
HjdETPDTwArSMP5ZyErLH5y/Eh9uiIhQ+0FOT2jp4J3BrJ7Q0asqyv5s/bx96HeR
SaK72zctJU0DrIs+ljCQxCHNHZTO6mU8rrZ2UFiWgXw/n4Nd+sf9NCgm445JEA4E
4MUkyJxPBAzrzMgO50w+kjfLahOusESK0LIreCO0j03Fur4p6WWLlK1yZDCQh9UY
H1D2RWzxnPenJUCPt2VA1ykSVLGnZ+GHle05I4abZAK9wJT8SuxUZ7Y7bfp/sJPo
IAcCGxyDr3oQO2kihAEhM4oE10CazD3NoA7SJ7vrsqUIqpDuW87j8/Rikjlzay0y
u4dmQoWQw0QH63PHbykXSKfG4r90iCg67JFBbC75+JZkXw3Wl+aLY36CiuSQ05+O
KWx6X1jdNPEsBS9tZ/k0uUJtY5pK7/k9JEkWeXkDLrZfudXFS2m4DjigkiNAM0nQ
yNb0j1r4kR8ugEaZ62lTFxE/e9naWy0mEWs+Wk715HWsWDjuWN4v8m8RJ3MjdR19
AsEXoD4rtPS5Z7ChbShwER8APJdYL24gJ75jKICFWU4IXwrNEqNVi5utwTvocZwd
L1DJyfgnWIF86bEq23IGmGxOPEsApQ32DM8ionKtjZsYfPZKpT12Q0nBzsM+9ZQe
4Y9KkAkPWyUVwK6N+NQ4rkNyU07iPaASFHSS8fvnbagPF7n/z/ovx3hTFsYke5oI
1U6r4G7EycAtCyDQdb+OVPLcMXFIP3ZkslQVxYTM9tB0opo/ydx2N7+6fSRZCTK9
zvJqJ6tskVGcTSQYxiA5XnxvfEswPcmstQkMdx4eBJpoVHxw/dvcK8kqir6beRZW
BR2rhLbCdMGYrkARqEmLKFaAH44xn40kVxWmdKYb3W55mrpGuckyqnq5M6LMh+IT
fgBc87OQiDPCLGKo2Da7PbZ1aMHQVEXUg2TDJbHuK0Kr7m2FxXQPAGvS2SJ3BQl6
rrlgQxrzSRr3TDTHTfrZif8nCZ1zW60ONE2LsGvfAYn3hiwQcQLgSyKI4GldFc6v
YtO1mep/8BspnYg9NNgXk8g8NatIaNXIrxnK8ngMN8dW+5KVysWhFZXEB5Gy/DYG
DF0BE1zwyQD5zxffMnFYWxoFz3yfy6veh4DHEyiTdbLwQLGafKidWiOpHoS5hOgG
pAHQbfiF5vKt8M4fugSG1Elf9rAdRw6xt+QGEgzCHZAvyFqzaD6P+mq+383O+Mly
2LYt7nfmgQPLYf/SQ4Gt2kck8gY2/4sC01rQqhkKB4Pq7LQh0VbvaPEmIf1QSI46
bfVd7Q592A4fmr4fIJXGAmybXJTe37hDBvxIlcNFiLwqVYURBjyRTlFEmak7UgTj
7CSUneEOhMilYwqakvt4up0Upn4PkI7jyNhCIY648eqmSN5t2x8Rsn0Ns1zKaLXB
ioEL5ItVXmfBRon3FpwhHWx2evQTELqbq+GuurOjGf6VoqJAjGxeAEJyiPyUaVok
ZYY0IaX0z4c4e0xthrrPjG7MiwtwvmBBp0txar0sxp5l/O4ZtE6ARTxZtyhMdFBF
iB2p0xzR+Xv5j8KnP/gm/TDkXZQhbFDxk/qXe2bjgcga1Ynx+wMZbXmnr+U+TGfz
8AjvV9lIGtG+xzh9+h6d1vob17nKDJPP6hnKyE+L72JXyOiYrLc5vf9afWw1OG4f
7PkXMFfyO1n3YOU2rxZBqwta/JBEU/gazMhuPi0ux1WL6Kk+tykc+EMwJpbFdOX+
jPoWTIGW7fRbyKtYPzldrMDKluRnfZiaX+lkZ3tPS2cAzvw4O7Gquob8belLGf91
ZxceDN1WzSKYgj0WdE19yaRaZ/0JiHsXlRHoDgoAuMPRgHEpKha2rnjXSkXLD36o
GWknDqdneXw9VLUnxvBOOr08HPneFItIwUlPNt8mc2UZ17Nd9mWfSa56+q4HZwT1
8aL1VawM1U0YmtXvyIYMHplx+Yv64aelpvFeWNgAj+HqtC7zGKxu2upm5t9S3NEL
TnPBNkTvKtOOXC5YqSIp4pyENO+s54+KMlsNOOKF2Xy3U6t3Ug4y0/XxoZ5C4EtX
iuLN5yv7YdTHXUVYi5+DPBoHXghKWUueN3tftqK2Y3tnLIhaP6Ia0DhTCEQd3kpg
YqBslu9zFhxzr5uwWxg1/XY2S0WMNSqZ8a++23S7DTGqfr4qyivrw5MfoKqGUXYw
ms8HAbw5QL7NljE4OIMmoecGf9BWNtmfs3uE/ve6k54fP7Ef+JGDJFfV6IOBlblw
WUr0kBK+nXyRHZ43PDUsCXGxVyL3xjS4gCvtfP5gmFAkVcg6ShlsySRYY5S6iaB6
cnTZHWrZe2+HeHFtlkuHWlUwqRutRDr4ttz+FHEKsTChM46cNZjdXDuFm4Hrar95
0INLHwn6x6eIyIPPLkKJJdHyzw9dZ0zfxXvMK4Il/mcsek4A44OmKjLMEU0MZwAx
XfrYmzF8Hy4BdfDwpabrTde3FGPeqIZsIF2/ftaK+dDZNN8K/5juhY5ykuf4hvIo
BDxrhFpHiuE2WQb1CxUjMi5OsvH82oTFIWwdyXDH3hWKuJYXIfcIxKvkaz4Rv/2t
F/E+NVOLaNxdM/6l1VGKVJoikkCj7Bfcc8tav+9R9w1noWWUUFqZYdP7YCe3b2d+
a6novHq9Scun7Yr1kd8ODNr4wf5TJ0iuvG5IV+ozsUhmlYqUWvKYUASrsh8TW/y+
GDnzp26uS01oxU8uBOvNiWnLUVDw0V+zzUo7pUfnohFLiHYaTOqMulFbKQHkr2Wp
CCbtGxkwuLgwa5HKtVS8HdpGmx8YPvHTiml5ZMIfDlSe0jL4q3iRXgOKMVyOaFRe
mJBxWj3MK3eb2OxELu737ceAdH7dtgjYGPvdGshnuONjjYUbwOhluYNdrJjeHf/j
TxRAqHezl1+IuDzNkS0S/HCGDIWcilrSTdtGr/whEkqIgVqVQd1jsydvxEmj5Wbn
DDXRqHIKZHMZ4AFhncrhkNrQk1RiYivUQKX36pQkU33wshUF60/FvROYUfs88eu6
af0I6wr79dXykCwi9EHRqZZQhws8cXqs5CWC1buHnA8OExl9337xAQHFqcGjhnw7
JM7Y5E9sQlj5UWo++fQgiAG7xMkTVQWAZRTSUJwtJKUgF+X0NQJnkDBTFiDuo5DX
8AtQ1zxNgfmtgt1SyrwPK6m/+yvEVLk73trNyW2pcpvm0hXapgq9psaVRoyFqjmv
KOZF7EqE0A6yHr7iK4+kbxxFnA2f/Sfn6Fg9PtNlKKMqr5vxPZk7CndYcPSorshq
NuPwhJrDyahK+l/NgT9qDooSgwpidytR3QWif2ynzL6c8JlpH7Z7F+/o/FDXhmff
gaY5W4au0JdGBEqN4x/pL+9Ye10P81w/ZnzUAZAtVFV623CEuk/FZeS0E8V7kz0R
yfmmcgPDKRjTU7bcMNWHuiFCQaf+FayJ/QRVpOJoyq/daaY9KSmPhMBml4f2YGwR
8Xx8he7YM0hXJOiZeva1aU1362cQTJupud/VHerEuxVx37KYoZHp/aFkxxNIOeXz
ZhtRDTBEGvE0LE6/H0zfcxxoDwgKWf4/DzRoBFgP0yPAhmB7PergZRuh+I/889HK
4jwzlyZeR1WwwgP7h2ximelQQaq+fYe2IP7Pyrq+7GeATUmEQeJIJrevfVzYAFll
SqJGTL5R3gsaJewT4PU8Jg5oKyA30QFeeImD4fJuZASLawXgGPyT4BJsPOdqB7kO
4jZ5uNyGm46xKALmAGQ1lDS6F7n9lV+sXGLDzBoZ3nXG39oI12Bk+1mA+4KXaBWD
JqREyd+tdljGeVIJelN0AdKXW2DrP6IhFPQ9/8YGbTkMKRiHdOhu7YE6DKYNpHWl
EJTLowPl5rIA21JfDVjmEvRzZqpmrANv4oUZ1BbED/5xtZHlWf1E7irxlv1rjuJ0
82DhEVsIqWg5qFskHZ6rgrvIMJlS11KjJXJCVVbx1jOBROS2imsk/iSgtS21itlB
Nqb8SaBqIdQykijnBaafoqBjLUmClD2fBMU3Az1HTG10kpeCyg6xaglmJ+hFXwvh
sVbZK3Tga0Tz1+dgq5dUOd8tNb1eYbUgdlBAENUao4Rnt75JIMQFgzUdBDHLlFgy
WsIL6M4P/cxopLXxUJo74iUuAErMtTAONs0Fg5F7Jq3b0zmcb67dDQMNiR5VxHeC
E19kjvFhX6sA8/NT9mksBA9kOM6AylH5Zu7VholPTNacRMKxTj+gNndrKXD7uZDf
msvMVZRYr4y3J5ll9YszaFU/vrNCofCga4jhb66L1lpyLu1HeSiHWFu3ExmRGRb/
VDv1Oohg1eup1PW9z1mwkTsTBTN297h1kS2YCXyTQtXb6mFuKt2LW7SptHAySo0M
eTef5p2ucnlSYL0zdOK33nSvoID+y8iVpGMzmcihA9mkpxeMtVq+qdChk23dEBEz
07HK4TEG+BKwB6y/lktBIJZTFRTgAPnS36dHf541Lz1Xy9EPe4OS/h16r27KtsB0
XqQat8s/YN1QjjUfcP7ohcQzZvusxu2nokiD+TTx2SgKeiEGVX/KR59n+/ys1UoP
dxpDAdaEPedhv5iysqXCLOWRMTE+Jb5l7mYEnDBAgr/LDRAjsXhrpMvQ8kJ45cnN
e+K4SGnKVFKyTQ8iWBpR6YRSruRo7HUFg7x21hDGst2nlDUy/IA08G7wQmliXjjU
sYGHLeDf9+lYfapq5J+yId2tG0UZfzlVQbBvvJJ/2YIWj30yWWv7a49fk7eGyUp+
LnGyQTv9Ieg+eXq5LTr5+blanusxVuZBWVh16Xj0T6ETsRzEZl7fayorl5EiNF45
RNqvT2sFw66gBVCUad7ca2pv/2qCzfjCKW4SEU9Fam6ARphoAiwsJsJ3RVqgLFd7
i/255IuotDfW7fKBy9oLMR8Xd5rnFcdtbN8KTV+LyEhrAOAynnD8NwDZircDi5DK
mU9QJfqdcYjCOo4R/UNQkmBCNznlQFEkRyfyn2fj++hNZf4x6QapMIgu6A0Avj4t
90vh+Tp2INPi860dyPypB+jnrBVxf7+AWGUBQh98Y7p20YdnhaHQYeQB4heR/2my
xTJuCm7udNtZQPpLqOMhpR42RNlmBBWv0nK1TWOPOd8hH3IZWUXzTkLmnNel5Ntz
G4eUlqklgGn3bzAazdQCkAoQVFGTlUI8dxdbHDQMyNeFQ2100NvhtvTHWv6TWrPZ
TZRChNrT7Ly/WE+oMx4ikzamRxMzenlYO6fMJ13fagFbP00vS20E6H8kXKu8Rbah
898q9CJ9V3yPhl84quvNEJhB9kA3gjHhX0QpKO8bgzJ1RFM4EA3fc+N/1Ct5D23w
mJkSFmtdDjKu6JUihWeKmkswDOfGaPnd/fdZwIPLkqZk871eJI8lTqQ6/2Gkdtwb
E+2n9/C9o0cXZYxWk0s3IhySgdroZxhy75FVSITX9Y4ompx7tLmjw0JJrD2/yJyq
2Qc5TsHtAY95uEOHmDu3vA4LGMB5XfHg4tQpi5P2+QkFs1eWLI6ZqE7q5gCS//4S
VqQ2Z+rkgcBilk67/qpfGvHbiITI+xEY7qfHc719D14HoWRHcdeYO9X2Wlyyxxdc
w0iF5zFNtyfQOoIxvxjkivD1xuog4FRPu9NBxNM2dkY8XRxhkJgEPMuh3jd7J8NP
hqJypyqNFdzUoORvMNa2JYRdsAVstk8yyQ+sI7eX0ukcFR84gCHP3FSDxkG1VoBS
TjVUs+JQLtTeGv+z+VH4xUj3Jt5UtwvWIyX+ba5t0LxsL46Rij43NdXRmZDfCCOB
HMzFURMT65A6FJwdzb8RL2Dwk9/u4dIKtB89XC9tmjaELfCK+PSTiaZgmulF71Rq
uK9PBZMXH6qiZob439K5gVwOF6CSOKvlx0VSbwy1tqO4L4QdIKLKO4VFlUVn/DU2
34cwoSf3FvgtQKTPwww5EIKzkJrgKzyRQMr1XKEqA5OZvhEKEAAqNnxPFplFZB2D
HdF99U/WsaYFzKpQ4KfP/8Exu9mbZ+SGwDEAJRnw2g4Uk7uj2c09LJrWOd0aWcR0
tMLwltvbJFPKnyH/TH4h4eTbhVoSq+V1QFrGKfU1t1lJstlYRdy1ApkEKMj8Y1PM
hXZ8c0nSm1iiewErcsC9lJGRjfB5sIGgfEXSo8jzmWqKkTq9KbMZsAkY0VCFqK1w
4AmptjkqNU866m9tMSfS9Rfa1s5Xy3nC0i0lCOwx+RKVM4MJUIou91joIzJe5Ozo
JBUnPTxlDjSnZMeddD27pYKv4a3Kj4BnatrP3dOq8HhtgUi3Taew+AhXLR7dd59M
BIGqN7Wbgju4PYvJZe6j4GtASGoCWM/Jex4RYMBoeR5O0o5qeZbiwbML5RcqWP0A
j9Q1PEoTvsTt7hot4e1XhZVLg0TZYgrkuqF53qvyc6h3wGO5HNUgVmwPcH0V/9Mz
7qo9XeZ3n04sB4xjrqdw6chIhQdyoWTRXGo0paWDPRWEXMlh00r2GjXczeqAo9my
3ccPuiYKFDGVEsO4S+0T4bPRxUi3p6pSyefst7mOTtBOvWvkRgi5pR8c3ueh19MG
L8AO+HyfQ7pqPvUERff7u3QBYlTdqMI25hPMnvfGTa3wU45hTjyk+TAhpuCko1HO
hsvJCWb391BE5LXoAJqlhbR0Xdgx4PufUQ1DhnKFhVIFMGr1tfMVsgwRTqgESdAe
fkF0X2t/qHzGPTLX68RhSVEC7tV/H79yBQAUGCQlMt3jQWlzafhyCUEY91n2Rdsy
PaFkQPcAZL1BU/y7KsZZ97PLdogx/k/wPB1JwO0inocecLGwCN85xZ0bioekruTP
e0YuJ8UMojUyp6dPGsoIlzGYPxFEYz37t3UFUpNP3ivcDERodUGvUPKmYJ4ZvaXb
l/sB4b4qFn4kLbExNlHBqeQZretU9F3Eg0ta9iIpm8RTX9JUcVD/hGds8h8D05/L
4jjAjJPOsAzDctgJcQONOmTvDy90CVxkU6MWynrrumlsbfw4Qro1A+IeZLw4IIsa
Jom8lb58era4F3+e/8MDL7QaodmrRH54oO8tvQ+1M+2u/wKuXI9WL/4j3rkF4fru
cZTyc6lHby8nGdyCKZm6SJt2g8Zu4FdiqVo198Cf18dhHKq7TkhRvGIbtF2NAU73
ujqJWQ0OX8lIEkbnMemIvqQF1tKcwPOKwjb5mdGq/s3DKgRiNFCH/vZ1nbhUyP6A
JVmSlrE2OjW6omtSalRJ1bIlR8inQ4xgBtTOW+1VSAKsgz4CRgftLkJtYOPXmRw5
67dGDVULCzj7gB875UERJWl2AR01+867a25WykZceBbTiaEzwf9HOtyrXMG30zCq
rWIhI44xSbVpQqzlaHwqJsKUkN7DpVglnQc5G2mi5T41IzgDGEtwvGoU+rF+GNt6
ecIhvtjdC6gdcps6ROXeNlMooK583V61SSrT/1A858kDYT6dFHVqIerBA2wGyvAU
bcYNdMT5EvOhMLB5y1QbAyAmUncoUoIM0cWi5CLKifTSWm1o71zmtZ4WOr5LwuQi
q/FUASciUC6XSezhykbq4oMLYiH1IFdZC9G1TRro4ISArS5gDw8uK70GsHttL6Wb
NM7Y87xVTpffTOia60zE8YnXDnsB90RtOerR34LBjIO0DYHebaNH/RjDyiksRpUR
ugHtlntCHN9UA3/4FM2fBjmdICtqFWwnBA74Dy06dt1GTkcujFXsZgIUP/xv8yF9
ODCOcGoUGXmLiUBgfeSMZ/DD9w0j92V76bewxmlAfkazwRFVzxO2/PjW5dAW2Ue5
/kGqDRdAdOqzvs7F4mD42A9YJLRg2srgqSAxSCt61BkECYf8OvktRJqQhyrDLiYe
9NQ0Wg5r7wTQNTRUzdCi7/G3MLmydsRl4mJXgDCudJMGgXgoir6BXAd2u4WIuE3/
zPV/Klyfr2yxOXX7BmxWQL7ei1x1uEG7YaclUmBRmTaDSx8YP/zzDeIKVuIW8e7I
6sQHJOuKfMyb1jo0olC869Ov6Ev1zekGviqkH/CvMb2XRmeACNHNIxCCzoizfJfv
/hKmdYj3n5l14rWk4bpZlugSQa7fajJDjudv16sfVytpakqiItxWBfXCwjwDe8kS
SbXq1KV6XVwCVDfqZyXCqG43ZsRU2noZd3XoGvKlFtGkuSJ+SyWn8vf4yjbsTW+i
onwQrSAnJkBl9U8+MBc5W0TNJAOJPPnljGibX9qKatJunidtA5TJf600redugHNt
gOJZFZ2prQPrzjoiAx3LgUwx95VhPq6Cleu9hu/Ekny9bZQKKrVICPUUMwppL8cw
kgy2GF37ku+5EElDHd/D3v5fQF92XdsXzczl3ZTPdQj6bZn4waj1H4GahpjAzaBh
6l/YLSlO3s3yQeR3yHE9IlywZj63mvJcUsxcBbOW2Vh1FxXYnjdsL9SJyzzmaQQJ
3tgsZ4Abiw18sr/1NBMHnCAQx4ve2AGFmQ3x70l84YZ0RsI1deq+4xCZLoftpqeM
YFjR7KNZMX6AonaJUShtvRZ8BLJGSWdofXsZYK/7Y4a209p5H2liESebDzQ9wW0a
Nx8MoY2ajxbZ4ieN/efIDq3jqnyssw6vWlpw9oum4SYNcy9nxO1mLuluXJRCMhMF
cH6d0nT0XGYwBqgEcPoVB26eeJaEj3VkM4vMzDWLmdEcKgjLIXs0cAQzMWax2hKD
oH9lg3h0QqLKvpRhtIk7z++pIbdrBKBPSqG/WKhYfRFeFllqyKQ2PpW3PdK5+eLa
iL3+cXMp8vVquGpo/IdyuxVBsUrq7oYsZgtdJcMdjhAJaH7OGe9XWs9wkNkUZ6PY
DOrLpxIM7PDOZ0gbIRieaCtZqQyLFO4rgzAGMQ4UDNkXoilOKeJzaitY56iDYYEv
jR6+KldQWXqysdqUYoqGPWo+Up7L06szeN0H1Op70W4Qy5S3Jgreofv9xwu9H5XG
4Ww0AW4e5r2CWHz42UZ6Zb2UYdNOdMBvl/C/sYiXQbsBd5d8hxeJRW7lvTqFveTo
M0JsgVPUcsQmPqOuviQhIcKXFBHDlmdP2d10It45/YWXQinh4AMdUpvnS+X4XLyl
ylJtqzHxgk0NotW1ch0/odaJtAUTGvXKeoqGJ/GsgmGAEkNn2Zfyps7JZkrd+NTw
X/+tORh5jntv7/BIWr4VUdb0G2FWpsl/qdazPJQ39Ygi1sbY2Dkxe498rmrgL0xj
kVKsG8AnngUiID2yVT+g3QIbBJckJdMRMzTRHsy4OXwjfwNMotlWhu3WWIXSNv3z
0LFFbiqzZkBQBtr4g1IfC9bchsDCluhs/O1jxep+o+X4MmHXzH20npdhULCO0ZQz
CB77m37xh8XT9qEoIuWu6+gOptPdKG7PibUE4WKFeKZhYfDQh6OiH39BDiNGVREp
IgZPUMHzQuJTcoYfgB34JHDXRX8FzjCSClXtoQYhL2rb7KBVDpQ148svJ+OngaG0
RyzcIc7rpPfcQoSCEmUGvCN1Evlt0xBCx+qDDajmJtmxFsXUad8vQBfDeeGtwfx4
M0fJWg/v2dNVS4F2iwkuDjCRQlSy9lECdMeCg2rX17VAFmuxa1jRssFme+Lr/y68
7gi56Y9CASKzKa8jR7r+EzVDmWXiT78/x6DUGv0bqudEE5n5of/un8LOskLhfDxi
XqpnapgqnMtMrrzV8jF/HVXdj5XEOY2Y6oMEA0D+ahy9uKB556BxM3lZ6V/xIiUS
6ZZW2IS1zgE7GW1FumrT+bvaNDtYKDekbsQgadPM5THJiAF969X1WZIe7LYhkXfh
H+lBcNVOzEAj2VIqtiB7BE8a6ZeHGduFTy2vyGUe886q0WdIfqAxBGg2Dj5ysPch
oSPVgZpCS6Aty+l2D5zjYrfDygjVer28QuujAP1iLljucg31cfKsfQzyh7+YbeHk
uopKCA+x4lqlaTd9RtlxR4P7JLHt/AU9oPXOJEzqFaGLedWk4970MzPv64sf3Tk6
po12HKufRlqokl3gCoIEpwVtqaPHx8uNgpqMsi5bg/a2m58OaZQnAPTZBGh5DoiJ
fjhU9iLevCR7KfcmrNVp72LWtZ+1DmSgcuP/geX4/1CY1uBBqVbV64JHDWxXz7Ri
QKQikDX5uEIEOJEhpqPsFFaLacP1IiABx86p6dLlufa3NPa9XB6kNqMqeOnqEPQj
nSzd3i1w2MrrH0jJR7iQbrkEBAkCmkXgOmwlH3bNBm7lFvDzUp94hED1HJdeBQ6P
T0Uv2z2lA3n3dAjQWhol5PO97UzQV8WBYeTWuPXTX4mWM7XXYnBU+b2B00hk5JYw
DnLSA50ThljIqeeRNZTldUCXZ3Yf7JChcj3AVDgZPNyqWL/HJRHXExYaNR/ioHC1
41tFWV95Jwt6631uz5ucePjbrTAnY5YmQ6K5bZvd+Gl5WkpQnWXhWkZUTMwhi4sk
r4ZCrvuxYb8NtA14edDiqJoH1IxAP95ck/cMSs2ej2epqIIHFntqXh01d9q0JYGV
O7KYKDOgqywjv1yM+gNUsyQtP7Bb+6LSCUrWGC3EWrNXafi69ZovsBD0RFKz6cbR
1oYVc6R33dZofh1gZrSN0c+HNMMhmmQewgj5lhpwx8l8EY4oNT9Pl0hCkoz6WA19
HTpzNsksfCI2w8OnaqTHF1OnRx3BEErqZboQJAHgW+c01/zBNrU4geVrkZzYRwAb
AbXQCUdr1YPd+bw1TXWQXbYpT4MdKUN0I+P/GgPBFwRVzRl2yo0Z4A1DK92l3HLz
zcVtI57Q9ywMitk3Rqh9jwgZbdcFkriCHvXnWnVzLlAiDqO71zahOlRFncekL2Ff
mU7bV8BnCd9mIMyM+uySW1/HBrGVE/BKz8sDQqqA1yUjSB8vY8qQS8lUBu5JyhsT
yd271cf1fB9tJyhg6OxLCdH1eZCPw4Z2Ebf9/xpMcKW5si0UV3tyKbZ8D359bjX2
2g0WLtdzVkWXcciraT9cXqvI791S1OiXwXWuWFCWabrbCcmHTl7R9AO0qE8ZjscB
2o1g24+gXJ3e59OWNkBrPLoVSgHtWuaOgvWvfxE9dX4hod5sczLnPnw3j+FX6z2C
MAjxQF24fqSjrfgOQ5ulcQ9GNJ4szVweasHpgBbYOpeGN8zSyEwtixgqIzjzGi7W
DM11C2cmZU01kk20c+2j8Yujv7ZERZ40G6O3pCPKqF5dxcJBva9VonkhzC9Pu6vZ
YzD391BB+SLWsu88g3FrOUtbIH0b7F/OSSzYA0pOwRbsDU/jLrhMGxQcCY4Jyn62
eEd9pnTt82YkrSA+qOuBATXKrIStxQSzQLNWoX0YCAay27MzYV25vmwDMjjc0hHC
UzUFlykHpuSxljdveGG6ALywzNb5Md6OMjyfBtgo7T7ZE7gFh3mpd0cn5J7F1ffW
dNLJQNgEPrxNjdP3yPJiwi/F0a/ItvAztq5aN3Px3CvmbfRGceHDa4YJR354TSYe
Qxi214aEuv5VC+WBmrLqvTTLJt0bICCRG2TdCWI8iH+YBL1BFXTxdlSuXdF2EeWX
jMY3lgKTt+k7kvn5WSZfAbpzHq/Xp/ehvT6/MRuxtjW98noqT4TiE8YFRnieHK1w
LRdRJFfvpq99lUybipLM4UmNk3jminiuQg2kFfjHN1ByubDUfjCFdqJKiojGTnZQ
XSxU6fo+BVHPP3rK1cCBAkFYVNRYYSupMoum42dpEqKZveTwvwfeAlxfYi2vQ4sP
M2tZQwV+4NZDqeI+CeBe9Qq/sNZdZeA+OJo9bOLdR+nZ5AKoKIrG0j03HAuUfsCE
v57t2QFIx6Zlrk9jcV6OFifz9+7rF8BbLMltqcA42vjBXB/1Dm4At8//Oynotnop
xjWuQQnT3xH6wq4Przh6w+nY/9es6HuPS2db+qSKRIRtW6LPIUvwWl+k8QP1VDnw
GxLpIJdZzsEaUbttGX48cwH2rxQXE5VzWuQoXrg5dfcSta7P929HNhUjL52sSY4B
qMYMaRD6jPtzG7cY2PToh4gzOHJayZl46BdOMT6M8/FjCGe4a91qDrdLZ4jveouG
kzuvqhmz1HTsoy+L6aeNcm3lASxPvPoWRmzKCypCxF7vAoJhFogPjO8BoR5Ij+zA
Nzv/RkFCtTEs/22BToKgda6tLzqYH0gs6TQu4vX0hJIMPQi1ksy13fYs0FXMSD9s
HABVLODm5H3haTvpY4ifNnbUDMeYs8mo5zpNsMRGv6rQw612zN2eD3JNmq46skPA
qsboYTFlF1cpXP+CbW/J9vGyBoUq9IaIrLpuJkt72RPgdVIbpW+9vXsBNGexET78
htrEhZupmGgGyOSSqYAYTgHX3zhiIinqVoRCOoBogDe5PFzGBesfnGGZO9GLCv8O
vUV8Nvflv78qI2hQdrnvAGj+qcX0Ob8Y+PpW0JGTCZGyjXpDtJ6vUgjObQ7CHHdY
QJ0OjJwAGUF8Wfv+wySRrbW0yB7cQfu8wNfesGT7zRrF6DbIMyFSUm1Qvnl4WusZ
e09IiK7M2LWOrPL8ccvJqeXKQE2zybw1usA/X4zIeU1oApi64G2ZiGbs4Nhc0C6q
bGBIipL3jUlMGLmoIQ4NpmztHIca5Erai9nm97exP6BhKER4oP8bCzN5JQw/h+CU
HWMQaiBxwMT1mnBjWhmICnbkejwzZBX1VvGvMHQVgeaXHGvJXns31auhG/rZZWfK
HJBWoN2+SGUxnWkKLLftj4/eMfri4e2BjycJFKnlg0qTZEqIBw+krjxap3PSN4uY
g3/ceDf1xP8rNtTXN2ptdojtHq8p5AQfZJyYudGd1KD9KxppktKW+zcREelXMQnJ
IiIwZhVDXo1TohPySGsJVYY6Ksjt19F7XaLZSq5ZmYYJpDmQ0e6PiToGrgvLj0rF
K66LjKh7y/4nyhWnJyHSY6l1dKf8HlSr+HQ6/qPlZsicHfnT4FYjNHVIfw9LRwO4
SdpPmPyJEfH4kHmoKcMLRp+OtKx0VhhA/zyiPR8FJIBqtOLw+zknhLiORQfHK/6d
Do0kw5mRLXMtajGKq2eiBC6XaKpoOgGDBxg+bigBl+0wWCXVK2SALySRauZEPLQw
2pp+x5qCs9ZpVhKz8nnu7AHZ0nu0tf3JTlw0Z3OaRFlOV9gepZj7Vb5oi8xPWz9y
k9x/J4FuW57jxB5ruptRC6YJ31Lt+q7UKwt4d7zRJFNvztkTeOPEpPekYZPQWyqw
0C60GJd3bosgnnDMyLlyDwmklsGEYfUmYocvgwXUbIx+UyZx4P3BIIsyd8TsPPLt
gt62rss7Lyj3XvPBdczfbcs1pwxQJhcZPYkluzwxAvgCQhuvi/GabmJ3BOqK3cKl
w31OJJ4jgJqfcTkVry844IhTvGUh9ZrsLuAVEmsVMWOjEJUpOi13gH8pgic9R2ho
kf6vnmJpGMHqiEn0YbLJGwDDfvg/NLSC56OCn07Ngbux1scz/j2XY1MFUt0Hg8Da
rWj6aHguhhMMImBNjJea7HkgOBhVO1y8GSxA2ahvn08sXkjoMoOEONj3t7wrr4zy
oVpRCHJfk2c8rVX9W46W097Q9KeGHDJ+WaD+582uhyyFEyXoI9WPTMNw1IwIbe0l
MqJlzsqs77LQFHE7mFDNJidh+DRuHfWGtGGD7/3rcl0dZGU5ywWTJ0lmWcutVURX
a++3HbsJVy0T1qB5IKupf6h3w1tr9MYIw9JxqkWMigFT1iIrk2/7K8VWPOFl8IsM
l2squWlPU3ZUfEuOYLB+8ZpC6DCIm8YC86iptnhtI+eiOSa1tUAJF1yROVuPR9AG
N8cUmGEJ01imE9eE3mNpj4TRNS024uzM2HxPEloy2kbuZAU3+2J2PHDP/vjP9Lhb
fdpgJelniEXY71QdCThW1vncElVMcxq77R2Nb8Py1R4lCzdr8C8tjw8lMjAdc+f+
HKG5IHekwFF5nApgbqyFn5ctMDwB/nZ0SDOvwb9caIXkwU19OpCCv3GyIfQ+KLYS
4acdmFqKAbxJgI1pkjDnb/ApMvsFWllDomrpUX+UjYgGB+yZu8ZNtoB/DLwnc0QG
xRPYnunXGO/zrvN+KVTiUWTvxS7SVA+XJA3rphTCaOjsSqRCTm4ljB8xqv0910FS
tcZ53UUJT38XyhTC9SXd41NGxpU+8LDFnNLjRHmudZpPDwd7a41dQeqDTjPovw8h
dX+d00+LYEHaKEHSVoFJkhObiI709kYG/pDNpjFo8XF/q2GLKNcS9NWiROHKIyEM
LkgYbb3WgtjRjKJe8Ol6w/hA+sWDpGw2JPiSag8tXj2lBxrlA0AtgQyRCaO9jNeE
fKV+vVEbOlwYwCMi/SyzKYIpfRXfHkaP0Ncn9DzIEFWNWA3CW8f55qLhTZe6jZYC
p1rOUmf1oPhP4JR9Btr+MwqFyqsQFg4ebzWSViIRBmv5rkGdmc/kSWfX21uTw5Kg
CEQE1b+78F/RlKO/HsFF+zqHKuzM4X/gLkn+NUro8WlSKZKY6aTQurqX+rMwVemc
w0THLzq2IUU+qxFdsn7LvpQOH2teUmnJB892HA+GeJsOTi9M9hu56ktuYkCQ5j3O
HfHyWofhKvmWvDI99c4OfFptOoHkXYb27AmXqtv22AY7/ATQTBfieKmiyPAtCN4z
o7t1saivVdm06QA4iSo1Ak16gKfUIMz9VVE14O9r55jUPSCZny5Av1/0oq/QygCJ
ka6mEoOPsEcB5e0Lhwq2Q/0PmsXyG1anzrmpTvAvkyNLQO4iEYXG08nIUZmpgDTi
aR/Opm78GJM62qJNtjwsqEzIGiCKoIiXL71pJKhxP5F1Wqi7H4vkq+oqbkvPnNGN
WGl96GapBpAgebu2H3yZkNbJZdJzCH812htr0Ojyfyp3OZI/ofZPtO0m7NsrKiE1
pAWmoxbix6KFY275yImf0kdDgfZsfvkCYShIaHlcrXjI1muGEdJKQU9/2EMIGc2g
Lchv5nuMghkCusCjaR7+0OZXiPxUmscO3eAKpqJo863tPu2+gRkpDNLd/1VYJ18O
zqgVIXDZgM0VzhNu3GT+iZF7WxS9ot0Sh4qr3vwr/UQilKy5yHTlExNhV6nEV+lr
EsdG9TuLVJvZrRNqDgfaKJ80sOuMoigYHcxm1zT/X5hPmRld/6sX+Fjcq1kzO0T3
K5PLDUGkpPLfu6NWlB0KPsceaAHALMt3etUzxsr52d817VUsLPcGzqVUNQKapgmc
AXWTPriru4ePLZk2zvbmdBpw9AbulGKxCRTVwz2P1DBubKcGjgYld6Ex8Ad12wp7
WvcS15yJ0rz8FbGB48QPlNEfRkL/E5Qs97QbFkr8ST7v9qHKZOLJWRJAnyH+GeI2
ZvB46oc550zTigIss4LxNvhZzcSAgDCt9T5SDOCHBv/1Z9WxTp3j37A5rzsiz3ND
ojPJ7LBFq6uZIrHpTp1QYVhnsv4Kd1QxcXEVEe5PCQ61or9zkXnRt5spGXVhMBU+
wY3UoKoCwUdLjMJbt30movW+76qWENEz31vwbMlYnrf8NOjeIaNeLUSjp2ZgUpQC
vC7YaOzVw+fMjGaidbT863WUCR2AkXdyloawh7YFmDxUIl+NaJTiKhqfknwjU8i2
WYyf4ZTnHqwc9UAOSg0GrPwMAa2Chu8c6ku/xqUkr9ziIMAp2a7R0BsS9rWJZy36
jokEOdJrDccpGN56tWz9y6pF/ELsNfFcPtrcbCIq5IhUivPCItZAsbSpXHd6tjot
wdeDAHMEnF/y3uI07jr2mIzuqtRP/I3fsghL4kovzZBNRGseGlj7+hP7fFDFzgyV
P6VBLzGmnwA2jEqmi+EZr+ZH/w8IA9ITlofM2pVhbHiSPkdyWzbjeXluhMs4t0ij
eJohht9TWEMKdv9af0n2xu8t2B2m7nUktpl+amPAYJCdar1ZxSgsSCAZhI7M69++
KmSn8cPaoHJXVpnX0ZiAQFNFnJYuUmjtTM3IkagRxovmmYkSWOxJrtOWvZwBq5i4
vFursWLcLT/B+bGJkyjBdQMOxXUD96AbE1gLIHAMxN1eYRX0QJkoyo9wWEHxO3jT
NNpfONnphlyWoJZEZ1fPdp8qv/Q5sWiOk6vRMAHrtE0o/g9UCjJ/gc0WHDo6cxVH
gxh+oxgenE2UUqEL3nRGU6fpJe0vjw56Z34ZNKqHtNOUi+z/9p07cjr0CcBlLjek
oclwn6UmPYlUi8rlDnhmEBXYSHic4weZWfLQRgmFecodx9Y3+D41K32dKLS04YTq
vJ1wDirtC7uK4GKl/dudHc3veJ3WskZMdrdwgMtpjqSGWCI2FwGaXNjwtLjFsgcD
dfIIKZOjRJ5K39uAMbsy2DkFnX/GTYYpPWgDhZjToef2kN7yCVyQ5rf+KED770Sx
pYKhsotDAaaYfK0Hl5MIq07jplXByMLuBG4YCPF5zNuxNS8eYWVJoYNOd7BKL/1L
I3Pb7cooCXKMuGiJZPfYmlcn5J7sbH2sdme/HmQkGK8GQLhvJS6BUqcVARQeV+Sy
OsWlf94tSCdlHaHXbJuJz4pIbmSy1CoI3otgiAAivvfNaQOm/ERajDBrxAfOc0ey
Cs3meO2+J2v5OBtHyI6tUyc4yf/GLAEeWBNEQNaATOCrz8sZ6yV4uE/KtTTnDi7/
bVSB3KskWjm9PcvBYptTuQ/xB0iiZ7gKn9pPqnnf3V+SDnEDxd8YXTcLAhMta+b2
uRoN4qfV9SagYqE6UOwr5FlFIyIatLXueGX+hOZr1ZFdVIig8PZU43oab6Woxgii
RUbpyfpBInRMmBOV+5vJ8y+6ekCpK/IuI2LdMzsgZ9FVow2+6sJ+IlBmy1YQXBj0
tRsULc9vpMV7CjmwMvjxgPIQ2tPpjVpLI7UG2r7wlD4xboEK7VJJr8B5bj2x5IAP
rB0ZlbA+uBsnmuFTaRQonLi/Ccc+lMr7E59cvKzqKH5/yPZuOHGloEdUAKhgm+by
mfB3PyRlLJCudlX+zv7D+Ldd4uSIf+5tH6+kFlRKvcTclpZPrSi1UmLVSte57S8P
UYSzWZHjkAUqpkXmtCzuntdkmEt4l4jeP9uPe45mPf0/ph5CCRpHyEmORm5ttgZT
FHZ3Hu4Vxmrv3bq3AgqtxR6FobSuiIW5DK53aXUVfYWyeqJ6PFy93t0AYZC4E7C1
9t+Rfpd1q6aL+SywPnn6+7c+vnTPtVRCfHMHY2VomLfnpMPUZk8KbfQpTNC9mdKi
iEmx5T8CZIV1cFcRuXCPQCjtpAZY+6D/8Lv1pRWDN9Z1AJZpH7teWmE9sPkdVkY2
Ahb6am1WL/RMI0LokO2ZkEA6UKXmVBbe/fcq17891GZuIzSaM5nWPMl9P6n7QXDd
zRjmz/j5S7yYh+6ns/HvdQ2hzshJM7LEFVP7n+lMwJO1BRj7xQqBnQ8n+giP4MhD
P4EMBAs/5k8gGjf3G5XVbN30Z9KnRUFPq2HMdXQkjVQWRUpwb2C5zzbKMA6Ay3OD
wJ+Zwr4uUiovOerZnwDPB7raexl5BjC04VRLfKxVx1vle+FvPJ0HFq1nEUSq73i6
UeRIdG4lgyft6fLrbZvvDXxe5GVCaxVLOFjvn6LUqEKiWgtT6PHVQq+/lpklMCJF
A12YSGyhrgi31Mul8bLrm54oSXclXxVMdBhLvnk7d+fNdHkeM4V0Rdq48fGaD2eZ
7VSs/hr0wCvp96ZpvxajWSOqe91TURoeLWkeoSO1Mg9pxJAN9XTlwv0Lie8j6Vs9
wymdeSV1DnZFjK4/rWqZhNEzJRl7ImAIMOu1I+onoJURPhgLELBXxmcB/pQd4P9x
oJk4u5hq2yd33FQzp4LqRoPRkjuqjIC6tdZf2TYO6i+XU4Jx1rwvyQmcqEQjmj9J
EvqQ0m4CLd2zKyLZjBuZyLzaC6lq9RjiDXmWmw2f6cQKUROLb8LAv5KG6LvqaKB0
jx0aQm6dVXkqJe4t6tWPpSMVSWyYOmOU0YMC91IB7Cte9gto5Bt/5lwD4VOBXvYb
vjuHct287mWFW4gAxRQrn5my8WYLnRBaeoeqTjhk6B9dI2Ff1RaUwif5SMWojAzy
GCuqxK3zQzZPIzmYRd2LCpkTuOMTJ+8CEhDVV/XLVZRD7BTsqKgWfXBcq/vYeoXC
MEWhmk8JYe1BW2ReeCyTAJf3vCVj+jFJ+taPlRdaSUQ4wb9Upn3Vo+0DL5UbdIxx
dKmzvpVyFDnMlt9oC3Iw/Y3ogCkTF70tLQKvKxYY0otZtZEApz9VHmkWSs1szh5i
PIjHUHM1dyi8P3iDAhIg76gybxJnsb2hnREwNE2I4CETD3k4VCdPUgtKeFmgfLA4
M9jG3Rte9lox7JyzceV3qWEIRTSOblyH7zyN9h8MWTMKyC+KiEYr9pg6MZPHhoxe
c5ahr9Xp6rxnbdFTuq2UgSFtu1Xr4QQF0IkUM/exFiGFqkcduKljKAGATqa6rQhV
xNI326xffZSa/4LVq5R8rniFRKO3bnbvG9D+sJu9H61kMzbzKLY/a523xwEglxvI
Prhjptwq8nqCesxPjg8mDyGjQAE5Y2TLzIVoWRNENFTyfaKN44Y0BDsyQAcd1ihv
6yujqW/Tk7yttybfk+ZTRPgYtm0dvQkYxSdVyp0GUumoj61zZu5M6rOGWSaEk7JM
+LNbqlsEqBheOtNS/F/8JmFM49Mc4D+/WtLhSCxy8Lrg9qHP9Q6MduyQSddS7wd0
KjHDVJ7hvL/Y2nvMhNoSRxzorjHeNJhLc0KR+CJkIQVDtIz4HLD26S3eR48tjTtR
EMMU0MBDZEWCV01wN609NzAtJYrvaXno9/61HvtlPqIP7aqWm5xsnSgWvW2Bl/MI
7H9RyhIo5ccKmJq5czUhFxup1Oi3+GS1kPQCYrft18SKQyFjysTcd0fF/KdmSPuA
vbD8OdnMhkyJpedSeY1wRDKE14G6qHSFMXR6QPj9XUASkPZZyz2HtEbp6AGQjt5U
2euRuysOYwbBP15uqAyj6rBV29HpUiQ7zlU3nfIx7zKAwzxg0tHx3g5QuPbwc59G
2XAF6anC+e8kB9FLMh2Iafs/qkbkFDO0/ERgDkmi6C7T6UI9qsyWpkeXVj8RZ0v/
jDtiJvzxvW9JhDL7lsEmkzUBA7ASA1vCB5B5CLYuI7FK4IR4W5Q2jOHqytJgZ3+9
8brr0XYoY6jI9yfYjXtFVaL+FUjVmJ/w0vbEk/1F1PbC1YChC00aR/IgcEHiL/x5
NVqFxKgArBjGtqHlDLbqSxAc5zZPY/K5v9a6fru3f88qyjAJafQcyqt8hcjpbFMF
DlrUVaYvgslvMj9RYwWD9vQemzppqn25DJM9HKHy0K+lNKb1M/auKl5uIw1ZyMM6
bA7CgmIdY+HBBJKVuWAy9ln5r6otcaLy8IFxGgMGGBY/TYUyEb0nECTbfD29BYsQ
UQosrZ+hTyKPa8P9LUUrZpjPYRSsIrW5MY0eDp1HyprseHl9IF30lR1MYVAiL4C9
q42X7XRYXTOWsKbzU6DmvkR7HZAxnZmz3f8rSpezUX+i3bHxi1FkoJ2M7MSytSg9
5CoksO20lwruP2ISuFJ3XE51+WjHZaR1wlH+QJaDz7ltzMZjpHnDabOZY4EFOLA1
YA+02OW2jzRpQN3SJR39VLsYWhMQH6vufMSa3++dNhYU/MUrx3RV8DVD2LTbxXwg
5gTwZYV5gXUFtSQsvZSIv/97rhGV6Wx2pq/OtMscVHkPv+1pThyjRuzZheNp4m6R
nvKKA0eMKhy1bl/6gvzct1XjrSznmELzh+b37yrU/GCC194bV6wCZnaUcbNcfTxn
V3HhWMHWoG0DoCdLEghzBPzddLRriRoW/VJtrB89qZQBS7B5llPKZCUG1Zt02lFG
eBptignQ1RvYa51AYDybDtCpYhCRej5oIqHD2rqsv9eYxM0cO3qEO6MbYSQGgSQK
ojC/4m8IuyHNpmsw19//yKKrkhldn8zzbQdYGEZxE4CRWUHQIcN5OhFBs3kVNKCy
7lM7CYKAjU6bDHSdgc3FXxx6F5xfKurmgniewwJJtnu5wE4+bpnhraiY/aiUJsxX
2IgyR0RFz6cEmof5Ofm5h0672vz9zViOsh6RhjPMqduPIySZr9I4CC3JSawdiRmV
+Kd0RsSOz+yhx+/b9rqSrpaVmceWbbvHZL5PgBvkzOlFwi2YTmbvQ6166gp65qOp
AErs9gV7JAk+tDYBTrrjpoQZs7UlEGJMA7KXFA18tLD2mQfYmnfquTnb/QNGgVY7
YnAt30ZlNUFG5N4TZQ4L8KnH50FUUeHTVA6Db100SadQl34THbVGVaf87hXdukQh
yBAWy+11GdaXvyHwAmPXPnGKyUpS5acwWJCGwtepsJf+9Lg0t8CvI8u3MAzKljJ5
SFeoF4ymZIZugMGC8JmHC7NmDZ+mJgH114Xi6ok2hNaos02bVKaj1OAf4Zsni9NO
Au2KWBYPrWVqO2yrrfCwXcQurU4YT/wUtEaI0AYWEx+LEXKGAkK+AxyIir4DZhAa
yM4QBD/cRigpxnqulMPKw45kbXvDRG5UoFJCH696AuEPo/slxJNGuWHNwkQt72ku
hBl8jXUAKOmYqY5NOqLp31GMGhyRLdpXCcOBBWflS4/ulBKkrM5Bjp+PRt9X3EIr
q4QSTZk519FGz/CxLmaUYQE/lBm7O3vnESyA2XOGvuZTqEnxIYHDnyMTz0CYIRjA
K2mafP/TFizPvbzLmuHQKXZcI+cUmxV83HiHXW/6r0Xz2Fjoaj1f492dHIaqzfKw
mwL9EIP3yTYeS8Q6S7fv0DIZw/7dsBiBA6T/8Kuw4MrwMjdB/9nR/YD1AQzJgjgh
NQ8ednPyHbwz21x4Dt+NrzTvHpJ0s/vT8rLmhOHXrnyJDHSg0aaVa1iBv/M1ZlbO
xttip8tL2eoE53sYwtzJ30DnvNVuYBJddnUlyrLWnQNwmabGqI5LkXcI3HeMNkse
wNCf0e5hzcv3K3KD5HCEY+hSZWo0ZWYlOU6HhdlncPuRBkSo9PHHHnQQBefoE54A
e77rK0xfIFsek9lDSNlhqQh6Y45LW8SEita7bqWMu1p1tSuoG8beFIvzL5XiCtzq
LVHyY9bZZaGiZ8QYNWEBFnfrg2gfbUEybApner6VF5h8S72BM3StxOaqsHF1dodG
ILnMspyjD5NP3RqEaeIGzXAIzfZgV0u+sA629Hhm16ayXFJnOoTkDVN3ZrkL5euu
ZuNVtBZek8cquavFhJVMxAj+5hpeK2Tcx0C6W2Ucgq0wdakFsHDiTZOx94EJwnZz
xTyoEJcoGrv5UCeCJe/LM6e2TN8ikF7u8B7o5Zci9uixN0Z5K8LcwmYvTkvyUpZw
i5EkVsEbrDkzoaUy836yEG8TshYQGXmHohU4zMzSbbX33+qvt9vm7Q6k6HKA4EPu
L1FUVD7CNDdFJyHDLrRy4oBdHAZhFREmbR902UhOotpX4VjnROcSxwi0jGYO5JfF
gJlXiiKfbrubyK8g1CEH+EK2uny7slpJcPiXFV4M0bXapJElXp13WHps/Le9HPRJ
5MFPoM//RGhc06olkwURHHfZHgA4pMXffEEFqFV3U68+nFgwe5BZI4FrcniOxkhe
VGepCa2VznDE8U+2o4ALBHJSuDdvu9z55GKnbhq90SAnUMYzzki3MM8h4LirDzOU
rSDr601ulc6nLOqQtkhtYFbGun2xe8eQcQuacBYUyVYIR+tBvUYoK1i3EPKkq9kW
CZXZ1VEDYM5sNFA9mfRe88qoOT0+slWqpY5tsss7K/Z2jU/2k8MrIz5BNtcLZjXG
R570CmkIyMgRPFH1AVQYO5VzJCSJGLBR3sWSL7vXeoOIL4DsjXWrlRDHJawhEKeb
/cexBdMvHPW4X7kIRY5K0OCIPFJ88OOXmNmIUhhBbI7hZotRmjpXVWNEEdy0RTk9
C+Z6m+B6NE4uP43rnN3IRGXxNr13ThMOYdq25lskXZ02DTzZa0rETNG0ipBv0/dB
0CCIuMf/NbyVEBu6aIni0faGgr11W02Ksf/LfIpAncyVZysMpCxI5QsRGUeIShxv
EcXcVSLkqU+e45f1t25+9W5QJKRe/dhUzEVAYkQrYTGcexquXwuyBGPF8JR9EG81
sn03I+pYy445mP/5vKdnJYP2DCXtpKlvPjNChWb4VBkMP8CG3rMY4IswQb0vAdBa
VNK5d6DMh0+jM2D4kNj5GNIbg20UikGyfxC6Pn58+9A5TpHDB+WDUBL7Af3XhoSN
cfaR+e/Dkas5wD9U4KpeBsZj9Jxxqvux+XJei5YnCAQhu3xTKpg3V55w6rZcL/np
u4r2i9gNjsfZIwUEStdSv42I60eY9AUvO+xtpcA908A/Y0nbUaJMsR8//t+jTal0
wSJXt/Z7ycTKqSEKn67GOEtzEMGlCYmrdWqzVTmV3wc67hYU7YcshaYxS42qglNl
HFrA6q5fidieFjmChwOfj7vn9EwxEWbzfYWwjEQVRg7DomJ88UOG+VISOfDrTJrX
lJVcgkz0VYABJmisRZ8vGnQeXBgbiWm6FEAV9zgsKUsJ54t7NV86ONExOLeWxHj1
0sIDs7e/Xw8G3AnN0JqfsxaC7PJ9+4ipH6pMsuHkwRk35ZxgUsKM32SGYeZhnk3j
uKsBeyhBLXs7sB6NlNUtKnU1WSErisSs3rAIK7L6oxpQZJV5CvT6EjuImJjoLdwY
WlqGvY966w6ExfpAmFB1Ch+e5J50t9s0/cuinKodT/bIDUjOVgIJ9A00AsXZNPOw
aruk/oASUnGxn5n87nxgA41xIkq9TfH4NlW7pU90qGxUs5oZA7gW6I9PhTSNSrwg
LHuvJmEunyt3vgsup57upnRSs6aYeu4dD32xxxG99uf3dDWNJ7gcOcfxFZX76Adc
CxzQUkE6sHbsI7ul11zRC3ykuI/SJn+p1FbLaCC3znep+WaI0g9Uw7PsZsvD+362
Mbyg/dV2xo7szWLyujCj6k5idaWHh049gsgJLQHNrNo1yzr01AWkoj98m7KX9bny
tKaO+Zyf5IqEa1nA0MjhFs4oGcFA0aB0dN67EH6D7VzcYvJqbfaK57vnlOFfuvRr
lF1ZJ8OSJR+4EP0Aiv/snAiC4BrBFGa9+lWK6cFdi9+oEyq2PwByu2jAzR5Jkmel
ctuMTDoa45NRqd+hJjsBqnWl4J6dxHmp4iaKVMPc1fK5hj0jC/jZe3dKo2V4EZWS
wut1fhRff4RFGMYYT5t/iaPqqHwzrMuZ5rNG+thOSc/Bg1pUiQfOuSJ+1I7MQ/WE
/tVdwg9fZq8K4F4n1VAYQyj2F1AlS/1Z71RjbO0xOiKCafJC3Nb1eUqV7hDMM7rk
bte0F2a7/lbbT0sTA2KAQC/JD/X0vvJM2SMuIRQOdolaKlG8ToDCm/qukJfGydKb
VJvzv1g3M0Aj/nua2Mg/7TNkHJufLBDc7ar25QIC3ANxYb/yECa9Vof3MVRu5M+A
XBesJ8PBQap7oYKddkaAjjT2GucD+Iz0i1pt3SB6bXvYHrh7lmx9HJBOFL/77BM2
SXN2MlAptJxHpEqiiu9m1odCWaVV9kANsGveqnAP/nCv5pV8y2CHJMbx/BUgejHK
5LukK0ErdVV0FFURhrf2vmiFABts+B0xzH911d8H74xrKZNXFEVeld9ulmjxveZh
/B2n+n1Qvqap/FpAjXl9BuOjL1eFnomdbr0sJ0h3Hi68RHjyaSBohcVAlh5j76AU
YRKq3zXX1TTWHExG+rmATgAwCIJoE99c2cshPWjEs5k=
`protect end_protected