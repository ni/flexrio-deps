`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15696 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
QVoh6/ZMejDNAJddTaZkN43b/0p314vzIUwVMFuDfSyDq9D5wSvlNAfw5fBgnd1d
xwiyVoLMtAzEAwvhT48OYb5ZdAGf+J6f56XvH95Z5jpd+IEqMwSrWe4p3UTpwuN5
2rwavKJH/1kozuhrcNzBSDbS/4EKFGdpdEsgFj+B9DfZHn3Ew/UJFDH+BAAzDZqf
8nG2CCktrM0E6PCygMKQDhzlOaFtGkDehrZS3UbYnsNZboXPvJmv8TWfKCLGPxAG
j2cvY8GYz13QYuksveU5wJv7DTQqx0ufVwttE6fD59T8iOpVyn4+13d7GjS+roY9
MOk8YS2j7N23ImFIaHujpat3IT3wLs3SLMiT5xeSe/Py01MN2DGKP6ebB02dWr0L
6OMk5oWHupNJVCLATKBvbBHAfOcA0ZVgJH0h1cWUG/hIFv+J4APDKT8yOoKmRUOj
J8mBznBwPQ1Ha53idMa5eRfbR/hUqVdyLNuTxRPZvtg8QKuG9O9KAYq0uwCcWKc1
yY+ngklt6rJPQCxmBQFtMjCycX7kb3IxG97gFnomTMsl5mhck2sGWAZMjIQIJF/f
NFf68dLGsOXyR3clcEyWuyn68Hg/Bv1OHqojyfgdfrc3lKPuqcA41B2hf2eQWJkI
SK0RzG4ZD1ll7+ZDie5fimRa6IeA+Bc8XO/Xa/5F2Fts6XTr7R7jBUftG5FVJ0h/
mqIyyzEs704ukCp4cSQIc+ZbbF8xkznox5smjvBM05048HNT2m1FPQJRVIOY+fUI
QGaxYdRUl6qTaqbvlQMZiCzrrbnomiwzKV0oTu4DtMM0O3VeHIWaoPIQCIkTy/R2
icEMA/r7m9uiQ0h29nvRHxQZ5jfy3LqLZqc4RWRXb8d2s63IxIehvg2HJCLW0GbW
pCsGMXU1JW/Cc29CSrPjII/B1VkPHWg6oAppiPDqIjvZDdceOW9CdTbJIG/3eAyK
d0DAQyHM3QdLJ2AwA9A13h1kkvrT8OIJ/UdSJvPrx1NOA74cndeP2RmveBfCAV+g
LDzXt9fJL4qTovgFCO4YhE0Y2Tixktxx7xAo9vTKbemgr8WRacXtlTGVFdeXRgVs
eZEoF7TX4X3djyVoTX6fC8YNw7goPU4+yx0URN7t2KlN6fEwscfPyQLntNJj1kXa
AwJ7gU1dZrPE3SrCIvOj+TsPqAeRN9/Ky/zl6iC1VtssXDtP7hTs2dNljd7mVgp/
MAXM9XXZS8HxBiWQnDWNibivvNj5GknOO3e0gSwr9m1cdN844W+9304fupIVBnRI
s0pIuhqX+r4Sz2GOSaV1XQ8FFXOl+ygusn9KYFWP/lMI8XMRfTROeL3pgkI5TVqs
LSPFeL2H/QuF61xzdSH+Fkp4g/gpHJqYy/ZObwr6JXHD5sEMTtEjTayLiDSqacb/
D061fO+N2zLNL3IUT43lIkDZSs4M01PnrVlfMrNgD73jEYa3LU88w/W3HT6/IXDR
I5inDOyFnm5rJt8yCKqGa82Z3latJiRg7+1uficQQZwnlvQomNtWeUFEQbMhSKyx
zroGDM8kbfWaLCEvsrRRLyAyjrDb7vOTJV3VVoOMGECsAcXOiaqHnJv0z4UvnwS4
g5Twn0cv3tzEtbqmpl1zlEN7bPOyOwqBd18doFwkKPeReFawDJs4ojvnSlooZcRy
AKidSgKsz7DTqI9R+OAad9JpfV4HHmv6bqn25wl65r9vqU57QXMexHvb6ltXjkZX
zkxfytnB++WO85qq0DD3L/8o8s4wpObW1CSh/mc6MxI8DZfziVxiBPoQdz7EWKGq
5AK4i8e1cUxC4hcu9SDhS/z3W/w/1W6rC/cuoAJToWVWE4K6OWSqw89apcUgV/7p
toe7hvV8PjfJOMFtsdd5F/g4eUYmW8f7b2+23uiraGHUSYQ0vfJxNQUsZycK7tcI
Oprr4VSCruyqSWE2N17zK7wnRjMeMt3c+s4LVqmZXhL4YCcOXWiF+Dg+q5OC5kdP
T7mX9YqKCHBGcFE5MaRZq73iFqNN1W1d7hO8ZS1y/185yTOQlm2IwOfDKA0+Tq8W
Zq8W0I2pvZRbgqBLU6jeTuM7r26gzrQn78BUOZOPa/vTwqdDWf2nX2Z78aD8kBd6
WQxCX7mwisedwpt3nHM9uwVv8L/6vq84xc8YC8cDkQvr4QH9RNseZppEjQdsgztM
y+g6f78YYwZ+OqTp0KB1tfKG+L4OPCj/D4P4hoOuKeMKdkdG7kMjwTjmfOfznNSg
zwcVfU3XOOswOq6c+h2b5DsHskRUv1HM/MZZjHGbcpZ6lmspTZNI3V93IMx9H2eF
RctpgkrX9y1x26x2GZrRrRQuc0eSRY9jMoSbe7Eda9ktsAVGfibggoSZmME8U0/n
haJfNx93gYuYHC6l5WlIO8DmRN90dBuLvCCm/j5S74AkOwb9zBQsQ6g1OMobKY1H
0XzdD8lJsXhe0Sf+Kakt9e5ve8IeAND9l6pwMbBY5vbO90XeXdgu2UwuUXAfqmlZ
LsySrz4eVOJHNr7m/bCHBzHFHi/aD9FUD/YCO+XuOkxAGVS0oCxtLq191fnVcT/K
kcuedchpvgtPTKccMUdSzhKWCGPvKUo8UYJfhw0eEOfcrKrlKEJsVSStlTtkbZmL
35lNH5oV45WLIaBxfJStG6JIaX0TBEsIel7oiwyVi7AmOEKMx4IMXs/WLZ1dHzd0
VxtwXcC/tsZFxgAQV43zPz+U19Xq9QtAixf2BGm8hO5idcB59LfyWCQWvtvupq3R
ce4SmtSRznywJkHoXJ5Pw3Zz0aH+DzrgJLQ6oCTkZeFShjhBywC6dBBpUuH/2f3i
S60BNn18jLEwX7UG26kPGcpqNCpVqx5fQlJQPBx1Vj3ZfoJotRFWIT1sZ8PZA05w
7ToJjmMmhdqkzj4xOY9DSottdCcAbVVcQZSygpEi4KZ3DZcBJHQtlyH1F1fu5QXk
GTkOHS6xdLGY1LT4R/eLGuMfEVrfehL34SvZOF211R3cEvC/2E0JQqhkzXhxee6w
rDmcQcfNPcbpsmkv5ict9LTCX5ZbZkNfpPhL3nO8NnGTadFiZ4d98s4pjtNdO+Uc
JclFqoGI3LDZuz5uFkkX0lv2H7Ifx94SJyAzknjMFf36OTBYgro3Im6DuZi/5UNk
Ct6k74cOgf26VPnJ+3RYEju+ekbunnp1UuPbeFtolQluIgfey/dc1pnNt/gDhb+r
xJAyLHG/dhKz67SwyrZqgpb4ljizCAwSMnIS707tQhhxbkpcBu4UwuT5M9zQ0iMu
zEr9nBHfaBgmuWpWrmgvnzOLSV5rBWqkfMqpfeenLCGSDzup0soamgEVzFhTngx7
l1o6Nqgv23BxjC76Pxe9iegiGJkPNJNU1mRVtmS5ESjyHwZxcpa8ken3L+Fcf9Ht
+dMI29RcXSnhdc5UZxwMXkQlx9eIqjKXAYcHydxEwSm/jliEKhjP0DoUYHrOGUJz
MmHh8kwWgxDzq56CWCQRIgL/8QvclIcfiylooB++qIf9GEnRNehj/gQQEo1o6IJw
lPcWdpAJTFYQtwineJUb9K+pnyc16JNike5f/c5nyWfRPqoe3u0kzo1hlJtgohcp
hoAmhChfUgvtGlrsvonojOITjiEq52L5QBfr1osmVUw+5J+/KkHZICKh8JN4ktPc
wVwKMxqGcHn9ebECkW6HGsyN97Z1PBksL4wPrbGgaPf7BVCzs9tlOZM1jwuc3Fhm
JLXKnzGF3RLtM6y9y2SpcoqnWRG/URLpgt2P1EVy9JWzD8om0hV8UhVJ4fCE+8u/
aRUJlrKzbUziZ+mWhHgkSenCu98uOKOb+DbfT4bp7ky9vD0zquUkVnndVa7ldIgi
CgVZ5wPJq+R2cZBrGJlZxQ3PYY2Aw2Z9wiHo1/ZufqkX0DjL+oWcrXdOhE5yYYaA
xBc4UETDI0X26n5E95me/WSnq5/LKvm6OHW3GrgUgolmOsbo3yw8wZKUHeQIWzEW
OaYTSabllJwAg1rSXTSZZvoJl2wu5U51Eyzvo9TapIWQlRG/b2xo2PtkxbQdwSHZ
8ER+httYYHahFh58mmLEuw8APGDN4ojPOLChwJBCbEd/trO1r0yFIXwvAlkgZVbm
6sK5B/oPN3t+LzrKf9Fpqb0BY4afRI5cwUo/OsN00vTjV1XPatSmHs+wtChg+yTT
YWhW9H+xWAAhqQCDrMdE6Ac1XeQREYj1i/LgrFZD5VGig4pSLotJA6T9pAh4LrG4
wSeFyL4UlN0zdpeHAp2XLWSuwA1JOoAxfzyxEc1cwin9ljk6RCtGOWnf4FGtdFAm
XGxuwvXuttfRTGaQhE98XP8FHcVCEF6Nq6DiZeWG9Ho84//pCv/8wSvoVQ76fPJ1
tOWku6erfZLBVtd7GTFCEn6tmxKWi8N1EWtm4KoLMAbStWGfkSEzUQReHZauwKnF
4ml0TCVB5GraD4b6dMG/PX4oqz42HhKGO1+daEpU5fco4LiP6iFTqr8NbHY7IZZE
7kspDuhRlu42wJa3ct8FK53LGUvjGj/pBc5S1VR9Z4u518rAhY+soV5ybe5gdyLu
byQNCr3WStMT2TvTUI3INhepiiJkg+wUmc6w0Ul7c4dGY/h13dB2k8K/Q+XG6K83
Yvp6sAW77oMvCsLH7+HKClCMpTgXTetXkvdbOAsM/8ENL3j/MMn3Vx/RkNYFf9/g
ylHLoNsaJXrAw8TjMeiA+7eIdwb8X2WHFmh1bcN/2HmlFIaescfM7law+3wWL8If
ZjCSHSYdcgqwjna251MneGY0OupCh2N9RnVpLNmiDqyNq4RFscsqaiYGBccYyEtT
ySCB4VDBYQ9GzaY89H7QghqsUj7ATUFJoVh8LhPvhMV9MqSsOChREiYhxil7+W3Z
jVOndCtoXib7l52v2XytUOn6BSR709exszjFkZdvD8CSIX1JfceHKMbWXPAqAt5+
HJJFH8IUgVKNiWWKyQqFJRKN5N/mp/ujU9EsWfCIu+LPBTZHx9OPsRhZbre7Ndfl
B7bwHgtJ+ImyqOUWxji3n6yZB4zecgCykhOoPjuNLx/9i6E6q9AC8IhwhK//lkAj
eyG+boOvlGec8FChAANuP+WpEDbhsbRxXwzYJxhOy0n3M5T4Fmtn/g4g+6xPOKVU
UWTXkkG2B23x6GxiMJxHXEbvvFIrj6NNYOPTYGJIpgP7oYiLNkCKMrJp/dwPd0nl
kf+UzP4FB0n5Wp/Rhxdt3oHrKn1p0R01OOoj0uPeVVfrddy5Rbf+aW0jPkxpAsCb
GrpPkOB4j+7ulJMb8Zf8gFxCOzt+5SQinDynBEWZ6NX8IRdJJCVzz3oUqaE6sWxo
3Xx0v0pUq493pWSA9ioKDMinAmHkiZbVuY/oN7KWCcej25wXAP1epzDgw8nqubAL
Z9W1xqqAuToSR/YuuHZwkD6DBODw2V6Gxw+e5ElopbudZpKfwHHJMM3UE1ev5QnW
Vq49Irc53OAPVtPQLkWZqxCGcEjMJpeS5pmKj677oXfroyVKUKCiQKPWFXxuYMSu
QdOyP/edF/waYEKXHaUK3kz51zjd8s19in5c02OA9yn6hOIkuUChvR1rW11SYz6F
USx119rWWWi3lTnnGjw4KJaQ7uiWub4lwfnuFmYQSYr9n1NUWY42Bn1tQxTCKhkW
V/3kbvvdweHsbVUhjqM1H5tXo3Y9fXWYpoX9AQkA+trZIrWZ5V6IasAEgFgJEww4
ms4WHzn6H0ic9QrLl98gUMaQAYAsHYZHf9ZaGUBb6zMcxP6wn54WsF9cUlFMAgJX
nACxcgkg8uUwNuKz8BeU4cCAiylNig5NjRImPh1gIKafIjXA+KMoSOIFPz2LNv7J
8g0PoPu+I4yF2WRM10yTQTYusKxhV+Rio2iGA7n2/CUzxBgkVcIIVnTazmwhkctQ
POAxJEdL2Zw/MkZDtq1l6aZOfpySUAzYzCEEJF9Sevu+DA85248Y7WIi6oDzCGvj
cldPNWtMSHZDC0Qjy/l/aAtFVoCmXcqyoviRpqJx8tWstzplFuIiCywueJ4y4+ap
d8AsINMsR2hTD+3ak4laoq/imFLYNzIyYvi3m1fnqeJ5z8YRvhHQ6RDWbmNNZPiW
K8x5FgmiisZlJesEt3gdyozSfg2uN+NC8fOL41vr4NlroP/yiC8e1vrt6X6gUnuK
pcd9eQx3R516MzuOKW9uOIYcamboUOQ9OmIe4c7r4k11tTuorYz2ddY51p3gxtcB
uCZPRCSmWaAbMO5JQtVp4PGyWkwzm7V/hte5GdpVUxZ15sxiIIxvt2G4NnSloShB
YVDPkoR7XENVblwaohek5wkSFUmmL0srHY12+FH9Nsq8nVeu2NtHUaZor/5Qjv6K
qiJ3KgihlJWFP+P/1+xSQVE/mdNu8+HoAzGqcCgQV8iphHS9a3zQOoqjftUIpZlR
ZtRRd4YFoPgpKgXTihVyegWP7/b7oDBAHpiGfogZOv4nt4/fcTpP1n8fPiXqCNmc
HmHGCr6nBXDTqtcNGtI6GoCQFWCy8bNNf8dCRkI8B2G+WunaBIA4pe6NFtj5V/R1
PjQU25TECnAe7iM1GU4XG/5Z0UEUvzUFXMgtFWJt2hsMVzL2Pu+wLeYhsdVIRqjF
JLKI/6L24KhJGItpwDYmJB9mHlwOt2EdfDdXx9Ztt87NkuFKApBc2yQkdAPEQxQe
wruG27wS0vsvRq7kUOJHiAaFhPvIOBabTuHXtloxmFmE0Japg1mRi5xW8M60ClPV
y1XocCJ+WmLf9huRolaPFo3yEOC4Bztk3v9FoW85UGP0dMSu77tkyxmiiUIQPtjo
pB68s2F3edFdFh9572rdghNjSZctXEMQhGpBJPEZhXAum5a/5PTKe3NnTOFkh1Yb
jK3N+MS85aJPcnnG4xBTt88gge1lz2QpU806u/Vht8cBjeAe7tUK5GMlpdSomHD8
m9aj+xvy0nqzwLhtNMU8N5QF72SM11zBqhlFZEoYusYiMDBEtFxMGNAal7FJM11o
Wq3Lwu0xWIxWXKaFVSwTMbWRMuTNZmeNIU16OySoyxlICeH1Q3c7nUXUa9EuN8UB
Ef51BnqhjOSK+KCN2/tsoGpIhQz5e6HyFljYzfTfxEo5iHVPAsRUIjHLcxN7I5nI
FuMFMtg4RuAWBnmJsotvvuv72tQC2DHSweclyDvgGtjwZzzviutnhowrVVHJ3b50
r4C8w6Nkvk2tJetlaZyGykT3dAWKIx+G3YR7R91Uer0eBz4WogItLNy51dlEzHVX
h4KBXhljrO1+ooYZIZBeiai2dcxywJMm77+3jeyQ50oYZSPBMkmGlSAGdBAWtgKE
H7UzLWzAlx3eNsSP/6c7ru1PryGGfqwPk9N40r84Ipz2DHzpuaj5Fqk2LxLXPmuD
A149XCx1xoBiHocm2BB5RIrHcukkvTwQcqgSN4/JGsHfHuxFHlKCtBWInyONQe+n
qp5I69Ei6u5yHURdXUCtKEbxWwfEgHcJ03Hp2c4zUxZ24rbcDpL47vWuhSPQiCuh
LzjeipLdm1ikSMSRxAYMgt9MKuljkQoqS1Is+FqlOSegxqL8jWD0LekuFCTdBf7Y
S8NOpQ0hJdr56gbJ7kPlEpiYFEEnFdDuTl/l842BIoEfP3l0kz67vYhOyBQIxGcN
hdzfwnw6WuNugKGwMbL2Uh3+I2Hnl9fWVAYzymBp818j/wtgYbXCSyhUm55J4yEU
nEtV8AVuXsZXhrIKDm6nYCPd1Hp+R8JVWBHow4LQqkGM3unLG7ghc+5dHzrZmy9D
9d7Tt+uKDbZ+yf7dDVXy5s8cAph2h+kcAbBvS9ylmPmDq/zXdgN1CYcIUpIQvZIb
vLIguu6ZFt1rkRGfwd4FIHLcfvWlp7ZCrbaM0DD+7MzF5Uv734IEuPuet0zK7gBX
iCAA64MqoKtEc0jE1s0fXpDbv3xq+DBFV/B3GZ+i4Uy6kUqOOT1rtLB0QxcUV+Rt
YCJJzO9XIv7cGXapvmh7B59ezNZwQdTTzeBObjgCGxaMeGoEO+ZoYkHsQpOQ+UGP
jxmuTTylqJNXfOCPZzbTWMr45fTmsZTq3wOI2xa2cJQNJOwSK8BCY/Yzhs88kHTZ
60MR5Te6snYC7kmL4Q/JQbSUsvf9v+FQFEC13rXbbA4DsFscZ1NnGFJQlZrMgzxm
kj2F8lAWYckTr+JFnYmresq/iRp6laAahOyZLtngOrmxsQcNkc6VjYQIJ1OZTdef
O/Zg4WXkM+2BQpCpFu5bFOSfXMI5NPzMTmofwIYxi8EBBXe43J5p9TyuxDOMUgWJ
KA6oiO1RymBxJy0bWtUaLrUzqOSNk6VgJGDee+zRRGXmaKxxVZZLGGyBCs7wGLTO
fJFuNVRk8zI6yWdg7dUKqM44YA8S66gVb9Hixx15nrJdhrxv5C7ZVwSESpDLFGpV
jLCudaBSb29UXJYF3HUTY0lCxIv2wAH2o8g4gvpSWCScEX3nNsKx0469Phq1x/2P
yyh/5Q8CQm0eAq2L5QggYX7mXcDWXBRt9W+I/oE6mrOtnBvGBmXdyFV+hrBv8T2r
ODiCp7ywMkc0hPFwewzsybyRVW0WCPeZN3rHYBBmq5ZH62a2cdNRIomBjnSSHIzr
ukRNLMX820rfOpJWGSj4ZSAYGeWVLHkJq2i6kDhmpXtMptb00TpMalXRIq+rNUbM
fqf0ye3WuI90Qv1LQVeyh5DQUR85pCLv++pdsWAy6ABGS+yjGMVgE0F/iAqrJXF1
nFloDlpsl5ZNKMDwQekuJBWvNWFaRilxGn+l9EapEmS9Qa5bEVYCWv/6Pcx1w4bV
1WZb9lxsDUxorsonA5nEfuErXthfpfYTYvR5QUjKybV8mbYj3FiCxLloL87tx0Yt
76m4Za7agLrd2TffefugxFd2nHB6EkxRGtYx+w92NuFydnt1rNIWkz2TQg2wZSja
QKmv3WRxajOhwE9Wx6Q2jlLVDC3O24RfgaroNHFl+EXwjgTof+wF56ssZKY4ZYCa
yRaAI/CGtnUYZSWjC6xcGS4fSadUqvVZeE7XFm6x6e/SJggsBDPmHFtz2KVojqBR
xTjEv5e/4uP+plhwLqdToGF5ayL7DDlh9pVHJvUDgNGLej/xh8iq8DV/SJCOo2Fo
6OJ5YpNz6++aP9k0389o42dnwHawgGMDCLwFbcsfpFXyB6pkermXhWzjlyxhDw58
/pYX5aOFkQmrcdAFZ05G4hRTmSz3pCrXAIXaj0SkaBe0INufBUzZzJa6SL/RN1vR
prTB2LniIhhpN6xmkBuvR37Ao8OD1oT8emY55bc6Qxl0AXOwMV9u1WBrpRwTRslV
kht5e045c7HzKn5zW1ot5px1iCJlGC7N5324wUTFxvUgOp08DVwZN1zwE+uwH+VJ
/GrZnM1ncFSTMRzVMACM3SPzLTh0ZxeLB3OuBflN3RNIvRXZ1SJGgEqZeHDGbO7H
EQPccV6Q9Vr3F3qkXcgkrPgkK/2p7pnA62sgjvmmiWxvHeqiuFIgUQh2OGm2r+5Z
nDTjcURbgneNZMi6ejB7Q4NHDC/bjSFUaQhSl6Ku7Kkz8Bp2Gw/yEhGKnbLyPVAW
TIRe66TLufDvuZsk6DxCvjJWAmOlYPhxpMFVy22OXZZqWqH7gsLs7eIA8Btk0Njr
N1B8curZKLke8jIRlNaYdHfNGKd+TUaSPQbILgmEftJe4JmrXSrGbFJsEA2+3tc6
Z0IXa16y0sHiGxQLmChz1b1On6s+e3fltKm6JF5OT2u9Jw1loQROfZ3Ia+qCc6xf
LTuWcZgnl6xtfWZp7Ttalq/qF7d3FGdGBT6+4pRmzTPVRXDVkJLBfdTPkDzE4Nsw
imym4WJmngZXiIwvQZ/0AWallXKaCW/u2hIvZWOg8zdEKTzu19iP0Q0pgEr9jOJ2
E7/v5iLhIx4QMm9CtjiZeccsyNjs1RnJ6oR+jkYbW49Nthuy1N1Al1DkVtasq1Sp
riDyus0TwqacsWffFz8umiJe6zez1AmoHR3nUs8VWPk+YaMmpdKo4huQj2E9pbWq
oj41PkI1pR16kQcxtq8ncSjEu7m603oAGapMDGtdML61334BipvHCYxrN/KABceN
QdUaqukq+RXgR5b471zgHkr9jDFN/IV0iPAIhqeBPJD4OYy7pUvKvLitSU1PnKjV
6Vq1M5PIvJH68FOMKnSl4FhkIoI1psWxLiavY6eiDeITzqFFZdTFwgIooFJrO/yP
yGxXvShH9RQSzQQI1A7DtNsvQHvLBiS8lcGqCgHji+aq/OBr5sK1Azmk8LVkGZ+z
nS89PcKfti0SeWGOj/504YgGiTSprH5k8/FzUdk2wCNh4IphAXD1fRiUqtXWoc5A
Pj9KTv0Kx+G+bWoWl0hcPR2FNCA3JH41IxHbSx/Tr6bTxIbJiBHN4JVfWwCWjf8i
3nO+zoMX53OOyn0gdBpvO2kRNqd9xB7Pegtgq0wZD6on7Lb3w0CkK+hMBCaEDQzT
wBVVB6/6szYnp0saQl1xD0rhuANiDWLG4PgpnGRlyXey7Lzno4wfMOhFO4DWSYtN
hYmMssRrzHife7bxk6xsawBvqrlSuY36fpkDLO9/+rtJjxm3PtF9cgNkTKuv6Ce/
HUjuIPpid3NFWpfLXc2TKu+3oeakuf4GpnMHcKxtjJtF3Q0sJmRaW52f/YtzVpUS
p4I3wz0uCS5TFt18iefgpaJYbo29Y4MMbuIHLsglecR6QV7FAN3FSP9E2iBbkUgs
AaCW6BevGrYsnxTH5fAuJeW3/wCHWZmMCDAeMOyRm28bcuLVflVVaXRzxpA0782Y
aqWPWnmc4QDMJdIBs3n+qzkaWVwsI1d6R2c1jCvvHzcud1j8oUqGsFa7xu9wcVxy
GzNqD5a8jTP1C0QAD3g4WvE/OlMFMELOCZ6lfrL+xHA2ze0yRnPg58oViQCa86KR
dMi5skZ2CVolJdg/oEewDIfe5Ne2ovO/RA1C0xYVNl1AfATQegY9xjKfaaZPZ4MU
6Gf10qm4odElUL+uEPOgbz7CuMxY2afCCUiSy8TesUHXsePyPsCYEE3zOg+69uVg
v98dWzFP7/VbjD2wvcn3a0Rbka/7lYHa0w4cnXPkf19zzrRaFIlRPs0b4djIuNKt
ycUpSuj1ztYP+ihBKCeK2wStH98YK6OldECsdi2FqMCIoRs8caiYR5kj0gGw/QKH
qZqr/9q5FJ837az/+NgjTvewTcSqUXiE2L/BfsWhVn1B/8KakSitvlOaTeEZ5JMF
H2/gMVQ10m6kWdMiyJrw4C+EfPr/rhCTMM6rRA1PF6qYEPkilT5fU02GqrkJZhIU
0zTs3cmiqQBIQDoUGYmHU7W+d0/V3DdoBX3h8O1yJl0s7Uqti9PVbNFSUo10jyaO
iZC9ciQyfT1CEaiaSPtIM27B9z6qeMnSEcJ04Ujmgu22uT19Sex9vb00ymfdHFjd
k1boBK04RBpp0mRqj0c6GIWY4xiLC00IKvmRHdApnvYUQavBmG9B8cGZ/G2sZCxp
YV+2jjj3QWPzxZ6vX9nIwmjrekOIcZ+52osjU6YWNhsITwmp05fZzh0wa908aeiR
9lqGYQT6IzweXRiA95ziTXa05fRnnYKSwhEbO10PBGjrOflvbFo5KvNmUmIYNK7u
+NaNc4j/L34vNPxoxxea083YHDoCe1tli2a8Ye/RXV20iLPTbhZz9j1I6Q/2S0WQ
OoRboGoGqToFXNj1L8opvxaYdbXZmSmtLFT9P6uDlcY5A/ffWx6a12u42oQaVBmV
t6Usd3LX4YJ8jI1tLzZHO1Z2oyiO4aHJvgHi/hUbZqpVjpi1zzv2boc2RjAPow3I
AsmiAtT3trGHGjkR0/Hz+a+fxwfE6VwRWgNNnYe5Cj3d3CuH/xBFQeKU2qZvAHFR
eT2cq9vVS4uiXjm2lWbBtD4VTjEjyOqWkIHq74PSiNJf+V2tL87hJHvljpn7X4Z3
cNhMj3RE0yhMLX+OPkLlytZA4ghfWXXvoPBZ7dSt+gIKpZ+voYVxrjmEiiTtPPev
VcW4i3Xx5HtAIoRQbZJLkk6Ixo5k6u5v2SqdUEz2+GmY4N2lEmUwi4zJcNCL78RC
8ESbG9QJs4tPD/AtYHCPaIP1Xt1Iug6rwt7MJk7fVnFvWji2gTViYDa0b6Ez8AiT
uSUPtkOeNtS/BzfEmdb9FXi1ch3VVVlu7UUd7mGSJ17rrqTpqMm2lhUP/K6OumIf
wtfFDmz7aA0j5RlEZQUhB4GgGPTWrYXNpc30Z4IihBguDUz6w3F+kbyxhpiexwQV
rNe2WT7TWWEIcHFKYGp4bTg9wTYE72OqRWw9ZgAHJVTO4vIpOM/LX/rEHvylNRAC
e2Rtz+vrCZHqqzJN68cWIcRxiANC0IS/UR3/jb07WuOYX47UVa7vMIp4uSA6hnx0
J5EGpUeN11pnysCxEftpf9z1oTqXePBSlpe/Tj0rAlIPtBCTQiKwZ0dLo30rbQoX
Mx7db3SYtEyLl36CwpE0AJB2ki/iza02q1Ob9z8wh6Y9rPQVyJSh53slkVE/Mqlo
ZNJ+6lGWE4JyVT1mcyDsbzkk7sIyNg9LWp8Cp9TPIAbdHycQSHVkuyZ4XNw7pdhz
qJT4toVW0RJrypaxaC1WD6C6yvWS3LKH0kImbaePqIdp5FC04SbOT/yVwoGAwHJ2
d0Av3+OkaPONiYaAAm2P15613YSfVpzXQ8Wdga/5JRs3XWnm5vw6i4o+vKcrbBbS
oP1PmdzybuPQztE9n6qG8JCQogBjS8aBQ9Jw8CMXxd+PbSFgP+LKtwzu6lhepDjO
Cqz5U2gprTVfd+f2ZqRDH1nT+TzUzTe2UXBVAK6a7b0RHa2V1CsoojFg+iRgkzJO
9WNvlIWK59BZKJQyrEz1TGvr/90yXJdLwnF7+VpoefdVbTVMlR1MMa4nWr50tM/q
Y/fDqCLQe9SaCHdpW9yl5w8oKVDts48JG11aRz3y8dU+yw73dvXFLghT+Rg+zv3e
ovQqCHn71yzeKjeyZ9kIkhD/z1hUNUWgSMsibN7Klpeh9JF6Y+tAg4MsdKmQ7eVZ
cqjviRlO61dtlpviR4jnJDpzemnUfyZU9fdU7qGFTJLcgUZIfJY7kAN9Pe8yrb7i
XF+o4cLWXqCUDVrVsXYqpQa++1chZpEku2ivsKfovd4oN16vEIZLMvm4RQyzSCIg
HlpWkzdo4eciNSc2Bpg9jtn3D4zfI1gzzMWsjQXG+h8BxOou3AllgXE2B4DM3mnY
eQrnFrheBiZj5znLPCpl5ZFNb8yzD0TnjdtrXadJf0jjzztt2rfueCPKgTlF7zil
51dibjXcC6CHEMtftKfBtEUtft0VJcsXyfe8aYqIr2xFdTW/4pXfNsOi8yA43NOw
U865oz5GezwHX0hF23AJn+pL4HfNcmSC72ZZrjLW25DyE+cdlelUYJLWcQ9oJfan
L+PGSZyJICLKjtRDauozgcYjAx6B4gIE8Ij6SukoJJyCCTASyt+jASWkytWZnFEj
+QAMJG6Vz0qIF9fot6aHE26XhGNe3ylQaA2j1xQcoTX+ti4mpg/ogXccLBIvNW2O
kIokNOSxBSkUkfRQmBYPg3NLsRlTB3A4N2xB6G64rySWZQ0SeE1TgRr47J+0ddix
pd3MHapzi7N/O+q/sahbgk76Doq/SIlOO4h1yVw2a5hGIZM2lBkcLiLT42q4oJNs
lIk8Tfguq+MTWkmKnaNE7DSzvIgRbxntF//KfNqQBdd0XOv1TRQBXxT2YdeSEYRl
g9NxqXNFtfBzfMj7G7gge2aozbYT/ojLlOkunQUY5IkdudMQK/lHofNosZiaK8y+
YvRtULqjYbKeiCaLOre8akyG0rWmskp3iPKtXK+Hr8Nf9PGMgqrbeBqtWZSz+Bfp
jyPKtR9fDsRDJIQMcsfEvvdpWHkiexL+EF6VuObNNw5R+xS4gT7YZWqyc3iy23Dl
msuJS8NldWc+EaoQeT/KkvRJDgKeRf9Wcy0hlJiXICHNgPvahm0SNaTYrSMuLZZ5
SvHQX0MQuhwqbIqKqkPu7Igx14I+TMtR3KzOcx1dEWcku+VHDSu9vEd4AcoUGuEE
rvb+7At042p4YhCYUTT093c6AIhxMOqiCidUBIZquGjVe3TmXe4JkW857xjEYyaP
4ngF2+479kAe3zmUohY+Qg+HnYKGPgWYJUjwPTDl/RWvhvxd0NfAO5sEXxLjmUN5
iZhlMsxuQl/tpFM+hhroljIB1ffvnr/HxXD1SbvZg3uybbCkfr6lBndXqPEM21Zb
NMwyqq2UKhz9VnRGXsF0qgg4bsI1RokcbJg3J5CzZpva2UifN/zYIdLereNRaP/1
GhGW8onNZNPcC8aCHlYyeMlI/kOObHir3qawp/Yu0aRTs68Pgwj++5gq03qcDavr
wqoYBPGTY0SHqIV3bzggTvlx9tWV3xOSTL251Doimq/zXR4adUVBEwSTn/H8H/6r
8xKA0pHEpyQ8+p/XYFkADI39QPjr5uDLCRTZlaAdju3Z89ptu4TZyW2htiR/G77d
SJ82Q2KT//5I2M8db9PgYB7mhjyUjQK2wBIaAapPAA70Li4/P0wuEScR67xleveJ
uDyyAhyPJ9RlF/ybO7+4B9ApZu+uu1zPwPlVelPrbZ+MX7nSaAvBkm5pGKEkpKDm
63pJiWxosMbLs1EJ5MR2OQxZtNUl9MDO1rZwiCanvKJYiRRE311mur4xETQW22zw
xm7hsfJu8M3VX2qqu3Q+MM/auFmdmqqejRbxXTxazK4TxxyLGnhtZ2d8N9tjgzeD
2rmkFTBIvywvpwHAGKBezcxBGlW3nt4UdEvtmxd+5yAbhqVeUJ7KbJWcE6XJZkHo
ewShNcdVLAS/TA1Hm79quMcQ49w4jFc/pcoAlh3il7scrN1R3e/W6veiiTAkC+a5
VEYQ36uKPPcohlJJl/se9WW4K3bJeG4lTeFFEjBWEV/NeC+xwHFsCGmxhHz3Uanx
l7pmhcDMYPyQSXhjoXKDwEG48Y3fncH3nFTEhKwgHZ0MEdfOwF+oaJp2AoPAcnMB
k/guR5I81BbwWenSsR3yGby3to+wl3A1AQt+TiWmVIz8Q5rbGbh2/MkF38Actcn4
TwzbWT7smE0MOnWaYfhc5/QNi7/GAMB5ajWSnmVh87SXDUxV6JcGcVFOl6MeqsHP
KHC5qLNbZDdP+lax+xNmhD/P1ZcnNGDiySioTuzPT1D2bMa/9N1L2D2QZnPBxisQ
yT99eqNCTd7n1si8RaHh+sxCamMG3mgV5PaHoPAlFRSRNGvpmW1PvM1EjD4gzDY9
spveDr2zdco2n/qp/1GdIoZ6cEIQ0qUemkFmAAsr+C36HVPpWNHDet5KQHQyFWck
RfTYfhJI5m5enKd4lWwPgMgPs4dlwQB6L4xc0snOVdmpd3cCCoDyooY+3Nyd05Dw
DHHg19Y2F5qQh0A8nwLDlmFHktDDLodkGDwyK4dNfxgYp0TQnXTVO0QxsHufH9wD
1ragrnGKteVPoDLJlyRBpwPoeee+X91welHe0NpQNXADFuAn+BD8Utgnv1pL6pQA
Gh2hY6L2NcmLc7P9SvwjZIwVBH8Em0UxfJngJqfGZW2kXvHjTvnvzf/E9WNjA/9E
Nu6MYcG8zOHpF/2IVtQYCVgKQ0Y+6OTTUpbse7J+YJU26iFQlZZY52kSR//LnnPJ
odorQ93N1Jxr7efnzfaJYDMs5FnzCq3186+Oct+EjvAM6TrqapLeG1vFWIpTv7z0
j88ZCRrCDW/ZjIDQV3UOtdNq82EFmJFxm52AGlLa/Y1Kprbx6umzsvZ283fB6CK3
KCAZ1BBgGHOolqs+ppIL/SJ5rnj6Gn1r5X6Cntw0PwYSMlN77r7BRB4ltt6ssT/S
/m0GoANmSmMWUwXBMquD7VPB8P8X7YvpARkU/Hmg/6u+u5FOTn902TwaoR5zmzbP
oFrG1riaZfnL/qHAq1euBTfVOFx5p/gCmKOoECHrIT1yb3LjIgEqYof55lMP3al0
oBFyCmy1yAq5uE6GINikG4A5989k61oykp42AsDho8Kx21eG3bw5Oa6ftEHfYlTP
bjl/NoQzlUHEhVPH5GzaA+WYcCiE+AzUdjHNtDQQk4iub23VWKvAN3CPouCqKKSR
nORSo0KeQxi7u0dgob2sRFss1WEssK7cd0UTTYjmB2RFJ1/zMPEFpl9As7tsQJLn
HH4WTkONRYyLG4ui7sF2f7HZSvFRkOnEyGlM9I9GtVwuiSOESEdJ2swPbgxoHg3d
y7rs9F0THDs6TPHFBh8Sf1MPfDsf+ZSznG12JtsO5gqHCquaOATjU0A2CgpoQ3Io
01/z2AFiiGjLJAIIdYJ0RBPPjRHeBSHcMNQxNNLVGNdUGIDgG6abmoPqAtm9PLbH
rYJRMFuRxyjCJlDo8g96DGe4vJlP3GA87MWrfEbz0kWmViNrAz4S4cKxph1jeWDU
c8eAGEvYsPDSpMiH5nY1RfBUI1diwTE3/ybnXmXEpXcmLulTreoBSYAtr6bU9ary
9Bq69Ph2u3i+d1AMijg4T5kSAqdScNuCB0m7wnWCEbGQljsRqTLYb0L7lUMMwj6X
38ASKoAuvwrL49P6PRia2IAEt5c3plE8XSXs9iF5b5Vvcf/OIT+zhFSh0RuYZYLD
4hp+luAt8rIUzxvIB1AA2gU6XA3xvEEgl02k3Q9gQQoQ48l+0jfIJlEFSmW1krYm
cI3muPqbwtCpt3VCjUZurakox0j+M3yqT0ZROZGqHsluxfgQe1sEAQF8F7hVLiOv
bUjggu/F+0DPYeIZrCk8t3Z4lirz33JwBS08H+Xqi4UJZy49g4wLdSyQt/YxdDbY
uwXPTm278rOpi4M9eZShODPIo99XaHZ7tNgaoM+P1d5mYs8rUHFra7QRRntxFF90
7gqKLvNslAsHKK2bPTjpr8mymVzoDp64jrZXhtLego1+XoBcLFRHTs1d7n848kTR
v/U1JtwmDg6ggXbfeCncsf7TCwUFz3FV/BjQ5vo7HECayJ5J0j7On5/X9xeXyjO0
TiMmmwHHi59LeG4srvWpZkoESo1FiqYEAya5qUmbtMPRFqEQS2xIPm4ji+jcjWtM
qJrwiNeFddmRiTnO7VypAqoHJR3Nu4jsEcQXrOogK/0WpDRunjtqvh4+VTtaIV4J
YJolWKi275LxD1gHdT76+koVfTJeSgKTSmF65pwl5FPNc19G3bDl2CYqJLInTjpS
cZzZEV00PlGeXfXuzwc6Zyo9YQUbiRInXsbMFl8TKEJQR+SMPgk9xSaTXqpUeFok
USE3W9mSsOapQn+PqWdySPoyQ/vKvaZh8GGAVFgADvtye/VwMnGQL6Udz9zlideh
ymJYwYadWCAh+J8lynK+4tb2ZKQ1KgJFSnqs0TLf0zsTHZTMedmE6mmalbY2kL4b
06frow8Ui9uvNYSrrjeAB1wQs5cKBw/VmHxQLuYG6ZEO08DrbRRkocuctaXI8RSu
bVIkogjyNsSVv4j22g6sUtEUMDobGL1XG0z2hTo1dIfuKnpSqKbye+G8o9LmDndG
aT24pNeuuXfN3L/dKYrGRcDFddT/gc7J+bmK10qc1r+aVMh5dMF7UOTEBo4sVwYz
SQdDVSJGblc8TfHtuwTWckr/Yi8FK/KbhfzdId9lur3m3kg1m6Tr4WHUkT2AV/Oi
mZfCqVY8K4O6ul7YfsriPrP6A466l/LmiR+sl+2v5lq/VmRPYkz4BjsJUHSYePnk
s2LoVieGe6xXV+r0aI/AsLqi+QLjZrCrzZYk5y/ipvzvtvXgJ8el1f7c3/fRBzfl
rbL4dm/KhQ4WT7ZaBmM4xbmiYEu2LlAzkEbxjAFKjf2x0zZ3ILEWwpm+Sxt5vF2r
5CG6CKMP4ZEf89IkMDpeWaiTWY4HU0+2Lb2SfEwJZt/2ccZAzRkWys6GAT/XfnW7
IogKJMJuzDO8iKxbceCuqXf9E7YZeWgCXoki0PGZ/xfJFBdU8+XZ4KR0GxchwUN+
hk3Wz0Bbf4e8aFFjNv444VcDpEnZPoz58z4B/8S0pEoNaKrYFPT3jcMYYfSPPSqB
3xk/iMeMUyn+N7N8FHuqwQTAnt0SUSeX5+hx3Ky73fAOKINOJUzK+stYnhFMzVCe
VeFBvRPn8CdYctAS+TGR3EZJV+LA3RqCUbfAsneXKcIFz0w6ALxXR1RfvwX+AWau
k0de8TWC6pJ/m9xqeE37Ih9LfI3g63FhnjaTpUw+3560EP8cSp0Ct2rsY7OREeyW
0oPicsBYQwlmFrUCSYANMej/V59zfjsbUAi2nXDRnFR+6SAIvBgkpI8PkXFH3xqb
4rIxUZD6DYQx7g+54Ks5LeLJ9dYYBkQeDGqWSQOsbg/gI52feRLQb8JxWLMa4tyz
KN9fZXNXLK0wOHMDifb1Y5m6IExeDNtIs8qWH3f6C/3q5bdwT1Nj9Hz9JbY0+RH2
lNyr9WCc3yY5+eoQHbYTCrBAN1ULci03ZwG9dnSB0e3pEQgMu9pwyQrGJaYQYmHG
OvIDxsDuXfE7J8PzlMhCByphChEZvcmjepqrH4ZheOiv6FeSXBOCjzyQdUWxbbpE
8UNuRut2+xkmMSY/V33GSKbBkCI6LN9BbcsWLQlUxuofr3aTecH9uV26DdgYlZ9c
iH1jCMhGR/ZbbXtGkV5eZQCjFL+ouW1CRrTxw9Y1MsUMEKYR78HbL+FiIlg9U/ly
TdpP9ZZ/V5GSV1Ud+gTI5jvqZhSi9SjmTaiElJ/PcMIRGaw2GPijExnTHhPLTRol
6DPBA6EY5bAsV7mMqYUSII3TwIah4qOC7+Kqyb/dzLDjdN+ejhisXH+n3vUPdu/1
21BBB+8X19VeVUKgY+yLKpAgHFSdL36FJhLOvlNYLAMxXCteYKSHMQRMRHSk4XW8
BGH6OkAK7hwcIgPPRsggllhuzx/Qk1mIpr++UmfrlE9k74GunjYF3dJopmzzEL3e
q4etJNWC0+aTkOOtRVeWqakcyljyZ9DamFm3xiNECEpLz3KBLpEDDVOXJ8+VVC6D
av3wRguB6LE7nPYVpDQqxw+69xLjGngnxIAxuSAbICEfR5DnlHWYMFuYf7oMl6QY
e8nH+kYNMhuUi6vjvD75TsMQl27PIvW5n1JxznEqZwXk4i0jP7JxEdwukH/lgjcu
p1r+K0q+c+EDUKws8KCz7uC4kM2Zd59R5lbwe14Zp4iX39AKG0BbPKN9vp+0avN0
YooKDJzLMhQ84X2xP+Cfx4MuLm8y0XctaB7bCL8Vl/9hIFz64sFNB96ZR9zmn+fH
zW9uG7ui/ypCYLhEDcUQkd0BCoD4yxVfD15G178m2xvzhg2YOMXBhLDXWb1gbUUC
C3ht21tUTCFtVxZgDs8bhceOQe6knjDHZGqPQ6T4Ub0JTgepYlNLyj6OBHRkRi2N
K6HJPNZV5/nSVO4yMwW/b+fHcuwFSR5LtdcCvYRira80v7FGavOJLYmvITspKeLn
WuaT8zV04kQJsixfIWb9IJ3kTmSM0BdLqzkb3ZanmJu+EJ+VjDAfTiI3KTmuvxw+
KswJ2bI7Qs+N95Sv3GnZewP91xO7JvxYkhu/dvI7xNxpF6yZWuXqfPjcShGiZNJI
78sGdNNd4wT1J3mcKQNQy7QG/3EVVuVJ1EO3xYm2vDxyubuAaYx+43AAGGPvoK2I
aWfr0eYIKUmzn4SzsibwZFsKiPn+uSpfgE0Mz1YGBW2S2U4OJldT0k3QirVuIlso
OrVn6CVk5WrNAX3QQTlUztD0FTFd0TeNVMmsKKVkw+XKAuk9kPsXbjfJjv9Tfx8S
g807P4I6kJLyGYS2gYxIEvSG79DcN237Sf6R3Zbtw2RUGEcgKPHBBJaRbWxb9Sqn
AAOhZAcwoYOjRPGOKnbcHVRRZx5fgTgWqi0nAjVQmDR1WLyDirEWuvci9XAUM46d
0RxzR3mhZ+z/4MFFMSg1A7RcK1KYaFP98recJwyq5DHR5wTR5ITeiUtre+GSBlwI
VnGt/xryVH+2DkJWMlvFanuGLYy0v5whiIZ/hptyX1Eljqf8o7LU/bQNQC7e7H+G
DE4XLbv64NNur5ds+UKK3MXeKib7CHV0+pWr3obX5eH0ofXZf7luwN58s6D9AjYS
AM+KW5bEOFS57nmpwORzzdkjycmcy5jqYk3DRPF0i4CAGhMaI5hw39K290D3V63x
Y1q3Tbml9l1Gm6g7N8FBXtEZf+vaxoTC1E9+2eDNP5sdI0pyUgoWAaMw3xMLgZTf
efjD00lRe3W1Nm8v80YshXpslKBrKdNtkR0BMjSMt0PZ6GVw2Z59OycdrySx3x2l
E6Ozw35fs9DJgVQ5ljvWX1cZTylt84nvuVOmbu3aT1lIcmbR9gn/eiXZ1H+v1MIp
S7Dij/+5Ddo4YsHCOp6y3qZ5fKx5GGhlJYo+CRFmxocX1dfIff+kW6eddzTDDgBV
fgKGmoVreTYw7ev5LXAYaAww6lvKVPZ8LD76iG2CH7XHBYed01Z/cjBgQrIJ4r33
JK1guX/KTCgLygIhyFzcPdGr/ZpBLaNlmV670Yq3wtBckDgcaS7/TnTM161H3Ls9
nWuCuXUGeWL6DFf3nMKasUCcfuCsvnx9XqrpA28tToh76TS9cYGanWw6DdOdSAxp
3qLT+rdndif5ZIVHrlgyNAxlGAmRhvtJ7eZ3662wLl+Cma6AAS2V+hJ0dDxfcv3k
Yfv5nUo713NYrJ5PluU91D1mf/xH/wOoIz8+aXFamsyE0bShMgDR9Ro+38oHNhxN
Zgiypn0GJp/2fg5hMNbXodZhbT6m/5qw8cUPbVSjeERsZOEmhP2nDJdkHB0hmmVW
oADyY+xF1qjeDcCKNDhiJ0/D9SM1aL0xQ2QBvSSmPhpCINLmbkRKBNap3kXlAw3h
`protect end_protected