`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8432 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JXz1+zHgF4n2s6TEZD4KtuQ
ATkS0e5WlIVeyjNZ91Ns36sZQfrQ9R4SbnYvAtVIyXQcw0dVgezYOkk9/8ZSqeWI
AIcaxqXHMCDgCJ/SFKaLObAx/qacvwXnWXdX/YPb2sPBG3CFGlmcbRKraOPywtWv
2OgZ10o25svwuQvjONk51JFbfFKOQVyl6n5eO+8YKTofmqCMbhrk+MzYKAiNVmzL
KmoMlMGHN1/BZwdfFbVFP3mFuhRsNsXyquUQ75SR9PEROW+4MmfFa/5GAKcWzzJW
pDmt7RZlV3qYBv2ERIIb7fWL0rMCi9gx992tDC5J5cu5P/H029oB+1RC2b0J+dT5
x79miqk2sZRQ+6aKumXeRe2fq+BqQMSHWsvs/FzndJaz4RBNTfzPP0jwqbQFFRyX
hrTErRHsfK0uDQRq+Q+hEMXZtihP3mR61OQkmEXQx+LfwoYwvidER0wdlgbqjKS0
Ko1MFKNbf3qkXUplLBCJuudfHWGUJ/qwGr1lv0Sxx4cMd1OkOOAHXwC5cOsCmnlm
V/p+6X7XEj+W45YGlmmwceEbwU/zbeMgZif0cKpYWBpYvpgpqTlGdT0A7P4Cx5hL
IEy8CZmlhBGj2CIDjBdFulY++TdAr8McVXfkPl/YZZWQvqPWi2pyv+KF0iX0Qay+
rbhJ0uQtm8Y1RBqfTw7kzyuvZCI95xxRzq0s5qgm0rXLQk/v8RFEUvMQqgMLMo3a
7xAhm3kHYLXTO6e6daiJlj/7arKUlQPPx3CfTI03m/se81yDCuQptmFcw+WXyWWt
vDxQozKZb7bVqjr1RZbDOEfezFdKfA2HywW4xYTUhDkKq+HiAMRjnDEGHv6+IYMd
/jiyO2eOySSnUe32wEpMsvSA+GwMTzLVMiURDWBbeGW2+N6rET7/NgImS1Io4UnJ
cTPir7PhoSMD/nGJRrqyGZ1nQS6Cfgen1L88jqDU4QvllSbThJst2HPo6yLqbMa+
/3ncKiwBFIYJfATT+WsW2MtwylSTRDds8FD9etHzirCOxc18FBA1kWIW2FvKO7/t
2wU2uwO6F8wJSgYOCwsgcfjyOXTe/tq44ljt6VZAbJeJskJirisa7kbNjPwZG8NI
j160ew7+P4cER+dIbKJB+0bBgm47DChrYweqZtNLqjqZcdovH9NF09ym7hU9qJ0Z
E6Vw3Ns18QDWJmHuWGJtYVFivZcvsY6xwTNWw4in8CV9mvoevb8vwpVCjHjT/LlR
lNId74DkaL1ltHouslug2fCWQ0mC/hrphV1WgpB0V9JLlzXvHDbp8ncZGSH7pKB7
DuKdgSGqc9z0dJIq3DGjq+QooC7UqGfSguBMhwEe+/nyWB15ZOU1aigCGpEPdFno
13QJD6N7uUIuk6lwPsOWjyjhXGjm101FWMUQrtwB3viKo6g05KTAet3Oe13v+5xN
r0Wwe3ABIuUVS5osJPPw/zYNDIlTIUKofx8CRl2OsIKzi6VMRN8V9OsPvjZu1hER
ltXi161ejo9ohaZqKs3GOg7YYanc8/WVF/GDT2kxDUFSO7REGqAC9dfo+vk2FU3q
1TUlZ0T7eZa2vr7q3zWsDAywVP30Su3m3VCT11XOk4gmEnEf+HC4h/stv7gVFqZ0
ZiHz5Wg4WDSHFaTy7EvmY+tLPf+xVijpOknPjrc97sTDSpvfAjkpp3qw3zuzCL41
X3Ij6YInLYgagW5UNNFp3enH69VFYXoXBZJwUZl877bvrJ1EAD9FiWxeo8536TpX
sB6zBE7xf77uhtvKUecULqvvGhkUF6jtG/oKxRu0/6v+ZhYc882dscWTRt/vqbJ9
F2E0tEcLgZ6Oc8YCFhOUJbXJ8tUeCecLATbvmE0+Dobg28hFje31zdsI9WoJCaSU
2w1IHRWLkMvPp1y8CVFoFG9Odt5A3wxVoNCT9hn0aqgKAyg+6/4zoQzUDFd8rUW+
UccudsrL0iIB3LziD/VYaErBp/odDsNdS4+jyvomQk44J+Dg+Ro6XkowPVyDTAl9
cuSc2VGVN6lgstZyj2QuDT6D5HNrc0dOLEMFXM9DAlbhI1JRMAyYeyPFFjHk+0ha
iKV6X83lyAkXhwdAow2/DkUOOe3/ezSLo60jaJGL7qNph6UHKYJzuZ+/AD3ZaLad
WkHzKzBnBFfABY1nuYD/JS2rKrBRbYJvxVVhVVk+lsQy0IVu+kOadtueyQnuQ7A+
K2ISgTEgV1e+Z7pd6CC+6CE2k3DUKRA5v3vq3bkgmUL4cBG5/3UrW0eoHwT6Gi+4
N8SzKvB9v3q8S7zGfWcpL92HYyZ6JgxJR9MV8+eBNEOThjiWcamnlPNJkRsskxBF
GXxJhVN/1sU4atsSipuwLJFommbtxAGgPcPz5I2ARlu7kkrBmCViWS6P1HThMqOx
Vz8O40UYnLCwWryqbS0EjhvBCEVI5rGBlHvaQwM6gaUwH3IZhRFF69rJcJbp+P5m
7GEFjaLfiGpeapLud9vP9y5EB8pIcHnYHCZ7L2eySeqzLwsoYVRZScesLrY1u1S/
BxgzPlPX7ekcyK4g0c0vLgdHGi55CEXBr+f4w/hyR2BfuVNwEm6Kpg/kIvxJ9A/O
yEzNB7DEWCQl3gFH2qjKdzAVh1euOVITkyJI4/RzvR/Yg+ZpNpijJtXYT1qwpntR
JVLCjc7DzixccwotU8WUleynYAqRPy9zlXDjw3BqefM32rGyRTO8O23YepvbFWdG
rBLPqgPzUsuDlqGzOzHAEACn7Yb4PM7GFQ86Y5f4K1fUIyeq2DkpQVvCCb0QF8A3
JA7fNGOYS66zXUdg9hoLA0eMBnew7NdIWttpvutQEleyG2nhQb9XiSHGJv058AGi
5nt8g1XDb3+fGabKZv7ebqSfGM7T7MjwIrFQUaEln4b8QPzayNf/KBXf451jFUdt
Ozha4xDJeNY1gSIr8mMJjaiNP9sv0dk/2omTTT9ijubcI+sKocS71l23vuuD2CGK
gBbtKnBdT+wLCLuS1kOwp5wyhregjMpdwotvwgjfvgYB2wm8Is63K2nMkYhUSMxt
xxZwHtKaNVDSvDSmaYSBH09G0ktq7BIkKaWVTBOtlBgB6Y0YqJHOFGspAVLiS5Gq
NnOt8gApRm378odf8ZpK2rzuDOmuNCIblCiweWxEO+x6K3FuPx9KQoj0pzOOelfH
t4ut49NKYfWIZGNI558ERIZm604OSPggwcODNiJitCdJ1QaETh3GmPOlMOYwvb02
Z28PGZ2CSipk2djHBRTbCNY+BTxbKx3GA6FaGUicOFx5zCRhOwPH055GZNtONNG1
ZYENkiY+9ILSkdSTRUW0woc6IaFIDIdR5eZXBG//noC7su0ABavFf9zwPsVv2gcG
cYYz1/8vDbo+USHCDQSoVOXBxI/py8KtbY7RpONziUUzFRJVe+463ItUM9RBQYLV
6VjneTiEOcK4v7QPkquLoq9nrL3yiMUcTYDca/LE0bP1woSioEUgIaAMQJGg08hv
PH0ScN4pfiUCoLrSX0l/iTiKmDR4vJHciNnuN944OdYsvEQquonVje0DQrQ8pXgl
fvTRZk5xe+/48PAQXs4Yke/PFfiSG2YXiWgMfir2X3bk1tWdbSl49ccD3tVwUPPz
fwbpc3/FxyPlhheSFgC747angfmU2puSZCVWletB7Im+Gbt+H8OSe5Vb04tMwTZK
QUjOu6D2FN407gOG10+SmWMwTyHAx2P9WqBPmC9q3pqlF6lOc8tesOzn2mtixFg2
t3cZSMBMZzczJhMcgUhJ5QoSjhxvvfZkij+4sG39e3ekGAbXDUJDd/XgxOh7i7vU
P6A/ZykTQOegbcHyfbhyew2W6WeUQREX9c42dSlE+CnktN7Sc3mdWCQ+y9j50fRA
7wQUcUDwBfRZqHnBw0/ppdsXMUmr0IbRKFwe3ndaM5PVfaB8E4OwZEYaGzaXbSZZ
NcusmVZFiGUnS0h0RBOtkE5a3ULCHxI59EsilRK7tPoUiuzTharg6TGr7eMKSJdp
u8uTvO5jnHES7wj6X/nZRVuHyIzBpoiFOOvdVgzsuXw6sUBX86hLU8bzTyGiGjaa
kyyKWSsnNFFJ751uyWCOFsJqlEu5PeTv+Q/M7yaLZ/8iHnVzs+vGUA677iDTfIg0
u5/V9Czgc/5csiW3An54alduHpOpthvihgRRGcExKAfSiAK1Hx5UEinET9cFxdB5
9jBBICcllDrJrdRvnS8LMX8e1JaQpuzmyAXr9vZID6J57GFXqZ1H/eC2LAcCBKbn
CrSuT8OvIopzvIimypi+rmAygioF52p5R3a1Xk3br6BzMdYv+cMygD4Dksupux+q
SkGhMqdhQdcOJ6puWsTT8QNIU72UhfWaIQPORDSeCmCwdhESi695rO4cCxMPGZSo
a+XTtC1OXWknkrUCCPnfiwrgv1yZmjhuhmTteZL/6NV2MWKgTSAbHi2prEP7ozib
PHqAzRJSmemXfJbhN1oGdissDMaHrbTlQ8zpDeVQIGi3H2ClYe/dU5h8bB4qkhty
eOzxlpC6Wg45M07HyiIovswTW9s95IqDcVwfMFfiWIG6uCH4kaAjS/qVxgzZoj5Y
NSXS8TZymmOu2DrVGbCNhzyTJSUMOxhtdDZ3FTzKl6+O4DIvhcQl+90EbYmnInlH
xgiT3WBh/hKX3eqvS+13dGMC2R5ETJEvHP16BVd4Jblw7RW8KhNUlNuq0tleokq6
UhK+U+o+CO///w7AW1qXwUhi/j5SNSqmhJJDf8X2PuqZnZcU3UdlibEmo/wvAyP5
G+uw8nH//LfXl0AVQ3N0+tzXMHFZ9er1JrvCz1IfLZ4H0UVVMe9GK6+Hg5J6EXOk
+EWyRS3N+Q4lcKnFpsy5BsO9P3sFn3grjKzVwUKOAcnTTgGQypsHeiHdzukQbY9R
UCunQyPyWnSzJGonrM39/V4VHk9/RIMPu9DT/ML1C4oxztQC6EDnFklNhg4zoOdT
acTT6S9n3B1G26n+FsmsdYnMq4zR7n1ksn9v60pioF9Y1C1G4AU53i9yqoWxkcML
N70u4F32WH1LgVE89vM0Kq4oPWIVRbVAyfcM9C11I5pWLDJY48pZlZWAuxCPlnJS
e5lCfIPgsOUM7vZgTvtxwe76FpZ/6XCxwiC3wHdeMIx246UHK6kWGtdg+66JWBud
RedmtmS07Ij/kLKYBX3v7+2/Ho+5KaJY4NJBT6b+J+5Kf3zSodsO+d2JWAWgspot
xo/fKzrQbR6n0XSir6Thyievra0JGKBIER6D1odFC8cp3gWqxNRfxb+RDtZsB58U
UDCXo8DqfyAAJ9dUa2IgjBgrNz8CI7Pg+Q1CuqLcHYEwc41z1mXcAZoI4Xbk0bY6
ZwoDmpE/S/U2yJhSWJkumJ7r+IBEjfKK+N/NXU20VyB+NoSCVxb27SCXRCZs1v24
KZNcXSyn3l8y9o4++mgEx09WNTZC4XJqfSSoG657LVNrNMvs1W10I7hCFEMNlr5D
l07Ygum9esCntOqPGXdq6oeZVSS1QRcs3HfAzbYQMSW+dmryPyXrHSpXazbCFmWL
iCZ6bzFULcLzS1m2QTwlJBRErJhJqtgwDmidLM4z80ukiKc7UWpjbQWy1uPl8gMK
EXr0hpplPRsJ0fqIMW5Y3uBqxaj22IxWJTH0MIoVy6cYMyCsyp6YJwLLTgdDlg4X
N7AfVpw6vrO5TSwl2ToyDaUzQmR1ijEMFtXifa6nP0QnVgQRqJB5UB1ZzxWCH4eP
h9kroP13dsCg2wljfUvm4++45yIQ27240Szv78uP0EMvJHFHzuUfNXYa40gAyZR0
AwL+7m0oKOPVvPdBd3RMsSMTg7iVZrhBYX4O5TaexnwX/EN9qR7y0pHaHwFTncyu
cC95D87mGwQGhQ4UBrDaH9F3MM+ppclXedx6hz6TUKsn1dA4/zOVnyH0M9Kafe7W
O878FylYl2zQQTXrkf0XY8f1Hy3uA/KPwSM+9MoOD2INy4WoVtuM10GRXHTKxA+V
tD/jxxoD+oBA6H8cwJNSFuPRyVlMZju1Icp6bQmyoiEVdhN40KmoBXKCRgo/sNsL
ihpUk76GRRxjL+DQywPR+IU6U1RnyaDd83Qfeb5tRamf3z1uh8/ozXeUkidVnlXV
KGnetQfjKO29/xWMpqKoee/oRD1wrATpxtcYA3uS6RL4+W+FqfFYBPkISiwtwn8+
gFoNVZX8OQcvYeDv26NjmcpbnfTWMCfyPhQauRTeXm3Sj8UEAsADC5OfkFXEQ8eb
slw75wE+RqxqTg74rimAnf1QROf4NNC/Kqb1LsKrmjeesNdPpO/8VgRrijpD2Gok
ghTkxA8ZQcjVrdSRVHSei3BRrnKk8UwawvVVCeK8QVEE2GOOp5VPyJJOAAPAEzuP
anw61X4VV7PtDh948rAPd49nOB3L5QbjEXv0UEtKi0AkmBwLzVkYnxTY3DC0u8yW
VOCEkC4TN7arSkZIRTOZA7aTgNLNJSmN3DhxlTrvncLKTkOzgMPBbZ4rQUihbS+3
29ZPJ5bOOCe1Eo9A8efCm0T/KcUQh7GYWh2YTbm/eRZlyUDRr9fMz4mnnEqi92S3
b6ljyi8vsRx5xBnOFEJdkOrEvmqyk79yO0ZOiwOzraWxldKl+mLNJYHzFVfK/R2G
1riD+XcNQfN1CIkDjJjA6cCZYzvtU8Sd3bB8DtFcZg1ftCKDRBU3ulnGgBYXTHjE
ZUrvHPJssZXJg16VSy+U5sD8QUqKeZOTK8hvVWVJEyel+ni2zC+8xCN+YJJmHywt
y9r/9RszTgqZXpqgOIcrMnTpry6Sbgle/y+UKJ77ycTdsrKUCvALpXBPbpLBe1Ld
rsIdbmGgYB9ztIRuRdAAyFxHXCZhZuPFxatYL+cM1MhKLXnMLARqyb5288iS9zYT
/O82jKLLI62R1LHRxgNeM+oD8sd4R5hQsVyE0DQu7ZZWykYSNOjK5K2mvpXpAEvq
mXdAeMeFu1r4Ym1mwy7lzEbgfFPATll4Ep/Nq11Jc1psEmYs0CaCyRtNt2DZZLmG
bav+Sk0BPlytryK00wksfSWD6Lf3BPOB5gQA71zQdvj4lOzOhJrSpaz0mp8Xorp+
ngTxOMB9gk4LmZM1/3GXNCGO4BOUaTIO1wvUM8pbhRyo/9olpGaZ0vd+202nuJ3M
8uxuvgRhtSRd/n5HeORvzAVJ/Q1D+ov10Wpp3LpBV5aoenfF1PtG97Izg44mHPLL
eX3LAmvUo6E1/9zgCYLMXh6mDM2JcyPFRsdxFNjkH+sng3lB7+zi0nnIqmZO8f6s
SwaVNd/GTdilyLtHp35vK8Ofax10N6Tgeb8De83fZSMSAMdOglNiGTDxCBbA2x+n
LChTykwIifolq3NxOMKTeUhFaF6PYich58zxRUwddCmoPYInHRPloIradUovccWH
uLSkMx59s2zFT+h3Hu7O7xO0iakCDdcEKUFjiUiBWNUAvXyXGbFVfQJGPeHwkZrP
EVBZBJxsClhEF+nn3kob+9mkiSUf1hCWfY5Js4Rt08YDVUV2acLhSrxMklZiqhN9
UEeA17RZvmG6g8BW9X50y2xRgdv7EEkk4d6KdyT+2Lb7Ti/Gx6wJwnzVO5GiDPCE
FoVAJKkWJy2flh4RE3FChX27QyVq0l7lAGgB3daLb1X67fchKUfTG53Gfk/LkF2t
nmMbhcqi8dSvLACB2zoTF4Fu6OgAJixWptniW4wndXsSwepfKtHgEJB5sADTSXzJ
DmiKAzcNGT0Seo7G7XOr1LcFIYEVzKvaKtfhpLFl/HxeGrpYXDdIX9GUCdHuHdnX
8/1JCPu4sQxrwiR57NImcSP4Pcbr9gb8+ypIus6alrIrnsjkYQsFDb+oULmDwzqp
tOH5ixM4AKlFaSWoAoz01uWRx5UM4T6ZafwJMasWVYydi14mlNXb5xM/Tpvri5lQ
88z1Jsl0czlvDKKtQxy91blnVzcrtuNOwn7Xt48lTMS6x6sieMdk33HoLHYjEAoJ
Jh3RDgtQ0sZ/SVRKoVjs2XQAyMPTLf5BLHNcPnyKpE8VkRvLyhzYbbY7gdFFfXX3
+CgFL0MHQ1hWIJ26iNEoIhs+aakoqebQLx+tGuoBjExr2OdQ5zREOLZik4T6efZ0
Juz3CUbHf80odZrRFOqiAfF1SFgzPVpkw3lF4OwYjzppoQKTBKED0xVV2Z55qP5k
Dj8gzj2BfChwDrK0Fp9+dUoH6kKkuOyOzgkT5F/0SJkPdxK9i5Fb2VIScMPD5liu
iZuU9llP6YkQLx/cgPUNZit+qbMdKRNzJN0ZpPBUUenSHvaNCBQkf8Ll7+oexvGZ
csEwuCQRVIn0CDDczvT1VytwMo42ZWm6IQh2V3JYosxdzCE8u4W2nKMDRqipf/Sq
IxlCE1OztIKeLEZxJtIRY3RYY2uwv7pQSdeG3K9HV4D1MfmjZSawr/KM4KWjnrpH
Zw6VaFuNVVVgN90rPXea7ASkZ1XSn/rFMIvJqnzjBkw7RgqGDL4ZuF735oUgCK70
7IGvwlSl4hvG0uKhn2qyNKfQ/1/jFIzyCz+cRvqD5FL3iBNMep08sNorNaeuerVg
8vOt7ISyMN/KuIIUpxisprEbbqAIDD50HSrCaPWpaFdd8U9FAMyt3N14heWrsjxv
AbTVHktmmt7TOZOZqHuLoqrd+TXsijn9mZMx7NZxdhn23a6iyO1Z4tobP+9aNQpx
LrorIuUWj66qbCDgXGMWCf7iJA1dyhy+gF5MLcTYpr+6bdtvLOzgglfBcDZtadUQ
jH8iz/Hx+rkmdghIx9Dn0F0mSyPi9u/k9KqLaKxK+b/mxSm35UKtQS+rqDXd3qBb
I93clBc+0Wgdd92DVhOeEqv39nO+Z5bNHeuSIK03NrRC6y8iB6osLQmQdfhwl6jV
FjRkVkotlNgwiXVVfGInrz0mwb2brEJdI90pae/iR9QL9fOmSZe26pTA2aFVWu15
LpIgdPbX8miJpk8DkSmG8R5YV1gILMzFgU8E/6FKJOjb6mXnoHBY9oMb0or4IuOv
6vnk1auTAkAmdI5wdWl5is4CJSs29LNWmN0QbeNJMVhc0OGsDr+iA1Qg3yrWAU1g
kXUpaScOS3uwvxlyW/SgI3JHdNT9gLpnvRw2PXty2d+24MHPcMG6fqRsv8xdFDey
pn3/Onl4D3/YpatcLlIFTxn/vVJalLPZgRyTGHQGOf4hs3nOo6lmdPftqdNqJBEr
p5l902IEYAhS4iZ18fpCR9SqfP/FP9rXrPwhEM5z95YLGRPP6cxBeHSkA8AiKvM5
jmtDUJmw/AsBMUZR3YZF2ltPW/ZIH0nB0QqOxrtoh1pjsOCoZ5Oank/+r35daB+h
1UwwG+G5zA6x/v/h8sSDIgN3MnoqqLUtHoPJSYde34eBoaUDqcmWLYleRqy1bR9K
oPc91RtFg5Ee0J3oXTqbeWI8yCRZtVU1NLkBMK1lqDZcWAu4mixrq45WqsSfIB4M
/TYwQmWiFNqOUtUC0eL800Cl4WwEtGtLLae6p8yIhUArhV9W3PUXPf3JjuTjWiMM
khofaUbKp+ducUsnm6UJBgRjYyN+MchP50AQlnBTaxrE0HyOzuKMZYJfphZ0+cgN
+d21AjQOJEBO1y990/FuzRLCOQNIZmYC0YkbUP3Y/RizTWOk73vWwFL0RjsgGHYH
9AVvWvaiotstAcDsWNFu6D38iqHr5IeqSNPTJJIH1hSTt1eHvvNlTLy9765oyQh7
6LQezs2qWJWt3gTt9Cnk7HFQFDmo0k3WpZBg95x8zN9SwIPXQLBHOkK8x00n4oLF
iE75SX2vSnetgPFzQlTG8Nwhn1Eqjr95qS6i2jkPM6j9fuA4NDl8SLlJompdy4Cr
/9fkE9276tzRL/w4FfwnPSoCVQMPT1/6QVOvE5gPOeAPk2tlEDpz4vNs/J6bWG3D
xHfOvmSS4PSS9BkvhkrQO0E1LyfZLoVqvSR7OzwtfJcrD5AMNOGstK2CL7NLCeKO
f/z7AHJr+hwzoUgZLseq3OwdDn17Jzw4t2kUPM6XZgQc0rjLS2FW44PiebfnYgrA
riYd+TrzJCyeZM+FTjoibzg/KNzi41eudmvrPglKYqfxWV45YgyCz335saxu50XZ
FWETzUyxaDIr9ilpe2TMRl5qQv1wrPNwy/52i4wJOCUOriYc2QcFkwohG8B8o7RT
xlBNpq80vJ4pChYQTavgXQgKSq/bXL/6a7Aj080bwBZGng1hitIOPg23qN8urw3P
dqniQDTVDtW6ADWEpjGXFpH80crQkNCR/q9wbnP4lDdbWW9+6WT/qYNUleeay1nb
1Dqlnlxvq6LiasuTR05S33PXtX3T2GXpyfbpCefPYVDx4aglkRP/Ma0Mad5brJvQ
4MMZakPbqCAHVNtzzW+2PBVL4tkFAaDnJaPjm8d3EbBI5muuK+ALtrAxyP4rZa6k
E3fhrSve0/CRAiITSv5MuDiIYlgMvivacLzTZ/X2Zc8SnPLN1yVeKyKCv0n6HKKg
Hi1OzArpCPLrHMUR+/Fs+pqaVhNO7nDlEWSrI6MU9aDV0bZ5zm3atjUsiqqDv6fE
ZfMSoXhbEhZJa8+LOde+0LQsVSVpUh7MyurudF5H0gE/NAyP/95F170WlRb0maLw
wM6tKmOqpCXcWsWxUs1FYj455M1c5jl4+MvAuQLrNepUfM8s5xLJht8ApogQoGvQ
0DvqsD1wsAuFeaAtgzRfvfdDrCui2mpBBt7unuwuF/32zx3XVvHNUNzA2P7N1++s
uAoX0WrZE9zpBRRjyAcQyWMSIIazaUJ9wvS6iQyeZNFQEUsWhGvGvbmdoPZd4USG
nBWzzgi3yVABRFVnzzl5yJzA2p7tYLCORfN62UgtOiaosWI7p36CHN+0WXXdslob
vlCHawfUTBxZp/tKLDO/1TZHJ+s05R9dOpPQ4C0MxY+ZuoWLrOKMPX3eOyQ9ItRT
oTBsyt2DT43APUVA/+VNFtTEuHz/9YlMa/x04l5FEMk2Y6zq3MJr7HsdxTJGFCzR
BooUFWH0Dzui83HP/P30lmuj16UfO0FrjCVSnyOn1alwQWb7iHq24GKnFWCm+H2v
lHlejhZFYp2gZUQtZ/Gum9YF3V6AJmakwu12lw/nZoW9kGh3WQi2wUvuT18tfhZ1
0JxYs7a59rgy9P22m9Jho/JtvCoH2LFBI+stdeMs18k=
`protect end_protected