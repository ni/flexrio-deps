`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5040 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
r0poS0ytQydMvF+aKdd0eIc/dhHihCiLM3NS0M3pwENdl+iA9bH2sbSINOZd7381
jz7pUKl6qC3208XdiyhmSDpWbNf386ff92QYPP6LJfb89+O2kaSIuil/b98yydIt
aZN4mizm58MIV3CyQ1HmEXXki05TUP7t4XBL58tvsdIzt6ytRPpcZ/zOCVOLsxLT
elCWEYpGrxWyMSoBANBJbOzoJCFNf1cQ3PYm019qrU0o55teIxnCJu7zd19Ah6f5
au64NQlVndd0+MEDW7wvoIk3NUFa8SVfedZ0wVBnEHVkAfsgdYg9zlphV3VeZTNH
BzFmBzTs++J5eBp0LVbr7nsuTY3OAPrGFEKZf7/DAejZq4+FPi8u2JkTs0fZm6w5
Oculrcwl8xbYrcRh/w9c3nfMMLZE17uxkKQc78imi1JGRWY/6xm/CykbVDuC5TLM
WLooCs+IxbTPyPhdWHz4eFPcrYCkPcOQca9HPaV9hntgvsBvhTWuv9dSl6AT2F6u
IsE6AQNZs5RwNSPJce2Nx7UruN4zXmOdGYHY2U48OCiqxW/kpFKKocL8jv3PbQXB
x3QWkF/msONkyIstu4miyaL1TvfL3jX0KwHA8ldPwdMj2NNBRoZXxFwYQxxEQRlk
bzWwPamwlC/e+x+BoSkJ5VLdZaT43cw/w2GG/DuDKpvTyn/Z2XNEluxWl2tkcCBP
X0bT0UNcOFV5rksv1YDiSEuywSOMiKnJftVgeOJ18UN4XvcFmq4267JOBwAJpppp
TGC5+ciL3yPWQmQHUke+jkbTz5sQijtVSTr61pYVNt7kiGybppr4RBBeKFry0+jQ
dFAmMnDQa6yLlLzvtwEYkOPXXW9Akgln67VfHkVqfST7YcVQcl8X6jhK9jT3T+gM
wl72ClFEdGX1BQk1GVL5TjwdV9VrJUR8O5B0+7C15SDk7Vf3x/60KasTrsW/mL+C
kKQochzhbHi/8sa1oUGCVhBmRmjd4gNMHTSus8GGz+du9RId/iHCcD+/Bvq2VMTe
/mvgjH/oMJOBtNgSQgX7NB2SPVihFVzeEK1qy/L/shrUDCRw8MTL/I137ucP6dDG
MErujRRjRr+vaOPOmq7T3Jm3n8VHiVwfecuuEAnNNwIQbzKN7vBFvKmuWDe9ZScp
kc63I5nfb9DpBTUEtwhEu+V8HdCWeI7ad2yvmfHEfCBQyvtv7PyO6QG1IS8jwi4B
nc6rHVo13JKiDSgSOH35Lp+nPYx4Ze8NYX4i5VOmr3QW6pMrKbk4FB2xRmjMjuQQ
QMkre764L+UU3juLT5hBxsGwTJl4tzY5fqGpsE5VziMYQEKIIuWeRGHjXKZSiclX
sx09w688iSAnqo7rM/pVpTWylPKeacMK9xMzW99I1y7ATgGGCQCaqkZMQMUA+p9G
R6ca5vDalr2oVathS5P0Pt0/99q/5tAOD1WBT1G5f9lDglV4a2FL/z1vD0ojOKh2
KCKleIq+1uPAy+b2gd8C1Awh542wXTCEiyZDT7/Ti6W4qDLhSx6qD5/GCGwoE67Q
ySWtm2W09xQZKj9L07y06xEQc4dTVfBIixdPDwr/a2TAf5qVBjrzwq4bi0OSX8uV
xriBAZarJw/Vdc7svbZMA6LwGATpoEKB4Awx5x2/JDr8FRtfCjKnA8QHgJVKoU9Y
vSKs1UvW3YYBDP2Y4j1rMW4ROMBkPTwKv1tITTzx+2Uq7Z1GYwhP9v/eUqknkUqv
cy2KLiOnWH/BEMn4BZeWf6vylWTr9+XmQ/XfqHARzBZtTooOqVnfUf7nXN6oABju
hpz8YddceZFO7T1nda+BJQal6iSdeWLRENSfjbJRdRS31sZPrS48YwwklUNbUdBN
QInK57Hbg7QEJ980T5AkCYdDnMr2DldZ9ZqFDuTO20wu0Y/XLh8GtW3reU2ZFdoe
hVV7S7pHRwlmJ6TopPkjK1sapZ8lswECJ3kPd0Z2HqkdZcrMy2zpypygt3MOBF1c
XviIbHIksQeAjlaNcxTJnQ5xcu++9nTpqaOPT1FalBPWL452IcEdPDC+VnK//JnC
e0tDVJ/uKnMM6ql2FWfjS/e316qc/AxwC73/1bjCwLqdXHaAGUGbk2d5t+q1AhbQ
3kXjil2sh8PswfFtwsfANDzPtEh7F+kyEW682eGR/sl0xfGSiecrEQUsBzxbeK7j
G0YdVl+PuJyVumySLtqJz9+FiglVTSKu1h7BTsPKZ9qJxWDDubi4yyZ6UP6U+9Xm
XQxjGSWYi2a/Mgkz0nANTrBS5xb9ohB3K2YQqVIE2snqOqns5gNR0GJsGtyONw2R
HWPmHkpzY1dBPkV/gKbwuglVX6kWEgW6mHpUlItyvh0tymSB9y7A3UKrgVSTK8QZ
yC1WQEhYYvYtSsWwDjsnmtxnqx+G8uIa/kl7tOSKwuc6GFnUAfSX8hRvi2mfepmZ
CsxOSSBXQGs+q2vMyCegKJzd3uRf6iQyB2ivNJ8S/6F7Xui4lxd6fqI8k70kdOwu
OyZNXEqRq7Znce54hXAqn56I4qOBJiGjXrn0EQznOGb9Z1vhNTWoA8pg9fpQqj1N
0N4To1KyVZAyb5t1DYlL048LPYAJjivUu9uyb/N6Ppy9yYA3jCq4GBsfkAB25X44
FFfxfakIvV9f0bS9SV66nUCFjACZj0g9MQBJ/tf3D9bDDhTiLULKTOMFG/b1yLEA
3dgDBPMSL532vHx4G/1LM3Wpi2pAAQRSxUz+jElsxqmYyoEwyjHv2/KlLGZGVk/X
fPRv6GfQzIz0hsVQYBFDvGUROHicQwhcS4HcKOVjVCrCP8YXZxzyt6gsyG5DCxnE
P1wzpJv6dbDs+mhEAfvyHMr25izMbax+Ww5pjOytrl0hatVz81886PSYkhPKlJQr
YyGlSzlFYQsrx+jdew9r6usMvhUq14ZPaGIXKnePxAP8CNzKjdI6wVIgys2ywF5y
StJdoMRgiVC0GfUVl4DB2IsVl4c/bhSpqs8zQa1Fn7a7OHHEUfZWvntofX51pQ3y
Lp+PdnazKINrt+I54KyhhAzgvcPDz+kfrzI8xYpLwcG6K2lXk5QYHBDCJEpbUOmp
4iw4+QwuVSTpHDopOpPL8KFyHJDxesK2OkOva2mFAGEfRAqCngQ2LDNLfpYfZubb
N0XjrPKxXd3Q7ZHUqUlLT7WI42ev//7ehtp+dl/2P21VGx9h2hl6dDAX/zIOPpcK
GJMJ2ft9qK6IU2YtcucWLpyPOyVcsCn4EcSgegmn5d1jKwSCcPK4Vi2TxjIFKDlR
wkQB/6glAoXheng125jkosCaz8Td4NKnz3O3374zD9kjwAIs4HzCH5vT5IzEiZ+G
bjQU7xuLvqnPchS5KjehktfFKxgjRkNAzuIb/4z2wSJ2dF53ZjaKMN7rcdXzEViy
os1GrhC1iFcLRS334uiJQfNTbwwPQfkUaFOKILoGPq6lirwW2WsPDJeH48DyHx27
wq4T7YrV5xMMzEe5Kzg3JKShcZWQg4mEFlblNroeV5BQBwlD72t+Zglx9Em4UVc0
PowGFaL1sNQZCNxHJRjgKbNplHp1cz9LrUKxj0lT6/wYqXs2X1sT1t1Q2us9jyK3
WptypP4uEHKUL6h3WFRxLvpdba/uY7kMD679LGNykV8+el8aLm/+QJs1tsOtmH+B
niYpK0NE8zofvOVw5whaPnLfqFx6CmPDzpaN48/GfptYyU/CnyUpxuO5CLZFGf34
snEswfxV1VXGLOi3LNVeqHdbRBBOZCsWtmMzoMScE9b+r+wwFjSbVww6tIu7eev7
kEP60v/wmG6dZfJms4vhOfKc0cDkniei1YiGlZFMePVAZsXhGDkAzcqXWpiIAHRO
UnU+setseOu0B2yAm4BFF9c7QSA8dNdztGf+fhcTqYc62rvs+0PCu0iYiB8smuuM
dp54+10muRv5icvFSRIvfgmkAzn80Uq7eZ6+mR+zBGTjtaG+GQZgmIX+tfVjrp+g
kz+d9HbbulvFAuWn7qY+A6wTYDAMZF7foFwpchLlFd7jDql7B7i+Lpith07RsJKm
AKBB8mZzelFRhPNXxs5oOnBCKVYdQyOEbsY+9TOHuW56KupFSSNVK+so3/bXCdqU
BeSglsicDfwv93wAw0CJE11Z1gr6FOexE+JDXkLY2giIn2pJ+UOH+xiM+7OW13u4
kzx0Vt/PVa8vJznQqOajImPgCcO4MT4cCTyQX3pZcMe/AowJ3xQ1QNIp4vr8Zswz
saTlPWPybzEG3IFpK5GRGlaxk54UOAH4xXPljJyPwZVbCsqL2HDlfPaAOls1JVFX
MpRJInTeKKwO9TwmrB3IexZtwCYxxD2fe/if8Xa7DWlyIAYMcHROJjj+BF3KHhz4
Iq1HnuN15Uujb2rlnDhk8QdiPM5dRZ0NqfhxdYGTaoGGJraDLSe3VfbmAGJQ5kqo
V7npZM1LWUZ3eh0DENFf+gl1DRvGsu+jcIsrQG7UJ8kb2h5SbHZ3+OPgRF4UTdBd
mAczdsJunkMTHYZWpDuixzWELcZvUpXPBbLJIjtSGaEcnAFMCjCT9np1CuQ4edti
76/5yvxqPRaQ60EuUgpZeBIJUgqo2dDJg/RsZz6SeNaWNkSX2H48h1foDY6JGPpw
wzX7rkCfSclD6VmlEEQYIDZcD3lkNZIJL5HgoKVmZ+Y7wf9bGV+CIb9YYZ8EL6l9
iBHI41Y4kcc8NLZXGZOw34fiVmaqF0Adwp3xbFaSveMQ22AmrRRA6ERyHwYIOH95
FpNTW/GccHhHuW3vBird3uC1Eb09SV27GPW2qqF94vIPHnc63UlMj0YuedepxduG
czwQ4WKXMDgG5PwYfvvOhDfB5AjarIZWWgendCIG7bRuIA02ogxTRokEDXZvbVIc
bWScihGohHT0qtjbsAv4NR5WSLVicE4kAvV3smuedNYHYveaUbImKPT0q1JWWcsZ
T2SxGg1aRYWbmfHsem60zPDvsnuYfF3oapYUm4OvkdNWnQaCU/SAPu1Z2TFFABNH
UxOoKXoNnLCNwcdxMjC7LwHI/5Vt+KFRRaF20lQGIOetHtnv7CoNiFN6JYgPcIHG
CJhNdGMy7RSG4FQEet1WTY1VQvMkEXRjWK9e5D3dXMs2VF30JDicla7RRCbxK3g5
uSnidzYejl6npnQ6d3Pr4yItMt2wiVtuTgJeh7r1hlMybeTVdjOYbmgHp7GTZqKV
pAglbRIN9eH4qKDDzrCul9F5ZuivJUsgWVlgdYlhcodHkWAlKcM3wx36ZMZCHUA/
wkbjZXpKH/TTO66xcrGjsLS+QYOCC08sCAhtXiRrOjw69fp/EKN1f0J0jwwAphz3
+xIGujflEnI0G1dJb99ckJswO3XvRADWIXNyRrRvro0STTvyfIfslQdjFoW4RHB1
HituxsI9RUBs/mRBYBiwrCGzhJvznoN2ZBr5VdvjBUaT8GPY7COfMzGiRJttX3Km
LwuvALdRZzG7Ptx+K4tiuH0jtMrMgayLeMWyc3UkA0EvMJcVrC7XVY0Fbko60Aep
0QD+PIOEBxqYjSCWrhFynZvdlw/eqpos2fHm/YpiXQx4xyGAPwE5uE6ghwhaDwhe
mYpiI+EpTnOMGctn5YNv90O3jIJXV6F2BBwaIN3DJT+5WVVJNOC10A03yWHTifoN
dsXVSpe7JvyQNwFri1YbkBKeR5u5UY7cDtqazz4JMjw8WKBzoVjVfnjdbqDUY9FU
MsMqzi1FkmJMapb0MZqVcwNZW7PNgbbllzo0umc57EAbp8OoaaDOCGbeA7VFloAm
bgs/Q15ztuQlaNmgQGr+uOaX0S88vpAri6y0GNHZavnClXkKHTyC0DBoZdg0VAxu
wA/9a519GrLmN9RwIfkCH+GkkXsFYxY/tt/ATDpVDHgNc0PeJl8AAEA97P2KIQ7Q
WeH9OUKvF8WGXOKgn6m5PayAejeTry9akJkrpX/dYxZdHiIYzHQxoUhFKo8l0eAq
Sklv/kMd+gBi5duKAR/1iuNFzgogZLP4MxTw8LY+OJlbJNxNQDvoALhYECgvJLcy
C65tYXpR75oWS4T6Sv9JCa1z+f1mcLJlMYDXsGVYhkituQmyeHv/0a532Gjne8GU
e4xtNOBBrvpPcfEr1TxNXBXrE7vkAB76IswCWD6Va3ybvDq6B+STWOhZ35FY6xPu
uC9dGEMQcEXA2i0mX0CBR4CsUOykaMu3ww54G7w6MO+fpQxkLlJ76+XVat0A/lJC
6py6zQsiAjvv3FYnR/TikDafxk+SrjY1fwCEEeHykOM4+MRRrDsw5j/xcDNa0fot
QbWFT9dvq411F+8bJhzovBI5GoZo5U7Y19BGoenumjhpiVn5jCNOMmCRVByoQVlz
yn3Yt98Zkn/L9qhK9VNvT71shu5Q3Qsz1iIz4CJYzLGFctBSSxFaAk7t4jv9soXa
ZmVxw+aBOsi4voBbDIPVD6h8/w5EaaTnDTrg6y87sRnLO4/TaNCG6pqTBaZMJhWX
QTzkAA58tl8pfs1tgGTvh935xH6+W4cHw7DSG5djoSqlMcame+8QfL2GeQbYzZyH
AWkRFBNufx/R/tJeYZQWnuB52Bac8mPKozPlNIwtd0TOPJ50Ab2Iuf9xyq0N+xZs
`protect end_protected