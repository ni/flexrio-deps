`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10128 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10PzJRff511XkZKpyIOZYaUXASRqimjT1PfOZJNsuiaG/
fYhJ6w5kh1+1pfPY8Yn+d7/ZmB5XpcDT/23QRArEacQzSsrFpNQ+r5A2UuAnkk/v
fTzOMIda2GhpMbYVUtT2x5fm3QAAczP7Z1YmsCpKIvKuA7iW7aq+tsF0dvJ6/95V
I17sd8SmlzHftj0m0gJ7/QwE03G0Y6FtBEWRTvX0+JAkrrsSBIF76h7IvObzjRC3
M2fzrtBEkthPMibCkSRfUXF3m+lJpLKtIe/YDtn/D0vNpzFigiKEkX9WMcCmIbBB
+2gvwDCEhMFi+7/8tT+5txvDG96WYu1iKKw7kdUtZwWFSwSxpt73Xf0antF0NLmj
sHDsuOCQoNt/fI3QHcwid4GaNc/SH45LZXkrXFeHR3ywFsrM9/n7PAMWoNX1Sn2g
LQ4QAyznrSKo0//Ch1bxiIBeF1+0+r6SGPyaCLpUxNTWTCUshrf6jhz5hbCJessl
IBO78rcG25K+MUqyk9nXxCwOkFg2yssXheQW41uf3PKM1NAMvKj6f5iIYlMdAF0N
g7T7GkJLFFAfwVqX/AM3mts79T9MRfSqklkq33s3b2JD4Vaxo709LPanbr/uV/Z6
E8ZYb3qKpPs+dkfegNsdsYg+LQQfMlm/98dGBB4FM4QnLQsNMV+AsyVKegDnXa7c
KNpzMRqTE1YMSX8DSvxsW5ZNNmMBBwP4SCFRk9b4He/AiREKym/jrQkJMoFD7uA3
te8SAWvmeKHe5+4G8Q9Y+0hBFjEexlJ6bkI4U4jyFkJYXLv44NkzZ+B8+3zoSq0/
mCo7DkwIwhZZG/odkc4uCCrJplFaK3UQOjKdIcABdVfKot4Bqsa95GCqywZPU1Qd
I7JS0+h82ZDzsBdl8FevcYU4UwpMY2n7s9szjhgVGA/J/rxnopfKyBM76W0TtNrW
OjBkKx7l5QZsdCzBUVtw+kpo1/c6HIn+n0dm4B4qkBlEpl0upQl1lAWrKIvmNTym
2pPyOQVuk6x0/ZJsHz5l3bBcpxDXzmVmLYBA7+C9nh7ypqjn21JSg5gG+RrV5opc
KQlh8AmfQmuDdHlBP5awL8PTXAdxYvvwd+gh0wed/YKshoCSqdQtTIMLZGgmgtOP
UXSQ46lU2WEZ1MM1sFoxQ9YyijMCjdoj83kPAThIesVaiczTQJQzkRkZKgYPpY3f
xuJMGFLDDTyBSKv8NXF1vPwHhGjS6aMyhX+mh2uPl3aSmYNjhbhObLdmLC7SAqA5
o5BI9BqW/J2XHwnVmQ0ZjqxMD/flx/rAPiIgXSjgsbnw7AF1255da+Riewb+Yb1Q
DwVsxkLKQx5qsf4TIk9nK1XSd3ipeJ2DN+8m/5vSoIQsxzLZ6fNaPBxEo6V5HvH9
IVRNK30BLkM90bOfI7I9JpDzCMLf7/edeBvfL+3NRD5Kcb9VUg+3WiFvK2v33ZuX
gkQYnO2JiTMDiKVwiZf1vj/LKMUfTw2wnPRdx4eCE82ABmc6mlW/JzoNi+0aLRQm
WL4qEky9t6xYreUa3JPsmbwk8Bu5mJ9Msswdu6Nb4e80tOnlUyJEFRn1IuOVP8D0
jjBhGC3z5MW6EC0K/k97dpZdgsP5xWSnXWiHnoNNkxh/kE7+3bHG0Orw8jMDk60r
eWcl1UrUGtnU47g3thlIpImoU8wgHkaKnUdiET3T/21PAsa6HRhpp60z3tK49vXu
Hblwj1DDe3+4dyDod3PVY46GMxC7RkZJcQbA5wZoLGHOqhijqr09UhNAkcd7pO7/
YopUWV8RNV8v98/njRakRztePCrul3cwSmxWkPVGw5R54PXUJ+YpvS63nLMj3dh9
Up37ZbhBb3MDW0bSuOw90+ANnIJHh/OwToHUevxTMXWl7/CIwIzfLSi7eixCfLOu
a3RQ1QUnlbtYi2/KjYDy22DXgA/dlhXgc57biESWElXnrA6b01LPv3WB2c60v/x6
RMzNU5jqvR0zoxxHsBEgcaOPk88ONoPw+r4CsdP6p2fwkQ2C77uCz8HJ75WLhDn1
Ctp9u4bnLBpKSxAB4STduhH91TgOpBlAqS5HN5pi/i7d8W7aFSV+AQBgNYR0UPUM
IqP95ySwLuVIT2wD8byzkhXkkzGrpVxlCTxdIa5RkDrSiZfBYNGj3Wwoafjo5ljA
+UUVG5RB/qAkdD3xOvBMb2vjoy6gTjicIf+EXfen8kZiztuNp0DbiLX3uA3S7L4o
a0yI87pEX+GZTVujjd3XF4Z0v7vf4oc+j6BnScADRNpsVnFpHxF8VY5BwSyG97LP
TSOTf83ghk3Kh2igzHuuladwFrY2st3XoPvkWabLWXzKkECka3SpPJZcJpy+LdxH
eeUwwserBgHlJL1eVOpljjdkBKjvlNH8U7fJC43xMF/r/NeOygExjzrsPEHFLihg
d1HPPhE1VOHSOhsR8LqOYdI/qXfErMirwAFQ6leil57ZHg7s4w8lezLMrnMFjqtx
rghdA0tZiQqeV12CGqKTKqyCgjkJCQnoymVCeDajRJdVq93Y5trxcBmPJdvDtyp5
eu8Oni0ShSuXCaxH37RGaB3a9fhDOoTg7M3DGtDxAvhPP6+06JF9GBXetBS5vocy
Gb8u0zq1xccLfdUHQllEyakpd+XHbeqaz1KYzqbrpgsrlYGcRQkG9SxJC57NucCa
AUZ76mTE7jEivAKaTdUHUI95QveyXXt7iQZNat1wJ+xZz65pNTJsae+qApsVvrM9
9ddKbKmCk7uFNP5GyyU8kNGWN2AvpVRTCl+saTqPu6LORZLmC/66IQNJDAH+M66k
4I3C0dzlEHrCEQa1vSR3O1mIUYRPKBXw5kKAKKa9FUjXAFq8koWc7qaxYYB2o7MA
5d3jcwJ6N5QGTrtFprCnzlwSpCs8xAGeYQrduc0Oke5Z/2WhibJ5mDDlYXCovNxv
cKkLfB/6uoSUdIuteB8oNLYONBpjI5BjbBmZF5DcNUzzP2QA6PLOM408mKjlZ6gc
I/pBL5Of/a9IPaHa6My7H5m56Ch0QRw+DknL0cK9nc/YtOPCckGPRjs3zWsg2rsH
EdMaYUYu0NwLOSueyKIRXZ78R54Mq16W6EycKcHKMkN95bzn7M35PJ1zZXFuZn6O
8AouzvAaBeLmcS76Nn0Vq8Xx6ICzVNC5xoTN/+QPoFl5h8chq02u91KQWU+vyAff
y8r2gkEurnIfHut5+WHAT6MWKbGxxBjmyFCZ3sd0gwNPCCYeFYbJyVGoymyPvhu9
swi1tNCkgoBugU2O5mcG4vFTwNC/UFVfuBf0+KQt3HKM4pJ6T3lSmjo7UMY5W2D+
89pvmFEnxd1jBzocsgn8rYvnyvLuk9k/wFcJ0Ga2hYm+u3UB4mH9i0w2Ws8uN6NA
VFTv0cuJi20PROO4HbLR+7A6qGDfrute1JhaevghKSWjTBGGiGaBkTkiFZ3bTkmj
6A+H7uui9MNljuN6gYFbOentMtmoxsgp2bwAHSiChnDK1NJ9Gh62M1USdNpH4v6d
N3/NORyCJ1IH0XKr73A185nWWjZNNV6u0FkHFVZASUdf/HynfiqRB9MU1Bvjt0Yh
XWcF/48Aav5ozmfodnA7xkebTSORZSwm3WcbNUE3D6l/xCLeTJxPtifbofpJGxDo
Hx1m+xCR/Zh/X8e5KbL8AZBni+9BxTxPwCOys6bYOC3l0F2ruFHQ4j+0Fr2umEFB
PjNSfY3gBzgCtF+yn63TcFzgU7dLSKDzFK4m5AlRCm+87BKMbDgc+EVSI0NHREuU
+mcE+VkAewgtvmTANJIA161LmJvJw01LrLQT16YZTjMl9xAWwVjVuqjcRD6B4IIP
akTEyIDwlHVifCgUCrBhj3SNHSpakNTna2lh3jYP3CQOPdA852sISH6oYFUIIPoS
5utzTLtIEkUaq75TuU2vgYSzwEuKin4XcWZ4b41pZ085LyhcmdVMw4/tbe5Zb5sR
Sqb7d1fSK/0AbjaWHWR8h/LXCXoRMMXpvMQzglIZDnr5Ndg2G/HU4cE19QwAr4br
FoTvDnx4cmY+HRjZggMwjgkDyit04sK9v3jKEKwy311KQ3DZkeWzpGTBdquAhUwm
s4CmRWUcxDCctZRtWeDSwHzxYr56UnyG4hmwejE/RFMI11Ep6SSS5AUG4aLG0sNI
6G9+nDkxrkRoIUb7E1wV+zzaG+VgZFOGaRCvwUMLiRMux+djq6fvpNK4U3hkm05D
fbZfHU7r2XaXw/LbuI5Rb2XSKJ/4zMm9gmerxWJh0kv7tJVtZgT9u3dDmDAb3Hc0
51dwzpfP8R6ekPJdtBZSgnBVhmhRfqmS3VLPRZlz3t9LwSBiZKjg/6twBB+/WpF4
GeOKVM6PRq/uVUTAXXpcpit3EYE+q9/Fh4YzE4ObFx+ty6iHDHQS24tZtf0nzmPn
ZsLh7q65ok8KBe5kiQ4tlPhB50A+41F4ip8pIj8iHIT71C8kb2MznUt/5JgyjtzB
5NUTyxnqpfoE86P9CxvHV+uzecXUBlF+GodFDWUvyITka0BBN8q3uq7KjN5KVMNV
pVXuYfrTBEOX9u7kBiHQIGQConh8PLzDJ4Yqcn/yki+c3V2E142QEIpnfpI7vVfk
WnPAHkMMtbosE8VhKHM5j3STATcWGJ/Tujd3o0U6oaXnE4qmPfyy4be4d11UUbQp
lCghuFGf93lkPKJB9MRWbXX+r55XVjICnWh2eBj/Nsf7tsNMe/DRKTSWGBZ1RfdZ
izzlJDx11QvuB4zydh6ogV0w6o8UZIKqqOpBh7RdRZ8IU5E6hX4U/sizEkfSNFId
/Ed1atQs3s3Kg5c3Uvcpl4was7HHCXcBfvOLc6LV7ysptJgA89GGFZt6l2LQENGR
/wL1wVCxfnWvc/XNDbnXvekTsjvyfnz+Kv8FuTrQHZlrXjE1IzZdGD5RQiInXGOG
WnoxARPtiBBzw82amEtRCck4IzvAdJM+jT/V6oTVoGJ521lQP2KJpOJ/NXyWr7ge
qjPwyt11wFcXicwHKUgUhibfm390xxTRWFuAxPQxBq9wXNJIcsV+zBZqIVaRKMRi
FJ/1Fw3/y8tZVDMwzXHkARFF2zoFFnnMeBLgXRNiNn6JiMVpe3hXpcysBkZgLmSF
cf07FBC8Lc2O0w9SAvg+neK0vlrE99d3ntg/mrvgph+Y5IeycAxjJlrbtwZKC6qU
NP0upSb1I+KLqYbKE5RPI/scIC65kQ9vrbZ/iqOLTKLrLeVUw5f6O6s3zlpWrQ1h
mUuS6LWcY9v1wYc45fQ4B/ucmsq7gfRkDd7NlWxIDVpSzePbJ+6sRjmMR+P7vu2P
GQ/YHL//DZC5ixykJ1dUYx8RK+aNrLR0Z24/l/y1txRG1YpRlefWXjvHj5GiwqVX
uMZbpLTYMRIWvZapxZ643CQ+JQou6qwyuZKYkbkSYQPEdwC0YIPYupl97u2tYpJj
hQoSQwvuqGt4mvybKAbl+yFKivbm0NF8kEQ/w9zFRyveehtAOg8BVigtndnG/C63
j2e2IhHlSJ9dV5Q4g9nBcRLYaTUn5kmmeodWHj7lge/sfSR8dctQSSD1u1VRGfw3
T/6KaybFfo5CtogzTWlu6zQ2Zj6JVezbs/VLnCRHTyEaOJPhNp99WZXx5FiYDPxz
ll/BBsGNgL16FkrBlzLIvDfkQu7QPoqQel84iG+6Ze0pJuJ4TcGehOEEUwSwB4V1
gVc5DCTDxSJ+XiOcB2Om0QJWKPWgEw+66L4jkC2HXfRCSGt7LMsY0sNhwzpGdQhx
FYNK6KjJ2aJsFSFGbiPe3CcDhPcq9gC5IWVhm7Yp7c4yIUf6DbfUZrsLWmUBfTKS
yOKKosr2IAZlQ7Q0SOTgWtN/wttqHgO8x1PhO5u/ZwXJUQc5zkmw8xF03CkRypPT
kDKWoQAJmXXr6dm6KEaOyLN8XTlPaLPzYf2WanmWpktybwBC+aOC6aB3+HRCp11I
E/E8Eo2DfQ8UxIN+yV3L2sYbrRuL4fff3NxLr4Gt0B119PwpwHcfp7/B3euaTiVC
fT8e8+yOFwz/4BJeyubYrtyPswN03Sv1JhA8mLYQRmDBkc9FZxNqzxmRUe6m5MqE
j4FhHVL/jEBzeomF/Wv6MKU++OJZUBca9q1g/oRFBY6ASxh3P0eB/mZUzsUU6lWf
7ftyvyl+POAkO1exOMBT172WY6DmlwZQf3Jo0+uD0nxQMV8lIWshBjaqx5W8683n
w8jqZZIfWFX0PYHd/J1KpNF9h8L5VGVZAkVKNTXHz8GP19CIrT2Yae1mwA70gNj2
+64iygNhvwbmLFEsP/jZSkYunsNoEhqBWdwPzmlkOYQH4lDs6o8be7yHvA8rc0g6
El+BSkjOTeaS1Jd1kILvEtjafAQOc3/l13Kx1ymD/1Nao6GiTvg0+66iArAhv9Sy
EHXvNEByXCYc1ywFEOklC/ge++4fwGd03/gIUevegwURTp1iXEvV3JpZVyZTpEMu
RFSgTkNVRv1YrRlDfWuO3qMJVpu9ozW+S81YnMAAHXaWNZXkzSQ/OuAZiU3CwmPM
qsrcIe+5VvpgdqeGpEhsZDUh32iqmnOdf7XkiWCIBUBHCx6vJYleTduOOQxn6SOu
f9NpQEPcp/SqIQnaBTqi1MxAuIviynOLSbeyklVg4njMkrU7fouozqKf8RBjKPAP
5/O8zWEt8frXmB1QqAJLpc0FwsR5YwFruyEXhf8zWaUfI+H1SN56/HC/Rzc45SSA
J3tl6FON/tIyQvJPF/DOUIN+A2HKn1xp2NwuaVzlgO5zlZ6TjW7BroKmC7YBhlHd
ywvFvnWp0PN5fc9OYgyHBtLHzxuxr/cm5B2GkqHd4+yXDw51y2t3tL5+CYs4D0f6
/QkREVQm96SSGPoXVAiPO1tOdmNqCwuh6IlPbxyZ1swqHP40cARz/XL8SSppTomI
a69F7pMetu/w9O7eEPYH1Af2f1+oozOsPo7iZiXOiKW+a6xNveQCiwLHH1IRolMn
JvXzxfNwjZ7lWxvu8b9GNxfUr/r7Zvjf3Pi01hJXUYZY6F+1dUhpsCzSqmtWQyRf
0rVquk83LTcvbdfaQgIakGbg0c/qf9xe8ahwNg0Uc+gmHMdLVUGvJ/xFJhMfqQDT
T4D4/E8qVxA10i1ZV++tlmLVM0b5FOvtHQx2eLbSuFBGuQOnM6mUhIbxIb4cBUQV
O9Tqlqx3cXD17USVGYWBKrxF/W/qlTMH0h3OVC1Es7I98ASdtogbk/XgMn9kfPJ8
p2ps9g9Tf1rnISLR9N5Uasxd/MSx8trO+d/4LudCktzJ11pYYfMEZjJdGq3ll2mL
3CvlAPeZR2ym6xDgTf86CmaRSHZplsRpa+oLtG/z7ApFwqQaiSzO8Tt8f+i4JcoP
0u/MWiQmElp4DkB4k7y9WsrwyigGFnmrY2meJf/2Lk768ZbFM3DMlHQcWrFM0R/7
STeEdJTiMJjMbxOhq6AKI1pfrDI5qaQmJa8SGH33YvJC3N9VIO1pJNjJVOT0nAxf
Slt2XQINvN97FZD0h1Hv0IOdsdU3qxPC5QGsfKsN7aBwNu0BmZQ/VDPwaOKDTBnq
1Li4vpodKAuVwjmDnsufvjUct9HJl1ppK13xSOhbHxkDzdAjvCx1yuq7ujKJv7Q+
+gqW4KS437U62RdecEGOExBzUwpq3IfMT0iW88y9OXcz0oaVDBIBw7jOG05alFkV
mG7bHNrRkPEaHZPXcBuGbGC6W2A5QJEbVuyP5irVIVZtaTHxmLyhEwHR3B+baaPO
/ShLButWkvPqhLr4drATTgJ130QclaNpZO8sXgDe/Ug1mtAz+/faMX7dyfn7WDnq
owss2wmC/ZfvY0VlraOTUuLlsRAArrOviYjPBq1bxoDQfQ40s30GqEsGbTXU7Teq
VvQyINMyvC8Uc6gTh3aXSo47oKdA1k/B4SG+Jg4ssZl4vXodfY29cYgWqL8VIG21
is0td2UtqEewcxnY5u8ab5ROmfTVpmllSHSbdsTX97xRkVtL07L5lfZSu56m/EEK
ifYaXzdDDj2dEDyAAEG6vbx6ltCZkKUB1/nR8kWeBmLxzgooZni9iNopomhPhJ7E
W5coUXJYR/Z6QgSZ/52Gh1iPfFekT1RwOceHERX8eCdF0qmMeukiCm0cc7KYie5i
miBqFRKxPUF604znC2mKVn1Sb37SPsn3w+dBnSXX/JMUq8BlzhYAbRSJuVBo5RHH
+GjrUadsKWdEuroAnjvnp4M3T9C8d5/9vqBt7xBbfoT9hKp8i+YwAn3zdlibEHZH
ibDchKEAaZRXiKjo/iaoqezraVA1g4J3MOqr6lZ6GF/Zz8tOGrfwsP3y0tJfsxaV
xppCIU2U6MwECNi2zjQmyeM/PjbIfBunaZv/0eNCcQKAwyAgBYUau3HaEYFL5/11
Di7hE0QoEQythhJDJ9rX2i1KfMECCDy30yfm8yAvPrrqW4++f0dyXUimrDeeJNXH
d8aGpoEMoEIzTtATsQDhNrbCtR/9dktmPlXXYFPcKz9sKKyjzh0UT2TdsvXlLcWH
IdGKBkOd9VULQ0rLe5qX5dEm6c/4FyUvLTzERmibUCX7TXUkYobAxxCEktzdCq67
tOtSu6soPuaruOI5/RkYS/r3OjdkRbYUTZPnVc8uuUoGiVo8ZglheWbFyT9xuL45
hG4J44dsrKA7sKMdWwtFvKY77odL6BWJLXnU0CxLPfWG+YVpGvxIbGM+Xd/Ayryz
ADBnJDZjVqNiiosNX1xypLrv2MqJTg/21qHh9LVlPeT+zZmDBjjATRQZfiakrIY/
3uoZbBPQIP+O6G+yiRXFeRYKRo8ufUPnfl/cRFS1wkSacCNvla/KQO/dAC1L+7+5
/Vez0qBbxbj3MyCxjagpTHsewJ+/vOaSswYFv2BaD7qOijehQ20ZgZCyjIRTpgCt
21TBCOLSWqf3r91cO5Z64ulgMpyc8EgSNFJhpNnxYwYIhJx6W+89KDiUlEufG/P4
h6D8QHRUfRarfqNOf9zoLNcKY8/0CeivDZfjrWsdwbCE3g1t2b6jRed5Dc30Fdlz
U8mMYzbkiSCUCmqztL6Ri7JlqB6TScpL0/5sxcNZrC/+w6HXdRTGKCTjx00jcJju
UByWqafp+zMvBWvP+mCXqrkueOZCaIiEBIV+wqwZv7Mck9QvfvBFmmkCJZJMnVPD
hTnK151xDWSRUJzF4t42sVhRvndAIz5bNsnaszNkeAaC+q2jc5pH13wUMwOuvz5J
C/a4i9421QPggkUKRE0TTDOGNXTbmkVgFBUIJRG6aaGYaoILTNBtUeA5ISL2Rfq/
bLx51Lhjmh5n96aUYwYr1BS7SGjcBHGWdyeZ3iL5vIM165VbJkQYenDKzsi2+/wb
ht8MmD7vz4snoeQD/IhNzxQlG8k7qEBf6K7MHmyjfuf4ZeqA0Kg/MEbdwgE6HJfR
vuN+yEfRRskSY/6+FnoyTNWVLtKpGdS4UMJ85k6WlT+w4DhYn+76KPQp4/fPgBAD
z7aa3zbJ/f1Cm/DVHS0uBEwptiGthFtVlQceVNJeFt5o7tgz0baqbBiNVkHXB80G
Dp6RsuBH4X/ev20lQoLpNs1ETia53YVDxwswoVScyv722aiZOAvP5tRaOqug7pQ0
wHb9qNy1I4zsNSaboY0Al0rYLdCMVI0JCUwVXNFGshJoqhHPCwudAYq/Obk4PVrC
+Y8Ah/Xd4SIkXJ2RfesNUZzcid2slIi/WObs+zNtLxymffD46zEdqV82oGokT9CK
LaZotNKsLeTXOwC1cKqIU0na8XueNeahSY3kHT1810eLxM/pOozSUPH9djrjogeh
OV1TYjph7y7qrlDHcSYEcbKylMvD2UbzxKhiIFFAnwWyPnyTagRupiC3bVcGeTZ3
7cjggZWngsOxym+BDizDIOI9OUGv9K4QTI/o9fAbcW9TXnF6ohKeSxebga0MwoXs
SsKtUWeehLcXUDHt++aj7XL5nDSzscaL2lppZa98alCgUUiR3UWAzVZv1OUludat
6NuoMvYF6hhLFI/8+GBf5er5ppXL+DAOx5Ee3Nl7I1eOLQp8BhwubG8SWzMxprw6
D7CM5eibMKdSXeFsyzLWTH1pUqqh1EZChG8bRMqGw7jLycTqHiggcd/CN9APUzQa
3/pVqtZM013l9uGzUSeuiTtqcxnVLarRK+dpMDgGY2DSXfRW1Qnvyp6DNfFOdOQk
YL2lxce8LFm6ht1p7de8cPQuyW3JoLaAE66Leq1d2GHs38G+ykGVk33yIJ2dgTYK
ChnKBdoMe2aHg36b1E66aCNsoou5qPkHXdBpr4LzKLYt2r2W9bryHrRLWd67NPyD
4DHqS68rHEX8bjFqH6O84GVV8Qvbegq+1lwbH/Nw2339go6F2JGKsC0/kPx+FYcw
pE800ZMJ0XulIuGDCZ7TPFjIWdrePKMxk0OiKyacNsxRREw+5gYzcW5EMqRpxt7T
TSRvW3AfGY66hsrY1XAmZoTVCl/jwXT38mcs+eBJaQZMBkc1LMxWynn8CyQojaYY
cL4qH0bRExormbfzqpx+L8wxUd4O0HmwiT9GbvUny5PTDC9zY1TTXHZTYSBcf6/l
OfVOj99tMfA8ADGBhs5gWBneAsvaELs3j1APgZewyn8N8clXckj/ZGMGXGjLFWkH
4dyqsZkeyhXSUfDQ31XNNSd3CSp0Qyov7m6oTU5k12/Ed52R3FXebSzjETNLuW8v
G1so5UMlEbd2rUggK1ZmbqKGgdIZW4hQsckIewrHCsGzFhCTCvmDDRyH4iabN2zM
lTHRhzCHPEq2LZ8kYeu0yb9Fmw0HWBZx+qBJUoQlWlQpYVUQh4tQwBwEy4K9Dog1
wt1kdRyIoLlOrROuovXDS+t3hnTBK68MW7OIKKhQrP6XuKgv1guLa/lMK3z7cZVo
MNneNOMjtOOhsUJ4kFsJOilDKtXFud6HWMZdoXNFcX7M6E5SbmF/9oKFoO/CfBNH
rio5fOo6J1Yd5PjEGdBjVvdf7bM0NFQzwY3K1T2tNqS9/umZF+zc/GKm+Zz4ZW37
DGwv7bmVpXO8/iv94L++CjjNTdM88TYxJ9JGExKt5BRYiyvuqLqII7zwOw05zNGL
Lad3/9AJr2TXB611LbQRIT62RYk1tuhpb13RONHTKP9c47oiyCq4umGj4iYWwqt1
bwj+kPFp2zXfPKvNTg5DKpHIDRscl92/9Sj/XyJ6Y/U19T3YgosVc/lV6HNLl9lx
nQAOFWhKLOazNf5WY/JRujmaVCoVdhjN5uqallDfFZ6fhyqG9OBezx72vSM5v/DV
VBYS1/EJSr2+HzJegpHlSR/atLz17BUERCd5G8eCR9S3LgJJjk/UPg03xJCjEpFr
dHz9icPz5LSH92nwhCOWUFhX1FygM7suSGXtp/C7pbi7hrYW3lWBdVZuLDn4cBUu
x6P8i6FyOknu4/c+KLKk+F5FGCsd/tzNIB6VgBCaqL1Ky0FLd6hpvlSABQvNn9ES
snT0+rt0BiwwsF3ZMzL4GcdhEGdlvrOmiV6niITJDXK0dMPmO648nS/GphXUhrWs
AP8BB8jP01JFWnZLmxhAkkmO0WSnFJmCYiYUA+rrJRq7qLAaXtMkSHVrdnPBacCY
xlbKWo3LHlUOPdmjF24x4yxHlEMVP/OA3MxhtizRTKMqCu71LjrqAY9+inBbvDgP
UvBPyXrKT12PxhtQAV6Oz00L0kyM1nsYCECLpJAKd9OOaNlFj/a8NEhY7d6OXCpm
Nq96w/oY/fLJaOUyQlGEyIquY+YzAr14bFohTQoqJBkPjPH38FSnDiATbsXBTVEH
rlpZ+SrO2whKOEpbWYZIhUBjcGsCkuke/xvBTgIrcjLrWR2vzYJtGAprNQK1Fia/
i0NvA1hafR2WVUgOlfFvSHZvt5IvOSp+eees40NWp0MZOj2CycDwI/ihV0rNGW4C
qI/7xrkeCpTa0eC2TTutm6/HgZETG5S0bPMdhv7g+DBMxFmKR5cp5QAjV+gZbqM/
/4nOvgZECQBN8HCOMgmiMCpJPIAoQdrVQsCLsKL09oGBOke6wqV8+EGPzJH7zEu+
ogLCY24zqYZkDSaONxPkhfOmSzTuLH9xUhKYfl7MDBYMtDrTebWmzAFT1n5aCEt4
orzQ/vCHLl0fuO0jEXNE0H+9HmqtnX9yHiK4YBxNungWA9n92LSW2WAgQN2AqKRC
EfpEKGL30W+Mb/WS/7y/0FFjO9B3SF0CsqPndJUkQpFLZeyuLgxYMUZACl+X0qxV
bICeLt+9pV6eLU0CcxAfsvqgQxQr2bOd3SYvebx4oUKEsNi0r5J52AnL9c0KNAgb
QzQqvCFzMku2vsiQOLo2nHXFkj5OmovVSRbWvshhRsr9aS9+85UisMxQTbynhtDw
L9/JU6pXSkOwa2bt4RVNfgvKA0lOfWAgvOdlGjbAHLI+E5NQpuiQgSSnKEVlNjY2
pJ+w23Aoy5jzzBcPZZ42qhc4A+bpjQ82Tpo9jNTeiucaDPSs/k0mQFCxvAJwInJM
eFiSQo8c6oDmDrFqlUzxXWPI2X7vSYlAu7M8QWz8SNzLSbN96T1cY4CId0PxY4Hw
HYGCoHwKVNW9YJJ41HgEc9Y4p2CIcPFO/o81B26dTA1oEE5CNZUeVsXhY4EXIIgB
vvuy5I7xCPUucA+gGuY0b3aZMmq/V5bkz9+0KFStJoHRst1jdbWS0eU3sy2J79PU
BCcwImMpBNO0+YTB5qncoWH5KXP/DbLdY5NzXixELZ5vwbv8XL7hN7oIfQvktMSW
LMOS6B33uI2O7JoA1rSXb1GhsqI2I4c1rKLIA12OBJWoxADvIFP+r8pkIzmqqClW
RnyfVVKkfY5VS3IWiznvMw1E0o1JTZd8ji8jyUw2alwpUfT9PyXQTKAmdUsOORg2
PhyMObS9RRE7wX2WWjplH/Kfgp5JTrBc2dadGuNxm5OKxUvs59xacW0/NmUGnVu7
xbOItS8Pn5pGx4nn/Qj+P7ZLajyFwZte9xCGHKHcIeL5MJRWW8tYgDZyWKIbdwkk
9d3MCuzCVYsf16l3X9NVwoSoBToqOclEK0dAuvMGAc9RRkKLJFo10+ShZ0DRLqHX
qNVa/+0f2PW3Q1oXydu1W6a33IBfbW+F9K1G8AYJiGkC9OUUnMvSbmnd3xne0Qje
/WGCF7vaoFCHTOTFVQXGkNYdYpAxkyF7WMRHIhIcuux7t8xkIiEWRGf63D6GKEEg
gv+qLRcm4Xq8hR64MG9m5Ym8x6WbjyKlr6Hiv0jkNIOv5Ehm2AmAdjZLqdocYbwS
RUXN8hf9YZIh2KMam0OFM8N2arufOv+LP8Ur0gugryC9pr21n/B+ee3YCD0qXFle
gnWjVXu7RydjYKI7bVupY6MIxO78PlG04GkaP+xSSOBlmUFQ7j242NzwCBZLfIzx
`protect end_protected