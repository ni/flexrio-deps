`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 200784 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
iga4gzPKo9olJM7FS8BWzqU0O+8WYOuN9RCSDhCRCu+hpwdqKSr41XFMRCltQh1n
HlfneL0Q4tavqqou84u+cmdWLu/K9HJujNaG5nzMgK/SRtVovJjFteJiPTQoyvHH
56zYaz1bYLVJGkdh6T/bnJGzPV2ZjfzBkGyaNWobpU8orMKkPVmCeaXWy6cMVvFU
J7BdQgPYmOHCiqP7O9xjSWQM8YLyXb9jT9U6HCXOcdvkqSKnGQPnga2yOaUKASoy
0HR9XrXn6/hWWvbcoTxg8r1oolz8xf4fEM+It+QEpPfHsNqu1TqCz9io40Sn/6WQ
P219zK7jBBOsWOP6B40tsGBKF7U10jP4qUY1JMRCXeB71YUBsfkHrjA5jK+sEpFk
Ox4MakKa/cbtXZPGYn5D7fSlzjo+6q3wYluJbMKBthQaUVwl0xj0UwEoPeMnhd/m
eoCXmH/SUlsKVtiSPiOUR9l1BkMZX0YxBAWVDZ55g8qZb0BPdWQcPQzReIq1TAcJ
lYDG3CM2De+oiK7WewTHMZdxZMT9ub30hbz1zpQIAwdNpKr7i6MCGXSuvivzj46r
mXZW+U9uMAxFFYWoZZvwRHrGjAz3z2DYC+X8AQ8iCFj2rpWmsBpQvMxwaolONC4/
llxRdx3qxL7g/c1jCmu95dS9u8//i3JOIsFtiYD19hkADDA7bTOwTTs411LpYFNT
3HUYNtucHPEy3bbhP7yRvghIy0JHWSk5qzb/YLVfVs+7dwgQLwl1AskANWSgWCFS
e5/AcfSBk/I7DUq8HlL/TUpvd5CHZcV0r0eIBVR0bEUmp5gm26de0wXfoc6xknGB
M3pP06WVAWPystuQMWKkzEx1XhiVtkArU4YA8JhV6I2OPdDKtkANXNSAzxwVMXpz
hFjX9+pFkO2W+G7M5p+sN2lKJblv0zUNvwABq4kvtuPPKBE6EU5xrmEMTuCxF+kt
7poQ5ewfwo0Yx+L6ho8BIthU0LCck6FxKJG3XDoBYccVNVlGxntFIO0M9J/UBFSY
efgwc4tV8ahENeKEABFpTnscONMlmHS/TJCJSH+4qdfmtCvUpK5DPnVMDal3aDNa
ADKkjCr1Ay0dW2IZ6/YxzVETTwShsWhf1TdOR5v45yauBIchMHNkvN8fn9wchMIG
/VMsVnERVFxlxBR9EG2YsvGSQpgrseeGwVcEjSNoeaoRSttX/99rG8bQUQsjA19x
EkN9LIetYqGudo0AVDfe6RvpzxnL1g3W13xLg1zMYB0b6F1w+lkd3nnacS+wCh86
oT2ZD0nAnVIEIXgiRFfL3zjLkMYKyqQP4RbyMuNbbBBoxcqvxdkq5WLAh+pNjJqo
dzpd3F9fwkUE8tRUCa9OoJhdF1LHY85+CCjFU9v3MKPyAMWEwzmKJeqXVlXUv6gC
vE+/MwSvLbLAZNEZ7+P5dTotAviPZOwS0lHIezDCjo1ugDByNKUVlYT1xuQw0Vq7
6RprK7MZyqFuUCRAp24uEhtLYhWHAjOYof3qphQLXSZqTas+7fkuoxxZ7RgqH24K
p2eSkuVjL6rSFvH0RIfnxGSS2cfG4K+b5Bt+Lv7LyLL7Zfe07TshC588/89YzENx
wHk0aGIFd+sILePjelM4nWgPNp0avKiS338ChGpU2uMMbPIrRSLBhB2BftrBKZLz
L4qjwfi7AYpLs/Y3MYL24hTMcefHcSnjl4AdejS6/xPtY5yhGvH9BfKlj4JUqGma
+xo2JYwD4DWa8bzKS5iMvNwlSUnJ0OkmUeHc6fueDc8jPU/qJySZFz2sjzgJbt7q
C7lcWsxfvKh9zkcRZoZWA4syh3L++uDiwCcMT4huIvR/REP4QtDrjUl7IJ4yPnoR
KTGl2lmshySVZhX4n4+wTfwnvGW/5V8/FPd5bt4PTOhm6/cQbLjzsx2CFWERWH2h
FW3IF4frRJe4uoJk4lqFDKKeOidChfUQ0px9KX85SsW/TJh/BL+pL2+FqW3qwTYx
gG5kqPJI5SPor1FZdRZ22b2Xma+LRjlKC+NxTarZucoz/ZmqICDNMScB5B36jN1B
E5IbBmePrWfQkamOXj9le9cSrMW5JYWZBVcFZvblXkf+F1ssqaBEwhmpoq01MSWK
dwJjJkhCWuI7gX4XB/0aSZVYIgh0dMeKtppkDb+IqHGoAxjTMmIJHl9SwqNiZiOx
j0wlFzFh8N21dcBifWNdEc0SH3OmWifBU0pS4yP+H4QhbZHZqk5me/NJqIg3egaz
psHeSxQZcfeSWIuRuB2zM6yeMAr0iro0A6RFBaPXaYRl8gl5xaeJeQvXyv2JpQ9X
8GQzzxMztizy66oPT6IRL/VRoPkTuIiTae9JHLLW73pztv2DA1IBVrELbHZ691Do
kY5KXrd6x7opJb8f2KKuou44vR3jdtXgwMpoQIns5M7MMjfAgmweZ6zW7A5h0HZp
ANcB/Ds9Slxc/v9FzlBM2QCFEvgcXGnM2Ls50UyuZvz8YsR7j0Q5PYf4gOw88GeI
/n4GmYc3fSS1QyAUmgifuXBH5PUAeqb/evutIg/2hReSX9UP6PYFWIfO3HwZ7VT5
S3QctV5lZ1PtF0x8HvpdBNBin++zN6fM3UhqrybFLnH4pAVxbzc3/cGASsm96b5i
pn0mYezwHqtT43lGOfxtWn3BB2eVIyx6pBNIDzGUsoLTkpJhOORtpRihLoDTcgle
hk9rQVn+Q6N42jmLYRIu+wHTLETdTSokjpKrLv3LxI/CSqhDE1nAjuTaZU0Tplfz
H2kfWVLSubA1quyc8wraaImB/oK3sYEUBV3yfla3Ef7XNQpyFyOaVsmvBvERaXAj
on0MlRTBEUhjUjfbtPtxmUJ0sI0JwP2nkNbR05iTCGAR+W9KncsPToPci3kqBCpE
kxuSe5I6ItQeCFPprZ7FpmigYF0Z/cFlLfGWXncoW/u/F4fqBWqqjVnroFF68HOs
sLT/JmVrczPQpvaYrlNCxn+6WkcN7NzDkWgM69Z6B/0WCGX4P4/8otfH9DAu17rS
GL15KbaRWrgcSMqWi3Gn+YL/uMBc5bwoIA76IRBdInwdA6L0JoFGurysj918VNSe
smV2ujZyHm1b39wGhmAXu5WQeOomIhJopOEIdNMcmvpfwH1XJnIarrkHasmbZURo
bIPQGWSUfSvp7ndOyGs0acY5SQHjtnnxt+JOC6jNJd9weYfMR1TTgOYQ2r4n5quI
he3JovIzmLog9iO4bkstDcizHIimrARqp6Ikrc1d8FQtl0rG44g4TX8bmzHWXrf7
UeBdj50Eh4s+V6Th/ncWTysCb+z+cvzgcrC1WyWxUcJmsndnPqQqpUH59A6TgOGn
cp8JSQMaGok//MQ+7CA1rCIWB5z1k44m7u8tRbE3bKw7eGFuiNnwyLobfEh9ZleK
3/c8R0yn5tOuJpkz44+2GgShFlaqtGBenOH5Ok0bH5YaVjtgazaSLi8KCjRRHJxe
JycPJ2HixSAwIBtPprnTSEv/q2zwJZHQptZyV9LhEasUqc89TgYWy1bgs/UJpgYw
pHzUYQFOalqw/73t82SYNsk+DO23MBKRVMsT/JAcpPZU4KIkgWeWdh+AwsdaIY19
e9LgPsMGzB67DFW5P89aGg17WXu6msfDw0MUt0R+DumaEAo24o5AUN9ootMKZO0M
1yh2zvdc/Kk/Zq6bpcBXbrZPp5ZVkgUezDIoEuytHQoNhVl8IJWebduyoSmmuiu5
rp98nK0xidzcXFLXmr3kLOArNFBywg0VHoXNx9Ys23NjxF/C4y+diKGtBlLWmjNL
6rWawoJEQgG0StoavHQ6eeb5CQtDXM/KnTIcG4PQXsugr/1CJCTMHOorP46NB36L
LYqoI6d/JQF7Rvzsb70in4Ap5t/SDVROC8iGeiqsZzqGaIzopsZIxmbmv+xKwwEg
STHQL8yHZTTr6od5tojzchek7l4d7tNcTJa5sP1upLcGDWc5k7fH9Z4zxhYeu9iU
HAI0iqG5zkVNpU8q8q5FT/dvYlIhSa/elQ2q9l8sDP9AinbNLsp9I7iL6j1cGOxd
2xm8MgJIVb0Hcnbd6JUnnPND5jKt1kwUy0CqXazv05Ds6E9upVg6BGM3Wecf5Ru4
y+HVDc7Kolr9sNDRLGGoYyMPkrW6kJDQPOPXsjRnaMUy41SYWfp+CStmggvk4LxD
SFfBn+wT3Unv71DkAoZ35w/3CFPK+n67ncRatHB8+CtaIdSoWpRMwS1dzFKbB16f
mZ0ak131XIal+nPB+EA3fixr8c6Yh8337Zg47q0TWruFBFIwyZ1vf4E1XProVsbE
gTYyE2NP7w8Cz6zee8JaXaCu5Ayu3E0i9xOJErBqSOsaBZmHu26/PM7wrBHKffkk
w7Hawn9fM2TGMfyvlhngX/tgP75D9S000VktB9vMnoko7Hs566dNLIXHSn6M4+AY
vcTPxAhB6dMaSrZSOcMNjBvImQec8qDAKqC1b/z60jq/1S+xGH/ES4e9bOTo656V
XS/lSLGksR8tuwssXPe0OjlgzVid5gzy3H+MiHVGcb7TcQKscWTBn7wNSApzxEhd
GlI+StRKLHHbD5Z2uLQL4qSNcI9I9vZfodfQ+mSQXWccnUPfEYg8Hfb5x9hEvWVo
H3XRtvQNSZNL1gMEveshXHvlIHeQBLnRbjCPB/Atbjb/E9Us6uJ8XYAjsqRFMQ8H
JXQm5sg8fsOlGFYv+rlB7DxfcIPqqBK9sxvKgRPm3M3p4C+CZh/kwJH8IyV0dUkr
Cq1lcM7PqxMb9t5FP36irX002HmsL2wIuzbvIXFzcKor13+IzHOEx/n4jwNbzYY0
Atj/++yQDtha77Hbx/icQJdcCK3+BS1kXlmQzQmZZDlXbuWYC752ISd79tgUyo0m
uYMqjFsxqS8UkDxopFET0U6n0S6jitTu8ByMJanvYdVWCjtpJr2J/TBJ9oEXxJj3
CK7wOJFBY7ylz8hxJBeF0wmx+s1/3Fr6PV0RSqCAGIacvEOIBR5G1gA3J8jzHiOl
+eebaMKS/tL49ZUMe+ZgZSh/zCidOcQNwCtZKfXSz01K1W7C5YpQDJoZIr6q8YpK
u+xxtxMq9vZZa7nWpvQQbAthzpD9Wa4jVK6dtYZn9ce8dFVDr6lVjb7CTSZuQEsq
znMKKSjCdEv7PNJn14E37VHuueZL+GooHT3NDXStNCC/Nn7tzI5SsNkKc37zTjtO
aG0WTYzKiRMXPcWFSTZEynGulGaOyt9TjiDdSIX06Q2M1j/gk9h3fk2/VxwvZ2kL
V4zpPJPv4MoJcTZq2VGHyDmWPROlzuy+iwDZhSzsOpaHhIu3dY3wbsS9gGer9gAn
DzItoVbewd+fsUTA6j1w6dTmSbawDUC6P7EkmQugJko1BbZ+dzI52T6+BznER8Dl
fb8WlPqYdw3VUFXRlfr/eNg2PZ9tXvtUSMVfn28X33SqLFQM/7yn+OSsUycPig2h
DE330qt9HC5z0AdZ2HA840hV0fo1GPW6roUAatNB2SCmIubfxaTAZUUwihED+Bpt
Opk5XomaYwsiTCuIah403g2rL+P0bsEGK9zwyuw42qfcd46vSpiHz6zx1LpcGt4q
PT/9mI22X2xsfFkucK/1ftt/zP9fU0F6TISx/C7q/wcYU8FruRGC3QSmHubj/tZv
TmfzDPNMfoTTTP3X2FupadLKWlQa3afay2mkJb9L3MnJyx+21YhGwCphFH9OIIZX
TuJ8jDKJXQXzrBdMsdMx/VMKf3dOnmle7tm96ZzhKjBFV0nhj9OwcEZ20ImiTgB1
whJHdXLC4BDNT7quYk4p8jpbJpDkr6q6cRgUcnwGzZ8DycOr1rE3s4K3hYNVPGMM
YXkq/sUlUlmm9iGFsRnAJOLjkU/kPCGcLkuI5MUHgW0L4GUUlezCN510WsR0714i
JkHgoAxEyqQmgcrudyAUYDEXOXrTSXrVeynEPmllwlm07khNBM1F9G71KjJJPKLc
HRxMIIb0dexIMruR3xJn/2fXVR4HAJSP5aBIWFtVz6PIKM1JZtAXaZpPu5bwDnj/
ueqShg/U8gawNmDyIQ6o1EIsokjkbAD3Ct5Cdb8eyurPfBOV4OqcDd0p3j5RwUFK
PKTjMeQt/QacmK3ydBl3pGyJhDAltyUh1fXDoljrQG1QQcm3MGJJzWwpMipmXntf
cbO8mJugso2ZZ96SEIkmBqWf5B8R0US5sgNGk/SGxPANrCi7VCz6QnAguKDiOj/F
30nMGz0NVYNAS5MIhR2NTqHJJgmhoaX888KyyFMKrEvzeB7T4QvoNS58lIjX3fo4
MHMMtJZ61V3fIOEWjOBm0JlosUjry8sga5MqleYRLxd7HGdZ+306SHuiXGdYUWGC
znhyYw/oLDUEprpzr7AiDqBTscGv1i4ICnrhv0tl7meh0FfUGI1KgnNZDZyQgYql
5ZIMDzLTuQq0yoRii/TMgUeVkxbcC+ViPJO8jxAGaY91n78xRrS1SRxXKEWSaWPs
orI6Hhh6TFXHXHWsqgu+FIalo/fDk+OKGZkYOisGnsTvTZ0eiX1qr6mLVauP6k2q
1d7FTPSasB4D0h+CP9TkW0ZGHo9jTTLQBV6zXHur2uurcBM8/1bpi/EaecsWp+Sn
nmcWSHGx24eL5GSaVknYHrnT6iqjzDa4JQzuv20oDGze74CdyZzCVY8FsNKes0pS
kIWkyDlcWm9kiUZRS0CllxvP12Zn1ScpV6VLBdrtUHLlj9WEDm3zriELuHAl7LX4
NMHQiI2pGzE911InVwppl5tFMqpB7ofdhZw1/qE+tZDshWtYVhBtvORM0vBKSnB+
DaAWGg3EN9RIjb0P08bmvBgXaDoySvmrXs2UDTFncRNb/WOcdN9woFftxBM2U5EA
2xPbNy8NQ+4rEgVzfdEQ1urE9QAv2fCUv7Sqc+W2GgrIeVSrGT6vphHs30A5tfoH
qooNf+iFDcZ2hecpptX2Y9jT2jLX/Ox5FxMqNUBFX2kCLOYxve0fYKCWg3Eo0/w9
pbN1MtPxHgw+bNEOjVfFqC0KhKGsE3camE+UG0lUiAzZ7up7K0EQXFlJ1/5M5neA
9hvZtJd8a++rAgXMUzLDy1bo07eJqivtBpZh34OIXCdrpWyJi67AnM4OApUOy0sC
9L2xJVrgw3Uz5jA0w87bN0HsX1Etc3IkPNmVFiMWlATM3450aRes7WYFEe9DBI14
uoq2QP7PSky/ZOutsUA/6pNwB/g9Oi00/CTtB1W4rIoYWSoRoYS5lAcMOImwDXda
h8yt0C+gn/Hjo8lPmT1/2Sf5jCaUJb2uoFOngpZcn6lXYu5jAmRN8WlMMaBBqQDa
mIeTQkkAz3UO6vYjjC5ehjo8GjzcEnUF/Lmb0BjO5Lg9WqowKXHJkWthn7d76Chw
ZINAPPc3Q+lLc8RI1e+wvphq1uKLbgCdRhatmlRx+WoHfNouP6vf8wOpqu22BEFe
heSvPFSwZM2ZxMj7AX6Y8qPswS/55A1nKcu0LDLd/qk67MStTN3yeroqz6qasXLZ
66kyXZxTXRZyE6zlwxeMJinSEymUC1OW4l7oA4W36ruAm4ZfGmNH6KARWPPx0mTG
lTH1m0BoXpsH4hEaqFd3tn0ajoRa0ChFBIXOfIJnRPFe83hs95syfdr6mlMgrTp7
jgyM8ycnksazXzjtB3cjtKxqy+BAPogYK6mrs1y1uiD5OnSM9xX3/nKk+gzC3jS0
RXTELPE148LyCnJe9T669YHvxOVcN4KXQy8YuV8P+tf9oHTT2Kr2380ORRZ0+xr/
DtnifEvBLGSY39Jpcv8PGRcyDkBkz/6WARDZT7G61uToJo7LP1MY44ymeFQBl4Cw
hyJOL6AuDZHo1p34vqDd7Ywg1hPyFX8EERH3gJmrcnNO6Do1ntBDRwY8A2+6G9U/
OIGwbGDymmKdPwXEx88PU4yocP5kqM0dB8ZbarsMBi5jH2L0IAZ9f9AosySpewea
c6hMN5JgzXsRmWTgaaIIFDybCFsAAfDkCGykDKXo7femAPcV6PsSoO92DjQuyQKD
30yI0d5ztvg7WE7U3qnyRzKrzky0kxb4cJvZ0pTh47JhkwjYOLuB6Ij6Wpk3Keon
5WNd3EDXKr3Ow8Z6g94mGXxbkhfSuNq1kvh51iHGqdwKyAT4JX46s3ZiUz5qq2YX
+Cc2JNsocOReEGnrBMLxdeKer4lmWEtUxqqcNnJd/mtxzBq/658LjcLpRO8uLQkX
FgJiClUpPJbK4j7rhvnB+JOc6wZRLrkmo3Qws+S3fCGXHrQz+gfeeYWsBCx8CIMd
/hr882wO4kt7USHnFyV/N1dUCMfn0Ch6gQF7fF1Gs0VDqvfZXOVFnd2hFbnVtl1Z
PZQN9esgVxc51U++TdUikOiA6yWtoj1m1ogO8q2qq9dCwcTwK8SBmidUb52uELb8
mmHm6G8/Acg/O8n+GvgVkm76WgRVLDQ+yckCz9He59T43yxT50OtzgQ6SHVb6f2O
HKmrkEGv4BKtNPcK0xXj32RWDfaUyS/khSBUEMdxu+G77WiEG4oB8UKTVG487NU6
EXMbqPVmAFolHro9AJS+7c6kcsfJaD8oF4cOHbwG7WMBoGMbdG39gk2W6pMSCNzq
EGgTHGrcXgrHb/IZ2GPiRYyU8Ll7GvOZRdsc52pcSkytggSLnU1qy2qCnq5KBcPR
IqgwpYItqf2VczMqVk4ykeV+1p5XVu4uxr/oJl10RvYtkaPsseCHL743/0kaf9k0
5gxPilsRdc0RxKTxdqvg9S+EDSXWPKtBvE+kFFGM9U8FqRTdQS1PY33QoNNmKECd
DA3gbWeMV0fxE/lU6uKtN4lVSuLQe/hqESQhLTLZtUa3a+j+R/8X7l1OpRNXYT90
jQhixn6J2JhW1X8Qm83nOd697lXSmpELyU86rGhOzkWiBXgzN0oEHC0CPmbVNMEk
JwCn1CU2sB8hK5voF+SfMDpL47Pyqe8WlfGAtTMlhm2PSXOEvQEkWb9QVmlvXVbY
3LY2AQ5vmnCHpec+ZdT+rDLxjA/5stVoyPkWoBhT7IGlBdhmdVN5QoIERUoC4WW/
Kp8jbkJJNlvvFuiu24lY3GYLKp4YO8tadKp5XfCd17lK9SEgzYOSymmbvKUBrD9n
3Y7E8S5aPRjqhcB/njDcRLernQsIGmm38TAs+eXr54oAw0AauxQsaSvPNIqvg063
FBikb6Ci3+7iEuyUx0erzEP+ncbCpE4t1Mn/i/25xvPZO3RKzi4vaRbbElxZa3AE
Dsw9Zcf+6x6H/9BCLM2eeH0g2x2bASlTLEiNKaVcpQqkdul01aJZ7FntTzuKGb6o
+aU+/8i+RCOP8d/aSS/4JP8h2s/aoIGO1hPqCrrlJs3PZkcx5gM5/1u8NV7TGq21
kB2caq98N51wvKNJNQzjBbt+Mwd9kJd9mDSUMvmbUnoKLyaEEKRmSR8Q+quHk4n/
LcebbIC3iqN6BuwTTTVe7kFbdrD4VQAHrxinQBPCcDkDGg/Kilje6yHxfVikbUu+
QjFxXA/qa8ovQ+9AU2/kDWH0+jWCsQZ24nQnyNM8pBj1J82Cch0gaCCmcg4XktaN
H2JDMPOPxGNu1GDgroyh+n+n8zG1uaTSyWM2B6cQXE8Mm/U6oyraXgYwyMkxdOIp
tpYwP7BEVHnt3/lonVjbskaVkWjWU+flCgHKBSHd6o12NDbN6gtYHyf3IU8hqLCd
3B4RLaqXiUP0XeFXmmi2NnA/nR9YaILFw4YaI+FG7b7Gbt3eMF5fimvesEvUMo62
daVaFhWH0Mear8DbkqZNI8CCgC/KK17lI6QaYUt/y8Kdt5s9hFyw+nEleAc/zddz
rtOn8tdktmketZTnDuOB9eJxMqUZJym5jtKehzRXr2knZPOAzIELUhVsB+Xh4v9U
8ueIABe+ZiYfBXg5MxPDz3cm46D7nhRRxqaer9/uVDJW+LqctqbKXNjMjL+4U5MG
aATeDCeWYYQF+f546CrbwnyxVJ7bDWOQoiRB6ajZf11cDL6Srj+P22KNy7lb0RPM
FdHOV2DniaJFPT/jyOiHa17SSHitIx8deO6ZOBVopWPN1p+cbIrDquLm0nhwlibr
tSIeHR3yMjHuLIf/i7WnpJEEi0jtPiKPI5KQnozA1mJCgj+98+cRsEwUp3Qkzu3F
W55+ejschAXCFJxjt8Y5vHk9tHiQvB7/VEuTkWQU273M9tjSMQoWyWv5RgIZZtvy
zRN6r7Brv6J2a+mlngHkpfHelxZFfWgkGGfj1byX2DC+ijogpn4oR/iwYlGh/JBx
Thh7hHwxhe64KdtnTSt0pgMW5TQfUcyfdtJkwu3p7zhLU0gIpYnes7/RLj2xb7nB
uenZNiZpn0BOgyfc2U1lCQVY+90e8RN6i3d90ocu1bJE7HVeIrR6XDOlV1AuCbAD
Orzgl87Uatsike3YJH3MBRMy7UaVSQwkUPJc/1btepod5M/CDEVBsy0qaA5mPm3i
E9SNjhQtMaV/dmli7OA0St4x9bAPp82yO77e4Ehd1xZ80Tow+GgKKQyiu4HWC5Vz
wYLEYLYKe9opxTCme8iFicO5IUM+bSDhC2sm8x2RcuNI9e82kK7/lC09EMLabpm8
4YtySuR2tPyfXrmiiaQdTch8hzjnEUL3BEM3cwlUG1YK+jFZhDSHNUHdxMIa9xI1
Ho3dQ+oI/fUoY1iHFPnQRTwBmR0ZN0yynkdcY7ZLxVR36DsLqqUE1cJ6T475YI7d
5dSfYU2k9MxYRwbKFp2LRonJjZPh6XfafKpPwZt/sy+lplXxFXe+9fOk6PIpxR37
b849u9xzmjIiosQu5uDICj1I8bXQYYg4ROhR7O3KSn9s+h0imzt8Qqzv/RkHS8wr
VM4FaYx0j9YTP33/WwWOcYnA+pspNBEBweQrxVf2S2FL2wvuNFVdLU+XhSlDh+TG
AEIKkKIQ9MmzmiwNI34Fvi/C+z+hLxdv5gcM7k4hX5hwd7MwXUyEEKIsnAUGopuH
p7daafPXiP9rv7DPvOenZBIIB1sMEQPBFzFnOTW1z55kzGZPn4QAnvTHvzoZWATN
YvKPa+lf7HCKCcFy+43CHOJPlLOB0XNYmeerMIYatyelv1BoS8WTaSpgUhoe1Lrv
qfwhXi7ZJPWkd1vKBctv4Lw1SS2o1xLS4PQulQyo0Av+wrrVG9JpHoGKrRSk6iJr
a7we8Q8dqoL/oX69bfGcchD4tY132weSRPPaSDSGZbk33EMuzQNeHHJLGnRFfDVF
fpMX5X1M36tUjczAkqvkJsvqKa4swnO1ZmMpB9oQYrUz+MHB0QWlOROkomZgF719
bJ5t7Nye5w10JkElk/RJA/WMPoFMVJ1QgyrRcK1Quc7H9vANHM1SJmHsfkcHmSLI
lW3ZztOmtCdPgjawBTs5fMXjx4+CFgZUICcvcjLRqugCrT4/J/Gcohs92hiHtpXi
hx6oeAZ65lP0sJ3drZvPnifGytjHE/PtCn7dfieg75wWZYb2muCmbHSlIja0rl6t
eop4j+NAygFIEihYx1P54HenENj2KzzGTTYEqkb23pKfUa4Qjtbp2RAnWNAcLndX
GjLTpqsOPfPZHvs4pwIQKVZdY0y4TkXLYhPnA2XSxHTt2KtMsWHLecv/E/Lgbe13
LCazUqFlzjPnnGLvv8gdnKmvfB3aV7wqpBPnTuUWKgswUP8XykbIbwDrROAR5JIP
a8gWK1wzLp7/9YFKb5+I7px06aI4vCY/PK9H+DTnPVTa2j2+P/wJrfVZPAom270P
biYhXhah57x5+puMkXTntf8AKDzzuW6931RfCKpEvYB+Pi91YagptfCB/WIyNAgy
HDgME5KEDZ6nDL4S5wV+H6JmF5Li/G3bAyinB4iKZM32QPrC+t4IzwLWal213ZZu
4g4tQ5/FHN9LkMJlPQdK7adqM/7b/pM1wwNIB/89OzrPr6XPpebdW8XdwWlV7awM
Wh/7QXahDSxqEEEUNv2QeugIC8YLk73x6IvL78ryzVel3LP2st1sD2I5HQ7nzze8
HJlsO15/dz8+DGfVahWmKqKATD3unfP3DqFaOsnSJyS5Yq+5JaclwZwo+qAt96br
j3IVoUiP9tYgLMO8dvR86hXSrNmtYxfH7c25p2WQeVq/SGD3K695efnkYog/Jr3O
svAFbVlHtZNDw1sf/s2A0kJxigfmRpTTQwx+OqJdneWmrESD1xQGFy6KDKIyRioR
92sAO36oMQlYKmjn/eZIf3B0exO7tWSupGnwmPsVmylLD/Yx5MLUTArSUB6qkS/D
Tmes+y1dNK+C9FPepGtT7XFwBZHNQ7m8ld6eWYY7mjWhC0dYhJ/+Wvynt69d0t+3
yYeBu5ZulWk/9l8s0Iwc5aCuQY8x6HeiMCrK3KLbLvUIcgTSy2tKQMnI55ZZNjjh
smwEDViy8E7jGgqZjRUlpHz1gyQ39BYcWMkHot6cVcwxCFqYtTqoEUN29RzmTx3n
0V8ouKDqmIjVTK693b6Ysvgluc5uS8OJafpQP2KspiriBjl5wg0Kh8ukXyCVsUMN
pk4RA4/CFKyMskbB101eWiuyRTUcFXp9ZfqdVE/ms8BRCy+pMIzbHQ5wgurK8p4h
LmI71rB8MSe2ZixDW1TG3nX/CETrWh1jqMaHMRUqFQH6eGPBYiLvxMD2w6yz4w//
3I8tV5Ar6iCEooqvevNt9y1SplDrY/1dM6ViFO7KlNoBRV4C2A8RX8FynKjzARlB
TuT03XwOinLeYtAvUSdAYXw3YHQ3oLPllrNJZAP4F0cXlZTu8NG/06lvnnjG6vNf
WEXNb3/vBTapRHrXz/Sg6AIiJRJ2lkp3wTEnDi/xow5JgADeZSg56YkW17VnnzFM
mRJ169zSg01e2NRjw29jdPhf9bOAeNvTdrKafgow61lbWGEF0QMj1YAmt/5mSaom
JyFa3tceDzrDlI+nxFnl2Zn/zhq7jhOnrt2F/XgP7TJNVxepiZV+y386S+6hrCmw
AfxRSZJD+5EUdmL3JEV+2z5P1ujY3TFiYJ2367QIEz0mEKmYtojsQ6EH+0BLchki
wNIyoIJNyAj+soLK1cau5iUcSXt5W4ScEo41P+ks9W2nrAwqyrducoXEqVdxko8i
FSk+cg2Gy1Ka3XonrY4zk8R/2oUOPoyDiP/sYJavu1a9xjH2g6haKxk7P2mlYGme
lwXnGCcbbP48wvA+xXgpju41hwwefWRDNkALB4kpfe2GHo/dqkjcV+a+3PQvgDQc
ckE7hmvAh6b3d0A2rxPFCWXSRZoHxnuW+RBuGQqjJVcfj9bZxeKNWJOhxK93wpik
ohPzm148bxGzVpOEmztiWgit0z/VWsVf/y3oQrfXwV8uEVw87KCj4FHjPb0+sOgQ
APZfsR5Xs7tLiZE1DlRHQZyC6GrWadi04CpVi354Yqxm9uwualquVuESc12ia+f1
NRwC+TJTTiQx3D51O7CVXcAE45Sz336FegWUE/SvRj8dyN2PCdj30h7kFk6ImSeZ
DSxrqytMLN5Ms+OIm8b5hflpYvxzeHtcqWWwcgdq02JRDjfS7i4LIjQ57KvmTvlS
86LrD7W7yngEmCRliMEKK2aNQhlDLUADUb+jWRNtBE+jEV0Vrn0MaIjMUYxQtbs6
rqJCNjlQn+V6mrKr4FZyQhL93ATR+dzGdYsmoRuxMjAc9dKev0j5sY4FJQylVol8
ChV5ISX82biNovTmshQHlBLZkSvNJk/1gcy8aLmbJ6Hj1TOjaZKpe3gRryHEFwQW
l1DrDy2PC2AmQzASM6LmT2YTiPNCHkL2gxnbPcm6YQyyincr4l4z/Ck5sQTowgK/
FFAKaB+LyKuzAf3rfPsdmv52RiWPcrx1zzwf9Sv7HKSrlmMM8u3TVQAB3WqUVJph
Em0VVprdWkh39TCh7qaLkAETn2nquL9pvLyfimcCTe2Ddb77QCZy8T3LvBZ+LGGn
SwKegJqmkG0najUWDueO5AETUudkib2O3vOjKaVsNynh2LcXHVFessEFpOkuQCzW
xGP+hkjktMCYdwGof5+oZouW4vj35biPeNrSddEpMtACiuTBVwnzgY10e/Gg9tlK
eXNc88xl1KScbw5rPrP3xtJuBRDKEjrbV1lpUkcGBc3/yyot/AvJz8PcahYb8Xbg
FWPkwW2QgIQHPjFAzHnazliVbc1XKc2GaEentkZW00kdOqq5DU4vQa/se3KXM0sV
yBJl0UR8l+5ef43AF/kRBG1fxMManWB4AxWWCfcNBSxgeo+kgUM+sHjsL8GA9zHe
wn9h+4UdTI/qA5yUPm/6A6CZiA0x1yRikhQOLFZRYdg1cCf0KvTVF6p4fD+alXCL
pU7lfXn4jMBp91inBYnkFsspo87uXFpLBjMTkQYRTCoubWtIwv2f9eTmNP62piGw
ew2Ax6jB7RoXbHUJA85DLt1LFWWckTL9LlChFbXlpiRodBWXU9F3VZI+gZluRm5+
anVgpSEcyomjBCVR95FJvknP+nsfeLfrjtjhqUCg9UqlMnvpWo4dV0e+a2tddEui
b/2SPGT6qOyeC155bStYQ06UvSthHYcNXhia+9Dxi5CGg3mhMJDa/7a4C3NpCn9M
ZHIMpg+KTu4b3XCp2Yp5iyX6UvDOm1izDyIQV2+gTBF+RK6L5vPO+1JotP/IoD9i
m7F84vX4GO0PSIhAJpuxHAFmcKkDYsMCz+OYz5mMGEVx3lmZ9N03puETYyUyjcBS
yd2GIGb0Mms4t2oIfPf4sgFdJGR9cq5UZTqaXMOo/QbLHErNyrCYk6L4fvOk17/I
ccnpHIkKiffGPQYakUbHM0PqRoViaNWPWP7kEh2TUC0F96WEWymBCDp64D4Qk4v4
Rqc4cLdvfB6LuppauzF511nQEV3YmYb6l05QLJfM5SzezexZXDghEmNG+xeyQkBN
sWU2g7ULQvyHxbaCLAiMSCDUTACnb0zGOwFUXdKjxkEz12IATHmW2ZcuNhoPdhEf
IDp/r6tFbOI+tHG4vc3yDTKXMmzHU4Fkh30f+KIOdlmTt7YQQyZpxXACXZWa6GgE
D9+d/HWWxz/7FiRN13/L85KjQRqhLNFD7IaTTErCDBXNR/RdQyLSn9nHBY7leg6Y
527NW7CpzPEU3bt6JklpnnOGt6vCMOjwFFyo6GZ5QPC2ktY5SmWLA5KJ5zO2RevS
EdqkdRZbvpGiEnePvNZXKcF4C43mJrKPLwbmVK4x9i04mIZC1v/l/vqV3J3cMxhO
IX8i/c7yDh6tLJe1pfivJzcGgzgR4e0rafRHcSAsqEJMIxT8ds9eRdfnvEIZaCkP
4Oar8JPF/Jlo917WR69xVT6cObPpzhRPLI7XtO3rdi/bOOdlR+T3+0D+fGWtaqFc
TznaQXQqCZcOvrqhwELcFG7j+kOd9v/f/lCOu1Vx01FyIib4BJ/u9F0UdUvoZ1m9
38rJ1Pv1HyDpsjJUFg8bdcZHZdfTI8f3+BnzW6Sl8swWVbcLki7/QeuSDv3KWxJS
N92HONx+WixHHypXLL7hbX7zNXrx844fNAMt/as4oARfzepFBaD09QZWm2sPUtV6
r+mb5Z3eSjnYY7e/fdG2PgdzwWB+1c/PZ0jQevrMYno/8p9qOwKg1qQ///T1hAb0
er7Ol3AGLchaxNvYT1Ms2aboRu4hTPenMuB7UEPjrKfNmSbJ0Gmv61BzDb3UUPTx
MD8EXoKtmkNbny/KPU95mP/Rk7uZGqlCJFTLiNEelZ8QBIlzYctrmWpck54VJ/Of
KqePK55KvNmsnp83S5OgpmjVlSkwTMFIBqR4XKoDMcOgwIja4G4ZzKZDWxBoUuVU
qJu5dgdEuj4EYPq5EaEK3n/ZoUzVkPuYju1V/uywrcFQAe47Zh6wddl5gREsb5uA
gvhkpA3TtE3g9Puz4r0pt6ny+jaLejux8FvgmSnfCouLmSaxAfeGIDDVu9Wld4di
pbSyNk0gcsODQikB5soA8HaP+0ZgLACzk6ZNmy3xCCimGJRf5psXpkIbLfaPHZBm
cVOfr1tOVOcQ8B1B0WFZyQlRSk91rk2IqxQE280u7z6l7rV+SxwIkWzpEpTOEd3D
YVldLIrGO5ii8Khn1/tTNNkMDW2UcLMvqxVqwbKHXlw2pmSFx0QyDCfgkzgd/oTx
uufzj/75wa50G2sUdinJJ2raMMg/alCLRgfAXjNumWJzIDrfnrhnHXvPKXxLZP8C
NudKNDqsrDI9fND8yMyAGYwYdEcVmIaT+ypZ587qWBfSQOt2Ut2THsQE9m8fKQdv
Nv3D/5G8cs+rFd95rQo44/L5OfyWXWpXtPyIfGoiVcFsj4NEmth71yUKRLK5TDBv
0pLT4W/u2UJxwp9w1v/BbHJ+MzYVPLxT0pXfIiFK+hDpe/BbHfjibckvUCM0gX54
HCJeAFj+181EJPxevCa029aPlKaCX53Cz7a8JfJzZVnu56nTAUYwiww9H0UVPoq0
zDTetrbKtCAya2FMe32E62pDEEk0ZnUWVax9wjh1l0J6Zb1DgA6ycCvgoqNsFwEJ
8X06iqk27yYMTsUaKJW8MvlpF7szgQOmQ7XtGezHM5ATYzasz9k5SjMH49srq+Iv
1k+f50D5EvtEuaM8cFKGpRXN+vdgTNGq2hGuZnwpvWuLYtWEbQRvVgddGPgeRQ9w
8U20TynD31BgTDlcMziRWe6vfCgUSikmf3Us4X8GKa3w67NyHz/bHN194akO+md4
jzyBzN64k2sBJpvyebGYZjDbxF+odDkZqBLeON5ho6xm/7AQzoZJOFsjjVsf/CFp
ohb2wqdQJBwd827m1kWFaSMMEKuOvlT3ZSTHXzwqLvwiCpqRqBGCvFvZXNyH86xb
b4ZB8/h9+tQvHCRg+LgCU1ra8UpdL0G2TGrd65XonB87ftrAueSmIRmAvSOrlQsd
KFa6BT+zdnQBNEfCyX8H0kIUbu7v/llJcPv6tPlcj6di1Tn+oabrMSHnhuWdtDp7
Gv7cS12vD/vvNbshl3XzL0VUVizWaxy2mWT99NsRcUuFCp4BGsq/CdzhVlwvJKO4
lDky0FSad6TFjzfrlYEh60WNAPV9B55LXiZ4nDxRB7oFj40kFnTe355doXxPN+lu
rv0b6IgUEVgD/rqKK6wejnilL3ZiHuqLjioKqLqFZPJA8nJyndauDndBFSxZbBZw
RCZUeVgdTaPbm85t7yKxPaGA/7b8kcjrkLh6jFRVkUkQ8iIk1nNGaDfUINeHiid3
f3rH+xstud8sl9U/6DQKHzoPSqDVOjDa4xScxQ207vB8HeXT13IFg+Z882+W7sEx
X0DqPhD23vivyGNIDt6z0UPpjQrabhzGFA3P1iAnuJScSek1T3P0sRcqnPBD5v7T
ig+5jw/cHhekl7vUW0RtHf76DgetzVH2li6N+2efrdImDr/cMEee77uzkb4LLNf1
IZd/4O3Q0q8yYPLCWaAAOuiHN/9MPJjjoq6cdTzU6ArYM218p0FrjuTkQYZsgaGB
Nj7shsAaE8MQlqQzHwvWwcIzmJ9TSG7NHks0RGE9abyLs0YUxSfBPzAqL/hN96Cf
mHsx90Ixb84xCkb3g867TXgntFStUq74P3fKa/arNPtvzYsel55dPdeIqv1LzM/m
avTOrK+rMZFLtAhDFNWaI9yWAAP/BaIuiWMinwTx0uqCJjhqzMFTlrAny9Zu7ZcQ
beLcAV5xUs1het/9BS+z2/0I4BPW3eYeYThtR0hv083HQLyfpNky92DM/k8Xq1lR
VQdWd8Nh+IUW5YqLbwHeooczP+EHOhLqzdyhr8JCuEc393RK1RYYgZVgg+eh6J/l
fsjDRMA9zR0vCRISHTWyPuKvyw/fcOJpiWnaUf+XnKwd86cTVkgwK4x1KWYvER5V
fbepb5hmaICEwinBf/FRsYitnaOoKJ1Xng5cDEl1l8KyYroI6GnDe7accuk3BwiV
taOXUAk6CtqGTEmWPq+KDwtzyjeFTr9kiH4YQ0kActSh1326uQGlgvWTg4Ckje9i
zv94KQL4ZwTyZE2RuxqKWxQAiBrwDtjOQq0RCjYPzJU+y/ozmsfQ/jPawmcuv+Yp
EUPEQJ1/R5UxOWeUivRG4051ak5o/ejgZKlgjDcv10WJFVdDWcca8X8+m6TPT50I
sZm0Sjis0GGiM9nEJr0rhnafDUNDTmYt4keFiJgUvZI8OPEGw0CcJn4dlSs4DSX2
CdI+3vkhhhubhO08LEIrPkRoWALTcddRD+3Acc5Ds0Na8k8qDyaM8lig34+mriNp
lJGSKN4620ShqW3Q0T+uu5tHJ8wfaXz63NWyCWrhvzN5hRM/L6dww5iopKASemvO
KAP10fEaZRo8EeD4qRuek+unjGyXxyrc0aoK3xdXq2zftNYlHyIVC+dVm2MorHQj
t2/PMJ9xFrY4rtYAW3COzSNqnQIvtqd+aN9HLj8Sc2p6haJpSsYMe5q9arqUHA/L
oIIv6WVFe+otfjBCMQnh1siqBuFbV23O5aUK45WvArrj2xE7+GMbfU200OS4dOqi
gGeLVH+JrAQk/+NHqw8emNS8aaCGVZPUay92g/l1bggzKmJIormpVFH703aHw3Ws
xIzSyOM/iol+Nqhk8jVKcx2J8WFXGdiJJ1nl3mnFv6obOcXUohBLd9GoCOtI7LqS
YEQ7wp96Ut37gopUg/Bzr6zb4cFpQe2nuPUzlxFmNL/WZqHdAALGVpDmZJVv5lOe
aBQkSrqL6nr5wQAq4f4DVa1bTDi4qT2DGVWDlmiftiKh7zH3oH+je3eFLIPnTCR8
Hlh23xvTD3/wYvA3/gDABR0xTWK+RpbGlW4/qPGQtglKc2ZTYFvkF4vjA/ic5IH4
BiXE2V0AOtVuta/ReRGn/u40321HETFfUn6qEVLCbGQdh604xoDSg0AgwiWRYai6
lO/GcewMnI357h6iFdYvFd3yZNkmdfezwQAokj2S4mU2UfWZWIpXUJnfr3c80/g9
PBCXFrL1fP2lA9pOHtE9sK4VOGg/07dzVp7IP8J+k0n1RY4Vswu4Y/oDTrJ/fmyf
6sEtNNAh6+tK4N5KsJQLLsL9KfEn/nm4eHPiZuVgay1WdTLOI69YSP+oz6bXdGpD
4f3qoMCFLbIQH+qBXxfqoDE6H5CcEa4HyxsOvpWEma4mN+uXl+vMIbv694t/OAM0
k0MEQ44HDcrfTEzbZiwBCMWH5eArDqR06sp3By6TegTDbWS/hljv0BtKK9f1S9s8
mQxe5bVT0ziCJnV/j3HmWlcB2/NBIMDoE+eb0SQtn3JN5erKfOEvKk26DD1a1fTQ
6cROLUFkY7r9VZDGfiDqYVxyPX8tMzJAZSfkiHbd9lp6d8ONSGlNwWcQr+kQ3NoR
aywYUr5gXeY9y0FD0pEkKG9hSchFcslmyKq4iKWKLz1RV+fHl8oZMhOQlekLXG8f
rMneTDwqzAjcmsDkYeWcifyKN9BZHEu66OIIzKo3tqHy1+w5iqbyNKThChOMpMjg
ctkNE3ARqnQXD5+4ymMRTHAOtYYrluGmntf88CG1DXziV9kBlyuJMIxvIGUrvcdj
gi/K1U3rlhaeMCSlyXCrAT4BW0HKZPti1INDW9ftAQ5kboV6kbL0l30Sg9w6ucon
N58upzgqYaB6vqplZeCPFsNzGpkcivthGHWLvU4hc37b/T+wWvo2QBsEwwYM4Wdn
4r2J3NJG/3JSDgTorsb4/MDo3HcXAktd1p3//KidvLouO2BANjQ4pmfO3QxL2bIT
k9Xod+M73gbU4UfsLOoqsYASlOfLPe8950ya8V/NNsVPnB+zuqKaNjPEGiuAbHsO
8ubxzqczRfFnwey2g5qP4giVCVLFknwPr+E252ZtFy/CO3jvW+rgc0TNR561rdmI
RTugEkvAxa5R+IiZfC8Hpmz304ht3zY/HbNkGinlVvmOtaZ8bFxyWJ8zyAKs4xMR
StxbbXm65YkYPamvjDSrBX184RuzhImoc+REFbxUJuYwvpPaHGb5rEwwcR2kDp7g
37T4+NMhzxryMthXUEomWLN9NmLBPmA1vYdxHvUQwmhShmx5SGMoKwJZ+JSt5QCh
ju6JovaVFRnc11E3QFaWAWrS1VyKhS1Qobh49AMozkUB9f1jq1wNSNZJCDztrc4Q
O1AZ2qv0V0lo+odkpQ/rQ3PAMopdVc5BHjC8zACb371u57PoByFDU2DGQ9e8HaY7
a9MkSws4Qdq7ZWa8lUlDt8hqUdiZ3cne9A6pzizsLmMEmrjWnYzWr2GmIMqSGxx8
WkBkWh/qz7+/ntyL2U/qQqKgMb6U1OH9qP3OS1spB5eTBU/HDJPM7yOqLpvS5wRt
P6/Dfx8bPAp5EXyjV3O/FU+vc/j7otQ0wV9rYuT+B57TNdqTHREeEhc4LA2TCy/m
V3GkLrSZe69fTm7gJaEQImcCb+GrS0VXnir5gIAePmhNnCqsElYGBZqZhuOwSFjP
zrPhZrSyv87Sy6Azvfvq4YU2lYBp8nGFWpqq6LSbajhEwmcZ69n1w2AsaFtBMfOM
PaDZx/piCmIsbnT49ctegoaE518IUR7VvE8UliY8Ce+Qo/jc8pjsTOJrqV0OlXrg
vEJVrWYj71igaqysOq0DaSGeBtKtGaZu1tDGA5/6oej7rs1vZUkNukQKAOsamR8T
O0ccJsCRm5Ome7UR5XWzdiEw9SxYZ/P/HO9k/ZJqxcv6SI4Ribwfjia59N2tEMwZ
rJS+DvCo66Uu/6yHBUwwD0y7/1jh8KO47yG1FsdPGFSRc+TCNkVfBxwBsWA5ZlUN
dp0c7MRJRODDPBq8MGWIn820dqIyxCYomwudSgXDRDcHVNh+ObL/RMBrlH++52LN
LKZZyhAhFNxv7h+fURx/xZvpKE5Khev1jVX379DFq/wBzeMS3Kfe6+ADrlosz6ei
VVT1gg/6opb9A5zFj0ZK+5AMgibd3MNeja0tF3X0Nvvv4IkrlWC4POd0daOy6uoK
o77Jd+Sh1KHrldWT2WIo1dZzM6SzOSkDItzVF+vXEkMA+FLP4OKEE3XBvl2BRafI
nBHHm6+cs7QGaHBsz3EPa3R8uMNBI3zfxH3iFziwiBEzMkjd8Vdm22BOqsU2c5ef
9rSf8sHd2Uu9YE2k1Qz6FewYk+lzVXi5R1U7AMTVCkCz3CMzr4zIjG3MM0F+bl4a
5gjECl2jG5DxHzhBu4DJvi/UlS8nxgLQ/0IYmdN9sivHJgB58uDKxf9Qm48s1lR+
vuCDaZN0IaZ+8dQaV/2Oax9bl6xsVCq8SMRwG+IGRiBX3ZreuAX8mtUJAFH79Qxl
Io86Cszw0Oue9NIaZjXdCDuYO84hJzAI7taBfUpqDoDGwD0dqDqarodh46CDGJc2
eFPfvCbXhuxvkVmeYeq4kJKMrsp+nDVeYZqw9ydwfGd9TpwElnM+N0IMk04F8B6w
tBh/Af5hN3KjDf4Q0s4pRbPN43/Lm9h/91mPH95/XC9uSHuMKRxXpB0+1ttXuGlx
RCf15xdHeYghv2d7a8TJwcbpQR1wQW3odJbxIte6pibeKDfTWZxaswm/jACsm229
8HCqoSEJJWo8mfA26ro2x26IUCnx3J9G8itumfp+C9isDjN0p9dEYozVbl3nCjmf
GUmEYdA13zCUemRV53J+pH3U7c0I2Hr+YEwnmm+qjvjKT6JjZVVf6QS9JgVmtQ53
OuJ33WBB7uwefl3R3Xh0IhTpkQdPG36r6bEoUnkY7lGNXsrPzzaG/h6JSnUJh5Lu
OzHhy5K+Ot1bfH46VWHh7Xyu5k50i8lESNAOunKTke3KKg0UMaUhtq7cC8RPZXOP
FtxCYR4jfI3Nz+qqtvIywwv5mYuomINWdUq20xa1hsq0ZKXofVlIEArxmTJI1r4y
29E4pXYOWvbXqOcEEMrYvndmA3ImxKhbA9a5eGTpfIQqTlU/wYdoZR+gyZT3SLYv
iO4Yok4Xs56DgC23Om/Oyp4Y+b1DHbu+frvtg9YygY5EFPXXKALPWz6oa9J3Kf8K
YPAJBGH3rFtioiY5LDuT33qTTHa6anYn+cMXRGJWnFQK5oJuHheZ1VgPUrs10ZbC
uPRVT8VusDQ/D4DBEhf4cpGkEQdwwi4FANjqRPfJ5Q6VHNDc/KGww+72i5hs194s
35rMkeoTR2ZHw6/Z/L/JDIalwkIRRBTEiINoRx/IyjztFmqscj/5ZiE3j4PB+46o
Qo8VR/lGxgIPLUVwvnUAj/gOloKUpcGO9aBbs7r3FvF6F6Flj/3aQlOfdVhi9Q1y
385qBo7/CGwS+2K6H3jgfDrTpVzemhftdm6kO6j2gc0HV0UuXUSE3HorqYCWsQ4X
eKEqaOrFtXyZqB1U5pqer0wlgGAa78Xtad6FJogniIBXnbnFImTfnwu1sZmVGVFb
oJ7BwTeI7i/WThsEc5H/+fVEmMoCo87kit1NFm/hi34TH2pxsw3fZ04CqZxATzBO
r0i0nWPAcCVjyGvpA9PRXHc3wP5eBzuia4OE5/AHrod5fhBIdVxwg4WoO4KS/60w
i0Mt9Ui8sPxh2uT4RJPvYIicyXQt321qQIMhzdpvHGZ+lz7R+P+Hnpi/1PhEqrVu
vK1UcmsBcnuQ+zmuTOYE9YU3CIdUMasoDCNqy090dmZk3+ts+/PNXns1k++20/hn
8ZLFHRZRt9vaM6EoYYIxnLLWUbgjyNzSOmqRgITkeiR5gHaH2N+fI6NeUDpFjnL8
NCseonDU1FlZktK8uV6fYwDSC5sTNb4sWuNqNmnWaC8eMP3XrpLgax5uMLCI5xj8
kep9KQLseEfl3T/5x1UU/OTACFZM0ChvNIJ/yJacUW7UIN9Yygn3H9FdMcyjSOan
/WDBG6vtlRDxd6Bvn3H5kqkaRpMREMIcm0IP4AcMFp6yfN6dJJbywA+6M66Rg+Di
LeLpgEETBnG45KGvgyImGfhNUXk6BKElYHmczdFT4VVMSxOUnFOruliszhF3i9sf
yJEmXN3QndfcF3DFIQE3d5f8sW1Bc5doje5RNKiYiQkKcskadzq3nLgtc5DVpncC
nST7EQLHz2JHXYpk8WyAdpG21ghBO2PHBMxAYK/zHBalPINXHzWSxdyoBckFctE1
H5RkXL8VaREsKMVCDi+qkxBwz5HN7G55uXYfquCBbPUSnLaokHZC5U/DWUATO7DI
UIPLz+GWfI2vH9gVd3p9uFdJrnoLDU62u+afDCFiP7bofelK6utrztIULi7S8yfG
vZIfM9R+ZUy/fLaoiljlPQ5bLY4TcLZBMJ/Tnkt/zE512JsdkRiJc41ZDiCwOM/H
HOC0hMkK6ntqbbYxqXtj3GPk2ENn16BxdDL6zrYwMWgmhnE6VK8xImYmz0wnFDl9
8W18kpJNncIFi7REMw9tQE/JEzY0ok7t1tkDE75WTgWGHeA8iV3O9WyhIhGdikNU
zltPhvExsYAbppBjz0i+Qqav/iStAuS0Dh9VEJMWgRidLOu8HblTLesdswZEcXEV
9s4VkO3/5zTRPJsiLSxv/nUkfEp3nMXt9rP7OQtmgscY7xg/ni3dX5WpPnDnHc58
t39BbllU8kumtsdZxuQEvW+Cw7hzpNhaEgk86E76DJnZ5k7360iM4RzhzAFevsng
F4ZrAqK0tNLhXzO6rQLU/g8+N5j5mOF6Gjr/jsFz5A6+daMrArg37klhn5DFudFd
p0D+P9+jDWhElO2IMpWVG8rPEg9x64+POKzDz0zIsMAmlS5TJdjax7TXzZxjlhoD
QoK4YfSyA8vn6D6/E9WiUUqALi8cCFzGwLhSOVq10yhakvZQo1VpuM58DeiZQKF4
siGPRcoGlCLQoMoRH1eiZHThcCIoXaCJRKvYHt//RWw6wUX/eDBd27PKr4xQFCc0
9AHDJpsWDuGpZad5OExr66eDvSH1NCz3MHXOAPnOI58McGQuBXu+ZwlDI8XTHDcN
cXrADYM47PVztzLWQzpdGEm4ygneC99jjY5CBFd25l7HTRyjR5gtnCNYpOENAvUL
HqZ6cgNE6grJTnEIVP4C/qbhGyz1gYWKZ3WkmsZjgDUZRsuohJwJ7tP+1S2aA54q
aSiJ95SP4kzVbNSRJDGUq9VpWFyVvCXl2rOI7qBSG5OFfeosWiSM4lRhSYpHHs5Q
wvo7xVOk5VGxVbpk4fkkHa75q1KG7NVRlzLYyLB1j0LtHb4qM1RRuRfi4XVAlStl
dO0OfD5GU95bBpnp5BXRCcJy35ccz+EhIXpX7OX9C+/ApQVMExwaCbRFaWZyX2pt
6gRlBShyoitUFKsRqyxP3Yu0ueydSKQbfbjSiSd9fH4V7RoQAQVf7gt50GlxurAQ
2yroqAf+rzJJtzMdyyU3decCRs7hXw+0pXS6b/qUGl0YEomf9k22EJ4kBxVkGIxT
F7Wzph4qFoSEtIuLcnV/H1GUPWVMwkl4NJrUgMOAk+DxKwesLRl+uWdq4gs8EWXo
QU78l9ZJacAtP+SIPJv/bf7+StlB+fYORoR2Cw8cd/pM+0NwJwNNU19c6JEObSjE
FdFS6CIDzkzhHUNUI/YxHN5wtv7IrrI/0MzuNYVJhjG9q9M94GmZds2tZeUNZlzB
CfbhYK3GghQfxu/r4YU1M3u7+M3wAFQcXx4eSYkccyQD8swrztla5jWA1Ge81Vqh
aZ1UfQ+Zl8oE7vYJFeP7Xnrp11A0ZgrCLT2Z8AxJ9JsrGuSaynOf6E834u6bX6CS
aXgEZ9Yb4TICeyeYHQ3tpL3z3LWXYCRhaczlMAWsCywBO5rW2YVAE4DQj4DJp04f
FC/PV3dn5m+m6JZwsf1dHpX865xwUAJ3o2uH+IktPUu0KnlMp9hk/iosk2AOPyV2
AQSVmvt526hzKIHFYd9Qnuo4tE2DpOB8k4lwNxA36Hg6mQ1TKJ0BHdSukhFZIk9N
dCZD+VGvhP7ikKdQ0oNrs+93YFNMVwzurucawcY5NPO29Q5mToUiuWy5J5Llmr5S
72/k02Z7bTuk/LHgYtlDJ+dspnLR85g1YLqZrnZivuU4v3nS3wkn1dR26xRDBfXk
1IUjCaVUcMX6mSc9XpAjxhJTdGnoFs2cpmTNx1+l+/28k99X/cDtr2FNS1LaVQQ6
UZb5CHrVSMREZXNSOmt73QgAzKC37tA0ApZSUsORrGAKYsN3FlmcrNOff/R6bHkl
7ENrFI8gLKec84DsRET+fHkTJWAjDvods+5p/N/uZzyt/LQmMKDeMVC39MXE3CLr
XK7keInXmIVEVub93GxptcobpSXBgDzkkFvPgM+XjZeMDFqWV+xxKfdzSWpWEzD6
q11jH9WwDQcoIbiAkKk0A8rWPMyePRimpU4zxkMFiQswCUupZ0yF1EraUYqn03LT
6L1C0oXnFLjuEwdpUQI6IxD8n6y9xdmGSFfQWhFVKcfCuTArjqujy/quH00XHrfs
UKiiujkZMMYXU7eM3HIlfJDqTiLZcIO+47xlXDKFhwpolqi2tcf2sw6lCdMyVaMn
Bv2Q0t704JOzUjfp3A+w2frVjnt+QTfXMygblsKjE77/IBIIWak4PYQ60R0dL0Ho
bnCJ6q2MTeOZJ4+zpWs/9e9J+OvtVG9yK9AnemZETvg8DEABPBiFKBFYVHDtpBiy
LPr0nOFSMZbxllC6jplsioAjXGerE+zMVb7eTfHTzJgS0J0ec9T/86+W1nGW3el6
J9u3l6Rk6a5Ch1M3FKhuoKkoM4fkllkeStwYusWt7Vn+t9og/VqM9s1xPbwHwYgj
lS59Sr96L/PRhZHPNijtNekjpHW6QnnFJnJOcvr+cTOvPdDbXaKC2uZOmZf3pTZZ
AlZTaPykXFi8+TpMBlfwd3kEiWw7nObD/qcd12jCxenLGMmMPNWe6BYmcLTtjPVG
3GHKcibr0l64L8dm+YPs0wSoirpPuHVkLlGgPRavW3YWlePxmsfsPaOAfXHZRn2y
bC1P9UVV7cBmsQlm90sfjyL4SIWR6QUtTlX4HD7vSSsDw2pEW7hELoba290Zvdkz
4p4h+K4/TXak50lFhwaZP6eDPNFfw+0JmeYVRFoAfIZA68DBNfYT06i23097T8E/
75T2fMyucYRg0JbZEqzIn7i43yPU6roH1lafYeKixK6Nl5QGYb7FgxUnjs2zz4lW
Lw1Tl25Lhbr3xLn8Q9D/ZCox01Gm0+Bw0QQjWurU4CaoMmK6IYQRLt4Lhu3xM6Dv
pCPRY8saWOVb6L+zvsxDMA/VVrso167O+LSdSI07VKMLg21PHDWLGe50Vm25crU+
GAXMaIHCMb26GLYLqBvkZvdAHXEEEApolmbH+Il4/cqOsm9vGWMJRB8B6H0265/9
i7FPuuH/O9TZL2G9cMIxI9eIBvjTz4k3nKPAKSWdgrn4GBVOcPZjtGCQ8FhlDOrY
i9Jgc3xvORq48kD33lET8jHeM+3uqjTNDN3GfHfCsZAmYYzetGIU+OL8UmiVFk5a
hTmnzyEmx1smSyY5xVOpXeZaKQkdplmyrifNVBfaugC3WCBqD3eLYRe9ijg243tA
eOeawCBKlnuzp4x6TI0X3egpezyhYze+LuuqfPBmomWo4eu8QZ46d3O58gHmqv/K
t6S1QD7bzUolEFkZOHUkMF8KBAn26RJ4EPIJsX+0pPz8Tp7GxaMVr+xzOnWiVoqt
qP4jxjUYw3uXkVJv65UYYjt0F0LZyE+QYc9whvB0moFz/3/4rpBsl2lsfZ44Q8bf
YA1GY6cq6+LZBlUtFF9AUUpPP/l8XzRjJATLW/AQOp2zLxHi3F+Mo3aW42fkPthR
S13BwR75B1o8KZbrNKf2WP+PPy/lejffF9Il173J6ZSSwzpoWzj+W4Maztm+VoVh
+3dMUZp5EJRu39FE/Kb6Ip9OpfCfBOFxxn4OSaGyS20TLmmYCrgrn9ABndR9uW8l
qk9WWOVH4j+hHKCMWWrDaD+BWDMIcMlTVXSasZFMkWocLDgV9H2FQgCt4eFMyeff
UZ6oBTrkt7EkU0a5LnT+sTQTsplUaASWLE767I2qbtcQitP3aIe+1LeRmeoWJj9+
cZNGZfN472MpWo5O13l5xnU07cWHI1rJ4CS2AhmbMh3gS9YqcNRSa4SxJIUFLiS1
rHVCiciqJjvliKdYKtndoD4wi17/A0IctiSeUSvWRK0trvsJ/MiKl4Kxt4GGl+zt
rtXEiF4WvAey+yWFTOod1e6JhXlHc3GgoIN5D/S1JzQXq+iWes3aagn43lxTlunj
bRwPBg5brA9+Nqnf3DJUa5yi+oi/rcR6Txky3QT7+5+hezB+XIA8SC4pRR/XV1zH
2/XTjq4m8LVlnVxwCjTlPm9AsuExhCqU22133KnsFM7tw9Z1hXDjTqil2fGqH1dt
JNWHGhSWuzX4T7kaXY3lt9/0E2vmmnh/n2QgD99j30hHEicD+w4NQyHF1RYkDBOc
2Nu346uSgWsg1U0v84eUOHP9bnfFnKfHfoUfCOAQO+1y1ZyI8DTiVGoWqO6W+wI/
DXffC2s72bdz81d9lYVtzQPLJ59ME+eoK281QExKcrf19xc5lJb8AjMF1iAZAN4+
nHHpaQUaGZt8ua9zyFwAKeKDzoKm8YxtLuaDMZTjrafi6dxxlRs/rMTt9GilgJ9G
1tvv+K2v65R/FkFqHZhQBBAvOXARnoL8Q44aZvq2h1LIy064Gai849UP8y47qCbY
LwM0ATEGNYLNPSGWYSnERDQKd7KYWAApdsYkfbB/jeF2OS3GTG1Nq1MBLhWMC1Dj
Hu3GDX/NzZh87hocB/kTeFFJ7SjWTQUec2+D2yekhzqXmmDT0MCc/TfPkNwZt9Lb
ixJWdkkxk4zfmSelAr02SRCPA6knCQtlUdT7nRHfmwZLGZnbA6neahjGbr+QbkrE
X+8dwYm8GUVh5UDDXv5SCWp+9UYRus6Zp6qheuCgFmaudZOy6szeBSpwXyLbyjqD
5ajMOCs+zvQD2CzyQL6XLUAd76JeOlZJS7XFIDKrVV+bQaH+4kUVipHSMy39VxoL
lS6AMLsuYNi1XSuBsEZLCq6m7XED8QnLjwB3UsgSCE6vKCZB4Cdh/XTVUHX9F0jT
oobBT47AODoAPYFOjskyL1O0P3hHOR+wwe21t4FgawGMnxnmJmi9boOrs6QdyFou
5Lv75ksoj79H6E7cDiw1wnXuNHdTiV0FBc/E9apdt2pe/7Qex2yGJwr/Po4mC285
kgJGJ+vdmwdaUrClqXpteOSumWzA0SrGMmLjpMmcvx1NldIQOyXydmbPxuW2irWR
MTT+hU9AX1gUxUgbz4wf0BuJVdSZMyOVxye32s9EyMvOoQHbnpKODg1JiK7l74u8
x2nYhV5Hy1RnnagGWsqjGXeo03QjojqO7ybNlVU8cy12x+atOZ4eEJgRCfxCckGh
HfLoBHbvutAAjDhoGZ0gXjicWAbHTQW+yAFpXV5B/IbPkBr5vTFVEwE3pgeZcEf5
JCnFthuNR1daUJBIcgeWI32aQqtpkSBjcnqX33M4DrZ8TxEW5mbuctZoQFiNgBdF
XPiLYPqRom/XqylTsEETHRapQuKPnIeNcvrJrzBQ1W7OimSr1dbWpLlgY1nAh58y
zX3M5gucqGZ+728tijtEidG2WZ37duPmQYI4pZQJaUuiQu1YRREiTqhso8hmEsHj
RgkNqdyhQZB4torTRFsFMcnw3ojfwa6YbUpRa/AMLJKKbW8EYGF8mr1MpQn0WBFr
PlUsg2lOwESMQchmV6nZyGFWUKw+fh3Tez+pGOXLDC0JLs9N/PrqfOdO+p3TWG8Q
D9f0i01nbHU2cHC4Q7/z+FY/fr4QvFPfpbtLIbXkAhqVnFNfL/mRjX60oXUWqDb6
kuiDABhTYQ71ye8CZYHtNWZGnD8I2nQbFEROqbQM0WfwLKQgJbDdYPmr4pz316au
adcrEiWz93cTUGpEttap4f1vupcmUfUlFsGieL87z7fbCD+cmRdgRODJ9dk36bRU
SM1gZJXlTm4Y3/SCqvdSw8QJl1rlLcmgln5ncT5narj/TWKYXW5tdsedusNZ/iRS
KC124qiKUvgla/iVTm5B1If7Vxgn/P3mpGd3tEBx09IzngaGn6DTF2OQAbnjNsoD
ID12No/EdBbOGVUIQaWNuO9qMThrca5EuphCpaC1ZvOxA+ZlyRAbqlJb8y+9L9zk
ZRMYv16Hpb2BTEhNcq+vF5qAJ3b4n3lYWpWNB+VbhRlCiWvXj+oE4kTMwRfdPvPA
cIOMn0rOnsFrnIyFagRu3naDFdQ2CFge/ZlsuGW+p0rSIyEONsvuz+IVMBPTnZFq
LnveGpuO3K1e0VZ4LTzHl4k0Eyj39IC2oco1jwwzyYummR87u8cv7PQbG3CuKeXI
Y5QaPgaft+A9zSRelGNMwTJ6V7IDK+1fJuTF0oFZVaBLQk07jz+x7TPHgQ69M210
Hl6pxHQDkdshmhUQWf2kVgosVPsy/9PNYb3DtuDTMDDUozW3ftPwNx3uMgOUzRgt
IQ5p/aYR5m4ZhCfVdRFgZam85CsCMng1N4x3Jzsz9JCB93pqQjy/S89zhpIHS/Rl
66kKKxnDWzNVrUuqCql4bN+iG0i7a8bqT445SwU2OVns8VVI2V21cnAc9ZwMxCv3
vUSGbyrb3SaDTXC6QOBt0f4g4nLyP5hEsBnT4quMz68b/Hz2iksKRmXfFk4Rz0+I
x6sZXGTlv9Xh+Mi41goeLfxH9PqpaKRxPbRHEOdt9oY4v8BogxbKQaIbU6V+ROVa
EZ8ZyF+u7LjeyYCuDmqlQ1VFgqN7ZG1ONKKWu4zkbfQO3QJzlLkib7MNeWbQlC9u
zsbO9IEyE6+sbdlT1Uj6kyWzG6OejVr+IXZyDIw7DRj5HVHjF063vgVju4Y9kyjR
FukprW+jaVWNmQwrxeKuQY2oYSf3uLXkoU++/5iSkO2XvIYQurLZaDuttyVzM5Gm
XUmj2mED8heqpTCzjV3N4600KJ5Q3q5SUJ5lzQukjZu4FzR1qKTtBBAmksVqSl52
nL3ubD7f0V/p3SRW38vU7M9tuRxYqJacEyVnD0aK+dFaZj4WL3Dnph2VYEfoOqia
Qyaq2SoLC0XzlIDztilkGgrGx8pd8z52OO/Rb6cXzZTpiFKcC/K6UVLKe9SjafiY
Hn1EjOr2Mn24SBOG9pP6fEZwUtgNdOWdoXkAwMUiJwYGjuJUgX33jNkOoWae5HMT
nkDKppsGXNCLEVuh16fSxDqjqpAuYRsxIBGrsb9Q/JrFCYhhbJPpFPu6gNkCNKAM
kdaAtwEfYSX50/XssqYzOsAnkY9HK4Oj8CLKsgrGKnQ1rOYeEHbeA2akKMdVWglA
pV8EpK4BoS7/xnA2JsfTGAnIYNt8MkiWdT4rtbuV77pFyTRQKkj2LdDU/kAi4FjX
3O+aPP+A0d52Fg573clc4wdKHzsJ46I6MJhW02PxpwgspeK1Zj0kAuOIz53HhWlF
z2ly8MsH1BQo02ldoXWs4gTNmWEgqDtfdndEeSTSWaJL9OE4pnu4XVBZ1DJnyWJL
DxaP/8sWfFi61eqw/QgszV42en8pnTMa39i3yDSnOelaEfqNbG6gvDm/WDZ/J8gL
I9rQi0OhlRTMKI1aMXp9Pfq/qkAWeP6YPgoG2y9+DA7bND7Mi0Fsc8Lj8GY6vaKR
wMdY495dBYD8Em8f1mn56vsR0icf8/eG+1jgCpWIdViHRvUqCQC0IZL7qBwRwvtZ
+a911by/K+pv9sI4mQZWf77ukz9q2JadI4TDflZYTCZDmRLzD2D0YXTmaSS2IVjf
yKOIngRjZ0jSs1k5vMkVcAIuwIIbnvCMuvWPPN7sSb5N/KTYlyYkgSyEz07ZRmz0
AnEd1wmK7qXde7YaeJXsh3jXYTPMXevoWIwGW/+PBKhbJG1mIuCuQp+L40zRr3Jx
YMXNrROlMtHv+OM9Y6yPg5hFVk+UuHvQDHZAUq9F9K//oS0yAD+6DUl4hirtlTii
5vkEvU8WpG6eCWXT5hAFBAn0f61RL2Dhh9qf4y3YOWpZtDXd2c1g0l3ZiHe+EQbL
OORuOnCGqLOMuBZXBMCAI/WyVQsvsTgjbCkgiqjDhC0BUMNAWH6FRTMZMSXIFoSV
7HH6TK7JkxALxpmZi5fuXlOUsMNws3xSHELWSi5cUanaI1aNEOvaJJ156aIRtQN0
WGvXDWq1u7RQt8e/Z4jFzWltRjvKQzYqNhMgOrahecLYmyUipXpfDBMz/n6v0vYm
Te8CHcS166unpg1BbkDIbzQy9eFBNim+aP/Nw/bxhDrjDOftks7BkC29uinNFpas
URWayNgzNn5S+Sf7m7TUsLRQ/aprLyfbRBRGFyrus5NYE7ol5EyblOvGNx1uNF3N
SoIZqY+HLT6G9XbpYfgJk54OvbXGywJnHbxKQyG+U/kKJ68YFvr56mSqS30Hk/FZ
wSVzNUgEUP68HVzSRNDl5ui74WkiGMQkOKk9UADCgsrdsFHsz30ib8S4HEPc3WF0
eUo6jT1YNNOBGBkiv1F7dW2bvadqxspz9Ovk6Z03PJ3WYTpYlnly1G3xZbeXErxR
HOC5ut41PcEAhHoYhvu7SVWPx/ETyLd/Qcj8Irhl62jJ8iHUgQ2xKJ4kiv/X0VTG
sGor4GQt52qNffH6/LhYPN29Dl5HqsMZL7KRZ0TV5WztSq2HgON5lZ8JUbkYG/l9
aucuNeYvTyXWwKHHTIIj/yJl0mYuJ4byEmFgZ6IbC7W7NAEsJIto9OE85pUkFLq5
5p8rncwVvpreGKqcVWKgqJywV7MvcPk+sBefsUAIo5/1cl1uILfdaGrUZ3q0vqgS
tgbC1O/wahsxPT6smGZ8TIZxkl1jd29qiWMMZRbmEYYhv1PPT6hTga9vCkPQa49w
Ah4ADiplGMrFWx6+xHgoAhyiO4VZkodZ6F209WySWTdwYJ076eMAJKhjzYfb9FP+
HbplqiAs+i/gfBNeDvH9L8eQLNzNjyALYyV+psh11sY/jH0Cw1Mpns0nExqfmbX1
M5NeyXPWwnSMtBK4V72cxfR5AfxIGolUl48xxjlRcPuNRxIBDkgIojZ/tC2CUGVh
s1m/WVxbvyrpz332pop7xeBC798OJUB9Vgvh4dcmC4xoVJ89F9EH1dBT8MnJ4Zs/
jtJ2sR9dUXUfGvv/fWgt1K1IYdSnPcLLofhU7sFsvQwtLKbTmzcAgylTyB3x8BE3
o7oSKj+vX9n/2b+7Y1rwM7c11wqtmFPDUfapQAuKoX6rInoRpzMHl4bCcti5GMze
hgXaxSXd5TIU9O+Pl2pVYWFgoMMgHT4DTFrmZ9Bz9aPYlVKHplqMmwb9IFfcDFx3
WhUPhYAuyg7ozRzFIYRbdHLrT3V2+fqmU82fhix/Cxo9sDlHVSS5L70fS5iuX9IL
mQWPUTVHn2KjhsXUXUOD0qHAqgWZamfvuvOIcV7IlOa8Ok7kth+djJT0E2p6VkXq
exDZdEl2bsu6+6q7ZmgEZfcaRDFakHP6oL63uE3WMvcEm6t2Fx69mMtodnyRuc2R
L3O4R/xi7x5VAk2Gc4znhzCIEh5RHuWzppO8aEEYN5y1WUW3og3TdAoelf4dtzOb
mr226g+7+JywFa90paui+k1ANM/J3zvb1SF4se7bS7WrdG2lv0Yg0uabqjVY0X5o
rdRrlzEEi2AdVXXUkBpAFeLE/aSp5X1GktWQAhsbv0wAuMnlCOv1f1u6YZDIUUak
baVWBwEhSIQYYthHs6cM++YWfDVazyc9PuX5rE1dln/4z+pYwdj8f7OfWC3DZA3g
yZvHl3oiaUaUYg6UG3XTyiGuljLNVwgLY9ny5E2EAr2BIySAqqwMZJHg8ab5mwuB
16OLL88s5sKR8zXWHK59NCzJiDeXJ8w9VB1GmdmAo2qFoG9SDvP3qLlslewlqeoX
8moH9u2dk3qHsbPCAdxMHG3ffuA5fKyfSsW69Oyn1kLAqX1tGy4S3/T1/2AEbtEP
kCz+KUG8DesHSgmyFiYwxyDk/bfF6/Rja8hCi3BtP9ZR7bVattPPaByNS086MWgw
baDD+Y7LS6Ow+j4sx4/CP6VwMCZiaNMfxhvEEkFsVfjFCUhKKx/lx/6DvLQhl0xm
1ub+DKAbK7aX75RzsTjgwqPAs/VXt722K5S9cv3dRyz9xJRQBWCsUL2dJyd2Y2BG
mif+F3MumyVF9+k1CwiXEiP/RK6XO4owW/MlvXW7QAzB766Thl6+M041CmAOyHrO
9ef4I5LiPrsIofm7YvhtOeQKLgbRG7P+uudgq2SkWY95VdniSl5NHXwGU5cVeTmL
KIZZyA8B6AUDjosOKWlI6D1IC0d3MDpd4KUYACZlbVcPcOYwnCGHJfva2dkCMNhf
N0DoEdNDd8wHyJTblgSToFiKw50y9F1z2hrVB2Y9/cJAFjE2cO1Qd1Vv/85JTmBZ
m7FQlhMN6HFwBq+qXShkHGGvSZKzlwbl4oS1NjKVSWs3kcK9JDzY9PrB4mRBrVsd
BnTlzsRtMk1r8UTABr6x7EcQYEgiY9aDbGLVJVF+1iFtvClaeJEC41l/VfKuYhQK
t5AIUnoH0nKmMeTzKEGCGXrBm4EL+lnNeM7LVKuj+6O4tq0bx9edFjKVG329AnhW
U8HDTglOKQmTH5vI/b0LJChT9bEk1QTCmCFYc1s2Umm2+Y4OHTB+Oxdech78Pbpv
a8UDesskB+alqYJ4rShLdxsROnweOeZjiWYuTuj3ziXhE34iHo4wcAL1zTcvJw4E
WSNvSlA5sWWlRPjjDwci28K0yJD6XXTbN8rAEoHEWDcVwvtYNAyE8z9PPbrJII/Y
XNUi3zW97chxdQfMSGLfRopVQ/54HiLviBuGo9UQ4OGO5DUboqfeg8SnXDgSamaO
dOSdv8sfP+SRoK5eWr7/z9npeJCB+0pttR0uK+ErofWeyz6rRsLSDgNV+aFi/P8g
Gu4UldmzyHFFJBOuUc5BrzpMxD75YO/ZcioImy9fGyZ74vFPe9ljb7IgOIrc8pq+
Kyka7HHqetXd2s1Crt2eQ5wDmmfCbVrTD+tv0O5Qd/5dY3+hF7CXP3IDIn1p/vJW
uMDx7eqTzY3s3bKRByC76zcScmdlOV0C8GhKAFTuk7+0o29nrMncpVyvNJ504c/5
3cItuFzt+CryTW2qcpmht9ipskW/rPsezadTvrk3UDVNN4nrrjb6pcM6mMhfBfSL
BcFL2j4c8rkOo5AT4gauPNC/BZkY5WgrgCy2fTqy0B+s9CeGVYp5tt6ex1M4udL9
h2nnvPjucbK0yKnr6plDFsQ1M4b4nzaxcQbU98Tu14RweRmmLXbhFmfQl7E+tSN8
9IYbBtkyJM7aRhOXongZef/Aq8rxcwc+kKno1+zpAJWPdOuu+/4dBRQJdhDr3SUx
F0DNSldFma5Liocoz1aRZoA0q4H4e49da4mItwocF0lE6dcnxvuejzz8cUbQI415
m8hqvLyi8F9sKiIF58lBjY8UMJ5y1tR5lqwtKVTJugncWEeN6Gxobw0h13jMHJhK
1c3OZ4vEmc3mqTpdJo5gcxVoQB48ESWCl9f6QGb/9Rg6wiaG1MCks57FJrS7QXo1
eDZ7fUio+cJFNNO3FTuT9SPhXIYcJcl/oIaPhwu/EuheoNiBddu5bbCRIvaIxG+e
dEyUw9cCXGGmdUTAy319Q0LziA0BJXoVlM3WlnoJ8QaC8VHGKCCZxRw7D29s3Mqe
74HRPd3OHhkDbvQk+C4eIFOdPKfvqUgYSql4U679R98TwyQ/1dYS2FOeCn27Yq25
5Hb8JUJOPQi+x30jqh7WWmJCqzGxlWqqi4eQJWY5ZvCCFD9aka8lybysOL4Fw5SS
DLJQa8sQI0JXZEciGx9NYnKQVBeOvY3y3uwgBPJl1dV5wmqWEheS5+dZ6lJvXNYV
9rmKx+EuN/1NjnDkntu/cxiH5eFSPVmCx3ijYPaCvKecWq17l1bqrOZ+/AKsbXT2
rA+38STRfj5TVLU8BzXAPkBjQrPrNBRgoB0YNQuJpkqP3sogHP2ClPFkDSLekT3C
SENEOTQ6N1qd3YfRXgUmGgHWR1DFLZuHHMhoKbGjzKt6kuFs/yAFmdo5PiZZTpjI
Il7EJT/7raZ4j579IW6tHOYB+zeH3dztBXtjTTgsJgate5ihg9IJLGcRFJqESO47
WZn6YxYSTTJSSk3rsn50lDRThizMLLNFoJGHzFXjrPi8nqjGXsqaPKkwahZieqwv
vOueL+Yn6jWLwNKXdZbiclxX8w4Oja5WZbSxoM2m5NcAIja9LJMd76XJpIgIgb/S
l77CaXy0762T9I86x0iaVl0fdyJWRvqIVPWl5KihlUYggEfzUbbrcVAbb4OSupYv
MZa9ms2JP+3vxewISflkAsVv7fExzhJ148dBQygtEbZkz5vjktxZa13s4wFS+C8o
WOY8jPeUBt1YIk7Pnq2jK0ZTBDYls7bNjceUfhWg5Rs9S0EbMMU7BDoV19QH5JA/
qoKkxSi6F/iVNMmnvjgwccCkXbdyuzDknSP976a//RxQeTl/DE8tuPtNpXN5NYf0
L+xPuLxtpx33DmY+OFHZULnSGaLlDaS3YeNJqV6aiKAkbsd2xgUKhSHa3CeNbsQh
uzPKshDYQyjbD+o5SI+Z8z7gqGKTsNGhov7LrQ7YbxQeRX8Cl1cOZVrkrF2PBDzT
UeOkEu6VltKOt79GfVfUWv32zbqLmj5gmJCGP2RMFYODopgzXjLqfiByRcWBqSQJ
X3IN6rPRtqYXPLWU1+xD0vrNJ4mWcJN5UAv3C9qH6/VSvTAOsU2Sw9FLvvC34veE
xRTnnGtnGCNyQ+q7NNq3xgsZUWSWB9h+6WYq65sISUeovHPo32yA+1t1p3EJRt0K
a/G4CcXCZNfK/B9LMgwJG+yjdWG/FtMJAoRFHMQshSSfl5RVCobRYks7XvPcWBGs
QgQbN+gGGLui2CBjgzYfdGZGIUBa0wVrbQ90gqtMjZp2OZShOdlrpGi10deryBQ8
BSO/JgTl2RmQ81MkYiySXeIFz8mUqAAMHx5QFmI/20lv7UG7EBW/ZOGQSCSYqmwu
EVIqNOP5fYx/N0y1WigoxhiPrwFpJGUyVobvtXG7UwmrFesnh+k3uyySseZwSXni
mEdFTAPazhUJ9knMv2FY86tHDJKV9pipyUk4uFUHn4u/qbGzl7+4MJTQBsZXLpMD
7TTUXXrvXjrVExoIOjahQF9PB8L3SX9DQZsSzFmt2hmfi20tXNukfEW9IzieFl0r
G8fNoErTpmOwEmdXgb4BJn7ICLh6/PJOOsgHuj0v7dQeaXBXH20Hb+t8R2j5YMwI
H8wL3vjO/UyDpypmF6d9sW7X7yTYnOJR4F8bhlZCfUD/yZltPqxyB8XbvTrEHTeI
3I5wwBgOq6J6MhjADM58ii8RteWY9kmmsNvbfuwgf9rYUh4dIZATrd3lqf1tzoDY
kYDv/oWPQfbUEaBKlWQ/nOOJvrO/kDRv0CkZqaz8QAVcc3xxgv6+P/+L/uxIYoZp
90RT8sTm1B9HQ4apMd2+86bMG3DmAu91DVskXY7IDmOZBbqEL+E97sx9Wu+SXS5U
WjqSk+AL700rAunCXnQiKy8FcDdL++KodhFGyIsLhyuGAZA/5Ww8uqBOIY9Pq0Oi
MAVzBHhTndN/yEmpFadArUY6e3av1H3xKtMZj+uDdezVCPMYsf88KlhbnpvQ5DDf
7fu4hliVPG+TrMYyZwjIyrIDvIZvvIN4tJknNVV8g7OJPJR+2bAsPrllGEResUhA
iyIEo1pSQwGur5l31aGDL+wX/vyHb0RN0lulvRccojpI9mo/sPwNztuh1kHGDhUp
a06Yr3WnWUM1/svMbrwkzbQzYNBGpppDxtxiPPa0iRTol+M8uM7S0sYXGcQnMUZe
zCrLxmbdvthK7ve0KIUMRPt0nXUkwPptg6/ENSUXKQ3r7WxIVAtWHzCwHfgA0+r+
pBPB4iq5PsCO2BZl7CAOf4ngaOigBNUC4ywnlNThbGX3zLLhuqN8L7nuVGjnf0j9
4BioQV/gifep6GxwriACH10na+EHSo3CF5gQkzRmF3L8qaGl4rzBzDsXGKJ+4Bo5
KlTc9BXAJA1eVPA13vyQfOCRRENwTbw4p9l7Kqie+23WDoupc3FIjOqkUNpirtXU
6jVpN9a6goiAYwKHSkQXmP7uuGI/eQKqdsOyGG2btgeZVxAIWQKdc0/5gWqT0L+v
+e5xRCYswaCctwEUlXSEPATWnJhXnL4nIlNeSmKiN9zLZpwCKYfGT4JhgZp2wTh9
wiQRQofPawUxaNnPSuuDKyTqKZtRhBtuDbmqIVM/9FZ4jYMKjr2zMPrA+ACChBqa
7N23ZoGce4UloJAIWOzbG+JBoKRkhRM13etrhfzBrmoYDv6tDm9Q7Z1foUfVIE64
q4BLdtDOAQlkbZ+58YwvF7UsKd2c6LBOjoHCj091QAXemCVnZUDeIO/BruR3aEU8
L5SB+mzkT2OIH2VQR3v2A/03n/m1j9CttWTihYMywUgP4NvUyLAV092UeOt9I1DQ
xmUCVu+5NDOqc6uTFtR/IAcYIDHaPv67ben4EirdZSDOWfbOfJQNdM1IEJTSJ3ru
qU4DKxUX5o/ksnNgZdtvjSYGg0l4KIwCg55k928JOHYLWw5FC21TPcr6TR6WLBh2
oIJTyUfyLbFZbbkRqHb6fNNDpcl81VY7dhmfhtiAi8b6PMLGHKyN2nNueTVbBFje
NIQFw+hP3ZxNvFdtwrgd07YFytdrTy+SgyErjarnKDhkYYshmdPNV14+7mKVr6wJ
Y9a9mbNsYkYLZYL9tufXI3UTLA++d0RfMUcknLQbSewsgZaGXyLf/DmXWP4JzQVy
MRVvYt7IphuqyhkHbLPTFN1j/1YsH4yjC8ABQcb0YJYQTJqLHguTt+29+lqit9sh
6fTBg161fWYuwW33dwNu+X4Zn/rtrKQEHvQJ5snwTviB3hqYLd4aJOzxGc20VsLs
DvFnHXnAdtmbJ4L3VQ1v+3LR85ZlNGXrPLRwSrlm8knEplB3u+1l8LgBnQNk7mBt
DsRR+ESHaHgvpyiBqHJgM5YL8L+r40JUJyx11QflWV6kxFq5a0Px/YHTySldvVkt
t15QVc+Ab5WFohkuLqUHfZLLLJSID/Q2FDDLzml+dw0aR44vSyyhtWgdgY7wpzNF
GyFJNjyQRJ3yFzlYraZU6mCZTRZ8tv1DHMUSqvQCb0KavLs2XLk3kQPbumKCSVB4
3i32G36ac/Uq17OU695cu96hCRglgjaCW3Ev4wIknGT0u3k+heOOEOg1LvFCbwsg
L3amu6zAdmQ2o8MHoQU8XtBkN56d5LAjRn3F31dKH785xkpq4FDRXwh4y7zGVdlI
9Np70L37OU9bul+/pcEotKf4XLSY4BCjxEhIVtag6gKBmYlhQbukjn8YthPAelyx
q06zJjjtqhfN3CkZ/OLEyeI3LSSKjyM2T7LNDhmABm6zJPnUjIb9m8dzSUin8EN+
h+REu9gZ0hKZT01ZyLxqcOdJcdLmToSgzN+fJ92azqY4eP+CykiSPuFbC2E0BlaS
B2JfQ3yFXCntZppBlgnecWg5+HqeFwW6dQz7hC+KFrUPxByVDYyN9WvsUvaP1E5G
NmUp/jNzj4bmQ/DqxhioEoBoU/7X6r7pq/kmmSqoAbe7fencF05OIN5sRq6zOl/6
G2ntsVBeGC6SIpWxrK4HfY3LiI83gKeD+uH9K/g5Yay6fgEINnPqF9jScBrVepPt
bNdGex9xyfpyzWQ2J27WQ5o0fUoHvHk0UqhJOeI3KFJgt8K7kgvtXaGyeqKh/gNw
YuDnCiqw3jNdq2XT8uhiyflv8/keTSWCYWSgLONgm8slEUfwm1SLjF3/IAi6A9RG
e4qLUXFfEJDM+2LCMESgN6uvSNRUKHQoRes4N+WjmwsVzI799/Q+OXYb7EMcUaNx
Q0dba/9vXR227tMts2+zGVREGWdZTi/ZUSEYHe/lNbv2BykrJzrbGgZZKCqV2RHN
B4OhUHlB+Jg4yGdCPk0y7QztcU3b70/InZik74n6wyhdVbbSkpfvnPtHPHEZhyup
Teay36NNVchYQHbKpe+ToSV1xYCO9yeBnBIcRPk1N/+qJlsI5wakwH7Od2USlj1S
NyiuCKGC3rXkl04tIx4tm5QuTihsZqkdNSbGHjLD6YiVhZj6Fsa5TrUNYJ9teF0S
V9G8YVLo+z4QFhyMwin/d1HR0DhdirLwIO0xEfVINlqJjVIMEY3XkqsWAF683exF
vkEHcQRrmgAAHxqcQ6okCasXIEP4SzDxJI/Co1/K2Mxyc7qEI1zvzT2IarQcAxQ1
gnsnO7V6i5EQc2oyQLz0eA569UlygrKf77ObpEjfhz0K0MEYi2gNmsAiy+rMJayH
fwvYkMgYrbNjUQQiXYyW44NvotlZP3RrBSzUaOekj1lO3CgYHk6N6acu/s1ghxFx
oTpss4jGKbysfahc3AtbUhckv0n/ZjIV9o1wxBzWdecfkv4Yz5ga/MxXR6yj3sbK
oeLgY+hlFSqigDwLC9i5FvLYQLY0gAYeuoB3twTYneRLE0g00bcorzCrCxVtSzgA
7o2NCEMD7xcEtjEVeDgjicXBAxC0EKJ6YKLHMaTz1LDE+OMG7yS6XC95LPrW8uje
fprfEKLs1NSspvBNksXCAXuZUZfZLJBCDCpGxwwSkNdI1Edv/78Im3IiFNHD4oiA
HwqYXcxzBVw3/YD8GW6bmKHSv7osEX6SiXtdxSRoyT/D9aO5o399cm1uiixmNTw/
FJxyKffNJg5VPAWAELuEY9u8h6Zw7N2A2WLv5+Px6HPYYx1EltkBtEDNhozgfVL8
3wqVPlFzdPcK7/0Hz9l+JhUtOyJRcysg9kWG641fEvEeevCluUuegvVLz2tZG9PH
RaFLY2WSSD5kXATlHYAYOfGbDyTahF3//CFco7v4tY+A0OURBGhOYu8faRU1lcgZ
R0U8TnJtAgtvR9ObJmRhht/f3Tkej8bOvQ1F7SnUHnkltYMviYQyA00KkYYZdQKu
ih8Y9ThhqAERfxpDEOGDU3tUyfZ5y2aApjY3q4o8kG7r27tM9tX1imlxDC+e+STI
MLOrLdzPK1d761Pj2WX+pT/7Ez7pZcsoIrpLq/sGREhKYSbf8qXhjFPLR66Mx+yq
DEe88Hl2/lsNjCYmOBR5ZEK6mhL/nfyRq2+Ed9gyf7cQazloecNJ6n/o4C2sLVVB
51mv4zmlYrIeCVgswRNSLsL9yTmHrmODvEXwiA35s6rMG+OkSACk7nZWf0mQS/Rv
DKjOvl4EQuUY+nlY1j4mRwBP2R7F7zzK3dAhiFRdd27bXFEUzyF2KlCUjhuCepDJ
VS0kwQswuuF2YZyd8SROHLyXxty+sj1XfpBDhVsfMsTHzHGTqbt1jlRf2NxcAnhF
pI+TwBQ420javkMtswz1p7rs6RRjdjSENdoO8JptBw5ceTezGgNEAW5XrTwiiZaK
f9pBuJcBxo8ZJtc1YQmL2i7a5CbuJxLFbd7YKa9iEGkgZOsZFcMj8XLg0AUI7Trp
80TkqZTMZspFjdPPdMcRiDxHuJYMc7eCk280xSAY03LDwZ4oZ9jBKZXen1ZLf/yb
o7eo3PXxBRbOUUwJLlA1CMRDxnSvDvyZ8z0IlegHA3x9wTyzoq6I8i2fWAxiGLTO
wIHx8jbnrmaATcnKWQc2KaoMNOs6zVM2XtdRDQ6RAREKyTCqlOo43Jv09uxaKKLT
I8YMOIs48yu+zr8tmxc06e22tewdxArhB9U53j+SSIxkSuZRGCyqNF2IyG4HrJ2V
8jOmPWhKNg0bADZNfNbFvZqrJCF97ab6SzIevb6MnjdNLxUrLr2RYDo/cxgJKCT0
zDHPWxchloY8PeCQDGwJvy8YnMc1MfBeSv9KvVeCyFIRy5a5R5nrKMFWFienNuBP
Cy9qWPSIp1Vz8ur6UYoweNoJAFYHVcDbhAvX+Q2k+hmVg9kwg6Jh9kBTMMw+M2/V
200G/wzD5gPLhqzovjR8Fqq7wFeoPOwOARUAASK8IhaybQD29KFJF5rZ+Lyop9oy
E9MA4fLVeOpIzgFfesIBIDmM2pzEJ3LNstXDKogWoMpDUQgBAKKSlSCHParhgzN9
WZ4NKo+CYlK0Vc/f34W7BflmEuAILg6Y7Ka/IxfS5OyijNjSQdOULqGhxAaKyca2
K2oCxcsdGAS7MTw5NIzxgHUOv0da38TNfRVlfWtIY9pHTTnR/j7UPkDoQjvE6Rr4
8J/zozbrq76YcxYyR9b56Y4RAyON7R0hKw4mwlA7jf4gGc6UY9z7uNhxbs7P5TEe
RplLWmdWeMWsosrsgfvUN4YEjuQtCWGlY2gdFF0LrNH1TneD4cDZJm4Q4qqKuM/l
/7O57FlSspPsc/cMeNSmx2F4abOHWtqK9UoEnel2lENVvv4gC6dAsM7WOUcPRr9B
1+Nv0p3UJBwBIN9N9n3Xc44ZK9VUe2tusL5RDMGvayYRAp6lvspvjninRVDLzBlK
H44ltBboBKmwHtGYlOnV5Uod7PityWwkrbOBkdVBWV/vY2+1zRXWgwBQn3NhADUY
wp6XGQqyzbyhSRpU+Rx2kY+rN5RdGM450HPToIFt4D//aRBZtPllt3b5YIq11xmm
1xFsyDGb3ZKDIb8CiqMimaccwGs/Gh0kE4URqyTISt5cqyGcBjYZhW/WVIMLfPEu
uuhyure88DGljgN98VhJknZJ8j7kLyzz7fqLmkBKKWnZoAbyfaFfvlXrmWhqllWf
7MA/iS9ZhEXoVVFwSYlHfN3QRZoPlc9APV/fNdLWHo15S4gGYQpZ831WwCz70coh
MDqn7x9ccasUqleImivP8+R7msrN0eZPCgzjNstqmCUV8mPxdzGN9xDLP7T3aWye
DJ69DsPQKC27Fma28KW8Tn4uEOyaI95SEQEfJ7Z1WWeG2sqOgtvO6iqHHHAPNgL1
dbO2sUZmrZkHShGFKALGQgv7YNhy7qhwC49tvB7zrEkwW+YtS5NQfN7c72XHOO/G
IdAS2mxNBg/XG7FCq/OdQnJQ52Xw8GIZw49S1TbCSqs4XfT2eZPOuqTf0KDGnJzc
Wmt/eP4/jMF3eNLwpOPPk4eTEjIVDajnfQW1ZpgI4QePKYByk0ILIFIKcGHISelt
EOczJ1op0JcfGDDISaE8dW+qPK7uji/3XKG2fUeiDDgPHCXeRJfT+XqPpHm+4w8S
EHh2NcmjwkPGKpMceYWn9vIaB2dDeKNvfgY0A4X/D2PwzVbXSKd/dg1kW/0OI5BP
Y1L/t3MjfWCErzVOKFrQW9pHAXWyoUW/NigaJBP/cryNGqoNzKowx8nNhLoWNdWK
zIdRBpUvSU/zyuNECeIu5H15rTI5Hg6MAW/XNRA235ca6KXZ0o5zDjHhw0h/oHtq
E1NupKFavH/CX9jimwpaCAFBq3nA0wqpeTpgK+ItennfSHxGZaripjiLg/IHjeTH
4ufseGDBPbN4BtfuStM3Q9lb4gW0tDFlZ1MZjNWALiZIJgW0RiYd59Fdu9XSynw6
na4wDykZrcA7BH0mY41QOziILcBlYEDh/dCIiru3GCB3HyUVvNrp7gEuZdoKfDSm
1BjDHknXMb4x2ogG6gkHhovDdnzyTPXfmh6KmgeG7ShaGb1TYjZ4tEkG9Gil0hj1
rfv18q7vu4AFsF6QGvafNAxzFJ5T2o6RUGCH5NXn1DA+bVUJD1a81jHKKVyv92s1
7jFOExGb5thGvYmBXRYuasAxsDbd7op6v8WDp57L81n37s2JvGlxmumYSvtk9o4O
teZeKDvjOKhNAr6qm0MuwMA2C336riobeodsQmMN1JryZiwFaoAeJFbvDKtN618L
gPKXUikLcFh+g+fhPY/R1bxyf7SFhJkGYsYVXbj1y7UIQuy9DTItlfdGSz4O7R8y
LKZRHbphzX1YiUmmIrVCHlE0Wuc9bDFIcCQ1XTFETMtloLX2848u/n+IQcgmLdnj
kpThL6whEA4rDXWn8Goo1QVatpSAG18jHjcvszkbHPi3QHc7gVY/y9DWWeQ2XeZE
7o94/YL2rY8VE8/oTdJie7DsMKc+DpxLCUECbcQwrW03W/YrM8rIYXu69HN/AsB/
Q4Q0uI20Jak+W14gsY83JYFS4PMWuTKkTyD02xfglTvWSN4yOPrjX5aobEi6W1/x
g5TlAPYHH5Qq8YwL4cNyN/xs+6s4dkVgFDTrA0yOOGC2kftuBVu1fcklODmN6HbO
Yjy0K162favuMDSAB4LHePT5j9/g7BMaoLJR8OcmPkObQt4X2ORK0UePnWs49mif
ohuz2jtl2BkPFqR6Xqk0lEZT+THH8z596IpN8G9a7SKExhIRS0YCmkS9vF92h8g0
0y5sLYEahPqW2poQOQnb5n8hxLkdxaPxsr2jPVUgABsAKvHfNWic16pBKM1jmqkZ
dnDi34SGUB1Uz178kozushk5jzFKd3e6vjDyH/zgrzx1utIFCqbKFzRXkSrrjvdm
z9wV+h+DHZ3mJS3YloxhEVLg27xXQ2e94yTpOiXtFC31vS3tdBEsgmVpi/uQi8hY
PVTYDhYD0Zm9jw949pQKxIrhj6BXNmHsseMMl9/XJXkfjuVWAEz1Ehi7c/oFGEd6
t/PunXNO0bqcJvs8oHjrSLSoJEC4b6D6VTm+JJSFctOGMAScIoBHkc45kiHHOF9j
khqrjtDPRfmOEMTIRimjk1e/WfkSlmaY5kyluW6oX0oiUH47345sMPxuFqW5DVb/
rRPFRmw3zmD15HDeX8jqjzbs6cvLEh3HEjW34EvBetbNf3BJ8/ZjANxLnxtHoV0O
tcLRXTK1ryFqRmveMjX4Uoi7Iph9sxjQ0Dq02bbP86Wfo36vetrJbQS/c+dtAi/W
B8COE1XwPL8IGaRipW27KL6Vv0RsSPSQpIwWl+6FklAA017JtbkWOuInOJUxkPMc
Nfv8Q6QqXXbEluR4pVvXI/GtpWKr8WjdjPmoEFF3z79ep7wFpDQzGbSupDaLc5vO
Nhw//6hDxh9cVh8vXywEH+Ft5HGX7eQclg3XwGjreYhwmgVK+6sFi6tmBtAggK7F
Mpj8YAHs5XTLml3dNhr3EHEhmbSBE4XfffFZhMoCPv7WBZyLYirBPWsf+4DxfiJE
GgQf32/bSNdsmJzQYNEE1Uw1TD65pZTAVhgtpw+0LS7+g+ifhMAF0PWmmTrVO/cN
B1E0P7jzf2vBAqfqhpAYpyGz6Qg/5IO464qpyDN+R8IuVvVL0NDjNwiM6tRENdk/
pamlvUhXzJgyQsF+8T7wkzTn8VaEosqQsFVe9qCxOSok8A3MotdSl8Hw6kREI7s3
EJsddhBGzqEcyCVlsBckgr1fGZ4UQLxjCRLymg9ZKO/YJ5A8r+sQ69BMfxtIIylX
oj4Ev304kGLxevCR49SryjCmh1uU1Jp2Ian0MGPV4fWWji9kjLKFkj0uPl5RgwFW
OtaMq4Dci6drA0CtC9xX5FNTv74Z4zPCpwdaFEeRLvWi3QZOc/2RyXolX+MaN1j0
A5SMz2+yKHu1GJKwqnCMZyv1uH6PqdsFKVfZD9f+asTBtql/JvNrTVD27eK6vjDD
gDwnxciQqlJREfOeIukD/TOa6bBiZd00674xo3VfqnwKmiK1Z6Gk05gf5rKiE86p
/VamNzlHTFrTrISs7CQfPKsUvucgCArT/VFQCY/Oy01/DI5JwP/ra91SR+T8XgTo
dykp6wqoLqkXfyIStqPJVzFj3drSK2WlzqqeV6MmemJwvuiy7lZUEfspq4HifQJR
XHfIr7LXOOit+7I5xp7F45lxT1p7hn/lwfusScrwr8RZQeMwKPvps3+kjHOuoxpY
ANy4T9Ey7+zWvC4QeFJ+fZImLW7kEzyw6REGdhADXZfI3A/XD8AHKy6iwiY+sYFK
GaYyGJ9NF+WPw1nN8K2hgTdVZtkQ7nfnc6HO2ovPfqc7oYxtz5QOGZCm7dlEWIB7
iFArDc//PrIgEwJPaO0ZqEfrDj7xW/5cTs1dinOpXzjtmYPaV9Gr45LFQBGbGCFA
XNHYv5AS47ho6eKwId+IbrKvP7N8R9CDKw4Mi8zGiRScsdf1TiUksGVxYfGBBqUV
q6NFIgPDPry5KHku0AvFeNirwC+C6Ex/l4iO/FPlW15hN04grNKZHqZaI/GZlDkR
eGG3mRcxfQwQLONT8fLMtU187jqcD1/U4TFn//sdmCPNQ/m9LKv7lrO6sZtDtKFN
ZHvoMzo9A2pv+/6Jf2v3bh5y3v2nJy4KwVDdqJnllfLAdOtSlNiGao5NS+J1hwnY
D2kbiRbtmg1ggcwA/45rznAdhY+UesKhcXvXg05opeswM9x2Hx5vRQbKEb8SfWFz
cmPSWSzccM6qOePtsIltUU6DGDHzpgmJhjSIShV+kpsclyuyxqiK24dSTefdc/7O
BZCiqEWFqmP/NzjgiIRKKu9H84DEsaoezTg0ONcYuCLz7y4i2O2cCDGf/G4ohknF
OG62ycdzgcTQLXmzJ0O8eEXWk/2o+ORI+aSf9pGYlXMlWNVP/W4Mixz1OBNQurUH
bRDGzCfNA6VtefR4tJaAj8bfxaiV6Y1JTDo23UqrG08fLpTBZw1bLY9OK8zeRhkD
nG7t8kHjsTXD/VpCYftQeV1eS2U3PeNR0h14b2W0R9lTUQVd0/V4xLxPa5dJwhLC
ugRhAF4oTiPtwnCE8Vixk/0QtjH+tQ/guAdpNrN2B4s6x25VV/7OR1mwlxdZ/hwe
GPxtaNo15o0BFT/WTcb1cHj++9axHKJap3xQySx9Ssii3Pje9+BB1ADS6YfRplh1
BC1fCjAbWv+LEuzvL/b+CE7XvvhSHK0LzNgGWBvoucg8G/OcDniH7Fl3+HVaWaqK
bHtqXphyxFQCpac+Ko28AocBBHm0qYCAmxpTDytHoQknNsvJqgbE2dVPQKlHJiaM
Nn1xjboNpyU0FxXhAApff79LzcS0yeOmiRttf+l8OwcSL2RHxzvAC6CDAJwbz3wl
HX0/nsGs30KaRauCp/7UlZxtn2ulQkVOCV0Z2o2TkJZ6yJIwuYBJtah2cLlHJkJU
TVeutMbSjuprBjQV7BbI7osu/xVh3j0oSjbMimbiVxv/oe4QKspNX8KpoCypRgez
lh43PGn5TSR6vy+Pv26cmlO7uqtA2Dpb3HZHQogv/6rJLvcNif8yrm6kQrVb1Kbn
b0mjG5ofFSPjDzWeMT4dVKCdr1y79wUxxDMBDKVHgwp9XQ/P93B284ZrUBs6PH1h
F7eytUwYIcgInwZHG1uMhJLBh2gxaG+qM3HYu+rv+u873ZHBOO5d4bfC69CuvLKL
JCT2/5Sq0yRKCzJVbYxPFGJbgQV8zzp9rC9PQUOHWKib12j03lbfLQBw/XHk0D/R
p02ix+pu9I03/s8mcQLhg9q3UVdvdmhuZs15i1Il7V78aUHJIteIijGZ6a52sWQ1
dMMhjpsL6dRN4fVjEAAdVOyb/Hmwy1PiAbk0n7F/1clCpSXyd8GMTz63OLZRmYxN
Y41g16EQEdvlGMOJdqRMIJnjY0+C+O7Biaszncbn61WYAmwRoTff+b0+94+8m4nn
gf/8SesSW/ktaQIxg1UdmvS+poYclNjJ37j8+K1+MAtRPQWibOUi/U1r5YjBKhgx
YlrsoPdPnOauYzS9tTtpXVQCUA8JsmUKEdYfJlCn8e1nvdLkljF53BnIAHMwpj4e
zoNIL4HFZ7QH29UtUZYmHXyJleFLf++b+/5TOfppBkwL4DOfJT958mJ8hhkFRB8r
0kwOtblscaBQTXK/XONE0Ud+JVpJLWpYcx3NubBWiP0vWbweywDCH+EG9Yki/vON
/NWE+45z5PbkC7LeJQbh0+7Beq6x286hmNLwNroHzWHM2c/znR8apBQRESN3WA2W
jlAmGgmVClTovEqLJmIbtKLAtjthh4Nl3Ama1VOQ1egOc/8qUo6KB1GXlVB5+o99
uvszvXjgJo+GaGuJgNBtKgqgzcdGlyzpij2eMumjbBYg7b5gNANdVq4iKActkvU+
ucEPoL+SKY1TnAdcvkiRJFLh22Vg4iNKrusB2epQ6MG10MhEmYd8Yaxz10ohKcgE
KkJcbwn+MLJJuqVXZQAHouRgQduQwW04lx/f/5gCqyPORYgZtps4WCl1EAvNGr/X
qOUCwE482vB/y+xR1Rxc/+FZCNy2AX21O36aJX2a036WEhbzLKcA3TYmWAv3YF1R
FRzDxbEVUuEKxVvQ9Ewdn/GpjUfwLES7noVComr576YayBphKWwQURfZlXJ7g8Zl
utqiE9eMWQpHZE0I2+Asp/aG6ebT77+jwYUx4nG0mLs5ItQ7xdVoE8ZAsWdcCVTP
Mtg05LfUip7aN/ZpyoEJDyZrJ6913nmqlfvcJKU3Ujp9cvCom7JCebfzr6teR2MG
9CW0U6+EWJoDEvVpmyAeLfVIt/9ntl7NyHG9MILhyqw1/Qm2yLGIa6A6sl27mDiR
OYB9CMdgioC1Vxk10fiJEpLdtVxJ/vPCDksIlsrYH5FH0mgGls21yd7Za15VQRKM
gzrKJN6DiicBBksb7HdJPjiSLYB6RqwFojH5+ajYFpTVgXodLUB0Xqf/yQnOtsqY
kTS9Yg+lVtauLyvqFn4Z9fn9o7f9G6sOUjmnwknmj/4knYeJaQO2Ep3ZiOOrz1rY
s99Yp+9XHt1zrqtaMGjMX0e3DhYcoH1DQjHgXkLVqzKHTpAdZ3avvlaxJ5+t0jo4
j/N5bHd1pXIF4uMBmGGcRTjcSWz2reqHDZOM53gUSSBqj0lEFnIifM74NBjwsX3V
32oa0Uxm6yPCYPXzrIrfDYF3Qvc7/NCsXStSleXP9BfDm5n95Kr2gbgdfHaqwORb
fVHZvdOwTQ51rl2rBmlNfSpAvAFEKJbdfS2pyBruprhe2WJRB6xS34SfFFQoRlDL
JHa7tj0UcyH6H/048MQDyntQ8W0vsIzJGXcgSVUBy5RKJbnNTH0BcB81B/UjvS7U
/m/fYrsEJunrOT7Nmv1I5z4k626d4Q04Zf2b+oq5VWtKRvvX60aCdRsu5QThrA+0
y1UVLaQD6cLX2q7iwa4jaxQmwRMDpMjdndX9NZPOayQrmcpcyuPHVIcSRx9Mitvv
iR5zgbUfQ1cv7+4UaflUTHhWVDeC8TqYpKSP752WYU5//HBfZx+BDe1G1QeAU0Ly
E6MPRXv+KQo3D6Kr51aO2Oi2/1vx+IuBibexBDZpuuTp9Hsag6CgffzIq1gehHzM
1pyB4+eNFNA/p3Pcy6Xu9jka7qM6i7C4r56iG5lwJbVAmu3p5rMc4hzb0WkJFAD+
rC19LLNEr/UKa4JInyX4V2xeytkbcFsTf9Lt4H11n9phfb8bobtpjI1HRJGCmqnk
69NT//+wDy93EzIlF7/Mq9hfwBeQ0WlkrPDHJCvRKtge1vaKJYBlFP1ZtaslJSSG
bbtcFPsrzQ3eNikTQ9JZQakv22S2nHo5V+U5duOdfjRmKEjomfSWF3dPkRZi5Egx
Gf9LlzvXolKp9uytQYGzrPEyil0Aisc9m/59kHr5dbCrXL7D69/IThUKN3N9BbOW
12y2MdXiRGr60h1r+ER1Tx+dFcTkD83fCA7y8DdM31JmfopRYvAavcfGN8tk1r2M
CJ9ECCUxSMo2d4b7TvB0KGwZyxibzsWqkxrgImrqTFAjW/BHz/X9VCz2pSE6BgQe
WQsJOgsOiAZmjtrgFCGhTDWI7Bg6xpYa8yo/mP97cR/aLD0CgywQXhDqZTFCRGOD
s9SP7bv1QehL7oLlPHfZawr3IeEEr8qGtLgNrS+Bqcho5V9sc9SG94iWAsMiv7Fc
McePf0CQ78RRNemvXgvqHxYjEB4Xx4J81F0aV3VUm24KHAO5H4Q9op6d2/oD/VzR
C6TN7mMwSYQtti736vAfapBe5/qkjZUeidXxYpgzBNdmLbUnJvfm77Jgu+N3rHM/
mitiaAiToJUV1rwVewA4aYr/Th8qAf8jpk+4jklmQvXPayAxD71pCZiUkMl4eEDU
WH8JX1SQweDHGJ94HI8o9mpDCo+Yx2qXYYZAYGuqxGBfAKUbdtHi75RUaKKvQ71T
jeTg7CjLl1E1B6cU9bWPSsQjRqzLUFxwRtJgLLPFTgqrTCvYTDUslYOtULruDD8D
H00SayShz8V3iDuT2F7RvjX04AV+BNkrUiHMd5P1UUiYh0+dDDe5iUNN6bCUvBne
s063hbt27eoz/WKvHQSZhTcbnp24rscdAvo1PEUn+cI2q9csSlvW8fQdutDOekEE
YQdGCZQczlayYiUIAfHG9sKYnAwaTbSb8kbh6jA5SKcMtX3HEblEdof0Hzx8tP+t
Pdd8XQRxxQaWgfuyVVIUN11/OXRztGTJuC/umhuETnvNv6WFc8FLnNtsGq9nnaRX
BgYzSePfAmfZsFmZVxu9i1P/TZGUxUt6HDxRuJsm4M1m7ar9tpCv2g6yGLhPUFam
IEJ7QEj+C0McqrZvhc400UTSlwsrLoblmNHWz/ApcMik61uVMPyJSDbsIiMSYtad
ESKaBFSSmsQZ+qDNtCvPb7dKRnx2pnLweQ9gePiw02LCyOx9PCDKEtGXP0Fdt0kg
zjQ0HbKTTqyQPVZJp4SM+TIqcTU0NYPXzKHZQUD/9J0unm3baSjW7MCmPHBdxChk
ctPiMeaXUKN2PKU7/6qZtYjsWpGZmVx9z0a5MprHo3OCUld5zvUoLOPndaLs3P5U
16pdlP31yJ7x9LsDmPhT+NBCigH8g/hpWutOItnfwVNL7h4Jr1vdj3hOPDfUW609
yAv/9PIOC9mBNAuZHmio8k/EtQGhGPXPSm4z2428rHD2sUGON9gs1nIe2V+ZW6XU
cdmyxiRKdHrs+ZEirWi8lWAivTEwKluHOyA00wMh6wYRrvjd8rPDB1EiKXnPJy9I
qfPLR2aq9jYQFLrD2nLY6oEEVKR+Dw+i4fG+VbOUHsOXtp6UW0BwTQgTj7LhfBQL
sEZpmnfJPDBU+TJer6wAMVZRZ+7lK8zSLjJMT+I9z4F7n4B9hfzskswFcK7ZuO1k
cDtWQntcVA+LLLDFIoVgkrQrrp0CuhV3DUAG45VHWSDc2083/5b5oMb5waE2TqAR
Z60QiZZAoYNOmPgyi2WNTr8cTe5c+wh1YLhJiAUqHrr7NlVly0TXjaqGHwN3J6rx
2WpoigZxDLl+N8GBRnCALCu2T2rgctB0sySxaEC2uA1Xame5X/GBjFRavBqYKa30
TmNRlNnIVktxCIrEE0tDp8oiExZPCHsPA0CEZRHL/J8zkF4hRwVOjzOlcis/el7n
4HoQoCOrDQJvKFFMXjboZHQya63QEN6OJZY5uRH+1yDBQezkTmtXBtEEt2HI9Hp0
8Q6zv7Uh62NC0Zb34Yn59yWVgQ11GZZfvoXKbxSiIu/cEKjVdny2k4AihoOR+QL+
ULh914UTOUDdknco832zMRWyqe4me0Ai2dFsXI5+9NEd57Pmu8LP117Wd1MEXR1r
bBMZu4ej9a2BxfzE6D1dQtZrWcPJnyaZG1+SElYVnbx4JGbtXFu1zIaZL6VHqjcG
mQIYT9HZlS9oQ5wPR9y0vxBX7ye6ft00+3kXIthXXvGwBxT5LM9TyezNxEIWu/du
8smcyHBSUgAbgNUmlSvaEeCC9M4/RdwDq5C7jRK/mlyxw8GpP80v38M1/+6I9KEe
jM2F93KVsXv0ocLE24/TVBr8YReRm/zF+CuOjYvxVP6Xr5TfzDRXywQk5Q2ggWCn
8yg2NQpxeRjqsmAMFrlsKLHzVC2nemfr2vOuz69pC7ffesALyPFVqNTSWJlxKndV
hRD2HmoQXTOQcw+VyaKpvqSnqJ8FyIBpfXG2ot2kbOHy6lcE1uMsPebiodrdbQtp
iulp502m2POncHZH9G5G6Za9bXuqShtV4YPynX6REl//9evpJ8zYcKwJMsH8gKJm
CX++Mk6+KS/EhctyfZ60yPlr2Cv0msWVp2RtLzm/+kmbnCQdqg7bjMy8i6kKsP/U
DKZvWi8MvbgvMvSenQshDrI9OyObU4AzhxpHjZ6XCjBylj8g8Q+n85YG9n0mSstg
an/3tFXeePBQn8qeiEWqVr3NXKsDMOsbuWVuC8Mb348VV4H0wtVBj8KBvyYjmvtO
YuR+dmmv0DetE+CnWt3bztmbY6WV9k9VCMZqzPmVBcly0F89RkKHQ/wkIcgpOJWb
aleFW/I+JcFTRAyLJNU9LffuukC8gi8d48VwLbG61Mm7BLtUGw+SyQpb0cqkOs+X
fq+Tcw23SXrBcTHrG6J4tghywZzzns7dsnOjZjbJb2pts+Q7NN1asK84NVKnKAoZ
RDStojAQKgyJsWh/dYPScFcX/IXZbW0/xPGCFmQo5QrbgdjiawppKakbiuHvOqoJ
wOmkh5mR2XJIVD3L5SajOPh/ZtEx9NohxiZkyvg0iqmkWUU+cNNNy+nW3lDKZ+qa
C7gJHxEK1SYo43j+bb/REfiiht8LyGRQv5ntV0gsPIMqXtXnBQwMfGWwsYW2KVWE
acRdLs9rjIPt349027zxmhX6ETrmwraoQmnYLj3bqs717AbYEXxbsnLlaPJ4aKJY
1HN2G0xYx1X1oBXwVd7k8SqGpuSfx1s/7mo8ePtHQvXRI5qp2MEVWTS0i/BikQ6F
YqU4xT153zjVaXqD/51aBs3wjdaQad/beNQmRtD49K3MolzR8LxibehJKaE5BWkZ
wPFAYFrvHp+Jqzp1onfJl20+hplI6ZvxWBog5UIi0/iCK9DQTSn5qi8yJcHf1n+8
/743O0xD+DhePXmEcYwjLp9KX6Vn/MljTNL1SZaSVMPfmc0XMoFpCrcc2v3jOqUD
riIOFJCm6UMv6FqJdVPkAIoGUCmvcPtVuxmiBKJ1BhPMcnRKCX3boEwVvf83CiLP
Z20bVYc/pGq95zcKN45um3Dv3LCO56H/XqYX1weUBQEikah/OFVwgmsSqOO3uB05
EQ3lgZ0BOTdPmW29ArEP1g+CQFmMJFWZTKVkZLhPIEPG0p1q/5Ai0QPt0Wdg5gce
A8p75SLmaawp9N4bfpvHOB0uBgKmc/L0ApHD8ho65toFC/83QXQPhuFsPMku/ok4
OoPSgwBmnnvntGATVNdq6LBaDOz7UYeFG75uH918CuAWS1hdOymMP4InX0rpKdEK
mxvNJkzAdE1uAXZBb0OZPeMA8A+zc7vrFRTD20YejEjto8/tXKZsS82Wszl41mVc
V83L1fC2tQwXRrF7R1lora4TGk7t8IdAv9ZDeJKlHGgWIYhYIJNKne0dMOCeM8e7
0fF+PY/KrDxM2LlJbP38zmpDkQeG/nDlHeJMOcXnNP5JiOsHRWnOCokkWzNZBKRQ
Au4tj2G3eOoklfWdERQdZqGZ0Q8DxbLOXq77auXLuEPZnl5wzprvRkqv7W9rXX+0
XC+7hKnAOLkPFiJm5x/ffJjVGCM6KgpmE5cBCqhmQ37FZXdu21RTmhnWBRKG5InQ
PUZQxNW3BIkj1hP2MRSollW3JsMQ6Re9yZeOCY1NMglhSCvt0dFhW7wiGC+rDlJx
IsePVXdMTd+upmPveBV2hCWLGH6mWc432xfeMWtuinoB5LapqDiS3+OFHPLrewsv
N+zf3mxXHHy3mQdqJvs5vnwN91LJUY0HoXRT+RGphdVjG/nuKyY99SG9O/U9WlO3
yMJdH9/xOr61I0X+yjkvCEBPMg8uTiSQWFYWREFAYHJo58SDFfOUaB6HDGxGrHjM
Cx7sy7W4BPtVHqJRSQ9EHKAQiD6Ry53Jej3YPZFA4QGH6HHC07zWKcRZQt2lIyFa
KmtpG01kphhw+FzwLJ4QNtKeEZfdaxl3UUrzUF1h3BE+T9uFZ9DSMQ5U8he1m+hF
WDVTN8Zz1QtOcRZ7IxJGkzWMiTcfECM0absf/krtSg+v+CfuHbrgAyuDhI5nJlkq
gCdsquylDFu/zuNQFIDpWtjLEuJkx3rJXvdMc4EqKHYKyzp2WLfVEpof623MZx59
8bqahOJBr7smH/rifvjAitAYWxKW/Tmkj/PgF5MHerFYxizzpTAEY34tt/JFcrZ+
fP2BrLZgCV4hzzCyoic3l28ru1vpHRV8RTyXQMDdNMDY7LL9kPXOW4aFLrIY8KNd
2owt7suST+/XcxvbL4NI0p6ifzpMGHZaEs3mGFH4Q38aSuD5V0mO5XDFRrFol4/s
xnxzP7ukd9UPRaM0Xrr5cki+bc5/GeeXhzuWWMJsDeLhyHzawT1PSm3T+wjzi/Wm
iIGG2JEmqD352XsdkjCKLQ5vMrMUnJnSLdvVWoz/uNql/QwI/l/IIc/NZP3jrV9/
IkkyzsjDoW+uDhWcwfKrTqfVNRyTqsRoGSjYDxXjxy9NYc90Oc4mtXGuKa6yVQwZ
gOl42kI33YPnkRNwps2efEcUs2lWB9/bPnQXdxYOb3j0g5y9vqmHVfyVLN7MmDD3
KACuX6WTo9T1A0Ux6Qa/GLvWdrRV8+H83s2bzSV8reBhNdkgzuUQOgNA9tLmGehl
X/2i4Yg3NjD+4D71OpsDISLIqzjQF1dgoG97j2R+XQkTDllGemL1YqjfG82eWzTv
y2IPVKDON9sbKN0HoIR/NE91nrpnERi1K0Gh6xKWe5jTmIPohS16oxQJKo7zDKsg
Vhh9yCE3G4jkRfNqw2lX5oKPge1aT3FzSAkR3WE6IxTMHb5lRfIJSHAyRuUUdP+e
8TmO8gfJ/+9sJjOdPlN+6Dooq9KrbjnAoRRtja31uFMt98wI3KJXMLDwCmTIus/t
l5ABsFHKYzVy+Jyn+NUw4mk/4uVRE2evS739CNgIGoA3HsOchG0wMJvM+az8Ftkt
tiAiB5fh6/2djUPuCQ0ViKDFZAvNK0QQg0NctAOkxQcza4/K1VRPahIqukqqf2/m
FkCl9amB7wzCKflA3ghiJImseGzRhw7nMvN78C5JDT6Ir7DsHfMyvF23arAOcBHe
BZnpCNvCtswbKkx/pBzm7plpP/zBeeVxj2bv/2ayIqoLZUBcwZJp53oQVEJpfQZP
mcGV8LaV1/hbuOUtiH01qTtGvwx2sxRZn7DpwpnxCTg7jxZu6kELiYlZ5RxkFV0u
WuoLiDXZgp2S3WxA1xIrx41vXeI5oJuktY8g8eb7KfWXU/Ud3kmPgN0mifZ89vaK
4dcWlLlmD9wPPLl/BfUw5Fara/oM7+h+br31qZAub9eNVkKJxPajpHYWd/fGxe/w
2pFrgSbHaXQcNvcu3pwd54rrVtdRflYHQRhThaUKzNC0rF4FmOEz+MqHBmPR0Aku
uTTYGM3Ls9ShDE2opcc+My5czbTFQZhTwq90G/8sw6Fk/b067G0V+z1LT0eAidP6
icVkYrRUn6U2KxiE17jE13jV289hETvBa1NXM7YtFuNfLQ6FGK1HfRwtZ7AzSSTZ
QmiKbsAZDHesOOzvhzelR21JPsoj7b3zsuy5W8WVgCgCkBL0PRTSp/ylWP1O6g9S
E9y/BluJt10lxAqgpRSdndXUc2tWFr6P7aB6qFqKxvHprxOnAE+OgZBdcg/fa07R
ilOc9aJjplXA6KDv+YAcfh5ccN5aUc/uE/fs+sxT+07FqV+IsKtX0yC4Q31jfkRJ
GGgkDy+nXsEXNXWhELbUHli4Bs69C5g4yu85c2Z7wRqQPnoHSWAO7gDy/Z62bUZA
qVbXYv/jX8NTzwrvMJ4MFGxJ3Az6TaXz4jwLcnkSJH7/ZfgD0AE0ihVp3uZxqZLU
mcISOpnfb57PM6MKkiz/tvAlHwHP3uebYGR6N0PCValMqcTlcNm/y90ufof/4peu
/MLqmEY0+C9xamxBb7yEqyTWYG/AtvHYReK2K2i+/w7eLMVou2qeo5Fv+07nr9ud
gBWzuMN328TzActdnDD7O9rt9g4/Ra+MHDUceMGwC1XETizsh3U+zeNse89k6/IM
4TFqu3xIl8kWBIt75qJOQ8cK9E26WrqsFe4K8Usdmzl8TsrMa2z3Uks2SF/UGsL8
xO3k0Jn5PJeGRv0YdMBg69qHpNgzJDpsYkSoCjFxBdLrVsMfO0rpopwn2xxetdKJ
V1KdarzNtivVJZdPYRxZGfvXFM4shffhNYCMO6edHGJ/cUgtVCVjo1slUw7N9335
Ubdnu5Qp0yKCKKPoBhR42wX/GHT0Bc+yYcg7IqqMcT0AHCKDYYZxdm3yzENiwIaf
kuyVHetJDQYFp6ivhB9COJejqjbUsdkXByg0eIrz07y0wD1W5+i+fApJ9pXz98XN
MVcDTVTHg0XZ714MQ9PJClWsuxFvTWg4T4AlinIhB4iEFosF8t8SZA4UJKzTj9gI
b9qhHQSJt8vjeqd7apUxTyvqt6MpP/RjI0EWLjITNyV3yow3aK1RRUeRU8GKKceZ
MD5AxsG4J0CWgY2UlWeJ5GuTW550jJEpbol5MoTleDkIr31zpEnLOD5q/23NZoIN
+w8KI9uczslIQ6vbnCvPvHcdvjELs4yuLjIQevEjQ4fN7ZdLREBIv0DTpVWy/5jF
pbtV4Ez08uYuEMoHCA0WrtaVU8Dv9vzCcYWSJbFTIy6Ojcn8jHH6656AHTuVelS7
D7VnxsxIw5PtTksDGQKPZp6L1nvJsAsorRAp9a7UiGgQ/nF6VHgC6koz5bLsAShQ
yXWekX1w3Qw2hfaZ1nilHP22PPS3K31P56v5Xv+E0tvEBvTOiTa52X9ttAAZzFSx
uBpjr/cIz9rynlDirPXcx8OmYJNB2H7p5FtDpYbOJRgnt5VTEhwIC/HnPiIYZ5sj
AtNqRR2xoEjIFhELRNKcH3RhyCZwwZM87hEcw1lUmbqlaKHE1e2mifpPEBU68Hsy
c8AptNtCs87LRcQhpRVP1pRa6eTcibqUbaEKqqqTbcEF+INtZGbmFmBZWoKTWNtt
ozjTiHVWEAjCKWTyw6yWvNDy0Gqs8njLb4oOn4IXuOl2sJimDj9ttjb08bQhCNRI
+M5RaXYz0VJqcsymf1J1kxAOnU8gzL0Z5QN62ZoaXWLBGpuIFreXuUFCSVkQamcY
JFB6DuVfCfrrK/CD0PZjkfQ7WMlrWcXPpAhs0iABc4UcT92WF2wKak4I3D+JczFf
ojtFOZAtusB0jZBCwXvCvQlBsjrvmQK3ERA5XF337ShT+ttzXMgRlt0Kq7NtBXfl
9LiqRPw/TwRw21jhowfl2TxHLc2HL9+zO19cRkzpn86ojW2IqRcnDoHTU20pK+FJ
o+J3GqPyAn5GITd/Tw+KSsadLQ0Ij8mRAy+2ObGB97si4OJgiaVhpQCdlJuWZFfR
d3LsI5M0FTTQvtIoO9ElUylMG+n8b6MqRe0hiiLMrUre1EBN4TwcjgsZpaX7wP+k
U+rUOb+cN1QnT45x0fYNUTFT/U+wEAGz++zqrCGV8pdmfQh1ODY37+SYNNvf5KoS
MuDb1XGUPWFeV98ZKRWmOe5ugxKy+DsfJPMQcDtg9ReDEfDbNlwHMIIPD7cfe8MF
HEcgmtyBdqOe5H+nKHJ5p+hSSguA9a5+sgMhDQnAaq41PeBdZVrxjoVwt71/kWdN
M4sKpxV/qATJYZfMWtQ/cPIlkLioslWcWxiii9RZ3TxPL4qSh1BxuI39xPKceMXl
guLoNYS8hyPyv1ZM5Bas0L08kSd2LxWNfZtUbaACfMsbmYlzRZAUKgbsmaYptkLl
0JhOxLU2Nw0evMyNSU6yPe+sAZvt1vDY5l8GaIIrMOvyjbiDcHbB03AFqcYhNE1l
R5jEvZFkIZWgvCdvp1aUWZZkEFLtCj1O5Cr//+sI8KcFmCwwUu4qm//D+MA2ahCt
0h+UR7YbKVqcQLHOrQivaV9WSSssSca13wJIrWpmS43MNvaROQflFBbIVS422NvO
ucgmBp8knmNP/pb0yRPDoCMQELNGjAd77DUlePea2dWiZwSv6lhZD87EqBejBquS
64HBpdTEAPjthvc7JW0qFiSxVKD4NGNXRB9Q1My4Wt6gY8nsnitXZqk65UElfQpv
wvBJSwALySPBRi+wW+UmD8a4vzH7UAk6wdEnyIiJCdGZQcl/grfIv6UXBfb8GNnf
FxsIjEfaeNeFINHgJfK02qnywidl1TdL09GdS7l6PZLwIT0ojGKQXfjIO8Chebyo
KHiCzPIx1FDpNCuBrmdNU68+PIYbgzGecKpxgvL5y2o7YvU+d44VgIlgOd/Paoue
P8YHywvXUxMtxWWN4D61N4qGYzL51OjrzwacYfHJPoaw4lfnp/hXiiwR1E0A+gg0
blHdjNlIgn1AZB5ldDsfk9bQ99yCoTx4myJWqhTTeFVqt6+lrQJSFxrAhSYbJ+8H
YVv5Wymr45dY17O8kuCDcbiYK68X491gwODcHgvL1pYuEXlJc0303ZdnEob6oM0e
lEQMmT/1jwOd0M4NIDeE/QRmNCl0X494EngqKHjQNIRCVFRWb4MlUZU++Lb2xr6M
hBJp2ugNssDqOPfED5Eccoz24C6jqgsNpmUEeZh9E+fKsV3dVxbej3MlIKrTAakt
dR6LhoR1SiVipwJLIuIfHwSyJbE7mgq2fDecNrbOiSx3Qd71grATij0ch9iKMpCa
/wYi6KgWJBkTuYY5VN4JugHXZbkGaxdGMu6uRAVQbutMsTmuSndInQI5eBfT8cpI
jr1IBfubL0xfATmNSWNKsMP+HlHTUU1sH+uCxl/7sI0SVYin8MfDJa9k/2TgdhSE
+6SmQ6ordvkDxrRk8UFdb/CbdfmJUXioW19QGXfVDWWwvQGBYV7fHCrcVboV+D5R
IMdmhgRN67NOKff6oVALOso5e4/vcRWQzDM+V7JKFOtX1CLl1JtKjvyTePC3B7qI
v6ES/DmD/jFni5iGnKFmJVyhc6PC7Dt1k+TsMNldZVOGDAJSHQ8hPphn0wDW+4uh
RpBEo56w5B9Zv2UDWmC4FkV/mGSB2gYt4V91k4QCoV3HCKMnAkbRRoLUYUutaX22
Rg1t5Ytl9VuHeBb19FyL2d1iZ5uj2GOZaXZtvZxw68UfOhdrVo0GRvd0zbK0/RT6
8H3Cd3yHYFSYDYSbYyjKxsIIYS1Oc6Y8UhCAioBTVTjwoBWnPkLAFI0MFG2Ixo3I
QGeaou2CskCn+nB5JLEDeu2GPyIfbYzGoIHQ4NHHsOVo5KH8U9DlzjyBucW3QAEt
zeR87/VIq1ImjP1MHjzXe5U/UxfbWBx+xdTRmOJ5iiFHhhQDJE8yabWkVPspNiEF
OSBFz88Yar0r1yLpz4XmE/ksl/Up800cMWj5bVhgzfUJIVKN73ZYqkqP4mSlhXxL
51yNtB5v77TXn6TQuOJfNDyacrCwI5FTsXf+GkG0kG4AuSWD7oLWOhOTUgP/5PyP
a3KeHajoXQ2EqYYIBy7xrb5As6IO/sHxtIi6wPjiNflzm9K0Iv+u+3QLrQu/DRgc
IpaJOJRacq1+H3r3TgcXLvdD57xEgZEwMiTt9kXHlgAtnu0je6AQuMc1iBgAAyLi
rBNYQxDII/PJjY9/yIgaHIv21SmUzSKawMBLPHNiKES+y9p+2bgkkzIH60qxeVnh
I4h/8P8CyjxkcArHRAz6Ywil2lTVUDLVq49N2evov0eFxZQx8W9DHxOfWDdzWKeC
pM4jdUSmQKXkaU6T7f9A8JY/sM+mIGvjHNDgQHC1UvlQ9mBytzdrIpBg+2bcx514
o4oYadrUPck2BqjAtOW9NE7VqToticc1b0PzJnGcV7ruc8Gn2g6a/dlytN23hlGB
4BvaP7vNOt/RsfDqnlS8Anqlqz1kwj5klbgNauU0mrgLGqHTXfUG6C7NIX/X2e15
C60rSnlua5B5uSe17haapOzVNq7cIJbuIUGIwnYVnBWWbY7MKoGmCoLYsSeenf79
djv8vX/od+rEnW063dGBFoLpbhyMn6dJ77RCJXWkhSa3W+G4Ry/lo3xmVnr6CjE6
V8N/vWorTxWm+ts+INa0OB6rwSp2EJOf4mwN1KlUVXYFAXnMT6TujRI18BuUxuWG
QqSKBoIlXgwejGAtrChnuhxMZxC2u5/sw7eIKHy0yIGhkcXesyJnZfPOcmlHBPEs
TuFUEgPGM6R3GVYQSdOM6KSKBAFLOyJ13KssS2J9KRwcXp9pFzEzlTtlz1Wh9MFP
iQG4Tup9Dofz9YmxenWXexMVBxon87bEtDTO3aUSc8xRYPiLosAqQArr4KhxUfzZ
1ZJGuZGhZ8hTGpSuqPWQ4NwyfhpDmpZ2vJG2JKbBSUEzVftzSn9VkNFzEbMZHDaR
c/n/s6VwZlWMmItILrsAVOkgjV2ca9TSN+piPfAbehvLIhS30EQWA2nL5UUO+dYZ
GSzOWIf1gm72s7OvnFDkQeqLcOueUOVBZYLTNpghdSKHWkAaf8nA0NiSw5ooRSB3
F2xfdfPfhizWn30+vlpg6WZQuR+WzkULKRDyj6G5m/OwtOawObD4gHTxXkpZnxBo
bEFGAsBOzs9WnxhKmos8muvHN2ps8snA64gxm28Klbaq4aFL/kR2fbMjYcsw0uL0
sr7CF7qM6T8Av6naMiEQ2CiXmsRwZ6j2StU2k3lkX1S/Aw6qYCHm3V/EGdHVPhjG
gwKFJyAM3rB1EJXhghbTKmjFgaGaM6x611B8C+7s3AYy23NLv4RIce8X8rha2Lh1
kWb/OHG7abB36vHnxe8tgvNK9Xb9wBcIfPy2QuGNMcZ/RkkIuK3adB9T9eW4hd8j
Cbqi3DPo9m/U+8okZx4JwJh1XS1buHInH1Uikeu0xlh4+O7XwExMSWqSeQyohrHV
QLoijmp3e2U8C8GfdSzLeQWsJJdHVj2Gn3ciaDJ/5ClPRm+qricWmX8NzEB7C+T8
cV84cg9U82y3lvBe67NU17sk2LxzlnkwF8gs5whIKuqiUvYbsM4c4XXYglx8ITcj
oktnh+0aK6T5462S9tvgyMoQ0OQJZcaOJBTGIoMaplhRbdvU9JG3E44CdcIObuIK
pYbNJU+eACQMV24ezxIR4X69YuzD+/7VxFyLFWlm8Zh++zNSdu74cbDnh4BzCBUi
rnHS+RxHggaXSeMazymrpMH2XXgaw//9ybp3kaIv3F6mAyz4h8xwt0rCxQ+4Izfb
fdFoAzGWE0L4up7yM/zDJfO3TzIOoHjXk2boMhzsjPC76bm/b0YPKp/1RYKN29XY
aGbdvkT4lvD9Fl2Ba3Xm6hPzVeH1iSP9xljyc1MtE5IIqion1ZFZ7UwnVlHErFxU
53D6ABBzm14QBIQU3hjmQZ2msVPFOYbdkLgBDkQJwFLR9rKBeBjYEJ40uciF9np+
f+21AlUyyWP1NmkG62B+sDutSw8H+Qr+34aWnWIavzrOH2TY1AoefmTZ1x87DFQU
B+SBLQjPFJkPsLCx7Ul1qetIwx0XdjdQdtNV5f7q5QoixHIOUMolEXnRN0JnRe3d
03fY3fdyiBzIOWYFNwVO7Wb1nU1tZBmIytgVDYKh+gC9Xc0R/kMHX2Wkh5Z7DlGP
yO0Yal9BLiBm86C2TiYBXd230cp6U5TAIJrT4eDHlFGYhNvs3WNtC5NoaTCllY/C
Yrlgq+ChF7LFCDu0unJGTSAfQw9q2TX08brnOInMr+xobI1peDiKb2bmFvHEuM3N
1DhxBxrtf2EBlPyyJbmpKk/e3wW3dhZhGJb7J/WTjPiXGqjH9LGNLdIkoO9E6ImQ
sm5EmNKiXO8XpaaF6a3Q9zxQvc4l9DJOgvDBFU1yeXWBc22aHeWFFZ3rtyVc93Q8
UC3L9v+Ycb8k5JO5D6y/hGhY7AqKDY0esXA4D6meWCdsdmb3J4vKP4gG2PiqivUk
hGaFvEfuCvWwSLh0SaV9BGsyc+kIO9RtSETwvnScLbMsywvz3Js2hk/bARw0PtQw
fhm7k9o5wtG+a4JKhiM6U5AOF3J7LdSk/5libmxR+rOnj9H5FkImRUMShdiPj9by
sx0S6zvHbkWzWJBFr8OazJM98gzJADIEosWgh/CdYpmIOemt1FlvLv9tz3Y0DJ9/
cmx5+YfXBDJo3q/9lcOwx053xVKfQfURT7bNLE/gp5beHN8nzqv8uVEwJomnvCZR
uJ++oXs1I2+QRJCc3289/WVy7tGVPscNMVuW2tpGZVhhHKJSxEeYMHHWI6jknz0V
JN3/1GsPFLgvHn2YC5GFr5w0CjCfjtQAW+MWMeOyvIGLi4QK70OTKpkh3Wi7yU7Y
qjrEnhxHBgUoCHa9jwfQJu/o+bj9mSZEt/NLth2kCqE847Hq1BcFcE+PpaSd2XN/
3ao3zCA44ExoEUm+0YQYuAIKis/aLOqrYPsXL9/+HP3vRICgpu2WBKCelPACtNjQ
Owg/GaexULr3mAwZTxd4S5B70JqgkCq4MziEJPD3D/GhqlE5gnROXalQUj2MZhr3
erMWMU8Vm1LGv83ygNvghpN3PLEY8NDEMYj26GZpnduparZgFdRyOdsPG2yZTJxX
/bHoOALpvKvkkyUrPJgX8En8UI1eX+Tmm7fE+2m0HssDvMWUk2NisnZXe5JsG4Pa
12JB29+JV3rgLsjoehZ4hl1NI0Fq3VREyyrhPtWjS35PuPdr7LGAZHnfvMe1geoV
csDO3sWUrtElRf6/ORozssvyStVXB1kLbSemSLQlHWFqcRXPS7OZySRjivvbgCeA
dBKA+bKx5ayMgjaGlPehXaVX5+HvHtpxVyn6iLXtC9rCSaBlTm2pGA7AINgw4Awt
cZHAM7bnYX+E140DTQHqh7Hn8x8zrW/hqP1J7BTt96p/2f+OsGrWHgTPGMedUs25
rgR5kKKXQFghdY6DrSazl8IcC+gAhY6SE14quVkwJYxTkhVn3L645kKYynVI53sY
mBVOijQNJSQ68e5wqajakYiNqRF5ThejxGaTjGSjrEw2i7h6gBNxJ9bsblqK+o38
vIuJDm5jxCHjpi40NLDuo4q9DYhPVGAmtRmer9pxCElKt7yQX0QnECEnI090fjYm
3ebd1K036wmyay0pJYOd3n6i9r7Nn3ckU1rAwwwylTfsEmXGt2mLn4avT8HnAzmX
XP4ED6DXyuWBJcGgZetmyPmZgYqBZM1bm1mGoHjeYIKKcn6eM1cuL7Q9CaiL3r3Q
4lKKjyp5Gc3oR9ryAbswZCOPEM2Cy8OdBA3Y40q7iyo6+RcB6SgA0A72eX4S9KwN
/8mGWfEdKPRKOc5BisfYwG0dSaOKClvka43BoG+fwW9AltNgZsVKZ6/+xbWy1xA+
jLhRZIteX3vv5OJ+XAJpYVQ6l5XNtWn1gUSl4nwU3RWaongl2yTHi+FBB/1G9GVB
E9jYAXPEhNIA89S3HAbCaj/Iw8U9XA/bS1GVbS9QfqaF+lYVKvUv2+aoYMbXRQWl
Dt1nd/HXsIZAA7LYOJLkD+2lgFf4pSZzUCgjUSI+fkwTz9XVWx0Oysf2kf1Cc8Xl
E4rZt4PddEjy0uxQvU9L48OhC4Qm7VnZ5arVuActabSuaAKo/BEmtZFF0+ExyRHe
gZnlts0fH2wD91TFpLkpLHbFJG5C5Ggy2JagT9ha4oK2XP1YUzCBtzbIAdmiteUk
j9W5bY0RoTY6gNxWUC4cxs3UWq24r9uA3cY8TQLnuNAsCoYMj1s4cBPOU4GH7ITj
aVq4veGuBLkdT3NxSBWiA7zzMQFqg0ub/PxIpZ41Acs+6eAOYZtb8BYogjeaxjng
lUzAS3dGoi5DqU2CSVVEgNZsdHLCJafJysnuLWinhlHUJVIcGktKpaU8V0a5dTJ7
aLTna27ap7lQONyfL2d99JRHyckIdDUKUkqDrx4rhRrU0IM2TK1wq2JYcucxl2H4
ryh6c85QliDZVE/AwSli7/HtAqxebGMxVhce/84TtqTpgrxyPMjUcESM+sWlj2vN
5Apv7DEsP7dO2E5uXVKKQOi1xxOjVYWrYkDCFEfsjv/z9mgyEs6MQz7HoBlMgMmo
Vt5O1S4b3qCj0LWSJXBbhw26WEZnTNCjNbZT2nYOk2PN74KYaRPXXpQ5DaeMJglX
fTxffXSdSaANESgr4Z98ZFiert1DeT1MATnswAXsF8RKy23gqYnKMP7Z08fphj2e
RU3JIlEL4X89F9M3sbiBuFvw3Icq8AB/PrixwxyosboE7iAQHn+RXqbBSum+voA7
LMzouycsX56VpPEXydlBsTWQa4zGmqRY1z7VKZT8pihQ0ONwhNgGHSN8mFpGow3f
1ugAzNiXQxd8pxj0yZ//ETglQsRBhpQC/mca1yOa/IvJO4X4xKOAwq0OXxvlfivY
C1tYBbQT7o3+Tkunya/Hnp/vMXZm/CTVdvLYNlZrUeJeNMIJ2CrnL/bjBCBrBE2v
SUo0tjnk5sdLvO6IdEO3hOwOqvsWsLexoQfCtmm4P3jVIWqNkrTthArvsJDvT5pS
0A4viPmFXwUUDdPS+SidxtcPgFx28RkOW1i2oy3ieY3fGhjUpLBbYvsdbA73zZnK
qLU2cCj0sp4+WSuXI6WFApvLAfZ4ye+ykeMNrBVLc9TmeqnwwvDlqeK+c+SPLMt+
NuYJZ1QIPFkF+2EsnwbzLnzNVLbW0NNAKKN6euJ1VmwcBaSL3MiGAa/xMvu4MJeL
ruHKUMUZTO8j1uqwRO911NmIenl39S9I4/vlsGPaENjW5bNJVtZ9vxNf8YIbCxQf
2Wb3JVUXyyNadQidgbfER7G2gKv4vzghITWWcV576m4p9XX9tkGpI3AMBNDvAZaa
GDnR6YnrRuB0wn05K5hUUfDvmUB6ccZFvN52MG4KHmGnmJr3UWzBpCtMAwPqBAgt
suRUGaSnnyjR8+X/NYUe/J3+gYCX+uUaeew9CVq54mGb9IHWFFe93jiZGkIUK09m
bCw/5Nv9+SGugSm/vEbk6DxhpV3ojqmQjNHCxUjdXMkg3b1Y5NcGDlqCAghEu57Q
wlyLHNv/Mn21SBVZFL5gOCYSM3Wc5HOUNNN2sEyO+NzqJDA/HLBhaPz3/rMB08zJ
Y2C09pdznzGCDEHkvd3myhBhQJ6OYLtzcS8/eC2X2/jVX9zT0PhkQ8cwBJ3nOM/X
M+68cdPXTzeI9f5wJfRZ/CAsncebfKnh24Ws1k6wfe4Ffb4I4lNdRffimvDHf4tn
JpHsXd/BBgTC9sWHI+VjydB8QDEpCkkb8ISrVbng8OUfvaXOyeesXnyfgtXIaA7C
2K/uMx6nkHMVEjjiw+KB4H+ha3eutyTq6+vl/TPD346SLcmIgE2qR185zYu5329X
Wn0hYwmMofqxOzyxBUZUYFtNKyTaDgOmCyBaiF5Ys35AbjylC6soZbnRofc+jiqp
6z1xlXC8vB4NeVkCpv1iFJ4zuqcvXotrNgAjHBoHvkQ3T6LMlZRiWo0t/u4bDpZe
jL/g4Y6DuGPeZvNHy4DTqh6eBXLkiUKrSNiR8Mtjz2OkKP+wY3BeLz0+2fQnstWW
adBJvuHDwJ2X7U7hr87BbCaUjw2fqtVdzF3VxtOCb26ECET/Ae27YfbTIFHOhmVF
oxhb6bmRYuXKhgfVeWGixDGHzbLDXRC8NuS81GvK5mje9VgA5BHzGLMrx0JdjROQ
+ubGpSOvuiXKd3yQfxqe5vFP3Wmev0PQ7/Yygqu8HsEqPIpO/GfY2GqN+YXAnsZg
RiCtEXqNSIo7N+H9lrTbgaoYWjbPehwiQrn9DUMpYTSuW3sZkbqpjP4eibDyRLb/
T00ffXy8twHUXr+fQmrpVyPc8quHTvWshpooN2VcigsP1lsf2dZsRdx6ejI08iO2
OIOnJANFTVgURD0TdfhcfkWcCN16FE9/81twxMUkaz5gp135+bVurIUNf0aRVxDL
kn9yOinXY4BYfi4G24+hEmiGJoe0+dW9bGeN1YkPOHjwdCpPLYTCZNpDcxKzsLNK
vxwzgk8MDS/xkvmORDHW5iE9LT+tistO74T0Wp0R/LeR76jZ1XWNlEwDthh7iCqJ
NO8DdISaZ4gSl+gLga8sfip6ZmrTA6OCulq24HRUwIMi8nV9pZ2yQXhKxf1k3g9G
P5OsZVGC+e5zepE36SrQBMGfhLuaSBf4Qbw4qkINLI+a0yxPfFZaNsZRD0lQE/Ah
B/5OnqiaiEmeLRVwM5o9/nnTI95odUrBebxDLvP9MWPeL8qQ6KBS8/1MGlswg8Dz
frP31g9NbWEU9OmR2/fjgM7bVVoHAEEZDlfAPT/xwVRxEIQWllr2uJqzD/4PgE/y
g0n2Scmng+9qwm8o5d2PzZysGr0U+pTKkPCQ/gw2ns1jaIGF+OXD87jQW3mWlovL
oQ4YopIDqxHGgtLFizg3rlHe87FuymCDDU6UwCCAep30r1VPKFFrTDG0h1xYskJ0
mdgIoPB+yFVCaxvM4jviask0uQOUHPgOA041OvvKEOKW0UxPR0ZD4ht8mJKTNZbT
qXA3zkeWBzaxJrs1PzFX4g6y2M8mk94KpFS/0m2WZ0nDa+r9lGd6la6nTrK0nBc6
zfh69X6jKlQYiDdoCpdZZIhdN9NVhU9jHV0OZNjlcT4tVWMtRQLTfEMioMCURgTk
ugdj4AvILw3mfRTyrSWjjOE3ZrlLi6gDCBFF4fTfxTMTHQpFyNzywXq4cvRuqBu8
Zh3bCYDJYzZe2J9JT5GWc7K7noIW34/KJShSLQiJaZqFENw7T9/KjpKqKQXmpeHK
zFBEMXsBbmxkcmjc1VnyOVvGNJerndZvYmGqGfuc4OaYJc1b5qIVtPWunXG4KQtx
2B1tRwOjCkP6j29AxHIr6qOBLx6ellQgk6xe5iUwbvKHgQg/CkzAQ6Cv6KMNUsk0
Xlp35iGQFYiJ1P1X4oFpQvX8LjZhNJJX2q/KAyPHvfCtxeQWX0CgWzLNH5evYBRn
B7bpV5pbXKjBUUsl7qXkZJ3GJEY3+U63k1DUxIeti7TJiwyJHM/K6nGNxysstTSD
xCaPwGGE3W9YgvOjmA8YLJCEoq0G8CsduqJFTiejA82qu0lDfb56sLVctm9QCuTQ
9ZVlJhhGgwCCNuuILhMiL3OCKm1PUx79AavgfE3iwkGr6yj+o14kTxp9o+5buogs
WNdkNQtEyvXiM9MFEGEV3IaNYGNQgLCEO6aGgTSQ167VRG2YLoQFfngPgUPq6iLA
qkauVzGZK68Rcn7aw8SNkj3bon4qdAkoOqwWytTaqWOZmftq0KUjizmXvpV8CwcI
i388AsBpZh20UAlJKScHtuDQR7UO2QOy9bX3pc4ZUFv2X1YQWzPdENZEwP6Qnk/B
c0baqta9I2An7UXVTHXG6XcWyeJQunpsEa8RyRXtUhmG9uLdgaSmFY1o3cVWEGv+
9ivKtBK5PqIBzLocLcif6C+mDg5XahO3u++ltibiymD3vKgdENYFcHjeykxsJ1/7
0JwPyIN92tsjIdzC9bg7bBKtMByDRF54AZhfx+duDYFz7Zd7pF7RgmAvcnr4uc6E
GhR8a6oiR7ir9yUrv/9yWf6awHOkEkV6XqPy8Qqbof6khfdhoJhTPR4fzhowSxWb
PmvM/NrzWqdEMTHnK3jcUeufT0ZwCBD7KkIj5Vs1g9iUZZYD1b+juFhiQX1O1wag
IQZ3+1E9MINHpPzrPgeOOr8NOCTSHSB+qTPKxFvhSnntXe7xm3QuY5XIRclvTIGV
JysnrrgFk0v+1oNNwy87hEHgENKP3/lwrVPNq9GJ5CJICaC4h21NaTxxmKnJSxZv
JsbvAiswLWKuKPgHeoMjnV5nccl4Jd4Vay5sYDOExX4Rc2mLGyz2zvLqIfvym2jQ
8sc/4hkn/Yki+OhOaKjg9DvgoNEI0vSBCm1Agm5eNebkcB8yta9pFydzb0v0grcC
pJecXvl3MVKO1ipEWcKeYfwhhn1lfwU0j6zuVDt+hLBTkmimvdhSppp8vCe4swGc
wfze/KX9ZSpe3hxYEPEFUywMzqxOFlqm/3b1A5aVXKB9ag5kqWvLSUqmFFPkKLHX
wieIFaiUXnFcmkRt5BY6e9p3Fu/agBQELAOEhSjoAVgqbIRphFiE7OzqWig3JM7H
Nss3p/Z0hyLlpZUVP8hx03VMY5tQJOPProOZLEsEpW04ra1XhoEvZ+U1DccOKeyM
xUGqCIQwYecEyBQO1aV72uThd/bnNLfzdgsFUyjOMCa/HS+tFl4vRZ4cZbcbytYt
SVJw0AmSda+pnVv0DWLzhYM70P+yTs96vmOA+63k8exsQWQ78XEnqPKT+j8xGzr0
eCG4RDrL8Po+Zd3Jebx1OXwR1r2mdKNPZu4VFjEh38zf/qnpV5p7GgUXwFIscklG
wiAtxbeb11E9DArhNNDzFs/Vb5sAcWWiwyfc03OLceMeTuJEC662ZSUSYfY54z6b
A2YYRdPP1Ru4bTI+NUlVcIYInNFtrHWIlGheeN/Lz81N12EtpPq7KFJAT3ZjXREo
iYq8c5QerzAWXEBpcVuLjw3rsYAbXCxSmVaZHiEWzund6iTfDqajTlw3ARCNjWVV
XXf9anZN6oat0Zdd/nTdMkOw4vicRATjPnjgVvKASW7b/VGUlq42SBqTI28v1/hz
v8/mzjqEodEQOMeWxTsqr70a1goGJdOCJge+XYfAatMcZovRlfoT+hRBFfPs4xgW
Ia+EINiFQ6bd9vwLrXcX8lkaB0uFGdVWU8kTpC9s3Sn/n8xGUntETLXnhUobhgtw
BK0aQ7LO7I+RwURj8DxVECcOx2xeGgd4MvNsto4JHWCU7Zmvn6o1X4LrA1iLbRKh
ClZs2OnSN+l9YAITOtkomhG0cAJ68UfVA9ppM8Tp5gS4d56dI9wNAhlV5ml1k3aS
eBtAoClNF06/7+rAKqCQjdWO8f8qwBXu1wF7pDCpHM8GMg6jp6P2Pl5jE6ZagR0R
qCPAMWw0mwyUgzql4taw7hnz+Kb6pvqz218JEQx4Kj8XFxfRpi9k2t6UJJu0bhk9
aJKQSNDzSJ36e/dJBsrwxHnqg4X+75eyRsKNWP+6RAosgHjH2+PNjlgWFmCZdn51
hqRTG4rJ+1Z/+UfknQJH9R48tBpP+Ia3M3Cj+JPR+NYYggcJv4JWnqo7pruxzmFk
xiHK6NnlEjzInzowKuMzUsUeLXMQJWj6yhLRAEKtL75Sz23rR5GWROspHOzU2F8d
PhjTKO2DS90/1OxzBc/9I6g4AptA/gzsD5If+JtOvuAfsp6ZCSIhe3ksy0UO2OBH
TgI1IJVFjCRTAZpCw4RYf8f6hp9oJzuvzm5okzVriSJOrHAIyRNvbqxqrtxMCwGN
DJfX440KC43OV/OhrXuyWCL7ck7r+hh7mZi5K4FjBngoQ7oPPvnD1nUTcJ7GbGrU
LyhkOW90ieDg8DmEy5z+ugCNGWYpaV10+Br2M7p473aaLJsmp3L6F8bs2ttKB4Hb
3IdWiCL3rNMOJD2e5fGbc3eRVMdwDJdb3gTLF+xL53SCfPbvLkWdJl0DXTddcMOc
TRBCrdQatXCyFHERqrTyknm/KvZmKQTlTKoartxEYXx6ITR1KRONN08A3IVzWDSp
f7LX5uKqoyhPJgtKNjq+kmIHNrELehuTkyA39b47XQ9K/5h4Aw1gc3IkSjfZDJkI
E5G4xJMjX6w5YFYvk4Nk3YoKpbM35tfSqaVJp+spfmSUUdaFP4YFDo9TXcI0FjIz
WSdFmwhK6Av0Xc4VLHvG4ChNyY3IxEybTya+6fsJb2KmiX+bCbnUjff8lx1m7NzL
czTu3QQhMPUgT7vi2lUrlW/psYqB372yV61XmeH8krON65dhz8+gkyG7kKo81vJK
g/FYlXbjv7FLbDWDqZa6Z6LQLyxx7/oqVfB9NVee27q5NGUasIENJRi8iiUj87rr
g89NX3xWRljJn0PpnEfK7t9t0RWAQesTK0U1ifvtsFeBRDbg/yiHcx3YV4TbpY8E
aRbn/hG27BeJJBQUum16G0hQVV49pQSshFrH+gPzyXBaRX77wOs0te1QW3h1cu4a
ptTHhYow61p+/+dciK1F+btdV8H9S7CC+/+72Vlf36EIpKIL2xLba6X02s/j/vH9
yv4rh+2CtpUNZL/i4550n7GXpeYNhAlsLsxxHX4KBulBmgeDNWSNMp6aDuxbB6jj
+Ak6RvmeqzIJybMerAiczAdDlS71G9xKV8KoKEzGjT9WHJisBh2gBW99lwdRubPq
rgu457vvyUrtWsFdnOatxBnkUpgItuluBxvIOVj4duSwripZwZjrKzJHVjvCctOi
iIuK1huBamCRdw3PPaTdjxVaXlEeGjvXKI52QRm5zh3lZ2eK/ssoHLCrjxXFC8xy
uo4nD6ulUBRRA+Szt6za+NTzjPvZWQsrJOL3j1Kp6zRadZyvCVS7/+4cxcP0ZNfp
rSUUDqNBR4HhTgSHQxwvP0rf9bQbJjQF332MmwN0kuwEmVO5mkEYOkMJ9eLCPjde
Q0xkdk3dHtYgplPNPRklTsrc9Mu3o+/AWI+t1VHJ8ZeqSvlo4YwehlTR1yJ40qHP
MpWcRqy4rNAa2wQjpRWGegIorERbTwymq4c4bEqaVpAoWhoouTSCkaK1Zg05m6am
Pg85AMnIo2hLHP4scob9xHvj92m8aQ358XFJ2hOAr5I9SNBWkH8weRMFGgAkfeoH
2tABJ1z0cgIcxQmdvJMocP4l6G+0xFSLlZGpWBAt+klNBd4sBFlZFHiUdvUu6nU9
k0QGw4U/JmX03v3R0nAC7jrr7BZPKl+hIIPRXoiavKgY5VGv73nRQ9EUj2P166oz
xZBrQesodwKA1uPJ+THl6osH8iiGN9H5oPJjuxnzewp9mHHb1PLmlyMkGoqCJVaV
BGmRg23mmTT3xEbJn6NaVoe2xvPTKF9GzqJ/hx9WQ2DMTJ+YyHzP4FCkW8Z+26xn
sE3g/BkdwzKa71vdwvDF884fWh8s7nkP20Wy8M/8xoyPEP13MrRfEkT9f7N2xIi9
HQtVfpnasS/6fLLSspiC2Mw5inYMmOt7nh/lDsZy90cI0wIhsSY187zNuZZBv5Z7
JQX+XX+0h+W8Fr8e+SIwATMkKq9XQHdZgvrZXUMZ9tm8L4bEh/rBnKYLJEvUfpNk
TWks0zzH6OH37DXqKvCR87em7x4RGFNTvNFnzJNPkYLoOVJ9dkRq9Z2Gffug9N9T
BaSluVr7THxbWDPBWRBVhu9zD4W+eTzpgKGqVJMejzJsfiOrs57SYt431EKTsgw+
JGni1mPrrPhGH2tV7rebsq6HWHyNLdreCg6ziO40OIOfbNfLj1IRGKP1qwAO65co
hRNF50O+ssdn5fV0cnquDKhHsJW+HO79H/3gb7O7vsA9M5Ztd5wLYSM7cxVyor97
kBGq7DdzA5PKVNp5+TmGHvUnQkBx7tP1Royv0KcHhz2JY4AyY9j0Gpd4JVJ4HGqB
JTDERzADYeYqr960kZaYZLLG0vaxgXjxAa6vwGEljDJ2m7dZXD5v0kEI0SmZdlAy
j+4rpvGPSAqqK79J5P+lct0DXnNEIiEceZ0yUubs0lwXr4lE5blFkQPLSM8GrCdB
m+9+O5cfgw011ZBDiQiK4rZJTpyFg0lVF78dKBiDBLk6iCrJdBnj/73PRn/iDrgo
VMEuDs2N0j3uaHuZINkQC0lzYAQC6pxP9XrkAuVm+ibmWjpkBUPaEI9sF2GebHoB
/5j6D+Tp91lwQfWJWSYf5lv0TZdpBBCmFnkcveU4uiu+WQQCLiTKFniwZaFpmiqr
Z1A2WesMcB7dIzRpcwbjdgryF6jDS79UdqqYq+QnJv5QhEu4m17sq2RxGm5NOOBf
NQxgdqIbhI58iMvSJlBK1cMSzMkoOGMiLbTf7YD8/lH7a7fHbA3PUmmnyrlqWWL7
L00C+jIWZZhP11f3LjcpQyV4GGniavyGvtNN+e06gMvQBs0OnlHpMTDaXsHT6tGT
ArApnkobPalfKyaKvt5chXfkU1tDdFQIg7yKMbJp6mNS5QzjYxrD0ISbnm5IwnYM
gDfGdxcUADFBxXY7/LwQAsZwODV6xq1WSCeC2VUZopvlD/ehHupwqF7mAU1NpKvX
lguMXgLUgLF7+HOo4/VGcmZRlwca2LMDOTjchbpJkXYJZKc7BU/h0lBgZ8Sal5JB
mqtitqU+EDy1Ky2pH/nbf7JhOkWdek9MeqMMAkxhipEzUDXIHUJcC3NmzHntourL
ZCSbgJt5AYkBZoKNloP5k4LzJR0Wn9wXGnsGktzYYKaGoxDOxIvgiOwO8nC0R8Dp
JeI4OP47+mOrtTMswNtYVw/jMDNl5b2MBQ50CZ86qdQtvp4rVQeXJqF5cMuraIge
lv0vFzl+lzd+EovsW3L7rxEEe7oHI1bfA6GVRsTIlsENSTS2Dlk74ZYNxYgzntqt
+JeGe2FSmMO4fvXApqOnc+d8Or0zplnd1J8SiZtgNYIcJDbbVgWNrVqn8zZfa1Rs
IXKXHYpEDp5K0vLyls4VggsqbHzuzD9AXVKPAiEUyWq1WqwSNt3Iro7axBWOg6p+
gWTYP0JFawPJtaZ3jY0A4rktufIRZvhcgIpW1bSV+9gank0b3rCTB/fzjH/wTbv9
4PJcIR5TVC8nVb7Wf4z/5txLheXOMT2vpQzmMqbn4LDk8qaChSN7dzAN7Pr6Vnoz
+snvMlPR6pQGkVPTClFsBi/a58+UnA5TIiUemxiQndOpwE7GFC7HaRSs/adldnpB
A2omtva/T7uCLrcXb2ZNkTunTJaXSiFlqQT2yTMoNb7ag6LzdZPO1pMm4BWi49le
kFr8ACCVB0KMKrfy9bprOCSpeNWd+crHVSN6X49+YOjkhLKi3hfXUvWGYQuvlxej
JyvRtZb7jTQOE0mPkKYYd4CHm1h1W67c0x2eIAKFVePqJIuxYFx7oqC0ONGgfSlV
BjsjwowBj8ysTTsE3Akxm/Fx3yyD6Y0V55uS/9MCW1Ueih6GpPVPrJhbcprdPX+v
+oMnDPTayxg3guO3utNSeMv/PMbJLdSQf6p8Rlj2VmeJ6QRZqjpdEZG4Ok3Qto8J
0U0flJEVM2wzidoOFRG/wL5fXUHYaE6DVeqfU7EYjQGcE6nLfBaB7pjYwLLiGK98
rQwt8TbviOZ87aV3+Nfu7RkRQf6E5BVKsgLTImcC0l4DvERfa56y2/rWLL1de4rM
q8hv8ZlEn0nX/rCkzWtwTol/RCuNUiXV0G/IyrW/LV80DCnEgUN34qAhQ0ba+n4B
tlw5nvWOWYhd5ReCr1SQSPIeIHCp8JOYD/IoZ1UAZu9GK0Drhwbf/mfK204cw8uo
o5w4+WlDYWtnLeZ7ibU9N115hv5XHI8iRhIOvzLWD8d2SoinLL5RO2G0shIuBshZ
8dabNfmNiRsThN55jl6VM5p0uLn4IbhDwMKyqUQL1n/HnAs8VkEJKaX5WVpvDkNR
FBAP+A6ovvEcY6z4eG18ZlgKb0vlUq9xJqfCVREzbVZL71iaGrXCHBgHiVYgRwQu
/4YY8q5lO1xu+G3TZ2wLcQ9Y+VQOuAtYYF/eJxFekd77Rw/se59bbfrk4pvbgNGH
IXNtounQOfZm9OvIgqVVfT+UW4W1rPF3ZDAfPenZc63I7RRjz30MbU9YfkOko4LP
r1ChARPQzLkZvbvzIqbhXIqlVtVtFKds+IJQY8OJuauePVLwAbHEZAAA1TPEpVaZ
Hpw3eEvgKMQ2uhInaFmwGZabW2mbC9lO5AH3n2OeManihNLCnmmQnZyOzD0AvYL6
0SmENkNuvFGKXMFnJ89BQSearoaiLtALvK5DAibX65jdNfORU7qXIIddZLwWFSWB
s+xk2p5RSY0I5B3EWpw6z+3DvCo4dhbTb3Fvgd+O4LnUDLus37PqHj4k4kOX60r/
7jHX46o4CUmheYXSF+86nPSDaPRj6gsL1AYsbkUaGqbqBc1fcY8sdDTdlSTLcear
VYdLJdZgySmBMXDU8tjtGn4LclCNPniuv1ffKdOIVl3y1RLx9+nfGJx6G6vSV29K
DzC3qV3WFoPzFxpTeZV87QKxHtqU22vCQGS4JeuOGdfCF2gE0kum7Ni3JzcYZjwW
90gcQXm4+hhxN2UA826zEKXnGxL5wi0Cz31UwO0d6nzrs6JSyMFtI+TR1GLjHPl0
K7gL6H4Q82E0OavNiGoD7GX9MJih9Z9rZPdIBgzaFebP8DyBW3UNc0TDw+S9EVMe
y2FggSQquaXuIx6cjEXDxwTozOsMg+rSt7p+qaYTBcvGJP0Xv4NJ1dEbpEFPjzIP
pbtlIaBDARNOVcynlwSmyihZlfcXlis5bfmc1ybUArmilX5sQHfAK5GnwJftFNzB
QAO93F1X32MujPrfyboRWEDI5ceko+cBFRccqyjlQvcX9JaQH5zGYWMwIzlf7pEJ
exQP7pzMuu/7sDK/77FTV6V6WOLVBrpyAOl5zRs9fzDqhwzv4MO6l74gBa0lpRFi
0p5sxRvhDGufde7/uscJX8LWey/99Ir5e8ItLme2f3Y30vG1rV+5LIPJqLnw/nAZ
WeUwhenVaHT18pk2XljFDBTZWJvwoE2IsBpuFNN2dCWQNu2K0B6yUhHU71DpxPvp
+QHpfWl0aOvS+4WqjG5U0owP+vrYbXk++IUD0uHj+6feMgpLLri6nuABzeSReeQy
uHzWr5rkfkOmuRjDAqkcuTLFI8LRkwq9SnMiy+R1lsys2NzJcvr+eSDhwhkSolib
ScWv4GZM6aNwmE0K4GCW3DAv+E1thQCm8UCKrPLos2Btev476sUFtJjaXCV0WuJN
1/97FSJCvgjMJPK1pj6Rnfi/TPffsNLnY8AsAejVLLc/6bZFnfMZH/F8V6U9XdEB
i+uJNV8hB1l0lCfgowgyF9bL8b0I8UaYLNS2uDWj27aEz/Q+s9fbwTlfFqFl3myK
m6f9iaRdEDbIWZpxHg/w4daJTYRBF2pe74oRdoXMdMsXJWiVK3PxO+5AsgiI2feH
dHYwPK0awfnfZm9Y3SxL7p0sd8COzlKV7LAaGHWrLtc8FCGOzt7nP9e50ucLm1tZ
7pbz/fMyOexFilNdr/65vQOsFWbtDGADCKktmEKKyXnALmE4NJpjJmcmJ8WKODOb
F4zh4hJ63k18MzIQRBFpcTA0+ZTP53R9KLjYlemnwnJTwFmb/1aBzvCJglTb2+kR
yEyvqVoB+qI7lCJTDiMPdLi9P+A9cu7631znnA1wAqFzN4sh5YXd6Mxd8yBhZSHE
lPVcflcLszuNOleKgRBmKgOZ5wh0EhSc5x6HDwIyYgc2gXhyIrd+AkuSwEeezmnr
gHuWdI2P+ZhEgRppX+8zRCZL9vx9IfqUdBc3Z/zoeJac3elD1lOHup280xQdgDvZ
DIkUsKacjMjQDCrvKmqyP/INjxpK9Y+9EcrufJ2lQsR+LVMUUo15YFMnBo6Qpok9
ZRMgqfvQVHviX8jTTg/6GeCgf4ELXab1XutSo03ES2JNSHe6DZiv3AJKfPX4RZhZ
ApwAf1jWFl96bdzFj76w8t/0en7nVHeDYZEoZs6oMNwRprLv0As/X9mbhy7JnC+k
guLFO5oIMhmPqYHWRaJYBW/K0f9Fwx6hNqwW8yV+rN1cErr9c14c7HQWnercq+iS
9Gcv9sbAoJmf5y/Uj9ZGBo3gnPtH4Ybgzd94w9Z+m86s5fOcWAWzyhg6ZurgpTE3
xHxdryeeGxmpWe8vd9IrzwH9pnRwBvC4bJDDXJzgxu4CdCLQtBjEdVaa16iK6Z9U
Moy2iveXNP2y9Z7dU3TmBGWl1RmTBi67/x72ZbS62AnEd8OW0LQa9H3+vd3P6SYU
2VCIqCZwgu24grNq6IecmiEzfVsBpxXyUYbm1vdykwIuV+7TTZj2+zqzyWX3mBpJ
9sORVv60U7wk1uQ8L532pYLeL1pGstQK7XxxHDMa3tFc/8+3wNZJjd9o7TgXp92I
cm4u/xauj1Bk2iIKu7DSxpAjRTo7RFmOA0xeuyNClL7VO5TPAZVyTlBjMs80/Sxn
U2nymJF/2VIEvVpsxfZ26xPFY18LAOZFdrDxDK/2d534HqdOhfI6ZY2o+X84WG/R
MNA4Aj/xdJx6sDFhj5mcPHI4tWD78m2hGYAQzHThmjoCgfKcl36Ap7Wp/XYO3+z6
lL2/Btag4QudkD5cPzwnMtYg/EWxWQapgnv0+BKj3529wAkFzaY12aTUsWT5hfVo
p9GqeRsX+A6sYHu1JVjp3OpD3jrlGcnSKp+hGUXhgqVqknV5FOlQAfViefufGi+l
o5J0Q3xarLvbDUL6IYAfjdmGat7XfOl9PGIhSMlQe3FDCTK0tD5iTg0mbzkSOOS3
Rw36OEAxqxIV/QiHboBdQCsJ5rLc5BiYunJ2XL+SVv7ZJ/BbAZsCqvrzrMusDFPk
oPdYoOIi6JhwlzjUE6QEblCx5ksNoxeUFcwAm5JW1bQ4RkMxmI2imQ68ApzWdUeR
x2wD6Uaww3VNKpFk4AuplwzCsfKZGXvajEaEe8fh61VL2SbtMvJ+UnF6q7b0aS9O
/vdFUehQK8QktFSRB7Qf5brlp5SnYUpl5LlVGR+bS8vb0KHhkgLMLkuMzICLm11v
XWz8aDNxiDynaTjm1IpR+jENp0kOxL6eS3rDPTBVVDbE4227SKcjF2r8Jyj4vU7a
K1XjMGL8yOrlflebVLpH/UNRzk0JyA0N6WsPegF8c4CrociPIMTdyTJjym/+RFzR
ktQot4YnwplQSy4botXV03sSqmx4ouzMtWO3w8Ade7ZM8d/iKr+17G3EpuTGmogT
FGAt0y3Iv3C5AKRN7FKONL0xlEuP6tkrek+ycDPto+rH1m+ztwIUPGeFSB9VIxTp
/Ccbr0kvUsOccq2sKcrXI+yqdxTnaPH455WQ2dTFsJaADdSuQ41trQ6TOExHXECj
Z3V6cEcKaHC1fcy4gWIQ7FKGsL9OJnr6CyzPuig5LMH7JRPQqZ5voD1lKG2PA22G
ak6YFTG59hgW5fgOcLpzOOF9HZpBGJBCSwto8jwjb+G/c8dwMXrocjL3C4ppYs+0
a4Cmt/Em2Cvz9b0QXCjo1i66Btk5V3WtaWm7+GT5Bac0K4b//Mtc5H0zT2taLdv9
D9zsibMMJQYcCqqA4dpUPzMoy8JfKcVv7AoNeg5owYdyrx0W2zHmol4Kq06mD4sQ
7joZqFVge4HEDg5iI2XfxEQZVaoccXthUEMH5MONg5suiZZCMGXrYcLD+4wLy+Jv
lP3YEyXbcJZELZs76zWHMipu4s/dhgb3krHvvm/6PwciyXOF5E6xc45LpQWpUnTN
N5340v0SGcZo0Pr27LoBulAMloR0zPqYA2dRJXAWQpM+V8zPlILKaNK47Zwmo23w
LL4pYCB/MXvXc+KPSquqjfHMlf6hTgxTjHobnBWy78N2m1q8luKlS0eZNxrgEPn6
4BuP2l4SIa4tDpm0Sc2ZwjWziEQJGMvQQDpw4CehbXzGw7fgzG12q1riUrn3Ne9f
D3cyyFA6r9jjN//cXR3vd5iep+3Deey7oQ6raL/MhVxQToQEm9icN5IZTpnxx/MJ
NHhIYUqVivg329yPZ7SVDIfIAhepxqZSRvzY4oH4lMa//rixERROlcXd9EgiOzUP
3l53Ba0j8NQOcUPB/FKfvh/6Z92RC+A4fqxJolw765CB4f05gNySB02NsSAVdwQY
9C8PDlOzcM+mkZaWozj588Udg6f0fNgkAc60qMi4Dqa9bcJsnAjZSvQt19mM46zz
yYZlZ4qB+Otd//JYb4djuSgo9CAIT7lj08kaciIKk5543tYkEU+rxEY64iJb1MQf
2lGcyhj7qmlAOwh7mCx0JzfTv0l6WTpEs9g0g+XKzaPNmkohvY5ZoYMdHLAg8U/s
JkogMuTVeqR9oAhpYt/WBo9TW8ICh4+h8f+QJmC/ZBy7yEDeVpo6BmwBNbStFpxg
zOoYWz8Ce4GLI4wh3xlOOKUo1Btwj/0uNw0nBKVPELDYRG8YOrw+R92QCfrfwJ1x
faKheiSm+C3tWZi+Nyn10BH6M/ZJPN8NAiZaxHUlU9zNCU4obuhVq89771BHRtMc
8BIvJFbFW/YT219/0M0/izEaJAs4v+lZXlblpLE/KZTs21mQC8mC5d8+TqGu9oe6
NeLPTCoVWPLozUmpDx8MsFJEKToVHoVCrUVQCbQS+jIBjJslq6nPPR0nXVwWbBqQ
O7CptRCtyvNUNxzcxPfZ0Y3DVXXb7PhR65Br9KCROOqBEQxKh3HBf7Z3iIUOPptE
GUqjvxcoGAtkFUE40R7HX0CM1SUxAPLmskyjY8CijrQO98Cx3x6pi6HZV4B/PIgQ
cwuC7LVaAOQDOWl/xa1hbOEqy+9sxsSqlqNc5Ph3lwRnzajKRGawx53v/I5flEZq
iqcle/55kL/DsjRp1yrj8nob/M8GkHTeJ77YketdFbMA3z/fnvi96cs2QUYDtHNH
j81wk6HaboxSBjXA0XXzguaLQIN6s9TVq+jmMhibUs5Yg4ZCrMuXDyyOY8VTyiUa
6gn0FBMri7wX9vIoBVcuglT5DC5yFgEB27nizTxXUyc2sUXEBKgs9Y17ThC9cJrv
a+lM4cOqUixPA0ngf5Pi9rnJp22Dhwc3ymG4Pu9Yj90jOiPz8cqNIse82Sp1G1Zb
X0nH87MlR1m8JYrWNIPw7hOIPYYLt6HhNzewwBaWc79djo3V3KclBueBoKY8LiGW
e55ZsvHH7LiB22MCjfjJTEPJLJAhj2YRyrYCrINw9JceldzBUGx3uhb8m+jewHlg
lh069CRnVlQbHTFpL65dbCA0axDtKc5hpL+EQ6FdxT4KW/JXGvW6m/slFve2J1UO
0XW3ai7XY7Ir1UJv3OHIhDI2Msx1T85zEWWRUOtqN+EOgyLNFNY0wdl1PvrOrAVz
S2m29/Itdh363dngrCloH95QpLpR7Q6koAnqEOOnNytSMjiZkN1vMPejro92xDIo
gepj41jdu1HHXbXesGCs+r8LcsHT3DqljEUQptDE8CM5+tIAf/8W13LzgC4WG98C
AQR64HLV/MsH/yronGUfelA3drqxrcw9Qiwjw6zEa/KIGwKsk1gz91jnqn0YJ+xr
V1zy4k6ev0I5qvdNDXJFy16W2gq5t7uKIiTvu20AfFu5QCEDAbk7efE+Lkvw7SbB
zvdEh2K1Xm/ddn5HZIfyEmj36EDNDKvyDTOmX71re71riEpvWqLyjQjzkEpFrMdc
+xFVr6sJiqZQKQtJ2SvqWBP0NpZ/tLu1CTIDkKafKXpvKlru+SZpS/LzU1aFl/AO
CwmrQV2USm90iyAMiUi03uPSkf3Q9e9D/gJI/a0mBrdIIOa36P+5ssUDcICDw648
gaQ+vPSZi5iDvwN8ly8bVo8q8aVPy+7AtjuyBMjcSOvgGrlCDWAQhB18Gz4bni7T
YVaUGjH3h2L3tR6QwJ5ASGWlr7hnLo5oaaCdPB3TCFl5heH7IRXbOi8eXN0u16y9
iuVD9yoc/6nYooEoQ+AvfREKPRfT8D8YbcrIi3qGrc2mKmOOKKiKpTTE00H6meHc
bWxJ7KtGhSrkr/FB70Mb9AYXXClMuWXxj9Yb0b0DUqJrPRrhQZ2MFOMSfyM7MXyP
M74fbjw8TkcDeb0VZRgMgxR/oSNYdLlteggJq8OGmNy5KeH7DbwWP08g6qiPse55
CGCMG2FtZ2df+bvfzpv5bJ1bSaEzIPaOpfO7JVU1zEx0UtMhcLkBV3tOxa7oRijK
6ZkkTakFvyJruILKso/UreltqndngSVZlCigheOeUAS84YJ5lVjmS9KIriX+OvPM
sefDP482QqbLQ5iR5dOAXiO6I8bJOKn+2vVswKoLFNQF4xQsYk0N7z8hN+UelPLV
1Wo3wSqtpW+oyrtnK3CkaUhqRiHtSnOyrwx3jo4zQey+rNzPFNgPj9QIS2PEn4b2
lpOX+VUobGqvx7NwgEvvsytzN7bZLrFGzn1Vew5v8+labJTDpMa4e//omLaY00Fk
9BGvCghQdvubz3b9gEaSHn2QoNgN20PSwtrkVk4FLZZmSxDr3ONCVdoFl+aFKPmH
D/EzAbfWTtUzcf49GcNeCka13DJkKbtujgrTRP4ng1ROwugnH1+37Oogf8DbZzEM
oN0Y3eB/x5Pxm2GslDjmILf1FsOdP6RrT2AacH8ZGoR0z8EkeCk4s1ounWIvN59D
6jiSPAPAg+zHo2rHUzGk4/SYeEdM9ntSHi3Zt/irKTD+HAvanLBCG/drtBwdOeHH
q6OSdsf8g5iFyXQX51NNnHO00F736M1gdJeb6tu/+ymzcC7aGp+ew60/zP0lKxrt
sYmqVQ5MwVDIqYOXXS/xyiPYAPJsepFSyJk0bW95btBiIRryDuoxHAnJBpzFSQGJ
X4FGWA5gDn176HXkwN3l9Et3dDvwTrb4AQ1vsUeIHPCfoi9FGwBaqrHJPs49Db9v
+0ihdDZymSclIjy4RscNpFLNKpx39oYuSLJRxA1efGpNgsUFTTB8360ucY7Gs2Yf
hg5y3YU0QxB6+V08HJEbyc4TPUxZ1i/Xx2ZATV4XlE0EgV/Biy5Vy9tNNOxtCIH6
N20N1RNZL/dxkBSH9jH6tfTSYJyQxV2I/r8FuSTdE9yQw4yIrRdZ/qI3Xwsw4gwc
VNky0lOKeJde31TeSwZWWp/AvPbwQ6kcu7BtUQFsi/pHkr6ejvxtjzbl9EwF8q46
PPycrR5NXkFTfApHfkiwYccNhkCwRbWAsXPLSg1YzkyvAfvjFhNVc01jQe/SniuE
1hpuARbgBDQrkpHE8ZB8V3ryQd/3MJBA+2ffZnnlvCSPjZpY99jh5gYvaNTadwjf
coUmrko8qJnLdXGikn2TtD5fdvFIFQ0dgCHPVv2EGkovaFaO8u6Dlf3xeeb0bbG7
x0yTWGd+IIEGZRO8Du699FQMzwQdO0O1uepn01Yl+PaoMGlo9bBl5RWiwdBpFysi
lPIqIf0tyoorf57WvghARDLDCv63qPivS3AXYSgsiWwc5+HoFelIf3+M7u11eP24
i0kdm4anqbx8ydi3j8DAm+LoMyp2da1pojA8mSl8ah7W6aFD4i30kDFVuS+XzTp0
L5Kuj/atnKFiQh8IWT/AIXX9gqrfwAMdmlirbpEUmfCB1NLt0c8OwRDEBlUV6+wX
2t7WGCaeB1WAoFY8kLAluaQ45FoEG2vyyUQpbAQwFEG3XAIYnmaUs/t+22WHQ9Wp
jNcAn6dNxgJTCTC/3j1coQu4wdxXKhZ8UG1rYN1HaNUMhwG9P5LyujUdxAxbA1eA
cEAVlSk02M8InpL/R10ok3GU+x5HSV27oR7xN8E+U7fEYexLzMilINBc7OJ1DLrE
TOg0H4ydp7SznsC2m0exlLoMqgVXv+K4CoUvL9DM7G8EW030zZ8Ia8oinBbXVCn5
bLlwyq3F+qw7naA1dkCKFlaW7NwD7F0bvAR3AewOm5mHdbBqku7bnG/V/V+cEZiN
Bg+bHCRs3IymsHLUCs+yX7bDeSUxPtk0pJsQFFi38ymlp5UuncRvNd2VaLtFdhRs
jYbRFY5NghDuK1BQACf4VieQ4qs6odI/QKfCp4loRFaRD6IdFK787sUSIiBLpC+Q
IBJ4hMb9AIF8zEa/Di77uCs/JtwzwRWdvB/Qh9bzx0/D2bfCWyz6jCKMZj1imJMo
+yZ4Yl7PQoHMLemGOu1r4SSvk7zXcn/AzHrv42MNm8ibJBrSJ7giar+RaEgxOO9/
trnvqvqi39Y1g5hQ2VbXYfkaBR9m7TWMjbzYoFGypgejP/dwKvzPSGP+1JZD0dKQ
IrXvUGDEohBYfB+GUltliPh8CEh3rxPXBeYO5QihC/ZYl+bh6ofi+eadxVSEbLpQ
+eHwMufOfa1JP4EIIcRnGoFEAWVL0+NHN0a1orcJQvgp/sut+1aX8oViGhNU5OMW
4yF9NHCQu7e/CzMMF3sq2XR7zxR/AZscKLtaU/ehSLiz2xiG9hhDP4zSTOE26QeD
LEqFSC65VLRaB+LpqqfT/mi8laqYMmSj0opYF45ILW1Qp6QAyLuyF3LNYSVN7NkS
AwOAtXrM52rD8Mc+I0t+B4HLroTMUqsY27woYfZXT6urZgYCpPlNc2bQGkZ1Jm5t
seD4WXjNOkI0hmEJE/dAzjOc4GJb7Yqqh9afghX1Aym6JGOSPLxB1RFT/6CJy8MA
E9H5l6WMfKZRH7ekSBPo8uT+x/s0zJnV8936jsnTjaQsThnIMRCLN+Zg3DjeM2xh
qeUYIeXEsTVCv7r02poAPuC78RBI6zYNYIn5e1GQAjw47t/Fz3MqKBzj/SsW3WV8
ikuodQa6vRWipCNBQ5alOiQ82vqtAdTOpai7vEUm/24c26cwerZw0UqBy/EHFcPO
lLDQVU+bx4ruMA0tWm9qz5L/4tixlSjzPBbhSM7tcKjNJfyV4flo6lJ9XI8s1TN0
G/D+N1Y+szCQsTd3WmQP8+Tq33dQqIuIY+ajJJFzl2T/3x5fFPoHNsQVMEdYY3FL
NLdoqQPcFNZEM3uWs5dOqiHL+r1fRM9MHW1xMdq5xkqRhO3iAzzgQBgCK2FcOWhP
PxTVB4fxHfX18PAxncyRkg4WFt1YWotmG+nrYIAGwLp1TQxjetShU8cs/idoDlW+
PJHbmSsSeX1xTo/iFnMHmHV9jO/HVXjNzKEvzr7F5uvUlgWbqxNbLl1YeXMg8U6c
71LPF//lG8uXalys4lU2JEMQFNxeMsLSIdeFTkFRX5iYxWcnMmXtpIYYJPcGp8Ub
PVQWTJMZIYmNE4VDq1VPmXINvQSdQr0C9tvdjFnArZgNAdH8UKM5hPdXksv1gvab
q6gpCqUxn9A4MTYEXMUvnW+r97v3VygiBhvt5VtjTIrHtyIhrGMpMzJIYbJRv9HS
SJ3FBOsagcp4tQHF7j6Xay3De6HJ73bwDPgqcxTd0R2gdtmcbLvmjb1KzuPO31O5
dLfIhPlCuRtmbR3p/qOPqUE/SvWOOqZnQ9VwZqBHcq4Cvtho+HwUu25fSWqSNuQ4
wYNTALXRZxt3LAlOLraftZb1K21dLyXacb8V1Q5350xRlnc4JzHI5gyHvZfegnHh
lumGNqemdPADCYMvP53OkoMjlOvZOHdINKKABPMgKfvyDhE97ENTQ7bVaHtl11+s
7BgRHn0r08UcE885WEjtJrTZKhcGjmcbAscfm3YhSA+O4hSVdumqWS+mmnonKqbi
Vqddywlux4x+x7R61IZMFLj2ydIq+NeiO8i+fCjazup1c8ZxdHm7MZ05ICr6SVp+
mDsxcJ2Ytl2b9u1aCsaJwx12voQIcb68EivRM9qN2ommBV0upU/2YiQcEdKxrht9
UUQX4g61HydQHKTKk3YN2kP3ahyqxjglZUWcZ3V9wYMG6Xd2DTOmbr982NJZU+rL
jkCeOEnNnI/gDYV3Qjh4YZwRUcNpGnHMi2V7DhIKUolglFZSTpdcULY8/EW6RmS3
DTlI8sYKoFkOchMRL/6lNwPL1Z5f+LxnoFEeJvMjGO9rnjgpD9bhy0I3azIoDnKU
Ohd+E1SGLVJ5k9lyjxqaEAhP5/A43p+wCyZ8eM8khMxAImFkHZn32zakl/uyKZNj
iE2JAPQ6ybbup2jxU6MnEeKrxR1YOVDTWw/yXnGfNl8Co8jfeEoVEDMHP4YZt+q0
5FWpK3bbyOIRCMgmoZmh8NTp9JLJBODXr0rhGn3+WSisYyXmivdGamqZDsCF7eED
wEyflEOxju1iOkruP1vpzWyI9yro4cDzUXAfV9PMbKbMwGbK0XcdG2lTTb12HQ8E
5hF+FzPpsVxDq4YYnDRN07WlQ7/vx+5sXWzuDxqzQjhXQfIubDCGuE5n2Vy0zGpF
L4hbtD9zbCQi02wN+6Ro7Q+8lQ6aGY9G8aCY+i7ZXmEUhClxYNI/CksjfWpOHwno
6ieZt7oQ7k+7l7e7xzJpj3zm9Vc5qClvOOkpJ35GMJduMDGw2C8xBhxejxGJTtBy
WMpGxy1CkumosMgt+r0Ab3NbT0LGKUQfP5IqdY6Q0djQ/oHBM+OAi6Kuuka3LDqj
CBPmvmKQRm/Lehwk6WzODCtEPJg+TCPK5xZToyFe1s1tKmdJGPOKlU8V98EkxA+k
gDed173M+llREoOtljcAS8hGpi05yYPHRfw4qyy+nWeqGm9UuBUdm+A74smtruhJ
lR1tkNr/xhZH6TkHMMucrRidG9B9AjkirmDqfPZ8AmYIdiG/NsC7mG/D2/BBS+3K
0Hoq6hfrl8TcduY7qyWCt2cGQDVvpjULpC1mwi2S19CKH9Y7e1i0vGeSxa+NWmca
DjsWPH3UhtfYMf91XwlEuy6sZ3Ql51+76wBoO3lFAifGcZbYguaUGkqoyQqIe0cn
6pX1sPfVfPLIFZqBT9suosWnFIQrG1HzgCRqESvTBAJatlqoHMPnvAwfNwaC/hTO
AsBI1wjRVT69nfcSvPT+fq3jWWyZ56W+ka1PqxOSGJQFzZgRyLYXQJIq96y/RKvL
Sz7nMAtmhd0EyXGU5FRevG0EUPzvP0J87DJuWtOFuyHcHMoSU/hhkZDGvUP/mwoN
wGOZAdx/3UquC0XLNsfIPt3/1YtiW2DvYsbuu7fbPabxJCWfsNV1FX7aIf/OodD0
i8MTwi+OSzXhC8qFgNjvexNXq/NLPQhOq1lZsJ2uv8DdQD1uIkO6f72KTBuuEKR8
8cSNkQkcZZ9M+sBWADT01iPAtEAi8oabNG1tMzuuH3Meeo2F/zdfROEfblF5V9hQ
gxgUcm+lvhiNe5lEMxn0jI7JhP0p+2H6ryFvrT8WllhSKKJSoyhjya6PWDT83Gth
tcugHj8nv90bx+dHkCs25pEPD9hX24Amrny6IY7wd/iI9AhO/U8jo9u0RGXnEkUl
NJZRluENwDCWLmIjj1s81b0zrlZg0ISthPUIdHx2vplpLh3cioGRlHmv3gyjOJhM
PHURkR+UvujEfVYXA875zGM/0+5sDOjAmy0E3/seAiivHUgVCwZ2FVchRFrAb8aW
Y20RfJVltwBDkvR8x2sRdjrb82OYAgqApG1N7umhL9V/gpkC+GcBVbaPP9/T6mXX
ok7BjXZvdJhUpQa+y0p7qdS4TfOYO8/3Nj86lpvKGoBsBwP/9L5BNmUkmpjrmO0y
cLDlqPzHUeJFT/cVQCIforGlS57r38Yt7gomK9JCZj8wquz+oYYiggtZlH5mYIMF
obyjdlDHHimA9L4QQh54MvnfERvchtJEBILedA9zfb3DdUQq6Cx8OAgQ2hnRQjG7
wFFEXSqin2DwUoVwD7gEXwe/8vExSF/HA63XZLt9556+TUPtbsqtS3O1b9XDrmDg
XCXubC17PjTWh1YKtS9X6ZKBAOIa0U3Z1BjQxW9xJF4az15rTpMiODj7pzJwKA7Z
7v0iDoV16lzLDlcHVAANNEEVjKeL8B2EIvoLtzObbftm0wXcubD2uI3zbJpHYLnE
Ieyci0weFQH67aJTdZHu6J95jjb8utCrL3ZCVIvnt0CvQBDYY4t/ANJzjVRWtRjq
G084B++YuTwXNMTFU6zmkuGJMIX1fID5JXJ6zyOk08EWxC/eV0jefrFx7iKkKWDw
gXQDapbsG/0nelk6pSRI6ycj9sA5v0WD2O7vLA9RdcICyKiQCiQ01jKMQfbvteTE
4TfiNsBokLPs0VQHAYboFchS3Ycmmk0CBcKlCeSnmV79oGyoLe7ftf7rp2hl1BP0
/yaiUfLHpklKFbTBw7ZYvJLuPhtmFmOMpJVF0NlYls0h4nYVEkHGNRUctOIp1HeL
yci67/0CprAkeJ5lWsekztv5PMldTwOfH0Pacyb2hJiM4e9aUEOlwOw9GtYvGUeB
3F3aIClMcQ+fArPAfm6Uzmiw7f+Z6z4DoMKbi4xX2GwO2f/XaOp6JSZXiaoHlc+R
nChf/p7dxgejcEPwoCVGZxYYOhkdYSsuSNTIEPtUNMjwHDcAqVc1/Gy5PIuqZW9W
LIYF5RbhKuIbF3VutvJQPg2K9xEGyeuXvyO/mpr7HkAuyVOIH7za8UAmrU1hH1s0
KivZ87aayjjVplz/EGPROGgzFgctTkcguG8mOoeQrF1Gyeyltep4Kj8SYoQaKV9o
HAA4yhI0b4P7xhwZYTgWVGSaTTNN/ZpJ7GvWFu4Qp9j5aPjW1GSnrj5DssTCuFDo
fFbfcMwJi1bgPXw/QYTIkT04QhqL/WX926TU+5BAZguQf7MejeWiZ5/YBFu50pRH
5KaJbKgoEfNaaftaitP0y3N4w2mkDJJw47AVRrkOoGvbO93keV+3rAG8mVpuXdDs
WXg6s+PTXQABM0ejH3Lmex79up3iSlhSgsDvhvFZOx500kluulaczG3LBWOiNnZW
xKTGzN7XVtqFPhkmkprcgquS+jnY6oxNFed/2eIxdTF3u8f9QBlopgh5K1GOEOi3
ENxPH5E/mAL6v7etq2P8vrvNIYUIuyp9suAB6fJUA6pIiaFe6NmJ9Ko6zVeNaUQ/
qKeIttVA2EkW7kzySDgRwO2U8bEysZzR+UhcjxjcNeU+ky3g6KjKmWFXkuEcWxgE
px2pDONdSUnHzJtHJDIDy/paHQGqZEDnVXXnm7+/h0PSn5qjTCs5D6fpsCl/9E0X
KAgYThFcyDnhxaJjbxWkRV1P1u7EEzYHmPzUQ04aN2yWW5bC3hyjgzrjbmp+tIAz
cLBZN3G0tITMOAQObpHYKQMzoaRv4VUAqHXekTsJHPGYN8X+SblFJskT/gKlxVV1
LND1P+8xZ8buIrRMwyX2D0MG1vx7QxLTQ5tUx+mZi2+mCNoizGGPE+LldfSIX2W1
eun3Q5asQ2QYhFuoRmw0oPP4yHbsAvLXC5HvOnFlYJNeDYTbEwdAYM3NHFw3hBt0
9dhpcJAny4uM5bB1Bw7TID9eRWNy+85URRltDEcmAXXuLE3OtxJyiySbvxV2szbg
J17yFrfAce4nv24iRsnwy5+sud2Fav5ZaVlgvqGHkkbgUzqewwcYGRe9A92EXHur
bv4d4JXUwRU6Tu5Oq2sT+w3To8CQow9vrdGclmKCTW6uswqlPfDWViO7rUb/L9nT
uhRyKorgCxQMByaL5nGJJfSj44tdJJXoVSVhqW02QxAcqZSBKnpVwfiefI9JHUOl
/GqLzNzmS+oozPzNwbJMuEqRNxW1W/Y7cC1PbmxxepwcUEkdTvtqUSsq+xHPFzgk
rgRFsfsMAjdGfqz82S/0RlgyajS43aX5N2K4eKXIl2ewNGWLGNFWiAWt7qG9VTAu
SI0y2bqqW4ynokk/RrCx2d6xbApyEpGbLm3HRXgNt7jk29oDOQdmz1q7H6JSFtfq
oE4VDN3RTHv4A5Covi1xRY1/o5Xo6Y37CdCD17Q36Srq6t587W1qrzCyVWm8upq8
PhQJ0NLQWe2I7rxoeGLdROf+WuWjYYRi+5b5bboI7RvNAO4CywzRjcHpN/dxp8iw
gZNdfrM6aca5cRhIUdBPaFrmZAZzpCNvNVy8HycbyU4aGT8KjYDCLxasz85INwXt
oae2fZ4ZQU4eaHX4rjEnNRg97yKnsGJDRA4HkdQ0MVU/IOAvj/Zu8RkQIDIOWa9h
CZ/PJceuZu7bCREjKOFpmUQK5KUQVR9MvF9z059sZ/TebIOniD8ToqJEYPXNMJdW
ZUFt0EqCAEqC4dr/vyc4zyz3gFhhn7Rl+ve4p2dYnDD6BqLc88/2mp8ZOUwWGyJa
4BzOsPPBp66841TRhIV/PsvrIATp67UL7QROcSFbg38WwN1Qp7dJVt+3nZSNPSPY
bTKCyv433W04RsIzkNVx9nSau7UgMKgmFO52ey7+9Y8BuLwSqYEglKGfB8e5vZ/G
dSMqzy4fgMJvvChBX2Wd3t44JHRJJEAlNRFKJ0LtsqrEv7lMJabj2q1JsfaAdvpc
B3j20B2mwY66O5EXS95pyTwYvgiA2WyzsAZBxSERUV3T7vhGQJI62uEunrR0Noll
cenvylbLVUEOpBL4ah6BLE2RMN5veJINSwoRBeZFxVXt+r0r8N2tW1mwGvnCu72Q
0YZrCfIYSRnyzkbn4PQst3/gvsnbfalfPfXSUZyjjucgqu3XXi1b3atPxU/f9Y+8
C7ySvutXKCxnAyqv0iV7VJoWBAYIT8V9IZBA2ONeafo379Cw5q7xi7gaE7kIOa1Q
XtUd3Yh89ieunI8ot3gkfJc3Me0M5CCAsVVZTLRq7LhgNmClv9uakyAlHV1DyG0I
PR9j2mnyhFLtPPob1UuOkHx18w5dLknWOVd70A5+uxIxEyxclWmptKXX9iTrXcmt
4jr8sv+wR8KiNa76fFBfW1mMjnGENDf2pSuSqw/BlzEkNAjXO6Yh7PcbwTCSsqcM
Lv2QqugfAellw5JcadsqGaK252eE2VIye6OK0A8W65zxl7o/LKOaUeEyIoV7b2kv
httJE6A55a0/AZqPbpwrTyxib2zRUmKjyztX3p4SoYEWjQKO+WmOd6YLnfVITu/h
Q+KD4yUAR6IbCkwTKYuPCYoEgG2mmul+EAF9X4THl9G3T3ZxcfTx5XYGPtX2acTn
x9O98fVzp/YX4enxHfPA4gXHuJES4vjV3mRf9czuALJ1xSfsHQn5rK5XG9W+5irT
95WYyT2P0pCvwsRN2Vil0YjRAc9S01bXQGNvcGpALui0YO2hiHuuQpLJvoumFMHL
ZvreGnDOUbd7HFi4LDcKfHTI/ClIW56s9joUu3E4iVfwOZE83axBpej2MYeG58KC
1u1Ki2vg4HRRjQyk2O8FikkW5Llw5LOPgWafAhnSZPPAnfOHAiqP1Tu+Mm9ZYOdZ
ux7jqqI5kQLUM08f5nzmrQGc7+WLT9C67uH4KdU5YPbhxEJMf0+5riXmZBgcDf2z
r2yqVQyd+kI9jtGfFkOr9dS8zNtzju9W/PbmXX86hXEWFGZcIHlo+SJZNrOAH0XM
WI2tFkZ3D6gf2nwYraftU+K/pKEkrtd2RMN+KZ7tq80eIgwmmBDMom9KmFxkki9X
qBdTyjzsRkiSmuKbWBKDVg+H4Em57GnmgUf882sr7RRMUq1zwOUF2m7xHnpY+wYy
h2vmYczko7mIrlJdQ4kD5AKTs/SoP1DYPXyAM33KuJ18xLCe/ZQ7CxVjr/cIMYnZ
4XLywnqz/dWAwD2MygaWLSgEC3qogX3GvvoamuUFu4+ZedhIHXiiRw3i1KrzKGuR
nrUhyzBm3cgg3tCeA1fyA6n5FB6Skd2ZcCq4gDS6qco131XvrCFArq70JXvtH2lj
5j9w3Ca9GZOv70Xh5fhVt9cN35cmi6fPdME79dmrRoJynHlPwPOt6a89avolgsr1
NisJ+K8dnR6YMjIW4x1/P1vpis6Yy42sIDm/Zd8bGStn+4AkItFqwK5OHc9vIPLa
9INUTTovmqc/my1mmXCzbVUWrDmtuZNzbNShhGChve5CHj7LFgSzqhxYya8/914R
4Cqs/GX7RBtainRSIZUBCeuLhFKte9wtXJAYszSqpYAkWvVEUBXHvVocRcHLo1q1
W7v/CbdYUmq+GRSVJ5jiQFp19bocbUyqKEqSSJOvJ2QKio83luNO5y/smR2QkBO6
Cn4kq/54gAC/LN2JJLMSloKFc+CSRfYLWuFOnCzCh8IxOW1lfjldxsxBAMrj0AZo
6NplpzVlF4AWMWhkO9wZvbSewh/Pej6qfCVCrH+Ra7bncdQLM56KVNP12T0oIWsu
vwmYkAidMXIa3CUNH755ZZxIL5bvxwPp8NArCMUrE6+jFn35zPeNqxGyT87UA3nH
42SV1Qa/HwlqQCfihAfifanx141B5vHvQ172ES86rOsmWZMm5HnF598eWuPLfyAW
anVT5VSbgguB07U8ai3Ly1PzEvl3Ynmn4fv063U2qupfkOsbMvksySW+0tORpFHf
zpasWj35FwsRCZ5ioa7CPKA8UTsxJBH5+kvh3k/rDvG4sbmMHxR0sslGYIxLGF3e
o9f8BgIhsaCHt2BS2ukgtIQ8rzYyZL6+IUx+DCVKb3ZuCIjUW3fF0sJ8Y/072PNq
daZTmj/4SpDdcM2TZCbZVdmQAAXrTtHm9xqUSloWDY1SGx48frd0hUf8NwE5ka4z
zgX8SZc918/A4+ive3HlFVgoOVpuNMQa953utStHiyJ4Let9HQscXB/JMzk7Z5/h
HPSI9Ybehya0bTqBvUzAf2x5KQoEfy4/vz2H8hbne20fpffDSCKE/PR8z+fudnaR
q6MXlu0USw2I/AycJNTV3zjxiQQHIee71ejeXV5WtU8I+vLI9ybW/6xz2j+7WSuY
a1IgWhL326HHr+X9e1wR7SMqV2391W1LALOprd3M80pbu221sd7GT8PKP8hvF1ri
v3qUiLVG/sqxV3w+w7VbLHznZT7ZpxC0HtFmwHboy2fskgllXGwNS0NtAFTp/AZV
XQWJvXp2sJmwazVZhZTDZAyyspwpOseYb5oIQegg1tLVXr08Mu/kh5E3GnOKqcm1
DqMndrEcxjbxAlmnxHE9AGP5V4pWVHyp5NeZXpcoxXGhH/7iiLoTLrbxJa8+s9HW
Zw45nS7Rcn2CeDUvi0KMZwGH8T/9tf265e0tWcJwpXGyKTFP+g/BH1IxODQFoti3
09yYgeefBzf0K5Bb0Iv+sgQvrAq9YWqEaMPNkoMUDgNhJDCr8TfiH2VQqfge1cyT
E1hdLs96TQ4AmUNtOmF72Cw9Kr5LVnnU8WGMgIskDGCyWy5xYze1i2f8d1blGUhb
2AXSINO5QMhGw/LyhNkSV3XxLhWG0zj2TgpeYBLXp/gAULbki/ER7slCvJiE1Rii
5iZa2hPqM7W30UGt++ir37YGmDoqLK4QMD27KmuaRyMVr0C5+fuRQ/3oas/v7DIa
16llqekI3E3bpeMMwCJ1NGCRRBW4okgiuuDAVrufEnlf4TEZvxiJoPJQCczvsJwb
eZe86aSOob5sOhxKBsTNP6BqQrHVOpXe+U+3nWMUxmM6xU9WsHnVQ4PRtIEQ+7KO
m/TGG6bvSorCRtxJhmcZKiePFzOcLvsUMBHJwMzCAjpFIGEeCJIVUOkpSx7LmUoB
3EwrBE8kv0WFtrODfoyHAL/HFvkrt/c2FdLf0rvsLQT5rVcttRHSDQmYEEowaq9y
qkhWMjSiiFQXrDBHe4nqwNJgQZFZougq7MXgMR05gLMjhiFX//X5kOmJxBBaJi0J
8soacTNwtCXBj1perdy69RMOabjPHH6M3c2fZr/1rdURIoEjXziOlsNuR+QYwzqc
iIBd6MdnlJxVLCtYIRKB30ZEDgdK9kJuqp2ohwsdhEoTEOgbv7xJCRr/uys1nUDq
BlCkyDQJMztjgBdLhi4ppPmqjUbGbdyh6kXDoKWtiH78RocEmLQtuTt/bTS54en7
t5xL843SJXJ38eoPcroGHeQevFQeWdDgdnwsRtT2abGjdTMDcjYkqrNwGufNaW9O
l4OL19L9YGj33AkM6QePNCModlnSRIjNmczhbzvceZBQATaL5CNAfzS3C0V0+VtY
OqaX6nakTMs/toG751UBFAYOcF89YLTnurvKVw4wx8JuF6z+Yc/OllnqHoSf5u58
60LsRbQoOoK8NLxOTYc4lUGQu3XtZvlWV5mX0/8tZmnSNsbqdyeOQTbuG90ghwT8
6pEmkZLUIOZM1pJBZzjdjo2W10FM9m+r+r4uXBxo39GyS96AtrAniRd54EYdiCDW
rKg8cyBfCLP+YUwv/9mk5+LjCgDfChEAbuEBO0QRhvBqplYD52wm2SxJvbYz0D6z
f9AE/fxArPnChUFWoF3ykvUDU3lbDlJOOdeM4cJ7sHCnkaSnp+4BTOuMhTOewKdH
2BJG8IB2g09bw8Oth7RSRb0KWY/J6SgGyzb056Opw+hJD9RECPwFMLM1qyOS0/al
/wlt74edl4E0aWEUujaL29/2+fS2xIDHWSI5JTR/hn1Bc7jf/G4yX2VS8FJrz7GC
ZuFqydz0n2CtI+W+AG4VQ4jQeBNCN9hxWCv0sA/VDk8RUMg2/LYmlEWX2V9rXFTG
JO4wO/a5BdTpAGDN3Jav3ggKHAc3ROpgYHXvMhrRXnJ1/JLPj3MzB+ovzQ30kFa2
lShPMzxesKHf8fscMv/ZyS/g16zuy7MoWmvcwM2MerFXT8vKporTyP+b8K+8OgQd
hXkZ4H6IlK5AY/T4ZiEwT0oi4u9r5S9dMCeyiD46C20Fu2OYOWaKec+uwgyorlnl
Hr8JfNBNMCV/A5II6BXXgHiI6xNd56cf+EJ4QHfyTH4cyKxxVkeBF0VKBMsHaZEk
s31VLK6LBWBizExENHGrpbY1KmcmBTFSSJhDx901xV3f9zaDJ+4B73NAk0cAAhmd
cTXQ2/HxdvLLRb5QbtSQplusxyAqBu8WReQ579pT/HMRa5mHhGsV9Q48KWxZ2gDm
fQeNsDZoZXkgDfu3RiMA8ffv2Gk2CklWFYnNAY9gGcRsok8o5fI/mj2ocI8JuYBR
w27P4ZqwTW8zO9qgnv6ZDOj/h3oR87jS+3UFqMRLLWLxfA1sViPYhBJSmURVhdOs
JIq3RkQzumh13oeqH0ZzYJrduxcyd4K0055cbFoqw5NK5OT7Ft2+vpVmSxqTxb4L
TsszDD9SHikRo68OqAcmlXN4kyrUFCpdlf8A8xmbINl5D29GzAu02F29btJv5YtQ
T17nbFpWd36KclpW5PpchwDzlUe9F7THufi0y8DJNkCgpWilkNyjzzrdpKwzORi/
IFyB+OD4upU0TNuiUslVHpL/VlUrqnnaQzBXUuDYCXcU5HLAN/WVJRWibmoDGz/5
ywTELAzKI/MJlJ4x77xWPGfxtM7YGEeKdBUf/NWNQxZ7rtU/lD+X8nnegE5yfIuH
BkoeFR7bXIdit0dOOxUIWcPlOejhlkG/dmtXCGK6Yq4BacVi4LxfGf6Vnh6w+sfO
64LGDd/qlwrolXwrLuQJRH5ywwuIwCM8cRDJC7jgiPgud2ujmDRIySUzFWotKgFJ
tmWZ0o9p9ffhvgjiykQ1Ue76IBNZJ5AbbWNjQx0hXf49o1gCWHYDZfcpDBMSJ6XR
zuQHf3m/soDd+V+f+NClLXafX18EknNshwpzXjzBK9YmQeUhZTnKEqygThyz6MfM
SlkruF1HSy6PBVS4loD0m5eKLH9XaXoFiRO+m1J9DRItMe3WHi8GnLZEE9n9Jhgd
5L+tkQsLHp66ba40nh+OEfic3P0wiToh012crruMU3XDA2N5iZhUqaAP6si3tjlf
oGoHxaS6wMtPQon3KnDYEsdMGqZrSb+SkD4MQouB2SimuIPoZaEY2ZPvN60u77L2
mXWww8DFSJbbyIcYc4Uoawq8EzEp2wJob5OMGvrUyL6XIOpWfx6PAgguDXwWUnLC
NwC1r58v/9/BTw+08IE8CAB9qKdFHOmwx9jlR+5xsl3bpU7/5OKlGxa6VmzfyyjZ
jyd3157c919xX27+bIb4MVQ6R+i5zdVvKB184URvB6CSPWg/EK0BE49X6r+okx9o
54Kg0vJX9jjJsNKhjUN8w0zRtIGQyfiWo6x4UbGBDbCLDHMbV0SiJeLL3Kp9GnVd
K3uLp722GwJBZOf+7SsnhqHMGfVUZJmt5ufSAy7vI3ACBrENVpQbvWg/8Y2eLm2F
tXcDui+OtRuWb7VLiooDUpRHpmKclwTpzVTjVSM+/AeIRB5YhVTs29d9k2/YLK4V
hci7qz/Eq/7XRgPuuFrThq57lJ8knhac4y3N/7XTTtpEVNQWL0PppFrsFTXoMz6K
i2Zy/umkSapIXzeR7wPyM3Z7+eV2mZ40MMzXDZIRISuc7cWyA3axGAaic/7j/2AH
ykYF0+z5aJvcQNMv7Wzj4qFqDQgr0fpKNR7vlIT3UzHTL7CHuOQukjkC515FOMSQ
m71eFuqhdfv2JmRuvGkLqACYTyMYX/lR9EhPeXcT3IgX77J2qyAm0x2fqCetTSRj
y8voI12SbpY157VuqeJG2b5i3dyoZx2wOM8JFj5xuyhR4/OEgkjUZlI42NKhsa+A
LI8itPufuh1iQevwU6ljNeFr3CbZhabNPqPpt+jChwK/4F5uU0pigiSOfpyp95km
LuL5ieywgt5N3kpYT6G5MjW904WZ1x0LaQ3bzoa4k4l6zxCcv8q+YHvx2Hp6Re9y
ZStHagyFiOyXxD7HhGcEtbEPDsc1x3in1Y1UtflEoW6qvO0WGNuHVr4rQKyvw57Y
kcBhewEIC5Pmp7J5sFlYubxL4Ha0kKW2cVBexXsowAVO95oOXV/TRDJ0C6lTwbKI
BahH8XBSZUKMBf4SEAD2AxJCEr435fPnVxyEaHvjid0FVFZRxi1AoZa8fUfSibT2
Qxnyycseal3UbiDd2TzED9x3qcmnozBOuQ+nPMdv0zuBD9p2DCivpSuRTg3Z5oR+
rj30Ud1Wu8jecmgojKzmkWGvcMpA0Jvs1/ydb28vGgKIdZo5aCO3jkcWxxJS+pP9
u8l7XQvyYnjb3yq/g7MV/ASM8Bli2XwE5WCgjxW7b7VPKo8G5jdm7ulwhcvYmI0y
ic2uHmV+KbpKbUUaTmJBn2SRhHJyk58ZfY3B+m/EvonSaIl2vitaAA0qHf/28W5j
g/GDklB54HnW1oyVGCGlE7mdIcJBXNWUgVEokojZari/bE4CXq+FyN5o2lATcz+6
KwMmq3Acm036trKLbBTTvECvgWdRN9CP7zigxmwIuCggvabetVQySCaJaTFtu4DV
q2epMO9M45v7EATKvnO/DbTZnNpw11Uf5cmuORMS3tcQJ883ZyMvn/8jljoPUg8M
CfH+SENLsR+pSj1dIH+UjJzpa0ixy58XBiZfw2fHR6j8pMu0uBuCeUK8qOY2dvxv
Gtd0IjCSp15kDNaC3vJgkmgl9lJKWrLnDSp7SoPckukLnEL128unkk8ALGO6qgRy
KLqW/yDrzhsTOSg6oocjmjAWxh2ol0mqLXy5E63mRJdrxAGAPCQ5YoN0JB7FPFwr
8zAEUgrqE3gShce7Z9x+Pbfrbkum7qfSqlI3Z+Qk/XGfPLD9a8cwPP1MQ4GNzWM8
KmXoNW5i0+4oIs46exaAe1ROWnnTdhMptv/RuGtxwGiVeqS8It6UhBpUPq3RmZ0X
8PDMq9SWBwZzHhJa1DKHFSVFAeYZTC2pyh1LcK0ydva1FoQhBQEq1gKwD4vOQNis
VvfZfEiZeIOQA0Om3tpKQJkfEhwqGF4neAOjnfWY6mBab0txVHjnJm5FvhC1e2wE
m8ARquj5aCW/TPc+4FW0/XlkvzZ0rRRamGJ4w/av+rjnB7keytq+MzVSeqgPxX5d
cP6njDPfp/UiMWysIujVI0zCSbBxWCrhgKBQzcPvzXtVeoy2SPDhXt9He01GrnCZ
XkFsEUWfs2jcgcpLpznL/2v4HgPLnZpiZUeLP2di+W+RTTsnVWWZAfMA1MDs6Bnp
kDUZDCGexeCi8AWNuLrbatQzjut4yxP9QeldATk9w98FHwAeCjyC6ZCRslH+BhgO
UWmOLin1IUh2WhDYP6BFAK7vVFQJI4s8PO3iQGZPj252VVEA1Og8VIeIhpQpkNfL
Luw8EUsefeCXZu+9BKU0t4HovAMKcm8R4LM0+3mvj2tNt4q4lco6u+6w2ffvKeGu
IAx8+kUTwWcwoYhUyxcoIjNOKfG3svixcsR84gOl0sKBqQ1eZWxbfhB3YbEooDKK
QzroQFTJwAzSaz4S4yEbOQPP5eA94Z+lR7EgdY/1C+PJJOrj4mh83rzDr3IYTZjN
7z1BcrqpImvycNaehRBbyVUGi6d47MC3MB8v5nTj1nnDgSvKWupagtGaHngTXBZC
4zhDK26/th/JdJse7qXRWNCmNj0/M5ajFdWtVPso9VsVO1019vxDHb4a0W2k4ymZ
v7+Vfoi3h87vvZHXPAZkQWgpfuxMhJNwMMxecfZxJ3SBEGyz00+kh0upjUI7XgB4
XMT1qyHBGmnEOWUdf2Hp1SZlLjL3bcC0HZNTq5H/uzqFZ3JAaCLbN33t0pP33cTO
6Xfcpuf4nKh20/w0NAMPvtdBr4UX8Ukd3FK8ejk3+0lkFcBF0IgEqEyv5jALRoBX
51j40iYnH9kHaJFmiu5yM5WIvBpSyDwFYqlInfFKXElrUBJEG61p1br9G5RgngXg
v56NjO5S121i7j75Qz1BDb+JWZLRZkJBG9MrDyfHEH4zem9oOphIn5e8Vs4ju3k0
oxAIN/95dcNpxBTgcpE2k4FlXi/d5eZYYrVOGRti+87NkLQtuK+xsAr2IOKgFgfJ
EFDQU617mEXQNiijOeZeJ3vUU9EXOiqdAmxJUu781qAka36zrgagu76RmUz8t2pD
NN/AprOw8lfVY/pawY/ZzQQMhKwR5PAhskCFEWYLHFF1foAJPbRDk1wv1dtyv4qu
9nrnHbz0+eGNeOk2IjAnUIbmzpVeHUF+3bpDtUGa0FK0RI4jvg9C71ncTlhHf1Ox
j4RbkpcQ53onBfrGxmye1nWnsvK0nIncMa0XMm+UkTg/HnBCKXVTrtxCHpJWETXL
eN6GFt5+UgmaSFwsisMm1+JbyAgOX8bbSATmT3if3tHX+A2cmE6PS2sDAyae95AM
IDJSAFW2gzYw7P4OdzqWsi5gYRms5xJ1CwQx2BRs6QJSQr6tJQUeX5nZwRJzeddT
RtdNXTtQVPzV+/yTNtoh0PHUZVbkVeGuwVi9I3mqbzLqtaMGNFVyREW1QrQrVapT
qZ8T43clM2V5fFOAE5QIAnr2RItIU+bWcI7pltv2QMlp/afSejsCdEAhwM/gnKTP
33vVSWQzTbzeQUl/uK07rSQv6JGHo/PPzd3kYDlY6GsCfj3Yj68yw6yULTuEBtsU
0GP/hJ7MwjbR/fzYPsJQc6d+YXSX4LYKJOPhVoWEVMWQiza93AW534TbqVU4FfFu
ZUcxIURhmAJoR7JZh0II3RFdaUz4dCvSW8SePrib+oI3zLYvZ1dkcNRpRjfAFnCJ
kxuU0T9ZGgjGqwdturCNbIcyXsob53SC0OcqZe0gA1lrDnmTeQT4Qy4dJ2AQyOoY
z0JJU1x+6TKYDfwSPpp8g7TtpmPlM+WM2Hd9VyMrVz2HgkvtgE8qVh1QDkpruEex
r1o7nqc5ZIXAEvy3schCvSwo1N2RpuzqRwKpZ5qua/rn07TQFZ5SRT9IRhAwTkXD
FSzrs8k02wc7P71v3lUMa3iA0TfyNrXCsyoV6qY3sTBwQJ7SgWHhh6JciF10G9Hs
8L4l31qdCbhA5SWizUomPQMPNFcdoc0LCLji6T2p0nNrnMdGF4RUxLVsTJkFtxLv
30gXEcFoPOBuCbdGKmq97rJL8jNADbmfPeMfR+xFdCopFhEbRVHM8L/QH4vsgAGY
mr6q++/5x63sQ4TK8UH7/4mn38gYIbwwsQeabJbWnwgGS831RCfCDe+oaVtcc6eO
dr/dat07AUB/XcifHlZujQVaXb/jfUylcAhF86vLuO1zVWmaDK/OtPVAezh24jsS
uwhYegayvC4bdASiTv1Z7GLlsOKn7LOIN/GqrChwa7DN53Gm4flnFVVAvm6vYREu
ALViYMLIRG01PW2PLfsYTqabZUYpoIG5uLQP8MZVxAGseq5FgXa/A6UERx+VTc8f
j/8m9AMNaI9WSqsE1OChv0jDxu1+7QjAl8+FytVT0WYlL1X2fow/xgzDd2tbIYYE
4+KX5ZKelX9LAROOtabO5rpDclF31c8EdxdJpI8vxqZic/SEyQftzECBF6HDFGNy
2mGfLjJn0uX+sHlt9aBp8oRBJm9Vo2LibC/iQN+rwpBqBUin49HnCn84AfurHyjY
+hHPmojvDSdZIwLtc4f9VNS8eYHWV0X6c75dRw7v/O1gYeorkm/yyNX00zg7nJz7
MMP0cEWHDsaqZY3evo4uYcaAmJpeQrpZtiNQGmByewJxb2Lf0c4fIvMumXhWwmRL
C3E96zw5oaz9pldPfjc1avCIce7H/jtXIDywrGKfejgDfXYOQQx60ZJKsHCA6rWQ
yCpsnlybWDOkdxtF65qH/x/jPj61YuvZ065M+RChhO8s6PdjCUwliNnGM9sSpRFh
XCQwBchFUvTXv+VLhKpes4vfD+PEEkoIu55sr462xvRNxbn80x0N6kMI64XYY4aJ
Q5PUzT29RDphE9WiejcN39Uno6wuFJzonprrSXO1omKQknARH9nZCG6XH+/g0sMR
+1wL/OzQCRgZ/leB5YAHP8nQ9b7BvJ+IN4FJUiOk+IeQxg+VuYqqRj6joROthiq8
gCyisosTq+mfgzlFLFypMwkDZ9Lm7wqVZE4aR74CkrntPHSW++7srdbzM8Qf6H7t
X9Y2832PlKyGKzBZknPcbD+owZrLelNZwi/FbAk7mUTQHK7rzQ+NLjERA/xM8tHs
duGfvTnl1crzcf4Fi4J6bhUSW5SVdm2tBRjvgvEJ7Mcoa51cELi5dthuzrmf5I1p
WvYGjDNI+I5o8vQ3r3afEKpQ1y9KOQjqLei1mDlPeuRAa5OkfyvNTjvbVRsBxYuB
zIpVF49J+KgQKcRc2bzqH7EtJfbJeGidtVMNXDHSSeWZOKo98uh68OILpwKjkc2V
n6lGCs2zn5FxJN5fCsvt+Uw3tVaf+0iwsPz8pgUQb7OyXp+X8OYHHvEDrsM2aZKL
DYY928VjL3gjlomrB3TvEVZBJi7234+bi+njQOj1noiswRGSdOzU9kXoZOWOupD/
pCvWYezYtIgEdC4CzLq7barx9nOlwkAaTK8/rgJMjgTg4Chr1sxFiuNjSurdzImM
OQzxohOwt5EqX7rjB+aDg5qGZ7fzIemyE6rKiiRUHwvxRe9irnn0Bv4s0jhMkvOs
1EwcFYOUJPXnqQANN6zmXlItg0Pg/sEw0XbRoFl1+iuUv5LPCQMgtZPbyTneXd5+
4qdSQrqI9rHvSXte8W4zwOF03LN+DSCNkghT9yR7jiyApEnZ8PNPUUTSyKu8mmJp
e7sVfZg2uBL02XtYBZnrL9MWiY34NrgAmzkh9rNPfxSlYCy5eZI8Pz5RmwE9UFPL
aUivEcitd2oqoER9f0AtkDF/aJSaZS+CrS1vVcWkYKpgqHPII0J+S8lYz6nfLRIO
0rUXL7PXLrlC9QyOPL3wlvklJW1ulY51E0QtU0eNNJ2xLZLYi4AOv6jbbIW6ADKL
QLHCfPrUHmztK/IiCEzzlR6Cs+FTp7ihmGfxrJC8OSf25E2HyvrJgT2Zj4QiTtic
+oOgdpqFYTj15IbdknBlrPlVgvOatw8FCNZHM8s+r+glinQVT4rwWozRa4dp/0L6
ZJNrpKSozvaHeHkxrCVCzNKyQPVZHFS5qeq1vF1dh2eN3Y+Pcw/gOSgcdFVFBRca
LfepfprtbH+rLK0gIXwraajC7Dx1Kc/4mh+dEDCB8nAPdH4jJOgjO4nZM69IOLYU
GeoPkFqnzTdMqqXUEXw3P+egvkh93jdhwrW3uqqujn4KAkdDacMPNzmhMzap63iA
8INd4BY4kEVU2X5P0RJqWvRcQSxD/JX4sLvmjKpMmknOmqGRNJzA29iJrEDdjMqH
dNUxUNyqHVh19MprLo67nWZQESnUEiv5Xy7WGJB3C93OOuvcsN6mHnWOzeRkLw22
DmRHRgU8faK0/ZIu5OYP2glou9KSM0OEerff68whd++V7BVoMZZPUbpMSf4iEzI8
+qNAqfmnl8lUlGEZpoIoxE37zOQs8dwM/U8m87vos2E6/kygWcqp5/aQUoQoRBMA
Epkq+pqND0FXRwLFQTq2RlulY8vZTGjtsksinf6tVeiK2Yj0g5kEH+IvxVtTmLjr
Ov+eAYPltx8dQzaaH8SSaK/7d/nU1lZ5DJyQmAEQRZzvQ0inrbfU27mzXwgkpwsn
2/5yhaU1HpzEgu6JBK9Z99fdur6oGaWU0U8D9ZMVSS8n6DJOoRvx7XJh5raJ3Wlc
5wk30/FksufXhcCkF1ZVnatvWZ9cRQWqVibQjs4M4tXUMkfNipY2UwtoEr9bX6LU
bgihyb/U1y4nh9yoDsRVlHMuuqLgxkiFRXGMVTIKI+gEEEcNLwndG2zXz8fxQQ+Z
gGJ6p52KHnSHVg5SgdSaAUSns+j9Uefv7NFsd6a9hr0XTCC8aa1gRHFvUQqfM0X+
ZCWkXd2oitl+9u2TiM9qprZLMfNkCgl+o9Si5CUt85L/zRknDryERxxW6ujzEqwk
yMKe6sDFSfaROzhcoJq7t2O3ByCmQudkt5ccN7oAIE974T5U+EaVKf5bb27YCd2I
iBqRSceLVOdQwnEqVxS3ls2Z5vg+Rhz2GTATdq0W/7B39C5etnDXhRw+BfP/rQVg
0CDFmitpa8E1S9SYDg6tKW4v6TKczK9pzydjzxhbADb9FaQhY8a7IFdTXqfmDIUV
CbeR6vNMAj/HTqO5ar/vKTYaa8DZ4HzZsF3S+F3yfqvBPdHsYbVdbq2JnrpOACDc
A8JkZ9LPp6wgs8ijzRfRLpJiqTJTmXScVaRS73WsAY1+P1JsXD+P42SLKVrPQTt7
FJhfWKRKnlC95I9VAx2Ms6Pc9Icg44teCXxBN69UeMX3WU7gHAVJnZE5zVHHATJI
4v5MbVw0PtxHIfaMgsowY4NITSYjyyWKfzGKzqwqO0Y4gb2gZUVtdhg/m3IaF9XI
aaCwJsyk16r/qHSYmN/6GcevD6SjA+TRJm6WObpD6Phh6JMNfDMx4+sJZsJ8hn6U
5M56Ab92cKx0yv9VA27vYrH9HjNpZriRUScY55tZGDvfBoM1wD9PrU1cCXn/pZyd
dmgFqYN+TPyWEcg6NsIMBhp/kB+/6QO4RQV2DvTcIJ0t0mYJAq7uWDbeeJY4EpWk
RuiIQDGDBjAsEgCYDZQzy5dQ2aMBmS5pu/ABCZ/AJ9nOJ400cb/SxA0zbBik7/55
+AU4IHbr1rziGsdhLRx+vYKt60BU/v5ouHgUTTBTg20m0hOn+g3VMYZSHWjbKLGN
q8Iv+2ArlgLwx7ekW3K0Uis+Qiq5UNGRe/5iNpxHJA1Z2b/K0cVt90Z6EOzraMMA
C7ZO7Fo2/MKvfVcO+MQ/ieoxnu/MKZeSBu+fSYWfCo9AmBIdgXHL9XB8x8yfaCrm
qCLt+3A8S3PpOCVlEle06VCEm3PbgcjkPJDje2YXI3RgXY2ZXMykCSz46W1XPR42
6gHZcWoajkKKCPatJhP7Ju3Vl4u+5dbKGSOoUhf5NxY2W3c2LPZCewAfU1WznUtl
N/sOEVpeBjVGfPxh2HhsbbYqrPKidk0Fzno4y9Ma7VmFp3tDstg7aLTCSv2dbj5+
14Xi6sTnkIzk3thFYUEJhd2MFGIbY/IjsFaKLaS6egFpMU7jCJs6Yu/RuNjkmuUr
257VBXvu0Wr1xJTbrcM7AuV6pJvFvLQ7bNj6TQNQxZQ4fbJ2kqG9u7s057KKtaTb
SNpRrW8+hw+ki8nmkEeoc8mEYPNfOlqFm0RoG1OvELfBs007h2gCNMt/KplCIziJ
Pha1v+AN1fLyynTp4GsFRI7V33X1BTKZVI8gxKsoQKP/Btlbo2CE19r3bh+XElEB
32HoTJHTJ760HKwqsP8oknuA+mLYl3XIF4kKOS+aaUz7K99rWxmZ60u6me6CB06k
q+yFq7xv8qdRJlzBFdkMR7Io9OQyQRfRHZK1LhPeJClddPwe8YjIdyaeh3Z+hJZX
4GFIB6t8JpdnlAvdAYaUPtzBTB8/2FxhaxJ9GOGG9kjPbZkvr+r6CKSrUB1EETvV
I/XE0qdLZn9ueklVagsH8lMJ3QHxKFv66cHVHnglZ0PXTGFYL4rIA8j4BgXJGwpn
Jer1BXDYHZtXprL3vG6f9EUXtO9K9UG7Hr9jXPNNusD3LkUE47NZHxFDtVEf3xpN
DYYQZ3CeG9Ul4glHT77i/Y7Ssx9WjIF5qkJJZvzexxOkYPE/pilywIlCLZjSPJxY
Vq2QGtaqDaMv0kMNNvsQbzy+1d1u2QvIRxCvqavJcU0Nq4tGAMOS18k4rBEZ4aZN
SrfZBmszAWlJMyEJRwDx1XriiEzI2Y1hG3G4uBrBa1xhSrLrgQt5Xz4A/CSnIKTo
P5HEBE+ZDzuFQ0OL/d+9HaRjYdzUOGluFwbo5s03aztRbkirBnnC7lXUJ6vCgx9R
rXoiDEmOQfdSx9gW5OnL4TWoy3NN2KoF1YTzMDmw1csiwm2D47iuvQM5ystoP1z8
fhhnhfKR/AfKDRoZH60ru+RiXnJ7+6lsI0Hoji/vd/eNqa9hm7H8+BaePllJ/CaU
u5VU1hbQwVJ4X6lKV7wrrSReqcSh0WtwrPBn6SkFRrT1mHinEw/WUgzWg/lNIOhc
17r1alnXkShINzslH+HWYo/8VemaUE10Uru5YsYOx5rY69r+ftbe0gQLqef+r9r6
XLj1rrfUuIdBZ6s8ON5PM+q/0WohvwN7j5KYNfSp0z57SnKtXO9Hpa782+ELCif6
hwSjBSbjlJ1OtRyx+7IcwUXUMGN1mDpI8+enOYkAhMMOJ3MePkInmqmeB3ChSvQE
RRVFVKAQ1sazVkd3hiHQVT+CFqmzec2oK5qquubBGla+k/OoNGV2gKE7BWX820fh
oIFaWP07ffTratcWp3dmes6u0ABEejgPS05Yc9SMtCSZRR/9LwgUKDl6C7IE9Vp3
SXsblGXUwr0i/oqfN+XYYAGFWsSOBbrJWgUkJx/fe4gcpJ8eta5LdlifEMsQ/NXF
HOVPKSIKZkloaTHmLYl6IwyCF+Qr41Z8R6BKpcsD+gsIelbiGf9lU+1TT3TutA+G
tygERGJRubChEKLdAtM8ftBQecs566wIKdyHAGOVn3Hb8Y9rp1GANPeHNNQsX+Qy
7nuQaVb7jnXZ+UMa4B0pCzJ9SU9CdvE+Ae78kvFPY7uj4ObrU8NXZTN5cSPPCHOD
bTd3CnPpGiYFqPd+VWLOhTLjaajvqjpK6+PuomlNZHhZMb4vei4Q+vrgPTKuzGW6
dre7Mjt8HgZ67GaCjJI6lPds2M4IdLvgZBZG32dURly51H/wNa4Ps4BQRBCdUar1
P1GEcZpobVZiTxBP/uCf8xiwPEbdeNDSpNZjD2Um98BNBMNwbTRQgclRWUZFSSzJ
KMh7FIUsFfYZT40DU/v/exkPr26Ootvt4m2MUfa9J6aG+orN98Zwk3MXnUegtr9+
B3uokYHAVPX2yi4k/t4CcfrkyA5YglibVRbSd6HqU0jmL/slGYTm6LWFxQSSOZ6i
AgykDDu20BFpnieT1AcwKydKaSXk617AwAqV1a9OSHMq7WzXP9QH5jvzLU35POgV
uEpOs+LUScdiaAh+4eApwgfvyw8yFfYD9XMfRMh68zQkdBGU3kjL/fD5SkapmDOY
n2U6j3uVeIUMi281SPqecUVuTuCaoEfgP7wCnNIxpzcL49gfHHZNKkSdH7NLtnlw
Hv+11P0WhYvXb3IdP8XMTBOpScp3CdYxKor5Vl/+OtCZ8BRZXxI4pV/TZCL8bXjU
1hLn5ihDl0wdd7qaKI27iwBSxsbLV374L3MpZevHMMTguFCMflv+SwaCHqUU5MmY
9ujufXOUJIfxH5XTSNMEZimmWnQzIKvDIZpEFLt/gd7n3HQGIMrBn/8u1OktnGmr
TVA0KK3V/2DdxbuB09xXYUk2S6hYSN2606cF1tBpNeltRO9V3YcZYNAvOjj3Lhj9
UEgVJ2hGCh+jj457qcN9G862lb5eagmPNiwxj6g/SF2TecBajn9z4BNwC6lCTqbn
Hi9xr7FYqLKqTHcrNq6VDI6sRf/0cgi8jSHVcXVTGCRW4Wq/ktjY/rauvGPQmyrc
h/OfgSV3QjSAMkHNJpwHtZH0lIZp9WT+iNr1Yb/y6OajvHxzSHlxCUNu2WuMYXj9
BOz+9cQj0PSo/RNYRFqha+I6HllchtLal06lvMYe2bcfpTsvTk1ZVQIWbcM526o7
2Rb+j5aQae5X2xj0nRuRfUw9S0XEHNwezU3vmQPFTZYDA5kKwEX2NrhOdRO3eVyU
uHLAy9L5P/f5jB/aICe+QlaEtY2r165iB5bOLA7uF3CKulZbwjkQYhkukLlqY45U
qB/fUM+QcFxGNRA0+Fv0E8PPU4Vn5I06RRgdq6FS8Einss0N9y/i+1QuaCV5QJng
r/igvNwd2VmSvemzb7xBXwSH70caGlhRlqA84XHRXuCifEltyQlEIvI5PSxVvaRW
KxMRws9jOMKa1LrzZrXQbM3PqbKrRxhLBwK9DUr2enlRmQK0/B0XhDkop+8EPxwN
WY5d38CD4lvv0jgpiJUHJicavHkKgqakV7r1+ht+hwkw49Vl7gVfZC8wA0KehDa/
f0VoCt69yfNLpret0wZI863bRoIuh74+dPVTJHQxZjlGNfgiiXPXZjbq+xXD8CGg
aZE0jOy8t7mKuTK5vmrtNeK5B/l1TVnqQ4jzA9+whR8G6dBH4kTgPwx0+Og8tpUx
HykHSfEdQC+Tk3dV3eM58Zr5jZGlwW+randTdJq1VSSYWKkLpfW9IodaGVNGhjRX
3prYS1avzKjWIIELONknkH1mXJR3kwtaBQtw1V09DIEbBEOYMB89RfhkBWultSow
wFL7zR58fOpZIFqJX2QkKUgmouryicENaGgqYYrZSF7iW4cmXjFR0akWCaw9/YHn
N/WvWBnoYDnkShUAgXUMxCgeoGEdylELciJ3QGIAtliIp6HJJr78O4rYUxUlOZlV
ZPZkx+p/1KH3b3iCbq+9rOLxLj0GDuQQ/g4mYg8uiHgA9hjeXy0p8Bs9A/uap94J
EK0ZCmOUx5F4LAX1b3zd/zE/UDL4S1ERtO3EoXf/uGQP/+2Qt7rM2ZhgUC3xvnDy
iM6toBbc8pF5iMPmhWsj8DJeb2jsJy8JWYLfMF7PDXPqemPlRSSeFYLZuBiZ7cCH
9m30AAqkGmnyBANjVtIlEZuGyG6Zbl+grc4C4pwvA0vxWP+eg7lacHDp6Fd3+CCH
P0mUuXK2AJKeCebBM6RzleXUXEpSs65gcyCVFiDnnsXf5tXzamMV4IR5IUYML4Ll
TmenqNTANOaStvAbGJQ5Zk7gMoLti+2I9XW5y8SiFGdAbZ+4qMrQwIfSX8+Trqh4
5poUa/Mbacufp9NRq4YkXVeXBlXoTUVMZM+ikpjlkd64Q8DeyrWFmAA57yFVSobN
zBgOuvcfGAFEGW+H6wKeR5cXrJZQUVAYLgElj4WNf0/wNv84665+jcXNJECtvJYn
97cbXMMxMeHrSSdNDMFj69pzI9aitXZQHcz2qaKwRf1QiTVWqIPZI5SuideLrxYf
3MEmdt14M4rzDphT0N4k7en6kFxgU3E2/QLuF+1o2wTiIrtPEMEY2/6Xz3fFb7HY
OEPI77P6O22KAgDLveDMpgvPBmrq8C8slPmTTwJQODCILjpnkXB2zjB1XPuYNw8e
oHmL/fbiBUDrRCHFLGhZSLZWDY7xCF78scPrVGdYmLMUnzFw3NtdoKlJjaasUgpC
Dy4wO7o4p/Ods8rJVBmRUl24q66WDirFJFeGjx5Yi19wVwLf2c/6/kLYpveUK/he
AR/XP8Ita9Oq5Xhfgc4DS/UllJqD2oAOEDx48wOGy6o4tfid1BMTm/IxU0dLRDoy
tp2LFJySruGFMrbINslHTStzsH3KZJBZvekye06OFvZwPUv1I6J0tuuLMP1th5Qr
e/urhFE020ccNWNxl6NVb8FuljWx3YSKB8lxmfSNK/tHMXFHBQ6L2NhFxZGOPJG2
mdcdt0S3CQZBKI8YbhiZphwYAEriKFTR704OmKbaSfb1L+3uasTIGvqRhEFjSLAN
i5ADNy+LJ/UrGMrQnnaoDe+1BiIS+6wO5HqYDd8lZvvYHbCLyMh/mkrXm9hk4TbE
0GfHDUccM/Vfm8TRO7E9cADChBbWEkXddoAQ/to1uXvd1bLLqC8sIjOzLSY+EVKg
NBt8+8+FpR+xXRwmC9y/Mu9Dm9Uw4UFnfkHMxm5v8cUkSqgZLoMEngz+g23oGCyN
W3ACuWdj8P1DqxJ6X55cPJlQimTNmlGe+cvNvAbdKfIQ//P0MU5oqtS2xrhHIPff
MKp3I/V2qyhe9qydp4mqghTOSY+ctv2ZdBl04akyAY4hL9CbSLHDqwcx55xFnEpD
4EPLWd2GBX+qqmbP4LncT1pvErdoRzr2nXBHnTvfNhSJ24SxyhEjgyD3NBRaYBGx
TP5Lr9Zi3L4jlhAOcsEVm3aC3F+0UeyyuklViT9soJsDJU1oaPv/AdUZmHpGmv4p
zIAZTPCqlDLyOICOSCR3XFNGdJjaRJtLtjwF6IC9WyptWr/5TK4AMvSk1EZanjob
rAKxlYHs98o9/+Mz0GQRzOiaIwvdk4z1yJRx250rU0cWB44c2LzK7XVWRQfLTxlQ
T4oNk7S4roU2XGm3/NSVX0fZOUkMz5GhOjMtgM03QJFb7D3cTNp+X18MVdYjUTgV
Rpwich3EoAUZXLzjen5tf7IFxFDKdJrbCRbYP1NYvqullCtLrQs4ZiZvjGLfqGEG
mnG+wtWCox+kNEQCT+k+2hlvt9q+AMiF2wP/MgAF8Bu5v/ntU354tmQvLJmRrVXr
J51eaHT9mmTzjwOKuNWSNcAVOlugU1BOTXTOrxkhxgI+AN70fHNH1/jH+nAopzCN
piu/lhKLnAl2xvTny+ypM/EYaE4oQruXaCjDSqvXZzO5XEa+wDW6CRm9J9j8DBLL
YHvV9bzXmC/oUV0gAWYXxIqZWNhC+ua5IS46CeZRl/YeT1hl9T5YFfqXwxawOzFr
XMGZOpi3noM+cX+kcSJIz8NmPMKSBajcGyyG97K159uOtNAmhy932Jman0pxpzTK
q9ptp37Zy0V0QA6xWETGFGLcvI1RPAi2vVyXKsQ7aMBIk2h0iN3qsUUzT9jvt44h
slRPYVmx1EyPq6KB3klOeVz+swWNDCD97nzLydku6x72M9yhuYtYtS61RWDex8Ae
uoycxORoq1WYczrnImvgmS950yPsihSLLkIimfISUdKhAEqLrgsEwlOWr4iZqRx4
93pMCjdIZD7DPwFzKt9va1psymsj4e5jIor+OGxb/irRqpynV998y7MjWMNpsjTv
SZQusTFYGXW8lDegyDge5QZswSkVzikUQosElBoATYJvXNF6vGygn6h8oanSitXE
D7cJCOpHndT79RJXXrHKJ8LGY99cwG2M3VvoRuE9RurBfAChWnsMLV+BWD0kHOue
NwZh5+QQ35j6avKBrPSUIjCP7X68AT9oKlbIZjln6Vhd+7izSe8/hk+CbSm2CNBK
L+ctzAqcEeZE3ODqH0puQwIZ44hDRHEt2JXTY9KvtCY1Abdh3mAtJnIr9g3hu6ga
dlfTip1QomA4HYbB5CXN57m5YEqV7Opm/ALk5CLX0c3QZ4E7YBQcNqkjHfhd7poC
w8gdRFslqp0yM1XbcG16SLIsA22xv0mFmbQjvU/SpWUK0poT2PM6u720n0SdE8dT
L4Ix6d1l/+CVhG3BLCStfgoLcDSuIUeTQKssXN2oF0n9uWUr9sxJOrqfkxZoY8fO
rrgV8buW0ae7aKCDQmGcGm5BdX5RgoT/H7Gvn7CUuhe+jdWtFcTjTUd1vKVaGWOu
hbfruEvtnY0tSI7FprxzWMfaDddqr90GNJik2x765YS/YJ+toSP3J7wgeLbj69+B
bzxvXIaCXxSOa7kczC4bRKOs7fvTsqH8z8r4/dJa2nzSH9pLyY7TpKatF/BboB9z
g1bdCyD4asmv51WDw009HJ6a+HHXVadHKp4MTeADLGBiPEtZJ9c2+AGsyDgcTV0T
G9TJzU52ciMLKhHw3eV4QkaIAbRqBnJ0LnzrQ19CPCueZFKLuUTSlsNwca+5ilBV
bjEIO6spEAxq+mW3J4v2xXqRY+AyxCnUFy0nLhfJvVKABwLlnIVqlCxu4DwVTIyj
jZFCkp7gAhzUP1WRWZKGNh44Hk9ORjl+DvhAuKMQ9EXAejuYXVIoRdalNNdEbatl
olODNDhZFdt5Sc0GSMFS01ngpOmZIwm4boW9OJEwXCybJkiWbh6L6THXpWFnhGyB
nQjF+XniFEHkKEwLZdh1BsQZtnhzxA6x82Lz452Z7S0goIHnvko2sRedJKAcYxQu
KHbdoFIiQuHAwbDBr9P6o8hUpFkaeszv7UV0DuTQLaytVyAGolE/lGGlJD80D8d3
yLx8I5aqtMCw8+LKhpvMMxXL6Op9Hkor4c9FqW0kV8L66zQ8sLILHcam4Aq/a+sC
oASxTzWCoRJ6zu/xzkk8yRraqPc4fLTy2+hk7nxL7+r9Z8CCOcyWy+/8d6gVB5+r
8Vp3dVnIbalCvF9i643wBHAMJ0j9/6D9PrhEztammw+LAjI+ggB1+Mkt//7Ewms/
OjZBTkbGeLPici9VCJpf+UHk8CW2pafrL7fK7dnb2M8Q4r0ny/sr0ZNotQ5QNJms
dt/cyOW14TeTKZCkZHwy8OD+VWEipzfFAaDyV2oVdYwEeuTDTW+TL7Dwjph2np0b
T9QPZq+84LTIe9/N33cwEmIl83gR/Ek62v5K2q3HaFbwiAcav0YJ3BZEBsECM98w
RasrZuMFlSBINatQ+rgDsLRI1oPdGyGa4bFY+UzjKuFivKtGu7QuVzjq7sgFdzwK
QG8Q20bHGlQVdWejfECyABSerhEJZvMKYh1EnvCbdejYrIa6nhxKSbxk68mplwOx
qHQtbK4O/pbfLn/++e8E9Lw75M56srl2p5Dg6T73INeBSMqBj3uZweu25P+a7iXL
hwLAxttRnVaHc3H6KHhOBkCeG4KedVgXr1VIszKvd2a26YT3AAAYANsMSjSN6j+S
jdC7jzDNgDu0YedJMwIxp5bStIDNyH/kW6aKkCnV8GVRPKebjVxoKv+AJLlkWckm
rPcfoE1gHgTeYOKR99IoyW/ysbtVv2PhQbilXlXNb25Mtr8b+cbDVN/exjpFzJ5B
LsR0ypFzQTDzA/5FNBrf+pb8D6UsKejAZ/rOezyRa+GGjLFxifY6l1is91clVz/6
e/zSCexYOnvj8k3LnT6WKWd8y3aRVFtxRIbH9Juy0WssPmC8B1uRxVrJPdpBOfWU
DS1PcURBXxPE8naDPEqD7DEw1JoRQBaYQc3NPnW02wVVw/6zBfqVcrtRGADK1eR9
n3GKe3341gpSa6J8zpuATlEcQSyuiuTQuZLupDqO7jpn0lWPdl7PZRRZydixCS6a
RLhWfyjrgHDv8/t1N7Yp2nTU9fZ/emNevSjlSQFVc9l0UoXdirKd3xch7rcg66MS
DRfZWRsWxAo0MrqWNMuodI4Mgw7hZdmbQoVmGZkX2ZI/2vvwEafdOxz66EEjuWp/
fqleqK20ctGh3qqdyXjE5wk1zLYDN29gZBHfOKZvbIFuckOV8GnWbSfKFrHcZCTD
WnngwG6K3y1RxiT02dXFT4E1tUYBZMBfsi4aFe5vO+4wgQxPZ9Barx5Ot0BNDq0i
aTr0HAkRpFgGE6oufmtR/UsRS7qF2xDO9C84/APxky+yFSUHBJksZf6mfnXfswup
TlQGp1d5Do8arFEq6MnUFTET9pqnpphfcCFoN3qJe9GtyfU8vNsknb8Cfqga+6Rz
A205V5cVb9T5cuifz9ZdUB3fDvTWPo4E+HUPBxNRRUiOR8kJMObPx2zVdSiAwbRM
1peHjXYEUyvjxWfyAZsmjh+O/FWYIDg3zjWV42HjPv4YNkeZHv9VDmPpmhg2EB5K
IOYnyQrnHlO12lTJ7RxNaOafyqOHnRK6nWAr4w1M7zmqePmpMHxDd/Kzq7ZQd7VA
6cS07PhZ0DHrZVrhsctut2DalzSEPUCbQT0zvj+yOEOkd+AZBQZGKWKpUDtH49sg
JzTdhW/YKgs3Kf2iA7emZtC6DevjSu8z6OB1ozqjAVyXdK+XF8GMed53igWJndQQ
SClX6LLPXPuMS9wsfsenP0o87Et734Fvy3hpk6Vv4ZhHIt3WPqeNYcb3GiTFRMV/
awDQfadmwr8a15Z4mARpFaJAvnMm+i4xxpBRrZzaUm5OI9JWL2U3PGHsjypF1yY0
xZxAIdcqOlaF0opIP18q911cp0HJwgwsf/IW+C1suEktzJ8UFkvxgpKfBunRnNNT
cxEBe3e0/fGlUBh+5bIZ4gW0dAJNYGOkKNKvyARUsiGSN1FTZ5lKcNHr24UeK4mr
wd0hpDxlJPeDBzCC8haqVJiH1Ugq03EI9rTL8brQVlwjgKc7bVj9sxZx/7AoCep1
lbNj4I1/z+Yv8cbbRJBmN3NYgkeG3Ajr+3X9dMRBkmCGIYgh9eHUzpJmioaWbjdy
KMRWU1si2atKwuEj5OWgo4YbMZovA4BfgMV1IkqzTxTTmo65Z9ia6vek+DvtpUpa
dq1plmQ4WX+43FAYCgONYX0s2UWXYr80zNfKzkJ3uFgyonkTzbwcUQevNv1k+Yw2
1GCUx3itlsTKs61jFPaPiCCyYTnlF4lHuf7hJOIR2yVVpEpL8CvnJD7TLIfV0QxL
Y671AJF/peQsplkXoAkY06kZ7gHZQ2X4ZWrpSCW6RONIPAW+fd83hJLl+HuKfB2x
iaOdSgLgwx4UYbJ6UXGrT28Asm2ZgGqb1/7jkaqTJ1PGdeVxAHLvZ/a87JJ+Zdte
aC0tpm0G3di/t6WuoLdnGFd65Pd+63Ak4/5UlRwl1Z0V/tko7k2f+cB2fDeUKemi
fq2jNGkKmXkzWgN+4JnIqbgpUJT06VbATsWjFQinNZfKlKn2o/s8V9y9verdS2xt
akQEYHBOQY1O+BQZG3gN1+hNGmeN1E+gfY+C7ihFO86ADDdELhmYEw33JGXL+PVw
hYW9PWRfE9BveSaVK9hnyfYAgSbFGcN8Iz9BlrLjtuCTDiNCyWyNnVD3UBE50gLa
E9bGU0eUAGqGS7XNGTBnnKc7kBvHEd5y7AW7FITUg7gzLmeBrhwOW3mL8Dl06cmc
S1MvJmBj6qNoIt0n5zetjdGw7LOnDg1AAbACgvrwE4h51+5kzP3wYlgpLhEUJL6r
yENqtjfCp0Z6jRAVn/hsN0+NG3S6csAlShM4fOia1dIj2qNSBjjcqcij5rhDiQvU
b7EhCBHtLlA2IUCWZ1fE2GBFNaIQtLjfEiLdWxmTmRba8snLjq8dQSg87iGMk8UT
lOfz/0Ww/QjEbZHXxXgcXauzkhy32Sa4/vlzYKdESAnR66g5qIsmqWIhZ3wGKUak
mBX4Bli9oQU6Ibs5zzT5CcmVC4aZbP4SXUafRJNksw0EltL6sXvXOVm+Fs3xFNYw
VRq5cwlHjs3EMqg1A8KVEVCo9NE51RPzlonMcCwaPxJupvmyFutynKVEmAc46Ijo
UxfC2ShlNIzYjd1lDwIpiWZzkAQxFJN4lcJ6AGflM4RIs+Wq8h3W3OEbxFfCFm3s
xqjreQFVY+/k3X1X3MQS21hLwV605wx2DgMM0Q73p5gylv4oc17FAQDq+MLjGYl3
ArZfFMqJ8xpT3y21aIpZuibimTXICgoB0QQUI2PQGL7nNHDyq2OENrfl3UuR2vMj
ACXfREblFNIVfJZSD+ToaypERRVWCQQ3L3AK3YxipAI3+eCJ4IPGDpSJYvrSvQZU
R4Z8WlKScG9HzWeT4rgMwHdrES5eFaHIlZmTLPYVXnqbAMriYyDEYK2yu2U15fj/
bzYoYurmGuSGxLrpg3gPRuk16QZioV8IqWa6MvnBoZewg0msiuxq3XSSYRM/nfPC
Ma4iQGkgqOj4snTTo6EqGiAwBU0CAXh4AcoiUKzOp3Wz9m75KMSFDp7VWLIRRypt
12ORZ+uhg+9v+2jItbI3I7+Hhswu3kaaNbtH/Zu++zbYeA9AxlXK1uG5vMGuorIR
0966G58PveJ/jizBvbFF+SIn9PNQGMC/dVYK9283k+sn1jXoYt3roYP0qCSY2bMs
WnBCkwdibpilqxNs97DkZ4K+WZdWQjFzO8zgbs9GV/VPR6+5Ywn3xDxL+GBksCym
yc7gxdjzO0Dm899M/SYN1A/JM+oZn4pRHMIDLRYlN0PekXIzrYwg7ZuyNOorrkW6
jXMWKzyDo2/Dgpd2/XLyZGBX1Q2x/UwB/NvxfNjPuVfrVNWLBTYZW0K5dghX3Jv9
MG2kuicVvvP3Kzr64deFNtmEeiArMz9tr/gu0vaUTFdDmZG8Lg6fJbtQvzeufDl/
aYtZXO2NtNOuBIKdhzUxLDHlcoeYSxXCHbeZlhR2YOah9ETA0h0W6mgcufxnvR2a
ztCAH0sX5IbrOSmMoTnrYV9CEz7qesGo6vHLoEX3wG4i7J5KzSoiV/huGS2+Gs9A
bnd6EGwZqBI1XmERrkkDdcjC1LYhlxEpE7/VoGAkNlo99QORJt3Q8tdu5zGaZ2uX
xXu3vdUQgwfd6HyUDvmxXm5p1Cegnf2pDAxsWiBr4mGAsi1Ext8lLFp8f9fpv2ac
e/QX6K0ET4QI9z6W4f4BHyvACKdjrjPKjOQnbjsm0Q0oVMoWC/zv97T7tdyMnioH
gwFJ2oT+bndsjixtmijU+rqVDTRCMAwVyeJm2fuiU+u/zoXyn24Mc57fKinYU15v
XUPZNKuelVl7XosH2kJ4Gl5CkEDdZtUPb+MNginq3Ma6+oc+/joa4v501y0a0tL1
GwDXIPsOpESCg3AVbdaPXtHi9rcPs5tF82lEydPH7F/8ED7GNr0icfnEXNPbekev
mW6u6DqZK3fN9pLF/7FwACz8o0aIklGyUl4wwME8YidTsKdk1LASk0jilfy3kWs3
Mq3/eBF9zjBrm9L4U0vee9jymJ1c1uwW5Q2TFFHXpB8SBOeYH9lbnh+ffAU5G432
ooVbY8D/6hXYe0q/IMdyYC3B96PzVEdizh1FaMJv8zmuNzgf2tfgjEXtE2HGJtn0
/SUS1GIY56SF3JM3BuYjmG9pnu4B+fIH4WVja34x6xBmvzmeZpVCULPwNfbzUolW
zKGB/daPGFBBlmvfarx9r77D5FWOtp+f9756SSUeKdZPavSEXaxANRGqeOYt60Eh
9yvniByV68Q76RTQK9uUI938R0YGKej2T6erg30mpn7TEC3jwy+z+r+runL6yBBm
hPNj4ZdXtI23fVX9F+/ouU5o7RAkNZqA2Gjjjc/fdMaBylw2FbXfmMu4dqhbcgE+
M7+SB1GZEZEwvcdP5rITWipxiPB674pG2VFSdUPNB7LKaV95J8O9GLl8stKQ5vMO
Kes1Mji1gDFGecx52VnmE/lREvrC5/SiXn9+b8pL8WFF0rTGeXAJhQJO/Iom4sA6
VS9IqqfoJdR/prCXOxhH2fsYHHvEP953KZ+j+WapBVDJtGmdrDsNkIgWzu57a6R2
VFwjoxb35qxwFOyUpZZMv46ebibE5gEVD6fYXz/ta1fJckd0cjoJYvDNRGGhEhVZ
zCv3S+XH6Ajtm89niVsXf5Ze24JMFPxOxg3bJr93UtbPpJ4i1EpajBzMqwgUgQZ7
g1kOVR9VUhH23+MhSbEmhb4uA890XBkpM+RSirAh20Jmoa1ec/puX4pC+/2blyUX
Be8g0iQOtZJEObFMti6nVfGsdtNGimcRGStwIdnTrWuAHyTLI+88bM37SwkJy2HE
XMAmYo+WzABrZGEST8afZrd0F0EJ10uJ6vrTWqe+Q7GLuEwEhSa4jsrsIKCAppEA
/FdZ4QVx8MqNKJ1Syi4znGB8DkUy7Po8K1Lm6kotKs1n6NQPB/dpH8HAyC5pqwdi
GYUbtuaDJBSieRC0VJDqsDuDsBwsJAxzAfHOyAFJHLs3HYN8wELqqrmtdyaMzP70
WdINWy6BTxQfMEpjxnIDF9z6eHa/stNcT8GTHUnNpkEJAzDQ6HnVuS5B9ysFxXLy
WKqS9U+Dw+mVhd6MBVi05GyoP98CvuNI1ZEh1zHVq/gv84uLp1QrQcnxgZm0fw1t
iuecRx8EXabW7Ut6GvlNWZP5aHL/sB5Z3uR83dkdP+eLzWpCK1JzEMxKI773vjST
Me3NCLnqNCsUGZ9DWZYjocaB2KjLt2ERif+4aZ8cRA85FNQ19zjzT+wzqGJCtfWk
Lbws7HvGZDZJWnjD1hD3SBOo1GEijyhQO9IWNrwKPqyl5U9jCpm2ExfPUsloB2Km
+PAkG0nBjDzFTMiF+4KzsLLwDbEtTVeWkr59tVe8nRXwHHV9LI6GG2gOYW3TszYu
ooipHUc2qdZA3+BAIWlGh5jViMoDSaqrbVpcSncV5PMJmHiT34D7hCwvBSNKYUYp
k7ooyr2LDCtFgr/e/AGVa4b92Vpzv4fJfst7w/t5v4X+ylEvdFGNtEFV1TaP6izn
i4CEVbGP4cMPHJsPI4Olqi6WX1CbxHK0FAEXPHRtmiIylrPKOFGAhS2xyR8Y6qcR
PgQqXVllLyE/OKSXNgHsHavU3ktfqwlgYCEcpXwwzP06kCpDFmdu+LRZNPIX8lIB
A2zCPbdsdCDovQny//wEYkh0b7n0Gbpk9NxXvMXBrBAv5cEl4LrX4tC4C+M1LNIr
hZccPIgwrRRj2dRmM2f0VMrpoldEjPZ/o5hC4fTX8CcK1KfN6SSrigupssaTi12k
ykJV76eeY+/aN+JZBzFYjqFOXHRibdrRhpVHks/k1FaAGaLwguAKvzPeMSLVQu4q
5JRYsE9SUB87dtD2M61ja+CWkO2lc3ypRTbbbNN2rxHA80pN0reXCwrMAVVh4tK2
0yTNFcA1jHpNdmLrqTbOb1E5rVXWpQ/H48XJt7mb2K7CPbcqB2GaOPdf2c2KYfBF
uJgkczTO0DjEKAjeTuZF+k70psNp/Wo0sWV7MWWu1R1Ythgw06ZPTIBucFjgodpM
D8q3WAbB8byHSpZXa6u+PK9k1YumFkFwFtIJ4tmVbEeEaK6EujtcSOuG1z4LSf0D
/c2p2js1prHBXGtGgJ6oUMWlxladz+DYd/SACtPrzcreO+TVjNF+msJKCfav18Fo
dJ+AgGfVadurUyd8XiIT/80FH+rtxRmQ1mEPlB2ZhFXgS6a8ANrJwIBQFkrqxvR5
hCOtvbeey/3CbOCw0FqcsXkPFODrt9fhcNDiOFx0nj0LEdpOKwTg74j2F2WYC3pZ
2wBx3Om9ICLuihTZrPHhpvIQKGXDeQ/GHJyO1LsTZ72QArz++8EzgYdC44dKk0zv
HtXQaAlXwV/S8PmamJW08sg39NcU/58hwbITi58uyf4wN33sEBUSTQRaciVaOsUJ
24XOognS4ShT1gceTMlfbvkTfzaX6cwemu2q1hAWwjT7ZPN3ECA+VTxm23AEJuWT
zD1ZV2VtJFtyM5F/oF9FnSAbqFet/0koJoCVZULAzXP1meaGw3hNIX7RBy8yjbqZ
7/wu2S+1gmTmQ4VXKkgdRj2BF2KfpzPKZV/s3m/5l1E65FedJalbxyndTeNBBTa+
G1GEK4BbuegSyyIhhQAWhM2e/2UyBG8CKYBgOh+Aoo45Z10TeoeFdBGhq5PLOzqf
5b78LC9f3by23pfhMy9sRaxg77g5p0aBdRSGfQjzrATFymKwrIaHw4mSKM8MgD8K
UjM6sR/sCCNjVZR4NOrUpEr+GxKCq+DrdANb4YBynZ1FkHM3Jh0o85FU6YBOhFac
DMNT0Nag4fvyEesapZ9h3Cyehu9IjqrqCmyNDvQbDx2GZ2DXI9FN5yvQ2E2zZXlL
7VMsAP1tu1t9Pb52l2drS4eTiOBj6V183rqU/kaN7QpYo/6gSpic6MzTnEdg51Mr
e1APbdw4/VSe9xRoWAn9Px/4EZ/ZLe/DAElJDCM0ILdCl+aUTsGUWU4lCzJ4Sx2Y
FRcjCo54DE9u1kgcqQtRND1rsssk0OiFLcWqV+iKbe7VCwlci9ziDpcD/u/ePCN3
0w5Yw+bITvhuV2sP3BKmAo6nqphuQVwbeFtIMWfJIKa1sdPE4R5aTHphrz3O9bDk
Pwxqy96giLPiNji9l1+NoiZBsIl0miYUMH7q9R6NNrzgFSlQ5iA2GedwDxPVYbts
+DKsW3jSA8F9CoD2AEeDeZToS29+NRYhL8AGOQ612ZidV1gzu66WE9sg9j6ctwIo
yetNCQOExU/LpayMn9Y7/GSdD2VSalujSFLpBcxCq9cordcx98LjhMuscZOO3p6T
2hFAl8vnOv1fGzelDpSDUtpw23kn6TMPL7xh3XoGdUFEgt3+GDeAXXHF0f0WoF8n
m8mPrLZmX4ZixAcm/LL30C7kEqGVQvgMo0L8Bib/kiOMPepdVDOtyNCzACHbE5yi
kGIAdSSVhWAvbGSC0VpBDDVVYoANvQqu6TflkYfEiYFUa5AcX0HJ5DuwFn+MpYFf
d2hesR+udCDtfAmK6Co9vbzkS68B9ukSTVdHnUMjiQFXwvKus/zI/klSO1LnRgL+
JmOFsmwYLOnS3oQBzx9kzwdx7dR1MJV5YQHAcO6UZDtTDYejfTkUtmux7N11j4mM
jsQWFB+ope6BQB6NriU2Rkb9DDTYZrCSHymNJY1Sf6bOJks6f9QIvsASEypWb/yN
UsKaLqC6NGo4x4B033uGUQfOrscirfjBsci4QCWZxSfM8T/+W5pUi/jJOlEmiueU
d/hKmbay1Ef+1hiE9v8S3t+xh7iFUOLGkJZTZMzKVINez7xwiotIl0jAzT29KJ3T
U07FkHUZBkbFh3lXj9scr8dDMXHaPCoubdKRnUquLQzHLeW1fvuJoK1n5VJTuVBz
pC74VjRCe9I/1Pp7yT94EYlIDl9IrX+k4+jyrmN0RoAuOS8p73NDQF+Jkj0zCXXi
RH4SF8CTGG13T40TfXgtPZZWiAOI3q/Av14JjfPNdXOimKcGGwWQlUe0ccsaAJDy
2vzLkChcVJSDVGkeIjNtecErOnMx25Odkl1i3dPR14e1Be8y2CLP8t7AesnI3zW9
CJ26IFnXzMlw5aAa2LDqkCjOaW2JbhKYjnPYmioz2hJJ7q1QJsh7oU0fRI/PAeAi
ZXfFL7M7YT+VUrH7ZhYVW3uhNvtSgZhFEhNazq9Hjc7Mx6R1uJx6ouL4BFdZsa0L
ospNb+K+gbBBrXziCIKnHqtecT3O9DPcKpcWPcNtAsfrxT20gaMiURyZb+6k9E3k
toUDEjBczntR/zYtT9lFttC65DyAy8blXITSg328rlm8DNzuwI3P7qJQTHKEZMB/
DvzFEZVx7M3lz54nyATdRNvcKwFF22LR5cXFI6jLInz1bLbn4l+430De2jmM4yF+
erDGsYWE+zAZDFQ5sxyGz9wAP5fK22yfXBEFTWqGSxrwnN4IawUTNy9C7eVLPvgX
SJajxYVoFz+kVjF2o2eEjezdIZ6q+Mv85EfSWh8Px8lwCylSBoWn8i+aSkpkkBKf
xwzlDyULarLZf1wg5w2h9CUKgRNRbwrU8TJkRwjxO9fUh71ZlKBUPrqse8ZKHoJS
g0o27uOqcSjhmQ5veNyiy/k11xb7mMPFHJsqcxZfmf5BZiD4NFHbLwS1SwI/WUK0
OhzDSj5bdi9sjx7aTCV7oQjxPiFHt8Ghvbxg34bh3Zb0wgT7VJfzblUXGqhue73c
X7yVrwkbiYU99toYOSFr9TB+xZS1gIkCApA7wDdYYvtX9MO3yT8hnnb1hT2mAMIW
pERtHYWbXTnlIfignaCp4n53sZzuEwRa1OpYypc8BrxwrD2wZDATrm0mkuwPGMMD
uug4gkoZhEAoqYLQo7PX9eT4nIJMd6B5C7rJPzbrBaZAMhnOvmNIeFwy9FqgSrRn
8WTP1vB9jnoPs8PUeAOR8qxXLgrmCH2fzOL5rvLYlqIZirOMY5vfaSoP56cko2RO
LZyz/ziBpSRjSEHt7dCJmqkKLsSV9L80YZmhYWairOD4BxxYseuPtYCqZfaJnXDj
ilZt1BFThnONuHAmtyLpDIqZdiii6cCjTAXh4Z+jKhEkvGrjRK4aCM2ibmJt390l
KZG1rryaaj3be5rQ4TA9j3E3tSfOmsijDV2u1zYqNeIYQFqBpDaF5UFsxi5ddKC0
0fw6rmTquF8VUsuyqIVF2mzC+YN6TZUeM9yrVY6hq1royP/aFH22EtRhW4aX/1BB
Rswcm9sWycvE0TnO++BV+qiPwnAA6kMiOYZhmwsHd5M9pppdYKGVRMWEDYkWgMis
A1NIc56cngwPLlPE5u3IPdXCwoWMfTn6acjZGlWjIIzLKlpW43qPlEwVYrC2+rHk
k9XPf5Y+9a1nPgLu8usielkM/cWkeMuuJp5e/FZpQSdvsZ4iTA4OLS1F65uEOhHS
U7qMUoo2bH07riE16deNgatuvrlsU5aVOyvVD1cpkd7VIc2ljUjvYnbABcSt12lR
6HmgH/PcYaDj9UFMKCoahZg39XjpwkTt1dNBEck92U9qsHtCY0o4CN/jJHZrIaOF
hgm0klJbpJvpLWotItjqzQ6vjzM5GDRHiJp2dNjW4FMu6ogT7LO3ohEu7Zczx1WS
vuTB8k1SdmvQgli9RybZE+tp86ioGY1uXsgzk1/9eOEQn2I1b6U3AU6WXfQlqcll
hmqVXk6aG8dd7m8mqOrDamGQfTUCfdR20qeim4xTlqMCEC/YA1Ny+62EnOLEFnsw
Nrzn32HjV1ifdj2Vhn5xsC1JBxxqLCOEl+duZcuEAeGh0U6RDHX8TQx4HT8ZS5oB
WUx66/wHRnhyU68nReb/LD70sWhpN4RtlOJRwmnpV4HbfYbYps4BT4Y8ai1igVn2
mwvtvNmfgJSpoXsNm4j6jtwqVzLEDhppfGIkjOG8gqeDbTspH7FwtYHHY6hgS3kA
WFC0N720QiytUmGkGZBqpx/rYAVCkH7gTdh1f2sbwTIB4h8OLigzt+9SyGI9kUBX
l/2hSGgLxhm4wEoqsVye53/6Iey0I3D30Agt+At7bo7mLoUweIdyJnDLQyqMnI8R
VIwJdjbMp7H+/H6xcTrPlypsNjFQ2JIg1qFgcwrbQ0cLZGxtZW++VZJ0sGUU9nn7
6LkffU8hBeGkZG5MRYC9WYsMC/DHyMMbV7RWvMkLcAMbJIqruUYRgzCIxcgn0bhQ
cQeJ0naPpptvNVz36R42X0Pzeej+kcnhYXdBWMNbOcirwd0UbftwOBsuql/vmzdb
h0IfRMdG5iU0ISDIQtQZqrE360GAxD7ppd7ton4yyTo87fFE+/U1TAF/v/IytVJu
igMDmcYFzrKAFZTsFHagLNvIUp49JVOvJxT9Lq+pTZ3IuESq0CqiDbiTn7r+eiu2
p2pqMQ3UJ1/q15rQxOQF1eGour1foifgypOI5ZjNxbPO9I7BC+AMcLtSQuvO5Rzb
H7lLaOcFPXHSmETj9VNAC2z19de3SKZQX3nLW02KM3QNuVoIapgQL0v6eSTrXgAZ
W2WfL52zG4rfQ9A1ZIebIUkVrB2JSXm1VxPCYxlFlp9OhHZR2nt+mI0M85+qFGku
LJIa6AhWnvNJoOApoQeR98jsvh5wupFm0F2OMmb6LK5JcUYLSMvBl6pFWd7z4gco
4tENHvqw8U9riOquR8GyN56qF+HWKPOByo4J0b45RV2ZB6tFRwfWViQjTEbztqcZ
Ku6Nuf+yuVhSyBY/Kez5kF+hiPzlROi+7BJf3HC1OUM8Au2XwZNdv9mCUz9krStU
UPyyjIUaaF9EOomIebCkKT8svF3Dw30tcyhmIDtCfSdq/ZqARXHDsjOcraW977Cz
K2whPjYibV6Rt8zqw28c9rSqBkOXjZZ8cmxqCAygl5482t6ZNIPuOuHYLnK3WU7V
X/kA4jguclVOe7KUz9oJGVsrRU2zoDij/h4kX0wk0bMZ+0RV1oyMrLFiqzrAO9pC
R/UQzm92HWyfKE0iud3skKEx7WYtwD40jv3lmFrcP66huo3fu4zElQ2ogTVYubER
SkTZbxYCzC2iOQTDFEObB2Jsz2W1VRkndQfjSUgm1lScgj0oDeavsErmLNlzyVQV
QqZPbUVYj3FWDinIrDU5z++4UzvNMXX98ZYrdeamuvvBvYdz0nwwuZsAjoO1SIMO
d7x4LDRgp0VyEFhUaoe1Rfs2W0R8kgnI0txhpyvz5BCMDnm1bkQfdJK3oOApceCN
UzytF+RkTt9KJhIq2UHd0+uGMEMq2AHkeaGT6X79cB6VvMjex0eFQ0y8A50vdpus
hUrm9EsT0qaFeE8kxF9smqPV6vacic5pNKssx37QLdseRGTseOS6ttWqnRR6/NLN
fgJBAZC4qdld+D2/WTN15lilu/7vOqAeE8ZW8wdzg1xvOxh4wj0zHdcm64K0JoZ0
C9ECbafaRUq5zsmfpoA2h5AaPnemYuxH02veLbOdjzT4WdEp1ooHgnQWSzLQba3I
S/CdVH3AFi9BVKr13qxb30hC4RkHH1zTf+rPAuOkxk8nhEcov5ZxdYogHdzI4JWq
B3NNBoqlfHojUotOGfYntvvO3cq37sQRvSSQ2vOtc2q/an9BZKQgXVKzYiQ32NUf
4A8KDT66ZrH+gyiF8jzlpgybGppGzk94UWQ+rHjonW8z3eCp+IchibuDPJjZIiNK
iXn5kUA9YR0w9nYDwfVDWwlhEaqfWWkIGSacREF80lILB7fJUbO9b3A+AH8JEamy
pGvbdE3EVGun6i5gbUJcWcWkDwqB6DfsZPLpVgU6T47mrHPvTvQITFOR6tLT8Nbx
LMClZu9uQFN8rtH2CHK1tTVsVjfUqSganhN7CPXUmfeay70pCIuR3ixoC6CLl7Wv
QnQuRPvNKDPhIW/+a2Ezgt4l33W2uDy/vH4s067W+zLdqO5CuM8q/z3M3pVATboJ
i/LWB8zJQrHnGLbz6s9YcJbBUF/FXiNCVDmm9tlsWZ4Whriu4mIGUJHg7S/9PVzi
s8XV7H71iHQ6mYKbSzRAIplojD7Pf4sZNnektypbSBp5NjYlkdYa8fcWY9Vc4Ch4
92rr8XzbBONMrChyTFsFpE19UxlrX6LOP6mhE7JUvBZ7rj/1Ap1ORjqiFH+2Kqe+
9NUrnzEEyu+7WToGugmPgy7Mdrx4DW1NlC2+EQ5t9iSZRroQTxJwEKihUn7pgTbH
kGvawd3ccbOd4sbd9N9Huw1E7WWRuAVfQsdvUL7JlrLYffeMtn3ISQbZ5E4DczPc
5wNdpBP/PHLBJ6/9q/iuT0HJJB45tZvjUmn1rUnakWunFkrsjbeiAQelzRLsq6qh
z7SLbcoKgdbsxePiquw1QpqmqcyPV9DYzGt/3xghTRz1OBhPfIdDXKOibjJ5JBSi
lO7lingcTyg1bzZEopZH48GvBOs/yYMw89QGHYG2D2eMKRxqh24bpS50QNkHJtUR
2pYLi2vsVDjIy9DJiyrbs9JHxnQHtrJ96XEykZaS07DyhOBikCxQcwj6rXwKGb33
kzKUYe1yfGpuNF7Wam+2nYW1k2/4QixwIeqYEoOQ79ZwFtx1wXPJ0CV5y1HfLfAX
r8m1+BeQ0JQbaauQsWsxac1bdxiwOMyvBg/DIWGc1H6XNZL6lH5zFDH2APwZp8tw
c9jJoCYEhhyrPG8pVf8dd16nJmqqdanIe4wj6jMzQ69VQZZ0v5r1bVHgcrcg/dXp
+PmfdFWm7DVJNWTze9Rae1y2UOZNPzhzeR5QGTshN8eHB14MMd8PdSxg7BoFn+JL
KwsllhMxM+luWxK1e+X1VZ7nZFlSj9iwHYjiyhtfNGnedKshE8HjsUOlxhLpWmau
NOtcTEzqCArEN+tuXTUFTXTsNnJM5oYMUBYK8u3PGsP513mw6zt5D81lpFgg7fkz
C3LtVHNERyuhuKNs6iNuiYl0F7NZeCsBPf9wHC8hZ4sExb+H+E6hxKJzPeFXCH6X
luJJinYVqssddz3sEag5iKrQD5KoiJtY2NJ/WuEHuJJ5SKMisCUdPXNi9yPwnwgv
UR2vw0CeZXJ5HDDowX6oH+NrEkpzYK4c+0AOJRpa4xGPeRF2t9Mhl3bM3jxRV9p9
keg1vfphjyMLZILqBm7fJEqGkGCSOm7JfvYzsnDq/cYd9X1nmEzh6VsaPDJXtB/S
swVk5kPTaOSGlK1otjNV08w2GQjzqyG2NP9hclP15iHyiLnJLSaHkP+mzKRbInip
zSzSSra10DcEaanf4AalRVuNrXKWzquhzo5m4xwUJBmBrYYvAIJii9dHnHclgILc
PlGwZcgOSPqhsADxZm7PQFf3WwD7wLlgaF9NP5F3kRLabIMramWJbzuwFFbD4vUq
gK+0fHO3JJZeW+lPleZiVN8HHJL1RIn+Opo7fZGYDX1MpA75tV64URvVPcwjoGIa
+lwo6G/VhIq6sYEz6z7Q/YvNiJcGjwvVPLY+AitetdPwRTR4NM3Bqw5LbSWdvGdW
5jh2vs/p9SOL+TjAihEC7Kus3NbMmtua7loXvZEggv1i9y8tChmo3RWkNa/KIdMp
3m74C3fW1HUii7k2l6DhzK6d9F4SmjR1I1UI1R4wtaObT8vGdWQFheM6bAJ1isBJ
LasiKFdW/2LPSgzy9PzR7sK2Y6cao4e0sXcSbfX4FCScxLBgeIu1l7ANFxv8Xgj9
WMGW1kfmVvUusW8bAyT+bej7io+5rszbyctt5FhDha6wVsrVi/iXuuFxqVuwPGJG
noaOzAseEm30QB4771h59/r5W6+EWxkRapcKPffZOR2N8IkoJ9iUOUuhUHOeUq+2
rWXI6XC4xqoAH+BSnkQo1qIMkEm6rzNe+8S5vuK0FwaqQrGBxSW2T9ajPkoJ4jcd
JCMrN1Q8vDLsblXg0B7xBpfP/aVpTUeL8sspOZUE0IK9GCzRDx0g0x/24gzjlpl4
fJ30R0oMHuG/o0YvwReY7TyF12CBjv3qB18559cfHJMMhoGVAeE9He5v20bupqIi
K3rwttRHXjMYsoaK1sm4y06yHhynfjtIwYmQfqIsjVN6r0E49My/2Gk2qG7S4ycR
XOW3YpIKDecvZkUk/2xp417P4dWAhVE1SPAVyK0F/t9RfNkVrKoTcI52U8obeYr9
yqC5CYzTzkXj6yasH1WFwgSTilUjurMiYGmaBcWITC9WGECk+K9bamLt+jkkc9Qk
sEpFHJb3dZwjo3lEKv2tgSGtqckKCf6V1bjnKAwbqv2C0iRERhiXMmlSJZ+wDeyH
QF0QS2zWLefnK2A/52mjUiOzJCFpvzM7aJhRCE7exlmDkl/fIjSoEqDBDixcd9t+
zk6GZMr/Go8YDL0kFWgyMrfZHjHhZta1F1aWCJtp88UvpyKAsigpAItbANjsYIFW
E31xOLVT31Tvgb5DY7RcdqCU5AngxWZfLjE5eEjkjwUfuqR32jNShppqf8TQ2B7M
OqDLBUVSBMKkN83Fh3cMJeFo54jBTAynwZfAyRf70+37ue1RcZ6IynYSVNRFkou6
DdK3aRa0LoXT4UGjRcKogC4RUCWZ0Nr6qL5OTKQodJOT+2/vJrLJOxS3vf8sFv1t
XKFK/nIqtjO7sXWl7GUlpG+IvcNZx362tLM6fLyDxw2tzbqYP11fmiuUraFmiDfp
c01+Yfvc/v7WlKw2XXzW/hDDx/9Ii6UWt35gAb72S4MTqdAVuPHvAj/iQiy80i7J
sGuIrzeusVMpELOr1zybbgfkw9WKt2im8X6FwVK/8jhBv8uxrrbh5zQe/dw0BX3Y
HfyPyHvq0v3qkRphvDhleQ5g3ZjUfgHGp2wdNQJr39UG18yLlptIzRbnBDdiyj10
5P44GtQd2hOe2gOEulXHsK7P8gYKappl7uxrXFq2Mfhw1+3TDODkw9qAyxk6vB3W
ahxcEGNZD0xqFyfiBEwEemBND6fkPeWSnElAsb9wz1fGGY6gjBdrqK95aJ5bJdFm
ZqpuKdG1gdvGkUYPDjafkYSJwEat1QdLbeDRO2PBng13WYZazYm/O2mg0jHeqsjC
jI+p3gGAK3rmFRL7gmQUD/urmZKhm2ShcTIhROaTFW5/RJtBtwObdD6360mYaw7s
UM0hlZ+P6R9ynlhbWoHfK7cFp+BDidm/iq0oUBmI8KkLWB2SJMRtQ1ZuSDXDMEAk
e/TE9hMDd2j6l+/aPP9T5tDMYsGlShooMPyOKI59xd4oNpcGwXKWGiizhscyz6CB
30CcRPSFu7QsYgq19l8l+iO1KEFGLTA7Nn8ePlh7+vDDm4878xZmA3xYZCRsSmUA
n89Resq6/OmHuoQdsGDCmFjAUna2WCv29RQiakydmwmtvO8z4sB3gkrBntSKBpJW
Y+e4QB/dj9NNRCOIT643FetyMv+cPr56Bt5A/vnPQPj/thLG0ZdhOd79tnY2eQ4I
6l+ADSRtESNGoHsHQDe+TO6ftpnmcIQpzMGt/TZkPVGOPvi01tqzpsikwjkKbVjr
lWUdvNaIiyYfBywWmYf7Ht2CeHA91tWJIeCNRFdsIizvsXSEbuC4P5Iwta4tyr/z
mYguS2u46ON7Ufwp/Q2YgK1xIyR6PO5lRyAsgHwFgl8H5IKPIidzPqv1vFN0NFOi
FAQSrd88rULnsmNFWbDhDHcu55vB3zUDeaDYrbEJ38oOe2mMPilo5c4vb+Au+KgY
VP6ObIx/xDfTJxC2St9PsEgF3p9S5fkeIx5am3vdEQkmmhm76gaAB72GxD3C3DZ6
EufOS199ZAcK6xMh38qRy8xsmlmMXfNHQ3AE30CFM5PlU43o3gQHewEZMA1rMStG
vRPO2rBTNKhCEWiBNJ63A/hayE3LkrKY1PvAUcRowYIvWmNgooq5LeJjK2noIUuq
yvSODZOqfnAeRohv4MP6XbHMPRqrhwLecMevDhm9nCZhwyD+WVuIqQkO4SyBtcLg
7f2XQUQjRmrSk4XpPgpN2ABLLlvS9cpb5bznEn5yXrSzblpriuqverALXq4v44C2
7MJAxDm71nbhiZ3YKYkKtp1ns/OviSd4bMMJTtXRhRylw3uVgMEqxwaY/4FNlGLs
m2FvuXpd1zhrOFMjxsbpOUJKhnm98sOrfmBCifTPUEcqT0YFyOl5oq2SgNZ9/VtE
jbohaQdvq426vr1OnJmgRZr0lawhYVa6OtjFoFmJcMpyquilgoqm8MgL00QQrl1F
HHikKoWkcJXUgUK1e0Ud4r1lQioZNiefBWjbtZdpqg7RUL95NpgM/snZi7rAeZQL
OLz6jRFeI5d/x5Dvekl7qOdyiIUAmR/tGf3HIcok9J9fTJCOT7mPyuGGe/A79c7V
eQXZY+TjzKD1bHxToW7zeoDylPBiGtL3vU8uC0HAi5Nti4Ra9+9HpPK3cMBDpgbv
Sw9gQyy7O82iXM8Hjv6vuwsV/+tSo0eNwKhfrMzYErrkjgz8GI02ajebUJ3Etv2y
9bBMxhNJQMqf0NIlbwZw4Oji1Maz3NTFrqOaq4+hbq6VNTBz6DhTsGiLzf5PnyXK
Ps/QaV3m9PGQ5E81txSM6qnxEhhtHrjY0NQQOI4JWdRs4R2i6I4whtDJYwPfyhPz
YrY20++015vV1Kv2UnXtbrbExV+aXMeUMTJEoEVhkwwj0nJafB5PWuhrAJZslZJQ
CC9sjSjYB0wDnGzg1jZSHocS/xAYm3v70Z5jR9GB+D2bBc9koN+9dyI+wEZAAhEF
zw5Z59VBqNrmGSf4lIl+sdEmFrF5dnKDcHZYScJeSXfAdntTlkf2uVFg0Ihg5wUT
nSnpJpt/ADgpy+wAASaKoXFdK/QDIetnDqMtJoUbEyBBV2APxa+S+IuLrgEcs56/
qtMrsBBz4HLP7x15W28qIlhvVSNbrVeX68VtZOWjbexlKYMwgQjsFFiTUr9VPVFn
ztZVVYRw/lVU0xeoIvPRYV+Qoxme7UAlAXXsT42dEQ3uKxYXpEbD/eOhJLwFAw/f
+lLs+FcHP6voC3JjlzXHkaY9j5HaRTa+R1xxNpaTZ6BlcUKX28eybiRyE8LG5NVS
NCsv+wQiRElZJC71KpgKrfFAeyevmuXhCbfjCsjlJGxRXmGkxSwqJobuUu92zey7
qm5BCLL5DYOb9fw1c6UBhRXTvcuGvlKGmgzMvDXoG29QE2JODes3G4J+6Ium5Kwi
r3bPha4IKLqKo9vGKUdR0BwusybZDXCVf6Cz6dmdAgplv1nrRMmSJA+JnkAv3ZAo
H1lZDGtjM48RTQbmlmg3OuLYInzJnX6wDsmygnjKV+k4J7qzq/hhUcJx5Ks/IaJM
PGtWQtC0jPofnng5KDeBae7tkqq2J/m4jj51UUhFhUluhjobI5JIosn6OqZh10j+
zIIXb+Qg0ezDgHrmrnVIu7SQ6AVUf4gZorukd+qtEn728KOoJB4lIL4IQg2/MMTW
/b0brnjkgYwETU7K8YlgIYvdzJ7cC6z9KGgNBilW0ma2LiUPQ/QUqlGHKNf+2vzb
YTrcJDn3SrOjkDAhd00T1dCLG3cJC2aYMXBgNCnKeB5r0Qpwe0loP0Ui1bj/8BId
QLgjJWu2zvgmzJgkDk+ekNZs1pfWbn8mUJfYnF5d9LnrdZKuLYGtizHStfOTLqn+
GxHgmZpxETxc/WnrppnPd4Lof79qbqE4kDfsxi10GFJsPoMHxECrNBiMyzTiC6NM
IkAZcKyJVslKcnMHwTYUT+0/LG0c4xkNzI6gOiSKJ0+rnr9ndAAN/ndRPICJ10gd
87xAv8idslJc6B55gzmQLwd53wUOkWQ5D67b5Pe49K/ExE7ayWp3mwC3Bbm0u3Cv
7dTmZ/3z1pZ3Fb6X9ebILqY3rFTwiUzzLc/ISzYBISmF0PGlswIYAENbMu53i3Ow
aell49FRBKFkFUCDZ+D4rncri/Hfn1N484LbUYDvOtyH6xkbP9hQP2sS6rlM9L4Q
r/bMTVC1Py+/vbMsjDXoUlieFN1EmiresF4HVJSxzxmn7/yx9LYbY9RNjj2I7+Yz
uDsKpIfuDiYyTJf7gwVGd4Tc8u5QUiUEl+qI2MN9Vo8Em0FryuTdDrRKNoo3lFgF
CGGMX3f43L2AEs2Cik2of3V0L5h4RqxR93fNV6zl+PMAyebhdSWUCW/FhZtU96BR
XihrfAuGzd4WFLSZbVsiz8iQm8BrmhVyVuvmUdCaPIT8OGDM7Mc0WEHTD8snndI7
Wny28GahSSrFMoilpstF4tiY5hQxqN+/zSKtfMVExpRA1uH6fVbrimsQro30XG8s
fGklITIRRBsGj4vJsVlHaOLH+B1vewlVY3KrRmD4VqXjWtXTvguZPN9CW6d5I96X
rJ0WoL1FeDvD7y1yZ84W2DgfjsiklaO+jmxKqPRbCKjdoFsDwujrx0S1zpvhevFB
uDLl3NjVSRwhRq2OzGstPyjS5KTmJOwZPMMq3jZ7iDykamc6JK3QNKhuBd3R5sNK
2l/9Gr1jiiXMFUUtaF643bL4s32mGnvYKxI4wErswtAMYev2lThmDBFxjDdUU1H8
+7jnFZQ/BucGrot4Rf7G8S0y5gUpuIhPlxzJ6zwIPvfm6YEqcmgijrEKxCcmZacW
owiBiVWGvMk+KJZiCwOv7eYNMtAGC8Pho77CdJjfZzO8+eq+bysB7W0Zpq/KMhWU
fIvjXK6TFMKxw/Tr8qodnAKYTTYWduozZ9fE8eAd5DFQkX0O4JeCbS4dFLMbiCQy
r6V9TPxPkMth1yC3dI3i8XnQsXFAt/3ClVuutcUd38ahyVb5kzxMugIt1X2bJBw4
rNDFna4ZAoasphbm7FFNoPUNnoELKYOfBc/Rl/Av0dlf+5xywwI00sr4maAcxyYO
RxDfLAgAkZhu/RAw6vS6+MYuQWZS1DhW14BLQ4diYfLpRbP3OerT2VVePb+3VPeP
Tlzbq2C3fbtt4DyNIz80k4Cw0K3+Jbj4T1zk5s4pw9iB6+xx+RH2OyigpmNSP7YY
o2xsicTD1QHI8LTHLulviQED8An87gigHkReQ2BW2YWo41/YnhC1yvPoYl7oWEyG
HSd/6Vg8++7s45EKC77++qp7hr2EpHJPu7cYYMTvvhBJjYQYLOMTiwOGIxXjcWyd
8ETijklXBgnhnk2I4JPTocX52ZWDPsxE9Y9E6wpVaU38SBPCNaVuoks1h71oEW4A
ixZXeKV2tXLL/yX6jYkoka/FGibyX0GpMrXh2cO5IMTj/xHsIyiwA3EgBKtfkxGv
jgm0teWgZcZkVKyTKKqUbEeZUcZzPRfk+XYfdLvGLf57K0m90fiMksrPDyuQH8or
XflAiVqr+u3P8U+Trg1HBKOq3k7z4cwB2Sj2xxzFhy4xvsLBf/Glhqqavuof/jKp
jrxIIrldvOE5jMm30CXZLv7J+ECBJQM18i9vsDHJfgx/c7KI30NS11wiA24GYiH5
/u6TU4NGaP9kgxn6GApITUci1/RgX3Lie8eQyDLWQOcKg5HsWW4k5L+hvhdO9DOz
kpiwyzsOF8wOyAGztTEEkFj9YvNMUoj2H2vGUvHJeHJWehkUyb0BYzH66NdImkzJ
UFPgLbbGlP8Kdq6c7g+oyr1mquJPI7hfZBZlPLEfJKjIZoE9VsJZEj63ZWhom1Gj
0pEtxEwYABh0s2AY/smiq9TnIGOq/uoiyHvm6qCESYWX/kNzKslyGhlizxcQVL1c
b5CkwED3wCVUJopLRnQ5CEGJusxvtgnYHRECC0lbvmkD1lqL9hYPCepoJhqInU2Y
4WWL3Asy7EG7fonkuHi3B1icdxPkjxGL+cOb++GRaOALUlfkLE/ldfv9KcM1M7JO
aEDL4vWdHqrIx8JJ8gQe/2kFL8GdSVx51Ml1rhIiiTTGH5GSiNqqB+ggAc0waiIl
VYYUUWb8eE+W3HDvCoZ9rp+2YxuDkdn9k+kzQxdASuXylPn8wzNKDQtE3bZgiYbb
4p6V3s5JXz0WXFCm86SZG+moDnPITiruTA/rLYNKWRtybM6v61rDnokhLFBGzgQJ
Ybr8J4sF3Qns8E+UrY2S190LVj3yFj7IJFDhEPiBSvVmQME65OJocslvViC6B1dM
/Q9UFQbOhUzpecjzEyaTpvoNL9rjkXokzVA4KPxJHWvf6fafCvhsvXOz1G1Gsbz/
dkO+FXWTKG+uCTSJL+sUQ7m6b6pAhb4d42J0aF8sWLGPZin/PoC0H6Tf4xVTRlBc
qshzlU2wfhQP1/KXKutSKwW7Z9GrLZBptPFbhxAIiuxZzFa9YGoL7pR9W0mxcpld
iXyVpti4/ph4VwlF2PBzjKQ/yr6jdiEUN27lYlxJkjxZ/cUfbYdczqXhsnzbJZAO
G5iLreWr03ICRDr+bKwLTn9HV8+ssOU+OQTuOHf888OaaaMFt/1BPC4qRsZYLvBw
AObOV/C2Y6lcDCsYki2jtFMxeEKx/dnTUHsik85oNPaRZC5SJh2QECZK8H4j2eQL
joMFl8roPP2hDfxjmmrOcOvhiCmlZvF/TCwJfb3wl0FReHMjdSDkJck8zYLzVx8l
HeRCfejtvmsxhvHKn1OXZ1wgeUwLIiu4HrTSubOeAT2uIdPVycEVHuOUW2Mw6nEF
pCWLApfpKGKw6Jia+8jV13DqQ949QRCWxurNKStOQmMITZhHQjrIo+QZjiJqRYH6
owvQWWBc3lqkCE8rHTPFZOl1m0/zdm8o3skenILoR0RLls07KW/Mer+A/Fa6oGaJ
ci9oCAwtXwdbhyMGAXaWMROPZ82WKPveq+SqeoKKm2GTYcbgdIwkqZUVI1O4LK05
ifbqjhr4hV3xkJ/Q+JYxOr+lN0NF7C1IXsl1K9yTFTVpx7SdjYgINrUFM0pTEbNP
zVePHcb/FdGeuec9ZCmETi6lNMnmZXneQ2VEq/2VdXQqiUIQ0PRNQT9Zy57oNyBd
2UwiVXqm3BB+q3szTHm+LwvYaebHSnIQfW/rIvkJiAQ1aGwtxQCLGo8TlSQE/p25
C0CdXnhoXn40z8uulwlIjCoM+6NHr52mkB/990Qw7Yq+QdDd/y0lk9X0/mSGlcgp
lNMRpr67ssdbzQFqZc5ACyF04Plug24+KaK/27A5RdLMd3MXej3C+HZO2sHPM9Wn
VXEBW6BWt65NH+Xr3FSw9YKV+8bzzcOu7+9+lW9KI1SrOWNm9Idr2UHDMGuhAZSA
IXbaY6J8vFWFCziO+oTLdlo3K3ZRxdbE1JC501u3FuBrBWbdmhfdvuJ0PXs/kN2T
9yFuDsxR4f/6IdOJjsDJoBKF9N+M7+uhFqc6cjL/d+Uy0jsZJwuwlxX+Uk/6JlCd
fFuINavSe44m7aEZSL+DLL4qAdHxJ4ZtqVN/JPmhApfd56L5JtnKpOQsYEB18IOE
hjkqASME9QOGGJFwDhm6H6s2Oa7cb+nt/DWL3CwQSl2pxJZXDrBbDgtpRGwaRxNG
Xn2KeCaS/sLW/16dkRN+DScpYa15j3Aw33AR/+yhHL7tRVHIC6+lZSXH+lRzgE5E
f3Lo9kixVofJk7+nTKKIjboz8Np/rTwqxujj4uYf+DvoptjhmbvG+ouOElq+PIgF
9K3j9IPEELi9ZClG1VmQeyQiYxUX9SFYmECTW2twQog3V6GnEy4/JhfRmmzcRGhB
zT6wlGqhF712SPz0t4nw+gB99T5JkUaj8qvo7/hTB1zPg+sD5kpF3xQT179+2aN5
Y3MbsDPS05XsMiBJ8oumLAmBPIV5MCE5SbTuP6W7ngHYDu2aw0i6wCgRCMgBwPY7
u5JH+O47qfRrWmwyEn/cTxNSL8tu6WygccGFIVw1a6J4nKTFiRm8B8QNMXgcbQru
YRwxn4GYhS0eVRxNfhh0gmHfZyMXJSiPWAJ0RsvPb4gY8ywyBP/6X4zYhwPc6jpn
//l9Upwpo97yLQk1SA0C7cDTisjo3gzvJ5tLrfA89HrxTMnG7L+qYHgM4sQcYYtW
BlX6i1GXS6l2lOEqJk5/ZCyQKKQBJyZ40Li/HaiB6W6drWsok1+Duk9Jg+4dhvFW
bXhQQQMXTU6ZoBTrLSgPnWeKvhSlcupz2VbyW9QPz3QRM9eGVyib0L4HpIZlQtuL
6zV6aOBkvzwh6NH6rzaDKwRuoZfI8vsMvHJMVTADedKcX3tkm1/WEUPBN+JNcmil
MfK6vvyj65bNcKFrm5pGzQbEnlQp9CS12edu0u1Vo3HyBm3Zia0PoaNLxZ6rTkmm
j6RmzPVM+mEmCnU/3NwmEEtbVSsb/iXSYjV0XuDb4XDgrTje/GsXVZPT1ySzH86P
IwBtU8Pa8mUNq1ZCZOqAyyTSWJJ4CNts9l8FqHGkzPDvfRAY3SNdwAxsAakTWMPz
QxkfXQaUhFMJ+uf6cbpdlqs8qKTxuAnxT0/6SZSKZ/VmCCOGKdRXaFr5sk+xHHyl
LMlQR7VYirAp/AYaaQYdcY3vNDq5SZ628uDXN2J3ZkIjMcVZDVOjubD1cvS+h7Ak
76xEBB2h4u+7P+18VNp2wwtMgStKmHrcHakd8B7NoOETT9XDziTgP7GlKQn6UVpZ
tjGH6u1fxLEseoV7YJ3lcakFajWMqRlzrOf2Adelq0NYiy4kMf0tGHVJpiKcpLdT
3UPcunWRm43npbD1Cjx/2oZg2gbLZ40eggQSMsCVgkfamDaz599DhsC4mVU74gxI
pu+2x369fqA1CBKjy+qhEQf4EPHKjcRAGSvnooAKA1LXBYyhHolzl14MqXg86+iS
3CJWfFoSt5j7UosDLOWXdxWC/BZitd7F6vHTkxiURa2+m4lDL1z9kl4tBBpfCCdK
6Qx/l5vaPgIqrWPnwwTe4dkI4sc4Q1M+J/MhsjSXUtTUPG+aJxX6h4ySG707q92M
2kaVWYxHnT7mLYsZ7R2hn631+K6SEtX0RfZ/hgf4Tvda0uT3uR7gPDzWhRlNDthM
crIulwU9ZdvyHsS6Pfmiu48idgXS4SipyLmgb0+i8e5UMPDf7HJgBzlJVmubsp3B
naTQw7nVE2+7dV4lXCL5SVmoopIZwQ2hMWS0idumYEu4z+Ku/Na2zInyr08XUwgx
Q9MW0vhPHEhi5ALAuxgAo1viw9GibomSkNwn6Ck0/Aaxwnk2qnKCj2y8FgDu9omP
lWpjK0oOORrA4hKYEiB8CTm3SDJgedlNxu9gvb3WToUdgBeJypg1JXfCSJJKMzJE
tT14sCpbWgyiGpwbRVtsF+UORfo+lNi3a8Y99JsAmG7yOS2yDU2YniAzaTejiHLC
o0kxuPONSkjTD2NO2tK/taA80IxdIL9R0cpjB1QsppJomCNoJibAvYfSiD0IFygz
KhOp9qaf2VjGixURxiL9Zf078+rDtt/kvuaGQ/9RIGs0/lLAMWzlEHT6+jztzp7m
F500+yna3PMrLKzc2H98hcAgxJwIUnJkOjWvn9S6qz6DIsXo7cAFOoE9HefzVF8f
OtVjIPBQkSX/OVaHzUb/KvxkJRnxQAM1UH+LCLTsYXsz6DpbjwH490e+2Q1AD9k9
GfmS43Zw28t0/ne5/paNmCCnf8QNn+J89DagH1UnKPNZcUnGxOeUrn5G7RsN4SVL
r6ITdRYKt1HlYowl323p5N8aAnSWodvxOSvsbWFMN80TjHg3LXfL2NqFDxiyRW/Y
k2l/b/BU9Qy5BFUa1tYjoXYKeI+1C91k+jGBb51q6BWQ+D7gGrxSHpfA+3HWPkGv
49DXAiXabSo6AifkJO920PCwYoBFVwEV8YfpvpCPIFIuBhErKcN+kGU8OgDwXx5g
RY2xPdg2YSHO/KzHN/grWWWM19d/bd10GBAxvavQRgXLCNfxrReXT2dNfCjeqTeI
Ncal/8N1RjheRONX01eMuDkzSFh8wgw/8u+Kqf5hd5wDdCNHEh2SccHEOwrmdrOs
ON7wSLoNgcB7kPAK9sIxubBg3D396nB0And9NlXywXNzaEuO5tqRclJeF+LINcHp
5YzNMf4JsoKRLkXpTdbx8eL7FVvyiZcbZlDkdscx36y9ppZStniJAXNEk4Z2BbRu
SpXxS/HtVh7b/3PcMNvpLHLpyovkAaWazrosQk5wIGfw3LnpzGCY3RBpIjZQfbuM
Ay+xYk++f5QKCB6wDKMTQL38Xs9vkSLiMglP4uvLb8q8oYshJZLpUkXUoNfMr8eB
+qmfJqjuJY07qwRmfWEFfqCGm9Y3BS/fyMBBlvs0wq+u1Ag2wahwNSJ4VZ/FOmw6
qAboDv8s8r2ASg2hiYFlEcQMJFwYtnBZ1BBpst7E/B1i1kOGxwj6lsz7Y1d0Mvf7
UQxj2KCrcBQ3dtBNNwF92YkrwL9YBP2O/9E21n+WGElE83mje7TDStHHXs/FU2aY
e1fVRgey/Q13TLGqYe1B8KcmNFLAWyWkx9fx642/ze0iNuHVYLnUGj0oWPFqH1mF
GNNo4/ykpIuGBfzHK/vFqk6Lgl6E0AIYszEqAFRgqXQBVhmAZd3aGf5Kvnn4MIah
U20IudaaHOb2bMEoe8fQs+DpOQyIlZUrxKD3gHvW4lU70RZTv/Vh4zcvVe8WN/1h
/1gQJgltbOvrny9ELfko9brPX0YKKqqBU8i/YP4H0kxkxO0YoSvIgcYaxBt0MUeh
YYejszJosKNG6BPsw83RDhfoeEOdm4i8lHEQuLHvJllrOCKakqkr6C2OkAIg3CXz
NrYtfpNeHVBWZDTbTkqE7lUZQSesc/BrAZToozuyCYyPciWFP7sDsW9m9S2I/pMX
tbgWMS/VmfMb2m+AIwrLDBQ8R7oec4k7kVaRnVeaWnpxJx73zestBLbFCxwCC/jp
LPfuJoftwvswu37+HamjlFSZuYnJ4hr6fLhzeKz+ky0KfUV+rtCETcOCLFUCBYPr
FRaJwOgDUU6Qf8xOu/Aa3IOKwdjG0SiWi1LoKGhN8QvscW4kMgKcE/uTZ0izN2oh
vtrhAN+13TDbRX9X6UYuTpmkFzuPQYc4kcIhEi0aO/efcwNMogBaU5EsCYXmteYY
znzzOiRAn0FiDEJ/dKLnzeYXmmsn+lrRM1v/e/a9KN2X2Ck8bBhHs1WlNYOSmylO
UEuxy2sNsPqMnLIvKiHTMtzOuxIrwK65FCSdA9/cLStKnjLH/x5ssBw8OuaXzsw0
cOo3CIghpfgdEvPY6M3LMfIQBZeLit78SxLp+GeaaC8ylN4FoYVdSRj6fIxgnuGW
MX2X1Es6gK1qftLAcaiLlux7TGvpegsMFOxvEu5v2Sh/Tg2Iy8ZofLyP4XdS5dN9
rR8zv/LeH1/PyYk/aSygvdmU1em84mIp+f4AZRD5Z4Y9AgtHaqGTZOC9Y9iMSadd
qasg/rZ25LajUnlJnhTrokKe8hNzAqLLGIhAx5QQkRZxll3jplb9pHjOio21N3zj
4JMHYKaftTYbwyN8Vxgc8n2fXvaMYqjBE5n0l4AMzsX298xcvMEI1Qjut3JqfRnO
SB7fPpm0oVumMHezeMLsGawYr8T8msuZ7ViOORwb9orMK4es/64eEChrNzELWGAH
17oM8ptBEByhinF+zVbYAZ00QpBoHFhM09CKsHWVa59ou3RvJqtv7hv26Q+n11W5
9MmhygU9uwPQpriH3FeOUuDXjEpKZFIoGkBQ9iVt4I5uokp2tCNeQnUKb/K/yO0l
JyEN6xncUe5NdmbLk+Fssb9fi9zkl20ulVQJApUvDmHLh0hszq/BsNmDKzqriLbm
mLhCNeBRl7o6W5nCaZgqzaJ4SNAIeR+UzPkmwJ3E4r8evAQyQIghxGZ8U6apx+fF
eNMzaiAGpkKHRHX5W2x7fQrMc4TTVTD8Et0ialfm0Tm/npmUN3ljugOX+AWC3Oum
g+QVdXPKiGCaYyAfEygQQ3POZzbzjuDtyow+TmhRePkUNApvoB3MtVTTyY+kYvx+
0NDT5MON7XHoOcQp1tZQYs8eMgOYATq7/MdxpvCMrTRqUzPy/9CWIdfbSHvTFlGu
wCWCyBvxJN0Z5R4TRQMLItsgb+1QHlKs+eYQSovnaps7mJ4J+b/6QByxLPjsSbCS
uRjyOdIbSHUkuwT4KqN5VzQUo4OE9To/vwTBzoIaYEDFpCJErQCD0K9Lo5ItNi8u
NbrlVbn4eHAhxhJrxhzZjhEWJeuT/K0O3x1xvDFFhj8vweRRR/4ngLRv6qnFB+k3
9A7qTf5hcP0suP1OA/y3Asjlq+qdXBCTwh/PHKylBeKX6ZiHBjdgezBf5nzrRZA2
DpH+XLkZ7tce0uxZt7d89C4vqWv7E9MK3M4JPsFn8rMSWZk+21pmmb3ljxK0ANVp
K/O45/GJxstTwjMVLCbM+GN6Encz7fAv+vX1PiqdlPlQ/quftehwe5cMyXT5jF2C
nxadqB/fjEpq8EQQ1aDfuEdEgQA8CEgtoUJQcDNRqlIEyu3r2kAs+ffC8/J0tcB1
V6h1c6Q7Jyy8ih255rKqgkjLPcjNL1XdUk1Cij0NGyXo3KIKlC9jJtYQ7SYvwUqZ
U1/bbBXPUpc+JXPrCGgKaM+jpiJUlKXE12bBo0PP8ZL/gqMBizRn9HF1s/5mC5QJ
WReHVeu40hKjV51xiyevLDNmz+E3jg6+8YJ3wPMuBrZtVGKDJCl9DM2loAFiWo96
O+tI7vN3wbFudkfdJXjq6DM3LJ7P9PUa2ihlDFP/Ht0MurU3ShCCuaeIWp2tK6iJ
G0baxcaVcnbXeMTRVgzO8rcYpWKLtJJnyCB1c3eeCUf5zg0WmyzemQqd4d3RHjqZ
NR9MXxcErW+1+syzrHHQbphf321QsULZ16lwUW8WiqDgfeWa0c3d6W8ExU8KbGv/
pufjeELgbqdbU1qFMYZWsuLYT0SNwmocwCnKIsxhJaP82lydx/VJwfd5xbHO2+Wm
UapbZ4nUGg3Zzvw+t0SeYWxdx1NPhObD+valRVS6NIj+IBSP2kfYXjD6DegOCNqQ
2ATPEjYq8EvT75VPUS07gI/QDMqsCpDRggZmxyOdJYagWKJgjeVPBVHiOgUV2K4U
LnTZYu6NdA7maH8dmBlJGUeMZX5Y7dDam5QpzKqe2rdx8JQIpu08udNIi9qJz95+
3KvlfOYZUQ7Y5fJzqgrvrvxxF7/QADdpcJ5GINdJyB9jAzu1Nyxvv2DG7/pKV6uF
EYkO2sgWzQ3ORTScx00cdLYJEGCxc56iiPRZbcQ+Y1iHJEfPj8ZlIk7v+IBgsFZ3
R+xadZhLQooIsoekjf2bvyNXhU3Woh4V771EXNMhFNsm3FldFYJnFwJntVh9z7Zc
2dHdsXIEc/WGwNMKffCjlop9+9szWRUxysPoj3vYeSq2+5geBEBxmR5OjFExAZBl
RtS+rO3xeHXKf7LtJ/4+X7ugI+ymQkZAb7ab77F1W+j8sLgemw7/YwoFperzgZkr
oB5jnROrWJ5U8+4fh5asXSRu7S1gq3cDxHFmAYuCtPI+jKaIetLL6KgtH40aISKW
8gh+8+TB0QEtc+QswIQa+zUyBLPQvWLvfR94Pv8k234kh8EI3BWaybF1vk2jkJO6
/2ZAR5uQwaCYL3QwDtE0i5bUi85s6Z/4acirUXOJMrl43WDkLUIlRkzbG7KQyoq7
lxglgTtpDt13kzbgzkA99oSAkw042RMmOUboN7jiG/+psPgpVKThrwn+0HcMtQON
EdsouubZ8bgmaGCprXaxKKtWLlfds6+oCvTBNpaDyFPYcPuHhw+I0XEBplFmQ2hy
m3CAU1c1s0/oTkP4bcXi536JlFUEP1zjHZxXnd1zb1xakd7K1Z+gnXHxV+ZuUbDp
JDdF1xsQRkcrd/rGEHEIVXfB/l5dFhfAOJrbB+uRXah+KvrxJ13KG/PBGah5YFA1
Jw38QTvlw68c5v+MCPf6OaDgUB/YFPaG66UzrUOPTIjofq4HhylUB9LIgNbpORoj
XfES6fnhr4xDDvHqHQ6DK0xV4F49b7ErxxOtMUvdzOBLTGn1HhXAt0fP7/leSLTL
6XcSKDrk1ORp8/4UTu0qwkbygd7BxcU2uVM4dimIwOYCre5B5GGvrjYLckATCBYb
wrOr7VvDwQmgAQqJMw4vXQOkDABGESyS0JVpfcJNSLMvRt7zMfRpEksYzK0jgsKY
cmN91BahfhedBH/yve17/DZhW1vAz1ZInjBFKsmOeNF3mxjI8vo/ChN5UxCicPW+
ALr1cYL039LB4Qi6O9K9NEp2DyznPqz8pfSmsXsS/Ri/8x8fcnzqilEIrEqFh7zk
iCoxlfyzRBCy1R4nbL2lnNHobQ3olgx5OxDmHHbSKp9aT+x5s3zKDcGZJFxslHTg
BkZ3U/UE7D1L3kmiTNjmjp4cscvr40KQ62oK7Bi52LpeBGCeW1rRM0xIS1L2AHBM
19B/j0Yor5K7f3bmcrN+uNz9WRN8Ikl7Z+LQ+lD2erwnbnFT2stWWBf2ETqJYNQD
s6x4Kbltu/aqtrCp7oSijPWObckfYz5pUDiegdejdbad7ZvuNbkD9KPs91+a8Qev
8ZiGG8k4K4xtN2urslTFzBmPBm2tTMz93brP0kCoMQyoERQ+3sw9nmTins+3zhRl
YfyhoXKZa7dRsm2ie4LMCS07s4P33GVXE4ObuzvpmOhOIiqEyaREjgStpyeSti/y
oyCJyDZbn5PsEQG988OEYlFptzYaV4q/l4dUc8vniktiSnIzOCuY4u8265BWN5i4
EDQKvfmj33K51WWyKUoV/K42y4RBjzjy8FNMj3Dcd2zHKhRj+iv8GYDqF+PTcnyf
I3xUlLyjDTYewjbJZkgh1V/+YCUYcpNn9n6+IjmkidPoCz+8HMNPSdkjP3ssbgeE
ni/Ilke2Mtvsme2gb6iQswi1q7yPX6k9skL4L6nGBFir2AJGmIplKITcloovB/8c
1xop4+S2hQll7KBbs+1+MMSk1LMCE12SZCwtaid2lqIRcrRJpFrvETYjP/WRPDrz
RbBIt5SHPMfsJrqtP0ou/Lf2fUKEEoyrjSG37xVOC0k5PwZEuGd5+jIWfTxyqEH7
8FmilZ4Hqpzkm/75MJXkmGFuXsLGWLr3hRLMu6IO07dxWvCIeMAp9mDpJ4fSAQmu
lQwC9dSSrygUNhHMQUKcHTU/adXNLzqzFb16htxmwBKuFZSVEUqdII1D3wsPxckl
Iv1fbblZDclULjbkntBB796Qd06PZ9JdtAvmKaiHNiLfaAii4KC0P6KXNInbUF5g
gnpTZzDdzcQyPbWzpjdVO6n4vyDAZjmzmJznIMmOIFaEsePdvLsDtjkGC/R6lRXk
mitbt7z2cuFgPIa80H+i/tvsnQVYtu/3L4pN8qlc6I3a/ejS8cIIChvdSgNS0s+Y
+hOcoqmkgGEjECDKyWrCTp+BFRiR94yl1oZjG9zx1WZ+uumOmQKrXJgDt8/qZFtB
i9ovIdPb3AFxtFpPv5ORwMxHNFNQckmAewGcmsd+/Ixx3tw8/baXptqY/p5zEsZq
EBZVEIaWJGlFtZmrek8o4SzFXo2LywcZ3n4g47e2MxNix6cdeXQ/++aNkiCWzUHJ
lOm5Uv+TB+RbdycKyPonxjwt3gixHJHDxVh56Ei+jQs+ucSGJR4NlelUugMXhPIe
wFtYpvlojkz2MA9SUjAEV46L25nO5BfIlBmekpg2nJ238451LWjoaA5nnTJkN7xl
0jzAuJdZNPNYKbo2DfTbuqwKROQaeysjgf1G7EFm4a4q30V/miqcM47jIQ3CD2Sm
NoC+4X2Luze2oyeYmv5qhyGEdmTPYhs2lDYti+kY4icIRRj2osh4/nSgYpEQfry5
qD7X9j8OQb3tQyIRZcbB3EzKdw2K2z/1c2cWmWV6Od8lt4XYArOzeE7yfiAZfd+Q
IrrSaHHyYlZjyQz9jC/3cD/et0DW4jkq6AIseP6FYktknopfix8/a7/FIe9ShpmN
+sqTQrwfrf/ArCcWlvXraGEFq/Al+NCQ1dnLRxMS4riC3CCZIfkL70rPpR+mXY1j
d/k7AT3KhIOmEfVC1ry05Wp/pjXZe+4zm6LK2vidhPjSpZz77FQhsObNCanWwXXm
618GVxUQRPAPoe3h6BC8tcJsvjtSWMxY6V633MOwOQ50tjgcFI80gwAr6+zAu2yV
xULS+xKC9pQeA/Fo3Q8hpuI0//8jd+VWWNkeSj8dHK7G5RXMZRNZ6JkfRn3ulI1X
DOZ+HoD1c/8TSG0sxN5M3k4mTh5FpRga7zKPXhR+++P7AwiEBhpsoHEmF1y7wBxX
AvNKUyx7zdtL1Ssf1o9383DK9M/w1a9dIwH1gFD5FX0JLhoLFe27hODbFHDlrclp
kPTz2oyAb9osp/EJ4JwdEcaPwJTAJWdiXIP6QN/9JdXfhpD3SKONkYk+EsR6Cm9h
0Hf7UH6MS3u3tfKVPsHirK7/aD+AVKF2kGNtbMjqROQRNn/5FqpJDL0nBWu/sCIn
5knsJsdtfQ7ANJePUrmMg1VvsYMKpV1zrpOik78Rfgy7xqAMMPU1guG3riC4pPt4
ieYqS/LuhQEe0eF7s5wxkuBaOW91xXdnEASI9wbS67THb7MLADWS7/SXyfm6LWaA
hXMI9CoK3QZAj9dXdtgQOqI+ZhT0rR54RDHafjzGDggkP4c56ILGbQoslVKrsRhE
QHivb3TSGTUBkRTqlbac0awdKw96Gi7gg+6i3ppFbGUFq19SmgBY5w968Kj7siS5
TvFyEX8giuddo6vQmmJqjBa9CNilAbn9xa3qIfeRyVU18kePlnD98RAR/mra0Oqp
i7dsqVw+FxR17jphuMcuIgf4jDFJG3dyeCMNtCdYQ2hht+OjNhbCwr3jCm+20VPy
3bZA6eR1lCGxGyZ/D1ylqMOP9JG8kCYxdhHSMNilmKmNMNL9rACVMzjF7+xtScSH
JYs4IrejHzw1eO2AWrknlEcHB4rhiSeNd7C2F67a+UoJfqXYhTtsNU9WAJPgCyOx
dgejLhrxWisGEYm6dJdodptc1WHhecRUHv97m7YbUL+knnzbQxgRCfUm6/opMSpC
IOBFCVn9/51v8Px8yU+aznjrAZQxqnoDj3DcyFagX8wzbNHe0FGcrCZOmVaz+Hfb
ZKNm2UWL/pQjDlY4OYpipK9Bwh1RVpXWdpEh3EvXpcHHb6Nhtc/vj8lVjN8gAT8H
mjyLf9IR4RDqRhm/T1zb2AzwyMSLR0QjgJ5NzAairmSw86d7k+VnRwRb3fVifiDi
LTlqSejfA2eNCO+CVjho4EQ0aHz5+YTH0MxovsrN6D3aiO9/b1i8RXJDZLvY6Ooj
QZjBOaVs/OzBB+RCumn+5y1WFA5A9qD3lGq6QGq93hLsCB+lWlrSDOsilce0VdWG
UJulSA+QzUNyzLwEp4HWwoBum4EHMYYAHe3aHB9bcUQM8f2XlZSCgfrzZ33wKix7
FLPMFB90KhSQJk/fuEeT0ELyHukXrCEtAgExRSxtBG2H/T+5YkZjiZo1mGEvGYsO
mkuooOKzFLsNAwQH5Erz2frqXQLAqGZu8+6UCMEN4G3Bv7GYAkjBoLcT2D2GER5W
Dy3jOVT9M/3mJTYWmQQMgVtr1mCtGoFtDcqo9NWcIIDjt2CsAguNn0RIpSLw6iGt
wcIwv2uJgVIC9oM26KKxBJv5mq9GWzD5H0mfHk0VVRUoPLm7hIBXFKVaUftnOuQT
nQIqgSPCM9nvVexYRCo15dppptAkWyYes0c0kniBf5k1GA5Yr5GmjmdJVT4x5qPN
RM7cxz4bzDmls2ahWxYBEXckYSJhrYyFduk90cTrpxy/jylbqvKbJa9YMCBSV6Dx
BK8G80ymcllO8nPpg8k+UQlIFlZf3hwulDD/kriaKpqAcs/ZU5gA7WXNziLCzPN3
EuYVcYfNelowJlWRBkHUlSFrqYOPU5c9kbTbpZwjfRfvOAFve4qe7RMWhzvOaGIj
AW9hSMNK0aBTOfUxdJJPUYoNPYxU02SjHWcSiQzy45t4F4VoM4gdr+I91ib61PiB
mGyIfUKZFdGpNCr71ITAZL+gdiNidSez6hIk+9x1FX1erJ/RkvUjwQJw30r+PXVG
RN8mHqltKCrE5ouTcpvlxQyuKBfgor9GHzn7yrDOn8KlhERzoiYfp8YfSt0D+gXM
qiDicfCW7ThBkbv0u951LweoI+otA+GWmyDCooaM871skAky0/OwY4iNrzojt4Xz
ZALL+mUraoUF43xFzYQeSXeDpJ6sHhv5GXSUU3aZHIy05jhjWjWazFftuC1F7zo6
F9NFXJ6gNmnFfmPDfv97xVqyPopCl3T+vEWjYmQiklksXUEY0Zeh7mpkBJ9QS6ZX
uLPJT4/ZwTkUylnrODQT/DA8gErTmhU9vFD5Vo1watqjekyrqR/HO0b9SZWh0u2Z
PBt2waiN8uPu1Rk/W32cHKkpSahWbkE76EUcKK6UPWJ0jpjymaBhExuIdz9GUFYT
cp1fgcoAIjb8iomvCuUJ3dEdyFKhgR5cbeIgVh+UvIlSx/cU5vINY8qv/YezUUTV
DG7H27/TA8Gt46YukWMFbbc2zUkZihX/GoLpSC1fV+0ftjZAfjxenJr8AayYzSCV
J2kdLOBD4DUuJLx8Y3wyTsyr+NOaF8NZsM0R9b5i2QCYOVQ4mvGo40/Pvnk0kbTX
1KhKkm5ATubJ34B/WAVye4fE64R20d/6Tuj7RNriQf+Eqz3yj+PX5yadWDchxwee
UmzX9IgaBO28/aMl6nEvCJ6eKnTXBOxc/Xj7zAN9i7StrBcMxR6x/KyYEEqkjo2B
2lCfq+o/ZI56YoOOcGHmcTbdLKL9Pn/WGkdzdPdZC/jrAUU5CbBjVuZAwcBxNU6+
Kr2TSKU1F82MpmtxW+yIFWg+GysC+yq4n9VcHCOBJs1WgkAIGtkYTwA0jnb8CfMQ
ykOI3rBSu/k9wWRMTsBSBXof84JC089FxHF0UUK56i6zMGJDEviQw/UFRxyb+cE7
5UIkUvqoWHTTpPxfH+3Zy9gTss8glgNmmTj+FCEig+an8ipR1t+XdSciIsIk1vNr
knRW9tomOg++tlMARXVycfR6QQghLSdoDsS6e13fQ7sQns4BxDhxqegPNpX2ngoj
lX3FI+3fCIq32XER++bcLqAXbCd0hLSxM5wxyK8g8yvUbDTysX/N0nwxvBd+qmh8
c+1KlHxAGx3HNDBJ1M3FrjDq+v3a+mKYdhtnLSFErzf+Vjj88KuQUy0X6b8WRef/
cjZZIN8d4xe3LdGijx1GG88C3SkSXs3Ny6X2VfZIbfLxJmdEMhAEY3He9JNKq9RA
5tqjlLbjivH2x7Au76aPEV5BDF50n1vG/YPRTx7SIIy8KPZ7zPlTQCkc+KN6WsGT
XRr61vTohUqtvWBrvOnEGyHPMlVKoa//cpX7sS0//uAimK1kSHPeJqreGbUWGJh9
142I471BIvAnp0JhyUbqKHAY9kwgGRqpsDGdwL7YOaVYIpyUm/2aMiul7rDE9a/t
2isqvnm8Wo9PPw8z2jZCt/07B4y5W5wLw+L1OPh2ZxgNgdCzqL5sei9YV16MoEIK
/j2Ow/dxEDmyWwiqyQJfrPYYF3N2nWmBIiWQVqAbuY6MyeQcdPizOLyIgjizle0g
dl72OZr5+mZ/UySkx4C+bfsoXDyhnZWHyeKFcYUd753RNFPz0O5Qlx9in1Pit9gF
0fFIfqhS8QcVhJZ28hF3DETy0E22WpbsTkC50FG5Rij1jfGVHalaKTPe1XrSuvdu
QwRQLqZh7x9rBgSuTd8M3GTdj/r1CbXhhClsEe9im8eVAEq1KT3Vie9+e2X7lIfA
IYYM3j3+04VxqebYiZpOtsT9v79ZYpaeM5KSsRTIyeI8q9BqHNi8phfQhtOi21Gr
nvEbBsBSo9ApzpYDAFuuoW16IkEXo6ZawnGwTX/T6lMsme8eGjYL9zBT5ZxMaws9
b+o+sj2NBkjyqjnBZJq7rVLsZvUU/RODkXbC1EJBlp0/R+0wB0sFnz+fcgMZqR8U
B+AtKTEj5M/3O2MQCpfNkKFTk9ws8t62cXRlobwF5G9jGx/JYBkiMe80eEe0IzIP
Sbj9Ac++72VYik/eh58dBCPa72axOHmZn1ktLM0vxkDhADqBAc2rN135NI2rtRC3
IKnAmxYwdGpdRHrOlFzZ4CJz/4pvEWElqxzCjdTL6iogX5enuuebqRby9eKZ/cS6
iwomAbqVzPka82t3plNDGfKzRBDrFr9iT4WWt/+HzIdtQ61sKWczGTbc17+orz11
clbgSSoQycEpM5RpmMP+/7jpqASMzZ7aBVl1VeoQLly8N9mDXHzHy8YEZ29JJDDT
52CUWL0A1w4ljusvTLdvWI1oLcWq/9q4RvxojIwvP/qEGJtRFa2nJUbSdaNdiybw
GQ1oMN9npolvUS034gVXnKig6qkHaUMtRMMi9wL4Na4wywHL9s5dZC8P6TltrywZ
GwC5Oh8ICJ4K/b6hxgpTYDq4Q3Pi8lnTNSYOmvKU1AFkiybFxPY80m0n6qBBowo8
RF+kf3seE7YqilkrciWuXs4UClyuJsJiSF8VjlCpbmdTGU7wGgv/2ACVEb00efgv
g+Bi+CKHvTleU194ePoKDYpYDk0jjE6MTW1sL8SKnnQt4JLGxQWMobiEUu26L1dK
oH3E/Z65fd8+3gYOr+7FJc2pzA/4PZifE+G3bYZrfJABZc8ZgsC4fcnB1KbG8Y4h
XQt4RkjslBQf8p46WzPuZn2DzkBLo2kRg0qopCshZbnT+gkLRP0H1mLG10qbWyU9
yY5R0xJ3X59hEhh7AyMJSKLqUC/SMDnUnqK9TkFWa+Fj4AWmZGeLhwX+4L8yI6WA
w2OEcmo6bb2MH58RAdbFoJOXwuL+dblt47VNBnofkuDJYB6NcTZYyXAPrfNUKX3L
R996MQhVS2ifx5VQtFdb7rNPRIwrXMzkBD7AW/VyOZbvGToysv1lg7O8ra7jy5XI
CLGrnSiRNFJAK8nklFq/goR8CSA6LLnprO5MlviZlL4M6UVqqsgxyw1uKGp/7kW3
A422PO47yrXwjmnl2y+6ckjwZ4O9nanSIWeCq7y+aeqrFYQErY4MdpDKL+pxmPFc
MeTOnyLU9sGB0Sa0/a+joF++pfbWKCcl0UgNUnmqjUrQqjbBjqta0RU3xq79+iaq
QZVj8ndhTo6+uNjZKN0fOf6duvNHeKmnA4+e6EymTTDR1INCpt++DyNZG2jvi7dv
pHTk5Bv9iZPsAWjaYWrGHnbLqZdhIsBdBBViY7vkshzI1nBp23VFfm5wiqGwg7rN
NevFJbJsjsUiUnvt1wHSwcpCoRu05woKB6Cv8iWeJtFozeOI3bn6P7nzESYJSUhU
68ea1K0gAqdR5PMjv8wG1FxDlRa+ZuTOlV+42wnPN8EEFfdkyJgJ+FBkJR/mfQrz
X9I97tL8KzrqcQ6V4pf4IVSjpS0wbm6aFO650bylARu4Qb58np/MtNcfc3ZPbKHL
QBYn/bKfjwdsHnvIrOknsfiv3ukjon/RgstZ3PhZi2JV5aDxEzdx4uiHgV8ziq5X
I6WN8ewkoa8ZmPuXKajM6wvNrFdF82HI4hGhvc1J3djQEtdibPImQBErNHBVKizi
hAuOyItvnnf4jDGw/tokWEH9IEx7sZCuqrt5avr4i0RfIzbGE5x+3+Ypvmz5dBSN
IscaMK6Ig0rAcmzTcJIh7Isi9T1ryUsf8r4lGPSdQINwJe7EylrC8Zl9U7bv5iNb
VaDiFPH3aFK+nJedMYePCHFFHqtOe5lDtAsahkVbFjCD0YMGgEsyMBc2rozslNGx
+OKO9yf1bbSLwE6s+9qVRDm/lJVsOJ97hmM5oEcGI5KKj9+lxMEkNY4Cl9JusZn/
afuciKSGBacpqbl9iqKzUcsICSvZ0gtWQGTnxjeznVo+qIbml0BNDWcGQOjAdmYl
8HmMAL6kjl5VI+mOHQMyIcXrY+yMAOb5iEXb4DjEaobvUOP/AER057mDYQhKXUFF
AheeYHMKTrALatS4KtK+4DNcM7pFn7HhTagDmKUEdp2Y9ebFovEDvdyZYc6jbC5t
mm/3JpQBgZY9HkhrZA6qV1Oz0gdnVM2W8cUiH7rXBkDY0ZU3JvVaAp8l8wQsIGzB
KbUJ1lCGkg1/jPpHcM3axDmGOJmuSy+NQHVNbpu2zUswYywoyFa1+HE/kdmJflAl
vntgr9WPUBKUeX01PTQwEbBk6koy0Te50QAlE5N9q9AS6RWAfK8Xpr7P9vkGi/Vw
uLZFA69Pb9jx0Hnc12dkw6eBOceXSSEwsEFVrNn+5p3u+08INWoVsSDTNSJ0lBA9
lq0uE/xcHhmE+YakjO0KxJN+hBlpUQ1WypR0QUPDZF/nmIeITOXbs8KsMImHiqIw
DSeILVj3sgVnk2aMuFEavOA3h2fRgPc5gKX5lWW2zl1z4vDV3OEf8UPUHvQpxqtQ
0Ggq+OQPlxYa48DbMJO58HdjU0sGdWDf8rQH7CzKB8xW4sRWhL86pX5R5WfAPaLE
9MV6Y3Efd6Geb099E5PsHVnZwaSMZjbAH1ctVtyJ0x5fVjKCv+RJK3t0vbnwYPcO
otdqyRyRK6vRGoYY5RbJ3uWrFGDKiEHMnslrcTThwCOBgjUKeUeS4UiVy+pxDcr9
+GR6KVRFm4CkUFNuc6TzDMAYN+V0HwEECfxkuwXCbvSM7MgqPSUbvl5SLi+ZEYVu
0R967LetBLg6lynhAVvabYJqWc9uFW6Uf6s3FzHweGZUSikpIwFDpEPKMWLmgJLe
OiR8SDGPw/eShNVY29HNlY8C8AaNWWzoWHYYwALXQ3LDkGX2g3+lYVzZzzz1RqAU
78D5m3EMDIwINJqvp4kkzYeM6BvFULzqJLw/iXYBJiMnd2K8M/afIX3+VHT3lSvj
swfh76LFbJ9ec0zM9YDc/KE5GxTIKG26SEDds27Ch9Zq77xHFPH4ndx5QhdzmvGW
LN/dHqOn2cuGj5wjXgogb3u7O6rcA84NyuJzrJyl0zDO+JPOVLifFzkc+hUOSBFn
jWXeuGKXzVrC7o5bMflEuaof+/393lmTVTIl3Sb2gK1RGQ4mmEKYmP2dSlMrZNYF
HHydKOB18+vvepHxjvfifWgXeMEKyCbo9Yuerw2XTsV6zK0qXG8fqY7KPM21+7kL
qWiZatv01n8gsQV+G4ExHzMG8fV1K0+9S2WhBsIbZloGpm4aqDufaPYCGHw4sAx6
oXI55ho0MRhxRU7z6a7a3FolVYnXjSk0IkhY1APDbuz9QTkJIPCMNuxN70QKQLPb
V0xcM3WU4GCCQlEcNh29wsyJX3srGlWTj48UheziSmWgifunldJKKTOqDZpWfyBa
WRwOcALCRQu6FAf0A+ztskPfAqnecbwYr/gYxsGWqvWltQXbBTENvt2bPtG6cNOZ
M+eH+xmxgrxgs599pj6vy2mn1sRzIs5h20yAfPynxKbYtGHsqF9YNOh6Vb0Xkl4J
/k3T0sU+IFvS92dOAlpnWX3VoZXx84ZjnEOwrUZFS3ZQU7yp/zzlm5HMYnhThezf
uRtTri+BSkuVMjaldiWTwQbprwLgUVXOl5RcdDwSJ8Apv09/7VlcqLfHb/zd3Z0j
Y7kv/K/OUk+8/HZWo8cUxtzKJohdrUWsKzl18r/81+g+CVwsqet7XRDSC24W0q8+
N4P+K+28AUCb+pEC7fobstHj32ecrjtrK+OSGoeivR4v+b0doREyxhq+ATNO7ppN
CjofWUBSWkjFwU5N+DLWQPUZprrF7ebekCnZYm4S2ThrnJKt1z4YgO5Z7djD3TLt
fd+cav76xTxBWf8ey8g6dKU3dZujr8JjgXT5qg17iD5M9+nL2QF+rL6JlXTOeoXc
6AegivOgEOR5rBecHwwCq+HzlDhToumTXFOUUoKfcng59A7Fangdqc+vSVN3Enam
Ni57A404w77a10bZPtLXGBmuvdNExO+C8bljQvwIUvfKlSebkG/rxE2E8ZTq3aKV
iDQErKm68lnKW1OJKdWJFZb8RyEOZbEEPpD53DCUZ+fxjllBsLJV/VYhfi7Lu8Rc
s8v7onLaiWpSRoDj6Qto9Dq3Z25JKtZOUeakEF2K4XswzgORKAqZEIUQ99vvwf70
vKF1btclF5kyvJZcRxJzqwyTNHOfAJnKw3O8ntsf6hl/EfuXvneFCoLIoiwUZdPW
HlaSdJ0JMsF/9HwZ2q6SGx+icmjY0EYu6z7WfWsT95FduRugOhH9jLC70iGp1saT
TQMnGX/8QFGZN67GYvNPn3ipA3/JK3RCeIU4tAMW96NqDsmfK4k00zU8phbFYyGS
dAhiS+pjUQwKmsZdkedx86qseCpnL+/LsfeADqIb/0oTtHdFhW7g7JEJvF7c7LGE
1zwSSIoPlSIyJSZGF8ZC8VmakoYAkO8Pep05hTFeMsrsPb0wErxRcqCGNhArfp5e
YJ6m1KoAZFxmG47PpcXDsD/k5P21KzVayOVciyOxLXUWX/FpKtizFckrDYknaE9l
esWozWnrXi6I4DF0n+pc73sCfKuhnUnnpzpO+fsE+ub9B1hVeBDzWM6X1l0SaiHD
QJOnox+9rh2t1fIl19glLVJmj3wXpnCQ4RvMbjuyWRXwZK2g1za5ZsrRtKghTskV
uy9e9gHGBTxIuqy0MoE/9OytUjwJ7//jW9oSLO6ml0gvQRJm0gG9ani/eIZ9xk+f
3beMeLLAbgHdKSHmF7v51sFkbU7pBAeah0oe4sFa738A7k8VEFfQ9I3uuN/eOjB6
UMsOf+NQ11FRw9Re8F897vns1GinZYN51GvtX3hg1FjqKSQJO0B7OYKJ3xYUUNdd
pg5yld13AeEFZjX+r2BuYp/EZCBq/ueK11l+ZeAq1H0M4/PVyJC07YitV+iE/DJZ
U+lE8ub0aN6yN+Yc2i85hYLlO+z+mS67fY83kkpUTzKHKihIsji/9E1IU1b3j3ft
7dK6xLRPCWDQnTlrCKVPfYVARoSvYxVrcdw2tblx/z3g3aVpSLcrZfKgGOqXPkwZ
tHnwwY3I78HXfKFLA2Ra+HzBTCMXiubvu2HrhbVh5sbcsEg3uFHKgKiAulqmoMpF
P9w878QqK74FqwX31vtwzH0KQQ5uC8vZb/lDQGLy1BpFzAbecM51t1a4grGQTKxJ
L7mo5AaZiom15AewZdEUhOhMyHJ2+W1SI6rxH6ZYiSwoYtSwaHtP59DZVQ52w4jB
n1Pcc4xru4D3Bp3+RUGIqbRcRr0fXFirspEpYFUI+4fD8vEx2W7+vkiOMyCXDugu
8BJzeULB2kz/f6sXXatTrx1PIivn2qCJd8VIPzJdzSsRaqE/jgg6zG5YkBKxWPMp
SY5uZ90kNktfui7RZXHY3p+mRrG7MJYkiirUQKsJqNT3sndty4s05A/gbEcxxMhy
NWsVCyL0r6gkoVivJkfe00kXeUxFwsi595iBVPTnFfxjzH/lFgoEIJEgy7V8DFpT
ddO6hGOX3/TY+DFyfHPeqfK1K8Dtj4JlkyYw0M5uJyREH9Uwx5bC3eYrRoFLAkOA
JVK0J2KD7AHwfLM1F345YAQnQf3hFI9KweA6PtgmMswzhSpcIeoJlrkbDj5i8u7y
r5ocIGvr0rfmBmKNdPDDv573qyD1gUzX7VF+4kBIiiDMUWYO0hZdi99jj5YcEHSK
l4RJTGJvWcfaI9wQEQ1JL0STTOoHQU2PT6F/4xt92/UoLNXJpgdQHMCvVXWHUj6t
P9tmvqEO1nJ5KrMk1jL8cvxZXx3zPj7T/33QzkuVNHYUZc3Ord1dFmm2vUsl/XJ9
I0/aPCNKvSN0cPFAX82nS76/FlZs7OIqR9EhOdlcSK0rlWoLzzHh9oS0EJXIh3e9
jSpC6ie7y+Qy5DCri0ByuUQWxWDrWfF7PRHgiOdPZUWvmva+IEC3m3EH5IHq/Jwo
4865z0DaZKZUvARpB/LsDa7Sjt4RkRn1vjrYncP64b2fGEccLdtyZC9Shzooc31W
2UL2+zVFIwuzsI+GltFfc/9NOXzWqdaKMdxze5mGtUhSaCu/x0tvDbkjgAqDpH3b
wF2CpV+6QanpKaH4/KmMbt+JXSIqkXJJhEQ+XXloaJAgWhmMFfG5tbMGXA5Htix2
27sGLYB2cbF7bW7QlBLZY6I/3lxPdgaDkUlGfZJvmpagnQcyqmNurX7Uy62WILZw
J+RS7lT7mPLY4+QbtXsb9MnFQV3PYf4MTkq1SkvPElsoGvplV5DHBjKferdE1BBq
ba/RMqQIGNd0CDNvjnshEuFH+WMLWd7AlM99PhK1g//UF5ZPY+75TRISDKz9okNH
rwW1c1TKtlIRb8yu9zcUStHv3VmzUFG06O/3sduPG5vsVR0qe4XpBCUm+/OdsSEf
o3yngor9yamu8Tu9HpB8flBlsm+Fnnu/zwu7RAUIDsNWt7hJRIAxDOb8/ROnIhr4
9xYB2+ldGE+Ux9wYx4UHT0jC0iaBtKk/QlUVtk97LFjfaTPnTWWMcVedQ9TxKs3L
vDGs+jAVNCWz4OKp/cAgT74k80VUIjwVo4E283e4ks0z4OKGKI58YdwVQvGmT6jm
A3q+d+2I2NmR2LCcqi8HUcTS+7CCJLy5ZF7saJ8A+vOnuDiWS6eYbCg6sQ3ZEhUf
H/b4R+btUd6fN9g+UHi8aTp1bkO1bD5rXZlj0YId2R8ANRKY12iIuelrDw0h8ubC
cHbZny0Q1W9rAmpQQmbwi2o/IqXeyoGopPxQFb058G5Cios2MAJXzCHR+jy8Rc+a
22TZLdrwDCFoHyQH12LIZzpwguvEz6oR/BzOh0vknO5znADRXF1qX+inVFaKpxBi
WxfM6/fNdiES1jfS0tQ8UdRBjE6ZF/GFE4u7X267LwJrYoQAbDQiFQuUHB6cHzil
aqhjAI9qshYsQlQV0wzoWN7BJqNOMc3i43aF/xMddwo3clN9bjf1gL08dhsscT9c
OPbbY95+1xbH649FzrOKU8YOmin1/e0AfCXL7yGtWcilBLL+mWdjcOIzBr3Y4d2f
NKk973fBBaoje0jD80jrL+roTt2IpxUb9yfCPyYa1vDNCX3koLFgG6tF+Tl4LuKv
Xu2xvgKexkCP7C47zEu2gdPftTxcxMuoOTZlPi7t+zWB17XGRSGOgYJuJTvyderc
upPTuNe3NY/PJ8tEXOKfXauyGl5e25c7r5GgWDcRI4vP6X3OZqH8DSrKTUbZDxAR
zOfkCwQoOFNhzQOYbfOLaHw4+G/FdrvK9jSfGWTmnc60/k9y5jUCoJW3y/sleauX
wOJFNvfDijmL+z4JNBSCMSgBE+uVyJ49qEFJeNXo8HSws65uKfbHlFQ9wspZ5n5n
/nlALOnNzxIGqClMOJOBNrA3MUaXuzjER08LMmzrGJLt3EgVoLvuHxM0siwQEkDi
TAIQ2AbtDjLQT4afp0p3EXY0F+PTSiUSS9SGcRF6qzXGGp1CIvVWcwBcE8CnGyGc
2BXxVkdUUxdqKHFRdAFCZTY50uSPaOBiAr1H4ADHOy6TZb/FWbHcA7Ubqqmw9xRp
Xq/tHhM3UPMrFSHdKvHe1t3iYmwZHw80ToNyTHXEeowwedp//QGNY31+QyD4Lud+
ZjPHLLQtbx7YfAdoc6ii3DUNOaSSnl9B1Qjv0f/9FH3NOP3pPVJxonTotUaibHMk
iaCG3uhXsEO0CQUzszorW+Xoa5D5zRtbL5m7F541NA5DXfUmHa92SIuJny5VmyGl
aNArc7Dj+v2lPH2Grhc+rIHBpEPy/ZzK72/d5pr6ZjBNU455UXh/mjwCPiGlxjo7
V37F4yrwhFCX48SNdX71dWbTZM02BIaRKrW9qYuGFZDIF9LzRn0ybb+DGdG3lnJQ
IOoTddLkX9h0mTBbF0PxeRKmCpgYYwx5t9AGtuxY3Y/5RPhluqfHUp4uQNBgbiob
FK1YA4XgAQNncJX+Joq+/SeImzJjwWePjqsQh5Bit3ny+Z+NDMBwnErHU9/R4gCg
k+T3fpTTsKmSeCE1K0j7PupPTPmnUSY/azDI6R3qR4A35XB0T9IuF0oFeoSAz8ZN
90bfEhOdOagIbiNtl9Aq8lfT/f4ukNsEslXoE4CtbhsboCkczsgUPL01WyF2eIHf
TZmjXSBauurn9aABn2lm0+9HpKQh9E0GnYvlW42SHdp5DVbytV/ABlvpBgoRZs8Z
axUg6A7L1Tfq7/tFYeakwGHkcCpd29Zipr739eQjVmTyodlRqM/KAlhEnz9at2fN
KbBUMqsAEeR/R0s5FAtVj/FwyMHCE2xcLcOFtUmq0XJMteKVDBQfq73UZN1U7aDQ
0HVhuyvWjDH9rZBeBJZ4484m+qxf6U4t5wBkO1YLwM9hg25ObUbxt+2Uo723WYry
zvOnwkjQH9Q2t1Ff6f8utOR7VyUBfPbtT4sOhxg49ciPB3bRtqo9qSSpPIxYgc6j
ctNCSFH6dwjOfJWU3/3mrLCCIN+VPvolJOdP92XzQ1gM3VE11xlg3JJv3yFSoIO5
9Bj6LHEdVOQZReJhc8Qv3rH2RO8rdjnKsbhrQkgvqUQi7bxhLyRe3GP1VuJzuQkW
vaBLkYs54sKXbkOExPFSMJFwSeqyW3uNhcvTVfpL2EdZuhX5dECKQeRAV9NwKnwA
nk2SqaV+5BKkISumbSrQJ6dkVDq1D4BqRHkdVgIbAsT/j5WGINkMq7kkvIFFRxkC
Ush0xC0Ye6bCsnTbWCjbMaETSK0n0CZVZeRubPcN0C/AIncmsl9aDAKoU88Fo/OK
5iM4M2AfxnIG4rsOIDlqLxznBECIEeOACVzIYGHu91YhC+8xv1dtKWVYCOGrRvZQ
PIlYcg2d3xShAi2OBsRYFZ21aYtoCCB1Gk5/x+SYQrULhKoid1lVGsAzZLrHHCMz
RTvLo08pf8z3GipzeDlUUIArrwvyMlK9qYOHAjkcSiZ9cKhEYLN2rkeUUuVJwc8R
1uRs317xKq2D70J/rMm3TsmIep9/EDys8W1fyzwg0R0jndgbhzVNoToClCq7z0WU
WVomnW8Vlt76kbUamIgTVeWRrLuncMOQrgEEGNYA3vgtSpqHYbfdmd8HSYbpEF2u
PRl2Y0VwhrFG1hvwW3tM4tNDN6j4a+0KvU074N3BpXpHYLmXn4pCOhUnvYUZeo47
Liwq4uEdiz1EKmiSZuXzudiAW/2d+PahdzbD8TDOnjs3NXuIJimMt8dl26ab4FzO
n+tVqkL/4No14wmA0yEdNt5kjUc7EeTcnGqLipyUs2QCaOfQfmU3MtB5BkxZsCPM
cMa5BB6Faxemm1NBNxZSKiFnKj3tyZSDLU60pZ5YJLNlH8QcQJ8Fv3A4uD09YuFU
4CRJKfpnSfCVs0E5AcPs7LdnGss+MpsoI2hXYhX5pxIZ2UXFbKSa/hoQT/nUucJw
2nVh20mKr6ESbnjrTkDso2066h6nuAEAw1ZHZ4+zsKtfvXbtAXK+pjtuNrbWhPvn
vSnYGlR5MDv+KG3nSkpQrQnFils+S2TYjj8iiKPq+8kGo9jFzWopmkH/NgZxqLHH
xQtLr5sBYPqNzA6GvXKrd0OM48XW3popEVh3Mf1cLKcJudkFGS/194Tjs9Kd3rrL
eZJHf+yApXYl4OnAqoKMWne7p2UJvpYK+FSupXi9nBVVBsE/H+FAAyjqBwnwtCuJ
HW2pKNCVJzXQZPjNgheebPct9av1QHAWnHtEI/GA7+yx6TUWGpzmqvsBxYirIItk
z+TZoJVK1X7y5yRv7FPJZEAt/x8imjb7sIZLVv24hr5g1ICJf+UmKU8XOtOk8m9N
Br3brVCeBT9vLY0qi4FiisB7rIzGtfcBZEqr+9ZeZ7i/zgz7vBawNXTUE1JKhzdw
jsVMy+yFjhTSZAmRr0Y0r884v/NO2ylLZLDXUhVkMNVxDHeSnrQuFHnx7wV41tYe
yvwoOWmHpEUipD6gu70H/gWS6aJud8vWQhgxLcKogajX4pxyd8dBKMVZFOZ9xA9z
czYMcspbZVAJ1Cj+EHrqFcQgJHMkZtuyM1KxV2WtOsw8rmLhXCdlPCpnjya+vAjC
lG95T2DXjoaRxc/8EFpZeTVDPqD6krVZz0rq6Xn0vSv30bp1oHUgvBwbdcSRDoOj
JLUHv2SXNgJqj+H82SZLh8EGRYRbOwAFIOFcqC8b0sauk6J8rped7fj4Gju0GowR
mP43FJxuHEuODXRDFXSQYyOArVdt7oAmpGdIkAicLXH1izD2ELhnZ88SE44p/Ja0
SjMhkud+sUdHnZeITOiwkQfvCd6ZWRXr1BfpvrOjibqF3uGkC5xeHzBFY2FMZCKq
V2cF/Jphdo0fR8vRZtfm7RY/U3Qce7VeU8EtN6rRsvpJ0+0R5ObuTMtO9L4fbU55
289dzn192SuHZN5JIurREUD6KTuX0+P94ylYmpN0Npr0BPBeIXmAjNgWgfLiNwT9
MC2IpGG83ql42v8hb1dwRm/LXRtdVt24V4odRlKetEewEK3J9BR06Z+rz5gOqOo5
r07aVoE/CYQGe9M80TF54heDdtEr6JQMrLM+t5FI++T/+eicmOc5DBXlKxaVf2KQ
VS4UbifoKd4TnL3ya5Cm17wkCqmfQJ8lyws9t6REWRQ3Jqalyw5j9Cxswp4AOuIP
HUO3/Xjrvvfhx3aCYLfwJGptdoqdlFhMEz3vYfT2+DdWCIo2x1JOpUlCnKaxvG4p
q0stts5ifn8zYWQ/OgRPzD4PKqDp+Naoq2QlcjKNHyOrEivD0mq3rPYZlR/0Ymg9
dk+v6eKROsbc0DNY93tsJ5gmIgBUfKxLZLDnrwE64D4BsQZ9EC5/y72H7mDNNF56
2d3Lk/tQ2AIR7Qi/kTvE/gnsjftmI8AHyw3XOtkY4otobDG/JtY3/ffsqGm1CvHO
1pGH4DlU6xqni1cGbbRKmleCzvZC7tqNI8byqT8ZwcjaTjdMPO3eOea0P8Nbus7Y
PivTHt35csLFYtGFCfR1gQVt0lKmVsuzv1eafdykcuU/uoBg54w2WcJ+G93EcdUr
j4z5myJqbInMPsKBJGewUv0Ob+oz+CQsFHhB+s2PpxOIV7MaKk1bMEb/H1p6kCgv
fw+DN5HUUuDQLeNDiCthXgjWw0xV+EjAa358TKYexFPyMj9fQfOJfH4iTSTpo4yD
hDdH60d43Q9KJQlxW4tHI9MIBTgcgOFspkpU0fZCHWf/68vymTyXABdr9ACXBzZ8
8Wa6aTXfwQ47ok2xgakcatY1yBcJijBYCMMaplsaDGF6uzQK8KKOHA3TWUss9/m0
lpcJrxnQduQ2OgteppzuoLd5sXgciv4QGdoBBfrff9kaHJ84S1nJq9c1cj+q2Cr4
ytB6pBM3bq9I9+j+pB7pRSnDipO/LXTibXhLe7Oa2xmDVZTWzAPBca7XAD0DhZuH
ngznHpQnxtlIbg4xHAX7Rx/JTj1E2DWCw2tFHgQiZbv95cxmpGqnvn616CaqWrAN
+WKUTN8nmDKMf82vSz3fsvyI3vmTOH5uldue3OB05YIuqcbf8xBo28zsL5a+xIEo
jSvy/ra1Tc1nUARlws/EED1L6qKOgEiAKCYSuP+BQjvS09l7MUu02iVbVdowxpxz
TohW/5fyHAKCJf+y+OuoEPyCQKfMCbxkRLiaDVwNp2D/OUVbnaiAOCEAhC+WdcMu
CS3o3sy43W99etxB4t467G2Hrv/3CYJYQTEkwuh9S+/a5Lmptd2M6Amfg3vgPYn9
VQAQY4AhI57nkeoB4lM454xFPWB8zAQ3nNBvJ/qmCxniGqR2XPH3CJOsGLZ2btUc
0VuFC0WYm/TcecTpM0qel01P2zClIl81U4gz5EHrIdXPJoHZMr98MTS/OuDHYIGo
jBuC7QOZLf6wmK0kYY4hJ6geG3NvhP0587135Y0dCI6IzXMsqc9mrx7ngxIYTtAv
c1lbUi1zxRFf5MdAr+2WwKq7Y0duJq7EMCq5yQGEcVDiyVGk746m2UkzilJD5EJY
K3h08oLs72lwM9TD3yRAFD3YBrDzPMWwK/ckhm6cNm8JXEspJIddriLwz/AgbJAk
UFfMUxQFd4llHWkJ4XYNzK5jsta06l4Mu00RTLba+2qO+TmAfnQQg2/bSSFoYBfh
JxRk2Jnn5JdWQ57W1qD+kEiiefQs7Nq/Y7u1Dy7BdNh/FCtoPkN5Qkt0acFp0RM0
MbLDGFf+7NNXx/XcPzgHggBoQTtjFzheS4Ro1/4PxrM2dKK7dg2L1TJK9BkfOfUd
MgaedNfpAZ0M0/2WUoZt+8LwPmxDqXaLT0qiI0cs5740zWhj3BbAFSB6tXh4UFeV
xB69045XW/B/uKLlJtiDisCXOItLirA3HAgoDpQhocD6swpPIbg3aDDrLX2HmrPy
YX/kEjZP1xn18KyciUyLiJcTN7FRjTQzUQSpyUtkqylo3933jaobFoDtAIEUCAG/
Y9x+HpekXSqIzIzXB8I6JgIGQkxAo48llW3cXNeu6yzZR22OracBtyoMGQEnOj70
NCWWxCriUBw6lGaISomO/ueuWpNq+zYSClw0jojmoBM9NEmSB73kETmr/DyIx2xp
2kd9tedHrTAEgKbUknjbcGYM63Gm8f1yYb33R42rm+GfOKYkLNgfK8d676GFjTRt
rSViUXgJKu20DSYUeDGQY6RlZqGsQCP7UBnoAwyI+3Hj4K2qZkAz4QtOJOjKun5V
wfmU8KTDB0+xNohSv1POiZycCcJR3hSJzkWzJqQvS3YQRl9xLZW+eeXL73ae4e0H
0AXv87YV9THGrXEGSH2yVX45jvNsvVDbLPN2VZfIFQShC9xLTPlsaCrByFf1pVdS
uH+/P5qHogbkJh3nD7bUrPq2cso8UXMw2w7RxtnWPok3UFOHL9fJQyCy2AhB7g+e
FoR8o5qeEIxNobu2xOH2iCJnEfiUq7698kumnAcplUc9ahSYSbvkTETeRyyh33+w
B4cKnuGjiNtVUe7PVkXzWXVVQH0XT5iM6HBpvLwmgfPD6c4bx8kg8j2/wR7zYlY4
qNkXly0ueBrrG9OO5+0PxZ7TySshdsKILZ4aqxDwb8h0bxVbVlKxWS+2WtfUrSak
2rx9Cj11jmZDw+pvqqswKyfdzgSBprfzdi66tozZYpQjXtuK+8Pyo0lodTvqv5ut
SwPRpuMFtSPPpJE2q6uWa4/ZeBMpLgzOH0/DtpZZQVo6G5xVC/PCB7gP68a5BX+E
15CAbfRGBOkGuMd3pZhd+tc/uRAdwp5BcbIAgJX7DB8FbYccX2qyv6VZW/qmqRMY
H3LPRbDfvV+9heKpk/NjF4vk+FQY2jl9/bSVLdQbqZFgCJn7xiDGkaqVg4kRIlcV
HdcnGnz+e/7c8j0aqOXn0322UajvaEzNQ3iK4cp4FsQ8OZzCg3JPQnlwqZv7vn5e
rE6AVLgvggg7i+0S4pznbd3njop8efUSVPgpPTO3v4+afNnjFCIDuXu0Ag4bbJ6E
s9VjJG5F2kqneWl1a8q8HgwyeoURHK7VPrtrpqN1Z5XSayk9X1eLntBUpKZuxniS
7Sj1eC+VUeu6ODPIi75dIHF4DKp8TjKGZ9vTHABKN7M3GV+DmhGjdyeXUfcLQjqB
8fjcLRT6XYFm+VIjfEA1DfzMtvqGTjVlgYSGX2ZWmsXBYRcw95b5GxM1PpnTlP0R
BuZz7+gPIfIgtLxLxrzyIaSYtDgQVFy7afPugr4rakOny27KwsjSyoIYfIJztXNj
Na28gT/Vp0Jgpr4rbyYvnwz01nDNsCWKtvCcHh7MvA2spLR7IqX7CjswSTKw/4cH
/7pKQpVj9OQPMrjlbC0QTWt7Y3GGOhLMbj3ZbZWZpUvF5ZQIUVID40p29Ovf7PXP
bKIgoPMsKyq+C4ExDl/Lzxltr8T1e7HUwU8CsbFpA+mV6RpjwJ51SCnyb2+PxSdg
ShSvyYdAPNEq4PfQZS69WNXurQXRx0wwZ9OAdu2fFN+qh4tyvYzM8n/HZVt5fzmu
SkwI2OGzw0PfHBBvf8fYvuhbuFHrEh6wyswV5eZhMtN7yBMnGbQEzL3JvG41FZ8S
IHI2rNGxmN1GL2Fn1VnArQHsMNLdu4PJzqPi5GK40QGaQu4ZOFXqjabrcCD4dIAI
ZXF4MjOncx5Yral2b952HKWP29OCVX8hsIm7QHG/bYR4SsagJx2B8SELpRn2F6cO
zCiGh+zcst0D64+TL2c+99+4xzwr4DZD252Hs28DtYmvtjlSML39zwm+RI5pjwon
N2/GEqPvoWtZ8MDL5OsyYt8jePfZRLpLeSja5p5tx4I1WOQKlzxj/cAAdlXIh12g
khDERy2U7JAncxOZxUm88O7L9Ply0yz/XwMn/A2s1FZ9Oh4Atn59LuBUboXzT169
QUHyjBwQFeVtu+OFPIyqgu9/g62T5L39gzmtGvGbvjcqFElyjCve7bNdTaYfDECs
tsJg2p4C9dqbvRwQfEmRnuxWQ2/+i+tycxOBrqI6HYh+TuLBcU7wWVfhYDiluvrW
QSu8EPctpEYi9ssPS5FKR9fm4yXV1g6Xsj0TQF0hQO7LUbsCs4dteQHgeUe5/ZiE
eqja1T/X+d4YuftxwLy5jDEm4HQOoebCFX7Nc8cRZC3O642suZTdr5wgafy/RDqe
cgFZ3gjeXM0pz5z7m9zCTtwb1qhFyw8ldhnGn8fvc/M3Ht1M/CTq73BcbNfc21jL
eSdI1DCL5A6s/Md2FNlzJT1ue63tHWW+KBZjvYz1BNhbbPnJiEckt/xK/BoFQC4x
ot7gQf2Xj72ngGhPpvSJYXAjvGvKZjQG8CrhJDVXomIKpSNmutTuSocM2UTJVIcB
Jv1sfGGFa7blevEWVfDLbLnszu9u0QaPUY89hDRUifhkomEIVWrIlfb5SQowDeI7
jk+tU71kpHLUQZxoDcNhl3iATzCy2+t4vW6Do3Ca3VxWyghWZ3DgGgzNlamsER8G
5B9UhflQ9gYCu5JOVYtci+0uGEJ9e+Mj4QJVMLjMhXMbwOll1zS//DzOHkpmD9eb
6Wy9peVL7cD5cL/W5Z92IQuAkEi3T6GJfimJWTN/U1G8iRnhvh1nHymFCrN5ibKF
yMLHsk+EbX3I4pSfD7J8hcn/C6FbiMxXTmN5JH005hLZfbWP2JcKhzFFXrhcDwmS
Ba+9pRPV/k5YBGVUxoGBriIi+VaWSY2IqgaKuwtCou4sV7aHihiYUAt9+w5vyjpr
I0uWpeXEsIUWi5up6VaPXtrYW+QRJgJ/X/AvEvBkaJUP3rsAyCGVMZjeAVq5PFNn
yNxAgGYEA4iVsK53J8T4pgu6V1GhOMEVzoBTRyXhsY7INNyDVyZ/iEA8A455admv
kNTqBW+7OD+18yHHvbXwGHB01C2NSgy+zZfkOpY2vTfmh1iUYGqoLRtrznmvK6yZ
mnWPrpgFiOWMqxhZKDZhSJnCURdp05HTfv+1vEyHIw/+lmSCtlbgnTsK1050Ikj0
PlUvJJvF/CBytAxYi+OYauMU1Inebm00WTPBYKi4zwCKWbzRv+tW7sPIKylTCuWx
0J8U9K2rSDjDbfROUlTp7RUg/AR2bEwyIKL1tYUFNtkrMDOzbRU90LxBH9w8IZq8
xpgWTP+xk8dY8Qo411n8BXMQsbNtNVK63ixACUrPQ7dwbO0yGhYK+OugXYzv1+Uq
IpkbkgiqWoDSGIAlswYj/pDJdshG0vgBP89iaHOWPUtP+tD4i/0gb8ynu50/IHxj
Z/ibjW1OhQTZQgqyGphG7YKlVn61+sC1Ww6ovPQznxjnnNG89xoUcD5/eNsivVYa
pz1GOk4BSZH3HQRxn/y/4U9lHgsrU0Un3+j7WvwseVTpEw1/U9bKcmrKEd/NIstb
ASMH23pof8QaNtzmEtwum8fgxmzDxuO/MCX1zUbQHlbSLRjGaIFecZ6qxT679dVN
5qDVxZYga5VJ5sg9E+DpdvfaxXot+uHhrW9/S0ephUZJ+tknkWz+2sgTgfSzujG7
UVLOlLA3d9j/CX+ccv1u10pBVf0/kI4XZ0CrB/FLHpphA5M0KZv+FKvl+UvvK76I
cIHgl39V882Wf5rc9ZO/nal3j5hu9xl1x7iQo/ED4NRON8s4alM2hPnwwsccjXYr
K/yzrNDU8bo/PbHm2H0G1tQCWddc1jfLMVTeoCj2siQprbXVO41Qw6KJq2a2sJte
+U+Eg4ErzU35lHsVPx3AbsQeSRBs7L2JSN7ILUwWN2eEBDaGsxleOJVONhfJ+Haz
RvwIRMqp02MyKRjocR9HE7opYlFFFm/Bn3CGj3qQ+SE0VmSZKbAPf7qUGeuKP9D+
IjlSF9+v/FNGFefGWgk/ynNrMwviVWW+96FcshaL7eJVtWRvovWVxAtTcKTkbA3t
SuGlFd50BUMz6ZDDDuzMl0kCgWLE7s+GE8MK/yn63V7AHsZfINK5C1PHeBiqeSLI
JDtyfWFUsoYBvgXI+DETvMxW1FxUc4LNcqjBByHm8d/3ZNp2bKCrsgJ4/GfQpEwX
ywPYv3rK1kbCHh4QNcauCIvPu55f4YA+nXCeuyls9aAj+paY09QpPTOP9BDZscn6
yXZtXXr0Huhhw1O+sZM1vBmP2Hb1whday0N1emU9lVr7N1oIwL8KIt6iv+2ansu7
Wt7npFMBNfV/tlmvI7eTkMdDKQrDIlgnuv8Hyu1yhH/Xlog3aekH5rmQNEAmC6dJ
JBCOi36OqS6ZdsdOntPy7f4NXbevy1wM05Ut/7rFeHhTPtQuFVY38jtij+1h/UOm
FUMmxhsG0/2QPVjnqqKNhwFudmW/3jWOZqdbwJ6C/4q7iMAnbW1N8jOqv1m3fVSy
Vd0masArM99SJjI0ndQyOi3xuNDBzWOxVRr2ZjBCa+rCulBxRnv7Kd4KoFwi5fyX
eFMvRLBWdgRvNwO/E1WQMCE/hNZ7kFYNB4HbxJpxuaMj72GVoV36124HzKWC0uVT
9apjbsGCasx3k3ir1IsWYF1K6T1OkFvAaiyKP2bMemIOI7UMKxVieMFiNp34N2rH
6bUIhm4mWSBNwM2TWwL0Rq7WRcD4yFZLCrb/4Ntwna0CEnwieDN+0Dk/d5XShqPY
Gqm9mp/cgvNQ14/TDfpIpFFhy/WMN9eLlH+n8Cw7Coq1a9nLdDHJzbMFzaq/N6ZP
FvsCPjrCMWVjTEGccQsBlwyZuzsKA//0Y2A0ELVlr4J7MwW/OGEBOEY58D9N0ktC
Kiy0x183outvnzPmBg92CH216nidKVRSdoBTRrDlMSuVKOYOOac1KHzU2Rxgjsxd
Xomgyqz8Gc85hRaRuCg6+tnC+HHy1U4Tkc8IUZk3rNk1coiwbWCGyxVqUhwrjJgc
pA9JnMybVGqMxP/Hts/ZKad+W/tfP9VbJ3flf3yyZfDNiOzOHva1PCd4Mn9MBc/K
nmYQ5LDAWveRn7Ws8rEo2ZFK4nmCNTiuGztZu14fEuKE8GjEbumvrwlyAOg/F4SK
FTP+EYEZxxeBtOjJapQHhadn+BsMQ11xCG8rCaAJkJGrmRt1So3MBh08lA8arOOF
OWmOgTNwvyRbOi8nwt86ZjELUBjXa5XVVz00VPQYFCyOdlNcvyydrGOe6ANnhtNB
ifVJfydwey4uAs5C8t1444cviW5BREvnMp875PPEbt+UOr3vUpzsDl1ouFEpKmhF
rbGHSFucRs/1LaWPVLJowo7tP6b25Hujgf91CYPTWKZvTXY0KWFail4pK8Duf8Vr
6nO8mcgALuDJOmebShGB6dGbllgQW9O6x5rgLle9LSFkK/uU/lfahrutseN2YyFC
KJkpMc69INrH14aVo96Hq8fQdmI1yz1YBV09hHrUj3aezGt1jCb8SAkcxjsGZF7W
sY/vI18DDKrzQqPnHgTOE9/QcyXa6tZFQt9bPNsmJrUd3ajaasAFKZUJ4mFZ+Uz1
5K433N1N3FQMMvA1Q9LAmL9SsGtE4/EkmVXbYM9ObLhOH3tOqGHZ5OsAG7j59IpZ
dZCL49BGoAGOdxjH/SteDpSNWzoxD6j0Q4buLV/nVMMl7wIhScSg1mWfAmCefjEP
kmsSgjkLTP2yyitVRE4068sREvNPK0A1iFHaezMdjPy6eh4WRP8iMwT0uXlR4y2t
KoNGM1BnsXOoln3p7ai//ksK5XpEEBT7eACr/e352i/pXQEKXHqWsASIsyuINBsw
dPz6r8AtXZT35BFn4wIS4XE2XsjXpgcepqn1fKZS6WuQ5nmhuIr+q5OB5jIwhOjI
UtR4D41AYxSPnQ7oIldKIqKdKZatiW587Uz0CZTeHur98dGAQt7X96HD96toxElV
kBdAcjJLQvTaB8V/ulc7pORXltSfXUg2NknJ9I/HM2pzGZ+9eZwap0/Rq5beRNG8
0p7A1n3AcqZfEOXpowlPBJfj/tVJk5omMAxZyDCX87/hCzqFMr+u6072icikLUeA
1dXaSVJlq65WSf564S42iYZ7YNYXirm43K2O6tkA3bSTxzhfChhf+Zv/HwiucyaT
GEJWGy8SefB39k+7z6MSY+Elf0mG9FrLfxT+zB7XfyQnmoOtTb3tLa6pQzj0X0HD
kVE4ISPjcSb6KAUKd0fHOCVBL0+MZsZdiwymf8S8m2/mmsY74oT/HILfo9E/aQ9D
V9SWpQqGHcDTkLLYgCk78hLUyIWVZyM0ft/shgkzctmGHEiXfxO0dSKUPjNbfcUb
qKu7WsE2ux54WzfxxuOHsUTWTlvHptrxS3QZLTMkjeQ+1JMRsk7Qbu1LF6IkOER6
i3EWCd/QOla2p5ULhxtNaRwGkD5I58lUhR1QBurlJXDAlBcxBZVKH1/BDdjSzcVn
nchNVnbU3wli4316MQDjTRoeH22VkfaO/Qdsu04FvD9dYZJnuNb1BNRmJkStZ2Hj
k6LA8R0BYGJpMeRtZvBjtAp1zjF4Bxf37yNJfhq9btpxI+5+MYGCgn6dkmBohnOJ
4j8AHziX3R/df3dTEFgoSeZG80WEUnPBE5nMjzBgIYeGVf+I2PjU2cgWf7NrbN4G
TK5Zo4pGuuWOmiiHsZqMrV4tZBEMdPDCvpN0LH5zRGYwBR/esrglwctkZrX35wY2
4X/+QOx1pAiP0Tg7LJCdMjdZ7GFUQPoIHedEBKOEGH/Dzeh0EqncWgty3VX8kbso
dtUq7FtsZvglMHaCR51HPhleVEd0bhDOeIb0K7iIivmy0ashaOAm1JCiitZ3ZQEa
9iTNRIc1lhfnyEZBm9A90LdfpbuHZ1WMpV4CqFPX/sxN1tJFFdCi/AF+cmPmUfZq
ZrhQCLSLncWvINsKOor69QWfw5XnEE5DH7TIE81a17tiwO6WDI+5bZLvv1OqkS8N
IP2llaf9ubMlmb3BUer7tf9V0TyRc5G7RjYteouORsLe7aatDl5n45mgTnxuCqnH
hvGVaaGUdLyBLpQuma9o+bkxkvgIF7a66wHFpWo2SY81YBL9eIiiznQHL8n51l9T
2mWSX6CkuxFhoatduOapXLLooKOaCwAQv/1mwwvJU5NvtuNomQljI4iXE+g/p7k0
1oOW4OWkd8yFxpXgDoZO56agdwf99toi9czreYFnpvQ0H24NkyqrN2Vsiqys+o8/
tBWcKGKJL4UuCqQi3EyyYBMfl/uSRh9x8WhYij57aEFgskm6hr1WKVkeIzPU6bqz
t8UNZVtlIDll1psh1/qaPcJCSb+RnCag//IRGDCYwPanUQ5eo5/iAymSkoPlB2rV
0LmHNZ2Nbuey2N5L3X0K+9arxmam+Q7pPk62QMARf0WATepz+hOd2AQwD3u7kpyc
wDNMVgW0vcKAKUDxr7wa9yuBrezazbA0tQRBwUMOo1MBPx45r64d4JSVZBQPIKY4
0vB27sK60B724nMlyakprpCCaB3F4MNDyVMnryTlZACsUdoWxSgbRB1aLA/BfJyu
drd3XUEVfJ5UwDc2e7UOcCNvs1UTJ/hNbuX2sGPiNunGoY0jxehqGKfCyobwHzup
HfixRzY2iwLg90hp3L6CW0qsja1Z6yV0b3ieCA17P5U6QUo4rVGceWl6x6LtI86Y
USaWkxcEQVwlYmnEvKUbnsMP+hDEk8hzmZmGmmtirXU0RhwDCqGI64ip1Cf9HtLW
CgkH2zOdjYAYIXoJ+FHG9fX60GmHo7MhFziz6xyc2QMJnhjnxF0ggNb149iRMBI+
ngIUV82UlaXpcjsmVYOvvG5cDyEmjdYcFO5cMRJRhWBY1lkvEy5r3ax8Pf1GWi/x
zZ7xkZazzLNPBZ9/ux6mX/qhn5D/0TQBhOUo9Q/ZbFqbyPfc+KCo36qlp/nnEBaS
ne2OCagI4xag93fF1XbUiBuG1XQ8chCxYIL7wO8bhn4d2PdR5tWijsfqGVK+7a7S
01e8zoFO4KTijuUXLpIZCz8gJz7jmtRgcNLEwcAwFwPwA8H4AuC7b/qU2kGbkpTc
ni7tpKKYpuAlvEG1cGZhhUDbcNY+vqtQflxrBShjmI6Lq8Or0k1Vi3pnZteNY9Lb
AUpoo6i5+dxfX9qGs6J/oUPIQTdiQa0ujngDibfKsNCaEPPbLt8SKW1ebXBY1c8m
uvDeOU881SVFrEaLvDb0SCRPzez8YmlhBerD5oLmI0dbzTwPlsXKCHFNoQEQuMlh
bqP6PYgnJaQM5U5s+kZGPecibUb/KOxcd8EgUSScaok4dGscIO2s9nYXVC/8XXTp
9pdgUZ+oB8rHFg+2zybZC7OnAtIjqCg7E4CXi7avzDpZDJp1uaSTLK4zSVaasiyF
i6zVHCXfUxXhK8TsN3KhOs93x4gx7fAbofn8V918g5+kX8OSEuAO/crjIeBW1tPt
URXyQmsBXFjvEIQ4vpzzy9HjV7QfYPi7Gs1NW3smrvRXWEymAALPlSHWZplztBvr
g0MrVrj53bou/o/7/KSMz9SfcDALcxcFYtya6CREnkvsaH+xT0+29+HjSnnST2l5
RzgPX9MrNnj1LPoJE25hLphV8AO64/DJvmP8hasJS7G+sSwqGMMSpv2qxKZSE0VX
tYYDuyw4JY9817Ny8WV41tEMSsZb14EahyDHqM0KKohqdvqXics24yaGquAfLetH
Tg1y1vpi3crKjc0gMW2lRtc4YMTJ9zX/HHjC/tZJG2K89OIFF2Rq06E5guutbcRn
nTEUPlAqqOvpX7CR/m5VgDZ5ERoMcO5cM2R0AX89gXAjkjClxX/2oucW0o0/Xu0G
VcmeWN/nmsujiG5MHoOQt1j+x3YMvQaBH4MjtMumVE0Bw9+gdwOndOeNhGaOwz/J
hRqknSGb2gT7wrn4XjvdlyhHhGdtSRQzyIoWOoumyV8EVwhymlv1/STRKZa30755
NEp2dpY/ZeOJIsQGPdgbkkLQh44kFXSIYo2/7QOR+Cdv4QMMiWfdq5IXDdkQMkWV
8ekDOpBJkpQip14EJlszSYZlkQ51sP1u4qBIP934CcFygG2BOVnIdNcW0LzIDFxc
Q1nDXEDb8N6UCHpWsYsGsEybkZVeA3ZESl6rcL6lRj2jXCRrfltDvo03l46AJGrM
MiOalHx72iejVeegkEmaxA9wL9NM3Hq2ypvg0lyuYxKbzDBz50QpHv6IgIukxfoT
vZVJlAJFzLmE7V3GTNbiRDcnH/tO8jMkTLazI8VuzIHp+6I3eYkdf/7JZaqZe7MZ
LqsMx+EuWmV1U0M1VEiDVi0sCz8g5g9UglbwIKnvaj+kEVkiT4RhIIErOpnXBjpB
Aus1ZcWrMIDs+sErax7Dwv3fmWmf4BnB2yX1nd/f/qQZCyCM0RIceMoyrxhghaxu
dI2GwmkZwnTUdbUL8hiCvFshB69jKZTziGq5umiX6RRflqYbIaI4Vl2GYb8HWcrS
cgVBD9m54UANrhz2qMmv9zwRI36ZG+UJ9A/k/TGREBEC3NDU7KrcOr63w4ZvLB0L
VJ89rkiINp2QS1c6A9so2bz3wtWOO98w3/jFTgpdKK2xuFjTKe/F4YPdG5f1N+3f
8OUzECzuCXs8MpLO74HDDZO8hi1aYsoWmlU6Rlz4PsXUOb2URn4X2kikjLn4rqEF
pdnXzO5BuRNzfJF+V6IwHh8Xre84XAx5FuAh11Z0k9aE09bSP0U3ogDrZ2MUE/p/
BK6mP8+GCUdCAm6fy8bSEDlOpBHJ5gsqKN5Bl7wi53bpqBjVEqY/chAh7pdrVEqc
xMRAP9deJI+hKEnR2FiP6nJlG57h4BTbf4iIXRc3+UcR4aKO0vugL/aIApw09ieH
zFy5MJ9lkK4DqanbT3fW9y/jdgf5qSAuYM4ahyaV6km8PoeuKdzMcI9OCNBGtL7x
ghFm3fnAqj1njCFZFg2ga5c/N9iLTOLz92cB/SE4nut7CX8K43nA/94W+rl07Yu+
Gbzjo9+tVecsT8qQF6T7VG7pkeoQJ8VK6ubDxeCR5R/lETp9X3Et2419UcZjYtTK
Dr7qio1Gg50ErBPHwlb1cNbnvs6ClVlhlI/vjbYzVYD2ZC0UWLlxDSPRyezgWytC
97TkFDyMXDBW9V/rEpi4DrPphQp9zMUAZxt6iDMI2coYCFW9NdzCU7gr4MZ8qW3g
dmXO+h2UldK/eUEzb9ZD8e9cPj6M7ncReoMraN8b+Y3tHL9QR+1CKRucG2ktXy6I
eLKb5OxmXfTL4VBtCcViMRmj+EVr2sVW+E+LpKZrxY3klGHQpFawau+y1OzjoyH7
dezw3Y1GrHJU1fmBSQ0qBDJFoC9lmgLvl9iKwN99qYMzgcQlreWmhkiNpD09F03r
85FNTmQLwtRMvX6VfTMD2iLQM9uVJsM2xFnmj0R3951A8ZJtYIpd4dl24q3CDqHe
mcg4H3e8iSMc6fmby54niLmzHlsLrvbcCQzAq7E2ONccYCysY3M9SPTGAf2teh2F
HFGVDm9Sa7tjasBrbsHxUlIlfTxzvNmaZJJyXm2TR0xjZSgF0CJ+t9KlmMgg26zS
gQpddkLcQHsXvH3acFZcmFJBNBfhF30OYNk4SLCXkm/3MMi0zrHCj0iP9jjKceAo
3Y7MxJgFOw9CgtiYyAKjjI5ASORP1nKhhZMTneeXwQ33uE0yvtifYNXJPun+0Pcu
vWiNG0tGWjRZTNXrmvrbhtFvEmdFyQBWmtOMGgGkKX+A8nk/bRumhSQY60DhCqzV
7KXqkM7yJGrSlN+Kb2xMQuSZkVuXRF5hqIYjRmk7v9sncntEY2McJMqJcLgdORB8
ZjA+lJLAN3P0BrwfHpEUtsoBT32pn/ceRwPUxrUrfOb/ZUXPGS+UanERh9Z+qJJp
Po6y+s2FFkFpXHic/J+6bz0gpHUUm/S8ADdBsbM205Yhp7ebkLkuQmILnfI0CL0/
A2hZth5oxfdctm6c3QLUruWnT/+TgkV2MT9MZjLrZmXFkkP0+mSOVA48G7TSNSXT
aKReRtrHRBr4hDvh3KTeq8XUFA5+ZpiipQWRkcWjHuXt5f6/bYvu5laxY9ta3N9l
6/jKxijLTinKpvTLUFKMbW9054AJ6Pyytm2qWbFY50RbJXleyxO23Jnviz8zMhSt
iw+HLL4GyenRw3oM2z2aYyqW8f81qL0/1fTWC1MOzzDtLKX+QVBavJJ3DFLIzuBg
EG6irJiyqCNxa89up3H2RVoZo58D/S0z+nE2YxXbO+V6aMPKMb8pQa2DDqNSl8ys
Xtre+GKKpH9MKT6EqE4yNM+b5YhzRwc4k9MSQRfW/FaU6Ua6QHmw15RBoR2vxxvL
9tRzlyPuFNjN3dqGjPPbzFqx9zrDWYXnews1Gyw1CVq2GtytaLMUWlW4fyW8sKn/
/CJnmol3ydPyaawrUh/vBV+/kEPvkjjwiz4T21I3hwg+QxDiHQlBc7IOqellNiu1
kd8WFUg1E4lTMVhSgleLcp5djybN4/FnS1/EBEG/TCc4rzyQFTtkRRARdSipq/tB
FYuSkQ9QysYAw/QOfmV5ftm7uTs4xlA3GmwZRnNOgw1R9r5hNurBbxyrMcc0SEyF
D23VVU2TIyOzaFo5Q/lsLLJDmbGKAyhsJ0IO3sSUaBZC9ojqFIwSAn64eW4krfgx
jbzKhGOVfHQcQuk8wyECp6w+Nn1srwubL1v0DcsGKHAHWpx3gKpnc6CncXt1WX1a
RLb7kmUwWaK5KZgqZi/xuHCvjkm776jagB26K7Ng2br4ztdpfgT2uJQSPNYN4QNB
V9hxODBFUgCmUOynhVpcHs6jVGdZPj73C8XGq5bFc/uEDkx1FedTT8y57FRk4tx4
THxK4UwAKmvrlikyuMEEEX9hWSdiNpv0YQbKA7LKP/xOeLo7AxxjDFOxdqLV2UKK
RT8qcakGSupG6OZSippfOqt2x1TEEfpwOT09Y0yVOp49Jfa8WfbMzunpoDJgEHvp
5qB2SJujT/QdXrk/MEoIvDN+vgUuF0NT8CDu2/7sIObeOufjkoQoG8um7KPmbkrC
huHTRqrDJIrz6wOi7jOCNdmneBfqH0rf7dJc/q1nBcerSgWnUJuHMZ/6VUKF1f6X
zMzmbJi7Dn4a7uklxocqz/WBBOoFsrG2kxjHHQjl2gXbPsmlysBCrhqYxtCOw9kk
vV5J8U8m4pvZt4RS0ZFU0+qi6PzUa+1BtYQMhtEFjs4qPbFyi/oQejP49YjORSO2
YejSQVp8rWRzw1XqsNlYL8LiAw536Ydl+EnddsGf//gKq0qJY7NbVxYiQzAJJ8+6
tBHZcoSax1oJWjHEWx7L0Og2CCl3P1VXAV/1w8jX35oTVLCWuztXERH6yF6JuzM7
xXK+B0P++HVCD5UexuGTfMc0r6CxwBGO8ZthF9Wt2E2g35VvGxJZvu+SBA9uw/Jh
NX+lHV11pv1dTCG8Svw1BzPVE4ulmkYKo3DzQBEe/2hvODuBFm+o6UfInwGCluir
yXoq/pk+CT6X+ZDUyh+qanSbS2q5PnXbazvQM6GhqMOsL/KE7gZL7fOWFC2fs65f
havJ4V9DpRlO/uvmRI1Zv4WwGocxV2HaGnBhpbI8fdoONwx0gBPTU7jBext7jplK
OeN6gBwyuOnd6EH84VJSUgtx0uX+oKKjGYRjMUXYAmPDhuCF1sRR6yyrkj/By9Xu
OA/smTPMzJxtuf01KZg/6PNVQ/IYLcaZEZYE7fuqPWQAlk9c+0lOzAufoeYpb8au
Bk99iLfPgoqBK4hYfmEcdz3c+qs+G6IRqrP9lfuFS4/LCg3KmYt7FB5GgCpgbqU7
5ymaUx43Uf8wShHV5W4qU5aCERhQ7HOuK4R+htJl38nMTwmZ09xjT3qcEfq/7h8N
pFl1e1me4r4v6gIocoUUkX8iujQ8sHNmX5PEjgY0xnNovq3Z8DUvFnp5iaepO8RF
a5hN77k7SGKjmD+tq5oIAW97NkilUx3o5r9s/Y10tNVNKgT29svzh1rNVeCvEuqr
K0WeycyFF9+iMUXgAjTSYLrIHrK+hufVLZaxBr1sTAu+4Ad2Hy4VRDDGcy6EghVA
dUei3xf5jBU563M1TuXD/ox3rh0uhGjiK+EeihF1PvbUwNpcK9xuzVz7fFL3zlKJ
ER8z2QtcM3947Mu6mmBaw4/kFfad6s8w7eDKS4T7RVOn1LVAb9PchEqx1o18554c
WneZMJA7GTWP82gAhFZKVpbKlOPi45KX+SDVZqJgz6/FrjL0usyi0rVHxsoU7biS
E1xaOeHNv3DeT3q/ax9TkcK+IdeMx9+dQbjI0tO4lQ0YBlSBGj/v/15JPX/mnAY0
PkMK48b/ccoDheZyo1JKj9gbWv9WbEWTuCZ0c/Mv/7ti5CQPH/HMnqbhJSa3yCue
04XJyxWv7CO/dCshJc5TZfDxhMgGZ007QapUf2wa+0lu8sOe2GipFh9t6IrVJqCv
Tj18Rp67LxFtmJeHrK6ZEt7sNopikG+34bkc6M3bjCttbq7+je5m4YFGZ1Rzfqat
XGZRSxO7ZvFMTL5PzGlM3yZoVN7K3tB4VcGiFD4bssTTys+fMHgHAqWW2hW5yo9L
+0htdcGi1UdRxYPTRkC0K5KLsz5jc3LEXz/PDPv1OliWO88BbBoyZvUY/Kv3DPTa
OI9/MnM6Fr8b5EZbus7rAn8rNNt5NzMcaVvQbsrEfpA3sOjP01+k05Ei/5xXcJ2R
cKh8T5luLtRIc3FKw7Evdv4+HONjczgQPTpqoi1xU44Q5pLI35arM0FChaWy2Axh
1Cyn0NInJgQRrC5Weq2JuhzBEpWbYqQTe3+zLRb1rXUAObkRl5zbSRdCEwgJ4mhi
HgB/4g8LcDRy3bMlb2Vkjev+2T3pyZCp6O8Y4eJzffNESjgkWNQ44n51138JeFn5
8URypqzUi1jDouxZHPBb6hJ+OPnnf2ryEqCH18qvoeXu5AZzjfKAEUqXMf3ocHyU
otEmrfEw5SLbmtX4GzVhr6mWdIwDzsRrxbBBwhzrepax+/EeFk6bJZKgd9IiqAj8
5a5S/51KXuUKmJy0Kox75PLFHpPg6Zcy84xm/5zzEjt1tuKOBHKQH9Sk8WKS6/NC
aNhltNSi/PX/esbt5A7C6kufuW+s10kBXEeZFltsuVu8vWoUCUYUEpVlpqrb6nxU
3NoqOmPxUGxCGUTIR9PxWWRXoZQmUu0StQwy7UDkIuLyaYVLGyWZqsynq+wAUHG5
EzZeuAjBsoUZFXrJU9pjnDC42K9RNNz/rJ47MoSPSCm9BPMWPwx1W/vp7O+BVd7j
NI2bP2SwZocposOM5uOO970Q3boyIvrygjUyeZCIZ4rgiHALgO7ejXnKZjuv9T9K
GiKEmXNNTV7X+w3GpxQnCe5LkFe2kQiZAN0hV3Jggwu0ta+ooLPid2IYmSgwAchs
AwGlneFUDuHOiqBQZ4KgrfuhPVL3d1qKM3aGQxE8S8edswZr+ZiZri8WKVt37Km+
6i0IsK8GyPKA/4QBYccH85VkGwQVCsuF+NQMUMDPqrO285YBwE+HQ61uI+rEfLj4
USxJQoGpQgpD167WdwwqI+J0WzswxQOQlbJuHIkJB1vAKolTB9pp4zti20nyeovp
D2I0zpGdPNIO2JEhAdZZ/YJ4R2s7V5FtYZ2Mk2dhNeoHhE+butG1x4BMgRFbIAA7
1Rr/K3jBJoxFY/rVhWtub3N+UHcSUfFRw+0uxD6d9BSOfpNDIlK27AzTCZOgSHho
SlrbwM/hnoCIOaHK1tWZhkznpJN/E6VRIW0QHgKnYZnDEjxaqJnTLl1QDPy3Hc7Y
dcKxgRkG5KV7U2LkSupsUYIJ6NtTk+fZXn+gVkVIHbDjEni0Ky3yavLON1NG3dPe
k+MJCJZ+H7Gvqb1ySjums0Ga1icfyzOn7Ybtrf6jHhawpoEJLvmGNYcdsAkKEmGR
CX8Z8/BsWUjZvXZPzS3oSs9nXFTfilqcE8Q3AdVf/sGtbn1VTWOHVrigxhoMs2Dm
MXZsVhrJ3V4XvUS/Omqzojpz6g+D6iIFNMvFZMdnyUNOxm2BhE/bEg0GLrz5MX3m
lbiItAL+fHj0pa1IhD0D5JMEMzobZdl/s3HowwLxkLjdUrHNKtBSYco1LL3uaa7v
qXhqFP9roQRhfXfw+NU7lI2tc/WyOTNRO1eZQWRcN59engA3sLuCIXMybmwLGXwR
TL6u3Vb7or7UIMq6//boPknEm4c1KsrluL1yaTUPFWZQB5B9jquqxIWfFvr+S2vb
f+tAQyzgCpoa7vB+5JXQDbrUxG0gULh0ZbSXpXAQOoq9liWjp4BI0IA3tbjWUhAY
0dKfhZC/4qhZZIcHL7+T14JghOEq5zpvmlY0WMafM1X+yil9FNH1r2NCEszoWmU0
EFkQE+TBW+KkQwSCA8zzt3SGz/ZMcsXN9GsZKmpUgBe1DXY6wjp+ihFsDaOCOG5R
uC6P2TUUc2LV2bKXIKKIkc6mpzEGvvZpbIuBXxWiHW2x1aF839PUAo43FV/C1HU4
WJavc2dwVppo8tTUsAyKkQP3ypIloGD/jyJHwZFWRm+PZRCX49BshB4o2tYhtAl8
9g54sElIJk00N8icbgVMQttuzb2OItg/M9bJVRCSlrUjIQx8a3wrl4QAZa3UX23/
xQf2jOi25vuP2AUpcvQKhXN89bDY+cCoLtuOrNfHM7KQ6oxzYfWeY16URF40TrLV
eMwFIB74HtmgfHIXPYBLYNPj3u7sCHQqBcElIaLv5qOXiU9JNwN49n609zm4R+y6
hWv1vUxAHDPLquF5ixzS82wKeK25qbKN4UFmnMrrHCAkeIraSV/61ba3C1QdOaHd
YhuR2hjLPpihSZImzYkQU6tAu+w6F3NicSqokBITqwSLRuckou1UenIKBqX3uQ4t
Aszv+jnxBvI2UBjPN5nIYvW1GUqbpqJU1UTMzACE0eBT00/R3VkLYedttsGAJOrd
C33XWHTZUSvO3WlwKJe7LbdfpvSSGa7WUJQ77+wu2HzzddpuZ2gW8o8j9sKPVNwz
LtkyEgBvOReN8CuxX/wSNynzvmohmeHRRvF38dOib77MDyWENaB4BSRn+lF/PYeT
VfyoybV2RIBOicLr5hax29XbJdMLPFbHvd6m1ov6WI5SxMBxloaOruyl0/1z2SnP
BEsRuRfOw+c/ODG8KClSdKVi24qil0EQSYPoA4q9py1GAka+YfNrDrzsPn+c1dn0
bhEZA0+OOQ3g/BxMrHSOcCmfNz+pG4rcE6PA5sTqcOj6i1Ayq/hDmGlE4kZojY1G
QZzuqyIUJmOIL90OI+8oR7H3HuGblULvnz3gJorCkdEOZGUCUUEjKWb3EvHb7KM9
nbrc77kWXLBCgJiZjqAjEIb0+UUzi2XN7j5z2tzAT9KAanNoigXu0CmZgNxIxGdy
Z4WVE0va5Q/w5jXnAkLWKicOIrclRbveuK4RSzBoQrBlLim13eARt6MNGInsppEP
23+jQDyWZgYDSZXqMsiPq0k5TCpBvb7alBEzqHuuktsMpQI8fC8XfJc94xFc3/eX
Mor83Kg/afirK3PiqyMXHOnWTrdlSCTE8tDQK4444Z4K/zUa3OT1Kt5jmXUJCjNq
b64lxgCK4JMK+yOq6j1PSovBdd+dNzLzWilasYhU0zC3FNECFEbqaXnWfCEBVVRz
VQce7JD4HqSpA392u8leho/M66TAarBo4dfpn/peHWY5g1Zlq61IP155g2EnyEI8
iQLffndM0Fh193ih6y5UI3X4AekKNcNoFHJ5yEG46F5eJ1Ba9Z2ZfpQ562bEN6gN
H4y/mKMH3EfYiYBPklpMAczPJWBzWEViZv8r1geeWb8KbzSZ5p4rH6b5vsZa4/aQ
JUw4roS7SknOJL+/zCDa7S7aOk2rbLWbehtQR8moD1K34S+KSrHgDasgjkGLknHB
6rioA4j9UK7GwCeD9fyi6zlQbCbEa7ky0de9nOWQyfPlK9wo6eMWvGSaD++SCdhu
g/iYYczTBywVFsHSV4twgYBhYU1/RYDYh3/V2pPV+kRUEzpPD/yFoDWwFejHbDAP
IDJNVd+Vtn9DKS1LzoXNd3C2ZWgdsQTiwI9TUG5MDPVCSAcfPNYPgyrcAhEIdBf4
wAWz/JWDUa6Ushm0bfwyI4GV+c4QXCnyWPMO/p1NZV77gXKV5lNKEGGhgHdAZLej
+Zfz9OkbWLKU/lsTaBfeFkOcqsTf3cHWT+XUnI5cKtXZ0bml8MMVq1h//uTgBOWL
kJIx7/8qNnIXKEXN7hW6Di+5NC0eNcAGOyS93tPSg0IV6CdG1xsWXgzPWKG5Y8PJ
gIEHcsn08qY4YI/EjKwnNTzzI65WKnjJpYx05eB7UHsibNp5vmJvgxBjqyLYf1mQ
wHQCjQNPPsgMOsWxYBLKvkymNu+uk9FDf8vZZC5vw5bjtGKzOJIqrgXkQMHl53X2
8VYr39vB8OcBhTsrL/HiTIOMtgXUSDy4s0Ui66Xbv7+qS1K/E6gqfUZTf9cJ/dgU
0GTtF1yM24pJ/NAeQ0g4HYEfy5rTKf5eyRaYPDR9BfQrGesq7IhmaMUhlXXOSlsp
Mji6aRfaPyRkST3tYxcFaIBhA32uZ4GS2yNGIF9+58tsJZ+9T6mv26Uh7RYfxFRz
MmtWuX8wEqvKZnsavmw9f/gUelUhz/dk9x4Djz96Rzx+dn3v+AxPeJikY+RuFA3s
VBFtpcjvRuG94oGcyGdvi9vXSPg5OGsIChZwuscWaVpcakLY6zETjskVOjf0Qy5e
r+dEfqyGQqxVunN5Tmu0x/tadQtbvlNbJiYbi6Ab4m881RpndMXjrjmyvX3JIcq3
Oqf0uHqhwp7YTy08/UeiDDSjsKUxD8216tkAQW2FFk4mb5g2kjzFH7cAj0ghX+td
QkBgRcfSE5crt4AdbuC8LFz98mEKcLCSWuNF/wn70wFWNbzkA0/pR4WQZQABHv1l
C7BgsXgzghG13vvp0nBzU9/R6kF00PSREf9Gi4XT53ysofKhX1No8k9DVWyf01aJ
uy1H+8D5GQMjKUncwJLGhHjg3OXSwL3tfdEL+6Xh2lZ97bC0dt2WYVqE5krAJs79
cUW0C9IWxkX3k3XUL3K7Vhz1ZIiE+2ZC/TZLhT+26lY95U41x0cDS8YDWopv/DoA
PXiOitjeoeeS6iBAAMtpjTq73c7YYnMnpizyj5PaXF+gpO0iD4GCctG64nbuIafb
Ory2Ta7rLdOpGLKeDoxbLTnFsYwtpKdvfa6rMVFcfjKiLo5QLdGNGiTnrrAhpX44
NhA4aenZzB3pu2qFYw+NP8aGlOssaP7WKuU4pUSkpHS1ot3HWXm+dDqkS0QDOGOD
z8IIBKqfgPYC373bzYL1mwuDCWPC91T6bUKgbsFjN3BCWbTMVoSebItulIRMTbao
sDMhU8HvFj9DYP7gCRv/dlBMPHgCSJsa3vr64j330MUfG03eozOMOsK6sL/06sZS
9dym1V4RhwV8Er95XcIN1ovSqPN5uM4J4dUw50G6Q9MW1bm2tP4USYWLtFCQ3EZ7
MErfPsdYolTIrpoxF+Iizh2p1EI5jCblqdxxf16ItsVsAxkv9zVpIQj/+UCcRL9d
ZEQd19F5lsmfpfEK8Wu4fk43K0Ar+bbz5EzoTpl40L87iqclzoRxmLjVqknPVYgN
PEuUe8/dfzAk4kvpHl6p4YbNyHPOyVRHkwCjpdRXZmFyhB2QPsUZpeRAn6n45aGR
xWNx5YTHrWeXMYJXISblkUrDtm22gKXimCtIKwARxHv48dPKgiED/+QNYkHxwPWg
8PbleJNSqX2vnQ149yUK34VlGZnazHQcRYWYtiF7GIiagwliGOhwQKC9Dp63wH04
RsWHrk9hArmbs0CPOt9syLnOOK7izZ02LVEOtyojABee+eoBz81VhzZ5ijNkElkR
6DJqNV7dV+21PLS/mcPifS8usOze1fmVLk0WuRHGQRUEF8/WaKfo2rK6J80mZEQ6
wV4qKhZAtJVaDcaHALoS/0ZA0tRpydpAkz94woPuELGtjhLJK0u+ncCpK3abOf1z
B9aI2+LsAGkiNnAHLdHSVdtTJEA3sxiHZils9eX29HiW6LoS6XYf4KQjx9riFwny
t10OjvmOia3wCz0LxzWGp884TOt4OwPsNCnBJKloA3g3ry8PxNuCtKH2SnkhBk7O
QSBFD6U3b0jqGbB7g34y2QII2fGcVYNfQ3/28jwP/LthcbAB4ESl/z5pF1+6Yczg
fav/NRPsgWRpdzFc7aRCgyV6IlxYcIwJ6bx1hpe1T4VevC0gGiSb1R3SwRDvVEvf
PjY9gA/NBugLe9E0ywcOSq2pf8qDfwS+ZMtl7wdw/krvMEchoeyaxB0CXuvVjU+I
z+XVcLgUsDEB6k49O+m7l8yVm+FRqDnUe//3A8ONTpMO2muLfEPT6BD9IgC0cfcW
9+qCrWtRC21jrJ9bg3GPzRJD498hCMjInlnOUKXCjrAXVmGOS9ZFm6/8rgqI/Jhc
F8/oi0cjMMkgLvtTr/D7Fy9m70h1JlSmz3lwDvMB9uBmuRmIPSwKSuoZ+F6XXVIR
nelUMh4CpT7gxLigkf6twitUQzoYhTs9EvwPsaPaE0GQh5h7U2UGp5lJ9894ep1d
p/xP29QrbB5xz9IKR3J9r2Zv7vKN2BKs8358WyOtsfb21ynmAgBZ6UHukDvel+Vo
LEUgstiLM2ZhPuDvC+pR2Ex6Y/gi63h4/JmJ53yfPDVV1zqzDkOmN6s88Q9PUnYO
WM1mphmew/cSy4QY6XP4OTzHi/tq7rJkWDQUgdMZj62BqOKbzOPwTsqufftGGE/p
+D3IzgHSOVBnje0W5YcLd56i4cU4KStdm2cv43JS39XC3rEDNoH8zOaUfu7CbV6z
qkfzX9lYmctET4V6kzFleRIsqAgVAegne2pV/6O6E3k+nkqoVT8svK0GVMYt/z1k
ncXM6TWjtspEMVzofRmpghrt8HgMcFdBfkVwBJ4bnh7IVJ3gKseScLmPFX4Tbwbg
Ru8sJyfpwLI8JghPvvNCFycbw4GmKL3WpCYTPaPQabGBPLB/wnKEkDaV+530ty8P
JcuzeXWe2cPXSQvnUvkprus/xslbwUPbVmkiFkteCAYD/5xXr9bDJyPYVQb800yJ
av3Cga2jhNg8VIgvTvsLVhCVg2RA3BFPwEcwrrmbKcrxaHIBD3pOOsmBvwMkft18
TDqoDfy5Z1cvMTUanUAwKgdj2odrZbDHOUicRexK4dhoIK4zFTCwT/RYXOnZ2nw7
sUyvFoUQlXg6cKFHE3QiTB0/63URuPcA9fnSzPn9FK2ejkp+II08ZYB7b3dFmJqL
HBJHXwbMC3jj57QM+z1+5P6jlAkQo0Uw1h09cK24dsP8+rEFqe6J7RClosRhj50l
qInvS/jlG+HpwlaQQ8/vsi9UqSeyK6RrJ0lgyAeqcjVfr0MMX8RTNBkLfTA3pxSd
zoO2dA0+sXjzWd5Xd1BhyyFAC8UhaOq1UF++O2rMvqJJn7H/hFkxulR8p4INlwzQ
Z+GmvUAqSVnz5ut9JB/dKrWevy1jtxJawbYUJDUCt7Xg+dgjl/mmx0wgVd8mz9U5
xq2iohh3KmRHx4892Zezq+x2Hv+ouOealdNKl/rEtUND/1CeqtN65cUVBM0BgAxO
mK7jH3qycgS2L70QkgkS+23gIvp8C6u0BnxNdCeU2iP47l5Mud+ckS9iEfd+VM+w
tWYUI1trPlh0tF702D483OfbzVs7y7biu/tPCHrmCnw6YKknquwsMSnwbDBmKa0Q
VBvwq0xI0gOPbuyhHEiPOKUsNas4HE+IiG5AxK1kMuqfMljPyYoZfNtKdGbKm+An
ahgNHWlUi2jJ3+Iy5u4jQY5OuQk88nF2OoEwzhbUETCvo4/B47BMMKDvCQ0qnC7v
SBfDfUD8fgGyuVl1SwF2xTXfzwpnrT43A8xLaHvxpSYKFBJubCOgFhiFY5rKBkuy
Ff/Ix/pc4oFNal+NHr29PkYJc+RQSkVzqIPLq0XdqO8X8XHx0Wzw5EzG5YgAqdsw
UkmbU+PTqX0JYArBTw9CI4P2xHyLNgRonQiX1+o0g6I6nBTYNL0uveKM0zS8R1/z
qOMd3HPrksLFJ9lmmuh2fLVJ2QcXq2poaf9t6H9Zko6Mr6z76UcjsFrro1sq+InY
+vxUnNvXSXYdanEOfEL9lRjbrD4YU9ZDx3InQo00F17VZvIaF0yP8j5rgUmQILBh
pv/iZqfEV9ddhva+WegLQ+VS8Mt2WJeEIS3Ak/zqjPSjmithaAfZVagCuEm9+ExH
pG3Yd8JJnSJdDsXMzKAf3dJDARUPU06YJH/nPBxLUoXYK0ivz8wD4uA1gi0Ahqp4
yH8kmCQKhvGnDqMtrKmtNHUxLdZe/dvqbeEG5530qcnr99kHh6uyS8HmH3jxwSM9
xrLTXrW8IxinAhULJr4cVkz4FdhM6u8S70BABhOvsrYUaxXUYrGi/E8wCGzS92YT
UZ/ny4IntcxserLFxH0hnxu/gZ0DIPbBI9SyP6NMrE9Rh7kzsKOp1WxHdfcu7tzP
KTQ33Qo8Dx2UvaLPER8ecqSuxV+4u/DdsmOKEGHjzwKInCYJH6uPbwzNsMl1Btne
W2TJWhvkX3EvqC+cQsBvmgropvF38uY2JyeDVR4wppgLkva+KvbLfay3Cv8o9xs3
hTlkP9SPB1y+Dyj55/K3jUoO57O8obOCudQKn4S58i/IL5KzcugnTJsI1L3nQdFc
JvVSGTI3oCkBjrGcjqcgyTRuCryjr0t0ZMwJk+RxepV6WMCwDddYJcUl9qvMCVG5
x12dapzmkID0GqAyDkd6yb6M2cfKtJsbmlh7nDVXZC0llDvMhwL1+xtZK0WWDA5Q
ZN97Yy0asgKyYq/BC25qerUoFMWmxkrRnmenMtVY31rPUa0dSUI9xTedyYQw7/3M
Ch9pGzv3UEc/cUOTbxX4KfNqqHDaqI7gua9yT2MvVcjulZ1dT/ek30z0J9A7gfiR
ieDAq/rka3QjRJozcVe2i3dPYeIioJAM1Z4+8P/6kjHtIL+7C8RpYWjBu+VEmL0G
ST5yQNfbdpOwdbqLIN1SDvTH9mO2UWgU+Ebz8Dn/5vnKrZbppb+pzBNtmewSiwxL
e6pqMMrYDde+u9tRwyE1CcvNUEF42b2hbvFQyLGQSmaNtDxINQJ8F9MOTBjFl42b
ofDs70+eixCdKHmP1REJC+z/vvAUuBYH5hx60DsLngq6OefDCyWxw8bFBG+SYaY+
uUxT/LutLa8EzZ/yF9aqry7r72XuBcWtzWIsbtgLXEFQ0JlAWyIyEsuIZBpC0C/n
QpZklsAHYiRz1uPzZfA4nR7m7qisPKHqzs0rzWmLTFxdRnLmzTOtqdlKoEly63yH
CaHkrp00nWKMNMxX5kYGrw58ShDuyvPbY0BW2f/lyexLvQ/nNnEC7wmpDwUNpCPT
V2YrR3MTYfijC7qpmjA6HHJ4VhvHbIXg9JxRh64fVYRY9QJWmgkKnAEOFi9ri83C
T8fXgSLZCTG7qt2QVvPSnlwIBWuBSuLD9slGKdtDC0yOf0n09gx8N0E74xUm5t2F
cz8NWbvFEWSs3sZlZNLfVWjjRfUU/Dn+33jjN8RrKvg2j3VfHqpsQPI5QKP/LSun
p5zEAiZBeGp5IrKZi8iV7YN+VcApVLpWI5K21WKc4cc1eFpSkunxcdN6n9oijoZu
JdVKK3TJglhS8p0lZWDr34wc9cZa3gSPhYkzyQc+PXWLfbbMaZiW6yQmYaqyK/ip
E+TOBGbuIRpbR4RMalPRIcMEACwpV4oGdRG41/Ul4crX459zXljWgT55U2sQUfJX
ejUoz5EZ+JZ1/DYnDT56TMcESW14YYF3CaMz2PXdfhVm+JsRGWsQQmSqivZHR/DZ
rJIh3Pk8bzvfOfcDX/UgC1qo6vydUTpY8nYsRY7ZpjgIRYBpXo9th9QxX2KpRFSg
o4IV+NnWddbPZ26BW+9Iq7nlfYBVu2oeZgxA9fAnR0OUrK9fu+TBxJWlekLE1ggl
u53jbXygfMzKZKL4hegoIUdN0UJPVm6poRoOMJUHjl62Rj5A4STwekEkTrjgsib2
ellb6QxxhsRtlnf4X34pqJsXhJqj4y1kDPNtgs+9R8qXscTNwXkBEvZVimAbgbre
k9lGGt5DuPmI7UGKfx4bv2pcRzz8onovkDeLo55ks/4Nw27wN4MSNGWzC6mhR5CY
Ty7um5FjgA8x0hKdte3hut6s+h+7pD/zMyvhY4O4EYbnFQBotUPLULe/jPzO85oN
/9DiQg7alL25fqtprjQ9lNIacI/4pGqTRzx3lklmj0JJZ5qmfCRj+BgVnViz5o3T
56g6xsllTh7vZ3kkS3EC1ihk2zzGGMgLemm9Qkf8tGKgKqiaNA1VHrgYw2jZzJb7
iYTg5frza30K0xCTIc7xxsgTcXRIm5qSJpeWfMwKniWNp2wm+YN4lnLQeEIFltyp
tzC9ljDmPvtnyF1fsDMSjm1CusMkHuu9b4+tiPuyz/WtgTFqeKskf4REPWQQyqfA
bzYeQtsUQ30Pxzyel5xBZ01dORMRUpjFXT7WZ/9RXhJpGsnnRFM3Eb7DT/pEbL14
R+qjD0OBdI92rWA0sF4xNmonUOKJpczyAfXu43wVouwrNEEwgb5iUZJKMd9j0TQJ
mjXyhY02rpaxfQic932+2fEnYkPGNLyhKqTmvuKRJrVbiODZzhINzqoXz+W3jkio
BncvUmcsAadpEODjFsGXeUZFQi8uEBCM7hJpAj6IjSLvkUXl3r8OwuY9uYnPwSfR
NsZZkzM8BfySr1LwSRhLF0dALH4Dt9lZ9o4ld4rKxgLvBjZA/l+KMuONhPI1Qkie
gqa5XvKAlgIXi6aXzwQTOpXreSW9Q383FodKy8kmVc86eb0aYaabILuR/kmwdTh9
x8PPx/zJSAgYWjLst/sSwGfAujl8J5q5j9hdyh2d4nMuqGXWn8lSk2vv5HnvGstJ
3RUtu7rhILC0DhFbP8gLL9GEzut0P1uvoy1K1+dl/rzVqEZgIWMpdcxveuf1f76I
c3HbzH5htAKk7aiP+FfKz2326+ifPsj5ybYBVG1T2agASzQdXcoxc82n9RfPnRmz
BPwC+f4wUkhlnaq+GZ3K52PpGGX14j6GkgQYyYjLSZdDbQYCv5nZtoVKsIB8lmMA
SOsW5zl40/cKJ5tArI/LdjQVe4ayr5+Ibon7qcONGhBupujqxL3RIHTQyYUxPH4B
hmITVhCxJDQtr4hXQOSIrenY790v/bFeXm0H6QCq0N8m8jhdtNXnDR4ZslIKluNf
QX42x9pZfGpFjwdKbiLwbM5v5429fz4LNVuNNayUvtXJ9OVpGJWlk2btfWMuX+Vn
S+AmBeNMF3kLK2i8GvrjFkl5dBqjmGaMT6Nkpi9B6UvihlPPp1lcorTgcPGhVu2B
4AWXnnWeGI+jjk3q5d3va3p+8xn/pkGLdfMwTVK79YnSV/aAHu8iAKJ6N+GWaGKQ
z0M/oj44MBEbHs7flkGUe6yT7EtGZMwACQglsxpcIa3P3OEyLiXyvD5gDikWp8ZF
faFuZFTZz7yUXdM716K5Wk6wPiqP2j5Dm3sKDoPUuixjf7Q64OBRWafhLAlh+0zD
aDs5Zuaz5q8J/I6no7iXcgKdcivsNYo04gMx50GOhxknr4y+uUZL33MqbGCc3jTB
WCf0E3H3sohUn+vej24WO4kGS5DUnO42xQtbMI/MuGEd9pPxiVIENgC8NBvL7cXs
oPhKCeFbQ1cdwFvxZSm3bpferYLfS2TZ7Yd/k7LM0KXfYLNFyUNPuN+xvzEjJpmr
Vsw5+Ey6Z2jewOlVOBCaDJmPDX6+OZkcRtaPLRctd5upZXW+uM/gU1WRocjDyQqF
2Zssa8Zi30ta0AMibpQIVjv0w36J34N8fTdwjjxqyuUscobHjBuOTQ9bNYC2zpLV
xv6yLPqi7UEGv48osNAjE29aVGPbOdyMeCk2DPmiHkx9zSdtmE9Xc3BA1F1m0Rp0
L/3+bKlxSSIYOI3MXdQNC42ok1MLSDeQhn/9GlXse8hbJegtbC9OxqTbY6t7Ne6g
sbN65hpEvu5CkISQwGqtJy4YRAO64DOoMkOffIrmvohl4JO57SeuMhX0H3/x+6xE
qqEVHQBogX4LGNopPUjL1iE74+eyXTjLZroZfSiU4M1scY9ArNzeVuGCjcIFJvbX
nhfc6q62xTu/zolGpIhXyLwgcgUjsHjKmd34IL4z/IVNht/ogciz4oTmFIt5AezA
cirDac7oQxjz3oZyZXuzj6UG+Eu81VXM9pDB0xL/0p6+qk23NhzmhmH6AYYH1/bi
tXdJ7EMevlaJTFFJGVU9jB2RdDHUC1qu8fIpLYT9KWwkCao9Fi0riwPBvSrIAuAJ
lasY19/uhm2DIPKz3Iku1u0zO8MkrxT++lurKpJ6u9WS90xDsumTOJnWb2H66kn9
MQgAclucApI0TaCkyMqMsx6GgVWz4okoY+MLHdezyzICXUvRqThSrIwwQQDnwhoz
X0/X9wBME8ggASZ5ono32Cf4bJs+9B4+1/pqlNIee5sf3tN8M6Qw0pgFvB1YZAB6
wWg85qRZlVEQYKQDeRmX29bvgY/LuvDi37V7a5qz0Bpi8fzJYfgLnkN3gc9jZ061
HNA2+vIxPr6f4IQj+P5jfxVwUZmsZLzSazouIAsum5m/pVm1SvNgXKMCRdOg69hZ
bDWT6pLBzCSBaUxhtYUwtrlh7B/TlJJVrlKMWlpfoeC/UlPAel+fU/geoL8saPqq
ob37zT5yetYPheYqdYMh/qHrWQEGsumAxFdvqtxVlLP4y2n+57h6WMVu/Ty8kCdd
6YYCb3oKAI92IjEDXd+ttCQWaqVyfLuqsZsalJK+P9661AjJLhA3LYPTit/TkeRC
PGWYx7z2jPLmVDstGrY6Kv90Sr5isC0tmhBB+NjQe/f6gRcmhfM38nxrhU2tITi6
FqybxDaeO8D8QWaKA/W8KP5tNrkeCAV3NB/BKj/7wbNeo96okuZj8hmtfu7+lChU
adjkWBZ94lf9Xi1wpMlYEHhUwYY5LFqGWxMnLq5U0amd3ahYbGh3WXyG2WSAcC7v
rn7QYwknciOv/oeIMfRDDsIvp9sR1QJ+01PJB59guCIRkHXkjLK2LsUmmVDD2clr
3GQbbnqAEsMWdmFSehKMc9+CWum/5bRdyFVX/IdECHH7eVdmqdQHO0qVUkTuvDUQ
7Gz8SETsjcyjU7hKqLegLuT4Tpa7OJEroslBuhCM+pt/D62xTnBtg4Qdk/ROJ0I5
ajRVFweIHUu5ybI4jDZcjB/ExBx2blt0L25aM8fVWVO3ZQRsEN4rZcvLZSL2rD9+
6IyGc1g+DihK00As6m2PPqF9QvCXL+ygDSztZZr0LSLVi1iT0DAKSR1xKOCG+Jym
onW8EnjVw4YFjiJKFaSBzWGTeRKAHVU17m/fz1kYZ6D5fjIB5g3TDCLRcwLzM5mc
1ZaXZqJCqhvfRbzFLoxo9QKSLtndVGdR7zeOeiOmE1JbNtbG3xAIgA3zHcsH1k+/
ni09b01fZN9/E2bbvEe1sQsFKE/XpzmpvrsHFLXfRpuQII0nuW/d+peMvxgqzQvY
3UckGU5197dMliSSiFIuROiPnEwq/+fUtyjsSz/Gjjw2sJ6iygfBETSoYj3EnadC
Yn/6YRxQHDuVgypzCWoGqqzbeSM/ui5BUZPdmT36AfTw0QXaEGCOGQc3KkUknKM7
NZRCGBOGreh7wGWesHbnQW0enO7FSGNnjebHsj5L1Jjmep4O3fh5BJ5Kf7qrmxxu
l53d8gPtyU1gGekfJEnoqsSrdeXGzhTJgzC8DhI2bGv78kuTl7gi4stqiwXw8Wbt
y9UFi1BQ43asGoohvVF36mo52DmAIV23y80uY73NW0U7rS3B2KciAyAsU2EvIBTr
A4cY1+ETMDA0KbsZPOWbwu6n64kQyqN6kDXdaHVUowEbBBX3kirlSg+XEeiLWmO7
uN7t43lSQ/MvaXcMDUO/gUa/p/ki8V4+vvJl0aiK0G29h+lW9uQ2SGuABV5rrAY3
/Ca9nIFmdvzEqfHfmKmVXjTS7TAVvjhxNg5VQ7IZkqmxxhf/3SPpB4elzzlLRv4i
2MhK3co3yTlslcqNoICJfYbUk2YEO7QtmoPcMUAGjxx/6bIJcIUgxD7/+vI/E0WE
zrO83tWJBRPybkDxtfluT3873VFd1DgSUGBWkmM33oavXgTENm4B0IxT4wSFlwte
vPq71tWGit25eeMqzGpgBeeaiF+nVIDMPh+pr1Q1lPe1x4q8+sRfgYjYwlvVruFx
2JDQqMglQjo5sFTy8nyDQB2ohIC60VNmNuSoKHi/se03yzauTCISJGn79kZvkCmS
l5EseqOYHfCPEbbF6FVYczvAxUOUpCb7kK6vnh73ajFFNnT4yHI1L3q92R0xtgUJ
qOFGTBPkfR2dBghxWCZVPYtsmK63iwcHi6fNls3tuR1IBYXFLyDfdqIC2eBwGKNj
VzNZ/9bRmhyrLQIbLpi0De/0h3WnMqI2oclejiPZpK+Wi+CDmmDD4TTGXyWtpyQU
vs7Yv1OXXRphEvtBGNpWral6OGHDVvxxYDE/iW8BMOGWADLlq3otJWx0S5haO54A
Kt3C1b6YMK+l+UiAd9wgUJnFmDBo6v/cM1UDdUuDS83LkUusFeayksfyHmlJTl8M
7/wheKCr3cgsbMQYt+LIV6YCJkuO2Gx8cM/Bsnh517mBjvVUiRH+BPmfdxPKUYbO
W5QHp9X05MQs9LgWQSgsXCbYYJtsfmxFoK/6O3vszCVK3q2sagehOU8x7Fc8xTXg
M+xFK4BHCANY8dGLQVPHh73iHn+y+Vs8kVhQFt0pMjmTvnUsbituq37QCdiI6Q9m
bEy7eqayhRHucYHoUPhhcQHoMSwk5srs9M20QF8q0878TLHW16ayJmWUnMOO0O/D
T88X2E08DLgr65Qz5lR5RgiM0tBVBKGk/0uCpnVEAN6JX6OTZs6Ea+VJKpS2u8c8
DOCzeYeUb4UaHXXE3GEGzMoTb9nK/v1SRF6GvITW3uRrq6xjt5IsclLQt5WgQ77j
zTmFfh/flUC3H99zISsIvbwO1xWqOP4hp1UUTVL9JFOjuLT4L7xZVGyAbUQwl40s
Ad48RTZ1ZlqHh4tpFYXCASheKFtGs1zL5RpE5UxpCIiWkESg/u3c2QFb+wDdT0Y2
tPt2oC6ap/HTC9+pXARuvdvjBinZF8XrPYqI24dpcvol9pCJIfFy5aV0M1toDUls
Ys/oNPJYHHt6MU+1JBZlTxgfwsNQcYZD2ILfn7Y0Q75qbhAau53z/4VKQUKimIoz
fFTRj7Q0sUSl7+7IgfLAzbn1XDBfqIUzosUJ3Sm1p8Ahq38vFF7ZDvAuitmDXOKF
6m+l5Ri/nE597uf18pG98h81cNUYSx2FTZads6F067Ks9AiB7qYYhNW/QVullyfo
k0+OmDqSaGOstdLoyEQZ5PXPYzc9P6WyXlMQ+cvY6WIBw0CTkkxtNk0etc3TDrej
lZWLqiZWxdWKdoZjbuNeN7N7hBp8LbAzLwRctfiVDfrUg/3y7IJdEOnz3cN+cHqc
OwrXfQjYlnxfoHngu5+BAi4MjlAwjv822vbalQzGAWfdqwTNysplin8TFkli2jq0
tQJSKdmtZbTuxldDhZ9ROTk4cp+7QX0kTYSD3eGGF76oNeEzKaXcM9xpIqn+DPLG
aytcjIFqj+rBLreD8Yt5Jq9JOABothMAVABiYtSG7GBB0Vzr11BcO9zci3LAzwjS
Z/+VyTuM7UC8NXKjS2dKDq8w+IU/kLoJq2Ql1H+SPZuIlumeT4T5EQIzCvYQD8vq
VtmuBuVn/hD//uok/CKb5RtqwdZq8XcrOY6IcZ8Pc+fuD3lXBBWMMRNetmE4jNS9
6M/YMijCT2cQi11mJecqH7XCzMEwvacLMzeaL9CBeUFXyhosUSKqTGy2t4De/LOR
7rDMlUUQXFxbDtlGuqFSgQBjFTLCGLM9BeS/lA9nWQ6MOBdbYob+kOMnCkw+6VZA
RbOzvWToTex4Bg/DkKcStS6lM2HAWphqihXeOcEbE/1Tf2YT00dXaUmcoIkacQR4
y7e2y3AVbLVtf1n7QiPXRVCwS/cm5UGs0E3Avnd5Kz37m7lfZbAJsLkqFryfR+n3
0wVXTES8pG7DeCbpwIQSLMYo1uOdE5fmJ/kC1ZPs0SEFzPPKfnVzk9Y6WsPHqDWb
fdVc++g7MOEI/UJT75ZGW1gfrA2NmqYHGKgbuehTsDXSJvFL5M+KwrNb9o03mZoE
SOmKujoGHCfuUUZZ1n5hWI2ZjD26B7j+P/4uOfO7Bw7HRtvqm1tD9z6wDontGycL
mjOw7YrY4WRWZkASFmSeKz6gGlaCIy3nCLV+eqvmmSOBDw1P58FuuJR6CdOVLFQn
+/t60dBRsTfU0Ce9DxyDaUsUY/7Y3dDSG+qB5s7TtJo5p7I/JOaW1E+nHxtGaYuZ
mz1+FHFJW1nr+aoRiyL1sqtzEFfabKSV9zU8qD41RhdSf95bsHOkOY3eUTycunYr
WsxJ3y6unFIVAYhnnWpEUpjRl2AEAMPwPl13NmXhFk0BHEWVXwiIiOorUHexi8hh
YNCrzw7OUNeIaNo5wX999ttSE+vF1H/T4CvhEej3/hd6ZW0PGkefikDTUOJd6MO4
B4YgoN90AL2dH/l36YKMl8GZBB+dKqGD0Y/Mt92pMjV0apF/ujJY74ebLfpPt/8c
pOaPBinwsaaaV1YmxvkCxtxbepcg8V+89AyK9ApRywK05xqKByvuvEPtU1B0jBtD
ub+UbW1qjjffgrKD7mUxlbR+nSnkGtrq/NPld191fQjs0hWeFjfjoC9GgGoiZQrz
IWfBwrqlvnlpSFL6sufNTv/lPFIfP9h5OQytcUWNQW/wvm9gR3GFSZkVIUlt/Wcx
3iTXI4HUHZv04awKPYG2APxM626Y2paM4v4zGaz11UDbB3TrQBOA42uGyn7BJKQq
iFML1+56skvl0q+2NDOxp5nvMCDXmYkBOB+JcUMglPp5xWiSTMFvj4xy/5Y7dBaP
T2TSAloauDHBFOnqBZtnc6ITBb3Q5N4ggmxiNsWO6T06YGFTk+lYqGFBiLbY+ADw
b/11jNV80MatIfb3FFpD2hoRmYlNz6DhmYRumWosfz6BbeVyUJvpFbSQ+/Yyo+Pr
ERJrELdrAfnrGPZdokKBRl3v+hLieCjccj+F/IV/d5oNmYlAkDEw5Sh5azgtY9FH
2uNICh9wUEIWfJrDVc07IY8gbrJ5ovEUwlUq4VVLi0P1j7YZDVclyO/yjDy/pETU
r5CK2WaOYERUqoUgMAEAUf41/w2v/iRdD6VZDywxujc4ghm/0aE/842DzMF4BEuw
6qEaB3uZ7/DTfFOpDs2BwdPX56YnxEZzi3GCkynbgusPlPXXBSCxZIBE4gzUent/
q90WDoMmQxTIgFpuVS/kd0z6tEpAP4kXx4hyENhrSGlvoWAOKcAk5euiFP8hlXh0
K6w7hd8O09C2l8WLDT1RCb+mvljsSAN3MtbgN9/S9NydHr8AFf/149jx1F8FirO0
wk/d1BckwooMAhL56i0IYGbCH1nhgHn4d/wObfWSjFAJA6ZCUL52hf2T0qfhe3nr
t5dXtQD3jFNpXxkZvo9W44oLcxynubwr1fWsTby6B0MInD9OVVHOHu8KHjfS3ni5
W47GazB8C8y76vSA6IcRx65RiLtJMzSpXjVJ5l+CWjnSqufwB5+oQOGkXxgMVfqC
/aNwktZZoajKGpXREobxYRBT0e+/qv16Rx4eHz5wv3BP501HrQTIrcwxbtOlhMqo
A3gaRKAfTJgsoD70+VBJ4fOEM2dm7TT8oNIYl1+/mHsRS4VZ6kXyKBTsFIdO2Clg
E3Eg+oVt0MA8b4vUwnCcBUaQd9jaHaLAOeWsOTnb/IxDNEg0IlhN+ZG96AWNsQTh
Tr1UsM+x4qjqRc9nZbl2onOaOfkBQlREio7ym2ZU1Tc01WsUggMK6iJmWqYxSX4I
JN/02fKRKKlL5/qOQ2KG6wMz51B87Kh6ec+WSDl8Q0v644+YhVPtNWoXvdyjfKBq
hg1mQ1c98bGWFVC70PQ4yaWlLmWnX0ab1MYxJcuR6reaThpCNoDXuIBUxTDKJM9R
Ysymapt3WN0gh1M0d0FpI3izsyNGszn1Myw57qhDOduwz1RHYjcmd5MRV4hrtapo
S5ZMahenhof5NLTPLnxXRdaR4MvHHxjLdhPiATSO58Ttv4PemZ/Df4P8bMYaQwdC
vBNKhtIiXXRL1YBqL2vxmvqTHyzMfaMwRmgC5koOPFjLQG4/uQDQAis5RqSOtUPE
q9+fnKjAiCh3k0Yb5wYQr3iRCURzU1CFZ2NI+HsNcSaum6o2SZtP1ZAsR3ZvgUoy
aySO4dv6FpBBQ4XjbjYP+sEE+xNsKGfVf7pfxW/v59Z++SP7XI1b7dsF3ORD9thI
2SRl2cykpCeEsQCS5W/o8c0Xr+6ve/icZmcbkbG21cDmLKEpk9oS/4d7IpeLOA7I
fvx4nqov8DrWHGm6aH2+UXtvHp+KeEuxdynqNI4YcB8cPIfWJPReE5DgmU3ETSba
AHu/1G742UfzML2unXxaK4F2OF1CD416dV4m3XoYH3jIrEFSsuZYi7ugrvPB1Lhb
roJnZOJbvcH9iTYbjumHnAgKqMJGRW+FG4P/GQHVasg1Fglfs+AVJr0/aYhfhrbO
CKjp3MA9F/UW8ey44Ti3oYAtXCyHqJofFdpcGd4CNAy1ZZl+0jYgRFtFscLuSyzF
z97FFqbE0uHIUu0zOxZeQzEibDXmvb6BTnSQkL/31++NpWixMZqNFar6apAodp75
l99s6Pj8pIxKUZN6vgEP+MEntcWAqx8MR28pwnmGdp0eKPd/YIRmXpv/ntg/eQBC
cN9c/OfIzsD4Y3JQVM0IjhJhvzaiIO8A2p4o9FV3QuX8xd+E4qYBNQDkM5A8G3n9
TsadmxO+P9om1lCyBWiJzmjNlxc3XeazjTeyoDL98dMc7EqayuLTD9oA395CdvfH
qoSj9WrqLhlXG55Sb0X94aD0bwdt6KpAN4xkSPmDpDQ2VUHPSHJlwtR5QCmE+S43
hlkX+pl9oGG9fioTs3LBuzVtJoogipAxdJjvw6sqQT9IJQHTkTqoLXvRYQDgnjOw
VAUBhnaPoS+cFMW2/jeDRirwXJ6E9V9Jg4URjiSr4TOHi9LVObQ5yq6epl3GRPlu
LRljYkrGsyJum4uTwjFX3UYaR+7KQJvf7Y92zViZCMp1s6yb5o6jtSn0Zh9glsPy
enRjHjHRwq3/StvwdcnEJC7UxZKrJ2IX38Frg3WEtOVrtT5Um5r2au0yPJxrAV1A
QGCPKi5bQC30jwjcUEQcQfJWREBFR3s1P4db7bPCDncqgko0tNqZHmPZsIRqdeeg
H52XJ2XRNFzmx4ZNEV3E6c9IeMQcXV79eUqpfRM9f7a106pPurPtWm3H0Yte59xe
oHAiysgX8GkzWkxwIvDhCqU2blqytDyVxNV+nDoT4A9jFx2lKa8VHgi9M5luC8AS
gqCCFSvJfce3QpSt4Ey79eZkqeujBu6AUZvGwIKhrpbVSvODEih4naNzK13KlPrv
IZHqmHfEvIOpeK1v6mCWcT32Ovxb/iCRBJSV7YNn1vvT1DaU71wAJvZ8dMOB0be1
h84ZBMT7UraZ0t/TySeK60clnwMqYsEkYY8AH6TWX4oq+MBF0Mua8I0sjrEQelzJ
TWgLXIDvoUEaVufAjtyFDZSrWEp1gpJR4W7s7vHNBeHPNfSPPUudA7IYptddl9/J
1poPkr4islqDf0td6NiBq7z4XQoc+FjXzNdzp9muKuS6byQnnsroz2UaRtiLmjxo
XfVzPm3LCgX4hduRokYmPtlk+8dKi/FkgejEkEySDYch7m4eZx8btRCUxbVfqvgn
rViP2rqrDvM1TQPbUPOXZtwGL+Sev7tmQ4UBmQwj6KOZ7C915BUUEFFBwrzxe6F3
uN0+/YC0GHHAq4TgyGkwNF8a99oyww+FQSkClaJBcwqUL+OtdQbL5swy2LOQOgjP
xUtYe6WDYTTKEZhvHlaKi3co9Q3LuNdIiDOpUwzVw+mLI1PcRhQEudQTNE5e6bvi
W7MUf0OpUIuxkBhYOKz5Ent4H87NRZuN4hxNC8nMyPetr2bbJbjCLLEymleiF4gu
hLtm7wE/A03Z6liXRD0VAdC2PszOtNOAkg++mifilnCRQ46wCn8/dDERHG675WkO
h7rxkRnQojIfshpk45fYTHPh4cdwwLktDQbPyKshD/pxvgiW9I3rx339Ebcc0RJB
pfkC3qhwc/yI9sMRK9NkxzwkBEWX0iYeSN2V4YDJGAKfbM+rV3VP3tT/Zo0Zyotj
BNag31gHoCWb4VCmOOb/W1Op0P5UHuEWjtRmwyqL9QKIl0cqn5JFaX61ZsBVbJtn
nkVqrWG88m+/VMKjoJfr0mDpqxByoVdh6jVUzqUQlYofo7dSTdaGQqbkTgxMqGBn
2rcL1MyjkqZiAJcbTIcuL9+lpFIpuuN95IJid9sLYCFDrH7u05XTVto5XXM48BzH
R8AzjrL1KhwoI7Jnfe/u1twn/L76SJ85BqsVAXzTPyumGdMh1/Kotss8ly+sT/Ji
zAKUtnXe/RAs+BZXzTRrpIMGfILgmDgzlXX95oEtDiWYBiQ+WsbF+OP8w2UFG31V
Lhz9Fw0EU9mJh9LUSD32lzCO/Pu/RSeosOc6S4IUZG4E9oSeEFQp36H9Y9boZIYb
c4frBaE6sbiUaBVH+hwvK37uALEu1Yf78tBpRHUfba0QWqEPsq6qAPFISpusknJM
D6fYhvDYP2tdqcQgwRy5DAkks7nhXhbGE9DcENkLGjKLfxpTlI6B1yioZV4+FOV8
1vb9kfYAQgZ9sr7wUPNifIhgboTwO0p+BsllfoJSjsGrq4WYYeAcp9dcT+g3tWF7
wkmIqEOqS0ADrmP3xkyeomKCzyq0osLoaoh//uIcwwns6Ywbcz00NcY4gmXVeY24
syIH2cFdApaK1jknz5O0hlFc4ARqcg0Jo0qh1ORDFfAb0cs/5nO5aRZ2qV5c+iV/
dx3RFY/I8+jlFMC3guhRTtjt4+b4zBcSLDYezteqOUclC6ttS2Win0/lAditWe45
UtiTKxK7w/ku+IAC7Nl7LIo0Cj390oNdHrb76RYBz24TsW0UXovnlQAQGMSswlyO
vK9B9gIO5yezsLGbdZw1PBTnanCyPsrSa346GDqdjwotrxm+UFSqowqWT/UvV7Li
V7hGElwV5qOSRtbm8l8/2jm3ICRRcXemGTr/xSq2ckSNa/ZiP8jf+IiijA7MCH5h
1aD6wnurtb3Shv3lkNnwGoWEsdPfQj5XgsvwCgs/Daj7sODlvGpw8xssf/oe6Hz8
P1ULY30/5/RNVQlIwjXdnQHcw5+VRvdDshaHViN8kSCbsLrc0YQfV3R8Hxsg3rWC
nK+Ap8ZX46aTObdlZes2aLw2gL1DIxYT21lMieW4kxzTHYK8NmlmDB78LEMOu39c
fhIGAIHTb5LciwQrcRwTa24IByYiPVPsn8GXEUr5pLADNuiHiE6DJXlaZz1X0kjs
asxgM15uPcXiEAy6NACgPVHFLvKZXSMxQUOXjGb0CbYJW1gS0sm9KX/ivDqG4yOG
r6tUVJcHAskcaI9fWubQ9C9pCrHoXfIHLIVUpLZWxf0rHaDRO8yTL5pUN4FwtMph
hvSiQUaBa9RnRFiBXzLLFYs8a30CogADqTC7Bbh+/kSHI0yH+939SWfJjXMcI+WE
WDvjc6awNrLw90hwO+YyJ24R37f0E8J4QJTr+6y2baIyOlSyVPb/pP4aLplEfXge
yE2oHgA/cwpZ3DXH7ySrqDUBwojnso4GcRtzwTQP7xyh3LpKez1sOHav6lfR4UMz
t/RQQTZYZM+9rhnkp1YhROTNqpVqMmu12lxIAFLs1KgJhAy3Fac0vSEJOY2+H+T5
G+pcElrtDYnySFwY1KuEouRr/nuLguZsjwHxoMkmLDnc3aE4lvHEgn5GUVavGHSx
hyScho10c0qOLHCoDQWB43qJ+L8RG8xAVpM8fLn/ArXmIzkIOua3xekCYSC2XxpT
Wahi5Rx70MNSjh48umBNhIxP8XZ10PIg1j1czZJuSqkvhKFZYi2V7+mnfzmBAJqV
W4qwIaM2QJcjEc3tmGtEwQd+gnJpezYpvF1Dkdfu11oIJzImjzYqieostpG/ML49
A3WaCNOayDrkB03MHoPqxaHI9Zk68Cz09/YyWfF19a6MFv6Xzn9LltqrxzQiVoou
QJmVGGK1Ocxg4V4grZDxL7WW/4PCGRlfz0SET18k6xP3PLOdx8QOG3DRcNhIePJn
KKyHzg6n4ZbTkDKGioeV3JY2cnB8ibRj8TRA+7QW5zbt/96PtoApknJAmj22hbrZ
e5RkAHVTNlotog8x0gagyjLHqHHVedxvq55x4kiK5erLbGTL+ejNt6cRnVOQCJz5
QeWhCDfyvfGy6y8kP6EuQqDiLm8S7b+u6CqTpLLqas2Ra38OCfNMr9FKi/YysRwT
BU5vMtHnunsDg1qnuMur/SnqDsRUOac8Hrp2K/DhIekkjOivHTxElcnV0bS6n/vz
h9cmdOHGwt8fGr1yCvmLlnEl9KSAorogFGzgml13fOfUmHGfKIpQhNFN7qn93Eo7
mgPlGQoULCD35mw95RD1tBhrzOs3nid5KjTNPe2xGeOTvjB9YaVMduRn+l6NpqAN
tDpm40jCer/DcceUyjxQZG21XHESeMqKVodaOkwzDlBUag5qqyXgqfKwdAVpsi3k
iiax/tYvwVwuszu02Wm3tOilQFe9egOz7lOwBiPxZzFz/oR62C3SVyOF/qLEGNew
6u2O5MinIEddBciT+QMAfef3YOOB6fQP5Bimpek71wuAobmN6Oma5RUdc5s27i1e
W/sFlkFLUTtTqKTM5hW8oBthHq6hnfmX/ZF9EGZo9I68oUtQ0rn7uvcg64ogBDWz
frcCl2QP7nexGLh9xAPeYEAOn6mKbCt8VSwPFUYe5yKd7+rEl/hkwUT1A1emQTSc
XNg7mLbD4e0YNQhaV739L9UjEpzbCHgLmCbZxgiUyUupuDYnxS4qHivroQ2y1bPU
mwzmrjqfQ7FC7iXXohi/jXl2MJxLysi6nrjE0fX09jWr1hDTp803RiP4w690y8cR
+JqrU2gtnjaWD847Y56l6Nsu1oCkFRDY7Br71emEkzBgb7UtcnI6bXtixKcnyy0T
WTeZPrc3dZNDcVzhG2j68h1w3xbGrrwsTVloYqPajaZq3ccDWCOoKip+E1neINmJ
uugEGy3wC2y5L/5hFIltcmFl0x7fVOovd0XwRwuuGGiE72VG+JRrbbg6fOFXTRDS
Q1lJF5M3EmE5H9vdOudPefJQRBKugSS+hloeC7Wh3y/qKZ5jdEMpxhnQXgP28hbe
2IuSEp3XCRaSze3jqHuB7KiIT8Z32ibe08JHqGi8Butt0Y7WErz8YLMY5E0AgBbL
T6joEqRgbQB9v6mbfgealIW7D3R8IlHcCU/Ee0e++34UlDGSnyuVibd9cJhxu2dT
4N/RJyriO2vF6RLK/+6RkkJH61+xvWXyCUIamdoKET1y4aOIIXa8TPGWpp4Bt71C
I7L0kCQAfQmjJWQoh+OrFJCTC5a6zPGv4GjBEKTM/kcd2VdRO5eKHn7RVTWs6ZwR
l/xvKuHD9i5P3wNEHQiW/jLFyEDIcS3aqGLk+pb+CClNw/3ybqbwyRIrIUPOKFbI
9OVdpkLYXIkcYQdYigNrF0G89OkVGwf2OIZScgB6cg3bZZgX7C7/C0gXdjxH66L4
h2zac+5Lr8Ij7xfDfHPLZTMzMW8SAxvrjNKgeyqkIprZ8PVxH7vm3f4Y5vfmgC2j
HQYOWOAL9VYe8jm/NlZnGzkkYAh60BaXu+jo2rNV5SOie+kNIAQTsnPpei70B3T0
WnFYlC9P7IEfM1oPXym93iQr9GHo1+GjMkxO8US5rT4HI9l05xSHqc7sftZ/xOY7
yr2tsdskE/SRVZyaZR48XwiMygRORtueHa9EHJZdOEBsz1nsJWeMeL/KoYbJc2gY
jlwNbab1lXhS7aszBy4wXQvRxiEQJDEfoBn2m2Mx1gyDRUYYm1/+d/HB92OV74Dv
dtdH2pdka8FT+edV1gV9zoTpA7btF45kNtDWbEeF+rgPlNKVuiElK2vVphm3MtdY
5FK+c9Nae7m13baUQ2BkS5WlHqr058T+U/QAzdYiKjgEWBsrM/cbldS5rzj2IO/B
+iS55QpfNarKKW800iVdBT2vL2HqJxK5IDVq+PXKtWdRmvikAdfhOeVtsKqcVM7X
tDId3QxHIvy2IOdMNhhOZvTuRG1r6LYax9gLY318FkP0iWy4KnL3G9OT27eBNFGZ
RUlESqww5F6pm97Pneo2ve7l+WE11AnI2CN8VYUT9SSgvgwaHWkbRh80bUSnUIEV
IUiukF+a/J77DEkMMhvC3/9UZ9JxMt+zBQUhPdsn62scsXNdpY0qGpxKDSPK8gxO
140KRnGFQcPxOBNS7oqmPfso03r/ffWE+q+ODi88BVPyPccG9mcq4v66mx1oFPVl
/cD4QHp2cUkfnjFYYWQNbcd1rW9FPoyct0Kq4+DWp+VQv4gwdFVadhBZJ/LzXHxg
Vxu3zd4vLI4Q6ZLELEVbdBDH9oYQahh9HwCWi6mcrmlhNneaxkV0ajMyujO6ODh7
dlbcuDYiSIVmvdlb2ggZ9xqhC2Ko8DYsv6zSM1OIhNujigs2I9/hKbfpL8JAqXhm
GTbFDhJ+pePBPpOPuhNANw+Xfts0S7Cg0bXZ7O97pK+Pvv6zcAAooo5divIXjdbN
71LR7HFHI1GaAwLZzv+1o3mZe/9nHYw89oGb98vHUrinWFrZY6F2VfCIfRiuNbMG
k0H7WHXZCdqwtghuZbN7GEDyr19A2cuTHgBbBCt/IhWX4Qf/TgGzTVXjTGcZJ7zu
j91VohuTXOTzWZ4UNmsA299MofyHCQUlNCR5piRAxXFQmUdDgGNo6XHxQ37YkzXP
pZ3xSgCUPigngbJUqM8aSMrufA2iHPkFxaq4sqU2rz75b7qxmjup1AuHVoMVQ3Ug
k398EdLAQ7uY5tf4qqodLM+G28XmFI+E7H1JsM8iqZFkktPL/Pdk4OmKjwdd3l/9
7Q8VmPrjTyInoGhOudRuHn36+03Gs4KEfdaATgPE3HfytggzVNNeDfw3uywY033u
oT2mIpuOK5oGvTGtw2gs1RA9tbaFk+iZUC6ukJ5TeXUYuuebK1RCc62vlw/KZZ0F
+1nhr4qhb/paz5B0gMZxgVynwFcy5qTQcBLs88m7Ccim6VX1ikhJQBjuWvGDJb02
a7+adH2DXqhQnLZ94tNDCTiGBAY0sRafQTREIzw9I2KZ78D8vOgKnTobbhV/qpmO
BQeBYq1pXYZWaHES/O+Pj/UgpMWwm8yXxCqnhpmCmmwZCNTx7VYgInV3tQv6PwMl
QgApZysuXRZICy7zgijDSXDTnNl1W+c1gy30UWd+7a4HpswRy4lQggbhgZYW/uZS
phk6yub+VoyZVMYhJR1dMmoY4FFcmTMPuxHIdJrGrgD2bucWrBDSf6S4VpNFqVoJ
7l9/PF6zJChy1+X1WnWNgIGk+pnCJAb+Yu4OVY7Dio6UhmBJ7NLZ1SpSIqW94Z0s
PxwEl4l+6RR29zbhB+9xggJvg2UQDYGCxigRZJDV3yeuzkDRWu05qMeLngFx3pB3
fqTttO5VkiMmjNeB4iYtECpK0bz5H44VhCnb2BM/WXKtd9OqXINwT5W2sMW0Ofb7
9BLq/FYu8H+FLGq6CH0+bElL+Y1RnUTvfLIdqfCpQc43ZoFOtbHINP0nlia2VeZN
20diune4Gb64E7uHxrd+35h5K31VxEk2FfmBTdAnwvJfbOnxp64DuRBM4HPTa2Vh
QfxSRymGlpS3dITMIA93wkwthwWv91TLYw0SLB6AvrbrGpafk7qX7uB3BMzJXIT1
4nwZe03jdKw4reVlNqSqmw10ZKO4Wkm566ShiEJAfq1z5Hov3c/kZ2Mo1NLYgZ/I
yIr25MwZRr1Z/ZtUIniCHkZP1bdcwvmr8NkrHmM7HmKL8veTPf2tcN08t/Uy9GAe
Fha52YcCzWKeBMWtJAd4l7Wx8QE2l2yCg12LL96r8NUNbYFNzp8APLTL6wEuMqiR
nqLvGJcg/fO8AWhyewSuvVTRWaEuJ3BWjEyUw8gQjhJVwujyezEKcn673K83X1tU
0E0/aR/dqsYaM4SSKqq7cgr3b7LC6T/joKbTi9vsGGlbgAyE7bkCU9s+zdu4lDw3
lTecWDlLFWwk7Z/tK4zZMyq5wfO1lP8J+KueGojBiKX3KnwFBGMpj9Esosj2K48+
ievABgt+9JPdqoe+wH1V4waL7XH+jz5WwUBRCaEdbAWGKMklC3pSQce63CztdnlR
nksxI5+SrYtgfdebU5tCqf+5/IaI9tjxekldJ+Muvm2EvVwGRQn9GWFYDaewNaMP
afj+EqJKph8HV6icaDCnflo46K3erfVVOfgvEEue7rzB4WLmHIyrp3j04LQbxjRY
9JANWIbZ/UkaWyxea9ZE+U9NZzpvG/3Qllst/zpC99WJhykOSkA8uLTNcZOlsA9z
LWVDGrRmJOGl3QKN7oet3TBZQzSeB2u8E7mMrlzTv9mLXkhVSN7lqPsDiXaLmawv
BQtdaeq9gp+LlgGz8JwLp1g4+T3Z1MwMSiZXIzuBRRYg14+M9/QWssD+eZnG0kbn
I2Fsr+9uY7bWphsD/ShD/lWPMVQ5R/dmnl0dD4rztSWqQ4f1FvREhN4/e4GyHSM5
CuX3//cKoogHDpPPYuHA9Ag+4iyFFqBnjQ5K+mQGjElkhmTvTHt38xlI3gEgB9pi
ybVLL7OKJoB+0kXpjXsu56fJk0Ieq7cCGkgpHmLaROgeQQJiACrpzNNUNxvZ8rTL
MLQiiCmymdi1OY2S4hGDdOS5zV1my7rxOx1tDXSzTgByzbGKE2/FantJO9z2ZB06
+6b4OvuACXnyW1f7UT4NbSBQ439n0fvNaxRSmfsiVHwdpVMipSkae/sa098AWaob
Mnx/yuIfUrpqW1R4R+E1Uakw2umx4H7JaN1u4v0k0GDzCvpYgY6bvCSKoDxysbTO
NpZZMtAHIQdq0ynhJ7LZd9Cqv/aczxyUvl7iyEp0adf5JULGUqXXY5mtG3jnQZBw
6p+oOCRQ/rNBNtWiF7b4jM3Z3u5wrzO+7Pw+Pt4BW8mj987mHfaEopmF2vtiIdeZ
Ip1nTPBzlaAex/HvQihgYc+GWYA2WH4n945F6+9402fqksNbkcDT0PIQEHXCHAS4
W2wF30L/DEwF5EqmkSuPHdltPyhwaI7C9KeecxVURU6AtZHT4bmUdqjESNPR64Q2
4sYzK9n4ubttyzK0z3TTZTg9FkdbIclZHBo1mBrWg7IYOiDnYzoXKeIuyopYmYva
VPDYCcTX1m0rlk4V9O0J6vZ/T99jL2jyov25AEmL5nRLtPzlFizvb6cyz6D3KZWW
e3iudJaJKgqyvxb6oJygU70kpKTFTGrht3urtddAL98McnmzetiP8IuI981amrej
CQXzVutxCO9vlTu5Dzt8kluCEohB+uBA07oP33obS8sG0FM0WNK41w6Gm0Emw5qH
UIfKUpcaNAzff74pRppRPZVf6REHcoM2O58sLOLTetJLI86hwjRmvDNvmCsi6mYS
aRNQ84mGf+212gkzdbe9UuHNkP1/vb0jf97UuFWvMDYaDnRGLGsehHqQa297pr3u
LwVHyuOftIE5p/tDgKRyMHF3/3nRMPvdnNmyO41TYojZYRpFKML0W5yd0oSSdHm2
JO+jFCV01hSIMgQNnaWiwakHGIQ0ifkt256VHNkkrlUsfATWxgHVdLUc6zZs2tet
48RLGYa9FSsB5qDoJdrln1rPzrwVg3e3YHzV38K+IOhqfPljPI8hBWdAgQ0B89lH
V+Dn/LeageVY9A6CSN7EIT6p6J7vgFV5zH1vLZtVvYf7HHc9cfPxZnuH6Te129Fp
211/8ZKwzJxDq3I5BtTLJ/1d04SGq6acVd1mKkrK8P+ll95eMU6DytF90cMiQu1b
GOV0SPUERvISngqFahJ9w+Y88ZP0TYD3+nOWkMkgSierp5zcOLEAuv3cHoKqjFR4
yKekvX0ZDXiSbNLWhu68wEolU/GCX1fEoucixUx2FArMe9jEMhzPRGVmYvfsLcZZ
H/n0THP9XxuDJh0UN1t0hU6nWDY1u1w7+HzRp4j6/q+xySPK5f9QrPviHReHSkOG
1O8CNcPOWRUVGCqjfuZ+7midGNXd+JaTB8mKXUpWWx/ALc7hlHBhdBGfuOLYxHC+
GBHA7U6vE6sQjFOEuMicm4piSKiR0O8I9zxTtuP5HW0sHfX/NIIE3DxJlcTkh1L8
W9Rkulz5OYBvza7ekMFHwb7d/ZkFrz5d2MtVimRzA3IzSLAJXfu4Ix3jo81Fb8BF
wEOS1A0bCrJ3DhpfXHmVR+heSxyOmL04UueIf3anZq8jOaZ0/Z5e/7ZdPSE5bTQ+
w+8pixpJ/rpeaNHejyuQfRVfinCjF3tmJtlmW1w3MB+wTTTL1EefoWYqWb58pjmi
SSzTJYOpbb22bcWoLbRcYMAho7geJCGesm7NDQ8CML0+fOWkyMs3GLwSU8ZdQEjz
kEM/K3T4xv8zqOtaopXAe2Fo54wt/BtJTSN4/Bl/rGr5Lja+NEg1tsT4nJXwvn3k
vZCSV3h2y4WqOmDsQPCKSkQvA59g8bqI32iV74rVjBbdAow631l1GZsi+JTOoqJr
tWO1qTgXs7WriYnEI/IC39/bOEgm5iakPm/9QOjIAnI2KHi7bw8JBvYJQJlkwhKI
GdTPrB+rmk99+vR/xJ9/ZtM1UORW2dVDT0yuFXrGTq84TBYF11gTwxZi+kDfZCIX
I/icZsNe5JouVDGVxoa10nL2QCwYjzBmOhcKE1fn3kTcxOz/Xq3TcxzchI8Fu/3s
MErh2nRwE5AVqb0eY4MyEknkvOxSRZURo3No4yduMV7xeJcFJqzv9wciJ9i2wr7P
mMFXP4tmqbtd+e1RG5DCuDwufB+GODa9CyHujAl8ooUVFuWwSVRwfOe1joHPoBy8
ayYoIHsTMetmiOW8WXjXGTG3/hmh1xaN8gOgIe4RIUsfFELcmmA92MkHCj8RdkNE
lmpDKlC/jDcWMuIMXWk/YirWdh+rwcKi2EEXJ4jp6wPuDltR4AjuVIct229LL9hC
Sc+PhP08yLeFB4Uw+fAP8Grx6w1c6F6lKk17IYw91AE13/gOwz58mrNbK9O3qADu
D+N+g3LDgfVIire2IW8PvJcLjlYLhpOTKI7cZgoGN4tjBJlEGx4XvYodWsMCNHxz
WxxY68Ab6hOCiEKJfp870DfkiPK1ZZY5d+95JPEvgwZAbSEWGvnGc4QLeQtWNYuV
dosbLs+tg2mk14MtTI3hFOyziNPTSabPFGmU6N7zD13a5zAmlc7jlYT8sc3UrRzy
uRPPEspnGfGbfiZnB6VVJdU/wVedxGB19P+OOcFgW4wkxZydqTWzmlW4wxqFg0No
yLjYr2A+uAe5Lg0B5MOX59mE4yP/6Q3XxWclQMhnuV9VvjbO7jhe/sepxXVmEnn5
NNws0KGMyAUevwoqX+cAaJR0KeQLKH6gxE8k9yW/xE+JK4oWeH+umkV5n8//KUco
hxqijU5rLh27gO5wHt7pmOUpVKXbvkupR8ACX9uXS7wgQar+KYLxt50Cn2kOajyz
PbLl3RZQh3KCPyyt6DoH4fK8xU80Qw17Hz0Cgxc8E6NOY6nn/6JdyaXDYXzFHaHG
ZVfuhkFDIoWWIj+GAQd/3PQmd4LVuRwcJNIxVmPO4BPJAzdtdu18XBGaawZvanVG
3mEOcUuYTsyOYKAdqKA0BYQ4eoHEfcIonVL/TKXD2C+8HD+WUhsVk0GOLkLRe/X1
9CLN3WjGZfty2EnJGK2kzROY28CuJ/tGWquefWMnOYGGV2WPZGsyk/Ke1a3lzlUo
36IExflpoAviFZgpbSfTPh0Pi2qoWEO3qHoEng5IgbWs5k+2IbOxYcWKCd0afFAv
xFzfvWMUqU+LQ4AREHjUdAAJDhKNviwRSNs883Z7aAvDWADKgWcc5FRB/uS5AsYr
2vtdogBXgm8oHaMQ5/6dqBj119ne2lOIj1kKiPUbpdFW0DgLGjtNj16mlWAoiMtG
q0nBWSWNwxNcaNA/LjYivWYap6dIe1S7LQ9I/Vp9ceFEjkLyAmRhyxXioSzxK9IW
MjNFNy4zzEUiWFQy9M6rYsH6BmTm8cCmREdmEb9QBGNaMCjjg54zz4RkPUFsgoR1
ahU+N7PR5wLrvDup218HPCls2+lQW2nDYbJoW0TAmryFExPuaKRbgJxeDrSrd2U1
QIpGqbQbrRewBaiWdLA/j9JBWQzWHvYQkmC/6f+VFRseLEvIn+5MLXgIIqg2ywRW
7skWN+IywCBhvVu43OtiN11zt3H49LWnlmhroAmq7UcP0MCR/8Xqt7XGQlvsn5Aa
bPB7zHl9n2Wcm6A8J3bDPWWF4VRTcAV+yEtXQk3UOJMK9J3VV7xnAxp9V/zwmcoh
9TxyXBA6nGO2LuFxXfu/6ApJmrdzHJkrvch56n8cWenNtgIH7mswEGAZZqD4KztW
l/5u9642OyjQLoL03RfbuBIuVsjK4B8/DjBzrN3JT9sGt/AwfECf5wWh0kfvM3Wi
oykCB8Etl53YLisqTpuZ9x4MSp1FVQVHbIJzDFA/Jta8dVSbrQCe8Q+mAuE8PuoR
A2kB/+uS0v8gA0K37Ov559me7GvOwOa7hJox9WwtUjq66lPa1mT15i80pV2aAwbZ
ki69pazyaUrQ5bwtZvV9jX7UJRicHGWwRBNWgeRy8SfPHdY9ygTfp2YB1wOWBkg3
B6QEi5HSAsNZV/0AcjvmMHX285TdkL+I5wUJBj09Odu9RH9vNgCr5WRF8NE3Utku
n5amF+31Uj774Ci39hsGm2QKCtewtvRaqpZvCu4i05/5YosCbOxad4M9SSoCNj3+
b3O7fMYG8Be4cVqdpbd/lqE4r31vOAMmt84TEpH+pWsRMG/3Ds+pX/L3ibo1pVMd
wM29M/uCT9sQ6AS2aodWzuSvGchXt12u8WM4npKhPb4Ob1tnsH8ySj2xx7D3Ucd9
yHOQOfLmJ3lOEBAbt0hN55n46o/20caah6t4LKZ3irpgRZo5YD6GmoKL2+PynVJ3
PiE+WD/ootjoXCGY2SIDKJPgy88MxOKzEpAJqtDNDEa1FxuosAjza5YIvdbywfnl
AXRin9N4DOHPQwcAKlo+Gw3+GKf3gi0Lb9VuhaTr1ezDzd88xPPzWD2bo1hPt/F6
Xplqu8u32Cd9l5AGoU79lSwQLXcQUXNL34yUIoJKvt4JrsDO+o4GS0Me+IkhL2IC
UX768lOBSvwiLgIzsys1WKe8D5X67xtSOS4zVr5V60V1bdEijukatuxCESzU6ko8
/vl9mfltqoBuJneEe7HzWd/m+coGyAxNZCKvrcEV6VYbN/KRc0qxS6qGq+IYmlWX
Q+NZoDBlN85k7OiVlT1cuXhbLf7zSJrKyDk0yxSB/J9EvBVbu+GHyncZxdDGZNFT
M+OFQdCQsd2D/b+2Edg3l+8whvJoKVZKLmMulO2puuDM5DV96nGfwV3b3YsKLbii
LOpKfbRkWxm9V60FZy41zcUBP+hmVdVhNwF9eiBq1nqzGXsVxiWzg5syyTtb/er+
k6lTD2z9Bww4msbQUOI6QTx/PWYU6YvX+jizkinS5y5Ik3+5Zml2kY82s2NE/nUX
QudipX50eEXp0VzqsBiMszo7duORwI9sNJqUVi2Xuz7+SXFCWeurX2z3tH1xuR+A
BGyUPk1rUqe7KvkR7T1h/Wr9t+tYKpTPtoXdJt3ITFdmyC5qcyCbuNRbK3LbmbDd
4jmXip03+gcWjNb8A9MbiRaFuXCLYDPZkQbvElRkQkLx0vDlnU+tEExS9gwN02ZI
fbatQ95hDk0EYywGqdhxqBQaNeyAyx5kfoTb3CoXizQIGtq5Rwl/Vcu+rQBSPgzH
Y1qVWoDousK+MuLAH3ggh3ZZOJY31SYNKwBQ6DXjP4FfyL8Xd4PtsArgpOd00JgA
+57mbZlBqVwgmvTuWiYCHUPx8juHWqNp1aFfn5Y1pk0lfYD5YDz6LfCc3aM3ScF5
ZvAsU2/CFYKFUTlK9opGVciCp4WfH0/M0MLB3WM+JDz0r0U7gCRe+mUFcEtqtFWN
JBCxetZ/A5EAJKjw4gQecIyDLU/Lk5hAxDEVi1pvTX0XjJ8l6wxuMgFKl7U98r1H
zU0YBG6SxuR5HCbDKUZVqEUYC29F51Gwdc7/f9yhPe7f18ht6QThmytsg6C8sVPO
zlf0Wt4345ElIZckL2dU52uwXDtDsHwDZbNqMO2CyQJPZ5GfjV6LIeFBAJzd96hc
atFbrZjgwMKMInA+Nek2K1QyNDXo9AkNWWY+qDHx6jMrEpMFmaj9iIoYFbn2ZFI5
uAFSTG0vTLdvD16qZYC1czK99+faWv0Ga6OaWKCxuVfF+1Lyy0KXvdH/FeoWSvT1
aE8DSeRCNvfFoc8szNI2grxd7kT638nR3oabcAOKj1MJC7LLm7M09qs8QuNIwS3/
5Qo+Ges6KEd3F4f1GwaMjOe9z5g8PqdkuQmQ4PsJgYb6chZkfWQm65hpUXNUW2Wv
6ta2724NxIazIvLE1PsyvcJ32sHUkezEiYEqKIikTBfwbgYaVSdrTpyLQBJiAibo
pQ8JV80u/xdC4Hy9Hcp0fAG/EoVAFwsisL4w+c13gI6uHOdUTUSHRi3FnlVxnxiu
24hTtiHWJjQJu007K9XnEk6yR/yh5+/8gAyhECib1vN5NTmbYJTU6keF07QkU3R0
j9i56F8ETsej0nYKB3pLEJJ9wXICz0cusY7lY5EVB+6RwbNDvuzfQwreLX8yIwac
kIUemTu9VbnLt7CIpheWNYq9VkKf0If8SbwtnT9AsuGRU5tjJb5WjCIoP5icqSlj
Yw64nENT9+33/WB/hoMacWnWDscCJHeTbw6y1w5pl1KTGLzS1BQzjDW4//SNf3PT
fnZHsMnPsaZZtPCUqMA3NOm4HX9ZxVUniDKdN79vT7nJOBWKAgUxMD+ANORQy2VI
B1vsHbkvHB2FF9pSam//irTe1KicZhrr/ae1iXtFCE8GsPRa4NtTyZ5NGg7MKf1B
YC+LUhD5O/a/tEbeTJw1htMNpPQqusKLP8NvAfZwJUNU0W6kIZogZ76gV1CsbiVg
CRGpGZSNYMAM9kbVDA7YbzD5wjNt+saWk8WpmFvOGjdP2qLZKPWOZlv/a6GnJLjQ
LudbjKblNP/ERZovUhX7vSE99B6fNPvHh/yjdIuXHe2NFuMiUjndO7wSueJPVxaJ
xh96Mfp+dXYOh4PjgM9/h48ZfUvyYXyzaukcrsnsbY5YGwGS3A67cyb0ftlJ+e23
aLiKQO6K/coQHUKy50Z1Hb/x12kHYFqU5QmffADmubAtqzW1W7VHUApLpApepW61
DJQGXEuiDkQMSgxYr+hct0p+SQBziYZZiHmodjFROl8duahmJ6mxvzvp1SK1CQtG
cbxnN8QRXmogQX7lOuCPNWUdFDEunMMiENuGpqT6fX6lWaW3faSGnNeaprhuog0y
jXNTmp8chPMIOlTxc0c/gyKPsgntE6zCl/NWcxiGBW9xpGxMdL3V24mXBF/lG87T
j0v+IucnhTU5mKDG9sAtAVwCB3IFbJzUYVO6CO6w4FdHJkjYaanBulZIfjb8Nt4b
TFkoxFO9x2uTkMj/DRkcBDfoO6GBvJj23jYyB61N8EXip+RoJRezn8eTZMToKew3
NlYVw0RjgI7oyg59H4PfD7LrzuMIGWQmD8Js63GOUkWGzi8qt46oJ/1iZvKrWY08
N+erj9UiqPIKadmpIjMG8Vx/JvzHRlKKRIJePIUJHb/BFUPHHpI5YMnrH985zO4m
01Db9e4PIR4DwrtRqFx4s3H3Jxkhjk89DkS1PGmdrIfl+QM+kYBE0FgBv8Z3HT97
CV4w13z4IgyLMFN+XPRUz9x5U2x9BN+YD3+9g2ipPE9ZFZXC/uEFHa5IaTXULd7K
bQCYu7Qu/tEV/LILucHw0pa7c3fQW3gNpmqIvjBST4gSZ1Bxzt0lHD+lI6LRr5uw
biXY1s0cz06Bdz7ErYParz3dOnY178WfPCnGlzJNW+BJgI9XugriGzyZdS30iNaY
ta9k0PxK5NJCrMPCfSrkCCoxCrD7X4rQbib32phihYTLt+N9Y1q5kgLlGhlj8jcC
9xoKRgsFFSw7dD2VSYtq6fqvZdCAKSjvf7rMS5920m19dnv7yYh0ObTd/1XuO/7y
Q2TzkvBKwZt9LRHk2JIl99MVmyJrt9FPP5PU3b+4AG8Z7DhzAr/cRr2GHGJMDh+F
eZhNQ5xJD+6ObPFbzVzO4rtOqbJ4Ctp/o6+u1IlzwqwhKPbbRZEUX3WAXInayHbY
sdjVV2DPG2UP/puRc1g9Bd+3AwkrHefkqm3aemySTBCGUDeAdW51kzzaTj+4Votc
K06mWbL4d5kLuBAdmvB2xq5v0YeHzA2c6LMg8k568A8C0+0VmRIMS848a5cg+tTy
Diyhym1rASyetViQhFgBLwnESVO0sjM94/OOIyP8dAsT3mse0OWMHwAZMiN4uHeD
FWaA+amHIXKSRJbi6S2Am7ltpOBoeCSmMNTp+EkchgdOI1ciXGQz9QrLlEIv+4Gh
b9DsKm/d6HM1TV1rnArhcMzTKihpBg1vTgGStvcUK2KzLjExbCLxYyOTEF5gEEKK
hX5eBdp3aBobCjdbwTbMDcBXmHRvuz9SO6V/j2pnOm5QAX8GeQLG2Kp7vZF7FpoE
HgmSg1VI4rrPpTg7bm8D3ft92T+bbwraJ2tfHHNGeazZgPQfD7d1pHp1BGVJ++io
P0o/X1msBtjOG7o40MvaK1ZpdQ0LGoRkM+fgNkDy4IePYAlcCHIx0y21nZAFjORV
+5o/ECJUhhBsqOlJGObMeUEQ3frVsgOP3PZ0UB0J9Pbbx4PaYGDWwFvSxS8ydVD6
WM5UsOTHx1Igfy1oZVrQ2B71WbaCYcdaluIJlPFn4UTjTmef1JltDAXcTc8A5E2t
2q1Qu0RucIJcDK3wZRVNSnCK7sBfSLNw2ASdWi3Tl1iop+HypgW0WKhHNGq73mW3
utN6HNxmoqLKLZn+5FslUY2A4wpSJet6ENAaCsPIqiX7YPvMmBmTeiY+OS+Y1wFA
9vdAHGAKzIhzl1Xht1inYonpkBwQmT3xet90nAgvkHiootbcHBmdzVyhq8xU0zfc
ipuctkWFGIFzz+6d2T8dR1phh42QRDXoSi250oM4Ios4koJBimchaQpUkNPf08MM
ncGS171YQ7ftBSNtQxdJVFpxULVgbLe6BsKCF7sps9ZUZmV9cs+cHzDhk8MpoTL/
SWx6fVxXhXoPZKtav7GPBSlx8I1Qvz7DhGkRtboalGKIr2seaqcQNU4UL21Y73r6
giiDs3Y8N6ruIVr7pbgzuwzN1zJnvomRj/BD6mULdOjViugghG68Y9jeI+QZ136i
Udrxgg/16Lbp6QrkN+lq9pnQnByRkq7QzQawlz2LeSv9OS02ID6AKUXb81AiLnrr
QFguNKqJR2Lvr8U6O452ipSLhuRGaTmSCO081z434vDAeWS7UBPnwpJJKpszQ6rc
G3fceZRxNBESUMg7iV3X2rxfyyNnYesdmw8YV439zzXrK3J80/I6RpEvB8tjTZIL
ly31Gqu64iZ+uFP2vpxzZOKI9QwNn6o6a7LpOTM1DhPFzQKsrJXGj5K8U2ELND85
SMU80j5HVd8QBJfqVpMatTb5Ar3qwtz107D7ELrsM2qD0ePqofqpmHl2Z866LHuN
Cu7No6xFFMng1dE1dy+XQJ26EWJGhkmhAdZCZJKkEbjO/brzipHSW8TxbgPz023w
Sv7SFhhIUmxlvxYuib112EeFSiHM79lwwwFwmOH6P5k1pP7gSKc1BUgBFktMrcA/
qMs4QtgJNGDsBtMbB8HI2lnx1ovuVs6d0482Rix9Ruh6jBtlBY0ILnaOpQ1N8CQF
xTtW1rL362ZUHrc6fYgWzSjeWQ9LA/AUmWnhb8A6SxBB+GeYW04431sDxDqYaeVQ
8ixL8e48peJ5CqC8ekYptuPhf4H+KFO2hP7Gev7uPE2yqSCiexSzrTbZ1+vlg/bA
aEveEgbOMoSrBshptE1ftAgfQ7SBRqm9ndy/bDITUCsPLB/4Nc/T1+sC8ZXmgcOx
kXJ+J+Uoq6FvpseeY/fF5lYYtagSXKATq/7aiG6xx6pvmn+s+EBPxzKpLTAtyVt9
EJsBT4lsRfe5O188a8B/UH2beAQqJBowqn9b2KBVVe7zn2VXk5eeI3aLT0xrErgX
tojONs9KCeLG3ZzF903xvgjYuEP5dWa5puVwW3mEbKx4UBXj/UUkKFl0n4Ezs4M5
BkVrwMTErdikOywJCFlDE3PnaYpLGJIHrIO1ezVyQEs+o1kBZqkUVPb3gcLf1fwF
vI/CA53L3LQSpJBcAqBJVwI+PIYgWZaXTcXb0Z0yZuJV95ZSEJrExjGpAS4tFKHr
cywAAy+aaMel86347DKqN1VwCPfRNDQcTG0y0OaEdXSl/qIxW91Smaena1teuSMe
bxYcGnctP6KcTVYy1viQez3KRYXdk4oZXxjYGjiBWm7f2ead68k0G3rjffE4pwOo
HxkrPDI9Mpvda6N4dzcKX0TfwD4kiaKn3i7acy2HEOqubZ1iLNZLItIqrZKILBF6
w3xxRA2WgAf5IXL9fO2SKmEFXOTVWPIdtuXZQmgZQalqXJYf19xgqvHW65lUdBlD
6KmIYq/ykGnBK/T5zXqmTeIfWiF94DnFiJBVyaT3AmmyiHApAdqCbP7XLuwLPgCW
OJyX0/j5hw0VyuRedRkZvDB2zMHT6i8I8MjbwisYCxUvh3jQw5tC456fSlK+hMTo
VkI4WBaQUrRBioXW1BGeIx8c5L8PPxKm6mIyrF+MOV4XkOwdWJSbx7/TrU/wzyJg
eKLkDuhCL7kNfGBM9TXkUGaHTiVXCof1rr7hbTrt1beaeYAY0+VUttPhG8HpCvwT
hfdcUCfvduTk98sCylIGRE6gd3DwdH301k3xoF+ziPIw3THTaMrd7rUy+pSbE6eX
RBet8AxQM9GaDaBRvCc/OnGR398TW0+VgXYEw4LVacHnryDokMKh/rVutuIze4dl
lxUFfpVJvyb5Q7lnJ007hNV5oISeypojlqJzWW0y8sGNtnSg9zmwZO/AmS0fukis
tXgALQJDIEWRViIm7NGLgFRl4AWZeSWUPXXvNFR/WWqEE2zKEWWorN3G1I1ftFyL
P5+BWK94I9+lK8S8D6LKhVaDINk5cZlbhShPgplmLksBL8tYPO5N0u6zxnmXKoWW
7vMZewIXJxjzHkf8oBA1X0NTxbVoTqw8++Qwc6+jIdIkCSzakQoLd3r8/mTNYiIY
VdKdThtYFct4H3SFcSHZYOuGoMCeICg0tdQZMSCCnwBXLMcl6cTcXY2IMxQrNTjS
E+umzUoACUmw6g0CeTZte8HdppRRQrEqZBkxw3TyemlP4CJ9UlDLDMVd4FEtuwj5
4r80y3236BtK3ov75PV8mGEfXxRnEqn85JLE6ceqG2iAQ7YCVkq/6xToLaQtH57T
3NweXysp9utrP5WPbiCuz2kr/twIAmPAa8Gxhi8kokXZ+yyrOOPa6ytm1oFYPlCV
ZNpw/ESd6MjQbwDj4bfmKccMsIIuIjp5CJkqPM3kI+dUenmoDQf1D+U7hNYAHJ3q
Lgp1WqRNftjwSl+iO1F0YuZ5DkGFnlOqszX/dQc2Zj80m+QY6a/Ha1w+pl2dYNZ5
KR3DjhWmSOarvNHB8AQmLeNPiAwBB2mWjrC5HDLMvw3pyrO1d4rJakUc+EuyvSvp
g8b9Z5BjmGhqN7BTrlv+I8h80kCTGcEBe/FQYQUrcojkz1uDW0sfNICkAKnbZWXN
lfglsn2hQVM6uoB0qr2hewh4Q5nvX0ev0ZmBMICwM/0kC97zcJY4yHEv082xa6Ww
bTQ+9f+e9JCqvukakYcY5QyOiTd1lW95sx3Y+8MbrkFeBhE3G8Gxfb26u+dDp5Ei
IpdK2TFNH1ZNEbVIbKp5QyT/bVoXB/Ykj0zZfKPq35XagfdVacH4sdtodZ+LOwYo
KEKlCFJN64Vc1k/8JlKinhcxRCObTAMac0vWJh9dkU8Qqac63C1/RGhExdVYN6kn
5HChv/9GFjVW1M4E7jKu3pNNMTUebtG/ZACYOv+CO1pRMRwurSuwaxb2FMEnjDc/
mNFuTD06pSHKK6g/bORPoabbYdvUe/XBR3fFWfy68ylHNQUpkY9bQHZ+sbFiu9Dv
XwRwA/m7pp/rR+wG+9Hlw5XNeKg47NOQomt4t0mynvLOhdkTgu/rraMdvMtcSAH8
XGLOvPpaNywInMMuhVRYEsePkE7yXBZTJ6mlGTYLmyv/4c6DFkO5Wl5ALWM/kKU6
Yi4DDcRu8A8pTmP+F8wH8e8q5L4FDTEbosyj7XqTLauk8vzGGH66B12xT+m59d0P
0SVjVF/FiO1hJMvtXMoh/7t8v5v1ecjpLlnTfR1pasK0igvY6WtWil18ilzkHVwW
dsZPtF5/0QNcYW1UUcKxcXsmaDGNH7rqVUhbaRNpd/uFcb4uKXq2kRvi5xxRZ8xa
HcCchuQKrDpELyJ50m26NbuS6AW5GmmRI6QBPxF6lTwbahlGsqEi/OtkKIrJZXh6
5PbBpzB3MeHKSugC1CPPj9Iv9OgkRmIwAR6HHZQyuSNXa/s34M/MLwWmODcgKUi5
K59AhZym4T9Plq+0VtdTvWkfeLNYEA6k5sexRz37oM+ACiFWub4HfPfPHx8TXY+b
68fgcISU+sde2TjWxG2gVtqT0lWragX+XXK+sMIUCxOw48YMsBkYmMw+k6dLFMs2
zCbyMzo4UB/yoiJhxncNhKzaVzDzfh5yL3Cr9DVfexatYkE10V17+EeBiGxunl6d
+sVjoBWR45aRAoWaPOrJyStUHzGotEEaV7r2Gi3xk7sIZDmSRzuWukU9ov+C3kFf
z45WtknnznwbFG0FaHp9f4pwlOwDB0JN3e+lYQuVl83/JcZzeFQen45KAjJRKzKj
2FCEVCDqiwRfJW6rhI4ocu4tjNkf8Xh/ir/l1u2Dx5J522lbqJ+wul+zT+eefli7
PF1rRG/vaRrJb9wCJUyMSC8rR4FRTIKebPU7+xtAjcEl+fMV4n5r1Q2IYZQFnTP6
R4RZ3+oJTrckH072J/DrbPDY9OvmesSgSdGt/kd6WfBtoYHxm7zsYqQtnNEXN9GS
Mhxk0A+MkB/enqgMyWL4+5pqVH0GIrI9tnwf7mIwcfo424JFzq5hujxmjlIOD2Kc
Vprz+/9KruFL1u1TD6eKvYtU6v/PIiE3JUIYThZ050pLwHLZ9NTZdyl9jUDBHyxr
Vw2Sd4veUfceWZy3uovfpCyfE7E5FaL/3rEsPGW+mFszkAv6qAxI5e2mXxHWG3dV
rGPKx/DNTwtVyqPN5CqqaJi3PtAafrmQQSJs1Hqn6+/2+px/BG5tSVEYs//+Ah0i
q2AyNP4IaOBGYYEclgEi3kmQE1is1WWan7uOV2YfFki6REIMgQVL/o9f13kbeM/l
eCALHk8T8Qmb2LhEDXXbQjppJrwgC6cvfpvohhebgQvoKYCMVeTjkoE4yQewR6DA
jmHKV93ER2eQGUVl4MZGtBClRcbwD9mdiXjAVffZewSpoJxBFrbk61hlvxm+j1Oq
ND+zSZVP2pmmQIY7oBchkujmJQeO8IcfTDhw6DiINQHZvxjZUWcC+3R8S3KYY5FA
eQv2eOTwPvq/UEtf7KDx9IycEwmmN6lhUH1ARF2A6owu4eDEzqR7ZkuzVsODwu6X
ITF0QUUQpz37pNl8r4E3SfC56JHnjLkFR13q66HiivRr4avutt+iEWt9FyMLPLzD
8Iz3BOcRwX9Vs4mjHpXGprJyScmTM2jbYN0/p4PaEP76aWVrM2Ugnhqhuhw0WZE5
w19DrD6aIFbU9JPSKh1YulODD2ZbKimHHIpR81bkHZs4mmNKIvftiKwPtFRKVQPy
7NQAt3SxRxNcz274hukGkyKA+SH+XzHrcHnXqP+AoewT1Mah0dhgIwz3VBhiBqem
/8dc/7Y6zo92sY34G0hwKIx7nPx2v9a4at3K1bVOr0WEHdpt5eUvPqOU+EftiXsW
O5KBHvsnOJp7FHRuDkKEGl/V/+lkiQve+QopCSBGel6SL6geI7guO/Ibgnv78p6/
QRdxRPhdKcGcKGB0yg8iQd/QujYRV9HZNPqYfdGOC5EVzP2Cf/IYD8u8iNhvtrZt
UXdfFivsyfS4e4esgFS6Vie/6yPrGBaVymddwapW9hJqbOMsE2sUt8c6KtXVyV3q
qcVKh0LcahGPpAp53RTXS/s5/Pv/xHvMgJydToB2K/z7QkpNWaRcSuW0SUo0UxiX
dq7cFzE29lVa29DxRaxFyw/NY/EhrevL5f42jrCw1jtSA3K4kDzoPLEuH34m/dU0
4M3uafVhrvML6R2nGW5B0Un9FQtCdMDEIVk73gKCBJDGRI3CQESe00BcKK6KtE8N
PltDQa7pnV1jUOeQF907CpeK8rPH6Zg7/YGMeezKK5/gi1E6tHMtCpRnk/Df5oIN
uSUb2inUNX0Rc7zHiKcJiy+NJtsgCBIu6rYjbfYjlOl5tL0edUgA/KOUlvflLyYF
dHZtlimL7PaCAqzHDsCecrNs/Rn/dEccHW6epMi0tHuuxuuVc11HtAZU3oBIV4R5
zkwSXNuyGXgVuNwYx0jRx78y2PqUi7RDpcwtZ2hsryCX/oxkKw7bKxgiRayMdY7W
r6282d1HWl0yElF8Mqwd176hcsDwwKvTmPphtridbaq/ntvBWvbHHwkdYqe1P58+
IkLQRBtkoev3nQK3H1LbmqHv1/tJ6jLr+UR9L+eW+eLgV2Oaj/laUQCQAExTqVUn
S46iVNOtub+M5CQEog8B4mMMtgbgmoxH84ZiUDnCqiMDQ+/wG6J7p+fvsP41BwPI
BH2i4rqBH75iCH1D6l/jazEYzM668sesMfSM6wahbhXflhk68e9+k5rZSe4jTY4N
K7bIPpufzeFZQ3mUqs+HsGa0dMLA2h7Z1UsvgclNmFY3EEI/ycRSJgSgKV1o24kd
nfirQLIUAbdWB2i3XYKIjxgNMenYy0+ElBVHIFGxCbHiB0Cg5X4rbAkzphbO7p9e
ZgLXmvbQS/bSsoegkSNU+Yg8mHsN5HJ73Yz2paVkpkKNDOIk5/gReuR4E/0+Bgbm
wyS5nJCDCiaHRHqlBBeqdR6CjZSnhKCMn/q41KqKxFXMDQz2yJ7rBvV4kkKlikKx
gJvtbV4xm0llIjtx1zbxy9YNsyjka6jbGmJwYbaIOn0oxaAFihhMOAalbYUqFgvs
im9mIIA40wshe2pYM2fK+/JKJXJ5ykkBJcj05sSPjbBKUcqGhTnUVTtu0rFsDlDc
4T2EhOZsfo0QIF9tKDg6+XKTDz3wRKkvqlZPdSSssUvJe7lWjj+3y8qp5soCGcjR
LjmjIOGuWxC7xFSAS4ei7utqaeQfWoyh3iD/umXddMZFv3NokqONjpTbnvlAvjkC
1l8dVx85c84oY6muOlHtvNAJ56n2oPPPuKnvWBt2dM8B7Ad96iSKhTYoQNsHBr5S
j4Fwxa+W2jbfbrT3i1uvGK5ZANAX+BNYADnOMePD3ohezP9ErwkKyO5Do7B7Aizd
AbaXRd56AWc41Nmw5ZVjLeh72TCdXs6im0P0iCktc/Y/iJbvhUnFhtqzCozuAAZz
mPCEJ0ORB5vN0ghmeG+sFVnHoaNXRplwUT/vQyaqMp3jaSaqp+2wn9PfRLCoePrK
fGNXIYjCRK5jfNo8XzXbx3ZADzkJJv8fN+19n49Fw3+K7r2kFWRYujLp2/0FD6R5
AmmQ+xqpBYnraekccV7dEY3yUgJ/9xB5GW6tprBb596JWcsZPrbmMxEGnhcIYEgt
OkVCnnXNN9WPMeGgwRQ42B89vDF1Jf/2LqJx9ybz8VZdWsMr9PASM4yeHbTNZNfw
HOxi2cWIpUEzWC/ZYpZm15wln2JT5lgbSMsaqwp1IQ7Vk5bITZSdY9CrtXuQXR5z
12rM+cB0RXuavZSXcLp+qwTnw1cj0HMjtlt1bEO+pc5AmS46qZ2kS+sKp6+Qe6FM
i+tb7AfaMjFgL74OT1+DANMqcpvE9WIIPYCSm3Z6zNh3JnjSRBBr3CWLJKsB+1oq
H50+Hv/5RHrAGGtdgfbBcTPwfDdVnni8QwCqiva8F4056Rf5PkU7ttKtkstZIRrb
B5D4NLvVp+5GhtlwzCnQbPYpcX9fVuiFmENyv4nruY7IKGgS0uRZcwHKowKwPtSx
zhAbx2aJcJwtB3R/VX2Ng3wmhaDxgtHOmNJWeAEdhJDjct+04ZrjBRxi0ichchR8
VIR0vLun32kBJNDsQ6D+4ml6NC4vKvWbw6qX6LfaiX9PH+AkBGX8YJhHZtsv9Onq
Pi0iWenCKapDg6Jy02vp3K9VUTFmA+tGNe/c9dkeYCAQXI0gcGS13t+5WaSajYQi
vPAKROpu3g19xmxzE5PTWcUOTWSX/+YUDUsbRZ0+yV6jZnQ+2YQDXfRww105Tpd5
aa/uiKp/NDEl9GIFcZjJJNCFNxR1dgPpPXV/6RxuYiGg8TgRGRdScGKG2IZ6Ji1N
bDSOO0wooErl8H63WsWpnDoe4ERxJ3MZzXKBuv1J6P/BDTu3vE2x0VB7YwcRKCrd
Bx8IPa+eaq4EtY70TYJX/waIkxdqPMB9AtfbDx/OJmtbH3xJz0uTJxX0uq6a5C36
pR8vhgCFewCW9oz3b7fOI7+tjUX0IcR0kIOUD6J19uXe1NwE9kBqJEeB8E6QYQ4+
GZZ3JOWYiil0dQLd65lHezLCzKUeAwY+xjzTCoR/qIdrCuryOjB7oTnxuWsEV0Rb
B17IEGfREAv9TX1kwTgT8C1Ou9ff2Z1SPRpkSx2ha9Q9rsusGhQ2JhNB3tpzZVed
SLPXi6HP1EiThcdTruD0pve9MjV2ACE2WlC224gSoHVLlNgEjsJVIh50wA1AUJx4
DVzNfeKcLJR8iOqREXuEztNg7j8nSKazg0IALNn8RHDIKaq9bm61dWeRARwi4444
szjKKePu4MS3530I+FYHvgf4H1zm8Je6jR8XRIMj9UH7BrIeMef2nbhSvrz5+G0R
4k4fHvYOBCVTrCx0aCnxgfRMyerFMR+qWEmAv4aHG0YLdKErVj0/Scmh8f+6U6fY
2SEI/z+6lbDL0H7xCdAWStnz5xY+wT92Kwn9O2D2RtjylajSijsIx+tvfOgmGUCX
l/mBxESmsrBJcP1Ii4JbqbNiSF3CYl8wzxNmvfKvW97LHLT0DtFILiZU9yUjx53q
KAtgfbnhwReNICvEAWdRYLR5QOsF3WQNNmKnjr1drDd5OrGFBJ3+R0Frg9hc9tBZ
Vjq8nwKmAzkcTpQymO/MlIhYP+mSG+J/srS36o4BXAR1BfcQkMZn8+kqxF7rxHMi
muy/9bvtgoLNRwXM+SCWQltGIjnBrlV0XeY9mq/rhYwe7ybsyyBAEaKAJot/BG2L
WlsFmTAqk4Vs8UBUnuFCNTdQZBNpOSPQaHqUHMbB000T0GVev2w1qrVkqaozSHRL
HjJg6sTbX8NfxcrBXgZMSw+kF/hjo9iTL3OWl9KoeebomrW4Hy6F0saiUmw5uZ3M
8udqoVpH01/VMucDQ59ISYS504vpljDS6KQPZEI4rjzR98iIYWup4YpZCkCwd4pV
9yXMYeg2FzW9eL83pdyY7f5LvigW7y3LavM2ZHgWpp5DI6a9k28samQ4n8U+Fswi
YZNw38m+I5obRILoDbIxJ4lsIPMQT7UJ2LZr1nIjePqEJ5SS+4v54OmC0t+hju4y
T+hRKoEyxOtE84SZMTrvzZyLkz86Tzy0Xm3gABOcp6plXZE/OrN2Ld3pGY5UUJm5
ZetKn7xfIHVJRwuH/JXZ5WTv5FH3F+GoAwhxJ82X9GMzk2sTGp8vRlprJ17k8MrW
T8JEb5dP+571G9TbjFbOUmqvflUsuVMLXcICaVcjfeZSnCb2muyv1OWYW923l7Iq
ufD531yCNfvMSMYtHpEnZAvIQcTneu+QhXwh9bcQYaLhGqFXnbmrXCH1CRLiKlOl
Xo9hfm5J7rYoOQLKSXDf+jnoT0vsL/1HCNz05EwujfcoKoiyA4u6RqJS/Mo4HuAP
bryoXSQ6KXFW6BfRjsXBZZ8F1ifVTdP46ePnq+K8aGxWvSTw9BSBT27UdbEE4qvC
mO5KMAwiXnW/uCU2RqLNzWuBjR7FW0OdjqNDsAB6Pu8eXR97G/3tGprnOK0aNBxp
oW55L/VYb7PdpUrdMtSA/6HqwewbwyiulJ+r3TTiyN1GluE9N4CIQtCfh0icsU9T
YCZY2NBedT1K28f35s1Gy4iNU55kbccdoD3y6hT8RtlDxUmaat3MCD1l6+lcSG08
Up8VQimpmsQFkg4MUWbrt64fHJRfUZyQ0ZXExHT+NqK8mt6pRaCktMBLHV8tlFLy
RrNSo2cFPVz4RwrsAC2I50Oet9UgzsBnpEp9YSBsy515EqCk/9pOaSpBytW6Z78a
3Hv066C9Hbsx/r1xpdDf/l3U/T4mCHNza//XAh0MIEWB6CA0ZSSEKHcUbauDvYUD
ooWbJJA+SCnRjUQYGm5KZ8H6XpF3jjjiQgICHseUtijIC0MMvX8c5eK0CAac+yAe
MWTpUWAAvygNJUf7AEvP/GFD5htaoK7rnHfdS1imPLaD/bsdTQy9mhZeXbybojo+
KW/WhHmXzNa57laspaeBZngaUZlejh+2AF9VzGEEJNu50Zr/qAddlwUaahXT1pm5
mHwmxI/nyMESuFravcggTVAXjBPOBeNZJc++PpnwjB7wrGPG1OWnl0V2LWyOcJbV
71OHYBYIoF1ggTl5TQ2YPHMUoXSzQmfsZzpGcP9JWMCUqrOu2IpYzwA6OPQiQ5jT
/zSIxNDMdjAAaR5uJAtw1m3Wq0UuBWJEyZTY0wS34XI0iF31u9ebMjuWdgoXbJZ9
DNrbMrDkxzONMOCeKlgEkuJis3sBf8DpGamU+fDKiHBnnMDJvc0miUlLpylYUhPJ
XAfNShSauhensmWbKgbetppQnldHhPBwIyYDE5LXr35y1zWuQbyW/0gyQRUwn0zk
suBG8wWAHPzXQ9nnla6edCaOahhshvX75FfVspOuxYNeGlYUQE7W2N+A7joywJfo
I7xoEG8dQGgz0E/eqiWLvYyfFJQAXUhMLi9wq1AKJ7DUFMHGfuv3y/Gto9GL/0lH
RVPXMNdBR0qOAOp1xE9ixIIkBJ/q9WE8HtcXxuq5HNk6mUeYYDlN7LFB11Yb+cvC
vSvUKje0SsD5dbHGtRPYZ9WjLb47cdqkqF6I3NwucWldjC/5Id/tQBgBzjzASiB8
rDEoj7pF6MeQ2LELGwZeueXZuRtkrxuC/p5+aqtXcHx+p/SBFjpxLChavIcqh/c4
qb9Hs9ExCc7nef1nEggcBYaA1BiaGMFdrJlXPHkZeW280i7/zyFDswiNevXSNyCe
U2XQz0H2aPHGnWtkyfLMyuC6cXMv0NwULDjPhSheeG2QjOiPCkBs71jn8FUWeP9l
qSiOyVZMNriZF2ssw2093CNxuLpXfmGWNUBHeHLYN5pb+X8Az9aqnOjvPmNRraSk
oDMeH32Sy9gWQmyndj70Dw/gyp/YHEMDm12IJ7kst1br2zUfUSigcWKtMWbZk48R
e/jMnmo0bskDuqc2gKeGJkMggzWvfwFroLNgfcdwXZPAa8itYoW4spjDwfLK9kS4
V7U8NBEX2qLs9lb+9HMawzARoy6qlcwZrgHKhPOJpAjo0RB12bgHoZdzaXnf2fBN
8/ObRzrnXA73pmXoBzXqKv1RbcwoS8aQLXmq51npu/JnvCXcvamgUYUnh8LVeKCt
BdChLv8Zlln2LzADRs8Dy+LbfSw7NWvtsq768c1r6hST1DdpDw+f8DjHLM6XMW2q
5gCpB7/17zs4b3wWhyDJo7Rz6zOh0uvxsloOUezK5RofHN3S8vBJoJgnG3fHEKBC
G2RDS7QLccR3NdtHw/+d3knmVNu3uiozZpT+ulL6uONcIWVqZoTVgHOWw7UqkfRE
ig5pF4hv7qmyDtPAHgYXpCP0muK4NXktA+SCHacv39wmpDPpPh25FrwQFwkl+nbQ
aVKaCChnrfONDFsBpFHmg75Uh08b5t/rgn+btOqcaNOdQ2ClGDOvv6gX9YB58qAh
ECGEGH/0cPQ8AFioRx7Z0bb0Bl/rWkVdAn/I7wHxDlZA9a/cp9La9KLfNdXUKJeX
B0+LyROIbBCwMVZ+HKcmiT8R0kphcckKsk84aiQZQlI18OvC/9egxXTnHcBuLjOW
MuP1Y4DMiYjEyWAqfl68oQg6UGPpM9hZk1A27mX60n7jUpgQCiKKzYzkzhIL1JE0
78cemSH+7agTi5J/PTlLrq0YCpoqAEyUo9qzU9iJqBbwWdtXItd120KXTXkyGO8+
4nTbWVEtwJhveQLAqltkp0rgWK0XY2ABsWovdtLkhWLsDuMqZ547yLvkKvyiL56A
wl0NK4nwTI8778+I+FvyJDV8jk0VMaJ4urbCXa5SWztgxKH/q4ucHZVis8f7HzCD
Wa4fpxq6tJUM2wUSOjx6sv7MMLE1V8WEPaVbZAE+4wflfMBVaHadjCV62sIrUQy9
iPEe7+PL/VBB++1uUbttT9iGXpctqbBnaQOlGsRLnKKXaVMNyJQlaWix+nKSrH6z
m8gN1gWuZ+FzjscgBTHyw0PixVd9JpuuJSKT9t+vVC1gRc8Q7QnB/zlbNOGw3Gnx
8EmmAJr8JOKCk8c0n3m9zdXkLsCJwIVWwKvH51Kiupnfrh91DblUfXV6ygsGiUH+
RVxIJOkZqJb9lfnhzgRxXa7sFEzOxb7I1s2HRh3VLVrulRF/Xjor5/p/c2UzCDax
aX7/9KrGEaAmJk05BSE514kL9bYo2mXBIjx5KhWY2q/KaGuhbayJ5FR/ixulBUY3
+TqdzQ1nnGfnv+wybeYfJONL3u2Rlv6Anpdavu8DomOW0x3DOE1UgznwjgxXj1gr
y5nQE76xnhxjs8yincUVJBZTaK9UxtmIt0Hp6YAJeHUn2QwPzIwZy+1vlC/Y0XXu
KkUXDjNlOCq/HmCnTbOgJz66qTsLO4Oq1PFAUw9nB6+D0uzWEkcFoXm6/Zgh53TH
/A1XmVUkwRT0JT3Ei0L8T9Lk2ZZ/v+/M4O6Ew4fKzlN7JBV2SvYIBmHLC+ch69YB
hc2MD4sqIIQlLxoC0V9O55wWdPW9f/5HBNCnfgUreIGrLEI0zdLs+lNafX7dqRwE
ul4VYO2gU1/54/e3wDaIo4JLTEbCMD4ud8m83k/oiSqm9GlO+GtSb2A0dZgeRQ7L
aXwpoxyg9kViGR0fdhkins1+uLb9pmMbTqskdyusitAJ1Wsh0CV4XnF9PoP+Xbyv
INgswZiWyM12uFSrvIOvxlSJ8YxgHRmaAYqnnn/2LRFmWzq+s3WiqOjObT4FjtAP
dzTdHQyEYFdsDIqwqR2iRi9qtYUyOwNgwxu9J3Q/7SpDtsYL4ORlR2j45iDSdXYh
ktTqsgq8Jcp7QsbeZrtxNvIOVKDmqDmeWase8qVuJ18o2v3KfQW0cbJPJW5E4BRT
iHQ8ZhRWx1SaegTi8DWGbW9k13PjosuWj0efOGIHpJMhAKAYhrNDG8q2RniC+6p0
hwYuxY+WcZXcxgpm+I29+Bwi1DuiDWPr+kYTkuX1WBjPzNdU4SqVqNY2AjcBp/zZ
foq9kvQMJ2bhskgWNcq2xC6XZkiC+IcgZ4j20rgnZdbz+7+JGqPwIZMzc7odRXPS
4enb8dJrsPf7Tw2Z8vbWl+zxvHrCntuivuTcjIw/X8ybJpHd4HZRZL7HxrOQjcNy
U9Nt1o8RQIlPYS1c5DbZnHEPa61hEEeMAqeMN7yeTJOmwwDM7ckL6dXwVNMeYTtT
95QNNkVnLNybEGyhg59/OoH1aXXnfEXM6JtA3SBUoy0XJ5gbjYU1lltuJ/Lipcvl
c+KSaX5SYVfI7p5Gfidw90SqH4fWppkAH6dO/k1fc6EJiioJwEx6eQuD1e8AvgrX
X3OYSeqleufpiZUqu0Lkj2cYwgbhEIZrMzbBCB2bi0NvUgXBDVkiSXeHzpGn6gJ/
aPAtJq830FWkL2Pgzhr/xc5epCxS3NoGOnppAWqxtXhq9x51aXs4JRnHqRYcNV4m
2x3cY77mLYLw8oqrsyTy83X0SLVPqwpUnzXH1CUZmbOiBZ73Ro5xpsvcf2qrgpFi
R7TS9VsabbUyji1Wj2AUsoHUuKZhbVpJxrHQ3o0DPHn8tgtbY2u6vNmV69t4M0g0
ou6rxvULO2m1s4HoPsmKM+kzRFcoQ9l7LcdCz86bep2/3xAFkXcYRkl/QKqTU0ev
zqXoEIjFMsKdK6EbX7y0Gs12PUImNkxIa9YmyM5xJVv6w0NhWP+a7X8xHJCZiM1P
1bPvfVpGNLQEvtiPdTkpHPkgPCQkjO63raA4Wzyo858wJP6YxF6WTLO2VTtmKDRd
dfcNHTOsHxNixmZImQT7o4F0XZJ+1/6UHrH7UjBRWARRbAYLT58asR1IsQcREGBU
bF5tjqh4ubU5FBJrD4E8b0+f/Zl8j/afoNy4WcYysti6JmEJoVqu/YNApgTLi/x6
IOqhchNyhKVz5tk8kllSGW9ky3LH1JqDU+GiTaV1CRGW5rbyvBNZ4naiyjJpT1Kh
x/+gQiYKKN1MIOPfUx5dWIFn27v3eavQSGqQ24gmEKz7iWwAptW7PYK4WAZBfksL
PyDbpuX0NpTfbVGkh/lzI9yqHIoIwTv1AGWdm0gFM5phKaI7hyBpykyP4IEynPsR
N+3lrjHzJkUdG9KyMz2ojk/0JA1oSFj5J4UH1ACOnXOdbda+OjQaA4GOqe/mj9fw
MFYWU3dZfGSncWld1Tf1jMo/dvoGam7kZALT//Ls7y2JY0xEPl8exPg3/hbiZwS9
0Zf75nt91sKDtHa73xul1UCrddhMgObTR0TOuZxCCB7XSNYnTOCZq0n3mNSWxFNR
A7gYr147aoIaN3A5BQuhoAY+Z1tX+vqJE7ahHBx8caU8UyxfGKA5SQSSlYbgfCRy
YINIRInYIJqbZSn0CjdJBhM1aUOiVFkJ4KmVvknMrJQXkBW6WdPVfLC8Duh4JLt/
eBuh76BedTaf/KrAGIebe3LZ06ogfVFyTGlS9oLrxos00kVtbyxf3rtD/v94Jufo
Psiqaq0Kgec6t4YgN1GDpe/E450qRZ233xqVBllSduAUIVEcMxuyZ/On9buu0aHm
Nb07ZR+3+IiLbFa+hZC2c/zGjA5uQXrHRLWiHxOCMp7n5VCea2+y5YYGYxwqzNP4
TPJpRBvX6OjHqhZQAfDO9RDJ9jAz5vD2jTJIe8Qxbk21k/hCtw5Q+ARUMEvlUkQv
rKTB/HehEGlpQksYjaIYLRbuMUYnYnfvlEnh9826O2qgMX49Rioy8K/n5vmBTtb/
eNpX4yfRR0rCnqaOHTH+MpwNkvH2OpyYrG6IoB14VKCF5EaLfc3eyrJN3Q31craz
7vTM1TRZIhSQ44F3p9qXeMjVo88EQ91wk8U+NaWnkryA3e5nVdE/o6PMnILymxRv
GSZu3LKfEopIyUxB9F/IDfVe1vQ7rL4K9Q+h97R6fPb/b1VqiqxSEIzoOqBU11tO
Fz/FvPluyN8WOGbiNO1M8qWs14hlH8quvxKowReFPKGG6a/k5WpIBVzccPKFKYEt
0/Cf666/CqYLphNfJ8bKkQiCyiNneIGj/l0iVSbv+dVqBRghBzJhAcBtGLIVrQ3r
MqoHmzu4BV+ztcWitObbUz6kzoZDUL3upntdmTzi0L4kJIqbQp40bHOCy0HmRlim
0LPK0qlRniKWDp0PsdNsgQ/iied+7zgPGYYFekAwd5NYPpukEl2nZuZAL3VuPIjM
ybMt2HF7hJOzhRfkKmFL5QY+EHSCfPZrFcnFaf4Z0lrBBlSZVWm6p7quH662PjQg
2UuSehyT0hYEl2eD36JGUPts0Y0FqmhZPijgzAE/xc5SwISSzSZ4QapYrelt5FoX
XLD1uK7rkTLg3d5I/h6jwo55nKVrRhzjE1dH2murleW1m7KiM1UDAl0cgWZmanOM
ZozPfKyaBYwZBG4fNiOvRghHHKdTwB68bPiVWPG4aPdBihiKnXabqWCkKsN1qxYc
mYnS86P9T3OfLWp6zZILd1ptqb7fF6i0zwaTchfWJHpWFibAAK0yuRGiX4VMaVOq
Niap87BCFl3Zc7nxaN7PofUoc1+p5zF1DJ1fp0z5oArUxV8BRM5VnXHtZYO5kOIv
dmG7yQRuJbkwPm3HofrIFsEQ06jAGKLaNZllMwhzaEMbk6fGL0ULxFFHkZNvDOzt
Mu+sXrpA6ITrpKedxr6Uzy8/ZZKLlwsKsZTy1exmaUI53zcGWK4Eps1HoAW/BFtK
Tiu1VfxoNFFOOR3NE57EgvMCOt8m9d6VEHpKzakpcYfI8o2TGmuRcKGRcGXHPDkN
HLliwzW7XTajOBCiokKc7yV5nf5zM2YbgTqGYX/tVT6a8nDfUz1V5sdIFRptde0T
Ogw2hrOi4ZpOz2jGtT/4Ni85skXD1E+KY4NVT5+HYzlT+gR9RByb1sxwgaO+g+fC
7llM3GQdO5zOxevNfzPSRUkVUIbcSe1FilCkyQXtJvhiQX60fzZ6V3mC/THsrKFH
XrdZaUwr3QyluRNF5RV0I/fqIqw7npfMZfF/g/s243yEOxXsxf1v8FQeAlTO3eUR
egFDvQ3Yf5RFC8EvH6ZfqBbj4CvgPyG5+DmWpFY4WRvQyUgSffCnSg14xbQwkEcA
LkIKXn0CgegC6sGZyRQDngXU0cj7k8d09zgxCZDkem5bXb+iv6crRxx/krKVIzdG
q5lqiZIVFuGx+wOZkv+Yeo8ca5bJyVw3OHjp7dl0afwGjXD6yPIazE9TJrYuL5MT
3Z6roeJwnD7oX0Ir8JsdMoGGzUpTlOH0RHDEShU/0L3j8drW2sjd0UUYIIozqycD
d+03kt9rlxgPZJWjOeDE87DmEZka6//ltEt4aQchaughYQNKQ3dhA9liHwE8tIok
DpOp6AtzqwE29p33RR5G1HMLxc1vMhuU3a4y1G8LI36OoPi0Jt0DXiEE1ZuljV+0
jG8IHSzaMWCIfT3AzeSWY/U0t5i8XKKFEINQjBZTvCwiVqd1csCYrxVlqRFLi4vQ
asjVuCTsM/khWswXEntizoS7z5JhZ3Ntx/1zi1VLNx2vEIr454IxyAlfMpo/Idf7
nFEGS7pB04TYprvdPC+PqlKsZ4P3q1FpMUPhaOd7w4fenM0KCgdZ1Q+MXQD1yuxF
xarnw4bn3pbuMGuvmvXuBOLJNZs9kDwLdAgoWUfMeKmJr4ui/h35WrugbpsZnVK5
QOh2hZ+mO5TQY3CxdKBjYaJ4lYQgd7dl9mZAxk7GXtIWWvBZlVC/TvN5NFuT+wAn
tCg3qYQIzl0DyvDEpzqCX3ICST5nP1bAXP6/VR7B50ZFuTAfydlMxlX4z2X9jeL5
nxMhbgIcrDVQ2v//RkEO/KEMuz4+ZM68kjz6S/+NGVTG6GO2ojPaHg3sv7bfXFD+
x+s9qYX4MiX31hweA9F4LSBgSX+2rUzoLvSVFICSUKbARF6986pAYnd4AYGocFwF
a04HKyi8fJSQxtuIkM8qTcTKMGKDXzlHAViOuF/hdVA7bxMjwI+4vNsNsA57DTsv
VLWUN0oCw9JQauZzESGNmLJCd1zQNfmOrh7uSe2ruT9+EIGT18SQ05XKKhcnOyxs
OiRhb7OsFJP2R/caW2uLiR2Wtcari/GnszGsIBM6JTmHwOPa0iqlY67cinP3uUxr
F7OxgHu2NMp6ecixJCG2QDWXxFT2odmpekhjo1MmFOowaxmTR4friryXt0QS5Gbd
t8+G9kACKvSG9Y/YvV6h57aeb4ZeV6g+3HCozmNXF4kXHbUKF9MhrGOsW8s6PLjo
ejzppQf8r0UH3e60KO1frwbEuo21SRnwJqAQTEY6whUWTth1uLV/MRggdzZTIyC8
Ht6mRBYtkg+MgAjTdgAY72Ny5qTtLDbK2hfIOYwHekyzUQaBv8ucZwN3g4mqIHKc
7QRp0dvkzYWQPCLAhNM4tVZdlkGeHhXkJMoSnRc4K4SvWRiMUyiCk8nLr7SbSRD9
9pmUhwu+v3/Q5VsGYuo5CKp4hxgjQ4pKVnzH5ZtJm7qccASdIAPbkso1i8okaPII
pnIIJLnX4RWM4itId+oOOS69pTt1r3k02yR5Mj6fGIz7mpX5LMcvCRazWy1wGniN
mO+O4TSTqltlwsK41cP9bQhtGqxt15/aF9TjzD02rSiLUmYxsaBv2gPVftx05pgk
I9mS0T0Ciq71xZJwynxWc3QXd0Qykpz7HghpPj4aSyLN7wo7Op5tHm4xguBJKYO9
ptyrnzLEuOmfKhWLCZOi1QSa8eHSmM/ZrRxZv3K/KmBWGR19Iw8EDaAegcgyZ8fS
XyL4lGAl1DPxMoumQw2LjsyFdsbfQ00Soegne3lwjIRiRdqtiQy3jNNWz3G47uR2
r2SQxoIPiO5u+z+aNgB3mR6U4vx73fmO9S9FVGRhY98zMENwzIaHbQ/EwyZeohmL
7IuxJFL1ie1m+qc7YYHnwmBHRW3ZTjsJSIdWEos1svBirBNJYXv7Is8rNuuxUex6
Afd8kez/UPC0g3FANaHcLtLf92y/OzftVBvVWXzeUOljZ9+5Ht/bKE6RoU6j+RnK
tRi3hYxUORUcWsNBQ9/EiJ8F05PK59wXfRLzT7FA7wExw0MZcd7E1ZYleUGxYSxm
rhaAdGNv/I3dR7ZCAFOdJ8ozHPxAtie/HlU66YRIsk0bDt3i4mvrof+ayCXDl7LV
lkkW54QXMKCXDY6E8YbqDegv/BLZrNCyR4H1eAY+U+IVlnWHrzAdPyHQ2iFG6RP6
FrLFsyRoXhlUQVWOiW69L9Ir965QYHcGD732oW09nyQnWvj8b8fZkD8SLwCyxLjT
5ALKnuxMFlZc3bLOiqZ+fzORjxVfsUJcfI7S7CItaLVslEwe2KNbQ2XQ+LpVLK1E
6ZtUE/dQWDZ36g0Wm83VFpa6BHYPiFmbaFOWTjSfXe/yywpgFpkp0pumak5D4KC4
JcSVDIZdfgcOqF9tme0P/KHbL6UMGK7ZNrkZBQaxKbYnF42+yfcyK6MIrjcS/VlX
6t42Bfjle7pVMGhHZfsQopxF+cpIKQDuScMmYdUYAbzd+ftXh8DnBYcxNoXcdvje
G3x8pZybWgkdIwyLIYLYCWn4dvL+qy0FCX2DwFKcenRLsc/DrTD/Zx+kz8tvrFKU
G6QN+vbegFHEOsNQP02Edk/9qdRdziOxUgVDIQJR0UAAB2Fxqh80poAdUnzsdHUe
KvBZYd80CHn4/AFna00ajQUdt+8gUBkioXUT0m0lfmlT079laKcXrrDFRMd7cPDA
aoW90Ybe/D4YEsJD2EuquwAGyZzYrCNSxlMFGq83RDPy6CBKB7OP5Gj+H/vVwWoJ
Pe4fiuRjkD+ZNwhwvqn3XwMOO94t2dHwbobk2vEVYLOEpk0/mUMH0Dhc1e3g/Ig3
6EaxglKFxaFuYg8AlcijB+Y6ZNYeqzMXo5m6wby4OxFCebIzh3VCCyIO6cfKDRMv
KREHSa3AFfP5/NdtUHsnw6/cmEabwtrFv05ZBizWRo2DVc3EggNWHgIMnLqBjzW2
EUliOdK57IWxdh17xDQqd0vyjMMF9U7BKYr5k8duHsJz280sbb9FxnGzgmuFK8ld
YqvIULa5AMHvgcEK3MudK+Lh+1t3Sj13mm/O8GM7TKI9HpDERun7CIV9Gf21rRp3
R556vElmZubbKqjvHe1Hzqrm3ki1RtcQq2Mni3Q6ne4BJeWkg+iM1rR/NYCUrMqP
T/R6DmDUBSjbZp5EVyfzDG1WUXIhW7ULXjQoP6JTVq/4q7CAzawFryrTkbd8jtdS
UDZVRdAFnOoI/DtHj+M1iWUUG/9CJmUijj/YU9ex1ZmJvxLGp3ij9cIgkS7/cHBA
5b0ppTehp8ITXJfgIh9y2uQc5LlTYGTDxGwBStGehVu4w8Vvhx66iZkP1aGhv6xG
nBO/QDMEfCBP2DNbBEPua60K/Y8NFip99W+VXhP3Uu+y7CN3Hg7WyXdu+6ycuUyG
uNjn/+reHsg6DsS2Ve7gK+s0o5jAI5oSopYP78uyxA3fM6P6BYjBApDfbOjIqWcd
QfGrG+0KE3rsGBEEBtQ8hp4tVoPiyLrE7Yu3buFGtbP6D8JnQO3UG2+g67SrZrg6
1r3qxMw7BjKQ/BsCNwE8punLKQG5s/eVl4Ezwypy8DSit14lmkkpAyrJxDb/gBe6
aqEeX9m983FtZDS6tJMGMO+IXBqYfVUBG/NTzL5vSmDnszC0fhjzMwKFKlFS3I7d
BjCRlvmUHElHw6xXPsETLNR5O5Z20piPwTx3CrQqyAG3wNdqKQ6APTooye1PJfbs
R+msMERhCAFGcrcyJT878JGbYwQIYWkTP8s5u/wbKxMA5+LTs0MJLenA41YAuOLE
dFScjCs3xYkCet798W1w/lYxMa7joaCuHU+luBwyt9+rZcRpO/xCC20hsyL5YYGC
LYRHLg135EL33y57sciT6YVRkiyhXm3LFtPw4wwcQfQKA8ji2ohktVFemOGGIA+h
oIsI12cfhXkMwQpP4B9PlNJU42+B86kKeyQKherbZe6MhXmc4rWESwx3XKRaHv6c
pZWbsY7x2xsYDwjhSpymeUFKvsOvdnbqPHigUDoOvdWsaJ0HmoYHnRdU4u3h6Igj
wZe8Y0bjBzw6ELhEAm1QVzxa/c7d0Q+yyxBOALKS2Ow58gVh4y7MXeNMgeuODJ9d
1+iD6yXyINkTByeHZUX/ytX8a71/hcA3hIVXCehxH7zJRTdSJkNf/RNwkgoQ24Bb
jnidoCe9zJFvmZ8oiC5ZOl4QBsVmSsAsEOTPoniWMXodxL3UytuHUZqDF7Y1YLAo
wrzD1bXBhfY1hyRWaZWjfNF1pPBXwBupjIqGYMzuhGhOCHnsi5ccykckO49cbAlz
0SUO1L54MtCw3TPl1CIppeDDBtchXMIf9VmBjhotI9kZvzl4USEs7GfAfQEv6yMv
pd0y9PxKe6itwBr1QCdFzbQR2t9zc/DalNshJ9Q04Sjzpl26G/EYAkMvOmrP03FO
4dVdf96kpAZAIKu+hX3fU99Z0HboHwHq9Dpu/Cuof/UjVxl8ez+2mGdf+MGBbhOJ
SHaD8ECFDau9X3SaLinKd+G8iZY1OiLUzOOtQ78xzkTbejE7Rl3j35EoEkdTRJx3
SWQVsE2zYF8GC6b5S93+zUzxhrMgH0k7WlMYjEr2tDKuB6j984T2httnEncra+Kx
fcAwHIhzF6OU3+JdDmjAZSbDA5o8btm15j2ldINg4knMCLLmFvvqfVwKC/SFcpx0
D3Zcyz2hTMfGeLfQP0D9INpVYPUSS8tab/f0LMPq5s6LQCRYLLue8d1LSFPE08WN
7I102jGho8VPnYFnoPJEgpFC+kKlZsz0YexEz7qBwmElpiB5+rUQl2qOda+YQUBV
XrJ44Y+gd28zMH1rs5T+EMihFOwpBkQ5t1x8iFKuVc4UOO9eU9PmRdT5rgxRx0GD
zWlLtSiSmcEtBR3SOixHNeeV+PQPRqcW4vf8IFptXYKmILTmbl44k+wdYE6dqiwd
fnJOprqkkcKSi+9/6QOWJ6VdsogPi3KLPemvHFKR7EURHaZjv5HcXyRw/TMUKTIF
+HgBiTenh6RRFNZLJ5zlVPcRqYE/h5TNLNw6MYPLfPMN9dQOA1yYdXxoiB0xvTjD
p4fWpiqzz6XAXXaSae4MN+poJXo3IUm7eq/AGc1rppWP6ozdwd7SkLS/MtOebxL/
zk1DCBACA7zGaLvq6fdyDCYlwuEMzu0rE5n3cYv6OUh2f18vyMBV6weklrPn/ubr
UxkAnuPwrZD/OrPC5UjRA/rOHsYHVoOEHEafRf8O9P8FGNNHbzV6cqxAjKnSm+rp
ZEx+H00sY3AioITorFd709x6HqRcD+Ih/kUNFUKkaGDV+ne/24paJa7CdJdXBwaG
ITiElaLdPW4GXQyNADAcIAceZ/aogSVbAb8LhNXgCzKW3YBKFFkY7yfFV5HJ6QFk
kGrGZNUp9s4Lov9K7GNpEdqdUKhz7BwSYd9XGJrqXZbvzreaBdQ0gOucRY2Mhmi/
I6G95WLM/rgX2aXsvVQl5V6jXuY/MPTiP+1YR4IuGYSnSsEMv9KIWYZgBoM3Xmo3
6IIQ5SVID2PrIEvhFpyZVHZVpeXpogwQBeNtWFiQSxVvXbIOxeNidByNS1WFnjaj
+riIV4NWGBiaLPMCpOJVqnqk7xzvDofaFIOcCj4ASi7IKVHsCN/fGsM6oIZK/Sii
Mv0Fti9L8fZdZFLN5RGupXJcxnCVei4u4iQ9aXaBkEjYiAFxZ/QBVSPuwDpc0Ntr
V1dXVmuDhIV3YjNHqS205U4Q4UpYFcfYQhVdEmFQZCjJj11SpnLY+GrbvOdZdv0I
tCbcvxdoIBVmPfxFzyYZnbsoYJimfJzrsEV1Pkz4TnhvleWWlV5eDkl74wk3hGkd
R/NBvZ6zb0OcYZUUlKlh+xflE9bnAGJmtsynnuX8Kis0Uzqg+opAWMzBgW7d7che
U+Prd0rnn/p3PVXj37fW27clQwySVo9pIi7/Uhl/dUswfzVaU2kmqwSjW2NLhxkO
lePCbaOCe6uPZwfZQSgjqCA4/5B5JIxJV7K55WlL1LWl7OSU27ucA17s8v+Y6FSo
EJn02bENZaSVxZc+AdENv4QRRXkHhgfuYPD0gpNbHNrAbspn3OhDdSHCTFmC+tb/
YQrQE4gjpn3M42XcAe0qf5zM+/R5lOX/1H5L//GQFZL8YO+twLEa6gcDzXHFKc61
to9yfghZ+Bv91ZWz26uR7QNwIuuRHsbf137TMS8TfhGsa9NCsdTb8PPptd2rvoNO
W35XY9HWdwkqyxjOeD4r09LgkuKQW2RO5PTf2fj6aeDtek7plGL3UtCAOXXr7tFp
jhS42w+1HvxN1JRWVYIJk4aKE7KHBZkF8nMlELaGxpvp5a5z5XePxPUSWAyp27Fj
dKBu7ELBx88TaiEm6IiTeDXhKqC52RlsKC5l+ThTWfuilqS+rvc78j46tW5hwbRX
tGBdu+u9rauHXqHKB5TXoX0EyroG3U48059S1hgY5GWI/Mdpm2EeE3z7fiGMEng5
7rHZeHlaVzyOrylvu4zJDVUFJPWSfdCVTuEHYNr+50E0v2tEhP8cwmuZNIzFnq3f
KZTn2L7akN4eansNyQNxHhehJhAqEhnov+CU1Ew3TbnP20D413VrC7GmyAljJDFg
HKoO0nW71CkrVGPSx2/6Sqfw+sWQvKKkjXF8BXrc29riT+GBDnjSkSm+XGdlEzM6
pClO1LKHdf5Q06fhvLw7oOjO284B8VlNTFciBz9V3rwWb5YqcPpTkhIF6io0HVAm
2Km4xBzJ5h2HzUe5bZCaT13oUStsrkcQ56gDgHNcI/VLat58rEc0Qt7Qm318HpsH
0jJpEhyvpoBINJwcduYQGb5YN3l7m3GUswfKHbDVCXRIGQkTgy2Bj+7hYMzBix/9
7T79bsfC3JK39I1OjyZzEGQFmjI0+hAGHdfGgh003VDZyIxFvZZcwYfWnRQSVTLr
Jrnrs2OoPkv3uo6vKxFgeY9UFvtRWyzWg8khCH+UqbTWEGy7+7p9tLRwQXI+ObMt
RfPniVNt+dmhAzD2UE8KL407FnyZXLQ9/hNQfWEq/trCoX3Wbdu5XvUedkmgYanh
86nnMRQHpjphcoFAj2oQF3/1igj0JR5qeiH4wMfa2xDkF2sDX1rBQAD3BGRPndOf
uALJI8g7O5WBy+fKtti08xKSfH81QFtUd5FBdMjHTlvm2473vP6hgGJ0L8w/Frel
AbktOc7rYTgNW1nlJEmpcVU049GeBdQld654gqcFUzplhZ8JRbjOTDht86LAG3rN
LZa3Mzu4URfrtIKR+wbBJJ2Un8z6OT+kMQHMFAk0gb5Y9R/SxXHFSZFwuTfdshJG
fknPQW8WDeHaYscXOkAANk5a5NSjgriSmvl39CQKrJKskUZf5w9AW9CbrmDlI4mV
zaqa5S6n/YVCbcE06sZYFuh8n1V+639Fa0IImG2ZQxSVlRm//M90wzTqSsr/oB0K
re1zN7dqII6IW9ILzId4/0dmJYJVXz++P/p8KLQm1ZpTSOXTF5AMdwDC14sRit4C
p1YE5JaFTGbwCNYW6P2qvDNsucpPTbgL1gpQ3hxSa6kadR4OW8VhyBUFaVGfdUKX
cCJEh5ejCZ9Yba4lgmQEveXsKOvPv2MWgWP9ny9AGxXuVSphhHPTpJv3VD/5XUM4
f2G3mJYAKTjOrhckx+jmUqi6caQOn6ByrECl8UVmA86BmuCYOyW4T4BiCclOqC6Y
jrDPPLJGKLb1PmrmmEh65IXB2kt9lJM0HE9BMr7GXNIRq0duNoVuYdV8BZGAlTpe
wrh7Fvh0mRlV1rhnGj61L6efoRILKSTqr/v0YTWt9bkOrwP/dtdOA0PXrCqOkRuk
ujiQJELHGPQZ0gMFYmJgz7Awz0UZjG0GlHE+pNFGC92KvhDBKw83y4bhFMJLFpfZ
wQo/WpxEQ8kadV6L2wwxAbl0ZNrH61qq6xpQ2W3o5yysy+DISe5ZE999k+pqjLjm
PSxNzpihSSqjerVhN+B1JnlAbbTovn3k1nRzAlsrmTZU/NV8bsy+9sjuC2ynI75F
qUgykI3PjMGtvVkXSP+fBU+QcxDF3+M1J0lOCzIvhz2cwQrRuuAvGjzwdT7kLx1u
QvMkJtLxoz2+HW2cDceb1QSoDriSyxk6+pKq7OT/4ZGHLUrqnK+o1P6BKwBFwuLe
RN2m3O+Y+SptHHATlLo3Wmbh69uX/WBtwdee619pfLThnvqEixqA6X7ssBnk8Xyg
vklK3gr2+opYkP4WOskSJvkI1XQNL2RBeltCh8dHtjVUYWitCLpm2kXmutpP592V
RC0XIMSlWiOMaMiVibKxPiXD1HPvg0BwZHZLy5Vmqq2bIhlmbwNQsihk+F//rc93
Bb9x904tHLbSBaw53CtEFul25X7cWUuq1nWjESHR4D3TlysAqGCVtZR8wZR9G0Cj
BT7z1twB/t6l2ArjGXjzJyCAFtc8GlxevvOhseUW0UqgL0aL5ZbWF/6mBJ4I5zo8
2McXujK4Eg5ky3BDrv4uEOsn4ImV8iYBZm9Q24Z4TA79GuC4xyoRAHnFikkXFDYO
eS4RQZJhXqcILubwoWPhULyuXCBcvvpVH0UAqaK8DeNzbI+k8Tei/kNCdfkbJi6Z
HA1bcPXDW/Pbs8S8pR+us8/FVFid/X2Jf6J9Up3200Ypvinrd5mUxEApT4iY6Jly
5G+PHmY/DbHumwz5gJrxLJeSbhxgBMBgnyeY7jfbPwHqSxLtFSMZk/vO3M/YGPhT
m4ypuIMNH6dHq68xhJhPqQKHzWkAc8/Bl0B2eqhpU84xAidfJ6HK5uOofFZmwuEj
/n+ruqBTJTHm/w/3jeTYBU/z3xlZNdaCos5ayrF2sFzr9Yte8kVRGiVJ58hUi6cP
dES4At6uATYB6S98DJUGzwIFOfqr06Zo84iPMl6SAzA87pb7pYX5y8RJtTrXJ3bI
l62cdh8VEwjHa8K+J9+am+5xgSEdKmtCZ+m5g/ulifLV1ek9iQBlV7JO3/bcbK1o
aMa2NMmGlAxYDTCq51iVBEorZdFXT/P2Xg0PPCNDiXbdktQtBsqkRAwjsuy2izjo
68ubC7lOr/TQpx7mg+cMOTr99UbuAPSS4PfZ3zkpc3Xy9nh/UMrEJ7Baq6R/Fguy
A7MLJgWEoOKBVEO+elz0Jz/OPm2u4Vxg/N/gMTfr2kJyWSYMQAdyMEoAvsYniQ/4
Oeby8MbIj7SR5pNge3cbipnPpKgs+dYBvW3PBGV2GUsts5st7YX37IGjRPXuseaa
zFI7zlnKu+mdIIC8X561BN0HGAi1fUPcheQwxGSiLO1vrMFjvmqGpWui3QXBK15v
46QZMugrfWkrILyCKueHm4WqpgEMIUgfTKlxH+HzNXZnsJm7aDB6HlZRk7nwsKtQ
46vHCJ/5jes9hOZjtT6tR7HUePTGrOhbFIBIeYC1WV/cdw/ZWy9ZPTJpEuJgeZ0E
q6SE1lG/cyAWippTyvIcaSibEMNh/PTIHzPWwN2cwu3F6YOfsySHfYVspQ/NPYeK
HIBrDohWrG3ZL1xnAwOELTSMxyixgH2SvI+r4d9g6FXv386MQLnWeexRk2jk7Ryy
QhEb3xQpAA150AO1gxEqP+pFWpRy+qaVYvFHttG2+xEoyQEdOSRylSOHEB3z9i5+
NMYK9qjoBeHdpkFm6ssuGinJV38nkvQG6oLmpLUCMmIM8YHoneHVTzbHLFpdOsNs
7F/+dU6suB4Rr+uZENibTQYKQ5OPrWMq5FaCQ9QFIdaMYlbhfJzwVS2ITGCJh6ov
FGu96GZ3tlhbxE9FTHzIcpsuG1wGaEOsJSKbtJt2SBplVGufyjvEpD2vpEmAMr3Y
Hezd5Q2PTmU67K/qj/0//SoIKn9TpVeDRAPpMK+usm+6OV+Fr1wZSDaCD9+uDaIu
n+L8UYwt6JIESH2cj6BwFdSYQiJ0RJ9tDNXzpIDh0lt9rIRucaeajd5H70XumaZf
8noel7EmFPu93Q7e0NMB6EDotG9weQkzsw0lUtn4zCBE228EjKN4iKX9UDz2zc0E
Ke60beidTw1ONJ7gYOWlZ5Ja1X6lDTw6U4khFrbOUGaFOLp6EsjmxGIAv6cezECm
it4sevctU+gExWMOQy1DX+BF8/N+qccpm1rxuzuP17UtAJLQoPTuqJB36H7ilj5F
G5v1Utj9w3/TJrQkitUIUDXxoGCyf9QLwWRFKYUqkMv46Y/5KiEBUqe1Nt69Leun
ExHA0Jv6F2xU2vnuvQibtQoMTWo4XaNNhEeEWZzg4oYyDB9cPFV04piga4NVk3Hz
woktZV0ABC6leGP9ap3NIhu+asOg+M4oudcHnZ3hjZE/SkCWCQoYCAfqTMs8c3m4
cWrcAh8jJiFI2Tt0k4LI+u3V3d1Ae0FUj3ka+rKPppdLqZ1o6k225H+UBYCcIivN
UspHrLxyfKql+T2uQK5W6IcYSz5ZMQQwQ0ABlR0ymA+NWm1M44MXMCuBePOscp7H
QZifhWy5TEIrOAbOIICIXeem/mbkmlGlkhk0eT5a1u3WQoJyR0fQZgAIf0RLJXdB
8cqdD6HulRz2yADctgVvVjdyM/bUzlK5xB98QrJPrXtkPAPw6Kktz4SWflLq/nOM
UMcC9LCP+rz+gFYIE6nIEwFDQpeORgIPNC/1YHSL5QkhssnaQL4lFgIAaKVubueC
h0mZt++bnP+0H11YWiKQdkSSuUkEqHjGAx3kPncMVsdNyP/ok/VAbz79rTjxYPTI
nd2K9yV9mEN/q+GSh9ALL0KmcXleV6reIHHkKt3fpMGKNo9r+hRJnEaw3AZeUSuS
yvbcA8XL10RRmLQinTrtEGSgUirl7xanp41JtOVpn1ntEdOY+EK4WCjyWxvniGeT
UuQS351FOuxoYxIBjgumgNQT7br1juc7zbu7H9YeTkKMdiwVpT2zG4dzMh0oS/QF
4L6RgJV+kPRoN8PhAQRHWdxkR2trFvSg8LSC1DRSq/jpdcwWr2De8iD/zGYe/Y3s
kVVca+/myxvzMBKGFAfLrZuh98X2CakIRjpoMre/97VeKWcG4Kzl//LEhclLjLZI
dZ4V4S2sAdaCpqWRxM/5z9O7nWZV4ZiBETIOki2fErLz9vsPK/Vdh2rXqHaevC6F
4UnD4d/bileAXoPqEsb22MFmD1/bkvYn2lW4x4S0ejX2FQsNDiTjrmUWt9ENRwO0
DCUHLdIkykIgKJX99H+uKU8goBMttOZHf4zeHwdZvVujMjBuK3BAjgtJornay2xd
VT45n4cO9G0n1pQsn9Ds5hNNABH3iqfLstARECDHHJkBkrbzfkzXIXipCemzpQFR
S72neM61Vk3QGzbmhLuXmSFg3Zvo4uNMsgmBrYMpe/yj/WWC66OUpwJnchxo3NzQ
ddS+00cqfERotCB8znhy/5730vSjIe48gKJCEDX/Jq/62xRy2Om+xEN5Cr7FymsO
Aij+2mMQU/2sij/alXH0YcrvfSFxz+m6NlID+rsybCF7XZjabDTsfY+d72Y5leBQ
sWUU9P14bHZzCN4RGW676pRpSq1sC52dcOcol0LvL1HbVCs/vQQWAn3Cf7B3vDRy
lPP9v73g6U9BAjHFPQ+/Ez09MWdJ6qzmJ3kmYlfGA09U8fJe5W7yQgVWTI2Fv7/7
pJAj5jZBa8y1O0yAnG1bqu1vxL5es6uPgack0ORTuW5qm+/gpP2dFfQ2fdsfeuaS
Htztn3hI3qqd6GHuGwP0s+S4xF1HUBz4ONpbQpBJy66ND4wmQz+HNDf1cfjZyutY
Hx1S8oHJOcujvbWmmO5YE2tMIWWmZN1fYfupRzoj38iuez3ovYpfL2IPRERMH2vo
nlmQ6aWVAzhzXz6JJhPMpZ57OI62z5XSAda0dU1kEsYdXbyOp4nsLIV+ytOI6eTw
6f6hnSTu3yei58aZAwFgcB9ZtQ/p34ArozMHXBAPQZcpFe00szdTXeNXhUuQv0tb
18/HUZn8HqHEkz+nbw9GyfAPLmYq+L4CpEfeZ9PXFcTuL8fwLHkbgkgavWrzg5Rn
SOT505Q0SkFAGeQzXoIyYqg7tpHqub//ds2t4FvWwZ3OCzZcI3XyoPkCFWLNjJtx
S9C5zT1/jdhdoFJXwXQVvIUIj3gIRWgR06EK/ACrJ34eshjhi+roM7lvASYQH+yE
TgieCs8FnPiyehzQmWVInHlZh143iKb2fvgjWAjAAyqrTs5R/jg41iZO0fn0yWEZ
GHd0uqyjoZSDBgDZpJ/950ydboqUcBCy8HY39lNtmLRdvb8XI2nbZdTUKpOfd5n1
TtorZtwlGyHTHRvBUDkraYlSBM78WD97BPMGelMRMlyQ8C+wpdmWf11N2B22YO3U
4vzSp4YvCGVV9MwTSb5x+IpqC4KLA90FOGzDFmCyjG/A/uJZQuBRn8QDhetogY5V
kFiN3GxeIu7/pVhNMePMye4OxgvRv6QtRpg61SkOxacxA9Wvy4neiB87Z1MeD6lX
MGZCcl10HtC8+Mq6g/4EX3vxBTCIDGuJ4dHBgJItWXlv6KfhwzrU64yKlYkvEEq5
NlKtJCAjhgnUX2Y0RQE1JvrqcnCI068yt0nZVkEPJkQhh7P4OJUlJk5XFu7J8/01
uNYnKmQD8IbrDudGf4RGtzXEgGR83J4qOwDklQyrfDIjE+pjmHGM8UuLJrNUR8il
xFP7HbAgyy54rAUoYu74jwmQ4dWfFanPJYJku0cY9E3pS5LGwJ4nwPpGbzd8c8Ep
0ohmMstH+WEj8EOksBE6jEFwPanoqomeU9AYpoMiTR5JcERjichLLfXHxclACS9i
l3kKXt2P+xQEb3KjDueibVn7NbHw6cxcfHPB4YJBxP+cHaJ+Xcgztv7NrBdBU0pu
wkJrDHIUq+HSA1nurMQj9IBYmGd7IICUmEp1FPA6rAfeV+SVTvBhjTX+kYdwspvy
+9Apg3KYf1TNzhlCopwfwU39G/pyPKJeCftLtjM4ZDkv4D4DD4a99YhuhbaOGroA
BqE7jH+kZWgNALa1zqN1Tz3tchS9KKrQm822jDM23aq8iugb6bngQE3mdw+LeXqr
XRrwsAWosSQ7UJhJStDavXVPLiMqAS81BV4Av8WmQGn6jUBuivMWGHyMGJF4XA1h
8vdtB2BiddUBIkMCP2XUStjuhH6kjmZYyMzp8gRQUfBwK3waCE0Q2DLnGuwDw65E
a6BPbgCD7DkoSL+9HkeEdS6tREaK2kkte7pN5DqqkOaoRRIe4QrsxQa7eRNTTZ3E
zKBPuAnoyBfLR/4d1HoZkTgEkk70estY4OtPpNiZVCOvxnM/QuYdVgzoh5Jk0Gfg
6e5aho975apo2Aql4mP0RZq8eGXipMHylDSkuyq0hQ2f2QmdOVfVouKLDXWKfyel
Xa3ZgsmWJq/S8h7AfCiFrBktveaI1W0YjKV8Qf3YfG27mX4Ow9HRkiTL8lQcKMEC
1TeBvUDwgKfr6m++91X92yTLfVdHHV4EjbzjSLk9z9c6Kr2ln2wKc5aJFFaGiATI
qCLpKeQ8qH3930kvmw3YuHzNvoK3v82xZoPNkb3kRP92qsoFw6EUaPVYRIzA9ZUx
SJrIDS/XKxSw9IvjYiPq4OfJRYY5xqrk0VMfBIXZwSwV3nTieLJQO/aejhESxkJV
e9rqj9ltLIEmiWi78lxvCnxTuA8alZjMMl02TX1pJQnnbEhD8+JZiX74FFwMToBO
F6RUE+JyH35L9hzLlsGh5ZLZz+qD7bXv88xTXX0OLN5aUqqKHe33bSbitv6E3eRd
rOyk1sj72zJ72znW+6kyzs4IYk0UW8LklHUBbEEtKv16vzumvrQ2bAEI1R6j1QDu
56uSUtEHQ4iPb0h3uxz+UsWguoRPUvD3RKnxwo+gCVqAvV99kud/tKvvaZy85YIh
aR1PdIRh416xyq3nKub8pP+aB/1VneoSV2PCOcUvV6g3lpOwD1bqHUkCiPbvYdqy
Z6pWE3L3p2R5szjGRqbX00205nRTkJiSpe+IEChpqWqPAhC8FyDGF3V3cCXXFN/j
nFcVufCVlZ4lA2WB62kBqz8D5wlC2GGmSwGZsICNv1lNudRPGL9vCh1OY1nGBOZG
peNZ3hAzyKoj7W+/YJWes9qGtV1GybHiLvpvlPDQ2BvkCA7TZTDarStPCdkG4oOU
pyn1zmofbT00VHfQ0GzhQccaRxS0QxI7iHSEB7kVM24zf8vgeWMI96309SV8rd40
dEag5WsG/SLFsU0T2c2JYNTfVPbwc8curfkuQYLNI3CaxwU6fvPugWc2t6jHvJHQ
apG2w1XxPoLcRDqNRnTPx00XxyBmcvkur8NgO+q4dZz8rb1NsNMLUtG4jVRDOlO2
aXtBs1wubj13TZGPA1gJ33NiuEW5bwwUs8/dHwpM3J5BkPJ9fHTVVaCu1sFMII+Z
rA8MecKuH61Kw3kjIrqHv1QhZGiHgWxW2yq+q18+C3cknfzA4z+KzbrWlir+9FaX
1hxGlfXAj2B9nrLo61dPPx5p03qs0LAKtjPcwfFAWkDyeYHe9FIhkxhMWPYCA3km
RZZJ3YECcKL8kRbGAvP6QBwfxfl9BKM+X/hNWbU5MLuIXDsygzc3Bg2KLtlBdCmv
R8HdCGZ5gCp5lWz6sD6GZ3Fx8WZBd94z7yVaHZMBXJiL+230JhV4j2jO77ZmoJ6n
5/YwNL2rZcC1qSYrvzcBWnS79Qn5mLbAbWxKb+UBiHCxuc8cxYhD79uI7KohBB9O
Dh1Ef0tx15SzRAja36OAJcJwthXCSesvHwYFWIBvDAdCPK/UhBPLcmf5XwdHUpMi
6LrDMRKNZb5fD5dS59ooYsiexdVzNRfzoxh/BW0bvubHJuk4lCrsOOfhfQLswS7N
OVsKIlJwYpdKvoyq9FOJiWX7RsZylDkKURcCjhw77GOcRKX3+VSJaM8PFDgwkqs2
yMUOYxoywUL8gIQNBNeK6VjGcBwG5DZOO/VYXdB75e0ZUGQYztb3KJ9JlcU2w7m6
/7pHgPP4QPagHfSnwIyeo2RakHe/lOJg7WJol9RnNtCHksj+bUJNhUhwR4ePa0Az
eiTodoQ3iaIsmk8zTDj6lLWFon7xS24qOZeQOwmxubUWEHN0E6I/A3VD3RuQoryG
rtJ3FGSbmCokKFsNUNv+YBJjh5EyVEjJd2q3O+SDNmPxsQIO0ng3NXdQgf/ULkgm
GANwd2H1fiEmLbVYs+kaoHZCKpae1k7VPurT7RQzG+o1u75eGvpHdZYuJP9Re6xD
4yK8IaPuACVZvxN65Jl9mmWlCtWRSWXbmyCyRSmD9JepwngQgukbw2N/0J4jk1eN
Vo2xns7Up88vy93Fkk/su1USfytI6IRp6lRjPU5o717SORKIrY/i6aBibYxNWyXL
PCVjvGLhReAB6PHurvXD6IPVdWGzu4+gB2XyCtoi7g0Ncu0GH6gFF04kkGisAVsy
j6wImZYHLrzJOyyBmqeCpnQ2cQbEncov/ozBbEFk958wBZyKo1jbMfI6ATnWhpQv
w0WTUas59EqoCYtBUX1WMJ0hQILDzr4ZmIwp6x/rNcvKMh7ISIcBXPZsoK2ta3A9
eOcW7nKudaPYm1Kt1Ww2hv9ay7nRMtrwdONDyvVsZ074VqEVtS2Si0vmW8WxjoWg
4RHe40zBtrbaPM+KqqBkcJvVkS0w/EMfBZO8WMrYepQPYj+XGTjN5KfM/lSbGsi0
KAze/4tXTFqGwAgN4FOQQlKIkpnuIQvELgaWspEdYetCicn6x1W0kzhTiqmkLR9j
sEt6NmCcz0Pzos+wVG+Kih393Pttq1uklyM2+Q2o753IOVvq5LtWxenIjMmFbnvR
jmI55U21/GjVB4B8tjXfaOlMmwzGoKDeyxLu6N6iq+xqF4Tegb5i/gTA8odAEvQe
i1mMZhAgNIauHDnCn+zOPmMDEztUiuhS8GnmtIRE7bGDbV48xhNtIHsRhPMSqyIr
pMyvUTnyLRYFiHE0ydcVSWM47nBDLxe6t8qHX+8XYVDJhLoVnXRwRZH2OF/U4ia4
B8lsyDmYTC9SmATjhjK22VXnXJV4f1VkxOR8mUjNK5NtpvWlUa3RXGhKxfydsliz
YM98a7ZvmIfVkmSMTTQFEKq7v8ox5qJezj2apaZ+kxdEVDLlsMu+E4kApY1ISVZx
zh52O3DGC7i+gZZwUmzrEbXB0WHmdaVSSXCCWDA/T2X0m8ybde6+Ze8KYZiawfPB
u0GJrG+7xG+uC1UJaWLeHS6eeBcFpzlOyPyKx7EE6dge1tEODmub/+DscKXybLNb
M+m5wLinxJIIIsrHl0PV4nmzCYSwnkveIwQf/QUsD+RXBZ0DcwC9bQx4dTi4ZPfK
FGyXYpq/eoGdhGx9VSuhgEokyOQLk3G/zTvSxBRqejsTGupXvTVTThbrR60KNlWK
CrQ1b8cao6Nfp2r+fD+FHHYbX+TEEkUUabEAunH03SnL2yubke1f9NTyN7vRdrBJ
+LWbYIEa1xUU4NNgSy5htP/CDeDnpW1vXPu47ZMiiRNvVGV5Dq9b3FstpGc9sA81
rHCa9aShOhT/tRzlXOzP4IaQoqyXLfhReibQqaSAcOAaw6TtdAoPjdGRrc7AtUCN
Yn6JfenHNhhxRYnmcf8RFAj68MwFuaGH5TlRMid9Lo1L56w0Af+Fvj+57GzpZK+b
lCrXQRnuJy6Zutn2BxcrPsmTdPfu5jU1K/dyqVJNes/vlBVF+e8qbNMQsQvVut1s
v66knk9xpErUvOmKJQTDAf82MBwZFCmPs2Mjxa8XVlgskx/zinL3YvRsmqKDE1A/
I/6B/FWxJiAGkzoXh6d7P0wzIfb3rWvO9OikqBj8khQ8gOpOvPLAhePdl5lQOn8i
MlOifmf8QnYswmZR76C03S92eI0TUVDTA65LaXyb2XS+wzhxGdacBvktnuaj5tXh
5gwZWJ52iZ8JkR2l1YWIulZs8h0c0dti4N7b6R968JU3XQTMVb7Us0ZRdkADJ8pE
1Mm4fy0yoHpt2kJi+BQ+J2P29+yBpXoInNfSf8a0uOhq/ouSpDpN9gE1WkCBofxK
XrJ4np8DGbe9cHJ5RcMdu6P4WJ4GPgJSrZe4b3HBdcMJtBIzprn4MJNyYG3M5pwU
61wILfh7N3lUD97NJTLYQaDEdo/kLLADVrnd1KI1WEBM3R9Bl4FyEh4VoOoB5u5v
Jf3qbzCzCgIRRDvAcw/uAdmuqW1O2ggSIuxfOQeCrd53HIVP7Ou89rIqFxfOXkLD
gvH6p6DE87EcoFs2torbbggSaGwmn7VEmNoWaZb6NvS1+M1hqNFVCtexKPU7IZg6
atZ3f2lOPC1MrLm9+SKMssZM2ajqHK0B59MuD/1zfivVOBRzW+wSqc8BgAkQnN4R
9NJ7ncnnKNQ5vtiqNHyBtUpCEMFTuE2cnn+4pid/edQ4R7a0wRk2MbjpIYVAGUZJ
ibPt+K3U+gK3SBMeBoazbW2byuh8rzvHPxfySAlGJ5jo0+MYKiObK7K43znB9Lzr
b7EOTGreOZhUBui9VPvFQb90TT/GymII2lBYfaxGARUXsEMo72Av/98Df5xLVqHT
Dljf1+VirKG3+YVzs6z9FcVufNbWlHd8hJ3WXGGQLdW2NXbkYKEgVHz/zrMxwmvE
TJ3uIB7YPj1d0jEQP4vek7h5zw9m0a4N5gd+EOmXNdl28x3eycmjvPr3WGj9tO6+
ZeTJpehOwxSgg0L4VK0JBxE6rPhcFfpbJuKyOYgleNLgS68Pk5uADSC0RgDW9TDL
r4PNzPcTYfWtaMDcpXjZ5IUYVVG1OVD9XMC0u+Hze/uhDoZl14joOIQMZIGU1s5b
m2j5B7NP9Xu2COWyITiyhI0P5/kTsJ1DrSkl3cDdVD3Yv78EQo6E61Vtnf5Sr1Jn
JT6QT2sueUkHjMBPWCALN7Ga4GKyyOd13MxAL+Dwi9ZYn8G7oGqFAQvEMuiBepOP
YpHr5G6dnRUv6p5KGGmkTdsOSQr4BriNJf15hBFSmotVw7qr4GRYCYKoCkOzS/6d
wIIn74a+u5JJhgntCnhr9cRT9UNl/p0lTRxMCtNOfZsE7bk6BpfrrUZqmGu/qtQs
8/Cc6QqjRkeWpTwJCyRMGY0t1BYV1kyUifxopKZH0hiBfXs87HOxgxFxNlL8wzAL
jIBzkYiqscGcV2otlc+D2ysdovR4okla8SACyuQYFtbvFFDOIKizmA3OlYt+0uek
KpKncejnMv5fUG47lQkEp6uYKKRyklOeK4fKID3S5gu0NUbAsTPMPo87gkv/jXdm
N2EiptdopBxF0/xDN+VYoqeKtCWW14yjuVUHEPm+gwN0fyLUUsoZh9qh3INZudsj
+p6rBjl3OWUtQaw7gvDJbz3j+yAL4RbxmcOZ5uAOq4+haf6oc+/S7o00Wkjt6vkY
/sFE++LrECjJdWAdKuI/pO/ltS+yR8gg7qE7aOwFSNjrqvlHEuKizcPKMRjIBbIf
IwWbI9ChzXp/dq0cAVFRw3TV3UQ5CkLkVgRJ9jVfqCgmG5NmEK9kL+s4lxs1NVNM
0dzILAfrdrsShBUHY00GcCqLCqwXgPF7LSHu4K+gc8TTan+jpqV6bv2bODPRKQs7
cCRn+36bITa/sGrHO8QaWPHR4xpDp5qfaCZMDNvYG9CGVV13i+MGFnzMUOQbIjvz
WQ9N20nH1GKpMC0fAkjEDaQgBeWGOctwsOkUjnrvVrZOE/T8Pio/3PwBgqyPLBsP
jzQLvUcflsemrmExXlPJCFZ6Pr6gWFwNYYSNqG18lcGIMCnD+ZTbKA4aUaHt5vJb
NNa3e+eDkQuSUxtEXk72+tbgP0LmsOD4oyjOmV+r+4w7DvEQdKERnyd49fbjPeYB
ibjiRBW1oSd590Z2X+1YRPCE1x4vGpca/LJ1YdZxPhq+LEBFD+VUW7dO4Irg+lBz
oUHIn9uRCG4q10WU4h+315Ui7BN7CI1ROrhaZqJGB8O0BDVXdLVlAapbb0Kn9OXR
IcpzF/+U8rLXuVBR5vR0snbDfjDoH34mCh38anxD+dGtth2xHe1PFlt8x6lFH2b6
AfySvEdNmOIfjzy+uP9LT+gqNWsEvhPXnER6QJ7JXJYKJTwto5fetDuS/ZNTnQQx
WG36BP7h50/T14uxIH6t91KcuTZXgTOPxu3pl4Q8VlggQGr/SiZtZvW/IxqY7TIc
MVQhgU89Xk8+yXRnoWr3ieLeG44fIpF8kpjRDffU3fqE9VysC0J4rM0gWy0b3IWB
DcEhNMLqFLMepvGG1XsiVpwjGIemPgQgKMkgLSL+LbDkyzqJI5w/cRFKdOQlI75N
afUx1MgK2S72HVK0MAcYQxiHcSQulJIsxH3kHUMe2vp8lc1Thf+qRBN1RPphvnVN
RJGeSrd9naAAp2KwjmizbGcW6cLukNRwOfy7vbWR+30lv9JKD2tz9W03UKP7Fge8
4zXaojvTYxWiy/elRMEUly5344k+n3RCuc7h6SXON9NQpY+fjUf5TQg34BPuJTn3
x4exucMhG3ucUe/jTsmI5SXnMnc5DXYHNBcafSvgVC/LaYNh/F1Z+2V48egWKfkC
OVLfQtYb2Sv9dzrCJGlRJyw+34fBtzQXkOFcv1/5anexZ2xyvi09WWn4udZ4crzH
O4yS9aMN/7oYRtKHYqbXQPIVzIhpV5DyQJB31d6DE5Wlolctckuoj4FuElGlj2lg
qgY0bylqGqIU7fANFIBooW7Z0ipg239aDEaoHCqCSxx0m+D0SzgiZP2kVST+Jzq+
83sJZ0r2hTkISJPcJlgsz4DadS/UukycbYIwy8aOIe9+f6aYy7JA6Yip4nxeG+hT
+Gaz5fuBzfA45SQ5/FqhSj4yYB4XYXpQSNGKYQvuWA92nO8gf3UnK3FXz2JHVl5g
ojfPWz5UEHmL4UJ1OTY20KN7K4ZShir8kiP8Mh+RnZSbLgMDAHYCnCXmjqSamVY0
GsvB9VdI/n9MHESGMnJ28pzXV3P2xqqNfeqSs/4mlNt6joUfVaB444l70lBC/+Up
GFyrRIBmQHzhhLFaUjrDdlYTe5os23PU2zc9/BuiFdXASB0z2WtMvGpfySRTyqhk
73S+GuLL1PNYM0qriAiZm3qXMjlxiXt28EpTu3QgHhaCLH0VcHamYTlWqvfaeY30
fPxSLwqgvINlXNtpeHIoiurEtStgxO/a2V057gP5us5YBZlb/8ufquY65POyBhTR
dELdBuGrTa7ACppdRB+IHWlsnJ917ORMXVXeAc0dNpVl815eytk6zDqpDusQt78a
r8vCzvxIew/RK/JD5hNQ9hAvw7BaWMdoIt3/XWKmZecTT6pRGDZT+YSIOOX1C5L1
DuS8nOCPkkPIhA9fG9IuGJvJ2PCVFqfCyo/s+deKIerCGScEQ8GCGM6DSL6aepmb
vW/tHZNPlm5a0o4SfL1Jak3l03HlAVJ7OXnig4X72//d4OQj6sLWHbcJgSy4zaGt
4FVGZVU+YJLfXgqabzFeg3DOQD2GQd7qey7Jn3YX18sfdRdIe+uAH2dEJsXXSaUW
fDiBj5CYX7rFfqBzPtwfR+R6BLfyhkrPt7fxPw+k/N8uYxBydQlBqydAPFs2nvTp
4rGz6zGLiSgjzPQ156J8dXV+NZD4J7/RLwtppRWPUS3rZEvAL4Enb7QZiqtgSwYA
aATj1RQbpjtHDNlMIBy0oF1UR6d/xNDkNha4D3mzI/yWMgvUxSszBAIebYBXyxji
+iIVC7Vcm2UhDvi+3ku9P6IRXOdAEZkfP7XoN0DGNybd/qcpAlwEKifrHQPQUaD6
mxwNaxksBtINNsEQpVQ0H42kpan/IyE75avt+mKddhg5S9fZ/Pq8EZR22DpjBAPq
05NVqsYI4AdK6fPzda3RsS4Vamndu65WTPWvtUkLqRY35lSmMW/ybb/gtmTxoKAp
J8jYn3u8kUO4avoAWdkctj8Ta2pVPf56BScCzDILgiCeZewTgbGG+AiBTA/04+PH
1TwgYnnL+MyomPvyZrt/FMr5HmPPEQfHd5bc3vYtoZ8rgniB1ZXbkWFNCwRKmSmJ
rm9etQqSKaLpBdl1YcyZqiLbDAg4mHzmQV8XHuiBqqhcQhlJTQs3b+ujF7COgJPr
MJ0lNWkI5n72efstA6mbDIORaNozqHgyYUQuHaGwrfPVDM7RU/IWw32QENlatTd0
r/cp8FNyS4gr3hj7W7bWgExmjlUWrWVqX5PFFqF+/vUUYYzv3/WmReQ3sRPu5wcn
WU2ew+6TcT2L4KyhmHQKGQoyeKRU3WRFXNUanA97ii8JwEXfqqoVzOqgoNp/+98c
d+EtrcEk/UceKM6G8po52Qjza8tetfjAw7+UsoxPxw/X8ROnpSPLhecLCWCHwrKB
LpWO98n/VVvAjc/Vx5Y7CS/bttwCaFheywMkeS47vevu1pcKtKsP0IwnYGLfqezU
m+c9REkevIOe5Nbw50o+x1aj7TGxoIZtEY5SA71gLdeDEXstKSdf87RME4/TKRMW
sP4fguYX32hDta2d7bRCHYEl8IZ1EiShUKYHFcIoyvidpLy3AAzSit4aBWDYRAr5
Os2D4GoIdwVkApxstgVAXHxFF7ma0XW0qsCKSlVjciFAtDTwii9EYFfmNKl6Wz9h
RnhBCk/nKl3Gb9378DB6VKhyswczHaatOJ8eo59oCciC5L3RgItyNEhR5flJWV7k
afFm4VdPX10Ru8wdpfZiKx2Va4lkP+GrDLGhbvcLEzcuZZ0FcoN93w+qcm1Pt805
9O8TZFvm2P6EQW9IJGPfLOceAfbieNXJpYxzogBFGHcJpc6TKNF4s4VC1/DitA3r
lLsi0Xp0eZnrs1WvvlqG+p/hK6MYvLH99bV/DTDkndS5f0f6owa8RUUtOsNgogw8
r4X4N3/Unnv/DIxu6owH7wq4KrYVH+w2ZiSY2sslT4AnVq/Pu4SDTX+cwWqqkBps
dqLDEkkRqfmdsoYT4GKDAt1PAFFb/DUkAlXTedQq/8LxZqzGl86K9NpqinBAhUFG
ipcSlMEHGqb7oYD9G1lt6YEEl46KnYulU/YLuPumyve7uhcnN8xkmjFsROthepqE
1cjvlyK8LmWKjHubgwYEgF8Fk9ntWZ8GQwrS9Juj4aA9V6K3QvRBL5qB8tajPN4/
OzmfVEpsNSAT6QAs8lDRx29nMD8KaTME+kLaumKjKnCZ09fNmt1wzahrN7LYQ0Ys
EIZREQlaYhoZyimR3tH5axqQzBf/Jk1L/4fzsAkh9tK6yhm0mGmPy43ZebviNicE
2/J7eAVefWLs6nOB5VLHJWJ64a1KpspZo9Wz2E35HkFnTt0K1BvvXLjfsBGFzUrw
twin72lxrBW82MciCWk6XE1Mjxk+b6Xg3j5E0MmFF56AoZRBc1Dkt5QxqJtClZMK
Ey8t5J6QmJjn0huQGuoio7uOsiS/eStRVQY7LeFQfMMWfYPokTZdNcY/LlLY7/sc
s1QJrFpyfF5Jg24QThYgs8ZCF81zKDCod0pSo4CiMhdq0xOwWG4tC4WuCCYph0us
gMg8AAe028lP2bQ6aGT52Bg1j5sKewo9LHTJtC30e+tKgzyJVrCUMXNLqRtJFYS3
RT0MwrNsFSJX7DZfagVWfcN9z/9GH3eq4UU2ZAqFhkP5jLr5kZeTZQs22dkjHYqN
y1smz7kuGtdkW1zaVpEXI8GTkHCppOkYF0M0zjusv9VjKH5maIk+Mf7kw0URjG1Q
sPqFWyYvLf63BlvY5qBh952EQywEmYqPyjUs+/xLW1bp9ca2yXbdj2nU0lM20QXh
DXOuJH5XXbbIIHn9H32VoZSfGdnRXM+rnHLSuF6z3w6fjSwopFx53nWcLWnAcvq1
q3cTBK8nx01sglPf68EVwXgWRBze7qxyemj5QPd0xb5PLxOvCM7RWtVB1U/JlHR0
RbLve54dctQNg8pq0Yd2ZbDHDwTrap93y/XTRT+rTr9ls2Ra8I+6pQmqXOumx1VT
JqJ3VgLfOHGVAE4UbwHn0ye40n+vqUbz9AcHUjJk8ePaoWrgCjc4NLohfdpUd1eA
JN862t0RSHzqJiJudT0jpGLCmjsjwlyRjnnwaFFfiN6p+6/6EUFmrTSmX/APfWyU
sxukK5jF8Dcmcp1SM1N8ohRflAcn3yiUJcZq1QqYf9+7R8SMkdjWUvYJ4DhlnlIa
o4T5CQWWoWoCNyLZqjttXogbYq7Wi5icTrwZbaqdsoTKljc+cBko7rPXGp20lZPL
wA43rMhYfVAcqAPpdT+XsiscHLVq29sy7Klok6oD4UI0ZXhyS024sQQHhlEy2n5y
Oxuax0fop4U5Ght56quq5sQgkYlqyS+9CfHHQSNeb/z7NcxTl7/9Eua72wEfAyxk
pP15TyNYoCFT4Wxx9uzwPbl3fFlWu9Wd4KhlrhFZgdQ6om9H4N/INpGyHfmnKOCw
HlryjFk3vkm9DM5IEugv/ZfVp7Ge08+vPv9BxSBdhoBWV4z761/h2uxXlYgVr1DQ
So9mqXKUV4C1PRacq9kgkZezdQCBHHYrqopI1s4ArIm3ZtBWPrAXca78+QihMkSl
lqmWvKO24QEIrN/57GSgBYYm395h5LeZ+5m5oL6kZgVNAI0f0fNte/BEQEXHxwaa
l242AHyxYrP9NYGRjdiOexaM8srqtPmMOBLZ1XvtEqJCJh5+de+NouOKcW/YhmU8
yuvl+DMaXlEZKPVi5AYkZ/UhbcO9+mEFiqG2lJPIqN36uMVT/HPR+KgWJRt6ab6O
XjfnMo9/KMLqErTGUkpu5Z1ohZ4gXdw8vB2/0uED1Q20haZban+1v9VAznG3iM8A
etbj7ARpETbmVfrdvHgqBvGs2Vw0PrqnJN3YbOmxeNR0RmgNQ+pLRp0QaRsE2YDv
TwgdCnMIEJVuamVtL36ztbNltLBQZcBzkt9crRFOCdvUEXEKEkrMT/TK+yHWRood
adDrS/D2zt0HzstH29GDOwR/U+VaWRFT8KHN2jKDR5vl9fNs2ItlIACd64MhiYFs
3kJWDlJp445iPE2+/W7IzAw7aOd2uIeCIjjcxZM1ciVN0um3roGDZhRIpi7ktiJ3
511Cwm9yvkmam7H5/69EbFTxtw2IF0XyXUhnITOueDpdhSxl8ySK6cSL3gGcgFq4
f1crjlXWkd5L9hpDe9UK0nLVQSukdkG6qVDpIqsWLpZpH5ZACC7+KtfObWyOTPLA
VvGUxbItKFGfVN7neybuO19coy28RtQF1jcL0JajAKdXUadqMT0HsfDuLaFjZ1rp
fwS0ffFIfrQBa/v1iTaPGtYRG1wrhWHC2CLmtSqnWWyguNvnzlFvLYJnCjS8CGI5
9H24c5ehpgFIS7yvdfKZpv3u2AhhNhhPj9RibA6wa2N5o1QnqbfgZUhuaScxiTPp
amCH6HBVZbfYNWCSMxNmvcVzaHJm52mO1F2bzgtBjc86+Pk1IFAQNqcjlm+4l/aK
sB8VMGBpVYI0OZCyJSYwDzxuLpKhzUQNAFfc2v7nY3PCKGeMBRkqdOaJm/3HFnHA
3M5a+K6hE+IZ68Wv+NLoxjDaT2Rl5tW/3zRXvA66SfJMENiwlaNyFxh1mRpm7Nkm
X0npB0zu0YC/yA2zmOVEzYTwph1x0qNytBOyRjjyg94jPlD/VNVF1DLPb/VABL2f
4GFHRyDep34wvrubrotlBFQ5Ahh+6diyJLIM3NIqZu27+mBM1ZI+aZt/QHSu2ea0
lNAxSsAro6ej8x3L2qFh4P/ZcCjzALCWLEqaMNml+mmUgRDquKpyf8/8dGzR+FWG
L/nSEnqb/OpxtrpwQXrweA7N96zM3egJdtLy7xIWXooc1dDMNp8XN0XSTVQgqwiG
ekrS7yI2OJ+VnvwUZSQZYc3OZqkrA6Pp9vkMqM8Oem8U6pIOyMGjsfVWs/O3KO34
lH5LMALmGwVcwQAiG5OwgkOiE/3xCUGWAyY/iunUsirox3iHew8LxEj0AqowjD44
BE4JKhH7oXmjumMX4L77FYLNgw7a+v6EuDvmMUNeaI4f5nRAKC6nPJr0Hgt4pcNA
6sY9+gCXkJsdJ1KOa1f7Vlzvx07lnBCxLtTctSt2+5xH5T2niuxJmSpImzDJ1JsY
HQKgdasGMYRzbnpEIAzovRdWSmamZ0nxYlV59KTKC2UaHu77UqPG7n4Z6duCU0SV
rLq/AqNssuT/48LzM+FrgrXFHXFtPHcKqRAfljfkcqK7JX61ieYGfD7hLFgHrTM6
eNGf2Du4pMe2D0Ja28QwByCAFOKm5hHi1jyxMn1R+iVj6DXwnvKPGmJ35nvvkaUj
1kWfhkqFwG729aYeVwv6OJyD67O+4462I+JSboi3tF/COzxP0phRdxSPoGzk3uyU
92yrVB9bswP1Vft+HSSdnaHabJhWoY7f2YoR9K777KzDFHfRCOlNlJQbcs7moDfA
QhA7CxjwHfU8Ed3NW+Yb5P29LzW4aXEyopAtKiehQCBD6K1JzgUNDHBk1KRG4iCH
mYpsfv/bicN5A40xkoi1/IO4o/N+QH0Fk7ZU7eU8FAd17h0MNH2AXTBCFxCf2y89
dtMhIlzRuGxRbT2nBjVtjDmt7svlbl3xS6nhOO/aG+oO1kkNFIPTWET/1PVknbVW
KWdO4Efu5TnwXla5cGeECwueNrheLKXqFqIvG2lp8vZh18pOj6WfA2HAMCFn/E7u
G+GlZr0/Aesn6UMXEOrl1bTyFnJXatCVUDGF7qcLwwQVWbuGRXJ0G2tH5ofqicMc
HTuEiCuRahxzGZvyniRekeyTe9ps3gL+gd1FnqvejmoG8eSPmuNO6fruOjAu5Pa8
9TBGA/LGNxJYLI8WlEqdow7mbk66/P5+Q7y1kt801GTeKTvumplCmhrYoVeSlY1g
/5PXTM86I77Qx0Nl0/WYEL5wYTsH5/n7TrIr7HhNDDDr+3mP8SUr9foEGlg47kdo
Lz49hzn01qtRgz2VcewXSDhkO51g36yuXri7B+NNGYIWSPZ5ZG1dL3v173s/swvi
VphHdumNaZeT6/IR2uXrP1bngFaubpFrrVvKMea/wntLAWoGodnlDCHpzSf7SkiG
wTAwVeyr9/9rBBRuzIpOr04H0b5+ZUMd84Z0myzsP9r7vFLCUfsfhEBCLqHq1e/W
9E3GJ8eQ1klYqLZjngK1Cp+LAZSnrIOpoAuiMmBmpr0KuoXL3uRmWeDXQCqU7h3P
kMZq+rV4IQAbhQKu4MurtFWFmJQw6yexTbfBov+yq+nHHQSypOCB8PWBYjsZhUhw
cBuW4AwijmAtm4QH8erRtnm50gcCE/8TFK5+wWlq6EPvbL066Dle/jtyhpysilN8
u8u84QJcCQTHrzU8oNv1AiZLj2pgLHWQfbI3jOUxaDxbmrx2z9qcPHsqXoKWToOg
4MWLi+i76oMJ6hxwZahLfTCZDapXmaGm820k4a8dsuOIUGdsRUodSLUUCSbaav8z
U38uVNLR25vvPoiCKdeB7K4Ud91A9RvTZgj97K/ZTEOynvU6BRZxK5sfiJqpEFp+
26gBUnXVtgCONF7WXVDRQPNE+xtRSZkkB6FX7Kk08pAAHXrcJU77+2lKSoQvSqYY
4qxCkb1Lg2e9HnREuIYM5SsSUt9Wh2rxsJLnHIrzHN8SQ4HRkBTV43U4BflXW6Sy
l/e6npAbY7vn4LmcAfu+AEnn0yjU3BmNFy2ssSlLFDPLcmksCnoUT2KITajt6AS1
dKXbJfwrUqVd9ldw50j13vUzflB0iwGZhbKIpWCsclsLqEaifv8nuve9tOmZgQyi
4myx+Xv/2d1LYSeEdYK9Ths81pXgBTgQUml1xYsAXyTUfJrI196c0UUrHka85RUI
8nmHYpDwpPhR5DI/0TdpryPmbPPUeECruMPKDLsssztXqs9jhV1GDo3V7mG6owXN
Gr6aBYO80alXngwFEEBRh+NsVNb6rkrulJaNV1PreR3PBpKXrAPBgaG2mK7Y+YcQ
ZgLWcyxwnY/7yjQj4wvXRPnSObIPyidZgMxAR0AIT42Tg10lqTavdFfUqTNny18z
yGYW3zU2/nWx8C3bjV+ic6jT1GtlNDWWmzbeZkvvmFHaX4/psUAmVJI1Ex/JwfHB
M8S2xQjVs9F/8T9NI2ABwjrtQt4EUrOgQ1kmfTARi6Y+lvmOrx/j1U+tV8To+C2n
UO5FR8ZRWwziA+qeeCFIJh+8i13dU3J6rvWqQNex6crSf3fteq9WEWgkSLi5WFm0
EKhXfW85riIeeoRyPwRMYuO94Qql4b1ytDrkiYAFidO9dwoubP9/v5v46q4O/F6k
7XQUz06fYbNNyrqk8OlJD2fcDiPlyxsIQR1ouuzVR1KJsB+pVlruhYAgiBgxVpnM
uWj4H9amPEUdHrfIdKXWdCVXi4gqIvH1jXK0hBllKBiC2U3ekTQAtkWuSlmXAeZB
k2lwfxZXfECiiLRWVm2QtsMItYejKVFuIt85V9xE+Kmq9NtRbM63F1RXeXsoM0uh
N/zccP1/faLBHlxWFil1nG9F7akEQQGUgRoqbQJAwf8uFWqOBIh+Lqiul4HVzhpx
S6gZovEYrqGU/GpvB1ObVrsdXsz0Q0ru+bHGy5Eeb1vRGC4ypiS8TCWtqQp+klY5
8x6QwU0/zE875e3xL0gtT3fI7m5ad7c0wEKVIlgRVeQFrTz1mCgEt3uXeopUDT86
vXd+X5BYPnwlpyVX/g5QUnzk8efqUJ7yaGjNjcOhgcA4/6bg5BiOeG3Ns+QHPchA
SUVCfi4SFQrSO9ExGWxSFl4HpUFFniM3A/VWNJlKZetnruOrbN1eT4Cg47FLzvgl
wOAf0Wy/5Y0JP148JNZBi9R5Ph0lRGCRLowgkE/6YL/L2trdutUNuH97/nj5XyFa
EWrsV8FyOWo6CMCEoNApi1WsKVeojxgWfpFYJik80Pg9UiD9ezxrN+Ew5aOA9bxZ
msFfRL0odccXyuaAsZ7D5jthnS6OQuiwmVKr5WuxzztRT9PegPzEt5xyMg/Z931f
nRzXIEGfMPRt37g8B5aea3aEETTrwAJ8DBIqpfUV3U9bICqu3mhPgW4TxRt8VcTs
LX9CccW7Dz9yTPsMD3D/RON97f6RAxDS+h2oSJKJeEcH1DB1BaVHZpkxzpVMvPHk
UZBzFvVeD32jhcVWlzQW52urCAs4Lh2OmOa/m2xuFqYePhkeum629CGhNxyoLlm2
WR01IXH7zpOnaHV8i6p/tjyBG1PcmJLxYJtpaOgIh8oe57bYcXni6gB1B+4Lt2aY
/19HVDQ9q9TL/fcM1TFoJBIKE5Gi8u3zo/1N8Dzu1wxwnRSSvUejlfo0BOjZNuwF
G2rft8Oy2cKv2YYPB9JyiDxoxKyQUJt05NUdoXmfsO5ZPhZG8Gh1lWzND+JljuoV
rW9g2purAQ1yRd8JcPeDEwZudgVXKawLBw1wdj4dQ9FtcTTYOQzbI7XCwv9jBGQk
CNsKcbcbmjDU5FrdPjGX99Vo+xYJ1YrciljkNmNSABIBFxGN+BW14rD9NfNsztCz
VyTCs94XQRPSrX9HzO8KEf2SmpamjdoLebJrGVm1AUlcdOlhec9U/x/LK9/2X7xh
egXfLZlqfcFfPQRwZwoq//6fzvoK9wy463exXfEHLK19La5W8EyrgBQzwyvPtX81
Ombkfa314p4mP5qVOAJbTsxQSEbrA4fBOBCuq6lyadHp66gooRXT7K+V7/n7YuTV
LhRfbmqXZPIwszmWiSePzMijrHb7k7oLPM5CYAupctdLoPw7dF3RpfMKWmNEb9qB
RKzUPxIbZC7gGa8bLK697d7koV8suAOsxzNHFOqtm/9Hm9qJswNIfRAwiJDntI2A
YoZ4oYf/yoqoPxpm/ALDezb/G5gbc5ROwm8mWz8wKHfGU6zFd4EzpiTd3roB1noo
FY0mkIkmVXRvfKMfttq3y2BA3/rO7eroJ0joRhYpGEesipI0fpM6l625GvZ6/dy8
kKpUrdG1+7WsMM0xyqQ1i6UFhoLezYayrqG2ASC8NhEVt0XBjIQldw+daC7Ixx5D
R6cLir1bNcUqFyFvzPwCl98GbC/TdhcQcS2ZqEOqQx7Giyad7oEXSejdqZq/8WdO
PTcimmWtmMcOZINpquKMSfIjeO7S1sOQEk2MZTNdC2RdIoVBUNOe0Zkk96vlv9xC
AYLaFEY/vZkB9lp1MnItfivm78XJwNBgGk0sFq7+BRw1hsEnBV6hFRENxC6cNUgV
XFCK04Tn+23c9FwAHEOUqLV6JUb4//c781QRZ888up5QeCRD+JFzz8Vmt/PHhaCd
OwMmv6OjmZBke6OFYUf+i9VnqN/A2cfm8wesMMjbrcahQvO1WHLjt4qf3xuTXnWA
lj+EYCZOtrdNrKdTlMnA1CpRFIAufhrNuiZBq/T3X2IJ6m7MhFvMkrE2kRadFi1G
ZcdV2pNdPh4Oeq9G4pshVRA0JIBOYFNdYPeK97e/1TzjuLxbTKzydtD31M21Qkxo
JE+10JK4ZPSwUg9yPhupIYVFdcGMn0KHPFaPcJ6mDOIU5i0QgBQezqgOMLwtFy9k
9HQYkEr3fJ/8f2IdlQnm4VSzvue/WhFxB9m9O3KaKg6HUlnv8HFa6ihFDb5u/oro
B4Ol0V/cu6BlULAxKnZpzEymawcLLUrOHR1YXw9FPx5RdUqlxO6f+cefF190Ns37
beOEYKlJ2Lfjre5UKAMGhlXUS+8qanySkWvHGJHGJmUcUO2WtpOybOyT+O60kj5P
RqaeTWhhWUOIbZmt6L+fiXDhQm9u5LxotO4dZAf+0KP1ohY/Gmi9PEtgr03qL7jH
I51tpVOLErYv5+X74jscVmegkHftdox8vwC6w8j68owqedl3k+h5F9Twh6RTgcGr
Cl5Nz7+mSuhZUqfAisLKb8/PRcywpplAfAOxZdKylmrj6cLDDU6LPR94jg7W7wA6
QKLHUZogS7Q5xyv3SQ1UF4oDzCYRYGD+9THTNd1/xUW+q/4luep04tTij8WPC21o
awHJdY3zswBQMOoWh1HeSevD9b4yV9zYr8tjGryaXvhmUT90kbS1Aci1oexlYbZy
YbC1VYVnF6j7WbLpl6HMs3/ELLACkMgsem4oTf+1IGA9l8lc6mLCZySdsQsMy8M3
Elpy5TnKJHepNLblxDAqPph2Ny742Szeu94L+umfHD4bgfJaKXbwNgA5pW3Ltjr3
SfqcgenJNqsH8wvglZmdG1nh61Mi2OT3ksu8wogyGOpqYYhNSOUT1ZprlE2edHk+
p1f3gAHu8HFK7pkfCDt8qneGp9M5otfa9EI1XpsdsXEXU8eYhuiWPh2iJVsKBMbM
fRN7rc/n2VA97y3y1g8ZZS1Z8J30yP5tfDbX23WfzehAzoAV/4NuHb88wRUURdI2
8uZHvQjVf439X2pvs8oMScjQ1KCNYGrup6RRoAgal4UCI2xYRqEQSyemLTpQ1tOH
OR/L9d52OW6o+9NAfeis9Sg5nUd0XAMilHYOUNSq4Ee3rPgdlPFSAiQbwVH7LStO
e5ajO9KQ7ElRTQaaGOGn8dhTaKKIE8/jUkXRDXhu9llEzHJIK+2hAm+Zkn+qWBRh
K0muFPEe01TbfqwcBqSkeSDjY1ZqDsUodZ5lvyh0+gKKPQNzgJ35FRTK9lSc+wrV
l4oUSpP/sBz5d+5cqTlBnzNKUl8iOCOAjI9JqXGzr1szjgAKdWwQW6lTWoOSZAyr
Aj9SAy9aXnfXJNaYIYYkSTO8IpM774jqKG1nD4S5pg2Kp5zIkkfg1+MnQ+YE4NZK
tNgbuoW7lC69/jJGATN/yWJdGUHOumFan6/iiOEqoPkqnotsvIFGd+pTp1MUlcMM
pkzm3xtGHXUlSKnKK+DWQzBdHSEszAqi+7MQ2HakehgDRSaI++7/hnSeBqUOIlWw
xhyqIeEB+JAV/9ofwfrMA5/7L1vp/q13Y28FAL3wFCUSLsObeFhrCqaO1KRO5D8E
dVAfZVXjxLSyKg2qwlnQh9w3nO92PYrK/efE0Wzv9me0FlozTVpl8rZLB+PN9h4o
lw9bvJn9azp9FybLiq5OigNkVQDBVlzCXlymCmK33MSDTM/9Pooe7t5QaZ3+HB0o
DOlxpa9ISBUKy6dztx1SKhWKi/DfzW7rnQCibNcQ8JUt8FYLKVeXEK7EWxot4fTn
8wJsSh8a3LQIRTF2Y4J3vitnQgfApWbqoB0+9csiiCvK57PREfbKxzScRmWL8dNE
VRRESRi/ZR1n6nkc/h78B/fe8PqtBsAbdXK/ZzlDLTBW7ggytVNvVumdmyK2MMyC
0okw7KMd59coJgVWdPIwaodIOPk0ME7KQhZeJDXiT/v3xNq8qB2lQSvwM9Qx+lYl
AzS/JfuLOq6pSMtkNZLhZ4PjXe9n7Rk33kUC+btKXJksSKbhacwHZEo43WA8qaWE
GSf2ZqtTZ75KJSxqTLwROafyuG2yhcfI3pKBhEKUJyFkYtO98hVtU0OBYeXWgxRT
htpTdRsiY6JhvAW6GFvBkdYmWYQ4M1fLEgwF/je4EjG0E3piAJrKZ22KwJsvDPhF
56H+F37/LaSS41GwhyldTizQggD6YOJsCMrQGKupC36ZZkWkfmNcmWIDq6yZbc9O
gNNUtTbxhQeMHrKixqMUU497ZENWJqyhGj6WEm9qph2xuoiuwT9RN34oS6CuZSK1
ju2bEPtTo3ANT2iqIFps8H9Tct7OWczp7HqHX1qGIx3hCUl1wGMvzyAEP2VskCKn
MUr0rtuiItXq8o79fr/jD1XCmWSjMC9o61fmjwUMpa0MY7AymT+LXa1ktw372oL1
hc5zutry0RTVaAj7rzhG4bs1xiNhpcazteXL9RH1eAZpTIKX+xpvJxjBxWeR35I4
uVHiKqRaaBYcGxXPykYoOyx8z4AKddYzjjgj67rAB2Vhaj8oqjwqjYMw2/RsLeFx
oXUEOXRBF/keWFInk3eH0i8gfhauOdls3yi5HKRiF2ohUJBSrfbdnNL2h0QgvbjE
VlYDAc0ADzpTSiHFhiFT02QNFJx/dPgu/qqnpSMasFpxfz3H6xWfd+dHtz7+4uTS
EBPb7Li9Eqhf5V+8LmknnkHYBCAPk3ktblF37srPgvN9CxzJIhtlcpXH3CiJuZi/
7lFOn1tftK+n8WwyibT7m1flSsJPFgE7JjhuzG4WIZdw4bLEaheVjvdGjoZfgC2U
U+EzX+D0e8Kv5fQT52UO8lxlB21JEFAUbP2XMTfkZaccnmUTQQkvJ+9ZxXp/t8yc
bCc06bHyQRc887GDGZtw0xwbVn2nxAKEBjeu6qL3600IEOUZbEUmYae4s262Gz2L
6k4ZxlpwDUdlM+tB3zqw9abyGSHOUbkVEkoJ+XsA6FTlvrU+BG8oqNg2f7RonTSJ
itT2dhxIxcPhcW7bcNQXGqvfHdGv9lGmIzBo9CRY1wzLKDYNTRSmUw4Dq9aOsVk2
fGteKi6NJWNQZ6scL0RLI2MdTKxpIaQoe8nL6Q7nZFuhP6H8bMTRN0LgfFRlJqzw
gOeXuvDVE+1cB4m1GwEhvQS/o+tPL90xW/fFmdkiM/OpMXFLt8r58JQrp8wBPqnV
ZlkEASrrCWnnEKrc2fHcAFFg3dDG2gxRuVPs5BohOj7ewF/G59XormjawOg1ZmQe
xgdOCM6B3up+3PsmiJBd1xEJhaZDTFfYa3vhfBeO2h3bCL+sF+EvpPSuDIxMmvaO
G0bKYSimkqh6/MPvGSs9vHlJs5GF/LRj6IJYATkxZKSAugG8H654DBiz61cUS4We
NNdLkcM2Aqw/qifcGLHh7k3rXeGUAQtfAS2/PZ2fUoUjnxzBdfhLenW0y7mYTmxp
k5nUq1WYOf72F3k4OngN+bjW4Hs+Qe4ia9KbnAsGiQaU8YVOE9/T4DnPoqVye5Y0
bZhIIZUmomhgpoR2jaRSiz5FXNE5JZY7inmgsbGb3cBH0CQWWVsLBiMQY3yBFb+/
D51F3KgIXk+4ESG7wKEuc9bKvX3fOo0xTEr8XgXCiHrmZtKxnVD1HWA+iV/7nmPp
U0k53ft0f/DtNEcTBR50DigYURqQg2arGI80vuKdQOpLDM4M2mIxnE7D0mjuQz+7
hThBwip0xOo9hA1sJ5iE0Smmjl7WCmlC/hVB1NDvFn5WXd9s5ipRZ3vkuj5jgLMu
umkmYeEvjo36s7pFGwsuPGLcbohFakvkvkdFRLUQobKqztTcjhAsfUzfcTj1hNuo
vT0fKNYxwnszmm1fDzUVKfxQjdUUiA+oufYqLNDITVgQcnZlWdBgHIx8+Y1Gu9Pp
PGgVk5g+Q3Hv8z3mkjPnwPYCNtAUR8TUQIaWSMUs84t2q4T5elc5Tq8OAQEX8+Ik
5+UuTmt+BjB+Kx75DpwOHz+B2vtb+W22c7br47vfSeh0g2zChX9pzMWzWzYLhzOa
rDr6DKty8AFtM4cRspsJyRtdEgztcVyZFPXeXOs/wN3w9wr9c5HzJ8gGUdYPqNMT
xMIGpya6z9K+FvLnWCdFejdoc7N2tMsR1JUhGfSKkr0JULK78BbMVWN2x1QlF85o
QcMeKc/Sqw1HuIQxHwIkxkm+OzwhfjGqBVXdADHqMupPidNB8xFJYpyakf2BhSvO
HEAXgkavT+qJBN3D8ZCfc842NgAUQ0ZF9LULwI3xH6V8wREcwD3AChdiK84jubfp
fO3NK93O3iAg8EHu96Lcxu7KvpN1eFueu8yuPt9lK+Fu+e8wsqFwAoIn0BJXmhZ+
SN2RQdzfWSYO6M3tYE9ZMGOVhPafIFnCVGkgCYFQ1dpqZjwWST6BMCG0zShBmhyC
hjr2/c4M+5kfBc15npF6WNah2TRep8Leb/dJwg4BI7gW0hHH8ZVC2rtxWNuI5LKb
yg7VSLpmuDvOT0GWOJaH7VmEnubTjSaaXPkxhBMV/u5+9QmHoD37bI2LGUKDrBVQ
/gSx4eStO6bVM4m/Kh5Tsm12tUyJGF9UCxCdQ/VGbz/Os/R7v+6LdfT7TGN5DmgV
2YLZgkO3ENjnDq+cvUyhhtCtDx1IeUa8GCRfP8eiljzxCRI/LkvMKhaVBOaM7ohx
XLBQgy2sUC2Vhn3zVyphR5LmbRdc567aYOunOkI5C8kx6t2fuRaECS/CX6ONo9ax
40Vhs2XbScKCdnML3EjTDl9RhQA5AxBH2W6npI9i3Rq3aqFaDqxbU8vM20NuR3iu
mSNv+sZpAC/QBOH+wlGepiDWhSY0p/zm1Dn0PUjngwI1/8XUAXJuJ8Kkmn2hT6zX
M9CBuTqQtYGu/hvW00fsWeqHKi99167+y8HacxRpFDMDfONcfx6ZtzQUEfyMZvwL
ucQAb7OjowVIEls4WVV5gmmAztp/YL1NpRpS4FZUEZolJzhC8f84eZbsTeUHMHHR
mmKdWMOHmXYF/RNyBhfYfeNYhUhRd6kBw1cGCJoVp9EcEs3V8ByxlzuDBGNLTDrd
hUcT8RlM42y6ELdIoCojoLla2d7fodhF4LetOrta1TBFrIOqCwRa+kW4hCpak/pZ
/wUXcnXqdFrEZ5HiO9p5/bcVgbVMBPvSICi+r40twBGd07e0T07xznROYXXDvTI9
hjBwlNvyh1waj5pCqe70FEstvJkheOiAYm2f9Y/ovTRYIUI7ENvaDK+d13Vz0M2h
lIOLQ0fE6kD1xIegslymPkybxth7+3q2HEu6DeBFvjflUebkjGHpArshDFHF0Ns0
en+sLI4TVPjvisXgux+2p4M2u3FygekhMTGUNTaFez8Oe2/7pwz+zYCZd1ZAm78B
+ePNswziB9b/50LlFnGaOewWn3AOUcDd0iPybn6P9yAxxw9Rv72JAoo6S6MWn1jA
tkaLR44/WeZoHccw9TfxiTdHHYnC+9o7go9IG3yGi0z7yjo1MxRRovJXb868tF4K
g3462RvHyQ4TZ1hGsEGB6t5yYgOmoeXHM1uh/eKm4KESJrWGcVetQHuFBka3226J
pvIKctY/H3CJQFzU0tRDjW8qcplmLgayv/eYb6eFUdfnlhnjFM20cCGrjdU8fyHb
vQnfdK7Y2mBrFZDZfC+OyPcsmcvGtHNXVKPZ2k5sDd7/VMz6g/AJoXqH3+ENAN/N
19l7Df9ZuJPAuAM01Pi3M5nz6/6Qd5EUQhTIV1cBiNhPLfdQcUhpuNxckxRlgpF2
D4i65sWP/otxkL8RSvAgI3h4vJ7pw+XmMH0vfzeSMGJcZ5O6xS/H1TyPp1OQVcYR
85oyUdRp7SwNYD3okf3uq5WtQlGjGfDIfw2mw7fYtxwm7HLNY05aNmyf1cX/Baeb
umytkkgpPv4WuMYcE46q0EJNq8ruRXIDECkqFVxHXRzSW4a7jy71pAPNF636pDUq
loNS13xFQSExDrqSa95S0RvRXE297cIsVW4s30iptFslkYB90S8h+W5D76YRun31
URfONmU0XaTqLoDFBNznnx5JHVaskl3Phe4H6C+aWKyf8L3AMk3kte6NUFat511v
laLcWW1TJ9Ql4a+8xEhuwEZrThGvGkkRFn8v/gzC+obANLSfgtacfDULU3J8tHuc
HgoYAa2TAx+3t/92/2dJrkPHDGVRgaFY26UxqlXLxAvQxNiu5WedL0lIDyXjw6nT
VBHE4cSqrWceH1KmubQxzj0cwDPG9o7S0CmrpA9eFQ/SCHhuYiCYvL5BEZHBpDdC
ZWSXbhJM95vtJcmQtXkR4bH7zZoYepV5aJCVZC+tCxjQJK5vwjbkgI/jmnpVp8cy
yq/aFx4T6asEwYxKLc2dCXDKjr6sSD2HSQOUxirkOBlCnqc+dP5Y5pn3GC8flDw0
QCDOiO1vUBYcTlAcSYcdkygE+ReeamfVy56gC196sQ2qlLKUssOeHc+T1eyeYrsf
MDMkGMfbjhXWm7AsFqK1Aa51IfoV/NUlyDrBl3FR+GF7WszsE4nWyHMycLU237yW
hkmzQ2bfQcReQ7+6ZKwU2voC6SEIW6Fdy4/TQ+6jaxW9lhqf1nOEGd9rjFrNoqal
NCXmVSNUEffSJbZOJePjWTA4c+nF9Pm7dgyMFtJ78tDkXqUA952ViP68qLNdxBVK
fptxD5I/qLMQjx5GsehvI7MvRZodW1mdW1XVCH1Q/oUfd0WcpxHh9MIK43RlXPFt
L0zNIKouEefeXUF5FR0Qh32+r7KVlrLDP2U3ymHRTZjhMAQSwXAJHMZxxKJ8Ntfe
xMonDwdTxI2Za0aSak/amVaJqf2/i941qogh10N+L7XeVORtexVaO+Q5EsujbsGB
+WVkdp0PX2SNNAxRI+DlGBSKgNtFyWd92DfTKsh0qAygbaQF5lIyuv/+/qmjyDqR
UZFyubJu7XJhYlVBtAVFAqOpzZRR2A59arb+qGFEfU3xFJIAJWPLuTpMFg/Qd7fU
l1fmpFygFPbV4yCDcneQjVX9Mv0zNfbuKhaDBykqR6pyXxPtTOiRcareyETDvyU1
5uz2jeJ2EEeQ6DSG1b7eyd9UbW/jgVP9OnQ9kwRqggXZN82VWm+2O3f6YUdepBb9
j1mbPJIDd08mvd43r5LfVbqcFcJVeOPDFfdKVE71nVmvdPnN+Co6HZqQI83w/fnb
a+NDz2A1GuiUZG5LUWbvCebpZy6DBOdKF8CQZ0cto3ggX+zr+Fkv026faq1PaFxK
Secca9+4ofGZCEOfjFEtQ4X/tevG6mT68AWQkZiJaV+mfUtkBjm+ajqBvE6BdgMq
Gs+PUprHfW/k2xbvF8wIJNa/NmsHAJ4f51y0AQS0ElMFz15akhINw9jSlvRnDX2q
CGgDC2ORRC3k6dK+DRPKbZmbeT5q+Xh7ymGc3gtJaK2UAjg2yx7RE8DOPbV11u1/
5hpv+ZNBRRytvYAwLJVn17UX0MDahDxQJnhPZKfc2d3scHlKHyMwzagE3PfXyWFF
oT0XFTo1Ypf2zKPxn3oHeBIIzox0U7knzJCvUl/n5yG/3hgbJCVaSek4jwwZf3oS
DW2bwKwoHIYfH+BWFkMkVHPWyuajs9zO2AW+ViY3kQ6We0N1x+TGiG+0tyu0Y36l
nxC5WGLDrblT57G92QKs7/KdprvT8aJCXKmrzFGz8gMnXKW2MwHAPsOAA+RaNSeK
02apRshbfScJwo02VjoVT6Z9GonrsmsIC2HoKlamD04Ueoy1TyZVjQGsQ9cBYixF
RDqjnw93SkrZUkj4PRQ5behF0lcUGQU+yFG60RTR2LKxQ/4itUbZ6oqD/XzjQips
JF4sAdT+6nraWuebNPdwRFCzBFs9NM+o8hQFv/G3NnPaefU++1W8ucQiozlwevMJ
mUqKIAaPXr9bFuWbFhYV6rCFAfUxsO0WxzjT54RRsObYtHVh5qwWREUTwu1i+W5t
9gtoj68gEPsPY/aBYj+OL966lJ8ZbjtC98IzUkh3/5fySRi5vyuFNomNi3E+VZ9C
tVGtFWpN+RwtdM/6ZbUWwzuF6+SXvd84wbAvB8N2xMZ0o4Uq69bMeU4ZoPpRlYvv
Apb/rFW4c7A+wztq3PhmTqi0eOSRC5jNvHgVuY2DEWFkm3VW9tIWSAQpXpx3sSy6
E57LqUSG2fHV1v+QaNw0U2RU+cbsEJPQmgDDxxkd4fjqMKKklt+7G4doHmYtytwW
Hy/3N3myIziVdqNyDua8eTFNCvPtN1iGrpcsOREIHxr9+K7wapDrmmsFEOdNrVor
U3rtXHrl29i7U+l6Z57Sog/f2zzt4sxYuaxlPq1WE0+iVFUCXK73z9NOUwXK5XJe
9HtZzV1vlq7g+PIea4asTIZCRFp3OyjobN8Hbq/vGtNiewei7hhzoZhJLzpMlqlY
cpmtfoNXbbKly51rcZk4qr2l/5rx9zQPuf3sfhLvZsPATJAiOH+PrxBOGFobINH0
b99OzZ1N5w7mc3DEqB4+cVB37DurqoW4dpbEkpZ3ssgqsSnXZbW4IfFma5PUASiM
m+zvaGsRqLRDZDURAFyo/WGRUjQDbOS0qdDfAqrWhI2iHumodxZB3fJEWeWKhXMs
YrTjc211xb8DecSwiqBJ9L84RRGUSHMIquLErlwFE4QdJBm1O553ea3QOtt6DZQd
sCSJE7VesrOM7/RTXsl6w2Y6C4mtCWky/nSFnrYDnIe1+/iaQ7juffHIamL65Dml
5cDCEZr0Oiu0zLhn813c0DKGHt4OgLh+FIPIAhsC8iSgYoLOdfIK4uoa36rD/oh0
VdAsoXdneYCYuSFxM0T59wry/qcTH6SVwoMx/YPO8D19v1lJ2ihKbiKX03FvoTpS
j02BSFxW3j2UwlbAg+dyzvohyswZw5OX+afe12gqbQdJeJqSz3BrSlM4xY8XkRKD
k1x/2ejmN7ee/NA0WxaYhzLnWakzaZcmq0PUjZOAZ5RYRVWqYL5Lhjehe1tL0Gqo
caLWSVEjU2XqG4Iclz/3VmCf7nUOpGkIfYt6IhIJR1DZv3usr8901rjipHyukjSY
uC4Vnf9xUlK4MfbfCfQtfwbwei7JtKrLG6Y2D9ojQrGnnoOZ/KGCk8l9tErezWXR
okWfAVmtqw+PhMs/m1sH4LyANaFn2EvOWzJGJkaYshTgnNe/RJOnETe4yg2zlTfZ
lr6ALTYLe4ZA5N+FMmiwbmkAuxPJKyxKHznABVQyCLuNY18oTsTb3RmbxazVWoWh
eX+y94Dm2yO9y5ScGzdwSgtfLA6b2brKVRMEHC/+TsA6hFAiXLK0cU4TWKC42956
txjUVJy6FPsDu1En0qMRsVB5PxVudyuWt6csFrUUOvJc3tSGck+tEJhpm7yjYxnb
yqg33gSiNQuIzjf62owpFrSqQp0QD6TFC252ycMgVVOBu+pe/ISivffIk13TzeSC
eEGY524aFcLajygKiiJrHU7aAe+ZlaSBiqBqpVg9LauZXZ2ri/ZJJ3N/46aHOt7T
T1Mab70Ed0EZ790lqi49r/Nr38jIc/ItslHf7sbHZCsMwpmXOrHJphE/I0Ag8fua
SNA2SOjpeE9XuJ7akXRjqMXu1dMNBFZwKfDY0Jj3btbu/tqOwQK9Y4kVXyBNOip9
eId5Q3y+HwTQynUCnmduoJNjmRsW2cip0WV/awEqKscNYFk+yy260n64ra8wd3pi
5gP70HLMGX1SScf/4v/1sh7jipTzQnYtC7DF/MvMOR9BplbUP5TLJA/+wAhKzhyL
rwFVbbCsQxsdMHuNM/ESpqlygRfaAjYheMZtmWn+HM6UGVEQswi8uX65dUOe+EFY
6wEpHTBjQWayHvy4jhY1/HAHDU9/iO8mniljjU8L/ryQQqFTl86ESqvb/ROHBqlB
7GOa4DoKeijmDmJ2x/pUc5WeGQPosopbX9lg8LPlzafv3QFV23fl1nws+JAdvTmQ
5ZKde8s/kscy30yxlrbsXoZFJXIW4BZFl8qzXq5EiuuUHtAovLvTPhUSLy8PtpSV
wdmWyodld1IqKURIC7jiItkPJG7/xAcwhLpIZze9Rs4Ur/Ffqs8f6Te8lfwGJ6EE
NhcmVYDDBjIJ1nsa8Nxw+lLSAU/gVUCcqIUfgbkemyrpCoxvuKrzzWSS5JDS18W4
/A1mSqya/xSqcaLYRwSviL5KAPXv1wNTd8huNpqbwNK7YpPBazqhaLbq5Xa4Rge2
cy8/NGgLQOPDI19hqJ7UW3aCcGR6u7DFgA617PQtF8/2/BfR9jS6XRblRkUMg+Ms
70jL1bv4cbIkZFAaJJ+p+YXmC2LJ4aF/TGz40HRKT/RtvUgPyvCT6rgLivazL7hu
H6XcKzeq3H/UJQPaLvY1ayV3mHmggP9aaq3XoRjl4Ffwz6MUwUEgqmqeVOZuefM+
xvvkjrfZB62newBZOsNrriKt4O76oBkKMmV4Xe795GipSmydNfe0i3dCn5EdlN3k
izklbx557weX26Hix03ROR0KnXKxX9dofjZv/kBWjwmrnLKshO1DHJ/xn4gR4H9E
4pGkhR6QN7OUjNAJ4pvMa0WZtQ+0VAJchYbJcIBNOhGMCYz/xErQUPCwNeerpjgf
TCTKROiewtAISNtqLHqifwKDdBmPRQ6xeIzdQr35TK2kmnHg4o22YN4sEeisoLyX
1IipjvSNDaHdbLKrfYvRTUQzbnPkcu1m1RzulrD37zglI4mxUXUq88eEz9U3QgZN
T7D629UVHmZO4fXNzD8P//qI3UEtenT4ny/962y+eyCq9HHRiwY7ouFjwInLeRFK
ItxFV3vHtpcllAGkqD/IPbwGPohBKhdoIJKPBoFJJzIWyAwJv3ZtAYAGeogzOvlu
sYfoXG7v83GRwQ08g6sf15szHGVxYrXDrkkbTNClH3tz7Ba/g8t3E2EwDJJ0Iurf
zqObtpLrVz2cH4HA1gi5ZGc0XZazjfON/8029MAfD1vWwTaO9XUenFQqdsfomdm6
Q8acGkW4myfoPvjk7llEXKxl1eYckw7kIkqxfQWn4oPpXYdXSCK2ZoTToT7BbuBq
c7tZ90zssVCFMnVVSqh7bVosxw/7M6/5nKeZY1v/mmgGHm4LGGIKX6ibUPiBc6Zg
7FpXFzD78Gp9gbNEtczN/07UFyJqWaRpBDEBRXX0WtmS3xinGzrHR7HIzocikIgA
H4gPoDlDMsaCQKoYi8iqXX232Vmn5FKIO+g3SLMu28tA1zF0uaKrwJ6ltEYYMOOG
5TFRHeG3z9ECSBcvfbE0bWuh0KFW7zmqooHKR5Hvig3PrM3KDBhIzqD53qIOGYz1
zt/o8LC3Bwh+TjkTmp2eFgb2+2KyktYcOjbB4f6lj/15qmKUBOdd6Xyk4+HcJeJu
VtLTxoqMjWb5WST/LCqgb/Etib2k9YLo0jxMcUI4gmeJdM1wmGnhuI8iLO69f5qS
N6AnaChk9MWnZSI+Q0CjvZ2w5mokglaht028uIPURVPW2kDO1VYmsBM3eyjj/NYF
6Yd11VbStl/A7Jhwbf79DUH4y90Q1uBMXX88WrSLoKmbaGoiqu1hdkhEVsA9WJiF
NZDdK4uqCHuERJmcskhCE459Y//deNZhdwirbD8IMz5jpMgvDbMckhO5S5+XRWlr
9EdKzPcy/I97xCnZfV+yjRY5982xeSKJ79yS9OBoPRC0zHKWxZ/BxFmRkoBSBvLt
WXZoQxmu6f8jJ0/YkH+m8lLYFRZokQBZ97hrwDdT9tdGcrNV8+k9ARo+JUpo8k58
AwcQBatqKeMwPPPM2mkRjG3pPo1qT3d+I9LWn1J3nIrOn2B0D69lKZDpHKpdEDyr
aOCEw9hdC/w/L3y0aBYm5G4sCA9Sb55Nm7mRjT0wjnDcG/kVPMmsDzzLpeFqwC/w
1KGj5KWzTyyvmhhVhftHUlzoE0Vp8tcBOZT3ozi3P9M+T+fxKZEN8clczAfAQvX1
+KHlkTnV5rFL3qJ4NpvjHmyn5mUTAklgDDMI+vllVy65wx9UyN+xRC3XOgdEKqNL
o/A+dZ17mQeU6JOUX3tHJH/ek7+5S3IkNYAG1IjwdTRqzjbzR9a72kECw/Cz4ADt
u7n5lGuA6RFT3kKc8JD1lGWQGQ9WX09yzhkAPvSaMNgvLWsqr2k6zTtMxCeWYwj7
x8xlD8mYqCiiPg75XqMfjghuyIPJGxXzFjf8h/G53iYbKgi+Ut3OFFCSJ0oAGmeu
BmT9AhvQ8GDmaJWAj1hLF9/cYathD7cDJBst49IScN5GduvzHZxmMfQxxpdGl68S
Ekf4KxJF7sTzswAfuGLGtHNQi1SpbISkSxVOIrV5HTfBKRjkQwdf6ZMBjrqSUiSp
SsgDJ7t92FsSCMdOBpshW0k8hv1H4PUObdXe9u4hO5n2N4wPMLqhNZQCEMCJk/ec
+rNiH/LsWsBdE/tc3/yv6EoF+hQYsYCa51JGbd8AQ/fxD5Z0/m9DRGywZVmsgEQO
TNTGbMD8rZmSZAJV5yeUO1Yqk2sImM+vaSfH6r0vnNA7vUglFQwq/Rz6YIkuM+CL
6cUqbnJP89uB48yl19RDkxPMY/zrVopoAf93N3AVBu6o5l2AGnQQZbVjBPHdxAYH
oxE+/nem86RHzT7SKtYNw9dtNVhucN+A/aIalu25j8IQEtNYknLUShKT+bTXxKGd
npYNMtWGpJ4oTeZBsKz3mXVBrRG+ZGOrpFEodJzrWUAY3CdxAO9CjfvRpCHmk/SD
2XgLc+6YfZOEGWF4FCibUB9FC2kre/OwfnAdBhkJzAg3r7cQw83iWg8wkKjzSgZs
k1fcJa/TvEIgG2hoxvOpbKzU+3XMMRS7uMzOqcd3qlfpzGjVoWpaq0tzrUm0+abG
BQbKOtdpD00PquDrXX22DC0iQv8uhVSauLiMegyXWcPJAUfBngJogaT0g1ZGnAwn
CaOIu/9SYJE1kUgL+g/kIS1dRfANYRRlpAHFSC+uSerAMPC6r4t/MaKg6nfFNt2K
5CatfuJ8QEU/dUgyOa5sVEjUkNsiNi/GdSoH1ngWV65QC/nBN0iFfYoe519vKOeb
8dhvjB2qGBvsDJaH2grsSfRIpqyfsr/tAm1nwWPGNnQwGuD7l2rJM6rNQvbmGSaj
wMHMHwP1ovP8KPH1R/0CTZU8RFLk1NQiA349/S66YbgjG092pPVn/s/nbIVR45Lc
SxP8xh8o3s/UaNdX2bY0p643kqxLQsfudMBTxa9tAEa6xMrDhqNhhOnicKLqrJi0
bGJj4M08YvR4/VQVY+WBHkChVlEa5hTV5SBuLKsX7oaO79Ulon8xjy+K1qTF7z0R
Yf9FeLQJ5W+uHqw8DF0dTabrzlAx7yl55XpxLURpbjyVxwPAc7alnXlMPXu/Q4/O
p9DRgtXXKr0DbMO2uEPOH4tw9Djzre7jk1ltv1vdBvCrBJJZ/M8+3PTtBEkkE+MI
arDk45zYx/uwWbgg/Brxw0sUWxBYJ3NeRlHzmaG97hJ4TGCjvf585h6zX8afSMs0
zmDcS19oIHEt3Db1WvEOEAgpfUYS9AgVm75zSvZ3kcM7FgkM6dkdynVHZZ+DmY6n
a9C3IhatNd/Yu0ew+8icZJM1YdUnUkHdhRsniTmGPzYtNWti71rzBT4igB3hxjvP
9U35iOaq2//iwDW7H6kWyT1N+3pI2ncq46g0Ab3y+xtpb0vg++Y9E2bvRdGIP50e
050BWnyBwf1yrijlcVq8WZoo3YfhyZKtrRJ8kDeFW6Dn/hFGSMjcMUfkytHO1MZ6
mj22cD7DGP5ap9zQoFORmklTUMzmRlqdeMf1R2nrg72KcJ03PpKbdsaNv1TzgO+A
6n6R/4DkGYm0FYC5PV3Uj5nss/2d2csSJkaQVdT0pVCWP8kGsrM0Oo57zcNi8/pu
9w7J/aoNbuhR1xzNo2+XzkysK2H5Nspmz1eMq7/8Tw0y1DTiO6ZxwvqVVtwBIACX
7YAXGchwxl/0Js9TSemX51bga3Y1uAq6ksgTpz/uYQNse1Ew52Dw0JSfKlOzZ+KL
OXT8ozqKyA0ww6xGhhGfxXbbZnEk68WSkW1w4PAG3iy4NUfs0XoqzSz1hJBumYAV
EK3ygzBVutwwC3qWUmnGzrRi4z+ZqgrRI7JBbFSRmOD/W3E6C8yezX9eyCPjTDGl
PJ4GoqgDEPGRUk0Sx1fbcNuzh+G8JMKph7dZV2b8r+ZuY8tjp0yp5l6ZhPN8CnhK
klOD9aXXVEoKPnAjNOMAEfFih84qPNY8BfscCIF5Awf+26Vfp+YvpH2PJITa0pYg
lFDGMNQnQcF+YV9hQYYRbkmdIJOpJPjVg9L9P78nB0QBSBqQBc4urXIhunxcqWYR
8QY9fMRxL9S73qgHcGtmFHTpS5XNNghqKSrK4MztssjYubx1f0h/V3PxkY3PQiux
w68PE0f6e71M2qAoZ8GUvVJiVwkWhldJB4mgRLznCAcz5+yPFii+dBfD2VuPhM40
D/WjpWa8+s/Jw6kf8ciz7stjY2ioVfTvLAa+h/kP7dxYTy052NuxfVTP6+R5eThN
sRX6gKOIwn+UZqgEKevJTvag9m+LHkaLLAGS7stiMpL6YrddQw1P9flE9sEHU6sf
70d86EhiLBz7pZksWf7eT2OieZHa4M0NYXaetVmHbq3EJIJD8iQJd7pwhA5swB33
kyz4a3kPkfAZ2V//wSjwf8IeNrtC9jp0c0KKiKBgqOcEnzdBr9J8MF80XaMiAq9b
k2A9+Lny+DikYOxtRwZuwgTYsqjnktctMTFN19Is/h31Wqqs+NHqv6nm9vJuKDJX
ulZL6MUzXxsRVreQ736Otq0juXO7ZkvcLk3RJwpV7U9Chg7VnCEzUedxD52p5vjx
IAuNKHzoa+JBUUaJ4+IQ9DmYowuZF4XJ1epbcZWbCjLavdFMU3VRW5/bimYzCXOX
OB5kuOdey05F1A/ykX6oiW0Otet65mehbSkI0DksLjy+1P7XQRokEhZBVsW6Kwlq
Xi2YJ+PIvANB1FfcQrxhplqvSRCDksCPMF/amlP3BiUjP3qE846lbiOOLQlanepH
UxxN1SHFMK4xAnoNKT9/7Irdv65oAYu3EahCHYtKkXyTANDu0uhVrHPSRgOpdKlJ
sVftRwAKeqlkeVZJfOFEE93+yOxVLjuKHS7Way5tpa7uN2kUvuEa1Ht+caqUkLPm
ikW9lqF6i8taGOMFyrv9pTXD5PtA/zqjs8MHLoyrHpolp+F2Xwf0a0RM9NPqDZWc
0IUP+XmPc34MAEHevAspssp03c5Gj1E6Y/X20e+AGCtyqJ5HK6Xr+nTVu6UOg48W
uQlg0FcyOk4UgUYp/l85huaxiCDwd8Xe8ArT5Q0t9LtV/UETvYtnYrXhy7CUkoeT
DHsC4T8MWmnUXAuq6mCsgnu1Jm1MrLebUp6V2jXrYdtWkR8qq9eIsiC9ghJonb/b
LfvktcxFUqwFC5284bTC84sisQAHS60ydTPKrkE9sIw6NlV+NjTDzc+1CF9XaTw3
cCp86qxsyPRQ7+7snJCLHfumbOP0KoGS7qXXg5h3RCv5ZpR8GAv8+UhEEsSYtPhz
avjL6srcuT4WClQ7q2u3yACqTtYGIMc2XsU5OVqLIR7IBxFv5EwCyqPD4FbVxTwi
JC3vfw8qnS1N4jZq5aeGe0hXQPfQtG0m+sFt41XY5MxRWjbdol9NyV/KzQIm/NAw
l8MC1VeC3QKb34jb/rxI4zq3Tl8kKmFObO5OuYHAufCuD3u5hjCuztX5pUE+CP/b
FkTzm1+bGLphK2FPQiy/n9IKh0/3Tf2wL8dVn93yDLfCM5ptHkh/H3/gBayZgvEV
PlPwXWwHg0sC5u9DQ+vLLiz/RhgWPv5Y81Y0DLiCpPIAx7NDmTCz/yL9VEike5uQ
8GwKSK90+5v9UJF8LC0JSkHKgbXv9ESneewnGnBe71SVrccXxNkKO8DUTTs02nbq
6q62HU39DwEtR6LwMQYq9CNlrPimumnOLSZPII1BnjJXChgip/c4WWLNgU/CqkA3
60I+652pBfrFS+XFUiilRxqSAdOvMq4DSlxKMrtydVavrjnaH423cY15glD3rD6f
E6my8X0GduUzQn8fMsvEGUEoeSzA+Ewx8w+g0enLcnDXid5XL1aWmf6ZD4Zwog+E
mrdp1N2pvmQdV6AhDlvVfRBXqcGcXDwAN0Mq4kfxlLi15IHU+l6n3KwuKI96N2DP
wpZGRYmk0j2oD/OlGlGrxg27cl92vZxhkg+6kffrILUav35udywVvZbsCDn2cLKx
WBdj9SO7gxrEtM44ghbIOIRX+RsIszButX2wyTKGtfMdQoUatw5Kv0weZKoUfVzN
6IvS29RJtBMBj30fM5iLh7MVJXUkLv6o2dPiQwHvqSOUmiN24PySwQyWZ/V3NVjO
7jynugh2EDp+TwZORLR8l6CN/yevQsZLZAcjfDs+ngv1ywSrotbLLV3Emf25tYEg
Mx4iSkKhfgCY5yg5VbEGiSXybIAo62ul+Kr0aauWl2GlSA+T1/k+bhKpsyQCPWdR
wxhFPf5/CkZAs+VVFBJv+RpHrxJhRFyskaDHYXYb5W7jo+f4A3s3UyzP5SMZDR5y
3tqXI+jnVv5d87O7dv7Rw/kYTQcOsLUHPZXJF0KVG5/Y1RiGlv1I84hXIDP0mT+O
8gz+YjghJdLWpa6H/PrE1Lfv92zuNHABpPBOCdE8uxl1CS+rhLeOX0zb9/x8W5DV
f4utKsCWk6GYiJxlmIJgz71M/Z6hK0hjcP92MFue7gk2/MD4zi+pMkswGC+DjBHA
MGOe+SSjjWeH/w4UKgWfri0eMZCl5Uz9BLdCuT2tI6ibna3ew1O0BcDjx4dnwhTZ
7ngza51kcMJtSIdvlz6mQgZzd4kh9W+gYZuPSAlBpzFgRkZlPnnXWbHS7N3mE52H
ZGTHJwmfjP99rbyI0KBKIE9+4qboNzXwJ66/HpYCxVENl6UGe36eDi89J4dF70mi
zINCRKIgoc95z0TeVKwQhNmzt+KOWpXkunMMmCHzQjVsXODf8LD6TEid50aYytfy
Y2AoqqjGwfJhtfBC53SszzsxDh0f3v17pwRjeziA54q1qjjDu9t8PNu/3mrnY/+y
6U8Sk7JNLCT/YhaiifIq3Kb80kw+ANPi1qG3VxJOC6or9Ajq1JQr6yfzvjjy1pNu
TfvGTjARu47hFgGAdkvXw3ctLy2XjAO2A/7yj0q3ujTRRQ2PDEDXTUxOMQ2yz38t
C7Ig3zrh8nX/hHt/TrhOETHLfI3sCt5AOBNTHHD9PN8uhWwHARU2Ou89zy0OcBKC
H+9ci8z1TCZG8NbrXxAi5g4nksPPLA8X6G+zfexnXgW9bGRrdF8v+ymKepnuJyY5
hHA4FQh/rjgv7INfxPhKu5N0scnTzBNTqoh9X3W1UOz+zqEYXZfwG/pJeMpx6RbU
m9IOzTre7ZEm5mFN7vPGCq00Z+vidpdj91st9JMQr02Sgbi2cC/hRXxAWoI4HFb4
2vcoQQsJjAA26ZFykI3Fc7/hV3zgoe3tTmdLUoOkryJG6NvFQVlPSVscBQhQx+gZ
mTrncmA7aVy19UaEPPAOeIpVGr4gPM2uVWJ3+4Glg7+GfOkPYI+UwdzP3Wem9yYo
uMwQ+CtQ9DyGNcYKjShWx5Twd7XJohibZ38OTAkIzwvZmYaD4dXnwG5hua2dslDu
NVjudogISdhMan16qlDenIr44/I8CP563VSf8eU05nBOBiG1Gc3guPaNkmYjClDA
ysD2W9zFQSVk07B8vKyo1nhU9kRmj+qxacORbYdBCOMX5q+6tZJ5iYO/yR5Z47b0
l4mJbsIziZMPQ0z4MZxvqmtvD6ft4YxuUTspwzkfIOiIsyosX0ct58328Weu/ca8
/umgEPhzRV8T3JhMXM1d1SmEiQK+z+8QOp92/WlRYRF4rIuak9gTVeUPz204H8bI
nxfTFv/cDLKuPBCqj2GozKDOm5S5n8emoqjcDMWPclXODUxT7EEmX5QgPAAmri4e
JD4niuSryPcQm6VGE/w4bGGX/J/llFzFChqP32hoDfEcWe57hKVlk5TJY6eV+W8S
peCqUpoqiiqeOp4wvbwJMzhVIAnLMaQ/w0Igyf8ZakTXGb4mKBbsVWHOBSUVTPGU
ynCX9HcvDLKB3DfG3J7kOqoZMcJEBfzWLLvjwLp4QlX5V1V4QSaD7iWXsx8Q4GA9
VKEaKo09ykqBW5TnPxKOn/pT/skKQwHGbznnV9frSo4Vf8TX7JT5nKyMXq7OOM+N
22yMaAWDtt0EVDIP2koFe9Q93Ms0NfmEorXGAmaEmfaOYJWfbAll3qiQ/FRsiG0o
rEGGB3bJVT7LI9U6FByYe0pmCire76j2RJ3WOpLw+yk98dXO4YBYCSCjXcrbpqOp
7yCjWglQ4LJcWG5Lst/2bX69jH/6QBzhXdEztatSTxVw8S3sRiLOrRGXbhc6BL5l
g7quHAokheqKW7MvgzW2PPWAaPDf0pCckrYGDowrReh0TQu9Pb6IhtN+k4xF9CqY
pqcIELaDPKdvrk5O6lhyPBRhQDDYOtVDaKxivd4aNOh8YvQ6pPVhrTCs+c3VDWJ3
doMZgYMFqobldk2uV3Ua3hpyQUaLS/MMqtwmpxF5QE5oZ/nIDHsSpV2u31vMsUUf
9fFekHSvu4As0Jg9tcNdDn7ylOn0SVBZHnYYisb/vkwGVO0Qu9L3mcQ7v9M6Inop
IEV59d3ZqQ/ZeX0skRLo1jmXgYV1jvLSoEXeHTAFz/iWIvNQPB7AV18wZR3EWiLE
Yit92gQonlgA/lIlhO6i6GtL5UqmqxgJefSDg27lqBpfQfIU+SLT1CP18JOkDxw1
bKn3Rz4lMXTTJP5yH+HgHNlC+LwNbuZbrhzSqjaZkW66+udsjPzyoYF2CZZyeGmS
EtJZB0g5RXQ/w//CEKn5jp7XM1gB0ZRV3MFHt+GhJVRw8DsSZksXFuFN7bXNCG8x
b2+fKGTWBOGCpXodm6nIyyG9J52fCgk2HjqYO5YPewUlKZo2w6zWjWbxF00LYoAD
5jVtb+8MjxlrBEliuXFgv/RKy2Jt+y6SeKnAQrOCn4BXdr0i71KEIW0E5/BFA6SF
QNCgbLnrUSmwMMkd1FCH+QhQL/TZ35mvp4c6HbFJk6UFJlz0M++qHobUI4OggJoc
FwIxIa6uJ4wYdRWxJWB1sq9KlLkigu3Gvy7AMD7AmL6lWaCkBc+v3AuCn0lbnId5
cWMHq8WKRHHilUH53931fmChy4GCLgOsYCkny/6q9/GQbGen75h0RR29xJr4Wqu0
Y2Oa5T12fgBZdkTb4wuOzyn4J9So+EPeGmCJQEUJlTXIPBeSHtyYaXn1wgRf95YA
ssZiEPdJiQcj+hDEJZxgc6YytIH9LoIDoHc27r0O0tFoIWoiNuGCNea4d7kWxQ6Z
yQsr9QcMDImqrzJngI2PiMm0pm8AahYnJRfvXHzl5YsKYXS015ONyYh/jLzxSYrp
kns5To8SzbAdwd0OewTnmRYsg9ZC2GCeSfHKhm2EziWyefScLLxKoBfcPiPmiRZT
lG5T4J44QO4nyg/FUGcsG5rAZKBJM+pIsxb1X6bXdID5PPvYv/tfjWzs2IRtZ2y2
0MPcAA3Q9j8hieNMxnFim8A+HvrVW38+3LWFSdC300rXhEBYv7Wb2P4b8oWOMfwP
6RfQF6K7q/Tf5Imerh1tEv86BucOAWrlEBHKf6Cj3gRssWwS9+pUCqyY8ChjCIwf
eleC6q6xB22oxjCr9mZiV/LPkHp2tUA+cvpF1aQV/d9gYslCE70KF0OgI09j0P/R
G7FNAdfMWSd1keapZlJP2PqNugZvP8xCyVxfPRKhY28dt0FMy9sDmqFvqgPdWfHB
xnfCAP/Eh7BgsVou4O5BpB2RMYjXj4m48d64RNThT+wK4SYZyVzzjpT1KE0L26Od
2ujD1y/bDBCRBkm63374MdwaxMVVe01xELZFEtT9wJQSL6VqY2+dLODWKiIH8VFJ
ldGwZahrziAWoOcpL055RXeXHpzKvNmg/FME/ZkWIeUBBo8J+I9EQhlANSHL3Yqi
bbnKHKAJu0D0klGmTeyeQ1mAybQsRj4koxlkmJDADJlyxI5giGDjzB2iX3FTk0x7
Z5QGLTmf8BDgefYprdXmRxgnn+LbVFlvVHX5gW95MrfwnApkfDS+BaQXjWX0tvsr
rUm8RceDJlkj32F1gEpnkHRKPe8A0pQVyqL9C3e71WkrfE8ojYoeuX1eXBx319zh
2hFGU8/6SfcV0YmAgEQlBLU3ELImIBrwzIa9upBO5GV+xXNUIqunGskRu4tzttRv
QzLqjUbuw6dhR+Zb4s+rfbnG8icUC6lIOf2n7djaO0hu/cUaQsZ+47trDryQezYF
Lry8SH+Guhrq8MHTlDTzua1WoPXKVkQMmfu6Vj4dZHJTMyFsTuZtBiB7kYzmz9Mn
yrm7Aw9LtXJNMF/QDe0arvwglDJWc/d9lFTuiErkBVtc5XJOJ3qK1o304X5ha2tc
G+d0RX48NCq3mN5djNSLIcdLy+gTENKhBuT7RaZnTZRF88C5fLwukNvAMfMakihG
ZzA1YAZSD5Z18sSZ4QXQMY14mNWLa8LYFfofc2RP4nznMCMxT0owRU8DCJQD3UIn
eEOHAzRxckrj8aiQi0n2UxuumhSx1UYpvkwws5w+6T6XwNaDmtcBM8+7O0TF8sFE
BPlQGCasns26XX/uoPpiGW7T9PhZSGpTNRWBaMJaFa47BvH2nMqzoMhWVU0vOMGK
XleprJ4ENo5vKA9uFQfSocrlyuydeduVezMHqzi4y9gH5AQjzjdVZmRcxjMJie7t
Y3ZK2p/YqzHdF1YCNddgF5mTz5s46ytCf8a8kehEpHPL2OEksfNtq42NShjZPyW1
+vu6DKakxHATPr2bDsidKal3G6UQu7r1ogRaZNTPwyESkAc0ko0f+lG+PrfRT8ik
rYGMVp4Eqvkj6xeX3SFUhE2sD9OvULRXJeN2cmnnT+wo+9LLHVyyGHHeTGizJEzY
ZNsqDmxErglKYGEMVTkxPzvyDnP+0p33OzUDIkmFwi1Q9r9a2+yvFK345dVkiu/r
TA/DiZm0BBDDWNPMYz3mmBLdWeqPir7df5JqPkivkvou5XJgDnQCiKoMthmSXOID
cGVJVHGWyUTpEdtRu789Mc2JOMdPWMYhv+a8Qo4vFuqa1cjwaS3c2Emf07B2ArJz
WJNnwNUyBGCh1Sd20SUTbNlvFiDyBkGL2+ir65qmBN2zs9GQsEEgOWaOUPweWn9a
g+bXsLOZhupucNOnFTGoaFspe3WPH4fWwP3Rnre06+Jhuvte0oNIHMdtYd/HvTfc
rJEF0Xypl7HqjEJakaM7P7XW4xwBBJUNAn3AfrWR5Q3nIz/vmescM9E3putPeO2v
q3JYiRtDPR4ieFVUHxf79XunmJiMEPWctrdelw/lM81vtU+XwsE6s0LUHvBXCiOV
BllN0+mVxlvP7WnmrCkRWQ3bXBn/+sUXqRdSRwzVeHXMQQxJ9DpvIJdNGnblPVJB
tpbaIf6lvzSOZnjyCNE+E0VHn1dWpRwfcM5ZaIjTTeI+UpQk26hAeZlr7S9ARYjW
`protect end_protected