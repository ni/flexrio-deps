`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7824 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1wB2ShNYedzmkmBWjqK4Mg3
8iDfXbv5M0vDNkp8sRs0MJKXmOhrmn4VoSp2HGjZSWgo7txfgaIW6DYj7qD1AS2m
BicfynXt40+UNkxSpzvWIuX5Bvd9dv25ibr/wdIzNxS0r1kPNhtW1Rzw2EuW16M9
ImOHTJoaFzMIZv8qSyrP9G/kfyiWl8ndSobJsZBl6ry7KNsyhSiAGvL8Z1T2CksZ
pl96OsZRcsTSQuY/3UurTQBjgdo/KgwC+k8QNC8ydCrKWNQGTdyAao8TYjxQZDL5
42cKWRmY6CRBEnJi0t8APwWTW8Xd3FiabL9vJHB4xOoZC0YYH21ZoaKCxG+QVqGA
F5hucVTTbYMaTU3MSV4RT2G+rtAwPK3CYoW1JcjHekrqhgR0LritIBtrZp2/RTdZ
N/IfvEk7hToFUF8BGT19I7kdwNGyHlTOiLAO62czsA8KlQvbn5KUhHBDSg1UZdr4
5pXg7gvLu7EqI8KdBa+FfwUJNsWmx6LzZk4LkeJx5FqVbg+vOF3I6iKvRxoFFoGr
M5uTWL8KtDfqZ7ZYYrKB9OXoHl1G/iIL40vZya3v9C/lqAh4lDCklC1SJDKSHsoT
Kw6PE+PMQ9xc7hps+82RE/C4Oj/modPI9925BXUFFadv0xo9yPzA3pxfKZJviYlj
25vzqkqcD5VytO9WStghzGmKMGIWwfPGLpsm02wRV8TGx1QE4QssUtrg2aHqWeJY
inG/co7DnMCQFEWW+1aei+b+PTiNmWVcxtbdLZ2VZyu5Y2kgy3pzZXWqj4W+2Jjr
YxFXxI6ft3f2zZ/CFbkcy+MLH38/COZRkva6IFhcfi/b7L6O1OO/M/Z7+j/vN4Tp
XoLfl6EorC/YnjejZtvDkomUqcepLsfJLBkHv03P4sH1mOD+B9WeX2RqSGpq5Qfa
SpQted5YwPCbe53XG2w96Tov7eQuWRriWHgMTq6SNJtLCdKNQoWI5IHq3TNlH26D
F+81xxsfgopB0uWq/CjKpvozRo7NJC68eR7DN33cWqg9Ve4vX6AoMDcVu4F4g9Az
Lrqbml7DoArDY6n1hgD6sEa3seP/TKDkGFWgfl2CP8Cz/mFE5LyrwqkcKNJraGqO
mHdQFACtUO6i1bsKHehr+0qN5X1+chtSJCB4ZallBGZzcrVAJJRA9UZLqiHcEmjR
oAw4Q3JhGrOaQOJ327TL41JuwDUJs+ZDpuq0jR+WAGTyJsBoyraan4+hhGb2qEQX
ySHsG1KH3ZNIVdOA7rMxI5f8JYz55G8hmynq+wcoVmmvfmuujeQVfGICh5y61uIR
Q49WajvBQznMAOh5U7Vw66Mjg8Hy8dmwGhDqUzhQ0ADjdgGhuoMw/2Dg851S9nfb
EE8n0lPkV1oibeZpFVZ1f154Sts1y0ekyDq13Gp2AUQ69yeA1KN6IBBaL6Wp3fiC
MaJtQ0JwCd/iXDoHIhnr7AWJ4rfWCrYgDKocgnLavDLOFBA2xl06a3yglHU1cJ+e
VpO4pKfsNdzxZ6KFh87wwO/DpuMrQggw9CYvIqdizonh44S2aLxVjJjNXOe7fx0S
EFIvSFA4gTQVWqMp83ZD2+pUep9F66orDzvVbA/20/wvnn9Tq0zXwhtWI8bbWYgf
JQ0YSS58pTRwznBu2z4Yr0HDk85H/YXqbq5q8CDwEIJ+iiHuk3RvkUWXUcxUehse
44i2Ji0gpeeRLNPCxswIdWEaj0mqe7WX56+YZV0ikYqhOnyG9o/3Y752+qqA8jRB
noO7NM80pAVDQzifOHQx7oPz/83j6Ud/4yIimLV7+9Iv6cENq+SARaShuslk+gaS
zRLmZYwySCiMBrTE2hWx2Ax2ZhtgRjS4Yna2K5ZVUBqvovH9v7q1e9DLe/RDQVUG
TsPO89XVqiEc1+ak9GL8zm2EhA9wIZF1tfdHosRei4va64EigoJ3wIdfpyongMAw
aAwh9DLtvAJWddVD3Ag+r6+ORaZXxoKTsK/auMTzkh/cLkSmkwy8YOa5fj4OsCVp
ngv4HCW+J9JGwCt4QYreZjoG8xKZDs4b6CkH7HPGyhNw7n5/WnpLXJu/tK51CtFe
CGdm/+CpVFadm9vLZpxk/XJZ6Yu4JbKRLWM/avOAZCVw4+5fwGTsxG5/gDpWfD/i
vO6Kd+H27r35ZtACg8LvGgCMIu48kQR5K62T7wYPZSRziml4QfM6CeEvhoKUtvhM
AHUqGscMJmMFHO/NM7KESHMz/rGWHxB+fQbzGhhDZhprrsj3UEeh90VgevD+1aJ9
We4fdE7fsKXPVC0lV6vd6E+SMRd8WKq3rtk0JBtrJsOfKTi36PR8qmkzbuopuUmh
+CXtVSb0sgvudshrJKX3tDuWDxgVYULCOOnNfYGT5GCg/nCPJxV09n3KDYXTZFrg
oTZc+p2xJWeEb8pTg4I8DF+l2/5Fgnd45atNwyDqNr+0fXFqL1BuBQPpZqXYGtPL
HwaTfJBMa3WyvLnxzPrgA5u6fFnBz5kU/V8NXZkw188I0kVsIf0t5gyRrQZY5xN3
liKGRON9HtQdQBv3SR1uLJ+mEG6hODHfWN1eHCJ0dxoN39Fy6sVDlhbXFMejO0gO
QF9+IpV2PGQXGTyGKmZ188VbySvfT478EFWyvvArP1TbAmTlqgfEDx9e5KEZmgZR
A3Br5qpIwLbIjp+SJiPLGLiBIk8t4JCf1tMXeHzzGLYztq2heyDJvfj/3iyoyVtO
3Vv3MNEbpfWQw9OBXBIVbB7z51V3Bk1LmsTosJxXx3ZabOt63wrPrCJb0tYrLvR7
YEsI1dripbJNZmkWp1DPAJLkz45h6J67KO8y1FAVdeXYSi3P8/u2M+9wwygmMhw0
E+hjAL09apzO8hLEi/cv1lG2xiEv8yFLsOVEoWL9cWD+DL531DKZA09iy0rxDgWi
eoINFewPpaCY56TjkPz7Az84jbTDe70h3od3YCmuwYH9o02n9E6IEML3SDhC0FSU
llF2/BBTnDngk9M73CY+4Rddi+0JLahXUzkuDhs764pQpCOH0zQ+j7vajwIUSUPy
mlcyw/Qz4JNvyXpbVBDtqXCgggd6/ZGw/c9jdd6a9MUEFPar1XS7sm/de2WdQC1E
MCrNxNje5bjY2cpdk83z7tD0PTONVVUQfOIiZQu2EDg8kuw6kUKW0FDz3VbIcW17
N6R7vdQWbrncsIfcnkVi9AgvUB1Zew34y3w/UTp+scmyWWRnxXZpdAADjnBjdTkP
GTLzOvKgbQyQ5iCtZcDW3c36kAGnjVsvh7z5djTDV5P/TIZfTmwD+9aQZFkiwCgU
q4bQlU6EsOexZZ2U4r4kNuu8nUVLh1J02cbIGyjBNTp8CsOgfAm4xzKXQotYQUtg
8+nOeeWU5UMssCCkPFUJ79OJWp7c4559BDLd2KTqg4ac4ILCZcq5dE8UK216Rc42
prBxCHJMWFDQ8DiNd0ay0U86iAqNp76El1TxrrlFBK/c/7O/SuPbuQqJt9RjG8w0
iiE2zzBfJlNmhTbNiXmeIxLadTnswB7PCcCVwMVI+d/k99Un4zP6Ex/Fqdx8zzv9
Ru0Ai96cwRALS+IXmcTIEZc1Oc10j1BFxI8hOSQkOiT1iuzIVr9jRuz0sOIRhbSP
PPYdOXQP3lJInxYceg3zeorFG+/A48zyAzZGRMM08xm3nNH+ktNGjh7jxINebYwE
ka9nssG3k5ebEhz79uHJPpqu9convVUxGAhA2JgOMbFaXHfaqQIJNyozu+n2QLb3
3VZVhZ4SKeN8Ryg6xb0+wSSLhqSF6WTFexBq12tlYQufbmWnXYP1HknFM37Zouo7
PmmS9ZbJihh3yVRazGLTNEeV3Xylz0KijhB3aKpaG95XG0TlIdtMFO4H26LjYf4T
m32LjzrsC1h8wcWVnExU519JhqDvXzxKXIlKf4WhnRXqRiMStlyCn1TshCo/eUyA
k+fY/0ITE3FmTAt6yIRhKJJyH84U3i4VqPwXL59P4cRwZsXc6aghPZaUVZLrIlnh
89O0eIzg5iR46ddusWKEh5tts7figElFMRG8TBpBjTWqlaSRpmIeDAEtdtxWFuXo
q9Hnit3pjG6Nm4gjBqsM0u5Efa7kb8TgJwQyQu+8lKXUnwBgwSfh/gZVGc7VkKHs
SKTAGZmIsBfLxWpP35arUtlWtYyNIixsY6yXvqKwAiFK4izWm3uIiwj5IBvb6cYU
bEbNUHFuf5+Rlpz/lf2DD5hPjOO1HAUyZCXGV8tor7khPNWealAqCRcGq6WSlSqE
IrKgTB4VyxjqVdLTpChPGQhIZY/+TYhQFLiEpMImpvNMh/2hQO6sMZ5vfxQ/+XV6
E1K5A3yOpOeainNepMQPPqbxx/dieK126H0/aaqmqnKKqFwKR8LPk387Evwagy+b
uUlY6ncNdmzUjwH21iPSZvbA7BqwnQHM9cUGuHir8flV9nnMEh2CVPw9XYFQ1MX5
eujryzkQcxsGq1eGLDNm07VAhQ5S63UpQOROdKJRSxtSRhHuX/LUSriQdGUwUtTn
IT5ua2DqBQ6E0jlPaheH6NQ/CDrlqDfJUqVCh+edI55i4k697uoNhL1ZkLjWMxE/
ysY+hLmuc5vGY3aCsj/VjhTxc1NUPNodk7n+MgzguA5FM1829JkymCZE5di28Dkq
3GWNCSXlF1dfFl931waDyGaPxFGIz2FFex9FdXZ9NuP0qP0lcQ/SJJwv+POUI5Xb
S8AIwQFozwHKpxNfCyYrJJy6cO+Ex+YtsEnTVVLjoZdM3xYNajZ+/E7BjS9p/mk/
GPd35wzsKT1eU+sJLyjwztODUQNxqJcbgM052hmYnHUKuch5hoOiXyzMYLXkyEvl
CWHufiNPvP+LpzA4tLYcsKr86phQdJKaqEofs8jwjstHoY8Zk0dmvWdPK6v8E6jo
SyXoHosHMc5QqUXHsiTu6M0jkhZmXBt20AffLHMeBTrSOR2180NILdQ2QVIIWyNl
kSMXidUtSdIdtiOx3iKvwxZLtQF8OR6xEHErgA3qAEuOSLXKWCNLbg+vCQeriFJ8
n34yLrXomUnSAIgHKh9fMjjqtvQpPeCTr6xsJ+iW+n5M1EoswjHA7N35u+orF9dK
gmJAtQIuegyrK2MWqFEftrO8axgLZgVRPPfnlESFqNcZ0hVmQE2+rBY3WfkFXCzZ
zCGK30i2F/XfcmxeOJTg91Y49QWTCwqX535fVv2YJc/j5g9R8YMXGqO20undSbEv
vsazv5ffkxoDCvyT/r0rHp3v9PM/SveZKRI2qUff3AfE5la/BzN5EeI777KriOji
CqXjBYt+nJE7NnY7t+cvHR1TwKwYVtSKb1ECcy0QU453mjmZUgVEquc2YPKkb7lT
27383+mR95S4LABp8s+CmuE/YuTnz4bZ6lvgCMoUZPVI+oVsMVRT01j1XTcnSL2I
41XqM8Wr5Wh/2GVX0hqn/vhrLcavzoITmYUsChdpbeXlswu+Rmn91HMcwpPq3IsL
HW4kJW5wH3XBbCshqH24has54i5l0aMWnEz95P0VHRjEAJSzJNFhDLbwJyzQr8tG
/7NVpdL5Xjlq3Rdf+iAJmwZ1nhI9uqBEhBmDop7tWcNayR9XQWxp1AYN9wg4O6Qw
mvQEfZN6oVhGtQLKGzpHwW21cC1bZ+FhfYjy7mZwI96+NDMDPKGojI+o1eKYXaEC
CxzLLGBn/4FQWCeaVh4tCUzJCu4Y7NeXmWixXkGleRQY8qepY0fcbrb1d0QpBAzu
2aq+KyukovpjAJU49sIWNIo59SCCK5wJRMV4qckF15LQB3ZJc1BMhb7SJGk7LRdz
eUdxLzgD2p8hPO6hqF5Y/mph4XWdt1kT572b2axQ2ghgyW5mOU0yWfTQKfX42yrR
3bzUxZp8n98zheIKne46vLPWAXy33JZOFWm0+thp/pUccQmupxYDFhbGp/L0j1vF
K0n0WYKlteGn0lgd4mlwqDf0KfyjkHNuuMWDAd+Egh5xs9KHR5yrN4MK0ksK/PS/
6uNySl+p0HcDKcAnSBle8HI4l3weXMQ0y3qXhlwbMVOY+l9FxhATdfqVCEUnLUeC
504SPfKKl7YS1I4ubjxgvHA++4nFdpN7edFSnzidu88yRy95NalqWzffYC2QCRjp
UVUcVeUCV7fRL2hXDsNy6IQNQAlCelKCohacF8eQPZTkll5BHi4TU9xkeCWCEwXy
dWIV64eO3Hu5bbal6+YpJGOMV89YUNlUdOFxr7DSvvp6vg2F+Q0c4cDyXTbJRStU
sqikHCMa1TA+/dKayBKXZ2fgSiybwbUGTOoonleS74wLFCvKQvnQMF049aFFcWc4
bduRSzW1qY9LlkExTo4Bsi5BimI5l0TXzUug8MpNzyhIHqK/VPsGtuYrzn80gxbT
LP/YEEv9rsQI36LPEvMTRyTdDtbJ+Nn5pD2CJf7Cy6TXYylkx+SZLacE3OtRJ4yi
l5tymibqZiaEcdOE3jYEcL72OE6ft72egyHunRxxfiL9LqT9shzm7+GKVa8b4jQ0
2OKAKgmNm/6aE2LxAD2c+W8DDugcJt8x9rvfkROPYjOlj0KBmB5EvUZe/TMBXCha
7LlBfRufLVtEIfwrNhxLIy5Ra0QSjS8J73UelWyHK686Z4Sqx3XmORcbtM5l0kLt
Vw0T9Y+n+qyAgni4cHR94KVnTedRJj8k57sUYavF9yotgeI84KX916jDsyVJ+821
0QtHct6l57NCrCnCtoVU9ejisVlVzq8pSCHcyRZewpInaVN4V0ukOKCjV5ojOS+f
2SZR9blGljn04KLq4E0zoCnRKgC4bVbdfoimWJro0nifJx0muTEahd6sMk+R/2aH
mzjWzYv3W4WhbMc0EQhYR8zMNmQKOByqcE4aKndBKOFzueBsMRKrxyO0fRaARz+g
oEnxVbgC9U/c6M8zo7xjmb+kJ8bjoAxA8pvvADalGRacxm/LdrV6tG/VtY4yNInA
ID6wHf7U4jBUyXn2/QZzCd48WXgcODx3ErTRZ+4g/r6w6WgkzYdlzpKiRILBG30/
sYF+67JiHvd4yJCsHmP0q8yo6Yp99SGJmwLsX6Ax0GeAu7ehVnrRMxo6Y2XSBR63
GRGzBq0ddffTG7BODKl5GIJ484SoDae/HyO/H4nXmpd+XcDzFWRgtWNmgNWkhsJj
mjknIrTqgVUHJK3U/Dralw1prFf5iMj0JR/6IM5wvf/mEI6tnoen9d8AwcUNANDe
QWUv9QSYLwpIU6xaU2pKh0IGJ6ncT/5m8D3qrSw42+iuLU34ubr8XCBIEnSRQ9a3
FXmjoHK0Ig/U8J3I0U7fUylX3En2G1dkP2J8ZtF9BnDJ8AdRV92aVsqY8oDCoxuQ
HTIXzGO+WBQksGKEbFZ5CenJOeX8Jix6xnqa+YG2z73T4c2/HNOk7nRSm0fy7bAa
oIlEeoxYj0Skf9Lh8M4gV9nnhZwcAg2OnUzkBqL065Rhdkj/dkY/b5BXdD07rGEH
BLfyUkvbWmmPXo+P2DqU3DgRR8d7JzBJ+rza3MeePYln/K5VJrQXfzWlR8IIRTu7
JZSWVo21czJcKBy+iyr2HI2USqoTsoREupwHXVxVXBk5W+6qpsZ5PTDZ/pqVPhaD
7/bzlZr9KTwqaMW87g76wbdIiKQBNuhuIY9cGgKuDtqj+vOmXoMZAomyFIC8Rnjx
7ScJgJhkILAMs1tNxYqf2JIQRMF8q5ch11swQVfKTYV8o/7hYjDWwv1Is8A8mdrA
0eLOwrz51J3K84vx489uxT++LaZCy1PU4NN59fgfOgtawmCpg3FVwOigCOwVLkhc
FB5Wb8z6gZuuh8wZL4Y+FrD0L92Yv/MxABDwcUsI4Aii8wy0lMZCzzTOya3MjF4B
QwZz2Tl/q/9qa57Kh5l1IgrwBP4P19bXm7pZEORLSSlxuJvo/F5Q/grHVW8TAbiD
kMv3t9cj5W41F3kGy3C62ZcmHPjh0tjLUvUNLNYyil+YuF6cvYZJO4KauNfr8bsc
bT7nHN9bzTYrLGmy09qGgp1TYs079izbB/FGRSrBHJu6hRrAcQTsxztBuz4CQjkD
uqafcx+qg32QCtcO/IuzcQw63Sg7CvYIkaFdEMq7aLr6vK45PiYwC/QWwezWKCfi
kZXwUrDtgFED6TnjiSqP8goPa5BTRyZZ6o6uDWPF7mWlmC/+lVua+ld4P78yQLhB
c09/BPEow+OzsAWCZSAi2Q+1TwaQjbAAEEvd5yjg02ay5cuiB3JQmL2EiVT5HBsh
3mDJBJmoWJhhYfAA9wqkSFyBv3MasNTWp+LC6ufgUncocfUTwQle4zv8k+rruAm8
oZZu+WKMWyRhIOParOABjx5z8kJSbAnIr7DhO3Bb07yIHaiBuOg0fLbYsQ0eiYh7
Un4xq3mBw5EZsInt+//YArD+3GgjowoX8owOXBvSNtp0ECGEf/N8geA2Nf8xryG6
EGFdPz5hrgNCj7DbIGRju5JvWqu83go4o+OJzMze4s0NgLu3Vzi1UHdtRw9ABNXc
FcQjDstZzBadrYSDdwY/Hqn/JzUasO8f2x/b7XshMXhb/XfxBg6GGw8EQFRj1X+l
Zn3Es0uCT9XTBamedGMuvCGAXE3p+vq+F+TiBV0JsJNLy96fJgYGCT6vKStJBFIc
CfeL+e/7D4LgsSHWkLrtn1Y2hYooGNSfJQOuUoiBpdYb+Dicl3rTACp4aBvcWoRw
BoKVESJ2EpEVM9LuiSKcnTXm7NjQuEjQ/y7l1Au/PdlZ43axaWfkk9HzBySFmhSU
zQP+JvDfvLHoSj71dt9CZ8XtjYnFar9GafPnWUxzqvUqMjZbmDxsEj2GT5hPuINC
y8IaKj/6txnHX+pX/ty0xkIDhfy5ElyQXqBu1OHl75EefLB/kQAX2r8qM5zqFlbM
L4WGPZ44hD8LjbcIBWSI8mGzFRyHms8piGIJyyh5SG948hiOx4VyPD4hxoXRz6t5
Vvwvsr9SRn+TaElGzANKwJDYUuboRuCwrd9qT0RmBwXhIo/CywmE0W0LhW7sGYxU
wsUPmc8Lmusktge+U/C7ZjERZyQBNH67oU1MgL2MLUNjks8nccPr4x129YNE3JLm
96RJWCu/hbWpNChUPJjfANPQN1epXBw6WX020potSEvA+VwEYYOauDzIaIL/RTd/
WMwPTgJYHFdqS/DmSQk+tdiwb/Mfxspfw0Gt2rneExQoHztu1FzDoFKeSgtUdBRd
7/4DQduCLvHJsgIL9TSHllfnR9eJGIy4zmnh+IVXsdsX2pasH2LH5TyAvEd0k4ib
fDon02UE9YoCdEJTAGokCXJve0H2YZHJdVmc9y2aTn2eMRtR6QXN5fza0aUPC+X4
ayTjP3uPQ+1KOTg1Ua4yUftoYOiJwgkjo/MhgjNHZYQEoJ5xDhdyP7IuRqBRfvy0
VoWtNFF3Ff/n5/S9QFk4w96DSspNHHmo1o9TbbBayl4WYOzmZyYsStT/rrDgBO2c
Gus+JXVkih+J430IWnqSUdKad6DyihpPX7tM/KpPnQOjvpHSdpyFUqRv2T9SwAg0
+gFHb2PcP1AYH6/4zUNYu04kGwkvAvLbuL6sCTmbT9IU4lw+akVJXC91uus1W5C6
6ljuLI6MwfikCsT7qMJO4y7IhZWZbUvQFTY8hMtpebcWs5HM7wdnZEBBc0IFlCe2
/PVeesjFKSuZzObxnuGqFNREIxNp2hXLYLOwrHmvWMl0aalKaVP7RDAJHlN8+YSD
bD+A/qp6WxwjUC37yZfcmqgtIwW3y5z2QXqRdMAdd+kfdboWP3Q968w4wIrWXz0K
fpGPiQcNHxjhsSZq0xkq+6wxvq51+625c7mk0x68g+BMrsjMb08XWA/kuwq9MujB
hyutj1EpQMDmOapsvBFPAmiIi1CpCRc3Rr2i12PwR86x9lNbxC6e1EnLjz4T7YtY
c+vuTOpDKo7eWyxC0+c2MHkVAZ2pyApR5dtH1BghmoW1VLxOXa/xPPwyE3UZSrNY
4dMpjimvnnigJeN8pyjIcjoPDAjhQEmlPAfSpYMs5KbP2azlLRP4S9OKGKc5+roQ
iUdZ0tF5yw8QhsxEvie9NMWTLsoNi7iVQMSN3ZB8RDq6aHX5QcVRlUKQ0Q9srGUS
fxlrFQN1gAbDcKXN1IGoSNfmhsDX5MdYGwGm3auRAOmMrPVk573oZZc+t13ZxrOF
6p5MBrO7/IN5poFF/UkocHC4LAMf6/FGNPlyrsb1cvc9sENyWrtCouWb5U+VtiHb
rPpyYn3e72frHEhmY/gdsqVZmdC2LVhM0yM/YX0cOUdFQc/JEnUzOgv4xUVS4X4J
h0AIFwveudxD/Yw+Qp/5AWoMWlxnAG8GQcCNsNvnQpM0P/dGNNgCnGiQan/RngI8
`protect end_protected