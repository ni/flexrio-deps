`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7824 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nn7oC/bbltaB6y9f4wbJdgh
0G6WvBg4Flfb54G2gjKn2w+WOPqGZIcqQrEZ0Nt1IjWrL6c40gXCAEE4GXn65IVH
j6ZclpNHh/Gxz6ON+l1qLQiv0BRjN1lCSZPcW6N7z8tkOqHb2KXIp6HwbFyEkMhi
DyUQxVF9Q9akJiW0uYAN5/++AD8MHiMcpwY0k/IBEcSMpKfZN3lZNIRx2vsWl2Fl
FrImrA6CExwrp2OwFACL3P/Wrxxb6veWWFmLnLzarPYl7hlsq/hoD66xPoQsAaP7
jC5buuOwDs+uuzWV5c5EdNrD10t1jLwjBxItowBfYIxET+y1Gw/c4EwIXGQ3pUMz
bTPkb/to1EmHvLRbNutGIJHx0mZcAR3R2Vb76dvpV46lYQqAzT/Ikkwv7oLMm7P+
KYCoh9GH2LCAv4aSmKPuChXLgLIhSPm1uZ6Jd8em3zsmxYRcHKg4kIrDwPSZIg0R
ikxUlvlLt+dwMK03iWLZ/+J2wxSv97FL3ZRm9i7ISyfLG8gula+UGNmY4XJkjicZ
WXyhjmqxUMGdjqFPGqJl0xe2VHvY6517ApmvQzUnVLJ15WwmXdMJhnr4Rt8f3NPc
tlUPwfnDoc6f2PT/6lXuCrYprVxmTQpzh7XsTkjdGjOIOaaGYwUUpiTiXBQejTVY
4Hqk9qufhgY+ueEjd4SQ6zBsxyX860/6Y0BK4RVS5zobVudu8akU6ObJ5kERDWPL
uVbOd7zZplKPyMUuEZaIa9N90NHIz2/NWIi81fVKXDGXhoiGdkpKR2fmDGYOs7OD
UavHxuDAyucim5Wi/7NchBKZSOpIXfkMFBDpUe5flqvo5qBz0YJi136M4r+yyEpz
6BlKuYh46snyR3MiygDOOnlmzJol6AFIjJzEviSBqiJWhDp0NaelEDUxAkSItujf
SMLmNeDDahsfbEL88XQ8u45Cjmvv6Tmj3gRxhBApBSltRuGkNBVP4/BntGcaE3kW
H4zascGjd4AsPzYCSEpoFHaJz/zhh/6RusHLjHzBcJOkJgRodJsaJb79b4RWh+WN
BJ6GXwcFdOIp3SiUbCb+3IDgs/xfH1qT4ugKzgRNFTYp04fZcXEkhIuoiWLpfhO1
LgKX+IzJJKvLSha33FUaF2h/JOXpbzsVo5dEr1yv1jVlg1sjLqR08SS1r6Z9r1ML
y91AAkRHgJiny+/GGaB3UUqkNkDZt/a5+y1tSUfwXqWIJjMNcjDiXayFRvWE3ElD
aUpkO78mgQ9sovznDMAzljBUAduYbJgYz3FdXJMxkufmdiBUDxcRqOuZJT5gaJOR
xX1OF5wWRvNfdrODQeO/Yr8Agic7lo1N/MWiFXZruXxGM2f5FPObaME2T1xD29cP
wyUBOYUc1++r6fdXXQ0fzPOcVBFIp/0bpk2niRf8/1AlqFRVnHxkPiusvZiE9oAi
Va9CPn9seoxuNEso98bfVX/05LULidCfe8bADdNMS7rTu/9GvhGV++uaUbjtVF2Z
fsGUWhw5sir/Y4pl5ZNZpoor/EUQ7gl+afwpULHUFyRzF6Mm2Y6W8PZ4MH40iJrS
CEZwfzt30eadAHchoj6zV7CJhLQfjjLak6UEPeAokgP81qHDA/nEq29SxXobZTFO
Ulqox/7Sn6HFLSNZTlp7RUWP7hq5LqFLfdrIePDGTQFQvX6kEARnbbJXeW9OOGWt
KDf4/mlKKwwMAeyLZJ215cKJU/VErRpRZ/1GVhls4NZW4VQ8nPkolIXjK2a3dGAJ
JvKKXU+EbD4NOnT+o/XaY+zZMmixPhAkuScPJ+BkUTcUEpQMFElxg1mtIuzF4bSp
V8NO+R6OeC6W/yeZu3Y2iezRHuMtFAhQtwS5WTuu1aiWeB24iOohXOdrFXRqZGzd
NfCFaAizc1E1IXd2+CbwE6yjGlNLdH1I0n/A4uDeTx1j4GFtc3DEg3E9JZLln0Te
SckvPm0GpsmyVUvd0FiVqdzgN/gSOim5qvnoiCIs5JfKZagbKh+qc83E/Tvj44m2
kvVARcyUmqFERj5wplqgDYH0V2oZ9n1rOzYNsmQ9S7ChjTM18mfD7BV+mLmYUkXx
NNFPIjDE8t3U37RADg5AvlYf6f06tZ8utPIsoweRjhspXX3KkS9UmnarlkcsmlZB
+mPY6souHlAIkT/1oMvdpYO1xZLzb276dd47qAsgpt6rlCqxFd9m7vuN4M9U0hZE
ukEsHaB/L2roH/tF5jX0ljY6NmChZ8IHo/7dcfDAxBjvQbAIIfr0hXt1FKPcgn5/
vzvx9XTQ+ozq7rLPgGSDgE51L9Z8FZLwSdTd1iBqc7x4zWoMNCn0U7NJC3VdAitU
xZ8mrcx+RKWIR7CFMmnq6lM5FI6GAadgEfTRgDXM9WRjBeC1W2KqNQfRH++y4RO5
NRHS8rjFYWepQk4V3A5B/sloUzKQ2bs4V23eaBKySQvtIgZzHfwl3tziztgIWuzb
2uyaU1KAasfl6tRVQw6WewNsGiycDOpSbceHvsF5p/F0Ighcsz6EtZ6kcFWl0Eoo
Hyv4SuwV5CbWYYDYrgnWccACCuJzx07KxYVOFFCrk6vGUfuEElyOfbu/DqfCmgXM
3Nn7GKCGaDk/RF5NddR8yyGplwGTN5ULSWcWccA+gJ7liT8DmZt5EGPE65SBlngT
jEi3R409w898I+jvLcpX/7xUaH7modPPSrarjqtbD42ZHk0XSXTJYP4mI/WCKaeP
VNlhOb9zIicXkjFXruKsI2HvS3+hlbodr5g6O1Lck5fRbUSZ/OpIkrYz6J4dmafK
BIeyCTKE+D4bIStacaivDtPebpwUFysEjsVm7hnoSsP0SUIosXwywxpfqIoNz/J7
bQjZEh2QLuWD/lMdj4L/JVU2/0iIVL9LfBUXl4Koi75KeNQbbH3dxckVtfMwmI6x
qw0zWcqCmhWVLqL+zv1C1Jhk+I3MAKoLne4w3V7vA/T+fyFTWwTy5E1XNbJ9tjs5
z9iIQ0RUWsmd+XtbCarESfVeGf3acGs8ftKQxL5JZgg+k/fq37plG8m2Ur0DdFlQ
uvQ7z1UfkIitnVC8eLxtVVqCswsE2mHdn1+o3iTDYq4hQgz7FX0THgtt2QgZSFl3
T8ZGgp4JDDpokae4vEPIPkSg+ermMsua2ojHRg/EZpGpD7aWREVrOlvE8nqge2AJ
0fkvFgZKED+dJ1bkNpqd+2ts+HGLRPVLvR295O17dpyeTYXZyPlLrdSVDBmGcb22
Lr3B4d5bnfZWgZm4wesnrGOVqlJDJHy7wRSVF5shT1ElltTfZES+fQEZp0Jg8/Dy
+DLmuAGtvHsCLA5NbVRqzwTOVCqcZGxYaPC7EUmMNCtBUBk+m8vnggxU+4cxalJc
lBGabNKvYppkHCJRYKjWGQJCkrVXRKHdeLrN+vYMoFs18usZdQonpUdJTUBaRArw
7dNg5e2yD2GlS5OIK7BIMOEzjMYF+W84oxT0OA8aWP5i/MT/ljZJ2LgNRoIYUM+L
0e7NPAdftGQZIzgJAKHva+ISmoLmvzGz9KlIb/El7/YKI2rLuWp6S8OGHj1Uzn+B
jM5ntX9BMEuGNc+sDUXcVGVm5tYGyDML+0xswj88+nWONjoxktkAEYtFKw5DSMMC
anURy6tJYcC1X5kh2Bnhl4LkVNLOx9v5XllZRHPVX5FSBN+PDOzYc6KYAhAASAYa
RxUZ+G8KosTN1gr+blU/spK3EV/mT2TXnmgxgxq4f1VpP67VLbHvNUlmi6q9jb0H
S8cZgI8FGvw3XFioissmeTQKrBNkwLnPXJF6byV8VYnbkOTA31yJuOr1cNFuU2hH
VBMZz8GaRCNWY4bD3E7AUoyDTb/YwDzdUOzJo3G0HWH1/Au7z8GnWNlV2yqxgONt
+A9azHhAcBZ+R4CMOvJPYPof4gaibf7b1uPspBw/ZTQjw+fatyJ/iahbXQp4OXvR
xD+H0abwFbjfVIDFTwl1nvpG9em+L9hkWBhbGtITcwwJ235FUJEhFE+LPjvTDHps
ViyfqjWon22Iz6gaP/i4Jwl6WunwE6T0lbRIQxWPKON0BMFqcHsrVfKi1LHB8lcI
LMy5wi9DTkDuqQs4lSl59HFPibM3/DR3E4L5iWqXOam+Gzpqk37qNuaBmi1ce6DZ
Pck54Px6YxsQvQw+i0c7Z5lJh/1VsY12npRK260abQOQq+bjNkISCjx0HedPHqDn
DGlWm2uqwaGj/3J8ZB2W1vQwJ8XmNzt/baJvIDbHmpz3/aOjLdc0ohuXpqjuOVBJ
bLkQgmt8egqPP6riFUsf2SVvQm5BlUTJ7IDaV7xaJMbaqJNS7uWnnlnJeUjkv3tL
RgnPUHsuwhUxzXfW1ibTsKHxLwh5MDqGPYWfFyPYEcvHQnkSxq6HQHeXYpbfaj/U
xVR61d6HQ5DHCtCjl5Z6bUYrXKpaHn7UsLWZi3bWSt5rhbdK/rbA9m1wXkBT/Z1x
S3v+OBDrhXBvgw+EYLTYoE2GcO9vqad9CSNzlLPBaz18te/N23M0xsXY5IgGEuIS
HZ68HuMn6ShkbAxs25BvxHJmFarJJIu4LZaqzAh7BIyURWGtatLzOfA73kdB9sHi
MCUEXpNBKu4BC/8EpCrdub3tD6/ybyJFaDa5ZQfhBJdmT0FpqPmFN7Qs/K5t42cV
DEZsFrNSHhLVhwCmqWT5SeqXbAGU1CGkpkVHNvlfqwi9RuHDdL97+dXmQfzWJLoi
5DcrGyvkoPaQwUBl679hCV8GeFufySihz5I2aGTP1cwbiYhiaV/7nHwlxx72sOJz
BC/wwb+/U6kj8Vin7sdlD1lsnDO3q3hy+xc+UHNZ0ou6Jc35PObEP1/FljmVYvDl
h5oAqOoQ0f3C4WgsjJYA+ygMzKf/lU7Y8A+l1MM8bpuR8tFMFC+Vs8e9RUJGyTYc
HBxxcOxMDphe2mlAAXnezPv/TaoA1B3fj9shfVXvYDcwJoeJicke2IC07whydeXN
pvJS0LIu//wQc04vJIFCOqbNr13iMT7OC7Iu+lgl7HMmeWbRVlXo0cYPbELT/DEi
x4p/PvKYNCw9id2p1zydHOc7TfIj9JOrvMw8U9Z5ZuTlu1UvdlKA8GCLcnJz1cPM
VxOiqPMxlS/EL8zuewubCLwMkE81PSLGJ2EQH1vIV5hNXila8H7f25ofvACyReBH
k+hkdfPfZ6ZM8mAZFmafN7Su6e/FemLKJPFTwtUBiyS3rxi/yoJdt+iCU8HP/pBW
wEyE1ERtX/lBfgzib7J2bxxq0D1N0wnRgENgMbgmvW1y32BHblHVENNoa4AxsQaI
K33EtziS+HfOPcK9vcAI9awPFJnbXevvD/JENqXfFp9YPjSYUdvlqFuDEop8yd7S
wLXahiUn2aAb8GRtzuq3oh3Kn6Cf3Ged2TBadZ9/Zlf0ql7FuHTfOC+IHYtXyHSR
MI8RrwnoCSSHF1qtarydoGE03I8zQcVgMQwgDufa2LauArczOYQ77uYvF02XvDFi
Mi9CpfFYM5fCi/1HrrZwK+WgUUQ8+mL5A+8qOogMClhdajkh1+CRLnxB482KF+HQ
xaD2kzAwRQSEfwH/z6/hESzlbGr2PrD0zVMDNEjXRm4m/jw1JfOXeo4ygSwNPJiK
320yfuSVAUz1SQO2dQG37SAmH1pb0L3pfluHFvekzLo9h5Y7i186Cmc/xmEAZUCk
h+etOs83CKmBqbAB/c4P1O1c22UpX+l7oTr2y6tOlbX6KRBzm4STqgwHl7ME4BGo
g3ksLHtyPAZAR+bGmxped1295sPPguGSzcFWYYaidsKlUxsJvKeTKpdYQqCIwaHH
HgxXWY2c6LChAiPKZclNg0sS2gLFWK1KIAjVqUlZ3q8VS1pilVT3L3xHO77sxhMz
kRe6pThqtBhnoojkmbe9HzIUJzrZ0j4z3iLxkA2CzojrzpmZUZ/3Sa31SXMnS9zo
BNe2Cg+DV7aCtX3+s0QVqlsybsHrLeAGyxDIJ8uM05flN5/Vb/RlaIxuIK/Z3QvO
c+ijTg4OkdNowufsOyd9zsmEmYW8TlMGvnp+0QYwOMh4x7hEk+MHaMpFpWoQ932w
bwXoNc4+hmNjwKQo/JZt+ZrzqwvkkEU0hYbFuftR9+wEzwhGFBl4lslKSKo/CbhB
WqDUDXbLj2Qxwpn3AvyA9QjyWuojfEUA8fzHew4+U/Ty7m9EejKZrJBE5YU/ZhtN
DuwVH1rTM0k0eabNZ6gNvYAl1oDCwtsfqaQakly2SustT61JPc+lmvocBFjE9smE
1orCQ7qyn9u2F949nl1QlL6Nq+TnhRXRTeCbfbf7ZBT2ms/zIvT+0vrkeztKauyS
CP7KgWeuk0V9szZIkg3cFUaqOSvnqogIJdv7CcDRekR5piqfPcXmllagB6CK7l1D
Z5BAq3dwD2sCjzgN1EUA2iYCQUwcv1iY8l8Y2ujzpP9FzDCX1zZ5RGPSZCHUjDlx
wuq8m3bZwjU3VLq/FnFBjghs2+evR+vuR6wRy+1le04sjmZHCP3D8uanw0mHSGbp
5DT+V85m/z2ZVVyC3RU2T1dDUgcJFf+FMfbJXfzrw6QKTgdyj+C+dtWaki7DTjHW
VT5q/zErOvmnptUCw+Q7iaz7O2l8xN54uKX2oQamV3TNPO6OX061XcOjpePN09Rg
X8EaAavtQB62gYu+rhVbrSEoVFjcEFg60dPvNGCP2VqZzri0/dCeE8FAheH4FAKB
QmhD1wWMkl0+jweyoQE4jkipGTjZHiZYv+f+jIk8e1Xv2Kqx+sq3YKegbWT2VQfV
BXmz2u0hR2gQaxCVShJae8LvV/75SoCxnxmpqdDuZIW/Wz9DYe9Rbxl124myoW30
jBKNyIFwcez2LmfgLnlyfc17d5tz1f+dwBGHfpCFiKrW1QjfLXR78Xb9fy7LZSG6
DFYNVxQmrKCnwD84A9dDNpHhQ8SwX7zPHmBQcTSOE0NIgDHTLYvorXeEGrQnj6Fi
u/7QdH19GkD40dgslVKUOwih/iGYsYP8NCWuBPEl0Jda31V+HkRi5Am/aoqChMn4
DyIPjIFH0RxR7nO6T5AooulVrcOxVg9cTxXchTrd1qDiQ9jupE1gm0NBbs007wrP
J8bTBlhrQwRlbXg4VH6HkHVoVIWHaL5bfkShVzHdJqVH37pEcKiYfJnQI8Vxafoy
aw7c1ojZ72VjlSX4hjNPRYlGwgfqfAA6P8Taz+QVofFyxSRytu/injxEym+0EveJ
wPAF2d4wJqwmYzFWyPWdX3jZxkFe24PoRmhhMlvMLXdg/sUyAOpj06nNPTcE+8aV
GEY0aFEdVNJIhhwn6mdenDp6/r9wFo5m4fLq/E2EnvXOpZFzkAJ/MzFVuZ2H70Pd
O6idhIiC/jPEgeNaE24doT/cvExZNpuXG16ubyvrrVwuTtZvLAvjFQlt8qKYsANa
TJVNUhHIdrvx/pYZ1vRXU/tvg9svdnaDKoiT7ZitCQrZm/RlskKYhBd0wlPEIeP4
ZiLdkTuWxmKHWAubsum7fAgkV0MhKBtc6TOt0w9Q9Ms1s94J2hQIA/wgmGez7/0N
ERQtytZYyhI/85PmSxNq3Heq2hFJPF1zJACJcgeqyaAtm64srpsMQj3bydenbwdY
ibNINYv0Fk8sa8PBnjiMD/uzMv5ZYsBFiB23OsHP9Qd7jjIDRrasVnvd/fy82jjc
iU8dvfclMgGB2jGvodQ2Pdvcg9JUH6+VaFxgH+6WzKmQOtXpqyIpUdHVmZXgrPLW
GKFT+K5pGkVtP/jKIhedsmVVPmUJLaoS0jmkdNJygUPTzDFFdHwh4OTjP+WBWVRt
KW7eWRCBDoF2AWBzhsYd+iaLl7fLlVT036j6qEOLjeiNzMzzXEf5oF9g4td9mz8W
xfUjiDgFsptXihw9bFxraubODIW8Qx022vNTht0hR5fi/m6ey+4Ri1J0GaQztdYp
j0XtLwibfTtdKr0rYCDW4rUGKUOiKPwxPPjtQLxEH0G10e7CZqTAnem1Upr5kGqp
+u3z1To/6nqiaPW3skedji+RMYPcguSsM/XxS+azn1+rI0aY6BJM8K5j8S5AkD/c
Zpdl5cMmBGbtIcxzH2RB69lAP8teOnjW3J8PCmf8q7yMrvcUIuD7yVggrdUU3MR4
rbS21PoAfzQAjVviFqD/DZPXwPD7vDpeg9hlwNY7rxDbUvqMvrtTmdcReD5HU1dQ
mCplfYpwFoCRDim0u471ZEC7o51BwCuFrC3kS15H1Y1mlEC47OmYnrZ0o0vyPvKp
/i5Pjvo74wLuJIfE94Lg/+CMGU28mltZXiDk3ZMo1i9GSeXcRHrPzKJGJn3Go3zV
bVsPJ/uSYaTBTgy1Hc1xu99GXr1HYj9w7iXVDiP25G8HP1YFrCvKVupwGK9/dsNs
FtMACkX4aGey3JN/tHox3Br1v586EbJ4aoNKz1+XOcgP2dJiv9wI1YbpiBZAwvkx
g0VyGe133LiSQ2xRTEh/HaoIZVeCJZPTRYKu8Tz6kZpXTHMgUK0Lg0XaQ0fyXhoy
EBEVfgN9ypt3E5N7NmHmTiip8TSxX2RlUTHR8xSmYiRfklya44+yI2v3D2zks5bq
toEVo2Cee4ZBJCAhXpngvzxsINAMFhT0dElz0i6RgQB6gtZtJ60CPoNocIaCsfAq
Ink7ga9Hi1UCq6f3gbsGIY95GMpZe2M+Oeg+N3wCyEKG34G3XBi2TCdV2w2RBMgu
LaaPK9kr5SsSgUVkMs/oKWWe2TdEPBrBHWVzSsL+nEfyON8INSOdB5Jp1EHWUqWj
014S4Hkf74qfUjTTtzNCzPsmspmeX2eJn7Qz638AkGf2d2tO1xD3pKjRUw699sGc
kMGnxcqyn0+yPI7jsksfwM5aCei4hSCOv9nV5wx7+wjhEkXMdZSDB6n4Nk6wB+1E
MncDRUtpcQy5/nDix/N41glluWTsOJ55hDxMgY/PIpdLQn9v7qQLATcP2Hm1rQF2
g18RK4hlJRs4z3kfbKjEfliXN96MbyrkuYbU6n5EQIzBm1652lsThdeO5xBt/pbU
yQIfdxg/4Tr4WqeWrblckaDtjdooBbftCcsut8CgA+iqwrr31PvkoS0GOuoTG1i9
tUZ4m0SfwYjyhyFx481qEXLwxszxEKEh6LciJOw/tlGSrr/ZT6RWO0kSjwGZmLjc
5KkZbVFDfEBVuzOzRT/TL+FsF8OHNc3CV8nHEkQZWRyiJBHBzopIiu365fO9xjiX
N01CUudkqxqnj/5rQfOpN4sDhJ4eq1o/aBNnGZ/nNAzto3S5xuSlcaa7k+TlGFNZ
yBOD1daTpZcUvKDeFF/aAOaCLBZkopHst918X3ui8lzHOLA2Gb+wy0xrVt5N4c6d
HiUS8aPTTYPbUWOf3vPo9YjX/UnuAIZrXFzjOIdHnlIdss5U1z/z9LGa84+Dohm2
DwSHUYZk6KjyWysVe5Y0fgI/6dYH5Cdn1t51kmbKRwIXx2H8p8cIG2lyzoBcK2fM
/n57Op3n3XI0ScM5b1/+9sLeYQ7pisgAQC6ruqwl9OSKzv/lR/NuuW3zj3LCP+mQ
C81p9f1/cfPeGUxrqWtm+MlLud952KxQ/O2DwRDKgQX1c+9H7Iv8j8PcHTgMctat
N5Jppi5q7Gliy9fvvd3xnjQTtjJH+yvZVV58/5b23VKaFpWNR+FCXnteyMY0boFK
cgwjSkhw5o/EmCr96QafENNgtBkkSKCl7dbsMng++a7Xbls/zBCtcJ+MAvdP3xO1
ZUqtH/skpmSLX+BJFl0YYYPWkmQ9QMnEnLUII2WcggPOgchKyeXz+fq0zWG/Acsn
JAttSQqq6zOsfpHThHap0xDLfamA+u0fp7kbl4HyohqE199A7BE4EJYjfSfye964
fz0CyWWhBMR9VebYVeVJW74XEj2s8ehAsO8veJsvOKPaY5DANaak61bfrvRXfVlh
9Hvj89pbY0S/sGEFqwXVhLQ3OGqOeSezimXIiwCo9JmfCp9CT57skGLtY+oRKqhn
sITiH8Mwyb5fuJcN0xhEQJOc0OPJs8JhIjCmJQVxT+RYXaiXN4+jJkCrgrDucyUG
M7YWusrcV4xnv6p3cGkYi7jG5x+nyJKiw+H5Q5ODsCBlNzlBLa9txTdU8zTJlzgo
lfStPGBExxJabfT5xF4px+a4rWF0m819LkJihFgnY8r7AidnR2xPsZzLe1BcwpTE
moOmTGOLQuiu4O0M5B34zUHxQxQGdzaUNUESaVxSAKDZ6GTJVkA4o6REU2UhFS47
kbsYKogbPH5vc1alPW1BVwMgkJK6O+RH3825gLrdX15C8XHX2ozPn/Z07O+DZBHI
YaFMRgsknPO/zU1FecBAUue7f798gFmaqVB1F097K5Q4x05XCs6d89Q5i1cw+DV2
`protect end_protected