`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2128 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
/8dei0SfYi/yIzInIePi3Iv0soVS/1UkNKf+yxf9BG3AVnkI9oxFYvIJoqb+5MpT
kIu0QLOX6pS2lqL9ECJuAyowYCWtlVg4iEn+zujVPyiMcnp4NhX4tu460ZGe3oyj
eJNcUnnreYaFNzXoeGyjhR+gfycPlFPZ6JFHVuDwHqzrGHjGYeXgRyHJRLu7ABrH
UxyLTHogeBR0lYjQ2DqY+Z97w4kRef491tiF+Tht9pZLV9ajhFC/aUL613GpMntY
JtYmQkaf5ygEutDXlGNLzrCL3GNCdM6PDr6NOThCz6FDPhYFSShHDgV4nzxPmBJU
hfxwHsRMVxnnzbeZdzfDgbFc6vHgjZfh+uvkOmmudcN6D6Mg8rT5FXtqfFvQq5GK
WJSmLYwo+pZfBeJvuxWlfp00B9uvwtvaV/T/GakyDv3E4vG+si5A6pJakj2z0afr
ikdba4Qiq6kPbaHEyGHKJw3//KCHhVE1eDurED2llvishOxICjgkjhayPubfdcac
tW5MHNCz2X+8g196whvYWRSAFBcjFH8SdDLKVcycq7slb1Y/lRkhZomKmOjCkovk
XWCJJUZHSDGSKdkGOioZgR1wst8JzYpaCS0RNZpsgnt2LtQSsTsyzgTtXyff6XbO
yUJpZJVl6+3EdsFtPf1dgCVoXd/v5ECpSGx++78KO9zG7fBygsE5w9EUPVnq7iqf
LjkOU0xi4dnLZmBrr9D0/kX8/rV+rJuSlg8MiqPzVPr4MEPwuPLRm4ZLzqTvjOpw
MAEgcdl4HA6ALS22TfGH4OL9+i6B/rRe80laBPPYw76cyYJVxV1Eb88TTUgnrcbC
GUh6AxZnKNntRc+WUttN4Hx7cN9mWi1DBlVKkTwZufvbLac5rb9pg2ljDew7OaoG
P6780DvAy3Xz6c0Wv09tgJhzTXQBwHDZc9LxUa8BJ3gjevPfwgdjhnaUVvaGXLXV
wRGpBC4TPz+87kMSs75MKHKLSwR0GP4AqtbygdIuZPfNZB4oocbNnvkZClKP7IrO
EEaeFgTkMXpSoNx0pv3rzmpkT2aKwpd7idhGRygIyGYGmVUX+H+2bH8PbrW4usJX
KkdHOKUvGrFZIX3uNhYNXZppsYjBzWIFpvYL1seKplACBOeKFhe2dw4ktKTv08z6
BtzKGhozJ1ErojBBM+a1a1ivIjs8ohO9MVHajiK360atRp7CCTRSSDAqdrB5qTrU
Hn4SqIp9iwmaqOMcpuI1XCOVlXe7f5LrfHVGppR5GueDFB8qoOQWyPuqcTrwPHgY
xFsIGZYl5L/wdSp7xzG112IEOeoXPWvmuiNriuhjgcAkQtzCYYvS36vvu9y8FlJV
J3KPY0yI6mH8rN3oz/l1SmRE3F23AH8o1eOVcrhhshNx5t/TtMrGEIgRBsEAabEU
qlesqTEuew8FTrGE+/4Wl1K/JEMz7s1jmy3OcN4sjXe5iG/k3nvjqFYdi06AXdEJ
HyZzw+ZdydkTVZVarePOK1Cuv6LqkdzB+ss13hp61y7WCC0lZzP/5SozYNKhJrgP
NsBUFB3hnmotz1tled+ug2NlrmX7J3OcKii9muZnfi/FFoe75Ew3KNvNltfYO+yo
RMuhOgk0Rjew7HRYL/eKKLPcxCtaFU/CIAIum3Iol+NlYTjwRJPZ8idZshFTXELn
8322zDuyqWXEsv8mTKbVhal3yIbzZA5oQHes8nzL2S5pf+9/BpUPE2a8ARQxcofo
IORElxk1P3AEGVz+YfXw4jNzsj2FmuGwdB8hltR0vbz7vfBeIRDJVUazgM49lA4d
ZU9/c1G2QiLR6jc5/vsDazlG1p2JGkCUMs1yUG+VaNhTnRUF2FkJctIvdcsbjWCY
eMEWBDww6ZAGOYUIvz8Oy+i+ehkFopEvGNAw2t8KWuG3LSe872MrYHZte9w9xWpY
Qcz7ihzJ5EnUieCi1s3mif8fm1ZGDdeIwQyfzRrXuvXn8UB28R+tSPGHJ+OUdN1G
P112oJE7ARXLs7/Hhp1aB+ZpYTE3eu+q/ubwKjmvS2GCuUdPVD5Rzsum0eqfTHNp
OBGV7iJgErWo2OhC3nIrChVa1Jb6MVHeopmShLMvGol7e+2JR7v84s4YJsmeefmz
0Gct5mcDlJHaJGn0Mc6JhCM5vk0MmqwyZBGbOYI6H+ixBeIuTVfu3hlVcl8MrmdN
iz/514MEY2XFRBPTLQiW8V/P498ri2cPwF/dHy74MDjzFFocwv9DWqUSH02tsHuf
szBC7v/j/eFuVgnY1SzA/7UCGc2piwdPPOkeDWGSa37eWguKW683rnCes12MBwaE
LeSHtzx1CIOz17W9119Al5HYtQkCVTZuxsihpKMz5GtY+kQL8WjSISTMC2riK0qN
F++FOJ3ySbJYrZsyI8NPFasqgV7UtgVCdmuBOnnrsYm+34GeznJg8S42w96pmZIc
IabhP7JMOtso+0AzanPjvZl1gDnTVE45N10lwlyAGv30iDevmMU2dGSXAnUSjWc9
r6Tl9l9B5VrfYTlbhHFL9FkFU+Yd0MvWQzIxVB21QWi+dHS3JaI8KPdTqU3haIRD
u5UpeM2pu+AJcWhTFcvbEuRmf+vO/bGI2mYeJH0jmNJueDtVxAgiXhvn+5+PP0lq
YnC794oCjMi0AbebA8eL4qparqKAws1FZSPAXlIfJJjIW+tied+7CTor2d7vStKZ
y3pqa+MlDvlIndkdB6jE0w==
`protect end_protected