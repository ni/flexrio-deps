`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
Z6yALt3nnSw9nTnZfQBUNTnR+I06uKzP8QjuhVpw7Lk8htv6DlyZtthuVoT+4blR
hvkaRqiu3gXxOzvpEpgQYF7JKSxemOGiNhlRs14ZC64hkVyhPrJFWvIZAwcetgUA
q5z2mcEdRrbp8mG3QtZNsBzqaRLULitCzbyCAlFhSEq3cxM2MmVzwS8lrLPflo6q
9pnsz07JlcgaCRfyatzLlkqajWJzWREqbj2SO0EPReRcjP1QF7Im2HR7CtR4ZDx7
8i89RjBnqr8bCv2sFzWlaIzFAV1IUQg/a4SdZEmsvHsHfhbvgLKqzBcHwx0m/uEV
TzbrvO2eBLKodrlb/vddLgpfoA4PNZ3lELrjVy0vVqUeNizZHOc4PNEAoPTBYkQ4
FpfhK7zqPqSdk+lr16vAnC2hQaumnV47ojFF2S5FnT+ZPC493OXdCrqwynsLhv+o
+2AAcI8+bYi4sH3rujZF0R1TSKv+uUmfSNplAjeY4ABucWfaugdXK5lNtIbT5f53
nF2yiHyisvDnmpQ3uLlbgi18y4KwH5cLpc+QVlOlhssx+6qBp+LFWuBzlIvewOJf
UCTZ93XxfdfvzO1mJbFx7T0dbOJLL0QdZbjxdh5OqzXvqF1uGc52tLOkN2aDS/Uj
Z+e6XTSBKEv6B3jNncppk38R/v5ZxFRS8GO8AtPQc2KSYSbYYtVMcH1DQ2Mo8qJ1
nGg0cHvvPx1YmteV3o/jkdgELK1hHKNc2TluveJMb3W1qJCv/gyULukxVhVXFZWI
2Sx7MbeycKrSy0SdlWGBc/DEMAEle5K7LVyiYtprsfgheioI9DYL1jrWPVVvBexW
uimI9iVY5V26EkfNqIOSKKezbR0Oynj0WvbSJpxzTliTGSWSg2xnSsd2Xobvjxei
hlSuLWyAWXHMIHd+bZ2IQyk3SkOfLWmxAau1DeRsIUG+6Y3J9ajGY8ooGLK30vpb
Rj6l5VdxcYkbaxmUc4P+YbkHmksfUKxAm2iyADtT+Ow7BVPAsvtanZTT2HBOhSPg
sK8Kqcqih4jML2TcNC/PqfMw3ENer7eBvrMkyop3kg0dKTQdbG1fSEgfuAJVbdXI
870ArB5PYHJRkQJ4ncE9DEUCLfLMR5Q1gLkWgJjMpgg2a76lPI6vJ1Il/zgzXIU6
xtBfC2K2Cin/wR6ZT6ncd+oGdO26zXTK2CcC2IRv1ePggYGVnAsF2NY2/8LcIVnd
xh6JRP7zkGVNPTunwQ+y+uOVnzcGzhlhlVnWih+YLny5ZnAlO0CVhJm9DzMn/vvA
La6n1d2G/5UlANFBAcd5NpjZX56MtC/n1WgbBKbxrVDHZjJYs8XNphzenmuMgYp5
AyIs+9PJ1gSf4dO9k5k6axVNMAOxbbIVJUkviHnW79jmxIgKUizuUfSjZ7Sjjfzb
VGE3P7kBIIk+eJnrDDaK1/iwdcPcnTvl2jxKEUeUar6Vk9NRSNh0wHZBvl2HNK8n
4bl+AYLNS2R2fmdrANwKNcqqEqc6emsEO5hvj279JPl2DUXpp33qXJ1c0pWXAjdx
c/1vCuAcApBRG7udZieET5/10Zu0hA12VtXQka6r4S/j1i+qUvMcyV97wQ1GUVMe
JMZMen2zM0wbm+xguDNAxo6iRIOaRet/XmHooSYQI78i7QTS1HC+MscX2YqRxZGZ
Imq+SHdlD/2f/Ylgpy2U9gj7gXbH/BufbvSwnru/vW+qqnJm47ZgBplwGASXAtU3
2UWo8qig0t5AGXX2z7bt3shPSfXdYMstcYP+PvNU11osYU8W3BSQ2sdOldh1M5Ip
baXwBvF9sFVQmOxOwCH6WDBAFnaCxrrrwI9H1gYpDwIlU9Yk1eXJiX3o9eU8bsBn
eFVOvY3PSNpQSaG70XXwOEe8u0GpzhhhCt5oEsUtt/RMYu45en94+NbSA5YInQZR
GSSMsMbU/GeI1OuRBcBdndaDajmEG/UlOudrwlImblfBdmYckBUSuo3GkeLckgJX
50B4Tk/L7h5vcEpybD96m6DBaJW4UREwRV5R8pejcr9buxfJyNkkRhhLUZYfjO8b
QxHEGi3KDfzFsA9ZNaIVPdALkJk1UgE5EsEQWOzEMHHrVSC4FATw6dk7Hz4SZHa0
oDjZreYo50lnldd5t5qHbFCjDA7AeolHTvvUpikfJBpFCPiiOyqNchU2Rd9lhDBc
VtA+q0PbhKkUDnkAOKvGnQenM7HRBGX3Po/QS7K14M2kpiX4MGl/kcgWhRDynSmO
DTOqfmhG+awNnEqbFc8Gns4ELodJWxQQPZZlCoLXYcL5sKYQFkXJ17t1cVI9gcbU
vF1ANACVaSVcUqdQlemq6nQpGJGAYwQ9IYlMY+u5r8C+4NkNp6VbWCcLVhIglf7q
C0+yzASu9QRaPRI4811WidluLl5AuJnMKoz9K/e+j582LetOKlYv9UssA3jADtlf
8Ot4iRNErbH4yLaqN/tBuKpZ9LLUS0Q6QU+yMMofJ8Bz4yVxze1Lkkky1L6ip/KX
hMWMX1lrxjUbLl0suAo88Cs1xWYu4OhKPB+H2ELm3c9wajP1V5Tw627x6ICNBDyG
ZML8ZlFoFnsX6dg2cfLuLEf36wkxH+zgPQa35s8JEPl6vHOZcfpsPLSZO9YKg5hK
f9+NGCtIYsNe5SgoqGe74+P6oylPw6pf1mnN7nQIi1T4sIJjGkFzsqCLt9lQQkud
JC3EewU7dOjmQrS43/tNHrnfEfXnnES9NTswks+hHnn+anrcwvBMrkl7hluAnL2b
XvlMtWgFd4ciNVCKXMkU93S0+TRqo4OwLibRTMylzj4QseU7DII20TcW8YhAuthh
pDmgiLKmEvKVGsFH4Y1UOtPTRrzE3Sw+ezPX6WCOBEIogb93SzBxeT+sM9jg8AlH
KF7+fP5tSDmV3BCe1Umz22hpawUqIlzYLZJ7lwWBnSJNnW0hAm6iBm2WUQ1zZEHg
zBsgHVa/9F2WwOlE9hXuQMP9qiuYa8MgZ09IrHwLhDabIIMpNzW2FoWxHhPhbi2x
+h8Fh1dR3X3/Jm2rQ/+cH5IjY4OuZa69Y+c6TbSgxSWeC60MAAILA9dh4YU7U5PN
fdZ5OyWpavsBXLKEcBRsyVSw453fEEXutUPkNWHSE5jc//ulndoF5Ts6iY/1+teN
B2hsGz1NL2XBSHYtH+z1+l7pTZhFEniEOgjJE1zdS1VaAfabq6ZkvxWIcL7ZXG6E
jnmWDSpHhWJ1DbwGYD9cvAlDv7QQBXC2e6j18Up9W8ErTRjA1+EsUq6WxMSPnTc+
4+yd4jT1ZIPBFbLTxM+XVvlozElzc8Oa9UT97rYMl5BZOAAloxky4GQd7h1VuUOL
VWIgGeoHVYv4axy0aWYrOrKzy/VHpZX3RaC7X5UQxdp0aOkTmZHHKdObFwhTFyhN
Q6HKYFNLMOxmH/tRCeLSdy/lNe7VJlUzE23eF19RB/Oy1JIh49n1oDTkfUHcbH36
ikZrjCUmCSZ6kM8yKVtOuHsnveqYqEwRDr1+tJN+pWZJ3/d7wy3DtIvRK8L8m0Hh
yczmSbgx57JFmrBS+0juG7rGC3WYAeyG+Zz1w1j05nWC6PGr6sZOYJGxdI9aXn8N
TT56WJSDyVlJHUDEn4fDh6txEkiHp2XSLuSUzSrIuwB/sjVv6ew3s4t3HSRNXsdA
tdkShx0ajV4vvI8rbh7UoNTvJhQf9vEaZutP3zse8BQnX3VVfMqXULUeljdsLcJu
KE4ElDqmDDmLf8ON19GJp9ewb2FDroLzKyp05RBjDOtiBYmUChxe54NJ2FtHSOaJ
XTaR5ndFk+l92x2snCTxZkXC6+L1zKedOrMI8HqkZZo9B9RHGdHNwkwnFKdtWMO8
lNoDsEw2FqY9ZsT3UsQ3Lq/1avew3t1yPifgEY9JgfjxCgiEPN8N41x0RnZRnrBm
mdUdbjGz53w5AGZV8VaoguLsIzzkEXlu+eM3kg86VURiYRtPqlZygVMflpUQDprh
XAxScllcqwN4YheCk3fJP/kuoTJ5dpT03rNRaJQfz9X8mjgFqHhG2zsPladHnjY4
XjVa3OPQBfkP8Pt2MK+T4LaXiR31anqHoC+dgaumtODbbThUpmkpgcc/lo+Y3DE8
T5Ufd5/KJt4dZ84SKbuVIBUgRsa7KYt+vKQ3G57j6gkLczQ6mdw5xv5h2B+ARCzQ
Bf+4bLZrhzACpc2ayQv5+WVCISBUtePb3CgBdRIDAXhlJ4XeWsIVxnNN5T/bD1+g
VT2bVi6r0YyZz1U0k4y6DEarU3RjvhaMaw4QTWc3wgw5eOLnuSvCMOvWHo8abERP
Ssajs/SKWDOem/zEOewhcnYIm/gSNEgLCmf6CV3QAZyLEoC2G51wucbdAu3QkAYb
NYqMVQ9hXzaOBVGZeIxSHBeOMnyO9nWIn+7nQGpAYUP0kc18uhstgn2xNqwDLfjD
/IMxJ/IUDsILuWvW4Gk7G5ryCAbquRnDv3r1DzQyiVSR/wj0wpmd0AbfQBtU5PbQ
IAYWimPgi4CalRyUwPcXM9lxMntKhiReB5AuuI59YtgdiqpBjDWMwRE72n0zhnno
flReUzIOCETeYDpi3/wGLUKHfNwd0FXz1gjMbhr5o/VGacr5zbqxOLBMjTpMfwK2
Hfy+1rRNhw2N9LBhsk6y7ZxOQWsOXp+MnMcsef3wgGUEX11PTcXDb3BLSvyv4Mz9
9KtCsdQbymqxfNCjbWd51ufHn4f6CoZtSamBVP4QMamqkowQ4B4AmSRzqX0JnGko
l85by/ceFuIPVjZrCtW+fcw0HLRKbfs22QKvwy4AyQX6JoyAg+2guQsHNkI0xJst
qGvSCOepctTRKI+F+JIuDRUrBIO7AvvuHF83JfDKk3Co9OvmDEV63i+cplRjbt/t
CxoiYkNHnSubwCg0M/5nZXgLSR2uZklLsVQT0+UAx5WYiBXjieEsRls2Hb+GtCuR
ITsix2ARE06Ue+c/67RYT/rYpu12xzl+pyN5FDkDGX9X4+3sado4Dn8l4p3qvMx0
wa2ffnQ2kNvbInqkpZVRv7yP4Fu4d3VfpoHaJ9tJ3/6zRKRkpuJHNl8myezUb1nV
9i0Lx27VRykPs1DblzVipveywenckOlyoF1gJQDsTZhXBWTSynLVuU/U+L1wDSkC
8fbY2sIF6u8ANuTbekx/+DDDzsQsuap6TKbfURWH1cYF4JYrhMi3VseA/17xwD5G
cZxrKNBTTSSURKMboMf2poNjuy5apvelvbJupFMJt7A1vSZuPLpOB2KrwmTfgpUE
OzWUhzgIIdHj5294qnSXMDn8F82ny+4ZfRwfoT/ELwgOwn7T5LD7YewEwTb7tlMw
uBrNlpN0VvlzifqMOM/hSbacGiALwRTezWMYD6pfPkidJRNw3xoWSa5w5v6utCYJ
rH8IzQ9aSPnwfri3/RR6425JiB3Ef6qnkxwBp04UJXHzvbAmNm70jkiRUGMVAzmc
elXXBAPEQ/8kD7uZ3QYJwCaMciseaNVaHuvkQPBUR5gCEegG6CTR+6Zzp8iHO/6b
BUFYO7/IOLmi5mvPLpYeLP4Os9399H7jiC4A8kE4i92s94E/EW7au1WNCO/LI3MY
gyoUg+C7fygkLICDEK9am3mYh019o6hTkp7s3p6m//p7V1Hlx46iBjLx4u9r8i56
BS0RACTu+as8uWF45Xt+o0fDxA1BeXOOm8rDhcv7PZ6SNPBH9RmoayEuaUZMUoN3
Z3z10yx9vmn1IOr+IIIae/t6MbRBaIgtFFdLRO6L83qApXudKDtJIAnS7XzrILgj
fjGIQea3ZKHgUVboXVpMezRyn8Ynax60GyPXkIjrmopnly8Ywt9UWFYzLdaOUGxm
CheHZ29LhhYdzED6Kh7hgrsENF+QUHcewV285gMQ/TECeKgvNslyZzyceUNk2fWW
Gm4JvCSx8Afxq1pWyMqoGAVeDk4xwYVDBw+rpykaKyymcykHwhZu3+IFUk88E8Cf
4xSM3Y+0nf3g4kgN55J3iuOPkfBeyH+iVUHCdpeQ82kXdMEgY3I3kSqFSJvgMtTq
10IP8fvFrvPeEwJ9o/I+YGVxeHE8/o8MOQOklk64A4qaUjobvPUWKPXq1npIwRQF
LMfvbwqC1jylSqewL5lWDaMRpvxp1yLf0/NYtB6TqhZCcQje0GMmcZzG9RySDBxQ
tq4ly3Et2TsDqJDwBC1a0urkqVoQhmuToQd61+8sBOjBS+2rDZ7OixIx1lgI21gu
NMqjtrYWirVsmwTq+Gn1sb2Q3Ickc2+FmlQW3/dOsrUop5Zcz0921VFLA34Pytae
gIIg/RLwt7pzchfBdbL7fOWy3gdHyLRwNCCEo//4ViHFABAC4BTiADD2sSuF736y
C9I3XSocrUW9+C/ResUZQZgpp0R4ZAGRjaCaKKj7I8tjZnFtpvQgyV/Y4iEev+RO
H3YRQuXxzv0GV1crvVfIN4YNNyecwSy7RiyiXJAJ+Th2Uj1JbaE6YhdLuWtcoS35
ZL0n7D7wvOZJLoymqc0mLiyakywaO9ZU2uqbbJB0HCplYdYqn6y8S9pIk7nSZaoJ
lO978/SzVyTWLdLIKiSgoPG6KPcGARb52ssM8zglMQJH34GpuK1mz/Ih/Fqu8ddV
ep635k1flM8l+NmHbDa9CFefv7Pz2Dx59whDLlWcsTk8s/TT42ZOrQ/WLPMDnmlR
rz/oQbOpc7c7zYNO1mS2zkmfqftsOCLIVHYTNVLQ27cHvctpqbr7y9VMrZihdliy
fgFmiImQxwfFNr13oaEkb+Q8+KfPlEND6ueOFbvYknIZ36nnIuUpB8+CNjUBbuLH
StAY8Q9jchBqDpeTWVswWyFhMpF4KNuEaJJZ5Y53pPW3AUX/O7l3+3Ju1onXNONQ
Cnu0usZlyHWZ/2VCuZhdqR41q9HpFLDYCd84zyuHVd43mAbtzT1dq5drgijkdIx/
CRuAi4QXPko+wmHCQapF/YAq5ybeehrith4vI4uKifs1y0rfHzsAsK9fJpa75Ico
ZpYCA9GyqsrgqN6BXKmltyDGfnechNFppA56u3yCsTtayy3nNNJJX2rjHiUc3sXn
ZdERuIqHdcNbv2GOrCcjNXHuDoFXgI7yM6HyzMQvp9Po7LlQJeyJ6Y6hSCzLfdpr
8Dric+6kOO6hNwvlTWK9WzSdb7GBgVa4fEVMe6TLBHdq1F8dqhQXE1H/TvvFz5Ex
TETwIUQFFB1mw2Am8RaBlIgg2RhKb0QOfoO/E86u9QaxXhF+7Q7VbhHtDuaAu2Gj
8FhlHlOQvsHvbl98TzOYpgTrHvu7EGPiCP6k2v5ehdChIO2Ia5vPyofKKzrrQHQf
DNMWsC4xnNV1arXpVdBaEQASsit7d1S7AIHhvuzL9W5OaiDN5c4vsJoslI9pJWuA
sWl4J9WAUHhkaN8IzKn27fbr+oe3LWJyQn8vH5WzoBylxdxU8cPMXJg6hbFwSN6S
xytwqhbiVv10Cu+L9UHHk38DWhZjdJ4T7wsGGPXdyuX78EpZEHV4qhxuX+JIdG7o
l0dnrEJTe/I1eb2SMndsgvRTJ7VX4kbKYiXo+woK5OphWayTJtziuWoRLf37jo/k
YThuJoY9wSaphQ/bQ2c2uCyBoN9iAcgCNXgDMOaYklsUauIRafOCORLGXAq2C5oR
boGQt6qrMsqjMF3c1sKROoRs75mSqTRbLHC1E083qd8uKqAWFM1JX8/qignLKNLq
5eF5lqKouAw66zAAqCtn0adT6FOvauthOFuITQi+l2GQtsT5DM1ZgwVsbEqfKGGr
2uBS7gQWalGDc0HaS8pbNev+dsPb8KLW+voRF9xhekNqHH8mFLyGUsd2pvE5rXqR
gnc0p85/pFp245LTpA7utEfC2nu2rRTO9PiT61o5BS+LdRd+ktI60+GYweqmTSd/
owqRckAzYNMzzQNvSwJqjc1J3+nf0+WEYFQP+yT1B8DZ8xHs42p3cBQIO/RkU/QB
MbHFnE5M30UlaUpzaZ347g95KZ6r3cPUBekS2KMErvZ5DYaa9heF9W4jqEjiKB+t
3NA5CPRfJHRKCJTSsKx6GUPUqqKkA6LPJPbOR6eiGaovNBqf2r5Gfb7IDoOA/Pcw
5Q86qTPfUlt58DzG17/AGprvYuuIb3Xpo3D/IBbFDfaQJGvwGAIQhys+xv1fxNvZ
XSf/SARa+ePUGm2vb+9XzfvNDYYzBKIBQgg8g242XZ9WhqUjSWkc9PyoWAva0VTn
eMETlBiB+i4Uwntt84qSCG4mfHXPXurk37QbDPnbYCDqW1R24KtE7gBvNitOow6g
QW7v83ik63sMokzO2AhQzd5gyXMsxcbs1gcXV4m5Ix1+Eire71pYw7DXE2e119Dd
AXpG5dtvChyTzSknEE/kYmPL8cKKAPKyzZSgxuXkp6YjyaN6bL2EmMzJiEzbxC4o
Z5f5jypZg5szkT3kntMNLGXW6la3zHXoA9L6mx9V6UX06gOawUQ1Y3bXwAt4HndA
HUEvsFCzt6MNFBHmiprKZLAL+NCdcKBwfapq/N1Xi10X5QfdpFDbhYwb0AIqJ+bu
8CaZ5551yn7XhDXzDdh+vMPEECjoZoouReMiQeIpVp/wSGjgCGbIPvs8/Z1kYdGe
TzIiPiN9qK+FCeTIln4OaqokVT++peeoqxbHV2RoNDGMndGTRDBOEE3TDdQFMBC5
08WPbgWrI7Nz5Mxu22+tvZJD9Beo4lO/A5xSDny9Q9QPBlLAaXXNvko2FBDcy0gS
c0UQv/ifHykHRAI2yg3hsN3b2OGhkNsDW6gurvt7c+1Ae2eT80LxCJUqNhz/MiuN
6rcYI03oBaydjcudQFM0aFkp+dLuQbvSSCCQMq0vudU3Cva/TcWmhZXf7SZzW8f0
x35arbFnfAPJiI0xksRepBFfelgUw7de/BbMo36Y65ZHWYcm9hhECv4N9fkIfeYB
ZiwsmnDwwpzWSoJtIua3BUAtZznRYW+vNawzw8k9LMrLR20iXUQzjStNFNzMDClg
XthmX+6q1HtgiujD4T8dLtjdaORRC6dtO0sQBA4eM8bL/LB/RGWBXpIkjP7m+9ML
CsHFTiLS6o/3cvhHPpYbRMaaP+sOTjuFMjTDbvtrXU76jfDZhzqeubD9GiBGwGCQ
25tZvbw65qdU1pwvrlDQMi1HnIn6zBI6Vh+tR6hV+ccl0f0yTERZObgEybvG+tMt
IEjGJFGvBAmAzGiKHoWyGU+GR+woWmR2ZUf3abslHKG2p/0I+l8MoUH+QDmWp0Ag
VYnxYEEEXphCfGqot1TF7TGjEPlWKW9nW0iHV55loPnGgfU0Jq+Ss32uRcxsWrOw
HEonLUhs8QbTlXhnqLUfcVZgE/PQveeDgbQ8V0O/tMx4nkEn0vl18v8CbJGJwMgd
FEjvz5q5wJYU3Sb3RF6oIKswshi5kkRoM2abyBSIv1jU3fg1/T88yvruBuQKuSD6
MVaWQqH4J+QyQlX4meR8JKOlP81EJasm37M7tm/GejGhhWbWpjEKJAU1NmG50SAD
JBGgOezcoMvX7lbj/GMk/FI+MBvNeqZF29AAKlIpIKSIjFsXqPKhn86/yuQFCG0W
8ts0LcTEC+hv0+0PIPw6r234BmyTyrUspC3Z3voErvzkG8OxYcG24Qp0EpMmfv5q
qr4rM547iCPghQuFsLfOW1UmVdZqfyhFXcH71/5qOPxDWgPpx4OGs4aZrWaHsdSa
v9c4yLQ6gq0XSuq1+4WGWtHhM6QCSsIP+foN1G9zRONrT+4q00WxjGs4MDh6KjXL
8191TmJDAem0NdMUTst+A91WBurddSiB7bg13bUGOYiud5RELSDPECPjFtglFXKr
jZ4oFUpeLynOqceymrVJaIAFwcwCevyzZQla0hyE3jWV6BG8qlD8WGEq0NBygTDa
VviUPZEje/x3R/8Aagr8DxnOWUWBoBdrJLgZfYOWgJdA3EUgeK4PR6AlTYib4i00
f5TEokTfGdsi5peqt2cJ2zbR5mVTZt8rlkotWZ/P7IbGdCGJX9RtLdadoZX3sWx8
wQHqAPlwZBiBFz9w92SZEWnBbn6gSnRJUaJRb8i3BkYKOqchyiCHzNL0UbzjOcdh
lVRr8U0jFpMnmeu7xSEfTIG4+066mKpqxqkqMM+hCRBfNHWRverXKu2Cdpb0TwRv
XV1WGt8N6cmVoSRVJCYs0IwlO7TB8RocW07VrCahYAqRi+4ZQt4Nn1nBSaL9IBbP
uUgA4RQS99PgYTdffXIU29OIGucEWvzPOlpaCHgnC5yx/GNmVCP42zIAXlrDZdf9
rqJ+fuuoyHJ1Z9DIi5u6lFBbygpOwFHd1z3AVaU6L/8f0fbtjI3vqiJDjoA5/Tqm
2q7XOQmsEXzxAB6iJzoUgzmxn1IiX93y1wrMIZf697eCHayScsL7WkGIFIqksTEd
C4jh3o+oyV1h+B/WKGwG+cquS1inrbKAlkdbKhqFMNXbYKCrTsk93lJ7I8VCdqWQ
iDeYYK0wo6j1NhH3E7iFshf3sdV6/D7Gz+eDPt2eUunbob0jq+Ot/sWd34Rvro0v
atfU1P6hZ0m0Gytyp48CKJDiZn3HV44nf/5e3rbyvWyry8qEgaP++Rn1fHCw+TGy
nhgd3Ahm8X/Lvj6Bbn2y1bYnmGoeW0V/zMWIk1MOAAXO2YYlkPcMxuBgK95veixp
pdYEAJxLlsgNC6aFRJm7Ir31R2yF1maDCToPm1ZsKypT+T6juN4Gy9aVlLfFaGwV
+ItQgo0s+gevxYasbWf0gLypMmSD10E92H+w9x5ZqKeyYQLf8nmBTvq0gGLNQhb4
H5RukUfm6+s/KlDSCJjqJKGRuOoEy7dJfcEeaETHXS6tGVMeXmLnN2UXnC2fHSD6
9hh2K2N3M1fimtHT6ojWKlV3bsa0XIWlNsANuw/tpxJr+i+DtIr2zcpM02e19M8h
WuXl/Tz+bsvIRY82uDv/VEQ9vRVL9nSNYt+0r6bmsaF7Rhcfr8RYX43RvS319pkL
qGksHBUOV6TDNriKqKUN4+Fa9CiU0NWtrs82sizkxWSnmPQD6PaYK++eR/19u09c
JRTbIWMwfNfL60Qm9r9pFQowv4d6dVW77wfeSwyMsqcXOBWoY7DDwJWLm9PASn/f
EnvTErCjl/PkkuZ/Bjkw1rRwC5U2nfEUscuAFrXW6PUjF3wddeR0j75cdSs/Z5lm
XWtNZsI3zi4ipQS73wjvcNXlnVp1mWclr+/oXUrr7bognPqtOm3W0nT2XBXyl4+s
gPruscom2FlmsesEjouN0s6/Qfq/d7u2ooPvcoZ/TY1G1yY4GtNsMDXZnt+Jd7K3
O6yI1/NNyIE5ZnEXvyX2FPeQjPRSRESKZCZjXpJkyc831cTtX7RUZ5XpogkP22WM
JpXkjt1Tw37NunVjeWTLvSJmOKVg6UF+15M8AwqWnwYB6v/ZIXUxoeAW2CKU/XRy
gz9UcwENnG8wJtWXqhBqQDhek21Z77hgcUx4p8Z7jzuFNF0iDrB/s+2a6d0wnNEZ
JYVzDBf3bwGy8XCewjw6A76gmGAx1oHN0yFGHQ5/a8RlWU1KoE/5TXjufonMOPgW
9diUGo6cYGhVSR0C/Ty66oVqUBbpJ5KSNrnigktN5By2YmdBGqmD9XLxIF7qK/s/
eHT5I0YwdIX+UgpcYZrTBtjkkq/nGGXydIu+Wh84uJ5U06SF2nnoFi9iup7Hee8W
/QwVVs0KWJTNuVQPBYkJ521YzKVlr3vLAQY996ZEY4lqY5cvEq5AkJMBVbHB4Pgd
RNCZRF/878kaFsIERYTLIBiof0ioU8fBUqIvKTlPYTJpHjoiuWfjLkFl9MEmjjTu
fO1UfVvxF22yOfZV/4d2isfjF3QQbBtFyrXX5SOGuT/BIRzqhn93pRnOA9zvaJ2E
rYWoBDbruuq/qyPZvj2uorL3PrK1ILxsaZzUL5OPiHrBh9Baq7wJkXSG08IUB4Pn
SGfedNZwjax+ZGLbQnhdhSCixWraSxUXvbsdduA1T6F/QDXS0jmD+Aufy4XvskBp
kC7c9C/NSuWZYuwdkKUajM0V4bEcXVqcjM08XgXf7AXOkLA2JJd3GM0EHid4/Mtl
LfWk1FBQIoGUTbk36mYmxY0ViSV7lQKRDfcICq4PXczCMhUxPDoLLN07GqJGNNps
/qooAHrPj0Ghs5DIxReGW9WFDp/oB20a+70Sew1lkCGhriPPC71YGQfRVVqkC5er
bORAZT7TuZhxAwSqp4hrZxA6P/pmNQ22wInfl/bB+OBDbTHqvMWJnZY67XV8raag
fvE4rCxofjHLZs8/nxzf2eKcMFJECad7lMyXLSvWvumfyKfJ7xzXceZJmZG9sdhq
fZoIcFaJDoFdU2x0Ane6fwAEbCaO2Yfbyd10f8PVLWp+f03ly9+nU3CLzaouC1kh
4Yxyn6WOLs3Lc+iPitcB+zuNiPAvXo2NZTKsfbTmVe9ZXDWQm/Pq9WwFfe01Rb3h
HARvSNyszCzyQl3f+3P5oE1G7/MHWEo2tXeC/+JwcCb8klYNbIeuo76S4mDgC6WG
/jtooOsa4vQA/uhe/RB+AhaLPXcGA2PXdymLgxU9Vhq3/ctpkmrDeMdDC5VfxwYY
ig9JA9p0RWaJgmy5GpagNGoWn0a5kWgX15RD8GkEoLSLM6fIYmHAm+Ue7Pitt9AK
HdgRRFJyPL3VSbLfJm7mA1b2Azks2oc304yF7VnjrF/er180GRys5ArtSPrchxyq
jjBVTSY0LgYhz0Hxz28zmoeMc+bsBcyPcgkMWPgfodR9qbtVHUFIPGKRTlYzhAbg
qDz6SXiHyYCxWCaRbjumkRpFPg4kzxZpACGGNHXS3jzjKqMPyWD9s9x4M3DOnJR9
NIsSRkvmWEjREa/A6ufULQAWy+peeLYE7sbJBq0FTKTAQRfijMhL5UfV/DsUrpWZ
IIeDWzFsbtUH2+AQFk6k0L0MNYgVaRnORB4npYKaOhCs5Z3OP0rqVq0WrDcn5bTs
Kg8ghs8ZrlKH6RrEE98oK5xngCRKoJY7h27/782ZATl9wUdnd/quuWwE7r+v6MmB
s4RghpOJOFhXyV0Gj3/UZZOIQa1M6HxOgxr2DiMFqfRHxxwKJo/Y9BK2M+0odWbK
Cm6aRwRNyY/djGgzci9vSEht0AQUbhmGfLJeDpjlSDGz97oZTPyuULAJjoURw2at
xZyMKmsUwFCUd2SKMf+Ra2Esrj+Nzq4EWD0H6EPk1q0rV/iPe/5o0XYggpP9fFFm
2XjlqhlsojPQKNlmyR1CByVGhzc61yXgsTQTu65CoAQSl44WsoMb55FyoLF8yXrS
KFOo/q5KqPmZPoLLFMTe+ZjIywa/899uz9MvwOcaAGT+qlsz6TupsSltIbKrGuJj
DrpYUvv4f2MSGKGWUHQvEWRgkjDLPK5PsEGxHs/ghmMmouQT4sBLyNRfm3Yt7MAs
DnmSdX2L7ZDyUUruIuskxizK3gWiz6QPHBx/ZYbj5g2y+KbibWrP7+UFBxHOolTG
Zj192B2VblsR/YP/aLoClAjeWPeafiqlbTMQoFC3QvcBW16r23zGDl1aJ13CYjIW
rACzGG7PtThHNbXCHuZKRR2TEX0Q/d93T+kcryM2EyjWINHqwo5T8hQUE4lagRHA
lQ5O2EH6IrQqKfre5+Z59zv2vyN/d8U2M6WEiFwqU064i2GJI3eqy274xygtTsVY
c8Dwp1Qxf4oFbAXPOt8axm6calAo79rueI8e3rFANnIXQTVgX6BFl40VzfWqoPx3
lRIFwuF88vRLj7vnTouuWA97vNvRhHehSRhKUn3OFJB8bXbUgNSzS4ybR7lSfE18
bE2klGPoSg+4dPriBzo0N/9oeDOIskcyIcMpxjDLm3O9T6zZ00pNACs8VRQOAUEq
T5wIU4BiKZYivwH5/xyLeWw7j50RmYrOd/lPXSeBc5FMV3LYqcWd6eHF2GDVFYG6
kgRl4JA78zTMA7fzuvaWrt/jBBandhKB3xf2Hts3JY8PLgLZ+G1XeRBhQkewtcVq
uGzszTmPR8U+V4AP1+VfbMeZ1bYg3XwAP27fyU3TaLOeDL5KDD3bAdRBW0RZfgL6
s/jpS9/PDcw6PJrrdbGMMwQw5WEVKP7Xcikxerh3pbupAgvk6qURE5bRcWTEAvSq
xbQ6FBxgI+CgO/+kvuUbjJ5l1vZUNCDZoCGGEYjgBKBTfPPuPrg/7+tRlEM894Fq
f29YNWB99WS3veeMeRMOn3eTbRsQFjBYB25G6TF4x1Toeer4Qa6aCD5+rEkyPnYq
+XsUHns1WG9AKKFhUDjZ3M7px1fmOYDj36bfwvEIkrhLz3tvQIH/KT42eQxUmsnR
GGCX91j+9MnhF59oHKmmmT2pmEtvowfGeXKH6xy8Bvm6M2JwkEqz0sk8M13+bOeB
cF40G/QyWUSpTXtKo546G5E25S4V1I2741ePvJKR1r90c9udC5gfZcFZCzuSDtaO
6cG2Hmu7Dv/GmFfYkeS7OM8ku+YgVL1XJJwDPuGVZHGWO4jWLq6QH6cniPPRGAtW
FoeOwcjWnkXfybeanrHv4RTfhQ1t5KhPtcQ62lQeuRsLVPwWybG0QzrlWv2LJZJa
04bI1KFbt7J45KpWymOpwKy3RKyxeoZwrQxmdbYaHrVchddKUZNelHIE+oQmA3sp
ey0HPLVy++WZMY0/B/Li6vbjnR16OqwVVgpk3HM+0z4mAGbnVpSQx6B9wW8IXMfY
RUqPvWEFxS91Lsw94G3FHpxZcVMHOHlGJofVtHrS9r4JszsN+sVRR38v869nvODA
jrs+xBt+mrZDA5nTUSDLkEXe/nti3mt6iO89/Ty435vozjcnTGQGBdlJ3KzC05cT
c/QtaiwQ9hGnEhdx+Plz/HMB4o225h/Dm/V1R+ItwY81KZMrIKvjb26wRildXil2
FE/S9LN27F1LQliu/JBx9fgEAMsu8rjKwmIVFjPZzRFmRHiUHYGjJrgH5yYKT5lI
hwhaTY0YshLkjWeqWt6K3MvjkENx9WAPBgNE6v9OEpP3cr+zXMIb1Sar5P9OcJU9
h6oSzOR/XfaEnmBuhL8rYIQuLmTJRd/Pkr2karX9dE9Vn45JPgW4vOcpiIpCYvCG
So0CLxSPp0rHYoO1wYEIgu6Izt1wVgCxTbiyEu2QI77z6QqB0HIxoFkME9NOOqps
fQj9py86I4us4TFTgrAkZgAcM3tFMSOZvcSi19be/+H61XdbSVPJ3EPlN7qZF3tm
TFQSmMvtywOOHwUuMi94uqMM1Xto7yDeugEhqhCuljeM1VGzP4t0tLfGsPN3pJPO
/l99dP0QOL8zqIgdc7ve2EOPy4G7cfSwHLDj9nnYSpIR5OwpTM7lROtPMs+gDcoc
f7AHpQU+WG9EAhUZW6EShb0dtGDo7xdmSZu8Am/388IC/b/aAO77GtbtDwXn/Dfk
LvgR1VB4hMh35GEtEZjHwzwgLN/b7G1xN1D6VE/ye/n+TjMjjDCzTiy6m1sUlljh
a0G0ZxI7d0vC43wZDphfdJi1deUoPiRkwimeqc6tFRfndPoC6pMRzygWNUzQwSe3
ETX1Wfa3LYIdWqFiUzAZQPXJr2PHymAOGAvEKl+K+hg9myAbSGQ/Cd4nJCiqVnL4
k+PgBov8epiuaOqj1tfrFoqgNZsckbQQ4k44DWTe9Oa6tDb1kePagjzL50khBtWm
RQPpxLCDK/4L2oUBmYQsd3DG8s7GWQLNdQr36WxKrL0+779+X9oURf16hYeEuBer
go7eBNZabrmkuqk5A/LwenfoNVK4T0wDhhABAAjCYVf+SyVWoLR7i8trnnIsWUvs
uFba2gFC+RslAjMdpWgQ1TsetzsmRfAn+gPLkZdSR6J3ga0b+sAA9DAko4HRDVI6
dsNJzwqnrOGEBUHsjsFOdE3Lfl3OzgNrEwKzyw48WlRATS3cq8BGwuR9mKD2zbdb
vw546P9/h7tDAqlMITm+JXb2CS3PtGGgp8ASzztZ078J33MTMHzWJYArk88q1fFi
n5cddqWS/sUDI6mS+yOHKMOPAq7LPPgrbSu5hx9EZJNHX7rW+ApzuWug1cQyd1Ku
HvETiY+lbWKQOSyUO7O7kBteBVktLFOKyMIwnzWjgklQnphtwLQmNdeuzEK5+ngY
35vpRn8aEzcdRTHpfyboz5yv/IoYoMWBvAHZnUBq/34jDJctQbN22nSoUYgKpMhZ
uzVZjWrYRiMoi25maGCEVAPqRBJaJMXH90tnXVZkLI4zcn+BKgnVCe975I59yGkl
EVCxHlssSK6x8rOnrOeUrI6mXLnRSnH7NDlP0Zdtt/Fy6reXMbjuqtQeoUkRyWGB
xR/Z0dMaAx/Pej84smYaYFMmcqKJhwqiphfmeLm2Kg1skSB3HcXW0UPCeB0oPtCd
4iw/cn7hsFlJChcbUArEFnWGfDAhKd2X4HIQ+zumj/XMGeUxXFxF816pthaK1I5S
ixQ7DWMoDe8zTatyRo9JAJOiQ/+WMxFOGXBksg/rzM92GGZkmPR8IbOsIwt03JQp
7sIo4JsnyvjcYHp2tfCKtNh865YwxJjgM71GDLyBd5Sqg+adDPXrN8Q/EiLGi7dQ
ZMHjL21BabUOTdMq+c+EI1j0xB5Xy+4OAQsC8O72wiI9XWxHUkaXiLNIVveQ7UXB
oaTSDTc4nmiHu/VUy+PpJmPg/3OMaWsRZCGKLpUTqute5R6wnnjDqCofVuS3KCKF
9XN9FNSGI2Rxk193pS0iFkhHES7iux+sSXvFsoc1bfG1Ou2WB4JSetTahRufn9Y6
rj1andO7EGCKVvteI9dpd60vddNsVPslnmrq5k5S3Xoo3C+2RSQzbUzvi8eMoGxa
4Erzj9hX6AmfkZGXEHCaUPap0i73l76Be5Wicve+DdU4yr0x8cgWO0CRDaeqba+w
xA0lF2G5dgIHJWNynDkOLJdK1F0Lm39a8l6BkpYvz3hJjFp9cSmTyN63Vx8sqy0o
v0cgXjvkiEZz8srf4prxoELNqh/rRebi/VQZFIj7Ka+AVS6B7hcMlkXT9YCniwIB
9+kGDizFxIWNGyAacJtQ9emuNGYgBLxCXPiEwnA7N8l9Shd1Jy9YgSJGOuLCvueC
ioDjfKrizuSJUFyXrIfnmN3aA4+FoJ103dh/nUV2uEMNdqa1iL2ewli0tA0dB4QK
EW4YbNCTR/5+9KpPEWTncuducEBfcVk7nCOcJkV6rVMVst5VMxdRrPcUqU09/JYd
42D7jLoUAnaiYi9DTev63LZ+61kXqd3oPYHXxSOLb47F60ZQ8dAiZkfpnWYWOCGL
VUW8WpkhVz5g2whcuDoF6lLk1dRySu58N5UgZEMS2tE5b4Gf5oPHlwSjzkbUEKst
WlH5sEsARC+LuR2rJGwy7A/uWucs3kqdXubM/xPdkPmQidCgmkQdcBCvCYAEKAMy
Y0TjpjXLUdt5yK8uPPkvQhSLmwdIlMhtbMJypaVImq3nAhpFFvzkocP2pU5edN5U
8dgWmtAqafPZleB6tS9N3ZBSAWehf3r+NFxA85gOaGkXeeVILSHfJH9jX+1KpExY
aPa4aQB2oGrw1wTZDOddJn66xOC+N4+N2xn47bf5MXeuLf6z8S3nf65zP8nfprhD
JPY9Khai2KOoq7rq0XGrzXw8JMgWJSDFEnMwrZefa1PhzwNk8I9xxEqHe6OMOgcA
n2u/tJCQLdDyy/dTmH5aMC7iseEIKgUiZT8i3qh3DFf2GRthhJWQMVMbReH1TmAB
SjJ3q9ts5vnq3W8B6UZXrVQbOV3rXfJGo0A/frq5fAoLJM2F8h/k3rLY107HTpUP
87fu6Up543LHEZVVdGH3Tois+3DraoiGtwlx0qfn5jTfQ5KisEeRbQrBMlgEZbY0
/seGOkuzMi9mkawAy9Ong4Av/qVzzPy+Vho6PyPnkAmQxTwfgKoV+AzYpp7mYGq/
yGsT4whZvAmfe35dOnjJN9tzy/Cz9qsT7os6KeNPOy8M4OcUC/PQSgjJbWZAej20
7hMIlIuuIMArMH/HSikMofUWC8KaG018CECA/JG6tybqVUq7NbITqH8H7LTGZPLI
MWOXrvs9oCD4PgcuLnitlBidvuVb6l3IntEsHkbUP4haCGOYAeU71pwU95mxg6vB
6Jp44fwTdOR/zoKLljDtbA08Tp5v6SjpVQTvUfAcNXQ5jZwCJy3J5ucuvdAviqwL
cVgLMi8bMryvwQICbBtSlgTgG/RjzBPkdnUY0R23qDAQtKrbpp+l8vDEyAbQ1nmq
uLFEBz5u/4qqYX+nrbCTcURoFf6V8eI7X29WTEMYraWxNcoKpr43BP8qpEybLvRl
ja/z9gFHsMDV5U5qSGTlTWOwIBOnRXTGUumc9l2v24/p9QoqewCG9CloMpG/KOij
fMH52A5hh/Pk5/FkKHiEQ1pta8UMh77Fiwv91vrLzKMShbyBUAXk0eRKFcm32H9F
ifNzP7V+ocDv2pXAw5apY+SZGl2LdLPVDd9uo+4wZPENtfbFRo8lQqYuXJbGPXKy
dvoXv1R8bICN2KqPjIlfDdvN88tOGmOhUm/DZw0ze1P52uvsRdJC6mRNHvypxNvt
nsjCHWdZTMpvZY3SFxqWPRqtyJ9pE2+QMoZGCvQCLA6r8XKINco5Y8pc/0aFUSbB
k4rtOT579WD5iubhEZJWWJIh9KJHs9aMRRnTr0K7htGIUnzPBcabgdTU4HpCQ6Lm
VFCKAGIqsjNdQkdIEjqyhi+ZCbh3kNXQ2UExBqq5xyvj5KNRlPxjnN2S9yjWPI3K
ncVi1J3DtAMMRnSPSP4rJEUuvYXvPVc6idXiTzoNYtdqIF1q9KBCOIfgyRJnES81
hjsI3YVsaLw9gpKYPBFDPostjaNlwGwpzFAbsByA/KYL0wgia3AFi0hBRZMjRfJF
5GpGetUjWJTXdwW6tJcP2W0xRvEMb62mLVTwFqu3CUCi7rNGZJF0ocM2PhgQam4C
PzQ37ugFFtLvbYbcdp4wJttDiGcB0c4ihBJXiSt3qagCT/HCviLHYfheLHzk431p
iBa7wRKowot5qDDo9ev3XhJjJWjT8piLdC3CnyDqbvP885Q+e2baGNUwC5sJ4pCd
6++U/xF1Igr+8qi/FTG1hLLXZxLE2Ak8TwW/OOpqk1mYapF+nNcfQPqaooK1lv3w
5SbePfIpAoIWoJtR7ultAVN0qYgCLpvbhLn2itBd+MdxskkR56ELaCbN81JdAKjb
Gr4IFqjDrw45OJdcP/Xgbbn+HNdxhbgLOw3dYGLySPGtLWzbNQ1EijALaLxPgskq
U1QuHFjbnbyMu7P3TX3RQBj7h0nQLp6PJXOy5jiO8G2d+6XI4EtMcTn7uC690ru9
v9lIP077AtMpsem4VKU0Jn8g0i/R3cu5d7tBbDmW1kVfkFZuqqfJYJwltN7Met72
mTpogtRyXZ9GLoChIg0xO3nlnzBdwYxH7ftaYagJQv3d9LzvNTsSUinYPMfADxEk
F8A4+iLSDQVum6J3niFR9iQObGT9Jm+gkv46AA+0ayBzZzM78AoiAk3VRmUlQIQd
SlqWObRqP/YmlLBnzmbiETf5Ca2s9AShgqplOytP3al1AZEFyrCZJzcFWQfjTcyv
jclXwQR63bYV45LlkDyHvVHCgFnDJvwWPcY7jTt1z1klEzgGzKMmiHkRSbUx90CB
7kN756IydJogvJ+UYJqkfGmFCeH6G685Z2m+8AFiJO5JlHduJ4wlsKC3CtZATd9S
fBQBLsmQb/nPtzaZMahF71RRgPTrWNarhVp86x2TXvX6fueagpZyetDFwFuR2v3t
9BCeBXT2GqDPWI8iMQ8oVCbDL6m4/9V7V0ZS0T5i7xKWaLneDVZyu/yubDpYx5Ui
qgejhwq16ly9qQaQdZqycDfyIIALbFWOaqe4UrWLa/fG3GE3fdCrUmZ6iTRdjyaZ
0ME/Rw8K5i5NmhZB/L89d7XO6Ryir+32sDBQWaMngppWjts22D9WlIMcUOKuxNQM
503woBpjtWBWq+327vGfW4UZ8aTCLx9rpWCDgt7sOs+QxSTCIGOV0sA8oB8xGFjd
rTFKeBcOno8U/7T5G8q/6Ywrt1VKFHncA3FoXICjuC63BH+DHU/Cz5yy80nwiUBb
IZ9+M+nR4XNrICH6zAqzkH4srxHoO/D5+jYG8cXjdeol5adW1jiZaSS6zEIjn+f8
Z4mwKET9TUpBEVFjuXiMXToi1X3Spj4Oy+TYyiF6uIz3Er44Is7BiMepyVjC9N81
2DWAYDspCsZdT4PYrvBHT/uGPJjlvqMlMQ6z5F/2t0OJf/XOD2uJPRBvyz6UWtXm
Zu9NRZuFQdsYDJdZXw5KYsaHzeCvfUEegxpnQ/vVuzX1x5Y0j0vAe6eZ6cXEBah3
WH3yGBdVqusc1anj5NFEQQbSO/LYP0ZFNoSUGyS2QEkoxn7+xTr5QSGm8y52FXPK
xIxKIS40YS+XlUOzL2Ajlw0pE/OwTuw1juqX7P4c9xkjr2plia44s1Pm07xnfO0P
WWU6/COBq8N6Fly4iHPzAZUY16ihzLXxIOvsJxxtKeF8mEBDhbJgTM0+M+JKny9v
BNli0egWAYSJ47QrMhtrl8ubnIL2NOGqf913ODLzzst1Qe11pl7zW0Bx7kDD5s2u
4k6ScESGtecbaetpwoDkRAp66T05KbG3eQKJh1kYsNVCqnz6G3b4VKvco4N4YNpw
hsmnu4SPIke9itQ5+hOJcgRuBtb2+A9XJ9yBdfqIFqqTJpf1461ndfO/iEATSKMs
1eVYq8n+ih+3SaiICIt6/Gg8oXxpsuhWLYfLXcgKGM3+wAKK9SpM9eqmqsBT7J+E
jtQ1kA1sFCdqculaf+MruNHoMAcuBgZV2Eaqu4BeZhLix9xu5vGb3TyxmSM9CKUB
Klh/Zc7MBl3aKSkAH1n8l6ekNOE4xFWwLjiLx/jlwvdEnRLWsP25PJ3tRd3Bli+Q
ysquQkrKKFH5zPkC0L0scWFfCW5RZh5xDMIuScfulm03WEtgpCKFyGYpj2GxC5W7
XFPz126NPMnd0ZSi0ID6aZQTt8EtmuvBBEq0aLxs6Os6ORAxZLi/7vMY07NrBcJf
5iu6Zn8CDrt7l9tE5M0gGnJ2KhGDv0/OwKeTeBzLVPrcH1X5ty6UeatBBFsMNmiu
VP1e39y+5gJbDDXhs7dPZL2HRy3unwav5++NihnlLkvTLas6Asyxfcyk9FYfe9B6
KH8kK7SWyG9iORbnEBg0KGW81IQDhNnzc2Vue4NK+S7R8vIx2aEGcx3zoJA6KeVs
R3u3bB4u25E0H65HbBagdNW0cM1Plpc3drtHUwwrx/IO2x2rOOcNE6V5r8mXgDEI
z4tezQwdT65D7U5D0h/wAY/lWhHEDaVuqEIHYkAYHYbzTazN+1NBHG9MB3nYzqCw
ceqtQ5XGkKmRfWtuFwNrto4dKzKYhNuX5VvosS2GzNyiyaSisATX/VNTFb8WPHVA
U4jKYZgw9PyiS5yVcKtbRJ2daAasz/FXVM+gyFHA5+CylXpKWBGt6yPXWqgziykn
xV1iwXbvCxlTYagaFQmVJbDcMC8hAUis4yy9g6nsdH9iZZe+PrvR/IDYWCtI7E4e
KhbIl+bx31/ATh5QiQ5ni9Ji/nzz30CqxmAfRB/GApl/yHubQN28scPpc2PIh/X6
8TccQC0oxZEueemq1zOTNIt9Sx3YbxcLb8tU4Uxxg5LjUUYwssmrUc1I7rVOQ0Sj
4R4sq6hf2nS5ZX4O1kOhsjW3ca4t92V0jNl8wv4HjNKRWHitC0IpkorqjE9Kk6vA
mYw4r3RrC8uNKtqOA9m/x+Q8spgsr1ZkGcjsP7ZiyxcXuFQT8Av8zHZwrFFp/WSy
VsLvxUFOK6QUr2kthPdiGtamtbnwi7vbUNEUjYes3quXRlj3ZO6IL3zRlnLeayBD
p68bXWyrGBngMLPpWeV2kpqAYKyJ1v1Aah2s59SQh5hZmwPQR9JySCJJC+yLBf/E
dr5AiKR7GZkDMIp8zfRk12GvjSr/86Cms5ZXm6lnLEksp3Pigs8nD/cp6OM/3LG6
LMsjCdR+1QthZyMYrsb30VXjnObHFnsV9tFCYSpzg0IGx1vjIZkV5CvI+PQiu5oc
tGuv61lw+kNfhNUzNOJSL5fpAfEFNxshOGzd1wArZZeMdI8ZZRPwYF7lLyqnK0g8
2zAxuMHyIescfJQbO6FTNo2VNbKF4nC1aEs0jlUlajpHug3F/mswXagPws1HyFi1
FuMZ0JYrm44xWuNRrs96zFJpccNOfqd98rC/QtNigd5ljY7Zq6KSJKnULC1uyd3N
IrbcyL32VyOtr+rIVC7Ytq4bup5OHkPU5fPg7D8/zG5Bxjqf80MouOIW87giaMi0
F+MZI5ojNIsVl4c1hX6hs0tn8DKVX6scB4y3K0j9jlC4glixVLPqylOMybw3Ti37
AoxUkqw8dH+PRtHzG1/JUxnUZG17gpyWmJCTv+mFtBOREFYDrsHigvjw/h28sK7z
AgI40ccf4gl06rQoorvfmbjwUn7oOVmjdC5pr75y/UB1oW4ZUbE/LSyevGb83y5s
YxTmcAFRUNHY4Xct42fbIuxp75HFRI1qwKuZ2zumCwX3x4RJIIcPk+hqBEYxPNhE
qaAeJA0t9DTysQH1qhWAger0S90XtK2x4SNMnwY8IO4ecKqroFWQyr/ki2hlGPAh
oQbLiFHPj/SVkF5RE8Th0fEm4VBD0hBR65So4fmoJJy+CUjmYjPxG2maHq82Pnu8
jkmqSz95q9o0zLi0uN6TxTj/QbiSdRgBhulGYwajmljcOqk8hN2Jk7mpINElQGR5
/FyS4eD5602oVEGd4zrcizT/rkedkl+ojvtbvCW4dDOJYevt/1QKUWfUwQNPnRKZ
j0yQvm1DU9y5SwqUzfAUPPpODrhKtDgu9ZQaBiNt4acGiMU2iWwlvvJhM9b3QbCq
04IDFXEjHxARTn5hEmBWk7DTyPLA6hgmJazllnb6IHoLSXhN9wo1i/rQkvyqkgZq
tQX60dLb/VOJLuKE3D6wD5OoGAsYGBIqNssIuaZPLg3JhJLuDKu7o2MlAWNmOA2a
j/7MLYz3VK3FsNMS2nc7bgkXD1Pd104ov6OAnqtxerAVdmeDAAm96brD+LBCx54U
r8zr+wuU3MMi80pJ/dFz1qeUFctNTjP/khLygbcCUAnwKz9gnYLUstRtb2CzMF9W
cw73hpOyih05kaP2NoNAtXzIrdprXOCRxKI9lX03NuZqm6TQEK8e6u46nC2P/7L6
/B6DQuy7TCHWlmou1zaEztmfOcvV+dEhxLoQeNPNTQp+8J8gaBTHu1UOLNs1797e
Wsn74yswR5zkkSY5ct/ycHNjV4Ol6gG6GrnUp11rtNF9as45CScIOJr0FyeCS+ss
CiZf5DGsy/C8818B9a12kRbNoYjaEuoADI8Kd4CWGE8wvwdIw96kYHmu/0J8mGLa
a9/5p6UvGPLwM63eMrjlbuDEZVm/WcNkrfzMP19/RL6QYtE/Vo4R5baef/ePul7Q
6byp9JgHzKEo+h7ZUeecJkTd6PI9ACeDGfNNC3Ok2zJ1v4/bsUsmNjq/XAY9mvTx
cNuPHVJrnB31mjbj/XcScpOu7+Mhh2iCYyxwjDmj6GQ6I+3+7ayl0fTb///4Ap6S
ethougBWNDJ8GNYbsaiBrN62UJo917aPEaTFNzZ1zHvLi3b+AgYhKVW5Ap4uJ5sE
ZydAtKXArI9+Ui6Onc3qK+/vXA/kxS0ugK4jgCMr8ndPMUfBOObRNrrExVPPMz7S
ecvVUbpRBO4rdpoRCSrXNxAevadMKAMsypxZ/klVu8G0ol6C15pfYKYuLMCzQUwa
F4qZtUnR9WeqqDiKJvkWUPsc/rKXZw3Twos9bNILowFDsvdXIUU2eQUCL65VwBql
m4Zi/+LFs0LgV3tDJL79YX91fAOXYKydQebnQ7JDNvZLSHZ/P//Du6JUG0JqGeUf
C/+pW7NTyXpbqdnGoVNa8BogRju5p4YUUMFt2Roa3Dfjy1E6IccecqKPyL7V/e+w
Z2cGizjI8aQs7Zi5Pkjz2QDoO9KFapfPmw26WOywqpQn3qIaz0DIvF2uNBTiwBnx
/0mVIfj5vj1YLCbuMQ3GilN33+xeyqyvjI/hgCnGyPsN6savo5OiPPQG/KCNCj5I
lJRILcLxdpUn7vh+ngY1g065n5wOWYRfY7F/byqwQ8gWcWYSsz3wMPakzozsnXQZ
AlRahZzTroG5cUR67vF/HnYxmtoZA375Nxu6EAHcXcmfOsuutbOBD+/gRs2MVrbz
tqFqJVcwvQ+4UIk0AjPGIQvccPt1kVrKkCl8zZASffxYdIeyC1zBqmM+chPz5LUG
sfviC16qZ4Op5GMqOsxRG1du0EdC1t5XJiPzx/EnOr7Ffe5oYpM7YnD1EKKGzzME
/0FMcrt1HCgkHbPvT89/zKfgIdXkzXq743es9lbpCoDQ7QHGnzS3BzbphVIIbuJb
BHapSnjg81Uw8FWtU+nq2wQcRCXnllDYH+r70rBbaBJ7RMn1+jGaXtVTfAcXVMHm
xXENhDnQZWgB7NWx9rQ5Cbjrq6IINrc4pWr7hmLNE9jfwIXDD8Conjq4iG2W0OnB
muuvzjty3Y2dyXo5KfK6ieZi30BufrrnrSHjQVhhZ8nbQ2RQzACmxHO2E8jhpzFV
8tnoXLN2U4O+QabEYoLdluCP5lm1gAwMZ0I60m+2zaEXwYem7YSZ2Cdx0O3Yq+U/
YzEvw5dViKbhEPUToymQKGAoSZhVOvhfIGsg6NRZELpOJisBYvVUo1V7VQltbnMz
b3pMhoo5TedvT+GGz8iDrJVgdYpJMrdx5SGjKSKdMcvbCdcQ2YwvrzfCyG/ey4DE
bQYxz1iEmdQzLKSiQ90dqS0xtVNoI8RaXFcbSktQYz4PTDrvMjbTArz4ajhEjemx
kXEusAvsxDahRt6QT5qUDVSCE+eOHv0A1VeqQS74G5D2GicJi2bDV9wrXU0c7xBl
AvW6EzbhV1WigK4u+fyrAZ1Sdbrp2fFjgjHzOc1ZSZTxG2iEvUJkGgtN2c8Cyq08
1zsxlrN2yfOJzMDvECkOOtTFCo03/h4Bue3Xx1yBOzPSSexNwf959O3JoJL0A8n6
kjfwuOHS6VnsglDZyMIHrZwAmDxpzgGHa3/o92MQSKrNSjLGo5nkhHdl/OFb0ESo
nB2r8MPeUtUc8efyJoEHRGODdm08tMpeV/F5BfmTE0ZkopCkKowt1FJOeXFyfRwC
xiLhd772vwu9ImCpCnD8szPiLQhPbog8UnAQrkIiYvi4MIgAcfpvFFRBcqvaDCAX
MfIvM0WweZqpFkkWDwASiiB9MTFNA+Owj2usHMVsLXJe2MkSurgy/qlmtQSV1GPw
jx49XUPoJHsPQAhEb6YXXRGTgA3zwKzZZS93Y0dtWXJ2kj05mdryyfPZQM3U/rwW
NmqlXXcZOMvY9u1JY30ZjqjmOVfjkiBnD7x+l5L6p/QGPmLC1+jiW75ND+hhFtWZ
9kJfN0CZ17rsKXuFWg6o2d6vaCHDIfxeUe+oWOMYhRlG137K6tZzb6LoXCVsoaRP
fTuShWSsC295sQpFl9twvUNddji/ry2NqCbhAvvhRbusNU8u0/dtwEvtGC65vdqX
6qKRpD2Qu/8MVEiR9QRTGA3Plz/JZyMvjMoDN8q6QO5XnP+jdtFyYFe4mLA+qHOH
KYGjugBywtYakJv3ROhFSlSMRu0p+pMalrtxjafIsRAXCwp7fV0/BM2ILIleZp4X
BaActJ1kK3uFn2VInaJT2iCE43+iNm+87JobA5JvaQEk4GEOur4sV/F4a2Vp8My4
qD1fWokFtxbMYpPjiU2tInt8GFG6dMrCRd1gG6dJ2xI70I3tcKMCoSfXvLSnPIop
gEbIzDP5msE+49zOCb+OI42OaVjA8559IXsgk/wzUptILqKxSVpMuCoLukvB3aB2
7uXqIa9yOKOJGaLbfIPoiRs9cOrcXJ+VRjojnQaUZ9zyNiw7NMCo8cyewuT6YEZC
1arN7EhvGBI9kzuX6jaWQ94wF/GUN0jg7nrvP0BYgkmWDXA2B+hh/fHHEo2qHlds
cjr8GzczC6dzEy14Y3uUcxH9SOl/NS8mIO0cxX/jpbobpezwVyH19VB0b2k2jN49
+7+2Wwr3PjGXPQ7lZaplfKOTNXrJ+uBj5996utattcti8tsbtfmzGNsfqhUjhgaJ
A2y8YWFZR4iDXlvlK0r9lYaWzFuKLz4aBtyZIqtTZe0VnaEp7vPVl/1b2Fdhki+q
KN4iKhRd4apee91KCD3ElBHvzWs2I51+L57fHc5OX9J7FQMtO1shxl+KblSul8i8
qb/lAhI5l48H6/Qna4/F9DJramVWZZIu2MY2anYhyPtlzo2imoJmv9tjJVvoLWBW
ZCmubrqSnb385NZ6jUJESu1VbVh+8hyubQbxxdq0nQRD7REelAdwvr7+Elihc/FG
6GN5Cm18zvKd0tD895l1eV7rHoQEK41x4fePvDobvwRGzFGivIezXGW5Nt7V1P3c
YNEXL1qobaYd1UaNgAWhjRP54+Jar8n/iscc3UodCiaw3IXZbXtslDZv7yC34vod
xfDoOSRrPbKD6eDwofy7yrGbQ+M86aAhOShV6p8FT80yLkuA6pBv5NCTvP2zkjH7
y6SvM643pVJAtBbS3931tc22qJ8I9jckOucdoMqX6A40jeMvrlA2EJWX4yCy0GZG
hrEUsdiqyzRlxQ51QPwGwGelgs+Fhx5+Knbc1AdsiTRK9FI3PgeRkIZITFA6SN0v
MZE6Us9D3B1PV/g5HuqZMpVrp3Z3LaEekym9tRZmPChxLBmF0Zy805U3ewLssJsQ
RW/tuZfMvBlz+gtB6fqic0P0oCkiO49rCPhm3nVL8QhZwzClhN8feyMBDXHaHOjs
Fuc13wVoBNLTSafYR1NZ5GYV4nZ0V4VnVa+PvQIVUDan6ncQ4c+xKjmfQXnqcVza
FZMFEximbqbytWcuhqhggwzgSP15miVYm8mBNlVJHYp67ftL9Ch3Q1eHFGHEsfYZ
btvaM1GHD2gPCelAizU6OdndYjUWg74T7VRs0BS4BJBZr4BkNvHQ4ewJd8pmlUQx
RqfusistalxhpeceOKjnM1PU/xAah1zQC41hNhZPkAdRxn/RA0b56icRj4sB1OqO
mLqyhMp+/DiB19vY4oQCglrFz85UJjpTZl99PXvrt7cjdFEnllm6dekvEpA5dHNf
oxhBu7/0zyup/5km78I3VQm2auAlegHRln6fe6Pj9rRRzUUX/goi03jmnw/Q5bfU
tMmzZQyljYR4ivvfZO9ZGFK0ddLoiNuwfxV91tKH0U/rF4F6q7zQf2uNK2M/j94R
bOH/9yuw3kXevnyooBewBLf2aYOVnhKXg4av81woKbB4o2dS5ht5ENbPjZ6Jh6I3
4vLFtidQQWaAkIZGJYsCWgR/BfaDXUr9i29EM2xqABrPC5rSww0MkAmEf+IcGztU
o647Ea9tcJwHGXo0Z7yUi3m/hCKC8anB5jAwNCqnWBt+mo7eyPYWzJj94YvmErNe
ceWE2DwJ5tIBkJNz0LmS4TVBbzgHeCw22B6JT89kY1rxwVJ36AYjrZhAibKgq84F
dO6er99K8Z2J57+E3I/pmQurrQHgtzrkY0B4qvsXMuRZc2lEku3nPMLfed89Kk2n
2i+CZ792dWeanQUdMr0ctX+VRb3/AQ303fV4Qw6QLSgdEiLigHg53k7Ev31mggTn
LddokQW7VSgg9Mp+xDIszkNpVhbSIwTGusKO+l8P1olWFGbhJ9/nuyztTD84P3W0
Pfu61hdDff8aI2bOKWvAV5lIAhtc14LrGZTqT9nXUyISmWWJ2AeOHcW/LzDb2I8e
hw54zFIqE6MXagacCvSYDqfB6YcAty5Y0m+1diJdXerdiO4QVRYgWpWWRr1i1n/w
M0f+4WeXact7sKtz53RdCeswslEcJEzA4YTz3qRq9tPlyRrfrXV6AFCrpsW3d6wN
m7XZfLIAb4cfIDmWvcKfirIn8HQqMRzctFRlmR5o+ZygeTooFIO4Y1gye875rmvd
k6nVg1Y6nptwm8oMSnQ0kLPWnpZp5auzn+0oTwDeW1vwTrUa+DglvM79BnhNpD/Y
3MlUFrsbL32XQxGTYW94l3q559t+f8BQzmYsq+ON21OrBXQWSvBgbEL9ukozm4OG
pHNygIpOTQ7WdIlou7vp6jonqjUtJK8hEapFR4rLaBCVGs+D6GkxVntVqO0+Z/Uk
Y17Pp3XOpZkwZAejWCRF23VwbHLweL6UieV+lk/ifHCvb2uM0lg1ptFYmMjOrxEd
nGyGUjg110WnFMiEH51M8fshwmJJJWfSIuAUsYNFEGQGuM6WbHc9UWxvyhoWBNkO
roFNqvCKdKXZ3pMbCWrx3blLEkwvNMaUM/0LxQASVt9p+iJym7HbEF4Yhi3o1LuQ
jxzhUQ3VWpA9qAEMPNOBPRgdOnaTIsTis8sFuMR7kstujFyKjF8FuRbbIIEahaaB
h8jMtQWUMlwSdxGjMGfvmtQdn4SgSg2EL8NpHaX68/XhZ57NGtPPdp5DDmwmifke
4TlIh93CrZCgzSF6iJfJIdK9F9UjrEwnAqmYLoXif2nLNAme0X3JhANntMFGZXA0
s/JWQzuZtGjT5fReQKLRzgpiPbThz1o9vS7E5G1SmYrbxd7AF3bQ8jhQG5bBdjmh
2CDUetnQUJEd8jVKhJAqR6Czon/sm+WDnQ9Su1+v6cs9m6LZ2WrVMN+WZP8WoBpE
Koe1HqeXjFq0xaLKTeqznzM0Ou1Spl/C7HH2rbijuJevjwjrCVTZZLJRUOTChYLW
cw99hoWoIwn1FvmyTzdjNorGqMj+CM+OmWvKEJD2gVawrr0kSHuLuPVNetRerNoN
5MH6k+C24d3L9+lL5sz2PEHx+cFVzLtbgNRUU4qoIwjkku/uDJ7c4crmjadQUBHL
w/B1F25WgGgR+xi8oJfnqsrjxxOLEx5YPKMMmjatSsQzOhlpqG3GXwPuY/C3j3DK
ak8sb0rUzjyMCs1lrnkMCAd/dPkpoaenPHVhD+g6iWRfrhx5awI6vnfTbWlp60WY
I54HUdTRmarAR4zVeIGllT9Pf5vFhBdzu94k8M9FUlm90k+FpjN5yR2PrYfYoBLi
1J4fqmXnZEk8Q4MQ47kXIYyWgwb1QIMIBkGj1dM7d8fSdoG8Nu0mB6EYpKDI7isP
QFC+StC00f95cMjBZl/Pdm4bQEakF8Gv6ZxVt4mVZz1zSaO/4aasJ9UreQQvN0rJ
oKCouzJcWvXoCXZYBzxtqK+CivCkDeXupTN1Y8g8WTnaBS1wy+L9gONpvmh7gNoR
sjBIw25soFB62kkNI4j+7WHkRL3HgblxRLAkn8c/bKHgdumhlDCLHjDEOV+evI+E
y8Mvq+7ozScVgjjx9gtn2XMkbEmTUpQmAKoQek3/DedM4mtuM8ZcGmgmTLsqyjXX
7IhTrrvJKDaDkssTyfpSdo36e5njDCS4syk5JhKbI5wYF57IgAYW6HUDMj7FnPvy
wOxvWhsad6mmaSlVzoFvWIEAzEVn2HxEzjDffwWdWcS1guL7dVXddE3BWBHqw7WV
HL/61DD65ctEjVluWZws/nKBlZ3q+tYLSqWnmmRPVoogrpJPRM7OFlj5mZCrnmUD
Y7ReAkuOurc/33ggNroZKiN6oszqzy0e9FO/eZ753bMX1pnc+LItT4eWWOLADOac
mEat7o3sV6yWd91hlc5Uvi73iXaES0GINduQLEbAGAQviAZ34LPAxcGZGjGodrV6
jrH7Jj3kPnjPnRVMhCX+QYENKvjDpknCkyST/xr2ljxdF5Swp//wJi6DGH45D+3D
fV5yM3+tA1QvVXZsH9MOLZFAeDuXBGQMyq2YNmWtvguCnA85mo59y/tuwS/h6V4D
waCAlqR1TmuTPubIrTxN4COt7Y0HgZQkTeqTqiUSvh3jH1o5ulb/OpS3M81UMCgc
jYYalCxav0HQlK/Sa/u+XU/DmB5PX3DPK0qmcUP5L915Kgp/BMHC7GuMV+ww/+j9
ZeafKJaAQwItW/PQi/g13XgoeQ7ET58UXrFqqxXtAkvwzvHLDgOYe44pyNFp3jAe
IU7fL0P7+E/KbqRxQhRAc2KLICZrhxFDI/2yR8CtPEMfOxQAbLICZtqMybZ5pZSF
0iT3SnU6k+CNouKUVNODRJXw6tULU71FmJJNZElCuq6FCkxyh6nI8uHnG8ixqz+y
ckxyxGAEurIg2QUVKnF42JKjj8MNlmOz7saksO5+52XelWpxjeQi91fFV3iufN84
AZjVMI0gY+jTmgZ4nIdAsoNMWTne5KZIK3/y4xMnjUVTAEhWIgXwBXxqMK+sPbpw
TvYO5iZsIstvYvkDOJc12QG/6s/tHejC9CZ7lL3ekSljI08NBcXWtcO77OfZhujv
ZxfHFqAVxk6hzwYJW82db1Xf8keaSkkLFy/hqp5Tl3rWgOiRwmnGKnMhV41xMcQb
OF95W3sjdEwqOrf9ughyLbzWbpxKGeSv27gSmOgJ3gbcGlFBQMDhNTGlKJ7TrolG
DwysQyFsJz2/lpef65Xyh9dsbch1ZKUmJ2OYG6BTYbAyU+h0y2zFNzYy8D2M6uI6
3ksgja1U2m3Ds8HOQsB216U3lQuUAILyZmbbWrlVQyq3x/qqXqorXg9FjY52Msru
r7P84tZTh9DaDiQSQTjlSjYMuJwULh1bxIjE7hp5H7l3dQYeQT6o8uJyXGaXjDb9
s4+MHRIXXHjKNwERXXV8+ksQvW5dbGQchYsRPxJ3zpBfJwrIUNrOodk0gnMpiH4T
TahoaWpLggMfYt8z3D/lD0nsJ2FYkfv4rbdUXyjTmIMUNLGECmYsvtamzlDNjlYI
VJY5+ArhQ+f3SnDC3KnOGwzYaOAr380FHhqc2dZz6FdDiR9RqEAoSAO6QOF4rEgv
P6D1Go+NNZO6KlZXPTl1X6kDfQBe1efwY3pPSc7U8b5U/iSdXPDnIyAOsr3F5Hg+
xSCg8OVADO5j+CrQqg1JnYPOBUeZ7daTlGIed93WoIJyznF4AqKGUpmegFDbhXoU
mWXX0OKpdknwSf7rM0uEGtwxO/I0YNkKdOt9hA9qI1CAPkOh5jN5g4TFcM08hnA3
qk7l6yqAiVcHLJYVwOSb1SwHmssCiG/L3jwlQ8pDZQgBMOovlPRg7kZ2qrbmeNII
o7Ei+o7Z7TCnNg8NnS8TA0GobAMSO0tTHS0e+VyFaPrbowdwXEOhpu7yeQ4xdC1u
7yXRwcfl8Q2Q9QFeelWEscOILNZffNKY2VVGNaUAB3FPbwwGhShR1Ul1mkBhBGVD
82vYkv2SPABEuDcaGKMMK0lBrhcUwNcZ2f3Q5peMlwzsB/nFOCz5Q1lu6hebm6L4
WMdvmbCY0jg57U1oiVycqXQLaL4L5tXWUPjtounUUYL6fPX05j26uYpsD7m3iHyl
ivGRpRh4yZlUTjqNku83Fs2O7FmfODX+d0G6WzdSVy3gjZuFXq/uPe7pDIS7FAC/
mWh+tMPejcELrSD3slWw/TFV8pOCgvz3KI7Kbj7BYMCtRyW7Nz3hm2mT5IfMvliu
45/FNikk07uCIBUbyGjkErzD/X4ZIMloY0uo98aTYbC9JcLScnzf6iUc+7M1/+w9
4EToN+Cs3HDhM7ajTQw/4QaJYhgtcpUHI7x1XcJTf0YXCGkthrH3RmGgAUZ9AakG
+GcUKuPt5Kf2siIpzIbpDAnHzmH6rrF6A0YhyHfF9OXlCkiL3caxD0LcVMaGq2MA
Jv9fWTua2uV7G4RACelgGzAPeR9oxpWrMGHjxmTa+ozLOnvQb0CmWlm1CA4Kr3Pg
6cF4rITiqVEWyRyFUWQsog+43Iu92SBPlMd+ARil24YXLXKWjob1meD/lNtl7tah
xfBs/ivOi+vsa7n+8iikwIbdrDyM6ZdYNclE0+dy6gVnJvnuWW74yUlN7E7ZHqeS
KLHxWDUqTxl9npHW3j2wrmSrO7F1mPhZJtA3Sbush8XPG+0dOVPPJOhBrjKOg5kb
p+QgKOxXXkAJdHTVqo0OMRtqjz8tlyvw5Hbcp4D6+M0SkAjMw5H11kxI5VhuVJvF
dQYeUWNltX5Uj/ceNMnPWRDzAw7cFfht+SMBPyHlCdKZWLJYp0craLcWm8EYCxKv
orD3tp12/3UT8fAkDDI63/S9iEqkEV/HRHGxHviLeUsDHN4vJJUJvKW3Oy2vW47z
kpskCXHpNZfmaeYRRbacrcSfqPjOTxwje5TctnqY30ndTRhkyz7Qf7GvCTHz244Z
PEJ7JO9IVVygWrtAQkIuaDIiOPDEdBDCeWhwli+oTYkj8PmqSCIUOnc40SBc4qVQ
ASpnKPL7o3jzbpKuTFUG3XeXgWDYOO206PBAnQJZjYCVm6t+1qSrV3fDgFuW2QyV
vEQW5Su1RcefoWXsSGU4RHcF96GAL9e9AHLJfnuHwYOseyOKCn5VRUO5kMqcZ1wR
hp3Y99UiF+lXKA1uFQIGFFflv1wJlvX4ICmpqVzEkfAtRU1Afl587RvGfeeKGeOP
oAl+y3XgybvfmC3umqLbX5Ag4uLEIis6sCwN05yh5/95sRwPv3IE/siZPS8NMVDS
eflBO8zGWcN28tDTu4VAxmoY1sUpJSZ2T4pNlQcrPjRnN8C0E4++F/bcIEBPMC5N
kCU04hKuEV08jqrgngsFTGqnUDeNIrhWMTIdmQYL49hcQ7VpV1z0Y5tKFkJFqAF9
v5VpjQ0eXbEt/wAOnJfG4QW5jh77o3249irBzK7qnAwX6PBZ2KQacgMtXingA4m+
7leNmEtZnvUYPj6MUZNQOPjVNC5c5C6cAmAFLxkDdCoi2yViaJJojjw40RJm20AH
TKIRmn7dXTJenhG0DbBRnEXjTNhwuaiNS4XP4qPSHqgUAIBAKN5TifCaN4/bQuQx
MoYI5+EI/QFALrEJh59TuJ6KWryI/Q994BZgAuhpOMLGSXIlKrMKPfkNOrTMT1dH
sXt6cW5tCEQyQFnwymZUXmZ48rapDtDxeLfjkry+z1CPn01nBa5ARe00NOaSVTFM
RxHCU+M9vOvc0cFRnmDnGr8REdqTpUuuup/1Nr63PJ8L+VttEHm4zBZKyrBWBJPz
M8htEwYnWac3SwnFfpUOo8vZIH9vBUUWRmps7eP6CKkIV1S4XO3IhTMpt0BNv3ag
ldRuZVnnit6TifKktq5xAJRwaO64vW5pos07w5K7r1Yz6M36B8UTuOLHgR+9OCbN
7Q+/l14Sqg6DO6Bh0Zr9gylsKpHgPZMNbQAVu4uEzr7/Zqa0gr7AL571VUup4htl
f6IzLutHQSjck1B2KxjHGnPHPt8cU9Bd0Sgm/mZse2UqUZyP07eGbMKt/pdzNv0q
n5x9QGx789gVClJLWtYdEH/OXMHlySEwmk/rEMx9m1ujFLhKMkD1crCoWI8L1sMb
LwrMlLbJMYXMJSB4TxhAsTed5hlbUtuJkQKhe9kMR5El+ab2Ax7M0n4e1v9wOciS
6lPEiW7jZtz0Mp7f3mgb0u3hFUMZnH02+oG5OxNzBeCh9EaNRsxPrUiWdBa20fSH
Y5KWOIaBBYj1zGNUPESsIcWKJ/3QrFKgsBD1Rdq2fBXi3qKGDgxHPHVg9pSjEmRp
aVcvrUXk/HZIPVHq/7qr0rcY5aacNG4cIUY9wJbtTjBeREJeco8wXsHn7PebhEZR
THc076wHuC7iUNuFeHThQUMcllJHto2uyBXdXCZhiTp60eYbAIYEsJCOO1AhvutA
uudrM0xRyXDQQ+A07g5Ba00633A5qE2Px0ANfC0A+aS9uEKNiqXEnq0TvgYiJe9z
vEN097exW2xlem8YJV/By/kdkud1TsX6/RHnK6nzSb3bqSVh0uEfhS8wRUxfUTNr
c3E9Zr0UVWi/7q92kgQa7qn94vsFuo30EdORDlp9Gev+Vo1zwqFGZj/QyYIdVQ8w
MbPIAmu0Z1gs8DHSvMBU6klPqS7ghhc/AV0mYDA+nSgp2cW+EyJQqrgNxZI697/R
7kpn0pRGCLIqTyMQLPlhtYNgi1MlqIeltK5Xrao1+ijrZjla/eSFBiiPL5OQMMWD
DebKCX2br57HguzFFnCHSweLUdoTQ0iDl/NbUuwWTktSkv33jZn8ZEHwQA8GQu94
iDIRFVIHkcPy6ut/pb5lg6cdtJrC3sxbyDZnaAac7vql/7WrgjQ1ni9F+K/xqdRR
XdbhOpgajkLJ9pB+TTAS0uujRm88bpnmfCnPmt+rBvJNov51kA0mGVgS0zAOHvex
eIsH2cFMUZlJjv5WxKHVlYqI93FU0oXd6Cj4EPTraWrBzyzxo6iywNuN3CLz6erE
dDm8/tla0jzx1kuCPO+F3xTbWOCRuFY4ZigEUKgvFSPFyjyX3LI1CKA1rPOgmIKQ
sBDSP8nOvRgEgTcO0M70CNn5qO/s6frkmj0xo3pQEf09zGfFw1kejH3RzUkx9+Zj
aSHHCj1X3VH0NN7M0jBD0NHXi2JzHgBoQYc+WO0YCfuvA+oex++Scl4+vZ24GbiO
vkxKbR3jx6B4i9mJ9I7tIHVeBDXbGut41n80Xa6epjdi7GlGvAweOBSG/W6Q69p5
4aciNyz7+gzqx+fB3pZSkM3YrXBnuULlHiAS4MGQWKTH8QwvM+hVBtiyeCJDIWyh
QL5IzSJ3uSQHrnYOH1mi+8CCzNsR8Ul0ubq2CYpOFbEl2Q6F31caEpjCAYvoF70O
nYySGlWAwK170wfN0WxU9fE1P4kacyn8/cFF3VK2yizsotQmZYOSK5A8cYWKkHvz
xW7lRq3fTpTAUMPRQnMcgCVKL1gmGd4IVCsdnt5V6etGud7EAXlUDEmEztv35yt1
tWH1C5B3XoMFMDCtj/jbo92g7IPV9mc7S3uIU/tUR6+/2ssGRcvDh9JQB4d28Rnp
Y0W40jompvxFLQ2LtZBKWUfrEAbsxLqzGA/dZr/3RtJ6qFZNZTnJlb2uWovLeTg7
cOFXVDlphfzyqKAUco179QU7+YJFrBh1o4I/Wpn5QFbs2RYDYMD1A14SEJd50UUu
YQz2xrqskj57GXRb9cdb1u8q6QycMTkIfYMc10F947C6w8HcuLZ87vFoRvCe7KtY
dtKHU2VDgco9rh3jn0bfot2ZkZe4T4xT8aLUFrOVqktWhuqtRl7ckp0Y3scyYE4n
8C/IvAddqn7KVJdkbD1i/QYtTRW2xoxrCICSuLGXbDyJVkytw8C8hVZpAiyWI2mJ
LKk8fAyelcg3d/razhQmiGSrE/hGq5bFFzbZJ1WcBwfbvlS/Runlt0DeDEo334b9
Feop5GUkpGs7pvxJnPEJYud52r+TVlVmk988UcK2tGc9+nqIuKoWoNHR/T0ieUO9
OV5oM1UpdjE3DGSI5slxRT2Jjfi9/yD76R0uVRQ8++KQ4dqp8/DFmtWlugoLbzIC
Rx41rmDBmeIQnhd1Koy1kXMVRDQJKqD1ocBsqlxPcWnBrb2Gvkii9kPldtgIFtx0
sOsGD3q/YmpNVe2/YAvg6oJcaDlRAbiMeKAoe86provVK8hW1jrvhwUOOm7YX/ar
THR7XAubRPaI/nRfrqJfXiRm34FYem49BaH6cgJlfrO5+ChKI2VP82dtza/R671y
f0xymMseI6nT75I4nvtSjylxSVMWmqlrf36Hx8NS4fUzhaR+na4LXFLlKHhPIJjX
4EWH4SwxJc7P/qdcWuCIjV4E6EuzWrTG+2+iMEI1SuQwldO5qoVtnqtjB7TnjJyv
62RmegbfgHq9LOI1qp6u4w2qut65ZCc5CXR3PdXwhoo3AJ3uQEAxRvTR74/43rL+
UA1sj6nZB/pyAuz7kPEgabfywz2SwisA5PEk1fqir7Wox85Rv/UX45J5/5KXrYLV
GgsVmHApggugJdsS4xQAyrRIvfTBvGxE5N26Xo6VfC7yVCFTFDLjsyCCE7z8lS40
2KYIq52tNy11HGk8HkF0bb3ByglHnMExJ/4FuauaUTxWNu4zadRS0b1M4Vjtflv+
ndzjVpDJFd4vyQ0OyO0bk4Bx60F6Z7jo9o9+67pU+WWyKjI5K0z0Cq3Kdso6wIyG
eq/FsPuBLJT5y1o3CEcGSboTO7JIOPxWjivrCs6nROuPvGxndAtU2Rr7GH532VYn
/KZAHivRLEoGROW9DIAqnol2XXVlu4Thg/xbL2jKVAZ2DKhTSRcFNTBD1XDvCAK+
ca9V10NljyjbzdOxGVemPgOM3Ei7Ygl0DmESbeW8civDQknLORESzxoEyAgeGtsL
DTXuXDRvllCqx/+9H59Oi8FrebuFSznGsKOD8N/+93F8nlM/kCy7B9uFtIagiHtj
0u/HuHxBr4UBGEYVpk91F4Dhi+3nPq7nbzW3kgcsG2V8uZS+g7Hy1+qVRT7Sjwq2
mt3le/Fq8DyXmxGWDQQs/mVASX3XltNPjSPCkZ0UasGigNNhHnX3xdpCIwJ0XVyi
wVnpeQ/CotUp+XC4Y7Tidun4iANf/nmGRuDM4y4tv1WDKQWxJALZOwdTWtE0G5pw
Zn9C/869S4E6u9bWxUhChBVCwti8as3JAuRFpStGtgG8FNzYo2NfDgTSMXfIocCK
GiWqCNfECx4yuwaxmysPWhhEB14yezfp+EDx2PtlLQJKKgvkZuJ3uDJBHuqA0jJZ
qhuDMgRYugnXvCHcDns/QtBUv7FrEE9INKuYdQmAW9DAg8cqMoN8Up69hzhuGSRl
YHIS7/dfvR1sqzLg8bFXTgCzIeIh+lL14sgzfwnXFNPgDhmdgEP5PSHPaAClqKUU
gQuU9mojV+BDQ4AJO21ciU2TMOZnCoIb36MpLIy2C+Cw+WGcqOLEjHXnskbairBF
apebicmCoa1dCRyAGH3AWXiWRYwIrnq/Xa/n16nFa74nwI/YEhZG9A2MYp98v51F
wF8nxDKN/jqDkZsq9HUBCde6HiVrjtFQICwuAVdhXyZ22xdGGplLppmpXtt/uplV
X+1Ffg+757Ag60hhieqaSlrWcU0t9SP5F0LVmJxVyheJ4UPpta6JmtYtUkvLTLDJ
y5kNwg3HP/FM+cbaz0k5/GZACr3g7JI17E/Umcyftz56qMdyIKM5BEeJL1mrHdh/
ni2km10BwCD14r7yKm5ZVfBGQswkBV1Gl2DrrwpYWt6yONlbUKuug781K+OOi16V
kmfgyOo4kZKiujujkFDD+TQ2I5iqPC5D+hegUuUK5ZF6tWfeKCXVKQwuc7xSe4SX
E0EFVdeErh6iiW2Rx2C1BN8ptYJymQhQaCLJyTyK2AjsCVw2xa72K6joBajTsvW5
neI/3F/SjCB/l9oXseaj7mZpnDtu0/qNQ8KFWNrzcoIybSwWAmFWNx3SMW71nbxE
Vd58IDnIBhrqG7FYPh8qiHnPclspa9wLT0IZ+Ezq6hiKe1RZfNWcgqn0r7jgLLPy
s1WWPmkJywkHGxj/N1vb3J6AvYM4pIXTps3sC3mWk4X0oTukCM2okVCrDuGXjqdk
MJ3Pfp/K9rplXd6jGrGMUyLP8lWf0NGWonpNfdveq8e1T77vxTOnEUK/txXlxqJc
DosEoxaewmwfn4Z6TSdJAHuq/zWpxFTm3dcITrlJ49G04Ohz1ThR8UCIACy6P4Za
Iovu9PUBe5E9K/bbr9d7SQ5/dZ94Wi6pGOqt+xK2mKAh579kZUTVJHOxy7a9ka2t
ytdTOl24tVuO0G+Xtti6Yy6kMQHXu/JbZH+hPoYzbHVa23mcTJl/vf1amodZ9GpN
9YARaLa6W8jHxXYwphyTI2hpMPFR3EAvzLQdm15UDAaVvtoxOrvl2vGbMTOcs9hI
AZ9PP9CIJ4lkCznnz5SMUlaYLcMvo/pem1BUz22Vlc2SgEvDvptgwAewJ+YpD48Z
CHOmOjJPmSB17NmDfJf0xNYmU+yJkNa6gISHnC9zhhK0ilJcJF4XL1guMBYibW6r
M66Tx+Ltz7yGwMPTjXMPrCgCMmTgOSjIuPStqHAZVD1V8/nhfAz7o777J/MvRc9C
7ANDPWcNZ0yEI48tnk2ivnMQoGEZ15NsJy3OpmcR5IS+5QeWKm1ojqkKuoI4/AZa
iJjrSeTvRvDMqc6c84evFqojL8zqe3juNL2bbxWRS5ppT0GQADAyBmiv7mBHGz/x
c0+nXY4IWdwjqvr+s949+ioZutIohoW45tOnasqzBkRLLefP111PKc+4xGbfzreO
56waSelmFGG/x+TCJq7AWu0Sqjvd5z2YsjWCEbglATEhbKU+sxuwSAcYWh8P7ky5
Dv7aIB1N/LW1DBORwyZeAt5+Gso3qdWj4FX+jYQxSTqJXcJxluyL/N14b871eBM0
FCLArMhDtaeI7QswFJVjUicqeB6KUTWKy8Qgr/JYXVj6sWSMzBQ4j9ZGdHUC9JZJ
rtfDd1Vonn55DDZcth/Ne6mCpsieUSgOcMeuALnTJ3t25pFbsDEKkJWgCkA3qlcv
US9lcoATcgSEhnj9vTwokbeg+j32MyP4b/hQB8x7zLTRRiQlwM3D5VUg1dpHbV9U
f75nX5wxkD1QyAV67/E85oVReLK7Bgm6sPah83wCh/1t/f6byMIj+WIbtFYgR/wk
v0i5PVw/7CrTP5AlvZJBwI5YkfjuWFfAliHqMFqwnXvOIKxRGidvOFxhj1WlZtae
1fmvD/TTfIVQrk/EnNPFAZk8350WrpMHHqiCWv7LA9135tI54F/4aYD7rjya+icx
TwmYTuJVAllA+wqj6ZbWLs3bWyUuHjF/gMTcToBb5KOjbs9fmThAr4isHF20tn1K
RNtOIIhg0A3EjSCs6Z+MGXZ603s7GRLDAqPfj2kLfgkHmJkpwk9F7Z/6S/6mzv8e
IVKMrX1SQyX5R8EMP7JRqJmhxY2ZceSnMnSthE6Y0+kOISSGvGxXMwZJjO302Gip
HpYNFhR8KQggal7Co2UJoP0+2H12a5/l0M//jjxAJxnyg+dMGvjYa8wJhWC+67hg
QklDj/cMITEcZQwy3JASm8XPzWG+uAwoSDJqNT4Va3R5qJ1vBds/D7ZpHCp52KLG
fZUn5u8I0nOmpz65MLV/sFG0RKwUNYjkAzWX04QnZP894XfOrGXqiFvExlOiXhX+
6XChqTXLYtzV2GKDOCtXgd9JNpQe3MVYRhQwaFowyd+dJNNtKonuxv8ABPq2L77+
NSjbC0ECXj9fJgivYwO0QmFfRA24S5ABz7lMi/4o6Dn5b/MC+j++Nr36mEbkTRuN
nB3YW0aAt3S4oHzgk3dDTlKXRMvJ6tSMDyE4tzUSk+4XlLBFQTO6I8+oDDuu3uXd
yNdH+ln8ZDxnW+JksKCLsJbaZv99rseupmQp0gP4VT0Ke7tkqDQ7jd1l0I3sTCTe
LnOKryxTG4P2BoEASsJSSu0nBKTIzcAodNTYwNX6V5rMq2Bfpdx86/CbYen94tqr
fomhezEMFE0u9S9tdJ97oCR2N0lL+cBSgUSWWwyoht6wi3r92sBggrnsZpD8C48z
BF3sNt7vZGBcvKm43PKEyACB2B02YZilmBgOk9TejUN69cVE6AryomuDySXnoItY
kCWhx1+mzJU1PhVQxJmfM85UkmxjFH+2NU80IXWejveby1SLFS/F+boJPZYNl4cW
luN7WngUI2jnot12UIC0DPXAboVZJ13S+I5NqQz4+z/KZ5AqCnI9NgtEeuKMeSgJ
kuMHaMHLETFipCL8IrP6DcRH3h42kBLeXUwzdSYs2BOuYo0b4T0EN7QOjkr+bBSN
MWUhg7GKj/hTqlQoePirtFXwlN0cUADC5RVsScm5Oi2LtoIZSc1CA1XyimHmnNfY
4yEFq/a/mdbYt//JJyYsIV68SN5WHpJ5W2pfQxqDz8OcpvLhCq4T3Ql/L4X0DRAE
RrdlJZAXEwrDvOlEhf2F1094yEu2HSlbe3l6J46V8R0zkuU1Ke4CtFo1F+CmNqOd
aesPjqOJWdpL32VXb56WrECaE3rN7J/jgTrvembn0OSkCbIZtG7HKIsXITInCzMu
RmffofUZ/7jOStzD6Qo4FVIXQeaITQO1B84EUYAyuXWYB/gbM3AZ2bRVbJg+INYw
rvAtbCOJ1xrefQUMKbjMYm8uFf9mhi906V2gFSCQ/4OzvcXT3ujeSfSi1JfvjvNq
d0zGSRA8Ltgn1I+7NQJtRz5s/T8fhPkm136W1ZnvTHob52mPIBy8THAldYvxlPu8
+7EEU2d9OogOUfNABORV+JHoP7OPqETtSJUrmmXkTtKxElYBfAXLOdjMizlGA4e+
Ti28NaQbE6c4VhvOiLCt2xJ9gdeQCk43sqe0x07gqFZjyIt3IEk2lfJVI8y2xocu
AGuMfUV2LKxScp0seebQ4P0ODnHjE5NdkhbAcmevGN2KPpkLNQqjSiscP2+KZPJ9
cBOxFuSvXKZ/FL6T6mKRQzSKDo/ooVsNxLufNq60WDDZ7zl7WP0XffmAYlGbdDxE
LOG3tP8Oq9POBKnQn9C9i88dD9nLqsp6xnPjmVGD1zdDVltARhud4nAfQa1IYjny
2KqdLEBDassFe1bZ/+lYY2cSDEuEukLWkBs8IEFFC9wpBYuMUFGEb+5H/r12E9vR
nvcWHtiqhfhMQMrTr9uZxD6W0kb31ceT//USj+PG+Msa48Kq6NmZC8sdYkRV3E4j
0TPdY0SOorLvwhqk2IxCbts7IZypw2ozX4WfTv7AgQkOEjcK06yvWZTauHj3g2N/
FP8WO6qAfXhGJGqyFghoZaGLXhecVUXBZH6QBcqLiyIhJlPRvw8hKxHKKb1GsNXe
tKMjD6BRhfAXPIL9A6kHzZJgysHE36FTotAFrbDekYdZJVtImJcNVjy/MTrOSq4H
aHNx7bSGOzOGULXhzX86OHtfhRBSRTkBiMchhUS/Xo7GGwAJRYiGt1PxgMRojIqN
IuRB6CCVho+6VuldkZxTLtVP+O3khKd0w/qQ3c9oXFNEuNKPFoiF82zon+dsdk2v
T9cay4Vj5+dd8wESnJpc31U/rG15l8n1/M0DtTN5/p2uGjVksQK+qumizZBv8wug
IVO+qk2GUxkTW+C+41Qd1OJ6hAt8ycHevGbZlxLPyA0HfcGbxHDGL/ZVUCjcouPp
CKe15KG7INk2DbNKPOiK9hBj16M7YhsSRJmMSXa8XHxPM737b0lfg7bhq+/ht0GJ
AQWir2Y6m0nuQh0SO83gJvf2WIdUQN/N5WuxzeSvvPOFIGgM1xNUWjDh0WJ06mjv
H3SWo2T/QdJNkdKmAaP731tJXeKMBmi4MlHCBCW/d+hp679E4cMlKw4GWxzK4fUC
S/5xdexjTQ+fQsGda+SL2Z2G6V/3XKAhkUnf2RdDA+Ay436plxR72OfsuJ894r3j
C4peZsc8McbQHC68w2AJ6zx0lfN/zd3U5rbLwMnyNUpidwIAKTywjG43nRwxi2MP
D2n4p/YrKVSS3qLlH6O3EduiD+AQiWrlAnW1GKiNmKlTH4jdiEdLtdnYs4N+v0Xk
cF+Z1k3tFiGUQCpqrJAWJtAO1/j+AtZZTe/mWMBEOc1oEj/MUdjrpNnmGjxbkI71
qnZR894GEOHxiVUiHj7jTe5OMblVKtrGwWf4dbcZm89M3lp1ltIS/VoPIYP9P2Tf
r4Q1VbCYd81ETvMA6RfNoj3y9H2FZo5DndbTAqKh43Fa6Iq345QTuZcob+tqSVbo
Gu4aqCS10DrwsxlyTfG4deizTR9enD3P3mZW8T+gJKI9UYVIu+3nQpVzYjKqGCXy
TUC1GgY3uPw1R/crDQtDDp2u06aZo0LBFvexGfzs2nDA8S06xpGgJ6udAPSLR0Hf
nA8+YpafX7mRohyJUsDu/sfGA138Ev0lOQ+XGnvFBCfANszUZbKuc8eHgmCaTGM2
6eTIN7aEEtVq7tcUk5vlw+pYFVwx1rp6oybFRyCwgQqjU/UzSiVZ5RFYV/TcRCPc
+URfFYYHWZD+7WPnSkijIuf1LAYApwJYyNhMDJQg4jCI32/r8vMNJcutqTDt3p8/
hLpZ4VpO8SCNP4W5kiX7ve3/Ftld4CH9W54/QzUpPdjpt+Noel28GMPbt7ZJYJq+
L1bd15yQx3dVccc5H16FjHCJPH4Jw9PB0i4v5qSDeJEnLX7poHNPlHo3A900oVze
OdzFjpyQ/Ca3eIQPSatYov71MwDYRrfQb0kAroC2Kne2/Q3VoEctm7/q2M7lKNRN
hqJZ71FA6Pf3Qsc0jEURMq1ZTfQvOEG/0k4JmU0cG5iO8bUv67hVZbRQE3YeJzuC
mXVG3HGB16Ps+r0pmjG+sZY4Lu0/88fAzr8wTJVSnSxXECxApamZAHujeKIdqxtM
mjh9XxTdgN7/TrmI2OjmT6Yd2XZMzzKLvDHuB3Xdaq7E9I3BcwGSnGlmvbNvL/ls
DRRw25+kmCSaFkj2Xtndz3oJgkLyPd8INc5S1xo/pbXs1Ad7TLyDxBxcqe5u894g
6E17ubRw8r6N7LSooGNGsQMZjl8in/VmVFV2uLiBKQ/aoLB399vcOfVmBiD0ULh/
BKcnak+f9sykt6wGpoJhXsAWoNTXCshasKjftFE4qWefRSIvq9p4w9TFZt8JSse7
XPUlTq5H1Ou9FTG5av69zevg8fwJ9pMFrnzHKQ7iSwbW8W7YPy9XM2vAiD7gxmNT
4qkvPrC6RhpXJvkeor/qCv1J2FZZiREtwIV6hERX/m5qrhlldXYUrPB4pubyde76
Mnm9uvcGwiBvV8tVPbfedNilwI42GUuj+nk++o+3KZrQwkiLWFWhzyD2WdMz26pO
XxRZknKR6S7r3T7IOA6Qa5kbzG3rIVbRl121doM1AtoA+er+/ke7IVysIR7aIxgV
n41XWD9eVH9lE/glwsPnMTQeupT4ZQ2V2Qt+9Z2Akxs3aVG058WnofZfRKUa8Xb9
tN7BdiuvwZoyBx1MDVZLVyUvrGnRmSFfKmvJpYfwjsUz2D2IvBuCQ/B92jfRbPJ7
4pyYmmTIWPo0H6MWbYa7iUbj0+SSdKFgT7Rwree1l3vxBP/4bkst9qo5Bo5YXvXK
5v5kOf3bTVhZrEBaBGVY7bT8WV79Jm3G2JfhXHIoJUy72TjwhYhQOL3VuASIdROS
HxVLwTwu6Bc9stXb53EVG48jA8kHWRjxeP604y7y9ImTzeDXowByk3Do/Whm8S2G
QZN8HdHQlwallJmZNmeCw4Lds8ZPxyjs2tPvXLS8Y4mLXU9l5TC+6o/93yQVoZ3o
vbxd7gcHbWlb9Vs+uKTTLyK1JSorswjUPEcU4qBNGi58LjkLoZYwo0P/axUPOWk6
YByMalwOE77wKltBInyVEA3QhWhyywiFzUAWWOC+xOr70VyKnfChL9BvNWO0lygM
Xy8Wr/XrFgHCZhLUxKIkOMT9/eDVk7eCx4cu2w5mhcpym08OPvQC+gJtLGHeY+sq
AuJn1Gi5EkQogP/FG6p/jn7YCJQj10UGI/97sLmzvoVwztxhgCf69rBJYCkU0QzZ
2QYArW8U9PA0saeIAlRIsVDa5sO3jHtkixN6FeCXpMP4mcz5HxS2OIjYN3tE3BlJ
ksqIzbKKXN71a9IpvWS+QM1Oec29p16v4Pxe4nq9jtfmGUlP8NkKxYYAGJrDop+B
L3FLuH132HHrBRt1ATCzOW9kxxez6lFyqIIfOfRBcZ+Fazb83QXkSGaSlQYN3fnX
eLtn0qIlo8LAjrMq/Pdiq/sn/5PuJ8r7V2j+bbATTvsCa5mqSwa4NvzLxZoA/F/n
Qzx4mdkr0le0q7bWXJ3p+RRgJzRer9I9hFIDB2W7mdp3VTeU5DpwkeAgVS4k8NxA
wEXyekJ5KH7FnKKtzPU5masV/hYf3nkmPcye7SAo812+ealZoQBtboADfFFaIvhz
QjUGHMwJRitmMGBwiglXMpVwPJd2THMjlblZVeESr21EvUhGuqjw9mFtiwlbO9dn
FLXUNs9oTH1kmUsn4PbwE5ijiCz7YQTCRueLrYiv1WLs9PU1z7wxf4fWbV/UDdBA
Y0sIZ5LggAicdFPV6m3wid41oYKoZIzkmqCo+KRhpGK1j2AebNPsWe2lojTAO4xv
P+dVUsdGii4VBHNhM8HTZ3x7lVgmWVcDskoIiEYueVi6fwEzPhcdXjXFXM+YmG0K
LjbgFMugenJucgLFsK82qrVngOu8cJChGO9jzq+Z+V15gDQlEv8W8u49u1do9WKj
azlgi3oKTDLymEy3BYePxf+7UZXB6IkPIaSrYBAN4wQmRrnvRtwWB0v1Tk9lI+Br
11g4yaSku5ZBDfoPdxVfiC6Ejndq/u32/mHajTZ1tj3dD7Di5SQsifLICimjCnl2
iqNBZy9CorgweBeRAotbFFd8jJw0Vb1H/yE8H8jNrxO+wP78k8ZAJAzHLp6N6jtp
7EvjN2LWbgYoM+8tkpRtMRaF5VPSR1q4RwJ4VXCNpr7m/XOqareeK+1FwqFWMquy
WqahJJzMvGPE7nLT9CHgQk+efchg+6Yj8f05uBaZHpdsTI+e8HdKZIlWt/ypBBRp
+4DcQwrrxKUipDgP47SuVqNYOBhwIT5PHNsubL+O07VJs9vZPC+37xCQKSjXDz/C
gINc9g4YT6k4v3I+ASdB2WHja8/ipp95ye6gxF9utX5Z8SUpOeVJ8XjMwhGWbRuB
YhaJb1oVZyVc2y4SKjEnp0fCnb2WYCnxecGxjkxJUS1gH8ETlaZCiclX5GdfJ52d
Su5xw2kOG4DvwRQqpqEAZp2aJf/A8vslqfP7dAN6FB8Cn+T1H/snexMVJ1tT9RNG
fF2rFB89yYhDlRWnFKd6halsoIf3D3C0LpLyPsnJ4MwQfn/79tdYQtz7OMmKDy5k
HzUPX8VSAXUlKzYENf3McwwwQJX1yYybeaxGVUAId8JYs0L5LqVuYVkjJjuQogZB
FaL4cQ93pT+mj8nRRBuey6y4VIOf6MeoXNZSlllVy9vyArBC4oitbxri/KEz73l7
7tqTWiH6H4Cum9E3y3dhExoJCeqRdBISpEk9GO82dPaVgunDcF8bi1kgiKe/LLf1
aQolEJqZXBgNGzUXZGvuND9lqbjaqMWhLmJbha79KI4Ys4YYDVJq1UgqycdMQ7Nl
UP6xZmlc2mY2QJk2RdM3OQJUdQQypR6dwFBiI4bf3NK7uSjvMTL2dizoTGIhUVHc
mqLQM1/MC5AS7CJPmqTGXLOm/YnGCNIH11Nbq2xAxzxkxNmM2E1/4uy8hpoD38I4
zmSUUhlqrWX6ria83ASNIkGe0ZI2TuX48s3YZdR7xxN/zyTzL4MVDHEkUYjZQwS6
3mpC+HWPMR/sqswtoC1GmQDpCBGTH1UCafNwoWj4aKhrnRGJnBuoPg3DD0syT854
/hGThtCy59mmp1azIpdzhyXCFuyaZEEoXpcQujDakLOqCOKUYBvXMXCi4VRc4FbJ
8LBl37FwRkC/b0FlmdVC06EtXluWtk11iooXalZ8NAEzZzpScawEojJuDg+du7ch
Le+9GYD/swBi6gCsyjeCSkSFW0CF3hagjxDVLHJ21QA0CJsV/L8ZZxO8gBpd9J2p
BTBqfLsMPaONOiMi05+/ZdbquzoKOyWeGG6qUzRBTIq32+hLot4rZ3KSjbR8iAUy
/w47HjGAZunPFfKmnjKQJdu6PkWGUi0H0qwFRRpowXWyAgRwxgE+pOMC1CbXw8gL
SIKv9mqsDgvNiuLGopbL/6njM1vBiOYKjXriMPQ/p7XYZH8kxdENxzwD522bn72C
LvBxcnvZwUPB3T5MzzyA16e71LsgO5vtatdr0csquHb6hrlVNamuE7hWpNpe0ITv
exwGHXazeGVZ53IjREDtp6i+X4bn48wg06IWLTKiaXsKOLy4rbisAnSmRSAbyb9f
pKQBgQiwow5E5WQZ2Hi0mEbPx2ZYz0YF5XmfWO2V3/DxWWdY3b0Dctmj/sww6unh
iRTeTSntc7tnPJHeZYmuKpMS4PJIO4BpPatFxigEeR4zYoZj75PKu/ljan0T6osS
GJuAPz73wlUweVoMIVCSNKiIvW8dFbsmNGYMTte+cvpXx5DmuFw1oIr7dzLfkgnd
pseIGVl980z512V3vf7Yqo5f3pA9rz+k4aLZWNGUItahXJaOORfNGCVYOc86M62R
eSagGVHAl/Y7qQJTOOUtXtQNOA4ALicTnCjmOxJmhhTLvAy1zi8eTG2SeRw2CFSr
HPeBj2hiJdO5d1bxfPZqjtUWip9HAEl7lmf8B1ZmN99s345ssO60/ZYZcsJ6L+OK
K5IVaAYDIIDjHocP6NnVobwGDCzsJyhuHRdjN67PsEEX7jIQKn5R10quF3SeJVdF
4lxN5SrL2ijFKupkvaMoFgCVjc6wPoITqWe74+X6/WR7UTekeO0XcGfRf1vDHUol
oKQIBMpopnxpkS2Ud4ZXADSPiG8uPqOCSskuf08yRAacKDzDTajfAlv2syFkA+ZM
NtLOMc48hXCXN4KrAtRuROiH/w3OQPJ41cWpjYNT9YHYf2oxstnFkbutF1vWl23W
oza3MNFV81gzO34jTuDUQmK8QnmbU+hGdd6khw5nNfFvZq7+EZGNZsza2UNzzXfH
Zzo4dCkf2/kme37QgxS+4TQSzh5qQDrTeO3vGClLw2sWi7fLcW6yjfr/MkejDzgc
wVGc5V5x4rgH+9KohADjFPhJTX/P1iiYiIdecz0As0zkJZ2LNv1sXyR8uKc9y0qX
pfZay0UqQrSzby3HOlGzI1btug64Dc2FOwut4unDWAqQLo3Dpq4vm1s4ovjXt2Ww
1n9F0MSkjZk+z+/sddPOephGVNgC71GtmzLWoMOLDNhvP5sxEwyGkXN7jGZ0iO/P
uaHbktyaH+ZIDp1c2B+8+DZFpdOM4xCuhVAjHtNHbeUKGihzYKAjxajI1By5hXAj
WJ0tGLoZNpuxyQffvycfwltYZVYYRptoV+92kUsBV0FVI8W/Yme8bOo+looDLaz8
ultxX+Iw9B2VUP5r0gXrtncfg14c+lWxkFvRg/4K496Hs/ldJ09A9QU+uDlY8LrT
IEeXeMz1hBuJgT6pJHfOTi2f+BxFezkFwLou7+4rx6jO+pnKSfYcxJf8n0778mkd
I50BAJOJKnyqhCaceVZR++kHLncT+bNdO+Oi2PT6HxR4M+PN2yQGQErkFE84PyqL
AOlzsZ2PPpK6avYf5MR94BviEkYtoYkTIPb/lzii7WVAsToqIV/N8z/y8hCtJ0BE
eddoQYsehA60k4ER7E/IinOHAqH0XlK2SOWb2sEfxELyZMLCd8QxcjlXyUaR2mPU
3Oup/VgODkvWD06fDvqboRBuUQc95AMGS+LhT0tlQvuRChe6RZvlX9B4Y5b9NaBu
7rhrE/ARWCJfKeBixGX4I81uQVAf38mXZdXeghZ3rkCzaNd+pQ7IRI7oQ353MB2i
4E1IUcQVlAW+v0xZ+RdUKwk05oltC/lAcVIQGvzBsDJJL/HFUhbogX/zNn+PG+TV
6wKIV8IFXUsBZBzrP41WjjM8Ezymdd7xIEwjuuUPyR7C+sutFpldBfLD5ti7As7s
W7rXPd8UlelGgailkpCsonpILhbtoJvxrGDJ2HPA5/dvXiL6u0OLvEP5ePEl9dIt
TDakvL8tITJeIu7NtmxAlAdsQMFNRLvilkBl1EUCTnBUnm+m35FOSvt+WYK4POcq
Rlr7IdsLM9qn+PdsC6/1CubwUbHeHiLLPR2DAjsRRI5ZqPWXkwwXyErOH/VAbSEU
5qSFPPEiFw2W7grWXZWPQ2Q4zAPkD6aYnvxHoUyICSB78MSrlGn6zA83NK0/vKmj
VNywtRcfLVen6/xqYc0Go3vZP6HvHkAv1Lj8CSc8xSgczb9Wiu63ZdVbVm7fjad+
2tf7fZFrEIzH3FOj6ix5ATV6Rai1v0HsE5Upma3H8sU/NuSewrlfc/+bsX1Xcx9i
4DrV6kRkkebpo+i+0pDrcQb4hbkJjXcaWuqs3NXJ+CiVrCaCBejqaroPURRFCmUB
rIw5uS9Ae9jojnvq6j7BwRHpSPGI17VreNnw+vdnxsHminPDb7LUwCwOQ9cxy2cf
HFXbxhM36ydnl3RkMG7dW+z+x9BSq/e6Yrz+JVaNErdcGMc/1BJEaRq7Bl0UApBC
uiybFhpOk9k5xpaNudpV7tOWo+AK1/IUmPeqzf5wWyTaEJvL6x1HS787uGp9l1nw
M29PfcLdnPtbK6Y3EeklKYlv6+9eYNzukdLsp8bdaxqzXAf8OcU9fUTBga+3hb6r
lCM1LVhGFBtU3AATcoU1OglV+mM9aMGlpTvpULZB6Jj2FO+HkxAS4BGCK4M7vooK
1+yZQXgWLCPCocP6IpfJepkpXN71UahC2FADF6VaU1G3vdy/VtWoguzWmgJd8mIy
4Xpv3HSMPHeyQ4T8N7dmui54DqdkZB8m1EgNhmiSSqY7jYhWdP6Lo8rgELRWdg2N
z7LKZqtFl0O3bbnMLco5qd3znVD/EOwmolqu9kSthHVQkAjGmlnD5Ju404slHFWR
yVuFuVKNHiNfxq2YXqg2zaFkg5G07ReyekFEla8a/+aKXt4RJjcf4AD3vFgx8mPE
dYKst24oqW2M5uzqw+lw6xwK0HTmjz2Mwkx49HF2SUl7agdUPNI2Fp1rrZkZZzTU
GJyBJRqx0VgW/OkT/cWYHjmuU09el8M6WLR6mNp4eSBsPBRTvaOCRgZD+r8F2UiX
kea2oGmSNoT7vM1ZKc3hW/1YzlSnO6NJ0xPNPNKM7sESMfIGrSMWkdRq0qj1dDRf
zdGWgEjy8Pyr0HDZFFReKgbPLpjNc5MJFo3aMRuU/w3t5hdOckPItTsBcOvG9GU9
0DhCKGODMmWe5pT60JxWOVomidDSQFEwqGN9DEkPOPnOBQaa7ZnDsMY3qEG8LGa3
I0C5SA5rsiKTLObDmiNOb++YAzrt8xPg6BQZNY2Zfo569fhXwmNOWKMGwLlI23Ee
jPbE1UM1a8rLrmWBHKsul0DVyXX1my0Pv6382H+UMeQxfywlmyOM2hp/3NbLz2EB
qT92SjcT7SbKRkVk2HybjI2Xi8QdHy6ZJJgwQ9YLRyQLjJimwrOJ6dIPBfB+EfSb
ZpeY9jLiqy+XnE4hy05aRnQ+cYitvwI0smOYmqf5HDhtmta3Yb4N84Hu8/UdsXiT
lnULOjSaS/g0zQHpvkU05RHPHYkCnWwBpRTMvOFGPdq0rFFi5HJbKPHdZjsMG8g5
rNwQWxXin3GshPBWpouKeA5zWnY9/SelBLf8EaOszL/xQ/oKO0XflTFoa2Zi2LZf
xTR8cm6HoTSRmLTmSjNlq6E3pr4iOfqvkWPCAUDwjXxBu5PTWQOMoQInI1egdOw2
2+MInSu+ml03VJhIiR//IjPYJ1rx/UKDlVhaIe1GmNhRT7ef3zYOFLy4EhtYD9+n
N2/3Ze1DV1rI2QYkJNoHhY9QTdsvzJ2sLgp2xAo32qGwhzdlcwJxzqz/jb9JIark
u40nezZEx7dYqFI6/5HAB8Hbow83fRp8rAsmzfF0klSpbHZOd1qpmHyGFC2Y6Cuo
94jIISnXTlbg+54m//fIu/EYbzLzhyRkhWX/WWNpJo5YTyuFj1Jf5I8TnzrKmD47
XdroLKcwSiTn6foNFJFx2/h54BFOEDnMwQ5T+fSbKD09DxAZANfWEBCf6U1HYxxq
LjJzeSZB7RHkvPtjL5dGzpk6X2tDShvIMb3UosXOH8YW+/mObf/IrYBwoiIbqDwd
7Pl+eAL/633BHGY3+kEQTEs9IeHSc28MEpmrRLQQ/C58+zczFXpj7Kxcq+Qx9fcq
L+xjpb0UsKsTGMFxb6kWvNIzT01CZ6SpM4fPyq4G1boYfsgRODqVCdtGkmRzAmR4
apvHrjGj68A9kuZ3trq9BrooBCuTvWw9d0keAOv8sXxJyx+5rUEhWGmkV3uw5VCx
JSS7MNSkH3WjeJFGvCnezehWsWyM6529bICCejJMUPVP0Mr+u4rBfl1hFeJGEjnR
b+cInWAbY8uy212GC4r67tcxnyKqnF4H6Y3TggS1kxrad1eIkfj5WTfPuNdf8s5S
hXaoXBZKWeoRBRslYfo0PMHga7hey3p7dKxBQTZVTcdFj5fR6edRVWfwKccdYHjB
c7Txlpm5I3XkOQJgnZPfuYVBKJz3UpeJRkXJPxEpezQav50lv3UeQ85XXcxeKOcI
AAQI/QU0ftUETJkPjE8dxY8w1HCpMqlHAUcsp/+bD3oQqY0xkew5U4v6piXYYosn
MiNrcrf2Icny8B3pD3k4KWuWUF5gDgnLMVvSu5YA4Rn7kOecDPWFqx7NBO5C2yQ6
EclZymgkZ3g3b1GzAsen+EXaMHuoiGxd/mD2Z/58RVn1j5qC8UI2mMTnONj8go59
YLcNRwpY8Dz/J6BlfNmWqhLbh+2ZrEw/gRXL1STEBy9FEQHuHxIY2fh7b9pMCMBA
DGeMufLS3UqzONJ4/GhMynHmPkgap9L2pUSbIW5sA5CDD8c7ckwxr55cUBr8HpkS
AshSuwx78YbEFqXx5jMEFUd3TU1TjThy/kNYiXWCriHJZ6eXUy5bYPF0cyvREvnk
OftmA4zxMe2lJLFWl9sAVhrhoGSq5pNTe6fJ1lHmLOMTUvVcDNS6hbVgrXydkAPB
a6yk+79vyrNJbvCaELCCiKGgPGRAQcA/lJO0BK+i1RoleQIzNCHpU9mO9NhkWmw+
ozqcoUZO06R7o4iQJacKwBBZNxgc+hyjkB6ccxUl1TRgftGeeLZxLJGJxsdzDumM
Jxb5vLmUJjOan8fPfaQDvNfv72bpEn4ZIGDj8liDBp1kYLundyTeqvp0cq6BNaLa
1/yqOegIvtTbdICPPk4uHsJrZMpsBJCPpAviztmtHMLvkOA141mUwpawT+LiA2/R
d6GzEZ3F+znkJp9onIi4YsnDI7Z8py4mZ3jQD678UQCq9JFDkRbFx7p8R0B6iOIf
0m6DK/3AG4VIRNDnlwwPvSbSjcxb60q28W7KbMHPmvcrIbcR838b6ap4As1+M5Mg
RomEnK1fYINmm4YBoj7QDrd0dfiAhzAoYmWXZmiKxkkznxfRIKSe0BnHqWDtes71
Om4Sn/VrFIY/zw4IeousFJKNq8+4UqY72PzSQSI1Uye9lz92hyiBWerOoYcBRzYL
dhAJd0VQhgY9L4eu83R5peOiYaNI7eR8VyNrJrtIJgdlBTRzKDQbT8nBt8/i/ySK
GN2PPddL7jjFhmgkjjIE0H3edv3eLwVO8TXIMzr/jvlgNMqYn4424H5tTm0mRQIv
0RjoQwW5t0VKq8XUdT7IcGytx5oEyFw+USxKLrDQ1Gv7J0IbM5SYs3BzVSv7oIkF
4GRPzjpzPyvsdCD+TfVTCvYpKsT0+uiy8GE15ZXMfEUmG6BGC2Hy7P5h5oNIiSkn
sIiYIRZDi+QwZTLmU0tkkH2Cz37orv+2uY/5pwYWCXm9YuyXDH3pgPc4TBzoLxGC
qMQ5froyd11BcbQuW9//cJFzjWSWcsmw+8s91stbqk0MuCOpwO9FkdLL9D2rN3oO
X6dMrquMN2uMu16eMxSN29WXBIi5X/MDauokc4FVLQOzjBt9zk5ykH2Souf2A3iQ
nW6i11fwRGFu0yTtLF1ZvAy5C4M+zCPGlAuLSX1nqA7/YR5jNisXK5ChY69bM9al
XDG7YcCAO2YLFFwNfxVoPUd384nFNBHwrq6kh6yEZhmFyYfBLne3qtYapF3hgiuI
vNr97yIzdhUjaQ/Xiso/XNh/XFfNSeUR3Oy9978KUDgwsoCxQTWVisAvIdaDEkjo
C1hCTa9AjaadUtUIu3Fdm9ew+b5dHYBObGbwZZc1tfGpnk6mYaFlc4wTLC3FlD01
/Y+E0sPEOriYifTHnqQNyU2YtK0ftS5LahsxheRYhVYQJR1eHuKRINpUTIa7KsMc
4Cj2dbOHkkLAbdkcW49pDJEbRxUbWWcvh7fSSdGO9OnoXh5n22DrDoMXilsabLx2
0XefTeZJ+GRu1UxXVCMNB39Ce8Ddxa3UvOCGEp0jTakZvMBkR+toaLuQarSSv09m
ysiZHTn/EpaLJX5mekCbyVWiiZGL+UzPelLvg0MiRVPXfR0SvfXwXdRS2Bl13TF0
KjDsEE7uy1120hu+aN/TUJGi0hh1ymTFUp3Q7o8vappiLgGAZnJgxBAT90ezOtVb
cfKip1Dhs0dKyhPDmoX56aChHBG10Lp+zLw55H+vkYMnq3GphBgQRUFrguEqbi+T
hnzoEIMgzHb+/hZO5IIYqM5E4i5Rhz0Wg2wB/fFSbOB0mPyAwe09dCTLevmceSnN
OU7MXNp80U6Ma7A69WLu677Xjs2kaOdrtnKCAA/Apctx1rXYcYaxFhjlYCtKm/wQ
yfrE6+sJ0Ljiyo7yP2Fnd3jJ5qTerAndVnI5ZvlxNvcW5OCY8kGrQhdvPKlWGKq2
tgQF7iE10a0PP1naKq+kX1OEO97Wya7p/k3t3ftrbeKwvo1EIwz5wMYrTIEC6kNT
5LK18QzL+7crKWh2hmxcJ3ig4hV//0eXiJfQ2wM15xd9URpW6ohEHHNoP73FA776
SBQsVfpz4XIozlc2y0l9y7KqdMpuWQo5jyT8savb9fKDhj7x6Alt5Vw6DCrrX7t/
vo7e1SD+DU1LjS8JNYXRjAjKPJb+UHpcakB/4m6X+hGortdadG+hfx2+F/iftDj7
AlAXgeo+c9cey0lgyeP6m1eKp37OjlcY/l0du2nDI2KEnmHP0r2cTotBuQBO4pLJ
iID98vsKSevDZO1P479p+8T+7j2a3ldX0iWW45kDT0qvsUMtt3ernThilo8Em62Q
5hPRdkhx5yjtDOEKd7xv0bcwNgGIfwsOZA5gZ7ahoFLzDm1wTZ9xEPnDxWN9RO8R
fnCu9tzv3FRok7biAT5yp0eQ8KyLFRnSu9lywTpem7IDAxD8EwZxASe/6ur+xWBM
50fPeneSRQ/NRUiZFDLrMcalTjjJAK0/0QB38tsfbMhdKSmUEBoh6lDZY+Mm+312
qqfsoURGzPVQRv7LWzifjuN+7pyH00RqEmrV9lKE4riX6f6jCiw9V1cQemAf97iZ
XEZ/q5lomsXp9pawu5RO1JlD2oLMkkpFhU/ZnR3RgWX0qTMxdozsf6s7tQWlg2Bh
By5UH5Oc9ptd9LSYmkifc6h+gYV20TGSeI55skfs5oTe6IaXO0k2oskobu6D0i+8
4O+YMfv/z5Cz3YMd5suRoiRYS/sDMoMyFa8moJWrz/lDHgYzCX8gld4yj40Xbceq
YwgcPBSI50MIxU3IYlxXFA0bfcooHMC8/SePyJYTgLjv+7Tn69IPezmIPABWoP3h
Hy4cm+zTODRmrgNxsLxJA5kLZSfaobOpiMOJvcfDjxHlQKmZ6ZEUuM4Uo7JZfarf
9X3XFEgTsWtDl0MumD8IQ/gxSFNrENjjcSBExEcE01g2AwhACrui8iyV6q+cYadH
JUSiyv1vSvyIh/ZmA530Phn9PqSnjlwu+vtLi3su8Eu0jzS16q8C+EjgTQKek3Dk
s8ekD3HhBnagE5GdjFuQ+bo0ewmJ96zKBr/8PGvMmJdqRCHavZQWHlOXz1IojgsV
DnUJqHk/9dzQx6YY+FPTH/6Li9AVe3qgF2KnsQChx8/kmCQIRecmsdPJzGKAmaRA
JumnVYIQwXAgYQ5Uj0yTNeXcTqXrzX7zFmshjaXKFfDENtFJZj4OWKcM0fhfrS3u
0Ukwn5z6zZlbXcc+4jrQe+boBi5OfM1A0rFYZV2EbTTa+316qaThRvcxKtzP3P/9
DOQTSJcmrcVaKO142elL1Ux+69IlYVVRhHvOLEe6S183dZrVzHFY0J06QRr7sUtk
ERYWtiGMNw8PGYJ779ZqWM+3oehC2WgMX2rQv4nBAk2XPqsfE8iHQ3F/MHLyTVhL
08eZaX7jnrVyPKRDrWtOSicqk0RrLUdDftJnvWaUlx6PuHFL/eqrbbyW8zmd++jS
BDZmDSnZ+lyTa8OFploVgOaJe4RDYlbdkYdBC9cxJ3Iowvh/BlYKhaE9AYdffCf+
M9tOcDs3lOrC29t8zq2Cl0JuOUmWI9auApQb4EN4N1u2KBFa6aojfbQzVAeFS0ux
R77FlpO1nOXgbusCHV51gJHMsvBe31aTH0qFivkk5CGUAuG3PNx9oQNual0ThBvt
Vb13Aw+zXJrQ8wsYPm2tvIXk7v2KsBKMeaxmKG4Z0PwwBhqGy4GaiWlUQcjw2QF2
mLBFxwaqBBVu2B5nCMAiScptSWY93pGznA9zymzEkA0mDzQlvjJWJtw5ppQEvsHn
98/O/wSKDxjrVrqkt/rdF1b0KyszylEGda7OdI2W/yoxMG+ri6x+Orz7q8rwKzwA
bnejJ78bfu8JXQd3XjZalRjgaz2pYncyaS2taZTUtf3mmOLCNGu6V7gMW1OvdtgI
PnMWHYuW8FrkelOXX4eULx1RsXI6g/Pd4+rMCH3ymmc65IfVyvPwtQhXur7z9OkT
darsBEqi0QCaxRxdx5xldegZMQU9An+O3mXNin1IsZsJQgWcJKuUlM7j49jdPmbB
SQWwvrKcFoHJ5yPQcu18D8RS/myxwCSyGTk3hZRpg9OQHuzmLLzyBIt4JLq88i2S
cCkH0X4nqcTF2rzO3X68r4MYerDchm7ETTd5nN7Btcz52rM7n17kKYMUvR2kmaLO
omvuWWJbvuvzLsLEEh0yzkE/zoJEEzvx7edDRNPxuaqPWfpkrZsmeOf9qRouanMm
6OSit8HlHmDcc+H3A1o8ytrGPbuSlXVHbTM3FcMkmUahW8nhBL1YdZmm24MSziWt
mkC0tinzrxOMo276zcoNVE4m4QBZkkZLqaE+C50uiu8qxDjD0V8dNEmPkCWWt2zz
wqHgkUk+tPu20jEmyUNL1q4SJluGaTuV2c0VQDJV2aDAK9gOJ+l7LRUjGKBeEtIY
SsnPwS9vzPv2rOU69yqQXWxC714nCtmS0esYH9BfbTHBSEu3fKrfRJKMDyDpbwCB
lftICX/SgNbndNevP9bmj3L2TZmFpVSsOt7S8KAkjs2azhhW/ccy443RwPUf+1XI
zPHE3uWpfw7XRcxNjEVoHuZl0BqYb+qHc2in1h6moqyy/qeUCEVqITXUKs2ZrgQ9
7DbWFIVPjX6kcw0VtsB/PKpVquXvucX6khaCdu3Io+u+OxY5yRliLSpD1ATjzcQl
s0Nvl/xSrG8+yuDcJXLv3x40PrHPZ1cTz1qPuW/kwJ9a5xST0mu6laA3uoCQ+Jeq
+5WU0fS2LIyaZPaugEbZ+ROOrnk2B07Dbl/A6BFivQae+vDj3aLroqdSe2Axy+Xq
x61z8g4FdJxAj4MYH3YESgz4psR1NdyXHDXeGYbGnXIN3v9asQJnJgkN98NuQPN0
QFQ6iQxwddFA9TsHpFYbE7FtFyWb76xbrGxUS/DtJKhzQ1OuUU0Fji38L9YMMfdu
yKNptP9RDu998Rs79oA/t8sCfbc+L2evIjijMBq0IuP2MYE01iareehYuoRNv5yP
oMuqkV6B9ev0iX5PwXNP29J1G2S/FrlCOkPTi/iVcW8KnX9UXllwNrbDzkO0LqUY
1kfvyFL0mzuraclczUybwkIlN+ogl9zIgycUcJQDEp/6HQC6M2h7Uu0/kU0+0N+K
IH/SLeHvUU2vqqLZlYo6xYVZ0l1ehPlAAh4p6KA9HD3sosOHLozw84XXMNEPX/6R
8frv/Bie841yY9Skp/1n2NAE/zoBtnqXG5qTv4lq/FRDNGpkVUBR+c5Kq6QOJxi7
F6tkDV2b3o3vB1wE4a4OPHxLw6uqoVTBNf3/AyCj9LI3VDSeR4tRgXwu7IwWsiF6
zFyjHjVxitMoklCsokjQA+BcVZhVycl1O+PxjSPpyaGb1FtM8VgdeozNaENAoPxa
Otnzc00cYz/PUY8Abyb+vW+VSSiFPEbPHOzisz6N8rknGjnwXk/xMZOtmT6on+MC
/UCeOkUI+0AIVcoFEhD4ZfGKlX8KPPesDzPibCJeLQKKUmjDDnB+ctY1aVgJDZBM
yOSiJ5BPQHV57poLVgpZ6ZUyzNlCipIVP5Z3SkHYisbxCXMob03aSFOHVAGVlGMI
3/AqKtCLnouFXL7Tne7jukPfpVz3L4Z131jtS+elkzOkDCuWd+lWGjMpr60C1mvu
iGDx+354LKwLs0UNvmyFmkCkPHesy20j8zzXN40diH4kLi3FCpXuWvUsO5Heo9No
sONLcITD82VoIy5Lto4RH/8nX9CAIhHpzbMDkAiI6jIsaLt/hZXdqJoP8aDLprHi
PIzXU831cUUposr7Jadz+PjJzD/ATkml9u09HZ72wLpPoAxAzhUed0BjRMThlSSb
11PXRbCTOob2bXRwqvwup+FlfOe7PeELnZaOBLvzGfiljHXWiHMejBPTl+58CP41
k9ieB2svd/BR/HBRX85vd6QD/i2Wdq1l0hKCp3+IjKPeU1PjCNQDyqwsNSLZ1SR4
q4bsnpv5MxM0NHucuQRjt0rWq2LAmXkmTkrI6kAEsWF6eT0VS4SylJOUY7PVRO2f
6Kq6kEJvBJY08naThYHAh2lNdWvYuLrQYrGI3zxtJ72JOm8MmSSXNWY2UrBBTNkD
Dw0OnkYFw4JDke4wnJAIyNWrmRwona0+Ys9lLyzHcXY4eT3SVU8oq5BbLcLr2hAb
kTCvGL/ITHTog5lagNJBckg1orZtEwFfezMS78JayLgrMyU4xo3DUsq5wWT6jCjS
4WgzSmyZdSoaUQx3l+NVq/hucc7O9HdUPc0eM5/825x6uESqLYL9/GwMic200ukL
6eYhMUQa5cpyMFnK0pMKtoujIX032mQWFnmh4TNBvuzHz9bAqexeyYrcP1sP9YJN
T/xCznvknzgpNiDAe0hqeB2tAJjQ9z7UDwEqG7QPVO9WaGLsJ2o+eqX2B4fqvwWh
RUo0/lB5IYeGq9oVI0J35sIHkAxbN9nAMJACM4Pc7m/UBgG58aYYRngHDQYkRz2m
m6oDPO/74g22GK+MAtaqtixHL32nWjn+NqvhKOld2y9vxqOP+PEMG5rxnA7Zr5xY
bOUI6WW8qeIdTXSKX6SHoMoJFV9FyPelniV0v7sPbaQlwqE95L8DRV9M/MQjxa4f
NWuo3NKY+vz87C//EJNlUrPgwz6EBL0NOj2GL3Ud+Qiss3PO8C+l+/Sar3wRoWou
DfpKa/QMsT+O/0lQbDKXT7yjhuFQePlNZBRzf/BrpqDVJb5Fq2EFBl4OG6GjDmU2
wFWgTCBdZnBTzeVkA2Da93XtsjvCQy70vn4Hbjij5UMhYogq7CkjtEIv12Wop1aH
V19pF55rXXYCq3I8SDIN7I8muvkw1Hbqwb6O52OA8FQkUzeEZPhl0Cd0Xj3bkHmp
w+NjgdprrqKuqDw9LyA+5PzaNzervro6CEVsny0omvevhXqz3xI42ceQu7/bvsbi
zR/hXxJxbU7ymAETudDmDLSeAFwr3AmCna5DO39PYXiPJtx3s1om5/jxi17qI+y1
2F30IDtNECohb8r391G/wDIhWzWg1qG9LMNG/rXVcVYfi/6UwHNKbQoonbAtm+xm
XscK2k+WKcelcV0OupmF6ScIuAwHsNOYKPdglsBpfmIF2Futp90fN31fD3Hq6aVH
BZYFNWaTp4HJNzNnWPoftvzriXrzVQ3szEhNM17sde4AGCYls/Zv21MGpXGalgRj
GvR+yFXJX8UyG/WcqW8cBefuwzY9jO1gOzPf7SDxCya0iKaf3yhwaHcetXZjEDWH
rhfYfiP+fiMT7ti8/MUcvfh17mpVS+16jEzRUk9YXsW06On9gncvBkZyq0Bc2BM0
wsQlRvcHEQqkWGKEtdKeQRiDK77sRFTEcPvwxdecSAoywwT82tcB8KsmSXvqZEvv
8neo8ci4DMoXktrauGn+5Zzd+N6NrmpmqKXW2S8m/ik5xpcTcn2H2pWAsVHWe0qe
ah6k3E9farsQ2WJzoett9Nsyjgxi7kTsPbJDiwAk+NHQQ2P+PHAa7Qj68U0J9PSS
/aOsSwU60V1IhSBeLeflt+Sx6OEaHXGcHbLItZ56It65TXYoQEVNDdEpRklmUuII
2ya9mVpaSH2ZHt4wmFBl63gHbkZp2q/x9M+OsTk/DR1bDrb8mI4G3X5t+Ztf98qY
oc3yPKib7ObZaV51j7xPRaaB0df1LA17SmL0IP0vGumRrXpq+yofmogZ/B3bQvUN
+ASL7PYw9zUqeDVAuyj+wofY9kALgzqEOo0FbzWlslvcBIP/xF8f5ivIaHI+X0fE
QCXoQsQNZMRLZjXxRNHzrSy4AjHf8/SFp3uKsJIumkvwqiuCO1I/XjGbwgTJtmYZ
DlI62vXD+MXA67pBqZlWCzsovdHDsXVmGCxdzYbw6ng8KElQvZ9E0Qpug+Ois7g6
DfLSt4RD12poaATjOrQJxB39L5hZOPQUl/ViIWcJe6mcYa85XeD7wnxZ6qW/1veO
lrg5VUEwCrG6lzUG9ImOPTIczqtx9P/kk+0tk4JXjZdfs+XzqQMumqy9VOnvKzku
AtUUqI6mXOq/hlgpb6CNrxoR7p0Rkqz95f2NJCLMnbK2cDhe8/37vA/33ExoYHW0
M1D61n0UzqqQpuC0kCZ9MqpErgdQWT3RGbgN16p/YRumV7qDBdgZgaGj2mo/OYW2
6sr/9XqDS1m8Ypwh1HJbdqQS7oh/uyuJtMthQ4vw3VU27C2f4dfhOtg1CWycCBtv
iGrH3eP/Dzef5O9fkkF4ME2P5ZKwuC9sVyYKtiO3vi0rjA8JWYP4kECkA4UtCY6m
O4ToRCh0t57np20XTgGMGkbWs5KKN8jfTUVHIHdVmXQYs0OZE8J0xOtrjvOjILOv
pkWYAY/+qgAtVSuVsdOmGVbp28IKBfngc7zSm9iJKwW3NZkw5rRnL053YiRTRURb
wPYIC2Co4L4K6ceXFBgVN1a5iazGapx+ujK1pT0wCQ7yBKM7YVfC0woOz2+s+aBZ
zdGPsG/Iy2errtnvQitLm5IIoEk6sd9WaNrrWeA0Y0IafpX4XXzrDgMtGcWUQuN4
s6vrGJDuDihnhv5dwdHfS6nRQ9EygVnS85r7FFqG2KalKLnSAdZTIeLbf4RAoueF
mMyIB7+20UQufR8AlX5LhPWhl2B5QTJIh2WglZGpnhv5uN6VUgz8SpFtJSNlDp/n
WBH6CPiDGmFd08IrPvzdUQ/55yDSw+GYZNVGkDdUre8h6uRlcgIOtVOlOsFr25Kn
pEUm+4hDnCsp0m3pgOj5NpPwVR5OUgxWZWBJYI1BXjWXSyVo+741aGC5ScYG3mZP
rUwWJ9ACPdpQMOrn0xz/zyZMd4In7rkkm8AKYer7n4jI0TlruDXg9M/d0Rr7WIoJ
LfDp6B8ioXek3TcwW/KRw45ljpH+rYnMa7xOzDZvR6i9Kkh/6N0gTvap3BdeSyZV
s7TQwMvQIv4qMgXJiQlHdZPwZDHJhd58RI8UiDIIZiWO2fFzzxe7lCF4fytEFqmU
ptWu1NmAa/4R0UnKTS3hulUZGk+4+doBVR8aUyQzF7l0b3xCJVg9QLofAFAolPpu
a3XroWx+7Q7gyT6LrNLH29ADeDaJxP/0xt9R63pKOm/rledPj/g3V4t7lbk0bLTK
jGQdUsoVI/v+h6h+wyNiX6wdabu67ZQ0IlW8U0wJSU6z1eG/YHrjdRl17Qvu9HUe
3hfV5dlE9PxgPXXugimBpqd+gbJ8FIXw2f2X3snPJT9QiYBS3Hd0x6ghc5s/INnM
/sMQSny3Fks4IG3r1Z859ZY4i1Xg/xDGQHLYefN970WEnK7znItXLzVMVfKAXoBH
nVn7rCpEsxwN83i8SuKdL235iFvDoUiAAHLrFPqS06y6ukiy7HKF2+ic226LQi5p
lgqS/lYsCa9eNYI8l/BHqsn3+H+YGpD5r1b8HArxsu/8ihYShEswEVWzuOjqo1Nd
CNcNzfAXIhfnxlhP+g9Vn9XCJ3WD988t/1/udyHBpN+1Fs+nq7+wLy6cb0ap6PeN
yVmj01WxaWnC0fYTkdmciBqJdaZiaIUpXMtuwEsisktBToyS7txOGNSy2ivIsgxE
j370B8agbLcXk22xjf7B/7pA/sBIx8WnPCrqB/FOnyMOiJS+zUcCiTIGV63HMSYg
ZLK2vQamPT/0X9+gv+r1j05JwvPgFcrAj1m0riAzATOBr5M9onPMHe+3LSi+wi9f
haxgRum43wHGaawy4dc8uzVVQ/a4s7R7k3t56D7jAxbObKM3Aw/CGlipGUm0EuFv
703XPCclo55fH5CCEy+5Nd/oEeOcS57R1MMpnHS+vk9MDH1wH29AcLDqP89ojEcC
zTT/+YhmTiqhlxBZa5OcTDgT4t+0OISalWd+FTZQz6fwJwYaYUa+wFORihY+E3kj
uLul2J5vtErKL/MqFuR0alygX0ZsGLkfrXbQdTdrNeiFCedLFBn4zqYgooHkDbPi
3amwNppjeI2Ie7sazWE2lXjP0G6nhw8eccj8TJLbnl/U43xmRCzIQEfkX2f8BXZy
U/z8tzD8IQJaip6ogymqZWfXzS8HvFkkzuWsFPhm7MeJyHujLQgLQsxvQpx69bfc
xIQb2ZkcHQliX90mPH52z6u8EEH60XzrQ6ypRy9RnRKVwSpkTPKSBECEEhUJQ1b8
/uiK5xRANHXYDJ5MnBxuqYnIg5+1YDFDuHJ5CJzDUB5QLF/nWy4GEb6WBcLxFq2L
HjjvARDmePrKOCSIIVT/6GO0bFvdX+zKxhX+R9nxkg50gljmukRV3oOyS5oGQ0Dd
yHVX9/UTTRX7OcMeM/i47wqbz4hTWJlVc+qe+izBVu/CGn34X+p6G99CxGggtZgd
+3y7+mSaZbr8Z0psGWYY76CMnzrRMdnfCM46kAOposueA5nH4fEcUid/YHXFD6lE
tAgpROQf/DBdaG9ti1ytvxUHZTsEB8gtCAWYJwYwkKODCRSB+QMdTmIYeHLhYnnE
vzE/1u8c6RzinHsJhSJY9OdGfNzZvUcSR0Er073VzHbS6hHNPNSTm3EQ5sUExYR6
16US0wDYVu+SUDMNWMXdcCJqcEgoLNKSiJRkwsaGYyOVJIUPJngTS4A+IAEf5T/g
hj9rWji6El+WIk7YmPNLrwXImGbk48Bflz0yQAfasc52pD0s+IgltiQecV7jkTop
uverrkXWOwsbG2wgjeMiHBwSn1y5Bo82Lw/eEzAgZWQKebDN3C/YUyUmyRLEt/bs
qPVGpoXj9Tcg5H3KGr5ZnFUDo54eGcUOEQmUH6JJbujxmsAIRkx+yfxxRCsxxB3Z
8wuKvVKE3rk4qO19LVvSZrlJMDNsTy+tzyScO1KhIaWU+ND6kzBM2cm3YV/TOgiw
TfGbvElE6HbJoQmKbrq13fi5qkmHnQ6rndJ2GblvC5EUgv4cq0FOI3fazHKbg9hZ
3jEnW6Q0c//nulk3ZWz8n5EUFFQ0f6frJ9jK1ghXoXpyOMYPCHPh/+jsUzZXh04E
EYBo8mII2mKFTGl6/jC5W7uHxA8939NOJ1lDQATvz33zLVaTFrJ63yiLKNWFaS3X
+mC26h+qkwvuQKYBHmlbUMX6mxVqimsbRScAHks8I5aC5mNN7mx7R3Mn/nFUqC8H
1Q42TS3U77aY8xy3zkkjaWz0n673ELQuQyko+vjuuzMVJsINj2hitWV8SVF4TthA
AbAQtmB2eR545hsrKys5q4UiUV3Wgn/9Ocnto/0vJWec2vHGkylcy0vWBkI4HZ4N
1v80h+VT2GjxmakMh7HM6xDus/haBVtimpMSDuM0KPh2yKX9UbK1F1WFLv254Y/o
x30cupw6c37jgWjhcXxb8Eof7U1lyDDW0jcGvOv7lFPHUrQV/ZXrj0yBomwiBGCr
Yd8e7caxuRMD4JZxpGqe355tkSEAQbmWVjDW9Izb08dJw+ThN5KnDS3Xs0KYdNUI
2UGrdZA1pTw89cr82t4dSlUkHNcQ2HVPnuZ1r7bTQ7NTIYyeb29BBpq4k4OrQqyB
Q2twSaEZZybGufHwKwqG82DcSl52WWbhhDkC70mWXBwA5t0qtgZT0p2KmzPShAp3
pOJ/tPGOZjWhw0cCBQUKu6utXLzk5CqLN2Kb3pArWOLpvbG6h7FUfc9dc5INayaZ
OZYQV27eTpsY/HOc65H6J76aq44lV8XmX/TDqvpMAR0ORkd5+kp5632L/QZaA+D1
qhqM2DG3z6+ADzchSQsBijnouzJMONwrJr46DrBNuoL+ezHsoISqXWf4zUn8cikz
AfGVpWCpuD78IGgPC+4tnZwOD3RwMwd65kRjOmo4+HvgfLR+TN4cpL38niKTQqoW
ynCBlEo6vMkCYw07tWnEPlHKB2+mgZYUsY0pLYXNv/UL/euLrjNMTlu+yUusxVrw
H5KXBtGH6ldMVzB/3tDot3Px/rdNSoo7brs7t0Uqtri9xV+B4W4a4r5kTXV9d/9W
6ZR7FGEVrLuWID3aqfHqIx3JTYK7C2CdrkZ7TbURHEr6W+uAXPJV88O2rPR104by
EjcO3kZwpHDXcdK+jqfy/pHLProNF+PddCeExLCK5FMZP/S71NXGmurDNEmcgiHk
UuFIBh48xFqvfuUTkM1TZBa93qwCIWO3GAZVkce5ym5Vw22TCTmQSzfjRa4QF5GZ
C8krTJ8TFjC2HSGOtxEGYroOvy1hSVG4apBT+gnRk2Vbkgdbu+e/LIv4i9yvFwtC
zvRdwVjJT6SI8PUGeLMQhTWjV7kbmb8zaCdLZuI+RaAgbibkBgIG/97idaZjhUEy
wVzoYKClu+p3rjyBNfOKp0V1vzVzRmWqdKz9xeqQYDNVWLB6lC8XVe1X/LXxJFUZ
R9JKtmC6QJhOStl+FDRpTHBUdJHf3GOP07H8ozYgeMvCFcHoFugeqzHq/p9Pll7D
wsl17FemOlY966DxP3ORMQnoFtf/zGYj++qt7wRXj1mdN4esGQXejvqmr8oCj4Jt
x/sROUOnXlUNgrnrFyrhaCqtr0IshJ0U0PrLCidAiyPG1mEdER5nusvmqUGq42Mw
lKeqfsS1sPe67wI9SSoXhWGdo1Ccb/S/YFAjpr8qBFYysPv474gGgyMBk6YopAb/
kcdV+id8E1yt5h2qpucbcI3phapDqPZ4d3sQXc2BPo93clLsgcjX/uVfvouytTKQ
h8KN6PU3b/mEvEK/zkuVngA3sjDVpTRMqqKlrrGXTs4ncZxmc5zNRsQ3hBsH3lVG
awDAa5E5tifpvGtopzki4NHERPK+FSTvpyRI4EHMeg3/vu1K1ORX//bMellWxqWo
eWR2pPlcaBB4MCdOuwV0rhamkYaHWVYQKm6e44XaRj27vTC2rZQCuyfFrse01SOC
wwGI8yj5Cm/RunGZD4eKHMfXWrBu8tkc6hbSYA8UHhw5e/vmPgWiSDtzeTPaYvey
TWZ2sU/poYHeZvvrJMBQveprsCs5CanV4SvbryUxc30xpTBJNtze/XdOhawJ4sVs
95iomqeBib/lgk11HArVnkwhReu2OBzdFWIcYlKs86K/ObIQO5AtBC8FiKlaqdnz
lYzsfXmB+u9hqNwbgiwPXLVh4tZx/COBr+qCk/5EKaZO9MPcr+lcuLFvSzqtzss3
1IVXIgX2Lp3vnlvwlmqxNQH4kAIV1rcIVWmJXjnwpCDbKKHRK3wKfN4qB3KLZs9g
LyvcQJQS2n+T9Zck2vHrpJL0UWW6sewHmOE8i4HH4WrcSZjtLEmNrKSzY9vbDjue
zFAbm+XVrsedpxdpVzvCKYMhpb9Ot03QCULKqPbGDmfgTwzgfbZ2zE+CejB2csIL
keJrK2DhyNU2mUWDMysc9tJymVkcysHNnKooKx8j5VFueG6xQpjHhxU6I84WA1OM
UwwWPdP82GnPJsF6Q+NZ+tR0+0OJMoN4SS8dYV97YW7kgjUaH49Mt3ibW6QmBFEJ
Z6PLa6T9oKyOq84J+Y9o421RsQASEPy/7KSIUHE0lrr1B5VjfZ+q5l6Ii2h8KR43
F5BDV/rOF3SD8+o/VjaxmpJfph5LNcLw7+uSzYQt7tsCjuqAHSd0dBfdI3R0tNX6
ATVpIbyFwVNw80Fh9GDvKNn0bqOYxhPhJFVczYHtLehdO3Y2YFpp17mRiAAZl3E/
gM25Lcnx76/OrlmDymTVr//7j0MjjLViEoPdiAyigv1zoIpScB+X3417D+58a63S
FWBzug5jtA6TnVH4My3nYuH2B3aErilT7CUatKJFnoHe6OH0XFBlJwEj7YyN4pCQ
JawnlgHrhOzFNDGgRojIvpxJBLmWeuc46OW7K2lH6PJ4/CpAX4ytf5DNWs9/m8pd
o+1TsnJ736T4RwT5K4gojm9QttfFgMhG4zGf/3YBvEYHLEHfnVe0WF6tjZ7JADpb
uM62uP/+QinFnF6neenE/9e2nQsA0Vlu5TLOFK43Ret40QHVXb5ZEHGIC+Zp/86A
oVFli00gPoD4XCWNFuhIB4F0k2CajmVGICqtj2fTdckGyVJb2lcvdSQNyBLzWk41
DGp3EYNd7qIx2J1FG6uFFwf8/YwkfGXwbZG5PGcTHJgjEIoLdIhNxDYiuysf8huq
DZzZNXr3JFaXWppyGfPZLjBrlAt0PJjgwYyx5RfWyjdxQzSe4pvndA+FpMMtepHu
zWyvTjiX+E6k4YK1UlDSCQI62VOyxyUVz+fog89WD+2mHC3KNAYrawbbhJbllqoy
j7hdtd+UbCjMizgFi/09YNe3EAjN/Ps2FAObtjswEZYqiYtjNlOegXhFNSx9EpoM
kfIveuLtzk61FMbiYk7v4+RoLg/JPAfa5D1K1xeP2S3VWBm16EQxKWYcNvmJFQyL
VrkLfyhw1WwqFdDVGY6m0PWlRdGPwZAtUrTFrSeaGABS3+nhClH+83Ctazl+IEyi
7p4UcNy8EDBbrA17aBNapjfkYkThEbnkvue1Ab4/luYCe+r/ReR9NjLV2o8MJnfC
QDPvzBBDL4WRIa7wIHpIvE8dkvvnKlu1Sb03E2YaHwWN2vlWqSAYMM7Sca42Nyxy
haZSUAM2D1PaJiqR5s7JWGpQ+jHIejEMA5PoDJdiRE+Vzf5n+87UGE/NlgMPGl6d
NIcXyeXdLk99ueY4s71yN7yMkG7VEecd529ayYP24Y+gNhx51pXM5QVSSOz3XdTV
xCmyjqCVhZeDF3urq02QcTHii7MsOUTLlF4yML9KWuQgfboVJWejaAGf3fhZ4FxR
A/Y1lSbYW2v/RQ7wb4/wBf6yFafJ68BwaXI7OL07F+k2ipPXxvkMEzs2MgGO61gv
wpYgT1dAQr+Ykb6fBUUHxnaB+LLeYFke7R+koNTyddd+Nqo7KLTiiiN0krfjV3z1
KhjAbRihgNOa4BeN5uS9H33pIVYZEctjFmDfsPQkMwUGU8c625L2fxWs2pUVQiNA
8OxkcK0QvXxQhVhE5A3S5AgbYDdvRTYv6mXGD1hkKXUGxdD9CXtEaXJ9mrMKFULf
UBPCcrANBdLc38GgPM3Rsz4xgEHFYrWDWb6jSWu8e07xWn5o1HK1A7CP5ZTyAk4k
u49+f6DW9pC9TfF09qZB9dj7k4vH5q9Px7xYaiE1fxIsr5Lc3YXcawLUqQI+hla0
Q7/vRaXwSFM4dIAQ8F3F5wBy2xteaIRE+EvE4C6lkS7TJv16FdJLUqdm52jmaNxl
iA8EgHrEqTJ2F490LCCLF+BR2e+oVr3PVtBnN1ajRj1gblDDvVY28BuEKSYAf8zR
wCcvcCjtzMQPX9zoDvEcJTw/qAo3wxPnw/oP5cxePwBqwJcRdhm+CyFXepwnz15Q
irhoYpJcj5YMtNwmbPyT8JAuKofoDYFybWUIWWYjqBlHVulnuIlzMoUco6m5IlgQ
Lf5eTNn65jPzk48rEocEQi5Wig/bAuP4/RftB4uJhDxq8ySF+cXRVPzvNLvQL/RL
zi5GHeHHL1R0ZtgsQ7z3wkhM4bybHoW9lQAwUHQEMI7CZ4rxxCVaRvl5cGMq8/qB
Pb3SaI4fE3Z6aK6emCyII6UdCZkBVqKWd0ttQiPb2fj8DdRxbrsNvFmgXdqxUieS
+uYrTqPE0f35F2vkk7xgyON1hn6MQa1NLMSkBOsujQxr8i0eesaaCW9XvA7rICha
g/Pd7pM6m5yVqlzoWZnt7d5gm2UaePEbsp5RfHrlFaAEZmOEJxXO9CPW8o/+gH5n
p1y6uCgr/M9C0BIZzp6OwsdniAvIE7OkZ+tQ+/NG7yvvuEo9HDfNbjbVybQWMPi7
u3buHZIPdnqtOdhIKY2XuVQLU3u0zgDxiXDyWt5Gad3hmXeOft1q0scmVGKZ09EK
5IPoCXDb9e7m8C1d3McHXx1Skmw7zbjGzcE4zR6rd60gnWgFoc2aEwPWc/yolzYj
HG5WoBXp4JW1fOeAVTYMnYZ2a37VLo+zp/Nnth4IxmMpD+ZGi3P4Areb3BpkqW4+
sckEdQ6ccFYUY583qvOzfNksU9m1t9upqBOse8UEuDuqoAwjBEZVNBi/1rmCTYhq
R49+yHHjQ/JRRiR5+os2YyjnMX1f18gn5Q3WFZvuEHYBJPbO0xCAI0VER3RuOqdp
UqtHud1s/bW1hZu+zXMvZju675LBROv2NpfUQqAHAdWA0/ou5Yj6W4WmgMQlF3i7
63sOFE+fFLiqwLH7/jE0/HY5+YsGiCP3vjDOaq653awrrbrdzpHWQW4VZlqiGVl9
91PY1DEPzGfd65ABjuYv/ZtMn4gIwyH5BJ45uhccyf9w+8D7uDjXlDzZiwHWulp1
N1BW+YO5sG5O9DE2MkutmXF6MIJ2XnnjJAVLO+IRLzA3/blgKKymLQIvRlzH8kjP
OrrY6Coki6e27lb4VfjYG9bUkjpUrqC7pjPsIrriJCAucVyXbSHXLBPQqZROijHV
ie6ldJrVTP4+VN8NbGE7qdJ3hbxaFls2ESNJB1yxSSz7sD9Xx8kdePF1KazUOZZb
NnQc9lA+YrBf5cvTr4AqIhu093VVYvACIbsrwVzW0jAmL6bRSH9pPRIUyzWKVHl/
ICuW7CBT55Pw44KFyY9UNceoRt+C7Gggeaec9m4I5K8PIpn+wh2QyrEPbIqYPgTZ
awe9ZsDBgk4LBZxit1FwnKHUjA++rsc8bEFdihXq8YB8kayYD2P9GXrUEuJTqeGU
SlbYVTXXCZ8mvlLPmnhn5IZVgBHv0vMXrTo5yRbHWPZXnlYcB18SbaM6PnQFrMS+
6XXg2TQZ18e24cFyf8J+7g0iRw4qxQnYdeyttKvm1V5p65QEyQ7lh/yZI7kBmR1r
9s+mm80h2enLWDzaxlIHsAwLqV9JkCY7gR4JQlpBl3w8VFadOVmhFE0wNN4zMrFc
bgjqBL7JEzRYfgOMP6Kmtv/pzO+dUighDYdiL8+0T4H5WVBGVA22F/Kd1ebbRM/z
uwW3oLR97mMueQFGcGjruGrU9gCUD8748iT8S2NLvWDX2UQgyOPN36mDVwASuhEO
hog5XXYKt0V8TCxBmv5YI5USjEpe+pX5929rxy8DvuO7aIAyMS1KywT/Y5wY0MfZ
VMxHZA1qoBSC92SEyV5Q8A==
`protect end_protected