`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4128 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
VaA5/k9eGPDS+lyi+VYZW+OHlIM6qEEwybptMNhqBqBktv8xG6uxd8De8LZvTtgs
EzyTO6tbEL9j8ursU8JwT+LmYgnIUpRNGhACaWRMpuvg/n1qdfreasQ3/5PH0cki
ZNYwjj5u3toZwO6CAh7E9pIRuk46UqFgUA7szP0gTfjpZH32duVwqoiaM353vA/J
xpYX07LgIG7cYSvMLpWmUjP/5aWQQi7YNMtaUOilwaDfcsRpJsA5EoHreKXAFZXf
h85tsvFy7LDG+VojtDRZGQbSb8kT1C8NoAPvLV0YazoFetH2jmv4epX0A+Y8qUNK
vktz/6Okeltxr9M/9n8gnuxmhjYo1cMLsao7nHIvqbO/UAXDgOdxbKYvFFYqIoJK
N+WS3TszoLuqxZrVuWv1/GEcRlDs/p7S1HOellny8CcvCAyVD2E1CWcVNkkaBTXn
7tYFXSwcDNHd0ZRx1LoW/6lpzeIBW9iBBMFYVODpu66X5xuZJ60HMjMBEvEQM9c7
3Te21fcWBzm5HP8ZfCHkBCrTlmmD6G65UmsBsDkyutA69wYXbuoVADeS4+GkNKNs
eRcytpOhnPdfpC3jgC6X1p77mHtDwJArLLW/369h7hm99MotXzzVxljAoJIKomYY
mqQ8DeEMXeP+Rpsk+m26o+cryhHe7AE+yiY9f5GHRyiHSg/xnnYBOR1UTF8dOvFh
TGTzgcrgTX/xPfOOBpwc2tTTrwDAOdPQIzqdF5HDBI05x/90nZvOMBUH2GHMC7Bc
qsucio/qyCwZKElBNmgfLr0Oy/wg1y1CZCY6FwHBR+f9f8WjOGNUhq+pQJUoKSR+
kTh+YkDVT/ROWOwt3p5SpZSdufJtb2N1keRzAqZJbcnhJ9NlwF0/SRj4AaRxPH8h
m0pRCpsL1DTc+26JkLXnxP/vLW3pZSC2ULkz0EH5DcRUqzuS5UPs+k7yfDVPbSg+
BmAzYvAWmxlFsA+5bzKt/Ek+BC2SxIVoPU4INDCRffHjTHLvANkYxBMd1vFIRJll
zZQ6HwpTyj9GQsA9OSdEpwxWoY1i/Es/dRZ5wPFqmOVwJPLT4pIOWPsgcSndlXKO
MsnOX1phoxKxhSoxtRgJ4cf5A2rMLZq/7p1hCGoMgvrrmwjASR2GcZqb/yA8jaCk
D846DYeUl3blk/SEIdrBOOfKJSj760vYCtDGPpMwvZwxcaaJGCbTlFctDSHgNdRJ
EDZjyUYzJz2gU8flB7GnJtAmsNUKKXgJOp3ozs7T9oS1EKOMLy63Oqf6ey44ea2f
uBcOTmKcEvYEcTNNsf43AbyndMKyrcgD0Da62WUQeav7biZGYEh2u5y7gPD3CiqS
Rsbg8wmy35s5UFnE16tN/UTsazPsc3aLLNOheCe4U0unt/GgNOdi9RFgpjDWvCNH
aJEhIpj3Fr7egI+yO7cnTqueOq9oj2yGUqkK9MMkcxEQ77GmmiXjo+40mDWkjEWv
yyg9sPwrzIk/JUsWpOPHSd1xbt517E5qEvn0iU1fBpabfmQnLa0DaF1GE8UHulww
5dI2YvbbfgxVIcxuaNXDjwxAJcew7jBz+U+DcQPtx9EnISv5hVSGNW/RG4sCs03Z
xfZl7f6Kf/mVwZJrqi8u7gem9yfiO/oZzluuCVTgBjyIT4DRfJNshRF3Pj47BSyf
2uQwNB9WzbOygFKNk/E5ffCnDyRNd60iZxqXU3ZaePE63EKF+I6kSi/7sbCsdHOj
jOdUVoltMmxHvdK+QTM0xq5lUtO/yQ1pjIpWDIQd5wrsnhNNcobWlTxyS6scOXsT
HTPavutiV1+fxJ3p6Uf2CD/yB7fohNyt671LS6Oah4NvEHxeQ+Uv5zRYirm7OwcP
5gJMb+ESdGKsNNyBkOAIO3qikR2t9GZr6MQBJhJYIHMpV5TMTLvj6bHPb4CXNAPK
/jcgQI9FA//OXRMBfaArNFvuU34jxLQuaUWfJlO2XGXu6FkfH4pAXutomi3DZI9i
G+YWvceMTFr5ofd6HILyQyDHjjBfEuRsuZbOzmijZ6GGT5jKmph4980pyo+Pqq1M
yLRm/KmXqoPLj0vY1YDGaPnkDXoOgCEYjuMK7T1HdIFhFSVTTvLDq9hKeJllXFG9
nINQ4w55YnwIFMi/kNpWxXdVg1Q68K+dZjwS8QjOjuS73hiQtA2idqOkEFntUXIl
92puzfxSWY1tKLHElCZEf6QGi6LPv0PALOsTeAgkesQhob/+8Cl/TLKtxWGL05GX
EAJ0+n7Kzn8Fd5Mn0a0vrjWjkYOgnt+s+m355d24MoYO/jdkP0lxBG2vfHCUnqIR
r1OzEgHZUO23V6l+G+WburKPUJzSpJs15ZIpw0puC12dihcM541gQ04RGItLoGDt
YSyK7nOPJ1Il/Je7lv3vr0PMUxNg65LuS8O+ycMRvOeJbwHk80kCb/guMplWXvcs
mQUfFIe9ynyjzC7W9jQ/UAOkrs6tD9wYibbxc6dF43R9KqTE+eC8a4/TcookLiIw
WAEeO1F99EMmhWEuUzTk10M8ST9ffq8F3v7ocTKa7RmYsThsz6L41eRBu8mbE9B1
cvipBqKdrpe6CzuQq/YyE4BKwt7Ij6WbBMg5i6M8+yb9cw1mpe4H33T7E0L4bUBS
vUPvQ5zRij8kelIMM3ZCiDrhtMCNf9+kmhPc4QG4n1zTpQnZPg6Yi8gMpyYQ+JOa
52eO9tVIuNOJPKQES7/Cac5ItCsi4IPK2R0cbwG21GsN/erOkabaeooTMbXfzjSi
BhbdUY6Jy+2gs864ttQ2xDHQYunyhIFCXtujhAy+gkB7C38lJ+JqSN3kJk909kNc
HWONp/0Y7DFW/Et+Um0JvVEzUiLHU4UFALOpLbcbSm0kY0jZsUShJUiz1Embb8be
/YaADcrmNLGOXp1yx5H2YS15cci63k4Kw/dUUI+OX/fFbmu21uj2gyLslqmvMtrb
/EfsTUa5pz+3ssI/J8PoQgLK65uDd0F72JY2eF1DMF4xlb2iSrnAwJu2GrcfJ1sX
D6us3fay22GDn2lxWn69ZFnVjtSvVHXUxJFmt0Tj3Em/MVGNgZ3L2BTCEW5k9gJN
CmOonIOJlTPIMoCIa2FcT102Yy7ZMMgswffr//J40KVIgHXneNbZQaw/aOV32vrP
3OAcrMa5ZIdfSHRcdEe03n8lvIppUMpeaMvYWExI0jYc+1TTRROwuAddY/5a/qjE
+Ag8j5vC+3vQK8V7uAHYJc0d+GGIRau0w3/HuEES6pmjARasYQ3FfGrumjvk8WYw
vdXogzjuQo+1j4I4NvgIefrvANyjM+WkbD2/SZHXEzmhCyMJ98wS4X7xUpq0gDhl
FcI/ZTdKPzOpxdI+gCXFhxxKcEhqj1OK67DaBZWN+r7c/UBemzgiId3LEC6j6ezc
N8WhAKIhw1TXGANepaNiPhHfIml1q9Gpm8JlkOkfGI+/6i1fUt0/TIZC066T37sE
dZangYogPRhSo0teCLg84xmQQIvHPRN08JjZ5nEM6OwxCYbupePCddM/rPdfMQKR
mu/p3HTK9jFChJ5ONmgDguyZUxRgyR02M7xxn/lgqrSKBMuBAP5sKua0kzxIzCl2
PSY65wBmpVtkNTauUucZz2vbj6sERYwNNiIpNvueP/XKfdPllvIhtXekvt1QI/OU
joH1gRsidy1Nt7urMIdxDpLIRDRQ9mUN7V4L8YCJVJISgXaCz6fp7dAnVoz0FO0b
Uf85ZQnJzvatXMFDSawEFZKWPNw9vMa7e5KKgO0PO0oRxBAdywbJ3sz7YWutHMsn
JuD5UFwDWpAanIf7Cyl9Y7fFBGpoeFps5juqccpVdZmQ//W29ufOYOi1DLpaaUb7
N+RyspurfyZwGfkDKwr5X3Zfltet5449fup64AIKTdhOnHPy/sfhGPjn0SSf7ZaJ
ZifeujbqrRgPopxAd7SXW7S+Mfrk2hrF4riDgj/Aj4o1wFIpKo7H9k8HcM/oHSbf
2X8njxSkVIaYCIpqxhL/iiXTg9ek2RWm5/kztB70LjHil/d7LuSbuuA4t3apks+M
+YF5Tx09bnVyQX88Y/Kz/aaylVj41IR3DRUtZjxzI7BdH4hU7k0aKo9IjXgBzeKs
AOYWno2WD+ZkxInDxbkq1YPE+9Cg7tuCy8zAoj00ygzMQNAkc8Nw8NPs8tREhbSg
M4YtZnASj++0XeqDvr5UWRkc/v1nMrhtdRTao8kBV95JG3M91/krrYxghW1DsViL
eMGHj1U/7NWLe1D2RAl/UtP6DTT3eIEdKJbE5e98J20lI37dekQbI2azfllzRKGE
Q8zZPcA6v1UMzKH6T3TpThk3wvmXWIU1Hg6MmGB3pDYwWlgNSYUxYgEOkM4UmLzN
vFlb1InghssyfaT2Ql1nniltwbe1jq9lCYvE+pynpoaH8VCcLyDFjT2Cy+1QfGf+
MCCnVdo97Uc2uLjnOq1qvgcArK8ayAe+PN/30Sg+t9MA5l0x2aSiHAfnie29v7Ml
36ig1HXif8nfUOuRQBqGnFr40wmTPeqZGJVTURGaGrikP7APzm58pAPkTK0thv84
PPVWl+9gtU5+Bn0OjltrskZyGErqmyh0oDJ7xTWeRYZqrxOUVJR0CA1v934UPrrv
Y5fzN3Yj6xTQpanKJz2MKD/N8NSUMeBR2t4ivzQzghpjvEeiXydZmvSsbqPDXFeW
S/RTBsTCU+aLN7cwFcYN1Ebzj84wwhlNyHBW8b1dkKqAE8FpakYSUi0xaHn2L7y8
qFIj6G37EzmzDvawWoJupIQOgalzhxkERso0YGOiS2xQV+x/0t4L0U2W6s4coSW+
Ot9qV7zM+5IeOtPNsWLkW27avdIeYgj23tcqf4ln/kun+yWoJvujrrD6rrbdHKJi
dlrMIXoIS65VC1SuM0j1BMbandeV8Rocf3IutSAN4ZhyjDITkPVX1RjUNXDpjBIj
BJPupS3IaKB8mimQOdfQStB9JYCuPJOZkAQR6s0Rz3jndBKoV1BDvF0Y3KJIQ8ot
WtEcf29mhoib/F2uwuAwLBcVJtCIg8b9KHs5JvDOG8mXBGT3Zyst1+0tudsMuHLx
t0ekOT+I/k3GjyR+3yO1P8hyep26i2vc9G1tP/41g4oUwKu+Je+yykMdpFpcsIi6
bgvZFyHt5MeeutdpUUT2k8LLe8Rm3X63LlKRNk0+GW1S7XsQnu+2GS2yBixCRu+j
RubMgAxWb7Z2Y6EnOO0p0lrPGiPIR1lqB4teht8OnoMNSJ8uCPS4JO4rBs2P/mk5
GRlexnrxKIDmH4g0Uy+XMrdsdOHMlimCJBYrZECGlF2JHp28iK2U0EDPVY2aTYtu
bBLMckSDWrTX0GHxADHTE0/O8ztdnPtDUtcEfHtLRV8QHNdAcHSuVB/6KqEZNuNM
`protect end_protected