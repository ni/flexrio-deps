`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1648 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
/vEkqJfyK/81z5lf9X8oFQq0iu+Qc8SYLbsZULSaEiT0mxWTl5PEfR0c3/Zrtd+z
b/4glKmQH7b1l3m2bxuIPr49ipUwe3JhzKp1O/c7iXGw9X9pnOnEbvhYbd27YLL+
SX4cq/59v7Z0+YzLz+pwSqdCGXbPanYo1IGS+Rcve6pGGxAivTpUfkJUwjY7/xvx
Bg1wlH/JZvcXKz79a5M+wFkfn9OFXGzNGSvNRgqAA/80qvA4xwkjMHlD+kpWXOFm
8Jr5nLlTo7tATV9gS5IJheLGHkRsRVpmWbHYV7LCcZsx+/DGyYhhn6b+9Wlr3KZ+
oVizFOBSFd4/bpKwYHbhGefGD3PUxvInVpcczQ7BbfVvTVhdg2Gbrpb+nntAHdqc
2IUsfUs39Q6c6bcV+OxqiRr3Ve5ovP1IZXQLYCVICWOzQ8YMlax1DaQrkpAVnClH
nFyBl6S73DalW7crTuUMOPWDjqQA5sCPNosImkOtFcgKjHKKWHThVnyFDOpgnJo8
7k1FughJlbe2NGsSaP97JQ0xAxO/QUEYKjXu2/YsgsahwV5cGSTsZRyvb5zfWTjd
JuA+unhoBcE/7RrRWviR/9fpNTjnlwvxmN2Ynvpi1PSahg2SWUKUyR9i08/0f1sq
N72FomTxZflhqPC5Kc8eW3+Uo0cQ32sXvIxP15DvUTbWtoIb1yCkqmsxS+j6CsFX
m/5unQNjSQN0Mv5tY/6Rta91iXVsiwMu0R6657imglGVCHAgLXuOGOFllenALGEl
VRfqOATirMIu1B/tRTKiniPalRml+3f7gAsbjzI2sa8u1N79KjPoWh8bvZrOBzo5
aEAq90KiBKeT16avxajTtpZkIUNE6Yx7v8beAhAkaFiTSyeLD/YkndOhzqHu7KN+
ruwGEWfsYqEVqRkq8EUnc9uKWV9wQOzbjHG+jK20dnwLBNr2qTBmqIzVxPv5A/ci
27XHUmUH3h5R8Rrrd1DPX9qcQZiWYyhrgvJZ05ceHU4A86Wum5AbULcxm+jRz3ma
A2Eg4dUjOy975y1CLUfxEcT195w4NnZD5h//CbsSj7cVLOocJRi+GvqoWGFbs06y
ruvF9lOPkCcQiI1Y7Iib7n9UtS4yK3VGdiMdqCUGcewNXMtkIzfnCTnjxeolyKWe
A6cBkYSm+rFoEjQpQ9eSg0G3W4MpCb5WrIPfleFueCRDcM/ihhF5F+xQqsOZhTbE
B0E+drBBV2k+UiLDHMpp5bVt0BQ1ZJa25xezRQ0Hc2qQ6BFbDhr+rZmeS/YDfWQP
jGyfMmuzkLLU4oZ9lYgPUVaD3+S4FQzIMvwht4mxJpptzItKDubQswcen3GYBbfY
WJLP6/lFb7BTu0oUsk2WQKZ2SyawCXf7soKXLIxigQDPYsqZRCWpOCddEwsEuw9x
1aLYSQWpNFtqsHS+J9BOxkcF3A6M4T2GXHzpKa/dLFOUMvBMmPhpA5CfPJk/yj3Z
ISnN6Eqzl/S+vhsioEc6I9s7X59bKMVIOlZYTvtgXmpVB9bz+i3vZP0l9t3OOYWe
k/fUqzWimwCWOjlJx/k9HNH46zHby58HPptxkf3MswfTYhjLj56tJfwBXP5gJFyM
wH/iZqTZlArRtq+YFRE++tQXDgLKZ3T9+IiXT7qo2+W5GInKL5s4Ba2N6GARa4aM
1PvFOjtQxFIiJcUx+Aefc9uc2+YFAZi8MD7+AvL/sxLv8HrWzMvC+91oVs1EKKGf
RWNMc5Rwyzz8BsbU9GL9PvafpniMp/aqldl30kNQY5i/ln3M6Hanz5kGwn22k9/Q
I0+FVufLiUWbC9j2YydsXBg38cephK70aS2VR/9u/chvCpL+JVKftDIuyzQKR2Ty
uK8EOw5WevHkv0nz3n68Rvm8MVzqQHwVIdvZtz3ELuNxXa93z/bwmci6Hft3Bq1m
si2oLP7/6Rb1zJcM6Yf97x90FZcFvS0xmtcX/7Tnny8+pjH4bzVnBHaMxw12155n
zd7j+4ia0Nf3hVo3tEYEMD9AV/IlSHvUmbKO46zqaxn6zxtYGHLHu0C+rULI7+cA
PtcnxlZBJh5V9Oh6HuvwYw==
`protect end_protected