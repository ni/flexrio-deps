`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10080 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMXpMQW0GqyMEszS4PQs2B+W
dAK4WoK8xrZgmxcq+ZCWAbXvSy/1enpUyXJQH5F6+IRsN/WxlQYYOoUWm9wDn9gX
Io1RBewTtCI624pCu7wM3o6o8jo2vpFrrXIHId0jaN4AZvTT0kFwIQgkhUtOk0Jh
wHrTrcWcI/2wHpNXsmPCiWACyDNnwLvOwwv6pK19yfQTzO9/uPNc2XQ5wPfzblh4
829R9lpzfuWXhWBHl6m8OUg3ZJsWcn72M/IH+3jIfxx7rv32kRG+KgSPofmMxvFR
HRgBCbzEc5N0E3nf+7fSRNgFslFRyVl6pfKQHLZOtNPoZ2YFoKbDYDhGdpO7df/E
H44yVHm2855NKUfnGJ4GiFS2g7E/NN7I5qRj8HIf8MqTNxtD3kBosFPtI3xtfFc5
Xz64wxTxN/nbMri57ahxIXv2Qk8gjjoeTnqlbDSzUOQd05je9j1v5Z6CvJ5rAgs5
ptOujTZT270cKUmij37i6YOhwvpiBWBlsTfcunjkhG3qXIsi9RQNc62Nj+tnsYab
lzfyt3lXZQfGjJnnNMI1Iniw/jbkFnx3EjBiSPP9uejDlLifN6NAmqK6PmYJaS70
U02aML3WGO/d4A8u0xwhrqw8NfwuBuoR07TXGekPOXMrWj7/hyjitRwql/xeR2DJ
GC700wX+kzPDajMQALBFo29JpMD5GES7FD30IYnTxA5cbiGNzzNB7F87KbzboC4d
NpxFHPPe36yX7Jvfncu8nTgO1kL6iloD9WtQz0DuIMl8yFcwRYlT9XDDfp0RDeKN
HVbJaQuRi4E1Driv4uYZSiZWwVFJflB41hfoW5ZGk/eyduoWvXyU6hiG5USWHQJZ
pFgULzxV9QbIRTahL1iW6sWkazSOgKZ9mTGfbzIT7zxodcLPyYDarDvZZCz1z9u3
w6d+J/qACcgigwG8wKCxdsJj0ptl67jJuQtt/wBvigY4zd7+v3RK2Tl0OEKmMHZh
ZenAWY6rZXn3TlWmOhQRDD5fkohZzEcTJWvlmYXcYonXG/vG9k+YSggQZgkQnfGJ
PleHxKow+z4aLwsfBwsNKPSQkAzDqxfAwzkrCwf1v86SMElTXA4uLFuJVR/LivaZ
6PQK3YdaX75RKthPP3sfbY5R0hXmLAZ0VTpcnLx7blsZaNcozk2iOTrd6VX/UKUj
3o3zBuLFKokeepyeH0ipetI2GnfGMMcj1ueJAtuZEN0l13czJSm1grDy82X1qzSH
L2ZIzeeAPv5swvNGxCLmQytzQmmsqKwSI/WX+Sh8M3gJqPaIhyqgq5tWwXVxyd3g
v4O73v6Y6I1h2IyG45i7auXXFb2Zy3aPDrkOG0sqf5wV5AXCaSam3WrwykSt0WQY
2r43kYqJ35Rz/HTfT0p1m2k41BxZkFIxhPyDg7lgt77GhuQahBkaZxPkMmULbOvE
vBJOwLCaqbdoOmMrwKTIXiIdq8n1HTmNKguJsoNzyn6ceoXLbKukG5Qz3J9cE/ts
eol3gnOao3hwjKhEwLqfZEaUCqe30SaPgFtHw1vtuheYTdrUw6g51xn6p0gOxH6t
FBWH5+w15yKPq4xHokNYfH4lWrldIYOUpl0fp36R8zhzgQEvSQm5kXBmRcxlFCwd
wtF9B2FswJfhQJuYT0IVYhx5IWLvwnxhCTITb9nJ4DqDLaYyahjaN66eo/LHAyxg
n9ZRne/2LEyh86L9rEPzDxWVefHudyjISAsh4KYufTCSposi3a5ECjwbL68VvehA
ATBGgz3TO8gDCaNuCq6ITVBNxfDhiwrxMbSgip3zkVk76r2HktB7SFzKYl28n3iQ
YZb8ALKGDVN9dP20OtWOZaDxzYEwHN6DR3ePDLU4NZiB8STdb78OqCOeQparqnBy
nQRLDNTygASvoQ+g7Azkfr5L9lOUALKxRuPHZ8HdBST6qINViaNM4eiw52Q8LwB6
KIui9AG/IwondSgxyWFIVCJYZjpHrRTal+0YZ0QjpjYGGjauSUp3oC8s4fzyMl6U
GhPVOcQ/MfIQdschPlzTJWT9k2uA//MAKzXoannolGxxWPFGo8KrD9OBHpnEfcgO
vAxyxs0CyEpZnwNHydzMBlP9BS8mysUL7ZyFFckuZ+UD6mlVbwOM4IM1SwtUH4+D
RQJQSdhQQBZxwdtxHkf9UbvMDI53XzQOQbk8fS9IS70HV355f4Gu9sGdErVsqfJe
a1V8SJfxSiDrbgyUdRNaj+amb3p2R5f13LlKukLrRZbHdbUgJKcrValywio8O1yV
TeZw7dgsBfL2cPylVwOA6FuPZkMEOOqR2TlyQSRVATcKn4sUVmziB/vX5mTocvk6
aM+/IsUzdFgh2okmuJm7+zQS3Gi1RTh/O0fWn/Ejhw7v3Ul1JMeOkAIT9rWANwcS
SBMGpdCuiomyfX4Ya1o9uxkrqwtz7GRI7VRcCmnE+uek5+XFrAvZSG7uZyLmKWI8
ComUatHMnR1tOFM+w+dmrNtDVyL/sBRE1EYc9OuqQAIwARnvpEK5auD1D5vKYnMx
Xa0HfulgJWMUimG/HiKHJF7gyNYNTMQPqX+3UioBfidj577Z+d4Fgk1RLFcFkioq
FRJsAWhPjECimFFBleMrXSLRZlcoIWfAGHGdDTmto+f8hWIsYxTtre5MwLX8J0cL
jrset5jvjfKTs/yXNQOoC9oCWoYtQAamobTsaYcMy7LqxvcKYpoUzsiSi9BnPrOn
Xkep7Iw8md3zoe/VAwqhSvkUJMghpjjhrBQ3ZUFHTiAqMqSqaHSkag6HPtSryiq+
UotBkkVNpp2/OeyJO7qbbWlSNDwGfw69aGHmJH1pOdfPOEKoBW+0UXzXnxGRHKsx
rcIeG5vDXvwBaxczeqIQSn5ZrsHayxE9lWQENdtme8JkRdN8lsAU4ym8x48/YCle
3q/XK1SpOeQmklvz9tTAXHeIsyZfBJX5BxI4iUj8sdJYN3Ti1/V0Liq4p4inO0sU
3DSmMe40cDvrhjdNYBXlPvH1tmIrPWOUpRgzSQqN+Lu2E7QNQZgA6HH4qWujJewd
xgRXMmLjqAZMXl10W/H9z4PEQEVdQRFJnZ8vdls4xD27k9eC3/Lm87YB/KWBFUG+
8ZvMtf8/SmLXdZuJ297u2n47fDuqH0u/MjJ2RFBhFc+PU2on+WWc6l8vOhptbr2Q
Hi+L7mIpOYiPKEY9RPBZpNtXk1MpC0vg4QqUrPjvf69kPPpimiHF+4OftY4kkbiK
fMpcgLYZhhuVuGqVEEACReTe2jfg17r2N5dTqPXop8tL1UsLUceSCQ5pty84YSGR
JtKds8Ucj+AHbSlaXYxsZhajCwlDgVhHXRyC+CPsh9mpXR4RzV2/CogVZIKFWU02
5j4nAiiEfY4fiqqumWK2/69rPKBqwBH454Zr/JoAb1eGVuN01a4/vRjm9bXvs4F6
BeIH/IlT+Maot06PhNJfvTOMwac7bAb5jTPLWmLCdSMyPqyP9xhoxKmLFh7m9NUg
fnF0fU5qXbknH5EYmUTRXhOco+z5as0n6916RY5hrxYqe0Ts5jIwbTZnjrJDzieH
lBW5Yy8I6qDuJ6MArM2gQ1jdFXAMy7o/A3FN7eIOmzYvyW5hkMuskGFBkjR1Mlub
vQdgHwPoAu3U+/zSZ5j1i1AgKH5nynGW0rshqWlR2PBtj8nDM1yHleq1mkYkRg2V
VBl5Lsl/6xLlEV5MkLJu1+soL9c3AmC31ClkbZNHIklbFjezq5sOxKinE89HkytZ
F/tn7hIKeCUO7ZaCKQ3cIWtv1tSyteHa95MPOBLSuA2aop1D2RZQMz7fOKsQMhp7
FgXamzH00MCsSJOMs9DpAUoEKYQOYR7lzRHEWQQ4CbwPxtwAPxUIkdXjW24dyFOm
nJvDKHXV3rCS8cjtooR01MFuwbBD298ZlR8DW/V/nCtTn3UjAAZPwlKovFwwHGli
p96lDTXN93Ggfy2f720ajwDkWw7W9Fz4zP+MIQ44OXd/0nN9YmjfWW2grN1zCfs1
zmrA/p2uBqScE7OjeO8L0O3zursrxgNKKbk0zjsQBt76ZKy5Q3loatryDU4eTZSO
xpstcP4neVJu/EEhGxc6JqLWOmRx0pUmPyktT2Zyr/NXoj7UOkn/BTbYM5FiSrkH
NzO7nVmNP4xK+ncPUQyUrPNXBCELMAIPvTuKQMvKQxxUt4z4h02Q+qaVpDAi0sEy
/ze7SuDatCoLM48pl3WFN6GjXmdaptSKp6KnS4Nyj9+uvxiW6X2HeuLyKF8bg4Iy
7wNrnfa/MdNTWabhcxSpeVPhOIOqBXeZDZENlyI/mHR253RYRp79B4QQxejj/eAQ
rq37qTPYDVaJtRY8MTY1Sg9UUlSTUYVR7GBn/egbw+Rt5pPrsJ4zXCA6m0Do5DiW
ILHLaOKP64EVw6fajySoHSfKn4pzAcF1FJpKPGizAFhyNDS/y66sl8ClC0k6250I
IkIivaT9mSJi4xGs5hYLYtPuP80+AVvxWxIhZQQVHhaQt2ua1qlFUBKW1tDKX8HD
VyNZx/zV12+LkVPR7HguiezPYhUigMmMkRf0Ycli/OAZLN2SJuFylsxO9Kgfslam
CJCz6j/FA1HGw+rrPa4owbfLpeA2yj2qQiBlTUYCz2AN2LaULmMf99d667HGoCgu
8r/6lQY4aA+LpnmN7I/dDODQand/mCSV4gQyt1mXZLSRjPtb810LdCImYLPug2OL
8DT2iD/a1bvy0wsNIgtN0sFjhqMTNXq52gJogjnqnzo1UFhg8RTvbAx7y6+aGEis
+f0VxKWeTDQ6OmuUfxYa65XCJ4Ah08WkTFxEwTXg1y4NG1j+iOxndOaEfFWVVSAj
+/7ywwLeE1rwmt1nis4WGT9/DUQH+cL2KbCrdMpd3aUAFpYeRfx1JgM3CGs4swjC
EP9ohLLTzyHtQBIyG8dOXcKKohPyaX949Y07sCLqOcdgUhYWSkwZhBX79AtLN3bG
rgt6inBAW1Ft7mrrmLiz6sHBMyziD8rS+2hNLjO7b9lh5Ct+E0FNd2qarh9XlWkj
85CoYV1YoajU8xTCEzPx5ZHIDBDgKP3jZMMQ2F8GRwQ4PRFx7b3WhUzaC/ISQe7o
d2wtT9aNwVBOaS6CM0j7Bi0uXDGnBLK3IyAqZ+BgnNKzPHCEpDOdVeIfJrMu6Oay
hv9uxqnwwP4X0HafipvOQz0G6WrYigwUPkkmA24ltVkNVP5XfgPptaUUaIqmKfje
PS8KZazptDPmnIkexZhq9CbQe4liugnP80mKPtqdtSkcTDeP6gS8dj/8+3Zahe92
mwNjvWkfDhb++rbATZoNBVXpzcMOGf6sF0Tgqx25BlpmgjUEu+tdSLBasmiazxYh
1h2KIy23X9TMfEzDX33CEJOc+B6+ZrUJT6tr75QWR0XX1oFFtE/NpADmoe/Hge6y
m/Z1TmIKbPKZahqN0UR5q/JxCe3QNMxmb81nUhUzn+G0Q/vKOzyX0W5tfKJ2hyo0
3xZJUVuqY01ouOXuCZusWuHTFhoRTBpXMJb7t955Q9R7xHgUpeD4eChADfpmLfZd
soyLoAQRZHmfY0R1rKYIfLaYerTqtkx5/yG7zGVtlP6vkgEiTBv5INk96rTA+8pO
h3wd5lpqEwioWGBvC5BsKTlUObPmHMg/xPTQTId8fynUWPV0/nWgSPZBKW07LBYS
9giRU8PaUC7qke/XGI2F6rDGLRoaTK/JlmSELG1+UC4EilvtcYNvS+yvIBRfDadK
m0GoER83L5/19HCW8Hq+G8oyYyj32xjbCPg5RXViloooeRxEfd8Lbg4rQIh3Iere
d6ZZNt1kGrVMErCygVXyW9ATpt0dFCeNmUAsFNq+WuIYA4pntEixZw72NufiWMT4
YzwZR9QpygmoLbWErL52t05w6AMgFt1sy1WyWCYKHNzcnG/fM7TB1Ggh5nMtPwEi
zywzxlvDBsdtwhG3tV7ZPS8AJnN8rmbVqqlJxcocQo7S8TPsU6ggUXhYN48DuPOW
KON4gcynxr4RXL8kBRG4TuIPDlqR/r7xvLVO8lqbpl3J70w6KldbJYHHBEX0K9Me
dzVbYdYE1GPxYoZ3YI628UYNfjGN3+NFHtJ2L6Wkc48ISOHumpyHlbeGfHUgbJPK
MRjU9uFPuNwNb2+8KDyT6a6llAoiDitc2Ibr6xeCsI2dhbARXzTtceq7MB0+SwIP
4M5CGTuilWpKTGRR6x4InfRQlwGr+0crmzqZ4wClsi+Ib7o6Zi85Ldkp3tC/wV8n
T5E8fOiZlDC19iXZuWQ/YJlBNjcfSPYRbJEtBfCAHh0X9Gk+QoEbm02OJy6ZP5kA
kFjmS3ry5UNGS+WkJa8xowLIeZFzfv8LjGHpflvLbFT9ZLHXG091PSwfuncumq0M
jv4vllXhHnVY+B1e+KfYOwq/uHk1vZDLy/sg7gyCqVG4O8bQtEM6zdZ4/tgQDrBU
12m7M+pB87+jL0QrHMcfeRK+TGyQNOUHlZ9Cou/vZahA4GbC81SSpYadFQ0EBpZC
9U5q7TsKXiGUg9UHiaf31vCbPwGS1N7lr5cN1630ln9VcXUIQE/LzE5mLtfCZfzO
hoo99WL6Pv960z50Jb8IrvAzNPq6JTBGy4VtIwveEjGQ3xg8qL74r3WliXjDwEFu
ukepIBIvXe2iRdMGZ6QgatnEjTAHFe7N9vhJiZBpFE8ULcl6HP1yiSTxSUxQWR0S
57O9SDbKpk5Hm3SVO9D79EVT2cKH1H1PA9h2+ul/ZGL4ni0O+0qX2M7B8e7gapNF
0EPs04/112lV2cwF8yMcFUmioRxXLxumWHkg57Ts+ZSq43wXd0Px9G++x2DIHAQ3
Dk2T8y9PNO5XNnhuXyrOmWyLRv3MjkwgXsf+P4uWvJsRsg8dSZImgffCqLQGBcPp
LvtHEXK922pt6Ar6DK3S4m0yXg97CP0IBAbNG/le+j8OqEpz4kHgcfWC821mwRlM
aLp0fJor/QkztESYpEJIkxMFHUCXI7Y9kvc9HyELRgeR0YGPSrgWw616tR4qftlK
qTCANBxfQ4AdJ2H+7syJwuquHY+S0w/1DxE6w/I0P1oc7v/oSkVBNw9xuDq49y8C
AFarMQagDGvD83lU4MI1OgynkFnoPFVqLzwnTbv+c1iDndFcHiN+gLNeI9jJnRdw
Gi6Z0mlGJIzOWP/tgsNvEfqzbDC3gWJnjrUt3W4PcPoZLtyjyNdYqGp8pUxx2LyM
kR2KTiEIQBySrveJbtQA4wJl8go9ibksOnPdAWkHkc86wi1f02gO7hajg6XJDAf2
I0nmM9xMeI7xszZMxzoJ+rNRTgjETgLPLQAtCUZe9htFUayHyAl9Q+o4+wruju0k
q4ZACWF0HBonCcrTU8TvXVw8F9t94BLQRZLH6EgKHXQgQfMhLc306EAYVDD3hNL6
bDTXjjJt1sZtfd4Besa00nFQsDhtyFSYa7zMNWez1d8MBYyZfRjIB2zQx74na2xv
HmzWA7fnhyk04Yao9k9KfqfCv7l45D150fbCfH6GS4OpAbgmjcBhD9aQtMtkCJyc
UDWrPjIk/QM5N58k//44KpmqfN+DHN95yT25CRbjK384kDWn9qdmsqoE+fT/oPFx
LeqbK5HjFAIMG6Mric3JM75uIcm9iF6FmLSrD/PXh5RaVq1ffnffDYwf1Auyw4E8
9gxpj5CwZAw22nWhOKlNlSpD4VlOwflys4z0ksxkrhut6vwtT4qN/suy+20T4W3Y
GxfiPH34qGBtI8nEG+xthHG4Zag83C8RgmpgX5p4TmOf/f/jwvGF7I7ZBrecS8ct
xqiyWNRtCEbZqB9vnUznNYbuvVGfcTNYTyRT/GOf7XTOoYISGVgpiIqkZ47HI/6Y
Mw9z7qs2smNSeSvPbqA7uLy4MrJwCT9ZamLj0d/dpKNjW3afYE7vpKaUCn3vd6xA
xJrbfwpz4sG91rCa8yY5aMvKmUCvH/mMaKD1sFGRJP5+bUJp9ZkCMkQVE7JMdMxb
WhtbEWa04paBSdD/RALpo4Q3+JELivu9VD+9lRMMLr8tkdboOWTOYqw0CH4Cz1Wu
s47ACpXFvhRYUBD1oM7gFghMxsI3BNUaqT04nSaI6qImIGCSOekdMLX0dApkLBSO
C5z8H+r1LoJWZjPajzIkD5W/0sHAcq6X0WjVdR+uFLS3gcU5wHkTex+6HRkWIVlr
ILM0knwfZ4Ghzkj9MFeV9b4UhgLlofbYwkstiPnp5JCtN6frHF/ZLwLSoFF79EKl
zrCHutBu5Wt/t9tMMDyzfHJD1irsonYbnvmV6e5vkMLG0yE/GPCy0Hq2FhLNHBrN
3dfpy1T3b5vQw+uDRO9P4QW6/GlXxDiHF6m8Hi6XYrOLYhk5JSQ54lXws+Qs28iV
0PUQVv8+v89PZl8EgiikMWroauWNd+bVFcVFQTWJ4b3kFrN6spEufcaDDnveJOg5
XuAbUTsM58Rz4aVLB6cFVTPxGPXvD5zHZ/i++u06rLUoZyutcMgZnpRf79/H+Dva
SqRaT7V5PqP9WbzVMTR6ovDavbFYmsf9TzEeBTwTSJVEnQ861G5u34p11FYLerEf
E+KY2uf2lq9lQW/0G4ozXVdC+Q/FGdTVpjTYegcNJpv7/CmYR8WVHx4W9JllVCgv
8vQD2yLdnurnYKuCl9Dosaf6efxzU0FJXP8pbEn1aE6rOHPqZSTq1kk4ZgXqaW+d
6be/le64OfmTLLfZSHjE+yOvGaafpTlpUx6Js5KpVMeNHN1GbU6PuWSj/RQoVxQ/
noGTLEBAULd62xg2QOwlkc7s10sPKS58YvqPKEgO/9voB50CDlnUnVOtpvi+zjIV
hc2HvQjFF8eqhrc6TwQbZ5YGjG9MzUAJosnTkPmQduCVGNt7IKQLhwWUlbDpgHQg
5jA7fqTGb5uBAOn2h2v7dxhm8I067XNzJyw6lcQvYTJlzqfn/tHqGDIQP7V/OfgK
OhTXL53uc0ZuK92y0VAQGa97wOjRbWGjazpql5zKTd5tnozmOsnxWbXnT1/WX4Vk
9Tr9YkPFxpj0vgbOZk5cK7bqoX4hWTF1YmIPL8Uf8X1+BAPADC82UuSTtpo82sup
dTK+q+cmakJCD6olyV9CUERDFJJwysiq4lmh85OMX7fz3a+12IRUdisXI9zGUcvi
No6qut9qolmrNvvkO/vGtNC0g94fRhvEfuw/TnXyoBpzBHzkmtPea/xppaNTZ7g1
J3hD52EKVhlumfWZccKPh6TUO6gw1uWYlTwzvpKRn59Zm36qJSYHxadiDsqnkfMv
GSmUNF03q1oqQw6xCoGsTV1aci7EFdPiIxqCqU2iQXlNsqF6mjlB1tF+8AqoigwO
jiKMWQ8kRcXP2sZE1EEnS0URI1SWwtNEWOHkSdWjAR4C7jNpM7gxkpFtEA0VBgea
Ii1LGAAbVvYi1iN+vDuhguVqMsESwBsQsgvtuI60mQCHj3Fz5EcSePaZCQvelZR3
IVvuO3OAKyRQDWb4aV2svMBo1GavwdAKIbZcRRWmvRkOCU4BOkalJ5uhTYgxsu5v
id2WJw9ROB3XiiQ0fp4g0+7pYJm+TSN2ic8X7S3fw5tjii4MmKfU8rMUVHEbv/Uf
Zo6qidkrtAdsCpJ+j4wNWC0xJ2Zv29fUmYaqXhCHE+i9tQvJG3tT3VZ/LmoZZYII
tfulYQl9xra6fuWu0yFn4y8z3Q17aI9uTk//VEjDHrNnAVlCrX5+yq1fs3V87eYQ
XgOBdber+6objguwcuXiHoayU6ASGNz1uj40quEd0Lmj1y8jQYcs275b8qabHeha
/9qLBnRmA22USHO8lLAxzT7TCz9U1iU6x37KDdgPo/iIRUwZt3gUpdLKwnMp+5X1
G3unboLlQseUU7OUJXwgnyr9x9zNWGmbyvwFuLg6wLUFBTgdx5co8uCkYzz273TL
LQ0/2xIYCJG6miqj9+CE1GM3Gu0xPnD/bKgM9XnaXyAKyRzjyIVWE3Ic0CklXFh/
c7m3qz/mbEpR3yBPyM0qtOC5NqEJyq+I5mblrTV5Ipf18FH0jGFisK0Bc2yuSoVi
oQaRixclSI8b4EIf+h7jOW+x7LI3UJpg0zhU3MnPDrLwwKYT5G21s/PXCMA/Te4e
91kzTCWWlxs/t+pmZB3GLmiFOJBbAnPBeOIyRF0E2+ouY1NgUb2viT0OT+Sh65tg
gCVW7weJuaY1Yo6qS41n8Rjmai1vHo4B1GHWiOu+4/fdNexwE9BsIC77JVDxD1tI
sVKNRp+pOObSrClKb8hxA/hue4cauFQAYlyubW37Qoo7fAWS7HtSQfVIJp8ps+DJ
+4cQO6eJA9wlBB+8yVpC2kMjecLwoV6N4vPVmY/s9weGdn12sTf1QZjZz8oezJQw
xEXMZae/lck7lyGhy5pEvsiYaEiBN5vdhK5fbIbJRQVY3iNAklp+jMmIApJ0jLeW
fA52Nftsx69K7qp6Q6L5MT1lS3qoXU59oUngb0ZbVsNCzvimlY2AdD2Ja5wR43+W
8opybaDrPP9CD0lls7mRBu2HTfujCj9BVM5ikmMD9wB15e9SZGyoJxFkBdYa6eFY
KuzzgwSsasStEROTJLuLQUJQU0rWejgI5p36gZE0pmsr8KbjYlUceu0G9UqOYWf4
WlozMXgz28v9NaftEX6o+O5J9pGPVKMXXfDdMoEFJao8+MTKkFaPjMp/14nxhrvu
vBnEiO5G4aDcCH7ebaJSPSOngJtebY0rkuhD3F3wDyz0i9RnF52+F7GC406cg1y6
QYSHNK95lSNp1ubtJ4SL4n4DIiZD+d2g9j6l2/Py5m1Ac6EqNTtVFqhkUVjqZ4Oz
K2Un1I9Vpd59hafzmeOfgV8irESbwYDsJSWsLdzLSOviZU9EJJXmkxakb+lnnHZv
z4Jehz8rKEsrTCG8VX1aK3aAioLnmVare6XctgBJaM8dN/rwYu/aZ3LcgyAICQde
HYW/zw4d45hw5J3ZW7RUimqmRN9ZdlXbCZ1x+XWCu6HkRkvSQiu+XwjjioLHu4Bo
wyLJrr4J55CYSSTz74IuiWBwg8xmfFGaG+DpKv3pD9Q6FO3ljny7y0gy6UAIl5km
vSFsa8YokYt2Y7a2/bCnqIg1NnjZ+jXDs+1VK2IiP85eN0EvGP5AlKAkfyBx+iVG
70bnFL7XEFWWxVIgYcsISPcuq5CKUPJzQ17AQRV75PBS9dIcSrIrBVpe3w5/SGxj
R6AckmZ6CoDqNE4SV4tBUtf1NjEkuPJHHuOHPLJcYIBIXAJwoZ7YxI0UHed3Dp1a
IGW7iCLwLfNqS+hHyfHhJ1aFOWxhZ+xSiBzQ9YyUdx0EAEZs6jwFh1Av5F7/Z8SX
geZB2PKwKbwWhVOTD8kepc+C/OVcuP2G+VqVpsVtSrdfT3xhrSKp7uYPpwOi99Zk
3JfyTLIaoL/Y0k/kpq2Sz4ypPAWBjFJmAHt3h/RKCr/Vw2anE12KgozXrtleX7O4
ovyq+lH6d9S+Q0KQMrVrt+BZ1cz8NyMff5Bu8wB3s2NFEjXOJ8g3F/0+0gzciUhs
mhKf+uAra5p1XUoRruDxfwrYFYBjMCJdwFs3I4VeX7Dwtrmtu7WLVqi93fKSnVDe
9u1bGdQGtdLgxz/FlmITUltw7mZWf8Nagi4nCw4H6oO46+ZqbVVfcrrrAKoMYfrh
sVlTbdr5DzfG8sowN47GdMNDUf4zpUjV8ioiamB27Go0/Z9zXahWzEb7HzT0zxim
YUbqs0XGgjrAd2qp5GgIhewYkAVfHkuq3lziaiB2ftxqdd5cnSXah/j5Sp62aGFs
Njv7MIsfWltrk3fxg8KWLHM86xNBw8eJ3QwFkGGIxoOHzdO+NwXCfjyjAw9T+Qdk
0CLCi1CvqLOrIvCZ51ZrH8JJiCq4w0qByKHzki08hNYkt89e9UyRsZkvreNfa126
Mp2orrw8a8PnSQdmzSB9YLUdh7PNK9yVne+ppTfNOClZMRpXmmLtUZldNayzRN3J
B44t4shF7bc7vs+BXoh5z5yJXNOf49awBzbgnPYdhSx7aeYYNM9lIT6srK4oCY88
jc5tQCuW20H3cN4INO41ZD6Y8tHMtX+aW2ALApl09nToZWYmmWemOamlwbLOivnC
CwcVBORiXPCMuRtah9bxQy+/2GwMuWJRe1f6cRphERjfMc1OrP7vuUr3a7+Nba2t
c5+Pm6YbKhjJXFigJKItEK3kv7NGZeP6fG+TEXiZ7qqO9hkMrMpo5CBFIaKVZTxG
+zdhZWEXF4Za3jMaLOkAtGU7yCbtkTVgCUSIyf7OPjOR6FNIZ7fscCgB3zbSuX4t
BOIfH5daDz9BHRDAojAYTpRSFQM8DMehSp3Fqqv3YGDY+EZv/5TLyMk4RZUPKnza
YgjUDEjUY7V0/LVYIoCT7k+3rUQz8gsVSDLqWb+0AFm+WqvwQvNpXluYRisuE3DO
jZH7q8AlQbj4xfSNzwCMhX35EhQUg54yjnEY7ymF9bPoo+m9lYWhebWi7KIPQ1YM
qe/hUZln8qDNj8VzE2JJdT9ujLvShYthVw8LjLds6P6BriioK6iVv/8PPkYvZovg
0ZKvFIIbdwdrcEerIy+G0UjR4yhcYKXAzNJ0rxQj2xYzs0er6BnnhygqmRPqSCbY
YBPkb5kEt1jXHAryo2cwIOORjzs00Kn9nqjHNMmhY5v5vT21SsDkBDBcxgN9+HR4
vyfRQfjwIxYMbIlSvMcA8C66/ADOV19gPm6u6z/b61rXxoaxKcdlWi4v76VPpVKc
9i6OtxbIqpeSqFvWUNx8i29A/l0KWWJfR7LavP5utYfSC94/zbLPV93m2NYHRYAc
DKPF8PM3AARnZVI0Celb/leVzPE6wCr+Fld7OLPdOgdqcAhqhDcVmEraR9SvNQ6R
Dd/30tltrymyvELP8odZ9YW87jXfv3/m63dRGvqXVKkoDBDdPxtMWz6I3VuWaLEk
qgQmSL7X2IuRtNerqdRtE9DAd1zzdqxOXQuMlqhdCn/NUn73+7vhkRUu5IsThWem
aIJu5jJPNrd3JAp/DA2spDS9rBaLgGUYliTbE+IMIalX7FVXamLiO3DOoVFVkdhj
tvDeDy/D85KQFMWFisD2bnMBh17JY3y84zPFZ3sCrCRA98zK4RS5xoBcSuxcsZT3
Qu/ixbZ31+/zVcdhvJEU5GP6AmQ9VvCWdVknmV6p+bIwmc/zfbO7CBZGcAjxOB4H
IewAOv9Z+pTZmM8ui9DCj8rFh3WpPvQZfx3Kucu4SNXDnxGIsUFO2hT9kcxxcY5V
NJWPiHJXBMNzDMV5H1sg2Hsdq+MgnWS46dGD8Rcs2zHleuvzHvyFwd2UgI3c7j7P
dg1HCW1f1in/H+rGJR2Z4IMSrxG/U7A0OgVCA2dAj9/ayAT96W9qREYMCbfvLOmo
`protect end_protected