`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5040 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
mvOv0qUqD+6HYGQ6UGdqrcy427utF8vr6qxaZgmhWKDKwvstoMYqBgmiydW9Fkz3
LAXfOWJIwxDN6T9BcVXQuc7yEM76oyNsFwny3JnUgVDxPOcmCtIz3OadmK4hOoek
FmRWiQZ+JQ+NB/TyQQGC6QF4FoJWYb+ymI6VlF4W2vhQhsb3rDl1Px/ozGWtjXsw
jFiVX2GEigndJmnjt1ztUSM+XVkPhpXhV8M4cKCAoNj+foPf6n65PCA/biC+1X2r
0LCmrKDUiYfVC5xIiJMq7IOqdya4zuVxmfGXzhPPK8OnIKMuIRH7IbeK+c4DZ+zO
+iGz+QiKsHQGsU69uRROwRu+c1WCjWt/FMaqAGQpEuv40kSu65PJb7SlIacn6m1I
Xitq5FZ0qC2lE+W6BJUPI8K2DyNhyU0RkTHmzFnN+fCSUvD+poSpnAxmz5osSArN
iLJxvYm9hq0EnMI8UQqet85pG46WcRIZtSbBiQXs9ByW6ndQgeOcvo5+LnQXfXGY
J1PjlHpFECUz1XWsp8dzgsItwZasWycZmyvEsvPYRlvk5KPWBY1mqUbuyjq6p50u
WqeoE+ZNt1+7Fc/CE+FNo4FhdGuF5SrQTcPFpJc6mgw47oMen51qipqcOi1KDsVI
Hk/QyDBue7CXBgflKLS5hkltq5b37LEpRSvvw0ntjOP8FHVIs4yuXmWGiLcdz+rx
18xzRcbS7cPekBEXVl0o0ErxMY1Ib2F4jml9Dnnjdj8d9q5YVbPDlVaEBG0RW7q/
hFegQ+50ar1oRIn+bafz/ZHPVbdkjP9B73ka9nzWxdHJhx3YQ+RCIHFsdQ4KwF2V
v31BBbc2Zc055H9R0xhXIXz3MiqnL9vbw3/pMt6dSgCwzaXP8K3hC0tqDzQbYawp
aiCYeekjZ6AqvD0XrObfDgtuV4eQufGCmSTT53sDfMAvY2knoOa/ejDzv3MbvCrj
YFvOjCju7Qpd0zswWAzWp+/YN48Trfv8P4pXZIYRKt81C7G46tKv/Y4Yre1ArfyG
sDWprSTRaqtG5Dgw2O/csiHE1qXXL3lmtMYTkCZo+X/aibAsa4HJJxVyo3P9X8Qa
37T+Y+Tn9eeIPDF6PGMBoZGUfjoMzhE157SvlsSA7Sx4mbYmc2kR5m7ikZitsV71
gi6cFrQSA4n3Yo7ItXcQBhYG8Gkgbz+R9RPp2pm77Zb7BJd+3l1iqy/kw9sLB4Ls
H70RcYjJ5gRLuH9YxsnxoRit7vnnkoWtCuT/NWJKxpirCCZUBHRgFsdTV6XHY3fS
Zp4tnoO6iO7dSzKWHv9ys0JVU3VGFiAu8KZ+uuDoWvlTWwi2vSbwM4st8RwacZ5d
VRjKU2ZF+D1EEweDCFh2MsJPu/wU/rT/XRL26MfJlDTr1NLpFKL/6UdI7pftMa4A
XyU1qVrkPf4ra0Kusf5xz3Bpk225vmWZSokXbVKv4GnuswxGhjV1l+cXcoM/WFwE
BbM6Oc3OOD3MrQz8u5i6rTUJyox34FnrsP45M6py+Yud0Md1CjHNMmtuhrxkItsB
6r7+oL03o0gumaCLR3EZzuBrlFngIsY3TLrDMIeMs22blEM5ikPwkrmyFxyEFY2+
1qKOiRPxIXd3LOF+yJ++heE5md4qjjxlzz3j6TA6Ym0tj+P9IMtWQo/lR7oc+ZfJ
ADAIAGmh1zhUKZPs/gJZER3g/TN0dEXqg/A+ursKE+ewBrhEDd9WZDsgVmBNY4VM
BFA9y1VOayYx253Pqfy3k/sVZWMhQGffAfUojAIvfU9cRKzCyHOxXWtzsx1ZG+Di
AMVDLNSELWZzmBhWCLFM/lk9p7W3GbCIIMjQEjmh2xVUqhNvdnYWcNgIPHkrAd4p
SnHfrGwWzd3cCSchnql+TaGhVI0iak/vqdEyDgp/bfOVtlr0EbX9kiF/HQ+2E9Yg
6EV0MWLNfrukNgssTSjH0oanMP5rYIya/hJShvK7hgS6slM1voncezCflD20ei03
olR2c2uDtmKuS6+KbhV+6Wq8EbTgBEtFXh1jREYoLl4B4uV80STglOWvQCjGDPpT
W41e/cANZjTXujweF9xB9v3Q3YgjZdtPeV4XnKwEuuEFZwmMxF2MxJDzNX3XA2tR
UlEtip36FycFE6DOZWwMOVEDWDHLHUoZ7hUoHVt7rhDcNgR3iGCA8CdfjEwVQZGM
UTCN+uydLbMkyXAA+Vxz55eEl9iQf6Innqj3zOSbyp4QPpv26x2PqSvdkXguhuXQ
Y1YJoFmkE/ZRzC6Pl7RWGoZOjweHnsygl9u00cKJcvUsac7BIyxn/3GrNcdO1Bkv
Mn6G1dbrRebM2QslmRguoAXQNJfsjcYPtxqE1BBqM2oluN2Dt0nIx5L8a1JsaygW
2ZB0k+/zUjSk/Axco1BLACI6Peidoo/XfM2JBVPACOXhB5sL6+pBVNHK+SBH1UFo
Ua+LIVDNwfH49kgnVsiZM0ZHMXYTAeugSyAJ6xbaXrbBpwUZbnZLr01ZdGmndlTZ
GfwSYgNybuCv1rzIu9f8S/rXAZQZEH6EOcs2Yj71xPmDmTmL62pE/obGWHg6s0Ca
gDEs6+1cqlL/91UwvLeJ+jvyBfxOCRrmdaUGYKCoDJaA/RUw+UhFKGkniwRkhD4h
ykDy6h0FSQkz60XZ1hl4LncphKkB1AGtpo/1p1u5oJE70nxRmZlK3ztUG21KBX2W
V7xbeKwhoBy4ftk+S2DpqvpDM6wRL8CWQMziLH9hQUKBPu20pn0x8R6RvWi6QJXJ
qaNK1WzNcW/vIkf8tdAq3YeDIOqhh6EMp51RWMnS2bJp2laROP7AIhlM7RXcwutQ
kY/o5iwunKqdlVLFgXwtU4cPF5mi50toCeA+f3WKtQRJyeUnTBsD7k/Nq0mnyjib
y16W9tHqK38dzMEJelEL/JjrmJcrzRl/J7CuGhy3gLchldhPAmxAbMCdZAI8tsAH
r4chlI8gpaxxVx8QAtj7Kn4MUP2EeiKp56i6Nzli42s6Y+wcEZKDpsdrwudTTZWL
tzg4BXxZtFeHhcWR2l0iWt6TlS2LbLFoLeFUYGoHY7pHKeFkMIwRhQHSuiskmbwv
FgKYlgQTPg3auHfXlmqhmP7yhj72PByaC/3PtbOD3vSQUNeF86T7cB7crDdaMVm6
mGlhPyt+JmPyOGSK/NEvSMrXBElMPIsOA2vyOmOjdmMTAiq9/dEFu7fG4knua0BB
ilavTG3iNjpXNG0Oc1BsUSwYoG+blXh8LeS78mczAqwBQzcfOEFGE6/CjNqaU5NM
zrzBmGQIw7XIzunsq7/eUjpxM4J0oVnN09uVy7tKxBmlSjxCHtzUl5Vsue7np+MY
HWSef7nABRKkzvbbfEd0nneHyH5dj3ZI3yg84zVYFAXjN1+wcd1AJJxQ65adaxjm
d8IUYjhRgGjEvQSiJ8HlaOBawnnGkLRTQOHo6aSvMuWqIcdVAKrPBH9abl/91Q9s
LdrOesf61FA12eawBwsYkQdY6oafuY0f/EclWLvBjCe9flmMrgonNjirAJSRbW8t
mjXstHAonainARKsqkl4gl5OhLdcoqXn2sKf4UPx1aYZmn1ZHMymfNKsEDEv3TF3
S1EPub/h3uNXe7WkuGdR02kLcqROM7pKeIvcXlFdokhoWDSODwS8GA84t+xiSZGL
8Y/XWJC3byJf9/BTFCc2PMCIde1d4kW2dPy9yH3JSYAXsRskLSkbhTMXmXI5S3iz
cVd6I+dLX4e7oWMQ+L89c75oiOLqMxw+JG2h8TCHy28ouyRjx0wJA/kjqi0NS0JP
sqITdTJNf8+elxrkL8byjvbBwvlB3tWHYwlArKzdnWi6DOq5PNZk2zDrDodJc56P
MQ8yMvspvv8mA9cZ+45dUnxiZCRv2OfUwxrFsrxetonyg3bpeCcqkkcGAaYhs11T
AEIdDTOsV7pwjYcQHOE3z2eQT6MVaMYbnlZSZkA9umNNXb3zwlslE8d2+DDKzpii
f8vUrmD0aZyXIIabuIUma52jix7ViSmdUykxNIVTPRbufm2yadrw+zqSvKKONG5/
E+YNtxTXHePWI0WM/l6cLBGjTtGUmqFCc/LyGWXVbc7OsBCmu6ZuF5IQgErNPc/U
gmVzd1chKw8r+Gy9hINPvqo1zhP9lRWdG8xkThGv+2qs/9bxUdtX5nvnWvCfGEJF
syJJxIat90xknA0y9PYzaHPUOLr98Ed7zDPTBXsWOTDi+NsF7H1u3Stb1nvA9CDQ
nNoROsT2yA/k8N6d2yYaNFS1H5Xs1lKwD2feMsU5Xm5Xu3MPS08xlHY26Chq5KBU
7z+VU7B8YXqL+xS6MsTznSJMZqCjV/SLvkeHcgkk8CQXWSNFEoQxsmkUaWPtRdaW
4W3VMz0fSAAaR4chwFQU7KK8NW8IV0TU761OFvYfy4XaBPJcvV1nEkkWUxz29c2V
sKhGv5sBk3EEXDJ06NICI3RZ0Nw5sDcCnP8+5Lg0ZOUuQoFfmGblQlDsVlUrqwAt
7HVeDP30w7bAkSk0AVgYkAl2Rr3dJ66YyAJ3NL99rHjcHuViKBpJ9+yVOFpCl3i6
IwcwRMw5dlnfztL3Zfg/cVMl3PQkOEoBEQ/cj1pHLoQOO6A1N9MYrE8Pkui/Z5wX
KrM/EFl6wZrHX2yRGfS5169RuhZxtmE+rDIa1OIQg/ZgSAQsXjZ1bs5KvkOiglCk
M9V7oZaObe1H4ZeTI7bPOobODIE0otgm5eDJwYvDO16DcPyMXD2ZgjVSWaZvK7jq
KCTol3MoGAU2Ihj1DPGaLmJ3+4EvZ8Bm/e+uNx6VAPwj/9poUCojWD3jbU79S+ce
nyJzbVT/TpRqz80+KXT9skgvyRz2Urf9EUd6hSZYjKIxH5HrpSIF+faE6PJJcKYE
fxlY3Hek+CBG5B62C5O9sxX1B6FUFya4CLZPpU38bPpoiKp3G1XdA/gcx+o1AsqY
q49g2G9HjKE1LSY8MpmgNFbsF0Aql2Pf87/k7zYiI65r5hWGwFZtWUpYbmLDoAng
nDxr/XluVKUop0AN/KCf/lAK0DTAolRkMBcFFzU2Qq8xXvNc0MIU+buGG/OfLqZf
XqDwlw6XT57DahBU5BMi06Bgi6jwVLLBaQRBr/TPRWdMf5Ll0l1AVZcdk5RwOyJw
iEjG4HErzZLXc6DrIqZR2UZ6k9XU+Q7fI4+rK6K4VRrVH4TvfV3WVHWBnaz4BGlt
AVcg5HolwuM6PoWtL2GZlExArjGRuJhIfTV5U5hYCWv1x/OQvgcupqJHFkiY+XAw
UM4Ur2N+BSuYVJ/o0V6XfPoIV6OfaCwLj+IkQ0DKqRrYOGg9jkzzmai+lTYpauAv
aJQGjtng/GDFjLdEpqNkiheBr+bpOoYltd4hYm2LEXFeBhEsySYEA465yCHcBOqo
vYOfbSfE9fl1FPvZjYffUe18ti1HPolQrd0/bcA6uKxgOhSq/6V9CDBywMJby5Cf
ffhea3SQkuBY0TAkcUBWQMRDsg+dOVcL2MnfLp+HVMDtC+pNJN46AwSpyeS31iCY
LLwiNvod7/9SEqRnQXSOJJ2XjCZf7XpAR8G3IyaDAg+/TSqEPTjHZQtixqnWsYSf
y6Fzp1hM3nlIchlrS8UAASsqv9oy6EHaUr72TXzuPy1YwaFItr+tGDo3XE3c4+7s
5vThw39ywyuSaOjMP/eOAYJJY94cAtv19fgu6VrAse5RgnHJYUeoKq7vRoPquSjV
uG+5OXARyuWqE/Hpguf5T456gq1wKT7+EeY4gDhYsliCK1XyHQaKGCqs8Qxoo2j7
FRsjcqoe3PX94kwyYfr1wuC9/Gkxn+ShzlhTMFViFWPxaNBaUIv5s2Dw3bJIHopc
5IMYPf4wZanpXK+QGvwWp74h7ciTpDeu1OjcW6zd6e/icbNGykAFMACBRRzBWSIS
KtHcNGG9KDOtxnGfgqHVZAPUZNtTQeEDElIwXAsBitxb+oVZcS37vxcSJ52uYWpp
HfR9YP7MRIy4JX8OasnBySbAIkSxN2O/dJoGxzNz2TnVA7XNSkhX9/6Yr165ANep
SlofoOoK8enCiPlrPqI24QZbfhebKKzwxxhQ7rKAdKvLQqKnb94Eu/Ux+epXgGh9
IxEhnjHQ7lrRTJWsWNRlGgEQs8m+UkJ6YR6SVYhz2JBKr/t9TC1PQqP3bUDqwmnE
oTj7qxd/Oh8XQacAH5Hy/Ji7mYtB7AsoqcCcCywtRfOT6fSFdRnUH6NXczMc4L4k
yMgB9UFxDZEJfwrjX9TxOoMun1yXdp2nvM5EOMyseBoAYNb9RPLq2hSTV1kGvNyq
TTspaHx/t06LNu7xg5cwwo2l1xRbxQHAb6cep8emtc8c+hjLWUbHTpHoTqLJEg12
VoizM9siRxXH8wL5xQM7s08fTlUmXXvWj7WnIFd+8CLbmiuJ2PQ2hbGGkuCKe+lT
ue9p8UbJtp5XxiqPtuzf2JsPTpitjm1brBBMFQB3g/V/ItAfHYiQMIyJ7JTc+DUS
rOhxFCoRXtuXE8CkL3zMlkbdXePheRMlLwu+FJmYoQJHS5gjU8n6CCdzHvWsEHjq
f+eGcCLEcQ4kVOqYWxkaQaXGZ1Xkc87b9tjHzIScK8BkcMU/A7tcRPbBtXWmEPCW
`protect end_protected