`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
0DfQnd5hIAXb2OPobVGJo+z+/IbfxvW8dMGIcptpCG4dKziowNKU4uGneXQOi+sK
xEaoc7WDcegBHnt3ogGBgnLMWf5jN0yWRVyCGxIgsO6+HyVEJugybJNPuTy/R/zR
WaTKYtpriHgLEi9V9Yvw7YNlsZvPgt5PkblFexJGudR5PzUMRie/LGEhYalYCLCe
h27q91C+OhRTpW0FITnXRbrOc7kEc4jO5PV2mIt//vOCWGCOkP+1/alExhRHdMWh
Fs8ofQVy69v3iW/jOvXcG2RHoowPb5M+5GOBinVYiUZ72lSAFzVYDwrezo06dPIq
XlMRJIkzgo3Yyotl5sv0wF9upved0GB0ojPj4vXeGCZpt97Ieqp46fF0xIhOQQWU
HVKr007lW0nffUAnQc8Bd+xtAbCvWPSR6+IxJ2F9JO9PfM5lndi754sKiOUQ7RkC
XPy/shal/TWtfyRXWQom+fq7WU12YYKvJ7x32UmVE8JQeOe6Csf9lMizNPRX9oQa
LYzkNlOMEVg/L8vkRgeIvcEQO9JCg9xMC9x2hu8ropMfL0NLChf0xG6BzCXCzuWd
HG+zTHyfdINZ5qiX6et2qkAZ+TJNdqmhP4BnXC43wLu3yR3m6xWNnQNxl8oIjmUp
j+xhG8pivV9QIBEs1M1HfMIos3CQbGG8MROZiXZAP4fgT9OU9UXXwQetSyndeUAn
40m9PPwoyufCTiuhL1VCtWHZ4myqWCPUhqvaUCFUuG0coiDk8hrzau1PkGeYwKR8
OVElPK71SXuXKlxEnDU8UbCWm9Xf5daAZQbV15ZQzguIUP+6++VhxJNJNsUYn4IM
AEzW5HKlE8OL6yRr29MnadWJMyDfA5lhFPWcgLkuxP/zpvdi6jrp+e6gG0vZ+VQz
4Tyo9OEKTmraqlh8J40XRLfTfWHbMic1X81VL7N4hlY1Xtr2A1pIxfg419yXSjDz
bFj3Bh5XI2Q71yUn4Xd1/rziTY+PqZfmL8MxtBF9zyTN+mtEIpDOLqruhS4h5Lk2
3Ot6JCEvJn5cuhLtrHCD8GNmn//OLr5V21kbcaU4j+DSlFtHbR5TtFSaKrVcOxJK
hbL+7QQxMNBIPrIhEF3UY88Wl4324omPaVV0crPMDzykHsdkv9/lFEdIU7LHbMLu
paIcrQhLxXrYlVtQjAZRXTT4vEbFCmEp1z0xjuVUV96JEpljDZQzV1HPuLyi/utK
kTHzVw7S0z1JiY8ngklnCmGIQ/JSNM014l4H6iVhATRGRtn8qh1NCCUyMNDld0Wr
2j/AKlCE17GiPYenXk4gv5s/Ob80xmsr6Qx7vLc+T0fmbzVg59MzrWuUsF2rfog6
dDxzVcbJqPG4n6oHv+wXxWHvxLJ9ht8tH25j/QMLKB3B/0Dbwi6qQBPyjW9FtB7I
BL55v4lqWVJzkL7tEyk5CTn8ILerG9xncqA1sdyqIHLcz8/KymdnG8PMpomB8gqB
kfO7A21bmCxzESJBydKRe1oFwNLB9qtSkyEP1AfVJbO6IGLstZRc1bo3DYYjrAO0
XqRmsxW8fUpz01c+eTvy9LIzaYZNrrV4UWM/gLR03uiKIUNtOFvsJT/z7AGYV+4Q
vcqY6baxnquYwjfc6AkjjjgOA5FjdpuL2m+yDlRgw+ocrmLEbyd9loP1WHBIpQ+n
7ANev81+aCAV1lqXSssvYS5bfKldPE5sfq1Iu9gs7jKprGQ/yFAEO6LL5drAoRur
EXp4OKjEvUGaBYEWvqcLXR0s5psdNSta0OaGkLt5eXiq7gNhFkZjqmIusmsZztMM
cmgqYBZq1aLvgilFMfB6FAs2IdJQGjbQAjkNkLTBw5vDi+I2zEHkIdlDQVsLY4Pu
WuZNgTR+d/VuehRrsPffjdj6xEUDohH4VC3PHku01lTEDVG9Go5r+SdwVZeel0gh
xIUak87NxDdvCIN+CX0wUz4vyx0ZBExsjgNx033u9DUdGwi9GzOQjHcK3FymUbjj
rpc9JghTUlU+JUTYACE/5Cv9xBEXpnRg3v0gP5zuO7ElbawCEnWx4JrHcZoitQTR
h2gcOYz9xgXK644VRL75y+lA/G1/xP6Hml0m++RS8MMA6QRDphXrDreAsUTVKC3b
SB2LyyXxftbXUz0rXW/JkOUKaMueIKhA6hK3TuEWvneJQewVDACF6q2QfpusGi8D
+85EktpKhD7L3yBuRmVbZ27ZXuoYTC20aKFSTBPChteziMLup9pddvuYgiqpdtvA
CPGMF3kqchkiHPF1VfrNPTEMMofbwst2urXDN+rRaAMEHTx2Z9jBgqhrvEPltprm
UU+mky1z8/rSLwiU9q/tMa6qecmJzd4v+pSvH+TX06Dw2G4jtj7G/HF/tACe8ad2
HlAXAS/welBlcM3DJc+ZjRQ9/wYkHqjBVWurgvnQ67X/+z/amJbIzPbn28jhgFEi
rGpXuvsU6it1k+5hz5yytBh6RvybVR18A6SYiD5bO/b/c7frB4YqG9jfEFi9nLV8
YJKGmh0U57QOALac2N0lLZJXKKnIvASFNkzLKS6ZWLnpW+Ri2Lap0IosGk/PmQqv
BgdcLO6gjmsu06jZxMuPoPO/57RecAZBJd+stKJU/bXp005M//QNDhv7FfmnC46H
52P/A/jkhfvjoe6m5L5zBveLaLUqbqdbLYrbE5abxmvFTFSQE6ii0TMMkiCwGonp
UXRRKylT1bPrNDC8UTWL785Ai2DHLLgYosHOxTzRMcq05RsxFnE8Yi4E57C8I1aD
vy6A9ysw+60f4A0qnRwkkl2fYdlSLkjarc/ZVcNGyHi/wphr6a3YQGwZW2ftKSbe
QOdR7ab34aA6xd/deNZ3FqSu8xRyePwd89XkXAGfbj/ZKVeIEI+QnTwRfFOn1GzO
fA5RIoP9TvU4lOiPkY/H5NTknW8LQBEWMkzdfUzY8OqJkromWQ01f3b1JCXI6LT+
TNgFD+QDlfnMGleWqGxFaHfgWP/htP95/QFDvtG0bLddPnIuCjqikOnhKvL7bOE1
2MCjfzurGiUSwaPtoxWlsQ0iF3DjQIHgwAdSxUt4CqX6hwbVZv67KFSNOMS08t+/
xY1X8w3QZM4uTz4NYxyzH27K4gDTvQvG5HukDqCOHBsSlLlax6ax/nW0tPjn0eqB
USJ/HY/R0/0lyOsE++KUVfi0dmpj3Hz8eLiW8eiO9offGO0wsW7FT3hRk/tyy0F8
3KSM4gwOStuzvIgVtldpHLMMU9WOns8NZBCDirrwHgJ7XY/1b1r+fRPF3l6m74SD
0ylklfj5OxiDMEzPfoYW3+0lthsM+4MsbwlfLbscsyzQzjeZSFE+bnGmYW2DTEA/
4qAO7tXrGGPmEZcrOGuJ83sX5VjgjW4X26VsnI9IyMvRW5B563EQEKIBnk5g84eA
dP4zwcr3oKGpWlUlEQ8gwBLVEImKk1LXmN9ZnmYSmkVHDID6/k/bFRGP994nRo+X
lIO0GIHwWeg1tfTqiUjxU5ML7eOA8uBsv81BNs2nkog65p7lmvTzd6y9MtmeWQ0Q
SJVbg++mK09eqABrY4p7md1llcCEUNQOEQIWcXPRzgRzwe6ceFsg2oM80bUebquH
FMlew5Hh3xW5gd0ydRe6ls6dQ06ejCdepTBJcCdezVBPnH/H8F0W2fmFMwXNBUs2
ruwpnbgeMV01kD/KqDvWuTDzFeAgu9J+d6WkdcJQW/XYlf17aSfzzpBdaETf6LiQ
2jKQb980UnOaBPFCLE4Ow2c6VNu/YpEHwOTLMbQIr8ZEE0vCtqIPTZQVF14Ogi75
P+XKa6ny+M55dmxTFHhBZcfsCaeTaX5wh/G7nNImNEsZSi1edMWwume5CVNuhEK2
dDiy8wt106AiVAWk3TOTAkYxcG3jnGSa3Wg2Jjga+aY+YOaB0slPKAw2G9wcioIP
PaCyPtkWI8p3VHW+3xuVYRzfcHqnpiPTzD6jXOaTfp0TzME/RO+P5/reP1NWpQnU
tCT6TT0YvRKr/1X+J5FmxOTTSRJ8EPQ7VZUfTm2EWXmELfmE4IvV/xUXRDpKjm4s
xqVrbK3ape/P6rdBPuTO+juViCXdNgB9mU+bCMJ59GFzafEsRDsXRrvqoDky7QNp
6l4jadCbWkJsbDiREjfFnXtdy98fH/bfPLUVet6zgg28JH3cwjukGxtvmV6MDZbr
ORTcMkNC0rEyYOP+iGRQ/aO04CamZtw7SXSgQMpnQzIQwRY+QxM4HlAUXjAPOI36
NGWVHnDip0pnSwfbEEbQNrBmZagyl31DuE8qZ8e69eHdBbzT4pheyEkDPTxA5nlI
V8ijT3UFhN1Y9aSmO7OhHNY9IO5x5KXqoT63AOUNn1XsK9M+vfk941kcBRF92SNE
6AM3ZUfJEzmxi3HkiSpjnyYnw66YnzEhz/uKtZvlY0xKQIaAoraXqJtbfCh15kED
09ariz7zesoxapWzoYvhz7SbKdllvhU3cXzbAAg2cTo1L/D4iLp9EFB987oi9/hy
nR+WZVtnTikho1OLypgkqYx/zFaRyXLbprnnvPLQseoGT2c1J6dMBfvxlA+Ylfa5
48MtuMQi35FBrS9Hzs2OvjYuUSf9iTC6kPrYRAmroMPcZAtGKS4MNqVVrMDcGxQW
fOw9osCptpC/PfkFzO625h7amr+LF94ytkKlxJ/CIVK3TJ6SiEhIk25GsQWVZfVu
8eXVH7oAb08D5JhV6XS21dIxwtEMr+J/eRvuHyQmlu97wt84qo19siHbjc4EyeI+
omZwSgULhRDWbgvhECg5sFTxRLtjquaTEEmdEadgzQRexkAzYzMFv2VaKvqKV6CS
UaxT8AafYlhB8MS1OVhh8ulFwjDcX719hYxk3aqJWUAUoxge8vuSZA4f+gMOf36x
9lUN+B+sP6by/XclTSjyTehu/tyxuXv42xl/eOS064JcWEOsEkrIsI8sco5PcHqI
h57dxYl6Ct91K+vluTF0D4fgDTI0L6/iwlzq+JzDbprD5Hs0Kl68U/aQkg0bBl5h
zqixENdjBWP4lQVmkfpoiW0c9bhL+NDJzIpZjgNYqlwCDHOBiX/rWMoPzKGi2l/y
DBB+GQOdcKRRhHPpyLu/CNvyvx0D3o4tBZxvJ+Rxf1vEUj25WXELp2W6Zh5YPOQl
Iaql8SM56HTAjvUHPs2OKhuBgtXYWLBOUulBFuKkwfyM0MCUqLLyNndnL3aGOHSj
ixKUsU3+nABPyW5lOHwGaaYHeA53Nk48SIIDHsSybftBPAPvTDRxEA54gqgBg/4b
y+LJ1AB5ZaRH0UvEcPUTd1u+Di1cklH4gFy5AXJLUB1u94jovOFeqDpbNiqBij7v
2SJvCv/MJtCytgSwJs3Uig3x/moeMzJfL6QBD5ToDYAXMj4poNJGOhAGgzT4Uwb6
pdeziWyMG+df6u8+pzYDQd8wSxP1E02bGM314u38WQHrA7tcm/Si6ibBHR46ejQN
llQxmqvrSaT846QEzm/sS6MstgMjO9iY7I15te/rtOvgsFM2ZFMt3mWlx6frwojq
n/vr6Lxx+d1RH32mdByZyNARzgzM9hkgVq1DUleB9eoKzKBBysgpghaEyQtUaka/
p0bgtCMBDSYohtxodye/LzX6e7OojpzQHS6Soe2Yohn7pmsmFUY/ypHhs0/nZ6n8
PF8wmCu0bIrJSB9ktMCWdK+ZGRFjKDPc7F1Fpf/a4kwWLh433rguj9eZcOv2x+Mi
Mc8Hpbmlq87rD+pxslrrNloX2iytNsz/p6dswqNucmz7WJdZDUHoubLreld1DpcS
Sq2x0YIz+DkidytrJRMp9UnQCoVJoQx7edKjYKpyaQ+p2PuQ5tTmZNQkinO9le3T
YvgojK+SK0jnGzUfOz3dpyeq1UMx/nDl+1LTdPYbXYqp/oSSmtof5oE6BihKIf4y
J2RTCtr0ArGVdhliRg+LZYZTkx9LmeCiOK7KGU7Wrngg69IdTXhytr13koEQfKi1
GKhJasE+q5VuAWVpj7TMGqf0K7mGISd0+OHe9Ri9XiZ8AOo3Alwm/9edIOHaUdMo
7LA9gYNcxV63abyMMY5UVbn/IfkPBANIbAbP7MAlmP+ilx8XIZfKoEoyRr9Ieurl
glUSlgmLVlrXvC1UB5tq1ziehlEjEFXj3UnyyyGVmMFMA/eIc2Cpfvot+TD7s48J
9D1O8ldIquInTN9+SnMxPaU+08LrZL3ig8A2ADQGtUmuLENGk9LoLbxkVIFg0+L2
ERygtBTWomWL+AitThTnZMj8DUYJm5eVnz/s2R+Te6tuHkIwHVGk0cElDLGu7X3s
A9dHCA2xtn8SwykhVQCLgd7zDXc667ynP06vPd2KMQbFAFVIoUBjC7zX5v87d0PG
6PuiZPTFxeGiMIMcCjAiaAK7nG1flDZeMp4X1LoIPpME4Ry3Ve13TiiSsKeJkKED
R+Lup/yv2u6LGN2pwPQWGgk5ukjvLAE/Zr+uU4eLFUsuArvr7xlbGj9zGauWu1HR
2nt5EbwYX7PxzDGDhWkUAoZYV5Gj8ZwtOPBTa8y7rd3pGtVVCwAidWQ+Dg3SPqt3
mb3C3xhvq2TrdwttYPL9trYbCilXMzRyw1pNiUlliqTERMMBE2+yGaWaVa2HJ1Z+
rNGx4aqQNuVtbrs5eFDMY06H4S6W52gaJtco+srsbfh+yBbhX3amN4wd5EozEQxZ
6ZlFu5vswPHLlRlhnd8x9KRiNPI3zq7vSpq20R94QlTbykS9W9++/WOn9pM6dv0O
y2/4Tr1ZK+0ghjOnOQL+B4dY0Ifyq+6ItmKFVChDKXYF1jNBFEP1/jra4PENf8Zo
czqOaJwFN/kfyp0Y3RXdCCVtmmoWYH5r72uItThLPUoMxj+MT+b8pryDdcujwx5I
Z+l9KtNrOkYddBJJKpPnZtO9Ezr/KLo2veOZ1/bXz1jGIDQznlJdHdGgutAGVgfj
a7XfwXPdiM0KGTtnml8lUl8NESTRJAbI1JvcQULazGwWamTHeeB+fLfHx9bEYayW
keIJOLpTgFlu0DMq+UwmAjaQBfa2NW3pGEjdDijQNngepGyYvRZ+52CD30mw9QEY
vq9fJHrRE2KSKuyzx/h4ynWlVNRFRAC+9EbxYmUsCm7cR3TShPcGlrJFYJ2tN7zi
grsutGSSkQPVptcG6sVqFuGCr02THufwj3uLfDnqqCRNG8S+1yOSuZtJZ+9/CUUg
ClPuILIWyacNAD00QLGH+BmuVSh8d4t1t+53DcwyPdwhIrl+o7TakGRvtZ8I73qf
ecMWdcTpHD4ZbtN83rI0qI46jjsh/yglOXTJwxJboGU4VD6rpVIx27WQshODtHou
9Hx36kiLfq5tETAIa+BfMRkNc5fcwaSKy6tdqrqEmp/m1NPXtVZKaGDukJxB/AMQ
R20r/A9bfJ1dAXDhnJlnDHtQok8nd3iUkaFaOlbe4tWVlVLbfjL9dfBfpLvX5jCP
5jaCUMa7xS9Yte2f4nM7ubAPXk4dv+4B3tYFW/Wrf0BVo5ZJqqP29huvef7xXA5o
vhQ/Buj23JQExGBrGMb0w5McVdC6PGAUv5XLMaUMroE3iwCLj2gtUdIDTZkdiJSj
iDivrAZsqG6qjEePquV3iQZVD5w8e6isHhVug++6o3fiF+99uOeGCvlway575obl
Q8Lc+gtL6pgD0XBxCQsbSVab99KCRaBYOkq1RPHy5a70gBkvhQ/4GELaZMFinSQc
2T0A9+hBDM5ZRoGlMGRMy2loYK0ApARJfP8S6wRwHncO7gyiRWTaQdbI+9VNn+i1
j+M1LcgH+brrnDmR9jTawEVdz94ize82kYuASK2oZZ3bU8/UrW7TDqPpCcz7ME+R
6QQq4BQcQHscZHmy+tpzGuoV4UKv9wCbKmac6BlOW0amfIPJniBJgMVG1AwxlJOa
cnP5V368Wo9t7tHMpxJMqsQPNuA2h1R+xWSe7p7czv1USvaijEjtqYgDTWkolCrE
859ExgX52AEDGjDrtIC5KkEmCPcUJnjc2qGYsXmVoatKs7nxuNue6acCCua7TKDs
2ponJ5M0risoHKmI6o1OceeONtoaKVP+aN/IHbym9LjckTngYIEBmUdnv5jr1SWU
1GBXubkpwot6HEWAttebEU7X1t1KnANP8xrhiKYhHlnp+crYNTCu/HLm98vDIip2
H5OOf3Q1xuelo+dTJ78KCxybjEGh4NcugKNpYQ9UyJqhwCYn2jozamxDUGSqbtDn
FT2Z/uFiIBE59jr6tnCnZOJFfJWilOhhD7avXHSLQCO89YjPpovLq4kyi8s0NU7I
AhNMZZXWOsm80flSog7Y0LGWb6xYx5JUPTWWiED25ykuHZBtls00QppGmjVGk8TX
kXcAyPJ3LG8sQoiK/clRbEUriEoUSTQI30ld801a14/xdPqD9cKH1fRXQ7RUX+ZW
yCFFYGLvNbt/rsCWbWnXqpkRZwvEMrue028+DPxzRvTfg1JnMiFqYaZnO93fY6s4
JleHWK9sDi5ZTH43AH7kINBxXvGjxkxNHaB8dA6VBIjU+AhCzEQ3xhNzkl16+inW
7k3R2Ocm5gQIGjowbOgv6sCVEJX/Lxp7Yv58VoTayU9Re54dbErus+rMMuZwsD7k
bHybckOEGqVHlmvzHo7pY2w1sV5zdU5ngk/4NgeCdtwWMKz1nbNqFPUUAt+HCS5L
C/C62Qv4ZN5FMatjCIJKhv+2qqB6ImqUEhCInoF0yNkjZYWczgIwhmnyFhcCgA10
8yTSsvW535Ts4hAR0veAvalPxFha7BkNZpDaGr/1rP/Vjp+rnEdYzBTBAe7nMIiF
6Ik+6u3hHZUq7Qe3a+8qvNstwoa4KWPe8KhqcOUFbeqTIwaAf4cFaSazfxgrCMxl
9hJfTB+t/90PGTL2kcoPkXBFXjAMed7uSGy9tYhd4h9/uIVd+L2oO8A51AHmn5l6
3J++ZZL5ZXkY9junQyC1PL+Sxziu/dPVU7w+1DVMxMf1hZx/cULeSsNsvCmtve1L
pc7w0e9minuGFnlmqd8K/et2QCP7qiup5m1FM1EbBS/yznYjiZvv6/1GYF4WFzpi
ZKMks8l9i+Iv1NCLAU95Yq6WTaw3U6i06CBy8F+bofnOcv/A5/4YFcpmQDnkBeig
SrjzXpSMO1bNdA8Dm+hr3U5Dpba9ZACjVQ0I/bTgHIa+/7HFlqBn0lzc0+cOkizF
GwiyA8flAWDAdISyI2kWHBmneVYM6FRKzCCkv9V8aLxWuoNQXoLA6q3gHCZqaN2b
muGDpBhcn4ucQVYnssWTcl37fQ0PJPpy3zb1poodILvzx0YbMhSMQhetXAkD6l00
ZT5KzdxdCH0BRTEUvtp+l8nWxzcgnay/0RPUbOTb7PJX8YE/u3+bFrl3Ots0GqNO
DO47CKsYTJcAFhJGQCjo2b/qP/D5v9ANf1B2tdNyUCpGA7Gna8gWWjDTjlTUzsfD
iJWcarTuijJ1R1y3eyjTlosTKWLmo+NrxSR5G+6VJTnxScSTgYuqGd6BIv0e7uXV
gXKtSbpYe9WZ1FDvsH4tpYQiCmUvTL+9+mAQbTswL5O4E2C58eC/VatcpZ9vaUs9
KrG0ckj26+AEp0vt5yJKJ9AhrsCkDL0xBa1ztcuTEmXzVffdRmfwHePM+rFU/EtM
mGJ60C584npWuv70bECq3bPS/f05bPbL7WiHLL4ImQNoup8T4p3HUDvbJY1k2ZXK
A7zL11vTzBorkaI3Khufz4HeEeZE1dmMu1StCYokYgHhsQCwNN1i3TV7IXwpT66N
/F5iv63g/DYiW+/XX5Vw46WjWObdidtUHfDoYAgsgpikm/a5BAVlAFgx7Yit1RDY
cWbrOWuPkB5x4trpPj/1oifh3f0JTM7saHnOZzIjjp6wwZLOfnm/8sY/ejj/n2+Z
gMJY5XkvbyWatFmQuDooj1OAcH22lyKZOIDSWlN97PGpACvyEvEmLcLmtpI3Heac
bHWaABhZvlKIqs2RC/rJRYUUcgHpVsY4WZYgUGn3zlniYDQI9WrXpQ0Elc3PPiBG
H8nGfin31lx0YmX0iOuF1FyT7/CDchlwuq+K4IIOSlBOyfV01OfEacWJqO07Ftj6
ytZN1v8t2fP7640agux2PNoSMV7UxQX6fWwE783YmHlkGccnprCBOkqI+obzwxo+
hXz7h5fr9jnynXfDsieS4Cw08knxoXymZjCNmpfysP8skjsv76D5+pVXkCnSa1ih
InujR6alCf/l0Ai2XTJzWMGs/ofCk3m1fPw9ulzHnPs1Gdj+Q7g5B+H6gn9KN2KC
zvgt9vmRIIvb3Thkmg0lKCDmre2PKK1w1osgsFTvwA1sLxRaELxQSgOvwE3HWWBs
H+XRXTIwn1GoD+psqRhfa5dz6H6UhHRmNBkBQv7IOpAxSSWA5mZrnBjx27/j9ZCk
lziBdRK8F854hYDKxIubuhngr+oLVb17xuYq6M/QkUtfRZhMWpWyVroOPzEG1fLN
U6+Yweh24qTcgHR0+/G9dOIaLblPcsT1UMLFkyFHVwkOqIDB0NMdJsSVVqxr9i3e
MyDlrMy9XxdVYOj99hUEFZPSf67+NjPW6OXAJpC+YjE48SmaV2tKcgs16Mo04Wvw
Rpa3XvlfqlojaADuQWoi20/GAuAU2AGApch/6hh3jAob0CZ969J0qhPXv4VHl8MI
8YCSnCxT73y+6BjLEPHSKEjjZYivU9pKJlEm08RaYEmhExODWxYTrHZ1BqPRGJaJ
0L4StjV+pP3EYCZrLW+TnrA6e7msSlqXPkWE/rSroXJ4cm8/eGzZIFCb2fTRgl/8
+GSfjKe+KW6rohZ+4HVwTodE5Izero0NMP54wWArJSk4k1OuLjqCqp9bFtFne2uY
yEq0R30TD/+/Zb96CnNqtlnJgnSrlFcbNJYLN7JivuymLXE33hejoanjMzDvzguY
ZjsBGDvAWvJ9OIEw90SjTtIRyrao7WVI3Z+jFXSBef+Ni7oKI3QSobbclA1HagjZ
O2PWK4O5m3jgMty9yJnTfQWR1mmvCHeh4uIG+u7yRucUbOzhPbJVyhTh2MaoOa75
XT4J1QkLAKctARO6Cmd6E4LfMkZf5c1jpVWyKHqMzrS4p1DVuwt1/QPDkVGid+in
QYcZanoNbhL8VnrQ622iz8clQXwnofuWzhlZJQpm6LMmO36NkfDy0pyDMqk7lwFU
n4lopZwDba4Vf0JbvOatqoFeQ9XjH4CKbbAceDH7LJkJdI7wMfBLPhKIIdEHondG
I9NuQDggccGpjxVFcjSgMGVR+mncCG9SqT/NLAUh9rzmFg1IEBxQAHfk/HpfvQeD
XhVLKTDAgsgCRVNiHK3RKgsV7bOgDxTx6d+gF703qer1u8mjbdp6JOSpQKd/K9M7
QQmB3njsh2UVEN3DllmSxzVKwKtUE4t29Md4/+BA9UXqDhhYRoH8hebrocitkA9h
4OSJc+19GQ0YTDkFQLo1cOx4FDen7BDyG4CN1LNjWoC22ZE2RtCKGiBMZW/P5CI3
jpEIJaSh8ycCZ1QPg4auUEaXnKfb0IAntdDXnjhvnF0lwJRAz46pLvF5WUT3zk0k
EeXs+GcOXCPc47Og1DnCBrdkO+pjXn1itAHclT2lyd2E7doBC7OO49eiqCvNfNrO
gQDSXYzqwttR83UCgswQYrT0p8JwzmQSFdnMeOhN51rNiQv5icFRm49MWcXTCRqC
RPxGZXwN3KQLsXEUtuqE1EefcI/NGGVUg/vkLea3Wd0c6YbCuemYBu6E13OQkyO8
K8f9rKc2kwd7RxrBGia3AkkJt6ZeyeJvbrxHNMEzyuaToOTfYEWUatRrNQ+Shjin
lIqBN9pz4dyLFLaLVN3vi6HCl46JMO0gHTLYnghdWA7UgNlczoQc9d1fNoV0uisY
WOrB7+ypy3L8ep07jBveK2gWjvtgt23wKKBM5xwourjOkbpuwrl2RSR3HtVZB7kb
mm3H0K4fs0WdEs0MdtZkesvdN8cLN9n6WuY52TQzi8l7XyyT8Qn4LU16Pf0LEBXK
sqEdK5nhdzD4mVJYTbZookOQy1RNDp3I7j9caox37a0LCEkkSoLlCf6lAHa8HqYK
vbGMU7xfZX1Hfgnk622WBmDYyJYEeIQNc1ARtOK1joPYCPZqOBV8cOM9KQsmC83l
zuUU0Ygq8Gpja/Cgwot5LDSrsqh3MXQ4mpbzcLPOV54k9NebSWe5FS3McKtxkLb9
83d+NVpMYwSjJw0g2p+zkQLRkOWZG89h8jKGFDRqiZdDJi6GVjhVO8YIdLEwelwS
PVqCxTQ5jLmLpB5EJiIpBIVTDwg6CV5QeOmSyXLMyEeO2ygMfTN/ebjG3ORWY3Ut
KIthQsM7jcxxUeCikIkhyBCommuKPJDm0t5cOjV4KABGUNI/8dmHyFkdeK05bwic
7LF1kx7Tic1LugFO6nsjpszzm1YSks+sHO5vp3qlTJAnOo0J3doboEhlc+H5GgWQ
4erxsIJ25cWZaMdThUCSaOeX2XfLB6Kmn0xa0a641uN4gtGKktPC3pRqM/Ev2gfZ
/TjYC+HDYo48cTaEyYpLSOBhrbrQztIsjaw/jLxgMJT0nlaAf3gHn3m13l8/S2cu
JCHF1tOP05mTiEuWw9RXSKZc33QkmM5G6U056qX5SZ9/vgpEU/HG+MH2rAoFEeZL
PFNSK/RpUjNUxIdk2tH5zVNwAMjfcpT99UYaY/4G4cpgKNBaTowTCjop0TKIX/D/
FB9iSodAPDDb3AA5SeLgIws0OTPQ6mvRUT4FtNnF7Wiu3CZ6bwchdB/1QSyVfQ4G
u9yN0qCfDYAQ46Hdmth2NPgggQCjRF0tkNmMH5cLNtGXOyugm35ML+Q8r90dB80N
NHABE6v7WX+u0Udor79bLHT0DXNFzr4YbeM6H/C5cM4AYC1yd/3g1nbZyI8IRbDM
OcEn37pgTg/pHZU8B8fFpmScjLBdIzQ0/NMOSlB0nYq/i1un5Hyxl6ZS+3w8i4m/
WDOARm2YPamWfH1W6qyQzZUQrh8fhk2vgx6/f1pmdEeesYJM0V+blhiU3pVdgXhp
DfUyeSWFrSOTF3N4E161TJzNSbE8jJb9T7z1NJs/limA1MScMZCBLHzredUftFai
RtzMy6svwGacjnj1qLZIZMUwrX/qUahhMk3AdyxrnGCbGH9EW/X8sajvDdQgDcBT
8c7MTZ2Z6eBR41bNEFEtK9/RfHQse3eAYNnAviKCkTCnttfnPxN8A/9xl6vEI5jj
4okzt+ct3c1BQZZOpBFMvmvZMi+nWYFbMk2KelZyoFboUu6RtQiXIyzUJhllS8se
xJb6Y5oexwE04SsdU6iSFbWzzEItAVbOuL9ANHyQUwE3EmGKBB52DiBCd7gPbsUq
DmIx7TOIIyT/VDNfipJ9ptWlR84RJbatMy3IftBOQD4l7/FDS5sDa64YOuI57XC2
oFu1MX4s3c2ewhAfV21bm7J8beSiPK6w5pZ0zg8cag4BKICW1WR/Ku6zKcOlKiXU
e/MsIPURD7W2BlDVl8dSaWA9ye8MMr0Jekw2beYNROZpfGxPRhViHUjWZm5420EI
8pYNcCq8B9AKDlQiswAGx+7cGs7z+nqQuim9jRyMoQ4tCCujNNayARd5gojjgvk6
KNpuPOtfO2UVvfXuPzDQJSIatmF5muhbBVtMXOm2vcXRTh1ZjH1NPd5x2as52x89
9xlrkb2xZ9bRO4F+JHfnHncysZF/kraYZk0mEtfpY19mZoan39iYJXDwkfVWoQp4
PQxbCiTspE2tK42WtSbXvCQYn+Etzx1qg6J9n1mbaRWGDtrtJEk1kkqs9U7z11qp
isI5hJ3TehL1pWZzbZR1csbHMzcMugxVEBOKQpPXikdwUB6/KwTgzsOzWMOvb7sF
CbuDUCuAPtklvjOnUQewvnLlNbLc48ihMx0zqdZMBmlIdZCfNJSxiRAvjDv1uryc
dE/WmmD1v3XO9GaAz9SMw1kEBT9eMH5q7wwMH/r8/g6nqrTPOkLHhMS9RCWTaVwX
ytlYVIRZEcJeJV6bwXGyl6KGFSCfrd3+mO9rkSuBHULcmzShxykSrdg0U2Gwl4Bz
xd05kbPRzm6T3kiZ09RMlBNjtgJPw/yurFjXpZWfBiXUdVrnZGo10sRv6aYLYOHh
5lnlgq3hVOsS0jB1+R+bgUBjU+H8UDDSOCscwn8ik7PtACOvAkDsKwv86MgTRtrW
t1m0bro8268v1RzjJiFOWpKXi1tGjMucSnYkS+vNLTWEBiqcptu6HdVgOfn0kR6o
3zowuvZ4vcrdSsLUJCiRSYoa80++vd9uRecgLwrNIZ5+3Dh3mZNA8co6yY7raNVu
3xo1c4/VW/+ccxCYaZ1ExfbBqHit5f8eilWj1ZWNL06V+UhcYEGH7m3aqdwX3Rl5
kJd4a3cZJHdvfIZ6+vn0/L8uYvBjZ/GsXRs0cG4Lyt3j9RoCU+4H2sLzjVvkJRqS
nFaSCQdJYXYixYpRDohEMLkm9p+R2DNXhVwsq4f/M1VRfXKc5H116eTknBpvPoha
yPbUnxHQGyFhMUQ4hlR2EifWW3pgw148c+ZtsfAKGbT19oL5UoNz7S1uAHmatrbk
6Ki66bgV70m4uDvWAdQV+UxjjoqfkuHTxPlcM4JMoPKKlzb+KTsdNoAn46Yevs50
uoMFi9eOiDvLsjiQ62+A7YkFCGDggF3bbQUfE23YZ72WSEr+pDqXwei+wXL6rNAT
mx0ugT+AG0PpLKClUwpI4wj5y0xLXEg3SGlpETXs/gKJkEhLFVGyW8jjy4r/BmVI
6EQHjjtnlTI/3pp0hORQSkdwjmi/ckHGmfyiZZQ2Z75k2qNIzq0Ivd6FkwOWfWYs
x5lh+42Rfk+FBJcZERlPPRzMgJ1ipcbl5X9HFZHld5PKRUnde9Hc9h5g4kIS1Ni9
RP0vWd+4pflJ4H0ObmYF6YgNjBCYezjQUdw1m9pla2nK+tDae5HaQ9MWe7n1bPHp
+n7T/18UKTW2TOiXD40SC6okTEWXL2gQH7gyklDlRwAKlR+Gmfz/Ox8D8hW0GP2+
9aHJ8cmewDHJIEjt4kdmyP7wao91jF1MPPGB3uBQgTLfHB17B7MAOCSGXssmh1rB
PIhpG3gIhZ1/DYmqljOdy6MS9i0MqG6UL5a4960Pp2pP/u7btEf4yaZxUnXN6PgI
8capUXnHfkLgC9tZcQCgFdkiVBNZ1se39gSDQZs9uTjri52PZJ/ZK+i+FD+GAd3o
fzoJIp11IZBX/0cEDoqT6fKqYbsjzwYkqWYxqoW1AWRREvuRUNVjjDDuJV+G+6AT
8sLY8FSKuY03SLVMWcGkkLT8lFI0+9N/ocvst2pOwW5rgglnYLj9QmWj0q9Xdrnz
qB3YdgOHeNGrkmYbUjEQs/QiG5N89tHqUQ5GfSp7+dhv5JzXGGpcyCL3a+7120sp
p7FblLNh7LGfNlP1MkjpPj3/0BPD3HLJDKr4+pqegojhzZcpN1mSwVGv2tKHJKlP
XWG5ly5ueS4jU8CDgDeBgmHH+ZWahzfYvm6PJF5jXO7D3JIbbSZYFF6u5CvPOxeS
0zfWADnQq29k4jCfPk7UDZmH652IWgkDnuRa7O88S1i/wt8IEqmfDj+XYKlIT/HO
46g8k/J1mV8C5lBW2yxQ9BnKi6SNHJY1cXnWK0JmkNB/rxj0aIL9Q3LfTEtE2wm6
0CiMKJjnVrHPPzlYH+5JHce0qOiPb3QiHfzzGJVyP08l/nypEDx5ef+jWY9NjUP3
TfYU8o1NQQj+askWEkWRUjSOlZwM71cZWWXpGCp4+0z1B+3BZ+jvCCzqtABl0Hvh
Hw6hbYmWOUKvT7D34IxikUcs3jwQEIrd9e0SBi1lNcvhsrYqYUoBLzdNYK+aJoRV
KqaiIC3+N9IkXIBgHBpPOfhneF30ShODhBjJmHrbsfHn4i798cnZbjR2zc2142qS
w70DtopShSTytHTaTTAaqIB9reL/xAg+4nVeG9G4jOZeLSDAOellxkug/+lD19c5
s0pY7HOXgiq2F4X0HPGp+Ks9YalD6yDcUpdPk/FJiHWzYCzcCplN/NHSmQZAM74S
+CxzLE+Cvdy5A16n+RkBTGrGdLOnp9/NrSHQYZcJ+/enueOLJ54wqyXsHnCgP7ys
xjMEqQjIz/33Vq0icVgMquled8QgqRetKMqG5rzIWK0Le25RF5tKoZyhdPbPM6yb
aL4p1c8/l5AbfByhhR9Na7riP2KbzlUWnF6qj7uFg7f/daohiwHboeu6OK9XNmzb
S0KKMrTZZiK9uRjmLnzDwYCKLrIaBTP5jNdgyXj11z1yv8PBixlfXKjQOVfFEOkQ
pepkY+l55DZCnkYqrhl4GaIXs3W1hVEZlw96YBvbYt6x5z9stsdilE03u7dAjH6i
PVGgeJfXeIejYaFcGwpDA+BLItTf6UfuBMDLt3pUM57yPTik84NsyDf0nFICWEtw
uPjjrujhK5zC4viN5xor0jvN3Ae/Jil1Q+v9gT+PsVvG1URLV9L9JgrvZVNDyBR6
BRUOYPsx/3Dyka6aVcz1lzGlmoQ4AkdynpkmX0NFJG7uCsltvIfXUuDvgsReC/kp
rO5KTG/eyN7SQXbjBhD3cEIIIEDhuDi6gfzmCYuhCUIM0Ap5V7sUC2u4sDGS/PTZ
4yjItDRfdtVxD7ilIUgb3kUDW8Hm5TUQlNDmPycYVFHNkVWiFxvRCNWfGuOY4VUq
ELAAF93msW50xS2DmJrJ7uYHPt51FKRlvVGhnahaOqDF28n+7xRNjcLKQGTOt1s4
DqhyYfnzLXy04923CrGWH4sAwzYo/cxP9Zc4YOmtXud6yag1iVK5odYz/gmnYkKj
JcTyxXKk9x+WG+BekDlrcGySueQJrX0EeB5xkkqhHr7SPk4clqXMJqpEeA8bfzvu
gkXcHKUNUSQUVVPa38hJGmXsARQmlYs/Bn2OL8O43aeeCC/iDHbjh1uCOoUWyuZA
2yrBUEVF79BXooVj3fFMJcMrWieSl55551f3RdIhgG3Mxd3e9MLwyoeML2f6uLS3
mDU8vM5yLWvVXDqFe35ZJgBD3nKS5F2u8/bitOFaiKy/KQ0ZHVmhTEyU6KWg4jD4
or20/BjtIwVvUTwINVkBPmy74/u9hGPf0jPxKqFmZkbPU7tzMuff90EMHn9KXqGX
cu1LX2in+kAvV21Pa4RoBAZBzkV8+xeRU0scx4Cp3WFJd4GQJydp66+tWhZhFcMV
fOZIh7kzdBi+YrR/gxmuOvYYO04BvbskbQKYmcr+PBX/Vo2bwkmue2G94+jpXjoW
si3/nVXXfy8GeUWsGcy488VKz2NsI3fHkSLhHhT+KZOoyNNhPRGNe8bxHGYJ4xBR
0C5WurBYw9ybWZ9bF+rPcx4XEa2tgW9bc+jjRKx7bn0Q/03WBn3ta+Fgmmp+aLwR
+lf4cu3HgluITdsS5zojqTGreoy70Dzc24qMHLkyZ0duH86tV9uddW01Q3Ii5sDO
Vv2D+I8PVFiqbch+IgWFBIJMQyOpez1E+77dMzXSUm6ckbLVcpAGmW/oj2MkjVJ0
Q2OcD4DwAiUd+aROBT19FbPKqzKrpC6UyCUiRuDR+OeNqNB4WrlwFU9sj2U4eyvu
9Wx0K3LpRf49tVyY8FGFxxWBfWnyNL+v0aBe4ILc9q3cuDIqBh7ZHHP+am6ukXaz
Zdd/SlMKj4XVrJHaIVYyYOL78R5W6SATGWq/HCUbkFxaYuQ6vhSOIQ4Kce3qAZhC
lluZbHA+4vaQLnCflvxJLvFEYMpHknBWXHn9V7qPQk4DZQPANhRo0scTNLQ4I0kd
2x/WFVwCSnVb+35g1dnTllTDghOMckqq58qrD1pnpJ2LWcYy/7CTDhAE55JYHueb
V1EghCdAhBydX30hqHKuSebpQNTX4ElVmuqDJxqA1HmlaOoFwPxmxCsctoi4iwH6
dFawZSSqcY8tp0C1IH8FwdddWb8XJ6JXaAaCuPEQp6wg8zrokNJKA+7chsWA98Fr
33TwwFcT4w2ujNn5C4urR3w0opfMePzFu5APHaLt2XdKxBcHa1mUncXfqhgEZaWu
6I1Etw0GeuHczLA28o3tE9ikU/e2CNPijlb8/O8Z//p3dzV73530KsK5j2048PcV
BggynrB65YHrCwAsddyeIfpvFlmsVIkCxgN1F0DmbER19e1+KyIP3x3ewVO5c8il
1yy49Rz4eu1Ep6xvDnS5BLgc9NShKKJyDgYTyHuYJF/zXpU279cWTlpV20FRRaYE
21QKc6sZ/IZ/INO1muO2vWbE2qjOlOL4ZfEOugLNlc/P/AcqxfsAibdTbdErf1/L
/O5XZftk5G+q00sayWtfP502oBwF/ifRe47d76inkn/IGSX8ehKdxGTrWpGzBH/e
eGNTvX27DUj/dOn93aIv89TbI+El6nJnrqlSsF1ARXfQEgWqFBXyy7bTvUsvNEM3
jac9FNAWC+IX7jD7pAIcct1ICq3JI2+K3/qiZ8t4XJ57sLD3YSVgD5D3l8y42ckZ
svnmetFxfTOA7/9knTQYRrjQAqi4gvD0k1YcDj40fqyqtFyWQ1RRz56yRVuLX0Sd
CD3McYMijnrv4Lp7HhWPn7JGrivYpeZ+neGGDTrsDWW2hpKGE3hRs5otgt6yNBTQ
6evLSlbbmiV9ZmjuNFJ88Lw+TNRmP+5nmRDRe17ZQd2KWcNQUoljipqWfjSyYhVX
x4a69Y3i/64orqxSPdIuuWWOftaq6dUwGOulWrhWXNtFXSDqrYMIMJBA6xJEYY/U
9YqGHVPcZbW1TLXDLG6poAiESqnNHbAj6BtcHadp5ap3eJ8Vxo4wal6OL6MJ05vX
02SvZrIt7R/+jMkR6QZbvSuTtfXtGgK9CRasGfQ0ZX2+u0oQImMeV5lViy4a1k5l
wW43L9w0lN03jfPBCTjx7lAeXsnCpdAtoVAv+COqN26V+6e10jFOryX5/bPXxarO
/GA1h3sXvswoG77N4dflfTiLfQ3sa/FJOwIfuo5J+0Eg0aT50wEDc2bU5gz7C0Dy
vBKXrZ2cKNc1PS4uHQzOQtzf4VvCs3v2iV8g5Tyx/Gc9sJ9iyeIPUhMqo5vzAdbD
4myli1NtOVgHIwOtPtEfQEtukc9bqw+SHtNamP6oFZZ81xoSaycqAh5QsrezwEsX
UnbxGX6TOmwCgxTkM5Vf5nGTG1+jr2m17+fq3NxndnwEI5GXwMjaCcdn0WVcqR2f
RcPVYCNTlfn/wwYoT+P4zTWGOSpeRT/o80169aPXwHwpkhYgO3l9a9SFFwLiW7KY
PvbWBewPZPSJQFEnLrw6hy2WDHBNsYWtTYJVTyfNfq3Cr+1hM5/5gBiByZ4v8t/h
jJFLTMzPHDih0RGVN+VzadMNLuNwAmEWHoo2EtJqkLLe7Ixccrb2KNx2ihm0ZtKE
n7Ky+FNG04gTfOUOFqBUot/C03q4xcrVTpxuyrsOLG4L8jQXZdvo0zaxx5ybz8Dp
+Zdi9Co5UsEWc5ADFJvkOCQlSp0NSYRepiAJztFKSDdbF40QGKeft8Z9XEouNIgH
yAx44M1C12wsUlVm4063SYyOtf9+gsVcArCj8LTxVca2q+nLP6/o9pOi/9B25PeG
P62hUX9Gv0w/qd269FygedzBcMM6Kt+ddVcEXPCJB9PeIUwLPeej2rlH3ZHg2g4A
tsvMPyFAGCq2mcmlIJS/yxYOowL1rFPQIpo2JVAkAfhk3dCt5zbpMck++UuY1/jG
6qQHjxtMJGhw7fN28ob4GuA8dWehHk8a35wkfyV6NkaWeNLxgvNbEF7zmFrCiH11
v4BM4FzUEWeoDyofH061kWtoYJg8Fr6du40P7fprOyw6LN1WwcgqsyetgrCRFdMG
LPnEvh9Sz1lP2gWzg/24eZMJUAApFOh7qXEVFVW7MPxo2Mvg/2bVpJ1VKcvoMAi4
UMsdFjThSZAjG5Yi8NJN3FWDWbjHrKOCy6GAVng8wpG1gusHvhmS06RvJ4KCz/VM
H2n9fZ2mwjEU8wgRpU0fMU16Tn6A/yftZJqAP7C0NA+eiBQvDADop4P8Bnx4IaWA
XFyY9vxQA0778zJtzRxlSmRTQYKf/BYawQyJBRWbCb00Us7XGdaSdy680YuvAUs8
ebhdZrLJogIS3hH398bekXZxFGG9undcFwmb2GFgOt49U+Qz2KEU/VZ0cOXXckv6
/cTvz8E7N3/WH/MxuISCmnM/CwoXdbnlC6Cp+lk2SLnwh7C69VZlgnIOMdzGmEw4
tqRqWAoKR4N1c6AOM60wvj66/+F28kj4q7SlqMSs/lEW/5dm5Q+G8w59MMxdFHTQ
Ecf8aMF3BQ8tcDfpxHGm+YdcHQH5CgfgDRCvZBwAC9093L3/YycEABKe3a/GV8Pn
EG2EdD7J6kYfJRkAy1CHfaXgJ0nchF1o3jyzXcFPhleghYttzCdo46EVm8hoTtiF
NLJHViG7bin6Nkc/qjHYZKzXUU2thkd4cgcWn4LT8kFI6q5y/AMric4z1Z6vegSb
n1C0cVAsGFc4KnKmOvsUG1eoCp7nS/A/h/BUgkD01hfUtiPvdbczKhd4yqqxxDFa
0X+DelagM33/xs5qk3ZnqrZahc82zo55hkiNPrOUbnLrVFu8BTgrZpBUSDntu3Ek
8J6lkhYCgjrwaeA4CPrQzZ5R9Ey6PfHe4uexMpdKa5FGpw1ETahzwpgv7EOwp4OX
mvyVOmrSR6vnjKnHFmP7GnNDX1PbwiIzQdK9N0IoqHGyr0avmqWyexhy87i2SB3a
fOv1ILZu5WW9QHslSclQLdDlVcZ0VRLHG2/54ozHdaXcn9XRkIKNDFIZs2ml+Ia8
EFVkGX5uOeh/gZI9enXpxOIECfF8JCvI8wY3yhsDRVxI9dDx4ygA+oO8CJm8aRck
BKIF/nvZcTk46VksrqGoITaQejXQel+WBHuPgg3Kd88+M3IeFc4msSMS2aOpdpZQ
UMTVeVBzlQjljy7L8bXjVmBLzpPEEWltD6vt/t6iGB3ppdmveV4m9FSde8Pra5Yg
chXhAIX+VIr80StxJYdL1iZgh0PthxpsL3TUlbtvSktqHX29DoeTFWliUx4L6/yG
TcLUN0WdzDrJ9I1GXFTgZzEpwkjDNV4WB8cRNd54drHzjLlIb6fvV8KWe5zEYaeB
iROn7Kf7Lh11AUfimmBRtZMPzH8HvvhVm8l3+F7h1JtwHxscWRC6SL2Sp3h6RSFE
woiWsignMXDdLpczlwVXaGKFlbymn12EPGpSDD2fBLPuC6rKGrXo/Om+4lpKSHy8
15HIbBzmoefDNsh3p44vfgETx7QE6mepX3lklq7vn0Jo+FN17kJmzd++zUMCgSqA
smHlG01zfXF4TGBERse97Z1Wj41KJhFslYnUO5EfeKwnWPHy7RY+sBX9Z8Q8XObb
nclfb8ciPjvsP4RmmyhYCN+iWspMwCKGf//N86yWvxXaIHqX1fjL0UhkbIZLC5bg
Oy1xZsbl7enFMfd7I2P+x5B5meXrzr/ZAftPjKUEOrmiN9StW3d63S+ZKvrnQ+TN
TVzyEke4CGtLnrZEZZYgMSCha82h8ArhHwfPxXV2tN3FJvKr4MU7jeqPuz961nJ9
05VD3F6LoHolgZfGf38Cpcgq9tTsMbGHiRMKnAEmPNurufjwK2jhsqOsFgACpXj3
LA5/UfLA7WV2zsZV874lk1nISuXHN/q7VT2s9U7xU+sHh591BbN2bGwW4H48LP9S
ZnJfj4maUGcjQU5Phde2NjfU3KfvO+GCXlZIddPTLErm76kPrqwMrsIICh7q/n3D
FNtDO8Ar9W4nuhixWluJIkXyZa0VEyJaDQUaHxCLCW4uy4JNjTh2+78pwY7aHX9r
V949bokBSA8aO+GG1h67Xv/8pK65b1bw3RvCorxnXCcdsvwzfDMNhsaVMmx0kSq3
qj4i2wjf9UXNQzIh+dNSCMKm6U3KsUqD36Vk+NlPuxX8rCAPl4SQXm2qdAXbraXe
Fp86+gDOLLj0ZwvYtdj7s7Gwc9pDuICeU2w6GTlteGB+71qgfR6eCzUMIVKMysfz
ji9G5DG4LAkkTw+ERKbvNGbdCA8AefBmuA7t1GuJ4CVxuCqwHi5eyucNE11A6vBC
Xwh9sKXoiUwKSQu05i5GSH/urhXUwcr5lPpM/PBu4cjhnpZFkgL6BuwrzN2beCs4
VOhYzRL8V23pfU+hXne9/wZwR9C510862uasY2+W/ZXANZZ8t9zB/U8tjzbtrMOD
gttm7ALeZ+9+vCGiMbgqjXvlyQhgB/uUue0YeSbTLuiKiLiTXVq9k7nJ7HQDL5cn
JMpIbLZnzhawP02ZrNlqA8/DuSZLL46DViR0ARI0VYdS2i0u8jfczd5DCI63LWKt
X+RhaIdNbApL2q4Ka6Abs8irqfNb6949RuLzyrmmRxkvKNp6wjNadI0PA+IUOoqE
Q1cEbm6ErQKPs+7TnhK/UzaVbIA0dIqASDzf4y/Kr7tp3ByxNvckyCoNNnh2O+h5
EKh+IPJ9/renlO1tPQO/rXIx+QnikalaFNJyfZGkF6GiKSOv3WQkjM1F+MI48Rce
H4mcli6d7M0OgRSWQzAzTgYFURnRk5RFyBdFBK3cV2MPsjM7iljwQvwzuU4mMAcp
Uj45xnq+xJZDWdDEfj6dKrApb4x4HNVraAGwKvmjDTIgtLrx+Rg8BD2x2Q0xmxpU
muB+Bx+jnW5zlZ43WDYdluiJUud7Y08owZc4kDiM5pPCHFIhlsirRO27Iyik7dPT
8rGeY4SOcsMXCOpN/Rd3kagc2xR69dL0EkxeOhCM0zGx6bmxsUsAritIY+kqvBPw
VDJa1emHmSeEzry9OT7Akth0PT3FkT/BfFvuE9uE2VHkEYdcEyfWO1MNdsMOItEz
dbkjOjgJSy2ES/lMAONzKWvw6eWmnuXSw0fLorIOlEy/v6Gz+0HTMGZiKk3c7WGi
IvMVGrgAhHShwJO7rSlkOjBzRQKwMrPC4uriNMuNWb13xGpYZWKsniLba8NjL41M
KCDG5XyroB89exCA4TYyCCP4Hnwmyta1bvTrIKS/zbN6mdLhelfKcfV5uY0wMafp
QNngVnfQHNNfDhBkDlo0Y2aJ6JvGPSWE4X8DIAV3JVZy9iISQ8WLEX9z0exHFK1v
a3mo0G15Skn3BLKs1a/2W+7o9x0cTpWcj2jsED3t0vn/O+Z8WfYvG7MOQ/PgDowV
f2ihpuXqQp+MnM5mTRUGpAMhzDl0TEpWvFmwRK4kR3rU2rmJ6fk9iaDAJacSdsw/
VQ1ZLQq6E9r3S7dvklD80cphA/f+Aw0dhn0TvVhcH+UVnBLrL/Zr/59TRzUiiZvf
TPczc6SXLxcVvvFs6HbzBhVwCiBP9HOpN1TFQjX+GjAFX5Nnc54VcAGw4YMC5H/7
bDAmVFp8FZYWX+s6vZ2Au8EP7gwekuRqzgOXZ5zI7JZFfeXi0WTNMZTBS3xfDBxK
bnYbsfw0ZFdveF99W1AlHazhNjToXhcx86cIAt6S85sQS/azZ9bBKV9/mjLmuoFA
CgFSx1GdMk2obVmUI03SV0XzP6fQQ0M1DwXGHUn+Mk5MjmHx6IJ1X+8yu6Hxf/0U
7WAzT4JMTHYtczjXReYx8dZrkVpgMQcQtXvDlRYlGEv8boCJKO9nIhpECutUZLMB
ubUWbGQdIsbxqklGiz8CT/Ubov+k259lpTh1tRYgYYIntfYElTXMmNbAK4H8yroD
cYR+iOzh9GghVm3KSLsWr+6AT/yS/VOXW4atrLXjwcdURktaVklVAGjkycARrODO
9QYHaibsH6UCUVKww+zfkrtSRONuIs2h5nHjUJdCsYpE0f4Ih1F+Kn16rOsDkzh7
d+EqlOmXFTGarB6hk1IG+IRxQGqil/4+lG2hobgpz8zS93Vb3sCp15PTXkUhlZ9L
8iNJDoxW5BfvEFrP4jSzSO1Ru9m3ANBYutUxdG0JSiEWOXXayHUCVhrbwQOBiMxb
pcLwh2NMw0XOHXrZwWGCDv5Up+5sxMeySxrJRaWR3TNDhQwcRH53EXfk3nwuP6af
IowlbSCrNtVWPhnXQG+qwTDfi4BE/w/4osovNooOUk/vb6LX1W/VObueXFmtmsPF
wMd1xuUhj/dMuRAKUGtvXRNCdJd0n/3a7S8FIYJdLUc2fvU1Rr+J6NEHlkb9cxzh
3vE2vYkwMBi5hw8X+6s0X/oGT9ocZeALBhi1jL3YTrDykcdO6oXHKoYsz6ggxiG0
2GoazMbZ6UpCD9Na12KJ2rttzHkxWpX0P1qQ8GLlhnp9gTkUi1hfbIhzgi/O5ZlZ
Q4+lp/Q+Z/DEU3UcENiXdgwDplFbHt/t+bKUxLAnUHRurPgJSieT2ROwrZCsPT08
6D19ol+2oWpiNIkAn7nillRjbohoG734o3+26mmFx7tuEqRZEmy6HpkhGjA0q3eL
5vX2W8FlI65PRNTLo0fkfVHb23ffItLJaR0Z50nvPvwUfI+TM+i5bKmryoHVuX2a
svEQ1LySmuedd81LwjzfaYTItgAOp7hleiTnz/FFh2nCvnHK6Ye03Yxf5p/EKP5g
L6E95g5GtG2iDwBkPrfUdYciW5hHVsyehjzSi+v7/ZiT/E6fQs+H2xArBk9KBXWB
329UAAYyOL75TsFsXiXSCsg7Nn7JXo/7VUkZODRPT5v4/vgH6a79nxu02MrdpkIu
asSrTMB7QkgswIeTW+LEMTV0nLK/ESQ8b9XH0ixy0/JNLf01ORByCLzHh/EenVi8
RRlZfCPqKjZIIw7jiv/vcPlv/L0EXbHRjogM30i4Wc+zjFumO42nP7ruaF/RVnJm
QvnxS+JPd96sYtzXHEqfycXZWUsZoWCleH85+M3wRl4EWuyqYAv2Qf0VQVZfhwPl
Q5tifuO/9DQrrvugopMjmREtawWoBozqJNbe68uDv/t8mBVO/giZzdiMiCVq/ntB
Ad52/IabFuSNLKTQJ0k0dSx0UV3XW/KhfWKBEw2qiJYSpc07LWwAcOUHjmKlrgLT
b7j1UWNr3Z5LomPrP3xiv95qhuPegaYb999zgAjaz8O0ZweMggM39FNHkUhVGqPG
sYrlIxAnHeuuYhrADTHu46ASb+0G1xI4+PzZ77xp2GVESyarl8K+Ua3aU+xwSSz5
PmbBqxNjdML2T4Td3OjRsJzh9GWoZjBzNIyJ/0iU03bRptF37MJQo5ir2j4LGeM1
0FuC5tQYkXeeTfcziHf17gqlzTEv45fIM9i3O9/2eYsKW28v36xGHRn6Yivs7RvW
wNblh/8RK4cBQFJhevxP3I+G9ChYViqsaF3r+mkyYA5PebFGPK0SoC1gj9142MYE
r26gz45KqxcOlRkatnE6dNUVxAeXmpSNKrX/0be7SOrjYqCeU+E1bHDEsYL7bT/q
pFud7pR8XyeGuMn7Ux0Z5aIHGSJoNM4jbPcFM8y84F7W5YNNrZ+y+T3BnpzkG260
6hKJerndp1saSy/KD4rPOQWx9UGU+bcB69SbY5l2JnIQs0s8TqFp7LaaCpiluPsl
JORNhvwxrLIKnl72PVFHN7bpcCgSZX3DpLlmL2pUovZsj2SxOpRWpcYWoQisKPQl
kZypDBiinYu0xZe92D7O4e7fAUv66F5t1CfRhSbijjUZj6bRGwdJZ3yT8Lv0BJW2
s64+FQP0afN0ufwRk3/m9NlTfGNFKN7KDPBBHwhw9V8+KVvA1AMhFJZSLomFTAQc
8mL+eLtLJkYDWTcqgY9KOhZdcAI5XmtF9pIi+gohQomo+OkH72sKJPr9n+YsyuW2
qmhcoNRGvh1hdKrNngQgZgyQxApJBrO4SEQfAphiXYu1UKeMbpAJb6uL2UeXe8b7
ztNdjKwAtAFrQsKGbPdx/CwdNgZz+LlyxLJxa92t9lBEBpvcKOBsoYaMwrhJ/N2Z
susua54TDINezzedSxpaxezEKg9HIpQ5AGKFPuj1zVeuKWADA06pUQKkyUkYSCYI
FEqcdB735Phf/HwTS3Oq/dMA+5o/gfmYh8OxGFWMzCJW7bUBefsf7zhagZhTM6W7
Szg0lLuRYoqd8hsOA9dl1ZBftrMGQfEJrMExxLfCd5UpHyiSMR8zi4J+xz54HeA6
ks2rrwc3LfvWEcDEQgxFMo3JY9gZYnB8LxdsnP/j70vNnEqN/qNCPUJENQCmbG1U
JJRdskQvTmDqZnG1oVR4J74fihTCejjeqjjzeyBFnf76b2MAE7xq2bE9gtDiVo8v
L5MLgh1zRNE3ZXZV79Yay6ybJEi1mUJH4snh+2RprdpmW4BlQobARHcDBpXXQYdy
UqKQ9lpToMuCsfIVBDh9SQifNxv2oM20H3FTZ3lIcf99j/CQnX0I3Bs+5+m3PJPL
K4c10iLL8tcoo88IPTNwReooDMebnKJ9y5f+/43UpKs9E6HFa9x7V+rguTNYAshn
qfqimrXig2jA/DBfFdzV/4or1/EsA/Bfd+4FBrqelv71O9FHnUZkbgQw3j2s47YB
KLmSTOK/RGazG1LpGUXacYguyGvlPQvrcx28oIGy9FlakcdVqA3jJpLkwUSKTrJ1
cgV+0gw1lTRb22Z+aGM/LF8yw5O1t5EjaVAe4oiRO8IYH24KfZFokClCxBtQvhyU
ro6pAA5seEvtVeJ7hV+M3tdPSz6ekFLjZkfCDyWd0h2CMFtTwLCseXTWs/vdD9Cb
+ZcY6BGEsRI0KQ88l/VDCHndmUeSsl5ml/260UeuaCo8myfUP0ViA3IRVqZP8pJz
KXrlPAM58inNqxoiz72EmwddhG/Av/OScNoqMWuh5Cuq7mCUjZC3WAe93likx61P
vcWE7TtozSs7b2t3j6QWaS0HRRHuwSKGNjzRk6PeFodBbNVA4Ux8KlS28RfBLccP
OctL4syH0OKt09XUTviDm8m40tefNxuTVp8jTEq/rLfI0zc7VgDs5mR+3Sac9uIb
kpDKB7JHj02NaUoSObqdGodOT6yWPoDzl8mLYgmvYC9sn0hxOyAZdkJ0YVXXn1bi
zu4tlpspt17zLdeM+HQiINzj/eb/witZS7tIZcPuLABkRgxTNePWuLbVvHs8W/XN
fbRVyOQ/U3LHmGsOuEvCIcahtECMP0oiISEbSN6Hw0dbs7hUelSbjC9t9ZcSDY1t
6WnzsYD/c7xxM+4hszjvmVHiUl7hakiGnCUHOSsQIZGwB0P2b3jQkZzsS4hhFZ9G
D/E0Gwt+NbI8tLCHWhouk0t3M4d823AxpXs+apKpQpEXsXo3u/hP2aCKl6wldxu8
1f+m4AIVXlu7y7DRmj628JZesNobxEVO+5cWhstS2WYkkmPvSqQ5Zl68nFv/lCfR
Z7LcxpDOn7oR1a+OR0L3Bmqxd5LQ2eDc0Ylqq05n2m51NrGgvud7CiXp5cNdTG8X
gZqyt/sNu/Wd0kp5UyGCpojSqXcbkFeYtLJ3asjTo9otFITcWjP4FRTyCCP4CnHb
WjIMD3KQT1Z2fPpN+nSNduIz5QgwLl/2EQLTR4gw0tH3Hy7mo/C0Qn1jqD1YpbZy
iHp0LPwFvASfqPxNomoYEmp4VAGPJ9GhSM8b0N/QNvyjOpob7hb4ebjH4dTY2fI+
sj9OuT/LyeMiDLLOLK0yAudFI7IF3S1GEhD5txcTzyl1RP9qtz37JDm/W28+iD2x
Cvz9++SuxMUBA4ndjOw2VVZ2g4hAQr2Rysy39kw9OGwTb4Fyle7UTb+GyG5XlUkj
COchpjy3CssUUhXl7ORn7b1SFQeLJeq/jX3w0K0g2vysRFT6Mm7tXY2DPkqnvWe1
rZ1Qk3Fj+pJt38UHvMTWnTa0bM+0Sd0ok0/ODkvY1rhACrbEBnHF4XRLfhyuLrVN
LyZQ8ukxsio2cM+gcaLumNgPIJL0aty+1gVtzm6SX8tKTWKJ6F8YHxugFgHWRIhB
iqScHxw0uiivggJKz1liYrGeA9IJSykxTQH8FrR7pXCEz3U9a4WIEo2GGZqYfIbq
NTspoyIK86DTahogv7IV/T+8FFJg/C+0y2J6WNUe50jgf/QfOloKTGXj493IDc6c
KrnGvKtMD1CesM/fJBL7s0FdTKjRjba8n0FklrFvSC9opLxVCnvQpKnBxU8kgc+H
RHQ8x8ZHAv6ergMlG6TECdx4J49lL2L0dPGYMEMrNyJKG9JFmF9p/3/pbg8lrwB4
3VPG8yK7n/zKuACxBRr/6md1FVVQ/QBFekR4bTuDH9bCvPNxF5rqCgvbY8ZhtaCJ
GnwxperfJcPHAWp6ovp5Cxlpf4Xq/SPbwE0ZElnMDrYOsQfWktetSXdTAo/nLFTF
moGR3gsk4Xupvs9xvKrGe635jmcCChI4GXGSD4sGQlnkAjAH+VCMD1EfXO1tp5MD
GbJdW5et1y67qvqRtv38vmiCUDLLLuJKNZVy9k3KL0TLcvZTybRBl1c8iAShh//P
q5FQSvcwvsu73YJ3hvoZq+ZdKbIB627n+S4G1dczGNdBulLZi2BcUBzodFXnb/LZ
4kcPCSPnhPpJmzB8jZNs1PTBYDQd8fQClxk26JOf29Qmib8bAXPq5Yz5PCqHkwyy
CdMFKQaalUuvif/57kfFF8cN78+FELhCgStSZpEal28R4O+Js7M8Ah03DKmUTnFO
RlUpiNr/RJ4e7PJm8ddhz0qZGsIH7wwh4+xIJvubdGA08c0Gfnd/O+77G8062UbD
6TtIYTkkIa1nyyMfqZVhzUPKh3h1+61hzqiXkzalFbvui7kzrZdyCDJh10Gf0SJD
9HRmNR7Mk64YAO82+IYrxLhwmR6wD8IoLBBs8s41mBxMtjCMDvnmKxEaA/1LeMV6
kWq82LpSykfISyl1IFDEvT19b3umyC9AdHtgyzv9APkDen8urv4d2jNwW7Hnlzsl
gGdb3l9hemygz3XXwA1A5P5ClfWWxob89E7SAL9m2xi/lasdwQJh4QDqWVA3U05x
SvwtEGfalh+OBAFfElMJJX2JLiDx6OyPWI15fSYx2J4UtczbDjeWT71UY6znWPVj
f4TrJSpEHiJ8T2pKV+U1ONDi+BCyiAuuttvmje4wEsnU/gPaCEe/AT7g4TLihxUg
LpEKRIP/WK9ucPP0nPR1K6RFcVSLmS9b/rmZjBWshVCGBoL3k7PB84lxAdAIF4H4
p5WFAaeg97fAmv2LPlx+cwMhHbVWgTMm+nz4i/pEmlwpvJ1kqzgOA47Pq+5uhj+i
L8UWaVe0BYc0usr+wEp8WTmiDLj5noHiaNi28JLyq1HR1AxWzGPgPSXZ6Uvv9sul
DEXiD1SGMM4KVQlYvDdXOkBlsfUTCRllu8WlkLkpbPPRdZGSe9p9UmeCAmIpDEpG
I3gn99q9DZzi8wdNUukVepqRTP0ziJxFzRMbiHiigpFzBvSKPNn7g9K0n57JbTvP
LiWbjB5uW8taJ8WD9FHfWh7tfg1roMvHMtn7m58PUcFvyYwn5PlanAWAqkUiWQo7
rqD8QqS3ZvZ2HB12rW0x3klNWkqg0fZpzNhYHipp4fWg/lw5QhXWki0B+flY0GwH
pyo7Kbmng4lOHbu0VRSUmRN37VDBtAbbR/b4hhQC5RRZJwMx+4jrGI5pJHKHTzrw
2/A82eNVpuBMz0lvIFKMDT4WW6DTiin4dj8RwiQecNsrjv8p5Re1jafmuWJefE4i
5VOw+U8okUgwFabuWqsVxgZima3S5Qi5EdqktllpJv65yBsHJQW8NaxcQIEVSxQa
3E1BYr9Nn3PnW0P47KdSUywbEnLce/2DjZDoB/BiYAToQKbI69+rmc4WQUtYoN2i
LnFWrtxmHCcwXHJzIw5HgxJl7srLTNPodByICCL952QwsT+Lwvf+V2QVY0uvQ6uT
Y0qTp283EErNLJNae/H2IwKsxxjvn7sF0oASEHzDMaUmsTGSURxidkqrLV5TwX81
nBIn2tbOyDRKtHwR3yyErg84RrNpn/8xbJ2XXSZxtTz1cNqZmb8HsPOHiCrmSK80
FoTkDhtqbCjT/r+DFt4j7ISQMVPaSks6ekKOMSWU4YUu/ywYRhjrEqdySImdI4Wt
wzzEkPCFP+0QxmH9HV5hNdyMc+RG331sjRq6nNAWJXf867JbAsILlo694/DL7mN/
aKIzysEHQk5h+hbQwHdclG+SYrjjsh87y+ibXG0XyYE5R06ZK6D5kr2Cxr80H5gk
7zwtLyxEH5hg2hK7cEtekvg2eq2xrK3OQT1g7VXCI0K26U3G0dRmaleFFJm3I+Qt
QXXF5vO2Eti72xyi+7uay47fiDSFSThG7t49xLDl7xFjNf0uZVl3UscgeAdhRWpB
YzZ7yWhkl6hTj9NTD11M5hBtf+vWTP+Pv7nGrik3P4vlBDlY9FibVBRWIhFj/L+J
VgrVcIhlC9W40PSuDAG4B4pxdVCxiQl/H6GszTgAedClFmtn+kbAXmXEi6oLpnGW
bsOmHz6K2hNggGIsPCBN/19du/RE20xP/DqBPKd6YLv+F/6yx8djucFbkEpRbLa8
1+i4im8H2/mNONBG5lMfPOSdfBbgvyhm0yJErlUyZHRfbyK75F/dR1EtBIdZd3C5
pE1fEznDJ0VqkFgLfBX+ypEx7BwFS8EP8Bkw0TMYuWrA/DiiTe6AydqV1oKpEtMr
TaeA0vaG4GYygEvZZDyNhdESkLqHwzHblAXKRGfVejaOOgY2CO5vSpVvWUlrYNpw
hvyajLrGy2CPREIzIZAmDiBM9Z1rfUYyPb7jjKjMbJdqCV9acrbwMesOCtnKSWDg
7LJk3EzF0I5GZMzmRIa1A8jXgv6JJHF4HRgBvf2+cZDRxr8gHsBD+5+aCCPdgZgj
tyHwEtraqHNl2YhY63LG9lBhwY8YR602LvA98NqZQI5Jwf///myq0TCHwYY20psk
pXF8+63D9EWfHn/CHU0p/SZRa1clkoAMZb/G5ugEHK3i8iBJYxjZBz7d8qQNvwtc
7iONmHInURkhvQaytrcOl5YRcSjhkbLYGagb2KRtF6pmgJMkozRCFS0BmRQUiuUy
qAgdH6yurbPVrbCC1GbRS5j57wlioICciibutDGKsoFXFYvkYTozvXAn/Nta/HG9
tWdte6UJFdbot4TiUCsx1W+Aty6WfVChEKaVlvQjKS1y+hqt+IKzZ52J4WURGk/Z
gX//iKYxaWVvL0a8Pe2KCGU8AMx1dvW2iTOaJWcM4YFq9BWjplYKNS3k86hQsz2r
CNxCWjY7swlyNwkQwMOecB3SP7h9/mZLrAiD9NXzCZueUv3qRGjHevm7imB7eie6
96jONVPZ8ji0rXrWyWhhUjuh6WCKM5iwlmiezvQUgmtnuCi71rkSyvbmMxyd31Po
6ptWe8K5p3lulQQR0dTOuNieMg1ISNIjLLMIAwP4dKr9QgEbcL/Mfj5VO92s7hYV
7BpYo6AcEkuHes4ZWfq17XRUKnfnBZCKTDiFa22S8EP7J0+oISjCE6nT7WXX0r5Q
SkqjssKpUfyloijGMmivA8cEhtMdazgOCzf9WB621jMym6jdTyFS7nZa1VGjm2QC
`protect end_protected