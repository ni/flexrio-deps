`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6848 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzrMQZYQafMf450Vd7e3SzCsnf1M6a70to4T10+9i8h5u
8fsmjq07M/elXXW9qKWaQSKDNoQeoxV7kMxt9Z/8wYmis4InnH2iRrviucJ9T8wX
T+mIQzWqF7SwP2W7NRico4Gup0R+4QBURbt+535zvaED/EREUlsQEfl7WrvXXGF6
i8ZfEZX/P6GUnBF1im35NLgkh+gy2cQGqb9QgyFFEQE4TNp+VfXCKKz4ZyJ4tE9m
D+IczNNJxTk+9gxEA9Zr/ElwYNWhfIW7nCiBFFgZkSR+sI4Jw5N02ROIxmSZScTC
chIm6Z/B0tI23Jz3mTaZ39VwtASiBzlQvftXht3VyWb8E61l2Vq01FnNKt+4+nRO
xmQerFSBQt3FNe1aFR6Fv6qDuJZ94wbxhYFg1qc+wutrsOdF7J1qTPOFhqkLqvyk
NRhDQPy+nX+Urnw0G30u78jLZqTic/BWPrh3VKpmzqtLLa2fiC3zUUX5dLK5qFwB
3Hn1k+Fo7Gibyrs9cRm02rQiztKlN2kIfE5YXQFHJaOwz6hsC2bB48l/h07aDSe4
uuXIZe2ifW2yDfQLTAJe7HgzZAJQ/iNT8Irxvw77On1AyFu5/XcSCHN/4PlhBAyf
eqpx/CAEftI0sf1n+FfYszF4BwP0qsfC9r16TfUCThaOE9ln55KnZd81g8imO3lV
8/uNZiT2oPXwJavEQcmD5lsEMF0zDxaNllXDfIHQPEoX9j8cN/6bliPHcTf+e6uS
sx44aQ8w3vB9+8hYR561mDk+2uj7Y2KpMgVR8fFPr/x6y7XitkDbFhv2/uu9CbMn
P5jOkg1B1QN8PyIc4rJAJ0CVocdHM1Y0FzdMU7MVnfKFNRR6Hl5tLhdywxeh1bZv
KECsEQB2B0bVSS9iHsG5+9G6khHlzZc2k4kx0yAeo63MaoZYuN9YiSnHNyx6eNck
ZyOIF6kJoMhDNZoVXT2x46dUYGYmpsTRR0cEaMvTLf+KvofeyviRVhkYT8O1MWVz
OvgNT0BCnnprYGLC5Cd5Fv/w8R9uYkgMUFa02sXlfGXFP8/EG7+guerWel2EXpCm
wKuqRdbbmvCdnSnyhOSPAUWI/32EZGnm/LpvT+ai/qR870YFQA7cYmEsjJrRmVdE
CVc8xCLlGYWhAEGL0gkOu6rsiEAx3cEKZgwywKvCHdgjoDgK6H2zNvkAYctMKpbD
1Sp/svMDYX7CTHQsXymnw4CvYVoxSqMy/ZfKHp/+XyLQgcYgSjpmt3QHP68sJBW+
/LZshO8WeQVwCIx7g/LCwlc+SF4PSQ+6I7kqqk4s4r0jEuhAG6YogwD/Uzn3Fi9R
00Awrxj12qBbnN6QNZq+NuRrsxrfvj84RaLBae53EVtQip2Hdl+zluxJUtJKBr4V
BiogBJFhd7YexOpXxUERpZFcPhGfKLBjGx4JpwssnfmWpUQZr4nbuOONYD1uBOLL
YIrYbkbhscjfFGg7OuMmryYiRszbEGgit6jpFbEABnQoCybMoiByHBkMfMx04+sd
D5KDzHNErruQCmxj0y0mI/g8lrL3LEMf7LW4hLCQMVvqFqMv0j0T6Aim/WisUaM/
6gvEwvTI8wK7kDU1H1Dbl+XuJ5Gr/rti7GJfgFhKrfXhXSWUjSJS9ZJdO74cQDIF
fukalZZy4zM5F7bFQopP+NvkxwWseYzHm6fkCdH7MCSDNG3GGK5xTteMVHHuzacA
9luA3Y7NtnnBWRgfM8vveWB69uCbx/8yHhlTHhIaMXwXh6Yqs7xN/8lNGYS+cS5l
MeXj7XuDa+CrZXkX5dyi/9u2e3BKdXd5B7L0RDIBs2NRgfeuoXUtIg2eZh+fMCNQ
Z7we79Ols3oxG8NsDnbuAuF+1ICD5oWjJ6yhCmmCPu/ipzaaG33eIxI9v3lnXh1Y
nMWlXZCnL68PEnb2NHhehtx2vk2wJEIhoyVbN5N+uVVS+2gJefbRe0dd7sJmLEmL
pGhTbLBpIILkazsLNNpPBx/FzpBYmfAddOPbOnnpSwTfZoSKkQG0GZ+Ijos56imr
OpFb+NE7q/+uCMFcLBBul5SSwDxqwveUz81A7dCS2nubUhkmC6GNc6Dd3kJok64H
yqyioHfbRykQhYnaDmToo4ly8iWX7BdR1TdMEGQ0C9E9uf+MB+0N71EGgujQghhX
q4+5taewqr6zFpz+9pyo+EkpbOsLYxvERL8NiG53Vn0fcN/USeIfu89YDNnvILOA
R+fCgCo9xUNh4yfvcG/vWnl+N4ASk6dENNO0mFsKTwKEQZ4S5Xs0I8+ec7kiEoyN
iehci8StASBeLxUA2zZwYUTZoWVITjGN3q/jn00EAfJ3F3mAnWhby1H13+C/xusZ
es7f439Z+O9+7TEuwNCB480kTJSSuAiyn2n3W83vVhzZrtRorhx7RJMS9wnPhp08
cG+ekrpP0L2rK/BfFhwWvlry6h6m2oH7/1r1vKr9xTW9UNSsSumKoFdc2BMBycTJ
l1Xy1OqSOPuxOzGypk6N4mxCAOdMCauJQb/HKHpgdfhthnnS7VZzC4jZjcy/Bux1
bdcobom5aDIzpgn2i57+oUcOf+HnGHfat0sharoUV6RtJwpe2VS6S8M7+Fhc72SX
XnU3TBcCgbNGZH2ae9ZQzb7Mf6AtYHtOlOmoGVt0AtH7Qx4JfyQoz77r9Ly17w+M
MNFHErSMy2S7oAB05TRGsAiLy7LZsHWQHbwZkA9VDhbDjQbmWhNVRHGqiQdBcie6
OG9QpS8UGglT/tjGd4u3JMYAk/SpOZn1FiDVIcd1y0AMzn9U4CTNvt5LrP4OnF/t
8G6+YpJXJFKh5B1WVpfEkX/RJF3rkmvhm5gAhuyftzZvWviT/TxRtvSye6GG9yRA
RjDJtR9FVxqyjAdjMrhYvhx8Wezgzzp+QNHq3BglXGJ/xe4De0KKMHvly+rRX2BZ
O4MbH//QEUZzM2M4P9uL8RBBkyQi1MKZLt0qbJs+JkR1I+2UMLMl5QJ8j37vS3RG
St/tV2YQa0qJOm/Si+w/vR7m1K9E8dLgg++0GVdvQQNWbznvpueKKCojzIQyVHX+
8Qr4FDVPpME7QuRooTz7RtHWwoFm6liu9Z9iaHJB7abfU5I9zF4wNyYtdexpntbr
KUtVHtiWvnzvFtpjs9Njd1yDGbmiNLD+DTLLa3rYfFZfIH935BOy9Euc+TlfXJ6z
ne6GdFDBPa84Vm1WZfgBxk8rjvxBvAtjkVybH3C4YWeqhlbRLehGLq3i91UtPeLd
eiCmWy94SrYu4tuqO/teirfFxGsf3B49ClF2GmyePR+p9RlXRKMpkZJzTFjJkPS/
FZIz+NFolWYiFanTnq/F3Xe0+1JS5W1nGGhk8UwTS2z65vxo5RJ5fpbLaULYP9/i
T3CeJVAfSuMx5vbgofSl0xWiqRGew+80Jz5LE3QFukb6J/ZCLXGQXu1aNBJZuXKo
YPj4svGhQl9XfVvFqIqiLzx0DBzUusKTXk2fviCGoSEyk9jOJ+9bdK7Ujm6y4JEH
Inetff/ZN2YCtKu/C+O6sKF1ST5b2nvQZo1jjZcVICwzNLuEAe/CsFotVMGb9FTr
Ude7BFKaWa3R1L3wXf0AhtvPkbXMT5eBgvXd1b3Yue8koOo1OqR8eteXijg37ivG
MN3cmtyw19bMbe+k/HlfHZ7KsmvncK7F92hBkxcbIE3r/0P+CgVbjJVN7kxxPlaU
NWUW56/HxNThj1P1kjh06VE0MAeelqlPafv7LFpH5zmpHA95FEq3nEBeeeO8ynOZ
SePDehkhcFszjkhkEK6hRYKlfkteRbQfHZUavTl0zvQJ/cdEreiJWs9BpF1RLcJ+
ACYmLerWX3xMShUWXLPGP5Zp6a55VboGTwLYpfeQ9y+Ksv5ktE+jIKdk1V1ulIWv
/rXHy/Y3X39/uYP/llLq0whpplRtuTGMWYIva+x9ZzNgR8JpKkpJ5xPAmfgvWWK3
v/H0XFh6U9EuBo1mZlXBfOyl52OM632/6XqUAyh+6CO/8goZmPO8G0N016VG98Ta
hsXi2ws7a0wruo31PzZF5i3f+73zd/WOsvHof8dlYO91NQ0RglHBVr1ml8ywdPuK
hUUluLKTOTQWsxZS8rYdjDm928qAk3nhHJkGqMopBCOve2iX5JOLVYplnbOjU9Pk
fyIXY99t5xub6utoofYZMF3kpNTmP55wtlJMtHRdOqAsMVpX7gD3F1KGhi+1jm0v
TSaGScWHFCPLoPz2xwW18RiR4pz9ESzyuBKh/MJhqr1osvXRdDkZZsS8L1mLERRg
5uJ+nrgrZF32m7tWsU1qhUnoqG1ZrSu9oZqATR6msl/OiSUmvQ5m74ox3OyrCyO4
k4B9l99NEVg3yZaqiXr6n9xXXRc6gcvgZLPQCqjUokg7so4PPrL7cibm9orW6s2N
seqxL6HustTsD9PbeUcV+Bw/plITeo8nZ8jb0xjTv10bDcj8OvNq3+HcbLhoXxIg
OHNqsQQTwid74KmhUmlVweYhRiyAQbQ65Q7gk0lIyNkWE+2v9T+/8lSdmN8jlsxR
3Plvo+uhlIyu9KcGvYQo/ycWsZP/kkJyasICeFHfRvIRKV0xl4BNibuwJqjBhVVg
6ExmIBIey2l5e7Juy5qSQcLoV+hxWfENYCBiVJz1ScsV140U49uFnAm3AbSYUN3z
4uJFQXcp1d1uacABQjXAHctahb/zh94YjSlu+BiKfKc22rT4UNo5LDPA04VpmQeP
YD7B1KJxUZgpP/vJk57SG5WrkwUfIuxrAeaCD7UPOCOmeNWFcCiZug34SgBhWpBW
XOvP3cOSZP76M+ujY0u6f2H8ti5bTYBNGBTswhTGLzXUvOZh3mQzjY0q/wVT45Ap
ZMqm1oXyGAbNk0piKj+dvjF+56xKIQ9UPS1Yydi1FFk5OIPRhrfsyw3JZyGe91R4
e43m15EIVQdBw49Xoujjke3301EZ1PgUtc0UofU1l9czwJbvWvj6898rRQsqEAqz
D5a7eoOCT9UAbB9/iJgtBGy5tAyjk8yM+iT1jG9okzoGa8vKo3xqQUo99/e95ISm
PdE1tj6q3EHBboeCxjFb5OJjMJtBU5QAeqc2fWE7negPS3hhKBPPO6T2yu1nah3I
uysYeNgbrAJ0m56k9PQ353F5zov4R0XoXb1iZvRxxTtUKgTfxq1rLKpgMRaF+WnK
9yXHiuk5bN2n7XJEMx1mXx+22mUTbWKI7AD08CNPp5ysPtbIWKYB1mTjLvO8GZqz
HZ/cXLNWM4/bOh5ENUQzEOEJm6t+QuSrzrD8zGe+veLqN5/UIjqIGd1+97SqAbSL
lOObwa6LlHBL4wk1jjTTrLAk0mnCX36iQkJNxsFhWXrLATxo22LRusuSfTEVMXDp
ftL4exhRFx21FofOJRRZjKrVW+yO3e1smmJsHJPsuME7OuowJT5lj+uDUPTrx259
F7AN67cBgIC37oBIs+5XcZ++OsB5OT460kzPdo912ZX+nhjG+uCTaYC/RcC7ngRI
RjADNh7VMKlUOVm3I1lBbf0fcTkJYrmcw6I2pXla1OrhhrMGtN282BLKNS1DCZYp
TYUJz166SAi4XUBHTaoyB74QO0GkW+Q9f4gXrNR/T9lpvL6sberxdOmWZo8b6Ym2
FH/g+gsLhfR7bA6Ht9ASnIAwtUAuKuH8G9KjRvZYnjyvD6bGwf0Q2bsuCL7BEOBD
1QceOi87hB1CQnZ4Qq+6T2LVAIg8zNnJxOi83ZPA1zvLeh3Q5EEtG5FT/l66m00f
HcyOLKabfbGGoFh+jUlzUzG0DAoYm4PyrCrcfPhQZ0ztSmT5Ebs+ELfM3kZDa+H2
0EsWNKATae8kBkeK/3g5RJYmD2DqC94zZ7IDX4mnFLYI/cHPAulTIuANNDe4b6UZ
yx7RRQZSFz2CA13KfQpkoFDU++NtQ7UgBwA/bms2XSvj1DWStrInu1b+CX6zyjeb
4qnGDKC5+LUSYDYo/ZiZSdguBsZKythI8ABVeTgtGOrXM+pMOnV7fgildp40fmY/
jD/hcrBSGfnAv6jdbQ0FahQtOEtMcbsqUnTY8Z3sbgHNmZD2H1CwTlRDYKHB4C/Q
V1Za6VA++0XiZZLtXo3nlYEq9C7qv8dcMRd5RSRXMOos3PeqxPmxYP6TIaAv9pV/
5qiy7qyblYid7JRDE3/nkleVVWIrkEarjEToHWVLZlL03OX0vKMeF7zXLrdx4PQv
CeyorTcWNwwY5OXTRLB4WasTuaO50FlmmlcmlqeZ2ZLIH1MW6wUZI9DOVrxeA7es
sFSSkUF26q0ek7ROD1UJ9HZ/URfiTacF8YcBh0uedEbvQwTUmooApgy7JzKA0fQW
GTyav9hYwb4urPdp9wvbDpJ4U7AJX7HscayA084gOw5MvgNrwfCfxgO7ehAvKiQU
c2/M6/Pul7sqsz6tONdxTmsWBKHT+0o/YT2cz2yH9zOejsxGGp5WZbaCdjK6oWVG
X480BagzIVArtkX8Q8PftAyGScunF7HDTeAhe1ScOfLyXh8IHEeZpo5fk9HRNs83
zJ3qqy7AdmYBAUHACjEtuNvfZsBVmMqtso5k6uEU+HkSs8s5R9aO5AL2a7KM+bBM
8TMCZruHWRKA9IWiu7kym4f/mD9Y2IB8qgmNkAmWu/WbhHLqv3DhC4f+TUsU8cL7
SNDe3xayje0nuDWu+ujikh1afyPuN3tMJw5AS2Jujgp+X4LTMHQ/I7L+SsuEYEzr
9SP0jb2UnGgphzyleYSPQuufFYH+FtWTjmkiN5ztiY0VvQIK6h4G/uXbpbPLxjdZ
t6wSJEodr17Bn7R+/RugUYKk/IHoyRMe/jtwzZTJdWNyx3y4s3+AP3OWRSAnJPCW
xT5/CYJU4Bb8zziAtlAoC0CihPbc5YkD1ri/0e0oLudaUgGFglE7ifTZJMBwEvK5
HwWZeWStEjqdtu38fHumK8SAHT1ef5Uy1OrnEM4UFKXhhck7EaRYfZhql4V4xHTN
6WE1t+ZJf12Q2EZUIbUYDdNEVSv3Is+YWtrTXybOjJJlMJ6MjvrgVv2h2eFI2i1k
ZaWvvPBMfFDGzpsBn7XPeRXsk37wPKAhoSVSC2bFsw6O16C96MJUjwPUvj1UTSXf
CUfx+eh2DXP/gx642S3jkC+Vx8fkgh4AgAmFLCVvUpFt8M4aPXekD3W9ftwzCARS
5ZUx08Lmdfnp0mzKoCeklYzB0UiAsDU77zMkp7ONSz0eoUZn0APFHZYvXpZxrq04
RNfZvq1njSwPzfBcJ9UAmnbTKHj3FfzcwRrPqOiQf/sWmH/l4FSbtfb16RwQgb9X
B8WQuYdnd5CC60aDyYmRrYTn9LfINIF3z0TsEw2jp93DfWnL5O3K9V1RftbO8nDA
ZdRWGOEMofAGXys2Rie+RyT5ocI+zQedQFN48f97xDjKS2yqX5ioqybZs/ciQ5UO
+NaDVp5iTyZxMMz7fHSGT/zMtHFf/drCiHB1BZHuOYfChFTz2nZXxLnP27dCuPJ1
gY2XKsnBq03JCWbS+n1DYQZFh9HlfgU25jm1GEHvTik48JsLf/IGbiiAvjGlu/f1
4ZQ6f326eRQ111X9+1NwNeKbYBMWQeRlY6sGIGhVIBNdTCssF284phyL5LOUXWHB
4bumTcolAN4TZpjuduv3RyydlsDnEJttEvKFIjD2hUhdWJMvp1+zgfltBukKua3f
5iJFJSaZjsl+KFxsyjYGznQkQCC/zEjlhJQxk5WTF3NS6ZRS5X6xOPqb6X10aR55
GQqgl6GhbQ3RtG+1vmjsIYeXS+sz1IeHlw3riZ987MhcY6zpb0dBovPaarsWls3T
hYkPMajMrdIbLmQs8DF67xX6dSohNuHpX2qn6ONIr4IGT/CR9gFbYBQM17iyPmqU
5fZcLA/pi9JXB3b0q2QTGAHkZVae8rVoQkfxhMtNw9l22wCQvLGl+6f/lP3rK+dn
WE+uY8P2nxAibgSMHgsaQHsq6K8/dKdPWH8bv3Obreok/lEWjszdMpZ3KVpsJO2C
pcPG9rJbkF5NmfAxcca/7XkJzIoIkVVaQx9VNS9Bj7D0NGMm6FSTGXARSCYxNfBx
vb1IXt7eF/tKvn7r2dynApZ6mzakcBqEHFoAwo/a9AMFae7S/H57gNLfg11Lkj4D
kuVky3FhXQSzdKgb74Xj3/fRHclmWhaeMSc0/+PeBf5jBT4BzXmYMnumiA19mD0B
1I2hk0Z+D3GAFRMwp0o3+AcWVWJxFYqcg5PzAqJU0pI4BM1fPWf66YyCXfcWcLQm
o5TDsJPVleWk8T6QO4yCzUnHYP7aizHxf9T01/pJRn4xtr1ZpHZCD5MqtkwBSzMB
PtmSlh53RUgkdzgHD/bGSGTFEPMrHvQQnsjO5Z30KyoEjOSaaJMVhUZXbQIG3ljm
kJoIxYwFMC0NOmY4f6K1CapjYrt6Yj0uaf/k54MQ2sc7f8HOpje3O2CxqDHvN2R0
giXerrBorMd9b5+cEwMTqpJGo0tB+1zfkVKD2cixfI7u632g7mJ0DGmOVcV368I6
NpYUdWk5pvcSriNz8MIzy0dYg7KWH5ryfP4p3/BOzIApcgAp1pMeICyVTv8ktBJn
ZtpDu3cJSIWrMq2Ux2cFbb08YHB56hofc0jgPy5g2cww4qJ7lnWiGYJpFjwKtAGI
Rkn4OVdUBSCH19XpHmX0rhU6T8Cb9rNZFRRPBPQS18yFItgrROhaVNaPjTS8R4eo
lDBFW9K4XQEJjgfXDGl7pR/y/0mxPbMX65dBOKxgKHCWqdTnyAzvw3BoiN75SSQ4
JZM4I8EbWFKbq/UhK5c7WhkX5vMujZU0Y/1AleunASzw2oq4Ryyd5OzV8kfPgr2l
HETbZo8of2IgRdk3ZUykH+HyrE79swhoHKeYtS4m5ZEJrBuK8p/CEBE2FTYddBCC
GCiLjSPBh1Uaw0zifXiPB7Cl0vZZk1DrNaDwS0i8BEHZtZjM9sKbvT7dC8txihJa
TvE4fOOMSNiN6pL3EHE4LU1Dt/V0MlyBk9bWbwnPTfk=
`protect end_protected