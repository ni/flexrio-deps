`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5408 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
XKfcKMLWLY4TfubABeEmfl7dfXW1qGE/uHJ6TxR3H93dsRTaWeW2BlbFotSwZ6on
+Hxa7TZyYKFpMXvPGNH/c4GDa2einwzS9PVj3oi+Qsg6F6vTgBjeCOSo1Qnbejq6
NmXdZ7dEXsFbntusL34lq0NV3aPkcuQbYjkKIwql7/ycn1y6wdS3n+QfoZgJ6TxG
7vWCghHQfn6/yZ3qPB9cn/1OzkjymU9mP8U7ADsJ+AEuGQyJ8LWRNwfEaQkPfGay
mvrzvWb6iEj/J5YnbT06fIZxcycEHjN5xt9FapoWPLJE9LgAa/OEsXEKzSXacuiH
USCLH95OTdT6hD1xYykbTcBt+rSn7NUvtUm7PqicXUe4KLrfloJVCLcHfNVVtI+j
tch06CWVaPpoR1UZrHHZcOQZKSs+n2/hoOgS/+RIR/boo7p4z7HWrMdisCz11BSC
uZo0Wm0hicA5NNsBfjlziIgzbFB0rsA9FHJ4XLUQHFxCFGS2mZNCs4+TosplX/Pi
KPJP9T52Z8RcHKbRp6Wc/iBTzc5FxhdkscceIAQ9eVM+CAfsouBbWdrt/043N2Sj
zhVmenfHFSKcYCK6YgvVMFtt2nqHjGynKGTPPWhS1jIPhlJ2e9MqWVOUhce2wfOW
pllpfk1ikBxyPBRmFe3bE5kVZijKP4cgXZpehj2tOvP14If0kWk2Zmp3l2H7YMZK
BF6T56RjJWhWldC56UtxXVQhM5K3k8IIdxpQa5B0gd8fPUIDN671QPGpKkduCrtt
u27tX4hXpAHy8LaBfnNc/9rp50FbgKWE/lX1k0UmnWtg/agzbFyyq5j1zW8B3tDg
vIEJfFBIM/uhr6VouBeT/Dez99veVPhqh98JG89MY3o7iJHr/mxTb1Dq5CXwtYQx
t3/9FfbJB7/wqtrp853nSuPecYutkMb7gcoV4NnL9w1YTgJIKaBj1Zl0lflaUqJm
6admR2fdcNKnQA1dEikDhLKrmGxx8qotlJK/+hrGJR0QwTkfe/q5LYvOCTjUeTMf
wcQCMFVYfcaQmzSg6XHdYENsHWnizL33H5rraaU6W7LW83XCPcKnR3zFL5f8rdyX
pRDgZSNecUvmk9rAZiZPIgnVDqhwc7GU9nwRrUjUAi3picdtGimIxu8lf1WyxBLt
YZwDQSKlMdiqcCxo/JZKPCddbfhvC15+4yslKtwVG3g9CosXpeUApzDBEwDF+FOw
r3UvFHa+f2Vr499EpDfK1UTBunr1btjbhrz/MrrZcqv7MUD5WhGKzDCFbtVXWR++
rytrY75NUt8q7jEUPToQ6G3P/BAUbe8uhDeu2N9QaXWXm89vPEAJpAtjVgI3Fmi5
m0h/CrrSA9ZyNIP2OCi4qoIKKp7N+v3xc3o6gkQ8oxkUvUXpJibxBnNMStbff4Va
dPyyAOf8VnbVfxbDz1I2FGiFV3IPomDx/JetRp2oI7Md/Sk4g/UNePVi/IGXEvzV
dUpL5WYHxqI2so3k4j7AFBJkJlKr094IzqCp0S6kSmNZRuX3lOWwxzG8y5wDtHzV
1LhJDzaB8Q28ONS1Y/mO3qzX2mVFQ4ASNbWbys9OIgfV/7G2XwCy7ZfvAXxyQ4pg
0MfPxsMxV+S/K7sXn2BiFms8sB5bnJWya0LoeDMT0I41JTwl61ERV69WnmSFwClT
7UMDatOY/yOtMMDKzc3x8vU7Qq1NwDNdRPAoFC4f/44ft1VDWpw0yBHMIldFg1gx
LzYQDAnDHSf9v9oFXbtlKBht3GBOhuXiocSV8kJn9K8cnWJN0zAgaw1ajhKLYbnP
iJq0cvaubyotPxihmHNiKPumMs+8RUF7mvRapHMJq7hQYUJpNnEwiNvOLJs8bEqK
YVg8MGjRaOdSMvG14i38DRyMcm5R+FOKsWfojyGeETeniXAMEEk4QVdmT+HZQn66
jMXT/w8nYv4M13AWK0Yjt0MoIP4yVlHNmD1zDWjtFdw4cRSHZPbRnRH6F5KFG5uK
X4NeQndXVbTlAfidxEg+M9mohO/dZ3gU57nxCO5sukakX2jW7LPjtOlLAuzDfRNN
cUZmRqA4p22fkq9WNvcLXmSv/f6xlY9eIs6uiAJdglIw0h40N99RknLHHx+U/au+
1w8s/SLNAifdJUC7xkXTSFmg5fxIEWhjWlO/I31+Q5+2mTn2nLqmj79JkUa2uxtH
DWI31sj1wfSzT8j+9Ue7M6IUriFU8buvdFfTbBgA0On9yJ6hxnJyRkfAd9DXqwMf
Ryr7qfV8UKHP0H5JsD3cJl5kcqTUpsX2FAFM2xRXJn5yuIy9feuodr1LKHXg6Wwg
vPbAvZjRVdHvaear8rMB83H776i9vLhPoCMhmMr3Zl/nBbv8/d8NWwAlcen3uWBC
pqKECLUIx9JbSm5ak9Ftwlcr2a8WgVXYIyGYlbhzGgaULI6IKaH94+vnwvXxx8uZ
iiNRfu9klOa/xsrTB+mg2OGRAqWBsvJ37Pux0qMJ5m9ktGjPdCKc9k8MrkYHUSst
xq4w3jW/MUOcNKhY3SE46WEcfKvMO4iHxQby313hkz76JO09MuOc7qECBxWzJQ+W
zcMviRPrUEfJkldVNYgkoORgLnoh6FyQ5zp/EtXdWZA5GAN34s4mCzZh02SkcO09
A/bizlE/eH0L1sfYmwgxzeGsZKOs4mrPMv5b89bEV4+xDg4vwZfy/jYKbGKEuQMI
ccLeJpEQasCFIv0VjzfpmFTZxWU0PNoNYR5dgRqMIjyBuUwaFPtDGeW9Irt7SW61
4a4NCJRosrFKKLnold8azbpAV46/fPi7AK/q5AaViMonx69nQ6uPTrfziAsl3ycW
WuakzA+2zWnNZ+KDwlw9o5GW+3Q3yUNJCcdNYw4UVSBbUSlEu8C1hZo0whvwxdRd
NA0ASxRIYsYnZ0p3NGjEM5diJxVxXUvaxSHWsayOyKy516K98YeCh7zfLa4zbrs4
oBbr9TrKkNOA9DSmgxbvEJlua5dKfFsbaWfd2s7LjPsiVywGf+x5+6sCPM9lOkAd
43oRByEcYkmxyxf20bvUj7BB+c/GBUd4Kllh02PXUB67iARxP06hZ3AxXsikU07J
CrUokC3c/j/e/ATWWFnzmxeQ4i5AG8XpIGaUfwLTaC9iaDD0rqTLNni+32yMHI+S
xvPMN2MYDUoxZi/AAOD2QRrt8wbVdBW9rkEd88pM+MO75noOnrj7pD8uHlO7faEh
IUoYWwK8uuVO+9zFr/0nk+zSjguymkUdwW32hx94cR+R4p6LSMwVmE4na3koOZAm
Hsw/MP/9CPbxs0x8sSETYmVuRLAC0FwXMN5ZgTFhDFLO3Tx3RjedPSqD1inE449/
6mUpq4M8NmTTriKHYxjdbwcwLOKx5uD4PpN9QE3T387AFYLahs97BVBqgpU0Ny9R
Xo5B8HThF0izLw+qVcBqCnbqLwCAWjbP7Kd/n0BiUuuT0Sw0Jmw0BM1uYtiOFcbN
Q3/nmtIbYIP3adAlnApsVSxYWXxFRghjSqQRAm6jQT9UhHn0clepqvmi7+oyd+wV
S//AXaC+YcTh9tVSowj02lPWqdxD98A/laHRq1F6n/z4Mpmc1qcE2Ah+IlPEOFiS
fjOhcyuOHdZ4zMqsEI2va/CumFnnM+ISxEczV4A0mQsaLRBvXo4NtchHSBftlSeb
fg0iC/36xE3RQC+5mzg52SkrStbnM5cTYkBADfClno/ByO6/OwREjQDck0bDe2RY
NXptqP2lsFYwHCaA/msgvC5bWZ6OmxLKN+1IDR1VLF1Ab5ia3lqBo1ls9Az5+GCj
iMM9k2xbQAFo8XQyX21lfLHJ2mkc/XGaR1CMyV0p3WlGGrsAL3ZqodB2rM0BWmUk
W5wwY0mFlavZNg8Amd1Uq7XhUc2wK/Y1jiMRAn81Fa9ZXI0aDPP687KoimwnvHJH
za6OFFu1aG1h+Vmk+tH22UFshbiO6dRnU2JQRGQ9jguHDkIwZ4wdvN595yee10vy
CShfb4DyqYtJLrm0GarQjvPydCq17EBMnRRqHUHqRobvnEQiubL7WHFBDMBB0y/H
knGCPXb6Lwqxi3DTGEwsjTIU39fbplbuSrnMtmJU5mQG9ZlD0iV7ZZYLHf4LYNOx
HHv0xC41mDdhVIfYaTBy271Z083wJCReJakh+xli4dJjbTZO+k+t3k8Ceqiuirh4
PLU9vkSiNEJGmJdGCK5PJfWu9V323f/MDTZYYkQ0FHGG7RQT0pWX29U4Aa70jy3e
HhG2rp0oOZpJlqJnQ01WXsTRq8ZxaxgshANwJNQC/5upIigZfQJVoJFSOQg9NEaQ
0OC/2PGHaSnP0AvQ14AQyFOYvQt5hZVpwUAxb4ZXkqsY2A85J7KhbAqL2HltC7y/
/vNLCS2lJ+r0gBuEyfJhrpVUYDM3JCPY4MK43zhKi6xPaq/EVjdKBjBfMNVcxSxa
utJeW3k+Rx+QBaT11ImlR+rm56esEK4XbO7rVkDMtejMYwyKLnl7ZL9IyFzsa20v
F9nRcvv8XcYvf4lkRHZ4CKVbdUM4OTSQfHGBlW3HXB+LVYMnzsAB5XZip0JPBC2x
BznIA9fbjoxCV6qs0Jk+ZRNoyNgf8jnFrwZLH+oJjlLml2Fbk4IE1jR4YLbvVBjH
gM5U+Ju65Ge3DV2sOHqv6zmwT1oyodbrjbK7urXBuXiLduhpvo3wqEci6JlLgow+
priJJmsny5dcmQ/w9gFH41BAbPcwEREn5SqbXpKKg5ANQVpQo3fcb33x1hOUrmeP
CvBYwgnM0ZPho7aMA6A2mzNkEshOkgfOp0M0AEgLa8wc7GBAqpr8ybocBzoASnL0
6czVdpKPQ0olReEvPrxEw7SgnD29cDMGZFY6XiZXQMrss1/X7j1XRlZa10inM1lV
9tsPM1VVfdltGYVhwE5ogbieR8spaWO4tjzJ4Ce5hIq7FpPI6jRqDEZxc/iQEF6e
9QHa6lXzy7qY5uD5TzWSaiBOnQyWRPmvwFmgXqCoMgexLQ0VMOhFSInjWiuwzS8g
ecnl1+HJi50Zvd7kQqw/TNUUFygBgc6dCDZ7ExnzNSRWJ1Ve3IQkPQVJmYGbGLYL
kulbOG/yVLnup5YDjnnTIV7LKsIBgn/seb8y8j7vql2tK8bpBZEChmK/YRBGNS8p
L6ElP4cqdOM6uuGGTZ/XZKx8mwM+sPNp38IyKHCvCt5jCTvtH1xjDA3MtAiMsLKb
Ioe7livYtHpZQYGXUxbozGtM05UVoI5/dkpPmMJIZRNNl8JRaWr3fT7NUDAQBYZv
8hU7HovA9kxFYVMCT07jTPjzFZLXvHA+maASeqe2unaBknlQ3d1IPzwm+l/WgXrf
aLwI4iwdkCyNsy+W+gTuNaHeDtMHR3YrRLVlU9d0aAsaudxo4MyjLH2oC0SmknWV
/RchvsNjnOSUNXvQEAiykDCeu7qNFpKE0QWGfn7NfSg4tcw4hnaD/0JPjdObjzxQ
J2r1MGX4wUZ2UK64GjCvQwYraIRafqN3J8FIVjzzXLwnBnUYyJOpuSKY4ijbUvou
/JCr5hfBx8XhUVDH/RXZp6b53buTAUDqcQyLIHJ3K8fZTqOIKw8mHUUuj+eCqgsh
CIzNum4NTxz33ov4vMPIisTvBeq5oMYGzjjNI9HHgb1GTzYsp4GOVU2urMUkqBrF
q90F3F2i0u2KkTE7v3fs80AR51/F5wVLtq5LKZZ/vqvgrZkG8Sb6jugXmbzOdugS
7Vbe7xlMsZSpkC8QcwNTAQgz2zI0XG49Fa+SYdQMOh2gHBl4EiMep5UhBQIi8eWY
r3usucTFK2uJfE+oLDQqRdZt+6A+ZpgftTKNkwfPO0Zo6FBQ1Np+hntkvxnPH6ak
IKn6wgqwY000kh4dcFL7u68s5lUYvAD8zmOnfGxHSOK0L9AMZ5mB8mEBveKepAi6
+D6l6IUl0u4L9U7L4FelDTtQdv6YuEN3McMwBUfOk/jDQZBEQ+jHc4Ij2mR4M/H7
SlskgjcLpXBAcETLD/L+dkQZrHGO0VqWiJnxErBntDGBLcgspKkMXxE6+Lt9Ouyy
0wC5cYgYfOoCMz/HpLLZCDUL8VF4w3jmRmBEJuGTKG5Sg7kANrnXMm2BqqO0HzAE
9ufH4rAjqWU6BVp3f1HdqsSfCXOVAluWBF+wmE8TdgtO4l1sm8QgC52Qih1WkOB6
CeQYgAg33PjjplPpK6QDEk+EGGvHYbbDBtr+mkCgWkM4vWzP/frujBFHDyX5bGBs
HBaWVRtsiMZWpb9QUE9q/0t5BnCk3A/OCP55zWWRJNCrSi5GDLTwfUEaNCX7GY3p
fmjjYmuHXeyjKK3fVi9KZThGmTMRTPEPDfyJs+vkXAL4D5BTR3Xa4I4OzqaWnDO7
rg0dnBycBNYonk6wuaFnKuz51v8Td4NIfUcRT9dv7DQMeDYpYw0YRQx+zfyeUQWK
PdaXiHt7uCT/EiaDTkN6CulMEkxhsDtfpBd16LJ/g1sfv229aURP/BMkAYTTCX79
2q2TY0529MUWxAG+CLAk2zQZeDZvLVO9LaRvudPcrgQqBtVuyio9zXtz+w5nEYTK
pwnhMsba8GFZ8F0jo5bjD8pMek1dNtSYPrkCVgy7YGtFnAPEqi0MoE/+Oqy42pAh
sBVyQZd47RukOC48mfLISl92O1PO/LqByQt88i5H0ZJl/0WFj5cJ6s3ZZr8TMQ/p
/0uAeqmbazw2t9mXNLWJWBGmu+9qZ/0cw2Yl6fK38t9AN61RH9ggWzyxWmewT/ZE
ZMDfQGGSLLWwniKzLqOUaPGpG+8sAWxqif2+YvWHeK+lszdwB6BQV2b1qy6ov6Kw
7PxKf/vWudw5qbkU/HdFhVSVy/U6lqOj7AxNZiePjwQMP54hnYtHbJmr4SHvPdNB
0XZ3v0gpVumr2PDAapSTdPHSiLmHZ+FZ6c3sy8Ha5cL8qEK5ALgtjOjIMVONqmRV
LOWBASpk2M1FC8V6fD3XII3dKjTE8wB9vwX6M7D/101AeD2PtTbi/adoWFTDJNi4
2MxF2TVIIAq1gVl/Pofwp+IaqyJ2up1k2EG897sxMof3gAa5ttQbdT2ID6iJhQNs
FD7dpQoLfK5T8109sZfIkTFlkSKuh2PiekxYDt/ESEE=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5408 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
8aCqQ2oUxf3QHZjuYP1t5OjsxBy/GOS+iraSqP+jOUUqJHNSRnXv2WxIb3CUWZqg
IQb885eLT1c+iwjnK40Sbp3d/I47Q2pq+zjtXwRVFkM1qKMdPIMrpZ9AMX7MuMsl
aztacOPLs2V2iTdwjuTLquFeXNlbR/HagebbLw2PQUMb9r+IHZIcZfYgB1bDBg2e
8CU0gCOnBaHvzqLPRSrVFWH/BZN9u5b7umT3L12Q/7tUMxQ8MOUg1Uda72gll5Ii
CGXBzRS1bqKtkYCmFgWFx0+3CpaenxbDxjvd1Bqm+70ohU6JdBZdeBiLqkDXv97+
wJBhrH428qlpKRkjr2V5TgdtpPraQp5whqm0qrgJuspvDENaHSYT6LGi4owcyJOV
D+bj57qIPBghm9tAWVePRZ757zZynD0qrmcPgAUo4ayUrJivhW4gbmp5+NoMspvh
HC84nk2n5n1jHK+1SJtrduZjyhfrZHF9bf/dZV+tgsbfdWXjiQMwUMVzYqAvtupY
ZsScEFFc4JQO+xo2qzx4N9iqTYm19/kY3FMrcc9rLhY/3To9VqyUREqxxBkY2YIj
i8ldT9CWJSbFniS2uo8YUityuOXB2dtwUDwAkn3bTFdqQTEg2CWaL/V9Jtas9bI9
bum3k40tyhrlbh0n3k7vqJMuv4gNGurjEmcBOs2la7U0GPvVHVKJAJrZd2jXF19w
jgR3VDZly/GsQgA6PGip0ZaNHzs2f3w5kwphLb9LhwjFVlf7G+gDMfeYiIcQ3V64
E4R0nEuhOGGr4mlCTMNP6YrWfy5zqd+44/HvJjtWVjRTaGMS13iIrbSHkpJC5AlT
4jMzBQ0nt3vq8kWT97PhDsfm6/NjvJwafHkDm7X23klA4Me1F2dKpSLu4pkei2Li
C6kE9/vzu3q99xlK2mxZz7dNpRaYByq2+ZWpysJf4UQluX/rKzZzrNM0HLUKHa3B
SsGTdkyT0RZN5URdMLZwE8LNe6cSTgDIIYAqm0vgX4jYMwOXPgW1o/v3CLCGdbP+
sbayULcXEBzMAPJio6IrQ0gGRhgbpMeqZ+p73+wBbZEyAcqeOs5zTpFiRQl2cNue
rBJ6CQbRm4ZVmYH4nQWytkUVIHcjpLtvXoMlLqkp5xa4CFDlk8AgKhLxce5cqwnr
O5ylQBnH2aQha1m54fqO9EqgjGpnU+rf319ArFe+dQRhAyuX1koLvWn6OagYVCPA
aANI5ZQ96X1HsBr0c8Lwd9dFnJPYVkWpXO60TKT/tor/OrwEngqYLuWXJBX/Nt+k
vY63MBtlDsTB+fO7h8zRCwLqdobBZEtvCgJiaH/zwtKg8DjRexY1ZFT741VFZj6Y
bz/pOe5UJ1eehj5FUGsezwAeerAPNJQkwx1FClp4hAeC+Nynrg2g4ezctTrpDYqI
5xhCCdsKFvdgc8fRwo5nbuxFev8/C5QpOvCEr/CIAfnos13XYw1auGR+s0UjuX8C
jW/d4C1CAAy4jPy8E+gq8dWaB/go7/+ohitY3MqMKH+DgXSqJNtjKgParCqzyOw3
HeOWFXEbvTFSf8ta0VVdki3L4KZGOu8p8LnUIL9PoSCcvI9CJqGjXHRLS6dIi0q5
04uTVFJmLxd0QM4JlZYS6mE36pTBzu496SxLSNBsoLjssmhcQF82j+h3RsUBySI4
WK0KU3JeDW+MOz/vbq5DEheT3WK0WpC+yNS/SNwEsKUZ4Zw6e+BJwyTo3wDyHX3J
AoQUAQ/RJVdtDOjd2CQ4vL/h5dScgciamLgJSWwwjIQCcra8v+9vZqppsAAMnmo9
hwG54oHNGIeJaPaLOtW+NznQN5gpl75YAVRgZoEPFxJpbrSUpG0Nz3fL15ad1ay3
9JgnR963olwWWMD40DOoKh8JCKWelVV5ZrdQM6Aa6csI3M0rH6d+w4W5PVcxjowd
QDG+dnFDGvZmv6DP0kCnA3G6WZM/ifz2vcfggLSWENPz83VoyhQw9ueiaTHu6t18
t5ZmybU7Ak0UWezWQ/fze6PzAQAX7MPqwueYtfUpTEpJ8MooMwIXyCOQKniN0USE
daaruI1LbkilPYrb8jmo6xOCUgAtgnlnVennMX1hHsN7Gr3LDjOnyysJ0MBMqeUw
BvVxa/d87W6ErFL49R+X6Dm6eXaHCNDnhSjzDnw1ZigiJl6rxHXr53warLxpyJ5+
zOo+510Jb0k008tgN7DNfqC9l2FbNrfbRxetwjigEN/gurxq96KrsZDC8O8edAw9
rVxisREU1kuzlJogXa+k3RDPlMzwDknHHO+alVZYeYxNkmBQCprehgx9M+A+eYEy
E/Y/nFEcMhcv6Hiv6Upmzj/hBaA07ff0hGL4U8e9I/PwrjmT3BGtnZ7YJJqoMMPr
98ICVBxaPjIOKNZK5SjWzXhNALEf6xn7pfH6nX3v8E+BWSvwavBQgPJNpS5ENex1
zpEjIo5IJGyOmrbcny3LtqZFJgnI7mbTUfPJGuTmPQLG32ENYEFThT7xV36LYvXu
nCy5vYDZ8YDHBAmA/bdqU1Cl+wFG02GL6Przf3PR02Q9lVFj7eAQ0TRDecNYoNra
qFMk2vs0e1fOLXN93tHTgr9eBs+tOIeATPisM2KTeB3Ciz9gikR0V/ddziJ5Lp7l
PK/JsAhLA+1Oy9IsuznElo0+m7tlyh0aMhDiGYT6mCzFCFiwx7f6vQOMCGR+E1ln
IVZLDw39dYF54YjusiTde8eToPrf8Oyq452bDCxJH7MYFyOLBVVd64Imv+OnO3Cu
dPjvw4j32CxoG8dr3B+dd5Qwi/sY2kTV6Y/5OhtCOJA0aaOLI58pRuW62tJPDvZJ
b/cZDSMrPVzl7HgaC6qreqVkVxL8yVLTUvQk1ONXahrzjWfrFQFNiBhWub7o7TFQ
jf3j+wIh8x/OwNBg/++8nshxDPkWd1dPydSLjf9bN3JhIJTvcCknq25j8vuX/OQV
/fDRUyb5/BKrcNNKIVQCyzz3L4wl/OTO6tu3tCuB1dVdgZBtCCzFVvKx+d6X0NI5
PVoTcp/rPxnXOJTkLy6zwsdmEbZ+YrhZIFCVz0w7br2bzFo5yLj06BqjxEA/I6N8
15Otw+VLkcWEbcPCpfrlHTgyXpQ3e6hvLGL3Y89/SZ7V/yiSnFwpdCoS2DrsHEQr
b9UncYSXGsT45vJFZyOsfW61Gj6S4OroK+u5DFIfmrO+mIiIyEvWeG82bLBWs+6P
w8RSYiyTItHaU/pY0zbXeBaL56K7wwilvjKWlwIeX7ptcjisj9ABya9pwzRGdBrG
toeVI3uJDgfcBxAzEDQJ/3fc6OVwrK3BLJ4ulxnogVOZ1yoBZneIhynwtmwy5uFk
mg8lYWEudG9huTSQhq7F2w//Haq/f4HN+WiDCQFs/hMWzxEQviQVQANWcm2RleqK
xIDQPPTMwlUw0hyfsb44dnmYztEdLPRX+R2IVvelPfY1rUTjF0Y6Cksdk/LWbuYl
cqH+Xt53GcLn4j02PzQrr8we6L2rP3UHRsfSRl0CgYSQPwe83ZHYDBn2jxykcPbr
qLGXF+WixkpCeOazqPogbHTmu2KWcqz5Ma0Hz2+1DXL9BqxGthHAIGhQ1gFzOIsL
sIS5jQVPzR4iahwfXNG4lU+i8CesbpzZ6rsuxAXoOVP8sdGBXvNL9GVR2QStmb13
XNrc+SnBJgBsPxaK37/T2v1YPSIOc6I8Fxd11wY8AR2WKA7uVATR2Gtf8vo6rKXD
N7u1SUIp8vH3164AfvvpThVM2sg8xyCNoXKI6in49UkSlJBQF+Arrx0opkDI5DJr
/EMekloqgZA2D5bw5jABRRK9zn91nkdTsCn8wfjMeXukoE2s3WgFILJgt5kUilBl
zkaqz34KCXQWE75oLpTJotKb8f0VC4Gj8hqsHPGvWiYcERKGB+phXmqzKJ2Khu9s
esvBmMVOgZyPHaiyX5ebC21wolWflfNB7eFUMQHequ0fffwkqzCQWvWr74Imhpn9
/HOAT0WA+TFkahWxTytuQuPY0JUTUXG9cfmUrDJcW1GVcIvfFd9APdoAPvHzs9iW
4xjGLwVEc4bcGFhy6cdL/0L4iUMcWn3UiYCSAbW/3SP7Lse4lxK8+4Ou+fJ3UKEL
UiRZiE4Xt111SNYMbM89usEbP8i8KW5nD+5TTvD9dnlf54kPSU36BSM2qSGMIQUL
4dBRmtjXJOXB5R1VpvcD2arrOPlu3uATraMxYDrROwmWCnZsiv83j+S0qqzkGKSw
aQeQ3ExXYrixmL/95SbLcuAHOVttHcrOJPoR2B5L0fh61508QzAJSUEQWjwtwlrZ
ZMBsySip4PuYsfezns7XSS5IguIcLzTbs/w02or002/ahMaG9G50hcMyeeoP9x1e
+h25QjU7P1kdETgKexXprN9fNteGnXN31zzMDCFMrkOR9bYAGXvVm8mEv7Smdmbc
6trggrldvGBSTmABPhC2lUZTbupxrR5Jx5IYvthF5C5vi+BxR+u7CgwqfDGH7E/b
5nwOk5J/MavDPJXMjSBFwR2/0vsrg3iPltvS9uJCB7B5sXgSJPpLRMjxzODyfi8s
Q/LoGrWxErowthEZG1FkyuC9d6nBzBDpiR7hzE/qAcgjaCX4FquoL2k99z4aHw66
JZiBGq2osBHMi5yuRq5Zh0kTFWRqkp2MPq7z3Ly7MuixdtsZzHfOHICYH3Z++uux
8dTy+lnZSU4hzqpy5r6ZhYMWgf9PuV4AmMNyqFNTCSewomPMc5MkJp8pPPV7Y8BX
2nqzOBzNiXUvYh5VT+mOBwZhAM3TEXbBaqtnrFk2edX4zmf/yvHM7wt5nH/uKMXk
2Nu7yiqJMyXriLBAlzqeuZe60tesTvZr+FzhH11yyXI195arOFI9D+PJ2AmOA9/y
ENDg1rxEn2c+vwKR3QGRwK3jXXfYhUKPED8qKw3j7XA8CqrvAT8HZ5PirI2LuaPn
SPqijEPdVAtExh948uB1JO4rkNCCtRjXqwhor+ih3KXoQRDpB6KjE6Zrdk5I9lcI
wY0HKOwwLaoH6xL1FkJTew04nNAphAakS7JL20tiyzzwtagmJ0LKneH9hZhtJUOW
lyx5s450+3Hn4HzWjzysViH1Hgtc+MwhoO5lIguUfdvRkfTXdEpurxKAzGUCi+4C
tNQyWvOcXiCZxFJK7jdallA/V8MTuEWRqt5vst5jFkqkSDsY2SGDBxT5emLoMzlm
Mq2TVoMe/U+SIiCVazznra1fufHJc3GpKtBoeYrJglDGjEKsqQub3Bfe/WKIFmPh
a/DQdAUJXi/b5pg/PsNnp+Cj99ddGqmnhbYBIq8CgypGtqItqOi09qNodR6Dbnt0
TME6jQeJXwvo4EeLPDseXdswL05Earq0AIokGUs5yfGBrsQ1naNdouBS2pARXV3I
Wtxbwjs/V/o3FoqGqByg+0FcEpECjXXXpoG7uAugnHLDj9GSvd+9SXBKBbKHAuyj
Xmu/RhW9wM2VSMPmMZhXeGkn3ELYxCkAeckH6Pzj9QH703Mwd9Q0itL3UxU7U9dC
D5TZUjzSfYWtiMjEuwEz/Gpmod3bQ6n8+xhQ/sovI+D/oZ1PVYfExDZGtkazFn4m
FKJgXmY8DxHh4QCXxyVgzjL1m1H6NA9VD5y5N36mYYVQb302bVE9Hye8SEqYGFjK
qnnIj4mycLQkby4PpAuEe4gnCfNs7fY2rp8DLh7aPLxItgfjjDihSNM1ca1+gxGt
X2GIM/T2TLMSQ9VYkHSdGUBwNoiDyCbXmTJZXhLrZnpgMm8v0GwaGQBQuF85Aa05
9jw7J6iwnpshgAQyxG7ZTajQ5u4oxgN5nM4jh9p9C+OEkWMBz9kZJg8uvDizcJwK
WzmJ62E6Qfmw3Jkou5DwkWno3vsvpi4k/3S2wHAXA+j/Wx4xEmqTaSVfBq1KW/KL
uUx+H4ofvgYmX9A9Tvc2Ccm4M9s067c7MiaasZrTNKjS1JFC7lrbs60l1O5PNroc
UMn+x2JPyE4tOR0QoWND0gacG3jtgme5PzVNxDCEsATgQKkBBGhMYaZP23V1DLRd
abO0GHEPiSWecPMSlmsAwaJuFvUnn0+MLf9Se+dRlVqI0CeEljZbq7p0mXNZTZx+
oI/oErDJYqpMYmcntNI/AGgluQO5pO5vCOU5S2HPZLwa+2KWjI2pqqTDEDFzHC8c
BwXIBL6P6Lej+UZCE6z7R7B9cK7GqPhJ29hGkWQqlcUSOmvTRt8tkWG/dw+nl2oa
uHWgRLM1bal1bsjcoixhCrJQDF5vXvnzKfKJS+IO1oiuzDA/I+zDOrRwVXpnXgaZ
j8rdOiEtgEtMQ6RW5hVrDJYfWiMG/qyLESRbefrioW5P4CEFSpfJRjBuQtj6FFKo
IsoIYdmo1ZKRlVrrX+tyB7OrhzJSav7hL11rBpZ9By/RZATZLrEvqVu2NyhUMq9W
Q4L3vD1Yfi0IfJFKlO2U/puZ/a0S0Vj0yvgvYfzCJ8ssFmV8ThsR1xbH2h7GuaOh
4zqXjshaiexpYPvqN8u9DKecRBaNLLMbmru9fBi1ifY4d8raN/A1DeR7GB8zr/06
4LADuR9aJ1mcpaECGqnuvXGrGkiSaQ9Bbl9eAMBy7Baun9Z3/DoS9l50B2xCFp0q
9UTWrqGh+0fyZhQZKHc5+O3EK1DX6au67gEcAe/yfYGV5uDlZuDeXfauy7cqzoYP
Pt5AzK7TvshsQVeY7AZL85e4NiU5KkHqfBnSEVDIHGonCX08IFNd3N3Al+rdHUaD
7uS5xEKwSGENsV2YjI+Wg0k4bSmj3/4yGNW2Gu0br0Js8UNR7V+V5RV6puiciTSj
DDSYLr6NZopeSjO0acEclDq3oypN4GNcXqYW77bfwhC7vu+unS6x+Pshb/49UMY9
FZyGLFtHRjEsB1ifwbqPto8KAzQfagT5e038mOl4E15iKhnIpKRdkuCtWSTcAjMr
D8FtHTMTgMoMt1O7Sbvzn1i2r1648UnXc/dT2JVKY49J/kAbKCHtrRffxOwTMN+Q
JGYlbDEn3hitHNZK7EXX7/FZS64C5V+2cZw9wgW3XMqm141r+VKBClCjjtZ4iMaA
p/uWq/CYLtRV+2gb0IgQ9jy9pKD6NN0yp7iaGN76Oe8=
>>>>>>> main
`protect end_protected