`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3824 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
L2bRNdr1lLBT0eERw3vGlI4eLEDE3nqq4kslHvE8qOZqmiEeOq5WqRg3sEl+ZMlG
I8YQ3aU9naZJ5oI7LpaYHL05j4EtOIKq0qMSS/zI6Y+EGiT6azZWdCD84yAVJqpQ
CMDqom8uu0TY3HetviFYm+Duir5wUTnpwcrPVyPxxBUiU7KxGxlf8RenKPZlnA6g
cHkaL23B7dYUPMFDm1OGAbHM8vyJsPkShwOAsMPQuHZL4+r0GdtKbC9MUdWyVkeF
IX0ympfYEHzXKq7CkICWBapqkOQU3f6/pi574Mq4eihf5Cad/ttP8FYjMCFBKobK
rTb54ehBwVVyTSO4uNdekDqk2wXwpTzVWitWhZz2YdhF2EELn2Kkg5HTYX6ZGguI
8KK6X3VeYC6HJyzsVRs1HH9eJsVLgF8VkGXKvw1DvQahmeWLdtOKj/TQh68eXiJL
49dWMKvfPqCUxQvL0qQQiLX/aADh4FqlghY+RWdNT/vaMkJ62IDHRioElEYUG6Xm
pbJvhEvxPm17OT4CsUbalcu0w8GHjHY6OtbA14aiEfcBO/igkeNlnsq8V8RVWVOl
0TI5T/lIbfvfikEfwmV6BNC3OBiDPt2Gg0PrzBNd7mysRCI9UbFpXrt4hgblTuu+
VI1jlFIA3z6zO9VDJ76DASXvFWdPBycmsRqxQIHLPLwh5QLyT2aTaSPryn7Xfdgz
fscU/hdxG40w0rglnNoEECFd1aFLsKuZanlGl0i/OBGgMeKbQ/6I+o5WRQT+XP8E
VYpiYotnpsiYwXFCp/X/WOkAdyCtpDkPgGkDm9gv7hzjorfHL8UQLKdC0hr5S24K
fy5PjfpUi0PE8XEkNfm+BOnfjNZBbsaBePXfap9jItyXvXsNgKNXkkMIa2iSkwmU
830pXljADhYbNwpw1vqa2TIEwTPrKSrFkwkB0U4X19AWKBEER2POq+2sbDRUOr9Y
uf8KWhjTN+ZMD+S2/BqPG2Z9vL5+83j+mjRHxBR6aK9YS0ls+xYO0C8yLgUec5zC
KTD43fEXWWvvSluh5lKfzApOlbh1RwbcTDzygM28DifOF1/ciJ0su/RNohLkayd1
xVh64NuOx1n6AghVyrdrPGzxCxrvePnC6jcMKM+3F0iH6IAjDyktJky5bzclHjeo
Shdx/O7d7+ttimpVwoxYynZzMPE0C4uKaYAC63QJbuVyP6eX9rZfEzleKKLspC//
QzstBbuIPnKXuq3Vj1t2R4PGI9ARS1lWin4ceRUgDiXDUOuPD0zH6yT4+DALQCMD
wIyzMBx7JuMSWa5Ld04nh/jaHV00yiwS+on/F5FAndaO4zWARM0beayukBnjq5NK
VjIW9uSLA2J6LkAeAmYhGDPjQwSFsKFOjynDVjGeC47/vVkPCSytqN9L2Y/wsZ4t
9DlXoZ9jm6eKEG5JqTGmkfMrjHHppaH7Ybw8M/1IZR4nYIkdYVMFq7KZsHe4dEM0
3QLNbo/1ykIoaz4oP06DA1cNGlp3QbWVMqI+rFE1oqsdDG3j2jNftyC69w0AWu5Z
PBo9V4G8GGJlIGNT6s5utT/NGFV/VPEbKzdALr5Ba9P1xp+bqWpZug4ranrju6sU
hwQ7jfDLAV5YBZwT1+lLhk3eTb3W6xS3h9dLekarA9f9fcVLxWGnOKU3WLgCzh/3
6bWXHDjlGZI4wUzFI08hcwM7qXfyW3BRr4sFKwPZMPX6sxW0QbXoIFi82cnng6Hy
xzO/EciyfsPdlrkoZuYkFXyRu0Ex4cZ55FW597BCKRPWVLzd6x8RwjDuP5BgAzUi
1IXyKQpQ9ICQj8sxA7bhGt5Ee8agajncd2kRdlcoPJWtd4FUIlaFHX3akHCfcOji
hMucdXDdvh3BFg9nM7HIdClutFGZ1j+nmgKKxgoYeQRxx9wQzRCjfoQsnoJeTNr5
iiwU6BzmMf2t9isja4LTOJRA/ph6cismtT5uHmJmt+FQtdZi6LDM/ywIKvA+M2/v
TO1xqwpHystwGoVJpQ5Z7Xi4okvGTIC3imboCax6Im8LnCuFJZJZtY0aF1yJlewh
38k0lfJim6umRuEtvBXQxtVcrvKGbJSmM2bgbAZn7uTT5l8zh5zio8IKO6nrwG95
ZYXgbrDJ7DkwnlcdgTduZ9FxIrgoNwAKFjYy73FjGhtictz2fo3koeFsKXoclspl
XkYfPmdxd6tNNH1YBv4GRPbmckssr/x5SYbixF2GuLnGil0zOR8RAAafk5XX2JPd
3svJ3HhkGWlB26CgVrzkWQMyEG4OCBZYOIXMEY12liINwDGfnSz1zR3SzdRe6HYk
YwoeS1hdpXxRtpOBx1W3TNomvNLxv37QdZiIGnsHmq5E4niw7Rjq9gKDD90TSSen
S8jDIGL2k0O1Xrto/SMVVjQrUAEikp5ylu3qSHAza3JO+hopI7ldf+56Z6X/j/oN
1wO8BfEhwxjPVTswSZV0L9EIiZzNk3KCTddyCH4oT6GK4ngiA8BFrUsh8NOYeinu
CyBViWR9Fk8InyM9ppTuzc/zqyOZJRiZS33rIW8LctQFy6yxm7064ZSoeYf0l6mL
TbJDzF+xyfMZ8JCOm2smbXl803KGtxPgp+fhNFq5K52QBrZGuaIfw8yzQWnkZiPe
7d5F0hsnqQvT12vYK2iYXmLKQCiQrikH5S62xKMb6uU14hAESA56uFT3m+semidB
iedoCmgolvwwKK3sQhhVgH7tUWllH7Zxq2rRov27tdD2h2msc3nEwn/KKZDJ/zJ1
3PEX/iYNv9ciy9GcOGgatShtKHhY7kx0QQ4n5SOSgPJuzjUIVyDUTOus0uk9bRTR
mCQciv0Zp9PbRY15SN8v7ycmllGxgvfM7GiF+EwIE9PLDQtik+dvxfn2HQLAbPDF
lsyE2uvFH61KCt2AhB7cIrMX7IwmgDOWVFhIs+r5eMm44DQrr7eN1XgNPEzeFXAn
LAFW+CW2AyXe8DTnG+aNyzGR4Ibaq12/PeKr2Ulnt2o7lUeBcQogjS2baRqX+eCg
sZpdQdWARQgWMZXKxDQA8Ll6eSwF3nGT6g1bbAh/HyvFydfoH9CrPtbhVXjdGzq4
SwqNJfJp7i+VtJKWLBKP24U2cLrjAS37Sr47wLjoL3xpz7OozeSh18tL0NXNrsJE
UVCNguWEpeFzAtq7jC0yYbOjJsDglegjUr/qNrjcbysgufXWYmz6LBLi+mifovmW
ajkoM1eAmdgGV/MHmLuDa9VIZiKf2cYsBhahgfJ7uin5wN5d3lrjwUOPXXSobSM8
lTyWns91rsRBrbLrLA76pJkuQ+4Lg8DJl14m5nzlAtTopqUlRA0G+81kOg1fyQmI
7ICxRBtCEMenLmeVFKyEYpH7uemfs7vKPWZ28ezUG1koH62Ank03MFsP7aV0YY+k
wQL7KbaFoNBt1kHrPEYVV91rKW1iFuyjX31Pv0JJ4qSvWPOniTr22rk0xVdToZwK
wts4/haDbBZIM7Ffy9jE9EBUi2nrIWwFO0Iv+5+5XuQ4Ag3j6XQf9OgB0p2GCvSj
Nm1Er3eFuKy4oVA5QtctwcFlHPZ0iZUi+4b8gLsf5B9+6oHufokYZdrbbic07IY8
1Uw/t08zDnug+NC1wrLTQXYeoCJSQ0lnz+V6CkKMCx3VPwSmKRkBVLGyeB8bEZrE
tvq6vzUeA/eN9l+6ci9Yp+TIOekZabAxF46iovQmD+Z6//MveTcAvq6Jba8OYFEp
sGnG10QulrcyBEZfu/3+hwZVmnMyQtyVDbORu3+c7bBjrJv0caZzZ8Ke1P+DtTL1
M5JrLjIKWAjlvaLltdy7YHFxeu3Ieko2gxw8C5UgmtG6nbnLaiUe6kZMGDqTYjxP
90rON1mleATGsxfszpWHbU+gIUrL5+qsgZGz7hEnJLcwDM9XpGkdyLSV9AE+jz+8
j9jseEfMN7+tJ+rpngdRM8sF3o23TW+3BTPpcZT/PG+HnYGs7UOjxC6Sj8o4YCjT
8WS92+OmMUOzztdAB/egWvWJMOhyeXCdo/65C5eZwyKDhAIEpuIqr5cahhW1npeg
9PN+qkfDFI9kob+F/KywGXazyapxhOmrtnYrT3XuyP2YV14z//fY+lwjFw1SCBcW
kgBTp0qD0T92t97AOm24tnnh4hfC4LiR8HU9iaJyqexvwoHIKelBkNSW/RR6EoWO
lMt0byHgnui2VI7pCnGH50rulEIgQGTl+wjVpLIeryHr3ukNdznTLrxM0ZMMBxpW
n5XAKGBtgxV3tNAsCueQMId1U2TkF5aiy4XNktB4BE8bE1/GsVoR1zSsw/gwh4Ra
unL1GXlN1fsrA5VQblmHXejFKvpJPjEsVNdYNkiHVNKxAYQj1tmIRUDqsKVBCnLv
B2kjt8XBZV4qLXMQ6cj/E15P6SYna+Vq4ocYe8ylJiAww6Cl9N9dpFtI+qQp497Y
SP75bYdFcZqzEo1d+gfcoGmXEwRsaEYLvkIOrtq1PrAxh+/m+bN8QlODQvDnb4il
+q+qdIHy8qDBbumtmUADXGLmYPC/YuMv3T+bvbza5zQrNu/0LcNaPbPMBzJcA9Hq
ra3Ayjk8eePxfEZIzL0sQu2k14JgyVbWZp/1kVnN/5bjq7GhE7T9XoK2xCuuFwUv
+jnTvxGs0qLXBKn7SqFuhW85OL618NgUzlCBnYjK9LufVQo4ARF1ZmlyeTttPI/8
reLFc6LtEB4UArnirhZ0MFSollnFjx7eg/KJhmS4GQ8WbfEsB50R1Ux0nGFs8ad/
+orOCKRcbum/8UlwVbVNZpBVYXQ57j7c4SGPEM9TU21k3/8N573029fR54L03vuY
gdVupTy95F9/TBwsc7/bYfwufthA15l2z2xAHzB7RcyFCQvjEnlX4MeLQzdx3jyX
2QBQ6LY0SCkF+PLOknGpSM5xRVLjaQFKgcHecMcE05Bt34mPI+1V+1CEjTOpPwWg
G57sm3m87aZKqcoGwbRsgBoSj3g2GXyGBOaR22BHZ8Y=
`protect end_protected