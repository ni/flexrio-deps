`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8224 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhBNVMbsl6PTB5/ApNH6uD+AxODPuZxQZYuFjLlj17wTl
A7UTN3AZY/Be5WwXqD4f2k0FG4yjoJUmHJYp5diUDJbaNMtYHJFEqhvU/hHd6huA
W0/1EbF2pQ2I7mITqVVzxySeUNq9jd5QFQ3t/IDWS5qElAZzc4EVk1WcDqZ8KC3w
74k4kLJwi2WO2IKnSlVldogFfaP4da53f9FGoKdtmwoweTTgDzP/cby4GigqVi1q
yjky/qnsI2vtrvAI7wflhHmfQozGn8QmCzDGDyjBKW7NAlATvsWZCWKR0wwetPsi
For6m0qCJix3WmYYD5675+K6YayBH1xe2oM1cVg8/PtwLnXQkbQTYWMc0b7keGQ3
hDGRJ3jQqK+QaBlOw4gE6ylNnS6b24X5AU1TsnD8MMACxsrLtbifq0/oov3zSpr4
PpQp75ieDveNb5IqmCI/EG6qHLABryDY3fZcvSJeTt+97VaJK16+/akQ+ug/4IyX
GAHL/YN4yIEWHSCCDcKvEoJWBQxhSAh7g03cm3BOWf38/Qo+pl7A0ZhMTiPhoWIa
x918joa5wTUpNr1NbDZQdXffFOKpquCr5qz25Mc+XF7AYCXugssH2p0IkzUVWGkO
wT71KsmgZHcU1r6iRVeQfpPUcG5MO4I1QsKpW7k3Vg3vZhifPO5mtgyWGyOh7b8E
4F2fgm8FyfStAo20KGMzd5ZQ5LYC7dZPiBSquZ/J9aD8KMiuK0OT1cjiVYkzHRah
zs8G0Ib1FpsEL9pI2S04Gw7Vm5fqXlkvUrENAkcZ5fSOiLgVWqQaSa+5wojuJ9DS
1Pt6sVpFBT6KcTk3GkCxI4Op0ZLMuwpkerq1c+i8wWlm7XAGwZjc3qbUTHzYMM2V
5QCDAPcfYtExP/tPRYPkyLJ1fFU4pjf1ZM7t5FCtWjoTdV83Hp1TlNVYDPuOxOyL
UdLqhzr3pI9bUTe5j31oRQj6DqC5po9eH0DIfqoaNiV5qC0Surkrfque1WtPjw3t
qkn7gQJa1J1AeOoK53AIK8QPJhcX4XiEchBruFR3dB/QQiEgA5U7tXL5ifQzx5jY
zJcfbmGHJR9oA7z+DGu5tP1YKYf3QrvkVEiQEVum+FvQYRWOHYAJNYQ8cL8KU+Sw
MAf01MOkkcwTVHAW60kZE7+aCREYOqnz5YpFjI6GCtxHJmjafdJiSLeB+3HEqsOA
hZQzR1hRVcGvPvdS2I4AN3Tk7E2HtL1RxUMyuIbCXJ+csHotsVe9xT3ZiMgN5Q23
LQQRtcGRvEYjkMivxDCMzUIx7fz400b303gEHp/vxjY9tAUoBPwmySRyIGuQWims
Qngt4CNUNiSxXmkBNluKBwPpRLFy0yU7TIEFfTPB7v9uLT8eEKqqUSi8A0jNsxMG
L3EtXwMAdtyVFgcnZKweONRL7wdcMRp9CgL9MNin/sUjVgzIhiOCv0AUiEGXyRZZ
iI3SRx6Q804MAGahk1IXwUZAFjQnxIG/WusgziHfHsIVrSwXwjo6uSf3ikiCYoqN
6CakD9hK9J7pqxQLcWkN5mAJEq7B7ybwmEj7N8ay5WKU0MEDEp4+JmcPpYLzodL0
RQxSWytenjI86MNLzf5aYotm8rEITA0i0bnTljAAQvEFgecZiQdkknfL+cH5MJqa
aNrfTuCu5Mouvf3aaFKSCFsrCMIm1fOuQL1blPdYdftmOID0EjVG5rmdcXRl0jG2
+gCZg5NvRfll0r6pHSPgCM7CVyXp7fYRLiPnpAvkRMrk2HnObn9P7OPpISNqKSgF
Xlzak6pkvfoGxnCLQ98zaidK6aCd+LmAmNkB/QrUyrzvyZpfHRe6vyTONCbLQAZZ
83wx/TV+cAybJIntNgZpxZ2lom2yp+Bl3x0dFfTvMY4VPiSiNnHOUexS5cU8AmUf
QBPGU9Hdze2km0Cu+m/98cRuOoU85sCS9VH6oeejoJR+on5SNqvpn1fP86e4oGlC
WpkCQMRtCFDxJbNmnShOhVfwrxsZwfmO0xThqK4F16b0JRM8dwNFbTIhwaGLV5X6
dEiohjbF+ZAEfOxyGA0Skpb4jOGVxern/+WN1JsT02VN7HxRsTOk/aPCLlIGDbbZ
kuD+otryho9fvXN6gjYYsXByBSjB/5X1qoGRFIF6kCZvAmjoTL3FoONWMW9ydm08
mb2uGb6UugJZZaHNp4L4fI36JmaYjVpf3Wd7fxNk3Cb/ga91ibBuYRPlLSH2i4Ok
MzUpAJcBi5Mb9M570VNfNeKWZ70mp5n5aoszxzFomUVhyz+hOT9KbHxYdSv4Ff3Y
159Oa9tGWEx+K5i7JEbfK5RkpfG/6STMJ9mNqMVKi50Pk0EBXMPJwIFUBHxYWG+k
AW+WSc/huRP1ZrBdpdQJby/RzxMx0m4gVZWpQ2UHL3+YunfB8xCPkxDLEDpQk2jX
8ZYa4AQhILcpaJV4z3mHg5z2IPbZAq7RKtk1nEL6j1g/avj7JeKLMOW2dm4btUPy
P8tsLT7Kj1LPNqPWWNAvXQFA+6shWdvl4bOKOQ3i2HUr55gJiiQEyyZvY2ohWXLg
XK1wuucw8S91fuG/Svts9Pf4WoMkogKYhjMFgQbbuUbzwXfQiESBz8NGfgrAkhoO
hf74QtGwQ6ES2l9eLbXZUDLWqe7ptoFaSktrxUU8ftGv4B83FdkWBPrZj024A4Kd
ZqlLKl5KqQWRYjEHWnVOBydWmaPPf119M7UvPiuOXxGLHZ7MZMQtsuZmXsRkkLH7
EtbPzamB11vfl5AV+tKoiHgXazlQCTAGeReHKEk8KVxRy9WxpuHf0AO4Ej0kAjRV
d/vQzZ7cqY0XV0SDsqV75mrGrpzrcVAnZCkAAkjTPXmm2MaWJbRxulFZxAr+gZrU
3v3BQV8m+vgbA0+JtZ/7Fo+kp9ceaTfR8eKrnuM2rK6ras803NOuIQM6JCwrCqCD
XWNfv7uQjFga8gxX7JLkeLmaCNlcoKGGZ0unajtTEOg5Z7nX1OHmPssELuGckI0a
8RSIL2k0599bOFXcXcV/TBlwz1POH1NM5qZRX8JxSHpk24gOa6405ukikEAAd1Xg
o3UPJN/qzbjgb0o5vKu8HjHHhI3Nmr52Y9+MSww2yeb2xQd0OYC8MzjCygmAyAUG
zYZxnNcr1Yf4YAJL4Wxi53Q9QaeGPnr9j+1bdUNEQH+iW2AkZw9yAYWv9ooD/qYd
XX1hSSjzpBUPQ473UFrJ95YaIIKLKmc9lmmJZPZHUzLEBLynhM8ZouSFaWUFxbdt
0fsmSTxQNTtES2b/bG41tcF6e1Z3GJsArtNYl6qrd9dGVxTYyRF1Ffp5KJuI25wm
8XPVmnl/D5t6WTLCKH2loUUhCQD8cp8/T7/svpYo92wU9gRKdRzVxkGia2WDKMiy
Srl06emPq6c1LXRSuKlkrq2I2cqBPvR6adq5BZS/LK7XkMYfpwlWx1xWhvJZofwd
/rx8FdmenkcZzUCdAnaNZVaCTQfS3C/7l4NOqU4g1+59gpyneFtrdzQl+QN0jsy/
D60IGYQod/BBqDS8ZpTpneAfaw0O7ir0A7/6BWpmj9KnHXfD+LvqOtP2fAflbH8s
KnkqTvz3TZYElFbkwCKaDI7wK/43m+RbdzYsIoym2NZ4upz8/VQxHSIT+rhODfds
7eHBD3dmAFWxyWo6FnfyUCEPZRd8559d+v9pVDVXSD+w0tP7UkkxoYzQ32H37ZXF
dwvTheDVz2r+QOgwKnMKUe4HF84oXqw0oVoQsMJ1MLhW4K45u6JCZQM/cirZDwBS
IUV1mgp+NTEVXtkRfoxWxUA4ymcR/ZeLCGZZUongJW1fLO3jdgAQzzVN+0ccDUyW
W33SB2mJKqRDfF6Psd2ygC2toO1i620G30IddiqhCkE3O3OAg9gMZGW7koWp6/z+
01YpM1X9/zYVBI8lzoDBHzqyzP6YYHTBRkfHNu7IF2WaDf2eqvjWOyxNZl0/DKbp
eJ/rQLHJuS5WYM7EREhCeNNZmBno3IFy6JA17MzIA1S8edNDHoTFj+KRW1UwJec7
NIPHRglfHJcMNk2o+vZiGL7zsLdzPcOjwlHOBYUEtobTPFDOQbo7FOAFsRhsoWqj
M4KJOkpSrjsUiihHkJ2Q/89hIzmohzyGhH12ilLyDJ4Zu2JbMXvb2HY78znqGuxk
dWnTQSPkekp3AFwWcVHYcQ3fecep+ZZu1IaFmDFw0coJEicQjA0vsZpHVpTRu3/o
yDvn1afqdq0fBDjmwDZohb0RR96TCtqaarnbCqQ6xTQi4z/UmqqfBWn31ySUCPug
qEn5XOERalfgXtJNg8ZOuGWYK2+sbR2PEYwE/9fufYIBe1xfEraO9ImKKbnDdsRe
vQGsT75zcz6NcQFDmkO+NADe4pb171r1Tn2c7if+Z9VRAheNm+DBxB0F39gBlbF/
AjziZEYMBYVuijhIPtXgqKxPd0Q3g/MCZhkONfQg6OR1rIQ+/ugfUdGS6z4duDc8
bNj8N8zSTRwfEbHdDVMhM0Zm4gYR9gYU+pKA59T7d+QpsGXUDSNcaIKOlrxsAYeN
VxfUnVoKsdBiQwGfqhV8z45BqqmjbByHuw1Yfx1vIFia84LfLApY39pZ91KfZ3HB
SmCTYa05cXpoL9e8zM95hPT/H2yDPmZ8EqglFLgu+UXlNrAn5y3xScx2rYZo2LQ3
wH5ARsmzGvsxCZFjQaVR3OTDjyLxh4Ggh3olXLteYm+x7jSBmeRD1csCQCeQGFUl
rzX3hXiAZqr7HAGXIXiCS2mPoYRuvcni7OTaJ8Mr8h5E62AjQrbqdqSoioVFDOOv
B83Rfm77XEOKYBGQof4+qggn/aJF4k7QoFJw2LhEyFCu8y4UmE61uW9NElBggWcA
vhwj7W6PyWud/sK7pURLVJtFFzaQTYwwXhTeToTjV1zlOcJYzzG83+N67JS1N/WY
59J2iS/wUcMB1s3o3yv9sT4H9hLG6QVeX+ggSyVgNT/RKlNGKVfL9FEmUH77RT+K
jIZoRCc1Rzc3XI+N+UECzBvmnteBageN7bjBq/1knJcz04312PxjXECLONST5F3E
I/G8HND/t16Gyv8jWDDlmaiK5EbZPYermCKo7i3Dawifz6KrocG9mNpZgHuRVJZ/
5iS1WCG2mxc+UQqZeubnxzmgKu2T/p6Si2gB01zfaCD72O81vYOQ4i/Go1CT3236
dpsMOAXP1wPwHkU2OvVOkpTIQlG92uqmLyCya7UlVrtEcmrJgDetE8vePNU0XHbf
0L0hQE3WfPi0QxW8KnlX7k/Uc1Lc5AurwwANvXfrywM4rmHXD5PRoaBH/1mALbMs
pG9Wx3LZeI/cbQtJs6yRYQh13zGAWhUi2IROB8ADCicWnS+13+qv0Sn0IXx3RiPe
NZu9IXAUBQlP9AlBFEF5MXSv6IzZ5KJQij14tVbe9mmmKcyuRVO3pIGClqWdybsq
tZmPsPC2PKQW/u5hnCKfTR+sBFhb4wkierTi6qOpvQvjjpv1SmoDzMG0WCkJbXiv
ADnlIMP8hmE+jGyuT8QcCaKdqV9KUrvpqb6uSBcTsiPFdTH+N9AM5UCD3ED/diUn
o1fTqd1RECcmvbur5eCXvU+kkvTj21sNC6cwuhGu2HRzZoWEZszROZSIVVdRlkhO
gN400Nd0iiLMITWVuwwasK05cWmQFDwJWN5nOeYMaAeSdcL8uQbNGTNgMeXp9N6l
pumk0wuGSDxvb5FNMrHhrwrqkw1A2ivEfzUJz6aXSDln5aKhc2cKBDok7sj/PTVf
TTeDKNfnZfhxNnLH6XoH1vUP/8Fkp/uR/VEkvTZsDLPYcKyFaVnfT8KIsQEz2jv7
xzCU8hMkkAzrNq10Icp+KOzex8Ek4l/MlcEYLa27yTslqdUsCQgMp95kJ2wyJ85b
3KXWW6trt2hecCR2ShOccu7A77toj+Bk3+3tf6gWOMRz33NC5kCbZrM4tUE6FImc
bplUloVvS+ojcFjpg4H50N8Aj4MYHT08ycGD3SSLeC9aeDeHDxclNJISsJ5Yzyzo
EBCDI/sFRNiutz/41BKUpbzvATdYuU3OXZYqC52KTywKHUXiBG+mGNuJsiUQDjCZ
VS7NDv6VF9hryOARzqrYtLPyi5cw7DATCJa6t9Pt+PEaIfKrzqOFHn93y08ZNqTo
+dIBKzACB7lC4Nk+Aur2109HO/xex7YpUdHdtJbgGq3awk2dyuz54/sqN9ZFoxmO
bEadlo04DwhoUJ3fqyz0FB6mkgG2pf9VgXUbZ7ZjCLiNf2pjx/JUaDt5wUm/sM9M
D89QrmlDbPaWReCcChm4W7ufP4thQO7cgDEtrOyMLwRghovsoeSyHuB/G/7mEiOS
e42SkUT+pip4wX1Ht7UwJIU1F5rW/nBRGX5rslp3a66yW7mDm/E3tzfsDFxLGwLV
1oKgAyzzpbXIp52Ng2OGMuPHzkDssNQScKHItPaSklnPFix0TrjSJw+oq3t19Li4
wCF/ZBEEkRHXe53Yjpz9NDq4qteBlNRRlzijyIoVXqs5UhA2TvcYrJdJ/9T4S7Gy
lnCYIC/x3TYIH7F9sXTSyNvoC6If3GWLPzDk8NwSP+htZIjhgokCQrYacSJ4NOHJ
/yAdxi6NNRpxNj8NfFtuP8+sW9Xh2u/wDqlHDMnltpTArZf9uoidCznF1+0kpwLp
ALh3wnDwgTZzkoFOIxYDYxu0ol1bNlZSFXWB6vVKu0jPaGxYkUZFMIcqPT7X9v2x
GbOfiXg7J2waD/Jco7J0KRXaWttbm59Pxamuu7H9ppsgg3f1yWWVaC9HDtTM9FU4
quZFtQorEpgYIyahtFOoRm5wJyXTG2G6+PdM7GYBy4ztWDvOcMxmp3ewmiuMiEIn
PyiKkYWvpEXxUEssRQ1Iin4ytAEm1upLrEM7ccbOC3iY76fSubrnNPb/I+iHubDo
D/PRu0zRDHVU4+SYb9VPIKrGr6+ZoL83VZZ4b2XJG6sNBRgLwe/+zGaI4PqXDbuD
zHbRfS8VjkcaN72rjh4PGiXSo80i/nqrgki8hKUITU7UPuPs1CbTzzUCuW0wqnmU
09hoYYZh95V9M9Mk8mcrH9y6TpKzT5gCry5J/5xQmFSLFZ1NwPtPPxnPl6/gyKcE
RBJEM1Yno4Ot+n740CuWQJ+M1NZCRHPysSfVeWqSbdTfw522Myvbvs0ulkqRsYmw
c/kSQLcuXBHYQpX1kOoaSD+BQF3KkFYePqVnRWftCYR4PYYL8vftp7esUCBcEbmH
95q34ZSuuoM9BVQ0nVFfc0D1OeWIua9zBQhvp8ZCtGu6K/erUGDQw4zcp//trTzl
uRqvhWKnKfCpKQ6Q7tkPla3AKYzEJNebee7PJX6kg1sxI/kxkycNMCSTzyyVgN2Q
IE211kwhj/x+tzIYzBz8OJTkqjx03i2WPITXQV/9U0jD2neBiirTcB49tVE8xkFZ
doVgtApGElts/gMQaOwrhvuCzTDmR2uYUj3kPH0PcXNBm7ZhT1F8OIACVTTOz4sF
kIet2x7LbUGbufeeopJvqAkFqDD1YqmgcmAtve4hU5S0uhl9fTJzEPB/pEj8G34f
9nA2hhFN2birK+2k8qc63e96y1gduAMq4s55gU8SQvxUT5e2qJ30Op2JE2do5VZo
yITpw8zb60FBo/uTFLaMvdL3JVPhfjBUkV1hW60Z8Co0ctw6bfvDL1T9cUF54xBF
Ybt4cgROiRamp002Jg5VGtsec2oCT8QUy896UkoPlHNYRJWTA3o3CQqtXTp8nGvv
nKdc4lO0a1w5ILz93H73X9gn8Na5tkZpfJ47ecZsG8X+hk3ZrEn/60hSaOYpIQux
tvcs9cNK7HuBLiRCmv0mWikaq6pJcswKD9wG8sEa5sa2fTwYZKEoYOAM5mwdZytA
/oZ5FIBu9gZW7Rvam4BYi+MUjSipfN68ejakWS1oLU0YHtXTSL/PW2Ls7dlQtrb1
qvRlklwDZkERI0V8Z6ILFKzeyWqLBFKV78hhx7ic2j7zcQTS4X6cy/id45xLSnn7
Gse8pqL7xxvXUk04L+FMj0LK2GSYytQ78Fp5iofEmUoUqZoD+rEaQe/mdW0e1i62
CpGdf46sP4dBHZwaeSGFXJLg/4kfh7yz3Qg2bP/eaI/aqKXSrrEm+bmzxFvheF/0
hJW31OfO0hNY1ay35ZmSEC5jZoEMU6RbR0aBfMF1VHYK+IJmMTud8epoEBDjQXkI
k+dE1FTTr47VhP6wpXDLqvmJuF7XVEYt9jXid9QKkp3w3VvxbwfzP2O40KmvCz/p
siBm9LweDpu+5T0NnDvjFAEqTFxxCoJ0LeyQajzkRFJfn6X9gMZ0EoI39xLbWjby
H9tuYsUwN3WosUZOp34Zq5+u9zVbPu0BqT+Wy6smGdgLRPS+BtE2crFrmbai05j7
y1HUo8mcfaMY5K7sFADzmiORLRnp+FfB0XCo7zfL772IKh1glUxgdGYmF19PidHc
h/GxemT8z1wUDjmi4wOMwnG3WMT72HiZZPYaqCKbNZGeb1EZ3vdlSafTlOv0mw0z
ReuWb2ZHwJQ5wu3LLHx/sEldD5eF5HsxqGF2iFgRdIaUfM7BOoyQj2JQrdHTuWTB
/ckjxsRzqWLNRfjX/3pTjAf+y1cIDFN8THLeRgl90taG96blntGhXRuc2h3h6NvA
efHc6qNPNRRMXjXsRGV3r8aEjSxzUI+dpcdJ+rsX0uplgDJkwsolI2J9ENN4uh5r
cUMgAyDLlh2tnzgpIR18uKcW0eh/PLL5jsqr4H+2AOBvtRj4uB4B6CzLTnwvGwYY
lfjyaMKo7K6myg7AvO/qiAxDLZdhHln1bRw00SbSEBQ4PKZz8hEGpy+mJaMhPYW1
35K2Q1rnZOeh5+9JMOqjR+z/o0BaXV/tMTuZIV0NnIjgEa8YQrQcwLTaxdcptxxn
+8I/oMJ0Y+3MPqBJgjQiXVf+CozQacYUcCCb8Xhd2lcszN2bctW5q5ye8tV4b/Zb
+LGvs5qq6KznHAUWuJIII82KtjAoEXBGRO01SiOz/P2XJ0woGAltrJDREEYTU2dV
eKCYgkdE8sXeE9sguwQaGQb5f45LVQudc8Kyi3wMmjZTb2GKazIVxW0KT6NSGzWf
i94LCZLJ8xZDAkLK72YrT63QPe29OMZ43WTNfzzhC29V1w4S+LoAYn7VtSOH/fDp
IJJZN2mXY1qGs1YedrSETk/1W0aUsETCrGZH2b20ip8zAwOiAFfsmNu3oZ/FauU2
NRWil6/Roz8QtbzvajZ8cIqlEwSZW+N1mgP70YoAehDLZGCY1RHiytg5HYe3qFHV
YYxwq4wnnWJkzm8k04EzOGaZKhnlUWrm00Wa8WGk6/aL5KSynKbTVTa9Vkfqwcxa
xPK59ZhFPtzhQnSeCw8h+2sYNMgfdPv8LAlLQBwfDKYp1n97S6QB5VxOmIRf+RFc
yb4cV58m3L38lkwsEoJPqA8shUOerL6Hcov4DyxjVXbpXksmOHAo1bGqSr8x8Za9
F+fQ+1/E1r/mdNd00s72kpUV+tz+pC8rSJ/lzi+XKSbjZXskpzWHPFjDjEWemyNx
wlEfAGbhEoOEZCSp87dvhTgnnbQq+cHlrq2iMa1iYrwBQEqGA4N8ikT3Cu4Mb1gG
lth0Yx/b9T90LlhMtUKIdVh5ou2XwWKoqvHyreZDD8g/dkvPbGU1d7EmRiWu/28l
cZHWhOTlTAb8Z1vPW+q5ojDsfnpZL/9IgYFh6f5WnZP34cN6CqIkQBfe9hRlitU5
f13MENqpVRJbRFLR6Qz5TEodrDk18d51mnw6x3LIUAaOXlU8LbxuaRVkBhZlDD/0
aO8itMvdDBWwMuhchEQlu9bmT2D+RX0/w3073yz1jZ31UQWVmYED4UY6qMDktbVV
ftPXPN59hynj2ypgmuxIyRD7yBrXvWotqhs3vmF+jU+HtI9vunw6bBoqyiL//KBS
gPHxrkNseNMQZ/tmdC+0DowXMG72WNZ9gsIhM3hXDmyjjgHR43Wo1COU5aU3vMCx
wS+4VIKaEE2i4JA5/WmoGaoz8ZWWl6Ttw6lm7CPSqsKIaz1uEN6eqSZ94ALeWHzP
EaYcZ4IWmREZPWoMIR3u2VbD3wSA6idmUoueEuKtnusi+ed5Du4qh1TQPsSYO2pC
pi+Rts6biE7E8nabpNnsGg+WtC1asdL67+cqKXsynBym53M8sADdG5LbuwnozpNN
XOp/KDUdEDPHzZipUaTdQXaUOe3CBjzHlp75HCVcDeeJ0mKQHI6rNblDvEMfzdyH
WWacBdfLuJxpmEfEhhajf+yVr/V55XzxusexWrNmgPPxoMFhkHb0Sgqn6v3/63WP
chvOcKHcQxcS+Ri3A5cYzrn1lyntcfYAeSyJWFOWO+7J/5+zpNJabgxVB/C3PnXm
+B4txEYevMQs06dSqFUgEQ09qYeIRMbSnGcAP0+dh2QKwq9imNo9Ts95hGFzBAyk
CNwyQfx9hUT4OuRB54kCbuXNZBNijMCwc+wqck549vebxhPpGwOIbW05hFvEvV26
Mmsg5mdDF7gF328TW+zuAPl1L4Ms/bguonHXVXEEzyZ8jT4FcpNcrJHyujgmOJLh
sX7vBGzbkkNf/9sYbq9I+j2WFKHgH6EMQMZP3khld36utpO2OU0ZfQRqIZAK/LnR
YE19GWoiMIKTfBgfrY4KerAvnMdM7XsBz5mTwQpzQ7/fb4fW2iFE0sTbsYPeYeFa
KB20r/ZV/2jfG9DdPLOdWp5nB5Nn4KjJlbkUgKEOK7G1EWFeCUBgAFwe5lF+W27t
fkzxFeOgg/KwN3SsaCTU8KntoVjYyeEm4Gwb3wiNEEhSEJRNPPUiJKOmUyC5a6sP
JBVW/E1yAalciXNyH1Zdcw==
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8224 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl7TOuMe4xzV7rdHsSWg325uRR93lr5lVbjRD50FEwmxi
VLE6DDpzj77rGHZA6wj6bSxvKcxuCXXYiss0e/kuGtdali3KHh/gZ+/KUAtg2aXx
ajNlx56XA5JyyTMVsg0a0+Pf/nYbEhGq/iA8TBSOeDYiuiL6W3KPMBTajvydPqWx
JMfHiZkf6/cf2KGGlZ2GE9sMgZSx+UXg7ZZomjQiEklWNPn+ZG8M4L44z4lL9A2V
72aWu549SFWAdA7kp6cmwRDHR/lwD+MC7K31v2eZBisXZh1mB2i0FjsDdI9s1xfr
FGwRxRt8pq7IP6Ei83Lij2RmFPkXHBNXMVDtiLdo11JIgqlv/6IUI47J3biHJlkc
8T+hXBc55L9efeJbQhSIGedUSygfHRjzyRECgQG18gh2hCybqDfC3uN4illxcvuw
Cju0R0184cm6lCoTtF+wMrSxiE+8nwmpDsf3/3U38gD8JUHjb8v7mzeHD2bDeZas
1avePlNwpo/TFlzW+HRU3N0UxJcaivryCfaI7ITnF/Fm+9D9tvZ6JKG0YH4VD346
Lg8wQsCt6F0KieM3HXF1InDLEpqKfFyc2o1fD1UrXIfde+Iy/zxhchOrZC2DkwJi
6kD4NvWUy286q7mpqUp1Wt8oG6qE+7AkoPqNPnwaKHF30uyPWFT8uCWr9LqcISwM
oQMl6AuC3cm6DWcLg2xpmyLA2rgtIcNocME57jcGVMcIWgJMw+xb/HxxTf9fzep3
Bgilr4rQZn4R+Ciz3PZgBFCjhOhfDPdabvJK/vaLng4z/OCaS7lWjfAl2bGT3Ajr
7ZXCqzAjysjSGK2Ni6kW0WelUlbj+ZCS14K1C6IbErhydzuOn9sRi+TaSi7/tkcP
fETpjrzujU0fVcgj3IVeKcsxK3jXUNj6S0ADo/JWZ34dkf2wOuln/jK4qKxtmaim
M6Mf7C8f3gGGuauTPeXlLBreB/lAqGxPVxj4gsnj5TVP0KOItd4eQbpXc2amABkK
K0U+6vI/89AP/SX9cjTWRZ/AlJ8Bd8BXQO88TD0Fan4HywIlnxD7CNbyBMIfyL7f
OZP45XgQP2E5OClQ+RxkrLSuGfpfds9njW3DHz+rGNkhfv04chszcfMgz6vialKQ
dsKFi1d3WB+SDQg9Eerw/ATeXy4KaI5SHNSRvcMQ3rak6LhcFKbuI1ubgU2bQt/G
fKgRZae6uqhr9B+tQRg95sryLTSIskrO2XuedsCCd7r92ydtrTuGs2gavReM9p9Z
EyAs176x1Rf1HV4UOsja33sglTjYCUIVObxjUO4ge4eiUe6yyJ3DBM1zeWkGStyq
StT66etGeusrcdM8xGeWqSx550HoukTXbGTF7EHuMGuIALqE/PYu/SfcZoaVceKk
Njm3lgNmvibJVPTWjfgWWOMOE6unuNi/uRpOIlkVklPg7uenjdSam4d82QLoT+gC
3DFCAf5aTOnkKDzLvKUFHagx+ErXW9w7dblTKWvPla3TaLYMkcV4x2Jlb1ri9pNU
YsdVuPnqUg//KQDE99G+V0axDcj9baSWDijz4Hsjne+gsdsnchGASPvGgEBu8Im6
ts66Sb53YWiAr5f3DqQi66g0iCFsoXvVqgEulZqTp7plna75fWTthQ/d3Alo21ne
ES20+x7MvEcow4ESS+ItUXot/zUXGHtSGlAJvYXyyjOKi/6DsceGc9HZVHiEFtiA
CdudLGHzf4H9jnoPcrKORz8looboVlxSY9KFaxOEUXsvuUXRexKo08TMgglonyww
fG5sER4BxNUUzXBxi8vKGtR5bJ3H9rsNiidRdA2BMe4xlOTjvxTjl5d80e/n2w5P
KhrmthtJLjuFEruUrEZAFzDWaAwxKRQFPHnLUxd82rNPel1/dRi3QqCzTw8jdx0g
vVzUhnNIckebJeoEz6NIonxSXYX9L+qQCqF22rg2YtH0MOejn5n8QnEUyb2NrY06
ybJURF00jks3yq7OV31uqcbiRCtCPKGraDPjMzWTbQ3Dd0ha2ZbVZpWAeEUBrN3a
LXiPewgJQiMYGj3AY38Sq396YYQY/DTs42uvekYmG3p5yvFD/oEGY1+pENLlspBR
JP8XGiX8GZwVOHSuQTFPeZdj8llpM+EbUDmMGaURHCYvSntqlCNFzpRz2lHFebeX
Be08bn/N9MG1iSkj6qhmBtLrQX7n/peIP+W4fnj0/7h5M6P4bHC9Ug9E6eYPuhZ+
o/c2vGbyJ0CwTxFGXuHfI/aXUxMNC+bx3vkr3fk9sWfi/4tkr9FfhbKfi16jrMDG
9eCLK8HNzuVbL/uJhuilUormoKOmAmPQB0pWRhdS23WVQQB2PiD3cel49+ozmu8r
5Z4/rSxHZF7nqAEqqZDEliB+YqXh7IZbIu12O+B9Pmzu4U1wnT7MiOX2Au7YJzhr
ifd74rAE8XS4nemo/2AEaeSgO6sP+/k3AS/Rwa3+RYGhXsl3p8CdcXcihqwxH9lr
ehHfiSMA9sgC04J00uJfDwLUSTlBHdefg452pwzm8og+UDxybSvM81HInxBc0Sqf
3YHHU8xy0pztDrvdZyljlRcBbEIIvYYiGF4u0JhCJKCvspxg6QGc9vy5Au5413Ts
UmJ9P9E4k/7O1sWMHkOaACQWJrkL7yG59u+Du0+81mtEj5K5y+eEvkNvlNN5q8YC
KzaaahFidvCGOK1lflWqY6fIiLhVgP6IlGwuF3keFpenvlW+RY46EM1TNDrS4vxK
KJj5cam39h+5d1ul/DByX0S1+4gIrJn/r0lq0t7SRUe+bVbT5hzobrqMhiJNxM0b
qOIXDnuZYes6XfTplAIQlE04EeqMnDoeuDJZZUnLayt2ltJFghj9aM9ry6jaIG+o
LgF+jUfi70uWGa93ELBpAG1Yni49ZQqtLAxQa98QykMRTjwjHy+nyfNlGVfuGWrA
xhBuTcy5Fr8hWrrI3gXm2kzx7kixhtfAXh+Gd5gDdJYWuKKotX2+Vg6OLaiSXjaE
2wlGlQkRmNxQy9H8QYm3KB+yfrEgRG7kzcdZz/qBOGhDPkBsy//2lMUI1WIkh2kG
SldWZZfxtRuocsa1BODeOBd04iM+uc3sesHxNfl4vg0tyB9uWTj4nw8clTZo9g6G
W8W1Gc2HjC+UyRr+zH/aJo87/bsjxnYvubbV/dRvvwMZRAI1t5jv7/ZWlzqUgGnR
0z5dJ5rg2PiguJEQ+X4/maPB+flg7sMwkRPzVyOxkD+KvP1TbmUrJK5TVICrYNOp
97bnoRBMp26W7JfCxledGFsvNPclDTEhN316ln3N/VPcFqqBchPARFMVkbIwZOus
NifRzEal7Mkk60FEvV2TmLVK+5G87q27DnMeCv0RXAjLcZkcCHWOsX8hwJ2ZzrZp
1jXASqmMIACmT0jN0g9azGfMSIX3ZNzciVG3dn22hhbteZ7vMplvUclJZ9bWWYms
RfksDGaX/8jNZ4FPHgi6ysOv05M4UsoRslSu1AYiP+m1iUsE0Eoir7NX8ActvjL9
QgrLuT/7cfTXUaNjgJLVE8JIfyAGaV9oHpKlCLfR4kZe/dGDJYGBSrduoebXedh/
wO9/MjWPAXDHVTLGFEOQ25jSOW2G6DAQXo9xOzIzhcrBCgN4rFJtoxjaZja77aUn
mJiHhYz3OcLYiZj+XTKnFRINPTi7aha/s//C0sFac+FNUusIdSLIa+qOlzH2w+p8
Sh56UlisJr9LSS3og8A7ELLY+hZhGGZLBLpbtu0G8D508850KuFe0BaZOuz0ptuL
Y76Mb3vZzn23nVy2mgRE7dKydmQYPDt05rOjGSgfN6cGn7v/qRZf3rN6TForBhN1
+F/5TquIXs+rNLuggUCWHjb7Ulj7fDWVGtDz5lNXegKrkO+KFYLXP4e9otABYnkc
GMK3+FIm7XDKcQrNH+78zLgLD3Uog+LpRcHLymYNgmly6kNZozb/gnnZgBswOSnl
G4i5WiYAWv/7F36Cv2lm9nzcXfWJvwOoqwxejK6dVkZggLJzLGhFsM2CHta0oGwU
ojTm+glpi3XRW3hW3J1BKbYFRgudk6FaXJyn2LilsBzPHdmw965ildyZU32/bwT+
/PKEM2LP696Yic3sRPmKYu+LE/aIHu0eNyr3PV0sQ6juZLxd2N5vmY82lWHx6W0+
UhT3QhEelL4cw3qLUml2iBr/Z1PYDLGbqq6jJbF80NTfjIj2XoYqwnCLn5O3lqxM
1dD+EHbv1djqF+HpmUAJzhiqa0312fcJVVnvNNLF2XDpTcH7SMsyeTo0jaiR5qo6
TsrrTj4O6iBnfA+EcMHORuzER7KaeXYgqYtEWkyCgZDxN4Aai8nH3seSoeLnZLC3
m2+Wb4HnLTuhUSGw+K1sIMYrGWDw35P/hrHTmdFNhLrGK303uERV+FUQc/ZG21F0
nWWVJPtDzK/LTkUH3Rkb8J4igDmeNvwDromlVKCSH2DfxZsyDYGgFPkcW79dmhoI
Asri2berfOF16CNtJZeRHB1bPzfRF6+N9tSvBy8LBRuYd7lDJKw8kdwCYXgZKdiF
FDBqXiTHV4xjghsD95z+7wAu12AKycjn5ssRX/HPuYHdY67RKUI8d++smz+M2zm3
1S8z4ocn+Z3Ouohz3wkwNLPoPiUp1Shws0veNuj+SEV2ByM6zDPGJ7AXQxAOgNwJ
ssh5iEqFwSkxHljedfk8LYBPtHzvQIYAIlnbLAB9q/Tvjf9i4SGG2FVpVjZY4G7p
PDDfLSTigBs25RTxoYmW0WtK7LNjxbRYV7L7XSqDY03MgOR5idekb0KAv+dvMVPz
c5pJ5l/TBQaVJ/kKyZeNTL7jQ3Go0hwe38H5AUWMDXbkwUcx3isb7KGvL+VGUul1
f3qs5uJLaYh8oz8qX25Wcw7MG4X78AyMSKSUivunI6SeemVWCHXE1TLJvAPprveL
YVTNsXZ4YeFtxcOdMuwCguzicsWa1f1qECHmzFCb2zguISKrN/bxaOwzK9LofN+w
c/L2MkIOTyUStT7lsQdBqxpOeLeiOHUWpIIsmxD1kAUxWDVSe+gQYwWXRFkHkw9y
YiQaMjFJErxX3DRCOoZ8EYj4uk28IOSDL8lDoqx8Mm1JZ0Nd6XKbTeITNiTSGJq+
wFS4CL8FPrB8Me8OBLP8+aeHk4DTofhvP6wO+4qai0O+VDPuYPoYD1REwoGAufaY
06INzk0bxpFxv5U3mR0FgLzHXVmR0/H/qOAd/SH7Fu1RzKT8aWwm9Xnsv8jH48Q0
UbxkwH+tTa9PToDj2d/qSMQKdlq9C+MOLvuCHgW8NSPISRQyCxKcXQlSXcwtxNNy
+g4dtNr9V5S7Ca4miMjo2NtwMSzc68EggjKdE/YPv86rIHas81cxl0ZEbzREP+rF
54MNdKFCx8BJ9OtBWyerH+Sntfxa+7NCTXbVbHZHmKkdjV2JdCWkAGOmEtx2GGzF
EEMvdAHCWV0desS8Y4BxSMufH+IJvw8mVZLxHOVIxmDXIQtngJVbPriTUWyRMdxQ
0KhKotI2eaFFl2++/R/z2UopHJT0Aq7cswtvGqEoxz829Qckhd+Um66eM5G3fgKm
IfJMy8Ogi/Zat0WZAR8EKAlKdRp9oGIxPWMqrbjpEu96q433rRZMm0wNV35Iou9e
yW904QwK/3J5h5vdWJUy9+j5d4oLxUHv+FEMJUgH9LGPu7S/IZpXo4/fa21FVZ0b
ZaxydpB84gwK6CNy/okNduwiQvdt23JZzoYcoPd8A9QglMRSRsIgO/9JufFaRl5O
wm4idtYgCg+Jog3SVoHGW3nCcsNEPtmRKH2ZCp7Sn1COXn8MCXfqPtJLMU1Gm7bb
XcdPhITd7F07MMM+ANb7TQSzOmEeMKyC1his7PK9anPfOXZQEkhyovYMqX1neITQ
8OnsomMmSxOf3TCVxyEuf8mwRJxRnauKP86QAb/BuvQF6HNTBNWaOV6Rek+crNJG
I2dni4hrQnnz+A8Cd+R1g0Ev50Ab/HltDQdNkVYK33ExFSmRn0MCpLFQcURBh9DN
xW205oZQJJV/S1qLV/1t5HzkYrOUeWrDv2tp9vALzLixq4Vwvz8jKvAChLoew30D
g8lZ8zyg96wNXMSZR+IkDGg8+wdPgDgz5cdxtKnlNeAIzdwwUTNH1+e4NOP0vtcS
BI1G+VXIY8VRCFxAbzQM4vXIzK+oS/GF5LcH1jTr5pthFe1E46bu4zY518Ex6UkB
/cZIzb2hrfiEVf7auTU9QpXkp3UrPjq98GKgjOJteeuznvDKfGGu79k1aK+NrqtA
XyIuVkngTiCtfxBIBdoRlAYEn5CcskztjjUA8/QCMW+ZAvbxVLJg1Q4gXNgQPAAC
fLHceD5/KtADMh+fio/AFgswUniNcvvTd7j7a02y83VeMNoEPGOzyQscOLgCgKgj
BzG7n04UQHh4wJO769FtlPO4s+i7dl8SMC1+yCgm+/Nz14j5Qgi5TqsBotuOhlz/
eGWApd1ETf64+jBJKi70og0Nz6hFCCN9zpmYyDxmY6fYSgGB10WIr7r5GzU6wYcG
jrLSJfIjgY+JLr8pC4LKTFjssYiKDHg4FQZoWN0CfOe8ybzUlaPgJNpgjpTgBmsD
G6x9C2Qq65aZG158s8mMFKgn5aBY0ZCSdVgYAmBklOevg1r1rCx4BPeQ38slFtci
1q9Ag0l9FtpeNvOixJYVkpU3fLA1EuMh5q3gaByM+Rh9YL3K6S409yEMxvLXnjdJ
vcVj9O+5Oxd7LRpi3cp+gZVJqVHGEltbnCrsRem6oNdM4mol6ewaeWZWJimoWeXK
9tdrrjfsm03ZAaqVIdTwRVG4GlV8VIr7w98ZabrqRLA+xAoEESwpUWzFAJpIsNU5
1jSIl95ZGwCNGsqPjhyFS/sa4pqcOwGng87eoFOZCcsjg2sCf+q9XnqFtXAGzz7T
iAAhp+junK3u6/30yXzldwmHDMwIwY89AKFAi3UVT5JTzgLeHCPh99UtYLzzhVvt
sFf/aQfeZxuVxo+zqV28j+EK9B6wFgxYzPkJ5tBCxcxkvjImuTAtvlFRq9P7+Bk4
y1opXq9EF5XfeSHyisgaIBgKdQ9LivY9LB8eWJ12nVMj0CezPCAgIuZPvDbEfz57
fLLM96DvXhOxdowc0jeXsJ5SEYk4HSy0ZvODeF6qUN21bTxzK3ep/sBjKM+0up3Q
QtDqm7MGDcgGBi+n4XJCnsJaMIQZ6RCO24UqxkfvazwXYlAGgZAXqSzqlUMwiOed
6GNqvJeWJMK9Ou8YEzamq6yqJ03jL8zCRMbju34m2kJLUHa+GoNAxtwBi8QMKfRs
vv+JYHrroCxmEXqdO//gd4xpghkC6TDDy5XLe8XJpy9wvnvzGYxZvdurze8580LX
urGWernqeZfKI/CDdePw1Ng++waZD792t6ge3eUYnnxJgIvC8CL2epH7f9vU3jdr
O1Vxr+7wv5ieSQNN1X/mclmTf+XnRFkkCdgjRsEAiAyDGBbYX2qluM8UwgZ/xoST
iDBWNciRW4Jw1Zl5uRmY7XLsKtvdQ/FZLR1d8cEny8eViM7bC+7mRq5NXkbv2bSu
YxYcIKSJ0L9e0m4OvW3hFDDXEPsdJ4+uJ8SOgiDDad5f9OD2XmmxmulK5/rTcZGa
CgVmGKXAWSZA76wgbxwqWPPRs5werQqqtfBtTB4BZJJXpg8DGRg6pq0DYS2CJA15
EiqiEuI0E1YBOkBRUkMVLTYRng3kF1QUeJqsShCwPcxFUvk7ZEsLn8WVbcxlVRfU
6wCoL4iiZOwT8e1b2lYjrQSHGXIRUih09+4Vwglz3jf2cKjEEE7pJYhebDrvyXry
hWULEzVMq/Zg8ZrQxsu9dekHYGq/4AWm36Jl75ToS+IJhhT9cdi0lrwESDsdar0x
bLGlkuIWP3iTGZo7++atPAKZl94mFS2uwkuUFPDbu+0E9T5F/5QCz5OueeQhy8OF
Kdqaj9UrajDvV7gUilL6SyAkejrsZIAS7h/U+Mb7qp7uCCUDt0SJ7r1FDVpCKxpr
VsLTXe0wYJtd3nO+xgorqi2ukWBP9YVsbSTrBkXKQSbO2ztadCQkT1RQ1ypX1+me
K/GJBQm7FuyjLhM5RWfPdq1XkaDX/bgDx7R/i6XOkDwZuS2Ye8cdWwSw24oNtpqc
L9KLQ1LCWKrG9RVjUKOweFAJgpfTbMW76PbDRhAo2G37TSt3HY5sIG3rqbRtVrzZ
b3Pu5i5Z39YFJzs8zjR9j7CzwDqZ2/YIAP+i/M9jahM7mHDOMGotPCHDLSa1DrkT
IygFTVQpHGsyWTujbS4vnf0pfhk224kLS5pjSC3V+CtedzKq9oR1JE6DrXi97YTM
YH1joCt7FlYmLmRuueF+IUwN7XyXdw/NxdGuauuOSl5PzZ0qpdN6ZU7Etv9aU+Bo
U78dMJtpBhYmTLbfZbeOwaOtYHB0uyna/PDAprrajG90Jx3VULU5xuW/t09MFhRk
UvPRmIvWeRsg3/pMR3+MNv2ceivToaovDjPlKEw434GggmZ8OQJyzXTHFQdiz1+O
4Zvq4X02+f1xwYMDEVDnQLmhjuaA2DNUAZ7b5gbfTFDJqxs+AhgVpGpyVw6GkHm8
gLMxqCsc2x1raQKXAZ6PaN2cBB/VNqC6J+VFFcxZReRuQwmq7F2Z7x7H88uRjoQ+
aWQCMX8nJ/Zh6f/Qe7ZTKEmgBBsMLjap6w/WeQXZF1wDHb3fIDRdg7dMbhntqa1h
jQxKlqG8td0kg8PehwhJODzOUU865eSFylE0HFq0W+roeh4cwJUP8j0c+gHrcYGB
GNL9Gu+3WCC5KbWSlTi3gV22GpgXV+8E6wOc/HkDP79GykFH8cKUdwkMg2w12jxf
51Dn/1bK/FJ9XDlBf231rk8DQYKhHY9TbipZ+tWiy8Hd5P6rDnHeN6dgIqRSY2Zo
/L7EZWmhC6HAu0TZ2kDABsd+LTXxVGbjRko+GYFI4w2uFladzldD6cL/yjcnCD+I
wP38c0gwRmKWMzyAPG5dZl6mPCG5miZOMUvRoFojclinOz8P9DwJ4l5oAEkqAcbn
resXorhxdMG8DebSGFwfOti6T1PgtO9fDmdPDikZPgY1ZEvEVf5nJEkHI0pnjBG/
H02rEKJVsCN+T24Fs9rmhqP56X68nO5aZkQ9ILno10ZsN8tllEl/VwdYJqut7oBP
HwIFCt7kvuL4fky/7o1aw7OoeZ3EueEivRgezk4F5fI0REHF6LAk0Z++uYmkuV7d
wsPAAWNClnb2Jx5S7+qmrbl4fIqkQK4xm+HqORBOU7ezmky4gBv7TGWVbnBb7DlS
29baQKSV2Y1yGKUiuBV+7hFB3hrkD8JUHXpf2xqv28H8WuQB+aOdc0NciylhyJBT
2Q8wC27H+8jxADMthlnAZSdLqj1AlZzBaZs9TFh89mUG8R+8dreQSiEp18OCVwtK
0tDKr6hTLem6rnfV75Lh/suXaU5Mm5rOejnIH/v4X4M5+Pavb9S/V1+EjPRc+WSK
86xslUDBUrmIAZZ/xIRohOwwQTDTdw1M53/FEL85jcvUoQE4OCqr0ZzZpDHw2yV+
5y8pkiXO23aJfohNjcbXfukQIQFG7Cg2g0SukRiXYcmBLqvYsSAfcqj4AyZOksIQ
tu0WHL5eFfAPLlAEV0mvTORh6NNdsJH5C0OlOc/kdtkpaViXTReLGVUliNYA7jmT
Mg5VCACXRG2yI1kDN11LKa/jHDikgoNp+5MUOlaCD9YwP8xATaLbgQcIvxao7781
O4yu6psCSroeCiKo0LevGfGOI4NMmqzo+3XQsluKIjmI4TNHErN/AeIMddW0zFbO
I3BlM+hIAIBbBQ3tWjx7PbwTqUYoQ5CjuZK0e6PznNqRBaxY22QOlaCnKjuSCdPW
THmK+zJR8E0q2xRV1uFd8qHUTY5weZO5ne8nbBWBCEi7hpvZ0ZUEx4XpdV/FZFoD
h5u+l6134QDMiz/VJxNKYxBH195a36bTRWMd95+FY5wNlX0zDGbI2Xt4NFbxrF5u
c9uC0lvfGQ/Wv6Ve45mTJZuu64rj0FEQxbIVR+lSQSwgR0ewrN+QQMAoDDtQ7MSa
BOO9hXgek6OQsmZ+5GnX+j3kqpqj1kzQnHo9ae2506mMg0+Q3oJH58xkwD0/B1lt
klMN02IcyY52mJvzGn9CIqtMXvPXbBWFMp9mzXC64r9IKV2xuHEcLXKlQgCb8Q3h
ANpbBuMaUpzUqdP+EJqWEioDWtErSkQ29oPrrU4YduqAl087aYB7YLOXUxW6xEug
mpA135BKE/M/OihmbWu+mxyIocgI/Zn2VGy6jRx4AP6hxxl89YGx9n6BpG8k/mDi
hpitiIiAIMaz33Q3l1BqQw11Wu07AJnDXR0D7yRFngvBX22m3BFIzZRs0nwsTIx2
dkCGINzVFz+y9ZZBCMTrESMPwOBp38WEKBl1+AkmuPImTSL2d9+Z5zQkiwz4+JVl
C91jGBGAD16/m9BHRKIzCA0YRBoUen3QPchFTc7INWdA8xele1AVtppxU6dr7eSR
eqHkEvyYMihKhHj5GATYQYsbxsh6IR5ChBQpflcd3nSBtoGUUBzM1zlAkCwO+zLO
yGQnCbNZh7LKbYzcHfw/iUsl+icXjCa3xv6RItftUOQdr54C+bLENHqYpSboXUCT
18DT4QpE/2AOKEUqYFlzkKIRP93M7iHjm3K/dKxkDNLxUgmvCn1+cxsOe9dnTTlN
xcJ+KSZyd4bQyX2UQxM36lAY167D9aC+E99XlEEDT6ncMjyA1hYbA+af8wCkTLWI
yYdqKpe721auDnKKIEgMsrpbxMYX0+GFjsQ3fwhr/1gc2/Jkbe16Qxkjzo4uS18z
ZG5xR0NolgUtX6welJOq+A==
>>>>>>> main
`protect end_protected