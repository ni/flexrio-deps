`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
L2bRNdr1lLBT0eERw3vGlLy2sUA4VsjnABTCZ3zt2gePYwxIUu/swhOW2UfiGFqQ
QVrgyyrj8vWba7fOd+yDe9761d9DtOarEtGqXQBloNLx/ODnQvzKrGN/H9W3noeB
I9mTgwNLXAGm5DOMhm4yNWaFWJKblKKLz5g/PZ6ImmJmqRKZu0BeM5s6MhOqtpS/
6Yg8Qg9cbZY+I1iC/pG4TheQZnMlxBSwu93qovCeBVXNLXcCCOeiXQ9nXz9PTuNg
OGaOzvek9mfQuz2pgQRv4lBtq/nHDymqu86PGtEldgwhpk/8sJxZMJ96otl+346i
5EaE0cSEHQLJ8L2b7uVQ/wu2mgVmVXtd/PqT0KfzsBCmoLC0yp+0PH3s5NmEyGYL
I69efjWlRD2skT6a1t+tfUn7bVeE/tc7BKAtqDkWGPDBjheBGiSygNZM6mwmyoTv
k0vJe82kZ2v6+RMLTs8xU86UYacamV7S5LIB1V5Lrpw6hpzmkStr+H5hzpfTOEvi
XR10PA0wnmrV7D+fCS5JMhs+mVFaOouG9Nvx1JAEhi+jf6GeEsvoOiTvSYWtsH5E
4H8y4xp+burY55yod4S+wqcOjo0r33r/FHQDpvdYsFPG9A3213qdku5R2SSQ/jxs
uYKLoNFOQY9BOxEa2vEc6C+BdB/WlLq+3655ZqtoNCCtmGwgJRTkTqZDRYjb3aDU
VEfFqi65oJKSxrBVz+TwSpfxLzhe0jbQ/b6A72Ko4RpKV8WO2GYTV9LODppb7ZCy
RF3vQT556s0rzCe9jjeG/B21L6cdB2Pha/JMQX7g7AWaySytPoMzj5aZnTttytz1
OheK8OWp3g7x8BKiU3ywCp6OFwNXKpYpFMnn+KpzcQ4IHcfA/Ds8VAoBIW2/wCq1
lCx20IaTMhhnKPSMICTa5thWP+dVwryA8+kRhVYymKgqLzYzw5NhbX50L12+Mzvi
acy15fMi+MZY8lhxDUHGNoeSKf8YTpq/76EZWXu5JgFX+syg4jUewEzqexM1wPIT
SZ+ZQrrG5HSCMOeE1NYG3JEv8lWz2L1xDG4tk1mcR5dR5ApieXfk2SXOK7xhNooB
SmJN2HUhHjkDkGtQ7e15LhHKuuhML6BAmGriGsoXS8XsrD6muIvL/vgajXdCHggN
EGyS+kEbK/B/qH0WZfdOFOKnSyRGxlxh6m9fj236nhv8HecLKOOG4RUzo+IwsjOu
PWS9oeB18PdiJ3iTTTOKP2JsHJ+KMZ+FslWxXuPBH9PD/MILPF0NNPj12v9ojX2W
H0LXBz4Y0qeRWBJmkGPFdDad62bI3sejol0o5cF0fQ8mpkloUi/jRvzfZ3vzNVMz
VxBJ6EP3WgXIY7iJ42aT9vL6a8NPjA4mEoWOa7+GnwlvSqYg6nZiSk3xhLndZrzY
ZzG2dqodyNv68aEMfvg9YrbyOOLqI1+HbQC4+OuRw5I9SQ2QDH76paY1BcQVU8cy
RXbIH5AGEshV+6w+jO+cui2sHxh49PYJg2cTsiwuyQPpwj5u7oRCxZo3WMLvGZWc
lEJTv80KraIzXggtZbj4qL4OKXYxeic4LeHMLt8DEzTmyFRWegIfiegQWSLWXD2N
c2w05wB4ZFCOp9RN+pkGxtlBeUsyWajhZo4UFe96P7EMdggiKkQmch4i6BwdUoQv
P2SoVzOBDmVQHt47bdZm2UcvOpA1WqvIdIR2+aA/ZYZzJeAwNkvXKlcriXRALR4d
rMQmLZRkrh9CeWjrOJYGJWh2rAWdyvn1eN0BZBpnOSehTDkc+4iiiBtr+L+AJJj2
iJkp8FXFJ+XTv+V54JjNv8B1DojfcPQEQQL6nkdW0wa8aBSRj6Iq6IYhkQr3bKji
CsS232BJhWqubl3HlSdq/7XR73I9xcVkOAv0jVlWOOeHnnfDJBZvdEhjFoWGaEJA
QoEa+sWWIWxXGeWcaWPBHg0JRjDegUTyFFMNriOqDugHhkNsmGVQBZ+RRTvKD22p
KY4u0zyPnIPtnZ6Gf6cBZ03gNaOi16Tr8zYFCCIl4d0JbiYPEwwjcjbPDQGYthRi
J5uQjjJpO9fzIXbOwRFYJMPC03WUUMoZDpNZuzFiqXxcdjw4qEvESw42Ki/xLL+C
8bgTrgu+9Sz8I1AxOZ5mgHqZ4i8ZXYgYNZiyU3FR4+idDp4sBW2QoVfyk9aTFAaH
Vf2RQWno0Ef1AXG0fB3JIUJf+6iRghPovAw4NJPETQzcGYGj00RgyX8EFJm0rFfu
NV9womCzSh1/yZwySINK91bPiCtTJOt+jnh5IivIMQETTMYMTLY//joR+sksm8/X
+JTDVpBAOiFqJnHK9C29wi84arUpj29s3euU5s/GN2PTLU8GOtArDIuIRMKqkGWn
el52DEqbZF4NIuaHZ3Q8IjkjmWMi+Y2XcuOPSnWxh8D58v1x+Y05ATi5isM9J2pt
lqPcmPmHWOBRQYnF1hcIEW4f8u5kEGCfjIjT6QBgNNb7hulicqibc/rN0S10aafk
tQybKscJidMC6/ErZR2hSmYmrc3MlPfJ4+COAp9UWBY9xqinUQKSNqYBRphd7pTU
lQKYLmJ8DRijLbpYEXmDnjJbfhYlkYYc4bB06DMi7GtnIWgnWF4mLP4qTZ7PVqK2
7aysjtGuBym0y8u9FAqbFHB10KIMC88ieh6u0uTdIMbKS6ApmjG/z5npOtKrvqUN
dTkHMtpbMV1j1diwj94WrtsM6tm8IN/Dln2JvrXNH2rcpGWdHkGpRgWLt71kPMqD
G5ApR16e/S7fV6DKIJNc7wlbES83tM1dFxa/msqWY04iDJks9pnkW10pUoeB7J6P
Ntg+yTUTJ9mhfqfhM4eptCnzdc3E8YMUVdkdNRyEuTQQ78lahYmp40W6tXp939GE
Zt32MlAlgjnDeSOsA6ab3u91rtoI22DgZA947Thiqg8slJBjReNoznVm2SS5XKC1
gE/MhH5eIXlEfqKS7Z6uQttWSQxyGjPbfYduwSDNGDA6+BEut/rdtnDALZzZtX88
EcwNjJteWr+YwQg0cpPN3rBORxFIRBnjD8lGVHOUrSxC8wAVeUuIP2Pa+9CUZQfJ
Ar2oZpufEhFgbeRV0opmDsH/ZnC40oq53rsNLR1dWQ2Q//TZof1Q6GCtwkcAWkDz
+eZkJTrk9Gy6CbjJRc6NySt7RjC8AtWXczssdXaZkJWA0Xz9JdT0zMYyheiRaq1l
3lc4EJ/c69C/7bRrT4zwQxAdUJGm0T3z7o3ZvUIW4rae/pZYryQlZlrzYCf6KleR
wCEvBapEgaAh4W/Tgcc/gj2nm+swUtZP/4u3fS3abY/qDQAdQbpKXkzMjeeqE3xZ
rsiNkD5twFsSSW3qhO/TFAjx93leedDwmUt7P6EMIhAim+bkVNapRxxYbRuulGii
eVLy7WyIJePObTlgNWBsihWvv6vHNY0+gXEO8IoFqNQ3mXF7xg4QCbBDJWxTD4oh
PqjVwk+MpcVLfy+tHLKMlKtV/5/h+KWvIPRXU+4cJKvirEMbhF1fy6Ex3VC2MpnS
ns5ghjq+4QBLdXNNfgCFlcSQbqitJeok5+c+03faP1+icHPeq0fjjERwgxJaCV7x
JZxTZzggLqfkFNlIUmBySEF+LU4bLbLSB9PtV7TRLMHjpRpCcPVfkgElJlzTcHGV
GjIgbcfisxtSSuTOX2hPofgRu9bGmuX/16kc5ehkizraXNTvQDLfZ68FbyBt3uYd
KJ1xddpFEA3aCwJX1tXdNQ2dWhpConjzYxQAusc84//YHUD+nXO4mUINku0+Vahn
/ZHWYCgWGPDQX1r4qwfaTlLdfO2gInY8IDj9OKNKA+tFzLBon99y+mSoO3e99fBp
f+d/TQjUI8Mc/ShAy79W51dk5Na3zIpSkhkAvQIN77tLNT1aV+bxTDzoUZ5nj/bR
/fHNURg5HlW03plPezCRNxZtjpmyhzuqo+6TY4/XqqGSChEPBnn9DFxX2IXDqGsc
N4dFVy0d3pynJRe6gbQrxwDcgdeZNz8r/Wo5TWcAtTRFK4iqvTc77txNvYrfyGZU
aFAQyo+sWjJDwHcLTCQ8ZUITAMCYG6uGWMMcOkHuAfeL71aX6Pi4v1LySS6KmCCN
F8iGdF9FBnM5lC24I60hPGV+94jMK2R6X+2AxLjL0QufNCYcecC6BAXelsLONupo
dQ3pG13m1fnuFwO3GW04u7aTl5bzzi6Yg/3wJGXs5s/+oWgW1eCTJphBfU1uMa2Z
97Hl+ROJwrVd7IahqHqk0soCbFCFcAF9gU4B6B4TE1FrSA5emCZvq1vLX3doeZ/b
kEdKdRPNiTqhZZui8RcnwkL9zwAI2pHMJLEWLYSw05OYAD8+EaDWJ7OlS3uWtOb/
6lAhvENC9qPFiyOA5I31sJEEiBE3Q8bZyY+Wqja34x7h6/GWmouGApyaCqVKYbyQ
bk6hxUwbT51uNPfLz2oB3K5aQHSTVYEGHUSwrokpxsROclQ2098HeUPQgGfjFC9/
0tWAzHIfCUEfb9TyJsFCdyxj/SLEHdn74duy97Iltv3q6qdPfZKLAxCw+NFm0i8i
jqw/6wG3eWP2Mm8zYGHHG92fgyYnrKyXQ9ci0zGPzSuBMujy7u/dz5geYj2KF2CY
IjPWQdyz3n8yhpNhiUgXKfmIBoAF/dQ7R8EJAReXCjYFTuiVfkxx91OlNycu29D6
GqM0ALC1Jgn9TjpWomuidcZor+1eRkR6cQ6IQ03bYbLuVUHgGXmgVT3zl+hrazqH
JbpO5P/W9hjgGACWz5b57Dy7Li2vwnRJLBf4P/gj2hzrmtZvKhQale3JO3knLttV
4vqF9MZLPgx0oEqSXCRZCXxu+fdAJziF4PPCXnyZiWGvWKgJnX1Vo09pSKtv+LyU
5ss1a0XebtfwofwsJ4cql27OAwbAPUwJ6S/W/5yXWY2Mm20LB2T0Y6B9/dZvqNjf
rEHJGGcx9qiDhR3wislVHiwIE2Xdsjz+p46ibEv6AXnloUii5roi1uRrfErCqGOO
UZU04lEanUtw6amTRiTarXBwP/mWlRC5HRAk9qY9RiRJP5Ev08ZC0MbRjaLNBpuz
K4ao9O1k3HBOLXxhJKR6Ll7BvmH02STQrmSFLJfEMmTVctlbDdwlNjP7Z8hQwC3v
UGpnESqFhC5ODCMNgavj02shw8JbzzMSDLRR3E2s1X7NiNGzqlXxZjYx3yEB5va9
g1Mpwj+HFbuzQn+4Gi+tfWeFnzmZS5fvMJSxjawDtWTerZ9SFFgZTVwoLSVwlIwD
FhPI5QkzCQ1eADIFRUrbK3ImqLEp46lcSuk6RcRt5fUoI5uzb8aOY1Pjy/lHZQpc
QWV0Tiv/Ww3uq5rU0yXgi0DBhajQJ6xZjFsZJ1ZQ/Mzaw8KNT0EsyLK3WMzXu6TG
XIla/IHxTYkz0uluGt9lcKNqFOXa1+9d1iemxpiQoU+3ZSCJ9IuBc7Tt/q59cUXl
gcNPG63ebKLWX2o6Vq0tdQIe+KBw+9AjncUBJY59sh5JEFZV8teDJO8Zv4ZIejaQ
HZfvogFigVIBYEOcHe9goLJHeXtM2sHqlF/RmBzaRDRvJMolsE9EpGeOXFzbzO+U
kD3uW9/X6vwohYWcTY/ueJCeuFxT8Uhn5mfX4VAUjgMKvEAYTTu7VLUPhigOPpzT
O79jJYfnIytKxodfM0bzlufb7zlCfGYlFPAcAL865bKFjUUoSjMNfM0sKGS9J1Ve
78FZOOZIhqjhZvpkm9jGIUpFCSwTL2Bly4yhtX6BHCfF7HMcPnCi3JwGMHYmck0Z
a59V75wA4erbmCxt2NQPREex7fS3tExfEfAKwuao/nCj1eCVhAi9bPZymJh/yDvl
ZO80qU4tTkIVifrExN3rVE0Y8GLmBhfB4QTG0RiUkRDVLxXeQk2IAVwsgcAdDx+5
u1mLVxiNsvLNYHVN4jmLAA2LtBhhKdGH7RHtQxAYvNuEioBgv8KCpH2o4najMVPT
R0lNMROX62k2RyLRGFhm7ndvY/6iGLXiR44EkDHXR1tWksEFqqed1eKRQcdzULJr
H8wBGBlOcVxCs3oCam5V3wlwZQ1MLR8U09X9kdLOhWsaYfOGMU8nZYA69DLnho8t
13jeMilIfOmCf2b0LkImM8xHDyl6EnfXQQPmbkqFg7bsGPbVi2351T263HzPNZ06
dKfyrkwMi2Jj6Xf6yHHPzvTmjG5DmtPMKP17NYQYMgddjFbLbojKvbJK+Hqn+O8E
iuyoR0Oucoig1E/Updi6apB0gKrSLJ6/kjZFAGhvGNZhep4MOaD+4B2i/z1e8vPR
lP8ed46KShkXUdWId/Qt6sH1og3EjL19/dOWTyZoflrk469SB128wRcmyr71Regy
UWdM6AJIDrwcm+dq49Obs/yYU1dF444Rh+l4myAR4z3Vk/pOaGaM9FYZtSiXT3GU
2pTM5tWgDfV48viAsDmWgf5trkApjdHk14QAAvilub6ZZ3FktMN25IzUoT6h2zQp
qDVk+ohMl/2Q+G+yd2HaneIkuP34o+BPTNrh4aKMBdoEN4lBRCrS0d/07JLCReMr
fbi1iY2SdN7EFmwxyjWnqe30u7S3o3jJqDD9uvgzAxVsZA39Q0oInlZ5Q5yRMg7l
YpwG3Xm/gMgZTozMcfIQybzyEMGy1oX9lAyb4jLd2GbN514HA6r/SO4poDSDxRfa
cN59JK/AJSj1wZb1ZHgbUcwcysZY7N4vYETIsTOl/QgQll4rTEOkmIvphfl7/E6N
ChHzDcGgYg/1ZnuBCleaw9kM91wLPQx8HgkChOj2bf3uphg28rU+UksHsXk7EfaI
7ecmm5mIcis8MBwZYeGCVxlKxoB5NUKxtSanOLvh4Xh0WfCXtTKR8JWDJHXasBe8
LCW9VWbKYTYc1VJQO3UeyNQahD1dSUUc9cMV5JhXsigh26XP2X/P/S4vWLTHCQX8
DknOHsayUCJn1SAsRMIJHA4Epue78lHN/B7WVPRYb8BRtn8to/7kRuAZ4tpEOT7D
NvryqVjqfE/GQcqlVCx6aAVuY+jPiH801geFowABSZIDV4y/KEaZlpye5X+JTUlA
yK74ZuFOp0B5GcWxu/P2YLujaHrFXtIrVHYmeOMdDnOMz/C/vkre4zHwK7JBQdLI
HDllXkTa+o8NRyBX0eaDGLi6cme7HB/8YvWabst8UWSrVZmSkbKTqtQNpa8dfTEc
B3GFiXt0gcl9CFMFoUCf9YO5JrGe0pNlsE5nNWOVep1RN/pWy7R9Apo2msYtyXXx
O3cUsAzhIdp3yx/XPL5s0PB401/pwwEqE5lBvUAn6/kccyJw93Z1Bsqw9TUkxMgD
KwXOvf/v5nsCPeEJNaPVKJ9xMvbeFmAYnnDtQybScisAnEA79kdOel4EcAkOkJxi
bjD6UvHVVzfF5a/k3V1eUnUb+CfsubR8jSHsKumhwwYERcv1Q52sF1mJZlr5aA93
XgES+PRJ+2sOm2I2dhZmsCRywEdTaG6q37FLr7MHV5iNUE1f8dLHSkid87EQ+xMp
O15IXoXiPsoylAwhSS62EsnWdTQ9JEDJr9DucVPAGUSqQ/aCriNDAhpN7GtEnwFS
2AKBaWKV7dbSF2Q6mrLHhd9ngO505Fvjs7V6yN3WMC1JmvhXQkL/KbnRMSKK6VTV
Hz7yqnJY6GRQ6uv06LuveoZK1ziPkzGX71PpVoF0ph8w2FWa5J36hyGd7zr6xCEf
KA2ngzBw1ApfGgcmqOggbDjtcO2deRP1E1ZBT8H+qNm2O0fBdbhkoclJfw4tkIVX
qFl+S5K23l9LlJpzuONynQOXU139zC79pUsq73UQbaqKiJYdoLz93nmTJoPCK2hF
WwaTmVoX0HV80XUiL24biDgyqgwGbEKFxEZiczUJADnEvmM5x1PbdlcyUuyMAttR
hTN7FA/pQ02HhB50e4+nY/AAwbpvoQR2VxqWgSP3IPrzT3vDKcwx5ftcZRX726vL
UjXKQTyPaA3GAGZiEfh3x6o+J3GGraRJs9tW643Vm5eV+kjShl68GHW+U9Mx8+6T
Fw2PYr7+cZ3bQ+RCc/X/Vwnxek0RrOszeCJIBVSMz8bK/ri9iOIMuwk8lgax7qg7
POcAW1E+S1d47mqERR9kJsPFsb+vSHNmxGQ0o9bSfi1/i60xs/FVjEroLGUZ5QY7
vGIntOnxBztZm+zlItHd4hTqvzndKdQJ4tnRX10G7w190F++pRbE4Ndl9ySHgVAa
4/LJQ6DIPAhw5TwcbI/7PUoIdaGFxoTSfWajSE49iENRcoSobW3ZzhCEncK1ge7n
T6/IYffWMfDjFTroKuGv0+MkJggyZTf13Z1JQS1P7XYKNIaBEk1jCfbppSJRTCeH
1qB9Ywsu9lhqNPNfRxyoOMalynKvb6mQNPwRG57P0Dx+Ys4yYmBXK/Z3F5P0TYJQ
kEGIpKbGhJQbZSC69gb9GnqmW1c0ntVDoEDMFUj7PYPakbKNijS5il7NocvQTmMH
RxrL8FfIaUPnA00TJFow+NkoBbQoq/dhHYbw1zbboE6+0L6Iu5F9mfkRGNaYxnhu
V8CRlnXP9qIQsrTWtjzf/Jnaib1sKF/AAGcFVY9RMbMvvuTgzc9WD3CzkjmuGvmy
eJdPAvDbtwUcJkja7zf3T2IcxA3vKad2D8nSX4qF2otZBoXiVvZQ2Ngei+Qs1HJd
GylMr5DwYfh6mukD9bpDdoinLzrkNf962YYTc8rV2M4d5sPgmsGr+ITFq1EVdoUN
8OQtClTOTIh9rRcihEDVlAUxywjSCH7i8XxS6WvQ1ukdTGjFIFhOtRu/vmfHfP1z
YhStz+J0tUGjLaFNyYgC7N3OMv0+tic1MvnDEiwH1lL605UDkllTFYLQBaEFOD5M
cLpDWfyhY/rmQ2/z8vrVbQ5EoDHtU9X5amN7LE1+Sq04siJG1TMybUzLh+LOHV5y
dnoJzJvQ0yjYD2gAh2emgSTzwX3ND8X+SSH8ceZhNruyVN+FCGS32Qsq/rt/F+hh
h/1aqXjS+XUxAsa18fNWw18G35o/dHzFTcdTlnmJF1wy1CQ2Bxzc2dTCTr8rgg9p
SDYKRiRndOBLPJ5jkzIFGhxzVJ7vCF18xplz4LjWlOXlr6AoUOaMnudPneXikU7b
WqLjuE1ESpBsgMAtSEjbhZDEFc0h8NRBSfKgk+RhT19vXKIMJ+82+rXuZ1DoAFbH
tt9R2ks7eQSOMntYjLIqcAb9X59Ebddmb9BZAufopd/T9uFoX/0lvUNPbEkjDaDm
LGY4uU/yRgrzAhggGvarB5ed0AeYiruQLwn0oJc8XsPi9M+P88p7WT9yhsKyW/Sv
cyKd9zmGV81LPxEddApaxyhuoaUqETNYv7PzyBWccyJoX7q5y20HrDNcMDc6clVq
FQNPC3AIbCIGCVSamL9uJwGH81qm0ZCWr7xCqLvXtGRi5IUmxZFrxA+F1rEvSpcC
ZKPvISrA+B21pZOpbA+q0NAtp5RhgjALb1wjlWxn3VcPsTq17ZvJ1fmEmUNzJeZ2
r/+8EtysCLJQ2GyIvrlRqgQt820cbHHFsMvC9jz+6qvh2XBRjBmNiq8iYbuLieoW
v7/aestW6eAhSJffXXVjK7XZmEneIBQf3a0AyBrvq792GhGuPK39D4/1aClF4UZl
SJ0SsrmDc4v+87dwwPAIlMq99I63ESID37o1q66Nur/4FIeV/QDDd5thRQt5WSnt
606zT6fK5hMoulLrXfYgQGRRRL/Q93BvsmHNG2hvoIgs/b14Dx5WdJpRVALX7YSh
qqSSQw7tCHMMWeoTCzASR5yCU70+YveS1tDQbQg5ErVKNdBy+BrhDnF3P4Tol0h1
pFAmOwzuyzfjYPu/z0FJM0emd63wVPa89ZdIfMGf/GLYQE0gBhcxoIjaavA+zKj4
N6t2l+fg43hS/oEgVZTcZ6vvQ/pMhExoa2AzJ54z4+ICo0vGC+yH9lPD2iQPzMUX
SYmodTT/r2N3FaFGuLtNHCbCM4a8mfxo/uFlCo91n6rwzRGueFcWaWNKLVbgQ82T
40fZGmDVm/Veqj1RBooXimcw6pUEz/1v2YEF3558vogsBTR5lpn1TP/6GD7Y7Xs4
UgvnXrwxN1MBOPHPWUlD50RLIGhK5ygqyC3s4y9kZktakvPTvHffEAD2M0wpCvo8
rcIh0t+8gcS5Dpt9LSIbk3ysAQOowLw30WZqwdMgdS2I8LqqbaoCJ7aNkfzTFKy4
tACTOlKbnkiA+3VY7GONpvbxrYw93mOAYhxgiNiWFat77PcnOqC9H9/vnh7gqmNB
7xMB8U5As20U1woAvayI17UDDjOCpiGWSemSygHbSaSg7jyr9A4HFZwEnG/eq/J3
UKU/sG9BsLEhYIlCzJJcq7maAZGhVmqSUUQlyXaN3UVQkIfrjDYZ2BvfGxUsoJWz
plUhV8gj0fyEZxLQKt9mXCTJ3CMP3OLzM1+bGeohiT81kPrIQDb9GRxyNmLaJuL+
U68niXzsJjuo9a2hRk1W4KTIQUpcThFIENdUpEkr0sP9L2YamuRngX5ck/ENWJus
gVaGVn1iWL6yuHE0pII+dDCKOZN/UzfdEozG/Ulkvjdcqzdx2x7j4XCd1PQq8KBu
A1mIEDGzEYYYXW92bJ+NuKLK7t04EPj8zzHQztZo0FlgZSktNV/9t0bWZKn4tBi5
PtLnbTuMK60Zcmo2yqlIOOOUDlogO18Tf28YOSA8BpsB3XP/b+tT9LjfEdQRROjW
eVYfIFMUDrILD9OvXU0OqyYdSwrI2ZyuC1gQ/cJv8kCApexiYDP7Tdsb9e/CjU6/
QqO66E6uPf1VeUfZ6RQm4PvSJGJqWkuaSnYe2v2jgK7MORPHtn7z0Xl7dyf7dSxi
fwicm7oep4ocfov+Rg4X1X3+Wbj5v6Bpe0/N2yLTbUsa5kgvLfKgvRcqjTbdxCfe
ERnCVAR8GE/tW65L888/iXIx0MiDwXdWhIdW4j0ucWHRfbG40HzvJiHZ/QVHPHOA
bQr/A3L+NOr1oNWK4WRET3laWkyrapN5A3/Hos7AYma/NG/i2as+Za79GP20WS2d
2QwB0UYOxQ/62V0jxDsEF7h5RIEsNyP6qtn+yiGKnBkGOay/lzUbOt2S0dfj/L8W
vWhWNujy2XYIzB4QL0nfYs1ZhqXwqCfw7OSFV5NlOhONnvkfYwp7NXBRZP/ZM5BD
sr8cgzv4YzYJ/0aKo5kU69IYeTf7inyWbuK5ttOQuCt/gI70lkkr7Uhqp+STijdg
gG2kUZxWW7Xcpj136fAY3JTektKxbKDfZt6OeGm2FJI5VvjPIEfuTZSynodB3Fzl
kp3uaNTC7G47lXRAJ28NE4O/dm3Xp0xqjA9dfjxTtxJLlOlO2rNxHQes3xXHXYZf
iMWTJ02TYONVGkeIk0tx1xhyATis/W4nbC7j2RZq92tKMHTMchrTJ3sE6CaEddsM
Zqa3K56abnZ8T8jrVSwLhbWXGxk8wEHxRFeaaL+mcABHjrNvEbJiDETabJcOfJRD
YQF1SKMpN14e4tNN7bAnZDE3Tyf4lj05Itf6Vz9yARUg+4Ucqhsa3m22PXfcQWEA
swc5KX+IkwnDpKcdRskCpR/0JW20ufq6NAJTh5/AYJAOMHVglbOS+CPQqEQ3eZgP
EnS6GjYtH7esjCDgddu2OTN688dAjzQbMsIkiMEL/TKp9qI64/BNAx4ghIdBCbFq
ld9W2WuawlYPfPmyXM2CihoLn5JCiBqLgqGyxMDTAgJi2oETRldfbgId//a6oxfM
NbiX9HCRWa82YXWpFnPAJkhodUOr/Ntv1kSdHXGjreAt6fY0ZPI8DwvRG/ztcEwn
7lIdO710Zq4wIx5pb+MdhcBb4UmRYEXdHgAVyNkfqZ22KlwVILA2bhc0VQiOqz9g
wpAQPMiOWSFKC6T3BjVhJbdYAOvSX68syIY0hssP3FMaodOv2VeNtklfKTp4/4jv
pvlq0U3CISimN1kYpk4paotaGQwYClaKzxc2eLVivU1X4VL8feK9Y3vfvjm4u7D/
x8Oosp9FgpksWg1iRAj18XyyYm7mSoCd77Xh7WmDuLmXMS9tGLby03R/O9bMKreL
pUVLJBgqUIv5o6z3Bl8EEmcKJX6Z2kZYSoqih+YQIzO3fJ4ykU6lfAUhI1rYs8HP
4Mvr9U/r3dlRbBdOnqv2tX6URKOmvzB/BI0OXWgS01nhiu1lRLRVClN6GfpQB0/c
QB1lxy2aKU+I3f+rkZw23MxAkLO+krdsosW4FyH1fs6i4stIfjmhU+qsIidNSFdB
yukR6EbKyJq5uWPyYohdMLMUAliJJUNRmWRl+dC0PZEBX2ykmzDHFmJm8grfx7fO
2Wj6v6xCfLNfiLpUzwjLqae6SwcIyBe20+CRzaW2nrNHVWFRZ6VJVLZDB17qCxjP
dYVUg3iuuzSrE629O0FKRTQ2TkckdLAiW2kz3iT4yjLZBBkMoPl0D9VLpHnp7lHR
lKn3gsEp78nHXGJm8LImtuuDJhEKaOsRuwnqxqkncub/RwYdmr/Im4LczNndK5Z9
dcPrkPaQJ5sWlzrss/4870UxngGD9KJMDon5URSTfgD7gebCBYB+3xB9YZhRlBtx
ESqUEgZth0qfj75WfanhieFk5kFyE2vLxt4Kd5qn8+gvmBTNvzLY6kBBFJJ7Wt/3
0Gg68/ADDRBrr0OIy2msixjXitrqdskXV2Ai4AYDh/oS9TjDWQKR26z4Pxmg9Gxu
FNKSRl5NbHRRSgBah4pqE48yCm2jnXbVkso9dKLrw6LHMLMWDrUrT6+HgtaQfILB
APbSZ2Mkes8dYzae/fj17CdI3vN8JkNUaIdhvK6VFpCnKX5/SSk4acNWJAQbqdN6
cT8usW+QwR6dSfybpf0yAAHIAYH15WYnA3iOBH1Yn3BSzhCRgh8Anj6o3PUixIOC
X4INp1ymu8gtD9n4OaXoGpvnN5F9HgR9R4dNvlkK3suSMGZZufZT29BItdB0uxR4
QzkOXELoAfctTkTRpw7gqS2S1CbvIDW4O85pqUOEq2YQq9LQazTXKOol23N4/5/3
Gce81RXUnR7tq15lvn9pMrvHnLDqjRTFYviiSdVgjYcyLemcL4pIyHgVOq9pNUYr
FKcCk+lOonx+SJE4/aPHBI0WvNGuKtWQDjN4Uh6BkzGHH4NzOPBBz9PDnn1G1171
q1/kofARr8TCRHMkNaE3asCnJ7BUy7ceV6rpSaYBOrL16X35kpOLJCnJhs1w33va
GFPd4g/zqkoLNNfFpB/+2v4baMUpQppuX/LaPaqHvRhdWzBQOVbs1TUaHEbDV7/t
WKL7KhePVKr8oh/MCqqNfbLQI8CZajKFQP0loGSMhy7TRwXg+fMCfXi7+PjZ3j8T
YNX7MAqej978ozUULiRiNvj36i7sKNhwaOF6AkfrlePX3TeSPP23FTHdPIM5rDLV
rnpR9MoZPKcbF8U24FzfYYmJ1do4xlH3MZ+JSz3MzB2mZV4/A51jfRto1gF0X+Yf
gmBKyqEZ/y9WnyRjOaCPl7SpJF9Fuqj91unxKn4eSWqNffvM5WpG/fNTHALOzWaU
DVGXRK5IXcU628JgzcwGcGLNSeJbnPFGLuIj7S0YCfgsvaSYA1OCHBYb9rXEGSL5
2hhhYkubgPEJQPtr6uf1ZnoeC32Ze8TtG74HN97XqhfOhd2/Tj27bzFHierX18Zu
F+XYq3JNG+j6lCXHjHE4vTTfJqlMT0B9S/A61DE5AqzZXt0vEOGIM8WuROLFpNy4
eeUgd7ISW1zc24QwCxHpV1r2mBAAYkt/mcJhhpgrOfSfCqEum5/n31RC3wifIf8A
31ZyWbFaRNE8zAHUxA//wr/+qkZ01qc4Xh7iW7mBxC5co8qzz835J1fjHlEOPYHV
ApgSMGF19dtB3N0oU7Y3nSZHEl6CN7EiuRo2CoVlnsM26eNOTbxaIiNcUMOOxsoE
y0UcmohUy3SeqN7K5MwooAJ+L/rSENfT9g5EadywdmzQ1GQ4XxGit4QuFv6wbMbQ
a0SdAgivnIcOTSmriVkmoKnQ/nCkjjvSgMmakivAoMM/pRm2zkhBpEz3a+1biF+B
seuDFMpgmqjvkheLcKX0OIHxWn/16x7myLcjozqBHxeTYXeFi6WfsILE8UDgvI48
ERzIEsdPqoo5TYNVNrKoGIvis+OaWt21Vtb60ylgMuzeNgkiafTIbegDp6A2bFW3
aaPG0Qfymyb7QgNRJJJ5wsFr2XHlPRAoM5ibWZQ2yRC8jFR0IYsnmdRoYmA7aK/R
f33a1CKb9JcgO2LzNOxV3zfNAYhFQXFne+w69GGkAW5O3zNKtErQr5aPS9EEg8OM
0R6ho5cu5G9nHyypZHpHTRqF/eBqQOXeeV2WNOUX5LZYsXnrXuBGgaC7ZgjyK+5/
ZxfAHXrmh0ZoTGOTAbS6DLbgJshZtRL3cXNE9mPqEazaO/eJLZYgWPusDkwIQGI2
R9cgfZZlXvlol8c6dHfcBDtwA65tOhP3iAeCbITl8bTJUmkuRWBuA+Ydmw2uEAqZ
Kd/2bLm9Vq0+VrBYyMWGgTPvdqUtzdJLy1JYc7VQQgUaP1qWtgqJgw/MgBz/B460
i1mI0cDHbQXhtC7zIM0VplFrxkwgAeJMocT3h/lG8a1QPZPDIIJwOeAUU7aVrpJo
hc/pFrJdXWtOjg32o7dyN1M+Xm4XnIP2m6Wefp5KZD6ohvkLELGF6Jdos/q7S43E
pNPhl5KW/QnVvf14rxHOXL0jpzaMVOy/fsg2Bnnj92LlLJFSfx6l7DHlOhuY5yTo
O+BnIWywW4jtDSlEbuCWWvDOzzpfkxpCLWoNXpUClyaUUMVb2cxB1NyXvol63rXF
h6b7gmEv9Cxq2SjpBFyiSRfsdPBj+/NrifQc6cIbL4Gpa6czOxwNaK+3I80kKHhu
SX8W+FUNGMjDH7YufmVhPRaSqcXUGJH/d7K609ZcOtUP4mq69UO3Kk0nii2vw6Eh
1gev0We6eIAznNQxSbdbyl7kUUDFVzkuy/eroE7t+d93YwRpORKQTGW1Mpg4ntm5
Otdsy6LS2W2LbT661j5XvgMwL4bksgHh+ORwApVC8JCpCerBq+T9AjovSpDxKRLg
DZK9UgwrcFVzI/WwtEpQtpwXHhQvKcB68FomWtsuDQ+so9tIucSAQKZqACYUlG2D
B8KoWYzXdIZ9qNJ1gPNYWQzIjbOf/ircG/TujU7kQrBQIqSbLYDT05t24KJHC9vs
b8ndNocP67MN2Lw0DE3J5Z/awqMk1wFV+g0lE1xJTkIS+GGxpUdTB5CMFB6FCL15
rZ7uWJb3OVkhly1ZFBqlnnIpiqWHOIwXtJEMcUpHfcEQ26hCp2gCwLlUv2R4ylTw
WONAJexAuOuj7xBjkZrHgBiZsxsdi/lkC+kfqlzoEZK29cLdb4YR/ht7CLMYROff
YO3SBEVQRSlT3yxpwAHSmTYMiqfcNinDtb64JWciZb3ZGZvJZufvmgMp2M1uDq1Y
kkNs756C8uOS4n6isMdyeK6mBbInKXcZUW5hLMEC4MhHu7AINwCuhT+0/cnFls8a
ht9otIFihZtJ3dvpIWYlwpx0AqoIH68haMmkUVqs3fha7F9jM1xtkfkf5ygafvtX
2V2X8QfCC4RX26IMKi+P+NZVMQF47LDKVe6oSQQ/pIlnSDySLvwc6C7xm8kkuvIm
lQ6unQBDHBTaEp7v0tvysqHMwRBcF/zYhrpzQyXxaTSq9AOVShqtq+Lw0nLS9AUp
5PwKdsaK2gus8UHrXbZ9BJsF+c2p4h3Cy3vTe7nkyIkZaGdexeCEgK7gOJwgMogG
hTAYCj/CLhy66qXHlp71jOr1gSCvbcW/2HnnQIoG1TZwje00WwOd1mWOOqTou8MM
D78EB27LcYakmP0figuL8+Gy1rx1sHWlgvSSwS8a5R4yhNzJo4IQFVa1shRRzW+i
gB55pD3CsE0vaXmNYYM2/njOal14Dy8cX/sa/QRLMXfUrd7oW4pCUZJqt+Qw/BE8
b9ycPvFHkKbk2EUDP2rfcfdMW6bDwtacLHDd9Y5xBUYunltZwtIkq9tvlKCdIFl5
YXajo5ew1mIR8NgGdx/wgEgpOFjvSH34uvbalL43m+x4eT2V/YBw44AiBereT8mH
8wj+0lloO2nzf+QikgxAMeNNgaatRSvgcnHSodEwscUdZJTV4WvkEsb6iv6Sa82I
GzTatulfSKWlCLDyjinUyRNbe4+/qL/1qh8UBzeI5NetQ5D/cJg90YOtljsSU5Rw
hpEVuJR1g2kSSepeqnpbTX2NH2O/TZWblgdKRKUZlF7TsBL6Rbz701wRX/nezHU+
X176kUBNM0+R8XzD9I9rmmh8avy6xdNPo2kliR1RDVG9FG9r+4H1ZgY9W5q8DYGJ
kE4einzKvIHBtai7x5AcWGrFwlPhXz39tSMJcTo4J5viqotGcCKf2nxgbHkoZWQM
ZXRtlOyYVpsq157LNj0Ay3ZdFzO4X75QwJc5ECa2Y9Mh+jwEtNv2XNSBL/rImiUb
NhYc9mhvXfC0YJ8WiVf7FwyPgmtuwspQW9vibfGaUirl2mmUbg0/R6IcflTOX8jn
AvEvuXyoG/8d/VZiLO3Fz2ZEN7IcS8j9fejTHR7plwMKVWk5mX3SThkxNRRwKbtB
CGcaCUjrqdQMEL67NM/g42NhtQteXxayDyhsvrhN1Qs9GmP264v9oKWu+TgqxdXE
2SWlWwur5de+GzrUU5ilsZq9FaiuQdAiNjoJFryrC1sgRyG5b4jgpff3llwEe3Za
CnSEKdo71UjKqTgNA07jbpYDtL5sL/8i1zEYjVy+DRluOcCVwu2NyWjoqD7bGGnr
KO9uuZJL1pNSelQw9NFheZ4I0paMBMg2SeCBm2eZqoyAReRRoM576lMcQCyN1S8h
sZyn/z1e2kjuOwQ93/Hr4EY2kioGNmZmAkNGZ64H8Tz2DbF1UpoXVUoTIJCaFMiE
Y/bpcgcKioUki0PCO5/9uAZg5C7uqF0LrsD2yXD/ffkQUf5Kx/BR/ClN16H/933w
Km9Ljtyt6jFWGR3gVhKsy8RModl1dWKhLmSHfpCXgDSIdfvtWlp/LnAyk0KJBs46
WO5NhkRka2BPT0TiGsrxqyjopoUgGe8+g13ymCCZeoUtNzU50GZSZUWU1ZgfD0KY
wZDwV2SzOdMwLFq7GZXXdJRfFwy0tMuTUD/3KFseQCw51Yf8Bhq2vTaAVGY0wDue
YzwQUnu/nXN3xMIYIgg7WDmC78gL9hBq43zYlAoVbK4NTmG7z/Ur2KEJ6VuK5Xw8
8OxkhjkJYzzZiaMVKuNuLgeh5FB0UQtUR72ZhG9mxPPyr7QsAfREW1slAZgYRGGO
wQRNSDh8MjLZaDmEhCR/BaCAzEc6sKPd3dnOam45Fzziw5yYByuaRy8HebGoWZAU
WeAwWZ0AJk8fU/1XhtaDzJgUI0TdaGX1KEvSaYDxjn8j2LJXWEo0zlpcJ8mXZVCM
hw3BrAuY1Bc+14/B7jT9ZJlVRYo24UooIZ9t816I9uW8wnyKcS/SWlzOfoZSAF6x
yB8Wch5GgSruLFH4zaT3TyO62ldu4Gn4OjXZ0VLlYRWH52vAWg33J6XAzRvDhr7t
7qH8/pVrW5OhErxA1am0aID7XKwrAWBQgHbYFgd2uR7yZ8EOSktBVyTFY7/UEOHt
SMkoJsaG8e1H7Faj70ujNcLrWHcO93Ooo6FUbWpCUpN38svmWrmoO0PZXcCV+096
n342pAHNgiHU8kkoEGdZ4aPKmSFpbOF4o4sHNZ26iZi3+k1yBq35MGDlOOvD0tV/
aKSrMPVb1pxfgny3wbVfZ7GP7bZwDcmsFbAHUWMc4FhTIVtr2nlVHovTMiB+J4I/
Z/tkLcYWPn1OwabDaD9NMKiLi7akOKQcDuSiRi+elWt5oppMhMGlTM4C90UdVnG6
LLsjQApoLt2oRhoG9wNyyZuKZo1s4tZFV382cPm7QfekW64czSwnGTh3zP4B7Jmh
k/IV/76WTSMZmUH1gCS8oUD+cpboDJIK8EdIvweYJxlGK7Z5/L4iqs5vsjCcv60T
00k+iV9H7qvSvFankK7IHRiI8Wka7zRy+FxwTlyIjGJdzaACv2B8O4vznUl6A2bn
7LQGL23Jd4D4mJWU3Wc9wFUdE3YGw3kE98p47UZFwKF+IwmuYukKRTJaAnLUHki7
2szov8pdmUqWC2IRB6fZAgqEMKH+f71B3wn+KnzrGaKf8Rwqx0XYNUNtfZOKxCSS
8HwLxG0XWoJKTR6vaIboKkpgGR2WIJZlh0q1traqO/ovgrwEpr+OTYCZf2hG5bq7
W4rqlCq7Bt2KIyqyCKd1lp8JAzF72eMIjQVr+DYaj1eUKqvo7X8aZNB0Ur4Gd2br
qDR12oTMMmuXGcIvoeU3wxEc1WudY8/F4wH/cmdKdquVWux++mHKUgEmmMnIa5x/
jKeiaqPQsh2o8L5dhkBPAwjzOpshUEUs8yu6t4bXmX85SCQBKl/RileBwIN4gNwR
PibKRA5k4eCg+q03cnimZ8WEZ6ytPsfnQx9uJlBfS2RKHInYLJ+OVUoADR+SHk3B
yxiWNMc0aXwA7g2QASarmrQlOAf2RMGCVSGZAzLCSA0EwQSwL2rr0XcsjcxCDnvC
2bhBPd1QNk42VipHfu88V8nWzsjOrEUEC5ATXtgiPbNJYiDsZYoOl6qPTAZqIWcQ
XQGZpUlWKCl77FM+nRh7wrvZ16nZGc+qHptcqCLe9xpnBc0vfIUbHAbuH9u1cIDA
IfLC9P0p1lmN1z1oKM8aoxXMVcLW3t9ZfMZHuDFYvZ85LsfdeSS02LeS3X9GSLFP
BFzT8H/H/uUOQ1CmqjLMrVXR9Evr12LWo7RRL7qQ4rlruFSYUYepAzzoJeNxXWEo
yhNEp0ClL6/h0qri0Mqrw8RXozsMUXRUswe/nCkmAg7mu9GmMiNSkt55ubmrj/wq
c3cIO2aJJi29W0ECv/720Tk4FDo/dGgGI3GAcltaUAw67C1p0trxMAsT446LDiQq
W86TBsUer68KtZ0YlsSWxZKuTvJYoapX2+rZJkdvzcN0dwXKydDPCr5T84IS7y8c
rrAYXlcRubIPOeRrUac0dDGZRafIh/4UxvSLlSr3OzPfJCZQHitGFbDzlOGeYndb
VbcZehsVYsPCiVTh3jtuLbvo3tVzU8QRT/V92U5NhjvJeBXU2q0O6S/c24ilZ05W
jkwCQpMaZpacrzXsMFF7WepNQDwaS6Ud5xy7mfXfcSyKDq8Yi6MnsOKkjfLWTZa7
FRZdavXFUNFLU5WOxVPPUVMp/Pr0WZGEeAvcamdg/vvfGQXSPQcztRu8sWo26ddg
pJFJVIslHkjryXfb0xQC8SIhGQStW4rwnbmpVfYnYMhb9VZ0JEtvkmMiy9LoXJZQ
PGP/R1HMGvrlExK+sp+cBDgj4cg3SodTxgYMEtVxa7JJi7CiaTMF+uQVRWPv8ZeZ
E1Xb8bq1Kpqqa4Kf4qVRWh4c6d3jwC1a7H+bjO93BvchZHmlnYH3UEqgT/B+DsvG
WzSa25vYOp+enbuFVCb8xQLDZqBOnjS9GzIwqVy+i/23ADa9F6afJaacGSMqqZxi
Fzp4UrTRz0HGLuBjrGvWoslADA+VBUoEP2g/ELQi02vkA8HnFDAS2C/DXoBJGxJg
aB1+JJWPT0qNXw2GQRdavp70sM77QocNxn/M/UosYPMVjSFuXZNhafTlS4mRAqSR
aYQYVlUsMmNX1YPWPehqtvL4SFxITTTyQnMvGuAcdJqIUH5t8R/VdUClF+LGnivb
e4USOzwIgNXkEmSV9Qhp3Bkuo6tzg84W+PBTNQG53QfaRmVfoTlzWk19DRk3HDzk
vBeGl5GPI08N9q5b18yE5wH2zu2yPwWvVUnQiUBmJTHoJq/mMnnhRv3LaC51RgNh
Osa9Rpx3Rp5Y9voiQ4RADnmWiAFCCphvzcERw7dUNJMtkvV98cXtN7AVFLShY5Zh
0tK/dERUv50dMp5C8p99iNZCBRVzJPlI53N08qBJP+OxHUzLQBGoXIPmliUIssg1
iJPiY4EgoZL2ZIqOgum4aPl0sin4b+KilF8a77vWhUsoEq9SGpPJKHYndeP9XO3L
lYFyM7N2pig/3Zy31MEeQ9GQbymfjAaA9jBNnWURlhOU8cyLmFYy8noqqTcwUgUY
covcAenGtDjBBBlXcnsi9qHNn5WBw0JputUnjSYSNAKxoyLvNeXHjMxe7N17bYOp
1FghafrsKtWJpEy3dSnKjjldm4AI2CPJXD64qS5ESZgKEGS/BFQaRgeSt4a4HDNu
wN7/+SbyXWB2v8Ikac6IMAnN9VhqBlImoNzuwy2PVf6maL0k6CRAEkZxt9bqB+Oa
ngk2ypPGStdX9kN16WIuG9BsRCkkq9A8nHzBK8AH7CHWpFy9gkC9U6YMlP+0a3i8
V9jtcdUmwhdSO7qQ6W/K5s95hxJgRb4GrxQxjv4C5pB7DK/xwjOqyDgnnqOhV5sP
E/cQSi/X+QXQ7RuPwumI8EuViNlp4jYsW8kXJgiDsysEWBQEGBjzut2txqtVOtlp
5m3uedqmE3URakzmG+BV1Wlq3wx4fymp2cFKJP59GgdKYoahBth8FPNijJAUtGSE
zg6DQjnuRabIVZzv2R5BwW2NqMXG7Y2lCntP6GcLwCZ0ggRxRa0sMOWmQs2nO1u6
2HMatOs6Q7XvZAsnw33/pknaClDX7vEcaxlAP89Cq2fUo3hJY2lGeotaNIc/5+nT
aoaJptY2/L2+saJmQzJIPA2Pai9R/IQv8evAfrJ1yPgRS6bBEWafjs6kjtp6uVZE
VEBXsh/mALoUioFuSz29BpUhu7NnqXPortBtkujcYmgFbYUwMxtR5aaqf7I+6voL
jQi5tDO8ooEgO9/St96FzXgmKM4M7AiWSBB6+zOAu5Es/Fjb/W0eNhiRmwqI8FGH
F1GYthrvyymTAhzH3anjDxcgvqe51fFr9fu2aLlRaF1aXc5xsKGfjv922QepbgOs
4j3ou4+gvvX5J5paPHt3lbXqn9zPWIHuVJqPJffy9k8sR4tLGYANQ1FmUK7G9yud
Zwv7cEnFZnlqcGhSnsHIZydE2yJmVKxwQI080oFqAiKfebsDGKdwGajr8oYp7Bgj
Oe7QP5NH5QGUHxYAhl175xcWRjrlvDhx7Aqhf+0NtWiRcwX5GKv86sCHvTHlL//+
P/lQwQtOdWABJCQ3GECQgHJa6V602DlH82W/Pf+8+MK+35quGGwKukk7/WxSts9A
2BxXPUglq25Xm2Xr0ra+720sMwmZC3QUGXqwZIt4ngKM+rsARAWOPvW+WZdeord4
xN9E3jdqHVl0Tljt6Mc8ey8esIU64g8kwx6jVHwoB1cOZMCt0/JBt/4nWyMHkUQP
VIdx8699A60bqmKoFksOsogmEQertZ//LiK/dAmEzNSYkeR9yhd2b0zRqh/Dzurf
XLe1S9xe8mAos07hnkUnkVKVTp7j/ZY07SvkbjNNfwW+SOuTijvHZ9ujKpGz12rE
FbAK+qVwjimKbaWMMfegS3onEes8XDwcF2DQ70MFCe3gipv9ncPSpkvL55m3dF1B
66OemJy/Qfm89/qCCwdkGl7P11HRgxmqLzg37lah2vG5/r4sW4EW5rHgM6YZZJvd
kD1+BWA1VeIgoHbG3yfCwX5sKTkWYW5OXzQl7tOBjaQVM2NMzf+OZlswt7D/i9Fz
XNgTwDU31Q3fJSmjWX30iLn76LAv9YEpy/1c1N4Dsimy4fGk3BfZFSeDCrCOkxvN
yvsYdcq5D+0/lbLbojWqcrmZg+xPQxoptWqSAB1a0U8npY+tdJrS3rg0fw8CdjjL
xSX0e9zfsBkqjlUcZZD+tF9SKmPR/Taj4sKiFfLdqSgWH5+j2uLhr4Qzo65CMipL
O4kDqaoThUawjnonOxoiz2Tzxgaml3LInFo05AavMjQcKdyTzXkfEQig7h4Yl0ph
kLPBfwvyTp3wnmlhqKz3TfyPIOpYQp2ZujxbYIemsuHs2KnoL/2ks+GEh8ANGEHw
Lqxb/yPB3hKwkifeMW2daJ/tasdfGzhm7jp9dFEdLXJJyYxU2FcO5MSR6VBLHoaM
7xdUghc9LlfDPWjp7aNI3hvmm6cXTS1I6aeptfBOFGLQ9tEq15uAjKf9CNcpZPCN
hvPCq3YMkTAvGSDiY3g10NHElNbRpV4FfAIdXDv46KB7V6kLRWR2TRic534TM/ND
fy6/jU9rCD9yvspKKyOYcwjAkUW9H/w21Mg524Uo75/FZePI2SkHEm0tqt3xaj33
XzbEL0SOn1zIbFRo/dE3F8vlEgh96DinHMx+6EVa2v2vgT+vYoD/Xtr4Z4b+7E+Z
Yw1+tUD8zR2JAy54PEn5EFu+3+COu6QfHPCOeRIF55PTfo8Iqct6geuPJ2DGckvo
YcL9IHLp2vGgruu8k9SSnHTjU9HPwLL8mZBuXaThdsPYX84ZZ2CBaxr0KDJ65NzD
/viXIWgKyk+xfCKYbGjeo43/zO0eACrjJu1QRI90NJAChkVfh0LXLr3JJuj8wXEF
3HmKOAmEGK877bUxtiHwDdzDPtKq3lsP7RJG5XYHzUYLs1twqSFtMam6k7MWgXnT
1NEa0vQni+s0kyWQNMIskXkBLEmEu2T8l8XOhuVtueplQiESaQdVfId/8LR6WwPL
ggipaQfNGqJrREOaVdgtWJnsH3LNagap7zS2wiARiwsyfYDGuk/ujXmCqJyMUL1p
rqZXLTs9iiFesu6TEtWEW2kLwNKLIjtaN8PZN3F0bo8mWOV3E70RC6uRMMefcrPc
bQoXSLY6MjD5Go2sbOpklKYMIR0wliYoOLdZUl6tZ388uCmKMiueHcYpiyEc61Sb
3s5PmoN6BOl7BnEyXoWVZNL/ThbJgaix/fg/g+ssce50SPWZBPF6oW+tC6cmjM3G
o/v+DsTGqnYl+gMl5yesB9OcIkl1lUyAZBlmga/Bhk+8B6G4Og7IVCdzJTVe3SV+
HWvy4J1ULBWYb69gUPVRRaLre+lrmeiFxpFIjrn1rKcTwYXaDA8ID78VQxX9ULRH
n3XxtAfwB7Md0RTkCwpE8RPVZDbtY/8EUTZKIzNuPwHgUD3T/9n8k1Ij0AUkQ0YW
qPrq0I8t+Gn56pTCzZst/fk0Bs1csVdiADINmnQq5rIyfoLVrCofKHIpO68FXN8o
xHn8t3l19cr+SnqPV2OwgWPDg5fxxguwqxAbdaYt6PDsnI8HF4XxC8L4vos2JJg8
+JwwqA26bVjuYUzK0l1Z6lNVTWIqzeL+Q1mPNFg0ZXQLkS1t6ZqDfVByM1aM4RBx
XoYqf68SSi4iNmFSxeY+J3b504vv5HF1K1CXguFLEFZTJQtexewjA1M55bAsJus2
thXO+eseyCb4938S8yqhSaeuiEA86T/Q+wgynoiK3T6M6lyfDGbCELyoflTVVK/x
bmdqpzI694JKgViVv46TqzecRkstbw6cMpDVGk/8RtqAxlBzI5v6Vdvtnel58t7D
MyAvYlnXaaDVRzR5tYlnhDEjMdnZQ2gNHbV5mO33Z6DZY76aIYNOQvXssfx6ldC0
b0ZLTmO5m20vo2Oy/39Ajtx++8YEilXRbGj/OFNoPpTg2cnt7gBjH455WX+Ne3cX
2pWg9vfryl17B816B7QhblWgOu8qhWWvHYI3n9ztpj0nWXWluAsYAlRF9strF4cz
mu5uaCcY3SalCqAAA/V+sUWzlxWLVB2C9SpYOp3xr/EN51qwdGLIbnyhi/K/po8W
nd92zwfXe28YzypM9fvU1j4XGLtYzuj13yJhT8Stn8JqzSM1ZSATrxkqjdvXDOga
JLPtXAJuLYBAh9CcC1aaaUu1bCVlALv4xR0B9hJ0En6yeXVYqaipikyB1SDzkFbY
FeqY7wDImbjbOvMPRJ+ZFfrlUoU70GAk4OWU6zt7ZBLU9gVH6I03jFzTYgyVjK9T
Ly7eUXCYHH5vaBiMFVU2cDEeyd2toNqpVBrl57e+pGKTKq3xfqpVflNT2Ofz6rEJ
XWOmyPWDSHcLEA/OUd6e/Ur/79RLzP+74y0Ai4p5U1fEvqwLYYDHc+lalKf8Nmb+
0X6bCNNgy9Evk29aOP/CR4xKNmJu6/LmiYcgDxn/sLkcjc4AdAaAeUvOQpde6PsL
8TcmNYj5NLoIqDSAqfcYYzEXi0taleZ3kpHxdo7jh8F4AJnFuZUDB5Va/duB9Q8j
80V4nB9YOWJMlNDRCCfwNyVeC+s57Sz+tCeylFnglrIZLWvxAicUfsLAKbki3DH6
MCbPZ0JjSfBUvUHG0AVJlVZXzfDKV1BhpqddlGijicYnMbGwVZMwa5Wr2+5yNaZc
o+jSV9d7K4UGNGD8lhUODGcWKfUAslbWNzw5vMSGu7FgJDAJ9SZWuMpIjI+ChUJC
l7igKAjL6epOJdoscZQw4lY0TekgU9wW4Fht5kv3V4NYAMNHg6oR7Dak95ADTTs9
AAnN91rMS1pyfCPIncme5AuhF4AyC6Dd8jAqJf/AMSyFc468EA6zEZfxIgD1yyH4
0V3ajbBp8G1f1kl8ur7ybXgnZKV549qUcXCNlm48wi1A9JhRD9NeXqt0o1wBRPoC
NGxWGFz2+5g8RRu2FKqiIjDsYVRLv+IyzJOEzAUHndqzUWf1AVVOqqVMlue+00cJ
H2wzIg3x3lmsbS9LmL3u0dRvn9c2uQrCP7w6hMxld9qAiYiUETKpaYmbZEXR8pe6
tHXCL0579pIjlg7eeB6Jn6YTkPrc7rzshJ9DfojTL+v+Bj7q17POkBZdr/XfC0cm
Q515lvz+LDc6+v0i17ISQF7TFKmjY1hlFvmZkH6N9Xnjh+NzInQrJyAeg2KAwbGj
j+o2bWJ+fx36nAbvU9frGrtLAOA0XKSKeBdSbE53tcfqgxLOvzpMmyOv0mOXHgej
HwUlgM0uqEh3sVYuJ6pcFbwJThUjdnqfVwN3qtflSqpJN7m32UAKJwxypoDFpK3G
Rbt0dg5+3ILc8hefwD3ZpuNw7ryrfsmiv4iz+LpKOe8Pwn7dTbtfd3u8QjH4IJ+k
7/rqqs4WhKNcSyPA3hSxo2zxP2MjEk5a13w/YrNS8uEJ4KG//FW3bHPr4XAWCGDT
ca/9REvOvs8NLWKZ25inWFWc2x3fUQUUML5npaD8g22Fkc0I1UrJAmpftlD1hCxb
D8/cjoV8/RJpppFbCsqTi25r/xd+5NRxxrbshYMCpA5ldLNqXXEfH6Co3MkEhZhH
i+ELyhQLgZjQNqL9IW3pih2lwUaEsusrJWQm0F/obVokchjUjyELbFBaqGPIXZEy
MufvpnSzDfhCzxV1lrM7EfpXjOfoUiSqA6efkOSjNebqqFX41BKqlKMwLYqgUwlx
q9kXBCh8Pdk0FktEvHH5iSCc5XRon7mG3RxNl5TL/38JccXz/3yBW2Ctskq2yB/M
puYLLcUyEX0XO0L965nAE9wJwJy8la6HFL7EL5muQm3OoCKcAsFjlx3de6hjrv6F
eC5Vvf5aat+zybJ+dKeRi86thvJxo1DB9wlRKgxQS710sfU4e5N9XkkRfXgBjCHc
j4sO0sBXtjg3jPKMNtx0dpJDhojoIjqyA1IeOnKqSo8+9hFnjC+muAKuMvzAh94R
IW8qAufQga3pWcUyctuLi8uHdmY0lP/CrnAPRNWfi5kVjbUp8aZclhF5ZpBz+Wx8
IVvqAId2N6hNlWT+llRwyJaHbB4KLAYweNo0PaJruU9advRjzUi9ulIPrrZTuyuN
PoLjufdxFyZrzTg80LXnBfPtv1wISqj8SNHYX/ZfQ1MdbzugTp34yAZnc3dbaqW6
58qCJcLVLmT/BhJshyBQStMA5590Q8JlPztKg/4AgUe3i5CL9LAYQ0qzE5xGuOcz
PP/O9Gnpxkzf4NG59ioGuzSNHpqfSaNd+AcOXaqhu7cOxUb7u9hfXcS0QUxs65Oj
3oeeej12f1gimeSdah73Xl8pAX3Q1acRsm8Z1FgVnkZFNsfdMlDaDlynCzHFjrvl
QyB3z3cR/M9MeKaNbmAZlAR5FVO/DQznnZ5IxtzuQ4CPrn4Yt1pdxDR+8tK7Yt65
Qt5mJFMuoFkaZgjXzzHFqIC++MnW4CShqJA9UU8wGyBJbAUxzOJkMJwfXz5DSYdw
PgkUg8pK4sZCdt6Y7ECBgZscQZ+ivxDBygZDwzbh2JlCcSPqanENbsf29LS2I8Or
tkJsShZOXslFiR5cRvSej43TozPrGtK33MHcBlrtq7Uo+GmZMsii6zq4bALdFVuR
xuoPWnfzAnZmGmjmWJW5rIY0BkS5S83ok4yxE9HYBDnHun3jEOKr1uCI5yCAoNZT
g3dVI/ANsYjanL4+Uc26IK+PHHCGNxQzm8OnwZS1NGa3UsV++eziudZL2vwnisJK
I9PtZltYhfcpfr0gtyryC+Tu/EXGD3YKv/D35qKubFRda22BrB32Wu/BUsiUySLD
bdYNk2vX4EUYGnUtk1wkncf2uMXZHzJM29R5FTTnnbs14v9E80r/2VuAtxp0vmqx
vILE4Fy4m56ovvGArq29+e5UBvoiMJcWOeb70Y01sF1H4XX/4h+dDb7di0dQ17Se
fATg109tLBGRVjd0KbIMjl6kqA5LzIi03sOaQMLpQaOnoarHJh5cF63B3I5tWBUu
/3tdsugFqutxxdRHZlZ1NewTXMeBpNTTS2R1R5+Gn+HteQ2/YxGwMFsHbtVtBL/G
fOfIVThKBdw+NPoOJV96UsNmHiVqKEaH3OHm/d3XCg+p2af9D0iiKmGFHqLHc/yR
GzfcORpk23pNsF2Vj1U+OMfuWNyau7is1zrUn+HsqsH29HfLvq5PSM+2V96v1RA7
rDjOWtHeq2lGyV27ODPlU/pKV6PTsapW5D/pKACH+4H7uxVHgHacV6V0h4wpbqNx
cyzUH1+iFJmAwGqGy5xR3L6CyoXbGDEjud+uXwwAM9oIph/9E5Leb8QRbgn9UaDz
60q7QBq4On/FFDsYw3i5vK5dWMz5bD/yjZdDJwlHUM7jh/jpMxXydizP/bz8aBx3
3SUoCTyvcbldPHKxJJ3fDx6/5b6LRqowInlY1K4XPuxtAmonWqD8RlwHYkDiasdK
gSRaHzqYxKLB6xyrBPfXbMZO5LPCA0jFACwMCGFfkvC5McG+6aclRQg/FoIjtipW
e38BS3NHPXaYdzIQgWFgnu7Ej0o2WHV5WXqSdwbnQZorB8165/QM5CjmMQ7goD6I
61sYJmIbxVpIet1iOAfyhHRtxUi8z3oWA/Ao/wgGVK6+XTGL33zyAIRK2mqymg2Y
rK+gxIfXphrHVqZ9CWEQ4eiTK9fzH8tuSp398Wl6SqRU0GGNCbrSMbVENmWjFf9v
zC7ENL6F73YblL3+lVNb4YvY2mqMMXISvtQZaGCxVC28aobuL5Ia29g0W3TVP1yP
YW5awrt40hNY9J9l9kzDe5purP392AKywD9jsV27dgMrL+pUEEuh1dHzSELBLjbb
GeGb9MTIjX+VOndu8CE5CcL6mMF4cOTKuFtM5OS8HmIUu8PAlc/qggMtMT9gccF4
qk0/ie4PnU7stvBCn8LVl9ZmfbYGbjWhgjhbMCrUUwZkgt0rSb71L4uEgv6j1mEm
40IejP2JGTU8LlUnZAcz58AL/tzrrW/Sl5szR1dTbRrhim/9dwlm03eV9HtXx/it
WouVpTuDMO357RWQ5WJhEXEhJa0bOSXQrs3Xj1jUZ3No12uLabYE2MxvMsETLKX7
8IZ7m1U0iXRAhxNmZj3e0ttaW2x0/tQNWDVd+Xi82526WdnwggTDh++FxwBZZbVL
aRgLH7WJ0W1pEr01qj340BRHYs0hY75qXRLCAwmVdDRfy21TrNgnz0MQz3GMFCVE
gTdQkLI8B3SdfoN65XXGbax7o+lLQ3FL7OMb6x2xEPK7fFpF0JmP6TUiE1PPWT/9
8IS2f906vOwFQXtKJME/DpES7sQhlefp8qkeHQiVtIJgnA2D5x5jXVgYtsFEVOQ0
TdhqPCbAQ0npD6DZPJMwyNnp4IkdP6WPgTSWw6blBq1gnsWz7Ywnzi99FiDuIzeI
5HFWP9diOyYWENfdmuBNE8Bold2CfEkqVCfp0kIsgIoKG8fHszIOg+8V6u0yhwlD
UNeXEmlC9Z3xNnLnR9NOHbRnVEPewk95dmGgMxCRbKO2igfTsOhUG+FWffyPU+KU
T1h8NkaM56eIHygw0YVuZmb4RQMijSombMW4maTI6qwNnHvU3urxtUNbZYisOsmd
p8JBSL8IR+wZqwlA64Q+X2Oz/Egg6Z/4jnWLVRnuCKTNQPtw45PHZMZi8E/c23Pd
xcFd7Pb9DaKe3OjZMbq0oiMwsnfkIcLHphV3ONvgA1DF5dyiVSx5KUBaNbOq2pE6
wi15K1+uk50AQBb08v5Uqfx3aE7EmnlWCO8jYEoCYe/0QXifclSGwir4mcZHouNx
C4Y8E8UZNZLIFgugIyFLbeJXFfJflRyLSpaBQNaDNg4UmSAQOOKatDi7UnvrxrVU
vgV9bYLY70svQXDPc3+lPfmQ6NYDNNaTEWUVaDXJULLgujdNbX2dmiHPPnt3I8fr
Cvbnsi3cL21FSnYQ03pbC0XOWmsnwkf5uXM5Cl+hl+wunt4kMsy5AJzTTANSI1/J
5gIjXcA5krEftqVXWGjB94oc0Cvo+udsKj/9WMp1O0VEwVoTt+3EP4frc9zwoCvy
q2nB3KD36Q3iICFGz8se41EzZz1dkkF9VDHAM+ngghtyst717413dTapdJKght3e
68jnwripCnauVtjy1AKlncjmHyG2TWZd9k/qQ3k1ITNDggpaHywMlv9HgxwfOJYQ
AmVYuk9Wx/UoDIvQhV7fNmnfYeqW44cLbXBlJmRibJF/uCTUQojTHpI1q6jrZIU7
tVtApG7P9O9ETz39sSiOWTxLytq8t4gE4Qb0Q5uNoPhExqFMrOH2btb2fdWE4yuc
2RtrTP9cDlxaL+WXPDNLJbY3EPsTz3zKbgM2SJ7d1f2JMQ+yJc4/jstUk0kxWDE9
s+qMMjZxo+l+d0NPz5kzwnd7Eyni223nhhks+F6dFOIlzXD8OUB7E5+OUYTDEX8U
3UiKGqBGmNClFKDPMsC6R/E6HTsnSFGR035ORjT16n7I/F1kcxNB9ZJH2qN9Tkxa
7YHPvAYFXheBvCoWKs4EE8BCKjzxjhd6gBFaQW92q7BkEgxNq02W7Shw/dZXy0X6
KXYiL3E4nMdVonmvom0WAub24rlQXqP1SaEXETX/u9bnPpaSTKAvAzdhrCVCEIM5
AtfqlC7kmj0LaiR/+Ag9peoUX7DABL2Jb3VWb45lkoQ5rfVqdQRae55/IM3wbo3U
N3nUuyGQAmQbDStvNxoGWfbs7VXibnUgYM8xREOJ1jRuwPTOWyRfeFqU6G6l1BFm
G1N0f7HuNSo7zXcIQ9oqEA0PInGnGMDAoN306JqDIZ7v5BZnJpILDUX+1rilf9xz
7c5WzvaupGK1cfmk/Tsb2f3t2ls0O/EJ+aS2LA64D/uhuvPjjXoU7lnw6lzJ+pYJ
yOXLUUKUenCw/yGmgSMTXgi9VRU0OD30ugrxAB58kdrFUiDeLRXvgvdthv4CoBBf
rK9L/ncu398mihRAr+6nGwrmvuWfrm9C+K1tJa1+6QntA13dok95GVhlvwwyoVGg
Nt/s6TtCQmCOQNwJ8+k6SZmhQl48DXeC8JUdpOWEKW8Z/Hhz1eweTKQs4oqcuf3q
0d6hSRc2bjoh1LazB83TJippkCHfOgN5gDYgLuhdUJGuWryZwGboypfmvh5hDzq3
puWIQ/ozfd6WZBwFjHovU0FZs5scPQF9DFC/D/QVOISe/UrSX6P/k5TwH/2qIQue
vsyC2t2HUpiRSg9YbjZ02vEeECx6V5k7fYhGLIbjIJeNWQEyJbjqKuLd9twGqJOa
TrhUQuwofyw+Q3x01CDzcE/KDogZvH6p1Dl+kFyZRwQkLH215L70cPsFwdYM0/rh
mj0ptsFqqF+MS54g6x/kBDduvhpEeg1GM1A2UBQ9WM+pRq7nNaXzQ/qzKvixVomH
orq5x4/qLOjnmRDMTbanbxHTcW8NDC/0RYKIZcqi0Pw61cBgSTrqchtglB7sj2oe
FzzN5cXNd5a/73LrYZvDbl53devNqTkfvEzrdt+kmWUPpa/DxYnVaMRASggi7T1M
b38K6mDClpYwvglvNU1JuSu/e1XoDEZrXZKM+sfxatA85brd79QPMjn6uOTCJN8G
Hr87Y601GFdArcpWDKmPqQBESY99XWSIBjDmSISrV1oyI6WBi/bLaxeH22xrWSTh
ha39+4R5q7l9eK0EcPHbIjuvUj4Vr3HXPHXgRw+HKyMI7f/bfeVxoPzoUfbdi8b+
jFW+lU1jkRlDuXqZgKg21IJZDmG4JouAiVCclaYRZvI5WUEeGjRsNkMxS56dauU6
YNFXdvlysz2qeJlgmJQsf30jk2VmDMnbd3+OnJss65h0W0OWWw8GWtUKL7Uzhtkg
gwvgHaKoSLUsYuSyDU28bCUyBVX6n0xuYGNehq2GoT1unoAnViCvZ5iDiSgRH6IG
lgFH55ynVt4IqLAYly8Ys/huoLHRLF90pL+Fz+78FBWSxadxaCerk9j5e1KxEHmL
P80dyHeTaPbDmsORi5ptaAK23LoF+i9JZ7ZNGLgH8wbnkNxM+eMdjpmtLi3nNme6
iLSI0cSc8SpZeBFs9fqNHZzFFs0KlD1Tsyemwb9qs1muujELn6uMuS6lFkWSf5iw
hj5NLzrYCCfspXMAekL8jTS1ZRp73N+49O8vNj5ch+RjtQDGpNbv2r3jsrKwwEp9
QrGXsWIdkiN+oy1/uAte2ScPwiemPxOQmXSKjRvPh0sNZLfMiydT6digCeqTNf40
+olAqa75XK9AohnnuCQTmUAbcXydpDC9eKNmTmaed5OcTzr3lIFtHt5GEYErHfQ+
bCZi2BpkEFOxcr31hQa/t4pvxX1BcEGErbXQdnRRw1+CZUPl3os8H0aVW6ci8qYr
YEkf+fwbj+bPmFNCgVmRuRGPbbPH2zXkry+mVlyrsX7r1428NtuXZGqOiHltFWGy
EJFI+KnBdyriwRVwkGX2mxZDZux9NUo6OPrWv0KoMbwZIcbzKItIEOSFRs/TB3/y
NIJemVXhC2AKtIOuJAfiHqCF+prSkot451aApGpr3sE2NucgEbagY7w5Z1cuGiu5
BLjyCVMrxP3DXb3s1/gFCvTiEDg5Ue4p6AOEunJqcESe0ggDgh13V0TWDHnEveaF
iRdXdJq7PleU4uyVrY1qGpObYZdZg7TxAOw6SVYHXtHOaRxGXsy7OGrFSs1FFeJC
/zr/JtKMp6gQ74anCbeVXhYCqxXQOK9VBs1jDmE6NawL2G0S9aza8GWdmzhKjTuc
svQf88gMvGrVJs3+OOrdCaIZ/cjPq501wDqx5OqVKAxPUEpEHGjPBhQhJLZy8fod
huP4F171nsTeBw/qnPfwy8M8h4NINt1XTytR5YxqB8SBN75vy2ZDNE1oW8SK2veA
wk0FmGE5pYFz5+REF4fITVcQB7V8rSrI0ugAeITJ6Ka800ervnABSIniqU8LMrHD
KGMZGc7+c+OAugXUZhk2U3n30nbm8fvqgnXGugTiUBA2CxIN2JRRGM6GrHs1R5CL
3/FHbXzNlkNSc01aGzxJbbaHvp66VgjyAmkv887Rw9XnB1uYq9+hfNsPctNAQjuI
w566cQlBP09mK/pxxRIg/IL5N2pyTY1JliZCwpggizVIymX2wHVB0XRvrJXRVIGK
ArlU7ChOOItcfSUB+coPtnic5IGbY1Wae+I8EgPzeuOm7Puh/2nBAR8ApOGJ++nx
MpkKzjYujTQNVXEz65JwPTTtCU825LJTKRPjAlRG3lAqMkHyLcmfiJnQUxV/sd8w
7Sl6Q6h+fMwQGNBVBx7AtwVRNrQLIWbrYdkmKjtXOOJgz8lgzt0yOU+iDrT3p5Q5
scWzxTeTuQBhqjR5LI6VK77vs3+HUznPzZQmvc/ulelAnZNO+YMKw7SGvTUrZD+r
y5O0+0FOo547iRlUtz8cjPjz711N1S7END+PvQAQCPD0E2njtUY7WIFzOYpxlzxk
PT3o+ayWbVFycG7J9Teugkogvdy9Qe/NCBJtzMWJCgzEnqpz/qD4rtg/oQE2lETs
37rx//KmyxyKoEYKIp4hpJXESwf1I+8Yg5afSy6YOD7hlZ7edE5caZMeXRV5bV3/
AsSpLkpzNd2ve/39RZb/RkRow2+DZ8MUPB49HGEMULE=
`protect end_protected