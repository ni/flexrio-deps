`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 232064 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
ShlXMv2GF102AsumIDG8qdAicolugbH4AoTe0nH595/VIw0XpYs1d8/Qd+BWB76q
YQrYMj1BjX7Uzbdwmt69hJuZnvRWH6/JPdMnaXfByxdlvXfEW/vDONCQHss0CQ8J
WbRElVbhMSVnGnCuf2dklIqlYBgJ6GUWKSyipJ4LdlGO2z3Ag2TphQQHDwTWzHg4
eAy9eM1o7ExjT6zC+apj6nvHkwWCkoq2bOpkDTLOXbJbIUOFQKGmSR69jhAqjQRt
WSxMctSXHLXe56LtNq59acd0vEGmhzip1nYwCWnkWz0a7B+C6Zcipx51xP5niKxm
PKENW2V1PeR2WVr5wAzDlMsrhfBN/69aG3bmdfyF9wmi4B1jFaoHriGxUu4qdR0S
RmQVBonYZBMdz85gsZWNm47kV5RIxnBYs4OBdrS+K4JwEkEZl4TqyhVNaWQ07ELW
wXBhaHz2plZ8Y/XrlAiL1D3ttltltQ7riFuBTDg7p2CINMF1l0r8VgROC2Tbvajz
zGo6KdWLAP4PP4ROegJryTSE7iEI/VfvcOUzwqAaq/dK+KYxcYCP61Y5JRGM4boz
1++gyp453tQr8KPk95Mk5NmxCy8h79jyHuW4mnaNZOVe9M2kehp0525ycMBteBoA
xXJHUV4lcLDKw5yC+QeKJt3ITW2ddWAwQ9xgtJTo3+jw3Sqye032PBNyGtL9XF/T
/DQ6XAugHuCRwbceT+GqfB8ZZwnA7JxECgMz2ZztZC7CkSngbY/Ot7vcX5VlYr9f
vv8H2KnY1Sju7hKVtO2frbvOPaycuav5rO2drfhl4ddaHab2Xmx13H4yiL5tfmvJ
mWuEOUWa+VDnURFhWAzcQgAlNMk+Qr69QLeoYdEyK3XgAVZVQBcNYQn4LloQ4VjM
mDQwExNZwc9QVEqQk5CJ8ql8KkoR5G6+YWJViwQQzPg/7090lh6v+ZbMGjJ8Mfs2
iLpi6JK7t2j9KLHgcaK/YYOjH1tm4/LoslcmvoYYHC5Ln4y5qYse+6d28nLkM2j8
BCQ+MoTEvn6RU/SJL9i1LBc5COuPCouE+9p8i7xa+3hDj2j6FLe53o38faO2/Sy1
lj68XnOsn3S8vewgKOb11S9uvhsCI90rC/tZk3xxUesDNemE12q8eKGgNtqsr0QH
i3T8+luarBMyUW/FOT1dLRuwJuomsemzxDuQKdcxNLJSnW6KY5ThWFZLl+znA69H
J7gg/hl8QLDzYlEL7dYHRYDGTh+PekNocCfykophYw6mLn0kaQfZ+qvH7JMW1kvT
GjCfWJvptv6vYpa0uuwtEaNTtqBJ52roH0Wsi4u8Y1IinBpQOXRilj7IK744Vco/
rXDkcNRXXszMOcQqis0g3kahse41b3gCX9O3pXKbyEF3zie5HcqyTlpNtuskkgh/
Bnh6bAZck8XzRYJ3skZp1FokbqBq0ydb5ImZW9PUXKajPWKni4JkwYynGYLDkOqA
rQ6egPGJ0u1pnNiZuW4BP5s/q/U7lXCEXZTscOh8j4cz30LDKCITPtIhSXby0cS0
EELymv/ZH6XetnanEF9bpJnWuKbEhpzVFALZA9NiJQzycGc/Jnbv9Hz449M7geuD
xz5LFRA+YERKk4u9KecMSiXNOT5vxAAc4olEyCozkNx6iAb09heVpHoyG2H58o0T
LK0RWAdBZybzX6viZPqS94oWpyq3Cfl3SMJodexEyuNi7w9/1n6DvRs+tocm1t9p
oB9RGfHNw8MLp5LKHBMwnrogJHbBckhkv7mtW9qOHw4CuPhNMCTRmfJiyW1TfV1T
o1qfrZyIZn72OssaqshWzEeyWCtCy8LUk5cUSkUOIw2Quc3NlcsvYULBaaviTSYl
8SNyfceK94RmsKAFPipr19o02lohTcLeptH0UFJpdsfZaQpnyMHnR/mggOpZYgaD
3Auvy1rvkLgjXzXFhgilb22R1lT8wT4jLG1NvVyUMULZhT/jHWgYv2uNvBpRe5kZ
Vz4dHlGMh1A8XPQ9gK485nUTRcUGl/qCMayPo2imUcyRIdBxUU675DfC1UsraG25
OcS5vk6IEBRSoewktbjasfYpKUKeQhHenvzfYOiGs+OB7zgTUzWnvFr595muB6aj
p0ThUGPSV169/1bJZVpd5r8gkvX7nCgsl2/28HP4/w9e+j2pk79U3lmJj2OQ2s/U
Yjcic/D6bb33GtTYvlHsAw5QNESW7EdChYvPpJu7ZuH10wuk3denCJ4X1PNpg8p/
zHZF9iKs2OzuUp8HVcMpX1lvZlbZsgj7Rh50W3V2IMDHosh6mefPzq8lUNTXdFsb
FWVQcmZltMjroqh+zC+1pSbXjCko2vHN64OOly7YST7b2dJ32DDAw28T7UD7C96U
ry2yThjkmeJcugeh8ZFRpjjGQ/ehyLe9Lc5wZ0nYFbmBZp8Vj82JaviIXgmD6xzM
Z5X7l74tQ+SKsAtSu+oQpdsgsOf4yur5VgsS1qGPgJuDD5dZ+mlLEPy0g7ouTAPm
d19I9HYu5FY8UM+q0TayTzDeWzRN00NT6Rg8MGqMl+aVfID7bjUuNGM1741uzUe5
JXMn8zv0G1ZrlOvOCBb8n61oM8TTLP7uhbLBg99GHnwAqWumJCwDupFyKApqqcA4
dMIKK+hLynGugrAfqI5BJAG9MnIx83XqZbCIs66DndsnWrmizYgWJqSN0gcbqfJc
OjfKmVkNAprMrpiZpdyXuEPXvuPXl5PAeOwrccWesWzholWoIdHUcQ2zteY5E5B8
yr0rit/wKGfr1Q09wRylGHxr5HNHTdFYmD1S5i1O6L6C0I48C0gJi8ScpMSfAYGp
txV5hO/L/K6K0VlfC2HcxuCTQEo+eS4moHEZIdmN+N1S5KlZIQqHO0Hj5Rcji42W
uXhHbq2mJrj1CSayB2An4ksM97IrsfIRVEF17t+FfjAKI+WMZFNtUTD2/WQU/LpY
1VMRnQXn4krisWZKCQIF426YvO6JsI3zYETP1XTCh6bXl7Z98rZx/CgBRibThFlV
tUh1O7+8JO1xnp71k1P1XtpBg+X8aWeFC47CU9OyM82nX5fv+JNHwRU9MNOqWgG5
jPLU8ubIpSUqUHNYs0xA/9jrF7LFgsaTlw70HfBKnffd8DG8rk8KBD9Dg25WcwMV
obeJVZMxETlloK/19TsKZpa8e6BaY4GwYbJLetKjbQVsvCBDDiaxrBaxcD/sOPNq
K8Egyf3/k2BFp1QRLNl2C7vc8cbIteK71jO3b2Vat7kVRFjnaikjbqtGEgtHnusm
42Ind0pY6+0TnwqngbWePouXqUXXc7V7iziSHTnC+n6GeeI4GifZ0CpJ9URPNF1L
0nEuHLE7zbTkCPO+JOMRsqM/gnBaop1mLqDp0xv8lSXAzRfQwZwUjT4V/WGe3lFJ
TYLV4l8HpIelAgtX9dFt1RXSWsbXUoAitYfbGRhtr7kEWxLHk0XBUU9xm+uvqWrw
lcqERTSPh/C16Tfd5R0AzENr232oh3IlW7HODXsXRFmdcn+0w+aQDPvpvR+LU2Tk
AuQeGDdBRbH4pDF6tzmTOkJ2Sfg4ZsW+GQWo5Z1rdEh6dOUlo3du8sQjbt3Ced3u
WbBMuOWf7CdIvWZ+HYAd5rrazTiQOm7bUi1MKawJqIkh9w0YKHutGRr9IThss73J
Jli3nBimmeOt9mBQmEu/MU4i2Jkfl3//pEy6pe8cRavp5NuwJw23MJfBNB3goEuy
90bOX7ytmjne+Ku2uN/2bir8pV+33Yf+xPCqm0/uVExCC5866BwRIpgeAWenXrPq
PIQqUUx/xwxTX7pPTv2xdNLUi93TzGFSX60O3waXBhyCu0EzfYhJRrgs6Hf1zEET
Lh6yedRYflhuFffjHo5jdQSMvSFSGk7I+kVaSRQ42vk1azR4pJQmSsSUjVi1FjcG
fwX9fMZT2k/vT0Kte8/MR+zzA/qpl81A6tp9UFMZQQ0wy/m2mzxWrwvtrRw/+7Ao
UolM2xnv4r/A0YDX47sp9fCb4MqgpEUzBcgrNy9zrk4qWQKZE+tOwKuzEsiw2Ieg
NrGorxHk3sV0a9vn/Px8uKZw7p4QK5A34c9Qv6XKxBO8TqSI8/i11wu7YAWleJND
APxr+gaur2nXhczfMc3CjUNJ3cpGT+LfDas9glHyv3+S1y+nSSo41cq8Rm0wkdE+
4InN2yhlQ4tUmkV6tiIihUMT3jhyE2yLTxrGQfBud3/ogt9mh3BzZJ5s7ACFzJ6G
/QP4UxnYdvS6k0blyB/8FqZxFHZUA46B/rKC2QeQd2y8xJpCNVV9SY75RVog+Vv5
0af9Ly/fFtteTC48EvfDMsmBlORkqosoE6Ndt1ajkmRfFipcjHFYM5552zJBx+FU
Pq+K192RcCgwaPP8dVs/OF6oU9HYmCl8k/buNm7Z1P4sPEw2tiue4K2pPvzevcta
DAhdSLOtK3pp9TmNJbQ2J+3nIh/Iv+T3tGij80c+whzH1aI7n/ZIXGx41ODp7W+N
80miM+YpwhmWHQo1JqnCe/K0MF8wP7mRdrt8kxEizdnhqTCKJJw6I4MWDV/1ZCUP
8tE16Dzo8Uo4muEpZJqRr8rftXy/Q10rNZvBYRc7EszFOdG/6MI3spgYjMx9tE1I
jpd0VQoot1b100KYj6vfkL2yO95LqElC8P+XkOTTXFXZtZ5SVS3As0zdto/Jiv+t
XJT62Dl46UW8M6dbtTcigpm1Doc5XVzSH9zLvojKyyUZ0skH1ST2WCTwX4Nn0Pce
3Ic/eIwTsYPWL4IIPghtaqpuvhJata1ZWZnygCQdy5iL8t17NWrpH51GANjuYTii
vOLDAsqjGsTU4ijOwofId0E1H1t8jWHwXH8RfM4Szerg9MHQY/FvtCcXFE0mhmG5
U+wP9Ulu33SkeZdTOunV7W4twO6GAiwK3qlbb1xnWJYyBHNqaaYtguMMXqUklyRr
ScpH+7wcOGim8Z3YHdy925vBE+xOTYD0P7FclQL8JW+OR3B+LuFUz8e418sZMfQ9
mZ7zF9BcFI6XtXnFhU3x1cWY5VFpEjtlFNijQ7tWsEa1PgcnvW3M3ld43+3MbetX
YJbBuRoA8IZDykrzijGCnJTa+E1cGEqEdo4TV8vu8IMI4vSCwECNYla7l6vIvj4s
ycfld/Azm0hB+gDWD/1al+aCCbE6/rmz0pqv/0W8ixYHzChoknH1HltOg/oY/bR+
aU6IcUzDOWek30KrsFikHRSAqEu/jNDfHwW2tXmHBPdWSgNJj8N2CFw8oCKYh1Ln
HrnF/wtoRCQe4NsE+jTNiJRVlAva9knBnW46gAuiGGFVu0BHaTnWSOWYN44ibHLp
swBj+nH22EUUbk801CwyxEA8eTrnwGxp0DhroO5/WWyV+9rJHJT4c9rny2CNUMw4
yfK/Le+enJ4CxvMsljKPXuuSz1gYVMNu6EhgfhFt/JkspuAX3ODcYaDycG+sps6F
7kL5bZDsn0pZLkhGYlLu2lzZc7H2+Pq/w3Iod/iuV2hCJ1p/YgSgW8rWlcTEfiee
XUXiPLcmKdBm0z9+3AjLVzQHss/3xRdc9XqgDmi+Xk78HoULWqthiyZilQ2nLKi6
UaZ+iNP/hgoieHkJp/GQQ8v476O24826wZ6JxVLdfNLFwLAd9kNUJYV24u8NA0H3
/TGvfEdIxORrhjKLUv5AVmxGvu0kK+q624OpHz0tROVGHwf3S7Q0gWwvruweOB68
BcQHuCXTcWAA5XYMghMNQVc3JvbKHSpdEH1HWNWJD7xZISolFaeyRlrG4dkYu7TN
WP+4Yzyf+Mv6Czm5+YPGHmQCQkggOY7onJZGYs3nSNNhxiHHKsk1HKOUpDpncwgn
RztFpe+MIfaBqAhLFlGXu1ZTsKcZIeIUQ75zv+amoRi8cWoLGJRB/vVSFf8ktReL
aHQJtQ3BE15xBx1eWMXtQyYp+gqcqSfzVUHHaMvyubA+mdPX/jBxamwXohMAogVj
r+0uuXFeA+vFmpurccI7UbniVxSByZiPhQvPmGWtMDS4LLtXnbdD0bCYOJt1VPyA
VzLj0AjQlT7YTgXteq8SQbbfOaVt5dcHQ6UHZvcHvaOmA/R37nllNtWdtyVn32qW
54cd6+UTl4Ono/uxK0JDx8OsVSD9YGBO4IKknHeF1Pf+q1EUJDb8l9Jo98WXp9Rs
TAGjC3iJxgmJdv3nVJr1CZ5xXwnUMrf+YM+d6j20ybDiNqx1qSe7naoXPh8ssE58
WnPQ4KCK6J7ZHpqXfpyeT3EGzdPkQHhJVF7hmGe9ygvM5xfHWYl765iv01ugvHBl
AWcu2ABU4MunizeKlK6Dp/niisqRhg1cdPnOQ1h2yIzct1jE3K8qojAPoAqG6xUE
P+l1yPHa2ykTlY0i5PohbvHDuIzCVAU7RTnOvpnpllGvTM6CNP4N45E/s9HJcvkX
CyfMEL/5TlfiezHWXSLtx6jfynnsYQpqnDY9GTvc1X4PKvg/pNnwQcfnvbmFX8+B
qugY6xoCz2BRffiDHmsnGnptvFhFAf5KX8h/K/cHUGBzkW9lhGH5O9hMxrmsgSmt
UBi+ctcr2U5PtHn7WPigE9aGIhzL4k0/g3yWv51T/fOAOlNW48WSGAwduCrLCn3R
lZuXGncioos8MImNz3yop0p1sRl97OxlG78VTT3AqYkAlJ552x89i/yk5w994J+t
CooEc4LjiiafM8ZQURGha3qx4e31TC3s4LRyLbFXjC6tUZBkQpsQ+2uhgiYx4zb3
FXK//1RfA/McrtXeBS0Zns3m+4rwkd+FAkkbY35Wij0bB2o3WnBBBd9RmCGdxIgr
aHoMzUQkyy4ht97yZzHP8fJqFsuYH/CFT6Oytx2DVvNFDbKugYcbhqBQADr8kGCC
+xQePzT13cZcKvFBpiU7voUu4iNlaUXTlr/qhgP+L2ZOK+u4TCLvSiMzJ3CMcBOW
lEvYFKtlufitE6vg5A72JIQT4EmEOEV6hH7ZmzGf+iXiDG3S0xlnD/JH2UDJLus0
bblokPTdNpbuceFuko9i7ZGgtreVDkA0O6jbDXpHbrlbvOmMM6L6GguyGfPX7qfI
Dxo4XGGfmCpAQYg1rlitAMvbquopQvUdUD1u3RiIB4eD4ySamo54cWTUUG7M30vX
EHqv8/dP4K+4R6vm+hk4trsRp1byNFWl2ftpNwNLd4gUPkiJUJxrklxxGgSULLRA
xFzLiPJ41B5x32TbWsfEG4sWt3hR9Ck1ZXR7YV5xb7Bc8BLbjGUW+S49lj24AzY5
127N3F+lq8G9Hyqqh9guqtbpPl9/HcPJR1cwdFu0mlcktfAs716MQLgnu3gGeNq7
RciS2p4fmwXdLwLe1fSCErotdnzgni4NKz6WV72of9ivMm3YNnGd4t0W4DkfLIhY
uGSzR+/9HJiN1MF9hV3OFsP2A9SskHHhARAmRVLUh7H3sSpdzR9ZMejDOXSWs4PU
CxKKxqFjz1cgLSb8+QecHQ9pyDQu9EShDql9njyKCN1KF6R6zA8EUKRHA65MKhQT
bHse5c0GHEaNJjMZcVM4Xvo5fxfgTrx4FFoZXAWQP0+mfoMtaeNHtV98b6xcrJKt
J3QmvGHvrPdnGdVrpADc95/haYpSqYAfdTTtj7eqTydIzQGDAXFJKNtt2ydYwPTx
VV6PNTGL+vJHSBbE3aYNREBW2yzRs9VGCsfbKNXkCNSlhqXaZCwLq06PL6wLcPd3
KqsAV9OgHVkyk4ckqHShNSnOcV9QNdMz3mSqO0aUwtGSmVr80VsaZMmmObw94afc
TXvUE+t6Q+2UuKxpZZ5XnnxXB6jIF+pltmO+ixr6uFCyBOBdVIQb4SsPaMWZXioo
FsuOAOuB0YdwtZeNgLJQ7uLNE+h132g4eve0ZUACstDAffFTSqyjjEz/kDqBuU09
XIMYNZxUulgOLnlR8coRsM0IxL9QKT4jGDa/XqGpFSHNrZ9YpffFkjg7DLEmDdzJ
6I2Y407HY7Vi3zKuNO3mvKVG40zvVt/TQUStdSDKol0aCYDRySwW1TLVmBc4pOdq
fxkBdi8DdjG5Y2x7wWRILprBux43nVfggHdWIhDb1dokCOWs5d6omlL4tQg42IHP
KWgx8MvukCkjP7VKJgKH/d0KLNeqeFWHYzb+m0bbhiWOatnm0HeEfCoDbeNgrNaP
z40Bf4co/+FCgl5g/kwvmw0F9RryO0jH+VwCJ3rT8Z2157Q89Dd0afhA4ptSA55w
CwDoDlX++V3zwBQipWZd+ZOHHtXpUa5/i6rlFRf9ZOUXj+SIhOtU6/JbmZ26JJHq
IHUD6drN6o+kB/4beBuYudyrk3oqBfvFo+MEkYnYuHJT46FlCPzOeCW3pqnX4hNA
GLGRDaZykgv4M2yM+vN7zebNXIUHsqnjJc5oV4M00NtDqL2hoTKKNNuBDO9r3F37
1miF9KgGNU8M9FQvXadd2xN5jZGkbjiTe29+tW6bA812ZnlnoA8HmYg1wrVsFxfO
PR5DYuyhkSVcpJSIuA+SoaVarryWWve36qcCF3+l/aEdB/q4/WK+86XLA89rcyMN
vCAttbmtAN5ONJC7deyMKGeF2iUIBUWElbzrR/9/Vxxh0FZEIQIeSpH9o9P9Lx0D
S4seNDZFRkQnv9NK43Xk970CHq3fjTt+AOfoo7yFD5tW4o0dwoXimZV10S2Er8Tj
DohKl2UyP6sJOmRCL4bCJ69HsHUWnNPoGRRK+5Bw86zX91Rots+Tb/ftqVtxoOOh
KktJUveVx9dFVFOZiNdBEkVZ22vdN6S0Yz1Ucvja2XkqzBRHuJG5SgzOHMNTMB3j
Onn/1BCyU+uG871dqccECo3VMzu/GmGDC//mfDBoXc4K1SKNFHv636tzrGJ4J27x
RHm0Hxn1XW5unP06rbvM3+Fh6Yfy24zR/FtXy7xmiXdHsA7RdNnSNTdC+6mxbCcc
/IT54/G/sS2m+V9+CkL9XV9mYO8c0bmR0HtSx4OQu2gjTF01ecD9deAHwLOncPZM
1Mxc0w8Bm75e5CLm79m1KccmmdBjfxwaYVwsBB77Ar37vyHs2SQZPj1b97/2quEd
9MkApmHCBV2aE2ivlp3L0zaFrtWn+aQ+qi6PMRP+t78MTOd4v/MB3FXA2/LOqSfB
tCDVTezHt8ChDIEsIe/dEzDZXLa7u2D/pHcx8jQN03+SZ2TRYTYjEueEIY7hdfic
szuUS8o0OO3XhXim0GUCxu85tnESpcUBSxEo/3nflgIWoBt2oVYXjUvh+QOvHboG
NTEZ281Z8ljiXscaAci6pZM5eUy4mRdNHQP1Vvbqjay+w4KiKqXLOgaUCEMNN9gN
kEB4Jm+TvW+tl3WxORlrBYnJ3VHxYx1FhTmv8hpnXkeu99ITD3VXLTZnLYMxfT2+
+PkduozwixvuJNZ9ZyHSy8uFawvAbepaF4QZCYvTP3MxlzIhYTMvyIQ28dQXhQxM
I7Uso9r7hIVyqzDCOgmL7D/z+0X0vq13vXpz4Qnvs0SAFxUcxpBMOmY3XfPMkw7k
PRHC44Idoyg3tl5rYOLVr61HG6VLxFxGRxvcxpJrmSLoBiUVItJuTvm+1m1M3Woe
DUPXn6xG664PMxn8C9ECyKqknkXVyJUCJNdv3OtdtglJJIuguyQQH62MzNdxiCo0
152qJpBqp1PlFoMbllTOlhPJvydpeELl6J/gEYQ77O38saWSfU5WxNPpeR+2n9AC
fRMlW4WHABLEZ6jABpeNXj7H+qtMhAb2z3cvFVWKlyr6miyTZpHsHxN4mUFPkjh/
4UhXqq79jHPna7KOOYQ7b7xLB47cwhiAguqv/7mHKIvzk9CWC+I321FZ3GAM/BlN
iZ3OSEUfGWulO9BHUj3yYmdl+dWY/vS3N6BWqenfCxmmjt8vput/SmT7haWPDIQ9
K82fGxh/Alyspt8KD/WWxJDyiX6YU8Kf8odd3oGGD5XqeF5XuBju1xsvfye/xOcB
H8HD9ScuuQwBLk1RssSff6tmSWt5PQ78d74GqhRsW+IhacOgtpshllHKd08SGdMt
iE1HERsXzeOlafCZVtuLjdxX1DbrSu4bO+1F6kWXKYL+M5cnjQGsrmZ60kz3KrQS
gbk3G7zMFi6ldFpYxjfvzbZIWAXryvHC4+pZsKRWbnuhDYWdPjvd1tTyZseaLPcR
5Rg3Fh+XqIf7M2VlafCv5YC8OmEhElvCWDWyY/I9XEdaah/8hQ1brCnLcYjdUEuu
Ycj3/reogajuvl5EnnIZrTGeUXT8xShBcvwIaxD9tR41l1P92j7rAOuB8YkreTxV
+gilRRMkor/00AWCVGZL+1L+NMn85LstUqipGt5kGNjn10vy+WIRExtP7ksYsljI
HcW+gIiUtp+2TATaHb27icpv+/ZP2JCo89JkzpIYS9xCyDrmN1g2GAh/tMdJCSqQ
ucEPtKqSt3819Ah7Ak5Wa5ud6i3dEqIctF7IsJKnhZz2C6k/KKbVxhxCVUkpO41W
bwWjvYQYcx3CdlVJRuPQnXhPS/1N7PChTuH7hj8JHJ85nkxThJ2m31nstwWjh13O
PLIaOTC1UdYVnEH5IsxrOckph7Y6ohtfYldcUHKXZWB5LfvDwJzFcNEmpFIDf1FM
/yXkhSKUxLrRyFzpclkMbKAZkVgPLp/9yPd1Z918p3+LbUEaOcQLSlvVswxer6P9
aslMlR6++reYFpf5Npwu8NztFkMloqxjCs3G+gmZbWDQaqRMV4xDyp/JwkEKwPWE
erIHHmhA8+cgiq3AjyFChIAs2OmZ0zzU1hgJu9RCvh3llErSXCELIl+5cLgfNoO5
uu/ZHdbt3UEYCTeGQQRmRpHHAPC9oDSjef3JYj3DDqwjG/MZ1WR5cNNVEftARWgs
T9xiwUQeaSoppm3zI4dQUUE5+YMagjKJUTSnj+HLBRjnKehYOxgcotAwlO39ke5H
n8Rr1XtFF1KIlJgwrvb9+Hrl4YMY9Is5nBd7j5Tmlbjw2VBoU0dcS088Kuk9u5md
E7N3Zg9pEPHwbKrXWBoBCdlnr5amgwI6rdckKagtd4FLENVUUDkQuNifbOIvPkvW
hoWtIxnt8L0Z628kwZC50Y4oNFODf9OeMobb30h9RAZmJkU+iQ5e6dzw8+NfB1Jh
2XzV5Ycj9QLgxfJK6XU4WFaWMVU78SZTAXl1GKizrbo3eEMoSxY+E2Yc70C1Ycxg
YFZr8lopdKACEzXPCvCLbvfGJUZ3u/3ZGOg67FPGWFH8W9mYOnKbNgG1A/q+gC6b
6yGLuuivkLVX6JfHoh25QV0pWhR1sxgI/os700qE41bSIB4yjN2xsa4JHn1LNasQ
hRuScXv7FbFrfEtyjk/5J8t6DU6Rfc4Flu8hLOdFksFbCxZsusYSrcFBKlgvNSVr
akcHLNxYxkIU1XoTK7BH+BQgEtLbOhpc0nCOeQjeL8maHJCpEoDKso3+IiuCUJIe
oWdqVr+XohMAHPpI/Gz2cJQk+WkLE+YaLfmb9njkNmGHG1vYvBoKYrIB31tXIUm+
rzdKG9mchtZl715SMgCrPoKhrl5lYpmi0HSMf+MN7/+2vnA5DsLVNHfoJSt2QWT4
z0iWPUPsyn2Cx0pdhnVN297CZHHMw7V4k6RsS2OZt/6uSINdyCwOehVfnWcry+Vh
67DsHHGeNqSDZm1nOf/QWGPX8MAyFtNVUIhxAg1VdbZNgQr7MWRSnlB2fqJPrHyz
s0iqibY6zv92/gJptLhOADj3itUsJ0mtnc87626tH+Cmld1TnjPN29xWEwsnsRCQ
xX9MQ6UbHEgfgB0CUaCEZ/SZyDSNyn6q9SRDF8P7TUH0loYeQ1Vnt28GjHVxNyQ/
Len1crhJEL3rVowp/NxXSmdpK45dDGgrT345Crzf8JOgQiND0w8mKAtsrUUYzIo7
bPIPuMZFE0MPgGPFXqZwT2MCPpk6Aib6HIXCV8NDhjGWHxhZmTJypSnQICfU8ut3
72BFJSKZC1uW0JuWGsMhrlvp/oaQ4hBqVdZPKp3U2WoqajjFV/5QZEEOilpHCmC/
BvhkROr0dJMEq1kvBOXEcCnwpx7fsy5Nn3GvZGaCD4RcDSeXiffJ+bxF7+1hsjZZ
Y3R1beFnF6nERIgVQODfTqYWEm7o7/aHPbdZjUQjlbWOlMybj4aDIESZIj5I1IAJ
icGfle8vm6i/ZFNuWPaoLvCka3otx+RWuepshjp1x0bPtwv0d/kkdWWy6HUoB0Fe
jcIih1dLzS+ZDxLkslMBjsLh4K3RlXmGKDm3tm2EQUqcl2BdU4y6ssnQ1Iy6R605
oymXncAMcxLiLzVOZd/mJKbd2xmk2xQvQYZKy6kQfBXH50hBalKBecsSZ02WRlYr
o741hNoDUCqKUOBHti3VSI4DQH6I1D6m5Xb460B/WeXwD3+/oax0PS28qe0fpndU
lzahFsqu3QtFYaCBC2oswJdj8CKKk+iHXl8To7XWwB2L3Zzwl4o9Jz6so4tLFE3k
gNKII2Ac4HxEHbSk7hYDyg4YVpB+8mnLVbb763Fpp+HRV6ahTLUeQZc9LSpZIIx7
eXrfSJI4ZyEwUmWafFWMhNoDuvTJlNRqfBeC0iyju+JULNaKZrtnfi2mQTh7g60q
jrChIhxqBVv/vYF8K0rEFG5puMmv0zmAjUkUg3l/b3bPAvpdpjId+VHe3jD8vjvi
3WnNO/usTk2eJBTPvTdO6g70he7RLyP6zbm+rBKVleGMqQ9NNhv88RgOaOUqsiTm
TPqyQf6NwjMMtn/36ZTfggGLa6zhoAA1HI1bQw6u6K7NEJNQCJxAQG0B+zMkuDCD
yp6FN3HR0wqkHRmCnfuO767yrrMCzfmvWgr0L9f3hDCScGKvkTvN4lX/2Y/SDkaS
pj+rzW2M3S+wrMVmxSLyjKkTwX4yAImIOTOfakGQ/7jaworCZKvuCYzFev8GDrcZ
R5yowej5Y480XOSORagviK6s1b/cTgW4WZs6kF7BWUbEQkqzEkWowakv4tR4zliM
2yYUCfVuLx5ZoDb7iKWa64dywQNs0otTXt38v4RAEOMDxfWjmEqSnPBwcJVDwRgL
Rhd/i1ErOjuc/iXc/RK+4MSdplPinshlSup81YmB7ROWaiv7FOPqoJPx4v8ri4Uk
yKCdlI1GmU4ptt60UcX2YzSpfJRZJV1//4cybEhXHpVwEX3P6tFqe7OYsu4hEbhg
WX72DXilZIm3oK9Cp4sjPOp/hmw3LTmYyE1Eo+lqUBNA+GapmE+T5TmhWppRjpAr
m0t6EcNnJYM4lp0d3Ev1q+GjUEhv+eDxDnDBjK15E/8Ba+yD3QuQszO7vnT+KBat
1kHKH6Wn+rBg45rI595mtAxUi1h/IndgVnr30KREQiPOsOfqD6rItUvfiQe1uNkP
BRhqqX9a56jm2cLsd/DzCNZq/6LaDuiUkqID1cFCPrkLo3CeEOvvUCgPOkhgNyCL
/OezPf95SIr9jUATb5ZXlCXel9QDPZQNzWI47nq0EOoryf9DpIAsvKMvGmtwwQnm
hCt74P7cc5aFr0zNANsmNnMgWNa8/PIo5K441o1vtCkCeYAoFqKMpZ+tHOuAJW7b
kzJwlewq/oYkEM4kZ4sKpuHDjPvZHVMwHdblphuNep1Ti87K9QxzYW7Dmwx/z9NP
BJ7g9GigsLZ89AJR1Yy0Da7HPMMAClwcXRiD3QJhgetEBLh4mJ5yZM0HUdHlxapb
dB0ofVAtW1aKcypNtBJWzOt9r9pU1i6/xjVQ0pT1cZUprJzONxSxS0wJ4V7l3Gi4
ulVUnekTRwphRB1FGb4T5VM8Z2+YeRCyrXwHvhopB1VNEDyXeEfB1MblG2mThj/7
mECcvOXIF5a4T8mymdzjATh6s7L28uOluvQ/4KzRdL3pJbSnmDU83igE3YVqO7Gj
3Ejz/SGVo0AEi3yco+rCFtk8zBFU5/7muKhuyS3QGQNp0pbntPIEtI7vujig59A/
UBTJECNUjzgvMNSImxZpymAi/ydgt2153WJgWodrn88HnOslJUMoj47/YE652dEF
3iCfrri/+i+Phw7xDJF2w6eDlNffM3Hw227Shu107e6uNHzBANFziAP4F64drmAX
u0HKiGNWGEZ4fWsozOmWsEOgJ+BLypFRc5XkcskAFc+Oe1VGxqejcyuTeoVioV5E
UJ0JcMypxSryhi8xyYCg0gEwFX3GARRbdU2i9IyEPOLg2wGh7934uj4ghQkQ3a7h
zMxECDqnHRoPR8FHbNsGV5cBZ2ZHhRQLB5SpZ8/TPGxd2lj/+ziu9V3jb3HEtdj9
0SWg93lczd0RETIX3tc73d6W2Daf1J75AMPWBvCkKO+6G59HQbGHwpNYk9Lix7Qk
YVkl+VoyWcFlc+H9DtAMbeUe1xexKjStEN1NHdsXK62p31rLKUZX6pfCEj9XPpaw
2zv3LK+c2gQLhyygPMFkxMC/eFwW8TgqnBuiWHwYSFqf9cv0vLJVgozt+7fST1LS
6hmM2iC4h0dtfKH1iUaUFGSEcyQB6Ztr5+m5CKTaEZTrPtIv0iIVdj6FtF5bJq+P
O1Y2j5qxumYvmgSXAX9zDB+gZZq27xOftgMCxRxPQ6Fo23lZjlyQ+pz96Yi26ueP
cCYpu0hCS1acFAUJq45AgKdppMBcM0hZ3dDBf+zG9bq9hvNOYiSmXs03O9qBwmFA
kMPTJpJz87h9yDwle7NdADo+V7TxMWc025y2IiWEAQZVyY3S7w7MuNRy2sBuTkRB
PtCxdADCjdjD9mmysGh82MArvRr74erbP9vr803dSdCI0Krg/AXDpypGdFfWphVA
JGHp+5xA0r+6vjqGIBD4h2MMwDUNEQBrPWzs4ANMCAr9Gnhe5Ijg7ft6woaQ7dIC
pSAmiUxAmoUzZ1uUQvjR6Dd3YyyAvXYSILCgEiYJYLuLTR14VA+zDIzDPHS+a/lX
ovMum/Gr7dfV3vrLFReM9EaVTN8pJDjJiHEoQYzxwR60h7OYzK2t/W87OHF42gBN
5RIuAqOM2sQ/Vsof0Xaw1hL/VPlFQqz6+jlYKkIR2HxH4n7mUe8HRtr6YM8HNevT
ltCzsZoek+z5CsDBVYWoU9OzW6pCqkqT2HWfdmAMilKx8pYlFOU18BCLmKZvh9l/
HzZWo2feMIjldNGHQN3Wu7Xwed5YzH+u1xMLijkz/0ekygcZq2+YKAEewj7EUsyn
PdkeL8ZalAO9oxOVyzpS7Yhy3i/ziLutGaMkKHEfcdlz0tQqUv5V8g1dI3Xxepv2
S+gJy8+ScNH5Om0iGDwA1wPdvoEdmfRJjDcGC52qMCnBKQ8jFbkFfl3SC2BFnlKf
r/Jrzp9I5fAlJYzfiZbcjLTPmTQcCzEqMyaP+RfRN9pWrkdAZSG5k7aSEMLAgJC9
QUWCBzRiCkASYuGmlvdcG6lyJ0C/B/jAXfeAjjvsNcM+j6fk5clzs/jWX7x9FtP3
qsQJ0u4BSZFHqpHJtgDiHmS/J0rHpRbUnpWHvmVcUyd0HV1F+snzMEjYmrh/TgTc
T0mpSB14KwJmp8UudQnQpgEctERwnRScAybrbDLB94JniPglwXFN7AArCgkI7p39
E2YvjMKWt411FswT6/52xjtfxXinmlpeYZebY9GdcWIcTAqmvgF1ZfYwenc9aGUQ
u2RDbCJ6xUupHcwwjtvLVuUxeIuSBPNwFkI8GadIb6+ZpM2THo0AWI3ocW6ljOrS
Pw2a2HD4foRD7Oa8aPSaw2LXJomXxlMgQpvReLxUeRBb6qmSzhmMZwJUGizQY1Od
K21xCzQ82YjTS5FIMaQUPjaSMJYMgtPJgPgYvO1ZF5/KrH5EfsecTXgS4sJS2Cw+
L/Kfg+86JM7gvS1UuoYkUtj04ovQS9uGyVUPIr1gottLXJjpSuldUGJBvgBez4Fq
q1QzxhlTXb87dY4wXfwZBseWGVDO8Yo28qF+NI2o1/zJPmlrxinJUqCqSMwdLUKq
I5YkXMRvB7Ua4zvjRy93sTMq9DyzCSjmGloP8gNkwA2Dhd2Kx32kbB3BbsvxY+bQ
JifHLZ46U1iS/XrUYl4crdBYHhaL0E169PXwp7l6jtfalbNbDnBxrAN6H1TD36hO
MGcWAKXb5QD1GXOh4CYThi0SEOaxrI9a/y7osKoYGDsnJHssXaiaX2RZb6xCDqAO
4IKNPuvfgkMli4z6lyBMBk/bYZwr/qg8P5t+rE3pbTzzA2bFrOjoaU04ZQivf1Li
MTGYbv+WsqBu7b5etAb90lN4IeH5wyTCHhcWIobSs5pgoo5comGE+BI0FqSv2F9I
sX0A6Ch9O0Z1e0kDmKeqtlwI2wXCENr5iwOvI7L+N/9+a240dB3yOQbWoXkZ/T5l
78L70g5FccsFhycCEIg1afnJVAzC+kfEBiML4uYtENFjT5IhClU47dqR+unZhAPK
3i8uiL+koHbYMKlaJK+jzICF7jt1r6OTBK76+z9gKUuWqaxFFGUkKx3TYEqHtXj5
Nld1ThZiSpFhCploeJZEn9AmAXlaqx9INwu7Y55nCHZGaIRcwOqomGlM6CAEMIq9
zDO9wTy+b1eAaNuO3P+hbPDXqMeeq4mqoNHPCU3/bOx5W8ppnVU/oY+RHwZ0/jEQ
CIbPm+EDhGT8yOgdSCx8UuIR9RnN5dCo0FauIY2QXU85lbcqXAZld9qKESwVF94z
fdoAnN0FIOzhYFmgenwEdkaBUfqrBOUEcWadLqKMoFEQreMVzgdtIEhpBUSnuY0G
0jOpg1ZKa/vzhovWwIcY1cV3jNe3Thri+F1tm1yIlUNhbXX4cEnWvQmGalXFJMs+
xudUVDdoywmfDEqj7Wyowkg0K2Tqts1ppL0ZY08SAljdoC0UVh0i/hFj8UCJSOoI
R0cSGFbU6VQZ76Fjp6cUNOfNoGQn3AEjuD6cC95wb2fy1io1mQztiI9wQNTRLadI
dRPivu37noUpkJw8guqHHvDGHl4xrbqVR9Tv5TH/5Gv+4DZrEdGle2XMZmCI7y45
5JEEiynDol2+ErMmLvXDvJk0/bbT9GAW0oIQwMaCJ+kqlnrPVmzkomCyb1E08XlC
XqkD/O8cfdIzM/3KJqA6wU+JinKpjjNYCWmLFAtm0r7PHAbKIp/fCFVw7mN3zLAq
Y+bpjhSrXK6nQoqsuB+0dnszDiQYItYx6ksGQVLYZWioIqM1TSazq4HyrkmcQLt6
uzc+w9zLclzHTwHnnPwyL8n+DE48E0wNM5e0nOmYxrORoo8hbXk83dzs342Vr8nR
+bRMzdP7vE2RUFw1mbo2v6os7OaGwddQs8vlGVFakSL3etCvR4kFYD58fgWnGF18
9bGcoZklyea53UnC9RLxdbjkiDPMrXtdi5vEdWT9TYZwMlHdynVFEpJzaS6uIfRJ
BLm+AAdrHWb2nPGxhW5f5S8t9lEolfDEqifp1NL5aAC+NrvEbLGoNzq13YS/y+lb
v5rlRjUPSeozbDa38xQ71wuI25Vm6ggiXkEe3yT+62pUXbIi6ORKwhidhzNH8V6G
oBkNxMT9a06VE+zVxkZ44p0lGKrn5foVEIaP3lzRCt308FCflRaAe9HHdp8fLEP4
JBHZoryZj6w1rzVYWMPLnCaSxoYDgx2IRc3HGnrX8tpoIXyJYIKxeAySSNde92mq
Za9m67FJ8QflStxHimKxI24GR28cxR9D3XhucVpO+kP6BD0oJkVKOn2Ag+cv/KRu
wmYG3ce9+hJi4GWxsYKgfGvNrEYBMfRwF6lxtY8eVvTnyBA3fSNt1oMDFfkvNJG/
NJDXF3e8Za52IiCNQIj9bix8Blox/JION41KYWbGB49GfwturvpVDfRKIjKDSsbC
Ar4cnswURPBxhjhcjEXqNXooidfvrG1vnk17Y4s8cG7OZl4/Mxf3MrkztpR6V6QD
HX7DOQBL3vYfCpZ40lXlF7YH/1VZ8eFEivJkgKSSVOM8bAwMR7Wep/U2hPViyLra
bsFeRlz57RyCHii8Y5hH5+aDqkgcEtYJ2rXKaKOxsgUNe6MT2i9R9fiuZOxiQe3P
/b5iajsstmIUH5wuOLQXKDbFj+gFZc9hAsuc2WIJIYnRK5U4AYVRTgFinF+puc2E
s7I6ENpSaLJBWgIzgHmqqO5+MQnjDTSUFKHhxI//yShc9yOU6oNslQ9Iw51rzJ7P
n/1+lTZ/0SHAsU5TlacKYYAf0Zymic+sgVoAgXNIwqgnS+vbkkWXPCMZS1sTkJ98
cy8NEwZpH21jecoUWu59PhWvzXCdVr1wfu5OCRl0GwGk8F83kOjpXEmFDxs9rVUu
W1y3q4qegH733uO7FNgbpJcNG+Cu9B50bUGbxh3BqLwhQIk9Z95MT3CE77S++LfP
RF6Sa94I0cVVUannk5NxdoxWVmtGNY3zwpPpPJD3AujWLqzb4DCberlYXvfgprXE
JslOX0eXHL6Ot00cbcvZzbwEfHxMfXSA/0wxnxD7OGG2o9XukhnBcwqc+WwPYHPA
TdfY/qGcwxQ1/3AOOMMsVJQsfTgIkbXnvmbWKtazkJqb8Fj5g8jX1s8N+aUgrP2O
ak3TaOAKENdLy/LyBEioQmb/nHcKboGrCwOsPcaUfwSWWRV+ZsGRfh0lMY6hVRpf
HNaPxkowu2qKKzHkch+HlWJaUfDb0Jy7iYMG+WCLxaPZQI5ct1C+sZEmPDPmQmJs
xNn7uR1mtDawWBNejY8zS2gmo3tuGd0h4k+5rYHbLThNB0GmjAMhjD/cw/ku24GS
6bK+r2sc5m42h9Aka1tYTADLfM9Q9jKhy5dZqrQn1r4Ic+6cBoxKsSlaoYzenUAN
3wxzgJYpQEJL+VtiuvQxx4phO66hTHXFZqM2utMBjUpWbQQqOOoWBR9zNaXv6kM2
v9nExhHyY/RPmxdnkrYhAXmVclg4JAFLiWlxZwaPF8Ko4BLmi/vhTUJZ5WZGsVWy
uEejU4UuvUdnmglr4cjVjTqKwC3yv51NlM3+U8xY3WUpACvt7NuIZLsQcM5PmCAe
kR2zjhBnagKOYlNX5ep+DncR8bD7QOBCSHvew1H7YXANZDDTBrlV3V0T/8rtL3QU
09aAL4Y3cIsdxetg6/MAArRh5sZkWZPua5mMxbp50eLE4Fh8947mmtR/8AZ/H2an
0uujTMzHWv81Bqkt5aZsFzGTfhjkxAIq98bWynD+7O3D0fC8BGHNqd2ScpxhveUZ
vkhYayZQWMel9iAm+Ya/ijs+h75flR/HTmLgogQ5+3scJiHUck+I5a9Duq6uxtcV
P7wYaA5gpXJiyeXn6RW3TE4A46P/0n4pN9B2yR2Jspv4XRX0xr7J6Zo0JpSSWlf2
qybciZO5rKikjr+HRPmmNPipAilOCkULe0xm3sfHmCGp+S4Pe55MhkxUPLKRLxjs
Fs28/Z57E9ulX8Ut6ljl+K6nqGse7Amfjwa4ZlTwZBFXHSiApr5rRiEk9KGPoHx0
UXwda8Cv+UzUtA8KClCPxJ2JrFzNva0Ao8M1zA+uJZ/1iRCLGmisqjBSBQ6+iQ26
Tr3pc574zI6irOYeStoZL4akh4V/RDz3wA+zrABqONYhddb+Y2sg14MpLAhooLjK
8BXX1yMO+dE8PtQ5NoIgEvaqSuaYgBO0I/V7AyJg8xQ6EfTBJuhPOr9lOP9zB99r
/L92tquWmR7nIVUFKAlLdGc+yDreR58+JoF64l923D892+NeyaPmHQTtGgKeLJTs
Yvjl6s7xUxnOsg4w7A24dimd1Df3l+hEk7AihP78tMV2gjr76Eqa3wtaZveB14mX
ZzDN5vpHP1IMDvbnTixlh+5mmmGvutYxCCuHkPSPh/Ptoi7REneRt1SHW9oAUh8V
f/cmjJxEQIFDCkryRba9DH35FooTM9bYgoypT3nOfhEpw2umoS5AtcW753Y2kjyd
WXmLmBrIng6IDPLGAnnUTzlTQLEo40aW4qZp0AIxyBwQy3P0usthy+H0M8q7dlBf
zIRqmU+2oyA/vBpVs0Xj7TCe0w2k+ey0/S7RDMXmCnsC5+VW3IXhRAk0DppILhRt
CCD4DZB7cpjAlZjrD5Zcpvj0EMeQWcgmWUU8WtIntjMR0t8tCV4wDFC5i0xuiRZz
3yq1TyuoN/LuT8Q1HG4yrBPjum3FBeeTQa4qnkesEA0Usmc2GAVgX5vVsOT44D1k
EBpuxG4yShH5eiCGYWary/uIcQ+mkJgFZzVpLRyKm8MpNvoDkhG66oN/nRaS9CdN
fXmdu4TJG4OCOho83reggarP8HiQB+r9bRkWQybxiXcAr7w6r/Z5cY7WB6uk0OrK
dVHWmhfPvM66viysujFDTYb/yIBYbdYyCqu8MvGmBjQKoI1kIvzLGRP/qvspTETe
fSkuHV2PtB2l+QFR4h00pJri0sIxsBu4kOyw39zyGN+VoFVtkVQ4ERtMIASXOz0t
0OIyujXNEYrPdJp8TakkWg7E7FyARPw8sUAiK+u79UTrk+zVID2yJ9Bi8WFnHtIw
0X2g4IBxKa2FtUlzBo9yMwn5G+gkmfRVtlAeDJViJJKMh2iPFtsozqXJoigYFgZe
nUf8jMHdvISL0kmdEg8NXAvUMPGcSKQDZ4p2tmomFEc/TUaQlDNWgxx++gSG0ejV
w/06/BFZ98BVlA3aS8bW8GV1h/ARnszxK8j2W6iC+LynRovU0Sv93xGmmmYbuu0Q
7dKlWbCKKPtfr+CnIBAENw07Vnt0WetBlKlDbu1Y87HmncKUhfvYY7Dkzujk1Zlk
5TMj/dJB2htaaiIp7Oz6UDWOT293c65C2KrZvKR6VJ/YFaIF63JvoQu9402pcifN
3+MxHRa3SRrk9JgR92x0DEm+L8+7lpzxEc3YGRbJAMTCHaOCMVaBsX15O10epCDI
SwX2soVkbSTUjzTag931KIvjKhhnUlhsDO3DZCk4Iw09QUm3bbzB2U2EWxBbkBkz
UPf4uKQO9xdC9vSNpK89URGlHm6YLx6zSOP9fY6HkEQ8WPFs+pQOVMJmryhWggNa
45tr96AX1KmOiPEMHmsdqegl5lF7ewTu8ZhqBtJ6r13ae8mIU+SHR4+vkZrpmw8l
nHjDjSRWrcxjgZoGILbGBCnJGeJc4mbJusOThTuXiNwVkpQS03Q+l1ERv8yyNaQl
QjaKfNV8hmyOBcbHlHp6yv2hlgiPQXIV2uMSCzv1W+ZjzOhbN2u1e+PLHYkd3+lr
01MOFgpwQHqMfOoS9gBBrajl5pugPyFOqqEbYwvnZRIOFHJMaXOvQNo947VgF8/R
6hk2YjgEoQASmPqxDprBCCx6Ijw+u2kNrw24NZmpegCiJ3Goc5e5cvxbwxc6E9bf
Yt8CJEeBkiW3LvLyhCvziRDaktZurNYROuShUvjYrSI5xEgis6x2Dpktqk0NHbs/
0F5tjpVJrtx+WEtPEGwBylwhrRJE2xhbYO65977guScKYhODZyHaOiPVGKndAIso
EYa6g8Oz/S0J7xPWzx8tZkS/6JMMTZg2MRF3kPsNUCehwmmlISqonaMZVA0GnBUk
ZBLPOV40TwPFlKRmlAJT0fxbCHGZ/rgNc1HSLSuwvtP3tzDCNZQu4mSE6/15/bUX
PPW+Yevl1K13aAoEtdIVZyHnxMLwvNgdjN/4+lu0P+rlvDUaRYN6anZVUtig3KPV
VJ1mhYayFlDV2pPFMH9q+1BRITl7inBxDvAl4hb8UD88UiQcp16Ib2mivra8WrFz
PVIIS/H+BKWpp0fkfCYQlVLf6Wub2edJkey5VloM3Dwhkt2AMapyFMIzPqnmKTYN
wMemDtJiqUGSw2h3R8P0A53e6EF1DoZA5w0nAEGkCj6QhFr/jE4sZH+hY+/kTLdd
wJt0IdF4Lhk0rl4t+liKiW+BHGWhXDd4F263ZKLiAZkTcWwCPJm5uIwSY/3TOA4L
eQkqNLqXk/2WfKWt0mdvzHNALY9GyhBN3AQaoqj0+WiHGfV6yNVKNgcAvhdD/dnt
yJw5o4R+3y0kiKytqjfBMf37KPtb0i9dFfIsA/M7C5Z6V6ktGULED1raVj8UIptR
YoPYKvEwjj2SNG5AW91p3z5fJe6N66WZ/59SBxndkUKTLxP4+AGf4NiWG6n9gUfA
RyupL4GcbXVfawEBzkvkjZV4YWWu4OXLFj3F5dILtLOj+x2PvyNI4PqcuH0A2xax
MOa4xU2Mdo62iaCTQPBwxCb03AOQGpFKaWBTaFtlq/g5/24F9SUDIvPAx2CVgkUf
9gYUvmfJdx2lai+Nl+Wo8gS+l1caD3xjRb8SW7rco7qJ9800q/vssibrm/AhHPZK
wD3fALkRf996Aefi0V/Vy8uo1FSVzH29OHEuMbF14NCgmA+I0t0z3C9+p/AAI15P
YhigSFLxJnzUEzUd6y6TZBT05lRyqh4EDIIYVOh8+ilMOw3/mxkYa/nuQJpFIzqQ
CwPAcU6DHc7YoJFpIkaPZIOmZq801BWNNGJ6z/d5GcGaLcJnlFixI+VKwb6g2Y+V
zZwcMp8Z057Y7ZMovh26iNxQbQ5PvQkOy19ovd58MwO/Zc1f+UCJCCDyugq4YLNe
0u+uOjcl8rnIVQp6STYtEwcszC7KI8iI9Zo7Hg0Nvjt5R0NvfmNKEk7j9NI3u15r
0OK8MNWgiJBKULgU8IwNl1UYUNpLEQxyROu97Y/LGrCFFlhbMvluUOQjCzfaZXEp
95LZYkm/jaiXStfOj6MYhcRCtWIfApY8zmnjTbUXETh7xYTfJP49zTZrsjx4jATd
2dsa7RKjz55Mh1o9Wy9+8/29viK7lZxelH3t9vCTNBztnGcfg4OfOGfvQVLEiFjz
RaZqPHUw9nu29wt51CQHv15UBeMEaC5499s3x5bYsgOTZnVF6ddHgR9pRN8dLXp0
uxyGsG9Yp2r0Vdc962ObxSjeZVop4R1gcZ/KkklTIksWQlW4cpfhqLjhUvsRRwfK
u/5oc9kA+yxOl1CJ7/N21k7B7q0+IejZjI8PJyDjNUfpUPExfG+Z49VPD0xPRakv
hsUNmNZRzEjWtoomdZ8SLvV80Ed68AoTqfwHAabVxaeRYFjgsmu8FH7IlIC8tN/p
NImv78tiyQ7tE1IrIhyK8s2ZwCCaRUBfYMuTtxNln5QSwvWtELUbsMfDqBrHScti
deC8vi3bUvxaPh3pMBZOlmvZlpRWEWAvP2LWYdL/gqfa94dGyD7VPl9apoLFmCpl
6vkCrYpXFQudw2Ob+KVEB8TzSTwu+BkkvXmD87G+n9l39ZH38Yb/TtRJ0GrAdEdr
vuQ1+nGCVSBslTQQlbrPKDRGm9zgt2qMYLzWjzdQHzfMlubIEWH5Pw35AWjgMiwI
fu+Sib+2VGBqK6DxH9FUsyse+WdfHnJHdJ585sjUCcdWNtrey+7DNFbdP5d6TKy0
DyGB5RTVj+P0K8AJ527z+z2yXjAipNqh05Nm5CDNgjJhV8LSPB4Vjmz2cKouOMAP
mSo2oZU3qZc50bWjWCoUBWhC4vVGWJy14gbbQdSi1FaY4+dCkDJfv7R6UpVUZEdA
mvh7cM8lejE1QIzCCEfQOCvkmAKY7eIZLUFfe1WBmXCiTT2p9+bLvOQBUbAQulSr
eWI2/YsKBMZROZeMAjuqt6bt6lFqeQ5rryeLxhynCh2ztT8i6mDIOYm64SPa9Szv
TY74Dv83ZAX4PE4Dpm4zeXtdCX1Ptp1M7l/FKxV/huc/fjDm6bk6reZXyDJLf5zZ
GWeZQdJTvIcCtmUl08a95c20hfYjFgU5MBTcIBEpupBXSPSl/5svEdz4Nlw5TgI7
T7709zp8k48rlcFeobKMSXHgDQfbDOxT5qxDt+vTduXlLRPd8EQI0fqZqGXA7yiH
5vV4rXE5OAL4b+s2WTWLb9sS9zVwND7iZfnHedByvJ3P6nCj5yYpx7o27eOh41aW
BJ1PGQ87qvOLGGbnyNKCiiipYlkQjUPjjQlAeVCyiJO4GxVgHr/b5B3+gpQpePcl
NoYhOS1X3za6oSVuYHiv8YkiEXZZT48fq4Pvf2410/iuKvjDRFBOHIjHfkvo6RHx
/LVRsRxQka/DG21WSDar+zoC8Jnw3yDy6y8QueEXMmb6z69CLb4JqCq6Q7xW5JAT
HBiuYDUsgSZCKXgrtHYVeD16Ht+wz0wFJhs2N9gwOa0kWhCdt1KAroXARcAEZLU4
FQoF/LPAiyxtKBPzfziG+bsCQtRbsXs7SkO4qgFRkMIhxoRgHVeP0ATwZUQLsXi6
4madXnM4E18BSlsuFFPySYuFiydrY7oKhcXhrXD+YXppTa2xRx0n4AyvE2q1vZSQ
n329PpuCFINaOsMqehM8I2EsghE/Or+imcpM12nXlxQ0yQmQVkNsBVK/Ckww51p6
BRux3yaOj30Obdg6TdWS74yXaASx1Ge76Weeoq6qS7CUhGLFA/PKu90PBR5QD1Ds
EPJAqqYIT37wMfoTFcGTABJKiIirMx7emMUIv9Xvc0wZr0CukDqRkQ2LeE9FYluQ
l/W9IgLEkGb1dBh0SMsv8YWnzF1hKa89nnlGCxbVI74HMw+MospsYKog5GgLqITK
mb6x9Al8MhIVQTVwy/j3hJmrn6tUH4Pim1DUYAXgHZXqe5yn2GPk7sP07iZRH3ID
4udHFVAe+8bvKDr/WBYam6vrpaX1cVPhK11BY84lNoqUCus2w/12wj/HNyIA7y2j
18j5UNk7WTP1DNAapySRwMFxidYbHf2zPMU0P5YSvZzQxz6rAutUIgD/qqGKdXLo
b6yVrPbW4K5kFwCcXnqQQ/UBdwIhpfh8JWy8lV1lDcLfgwGdp4CICE+YK5PCh87K
0ZsfryWcpNJeiUnC1EmVkOKtwFbJcPBQbO33HNQqBcPCZV5x67NUowseAw8ESqPL
fDM9D7KIRIELKhQgq0adT2+Hte1CFYWTZApGKtQcrWEwaNCBYDnDFKKqarz/zDzD
ypjKSFoFPfIemNxDC80gWVGmY8991HiDkjhJMNy4YU/X1NXZzQKfB+fch4tfyJVQ
uESop1l2RNLuYRiKPAKYSwKJBFKehkDRSZP2/AQ3BddePQHI9Zvj7ltYSqjiASfw
wONpATD8rtkzHzqc18zM+LJ7QIQ66AonNAXZqHwjLbhOkrzPq4vtKytTr7AExiQ/
5nn6ZjrfMMsYYsN3/bPKgVEhhyJt4Z6YMAJaDupmTLu8+9C7yQE13ddcE3PE3Xor
RNZt64IVoZTclyFJO77+U+JBW1kjTurGt+LwDrOiAq7e2uMbAwnvnn0HgdtEpFbB
8zDYs2B4WcdswVoK8PZuc+zH6DJAozBEfW2Va9YNlyld8oJUEG5zXhXWxJIQeAv3
9tY/RoK4EcBBqx+1PZuObn1VUHR09hZueb+OGSMgrUPGJ2m1g08PHCov+ZESUdLi
Q37fz/r3mGRRg2n5Vp9kjusGubuiAtzYgGiweY41R73FvUmxwjentkWVafd+gRiC
dIg2E4uH1EE05T188DNI6vC659U6OBSGHrrFquaPQt2pAVK5MltxcggBnVA1PBey
NNaTAF/mK4cRMdMv1ziI3Ofjo2zMi3mgA+2NCrLdKM0W3IkRPaJS3AFZBrZGxorn
OfyU1/JwGwDmghEgWCRyE0s+EkpODDHLCpq7qiQOjirU4/Vq7xBbFGwfa43uWscT
PsMFpM1mVUpLo4BrwVmT0Cnde10Vy8RAdo809AVZ4zFVvOlhg6As/JPapEp1X7yt
32Y5hdixQU08S1H5WMJ2/vk6CLDnfkWLOZrEFAHMxEdz3OhaI5zjbtb5BvOY4Y68
bovg2jP/6/bMU2qfVLKvYwH0tmH41UF7GHteO57krY00N7w2Vf3lDei0avuwpiQ7
r2Fam6ogEVUxbe7vTkgAlddBp38HBs+oEf71ZiCFrzjc99am5lO26CXyTJjnY9wL
wfmSTzidmcHN+MyXmSg2qxUDANSMnQ62Se2OnK6BaSIgrPmObpL3z31hip+YoLTy
VQIawIqvyUv2cU9rdWNeyZXNQHj+A1yjL0Rx1G2MTmaG/kiUZQMOnW5MNpQSgT7b
wJgNfdPyzKhMHVVrJvh3bpG+bkd3QWVDUjsxQ82CI3Ivhaykv2o7NBdvnUjI7kGA
mco5265aJkK9ZQtY6yIICnT43ND4OpgBZV5jED3/SIRLAtPBykh0wKzAL69a3tf9
ApKsE86Xcq9xTTAkFnoizRCeK8RXlYBWnvWAE52fICiWr3zAGSSJ6OF/63yb5fht
TsPsn7ylXYtfM8sZAOFL4Ut6LYT7wZTux+XaCAe/9mP1lI7/vzE2xBSAWygu9cxj
+664VXtYbB2+zMf+bpkPHH/SxqN8Ai+bObtHSDVZ0TB7YBUloO24ZWxVg5iD2fdW
fzvVT5S1vq1YzrYnlVjPaNS6STU3qW0e/eiEKk/6IefwWY55DK4ANttxgPLAJKPP
A3vk18qGvUWuM5Z3sgLFSEHLJmbDT0hzdrh26D0FicLLT3UAD0cAQHf3NExXyLX7
5zydA5GGzqHePMa0MrYND/ymJFdemYaXj4leghWizvuROsBYXKC8AE0R+2ofduns
cP5WKZcxnxhwNh9Ht0Iqd7ZfWOwpBOGMTJW5Yz0WEfTrcUy+P7m5Uc5S9ZAC6SGk
ey7PIO/RxLJtrbua+VSurgYl7XVg7jBApG8kjrGVMPaxRSFI+ML8Od/mxsllAs1/
WiaP0dfnupfcEMqaDhF2XTNHchTAC20zdwImXQUIbXTspMqQvAEW4wE+OPK5B3gE
TGFUe7sssKFpkKqAOc4dExFIf5SLyRc5keWVMzpfHyl6/l+k1WUhyq0BKOsiktPS
V/smB2BgMKstXiFwdyFK1qtKSBLrOAhN0HaBH9sDjxrf1hgB4olCQHcvdkYrhpDw
N9B8gk9pKp2YAn4XpvmnoDzz/E6jy/ncmd6xnuE5HrCNl1t4F0z8N5pzl1W2DgOg
U1zPoo7xdk7K+WfAdmxsmyj2yyAzSc3Pz3hckQHaoCDAJ5Kz0CzsMqOFYMDbJ8ke
BpD1cJX0FbcYMiVbYmjgPL8zxImacZIC57roa+XiXBlLdBUJuQrQUI5rtB5R0RwW
XmQ8/oZa+DHT9O0i/nD+FeS6enNdlMZMqU5jRzfPOQfqf/w583/yp+S3ncjz95Sr
0Y4q4Bnly/+WeDikoGwWzzYNRmMGMJBVTUw6PHZKsK5lBbWjtzlFqlljvcIP9bed
knSvwuGtjis8x9Bz1vHjXG0a/DSEijiFQElHq0EZe7MKAAG8x0oVI0xNZwdnnkiQ
cwEzjA4wmWuoaBqAvmrsIgIOkvePMbwg66ywOhiKkXkO6nqOsTioHomCej0M/j5g
SzMTuap7Mhtf2dvTyzy/9gCbtqu81VP2w5bBOpU6FatKy9XMGlmSa8XX1ba8TUTq
F0GqAoOb90r7QnpN1CxsyKmrnGDKN+CtB0EAInyMWKMOpd1EPa/QhlWz3Ym3q6J2
knGcMN0cbmFMDtq8aaiK3QRsLSci32eF3aa4r6dfUD9yJ5tCG1JSA5Lcjd8HGbzK
qB2hz3Tbutil3Ae3PrPRAMehoC30kpP6ya7fsw6pyugRKV3TnDSJpfv3QnIiOPuu
DDlgLIn8/HG/AeVlro4fFEMbRBVroBKHcrvaKEwCwHEGnbTbLORdfaQFQfc3pxZZ
UqwjwogJobHRJlUpONUQkEMdhnwVdoXRYcwPUXnR439MRKSGdguMQWA6jhcgU2NN
RPZDsRFt1ySb0GfduCBg/27YEWN8Sg+pblh2u0XptxXCBwl6LGT896z3A+dKEeXf
J96yGvPh9+otX+6U4yCfEMjliJ9XukPavoz3eK+dD8kigBS+uRCDsX/oWovK6t9m
iODQDfyS3hACJvSIAciK+8qWOKBeQLWGs0J/4ESSdcMY48nAmkgOUmh4195rFVeT
ESOe5neR0uYca9zP4MQFb9VdqDrL2Yp7s+13fcwbIn4Ifh5DJ14ImbQWvKuwiYiA
D4XVhyk2H4pZGKPqtkcfR65U/TtJbfW8FUtWkKoY9rM6JIPjA4rmMPE0Vx4rdet/
XACK2tYAIWmEz9G2yB0LqKWEnziQvMCNU4SR5RRTvaFcD60Cs3IJxRDzecrLgyFR
OTqRJQkJtc9yhz4sQqzHNPvEmlMaJP4OMHfGuSskRIFim29jhySepebUMJtSlpv8
e/sd/afeyG4eR95I2Q6TLRWMTD2Ebq5QigtVhlVGIT4+Ob48zqxnCqerzY+nfoNy
CX7x8TLtp0w65xhb83b+TeL6owSoOpv1zER4rEfL9Wr3dSXcSxJkoOCGzw8TCNjE
prrN8yrk1XNSE9QeEwKK2Kbk8Z+99wqmEUL3T2OXCvHyUAihCOAnnrEpNn3lOJPf
uAR3IVozWgqr3w/a+jQvvQoWsWSIVgjA6POiDHiSCtNesDy/3veIKN9gdPbyzeZ/
LTpkrcR3pymxkaWr47utrlb/h5uFq/sPES7h5Nt62emMbEaXWsrbm2Z57OzKcOts
kmKqLBuVT91EJTpJLhFVMJVwi0/pqqBIBKGZMAhzSvbuqAVh6yx+nmsy5NHG11jY
8bpXPDGrQo+OweHSx8JopeOFjONWBilDzuqbqDH3ObBc5j3mLiHx/YCHp5fOAyks
FEFuBEyjtIrVG901Tox0RGmkn+mpgdDJoP1G1eNlfo29OYDciF6QZfOjk1FeoJkq
DUaLIH01FWjJClmzZi9v5vyV/wPVaUcHS+vneHwB5uwgjwvrXOXxidr+xYFefrni
reqbY1YMyfB4F57GC+hTMRfdOUtR9jPCpLGjT4iTPXByrxYPaYEOKAAw6sscW31r
YTmVfa31pflZ9AKHup9ObK3W0zjKgx9mNbZWxjG0p+atkAkNacx0Tj5hl1SuzFjF
qJmL74X1UZEdaZb8l9Ou0h9ik4oyGcRcAG64TEMxCYM4mCTNDRTskTUGnbKUBDw3
XfctniIRSh2AVmISkgLrb+NW4V5axiALz/aqEzQW0z3b45Omyo0vyzy/3vncPh5W
2LkOszmm4H7q+E4olewLyTM/IqBQzP5dtBPJfLlVEyBYAdyAr9GNW5pLK2GQrV+z
oYLrz9vI70YeiEPLj0RMn8twWfmE8vnMvtjvPL5y75UmdzQQ/7JoeMCsNt9m7Yc4
MqG/6yu/ORuyiyis9iD3Ox0VR+ZhtJfxLN2PCmZ9+2D6Vx8CHYUEOUricHq/PoE9
nmHH+mwXPz3U4IR3yH/zkkyZlt/BX3QLGJMpKP975sC5Wp3b9wfL+0wyHgwlBy7I
Z/YPctW8q252W4VH5kH8HaActGOrZKMVBOWzMNxgrmNFc6m6LKc+s/kqc1g8h2V0
5Gh3dSkN7FDvxruz8oSIisUN5EqYYVGPuUuQpRgiAr/SJoyjcqj8OUImnjelqu5c
2AEaLroDK3lMCE0cEmsrEd+WN+ywdT6Hd1M/pnZEg6V++V9rb/IxM+DUawkE6+IM
VqydRftLNELSPnjxXwVZh6BBIjbDcibuzc8lxkfxPFJ8Z3fx3hPwR4eHVHDNUUu8
2ERt+FMC1jLSWBjHfkuw6fUvUhj6VwJ5ztA7YBzo7acT62HJzoz0OMVxyC4DVyjI
CsRslcL321TjnWnIWZm820Hl+fEAF1a9oeFUrLl7snpYIsAvJCIi7xYWU9VOEI51
+3CFE4pcYj1ODBE8Yh9j4Iv6BSyXUAUfTCme29F2OMRTnnX1fdoIIRzEyHlIH3b9
q69qYvjxyiUKXnKz0lGLYQrINsgt1V407yU/pt9QHGAFxyxt7sAsRBMQmgU7TsoX
2KtGX46zJDQAS+bONZ8IqHI1LGvYI38H3WszfbOva73OS2FS/CXUHOKDty7lr5x0
1ECSuD2FKoUP1p57SYO6TPAY1pbqdgZ0x0mgORRSI5tDgZzKwp6mUqi8O2OnSOPO
nbyv1Q5fnhhv/1SN4Cv3XQ4pfTKfqNHvJ4f54ucFxlAhqCWPaRkRWGYE6ZT3BPZv
fS3W91jWTJBAZNcIa9s0fKyoQvZ1clmW4PKR9f6bsKQkumfeaimsJZPFg5YJsrLK
R0sCiJtOUeA0xs4qLAVWXGsWTFDtOfY2kbdlfPnO9KelFDYcTGaBktg00AEmR4eM
uxwL4lKuWINqAokgOWEpqasZSIWYoK7A+N56yZtUq2W5MmnqoQY87fq+/kClzCZS
CAnvmWm86jDKYoBtXEecoGfjzbAh7DsPWxgpEig9DpldWBwrU9tR6dZh+nWbui2t
JR9Exj44K+uEeznM8k8/EFNKX30P3kMgVzhOcZId2KBAQZN/D53aGmBduqUtmfgM
Src4+aIkPd4+V1O1uSdZnssOpADCAmYa/QVwWrefMhNmOI/7F0x+rYis1hWoydo6
IAFg/5mpeebS24B+48MBmh/UAp8dzAewSN/us8DJYzcZzoLxliP2k5rtwxav/HFl
c4tAQG8gERky4CMMNu4Xy6OP0D4laf05ZhzKSbpRqxoSUQ+ESyQwUES5Y5+tZsKF
cqcnoH5cxUm52sg91sAttT3Til1rKYEfUwhl0DSumioOjyjHcWbCIBvqxsuPLpAc
hucqK+nXCkkbG7Sd4X31y2krklJO6WEG9CAu883OkZvTnMtPbGo/e6YbKFM8JxGn
zzcxmCvaBjHc6qG/FEbCyQyI2OX4NueCo9vupl/f7dQu2W0+4XmN2VZJ4epaXqB1
lc5OrROB829GKVGkrZlNoGB97pqP+c4RW+kcpz4WYX4aYe1jLavOzhuIfPlMXGxV
2kA0GwjQQwyjNVS3Nj0D85kafxyx2Ef53OnUe/v9RtL/EL2ookSjCrXXW/Va67FT
n4svFmYazgfP7VAmfFPh5ZJNeJmcwewwhQSacLl6ybgaqPgeRDKMA9mkFogygl6k
nxH5Wzk8+oBU+OJlbik0a0Uo9SwbZMNV3U98/8H9+ryhgrH/FShhodFdt/SqiVyB
8TwgmdNbhwwxhQ7jID2fKTqK8Lc4ZsRvcRG/ErABeU6/ZU4CYkSTBiVcilTUQT90
AWeA6MlEbiWW0Iwu/sGIIgFFgjRnCmnf1MuXLSKggASwaT9zIk14+e7OvZXae0zg
6k9ca3A4hWuJlLEstZEc0fcT5jjayViBYwCOpkC8JQ3+KZN4faaxQBAQ7SZLZ3Y7
f9+zzKXJLuT8gFsVvcTz8UPOvHytnvZTwE7pJbQPCxbe4nmuaa9tNtRFbI0lpQM/
YJqf13Qwu49brHZ6VDLlaNNCgYkEANK8YZslO8ujnHCj1PMR82kIZejVb0Qfcs+R
d3YnyxkmTeBejPc35SOnUP/sqjBx1xtOdyAl1UxEBaATfJub6cP4XPpMX/uB7JtS
os+Bi0IUVvwn3pV3Gg7TJiedOoqbKCuNbSxLUxubRNNJXkUEQNa7vUXoUUTslJM4
V2alS9lk25vIxN03n1upef4upvLcoflYakxK/10v6kkTBkDJs9l5DwK20Y0cIpY1
YCpnH93Yy3b+ohxNf+gQr1xs1eKcT/OgTKcggPSC5oYd7uM+1/1iYCFUe8/RND/1
Ple0YlPdBc76Wd6qARpWN/B2qHoTy5vrMgDInbDOYIY9Kw8APN3ChZGrtkFk052v
UuiF7wFcAdI50X71wSGQ58MSoO9VNioDmTxx+4Cve68MRMHlqF+MrsK/rtChymCK
kSTf4vP4mJusq42EoI7CRH7rxmcneBEdw+NYS55YQqB508krVkhLuGME1iDVoHLF
shZOSk2x+j4jgK7GYH7QOtg91pvvdz/FYWyOSTfvl5ZE4BrK47yUpSJ/s1cCx7jv
8eCnULvdW3W138y4eW6tv7wWfMaYQxQnLoFfG9RH2bEoWGhlUWDHdG4LUuxp3fj3
mi67pIg/0TsUkrwqlrFO2a9DlYvOdYmpOzRmQrGjfGvoub9ifc6yqD8S1CGubodP
bA/NJ3NOjELqqlVUqS0wRV0R3DTQHD3zuj0xLYaTPrGsFxAkOJ0AzSk4juUXZDbx
06Olhzbv7FNUQUpf/Ply4SrGK++oIxC7Kn1YZOCPKFRfo5n/oqL00yT9jQ7sDyHI
Dgl9Sz6dGsMt95dPuWZsEtgbRRTsGF4dVMNSLr+wqYNwQJk3lfs7Mg7n6RmNrM66
r1E8kBSQ2faI9y2CsK9Vwt2WkUp+yQz4NVvz7bGRQbuS7/QgxO/UG50jxzwebKdN
xT4SkDS7fRX6Q6NkwLRiULNHU2jGhfR54dSR5Bjiva1TSDFUCG0TraSM1X3s4W1M
aTJ52SbaVV3bdBp5KHl8J3BH2D0Nk20piuDBcDgmH/X1nsckuUdOPM5BdhMjAMOv
ZRGzqlZXwElcortWvS8dOzMtCGSqcEayjOHzDYZ2ibRtRMu9NK9Ry7HpZCU8bTOA
V7spjSHytafSPgDFJeZhG0gGDvjYOFNS6TzjU46ESg0fUvRKzH3Ik0hixMj2BUoO
6wTYzXbynGjdZW+ewWV6sAjBeWjMRTbDsH7v1exWENcCCXxAoRamEy7q0P1PsL3I
AbejzbI/lcpkZmeAr7rEesOFNk7mNH59K0UcphPGgXqCpzDjtGy9VUFR4EYg5VJ/
+MZbjothzLJF6l45ZRYb5H1QxwNfHiY2SUsTBaE4MOBD48K29kV8knG8ppnit9bG
pGfquJGc7jjhHKTEs2zrF30/lBgzkleZ4SUnF/tG+kmJJsgS5PrULdHE+ZJzu2/2
79S5Cap3ClEJdoBoMaHHD77wS19rLHxcb82mhiRkp6o0DaVZ6Wxft/GXGn8Nace0
/XRpMDTmKN5sEAMhjROp81gS1e4EyRp7P//AOoNNHuGoc/IoBZsJGUrtkbABwN6X
7t3KviAM3Mf1Yhst4QaCi8ZysDtrVIwFRyAD7cSEtgRpjkF2E9ED7CHIvA4F5xbn
oeVahaUPhmRLrl7NSVvtEuWS4YJx1KcYxLwKri3+WuzDKDvv5buHOp/wPDD9MToz
spIF4DbSZpaSB0MecH/ui/VIl1nj7qsaT6rnc3ybdQd0aGmxzO7IzJxXhjMGvTXG
8VGmhd4Vvg+DZODIMzUAGsru0aA2EaZIzg0z9RZOt5P6NzFGCHvM1114z14hldNH
pcGK1+VWdkbpSy7pHwZXDPPEPiSux0uoi1iyfhOb3XHH5gGlg4Pylic3Z4Sq7mbD
Gg/ht4NtGTvmngi3YlFtkM8SmNKisfScahJyo86GtmZ8WLXt4xhwifPM8gnEFvVR
D4jx0R1nNuRKiINPIjgDopVYMZGmQ615iYJ29+lDjWnRI+m9aBiWkBkVGFXv2HIs
z13im8U1hkssnTDLD8+oiWyW44pVUqqbqMKQITbrxBo1nfJORJunCEhReDWtu80r
nXYxC/8YDtlW7Qi6r9arsb3/SomoQr1W/8YtCx5OeqbjZo3Z0kdvLYjOV7wg/DzL
eSklc8/NKwvYtuzn/NCzBTeFkWPwdDftbetiefMWe6ePWhrJf3beldAL9UxzsmGd
Sb8rHbxrZPdt+Ayz8+V7+cxSNTpqChJscuwcQJIrooJv1UVhY0sWXjC0UW0xfERT
MleAKTOb26KMz7HNDvAPLCzbKDUL6ZwvItpmD5FiPltKkvqkbzhJH8FAfCTQeLUK
/+l9bn/zG2bCOBb0lIOgSwb5jQsiDPGBO/TdrrhTGpnUIsNQqcwmivS7OacFyq5q
cCtM0GpStT/DcAkvPwPuu2OstBVoC1KHu1/D6pwah+Ap2LfMkTO6fseWVv0l7MUx
PzKX5YBbEnZ36cpW15CQ2BJ1M+8Q/jscMEGMs0ec+iJaRQtObLlszC16g7V5lVmE
S6z0ArfQLER1Azw+rF16rRj2Gl+lSatbVsdSFw9cQVcr4S0u/z2TTvOJp2fZMDoi
rVNH5uzJ1TP3GQ9knq8SGECT35V3kITGt9UlSE2D02BbgljaXc6ejqGMX14+S9wA
JNV6WbeTOmi13WQ3aZi2ydQwa1sgmURu9yLdGY9Wio2X1zQ0xz9iUzjXr6p3bAr1
iF0E24pHALy682f3frW8bLPENoZQCh4xx7f5MIYJDrnEmSr+4tMAq2fO70B4SPjv
99jLdOw60UwByzpvDhHZR+JbYYFTnT/Rej/Vh7aNNvOYxbNHYT9nu1e+gmpK33jG
jag5w+G8aElpgwwT6zRreSCxlig/eesEeBmlTDDi2mLoRc6NlSXBce22nldK801X
iLxLxQ+UiMtPw7lTqlawhmWIoa3EbKh1cMbFVT1f2dHkHXN/OS9FQw4lkSswrn8F
cXEljv9hHbviOOzewn1Awj9Y1L94ZzPcW+KZWr51ZnqauAVeOEmrZYJjbudqSdLX
zwwp1Mr1VFfdbgJ1kjsqT9Ljvz0p60J9JGxhoWq25h+HxFvMF6CmuCDyl6I7tXD2
l9MpkP4+eadOu3IJehQmV8395nP462sf04zW2QXVtNjEh4xHIdL5o/cH10ZWFbtX
VJtYM78/eyIcQ8Pi26wqxErwcq76qpaSv16i/ETmGYmPlfVa6Pmr3yBd6EQsMaWH
24PzF9RMAUBqIUX0H+sEe0I9mi9ixbrK0dnTafeThLFVNswKE6AnSwQ8QmChna3J
QUDn6h9F7m8n0R/7r1XoiifOjW1wqR7PyHfEIsdTI9z/e0w6cBaQV2sUgCTaXVom
mo2jnxX4SxqOJSIU8mzH2As47ZoSXawGSYnnD0LB+UrWnFJNtHvuNMUQpcVLZi1D
cGBZOf69zF5e/rD5r3iP+RV4X850nXO3nzxOr9S3GNaS5Oa8cm2bywHEWN10wUA6
yCTl53FNDYjkoZ5NhaCdqL39t4hY+B8hLAAzMKA16WhUV+Hv89SWxppYVuOmqLrZ
GAvp2UpzvBlzX0YYxc3n5vI/6MK+SDCjqTWG2QLYQns4VaXOxrksE0x25y5uegDR
bKuh0dnBrblpD5HpAi9rRd3GtwBhQINfEmyUxXuhtof6b6XlWWdzzZhx3zgyc5Mk
9u49GnQY/NCLPvCvWbHj4SFUCX8Vw13UY8YWvYOa8l5btG7PI5/RBZeLKOvmmWqB
j+QOzpFKn4Hzag7kYkHpEpsO6SU4yiX5OxaBs1Dqs94mfuS+twJqs5qvgHmJlxgn
30z9RhVXpGtFCSXVHa37SyoFaxKO4hyZQeY7mDfhkyU0xiXBf7HziusCciKNQmkL
yPWupSIdvQsGwpJkEPZursqbGld7iA8wq0xDwv954bDVdyuuFNdiVXGM72Qt165h
YJCUf2CNcAba0w7w5/lJbqAR9MKrCB6+ukPV0zFvvkA8QV4nVTwaLXrDCd2JbY7c
qQecqMnloD8eYOMjVz9c0S8hXxIcjdnBta9a/LENJDEwJMlUSe4nxgZH4R1wcc4r
0umj3+CnJUS9z3sK81mkT86HEiAiCgT83VMiOGx0quTGJ/AXRgrrEbl1AKd26cpt
RNPnZzTz2aB4yC1cb0tr41HLu4m+FYbIy8/n0FxW94lk6gXpB/cwAKSS0CKYH+7y
FVQXzRgIyEIpB5GhzMAq/IG+Mu3+p/DC37IejJQGZRwpQNzm9xGER0nPJFaFZAMu
LTrKiu7I31QYNMVW1M7MXNj+NyhIGlJUsLq1vRXv2Z12BLl6p2JYM2JaiCBz62V/
+2gTeEafK9e+IpoTERSW0bueAtYlwIrwsWBwSk1M+WbyxKnQOsu6clSiLjMdMXIW
gIWlnIQfw4apVD5LvbfZA8aLooXxO22VDibNCC6F6Yivt9t7S8JdpJMXptXlqLLL
pEpaQk/7kXmLob40sQa++hY9YJh0EBtOP3EVYtvsIZ2sVF9NBN9LKnUD+4/v1JYA
jbGHUDCErvZk8qkHYPj9l6IC8Z7rdFSMc6Rl6j4ODYxbUL/zL3rdG3yNLtLGfVqO
nZUQkwvTNnmJt52Y6mkJevgDfKWKfcVvcDpoTj2aUmUpmazPyA1M6eqGDraD7efw
Gu7WrxbGNBEYIVCEjEePz+ec673wmMMmsfr35MU4GEZ+MCWWKinkFYf+lR5cE7wB
kUiBtxtgKLj+s7qOLpvuDQuNCUoh9EW1EPNVGef6Eyu0mZELIxvavIfU1i2vSnWN
j307c8dcsgnpKIYNsJK5Pj31dVsusUyGLKSR0zU6lY0hq87j+bIItwwavnjDoDtr
EqDkhSIQQfEfyndyD3UBSPGYntQJdTXh3q01/VZqDdy2e/o8FHTWJTg6rlrJFIxA
NCP4Csom6IrzF7rvJQBRgTz8kH7Nl1NjMoHxsFgV4KR14QwHmpdhJrfOoTxBSE0g
slF3eV0INNOH5wjXm0PrUcbEqpF8BqYkFoI2Dgti7UOHTU8OB0HuyQ9jc/Is9oCe
qsujaLTCj1ojvvmqF01LS3H6osKjkoyVGA51RiljFhPn+sxDmd3hYzwONIA2UKtG
/wSV7fimkblQov66vrcuLAsENocvxrt9cNaFVYKx7XRjrIM6ICaZh9086GD4f+Wr
Q98Xpxke5weV9upX9z/InC4FQnNP9biw/q2hAqxicyDF7a8cyVe/xkLEQfOQhYPf
ooCx1Mf2eR8OG8T7O/tkaWQFUu20J6I4GqLL4gFklK6Sjezy19ejPgeJbftWdQpv
xzZNORTqZtfAbEgl/ydywsMSx3RElloyWVm/BEOpipk6YQUHfjuNYr+7Ho6MumDP
URDqeDn3X/m6Xkj+NxmxaBk9ep17Wtv0NXlcwLeaouEp8+l6MpxFXG2fsqX2Mg0g
m+fK+3pX5NWG/uaZLfUqVMAT2PRsZXk/l3c79tJVe+Khp0w5qVkAj7bz80Ak8ZcA
i/plfHskobZMzDwlXcYwdQQMNXoGT+aRhHzD0t6j7rcfVvTfPVzESz96KWe/Wq07
QabvwWA+foOkwN9fGT4+sQ5yLkcL4g5FxbFXPzbv/UvfswljGmOHGkYV6w/aGDqJ
srXrTV991DWrh4SDb/gpwG+lOJZiDNmB/Npo9M7d8NOHYp9uPIBELisDZdZ9JKwE
Lx+fz5vWmd9zB3jrhoA+0zzP9sx8zlDxscGS1SLsEGH89Aig/9kBt8KP9C2QX7+6
uvCEQc73cALBxlxdrRpn1KniRspkL74iCoF5LzPV66bZOP9fZa4VLxgTxkRKmbmU
RiQFkpM/6ZNV50irBXNam6RSweQELSEqpgkMjNJKNt9ZLWWOzUmYMO1GwBoLixFn
yPagXP1IkRvVqp/Qri6kifZ8YoUptli2+4/f30Zy8blGBAb5BekvXJvu0sc4bxR9
DCrww0OQcn1kCv5ybOl1Xr02a9PQ/zPgkMT37bcQdzFlWy+PzixVM2mLOir58Q/e
PAZerBSLuXiiI39HBlnhWMfIFui4UJa6ZqynKTRfNqqltlww0bOUskfKep9MNJJ4
o9TyQfDupTvsxnkLiIC65OfmWv5NzpK+l1dhktVzhHOZF9YgbRk81EqwJSnGFpiq
fagKL55FFYX1LkmV97C8tJoul3Yq39FGxq6n9aDpoo0oSXYhd2XVyOL3vQrqzHuB
NvI8dPTh+954MdDkRMG1BAU4M+T570zgMd0M4gXrQFGzXGl/sTBKqvu4t4Knf7P2
xQ0H1q6kwTDwVvh7vR7RN0T60EGoAxVUQJ/p03DN4s87bzQB7I329bUHuWC30yW2
OpPWspwDh/61rADzU6MLfm1r8tAPmja8lAU6eYvs9yXQFWMQh5pMHOdhP6/hV8cj
77DOxaOZX7o1VHBoS7X3vq5u2h3Qbs3ydO/zUfItLfLXCXIDm9mY8SjDOnB1p2CX
awGcBwi9AvddVrL53TYHrtRjHTcyIanWNnQ9sMhhnfxU8tKkOndpNu3gQAZ6VnUr
+8kS0xCwYfdqf7m9oSVuYjXGthlo/iNlQXDFfxtqpgxcS3G0ZSZAx8K14QLIj82p
udNeYFqvnOtgcldkv36hwINKN5CGa5Nmnh0bcErbxxrhySf/qjP6qaN8mwB5RI+V
82UpiG2tdkN5szZrt68ZCeypJsIAa0vwLYcWRDa/ivahEdnyeAOhDgdemjDhO2PS
l43N/ciMf2ElVJmhXotKadgF4nZHobaRe49gT5Gb4XgApJ9dX7MTyqGbMzjBqRWL
MCcCOn1TRMZm/tC8ybadhlHYcL0E3CdOdycQPJyi+ia0A4xWRIPVdidIYsoPf4s3
eaHHmWRpBJtkKJQ9d0eO5XM0kb9/gheJxoFLQG23SNYQ8guPGqVb2UrKD0nzgS5V
L6n6sFDr63bvlgSA9vvZawwf6ZWZZHktRzMhJ4IfncccYR3S4ZWM7eH9lOM8kKdY
TvyE8D3XxB3BLzOmf5I09w33PuPyc4rFS/mLTTU6pDaGXfKtVOqZfRspUvxGptuP
Lr8fcp/+6flyQ27DPGYI9h1p+hftaRMWZcCYGFNHs4G8IzPPsQLMzn8U3aSNHhPo
7nUsen6qaNZSnNeH8kWoeMH3YlHxiaR+s2/ZKSIzq+mJZC4o2IHHGATFTwWdl8k9
mQ1kuIKTSeSC8CubebGYFJAiiuYXAHG/hFUDlOxW72YoZ9mrAN1PrERBM5qZd+Xz
IztzW8sGdNACHY5knhdjAO4X7k6uXerjiTSFT9AWDtW3JvFaMKIHTb9LVuQteVPV
osFV8+K1Wn71XEe2E3fp92Eurvfo0mTwEeuWnLaBr+8TkIADCamIg+BcxqxsHuI/
ELuY9GbRFuYo+LHlDPUTF8U5d0idNbXoSQVZYFB7GtycyRcYeW6j6dUu2U14Ja/c
HVa4CJpQVGAbMjNWZ7vSc3XSErXnDKVXFFVl3wYcnSzlIiwxQZTu1mFy/vix8nua
y/gclu2ZAO3cq4Thz8+/yzBIuoTsmJuZgrl8J1pj34ELDEUCnyedStJN0TQqg6Wc
ci2ikQV7xwx+qxa6GzfrWwTWFDcdE+WLsvReWaTAwJSwLw0JAPx7NMAJxlfAHpwB
Nce64/qs4CTMimGWut17kLTOGsuNna2g1c2KshqBkj9OWCNq5KXybGt8/VWW3cTj
azSVeIxE1kjL5G1+7We++gk4l+rCWhDNb7+4FuM8UbP4a5ush2+hRfbEGw6NMciR
hCF9q7k4RiL1pt1Ev1x8mhYwH+QMBKtKJXspPrz0TAbq9aNiL791m5Yw6ynEjzkF
6itTpGfN1eLe6AmUmgzMGpxrTl1/mpID9QC4/9reQPFpwXF3I/z3ASJkFX56zK3g
/6lCiWHGXEFA5gP+6hmVS2P9JR1bX6oReUBVWt07PzJGEg9yufWuhMEYz2ZAbFgQ
+Z6bZC012+ODz3xLe0Vm+Qh4xsqDJy/wZeA5sROIUzWPkyEXt3ywrWzf/qsRJQR6
XR3cMzDN8HYHqMAE3hDSOL1HQolgFl+8qH9HOu6LztGPJxVWOrrMdWu2gAqsYkU1
0ThswJUkyh/97Hp35kqLjq00AYj9G/bwT2B5CjvIOjJemibLmbPBDs0wwG9UY1k5
C6DlnwKxasmKL186gsfS3xO3zSm6eUR56yZQtIGnPTCyOfNXVb8mYQXUgirEoqzt
z1aRoy8XCOAPL7iK/qdAzmsonX4NguE66zk/INk7dEt12ehTdImh6rEOxZnn8qQV
VY5ZWaDeHnLfDc+UgXCqz1wsfiKlJxh4mBSwgAp3vJQrGC59mQSyNiZsmBtTuVje
4YrA9OYCkA3mQ+nBX+OMFLOI5b1Mt26VzoI70jHWz0orBMH73P0rbZp4ZHeibVS4
UK2hIJ4Rel41rvXufnbTulgLTwxjYSHyXicd+beMhox0ysUX11pVu8g6fWkpfuPa
6puL0p9TOatovMc35Jk5WCBUSaGoTsZO212cS1xJHBbnyvfxjhFd99LtdbzF2wtu
FDabnGiij1uSgG6qCBZFm4Dg5UzwmADDPUzHNd3zfm+Q4++9MCxt4IKAoYvdnEOM
Xpp8tzVehUcr4AJD69vUFFubXwoHNZexB0o62COnnPagYNAq5c2BGIvwTzJxfCZ0
RMDhYIm2ouWe9pjFioy0Nbcahgx9Z8Hx989IAyGk75h86FA2N3Mc3va2snaPkaJL
W1oYe8O4F+EjvIEgB6S1Cv5eEhYdTkGpWP5gLM0LjHVgDF9A8y4hNgR8T38aQiHO
9PE32EeCjoVI+9Egs59v3QeIlEJrrNjjIE7DzBM2x9pK2PtyXsjXz4pf9twXIexZ
tZ2QVyJESUQcN2ALG53lDzA+Zt7yrsbDx2R84Ag8ATrhYleDnKUVaRE/5bNFv7gH
HKS4+7QpkaJNdj4ZaQyfgnNSMfbRR1AKV9yfTJwltOEroCD2qecY5OcME1fRaJnW
ubGgNRP2SClhSHUXN5sicvQMmkFQjdv/Gti2T0osJQpGHgtoqNlZT1m73mskv0++
3PAaoX0RLxzQi+6ZhD2sEsIiJsCmxV13VS75t0FgQPPtzdIOfcatCLw+OQsRZWPi
I4PIS47LOz30o6Eltm7rmZYtQqbRqL+fOIiksMjkzpEqu8GOxokzoHB9LTeI6Zib
KrbWmn+hBU+/kLoyVR6A5u4wp7W7NTbiUG18PHgiT9Yo6gYT9pYuzp0wS/4NwXBr
iN3N0HZGk4dYeoQN1omHgVFHHlByC6KewMzGUiyND59lHF9JZJuuSMtAURmvOwCN
xg8r1xJgdH6Jsgw15vwp/wZbRd/vDg/ZyED4t843LVB/symth3JFMOCyl/raI04s
gO58dn6tBMn8Lh/OyKQuLcqDHEqkclSvmpm5nKFHgdSfIzfOhxDlgtn6PWEWrBQK
qaivnoqr7S5h2v4GF6rqj5x22zpomeSTXp2nM1QcSdJzfQeYWV8IndPJrwpJoFma
QGJcLk4RUf5ZljW7hSJtrtLOUjHfjRxbitHWIve9cST5AiPaX9fenLOtvKjyWoMS
Qr8x5r8//NLnVMwDvhUH60i2g1KWtI/J30mOGq/ydO718cvU3+rnSRgZsBZmshTB
86mqPGGpu1Km6XKdzAdaFjlEfhPI8m6s90IQIw+7eJvjP0Sq7wfdlyKTiQbsHLY7
QyOwBWWD3zZZl4TjyDm5RXjGDHR9bRs3hO+11zQGyQn+C+COG5o6w3/M2ZjOq3lm
E7Ck/4RrWf9pC/TzKuq5U2jGiKDigdVpPE7r/h92nrHv7DYLeRqXA2A4zGjeMTi9
+N1EMQRy/701JYWpQszx+0kBSvHfLT0WoNsTa9sjFbSHYkEf5x0dTrYpl7pegN4/
hs3qSJvaQQN2U3vvUcmu7WZMc/fUfGJxLvAgUM8unCVjKm699HGQYEkE4oyRETlV
MUIf2LXj5MYBvUzyV4pfjh25Mzoh6bJ5MTIo6F0+BjBFyUgJkfsrPw99P+ICh5CQ
sQ4vukOnZTdxmHSzP9/VQaUSWBXNPwfTseW3+hcCD5H8n1LhmrWy/PLtJk4L4Kif
hvqLStXNUGrh3BSVyOyhTfAtY9pyAKW669a4UkSkgdlmL9OLRODzrXFVfofxTf4k
Kk9w20jrA5yo8ruTOZ3zs/yBt9DbBfbcYkh+5iFPtjA+VCTUFylilP8AAvHQTE9U
SgKstJ5ehATkB8uxPJs8/qDICME2Sj1WjxPInVHRHUs0B51IXO/ABcdOn7VxasMO
WSTv73xnw+ouQtf6ugK9CokZ3Npw7FejND6pniAqf3sZ/7piFyrNdehrQ6lUJrQO
9Uzzbkp+wJxnf0pbCcjwx8eFsfOtPrKl59jZENXozSO3I2LQDNh59YZoq99g1Efb
JB9d15tMYyMDaXtxPy1iXTuSMt1yAls3pHD2qzsAYmjCi1NKbfgOnsEf8uLKl4p5
/FjvwhOtYJxqlz2yLVtd+ek+FQLoM/hL1pLkiw1MYR78dhpOB9F8PJEv7lw9+nFj
Mc5loihUsXbfrNiM65Dolu+Knh7UJgIYER0PNyVcSww6K1EJJZdS81zYiVr4w5xG
aSL03MhcDj0mRrd1s3u6exGM/UKRFusTuorKj0z2LCg+vAAlHv+R8hQCdpuTvof1
EWE4I5z/Ux9aQCRuAmXBY7lwRb0BMfOKBXV2iUQsKoe7MSguB2q8K53KnBqOMYNH
wlCwuBUoVgOy8fCTINdIdJcIuFYftzmIQ+uEgqyQJTiCY1FOWol4zfMF07kHi7Fc
qY42HdrFCs9BJk7kerA6ZEF2Zd7s09Wnxn6izyHNJY3aPwDJX5PrYoEnJKRMD65w
AD4CSzJXmnVRE36eHWSSeEM5HtWW9S9rWcXd6W3o8T4t/3bheI92wnWvzH84n4zs
CLiqTCSlwoVHpPh0ylOJLdhwUZuGl3/dBvpMM7yAbv3sn3O7OlA1R4iXJ5qkTrmH
ozp0EhXr3oJ7VlTHkcpDpZ1B7VYYekiePlV6qNgadBJsmZon9727U1Mpl7jim7bv
XtfV87nQHb3RghZf9uWS6gFOOjK7YsgPXhH7GQqKVsu7g8T7fTCwqY3RRrwyBrrC
lNrfv8lsQ7e/cAstVYbAzsRf0hLml7EzbHQxOJKXN5gLhbW56fbJWgDC81tlwjO1
KwJnpvsDqV87a8gpBW8rbMtCZN9ljyvr2uhd7iKT1/N/XpPaPxXYj+W75ChMBion
dXM+5WH5tfDMIMEfoKC8aRLEaibURE5avr4SmGdTihCHceAAtGadbHIaNYqcv9bo
Im+PUxpnQTSTpHwN9skRMZbeABdhE5cbDyfhB/Pp1juPcAHfeEoNwTKXYveqs8x3
QMx6jB0JIq6Uwjfe1CGhuFItgB4T+CPDmCCQzM1EBhTOyDtSSALQTSBcGp5oh9Zv
XrUWKzVk7k6n5uiJpPd4XX4imuH7joThCyYThLL5FIZeLRsSQ78SU9jCVGWyUdZ/
uloi10CzlvXS66FrBOBhnSNtplRoBA1mARzHe9La2FzltOwAE2xbFgq8ER8/DD4v
IZcr8dHBFF2B77YfkNxfByUHvTr/wgT0wEzIPYNt5W6zymoHShHHsCd6mlrwJDp1
2eHaI0wu8LwgqmwPePObXmD9Ek3pPhdPYB5fALCX3+Q4iYr7bf049uKif+cuJYiy
VCltu27sqzCXk/Ipkx7bgxgcQ7pEvOpBhV7yeNiNPT4jg2pS5UBW3oQpCBtsQ8Jb
YIo+j5aFFQvWDpOHAfCpFy1ZYIuqvwyHFi1lGX4KA0BEzC2h553TmCJmWlt+gYR4
axXotYaAytRjLGvOESOaBtih0fyH4hBVeUMeaJBP5T7TZRYwRslxyz/uyUkn1t7I
SYOUm6GNFZ6aFaBs3qRdznYJfiNWntDWiu6zzJU49kf5DVlXvbJp8pZyE96qQw1a
ry2rCgRoia8dcivwFSsbd5IfkQ+SHvw0Ios6RyaM1qSdM1ZDeT/KY+DHctdVWr7Y
fxFm7qoTOApQ48UQjfBDmX13AVDRVQvPeHtkZDPJ23HlLwCITF4HPSXqIePzqFU7
nBwKw59h23vdDVn4xcxCXFqddY+JAgdN8AyTXfVkUog0x7EC2o0lwBH5qp6+wU+H
V1JOKaUHFNeGWaywpIS9MgbhDQrKCBFKsBLWHOZTZBV9IdiHQVd3Veg+sxWKbvDE
fQ8sJBJ39hWCm27k8mVIXiLOvTeN5dD5SKuLO3S9iD3utDZyK6cZy8qupsz72wG1
B6CFoBuz1hFZpLOJRfoy0TZ8cfK8WQGmWqXlCAdcRlJZAYR7Z1YcKhhl00vF8qON
OQgWXc6Flhmb8F8o5WA6wUedf6FnwYvBs38CKeWMcJUSXUYGu3JD+5C5YRdeOEkD
DRCuKSKITDocMdo4YRHzJOuEj0BLRkPfX0Ev7Yn7RlD+MZ5122HANRvisZuu/bxY
smUrQoTV7h7ze+E25rBJYpw/wrUfjniuvWhWpiFJJheB+R5T/fZo56M9ObATy/jK
7y32TFL9dGYksBNuQ0whQHFBZJznUNicY4bI9rQ/cT9sha2ZskVobMMlqjvZt540
k65b1Wrm655lbx+nfo4YMsKfrGwyrIIlIQgqgNrSkxfzjMTTVfsdgMhWm2efSG5s
V1CELzK4fmwvAuqCY5nWHxMCh2ZgSQlw4YuO9BfNtIt0y0rgJpVutOxL911xGw3z
r/I7DS6VvgnkGrCAbsiaEkU1g56GwbdSlXiJ0iagvpbYtuGGKDStillyfuftIFY2
Htw7IMtW0rVtT+VqUvZWqjaDNCuQlFO1SM1Cc+VyGEqrwooRaU6sGVxNH5oFj2j0
B2Jq2u8nmHMsz8Ba+liGG0KKSlhFA2NdVcjw3SbgLeRHwyaUc+/rUF4IM1I1r9nX
OyTEPwmQVHVlFKMop/0AkoH0LI/RzEXn29scYQX/TCLX4RSf5qOAS4fisYeLkfvm
D5YX8Zq2/xdP1/pVeI8kougTO+CMno0fMpflmmTEgoP49vdycN08oXfHUkKqFuAE
vEhBJdmoFI4SvvT/uXOnzy2CqLyE9kcLotSDcrGGJm9XYQXqlf5ahyaAyvFsvL8H
6jsUqKs27wYprQaRyxJgKtuD10dSShCXWRTW7Fp0zfWShEl0DC+gSopqnCkgsmx9
wEw1XjWvG7l1k7IsQNYN0Lmsrj9kDzDJx98LuOCnZhpG2+Imhprro1iNHL/kXI2q
axBVwjURxWCYIJrduRSDKISHIPGTOvwHuoIyWX/dJcATN5C5zza2VZ4qZd77Favm
p5KaSmbO6ARa/BP6zVuSlEyVIyD+82hHOMYmqKg73THoVFVWPx7aqKmucjtUI0Pl
5i9t1ykxnRDolYIZ4zCJwpg2Ni1VIzmOLwfm2bnKpM7TE/5ORq4rpLBb0ulMBvEa
K96yA/6SoTFBxJkyebd3pzD6TwxoEC8uSkciA3awniUOtb5zSW3wfTiu1pMig1Xy
89ACynfpU+6jwLDaCBWTaDTTO/xqzVtCPkbWVQq0t4LWrFGOXfXYvB7cal/CdR02
ZqnCOv0DIttozlpQ0SOU9tXI1umtimS5Dyoyz1ITD2OlBuM97lMO/aogfkiknSGK
79Bk0OBKWOX2h1NP3ooKgYgjWuUA9VleD6FAuVQRXZI85Dj4fLEpZv2tvqZRFw0f
IKvUaLrn2A5/PMgsEqDzP//bMzHSBaR4Ml0GFMsUAF7a3ogmi3H0gBPW3f+q/WMj
yc0KJBO/DKaCafRc1Z23IuIHxOmSWSp5T/oJspPFw29e03luzNieWSB2+OX+Nigd
U6NAGG3J71D5X9dqoabsYxVFV8YlLKR7aQtJYmSCJyOwXkN5mG2166H2fNbypRte
M2mjDIrhhUPQKO3vVRHHBoO98AjzRJqgA/64GqXvrIEXckL1X73u5M4Qvc0oLhG+
Nv08YGHZtlyy2F1aTNGsTHLN3MCKsjZSnVR+g86ZW8cshf5vueMD93G50hdpUcc/
RnmwB5B5KMGQ4H7JAHH1agvlPYsfH5xPHwVq0O3naNF7RS3gxqKXRGykOLJI+cFa
yeT1ha3IcSNXmBgt4czhDC4G6qSAMzGgeFcfvkXzrawfJUeciZ0AovHMGJdlOFy6
P+orZNMrqdEJeNnDrxKEYIs+ktT364ygNJNNGWYH5OBYIRA1lO4dgVzxiqFUyIiu
GBwL0hAEIGlQV6aMW1UT00yJcbV65ArerutKjMbk2pBCa9ZPQ+e3Grp7izPFF4MI
+qy7yGu9CrdegaDY5c7PNgOB0FoIpsrzMMZx6v3vEZNbVpMkChyTq5YvF1Kmr62A
xQrg4PXG/VOw/dcoOMoCjofLGn85pj2k9Bs2H0ShXHB6finlHSNGNCbUrkqwZ7PQ
H2YSa8A1uHIduA22JYHEiqTDU3A64D9+zv6id/qzRgYG2/dUajUXRF6jaWxzqHoU
TEmQ0im3RYHG/wUL/ZZbwreHtRpl/iauuVWnxWnOcXINxLsKlgbbY+wTd1P7UE6/
g7nCLc6QD9ADYXgiyiIMzMh5rdOwkpGJhZCmeGRfgcz7o/YjaMweXhsmMnoEJone
32Z9fcyue/qlSvJUQxNa1bXoKZdqDVzWGq7hDHLa0DfrBqo6sVof+FbhWmrIOUmD
gthPGwO9mSDK+LDZi+3AfJbdHcSG1zpPZNiPUKxe4dF8NT1cEAlXLc5n8QG14ing
Env64QuPgCpjvO1HjnJp9GtAvQOcwFnMVL6LaOqLTn80iS6BhyMcxqfDcC49JD6z
qtGnCuKTQ3y9qO2cjRVHh0Bdu+QAsBaj/FN+buoUo1OQqYQeHcDmsYZcNNEogHx3
iqPPudy+Lsgv5ajmJYxAG9x2uM81GRWeXwk+SSlm47s9MvFR7+AbM3KVMgyylAbS
/RgCG+CedyzltCMK4SyS0OqLQbKAguN1AIRQObB0PLlUk5AbEjhyEat8XKUVCX7V
pp9ExI7xRN/jqV3nK9KBOlhJdYEqGSCPoMdcZ3MpPo/T7XDQgw3h+3Sye174SDRi
4WBi0X8hzLzzumeUjiroyNHyDJ+qYEsrO+ZsU7de6kxjgC6jg2t6OgbxCUkteOfy
BHY8qmSwUwYWFPOl568aLBDUW1cfePqjERJtu4xpms8seIBmpmcOiIqjqI79lDMJ
+gToDZcXwrKDPPGir8OUrtyHfvRONWG5VcLmuOa1AyqcowM3a0SAZaIby79zAua/
6i+aHWnQM9RI69t24GIt4L5smNKbbR/fg+kxjqOAJ4f/cGG9EOu4j8WKKkI+AB35
p10TZ+jBj3u4rMqe4iLiz4zBh/ywJrQLzqXr/ebJaalHlZ+iUwFjmJVs6IpAUVk+
WrUpEHAeX8lG41Ixie1A5/PHdVOybrs4XXdSHG3WnsxnXvnpuXEccJhW5OeqZXxX
QbV+CnUKegrJV3XRMYxuNw3XZKJAOwRV+M9DS/jtCaiCKnn8qLkJwsvNugT/XD1A
1BzBnkAIaMVC8gyyWzUbhAsYDbVDijP5z4qkORd5kL4UOFdJBuhPDuJXbvkVIvH7
T2asgnwzPXFPsQ25eJg8DCuSlXJZC0+1RFIAuIIA2i4zBrX4rhykrJbLbK9ksR+N
qkhTgH2odHrEWd/RoRjDrHjJK8+3FAZ0G6HZORCTXejJkOKn7M5WBqH8p2mEFAFt
+f7tL0iWst0yQeFB/d4T2w/6SgwHCtKIj540PGGApYCZ4tyR696S0Lw/K2FUHRLU
rfVHLU/zYoeZmBsArgzUnkD5Pc2DKjk4QOdzpvXG4UBmMC1pNEjSazHxXX53HAiK
lRN1MyGDa52Xwfuvv6cqna+2cG+GbBKAV9tuhR7XZEQhwK7za1ikBmmxASUxB6Zq
7zEiLzEGWbJCyUlY9CbbUfq7LDKsLxTjVuwqt2woIgwwHar4fdqr7CmNDZi9gbnX
0C+tFwPc339RAqLDa6DcbdKgMS3Zy2lt/Uk0t1/uSORU9tP9hrGQ0NKBxU2nNC7Z
TZfblU/X1xi0M/auel4r6oI3B8WS4ZfVJmUJoJ758SwvCha6iV+0JkGRTrNUlllA
P2fgO2Vd5TYeAkIdjDAISBxTQrRDugp4buTOYYH7+81BjLDiea8fa4zdsc8UKYBV
qNajTdIQTtRMWbAGtZIN31iRMa9FdD06l4dgUVIRve6k5M+4MrWJ67/jZpduwrEK
bTviW+HCKTg3urYNXKzrHoS/5fDe44+/gKkcot9o/XqHDwbhXNyGg8Y0btUnkQOX
m6qghr0poIcXEfPfes8f/Ne8Vt4cIL1lebHobOkyAryew92qcn74QVoSBitGZ8IJ
g8a/fmQKaiHI5fo/GJ9L9bi6xOCvfK/23ssHu/KoU9NDEJP9wdk8rhgqiSG7gTrH
4ldU+uytLAUcxYG7TFXoMiTaLpZpfuhu+Mg59UZyPnpFBgV2nTqQcSXXNDMuNblv
aqw9gCGFTImQxkvWm8j6SaC77KBPyURs0M99Epfqe/+yKCmgdyH559ilpQP+S3ba
bSPCRs5pzwbFruUhgjUD9fSInw5Psr0jRwh4ohL+EwvqzZ1TQw6twP9H2jgFpmDS
ARZqOhhTHhc/ifKBfx3IrJ7mAEwAHt/zP1UFwOEWWwOiNjwhm8fbB2cz0h+MGqW2
89fo/BmeF6f6FsLi8IYQAc5AA33+cBWI8OysQKDjR3OLrSUv2jwVPThPkHllwLFR
2QtTBY9tXkw5viyCK8KVBcMJtUqgRHVVPAbUu+NPQIlkwBGbJKMHXWP+EPP7nSAc
NkPSlzaGVKZMrqzJ2QOrWScXfaFfWLSVtYD2gsyH8sbd+SZEt5taM+Z+9zGJLdGa
0/Qi1rVf+LnDJiuCk6aGClJcQkBmFSC31feGiRF4CXfea9ZUJOFxDIP3Nq6JhOi5
VlQNcl4JiIYPhX2clqo9AweRGgW6sAhSCnJRgynHH9xHvhHDsRW6A/9hDBWrTvxZ
Vdva2CrB66zOt5zu5EbKBT49qnQXwdxCLn2pL7qaXjMXydIIw3ecvZTEpyDx5Uo0
rKiCGeC4g8D6j20ERpcIAbiqTfeXlZ5zqKSuDjxzufUizZsjFyvS8lf+Ysh5avDa
sfe0VNoNjxVqdcRl+BTP2zy8MskScP8i2Jw31z9N3dYH5+xF9/NwzeXhsImBujy6
OtBhbnAB5QL3yN6clpG3nazYCLu8nA66FCD5kfBpmCidc5tC/qZrKAYcNyQOG76p
wuVOKTz3nWi+heHe+ainEQm8UtJDr5RM+rEfepLgW0CddX670t/HcKLkl7ccSZ+W
uHJFbwYx6zy3PeY2zWce1pzbJ6cgmBFDYKUSaYlyVx7ys8V2xvhCY+QSJJ0VG/yi
QiyHWK6Ur3aWfDzL3biKyFsjYTqHKUwnxfoqpWDsBhzYal0ePsXaLgoRQDFbJ6eu
DlHakcq/7vFTWVwu3N7aCR7jE+IaC6DOT7FWgqSMtDMUEKSCmyYJb+Zzo7RoNZBD
c30xMinp2HPAwXIoMpROPMfIfMEh/mmoVWB2jdtbVjdRPgk7itK+VAeAkjNP9EPO
HHq0n1jRs0eruKGY+lsUGdbJRtXGce8VOvvOcIr6AjNN8Fzhl6EwKwJD9A5Ldq53
/uiYcA0yS0sy3a0Dja2p2Ub9VbAqWBOf6NOoCI7uSuONFH2VUcAAsNeHLdFzE6wn
2L554fWhuxKUBX051efp7TmIp85AibyESvEJGYWGnWZVUQyVGF4yfQ2XHNxoNQ/e
oPGoKxwdazwdugjOSQC5ntTE/S7/qPN2vf6GMwCwuHzInzUcZAm+ek/DizIFsJYn
bnvy48Asd3yZE1OLNfPlAWIZvB8PmUvUZb9iiVu5ejOZhSLZGHW+5ycgioAo5WF9
NmNmagHfEfkwCTvK/oE2v1JFowYu5Qer2tarYSKmZhwFeGj0oBiDSMRvXLWgISU7
yri/KsO/HocOcfHIMjQ47xCCW5BvzWwOZXg9WfWrB2BZdPLXSK0Wqz6QLwf0AYRu
Mgsrqz9snTknE99HWo6/8bMZOhpqkwQbH+hvys4lxADzFTFLF/dKlpEG22a1BKg3
U32qbZ0rzmMNLM47I2mjDwplGDOXlzhXm8CVG8fYz8MQf+wVLmQxhhhPmvy7u3bR
VPrLKC/X/y62KFTDlhg8ihtDeywaJbovWPUcOnKbhwt5yW9lwNkNFxZQZFEJOK7G
OjKg0wgxAItwb7DOzZWJEVDO0SfpNtd6Viqgq4PuyW59iGZ2tSgFMg5C+rf39DGZ
aQUncu1+d51kYItQHqdVZDebSE+YwGhgc0WILGvKc4DuPoSqQM9flfOgIVlzkR+E
MRyECz5aGngcQAER+rPJAdnL84GpYUz3OEM4Qb3g/rp2JL2X2fqjHzjCnm3Q/Avf
wMY2YPO9UHQHVJQRHF2o/pheT/Fs4k1ksF4S7t+MWc/iOj3/8QE367vI75VaX12w
7WoCpUnz1WPgTUD6AL5Q+2/kD096NtxpNCiMD/namaQfhuy1EVcZqVrj0pLMPySH
ZO6DlSaYn2qG5odD4P9FLcCgtGQmXbiQxU+UzAHj75bhacbl43KVS9fBMVNjILCS
1Og3OCMGc3BNzXWFGarSv8HEVw37MNz9iv5sqWiOlZux0pYVIDAfoYt+Jnllvhhf
cC1OshdMxTEQX3I2tql8HWEwwiwkMAC+K7BR/X74FswLQ7S0IvbSl209/SG4GjLP
SmygxvnB7cdVDT68XtKR7jc7X0vsRT74F2yBOCTAS1JzTfpypTO1YcibEFR7LOVm
Q1F/KhZVqcdkuPbjZRl2TPpX1M7YjIIVKptc9ues7piWcYriHbA7RE/A7h5WgRhU
dPC92RjmYawi7rc+HwDya3eDMsTSSiwqpa9CDMgIY1gTlVt+6+98JVBxVmGknkI3
WnAQrZersntHCZ4rns2WUhpeNrCkDsX1ldVuQcFVTISKe9dRODL7xBfgHHTincgo
JIjd1kaaJ5x9/7i0qrKboIb7u5lUlXiehdYr5BZyMrECKMzAtVWt2f1q3c35jXOs
1Csu8UIXM8WVUnrkN0HPQvI7begChofD91kPnJXDRw1Yydj5evhxqYNu6/Nz5UJe
+8Evwg5797w95bEYGC4RgRGoCHiWP/rAdzaTqon6EN+mCx2U44q+E8586Q9SeIxZ
mhMeMHOXHgB+8N1JLvIBmk3C48kqNNBVYTCcT3bepR/ijYr0L1gkJHUzAnIQGKPw
hrkUFDjYyr4JcjkC+wxdbJHv5NE/UPUHUTHJQ7yCDz+8MfVMwhV7nThrcQYiy0rh
DXGQSyqzI6xlzYhrwE33rd4GwC6yv0yivawpV8jQwfez6/nSRWU/UrDSDEAu+uhe
Yw/eyxQBfijcQwYRq97DQJuNxDumZHSmcuyobB+eCEXWH2dv7hrXqOyd0oHiY1Nl
WTM0AKJ6evf4jSAoY1Ru7MIdMmdlwjWSFQO671bB2QdJd0CRGoi2kkpkzTYkFUfc
+8vTXEq30p2GU4sT8USP38lTjRrqDXSCUPgE3GMuWb6CjEcKXOtpAmZd2P+17Lja
YgMRC6aomYTL3q/vCKpYFFjHXB70EGpSTstv+d7qJriqttYkRMpoCpG0fGFSBB9z
qb7qNlgYSaJCbpOqApJ2aN4mKwrqI0bXcVM0IRRiJVIHupf1pz/OlX1nGd1PVaWg
jJA3+J8VuBEE0n8YVBRpnRRgAt8ibYmk0+NeH7ccR9UfIT+1ffCriPpOsDrFul6p
0PU0wl5sJmDHsCnFxw9V4b3hQHyN9IVyjnS7SOctNCbKKAjneFHKw2sYpGoxPlkF
mVSJ+gDaVlRXvLf8mPnQxq3gDGxse7yzZthKv1ulQ67tudaDN8dLjdtR7AWHysmZ
hLgkTQokhPI36EkCjy3lN4j191l6wxXOYq6xoWyI4ZFksIfhOS41KbAmxoJRz7+V
pVXgxEcyAaRRry/DKrviEkxUWwQXHdtcK7khqf2zVHnLJyj4blifgxQ68GMDi3yB
GEsaOO7Sek42Q2TQau689/NJMnHEBfMuY9Go3QXWspa1sQNCqnG3f59Odz1pb+NL
op7m6cLZnv0KbwQRGnA8ByEuwHo/JJokoYZbs3WnmeDIhb5In/Ipc6WCqZVvcVTs
yyK7NmLGWLuZU+ELj4S1GaAC3vIFYJQVShwbSqqyajExiUhVxaEOBCefIAbSzTU0
WlyVXBxAGHSgWSRcjAHT32JA6xlkdTw/NLTfyRoaCr9DMUDJUEM41NjrLOfYPsC/
boIx6pmoUy1WPPlYBTGqVndPGprOlAuUpdHyWTR9ZRnJ6tvnJtI2mu7Qqq3jbp2u
05nATfUkUf5wt2XjGV8hds7OPAGsZYBJ4uwGfexnRXCAk77Lo7cUDVrtjdqLw4sW
Siq585byRUEGJ1xjNeKMx52UahZumnQT6cAvd/nrn/Y6oWx/PbLDNrVETnUOug/s
kDdJ2FoIK095K9/8aSivzLia2KerwZBLxPNu+vZo8UJgu2jyq0nj6ZRkUuyZHQob
PrKhMBLjdRus0Z4IQrfo6mg3SQQSqZ3viGK5pZCdDE24r2KlrHRAjscUJpWQdj+s
pnCU/sBpCW/gmyN8UYun+44l4tgNBsbOaEhXyBYugmoauYjwZNqRUyWRUU7iJbDT
L6uzKZx29ZbfjziIu/My5ygmb+7jfcuB+1RJ6DTJPo7oHIFlfirxyzNw3kv/ZdtF
CLngevncd2DP9UX3l8vw44ldHgstmjHMS3KyJWO7jCJmKhEWDape3V+fEtxjd2Ls
WVY9Mx8EBynvhELYTxTdvJgFzqNaLLtPoY76e8rOOJaMNnv1OBhcsPFI3BnWneoA
jvDRJnRoH9x5tgzYa1j+V4tSnQsELwiN2HhUR60DG2WcWEAZm2WLRYeXqQBtFndh
efTgIuRGLhDem4VQ1HZh+VIuY3xSwjRGLXYH1GRv9XB1RCXDFk/NBvbpUFESzAQI
2KqdtQtI/ub2ShPC0lHwiLFg0JqBCXIIXcYHaZDaHyUlVjMsG6tansPfCLqzlBYR
67ihGxt3tSUIkwDhjlZm5bTs95qszgFxqm2RMOCERgc0N38wYJw+jsAr9AagFTMA
jUBYT5tak2QiDrsWXvflLdD4WKDDPV6va3/iYwBfQEnODUxeJjYVWuBQTzi3Io4p
OZt9mP5K2a3h5LyU65pLxgSpPCybZjr+IRNzj4DxGIC6Ik9tR7MIhxSV3sZfTMef
L3HmA91m0YPX1c8CaFxBM+ZFPbh4bRIRp9XUh85UvbaJesMxJO89zWA+UtPG6E5P
L1Xo/P1aruvdPSlCPgeU+S6Fkxo9vSHfnaMVaGo05a+BQYk9QOlzUi6vUCraTwoJ
eimSPxIQ3maUpBksbaIsfuoMQD7Px1iD2S1YLbyHqFlL0uuBrjuMqGWpv+pfcPTl
BLn1B4ERnxnpyFcBeT7bMDE/DyiBYVh4JVhEo42M2i0kaMq4H7k7OxiEw+nTmjMH
+s0ElQEC1xTGMkjXhXA29QcjYfq5ckhaPTrPRNDlO+kyXkUat8pFS/SzxpK8tRD4
gJwH1dyw3q4nCgYhJ+ne3B1aw01DL8kRT/cP2YhhbCfZsSSItdt1AViWJF4BHR0u
LJFo6x8NxcPJt6Ln+SjVecDzOFmw8husxEFvXm+iXWwlCXBN43Pmyr2l+stWwr88
g4YpVvDliA3bwnOLX0bwW7X58CZz+edQxEtR5J2JzpXn7qSJi9ULn4r+OTjcxJ5M
f6REvqxG2c16YXHe5likWjBQvrvjV9DGSrgOIgTjqF9wo7q/hZKEBPGQDFxMrRc4
qkprQNwt3DkcBSbgHvHjVvRz2W8g+eehIfKqVZ0F3nvfknqy34Wfa16M+5flo/Un
0buQgLo90aUrvAP8hkbnriqmo67nHebG+GYrt38OygWBqORe+OECzTuBwknjsi3Y
hRrkGXwi24VFlijLgx/V/ZPwZekJ9jiLlgxNcJnVz2NsxlKwPfycCkqmeBaIwI4a
5u+7fmIAFrF8iUxUBMvZDZiYCfRgd+zuax4UDAZHlHodQjGuCk87y/CQfBEV+S0s
wboYykJDyK4Nbbpa9tyP7PvOeAvEOPQ//Q1aPnXAqsebshbLJ1kc7Z/0v614/rCK
iQsgoQ/15ybeLXIEwABDBULukr/8JYPLlT+ggqmVA5hsrvrv1rnjwM5hE3sPzRjM
Gp1AsTIjIPb0D84qlslL0SC+6xbNISigq83hIeTsBzt3kvD2s9byHw4l9Zex/uwN
46ja2jYFkwk1NIFebHlkp/rSmYwm4ijH8IDkSEEGuFWJwJOSzAgEOzLqS0+NpAbu
2MXIAoqZZTRjzG0EX+8vMFqLUw+a+IiDbOzxMambp1MGGI0rHHIt4vy4DGziKLAB
RWk14jlgXAcfQekUoP3+RCcldOVbR166y/BU3xi/pqukpFV6GzG8vt+v9gKXmbTq
3jH8aSjKy0bUwoqbQubXi5xHSLRC4zYBodiUKVuekI7iJWHYCXDxSJqEAc7e0KWj
w4qao+dUDjaJ8P0RK9UfX/PRekiNp/v+nUmp7QPDlSXpdzCP10lVIAjNHJSYNcUc
JkCa44eeXPUBvNncQ/wzx4Amgjt8Usgy4ngIQfgzzoPljsrAM7vzk9Tzezo4VBVQ
lu7x2EJNdfl+W9CKoNNrwMtI1NWGiM0rXQe4dsGqgq80hnJAHD8aNroIJtrIqJrQ
UdJyOhdYntF1dv6dg30c7/PoFm90jO9OmC3wvi8gO4tN/WcAY3q+AXV9INGhMiqn
Dx/VT5P3lo2dYY0S5Dy5ODaZC/R0n642KkQxbspiinI4iiVYgxE91/tdRVnurVgq
11OqI3UghhEuAohXTKZtYnlYYLUW3nSH40MRg/L4BUOdUjzERV0+4+qWrQQ/Eg75
7afa+1pHet1wdgHBIYcIJ4E0fVRRFCeaqGKhDqtafh4LTGENO6TbpvMEhyI9fh+8
bsgPGL9Gg8KNuaP2n6ZEti5X8EISWv1FaANzbLsPyN+VMjkdG3p/hYd04N2c5JA4
twqlqvIKNN/swK7GIV3nzdVj/CZ1OUTqkVVFVzvQklh//jvZmLGVKmkTfUJjv9tN
0GBfau7ytb9u3hRWyxHcc09fHbiECcfRc8KoMVA0jhErOhtaYi6eIdYWYZHUsTPO
LL6bGKWdsoiPdCkwNtZ4Iyk2oe7X2rNUKYPjymM/mge1aMO8SDm7xEw2O3iZOtJ4
J9d+nkEJWRVkFGv2pgULBIorCccJVVX77mTCcfyE5eP/abn2qTPnewzBm83xeZXk
MiZysYQK0Ec7UYNPjrOzF2+MkngeRocadQbxv6k1dxwheEBEZi3DDfbqXuBH3Zra
s9+PLjqffGWOyCERwoYmKD5Jg5qyRj4R7NjugFnPADm+CkygU47ifnUJNGdkTwJX
A4OJwu/QXHCKJ7XN33hzESW6+Kex3GfZcv/evKdr9JpOvBIUqb8KvonCaPUYUviK
9m1U8ZJSK7qEzjIIBRHLOFcaYz7bY2+gMWJqm+3+NuImEBLcwsMGz31suuGrxahs
OsnzdsMGBzC6XPdi1H6ZYNNTSeiV1xWDMDxJCi9bCnKM+PgdYsp/0ZvWyCvQhfH4
luBpzdx0GBI8w/4/apdTFTOpgTzU8hO4hMf6bJN14qrOwEiakw5o8W4RgYqLLdpI
3NB41JVIhv8JVC4962yOWDhnta+dwhpSKGnjrbctWwc31yT+8cvEdBYrNBT5JQ0z
nT5AX+fRxcEdEESuhWsZ+na/eHYZLX5s05MInX8CWs+W6RvCEGCLa2fSu2IfpXs3
bDPKzDCyUMGuk0V7xv1lGMUEdJ0rz0Eik/ZX5aY1f4Eh2NzZ4FjGzoWz0xF3C2Df
LtDAjp/jRunazsdYS+dQ6pLsZHt/lfwWLfXaG51jRBbihwyFXYS1p5klWu+9vFGH
l9ExPH1KBRk/RKuhEUkO0qECpLGUoZWhw/VK173Vy3eZ/VBOtutIMe3nfSP4AjSn
wO0Mc2fl1ULZOXk+CU6X51x7xsnqmk3JpASy3mUNa1V0d4Rp0yHqKCKARlWeMZ7y
0JtJ9zlqqrWE4xAlZJLJ3OOk4X0xnFFGdZShtT/UkIEzIBiERt+z0xk35iakozkw
LprDpyAaVvG9Um2/54M4VkXQsDx1J2M5VKavh5I81PLd1rBDiY5KAg6lejaQXu3I
iWOa2U9g5wvKJuKB4BgIxCcJnu9K9xBtB3HLlOviihL+qfwQm9cpbC/YjOGZ3Lxk
BO67TJPB8a815ahVnjaMGVPGU4puNC19jGQZf8WtFqMxXoB7N75fCbWcQDtPGg0j
MFtmLI8oWZ6C+fEqITVktzUgyrU5q879bI2AcPH+emlQYmRGn3vDgQIRhGnQeCNg
DQnnarKPKgQ+z9nqg9q4OuDq4+w66ZQme1kU6okeb/Z69vLnhoSsqR1cOeOT3XHI
19BasJW5Y84+mQOYCQidSJ65BW1t2ULKR+/OGaqJuq8m4u84q8wsC+ASX9pjT1q2
1xIzxtN2+bfNSznx4sTITV5OUKbE4EczHA1KPp3EroXpam9USBvN+6faQqX69eey
qJgx4bmPDegXJ2/A6VCs8Ikgg9jplXr/YFiDlPAmjF6PB8HR0p3QTVfUMLD7Q3tE
AnRwj9dWYurkACukbKWgjgYiyeJunYerfFLEqEp2IUjIHjFmf3nnp066/LQXKHgp
MLeMLhYISZRW9Lw+yhsRoI2nS0Q0Z/qGdlYR8kZiM+LpHHr8NA817WaogBj4H/Yi
v27hBeu9UOlzPpdUAHxos7pBe8mPV9i/SVJDvgTk/cw4Y4SSuaHA88d4IJJGI0QQ
0YdGfYdRbRy/5I4JfFquOybYJN7HpNuaqoBZFQN1LQa96N2jJfg2x+cLK3jZAlLN
YGyIgkuR110Whof12vB8qKq1k62715YQOq9Dkail3LrzMfNvywI1/TjeI/WvK2gF
gl65ty5RG6XkWpB3uBH+8N2onwjAwbRRvRI676V2eb9zAMZCM0K8v1s4u+sAXod2
XdVBLFx4VgawclyGv62thA5cJTK2lO+i/2i1/WNb6f/3k6Kh0NB9MYUS5DpNokvy
vbZy5dCNZ7WWqRaBs1qNqz47GOm8HLXl1yrOIKTEgrZ8zHsAMU1UBRyYnXXwAFTS
OiL77vu6e//DAQhLATDkho9Jy0MmfqEuawg7QEqT+ReRi5EqbzYhHdybPQkTmw6M
gzv6utK5mapWtaPND3uqH7isuwPY32Znix5PA+8t3up/NhhaX05Tm9Xv243PDZKa
37c01FDNdUdhWYhyYNxe2qmC7OQSn+gvAPhK0RePCj44AJlIqkUIUXR8r/3qkhBO
9B6wtdQG/Wc839LcaDnTleuXFZlfqt2Z1Wuc2sf9dBlSwCB7PVDGQDWCCipNrYur
JzL8AXBo4nfqB93HQkqnyneBIOp2F7tlv2Dx75F67CmiGZiyqco1r0dOf1j+Mfzj
GxVLF0CilJJBzOWpLunO8hD0RkBchpPw09jVdhc1ncXJCa2HlPSiZ5Eel1LpMnHx
M6GUYbdekzAM0fggtz+oP5mQiNuEE0Csm2yZaYWgwLDPJEGJiY6gHFesodJZO5/H
i0yTu08ckXB72Q0Rn9wlfWXXCFMg1fNbfIeDrhPM3++N713/Nvr1s5y1tv5lHS/E
C06Gm/aoo2BXqqvYX9GXiG28IIy86kxQg/XWJsOIKCyIneqT6E702e8REAi4a75w
jtD5e3HcJm5OLtnhNcIEjIBXfgigD9+zCvTCkP1O7P/i8V9DxbiiRUP20nqGdjVW
l4WskWzLeO/TrG0wN/fcHT2EQK3La8OK2cpR9nRt1DoViFXh6GNBxrd6AnIsgZum
sCB+ieOGbQKBCOCjsZ06Oso2NazA/9C8qLR9APyZFpedqTXyWCEw0lP7grG/bMU1
ZN60ckuo+wXZ0NyUpQ3d4Z8mzuANFxBXT9EQHaeUvQSeib/4zdkYlBcoJfaEH+be
f6WKw5l1QkDSCbITER7MFOEJXGH6aBbWvm5a3b+lWG+PaGtyYYFMh5Ti6zXneNfT
G+6a+91pBDgLJWaclGOV9ovaKRmd9Buf0oC3Av8iIT+0f1+YtCD7+5FaQbHX+DFs
O8Ngua2FXMDw603/pgpLFRzVU6saklZjtI7SrL405OIqGqUwjTPZT+xuGhNDamVw
TaUFNFNm3dOKsFzLRVrq8VmplgczJ/IwyNBLRuVd2fGOnz+pHc+UfazmedPnYmjB
ZYx9qDrVqOmmBHtPxSrTeD1bwuxlhjv4U85vtz/YN5qGjNvSwGYXDQ9uwd8a5Q23
w5u1RNgyhyTlcdi+Xl3tlFRMSK8Z0fZw2E4RpLtZYMh3LtnS/Yz4YUxqM2D2Ani+
USGKrtheCYeZde8ZTYHv3Co2cpsyJUrwqxENV5uaNR+6TK+ujqHiYZoB9rS8PHZg
UvlDG6x2lCaPRUzXyhzUhtZKPWMmuyU9jB7muug7juJ4QbyCAC1hGu1CQtP/2cBB
sOtj5lawG/S2tynZAPSekSMzM3bqkA4/1FZoQGbDMO96kNORw11umn5OsyJLt2xN
DlFpaLIn37/WVz/JP7r451hWKkz3UwVBDyQmuGgiydfLSGQfx/+JKyqLfb5l93nZ
eQkgeEv4evclQVR7iXTogknkdHVwXSCDVwnpNqIM0VDicFwJQgbSiTTD5Kd2Un2f
yBqwHFvwe/wqhCBg5utdIXJ/K/7WN1TfLWVMJG2GBdkWABSKn+WQbbe6l4Qa5G4N
uQRmZmf7ErPBtJCWe1Hi7S3GbMJO5ltcc4ZWjVMBmiqx7eCLIE9TWNpa0puwVIy3
rjO0/RCY/0JdRQbo6vEtpKgJ5PiApj16CchZPpbbNtIQq/f0nczqOk43OTPoKUMt
XfWwXkp8+Mutz+u3ZqdpSuMWg0m1+1YJVxxFs1Euh/VA0HNKFqS6deLGyIUzgnTe
C914PPoMCNwUWrSFYNUjI+yyN7scCJAqMB/2SRMH/q/1F4VDNV1uUUKDQ1QwnBgK
Rj7Bdy4sy5bomdKGf2vfOjtLcrBQaJfvwKbtzLQt2xW65mTYarUUJOrZ7+WEZuTu
+sGTQHu+PQQ3m0O/EvaHtPzSZAVofN+yq7dHAWLv+jvHxPdpMLeon9VP7n2Vc5YF
/wD8KTwzbCeUEewiUeEECAlUdbPaqGpHq2OkV58xsXWO16Nm0nDg5A49Xfnt33sU
O3zamOYt5nk/F14IamOgX58q8LAauw6KEb4gv+DCZGIrYjPv8YVr9qAL4eeoGbMU
zC9hs9L8V+l6Rx9fTEH5lWdvx0/fgaCRpkUAieusoNlZUjd43ijUOYVxR/pKb3T7
c8AxAuMMw9z11A8hf6SjMER0+fI0FhMy6r3eny9VZ1Rfyu51BoVmZekQMpn3BZn/
ZPKXaKju/bLy2CmBuuZoW+NSesgbsG8OP0W/L4M6OWEvs8MnEFDN3iRzTEGVEeVk
7kVffbauFk3VA5xDhWSpTV440q89lLfOD+swdenqfWZh5vTbk/UbJKiM2TqhahtY
Hxmn6OrfNe6wKiKSG7J6IJ+31X0kuMwMe9jo9+F4eBCmu7KYS6JykeAUh1cKf/3+
8qhXfdbi6SpRTC6VhCvQR3Om8es1Vjy6g31sVtxdVS71YS1OYnw5+hHeEMfB2uvn
ChtCQf661lIsmy3fSv8SfH2ozJLzdU4yWqB27WEo8aMC61/OZOytmYSSxFVze1I3
RDW6NFfqaDA76xCpIoZMSx+ionhLAlbLypBONcIzllg8PimYb5iIBOpi2F6lh5KH
8GDIWTvOKn5pszH+T2JzsLO4YkLBkzekFyWEQXVm/GZT9xSrgCBA+yvAH7zvH5t8
4jpSutz/DOL4bfLiPH983Ia7CIgzX7/GpElwvXLxXVVqz3CaZlaMk06t9yfmCj4j
JArLCkQmDa9DJvXrPPca+V+c2YDn1/gV1GSN7LN8pFqUHb5eNllzwCKxZ7nF4G7C
fS+D6Up7iTru0GmWB7Vlm/YSv3TMEN9jdeC3oPUIC3yRe/hEaaY6h2S14EzEr5f1
2ZMruujBek6+pX2+ErXpYGxU9ewvU7bVP0WsXRIGB13RI0dS6yfOs8iZ4GMdszEM
vFMY3eVaN6lWPZ/x6XpPDVzMqdZ4cJKpPQ7N0iCehacoTbJS/xdM0oNamI6d7n6v
H/97yPa/ee2JY0Be3Qg1tYsHbhS2xINpMWbfjG8XalO+GvsVl6tu/uwbydBzD4jy
KcVomOFimRYJvJ8Vy75+vUdnmihxOhXxBDEJAxAIPvoHgweZo273GFrLD0T6acVE
A+URSNHlq+ToXCImlRWVxOJWFru19R7PG7rxPgOXFiG75/w9qtVzpeLHy2KNZRBk
/fSfdItCQThtWsybFOJ1ze0dwdsgk/9dHlO3jYAXCn1jS2U3JTB1HGnt2k4hcBke
pjw1WTblZplG+Qigtf+MtcLXxLaDUq7utVs+zeWBRN4G+MEgiT5oScoYNvwnsnAP
m7t2tYGOimu+NSp7uYWHWt0LsUr4CREGFsG0NgZgcT/ZVfM3pOgJgk6a8VeAKXqU
uVPVp08xGjQxKjTNj7rga3jlJhZxNfOEhtGRC0zTIBMHtEIvqrHjLV2265R7e2DT
jO1xVaPVEXuOK70LYJlCLLkRc/gtp+uVovKexrocGO+RkrD9ArJsx6l/QYsxKArx
9720CoNgh66SHAk/dQS/vm5oAoyyYEM5dtHiorrdmDba8NrW0cl3gnaGiHLRe4BL
bje6qo4KvmTGpQJKlKtN+cqOfDKLsyMGJIfr77eNIWGVlwC/6pxpVM2MQnSTDv6y
rOzYW+27Kgj8zG/xanoLtUyjaQ75yR8I1r9w3DHf87vNGrzYByjlyAxP1+dwHoiv
whFxrUTynkHGWhcAM8waziZMCMyLweCps1R+ahRCq72xfjBa+Q/1M5KknvA1Xzhv
HjFr1p3bk/G58JBfHVz+KJQ2HVtI3wsdpsZ6lnH847o0VIN7MUTIcuMKYGMuuiXE
80XxFruhwhCSKOs0RY0nwHKOYVWjCYChORGH98n8CIXSCXi1tCKpG5W3H7qvLY6h
fCkBZ+GkbBv+MDDT8Jl0qydd0mbtCZzh/ShNbHJ/EocEv+ahQbC877476oRHmQg8
KlFrnSs26skCdbmNE/aQ06Dim36KfOauKqdmvkY1B7ry2bKGM89IOFHtyA8RqL8h
l4Tt8iGWRRUPH9npGSb4Cr99xOamSnLzADDQY+rFJnwct+m1vB9yrXg/+yfYfUwI
gcT+DmYDmjW5ADWNPgCgt9p78WuiR7kPzPrzMvvJqBsn4a4CuUbJQ1TlEJLADMa1
MR4EKEvTya/eRNMV+FTjUSxKj0SpM6S5ZOa2QnAYrT9A/R+SNh1WF+f0cbKwXM6g
1ynWg7x7ifYMsL+q28QZAk8mV9aaSTK42Nxv22oSfhAd6tgFgjHjnvqBhmmR0/1v
E5tTc6dgHb6UTl338G/HC1hZpW0SwwL+SNwkKR1lXr0BDbprM6HR8CiPEdM7VMmk
5N71W1xZ+ke1HPEWKRLXl/VUwyf+sPtMxLGHDQekkBcsrrL7CiuL6gf1nJj2PZT7
YPb8SRPOx9qI42fi+LaCQVAoZvHOzGXf0ZSG3FYmfKoSgAwQ51+TdakegoFEvFKu
XgxUwH1dLXZYqCHE4O+4bMG9fP/J9Yfo4h0JDgfVlI/Ma3aKo0NRlSFoPvWk7850
MLplKfEzcl2vPLp3VH+EU1acF/1BTXtLDaacsNmUYDqN7CVDI/wYoW2v23SsSjHw
DHVSkdVfWh1TE4DX27kCBZ1v2vt8OktLJVmQHw5UyRPU08TVkICOvZeJcZtU+fbT
DFY03GlMi3lTl9ULAHPsI7k0LSYI6cA6rw8NtnLyti51z1NjyJpQvv+liQbMj3TJ
AgqxXycS0hGTiGJ3kkdwUCnlXhHy5rNDRn97z8uOOkyaMTuSD2VlLZ+w4gCNLFSn
S9VxwumwolnVtzaCyTVDnTKmfYK+820I1C/Zqhdped4T9z2fL0shDk9z190m90xh
E/4jkiwGVEu2FVWA7W9sCwPWLBWE8qDVJ+mVQhLlcLp3L9/GWgyzuipPARmuFt2j
Q2E8bsKaOcCRwtH8ZsV/sz/9PWyeUqMnIrxXZFfvPBpOCmN335pydwZJXIDeKOz+
Sl8PX4J5FCsGoile2SSOfe7Ow1XCGhWKeR6YqvTOmysUdYRYyeXVxjHRqke1ORCn
SVkW/yI27ox979ErSpZFDXxrmkaIXqgbvlAkuHUpIzci4F2uv1GJlACE9YyK0v/E
ALebUwU3M4t2D2gDs8SkdmI7XeYxUSYpwqIdI8VaKI1KFNo9o+hEGspHofZVsiqZ
1FCLetuqbxzEsBlzxecNoAiiGdnJKeBCjRpNgjbw5PjrbK8GrxOblVEOKl9KgiJB
o5/pdRIe6cnWSSFT8+ad9dF6mzpQmRAeJexI9Zm7tQVYmyS5Kiv73GjdZCFLR604
1mou8CG/7P5j3i2SBByi7P3o2466RxAlPhY+Aa1ROMCaLkzv+D157cmcVrBkDgVv
tlH+/+1oQt67FiBEDLzsCueYxh3fFXzk7CN/954USASD+zNvqunOhGh3MJAdHd93
YIIVpsGRrYKAbW+dtkEFVyPrb3SOjyfwP30ZmZGjSa6Uy7Pgr/J1jpPbCeruk8xZ
QqTwl8lT52ww4t5F7NHhKJ+rewGceBm1JsXQdDmoxLIG8FFygeHmrD50r3AVXb6z
2QuYwvHPduqYU2gKGQe9Zf4STNYgsKvVU4M0q94CRdzxCfsEzqhxvqiDsnhMZ1b0
PMwL1FwaJEHdU/iAZ2tQbkmuD/Vhq1jhhQwqfs1thUXBElNiBViemz9YaJmBrUAw
LcaVH/KmjRPZvVZs36TdzF1umY3R6ZxcVNjCxRXxVFkqczB03Ird4RyKz0b1ZgUH
h0HIYsQIuX4ysxcAGH/WYpADRjtuvFeyYELhjs7q/YuHj1t8LWk+sy3NVQNzKkNH
4hLoDyki+rkicZ04KzyaJNWeFMcQBVWiUMiRa4J6td+mEvpCSDXBqIHQ+XHeagi5
3LAawUcxzbQa32mMgekj/ymJfb2K15PavGs3M0Vrc1FEtW2PB1FpBjFLx1MgIz61
8utCsk4GOWOpWvXMm2nl26WKT6H0PCDkT+8pTSumiPPuruXsxzjqmsuxSwKXMM6G
0WqxNS1yZT1DhgM0HaLYycbZ22+gCa4/pvc6UMcjKkFE/LRiiN8m+BLGO4SndSCY
I8J19ARH/7JVMKiO/FtveZW/H96Cus7ZjJRcKFeb2v6Q8Pws+/DG1dF7swvyfBSI
ZRN0dmIB7lKr3BDXcq9ewnNhw/UE9KXeyoxx1lwo61s6Rg57YgPRBklnA++q+UUr
3RaEctAkZVe6vmzjuH6RuV34bqZwedxF8u385da2p9Yxu95QZawNYC8dmA/0HVg1
LRMGqEUq19TnB7dVdwGIDUEFE9nf0ePg1dUe4ezF7FC5znHCpEKATvOlKvIvwA6L
QMdXjpi3BQxpINyeJ9QAp6TAtRneMn6ndszPeCGDHMEBdychdmRujHY/ykV0KbnM
K/+EiZbFHxqPVjlLyWBJHcpDWccU17rvk+s+2Va4riC8NhB3Ng7ncdNv9pnj74aD
4/VYSpPQ61Q6Yzekv+Rdv6lyuJqoBQ0vOAb3JEge3nmbkpmM6Alnm8ojpjWkGIZL
yNkbYv6DaGNEUC/0mSIQOqdZoJhPaUtA0cOiP/97Mj+dGBeZ8C0er7s0XNtZbnvh
EMQYK7GrxY1A7qxB72EwDQKeXNQRe8aPmMxqBD2F2Z0uCo2YMi71epqt2lpn8l2F
bM7dR/XVXFA+kcNzQLdw4exPgoveNkg0pNnXCEBDhWi0mkho9KguhWGUGLUPLWhc
/fpEJC+fpYM5AYFukit2zZjan/9k1Ib1vcdlSQ4Tq1XEuQbJ1NkxlbgYuYhdbcTz
QnvGI43WphdRYSd2WBMVzsGxNRDoe90ZXT0Wd99p2R2vci10R3diFG7Ut4bkbdL0
xu1C/6jCzzfKT9YwmBPsNPMp8w+I6vYwKRAxVBbRQmG5my5WaJr+WYeKvqN3q9vX
WxYUpqdpe6wcuuPvOFbm0nBfkMQyLtUyj5rxjxhQ1D+0xQTIQ3atTpsQE88kTWNC
IJ/uXu5bxlZNjxpNH2NqdhJgcSWLJ+Axf1fi4eKkW+QUh026KOxf3eUGVHMbT9pP
bW5hY1pub/oqGib10g/UjCyj+uVp5iqhTD6u4v+ZSkqmKI6lNlWe9IAJ9Nbkhgkk
6vBEUyCEsShPTPdFCkMG5bQBl1mDQ5q8lfW7Of6PYSICAKnv71NqslhuA92hbXcf
dMByDU7fL71dXWm8VFdxuesi+1M9fXPdYIREEg5/u595dnMB+D7fSXx2fN5Sz9Gr
W2Az7mihy/YFYe9taIKjkyKc1DBXpHjL+fHv+l06GnM1QpwXhFHoCLXESIqK8790
WRbCeVC3NupEabpuvF+GV661RmqpgZ7nHhaABz397OdPmXOXbCcFAVidCu/jzF+H
Udcr2GjQzzKKHH/IxGO2xV2QBE+5+Z8QPlp6FjCCVsuXWTbJ2ujbLRZuOSFDhyTE
t7rkQauMZtae1uA4hOeychiPWajyQ9pJzMBwzWonpqe66bp5wfrSNYZVqKZr/5Tq
U+pTQW3CoHI8PqnpnphyxQVDvlImbwbK5eosGdrIYv7QYdbSbYXWmuFri4FUd8hh
Suxs/P/ISFYDkIhrapTOsVllCe+WNsLrhAPTz6ELAM4lP+A2s0sJYZpM6IVqqSq0
2c5RFNAeauzqsZu+HBel28qwHF9hVVH6LNbeCRGAo5orHsNF8urYSVmpHLLJvxYs
tEpung9U8zCxCtcz4A/MQ4SGcmVICSfg+MPqyyCzZMhPt2AsnABLuSIsAzIFSMNC
bt3cKtWUPydwWmLO7od2hShikOp6SQ+QEyTK6hokZO6m0aC6lEJxJWluBKB2D6KX
ajdA+Zkl5ziyVpyyQ9bptIiLAodh+J+xQmOsGzY7sXj21oaN5/Jv25+q7uUot6pk
MbmOPD0r2fHMqYUSYXE0rYr1hMOzURQpBQyFvJOFCQWoznhv3JAk6wOvuTdeGY63
jpYlsXdtFZpV3p2pEHIi3Ot4NAeSIdq2oaKvhUmJSq9FYvN3RLYGv2WXSZPzQv+W
+Kwi1PrEaP+bq+8WHv1ie743goFQXrMiKIurwpletIMz8obkGRw1dAwGR2uuxljQ
F9HV4U7gpqmj1c/NdjvUVZJm1IJASFc6HgqeqWw//ODe0SowXlMBDpjXuGPBqIuM
LPN7qapBJmeYdIl8Mbi8+pZ/XMV+rC8+zSv3Bsd/Kaz4C2FG55c/ZjEC25iVe5KJ
eHyC3JKkH6UaWsMcVVR8VNVjoQUiJWjWUhGUB7G8HkVFXAROw4przi9lQ7nFyJM3
g9AGsuV/ZwZzhBGUlw+3BsRGdKJm9318l2xZONIh3aNvHx2xn10N3GGCJsiI14mg
tld+AvSGBPmeB6RCZlrY5pamry6zReNg/fe6Qiyvod3Fk5tOllEV//B5zLaFCd1A
ikJ5BUyM/1isMmof/TFi0Zo3yYruTyMAArWxuLihC1GfW0KluiqHmIO+jTxvyMIR
VipTC7E9tiR7MRgO0YG00nluu6shQtcT/pvA5L9e2YgMmtYWVopkOcP0zqJAPEQk
o3zf89rDOmUTsKhGh3Jx7XiACu82oifkrLX8u9S3minT8I44dOq2iR1ERDLzsayr
sDsiFllo4FkIemcsTrSCnOlC5VGpQ4MsiZqLVFjXCjwtkt52ysCOphrR3ontH4W9
ZE5Z57XM2eYWNSuSo307UAXcbCVVRgzSoZo/VLH9SuJNsgYDxWdmTR+xk3g22ga4
Sf6cuDUXXZcto7ZeFK0yGLVnekoWKVc8ly34gJBRbKndfWenHm/vwOlfPVDeL7k8
MyQu5QU/i17IE3XTkcuUK0Gv0OMBEf4vnO/BiWGkcQrMgRZOLoBUpLBFNZy6dKZH
cuQYEuO67kGwNUmXt77TUC+fD7VR0jyFjq6Nw3UFJdcfmP+3htFKGxhtikkvXj7a
t5LEp40f5go1rbU1JJTsO/eHRRBvAHajp+wC0fs9A7tUQu5bPdmSnI4q98m5VRsV
wzAIwvAu3xO6EIxFGsjKcsUNGf51Nr0nglz3idNJeIvH7WZaf0BFmtj37GGEX7tf
ExyryNKQ44oMlroZtOf5TYWugJOrp/WjLiAiKoJixZTIbdiIN6trBw9lzh6MsDWb
9o9yc95SHjQZL1WNjRKIn/GqullPws+H9NcUiJUO2A3OlV+IHVpfFqn09T+U9Kty
XNWRN9bFVX9UiXs5egtudkLJK52/i3FZLvz1BKCWYA41W+xGzq8iHF4qGds19yoX
vWQR+YsUbTr4qWkVqHVRg40UUZzDhbTOq/s4FLOo+fVUm31R2to26gclcHNaneOJ
vaj6HcHznyKyXepOAcKanD7U3GHZrTzzdNaaw4M/ceMtb198T5KhfOUxCJTpkSTs
MG3/B8qc9XneeRDYAoHbAwR4MBjTt4E+lR6uGGG/OG/fidoCl9dJQYsf22jb1Mvk
gTNp8w5d8eJaWxx6Oerjw2xVo22EzG5AJ2g1IeYSd/J6BmKXowzrE+6AaWID0OdW
UemKyOPdStKdZxnUAO5tivVfbGjAivpLtBzJX7rohhHy/6YUCsZ6PD7OWQOZtkz7
u6GlreeF4RJQkou/Oq90LgAqWRM2vbPtBKHrRQr0gt4jaWdXYo7GaZNvsZ809BUd
Q8s8w9kt2i73sgG4PtxFDWRzxX0vZW8fDvDWKxVjhBwCWlGkI6P3AMcOgT0rgGOn
gsmi2yWAlcdPkBziOZrZGcnIX39aLAPcKcv+zdYclL7JGKKslUOG11PcS2ili9qL
aCkcvT6dm+hvnc+gx6nKDxUbVxOvdx5P1MBSV3J/3Ys0KybU6tf+Iui9x3Q/cayh
4w72K/zkaUHgM5qfph5+S3P0Ujd0+J710wdF014TxQohnMgEd2fitS95Jr//HNzf
3hMVC6LT/TmLRXB9LJpkmegWyPdB+TYE45WMrAEdM9pDaxiLWfXquZY43yzi0sMp
Peqha71u3gMJKuoro30AE95ojaDeWVjpNKCdnonntrsmgxCdoh00WAGZ/Skxz+70
9lXf8cuADFJXhZkpB8r3ZKsgo8iFOzwLuWx3u0iRr99VP2yIRRtGRJX7hS7aTPJx
DaaJoxBgi6GEufjcb64x+zaRL8PgIlcBPxt7j9ZZptdaCnLZmIkRPNxUUpK1ALHc
ip8hm5Prp5azPnopkHnWW5r9Kpx04xXX25Pd9nSCH1QOK/7aTxCIYaUK34knLoEU
KOyaB+E5R56qnLqy3vgY8yWhC7cOwMW9zn9pfM0mJ0v3qSLbxRSp/FY0LtobSqvB
mEF/efihbjU6ENi86OkMeItXlHsaBPmuCWAY8nKW2IEzVYO00v6l+O9b/5/FJ0x7
o8KUZ3YHqQZKMLO9BdrNaHFzHPR7SWTqc7ktVZUYZwuNEDtA9b17O2fRuYtKiMv3
YpeCdW5QkIIeg+2sZGAg2zK5GkaN+rjnVSVjemLP5/1ZNqEHASfi9UP5IMKQhLOU
B/vsK5BEi5Afvv7iwvjcqjm6k61bbXZt2gdRxhe6p9ggZalj8ya8kUrd32UdmC4d
foCs0L6KqWq7zXHUQvR6WHvE/bcYCnvMPOgM9z1P8kXcKlAhJrNKVnzLAfIYKon1
O3/wmvle8L34cypKb8AVbGO/nKL8E4fZdPeakIM446U/YA3r+msa07x4ZL/i2chE
vjeXHRRxNOP1/W4Rlea2eo6Of8qzu4vQiVmofkGa5iWGYFSLd7esxBdiFZQqRCbN
O2XQpXDsycmid9uO31WSVJfSFRs/BAAOsq/K9mXIN1uK6JwCev50E1RZsO4T5O4Q
Or0gg7HmhEXo0o33M6YGS5gfETivSMZ7oxlJoNiw8Ze9TGzNVZjvV+KqJXBOoHmf
Y9u6FYNZAcMQMpiAuph7QZDJqivrMNgs2aBYCgnI2FkgwvB8+8rfZlJ/XQqTnw/Q
8rnNlBZyr6Xl0fEVOa9tcYkaIS6z0dRbO6RDBtwTE/5xX2mbFTgEmlLsrq+fWKMr
9BTf3DgcCgn6XHNEQecwlXMr4Qed8+myHNar2dqrPr7JKg6oWSfneT1e+iTDtmKJ
P7b18peEA83l3RkG67678GWiSBkDBDkqi7Fv2X0j80SHbd3Rqo033OaMgqR8wUB6
s7fyLjsCG6Na+qF+nObhC7zNdr4pK4mjEV6w4nIKCWhUyATasd04DBLptdgYJ2Bn
5pQ1QGJ2kIMTOIi/+enSA6Pn/eUsTvLHoEGxMss1u7bNc7CT27TVFUuyKC8wYApq
KuBt9FFOivTIwqoielgixn9Irfj/JASwTdX7nRI2XnXAsyaY4gEGEM9exmkESXkK
al7GNZQUMFp0kY7Du1jiwXWnFZyo5hAF1LBhPtwD5T+sPO9XdwN/n5sIZbYnM9W2
PAEB7lOAkIji6k9cKmIhsmuQcuPOoKxZSqizCl9SrxMZlo0FdMKWMZkNR8jBtrHW
M2C1lpwPWQFlo5lSGeyneIK5bG4My58V94fAvjK9whXAqXSfNXvjv4GEtB0z3dTp
x4+Z2/XETdwVIocq7seQdmOhI/aFlRYpfWqo9zBAzkSvoM11d6zdoWyQcjcXgZBk
rBUBDMJfIM3kIUMYK4yKfj2IzZHo4cTqYC3QnpHw3mSeYvl1QAUmLiNcHD31TC99
+QdtAKHcRRoqP29po3nkQvm/QomH1GO667EQpyv/y6os+KZdNQcWIfCvdPJLTlZp
bAuwxeUq/ZE0RCIeiHRlroM0tSH//CCiPeKD9Yoz3lT9psLPUj2geRpM3d5yWCYQ
09mi13YIGiJ9A2MoWadwXmyKD10T8aDZCbwFIpIs0WlEgqXQ8q+82Jc4s0J55lh8
FvOvJzQcC9xpxkzIXos/uRxUNQm4Yk1RluO4QTb0fU/EnyAXa6pKAFwiI1uSY+C4
raWcpgKBpMIjVhKa4RsYdiHP6gRerQq/qAfLajapD200MPQGZrL98jU6e6jrZT08
66Etcip/TwiVlHTjLawMt4/mmO1zfhyEnDWc7iT45f6J+M7DEeSAyJEs78kqCfrK
aeO2o458Qu7W7/3aM5KYD3pAQpZNDUfIOpNc4oxqwmoXdQWzwOcMz+NKNmb3H1dq
d7dEuvB8IL4oRBR+7y70JuoUOg1QsFgEerSkEg39v6NvTRkNk2QPdGcc0bOuGX+o
hcziUS4h0NMCIkogth6LGEAswTX1CiFcUnLCWwh9wQV+65eOH4zltQ/zzjbXyZyV
masEyoEhAiZFlKcxsl6LjZ9Go21UfNoKzcbnx8/VcCVJy9SPXnKC0kKAzeNbJHwJ
1M42TSZOTYVEcwSyy4i5XgDOXewKU5SnhM1ri0oerd11VhNdVkHoHohah1K4eaja
Z7ixXy+jO85gBUd37Izr2I1dIcY8AEnb1/0Camz3KeM/EkZCRKCk3LAFohL23N3S
p3Agdz1qMOYeM1NWNPUJnlqo0ic13djAMBQHEk8xWVYyTu8vgQ9oS04fSgcdz4rk
1pzfTVf9bK79aq3LWzFUcJShV/gmm4YsJ9f7emXGe/iD35Z4x8zvvTB/VbEtUmWZ
aCBOnGqmNTIJCrIJ+DrL/OcOY+hDIhtSTRzydofZKU/JclT80zUugeWzjsaTu6uU
b667U+1Jl7A44hssy7gMrbkDdPQ1gsyASPYx9h0tN6FygcNF/bZEB7sHq+jXxFKl
jelcftvJ+tDg6PgAKCRWSVveiyYEOASBn65ppQjOz4nxcxujuBL2NhIcOfkJc+i1
H4cRqVq26D9UZK0/xvlCzVxWlwHLVE/1hWlglD59xtY+gVeC6PLs13uo60WiAoki
eQBHL6V8yIldLMdLlcoO6TlZKPmn+yrOQtwhXDyii0o56ljtknjinm117COXKz0w
s+QpFjcXgXP/syNqfWgdM5Cr3IvS+83g132cG4amk9WOEwd2s/Yvw5/h8i/6ZBNV
kmcaFwSUqQlrcgC3ebScfPz6zfPTnNi1Dn9g8KAPBsFre43irR54XAKWULneHI3S
HB49yNn2RCyBG1EU81qTuZeUDZUKTyWdxy54V4Eulcqkvb+XfvwDC/ElwybRHFB9
HVLzTFP3SVbvrXBVsR20RYpCoog1AN76kPx5PC4wruPsvRWVbk3iyoyij54Fqgco
OODc+zCpchzC7u2k3W10QyprGJu5+aZqbQvA9zPBGrcJAc66F45D8HTW36wwLwFx
rZW2CryFhRPLgF58451Q6vBzJgkj2LwJxhMutfvm/WV2vqbOuJJuODR2LnCcHH83
Dhj4BnlT6Gwqe9dySLynBQLLcxOGhsnDvv7M+CZNhZANob9c2tch7hDBzWYjBraI
VuwVfXa/2Bl7i0zkWXs7/Gxecdqwp7IOLNOKJL0SRdpSmu5Q5OmsA3XDped3ncOI
V4ez7sBtbTU4J+mH9/bX+WJOSRQySeLBBGGZLkfLiPZfbB1s/ZfqjMSA+69psQw/
nTVGwrRaleoGkRXIMOzUZbS3NL+d98wnimbaG1UQj/Sv8W+Fw6IVshwgYlJwxg3s
ftMR0ih1qIv8dZV7MfMMUcRlle4EaTHqJkkGYXNMDAPBUCsgyoHchzWjZrtriKik
72KTvn7SdUFVUfYjOX7ZNBTFYn2/TIZF4fuUrXV06Yl8Yc//5UdOybd3lbg2dsBk
3xoM7MnI4o9VCHfj3WEpq/xwhD3+tlrGZrXu326Jtzy0qKQksrmQSYpxERZmtM1Y
rHpEoEDKbAFCm8mGvvP+UDjlJTHhB/R52iuPlmjlKxfAhfPjcEAPeQ/pxVn57Gk7
68Xhreo3I+GZpNfcWqBGXBmRn9k6UT+vhkCO32msXubML8qIQRZ53uGvdLmsf61Z
0vMrT2ChcEmqEvjza6/d+5gdn13jCEFZIfEpsz4tJ1BjEyQ4Ek/xhhsU9we98zfn
yw1RcatzVcc3lfGVmbuRyqffTSpSKmraIRf7b2SW2Yjf6y1AuqffUWhFY7MfthID
ou09hNWqq3ZCoyu+ssUxZNb0yGHrAS1lVbVm6Zw1fdIAhJ2EfYptCxQoB5zZ8BBr
QU1xVGyozHdCWFI//VwikowbJkW9G8R++PS0S9oM2Y4ZP/cFEp1Tzqxt0ic+J+Ko
6/NAuaaMZ8OHhTBNsF9ZihLARtrWpv43ZKSJJRPXnfJc+dV2nfXdY18t5nMty8fr
ou7aP3zZ6qL5l0z0ijInOXqxBoR42/zgcVi5bx0lrVS5pWwBqngEUQ0YpvZamZrm
APtNN/PKM2KzrcSF0XqA6nkmww+YYUod+rU8r6hEqHgRxnPgujzSF2H1SzPlyZLu
q1IT5w6iwKlQ34jYoKA0gbmmKQetXfM1LuuO4xUelec2VWhtv252MMk8c6NrbBh3
aUF3fFzxIiCmKMoySTtZ7vWKfG/jta7Ph1Qn1tWeMvkfdzxB1hyWgQhIeAeE1lVS
YEs81rrcrLbODWgfDgGq6tYLRPFjmf92GymTzGM+qaaDsm2ca0FAKjthO2yEz8Wc
a+MFxUpifGDg2oRc/NEBwd6DuyZFFe687vPwlQkaOjQHMmBmiyTf0uOwcOS9PUyr
f9A6VFJ71h6fhPAeuNdV33HqrVLl6WuuPb0XvnO2pykQDNvJJ8bFMsrtgXstrVbR
jY9EQCL3UuVdrue0EQMEYLznnBc4Df1YE2t3LzOCWlIc82LLyyZ5j3CiZfApCLe2
qVQBtBZvBLokpdZOc4JiaGWhaVrvmh3+BOTVk5iRLEMpIyHNO80hh3eLxc1CX+Y8
DMsTH6J+4alwCoAbFPXzlAr8sAOl2Jja/yxjeOVimjI4/QB7vUGxwqW4sPHBcLG6
iBdxv6qfD/QQLOFRYhTWfd1txGoHxVMHZTjCq6ncExjR6myhqS+z1m/bBb0ERI6o
SWeRiZT4W/x1cplQI5TAZ5kuYlD2joB9bTIC7DJWt32rnXBxRxAjnhcNStt2iIix
bh64Mn6N+5Vj8WUtIcXIJWcJAlvuosXZqsgGUUovDhuCveftSSRzF+MVlL9hmV9o
qW+4cFJtR0ZAlPeTbr/cvjdCuOyyqdK8z4FXPYHbQodEOg6CNBjeFZ8Js8Olm5/q
86fbyxbITRF4g/jjmjfj9Opro8c7+nj+T7qGxVv8UcGIoHCJ001uk+5XsmxlUklt
/TiRUzsXqauK0A+eZFou7KqmZaFOQ2yuOew+V03YoJcr6Hn8iBWEEFK5mbIfYKLx
qHu8sLf1FajQE9Vv5C8H/WuoAqYrySuAd7zRgpoZbWeUZvXC/0672RFUJg13oBxK
nrmqNaXv9ms3XsW0KbgzjWRFtnKKIfFpFS+hUVjYMGRU7pR053YBoKe3jPH18phx
g+QewT2+CiJ21B8EVhxwGZas41wBUdT+BnokaflG3LoxNal1TcMAiY5ruYRMZDT3
9IJ41x5dgO/J2yp0EybHKOG76nYE1UeEHPoXdYS86fXiSfT/4Ym6dAqjT6mJgwH5
gFH7XNdrVdwnARhkIz/cOURZt6jgMHkV83N8p8yA0MVBmVYoSs9GHKZ6cX097SdG
IKkY7v8DvE+sndxGNyn6Rv9bsG7Y5qZYgFoTyUxYTyAT8/oMszr8o0Gri68/ro2Z
novKQTMyZsIrxuswxiznvNAIIv9d5LDPn2jJwZt0Y/33lZXBt8/t6eXiAoiC2Cyk
5d63SK/M0TESjmPxONTS5RWuJgEckISqSVW+6aa45YZtEoLoIGkZ7LwjHhJX61Y7
9M2I3X/OOG9NAP+iUwF++ctR6k2uUyTY+x8R5rGPD8hZqpr4QTwjB/yK0GeF+QRR
DPqYBTDzNZ5JiTh4ap7ge+YYcLWlgP1/Lmxu8QGN3uIqIbN7wPla8TTUDg01uaiG
SEHF5Ad72uJFtFClWaeVLRp6QXauA8RsncuxwdoICE6A+BJefCaHVND8HN1eDjN9
EZ5mdlWpt3k5vU5Z7lmmSFUc7krEQcYxTQJ3Z7hHl+0ttouNgpU8bCwwgn0rKn20
nJRV/CKnBBqH7STCuzUc0IyUZDBR+wacQ8QuvY5QPfzT/4eWnAhVdYCwe7/v+gY6
r1gNzMRAqovE7e2Dc1JElsS49PB3sG9lOHDgX5F4E7QrjbbbLwq6ZnkTUb6KeTuF
eZNK9zul5wKH/nEq12vT8ekRCMnLXdvwiC1hc6jk573RxGEvJi//fPhr6HzWi6xG
uqxoWl+iOPrayjUibsjo//L9Mhjo4yxe8sTT6OtxpyhLWeIUL3cuDS0Nu2I3r+xA
6ccfFKDEf9Yndkib7U1wD+YYmY6EuhfMY/o44TDGjsHzWbHlNnmj/ERsL6NxKkep
YttYGo0aMZbc4F7pJCgAEUK4mx3DycyvBL8/J176wdXwQWHwF+uMt2Msi0ZG2zP+
ZXLxqp46JAJjMOIkdl3Q3EL+nlkrSVby1hNIp5DPaVUtMvV1yP2VnorE5a3fNdjI
9eBlhvj2UKhYP64NcXTJwNH8dJuG8kp6ULZ1cu+l3d1C3CEBPEB4oouk+4TGpY2l
KXjVaZzClYMkiTj1bLMCXU5tLX6ymhdO5kdW850JuN8G1Wtra2vJjwSDNK4muAzP
LTwsFfkBqkjUPOASBcQrMllRoyTvXG3AwfSzQ+vVoAJnBRp6xNX1RlA8tel3+9Kz
5os5DeeSfA3dxFgwfjiFP8gJfaXs2d0p0mXUOxrVB0VmP3ZCoJ3aWWocA99SEv5Y
83M/Zpr5iWkiT2P+8ecTUh+HQwfp0XpKGadYHihw+fxALOpZR+SHdfSfFrwjx0/Y
vFylmxGnKdWn4di80Dk3ebSFcdw1Q8VMRyv9GorcElYAuCaLxmjhdSjHkS1ldnkw
kqRySTLIHoYaJlbs7XHy43eUKU9zd7ux33w9HGLYgFX77RPOKNCD9a1Eh/h5r59x
wJDMdx0/Ht1li54px27XRwLW9Tn1A7FpYymME0j3jKbA4OPoaqqn5mLwEtjvd+4T
cHyg9mS4fgKhI8ANvidCNHmaCy1Kdvtj6OrxsDlpuVL2smqDLRzL5JFbN3+VijmO
ZsiSC2L5Z3rZRif2ZqL4Dp9mO3qtluH5YwSfBQphAwnAVY+/gMhF+h0jwb5EX46E
aovyEPaHg34MLPQSMRAQWtvzcSM00FNTMt/+tyUY8e0ZgmhPzYwJ6E5fiG+WfC9Z
0Md32Jd5aK7hxk82GokYEzf2QKOV0ym/RE9WIg8pnrViLOg6CJgP/x5sPN/yjoMX
L5tknzs8dD/4nHFoCbOwqxLAl0SvYo6BsUyjSzgYOhzPtT2r5IW3KncOX+0me9JE
vKh+zL/ZpTYONtIeT1pMhCcEfQA5VkL0kJph8JMKmWmrv38A/DRM1GUHgtCpso+e
URnJY/1mXPOKyAUrk/mRsAEQ1gMrDyW+wcJAw6JHPYpTz/ptJv6p5daYE8Lj3zJq
nZZoa9HLaD+R/5XgNlIA9pU5zcV+Xikj6Zg+TM5dqA9zE/yNj09flMW7BC/vTheA
dVt5u/ZxaTJA2bZxUj6nMJ+pkkAYzd6XcCB6TOfxbZ2nfEedugcYYtwmjimcyKaN
JnBymrN5gbnZG6Psh9I35qjo5YiIS2brdTHOpi41nma6UYqkG8IILz1hMaKFfpZQ
/K7fZDOpfGHopRBKqlyxc0YPtmnfEv9mIeGwQq17ej8pRIEMxuERZQDjYZmSNwPo
35QwgpR7TXw2dHfoMCJ1exXdOKv4kD43eRsspP9IMFBdNG6oLhrIBQoeTRt6x9Y9
ZdV7A5fRyFTkV4iHKJ0Dn+psCuoTbGnOIXhbI7IvWKK3TC9tMVpeqscD2dLEjaJH
xII+uaxGfoxYlcYqQUHhmWaw+7+n3RWyovrLkgTr/VH3PWQzN41GEsIFyG98fzFf
oPcQoTXDYjguyZJpOsxW/cKCcX5rLsZ/uWQKwjIBZE1yDojerrT2ON5tIe1dIo5x
QdTzjzpoB/8QuEM51IxltsuqIsMtOa0722YLmRMncHsfexRwkyiZKkW/jKZqp0w5
UwJ6ynWRawRGYPWb8UhWANGoV0AATvXWFHTxW/AVxDKmo16WqPqFQgy/w87kT7mc
H9bkiIYCmyY3z4dwOPGDTDDC0efltmbXoDfG1ku9m6JxqwQmFGUqhtcJrjDiYEp+
l03OOIEGlS5nJy+Mmwee6wSQi5XAA/OUdSOCdH3b4TZhYbbpYflkx5ojirxx/T/2
ArxOVB9oXSO4mCyrVxL1VmHfyodiMbstQaQZOALhgVfj7LajZcd1I8+kQ+eWld74
VnfYcNUqK4y6SlB0R5oAY0pKWyGcWG4J5ZNHpFnDi2DxsVbjRZeOrO94w6rZ8iwr
FCm3MbpQivRQ/7yYAjswHcmM2ZCIVYF4fXG07AFy9fNv2B/F7MQ7u49tLgilVMOr
ql4gKVToALhOXrNu5d/l1ufa6fJxp+stIThDd9a0OxkDKpkjouY7g5SG8tfXcs9E
WdYKySgxkqZ+9bGUSUL9nJDRapZfUb98XjU+6+TWMGozFNXKdqTUlRaPAN/oWgDi
67O7YWnQ5EGUsvb3n+43i1dd85Voko5VgCMNJcHh7X3ggHAxbBQz0PEUJz0A/6Ku
xsPOmXKtqKXSTS4/kqcS+7d1Dpb0tsaDN/RWrZ+mNsz8b/d0QTMVZ+iwipRIkzkA
GdmVDI9UBeehysGPbBX4UTU9RxV2jpTal4j5xRoIWkv4LOI4jXYEh/VlP2GgH1Q5
Pj0k5WHtrTrallF2Y/uGtpDsEudLQh915KFX314JCFz8IPH7r5FJjBtBqC8SLI10
KZ6dr+G3cBRXwVp12y1yuUq4loMGwC90/kDXh58zyMM0vg1mvYwA38aZ7XlGoAgC
K6xTERHqG3VPnKNMThPH7guaSjx8KRSerslppIp1rGZQoLNeQO+j1dCkzTvpiQMp
7h74UQLxOlCLMWzydc0cIQma/L2DNnJao1dhpAxKIVX1zYaxrS+fAC8QLWCHT85Y
bTKSnYS2qkpANNt9m3DzRPiKUFV/qX2ibjGNdGqzF1gb0Vz9VIg89CvVA5yFwQJU
WM/HzkPa2IarUPwvksH1ibfOOD83np2R1AfJEneSiHLJLZ2y2db9zHXajYg+/wOd
ElU5QXubhyCkmPkl9Bbwlpv6z9rrWevjVs/b7fUEKO7P0ZkbAvW7dNzjqqH375P3
Q/4JivwqEFCxIBNIJ/o6T42HF7TMOuIiRYmmqqmbqtA2w0r0c1okXBmgVBZCwnry
69+jaF87NbzRqLD+FjrAwxEuMihOiff+DVvazuvEkD7cQs/Hoi3Fk8Ra2JZTYEjm
eNn4PVOeSVKSLSW7KCI2mDUMyIlDL3emmyxSsz072lcE5P01A5mjuc9XbQGoGSV3
9py0WMDuLCBJDu23Q46iklDWlYC2SMfhF+WfkaxuseLRmWRlSE/aNGzD4oseF/cQ
+EdRJX9JUiqDqoE3eb//0/TTlgMLySPZpPT2SnSMCAwvCxvaKuyde9oCfBSwvKLv
aCASMQC0iV7rcxudDZ9h3SlVfpNfct6NP4HglK7ZwAiMY4lyiEK5hQnJ6ZN11SB0
TP+qCjLvYlAqyDcoqGPLmH9hVn8FHitnqo6BsjR3dM8cDCK5nQAHw0SzSlWyCyvg
XlQZ0AvGjVb+a1TUQ0pU+FM9CnYcSzKtCMGIomfd/CLb6XVOn2N94BromBjSiFVC
lDW4OeeCYt/qcV12H+9Z1Zr5SsWPV/UByHzGN/UiK9oHdODrtfmn4CvRjvCwfnP4
K0pYwD16r5l4TsAYHfyi5r9CK00Fp5QbLRW4YfdR2xTDMLs6i1cebKJJAszWpjK7
2m/qrABJORrmkfQN9L1egV/CylM20XsmMiUP/VpeB9fEMoroFZaosPtWHXRGf21L
Xl1h1fLAwNhkUzMAT3J9bgT3Dco2WGrcjRmH1b2rmgiLRj+/L4L/3tQAWEWBd7RV
R1eAL82iunUd9FIpweDqR3uunuJFmc9F0swwYpTHOHooAKVzeBdVOKy3YedW9Lii
AK73bhiFcEc+grjoipkJftqe8Ihjb1FSewVHQCoIIoh0xR6dNcDiFjjn7rCUC6UD
0ijsn0PvRC09Tk8Bju7mk1TMqBwUoQKAPrIkbZV6/dMBC9yG7Sqm4CKN1twpkpiV
EsmY0sAdIOwvSsj/GxfNnADpdclFU2S/qfyOueOS0GCVniXIluD4+pUPDNeD7huY
QVxcObbGLFQV80/jr1PYu2AB1VfwhK6tPZwsapnjesiVCOznjEdgYJ3LH46YLf1A
9T+I/TJWaiHU+yrRXVubEyLxiVmGRT3WMWQDdYZjPC5eQO7gvlpOhFgy34+Qtm2t
8qNzFhU1qeYByeY8b18+uUPzpTzHArUdexMbnAVJSjc+ixjOOVVFjeA1VaNir9T9
ENzJYY0JK6i65NCkyYzEZwCuWVKDE5kTTMtBS/cIW4E3DdQAHuFRauZ8LjKwuCsh
X33mhAIzmiSCLBknK9IYYb1TtN9nYfKaTKawCS4lQAH601S0QTh25Zd1IbO/gxJv
1c9MLb0O/QRF+9wSGE6hUz3o36WHBFiKpFN29HrQije6ImwLLPxGUErEsLO8cqoo
DHhZSbFaSnos/rdTcoCycywcMykURVDHNezuLe3YqAKmPg6ns2X/T0cJYnmcISiP
vBX5y0Iyv601ztZE/BPJZxHbz1+3YO64F+QcuaphtvJBqW/7Sq1JpYfNM2DVjDa1
yfznq2FeVbCBcz6Sts+0kjZEXh5qQUC8YqMj5duHzh3VBljypQGyayoWdgnIEKYJ
01iwUnNtMc8lCZ/vCvnzjenNo7HJoJQsVqiAab6bQisUcfE9kX9BV/eCUbkmULHu
VEy2d5zpt9oR+81yAEAZWJwroFJXTEElnuT4xC9byjy6FMCyb5RfsXVGDwnQVPvS
EhB9aWire/JP16X2wSONrOKXYuk4TPYlDDdGCjeXOciT94LPSAxeAIgKcws9oNer
SV4nkEI+Y04o6hqVI/MTNO3/pbbuH91g8bt0st0Q2tmuDFgDAUrPXiKgDJ1qCNnF
GB16uIsSO0htDMRbuTdXcXggULKnZliTYi3jT7lycSSxNVr5gPF/3/t9hsqMfc4r
RT3h53pSfKAqoH5ZvXjLSwMEpOlf5UisO2z9e7YMOCOyGTL+dDXdvb5s/b3/tXzG
tEDiacurTz9GWm/TOQ/onKOHOiP+U1hsDOcX04tWF5keOQyWHG4L1oaAhevj0LRl
6tqmMhd3z1e60cczKsHgk4SI2lwSbQeGubeUE/VcGgJqK4dVjOUUO337xC6b28vK
VuzfGbEVqAX2IL51K4/SUyF8zJ9rS9BjgDzATDATXS8JrVpSbY1Cmu5cH5SX1G0U
0+cD/5MEcTpvaQwn8GVRgmdnEBeKs7RxX5Z30ACJxCvO+sJ9pUYXTp3umWixnQN9
H5fBgZ2Z+lx1VhRy6OZPSAzQaPMhMuh7WUEUyOJ4bjHGfKokcetg52+pDFrbR10n
wYSxqgqH3Hg1XEqATO/+QTgukyTBLaL6fYbc0yKv0pyP5+DVLs1tv7dp9kMcNTRq
Igf9axs0n5heO6IUpgu1A3VQmDF7gpcL8e3dlZX9Psf+Ta+57ae9PqYY5keocNus
h4ri07MIhTkPOU/LLMbiMMMqFQbHhImk5kfbpLosF3Hg1gBxatliYEhLKtAnl6wn
1SdSIIi/fj9dDWi5usk+qgDDSyKosjNP6mmcDI6LcEeUvxRqXJ6hhlU4jK1CsDOr
90GB1hD9Z90u7B3dqrHpHtQkC+y6kxOEDO1YXYhcjegU6H1rUs1E3nx7Ls7i2+RN
aTCE8mWvNJF5DE6oXDhR1JFuwr9EA9vMVTkSvkJVAEF5Xx0wKkEel4wzu/4ra2ln
eHV45UC0bsG2d19ZwQ0vkjOklzW8iJM1XCif/8ITswjpHcolLnxK0cG6HFr6+Ris
3xqzzOej1IdGC+lRlsoUyVxJs6AThixiLcxO2T/WzA3MEUEXHYVLXUQ4HfZWRpcq
0N0AUtgkkiQ2ru0pwSi+iZ4m5OB4hm0L3vH8ym/kvwH8vnnCR5jvz0S4aSu0fHDZ
aZvYMYSFeWDhoi5L0cx0C+0Gj3sX3xk0AoucnG/3dXrWvybrnvJC9/BedVYyOnAG
GVfAd9EhgEVP3IpGJJrLUgHgbovLh3crmzo4+qLEVXVfBnAfeJWCuXI2qRCIzhWW
ynrLbZAHOJda1adV6vIcF8+gm2jr7qS3sxnlx70Y+qwfA+JlYx3PXSlBtKbbZSbm
01ldcBPaN1XyI7+qNCZhDUCyGKvH/Q4KVfNBgk3Fujw+T30WT+7g2SOmuU0V9TPl
2OQgBty4JfINRiGEsbUQZjVgISnmjMOEwur8fzftBAwx+q5Z6EqGHs1TNPahVuT6
KFHnF/RxTGImJoRfPGAhkmMe25x0y1cbu7cobzCWjCFzfAeMwC2DcsqCpmYp9+ry
SmBbHRldN9yrkkm0dgdwZ1mEG0olNiblHbseR99doG4wOccW1Yz+U49TZvKHpSix
ZyaYIVSz59BJRjEfYuTgMRoDptKQAht2DojASBbMScW/UIG0GWieAxFRt4VZRV10
Cadzkm0tiu8sqQJH9WpOsYHsEMEsB3+vTjDF7BWZq9brTRdYBHLhSakJgU8UjYWu
lfv2xqZk5cKWTN1c5CU09C5AaqK6zEXFaE47tD6Mp1Z+oF8skMlhvRMbYYhngw84
kcMhZJtiC8Cj791IGya++HGDdYEWT6sj+gBV7VK77fHYpXSmcauAnlCOnqwZph7y
CX4aTvxrMRhGuZ+xuXWxQwvNOzRBsp94ciK9z5AtRJI0PVrtkSaux8Wv49sQ29DU
ZfgSP825CaJB56xrGBpGOHWOg+6zwrVCvuyJsYlRf/LKlAmTWf7HIwCyhQgGnekP
q1i4UZ1lmpE/3z744a06K3wM1jK7kKGodPrq2vK0rwMCmJmAkr1Pm+1XCzl5BGff
mKslazQYzUS1YlServKkKWiRIb3xWQSRZ3cO3YpvAWV1za77ajFR81ezbZD93Fyk
RzSkNv39JIaYytxCBIRzgy1jnyASpiH9I/XyL2KtRRlDGbi1B9gTJ/ylCO7Dp3/B
sSSzJc4UZPB50qnAzlRADI4iowDm8an8VWJCMnEEwKrEavbPd+NwoD563t0UdMQL
x1jAXjuD+Mnq4Zpu/l0x4ZS57MtlKeNp1TgJ1rEJVV2DuGGjvwkhw3iLDJMEZYjf
HrEN/vTR4SeAoXJfflXY66/4r5N094CMPLXsXjQ25zbg5q4Pxsx3hVTPb/ZSn7w/
BsPchF1m7zLXPkVOEuIMR90hGzdYZhgo6dq31BCdS71hpkjoJMB1dgmlCTbzf3ob
yiiTMdECaTdZQ7MIug79EoLkaTyaKu91bCtYbWGAFJAijQlQqrbgVAj4YseJOoCt
dHIqEqFZjwcS5PiRsktbxojSaL+ek0Nq3i11r4Bz0cGaFHyabNhxjCTcd4GGFNfq
B+bQxWF/V/2BBC4Y1rDMaa4NqBNLeWzO0YVha+YUCMaviT2+ra4zO3lyT6bEvz/M
OI/NfuMWABgB09haifCWDaz4wFbZlfVXLp/5M+dDnkAxxcU+LtLRHihnFQNM7Tsq
E8d7tLV2Q2Rl/IyEflD5xJX3eMBpElqArEPxx3Qj5DCSq5gzninws6bonpuOG898
7YVK13to2Bl90iRQSBSxBqgSHKAL97Um1VmVjz/X9stb9rrGfizEeNBfVQgqONTf
U/B3Cgmv8xd0eA3RLCh5Y4d2/lK1f3MDbgWhIuOchZA3Bn+4GHheWvlbch4n6I8G
kUgu5WnEsZTAR2ufvM7XC8Z1Sa0T5S9tpTpP1PgK7NxneNlTbHMpljtrxChZR+dy
joASL8SE20p0hn49PGSWrJXGcX30kE06M71nKo43RKJmZQzFmxSlP5IiVSqzyULO
d35dN7vv0TTXpsUTv/JwiW1pPCKlRdeLvOsjl26rRusmQWsUMv/+dKOQL3CqzoC4
ioWPlLKc3GGlnCuV7YfHitQx6kGlaQyRMMP1TAv6hb8d0hZboDcgIP3tfT8GEOSe
tPKK7cjjMfOUzPwwz0H7EGnwCvxa51nG1IHdBe6MtqxHt0eeqeeYvo16Ts+8trwv
jP8Tj4yIsffS+/6p+mqzOTklvpyL2utGcN0bk23hAVuc99WAy4S2SNzSzDrqmlat
5KfwFetY0+KII360iwhyt3sUdpcsccI0Yefn89y6Jq3njxIUfJpYg1fQJYzAeJFv
kd0sKG+6C74XzVgzcFWlXPfrNI5JgCC592qsYT6Y2EkaVHzLcI8pnqzUNfB6YkRE
3M2GBr7g+m/brGM0zvGCj2d2TzdEm5TZ/6rtswsMf1UVCVawaDAGPMFHEjqk+1yb
BKjnz7t/WZrpzvW//zG5dn742uIOwQQQaaiGCwa9NLyn+NjNm2bDsrVwCfNU4HTU
n/3yO8IneEWtw5W9weLwVYVSIXgUC/6xMjYqVRjSpEjKu4mjhmSJfrQf6w+4DTQh
rEJfHU2AIOV/HvCXkNFv8bsfGglbaCq6gzrGiG3vS69bNUUqtLWqlcgWlAi4+UQk
baI09oMzNSjGpYxjqDabavSrdnr03J00nZO97K/eNCUonA6nSBpNlPlETINRiqpk
gKnEpbjOP2IqBzbQAzyTMeXJTpnPViLsgUBddW1Q6gF6e9PIRc8OPBkN5WdMvdHV
WBCLbC+QajGiWBftBODaZUhA6jVxiGYOaQ6ryczHYXqz1ewRSYX2Y1cYoYN2kuzI
Gzy2VrfQRFL9PGvReT89Grx1gdhQPcxxMrtGIC84LUVJ6VPqcPZH6V79N3Ih1F90
uTA+l+PdzM8kfo9wDniw6KQBZXW7FaGDGxE6oVgBYSKh8kcygH3QFOpoTEp389XL
JwFcFc6guZLfwuNPwR3FUM3Q6R6A/Fuv+zhapbCenSEiRllsys0GlC4uKJ+JJK8r
67BYUEuDpWt1Fp67Pr8pjjTiE+uFqU4lEgEHpxyY/FdgJOBjI1e3UTa/wo/MwBwi
S6S+fLNP5YCdLyRzqozTF/y3TF/7jdI4ueWOHefX1WP6FyOpJCTKAC9TA8AsCghk
3+RMEL30OMS3sMbrGXiL5nRMPHxfs643ouQXipb6/1np2XRu4qfF3sS9GUTlAWny
tlyORIawCGVdQs51xvEQ0NKioccAIODOONoBXHeRYaxpDX2t0OqSn8ifCVwF+171
apynsSbkp13MPyahCQVMVItt0nsf0lOVY+GM+9oh/NROb0bkPrZrFRwPeXHra0OM
X8n6aOG7hGW4aLGQIalCMu6SQOarDS02RQ+BcC5pioSjbU+6ScPHp16tniPfHsUG
7pyVOZWE67+IbSXiqChQv2or1rwtlmgxFLwb0bbtkO31WcMGiJFK6te4DZzJbTaM
myEFssPCv40oCCONeMPnhOfufUSGcIwe55+YLl+vmHM0pLdt92E+rkq5Rq78rgs4
Lfe8f20wloxF1KzfnD9h8CzqJRMLovzlkfK9ORcoJsirhbLVTH9v3fNpCRZ8An9e
JXygVTW3s/cdSf4p6p3tE1+Y3AX+tfVY1xNjKdBvXKR4BLXZF21q+TPv0RaqTaqa
CxpygHKrmTojoP+/sXLTcVpS/Hw07+Dlu6XrhgEb/HP1uCpXxZsV5l0mrps38Pmd
w5VxYZb9WBkTP7GBjJhI0IPKl6Db8uf7QZvHY6u6bsUACOosBjBgPl8TvmG59grH
V53J0rMMniKY96yYerUOlXruN7nHCFIYWuvCFgCJXlo+Vz5Y45UqwfsTxOsJPZMy
wx/oKNRWTZUHgb69rSQjG7vFQer12mgwYah7jeXkIEJK5Dw/izjVY7CfPJNtOvlC
bqPrrYtadNWEGMnnWkdhw8hc0XFc34c/+Dm8BpdEmZbUv7HwmmdfVAjO6M+iXY1F
R8/Tp7xKf3WoiLIXtuTdFqzQZ/DKEHlrOgKw8ldJIA7K63XZTzSP6mjox3lnL52L
QqeTDj3UftSMzkASFaPSMPR4aMIff+oL0/CjSZ3I49BYVN9hO2WCLEymFGEaZoa0
1T9/bzmPPxZgzSV16VUCUCsbTMnY1MIt0rWDnQiy4hSDBA8Vu+532zUSlPfXqhEH
hsE5ZdzxH0gdPJBYVkNCd9ayLS2NcdU+oD0V3EC1j6/D0kFHjKOavCdeEbVn+T5A
zxKdlkT3fEUobIJsQ8MdlE5X/u4TcjEB6c8VhvgEzNfHDiaeJk60uUrbvQzrHyQn
M3pYeXZAtQNJjOaixz9Vc28EOkcGrvLbE7McxkNnnuX3lg7Phfx5OdO/O9WoEZOt
1GIL/l7Ov3AG7Z+Y1AXC1n3Yf9aid477ugqVZSbBT9owcbnaw6pGkVYfzy/fJpF6
p2cWm6AXTzKaCR2awpiUwowxE1aEWdqWLypsNa9DSGqBZ+ES5FNCMAjiaDpO6YwV
YIYXeqNnjgl6nfg1Nd9G7kXUtcRMx7O4B6J9Rw4OPN/TSFmmfgy3yvW5b2JHA/W6
u4TcHOlASBoFLpsudEaO99nbF55oNLVclEHW0HOdH0TiDB2tkUVIQ70c4lc83FNn
W3k2YJj4ALvUSHGXuNhOqVAiPQArYwARu2rV3JbJJdLHyMuxVXd4M/5uQplEHzxO
VU+FCQkJM34O8zDMdHlO8ZlLwDFXFsWb0BDcxMxl309CsP/+qk9Wkn8rbOcm4MPE
TCIngcK17Ya75k04BBZqeVGXa/joARJtnQEZdRiWMPzcV5qRQthPq+FnQIQ7O/7Z
q4zvoHBqqBhCX2wo1rhreC3f13u6xqqgrlb8CpDZM8bnlQCYgfno6aCqtxvX7T9a
UPl9FOoqw5q8zNUfRXrY+9ljJl7FSuDxFH6Ei80YTnWO4Dv6e/y9bEByqroouPMt
yaebPlB1MdjU5xPjHBzEhFYgoj09KSu2O2AExuAKD6yQDdmpSC3ti5JjTFjhTQ+9
9pIR/G9SUMCx8/2a2aatKkKkL9OvgvY9Uskz5FW5K3p6gsWLTpsQGZI+9m9vYlDg
Y6UGFlZeeJHpYiwoROkUtFm3UOnb7OYwclubowakWMwbfdem63w6x8xhiohlri1q
YTiLIIlkbzDEpvEC0icE4YN2NYHJX6ziHwmKooRbnxVnqKzJevBePiT6BmhD9ff7
2VZ51fHBYOHVb2nD9bQrfCmqTAoJQ+50N5KsOZSBer3DIrhlyUShg3r6mKGQIzw7
1Db6yn3LZkbOZTp05C8Yk1VXarKTSnxNwDNKb+UVctLXTjQ74fhZoRWwmbvPn8MZ
v6GGxEAbH547g7DrAe6sNLKZ2PsDdN2HimorU/g7j9GTr98vlNybPczklqsfyFgX
nQcJIMi9gLQa/5a/ZLbBvpzZ9XoS5XTVvz19m6HpczShvTg5PrIyPbj9dLcdZUWl
wJgVS1EpmSGx7CpJCrX3mVv/BgzUWa7oL960eHxQI1u3vCceJjTuUFQXfA+/JPOG
OPuqPydXARipRH4IguvrbctEz1S0qnciVz218+TGIRD93Ohz5kVGsk8ownTH8pO6
iTUrb48P+pcdYwRStLHVFSHgHFGLJkRmfOyX2Hw+nYrkBbN9hjca2RYWQEmdYU2K
OmWSwMXaZZLIW7OMFpBVKnX7jrDbepNIxjflA+mw0U/JgL2O3kPYeV159Nr+jh59
5KknybwlMZ1AxE0P9x3K1KNP21YnJJrcPwStlOiDMa09KiMqaWER8KTvxhcVl4pg
dZ6Wrq6zED0GE+vp2oRibJZoJjQunaWswILrVJHs8xekeUOtKx9MDM3dG12ZgJEu
qnb3WsttxlIPr0iW1V9AYUZhjAIfTvEB9jMcxjH94CzGGChkkHIacf94kI4sI4gp
DHocg3LeQ9Znxul6CVHirnbd7Xpgy+M0hKAgp0cLfdD7ZqsgKahhmrfp5mVrUGCO
0cdPzQgRbUiW6L0PLK4+kKk95+NLSEmW9J0E7NjAQ0ogyZi8MltxJWBpoTP3n4mn
YJ4oHh2/Jd5UH6VSWaL2yIbjeX8KHxLGkKUaCcBFwVlt9zkVdgSGpTPZBtH2v+vu
SnwfVv1cgDTSiy01dH/1kg0I/BoOkhfffuTHdscsSgb2mDU8DzYZbAQtuaPkjOon
XMz808iMRVGg60MSWudfKaH+wff7H2s/2JBsgAR+D+HatmZkC1MYu5ok93csz4/C
EI8KwAUvxlBwU0eDIvKEYy1RUu42zJeE2nBlv7n5tiWxnwJX8fgveOA+XB+4uGFR
i1CmJcd8/TsNeAtRTIFBNAON/TIPsEtkkmMrj47i8rcGbcJDJ0eQ/J9qPy9+SUST
7V3ce2ocxBtpP/x7NRf3ZKj6CBSF3T1Pw4c0hXS43GkHP+HoCWH9u1Sf73gXcNoN
lAMzDwgQt360HnUj8qzwNJQd/JU3ufoO864l4Qd+/ENftA536vuGdYJukROGR3I8
Ur0bymAZ6uHIOLEvGI8PlKFOUy9l41c4hnF4nCBAA0IxLa9Zztf1F0WRJVt3OyZO
yedBXJFo/BnC7QenRtI5VIJ3A/z1qRsd2JUsPTdHlXdFSvWe1pVXH0514JfkNCvI
dpu/co0PP3QvDVrVEtRhkJqMz68oK7hzPH70MBYDK4kE3K7BwyiAapo5O9aDxPRb
/oX82MzAz+sM3GjZ1S/n//Va03f3CNwuk0cJX8meUcaj/KfWxjFhSMPvzaWVgbOd
eKlKMNQTlcDPoVf9AomYhjM3bAJ7OQtMB5l3XyzFisnc2Z5VYWNZeEHMWhEzp45k
6+ZVJUv98rxrfr0+icseYnQ6Kb2qaWhUdmxDcoMY0QDJaQXomN9vx62qj68JUBD8
cX9H0sH7oNuBuExdGK9X588JKfDKXqtsHxSgbtNJKT3ikgE6bRVNkMZhsvEtaPHD
G16QLJ9mTXfPC1c96lNAHgahm+MhLby/vvh0eyqSExKgQqpl6FGSFI2Yz9eZWq3O
T9QzVOEIDmLl4/upcDomljQMcxoqrBtkQHdAGcNPy+Tz9fw6FPifT7/u5QCgbDZR
4t6egYq3r2oloQzQQwG17hKqzF4e+S0407W1ujRI6VtZc90iZCW9n5BjEy+eUbzd
wbsgnFdfql2bXjSiR5sLEiKE1PrkxeO/zQHwrSb0tlPiS4MCHktaOcWq3oGGN/y6
yYOQ7x+g03khnOH7R6inwjz7AJgXXWuLJ+XDoZQKgsO2cbXC12fBuIqZGTghYJR2
6evjrnK4r9mLNsKxDVb854tWq7a3VUOcUIBW0m1zOUAVVky/wB9lV5IxFFSLtDYd
V6ggxJgYEYTkr2awhhaT3opdSeJ0+wufwm0EGbFRu78qKKujrI/2sZVSO96UKPzZ
w7c4OE0ppOPKoasnZWZDO63x5RCaKSR9uWJnnph6RWdiWWoZdAzxzW4dardJ9TrO
pDTHEIJPz2qjbdZoP60JlDQno76Wsyy01ozYu4aZz0DlBb9h/9EIZ3jDXNOQWGim
n2Y2QkpzANlDYDwiD2Wiz+cyS5Kp9j8kw6nUOXs0RssmZkY+Ywaz+FU5hYItIQZa
O7as+QLaqF/AGUgv0gQumzS3fAT7OX4jdC8O7dbQcWvoqDnE3j3nv4Weq08E2JvR
jK6jszZJjTcsKVGAXJNHp09oJf8PtfcolC9g7+0CwVPU2lNf2XU5tmR88s8kdGUy
c2B43B3jXTHk3zKjSkBmjE6Ut9SiIzPeSxAIwVvcxLp1Xgm0wP4nZQpYyLF5uhVY
SAp5YpEXNJsvOvRbQEbGtk3XFxn5819esagC3n/xw9TSavK4qUg7j57tRTeBH29n
AMfrLJAb22iAAcI68E7vdWpC8hU4nAn3SicYzYmWlaonWPhfU0bBK0mMYR90iJCM
UQviMTueHJtCMDiEsbAOlXvWksk80dybl+z7KQUFZZaKIGL1MpvcJG9wkpdDiEUJ
cH1D3n4YMeord1dZgpXNFs+s2vNJZnRtVWYkG2zGZvygF9j+D8CKX326xWKdDcth
Z5mKk1jqTLyMyd6xjCLy4h6On2axdobIb+ZKjxt55/5S6O9Y0QX+C2qJmVsrTmmi
nGlf1nd2e6gDSlju1sFgrIaSsb8y8te8bi24w5PS/XIXuopD4LAoQOUksRr72BLl
Gmx8mrRHMArIORT5FCoMFiOfKYZtzjc4rXmBNOFvi5OMCjjMg6Ej0a921dfZ8X3B
orWznBYQ+32zObWKcyMsJTgmMV2x3BI6vWcXZ1OI60JpjrubihXH83QQVk+KW5px
2Fej+m82qYNjlCq+AM6Flt6AnFS5UPFd3Z+AVK51KCxWtAx+f8nItsSrVuuFC8FY
G/hrDsjqZqHflvyDuuhoIG08Yo07vN7Qc2W9K3bDnXZkp3PjECSTpIahKrnuyDuh
QBrSVOqAp2iSryAfEM//px0ZesZGFhMOVZrAFCgosdjVFn1uUvHmORYyHYHLeurp
Fl3rrLOiCts2uz2Wr0yT+EeDh2nNQKr3SPONoIT3u1lj8hUJ0lQd0zU6V6XSoQye
tu1C5d4fMTZSTK9ByV+CyHh4swpTFG3o4DYJpSulnuzrLmjABr6fAmaQVr0FUqMS
OTCQsXvz5xyDvMVNQmho4gsyJbmnZAh5MrIs2smGe5K0PAOoyI+f7vKGbz1FLgKz
+rVvX3Gh8IOZEd12286xdMblY9yNEUWc+BRCFtVohlQgjEhf97Q+7aIEg/MUnPJQ
AluFTsh3PGMjcrJCmJyjX05jikZXObtmcKdMVJK9rmcCHJ3RSsaS0glhVV5aUcjp
5SdtI3xOCT7fc27SrAORL0AuBIYTEElmiVxMSVzFKEeFWiEu5iykr5U90emjHxIG
+ZBr9DDHv0LfXxiqdSAkrBsaz/5wkwJ0dYE0xiN+rwEp1TTARtlDKlU1qKy+ZZA3
U0pDLsm+umqGhV8duuPH7KGFSPpOXQCWhLtl0pR33ebYH4BvZ8JwaslG8PtdKBCA
g2Scsn3c88RyfP/RQmfTK1CScpNnWfsmzl0c5E++2IDFwVtcloELOrFsRwcfY2rL
yfbxDshg0Sz8M/CmZhgHnwnHtt2VQWEalY12fC49FtD4dVBYGbLHYJEi6gxSEZ2y
TQrF8C3dLp4tm1ClkWPhNmSWN2iPlryR83bA861ot8sNiQ9T09sqmS7lcVabMeVX
Kd34PZieWKkH0l/u69kZmqPWFPmbGEXYRGnIi7u026OlQZMYvz2c2RZGhU37GMol
RxwrdiMtaOf9zpWGH0R1b0xlarnFtPGa/e9tHu4XmznSrDq8tP9zMiNoIwokx17U
Da1J9lLcvRAx63I08wC53c309LdWIIpB79meFTWgUllZtSit/MX22/iI/h1NPXcj
wIOYvjhZYnF8Bgs3tVIxqzKbGuwTLNkRy5yuoJI/7M6Xk9Cc3zuZk2f38wqGdmsV
uDOBcRIPlwC9iG5ZPDzl28H/wr6BLX4om4hO97KbPB2zBgCUD1dNuUqyEWaxXyNm
uUMAfcs13p22pvRf5iB4iw/MDEjTmQ9ee12XsEy7CZXZnnDR+bswc+mgB8xzBCMg
WsjvMePy1Q0AA9RAY1iecUlMnR1+iLRPUIVoS+gLfVbOoeS3JPc1EC+gfE2nq7Lo
rKuHt61Ok8XLysjeMVdlgShe0qUunju+xHXktaM5Uiw43p8bGZrFrTjfo+7vq4sn
NLf1L7l7XRzI286tP5uvMUUxE/9E0LmGrhhT24Va3LDdU7DaAySd/UZ+rIK2Sr0O
pyPwocYo+lEAERR57yvu7zNHx9z9elX9ScYbs2zre15OdWfxriRwzfBxKeOQHKLX
q2O7pELEr+oOjzd6QZrbKW/6OwzPhiphj2ZmsJLRZnEUtp4sRgIWysZpUA3vofK/
aHUeroqE3jnT7JmYhsOfqscp3ZAtTL/yISAggtVd3AW3lc/SyfkbuHI1z3zD2Ykf
uIX5BxZuKmzZ3oojGpvwuzX3OB7aVXaRNnDh97bQ17q1+n2xmfx4z4n9OsIvQzqd
NTPXk8+n+5MrVr8uglugudR0fWuaEtygLjdZ6s5YsO++yADOQ7swYx0CtHN5FtV4
yLbfxGqI7rH1veu1UFlYCzDQGQRnPdvzfhYkY9x3ovT68IadvhCrIcgtj6T/RFAm
Cy6KIgHuUmH39CV0UwgvWOKsS0qCaXhU3YKBDzMDBvDWpmAOwnc3CmUq0qWkQ19T
KoBPNIxxG4tacU3a8KKm/weTTXd6r1aHQ2S8VPtgR2dAjfrjqV1NSCD55NQWG09M
buTyEcxrMMbY0hX53KhIFPsRpmjgsuIVFKPTLvQ8vCQjmG+BTbgy8Gs/a1Q2ESnw
UHN5C6cjEHYZeQhjmOYLRgTKzTKRx1By7QQxXrv9bCCV2nAZTqFaKutM/kF9zb4T
tA2BxU1fLpJkCIX/uoXlecn+MyQ47Bbyfs14zKUtiPfRTHQcq6zyeWfVvcScgMZQ
MWLkpSsZ/lletjcte4xy8CFi/WaoF0tBmPtcNdZQx0zHaF+xe3Rpsfxar0pcuArj
1UIJ7GBVAri5ZdLEOUoBVEotPBAcIJSpCn3d6n58Lip/i0Zq6tPSSyI77y7TXodo
vI8/tgaQhoaMKKrMQ+gpEaG297rTvsIdwVZCg8icqOJNu2W5rq6SBFsMaCVEBOlZ
FIKdVfBfKdxbLQ0/ebpYv65lhEBJbYikm8UvcTr4+bzZ1pjqVADncSRt3qoy8Mcq
H4Ta/No7OyNR1dmd5YBfgJN4jzi8Os3rW/nxeo5l9AZ419nYjQXfKkiNJymv3Epy
rPSMAeQNVLZgm8h5rVB/y8bsdLqUKIlv7QeYTLQj/D0wmA/hoguiqIPZpqbu1fIe
KNGAG/TRjCrGy6D7ZrAt064tPHXSexgixydiTea/t3c9XykNc5BI+1E2GKDmAeBX
VyFz7inWeY0cFP2IdOQXklnqqqXC++JgtsTGTLU8mX38oxI7gILxbcNXULS92sBi
hat21EjsoCI19WqEASe66NgDg904q274RafRQhysqRQaUmkuCb5+OMeUg4wPa7jm
/xt6CwTO8lXx3ohYEWMqv4TjsQvV94o0pmd86CpYYym/IbnCmbV5PRNOoIDV8b26
RvkFgsmUkvpNRelP/wmO7ZqXQCo31HFq9j+ukhArS4mJwiGa3iTmgostGER0kGks
1Erl6pXFj/CXXLWbeLYzYCH9s7oPD8nrlUkFoS2eXKvCwmEEU/2JiaG7bNwGwhEF
j9DZJktLoBL5VtT35daNiDgP7MMACX/3AvNM+al6eVOxmc7UR5AWm1p/3xg79qj+
Zl0zWeYt9oN4F0fHanG+fbqLTfr0dW/PFvRSZxoufD81AYfRkwzg5DZ2D/eKgSWu
J3FMy+GMh4gkbSQCgjcszfwpWjHfC0rJyI0TaDlyBc9VCt4aa33d9xTJPOQ+W/Li
w7R99SAWSebewCsMf/obtXsSkioU30lsSaxGggvNvk1u4iHIKgfiThetrmqa9NZa
Rf2ZWle5lwBwrG2yt8PkHZmow4++3i6ZYiTu2UvcZXuENTR7Wb/46snE6XUVM9ZK
yyt3RniCZAWGbZL2ykUUoQOIL8nXSrHB3qpE/7hvX1s2FCHKbJMeVzopiTXLPWxJ
ZTqAYzoFR5ftfGvtDa5aYeqL+PFxXFWjhc0Dw4mPtvnS5a3NVllEiROAYf/rPDvh
vF476yKv/m5xjCnM4mciN7EXsWO2yMt69JzCOn7opiGFXvQ9IVkahKJtzbSvUmKQ
KYOWmObsdBCitlL/mlgTmSMgC5dCvz1p4MXGP+12N420CweifEwymjQzI/9+2AVC
LlrlujrfL/F23gqBs5cUtdsPpgciRCfO+wtogBSGpFkmx8OTkerihUVfqJd3Jlai
i8A9K/QDGC3sg7lb+KVDVUv8b7qLFXIt9AfVKeJkFH7taAK9v+gZYgxvsOWEMz5E
9h2+17HxlpN4Cdft0DRTyBqGW5pVNCHfO3Y9atUq3xe7ZxZkoX1iarJ/lOGJUpBP
TY/ExgfU0F7uAIRaoC9bmie+1qcWnOzyRZZRS/5VBuuU4HaRiOXt6Kbyg7mB3Esp
CNZ58Sm5RuKFWIsR/A8u0w7T/qYE4unaRQaWtCiEg774zsKaswP21qUd+491PaNC
kkmtEJi/jIHj5ikw05JnPYUpZgSlnQtFjaX36QmO40Vh27TXUy1FvSyl7Pq8Q3YX
Jams1fLD2yRddwnf91k2c4Vc/AylRT6YU6JDSwKtmjo6COC+CQmRnW3OOa3xCpow
VnN37uNRuQ/zmzHYgzOnvB1320bjcE/0ygou8Ri4dBoUYfweSG9VWRrdtdapvmDn
UdzXo1TIQvEttqvwmCJyvEmOvlnQVYuJs1XsEv0/Z/hEnukFt7trv1YqtC7fuZuy
DtopJdLOrEwNesI1pofL3HQXUmbnuHglVv2jMh2oAv6pL6wdcfBcxh4Ch399s0lo
8ZXYy1pEG1BwqeG+P9x6it0SDUyp9HfY8DeXUpeHDoMarCYkMBYMQD1PxEh2XKDw
oV/pHu0Fr8/6HDDU03obtaBiJ7scHhpQ929Tp7UtDcMTQ/wy/KhuW6lm34a3+uQ1
5zwflAWMra4xX9BNqpesYXDWm4Cu5QuuPa3O1r9nS/+k46nx/38bdJQg+lmDSo/m
1fGrZlXyuiMojS3ACcRYzqx/9I1Mgjo+JRJK+P3dXYexL+IeJMMmcDXssK/OOs+e
KRf5I2teA/Ace7UPKHjwHpm2Q0SqHwQ1BGhkwoSAnDCiLCvE2Fxpxf6y05NEXwTc
0gWr2DZwskwbUPgyWjENEUz+lHy2noOG83Ptz198XyFDYKQykwdIoGiROELB0bbA
HZyZr1f6lyQ5SY+BVVMlCy30djwhyYSkNRa8oBBBJaO3OIgG2GUebdQiSVOliT60
WpTyU2BsIXUCfJD5D6G4GQ8Y5SNJTcJg+ypavTkcPwG228beKd77+2UlH5C8v/GN
FHgqNDKyCbIXLUtZJ8qkOHRCmfzZDR1OxPDKqPqy0jm4N2EDRkOiigq0g1cEZ8+g
C0eEXJ6mlYWT9StOT1/rARz7pWnjbH2EbzKhRy3yrYMOC/jGecJu3CGYVVhCrjA6
ZmvzTvdtbrH3Bj66Mll369dsmhTQGkC03bzUpH5oIkArhHQlDJP37l0xO0coOw5o
oHGzcAvlnB7hmsGTsHpv/ert6qvoaPG/OpdavHvJ4inP04N/OCG8nYflBJpLy1Yo
WsPnbs2Td6xGNIQiBL/+S07e9Uchs9ayrTwnV4F0vFvmmFP0CCw8JdL5pbyXV+fr
qdM9FdoRskWF4Wy7dyJ2UH4VKv+cPp49SNO8AZ6PDBq8S8E9euKDcYAVuF6BITFO
B5N9zzZEPmYir22Yu56Fa5b5apfjC+Lz5mJOd+rssvSrHMC37PoJhV6769a6u+fn
4m3kU1Lvv3ZIctv0Ea9j8+9BQQm8osLAwtD+JT6vtuZMf6dzatxF46dd7dTbE2SY
PIMR+HmRhOyzgsYvYx3ETLCV52e2GFHsRicOZKCRM/2XwFElx/liCKhw94nP0MaB
r3SnPhjmmjXOuHfxy3Bg6uuuOdRpPmV6DwWu+iVs2IW41gvdy2cLhBpkEnA5gsUd
lV7AMB+p7J83qtzZAR9+sPUlQyNOaBa1Kf3eUJ7/xzy1Anz3VpXjQEf2FTiB7MjU
0JsMEkdEuiJ2/Er67ly2pwiIZiintqztgs4UbYbMh0HIlSGoyd+WKMzxKETSUgsO
IauDai4XFGRedSxgm9OpvwkgAZNITA4IRVnzp/i+i274zFwQUjmvDWoaUM4fbI4m
MyyJyj8fFfuolw6c2x+tKIVdK29dqC0DgltKkUQh6fBhDNU7OBUhKkzCM7G69c2h
fRYNDmnEBquUpmOcXMAhNHw5Cz6+qb/NB5oSvyKRqfTP8SRrUO0Xdo3DENZaF3y5
VN+rTHJf7z21gewQ8dHHKUbNFHsV1R+4FHj3EUVRuxE/P9SJKXBeVmi3og+H/94v
AOAXs6LWS72M8gcTQj6HoajNZHiH+tPLU39h6/Vsoeat7Bz6NUgWjSgC6pDqFZKJ
KwF/8wjYUl9ynZ9Nv7+BuRdIO8Ys/fRgrhshR0IUEAri66+v7Jp96Adcab0CpcCu
q49bk72ZufRMbl75ImDD4CMIAbGcOoCHAPtp41ibZiRTmg4KFO21j529ZCWwdsJZ
JgBc2UZak2a8ZJTkJQkevgs1ChXBAnWIfFtB2kq1ID5k/WCnqxlnP5ZNtBIY4Vi/
mN5l7Ma0+3vmWcIYWd8Ydw2kiSVoTieoWAXLYz+aJom7EQV3qQW3hhyfudHoJpY6
G9RgSh0pNAyqlESjYwGka8IzySlgO8ma6K01va2VuT5Lm7FNFBh9hl53nIapqQLi
ohhSqrAS9C16qrGOniMF+/Lfn/S9P7xSk+MllZ1SxygsPiZrtA6pOGiFvCSWOIuS
K8sMmEPKzQsi7XXA+dLw/Gg9AP4fcTsAqs905xEzWFCOUGEyXYtfRaZ3RP7gzMM9
i4B1MIlmP+CZ3rDbq/kUTi1K+aSfANJVrUVpD1D/tXLw2upd4eJGjeWOc4e2531v
5AC5B9W00luSZGjp7eDInjxsX7Yz/LtUSA6NdEPXWq7M3ei6IKquGmxpzZRsHAsz
l/Z8qFvRHytjg8WxHV9o2+jh2y1f7anzUO29/rqtzOwWpY1IfIBtOV4+ZJdmFyyf
W3Q+zYEsGILAb2cAQdsW+D8PgPQSP80HWt12yAcyWszvoMk6SuZX4wVU59iZOmLh
kzvBjWDUz6w2earyYVqti5oCEJy75IGY5uquGGBBx6tY4W/eifKS21pC591CNpun
8+FpGBZNqfg7I90Ilncxx4xbOxBi34h70Drc4qF0S81tILT4hVnW5DTsN7X8vp+X
csCgF0gJ2ZG3PsZ+L/EBta9obmIpvPq0Uo87bMjb+ZQwmkYk23c+klmLacjaRoR9
xPidGQq9xmFps6JCDk2EbtXh9DvNXzFofPB2VpIhwmQuqvwGf8TPdB8P6y2pYZPU
B8i0NabrS0YKS8sWCuLt4zy582YDd+W16VwTnOQlSG37kBoea4TkFPl+SBMrR44f
qCc3kUDMBOC+N7wa0KSuAhe4s2ivzTs3ncpzgktooUCurLO5IqSk1FXdaOqsjEcy
xt/2juLwG1fOpeKo7ZLh0f9nL62TAd+Nh7/CdbPz2IZM4XW2LsqD6qpov3vFFSbx
rDBPUf3ffRqehYHeZKtMfPry1gBPDFYycR/7gysPMGhyOknID1FHmuBVVCtUk2yV
eqprIREHDG20cU2cQnpWQmaHYC6Lrduu8WuKn/YMX+DWkEAwem3LypLWMTvpbjt1
nx9ZQ4t1vPzGkxpTvW9qFQtxKzshXD7aM4IklMUgO1yEkAoB/O6xdHIl+RIjFcY0
ELq09ODlgmNsVKQsH0S579VHnJE1PYXuFc64JTURhsR5d8oMN+AZG99EptbegGdG
eyHT1RIq8y60VCfKLlH1Vo6KdwAsJGihMikSV44vSN7H3d3tFhIrjqGgIK7aNjEZ
IG132fXiSgfOGboafASLQy9AmHqwFuwdpXQG7CoXFY4ihINb1/VkORn8iXp0gkNj
RNJwbTE72VnrNHp5dzvCpzZ5WMQSz+KM/8BmdFERcoDuiliMwgqCVoB2vatWVd0D
PLgvpW1RgZdBw6ah6/JkdBB2GQhBF3LXWNKH8Af6okoTXomEw9aHleVj2qbou/jp
obDOeBv/eAMvCGaUqpbNxnl9jSj4xfzeqFugbUQDSXJN05ZBWJHn+jFP+A72XLWn
mt0pJLVPB1Y5FO0kY8Oew6KlQWHpboo5ehg1V5fwO7EascsPIIJfnqT1wrI+31dv
NTmu3zsEyhtm186Y1FSZ2uTMY5yRrMXYCv7nrP4Efo05CTSvvlTKemWNHPN3Pz/h
/yTA++iXf4JofpieiQLWGaUJjQrgmtphMxawsEVRw0n4QGXtDg/RBKaT+X1fIMlt
MSwRG7Df3UhqZjDX+oj+ue2+wdaxINm45svkB0mMjiycK1P6/q9AlwmNH8YqAzeB
j1V5LfeEwP15PLEKjCw69jFovhDKhxF7NI2Ax0ebPhKfjmsRqvPzFZN5mXQXB1FR
BU8Zh+FnXDNpgZpAeqSTYYiMCdIBuVVy+K79fKIa/yNXCrtEl0CHb6F77IQS/9tN
nGFHB+ZtU4AGhojhwHX40Ka2twuO+x5tJci9VrvMgJnpN+ZBk/xp025MSbVTLsjk
VoG+ZDgCU2V8wRG8bV6gy2uQjxqRuytIXcIWp15CNb2wLWDc5+ldw85l9RZyKKIZ
+EQ9DWMVocmVtMEJtuJD+srJu3vvi0HkK9aZ+FR8oD+sU4T7wS8Z1FHqHlY9eOCb
qlRWRCcqWYJXJEUNGi6zUzVQLn/EsGMOe42j2ZG46a08Th9116lGv5YD/J+gXfMK
rMFf5dx5NHaXtp87x5uBKw3jgdkkh7prdYHJCM9c7rfCBiicku85quZTI2tFSQZ3
wPFRek/K5rxvxUyBaEKIQORVXMVFrUS5i9K7F2lhmnl3XBvdlZ4DTUV5NzyjTYDK
vLluPGfFux+aX0Nw/ICYLaZh5zsJ4+Qd6VMStknfRm+CGnBpn+ueAhDrhh43aUv/
38jamtP8nMuAvn3kB7lW8kOe7DUsgtBBISmel4J9ReWJLebjRk4RWjWPxlMWhauq
uEa/DgFGBLpe++NFuClyWdVl/2nXKuYn1vsop66lLc2KqGEdEwWg1EgIvj46W6Qv
DuYqsHvUa/mXOTdEl1mDOBIlkxMdeTM7qo6LfDFE89N91MTTNlx5U8ynzVx43TqX
UFRh5Ub4Z9rxbe92ZF2wIBqNNBF7W4KpIOJOvca3AJW+SlOCDP3WKZILPOs0QiNp
uISkK+bo4NBAF2F1JxYl6UYRdkVQ8uvu6rtMT9nJy69mEdPmmF017wG5xitaIlt+
2HVzcFpR/WD3fhQKgsTsS0TMSPjB82KYD5tw/9H4a4UgbmFYid6snt6O9ngz28Xm
ehL76ytoX950a2kGc78Ky06XlYR5fFORJrAkZF/N64yimpz4H5WM7wqCMSxVa+gB
b7DAod91TGjFZ3iSZmTUNwp4naJXny3QupM29Vv/tnycMoaFlUNHYweYNOqgFL2f
vcv1BXYzkfLLIg5ZsLbkJLyY9lbkLYLvU+VycleWc2aFPTZbGdaAuEORsKVbuT1k
8hC8XpbOMS80ca/omVKZF0SlDG3DjS59WpGEoeiYSxt9mIhNqdldkbYL9RvqM5uP
VqZ+V5T5f5zqH3GzA7KUgOJZlTp3aFOpgcfFAMu4y8oEZk+S3JzaVp3ln83ojX3q
qdKKE2LGT47fgDMpJJrEHOAin26siGTS3Sgs9LjL+Ju3i7FaA02gXtiSUEqnYomA
iq18SqCkY+I9TE8kBzSgMMloF+C2E7/XJHKOZHaOHuUxPUG6w4HrNluJpzESdKne
hfFQ/jKPWM4knb2R1GjKMX5999tpaj6skTbBCaA/P8m8zd66arX5UHTLjvZyPkUp
Dq7/cz2vijv8d5jEp6s8HZMhjjx1ZMVI5D9lX00NrPt17gkapGub7Wdo0v/rQjlJ
i33k6zIPFc4qaLWrHX3H+pCdoW2FY7HIh2IWU6GsQadpkJj9/YQVkkhnYPQhT6PB
+jlYPwvlzhECCWsF9JHbsabJqNPysbVC3dXo71yIK6Kk/phNTy/Zdlp2yP4Io6V0
Gdp9qH7NGOzfH0ZUn2Rns2nDVuU+2pPDXoNo5uNZ7Z0H3l4YIyzD/+KbUm5+kBoM
4ikhUP/kH1knlpyZdmi8aJz+RTy9JR4LZIfDXOeHrhs1NlQMt6c050yTL1XUPx1F
3U9+lxRLUnWPI3jwnzDsJwp9Z1WAoecOkBl9z5C2Dp/DpcTtrk+mw4VRz4UFrnQ0
hsvOmYlWFkOW1lRUqdbvyjKm1kkwcO6O2WPH5bj04JI1CHLdfa63bJk/AAqqtMRK
83OjG509W0+/Kpu8COkenvTYNLuteLzy7Nn4GrKWWk92f2Md2Y9dhRa146qo7c3k
yRG8iMa0lOaRBJ5Zx5gmix/LlYcCnKvYl5+KGPe5BGK0JbeoJGsKf0ZTYAURXI9t
hCXO4L2K41xvUzaIgfrM/b5pm3kEjpkJknbquXR4kOHnplodG88Qd9Aj3jJgSqpl
kOLirYQF4ByJknPRb+zWcRKnS8VJ5nML1Ucm9ejK0BqAMdtZIkidEtoLlmqVepAF
ToKheuFxtcTooRL0fuYrOqzggH13B64Fs6EZR59W+PH/HOrGc9NAGqY6pKs65JY9
gS6AV456mtxptE9oGMevaRnfDUIlL6h6OEhWZzw2gFpKFCzQTvQ22lqNZW4eVCoB
VYsn0a4MWDgvogOC149zOdPDfsw/cD63zcFeuc7qio3ZHny7Dzm+fiUc/nLlpvjL
CrZxhbkn5PjWS9MKpC2IK3uUPDTE8l+dK/1pw2bkSQnsC/Efe6nTOPuLnMp1WxVi
L5f9POhi+zXyN6/OoTg7R+psUgAtib8rkUFLMXIc/PuMm4Hz4dpIGPfAPtBqvu1p
nZ+t7D8SpBROTa9qNNce6jVzAIWN87KIwNP++fPHymezh566+Jzhs17aIQ8IyCLc
TiHVpVIt2vkKTPoFrvMuHXoVehRgoVQ7LOXLJH7ln/x6z8sEPPebg+JkOqosINi7
4nyzbC2CJ9vhwtgQ90lPibt5U4FocMtkVU4eWLWwe2RCfHiX5yiwwBJodfE1WdYY
APC5or+5TBo9XRX5Nl250t9/7SVR3UUmPwtJzBjndaAwceWoTKnGbHj9x19hBIOn
62fj9n7XEhEnFa72+DYB71YAA2/gqes+EbCsu8S14SSnyN4MdLi+OFBIIotMUewc
gqFE5O3GyHrfMnBQtF4IAuARIMDtWG+SoMlvGWGvgscxOEZ5/N/MAOvkUmIQzwKo
oxdvHE6MBORlh9N+RLwpo6xnJYZS/u0+eNrLUQVw1WTZXJBVLQlvPecrCE6ulOX8
/kr6ALSBtI1xu7P/xbPIGMUjFIPCOwG1HyPYni7S5EkobMPxpEHTYj+3GfzT4DkT
3VviZ8l2Nro4VfDVZRw64QDU1kF16Li6MsmuRAXnWmM3ZzG7inqO27tP0hyCsQCb
urysczxyzbBE5wB+h+JTStrbWx1QmO+kZeh8D34znE6j54Iz8t5gWmLb5wpkIW7U
4UNkSMxB64jd7L4RXeb7El2PEWQs+3i2bPnR9qBQIYZkbcgx0uoy/YBD0Yyyk6K7
v7yL8J5cZ62rbz3OD017ELJ7Op+VwIqa+V8H8tqQRHC48TCSupHz1LaGdJLoZcTZ
hta2+ukxP+/xhTi4Cree5zUsEMd9ep52YSjJ3pGpOx/UWeBUc1FnLoXT0KmsTt/h
BHjf9NKBKDSIZx8TJn5ZI077BbDC0m9QN/tU1A70qiPWG2XySRVN/7ccbcc33xl+
MxkgezX545fg3U/ZWhT366I2oyLL3G/OGqdPd5RMLcsaMpNqz4QgsNzBYuovIqZA
sBrEdEFMCDCrUPuDGuOnolltDaxu/h38jbVk7U0H75D2a7uX/HQBnQKr7mcYZm3m
jypYWiwzxQE0WL5RVuSWMXjwmuqJXh7ZtAkfg5Ukuvt03GnNWU6TbpM2iSDQSL6u
Dsx1rT13pYX9pYZ5ELEk5nMjbkMO0jgJO7qIg3FlbljeY05dHPhwcR29Ohc4xYKk
3NZffEX1F/M2TpjVevJT52MqhsPCOv+kAXvpRmI6FxNh9GAMyH+ejBIsT3yNOw3e
IwrUPQAqwDnOyc0CII3pBxcCtDfgeLa5l/qHw8FDCfW8lZ5J4UI+nSvIJQQo0XQc
q0lQLn85UIggWq3MrD42WhDQCuezzF0/NtxGKkmEU7p8r3N5BW1P+NLlN87yGS5g
KBbkArZkjXemVAov3ZAg4zB3y4VZmeemkxdPSoT34iK/10nkZ0jCtyb8szL2caiJ
fNeJrHkipRoVU4NqOuYkkobWocMk3C0JSMAyrKDXhjDT/VMCBQbmbt2HhnkAvnD9
1D+Nn4vVAWFBwaNKfJysbhMtHAayqFa9D4FMzG49uPny4C9IKDG+88tBjW1ohzOd
lygXGYC0MMpwRb638vaPDtal8Ogx7mLXzo4UCP4ROskyO6TGZEydp3jTaGEe4Ynn
9XQscxs2hc7uHuCo74zRWP9Tneaha5RQxizw4QuGJyE5itraaVkALgXNolhE2CTr
e3kaFUzTvCnnFA+YYttwX4nBBjvmvxFGsJaxKi1o0JFhkZGmIj/XEObaX9iz4+eq
T4iasogPCkVvHfgRd9zej95U8iMFZ91zl99Ewx6rX80+pihy7zadkxlsQN+Zniw/
DOZxYq/G/Jvn2a1naPrYuocgeq9+TaNI8Jn9tBZEwnuu+FHikAwx+RVwoddycMS4
HZpejKr6L/wAW4ap3nELp3hkhlY7s2atzfg8VZd6kOxJM0lmU0rFxtVQByDEKPfY
zdNEDX4N4kmn8gk7oDmdolO0s8epMpvZXWfQi60OqoDDp4DA6hI64of9mXUMyBku
VlWsh9NKa+OB5aA/1kNUT68yEamE34cNRIcjcTcyA6Uom7l5Lv6EMZcDcHpIE07H
wK5w7yurPgUGY1Uq+jx3zsgZvhXXdulWdQ3WaSn9Vwbh2v/nNyRtO8QD02atkHDV
a88ivZbWn1Czaf9pPyLDmbSncnNs461LIxH/ZBLw6BvQuRGbDBfJkKJOkFP3iEP2
z0CKYos4nfoXant9VULvoj//YjEpYPRy5B9TQN74YXtj8M3gLga5R5uOdkmP5d/V
Jd9uzrmtj+NcyczD5raLI4beXzfZ6xW8cV3nhTPtHDxZMscLAcydz/SJBCdGlbYb
1KUJ97p5H6O0k1vdHO6V9wXnKrm6o2/5+8knRdq5VjiIYLCXf4yyyP+WudfKE0Iu
cNFgk+yKG57tUue2a++wRp38GwZ8sKqh8ckvA+fkSL0uk24oCPMs4GS8Ers2dgK/
UXPS8nfjK73hwp76qoMC4U5S/Ck99RmzGpAvHCNDJjz7TJLWZJ9ys0/K3QAocZRM
McOZ7SvtSWnVXYlQ9dKMMjdGJD93BY0aTN6B59qjwyKiTs9T0KvKjp2t0gC5ewTx
GEr1ftfZ1t/4yQTQm8WH2+p35r/qu1sdvhxRXBIJgF85/J008xdRCM69StujblPu
aUqayVW5LtEg4bDm5aQgoQYeOnwkicT3cIawhpRgzfgLatf7HxcvKyl7KrGikMZg
a6QyVYdc4Au/QSVg95oGJarEp7a7nRqExxkG82kR7Ei/rxmYOYe7dLpEZoI17Whl
TCFMRsni4H5snyDu+2e4c0TA0IynRYuDswegYUtNfM8OXPJcLy5WxFLSaLCylbvI
xMWCIYs8oJFOIVrg38UDH6nHp5k+jWvoVuwZn1NkgGvhiUV12KfMkqafyyHdXiFt
ZhKdHPN5DaRFMthXG5V8p/HSli7E68NUnbichailDKWuG9Q4zjwpYrZJ08KFC0ir
NuPQeOVd25FMDkpU2dGG0NhiASk9Bft33+zdwxoJduxqF5RXjX3Ef83C0XoiAkbI
2zyTJR9MRpC86B8ZfmxZgEzZInONiPKxPul2l375s6n0bpJ8x/mA0i+eHf6nUJva
AQB1KYS/jOo2wjyqIoFs9vP6bZeFPDMmJo7U0t8GxxYamuzmpUT2OjfmVWCWjFph
9UW27wW/7mc/MyBlrXdImiQvKbdnTyhmsf9TnqKdjdFrQvfIRyA84bqPiEuQdCuG
+Wm2BGutwaiMMzr7ELfDI/c222K92wqp0nkA4n0rzGyEXMEqESx8iceH3ve537S4
jLj2alMFpD9k4OrBj7qiA4NpdZ2in6B/Mr/v5CwthzR5H8jfipsj6KTsSv1WIX+8
0fuCxgD04rBFkKiCRilntcb9gMrejAEuCNEmtyOcNoesJfuEBycbpNugPww2QT3V
JJAojl/Qtb9j0sjoM/sKrEPdswP4sTt/my0qJhnrTyv7Kp07z3dO2L1OuTmYJQYJ
zrGIsb83YR7UGsQmiMX3JqySC/s6dsZyfrSuFD0Kzf7ErUzDoEp7EMQT6CGupx71
kEOJ6KITUEIQa/4I7Aw3t3QNX8z9Dq2xp0AaLLrD2tKmI/56q6TN07tqDLtNfSSB
rKj1d82xdszYHQV6nR107Y8lPzjTAoM4UFUUHpidqipZaVdPC3qb6xPe/g6yfFkr
i6hU17iUMQ5EONBmMBQls4fLpvzAsHpWIGIPaM6O72g9a65FE1OWDgc9ydBy4pTm
txOX12BEXvnQkw2cVkc/vmqtgu4dMDbPvJegGrUvH/Xvi08NpKwHt9lgLUfHDKQ6
qpnd+ZQWRb0BFfXG738aV422nmUNaVnY2Vn6xod61UpY5HbIiGRYdvApVjJQV6U/
FLobCyjxWyiGTPPZu9gNxC5UGkP2Ro1LdMoNdLnmMJkyb4rlJoJsgGZ7kotaf55B
XkDD+Ufg5JA8vRPDU4Rc6k1ndQ28fIRD/yCFguGcdD5BxDd67oWyJk66kr0tObVM
tkvzvs0X5xkp2L3dIp1+KE9rUrDMxKMYhpOmU+UivyDKPZpqnHc5v7UVOgaXddRb
LGliAYbKaluA9/YbT9laaojvefENR8e3/pA7CBfDCIoIEJldVVvja32qx4XkZrCK
QADdwNtA78idlX9MI6omT8dX3Jh95iOE1ksp9hQfuXnGuspSIbChCHx1OLDyXYQr
cO4WNMvh6fOAknYR8eHYfMCzx7W4cc8AYf1ztYKdmQPz0V0pVugWNOfsyJ6JELKT
PRlyPX7kDKVFoZ3RxRMMM4HTaASIqDaJuek6EFjjWZ0fS7mPtQxU446DriUGVXi+
c+Y5jNc2U5NBkvCwL4OESXh/yHKtzZm2ORSxY/nRU0/4VrhyiB+NKNd5kGcXB2Bv
7JRAchksRTtShi3Qvbq9SyR56W7OXMAUVTBzOVe4OPgw2WW127y+IG9H4n+92N7x
GLUyL7FUGWVeGRI/ROEuDiRSeXkyRlxyL3ng/VS7kugpF3Pf5gC6mJAKDlEX5o08
hwZtpW0ZQfcu2zvHr4Yb9GJOObzx6BySMWjTFRVttaSImL2ZA3RIFxXktbJVPdRb
yS0d8PoJSxZFsFXFWjEqnUfTNlvT7+c8EtEieI05DlvsfFaACSl2lF0AtjJQFla0
0ODP2m5aXVvg7sR4gqtqmn7AVdV1ezdhA0+G+YTx2YMXnviaJ3tOsNgh99KM38Kc
Rs18vk3V4tY7xbP1F6K32ejHVzSW+DPRPVA1Jy2HLSFHl2UmsicR4CnLQDwHh9wi
8H9SGC3PxWZoLl47FqXoZceWDbuCDhKPQKgXRtwZ9qaqQFYGJmid/lZ9aDlZqvjD
ExZRlYNrjUGbqxrfgZqq7aYRaqtjDXiMLQmxJiJQ/VTwHs08gPs2Rn5Ytyu3JeFY
t5PG6r0Izk799OLfcsi1Kj+UYCKhqp4kWdR0TZDoV51mqwqV3hBPZgVZafPwzQ6p
zCkqBy+BexK14IlkFNnqwcXk9gT7SZeLK8kOqyAW7jQyRbWWuuhWTsbljAEgRdjY
t/Vgv1s/3QG9TtdGxtiMHuwL7sci2KlcSofj2Iyly5JywOmk/L6klGpeexraKbfD
sGv1h975oc22RSH+IOpGnRAT0W07TJMuGDRTacb6merjjR+I3b3lrtUaUTCW8gc8
j2OJacQA3fv9brJray5DHTYpSJiq4Utaz1fYK4/lzYszm3X4MUzx0fD2sPpZPh5A
bkEIWUmcZZmkW0Yo4s+uEhktkBG6Xkvsj+8aMSbFfgq7UAudEvpyvYtlNuBTVGHr
RAQnOkN6m/ed23uPhm/fjICfSctGVbDobDFOFiqX1ideBn8BWuQoV9OlB3gN/m/u
G/6WzYqJTAhPaYL+Ef4RIVODNJ1hL/UHOuQaL9I1UNNyuptZodS6tF/lPjANgttZ
LOnHPjnrdVQk+nJqmfsRD3C0RWgt3ZESwch3uaWYwbaGBQ1eYiILpxj1oi9Uzb7C
+T/O2go7gRqtYd5ZAmVqxmCwWpK3S7sjOwJBqPOWWXVZxq11XBwHJ4mVjX09D3mW
J4MsYVyhUli/IlJ7TbxSkDnPdZCNK7SX/u5vU8Qr7woljThQolXYGeB6vKel+7wm
A1PWzQLUHpQGQh8rrwHfEPMI5Mi6oWVukQvUhe3jC8f2g/bXHllgvnpdFcBWYFbe
7bNx1sASAiG5b2mVRhFimFZcg4A3Nmm+KsEPJk588v3QaaHNrmBqKrs3VZjQemVc
qqNH898uMiXXRC2koFBCbfLyOM9cAlL4zXHrJkEYmSWq+GNwRwqhVBME7X3cZFhR
1EguPS8/fjANH+KNnvgJaEVmEiB3fiZm5Juotyrk7vEZC8N/YuQm4qizTkei7/UP
+LwG7d8bPeLOjUfLEfdOOJ31nJU/MD8wF9qRqnvecFVxsZPqxhUiC3/sBT0n/iHn
lVn7fjMt2sQbbpmn16fTP9iYSQYj1zj9BLF7RT7VvaK73iLxi/0zIg4+kti2Zy1j
rUNgAQgzAo+rLxkGjFr96wmIkgElicmhkdGGl3/knUvbYDYnKPm2ZBTJQyWl0bz5
RTaYkfuyuBq0VYwApW1FynCJzx47Cu+HRFopWWVgz2wVhspbNS+6zljngM3wM1UY
AXGWowrqh0xsUmKds9eL0WDiMT2w7czFJBuE2BE0ez8w2qHhM20Sbo/loxlcmIvY
hnw8xB3CCt2Onxz3zx79Z1KNsrXX+/gUl3E1GoyR2qiAD5LC3zaRydNjmCWtUmCO
mW6JbpSxAvOGiQadOvfV4j/WKAxI97b+Lo0EKoJX5UrpgaWxnZFKjAx20hpS3XnB
k3eKPsoa85Ne5Yr7SNtCDfL+UglsV/SmUCZ4qymEIVyD1LyItOy3mS2VvjooWiEY
j2Q5whn1qioQbWQtDbxOBpyXhy4UgBJvUSbs0kLgPQIhRNXvQTtbNcrcyfY8pPGY
QHkn0RboAa8h+tlhuHhlYlk2DEc8vB4VgqLTDnIkbp8nf9RH1+f8HJs3NDs9K/CB
eqPyfxpAdaL7BE2dUhUDyhudOrN353OZCDYJ7EAjFm9IixwTtFI2lqKREDZsB/Ac
nZJw5AjroWpgBPe2/rNZHOkCseGCs/f01envkiYEBuPnIKqxYa69vZ38Rdof/bG6
gz3N4nOiEsz8mL9a0oZHAnXCIVLY699Udym8vkf0zMrGahrD0YQp5lSFv3LfD9kk
vgmdD8/jscCyVXsWQP7FefvfXsl6hra/akSErd+7HGCDfRZi3ZxPsF3YTG108aVh
DuanqobyjpEVST1gq8YjsFlgrxpk4FRU2s1bgs9saAe9LPzlZptcHL7roMG2RY/9
ZzvkUcWep1x1Y1sT/3901foi8JMzW8nA0t4CToXUyz3eMr2UYzM59miV02ESasJW
RrBPvl4Asm7hWBDGCZenBAAjGgN4tjV+k5YMrTv3bBWGL7cqSdrDAmFcHO9HJEVy
ZLJxy0Z9uS6HqkCCG26Kr+xZdrCt9v83o+olNeUr2UYzX/fMfXziC3qvZbxwuHTN
k5zZ3Mtjz+j45fj/LOIrpAyKma0VRf4hk9hrz28KWuC5T3nuyRAWn4ZR8CPINpwz
VRVq34fgkjBpAFi1fqzOC2x8Io6J3UiHSpAaS09urqqb8Nce2H/4oG9/V4dNJJZG
6Cse69qKkPrLEWnYUFwKYAiKvUbnf9lEHLMjW+odgqQml++odZUcPl3nPHtR6WyO
n68lq67sKf9TABcLJ3C8OECEVs56B4+RJm4PRiK0cQbzdQvx39YDE5/CDQNJmjF8
bnkzS5ewiJbSIOVAO9BCv2cen+R4yu/ABEfxCEkXZpRojNrRKIhVZD2rRFJ3uI+N
+8x+G1BL/O+d/xnfC28x+NMENKV5VlN/T6xxiREdOjHAwASlVgACk3RRsHhe6S90
eYEEJHCnva6hmFMeYGd1hCDFNru5wp2RbRKpNlEc0ftUxiUbP++KsjrNNLw6I3Px
ZlEK3+S0yogsJohLTi0QsGm9JeC3vAmNky4BbrND+6rax5mzXMb5RM37QYwOgHXF
pnUrrSioAUOq/GzmM04HtdiRtZADSxBmgCJ+mvYuDr49q5b1N55F45LV2UnwINxu
9tdXv17tJFpEaOgu6bJYAiOoy66ik3nnyiNbDpL0qaHTRmxMkf1uQgLlIyhoUq+n
SWkXJWGv2NxC0ShJlthw8VYslVzGW3Nf6RcVE0K0plQjjn2ptLlfbClIw8kWVyPm
IPMIpoPwItNrqhfzo4i6WpCdS/6Hs0Uw3Ad3RmMAz2pMnb/vvF3hfKhD0VXm29hn
9k2BgximEK8Tu/n5kxB8iRZVT/ffZHxMIUWUaGwijPdXlemAhnH5Gf8DyID7NIac
nJ5d7JDNAMf2gFrZm1MI7AfX9ekPSGYHEBkKOs2gxNDnHDNvZYirogRLnh82uviy
2HI9O9ODabkI7Umeu6uIrtc2vIPZPT0RKKC82Z5yNgoowaYGXac4xMrsO9lCGYcR
APv5ZA2t7/EH4ZUSyUm6YICUhC8kN4XwAtl4LmPX2NuTD7eg3x4HZlwBmOMP+zcL
FWGhSXG8gI3Bx6Ld1gx2qoq5opxTQ7VxUdqi2Q8l7iDIABcJLLk8/yqWjP43XFXU
NSkufEbH2M+o9XVovRBUGn6J48mtg8iGR+6Ot2LrConSZb7THBqdKaGxNKjaoyVU
vxwrY4EhRXIIAyW7y5jq1PFI+sXij5JJfC5xdj1kQiZyv2AJ6kvpdjUp1VXIH3Iy
QVMlcmE7GPl6pjXFV0S1tEOtHSK+7LLYFe2au5f0QxwvWGCf4ovto2GMuml/uKe+
cbe1zgJO8F1mHiaatkcmsNntVelAGYrvGsxeXuBHgYqvmvL9V+ELcDrndqeF+Lne
vWkgVWR3ai7v9owXFxGYU2rzJsOSNIoRpAP98wubNJWEqYXPnVOqxFwBMPaUOSYh
bhGmxpyKhhmalvKC8yw1jukcBybPs++OzvnRi3pSlqKPfjHgbclqwlI43ltEcLaX
LWOPg0vcGYw8gZZ9cs5IeJx2+6iu2ASXs7gBmkVRn1x2s3kcFvERfQ/DbR1trHl8
qp/nmkQ05t5QJjYSdILsWmzyrA5bDFnryC8OX+6G8sqOx11LL3dcWIv6xS6B/jWf
h4rzuFpT/Re8nZwSaSlvx2zrzLuNb/kCUupzBzsdmbC3OSrxjTTa6d3Q3h7PmA26
OFAmPz/MTG1+ZkUmZdV1sIfK8aHOJe2ouPzWGelwaC0cHnFeizega4mMCdphMzBE
zNfCoS6OUml1gKh8i+WggIKIYi48nfZuy2QwwRJYdMriQp8V0uF+l1CmNS0cnMAo
od0n88dOq2gkKLzdaUwlz3jaVAmXAnLhFhByo96wAgNRcNcZ0iKCQWrtRlIYkCfy
WLd4I86++KQKK2uhQIQtDAkgP10CTIJqKQ7J2dTaI51ytH+TiORvLlUomblyy5rw
HS/9Lh08/qbRMdxZtiTQCjdYMU8aYrQqo4dBHJuAcoTr+K/WCig4Y8tKpWlzop+h
mnYnnbSkwVsHjd2pkvQlzv3Hl6W6AZnhWdmio4o6RwednOEi8FjIB/ErjmSo79QU
6wFLroFkmp5d0VKlb+oB6ysxQNQBCPK8VDJOyGr2ampe2hU4f82SCEaWWD/zUI2b
PY/eQ3ZYELf55sYHiaCMpNzkR8LWp1/GyVuAkpxLMbaxpk6YqNcR0R5go+A0O5rU
IjJAxiyxAYJuOgf97VurdoyjPGGj4W+RsdildKgk8lvnZldK0jRgCPHCIzDTLoOr
bG4Ty8OXtN34quwCKZFOEb1dDZR0TthHx/WKE3J8qomC8m/8lDnIs7bUaesBfK46
pGLzDuBv3lRFxIysH0XxwaiStXHJ0Y32qbreGFILFdshMBqubtWpTxKTzYh/dJ/i
TyRRynvteOBYRLVMHTmvJp/0AHsXQoBiNbkBwBNSyu049eek7qwly3rnqofIk6o3
Xt9T98ARyQBRDZRCbZFujX+2m+0BN1dN0ILvWKuHot4XuIa/YAmervjKlJjvlPqX
MEfNk8NK/l+p6daJV4yeTnNiTwDK7E8+P7v5RnpbaB/mHOaEWalwGBX1JKJ0N7FY
7pJ7W7X6Hw46S9IzivERpBNibP29F9Tow1GM2QJ8T8HoZy1eVIb6liI3+LQKjedx
DeTRAN2jqM/cYMJ4B8zLrArbwGCotP6ep9rqsXcn6HL9N6kmW1Jxlztd/lwGxQYi
4N0QNPV9MKmjSsNXOWpTZxwaXo7xWWCpqqx91W0Dw7jYyBql+UvxWXlnrbmkaaex
H9OCmWOx9ma9FVVTqeMoorEi13DXXe/OAo86QHgqe+ym/uXjEYSGpSOLQd5MyK6Q
EWbzrRIKOOOiSw4nws+6aWasxhk/nIh5qKH2odBDdYGupzSf+S7D6+INnUQYtWU1
8hSO1iSJws3G7sRfFfYf3JZh6CiBlmf7WEr1M0XIwKM/OwE4oBfzli1NXeEIUyee
0ZwQkOt0B7Ct/oh4AsT06IGeC81CYoxzetZOMFhd9SS8wiGyDNTWyQ3tbi6VWwj7
uw+BoOQRVb2gxskNMxOPsA62dpMOr2VC9l2Dcm32fSl33HhUDOxcko8jq27UuYTe
2XKO03KH3aaYkZDYhq64ElJ6vPDVTR+XZOYy93bspd+LMZezUsNhT/k7MKMT25p8
vPzmWKOOe5y7uywO28meeGHVsv42EBz81NYMOfN0ulGTzhlGMyPTCP693IAzRNgP
rc9aN+nI9iUcdoDglgEy95y4cPaEaC7jBa8zjOjvdStOhVMXYfTzmKI+eF23zJop
kc7DlPUwB0adJEyOSIfRKnNMAMk0FsY52Ufnf37biC3XuSixZUVIeR4poVfuH/WT
qm5Hlfyl49/8o49dDGQ8Ls4YXNfOtXff6NJvoVkaduHXEck96FPfSG4Kr/bHyVcy
nD7YVNb83uTXFD08U0qm88hBlgBFdgicF4b3bBIyj2b/zVQdZAQ8XZAfz690TtO8
C1XhX21Ixh5TZWESLtCuOSHQZHY4y7ngg2MDRG/zoaDw0hyuqBHLkkMd3l3DBlhi
l2stwrq4ElaQC8oFBO8LnrYwDmuh0xvHRq1umFqDBNQNJcuATIkWmha9iCn4u7l5
RbF4HD82mIXhxstE8tU5YfOpGNIDUj8EgK6qPL5atU9/+e1FiAz9/+AJIdSOHQiT
KoOkXKLudcyMwDgoLNHPGqv70Fb9L/N8yCvxni6A53osDUMJBxkVgbcOchcyfvPb
HXGrrdXzHAfTMVgu59TbQrmJHPvkz8tE2EbEWW0WVMV0wJ/hPGzIPr9H5nkJXwCL
EeVGNDU2aivAnfWYc6iBSSrG1cGOk2lTSSZItkaxI/ADpH9SCerj6ETLwBZ/FP9v
LOKHqvI7teE/+YEOs+fCOPEqCqy50ZGy264UzVM16CjLxZ6+pB6lvARamvXsmKzE
WX8WW4gjWDTdtZoGn4FANVODOBt8xPJbjPr+lEPiC6enf2tnfCi8mCwQtTr3OiX2
NXXL/kV18m2FvI8RgE5k7pxhJw+svXZICyyLNx3EBGW0Ml22v4omiElDDSsUNVxE
geA1G+extucSF3S6vSom/8JxnHgl7qHn/xm+VduOn2luyv81wokdBBoX9bXQPHDd
6lhQFwMrteLrJhBsH6ZX8h1jmg4RwPfWBixjDoVndnFjb1zYFeo7i3v/h1qg9Itx
sFvvtNA4prOh+oCQfj24UAMsqa81R2rcAnYuA3legI708nbDhIacTlTSuWGA3VtJ
BGTWOgKmS2WsVgyypYrErQF6lHSYyblazTuWdX9NxdfxAi9ru29KBKKLl4n13HYC
K692A+17rkz1YkqG33mx5Afq4dc04Wp6KD0o/FDwf8lJUfgCoNEAL8QK3xs8rptI
UBOsREHwo9Vf1lpONx8jnqc8bs8oZaafkDEJjyxEH8jceuydPL3SRlCv4E06c+QD
V4BqhhDkuZRf12VdT+C1mP5Al30SEZx3b/+amkaKBMDFsg8SRMgu80EwufKlcvr7
HcAzt9rs15kGZRHqo5nSytEY8+RwfMS6YzV9hJ7WT2+0xHkJZwF5Be7e779dGlH4
QCyHdqo++ALJYu54rDHRusGeO5P90/yaIkxdu34wT2TLL5+V9fY6raB6hs8mJhZx
6Fr1DOPahuxrUEGc1v7SYm3nBBd6upUf3CsiFOpsHMEfItwDO2JRfjaL6pqBqDVP
/H/bL1p3hoMHQpWQ2Cgh8Fhjk5HbqGzTmdH7AELu+CHIsARPXa+fOG18wrNWinIK
dPN41tt1AjqCPyHLyaYHbbkJ391dJxqYc+ZhElF2c5KRMjd4BdBJlA2p3xIAFMhu
/tUFNnx0U2oMEPhB/8kF72WpvnG8r+yD/UIQlLSB/8E9V9nQSKzzX/YY9rBS6TP+
nyvu7wQZTTAAZDh3WWtnuNx/ZHjzrOKHRLdsymaCuALCh9cSrC7mvKlwSbImzQ+s
l80l1x/kLRU37UPEQHDPBoFlGVp28sgMOEVNtyoZB82mo9CJZ20sFjNMCg5oHx4Z
H40c5tfSa2cnxR7zsbcd6k9/vQrXyTANesQfK5MbKx4Rd2YVhjysIedHaGVN9cOC
S+fJ/iupBcPEFD0mEkXDbrZFWGpgCt/OUD0c0A+zzFCVI0eZ6iPCye56JN2j7aoz
omSCEfN4Qj0cN1t0WpmCcK5+RCUvpcN651L/OJfG/rGCzYqLo5RWZKl/OKYs/0/6
9EELbBwDaz6V/At/6Act2UCH62O7ZaMZnCmGuXQt/w/bD0b6f9zZtQ/a58QABAs+
gI7hwzsQShVGLpq0QvYRJNDIT2zVPX2g1ZGSQb4EoFQA+mw0Y8RPyHsPlYVCVoUs
obDv5cZAYJCmj28pRb0P35gKqR+TCXkRVXGv5aMz8BZSBgpshzj17h3UXk1Y3UbK
RnKRlc3eUgzYs7yfTs3LQ8Fj7koEpf93NLt0LsJcnslOqsotZO4ZFkw0COd37WQT
BvOPy88JY9WZ98Mp142jKfY22O/EKihSpEPts1tUMx+W4qFvb+yAyVf0Cu6XrobA
4wJJs9n9ZR2PPujWqfJyEnoUnxVqsK3407Q2cQasIsXLoOnG+qJf7clQyJmC/Lxm
onlvXxnsI5i1mTERBgmOtyH+wfZqrn0r/Jo6sm1itOSQeWVblfMWGexL9citTBFA
9l7xSgnDqGcIQfhFIJM4KEQwqABruOWJlguZhgaG80WSWy5+PKFQrCNUZAzANEw9
p4kJyOw4czemuH9uAeQdejv4Z2XnwzolriN0IZL2ciDH2mrl3l1+BJrteoCzLYcJ
blFKnllWf8pvj/CQf/EpJDOU2vGbuNQIvafHU9Hs8gmaXaMkjIYBw7DUjwuGlJq5
v4icXC5eLCVeG6ghw+V/g34I8Ava0AOph/UPikCGl/Hv57LlIl01+AYhxWKpXhLx
W00Gs+luDEDSoxPF6NTRw+jgaF1hMwE9aYbpiTXip8rXPNzkE1wP1LogsjV0fNlm
rkHqguE5B1gSN3Nsh1tBgfRzoEf3wqT+FtE4+wjCl3rD1121nzXzBLsCTcwukTKg
ArXNf1yyCISt803SCVX5a3jmngmJXY3Ryw1gCZZo7QwzmpTjR6NHSoJegvm9uNOL
OafFPE8xbhiaANaw6XH3ZRAqWhQNltXiN08YCD0Ooi/J5B9sbVDHd8Mz/HovFBUu
hmMhrJ8BXJkTWOwZY8v8fXc61dWHK+ny33FIMtSu8sNWSiT0H9FLMKBf2A87I5Sk
QDubuVlUwcjn+uDjGuEF7hkxvAuoy5FKTYiPn8YvP0qMwlDgfPlR2PMDBe4TKki2
/y4t/VQYwu3kJ63adC5QpYvjOEci9g+PkGQxLDvK65LmosuSdp4P1PQnBMh10raX
6V9My+Uj4YxBiXxASufqAp00T1YZienCtQq1Z3z1Q75A9+RquYQwkFWDmLsY+yUZ
r8+J4UeYCWWZaHDllAFK71mlohhsPhWKVLS/L+y+nFp4g4QmLK2HXNMCVLXpDUSq
R+VlwEkQ8uz3EBcLzOUR8M+bllg4hvrFYMqQEHavQGOGG4hsxQET3CTWvmEfHyEl
qLOHnSBjDR2TYUnk4nFBTPRYrw2Ij74gZ8BnMpi38SHAfBwlDwqpWZji8DERyvpp
xRlPRhcaebFIGm8sZoTweDBWhxwCPpCaBde9ZM+MFLqrgfX0T33PotSB2kfGJBSJ
0UlRoOINRZkFERFC39tUYhGSamoijUA/Lc/jJvpf7b+eIPmwUi4AFHOgIXUr71XP
KoYRCByf9HGvhhpMPBgaK8ZrsfxjOh3Y9i6fNCsGqM3994AROX8UG+7sopvBQZcv
xyq02wtXVCi3E3C8H+nIzgzo22faZFdQT9oqnHafpFYJHnzctLydhoKrjVxXg9tq
5jbZqGh4f1H/g+vOahX5cmdnOayHNByxcT0qQsKR3efuXGtDWc4rmEox1cOMyueC
hB4/8Wqw7/+pZ6JfkGiy2uY7K4f+CjogLxYkKde3jVjkNXWEIUlHWnG+jWNch+hR
dusavVMOaStKpKnMPQp2aVihzA21x3JwEUul1Fl1ZsjXvyQfc64R9efdOzmNtAPv
qJ3pZFrELRCPq5hvcDvtMKex2fwFGph2+9PFVuS0yGSXkSt3miJwojiO5Hv1R4/g
s3NH4FQq2qxx4ZyiMfr8SUhPAbVoNTigXBWWOiGuio5LVXURAuLZryipWbiArEnL
KgiFaOj+ubn148jQOdQXIrKdgwjE6Zb6lFOwfylwlYO/ony1KTvUGi9HSfCc8bKN
tCYsRjvYoA/YQwsDppAv5pO+HEaCViXdHzkDRAFOiYeHMGA7KA1E0NeYqoU6RTMG
6BzzfnpIGGjU3n0HSpyDIxk8xsZ079HoxZ6z58tbCCm+I9SeeYM43vLitHf6oo5H
7j1PIPfDbgRkbp2FK7VWXPSh0NwNWVPvqhRqd3KX4q9JhBCYpcykYgWv0s/JC4F7
dVdO9AzQm1rCfk8YTYqWneq8ymTZxiv2o7WHTdImaXOeBFhbgUKa+DtLWZQiEC2k
B3aHhyVdAjR5vyDKQgtAcGyr6/MTIeYffPJC4whNdaCmXw8+xNRuwr5heAkq+gRG
POXaWn7jcPAkMkY7JQtwb1hIpUBbRFY6QnvOn2sHegHAgEePScj+MIMfmqWdlm2W
7lNOBqCc20phdh5Q4DFFPd2vk9gQMq9JJ6UVgJycNvgjz7iDEOQpoG8rfdyVsQOg
F3VuROjKQZFUhYVQaFBmvY+hnxaQfQmRGW9c2r4wwXKy14N6r9mXbBNokyx/gBep
HhtQJg5jZPqWdDPNmwVEkKNHwMDOdwa5g+PE/iFnUPhQpmv875wbfOF53i8Uln7E
JODSnWX+7yYb7YA/MyWxqK4q1gN6bjiGubicjausSoURBSiqxLFbNkdD+rCpBq1k
ElE6BQr84UUNGayBReR8NwZc6xcqMfi6zc2R9G7C7OMayHuZ7xfDq17SvD8TSFN1
fqNqKrIRejHyZDzAqkBt0MarL3XjT+R7r6wedN9S3YK81trFE9yf1MrUiTSALOuS
p+xlfuaYSo17gMHwyjoUpYvX3ZGUKRs77YQ620qV3lR+21It6H5w3z1rhaEpGbL5
TW5lK5nNee/JkbrZsuqNlq6jbQqkLqYK8KXcyot+4oAlOn/zR7fhi4g5GqxBzAbN
bGh3SthGBwByo4QEiSh9/jEwK9wZvNQCchcpKaGYPR10ZiMs290N27aznqXq0hSW
yNDaUGI6qjMHB4RlBFlpufWAZFZ2NQALEYWWMFEkQQDM1AQDZDO5Fhdv/hGjEGsz
FBG+RYcJyLBKaHnvj6zxbygB1bogrGoswKVh2cmDZrk0eGJKJDiNbE/NPj3Ku/bP
m9CBFkAi6NRAy8bSTgYz4PXqAkZdfFwj5YgL/MQ++Lt4GUITobmtgv7WPBRbIb2S
cie3wT09Or9/Zy07UA70ejo3raxZhLyrKrxrRbTTtfw8+XaMOGhbuKlnnS4dw3Bd
eHqP9ZAZalzXTEbPmNjj5RmoF3tubO40k79p6A8Q9eHHZnWNFznTeWiJZkUbNlcs
D+lYJWnqivWgiX6mqEtvwQ8iPkeZ6ITHLUhqLxnF2i1OE6451okZooTmcIpk3okZ
FMitxyBBZWMzmgHHyRT0QqaA+tLGMPiFEVzUpUDplmT7yk6p3m7ylnlIO/lHHKhR
4RVwiI2Eb/3jEvQip4RyoKFHj3GfWTze6XuhJ8O1erNQ54UReT97S07CIjoGzdBz
ArexAQUwYWxJ8NsnHQiZLN+o/rar41dY1J7Is/+SIu4uqqaehpIC18cxOPXTv9Er
VvCQ6XGy9IE6MJdFo6fbsG/WkqFJuFcTcsM6BI0Tu11v9bZA4D+49GHCH03q9ODh
a2XDJscjXDyYQ3ugHFlwly4vpjJpFliYMVNp41HWR2uiUwARgIJrzWVPEbUOvycT
8zTXX0JQnQhWX7LMmueRQv+y3dbUjR7IyR34sVfNAK/yH9tagLSB+LtsASWfEZFz
FN4l2tPR9sex8DA8x3Y34lq5ETa4MMlirsiMCaM/uFVOKjmo+jpZwl1f7O12JqqO
F0lyK2jY9+f/YuHom5uP/tSMI26/Wy9tikGCaY+C9E3Nzcfi6PHRS/N2JrPiZz9/
Lk5wMxuvcSb7QNASPbnnZOA0tqEFU/FLfhE1QrRpneT3QsonKCLtVWkuDJcD5Nhf
fKiReU7014cYHFaYKNdVZhW4sjJxQNcRkUojUd/d1sBhnDgbSbe0p06SgbwMDh+L
5Tv5zAQDCCnUPnfNQJT90MM7ZQ6H0uPTIjAKQ0p+xkGv2F9hF2Xpmv4lkyeA04T6
N3uWodc5V4NXna+OY1GNlU/Mo5SZKQJvfjc7JAV7KpirS71gQeTEf/puEkd+WLM6
rtIdGBo3sI6cxeR+rFPitXPxPOSIm6MhSmKN5Hf9bzOWw1zr+kWaisspAe5K2hD3
TNOA05jcMiwvmbntIIcp4VIMZ/6orbNHPkE+9S18wuf9DWUxBrYMDVZrwASXZSBl
8yFY3xrr+i76D6/2xfAiU3kZgNLBqNA3ImCNzUaw/Iqb9Vom6RuBJx5p+74g0hqB
HWYuyZpz4vb3nsxDTolb7UX+OJq02ISMmn3Xkx75+pHP+y/Kr48KUIoQ3APwNdcg
/PqxpHkjXh9I3treEhNSz0lZTZmGu63kRpAejxcRIKElL9/ABV0INTsyh4ZGNWza
QRXTCUT03sghkvoZQ78iSQ1CEZENGKoDpwid0Wyxy0qh9BIQ3n0+xn68ZQhQIgVP
xpZGa4LriSGE+1OYa/BWoNbqd13lIzIgK2iAbxJ4V/PsmIPzWfnqR41wkZfkIyDd
DCuSBXR9yz/vzqqDlTltqrt5gKl7KMFdfSpO+WYMwCWeBGTwm2GP7R/MEqR6DAXg
YlYvBuEIs+nJe4nOMxdhtCX+q6Gl7Spn8M50Mbus/63EQ8Fu8/qVU1v/29AI9W+m
33rTZYwESoOQCM7D9qEjmTdT/erv8cQltFipH0EjtDlHVaeJo36hdurW0DI7Hfcc
0dK5beed2W6E43UTVnbPl7x86NSsVpTmwdqSoSrOpYKZ4cOas9Jw4v7YYrRvwiCx
t/A4yi2EH2ubWfJd6pRFg/LpZ993RmVjS3HiOj/lCAGtktE2vYbj3HgnyTPySczl
PTmOvGWOtabxuI4U5+q0fIMgCp2MeMA/zomwX55Cf4P4FHM+bmdF+fFcyzh89LF3
EQ2az/ztMXjNsnSiexlKmNIw9U9jIIamgdwu/4OlKhLdhEN9nKpJnldQV55gOaTM
Yl20iU0gLk0cO6gDFrJ8CxiCr/eeOO9LGJDCnTcudNj2E7ryDq/Oo4XzmqwwNLrQ
fEyKY9wYMSK5UxDq/vkXSEAmRUkDJeZL3T8MFvHq7O8QZ5d4v1fS19N/+k6cKOiO
fIbflTsKg86I2EUzD71fYhO11BxWkPkh+7wXbYTkEmm73+RYiPjWn7PzGNVGHBWR
28L1pAU1HruCggkhE0Q+zJQmv2O44BKywx8rTxa1r+873Q63oyx/fqrE64H4otaG
b4bOvTM7Y8saO6vvR6apG8fjtbN5yiAQ+/XSgKuLocmBaQyfyEB8hqkGy3kP64oR
3mKRXVGadwfvSUVeaKg63zc6kKLBzrbONEmvwMYCdbSL10HvcnmukBY5w0pb1u4z
ph/tvluszGzfVigbv2R942GnpvoqtR3ivBaklP0ugOGanPmOdcXw1g/gnWDCAkKB
G7QUELnf3Ax3+xdpRT5fM0G6dsuOLuMY0VAkWNuexh52Vz5AV2Pzz4wBW7VJeYIZ
l2d823RD+xxEMchZmyKw/Ngeazb3jKqs0MNLU+Ai0R3VgcLmWdIECdDkVTcoYETj
WKaOOwA1GeBsocj+y041hCp7Oc4NPuXYaEo3tw5ZPxf36ZzullI5Rtj84YBlas7D
xBuDb3B0c/8z3ABaOBnAoIu6EsNEZjGwCjN+P6TzAi5fiZiyrtBEsB+c8acWd+QQ
PSzlNfvLh5tyaihLPIDT2jYKTZxPi+w5B87y61Bohp6TRMUEMfwj1t8LosyKHo4X
Vs3KJuDOdct8prcxbz092jxgQaK2lnuwg4dlBKZZUdwnSBv6rbZ+IPdq3fW/SoOX
n7G8+LtDRfJ+4uJ7osp8py1+c1iBzegxlv72bKvIgV6dVpGQdVp/xQJNrwqRwoES
52wrvvz1ySVavie9aYAisUmL7txF9l8nhHYobZaKkQs0n2geAgSbC1UDJTt+KkiW
okn3Y6F5EfafQmPwdUnS7Sdvq6eRzJMQEW9D2l30xkX4wGar6XrDs4Hn2TPk/8Yy
CyKZDT0SKG79SIpkRpt8ob0k1B/i28Ff+vUAtrNFH8Lc5BkkUm7aSenDvjCSjHLL
HXxj3xxa4QQ+sxpgBkkpkEcVyEIS1mTEn3Ioq5W3DtqpPmEa4sbHlU9RYLQ97KSD
oY067zWFrEmlAnMOhlOB2Ert3fUQYtYectL1q6asUGA0qHlb2u3r2RjeyFOdW5nM
vyXzA3tabpCxH+MzmJyPjKXQBgMb+SnO8/rwCkC2kKxPKb9mf7JmCLCMeiPQ6/Mv
U3YBd9mDXCNbST/jzr7r/t0cGjd7jpMIdcfZMzYyM17Pwr1uQ/HGZPuPN+JgROxu
/8AU/R/bbS//R6fS4klSEnh1ztiU9z4Q5Lo/KJ+OZvfwifEODfbf9EUjSu+Z8q6P
IM55H7F2pC+t+UIczyCodvw7Nu1nGIOAZNMIn4obAqG/CyG3yOTOks8qOiccMmsM
AUlucMgMaVtN0Zjt8Y4wOYfaR7Je2obB7hFNj5NQhjFQUK+O3VxQ+AOJMx7/O7gn
GcEcn0FZPORTak0oWoSEzL4Y35eL40EkYJ5PmhhYBCzE5XrvHLSfUDM2tc2jhmY4
MtnvzdYyrUm2QN+OpdwXfIPHqS12YrS+liSM8IPYHJAWnK1EQdoF5Y11cqAKSa8j
Xp8W3fLTbZy/aE/+pslpj3NCEzp9XNjVjUaeuG6UIl1BnKmXGt8SdHAUU+zD5Qnf
NX2ZKmQVtYKf44p7YWCWBXXKAIstcCscPpw62PonOSaT0HChEqCBtS1ikKq2sYSi
4U4/9J5zHAW/I9oQst9sz6Z4ZhAEuz2fsE1M7uk1XiYfZAdsiVSbqrfglGSSBk/4
XGvynP6X700WQ2oskAknesk01zCOz7loO4kTpioAaLSQpSPvUQBNXUWf7wFILanB
TWw9v6mLrzVDw6UB/YyPjFyA+3fCcD7F+rxJc2XyI9SO2Hk5CF8q1cfC8gCLttkK
0WbjUVQj5fhDwdg/aH1VYT4vtUZzZICyis/o60oHlCDbF7QHUHWxae5d/IvTGUPl
+RQj/Lo2eR0uWptaJNNsswQdtn6KvScyun/8jfF6PuAcvMfUA172e+6Kjkx3WClN
Q/9UNq1eo/FKa2E8oe4B/9Z1QmrdTK+AyWBaz3xHA2BVhkkM+dKpbrSNyudgRk+g
VY1w8OY1bkkm+5WL/9BFTQlf24NFP3P2/kQ1/j9VsBUT/nlBlvrInma9x9O1bGK5
F/QoayhXOSi/HDUxXry5wRTuXUHX+zFoW/qVqV43QiFqESrKbn0bCvg3TLnfrCLj
UBrY1bSz2FicgvCk0EpHqYmce+U+x1YTMBnydLUhWVVFjCpnWZghzILb5uL/UYwz
vLXaosr5t6Xtj1OXrt+1jPxa3qe/qC+2/f/QPDY2UgfFK8K/LfiGhxCnJXDWkeSw
aA3y6kVZkBRpqeWAASsF+Hou8kEp1WdbwXD1oSWTV1VULHCCNtgIdEyXCWjzoOCb
VH+g9F1GbVKWjNp4kt9gwvCT5olfWp2GkZfrBasGZ+HFyJj4TXOJ0JWwc904LYau
8Qy/Wrbjwa5hU9dSem+njSyEfl1hox3+M2y1BPU5wYLh2z6YIyLsI2cwKQziNKo+
lLi1RXyFTlXMncJSXT90SEX6+4F0wS9LP2zOF5fCqBx1bX67K3mQmpcf2BCsptnx
YjsxAan1NKe4HkkVgytImvsMK4oLNRuFfLZBc+1M3Qgjvu1S48yEn6Vk+UhgJHoB
ycPXYMY0/pQ/hh1lkNlcVMJwJ8hsv29L9/N/sv50Kyq8DniiQLbwaDfR/DgVJHuP
woCBMylwo3pYtJLbzIzfuCaxVUsOoSzhuZqNQtRlc86sp/ZDo10S3wMyf+zrdtGq
9v2U3ANnHoJgjYQOSmVgMTGhNUbVPg2j5Ohs49cnqM0ZH7oVrmmqU9+eROF5eH9f
b2Y9W9oLAlEWq2uc14Ui8Klj9khBgcgAAZqKru0Da/MzlquF2X0v0gILnXpVJwaN
6DN1nX+OqPkjUn4ZrwtKzCCYzha5SbFLN2/ZWsk4jF1Xy+uFS0p+6pApBJlxrjZ3
i/QzuCPV1SpVkK2chqBfklEh8GeBuCAg6BPqKZr9dMsLupjLbvZ0BPAWc++Qqbtl
yE6U8hu8eK+hIIrABBK6jUFiSK3VD6UVeVd+dzb4YUp98rBUhcaoJADPBCqz/sS1
eXJiSpomlx034aA4kZCX+y6avlMbVSk29PtRq7BkPLSMZsARMq7qWKIQk/fkCmdF
uloNyqhIVO+WH8Is+JqYZ8ZCiLapdIVlsKrfDeTGqK5UE6yrWNDRcqU5AiD5DIfd
uJBDh9kCL3eG0TlMnFK6efCISUq0kZABEbPiDJffNMbMjBrRbPAssoQd6nU8FEtU
VhosQpjuJP17DEVTi6FEDbh/R+8r2eZq/0JClRM6Q/DwBROXBKwrt1HSmFr6/4KH
/Mc2LdangVi8EzbmA9EAfueCIFDABlGR20hNHNHL2YrQjvCkkkTQmkahC8+7flHa
AnQZ68tstTwTB/r2d4ROBc7XQa8LRDPuInOMAMxC8J1BFCZm0NwoKOkH+Zh65WVr
sc4/FW3gRnidrgo036pWCUbVrakIYMrvkqWLUcvFE50FLLYFsCee5BzQX1VXbK4v
ywm1rIU+tunO71pTa6ktwt+FxjeR0RFokwBGcRNoQ79vpldsNLjNmcGgrv1RgCgg
AxetsUV/krYoKFKyGlMktEqMQ4pWoOjwjflKvjo8Oogd0QSjcMoocHgIwGV0Q+4q
+Hcn3O/mokgMXn6MVSYdrlnqwO65BfPaWbC+Ed14Od97rECOK8gxcBaV0BHPRaYj
ut6Uy5bpo6wbPtI5QhudZfUhhuhHxwsPzxqahlsr2EBLehBNZEmp+MDhk/UQWKeE
v/Dfydp/SomVB1RvTHarCHiGpxbZjaQYS9ff3aaRH5ZDTKCPcfCfJ9SRtG50IDOj
JjdvedqQ1T/aDPB4O86f3fLhGeJl//2S2k/450joI+ekQZdsACL8QgWVloKW7u5M
rr2YCnDjWkR0YzjgKJFFqOCc+arntuHGGoWuzS86vcMeiyJnSqRtjswQCS0PMJqM
azZqbwyY8x2UbC+89Hc9q61jb4jiluTz08MsS1kheLPp14CoZHxFv/2BRNbi0Lxb
UHo4JYS2J3Qg7LH9sd0oB6bIHocRDSghrClcrv6KI/NqI9WS2gvRIgSCAmMRN5n6
CHLLk0QTbLOavA4MSlaSzRMYPfoqHVHruoIOJuJU9M9Jid3o4EMpWsMyh6nFXf6f
E/mUxQjIFGieOJiyaJZn865F3GuRvYLqPwDDb10esMIU0959tfpN1djjhYCkhY6P
U0JYvzFQv4gFtd4HLudG9RBHqQnhzUStpBuxwJN47mMPSpQhx5k078C+imICX3SV
dQ3o9i0HEWYyrdwx5vPr1z8AHyB7LcH+nZk6i2CS7niui0VCyJY/cyC7NLm5Ub1p
wG4xClhMKKHtoA23F+VeTCB+Zwcjdb9I/7DCrehJdQxdQmjR8V8UhL3O8YArEyOp
31lgccWoC0ML0jkAinJ6JjUqyAb/4fOfE+9WyUmn87iDhiXTW1X78eEptPI4Amsn
TTG2Bc44Q6y6IHCVOAmPPKAm7P9QFCFRVhMfMrfZVfuquA9uy/WWOEJtkCXNc612
O9+qrAtlfKC7nJP0EkLOQSC/zQ1m6nbdWU1T3/79/j1PJY+dDd0MVo2d87RPIEdm
PrSohKr1LjWguX6LMivNfbTRbb56nWkwN/+Pur4ouhEVWo1u67427/FdPCSCmPOp
mId+H34utPAom2Svoe/BGDgRl48gFUuARf9eS/1ATP8BctXb4roan/yi8icOtzDD
YFRD2v1lMxUW7Poer/I86Uj6pE4fPUADzpxrvr1q0C/Cjdm3/RNgqLtCrYKWDbwn
QRPKZWl4CsZ3UmUs7RFVgzr3GnZtYG6+C+c9jmQKcIp5snqg8SD1xqFq4wKFXBFR
1ZpHIReU50DEqifSeUn+YzIS5Ulz2GTXUGSldypdbfOxVszbH4vTS7MvDJPnCXXq
Ymt8ssNBNxU6evkuB3dgcDpwiLbMF15z5kW3A6/+m4tIRTHbuCeb8xCQsGB9A9n9
3fdQE4UdvSRS+pLZlypYA9l82Rs2iI2fJqZrkzdUxufpo11Wv7d2PB0BEMo2gwnh
mkFsa6/qnqJI4Mg4cCKIbkfJQt5Qp+cmjqd2RM/YMen3b1qrZ6fKWHuZkuBH4eUi
2xmUekRVpWBzVVhjPW6YQ5CoKifoAZWhXpXWbaMoGvHOWvZF1suNM7ta0cVrG0Ic
9ekpFT0ra9OiOT/ILIgA5juSoVRRJEe11nOaUCQnYF1o71QEcI+T9iOWsvogv2UI
4offtfyVtQxBngdNnmWsx3rfiq61/K4sIiXqJ7tircKct9R1+sRuOQuDdeIr4hmU
3HBgzkt0pibQDM6GiW4/M/abvkpZd21wxpEDqCA0/u/HYPJyb+s79bQDzujpFvIu
wBwKSQSRE/laMB8uTv0zvN4bt2iC1aYtT6aRBZOg8nvSMqlTEXHd1syIOgh/jvWJ
WvW2wk6lWCO7QOTrektNVxoezvFJIJTeKILOiI8VOKuDY00eYS5bvu+W917FR8M0
FdDjznBP+mfySgS+L54DlwS0uCpR/nb3jSvLvoPVYjFX07ntNhHCQd7xq/rLdfpg
BzCrUSa8sW1E5wSHeXabbAfJ75j/j00R1yiliOnR90vpV5f6itjpppeXO4SfNLmR
aFDGD1hwUgg7zGxpR5IyUp7PPhWDMOQKbPBBH22tvuF7ortNj787PmTe9RK+LBPg
qiuyvFm1rSsDVCBR+GCHiYfO3NEf/ooSc4e8YMFZAztc1qaFNMLooMgBY4Yz7/it
uGOjJJRnqyXhTqzF98ZytPQ/8ShikpEgNOteMggZ018JcYw3qY0u5cFsFeKd1Z+e
FBJkgxNd9MVStlOn7EbC9gcUePo5/ooS/sN9tXXY9xkzD0rW2sr2O5XDJW3ctkrS
O1OGqnWiWF6F006a4gREuADM281h5DSDPudE4oHmyIeOjD+k0bYcU9qwThVvw6Hw
5jj/rVfXjzVEBQ2PR+/hAJiY/bXGqCmBnUvAJLQF2BbnlnJjJ+2p38187q/un8nG
N4r3F83FkCIQwh5xsR70kChJ03cTmrIKb4jsnlRyBytjLYBXBJCpBioOpSQPpXhg
nshtzR0nBuis/ADITvt0bb4dd9/A/qACTl+wQh+HWW39wxaqVDAISwaxlsAc0ugt
BMH7mmLofO0OCiMwuZywXDAzDLjQ42XfwWSenPFrqq+eREa87tn3KFcCbPRC6LaO
EFnTDvDyQbAr1v37QrmalPhlmriOzzJpaE93MG+WsVTcV6xxDiKBcyefJsxxv05+
9EOfO7lQXVbLiDyYF30hPQzhcvuNSJJTnNKlpCg9uQ2D3cJlzMyJzFBdyJtmIc2j
2HyWhDvoOWM2PmiVRuvBSzXsWnVOHNl59Zx5f2IRUV0HFT0Za/dhb95LYEnW5yyP
7EyBhgN6GQY/HVHi4oWawCf+ziQ5wzv/EtcSVeWein0Jo3Fy143RkJ26IZiUVLWq
1ts/W4rA/UBEOxfAAT0x4hMaLknAgztewRkfl257LmT33kdHr1fMMU6Jeyb0XvOM
65NwTYkksc6dGAzrsE+mla1GPoDE2XZiL4iC1SRTkqHm9fwqgdYzUyuh3kNvP4V4
EkFwn/UW7WE9UlejcgvsUNcn4DJZXrME2L6PzIansTYlIgOkK5nz9av6iC9aTztJ
18t2GjDqhdJP5IGn+tRi2Fx1+2FFqWmi7923DWSRv7LWgQMjRSk4Dp+lXQAT+Xlx
AcL8YeQ/1zYhXC+2G9V4h2yVsSG+7U3tZYV/f871SHu3GEzPXaeQLFwsCvOESCvS
lU3gGCyUYVI+/VUEgmKa6nrGFS78iM1iblaFz6u4UifjWsiJ0macBB4b+ye/z5GR
b8VOXbpbKFwB4O3XMbwp4uvXk6RMrXfAw3ibhTdta/vNHLL3G++CdGn0deYqIonl
Qnp3XIK8FGlFPOiM49hr9iXqZYosOKrhT6EOoyuPDu5dQcutMVtwmnqMAiX/XpiV
Ra7d4e1oHd0j2/T54pGtZokQ54MSdN8S6v6esBlxN06Z8n4HyRY6rm1qjWi6TpBy
cSp59BX19HjkgokZgiLd/7WWqQUBYouEA3Toq3L03UL07pxdvp7F3juHNJ45D8ga
dsefxLjfCdEmKJ+XSc9GbC4Xqx+fE7kKx5m+CY1+krIjlS42laUR2e3Mlubgi/yj
wRhFM1cmwvz9zt0Oio+lIyM2qQ4AJYyjdfOu7TvvpnTVH93Aq1jASJ4CA8g3BZsX
/SHLSFM8XIMjkyDN2OlevnnV67TXAqbzUkna415Q07yNXUd4p9/PHEiTkaIRA1Tr
o/TvutTxwpLxYp/Ga5YWBv2+gYDmKPl7EbHERjqQ6iWesSXbObmCoFSW2MYYvrHz
Tt+6pF6mYnSOUtCR6+SV1y4dNWRV+rKRbOlVQCLb6VS6OCu0DwADEPbcqTGVSSCi
qE4wagWO2yMmMZ3qHcpVskNHL9PJabHcpOrF+JESk+Gz6kcsvqprQn4u5APKE7k0
rnOLcblFK8RqNDpM6X9ZQ8gI6SobJZZyBF9HYESaEJ1CQ+sWV4652YvCnxBI61bJ
mKPQAmf3V+X3yJ1YT+0mEWf10k8uoyBXa54EZBi5AFYEsoHiEt0EQrDQYm1haKJ+
eOqUL3g1ZknU6RV5sMVl7bzdfk0D++GAVhbS3d15n7HuxRAgS91GvssXxWNj1ATY
S5LzswCmuJBGK2/WbzVYCFS/JcKUk4UstGuQuoZ6SDuMLZKejPlWhU4ZtMXdJpfx
vi1VoetezKkqRclnDFR3tdqswa/SdaWXPYeEZDfwSaWDft59we65njV9OlGlsJze
VDTS5Hiw7EVQVWnYU0Cc6vxL+Lsgg2PT5j/e0FHHy7cfB060Pf6g7wP2MxRx0P++
cognDfwpvddVxdsCTvK8hzJny6Gy7zV7vEwgKKvri/zlCUC2T9+T9q+D28Knxklf
WU/2MLRM+o4VL2bXKd1UvmvKamK2FVVjC3kin1D5VvqFy1alsmFj88u6nRvN4cR1
/+GERF6o3Ht59jN0f79wPJkbEPH3bDndwd88CTVlaGt0aSfbFIofcmciQ1xOGAZZ
7guLDkaJjtZQiqP6kvcjLPnHjJXhiLwEVYo/LMOcw2f1a2N9l1paSPJbj/RTlb9O
R3Ig7jvBBzetR8wgT1OYrVadoI3X4tLZDfBRiXrpy0i2OZa4+uKTvHbvnaiOzNes
mDhSJRPvFPVF1osSI/iKWuOe427epwbVUiyGyaygs9n9akcg6G2r59PRf/BUX2Qz
0CqPcSypCYbN7ZfyStQPY4wKsAXmNoY50sMoeAGNQKJEGrcKnN7NbxdugR3pYFq8
wxJ96JAk6TCsDoy+xxZchIDZfWhyWVbC/3HnWlhkQ5afbWfYATAiMazAAijyjyme
3/OwqQpedbgW8oFeWrEeMbOT6YoLeelcUxH3Gunu7tW/IbfWTjWYlDfqmHFml8Rl
QOhhAffX3DPaqw05tAolTlhgX/mw5uw4VjXdTi8LKjJcC8nsMltmw81rKIMbR9Vc
p0YI6MQBxuxTDpogET9mlSF6dVtBHb2WtrIftt0FG8n/Ohk1ee187coHc/taf35U
vVKcjNTBmjQ3M8+TnrlAzoDqGsaIvr+TdK+TZlSR0RO5ISsjv7DM0CAwTFoMjODD
nn6NprjWJfuf7ypKhBID664KFSAb9mLonoJvt9aMH8Q+shCKWzLpXtjmTY3m3P6N
gbeGtybf72k+AkWhigVttGImgnWhiGm5wQiHjLoeq+7nmm96JbfJq7ftaJfteZPN
TmyezeWyxVxiuRzMikMILB41OkLL7ZCJObx2XsPMTwJnc4GmSTmdcW4i6lkg/K/i
HmzxGgXpFryQ61X5wAhbovzxlJSBZaGzUVvjuzuGKKfkEx7fAmfz+wpomqWByyo/
HNTCEFxF/koBYwlDjlj0hKgvImOvFjpg16QXs3UOhGOYG+T2GxSaYvJpJX2y16zA
xOGrYtk0xHduuiiabznkQZscQQTmbMJ4og2HQGpLvFJYiELukIHKVn090RhbaOqb
GaFx/aShsabOEXTsgqrZiX55rj/l+pdKGybvVNSbIOi1ujacuWFxmtHDqZnkfxhc
nnQKFvZ+Kacwm7S2qwwm5jXn+oRanfKj+JXEIU84YHIOQFIRdxgkGNOjYo2PZ+nz
+wOL293Sct3G6jeMHuGQPx4wetBIzCHpyBE2mONWxDDRTRzL82ijFTtXltQDEPv3
0Do0XzFjNiG9zBw2exXvtfZsOov173WqS2CaDK/ojqjmJAPvL3iEWD3Xyt2lhFGV
1FguDKifQDzK7B1GMikfkOz2Wq4W9JHkaxGy6xeT4j50hd+jIEQz5QfjKloAJLKM
KMKxobeeLZUuadPOYv7H7aYPtecX60xbbBJ0/Ce5uTsJ1gUhsZzYRgEMaX1Pk591
CPMh0HuZoK3DwjuDpYOGHhhs9msJUH9jEgo5XdvjZSX3TNPIpAl97Jh0MzW4a4nf
R1NsbAEXmkLAmHRHOyUgoslWu8t6QPZLpsjKktQJlM9ONXeiDNstFx9ZPi/bYjoc
J81ohq7oC0+JBuLMmTRezIPtz4Qdqzrje7U+d/t9xVXoP89mFb2HQ3SnXRMaIpAB
520cIBUSnB7652aGGt24fZg+tYOJreAN+iDjYKC2XlMo+2+ev4EOV6tuE8O6swa1
AmI9ctQ7LWupdivtOwu3MnEisZ6Q0TXdPb3GyGGQHRnUP9kfncQoKGYTLIDj2Awp
sxaBNxWQ3sZrDzoipDwN87nZ74a+NFzE7v6Ntf0u3+vEyoR0Opmwgsxve73KkkXi
/nVV0HE+Xrm0tWtXRNqvK1+MgaC3KYnRLk7yE+fiHDTdQyzxPnvuBpQrJOGNaEfY
Wi3/zCV5F2u34alE9FO6NxDTFz90rNZvC6TD+H0oZmasRkNMGr0QleBlWUu8qKf7
4CPUSwU73LHYdeiIuEHYwQJbSaGju8WvQJ/gKTQDLW99iksLV27SmozSQjlphcQU
lAigEwpp8bmfF97iWZV5KaUqFfK9EQXa73G8MmCNKjETvGXciI5EqOHnkbspv0RG
3s9Jy1UqJWyceLucFezLKuSRYnco6GmWdlaOT3bHg1JyhTaMGXL7UBZf6C7pO9jE
uuY+Vy4Ec5q+9lgrIdEdK9cECW3aW+SQco2G1jMEd7dwL4enBRdFci7X/gtiDhmy
s67zEQI+vnL817UXtgW3Loyq7HW0M48QZqOAVZFh+NyldDwVazBs0WMU9DjYbHpZ
8LK27N5uKoAevxmee+LI8ujPIyF2xr0m77SAh+fx+w91oa66fm9HYaO/oB4VZLOf
ak4nT8keJ9EAlSmpXJqPzecEmCCTtYT9oAIX7H18akAPSfVOyO5N4YJuSVm1aDuJ
GiWbj5Y/1IScTCgVfvRJbnMZ6tpzLQDbVJyknbQQBRSraO8Qy6BJ/J435xKXdiXF
4QS2+5bAo8QUnagJVAiQCf344AHVIFkAp5apPKH1+6N9ajhyRuTlckmcNX+SwBiX
0Zhrp128Y1n/kfC3wP8NLvXavGXsKhzGKmkpnMzYz/Hv4nPgssAVz41C5CdVVeXl
vzJU7KNR0UGAaSLzJLwc8QpaQZ289ixNCKUCPYxCeThzWNeBzPFpqE0DoZdAPckK
pUyQUiPG7Wu3ev6xYi3nC0pUi/uvRt/fxcQTL0hyUy/fOO+pgRnqHjeUCw/rNgAM
X2ucQv8Yd29P7TGIfwA0K3/8aQ3NeMguNmlABacisY5cPPwxNFhmrZQgSm+ElYt8
FDyjscdE/fzxR8fpDQmbJ96dUa6CwC5AaCfLI3maps47mjTrZixsE5sH4Cawdrni
c/3rw39gnEKnGYNYg3nqzdo68GlBtobjgew3Tzp5g2lyv85mqeryocHNEWCQKd0g
RXx9h0OBhBJmcWKBeXIZCg8wfqQ8gO3+7+BFlUiOtYuIwFT0fascw+TKIJ4vBE/Y
iERkTDHg4ZQpk6ZAe6GFX0jte28kTF3PlS58XjrMKWDdHmw8mcClD86gMYxHDFHj
3VC9ttMgvokxo4NsofZgtgJk+grhnGzMp+KwpuSbhaF/OMMkbXHvh//tzR5v5mjK
BIhO8Dx+/jm/S2F0NT3SMpiq76I12ofJigKRLx6LK+HMuZAe2y5KDbdCIMgGy+kP
twkvDhRLOI5czJ53GFH9SkBzUBpZgG303+sh5L7w02EdIygxCrig2FjqlVM6V8MB
E4Ia5z9ZCYKO7j3oN6bFZ/IUvdXmObZtu0bNf/9kKL9KHpfcnCWH46DrnVi7FkUd
H8w5yB/yvltjbBJWjfw29vYofnyp4XsdOPqD4ubmjbtEQgvFTKt1Kn1JmTCvq+Eu
4tYHLhovYO0nKNag1jsumuYXYIgOzyM/201N8N0uFVu3mEin19QVzfnAXCmGrQrx
8g9P1QPf09lk8mxVdYclRypjCW9pKi6B2gYlrNEKQlkT6TwWDCSWf8yOIOtWTYHc
3+ymyqKGBAlv/Z88IAQ7pecgVJDq9kexQPBTo5sT4JSZkTuXXGwUuJOGS87CbTpJ
DvrkZGlsLl/bZArZ7A/RbBkY8QcahpzOp+7v6FyF/X90HxwoACPaRzTLPr5xkgzJ
sBcoT+oi/k6iUWAtg57PVq+3Idl4t4NVddxw7c5XtBvTXuHXlzSP8B7PeHr8TbxJ
9+S8RWx59D0hTxculhf7hmXMkDusuNVefouf51b/I5UyD6ci324LbiiDB5oPnaR4
sjDJnGrU/O/h1zaNjye1AsCZ2Q2DB+yhbyGBPtFrPMLcO+nqntKZEq6WVV8DsKYc
eg+Ikc9+U7YwQrp6QHQh7jK/8X8elxxU5GFBnfAe2NTMbOaf107/zmkDsneVxUgu
LcxpYtxpstGPpchoue0KYDSwShn7SrLSJNvkrHmQh7oRfFj6avmrBX1L5iyIZU5A
2zQAWDO+4EwQPJPyQFYW+6xP+eZL9wQ5bZBiIfP+pdnBelkSP1iUcQq17hMHzxYX
5AZD8P0eJYLocIXVpZxR5TveRlEFCY+7FEi/p2JQhGb4w9lWID+001C1CrPDVTtS
BCejBk+YOPa34xO4Gs3miZpqC+eq9oWNyioaHfSYQgB4O9mJFAHW69/OB6K7Fbsz
yH5la1z0WsjWr/MyyW7FD8hDiIW4FOq+fTGhxkkVJuz9g9ci4VxSgG963NfwoAS6
a6ukmTUBNzsj9bIbyNSEFQBlI8JeEL+LoQ4W5drhZekr+doXRSHStq8TMypHFNP9
GrqJ5yXEguFpaCNIm6IA7gU5yp/hGl7KoM6yiCxC4+1Ssga3Dh/6l9KfYMM3LPzY
4+aH6X2j0O5qxRtqjN26PaR3L9xpfoB8O+Megvc9lHb3T81cqXyhUpnis+GEhXvR
dli5ERWYxupg5fPF0gFqhMhUt6niawU2LvmIYjjJOdMM2WwizTXA18oqVjQMIzF3
2DbgvjyHMkna+cJaLcfUHHgdvQjFt0T59LWW9HTKzdFSBfdEPCFf8MJYvvn+kVV+
+W6KJ7Ujc7Pycm0H+NvuJjtdQ96NLeJuFt1VJfjSt9Z5nl/7uc7xzUPgOmpPOjKN
arYnto/Y04jCkFb+6VNBQcWUjZcgj621Gw6deWCuMU320rDpFprcIWgbL1vjNi/P
PTbondMVafhDTJNSOU6aA+hpBx1GmcEnM/lK2ZFy1FClY3bjiBWpPY9MX/boPwcV
neZsa7ZVV9Sn1mxhvze1r+aav6an+tUTqR55U10vOjWOTpfTCSWK883F2y8KSAWc
CNe5P9gBhdynWUXHp6iT0DmxxYol1aomgGVTPNnp2j6aap2/e2AJGxAr4jBa7SBt
tqMhF5yHQ1Qp54HBnPsao3aqaLPPMIiI2elw5k7YQFzWN0+itji+oNIK+D77HflM
h2y/+Y3hTS4LmjOse9mwHxnP0SbfESUmsApoO1RHZDqq8t+w+eQR2qrzLeDPMSrn
bGRytvqU9af4IHqU4xuFLviYwD37Um/+qufqt6WmFTASRaFMaSXUtWPcpz+Eh2Rf
n/Qe61/+mHUPN+/GvFxvo6CDxWtEZQsFvRpxMIX0uIaZ9CchVAjid7gF58CfAOKO
mmjD0xaxiK9q50VIixZ7LT7mKAn1wNOJ5Vy6Y9EoW5mSwKZT+Ye0/Qf7LnoDTwIT
z4mThiUduUmPB6opUCPAi6NXJ5MqJOwSsUoYxw9Z03Hb6WikNb2sPbfEHjwbAHyY
KTA4iE7g5IKPuyIagHE4cZFJrA8Y49FLsMZ7U0HpyDOFv/GlrotlVY6/ahDcqs5i
zoQakEqJtHP7kPSn+i8Rk56Of1ZoLWeUnfozndbAWj6VzF65iBNtAgQBuxRdppmN
9SAQ/verm5qjGrp4dALwYYLTtvvuQ5aYO77hz8V+lHhocNOHRid4mikZUdUESgLy
F/5jxeurKj4qfXy3z1fkTMS0Gvwfzh+pWvt+lTyFNAAGkoblBC9L67TmjX3XrXM8
kEchLw8CblalGd/8B56wvAGmoyVq0XJD14IL5MAUjtQigIKzmufveK66tZdTN8Np
0aX3hbQOm3YmzTjutpnlGe8jfb/myclX/ex3X3WZqxlkqBf47Wy1TMjPARxwZqD8
T36UZcjUR11ohQC9qFxQrALDiJ2BFVjvDwEnAiT+PJQ6yYw6C38+bgWTu3TUZlKf
EzCEppXSHspcY2XOAKMcC2dqZ6WHXdaYG4TivjuANDcBKvyMfRvocji2fCa8Xpc+
hF3GLLun2oWCyHlN0+G/tXDpuIRDo3tpJaLjIzQoKI3OrT20I0jquGn1/eUtC9dB
fdyY5Qib+OS4tJd8RhNOnxU7I+MQq0FHo029DznXL6gS9Wh2fT3jGmSok4kdYGu3
ydv0YqCrcpgtJid12X2e41wMbJKzH13T4UPtJQ0d9uV5lDR9zJQh04nDbZPcKIm9
kWqfqj3KPgDBUziEVQcgZUwTomh3T7h7sWm5khQISPaQIQfEi0a4hP/q5mKaEEmp
vfy56djQugLHhUTo+6ZH8g72PJ8dGIAJ9ZuA6CCDdtWaZQeOFSVm5D+KMvoOB5kN
rp+rKcScRKUAIMQeqKNmPg08Rq+T+Fmh8jGnYoQ6LlZ3OE6CkPGZ/peMlVDaOnhI
yZRO8v7GyeLJFLAvru93wR77KXHoW4ZF+jLuTM4PTfejPwKkFx+yo5/T0uU2mkB5
fJeti+VKuaZOh19oeZENJs9K+4RbI1bSDfbc0wTQZHeWhW9bkfCOCtXKMibwsXpC
frNBDweJCByP/kidilHTtQW3u4IplsZWiKFpj+qoYYoRNF3qAVQk34bYC9tz/ztr
9j9GPLAOZjnB+ToOaSSCMlPlFRHhD/xf4GDhfthEEsOiO0oI9hzi7NnvUmJLBLUB
arzQ9B+9aIsp80uwjSK7LDly3liq5SBhtqsC8pj+D/5qV+n0YJdEFvFMoyrBxjfv
NwT3dP9uoXSp+JZsg9PDWmAHhusr2eO6hNm5tR/TWujJqs8wwKm1+ZIv4Ly8GBVy
EvF0VR3HWI4uAMxNE1S12P6/qg8AVY0P2Q85JQFIScQGZNsbbPjrtlSYu4xFLsQ4
zATQFIUB97bj0Z6b5KVXq2kUmC/SOYYpyMSnh+167x9xHiqCiXsU1zpqBHIQTWY8
YsrHUyMX7QklAaQCBDRA8BFsa0neKI8LKFcNh3Y37zrLIIKG2U79Ff4KMm1itxlW
DCHUWzY2tAEcQgKheMa7+TG1/99OENOfFADzgwLWeB5xisSralPEkbWqvxcNhU5u
zHtn5h7r6DhX5fcVS2xEBuCmQgmft2lJa6p/t8Y5moiNpctO/pD+kus+Sw+NBD94
8EHFOyiNY+LsiEeT5EetNkZLd7knZWf5Y8JlRzDUshbdUY5ucBSZzQeSMjvJLdcp
GIbw0P6t0PMMosxtc3m0eNdvExvuZvRjXlCpBb7h2BIQImrLDieBvUXWvyFMZM/j
OmOC7prYWF0Uuzd1ZMODo9MYBS6gDP9SAf5JIdvPGbebPpncreoPKZ0z48uAtBi0
jpzh/YG9bhuXDq1fuN9Lo1OarlnYiuH0TSBYbauzknGyQC0DjmxJEMv/JvKT75mF
xASgQcxLzDcGe9VLByl84WBADMY21QEM3VREm40hIV8clfaDRNEqTW7wGSt+XO+w
6/U8PBvR+0i3pd/U2IAQhWXir/6/08QUmV1D24POMDkkN20CzmBcX7s4NFceQ98X
ZpYpWjJzSI9FlsnHqdlXh723togR3mbIfII0pzxWCZCgRmdeMP35YJFy+WIwqibO
/FXjWuMozmWv4icc3HCVxkEoWcwSyla9af6umNyqpHnlSGMSg5Bfi3H6YDWDbxbn
y5IySYewVCA4+5RiFm5BUwDMiMvKm0hwkiCNUEP5dwaicOONkrMiaE9j2mG//Omv
80iL51X5VB0TY3ax8z8pwvxrGxJRt4J8RwSG0mzEjALv0rCL72RXbzBmh01VPqoK
2v3/duWBkgFcfn+gf6Yp5zFiWQIRhhyudAKs9FcB7x4HoJVDqrcbInOO5+dZCci8
1YZnQ/i8ZpHb+1rnL4JY2TBUwhddNFTWcuQqqr6uHNEyr8hH3nt58zDKrgOkD6mX
YvgCVmjeUuat4CtiKd1w5cnuvN6JT0b0uvYNx4bmjliyzp6LYHnjK3UIQXbI12V1
ze1FT+6efHUzhkt4hMPgBZcFGC07/lFQL/Xa25uwJkTW/8uy7Vl0jWrZeoeoKObq
qvkfHR2hSFeTL6gfiOmUkGzc5akn3r5Rzy/sKfr6D0BZByogn05S0U3XGJkMk9x+
Q1P2Eo61hLthnio5ydW5ob8fV6kkxBcpyyfI2xuPktQ3Lru3Oq2kU80ACNHDlMcU
D7C/VCK3QMrRQafjV3d+4fdoXiW35bL8RWqlVCtcva6/2vj0MV0ZTBttgDsn/ZaB
SYn4t9s8aCwHGJIcAu+mUvFfM3R7jO06ectOuvP9/BGaAoPWDZGM0pv3ghbe7LAN
vSuDbC3ViXHOWSshRO22CA2b+2edsGyp7xvh54JfBfVUk1r8y1cU1Vd41Slmheim
VlPTrXT1ze+54cABWfSCoQGCPLCVGZ3TL5y46PePXOhDJ7S9zQGX6KtcYJfN7gUg
jwHkZPlHDlfeLKgEUnHn5hbTwzky8BPIMPTb0Qp2nH8Cjv1/xmm5eGpHh2tqNNRc
/i8gFIVYywWv7uyTnQ+iYL7VARAh2mrdH5w2DzUr+kcdCH81iVFZQAj0tLnEYhDq
DSSy8YEw4fNPxFgfRVKDEUOGJ3fEaKKKjGAgO4QIsQ8VEj7rcyqeZ35zJ5KJGndw
VWmTEp3NagVSAwMANgLhSG1o/qL4KCoSzphNq8bnhv4PNy3x6UwxXi0kB8kXOxsk
TwW3qhYo+9HYBKte9+jn30VOw7jZ+4vfsIX8Pw0rZRyTOTzYV26GuQR2LfuzXI+D
Vqk4VZls+3mHYII/YnnviNqNvi/XXOX5xpbt/PVgcfJp2ZpgUvaNkARt4ksdoKe6
dZwexqTVMEwuIxRCHXvFtd+4RxDZz3QJg2oXrj4b3doZAOdV94aMtFB7v2++v9lC
V1RAvb4DiJsGmIzf+0cvLHEoB4ZTVE+tWXxnnrbVJJjvwMC655Jocmr11ilUSrzX
C1hR2qSIeq91oz1KAaxwd8rysPsHdSQfwmUMPKZOe6Qu3YhMoT9Fe3CVEFSSqZhX
YdtC7/q+99fdSeviDKmydGQnbOQw6H0fG7u8XXWs/qitGTZgHNEEJSCxS9lj7k58
gCtDZa2OrWse+QO0vp+kQMXfJWk1S1+dsfbflsMK52Gt2s5EGn7xWMKzB0SdGnp9
2Jcrdilrx8gQKkZTHeSFR0GlzzwbKaQqGRdkcmmPZhoL1bdfMHsAjRf80v0klC7T
fm1fEgjMrJveQ1yoaImZpzlyCZe1hCMgHc4UH7BPnBp0jCYnVaFLj4LGIU+vAaIC
xP/DE4BGU53JW4ui7EkQKYxGO89i6F6Um4ic9ZT+xUT1OacWKtzslk1WF8sUx9tF
Cu/w57kPF+SChnEsyJZec/b32YWL83EU9EseEFXqqHWCtzOdgF8xbs+fEkNCqLaB
XLRziuDA0lxbDPjdTI0+vSrIZla2GO7GFBV28KWXZH0I5HM4EtI4+ALC23mYmkYX
yuJX8vmviG5sHiZeTTUBDpxxRYMd+JCooSawhvAHRna/zAhIxLvT8dqxSxu87en2
Dg0QW3BekalWU430mwfNRhQssfEB75j1aUnxGUnSOTxytwxdKk3VvXcPHymvk76V
cleHeP1l4WfSefZS8NQfnreHYyf/V29keOZOwXJL0MlwieU5PSCyZicPxHJStRl6
ha3DV41Y8i2f7Atxuk8csJ6mmg6ye+Xq9f7l4P32HjVCdeCOSs7Q9YeaQcjmLHl6
pUMAcFWij9naAxOK/EP4Am5JX7xW34v0/9fCVP4znB5oWXAXJOmNU5skfOwglaUZ
xQvNIR49zKMZNaT7GsJ/EAHKBJWaKpAIsHr72DZRkwAb3YOoJ8XylBm2f0/F4pz9
hLHwIDfNFLjZIoiW4q0nRbcenSJ6o3SiVSgwF12fUOr4iz0lKQMCkrtYuoUxo5KD
H5SfABHfKRODHsACBPw8EufcwTq0FrlcAnnc/8+81CMJFIh5FSn4kqlnDRWE37IU
jFtRCy7xMq3V1ReDyktXPQ7PPA6rha4+6/dVUT777poS6m7lJCGBvuAG5JTWwjMx
B0fQmHWl0zIcrpLwje20WKDG9Jkx1LDfAtWKOdhOd/hnT7Wn8Fw6fj6wqNQ9h2fo
Vu1Oz7imVQubDz/DOC19Q9rFCAiQf8LvWyuMbgwP9Poq+dXRaWRgaoslRKcgea6P
DMbY7BDriHbU03DhVgcuIf1VD7mdhHlE6j63+3DbvJ64JB+ODKwnFh5QixB9N8qo
rIJWWy/Cn1YICKy3Oxq5KuMq+8YskpShS0BXhxDY8BOS0e1kQoTzosH7KT6IVsbo
4Q0zZsS9gLbIPzz3fnKvpDUo0ekzz1VpFNbWmxAPy/5kheK9sY0ZbWh/CDYtra6R
GeUyA1njtuoswOIK/Ql+bgtkrp+RMqNAc3RGhgD/ucb4SkiCkYs9d+dCcJHCvoEq
D8kuD5Hs+z9UvOsK2EOBIezue+a6U7EkN/qDUHCBJrBJjUaktdf4EpJdUQJAy5n2
34DUuBZTsFt9gD6WFNb7HeJsimf2TqnlcHy2EgRwxPghwd8tdfP9Xlfm2jOukC9E
J7ODH2IINjybtI+HUHh6Vl+VZ5aO3RQXhNtE8ECv4ycWQx9ie4CQhwJ0fSvmCcSP
WUBsQexc/XA8ND4zOt2B8SYUS+EX7Vj6ZzI0gT/S8lzrVd9UF7/2NZsYJfheZltx
30y7oYJK2ro0sALw8Zl2xVgTiWjoFlYk/7tJXidfY5FfZBqAqiBHFjbRxKAIaEqL
TUWiDmUz7r2WTXTOw4+BqXs6njjDCKHXaw/ndVjDoaU1TtR+rRZc8HhmnM5E1hRM
xY5qmM1RGbYbPEyVy5WmFtmZ9k0kAvf/BJRg44/hAI0VFYog79Qv6xkhQ8vLCjpd
MemI9BPrwdtAPNEeYjXLAZtuDTtI+MJahgz+hpr7MT77o3g3hlGy5EkksFnMpyE7
SF3NVKgAywZK4DOS4MCG9dJotFPcLFkCYb14AO00/VdO0zvGs3CR4FNpgsOEetTU
NPDortf2LnCfj7N3wmY4NPq6fm+PBPUhRHX9U1w+3pfBpHIWx8PnC4XypDXxrSHv
qB1SC/s+KmeiNKWN/endBRkT45KUSRutr7m3+rPoJU2kBVgnmQdA+kslPIkgVU4x
//cuGksA9lXGSsgZnIhb3uBR6BjBqata9r63KDf7uuNGCjyJ8ohXbO6Wk0TvCKz/
U75qLRcHrecpYnnVOE02b7w78ZZfZRMyKnp4o6YShikLiRJzT/JROdBRTtr+xtEo
LQ0zIMpYWGuKiYRkTOjzPwmQ8Ped8zmwWqn2weshBaoF1uE/AqyXgJR4oXiT5f/s
xywjYZsveale0cP4KQjPXHx+Bjwj6OHWGY4CKusfJyI3/cBAi8SBifl15FZz7TJZ
9b+KUeOtRcRPUJj+Th9fyEXTRgZ7GBmTPNL7uOZJuRNCelmaB9YAOkM1fivzF8TL
evjlL6KLhd+Airwu8AFxCy3BYjaAniTan0w5NMCNZ1qAWlEOY6s+CHaVY5XDq48P
DXDvtZI8GpmrOKacam/NV52IHcihUrf0GcvOIMtd5Xa1LoH/J42kHzv3Lm7fcYew
y9XjUcSOCWMy7gQPLM64pxsO9akHE5FeKoAu0FTYweHEN20vOtG9XzJs9L0w/e6O
/v2ZIJAYeoSYoNoXughsnoyQcUNBqknZUNoHgYLoBCRrwc0R+5kuzAtnwQz/bgAj
t3MiZmdsGzgUf0GEW09M/4Ilwkz/kxBXLmV2zMyDr9xoHoKIUlifX6lqcDULtsnc
TnJDAI5ImIUOAwYCMntIxqZz06NgQXc52Urr3FpvFO9slQYPXW9FuDPFqs90Ml40
dUooDk+IhMMusJ971/DNmjn3SZpAlRkw/edlC12PPEnUrzXEV3UpVc5a+4Q1mBc6
TFB50VhGUe8HNEyWjpFdNkRCzCT56lUwTzoIDnKyWgYsY8oVUwjziOYjJ9LI5nGr
2nKX1XY61+lv+tC8utCiou/j36Qz5i4hzG0Ojrp1CMWXvQ+uPAh6LNJz2oUzZhAJ
N8nuasz0YvlJ1bPbpjFjBLQkx+2h3vbARRIi3THXXMIotimmBlLuTTQruABNw8ra
yktC+B26w5TBXHj7dCAC0A5CvALgBnS1/KdyUHqaPZMkcYozJbcED+QfekHojccC
fIw89yy+Xkv7AW1RApGIseVz3riVTSyVi2d+BNk865xAG5kCHF6DP1M2ZQpSQwRm
A3LDPS8Ee5D7bgQjclUcWPSxN9ZzDerd29EZaammUlz/FIhJF2OnjIHAHjUoVeoa
WAUsNAma/N82L2LslKZ0raA6MCFf0j0nu5tepyHJJv7j/hImjYTDJj72O3aus3Ig
hi69RBLh/FalWGKIoSiKkXQrZheLbUZ5B33NTHFb7aUXM4Dw/g+ALZJSSGuj3z0R
9zEkkD8xq6IU+uW6dDofcSSaEE9mCRLz6HqxuK/wNe+8TomicNNV9VPjLeWSfFb7
neWY4BkOucqEguKP5y3s6QEvnFmR4v+3Or3Ej9dZveitbD6WousKmbJUD7m9uuZd
bDteZRJOyvX9125PXkTzhZhBBglbz8veNjawhJxI50wnr1WlHSCt6HtlYKuYa+kb
FyQ4+S+8lktQCDdBCll5ZrqXE7KWhbbG9T/fJGWShiOpLzfKIxNJV8RMygQXKM0b
PM4NF3xyA8hfXHEjJfXS5Bt6zkeklEUOF4E0d3AJutRAPzxMkrrfESNrDXwQiz9S
AgJtcQ1J1gJt+qq4oGSFlsudzGiyB12eE66/3agPY6PpS0BUECb1F9vrrDh6bicB
ZsnDSmdNKDY9jvp09Zo1prPwnp6MTiMNJFfcRgeHsosA/XYbVy3RTeXC1Xkjou00
VlGjXZ7PGK5tM+7K4bTjI9gbj74Mc61NZ8yatO6DC79HGo0VF4vHfY0zBE6ilm6G
2NLFwa2mrI4Jgg4YJpePAHqKxvVOguFQEM3vr8uevPxm76QpO7zpB/CIkaSqgLir
qdF5Am5ycmsyTb3ttciGbvXbNkBPjiLS7gHA5GyaZCqfyS6pWG33wVmhrJI0jW5E
BI81+7y6uHKAS5H4aFXpgTzniNcP62rM/DsmGlbsiY+oYZaBzacLQd3ODLKGiCh/
HvpUx5jeCqRKQddaSWN2vAuPODmPcrqsoilY/Zp3Ub9lrmO1scasa1HSWcnIoXnK
ZHrp6qulZfsWukmSjmbxAr6JcmbnOVJA1bXvXCX60xQLuaa8UHN8v62T0imNNrUj
ilOZ8O8GiVZjZixPhBbpamDw0RVP5jsbwP5MvgmYhVEfV19bgt56JH+M+W7HbTPA
fxplZtkvshER4OCcnoOhgRWv6dxybM2WpLaEPYbd7hpUdLALMrAG2W8ztNeZNviJ
9PxWLQl1VLVmeKCFnzeCfw9wPTh+/sITM0sSFFp0d7EVRWwAbxXYR/zFC+iSZnRy
gKq1iYIJcB0WJYYYKLldSUU3RBfsYpz/pijE1m2Oi6p38s4mcl8zmmVhUOV8c98X
0IdVAasx2buB6npfnn+zw55iCwsJ7YIOdGHVOWPNubRl8q1giN8KIyLQvGYu/Xn+
adZdZoVmQsHLEnJ76uJKY6dNFcerU87RWMtnyGPi5MGUnCyiwRev6N1MDR2TTN4N
GBR82qw9V2n5k1ULnR6nbd0qser+P60ozNGDO5fG3esnLVx8ymkSafZ8MQtd147n
7zmh0m6x+lAElOi3hDcumhtY4zMvsNLrPw4X8hCqn4fKsb/mZKXk27ixr97Sa53Q
0BSKasJlgJnpduMC5LdwzsEaVLcx9qKMvejN9wiikKXVrGP7C16jfiLScB0wt6H4
Eaw5DFeqYGmWZLoCEua609DTXduy8R3ZY/F3Z8VGYGD+J0RyTSF+4v9DSlavpFtQ
svfPC7Hr4xttIMz6k6JxFEp2Ld+UkV0PfEHNWqB8bwDMKAZw2FzxhLZMsPCOblYM
i2MutWn7XcZ2RKGWFfMRdjOobeM/sWNfhOpoYern1C/Fn60B30nVJqjl00d3AAsi
wF11eRiZpyc2xv2SCg2WhhACFgEYxApiulPU9YAB2ZF/l+KqSC5H7rpgJZp66Q4w
cJjIdF7DXstGYEl/3ZxUyy0cQy1fm/D3w9SrAh/BviXnwsB6rNg54D0tUgPK0BSL
L2ZnEJ/fds2lhxVBHufI7Qx0Rg4trol8NkwdIaMc4UfklfrtTi1o7tjMJR9bKEun
r93d8WRpkah+OwsNuxe/VdOhfeVI7OfCH9e42NsnsVudkZqSxtXcGS6V/7PC4Sma
HoUkzCY8+gBZIoINIo8zmH/qVYpXD36sonLk7K2PEH/HvDVOXXR+hI28SN5ReYpF
pKSsEl8FY2BIP5XYy+D0AJnjsx9nduRWgfnx2zwiUq/HaSZXO0V69X7d9fag5lTr
4RcKNIqrsSnbKudo4i/4Rx7K605lvPqkq0QjY+uHJoYHjfbfjtAef/gimDRYf45E
zBifKd+dBU1FVN3Hh4l3rfEoMpaoAHUuR3nm9pBJMg03Y2g5vMuHr82bYcVpTyth
feZEqygRJSlXLQ2l+k2ujmTSaAMO2Qrmvk/uiybMkCUwc98+k4dsn86Z8yT39jl9
ca58YgG5ceU6xL1/PGPTej+Uumc/18juQE8doKDq5JqYLeke1ox3bpJzOd68kvlt
/kj1JgugLHjPc2DQ9TuDRot4++w6xIyUiASDGEkJXkz4q4ulw6e31p/rdl15uQSs
kfVVfc6yT2byiCM8UxpGt1MFIQCFSEghW3rya25itRG31bsx8Lh4xM0Op9Us6KWQ
ClIn8CH4F3EEiy8QqaigOeXs6VJ1TIfvyVzWvoxF6lFH0eesK6YO1Zdoy5PqqyNf
LUtoQS7sTQBq4ctdZOhbqJ6GJAbREco5Ew0GVV2CSZLFwt+PNHdVQYexAXUMaQrB
dTi8umDga3Xve+ozbgRkFGtjWCW5wPudeqhD2P4s0Bj9JV8V3ALPGqpeKbuUgIqF
PmzUpxau2ZhQeZGJPAkaLzw2wukrfKF1Je/7yCif6NVU9KuQiIugDhxFcpIeFbJM
TUUNSgkQ6dlOANHggBNH5258yhbJzPxkCcmsyMHSugL7HnDXSRutOiRHkkfndek5
yqyxxt8FOHDDcrHOL942pqFheSm45RSXDtSYXYvLUa72isyzkGyTNVvNxjKay6CN
xa2GtRle2YPQoKsVcKIDoZ8UsoCpimqn+t2S7YxFjvbqtz7cJitxcIHe0xVB0D1F
miMsmS4LxYeChxo7Av2wk9W7ip90GddiCzCXo33c7vnsa2H2tJnN7V7uQcVNl2op
U2ohMmhEYL9UDWE6qjTIDR5psNf9ewDUxDe5Wk9C4vF/ijafhqY/73o2Df0bvqb8
0/DcmEU6ruNudvsXProzIet4tVLRn/rrnDIC3zvGsInurH7yE88HWh42CCtlILU9
jHGqxfpB6HvoRz5SFz3+gNm7h4Vm84yq6VOkeiblM/8b2M4bRWcG6fvbnwq+dAcJ
gPV2GHNooNU68hRML9GmIqU+3Uf2pwkwX4RiCLMU1x2YCbVJTCTGLUJ76eW+dlbq
rA3KShHaAOE0/VBSPr9yr2lUvAR9QQXq3KFcG4kK0VAZT2tSUSxrKlNFLV7FKn9b
ONyqcJ5XwkCW1d6x98Dd5Uilue/IdiYeAtFKmGKLZNfcgkC+xFxh3+vK7cKVaKMm
k5Lw7rlLbbb3cwcplp6Yo6CTrIUFs21yWfN/l0SVCdMUXi+XgjkKWvPFtEHgpVKz
1IRa5q3qzrjptqUAAK9m0K+BAgmOcMp4F0fw9dueOcQGmE5Ym1F2ivrmpTjVrdlH
iljRlmi4xJUJAVYIOO1lkNNwrjESlG/Tu98g1dNIKsDY39sMv79Rdho0ocTC0+if
9sbnTYQ+t+4kIKiYfcE53yHHEBIimhHKTjkkW1qePh5Dt017CUnyB5Dl6Wp3NzMd
U+G1jakVFYyUIOjQoyMWB3kTjGYzS/qDSFLIAut7mRbjnbQZVuJnhqhIO8xfwJuf
IPqtKYtSOQRGh+QsnzMTQA6vTGL2q1yeYQ8PtvuYkIMp0aBgDe0NPYRofoFnHpmG
GZhaqrBo2/6CsKP78SqcLtRPCDQtUYGVGznY1ZRXDwKdJuKSB6mFgk2+T1S+tvHI
cjMjRDNH9vuJg3mNAYQfkOQ+OC6dxXXu65xT+XdHkS6tvcf6phXVVQS7O0Pt+LB3
gjtfEl+BT1Sbf6f42Iug4eBGZtt2zDfx7Tb+7SheMnG8AjbQfyGaLqA0G/Bz10Ew
MlnA9iHKtO5B6ENgY6IS6TxdpsMcglGfJuCnmw6WwLzkSR0LJgU+ZY7cD2bCNmzz
yLCe6TqAXrwqUjBHl/QjQrgpwkMpIvXL+Akxi7lb9IjO8VzlXrRkdClqJHvfiCaX
gscNGgOgdIyfFrJwjy6qsOkg22JlnztUMNg8B4Qmy/QASGHVon1N+7ElfEbQuR6O
xlBB36qiR4DalFSGgWLb9Atilsf2u5MJDov0+b3piC0EteGzD6PibsqbRh/r2r/3
5KBdKxRX/tU0r0XksLSEiX6bv/PJQQCjs2j525LgOLoRhrJvbw7u+iLzmMgjgB2q
3F2bKhAhmvDoINwW5oqrY9lBlwrzhjuhcElpMQfK8oCZzsb99RdC2n7weIXSVcp2
NRLtDQE2Cwr33FfthxgeAn5vhWWVDcSUiaEwKf4tDMMfpN6jMQB+5Z6Lqhpo2l18
RsvD2zxtJ0CmBIlgKgezcrr2goa/++N8rH1bLT0d0Y/5NGswArM5nth329bg4NXY
ZP+0k57zLAH8SYOHbLW2ZfWgaTO8/DXuB4eXP57cghZi6mirpTOV/MQNbKIENc21
8NVA7kUopF4RC6RXvRjLm8dT84TQbGpT7IpLpIym8B6rWFW6j4ITO65vyGfgsfDx
7GBDTw7uZXByiG7ijfSmdBNQXPx/dxhYwOgcW1GON1ClvD66i2JfxI8Pb8bIuLBA
jkv9XdmbwL+Zwp57BVlGWcmfcREthWTc/SA/ss8wpeZGls3v2rzQYhWBi6Es65Jm
xQwlvh5a5lx8hthmsSOo+8FEu7o8gL1LORta0o04Q2A99zQDH8T8VW8Hq3jkdiCf
CkZD9RpG4mxWmXg20UJUj/QZyv2NofB7Zhz/od39jTPScdQups5zWdikIdmzu3CV
DcSBoSsM2Un/62rSzEJBn6Ah4qzqKRXSvm4jTC8gtmvW1q1hFeNNzDHiFepIZVPe
howT66EQjO82LBl+GaoNDalwy0sV3Q21RYR13CFS/++bk+lWsncnSgx7t5kHQDJ1
mmbrcAfAkmZVPWxRZLIFzKiHITiJP0zAhNnmQIsmHNNxB5mWCrRqy5lT7+KlN6aw
evRIkF+4nP5kQH4y86xfnObi/OJD0mcVvOsdLmhQV8jHT9xQgfmtaglfli7shN2z
Q2d30I6hxg33tZZE1BVaZaGYpRkGYyoIn/C2g8qZQArLKyhGQQ6y2UOKCNwn3yFS
jX2+rkvaVK117x7QTIMxOoFSpOw5AQ+yIPzCiBZPMZItheDawzE3W0IOF2DdFnSb
aDZ5jsnYYwZ8vNvruxXAZPZ9clkYxtKgIICLEyMjIQpGmLb/sgDlxTM6nbIKThlx
MNbfswKCbZASXTDEXx7tQYg9xWY++ipzoy0AFurAZo8SLHa10SnJf0gYbcfipjnD
iZnF0MvliMcXU3CjD700weqIW/fEDGhO1iEnXa8DF0flfbyDeVTUs4sz5z0tcRhE
gdpcRXHeG+my+Umv97/ZiqajZCS1V3tdHs7+lkN/smJH4lm+ihORUsfiu2RhnrT0
qfuJzuncZpN3cjaYP5/PjunJCgtM5ExjuFf+bNOYJHT07sAt7q2ctIhpwJ078Ypf
mpGwtMqqCfL+ec8DN4ZM9xHPxLLNwJGT3l/qmLuuEZwn3Ug9nuCqvpqU3F958uHa
nHIzhrXpgUHKqAVUMtxthMcEbHG+UqiNtO0yYDWeZU66iP3i8+oFj3liVlS9bvpC
ziBi1bfWAS8WsRiKzUIIEfuyO4ptMVt58Wh1tBG2uO4uKXSToPtfczwR1xjclulA
z3rDvO2cgpkSNsUeWD1O/3605zGSTj/SaLGxkg49HMPp0I4jkhQg47SfLSJRtjBH
12h4MND50zP/YRzKYNMK2CrZCWpmTxJHL2Trac/bB6GYd6eIvOBQXuCkKwYAhRKr
3c1lG9uCM0eYxWPbe+3uJFdV7JJH9JNCWWqXTeL4DTFBSeB2Aweuz24De+AYN6hy
fkBQKvvRlmU1fZrFENqk49vONPe5GhCvssTUXSSbiwEninsFvNG6IUsoz8cCNfnB
YWgX7L3GbMoNVS4icCB4nzMr1TxkEWFfKdPr9Qik/sg7b9daePgyKNe4v+i9Deji
eBLdb/LuzM0wyCQBaaUXbRX1xlxLW2fvcYqULU/xKAZDFf1SGyewrCwPEIWRFjM4
MigywuWnj1yof4VP1NYeKG5M4IgLVCDr4yrfnYoGAqT1bkqznBh5QErRP0AHXlub
A/u/EYKWH17xYwamUg1bXUroZQ3nJ0W5Pf8v559qWBP8TDC6MRlAislFq1fs7Ag/
o+5+YXUE1C+pBlPaKxdTCXcneZRBDv4ce+lU8Wl7Z0bZrsEv5/4lPelFxoVK8EqW
/78tAfFxLRXbimBrwpuoRBgEV0LnQV2mR5Lp/u8U9PsGW4yuVVcHh+fcTnZd/piY
yFzt8mOWBsgY3Ni+4yUyCEO2M0tql26ZHfJjl5jWW6oKDcWRTyhypwyflRb8xNo6
Rp2qL55Cx307ObjqQaJp2+KNAtxk+LVevfZM46PbA5gY0x8Y68Mj/JRJkPcv8/gk
/5YayWktWKca6jDvfiEE6n1Kghu4/JtKld9PQ5iuKINWUYx8eQmdDd7EDRZQfS+d
k/Ri0Yi+yOVOHV8I+Y6GpGQPzQgse0/B24NsPnAFc3DCwqJXTCMPrrqijB6Q0/qm
Wl7Bj5YJnYsCEGGsrfyjVt7vkayYT2y3lIEiuro+GigKn9td3/jdGK9LJP6RenbM
+aqATIfG37K25jI/cNeZrwQRn6ThtpXwG6lXpen76jO/iMOUiPjnx3M+PoOypkIz
F6YbwXft+Njdr9daT5KBXyJ9OBw0tEvX5frEeHJE7vtaPxsGd4IOwie4faD0LeXZ
prWHZJodX+s7JQczQUJyzR44adJB/gV9SlA+o+BVk6bD3R3u2EiahNhcOBhce2JZ
0ZwEAlsF3/3ipp3GmS+OzKmUMF0va9m14kTRjK74VME2HIfNhUEk7zX5RMUv+BSc
fPrF4bGJep1Em210eZqBS9LFRJO1bsc2Rku2enbWzSS/Ue42RZi81al+302zCyVi
SFSzdyR7j2xh/I4qaUfYxbvakJTUBikuhlwD0unyPsHdlaryvdVEGbb1v4voMzu5
c7ooQiYPTfluOucaUT9iH7/vAppul/Rv4LrvrJIfcr/i+PceN/yaZRPiR18ZlViQ
uvBzNJT8cT4jQkGx8iaSvV2+l4klnixQJs8XqhXbaJ2kmluJElNn77mP5ruwO+RP
6+pmTUDvNo+8kHO+9/xahrxTxrpZkQqEcuN4ao5itagbbzVqPBJrZc67aw7M0QCa
ptE+Q/92Qbg3rGSoczxvhjDAMe2hdRqH3v4mqYd3CM0c2m75WeCRAJB+ibKCHX59
SVVr8Q89PtLV+wDRfAvQHFjoe5hGA6KlIQ2wozVrPcVdhVKk/ENUhXYRBAR8FUkT
1VSARLsehMgwY2W5mcJMtAKP2OArrxaKLovSM1ZUiNIIPBPEuzCWNUX/Y3Cf5q64
a4M1eBPeRzKJtgP+9MnKP1d43UJFkOGk07Jp01bKLR9jeS/5Jl4EWK5eqRt8TMpa
GSoZtuR3asx9VOnTKDGGV22CIxcJCTpUxQTUIn4aFVcRqn9b+NAgMTI3KZmcs0Je
054m6TY7mskP25xA8wQYeyNW14qGc6wrNQBIqwkfexLeQ4Aql+ymkd+bzrl11Jo+
n9sBVMb6jKFUHfN6Lxj5mZC0kGiPAcY49uG1BGFyFaDwDB+LsMVbegIPPaJ1B7NS
EvN6EqbBr3P1QFtdOyf6vh+gsYAXxn3S+w0Vn0A3GV6/RLpQgZGC45EHotQWOmX9
Ile/pL6ZEwEjbSalRo1ePNaifptnQ99h/lS0Z0LJ9s3NO5FEyu+0Yjt/F6brTkSY
Mj6+ls4bjQECqvV82ec5XmoJF0ePaP7My7U60Hy4yQJOIK3Hjn/6II5O8B/ZsDdz
ZQS9H/fTObyUjmdjUXxLsjVQHR1YKgtLzlkib5oczuRjT2eiDiHwe4a+0fSQOr6R
m7hkNrkTqkNdVTQCjWejOrYqeWTO+6EP0IPqOX1Oz13UQYrPJjchJwKYlfWrlMbm
lYqSFMKrxzskRmFf7hrPG5sZvvrppac47oQxvEVLJAedVc6j/UsYAxt6UnV4LbTu
ad33MbnC1jQxqRG7gz59MU6V/KO9RYZWiSLgs7VHiW9Yo05paxjTltTUIVDnR3NV
N7V8ww+bTiGHZhR2gEF+NEB39rR8PCXiG2ugj/oRohONtBHNgkxlywykGWfMDfR+
ySFi3zSwyC04l0fJLV5LxuruwL2F/rOIK824G9qlwkHG7DM+5Hy7siaDClj6yvZ/
zr8msLijcrEVWPt2eba4N4d2TSkFqvE79tfFQiK0BCGeea+Hscz/TKYD6Pgo0GM1
Jj8pJgvrdSHInmhaMcMVCeUG5u70MnwfBs0kM1LJuNFzD49r4Gnf/VvLWkbjRDz0
XZKTX65XJtgZMAld92+r5qC6gN8DmaPFejplohY6YD5oxtO1vB6hbJ8oRpVSLP9y
ARvvNePjeg1uN/TYKF2YGooYVdAp4bI6/zHuilkQC7Maw6bq/Ej/KqWqxOU7f4g8
54b9hOXI/L+oNNI/TipYYibrnB6EzVg5KSSFvYS1tAOIbrMXjroNhJng53gGtqa6
ouYRRDlyGIhL9Gxbkl9JCLrQdQy9TfvjzPI+ceMcfz7pzMk7Eu7pgfqxTkHKPzgZ
ruM7+TXEq4Se9/WBq6+3M6DVvRc3iIJ8KCJ/SfC4AFKaQSHvl6k2YgCN4KvgLkPf
f6No5EfdQeA5OJTFAEctJcd7gSbdGQqJXHAVHxDspS+sq/r5yO6AB1PjFX5s7VLE
5ECoOcL8oBi6hXXlgUng+BtQNK4KDX4p3pRUhjtShSyskxq4anqNLMoZB5X/HyL3
cJfyUp0SAGIMoY1KiEj2VZLLqQCdfwlCHs8O+gpXcH4/8GsyFabeOSLeMEv4PcmY
4FLcpJWPYODfJckr3T94R6iHUp8I55Rq+D+0p4qxgbs+Kp5QrNsJyyOGmVYJle8S
pbL3uF7vJLe/AOCuqjPxV+pqnlAc6zeNTh2oitqNDXP8hMhWQ0JTJSjlf4eFZkg2
yvf5pUjctcBB2e3zzFwBNaBoyalLdgEAS1xPxAwythpRfSHMQd/GdxWtga5YytUp
znk3lbLO7MiAAScsLbN/5cXPfTq6K0BT6NW2ebf5dywfagtN2CysWPcxTDSAgJDg
kln+lpPiZiaGg6uBvDimsOCaKwYKYKrAr8rT2B9nYLYAouKr1esSKH5x24eK3ow+
ouclkP88CeQi8EH8lByVKrZI7azCnyzVJCUKgmSYpIl9Wtz4a5emMdlF+1kep2JE
mgF/RuNWHhMy+GwUFcbIAOGj0fnSAtlWULep5p4g0RIrGqGx+uabjbTsO5eJ0/os
4yGCjzcMuk/TruE4heXgeAcCm51N42XR/iPrsvXn5kxYLuuq4U9TOj5GD9uY0AKG
G0kxqp01PFJyOdXx+NTtBHGWXAe7zvMUjMmV4uQjM51Eh7PsPb1u/x/His41xWI8
r1xC+lDXHjxcTW6j05jvy8zmL/fimqoempjd35qwiP09dbAklGV3MDOIU69+XodS
v85Vw2kK8JE35FF877PnVEh9lCZgVgMpsesXRfqVqPn6rUOYmd7M8qFrH88XYsaQ
pOQNNQnJnP0HLWlrDD0PVkyR59xsCMM26SlXBTKpMkPgwIyKB19bOuV5AkbLLjM9
fHpIMISBSjqsJhXyApHNUdkjq4a8tI6O3szWxIR998GYGo92DLcWRWxidgcSvFTX
eBZjGN3uYnHz5Qc3tO3CnPoZvqrvbLavGjVX0q8OtlgLSNfa1BIbUIUmN0Fnr+ge
yNk7B9S7QHbPQ+YyLnAHkSp55z1i10pK7kEr1lEwBfhrxwIuSix39vO/Fih4bblJ
CLl/KylDxA8jgVyKMwQbhkHmqDRFT9Erl4M5NSwA5iUzvJxL8Qe/PW1RcoVaGumS
7t8BeC1EznZm5yahHmaYWmD7kVwzkCwbBvClfw9Co9EqzKpnR2RSNYSyp7njVuN/
P7RdaskfQil6Xc/bPCUJ+jKRNZGXeygsjepVR8iRaB2CQfcbLU9deX/7WCP1uPeh
i2W12ivYRy+hjgSZ3WkTqLYq7HeTxhAfo5cWaJgLySBGmhEqj2d69Uy6IG/ohzX4
aWTfvlTfZsIoYw+ZXBTJbUJLzyJa5OeDCRXNWiwWBO1yec2ywdyTbMwEbcRdRUYu
zJhC6vYqo3YvJDFVtj4f2tYlTfXeCjbC0KkyuVSNGcTwmTaSQ3IrOZFZC4X0e5L8
nfs5TWXyNyWBarvzk8DlQ5bCjYeyrvwtywRNXof/rhcFZ0F3cuLnMpqy++tcTkFe
/TBtyJ6tWYDoAQkV0D57f3Ubbquu5HXOsCj30c2YBhihz0gQCLJznykCcWo+ysIa
ZIZVWp/bY9XlGyZbZLBapLDbj8fh4IU1NL2FpbKXd8Y4fJfRIUmJTIiNCvDmf12a
a6YGF/nmB/Rp15Q8V9ghkRHfc9JfVlrGNYWJkpAkXGqL36AQeV1US7/jfUDrq/Eg
QgsCceYmsYnVfN30kRJiPIbOoSTllzFJT7tkOr9Uyy3L43jYM3fYreRPaKPeg+gl
Zm1UlEom4OYpdZ0CE8rICX3NE/AJy2NGNFYLwm859Xok8UUHSf82GqxmRWdyqgK2
cNK8nAFcRnNH7K8TOk7NegvuZ8NaaSEN29WzbVGdhtFpRcRJ9T3tnlKdF3g6+iEd
/ryApHQMeGGEuYbsXYVYpyNQvmeDvWgQeUwf12SAsrDf+0DTQzVVgpXS/SstaSIo
cqs3pHyWOcjCgdmcdyF4uJD+BpqQuBUx8yHXH9WNk/W8oyWZB8xYiRX5L6lZjOo+
TO7vjRVTPEVR/Sdm2U1SFDNX6aupOBRP0SMY+AxzHMIZZvWz5B/rqHY9ZdHzD5Q0
mpzavhzJtEG5+4tpHNVZcFdO0rRL3NApanoHnRBBYlUsaAWzBr1jLPc/LQGxstCr
bpnvZSY0berQvWCwWELa3efu9ekEK/grOxRKDooX+wx6Z+lr7H6qUqttONORobMe
msnRa6gKqDcFNUUENJru1rq41k58QOb0DrEFIjO9/nu7dhipAMJlOT2UIOSKFOTn
Zbdwu+oBJnht0dswITFgkyoOHX/h7Q7Pw2BIRnLYHA/GF1YLE5xfV3KHCuuMd4HO
mTa8asFIvNfpxHWalpHdEimibhjXBb6HmJcSr5OV+qcgTMFKLrKPJu3no0z+CiJh
2/D4n9eFp9SxWzo+W/U0osPYg9Z/tY/LEqh1WBeobj0J8py6kleRDTy/qGLicXff
KWFPMrfb/RuO/k46nuMpb8jX8IcDbRsWiDtsNPzUq8v22xXcLFZlX0zzi2TpC5pz
c3/Q72juUKtL5TXMBbm+YvyLaBAezpYnbC5h86VjZNXM9LmI1aB1HYK28QkZM6WU
kkZeLnEG3iok2/XU+iXjvXEWk8kJGsWqgGwjWXcwYgjpiXyufpBOV8kfb9fgKAZt
PaktQBOMl15nMx+FEwnqgjctOOJjJUrqJOkARrzB5StfzOgNys17aQ62U2VeqoYL
SMDll4y6u5NpGP9DIX5rpMGD5Hf7oSmGcnTxGYqp2UeQg29GX9yXjJ+gearIHU5I
K68oIdPCWRj7co9pjOcxzl+naMFgTONd2qonwVK3/htYMo1LkgrEsufEY18fDpvB
fI5CwCRy/VlLIQMUIHXSBgyvaVDy9EhrX9PrDX5+t5JIjjVjO6BrNcRKaRP/5x1A
oj+/JbhVBHOKYmlEZKI8UtRX8tmb+BbAoa1KsFGznI275mATx9N0KUsjQVRW6S/t
4S0wamyi4My6XIo+sPy1ivsvZiLr1veYH/4Dee08pHwHxlvPEFeAejF86vHW1Ms0
fSr5jEbrWZkHjTIF1C/2HuHG685NTCpUSt8o2CVWAhLns/tLvoL/0AUoYcLEIF8L
1utd++wvuypxyLmUlEE38Q+UP42Ah9mMu2k6epwk6zHZGlnIsDntueaqhSkp+Lhq
L8QanrcnqpPOuKvw1v1cn8aFUQ+0IbJynTMP7uWVpMRafkgUcYGt8qQB8EbdNUql
iusL8pkFCt0TIVgeqEYsYe8nVT1t1KdhHfUG8vLdrKm3KjlX6Vjm1hyc7JhTnU3n
m2jwY3jjWA9EHBETHlKLDq14hbaMgmz6gTblGS4W2BhBKUyTJPvmRjuXEf8C+5D1
6PnuqAkmcnfdRgEI7xmV68OkUb9vVXR2/LYLH3LaGQex8271psnZ1jE35a48dkaq
UMHO0B1Qyft3F+CTsOQ0UW0LYlY26fnBzbjSsx3zMJYxVn3TMR5lTUCq7YYXLQcS
DAiF/cdcKcwKBrzV/BH6IGBcsDTMUfDNzZXPiRiJ6Y/+0pMPJqiH1fBtDkJO/zU5
ROmR6topIKo4WIIySZ7aGD8+EzM51Y5aKyJwxcwCh8MLM5aMxfIF7l0u2XP1pPDI
jy+nWvFPcNZ4F7TqyEOhfR/CEP6XMUcjTpX7jcs3PVyKLTVRTzqrbgm73lNHx3zx
gF02Qd5BKrNJn/j0TfdK0cYfk1GSHbG05IPuYRTALnEt0DY6OFEJ2RHvfWA7GWUv
hVOMubD3KgBNMk53VuPbmAAL1t4Y5dXL6vfXZzdOygeFRe3BabvbmvKYzTIXV3PS
skLalnjagHDrzl+iIcnCMwfzelrRipj2UKwFK79Naz3JZFcVatoOeG54/FFBUhMu
5JhCF9HmvY53gTFR07Ca+il+GoPPDyH7Do+bAY6wmIgn6EdRdJ3EN+109YIBKX0p
dH4dl7JyI3TS3SiU5/aMEEPyNP+2N9N/FAbZIO0EJu3dZ+eeTmNf1d9spEJjZRib
V4nI0UuAyVXVCSFJ5Exj6vhPLHGMKm8XoYm7TAwg9gvParHJp2h892Nbx0BWIPFC
ro1kPQ3/v7ZGZECALN4KH77GpNy+dXud72EDWEf/7kV81MAEYUK7YQLPwYB9lc9a
q9ZODIQ8zR0XbkRP+gqNv0rYOfR8bU2Wtkupwe26rtB29vSXeVD8G9v1WH5/pb5l
ushb6XlwQBNzIq678pBlgaWhYGGSM+v+yCMQAgvYJWIrUOtTtrjCUoEmjw3xLxso
WYJw/58G8g6d3fZFQ+UE6skzmsGrB0O3Bi4pajk3L1zEwYENNNo6NDNlxJr5nTP0
Bz1vvR6m9JeiDajyzCo/37YYqlXyk84LpgzJkxrVFQAsPv7CkLfgOvvL1+Us+Gjy
9irVRcF5mT0Sh79DvaX+l0PCmvSQRwyDebJsvN1T6G8KkU0SAX4G30aAAxSEkNO7
cegKj20llWXMdgLcE1mbDSaeOna2zTvi7ysBmL5mQ5PHDkpCQQrRaCTUCLIcQcSI
qa9S9uWG10zqY31pMA1+1mkHvSkXiB6jnQoJj2Tu2Q4RVCTi6LUBNj5poG6Gqozn
gsjVdve1q700JjB/m6Zdjv4Uxet+hCsrEoQTvSGoDqdOhvqd80UdALdim4C9c7W9
LVyJip9z+1DLOCUmV8yQWBNyvzqOCrkaZMOhoZh3YPkZf+L4ClPmLW7wyM+pGB3f
xptCOgkXyASsf4eFj/bTf1/d+5l5kcnKT4E9S1i1ZCCQg1A9BJ0FBRp8InBE6Oci
I2J1saff+9HzwzKdi0s8SeM8eEwZABtfaoS7+CssAJqX1C5ymHBhBHgcwsUTM20h
SvNIWY/KW/c/otcsn2vQHlZvmy3N02lN7FzRegmgqeBPTHYcWApp5cLwn2OGTUm9
L2r+hA5pJH3Pjmaz1r2mgDU1tZKeQJKBoTrwKCErXTOl6oqrlsx2fRSaLQMn3WRy
twc+khfnP+lWB/od36WtgiRB5ePf5c+FOMlM4ZvF8Wvt/ox+z2Vc/RhCLW/ZZDbQ
/hUK1FLP/7I/UnFKFIhAJtZo7vqv5jojcFtvAH94aWmq8WR22V9qJf2ktSzM1NMB
YEpP2i7hPIdvmZaHh9u7HRgwRSFt2Z5sJqurMNIQbeII0NGEklGny0MbXZyIp5d9
XC7hFP7lgQ6ZivzEOEJLvPMDVhClKbCV0QN6xnzJXcgP7w/sALcCHRSAzw1oMxcQ
Qn/3DVY8EUWtS+ooQG5E+7YN23BXaRNSgnQV6jmIKZysq6zmy8VJ5YpYPkGx+6yk
pshn3CVvkJnKM8uGINz7KpZiuNOD/5OUruCgJTCaiKKp4ofyBHiCFUc6cg4Y3HRs
rPq/Eb3l9e/I5IQi9+4G6+1Aa4DZsQ+8PGXl/kiNCAF9+v/SjRaEcyVzcQd7yYZi
+xGZ8dleFH1mY2VGesOpcMN5RFIZhbkV6c4w8j4jU1mNmxVeCtLUawtQwG+J1X+x
mxJenXsIm6DrgjuOQMfWy8GT5EXmaBV5cf4CVKC/5m5C3NMU9dmbdJHyHitfldZf
bdqqez4QHBXVE//nzgUvkK8L2keurE6oM0cdjXm2D3xmSUIr/QRsudvAvptu7pkk
sBtDBGwgGfWRDXNtAxIHb1F554zUdPYx9BlGEQgdQmNxzU3zViF7ZhXF4l1dGQVP
GLVYt+jB/vw0AFOmK5LYGy5f5SBn9J4AkWSSUV/5DNFjrhZGWqnyajX/L36OZWCX
VE0mASnWPIUKhS+wSxxh/AcmZ0nwMBiJneh0YK3jMZPBXCAasXYiCMgaa4ffmSxE
LKJwT2ddkF0a4KvI7A1dJ54o4Mk8sf0gx+nKpacr0Vv2TbQTpkopX8/5mBGT7CTS
u39nH9HTR/VlfMyg745SvV3QnjgagqfFGSgwQDE+5xerRx+cvzsdej/PGUebmOa+
7AvCi7S5MDARIfrQht8hA/wmCVqvf1WGRh00JMgGWiixEOSSS4kLZ5OqUnOSXlmC
jYM5GSH3gBMBOynTSSpJ0OAfATnXqNXJKiBQ5Ph3neM4/2bzBYWO9q2JWVAGHA1b
ukA7eHhATbM/BrLeq/9mojnWzeyqEEctU1GK1oVYscn/qOa1nSb9gex2s0fCNNXi
nFbT9NfNFVRLJQctYHzeVoYHMrqpiUb9rZ+dgj0LQHrCiWw0FLwXhWWm0voOzaij
Dg/29ZvcCiMJ7H5gOLMbMjGCg6Cg3aGHxGjRX5Nu10b3pXG9cq+C+1Alsr7lNZkd
iqwt1QjQ+gXWyC4Y3QWmvD/IuKbPr2Dzh3b43/6jp73fWWeXLM//9mfzbrIBP0wL
zRq7GiLDo/NztcHBPVCFWaGorhebu/L4o+85IAn97wehLVLuvWTGgtw+V8Zp/jm0
ayLyhhx7ko5VOWb526Nyi6CAGSanTvVfAW2mf1D5dIC9bq3LVDeTbTd54xthVH4S
PK6huDGTz7/R5kpvJNxHBWmRYCNx3ZB3pUxu3UsuaVyJVX/10ZfZjPzdr7jjVXlh
jQJaJJIYmZ1lmnJ5hWhwE+QTIO2kAXU7wKID5UebCy/mCLC5vf6xgSZH2ymU1fZ4
W08Bs4IywG1OxrAElVOETmfDSsMuR1XyOfuNpenIzSF7EIOsgcCItJt66MmXLXQO
jXQsyJgFb9Eks3IOgq+kBndIKfyFbANKLbQeP8hSHuJVx7jLkTlbbZDOaNNRZr9z
a61LwEq6XxVc1xFlDT6q8M359WjOU60WZ0fFP0oMznxnQbl+0FlrRxqVUBpmrC5/
9svVFgLBAPZOXjR96dZo4GDjVVunMWgb0+dmnrjD//QTQw00pVIHScANOc8q63/R
6ZP2u3vo6S0PECNB9BF54rUVeyUd//tlXN60Taojug/a14VypdBCshIZhvh66OJQ
if0s0hTKcaPbr414cw+1wrE1m8xi+IZmKp/RK5ZAYtdBR/CyysAuiisM/KYpRx18
wV8ZrkyDko/451mC3J7SmUEO+2vNR1VZc7+7CsMPC7mIgO6iyZf2sNjJEyK0gfL5
b9bS9f1vj2DfQ14QGCd5oMqpGfPNL1+M5kBcOKO3ACCF7l3OF9P23YedE3yYowNi
zIlRjGnuGNHmpYgIHDghzAcmkChrqBG8vpaCj3aqSAKIUXBzw5l3q3SIez4MqgQU
QV8xxvwRYaB9gTt/eLAyM4tXokBilDNFgd8c8oxZKQy0eIifI/dY2T2JKOugIV4T
nBFVZna+dj2/lhe1zR6FMxnAF8duHsGeMg3uKQu+fGIlbdbgPhwwlAUc3KjTRyWe
4PiT5lwmmdsxEmKxNzeAo/BEjPJJeG+p884i9HZ1B8fKO4FGiropm+3Faf7CWkA9
mWFUj/HM1I3HIFPD1qR2UjCVXxUSq37BLIFi1ETdHOofiSNzEGLe9baKV3JzEQCz
Wg0bCOXB+qqPOkrqXxMr0hQLVvZH+WTbPj/wtVU6mw5ci5PvgTGg+ex/rfycFb3s
kGpreIjgKl6hiGF/tp+cYOQoif8iyhvsc93TWD99b1LUsXEzREKZDaTwRjRTJ2CL
jiAh7NSHX0Ge/IGV1igI2So9dWxxOU2lNZEGoL0Grn2QcP4ohM6TeE1lg1dtLVlN
3TroosVSy+ggjfoCJHzRGPW4G772pajtgb5o1iaW8Nre8M5VZlliJ+iWVYq2xTUR
amWcX4GB2aEFzMbPJrBVfnKnG3qovW3YIhmhAbFTiFyUMYVgnOAAuaCMbLnOzCTp
CsfbAbloDBGeEhwqmtbznrAoZL3eaIMBOHOOi38kBOUP04kQntX/qDmKP5NPS/wc
AZtaNFl5g/iyYqaUyDXcOSI36GWPp/rK7bqpHh88l1PolXmTWkTap5c5u1M6X5CY
bFYbayynLx5pGsHhOUZlIyMHTiwygeISc27ssH2+nnNB3ombdJT4O61vb9goqn2E
Vmh6oKzLMCDT06UQFzCp3A9qyb7UF/ISSvb+iP9brEXFjdFQUuAa+QbWrvpddhRL
opD8cDVf6nZjFS0X/aqhVqvn5VzqtC7bvEIbxYY/7JNrdUw4/j3roeMMUQqP5eG8
mQFoo4Fmqc1U7aeld2vJMTjhArB4wn2GtthNznx45vw9MFgzh9+YmG6nDLCJFt78
vK+XRwtRH/WBo5ny7T39Em+IoPNn1om/0CripFC19x/KlLgm23j+K7BJJZosB1p9
K1cv6sRSWJUkAgUD00NJ5yMxuzOS2IskFbhHpbbYbuBTLJXb/vdbft/wyonlenem
eEtswtJG+U/CRaOm3scQ0x4dTIwfLHX6Z6yU1JvbOnc42zLzeHHq0NPXlfGS7SxK
1RCeHRtMR2G5a8pWr88qdOYW3p6Jakmb3A55ZN8LBOHpRomio1Fu8tzCrXojP6gp
5Up9RBMpVvufw1ydSFQfNzAljPnIvZwGue0f9H289/o3WFTYIyezgCAz9H/47kXi
BMEZRWnPEkoYNBPMrnFbkRVYpXMYM7xBv4oFs/4SxXc2gAwskjS643wDpWjiijzJ
9Oz3ohz8ZC0XaPQBJyyvFnExYWczyfsKSrmJGCSIlaKftYQTTaVO/oqCNBdRlKQx
eRlXO3e8dIm3WmrmKbQYegjdwmirX3F2BBPqaTXiGD4pZvUSnyD7Kt9xq5qdMFNs
54BWeAG5cl4jgDL55DsGsQftjvCOSqQ+CiEYxajolILU5jiJys8xpD2viypf+aMZ
lA6P8q2bEum4QbIaLkZCHHtLmDvPJZ5l3yQnBhaKqZZStlBIMvCz5dv/YcrJJi+H
Digh8GgQl8/3vKj4NMvwTcbgNGXAi2Cp1UDqwC71aG4yjlFfVPJrG7B8B4Ly7rZb
lmARK+2yWNQfQ6ywI2Lv1znFar4erEqP9bzNux0JjChIJS5eMpsQzEGScObYETBe
KSKZuQl8CNU1YSn7Lfma0MyQeohA24RATpqWCiopGZh3jI0qGeUT0hO3IXHH4PAh
nY6RNeEndW7x2UetawmbdxYSQ4acAlazFGyw+oFpIj8p71F7HPgnvCHDHBheHwBO
QyE+f/Tc26kWDWaeJRMZmXa4w513uF8hyLPIJrHordizoHw+RBKwLInjTEu1iFRe
NRplzfmZ7wZlVLu/6UwhDi5l4XgisjL2u9qgj1V35Rmz3eY9O7VJTG3QDtAyFal5
qKH5QBJOzUpddqwwyMWqiofJA5p5rHLZzlX/u/T+sAdEawFyU8bRrxTLvcL63lBO
82u9UXAJbyY3AWrk1lRpbjr6mt54wd7PEN/GbDG/SWU77gtaFOc53/hbnYn5MEYu
cFgmX4HhdLtKUg9TBCwka0KOAJGhW9cP/Ku8KSgfIbbPhD2NdGBFg5pE+bkj3cB0
mRcSmiazFZN5eeSC68dkWCf3si3SPxUzxxvRtXLQFPUdL3MRNUJUKgwuP2LYIHgc
hV46HQ7nxYEbVchqwP4AnjVtOxDUXmSCGNfEsEXVm16me8WyrGaLQ+UB8UgdJ7Ne
yU75sYgH8aV036EtgR/uyiOax3TVwdWQl929A6LpEud/H5+cYj2aNJMLFZnc1PaK
ooQ4bWzoTialTvxLxfVAQMN+5P8LIIyEhipbNmV+y0QsSrN1hyfNNvgRsHhoUzs3
/KJuYSakGMDYiipzDWd9kMYQ+t5lk/zZp2WLvX3nbOLxOUTBk3imsOndzaQyt5XO
FgLEbiOR8aARNu1OuMAb7WvxScFfFmXySBXJKzjSZCvuh0zHQK+i1e8rEkEph4GD
64AJNg/juIXGx4LpIG6n8JI/HrLDdoaB7M0G3eickXyoLQfQdiOYKYNKLwWPHabw
IjW+T3ic1Gzcx6DTBpj9RoWpE7q2xUVQwMgbpjTTGsJyR8EuSmBx/IqkJNqaWsZi
VtgUvySvZitL3cbqfVlX4j0popEKqo2hvn18Pk+WyKZ8gd6WH1vTCDcLgxUD5x9U
SzKm6qH4jSPdLLSCYUhGWlNXtCoHj+qGfM7iLvQVoVesoiXUTWujKP9tc9+Jjks+
5zdRYNxRl42hx1soS7H1UvDAkTDJifIynhhj/Kxtxk9HCLGSY08wefwPAnB/yOuz
pycts1qFdhU3ErG9h8oCrWarza3kEyWrJDweQPIoNmfX8xjOE0DQvVB5Jy1Ga7VT
Mb+YNwE2DYfdXt+MEFNvstMssflu8BnGp2Fb1csZLrqtce6Ut9Dg5dzo/gPQh41W
gpGav5zlvlIiGrimcYF7FUlVNMG7RdBFh/7yakEqCl1OiLXQK9RUF3NSigQG5vm0
t0KPDk5CX38uVu2aDUOGi2B0D+Wn84kcOb97lyew145Zf0cXp3MIf1pkyYxQsg25
et4XoXfBvLe2HEwE8LXwkG9wMNgMdyosuJsX6ooLhDERv3QnXHfgEm9Ytshh02RT
tFFv0zaON2DySMinRWg1UuF91ySSMJGGpSf+QrDDu6Mheb9QIEQE04nQGB98gtQ5
og/UmUqeQmNs+faRRXG9hdv5Ebptsmwgg1ETvcnAgkfAc5vPi6EbCsIHP7xpXL0M
zhaEvbxMi6aNQmSub7aeg1pyOEOk7OJln/NHiO7AxMptuUyK6j3a1Xv26MX1Qwz0
x4jGSJBC/dq3rbnTdXERN5LmC3qB6dNa2l0Vw1WHB+SzYo6skwaWdhj+oinkzLEz
JtFmEB47Mpxluv19N/c70UMNBd/AUo9B3b+8IhtLvjsjE/e5k3tWo0uQR/ajAeLb
5fXWtAfuNmm8LdMhbpodPjH50Mj1u9t0lkBXTunrzLYWeK6Tjm4hldrYRjPBXstL
tmOcEccGZAbwUYAJBMuNKjGJTlkWYoI6GfADaE4pT0OGAyYruELsR+kuiXRzj0of
uUrh654x54zcVGlCFalTcPe+ePJLZZLEtdiVXbCPPFbmP6PV1wVmB+FwT8KmXbAX
quN3WvyqdDskldXHy9cIkBHS3CBSRm2a3f4Hp29FlZSd3Y98xrusm3QO68UZsQPe
YP1VmJf/Egk8Llefq/qalDCEHyUXpjU6tsBxLUCqXeNf0tGRGi65DzybenmYZ+MM
GuQc8lXvGg39bQLb2IRb2WiF5SehY6vLapFGGZwae2kT+WBZ8s1z13OaGAHXo6BZ
onHubeWgV6ePHfT3XHPl3hGJedKn57RNL3PPg7/ZfaED4MogjLJVcbnVN6VPumUY
HrPST5GTIvzAGc215JLWw7ietduxSM5+yQBgOHopGAopyr6MpGg4layOkHTknPWe
OihcPFll3xJphjOb7cnDym/SCiPQTOurLWiZLiQsRjAS6TfwwTlP/fJVodIn21o1
IJ6FnNEY7Tp1H/D4YibiFy3QYVFiy0donNEig8m7t2dr5+eJ/9M6KihY5uJ6O3LT
41MfQf/iVs7MzgdD+5dm1LIjZWMmKTfNUCX9d+lgZns0NxW6AT9MbJX+gFAONWuM
5Y6Y6J7nE288FVTBDS5yVf+aj3iFLh3bufvqPBZwF1D0FaaXBBdeaCQbRcqUDdcj
iNcbmHzdmTVPHibxNkNPSusf8M6Cib1WhA9Fjr46jNSRW+f8ZMU/u1But8S2ezrW
5gndtXIzBQQ1VSriReof+GaiFGpKiQFtLzslOub+/rBnD4Dgis2zSB1w/UhXdVgY
fgbSjV40aklgZGS9QH9VJVvR3WnsZXkiuz5GmAy3+Fw2IJEVH8oiYmmjUKdZjxrY
Woil3mSsnZBX8TyrIlqh35wKFKS3xkT8nMVtcTEhxDLeahpxS+jfRDwysXeTgbH0
sihDGLBXVYMdTuU8A+3FZowHI/mciPdy4eM3AVjX19aY2lEYKfaBUIG2ik/917qL
2n1wH4zHf4l3yYxn1sBJ4MAvSZeldo+EFYNASWBxk8A5gjEv2rBWuhLpqT7Bt4JL
ntKRgcYNCcNAr0orxvIn5ETiHqyOzlD/ymjh+LQ1LUd92Fqqc946Tpg+FCe6NjGd
Bxf5qcIDZkzDe4/B8f6TMPtKLgYauGqmY/n3fXExxcgG39h3vt8gfnAnWNO1kLgt
a71XXSZcPoSOx7oukaVYvjqRfFbLPECGdA8jVNY+IpEgrQ7qj7ccgmGAb2YZ941h
KgbPpW4ZWVhWH0ihnetvgdO3Qx4q7Z46Vjtg+mq3W1MIvQhLtvWPgbq0FQreNXCh
LvlUKV612X3gjIzo9IeVfm2JW6xkdqxliHS4jk7oGB0bY5jFilWnXtqwKrHnPB/p
57n9TkP2JiWrHJR8oUfkVhsnsixVr8qsmCB+7cB9TZcfPPT2bmo1E/T8MoC3XQvQ
3aF0ZLzpBCVNu5+O98FVWi4Irm13Khc2tQNswj6m4+olek/bumqRRzOkp76NgOPF
Tw+ncNnLapKCZpR/HVaTeRMsxbnWrrG34xuYxYTqmRh+/ailHHappjDI/bd7v9+l
ADXdRUmMZGNClQjC4iVyMMDI4KvuIpkfMj2tdSTWdCuFH/7BXWCj6FGRImh++F4Z
thTNLShiof3Z3YCnLAcURisMq7sjipOcObm3f7WWwECO4HV6gsKjRIHpNeidburv
lwKgH/txTtj3x+RPFnSdFRbwAygB1XXyF4zd9KdZl873txT9VNFrbPqLhy8I+B6G
uJWofdyl9KP0FaQ1KVPXKkquXtPZQ3RzitNH1KNWg+7a4B4PJkudOmJUb3Jz4CmU
lzZtCxCznZU6+o1C4G8mCwx1lmqSJixSutaVX7uuu5zAthrXcu7qCKnlF2JE4hdt
7TmVBJFmxFATqLKrORg0r2UDrn+TMVOrGCD22/KOHaCo5xMwhdPr0t+PL8IgURKL
h7A4A2cpSyh2li7mctJ4q2JV5z0xwXTi+0teKMoZUBlC8EYx0d3FDt3qQtVcebSD
ibGofrM+KptjFjdGd2TS2/Fu3dU+rblZidm0whsyFzvi2Yr93hLcjXGCnyRKX9/9
jg4S4QehPf0DCIg+H9DrJ5l39vV8ToD20TmySRs/doobXh4meML59KYn+/ln/PaC
ZfAthPVPFu4Xz479axy/OVYQCUKNBV+QTYC+3ASCckdupCUPnK6lDSO4ieynKmOX
sOVE6wQ23BBLJNmOFKiNC4v7xZrUICjsa7FWfjkcFnsAUQzCmjxpZKt6alMWw/S6
JU400hfjF6D7pe1q6ptb276p0Ir+/OptSsfDTxTdqScbbknOqxNJPWuKkm9OHIQK
BFhGpxnU/jYqhgm23uT9umIWPzDjNU26rOlUkoa24GqugS30X8JxLD+FiHgqUsz4
zBRaIo3OMONHkp7oyzmu1lCdgdLaDQCx7KyJuOfAUCr/60SymBlSGmgTyTKfQPUN
J/C8bT4rM98ygUaYXxRMtEAgSrszVWz9OLyf4AIFmYGlhUdXmfP2GzbNnIcae5UC
Ur77PdFVnRMWfFWn+0HsWd+ufzavotZAyzbpy16xaQLAs+MmI5im+79Dmi9T97yR
YnUB6qWAJVlulFo0+65VU+qoruFOYktfSzpR9ZjXjwP4vqHMNbtavPoRH/09VLHE
/hcfIdMVCnzhpocHK0OVvmK1npjaEgwEniq4ZPkZyu0DT+laNpV8Z+UKBBZXvA9W
ghzrV5fESE76g3oWGchPzxPvRQc98ZNohUfKat3tzT41A2bQ8QpQ5ioyFR8atE/K
VYd6aZ2yWNeWJkyir/eRNDVVt11H3Kh431E+5v3PB7bWXZCDkx2RRI6XVGd6D1ZQ
wFA6emTjGLcOHzIZxnN8kS0UBnhwxQVJVMu9hnP9+wBI0HxYGrW/+In5pfavLl7I
VnWhn4sSQRBB89kFKbDd8sy+bgi5bB3XwD+caOYvMb4E0NJd2fWoO1cRUep7nB9K
4vtB28upbE973O5vU+qOSWAQdUBtah/HbTciKTp1LWoRqdYG4iTGKa2XoHFuF0oT
QHfcRssEJzK7NktgFWAw1gV4dG+16ljlOXbRWjqXoOlGnMjVLWmc1Y/bEILRDd8k
wq1vqjQOL+8Rf3suKGJcjIg5zf2cT77WDM8S7gjzSULlyBujbdm/yBRSFRPNZ0oM
opPn71pAJHjHccGPp4RCpqseOp6OsWW91NUJg0dODX3weJ+G56BpPr1JRABu/viE
dJyvV/192Y1XtX0WtXhmQ8cUHdLoC5IRldDkpEXE7QBzQCKvHs1edBB77ACOF/Er
RspONafPwq7dyPmhtArr5KkiJNZZo94cgmh3QpMqjkEyOp4HL5GYmE3xNL7kuxQ0
QLDZIbR/HQdEoq4GxuhRYPGFXF1QT7rC+442wknMSMtS1TkZTNDZnvr6p27IDoxb
9VuL2IVNyCyM+pVAg532CzxRxoSBYNYKKYKkB5uw8PU98aVgdKFCeGo+iJPBfDaf
DueASrSIKbymmy+jyI9HQEI+hnHxsgeSwFWzaUSyyG2XzYWPj0GN0GB0qLNAhgqR
jih9Knv/99XcZuvGLKRb9wgIq7Tt8OSExHER1SKlmcXDrIExK7UoztChPB0/jzDd
g+sTUrAVMnPFcdZ2ugSPWBWh4Dx06IlevRxW0oJW8euw/TW7TKyDFIzvHqRYqS3J
b/wBEckRW45hsyHCpui0QENXFsNh4lFdAKP4/O4UEbgC/kBL/xDqTwAv3cqTrfNS
ZPVIR0bd1XZNUD2YC92p22vwRSJOjWWlKQ4OPOOnt6uWgJ4PyWzIT4E4hhdN3zWR
VrNVGPv5gOEc4SKxuytiHHN62yXLjA/fB1WbcjkCRdPqAMo9GRe3ta8FReGMkJTf
4drH3xhClAzp8vdorPAqBxRUeU2QF+l7KR4fGyp0OWe5eSBSEtTzG7nWY8WxSEr8
qKgGSZjWlDdd0mVw4blF2yKiegBB6uvcyh4TQM6dPKLhLLTGeB/e8ZM08hloC7CJ
9vOr9p61e66JFGCvRrELzY3eBIWYqpIHrSqbAXfh1qIkqPBqiGcCNMS1T+Y1CBiI
m1Hd13fyq7MGXPJI0Eco+voMgDYbk5KnP8YEohRC3nwjTn222/7XGfA0Y00FeToz
+D/KAzrXa4M/4vJQXoMqfip0Ty27VsSpR2GcIyOLDo+aVOObSRXFqZfeFEkW2dYR
YXX+tydyykUjTgtI2MucVAhrHdt3D7GMlV2SGgjielUwZy36yM8iRbYKWX/QYOOY
SAgcB5tjcl/E166P8wkccQ1WO4stPSAU1ADgnJOu9wGWwk+jMNQG8tNkPRyGHxdh
vHeia8TyCt/shLiw5SYjRTJ09v02EXQddNQ24TRhVSfqigE31CHG5hgbZ26qqS5V
kTaCgMFVRRaEir3Bg7mDYJrKWTb38Syxqrqgxa5YFQ1DCQblYqsm5p66oqGx9g28
prPFyxRiMgFJ5IEeCogF0djU8Ho1HGqQXH8ToewpSJC9vN/VkZYFBSR12wymD6S+
4yF01RBPNN712ToVC1BRSoWlVKCJFVFlIyh11Z8WLklzkJWFYoILG438BPK14Uc2
Kd31c7b8FrYTN9XaGpBLXlaXYY1Gr4QxIF1WtwCIXi64bkmrg2zor3E5vHc1q3ZY
/w8s7nknhgjeTefCNWsewTMO2IbnnpzX2Dwt1VJErED/XLje/I+g2XAmBivc3AKm
xdfm40gdwl760VCRdvpmo21bNQhtN4jSs8lLn5R7tpFEqDXEMK1T7cXN9VWM0kKI
AggTpTjpv1qcVi8h1kcY+3eLBF2Z9K7xC6MJbxozY1Qf6uzdS1zL8atOaQtvIk+w
7DgPMoA47vP3BU16+o4uzuyw809d1hPeIhvUrtGYU21+KtVWFmRm/Ha0eEE0Xer5
7bBy+y55XG80rCdql7DQPHBygTMRqwz4oc4vHAPDUZMJDykgTAEsLRvtq5Y3vvEJ
asEpIPks0FqqhRq8Sk/y5FWl0HrH1gIxBNFrRp2hMYRFvHlq+6BlEaXoXZb2oR7V
NOE/r3aSddJIg7u8fe27b7lCWkcZNg+ysl7NGcOf91DowzpcKDOzBZd5r0/KsB7t
Rtd3yfizBctVkZDC1EYyUbAebnnkxhmVVO1fKZI+qrpVYamRE9fNuvEAy1qj1DWx
/PcbQrvpaWZzKubxJFHexqaory6GY2w5AOaxPMZshkLE+BV4fNJxF9VQK9G/Tr1n
EjVZ+qKKYet+t5UHTE5VkPKeRolwt/TDzHiw7WJIWgqJSR6ygp05HS0i6WM004Q/
mTEzjlIXNy36AiuIy8D2T0juII7VIVvafg66TcxXKpMJ1CXrcq+Psir9+eb/amHR
LSGXrhjHR2M/lwiq4mWi19gsHf8qFjqlaX6pfD3LdZRaXuD58EEKpVO7FFnBSTe3
GlFg7U1iR1ZjHetOg3owR3gGIIYh3OlaqCQkgUbfX5D7eNPSVz3FZX80oyjCh1Fz
fHOgpTw/GppR5Kj3n2i6d9wRKAUOfm4XhtBA1A0kk61NUHvgTFU5nL+B3R2IEKir
do8vx1kr0eREQ+PQ9WlBSU9U4eQL6CuiE6ZJmFlWUQZkYPC3o/eRT7LLflLXXVZJ
0EvoAtadCX5ZQ9HH+t5LbV1MmypwOC1gLFkgOJOBTBndnrasry45ifxysqmfc5wi
DX3GI1aioiJaMasvxENP+MJfC1rx3S7Fj1qH0SH+oc00gj6pHRsuPqjMpiDBnW1n
MXeaQeJCmXlT+1UTsNBVYHVaaAqWeVhcDpdXdPvLZsu19XP0t/IMJi5kAhnOxSuS
8XCK1fdWxqUOkScy6pfu+X6rk1W9LSfq1+ASFmL5tcOW4TWPK1PHz2b6VOs0v2IH
PH7FyY4SgjexycVjrPQsza5l7gHvSeiExTz0uEHgSoxi1vThKPtS8mIq078/XvMK
5jqbDvcYluK1+zOHjHEXTvr6xQa0b3T3IaFUfaH30F6wyYrDLBO1NCAVYHZiGWvi
Zp1L1789xuuj8APMXKaocY6u3CvbGhIhX9O11Ifr+nF7Cwlp+tCNQrtUwpJuKpZ3
5f7WUlcCxjpb86BipY5x0rpuQQgXD11zJkVb7DXwTabp2YCoe21Su5VSuCLXM/BY
GfSbbc+5yiXkgAJxieTCUjuRwcFcSKEvjDP1egv5YVCUbgQOftOpuJIovskPPKDD
JDxkTBg6AHw9D3BRPO7tMz35c4ZZXxa8TgvrVENmFcv4t1/fT5ME7fmgDf5ON+R5
H3CpmChv2+Wt45uYx0rAI9JuKpM+OK6oqo/cv/k9MUzx65bebviWLshJnWFHcWbI
3J6HGiOCe2BKUnPnS2ulA9MEWEj1okxW+72/YShU2f/4ADOlmy9jN3pnocjdWO/I
kBeTMtOH6Ts/mNuoaOQNkbggRYA7eeRQnCT3oeCf+DZL0eI3PnYh0fqGOKQJ+Gj/
7CE9obMKM10XKR2zVzJlsIJ3eOJulvKuCO1hLjHBnifwZ8sx35x8gA6ibPTV3bmn
v3dbPDjnmYC4WxOoJ8EmZ0tOWqkxcyjX01L7f2/uJ2PP8/wXScr8LWVXcYJ4hdiI
ApcQMRRkObsnRpZieCoRm/kygNGm+VLPQeBp6nBEBZCgSInh6J9mkMDARD7ySwgP
57xGvQXmpeHW2LbE2DnfBC3KsyEdvORiRR4uR9rzn/QBy20R7toi7RNgJEBUTjKJ
CylzGW32qNEFVMWU0HdC//Sc1L08y34I5JYvMcjie9HK7mhrLQbl9L+UbUV+ILzw
pCllxQph1SI1ZCvB0CSHpO8nmPCpUbx6mPzLNsiL0mW5d9Wsu3wF0SRVYx/cEEp4
ZkgLDwlZy0yG8+5tfTt5tIEwWfWMh8qc0RLeO1rwpJCT9cPmCag+9zfT7ubp5Grc
snb3IpX21bOtBE54R9NqTOoqFAcW8+odPslwgxVF7tZ7txiXtuRzYPYxaqvDtnYQ
gWEderxNeIA09HgpMSQvjJQCjvTBgu+DkajP9TkaOeQAYZWnn8boymzV2I5Uw8f1
DR6q/KLDup0ZRMJN2XXb8Q4kb5VOagW1jqs27m6UVho0KUF9pdKbJ8/4spnNt9Wz
Wz5sJTijk5z9GFOpDoCKDkmpgSCS2W+LzTOmM+XMj+hMegi9D7wyx5RL0Koyv2E/
I2btLtl5Eqva5spFv4HL01TRhXjjqBqB6KvabBbbIZG8CqzRkFiTozf/1gFXfyFF
KPwpxk0+mahf05ONJgD8Q/b3JRQVqxhv6LCA0ggaEFySCyA/o9u6su1tsxbuQzdC
NFD2CGGhmEBEn7hsWzyG5eUr1XTU2HYUrFL5IA8SFPhFiv3m7JdiuGEdrzHJh7sb
ZSJsdbQapgiOR4LJXgY+aLniPsaMKdAJcC3bvc0KJRXJap20zy+JKmUgNc38HuM0
iTJSbdtEjiPxVsl4V43ONcSH7UDTKdBY9dN4SbCctTvgJb4X3eJZop17p+piQQam
wMc4wg87nxumvGW1ibCas25GxnfJedS5Pe6kFjoVgeJ224z1yXa9gL7mwKtCdMea
UoiB3Rmvs4RLNxbU9bpogKGkkcRbS53ico8x9Ed8heOgCL+Db69js/o2yoq754j7
Y2Cvwz9gZKviTp/HO26DcOYUdEcZTU3vvdQq9LzAMdpAJbU7GFZgrSKvqcPjXtnG
YEi615YzAnxjnwfYZtWMI2+adACE6SQxZEbCjriraN3gmgKJFNvF66Pqq/MIEWB9
fVtb8MskHrU893USWF2Lk8fCOJu7+F4CetPTdauT3DcIwAv/rewfdcYsHuhHYx1r
SCDfo3D03sPbSH8HDvY3PoDkXjDjdT2N2rWqFhndECzoFiZtTaktGoL4l49U0B5g
58Ee6LptO0mmHGId72vs5Y8Xj6bFLlCGMmCaxuzLlaOOWkFaeK4ggaPR+mwHEx/Q
Stt7s47ldLVH2ehhet0wWLgXbed2my8cMnUNAC0Xc8lmM2DAET9ZHtzJmBov8mVH
nxNjmmTWNkANuAQ9/aRm2D/D0pKEQTwj6xMuoJbD7Uhrt28BF5sWuQki8fntTR0p
DvoqIMdGDSUmRgLVwLTRtmiWXlunKb6LgaLibwMCi39TIwkxTDxQ13yq9X8dT4i0
iMU6XEDhyJl85ZTBELEHFMGZRGsWRK9Hdx3Ii9M1w6Z56dqm7x1Xp7/9w5hp4uvy
WdZpURa3hlW5/hWw0/5Eq0AWmlfRWj0ebFgK/1CDWrueUVF3LuRW9A8BNr66CaOc
OZKLZN8Kc43iVTJ4CSTXDYqfYMj4mm7Yv8qGxweJ6YZKiQRftqd33sxT3Ofdea/t
i0WG+y1qYRu5H9KIyDTlXXBecPbVRDDCiqPEMd5xVEEmiQVNhB2dsadcX+cL6+3Q
gSMl51M+tkrd4eOyRqthLfpyaMvnK5coFTiFOEQ/C6jHtL9B6nw1GmUgK3cFQDru
36LP8lPfp7pxcsZdklE3vppWBntj74kIowCWX3fu+Cv7J0gIu9hTmcnLnfk6fF+X
aqTQCpJD8BgvWvD2LNnBFPtAQo92Vh4ev644FdJYTfq2w1mYKBFbqC/ZYaGqlG2a
5PlHCmg9hkiyAlc90VBSc/0zZ+w62//d2dadLVIKeKezPR/tS7bkRISFTdbFSE9M
aHH1iESPwc745HcYb0lcwTq8chsSdbqyh24slMcJtUVvWJefJyHO/llu/UJ4pJaJ
hrYCh+7CP84ibYXLicg/t8UI9JS9X+p0melSTXVZl8W6Ow2WlnJFJsjYAKeUJlSq
Q1MMnWx95MOUCYGPBCV2B9RwE1vmnqoe3WmaX+RqutGAOVnm3DujO/gSUo3kVUp/
AUFG0n0ygua22UEmu81SKcfHufcPOMS58wap2+1kIJCanv9U8ckmOzb1llnFFK2Q
Kae3/9144aTfjvDTkTV7bQ7LPC75IE+62pGDO3LZd4U1YMXCA0OztqpQ5fN+poOf
m4WBrFrdNNVDbZ3yCmXQIAs8wiyBadZXX5lieAV/Vd6k6/4ixdqsSv46kkoknAMF
vfejBnVGuoahSbzM2XKcVjFArx6yZm7DLNOIWmgm+3p7AUwDzBJUL6f8RD92sWUn
lbHt5l5rXTDhm0BeAZKQ9HhDjmamqQKTo4d+58JuCBLfY2zQKWdZeQ3nAmYvS/4D
8arMt8BWNoZEHq50QwzgVzTEMq0ycOFshgIGmSsGVEq3YbPgXYflpglNyKbFEt+5
ttcEu4/FZorMcToRQbSJRjwAu6U1MY70sq0vKSy29h/HhXboWbQFmV8tigHXxG4t
YVoyIpJyLGJEfI+aQQTimL95MRYjoW+waYvs8ArbVCa1B1ZM6VQkmKYpo1EI+2Vv
jd5+mLyHftaCDL0cgn19BEYYT+O/BYSBr5Wzq5uLVM/0bxrRhloCtRNn2uny+NB4
KNSH745vQYZkwNhS5O8zrJD0+d1lWQ/1CevpnUm3TxROIBaJf7Ttt9mZCxawxEBE
QwuBMhc3UGmyXUDcwlC3ZjzMr2+dSt4qw9w6Elgq7mNhLG196BBE1QPGk1S7PXmU
Ewo/Zlm+bLCCMi+YvLRGyu5p/i8zqnnBiwqH+slXB0zCzvZOXWvyvXSDQ53C+rgW
GLFdyRC8d0XGAn/vFnrK+J2aw4WlwLvDuHboX4xZ6R0+OGqL9Vi90iHnetQZOJEP
12YU5FqzjaSybF82l90s8eHoNGSmq0eyMd8Rgk/jlphLa07UIeckkvHJ65L3MmWu
jAUe+m2SHX2Y7dhUHp5sSrog82fYb8uFSW5ydBkjEKHMNE3LkmBtD7w2fNcKCuF/
1iCmwWydhmAXf4XNkjwxSQ/DiRRBGSZg+cyxgnLWElEk8EeFxP4WMXyScq1xHTks
DEDhsBCz31HmYeU8Dc/ErmY0Zpitf5iWcttbxHrHwzG8lTZXsrKUDnJ/cwQm80dN
No9pz/2ryN9LhYXbjBrbNGwsuoBayet1cpzzAgUU7/p87LEfnds6caTELHSIbkgy
1e0+KmFWfCjnIApVsy3QH8/B4wWoIIoe+dHnzDSjU2i8yU1hopW+szJom5j6aw3u
vRmGDfhWvA8vn0WYdtFkmxjiEd+md3HdZr6BtPASb4MKMU3a7GT/JL1TLFRruO84
cKsV80B7C27hRKcD9K8/RK7tESF/VVr6LAukBz7EOYyAiXipHl0LcZAaV0Nm6Bub
bN8Cnx8ToUB2UsaITOY26OoXT0BQ3oQPVCafptN+n0DSjoOsR9CuAtrfqUrwQXDj
xh8Fnd0cFReSomAtrmCH7Fqqy1WDpzs4J2+a+qC0mmppsY1AJc4B7aKxtx1EyEbN
hbtfLfjTE6I59OCcSZzV1xNFJIGyarp2w3GcjOqBnq5QvRXsjBLM3jgA5zjMb14U
+r+jSlOdmxozzc6PEp02ajDAn3CJhQZxSwNVSFnejZWSu+LeIjWPqnvJuPTLga/t
O1Ddtc23Tah7xGLSajBtUMWYZvRppZsioZSJS5v+Qp3ouolRHJz7eosaI+SD5Tjv
E4Vjm+itdBczd6g8zRUsX/szwPGGIjbySBmlwanMFZT6k4A12kk37da8jQljeTZ3
trKnjDFyIbHUuzkAolUqywWgMjaY1N/9l8I7Uoz05NWC1E5fF8z8tCICJryWOjIR
cf6tTLjYF17GY3zRUZV3CsW/K03D49Sp/bfwzbr8uBqkDNY2naW3xT9tVbTK74zD
O2fJOic79h98WSVIAwIAEP+dIUTKsp9vYKsS4DEICA1Q6Csc+YNTordLLJwuGGuO
dxpYKdc2NoUEVUs0veJfM3K9zxNK1BvNpHMV2yT76SVjDzCWZHQRLb199+EaoNPd
jLxJLTSNCoR3F0eG1MCIN4BDCu6/woocGgXFLaoNSdALHmWIN0udiKK6bLba5fry
to3913lI+JqgpO29jjO4CI/UlLVcVg2ifbvvVwFBLLH5alSlanHw3uAdN5zuLqNt
4IyCzH/+Au/Hgdjwp1E7rweEalxwrYImdK0Qh0YewtQAXM7D8UYtcufiN+VjFWg6
jXFd2M5rFvS6rHww1jxLSy5TZTi68Rk6T2cgDaESROAPG4kUy/ddo36LFs06nsU6
W5dzBgKVEPMbwNMZAZhy4Ivw4Dzldg5xk8AujFc22WOcAY0ugtedoar8n62m0jqi
ufKvLKNfxIjnSoL25ugZ6wdsBF0Ol6+Ida2wE3QjrT/qBGWW4zuEmIktbyp1ltzE
4EGyjB0+8PC/nAA3Ts0ZiQPRIQtgnVI52s/IEd3dO5PCcOixw36bP1U5lzOSgmNC
7D6OH9axUMqmmI1S8yCohUU9yA5XwaiK1PRRudk5GumSjzFv9Ecc863Xp31ryhwP
SZactdbnxacznkMGKVqSSnza6+nRa5h2tV/A3hz3DGTl4ozWyhq/2M1lGelDNjfe
uoVYuatXkqXIepDKmGCT5aUjOtUAbaPJ9cbJQHAMvl9/GY23KbpyMpVWCNwDu/nc
Nn2AhwFkixc1IdYqKKuQc/KlND2b9jy51eAX1WYjC9p3kJt0ZKWw5xoHvX/fhfgr
gkd7K2ulYxLr03wzCB/3Oj93rBl4aFPNtNcmQYHRK+iwi4RSvHN0kx76JvxOjLG4
Qqq7TUN5WdGIXILCbg4ShFgkxnYgjwH16H2ofHeoJuThk2xJRFfU00SYXeZLjE8M
YqeXDeIVW8HveeBigIXWrDtYV7ozHTrU7UArCulIM3x5Kj2K8HokEas/I9HTfDpw
KH2rDzu8nCNum4fXxpmN0xadw4QAgPkj6pVr8Bh9vJA1A2k7QEfZFWThz+Z5uuXr
fRs+SJiKT/+c7GdcCIcdQTSAxyfQHpmbI1wyAKpggd8tcf9ST6TfWMi9hpDL+nlV
WrJBuxoOesywoOYL043uwl5sHJH1JaDNr13s8PfwgGCUUqPnsKwpEaIi26/4dQo4
QiqNkkTZmGY0KkPbPVOUMCiua1znM2FPuACSDLoX9DgFx/AGmIEyx9G+auOlZvtG
+/GMXiOERyeIbKUDfeiJ9nMeKVf+Fx3mQMhR3yTpsWPAARhS9/x94ccK0BSxpk6E
1QpTQ/ii45VtDHJd4Teu4/H08ZQPUm5xjcGICw+jMV+dxfui9crUAfIIJxXC3ui/
7Wo2DicooYcqXhWA6rsL67V5BDmW8LeM4CSmgL6vmf01Lk47JR+ReqiejU/PXaV9
29lsIOHiq2qait+RSHrGMBR/xERhoGdp6GQyhAXzJ+u4ZCluDi7cNuXQU2j6SWcf
L8XhiRJK9LJUEi+9K6jjXTmk7V3ziRcGo7Hqx0vHDOrqDhQGhiY+JGMcL60EnGAi
Xej3+5DP3qmbQgCNWeXh5mLsn6nsX4KIN98pzn9JvUb1unMkcUcmF4jErx7uKwDs
QVzRlxzDYhJLIAK6KziBS4tMb0RQ+snnNbmMPYuTHcu0EgOGLpTKM6eMMWzkf06U
cKwdwQ2kMYgs3Q8PXWpYQEDfw5kjjZsJL//0xnm2YlnDZ1g3M57aTK3Ttr4TGmxR
e+VPNitfwB/SkLLXe6i4p6BTFvpzVM0FdiB8yS4AIk+LlmmZ2VMu+5VuVa76AwW5
jiVAb05sCMKfJyyn/ehe6sQ2cXKUSsNyKucsviarwhvd75vzK3GFmoEu5PMKt2iA
uf5bCCo1sjA5JAyrJZe2zgn+Ty7SZ9JFYUTYsQxJqwEThtKRweTXBhEaUUIPPqWQ
HquhQAqbsChauLYIMs3iakqrtRa2u1b4YIu0nb6eJoJoQ6jpBadefxjwd0EOQCIQ
ba20oRkzFqoVZHt8d7zoJB5IWFt7gpEx4DEUwjWhRul07dreE+yvPF7gYb56lPDX
bpGJMLUTz7b8E3m+OnYXlxdJOhWwm8zggxluV8iN4d0A2jIC+o/EnlHrDWwOI4v6
7ts3ihiQmbp2BootCJ9GhR2VB5Kw3xcpgz9WHiwwewXTWPom5AsO+p2sZ5Cavv98
aiyuaNuMZ3OuMbgHkbPs5HGPVlFZVjQSHnnPh18LIw40six4zX1kIBTYy+4W3972
Mir6nxTXBF+XNR1IlPsz0Up6WhDQpF67iWxiA/Mu6F00Cl2KWPqoIpxKzIxQic7z
0yVNzNh+r+/fchAIkoy9u4dXrmkUMO2JNuQQa9B9q3joyctxauKhpoJKz7/uDnlX
n525w2Tj5iAJXHIQIuXE7h87qYMBk4ez2dzJKfv4uREMK5BHwde/ySmfOLQPq9DQ
woWqwbzcdgvaCL+Ta2n0FlOxkQ8jT8sNXZd1ojPGyRiQwZ2rHWTj1ID4beRsoORn
jEiboBTd+Vsj5kMAtIBiMVUgUMRDWva+r6pWmrUvWuniwcFRfDbLT3e+pTyANXgA
5Xh8Iv4Mf1GyGC2eLJ6l9+49/C2aoqp119+tHkn6tuQWls2lSRAxi6mxMBvO5zeY
xWlyViVDGstzP5WpjqX1pSYKvA74BxMAB4suTP6NVdrXfL008UnJW3yfYbuIMC88
6XMoIFBccBmFzMX1L8tgP8CcgOjf7Dj35kjfdxcaOa2a/Fdu3vP8BxDY6tuM2fj3
mqWC6WVk65C6RnanRC6XuEEs2L1RFZsxn+Qay5u+k9gaP1UAjIlokDldEcElDOzU
1eIyV+W9z87lyqgskIVqwORM0o6LllM+LMx6OdJcsUYEn+PXwLXGVEkLojPJqRWk
J1EJkAoDgiUmzRZnBXwJN+ItIwI8wCvs1uUFqLek5SlmhZQ9K8N69HxoPN4BhOF9
Rn1fObzGUn8rIdQlb9gRRbA3GNcyYvhzCNUvj1B5J7QnVgSo1k5TPv4flyA4cQxs
Te1GVJ3te1XYoPvRcVtoUFhRxLpMrylcAfdjf5vaCawLa4TZ3ImQdq/g/Jl0Jn7k
yuvHgFl5HPxiX7kzF55yiom8nYm1exzQ9/s1M0OggFF1py2+9jS91SZ+Kjpl5Afo
vemhmmPXUZBzFLkjMg4gCOSc7IRt0jh87rnA+HA1S5B4CSYK7y539/NfOd81e+pz
eR7a9Kf8aqryESfKF/1HyPyTwgDP4KVIoCjKcRBz7B0Jvcnq8f6FtE31z8DaQodE
zTKqRKU7ae0X7dsxovzBIU7V/NwiPXy96q/i7daEivTFEdOVrCud90bYy/UxMd2t
VmJ+Ej0V9MqIYvjrsv48SZ/DOntWfkd+LSAJ0a4wW2syWvdcDVqEg0nizI45hjiV
ErInVEtoh+gg36J23uzax/DubZr5ZcRv32uVbF09I6APyxUzeTCjA4MUh5IRG85s
LMd8+ImJe7kD8yE7vhOfbJQkWB5kTh4n+7KmfIkFMmsFYKniDNbpQTkJTJHEjnYr
2+a0BMjW86/QcKasAZuHG3CBwl2yOqzRHJHbPz8db4/xS/QOxSGlUtwUdUtCS3Gg
e4/lcrOtMg/i8DTVRAHB7+PjWaUL7CE3ylbeXEeASoL5dJoFlBV7tpOFhEIOWH8z
yZvcEIPb+dXHpJ4yqby2s4JVz8xAe7EiIdVo842cdBtNeiZ/n5FEopoHIjUV0gRq
jp5WHxvSMkXAX1TZrhLW1EEBqjT/3p16KNvPFfjAeYS3DwjQ3CH18EYYC01DDVUh
/Fb5URQbFYfB6WqxRWJvSYHmfmQ74hNssQOW7iJ+D69ryA1JerPYXhcjpGlYg7xO
ZPN9/gTbz0H8ToMulIZFAbCIJfh3+EvTYF2PAR5xODsiYqnn9Cg52dQAXUajTqeK
0BUbJbip7CuPoAocadJ8BrnBUlwSv1B2+XCI+kJQkYywEyzJzXihugJiDfy2zFcu
3VCjbjaTa7JeknfVEq+2GWbx9Q1Xn/QmdmaEQRa8VudsLvQ2OSvpm/nFabc/jdHq
FpQlguICuDDp24qyMlPD9qfRiyA+gPIjDuckvbDTZV2xia9BOINMsCyBIYEMhJ6L
/jRmWYjNkA+jU/R3pqmm7R6Qx5dp9SsI3scalz6Zv3Lbt0j1BI6c9N32ppkAcC3C
RTGeShEu+0e9ijGBcXwev4+NeEghfsrSubEzMsNUEhlhzbpBFqbdkECm25MvPEpg
i9oz8SvTXkAdY/8T7IhPVC2nrZZbHiW3hRPrfLgP4H0ku900EIJnGL5txDXGEztF
/qAK5pcsUwMOqgfGXIZ4o6Onu/u+nMhj+ZjlmVZ43/vwkm633g151AMaGPTOb6MQ
wXZ39wE/I4TymS0KGO/a8f4y9K8EU2C7+QGpUzp0cZrBwIx6J2RkqtpA9EYZJzFs
7qGSWhXiPNfKER2FyXxaD5S98qJT8c6qxOlab+0FlgRoUvF4iHMXYN9GQ8tQpTLw
enVFNB6HwG4QlK4vyAppSySXOR+2TkWvSjOlFD8E4XsuznOR283n19L60v00uByE
9g3Ej6580fJMYNdbian2CWS/tWY3Ke6poO7kSTDfNvyclc4T3Eyw+JPrXHuTU93l
t8SHHyV+ecuSlQHkJ/Z0SdhcLggYOpA6+ToyfVbbal+68md8dOZjcl/EX3+WUCDM
JE6z2rGrIGkMpyfUa+yEe53fEtECQwEM8RBIcLuG4xwEfxDzIA5b1jhOmlhg60KR
vkcmJrzMojYfcrFVlhGT2g6Ct043KXOAfb2rFjmpfQszhwZ3pGoqqmiD0RseehBO
oLZEfb3r0KnnE/BlWY4ZQ1iaCEEHLHPjWEiqHpDNWf6pwUrumo5ZYi9b6dqCJ4T9
aXY5kPihYNtebTqMwmIWLArtgxHZ0mo9V/vI/4IiuceAt00oKunNRoIK2/yf2iCZ
f1L7NeBMFypuNgJxa3OophuNBzMIKeeJ7gPlN7DzssD6Ax9mPOcu5SNQIGKCaKOt
5fGVs/3rDbx6jOqXV2tPL9AO1jqX4lUVWjonYg9QrtC/Y1iGXGwDIPgMR87tQhwq
o+eFxIQBcASctG148xtOHuq10lvIEV9IekQ378eKslbyemD4jhPUpYqhhNzLJrZi
1zQf2otbl6RKyH7xpuppt4YB1ewgZ7neRXVkHeHiYgXW4tTH0C6G/tK9F1kPBCsa
vLDnRDYx9OxOGvyDvy6LGgoFX+EDshiNNIU+eBp8MpTUQXWQRE4FsFSO/NcvAaeu
1de3fAfRikdhh43xR5pI4kApQhr4+tup5JWSSJ4bV3qoGiZrCfTeZTM1niKLLpao
wfVU2/kpk/HbW/ge55HdsvOmupPeWwxTd977OqzIrx/RCS53/vx3F9wXeh5YZ5WT
4yA01u4qBGkyhxLrTe9B9vQtUbQ/oh5vBRI1gvc45aC+mVAAJbsUBgK2QVOrAGaT
xBe3W1ZGFgEh6n9oKaZAEfc4Y/94ePAn/Z7lB1zVOms8kYBbJfgj0On04ev2zN/4
npwNWRrj+ICXf4U1pz1Mds0Xnfd9Gr358bC2QaXxSrDw34IpDPt2UFXA5YPVMeAB
J1SVAzMWcGDMNse8AS2SGW8qey22BingkxC6oxjAfaJ+k5d4lFXNO1jALfD+V/um
GOYcavOP22WULrdc40HWXzd/qeREX60juISG9VBFGkFTMHVEJRudnaAH1owQdmJX
9vw3+SIKjd5DDeGJieQ+f3UeH4ikNG1VPTqWGf1Wgq7PHUBOOLG+nLBya1iRMypN
iKSKE3T2tHYu1RtEipKgGbZ7O0Nmnc+mVAejRkv/fC5Y87a29Xm6nDVlwbV2NkAV
LRFs+Bu4AQVKf6CS3ceexmuOVqZSeoaW4cgDOJ28jEHX7dCpXNremmOZHzYHFie6
/0ikBfncHobeJ/TyydIHER2jpNiOWQHIPZZcjCTknVgz5+I72s35/3xxcbRULMYE
tAkElechQCnEKISqOlVdoKRno2VzB9iD4bX8zgO1PGm9Bvaw9WxSMkrOkRG7+wGw
P3CxPFpkExQLjKUdaCsxpSpLYYX5P5bvOhoLRW6alqo6GjwFAMIyDmTH6Xj6Hxro
kk8B8s/swcte8Jq5hQfmMuYpwuhocESU0A4kTw5QRcS9GnvJnFPbBOdk0io7CLqU
5Hyj2RV3vR0VvLVu+MbrmkPVdvEFjyhqfmxRiITqjJN8g7mTl3FvKXhgLZEyV7ia
WBj98vvgG6iab1jD18WsYOq3PDI7g4gCW0xnM6nU4QAbggKRnPDmOspVkFciEn7H
WkRVqoTFMVtNPFNkh41IWTzAr8PsM/v4+6pKNRhIQlRSDrqNfb/Q/LUtX0m4tv9l
DDljY7BawNllm9wg5ncv3UEzOdhQZzUBg4jVBr33z/q4TTS3bngJw3iWlB6K89cG
CTQekNSlFy65Xs5owIuePIvhGrJ8xCwyWGFhoAEuijNYYE9ALpCJXCP2pKwqKOY6
7sTjuDxYrsmu3UhBlJZS8MOYRrm22kHhboj60FUmtZY1fRRqJwWZmqDvSr1B92GB
1SV5rlAJNIpN3qqv0COX/gXfDakpaaShCwbPj/CTqpmetr4CAm3unulPnjSuvgfu
99XQVqHgwrA2w8ZeMbk7+joTZKzqWmZQh7dGBQ+fRlcJXTKe/VDDbFmsxRyiK3C5
wv/jl7tjMdGeriDX0mYN5zagf7QLRG9VIO95n21JUN61KUfQNjO+CBps5G43v5cG
7fCYv6kSYLv8c2HvCY7XVHBYTObnrEbtqThf+N6ukggHneCOpaVt8UcsXZFvhvTq
cb0G2/MW3sFudd0G5LrZxocN5+wH8DYewOc/BRpNU8yTrBK4mEJBTl7FG+gwzIL5
BjDRS8DDRj8P9TkjRCy7j+t0sdYUQb5EfcohogcFcI8+qD5lF9xpCxV1AiAdu2cz
sAyt/s4JP/8gtEAysMnmfbGZubZ6X2Cz02JNCcqxv7VAGX+g5oP4sJKSmxOI3ESm
LL1mFJOVfVMGjhs47F7K272a/ZaHMp5zFayVDQLdCWh1ojI1eXpWoL2ACVai8uuO
iCXc4oZk0Yn8WiKyfsmOjebH7cxfl0hyoPZMLO3GU/yMSNWScpMa25R67ITvmzN+
MoUPfhMyDgo0KNi+VGqDqPpaGLMFmLL8bCX6UPT5BPQ8xbToAfBVqZS9G1sT3nty
ZohupH3ydy6Sae/GRqVzCNN4/hJcCXAkqPbWf00Ewvh/Sw1izrtHMoQYH6o/HUHb
ZW/EwzFEnoA5I741SHUdGiZH3jFPaQm36nFTsQvq2+EpM4E+aBR8+BMJZUrjJcD3
jMZxXlotLs1jD/RVhahKJwKRcIX+DM+YXjSudZro7/TQorP6/qIuZLiTDBpc/PEV
GuyucH7z/V/zeVyMWe8lSyatVHHl1Eh/UdKRCawxP9okO3oWQPOrfEGa3DpAKtYY
IoP3wf01YoPq2ZHxWa708DQoVz30MJLkRTKp3dVD2Mq8gyPXhUVzMIQLO22odKwy
suV60aShFds7Nw8xvP3P5NXhLrVbqlZjJZ5CUOx6bkIngbNv0X2EWJEk4ncE4apv
h7QXpUjxoBQ40wwj8rLCCTDh+KGaQMSLNihnpcVBHCo6OJiaAJf9QPsoEfQ6oKh4
zXFjzniYXhkY/Iu+2f2vPMeXA0cgw/4npzFMt09InwjvzFfOjoItF5BaHkEhVUo4
GKtGzZ/KHF/Zgki8bZbJFagkUPNhDOrZCepDoNVeyv2ztmHgU57hxBFHPEu0Dz+9
RGcVHG66lCyt9gz5vm4GQ7m0dW6vgam4WerS7FJcAxXXO3ex89DGjU3Ucle0fjVv
hNp32AG6Z4PnXyVih6r1Vot/r6Yqdn7j8VkXeBYWsJRrXe5si+xHxpQy/f/KSZu1
KXM+O+WNlZ2uLeA+55mb8F8jBJ5UCS323EUqkdP/Axefr6q+fTZlD999FQKnmRIb
LJYVZhdfO+0rIEM7GimSW2LRnLg4vzV8sxC1YOYVAWXbJwqIeozetXqfrOgIjMq9
KzsS65AcLL6f7JwvsdQD3JcNBguB8aYPe8RLxRjaKN2h5q+gqXgD7uGg9+JisALp
SYel9N89oyOAf84+kfftnWI2adv0mESAgmmViD2NozWq57mI4+UWeExv9BmLIHmX
RqKCsALmGQFENia2JSmc7l5QEAWPZ+2a8/Ur+49dzUVdR1GTvtfo3wTPJAp8x0+F
JagC+HvYK0X+QuAXzZ2WBPFfGsiaHqRA4Z+pqVJ8HLIOn+VKjrmb3H/AE1QfACjY
g8nDts2POgbTg1/iy3pWu4Qb+gphiuz/CL0qznULJDVzJOV7UiF6jIr3Ec1uL0GR
XLWyVIu6QCMlO3sHIPQBm9ToT8at4oUj7wkpvlNGfIt6/1bGIzCOU0GUJyZdxrAp
GzHGs1qSk+CR0OC+8M+kMHVXp4lJXgzSYmD4exknDuoZC+4rCg7jmXu2ssegq430
2IiHdoSKs+iPHUgmi5X+UgtFk0+70HOd9JdHSpqLmTUrplPRJI3tFAxzAH0uVL1m
ckBmp0dHEb2LtRPo8SLx18VYz+qxP+/by3n4/AV0PSAQheysU3RFJD/2FtQ5hfWk
FigbNZh09kFlpuwps5hBqrs2GD449TJ2XiEHQj8DDS6iDr+VpMUCbjuxC/NULgtq
cH5WyJWQHf2Ay/MSPBfHiSOC7q0AjJyBC+ugnJ4KNgptHngG6YUBqcgqDA43KMDs
YVJr4ziX4R+PsH/xT2t9JyeHi8EekQkfkfIN/s+hYD2ex1q5Hvdo5p30PscQkPM+
cof8p+y9ViwJ/EjhKCTaY7rYLt4jk7t6w+odxEkqWTSONhrveZRU0bT2rYat3jas
c8aECHslszms/q6LbOvrdcKVlu5Z2b3rioUMuMfXzCL0ogmHbBVgIPQ3D0QPSRjL
B+kK+xUGAoJw9mE6jIEuRj7RCPUeZA7/jXwcLm78wQM32+eBB48Lm5Meq8YmEu4/
mRWi15N9V0a7wQojEnl65hQrS6V57ni0Dl04HSd4pk3VOstecs4AtnFH8FmCG4Qj
C+ja42fdLKyLy+I4aP2JYNBMziES4fwKpvWwxMz7zYhLNTZCuSdr/eqYwCVoHIfv
7g5ZfDbfuBarOzvSCJ4qomPTaa3dhMCfKDEwn0W1eCg5tUamI2MYVQkJmd0U0FoG
NPCGzXGtpXybQKrj1w/HzdSSxpOmBccA4vakqS2Ip2PhrXoutX7t4eiweImX9VMN
aOWM49q5K8l5sodY/HIlWLZT7BdaxjKgKqikm4cZGLVFokGBp8yufNepAlPStjwW
sml5mIxpLwGcnoBqHnBVp3c9xfXm7w6hX7z319ymm2n6oAw8YSDnK23mKNuXid/G
4Sp+MD906+8gNnMkxquyPAqZ2SzjeCrkk5w7B49bgwJIMYzP63MZerw41SpTPlmj
ekzvKqByem9s+oOpzGiDXOPz/vvXmAAh9SIo3j/GprC2TPR2S+vn+b+G8hzoxLwo
YKxyHcz7rEfvdu8OBwzusePstCN4VwDnZIgTghlZ8a0bz3jtfGialOGwve4fWjox
CDinr7XbLw6Wd+6XfxiPm/0kBVPtTNlA0gLVsC+CV15Hm4od4W+Vq5/n6u7bNGto
sdVepkSaYO0lGGATG/dJX1mYeKpHHT5GUeUWz3fUb8svJhCrK3sF04QhXMa9eJ7A
zagQHJL9TD9scjLvJc3Ngf7yCpPBF9MG3mBaihcJ8e3BX0yea+REg8FllhkP1Paz
fOzxu+I9zVcY61HU6ElfzaFXpw639EkDl+2xNISAXXGmV8yFo5KC0QPOL45v7/U/
46kfVvFQRRDzw0XynRen+SBRE15cpEgd4imDC2bMfcxqalXq7hD1G8aOZ1zWnJR1
vbEfHlusBwMD54Y8NI/jJ6SF5Me05j/4BOE5ffkV/2Y4QHgWET+bvHD4Jsv9RVn3
l/NmUFRebeZ/ssB6bAopAYg5y3J5S4hXDLTUxGnehKDqDWZoNzgypJ8sMBEGLQKV
EFa+FKtHu2Gqg0JRuwyCbuEhvnRqvO0LOOVt3vKwcuk7x7V3AaBYVNnlyhSYhXWC
Zq1mpzQerHRYpzHk7kXT1/y4zEeCTjr+P+pnwm91q0k0dV0rCFqIKpRoHsLwxP61
w2GIX0XJaovEpxCCOIct42YbSqzWSH7LmJZBag22NQ9UtdFFq/KJS2nTNRLwKvvT
Fhbtq3J3jANsDWhbANQdpXZG9MTGU1xwL25U/ACECFiLr0aUYQudMOls2CodHNVC
YXZfMHvrYZoDpyhJfYO8XX4vnS3pJRHDv1wBbkeJ5u3KaFLizy6/lPF9Fg9weoTv
DXiHH24ZtW8RnOBNaFUsEPEyNyxtJkghUTBpsQlQBz4X1Ulil3fQYI42N9K7wTrp
BW/XIDt8GrsUf6mQsmsb28KeU8DTnjDadopHCOtf25ZHQQNf1uth3ad++u3Xb1Wm
nbzPRrrBft2WAtNEFhXOCAnRy/46Yb3Fm5Sp8wm6qgVReTh+fq3vNQiWh9+zI0GR
sMWOnDBa4xsOAj0ZbcAE/qBIH9UTxZg32GmqdPee0nEm2zEuE7lfxNoJP0xyhGfJ
Kn+CdepdY/etVe9TM3R+hME2a5PY4OPqS4Vlr5SyE69mE8Rs+V3S1KhYBpnPAZye
4DfpTV53+tHdIY6P3hICDjlmqelkYi97EMIuOUW6GX6KA6UzKJTLW3TLVbaOHqid
bEMNa4wflZ+lCWid0OrzB0GS8yRa9vqi6eplzUa2hUdYZVmWq2yEb8GP0VzMKYzs
pPnKGWrASCX8px8uA/FaAKN0XTvhZJms3s7J/BhrSiwiFSeanv7loUvlKQ2lBgpl
bHKk3MJRqogSxN1N+O9TPkXyFBclIW/HKK7pz7W+OkDkOfLupvsvfv5fcExKxQW+
zkW53B544mTxMIMaCHBrIA73UbcU/ZGfjHAi++MEhkvgRzRsXM6Qo1CioQCGw7wA
YS2J8Nv8DIiUlRhv4LrYzLFgu4pdFKDjshocv3a19PHQLjdwSS0MQw1KvdS7yj0r
Qcp3kAW5WMCd/NWjhRj5XBxEYMyqFM03+5yQj3hfwxjuhz+IDCh3NcX4nVKdlCqb
u5f/IIkHaLC3s/RyCWTEyCx1i1Lbx8EVvCfZChemlOoiEjm9uguyaj5DPorMzv9G
tihghclp6QuWtUcQ93cxRMcBTY+W0NGiuUV5SVlL5IOAd7ISW3PctSaLibuC+8Mq
QVandP3AkrK2iNSe4Xr0dkS7mzBg8+oMFQ2fmbl7bVSWOwcS40OI13NXx6vbVcBM
mK8jMqw5Hz+ObtepwKz3jaQm44EzkIv7A2KwATzznaRx7U09zYFueqp2CgZEq5Si
oSo3sL3d6/wC9eHu1KHllMI8Zh78v0W+jA1c3poIIn37+t9U9BedcVGIqrmWPWnW
+bsLMMsi3H/XYNM7+ZLRZVFzsIu9s33BT+2XHYRtRCH/BiDBQLgbcqDsdIw6CLE2
PZTdDnpvfFnPCOGyQdSYR8VY03B7qeXRlNZQPxJsPsfizccsNAe4fDRTsBEocyNy
SPhuXDlCkhe34ejgiy70PX1N4FgvdCi/uoJldUz9xhwIsPY2b95xzhZ7G25wctjz
1Lkgh56EaoBm/TP4O/dE0Sf+DuFR63BOb/stuS3sBRLC0gvi0W8XoSBcP5/6zA4m
bPvNJZEMgGjLMuLAg06DQwdoqe5C17MW9Bdd0PexA4o7EsETV7dxgjnXujs0telK
ccBWPjyVuD/eLwEDiSpBRT0WHC05R3kKRzVL7zgwgAU1ttSXy4Ou67RiafQ3GVHF
YoLffnC4r8heLyIYbU8cJg5UsSiYh8iZaAhhSce/SlG73AxWA96v1S6IYzZUq0gm
gYaJmjfN4wEhzenGFl5DNtGS7vBEIiZaIemZQnGjO7zmAqB/Fss6N6Hu0Lb+Ht5z
UmkEFHZ2wSOIB5Hgvw8YhmwrVwqVlBuSM1L3aXr/D8piM/+mTgduhVvLUu4T4Z5G
CV6Z0Z+g55GS9yBZJYMGm6XVUBCRtU9OnpLydu/jVPw/yRmj8tffTgI7an3WlBGw
0U1AhJNZnp4qGmN1JeN8zWajm1xWNoASHJ9A7zrfvoJFMR9bNiyicP+ujXBdhPuV
kvhxGtEZ/plBA2yGhP0aE3ofjJWjS4Kf1hKUBIGWizhy0/4oD6mUIDUB8/pqzfNM
DsDiQgjMSiOSVbk/hFM9+bRGkUwqpHE00mAXc0PyZsX/uHS7TgFpTh4aTeO+ZTtJ
p2NWB3KZVFc60n2IKEzSe18BdR39w4h+Y8Ekkr2atFZV7UYA8SrgpJx2V1nndJUC
VAa2pYq2JwHDmw1cxgoDhl96lhePi9JCZRrrS0DkmZ+KVz8XK/GaQtLrDYW4CzGo
prHGRGPZ6Fgk3SuNMjolSHOzfmkiyym5qWWgy8U7/9Zmaj9yuLM3ZWupLyzEtSnE
lJGxS1SEMV+s6cAmT+AvgGDvMfBcqrYwjUYRbic6WFf86rp2q6AASeUwh48Jh6c3
leQBUyy6h5Vm6B9ZdeHqMo5LhzF0yLXS7n7tKGpuLohXyOOiOvIx46P6zAfKOMbr
z+7v1l9rVcblJC6XkO9M/ssbri+Kypb2vOeHvBsijsGvZXH4SLCWxXEc2/G9HqrO
zMJXQapUy5gpOgA+iR0KPsKJ28EpMC4TWNhA1myKgfa0MWP+jHj2+w2zvaTLoeRi
1GP0y8ZUVj//ytSKVezZ0Hmp+TZkYfbTPkAfJzUwF9WaLeT047S5EcAKYK+xiX6f
IbMV9Dow7nqbuvHex4SN+LqoqYOjr+XcGhMRrXqo7hawzWNMhut+Ov7XenhE676F
RpjKIkqE2QARxUhdKvpK2UKPwktPh9xDspJEoAWwiKV46xY/q05Rvfp4pGTR9ZaJ
mh10U/Z2gNdnmuRfyXTBju3cugtZ0+r8Tbg6yGie+xRwETVWhT4yom3XDl4NnrJP
o9KnPrwEa3M2J4YqeArRYuuZQ7qYpwuJyHNGKWdpfNMMLOo/74+e7m8toyPRkItE
XR+bu+LJTGk3U+K4m9RACm4UWR5jkg5ygyVoTirEg4cguFdAkaKUn+plUCJxXd1x
EMezqEggNLq8thuMqqKjPk06N3s649hG0hmCvecGE9NmmOsm9guMEc5lNQi4fLP4
rifxQhgWBWdiqXiD0zNNueaR3hLqOaFJGxXehIxzGQYwdHinB4OGD57eSGyuM6wq
5MAsWzT6nJpSXAkYRFcnaaAkeaQVDQ52HQqzSop7DyaMTQlqfLt7wxYFoXSR8dNO
NSFlpr8pFIgVuR3XApvwdDD8nVKO5+IaBVU54SC2Y8A7SSk7cXUwLjKOXsX/f+qG
8f9qh4gvzw5dPo50AZ7Kvn8KUZv9hbtpd2uCC7zrwle9u+zIjq3ipOop+tqSIBks
5S45oXwezdxxE/Y5WMKiBOGK+ig+hN2MwHWhtQqgY2PhXqNyjqOnlxqqfIASFWD2
jLk0rCpwsJ/QAkuOC/cZ8M1/ekCefu8cleGMllyHJp1e2LRDNOQ5b07hOQgvvA8r
+YRoxQz8rZFW3LHINy7AQRT8ASBr04UTSyK/DXFGVk0fCKAPELGoiZxgaSPnKL0X
6DNjYWXNeMNXnVVJMIWpbiv8FYMLkUEbJKc9vi7gc4sgXUv9F7bx/Ys/TXmPctD1
R8X1prtafdlQAjL/DOGpLQX1vSU3KPAIQU7xRRuZxiPzPjLluZ7LA8CVO+Z+73RX
DvrPAUgTf558Ca7mM3qnXKqhk8shZ2nVOlU+ZFk7GSYUQqjb3edn8MtpczkYW3bi
be3rxkWjSXgA1CZsVTlu33WTXc0iUMzKVGMGguWLegu0vuiPk1fRAPZjaX729lZa
Km6GJyEFdi3uQWCMTjAJvA4vHFcaQX+yz2Y+flHlBgvDbAn/dso5gSxUAxeh0gED
6mCHHPQMlbGNg557RKFlwwQ+Iv2hg+iiIn5Y0gxIWVDFx3sj2leDuaEDy5uRpR8p
r+WgQyYvVKtzuff8PCfgppVlG9DuH+7IgWDvGKzZOXhAu5wIyT7zCz9U1oz+jUlD
V30KMNkAp66geYmBUIqVPB5pBEKv6Iy0UBkciKov0pIVxDQUihcmy38L+tOCHGpJ
vN3VADH/Am/vvYcHNPwPLjS5qX4pNlipkfJ8Jhq+8H4w12BDzj2yfqRZHw+LptQK
oKPzKY99hE4yXbQIAIbw2bQQi/z3pnHZUCGgkOpFuHDkl+vZWaYrWXkhdDiFauiE
nzY8K/dmlZ1gjU9Bvc/nagxn/bbiQOm0NXqBa2lvcM5Yi5TihZABBb+iqevK6Knq
Uuyz+8dMI6gmqPJ2Ufd7hk/i/DF6V2BuKphK7jhs2naBYJZXDGlh5SHNFUCWPans
XqwsL0wURk3SZNHGPkk3tKZjpw7wgrSntJpAstY3WhqTvDudaOpi2cKC/8XQI6IQ
DDuHJlde27W3LRlakNQa+25mBWiC60gcwj++BD3iNtdHrbQsldJOIECL0WWuvC5x
HfWJVNXnIZmtuh88e0UFUKJw9H60fsrmcGHq4FXPFv8gntAg8+fLhK8geCjdGsfz
Prm5RGBkEr1qh2I8fimleJa11CHmIszJPHb8hbX8VWLbUJS5L7L+6ZRDAkuZgSpS
LT8lRGUKGH1pHwXrI8BruVC3bKCKPsU1xuJt16h+Qr4LEu8ln/Mg0lOZ9JmYOGqB
DYVT2zjNTrflbk4u3ZgOv3W1megVmmz/9ob5ZEbtTlALfwnfNjCqn+WgREskgzTd
J5Qu0ZxYFm/zxs1+ys43WCfRK7RSjE1sbuSj6e6CSN9zVlFgCFWzyXeja3qlAKcV
baEJmbwcl7JgD00VY3Vk2rY2vEq+waUCYodYdu8U3UMd+yCaT6z/5z1usjlW3A7w
8LO82/2iZXPATrnWxnqWQv1yNT8xwdgqeNrHWsSSA1eSyV2puRrX1d5JBFD0M/Qv
4sQuGeFGrI4sVhA5VEtilUofCayLyINOj1YIPn0CRVkX6Fp/BjKW6yU9y/V2Fmxo
7qnFKfJaHPhiAIfuFgY+QW+9V7CCloJryvVEEcX+SmwMCrsePWPtHAAtwOa6PCVP
5cPWkLXJ+eVZ8TfhkC/JlSfglpLy4BKG+5/xVTTqXMNzczn/yQXetbM6+CneFgn9
ISI3eCEVpGvOZ8ZkLdDq9bdwcgCvF6TLIxL2/OF/DyLTsSVARbFschG7S0uDHP0L
b+gLjgYNEsfLWq5afqftTZveCOjMlR/A2UKW2+G/YrZlE9IfraYizSJvQOlARIgj
EDcbunFaXUt1kywchcYvwybdFtWt8GtPeh9gRtcQFQJgsIeDvSh09LDvkr4F7U58
RElnJ6T5MOOi3sjKQeN5+I53P3LLra5TRN7TFdMZ48/K9VkiKvbWYzd2dsckXMp2
uwSGCnA98i8+Qsl4UX8PByLMqB7UtvqGbKiCbnw+eQYBSTX+iBFSuuiWPBX6c4Q8
uDvo+gmo7D7em4AET0oeXUCT6K4Obgxqu1yB4mo0lbX1tZs6c1KTQmZdWxTBXZWe
89U2M5gA1y8LrtVeDD9+yR2VwNJjpzACsSbdEBiJBqk2NzRQkeJZ5WTcoP439jCe
Ttz9UL5whbPC6kRpFv5FnDJKSd6z6Tkv0Ddo4sT8fer60Imv+dHXADEIsgjDHV5k
vKnln2logTo4RJJ+TNXK+llqNWMm620K4lkGhj2f/bu9Uf+bJY173CngvHEgzIJZ
Cz2gTd+ECwbK35wR31vQyU1WJYDDNXcmw95J0s/nkh/XIjC4KcPH014rGOQUhHLo
+S6iUlzMbfGeFnM9c7YEEVMbusgc7hoYQD1xRxGu3aaKC85NiwurfJ7SaNiqTO4j
LvBVKD7maySrYRWl5H8AF8DJ54qldyC5Ml/hgXS8PIU72COCVOfqDZAuSFksf56c
6O3mUkSVjAXS6GGj6ThwH/nbHuEQqK8YcXWeisqooAxOhqRTiGKQKNUeBll5Nn4B
RsvAQxoh6hu/kn5mWF7zsTWT9w0WO0+dwQe68BRsn6LMep3By0niYN/B4rkCaDVm
W5SepNSq/xr7z1SaOUFlDHw6i38DqdVE1/SVwjf49iD+8lpG2shwHYGWJ/PmivCH
ApIEKFwudbaEYyNaakXbENcCm2Q3m5dMrINyzFPLDQ4nRFo/wQpr9q9IGqhihzQO
VX4peBaxtisLvoMgEZXi22ClHD1wBFtmzbSfBIc+rXbirITaPjHCCsJpnlhT5RYj
dYxzhu9N8wRN05/ouJnhjDJMtlWiRPvoXsCyvcS+CYfrHfQpUluj3dlt5ifP8CUf
hgs2/t+nEcqS1fbwOr/R3Dt8eX1mzx3NOH2t83lrVf0JZp94bZjmjjN7Zh7nA10F
ouO+5F7qOAZ4b24mlFeL6Tw+Bs3Hw85klbmYHKdB82hJZAxIypyaZ8fif1P9O357
JBEsc7tUhr0Xhbi33Knkr6pfPv3UEmLkInkaVEI3xi2tQCt3431lnS2vVq07fL3Z
JBVIujh6j50QrPkwQ//dRc6UsNy53Vn7HEfDkLNHyXj8XI6CG0BCAzo3/ogRoMKy
wg1KnpiTmjWcrh5XwBM7WDNLGM3GQ4RbpExF2QTr2fF6GjDxgLKItWCWri/9NOHS
nsitcS3RxzQ0o0NvvycoPyay6xUvT7nDHIJPNxaJACOe/q+cF8B0Yyuex0XvhbyU
XUTVIxmHeZEs9fw4t3iociub/MUq6T38IlTtz/ZmRUSHiPIaz0Ua7bkFofyifvlT
lgWpTAzkjsGo/BGZwNQflSOUjY8Uco8WndXi5xwk6MHlFo8Cf3PB8tmk2DBQL0Bc
r1i+WrKVReb1/ZNJunVBTIRJZ4U8is3t2vRXhYD6fe5cJfjeDJeJSa0hXW3m0BnL
/ZljNv6uvR3nKKeeINJWpzKvXcxBAFFJNxmC05RQw/jSAwP4JP8XEWImaVLqC2ri
VpQ5Uls/OmJFPfGiEkU50ZKRfngMJCF91ZgvuBz0+IIv2aOCzWYNpMnufyjFn/8z
PQNonbS4cl2Jt3ClXZvbTZOP/uHadjm5k7Kmtx+yk1Xe3O3PPhr0n6hl5AaODqiE
TbpV31HaiyM4/jE0LSwmLunvdKrUH/YbPxJNFcb9V5uk5DPApDc/kRTaiXifjRFK
4I7RHPw2fN8aR6Dq4UhdUQZjFDanKk4D4Pbc6gWbXc5dbFkZqX/tmf7+a8UoLux1
8I4ux1XVtmhvyqXeAA/wzBkLKAza/5zNg/j70S5UNzXoMcfGD5cn2AgxIvLDJ1Z7
JQEB/CjNWHLvgxHCBZx3+OdKpmsJAhsemZkX/eVByg6VXVRVnp8EHJVYIE1WmkZD
9+jG1yCIhbF4QsK53Rk5h0iXoyIeZbUwvoFrY+e4LXH3IR7zRBhOIJMfzVXpDoT4
IKZUVjdnEFMN8VdvbRm928waai0Uj/1ATaxqPMYyTdNMwNnJiq1XADlnABXTOZTU
QUcrf2BEhLu0fgniRUfaF7zaAKAGvr7CClmtCtPaXUxDxVseiWkY+V/T5nNX9Ljr
7SkSSWF0yIKriNoclNjV5rq87heNHkw6Tc0vvnpcNqgt/bc1bkLp7/InNidOhdqW
2M32Hv7evH+i916J3aD8dVi953++prDlpV3C8bHsG7XExRNAzKw725duHAVUYeNd
US3+3Cb68muY4ATb0v9RTlEE+beWLxEXNGlzRWj/c/67GlLhFFI+QqhaF75/dJUp
nAeDuQdxKni2bHLNRNcKcdJEmkVJ87BUgxl5PENISR9Hwl5Q0v8cabJ1thdFC9iz
de/uA+qX/G62t3/PmezxIZpcjJMQXIa6TkF+vM6wr2IEHkRlEDdrN13RF8iZeTLg
R7nSZpJuecGirZxt5aaMBc9f5nmlHy2x1447FOzZCEfel3ZwficKJghynSgsY20r
AZhusc0a2IqnmYM5kIxphXznwv4peyy8M7Av+DHswpwz+OHOo6pO1+itbYv02xzQ
YnhlUJmrbbbC6UFnJDi751hw+1u2GGk5NdPtWcxzN4IvgRuY0Ljx2wW8TT4MlusN
Qn4Lw2M4H+6AUyo5rtimmynDvWlHEVmWzhewkrffgNd6odbPSrEliCISSKr7gkwA
FF3auZoUsu95V12Uyej4QOPFML5ys47aQ6gW0Ty2igytF7GaRW1dnCFMvHZRzry5
ebREXtlG9r9RP5+qNnT4POeUDLJ8HMUm5FhPBp1FNh78L7u2KRNQUYWeR2gmys0Z
nCHBtszp2XhdLFWIM6ynFmDtJ9p/u/f8Zf7CIRnH1W2BSGjtS6poXNwRyiN4sJUg
I5diJwN34Y0LwUJSW0pfxPVV9KFcKaPfBKYtJd00C4wZoxzUAeQr9bSBU7F7rU3+
ap5Cl5phSLlYgPukKiQPBd2Zd76B2vEXV+17y1d5OYgW6fhCcAtp5+yOvcfcWHlG
sU6wDZ2/DJKSiLDPnOBxtwNoupsC2fuPHZaAfRE10JXPP2IdyGOmucahqraEXEak
OhQq1aMnp6C6fxhYRdVBd/L9jIFjuVMBTLlVHsVwvYBW1+tD+BLnSp+rR9MnQRP8
cOU1j8Rm3rWvVq2YBu7bGYYGgNrtlxwlidrGHgrC5ICfkVVRDcvH/hV/cMxOHbfC
yRV8FEN0ZaAnWEOP8FXuFD2v8AYwuy6lmu8/+AGkP7V+jPdIKdLv1ccw/Ue1poQK
gXrr6mnHdtsLB8A13kNfJojRRHXoFVo9nsdT1yxC6eL/TItc2C9ya58s53gBRM/T
8g/8GEotARJPIfug+QQIbBHIzMk+XdZ2tj64Bvosl7wb/OE4X3h0Ffqw6eMLSV2M
Xmmt22kmevT3owKlPoMD6jqgwr8FdHaK9z1vnv8kQ58ZuUFKMviCmFLkzQKcCfWI
rwrVIMR5yOZwR/dcarv6QH+cMZVeUQwuqLknTs9L+oyPUMEmsJVKMWuCvaBR/t7Q
V8iF5pN6noJJkMa/434whfMyNN1IxfJFpDCfdLhli5MD5HzcHmV+/7KxK1V6gi/Y
JI/oh49mVya/tl6/VgLoV3xFS5NIy7X3o48xYsoomlpFkzZyIVofrqJTCRdqx4T/
fopfgndVzgqfdw3/gdrQzP7TBjWiSvl5XsoT/W8BKoSrOhO2bu16OUON2t8Q+66g
tHUs1tBWZeLRLINeM6IepkM21RvaAEBqdVX0nMw8ivt0LCngTpucjVDKG1pqaJ5J
buR9ML5bO6cDzk2DFc4awM1gEu+eWanaCSrjqzeBRrE6FgIELWOIMOXgSBtvb+Qg
piruDIiqKptZyKcUWoBn4fTIkmxIcERnwp7WP7jCIuyBIsR1Vw2lHYXU43d6qqZh
3HejP5eiWGYsAwMGMW8hLr0B0ZjnYi2jjT5/Lk7HcbH2uUcrWz93lrAs9H7+WlEH
5WsYw7SA6PEXugLy6lFZ1F80DD7SGQuMrYP/xPQe9Hd/SLZZOxBYRC2jjfSfhHDu
sFmOUcYiF/OrK8vTyy0b59R4/6n0PGbTWBev2bERv3vIw154ydnpHvxawR2U7vEh
UT3HEOMxLchbakMZd7nkf2MkpLYne9VemZoCjroRMESh4x4w7kz2nXxD6OnABHf2
1MkLnAqX8xGw26JQM27zqSFM/nyV4vCrY+7BZr+uzozGb4g8PYBTtYUKKoEeUSIW
NHWzq95s6iHSJMrgvw/Bmf98Fh7bhUQH8bsEwF6ldjOkEGlmJUkTZ6HlFvbEiWYO
YTOuK/ko6kH17RHEt4Cjf95QoUKvBKSzcbSu1fBplQlbiiP2VoIEvUcCGzYFemRQ
/73FKAhcBENUxyVz4p4hvvzw+1uoIuO3Ji9WbEnS5yc+I77xUQ61tSV5+z6AbhLN
ioptEXemeHH03+Djd8IDmSRaao8CiuJy+UaFRj85aGl4yi0JV+k0OzrnR3eV/a60
IKZrngn4dcSUMkf2ANKWCMLOuvFavIdnmx8j0md84QCajAGNrnnKsSu3i5SNkvPY
3gwVHo/E0n0GIpzJDCyqPZgEdoz3wScYkEPVODBp0+5LP0YhThAKOfpIqBnV0n4k
WJgbjPmVdG08hO8ydi8Z+MJvQApNoDGj0eUEnqJlCi6EQ72OdoYOW8VynrhKY+GH
fBFPUWU/CCLaz82jfFngHRFMfc0C60Gbs42/8ZwlRrBg5qd9iwsQrJ7M0nAkZTxl
D9BaThkoB+XMwA01kE+PLSu2Tw72RowaCetfKy6EuGLRViWJ6twG8yRu57jH4/pU
LZaumtrenoIi+3yB7RVO9NPT9YugnT3945RmOzyc0rbV/8EOxxSsx8OvLoaxSj36
rccTGoMjM7I5wmkf4AM+c0tE8UqWGtVFanBOWRSeYUhmMLOAzQlSHg8KNkOLi6Tu
aHM+mfFX9DCB4UemEI1++oPttAj26eSy/DrWeyhtxJpzRd8DLtHn7ELXCrWRv8XZ
Dxf9eVSoLR7OK6UD1HlNYogMUqO64WXALqzIZPmANU18dOjE8UUpIs86a8udQzVZ
sALJbQjXdXH5fjW7xNUSg1I12nmP1d/gb2T3JdM1kImdeb3XeDZC2HfhEKhICFaw
t3tjEP3jcnU4/h5ypIms7pdhLwy2j0rLpwidbFy+5lluq1Cd2qBJ2UmyuthEAV/k
dFppxAQyCIaCXs/l0mFrcmbGawkq/AZNWWUg2kCQA4vpW7XK847kV8iG8CMd7BJg
WyTAlwbAXI3Huqla81DejbzdLmvi8jqeQ2qKEmZUMF7skn/sAgN7raJkbxaVrFCQ
VDSd2vV4LJ0xWv4wNzJhAJrdB/s2jmRKWrlQIWkE7H0fhSt/4tCajdV8548X6O0b
0TiU6KSTawHBnMapxmUpeDO83skMWqYsmRdodhw8hArM0X05VKFik/eyUxYEszAz
QRNv6ZByby/rpnuatrhLTABjiHFqG7NvX10fxgEoY1DdyYp+zfYmnmBJ95+kqu+l
SKwdcsWdqU2s+bzM57dHcW4Wg63eBAmGbumiR5YkrgZbatBJG1KrGgH1mERisPdu
u/ho6DzdbIS4mM6hDsJ5WWZnXBg3u9eJLhEMJI9O4zH7EDAXiJHiazzlQ6RfL2AJ
PKrE0DkWGKuiuKNcJGZqZgXx8AgGH1QS2yhI6C5MCQ1YZidM09CXexOIugZOp12B
MydngFxTuTXRHlHag0FSXbz5Ap/XkYLq8UNjOQ6A0Ea8s3tSScilYn8iJp4KF0bI
o1zqGxrJtWvtNAi5KtaDbY6gtM5XNiKIIRzh0mak4Icn+0vEKKZVUCXjc6SAogsM
cVCUx3sqzLtyJ4ZdLVcBrcD7iGUc+MeEKbYlzKzHUWWGSENxvyfEr6obUU+UI+sV
IpMQBWHQAeFITTy6kp49NmMZJ0h5KjVVsEFjQs3vmj+QSQWLTeZIMeORhDlP8DtM
vOGlCh2AyWNOWQiWSg+A7sxVy80X/SjdQriF3UI2E23jiJqj9O33KSKVZbSk107W
mXBPdOgMbKy6bjcOsiAhRlY6nyMJGys2gfGpN0JjOsYtb9UQbo9NqFBR8VUx61/m
mLxmVZQwxIf8ry76I7Lq88Zx+gRXOHB6pVBwplwWRBXaiNPF/5YKR6Eo1B4PDTW3
wRzuMiGhXcyS0ewtjW90evTslVEZqAEXiDssPPPXJB2UC06anQSvn5+X5myCzHdb
8HfqdSJrl755ESADEFNWEGAAk1b3RN9intnoIIwIr8JzHVb3Si1Un+PPLdnlz/z5
f5cGD4Yn0bYPTrW2Oq6pkwCkCmNFFCZj+NQqRovBicVZTNcdHmsB/nWv5mGPp7ka
cHszqI5Fp3xOYi2qPTIvaQ2wKmxfNfhkGH7y+WVfBkXSsAEKRJ0mdPbShgGEsY7L
fEb6F61VinJelOAr3UGPJQVi2YS/VwHf/fWQ0buzQtmciG4sDDXXT853x/TAgLPD
HJX/XILdi9VBLUF1MuNkZK3GdvbfCFe634X7b+PirhxpiR+0CtCwGttU4GneVvzZ
q7nuic1OpoDtnAq2oYlg3t0QlSpboQ35yTUnufD1n2vt2RgMuYK6UnbFwTAGWdNm
rEKxdf3CL1DDKhz5K5cz/pHMWSGOrg36wTR5ALvIsAGx9dEtdWyeqzVeYDzE6/IP
zaEMydOUIi0WCKjv5dTllyzbEUGu0cqPyUKF8Bk8f/fXbm0H7XlDenPbmyHBv749
gZRNFDZIUDIu/CqjOiRfGvRB/+inhIv8CPdoRQP6Cc+0XidSgaJX8bcGeNGjlFKQ
JaTbfdclh22tyVJ269pqwh5/Ak7Tny1LzgaSc4SZ8o6EWliT4AKoPhMphEJ2Kxhm
G/65naceW4868xsnEVcY8rU+RCk5JwHuv3yefAy4tPGLCN3Qsyjn1IlcQ1bh8jr7
9Im7Kh0nzZ5ZqBcawRj/tx78c4Mg0tDzd2Y8L8xHFJbzh50onDVISsrXCZOW4ZM2
NMmAF28cYyaH2hHqK4W1K90ctH0psEwVpKhIv1Z1ZTfQeavGYt3zRwD+s/dVpRpM
5I29DCzOaCRxoJNaz65BFYPViIZSTrgihM26RE/DmVMm/M3hVMd+iwWvJ+O4I8Sg
uIqlcrpu+taQteqHed/fkdu6P6Zs5UH5Yq6gTeIzHK7JILlsPbAQY/ltmt8Qr7yo
kQ33ejRYqFnZXF6DXw3GpmsXGsuRbae5x8ADvlicU7D3AQrBF9p4U3BK2ztKlf7z
x5GVkYmK+cBGNjOsxZ4DTJQdGyySy7Jel1lYuQuZuKDltmzuedoufc9zlX0/rMfm
YQzGTK9tcU5SlOUUB6qD+BoqDfqeTW6/aPD1ONXbF4wNEf+TgJSi3e1RnNxLXVm6
QXEMdv1LcebKkvQt8/PIs+hkmt+9cXpRJzQZopqFn+0bcjprxZ5VoLEiRZPjg5KR
q9hSU+zel44B9d9ub4vMdyMca7Y1pDSciRwb8c0/AS97n+OwUG9vSZ3vPbAD+hpY
zweeC2nUnUjfgaOHS1b9VeEbMoFNdOEXCTCaP+WfepzZ0psCNLv8gJiBocRsa8VG
hgbWoMBAXNwL/QuZLfYKBS3nVe1e8V277k2/90cLLSTDOCY8iULOfURVKup/qxp8
df74sZRRg4KQ6ouywmrWHFuKWokw6x25esuPcQ1VIuf3EBE0dO3wDtCTVrW4xeR/
t36Gzir1t3B6gSujzQzR93O1D/4CJ5quxWGtyBRO6+o+mlf7W7DdHHTA8hojQkvF
Mo/p835owE0Hx+l5j9lmKQ/lfZ3q5j3+MN4JUw7YjCjP4NK1G4ZYApkxSTVamo0b
mKuo6fa8UXiiSKZ3nAvhkxp3KNrequzKKcQSwhdzwHuhM25KIDpOzD7ksqMCsw/Z
4DvZYXqKWaxQjQHjQn3vcBFhL2MpAvamAYROqZiDXEka82doNc1vX6TyyJkQy9Dm
iI1v+umGknHgSHvojsySCJY8fF+xRJIm4JBk/wSElYl/XYbGtGnQfF8yCRHXQye4
7fTXi31uN2h3NDDIX/8lxJyqgcCQcTom3mA2c3Yl5ueKqZGlgJpdAmoxF85hp/n+
c409Xb1Qt7QXixnA/Orz9QjZxBN+1eBB+otepsxAxLzqlMKkPfuvTMx/SuGuIM8X
QI5cZdMKIOQ/6StOQNlPMR/mFRPbH9MB2NJpEtft2UwuyuFPkd8MutkPhQ63Y74d
tcejT5lkMlMqeKgptcc13TnWEaLqtDptF4lagrvTM1k1R6wDEq7r0OrXtX4og+rq
zxkBETy3LA13Dc//Auu20EA/beemPsAuDlURpMdihmtB13FN6XHUq1EmL1FFAl2S
hP4V/mDl8vcyK2FrUt6Wn5nb9zMUtHUl33YHgAHupSYLqrMQDWx6BRcob0PS9bSd
uGgCyQIxKOPOhfR6ZZOi4ilbQRPbAyODXSY03iFaSxk+BDBXE1haC2gtFlGd+sLR
nDt6nZTTyW80MC+34shb7+YNDDQDCIdeP8uQwnjNaI7hGCvrMgihFQayOdJvX924
M6T6qnQOl/0Yy4IMMhlqfcGagh2djk6eleCkLSPa/z+hmbFrkC6JXY/yVK9UaVGk
Phjl4EwhOp+NYKqkTIOPG8nt2k2FMO/1GA/2G/G1qR3YJTjQx3YDThvqy4kjtpxj
A+HI9Gz5+YAgSwy+eO6zg+9bt/xn5ERpAwQwY51vGZCsu4M8LRmsTlsxghHi40PW
AGW8RZ280ucaIyXd0vWIHw8PAXXy+foV6NiQEGzn9/0YSoX01bJezDheMWD9oE7F
YhWxtJ8nxt1ZFVl1AfAWPoZqtuuYUNH0Q7ab0nMog0pIiyCysZmdaw9p4XBEmbhn
vvfDwZ2KSbJqq77diSAtXFaRMXUgYb+FboBJIi2WOh+uqJ3oKSg6oC4C1ObxaA3S
BqPgU859qz86c6ACqI3oXOiv/fasa+C503elD+KTImieT0VzdWtSdvYkjP42nAVo
xiJ2Uacjx6cCiAFTsiJ2TlbM8Ct4Oo+BOnWNsvw56vi2TEpVFgIfRVcEJ+Sr9HHV
OXmW9GVPhK7i3R5vmqpLUEmQx98+WZVta60OXoh58XC1JIon52qKFKbBcxA5xv4t
tTW2q1y3ejb7QRuLkjKCB/A8RU1g2CctVH8HB47KzB8DmKyjTIfoflH3HX35Q5G2
BbhwacmUS1LE62R3OW1FDggd+/aSR2vFkD7Ly37nTXmWYtdPeRrm7NxSjXKxcccN
Hg+GE8gzDNGuFW7ckyznzwjZrmD9L0kE/9jbRKzfwjCvcVSkQi0RVaJvwlqsYWVv
xYaj/0PlJQE4zbE+OXMUh+ezeYBmZxeadyGHPUJiEmZ/A9eOgZe8wb7ANsRX2ppw
HuPYSXKC77vsA447sl4dd74iK5gRjktJmdjOuBEQHlD6QKk1/6G8so5NEZZaUGhx
JIcXsvGKErJNh1sstpn0XWg5XijKuKdAPbsrQclMTDljkek1AnKxeOxO84RDIBjY
SqjV1cA9zb3GVIjEjsMV2loonAastH7BslbCu1GVHvFeyRKRFKrsRlh4Lt5rWzA9
B7vQbiyMh2OqgflKbDxKFRJcN2Fs2hI43yDY6o/FPddmC1kHRF4FatGnn/u037Dp
OfPqTtc0FYkS2Q23ARCTSa/an0FMNt6/HrhyVnH3AqOn13yYdb76Jek58rPmALLy
BITV90Uh7kh/BuKARH092s5C8dmsAue3DhRFlfT4pTHtxqI2hegWWBeCLXc19h5X
6Cyl4yg02RjAXibSdsfD3bdzwmPkQNBWiROe0pQ9hJyKyAZc/3kRzfp5BanF8L2l
R3Dte1Zh+dHX5wvWdeCo1HJGKnNamX7jM+8i8qk66kfnbFLgXkWnkqyaFwhaRmPz
XJkvh+q6lLD4mNb28Qr0mtTDetPxlKbmb7aboHBtAUx1gAnMJnqjwjnFxUrdusCz
meflxUjspCl8eqqtxhPYOYG2tCF/o4fR0Hf8WD+0vYK48wqkXsurBaBZb1sx6oGR
nVeKn/EWQ+vfs3EKEDdmWK3UB9NnCwxxs8gsHoSCisdgpQ0cNjfkVR8kdx+QAlyn
Cu3+XNdB5N75jFTifyNL9JFfBlz0kCn4r1JXcG3AjXUfq7UBHKEZM+Rp/g0gEyFZ
NVcNKwy5v5oNrVHH073PBIHSLwI8PL9hJuCoOLbQeWi5Km5rJOew0TFCD2zD27zN
Y/fOt8Tp/kFWyqiAva52gGeeG+Mi8aTm5M1HdUvFq65g5rK4iF2EIFi5LPTz6Br9
yswTDPl1JFAtYeBifVnwC2759JoQmttYVXeZr3Fqat0ftxxAZu2ZhWmorVVfSTAG
cP9iUYd5yH5FKrN7+5P7QZJcKCPiycw/fMxvvE+B8WM02JwPSwvDS1Vd5zn6P3zy
rmIsngIEhJeToacg3x8Gw729MGy1iVryEW9/FtmxkQA6wQUTHdwD/SHytm8YGx0/
4gGVzoTr+GXlcuiLwgwaVQGt5ETcSnjHaHKY6dkBL0GTXgMs2HmR5c1Wq+IebGBH
urAvffghC5H/OrsmkvV6hdkiFfo6ShB3ua7ltP9gm5ghSA5uHpH1JHlfgbOARc7V
/Ea3+U8MerG7ybvdbLn2S/8jRF3+nRpFJUi7Dms1L+umHLZXXAlBvo6iKZNw+P0p
4fDhHxOGDVSE4oqtrWwaVk9UaxSDMbJ0GjYZeDCMVTUHw5MvCJb0twToK6CxNgSI
etrgM+4iJQph8rq0dAEfeh3jZ05X54s9oJHchtlskfsBY9sqxbllMVtzs4ia60WW
H9aiAAo3KwWdTsB52Zkh3IfBMvoTij/FB3vLhepQft088RC5YgGBPEfJF/nNlTEY
w4TVuuxxt9MF5qEpgSqg6LMec2yXj2ZidDJVsEjheg895vsluLSOuZQmMGXJJSLI
MQqb+OXHwB+sfEeQmcDxmgUr4FCz8TcAdB7VvCS43xn7I4gOksEbg9DiT79dC1Wj
e9w/qfPAFlhBipxDzXnTSR2eTfzqwBX+losy8k2MTKHVAEKQi/A+UI0KmalkbhMW
uhlOiw5PYcO0CtwAvuu+VFVZbWQUW9MtpcaYtQVFWwEttmekxXiTqpPudhr0DcYL
qOJv2J41Txtj+at6UxNGBTMax9o9m93cKmlFS8P3kc8NC/RVGxSUP1NMuyYV19hN
9GT3s55gc2i8CJwNbZ98WDGYyDjeVNuKIv89IKYYMN6hsrbBRxCVw32fyvx4JX9K
jPD13JIzlBratZJ3ILeXvRvfqmQfhXFGObZNcp5K1nvUldOeqjhbO/DevgNk6+O2
T1yL55Q9qR0zANib20Q6PwE3sednQrCTCZmdYMuRc8tETmslkqMdKbbsA6yPMJm2
U1DlrV10cB8lkaRJLmNOmKAY4Y9zU0Okpj5lTw3ohfKnoDbWzA77RgIBNV5CWX5G
RqE+rst4FiARoD/FE7EUVO4fLq9LTMFuvywl71CGQw11fJFpPTS6BOkW3zafPoH7
qetCI6evzKnsazOMmjhhOOro+AI67FdXJ43KzF0izrHmP3nr6G+5igNtEMftZte8
eAY90611lg29J1IF9CDnkjLqBjWC/Jqvn/jo8x4Xv8L/pXuSnJIRwPVhRSEett+G
aYCQSjfAoN2xW6zHscQhzN1BGiCz0iZaItJUkI1luelY8GaYYkZBRokOSbb6js7N
P+ezGtys5n+XBhXFdCy8DtvAtue80qM6uyEXwmqW9318Gqvxdv6KbBuJx8ioGxwt
/XoxcsPTSP8IHbkC+wDjVzuql9uAfat/gSbcrlYimrdmyHVSd62LAivDwwHMcFcN
b6De6BxPmguIL/4smqFc13yxtuSmc9EUBATOJKkdMtVhjmZAwe9VN08EApZXNgIR
wQ+vKpFFldCMnmS+S6Sgkmy9QMm9NCt86TgdHJTDXeF8ne2XUcfyAVQn5W0uyTnq
SuKq2f+C0SmPUPYKSs8WU3NIkRMWJirmn9Uy+tdkioqel5lMkLg5c/M5vGf6r6ql
6MR16ikqkYoOFFwFl9uS75k5UaQ3MnuqtVxrKnBSPUZOhrp6IyQI1ZZt1j3XsPmQ
G0UFayi0Qpl7KLRRgE6ZRtEk9n9daEwHY53b3pHXDDAItjjrjcCDGAkhFkZTChcb
I1/PERzN2mKxnPnaA+sDp6EXVyGhcSXeuK5RYd85V6r5CwjGNghcY0pZczcZZ/ve
5OAom7sa/1jilIZbJFPmoWHF0EbZX4uy8t/CiaBFnFK5BsICz16Gf6xZE8AodJEZ
L/FHYyMysfGfNcAQKG+FDfCzZAS8NfyaM40a0PAxMB+8ZymERuEKRqSDheAwFAiR
f5wKvWYq2aVeprnYp0IXCk59RTNAfq0eQN/nL9X1o7lBfTULQG/9pLJfdXRACzm6
pRazEAqq5ZNLZswC6jo51n4+xQZWGp3oCQgYDfkXKPqM9tGZrQf4b3vfQQEPehnL
Q6N8tx0B0qaUUNDy4EBlGvHn7PT85OoAwGem6b6FCuPi4pOfrtiZ2M89Jlko9XHf
5mDo3n6AamIAHBNs70/to1FVKjxu34cNAaoTs954kEDoSJgR59D0B35YqvL3nuhM
ny/Xd2zx/GakSNsetmFNmjHWRm1H1UgtetivtdCUUCtKt0/pyvzNI44w/FWvRDWO
zww2+vjmVotRBcjZ3LvRnWXTZWefei6DQMNXvqluzwsn5CPnRLEVhcuS3cy90Oeu
C27XtdDTzqJGfs6gQykU6KQN1Ld6cmLTq41uCH85JzfzNBtm4JESX9jk8RG3/N92
cYNHuJz19vmiGuUH3Pak26r976055YxgpRgFpqSLpvvuIxeQHVxLc3eIb+u077ts
kfNrGNo9nwsiUL+xRPobKzQQawqNtPs3yw813LB9zqUaZGwU3SFvrXoC375XjJt2
l34Dweb5/fK+hAlxf+N8PvifpDFnbOl+FnHWridYg/DsBIXj5ehuGThLVIQpG/Xj
hVrZBvWvvSbNCLmd/b9xDa7JxKhOv+d1Pc4bnqM/VfmaZzEh6OMm4YH1UDyy7s8r
V+E1UaR7Q+4/g4zoe0qLtB5T0UGU/ulfvMAfokms/DVR4DnpOVjbWOWaoo9uP66C
SSNHwanbmfdZL90vn9ALRd6eqI5UhJTR99XtbJre6pGVS0pPQ8jDu69kCWA33f4R
g8SoRi3OwTLk+sCMs8MlZipO/TTbJ2/2jRK/VR323SMNS+C/krtVZe26F3dFTTgW
1BejL6kJ2l1m3Edop2gUbeZ5cOsOF13fEqdMnAXJ861R6s2xWkHDgxGqQbCpNNSV
MHFFD18r8Dk6R2FHNOqZpl8TTBwlL9U2yCRnPRFEHAKOlrm3lxbDnKbYvrP9KcHt
jLToApjXgMw5WAoT1QWu+OQ6RA1K2as2hwy+XqzoT9zozZVK24PryZWP/xkvXd1K
W4oVbEEF0Fv3+pK8H6AGn7dETvq6YuPQ+WmBDAygUxe1t5MiEVuKWZpRtm6iGMlJ
kV3+IjMg7sR9oieMVaKWI+aFw2l/lY0q7ha+FufBO6j9sPrHSz+o1r6f9cJPzmnO
OkspJpDBTSAKsXd7yLrtiX2YG9M+F4ArR2ya+fUi0OC6PUOYpd6HobOqv5U7TLMm
7DgtTCAf2N1/Pb2IEqQiHg2VyBs6G5xAWNVZEfIfJGrI2i4bGB/agMnbtlAbDk0i
itNsaqf7Wm1vpTpvC3nr4/vJb2K7kXSnwZIDzn4+Nt3/x3hCmPMqdp2k6d+cZOlg
vs4oDK4NyOoiSrXTnAK+XV9nCke2+W1cWbjrD119X6tIIG0OkjFSm/GcT6MLkZ0M
LgFBjh2F5NKdLIEc8LL62cRVVI1nFZSt+nvF6cHPyUKNvO1qoIl19Ieg/2bQtkB3
CmKZ1srZRB+Lw3/GDpZHUJiFxq0H/AsijGdsiTt+vhlvoL4iLtGjluNm6wIsPqK7
8OKUgQBWbzAFZq+XAZpMWBplOpsGxEDG3grdYDMW5FDFFdK7mDN9fCKR5IcI/N39
yX7N4Xz+Ta6irvNq7b+hZb/FI4WREWyQSkQnZjNmp/Lv5C4EeBDEu+nDx2WBUY2a
ZLp0lHvwyJjUcODr8C/qF02c1xg6Kpj9ZvZYywBNnzUpChP6rg67tkz1gSR/BLcl
RXxeXsiIU/816IgW2fpxPSahO78Ism9P9i+aHkyml5ynWlU1386GSF1Kv26kZKFx
+HyjJyRjC7Kz7rQOA1y4wL8VL6sKF6GEhsL3rAskEfyLk30QhWJoOWF0rX5XzhqN
nm25hNsJwM7nOtuSXi/K3ugSDmjox3SZFg7NsTd68LHFuU4aKrM0P0JDextV5pd0
WgcWKLqC1whMMmK5gdytKE6V1fAwOHtBlAWL06pcBPDI5DegpHIn/v9xUocXBlmq
84qmSi0kgU6lqW/ba7+SLUWnLSiAT34TMLQChylS/1fN9woCJZfNj/rhw+ON2Ufo
5XVQiLj1GCvcljsooCBVD0pE8W+HjUCaUs1nCUbJyrVId+dAEX79Xsd7tCV3c2UI
WXPNgoIG2v5y1ZB2n1nsJ2vH1RdyyjJL6SHHOp0JiWRWCqJ7fneeqOiy3JXMoXCz
fnRNvAQngENU6RfyKXdLkQTovmerjAnIGrOmP32pKpLmAgyrwJ7bGocIoy2b8FAn
h1V6W2f0aze5dXu7+hzqFxhfQHIaNsT5gEVjmUsNmDZ/F57sX0aZyAnyBO73AKIT
rwAuSEB1RJHJ+yw0inBD/sE744uCi7WUKS8cPyXsrgSWtUVW0k5SbL70Oi1GSjHJ
M6ICnqzqe2lnUcXkTMuN+2srj7QN7DpvscGEYK0SEKen3CjjN74Weeow98WkURfs
hiI2ofZN3QxLyJ/LYTwQw8rpbcs7fGaI5mpWF6Mj+CALaBAwx8wOueY6M6x2AWjT
dkknGAPb3h4BxWCWg2EEdeHXDZrbdk4/mt+u8sHO90YNg58HI4/nIwYVCKxXEbc8
pL7oDQcYlFIoMDaXHDcgZ1A+tffe62mKzHrG43t+IT9DDXh31ywdUPUs2Q24qiud
t8LtorYT0hEFNoxlSfLcg3nfPBFY+Pi/fmXXnSOmST4W1bh3OpsHRQzJ/1sTPHye
dfb4mJpsjYNGDmSba3fd+DnYcwWwOCf1KsYhZN5njvYYhoO5AAf2mW1BUCq8bh/z
1MoaDHvUS9ZXwgSgDN7UdCgergRJdvTRnqE5wvNqjIpfJ0bnPAAK6w3ZpinNszEc
1trDY3ykf7Etimc6ugaHY9p/0cAHq5ehy7rAl3GSR4bsTGulmvNbJsiyZPUUxZg9
J0t+T8/nnXACcE/nrM0vWZuWB8KYXvmAqYsjy9mo2BvFU3yHIN032TMudm18NV1p
m73cwB+RvSRUwFdvMtgV7sXhp5O0OUJiTHlrqwSl6vOcRic5X9MbBKK1jmQT27Sc
6SD9FzynLMvZPmIvWq5mXX6TYA/pmbRcoQTdvjt2tDrznQj5ytH0dT44qkE07LWx
XXj/4uxYx230G85Lg/orr9n90e2ntAZR7s+o4Lhg71NsJ6DIAQO6fOEiOAI3zEv0
d5r+0Y3emJd4kHoNpu957jIVp7Fm7h+cpMPM3zpxQ1BLbabkUJ7mwon2IzLG0chi
PIm0LUJ8SZYQqaosFL/hkQr3cNN2kViwGDOanljkeC9SLGRZ38KNho7H6X4GxA/O
ac9YJSgZFuVWcOOs9BeHNsUcHC4+nkS84zl9I49mbngJnli1ZrJBcBUVnyY0mzyF
ErwAOoo0DGdWlFoCg+X7GnEWZ27T2v/8WZ1RK+w7Xbo3y151j6hrNfOado3tFxZF
FQdp/CfvBKWt8HEoxhYIVEsaZ6u8AApQ8dr6JQrATHIUekvA7QlqFbsvy8GOZMVF
V/e2Ytn6vbe35ITJyhGKV1KrWSPcvCgOVb7rnUzL7IusHfK6k67TxSzKdzvj4Lyv
mKnuaVxm3XKG5cioU+H4tQK5sn3OqE4bzUhG+Gte2Y+gBAGNhBvrYh91fpssTJSq
WcA4Y+ZUt4xcFsNkgeEjy5cm3LPsGBOF/sFq0zDloIR1dFkxACQ+htdBqgbl2SNe
b1EtMiFgvK9JhIfxkJXUvmbHZawDy8qJ//vmh4wJqcx9J+2OryymzGJH8k/Ax89U
XC0oNvak50anCqbmmZ5QlLF1bCxOuWXWMHNAXaEcu7yZKS1zkf/goSuyng4WGpYH
7zdLLf/7/OXM2P0/r0HIJBY2etJVrg80xyR0NTMBeB21jkWevqvtdxke/xunorqT
Xf3I3IZGv6Mh6dYK/kVDcV8VOdHwIeRqzJqExUyqOM7urQsyxbtsGHEDnQxCWeRi
Mev2VWXhcxY//BDyy13njNGfUSGhC/0aA64aHdFjesTuT0QEqQ6CO8rcGhIHVb0Q
MPOIFg+iDKbLi+5fstG73kO/pq8snKi4m8sTs7AOd8fUVVeZnYVmaNZtxtjdQInQ
bnL8RiyPkCox3IZBvs1srhtjkqlJRXnHrFaF7Qi/YXPlHt3IBdNQVIidRJpBRSEp
gZVMgipN0iDmSBF1hyI98RyACQnT4ff6LBci9io1Uga9shfIAMisZsU7pAcyasgm
WQPEbRhKJFvIHTTF0rCdXOCP5nFWDCy9AgVv0zRVyzELOeMSsHLj3ws05yaef5Na
3usfnX2hfHDBK5zTbQTX7LVYBX9KSV7qWo0lln6SybItJOyYIMDpvXWfqi2bbCg+
tthrVczkQ6QF+8fZ/lzSfLgZxWcsA2NM8OIKJ7ZTN1ABAwUAut8pG6GbUdltJTjO
Ishv+tepbHwJDFgUVCVlYSOXJh7ht2vpuo7QrPrY1W6ZSOfMLGqnJu77KxEaqCxr
E19xUocjWWNfW1RjIhgGOwaZsoJ341PMDRdayADx/Bmlkkqx5NyIIT8bVf80cqTM
c2w4lVao9ug5DPgzNLqygxB++W9+iUBtSGMQQnUstSCgz5xeNbKT4ukcL2H0ltCj
xABkJsjr/QAMXSEGZhRi/ilviTaWUMNnYlPF6nm3r3d5nEwF/P6sBEYx5c21IRvd
vWc62C6r8f1YvxEhmomMqD/TiaQ3mOjTPEruyS63Rarg0u0pvxY78rAvtokfT+Gv
9e4k6uOX7/mVD0NOAZOW79EixarEeL7eap+aOuUzdZwjlWLJPs2+B6GO0Nqf2nWP
LRytFrqj7myyMUlicY5AmEzJRkdRMcpdXOu6c/9AtPUTZQZrSg9us4i+YhgbaUte
6BPtX5DgSixyIZ0yCIzP1UIgrcBxbhbMl5rvZdcDgTeLNDIieHkCz5GPBUm6IaEU
bZjifT0F56xOPODehzz+e1H+r+I32HU9CaLQIFphLyAHejpD9KQi4FavHfYKfP7Q
rrP0fWEfgQhlDU3VOcWYPQ4gRw8uHh2E9Sf4oXIe8gRX8mjq3EldqPXtSlIvdWSm
sLKgS6ZgtB3FTl3SFw+CgCMl7wanqUMxThQmnJ+95GI0sJOtN0ZS2zp7xf9aQRMG
YLJJ7fndhDNRxAifJr0d7P7EmGpjakZyf0tDXAb1lMLYc5E5IzkvKPn4krI0N9J/
ssttM8w5sIfc4X06Mz+zbfU+N4bBNF8n0wis4Y19b65BY/FOqKi5E0asxWNaNYxp
+0psKxBBQik7yh8wVDtg6cw8m1PRYsYGmB3BKRW8WCr52EmPBa0YyJLHrOdojtUQ
vgIRcS29Wp2FkfNbU8sdZfhGjzMzjyBFcztWith3o4mL/0XVUs8kaTPwEVDyIYdY
nsFNPJUkbZpfiPdZNdl3FXQ2fYium0J7dOeqbJMmXB2/ANHMTBLZ28/63CCiFT/h
BjGGNbg5xMCdYpwj4rX0nO4E+kIYBz8hSACHIL0+NFNrjOYvSV+j7wAe4gZBVR+h
lJyFiyjvpqRuFtbuNbdNa2CgESxvQmRHevY3H54LigSiz28EqLMwiwxbj1VDNPbH
qsg8T4fn7C219Jq/yJFRseoPxAmsc2rxVCkfDfZ0uFfSSVN5QLK9NDzR9jUZGgM4
jwcmFmE9XyBU1qX4oFgDGWqmH4EhJwnYqdo+0xJRSeORPpiy+ELnlZYCvBp3MyL8
IlGM3e6qBYw8wZCtn6n40kx1cj7VK2m+FIdTsfDS23kyolTcoK8NLPT2oaSjEvhE
rUDiNCSBUtmJYSP5x5Csw7G9wJg+o/SW2IOY4PEPkOn5xJf14jQDkIzPGYDLqud5
efx9mppL77vr7zw5Ab4jJ3XiNoNElvvtQiou7Zu2h2jHtRWldt+SRpdcDoNXLZdV
klf7FNjv9NtErr5NGoqcMBuVWDOUpUoqBzIxmyg5DvEQZNqR3gPazp/rcLIdjAOB
Z8rN+nRRQyQ63wxnp3paU9IjsOejH223J4+9/tWvz54RqDdNiz5iN3ALNzmYrpQ2
RLZGu9jF8Mq9J0+7OS3sQtu1L0bZObfpJVa4myUbev2zZaARc4vSi4ChTU1WDFZK
sSHrp3UWel6nbydf2Cl9Y/PjteVld+Lr+rlUljPZh7caBq9s2S+2lSlNgyhzx203
ZjAvRrb23refH7iTm15EDQzF+MjC3xBNKeFp8fCrwU+CQowKA7Y4locIZ/garg7/
x2p5nqpU6a00XETjK52L7wJDeJln5/NQusNIdhHexoFUCqzDH7YPtecKNmYZRAVo
vpSzy+Een9etOAZpGvv3rS6WLoslpKHCnQEep54cOg55eci00dfd89BNrZsJ9fP7
6iqof7qBWJT10XO3VJMxwJSUNiD+d5bnKu2s6x5uUz8fXG4Fx+1vh5VRJUXuguos
j7en9iBjAKa2V2noVzS8U5IgXWhmBTs5k4GteLMXpyyQcgLLM7ipU1AVeCQgFWG4
hhYr5QUPfxfsceR5anJYHZj19V5vNVa2qmQrzKmqYUxDvBgH8GC32Bvq1q+wjRD5
f5mc2ZcpObflFitdkXDVYm/VeqlB2sy/OoQj0vN48ojlVfgYV/EXEZqwV0K0TrAp
Ctcflk3xGWHlIOZkEtgFwIWrVKYik7uoOfPWPuIc791YsTyh/ZdOIX8WwCic1SDQ
2JOFbCAcVJAO1EOA/bEMlMHcQAM8adR9sbq4fi6hLDm/Ex93/t+R5yhv7HLUsIr+
FxvWbFQEKtrl1PzR8TuvQ5aqnw/8XcGWNnih1I8GCiC/h9AxnsX5Jsnt+/Ik4fUe
9/nlgFNPpZZkwwFadVkdWW7tdBFS/ribz5WCC1Cqj46KV1N65yhpoJtReB7v7CrC
SvdB9AKu4qFqb4na0SEnYzABx1+qPIuXmfWnu92YtJ7bhT64TQZjD2rRQEu3Bhle
K9gcd7+r7ptlnF1bk++LY6jo3S4CpYe9MYo6AgfVPQQoLfGNPBTjd6PU+kniC8bM
LcUV2qbnnzV3DMrGLsU4ET2ejKQTGLlcEX27NLazGxrR8W6kxe78ftuqBMlGfpoK
2yQaER/JYLtyQK9jFBdP/ynqSKqgPEssYmlDHY/Ngm0GW1PRnKcFogtoEKS/LPGt
r2tsD4Vz9EM3sU1g5FDWzK3DK/gMDYLiV9ZIU6tv6fLVP8bSaMojmbUY7tz+Z9m2
qvykEssIG4u7+VWZW+dQnkHWWIBJzIYHv80vRLc1t1yuFcT3uujnpww5RB/nmS0i
CzISU5kSRuRSOgYq+Fs4bPdig4YWa0jq5Df3RdMPlaoMvpPck554WLo4x/yeWMDT
uyC3Y3jaUjI11bOSAsGKivBaXijJniwDopam2UISPJZudwF8NmcwHNQBCz8N7Its
yOoZTtkUsXAzQl5HjsS8vn07qWioMpI+iNkNfO5tfharoYmb0FGNrx1t2sjOQEKB
IzS16Mt1YGwsx5LmUzUpKSYeZ6bhaoXlG0TDAQmmLa5cBx9tVu6PasbN/c8olYvj
EWUbqrw4ITs4htoZ/bYfV97Rk5ecvF+czb30DK3hfomT5cD5l0hityslssYp6+iF
1eH+sVpYCjTf59vVcjTNJAp0ohUT/QIrwmdrB1E0CcVLAnG+5R6zRsQE/ujs38Ak
3HFYoVV6ilqj+CJqePtAQbiQ+mDa83itr12svly/xZIpYNx0XYClFKkH6+OpNTUk
xg6qnTSMY8n4wSyy6D7wDLTQUSfeM/IgGnUZ64JighHCHDOCIHYhLM1Omqht92x7
zwaBS1fBqkCoSDbB4HswUF9XUDMVs0EDGTGWvrELpWrJEML8zUGpIQqf/BEMTH7w
3xFRftR0FcbaFiWL/YiJKwcu4tP3dd8L2J6eV4hHO2VCI+X9vwxEI5AqOf6x4PmX
tGW8QDt80n7kRlXRXWimwjIZ3sIi1Q50Gqz2gTG3uWvVXnKTNGt2fJyTuqNIOU+a
AI1lXwFout1OmqwarRGppnahKPFrSuNwvU0Qfns04rVYFJLj83vIy0zFfm9UUw4y
Qag8u7wTEKtBThVs0UBtKZS6AdFWKq35HHwzlab00n7qYDsdIEMRjLJKV+qVaQA8
A3pPbzZ55TTSZw1Mj4DrjiqC+GZHkclOVuSeAu31CK/pW+4nSPCScC44dqwQq3M5
4CEVx8p5fdar4mnDyA4A58LYR7REE+gvA5vCJxsXb2k+h1PVhHyBLnV0SF9+CPSd
uR+CHOUfEqEAER+eB3K9vIif+4IFtYBY6wCYtazc6TKHJ02y9hw7bZI/2MSyhX1i
vtPXw/0RW3jX5F6we+Q7PwxlCNOokd8Ztj5J46c5SyTLrv1ahcDbl+GMEnlQnX8J
3qBbMZRjyGta7hkWlY5arcKqBgg1vgUdtUG3JhWSwcOD7bRZBqI1PDqhbXUmjxUS
u6E6rzppb7JhK1nrJSUmt8kno4y6VqR/SE0xxIOlVlVazFsUVhpsqTGPi1XSgn92
+I3xReRCp4r6r4WFmKm7tQqVaIeK8ZTYz1OxeFzK9Njn1McSzUwTq4w7pvw5RhD8
Yvog+ENM/lhUhARXclJo0Qh13ajd4wIk/bbIXiFV/j93BJWTPaCVHOimWTYwrJ68
lF+FmQH9Xr3ULWdslZr6+FHIsbv0ejeSKkMSljaG1FppFu2wmF3je2pZUdVADydC
tRSULG4dep5S9cNqpthbqCQGfWeqYOiQrrHzNbGpEj7vMndv1auHmVwchnPoJLrc
tY9QHfbnRIgKzQ+vR4JJp+hiiXPFUY9tUZYjwuhlW1rv2AbslF2JgLn14Mzlu53X
pZTh6LE7gVWmSmvWMPejYQQvSAob1i8TSBA5me8JO3548E33r6i94k5Ypdv+Y09E
njVfp7F75rZ7tLamwyfV7YPlpKJkJmu+oL4bTmpurUjlUAkQ+6ezXslK9QLMep0b
SdUKNwXV8PIcbJkI8xqhKc5+NJDQ3ag0O4AM8pnkYLZlQ2nJFF0xlhWrMAKXVCwJ
cM/TbEU2qwBdsHspYsqQPYirebkaFWl8lrNmvllItiYfmNFofpLjiorue2zTwFoP
mOBnYB3rwZcxSmLAJCmybmLKnawFVH66zvq5tUvOo6eYXzUfCWl5ZQt8/vIxYNzG
f2AGf/rWP61ulWwjqa/AlN+jOFf+xXPUEt22jrR2T5cUs4OvBSQ/fpfhC4YhMx9F
R+NLfmbxqkhL8iF0X+n8WC4Ukevf55pi5kwlgIRI39ztuSgm94ISlTCs1gnLHYWr
2YKi7CKJ0ngjEIsd46YFa4nM9FFhzA3NnLZ7NN8sYP1vPo33cED5KpgAHx9diJMs
KSG4lWzeRuIzRmq8xJlF5mgrD2h9H6FGrFGWCKJWfjrBcA/Q3UVHNqQQVXwe7juf
HGNnCjKwVle37tsNf9qJ+WFvM7P2mTZo0rSvyHewg/k2wcOL/eAbf8jURWZm8n8C
7qIE63yJgQjImbqqs2VS7OxWTciz/AZ7QAdXeNGcov6QuZPqMwGbrBnetV3V+JGq
dWETJLIAHR2pjV+HYrD/hSTz8fT0VrZAybfey2MwV/nd0Lg7Os1XVBjKAQLLWZxp
mDywIK6TnBVqo7r52nejH/Lml3Bf90x5Wlf9WDItUWzDAV7KpS2vVBUPc8f8nd9g
MGhHKNmKCSWuCSzFL7i0FUn7NW1huyKUrDDbmUP6mHco8LquChEHYrIQxLGEYkPr
qeaV3V14w0KMcfbFeO7WSWUpXh9WiWZHOGbYB1dP+iIztQpzwjkspKmo9yNSFcly
zwQrIKK7bhYd0RqkXFPjRk4F/KIA15sY8kTp3w97aIVPw9WE13ZTiNWTBPB8qyM+
/4+OYhJpKJVrGbhBjH+BPamCJZRN5D6DLMBXXQLnzcHCDtTDcRNrWfO0vh1Vt1VG
Jzzmp+NrbOVeaw+pnhUfq47h9jvqEMdgxcGD7qxECys2z0OSQtVdfKIQf8oJUUQt
1CFJWhBI8glKVl77q4sZgZ371fNwcMZ9kTYAjYH+mgR+RifAO5twiP2UHZi4Qwfm
kCbGFK6EUOGfhNGU+Wyo6VlabELuEdAweXj6XyHX1DJHWe/uybj9up7uo7o/7SMH
840m6ceMReXVEMaQgykv2s47kF1BnhsxmYs4LCKJQao6tx/Dnv4Y9FexxEkHrftu
4q2almGnHFGwLJrUi8pcq9kbBq2RU1tHmgdVrswF38W9JQAFiTxwNE6QBHiae+ku
gVIsEZLDsM+cNK9vbdwqA++Bp0SWj9mNCS4IqHBBUjiF9eV0fwgwX+djSQSJcj2Q
E9+iS3+SMJqUsq5CsCRLo8f/ktXjIY81ajoRZ/dr3JUiIUeedWY7JXo8pGKo+CmX
N0QCVNLOmWeueLFJaeyUnPlxonc8t6hkPREFti8vCOR9um6WD766yvf975IRdYo5
GMcVG0iEm6LQ5VQPJfzZAWrwzjsX/52zSczTuFtSmrh6KcFmV7CwINYKXbHXSxA2
/lDnz8xmB0IT8q8cIhgnqB+xXNTEpDeKJDCY+L+GouxMiu2u24ahZ6ROuHQfoPf5
EdBpjQrStyroTtoy6gZe+po3S7mTZLYiludlkF2e8X1aNUllSJ+wleUdSBtyPYYy
ypeCgr9Ye1CdEFpAAhexj99l1awlfvwX3A7p93fKZa73vjzbeNdMemi9gA8VChJ3
0Y3GFwA8hB5fiePnJILXvXPatG7MX6wV/8iD6tzTtXhYIfQKZAKfAbpWhW9NFusO
crWf0rulRoVHYUjHsrm+n8au9PK5F9RgFg+Ij/UWg7KfipBMWn86xea9p/cAuhdj
46LTTeBZvauTapq9Ly0bCTgQyu+utOakHcMTY/PpyVRO39zicZ2I7G3n/wG2Hgcj
5O9VkzF2I7L+wdQTutcQ6swv9ciqz7aG/Awj3dBZeo37ihktVmSaurcq1r/U+XTW
ohvZ9+DlV4oXBbr3+KbeeijbzIrpqNTdj+Sak9vuMTgxj7Wosfzrg3xAbKkzM+hW
42J8gziTgfMRoXUQtqo9MWM241zcRCUTlpOCr+vdEFN8KhBWI/pWqhEfwrGzc6gM
R5Rli+PLUUHnoQpKWmidzC0rKh/RxhsGT1gwDAiaA+oLbZ77aunYdDv7SSRx2+wg
ghyVK986dIOdU0pF9LxfiB70wlWrzp7yf7TrI7GFsPASqEaIa9G8NLf8cXeBxIFi
e3zf2Bd9Vpw3+kxICGUNxiAb1V9EIp+3QsoOKsKd/cGX3wCALX6uPcnvH+VGcgMs
fxaac8d0fOOV1F1iJ18gD1vG/VJtIHTaTVcbTJ3c/RYuv4wFlNwtu3tkn2ZjLHLR
qFfyYvFdGBqATCbXkqx4mbsl5NENCeE1Fetaa473lq7pHQo/CJZzPphOVDcFV2Tc
Epryof4jszuNRp3NTDd9eD+ZL+F9p8eO0vwFGRhp4tCGOX4AzHAHmPxXsSm0P2pk
otrQPV7ltwOCqg99U1SPzRMSbgYSnUqa0E44uw8/DMNn0KAA5Xo0hMyIREpUWJQM
xidKQZywrBbXWTTts7nVUk6dup6ZME8xTzoVJByJcRmdatkVWbz/mJBkLZDKffc8
WBoCb8i2kZzbkiafo2GexP5/ZMt1sktSV3EnGTYTDT/R/fe+YfyE5U+m/1ZDI8G7
6yoamVY1MhYfgAUybdysJJYix/j0Aa4NpLYt1Wrq4N/s4Gj3G7aOG/GgDyUZbut7
dkqHlk47C0Wu3gK65wYmxozo9Zk4Sv0Qo4NMqMgrlG05xCdT3axji2k3s6gFXNWA
tCOrddPJCtTEWjYV/Hb1fNBKo61orZOJCbTyutuijiX3t3LaYfuj/jqVPW2yONPW
BfDrfXW0nxMUuoyQLJF6fdqhSMkJl2R6iPQKetpKXE0pJl/fPHvUdtvXckrFbl71
i9qzCWCFFIE0ZTs3xwo30FrH0O6sOGmH9yGA45tMTqy/fKkwHXohzlK+ZUERYYVQ
+vn01zRNYwPncXdrWSRvg/bLACao1fLdH9Bm8ysU84okS6NROadoIsVXEixhUQXI
czAaWg86ViWPj5RO5EX8TLBlcR/zhgoxMNrZMEPyB5Br9k6FllxT8btLJMaRy5vE
y6s8+P66C2iLJV5V3B9rShaO5RN+SPYytysFLAaB0anNiNFOQN+lDBr4ghycgAgE
4OxgwcijwCrpEesfkouNNzwS/1Ri+OVZU3SCQfWubHZQBUODCCNmmNq6nT4X2QhT
caUPy2qnaC/8XoNGDhtbJKn2SD5Th3Jju0nlytz5JzLYVfywJFiWQOGqX69g2sEg
u7kAXn6g8RpumFh3YnooFahuR3chKFC2YNrciZLeS2riYPkd5ZbJ9PWpkiZwrjd3
QLn8fZHzrZ7H+NqJapiZ5mA6PtOD3F+QkvAL6NpPV7DWLzXDPHxOic6OPguRS2CA
q8J7GiUeIwPtee/zFMAv4iHAlRk0xD14AN5RmjFGN5HFGwkbIE1mPpJv0hW6gvLR
HBntnwgqNYx60koO7i+7fZ3rdr0Iqcb5J9sqGRz+eROAIs5NQ7dDkQdYw9vSSo3o
C9l5knFodJUSPUMeYnNIxEpewQ2o6Pr4YmFchZFiC/dTakrqHNUtkDvfP8ukcsxw
O8v0xuny7hpLEUNmdTGL5BsGpNsWRybSVXYkxZ4fCaPetMJI571Uh/BzXGaZkBB5
47aB9xF6p7xBU5aAICMxTiEoZfpS7sJoCcnuAbdu8YYgYOJjqgcESFUujviPAwib
+yvkMdO6qEUMBEbDh6NdGKH5r4A5EC1YHlx2366o4oYoKGZJ7kCrH7d6A4FWAirD
oDsFq+00QXrNE6gBu190P+Zb4/CZdseihArvpvc2rk+noIWG++cUEGx2GXQBNxDq
H/LiEwpofp9ouU0ZzK5Eqyzu+S0bFg1ABAamnHuGa2+JeD/kJu7Z6xOcC/2HW2H6
0NsyKFK05t+PTLy77qgic/LwVf4pTvL7OX2C0UHkjojZ9MFsMyUU/9NQmEjbOF0V
5zwRh+89vlClxI8QzMP+bTSGYVOXoAnvZxWB6Vm64C27e/wLDecg0xeb2XKPY8ia
eTBAuvdY7tzJ+Qyt+CPhIbsAiY0hACqd5tAZgVlHvqOq+pFR0kc5VtITyR72EOMg
j3F//mWfD4m2RzKiXqgtgTsR7dld7dx/WOVunyEU4fb+xpixADsKct6VUNQG9r2S
N9aPhedreuq167FKoJN8oMA/qbz1Cy8WeuyeMxP4OwoaKt4YkpuAOA3Pm3NRFe+4
HevP+XcfcnrHhPRwVGdSCpgH9Q8n1j/ljDU+1KfqyZWFCMEB2+E1/iHOvNt/kaU6
a4+mKG/J2QBuHyJOURybrLVOpwCgEJHFm9DOtJYQpjvHpyc+QQtF10JsQO4E2kLg
xDVPeQzUnhE2kH8hLGBXSPIZTjO9TqHlWtgi7Ig37G6a7UxGVqb3CJpn+Sr0EbNB
z/yg9oy9C3MvjqeE9/pmjxESnLWVPIO6+Im5eFreH5Dyng3yqx3kw7fIVntZw/mQ
jG+7RA7Yk/WCCvmr7IyulpU2bcCZRUWIVfvgwSeZ4uo6Kuez80TVwjt2yxMPHjwU
nPvYhylfyH2937CrAEBcKngv39GRAqFe8LlVJ2t7N3z+ZQh2Xv+/RXQEVcszYs9Q
c5Vd+aubZHbso6uIjX5Z91d6oskm3XXK2TzwL2qIMwHR76v0J1Twrhe1iejFzkhs
MsfMIgN6Cazhmayi3mz7q3/mkRcqERJ1krgz/cbv+1b0nZL4HNwv6A8cBYGDhhfF
eK36+O2bRuo2nPFuEGbWb2N2p2au0VsV/nKuI1nbm3a7wakBgxH7lDcXc/GWZ5Nj
Kh7iABUQ1e6ZA1iPM/nuK9Qv0En3Z264rR/UoKdcThrEsIwxqvmX0go5HiO+Wvos
LFqakjhTNtytHH52SGyydrPv6/g3a04IU0eB9226wbpM3C3LTKBm+KCfG2A7/xdc
Bh4NzIO1SVzG8hkecQ0a4IHbJrScJ7KCvkZhoaKY2jt1Vmkzkv1JqKexCk6GL9k4
QlK/aJc2Wj5M8lobYrLblmMtHe4kduNrNIyzepp/Rsz8tDI+lcLLdST1zeouqfl6
6wSEUZUACZlkvOHW/G6RbgsrezUykpMvqHhpkUUqReeBA5rJzyusAX/6MYltcLJM
dQ8dkyQWc1xONWS7dxCuGR8w+Df83cCwAtg/cJrfbY53yrHdaDiR6KyQVoX5WVvu
zCtMUvAzSCB3v7YK+zGsCjPHGArjqy5KBbUlMADWOTP2wR2Ia2FgOE0wVCNnwqPy
wb01JLUfVNLvSY2JKXPLmDWU4cmX1u3iQ/M1FtPbKeRg0NyP8FFnQsPiFAnWGigb
CqER5bl7uwG3bEXXImBf5M6dKTy8MWh4SvjgLeGs+wCH4+57miw9uFNWWmgoFjuc
nCaxHfBzhlnm433wb0vJ4wO5htGi8njmibI6SBd5LIEIYTz3dkNG6UuRsdoKXG8l
Bue7qneVHZExS0aytDHo4ody93mfu3TgKzCyjU8P/IXU4q9nkANVn9DG+olgTqw3
kYAPcmwV9iwV+ACd0NnipC+eV9iNeNZDm3EaJ4ZQQwWbKAJt3Esn5P7S77Y3VR23
rG8RNEBNlBufVScVDLTn3Qw7luukcKpl1MZM2ZoGLcLydUVRS5uU7jYzDjiw10SB
z4ZursesAua2YxOzvJS3MZB7OunI0JuDoqExSIZErX13Fzbhcw57VAvSH5+/D0Zb
QZQwNgXJahikqCsTCA4G6oZ3hI4EbGtYesrGV2N1ubdb4u43ETcXddZ/TelXghMH
nLfRooIHJApVGgIiZSnKSZxPqyE10RPzhW1IZ0b5lGM+XHXpw6x9SJKHAhjhMPqH
CKzQSdUX/KA2xbk5cAmKuimfNG2HeezYG0D3nddiVAja7Y12O+RAi284nNRRQM8I
WePQ1qsELZuIdwl6oxKWacIaoNLFqZw74Mo7Z4Wq1tPxZO4xOsaJ/y7sPZSLMd+U
CN2mrGI4FiIGAz/qTf2uBTyWutoggebwSSgGUWU+qhiFrIGPoOYIZGBLjPYMvliA
yI8VXb/1EXPM/jzu/MLmFTBEElTSP2+52t78fqiaQKJN31ygBLN55jk3l+TpVKyr
2xJtExq88wwFu3KgOUkRIKT+7albzQD6YHBlMSGhUHdOnICH2m9/T/E0Z3UHivHd
hOQ8GAfiSo1Xezi/PX2Kyp8ziVjl8OGYezFVVvVPNRDAUoCnWW2pu46cY2CZ6xOx
+sICVeBoH4srhoM46dwnqtEMBdD5vnXYO9rFnSj0EMQRT66NWux9bCRzldmtDLEJ
bxDllJo0sZBCeVtFU3LJhE3qGcswnWdBxzxySsziBq09rG7Bw+Zi7zs3TJ5WpibP
nw2UE0ol15kHyRTkOouEyX06mbdeTs5aiBAU8Lzmpolqh5eq4OXfDVt5tXZ+AbkI
gtEE14Un8Udus+kVUzb+cEgNPvV+aQ3sq+FJ9p6UvMZSnQff8F1EKomvFfnAAgBm
rCghsiiLYWRh3MkWo6IgWdX+J3bpgL66Jzj4MvyR+Ob9swKZ1cPtXGYf5YjjAM2E
ak9L3x0Vgin59UF4VcOr8RhlOMTBRTPzLzNY+16smP5MFvBHe09aIyCu2uI9A3tH
mFl+RNNql6lkCF/UGvBzreVH4h0BonRJSbriH2V/9AFLf1unu93SmgQgZc3Tbh47
Uu4AH8tZvVhGr6SHx9yiPC3673c2bS2cwSx7A00im0GeI3ZK7tE7nAHt//IGYlUp
G7Hqd1JCvXlWaqgHER/m28OeR+GVPFgMfqrjLUCkThha7/WLtu0ZaBZMfwnwlnS/
MnvWIYYtgQJtx5Zv+3LsTleR3VDJEJsSmZFGAz5fecKDuKia+c4eTl7S03MUBHYs
nyJ/9+vSuj0m8s663gg+vxdfnV1vej4q6BDoce2VL5HIKvaluK+TPrBZol8EJIXS
O+u+8+XTAnH1VhLTeMU6oWeO9lash8fKOK+CdlLhePu7vKvIUIhPVm9VXqDcXAoL
rBszvCahKwB2Z4O9QQz1nmMt1DZXw5WoB6o0m2jMYgU0fKDCUsjqssIECcyyOLHl
idQycWisKgYvvikpWr3s4/nts5qKCELCATMxmAqRVr8HYmw/rYO7tgNKGEyvuOO4
yk31cuSvPpJ5hVUsm9LZkrE83sYaYeEhHb9b7n1l05kQQTq6AAIqLreiDtsxY7C5
RvdhLqG0tG5kJYl1hK16nJMys3SAC4BH1IylhTwyWFiEvMkUyPJeswKj9+fUIfAF
znRqrCCod9JUPENARxLUW5r/mXLCJ8RZ3WD8roCXSCAU3SCz4TLTnMLxBnHHrrmx
YyHWv+CZ3DId05Bp+ohXQJDtzRb7jnVRvOD1wDiBldb9e2SVzSfah6jASrA3sG3f
x0IlrXJshDbauJlZHlYOhbcSqL3j7rWzXG1LIBfzcAx3V3mrGXiEvle8g9VE2u9B
2cAcS5mOsP0u/nFL57fAaz4gmRbdNGoCwpAe982jpy5m2dgvr0n22DLq6yMve1te
WwsRdmfFqIBYPiV35pFlSeheamJJ25YrZ5uuKG4NzntBdWlZ2KBZ3spm2tKJH+SK
9i+oDbDOvXT433rTTukCrpzT6EbZTCDDIWO1jT+6ciTP9avuS0H1LkPvRvq/FmSh
iBWHce1fXsYHpPYIhSY94juUYY8gblYWrZdXKgc6DmK9pzzuOeWr4RH72G6WTSIg
nXkhEWRC4Sqb2upCZfJLCAn/uEtuKStVJP00gSZ99z0oIiYA1nJWHSBTUbe+pNIy
jVwsy16KUbZ0i3b1aQjM4Jiz+5ywDFAlqYw436wbRNuq3lY+UOxHs9QW1sZq3Ha9
VKRdbk4noIIcb2azKlO5kCPr2n+qkNADZasJOHRjfPX4LpEHH4ymVsW6ZXtGuCCk
1almLaX1v8nR03WCvjWHH+Yt49Mc21nkw1fxwvHizQwfGIJ39qiSLfzZ0fQcSpkM
QA2h/m5EpZe/DIZXiJ8/KqMmaB+31g+lqY8kZKacUDHuhumgOg3yBWgEMnYAWD3/
FXHcO3A1ZUMWFuA69qXr3NuklG3fWB+lgGjpb7BgvUV+/TXp7AnKu8DVuRXgb/Br
PO/+yMXiwC+Xy/rzFFNTb2WAshHqq9Jrc0kfg37JF2d9p0De3gr/oGm5MbfvmsSh
+ZRGmC7ar8AiCWQOJyv+nWXz9HyjdQt+c/SZiKozjN1JqT7Nnr9Y6j/S0SdH865I
9Af0kjSEh3EO2UFtYCSOdj85HHDbV0v+ZYEFSANiYcrTJ2G5ke3kWFJVGwXBInTk
vehG4vwn1krTAS0CPKgao9frqtjHc9V+SsFWF6HDWNtHecSliRKiEuXUsSw63V6w
ZLxldiJdRwxzCOKIeukbFUTYSbv1Gj8k/crqymb2VrhZRBUN7o0UdItb1RLkHsvp
ZKdxqeJcmVjjx9cYt7/Am0sUedqgdYglf7sl8/x8ziqsGgH1aJNpBB3mF6V2BJv5
SlN93oThOCAyopyJFjaIw7o9svdIZ84UARfMMkXDLhbRlBELdam21Tt1+2o3ncJP
8+fWH2S3UuXFI73zN488EQh6B/G30X/yXWqoZHk01hX7b4QsX6pT8NFS81rG9AxP
qoA1jfc30c+g31rjQIweBjTTmqFOu3CXyXojxdlRzoOEzkQDFKXJ/6qxsgLBIObJ
BDvj3KCHfx/MYIXxD3nGbMgzAC3E7fbE82CUnZCPxjOJw9gVx9n8rIX/GTLJxzc4
IdhYRXNi1Fu7+hqHYwlNHys0PqLT9h3rOWK0bwUSi3wl53yS/4pFChVlM6QOwIQC
1KBq6mDXxh2jHnCqP4O/e1jK42NaRcEMOXRQGL8BQmzBlGFwFAietGb/LIOw+xYx
UMQ2FY+3AlB9z4hsj1onDnGx344OnCnxo515rcFQHYNffuvqnenqIGXRIPjp9YS0
3LKogh0mRoqD4ZlNZUC6cH8QAVmBrjIk3jYCbE3ktAL+wX538XpW5FJf+W6n8G/7
8phW0YE/lPvqZDfL8V4INw17BJwpzTJrO1BAqTDpHNszAnuMevFGWNXWnDxP368d
X3kFa18jFhUttMaJ+BbTYl+WenZOhjHFG93OPoIULXxccn/NlMbWfHS6c6A7TN7t
tHOAAVKrTeOEAdDRSn8tbz8QfYvn3NFgy52ByGgeD+e5BXEIGESnMa6JZb3sloHk
0saMQiFkRTFpFnEcykWMxO1aIyqCeDZpu/SRgg8dhLXIElJ/m5GZkd77lbZ6hbYo
hCyPCjT3YIZ4AYyo5kIA1vk7grikBAsQqx2FeDLguNXFN+Vr4JFIV0hZeYm3g2M9
OIrq70B/jHm458urOhDnHp/vFZNli3WfVU9Vn0hSNREtAevgGmlDC2aSshw5gETb
trnrLJKE7QUisLIXYGoglb1+O/oqfQTMbFyVo+ehJRQYtVdi6e6+ennK4CKSu5Y1
QiQc2ExNKsdmRXrK2PjfnqeJoxvNPOkTiuYo9Y3xxtbUOv16CvhVC5aV3qMwObNb
yqxzLMh3iDAqsVYXaEwMxCsMWrvDqmXyf2x5W2x0r/n9EM6RIjjIcqhzEdJSsxwH
k2qRSiwwGfFu60OxAiqiV/xoFlrbRG8rwPOI0Ng92RpkF9A8LDMURzr8kdepkNBu
eNzXTyT6UA4C6Ms4vfLJn333BbKDAlCX4b/5iBCtrQjg45muencU45rR15f1e2m1
JvyRp32kN4jRW2AakgAX+y15zUxBXY1OctAtIvX5Ae+WIE/5whH9kig24Wwbz1hC
PSwL/DTdlcNK7HYSVTuBegV6eFDxwIMc0uSu3vVOgAa342aX3RKW8eyY6xIJLjx+
ptcBz4n3jvwK+NYnSeS/v9F4O6Pjn2k4CwAE0yoUWEyGiJsFkR0BBaZcxo+wQ3GP
3vQ0giDrZBJxZ1JKSHsTogAoHBIpZ/vCHkghXziIo2dp7ftbT2atoBuKccWcWxM9
UyjGzw7Mh0Twhbgm7Je8abxvvB17y1WSueC9PdlTKQ7XapG1O/j5wswI4XwocTxG
FgeEC8aGnX06dvBZEHaSm2dDAE7iON91p0gS0QB4ZSoyJ8pXqItNprsw0gvvqnxu
GxlCuNwWevCuzkC0SktdZekp45KM2GFdNCnYRZiG+6y0ZBdf+OXrzLdakW73meoT
ikKQWchLrYjXs8b7bluk4Jtq1z+nqq8DM+/SGQW1WfK+HimYxyEH+bnvysFxARNf
z2xRlty1YCxggc4rmTr9nC27FnqChuFF7OeeOB69/9XQTrVYmDdbaaKKi4KuWTGp
1Z4WGyx7rbRFJXwKUwlDYt8kzaZOnKRVieTwalwnmDiOFrKJI3xOkOWVyuIYHJO1
2iadAHuSGPuNGMN9PvbZnOOjKKSPVSxKbulONvvGISlYYhd/5iVQjUCQOD1sDJhS
Bff3TfKSChXZvdxcudHRDhjH1QrT4GuF0welH+QbEkYbQyqHxWMwyobNXZN6SbXB
HDQled6vaUqCfjR1z1iGVxbLU2EavLSOStPEIqn9Dhl8+EK6i9x4i1n0geARL0NP
8XBMIJl4uj7JRIPNBVRvDGRUMfO+QOEEbchhUCnlKKYv31NaXW8QHqPKkN6VRfrQ
aGtPuSIWCcgPg7OlMC1cgvaxRB7nfAUOtfcZ804i+5OGmUvKRdrke7AopcUzVMEj
Vi+fcTivaRJQ/iJ2v/RzdqBKCkQbtcUFiEmZg5a0zH+Grj38pJXOw4oinia6fF7N
W5yCXZqG+F40OK4khlM0Me0nlctkJge5ypLhqlMD99Qqo1KV/UTOTGpaOKGmWS0A
2UPufNCoRlKqIkyx/C3U0d6zQP9hvk78di8TclxLmffZvBpzFullhNT2BczVvfqd
kccbPjv+KON0JIf57NEACdxvTCFCxVxoAdSc72pYNcpgmhk0ZRGUEIXbfwpyliVj
FcewWYtAYZWy26qh7hnC+IbHOvXPveP0soRORWveRC8ztuqWdsQzmtmjX60UbDRk
EWOa+Fbc1l3ese43TTCRPYpz0sJMutQhNx2gSGT5F2bE0FOM3KrYojA6htothn5n
o8Hygn+a8GBK4O3T7hURqgSrnSaYMObtQrPRYcBF2G2pPgJ9Em2uCw0OJ01I47qf
kqOFwYI7+eRJm1OUwG6jTfDOYF45b1AMtfh3zxasURkJfzjsK5RIbBetTZSeonZU
AgpBWaSqzxq6oLj1Hwsidesign2xf2+yrYDBkMhhARZVKZd0gkpP/lvKc8Y43GuP
QNBu3AS7mHj3FkLK2q8+a1A1zowtYvm4S9AA+Vqr/hCIA27PDhs6kdKE709PaDE1
y/gGnrQCIoWadcJP1xH40DahPTJgTRG8l9d8Zbf7wZUAwT+hQzGNBkOJCcDsdikT
5pfNqffjBkPszVFJTxej5eBPrl08DCVuPOtLllMr3nnuwTfb4mzJvhgY2w4kmCtK
VDcCRallQBhWBhPAppP3r+Ze84DeM2uxjanZ3S2QIIPfvCCAHz5yTMjBexP07Qpu
2IW+kIyq9RX+5NxcOma85i/lhvgSNRag1HUAKSM3dXH6uCIPYzGkuFGQwJV76rpx
OdBVgCxz3uUIIdLyezQQo/FreCYtf68milmldmwZsCcdwmC5XVu0jaliGBfDSUBz
x/4vfY38pJlpEFS3njjtX/6XxHpMhSoAjlijwPKOAZYA1DMWxTta5kKlMPSvvYg2
UIEtAFoIAZeBQZFKNH+WTDkRf8Ass2U7cHxbV223zwq82CF6YbqZt9armqlkF9v8
7kMLTrqYat9x41VQcgrE6Y70375UZr2JjtavoPhfXP7SvYXN8ZdtdJmOJWu71RSt
WuQsM5qjNgPzmYFH2BTa8mEH3WuOz86/hhjWeNNWXp3Vw/kMv8NIfN5RImTUXx/z
H0J6GBLGya4A7wlF826BV1HZqLFHU5t4mJue1DvmZLYog5nWwB901PdkYtylg4Hj
NPFZHeOS5g9GLW5msFjYZGJf2MdHTGskLsyvVkupMxzjPCsB4iBj7cvVDbaBxpOA
vLSc3qKIk1Q2MNrXePcuMqzxGt2W/JE3Y+iuI4KmKuTvZ4UF9HvEfge884TfY3xf
6BKB+QkFL2LcO4d0uzmA+G0hk6kcCVEC6BckxpGZ5sEpQdiSUaOOFHUv6abYe502
DlsmbZ9RDpln8CoVIAgxzW+hJrtlBn1YbJIFxMMRHsT1IS1uashAer/8U/U0x9tO
OyaQq8pcWy8QEW+226NQE3m2nanftDKLv1V5zY4ZCDKEpjn/CJ3vCq34DwvAYwRG
KEMwdyW/SP/HpFWDO1ZL7DFZQNSdtWuPJYAl+8UHUnzh0n8W6YPKl9uqFIejPAg7
7hqi/c6r3ExW4EJ8lxRc6hEOIN9rUxy8ggwqrN0oC73V1h1whH6aHT/juumOLB6Q
7EnxSOGlOz9TD/ITVWx0EsIiFjt6Q5IWpAq1jP47ukJqgifC3US2+U6pTf78c/XY
Y2V3l/VwjR2YAJoKSNqnmuJmdCU9JF4aJgWY0IrcGllaAHEzT/bMPt9gnZujOTsL
3qdQskPDk4qkI6RT8hM1LvbzgTomwYyXTzMIJX0xuJkGjp1k0+Hsh8B3Zs8b0Dk4
mjGnj528rNYCR+BzE7ZOGTyp0lFrx6GNNTZOXpzb/xX/btnK/VFdIp3+BNrugE2p
cYgVvVT2/4NvTMQAi3alYo8Ev+XMQPYbyjntHcTAlsrT18xMdZD4hKxniszJrYGb
c6TdOcjSSZNsQdjoIdOghhbnt+0BlC73D55vLOxTvPfmIccwNHD0B0JAC+CGLKre
ERAYxI1HtHF6/3pSDgESlpObkOg719tGCep2rvrcxcSt2R1mca0mTD9kAfbwIIph
OcKHe0MKwO2j6BlBVbREyrcOThUcc8zLmIpoS1xpo0+8LwhLys0/wzr+GOaq5Cbu
SHRD0um81DawOKO886+8ax7bcV17xLkIYA00yCkKLLT7nWIzkkyvGxBl+mouvb/8
K3umokzEcNWfGMHJYVlX9NDHTbXtjP31pko4ayJ3xTQ7K2Da2nTbSjnayTSuJntZ
YaQfP8Hynx1sNozD4y/5OurcICCaLR1zFXZJUJOGSXjl7UZxUkU3bX0k++IPN3VG
Vs0uUAWhUJ7A0tM3uwS2tVQop1i4t33Izbcg3LXFTuABGkEScUUBe8EzzqWykBXM
Ng46AljthIHk38XUtHBC0hrrjz8eDX8cEqoYJ1T6N5xANWgrqP7XB3hNVlY0z4e+
qdByuFX9NlB70iUz7pUWZ0dD7i3X4GtBDlMYbYS17XUEqzAOeLZmEFMQxy7WZaV5
Dbm+JTvlbVCho4QUxUyzNmSriqgJ6L360cyuwITvII2BaRHl+IfbvhwJ1HZOdkgp
pdYjOXEM/NzvdS4nMinQePyHvj5eSh54J5gq0ZuOn3sDzlOwX8Chu9rKuRJsrwvH
WnLxJeBIPd5nMR8tAp3dZex0BlW/bhaCjcOx3Fuv4x0oDykHJ0ElnTIayoTNX5dF
iyjoY7XXh4pLR/UwplyNBYwWkoiET3tOvA7wHxQcysdmlGNZ+mTm0qmJ1awPrYzr
6nYUgis9e0GoTvlCTw63nX3Z3a7C/46dwOSYTnHuSVAcenZcFj29YDLzluctU1i0
OpQ+dHW0NycwzvpH5PyA1AIlgkgw8kQUi+l456y590EkpTLOkYZ+AaKNq6z4duOe
j+O0zt5+6AiUxNooSqOC/ND7MCQSvRhWYkjv7v/8AzE8ZhFzko3qNeMsjDwWPKMo
mJqPzt8aDZTvcm5W2gwAingvH2nFyL2a2ZoMD373bFiP22HnvSJSBCLUY4Cp0RuW
6WeZ/LQo/orErFiYtI1zdbcs9ZoA2S00UeM1Xw+syX0qCd01SYsFJx9UbPcbnVxT
88O0c62tHCa+hJIndsVZcMSHQatfbvq/pdoA8Kdm25PAXqs1wog5b8n1T4M8okQL
HJDPdiCFmraO9cW13CjQarqQVawtPGrDnY1wWGA+uhJ9Fx5CbZd7GrGAM2Y6aMpO
CLuq8GKGm+jZYwmjUljdOvnnfGGXAarrLjKaa0n9cBr8EEk67jFPXTTrfZzGR6LM
VgxMo49O6j/iCmVScjkkkxw8DZnkehU4SbgvSbmz2vboi0bMRFzeV9NUA8LL1aCt
cONjMz1FS9U2Dvrsaq30OTtkUOcT1PYTr2CCVYTNlmb7B4p5ajAq98pFrVe3O5fs
W52yL8VlNow4LbZ5SodCGpUl0/uoU0b6EUhvkT7m4qEQ16NYsjaD3zRHi0t/ohRg
cgkr9YHTHKjgbXYoeVzi18o/gG3RmUHoN5buUO3Go7JQ7bIO/Jzkv70KK0k69PjY
JMnWzGhIAZXRMOtgWJfu1Q90G4qKGuIYFTUZhAVDKRWeaefphLzwu+CzpiOIbhqj
8LsRNw0lyTCaR23RgasXZ9aCu/xnyGCSqCPIWfJdXB5BhHt+C1SzC0tCKrXYOX1C
NNkF5hPdz0++8e+rO1rsKGDgYBTTZvs0aCMOTUP2nF2QJde23SU7/SdpoCGN6iZ3
WNF1RQvli62DjSDS+R2mKuvq0jniTxjTAL287HZ9m9BL0JRSlUgGwLYRoRX961Tn
QjPKstc1SAUsmtMmePBkpr21JTmHgXhoGLBr0QD+IaJ681Y6p1FE0kVS+bBdRhdv
uIxjcUzWj5uAIfiCw6iYrn8uJ1oh4RuNgiZs9JjXUb7tSset9/4Lv8TC7QbqMPUB
DZnGvqB2RvgZ1cpDTOmcDkTE47ECZP5FoTizXfOJnpfUjduVUMro4PLQ/4IcB54V
8cDyvWdUGHY851lxM7s4LMhu/zLcZrj9yNLc/XLKobAANkc3giHyuPj0euH96IJ3
3x6rLnIK5wHHExEOr/28OQ809KYKOnE0wipvZ7H7fVsdK5QxeUXZ+sQRZ+FU+QbX
7EibxsQNi/vEJjOjutFhi0+AQo2ueb9eaFpvqoPkJlYyB6AWKCRflvFIDBN6kA/y
zZShDitYefoAHsYcpu4B7FNlmbE/weyck0njWBK7/Wn6UrrnY3wUmmyb788C3xDz
1Ql+KnjWDR5dTi4jIRu0uRE7kx6uFWpHR3Laaq4V+rG8/OW0+fHcpuWPsQrM3Dug
AdCpcpN8tQcPMR+BkE9dL5k03BaXlPE3siLiTuydBjQsakedClvUb6FsIdK2dyJN
TcksDdk6gCjX+PpryfIXwF5WpTSL0iSYJD3ht4qjE9Nsc/q1tl/WJfdKGnjMzxmW
d+MtucSYzCy76lJ9kuNM7vRx/e4bf/JZyGH6xRcbcrzUxLWWCHny/z3LtmY1rl5g
pOfpUYvc6qyxBgjFLVDDGOF9+8uDHYfej9wJ5zOym0rdbscoPENI/81RLtEX+NQz
s42ql7n9hAM0AlzFqXzOwACULEh98Ye1Ss0PuroP3dde7LRGOWHNZ+1zhK7pXXTz
S0JDNyhl2H/2mv6zmetHmBUJzcbFYDtK0gBCLaQOdqM4+O3ddS3JyaLIiCX12oCD
k/wGyqG85138yxjUPRAi8wdzPwpnx4agWG8nnXOR603wfTVfrucJv1xeXJ4G6boY
7vhTkgYFzMCoQP7nMD9xnNL4fmOMepZd7aDExzJ5raqHuFJQMKf8X6pijkM8VZ6g
EINTpL+STcGZiH9+ZRI6Kw7B8iY1edgdCf0nrGZq1a75EOw4OSzrsaPfEe0CfCK+
K/1K27mmfJasWy0bUiXoZjxdn0xwNsCUItjIoRM8HYmrKI5dTIxm3fiZQ2ls60eX
nQyK64XuuSP1dAoMf0tSqwn84t994Y7/tSD0vnpJeqsTv/SrF+fvPgKswmehW4s2
nWRfY3Jf2wyKD0jGi2C1e7D/aamMrvVC673pOQ/IVlad02STkas2ZP0jsWsRP7se
mQnYRAZ/VeQWWnCYppREesF2JKNZEqMcMSwqK1yzpwqoFcN2Phq++yecIFeQG80d
W8DnabJo5eiOTxJ2mjCZJ6ntB2RMuFceNxPpv3EPVCMuR6y9dqZoO4dtjRksILRd
pb60kji5QilrA2RXdsVO3baP6VVLfIfgCxV+AfMC77D/vC5znMWquJ3U1+frfH7w
c915WBKUfjT6TBvgKSkLxtsFaU8z06o1C1TVUXkcFgqDVoX37bsGXrvWHVQ7Je5N
auhZ/Tu73QczMQQ9PE8lIReOuAwsBCHFw4azkPdb4NGxcWCD+akIGO3+BORTSOw1
NjuAnMSN7dQtkR4JhUx9aRXLBL7aRlSSLI7rjKV0fLLttqsdi+LkYa/G9JJseHTN
sIYtQe9foQx5nFiA//qiChN11JuOuoE7pkgVRJntwoJbetaSMPo8P78G+KgUCzOm
ADl1bZSHWgIxqgVcL8VBSbCIE77UJJnGScFOgeaJpxSLE/6WdV3vvCL7ph+grhad
DveTAVZ9ukuKnKTZeoky2EFPaOQ2FvaAzQqe2Mg4TFsfC+Vkj671NW5o0Rqvc0V+
am893mPNNfQIHV3fGdm+5RZvG8vM9ItCQNXSW0cXVOhQuJk0veOCk96szPvc4Q+u
XQp1scduCoT7vNUyWGNZr9+olxercclzOcQYHWK8Nrx0PFIRjqymwmmHHhBMaqw0
eFkxM9QdK5juHCOVkd0on7D+FnzYL91NjV7P3Jn3efzNqeBvnp77gzx41qUxFAmO
bRPeKvDRKCdTYtXb0yLk9LK1bLgIM7PvxsCbYyE5MDk4BgKvOFLyOH7V7Qq+T9uh
mx6BQFAe/Ps2Qw3CYMh8lHO7YM0i8bkep30cln3s6n2am2YjifqX9m49QE631Cpa
BphAfrQn2HdGdE9Uw6qZagH3EmGoXs20BnLoSVksFJ0VSIIQ80LDmILVMn7lGY3c
nMXRKoJjbfBt7vZzYEtt9CJ1yir5KPM13x2BMTLK7ifeP6JhCGwWLEKLrKdcmv1D
sUhUC1SsmY7UIRqJj2beGZS1WsEnVdp4tDTcQocsCdTxWytfvfFK71qwcxR6nd+j
U3BR1REVvKnc1yo8OHgoWKYa/yB3KqIE6HFdlvaiHtN4/bBYsz900UPRrXLiDo1m
lroVk9Wo9jVr/R9V3UjsZdxXzAq+3VsnpEHYymv9NWc+7PM6cm42XqUdmfEUWWlo
3d2KQJ21Nz3Njgp3zLbq/vo+Sk6cFVOJKXTIeCsQNsDvLN2qs2GOB7xjE0qTjZot
X2ISo4Gubtr+74Ta8/hfBFUs+sHgVjyPYDi0N9N34wPMB7dcfx4hU5j83GJISkel
jKkgk54KkMFAHe7l6fhB/lPGp4JymuRZj8GHuH2Ymle5A75dbwk7PFnEUW8oQPQU
W39yjHSPOa7m1uPZb2MNDCuIHWa1wCtfLxCH2RfqqniDe2SLTaOySMqLZCOF4WoX
si5B6L4tBMHm70ZQquAHuT6Agdf86c1KS/zbEwlQeIsmbaDxqmhcJRJ6fmh1kwB2
tZjcwngmy2TwrKSyrKYdGpMnAQnsFrzYAzdDSrQs/ejj53XpHqD1W7xdJK5aNw1y
Fo5u02mbhN+79ykeimJJ4HCe2iQyODzJi8eoks5jPXxMPklBZIC/X2pPfEEh1hcm
MmQthiveWZ1i6ikLi3Z/tBr9JXkqEJVamnDjIWDoy0VzY5QsLskx56GGpFSw4gbw
qB+ZU9kpiQ1sc0Y0Ffbzp9QskBdyKFRQsXUbVpEWSVC+IqI4NjzOpGK+2daIlq0H
+sEYqpIksKgHzG2qEmE6hrkKcboOhiFpJ/n+UDJo+PKGkWEyKQgnWrijGhoMW7a6
6l8sQ+QpBDyW+iWa8sLHDOmny8wgDZsUH6i1AXeWe94XFcuYVi4s1M/vZKDcPPjI
CpEiHEgHrWj1uaGPkXbF+p9F7vPnIDalM8kCXpY0frpWpCrJBY0OVE0J2rm481ut
OiDdofd16h6NZr5QizuAA3Du44uRPHLTXuIwbJyj2M+sw/gv+8ejzYXCFfYgMjK5
GxEuVk7Lxp2IRAn4tZLXZOKgNETYuOwJiHOpY3k9LELCXi6HZte/zSTmk9HT+ddt
4ws9Io9m50wzWszUVPd5xKKBFVFlRnASeUCnDl/rCd6G9DAVs1rTMXw2bJ0xXXDB
CxZHcrNJ4DineyF3mX0qJu2gvRcj9X42Ber1KRjFUmXfodF9WW2y40Ax254PN+Xc
ERl9rMBHMC0Iypj+cjKO9Y/kydA4hwySlveoIAq9uE6wNoeRtri0h/1BBiLpkxnN
6gYApMFdySO9f8zjA6LoP2EaAQR1d91f9Csi0cXph+cPfO+Bo7O8Z7xo29zLGIqR
L5pJAo4VhWF8d4rEjzsyE8te2nvARX2eCCySh8ouCxmAh51eLA+wQZUmMCs1wUO+
BE5Df8F4dxxaelcuUL/J2BKZG4ijQl48J0ZDNfoljTuvhUP879Vqd+j1jJ0xEaPF
7F0l8+iQorczrq2kre9jAKWWl7sh95FYqNqvgUHLtiB/MT/cpgmur8qKhRpf7Vn7
Q3RerFGQ13wnxnoq+f90VMKG0fekpbPin9e50OouJMGXIShPy04kJlOmCupmDPJd
44kYn3D46Y7fMxnThdkvHT4UCEfQPUYDD/UUnvi4E1sNYNRcZwdJHUHGfp/iwxN9
Iod/pkbLQlGAE9WqTv29KRjy64fgZbjcRDmBuRHfw2t7apGe4KeKbXDSZDHR03+P
S1Xd84LF9GBh1Zc9hctNRL0y9A6MQHFJo4bmZfLAOD79Gd67fZxEHF+LHw5JZYgW
28GHbmZvXKCc3klGeTra/NEyqhB//qT8U8LyneCtZO5fMoyOD/8gIsIXTXCxlfjT
FPW4ujM3CJT5nqQ4xsGzqZwIvQ99jSPYzBDXrEPmrtMIUsFXu9cmdMmic1EKpwld
/Gq0Ak4WM0YlpswMNh6Z/zCuePNd4hQCliVu7b4v7RL8id6Q33Mwwc45BBmjXp7n
wiugY+I0v+1foM7HZWyXbqBVsCTO/Gi+RFra65iRQZOhjeyJekmr1iz3TbpudR3W
9m3ddtedH7SaCUfBRUgMClCS4ZRyiLyyfwKpmAakrc+alrNDJN0azSeHCB8mHSvj
Au1RSRHHlglg3czpQ3i0bZ7hm4HCQQrFzXot3Y7Oz9AiYBCWYaXYtT1dyCyv7wiC
J0hGiBz7YzwZvz0g/rgjMrj+qu3IiJJ4F2JTfCfs2LKAUyiJUvN/dBk0B8hYw5xy
bDXb4BKlhW2ulBDcNf002+atM2D7xqFdTjLG+bK7xKsSkBAa9NSdPCx/04nQDrTg
KvZxS0vQrHJZmEeNWpV/INIQzgtvd/u4v/MawFhz30AXGWrDEmFSsQF6IgcYcZMU
gc5PzyzB85FKU8wcvCyBMrfD2xWVpTohXBrubw8DRqFuck8geOG6ie9EA8Nw2fC9
TFFCxe0LV2oQNxGgKemYlGeCnUfLwW2lvLvgXMjQA0LcOXt3qg6S/rKfkbslIAtz
8LW6PaB5xeMz5foL33bt697oQxPpkF0OAamcZ1WSbtO+LGNfUcjqjs8hP27a9qg1
7eqLkHU04SOrYBLjFHFN2XaGneF4KQaqEGcvRUfcZtN0e3IZaO5/twr2qJRk3JiZ
qoCYAU71tG4cLkeDR2R66joFFpU25AWTHEaWcKQa7HrDU5EKGv/Po99WFmrYPEGf
m/Sldlx9EVPVjOmVFrIKDc1aM1mcFu2ZGdugPWnr+mHnH7BqqfiKwDIRH2badPTK
DkdHYRrlMTg/Y+ajSnYhbisj3EIOdFlocWwpmL0QapkLrDlIw7yZKv2o7/LCOcVj
jNXAiNw79OYdYTV+7s6N284dGKQVtfFexwLw9ffoCqBsLrJypF/nzp7J2QcU2EUe
T47BsK3iAu3Osnfb0cN87AtamziOoI3QWwJpJ/4LbWVzzohThkVWBIzwhCn9pOiS
cPK29nsZrlqm6wv5SCvDC6l4EBrTIrs8wqxwF62xPM71HvvyijP1Q5nIzLw2bcWl
Hgy/seX4jO3J/00xBgddYGrXX/EY0NlDexws9QO0dQjR0ezZ3X8Upy2E5Boc1GU7
ElEdxBRCgulCtmotGkwodE30nzR2/fUr0vvT6h+NUZzoKbbwTa/UVHBE4j0Hh8mO
5WxKJleeas/C0rZIbzYiyJcXdAfrxuDGxw4yUlSEtnVp3oBkUvd6ekSz1TbPnHHr
7U8PMpsoDH+FDAXOziRDKLZQRGGs0J6NHptptCY1rpQuM+peT5pIWF8vJ4inSGxz
wObzr1XHz0ERlswwz+wWsUO6VFJmI9XI+9q37w+97LqUWMLEtFNc18DGqsYYMGeS
GxCb1wyVq2JDBrceRjAHo74fbuLHN24mHsAoo8TT+yTx1JHRHYE3Wntih+RHaFAa
G2yOUJeIr0M/up+R0UadceSEe47PYMWIK2txzacSwPujoO/xmSmIEEK2sZd1pLJD
qSSXAl+ZU20nUImycJQqUEj1+HB9wgNrpMuij4rxCGZ7FzxfAO3yerXBcYW+NnYd
qEAPuoNbGkNgtLeIYGMGXm02UT8XZXhae+P53MIY4IdQjZHMScHqRX6Iq5MJQzbK
eeWf7VhsNUEXPMy2SBi6lMDKl0Pz4mtqPSGJQRQTwT0IZ4MfSRPFdZeR2NtIvQtO
cbD6FgKFidgC57VxVJo78uWuwkfoDjhmg/6VodOjuBDW+lRLmXkefJwUzWTE8rzy
p6L+MvvTt16HlMTCCXlkfMNQxbk/EE96rYsvFDRMhkuQ0ikaWHxITHDL8BQcyGbg
Qjbx53qjPtw6LXZS9NAI1fSTj+hFmKfuK5t7BRDCBNHBAZAXkQyYtUycmRUsx9j6
X2UW/dRlUy0gECMlCpD3Ds0A4sI44e99f6kCaRgQ5P2/O55SHHyooxShrnRFZj/V
f0PE+Xe3H33OyIzMFna2VK3vFKy4oPkQdeXYeZIIoJnHdzs4ClPsLak/KUXIsfa+
74Tuyrqb+bp0H/gvzNBTqpF4Hlm8cT5vBZZlY24uV/ob3T8pD2f0h7fGFjGTGrTe
56PT38HRVisvywn+2nI6HopZJFE2ij0t0AbSUjGPqmjsfMulYlg1e9kkGmX3Pe2X
PQyUvhBRx65y76Uko7fO3fNBfE19KLHg06CqbbGm4iEA4FEZ9PQo9gP4LWwYFxnJ
PY/cuarPZ7AvNb3V8zJMFRz56NRNFOVJnn3HFEslOOCzOepzC/A1UJzZRuJq3ANy
Qv/lkdq9QjYuCFS09TtNhAvC3WyY68wm3vI2OlnTnmnDlFiJ/JxozMpkCR/bf9LL
0bCPmsI05wM44fNy3Mz+DG+3cdQmz1tByBjtXDSQn/HwhjcgSZgzgOwMD8dpNKCQ
Qn8HghTnj3JYR6VLBTcoYF/WJgQjD7rZOt9p6ia4fiZBrFiQGUI08o2eMj7Ivqsi
aLSe9OyvgNpcyF3+hbIcuDycRhGpoocxStiN93QZj6Byiz6cwqvSCLLzzmoVWc11
+MxxTRztCHetBeQFbZOcFa+W6HX06i4vVvzwZmIr8TrJv3qWWI3htsMhDMXHBkih
Lw8Qn2DgRTN6GAsXZYfvP/kGVW8Ha5I1Iw+3MfhhkUg0XnGfMuxkv4lyT2+0E7WC
E8NGXcHojbUlVtg/gXzeWJgeJ8uBGTyyJO9XH3n+EVs0BZewn8c/bYgJQlSaurqV
YVs04PnwYgTRtGKHJISBsaBbH9+v4WIs+mAtjMxYIaVWH1PF16TjWVSmkHhThb1S
aTH2jWyY6zn0DOfLzTK7a2BCyeOt2jJceOdjPM0M7kcE+excz554TQhEiDFdhuCs
5zwYnAaV/cw/Wa0Nx6MH93JPUyqNod64Bn5llVw+TmCGYV7s3mWbCxgXFuK9dvUY
PvGu+Yg8EcwwzAIWgRVvlTcwf+BrKAFhQa1S+fqCul4a0Zdp1k+yJkBdR6EEBBCU
ucBFO1K4Ua4CDSpS8DLn+26PLq2vNfVXLT9IXcCGOW2cvUylAnC5EHWwFwzHjnpQ
Wbty9it37plsiQG28TId+Gr+TMUO5y6taONKZE5yAtlla5NXUT281JKO6eIR7RvL
MCidisIQekwu/mZ0imw0VV1xYGRQZ/l3TdKiCZTn9r7D/EzyYNW6a2YadLeySiIk
LTyBm+Anhn5I2Bihr/1ccLRZE518ibr6OgazK/xChxtGWwzgbnj06Z/yIj38N1Z7
Hz4DuJ1xJcEiFOhIo6brbIEN2LTxoIKzU48JCEKRoWvWgpcdUNVto44IFxn3hd58
U4gqg8V9AyM3C+Pz4aDUQ2RwTyRiq5SmtUYwcrlQJuRIfn/vXM9+sZ1oKTBdmQzv
QuQxkUuFud/6RaNCxC3OGJrWi13xniu8IL/pSqFDN4le4Zk0Y1PvoARhSyTwBURC
IK7L3Uil9CUl+dxE7denWe0ALcjdCt5xz8C7e9s9Xn9fv5z+SoHIcxm+IQKWQvlh
8Vj6OgfUzo+77EBu5UhMevLJkaI9f1JvR4N2o5ED7czcagYiuxuZy1p/TUuApNx5
gvanxoS2hGcqglxd80y3b/cGgLTvv2vEOA7NhZFG/2hQZu8VaAkgZZOQh+0qhOGt
9VaSH/koTJHLyD2YF4Qm9IhGZBBmVissJJz+duTFoOddKLjjwvA/hdf6K2++y0Lv
0rR5G7InW4KoRLZ+MHSXXh7v8ccFUCjSR3vt0eradFPgCv8nHXi0sxjpkFw+qzby
wY/2xj7IMaOOLX5Qc/vmbqfz+b2TP5YqA6P/d+DOUBJWWVvs/mKh2plRDIsmDDMg
6KgSeyHnV2Cmp/cmBhwkY8//2qrRmptsx1jqGVVmIx6zj0FD1RQ1bkypx6ZpoCW1
yRRbrWpUqMOI5LR/yS+zKD6P0WCT3QnzPs8KTdyqabm5HRcpPte69F+WgKxyu3F+
eypRsRhDZxqiKQrxK2Gvik1bHakDhDReUpQQUPc1DF2G4oKyULFTHL/Yn6T3rsxg
RxkyQB7VURol+FRuQdoYARNs67qYfae0otOoOtqdzlO4CD1vBD5eC60c3DYWehW/
g3sjU9PX6VXb464iNWdcceTcr74tlJC3b6m4+pCtUfeE8xv/fVjCPdTKhjLeoPUs
Z/Ye+8CPPuO7LrSa+C58ZT9Zm3FgnSQcdivlvJTclGps1geIHGdbiD0Gj8jeoZNk
8SFbau78knXTMxFlv1jaZbyACrB57yiO9bBf09hhma40HGwpYCpOCwHyNSO9VQEc
hcWTcJ5gBLVIpZ6dw/MXR6JKAamv0iD+vqRGnnIEwiIHeSU1XN7IOWnKhHxuHeO0
BMr2AwtoGwb2NyQFvUaR1XVv+3DGg4q8t5FYXXY9Dp4rt9kz2TJ4pQEmX8a99Fu3
znPzWRA0QRkiIKbJfGYDrw48GuYqiFMQM1NdGaZRr1/CEu0g7il3iANJbgqidBIt
N7pBLfA7ZXZaW5YbNXgLqeX5LYXeuvlI00gVMLJgJWCZcqe4AZ5lYZaD1xcZW3PT
7GhcfGv5L2q0CoiQplYAQ5QHVUWKcxFFSviwXS8T6KspD+bgCVM5eoT+VEbXCXhY
IzVMO8naH5rjvpZ29A+1lRSFFyez2UXXNqXkkfO4klii/19LMiJySzkkc0xGDmne
W5DTcBnUnYh42PJKvUOh0PzBFVO8BWdAdVWM7t3VNDfA+ZJU5t88uy94o58FCj/K
d4JZL5E1g6fVENz8lGtBGBN9FA7fsyAP4qEHL6m51ZSoq2k1FDbKUXWLp3XXtG24
xdThcRzbV+LX5Tb2zRJyfrz5jgTAqNzIdug5RGnQI/Sq8GznEcr7bq8bH+A80H70
fz0ERcvENJb7fU6fsRt04g4nOMoy5iFJFZ5Vo3r8gpPZLXwIuYXSAYimdh3N1LVA
sra/m4EPMEZ6pvtsxQMZd9hpcMpkr6Pm7Q/9fYyHWFtZ4NO+K3nDvV1MhhUaxufD
6gwxoxLHjt/hb/JddjAQnnYlqDq0Rd0bdw067v4ql1l2L8LpEH7XL2uUEZOB0qFG
CVH2zb8phb4MqNJq6XRwMPsFy6Han+2Ox+H3znLxLz41kdH6V0tNs3V1UTu2tWHT
/yTcHhYyVqEzHsvMll+Tkb9Q+7oDqqlREK1PbLdR9Um1Fdk9b3BzNMiu+eQRgGP5
jGSmijA/Cjjq5SZnWqX/XqSGQbiEw6dwre4Qe0xsaY2dIoV35NRXXJivYUR5Nn3I
HrFr4+kXeAwtWTMfXY0edWFmdxOiIQPTkFlBe4KhtXyNR4q0F3L6/Lhs4sSoKDut
g1tdLm5wvoitmo+kdBiFOL5BuxVHTKuf7Df4DJputCB8gc1UKPlfbIMDBWLRYCLK
2Lo0nGOlNWAoPp74IO/r7X+yKvhjhgI4X2h9dQvpZ6TB91+TJFZ+VlgFASxc+Qww
RitQJ6Da4EL75RFwRDFr28keoXsjR5pq9zvkgci20uOwkf8TAv5w2K1MpxkLbYq9
9NMTgl7S0FLvpINlpMCdIXr0k0sRVz32uKDyMHljVjQ0QEjFw5PcaJXy+XXQFa8i
3B/YK3TZwGgvlerFbW5KXCWnjjzgMNZC8cAOLktqXo7rEszI+hJgqBXk27ogsAIj
SYDqBzi2ou+2ocjl1QiNMPgfVP61bfV9p+1Q00hsjJkvSSc938KAXMgCOcITLKMd
7Bp+LpyMPVYmRQrkYG0Sxf2sSwXwAXtuxaH1Zypjiaq64z9trL3W0J4wo5U70bR1
tKeQkk3/MTOUhWYgrNBJQzruZfngoz4MjUsOLeqaxVP7AdOAHBHgZMoVEEkATCPy
xf9FAds7ty3cu88ZsBysEtpaELbRNz3gX7YTrzaROSIKgqPeCylci17sDYxKX3g+
rPMSGr4weZZAX9BmeCI4bEFRHWlgfWgcfcAiwhkW55/TTPOg27R8F5IYmfsg4uXQ
ygSQYMMJk0syYp+YrRwHpOhb8Hi25pkEuCrSn3FFnt7X/cMxqF0wm1KMqPXBQEzH
Fo3Z0VxCAwlCCsZ3wst4e1oEVezMxWLkjVK/4+ICr85XNOikn9t/weDvN2CiB0wk
QTaTIgVh71acYs0KO/akAhkmDQwZYnEM0qKSA9mDCyyKeFJxeBLR0KN/NjRtF3Q0
St8G9O/sY5V/x7Lq7IwlWnRt4SHkl/xnGhbr3SJZylIj6jjlra8w7+kUPNLpvnHJ
hucJEBo34UsmWkyURVvrrE5GYVoQYVIGQJDqpMTpepCxEHSXyS8ljRU2BlnEQ+KL
jueB4OgptvJvcby0XGrbEFd6yThN9unL5cLY8dZ4hRbSNV04tArpfTjQyp1YOs3F
7a70U60FVwCNsDchcBoB1d52vttaZ5oy4XqQRAjFdf9E8qvjHHcLpcHmJpbcgZ/C
cJAk1dWqICt3cZwELvyBwScHY45WsAX+bXHaP2cuko0LsiCvXSwmrHfO4+GTySnG
B6E4+e4W6MSEEkaFV4OQqR7lD9RcVPL7UUqQ9/yzwl/tVxxkUTpqZZYmZr6FJOIW
lAkv3Z51ijr01LoDew2MoCTiL9BZisBL1OtiIbP5j7f0JRfTE0OOfwMiOJBNfm/a
YRxawYsJZLeN0lvkgAOA2kXJNAx39p7AxXfGtmIAUmWfuMnvmsc4IpKPSwlrw8d0
gdrqQrGdGVFH+Jbu/bQsVd8rcBnlxc5YXeJpuNVPYday3DsgE/RDOZebGYhkTJrd
Hf9mKrJWwlBjBpEYTjnQzefc6gVH0Pqkl199nNqriLgtNwgFQL1fZlk15rDEnat8
BXtMx1aZ0EoTn/FsQy5vn/FrGRcFTzAGPxjOHOk8HurvTogR2gy1KmwnVfimOTw+
ebJq6GdX11U6Itf6SN2cgVTLv/2gS8gw2uGjO9iSLwwl+/+cPysMn3LefJxg2ojk
iPhZhs3jFEoJkeg2nwVqHNQRiZQU04GB2FKAjXxk7sFeWr9D0nOBMXXZJo3lWhZj
KVF38xOBfH35fPU3ZsMGsJGmoaHdiAcdSzILBE/ziuHUVkpKUt16AFhzv61RVf6d
Po/os5ri81jWFvqeoH9jleBSSPTsB2kMIz8jc85KfjZCUElOeUevv0vKROpth4//
U1P6jdQ85jzOd7IQsthimjxA2V9Kh/n2dZ//OTfrLtztW9L1shIL3X8Ntiqc1pnF
WCS+XSMEeHzh484XH1y3lX7pz0WbBFIOmp/ifmrbl5FxMnm9S26s05elOOsSv7Ga
Ren+wIeo936ESHE47fjE5F9v+ifPokX5XzowZSQ6m7XpciLE9lqCe10EPXIDHf52
8pqcDLESgxzFjlypJt+KPER2TZj10mm4lHTmYBVrvv3h+9Qpq8D5bB6nRbY62YUF
WfI9lw6MPgTJxwEp+SGmruxixSEq2ODr9OakOIo9ZtNA30etVa7D6BYtMERVm26z
mJmb4ZCe+EwetjgE3SDFbsJyc57fYOYoaM0nFnk6dusakbAp0qiIVkX2Rz5mj1vu
d1eBOQNyZm1/Jd2FhSaMUUhFNOaUDjq7Pqj+VkZTyxPVA6fTfV1wZovAfOdpCPtu
Hx9+EU//CmBDkH7aHhL5JYB4U1yRXwy5H7fJCvTh+unXOrKhQ5+HSTYD0JSPo5Y6
L52hRYaQsuSTcWRD3gAK3sa3lJcc94H7AzpXU1fn6iTlw3hSTbJkTjn5dFY16h0n
d+V198Bool4SwtkD8r15vIgJRFI1kVHo0y+vC7eIbHUN6i5eS6HIrNpdjS/GdA5Y
rJkpQSbcqmj8kC06mNLAB0mrjW//C932qkNGLmomycvlId4jKsiMy0sGujHwJTi/
KCK7k8kOromAXymdDgeJs3x+Nz8noIaDaY4k7QwJMxWtURgrJVMlKXQamLoYeupv
9WnSf2ie23FNWFOHy8yfOtdie4K35D0JGDX2q3IPKqXJlfSzUSj6gF+M2OYJ+R5A
mc12l9HjmXh2NJK/Bja9Dw9k4o6i2t5ihXpM0OfztUhDDkLNpGclM7R/8lkKxUOC
37MI7RSka+juqS+ZO6Hdk7GL/JrtDmjZ7k8EkYyVZDUkbW9J/yMaMlWQHE2qWMCy
vSySfcF9bbJVFateIZA36P8UrClubsduKlNCtlSjC0zUrViy3uXWdg7e4/Pv2EXJ
22+VKgvDZHOSWeYds+T5Z8msKijm5ovGhsstThfkS3NDfPFWWJTnx+v6d3KuQePR
4zCLf90khika9FQobOYj6J6fhzrEU3Bk6gPiUfZzkfDt1RYKCwXm3CMI6Jcykyze
MD1lYz4sRmV6deOi7Z59FRPjjLoba+9/P5CwJYfXvb02La1AQNqypt4WGGy8lDZn
Ju8Qtm0R5yTUuxaWmep2cTf5wqhyq+oCQDSrdIcyoFb7fy+39um+8/ugOmOVyqlB
4WRm7t8u8ESXkOU2eswDSpM9McvdUJceM8Nb3Agi4u+c09Yo6u14MM+FajG7T30l
JtR6jvU1S4GGAbKk4dlEVndqhG4GFcSHbcZ1RxDd2b1X+J4eRmLopf1okG/Ndgf4
lO9OP6KcY1ETwrCJc7S5Abgq7/jig/K4R9xWCGeRyVrAK3lkWhcWLzuyurvb8C2v
xWmXP24W6AV2Mb64Sj5DTDKS0XkFbP2Ghk1vHn6ab+DfWl+DsKO9CBNqKTLNA0iZ
a3u23M1m3XHWzcLp2bWgkSg+gxIKZ1wWpij0BAJ1V6OH/0AZjnL4vpM+dI/I20gT
PSqK/qnN4QZAGmwJ5XqpnN6N2yYwrVOetlvDvisVA61WfEtMRNjVCjQJJEKAGOXn
EEGgi6wsmJ2LNAfuV6615Q2GNOTFZJ3Erkn47Wc2ENdyWrzJEJj1xneFqu+lUobS
r3jUBA4w437UZ5HVnzVm2ClB5UJ3WiiyknLfk1HEdoW4m1fgGti3/qiS9jE/h+bq
bN5LQaPFJR+v5apgbNYyn3+qxkS3HKwvy1wG07YtyOTnefd5RFGs12o1Q427n9Ib
k+pLwMqL4HxzQOhsNB4KM7Bcu9+72nlzN/ZUZJK/6ItuU9RPCna4D4C2KrACrloe
McNnUC7pfl5dAXZOfTVK7w53eQnABYOUJPpFkHt5VlFwEH8p7fG/z9sYEksz1wmP
6f2GV1Ob2bSGsW7k7M069E3J8TJSj8nmXzfDk//A8iGn+9P7s6+lNoeMSqJJRYPJ
G9v0CN7HbP/1VrOtcbZmcxbr9B1XjrjuExcvyOlUDOGacxFOSYwm9PD/LMLG3xc0
sjzgBXgb14+QwN6euacxdC6tS3DLiyiy7/jr+8YnpPQauA8FTeTw2AqeRBDiD0U1
aadrcgR3i0M9X/D3GKeIKTBURq5TPSGhfwaCyOC2E2OG/EWTFQvS3Qd+GLPE+c9e
21c3fiSYHTpzYR5tVu8VtpAZSQciWpZtmWS9FkkJnixnP/kc5DzI4IkOWdxQsdvc
YBfmwc0r4vWg4tnA2y4Tt+OQqNa2Ulcd5+qAHOa4btLrBwwcv2O6iJj7nPBsF+pe
6F9V/28MbjpvxG65NuKYA5Bjh1PK/kdRoBllNIUeZKjo8L+62pp1ac0h2zewPeSa
VJpMACFFLSds60qyoJgDvYs+Z//oCg8Rv5dNmgTvkGZIOtNpat+WBtxff+x1eAXY
tkoT7Abcop6gqCAwCnd3He8VYKXvUxtXgFIlnaYLuBI2eczaVZX4Fmr6uvqtTF2a
Xp/2kRXjAHzGRtU2EIYrFKUjgaE/X4orbbKsb4cueC9GVpAfj5XKy0hpbbay06pw
Kb0/vbSTXBCtACJLfkX1YQHpbbTKDJZTFNbCgRAPi4Hru0zBH3yLXZfGA4h0f2qh
XIZEsgKqF5HSq/jnwkOhmzg/T14At2NVqjazyRtDBTTUksdUyj72gwt5YN7GIZIk
7AayzGLPTXLWRKqRcNPoKpe2WgxkUPO6BGJTgoy9lnr09qKHWRYUrZZfGEMnYiAD
eH3S3Gx841oj7onfxrIXj/mSkCtt+WrqCCjq7NrESzK0hfTNlReiprRjYT3tEK5d
4eglzDIfoxmJ3OnD8mYan9UpoR/z2VmHRgELSNSqqczfajIywgZ8xiAA0K+/gFFp
QqjzqmciWcwhAulOj/2S+XBwGb3uaDAJkwp0HPgD8xA6ALs3zE15TwqVKghSmonG
W5febubG75KlZ88UcgsknvDVZ9mGprrJR2ifhSpfWn+gkp8yS7edo+xNeFfYWrV8
UHCS03v9AxwAkAINx2AzwuFwzJovDAL9UP2C61Df0yjXucIvyWskWhMtTDgFVY7b
YSQXPISdueLXvGGxVKu+r9Rog0W1bBQ/KxZbpwW62cBmD22YCZbCh5jgJW1GJIUU
rTHBcirwCHqdb5dYWhFx0ijhrAiqE/bLF2AWlEhirzkbEVwqDUtI8yGoEHJKajEK
rbZpHwDlxhNfh3vX+mDojaSJeMPOTejAKxukS8M0UQfR+9DqKlIlTZsehyIPzZKX
LP9I81U3DEsYQKviAFKS/kXBlgZoW68LpTAIfCOx9xjKciWfdgj2xg3JYMbIyp6M
g79eaqdCNwiSzhg/Pic4IelLND3Ku4UADNPpyyMSTAPdRIXqC3Q62ZWqjrxESWIz
/4giPiMF4WUvAbATQ5y6N6dlu3x20BgaKMEjKvyHXZ6kp6UTOVGouctv3TRSHFhW
jnhOjwwg6Ms1Vy9bA5U2+/tldIEoWLr9/ItmX/3uhmvb5DnJOYu4UKYhuPuoIfa1
/loA+2h8TK9j4v812a1+6N4JWz+e5qwBpJz1WPzL89KScDSWQTI8TGvCHTUNJifo
oftigC9xN5Gvx1a5ng/h21YsSc1EBOTBfrJbx0oWRQUzZFfokIZUmFjIE+lRsVy8
RUcf2UnjY06UA8IKQFP9kI2MKvChw9fYI1TJmwpGSPdEbc7I/FqSadF5qipo6rxL
hq+N5hLjzGc85WbBztk+h35obJkHPsQ9/zEC2r7ajjwABj4ALQbJtckV16+NpvfC
v+M2E7G6iqDVJ6K4mDtMoQGRVc9mm07gUPjPGEzyjoEMx4cOrleCjTsZt8VT4vOm
UzNSXg2ZKIPaKoqVuzrwChseGGgRwx0ZGoCC+KHiqkoeLH2ju5iMqzkkFkCMIIkK
Da6XyeBgzhduUtu4RMmygJzbBwFgixZ4jbFLZXbwXq+y90HqSo6U4dR2TtcCLiQ5
KyKUS6/QcNtj5AxM0iBE/uwFk+1FxDd1lsCQbqWJxouGRWH/ecPR5sLruHLxowj0
Uj8S5HbXgpeUP5R6H3usGdni5GfwaTd1SL3YfGWSKrk7oF8/3bXf9Nz8qRtH7qbD
mZIZcjTc059qJFaIsixMYNb+nOVlp8prHmwqOiUNxg6BlxKjJmsURp2vl5OcMOyI
1NfdRh9ajgqfcUK5oblRYuXIW9Z+kPRK4uatcWlB88WGIP9uhJwH1a+nn0J2h3B+
AtTOfKm649jlukVQPm9TUy3Izo9jtH3D4KeJGmrdlN6xj6zU418RqQ+oO/+HbzJN
5ejrOkIymunAoOM2x7EE7vzm3a7fS9c+j67qZrcq0xgUrS+e0bJ5riwr3L++JKzB
eA+xPhRLYnTQWXgtmxhESMptd5rdmeFJQWpT4sdgYNU7WaviX2Wd1l0CVH/d0hDu
cjw9nnDFO23UriH9/lbnP4rGQYoA81LF7MJVFlAVoBB/MJUFVrHcrIefiurbKiUz
1xrZVRuwjeDSKGNQe69v9d7797GAPt7/CPnvoqrKa4gYMP6pVT1IreRJRTGpj6xl
DZUxXlvIzi77LdbbZhc4qdmhHmZQzetBGrGDF7OpCnYiey5qVH5l0wbENXljbzil
iSn16IoYotZkomZPRn3tOTkbqWfet5kHrQpc+9XPbDRlfOvRsRQc8VvMMRzE7KGR
wQzBlsXH8Y4l1+0mFQukmSEk8NFwF+4n9wW7up7sAhGpW1l0Dd9TBIelbHfBRPlY
LA/vZBgtbMr/vosT7iXqMk7WnqF4rCfdXgYCtYMy+hgROkddrVJIdI5MytzDmdT4
IYlRzETaHkXW1/apPG/kzuBP9WZ/iiFaLQ35Ct/gs9idtChBbE5ClIQYpw5D6fsu
lPipJ4lYBge30jwZ1XEG2hHkLoTt1Qx6aYc6jsRf0+wpNgmxVUfq8Ug76jR/0dym
mp42OqYqbNqa8k860K0i0JPfedsgbPdzq1bhqcsJEU/TKE6qPUYO2VxLNNibVkHB
yCKidTX/wHN/7jaqiwsO/2wm0kN3Nsljy8i8HbTdb0HSbOziIJE+3K11GvUvw8Sc
QlaQQNpZPX3liO4uC+slBgroP21g+nP6NTUVkTnj7CwD14qj0RwFFrGUBielelvM
rdiZYaYF78pGTktMSCiCZkV+DcyVA2CRTAhXLMG+7TOCJknK+/pQm4lT6hsosHna
2eEf78+tTpOlhkgnSLxSdAFlRTq/Vequ31DdVQpeozYnFwIExbvOqDhWnpy8+cjT
H9Z0ZyvwyF+InD+tV1HfwQ2PKZ7T154bZYPxkuL6nQCqYjk5lswl0jpZ6Fpa9mhL
iEVWnEAL15ri6ctwhond7OXFWuuL19B95RW58623XvJJAkJadtmPv8oQUZWJTVS6
2ehap7cZHs6B7sQwt/I+tZkwAxbG3NDSn4rmNk/9I9BgBlLxPwvDCLfHn1pEsrL0
zRqO/VMDhQ3JxJ907LI54/NVPOGMTqDfmQ3NW++ymzP62MvXl64yi74uukRN20O1
I30ofyXwmaQWEdR2mkUBiWXDuKAZOU5v+Qb4kxPcx3meil57rG4Z0M43afknD9cq
pt5s18KO/mNBOlUgnsH7d5/FA7+Q8ZqJUIgc9Frw8cQrvl0LEFNjPo4q2n3ZnoCB
xW/XAO0y86FrI2jsFdEqx1QbUvs+cAkp+c+YRRRJnyv+/Hh7qOLO2CoBXTOgsHah
ch2pue0+ti/R217ErJBZmE2i5acq6jaID65js1sRiHXO0dZ/rD/p9nLSh2n+BR7i
y4Lp591AiJXwVjIpXeCnXiqZHGGXJ00bspJbrpqJzYkW5r0EqSj+n6wosD88BX3h
FIgj+ytfrcz6gUOf3EL90obpL5G7PaEWgFUNvnMpe4hEtSt3UkSyZyQIoT5UQYuV
oRRUJDG/vZhTDuaIIzhuWD7YsWzy1vkjAMec2uXHTSKGZnYrA71NJWJw5zlJN/yh
VLGd5IuwpRrPIb0TOP55CJd1/Bz7J44SeeA61P7cCERdLZ0X8fuayu6cAgpmJ3g9
896M1Mv98E980fBFW/Qe4txVpHNoieI0om/C4dG971MRxcqZSsz9w5SlRCCSkB1M
9o9BFpPQQbzjODhDDes8A6pmvVT/0yYAkq3U43GiTQPkuofPkqNTRpC9YGm2s6xh
Aezf5h9EMzNjE26P7rcrRNHg6iI5BXyOcwG6PtCvIsW2pDmlpbEuY90p9mtP+NTQ
c+qmugXnUgwOXa7FWvVROL5Wv70VLItKJflMktjebLQR3MTjN4qeW+D5wXecYgEh
P2Fu32Pt0kNWZsrN8Cw8jojz+mRbuIbP7DoakmxjKls06ic/n8S2U3PIXy8yexP2
vk0yxvfIsz5hp06gwgsAkPPE1HLrgm541SUqSGbSWrXvLwDtvUWVuZlNFTu4/wiQ
/3hg8zJgbOv2L35oDRLGKavn0eOmCJsJyiPHWcRuWtl8PpiHYI0S9yt/V8LnR7fD
RuJxOgO4tje5HGgtYOxG+qmnv/nwUW6mMp9lW6drp6J+jSSGbp7JlJWxXibP/vWg
xXf23KaIkDN+Pn9YCtLkX2BqzMAPoZ2pl7Uczh00lmUL2gyfzeDgu9VjKrT4WHEG
HLcizvnD/A81/awSuTpDJK3wji8hnj3ELVY5EMj/ufxNVRgFamqkqjm4AaEFX8Um
nTL9XiB4H4i1M5WH01Xpr//foT4sntZlJq4K9iBPm+3ObeSYsmyi7tqayZFMXIi5
Kh4gARTuFX7J53pDPnNx40LLJTGwGFvhitOoGwJj6W0fSwZVaCUHwTaaG6+NgphK
PDqtt5UunTIt4+tjbIkhN3KJEm0VMVfco/OgjpTiz9+CgVdcPLwJURO29+kMxkwd
WGian3nFnc5xcRYuP8rc3hEAswBpeX6D+aeLUxsG7rIdsTfbf2/3z++b2IcNEOFF
yPusAwBKQzGA8lXekv3sEEqLRVl2EM7IXI9E2gfepcsEIheJD/FI/bZ10Ij0GKxj
v31kDsjKHwIGMdXRHst/6WRj9yolwvgRzEyW1tQhhHe8Ip7KJSaNtnXDblQAcrKx
8a2v+AKwANTx/gEkgPvtJAsVaM60vxORXb3k8hl/6rcGkTTqioWni1B5RaZ8bFN2
083BOgtqj1Kc7e9cclY2/w5DttjXMVlw8fB2VWEdZbj9iuDiT4V61yCN6ozYSeKn
CaDY+ExeWZdTkKOthnBeYLB+UiVNoyLjOeIMm+pOjGFLvJ+EDO6VI/Gma2kImUgK
tM3O1puxfoBFvmnZc5fkTIW4CSXXYQM/U1fj2SI0uqdg9yP2v+QDBh/1vSf5JGQs
PrjPzvVumxZaSyFAsVsmhqKDJjYeVa9eChQAtxth7q0Ix1R2ZSQD4XZaorpU554/
qtl+LRE2w5wcev+ibLNsAbhXHrgfDqXjYG4kQTrBHv9pw1ZIxPef8nWpdVKP/tRw
W1S3H47YL8LHxkPdQA3VaQUr55Hnbt5OKGMntgeLTrJfHGaPcHKuF0nCvlplVy9C
Mr5jW+xVHZD9OMcnMcSM6uysu4svWByqtJqg/M538Gews/x/3I3jCueh5cM9582L
5eav5BYJhcdBoY0BonY8scjoRNnJvh9SLzmaaEMQjTeVuBKWXCnzvhFw6piYuLsJ
eoaAJInBLd3u2gDWxJ12fjQaCf+k4Pe8LmJCAV5iNCB5RE9MmmjHXsEbGvzkS1M4
silfWNTyuHpcMoX0e0L++Fnn8g+cQvnxpDfnSsz/JNNlpADcxWHbezHTf6524MMW
m1nAi6DSyiWji/ASFCC0DIEm7EOae8GCmis3F+6ZWW1gxWd0hngNZRthe+F3XJxz
AhzRY/+WraOVezLXpReod2+RdEIhBYDMmclWh0BsQ0gYj79vGery7olHgAfPuPkR
ZkOcmnv8aXy8CMOHeRL5pgJoeq8AKYUGWC3dE+a3wD1AVTxFCA12K0B+Kwp+gNyo
NYqCmlJPOnTBGOnqtXFvhhfeNy1SmcXSjkobXTHS2gsFEKFTH+lTlwGMfNVDDLep
uZNzUJSj0dST63h1e2xMny2wrCJ8XMKZm/6i8oxd8IgeIS0hrhTh9A8+uumIExgF
bTOU5dYDoUHJxb47dUZRfdxrb98bG8OHI6ds0mm+G2bdBjQVauwsgk7KOEJnBoUR
O00VHT1ekYc9nTuUUjgvgwfQ4UrN4eoVrgD9TkZiNygvk9sTpHM4Xok0oo7PWtil
pExZaPym+If0RPVfv39TwWjb49xKallwnZ2sQB4/FV3Y8M/GAEZLWdqc3TkHWM2c
rnu4K+zj9N6+a3xKsDyYxQ0nedXeLtDr5M3iAKi1mX0Ykz/8rLcTSX8Gl2m26yfU
gVUcaUm7y3UG5MdlfLh2Z9P3EnFn3oPQ73GNZYZeYoqYho7Oh8kpInHhOE+cLpHH
4+uqcYQ4vcWNV4PiNWyZjo1tS/r3jEg5d06r0axgH0D2s4z93hHxaKgrVY1xwTzs
vHgW8oVneGt43V720dqxsm0on/g35kqUJ36KDhl1xYLk6ghHxbWZixcroMlCLAn0
6PHVdhwnnIoUEmQaUaIOeUcFOM6XWZXwj3nbc/1Lzr4fCy94DLJcaal6JnsMneUl
BtmLENB/VOhI8WHOItK9pVs/sAVwfkzlFMOxubNkwC934WANTvzHZDHmAuwAprje
pp5x6EtHFF1c4vKY44zHORa6b1tpbnKrQWYmHFvVA0AQESpwOvHe+zb9KpACUwe0
0Y9LDquGP/N4oRfZZLXi5/PzXa5cqKigOgXPrz1ieNUnyQBFjGHYUt2oHqoOM+Vd
AtL4wQzT3wvEcJY9KPqdDhcGMGpRj0S3hQxne/m54XuIN4bUY5nX7rLr/uEBvxEZ
aDnqjNzBB9T9f6YZG77B7qvUUjphkc3uhJ2g/PeVo56JzCdeR/WckRzygHjZvvNM
ej/Zr9aiXFWNqr3cCewFBb//6VboiSu4RKOkBe2mw0vaLPELqsInccIEKdIpn4aE
S7pkiGKEqQPskblVYaT0JX0O6VegMHmEUfMDpzzs1lnG/2TNJHqmnCDw5kyrEGs0
D8dRg8J0z5FDg7L7WiiXpGf2dRUS+I0vjpqp+qdWtt9XQKYDS+dS+rS+kSiVa5cC
FuK9lIngHqPG/cWL/oC1RFqk/6sDVgLx5hcgHZGrnMMBL9QsBxL59vlxtPnjZIIf
IBd+Jh1YppfyEGRXtqtxZodPR7ioswXeqCsmEz/xITvEJAV0oDjw5RwMDeyEmsl4
wKbTbxDwYLOHtOpRdpAbyfm4EAwooC4L55XpoK0e0epNyf8fBwmwQEpHMEzpBc4+
h6xLkan8bAU2ixsmFpAU/mT6SvaauW6/vizLlG6+Ac6DVfOhhn6rkx1JGAcHJBP5
L9MNjIvi2wkiqDT3XtrR6Ep5Tv/Yk+KR/SZ+9r4uDbX5ViJEOcPyOrc3mQ4P0Uqe
D5N8AifhZTKrx13LTy0lG6tM6zhThlb3wdupfR/Zz7HrCWzjBNC3lLGEJbVLwQBq
s7TTVHz7w9H2R3JEw2eS32FAO3YjV1rOUxu2iLCMZiiy8BmFra4M/JE6GSlAWbiw
sPUJNQrUg3ftkJjS4KegV8bPPJcAjNBEGTwwSdKjtwnfeGGEQHWW1V8Htf2Po4pU
EbnHDU4B4fQUWRyngpe9pILGSlkxiOOUao3O5PzFKphsKxhi1tBVDH7hRyUjH8a7
cPPZg+UoWx7EnCOTBlLNo78YsUCRrb3kLEoDtCmuWi5PquvtE/AE4jtKarKl3+K1
IAMsAhAH6rPDZVrIUPIYgYiKj5ZXubJXvpmUcB8EUm+nMvkBNqkj6jwd9bC+wK9L
k0fCF1kFMdHTaTWqMxXCRgqW3DibuSp+kNpaCG4k1mF9gaFrHNmNHyoASH+owLM+
TkdtdkBoRUf3Eu9igiX0WoyYgQa5VP4zWVg2QoJW4HSnbvcRhYqWEWVWZfJlqsP/
JG2OPJUqChf0O9xHPT3ayPLgz8d5JXdcIGWsqMK4KmRyS843x3MZGJP5Tx51o6Nc
Z/ihENAzgJh22qz7Q/LqKnw6CpWlMjr0/wS10wJalXtM9GHOo6ZcMgnALhezji0C
9w7u8ydikJnbksnJfDXCkNXCxYfdygf1Geqs+aTHs82n/ft29kxiPTeXUkQe8vDV
lYGdcHZP438yaroufIpUEVnPWIQlzNumAUDU458Jd1xgvtsMrfwm2hbPJr1Xp0HJ
2RHZ3FzzRA77FN2PvbO+8VIAOu9jSn1eQrQZYwLbcCHBmbuub7pXJstSJQLYx4e3
PQe1pgkyOg6dW+a9t8FG7bNvTEd8PFbCC9i9LcgylQekxpq3xXEUzaCUXwLL6Rx5
W7f27gdalJ+TvIBYS917MyqO7Kn1eEEe6XVn31tcpgYNwS64DVRqvu1HNc3gouUm
Pybq3G5LyUnbppQM+jTubgiCmQpbgvpPdttQX1CQMXT5BOsPRUarLVFVb3+c0WEy
U7GK2BOUmLG8PzyrqrywnCgY37tcYRCc4Ty9UmTOaJYozCS/mNX2tT3N0fjO3eS8
yN5UqYP9pv705YyDMosVphds2AmEZkNLgSXyLQ8UwdGxukoJLFhq9mEhSLdkH+jl
+lreo9KewE4ECO/2JA05W3Bu+TPuNAaPPgjbwKIzxMrjgCSRFLs8peGhqNWE12T0
lKsx06ID65EvzjYuMwDOM0P3KkPBfTiNApfXEEGOKxgSKh08268N1oWZxbdwBWm9
R6al7S8SQtyonSPLeofNRKeVTifJMCIggHWDKRKAKt8Lo+NKduHWsvGKmCqh5FRF
20eIZCwxerFAc0ClXeFE/qY0b9/W/fQZzZ2jiyvpm2SO7PqHkPCVyi6X/rTBPWci
W9BvyylEjSESFgHr0RlycAg7zRHWS/Gh447N90yZcISEyIuG79rUYyap8HYpz55O
PWQnU6vs0dj5Dk5Ki1OoyVisVag+6Tbp2g5Mdx++fkQl6Bt9T2szuCjczo036s/X
R/LEFKDq7aYsteLwbBHVcHaU4tBys1CE4YFjnJmxbEwR+qCJlrSwroRxtjL59/Vu
m7mZzeZLXN2TLdED3QjFkYZs/LwLUVLkPa3IjkRPkpbUXuT1sd9mU1cHRf+Vp7fX
Z6ucZVBOdcviQiEl+PXAIPEFB4hRdtWaWe1tb67Kyn5Ao4gVjSmVk2kz11NURgiE
n9TRuoFx1mIByQ0BNCqsN8sNK8zn8wytbMFMGVeX2CCOZk0hxOFBzuHgLNrb06L3
7h/bY9lCMQ+9uyckNiG/szJc1azyirsxptdTjv1qAlpBS3mPVVMm0SOM886Fm+DF
r33EHekUFLBLM/91Y+ZeqRJaSWsQE6V9l8abyW0biZ333VP5tcUc2pFVA6zC6HhF
CBqYy8zygxu50sluw+52yjMcm7F96EgE/qxSNsZEbh3tzPda+i30rd/NOX64caSE
RCZIUfhJoLCzwUTS8q9FuFYJ9AboD3TnM7JFY4eI1j2syZ5JcqWFe4E2LheoT34/
/hCIYgH0d6mw2OZw95hdhR78CET9GrqPfr3SpnyfQx2cDhkXjfQ/cx3YUJEgWvMc
fkJNV2DfTEE7jMczgUIilbfBdwWsox1jrJ/gRjL9h8mn30KyCvjtvHQrHBU9zTFl
ZC6K1uymQw/R448Ga9I687m6zK5IP7Lo1aYLaTkAty3qjAfTlLlmIf47BNbay4ux
gxQ9ALJihzmLZlpxq0t9JS014eJCKmJl1vyEvz1SRqN4ympUrG6Dipzx9FChVV8X
q9cN4UOrUt+oIOz4rdTsj46zgLHx2/AwOcWUz6jbacCM++wXuRtPEabA6AoZD1T7
GdMVivbU+NjiPnAq2Ql7ZJLkI5r5CB7cbC83Bcm3WbU77ns6mvxCeVWdwQe/baDJ
q0bfmX0TfkaYBvESLV7ikdEuPm0Xyldtl947iWiv3Xr8CLaHGyfgOIfsd9jSUAhb
r/e8iHj6iru4ldYmVggiFrGlr8NLygR7nLTGvgMAFBFeaRX/3RIsMySQMAvkrMa9
fcQ84zNgwjcGngngBe4P3dn+ceEdpbOFEEDX6iCHbzh332mi261MTc6dngM4pG+r
HdhiWxawQZlwdYQixOSEOgKoYPjjwZJUFh7F/fd+KSCKTQP93vr2Obwz4O206XA/
IB9DoZIY7veobfw9EMf0fZ52DdekEN3st4/00nKnqGIeziKwOEyTCNYKuKWT/Tjs
4tZA0L4mAllXgwL7UM/yrPRSVkBquDlmAU8S7u/y8HCZev4hcMY+6qmFXSVXApyW
IgHRs7XLF3L0GDG2wrfjK2nPMiJqTglCYkO+3FqoZ3ON62R8kYeHtjBndMwNzYuj
3eRl9ijM779ItwbdzlgQ9BMA2QN5ujO2/DAHlMPEvy1lrWjRqtAKtsFlNFf0D3Bl
zUEiBwXuSKDGGDIrV3JpNEAOVlfEaAT40bHc27w1qAFC+RBNIX643oEkDVzxq77Q
VCDLrlfdLYlPW69SKRagdZN0LgRxpLbF6cFfli95IL/RXjUkXrImF39hjyjZN1pj
611d3L0OOcyKkpHHfgt7KbOAbF54gUXvwtwlDNcjVFai2YlLn7N9cFU8LZCe1PI1
rQ1EBsPmfO45XS9LgCFWktWTkYvFJu4Bcf3RgJyRKoZN21DPn1F5lHXba8cWMCep
Nnw0B6Ruxh6Urmrkoiylrp+RYNvQgOw1rZSn90rrQ4Xp6Vsw00q8jJPQefTP44pe
GLu/MS8ytIko1PNHKt5IMb6S9oaBYXV3tu5qpd5shthrgCiBXwpYIODRJfrAsACg
kIyKFSx3T38YzITPseQvEmipusXrDK/g9CsqnWeOMT7n/gFdfcCqTUjAKcaskkvF
q1reYGeg71Ac/ywtawXKxzRJBgTnRjt9/siUv7F5Fj9q8bP+jXX+8ETBjk8P1pX5
WOzcINB7H3WV4kuBlVIMHON9qFGSjJxqxZd2u4pM5tYeNAOyeiFFeu46hA2TazNI
hiSwt2lJc6mhBCswpnMAi7nPHRyFy/UDwjA+Zs70iLdh8fjAECsdGLfI+s44x7TF
2qtFIkEZF3oRNFAjtu/fHWyoU1D1NN4fwk2yLzBZI9M+Q1kgLuGdMHPcwG3Hb3JX
exZiGyg1Qv5mgjrXrBJTwh3nlwub3Rh5PQRWIKPP+MH+vsI6tkz10NCGeGd9rIPz
7mBiQC/Q6ENLjrSn+YMVAirFIxniroB8DanaNyYjyRKts1buLTZmeEvQn5CN4SIm
BAWpGMpJwDWDkzfvABXuhmyy/xya6Md8259ePv4ISsicUJsdrujLgay5+d1x01ff
NIHsxK5H7VagQg0MsVdOid6GB2qGJZz2T4yMou3shXCLU5ktc6E57Qili1MKWa9W
Xe/eYbaAY+862+MG/rE8+WRIIkTU9sKt2qZBTlaQxcnrKjXOH14YLXAJujhutfMt
tPDoJ2l5jCbUiih5UJhH1A+HQ1T74gDANVvM25u7bmEE3cdtzCn1wePJfTCLSKSd
3LwzEU7Dcu149PbcN1UMFDGvmlk7JR7RVntdLaOxv7sw8cLHKx+gRdw4SqFH7sRL
dtRHWZqQfViKRUC9hJspgiTLyuxIVG6Dtex9T1LpHvdzV5hRHT3Itut90iJHpcJD
dgHQJWBrcA2mgNHF5D/JOUjDJjoN7mmO6U3SjMbAFzmsPJRLNx0ffAbWgVd9KzQD
vL8+SN+RjeAHHd+jdORumpkgdEt0FU6e6ObdYQ49unWK8febxBLuelSEOrqsj5sH
YfwgLgsGBWZNfng8tczfZm0xm+LEJignvCI1Gur6/29MBZhVOKARiI22crbI4l7P
9hphZeoSSlSmAErxUrtInwl2uMqyGKQffDEIDyBNCTZMvqAuho5mqhNKZdCKJS02
QwCjc8LcVNEXlc0c+m+ErycgjYjpL2nz4FnHFFDzFLB4toiUL46Tu9O/14DJfr9R
1ClyBOk31JvbCxE8CiqZj8nZ9nbmT6uLOjwF/5+SojXi83lpzjrQAnbKs1bvdvtf
w29jvFOINZ600xCGMdo7OJm4EjyHB/DnljMa3DypW5yAD/AtjndvkDfvvSDqr/l3
GPX5MLtPzA8InyeqaWyYwJW56OL+ewxjOD/DLazYCmiR20V7Amqj6bDNkhCX6FpV
OZs020Ju+oIw9YV7AGgCeiNfgonpZmSIeMiKQS/IDsz90J7shbLFYB0f8HQkvZ4G
X9GayGzCTOH1Q0xG8QaS808IBNi5QUO/ByXxtgjylkbQM8/J5ksh3Lx3TGj8kpcI
fjNqulwHnWoDuvymIfhndzOZr/5kW5AgjWw2ubQxW2SK2zx7pdWvUmQwXq8BKkVR
wIraRCE6TVnH7HYtvEUZBmyc1wetFRlSgHuhQMVMoeOmP6ZRIraD8icq54ERiGfi
+h/qqH2o/qsmYFdsX6UWC+FrKUaTGISaPNp9RrYU0gDj2tr+cFxx8AUxSxqDDfJ5
55+U7+hzOOY1YRldxXtS8U6sMXddfJXACWtfnblv4ovtKNpbvxeqtG96Qo1nJoXq
vCWbSICdcUpnrSREhbuXWnsYBMtrRJOM/INOa6qJfoNQBytGQ4RGovKpwoZw7r9C
TS4zrIfA+A22Fd4k6lKki7CKzvW8WIRpbXtNXbT44U8iOjP9DJHZQjvl1B6gt0xm
+QwD1LEzFUSCp0ZADcHf/dsxNdyl6/i2UJ7zd+vwua8OJhprrbsOw15nJZRvI+ut
U+SH4yJYIIG3iboY1b0eWL7+TWujiu6XJzKrEzR25NFRo6Hf6kheytaxjTDyM+ZR
+Z/z1o1tiqIB4wmnpRJimA4thuqXC2udFogct9giQ045bo9Jg31AQ2JYfWLtZZe3
H+0nhmuiToenY77RW59HN7cvPtfHZuBvyNlyGUJi75EqlN00D/0jIjG8JsFnQWew
XHxGXTGGVujqEUVClehwRkuehGOgBre5X7RTQwNQ8VHnl/P3E4/mIkxxNowJTvSA
Kz6gDSIftjWLcUATnsz3WrRie1w89I9cg9RkjmwPu9VFhWo2ZOYB0HzknHoHfV/C
3kj3EvXEh5wCDS4vsfgAEZL/+5Dfc92kg/Jrf8DFMZ6ZMVoNd67MvyWk82fFLLRu
tj6wKLiiUCdH5VExqqkpD0NggdinMhNGw5zQIUhGg5pKINj/Y9/2GTfS206cLCCQ
zELhGYfG26SR2OORau9JSnt2Y0Zva+UoVZ+vjomRA6G4yeZ5FB2zuxeuTEjr3Xbm
FN2hbi0pPeWKUCOR/Ic03cq5d4T2grUqeFrNch7SqR6+wQHnx8zZguXZTBnSd35Q
JbIy2nhR65auwomqCzRkVSKCW6wFFAXSngAAOA2cxrq76X9+AFCXVwEjDB3NnfjQ
8JlB9YsSFHsTBeJmWDl6iibgQXL884xOi8LFICfMFjcvoPYt8XS2+h44kwsLiOXG
xoesdUtwHCSc2/zA3j7/ozcM5QTJlf2g14XE3O9/YmF1D3gLXnxPoVcgw4Qm/j8E
nj8Zf6Vi9hs1nH8cTIUoLf1cRdtNzgVFDmmCk7PgmxWyChe3JRdJnGFwvKfzAZVw
tpuQiPRSpsRqCNLfrzS+m2r0TC+Lizj0jh8kQUhkxtaJPikBi4amZzL994oPPOpw
a2V6V7vStUUmXHfcvaWsDrI+D37113VHCV1mJFwRZdSiWLUM4+AtysZ/uIdFSjTI
fKbt/TBfeMlhmuMGs+38g1vIxr8UsYhne0cv6bx9XuN4pAyqULm55c2s/d60Uj4d
tAT0NhLoAd5QWqcIvwiIcZdxsjYftNIhL+1pxXJTs4cd+yLhQCa0UFFZBbItReCC
egU7w9pHFkGX+WS7YHBnkLY3xxlw2agNHnkrZ4VvGQsPClbjXjxPBYX4kS5V1Lap
6SqjW7ug4x0/kNMjaJGEsU41/nZeMYv5jDa2rzPpJYLT1hwOIPvqJ4D9A5ikzAiJ
Yzi8vTHDiNynzXiwwi/zhz1gJILVkQcZaGQGeld9LU1XH5wDQkXaSbU5bAcZ+6rR
NpLR9+mPomatSGMWX2P/0ws8q8tFqZ6Kt1vHVLbJhe0f8Vfi4MrB1sRbBUMA+xjo
/l+8PXami68MfZ3LN8RciBw/CmCXLlSFHwaUIeOFDUQnhp0hypOLtljC9jS+7Rbp
cViJtvz/hrOWGeSLpWaXm9L6t1iVp2fWDdwVppsIr4TCTnOpWUZEarfwIR8mZboj
A0rHJPo1sbmuiQKuTo/xt1xPCVxXCEyU4YWwi1cN4PQ+zg87/61OD8irZ+slbKmV
u6X1xV6FIjfK8b9/QPGpC7L+mUlV6QLzfUzSPB0SiX/y4fwZzl0fqbGz1p39nnuR
lgV4w2E+13zsycCIb+4NtwC96rfLj66CQt67Sanayd1tXCzXN73RRjUaY3bpUXOe
ofljL64mAvhrebCBEiUeNj4XXMcRzf0FVyTiri4B6mCo+1aZdj42r1C1/TQl7xoG
VOHbZ+VK5IdLiUMFDJ71okjoom2nLQQtgB/ZAip8DKaiVa+fdmP8eEW5NTv2T5Ne
D+Fl4tZkdm/lK6gK4VVyP91msOFiRGSNWmoYbHVWYcS2J/pTm78Qe3ig4Y1E86JZ
uV+FBZh8isea/2t/s6bIlAfD4tOL9rsM/+6yX/7ufQnkt/8hT9MJ15TMRfiC1kDa
Nbly1skWDvoRg6bh/lSh5Qh0kyfdgRSmw+mJF9sQwgSFVMhq7KznZc5VzJ66/j5M
6S6ZkIggtBs/icTqURobvLT7J4ZsWE/dCwz2JktKAFUdxVSvN3GZQf253Kk+jaX8
8AYbDAoKLtapqV3NmzGb/Sg1K5LNbxashJ7qxhYJhoj6xXRkKuxTntI/OcxgNAG6
V6TU+fw7J9tVlj7wy2mAaHD3qs0GmgwQYhb2cyxoMm3jVwOXdngDVRqcRBSuBT0j
Ouhek9huL33YNvNifnmviyL7U9tANptytXwa27gSTROjv/G3ba/qOlaH+9kQbqT4
vawpNUSkdnH+HTDe9sHdl274slfsyGfp7SVoHfH8l/uOqXokC94UAdZFrQ3q9dCs
QQ2GTvQDjOHBKuYd7d09VxZECIHDYdgFPobOqKqTiXN4E9mBpnBX7Qsz14vtLtAX
UBMRD/sQrVgwzXYClDoFRoSgiLMt6S4U47uqGzrfh/avou0o5a+u8N2mPfaObYB0
QMABo0o4pbBiFQUCdugtHTH/FpOgmmRB0pHuYY27InBtTQbUOrDK9qFYeu0GW/ae
NDfg3lcG/UbPnG3XEo+itLf3xjsp2XzH+Qg35YdnOE1Z+ejPptSIYeSqdamUJugW
oqTsXExgJRxl9p1m6w/ozaSaq9GisNJHnrh6ec2Tv95dCz6Xc9qnRFzUXXDjTvJV
Ms0YA+MwpDZUMbwPtNJV4S/8MyLm0pFYAEJEJe3p1yiSMpQWxq2pVPXMbQFvuyBU
Wp1YKDzi0U9W5u/GnX4RvBzZx2vSVNw2YQeuxJJOsmEkdo2ejVZQdFWS51RcFsYJ
ZU3PbzsUVRmUW2RPbZTrHQwWqpzTy+QWkgSIVLnYI/CUoPtIwFHXvr/P1W5T6mNf
GY8iu61Hu3GCsz93LxWSqn9/WIqdXBMoQBzfVJ8Mejamsp6MnCh3MJlk+TpCrQ2v
sjydQOZ2bnY9OfIXPqLQGrDBxV6eJYHU3NF2eKbPf/FaXRM7Crdfaq9UQ2wq+1wy
x3F02MyrxjCtNB4XDyAee0uPlc3NsHdddLafk1gQzP3gDwkeg8SCX6+etuJDkNd3
F/nHRrk0lIAb6M1RRu+5rW852UNNm6kvHo2p+1LQoHk7q+c40qTpxKFhxcRBy7Tq
+zlxtcQ4/EfTFoLO4G/Xb7AnwvzssP2MEaWci+5XykmCDkBBjDWIQMinqBEg1C2h
rHE0mPTB4YgxMzAIesDAQRacNLmsyPCxfwi0OVPeLvNkMju7alHlsOI/R5s5QIQw
xXQ/xRCdC9af9jWWVGEkGM6vJgfLN/Kote+caSLwSHITn1fMrb5taYQKC/TxUeMN
BSQuzo4D66SDTEe6PTNiagJp6u6RcgP/RqnB8Cl1RKM7uPCVkBcvRnc4X1q5GlZf
OWiFAwYJ/muo3U1XSbGhppbS8gJ76xT4NJYHHLMKfDYo12L9mLB5WsF0kN9wQwYe
Rt8rzF65wcLXM3757cMlDPX23pw4yGnpSRNcm9PXL2ozU3XCsg5WmS7Rko7Fjpbx
2wpYg5ZsZEJoVNKVIK4PIUI10jaKrZ0ouatxdwPKUe1VQXvfwBxAh0L1dHV4n48C
nxrxl15HjurrdG5G/5AepBIu62kps8nzn04ojMjTNAbYBwXvrr/HxyrAanUg3roC
uJYd4YEAUUgJk3bGAwrcrnNKG1PpcRMNrqEP0W357jaZPpFvRkKy2uwExONCwLmi
K2AYFX2I7oJ42okH6uc4wacMYF+SQiMIbg7p0teTnVdXbrlXLIHepQlCPJVzUFVn
V4pMdf50ju19xIagO2zt8q6Z2ZFVrK0NlDSQOfgM9U+F1XdeQphiIG46UKz63N7V
IF4LSiPzLyMzjkIxdcmVCSvNPytXfdkbsXQSXF0+Ih3elwAi2y5IeKxP6lQo1BZI
SHK7LMZbHpxYFEUEht0x7ax3Kgnxriws9G/ywsoTG1pskTA/bHf2SmT0o2DhCbKf
C7LhX2NhqQXVUfpjUDCVOCucW+3a4PUsxVEdxpy0GuDA0qHb3MrveYfDIuOzBw79
sW38v3zrBcdAsw6guarbepwwFufwRgxEEoeRyfXhHw5pnKWnsUEOxhFBvAzjKibu
J+pivgd1jspk6cRfg0ej6MdrJKHRApUmiA9jdiXEf8uVWP9x7j/9kb4XQRSV4fUP
DAwakDtQbulqlqop31B4Zds0+Sv0VgVyaffic1e+AJIOxGRTK7GpvpX97OhVkT7d
RW14smyVfsaJ7kr0a7qTxR/uITYlMRDaxmpxEndrz1a6yKoCvFPl37pFI8YdaqkK
gH95sAZVuQjGuMdjF5sil0y2H77DyGfJlEEtTCF7bnbxTyeJEzc8+mbyM/W9yhUN
bSpW5ZJGj0DhFFgaZWScBM59fSmgwX8JGiWXxYJZtukGYr6jRMRVDtl5zVZp14k0
x6oUPhniG97li+nNGLIBDFUCoqZkVLlO1G7BnjuJBjZSDxDwuMWfxrFgLl7CrIQp
+xAzE69GOu/sNo3N/+l5d8IzZKD5nV9LZpBE02/yDLi5NFVhhODbbJbvsyEu7dq6
cSprEt8YUu66nREQRn2dXEVCpPVovtnSRtOb/hByCWpyVFymltaj8LM/zqZVMFsG
M5hW6QyYZfl/E/nnric6W1SoYXrPCHJn7wsRz5kKpOyoG1qtYblY+vOc4wO2FD0O
WDlG8Ko/98k324oCjwiZDLLPm5ln3utGHLwse6AWBtdqHMo8jbpdskLYw8Hoanbj
ebv13eWq7d7DR7lA9e8pqewVaJdOLZsCZSHK64gjG6B0m62S2P+zjh9tEjqN7yAr
cxFhOwUEb8UiyfsykdmZIcnW3URRG8JUblr9Lzsu/gJzgOJBofSiXUuBWHx9Aln/
uxILUQ1665DFRIlt6vFCVC47Y5ZtvQRRCyQUeKY87i+4yTVmxekYZwyR9OGvpGx9
4q/kY3DneizDt20LBbP07p1rm17vj9t1xxOH6ES2XzKYUYMwSXABwujzl/zgJOtj
JTYDxJb+Om9ycsilgLMLAKf17Uc6dPkC19TKSmn9nrLO/6RYMAWx5yCcTCCD1aWq
u1PPu1yIYtPM9IvDCXwenl62aXA3EiQgQkJR/kjeweCQ7n4xVy26QQrHaW3Salk8
ZV/eXiQtQPWQXLQe6zx+Ka3+qxdudg8qtfDcbeACroBoT2BYcHMgT4/K/+auQk8J
ksGrxr23B1cSHZC93VQ4gU3I2bXSS908j5Pn6ebqHZ+Nl7gjlF1ME90e4l2wbx5i
9AhjtPyVmZIW+fkdC8pmuFgyBkxF9TQ8cUkH62tDu5H3Nabf2AajqnMbpIC3J1me
/N4cDOobfE+9TOqOXBxFlwfyJacvFtQwGuezG6dhgaFsQtW9Z0fQQ1Dc0rmPKpqU
y09SMiVkmLeD0v0mJ0MHtTD4aisKIKvP8RP2vAoz2uGX/De/2VMjVJUVP8SJKfTj
rFDV3DSUL8Zrxmd3ucZG2fjLDwrYsFMn0okDWb7StEUQYNGjLqWgLcZODlzQyBdi
WTy+D3o9P9Q+D+gmDM5HmzT08E0D+7eZEEoeN61Gn0Uo0MGj+WLm4zifLoTaqIww
HMNOZv0j815y1YLPxGWLZwGq6r/ZaLuxQ7PIC4mXUtGKFVVk6Q3P/jam6jGKyPA8
qQj+VQ2PE972TUqoclx2t8rB7amhzulNcOnGDmQ7JA5va1SMnc5v0vCn0JgJR/qi
V8CoHonulR2+YHCcWqp5V+MEB1OanFolFBs+LdlDrC/Yyx/qWLdYd7VXe5i1AYkf
UED4u2nHLwNjLyJ4tuPJSxv3RAG8IWvK1PVU37kS4r+8cqSl4wPG1uLmw7Z2uQOE
UCpkJMJyEHwPBp70ql+UAv817jxWJRPSuOq3iTPMAH6K++z8UwM2aHgTgd3Rx31R
ZY3AgORqGPrn0qoQRWNdjG2xufe/QlcjmGrdFyQpwAjXi+rMSa/7BhcfkgVVe9mA
CNaYtYSyN30RUiPHeVbZO4f0O0+ZbE6ZsJVCl5iUP4bmabXSzL4YUk6p6xksxDmr
YirKUic1KI91kAp6gW17oapIYBFhMgAg/3TpFLjBRoEW31W1o+1cjV/52xlN6vb6
mxq3o6y6CCPjP9wtOfDrO0qlyVptxsrIx8YKG/OMJO3HftfeShqt1/XJ1+UZJ5op
8Cq5Uk042nBbcEQ2SbRB5XoDCsu/XGtDOCJfwFqAUGr92raGoLq5gzUecP4oJhX3
Gi/26N+sRUvDg+U+6Ihty9KhrNNk7Zu/dmcc6HQaTUZjhIpUenaTuWyFVyB2UAG3
A4GB2NykMRVOjoBR3I53AZ6czuQtdSEu1PaSw1LIaQIuznshhCjcmLpkr/4+kIgV
dF6p/zzaSd7Ke+CD4wXJowP/gKRaeSuYQMDwsjZVNDUb0Q+OrjZbKxaoHYsMlUBT
R6OO1H4VNwKsr9rNppzwJidJOoEbs40IwebuCXJmgjNqqhIVKL+3iCTHqjLXdqc1
1fxzVa3uaBvcOR6GRE+x8rXBG70rFrR01Uf3ZDpfhXDH14Itj5SspTRoTO2GWR9m
RSAQ2/ctuY75vFrJs6AFM5yz+v2q/jUrzCGlVhpFHkXVrHODPccZtGEc2sMG5e5/
gsiVbgP1Qjm75/hJMJbpqfaF41FNWLM0sUCfD8OSWXxqmKvwZ2fmmn0UdJWg86fv
u2NfZi1UbDxrDknaonsiTZWbxVU7vFZhprXostrmX3S3N5sM8X+YbsjXFvSe5nhj
D+9wdAD11Zdn5wgQe5OPo8RCRcf8lODLuw/g2jdoClOy76+wxAdj0DBMWitTD4CB
B0cGDd3bqlbUG1DH1Vrlm4fo2ABgdcCEoaJZ0fjmY457KJQ86MmEZKdDAG/LSvRr
jSjj1/bauU8dC3JlaNWWNOIXL8pIl7lPmdkNRxebT0VIrEeYf4jgxlF+oU5tCtuy
NVdPuIfORnnMfhCah9abk7Xg/ZUhup9rx2HSwsI/FVNpMCY81clDXNW3pnvsD63K
jFl5nkkJ1LVgrir1BfKObFkqWdGruslbbjmtgIhslFh1Ebd+eNFdRGS237mk45/w
UXWId2VNhF2B4a6hldMzs04DtrjVF4ckyk+oDsN//2Z1caVPnY7u5pXMDFCNbwue
Hixj0ryqruiyjcBADielTMeCXzEKEsnE+WhdlXhrY3rhqPSHd1H2Zke1QenIzjGb
rgOJE/EkpPkuzJHK6nesb+vcyI1MX7I4xVTywEdqJ+8uKkNLg5YEvL8fib12fvwx
LleK1WCwlI5gBELr0uEje53nHdUhlFAB/vIn4g/9Vx0SRAmjWeujvGJk3eiBQzX/
1FFrJ5rVxuMIVsh0stf+pMuUmU07C3eOAl5/KS54wnWubrLxRg2W1Pqb4kx/P7Dt
BZxH2vEXLdMRZW+Yo3+TsKpPNjXmYhCYgVjveVJs+nYT0Ou/G1aERTndefGyjFob
ZXDxGs6sbdtq/El14lEBwnR3PuRrmJxJ4ETWUM7bC52Ra5+nvynnpPO2ytturIuD
ruLnIDVSVxxQt4T5zr6lAbwvbjDqykNzElyiIC43bvPRnE+ezmDtxJ0/TLN5lFgh
YZR+rNx3mFWcwJRXf7AVxWszPuUk4L4eTVcSxNGxcTZmsW+feQcNfbxr7A9/W2Gg
2RPt7JveQP3pzcqU2bjotk+lxZZdKc6ueLKckz6+BemCK0aU++QcjnRvgP9hUIMr
U6XWryWrIjnqQs1pNw7bwqXvZhfP7mhmwJYY/AW8eHJaLtz4qHoE6iDx+iBQ2Eow
QtcbQQI2modRbdGsGLGZloo+sXimbHBzvV4PRD8NYo8NI13RklSjngBVA0Fqk3Xk
VWPxzPABKsv9akh6jk73bSjkif0GeWOPMySuONaZFoKxNkMXXXXjkRpBt1/xGT11
XkVcAVV11hcdgzHaQ9Do6Wb3GMmdO54O39jiXilv+44jdd5gFe1YZb5ZFNaWuZa8
wYI0gPmYK0YGQJYbshJejT6UoDzgRlz1W+lf6WAyYiZ58TvDa0L2waK9o/3a42g4
k41csmXWk2Kfv8C3dHfJfJCxrQURGo2ckVSCHMmB3DeTGe9bO4mfOtaL5kpgc3An
JrM+/620CLOrSdNxFs6s52b9htcLPrfXFCuKEEp39lV0jxpBNR9eLlruHFG5magX
iKuchjKkKShKbHoIxjF8XFR8P0W+WrPI6W/t0z77Yred31RX7Y2E3q0/wgsOBRu/
rdTFNH9H3X0o5443Yjw69P7/wjV6eIK3WG6EEsKtPMEFSgUabF0qcK2osemrRex0
2N9OSM0u4AI5JmVpaMKPvbP0iZDK49o1xI5voLxUwFoQ4ba+tq6yH6T0rt17nbEk
e0idFUjOOXBOQStADGwylkw46Kn461FkSLHKpor4ME05XmyQxLuvNr+C+tNfx236
Dt6Mb0G0kiOaQ2kWo+eK027UMAkuhur9K3maORb+8TiHUF5zDls8qENM2dr4PW8D
ZPAPyH7AqaQcK4vFZh0NCJzsaQHW+TkFBxKVJ4H0CqEN3ssEMPk1cCbpgYsomj0b
K+BCP0mVy6qDMwpnsMeJNfThXnXGlp1IYgjdpo/wtxA5Uk99R0EEr189DyIiviZ4
c9ohNudEzirVW+tpEGeovk6kX51HF8f0LLJzcQfx7rl8hH0LSoVr7Aq/7mcbQYfv
7LbFnDTK+XgmZ7llVqvnpG0hu837HmXoygmIy+Jwfgv1BLUeSbUAARu8cslDmUxy
I3+3oGrqJFeo4CxDs61BIj0/fRXX7bCR0khXBnQXIgmV926sSjztBrrZ9Pk3Lwqc
vEkrMxyUw709FIm3mFM28qVyvrpEKZ9DSySx6+WggtxACwtMqyN6dHhTZDeJrshA
qnEZPDzhG8V/Fg/gyOPn44fqNxlCnCPgnvOk60/XRPRHG7CGFKsQ0C/9DS8h7/AM
NiY6jdIHNH+QcLPaNIX1gaFnC0CQE/DcWPSS+7TFRZSA23XVd+eevtbySVR4EQes
9lUTiTYndX3k2VepX/eZj2sWW4QqZEDjdoR/z1JiimuQ7twWjXLPQi/JinI/BIuL
61Mslg/ljNhfQ08DvOGjRW3chiV2gQWzVAv6pk0Xmkufid+UugBijhDFxoyC/OzV
oQEUuHc1OcRHrjSHqHQOprtLyrXNjbtH3cRjDLhWEp52CxJ29SRgf57NG8ma/Lbb
5hsvDC6S4Id7nsYqeBmzbvBElX/cZYGmWb/q9x2+TUJ7pm0bJfDYZH9BJfcLgRzA
TBKkYVFfNypkP0PQFgy5E4y3Rm3ECoT3y7LC9N5L2NoiyAE4rCJ9g8iN4Ntsdyv3
WliiGR2k3L+yGxg04pTi5bgH2HF9YNoq3ilWtwSniEOctvBI2l21AX5lG7sjVd0U
6lg9LsXuDKXsyBokShY9pf8r2Iz4yoYTS0y9kTXqsAsgED3OnenCWzTzmBlvrlAZ
HiVqbH3mrvZ2+Lfynwnvj4B3XGwKotoRRHYjhRFywsUAckgLjABfxiqIkV4Xb0ng
o7y/NnOjFZtIO9Npm2LEqOia46kLbgjsh412vU4RrJFxncD+Ljqv5zqmzD28qU3+
N5kTnNPRDS3syBN+P935Rdpj+rUorbUwn7JrwDtpCckIAGh77XTP/xHZgYjTlhAz
DkmD+ZhJdpI6Wo9vHexcWxJr4CemfzGYkZcjeec9dLoSxKrT0mKipaDMaY8keh/5
ux3CE3K4sZp/Y1/SUiY5V+eoJBI+ohHmbeyKabzZfBdfxQigCDNPkDtja7LbB94y
wjcsXsoQ6Xq31mYOZQ9cuc8LczKQL+xCDlReoZuFrh4HWL7VGKKLbmdxR6MSsMNJ
bk6J7D0FbMrsZ9FaCbMPNe7+K8nxoYbh9/CFcUhjoJOKgCXqlTrxzF3LmcMEhtVi
LX54M4gexoPEhM9Tz4v12ZbBwnBBJ12SbnIP5+HAoGOPuvXHKMsyASV2lZ2nyW0b
48c+XThyEKhzy7WELVtZd5iNGLDRUuqTGboEK0kcP5Rf0EpAX4SR1eJ5Ui7IbkLG
SDNW50kjTlYgIdkNNQN41pUzzR2u6LUWFbBOKLiN8TwJMzhILR4cJ5yBcy1XZVFN
CjIUKV2I3N2am1r6zhwJxn/4Zg2nz2GKj8UO9Z+2dZT1PYwlSv7PnD7ibCOwe71g
ShlK6LOlLa041MCN0QihfubO3JJ3wQuhF4XS8Mq8Ef0RxiEbmg8sStUOYnk92hU+
Xi2aQXG/eXvvq8b2qMexcwI35V8mPLiN2aUaX4maAVD1+6HXBb0EQVdKhIqg/4mP
W7a37vT0sPdJ7cxpKrQ18yvuvn4+ERD9AHGBM/UtXxJ1ge8QW5El7Jax5tre6bwD
sSEWKFZkzNCNmAPbqlp8dmqx8QtruUAOtNjvN+iYU704xspCM3/BAGs0Cu/lrnsl
di9ZbxEbhkDL3jrp7omVs4DYws8Y0xjnfhSZp5J0cX8MJmAkfT9bBqh6YdvLw9OQ
LOeovIrQTZdnOw1UXC1PM7yNtsfHw6QfcVjgHH3TVd9xYq6DvLwuqKsqNDwc2GFr
2sWecbQc7zHmgAGQuTa/dsC+ANl55VVQPw96c9ivTMknDmz/LOWym2vfP7649/4K
uBZyMvfF2lF5CR5iPsDlkUvwQV4Gmo2T3oQFrqBOjsx5YbQs1PeNZF0WNvfM9dMV
/m0+Fq1aQHK9IRD08ZXfL4EkVzgWkKxgTzW0fEcdb7K/9Rc6QUuIgfVL1Plhk/YF
5tXWgdW/vNeSLi1jc9FzbZrl/dZ43eCoTWbv1Qc2ZSluVJNueK3PTihS8q/FkZaF
FhTujPUQNVg6EVgvdFARI2ZCvVbqv3qmQOCzB/zMO4YwxuCxM/MuS9mfA85dIIzG
y6ZT2/A/k/YIMXhybXZO0gwg9YHit5pskSovDLgPbwUJUdS7D7jj1qZa1yUhPE2U
GybFMs+kX1MZa7TO0g/Rvjz6uyUeZhg0JmphKeI/S83TXtKdtaq15lMcrXBjvt4c
JQSFQ1epPfQT5hfMh8xBtHD6VDk9kPibB8QwKaDuWpnMCaWOGUMQoLBT+WIuaA4J
WIJf3nTShZWUhW6WKBpdxZNinOU/WpvNe+KN/io+7uchcxtAdwEotFKkpCOkYp31
mIDioo4m/W2JGRDlaci0I4eWLGOlWpPWq72xseWgNTwHdkLCwlD3b1drvBCPUSvS
sjSwpAXA5/LaAExALVKLG3KeZUoBncigbrmPpNHfK+NUuSsB4ECVJzjFhxMXnkd9
s1qqM6EW1KduP0/JcYEmzlzfBT5YPvpkez5cFA9g/kNgdunOGXuO/psSNVuT/vzr
fptmY42w8LK/mWikMx++WTr2ah2yUBZjDNdlGv4zeL7k9/n1NknfQUfpJY3iRqoe
JCzRUkK97EZQ6CzjINoDl0lqlWwdFwcsD27Y+0n5dRLP/SF0eNiDsfekE2/FJcXm
BxN09TZAQGfjt9wxX+IuNSUF/UiNc1Kkl52+jq+lZu0iZAs7Rp7ZjU+A0dbYM/h7
fEIiE55Ylk0H8Xh4pCCdP6JQwrAODh3z+ptloi/PZIBKVD/ALCdZVNRI6j6JfKhw
FfhCF/AGaRLFry68ZoB+nyZpsL3y7yh+TlROQ1tQOB3PA2VSMUD1MakP7gWOx+dc
4ar/SaNojbcujfBTQZBPyS27gewDUHUqzGAiSAl7zwzcS2x+gEvnFPiOrftBl07d
qT/8A4IN4uUDFyEv5PXlNmehDxw+ka5VQnrU3klo5xRDMO9XrzynwjgQvlJSCw28
yrG9WZVdUgvi+5wFsnRN3EaNKqriyJo+ghCiCzAMrPpQ7hO0Kr3nd1TjNZNkP4o5
B+t8tlXoh7NziEroULkhIpICZePfLliQWYSKFlypSElVu1NYFtvXvJZpxsXq6G78
mfMq28LpUZ1EbDIk6VgMHt7e3POYnuuld+YOu5NeI61DiaVdcff5GRVfYFCSVPL1
Eu+M6I1kvPS/GJm8xAPnOwPmwxsY7bW3Wb9g3HG0nJSUIwpeMv/BC6vuxQm4KeqV
PjrsBgInFSf5QSHwmyRBiPpAZIqW2bc7qt3aVY0WLD4CBO+4LRfr4RGJobY6SCtV
b7OqWwDbgl1TldARI71IW6k9ejBYtwzLSXJ/cR3goxJUdqyyZFmpr1OENTOMaz3U
5CKifr53Mtfagv0dOptYwNxFMt2Yu9DnIzD4UX4LqUMHyaE44kgFbAQ9xYujvDQA
4vMuA/lLZW6BicJZ4yMVwB6acGDDO+VfuUjpfgnF87LiSCEWJyNs2EGPSZxyqBm+
v8hDjopjQ2g2UTLRFWNbcfKguhmOa46tLcvIV69BUOys57pNFoaY/ucSVwP2z+H1
3AVB0xmTK6ZCcW0O4ODj2wFkz4GVldV6/pSZ0VtQuQaFlQ+XVoGv/vEacp/Quos9
qlRU8lVaQfIcBVwjoKnPvMTTAUZOoNL2pRfrjAT2XKRXoyX5qN1L8PcqzH6DhuPq
gqEhIYc3bxpHMziDhNKUk9Wx9OmBimZoDO/tPl1ybpjjppKh1pdCkKBULqQZ8/Kn
sKCyQ4qq/iHNhGw5oMltdNroZKmqrX+4fX4pXMB18B2y4DjPMwor5dfR5/N/9qbR
NNXkRt7IdDSNzqNzXUNs8A+1lKTb5jmc42owkSANeUQCu6wWamz7M5BLIf3sPWMk
RbMf/DgWBswBlHAFzw3qV9K62v/rwYRlwMq1tkP1uf3w5qNgAiL9Rh6gNKOiVbr5
0Er/ueBLFImPK0igzJ42AwlMqVPAfiQu5KBK/8TrkoM24d3rdfn2xnVPum+Pc9Uu
AmSjXac3kebMIfYAFQLoUKfa7DLGbNzBP4YoIesFdMVv8MFZtnfOuHYq9h00kz7F
B3pI3ZPokwTtbxXWSntbmxhGTbaWEzcS0mwfIE45PjY3xohSkl2XODiN7niIbpPU
JCGezsDzVIhPx/19LQBSGsZ+xveyQ67/slK923pAnn5O4EupSFde/4WZj/90SQ4F
xkBOhWZarQs6PPgjUAuUeAqg/cKRwcUaGZkRD3QxA+0rZxEy4YGem4C3AIkylZLX
ZthWdg15jVDic0CIUozWgYu4qB9pXeK0I66E9LaoYJH7PyD0LS328JbORfLRVLsQ
yNn051FE1CIYUZB79F9HEw0k5HYXSWI0N0UhjFe7jMnaXp1HWRlROBn8DZrU5qAh
2A9S66JNHS2dtSEqqaUj4RMhDNuvswAAugUSJFUrXqyQZyh3z4HpT2F4QiwMUASa
RDwJ9o83CR8BQgl/YhEjPOKj8Hlmh2g6dnOBzCSwXvrVOgkc4vQ4MMJHea+4FkSb
sDfIPNWdPK3RzQWyEgR2pRyy5JvzHQ+7d2mOvRJVgABS+I32V4DwsIxHMPmb2KBl
ven7LMZhPPgSeE9e0GIUlDl467rM7KtPnKKtLxYQWKv1MWP7XWvz3FItUiZpLOr5
5q8Q3CjOjSiO7bDoPQOBQxG+XWCWMIFT5hdQBbETxubzdoxu2wjxbAUZ6X/4F5k2
D96uwlOme1Y3XD5tSIEt9ayuwO9kSnE6a6udfP9PsnIu5D6tKdsU6r3QcsIt6vWG
noaQgPDOewD0ytsSSd3ZgEMMuB0+3TQhLUNkmfHRuA5kKKQtdTjpOJ0p3HK0/iB3
5t9f+JQ3d/DzuJx3HXDuq8gIiC62KQNAvyv8W9CFTMYHpbKvs3tQOHypsRn6wNek
o1IKwYkoZrzRxRxy6F/bHqUaEX4BHF7JLrrtna2fVqymGTsdZVLnx3J0rgdWLubm
UEFh9Nh2Lxa0X4m2ApLNFdiCgUncILz8Y8VC/qSNiLOQ4iW3vBCZyxB1IU3fW1bX
393HLMeQoHFMmH2/q00lyX3dkZ2aHvfSlBlgFCZ63qtRPeSNyuTDaMF4+wafTgPa
P+n2PdUFh5iIfEJEAKNqcMiOnG4FGSecaYAqYAUpEW3GYVth3LIpVHv2bO1qgtjI
Sxw9CSSMzi9fZDJWT5L0Dgt4v0muiiXKjCctpZA1Mpn6snK5ABR8UVPLyxuPoHXO
zBQhwLOUtVbOHdBRBcI4ONyMoNyPwv8ElvwsVOhDKIHHf5TD+nkzj4WIJctjtm4N
bwH9gEdcw2q9gw6Z//csr135MV/WR36LcFA/dSql8YQajU/bGKtIi4XMMLzbYqtO
x0Yh5iYoEJ0C3aN0YR2sP6kX8cUIwVN2YMl9R/Wd8EaJfqGfPECxMtf/xb733Qtd
g3+8N4SHB2XGmaIhyARUkMcor3OWkbYRIL1BRonDqhk9+VY2ffrBNxMfK81gG19p
GStl+M+RKHLki0OM5W8lhlSIN6OjiJEuqQjAzC8ZUtM/oQamfF4mGRe+oWrrC3Ou
zlXcvg5zMUuSj4G+1potK53dON4aTpePqn1JR//KohxP8wObfUp3aUa9sQ9UqH6l
SQxdSxjc0b81VyN+Zrdyx2t2Nz5V/A7MDYxBTZp8H7KwbskR2u7nWM66jNNqwGl5
7mu2SFygbW6gG/LJfgsxT5tKyvaI7mswq8KvbSpGeOFTrym8HgdyAcEbe/vDUJS1
+MdAo3uikVZwJO40eKpXduA7isYMdjwSeyPw056zZ8gq1sqL5W3r8mdqEhO88no+
o5LBEJC7Mnu7rRDdpNJ+Qgy0sYAZdgSxZ4ysF6KxWCW/HOsctasa1smKeLwvM5YA
bnKH+vpsqR/lt5gMFgT38oXxxU0fwNmItSXqbfoBKKEwCCe4BwUcdKqOWPJbz9AL
fHgiAhYkUUE8e9RGAdOSD4JrV55zPdgPIeQPnhLPfFY7EzIUZIlusaBtLb4Suywf
pb5yt2LJmB6aWnwh7gLy6DVCLJkw2liOENYIMP02CzveFqcvKsw0LbUSTipF3uPq
xqfckfeqRffSyH1CuTtVEE7acpnX9P0WqsKhiq5CHgjXCuLSA9RO87PH8kWVYDJd
7KSI02seQglMJC51PZrqwSUHcASsS0rKrsTv6dlL4br3xWpwnJaD33KPQ+0x/yfP
zjej9Au2UaBHX67NuPNbf9ebahINIKun6PlIhU31Vchjc0xkxfeXCBAFeFo0syqj
w+pIzxB6yymzMNv73QURLU2uRE41PsPs9A/j2c+/tysdeB0Gk7x/w8wgltKTvBrI
dKB+uKiI1Fr+G3iNRcXWXCmoHyRcmkqyDwrgHCA3NYlzzTEexgT+3fK7ltigQdT5
UoTBN2HhxLNeEmynrY4dno48fIwBbbhsEaeTGMI3xCX4AgpmTz1dSufz9x3yhQnv
Brmj4pVS/DcNrY4ORiUneBjpDvo23aRZPKe2YeZErvTjDKKRNHFLdlakTqjWZa5h
wqVFE3RLZ+svzhluauZdX8K5DMo2CIQvBT5diodu+kD3Al2Dk94wIkz1P4CW+KMJ
8J+Kqiqh44tQMLGf7JcMRA7RCK4q2O8O4wJsQessTfCQ88iRwmnZ/xm+Sok+AGiR
I+GTcSKk55S9W8w6GgVybTQWhABXY4x86/x3b/sXQUi6hSngJdBHCT3dAOzlcolA
vtvZe43IdyZ1E6hEjH724Y1mYT5ux//JTlE0PkeIn/qDadpNlKsog92Ke2YSqFyH
pr/szMTsTrXSWOTceDK4AdZUeb6s0VCxVDOVulcpX8wkKLgG5zKn4vdsFM2+9457
tzvCSUySKRjnOBTW5lpZTZjKwrV2LVcG1mnUdQ5zJ+ayAaoFY9RTohd/GIPGHLP2
hYTzP/2QUZLyMlclwb2F57amctxSr8XB0Hg/woij0Lilfn3p+uUYJJpY5/TsXCOL
fk1/1a7F+azvHEdFjPoh3rosPpM5KbvH3TUoe4pUc3EWilXPyXiRIOzk5AvytcJt
wqSpKnhhIzTVh4AKl8NhqtWF4JtBtwoF8UPHUAtGGsm2U9XBbfV4+A0kamUf06Ci
m6SuPEYJQ8zG5aQbPjp5aSiB6bVVSy+tD1meLceRdejkf9wGy5aJMFj4G9zOTnre
xZKW0lvwSMzBHpqbVVdz4+C3k74bQpFnrlvXObTrBfK7UEEE2zAAHbKWcyjYZrgb
9VH1HPMbxl2jMlbGSfO1vLzAwshM0qv7hmerq9RTaCYNgpohoAbYaRSYEZHpJfx8
nBxkjo2Pgp3cuJ8jWBWwHojMyoRtWwLH9mkX7mNGapeoOlNNgr4gLtfZtqMlup8S
NPVU1lh65OuFWxu31nPaU2AsJ4MXloFpN6fHAvA1dOODo++0UwiygOAt+vsqLi2N
2h0AkFcBBnmpAHvg2YC/VLXzscfOmf8aaZ3DdoXx6U+XA2P9mCnu/b0g+455xPaW
cNqbTMI28M4RwOr6ouv6y8alGEPXIrAvc0NdbvCpPxbxkUt0CRyxrBtDU614IuFc
IKBqeoVUULoMulcynGMw5tkhTLegtxwLnQ/9eYu9Ib6tNRv8KsjUrGUES7Cc5Rax
Gm3iwjnAMZG/bjCPAErAuV1EwM/06ezInT0/gHlbNenA6uAj+stVmSwGg8S4B30s
bzhRhLW4++HktYamcNRefNk2IZ9jtowC8b/+yZ6b/tbm0LxcyuMRtPyE9Tvh3yAm
tgpSYoIje5o7MFdpENqTsSbmd6nRjZRyiNyqRcscihvRMFJ43XEo1kt2vfPcjgCN
Dy2+IVdcnRD2Spn1DackYUzQing2XAUgGVeaNA4gMrSpieleR/1mzV3Lkbs65meT
QZJwGspxcr31WhZ2SINAFR1C103CgZ+LlT1j/o+Gd+JDS6NHZv/I39Saj9jXJRRP
8bAV2npYQjZK8jVKDDzUlcPC+m12mW9Sna7tT0FEcAZvlbc3q611d6WVGplZZCO9
Cl0gzEWyRn0bNx5ok/TaUtOzjGAIRlp6uvqIxwNmbn6kaBvyMeafsZpZUFO0ekFI
nFGmqpq3KTmTT+q3yuUsipY4BJWlgkdvtG4f8z+ad2MxLk/1Sjm5Fos7hLmzJWIU
JrUzbYY90z0UTgcaOoNGXFADV4dDHhvo1ZmWVls7EIdklPPGJd1i+iKKWa1vLA2J
i/ANErW7ZWOtJZOi6rioAsP9ZNDBsQsm2yRpB+HJR+QkxfEcidkw2fasF17qeUE+
10qNylnooB2LBrwTkEhzCi7bYeIzif9QBHluJJn4rro2xwW2rUKSd97VvqqOWTpw
nFu84r5ibYZwUCBzFGArrFnjpbeSY390B0fFYjV9OxyLUCsI70UNOJPgecOZO87k
Ssm3i9pkRIj9ApV+Xt82fTcXZP0FIqgh8zw7yEnR0qIjKVvqbWEKOXigbK4qwOlE
p80V7meZLESpCEMNifpWCvzevBYjE9F5ad7N7LNPwBFGX6yTjCrE9XX1XJOhiP6h
tK0llfm9qiQLH1EFFr8hHaiC8bQIjmWmSkGSD4xsiG2toSaV/XSMikWp6GQdRr5t
P9hw/Q1z9G5Obxn/s2bC6huiaYK7cf6ln3u4OZIK5P4bnZWn8Y4yYSwk4uDGK3Py
dA0YjOCj9mtRIhvN6y9/2xIeFEBcA1ZFdsZfhpp7jXF14oVgodkApj93EOvJ6AC2
dUO1Tx4YpT9jawwzlDS/EUvLpyfxe0rkfEF33yEZFfoit2iaZ3ODKu4FhK3kbS7L
0tTX477OZ7gWVUaNSoAOpSlDXl18cX9Z3RVdlQZ86qNfqlxCm2e5UMT/ZEs+eUuV
EHoM17dFrG3fisKXCW0HVrwvBRwNOPZlxE9ap4QjMCBElFc44Rcrzr8FViGvM/4X
7ODJgJizVEJ++2vFdJ4s2G9wRGMuxRQwKEN8ZqMScsLE+/qmJWijv6nTbmFMKhGt
FT0LIFZzbvnxKuaSnfEhU3o0QJEql/793yNFIsI2UeFjKCiTkIIQkCcOvj7ewVq8
Wm9L/4UChtfgWHt0inxjnpfZGjmoP5laF1hI08+n00CKhi3gkFZqnNhTgVB2PcWO
VJ+/Xsjunz3d6Dt0i2/CTyMtLsK82/J/erZt9FFWj+7PVZDeLOPqDMD7aFFUZ8iV
5qaC6B+9lx0TnfG8+KH53HLZ7xH3MsNqNAaUQexK/E9W2QoxUUd04rkvwfVFjnJN
DWQ5PLQyKZCShVohDgXnfNTf5ZP8JbTe60LQV20FVAqt7hHo1D9KpUUKB09lfdfq
T6/Rp2gNUmL8x1TbBr9H1jy2jtgd9RgkT8MOHRmXSJu+JMJBUgTICYD0oeF+HOOK
RXB2fpOFrGX+XQjFINFCM+3zF3BB7F7WbH6OMf1a2kfsBhdKnAIJarA9MY/3tJVu
F4Zu+Mto5Rnz7xAesKpPYMyZGjHvwwdtbyEgHPZ8A95BKfp32rH8RWGPJt5Uuk8r
kZkEaMRs0Y27mtrEUJ1S9hu15yEQC+GgYyMHGhmNsR0Zb/2esSamQ9BsTEj58Yqf
IbM53uJJJhHlhzwKiVRDleb8ohePwSAhY2PO5/nVAxe/7CfEuiTSfFmNa+4ho2l7
hvUe4nR7WjyLxI71OFzlPYYR3q12nqLSfKBPwiaOscMFVBc4mROXMYPyo5Zbbk5Z
m1Vln+WQtAd2QlIjheCsSYyrDca+yC7EXTWl7kz8J5KkgQE6eH+D3SSmaVQfbjTZ
dehdSWvl4dQun4YTqjMmNfzjWK0aE9Tj1V23QW6LaPKjOMI9fInq5nZCgGOwq6P8
r7hhUXt9sOufbL8bjknRRWpMJdjlHYjxUgfC5RqY/JJmTQtA9tQtkzzn0HOQoVL1
7AZmJ6VSyx7k4oYO/5uMR3J34JCeinhIQtwshWDNrNckFwPw5kz55Pfaqj2Q78Sl
JPWDpItySKi/ZS3Nn8DRiPXQZIEhmcjvV/ESTXorMKjtRogxb4iTgF+80MeF3xG3
6d+xBfMVH7qENn44LImgQ/ZUiFxsUHAXa3M6+OzIpWtlxxgx/XePmACIAj9b7s2A
fo17ZPHfQj6EPIT6VMBBr06/ZTjPt+12orTV5Q+vRYndqcbQc39gPagl82Jrs13a
JXt+0/S1ja+Z3kH/sxBWrmPN+M23lty69dTg3zMI7U3QULJSnSUjRA+Lw8CBarJG
8fVOIKlL72OIEvWt6GuU2aQGVwBGYx96yksOG6hTNkzwz6qM0Ahdcc58BDjE3M8T
0zwnADDN9WnpZQFf75FwWNRllOzzDFKzqIzeSH3e3MhRAKPjJIrjK9N2H2OjMx6p
r4vCfQQS9dxgITaedCoBhqx5c4pd02WPn6+xUlS6D+P5gZB1g21vXHbh3tu5dAul
gFVhKmyHwyK8bvWXH0uEfQYxkTO/KjFjnM/IzIGGCwWkmNvAhdaZ+Nb5GG3JeKmG
XfIZgAAT95O+qDxxO8A8BmtXhhke4IXuBT3mrsf0U86HRxEbFxTVzGpIRp0W5duY
FhMUAdTvLtrvtOYs5jG3crIcJ13WEV31RrBh5AC9MmSYCJoLF+NU7T2rL19AUBiC
wQXwi9FDhsGQ0aKU9DnfZFpqViOmfM56v/siUNDSySOZu3T7HWiJeNf5smpmnDDY
aSD2UcxQgS0jofcrg5nYiYtKb0nhdkGdjF7NSq0KEzfl182IW5ejrYOGeUhvlsup
CkloCzljoo8nbN3P1cNdwFkYiU+vXdVP0/MWaOKrgafEVQccJTl2Meq0uc+knz10
BYfeqp4m+P1suJseR5TeFO32gxptoUVMXHycEWyqc/GjPIxsN490G4BDxNTL0Wpd
HSKXNVKakJ3nVE4xrPLrKekT7myck4d8aaQTjQmo6YDE1vqX51mUZBocK7Yw/enr
61ln2ZW/R/MsTva5jx2EQDV5SVfmlV1oz5xBf+RqpImaVICKBpv9/0WzHeqfgZHT
q1GrZ0miQjXUyijWshVZ1vlZPmMuw/85sUxN+ss8oLDK+UQwc4Xnq2wrdFA6URvz
180g1WN1AkiBX8Cvd0oFMz29DLugzYG2J/+FcxcLNo1qOlEwkT0i5Nvn3uihwRlP
fMLajqVjghxVaBal0uQUrxXyTnmrzuPuzah9faN2pFJLbt9Hi3FNgXWjQBoYNEPm
smZqmtTrQKD2bjoeKtG4+G10yqfRrFmAPDEuj2btWGtEJSK3mlA6wDQKJwdXNDT9
7eRVuMEY2mO6jSgm1V+fIrucxjTrndjD4Vgf0ECj+9+SZUI9OvHdqlleWkwGMDLJ
1Jk6AP/8NfQV48698tz96RCejQgW5SHwpPktWecS4frypdTASq/cu86mOmttZvf/
YWnG60HjjywFtISWIvmmDHn2MtlDd8XgEl/7IyXwREW+7LyNPBrPSCKwhI74ztDZ
WUSn8VLPeH+IhkEd3/ZIfR6mmlO2/KUXx4pNL8QtcidEK18oxqQzDfbdsWGi1b8S
m47DXwmJBpIMpvg16K5Bz9V/5jt5lmiQze6uNYyakBkgxO6oE3ScOkxoEr2jMj8h
EoFGwlGBtv9MW5peKzA4u8ivIFrZhOwI9vfyoF+d/wlXXSX5nWTi+e3B8Sk1uM50
6P2RpnBMohlA8Bh67FvRa7HyeW1yjW3/9IzQjqzu1PPAPaAqw89Ksw+jolDhXixf
UU5bmlhhbnR+wlplXsv4P2SXiZcLs0ZB8qEkrTBwAmcgaJEAiTQRuoh4hgUU0X/n
fOMOYhVn+7H/QDXL1nplGRNSWTG01PtQ92UpSibN3HHqd+dOFCFk+j+obz1P/FZ1
nsiqy746YohaOBzvoeP83oXM27+af7HtKqJj0oojUCDjHexgHpkbIomEVYzFPUFU
6+kOwA+k6HGE89AYcX+PownN1jGlP9Dzkg5AOKFfgxdfCHNrfEmbsKIeQYoE12KT
n2xzfP5RCva3V19m3Y8/fuuRI+YdSsMjCFVtKe4yBSNXJjTS03HgbQ+nPq9uonS/
eDtfNxQXnkfrNNRRzet+GWtskLkUbVboTwp1iGVmAEj1PJFLjQ4JhreC42x6vLe6
Uq6RHbpQ/vXpnL5oXYNHp3+jXmm72nKAVMjL/3u32l1LgyrB9yCiVnW5zKHAECzC
0XPawT+q48eBF0AerVqrrFnx0rv40befbagg0eLEIMJQjLN6J13ckC1wB1X+KYb5
GBSNQh0Ob9wbtmzFh9aQdAtRPmoKdvb1Mh0WdqFB99KaxndrOa9S2u1v+oVaPrb/
5S83wTSImUADFkrWOkJ2/vo/LV4j0t5WXaNPUdJ4qqY8JbQ4bggsTW+j1vOyCUkN
OTiAyVKX/+HPcAVuyJ6GIdbOdQqP0aJOmJ9DHLTN6pyrikuYjkIe/o4+QKy2gugN
GUJ4WtTxNQTzM37glN2Sp1r7BsgCxoDUgDSQ5vVbu7qa3Dy62I1tkifsaN2YRpyJ
9d7bz0C9lcppZb8eNEgNka4SGz/UVHQgcNHcO6XVNQ2Jl448716va9hEhjqBYLTu
YdYV2uFRwNF1TVwIpJ1XnihrlX1nXtF5e90+jo1lJsZgt6odty4rCb3f0B2ReGQi
spFQvEyFec+J6Wu5lw+A/mrYOY4wWn4Z1hXyFjXSTMUm6j+PtN0K0QQdHusex04w
4mK7i8NcACEH2JOeQ2cGyE7jGyy9aBzfZo5YLppok5e2OIDPvlI3xfhClruWa7Yy
brikQmXdh38QXK13Xa56Ul0lxpMst5YnQC8qn5hSHApzUHVIuVa/P2TmlpdHWocY
TQ9SRUO4OYxOl1iPemExfcBv47Kq0bipyTUTSohyrIRw/GBWdj5KNMpuTDlQ551X
CwVk9lbeY52vIXFIrZHP2VV7DHRojknxtHUebDlBGgqnnwBQYSkqSqbdUOKUJRpp
dfYxJULxaCs5zqiGRo5RQ92m6wpwRsqa6yNbmW+w5t+CpeQbTv0yZNd/qTOBkrsV
X1G8sH0CisRQyY2EtQ6q8IsGeudwrc/tNPF3SQ2Q7eU/AwInnGAySeKqp8Wg9uV5
2Wj69y0tzjzZ6O9iPL+nJchkGOTfa8yBf+0fA3J/O05XnrKmmWaDORO14jZDMJ76
Iwh/Yg+Hllp7gKmu8Zq0pI07cZqEO8h5zGK8VNrNZr4BdtttCE5j2bHaDtPXVQio
ffHl+zFmks6cLnOAQKmdajHQ5MqguxfkUab6lfZUE4rYLtnZ9zGzFXBwR/8NpkFH
hLAyOUfw2H8mOcLAZFU/3y/YL1wTmpxK18MwU5i3ikays/MuNA2JhtjhmMahl8tq
Kh5P7lJ7pP+zTRdeRGfXW7ZkRk4Wa6KVdeqgeH6MbRDR3NmnnyH0GtmmE/JUdP5j
bp46Oe039oyrfBBnhn6BdnjfGIO7B7SHYZPbb8oIicRbEHcHVQ2ReLznW0g98RhS
Q3ERnr6dtxb+nEkpZM+lxBT3Od7KYF6Xx4AgT69kDfpNuCT4PLcsYQ3m869DVMFK
Wv0DdD3xF+Art43d4Tt9zmZj7sUXX9aorkZV+djXOlHAXohXPA/TTBfkpTZll/Hp
nGJy2l3ro0UCvb3dC1NAeXc6h36yYM/wNnqLcvO8Fz5otwdxX7xRcrj7pN8gG/nI
kP7JJKLrJukirrAEVC0tS8YxjEto1yUOU46bdJyKFCRxwQitsYYSu06/D4vD/0/h
q+/THJWRTk1/50bnioZWE7DZaTwrwg+zS1dP17IS/iO2FLma7eu1p1Dy4b6CCg8A
5ZgPfZUSiJ6oFdbmQDewQCQvxoMn7jnEdc0ka0EOQBIBNLfGJK9fJcv1Kia7chD7
adsRIUWRDVtvWjqUFJE80ted5ayM/hsWJjmwrRpA4APJIeTnVCHH8mIVMrGum1Vq
SW3Mp/+yow8eguetEV+zlhhQwG87rD5FKPGtM5T5VTcYrcZw424AygUPW12Vcoz6
6kaxr5DV0+5oXjK/ufghAt7bjtrMGyQ8TFMzEddEAwZRxWfSkEvZSKsUcwPTslbQ
vzT56Go9j90N+kK9MVGjuoGnluQaxu1eyES/M9HUWNrw5Ft8FXCnAtMcDRF1uGx+
GiahXQYpEM2CLtuuvYP0P+R5DZRP0AYkc6KxuW3jB6zhrcBZrIXCfMo7mS7ug/Hf
uysq4xMfbauouCwkej+XD8BE0g+fklqHMHm/+WiYTZwPPmZSdo/LKxan3dsahJ3d
USZMFViyF6QbgBjLTuhMAC/cTFNnbrME7XLLAUvWHF7Th4UP+8ssvMn5ymBPYGIb
SqCKJpFnMroDtAh6Mn6oiKh0SQqwPYwqCaBR+x6neYm/bF8MYnHJ7gdAG1U65Mex
pzlByOP0kA3NgiWgZbXERbqifhSbJfQxorpPiH0yyk+2AgLVvzBON3ZC3xH914kS
gn0Ln0gPvAZYuPPPpLhpG4gxzvgoqSOtUoLkiyBbzW/6mCB5Mfwd0jCLD2+4P+J5
e/qGjcaSZGc2OSym+xUspzmE77dJti3pQrB8qaODjuaOzqCrTm8wrohcb3yzn77Z
KKJDF/x/PUoavI3zD57zB/gyK58Xv4RbHLjogFQlbAtO43ulbddXvL25O/C8vu01
aDDDbwCO/lWDry4NLLqJc6/d5ikX7pqdUqmcfm3VeafPF9/yv5a85z06hWd0DyWS
e+N2vOkYvl4dHHSt2nWzfwgU9KbeGlI6mtQSLW0g4qvuBABvUW2CCoVBMoWB6aCj
bht+GAjhb3JcVJ/2hAE7m4IidgreCPdTliNNEHmqlMM8gV+eKwwo7g+j+3lBQmR2
8hZIY8/NUQAw2s/0dGm/eSTaj61mu7izeLiPyWCDANWZOzAtOrjnna0ll6pj8ktR
7dXOF/ooxA9oRVE5plP2hzKFeUtGEipaR0tSCUYnwWvJ3GzBUBlQ+4wKguhNc3PN
o6k/BNO7mXcbRC7/Fkeon6j85oa1kJ5CgRPEXjihte5+hxaJ5fkupuQDf3gdf5uy
csblft5zNhxGj1ngkMPn7hBtp2uqd5Kk9kJSFLHcg5N5drcOCaqkfeuZS2LqNuR7
8Rvyxh342WYlMKxbIyWwwT3YlCk8IWdrK/N0s7aCnT/OchPxrK0y7PqXh8e86Xo0
opFabE1IyV2GVCvBsJLd6+rFiCSijxmN+nRDx5RTonpmD3auYy7zEZul8E0SD4KT
aua/tASuLe/7VFRxGBngHHs2v7YMzNaR2casIpxF/BybSjWcNHjdtdoPrL+r3SLB
qxjrVG0wu32pvuKwlYrjMvj96eB7m6i5STka/2TIBA8Z3QpJrsX/S/9BH3b0rBoi
SgrZB2mrjKLHvQESSLioC9I6D3Ho0JKOXmbaPkUdIYtZKbsAflKkVaUfzUMK5xFG
nftwugjJ4+JTpta7kKifnjiL6FDSKhMqOEir3qJjO86o1eqT05CGJTmKezRtHDVB
SZCWI4a2qMIXAe0XABOSRoQrjAT7LLO56NwEo4s9/dMwm3vC2FXROVQSztGB7i5B
//QeSZ4thkhJl8eIvpsNTP/RmI+odRLKOOpNVl9dgYHZYtdXUyWPsIBbqIXlFMrE
tenGYzE8d1xKuXAq4PgjaLEzFvgakDRLzEgoToQ3oGJL8PCqWPaereqsmTZrLAvT
htA8gUS0asR7IqRHssKIfRfS2/lQaYG/QkJ00m/SuBKPYvsa1Gmb9OqHQJt4eoQw
IN73QfeQyhNYxD6+bGdEYU2Jfj7GUaI8pDX49x6Npmi7NPnUwT1R3NE+cI+oc9J9
GbrHDaBJashpZmQFXOt0Xb1YoR6kVnCtXfhi6oILT90gkITFErAJJTEALDf8dPH7
1jRm3UPmOnwW6k42P7LfE3NaXAoIlmxHHzU56HInr9qhVioNHqaLiisFfZ1M02CJ
Wm4xghscoVEcIxzJQT4ukD9i4cB7bgWLcLU2p8kVI5DWcv/jKTF0hKcTKiRqdBJY
iNdlsUd1nzeM8N7keD1Ilx3P2JUK/p68MUov/ekTj4CF8rr94pdgfnWLpk9My663
8YWGvSv8EjxSL/pi6uYoSSIUNA+fUeTr5t2c9grimbXBWgMpyss3GwPMuKhhi8pO
0MNgNp/7p2N1midAM6BiFVlRXpoScQXm0o2WMABhxpDfBxuLaIy2nNGhiatWkcAh
GzvETIYaZs+0h9eqQUOlwlRIJiboBHfxpbyPrtFRqbdNtblahkT2C5Somaaz9hr2
D0i9He+Jtag55TOw7jP37lErCIaB7oP1m0VVqVkNj3iLn2ZwDYWx1UT58zn7AyLK
asxw3ZqPsGAxipHiIoXOjHQMCSwC6PKLI1wTiX9dg31lQkEunlplmLKmfruo9wa1
jjfuW4JL36oNOsNtAA8+sgK3/NICHH0uZpy0vm3Xi8X1XMWPwKU+FLWAg8EAXNes
WXgMI+aFHpLqz8uWBbFTUaWlU4ZRCCSy3+N5d3j4CArQeVCaV28NoIdSjp9hRU2K
tG1Sv5MzHsLx8CsB67PpTldRNpHaDnXmae6iypk89E6iyGKFGXFe9wpcGeeOOqdT
WESZQQJhwVfxRbcBlzt+5yieUhAhCBU3hhUN/aOcpgXeIZ3dJQmQ84zpynOQ3FLn
ILlXdQ8YRCuXiKLPzG7PpUQBDwg+fIdfWROWY+9Q2EruABLUSO/JLecTvXMxC51i
p4zzyzbWVmPU+lqufCeELwXBLfqqkclBbbb3NpSynyR1WDnl6yBb4VPzgocN8LBr
Uk2TOkRFgxLLU2kyv4SY7C9eTYZWULdNdqq/hvEU/It6uflqKqhjYGJmD8X9riYz
0auCexRfaK14rmwzyLxRlStrcFJglCuT8+U9QTA5+IV5ktvwyJpwQukdH9lPnm7M
aG2cZqBcWYMOz6fOHbp5reJvY5M+U6AC9SiXQ8YFe2BEhmOYopKX6qPX5Lt46bNE
/4+bP08vw4zZP8sQ9v1uUHqZApduEj4qE3bcQGaADTtIOjbKWppkIGtev7q2bdS/
EyExHHgvJyqpJ93Emu4+IdfReakZOhnF/jB+9VgLI7zfj1q51lGSj4r5T1L2Ylow
AOJvhsxxq5T7+k63i4CH63bDBlrDmDTj+Ii/qxSprCJ710WLJ2zcrPLofdI/5CF5
dXR8Yy8tiaTqBybWFP2sOyy66b2W5a6ygTYuCYk/mg4Eqet4W6tIZwkqUpu8yxsl
+6TZOWfGu5VYf8BkWvkJPFn0OctogfJSlAUllMOUQ6LLnyV9Y5QVnDpNCNjaCCFu
azYkaiRTr3aO90dQjcgYljfts/sVRhf827BiOicd3owAQTTWrzC3onr5O5CakG0Q
gHhtzqxNOu2nOZQ5C5q8yw+FWNzL3WOm6xEN2gPEmzWpNrr8BD1jB2BR0lujSYtH
b8yc8q2qr//pJbfpEkEQs8UgXY3MaQ5OfdXT5CzXqrzc+LJ3lWFYBs+Up078UOZc
3f7NyZEXPUcX/6FTlAXjYh+YT34IxYueAkT8fIhQ6vACabWPgG4pec40N/PB/2bq
ViFCAuqI8E0zFSeBcMCaA2gZ0veXRLc99yxwriSWt9txkdmJjiO4FVS1OxYojLbP
+LNvVq+01NQxNsmYpfmhi3C7UIcK3pGuyIaO/YuId2qVKO24DhMvh+HZhZwBxh9c
SIub7Di/WjY5mxdQgNf4GLtTYmPbGq5DGEk1GPkrYyLXNmhD8yMqGtoCIFk8c8HH
R90q4pqftkVhF6GhV7n4itBpLFooVJP8ei5lXqSfZ7FDziduuKzolX3fy0cdAZic
EUAiFTd7U24BTPoc76Yo6dbh1nqGDQveSXeZ4PZ/Jf6vv1XbzHei9RJpnHtTlOVt
mMKxU678wtLxTZt4718LUUES8fBjLodquyzEkstQ4qkvY0xOLU1sBe3cH1z1A2RX
rKGDp7OLk7piQy9Bpud1B4pfOMhlMT2bpbGWo5P6y+GoE+HvWKGXn3eCZHbu8Vt3
IWktJTVrjZDJrxEzL70vkVOSw0rGPhVjV/q/rEntB+Lqz/VIOppMkTLhm6ufA/f4
ahqjG1T4aW5cYaqmpLi++MeKo/6s8NR60wqgaPkXxIJA/6Hce8Ngq6+mf8dOndih
wnmV6Fylrf3v0r9weNLaElIRs13wV1wMkkD9mgFRpeF5nz5BvmppYEbSWbwzJAyZ
r0H2afxZR21Emuj/fBVtfvWXWNVTkk4GhRvbWF/NxO2OU7AO99RjG+ac4tyevmfY
NFL/XHw2tvj5dpxVu7tsd/hkkNcnCZekS+DLqNP/3MTEzdCqxXERHFxrm+OeHICW
FzzgDUv+cFw2k+rnk/7Z9NwIo9NoltBzppbf1W4pw2dZQXYy28F3KW8FvGYCOLT2
sq3igzttdja8l1Au2pWldwMQUHPzcJNfwIEc9++JVO+PUXo6zaC2OMgqztsI/6Y1
E4AU97TvXTXAe91o1LqHoduEFtmrG4PdTF1lFW8g4LDDtyGm2Okg3hP2FyTQuKDY
CQmyfKslI6bMtOeDfRFoN610M6MCVo2Po6zgGcOV6/sVP82ddBBoZ0k/xHCf5sfd
6svUHJsvZ69vCG0r26tarSPBhoCxv9LwyjcPbeLm5HWFXN+bZyb5RaVg9TQYEjZw
E715G7lfUa+17ROOTTtgV8IBY/nJuV5ZGKO5OW00m5mNQSIqFWFcaazKl2XKMVQV
JiQrv5O7XgvrPYU7al0r2gcSpij4DItts7ajCRJWPuoEoLJJi7XEqROf6blPau4j
Q5j9Jjnh2T6ahklZDRhudze6Wu0STz30/gwUqlhze6IO/GbtpNFQL4eLFvZ0IyCu
wCJeawjXpN0zF+/Vre9h7+JRxdwSdNX9HqrfgdYJnmD4+1jmWaNNv9UY1O9hF6fL
hB5YetUDXF1BS8JM6jMlVnJr+UIyGSYRf1Tk8Y4TwGqWy/N2+WogdF9dtiEbVRy/
9UO29deksZavsr3aj7KvCE0Ycb/leLwMYzUmAOociIj5oZjeuWBeFhrs5iKDMSMI
QlXGCurkiO8KaSLgy5ROziGLeVqITooRBMUYa244JsnSHeLsQyccmLIUNSNxMUss
TdJ7pc1pwVvfC8yB3G9RgIz7cdbD7q6LLMAWtJRN7y1RYOU3CqxlT1Ff7lpOLeaR
0/IpXg/Zfq53+OxhJW5D/NaitHIUtcG9lDKh+DEkDA6Lz3q7ZtI4HR33PLhWTfed
QYi99AKCbIkn4hWaj4C8llmfeW5+25SoQxWmO13i501U+a+Dyqa7DT9bmP/6CDhH
M8RAaqtCLwRyWS0wbhDfs8IWsWw9PHWCsMZtmp6mcPkhimqxSpXGNzfJmCOlLdAp
fQL58RascEYgPUaJtdA67c7M0W3ssXw7iDG/xIxGy7kjWXFC2FwPv/qE/YQVJ+X7
DNYGWJh6bhG51Qd/mUI46OztS7vn0+GSw8i3/f3MQwrncg7QUhKuojh9K07Fjq4v
w4xYimCLDYHxcAvAdpxICgaPFSWpJlsxycuCgGInOEc1iPk5UV/LSoHNegGmKVji
BhGnSCoG9w5z7Z2DKncV+RQhGVO5BXmA5Oz30FOIxPg5kXQkRAi76W+A956MjSDd
6Y2rippxtAULHtC5u2CwADrzcOqg0nSvqalb+q3z9iwy0jIGbFP37bBAW51xexer
k2bWpM1RC2WpRY+NdHzeVcT0eQycmmihX9r+ETQ6FEhwFIiEwABp6yJnRwma3X96
bzGukIBCLWHfGxyz85W5rIEbddsOEE9a0qdUtA0pMpM9TyBd+HZJzLZ2X+anxaSj
d62zt+4D5YKPfvxQET6uwxcLayNAT5VQ3cm6wbE9gnEt52J2LHSLPvdewOhgNlnG
BQY3JhopNIwvNm0KbdOjHz4QwEZnQkdUi6mb6UZr29N9bGU445A/hsgufGnlWUVZ
s9b+tWiG5fpFrQtPT2SzoxFKAlAyVua1a5EJdma21TwGDA38j4a2mZwP7KQkYTKG
/C9pArtVIU+lJH7vV16U0aNNPCkcGyED+eIBY2yF57l48huYORXFr8eBmHh3JJf7
Yk8/H1SpXsOGQ8Ws/QuizMhkINGo86MYRm7XC5rdD4IjygZCdx5SdL9G9GhQadLc
S3FSVHsZAKgUJh7iMzuDGxWPZ+9LBDKry3SMq/7bYWPuPDWqvKnOJANYqQjBDLMd
+qrP3ySh8qC4NVEu3Gy9GzC6Qu32NRvHTJPoWm7p4lxSvpQKc2zAEln4qFkLCw8H
eK4YA6x8FgZBKk2TtnjtYf/C5u2gPUja3vXkzFRLscr7Q4zOgjJo/UhmX3s79ecN
tL9V/39TgxaLAG7oFSx4GPrPeD3aIak855NkPXMlGhcx7MF7TRNw8EWukSofz9zU
q8pjL4z16xurdaGqvBpmkcQ2Do2GLk/MYpXbgFwdPQcTbAMPmgukgCvx9Gf7IxU+
GxlmCwmF6KQpiRupSLSaURHpKCYG6O4WCdKwfb1wL7N1sqRJRGnwbPFQAN/U7Bau
yXAh8jmEFKotDx3IBhI0QjHf5eu8REzV+UtWrThoP8OWegj1pdnGl/WgMqqzVv5X
BE2M673+IVuFslJ9ZBJz2cIR9qBXQO/PPWrgVz69Tok5rW8kvCg7V8IlkRX1yQey
BS9jKON53YsnWaUPtZBpLSVcoA17vxB2ECXB6oLMe3A3t1vF8BND5uj0OMRVNO29
d3t3n5sQLKQ8QrbMbrQn1CLnEAJYgw/05EziXzAg88MpPNT/30irnOpaw8tn257P
GqU2toxKCoOMr5vcRE2kKw15bs0C++z2iZ2oV8q00pZXaZNHwxsY27dHHLRvRAlZ
qYHtKKhnnMJ//0CdP+jbsp1KaLbw/0rCrIxIB/uiPfLBEj31oykFPZ4hsv3wGLSH
XkIa6iYdWWvvmbqNh5zTP3bmrdHSGAviInMmBEiLoFmn8TzaRJ9W3aJ1LfNI9nYj
YMS1zfhnQB8RWikLpPiVrJ0XEvDi3U2DFQWos/lh83tH7AxiwN7odAwa6WZJiXTY
m4hUXUbcg7bKFiebaOFqjz1cYTxU55nsjgpZYJWW8Mc3HMvJI3u1V7mMJ200BdbP
z14c9xYbL+x5UVnLIYV2/YqbWWRkClbZ6zrvbAQnVn6SIVlK/LzZAE6hQ9zx/7kA
8STk+YpSDfbrAM86LIAqn0rGD+S29QNMPlqhg0To1OIWhfHmVwsq2rQ3C8npuNR5
abP6O3ohb6dELEYjd8MYI4O9iyb/O8SlmkeGnc1ft5X7R1ytrNlh7a5XaUPE7NSD
0FoDnwFK4run6ICa4AS4Ut2GojgXsRt3FszluBbjTvskGocKGU4wcKDfMJ6G43ph
6BbQixj8iTzoF257sWEGmHCNxgYXv61P2Rz007+YfpxbCzUhsId4L4jUF4LIgXNx
xNOblLgk0Kji/QV1dTlOFeUm5988oK1K1oAeQZ8RGsVqfHEw6cJ9bgxmXqvucJ2B
+gIkjOzY//FSb8xi2Hl94ha+XLWn6r6is3eTz1GmsincEhXiOfSET7eJW6uzl8x4
Q2FAlB/jSOZTvf0Ijge7C3gSm1H+5rZOSV+O2mo810q4AnkpE+hDkdZYS16Z6ZpA
nqP+lZ1kjAm5Uth1KsxAF+7OsbieUmoa3F6aZXqun00YfEVM2QnFsAL7gu5BdLOM
HQrsJ6rPaBf2eSRIuGL8A8Cp8j2aC1bEcGfWIZv4bi2T8etx/AcpQq1P45M0zHTv
Og+syriEy4uslUTTQ4KKIaYpmvQ9vzVSisqod/RUZvOXi23aI2r0s/zFYQVUr510
3XZoj924So5UgugKzrgrGzntH3dBYrjqG3GqZxub3mub8igIyYwgvqksA3b762Ie
YN0lgrk7pekbMnJoPevQf/4GT1nmmVyxTOINasN5y8LrdrdKj1UnI3DBKCe3QIu1
B3y8pchZPA1y7EF3YyemBIm5JuKm8zOYL+BSX4j1b4jKZ0a0PlREHQSz1p5x6OVh
/SccLHA2T9B82Nd0a6MGqipMcJjHhUI2Kiar9uBW2eXnkSB95MDPXziuyIZnVdnO
GQGq6ysVhyXBfvJNMCtcK6tgGYmk5ycJiYG4I1d7xZbRdNcXI0VIz/q/0b/wHBg1
FR5R3ALx1AKMgPs+lZy0ZZDEIS5WWWE0N+59dFynOTPLFD65O6mbSXf9M8V+6ChP
qhtsyGoIs/uroMb4CaqqzUmlhIWBWZaGdkDcMuvvyoWvBjPKluJQaEMNXauutlT+
IFVhbLP6NYdhhAON/F6iYPukI3eKx5MAyZ1kI7xk8VCrGScAruZs05E13sFgIw3S
MUEkOPqIvLmJgtVbQOoFd/zq41HYCn5ZRXW/klOFqf78oRi+p8o+q83gSS2qZgJT
k39rIX20JW4YtOVsA/Jjlp0fE9zZVxG6uiAF7wB0kzuXUbsem+0xYMRj96d16TUi
eVxV4G8oYJhgYbnBGlCVqRWbNaLl9zqC/vMneMdEvBqNCh0u+e8+O1kQNcX+0bOF
ZUsWTwGqyEhvs45jPCHZVcwdm/B0F/RmyMz0lu0waIXtVolUJ7C/uW6Iab4k5qt+
Gl3dhJgtiZWTDdhJpCpxsLXPZcu8qNz9cnGGxSK2oPIrHjNIXkGCAG8bSWydyRWz
8kzpE5P9nVQfwxU122GeWny/G1z6xCR6tyN5uTf6IqeBwN5AyAJzc5fmSKyPzBAe
7fJzKza1O5QemInePS2QGnFgx9n4MGAxeBCVjOvhpnLS/yZeiF9mzRhSILI8pPvd
y6ntcCgIiypuGvYYKq/aIR/MuT8+v4EjCSyGPht/MKp/9OmVuwkfq+6nGR/C2699
h5lPKBEvYi23KWgpGmMT3FRcg4+zByQEcACLCZJok9iAoxF9yUiP2ajqjkG4wcVb
yfPcEd66JJqv8oFAmsLrsFG1Cg4vhHp2WN2LQxt4/5Tu7qjSlZlLz3XheKXUweiZ
kD9nwjiX/yPM7hgl/slUiHPYf8AOhlHmS18byVg+XMkchc/h/uqYEkV8pNcUurnz
HiC3iENaV8yUOYvlxwMhJVkiFPe2ZIFZNk8Xrko1Zro3Rp+B+aCRRu3ldsOfPNn2
yR4CmxpWxPxl2x2xEszYWS+2btr4p+0cR0DUxYl+XsB2E4uO+2T4dAFxlNiV42OX
1kjinUKQILwQXyRPK41cXmUv/A9IsPFchsDBtzJkxmBbQjnuYBCvkJsmRUj2alB1
sQ4zGsFTZTe+uY333f9nEQqkGv/UoYWkiPgXlklsarBO9GVxowfh7SHl129mHQja
OP6qAHr5RTzx+hOJ1FSVgliOxJPepQRvyF8slwNyx0ci4fCUW+g1sYH7kl+feD/e
gruzDGg9fADlu62vj6M0V2uejP8UfEVe8jLKfba0n6wVJhXDk2HrZXiCGeSUYbTo
f+rz1S+AWLFT+hTIKjBNwhZdkhXmaveFzSaYT7fFjJJDfSP8DUgaisfpPRt9I947
OtGou4anBVjeBDjoK+GMMcIjOFOYEC5TeMVXmDO4hGkWQiX8d7CTqA00+Qp3SMpV
1Fy3ZlmKNDerbkuAwKTnRLj47uXOLrHyOhSjdNtxs211PpMyV2bcpZaaoUgw6Tu1
8WnSIcaXbDe7DeuTHX2+fN4z1e5ZdF2j/OcePk/mYJOE7+Q6PvFVwHu7V7brX16g
QEL5grj8j9cdqFN+OrYkQqEoJ6bNR10g+2WSh9Ub4b/hw1L6DolIFdy9c6I/e/rc
2Byb3nSV8I5TVtnYs0i+rVKYNQzaoc9mDMEGCt58cwWf+3iumPUOmmT3kPuVG38B
gA9gQrH5gonLVMiubL2rJbj3/mDRLqjJZKJ+7hZSrZ5670OTDaCT/ek7iVa8DM5F
iGp98cFLXQIZsZSY177uhmwbA22q0QTQ3fVXb99f32YJ552cBSe9AB/C4IuZIt2/
EcriTa1Owu2Il6bYvh5Wey/z6RFF3Opby2PefpU8kLJGKHd+PjoMaOCy1C3tZgYf
IyaYTalauQoDhihYe1r1ir+T594mSn43NE1xekVS1UgrxWyHW5S/tu1fk44jPQM/
9hNdy8plmWO4hCxfW/Lg5jspkh/vWti8RUFjtuAV42Tn0xnxT1zsse8yJFfEPCen
KSq5g5ai9nZsrJVs+GCtZkkW1dqZsjlZIzm3TnZ9gI7LU7CXWiqs5QX5MjjtSDa8
mEOlgbAaaOMqb2POZ4UvW7GkBIwoLFxjmp9Qlal0IEt6e/7J5QbSsq2qv/NlQ/0s
5oDy2P4g3fpIn+nqZIYg7aP0HoFzS69rp6Xo+tEhXjk4O4o3U6cHcIOD3XSyiATw
33KcEAY9g0KxRyFHeBc6ZpVemwIXSS4kHAR2Sln0RMcWJC5Ka+UU9I22F63tSTDL
7a2OvIDdplZPJC0G/u+n1qpAY0koESscqpW1+mRfIxUsQu0Y+jlSinvS0bNRCOID
4JCv+7eBeN56MXJ354UZmujIl7QHgBduzXBHTFFsrhfKg0baGY1XVn4o9IFPNgw/
TTaXAnn9rTZ7WuqpkxeOtynL5kRGPQbVwiBTnJssDTrKRuiRk8hpC0gpNKYuPDhe
t0IXS0CNsphBaxxEsy5uaM/2L4d3B3t2xl3+9FjTBqZU48m4k+qWdjTziQszLooi
tEYNb07uEujyVApbX7c50FHVc7lvzp+CuCCCNr7N0wZt2w0ulJzsFLmYgFX+BbLV
RN+u/HBx5TCxHHlrUWpLxeBhS+0UJKyTWxa8LP0C6sWHFvX7istOFv4pwXU30tU8
kVOpuan1oeP/7PHU93xtdR1HtgNPU2NCb/tbAl4y4upZ/x2VCjlieS9nouRvnjEm
hP9EzWOytRc3KsmY2cXHD5OsjNKBItwqUwWNga/7lVX5/GEh7SuCWwDRgBJ6/N59
hy4SmTsKBsupshK0gUNmFeJjdfy1WzBx0hVy30mZfLOT7Wg1gojxIL+7ZjJEFwyn
eMfBR19c9lLyJj6HO/lw1doJd/FNUQHOQAA4JB71oYdxU2Haw1kPBuzDFRYkCK5J
9blJkxAL0SgQZj6A1Kg7m6zKdt2yNUHGAWxNcAekUjF3p66qixnQaeFqzmoTKKo/
cS4VnPYfIBFTdt+lFtmCb/4nOpPscKPVifzUL0PXUG/00dq5VTw9Vi9Ka6uxAoA0
whMd3VKEDOUDjoo3eF6/EhaSD+CTJb35B+DEQv9RZZN3Qq4oAAmvga1lnDNRHOEh
zMdgiUMh66VpCFACRuhWRiuTF2lWHtpefooA1HpU5ha42qYLBO08+yeIGRRjRcGp
C8wXzicy+x6kNdPHQwgpj9RLke1u98Eg4eof68YmCQ+eaEaY5S8WiSGvD1QaprrE
s4dbqZoRr6hz2KB0OC8msjQ9CqqrDqaEZsNjjQLE4xNBrJxElvHR+fwTmRgq8EI4
ROLTdd34qpHr+jBLU2crKWMCcpKuW3Ah5dq7rAatvhPk4L0834pHr7uScHJe0v3A
cMrUuGSokp+A1NemJ6tNFwRdMgRamTdT/aZ+Bh0ZsBKVQTjXVIWGF8K9g+Itt0nm
XmDDxD59A5s20qOaMAY7ZP7hYvyDz0NqbVMKoZ7NrVxz7gnm7zWS8gwajILYHU/A
AvbiGhT2mo6porWbXL9TRBfVQbwG+lC7KoGuFKaaswQv9eGeJk15n0anR7E40bSm
qUaA+CEEth+13KWsuhHS5OtOMI9SuA/gqrSMXz3iYLpx23JxYsDQqJpTvhKB6kOL
/s1Y+Burt95vda3Pms9bTlXMdmfpPR72vy6aJuAsSGjsd8PO9ckkIWmP//i1IH4t
UWX37dcPaiTXiJmJFM1C1iqnxzjQl0drtYFKnitEhH3dE3ahiJvRGodWRuUcFy0j
E8iIqfF2o/2M0sP9r8TSGHJKtK/pcbVNck9Mv8LEhWDgCRaiT3iMca2vDMiNxMO3
K6tuDwMajr3lias+147+KWqWneg1tcKCCnYPc3srAmWHz8NFsVoXMaH6uE4xjemV
2WQsdQVlqluw6yY6TJpAdxrq51W4dT9rmypdl0EjWfakaQg2fiHH6NOLPHDjBwa8
K01JAyPph8bE8zKisS6OKTunpJ8QUm6PTOHXNZJrXhMvW0k9W2dz+cKq9Or2KeGo
lcETJxJOrab28lEKeP3mDeuN93KxZnPvATMRV75e8O7S6S86o3AbCWu99vdrnNqE
zNU7ByUAZoB+dRgY2kIl321qN7TAEPeisCyDUhTijnscnureyatzu9z64YAgYsIq
zdlf/aMp55xVdbeuK1JYSjQn6fTyUhmJ0uahGozygnezwv/PHV3v7QX2SaDo4u1B
vuTPY6XcAh8NAsRDhhOe/dDNFoaYVzWhls6+Wqq/WlKq2yv/8ZWnM7FSvarW15d9
l2DPZL9Muyp8CTlBQARquitVbGyAIZAb1jP0zacJx1mfNL9xhS+RZusqtZ2H8Ghn
TtTYU2jk+SJf82m1RZMGWp6kseOOXT83RGdkVCj/qOXHROCMDbECuu8FowfERClg
b8V//2SEyCIhqgyimgx+01QI8ywsy+ZV4xGjQz7ZtZ2IAsoH5RE+Alr7n+qVEgnB
+GZdun1ZxbrVeSUOyMruc+HGDEWHr6TwgNBxS4zQLfcOS0fjNP5fWBAjM+v+fK2I
YNG8fTQjxjPGpI9baOWw5+OHg9QOnzFB1zlH1fgtFHqb04IDgznWsGZ+G9QEZYCA
X/1/faUILTKZj6pa5rM4pSdzPEoe1BnRg+gql7r2b6tFezhNII68XedpzNcE1SNC
YpRZTiaJp84m1Lgy3zVD70d6nBs7PT8+NHh8wjCCCfHw8binwualad5IdmHckuA8
Tq8AqIxsTEFMZx6MQdvgaBLfO2z8rI8hz6VDLoxxopyCnmENp4fE5jzMp6zm1msi
CWV4xJNu2MFTSNzDHibyzzfCtj0ko84o7jSWeo9Fi0jlkm6K9Nh21pk0H4OwZcPU
RKpsZa0f5yGDdOJtYCQSi9fqdaPOtfKJ6izxi6O1yiOp8O0R1zE5HbYWtF+pXIJB
GXTJYi+OtoPJss/tzIK74ba2apqiyxyczKJTqW6E0QJixOxtrsnb1TV8cCjxcPBV
zVoxCOctP4zLI/Kn3CBXiVviUMirwiDldyuoz/7tcEQxgqfwvA4sgkVzm+hi+DVH
a50GrbUxR5/2o4SJ2PGyi+eazkd9JdmebyKQLQ8lSQMeWRiFykfDViiyMlQuKKdO
JyWMPM1KzeWMmiJhLDTfRX4S21qXqkwN2UlwkeBAix2hOKuxS9EvW6ToDiDwFImD
vakjx6epzCasmO3XsFj39LsM1tr3BC8HZDUlIDwHV6fmS/K4DX/vPODUdcfqJE8t
frBevwaHuFl/VDe6elnl2NSoxw7ORFzMsbZmbXTV8kHs0SGCHRLUT5Mgi06edT3v
t9B4gSyuAxhFJd9bNeSt34wg3c0a5Kys9lDAv3O+ZYW1ynMXzBgZXUhHd18FZbpJ
npPzByQy9VUdbC4NYI1vrVODEq6TcsKoKUeM+CS4N3XQWAbgS472gNCN4qfU6kxv
3EAqNF+hcEmor1LJ0CXIaaYA7c3nRiSydwJMSIWL7B4foCX9SWo7SCX0KG/k9gSR
MOs2bmDz+n/a3sR9vvRlkHeFNxq9bmWFJLqd9CU9IZ2ZcS+qRKiu273YYMsGCcjh
bauFaSPNxYPIp/YKYwHgAX9bb+XzGKauRZ7JWawYWiIWRVyZY77ZREVcBL0jY1ig
cDTJnhUFvO8bwo0qiIIFa5LNktem2l0Y562JkamkY9Ii8PtxJgX6UQluD9EMZsHP
EBqXLu0SNCoRKKu/tNDMcFlX+iE+YsYsDtCIZ2zTlxZr/bZYCGdfTHMz45+mlFEO
MPY2EpinOY9xfr3EsUW37MOvcPkrHieGQcgw47b7i0QqqN5KRQHsXgbwVF2NZE8N
ZImdmJuEgBNvP7QOX4TIbcJwAOJ0jQlnWPTAcqMvVvTIwhLlWT9TO9R2smj7H3Qo
TtVTwXpmeHCAIoOgdCW6PGvg84U8nv4wNvy0mOvA+zZcKWrgMSWKCGQxnxQVL9ne
SLRdg6sdVvYrRpo4Xiu/wGgbH0p2qTQ274MywjEzBCbqP+Sf+GUSHkXtInvHt4Qp
Ilew9vHkeJDfVxJbJkSH0peeNMws3ry2vyc+KdS6zjOkG5kBWCHhcL8crodO0W7M
lR4TwJwoohSUq4/MkKi2SbeKD3sqqMBWs/UJ98fwAk0SvWqozQuajvUT8P45Vmeu
iwgyk6y32BGM5khHoAeQiL8trJbDm8WeWJlB9WEexl3y3Em9dj2i4CgJnh2l5Okg
uR8U1BqbwQeN9BE9QhDKd+LSc7fw68lcVZAMu9pE5vrKgqTjvKLl5DHo/1hfzwXG
Vub+oCH8//AJzTy1urTxlzYVa2/ySJd7Ve2O4KiXsqmzXr95DdiJfnDqoSsL12Rb
LzuNcl6SlDUu7YYAMsjiD8wwN68P6F5+/Yz0p33MSJ1bBNi3FrhrrDFcc06/PD8e
U+RT0z5fE2+ZB1KfcfyjSolSBDn1oiiz3p0ue1Tg3FkZ/7ev2+xbrNg5Dttef0o7
ft7DVE3Zn8CfV38zDot307uJBWGH1l+L54oApDrYkIOAVivK0JFN+Kdxyg4683JD
iuSINc6y3HuJq9fsO7Mwg+vDB20EDo92ZMMG6CQamqwcCIUHDKDHijGjezh5CknP
8jF7FgCeHvcBe0awvckhbQLcJpV7+h9KKU6ISLCIwzm6V1cFkPiiHWjavqrs8jx1
fxvpUF6qUyUHvj3klARIbBeYbzRFRqIwAeF7Tvo5lGHPCVtlUzwQkxWGWlqSfbVr
8I1dau1NW7R44zLuDDMFBWozENdcrEofV+IfuiofETYDWah9/qqJbgv4arhM+ZIW
oR5hhrWxTDLwFLfKJ4+tbFG/XHQNap5CmPmKtl72ieMovuN9IDH4hMX9cM5Muuiw
mSCPbOpei5YlM8qJ/J9f3HxeXYbvMwI6ukctA++Cvzerf+jZctRHgqLNiLYR8TZT
S89K5L6xg+faU76ybmJ9V4BiF3R80pKc7QYzilQR2tbMcouBnXcjb5m8wJuH5CDV
m0hSgf6zoJWIqSrWhmu45XfcuBzNU98Fs0IChvBYC5nTqmJBPGeMzpIlv8+g3ZsT
kg9t828VDbEPRoiwheGY8Znhhu9mYFS+ARQhs3PpnfClPzwtB2CpQEt4XxI4lbw7
DHKLdsMcPl6lQ2bCvIfOwLCn3sLp8hT7FU9RgO89wpNV3fFYQSAyvXNOSjSXnNzD
XCNR/ccgD2df81GS7y0s/GbNjBUDNgaV0kuVxPv/1H1/y6UiUt6ZiCJRDLjQmhGC
i/Z4ctVozJ3Z6PlWw9cfWyOCXGaLTxSV6YbPZOW6LMA9Ixn4RjxjI9nF+WSYZbmi
dAs9MoDO+VW9+s8l0ZcEj4u62Rq7LurwlHbVdzKfQgiRwJev/bitutOLugKr9z4I
ci63T2P/sc6xyqOt0WpxvT6vr4gx1D7JcRZUePVWHg41vYg8lEZIJmBwLKGq7toq
Xf1xpnOCVUDn+IFzR6YBxZsRgz88sM4GULsIPlymQpxDEMcMQ9DdFCdui+VS0vnK
ORMbYgTaJtHJG5gLonvSW+4kIETDyvTeo8IX40PTGB5UYTM7+UX0R9kOB9vjtPbJ
k5ms3UIXMvAAFNTGRgmOPO9xcw6F7kvaOPWPYMP7KwnQfT+fVQJKL72/oH6opOjc
1Ez/yZkAhLIXWfyVIeocv6UGtBW3M6fIKgh4KJoJgKmZkn3ZgN584+4iB2vPkuy4
Ei9rmRDJEyDaNNU0bFTOinWFBiOxv8r6gQeqA7Y+BuBiHRs1hHW2F26qKXOkaKM8
UibSb+e6Qb0Drowx242eZpUIBBQXauz62rkqCcWd1vD2C7RMV/jXghsTKSAY0imx
ytE6mBOn0pNIl4e/99/KbiYayrWWOx3rXKYWtzxJLnvANe8enH6h181ENZU1TRUH
C/vke+P2fdEuIj/IPR00WuslRa+STgB9qYBzBC84rPgdeYqy1FT1f4sJHDIhEH3R
i0V4LGkXXrrRTShHrhLORXh++LZz11NrF3Wg7gibNFixSTGz/bTd+XmNkyJfBNMf
2tkQf1lDL+ElA7JHjGyUFstUhTkJYPUd5KEyQ1RnNbB8BSQmkyUQcK51dfJx6fFF
bY1iOBIWtf916NPXob726dfOJmRX0QxMn1KZI8FSJIJZU9Yj47+5FJHZiefp95ct
eM/CS1izb8xCYfbWFczmmySzV1j6zN1NPln4jpl53aqHLmupJ/LLuaark++Qc+0m
VAqsOWRnaVUY288yNiRniIr0O4AHEEB0rDYnpfonm3lni974t5vwoHv+UnZuzNE4
3oUNZ06mF3dwacKh3en8qH4iOC+bbTW6kfBWS6qTD6aGX5zoXOYPV+fNMG6CzfiJ
7s8aJ1a2XpKRonTQswd1gQEp2KHagpRyLPRDW1Q7jOsh0sJDpRbDlgpu2w7U+rgG
3TqalAshTUhoHPMKkab7U2Xxj+Ie1754oGHtPzqgZcw9sm5mBEDXGu3+dlw3DNdE
nVMTYDzGLMGm66jGCz5sWtWAjuQu9bdzToHJQ7YMW3xVQFBWoqABVBEQ3FSEay6N
sS3fzBgTTm6oKBYfrceb0iaO9EbAW2OkfOVvXX0XNhh0JtapUGQAajDSItJEct+w
LDf30ijonPjMgup09v8E2CAMfXKTmcrFCz+lSbwJXiJVf346sdG8Ca96cGQsGduB
sujRTf+gn/ED3A7F76NCwroHtFs+WMyl+kN75QJnM8ggwElnmj+LcquNUinJLDAE
l6xaWgGRbWcVaxDxRmI2Mpp5dVH+VOkjztcFoqqcLiy9aChy7u6ZNegqHOdTeEPD
Fa4nTT6abeUo08wB3LIXrQKPH74/PobuQSVSKr0QoTpKIQ1TXDfC7vuQUR5pi+BS
zHovhUNvebcg1qbYV8gwQxOnl9laePOm1dAU5fgyl/oUhMKYydyjHn8oeH1aTtEf
e2sCMp3Ekcj0N+Uv/ptTzbbZN01zQofc1xcwj1NBQ12jST91V/0DbkN7JRMECKrg
5Pfk36gq1ueqZW0RujKg6Z8E4cnGYV/k/jieWQy/SYLC1zSONxcFhDviZ1bjy5j+
FmKgp0oXsyz0Yy5OKG29KXX0r4yvQQGaWCaP3RlnFtFL6H8uqONorWb9ClZtnWUZ
OQ+jE4BePJCCG3CEWzS/6mMmUSelqssaAn1AvUcrRdbhU6izr55xdc2cXbVWh2L9
AwnaiUsYlE6GcWuq48CmXqdbqQdLgAv7f3YB6X37PTVBOsZ4ueFO1W/LtoyY2mci
W0uFV+bYGYoS7stxAyPlZODDeiwNaxz0818jxFwEaS5u4bs8wExDuYUCjPeYng9y
Wg2jGakGMXsiI1tOUPP095cgw7AFwHUkQSA/lCl8W/ewVlb6pzQaTEV63U9+H2KO
9Z+20AXMvWJIYrY61BH+hkrkSm2rJMjExEH/V7Q0tsSfqbCYEpl2paYxCtCn2z+5
wubJaP/wVyY8LRi+/x/q+ay85ytoCVnwAGVRehnumF9XDRRkVsRHiRWr+1JgJ8rx
IZhIZbp3+1xfZnFXW4OqWRGfFhzrnXCRc/NVmrf+8B/XBXF7ViMPoUYYF96P6Nuo
kyoVdvFjMyDCoAUhfjzldB3eteV8iANYvr4UEYE7AFWoIv1fsoIhWhU/P0bLsHQi
rLj2PeDAnmuk/l43Ks7PBdscjXyoijM909E3HYW4z9Y4jPU/Pigq++9z7DIKntiY
G5DdSCEyhe2IhVyMNJL3tMCiqmJNUIaFYxwuv/AEELS5YQO0QHyulcGYQx4wK6TP
wHBHCUhIxd5wHxcOihzmbQQsu5F7h2ImwK52GSvppWZP3Hk+1XWaW6i4Tv3OQ4FJ
khpTSkQ9pIMZqVzEQoZfB6BSRHNppFXk6V3i0zuQCBUlBIIQvKnow0WWI0AvVH0C
lFdelTQeqA5hAfKo4pdQr84vBiLYcUgLwRqKvDIZq4XbC1Ki6XO/kDsN60P2/wDj
0FVW5w3qK98BG8HhST9HYvdot2u6NDY0ZWGU8Gbf8JITyJ17IK1WY4sa/85M5RY6
LiXZFgKQr/cQsMDr6iadekY6E711yNGwiXY0DVb5+ACfLx6qjuXHcPrgOLEXmvMn
YhaNEZAw4MerZSKZEQwj/S4KK6Snv3SlHCMNFvCqdzhqWq+dIJBgSp8LLgH7SHXt
d0+t6NaJ0J9Vz31m86Q9i+Ii7d1v09L5Idb8kVG9zM1UDrOhSokqAnHBFKdgMEBY
zixIS3kCYsWOqvHPCI1wahoY8XwUHXxzsPccZjLf429WLWMAU12itz8ZrmqV0faR
vlkciSSfc6WtV5kOhe6n02WMPsqhy1yzpN7952TAx/nmDhzbKSJ0Wd3pHZm08gKe
pzmSHJB19oOfD2J1bXH3334wRa/ez5/srKiXR1vAjnBVXKNbVVYw7+4b2yIEtvAf
XS3jRMGmdNKj0US47ErqHTGciwOK4FwlhJ7TMK+Xy77RSTAGc0u9ZDRMkEhhW1sY
gwTzoooEu0xiPEjaqgQOxhoMahSenZT1c7zznUq9d8ocqzSlmqnPQ3kpWV02FdtJ
6jfPk84c/Z5h6L2FsTX5/+Pgj2it7OuVuykno8uwzlnEk0EYSdDnpnBzeouRW2Cs
WJ58iPMKjba/L7SCY0vHzO2Bgk1ojdq8BgNg5xagjfhIy/Z3gw+cHJZQOJr8vTWs
lkexZQHN4bB46qaFsMw1g25LtUiTvWMJ5MsL6FExoOWtAIPK7G4JtutM5YDNYSeM
mhKqZRNfQFOt74yCCFDyHj2WHFiD4HVk8YIYbSxoKGW07fL7uMXcsOKbc+2e/P8X
R0s6YV19ZuN+6vjsB+UpNUOP3LkYG74LcC7p0LDb7ZyqDFfJZ489OOoqWltFW/Qq
9LgdaWecbm+ZkZwv6vjasi0OSqYVU2ShGuEsdQJoIWIG/2RUHObwWe8Lu0uIwzqt
wyosWc59gbsh91wrqmQoWVT/XJIRGUmis+xnhXUuah/kmZUChc/2HG0Tpf1lhqlS
KGt/xAJMv4lnZaS/sYBy+Os8s12F0qrT74uPZrJtJS4XGqm11PoYKhPnRJB8sApC
LzaJDcpDk5qPYIFWbux4cm06H/J04iiwM0BCywsDK6MLhTYsVXXM5iqFjAw3GEmn
EaxaIw+vWawQWOEbhcDC7eqsbn/IRIGeMKOdxPCEEvTOPs/Mtsw+JDx6oX52k2Z1
yQc4yi+Qnd89qPTLfuOQLTC0qOb2qUARH9osTaJTTtpw58UVnl26mFOdiRUEYec5
flfqmPGVjMw5BX3J1yCxnIBdMntnEf79XMb5U/TFBMapCPB9zeXfh1EaHwmuhFPk
/uGkbXSCdo/KO8tuxuMGFaT5/pH+dY69M4jh1eAuwAkdwfoNUFRaefMwL2zDLhfi
cpXthFDtqD+1wx+3uK8kQv5mKnpiMR1Tnpf987AINvUh4nAyvTwe/x5PkGBs20p3
LWIbONOZcMo9cbYQ/ybl64eXBro+7U2iXj0YmPz3lNSH+WybPyMSyfNGV9CRVjR1
spvKDGFF1aw0HmkJ9u6WEa5abPhdNEy9Acu4Jnm9OxSoYe06KfwjtcP9nwnSwYMj
SsFaj1pCw48p8wdYN9JQ+sujaE7dI6/TvHF+ikDidAs+JXSRYFbYDAdx+wrkUzfQ
HpWXfyX8BfzyFMPYBkiY6tm54eAy2ZVEL0CYOD+V5LPIoWH6ssWvn3kVoE8OZZfY
MTU5xo3fDYmv1mzv32S0/Jfio0Sed6o1vKgft4qj0UTqdANOGZnCe86LuO1BML7D
zAADxqwizeyv6PMZMkafhReWAPBuCWjBpEDdxlEzO0+UKxmzwFgjHyUezpedgZSv
O0KXKg5B/fjil9kmFy9WsW+C6J4EmW7XsKCioBOxbEHf7GQVzKg8HlRlrSNIBAS0
8Xwjy18ZtQvU92FlPNtslIYfa4oJjRVuIlsGIG/FnUzAjrRZoit9OVyb0qJvIIYp
mt5demurJQfdFZScM1sgIWwjXzIjZFDsLUzqQkAl4n63MbV1pUKXA2Jh3DJPpZe/
Rhy0yh1gXPz+pCZtLQZt0cU6m+fu0830kbMOXcOFUKTnGuAH1hWAL72SuHlHSksS
830uT2TEI7afyGQSvlQqDpki/WA9WqgJNupWJ70YDROWaI8XxtVGYmNOWt9Pi3iJ
4cfXZPMQupPUabXxWfXfdhLDhXi2klfgDjEebSKE/Md/t96q5fLRLEmUC8SfaIrF
Y4VVF+TvVU8AAGp9aVuo4sksbFhnbnf5PKL1aolsj7s+iJPhvEnQRXvnilf/oI4+
2fjJlFtQBZ0uWDDR/tcvktGXOUZ87gWbfzigWdru7etjJlWToVbkvH2Tv4DD98OP
HROK98x78Y/kBVfnJWW017OulL81akbT8VjB15yutniOWfowLbPRZGQ3DuUGoS7/
6Qt8AMRrARPvqrEQV+buW+togVC0RxQhqRwDXLqK9T3oOQgSNFZM38puA5HBlkqU
RIlf9j9EFW0D/ij/cH/WeVknZx1lKQlnvOEXk+Y4cxtq8BaA//4p76b3oGRc+Su2
6BQ/vjCV8z0nWwQLD2tikxDMxPyHDDpG06owfAwFdjTLs2HQCMCL+hJSJYH5d6PM
DT8CmizDnpQtH0HHA/rBpMtAtRsqJCLon8+THOCEPW0BhVWbLsyuGI2ZUf+dViDn
HeYG/WInIPYPatd0jwy89RrwYXBe5Ujge3kJkg7x39iUAXWg9M/eXqKmjHKf6fS9
/NOgCVpBMVHxqt1vs6PTqOBZIbL9nmzgHxm8XcUyRLrRgOk1ErrBl9txdKv2ZxOD
Q0LBXWEfwEd82eTnOKO8oF93cXg9AbPVQe0s61FqdA2whOkiAaJ71ZCTKb4VoTU+
D6SXK1UFro7ajpXzb+V+i9FxeZNK3akKVnLz/OkkPh/3db3qrMj2zPQybuxe/5/4
1N8IH8KlxB7HDJY3m8e8kbq5uh7+csCg1CdWrDYu01ZDSxqvcgrP54F8nf+maNWu
k96LFXyVFIGEiBAo2pOZ3mOgnI28pUxPjwdjQvkmTCBjuJ7IvwOq+2M6qxUurLuC
YlBcebmj2SE574Awo/ml1TbbcBXvk28e/VHlSD/1I0zqQfHBR8y6eGsd+1PeR2Bo
xESFo5qBu6zigqrf/FrCRVragdWAiA3m/UohAZ+EueP5RNzCOhSfK/whIZKB+RVB
citIE4j+9xCN2lKFZqg9aeQ5kOMf5nS7pexaVXmixJ9O8QtCOEmGM+6tMfcNnggH
AGL4y7nfLaCDJtXrylRKWyZjlLPwAy7lpZo8w2IO6YRkXs/XV/t5N/5eGOamGmSl
7NBoildZE36Un+kmpMXc3yADGqOP8XcX1RMVAUvayfEvGwpexapiF6Llk+VBdi6m
ZxLi/FWI1FQ0Ebd1c35/OfZXsQjbvtZc8sn5PlwGfWCb27mpy95zUB5l/nyuC7u4
WyF5ty/38Q//d3vA52rCTJzArnT+eR7Ri2WL9HD5pNFdG1N7bDTbGJ25Ad32PnaD
4WLALrtM8C/5nNRbZ5JCAYIDLzCzT5/5E8GDAVVullDB0+T92F0mSSXBqUmHpmL7
e0Ba3bW8CKqaLqTuz92w4pTHjUhY5cyB9CZ96UDgXO/kBzvLSanSQIBaBGO/oU/+
WvhWs4N8NK1yf5FDAJYN5rb25/pX/ue08mkvoviZVxuFU99VYHXks944cGmP9R1H
Uu0cT49aNH4GjO+3oO6DUCGyLl8GdLzDvrW8pwJeNZSbTXgKaAVpctDh0x4p/zCD
figXKiiPomyEORfQ4wN4l5uBtA8t5jhqMHL+sCCXin2P3ke19z/qZnEzfCPE2fA3
HYE3Q/W8/jiCYv0S9QMhWBg7pVNK7nz/WBRuTp9Kqdvcc5iTG9MyVhAo/wCn0y13
9flxOVt+GjzKSEaczwaKjOYTucjzuQuLAKF57KzUhkF8xcnwPL1lXBPg/ozAjxDN
rpD5Wnn2ckjwgW5qJgpAYPV3zqfJ8hEruelZFXPsoI9TTFhT7gsD3lAqVKS/q5Qs
0lLHIOMu8dLcwgwbpfzcIO0N3d3oyWVCYYROU1PMSiRZ3AxXFw9muUyHnOIwAoB8
JxKEi6I0+Rbnfax5yzGo6kEcov0nSuXLfh1V/LEF0ZgxLeoMVGVMG+U6HRj/AdAv
lvOs4+5RkePy+pUYQKhKCre2XvZ0YDIJgdqAp+sS2nqxwfBda2X8HcSGxh3TSgxs
DL1wjSL1qNrgHvhiInswFyjpozGbn39Mq8oOpdOgvPwv5t7iBkgCVa6IMUwtQbBp
xYvmyIZLMHcD5ZRLLx5lhS2tGpGspewQiNfTBLIi3P5uEOnRi3LZUOZWO1a52PXH
+3IvLGRVCKMdrpsBfJRt0zOOOYHetax7oN8EWaHwSYINbgH0t/JLebUpQTkDPzZK
yTrgn/yIDwSljgZeSU6+oa7LdfK7u3LhUBizby3Gh1aABNvgrr44aTZocHD4n80l
0Hsah9lTZAyVZIyGtZR1z4s1DGIr3RBb27w6mjWUYZxqiTfko3YWhy9/cuCUjoBH
KOwS40Gl+5kPqvqaGtuks/JtYmcyyGMBd2lxNcnCy7hud/fzK0L7wxsDChWfboSN
0225HFJ3uViWZQkzJENMP+NbNZTd99DVA3B0Oh07cXhiJzteQ5mATZxNrR4P/dR1
JU2npgUhsBoTDkgJPx+MvtG53+pyn2TkKNGHXYPWd8jxbrN5TimHzvjmi7EZZ3BX
fLxEyvSzDypNsuE0ExpT0zad0Yc2lhEWd6FOoV6FKzrxQLLD2f7kxQ2ffLpRMl4l
A9y2qXnNFv1pjTd8K725ve/yOyOx73ouWt+cLMT4qhaDGtjnry0C+wOQQjGwaCqV
kuqgs3vzyMK01Su9loYTIX+AxZ096vdPls+8a5gs8qG23EdnbRaEyjiIw8kcKQe6
w9NPEuWAfP+Zu17Yb17Ok6U3ZjPZhdx3Hde1R+Sm6cY5qceepYmh5cDymkl+5YdW
ECvfnw3SanRPLW+5IPrmoyUFEAk9I1yBGgbUs5XN8IbOSrh2bFgAutDgGET/DafH
QZpSqyBWMks30W6UKzYjGZuXkVEs3bCAPdoOiGmbHF8nDr+cOeh0Q9AXSV4YNmK0
+ZgGEGNTS6AeQc1HaamhKujwwRXo5FLx6aTUfcNhHZ4kHI8bo4VGJt6uHn6mcfpe
teg3oKWlBgKCwVTa2lCUmpDAXwYXDLVPC0wh3YRxOvL/O17LNel9Zw14+EOrjzos
cPl9l7grVfTxyboHJU/ydeILU70Ziawk2tnot+H0KZOTpC63Y+4G/OadBfR0s2kH
/0TbF4pLHM9v1O29T4eccsNXEf07cAXXT0abh8SuTasZ2jRVKvTkrQEogYFp0ig3
gsg/P6mY9Gbw2Mdhtm+PkHL7RbtLhRCl3cI6vnqKgGdymcOtzxGvTtMhI/74c4Z9
mJTv7TjMnvndCm6kvgMEOwWQU8uUy2NYtPxypCOZd3SmJLIj1kF0UaQxknxEL9Ul
RXa7yk5BdxNcIO5awNn9K5zcMk8Of0NIs3tw+xSrBupdbs0AMN522oAkKgeFP0qT
5hxKDk5SJG6t45jkjCBborvKOSCpMXxLu1sbYQRvwJbTiToP/EG1onMlKhsHeIDO
ijMMjd1Gs7DVhczOliNrN6FCr6VoVISQMDIbkPutzSOE6eaB44sYVWaSfFbGA7Rn
J+bcKms4azMeEAeYbVGYrxheoED2GDWE4Sf0y4kd5U9map3sQMxqmEf/onEpMNvI
HvKQmEGHtdoXntPFxZCwB+ZEBxrNa7Y8jSW2WFiyOe2DuD463FFbJodFpku/Hw3S
DEvh0NKc8aZkgyvwcOXZlBzxtBaFCTg4dSowx8azMlnnEK8uaSP0xs/gFPgZbJIE
g4pLZv2D6iyhkVOGfQ31VGmL5C6ZqKeXF/DXx8m0ZrFUAFFa/7b9boXVHsaQwCW4
8SuxjU0yaggkWuO3RCGP8pgu3qCHAhVpKx6kQceLurvwWd+U9bTzvkaoydR3BgS0
qMRzoINTUtgRiftnvH5caAxJgkFEAXfdHSeoAltIUTDsJNbWSVVVyCpYMSn9phY7
BJflUtloRbXlGimLZUvqSIclF1HqqcxV/oQ0wKuMJ1tZHaCdX1nWeIdqpqEJ1cuR
npYDqsGuTgZkkZab/8rKrH3xIchiWZBAOBkfbHdPDFlF27x6OPqi1rntZqIhNj3n
an6821cyCMIB4GuZIYcto9AQFd7tT/B6NGOHsXzoaGnLp9qeShjnblNZ2mFtK1yM
L/XShAMmvDrTkY5gOLX0cIbCDjNgdpCll5NWin7D2G5wyU8ZQI+qyl352r16zZwW
LQ6tILAP9AagN81d5hqzPybwEe/F2jcOKhW8TzsQRFUzWLOTcLJUJucFGoMLYnd2
o5rXv7FeGUYzI8rtiYCNB0G34GlLp9nFHdJW3J1PwoGWinB8hqYpVGCFVVl96LP+
CFSYxz9SeoMJQXTkaDRMz0LiJOXoEAxCIOihtZxgHR4ZqNSgPwlyVDd3VaiC5RDj
8Zhyj5aNk3b2QS/krfhgyizbQTKQYgr+H+fWiJHlSYWeUPlzj/DhHQM3QajrBe1g
4TJhlO8E6rG29Lu8gEOz5nRqCxuOcaYmhzL3Jx87f2CMsMacnTIeITL8YfEpLMQl
zmMwep9fwYJs0lkDwqybgbhFoj8Dx/UpO+OzUkq6kO2LNcjlzk/smTM264p5/MDK
MZ4evnI572yfK/0SNlbjJ4wA6sLI+9xuqVAcysK6wSDGbPnKRE19p+BHU+feRSvM
vKRUABKO4/ZLX5R0KPMSSHjUUZjwpNgrPm2Dd+FdrwG6/wXLbTrNBqm4kW7IhgZm
NOrIRBUJvx1VJpQR/dFxV0FrkxQ9UpF/vtRZqFZlEmRX6Zs1RYWUxiPRIaap5ud+
2FI5yzRyjgg/ocdot+VvwjuYXsOYPo3Q1yHECIhOWMiLmRE/P7B4xPDvYoOYNJld
wCcU//rLxrEY/nLo/s+MOjA/E0jc/GbgOaZxR8SS/Aun0t70D9qsXjB+T2+BJ3ZG
z+86sOQNyNL09XHrVkRkbc/DFFWzkSk3rCOg8aLAO6eW3qNepk2a40BaWbxRhtxe
Ycb6AFe4LYeo+oFYhq+bQbs9lOvlRfny9GBft3laGsssgsCgN46z95XTeK8zFD7s
4LYnGgqGf63vV2G6zWZu/2iLYxWnKh5X/H50GqSRY2ZFIH+TgvFV18ppMMw53NlW
+/atcc4YllWvGjnHBsHrq11D9o7aeSRHiPOSP2kiskbgrJg34cC6x0+EonYf9u4P
jMr0R9MiNhSRV7Q8blKbUsJeXOzAmR3lxctLqG/wwm/nkuxjX5Um4ul5CFKu51oU
054ZllCNbF7fnmC549l0iMdJCzBLoyPe/P309Kee0C0V2+i65CaxQ3tzeKppP6sc
jdrKg3lt69NKUPKDjdoy5QghpUk4I6U0LV5Qy7PW9QsUqwBWe70rPXaczk7kMrvO
CZL8u81/qkPKWN6N/EHUW34YdiT7cHnKpQsFdpEi1rxqQc3IqQHvnCZ7aaBWrs+j
vjsI9MaoecoD85l1RF5hVUfLU5ejgQcOPyaEILgW1yCeC2rqzvq5R7bfxrbwGPPJ
bCL9pf3VymBg95oHMpVBM9ibscSAjOL+EPXeoJDZdXypLRRmbEIOanNd/cH/nLS8
EalWTqt+djZydyvYDBuj4GIMFuF/KyIT0/VbovAeGxZ+GxO4fVb9rAyiJKfNrf1j
7QATFouRe15Z7plCwtBnlHMwgi8JoGrEXmfwB7AMJd50IPrPChL/wqNgOYIQ888P
ajfa8IMK1jbdycqja16Rb+E+iA90KYnAJhJ/Bu4HVIUbccQk7sw2uB8UuN2P0g0j
IR5kFkwF8dVRnaVSfrc5122vtHRplhnwJSZSbKpVb4tIKZXKb2dgZ1CZXgehUZMO
i93FqpxlEoZ+RfrvR83LGLVoLW3RUCKDbVZ9u7eTv1PP28uC++3B37VuitOYiIVS
aZjlmeJpx4HRMMPZfptE8xY1Ga2jiqIXBqiUAxGqZhqMHu3Es2gA6QbaqD8sGFAN
MXWo9yZh91C564bhFMEa3/5wZVwwElECm523HL2rVNPgcWj02Msi85lHUY8lTlFK
OVHZnyItchXpM0wkWC/9r6jpL4dDVnToSYwEizTczWZs+UwmEkSOV5prnCQX+DAI
KKEpHQtOLtpp1WjEZoCN8fAdhYLRjGPW4sFM7ELeEniz5AyF7YCGHsOv1og5BvGe
VUnpll307P9WGnIbLpinPrDD9zl3darbkL/JQ2AsbjSAH/QPzhHQEUX66LZb9N5Y
Kt0YpkkxVPCcHqbVROI03lWbZlMAU1DvZTT9GDS32z/lpz1dIRUiUD0WshYtmo1E
nhG5j9xqN6INPFsTtKc7CmCqT+uIV3Wgs7gJaiA2J+uzLvDHxD+QsCVfVWNcqAK+
o4aqkmLZq898cHKipUO4/xyhcEjXAvgNks8p80CgOnjdajmre6HWzslXcC3Q0QMK
Q2lXyRC1osNwK+C42RPIb18QAf+GnQwr+K736L3lEqcS1Ez5pjAbEZUjlYdt4Xq/
fEKzu4lCr38BG8fhIj7mdx/AWbzod51wHTPab2/UB689xxz+8qrEry69OL9Kw+kD
Sdr4s+v5dHq6ExsSyiyr5yUstBjMM1M706OXTgTAxqkzUtIbh3Z8k7fevZXWOz9X
WdFpMd4DIPz2lea76KSiJEzL2frI+UWw++GRb50RLO3i7OOLfgZihgP4DYYxpN1t
jALfil2DLIHDWk5i2aOgJe/956/LZrkIFLypG4kkBqPwrXmrRhuX9ENbRs5FG/M5
6Yaq5XvL5eFu39I+u3TMjnldYMkHquMgJqgnNHVvPIBBH+dsKklQ+Zf9kqIgT0uK
rVVyUgNejPKGmIIkSu950gke8kTT1RuZPxiEjiaFgOFWOYDPfvN3WcCfssLKZ9xC
jH1+nR5NvdyBJ2jMc9nI2T4kwCSOkBhrB8n1AyHGNaeDUtcyXNM/A4af3K3m031K
Q6kfmkcjXiE0+PDnCMA1iTgHWzPyjMWBaIIpG5o3m4y+ctor61ZcoOMutklTj9yd
r531fopdtAyOWNhVwoIu1ucd+itfAEhvafA1KOJ8qS9E5tRYKDQv7O7IMadrgoKj
PwgtVH9rxe6CQBKR1HuVMPrWUOd8uTJhhmH8a4tBcz87Niru3XSVoDSNqPE4o9b8
E75S8jCZF3fNuPIMWoCarh1xg/Ce2A2K3NIDn3+RRHi8mUgWayjokx3fkS5rqOVA
NGgIj3X7sbDG87WYFhb/Eg6c/Ra80zzj/uiCr+4z7VUr33DqQNAMZ0naVZmoGYTB
QXPGMufZSJA/ZWjx8o9RmjDem+LkzPaEP662+jCPZdon1hJlsL5C9juHA/PTiW6V
favK0rusVjj9iSWmKtztLTBGnf/8PPpRJXKbSGB8gquSCQ0xFK9Avcl8uU3lUyjf
SaEHgPdI82N5qUvRqJnONwPtAVWgvehnnO3Ez/ld2mYs9GulY3pEc4r/eimCznRM
Pq4k/dOYu48vaR3EkbGT/FXo7lI+mF7WLxxI+nWK3SPYsJ02PQAG67glYTgVwrIz
FE4n4I70ob9I+GBrP2rzaLvdsB2OU9u7/8A/dIqRnGvOEzboK8GWnV0WlS2bIiX2
sYhbFrI5Lz3oqei0ytciuHiVUqK1s320e1R2P3Y+Wsm4gy0hodO2yhYv3JCNa1fJ
TEt+9cg6eQ1SE0OwdDvTLZKra7t69czf01SYKrCGM1kvvii9q0nSJmgi0uwM1n+S
f3h7e2A1gff7TTz3mjuXC/mbSMdHBo6n/UzakwfFpZlb9fJTOyZQ8CJaGNKyDlE3
8gVURxgx7Gq8wSrKxiws3nvz0/BL+KsKazMxulG2qX6hWJLbbGr4SrTJooA2DXLj
Rm/zLbP+5pFjh4ZCGdup0jepLKE0oFXdbfVz9W3ciS0tUYIjrZXiHTjBFDFILLwn
OEuxryz72QAUfDrgZBpgvpFnurcWef8d505fJtdxv3hO25C1KYtD/HsmFm/O4Nz3
KE1LVHn10q5cIKj2q6uGd87MunvGDwilqGh1CIPOTzrvoxavRSjZbkzM8I/VE+KZ
dwGKpvDsrEAPvK7KzFOupGdUCc95UUQ1njjO4D15tmwnEuZItYe4SsfzKCY0UGXS
UIp4lqrjo8BVU+zWc0yFwbutnTSCIdn7Bl66F8YyL7w2UmDjP64aCekl6eiGSn2i
vLOu6/iMmddz06NCUAzD4MMKvXN9liDxq8w3n2xI3avJcECQivvfQjAkpeMcDPEr
A7TTzTPzo09bFfRQFsCJZ5v683l7L0sGLsAD4reRXCRMdVZDmWhDs7gGiztMCQIb
JZrEuB3CzS58G7syE5x7PTFM3dl6gNgrpuWQcFzMPcFAvlLW6gFeGYnLbFHtjx2s
hrCv0N5CFt3B5Hbu10qNlWteWCp1f6jro94ZuqAd+VqLaZ9M7bHfsS8L/OrtBRZg
JHRBau19izLqsBhff39nGwFC/yJKro2HgyLHA3JMaQNnSuQswZBAsytjuILhKA28
LR56Ts+7tU3ky78F2fFrvFZUeTh/aWQiWZ4H35Hv1pncuSDwTqVe7pC/kBbUsR9L
fe8ZCcxyi+ZO8Myky7BUWwV/kt0BHeHT3nJiaMWgoEj58OBTt272dU1eAajj5U4R
+G4YA9oDkAUUBBO4l9NA2W+2ZoZGsGvncBYsLYiCwGT3W2pMfk70RNw69q1S5IHT
TvMONMXfbskfXMhf8CPZ398Z+oKwiq147uExygmJAXv7yfphc6XVUIAVC7kbj0xD
LT5as/h9/cosdJU1BDAL4M1LJl/pHsUNosFLaNsMqn9PVXEkF+Pnha9YxBhtctPp
kxjWn6DQpE30CwLuuEv2Pu4VxMjjM5GUAynFSCe8x45BACNthkvB3R4nFb0ryOkv
E7ZXYdp55GqMxVVV2yaWav0gPFKMimyc6aowRNqFpsD1CrkB9OY0mEh5wCYgZMKy
k4ItbzOsDhIABKS1O6ag9PQfnfdj/U9kpVaJ4AkqaPIjyvCQaDh1ilmcs5UQH8Qc
jHgm9eGafuEqrfsuN4YZSsa7CEo5Q67C2Fd6/TYEMBZJ2cC+kVwvQw2fATdCdu/H
7GYxG+QMy6UqLngqZVenj8sy+WIGD7N1ryzIbU+WVnW/LnQ4Zx+pZ3og2EA9fPDn
TVc8MT8YdJj3CHHUlhhUksWSsPytsKFMgBsnyhGPhKxbV5CIrstTsgzHvrexjZPB
Pzg9Cn1LwZit8b1dy7Vv2VpmZfprxdQcghFrleQTh+ZU6PRpYBMoAEBz+kOaadlX
oba5J53bp7waGC5C/XtnF+qOVVvpefRhVUIbzaypUd71G+QIVrfzFysbJwCgEmlW
mpoo0XBqXsbTPH1GSe3Sv+XeQdBXgRqkWCsVC2WQVRvoeNZuDtL22dirrAslv/HJ
eRYvqHE3WH+SCmB6ciRJbcEwt3eAH1CZJ9Mc0ziTnaDtqBnCum6oA9PBn6SGTLH9
3eDilkm/4BI5w5IchXp53ELb+oMk0ChbkPP2HOPeOxKCJsYaKORqYcTDDe+pUBXz
5CmcasVYZ0eABo5q8CPxlOHLzcZuIKZQ5W7qOQjpl1Y9qQsHHXUx+YhnQVTlVzta
G/4lBdVmHqqM3SBgzdw1dckrMbpTFP3aSkuCTbD5stw7EeLHf0cRQWM1q2Z0b8i6
h0OqFKMyp2lIeRavouA2ZlxKQPiXCtw+pID9I7XBRtYBqbPDauefWvdjwxz6WtVO
VKZT03k9WUbOXf4AGbaGV36TrH8rzZRx+H135EYwKseuOdj7vH47NgsTbWHCo9HZ
RcLJ3aZlzkMOdyUb6lUP8nrYQ32JFgPnttSw5frklmQwLImQ5VuY0yAiWCC6u7L3
L6vJVTzJq/+lIqo2SoWTh7Oa07RKaeL1mypJvDVJmt3opXQ+yjSmDmOiqlVy+2On
olK2YOCUsC7MhvYNX78S0C6xesLHaFGFjhWWi4rslYx1PyrWK6036eukLb1eNcTc
mwG8RmJWkIWULQgER9/l5UmAnsZPRIQ2Q5tqaWVe9E1BtVOUhMEZJ6LFqLAPGPcm
NUmixSqKwevvw/qW5atObIam8v4OdgNXdYNb8fK51u5XY8NsxsOivsLaZVe8xy+S
pRDgNoPpgHjleXzoR8KSlkVVlqXVWcO1cznAy4j7lnIDs0tiW2af9eAP/CttvesS
YjXlKshbLzsYfiqp6J7lNSe2XpgVNmWhY00DsXJQPiH6t2MPi/UZjgm7fpr3Bxav
5Ww0dQert8Sz1IU1as/nIuM37aVWvXnXJ4rZf5VZ/R9DLoJe+wplBt1UTIW9J9UF
LQU6t2NBmDixBKMeWCazqq/U0D7HT23Y+dtLCL2Z8E69r6ZvhVf1qNBQREWELBEj
g5M6pk/f+nXNYhX8Pt68w+HkzH9dC/CCPmzBWONAKWC/s0+b96DpJGIMa/LOO82j
zGCBQEmg8jPDAaWE0JLi4fUfA0qMVuJINY8fSlzxAUpF8GeoMe3/IFEmL01FKu6/
fIAf2AYX1gEtNSVWdekMFSGLM8QvSK4NAuTyufzlmjniZZU5Weh5cbHSeHEpOGp7
CnkRG8G0axb14Ec/QAi20YXLCkTk2l6iRJYY3R6ggQ/R7zFFPXv9YZ/K1em8z9d4
PYNZRkqdvWHKLdAaqc2ULWUyna/qzGCIFMufRnE5TfmE8kWavxS+lHHA2aWIBE9+
y/6QCifLs7m7SwtiqBs5dnRoRwDi/MKZPg9VLfTH9lMEltFWE6mVJo7OyNY+Sb6n
GVQdsvzUQt4bzYvV3HJGMQjMi774TKwkx8QZIcsGpH2humJ/cXslqawMLPar4+QY
471BzKdAo7zk/wtTs6gJLSllEPWCt4nbmfebKqtjoW2twJdu0+rDxU6rQLfhOQ25
N59appLh3hBiJqIudLZmTbYLfk7axRHT++2phpe9Z81WgwUJy+M+Rp44pizWoUg/
KIyA84Zd1PId5vLDMAmna1wAt2qtqPxfIClUTKT0lVju1oUV/wIj9kdwcpu4WKzX
fFke2ZC+EsHqrTKXYHWEss+onp9iGBkHvC2RbFWqFO1Sbj0XedcfRxMKyqWe+LkC
us8BRRUWhmyYYov4Uu72b3Ke/iBwRTIbzpJSwwEApO8yQOgOAGsdb5u0MDeoOwO4
1BDD0JcudVJcUTzpQsPMgIbfBMGQmUNGePO0urDVpDcLQtY4rErHbtYeQG3sJwLO
s1GR4cKfNg7TYFuG4fjToMJ4/71E3Zo5UUiq/UMA5iVOuIoNTm8XyTKMOqv4rypa
cYKTvPX80XIoB8Jk8WDP2kRujZ3SFY5fLcJY8LZghpc6L3LUz/6udUHVmdU3yzd9
TEWkaNBcqMSBPQQdUI5bC1XU5BYyesdUQO/HqOhE0zQcuBv2Vo6Id9c1yuQHGFVG
+IcInUOpALmqkKfQFIOc4v5QE4ZQnBMXiPfT/wdhB7XLcz09jteIyGa0FSjBIBL8
3jRXU5y1PvtGdIgiQ0oI+O9LfA7u2o6D0bH8W1cDZGfCAfyvP92lmNzpo7VSuyk7
18uAFjigMgO64TGEidyctMW1lxXl+OoDHIga6icS67wAqMZfoKNMoVMMOsLyYe9N
pRQ0YI6tBxh9fTjjfMHXmvtoAQkYA4w9W8uQ+BGjLBtBmRx/BpaeK2kww0EcoXpk
zpNFHKV7JOOJnbQJdJn56VFsEEVTE8bk4vSbuRtFUqnG3Ym4QnoWK8+1qubNZsQV
bP/CsguLXZJWuXTZqWtNpPppv+BsdA/hLwgr4HcG+EKu/RqNDCVd7kvyvoWS8Ysl
RcQzjRI37iudDNW+vHvuhmR5kyPodxwOvoYv+z6hXQ//fR6LQMTskoJULKjFRORD
hmhKGD/LM5UyjvGb59KSrCAhibx67j3sgwWtTfqbD2IFBUyWpCGrClmeUh20X2ko
E/GQOaYvp+uELpTCw+JcbWLo01ggzscnilQ0mCXTGsqwFcs/mBKw+Ls+2CYBNkui
RLcbKGQHA4KtLcrQDiw9gxJ50JKddRv5dgzLvwgglzY2tmgG8rEhvOMuO+EqJvm6
MTBHEYo6DUDCJJkwxEBcHdD3SFIBp6yatFdGF2LzikXw1wx56pijkQSEmxOdqdKY
XSah/StN2OnNSibtNhhlu/v0YBiOW43pQuiIbgINyTY4StHS54HCWaF9bvX3Sr/D
KHP6p+mvVgUxgB7fOWHXVmUVL6g4z4cWSLUDanwhD4n8sBpXl3XclH1N5G6x+pEC
Lu6gQ/l6DYFd3MvUCTFtMHeYkJgqhvupP67jasCAXkFz3YjUnryZnkCgoY/ffnfK
e383fl0mYI3rP6/N0+N3HQYyLPsvBXnG8ZTy8Pndl2+G8yrnyozJ9o8aN6ahBaGC
dN59jC5el7oL67SCVAPVcWZ+N9PsTyGNzGEul226ZaOTIWescXCKA02ft2PvQpT0
pF2AGTDjFLTaOM2dS9hMJcF5QeRYXzNfeWzb+7muKCdo5DpMAAMs+IxrXHwNPodd
J/2olNIj/L61KvSUD3sYZkikgboTwbL7Ne5MU7RvjhPOIDmHx+756oj2X7FeLd0D
acddxf9Y77Q52hxDIKe8ZkS9tkzfqYK+zfgtj0su5w8lmb9HaBfJa7sJk1Q0fmA+
8RUCS0JU8sO0c3Yxd04tBJ7yHDgGTY+YfLnl2MT5ALOX+rDp5XLocKlvKDvD9Unh
LipCHzEjz6QTmIUJvjguUy2fotNuxP8cdD2L1SLutsFE11Pl3suZYz779MDj39u+
4MyYQxr3nXW0ZPOsyfHFdl8ZYfEX/ybjl3WUv+gVN32wQ9MrrwnPmPlCIf2uQbxK
B3IVcrhNA0Nt1T3a+amWM+YIj4kOiZmoMewN2DHBXP36FNpZQTiVfunRt1fh6pVs
Z54A1sx4Tp9sWS0k5wOY5xQylYvcgu1MI07AYLseFSVjYUuAogWOtx3MgeuNKXBZ
fBw97Hu3tQJcZCnnOpN0jTsYI336B565zcFRkmdbd2mYoQml7eyJJjahBkbIBTPw
fO+7o9FEGVkSJTf8n66cwSH2A+hyewkHiPHHDMDp5pKnt11+hD1NZHL0GqlG7Hdh
KX9UBmjE5bJ9R+SB5WnZZMZCj04kZCi0xmU+zNlf14zBZyp0BTf2rMOadOqxctgj
2sf70sHo/kcY4JbLhDPTPWT6XIxrdFTendM6iiJjvE0ndVoLdr8h0kYhiVt4CNqR
guPhxJr1uG0I2rO20FcRUDuTPPaGeheFFxDUnEYE1juuXTpTPk4gYh/ngF5Knjtf
P5K4WELxa313LKheSUWN83Bn5PTHrK6Jr7kMWYssKUE+0m5FCaHHbYx1Wg47LiXE
2xXtwCIDp1hohC8Ak5EtO5EJQLCZyUVBuZuFkTgDU7Dz5Tl+ilnE0c+9Hlyuzzmd
VpzLrW0lencvvZYHqpvvzMgplhelCQpdsamdr1xY6T13yhZ9SrKaGYSGuAfNRQU2
QYNo10knPEFW3WCud8qaEDxLqAFIAuxrShr7A+bmRXV2sie56DB8li9OHVqhXS/i
FCi/s0dAzyPNjAx3oFy7Cww2WYL1Cg1jQ/8PoTgG60rodUumsdVEw6QCpJsLRhiu
4dC0KQ+ZO9zFmqlDH5KxPr+RAYBvrQcxlQH+16Qh3qbEiKg5bkno9UFXk3tdltwH
kJr1j5XPrXJ3uwCiO0KDwgQJCf1yFzmmLDzb+60q+5A1rc/ryOE8URqdVg/UV/V4
y7fz9tdWhg7D1Pt8/ROk1dCqZRYQSUMgtSNQibwp/Fw1RLqkm1eioz2hNoFIkk9f
sJljOyPqxfH0x1LCo2TAhKgBmDRb6vKjVj4k5LQG39t7DQl3uocQeR6sSvEhhRH5
RysfGZdLJyE2rsA5rmnDngw+um8CumYpcUuEwnFKYnQv0YAHZjJdBi2lOnMQFR5+
GSQTokDmiOwri98AaDFuH2DfcdzEiTQXdAUdDsLNEebIRqvsEn/s0bAgxSTYYwf3
PdtqPZDFK/NhOKAgEtt3cTNmws7J937DLRlX1KYDABeBs9w4x8TfDCToUItDmuYv
lPkYZVmDoX5SE4gfoUdEbDrFDMd+QJLbachnYINeErTTwYvwfWuuL3t2HastpsIU
oaTV4jHsOftmUY8pB6glzNl9VRSZeX0o4f482SEPC/E2E0A8fd6hY4h6RIMqWyP1
Dwe1vkdn3RApL/HhFzBXj1DGb1omWh5Vml9McN4dKzfsK7AGr97jJ1zxQAkyZjyp
EHd8cVmB+Wc3XkxQjPn6Aj/p4Is4DiBE/zHrMdKbNXOOCblaFrSzuo3YtIiyW9V2
qdFRtsqntW/1jhpdR3XLBfK4CNAfdh0oVXL3qhWduJqztGDnRNqAEctCtdz6YjUm
Cj++l6WUNgvIxup8xQupufO924xzAIAgMBUG/oLVIDDNdq/hDYXNwt6ZYKZfuQfd
VjOkMK0XYjdkLaSAJzAn0hZyZmvLuQN0S8Hwbis9A2ZJTAdHpXgYrlJKQqoOMqIN
k+34FLtTH9dwyhdu2+a++Rgr4p14jFKrApDuHtjOTQ/xl/D/iCzYJaJ4W46xV5g1
cSyE4PJnbBHo6z9VvGRBGuTnLmL2DyAdLBS5qssNNO1qBdvxYCZfH56lruATYHLR
QE49RYfgvBuITGBpniW1/T0w4TOLR4TCUpCRd3saU7OVECUi9OJkJQWgPuNi4NaX
UiwbTMAEhTqZyMd9XG8UgkR6AlvWkIO/JLUkpbfQefr4VHNBlkxDCx/riu5B3yfT
t1RK1P6M6Cvgvuo/qsVJ6w1i+HO/QEcuhSq3oVAPILKO1uPn79tYljje7Yr4Ef/x
IFzxejSNDrfBqqsdmWxPyTYfc7go9Ek1d+zpkwbjiq0PANw3YW+MCM87OZ25Yb+s
wlQRq3Rx9upseY3dhHpgl+V6/+NsJ036P3kUK0FrocWrb1R/eyYPMreM6+A50NyK
/hh0U4jqfC8jkD0dLF14NlEUD5wu5HeoDsIwyNowm3kJvp7DhL9ZLLCxnHPASkD7
Qvyb2b05z1JiPmDVTUA74+X4fE+oa2TG0wlu7w/ydQcbxTzZ88JxmajjMtU9P3LU
s7RSWLpssdULJ2HsgG8LFBQCwpUWy9xBOEce44jx810EQQHm8Gg/rltoOLnBbcQ5
7XuMuvTn6fd8PBAzoRZKu5/7iBFC8+oHaL1h33kY3B10CO6VtBU0IZXzYkS0Gp6Z
3R6JZ/vE65F337vb3kG+hdntugvTxOKdylVrrP+TZzeF53oH+KGdweJIa+nb2LAD
qDTF5jjghCglh2xC5LKtkn3mCT5sBI/gpfjnPFQctsq+Yo6ZB112Pa05w+UkePLi
/l6F9pE0nL6h0rLbyu82lDsPcrzb1U8HSaYK0rGchKmE94KVA5jtKPuHETXu/VN1
buSy0I6J+Cmbnuf1ej4Snuvk29NQNhKrprHnJXQUkHabMLdLw28ibQ+AH8ErLXeN
v6nh1Qxhml/ABOm8Bf7aQqRhQ2DSCb/oO2Q5oRKo0j1n3woY99b6CokJUc0t1BjZ
ruxKM1vYVqFmVOD8GfT+2Zvx+pmy9+7zWRDEsQ9WwmVbzQjSFQ4Xa8f0c7uBcbkq
TIROEb5FIKXU4KomgyhKRc9u5qHZh2lyimLX21zedsChqXLvN1D//Z3z2rlgndow
hqbaBSYMnQDkanFWv4XjXVbZPB9DzE+8DfpiKnTmFeSV7LpRkmHEglB/O3NXYNLq
JlK3td8AB2kZ0YSS9zmXYFQoZkt7zX2RMqKMeRErEiiOMGfSHLHqhuD2KTj0lqBs
KKxll6tyiaL+xGiLSw3yczF0o9HbaRyhVjp0ulwx6gYpayRLlJ3zKr1QVTzXg47e
AFaXfkVufuFZ+SRCL3gR2A/kkX8K9QQCK0Nu6+PkyMdntduPOOPW2j/Ifcw8FSEE
/AKapZKHsPuEyDHIaXFUZXPQxItOsXRyXuMdmZ+l3Sa/Zda4i57cumriIwfNDdy8
uIvBjL6JUo6VIArhKQHQ0ulN66MxTtxw1+EhFfOoAbuvG/O9k8LNgsDW6PjThkWH
B49fsO5aEr4533zg4S5hLvm8qEqwbUbdc9OqtRg5Sl3furJM8wg1h2YkH+lVP+Sp
U542FMamhphAQugHC56CwTNQkp5APydZjEOgV9afIV/NV+zDI8nU5yahY8frZyYn
pLKSgoxO1XIXvAqmpQUrxhbn4gRKDK4n03m7ltOgnoI3jzUhuLhCRG0zpfYdYICW
oTU5P5Z84w470bJT/xSHlxuS+xlyfyg/CjUqWBC+x1icmqJBEXuOGiyO4uNp3HAd
/rf4EAYweY6RXEcV0U/l5eKSTHHZRx+7tgVYguaY0clKPRplSm9AABO86nMI+2VF
Vh6L2eFJuhqf8YR59qOZaGOOKRrRAWxReoJdGNe7XCTdKUKWLcFNFGzYW0WaBFla
GXQpCDVCAVwp+VUWN8ZL8QpZOkCBLcVxugXjikWyS6e1f/7CB6FLR5WabMNnStJA
nGq+ZW+4zPvxSxMlUmfY1RoRwTHiUMB3KsQCd5Y0XU2k0+1ZDPldbJ0/eJ773xzt
HS+/aGn0AV0tiSZENFltVNpYiFruNI3fF1ZdVS2oysa6BOc75qd7KHhO8drOBAD9
EJm5r8AWo+DSEgP3c+SISXM3ClTDJjM9BVQ0oHHaqpdh1GhQTi464zEJfW8bOnG7
pzyCLsSdv5jR/OhODAZiviC2LIjJ5ANESLgDlJfyvFY7UkBi2A9DBljn0pdPoAPq
1+axMt2Lre28n2+GdABBhUwWBqgWc+6gNTaU5203dpFHkTPyOXOtw+rSnF0lt69U
x1YBwBDOUl99ANG1iMhPZtdXQrmpSXO64GYIv7gdPwFvkbHraEQbHBuSR5TJZKBw
cGM0E/nbil55giA5HefshfF445Pnd15vOnS4xqJcN1iGPqRjE/tgFEY3zYteQxfc
QVsDShvPrrzKrvnBpL1xP3mGxu+Vf1kaqJ2WEAaAyioTKLvBgfg9qn/h/j1b4k5w
bWlZb9f1ol9idPFnQLvcF3olsXhwcUlziDd26uRGxsH7f5gRA/+MDj2qm64ksRWt
AMnUutQtJtPNI8HZrFDzWfoVnclZnsltXVOifXZzt9YL0K2ZrrSv7skhtlfPsRr8
VmqlABwfv7EfNGFEKyhD5M6I0bnGZNUtj1xgsafF9f9iZm+ZG+NaZxGC6ZLCWwGm
+HSCm0p9npSiTrn3xpx5HBw/lI9CQiZOoUcpaOtnUoa+x1h6HQKImrTgz3b7JfYE
YYF2VmLvKa4z0Yrch9zt2I5m4dxPIH5C4smJeFMjpq+2D14Q/mjcWTiGthGXNEkt
bI+f1cn9AkyUb0rA+ErovsXvDvvVQh0gp6Ig8UMgZvDwOaz9nMh0vuHAxPFWiroa
AfseZ/WItgg9aOMcyLktbDvV13GYEQi31m7/20FdP5hSLdT7GqJ7s7QqA/yBoTET
jCv4WwvZ/OBJKgFSi7TrZSmKjJlQKtakYLrocPss2jNwB7sgd97R0HGaRuEfWg+e
NIJWPmsF2qyNx7/2eGoAXlEqPd3bNIDoNJmnEDO0zd/84Huq3O8+l+UH9YftkKBc
Q81cI9na6pjTNIRu2bkZctLIgupPOwbgA9k9HjMg74SONHGdJ1u998n/wla7qcQO
+tgMcRWCUwZBg7NeWgO9GKuwoSB7MAwOe/ZT0WHdOafM7aEEjb0j8PHGmGol7ei5
yeYdRCABGPrCJh1DRq4KqUHISvFGHeLKVXMEQdJGAmXYEV8IGV0+jHhMj5jk3Efl
AslIc+LZvXaCPXhejbXE/vnnQnU9/sWHPUvWV4dSehoX1tSbT68IsLTYYu/j0c5Z
QR69HGyRTj6E6QrS022/F6XKxshZ0A9V6MRWNXsNyGl/QsxSpd0hVSaKysnh9HJf
DrXWELOunlqMfkeF91o5YwM1bW7gXDrknrhEzxZEmk+TgV1AzgpPWrIGdspwwzTJ
CI6E9tVz7UtEPZb2aCExNHVwgXR5HXwnYj4ORqu/fodVKVjAsziSMe5sHft799O7
Qbt+wlzLHxrZUCbykcjSvXxun3JAE+4t72JfCJVqPHNLUCDlaNkp0h4bwdT+w79T
FqU6/BtIJOCd+ojDX5h7XKNpzEnvwr+hgFLBBF7yxC/6Mrs84BDggqKvSLfLZJZG
LKv7cPEukSA4uz5V4kcfCT9KD9jyZ/PeRYxAp6HaJcvXvIqjqXIhy84LMC5oZryI
LtAhlKgBqplVP+/9aCLH19HgiBxWPBVzKlH0VLDXcp1xcMLKDI3PEdIYuWNqzFJV
u2FV4LrNzABA/Og2spvZvVC7hmhZAGLFLMbkDhglAjdeR6WOlda9OJW2Dyh7vSZR
It7PGM/JlcSJs5ns0VW2vosCtoJ4dkYgJ/BeNFb7Inj4UqQ6Qws1a5rvrg6QLRV3
it+2vfaoMMD5519c8+r7inLpLJlyV0P3VWcX20Fx+cUkk4BZZLvM2J4ytKczFS9d
wyGuKuF3Jf5SyC/EUBFCfcEXcACMIBqNQaAupWwxueixeWjjJPjGzMrZcVmf/HL8
7OW3MCbUT7oWrBHmrjUCPHU40v8KLZwq9WvP2iAQbziz+5GoohFm95Q3j8FbWB6e
kDYRCz5HfBbtzxbD1OnyhPkRoYfSyMRWxzxW+pO3BXerzSKasXMPmKJ5L/2zrthZ
ErgpgXWulkJm6z1WBfuv02/NTlHJNvLwqOuHc0SETmrQ1rwJqCVmX2WL4RN+gz+l
3pCPXxFcYb76nCdX+KVevT3pRgtrem3MM+b3psjp1mVdcnO0Mw10DfhbRlLAglqo
vxHn4rKfoiAtUblZL6tlM8BQFPiXexqLp9cfkqaW5hdvGbgsz7XWwA3/w6a4cAFL
XQPmR+KywVUMf1qSpvp2b4/j8R8W35h0cJ7dns+bBdvYtol47tvuLyWq0AaTwX44
FO+GjB0gtyddcXgxj2UKjIKnPbqqmjOce38JLFrEbs+lC0UsYjL36hz6Yu5WYk0D
AKWHt54d2CZiZVrbQSMJZMzmQfqZFrwUAHOjO2o+E05E2btgyReqHOZw0hm2w9hY
vjWn1EABU3y1vVzoQoY7893kOOIaoRvrnwXxb/jM6wL9h5ci4LdpAbFWOlDO8hAG
hWzvxJF+S6fAfaKoM2xx2Qiyk0gOYVzbpLrKXEgACfai8UP96N/EZNUoYxEQXr9t
qtqGlN9YPzlFE+iLozIaLv/kPFAfl9xg9+51qTjM8qFsYHoDMBfSBhsrA7iNqFtJ
4UxE7R8UOOjgUYR53M7OD4M8kYXuBIl0dOlFbzvJ6ikfWmFFWonyvwNfsuCMEhM9
MHLr9XvmUWNSIVo3n3zg6ZdcFkMJ0sSf5+bNAfJixZhlDgxIB/A3Mni7kyVDEtdI
XnQWr35edtZNwR2cUJrN9O88F3PvB16pHDOPgXHAwO5z0vgdWWEjiOjupMsnu51T
0ZRLx7bdhjNJRmjo7yYjoa5NkXXTzbsXa2kOkcl6X9yWOgH+xEtBsRmukNaLctNZ
CTlNePDH3Z97Tao0MQAFzMAH+qF6xtwUaZ6fEE2fTVAzV6/B5ZR26zs437Zyxnyh
kxsSvKsSKNUApyuzKDPmb54/KY3xLzqcfIX9sUP24CO5tQwxGTz0RtKTRbwL5vgm
8uCydNq4xYKwwsqUydN9vpXia68bXQNfwfAioWw2au2lpPx/e0GErLGg5lDBpSYI
Tz+hi1sUL28LP3JvN2pUMushrtb4+/76KP/bo2jYdXMbh/D2SS8ni/s59wBVMZBW
uIY0MZb2OHLS8WwpHqDkAn4Sg56BtcT+ngtM71209zHDQpHOwWb+Oz49qtf9S6NV
5lgyV8M1Wu5hdaG/giEO1Yl7xCImK/k2IQlHSgVXeGTkGp/4yxCKK1FPxivhXjVa
yqWAOYMreMEC9BqCQyKAKxRyDJ8inKDCAhFaYm85wd7VFOAzDQR+qdTas9rvjKT1
P7f7Y4qbLdMzIjAw2p+s32+ygCPhzTrSitcrd20+tZ4Hk3Dl6yzK9+dsL6ddTz9X
PQigyWEgQykAQUhsmy2XMRmxKiXH4VDR6nVYpJUr0sTJrGUXR6/Suo/g2W8pQ070
GIeZzeFmywcsxR9BITkxNJxu+CDHtGkyZF81+1d0u1fph78hjV5D63XtwC+nUsT7
E1KUheqHa864K7lq/ZXuv6RHpl1Q2fneCt7/dO4GNaMoUoqAWer87TCz3uwKu/K0
1MGB8zKIcbDWsdYrvcatgJSFOYO/Gbn+Yw13cqjaVstVrrz4965XUgRPdHmQY37p
aqlg1QMW9z/du1MdmjRnKlkOmMiw2Gor5TB+k7vd72ohYf17aKpvmjX3x+aJ5jlr
NFOOpwAo4eddrgm3VGd8xrIUBjsUXzJCzgsG/AmTFSLk6iBQjZs1pPsKMWfUmtcp
qRENsJw3CNd+Bu+ZhGVWeCH2K104sL9F2rJ7xX+9FR95KQ/3PvnYWupyOdvwIGio
1GWM7fXmCvFw74tohu9JoG/cdXiyk5ppiPStbGPPYl0t+DjvCN6Uq3k6Y6oACfbU
t0Rro3BD6RFelcpr/hvLnAZvVKpzlv/WiFVdCwa5LgvgBuCZRatKihnA7KwM7jsF
gKtDJ7AeUa6y1eDtPo17VJHi+JLp/tV1Wjn+yauYExfLrsa9fMlIbhZAN6E02md0
5/AT8c4+1bYQiTRCkU0Sveb3ckvVmIPSrZIRxbV5cb4RMQEUeCoh8z0+L7dL1CCF
joi95jN3ZmqizzKeraYEm2eCosGX0dCoysdv3JpCtiMw3w5UVPt3u9d0jw+YEup3
bQZwZbBFJm7V3/FrEm3A4UeiqC/8Sh6vJru+Ou4KFb/I/TxB94YZHA/W9wNkxZEy
QaE7TU0F5cA3q/3VUZjr1kMSEMs10blJuL02ka95Do4daTizTF0q20Bz+g4N2xS+
qSahSeOSmssCsbOFViJt4NbT3eOrTfyljKQH2Mzi36INmvSioWd3Cmwp/GzMklMy
Cbh9GPFrzRUBQ4WlZgrWk4lDYC/TJtbJ0UOv8ZLphBLgrhvuWrWABpltMClveGT3
2uT8iLfrsh9Y+SS+GkUQLmTVSaHkqaRq2/wvXgE5RoFqtVyYv5SG8+dRyn6I1hAn
OfgoOYaV0aIwAWmEVFkfU2hpzs1usqULR6HNvNKORQqzqbzcypmJvmdejVI3n/wH
bIzgG+NVwuwZnYN9aJfVzQ8bw+dWgJ+NlgiyiZhFI8SR8JJ5T/DK8WGWhVJqjrqz
DTxTAv55kNVv2ziBv69dF5WWLQu24XChrEIqXvEDKlLxbzqxOULkFPdkeoMcQWYA
u+nj427uNrID4V7Bp6OBBPg0WYlyxV1jkwQv9fWvRAzv1mn0Sppr/GqAh61MSIN2
qvvMyZnekraY8xt3wv5XPJA5xzOxcaCJkrfRCUklb5EP4RMsU5ZhEaB6oL3ckExj
+sSowszFWjWP69Hb2iS8EuPP0Kx87sLeXB4Fe0rnjojY5Y5fviyg2qc9GEsn5u7y
7BadagqW+0l0wSmsMnez/I/lEaEu4ITeOk+A/eRQVFHpuVUx3emHdI7a9LH3wMgS
PPONlY8B0J7xtrfXHw1NHmdHGYTKyoUvZz1mnwkJtDHLv7szKxc+XG1qsSOrpken
vQ3PEKL8sJdfUvDIdPFEp5RugJ+6rVV2IFMw1U0Z3K5HYfESy93fvq0i36fw0JJN
XeBXbOqlS0+Oua2IQ5UxOjl+OPncE1qP0SYwl3YqPAoeHhzYQev8OSjLIwnWr2v7
isWU2IXjsXsEFke7rFwjO/KTFxezVCC1uD9ZEnBzkdOnF/mxg4GqChKeRi+gB7ae
zMr7+3JglfpUYN4KvqiVGK1MmbaZdgM/8A7TfwP6K0kU8yXaDVuaXN6WqQ0GAVAJ
awYPQgpwDYZ+pxpAE9YInlgiDB74VqVVysAPAqXZjNFngWKOSj+ngvAdXa99TDTb
tiulZGVU6b2+akOW5SUsr0Ir5Xftl4xOvA9xPgwTjmjMQ2i9BZz+1MwbhmjMgIil
x7ywxTLyPk61FAUsaSB0WOhH71vgRUF+7frcGEpQOiPb1im0PbyGfdKnvYHS9jdc
a4r7ORRvfKUwPQ383xb0/gVfXrD/qvy6gQf/7SuxTYK2lcf99SwLCSIzSxW5HSQd
5sWjFenA2AwG5o039veDYu4Czu0eJpGTaQTimgwjs2yJK0gqVVynMp6kjHPEBO/r
QVYvVnHt/NQawi5XuLcJLZFZv4p+6fXQMEb8l8ftXQes48s6N+GCVilJM97VOpbo
1j/ddmuPHn3sIxhD4jLNCNbmocl20t+hSwAsIsRroMlfSuNNp5XXBSLkhDbXJzPe
Mlwy0wUDznje6/v6lf9CsWrvRy69em9rGf5KygkuK7UsjYLUUWGfCaq/+LQZG+Zf
PyD0wPMuD97gCiRYBHVbr8crbA/htwec1lscGePgWwad2yC4j6Ke72m9LkuRroGM
AllfD7XPuxoUYKlin6+s3YVVK9bxnOJBNCGlO+Bm1nVEObSOrfjts6QIJESsx3VQ
Y2oRLKhxerxlYRBw92fmaSk4dvOQvC3H/rBOSNTxhuYXcxr/7fmFdaCABKoKgrRM
4RbsrRlDvP4Hkw+Q4AlrDHz7y7XbfV76Ih1w7YaNvc5FD0aAYSt+DDL6zvnNax07
VM6TweKPjo+os0fDqoLR/jLHgFrCYMxoHLbzxb1HMODtdOSq5DQb1RqIRlsrLX7/
ZZQ3kAtZ6nRSMVTEy9W5t+bhzz0RDARqOgkRSEHHXpalE9RjwTz5bP2dVnFcxWjo
DbxolTuWjKOI5Hdw44kQnnjEPg+ZyNXy1QjvExYHobkkVoMKwOZv3Q3kP/F9g3wb
X51oB04MxMJFx9aHxPyW94V9zVQZCxBzA26YTQocv2gtlz2upxyOpTqNlXD0SS3T
25R/g2bt3IL6pGx/5nbpJaHG3oken17ORTXFxu9NhR7R18nNl9FR5cN6koMX/3LL
A17q6bvkWIwyTRrIMNkabsrxT5K/EUSTPWQohAk+eVz2a+rrOacwpBGkZ1APMrwT
P3eJA1nGT7RDeFcD7gRlMOQ28+3YDROppPPeHixq0DsffohagLyEcWa+V4bwcyiY
hiGxSvYYwa8H1LswKtBau/eo2El/CMBOBtXiCkcxqaPbM9x89QjaIOHnUSDqdXuL
ZI5RarCZJHrkDsZIeC8i7pdJ/Nr++wIHDMRWHJj9V3vcGIk1kiiJIXLtkd7QV0iL
lBf8vDExaN8PU9Y96+l2jbQz8VKLNIKy6/HfJb5cMjHVdlCHHQzO+24yybF3rUPX
vbFgVfOKmy/qO/R9kHbLMqwiPTQeZaJuagc1SX+lbR+rUZUozYvY4LLSgStX44il
3R3smYw/8e9Iy1BUPfOUg39JUK/VhyW1d8tV3zq7u9ZqAYZCkqT8J9kg+V8IgJPz
OPEKG8xPUOIP+bfYrZnuZdBGS3GPfHdx2l9ue6a72eqIQpsZbQWvhYUrgrK1DxSW
LWh6/e7RVXSCbiokJthV5wPF/wAdsgcuSHyRuJDe02x0QTvmHG28ez/fbGlIpnGl
gcOJuHTEpwWIuUlT6TTzaDXcVEgWyDOGtc4u061eXLGArzg3MhKH97WCtfG+ZFzT
lKX70j/02PQuSeggxSzlw7Qyozrsd+KfyVUDWLA8yUDVq4sn+SMqHwbpS2j+N8wG
Xf25f2gHBS4343wCYVh6URMKGI/HNV6dWvEOykagnO+INkG/cmtRZapBzNRTS5Yz
IgWmMTrIYeVUV0h1mVOOFpTVSuTdnf6RS32eo03X3ndvP/JzEHOFdfuPrTUaNG1D
MZYgxv+9UC2Wb3ZyS9Bj+vfTLDhBfTSCxnkBOLt+P+RO1I3VFLpbr6iXMYb54XsN
CXi1CEnqmJ2mMfXWK+HIlCi914lbmGMQyUR3WSO17xCRJPmB7GVz7g0LkizJ/e1k
3gPjysdmve1UC0zFKDSl4waZwgpL7cphjRtNscCto5CDCs78cJYf+GNeHh4LRnG0
GmY8ITTuAczzIViraKTPQfOZwNRY5bIoacx4/Yygz1GqqnI3YEVT7j9WVuujIh1H
YGKv/T9NbDbzbM6C5dMXQSltQ0T7Q7ZIr8QjyzN/NjyfP7arrg4Qr0UF3PT2n3ea
rWOA8us1zKmGLP7aRZMcSB6heX9npM/muJ3v/rd79xMktoxFXxy2UfSvJQeKa+v6
U3XAPlRkAOLKbAMk5yZ+ubdTsGU6cnrup7nN6kwH+ickgT10YHv85Le225xMCBdI
qM5Rww+wX1OiYcn8fxHfqQbzg81bIk9YTMoEjSzUHLEpu2VeNApSwrf1c2nm6dzs
Nd8tuIoYD1woHVfP1lklEg9SEH3vCx1ZEOcEM8aZ58Si/kJcLxN2F5Ad0bEJE1yF
DveYeQ+nVZdVv7EfNTHRimWP3FJviTT+YfBJj3zWVkfpcNhbaI0L8IxLnyW5Cokz
daDWLc3c8WRUBfCf1XNVcCTJkTlSWcGL6iQ9iiHJ6oLQJEOLSKE3/610v/3fvHI0
Bf6f9DKYRN6NpojUaS9wkshHnfMqRO/6h1cghjUd5DU0jz9b3yFdHTpXDYkg5Xag
AGCOLAVLFP3o8P0x5o85fierEAS3j6Z37btWJZYECWhkzl3Al4HWnCzeVuM8C+Hz
xXcYQonOgTCdIiVLg6hgizbtQ0Maj3txqO4HhLLl/tCHqaE6CU1rh7JBOKqCWo6X
W0+gl4+OxHge/53SslOFnfBqOc6JjJ7ySz6ERya/g9qX7w0E23AHiEMm+n+iCkii
4HUb6xvw3avrOVifTvlg2itP9mqoQbFyUctTq+f8WShMGYOMUSEUU7q1ynq3CKiu
mRMrGWdIRValnTd19KbntlBMUFbU2bhemEENCKBpR/yndnDtM3+AWr28JAkJfXZN
N2MPTlkArPqNYhNPmN1TrXUouGzzO6SXBu9/ag+toiin2zKlMgKfNg5/KQf6+LEZ
4d0dJWvZCJznGAbbnFVkBCLxhTdv6td1DelRTaXxxsA+g9ACbXj7WY066Wi8VXuh
2y/9OwR6KDwO3y2C67eAasX36tseO6/qpB0QoEDM/g38B/egBibmExdfecBpd+ci
0Dff7YHyv9DhjaV+7HUKd/4TK20UGslb3S3Cl39Ol6q0F/zVDPpxVqH0A3MWNC0E
SstkrrvdwDYdVa9mHn0HHdp0YWLHz12jfeuwqum2OzNDlGe4b3QxFvjSdL3/rCQ6
+QimcONi6KYVnugWzFNsH1+BElHiUn/6ZjSXEAg3zBhMepXVw6Zo2eQDquYCuJlB
TbeFI2HvAB0PQEs8I+Jmc87oyOh7xweWVlq88dxtHiuGK84ho/gpPdW43UXuVdGn
g08zQtrdG5p7QJJ1wJgcfghzyad9z22+YFgUDKNvNxuq1LG6FMpfOrKvMz2db6L7
pIzz/056H5odzPSOwk9sG60yHs7QLFR9OEqPbBZRekgDesMroOXV9jMaTBgOleSC
OPjzd6fcbyE7bCnt2kb/k0hPI+3oAVNX8hgWT8uK5e+QoW2vfakIWTuaA5mKWO5f
HUu80jIWSQqOZ8HDAkbarpYxdfafHq00Z88cfc7SOWcO0M2DGeMMeGme2X6k8pbM
CYJnclgQLpqeWjuJNMueYBERvXyNWCPiI4xv1DzopCuyxVx/PIZnodN4VM6qe0eD
ngHT2jza2xdG1/i++G0oKh8SVIoUOLN4XXUZPjGrtqwXSHdfGunntif+CSLpNLsp
0MGt1KVPDZmnAb19j6Tv0bF9++F2g0HB1DB1FhOlp+v3f+YsY+ZwRHjDbBfcFiWt
rK9aVB1SYee9eQSp172YPGyouDzmaPybJ5e0qiDOhzk=
`protect end_protected