`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
hVdJHWSfELCmA4ds+csnOQAALbB3ps7EiTSHEDd//nts1r+JQrRE4d3bDPRJpiX2
Sl8d+xAK9BIi4i+3ruAzYvB6kuD7r+gs02Jsvd/1kn7JYK4xBxCjtdDFjVHOTEl1
sSh1oNiYUwLuwR1yKfP+xBhqxD2Dv6pCKhH1NdGilpJQ6cvivGkSunAu0tzP76T0
4x1pB179E7uIeRplfHWX03KzEBF+eVtfgXVp2W1BGjfAe43y1pCvNYZOh1+TY62g
EgAFgbo7pAujZxZy/YSiZjUr2mGp7o83qMXyusx8+rQ41D3X6rxfuP0RiId2pOpC
6oq5Dfkx04a1dk4s8w8cVg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="Sm9DkM+kBxuxXCFA+l3fFkxuSWV4xqRc4Nn7Ji3ukao="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
m2emGBqRy4AuduN4dffN8194qYvc9UXRqiQc56IrQYMiIVQPyh59I8SYabcDdspI
7AFHnvKD5YaF6tQfxWm+mlcmMEk2Y//aUjxeiGGs+RkKgbHitJF/K7nqg1dmKvDg
a/GaBCq4Bqh0EehlN4ntP5HxM4qcvSfh5m/Coe3drc4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uG91daMWA1mGkhgP3oZKMYye3UAomMWgG80HuuXg2E0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 26864 )
`protect data_block
c9NqBF2D1wSep1rW7utzHsk2j40aow1MnrccxUTvKej2Q1cyeDDbgAml4eTSXI8z
QYgCADtWi7S8BeChdv4B2VxKcS7CMq/DaQrOy1MKTfQzfAlK0iubmlTkljLy0Rwd
qPJokL5dgHaoxHhpf4hHtkj7FMpbz6TEPKwpE+S7cAc1nBwfhGPMlT7HmlvONncM
iycQLJMcqo+9jK9pN9FTRzZcxAUXwRZD+t1DwzkVXwouG0uTDr/EM2cAkqvs9FOM
vqQplmsWumxv3mPN8yIXaTRP463ogkbef7zAKzPmU4Wg30S5GL3ZNlJt8RWlWVvg
sV42qcit435pCQoCdJyina70y0aAXJ2F9UWxh2ErkBqUaAlDAj82+n90XbakEgDx
Io3PnTxF0TLClOhvmtqIw/jrwuf1w6LTZzrXJNQgc1GwBPc78wM1VgquYdxg2Xdn
FiKF0Q3ccYy3KiwwGubHeGgHu2u0pWMq1cXmbAdWk0fMn1z64e/5JIfzlYAdWT9e
xXyesPOdjveGt8fBNc6aRQ8Hq0l92ILNAYiUx8bbYnmFjVHVqy7uhtvwksw+a3eh
okbTrT5tIXGRqvwSx7Va2X8i9516yxdxY1VKio5YXOb9or4JTc57Lg2FnSD2hqMR
Sc8c05HXmEnLbgKUZmyOQ8JJ6bMnDhubXPW00FcOnTLkn2DqzUqrHfuy+4+wMJiz
pVO3xem076Z7UtEyafzk6xkIRzNZBQks6XPy07llGmQyBQFTxzbtI+qO4ibrw2mb
yomM957krB4X1zjQw24c6LaTbfkzW2fEJworY8aUg7pn0n4iwHrObIuH+9nmNmmM
exsjQjobx18wc/6QM2MnTLttMJ675Ioq9stR2U6L4sb3NPlm5gtIs6DbE8hBCIDn
MLbvFigZtAluWxLRcGNq9+XMUa+H6KiqVdj8Q/VdyPKEj787OXAU2fcGKS5OyD8T
vQWEPFafUmCUJ5AMeS99LicX165f2JLXqyWCEGh9BIUT3FlsE1xtiGGYJa5SCOPw
oaPz3ZlIdlPj9g0un9krB6+A6hw5dllOL15vjTbWhrZ6nKJIJbLSz9pDc8zYbg5v
WNgp6F+4ZNCH56b0kIJbeFir65jypVspKM1rWwCD0AaXGgHubBgUgv94pxGb9uJ+
pqNmXQmJ+ti3vPLimVwx2n3Ivm2QvhRPBwEz8tGQAMBaYy8iAO6PN6V3WGREQOJW
UlG182WgNWneSYwRJgMpfqllcNAaRDFtP9FxRQ62Xpo3F9sIHsPkaUEc6Wcrx4hB
lyKclDrbvfKB+8j1k0aG0LUL61JQZaj6TcvDFEfmIfr/Hm5swat+PsULLBOMtMwB
W9YGvAN117+l4nmL8bCqKeKHylvOGbFJw2eoUo4KmKaQhzeSPuaxNgw/QON/9rNA
vRgPZ1KfZ+2vYjBtDE3DOtONWr7l2JmUsyD1EY7DBXzdVhbUuD+RHlECV6hxt1Gk
MFR6RtZ4qWnLjCxsE7gAK9TbGclhg0qbgD+OIkJ0dItR92EoxUh54+WV3RiWvVsI
SgElpyLBaF7I4xGqL+qWjxcPKD3LwylqggPLemWuvP4lA+hQhLpJTzv+98pX5EQP
27u6WpYkeVT3DZSBkxFanuHfvPNOqJY5U7PYrakKaRpH5Hblqx2fVTHE0VG4Yo3T
W/H5IWh8GyKgybQ2dlizSUyO77r8Ww55/MaP9ij6a43nAuTuMHovso7exvZksZKo
6zZHfXwRJ/FL9V7m7Mm89vxk5hpgyIWBgKK2kftJ61pjJtNhISIFlh+YJOhYATkF
3Hdirhzjxcwvu/nqCEX2WbQHFhq+O1UNGFQN0wJldiYjx8ktHLlFRSSD7Zj/BWR/
I69qBR7Af4OZAPfxwnQU38jWVIQI6YmQcZ9KMkHU2WFmwwb66WuLKLzqzjD0DzlP
TynAXa1rBXwbnv3DALnWuvQBMdj10VfS7E6z5jmzIv/s4e1dZ/9Ps0wkHQcIS5Sf
OBL73ziUIatXuaPVDC7SCZx2JoqWH709vB74oUlhHqR1jfVX+kFy5yj51Wd34T4f
BYnOm+40v92brzSmIoxjrDBd4jrOJuLDsB2WAd2mU4JfD+c1tcu414r9bf7XZJ3s
jtxO7+aBY0WwisPTsN9by+MVoomEBwjKWCwWTGQHzA7JFuLWE1qWYUfcGpq3eLYm
KkulezVZv8koCVFPXX2I5jd6Tol6cOxjJlmDUAfhzPziT9cbQ8a7aSrJT+mcP6bU
tAaKW26QdOLpNSuE453yVGH7t5//COTJOxFgrI5gDjG+JU30zTKdeM5pAGIrK9EQ
JbAfq++o8g8AKbddSAZaSqLwuQa7G2/H5k6UXUFzoT0aJo1Mc7A6f5CRphoF2+Fo
+8q8GZGUfuszgGG/sCyLJmWrXoyo+H0mph+JGf86lGemd9meYf3942xr4xiSZDq+
31Il9cdtYgrRHRbgz3XNbUMyuRzpHbLY429aOJqJJfywYqoKyvJDvrvsz6yL7MEl
DheqJisrEljXvvJ7XtjtmCqnoWIBiyXyqhevNQ6AYCf2CCZromQSk/hEN5YNHhuU
dSqrDi0pBXJjNDbSzQpQOUjt53invXz0S2u2w7t+wjUfWi9a8JKWEDJcQe7AvSSs
DxUTFPYtzedfQjILXHCm20grDV+CcsxFKFLlBLJZBCTy9dYiyu83KnWJI3/6NRIi
jk1bBtA1i/XA89HFV5oRhb3KFqRwvMbCjFG4u//ygcFr8833f2Ezy3RAC7l0j0xc
xGoITNp3iDukp+sYbv3cHHYInYq2syY0BJykrztJvEN14lmOyj/p9PupNSX5aHA5
dErfE2rNdAXeI3ZphKL6SZs7ezIIWXK/7SuXmxy0B7l9A2le7GR+LxxSs2lyAPUe
EaHkGVvX2/tOcwFcDAu4itEHO/l5UJSvnENRm88JXmMPx69+yvG+4DK7ODVuHqfu
KlR5PSgw/vwRa/KOQx9zQd3xngWx4z2ObChkYblEZqIy2x/FmkjkIdLP+FOoOrFV
mMGISp9RO/BwsqRQbKG2blrdc8e/s2lv9OV+HSETb6yW0ukyecejV9evOZ0AZOYN
FdJQo3F8ihpsCqrLZtbat1xhz/rpaGb5Rm//DKTyYtBIplB5cL5TfWQPChfspotX
IO3/PxVHmh4U05u7U8o8UWojGrP7Z1T08kpqEoBMc4jgvsJsv4hyGmlC8qLxIniS
CfGd8++rmD4TDFUmFVU4Sf1qdmISRueCAlHC3WQoKMtEnxVx6M0K3mcyfM5Rfocb
G7eI9c2ftaCybuOFPfTpr7YRaj1Tgeo6y8z4jPQOzzecGy3qhC2LhwatAiwG2Uxj
+W9k7iwtDcFV+mNw4SChD5zQPoFtYbL0EWGSO8Dnqd3SMd3TMzfC04ZorV8wvIY+
niiuNE2TuG5hemRrhaT0MQZUMLN49sm5mTVT7UcjhY6eYKKwI2Wu2b0wo84djWO5
J8HFWGPPjx+B5nx2LyyAquaXsZ7lGUET2ujPuA0mtf1fx/WXlHlNlY7xPcOfjnVU
c9gRdvVsoxvDPEEipFQj75GpocvusgH+wDsdQRYprSnZwtbaK3A24eLJFZQmV3Bm
Yw//HtHf/LuS1mQPpfrEJOpurN7dirgGTQmlbjs6gfIJSzml6OrMMCrSFFkIwP2W
NAyIqgYA/5F+7aC9nXwNnZW3vD2zL9ZOUqiqGQxGQki3kxoa+KDQThHXNIkCdiQB
qDdLwHkt/X+XBFYVJhLl+0OnGAGTgD5ruRQiqkVSPSvLKQwgm3SLsJdK503e/1PM
zuw3JqsRCTjLt8cArvR1WpDl8xL/XlFVXUg46xqJSoF2QeiIFhNPqVjC2O8yEywl
j109+g2Mg2vdzplV8VJCt60FhLCF/bep/+ROdAr26GRLrKYY96LL4hB8wskLcyBf
NC7WYmIAE5w6YlOpNrMuc2A0fWH686ElCsBlwkvi+NvwGUbFD9EuDrUpX8HSm1fO
RzyJiWB3EfCg44dysBOVKjcHt8xBk3eV1fviAYAh+cfwxH1iicQM1ovWIlWxWx10
yEIeEvBRT+9FP2GzdgZtMWim8ktcj84JK3Q4bokdrb9OM0wTuESvKBQLf++N1eBN
+DxXN8IgS5Jh0buGHsyfK1bOhN5BbTAqK9nVGQQaVSIsheyk9RY8gm+0V3RtQAZB
/tTo73v05SyHxIy0eZ6eNUeATD7kn5K0+4fL+5wHqY0X+NXcDD2InL2F4K+UJt8p
vrnEKFTEsxdh9D9eYVPRHe1cnqPIaelOHqh7Xvt+e+DFrGB9QYx/BX5PLGnFQ1KY
Ca432tPpDL3IKXRKIlGN7zi45fb56668dA8GtuUOsL7tTS8fzfU2UI53bwnWOAaF
79bqDRBJOb8UK9AKW68NqVxGAuCyn9LNZiwgK+1rP/vsGoRZcM1y9fg3vPG+Q8M+
1UttbGeF7/SAAg45ey6ojXN+lXHDTN91AXf2MNWHuEj3/W1W/WszZ1WyI/0I+5/U
GtDsz7Z2pZEK0s1N2AM0bvtnaMTlJ0JnTmHWmOwhdYHKugfdCxSfWwn2j3abaIXA
BUZ0leDHL1mmAm+XY66l0Atl+FxzUBgEzyzdoj8T/ZmtaD3Q+cAXQzZG46rCfiFn
oEbVo4NS9ZHc10o0ehP2CqHlXP5u87I2HA+iV6oMtUtGgrE8gcv9JR2DZA3kZTXj
9HbXZ6LTC95VMmhlaA23H2zO4B8YCr7hq6RFWpE0COXZVLwMe1DJpaHO4Dr3NLTF
I0ChUY7f6zIso/7fQB/5VglBR5M/qzPJv2jUe940YfNdPIwc9JU/il2A9/ey4f2j
J14eX1+MVezQaUNXoe+w7t/AsnLTM/bgWUoXGE6oHqEY3+9L53xZfYVbLRLgZpLT
OOPVcZk8oWuo2sdlI80lbQEJGKkYKrIkdhKqhM2Guc6duiz4Gm40tY7hFiS5mo8L
TZlgL+HbMdfcrUi38wkmgFq1GVYW9EzKrtNWw4Ua+9Hc9ygRdAXUBuvheZoRPZyt
elWsf3lA254jianxRhxe2z0mZQTh3WdwKr6mYDLM5UFqRLo5W43mfRLKIK1VKeoC
YPioOq/oQ1fu9tQ6RXjnkCjFS8WqBV+4EBQO3ZF0xiJbjSslzC9VzuDF6ZGm1c7b
UyXolqJ5ZcDpTd3mdQO/zOAQfxsCdEAAcma0nlTJRb3giRIDLbTvrzQNCrS0L2jE
w7Uy+ha1xlt7pbejBk5nDWasGfF5WZwZMTVcbvlqRpTdXjb0BiXotuEmSyd8weCX
LzCMwuLYLXND/TzG1A0g0I+SD9tq8+V4q1mvBMP+PR1uHNcma8P8uSOvbJezozUa
asyaQmkD/KG+5hNweW7PQwNSUaulM4NnkK5fiyMmQiZXgthh46a+95GURRDYXt/T
rI0VXV/ElwjAV5+g3hP4+6zo9pqZ/T+aqsd9X7Vn1XwD8h87XurQ/NtvW1CPVCFr
r4jxUUeGdfvVK1aGiXPj8vtJIziwbREbVltwdkshSfYLZRYyYul11t381PUkAVRV
bqClS3GU9/mQi//b7+4Sv3BmdS1+wC4LTm8MC405VNpZA9dUOQhMyuEdLzTfuUhO
lPTYjPKVd+Kt9Ral+ExT7B4G8all8pwhMZkl6AzGrlG1ReytIKF8mzj6Isi1RdTw
Dm35BBk8bKNLjDO+TLRUiKO2BbFVNEiyZ4R8d/0nFfBxyUDBVQEB+oCe4yizFMOu
Xdci4Yf+Qa3dqIDq7/DthPsSHlT6l665I0mIUJ4CqiZMCIalseBs+KBd2tdfOkCK
Oh+pT8I5plR57s6bISy/bcFPEpiTpUTSdD3oD5wLoIEsvovzqbxjlN+SWEL84TSW
bv9vKNBJzaLP/+J9IKIcqYc4S5n9DdkXz0yKUKsH3Zqzhq2U0W1sALq/++PjJAIy
2/VYes3eaZ7BXXF0Lq8acg3XMvolzJQImhtNXrTi+9jYjpGuLc9BejftHJbQzNUJ
2M5QnsY/S/9VrZv6tyLAch4EIyniGifFJjxHWigfBc3VfR6X+X0Z7WPLyeh5CgwA
vlioTgxweU3PkxmGLWhzDl9UM7e/dA08X3J1OeUHyU2cyvneq5YM0qY7nwqAcA95
jFb/e/1mq4EOp0uFclE/aTejjipFhYUMO73E5qvEBR4J8mgttbOcElsgdAtp1UNV
7ZeoIQlEAV6YXPJOG9ZYsJZ4ryp7/zHN2YhiF/6vfScBFwIGoMn6xSvUpHaWrngv
2Fqroe/iMrUoiUB8pLzt0c7eQgrOPm85YYfIODHl345oS1/suvlMtGCZNRwHZ3r3
Y8D/H9sGWXrGEqiWah0jzD4vgDRo9j3a/7Uoq+hMtuHFYBx2aHWidpwDauWmJTRR
JUIUsTWzZRJLPIxBgud8T9JpAknF+KDPv0irAVsfU/84zCQrZKtZDzWagVIa7nMY
CXfn1Sc1KQWUE8fsw0DS7I1OwDE4MwVz48Xb/sY91F2ZEnRTkhnesAGBvOsCYPEe
KRjnSUtveI7iP5r/x2IWxtd7R+1HZzLQY44UiCG8TnVnSr/nfrpKROYkAsOJwQSR
+TP/Cjr7E0fLRt9zxUMhp03x+9TSn+1tkxmuP1B9x9LfT1j52GW0Tv76fEcVtUSR
UQGQIVFoKSinfbhm3MycgaGt1q8OluoWTasi6CwqHbjoRmfOtXQ/LzR7tUtL8uU0
iYSvNzNYYrfYroQebWoDG3qGX2pkN709uO8h7Jl1MZN6n3s+DpZH3xDGcIulFZZv
teAaFDVsvQa4UhKJbb0SbuuVl3ENwjT45LArfc8dxOkGox0RBmrse8Uf7GitpvN5
VR4laysuuimxziyxqIaLYnXcgQv0xOJ0283eO29lD1KFV0/mv4zNCSult0dsK7yk
2T6niBwerxjJdXBB7F5un4MAPNLdq7qATyL9ES/0VYQEQKZQw/kTImQF6FttQ5l4
Qntl74i3zMB9MznwJ50QGhajo6HiSt2O5C43S+hfrqTf1QcnlQDvv1A3VJLyCZ4t
TYHnb/iUVp4REhBbvu+fMurOQhFxQ16bvDQC2j1E8k3tFSuxn/Di5l5HrgNPmHze
Pbv8pbMsh7uJes92pPPnKWzGGwop7QwF/uHLGzwrRikdS+p9Esg54FueHOSmSgU8
uqbjz4tu8Y44EjvRrH8I0k4fOpjx2SbfvnpA3RF1+DS8NeX6lLoAPV1z0NPP+R0N
TMmwRvm36HTZysw4aTca8FCd2JelFCo8eAx3FBE3scV2QrvQEtZ6WKRCbkviku4o
1zEAxkcoTmaN6UmGEI72dNS/2GvcKOSNWnFK4kzf+1bFx+u4+IXkfRtwmTe0GuDz
4zOQ4AB5GxIn12jBfNWrSJ6pXTUcqcDl2gMEqYVZcu/QMgF1vsXiYVd8UlFjePjv
NoilsIhi2kHTFG3iZtqbX3UoxihcEOHGl8pWG8PjbNrg2v5MNi+4yiC2y8WvbZ3/
8lY7lS5tQFdbAwL1gmTZOXNlTrLsWShRo8Hinx63GwE7hNdUXqB1fqvSuvlXBr3o
vXiPi7f8dtWMh5cI9qaRQ05kEiMemWgz1xdPO4myqILPO/SNDATCwWL15Z/f3VYe
z3COHbRYYJ71KG5mImM+6wA2f9GrNhQgp+z7N1ocQK1ShaVgS5PUIyLYHtGLVSMo
ecSUtUrnsq7P+89VTBW+6SOejU4Kj75Ex6Hty0ChfXAszVd9pDD8kg66sN6HRp93
705bXnFNkniLk1Pdy4hLRx3V9K4n8GHJSAKi0r5PUGTGRSgJkYrP9+/zRv1SNBtg
QEXEjayJEqSumDCAXd/F8qBm/nGRKm8quG8yUNl+JRNltQyZuuelfz+4UNWFJgkl
4iB1kMqamUJl62xiUEeLzZb/1iXNFyUM62U/H/WE9m24QDh28h5hsBlUgKHuRFj+
BI+s0POEeyp/uJ6U/JwkNNUaQDt0PcAGQ0IVGBN9c580H7WdPFUdxRkLJqjhPfIr
bjpyRXzvxVvLkmOW/e8Kg93vFxx8eorQUiaEA6tx01ZCY63PRooTZGU3DXzzZlVQ
5rLgTrErp/ru3HX6ZISM9IT6C/BS/lkwgtHwoh5e8z24p37wo88A528Mv5gx5D45
gNRpXl/T2DPa8Nl2p7Kj6+GO38ggeoKBiCVpTO6I2kGf9koF6wEfxsSOmHbS3YvM
RITfkVIZ+XUr8bVf2gX1lyWsMpuByeburANXlMArmk3TstT9YZ2cBbcRXXsbHQGn
Sj5o/1HKJUEmhUpfDw90KmFtuRdA4dUqM/G/fTJM3LQro36A5KhEeiv4aLUTlyzr
ZabAqerS1FKYnpN9ZFr5L3LH/4DFrpTunE0bH4RDNCi4hdi4U5sKm05OSeRqp96D
uPUMi3f2GN2NHWGqtEH1ifuNRSIrlzMqsQDwMIr0Yv3it4yRHOfFkbs72eus4Kuc
KprNVD6vr1Rw3wP2XBk/Kb8qd8JKQ1Im594dO5rbtD2yEWSsAnH2t8mpM5Vi0Bb/
zGoR1e93fvpEvdrrMVj+MTLRb1A2lFiJLyBM6V6+nRbZUwOsK2v85BjYDeFnLKwZ
KTYR6P1jbqy89Ez+wvJ+UokK8JkXHiOMqvoZGw0K3rLcJJv/MkrSl+xJqShP//SF
htCjgGkCl1vgGEhkto/vedA9EjDaGawLVSnVRj4KSwkZGy/5HTKMgehsUuUaaB3M
PoxTgfQxQgbhauntAbdTIOcGmtEKLjYVWJusZS9Q8lJilDff0bK5oS3Ft4rSwfv0
u/qB6L0i3Y/0Y4BqTGvmlXuTt7lFH8GwuDTH1cxdh4vQEqYsI4vQUqmdSAQ1chA+
pIWBDvM4q7FImPJKC89yasmamwiWcN4UUQsWvpcYsDIEZJ3MvTa/MLV2qh/TJhu6
U6oeV7wxPhJ2o16oPQ44bC6ctVGc8G/Cni6Qn5irqcxNefISLxPAsrXcb+VFlpLG
+KUEP48ZU798WvnwnriPelW5OhO5nkxvDY1CpBWGMyQqxgDP4NsePHOHjspa6Nv/
zVOBGAOaY/oY4rjwf8lKR8wjxyECBpAMCPRFa1IswfeaTHPK+gyUQQGUCsny0dEr
bH8mOKyt7d4UNDue41VCP9eE9gXcMalVEke8FJ9HVDj+MQ5iat9HBb5UEFpREmqL
AgBjJw5U+iyNH2y7Du5NyYNlFUjg54vPY23s7+As1Np1Deje/jMTYNxMHWGRLsDl
BH6tP2i2EyGA6e6YyNQoCu6uR8p/nunjXzBzkXPva73ci3CbXy/g/2yxutAm+oWG
AMwGlcqnm1QTKCYdjRoRhRn9wVEgC4eS043Wv9dXhua7lZbmTf8YIlGGXdPXoq73
BdR/CMcYxEqPYUh6b9Do3LrrNhSbVOZet/p8LNuFxWpJhHpg2EigjJILcmkYuT3Y
Br78TUXzDlZy/DWfFCiCM4QVp33uMJd1qGmNcirXuakiFaV6pmg/kMHcnA78wkrM
c6LI29IAdGoCDOgz1I8lhrlI5xjhi5gkIn7AQVnStTzPzLJFq0S5YWRUnSL04NFH
gitJSthP6Dlx8I4JgewBjzFwXWD+qFLXHDCNN53gPUmKmPE9S6TIpZrSNyrbjc5M
dTkapF1UmWGWWt9HzxmxGqD+8x7abBSl4gVFaCLEZyB3A+jjdPpuVUydvmGAR/0I
eCvqYfpB84y2C2V/Nyn/JTMpKbzvjba9uhUGsrP+3oC2vQEYfSPbgBcZjBuYRQgR
/tkwJQqbCzYD68GKw65Uxc7TDQ+txfUCa07QoMjhbQrsDHhLJfGXEvQ2PGSJtJiW
05sBQed4Cv2YFs4USvpmQyP0swmxlx1gNJ3rqzmQg89Bba6q3U5sUYa/4ii+m9Fi
G3sJVVkyri4vHNbdZjFjqqsFeHrmqINgSKbrBRAqBH7//Om8sILw5Z8Z48uOnt0a
gonmeSLDAa+n9YRLx7r9IkBbkI17I0IWBR5zHE21OmBoOkD67uH9N6+finL9D7rN
4HbSSwooSZSVZcwk/2tbS8XH54sanMciC2dGkFH8vfobdlSQN6fVYcihvqYrMi1b
hdd8enDrgv9E2PWEV6mCqmTN7h7TPohy5m1wNdL1SIiHcMQqdxEwMIsSu7/qLYIU
GxDYwyFyea2fn9z8DGnVgffTgqeby0zTxSUvVmsvXpiWY3KcBmdlaZEwzU0+M2qm
o8wVcVEm0gk3DhgvQpDk3AyOvz7hrdacAcPFcLKurWaPsYhHyp/FTJgetdwDyEER
MDAyWKKFdI2gZMDCWXoNQkflA4gM6fR1w7y/iwb2/dn3EXK+apmxRmlVtoOyocPf
9Wtr4R/RG702iFQC+Tm5fEQStXahCv9Pu977AXATN7SiCzg9Iu3okA5Thp20VEmu
gxzbKVaW6k0vMdoG/T/QITLju89L6n5TKkcKWki/ToOOeDiAWIgo9g+wcrMS60WP
SiKXj87+rHtUv0wegOxZ1Pq23Gzb5kOPyb1DpduVVRmUYNaS/WIJIzS+te0wYq4F
cL1LseykyUVKmbA+h8zuaa/3QSo8U+7IuYctcrBCvNqBLfd8GK26NvSc+WO+XRwQ
3xE4kjRPA/mP9mqOJxP5i/j0s5vQIWXnycSsJwUQ/7cU/4Q0+TCDL8zNBuzEzK/5
Wh3XAlL/yAI5PLaxzezxpZWHbs3Ob7XKCo4o/z4dWdt5oEfrRo4XL99oTDFJS6uM
ZLwNsDbBqYlOgQofW7S3wtqABrsPWL6LNw2DCUZgysxLkd5O0HheRkI8yuvRs1DA
4dglywEXBhGQvjVwuuVz5FFwswWKWsaegytPxk5enEwd57KzdbNocCR4A9JjvdM+
Wo9DBdIU3UFpjMTENcsCRCoCdQdP/tQqbNCcVyp+FLxXuFf/iPHQAmGs+2kahsVx
Mx4oD0ESWonpCiK8qiXgR0Z/tsGWi7kFLZ/3FFo/S3n95DtH1x4P6k1VtbDPoqnf
pg1bI2+tg3VnASiPBZ1+DZC5BgydU9tE3XbQc+iqYETSMGMa+c8voQ9Q4+FrHQTk
VW0+pNJfEQzx/XovbBEiTRHACn1ycslFLNp5zJUnCugOTezhxx7fyB8dRFx4Y0U0
McyOtdM51Bd4qglSQYN7pLEzgyZLWu4zUSEV1tWGIm5lWWdxXuidNy4QZhFdnSFZ
Vv/nYYQ2ipbJDA9l0OV3+T/rUQpUcsma1WdoC9fbSO+EeprGs2sk8hWj+CdNqI8i
ENWpv8gmOn/G8goPGyjK2ivQlIQNtVyJbUA4hAoDI4vs+EedCnfC+DyIS98xfMyr
HYQutPASOp3VHLElToWtAeNMb3XVucFY5jlu7eDBDL6mefaVvLUvlNvODsFMky+u
GhSJWvaDsNDO6bZjiW7pf1bSRL38t7+6EF9MZ13Hl5CQ2xO5HnXw3eRIAnl1nLRs
ry0NkFS3Jl7LKuDhjTq3JAoo+GARDvez6Ino3woYM9BlpJaCcwXW/FL2C+kzx6HS
D0IOq9FHtGvyMRTLV+03z4jJW9aWfQLG63HdjJbBMzhKB8wJyRi/GD25t2IsonC7
LPkxzmkIKIo5jTnNRla3Qk/IaBrr696lqBFH1adaCS1PCeQJ1QIpmxS/DHrPz5JL
r60wZE4a5CLjxml59ECW5x0EcN3IcCeOCgjO5wCFOgjDCriUwCszyJMuDFKx4CLU
yJViNt8c5kcSvBuwvDxVbJgvFkDo2msDjWD1yrZxdOyfoY67OVAjQnzCCXTno3aK
M6fzcnT+C4WoD7k9O0AmwuXErboVKw+w0a2u7r5txwHZiPOdnJ65bsWpH0IQpXfy
JtyOMEA1Oh1xFqdve+CsPkAZK0XPmv9qAyapgpTHdHyLjHZeUxRwgS/IX1J13phO
5zDWKqzqa2uhZHvjJWAA/t8Ve+x1pxK1dIjHNkR3JXhPtudmDPvGs3DmUeblDz4U
pyg+7wbpPgSOZCSxvrJ84tVhC+lYDEzlKINM/jcJUp8dwlq0/20eRtVwAPDc5PZO
hWqd019Bz9XVnMowCRz3mWmSqPx6Uyq7ZoCdAVv0LyDd22F74LLZUubPLcOtOfC6
q3JhRZPn2pBsrFNMfA89pCtwzyJP5xvwfSs9OH9k5MCkjI8P5Ao9u/0XCHyjvjl8
TB0f5NYDsgU02YtD1D6lbH8vOWb2UbOSLjwWqGIvmUNdO2o0y1BMX8WvkhFDYldm
/uQtp1ULK3raiaINJSbBd/yofxV097capGlPy9ffxS0Qe/hLCP4O0G2q1LSbOLPG
olZDATAXA+gr3tq98i/k1gNSuY949S3kju0ykLwLThy/DPluvVcjzbd6hwmb2tTv
RhQGOy8XAorEFQY2YTy2DwmeZS02dtb/i2m53oo9M5U6JVtiR3k18MKZq9fcC5Pi
L+/CtO3Y2JLM2eL5754be2BlahuqK8pqPvulLVOsQm2DPnRZL6sQ02fHI9+kvsTu
VpRj53OwS2/F7hZiYRTwvhQu97CycjZe0VYTCfev1mmmuTIP/PgdfG0ga2IaVu+1
Zog/MlYlUsHjmoFPFG/xV1j8tarZslK5+eIy4L8QnQOmFIWr4d4razwft13+qCim
Hf2HcY7bKVjGesgP1X/aKQ10jRi+/vutf07Ipo1E+ANhk2ECSsdTOcfT30ourc+z
qC1zhYnzWiKhmiZGLRDV2+ijEyKpI9Cdlclf3tgPpxJ6GYRpzNROu9Lab/3XwMAn
STuOVifBsTPp3zFGf8Qt/5uAgHu/5RXyjNu/kFcQPnvgJHppX0XhfgKFulziPzE7
FFaGbXfnLbHy9zqKhhphT0tHESLvOasQx3aQtgVXl7mCqrnuOnuTVc4pLrhNt+DO
6PdbPdcmlvraMGY2qBA+js++m8ahuKJrZ+qQdkKP2qi7ZLDcnw2LxSY2mqPCdu6J
ekm1ZlPdWPm+oOEZ7Ak8DEvm0U57ddtrxb9PLmwSKKvkdxG/lkHUAwtGb7G8mn5a
SKUCRQjLaGjgGrB7JMGBIVe9fhJtdUnElunSVRsIMGZn3sid+OvJubFWNWPwpK8c
NtubAY20Q11Yjaj0DDEKWF1jkq7aovPjZ5eeC/p+5DeoOzt4WxKMoSGgAq4GCW6r
XrYYUUfvrzSuo1B1VV6CqZwqO/Tpg/6dFyppqSJE/C9tIiHgQpUjvRIki8vrsr1E
dwMi3DkJEXaCs+HOWuZMzqsoilUTlUr6hFv/GZkqRNlxheb1muuzHAQLmmw/R5Tu
QlRUjkEp0fLPRWWpLCkhn4D6lnrn11BmZLVP8zBLj11xBj+1Ml1oQSwybeumeDzC
Nfm/WL0pQk6G8tPhkU/cQbHy9/T3b0jsRHz5krFeU4SRtijTYOcppcLYaon0cEqD
gBJSISMdK2ihTpMEiAphL0tXCLoI89tyxSFHbn0jUKtI6XH9Ph6/Uz13SEmNHTbo
Zv2DxE1/3BGsdzV0WsN8f5mTql3Iho+toCXaD7+a+AMVSYdBKXfLwU+ekMk8gMVa
MuhcOv70Ao92GGEcQyiGWe72dawvkW/LqYiwyuQKHKMMH8O9VcC4jgnm0iugwUPq
zI//v8cN0H8EWNhxgw5b/RThMAJDe77cHaGtyBXnjwqACYd72uDlFkcSSO9nurbF
rnNKBps66nneJJIB4pBC5YfWYP0BgVn1smtcFbAW7I6iTb8jrwpn6Ge9p7Sum4kL
gWZCWFJF0frl+xam8Rtk7dS42AmTfyYpLjXnQlb8AjwVdf2OaAPgbj7K4mUQ3owS
g1/5c331Oe0Az+b8oRX/tUQpScTDJQXoa54tlsivChczm9Z1697ENIeqNzj+eSue
9mc6zoNqT71Yh7A9xVkWAAdySeCULHzGRudsn63GfaHRSra+T01wmrSqwB3r3PBa
SROsWNopEcKqFpbdq5m62jCzrhw0DtHlqRFda6naifKMEB8mtbC1kdXeb/0mmAH5
uFYBxY/dO5z66zOO1gA8AUC+b+0ZRK/3e7MndoZyoQ4eF8eMKmMtpqv+ou9h/MWv
7pwu7GLZW/ZVWJyyXtP1TBj4/f6MLehs7eJ4cgkX28dQnneLbtYavcN9Y5z/HAG4
hKavkduw6VszxYvROhA8TzMoD8wRwFZv+cO1S9TY4WbZWP6eP6BX52keiT5sMMGk
kjP6nZEbDLxG7MkFvJcrL//Zft5siXh+6YVO3XTOVZ2ZQtHR2fflESSEtW1Ka5dh
31J7XW0o90RYtjH3vFKV4rgIDYbZFCB/NLHmPVOpEf02t4yG1XtCbMjqvGAkFGGo
I2k0eAsofyy6sOxael+LeZjyI1GvK+mwVp+MTQD58GRC+1pxgn2ryNUFfsgym0BS
yYbXF8Ln+RCSmrowAe0YkiCTcoo3sLDtqtEUge2Lfjjg6fxVFdSUEaxIHi4gT6Cc
WIMmKmu3KR0SV/ZBdgM6bEwmUd4oXWx9Sql7MkyiZOg3d9352BjafX3tFYRGpo58
2SSIuKauMkREoXEtrKc0u95Dzfbe27HnuHv6iLghU/7+EVG1bct2u6CiPmwrnC11
URjTw0jZdlweW6wh9yH4I+ZNEf9SlE/Cu6OQ46xTu5QZflVncpBL/d4D4BGjBBrg
YW7nJG2mCd6pJAaGGI8SQBUCHtousmKzgnbX7ydYa2Iql5DIaGMis3HBYXgSNLnE
b501YKGgHT9GxUruq7cr9lk4qx8cWG2R5U1dUhzgHwJYJo6F4CdtEEqBvZRrArms
2hSCDO4Z9iQxNaaMz6l6qXeqj/QbEz0uRQkp61+xfWxC+hMX6Qbrp5fseh6JX6Z2
G3ax1/ZVaEGAFVcvvF1NIAppwDuHn6fbtOLyeb1nDTjTR7DQFFt2GhqrnHD2y3dY
v4c3q3JzgwoA+0rJGsVO9O+bpKTz3zbt9hbEh6eww/dYh6jtaLlNRTxkLW1qI4wL
gIlx5cemxFdjuKX1IDoSL8gaNykESuIAmDbWdOf5uFsEJoF0n+iZrfICO+zeHJP9
vsUFzlfHZs52WGV3xjy68XZZexwO5xUA6PnvRmVKYvI8pUVyBaSP3HTPD2rsdJiX
BP1egj8wD5VB9X4Jl5kXuexSV++Gy8JNPziEF6MB/1K8Q8dUgwxfqckE9hfq6NcG
0EZmpPQZg0/Xkk3Lbk2ANJRdrr6yrsrbyLnSWZhCrVuyknst4lNV9Pq/8YFVUN2u
m0NEDCtmfgta4MNaU1yrjuTKXl6FU9LMtL1RpC7dxeT/qMDNqzQyYNPK5MnzLqqo
bLWpwACXgJ4EhsgdN5p/YUmXzZ84rigOjCRSVTYiUpdfpeGjGkQQ7JBBM6wo0pzy
ccOVpUq+ClVSFWIZpPUlP+Lvmw4PPyA8WgxrbhbElX30cy8naWoCD1FkfplHxGQ5
Dca1CZBSJODqg6JPMIX2B83t1iLeyQvEfzbNCEfGSgYmSfoGZdRZj7mmFyvjLnuO
Y/qnLDRqKpp0yL3CM9BMZI6jZSXaNPd5NDXXYb5nPWL1EcUNG6hKxLvR4OONU97G
5bDSXYnGEmvBATbKTN4083s7QRBefvU1iqM1LwidWJjiLYRR0gmHeDlykL7ZCIZK
WK7hQ7c4CEiiIlRuFQP4IxVSaXo6MEE7JwPg4F0wX8dSJdTI/7jGUenmdxWnzY8S
Ur3YnPoRyutKwSphoEZPNPWMPe5GLT0koiQyOWRc/to59gYp0o2hOIZC8VsqSWha
+mJuwXoGLNZMG/HO10aOhewx0w0Zmcw0oQ4DIpINYE++ZGydOsF0mWUps0QytT+i
Ha8XpgmMi55KMxkJoUHGbNFe4mOS0nkbbeEn9m0RwUsQZm513f62HBQ4L0oLPF8r
0SfvBBQSS/06xZ6qn0FzIfiEcreitckFecb+bVYb6Zfs5ctKOfDau1xpp++QAlOu
eXMxJmcNaratJ+3osl0HzxsYJDKwRZ12Rvu2nhi3Z+yu/24itqIx5fRvj8pe4jLv
auqK/FkwLC6Xa1oEqNLxjC8pU7v704YfjJmOVK2ZjTiPKjDZNhK9PtlE8TvXF+Bz
H1eTLpCINGjkBJAgcUUfsxV18H7o2nCUE5+D+YAEaEH2NZ6Oo7IBgZHEpr67jvS9
RMzQeCTxemfjqtsnJl6gvfLHldGexRvyVIArd+KQmhcDdBwnWcsDCAzPk14zkWWA
kFU++8Hk7mSIQLs/bxckpJBuORD4269C3P66Z3gp/bARhLW4trXfexd/KIBUvwGY
KP+BYl/RcVzScirQXc0WwpFyLnI57ikGoPbHfWyOd4uISs9zF71BNLJlwhGnFaoi
lWjIb7fDpC/QpZ28zAP+wW1JNjsWP2c//c92SKugPGj4/JNNFm17bvBHuJnZS0hM
JFSoWQiR1OMdGNR/sbWoZ8Oq4Paku4T04ElEUada9ENUQB/9jon86zCMDLQMvyy5
7i93fnU7YPVs6dc6rgnY+elZwia1RO/JlJEsJFfn9FUEELUKlJYiBVzVragC9Wfs
oBB4Je0z+aFj7orwFhluLw4zjRkTbCgtVZ7+G2k4/wiPzbNiXCQzeYsscBDZKQWv
Ri0S1bXepBH4JCGoceTWUF0pT7GnYgrge9GEh6jr+3JTZYdpqjCArwEbVVF39EME
VLFLE/EN5eFqD+6Wg4ZITWqZBrFE/IR1QV12Q4WNweyMMINI8u32CTLKjBoRKN2Q
+f4DB0YffmOqUaayQCCo5E9J0MaV11E10L5EMIHhUfdcQTs74ADXI8g7t0qNiGjS
M43GHj6BECfj3Ws7LoqoRsl+75pLQ5/asanK1f03r3TJ6gBAd90Da4xnryVq44wk
GDkBI/NYXkg1/02ZCXyGbyY6joLcQBCHskUoZqmirZxYXKujigUx8+qiRJK++g2f
Z5jaNwjSK5BsxCJGxuDmVLpQGhUIXxThFgOI7+0T+xymJS2O3cZPa4OUTokd/9qU
0761NFDRLev6AireBifVjc1+cBOv/vdaaolIoOkvAJhhOq1hmnUfyD5PsGfLI66F
ZiSXNmxVUfQCpc+XdaPBevHngk8XNuxysR+Z08Tz8uf5j8vIb/We+WEE8B4q84iE
6OedTtDXzzK9yQTdXVQqVslptR/2KXRKPqOVikXZR9v9jtg9k2bvoAq1FNgc2w5A
8pDGdPpb+QrZcwnPLzGvYlSjTIR9D7JkzpptLiFxGH972rluPNcDjMUybesfKMoO
mBE5yn/ziIjRVNIOjhU6+5bNNGFWbmLL80jhIzdv/96J17Dd8J6tzNFzvSXSAUin
MDVmo8HiVzmYE/6pV74nLVp3fYaugt2Fi4Xo2kRMsoub5f+5Da+y1gNpVhhGKwan
HYoeHjXYwE+ncl04mZD2WWUhdb/PQ4LTXo2AC6afd339zZcNqp7f+EJw0kJXI5p4
BTZhK4eb81WbmJW8nb1WodVG+04sJq/HxuSI3arYZ+fhjPufsIM4vo1d9zPPMcQb
XUbx7nbTuETbmKRh0X4l6d1keGwGRF8ent7az6gYkMWWOG9lPwQggJnwxPTRLpw7
HTk+dWqRI72aCxTuZhSWrAM17IvHDqjIbIGKUETK8SkcDVzvBwJmDwJf2wSFDswN
JY+Y3rbUFpGqbAWruZuIcuaEXI74AaHjUfX8ajibwgeU+qvWAsHUjJKDPHY9ytU4
rRnC/TGw1ooEW7rslt6f3nPYoi+CqrbijcOcOysQt9viDaQTdqDM81SV4ViAFQ21
P638QgD05yPu2R11MB9iClCdiCHJsuNiIzqh44xggVgsTMAUqDL2C+TOcmNu8+2D
5AoolZhDCDiIlSf/t49I8xbK4bD9wO30It5YqmgYcSsXft8tE9ldcfVOV+Fb45wO
RmpNr+Otu/VMFof23zn3X6hBTIzz903lO0wOSRUEvH06O8Sz9L3D5I6B++pv3KvD
hKeFGPwRUMErV2/dWsLQpjIzUmiXvl3FCh98vDdFh9G4PIujH18qbCyYE78JMS9m
iq+5XScp9wC8Ol9cf4HfiXKxXZWJeo5VBua+dFn7k5lV2v/yFSCNcJXakWj1JXoc
VycjICAAwbOQ4xLHgYv0uJIahGoFvtjkbkqKXDksfWhhYsO+Yy0mwrH5bl97GEP+
8Amb2HGgMwpEbWXlJYSOgYyEFr9wOASuMAIHQBXv/HepAGAdHCTyIL8lnjjk7btG
Vz7ErkxxQhTYhXQIXMvFB+FccUjkcgTJCqTBxXnYfiM0LfcdsVd/cha7Lj1UiOwX
eYqKutO8saxPrq6ICPGgWKlJzsepyH053vgzBtK5zUmQYrQrI/wYdGUy5mbMNufF
OJPf99EX0EBNnA6I6mQcMR3lUCM8X95CeHQLDjwDxPDOAbebzc/E0BzGiXqlcGNH
DneydSpyUfhiEUVFTxodEvG7FxoM9EB84k2xdaQtGvXD27oYEmprmW28Bqk7tvgF
Lx0x91TNcOabvfXlhJ7bW4sLpe8yGu1HI2x4OBvXnYx8cgBqnS2SzNzC23XtpyjZ
EKcP+wtxFUOUTYmZ4q/hy2KOqkj92xpCkUQ+16Phy4IaFlPJOwyC8GzBDVjgLUcn
wTkbzhVV23Q/fdxh2HQnkT2QqKm9AuXdNAvzFOohMrqYWmRPn77uYU5HcuFvUPer
Jn1kLeH1UnWenyIlg9h5Us/b5h8vALrfQmKNeMNgi2S6cblgqFG9j6ehFJXLrPBE
L3tCYtjcNm36VPG+/DYw0qv6VNbs0moPwk2R7voap2CplN/lrA4PZH7yAicVjw4z
52lrwIQWXXaMYcCfw0iPRj2Tcwj/vXiftHqypYaxcrrCWHT5BXpgGv0N1FOwQ7mb
8YRJljFRjeK4uKvb8MsqCsXXjHTOyGJPp5zQA0LKq6NDHd3CJLZ35iKGvObJqEKZ
9TERdByMRQ5Qf9SzAqcigVJx2sYXoG/iL7dG5peqxxHSGfUCxNvNtLjFE749G+Kb
DQgUHmKJmslUgcbUXDt3SGnaezVoXhGAy1olLmD6WRNjkcyu2ivBboRt36Chcr8A
EdxUtCVT9ZcexbwrLa3d0GJH+Gs+fo0gg1msIua5AKDnGYKvuVK0ZTGfsYIuYFEq
6GewTb3jhAxkcVJnkevOArlRQiPDOdTtl0jeUnTdpUMLxmi4tA2BHfGI/ielLBqL
8UIz0nnGECN+0c/bfGOdq94KAdPhNVPadNEaBHDaBxYQUM6xQVPOWOJ8Es7Ana90
hjp0xTk31iR2ST4u7M5/v789DNw/7xvTPUXhbJcTozXCyP3hdmMQ+mw8P6igUY1W
JqW86oaw8tvuA4hV3Eg++wMBS4KcjmY8UTluArXzf8e4HklpNM9L28sgfUcTWiS3
pAwv0j3YE/DwXvZLCS6auVXel3Sfhvo6DWajdDn6aXOTwvkAghhY5R6hpngyndMI
+aplzPzqNzKrLT9TL2IVz24Sz86+TCboloZVLKK4Jns0IxZDmj55rMayxTaKOrxi
lDkhmnDBHcujQjMqZyp8/BrM9CSE3DP43R4Zvgk8RTJTMIc4wJNIk75FwPvMs0BQ
giM8JcuwvbHAm61opWbQ1vt/C8sRhW7kurEpMX76uQxVPy5OR6ATENP1Q0Di/a+v
PAapEgCOuiFsk9TrH0pzd18g9oT3q95GvMIkP5qyLdDVa8P6YMHkBAwhXDl1g2Hc
PdXideMxxzLqmFLzV4Qp+o7OpJW4GVVF9i9SvMVxLMXcwDv4Ph02XXOYH4asWacL
0KKyCItczkC9CAjTFeUbtZCbwLYOpoijT4dq5Yp27w4yVJM9rRG56B+ot3JfdswV
kLX+MtPDNmugOCstD5ygjzh1zYaLIEBWk8+XS89bMhnpt0/dg9Hq2T06huvHhDqR
5nEAJGQ8uqtdBdscUkx8CxpfVBE7FDdKNqjbmGqyLC3L7ZacqwAQE9KRnK0Z7X6v
eDHpJsIkJLCPwS1p7GA+Ex5n+T4BphTbPPQXARZSY0jwFqCDxg8jM9xw56cunfpF
2tvMpIWnCxXJpkMGbQ59dO8dD0mux/Nk6xba8lzmuSM6i/2ahBDcsXRHohscSJTg
X8HkaRNmIIPTBJm2ifSAYlj3XqNEzamOaze8PcGc8mXrOQlt6bycCo8fGCBY1uZX
37onSRt1kh8AkVaspqpsK/SuOhW7yDd/qpV/i4lBqSBpPvZo5DpkS4MLVETUf8r5
7394fBtQmOeiZ8tNA8J/EpcuPm7v7dTSX5kL386lfppu43kU2dtTKYDjvxOarYhD
MTs+Hj0a3b3xFUGZwGTsWm/73FyPKtTtm58NwSWZ01sPUySS8wa1hlyzCengP3Vh
//JdE5wmjGvSHGfRz5nQTT8i+fwUJ3d/aXJ4+GO7TsEuPwIWJjDrssfqJvh34J83
14/Ta5f1p76tRGE4fFxLk+DG18WBbe5SSVXXyfWzgnyp0oW5GPDNNEFAeDwuL+sz
AyQlohtK/l41e0NmPQXQqzWy9cMO2U6RuqlzOaML65ib5xYU4Y+cPxKbQpMk95eK
kmdkV8SWZaiYnLX9YeIiikgQoPF15GsDWF4vRwXFj5HSrl0kWAaJ71nnJ2i9RPKi
QawBPADwL9hYLbYwNZnIoyFIE3fofmL+ZDvUqvvGKLXC2ZUTLtnDMzQegL0MfKS4
ODKqASMgiAFmX741GmSmeQgojL29eaNlb+EWxjIf8MKp4Bqbb2yKttmH9LmaFyk3
HBMlPmYqi642K0wCHn70nUnSJ/8qo4t1B6WsSC5Zd1lGQiHru+StKPiQ0PHqA+pL
XsK5y5QhYCpvl0ffvAghtCzZ6Ev2ypFdtuU1fYSeWHHFDl4+QxcWaOHtHgBGCrWJ
0kjMF3WLmlW/toUh+ZQYLdAfb5DPg++F0j/eeE6A5EKy3zOFUDzEapIYxMX3KFG3
k96GCSyhWbcYaTEGKCb5p9daJuu6K7uUXIox1UNONE/dgZExte1MDhKqbOGwAA90
gS9LG3ZV8Kf7wuwRRJbOMI5kdJttAQqlr+EkUpCIM9KlI2M2NC30MWk/yLiLDO6h
4UB63mXg1JDAZMnraVri7/uy+IiOEbXCiryz1CiA3QwIY45+eqfg21VAk+/cKJJZ
de/wx05F5clc6IJ+XyLS62z1NNlMkasp51fECNbuHFikTisGabCFcPMmw00DamqP
l1m/3Wp37IRUmXrYVwgQ+prrgStCDXnQCSbyTeMJbhy3tLmUGyGQ0Ew6Dwr9lSGD
APUbQ94lt/ouZDJYej98SotGDHxwxGb1lEs7yHgyFhU0a9M1OOCeHntS01YyUim9
U4ZhiXl0WeVQgRPumygvSp3fzEUL0KEi+av0f22NxaosntiFv+O3RaAp6OXZFaTh
0/LiLRbSot/7fUEi+oPox7V0/ywdLpzH3l0ob5oxzHClAfitfwK//xjqWPW7cz40
uyvtTFw6sgZY6IOnqg8VZKitlvWTrULEjwheXNO4z0hQyhjmTBr8jaSR34DnXjho
EHc9wUwL76evQ59ayUfydM04NXgimbR4SVfY2APfol2DdKw6AaTrPoWCqChg+ncM
gOyKWvE5AbzaNyhefIhjNWQxzW2LtaDNOCYkBSPAaB05F92pBfwdQ9qtvvPEsBhR
6IWjydFoDnbHoYypayhe8lVYhlmjXYx6etuF32+h8sZTj8qQtwwyr0WdaojNGwi/
qPZ3PI56RaOET3mioYXogzHpLMk84/7xVPl2ImnBFESxxqBbqHV83JBntnEQAOsw
HVKOVpeTCs0jJ25AcM+vXt/mJaKjJS08HmNAdDAEAU07iv9ogcqvJ33WepI1OET6
FZT5RbiCFAZ7GDx6JkQvACh5cHJ+R9JZKb5rjkPCxBurkTyIqKmRFYwcZL5VysaM
eC04phgJ49MPCYVx7ENdskK2+/VO3w0r8Ii1oE8q8pEOAOjB0FElQfUPdwKdil1I
nZQv8iPag/6FeuWVNPMwW7xNmDDuh1cTC6Vxbq5LBS+sZKCnOdXwRkmmQXHqYtVy
5pmZVqFNRuVe0mDnDn6PrOsaNha8nRyH1xlXoZzqw9C3WPb/krTI6wf9uodXeTwD
CfLkHiZD6Ive/lnAvQamq0hfgRw+XHeyQBYS/m/qrj562YQEiMyYzA2BzsZkA8qI
ZhJ1+5byN1SVMxP4aS7aBONA3TySY1hq59Dk9SMXe2VAuEq5HIZ4R7V7lQe7+ZkY
mDBwGHbyMsgSkPfSuHUNaCHfRe4XPBr3kMkqoexnVvlnpQ1bNEZ6n4YDs8EC6gG8
9tEA/GRmgUrVNHK0/z8zAcY7OgLc5ba2v+40qNATdzqLQDnnCBeF3+3n+dSmPR+v
aMNkbfwoJD2BFAEqKN4KD0OJYkjn+ms2VB4oK4HkMcPCa20yehWagnV5uW613nzt
4q5arkkKqdO1PdarhwGxoRxZ9ggu/IUpZq/chVGkMh2+e2iLCt1uCcmMu+EL8Axq
iPCYvw/EzNZEpm98m6IjrQNo+OyMgGIsQNN2Wf4qUlGZ9/qx2Vg808kEElHFHOYR
Qwc2tH32NGb8q3B8qBrKD3lD3EMlxCzqExMNGgzESo84AhDhtVAHqMB4iTia7gph
WPKrmtVO/f07xemaXu1zZH7p30Ov/0SBu0YpbWcBhVNd7621Ok20V/ka1uKjxtP7
jKJvb4qS6p1aqLvGS//YH7hhIOerHW9cSzGxzgtyf42JGKEF58hJx7mRfny0VpCK
OhM6hQ2A3Q8wKwXb2ZoNQw0ETe2Q+7V6qkvbeJHtow/IN45yFWK0Gd8AY45qUR4q
cIiy68Me7TaztmYiwQ8Ap2W4pEmwez1yzJL1fNgCrf/MEJ0V1+eFLJlw/V+GwDCH
FPFnXI/AThbSYXbvrx8KagcuFWfjjlqFi3DPzlc4RjTukjLfaI23cf5MqtUAUuWE
oxUPOkHQQU4z2E8uk795zOQmm2OgFTkBS4PiuWop+MsSMoW4gGDFGbMphlRlzsmm
bO1Syc1w1EVa7h/TCPY+gm1t+G+s5nAsOFWemDZcD6TRRAXx+f1KzG+y28krwZE6
oik+G/eJ+LI874gP7378scuLMpTgxTOTElxDxIs/73XHXkde3alj1E8mqaJHSIRB
amnYZDNzm+kyl6YWXiY+1NJRBQT4zccHvm2+JEIwglNWCuUsynn+Vty0Gam5E+PX
j+9yl78hjPCLILyNGh/SyMG91SqfbIrzEWKse7honO3o7kMgISEQxUtvxsiETefT
zeyAj1OKHXYQmyzXMLwSvuP48R7RuTn07ACnbTkRqZPItIA0Xodde559eAMkfKl9
AJh7eM/D0k7cPAQzN5c+B+U9/brRnofVg/IYVcCqYFTNaPGKhf0QvH5KYIhxi24j
1NPPaPhXu1Q0k3HQ1ee7nbIvvmQuIHotLhxrZXN3+mDYe//iXPTcCuFJHI/+bwFA
MDN2MGa1zw/HLXihdd+GKKEiDg5gOrIMXOiB/aYqCO0D9OzFJZyTT1+MoYagsAuU
q30B6hzavku3xdodi+rKvTZ4qLNYaKMGVwwiuIElXxirll8yJK1NVxYY4snwpjPK
LAvltK5xSrjqOzkSC4x6IXpJ1tWfI9qyZhP7wqj2uNIEfq4mS45PeI1vBD8q0tiv
2oG0l5b5hCsCvvLxRx4j3v0er8LRZB1yVH0SRjcIterNjOH/bwA1WR71KBiKSuxA
SDQx0o/IULgHPiBlRCCSVVngzTCAYZjJaf+EawhqWjkHvPT8NNlkxNyh9sJQRBLn
ZXHVieHphPwyqsXlVNXKpS/D0OP2wHUwfSp1s6XTl9+XUhyC4Yg4/PNYDxGJTiUN
VTJjBSgzW/nI0r5Bj7wqQATj6sd6nAT+9fW4oJQM88YlNDVdUvsxK/BeSBrUuFTM
7/ikPI16LrTJexrJwjzqzLJbJfv0CCmIrmjTlfcSMfFSCgMyk1OPl5OR9CP634xD
HerLGysTBtRF9hwMWKP8nFKeyPsJfrjh/WHttfMIff3yeSlqbOGWemcxmIZYOkze
VW5hTYAhlofzCLWlOGaADj2mvcdJi38rTsSMxyFcicwk3gkF/XwJRvQzYCRpHg0z
r6gJc3zF+cWDeo0iDzHqwbE3DyKSrVZdX0zHrXWz6nYv6UzwERRNiu3Lv9yKsOTS
ekUwO0a+xg1Vb3ulj8qjXnrq0V80IFii3WEq6C+z4OYfe73MqnUGy2D9EiPKCkCp
aXHFh8yHBaeDfX12KKafOpSmmbimBIXDL8iXvrc73SfWgX/lum6RXoLZztiIOlaE
tIN0Iomc7eT62ZeJB6e1R2UXgaLHT6aVk7IjGcOeC8+IRU6W2wwKvVBiKtnM/HDR
njWTrsxZCiZ5NfR7uTXu+0VwM3udmVWMqJYD4UDpkY2SSrRI8uh4bMyoUaykkVoB
CJtNIrHBvCqtICEXL7wdoMiZOU/tAc3Go7qCC3gffdEJUb+wGxAN2sB5TzwyDu4Q
CVMFYoWar+AfqEbNfzVhYOsjdghaVh9j2yhruRArmfaCKxsA+l157AT/kJPIimxv
cKfSUXsWSVMXKHL+zxfBV1K0+N3JYZz93MtEdctpED4rQmq8xu5f7RlrjLIC2V9a
IThW32gTwYFAqyLCWave/jN5u4JpDou41kAagbcGpdFDJUVLuX7HljpPTUi8tAnI
wOuzXimpwaH6gspq3xO0IIyc27WruRZ3V9AOIpzKrULJITLoCairewg0fnXxG6m/
mg/bswJYQGq3TgmEnk6z6zbBG8AP15iEVf3FNpI4iQsArWY6Qu2v4WN4WuwXXNCi
tUonc8taGSuYxW4ck76lHMnEugcqo/YVHfZwV4RRpe3DASuSvp0q8UIVImsUXPVP
FjykTYvPWXN61GVPxjykX+IQY8SVz9Y2Y7khJjfBY2dtLzYO5GAPaduGIrV/YITI
8Ji5DMZRB8TbkGjighm32clEt2eYYKzk9a4a7CbtlhoDj4+04X4W0L+Yjqc4nIbG
AIPINlt+JdEVqxc/FDo8DsdcVzfQ/Y8vGs8B7O7m+8u2z6iwQ33V5LjFqCdUr3tY
609LQv2haPMvSBBQYTDh+CiRQu/GutAR6g+Ro0vMkta6DLEqO44ejxUVCW/8ubg6
CyZfZjdNH3kUzs3leatTorR9JUxO8KsOsPKNBRI2JPjQxEjlPV3WzpMgQIoxszfh
QK3lYtQOXVOSnKu9tAG1v2T1LU1BYZibYfU9GurP8DE7p6LkluECswWAtq5Fgykz
r5OWxiJZbWX1UAEfqkC/c/FpKrmePSRA+dw13/BZtmUFwOT1i22DPqIOe5uH3LdR
Q8fwPxU1X0YS98Kiy0wFAoGu4XQ2MjxhWDSE7gDkxjZN+/Y4Xr/TwUKpMXOsvtam
Uck3kVyssctxC7XWCBudoax1qyzUkUjKRw9UAumnK6Lrvj0rQr8O+89v8c0QgIN9
26zkHEjH93NtBreRK76ixT8BP0EJA5y+0B9tMA6gZhX3sfKu4OaJsq8GgRiHgJSB
Oov6o3yaCBwEWTCUyg7vv8nGcbZpb0zlhR9hIYjCwJ92+5eKKD1Xggghg+b1hUJN
uPRX9alrW6rp8OYXiwkpskTWOXq0Y/I7fA53IP7HnPUK0zfdq6ZsSdAsIJApErsH
PGXs4dORfj+2r/V5xJvWDvK6LAmdTrpJTGM3AqvUX3QMhohEzw0MiXolE+iHPSZ/
sfgCWK6/Eniv7elZDBQGW+QxEfHFcF5Tj58+AukK+qG/UnoTMY7wYdDtHVlTe4wF
5/T3wdaPtq+X/4RzeYAgMKpZi299pUcXCg1/HLq2n+0fi7gf4uM07X8budkbR3CO
iFBNo4F+XhaVgOPziS20Lsmx+iG76OCOSnDzQWT/Vk+B97evB+Edv224s/3etBcl
zbI2sjFVFMeK4QKSjhPQwHXRAF6eoKgEEzT5cGIOMgZdFk5r5QgXZrSbc7CS/Gp8
qxqCDEaGDv1tjUDfZ02LlIR1xbORxaRtx3yyqcLNFvItdK54oGxGbp1OLIcyAa3W
XPb6HzMthSihisur7vSXoctIh3pf3Ui0RJQY730Ual7OhbEwdsdO137hDHDHekkw
mZVa9oTjsrUzxiSZhZcllgyfkK+nEG4d2xxbSu9jzndBUL6/LeyA15vXUNShl4tk
28bZzR+uTrbN0zepk+rK4jQ8XZBV4DX9icPKakdB5phe34Zfjl3s0LR56CicAfKu
jjKAphH7eGg2QiseF0XpCvhM0bH0ktrGZOZQH1YltOeYWczAJSJJD3Ar2mpA2NRt
vBSUuBuKXwQGiAREUpQtOPZZHdQ0UUj3W/6xFYhIiNBGaQuTYvVI8jB67idg7MRE
kvKfHUzsfJ1ERJW/mTVMkuyHTfpds4/YyvRSCpQsJe6FrHvLwRaPZKdbr9ojCWaK
NY14dU9F/ca+vi8pVc6xGRmJ+ce3zjbd4xy0fM/4FGcsobkS5Dk+BJH4ZfyeXqdJ
VKJ+PeRY/eRY1dmEGTmC4fmNphGUhTKWt4eBOUkbcFzCX4fUxDlIfk6+3u1qP/EF
PJuAoWWiAd5AZlxWEb/d8MRBDSIcFVLdG7iT8x3wlNWvLMsmsBlTMBxxHts8s08u
ajVc69QnMVhdZV3GZw3KCDhdEbNY/z00F76vWYy11gJvEnmqqSW+i7bsJNZPMYaK
ZRmVB7RXDlnXVbyuaVMBEpKSlTsHUBDbqKuxrWeRBI8MZTVeBAhulhUKWDk2E6bN
Po0youxnJxgTzaTWWzNlwOn4wW5XrDO1YXeDl8uJvkNAqPOopkBS2ASDqFD3/P1R
AvT6YhAHf9NlnOgT/WINOKJVayxn9b3utk6cp9cDXRZyCZ7AdaoUTsnymvPsYCuz
waQ7qoR2CVoMjjrTNrosNAXpiJzxH/MVCXHrQKfQRbA2tUvcLoZ1XS2VBTFXsXeZ
7Hi1NWIpHU+IpMLiXVxEhlo+uS75ex/YxELRL4hLIiAHi7b5VDeV8OcdRkEfrB7B
L11G0terfDd7snUBMU6a/eCxBrnQP1LEi8rQEhtdZv9lhvutb8XVdG3fRBVShJ0P
s0DPYqvdFFqQ97wIIsoBeA95cI7VdRHgoaqKRNIkU2DO9UQMIVcW9dP3SC9OHQU/
6boMLho9JjAaB8Cam/Zv4miD1CC35B/pfxXIGpvvfqMrPkmUHvu97DjJ4W4bs4fd
Tq9kLxVdu8Bn9hPKp5POIZ62qWnvA9HdPcykSRFEO3AESz43Qydw8KiCN9paJSMH
xk4ahEITlt/pj+xstf86Y0h5coCw6rGLj6vsBBMFqT72ypZJ6bCJLjP1vCY3bKyX
VKo8OLtkx4wTlbbd53Mm1LraueZZ+Kd/inBia3s/WkcFsmW/XgGDdWG9DfvrLH9u
Da2+epc1qXRVuB6zefRAWb3qcvf4MAJ8grmFeNyDYecSLIOS4u0LVGhXN+vtj9MI
vUv4pV0TomZld+MUtWJ4qj08mlVkc/+SqusmvZUqwvqmEu1riNY2c2V5o0hIPosU
8gRKnFC6KkETrsOkJCD9yzFCVqBDWfoaxwvESWsK4IR+cJ1HNUZeZFSEQjhwJTGJ
ZhKvJD25DMgUiXDU1Q0xnu84EvdCDaTVrPWYm9TgAWLaswbe3PK6WCajTN52q4Zt
xte1XuFcFzWKS9vRtU7VTmg3VDHZRZa4JMhapfxlxQ1I37P5CdpUH7YfnJosePWr
Mgqif5w3flwRCrdy5Y6iQcl0+WgkYOaOv0bYmZ8Mu9ovLRBFy8Au5GTktPE8z1rc
LcfJv0yVh4/VZ0mK+k3WYmL+Gq5FqABpGZPqOQNHabGHKYZBSSaGEPCCvOqfRnHe
/hpcsVXRhHUzMsKZMNMu85Zw9fP9omOZgEPPrnTzsujRHW9ppVigr2l+/auCR1dj
N5qEHEL0Rz/USyOyI2DOMq/FG/6I389Y9D05CJjN/HDz6w6UVbI/JhchCry96oSp
Ujuq99EooLJepkLa5w0Dm87HfgBTbgWuaq9pgM4xHljVU/VgzGUkOuyNuTeWsNCB
4GlEZqJhlVQuMYOIAgSn+ilmqKzLflSu8iEsftmxmwtSi2aJ8V3OexGn1bdB9LUn
0S3eM2VE06Z2bAE77dnVshJDoVf2kcWk7Z4sU9RfIOaKq7ov1HF75gYbNpldXUGu
Kq4HpPqe9xyVJPNGvTLsnSZz3NTLOjbSEaA70gjptue6HAiftviBjiFj6g9ioMbv
436sDCUWNnneGqcFBJXbeLyvGLAXRxVztt0MXgVSZeF5iBZ/7yzlox/DYEH4nVSJ
nOaCFA8NP94Ni6zYnYQKXnpWThzL9KJo56W5vhKzs5Kt2VMBoUI3vFBreze9XtdA
b/wW+ss/B3oCCKemHyAffe+f8aXsVqtC6OHTcqeMZlQ620qLN2/Dh1bB/A/xxf/J
97wuMa2xnJuyGYbmC3BPS84VQLTQI2bPrX0dZuCYQqPLs27+iReNqDOrJ+5hdN9P
0YqhFbIhx7HT5WhhIzlBlYPNqXC8+KRkjG95s1WAkB+7C8hBd/UeTrRyLvJF6ZfK
OcmeKzAcw8xuJi+RSUSLuimaarOXrny8wR2Nj5qUiOrKkqShC/hPXMj81IN0prjQ
ecdbURzYeKUy2HAmQI6lYLlwh0fRGTQU3C2p5lHWcyJYoKteHMGTKeB+20v7VqLR
4OrEYn2gur2TsRKLakLKaygCFCUA24SdvHl2UcjRTCcgYuR6BXmvHwG3ZlnvnxVE
phNuwAxGwtvYl53r9Yn9eU/DbfqEosrqAVNMNwCb+9yDm5wxG3uJbuuo0csOK/r3
WJwW7kVh+JmJHGNhtGGCLucPbAKyS97g82VHchLbrLb2zmEQeDy8LU/qSKX7zrRf
QNpj3YPSnP5yTJEe4Sq5KhmcmtJhcfgsQNLO8/reMZZhg1oBgbgy1BdgeV/VjWYo
iozleUZrfdsAdzmpWSzj/ZhlsKJEVONuNSUF5elJjo+PWkIfovAAl2pxy26Q6mkB
2qMp8BzuBGuNHz3s+QgZUeEcy6vQ5Q/QEK7gXnCaCax9TLPX81AZlMhSeugRwAW+
6bB09GZY8nO6jBo1i5OBxoMq9S8/oSlRWeb43u96mGtcL7RdCjUi9EMjTfekPIP9
+0BEVqWeMYrVSx3wPREmTjdXBcqy9Pqqxrk0Hm928lR31dP3SHXFM9t62ICJiA1H
A/ITrFzkFR1UqB5UBAs91KGqjsE8EZ77msu9deuyh3WTDgN+ooVGjbU7Ywv5VJsc
fgNgiunmdFttJClw72+Jq3U9fJsEBu+gvZcv8d87BVqoymnWd7PoSVHlUrGOCKjK
PKhrKXRhn0EOdDXzvIT4ukZ6QSbtDk7XlYJ3LaC/ry7fIX8rlsIpsIHWj3cZxMtL
ypeHKCikVVmc/7K6V5q7ge5LnMd5FfkNVaJqXkJcVCnpgETLMRsaGI5GY0NWnhXY
N/Em1vyoTxTnDWfVNYSKO/j764oesspE8JHIzJ6O4qR0RrYsmXgl8rsgbXYLyNBe
WSpI5J5kFasNkiMXWPQioLfZAmOf+BOpVagmzXpxXm8zDVyFWX8UOkcT2kMdbj7a
qqeyeEXUIAMHUFX7kFSY/BwI9YNDdRlKjC1T6sD5tJOWKyfu2JW60It5aSfxl75r
nMHiHWmMnPUVXBv3mpZ3Ii0QL5cX/1fDnPULnkRLq3I8SJJyAOk8dkwjBqjMLwj6
CFaEZDxA/1rrjxHEBrM8KqairDXf/o2hcO9LiAC/xeRAPF4cJCYqfGkwNrwb4t8i
iR28lLzhV/zIiSzxa0jkYprPbKRS4Mud20vgVjVpdzj4nuLAlRuSYzEl/S2k8NOO
H0DGC7Ce40rr75cg2gkx9c8cGyYJKcgG09j0qeZmL9lP1r5Ow46WSqcPwVrms0CA
j4mhGSnhZ74KyA9vfe97J+88wC1Ns10zIcDlN7euZpMPs98xW7uojtQRh0rpurd4
p2TWwFE0KzdHsdemmum0kWSLFhsgVJzBaJRJ5ypQbOT+HdDcNIlkgK/NsUIPkp1w
lHte64JMxwUWGzFmui+E9fPc/gWB4/v+QX9BnAenUR8OwlZ6rq5ynZARTtYMisad
Ss/O5dHVvKyGdZvFToHf0Qg8G43KTWyeDtNau7KTGAErgzuOJJKzZD3guzjEI7HE
aF2nt+KqVTH0QZNJKwG030CNvg0iglSNEuUBCqjbR/z7En2XdY1s21tnLxfi0pl/
IBqKnZva3rsmBHjePMJfK1V76dhbB20+HT6anJXLp79DaXpt9+7Nt/dfSaXA5mVl
gsAlVIkagvP8jm8ZQmJdxQETdvLgtcoDNnY2CIe/9uNlVw9EB7wUPd3rJLcRguHC
uclGgjs0ILQI3hPapfbwMpfoZRLpsPVfhXlwv5s5Tr24oqWL8uLp1P52643UBKye
agOGrouv7qKtMXlXll3EYrpHJRLNqKrSiSiijWBvYkqFqk7C3lnfxYZezy5/OHXF
nAjgxwuoGKt5IFycPDZumAhWuOVaWYM+SQQclkFh/FuYo9z3sq8w93RZnGxfoQh4
m+LByZZBCVxPW4gS6ZquPn+tCx5tPISZL4jaDKsykYrSiXTMaNpm0AvAqHsWYxtr
fao0pRjmynHrqFhgIE2Q7LJy38NbczVNrEqREwIGSB11D6FfZGNaKuckg1T0amQs
2XvXKF7FOHDucF7wu0C2A1+LFo7kygQTT5da764+0uA8Kv3RjJvbLmbRpap4Z8Vt
MkbHe0fRSL00p9b35KAw7iJMPRa6aBIFe3AGplXOqn68jD95z2TSp8W/4gtKIG0V
cPi1VSnAyHviiKUD1YYX59lHgBEOoeI3toGyY8fGjYmgBxSxgLSCV236kQm4gm+d
eHJaBWA0BxG/NZtRGLK3/QEFyqzCXUJ2J6ojC1ZEQ9twSAS/xjA65hIo+Fz3/QKM
OXLt/u4lEz6gyrrmYVzN7lfxCDSDzNNyOMlCiVFWOmz9j/LWzf8l6jJgm81Qv1wm
L0Com7jeonLdmiqyRo7c0nF+H3rsPR/rqS9gOvqh7kqtBCGeNuUOG0gVx8/xZJBc
9cuxXiuhPeTbrJlti6IAhoIIqOqHNssE/BtbP6Q7HbVbz3T/Fto+BWSTKMq7ZyiN
v7vwGaycR674B2xi+gQfFtg95ZwAsYoM9ZAi9ktoCeon3cYtrzaN/YHNym94rX8f
h7nhQaLOKPxVk4TJtIJoydyWLYB/USBXATwD3qAFXD7lr/rTKIdjRfHVyOnjeQtm
fz69JE5/vUxW0p08VFO0kNMFAStkFA0cnQpI71LkbZYQcrY9UHtKZSsdzJC7/ekM
DqgIU3lEHzB01yQW0g7DbJpZ6umqtjSptQe3lZ808g8AbCNq4izy4FY6YxXz/jpg
FhdolVxFpS0tqRHTXDzVE38A1BCffvu5gUCNdyRtq20tk1xIuZjrwmx2wGC56T8S
+LdlHZ+P/Z9NxnMzrbH+IwZ1+tyq9/333IxSqRgsFrC7H1/VWE10oLAHp+RvgNng
tVem1FHO1eITDdG5SRCoW/RwCZ0wyKuAVGpTNxSvDj8+y0H70Kf3Tcj2Z61ZAM9f
4L7X3gRAGYd2u4WSU5/SAdAIY5YuZMBlq1c8if9EWwWC+781aOm3VPw/4Qvd7EkG
W9CD1/yyzOTEqVPOkzfjchmdCtWCDpZNgDMrAzNLFDnMy78j0CUgCjs2EgJFUdD8
FajvMrmIPRT5/ClM3QuiEukNoGbUjBfklSz7Q03AVFskmZkttsg5VcLwK0Q5Svfo
b5xHSrT95ZABMNIMzN4UPGUK4XESqNUhPH7jRXbFImLPv/4KbNM5YVjER0xCtPQZ
XWjwzi97zLn+GBUvNpfw/rI3JeWTMSMP3pndkMdrzVsoEmc6bbzcZWc5e9hjl/Gj
VQZpbFSgqY6FbDD7DG9rUjNnYmh+vQxi4T3v7ZF8dYoaFGcW/V7Y1NL6TDil3/Qb
dbomc2M9Bv/C8DvdA13zZh6fUQo7YtH7KhSIn5fFJrycbY/rVlKbWJh3mjd3kUD9
0W0eIA+LLuCRSMI9zLGTIwajMxHtH9/yhO7j3Mmra+IOGX1rJkMBeX7HedM+bSaG
mVAgFrxTz0kXomS9dV3qsUgeDGsIHdUXL4D/frFXOlK9RUybfzr8de3Xwnti55V3
9O3/+PQt23ZSzdrtTmdEeXZW70bLSPz3KvyrlaVPj9UEmD5gVzAJR1G0M8d6b6y+
9nwFb28NUH9P9/jlpQlrhLU7vBYqaiu/c1z3Z2dXh6X2xhPQeGi+ZBncsMdinBMM
GEjCGnETJIBXCHetsGkeiikmngJeUU/MGCK/quJ76f1+5X6WCKsFMAGFkFGhu4Pz
q0c7I+mJXElV85KzByV/RCc8d8B3xEBvmJvQuBtEPoCh53MVDn5xo1Kx6yg5xCb+
pnv9AaU/eTFBt7VKoxZTlE0je2siO/+CQVvIcn4KjCwXZ11Da2W8EZZxLE1j3c3G
ZThUvvrsARzFJ2HCxio0fMTiYyAAZPsJlqc6oi2CyQgZp0KEuUtkY6H+8I7F66TN
ocl+akIjbYbFPq2KIHNaO28ZXqrpV77/H1ZeF9A1wKFF4yauTNcTTryvCpg4FpPX
2Bp0xZT0c7WL7HerwkEI2tIpPSd1Q+hfBIuT1YbHHP7/A6gR4IWxeCdfkeOdRQiC
BtjtSIKPboSGD32Fq3VK+68zunx0+OBxChPsl+ki/mYgMu0tFVIEOOY4JjW6ILYO
3KGJFKH6QcBUj+9qu1+5x6xbQnW81bIb7hDaH7KAGbZAvEGOd6tSSSrY7tNDa+/I
5TKelJzD3hliTSTmjmtgkSwEv7CpYNowo5/opsM/GOSaCu0/JUGCn8lKnkI6PaTG
1o89NY+BzF2btZ8NSim+1WXpISLZ1mXrt5zClQNW2NVxeACsxydlOj3p/jQnyTgb
KDad+ibE2bZmVc5OMrDg9PNep1EW+AZfHTS6HyuYT7Xap4MVws+BqsElnsiB1bQk
iewBqqIRXFmfkkvCi3ekMB2I3Y/fVrzAOO0X9HLBGKNXSkYjdwW6HeCjiNjysfTx
y35C7dEgsxL3lFCuXSwCfHOYheNLNOkaGAqdLpYkF3AKOVfMztVMlII2kQDlMk9D
h9tunKn4fTuHqWzfZbhH92EZbhwyssu7akrvKI2kO62wtMHQwXNdgDmVYFfb6jb9
WoS+fJtACux2lsm/DezbJqHNU28KBbE4eYqHLRpJIm4FNPqspx/E+Moz7sp+tWiK
XzjVNrOHDt/CvgYm4nbT1HkG2kGL0SAQ+i9gktcz6h2P2Cf/eGEn9CUZIgioPSSn
Qt5G4Jg80dMFRScjGAWmvGpTXn61EUVmlMboUFEIqwpcixAyNlxnVPakPtwXUI6+
qHR1OPrGMAk0Jl/pd74/yhU32u9ANSeyhKwNUUxy5KFB0UxlviI514Yf+0j6IJN5
gNlZ8fncS5w/ZM0CRaOnCc72nY4pGzT56yrALkuDcAnTQqzIkznKk0c64LZ5IXMW
yLCWCKPU3oy1GslJ9tTBz3om5RHuFw4JvnNmkxKqZqhAjltqAq7SOjVpgmF8QuTG
s2YYu9SfDXF9WP0xUV7DgDdQ80h72oLsENxrN5+mU44ThquP3e1hZTm45BWdzmXI
W3wAT2xNSFLX7uj8zEwPCmJHJ1Nj2SHxBQcKu0g0hUH+CO4U96ZizTUq7GtdDY8R
8Eh7oFweGejzQ6W7VsBwYS3H6l2x60dq8pWVvb0T4WKV0h/xDZ2o04wI3D+Skjg9
1+bFwak1htOnQ+5jGXCopqQh4pv+EAdg9ITHSoYttM6v1cSpDnYihQ2uY2vd4ft1
0wvuceBY/NjIVwnyQQMm4nLZMJVwCnu83zt1EmY7dqHXs6LtSl7n30hL9upXlp0O
+d72vQEe7Xmj2XZ4UWhpB8THaRRqt8wf+BksNs8spN6cuti0tS2yZcLZN1YhPry8
YokW5CkwZCsaWjgGXvPqPX9LsLWCkH5ehQbwTujtFR49JI0YlPYAZ94HiRhzgD0P
wcGiOWJT8iLefJ11hj3+Jah/qSO3lrq8KzZJxXmDzxa4VUTzT3Hw0KPa/QdfTubM
e7xATmK35tzSJjd0r0iaUOWdv+KOyipsSRo3uCu6/K3O4zMs6vdtc13DJ0xU6r7a
sMDgkd9dvWAMRF1KThqErOAD0KN/7Nnf89OgWUNSRpoMEVOVZqEJtsx4td4ctLhl
bA8h611OpKnrtjNwTTVy8EmJzSxUTZdshdWHwbV7/3rJncwKu67R+FcZ0VcieHWi
aPHaSvqIunk85kPVNXsYsUF4TLcFzLroWYBr3aD3h62VimOYsakPLa7e3kk/XBdU
VXQVf0sgNBewjwi4xSXuMCTIACdektddCzgzxWe/nIatjCZC2ctmgxWnd1FlXeGL
/U47ls9RwgdaGFeNoEhXL9pcU/bHIY9gBtF2OCtcZoXKUywI6JFMMgoC/SkYZqA6
78zuJqjn0riN7tBa5BZTXqaIvr5xc+0UGJxrqtaZjPd8xwJsO4JtUfNEONbG+QCR
vonojKTo4z2E+7pAZpozVZ7s2z1mlBYggM9mnQxSKI14NFu7gDpG/b76KhJ9X4Qb
rhZ1luhzdvkEmHXOLkCzjubSQQ214qkfjoBY+AUzSuEGEwd7JwbKGPXbf4IU6AwD
O6rQtU+wq63VbYL5JB1znJZxbMDSES2sfDBYrOBKTu11fz6eCpXAkxx+85YJGT08
CJaGjQfYepqKNi2Vc0T17wSeuoc00vWJVa1eMmTlWv5gkkhzttDiu4v+6/L5AI53
ooYKkhuS83N4eE12GYqwS5aZXjyW6mX++Mk8qfH7d2vDEi7D/QpGOjoDrt1VzRV6
ItFfytuwzFgDO3B9mpJ6RssbY7WdEv+/uFnGcfPlwRC94L164Jutr0TtV9oI8BV/
85Ccq3vHmeooSy2NXAp9TI8wKgFdZyA4QkGRpiyS00POfwln++TXQLa1D84O9SRI
HcMwQApWK7Su8+7mtK6t/3Wmp7R0yAeWvXo252LqGwdwl/FQ4YXCAXBwde7N8pjJ
cP/N4dhvy1cvyBygk9YnjoV4hgCeHgSbhoQpFpdyG+8TrobwoAjrR1tiPRFfXxft
+neQU2+JkJikhbZbpvj5HwQ8DvqOikAzfDc2qZtVM4hxGtrFpSQXjhLA/mEvfgam
zfsY3Xob2HG/5ei6zRwMJ+pq+1OyjsdJCjHGiP7tW2Q2RTK5oo+kyL+npRZfPC5X
HiD34MQ+EuarO7dZGMipIgxIrfSiupm2Sri2RvCdKU16PV5D8vznHqZgSxc5yoM+
XqC+KYF5cv5nLY5Vf85tHKg1/x56vb/Hx4BXfn1GENMLdbEEIwlkbNMN/JQdqkbS
u0dmdhBNKqRs2N6sy8kTDagZnOxrPoDPxtxA/lgXTsJ1Nb/IX0Bp6D2771dYihcY
Ty87fyKjfjISApjn4PxhXT43OtauYewzwRV1wyQKzdD/bzEXAIijzWBj169Jy1lq
8YRz5eCjSpYHqRny89Mfwrytu5awMUxKiLs7q5Svf+yJaOuhiqiUUHYqJczeATPj
gPQM+wA82QplGlR0G1mhoa5/t4cWjEFQE7q7Y0OVT11uSs8fagUsOdXL+8p/sMyR
q049JEGB+KVUZ/0bE0hEavOB/HK/l5WCrPx9iZaAIysdv6CtNE8z7nxAJDOpqHnN
eLo5h20SdDVKcxnPXsChahNypoDUKadJkf9e8LuIKESb5cOBMhDcpIUovQEjdsj6
Mv9bc6MdiwaVo9jDnbUfDfxYsXUrMI1CdFDA4g235rM8pY2nb1ELlYj8qc8YBEJf
tQAXtWsGJZJpTtrKc9SyM6QqzKr+jBpKEKTPZhaP3aWqu76v9e4EjP75wOUFZyFX
+Kx7TxAmuKQf3RA3KKL67BQlV2xw3+d/AmhS/igxipBXlFo/lpLag1GXIbT2Myij
pF3xTcK15q3o1S7tzPK5PtrgLaGE+K6EVbc3+4kxwU6qwiqn0RkGQM5jcGBqQ3dK
X/TsblOv3sVGq3Rok0W49z+hrw/2GOKKrVmecv87q3XrDnzyFYMghUQFRem5h/T/
p/U21lCjRe+vbXpbR5IAiR7orKsWMs//Oh4jiZS2XvDJ/CXRVWYZEiLcfq37qqS4
frRbCSe/jW9mm0uImlv322ay54FOa7ZLGLocmETN2/4=
`protect end_protected