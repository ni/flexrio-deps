`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5744 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
GgG2UXwpbWAyDgGIJC8iiNsjz9F8+4DCIXP37LWaPmL0RU03UFJ1j0xaxE+3D/+Y
kAd4qVtUZZUSER0iKivJE1N0NhkKIm7qFrecwRa9l9RiikVsTgwM8yb+nKAjLpVw
Z6LQe1tu9iG32FDjjMTJEIEgQf3RKO5pxHy7IC/P/AgWxH4w/XBLkUGigHe4Od0w
Iuf8p+8aG4v2qrUMf9OnghCsUWs1XpMNzFVp/jwj0ZQoex9TAXEkq0Q0fzjJR6z+
xUoNJ2BmQe3xhdnV1kJyuNXTIGDVG+HHnAtSaglHGybxXt3LLarvMfVNN9JrvQAI
d9EzrCwSypKwdV1FooHuiof/1h4ZhenGLKrs+EFqJOvnv3xKj0AFkpLEvjDqXnkF
aLPGgZkZj09bFmfpBdeQI1YLBmL2Zu+jKNTYWooivrkHKiG1UcpGRvPxhsSAFYm1
LEz/bx9VIKNfPfn4Rdz6LKIV0tD28IG3e2j/JQ0Yt5xHh3AZEB5LAchc82yjmvaX
yXCYXagaaZ4SaX3Z4JydQTFxmaf+RpoSLjPjCJhus3by6Tow3Ri5F0C46Ky7c5OM
AkEtyxw8N4YQ+ojlicOpFwbsViSlXTESboxPWxKxRrUVz5yUCiQVAsCHwp5ZC5mR
03BpZKTuSyMk9B8iYgtzTC/6yNYmg3K/OG/Clw7cAJFcpNm9uhG6vSLHO39T8zhp
hFp+pg/teGNqHVgAAeN2lIku46hNjP/HjfnJFNqHs7KeV6zx7poB8uK5LSDx4fgQ
Y9ld3ahT5FKEsVX2nGkSs/upkTz3OgsiG4N1k5cuqOsSLULSRYgnfM9VvGmvStR7
MszBGURFfr7a7XfqvsIsuMFzvD1iflhRoUem13uDr7RBJCaaDWmQFWY245/ssVke
dcLvxRGFVO4l5+SxLsLTTXu3sBQyEA9RQdHcu4NeP8n6+2nzgW4qJ/x6Zj5WnZ3D
hzaz1mPA7YxAhNBSwJw3FIRRi2eWHUCl0GxcfKIsByfdFh22e0XkYyyK5smFsYW1
RdNdky99Bcp2SvOkcqhdfCh8GU8y5n7SfUvXKMTT1cUQp9C60J3jRkW3U5yORR/V
Kdim6SfQETnrf0MMm6UjQJZtocZDivY4QMHD9nuimUFhyRrtt68JZh5SzSYfib1+
rFN72tSh0DhgHVbQyRQO/UR7CJbQdl2W6iYTqHUBEWR8IDkcvPDPrTsqy0t9+xBz
yJbLiraZff0YQh6ls1EXp740koHdi/5RlagvzrzpEfGcKhh/1AeytTH+e6573eG/
+itu35m3Fw12mduBIJ1a2p7omDwdgvTYHtcWU3nWAPOEvhskdaUhryYF75N4Dfat
QP9UOwobDbmYWOAyXPLlj+mDpVvPPQuhOFcxf5UYCJ1Dhh+han5zkacT4RTxM0PD
WwP9FpoZBNMgNZvDxB17O8b8f0z4B5QIWmJRxLMRB8zTJXd4V3g8+/KnwDRyOdQ8
/+om4CJxRoYGjf7kmUNHQVKs1ObRZ0C1+pRc6uzIixFDX8b3nHZgZXQTHPKN9R39
LhLsbrInxI1xqrKoAz6T9TxHDAduZXITIV+hWunadqxHHimJVq4/ReY0xNoJlvAd
fgPVpYWeEM7zkHhytdcJbihY5SMnH10gSLFTXgpoi43Uocdc9s9m2GNqmp9lB1Ty
SIy17Ak0AhsMjQ5FdqXKJrmL3DKGicdmuANu4jrGKVXp7d39F4KSSb32IAIwAXAw
DBf2N+uTGaqMd6k8Ix0ap6pQNsTJzHBfAbW3uGwvwdxMyW1tPldq1KwmidM9LNyZ
ePzydog7WHwpEqqIpyn5xCh7YuEo7OA+lwnkFONXvjQu+St5Qkr8Xds7d8u7WPUf
BshPPNDwaAtrXKHMospWShJG/YJZlqYsV1saTnKbo16XmExhXwk/7F2kAUaM2kYM
xzwE3uXRUbRL+SsJhVjL96JRQd/qgsNVacGEeJZEEwwHZML46VqO2EfUig+V2CaR
8lITK8EAm7qpMyrKAmqN2a/graXuRZGN2vuHh/o9yVAecoLbWVNtr9Q8qoLnd+XU
VH2JaMSJ6H54/WLeLz28p9+/gi6EcOO02QJ4SpAWFzF1/Wl0DeeEHuJiOv/TJUjh
jZvEeTrQmSNdG4rctga8+FyAisOgBpK+a6Z/j2NukUcNcViqKZkkDYiZfFu1ggYF
/Lq1tAr2edcP4Rfc8ie2U9ghyhwB9QxyM2G/CtJ+7/XjUhwuWKus3wC8QIF24nCr
c4JcpYk8hdXLlQnI6HJ2x9KzXmO9X95Ipi056w3topuUq8xh9xEiynquJWulE5yo
VmCktH5fdiQaMKzLNiporRWzXIlQwDlH9Ezmrnip0msRQ+iaohe9rjKhPSE2FdEE
IPGyBjxWlWikvPBfP/6N02tLssbK00/knbP8J9hZtUcawkbgwyE9VW0JMBsABge4
NSmcRBCn+fks4NMCkw3pKAMXVFXLE3VgrRVY8jVlSGop80DbXO6Iu+U/jgkqKRc+
qZ0dac/DpP/R6za6rfxtXe63bZin8/g/i49eepg8cVOA4uEcNB96mxQdWBcB3rYt
3R6yIM8A9QNKzmnpdtv1y1YVJyg0zFwJeEOLEVZtzg7G0uELtPEyzkuSIDNwdeEn
DQ9yJ2KBK373/5zlv04XUga820lzfU82biGARMFK5YT2ha7MitOVT0JHmTbFRWfJ
ZLLhx6W1vk/Z6hPUy+qg2Dt7Eg8TOAjBWLUeS7Qqqk0mHEhs6h/2exB+u3EZLuem
PLP+OQnZVm/gmPBnQXxff7gQnxEFXT3RTEL7k7G9PHugb8oJDqm0LDXQ6TosQ/wO
6D07+QItnYZCcNsr6+r1KAQBbC5TYzJPJNF6i+D0doupb3Ee1A9Q8+6YyPkdXLg7
koGyLoBDyfE0r/7/En28I8DOInf5TmXDukM4RUG1PmJlHf0fEHsvPRDdab0CFbeY
cqwHKK0FVm0ZEBCp5obJw8wgqZPktFE0tPJTAZShqiQshGWp5M6RtOaiLqzovz4b
MrDxg6ojwVssibk1jdsHj51DVYcYpf4zV6A5UehVxlnBV6yGNwOYYEXwIjJ4Df3p
i0gIAF+UmxpntFNh8gp/mXX8c1pgp5fwlXuWLZFBWofSmD/gOTQidN/eG7atsy/Y
QihARNPHTn1hZB3iVrm1lw8OIvRGt7NglJrpb7ZEgVVRbK1WdxlgBTPTPuB87+LG
mMT/Ny31noTu316IJDTQqirs83rGmJXqy2m1kNXcHK4lWiCGxEpvc/zRuGM2LTcl
Sorn5OCnBp5LHFnOnYqfTCkC/zQIJN40ZRYlm+kaNaOwet9I8Xf+6mBzEJ2AzZLg
WoTY5KHJddDtKvgqvow4oIzlUnkyI4TiRL5cxrCxYviryk+T7WRkmHiqmWRGiAUE
yqtuCewXhQn/js/+C9FkHJOBsc6vxLH6Y0Z+V1VlylI1rX38XOuGjN3zzmgn/t1q
RW8SF/aZzJWhK5tj5K8qPVCmCFsjumt8B3vNo8+TC5uvBaG0Gl4Yu2oSircU5y9v
MKpNSLg34CIh8quZ/qUcpa4/CwcouIaCI1anW5Nw8AIjg0BN2Sx4tPF8XEzBc88d
k3zbwXBBxf3JSNmTz2X6wJyw2vl4R3Pykl2wBqllX332TojuDpBUKCvkpPdUvZXY
0zK6yIveGG7FYuu4phcq52XZTx7u1Iso5zZEiuyTkZSYCnAj8qy4UrwaKDTsVMUw
lSaizMnOB55YsGhORj63iM0XQ2VTAaxzMzLmpzZTQYnAXk61gKxE+OKRp+772a1p
ars5cybn9+lt0NqqYgn7xl+ZAaly1QQTgRAZB8lrD2O8XhodfQZp8ZxI+XTle/gR
zTEkdcCS7oDAka0nJUvFCKkY/TxbYlZZZjd5OStOldD5CQdAXCFmsD6qhfHL7Vq2
gDHkm7CZhpqrR0PhiWJJuuxPMzDbYKF7h2XFRCs2yHMe5WZy7jnCFFw/u1Hl+xiP
SdYqUZDvyVUgkBSjE0VxIVaBGoaznU2vty5jpifdOkYXYyy4RSc1MdYPi5cWas6P
d9KxmF3V9E8DzKtMKWRuA+Ef27dknWP0KQwXvqhII+JYhHEuH4uyLk/TuUqZ6d5a
lhex4bqM+p/PAMOfiOb2A3QWXyS/auSWzB5ds3H4+sLvpfB+wYPvef5NVNdtNTgk
Qewc6OzVrj1vW839qvFnqWUX4QPXgApIYrfKtI+c6ls27GzdVHEwhRlud4K8Lbdh
Lwo9da/NoWfzLuRNsn9A74gFuujd5cMvs+TKOwch3UeGhI7hqbaug/B5T8rcMtlc
kCwtghREG6DMzONp7Fop+lyblhPTGBBve+Cx2NlcR3jJE676HAfxseqc8X4nNIAk
bgBlY/n1+dA7zmJNquEmiw7nBHSOiP5j5OwME4qUVe00tJjoI0MxaFFjrHAzGvyf
44U7JixGmdB2dI2gSqUbJggeo80+hmPClHFM3i3Q+uIBoI83AoAKMPZSAiB9e3sw
7NdTbG3iAfDzhh3jSN3YUBVpr4wD8ehX5GYea7pdkt35isKt20xnMzXeGadSs5eT
QLxJYFjmmUzIo7lHFTcFHP1E6b75AP4AdxZ5KwhGI16TTbdXQ/A4z5YTJSZtxOhy
/VWL4dQfgdsjU3KhhjsO81ynfwtGHC+IsCKlBrcDpCbbk/CHL5pL/jdTenXL6LQ9
gaj8hmH3ZtyDDxEZmZFP2MiaSUyHWY28pTov3ExY33EDmmnyTg5HsUhAZIU8MLPN
ZdjjG1+bkliASbA1WRMdo+PHGXeQtMejnVv7IGmNWfI/ytmN5q5vEkYFZW2lB7f+
mzJjDjIQpLXAjs2K1heMG/hympDNRsesOGmcuVhaaOVfNSFD7SZNNPjPTxWxAELj
XQb2/i5Zdh2v7AhKPgA1zy9JZI3YuvtQaXHeuxmbKxo/rrV+7c6NshAQ7dFvLI+2
IKamIWeYeclcdjYAEgeB1VWbg7xVPEvkoID5oSsHUiW8bKzhPlLS/z6QWZcxcVCF
2dg4s/sVcrmBNuZ2YKeLdH+/kCSRTgd/XE0niFVsFkKC6GCEXc0dws5kEOOCr8uA
UaGmsizblgnhUQULvAzcNkUeULFJmCpQpSEm08OmBSqf09mZGDNVq5NM+r19eBWC
OUTmf3f97D/ecmtEMywhzNG7d4QgxW6BYI7i4nWCDwLTZ1Cq1ncKp8pv8yCo7LhE
LdGUIPdL/p/3UywUgetUobviSyNSLo9nUt/AqGq3vsPzbZtX5f1ED7K8bbBiYSKy
vtVbJNlM/eCkprSD/Z4YBC8wdagslJBD7PEgN1pm9CxV3o+rBysWXSBIvNPH/C80
gjsWbkGaVkG0eYqAA/+ksdFiVsa49O/SLqM2GDRRf3HDwsALEydy8p4W4+9Sr4e+
SgmzTh2eriETA0Kg+H4BovNr79xC6AfQ/iZBlQGKoT3BkbO12HJ3NDCk/WzopA78
+JrUMlDnY1Jw9rO+0NEXTdc1TubQlSHD+/UqiPrEWk/Jd9WgKs7hrVbGHzi6YHRa
7be+FutFnkq1N4oi2zG4PGSqSN+ml+pGEvl0F1BAb02LNCm8WJwwpNL8fIhjwa4w
7eJlyb3mO60/UJLfHDE3DxJuJ08Y85Y/UR5+RYVevopvhTOi9Omeom4ppmuuoLVx
/hfSm+Gw+Rv9UBRYVXg9wU0yjXJBKea8jI3QhXY2wyGWyXAEJteBhY6dNaz1ufXq
anLMalPq87oB5vjDze5GGKGm+y50afyA/2UGCsaZ5P+8c+2cmt/Ab8pruDtv3Q5y
TaZoWkHOl5C6rVDQPehdGJzxPm1plv+HBhY61Onwinh6CgKJdgx6yvh/iUzz5c5Q
7zFHCye5HT5W6JjFy3Z7VNW8vZ6/T4xtk/yC+BdCxWqOVJ6I43CR9tTZOrolBaWW
JjyszPtlG2FrLiOe2UymR/iHoX64n4MCJ8knZ6c7AiWVHDjHDZgZ5CaAKvhaztau
YYf4KiDKO/ke6NJPpm9XYUYS3F/vdVNdbugfBIpbhdUXXeEm0fYNrJ05+DofTxzl
PUQausxe4tpr8hpIwdH9V+llpnsTmOjq2CoUZFAKzzHKxG9Xe5eyABZTXufAjPs6
KyB2qsNMkfA6jbbBraVkaechull2dcG6w6raAWM5DPUfF/jI8/1a/LJcXDyhMUKl
tcfVwhnsBJpok0h+oWKj5ekE7t+3v0mRC9g6uA6c7ieb42rkIdL/Sc+vHbEfNnLx
WilR0ijFSp4Jc9RW9ZQC4s8YbgxLqs6CJ8hkPlZ7yrEms5AbpZPI7R4ZCKI3dtP3
L34zHzJLp6dCwDbuk0SONDPbI8Y97uVGx0my7HS+MoSggw66PNesSvgJoWaaEiZs
LBUCptkiHVuJxmKYJOh9n+mlDvyjQkKiX+OOby7wxFCpyQxMW126G5SHXMVsVlzr
/T+ItGAQ9oVr335Zs80YAwjf3GN24PcJwVIDx7NqS1PkPP6DSQGA7QFpueH7UDM+
FzwkJFHCiUAdbQKTLz4nuy6qFuzQ1bYwo9+o9rwrzFm2vB9OVMKIRZCDmxrkH+nf
Y/dJnds4TeLtjDKVNSx9PR5CeTA7BJlI8n1H7hkE1yy4/ZsDR5dDELMckhxp5Wwn
4Y+juYEb6/GnX2lbyupAokCSVPx1WIxe47cvHPydDFf00OKKXzYqCeTp9tDspsgM
qzGLO6+489LM6P82hJDw7a+iC0ddbuwiUa8fB0eA+v84sjXh1PnaGSc1lCQYb9+M
kk7hybkgtH3xWxE/Df+RfEEZxVM5tZoQUlR8uTh6wLj9NDrkaEpnP0bHm9TCnoWN
Ajwf4sBA/iABbifzl4ZeNbtyBBRUEP9rubRYrgkIBA+LzoU9dcbg4tLyCXvgy9qR
IE3l/8e5htNUhonWiQCfW1/Te2KawORpR8E0GGk5gUPV2HX0NHDwJRDG9lZdoWCK
zGVyETLcP+RcorbbG1iSB7JGrZR/5n4tFRBmPaU3GX1zbFAkbfYOow6yslkPlYbu
Dg6fcRbxTqFm4NaU6ZbdnlapqwXmIxvby3ajSmLqx3WANx9TtWG2jRlvfGmAJ865
p5bTC4BN0RMDLO96/qf6EwDyKaMLwUZ1e/HW/D69tZCg8BVETTePI1QNTXP8RvuO
LyUn3KGTwgNtB4iOOQCqYrUqR8KxCbZZ5wRrXfZxz/iEQTgNvN4NGtFVySfjP2e8
U+t2EqiLopbnzvb9lBB9I/hLwmcVlrkBUA+5yrUiVGv4w8PA8rJuJsnrvzaX0SNm
NaFVi7wgIGupVUTIcT0uheisA4aSJHUSEssgIJfzeQIZV38yljezhwSFRpPmYP7w
GELyvIoqjjjP2ihiRTaiRiK48wmRnvSU0idNwNDVJypK9Z8tuE39ZcCkQ6MkWTVF
95m7pledPaWF3dc9RseYwny506MAu7ggGycTxoD3LXwNV9HvIwz+t8ec+AW5pcoh
fRpAucUZxKa27Z6lhqCRgXLm7PiQIV2+wUEltzMy8PPjxyTCGdwrlaSG60wyD8nl
k6swLM3ZSY1YboNR7Q7Y4G1nbPZbxzvnfzcLApttDIg=
`protect end_protected