`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 41760 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
akBpHK9XojjdOyFTP3pOwmQwyndwquh0hwXz7XaPCuRG7FUr92Wv0gCLf+hrjQzY
Wdpe4DJjrduvQep/I3pCiO/K7RZJFEEvuVFMuUHKQ8WnqphKV7AgsR5QtDwgrLrz
7l0yuOhCUAxucRLoPuGuwj+l6nQjHkzg9MBixZ9spsu7YoFIDKIfsK4vTmqRp/NQ
syEGZbHIcInKNfel9Z6K62Xmt1s6YdMmrnp/gsmrvXE9U/T98QO4nsf0sjthS442
GwiP7QSy+t/1rRE5XP3acVsKlnjdfFHLSkxvNc9PCMcDAdmGd4Qg9Wj3rmYuT5BF
fmLfV7c61z808zFbo7rY+FNlYkdkOdJ5SFTPrqwi7GcZ7t0T5f9xc+KOecc23Yl8
kMXh/Z9Y1Vf44It0R9QuP0Dfo8Tk0dDtEbx4tDbjXCEY4455Cawuwgcf64KgVhcS
ffexdcQGyAgTXrspCFSLs03O5DMQPhhnePylV+tYYqdnCjm5MihDzVfPh7ZJjNOx
S1zTFzTG5DmSVNuxF1xTuWXUM7i8PS+shgbCH7D9RG4MjOUrWeIs1MWs+P8OMYjH
vF7BrHWu0dXHD+ENl1S7p1qBwWI5R85b6KqkfTU2p22OGZ/NKpLLP3eoRTKC9ls+
Ip1w61NYQmq23QIeOsiDoR/ctMsWfzRWcHo+JijgN8tnZC1K6IdIfWfNnBbD3C0X
Us+zHspLpaeRqxUkKkH1IcTG6KIkD9xPcc5qtxD+qsSWh+VpC30K3u3INcZqGX/f
FRmbydEBjXOVlLffDusu+R/GOWC7it0OIMPivhU6smq3llE65VfTwL2rj06/GdBo
g9uTBZWM2PpGKCuOhr508QLTphMnuZugRzq0zL5A8g8lIj9ahOj8n2iULa37NY1e
6zJC4Qz7znZmDJPJNKuHSMitx/4nf7UxjMEi23NxgysegP/IxowGvOozGZho1n3M
l69We5d0Or0NR8WqDNANdgqfp1Y2mzSwnp9UOflpf0/sDSVPDNWkP1GbLSmashYl
pJCrhEZuaal+Pn7pvsZ5Ty1cXzQTPF1AxX77cWmYm7zbZZc0B1flU6BSV4kDf/93
4i59PJyVILyGabLnhD1CkcsMc/W4OQkrBp8VsZcFl3124opQx9sAFizIery9OQAV
ExU/MhnvD+BrESR30TYDMI03Uz8xye2Nwb1OFddj6r35LUn0LYIQOa6/zvr6yiLC
ivRVUP4AdtrOkw8/jwHRnBWarnl5iST+VqlG6dmq+BQQb7Kk60sUYgIvcWH900ux
hIo2B7Wzps4YvsH1qN0YYDYEkkEK2yRwGVYq3X3ZkbANrBmOiJ6UrfUFWadCzjr8
xA5Bxdt1AV8H8WZUKGELhnsCWvwLaxx7oYbdfjiC1fCvaYCtGAMxu40Ur98aTnKX
nkhuBqEJFQWLS9rpCQ59hFO7vIyjTjqgjzt70e/C1i9UEleYBH9AbefZTwJlIvuD
6J5SQ/UKWSrbCqBX8zN+BD2j4P9UcPZhnd9La+BKaueA4R7XoyJSRCrVIJLlq7sq
t6Ish8OsiYIOZaOchWaw2P+UkUNbJDfZKb5iAbiYq42t4z7N9FK0mf21Ym7IrFZR
NP5YW6okBUMM6+T7E38+CwS6P988bQmf0OKune1GaQ7vfZY/AAn2IsRZ/eixH+Z3
LDOu9G1BBuvy2EUqozEn9qFUihnb6FaO0SFzWPF4DJeiEwMfgCk9SOf7UQc6XUoR
Ov0+RtehyQPgZopj1a1T3TiSiPt66D2KJK7duQLFzJ6vxFKPZuCf3CO25+QOS5oS
rEicfUkH+Zc46mSNzVC9n1wGNu6lhUdOCApX9Po4mY1cNYZOMwhPC2oMp7cdOO2f
ARn/0dSZ7qVt9f5POdFIIISUWEBgjRCJMlvmXV3HmovXTJ/gSCuliJt15SpruKyX
ELLz5JOUO3/ldtiWw4444FZLWpzhNFzGblfMe6aq+/tc9sFQ9KXWCLLHgurky3aD
Y9yHYAUeB+YsAsSz20+brDF/dmrorUB3gDdjNUcqJ44IfHW1pUKf/B8490QfKezT
tq2k+gthFu1tvizBAZ3UoUxBEUj5PZtdwiU5aXjhWGYsAPIujVEMTM5bWTCO0XD0
3NRvnQ1JdN4h3AnTloEAtBoCAtamn/Mcit2i/gGzfguPoaNnsXEsXFWCKMSnvVNA
R/cJLUT8NQcxppZam3pRBMVq1w1Hjz8OC5WQCzlIK7ixWZWzB6ApwFgof5DsH1dY
5bBpO1nh2BQda/6xd6m0e0Km+ZfUjJV3uzlJKSugYKFQ5AiKWFh4cjS9rAQ0RngO
kqIq00Y2zUyT41OD651/JOHbljxkZuojbwtw+NP0gRhrKBNk760TUsXO29gbdkBZ
EGNg7owX5kcg+SXo0AYlWj/UXwXugFgMOSo+8x4Bo/l4MpbhMJfQ2bYBXmcSJ35J
QfHQS4ELTeylZnfp+QUTorTibt8bzEG/sPBoDJsP/UIc5gcWGOVp3AJlPx4ASolm
MqaOIIY1se6/fsztUr8ceQZ8zQvzEIb0oMoNn2PLgnjrrJFr3UCgx9874qqv/Dl7
lPNpeDiRycsHU0z1/eyDMAOr4rYUM8SXIDJHjomXFdMvVhPvo7+kM3wkH57pkPAt
+A26ruhZRIhY+Y1avUC8uusfh6lPry6d8fnxPO1NtYLxPQeSAFG4/BdfMAYiboMG
GeSM6UwwBupzYaipyIA+TEljGKrj0dY6+FUmzgWCC1ECSKf6vpNXMc0owzu36tXn
uMgcSRpjjfz/dDWzmP1DnoCtef8SGZRtsXUA4GD/J7xiRfMFbEjJCVdDE2cphMom
7lzMJhP2fOnGBI/op5h6DH++8uSiGwt9LM8EiJWH5RA6xm6R7FcLMRhWEu2e10fi
JH+VglnnVmpgL79GtFoPQucoHDMY+wH5vjm8kjij2MXCt+faepIwJ52apKDIx6iE
NuS3vbyrtAHmZ8OYwaQ1B39D/zb5cwstoW3KzjHGudEjSTRY92q8MAZZAFzo4udd
OeQYY7eToTqfa0uGgCkUTgb1fKdyOCAD6GhSjoItY/O/ELgXbj6JwxaXLOwB12uB
IZxOTGpaW/nghHXQBiH5GAOa01IBBZcAbgIACX7IJQ1ZRssvmlaDWellaisS5Bca
RdExBBgQVBRmMw/mE28cMw1vUI6CMM2y9A94gZcuzRb9Uklb3zz6S/YKMl+nCsXg
3GY3oKbJCCdRf7u0HSJ7Jtd4jMDP1QrCtUk0AyC6dhJqHKA18t5jFCiRb2eeHJs9
kzdDDYxjP158x0YJui4ZKeVkfLTpkCDHGJugk4xd4mZZvr0JmGjif/0+pnlwNPyn
HmtA7woKiSq7Dy+1jktNmYsqf+m3iiTjf+J1YihmTPbO7y0DOxgOIlQ/ikzU29Tj
iJBJiLg4UnUVNO8/brKkEW+9Y6NjUvA4ntHMWKtPsvcqAdewZiCKWSQLl2dbr2GB
ri2dvI+zXgS4v4CV+gcC1i4RZV/K2hhjj5lZgMLzra1oWC9Y/+wGhmKiVXIEyLQ1
J3OzPBDd7Agmn31+SofE758nYtDyhAEDkvzyTbY0fdMyCLM9P4+Cc7JJ+5CHsk6d
D1uE4tROqc0yIAwUXT2MJE4YE7ivvAyddSAolDHepQRFnNd4jBIQ99e3f7/Etsf9
ZjXWu63qRGTw7PwYHu1znO4mWJswIzSGrytrkp2EZLet1I8IsYvmEcHvqJK7/vbF
v31Rd7vSyllxbMCc/O+wGLiOggZ3bU7Z1X+nr/1yWQXHk3Mo3Ynjv1iYTRePZS+5
0MckS21WpA32P7X9oG44iRB9ygxzYUD63xWfWv0QRNDTVBaM1RrHZW+tETuUwEJJ
Q/8qeigCf2d/J4LIoZ86z1dfAyd78J2ipeWOhxLHn+Y3KoZXNFBiwnp5YCxQhBvf
XqYr4BXupnnqdyq3T+YY/XS2TODO/8aCRZw0cv4jMH+S6abNc5os9kFI5VgcInYg
r+fqfdOSyyeXuH77bIQU7UiYo5GyyWtRdDZAVpOM9dwGZuYrL/zUjBdc+eUD7Cnv
tNJzErPc29Ueyzha9oTVU/PLo9fJYLVTwT8qEccP+lFoGH4/wGXU3KYjIBZSnGhS
espFRrRLrk/mUEMqg8Wn1so6QtrOhD47cAi/Y829NwZ4qpEvyi5BienK0HvpM9Jk
OzrXITBZlTg3FvvrKMsP7avlt0ArzcaIwNWj8P9cysMPNkNZyvTlIqy6fsaDCMC4
XWbos3bAUtxx+ndUIEHepUrRdU2U6M2XKpD5XUNrBD9lzLZVkNpfAbE/N+rZ2kIf
6PGBuAB/RHYtfdbtACOy3maJQmYPLRahMOzuWeZsDbN3fz/AckgUWFK6hCVdR6Ry
k1kYtDhxwRYIVGvIFzAJ7P1xQaQEJv6LBDgRavESrX3PWWNhA9ZyT5J8PPqOaDje
ECNn+BdoC7pXqoMxegjiljG11UHUaaVrUiU/bKrWfkQwkb0XoaqDF1r+OIln4U6O
dTZm22+b6IP7FJtaGjetTJRRuNW9/ru8yZxBMBkLNLk7/T9k5APkgX5IrASJD81d
ujvDJ6zJwwPBAv+jRi4wPTlNYkeygsCBvLgHkVKIa9e8zOwA0pWEPgY/AwoOTLap
Eujkp7keEpFlFl8iHqNf0xrZ6+EpWxH5eucaTM6GEZfFr9cRo6LdtOBwisHi6R2s
oWHlHMA4wxeVoCZG2IF30+I3yx5wBC74+H4zSQ7a7ETjkLLv1ymvQcncLGBWFhAf
a7z41xi1dGK0RUzQTW8seVr5tC16AYEwoN40aZ0VOzrbeoUVXuhnSUzju5hmP5SZ
rTNkaLePo5JMkjdrb1+I5aBif7ID5iijq+HNCr8pE7hOclaH4MPGpPS8xKnK/iq1
6k1BHhDcUaYFZUDAjqHO5cLctXR9sH3kRjpIZrh6v2b7SohX2sNHRGvelJ4y2z6z
CtRDm/osYYT6dSFvkTbsSPoclUR1tvVMBVMEd+pWmvOxfA3X+1Z1rTkKo2949Zm9
WoUaD+F1cBgtj0kitWWiuHgXltVXm7Jk3hWRBfIXGPYDAl8Kx72bxpS6x5AIZv3m
55BBlmVJXoBScBN+1OvTeJ98KdS4ar2fqY41tCxDkAICEJaDVH/B82QTk9M0VJPc
sm81DSDa7CbmxreZ2md77JNgi93N/e6ipIdEZqSxqWd0UXz6JY2hGs9Z7mhHsZri
IyXffgp3yWKT53fpI+0pRfe9Wpnl2y/nxGzFy9FS7++Yidy61EXeMA8qYH8nWw2x
MQ91HR6YKgH6roO7QiHRqcD1g7OxHVf48eQUnNo6muTSBWD3ZElv/RSTXo9XPeRB
d6joPLxRhMCJgLz5MfHpIa3R6YHQCVxmEwleCRNpHXt9EmQIHgOuH+X2jOJYM6Vj
gd5AzEpZfKoxv8E6srjmlPB7O7d8UfDWD3PYa4KcBjFKPCAosMkoFFZLOk6Gj6Hr
voqziwZZ41bE8Cx8RVZUzAM5fQcGO9BncBRlEAWlZ5sFdNSmw84lLIbieBBP/Ypa
gxBqkxVycwYgr1OL1PoS3PRXk2PXybH5BQ/l22cN+egiiYrthff2eqojTmAmq24n
YRBD9XrOZLaQTMpQCG2l5teoy5/AwzJpmOsFt5Fgx1MVdoh2io4kCscnbhgThOqn
zSFhPfIH/AJwO9TfEIaNkryBvdai/RVHkkK9LgrXrE1nPVTC6X4WvA/lb32qYtYq
eH5a4Z03Q8gQ82Qw+2Aij+4FqW1fS8ASwq2KZyL3zg0AWFCdh8T5+gMJ8mcFg7Ia
iSe5rwDUR+8IH8cvKL0wMbk6B1uOy4vh8MZt268TcVGZR6xrTuGd0yIvmkjZ2Dxe
Dcum/032C49LGzUOWK3QCs9l11p9VfYK7pTCMB7k4xEKLbNfdrJ3qtW9Kigf+e2N
I1LL91H6veLlRs0na/cW2oKEHG35ps7F13F2VdCsq6cJgHwUMxqirb5CQJgbLeOA
elXmxod/mZl7HQQJYAiiK0IMD4SVmK4YUqvLMURRmikwGEzd1s0GAwLN6PYZY3eY
srriHeMehP9DsncX+3iyxjQRyki5axsDYMs0y1hxLA4MV+jm9N5FqKkJse2IAoZY
JqK08H8sUdD3CjqpUcCfTqpnvMgaHA3UaXZo/LkFkCDsmxrYRW3365mgJ/AMpVn6
w630qPeh+ZVclPMO4OmGd+Vw9/DLGlCAkVp1XMWAG0OGGmgROxFbhr0KGRqPzN/x
7ELvhyWqjcaS3YOk+tSFIMCwFEW4mgM9whM8qvkdbpFA2rraRHR/JPO3CAWwCMus
dR3v7KR7tOkm6Jca0LOpn3PMw+YMQQnPasOOGX80kJybYKBGExTu3B+pqUmzYF9T
S1EWAWd6iz7C+zBQ0E5YIB8vnsO3MltWuinviGAq8zbBuU35jnBgoZ/Tn34uHcYw
W67ntHRmROyXqifrhfF7JOCkpksPYspyfvQIVLAt910PaWYCgKAWfub9e9hkSpW6
HHRwm86hyDye1jJB0WjXJrDlZBshVouikkO842HVTK4dQkaibU+9J0Stf70HJEfq
VfYK3y1eJwkRUqkY9KcU/tbEVOQgVFjYGm/x+2W3NTXaRUqEnyM7W0ZuEGq3TjFU
NYKxPHv86qjz2U9yXRiFi8VIgtB8lHqrqeeULVFUVlKokgmfN8CYwZMRHqNYMxvJ
9BAM0PH5PSEQsI0YfGuCQyDOk9Os5j/B6YvimSDNrefHoB/MZlYAHaj3JCUFcmkN
yTOt5/BoV30uYN65Gjj1RbZI+1uhwnNWzaxg91wqGir6E4RTmuKRGY8E49LFjKEw
JVrfN3GRI6vn8LHsMFqqR1ONNygI3c8aiPn2FhYslA7YH5KaSi9P6csodw86CMUa
lX1G2MWC8efGy+1Ax1GxSWiSE1UhCSS0Zj1gVBKLxpi7dZNnzKTKIKd1fF3Owxi2
xKh7FsujZV0KQ9KGOtKi5Wc0sI52NTGG2sci9QZkTh2aSdtvDuZBn9z29UGlj3EZ
87NVFgfkmtmkZWBPyM4RdkVhzaayn9QAC9//dkofQWz/iWJX0bSOr8V/wSbtHvYa
Py9rwelJKTH+9G6oC9eZ6cWP4w7VtIsteFYzngzg3jXl1LSmtJgnKyNb/a3TQBFK
lQYn4Icl4HzW2QkAppP2zUi8ipM1gIgyrfgmPbT4lCjSGJOIr+b4dEigfhENjlvb
P1MfRr3V23V3VmPUf3VYub0cpLtldx8+CAJ7tBkRms+VHNFvCr18ogcHrIL1VOx0
S3QkkoSf3aR5jP1GXG48APE0ELHJwjgdAcRZbWnOd5MfaD37V65+6aQrBk0HWHYg
FRLUk19CwVLt8CJWaYq0vTQ5bsi8zqMNDISauq2bUofINt4TkDbMDSa0ZIlsGAVQ
uMaNk7d/hwJ6sV2XMorRSXoARb1xJQG14Zgpx3iRpu6bt5/PVeVJ/9t1VhCK+L99
iKTaFCm4Uh0nN2c1G5e0p+phaKO47FZ0CQDYlYXn+bja90TOEXH98SLeHDvZxt8Y
TRarYocEWUIzj8HryqPlNbla9QHG1/xf5LO4e97HnKc/DdcAR9PDnzuxX4F66c3j
2346cZPribJFCOatdAb3NIfIv2UQmJlqTqoPhU52U8UBn9r6e6MZK9BL/Y7nj966
khz8n4mHyqBqesfNtZAVqOH0Y8HYh2SV3trXjdbVgHH6XTv9asy3iiVkamS2cho+
Gy6GJ1QF5WM0LOKLBNQO1iDGV6DHUCUT6T0orFq5Xb5keU8OuccoEtyIBCJyuuUe
Qn3NxDdOZ7MOUMdDmsM8W6ajDLIMaAmx2abGH0jH5nrrGDwuUwgknkYtwIuAg/uL
E9fE2KL2XrURCBY8ugirgwnNJZaIwMmb3LuhdTVhkktLUSXShx1e80BWUfcIEbAR
UdDGzYJIfDyu8feIyaT1XEW/gpuXDUpUtG0E30rKwh6xZ3EegEmdrxPzYhbv22PC
HPs1NZ8aoLNv+7/eoFmUPMpxS2JpFs1nnBqhAUXVCikA+nrNP5UbzZj9pp+Ox/R2
HY7sdPE8GjzDNYXcHAUpB/tJwNR1AYFfkU/hCBqYDPH8bKo2xc7i5vG0FrIvhDeT
TGtUBhh69eEqxMBB40cVPp9WBACg3yHLaJwKm1P1JrKFIYNttLPewqTAgzX2bnoO
wj2FLVrvU3Q5Xp7LXeZ/jjZZZQkwwmnfTCP+gTIDL8OyEIjr7F2+ETSBUjQ0arsf
k+0a2XwNGEOVkOXU25Kf54iVpJRkvzD/vzUeAsYZzq9fic0RpmztkRn0HZzNL4CF
5YgAVqxVr1MMjkV24VGVHBQxliFAJd9tuoiD0oYyAZOmpkw3d2Px219ULz64BD3J
a4FTn+Mt/PzgZo91T9wMV8ogveeDVmy8kiYKHkgrbT8zkTVMfzI5LfqxorpdOpeH
pMn3XMYTNCCbVI5Dh/EcaoNTCIF5JmPg0A29huWlgdV0gLsnWP4z0gm1nqsVID+r
VfQDZU5cX7sSFQelXUUx/wYykW4k3nSrHiZ3hQeN1WkgdRBPocZ+YjcLBQ+paDHG
IUrZu5H28PqjbYAOgWF44JaCTuprH1ye1MtORcgOkRjTxUaQzGB0M+7AY2z+b+ch
XUhwb6XiqxLE3ZPTi7IQ9ugVvE68OC7gs3k3Sw9qvEFczhxxQVGmeNCvqYO5KRwt
921ZMjlzkqUi1ygl1lgGnxmXp2+i2kqHYTqY6iSQs1pOPdCMJZgXF4z6g93j/Jiq
ILQIlvI4g8mFrny4+VpkI8+ovEAQxG7XuBjWFcfbvMngQlrU8EDqj0ljIZSVzCD5
oBpSsD1sCiVRYE8TGh+3ncTDWXIhDOnV2qPdqa+G3ZXXExxqR4Ai6k8/3nn3/6oi
OK1RUioxRP8zV/q6wQvvT3Rqkdo0ZUtXZD1H2XJKS03hNFeZjUYEPM3VU4B656cT
XhG+0ypL9m13+eCkJAbh9eT5vmG74PMOcM6gMhbSzJdk/8Jb6hf5ybC/IWuUL6uK
km4zH9WjYBhRRrgxRCGney4CcK/Q52fTvbWYj4x+TqbpLxfgt9vN9dWAedQJCv65
YRIXYydG2AQurs62ekWC19Drm9ubO6RGWH7J8hEI1utZF3sGtmtT8DzmXJNDGbpB
SF8jm/uWLFZLCvFe2uANAG/js1fHNvKM5Sl/Z7N1Y0LBsP2GSylztR2xj5/wpAcz
Cbi4HRa+8a53p4Mt9osBTB83aK3/ihoguMQtpnOJ4kB9wj4zHgkEDBy2p8GXVh47
DPfQAMBRHRvlteYFrdVYq7F4g05UotU232R7ssGAXDgbNCfngvErDatvFGY/88JN
bLoek+NfgjsIDZ7OKGn09XOxNQAzKbBzsZnEZh2iL5bba1Z5BXNLkZW+lts4tDEx
OCNqQTrdIpIm5/uWatM3Aaq6b0gzQQpBOyoX/GHEDpXlglm4t6TkJU+l5L0hQh5U
seulMmpjbbG8/kswBD8equHAOFRCRs+ntFLWaxpxlqTJ5rUS2bTlv2eLpKgjDK1D
UT8QIC+zJ1nNTMX6m9s2uzEvc3iQoZuL7UAOLqzqcvq4FyLPfqTvfySayoXgiA9O
zQ23aPp+BKtng7pil1KymH5RrZvJJYacw/QDQBUwkVTNGL455L5KTVIQvDV7t2GR
NZBUyd8AxW+ZUYnrmoDRn63KwhAHXNY/nlIWJoSar2pcP/BQ/HuHAwOFDOJjt1ul
mJ51Skm4XVzJ9ZOxXMDfwBMNiyDcLmn+vAb7qhqmta8KZcLQQsFNMW4e6yon+EBR
d5R2qiu35MMN0gfzkZ6yefFNWZ58JXNzIxr0h5VA/KAjC24KKC5qyGvuVC20oxva
/NXTTzCkE0Tzd4Q4+e8GL3tHjR0n4UiT0eTI1VoM5KJi66PbUgRfYpUnb/m4NToi
e4ywhTuNoHb6o+Ka8TCR4G1ZzY1jieRzBl4Pg5/xcYG/EpyW0d4C8IYkgvthp8rQ
Y25ZxfrwcoQulOZBgpJ9Jo5w6Yx5ouqlvT+CUFND4it4ICdtqW54fCBxGaOrgi73
cW7rbpROt7wPP5d7zgdv/Lt32B/+I9ZfWFnUIn3zDjmP2kGafun/O6KiAfpp6CwN
9ObSRLJrZ45ZQBnKpGzYknRjOkWpR2cS3QNdYSSu1lhDTrZaLaP0tSFbGpV+TRZD
HyHYO5STM1X44Kp+vsx45qd7ktbjLY1Ne4KLLIdKJQ+gG9R/fPa0Ws2aS/hI/P7P
pPdSH7ONbYFFNnXj9R11B/Nj6jErGU8wC4Mgmuc3cSXp4bMHW7a/Y+kZslKmBjeW
hhoOzsTHFPyKY/W1Sc7qYjb/dZZ/gYE3/g8kPIpdLZDYtQN834Ra12SDFRoE+U29
0Nlwa0rQTSDY8ELpi+snyU3S2eEaD67N+w76aMIpP4CoJy2lT+over8ZR2I/4sby
zq0yGS7kLIDKHCckm8nb2i7rH/u3hkWHrgKqDUZg71/lurnOV1C0Srlfi1n3B8aU
jR6OPGYTq88jkPL4wJukQhG80NgkuKckIexJTgXqol6MHyrrQAY+IwVuCyb7DDyu
hWwhEO0ZVHn+sMCKCYKoUvcYIaZjteSmh3yqqwT4yLq/IxzF8Cf5FtL9jXCxk66n
PsvRpOVX6Q7m+KDLrlQiBTuVUq+PRCKgko71BlPfShF3XyU1strUrdbJHmN3pNex
hFrXdbmc6Tw26YFrIZWUvnsm2DSLXdQA0v07qj1RdgEaFqPlJHkUTAwoA9DJRdCk
9uBvzBpdbPjK6LQQIHpk/iB4oxBwF+akQlIx32Lfk4A4hMNRkRtU/223AN/rjaKH
WMNCJKulk77jEeSLNhGGwr7VPNQa8l8echW12gMhNloc9fUOgA34XjBksblAaiMP
eGw05Y+C4jUyQp2kfa7Y+H9pSvKO6JL2e5880mG0AOIxkApw+oeAU5mSFVcNiG+D
7wPS+dPmKifRHeMGbMA9tswabDJaSyMKzMUMrbCwWjtKmGtDax1ruCO6N6YGZVG8
zBh2iu5ozub09FweMoGE54f6kInPBvJdSjVNgRPpBS5h0xpXXYZmrm3x5yHvfcHm
29XGmVaEnvquFLnqjuFZE1Uiak9zJnak3xWirqKmAA9WpITVjc3knK7vXHH6jqn6
8A3khI/NoBB2Fv+y+f5fmpLUM6kVYthpICJMA8FcuCK5X21izb+TJ+rZP7jPM7Z6
QnLSNPruhc4sjon2+z+JwEZuLaHVqKo3amXHtizh60eTqf4H9SXitLy/tAsgyobY
VF3yWLwDBDJWKhXui3XGwtnMxbH/mXEqsBjLxb9KUEThZ31OgmuswmylI9bIDiLi
e7rSjxZclwEzTqbaF4tloiLa5CmY/JHfGXbs1acfCAedCMFVS5T7Qe49n3Z1zE+N
f0Xm5ABffY6UMQfgqsEJJ9mB8qXVUI+5+DNnrG8aF3rkoDCrOtmlEY7bLfLWrnLp
oRd0DlnNMIslzF3z0izvIYoXKb7ggzSx7zPUf4b2coIhwnAp4tz0Hg2/7ueyKZCM
Ft1y8HcMlseS+VPkkUjFTYJwNDEaAKYe786Gs5nED2+ESAuvFK6zCyFYskXGscRO
ptLN0SFAcSghtyntFSMlrctM2McXewTkffhM18JiXjSNDLHsLLL65NK1+3SiYEVl
+949bEOYvLftDGbL27H0nWat7ticxsFMukBaRMKosqCOiis2U5ua+5383jp5OOGj
lV0ggarQe4+ZR56VTKX57yOp1hKQk3di2V1imjwcGOtOmwGCo3oFLpnRskuncZ5/
tHjLLhiPWa7/LlmjujvNtAKoMgDySjyU/zZJLQBKkQDhIssbj6U4F2snQrxwOPQb
PdDj2189XqpVccrAwhMB37xizKVEvyZoJXR5a9nei83vc8SdyXYc6DWQhKoA8jzX
AeqerNeDRIVIQmgpuUxEZyfX9wHziuHhCQFQywkomne2sQRIPCVlbTBNhWpciznh
FKz3rQGqOGCkZFW6Fruo03oC30CSMVsAnssQV6Wcf1vO5M7M14nKsWj9kTsqRlui
HbENDWvAGE42t1eOnRAPeweIwG22r8L5M+HuxQVSIXdZrsJkBLYcuWYrpa5SeY9C
Dni4s6OwdKXFE/n2XuG7PgTT87kgGsJv4296i1qA0IvpRMbRkbWMf108bIVprozk
DusNjal4nP6eY0tr/sKYHhAIJfd+uZiEm0ZOfWJjrjvlG2r6MmCEWwdIUhR5Ozyy
7DqRigUCShhfeau5wdaGnqIY/+4+iPuH1ZOxBt3nYaFcwcxSx+VrMFIXwpeRzKJ9
HW+sy8F6CN5hw75gP8sMYpg65j2Hleq4pcFOLt6ogsx9uFqM5ehJdP5pK1PrZjd3
dND13HYDK7vKKgfe1tTxej5g4E78s6lwZw4v1to0/VQPqXqz5Sk9eUdAS1elU4zv
b/hURquZJo47eoq2L6q4oyHqUvFBMRa7DYWWrkpZM9Mc7JsiHOraAquzwE9Xhy0v
tmQCACdTEDMqb3smVaGUbzlOgzLN9TnO4oILQzdTSolPHBFTIIM5GuYWQf5l3Pbo
ivaiAzUjHrkbC0m//ujQVReAuPUDyzvfat51OoBbsJa8llOOlCUhOgn9dSfGnSm+
ZfqTJ9wfBvkbM7tbrSyJe1DGJM3yzqpxsuECVljHOByb/GbRifenRLG9SssfiM/O
B3Hz9/WQwntDXh61yMpbQFjUHVvgJBVYKrpQtzLlNRB/aIknCZkRG2i4z/gx2XzL
GJyUONzVcNWYvXj1J/B5OeC0AM9cDWpsnQyft66BV742rFmXHjhOBNWZrUCHpIz9
/u+XE1fkvkHklodbETNkOCfXL3uAps9gxs98DjaLUxJ6MgR+KjE4yhepqtqi1xos
Nm27jPvpUjDJ4B6JP9ojd/ZAFWpfIswVIAkgOCkiDsSfNnkUblpl7G//neRwBSJk
yWq1MlwMzyTpSW/DIT+9LZQPF1q2doJmJhoiaxgdZ0vRJVCpCoQKceJfn+R/humf
Hk1NiAHXmLQfu1B3ycmYQRCp+ysT7g3mMWlCDTF+8I4jVNHpHyeyjl+bjcg+sZzr
6xN2cYMIDVuYZ5WXLUz/rpaaFdxXQkBNn0syf7hBRmQLZbiWuWHxNmFYJBr5ZhBE
vj/QyB2j46U/JngAa+ivVVgp7jFHEMBc0t1G5GdINZRRD3ct9NxRXk11mJr7ZmyN
rDgLPaV2WXU2Vy8VRk+fQKWKgJhbqBpu9ZPfOkKrHwpNyA1hurbSR1E8uy35MtuW
6CSvg01dwfEgmWvXbx3j05CM174qf+/NGSO/7XZsGgbDG/ADd+h0WMBB+Hz9B3d4
LWGfOisLRPhtHemsniu1fa7zu8Netps/+e6kvBrHNqqvpsSYU7KUzDJmIvI2AGOy
mBH6XJ4E+PWmQvuEzXAjargs0lLPJUqlWsq3l6Pss1FRCFjQc6zHQaPoUCB0Jzb8
IcYZe4RI9Q1h2Tq5GuyvyPLI1ct6sVEgdqsgj6rLvqIlavbmOGysmj+SePlzjMhf
b5mLwsAJ10kaxrfcAXe8yE4sqTG1eWUWvdKCkaBmup9v1G/MSgST90VPc02HZwhA
Mb14DrHDxCO4G/Znzk9joycJ4BPxRmg974NiJBBnxczGvqu4sQjk8uEJLHKVT4Z4
0+3X2+faijU0jSAJaikw+udr4KvDXMOyXGz7kQbAy7nWuw52i9Bd0kUMoBKa0S2A
xHl/weWpGRk+6VP3bD3LDk8PH1pbqCMfr3QOW/Bd1S9HVmxeaoPIjpgWVG2AkqSh
93Ha9eJbz9YHCQnmFCulfn5OCBvtjK6psHxZnnZ+PFUYaYb1VBAovZVwylZFmy+D
f4bmIJ4InqnLe2UiyWhWnkjacIMKQvPmUVCFNQuL3tc5WHasDaWOOuQIhq1JBS7u
bUaLTQOGj8BVB47fpGAqMXLBykVOO5cXTRMMR/D8BNHvzNzXNMMJ++7ALkgk/fDE
t8OOt2X5B8yWfuhKQkgaIA4MpJUtLcOMGW7BsuqHTQIdN6HDLxmiDmXca1rnh4BY
njwQ/VBkbdOPUevuFNCRTaHvEh2eqaIY+DfuYddFRio9pGA0fS+3v5BzX4rOPMGB
XBiZNG9bjDQ4es2enAnZgeWzAYLxLWpn27WwzTvhA9nGivEm7n7EirNKdgNH+5K+
uMs1fsrvDAi5+eXUcI3M9SfCcqzSTfRgdDFkQOhpKnAFPXNzJACy7ZuSg1ZJJZCe
aZdwUV6fzhuq6GlNI+c1UbcRi5MxD97yOuonS1Bybu8hqb12/nupCMUnqZi3kPRD
8qBgtZgQEOaGLQxkz3pc3RuQcXh8J7b+rOMZIyp/pMaYAtCrgGrnlGMi6fnwZ9Sr
N9EEW/Dux1Cnh2a8O+3Z3J2Nkc89L5S3MZI260Iwa+2OVHqE8mPIEIC7ovpF7go4
U3TgNyHMus/F23Au4Qo3PGdzEeMc0RlYFhm7NQk5ukNdXMTeTJC/qnOr0jLtLvyk
cHBhp9Xswqp0CHnEDmUc7Dxyhzxbln3ZXkoVyk3GxWarnhgvBg3NNNZj6Ot1l58V
fNvHXjEsgAZikY7aqwgy6abX/prgRawvU1xMotRK/W5I1443IsmhDhkReOjmrILu
x55cpQ8VjIfTyFsyU+RLqGZy6skfeR3ZhTzSDPuEXrbKlzQI6MvE0/w5dtfWhUmX
lxgHByyEq0U01erF6i/S85lpavkye/2RbvHBNfWN6vXCcszJtiFfv3Pk0ZaJtmsP
9YT+fZoyAtvIRygvyuNdv5WJaC+EwR+ExnTm3lBc6zuj5fCdlBSPULfJ8SSr6WGG
bLplEt2jQUSgBSaklprLHINyn7u/x6+Hxdhd8wuVwzPQrEpk0d4nIOkxVg61sB1k
XHcw9Q22dRN5HZ4E8ZAJgQaHN/UVZKCY8BkbeDF/jzmmeE7VLdoFcUyBMcH7Ejx9
9p6jfWpRWE9lrL2QfMpxMfg6ZjiABt4ws1u9vx8f1tmweptHupRP1UVfvBykZJz2
ACLrwqn6LQN2Rcs5DnFhMVfNNVCm0lS9zL/nKUzqameCYjDOpJaa6K7wd6Q9OCso
ie4dAZlvFJVZuwQ7jvwYSKYeWiBy51D5vibfnOxHHuF3c6p9cGfWRVfagjf9fLVZ
Sm9E4i0H7eOxm/VVsvzg8/FGTpUsdOGvGwcgOT5kH8EE1f4qrY0lKP8Q5JX1RyJl
uo6j5F9E6vsXo9cYVbFdITnRBgk+sVaHv9jdsPeHgSu4ybWkVO/yPYgxI7NiM53h
brEqRI/2Vao2SdbPH5fhmJc3h9qix1quCTOIdd07zDERCOu7483JJGL74chSBC7w
BANhPBvO9WyDlb0e2Wsz4jn2Cfl7RatnItJ5EsNXh/PVBeviw3g/o8EgrdHHvxaI
wqfIG/5VOpqBlPOiGmcPtw9DDyU/lM4WFyRe8rGRO+nc/jg4RNCohRhXbRf2bVMx
oVZFdoAjm4XpoxMrYBpVyziKp09zEfyMIiaxqGU3fC5x/opVKe1vCiJWc1IxWQ1X
ON32OycjlUz/FCoEzLgB+BLDnKZEaUAhsve1Q5ZuhdI2SMvsyvJxq0Cto15yMAVW
v3xi/Fsr0hQds86f6KwY6fU4BOAq37kmdpvYkhULQ5nE/a4pCULvPLVky9RD2cu/
1pGTkIpqbyW2aIuTrhpNis71HDUNki2Dd4i6NfvQ7SYoW1i5D2f8h6QGsgUtDhrs
jMuVcwBmcDVtYg34JZnLnZQukhSbSj5z+FsxfY8R1YPxJPHMiQZXZ6g2b6rg5D+8
h5tYi8qLTeC33zx5vBZRsrrOFEu+DbR4cblnVX1dPQLNEcdfixj4HdyM1fHybmPr
fsCbV5QlAhiD7MmFbm2I1S959EDuGGQ9QIixWQmqUsdPrhsuTi/GZvkBUuir+wPW
BczNeQ8t5t48XL8feI9j6GMej6jwcrGQqp7D6Dl3iwy7ZIML6o3+2PfOmBJJ5pqr
BiSF4aj9nLOSdIpnFnmxhImS15FQSkUBpRO1LoXniraBSsAWTnShp6DLT6Xm0UYy
0MScnxGwldIuNw4ynpHHsbH1ePLb4fwCH4YSUQbA8zzAM6wJxvZIhub/NyjAaU2T
yTPxO+YPd0NFS7dCugK/t/MG7dEVucqOGGcIxOvq8HQiiJxHKWlx023RShY0Vrpt
/Jos3fJ8/yIutm5o+cvgfbQTSzdpaJk3LKr+403ZIxcVbx42wmKagL096rHl7EMf
TdQ7lYJ7DKYTVxnixuBs8KXm5mZlmn0KdbXHRIxm5ZXN+ql71grsWOEV/S8j70Un
zE2uPvmMVvjr89ASEhkeait//nY2jqctllFpPRIYyjN5d+bh+3ZveeopCjD5gxjU
cfhJpvpKxa5MAWs6c/f6Q0DAL0HW0zzpQMlou8O90Zvx4DpDlvULIDEcRN64+Wi4
sLhUU2jFF7lCRpGzBNjAU5TLRTFG0ZHY7WdCVHpBBYPuXDlgqMIALWRe7FLdn3dv
0aqzgeWUh8XLHJDHP6khRaNgKXXwC03EG1ePigPCWq+y+7elSXv7F2bKNS7KI41h
IcA8crWPyRhOY8gCF52p7NF0Qpi77LNdGOzU2yAWeihHQ0eu64VdGxLBUkn+r3GT
Y0Ki83w+qJDOjYuEsiBdohFl96lx/BeQj064nCzYNBhh9IX6YoTc0E2tX+Q0T1Ds
I7Ui+IRMYFdZdv329XDZKoj6RVWahaLB+w0RS064kGxqzTeOkNDGxIXj3TYqs1qQ
6bkDoAOA/u6OzEl5yrapwzR3FZYyPj5QLFdqfkntCj7tPfe0t+HICcDmQH8F+bta
3HGBn3dzLMpQ2gRC0sJ9/cpa5LBAnaH0YftYZHzxEk9WKX2SqSUqCBkl3nso55IL
zeWRmIxdJTeVtXB/9aBjMFj9lLnXw+FSPWKi6YSfSuQJGwo4iEkpZ0HLj8iDARmR
mfTf/ycYXi6yyxC+xWz2azzKL00f/bwu/c+QX7plTT4gPJcM/5k1RNB7gFMxHt0X
GabgEGjmFEt84QOHflblyJtYW+H4Y5g2JZ+Ae+7ODJb70vgIUxSQIBOxongFuzeH
1LFvWpzxW5RuuZhax1h1iY1D8//8nXRvi1+KnAEckmGQ55QOc/9AhZyAB31MaNxn
P3+RbWb8zam0Uv0Yyb6UUIY+RUegSHp6CDbCCQhRMG9TsO/6czkFN4PcG4yJV8+l
s0q4i8nXlH6Cqfaudsz38tmGHW4xbc6s4EsAxkc40xqrsjKo8tMprAc/NJ3jHULT
xayawJQzABJMfVx6HKaYvIE8d3trbrtmo1w2KmurxjvW/rRKiNLtBY8qMgHezrpk
AQIA/pgLvL3JANqPVpQHcnw46T24nBfZSJergyBAPdOQ5gtul2+gcCO/9W1OVams
4S1A18U2J++jG8U+YMzEH5vfPE/nGBtrJls9yhOVeV7MgyKZ9LmcnKd4JCe1U5pP
KVdaMXHA89GYISfXztJZaRq2sQUjwMmgXrnCppj3sFnWWsNUu4Ge3pFRI6mq0Z9R
f74Geh3v/+pnml6X9RGbu5fdvogr1W2OBXS0rDIKLsdD1+wfz01ddeOoaVMCfGNI
3Nf+aEC31ZwsZ7l5sHH5WgG3Azt8Ujo2pkLIDyHvUpVBrkerfPFFQ+15ioAgF8Jy
b+hCnKgGgxxxA9I1pxo53ghlFxyZDhKYFyUEA/MIHleyF/GGWHy2a9ArzMb8Zw56
BZkYQqRwAP/gMemKDia4XLTUqJUAQnFZNuGI6x8mk223VEzj0QLi4ZPqZTSBtSai
LlXUVs3kILit2uGwggABJI/ycpOehujr3hPHgrDD54iaXQYMhTkEqnNKz2GWnTT2
5QCzmI+d7UsrYlh0/v67MJRkemqQUqYUUFUUuyINRrUavtyTEyBnPOLjAlAmTWbf
69ZOR7kHiMd+nu+yNf9F3NyPX9AdZ/pmyHQRCHU+n6T9f1H4wOBGRzjTr3V1+l2n
q3kAf8QF0sWMK7opsqo2W1exwXtxy2ejt2+1Oq5PQ9oYovJ+uARE2wRtRXuAEZFz
xqW9BwbwTQak7/gPT8HQ7V7b1vW1gLMIc7JvtloS8+fzQQsohs2uKgrmNlynQJ2T
Jl5434/TYUUQIWV0WlpE29xstq6HnJTHkJ/+2Q9dRrRV+n4bpV/odkNyTT3u/9BC
Mw9/vNaauUnukjo4RNV1gWy/gatKKL+JouiL7G6FsO8Oplkpp41tqwpYxyrMRK7M
ENeXaA43DE6kjGZmgaSobb3WTQLWFKEdoVas116YuYj0RZmkKSiinbhbpMG+l8GM
WK6oe8XrkmPaByJ9Hnmhd780nBds6RP8cr51uKwvyqlATOjhLSbelEqrW3vDV3rV
UToP+dEQ47UMXM/Sm1MF5tKblhMfunG/MMYPJfbGze4OCuHI259lcesSxizmX1pN
NfOmzoWzdiIhMucs7ux5cinocmbfPNAwdTvrO6jdy+x6RfmcH8vKivoI0eeXrmGM
uL5Rchvn6VcEjNEc1fq1wGVq6jFAHxpC6onoES3HXIG1lh0LfOuEnAFCk3FudMXh
XWQfdMpSMp0R+I6KqofnRnWBZEUDg7jNcfthokUKdf1XaD5OhtL+X7jVUufYvw/Y
DywXhbMEhrID1VACHEtQfLfXZCox8g10AW3DhCZxhfXNXSAvENGlELC36XwRliPL
Kv1aIdzL7cJQ99+YUHztwHzwAd1iosNHxA/IT6UknlXdr8xylSR1t9m3oyG+9u8Y
fAx/o+YZOnxpVk47amoj5UjSspa471Mq2TL5zMtyVycHTJCSmLkqKVEZJcF1wYBY
KOHNhZrTIicJZncK+3CGBKc2a5eb4bgj/zlh2AWnpuLnUjB+hBvkJOoUY2gEq/h7
CxB+KlPsj5unwS/PDp4ewcz2uBNmf3WmRD11vOJTqSs2rXCNaGydlsop+KTaRPS6
U4RXmU2SAmLeV8I0d9Rz4omuIazPo3EvCiN5gE2gfUFvM96gSj1+tJDWc1tcrdmy
K0UbMeMlhHTRUmakwkKMZ+7+p2o4BSCkYEd6Zwwt6Ag1gfLP4DoUjboUQaB1uiu0
2Y7HpuwXInfZnf0ObaeAFP6XZaR83l2ZZo8LAnjl2I9639X8ail9XBs4E5p8vCSG
Tju5Y7wrE/4xVxBWjlpkqZ9f+B/AFSxwf7hceQR6DEZUZkiNtBk9zT4BOlRrQgvt
hGKB0mNObAcTv9bx43IWHCjvzL9sCxBlbkJl588fKRg0+cNAQBMJdFLjBNmcMl3N
Y8ODGGBb5xthqShYWYo44hGbdcmEpoOwdR3GEv0PSu5TqTjz/nM2wTPqH90mMJyA
u4874UjdLgo3vc48snpqKGtVPSzTDKUDYZTPcb50+PU0atCrSWnH2UFvvXW8hlXH
pNnGYBlPhvpWEUvbzuPi/ZnIzvcPc+xr0buJ194FETIZaIovQHHBIEQiA2ecJfY3
MxN+dWMd1gwjvmtFEjFgdKhkVUYPmeAiqnA9Ue+pMNWnGkPa6lgrjTxFz/0MEUoH
tzfKoHnAlKyWbywejYZHUZWcZH+O8UG/k+RYEP7omVu1jZ6koU5mHTkzttANeP2c
m7SpANwwSqJNkrOBlsD/6dKMIaYC40e31OArTmF2mbs3QktwSs/m5PseBiT8HYGh
iMfu8aFune5dB16qCq/IiMLuKNYexXqGeMW4W28EuL3+QTIqLhg3WWC0bWAkbod2
O/2p91dZUjBi4TlE/E5n7DqpdwGzp+sveN8F0oVetdJdYPEBvdDASunLeSNhWtYt
M19BA7kHeYBbCSbFQPJCz9Mj+/KSLoed4KkFzUOVty88tViqPMG7hCooCWcg5BKo
XB/ABohjPSapKeKIebp/EeyjMtgaldtVjT7gR27Llm+261EuG2A5WEmMbhlbfNHf
uMwxaVI4Xiy4Ah7yTB3Q7vxSfMoQ+VEMqcuLGnf5EhGUPtBMcSh5on6Zht4BL4bC
c1cESN8gACSZP6WDMcNncKvL+Ypw5JDf/RlDV1AyFMJ6uX8iuYo6WIF1T3DhI4qv
2Jfm5P+Xc8Q/FoaQtLXZBa6QjtCWDElPk7TMAtjeHBpTdt0mvcOyQcOqcU9HhhbO
whHIYxsnq0+2KkMtWBlbP+zlaByEyHOJIREg+GvoBSCIvd5/4JvpHTrXKgwDoRh1
G10UfnZWlQNXjt+M7kjC112WteGbkqWPEmMVsFJ56iz+WmyNSn2teHYY9cJRN4Dg
hVmc3UFAMgEwZ2/1lgkyn0d860MVcaausveOvFuxDaTBuHt5N+ULzKIMrN80tBjS
nr1aIdCy4weULOQCvrUaFv4PiuEom4/Jd8C4gVBngyB0q4cs5R+eSlWVInJn7mIh
EHzEkE5rpRqmwjJUG6BBatc7RNn2WXfFlMxaAuaeU2I4U4mF4f8pDpbu1Th/GPER
Xv9M/NUnVEghYuYoHJHRd62BOX1YEPCWjmAVhqpBp5ns2BUih54Ow52Flru+RNnA
jyLm067/LMhrS3tVBVdoWCUgJthWz1U9JZmSBrplmXB49LIBmnvV9OwVozRX3ozG
Q6FagJPkJKUyomAX9q0iFZ6UwgQ9O8FS1Lo3pn69oZgrob5fmX8WTsUgbM3pXR24
TFM828QJIy7r43sXTq8LDUSgtRmXeR1PTjxrEOGyGQVaIM/2GEbu7QPtxlawjARp
AlLTbrzQhX0MSLUkTvwqbThyx9pHTQVFXSlhgb2g9hmufbTDbgnElw580GQhWtm0
AaxLOQsgWW9XgDHL02iqv1HWa6X+p0GVbRLIYSwHQ0qcgo+83ij4vAgv/fSOmHs0
ox8sYxYwMP0lPgSecMzqtc1RPE6q1g+9FsbG7bs895xjk6oF5fZznFEQ1d2ZgJJs
cURI473rjnacUtLFBeynm7tGGV06SRJmQ2rn63QdpWvJpop8ff/eHziHQYMHUtXG
p0Qhe7gR2KOhh5m3lozDP39bJoVWNA0U2Uqszt8Nc+nXpzNhKThAYsFMHADRgsqG
JvWnRgQpIJk+4LIQWqiqPc4E3XcTHBiZo08BEJkLVouSp8dVLia/GqqtNuMHVCWx
Okri7Mig9u3o/JogXNLMpcFFbLGPPwVsiWZYNEBzwtVBWqiGnZ1A8aIQ0Rpv1iMh
bj+kK6pAQ8EE6Os6QCl6OaEjaW8UB6PcFVRBaHwaraVPnP6pt1eA9YJBA5jWATVv
SMa5dRMbtXU+VklG869Epq4jc1damX5u6zTIm3q9sUeJ4X+MQUPNTgH5qsqLQ2A4
vMe3PVytEN5Iv5WsgN/+QyXG+QgUg4vlGn7xI3DBlycHzNnTJ5izaYvAahUANw/A
ClDq3Tj9ZjNfSd981y5cRanlDsWWtPcG2XIoS99c8z7ocnLU7HMpdeF3c7rs378u
iM67Fk8IMo0hD+tdbstNIcAN7K4mNpFc9qU7Za1ORG1ak49333aZqhzUg7k9lDQA
+RKblTftZyxukOiGxuS6KVGog3L2qKMu2HYRi28vyeFH0t8wwnyyBe3lxdgPkvuQ
SvQMT2PxpNKG8Okc2njRfbXz65siHW3OtKyh1UN1GrDgwUYalgTVfRK71FQuJ1YU
yb+nxTapgaLe3Napc3dcPocpQfgTCPcEsy7eKaPN0+90T/9wNfCzlEF1PJe700VT
QNHqtCTSjmYwoobrfostLFvhqZuthmWZBTyCM/zRVV7v7SMAUkicqWDOqi2S3kIS
akXoIRrps39fcYtY7QmdJZRpWKyQg2DV/Zh0IeGHc+O3QICKh6uAEFEgvklcKthy
TZMi9DUB6jwM9Df1SmaA9zeEtESF95fQOZL0ef+lUpxnhbeMSva+jD+7bvP1saRY
TdrlEKcqCUO+VerLwkWnQPcRSe3v+b1z3y88zH5df66bz9oqULTX7G6HcNJv7liF
5Yujx9aMuvUP2catYGSQph5OMs87Fsvxy5vjEV5TAFXqUyd/jv08+C8eLmcGZDDG
9vj1WvSrPRfx/oEIM4pFGfRwJGKODQO34XlZi6mPum52F/nXuLDy22fQ+uWLO9Dd
6L5A+iQhHkNGJWrzPZnsWwc5CUNq8enzhdfZ2uthktcZurmldSLP7P+bY8YcvRWe
XSK7Cdy6cdWBuGdxewbVX/oBGYAb1hCGb6pumOj3IDb2Irh9ZnatlD6h3sQ1zF6Y
WyMj2U5h5sGUqVT30FaNjpQY6SfcmBJHf6lijksyZhiMi3rRfsWIJ3y2hTMAFzvg
eFPh9WHzRGQrS93HuVByBMKTYWqCgjeDYfECDL7symLHi1lUVxjV2TwFel63ocpp
14jnuL0kW8b3WmYOPQ5PcxX1r4gMb4GVPWY+/o1tChrHDo+sBybUu10t9I3Yk5ko
+76OZMFdWfo5EWFW/TqkNp//Gv6VNro24iTTUF8Z5YtdvqgSgKL51uj0F/p3aErV
KdcORgzr2wwfpUg3T4WgNlkiVDm1VxCD+8h7sLeES5rfq6GM42itOp4d+mPAPhhM
Kfst0TKHKCpHAxy8GFokhsObuxySx1bFR2e4MF7ssD+Si6uUE/lsI3eUcjn8Bx/x
OYWusm8Lcu4IjIb6op1oKW2pCQUEBLL+dBRyHodRus0LEkQKzrmeoDuj2IIXLiEt
ErrM4mhcj4u3uBuG1r2fo7ejMTfMPpVZdjUbkI3wlA+1kJh2rczhjHBAkDm+89w+
NePL7pCOEyxW5iT53a9mGlbVf+gFdi9lq6bB6dE6j08xx4KJD71G6geFQ9q6J4dr
smYCS+DgJK6H6NAhtf0l5Jv2cK60zp74Sut77ei6JO324vbDnSor4udI9p9pus8y
uDqmkC8N0xp2SFxdcv0md9Mamgm/ICVAoGpJx9aggRxAT4AYfAcnRFNl86uZj6B9
Y1GZnCoTpBsBB+NxfEQUQOqjBZBI/oqbHuNXHaayHPUh7Yfm0dVP6JquRWPgnEbE
VsUQBWP7mCSQTJ4SYSRapouVBJwx0Ry0HCmT8K+qwBFEp2ynNLt21fzIZpYkbUBE
f7PzbYCN7mwUh9ndM+48UQ5tW/7KL/5RPLNk6a+lZCazV8wclycXQNfcZFoOyORq
s8PbeiiGo3e62PdKlxliG9Qk5B+qZP4J+SMFMBPcnX3gGLuCa9VBIQIOVOIQR0TD
OGAkE/z7IAbLHgdjbaQNCk0MIJgLBWXGC+esTEEsJoQvevDTpTZhvByG3lmGXHI6
X5su8yLN2A4F3tCmYYav/wA5z8xFTZrlR0mLKGYtqmSuC8pDBjQnGjsAshXtdS+C
oGl4AuY8hc/mThmYCINIPdgJ+Pyv43x3Ze8RYHKxksDeYlmSZ0KFeFMA3G3ibCPB
RUpEUC/pXnnL1kCRApnhGzIC/FElnDSIosL2X2/lv1x+BLwEnsm69ZAMkQA5bEXU
owWvAPV5q5CafDn2/DvD4/NE3j0Pivwx1FXA/x3RTF7iA54+AnjShEqtvbE2R17F
PltOLzpZyJP9aupMcYXgCVDm364SMFn7QnP0D2//FoT5TwvqSEACOZo3lwXowChT
xiwTWg4LpRMWBHAKMohwnQ8h/tRONqlcEoWEOkj5Sfwg+r7CTHjHS+rTWTpn7vgu
w8oo5S67+wofzlh8OMl2qXcSC5G42JyoIjhb3GxbRhYLghlda94wHMkOX7l3aQQ9
1dNeb+T3JBJiaegGcO7Dn3hKCvWVUZQJIs2878XnzjV4WeSbPkjA8C31o8JzEZG2
pNvIcbX+RH1/lAWWWVp9Bxj5Y23XogcHJjjyM7AZBkTGm65Vs2EZtGfAONEFrpL2
B29siFbR39k6kFzRh+sYz7pmYvMjgPx5FRf3NiQwOlBWK4Bp832z3jpTD74heGir
d/GEbrfUSnk3r2H8uLe0O7rH8Lh4rP4FK0Ap73Pm13/3QtEzvV73iYBCTtk9mM/W
IaQeRwg8nDWzunWZrUbnkHMCGQhjbhl76YVxkQioogR01osmlXwW5X8BTYTGsL/m
AhI0eRKDEr9cWU0M7g6AjPte/9ARkiLE/Q4rz/fWz+Q4vznCmJQbi4BRnVKzvNU2
FINQ6gcJSF2jZj/0TriaoL42hmwjTc5vl+TtYmIhH4Se0jtgF6yZ44WQeHsoEyco
nF1Pj7X+DfGaPUsx6czckQrEoN6gPrkfp6sE0SYDOoh3i3JZF+zYlYCT6dVAYjFG
YS8mgZfE4x86PWnxRc+TOMlCGJIPTtK43f/D5C/ieNkkn/E2axSb8KMgQBLGHZII
DC8pmzLaDVARWeP95k4mu97EG7SP4h4CvEBnw2NuL8t5OR0V+kd4ajMMTR0WVwYf
ErI0BVS6bQjLGJmWmQqdi9ep6TZQ7ILWS//b0k+osuvmZm6ZB1bnFi1Ck7Gyea/8
ZS//eN0/DeSwwIuBG0N2RCg5E0IUPeLjoPK8xaBxMOo/okGs1AYx6uOfpJMVzV7I
VLgOaAX6bLjMdmzJWmc7uEFsL7GpwGxDl7aq5tZ0TzBiqdJl7kB7578k0dR2iPtc
69eDsS/UGNl0Tv5ovM0T6obQjCI7R9JxaYTRn1JH0s8Ur4jAwQjXYF7Q5EfvGtQb
F32huzheoWAg/ZcW6R0WFe+8HMC4C7wEhmBvbK8vJIRghl6qvTZ0+Xuzp3Z9d71n
TFxJF29j+oZINIk7BSKaujilSastajKC741Wo4q6Apw2Sb27kMwKVNV/qS7U5zFe
aCagbX7slJFMveG3a8X6NQjKJH5yIn8xkkd2Bs/pq9rN99j5XjKZuk/A6txOSbAT
0x2FeQ2XLNYyNs0YCx9FehKySsw9xeCVWfXr7r377UMTu768RGgImfMz5F4GuNOA
/74lccl1BK8tqVa+aPR4mYZ7Y+ILO1/aFXHbj/A4k4oF1kRStQNWopOWQoUa2SuN
p/0iuv86nM2pu63675qR/JbR/Oc0bnqxeFjlmHFs0EIPY4Kba1XZn/JowVxVM46l
l3HOLZa+IqsLsD5emImpGjwGlsHnRqGTXDcrAbzZTtJxbkAGbqqjYexmyuSsBCDs
VVta2P1MiVXD2IRzFvGytAhs6vqBToSJNu18bY1bGdRmNdVaKeAHS2seF1VHew8J
2SQ+Rmkv91+ypLgYkhydtjleGNEWJF2L1RowqTfZsLqzvatikBowGaqhMNp3sHyi
Ssdp6GI2/dOL7J1NdXeU8YWcJqDMQV8JEIeQXku7f5YezTFuaAKQGrg4d87AYkrJ
Aj2sLsl5dkfm6G6rb5gRATTDKnYjRv2RN64Y8br7GhGATee967kTZADqX9WnuMK1
lWI9FYqsd80kLZXp6oAtWcFPaio+u6R8/CuT3v51LGiz6VYwYghBmyqomx8HZiVW
0yAxp7+gwG2YrJ75/wdWfJQrI/p/VbHcDwthuCuIflGzVzYphuoBkWNikqRToTj+
OXROz/JYi1jp8zKhVlgyD+5fZnxu+9pxIk/27yFSQriT2/F6q7K0UU0+KAuOOY8b
NwQg7wufcBzLGhoq6vV8wbA6tRaURpIi228VtzELV4C8T2JCy6aRcZldyHva++YV
+zvtAiEsTcE2i32VIQ95e4pWsKWZ8Nr4iFpUmvuu/PD3ijuDJoB3wuC1cXhyaduV
sBA1Qp00yfr226ARHYg6Jjp9I3c962PnoojWB7mZC0xiLw+yBOaqHjqOIdGTsr0M
U68nVIcEu94cAjTRJx2qxWPsxDN+sV1ATa4BOUL+OAo6P0sOi4lAz8GRs7TRu+ds
Zg50QjE5EpJZ7PfONFdGmVmqbWXTvkdh6R3uHbcOuFYa4qDdG7oWN+521jz+bRe/
lBiOr7z/mE/YGwouB7c9Y+btr+YM+A3R977iIWeT4z31h8kdrHcq+594yyUr3m+Q
5518S+hEZVRR33D+/NouVRg7Xh5bCkStEEeYAolE2Cs3cR/uibBC621Uz6wL5fWt
ODuhmsKY9eHjCW3IY1U9wiHToMIv76Js2J1FMt87gqyVzb9aeEgy9xuOPcziPtGU
46w2VDo3A+UPXuBYwGQvE1MJ4q72Vh45BQd7VYb+45DvQ49AIz16QdtbO6n5fe1M
0hhB+9glWSTzfYKl4OOdS2QQrn5sPd4A8Sov1lXx0OyBfH2yKxKGXsN8vD5tyKwm
KDP+2UDQEvVrf5bJ3x4N36N2jiE35IJItuqZsQ7fDH6dNAU8x1ChoZZ8nluUzzms
2s24BRKVvbz+04qpcsgQ4ielgANh009DlHsVBPt9mThHTm+PKTCCMU68PrrZH7d2
l48yonhhb6tP7ce/+rrQLDkiIQRoFBgalgUR4zu2m0GjSMrfO7vvBKayqEvtl+Kb
6FEnn8JUGZ4Qyl91rfs31MsDKAHgdusAdnllPWLIGvcf9CIRM/y0XFexPLtTavFW
glF+TSew6FsKJgnnZQYEOhELN+bwXfPojTzLlDEvpZ1xbng0FjAm5Pv9RUlM0f57
lL3Md8PVELLxlbld5EiXSD4gKbIYz8wMBseUVd2apAtPDKYy1N018mDCwvJr5Ha4
jKYO8R/jz9BwPF6p2FBv+RiA9SQm8Ph06GA1o6EFennvqQYUZlahmHQ1AXakBhej
37lz1mqyQLeubZiHjJwAxFr3TI7pdsKYoeOE8G8E+cYzB7co7qtPamwXfx1Av4+A
/af8q+XeBLZpS/f3HEeKv8Jq5wbErJ2vPLi3KRe5IknGLoyeguQpVh1y+j15upO1
sblUKfsvv9SNgWs/wWwPlwYzND1srH+R2TvUB6BwtjpP/oS0Xzch8ylpQDtFNanY
bpybNJK7H8Eli7QrYIJJLDB+/IJ9A6SeXF0kb7jKFNKCpx8T16O7aOmlyQ4KoZrK
5j0QC4tbTgnNhcTbP0TLXgRXIdLe8RlGQwoQdXaOSvtLT3uL2+lPYuvngPyo+nex
M/lmHvO1KAd5ahXWwX9sF2+FKF3vPWTctJLSypH6a5Kq/ADVfKzh3YT/z0beKPbG
B0FNMluRwcLdry1RlBXo8v5OF89xxT9SufauVzgpF4SWmBPQTCUxNs1QOBJt/h4i
3DL/XWS/WXYEIzusXDo5rTV67qo+yzwONvP99cPFpmTyX1kjP71VNMaziCGQzg2w
7NYAPS92WKveFtWhp1a3VrBFsl9Y7Ctk83g6QtFDgTZhRSU2UQWzB38QTiheku01
hYYLyPRorhxr+YQu0l48F0d+xHL3bBdmIWIVm59ibnI5lTNRXOFzeMkE3wKXRm3X
5W0bb1A9q/ViY0w2Pnx65CPerVNjxqSbbz//AwNI+KPOBBl5M1oaAJKgcMuzkEFr
aNoQkpWrKYZI3YqHq1s/BcBh9o5f+P0vjhmjlHsJk7qGhovwD9d+Tjm2Ew20Tsm5
bBwXiaCzvyPc3EPmXcxG0vImulAZxb+UuzrjMUtmNZCqPdZIsiHqDombJiEdN1is
d8NcPu3lxJ++n9EcfIpVksXDwYNT97ywca5mrC94+wyZk4ESOldeYx+AdBK+ftw9
w4giwep8FkCezSlgbEyuEFkiT3FuTFpzY73XA7CJIdAxctY9f9jmgU03F7KMn+Ws
cawfs2/LGB7dr6cQ5tFh4yiuUqmFKFXeqEZ+0t2meVl1fTf/UqSt68RnUgpgBFSR
poAQFsFGgNTNj/zMQee1ZAzKTLYqQMI4Y2fW87jolrz6LNoV/L8A21+hsahwIe7Y
v2R2FLokYSMZBVcfkJFCPadStueKJu+F8mL1mnXQZV7a+s5/+xwp4q+26fkjfUTL
cF+Wp8+PjQVSM6aISsQ0pfmEiRP68pFUodKaSomWyBNwyv68hZtuhNr8jZAnIyPe
wEDKCV3K4LxKs+vmNZQgnhaZbQJO0IbYYbU/oWOZGv3UZQ1zTM4DBtCilJ8LDWQO
ea+JgAXZpBldpAHGOYpZjC8Bn9ZfIYAtpw1q4pgqNz2u3FgTpAuqcmUMz34ZfIgj
FVVAVJqFgDk20oDohynRx4KZt+yahYK9+TSvdh0i3g+hCgWInNvME65yWwDVZNNF
Tmxxno1sYbIhARhhO1ynif+MYHGTdvl9SpXDDtZc8PaP1V9hxogh3uRqd040eKJh
+9Xzopjmh5KmlfQcqPo70RDdys3ga3o8KEk1coeZ3wnjupIjGLlos1jA068ptY2f
TUPtrrjiRDGzc1TLuEHZQPwummuSR22XV+PRbDts5YgM/HPtLoq8vYXslTphdI87
VJUBw/C2afu0k9JgT3ykA3OpBpVzhlfNEryQovDWowOhrXArlvk5gVSNMVnhW8lh
OtlyzEpwL6VV54NmC2sUHcr4dYa0fvSYoJEY21Z84xZOKPfWKO1xNcFllyGGlG0r
5JKswN1kD1P+8KYt9VptUXIv33Q2FeQ+tCapeUhoXcXedrPAOWa4pqai5B3zRTTg
psuf0VA2DC87DoZJwrfzcnhD4fHtbaVJhSvaFhHA91AESwZeD50cXU2R4TFijZxP
kBarxACXMajoMivDn5MSIjgy0L66ho3NHSlE0ks7mkVgoLtWCMpSxTmx+7q3tR+3
KiqX70OPCUH0B6oSrKedd3pNDK5MhxUPMfxlHje0U6R6u+U22cjfmQaEfYVzkfX9
XHMraCjJo0KVqwULsUgr2mzh15zAXy0kFx/EMBBWvPJvcsiX6Mbkb5NJt1UDEiTO
4L/Jve5WmKSVcWDe8d3nslFXjToSC2zGmHtsiOac8n6NuPpG501DiJwyIKWjlruE
Hhi9JRWnSLaJmTrj4UC50w5PHrQsBLD/vk5aYgKiMJ+o1BSo0fTOcv12XRhjuRhD
jOAxDm+P+kMh5Xn0XXXlsDIgGybqgwm4Hys9dRbqjvnTFCj4VK2BO+U/B7ph/BIj
Eq0usJMAOFUs4+qbmtkWYWNbXQM/uJwDkBGs9adKIjV9EMbFyyIacVimoI2bl1L9
qV0yhdq3Are/oFvtQEDga/5Ao5TC3Mtv4+q2TqbnzXCuFiT3IlsM+PDISXzxdXju
VGNxGVDD9RS55clAwacOxHmxZYcTitporfVD4GJHZBYdK8mtjLqm+l3U+NoVKfA4
EE8DrvFM9Ot748GIw6ooaI09KbhAw2FHeOEEfIEOme2CFo+U4fGFno4qPQMXhN56
nHsNbfu830mJug+qgqKh23+LzWeA4grS/86BIcDOoZ2ZC+UDR4+HHeSx4AMT7Zew
+2dNTxijldcLwYTNao9YIOV6HvaUPG9IeULNzRrL6Ej7qFQhzg0obD3qWwsUv7XK
wgnf1RejN5NDBoSB2gZK6sso3+raiDyLwirbh7kBh4rFtMUKu7ufGRQtwXY2jcgV
NwPwAjiXn5jBzDUd2MLDzS8cwPsyeESIQNfiml2w/cJ3mPdDXr0oqF6zBRwiyvZn
x3pJu027SNkneiJ7EwwDD7o0Ct9HQWC+ZtF7SNfGNVPzwhQUPXrzhABSL9QyzM+M
Gb7AGDdBIL06gAmhFVuCHqPotv40gCtKRR1f2HTyi6GpSL6x00B6X9MbMlm0yXH4
e4iiqsmVc2MrcEsu3oNNEs9atwn3YN1KWjaG0ZVXtG76LVCr4woodeOXti1YPrmc
dBWEcxjqpbSvWXBlQyGOklC1+/uanUdlEScd1D+y0cbtsqbEXmeh8zhe2Z2TwQqE
JaUOMqZLftktz/+jkwCncKQq2qQiFeyQ5nJkXpJhYPjoVWf4YgZZJkUtu9Q7A6fm
i85MqjeZKe+VzBX8tdx7XN8PYMtBFGSVqI/bvXxTA82OGv58gHhuortQw2hMlEcK
iEujJ8Og09pAfTxHBuxMYzhc2n/OPLoBZbrnslYpQn1OdWcZpABt3UvmL7JmN6Uy
c5+sUzTmzz8B3N/VFNShZHDVBM8XknT0cmllK8h0syneY/h0K/pPKQR8yYIXPoqw
qNK0wLaTCsqP1pRHBroic1fD7XLgC6h+kkXLa5QHQJ+FCd5p6A63/mPQhi4rqIt5
svu8tsp20qKozs4ESo5/YNpURyXDpd8npA2wVrJph9eOKUoSRdTM3Z5gdhApxyj5
kani65JdVmVLe25Fg4XWnelvp5nh3hjr/5UXxdrQeZSNuuSNPBNbnJXMWQsST2H3
4lcpLaD8LlLQjAh1ugGgi8DI3iD99200nMdvP5nzsxrc+QzE0WKJkhHVQjOHwvJU
8Ze9yFzT4ksmmCb7gDMnFYxafsuRkbilI+ph4LOmn9N6REl057RZvaA/aF7pFf+x
pd13niK3vl+ifIWRHNaIUmBtpirFHKWCGwR3PMprF53reA19WbnDiLCnQLkbmGS8
JThsLxlOG3li1mt5xlLudrKRF9cSLNUXsAfS4gPsZY5xWhbi3cUaRpXeyaBAC8Gt
8mWsizBIOjL3AGHckLYcyHKL3cBeXcp34ImBqYqOv3zUliOpLoGr6Gh0X6xD/Bp6
yirO369RPsvtgrLuR6jZicwhm0ATAkma9VdEenQXdlbHvSnNKreg/BgQV/lRr0kV
D2r9vCHqVQdjtkLNGSHVphvxVPBeNoZBH87ALzHqbpk8KE9oqFXytFxJjruDU34Y
foGVoFHk1hIH7BUzadNCSEXBSbjxRIZr1snh7mSfAhYsq1oS0S1clK5DV/H9Ivms
CrIXSxhIhCfr2VHrmAG+ZNxsM4iE1OIZneXk4u2UXjf6FF5HOANFdam1ccKHo5I8
bd6FEl35FUvczqhY/C0ZeDkwwHlXaP0Kp5X+CIQNdab4dj6KW7pGxm2jsu+3hsiL
/QfxWQ9uWsP5pgCv0phgW2rcEfUYZsmVBSmmtQm5Z0pLSK1Dpx/DrmR6OOpCJTit
z1un8DAeRItiN7p+T3lSTjiZ5B7iVTYxhTCxaR2ufUgf3VFR0NXooEXjI0saD5pH
I116Z6lck1Ert0nIwVizHBnTUblD7wLUj1K0jMKEzM7gLZFsxJFyJG9ieA588An0
F1QlsXvXWmfO1+UQxUSKHd37hER2Ef5Csf/XiC/JgG5bcPTRcRCGq0Z+DzI0oetm
mtP1oOyQXQfKPGEcklmlwJpBL3hsMvB77+4SBPJA0yXzhoOFFfeIi4nD/yDfqVEP
TMsXPpQO0JdXV/OeJf2kH2NuiyEX7rOca1LpFbi8iUmAe8bPgv9U/Hj4CJbftQ1J
T7c3XwAHAK7uwI2/TzNTjeVmxS1Fx0wkW9Sia2yyqV8dCo2uuwz6biRxdEr8L6vg
dy5rN6Kofx5X4dnfDgb63M9fNGYrOLvb8eNkSQLDG0NMUOZ1KKXL4gOpa8u6fqnw
ju804YZPvPspILkdtRdnaAMCfXprX56CjzYzQPUZqp2jWG4srMNW9EyaUOEPHnyU
mXmS4mfXSsyvSu41h0V8rHu8FqvM43ZbEq8ER5e0n9D7VTxFy3BdzwDhQ3Zywces
KoCkt8jijqQEA7sWFm8r0ai8ADLJx0wdsx4NVoMaPO0SKdkSBlIAWOj662tpzUrg
ZeQ2kd61lCWvaHqf2JDmuuvcYj6xcZM/hiUs0O0q73LPHaNiVfC1EeMbQNgizdZZ
gXvAYjhOUGF7iXrMzMKFPs48wbw5G/UFEWMUJvEmzVcm1y+4fcWk8AXzIm7yoIhL
NqXaqitlVGgcPA1bmRdoZluANj3Rgtqlgyg0Pl0/EsQnsdTSVsJMS1FsyzgJ47rA
ifOeSnvbgu0rwGL/KqE6OwYYmOXSePsVM2iqjWT1ERm5VK1lgVBCshvF0TygJsdg
st1hb/2pqajHxy2birsbQXB+DQqwfDkPX2dUbp3rnqxTfUH5V7WC4LkZ22tHrVdd
InqXl4SOYmpnble0nnc70LFhlRXqmlXDQlZwyMK6cEdStectclcxv8l0IocIUW7r
m40SttAbCfrLoB/yg5Gv4dPHvMWJOMRk1h2cK4GlMQXUpqAF1FuOQR9G6EDHxsBJ
pqd2F+Rq9b05sqXVyWrjr686yub6xFZBXEcfG8/CdHMUKB4VvirDP7s8rj7+x9je
4e9JzKP4I27NCZeuSXgWflR9N+ysSwkAnScdaTIggkST/eHiocSQuuGz4lFtmFGy
LbqpSXzfVXEpKSjMrHM7NQEY52V0szKpPa3qUdxpttJ5F8kaTrJBgSa8Yk9BpM+g
Nr7hOF8R3AHMej43DjolYoE0eU3IAUzp8k0g8TqLQmoxMGDyfH0uLQjYkoIx02W+
/gFFaDiNeEozRjyW6Oo+CQfZ17FV7sDwKaDyOK7ARHllPPTCx37f7E14q9hJBSZX
ey/I+p1Xy0jIXgxZmKzDBVQIYRwbedv7QF/E5+NWtSZOJTpEJ4l3zmKmVgGgJUtA
sxAHzji5SZMF4eb+FHCF1G8IPFKi5r/WgE1CqDoej7cTAlZPdwD2dlYNNqsU5dtd
zYNWJJvbvpEkkHxDe1OJJNjVnFuM7D2TQelYbjDnTSDsVynNwbDhp12htEJpsD3z
Vy4j7GS8usiu9EUZS1T9y8S0fXfABvY4UCRlMVh5YgsZftUk/y7n3nMmwqHttCL2
JIgDUa2g4SjshLECQG5vWzp2In2c4oHWE9FKW9z75PXrzX868DJfjREnIbXr08iV
8kZKU5sh6oNUR4AFixK0nZIoazxkm+hiUHOFF4+0KFl0/YKrc9lQOsyFXJeWmRIx
dYiAoYOiCrHO2yxA/rRG4HIaziX1pVJsyjQsK6JCNv9QGwGyOfETrHC8UI6CDynR
J6yNyEw9PywzmT+9bw4al/A5fyF4BYZ5JPFu6ywkXT/q9RebRvP4RKMUsq0v7Xqo
t4diLQhk7DMzy2rUpyDHZ66SLpJt/Rdzrf0PrEglmQ4VakPml3s7s7bmv/vN16XB
fD49VNdJ3NbT4hwLBU5fxsKFPW/eK5phNJSnuxWVUEx3KFUtXZIFqrotjWs5MHOJ
onybu4Avwj3M7Nlm9tJ6hOS36M8aEh84utKJXkFsGHA7n5p1A3ny+3+leQQEdRtO
n0awDK4pd65GEZYSVUwT0oTWLiWE7BIRyq9MwJN1hRnVX2PbId8C5BNU31GykhEY
vPE9Y58OetIBP2/meEUGy/jLQwAQN5g6eNeaW5XUfkhNyZYtcCjcyFJflaHAhBD+
qmkfVaUGbqaC5TLIlluPzln5WLVuuNtXxR8PFT00zTNfVuDpFdTs2ULASgWt27I9
egGQEqdvaIFI3m7+VIoHLDUraxUQDmHwcOQB5OM9TEQ7q2DarsTCJacZdu2ZAh4A
0NPRLGjdH2N1cqs8xndbBwyBA1H3RSVSbcYrkKCBUzUF6jYR24MVUhS0Ie6Gzt8V
POOfBW/Kc50r7bmNY+q+yiZ1k3lVWISWksMHYijB5GX+VzAVi+z7huyS5YVyj60k
BQVJKnGjgArgHMB5G2YF8vjrWN5xN/kwg69i3DnganKQ22WuPcGkvQRRibt0eEHd
ryQNgP3nIcYWY1wB2S0uCG3nMeZ2GvHcpJKJtG3QaPnqcNIAHDtPLRhIUG40P5GX
pTOqEEgbnNM4RRyU79VDPmlyMCmiUf6OM8UtTR/jV0UMZAPT8BGUnZYS44KR2r72
BtqyP9fddEDxbv9VGrmw3bIT3VrgmZ+JjQxJ9Hy9Qx1aoTIKchMyTNJLrLhEpIEG
Cg8f1DxF+6fl60+TQrLbjRnj6BwEvvYUClOpAzICmfLWG7/7wn6RnMo1deCyZMYy
FwJhE498hAApoyRQGtyLErrw1gckOUJ44zgseCThmBpfjUXeHtSytdjT6VvtrMll
NvV+P2m96KaqRI+S9R1ZJZQ3KlCzjYAVSqvBIgn/idhxJR1qFN49c6YcXDksxrbR
wVx+YNvWnUM9kXpiM6rArr8YVVWCgHzs9q4hQQZQHUcF3H1HJzc+RXvOINsOm3nb
NIeZouM1TWS6hFDH1AbEIR1nOcpbJQhgDGyL1W/WUuhj+8lPnY3ZQRLagpvHXU8C
nccWE36bTQjXzIcWmFdh+ktCQ3P59HgeRPbSPnD9nIQd0WXBYaxTrqmrEoNdad8a
Yz0iG6i2gKvUyP70Xr6rtqnUANs+LoMdAvugmOvKipO7glRoTYTSD2sSEqbnHRfW
LXyaFWU5pU+DuRNb/7c1KSxj9EVDSCIP4/GrD1CHneD2jQF2hkztpPsu69L1w0Mu
wXiHv1wjO27TRG844ponGgUdDqXtcrzxU5s8fcUY9l4s+FgCM0aLRdHZNlXaSdhQ
zPAu9lA/yhUOUjO4ukiL410fPH26BqZ9OVD/wDH4jk1ev45Mr1gdnT5L7qew67mF
DFUofA5fcFDF1CKuabvDw/ntFr3ydXdP+qUJXAwD5G87xvzih4zbJQCiIKLAHcXT
sYag2MpA3qDfaxR/CyVs/UuPyPS5xvBAQfz+PQmtZ4kO1rUGxxoDxXx7eE6J+Pox
VC9zS9ey9LOVr4jY7VLt9zAGAv1dZyWXGOfYTCblXyV6SmHly+G+jHz1Gj3geuR2
gRIVmCOG6l+EpqYKhEOriJjUpLvrmX27HRchdJFO1RyWPgpXYGgiSoEXsUq2wiu7
jQT6QJC7KfamjWkat01ugl+KjNEx4gMrxt5qr9+d5vXEoqm8uWN3M27ssNgaTAKS
6S4oBlPF0yGAIRl6e5NfLYOMb3WCaUL5jZHvRNwi/vPG9P1r5ETimczG+HkCpzEj
dg/ZjNYuvRRz0NTWfkibewl/FVNWh2A8XjGu6305RXiTjzJCGRpiBZdLf8TK6lrS
UJu7GlMvD3HTLNsjLOdctSIATFkCtpv98piJnJutR7KS8VqiAv1iPQAB5zXneIwP
dWm8kWJAVEjHQ1taWV0NVvMnkMQ60FfFSI/tSDdXuUnufxVV+6E5j+KLyGe5jCzN
iqoLZBOhp5efkfCm79M/AFZj70wxNCdKyHCx3pLkYRH701Ot31t6dcEiqC5ElO5m
L+Ssy1Fo0ltbG2JdyWZayQbXEFHF7sbaix+kCXaUala6i3/MGSyeTq70eURdchwn
Mt2a6iU3L53uzGQMZGGSpas5r2pb6z9JZqD7JtiCbu1jxizclJLCHp8Cgxr4jKMc
YHTRyrtPCHpA7GG3VkYytcQVYEVIkPVrRQVPeYnkG8ii02O8iIJWLP+5lV0btMzS
XMWd9d+JSchHp86CAk7g2JILMjSDywVRCj6XNqWEJmsfHUKoKSXjRHQlEinrZYtS
TNhIB/gQ/8FzJ3yEb2RoXYzMnjlGjRsknqoQu5GmhOSqETgzYFd83PkgBQOu6Bm4
gQGnyT4LhIF6gKTZPoDN/dq/aRP+WYLXY4tXuvYpZhKtwslmVq2wjXZwr8Yz8all
3IMSa5LZN5p9vNZw850KXRBcQ2hQ4ryMVlqFP7cqrllq3RdojapVQ6ssmu0/Poi8
Vyfkgv0qcsS4yLMg9VSS927Q9FhdkxUAlxGJ5/j4EGyjYIqgj2Ledkwcm8E+v/3k
P4B3bXmppQTMnljPo3q+eX7XPFfb2jtvbM+hUaVCA4towskHGY+FIdK8iPy0PVAk
Kyg0+A4Jlvz+cxMTXCJsBXQujtSDshw43F6W8N/8aWPhC1PB5REH22sHvQZdWAH3
kvvS1rGjR4D0umQx1yCI/tT/RmpszqVyJ1syblQjBPV6v4FYBEgUnVbEfH9GoDHk
wpsK0/ztBogb07hT1O7XPZN6osfmqn+SOFRvM6DjFgjk9Aa8aHBl5SfbchDpttZV
l7qAskjFs3N53Hhev4U3lRb27u7g6kPfnjIqhITiURkaP1r5evOl8pHbxZPUTxQ9
7P/6noZ1viUZeJhA+mff87Ooldf6k0+nmtUFlWP2NCTM47tSs6vqb71v2RKWLdb4
kTOt2F76pq3kb3ji913XY+eB5vdPAduyM+trlEI1dC+AP6rsJGleTHd2vA92gWQn
6qonx03+l14RgkqvEXu7UE33O7WXzyj3Mggc2j0IDf2uyQyaDgxQjfBWkx4WaFGI
5rqLLwtvrvl9I7ISfhCNwDdB1A3eH14gB0aQTpC7zpMC/PTslxErHmVCC4q8B1CM
tr5Je3suJr80n0TfOMpOLUo99YiZilOLsS2B2zb4sVbdIEVpGPscHbJXMs83y3Zr
LPofCbBHYmc5LFJQWtpMRosvAWgMAbNVehSiHd7Nf2wquFWEMgrIN2x2LAt/tYXN
nxOh7qxqvQVp9SyeAh5lsLgqkR9ThvIXDs11z18icPBu4FRg/xAQkDXeb1WbZthz
ZJWQfiYeJwVb0L30PNnmF/Zh+dfSamTZ1P06jNbk9du0Wi52xNwpKB/yLHqE8re+
1exueoUyD1vplGp8RvfBNhCJJ+zQWduNL1oMvDGoOtdUGUge8ugFTWnKgSgLIu1K
8lgx+5DY/9tAlt6ywxmHU1E3p15MzeCUBJ3C7T19myvxHOLwkiuKK4JDHO+XjXFy
GN/B8QJ4ukvJcBW/52V3ExyhMJa5Zh60+8XMB4ncXZmvzK2hPU1UU1vdTtbTmmDH
u0/xcwPkBOQDKakO6fA5WFSSso+lEh4hCxKu4PkhsMVVhmNwB2/SCb+IzfwGA9SO
5008vvKlRsHdLgbBYR/+6XWA/W3eGjBaCTkYJs65w77hBtgFK3fDzCY9A8SVejPe
cIqNzhDK1ZgbmUMxqwvsjUHuh7HXjAp0LeRpxyMaA+P+2uh1/PNaYx1L4xnwXWIX
cL5ziV3eyOt58QGX1/xVCGHPBVQretudoGKZK9kRBYzAiMIKErEvVj5Gw2koLp3W
hOX9xAfUcb+SYHYDFjsSR5Rj8X2NEfzBf+vKc0BvL9+jpLD3w/JNTvAZJfDSkGAM
MeV1qoz7z6Ljz3Pln8AWtp4WNeXF6VPRq6uFwAm26mNQur6K52QYme53YTrxu/tq
emA2olUVg4sYBVZWf/TzYeHXiKPZWb9KEHjB+zCS7ZH8GgOf0x4ZKDsEsxpoPmhu
GyutEdLoymT7HN34dHV8b1efj7nwpkSHI1BmF4ppZtv6dHMutU7AFGK2LHgWmyqz
IJbSmofBiIzAUg09boXBHeM3pifCwu+UmOrUs5trlz8ZK8VHmWHjOTHle/PhOyuO
FyWWOgN6XbvAZVpXD02FHwYhbCXSrxKanmgPF6Z+ne1IOr+07P8g8N5BVIMw2XEu
weIjYvmUMeJqnXN/491eFPn84DSG0OS53fxM3dKW9M05Y7+Tf8TxNWOeWe2Gnf40
z3QLG9HPs3/TveQmAXYbpo7vdl/TwIRlbJh7jgDHfUHKAtJnloyclAxNtw/EEjIl
6jG3cp7oZayTqhTHcH3cFinF5ANq7fHlgiKhSmzU/tM2xiN8xoYldLPa5YNagC7+
B0m21bHPcQlHIFjorHo59Wj5VSEJ2wyOeb4KbjHl1Xz+uRmlteqi+Fk6XeRUlA8w
t4LQBjWZu3ebBiPMBLhzCkAaB1N736FPQfxu8vd39eiGXhcUsm/RS8d9VuWqXg3M
bG9ftC/atbg8gZ3FEZRQiUKGMMuU35yMe1DxDXz+ssedA8vTlEWEBNSa0u/MeJ2d
jo0weAHFB+Y5LNntVieShj1Ghifgstr1CWwa1ZESo7huojynoO9jMF/iiYkWovTS
hNPGyHe11vIrMzoFmva5+Ke6qON73zJx0lkJiZLG1W7TMXVRe/nOqv7cMdwvFnN3
QnywpF5exDRBnqREbHP/5S8sjHtDqm9EOZlinb3/5k2670YNTxaWo3xHa8wiSQot
wIgNhStU1C3/s+BfOguAbVdBT5tC2mKX5O5xywtCJ1yQzO1EM7DOCwXddL46kQa5
514Ci33B/g0WPGs5KA/eJeQ8OCVSIgo8nPQ7nJVKtQVpL1EHT40Okjjx8nftpNx/
NVI1ESk7/BbfBF18zzSnk/WhJwLHJbLMBMl8+nfIXRDy7gSnLe+q3Vldi5Zj3fib
t6yLaZ3c23kJyIPzz+BGR0dOPrPEzfTw0J87m7UPayOnAf+o3QFDv1Zrs0O4D4I1
aYkPygHPvmqvydm5rq8Dtrp0lTiZU0Kbyj6nfbUjM7PE2IXiX7jEuHAGMb6GZmKv
H/EnujOqn4OMYoK3eQJAaSQehLD/+qiPV7UPkNNCw6QNuLyveuAA7NeWBTAK44dI
jV30Zn62DbYUME5wQc4TVJ1wZ4JSMdzxmeyIBoCSzRMVBqIOSr/m0RedU84Pcoba
zcOvWHkMTDF7/QxP6Yslvk6IZwxtwhgH+YE8g4JbQq9/8oIU9WrCo5ko+DnxS6UM
n+e9iPeyHTYqztbCE3GqxpHwGW2AsVeGF9OnhStaDBtP3FE9SxDltWiFxTZj3vV5
2PZ3ly4KMWQvqXw7lo9rcAgo2gdGof9xfOgEuVWwMLU0agvf61vHHAaFrrMM7B6D
EsWfdtYrbf1gwE9r2JZ0Em6RP20/zPhxs7p2xG7COdi2BgAjen+oy2luoJfv744I
y24FsdlQc4yFOhKQDp2s8fvckf9K2NFwn+vwtKpZ0S5z/xfzznONcy3DIaWS0J+F
3+UkIYucqUTLoby+8By9Q4JufXRaeipE+NZ8EM/GR8QK7jqdX+PKlX3lesQ2wrhm
XnQ0Fdxclj8cfBNduTmIzWaCv37ZQHOYGhjjEnUD/isL77veU3WRImYkymPghzG3
ikosnlNnP1fJ5f79ATN6et7pWKcweeDa3AJn9ffD7idJSm5Pzq1V6E/dIpEe/OV6
jGB4NCQPTt/m+MXnnryB/9+juMgvDZevheLJyWvp/aO1zEhlFN5jpZn3rmMfbl8E
sP2SdSo41db49U7MU9XRPI4FqbLRSpR2ZmYy0+RcDrMjWq69U6FF1UHwmcmbTDei
vpmYdkE48EINcGKs0ExrTOlI3ctbOrS+qE3VTEoxIyTGjZLLSU/rFdnmGLMRxLmB
Gs/50+4fzFJgurs5JsdfBdOPy+wF+lhlI7k/vDbJJmjKUoCfi72jV0/oNfFJl/3i
8AxpOgapDcMuXyJv1itBOwj8aVfs85qB4UrCrsVWH6b37do/Oae2ZrHGreyDl1kE
Z90gdwAa7PNDWJzS9mADdpBrlefpZIIWxZwNEiWRDymefeNNs4fU6pVzZ4w5/Y02
57Ee/qHmsdsoGzRTbFO2pqxdyT+B300xpubrBQCD9hk8f4U75zqBess41LxqCCac
b94KEfK+3tdo03XSo8rSjyB6jR7fJ0ELs3+jbvnB6BTTijXvKGIJDvvSDYLoEehS
uTrsedV76+dEPny8yWM04QLjoAjSKVWvD0w/M5jamAa9za1vL80eSX4tM0FdQ6eX
y61O6KiWohGRb6MZrsKmbSLCH0bHJ27hPred8bGbkRKvOFmExwSuC6w0iUPnrEwT
xPcW+5O6XpxLKTlvrQnIP+vCOqyO1PpK99taPd4/tsQsUFB5baBBRQmt8Mbv844a
OYm9Qer4iiWqV8q12bzW4neq9hkRJogMQeOeiJl4XujPCXQlFae/sGf/EcrVxnYu
w86t2tZm9HUWSOQu+7duFRJSIUxUwqj7h9YhU3Wy+Zr6zrkXdDo7LVFE2K3kxdcI
vyMquFPJJAbWMd8zSe5fozKblnzYriMAz/IGlggwny8Lqfo3p8wzkMxfiqQQEKat
QALgrC/nZgAlHnu2yf0deCkjl1BnI4Pjzy2YaeKeDCy47yPZ4+8Yy2TorMu5qbjj
KEIlZVjLI8KZ25/LzAWzuGhqFbH2bWgzODDByjOIqjIQmSh8InfQM4//fH5t8kfE
RhCZ7vdqu+iuTcEWo1u/98ynOlA8CW/AhJCDYDeu+uxo7fp/MAuQR4Zimd9hWIWE
jymZd+PMZtmKoGpDnYeOMWATlKUBZoV9Qd9p1BJeJ3ofUuyLt+83EilxKV2OD4Sk
DJIsZpQfiYo3VacN6nXhUi5jMV9guCm5X1VDC7XqfHZ3+YYKgfxppWJfItv+p8Gu
iIhQq3WkDPoPDyzIUwZW65tp1Ns0Twb5DZDkxafyBaCvCBoz3zZUkPWPJbMkCGs/
U2L2apUvKNrPQf+oLYbteQja67RuTrtJLPcyYQd0FMDR4FrHq/1pgOegf47GH67L
leOhIxPhTtxBbnL5fGQEef4nUp511y/hCtsmcasNFbeoMSoZrQ+kkkCjLYn3HOjT
zv5nTWi1QzOM7Sh5GQ/z2uAlpUDVAt/4yfWYsnMCmjZAG59b3PpfWMFlKJOfAV4m
73SAo0BaJVWBLMsehlJ2WTtoHozm9/tbJ0pz/qICFlxIfb8l1Yk/wYTCZCDou1Wy
P2WHobKjUgb5J4DgLa1Bu70o7OA1ylB9abHSjMQAE3acYwnIcPKGQCLUxphy4Dq4
opqCmzWSayG5UzERLif4ThOFnEOZu1tEV9Gz4RjWKaSfOmA1qDuLSSypcgOHb+eo
jf06a1pbh5TCeKpGzrY7489eoeC+usDjGH/6Qru7hM6U4YNj/CyRao2qd/DrY2cd
trN/baAj7ifnhX+poGZ24CvaTEACuZx2mKsuEWEuks4W56KhN3i270xzgjCQZ6vY
cI3yxErx6fvf3hXTfROuQS3+hZIS2Xyynylm7DcX1c8iqHNSej40Pb93UgkQeB62
fGjUca3JWIDutfMHfblVfqQ3hgBbQ/ELvn487fpC/oom/ecNQI55R7fYwxkxZcBg
QausBUalXShyk6slIIjiy8mMXgMWoa/5QyFqA0gJfbBn6hn06E8lpUavHLXAnO8s
fDrLvBff5XVE4dVpqoLVQYWhyxOxc80X4CTLN3TTWPrjAnWcmZEC3cr/2qf0iFGc
eS3zCMSU0LuSIwgBIDrCeUBZXJczJbg0IH+r/cx/YtAtOgAUlKXq0b7i2IyL4ucK
varW6qz7tYxkDTv+jg7Dhn1boNvYnh4z6pOCPKxIdKyW9EgIpukujMUFY3Irbr8A
noigXxY62GZ9oUPV8UK3oFDsTT386K7xOetzp6t755B82yoMMKgX9xsSGKkCty4d
S1LlP5ReadouPhvlxJ3ekY1wfxT3ezMsJkZAAAwS2wK4d2ob/sMFnulOVC14L94E
qOnR3yZsJFk6Dm+YhB8nXC3J+I4fY5rdqBgdqSw0G/kUJ88dXmGgZsBDriuWFtUl
Hp0WQVn1m5kB/jMzakjhtktV/1wYSwYCc0j7CQkEN+orrXu5mWUnAqbecE7xM6VV
w9zS7GCdplDz4ClFha6H8ieRqR8XkosEQZpt1Ts+ISO1SEgMlV6gnxjzUsEXVjqN
tK0oyzq/2JqWzwo+KJrBo6DsAwOsKtZ5Q/Vqu3Wh904NYEH7jnAfW9TKTxIKnGW9
yjLqckfOW45Bs9Hs9voW0TMphahOoldphhfo7v6cZQaXGn/GLt0U5sV6QbFT13wM
723j55+dpq7t+ADHnVbKFLdaWwQ/BfijcB1+GgpQIF9sPfXfP7Dxo9u0MIb9F3ag
pKeNvInmiA2nlo4PATyPRpWgxEqx1nQARr4jXPkx2DSSEKySFk7tIEH2jKT1Vj48
1KicFySWcqX5wv2U9YtxL94dOr2RTrqtviu+7ynJnZlDRreoZBHD0ZgyXXbofGSY
Gl2RQfhl0f4bkaubxC0cYWB7plHIm4k2nVd5gToVvEbcD+AHCGnoVu8KxQBIP/8t
1xGqIJTwx2H8cxLWCl82HoG9Vi2wYTAEspNJtVMpwJHFghQ2JXKKn+BtLcd9r9JK
cjJeOsCteQu2iFjz55lhTO/pBzyelqe46OP4S2BnTi38YhC86OxrDm20JktXW/g9
s/IEEtd+39sLnJiQobBkWYhnAuaN94weEk6QPwvaTVpL2Cko6yZAivR5uuUM3vmQ
QqksmR+UzDTxpn4atWkxud/fPpBvfy6jA+l5UMP0jdp4C0+Nh3nnOxMfwgMEVhV3
zJT9vykEUL02OO2hOFHaam0YE6Zc4ysHVqiN2zxSIywK966WOfauM7+UEd03qhTj
UbQAN56gsAHksgzHx68h4fnEjvqjqqEFKMyIdng+zkr0sjbCPlfOvfolP20FD480
I0JIYwTuzPiu6RshF9Mf9MYyG0O47zSTD65sdA1mgxpkJ6bluWROAZkuSe2hhQ54
zPPFML9hm5TKE/qle9+c720Xk+9EHvCiNiFK8tFzFRqATwubEEQOfv5FG9ddF4eL
KjG94LdzMjSvG2O//8/+JdoLTeewUaVQDRE3SMpIanZN6HyuqCOvdQPQwdgNrfpn
WbbPn83UWrk/tKESmBWcbYzMLNz6nDuLcJpQMLpSFbVmTFRJktOqO+u32inEQgmI
umtaDXLIwUW/KFkasmeSI71sZG2/bGERUdbEESE2u69Vyuv+48N3pXcM6ZVaZCq9
FnZfxmQylg1DS1Y9Xor7zfi89GAaUwC5gdABRtWbMkTAY4tojLuY9rHkhDM+V+oO
IhTVhcCQmSyFkWcBCXSPzrm9DGtVm5QEBYnHVlHc21/NBbRGAfYLDSOX0fuY6xIr
ZQWDW5qP4YDdiU9gXMQl0+xNB5rk5fYBCST1UE3GdtIYn5DgUiMCHoi7LhzWpnK/
2lwQDbydmSwGV8gQvuTYwW4RNFqprX4FGhCGTKbxBLOtSvo30nzF8ullGKJAaFye
ZCczrFAKrSHHrQGvwt2iwHNjzmFt1jG2XyqYoUWiLmAJFa8MlygmdzU2Aomfrddo
f83RnzZI41urJFEfZWiTeA/Xe6DZNI2iHo/6I/KuqRvUfiqgSm56kjD4Ozw23VPO
hLH3J9Eu2AF4LQve4hD00+iVUKYX1IjXMCOzAjcdy85wIa1eVrA4aWkguFSigegD
cM3zgSyDBQJQ9nIPnxEQTTwnizrSXWB731pMOAAXp91iLp/j1wo5NPQUagxfSch3
fybb15dpQlR9P/pD6ebW8frBtAlbtIvjG4EchhJuMSvcpCEOLPHq+axlSQjjQaoI
HTiaLtIth2k6PpvSdELqn07EK/USTACQKA/LypmiyDEO+IODNjPIJ9q2bzbU1ADm
uOiqvKmzJ9UdW+SnomdNBeA/gao+xJ06rMbxU2AS1jS9Cqm8iDAh/An0d+ixNJ7y
2wMWeQiH+7oStA78TXce9KE1qCjn6IaxJEUpY/obSCQ5Z+DUV7eXEoT3TzIT8KBk
MLfDmDUx4T5vVA36inP5HQUUcxlw8yxsPMBA4yDoxMgl87/028vouuA1vCOefv/T
JtCfF7+w2qDUhEdRPJ4BfpUtjcJx1WA2uzN0Ig5/prHtzu5sMfDzUyIU0/j1TtUO
+bDo+2bWY82zqubm1s6xyDTGMjDJzsFtF3aMVp4PryXy45kR5picbQv2MIQLk2Di
6EATn/0YuZYi2+ThuES5Sz1TnVYYjBpao/YD0w8IpYq8L4EbM7IrRdx2+1aKGewy
PkvKT9r9KKBcMoKEyMkTWvYE9LoRnoZy9kMvxbIkLb3dWY68zXh/ByF9/oMQSbcT
6jkW3AW5+Q0Aw3WNYCVq3pgZ6xMHa3fMvfRG/kEkW1qCqQLw3HRNEXNMLI5i9UCo
xrfSXhOWOlhKTgvtHirQx7Gt2iASVlBqtcrcS4G3WRPareOidP81cMcocRVmLaj/
pzlNz+zHsXMbLunS9AU/TDexGrMOS8+Gq+ZoY5tpwhqqJoUGm9jNllbcWfBgymuM
a6lx8dSB6FPj8E0Vw6+elhqQNZyfGw6kK/9dTyc0blFUfQe3HaKSMK+fiIN6uVjV
F/mNXDd7Wafr3e+vlDxKRU/FC0KVJi0aNJxDiEHCVDpFWaCyWl/yBj+Dl58j/6pz
LC6QvDo7NP9Qc9sZaa//ngM7IiYPBarRGaid++zCnld48xzqPv2+ykHjLIHZ0jT2
8Ng/z14pmfAcW1uXx6KO/slHE76cnzu4osXcPPTfII7gkHxe+zhkxnJ0UpudLZ/U
njZd4x9cDZQomdXwmoPLgJr4qmDIEe60cZzBZ9uoowbnn4WgXEY8eaLE31g08Iuo
XHImCOjZk+EPu/x+z5NTEqjr10XUL6XVXyABmNj0xKc0+euU3gNJGl2e7tTH6d0i
9E/rfW9TwmLTw1es9DZNGc1CUAeItYykjrrFwYgxFryv0SwGZR66i32vWgMdF4t/
FLahfeBzZQeGUq3PzGePBc8Kn06ue9Rh6riQgUAjtZ1VmchhdWDv6r1XBmVU++wP
6tFLkCu+BSq6bYvcg6p68MiKboEyk2vSO2LTle6sV6KjPJqONwIwbHBQsnxExkuA
4mvFe2MQeW8PW8SLKIJZ+pWrycX/GHeXepKkxPDV7Dtsa3dZ3MEYDPGHN7uJhPu/
d0OTzxA86cO87TXYzZvH7Aslxyy7rgIgFYYmH6PtMk25jQi6ktgV3IYjkvAhSlsB
NXJV0sVRk94IKhAKlZU6R3PxoZrM4SoGYzVzCn7GXVoSXGrlpEnT7i4j+EBNa9oc
QyxZS/mWFpWoSBN5F/Qoj1/WkbJNpTg+qI2dwRhg6LcqcJKAZHD4VumIxEobPHyX
Cmnb79AN0UcJaLxE/AcMSypTt7YHnHk0BZgrhQx3xfdm+Dyn2nPeh99UoYuZi1jq
ytF2yvlq0IeWURVCK9RHag70ylh8wQadsDF/MB+xiLJ6JStmcUJslRVjpRtLiAPv
E5JkWYr0xefNddZq95Uk5NyuuQfyNFuTHqlD1F1st1ArSlmlRHvYDKPTHPif/TKx
SiYxyHOIRM9y9e4QF+LOESC7pg9F2AmMDJq9it+0sbnxOm8yQelcX+TUAASP8kcm
igmluyqRGYErThCV/meEpsZz12947sJOIgUvmwUoHMAG0XkWLXLgf+phLof5jxdo
BuXoFC9u0B0INkbw64zfRvUJ0ZjZYCUCDDXnlhZcZqxl2givpnvrPFVUaoO8OgLl
g3JswFvXMrQ/h9lqePGn1fc4cMSAQcSUJ9SXWLU/AYLQCkAgimVqYYm2Qbnzxc8S
aWAmnsInwQwBtck3H8V+lUOvzeNM5SJqiAkBkigVEWC82YGDnKTpmWNEPcSgm1pF
5tuE9BdTCfkOSFJI6ebC/JDJIhb4blmHES6b2GStiwW+sWp27V83NU1mPwh7cwIE
HrDa0uYU9SiXiurf7TYbVhFzO03FHf5ZIuk0TkOh2hMuxjE/MUwCNEE6pFUzTJPK
pdOzYM11pEluihG30VC/tDrZwU4ddp6MMTa5xau6YHpEexhnp5XO1pvyJosBTBGI
irxOmiCk/1Pw+PF75juMwETB9uDQbaU2YF0BkUwLyvapNAAomfUy6lO8N2eHx8qu
FmbZXfLHpgvrjpY8yrSdPL8Np9/VN8GpVTKXKobLqwcVwFBSIutLBLoTPFcvv29g
MPVXbfFqls5xi2Iqf6T3AH6xo2OP+XK9cpYGVcIsSudvTu9yxb2rC+Lz7knpJVRl
+NncTuTRp1Uaoe1caL6ARUTN7/Jx0pHJDAcDezzzh9ih4rtxQzwQ1/hci25T/3QN
gMLBn3LXqwLnVesjx+ZBuvUwu3gTesjX2JqISQXK4VjOCNsPlwV9z0BHAHpT9pNT
wiCesyhTSkxEvsOJMVE6mxfsAdCF9kpXY5Ig3Xbas2JNm2UQJ+2EiAvskTDnYtd8
SwpeOSLPITxs06JNYjDvBbAXuaO8/cK33IfyDGDIfztoN1EANef9rLaQPxYmiu1I
6U+4VPMlUur1MUQUz3Z/fn3RiIJvQKjsxEx1uHL/mdT5RB1f6734rmBXf2vLe6To
NBWqSk4vLSEgEWlvSEfAZH9hsnoJaiCTbxdK6jT28cOHPMJnGgBfEYgN8Lo+lWNP
URUx02+bKCnmxqCOV6EuBn72PN12Y/FXOZlbKN0aTlMeBPt+v49QEAU4y1hY/VsK
dXIG7zZZKb0sKJrWmzHP8cGzjLkseC2wdWOBlnPBj3bNswz9waLdHqktOjW52ppt
bD0T4d9kCuRdrC4//fivB14i6zXlX9QQ0zX/ImYRIvlTiLRxomzaSThAG41aUjXR
EcUeGB9pvl9WFB9dT2XbYNqZlcvb2vKVcRYHAsKqaSR4CxPKeIQlhK3g3//DQ1/E
W29BoN1Co0yD6ae1Wb+avnLCWmCilR85PdFLKPoGd7EfR2aeBX53nWBVNT37rxpu
OUNKd0DosUIztX6FREYZiDN889QavPVjh+t5MeqAazUO/cyGN6Bf1WLM9kARE7MD
ntUSwitv0kB2tez/ZAiFawK99vvJIWL3grPkCq1O3sr1Ox6w8JiOyx04HaIR4quz
mWT/4+q30OD3bbSzzGCyh8z+Kbnq0fBtQhUQto4YEig2ptlmrEWgebaPw96Peaa2
1uTg6GOq3FaXNLHexfhCHPLX3MfgfX5ifsj7wxgWMx7K64LmhxejBz6Z8r6WwO/b
xTWQzYkVMl4IS5XJKYGGXtmEowRaOP/K0+a3fW+rbwYPg4W3EiVgULP6isQmZUPq
V6VDX54ePFIDJWEJhwzK/wjB2yQwdzGIvm9FygT/mkUyFBke+5akmT4rRMWI1xZE
X+7EWwpLdv2WMc1U2dcmguiZKXidSpIu1X14VZ2f4OEtfPUZg34/4TczPO+7Vq6I
Lp3IuDzffGve/LFaA/y038EDu8/A4ZN3FuYeYR85jCD6JWVJ80KmKipjOP9CMEbu
7cfZCh8b7wiqy3cEMiJzjXascdFHrGXQLsVBYBDW3vtIfg89bMjRWDkjzjpRLIvg
83KqgJnhNlNPtk+uKxvJo1uzkhN8RmfSQ6Yeq/wNLXRWNs7bu2dwtDUgSQ/aIMZE
GECQifefTcZ727cn3sN/NE6xG85sIkOatNddY2Q+wIlwME27UE0vJeypCpM6EPq4
8pLNWBGLqOvnCSl/T1wWDs43YQBo7uhfqL14zDkvt3CxGkyAfyCn4L4dc5JRG3wW
UujQtplo/ai4HOQPo8GM1KvJUo/iXqiszcbbVjX+dAOSKEYm1ReyjbJ+Jd9lMqX7
5pP8g6wiWamIqV7ToCzpw1GSveQy99cyO2BJWF/qKot5nitGUeyYyy9xBGdl8wVA
3trrjQoI8wvBweDqBhkkfrgBH/BUYI1FxOEJkQ0NE+L2QUe1OEy8HqG2O7wK3RD2
eyf7UkH1nSGzJnUjJGiHzKM0un478p0clEIknaHaOgByOK6zBU2pnlkW9BHzfvzv
vRleMrnSGgowWcjSZStAZ3FcqO6+p8UN+SKUz2KvnJJ6wnG+x0pt1fnHe37HVTYa
7aULS40oqqdOy+BZbPtB4ZQC8zvW+bikhxYkveKLKv8zzYj7I8nUz/S2MW5j0TpL
2oJcW+yMSvz13PdlO7fQsQunDKyYUVVW0BinPu59qmoj7zs45W5IpDBj4IixMKN0
ZMQIblDAVJahvMilwoRjqXO8lPOW6sgBYdOFkcD0WbF59ff2wZrO3qwLlZ3gwtuE
mhh2arCJp/fFWzd+swedUajqxeSKl+PYW2LeAbfB2gcaJG6A/OjuU11XtgZt43Y1
oB+ShusDI2kyqFv6sL2W9hs5bocBvu8rj1E2d+QbO4Ht+Vieen+u0/56UzYRx9K1
ApNU4ADEl8+eHVxTAiElO/gbmqLe9kStnxbJL2A5p37H9co17HbReHlg81lov7BM
/LlRh0XM8kDKJr2p40n/vqmjkL+i3t6xImlOFqU0yGu+WZ0l+0TUtuKA5v/H6vxd
SyZrq6TU7ZxnJ6I0Bg07rBlf9qSogyyhDqllef2Bf/qZvEFrXc9qTJo62aBSiC5N
mJNs/IEs7mkDtRAlcWYFD21ntkoXMJQtSuUpUkqp5977hIYQPo0RfIrLm+3djcqI
SrDDLlEW3osiJuBR9UGIOpBtnNBpzTE9fr1jq5uJwLAFhru438VzaWYTEGP7El1I
RQ6ga1/XBpovzlZ1XPI3uVM05oTI2zkJ8Y9xicMMf89Z3RjmIqUAoBqyOs+X2PWS
WF8FBc6drAgC6g85+hPfKYwUuSxq5ScQsx/ChCF7kVBEmXVJ56Mn48pU0xKf0uPg
aLVeggJXGUWs1pBqvDPLacu1BrN2kPYO/aSW3kAlKEbG+ZLC+7iLZRUbxI+C9bXK
xZjN/mkdq6E4nIj8kcfKfm1A9WwqWL79XwCrJV5KvRgj1aTB87Bzio8mp1D+Zs7v
Qq4UOBc2txh09Tap8p5B+mz8/kmk1wzZoxyexNLNmbrhBuh39yPvcheL55rTEv4+
khYJpJzVQXJtXsXbcAtx94BEB37uQsGStYFwBmeRW473iTAt9WnxYHYYmfnU9IV3
llnRF0xXaCZELFVxoZ6zlDU9bcHw7FSc54yZJCTfvKQOMuXtW4az7DNmvRYVX2jw
3ZONBlPQ2L8U8j/nAHUNDb/uVF1+S1xjjqIVCisxFA7g4GnZCdYrTuc+W1YItNup
DveoayJL1/sFTxVaXfMcVutrhXfm3nTARmZdp9PueVzgzxQq6LmRC/OGvD08DN7e
HVr3K3ZAPFH8z68aZPXfQ+0O7ULfqSBcl++a6hxUNcQ3+m8O3YWSVnlK6hc2hBQn
k0LHtBwoq+fEdm7NAijx86EIAaGwuKl0mrtopxHfG6hZB84B+4QboLFIp3a0+3q2
/eCufPp9PA2voqjGzfyTUqEIZ6D5XD/2k8tGg+rOy7cQG7Eocvw3X3PCzsIjls8J
wXTjL6af1KWNIck3dqG4b8WfS9x1leDes05CMw738iFI2DeuZiJA8ypbTVgLPi6C
yi4KMBhTz5sqjj5H1TAtiIQbrcieg4Kvk8yGDO+YKw9BSeJtM3V/iFr3hvaZousn
q86v08EwWMZOSn7gAzBJJ/Wb2nzDCChPqNC3OKT+OyS0XGz8SqExvHXl7bzTDLgs
PpkWsCNoGRblsnFsxTvEw6UN0ND+C5St3GivX84fDB5Toq7kJpgONXUVsTBw/bnl
XcpeXzLpu2bjRV9aCtnc5pEZADRi7st6+W4TifK2yVF/n8IC7o+vnIn16wHNEZNw
ML4sbbXnFCCnd80ovSmYbR3nf7/1DR0yZFnkOky4eAokn0jJJIGYm358HDhPwmbP
Xlp+jAF/YKItSrg4R5019K4wZwkDIjHW76AwgF5QAVNXMIiZvow1PI77PPK4hZYm
OWWIQlv9+PljZsq+olCq9L3XnFAWzIwG7BS1COeZJTGH/HjZM5ObpHON3DoMQLrw
r0CviV80Ccw7UX0s6fz3iLLG35npsEvVqLV24++VrSy+iN9bIpwkJByng5RgLkQY
9U1BsjC30PAUFAptAXTrWd4EPcYFFP9sGhk/EruxPY/AipDdJ+2XJFHmuToo1Vsh
C6rfpIbeRhLM+BFTLvqW7BwfdNa8uZxnkqt6XtSJpofQth5e8TYLz1HY6LglZ27S
D7/MQpHEo1aDmvV1e/plAH86KIhuPfMAITpEMirj0daesyAaU/pzVzkkpevNVM4V
81kKxQBDS9WD/7iLHqLzClxcYtPMwOS8OC4WoWJIVZ77TesT2X4qr3fUOG2C25Uu
DJloHO64G8+IRK/ir/xj2sI5Vk+NpKPuLwwxwH4pqu0g5x3rSpZxMY7zAB510BdK
iG2EqNTgj+w1lrjLpxNAtgy1EUBNoS+pkS84l6vH6XK5B/TSfre9xpQE4dTU9q0M
AR4zEaYPlc4hTmKAV5/i/rvbF/HMwBZd6EVBU1nOf/TftRmgkMX/xeWoPHlSpqa5
Dqt9IddHCOIEn36ga6n2FXX5rKP9IDdDvA3/X6KPGl+3CJg1bSbCOWmDMAQJ19w7
qOjUrdgCxn7q3YJiY8FIvTYFENDPvSKWx0Vlw6dyrn6fDq1fQUpwWWOGdmUdS7pR
/6uY6zoLbrDQUqBXzhTlxSbOX2N61Z7CzId6slF8Y7ZZ4YM5GdYr0tlN/5tsH68s
YZo7hE7EbYy+S3Rx9JHwCFr+G1KR+2lwIHtweXu+F2m4Vtm1M2av6AMYijAMfA1m
fJ2TxM9PVarBOAFwMawcY24kucKgbQzIXNWKem2PvBLXbLVvsYjk1Okk6sF4v/km
qfADLdNK3be+RRlcCzPRnS5pwhLppK3oiqFHWBG3V26N87uPjJYlOxG9nC9LNw+k
Ds8lsn8GKBQJoEeY49ari3REhgWxdHUqLX9eaUjR53je3TS7B/zTq3Ryl311SACb
fWcvtc0KI/fRl/Q0Qw7Mc1IMX1lxe1Ag7KreUUfDnb3hpKY+IjqXOrTvtlfiv/jq
v9xd6wTwap74t4g/9AAoqBkl+LrywgizMacr6loGGREBZahHtwHpL21p5CHCpklB
4qgr0+6LfLDOXox+hZbN/vNNFiKRkuDjmgVqjKi/BLZQCok2VTTCCbEpGt8ZFqhu
HkCtdRaqWuIqZ6Iyc1wLwa1XKPRshBDHV24HcilOmX8oRe4BxxytOIX36qcIaYDt
mFFlWhzJcLiym6udpo5HTrVGLoTU4tUVDaY4GiKODw4IHTuE+g4I7ij0LNTwFFzr
e8Z48ZqdoROAad3xEYOQt+bXGmknjIJrBkvBJSLI4W/jO8sdwZhS7G8GUQhW8k2c
8WwqX1BvXDARQyG8Pk/47tjRXbtOo1AOXBwN/drX8a6dCLSKV7S2FNFWgC/9NV0Z
pr4cRRaUmRRNbn4A30CEu1WWBrznvJ2B3DUR+p4f3ctkl6RitOF/VT5T3SrTceb3
XoVlIjzNdUInPLx6Mv2vvQhxUsPYmqdqCzol69dbDBX0vnXqwioJsIU9tx8O5cs9
0VH9GeM+MXlJ4rHd5qijqf+yuA6onX8AU3KegHHe99VyDRKIwjrPs1Ivo1t8jkkO
zLElPptXumaV6+dbn5iHGGEwJo3VeChPUUfyB9AAvaNio0fHsmMafk58xNK0oc1Q
2lhFxPFrsqy4EqnNbCnknVNNpk2b8MWf2qIK26s+vtn91FKBQ/sYKzDbiXh0yuna
Z1jIQ7nmUagKLSzCWJuTau6hNgO8EEY7dGORy7u0A5Nh1xIWa7dHYNuoEBI+khIk
HAbzz7wb9Vc3/YeI7kXb5fwEylZWGrlAWSWBZsDxExd8kT5oqwdpbDonFZM1m5FV
zkZFp98ZuWC99oC9sckS4TSUwL5nYe9hnI0LNJGDrrj/HO+26GUbEpIVBGPPL1tH
+gV4Zgq/Uly7WMYrQUrbml3Z4tlrH+l6LxoFUA9S25Zz42DuatUDuQEC+G7AdgN+
2Y59MnGEEMsNCRh+T3d1Fr8krjao150d+6gOed7xm7WScucJWV9jeZav6bmDvQSg
11ASyjAEYVV5cCORwKJLLzjtHdG7hlHDJLsVDYmp25OHdUfOpIC8O/0R49w4B7Pl
ATXzMY+NhntVMGs/FSuLQwHX+JbpfLuKfycSCmm6pSWcXu/i9aUkN6i25BY4RIiG
HC5+voYSvc+eTwJqou31S/XLNkk+nx31UFNtoQhE3vxWnigXKxI8MqGbg9RS2goP
Nf9QxBVXS1UO/D1sBHSH8s88iwVMSKuXxyVTUmkkI3vjuyeufLodgPUYpwsInrwd
1J52NmFSJZUrEXePXApvkkXAomtyBCLmD3gFb9AxGhL3WHh50VK4vDauyYZz2HAk
g7md64GdVQ+tb8uJLfY2/rSQ6mX80azj0PYQ+k6Ihmo5uGaFSTFumYS89HCLeQI0
u8fMNQ5QjWq3OCFo3suvzUmokJjUMtSHhoTyyZG4qipuYm6akPYvjOijRpq6hR+D
uvvsxAi0KEfOco3eUmbDSxMq1sMO7lGBomGp0uWivjHvGOTVh8ApJ6YwJISX48oW
jCUKmO9nni7rS9whZefMtjqciDfXd9YnjdR86Qd/Sa7u2OJmlq3gGA8Bocqemnls
TujuCI+aDhz4vF9o8T05Zpq9zt7AXgAkhwBgbIwHeiE3J6G7gbatRcCo70dBZfcz
sW+gqAiODMqgS1agvwJnW8fBml6M6dvdnyVzYyy6JNncucpx7X21SyP+rvRddOd1
vVR0hkhOD7bkvRVGXWYlWv+R+2riC6tfWYnJBrevsAahqR07d6wDRxwidm7N0LqE
+0pfove1Ilfr/CB5gVhoadygor4zX45mnThJLy1S7hPzMqB/o3rkrlNGRQqay/TV
S0FSD6K2PKxg5dgegK1Ot9N/mT6lAsrdhp+6hm4Xazd/LsjkbNgLUYm+0KUSjwYM
BYLAecc+srbQ9aAJNddGuIxPMTttc9Tl8Qf2vziOAekeq+dGi2WD+w5Zd7bLRPP6
/wc/4QLP1cEBQeiSth9eOCPJxxxGmkQuKCrnCy5UsMKfohL3RwyHuv2uyWuC+3Qn
rAeDXy8TVTMIUk+NB8oDT/L/sofHs4u/JQWCCLiFqu9cLeGXUe7mlKxF4DN995+Z
wwvY44/Mt0ErfrtqZyNk5L0l9rAPahccWwpQ0DCCrGmqxZ5NbOKni685VTnCG+zh
A23/g8I9hwPkftRGHLbRQUa0FGxSktiCfOWB3hIDvJgX5DJdd/Qhq7vb94RCOl75
MpeOOXnv16nsZbyYxsPxRVVdpODRYljfQRq8hGlswWFwqjOaeCGyjVHc1dIZiqHX
MaK/sLbM8XzJvw1ODJgpn+SXjibI3+rxiM4QDEwIbMvpvGK+GNWmvK99g1ZCpRNb
adJ1AcH3fyMTr7kJm5VNr0ZbBoigKjP2VMIUSOgvMahNrcO02xQBmosAaja2B7DO
ogTCFcdS7dSjAYqHF23GvQ3n6ust2dR/3QjZ3vHSyDGyH9zzTY3eB2gbcPVgKoP/
/RJUX1Bte10Vod7IQFP7vZUShz1yjpoICZ85hJtPFCz1lReUYr+jfOzSNA5DB9pk
NMnxviHvWpPHQxF0pu55Hxeoa01rNbEtapOYwXJh1C+6YPrtmYBEVFlDrv4sk9hm
g0M+q7Z9O1t/cn+Nb+gAeVBKbH8YG7u3ibzM12zqhm7cznYEY7OCKsj/KIvs58cL
Iw8RYGt115TvuU5l+ZSdCPQ68J9I+gTwHMeL0I3QtA6HDm7aZxPEl4+pXm+H3zTY
2iU5qzJ+L9uuGX/2e4Sftd+heKroCgtA7nSRYUukmfFrztVeYOptOETMEyaA+uBe
zJNQNXq42bkXKRq6ELRxuK8uNjQPmd5Uw9jvVTl4ZdjN84g9ElW0VrBDdeVnGoky
CauiT0rty6fmMoTODlnAevSNtOGDzWJ3DCcCFSGYUeR0p20Zx6fEcDzhS86j/nND
QIDwaeKWlXK2lk92PSVZ5TmxanQmIddCnyQ2uub/axHthzBDOfEuTlsVkXyngNZB
EQtR3Sv62JqYnIdcaqhpa1/dKohkxCOOubORMOd7aY6dKdD3ZRAjMEPqIQ/5BnXT
y/eJ5BNrdGhvTwM/xTV3+nM4UzIJKYP4U/WnBrEKnC+NIpVUUYwNRvtUgkyQ7fSF
TNdgRULylrUU9gbwP3J/iuYiXRs9a2qNNlkvaJpqjsnvHqYjDNGRR2oqH+k4791r
clJyQOwmRVgyKHx3IfAjuwVaRO6zQ4vxwkTh2Y427m5KfvMOpgPhHxR3TDYsN99Y
cfbsy3UJEzu7RmceLDgj0xAYDXWPxW3vC22Cx0CsMHT6zImwRs+sPsg3cSyfvoO7
xVwLIvCUQiUXAAzsvrrglNGVfn/MlabMKXDUmP4ilvogf13jz7yvNaMkf/UbMdkA
nLZu7diVhrRA1q8/IOrGjtUK3taIon1JOPcCCAiRweWx1ZxAqfN98QNSJz/S29qJ
pYaor6FmG3hjaQ/1XtybhWJrFgzUETAJJWtVVeu2k2UoTGAG+Ub+EHOE4VGq0uto
bi3n0mx9B6MTDvQ5xUF6UmXtCSMGbonFdPQ8nN/yDkPHldBGNzow8NfdxslTi965
el5UvgIFWe7F+2SogWeyAV12LIQQ/g0SlbD6mYY4e0LqRzTk8/+lRKUplKg8g4FE
1+MixwZtd4q49LOt/Xfhj4btoc9aF3h5oZ2pZXAZ7HWLBwf4cL1QIgCAjx8zmpjB
hm6Sy2XXPzod9Wm4kYvQWTaFEcPvc5ulQDIwh2GS9CiR/DS6L96PZ9uwKFgMAx8e
3XusQR2oBNQ24AMsQCP4ovYWp8l3b9H39wJl9L7nShl6FW4NI1WmORLo7dyHaGu+
nsFpe+sy/TyhHNEzNcReaqDQoQOQtclm6hhVNK6qAuLE2Ok3D+vrI6YwJocIWPS1
WmpY9IVYyphIKEKzHTy2GOw4Wk5z+JPfTgrZch6V6i3W25L3jjTDSGwtqacQyxGr
xtmYkxfpAtyizvDmOaxTV4Czp6cRVdR0F+Sy/prq/10MfbbM6nCxGgUItflEUQda
3MDns0tTZFRfgar3z6NilHzIx6A+zlsyI56bIjUpvzl/zdgYfEL4cuIj7FyPhr+W
U3KxtuqhpHfp9nsx9Pcvv15qWcbgYA32hwn8pvtLMl0wdAxwWSs/C2Ma0dXJEg7x
dNH9uUdhhO7TFZdc1Ilu9N5JLph+5hct3AMQo+QPVg/6+BP411HNfm/7ShgFsl5F
XASN5fc4WnpCzDdyNVL/sF7gKhAkd2Oz5ep5J44hvCrHtvukVsVGy3uF/QGoaXvA
3UdbnnuqhNoWreoNg8SG3kZt5r9iBnFph+C70kj0bRNI+qygMfI/9XjUcaIFaVJm
46pNdDtxTquf0+YeJJ2kh39DYZ2I3BCmJdI38sF//YgIrm8wuUJGWQXrx9EIBrT2
GldPF8kvCzK8WeigszssPgqoJFrpEwMeFHtrAm5ko4CPg2qMryiSBAsc7NZW4YKY
fZrLbpMwMEjsNYGNSIJCte+Kwd8q31UlEajRJ4LnG+RsGxfLqcdJYCw6W6qhWour
fcNXn2vN0rZGNSsmr4ev4FAuZKe++0GhxTV3Z8ojtwXEInOcBxHwDd7HFqXgeyrj
oFazo+1P3mAk9htUY5GL9aG9fLPZLlMXUy/0hYbxy4kHwl0po1p8ofTrBU86I9Vf
tsZMuIK9AWKxU/wO9dqiDHHcb1jwrN0oAAZsz9QTp9jq4CEbg9wQmnb2mRzCxUxC
xxHtDUdYw22UhMQtpJIzvgyUWLAhX1nQVT43O1NbnRHHgGbxQUI5+OnROhLijXzA
Pb5vxJdxx/tCsFh2SldfREp61THrp0TWLrklBOqweIyu+fiFfhSSzswNJMmWnOVT
5RkY00r3FNgbyxnBMtLhuDIOKlD014RdpMUH0Q6kO1EZ8HVuxUd0LecMeDveRHI8
imYJtWnP/sMDoX9G9EcEkDKBurqXVHtQOktSi0OHEC1WHc7uauRMpcJf12b7qied
ohidn6I+wTjwfAqLuEh8g+3qC/Xfc3xlWO9i2yRUhuRDmJeaWz/ru89ics4EYoMq
PV2EAi6XuiAaYHvrPV0CDJVNEBCLurYbJzMSeoAsxzOffuO31FK1zgZ2blvQS7RG
8GKEXU+ALM4T3iPfxyvBUTFMwXpbXRQHiKxzDzuVBpj7q1siH/4EeTZFgkTNh31Y
84Z4ZIiLy6uyFT0uqbhUQ29XkjSykUBwybOHh8ZBBYBzptaPjF7EXn9vBFDgCxJC
XmeBoxG0ZHXiv4zLw5qeeuWIpy8ekR2oyQtxNjRix0osM7ddeHYY4c2xz6GHd4W7
B1n0sHfMp8+fOCuWtuay3moaTeP2J3/zeN95H9CkOilBLa9DDJR10ZgUwlGQ8gO0
mxtBjGN29eFmFbKP9N0kS/5aN4YACUPjQFGT4cyZsfSGaYZeBbOHetmryIdeEqRz
Xo4RJmmzKF8Rd+LGCjElbV/L2s/dQti4Y3Wmu9+luilRrl3WOIXX62yob1sY4pFN
0+IWcD+rOtdjWKuoXN7FhUuW94IPBmh09eZD9FQOhZAjzHe6ofzIRpZE2BaAMTq1
8Ft0XRR8tdLXCiheZ8CTj787gskh08fBuQN+LnKyhTtvDAInMFTdrY7TW+Qz4Pek
QWRZ0t2l9TMTt1c7oLCd0GOe4HUJ/Mx36jF2XuJj1tZQi9+d4q+gV8l9Zqo1hdiz
I3g8tu3LG9sO/0X70uu8ndOxBlwxj1tJt+xQhffrVtVInQNJxu+TA8C7pUVoGws2
/1hkt7p9ey8QAf5+itCVu4gRARzxEUm8k2d6y+Xuw3lWXDjW/HsATIVl6gbKGJnV
YLoeZ+ecsu1iQ5iXv66Bm9ujCX9a9cvP80jz5BTvIra+qgj5tvkkZP5QtgFPuIAR
5xzCTnfXIH/tQmuS+2ZmwEjgF7bvXhvdAN7uIRDKHLjjju5/GefbMidjUEYC+Gjm
`protect end_protected