`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 17440 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhIGJnlxXbtZK6kxweF8m4XbqkTa9dUaHpRw5NleAIIft
yWLg/vY67d1dIwn2pN019NE0h1enLV7O4WHJ10MM5c6a+LeMmSJSDglf7Vt5nUs7
bRTrQYw1chH3v0cVRllm75UtCIGHWEmoHz2uWvZJHeLJ7Zuz856YVybvNJmjqB+q
9I9FBnK7z5xQaXxDLrac5teT1oLdr6KjykJTyy0dlQEl6M9OgzWzEYbKdbkLHnj3
aIPTHg494VrTx054l0X36ADGbVGx4UjyPabdpw/b66CJbhNVRPaf/eDRyH9VbZzK
XDjunHA/exmVJTKJ4VIJgZcRfju+7rqGkRH9f+gWN5Q7TI9r//H6xOgvWR+h6DSb
7Cjo7HNAXWMranS/5T5dJbWkT820WFuzaikKlRb2gEm/efNpfffSEvOIGh0X27Jh
1Y2pL6tubXjLkW2tXZ9NFVaD1O9n7kHL67/cOrp8sL/uDqrLg0ymxyDEkigu44zt
CqWlgBTknCbc0zljWN0lpnqM0Oehc3/QCk9pPB/O/5gcho2EAt8ffbzK6ApJPCxw
laIBgTcxM1FKXRzU0v+CyaZw0lprq2bvaFyjRYljW5Z9ki8qSdbMdgdsvIyJisMc
RTQgiOYHyCwCVM5LQtK/RrsgVituBm/N/OHQVug2nhQX5cJxic9A1iEgGLUD8VKv
W36I7GYsCikDGST6v8A78tKsfzc7MUnvK2O8cYJPsKA80dmQFUbEy6+CePa8Vdt5
FSAdGzYt4pb/VoyfJzcp6JxocAFZJCQc8VyaDYNbAlFZt9m1dEdFvSqT+VgOITHG
ovZHgcqFp/3cqUZL1g6YPb3e6srw8gqCbwUB3tR8QUkWFAuw+P8vIcOB0lSSoeUd
Ua6yBiimjZyz+8ztW4F8N/qaZwZTTaFG9RqSYXBKRUnzsSs7teGSaaE1SzCuTEEJ
DV2vrtAiOAGh05aQufOYmCjZetWZV4cVilOzmoRnK+N9Mp/mLZU48FdayrXWwEaU
UObnhRmO3XxbyOXLWkge0yWgYq51O/KBYA4RoK51A6AaKHngHFG1QYN+GID9IN0j
P9sQNLl2QzzvDCuDKEAxOaOIzBJgiWNz7YzxdfRp9nBHRLdgSCXqzF+dbCcCcKyY
FC7JlbhYGXcFqAZM74ZGl/HGGepYbp84xAejvyZa5CSZ/woTEXyNUmD/w/aUwJCl
cb1e/uMLTSjrmeHD8bLbBgRAVwrkIaa7aGMxtLOq61hPQqPREyCA5JSvMlp4xh2Y
N12ZB5+BZt3HoqvRtWL8wIMT3rYl34L5gVNFmfNeWk5hX6+xCJFp72QnIKflgQMp
+zRDi/7JcmR0AeCyhfRLmZ/O91JJ3xR1kVhRq8D8/C5T8KDmnJc0k6dG5SGheC4b
RmHbOyc7/8rHqwCBx7xlpFteQxplpvLY8NCspUimQw8d1T4yB8D46DiZdYYt9vyI
9pT8jg3O11+EHWlDGa9/fWloWA5KdzbESIZbJlL3v29MvoIQIAILU3z74+gQr+9Q
NiXUaA7tynb/OjaPuW/3Cx9NXPmZP9R1/lmjBB5YTIo4xcDgDD8Vg9RCd2uMInfM
D6mMlrIeYrnQEVwpTqXIb00bD7GyaXYKfWryqwW3VUBYgchyrUWIKyavgUzTOfz9
JcVpeGX6sDDMtcILA7rGyrJ5tkjStMaoRa+zFM5tkRQBoRIgDFSw1pdK6XDMhPDY
+A5AlIh5PHMpAZhrSTDYY9O5vhQBFuOO7nOTAFg9YZn1PEEnzyYj9bXDTW6GzLgr
SgTgqQlHFHW6iPe6izWwHDIb7JNoejdudpiKdo06FZdgRfwR8xRIXZx7tsZ3Q15O
mkE0IUlGdfDwuKRyJCgS8Xv0547ehLJuUIS7zX7q9FuK9gMBnjCTXEB/Xau64NUl
bGtau88BS2s0H5jMgmyb7bD0iQjFEGVlC0BCGUmJ1QQ77NwUeLAREQL6LE7bVORE
CheMYT0ucqZ7hUGFWxP/Gpnw+heb9FSeqU/hmsDekLhQl85UaSZx61kMxUwChKj8
J8I7Wo+XzVKl0G33GhSYWCBbFXKXilvuSGvu2sPYSgiYv30fNECihjDYrQVJUbZN
5nAUNTJQWni/bVSvzmOJ/uKruudA7CY1LNr0QxkaQ+ocXN9DI04jeRSL1T4ZAt6s
+5AOR+TOELG8nVGpIrBiQrlleyA6YZiUyBkz4L7huiP8NgtfsbJLMfHiMulauZLF
+vgrbyQkXymPnUTz4c4RNnZiGggjxZj6IF01H/XqPu78w/mlmiDYzqiBmu2CREt3
KsGbu3KArY4F9TAo6UuVq6CV2Sq8OzPmnha8xfiaWgv7JGQ2/4HIUyr/6SYzrwvV
zaB5oy7plwPWrV6gIp/lQl4LXLewE7LqCXQUy6cvp53+ZWQwqV/jvroJmjak/fbx
IPOOjf+QpMDHvwHsqJCUNfk2VTtcDMUGOVH46R+CfLEFJfrDTQHfwjgAAAhYEskK
ToyYKKuiU2VDATdVtBbAV1UHgqyRkXqeAAYJQG57ObTQttqInUCYFplyoCBDxAtP
j1oJm+l1+7MD+YIKjSQXpRWpbKTNGl3qSTLw8sWVE1DjrBl5gLkcBPH6nG0Ocvb4
B8HAaeZbe3Cfh8AedfiQZlkWACx4xfEhodbeommCpfJV5T34gm/eoHYkqT49Wekv
s1u+K9y96LP68m2HGFInnoRJoYeAZqZMzLq/htm2E+2Bga9IIrLk5StdNi7LnpnN
A1yOklUYJRSP5d7kkbY2lPGv+C5R3rN2/wlU4Q1Ll0gli7HohWjQEZh28zd/dqae
hnbMjeodBpAqafZLc4W2tTIMKNYIz4dbKddLUaDN0Kjn0vbzS2PMKhpC+wrdouxL
uzXajyK0rq79JEwP3jhvz34zmy9yJeT36mDP51aj2ftFK5U9G1Vgd0X657aq2TEM
DGjMgbIqTU4z2MH/gNn/5ssPII4BSpalq1vovc5Pox8FYgNhZDdnJvndhhAEauXF
TOOlIAu/1FRqbRke46xCgnoGAWIhjhOZ+XFIoBDOsBeGHRz8WYnlwQDosWoKSGc9
zXCCGQ9CEEaimNakNuOPu8fpoURgDx+r7BrQcqlrtZP3oCClWPJ5j6aKr49KYEsr
lJFomphy8Q9R9IDSB7VcwLvhdUInj33IrMg8V/EXRYYTiTOGQXmd63B2gdz47sOR
W7rvf67ADDswa5DqOxAmjVaw87YKqiRmiiW5P7FcgVitmiO809shDpyen+oc5Q1n
qMat5NuIAJv1hVxQtWTKmk83h42OXR6YjxAvjnxsxDyOThZR1Pc6zkt4ly7DjtfL
s6IZLL911rQXAu4pR9mSmGO6FFsQCoGSn/iRMuMBYJBeiQYCaat28PxSWXfy5rL4
l0zIH8WP7e8O39E7ud0qgYDD5jNpRXFzKpmO2C9VOp+J5rWlIBeOLrgblIwAtrSL
V9R8/w6OBYzkVctYPlcURcZLVCCj0ah+OZlTkIzFptDy8DZg27/1m6P4o7O48H6p
gbo/wMsx3r+lMCm6kW9x55QJT9SYGwho1AABeu46UGSNwRCcnW30btksiRFDQ3dh
NvZVx4zHVR6NVnQ2bdpXvALFhy+5gfy8JFkb9Ga1HbGAlVskQ/oZHg6xO9QJBsYu
cksi+KoCbK6/X5SwIadbJark+kEJwWbiRTyQIN5hJ51/Y4ZrAuc1MarVPhE0u0Xs
V845pAvj12ccLbrupAgAFclB9oR06ZZ5WxC3BvG2Y8B/tc2HmQDjm3SqAkrsfehn
/CaJooJ/KOs5aFRNviMAcFKZtwlsL+kJ3QQ2ei3V5/oqg1P5lXHWI9RB6dNO+vNM
T8bbAMtTJ59oKIp8mj2yGEWEkHbJsJeK0/bjpVkYNj4nvyz8UyiJi4CAGT2BVbT8
NxsrAX5KAjJ4RBgMg8ymgTXjGfPSU5aYqxCbFLH4KpLeKc5YhNfcZpzfclWvTjy4
aa1b/7D3tY0PIcJ+7rGwzOIw1XgNoZzZirkiPOoALxeZGUkiHJHNvbSY+p1syIh1
v902O/4xdiFdF4AuJ5n9Z4WIvIZCMbLPO9ZLVUzOK9XzW2pSUvfQPyqkt7jTqcKu
iR07BrPvRZpJtPBU0yZSCi5vEeMl1lY0Rd1jrl8ptwqTI4sq3fn+u6s3hPXaWygH
auq96s/qmCfrJFVOxvFZXTSqFCHkALw96GE/XEA50tC7108LUxxanP8xkD9VywMq
dCfav/G2niaEim5FhcVMoQNwu6GgtCUSNtR3hsQYs2zzUT9EgR+g3so+35W4bqoq
7KLLMk4JOtSLKyaqu98YFwaxsEVnYxtgClePsoSuL5E/GuoSwjz2E2/JbLVMnugI
VXUDmRBf2OUo9Ib022E15lwgW/epWQ7E0Jk7bBIK+B+Y0xKO2Zqp/FuFZRCZVrrF
6GZraNwiQVWmLbwY5u690PRywpP7VwklK2B+1ntrp2CT0ppWHJUxYEiS4hMx59lP
x1jzPtX031e2NzxSS6qPg3/+gQzxd2w4+IG2hNJnxxyK7xjtWitf8uLfVkeWoJdq
15HRkL3xVakNllCtDDZoE2D98ZGvNHXwSoof8xuolRgHKq9thWHqBlwnuMLA5C7b
nEPy6JtSeRFDwVDo0SM0aILhL3S7rcZkeKwFoEuiSDaRzV1+S0rm3hY9DKZbhm7H
l2ROj3J0nUBTzu2aD+Fde/ediFo97DxCGJhUVy/B1xh9+g0uL/hstF39XjpFpOW+
VApXGRBvd/C/ORLKmrcndfbac88hdk83SlEsZNZIlBoYYE6B2gYCwb2d1Ym54xss
SbcU5/rM9dh0BhfcaLhx+xEOijjNpgGZLRGghNGHz9I/ufJeGvnPmP4/pCEpROlu
D6Z0TIsSBOB37tjvqYk+TEcdTOxe0YzhAeLmNmgSC+iZRz7+Y8WQGkfiZhLAsTDa
iGmAWA/5ductZ7EdtGnUJ1+S/jXvvv9aspmDoq2icQG+e1Wa3nXoF0nK8qcoVrlB
NLf4ZRT4RYR0O5sQeenuBuqM65WxB1YmLi6+RQUbZkasNoaumDZMJ9ywXcVg/NkR
6t17cJuTlcAusUQ4t879x14TsvJ24B7iR4FuWfqm2OcvtHlfOroTJre3UwVioP+P
k6mG6Su78Lkxa5PGepMv5Ux32ZrhLGE7cfxUmAFf2LidQ7KxZU5+AAIDlCFrSOLS
BpDJy39zOemC0rbvk1YnoyuXLnc+VnPrOeJwLgaC1nSHGnHlzJIW7vQg86aRy0zj
dClTnMoQk4DXUoSuOI79ei1MT4MTWBh8vmPv1rhTg17xS5mbLR1xhFF3xWWpi0D6
PcnQimpZrS+epGcRh9p8A5ehDdaMEe8UF7/KejpNiZYE1azhql0Z4vJA3I48DzUL
Tt/YxznWab3rns01ovNzVffcQuZwrp8oewoHnDtCmUQ5lwQ77LJmwC57GQ0JqCYn
CMUEs+1ZcOhVpILgrs1C6wyUWqfvxdMVGlspUTz0W/BWfdaACY7Eo98Zovg1f+wQ
plnIREuJGzzLwY3yDVccf4RZqGulSqEi3dRtAbG2f+MUWIxBX8MePhKe3RYQYB8Q
eWxDFcIRVKuYZnDSg9+Cbi3xI4JB/M/ZkumdRcSf6Q/WOa98jtjH9HxvURrH5D5Q
14cupi67TdWILkuYb3KwStEKCudieHnptYmOFGIDWUUODvVqiAWMt5HViYdk7KeM
2YVKeZ218ZvlqRfOZ6QGRUKKqSlBd85VTf+I1Gjn6sjcbln41VVkkfucPX3iLkXS
xDEoNsyoOlrMWw8aqQ2N2GALnTovbGnOAnse2oCjf8vL8hv3C5Qh4RRqIJh4IKKp
OTKB/GxQK4SueIwFgtS/9tjJuhyBTRi7NduM9Vr1O+Abmun5Afv3yDaszzk1a57y
7tqEQqt0kEI2kL0SFpun+sUKPoFJYwz2yOtbeEeac6oPvUPmixDVA46qdUdtRN9C
KHelznVdaoc1IALDNnS7OxmR7zDxFAjmjc80qfOZAxXXPAEq1JZO1wDONLYHXHGs
8IHhRF11UZdlygnIJA2xWDz6p5LAY+goLMOhYBZKO3AX8eUorA3GuF/8nXqD1SUd
8Z++bJf9ltFqq5v8ixeRmAsduXKMVswBOJGRxFkZ4ii9fpHlrFtlHwmLbGOjCKZc
1vdlAiRpiss/oNOqqQF5EUGGOymUB/Va83KYRdEtA0uQVcakS2OpnukeeKmF0nAU
ljjG4hVKnSLoAn7Q3iRMbMquucqJuzKhNg0gsNKKwezoVU/j3oaTgm9NNYDPHwz/
eOeSLj4QH/JiZVhM58Y1kugeVRY4IVehS7YBkJtVdkjoaFxzNxnKiu/Ce4qEjPOr
nlaV3Bh414/6cKWjXMawyuz6CGf4ds+Hw3B6sjwzp3HK3kr0FN00TnLLWj+LRAym
kY7EG6eUgdAq+Ikn+XO7sZcj/LrpesocCIEwIzf9ofCzB0WOGy5ybopH5b3oj5G9
nzeYDIP6F6wjjh3xy6mzGMd9PCO7mdO4BZzDQxieIMWw4i7SAvFPWZcDF+dTg4TG
eJG0Mb4eCz5dOoTk4YNzQp/TLQDYRRdfaEmsd9imFp7lsAdijKfZ3fl4b1RmB5cQ
kWiayrxnhm5XsOM25rbJjhFLrGv0Q6yJ7QypfFiRia6yRbkJc/aheBB9xwSg3cyc
5xORwMGtoIZBgmEAa9cEHVMopLZ7TNFTevU1GnHkJwBiL82JUJxKV0pBeqESLK7v
47EskZ9wxMvxwAgdePpaxwXU0NflXsh3mdwJMjf6sfwKQAzEfRXy+GKWyDqRu+r/
hmPiLqaCnlvetk1iWGyKXX3tGM6CasOSFd7k+zC3UJ8Qo5fcZZKdDEfvaLV/eKvO
CLTxgvlY/0Bs8Pg5k8d9u08Ah6ujn6QSLxTuwGcJBWPiK13ee7oEMuYAO7LQBs9g
6b0/vYQMlraxEuqB8qxdropYvJcaesJojv3zFT9fVKLHymuHMuzW+mKMybzv8AJT
7bLLVIVyX3XN0GBMkPPEN6AF8NoV19rOpehXLJlVtwu/vy7X+TSX0XLY1ePeDJZo
4/UxmqHMSqiFwJbbRlC4us9chT4dgD0K9vBynIuTspk1BSrvb51kFEQ/htDi2kkj
KlFrV3oGAJ0W2mtav5McS4beUe2iqAFFO0MbwN1Ta0c5DpTSM4QO/V9LiE8XTM1w
wXpC4QjglfWJjDNbS4ITBqIgcKaJVBunxyalu40zgS8NN5DYg2+JRZ0fo+ZU9tOb
wUo276Xx3z00jj995lJWqx34i6LCwAekC3lzNIn9Jl86VZIbEC09KjRhM6W4YVIN
yDmY1VL8ao7XkXYL+UhoC5yUAHQBVqcUUaLlBaky9bIK40tLkK88i8xwBX9mdSIq
qUOOFDKeFzDwuxFj98u8m+AT/X1jKDUviT+wUdGdrgXf9kaosJWQSncO9y0dqrur
A5jhEEAC+LoMDyTduTMFynqCccCtaaAI21/uucr2uvNmWLa3jMgtM1640oB2yGQt
5iP8FfigKSGYXQzwYCq6Y9HX71GZIi9XCL4Y0hbWGpAc64HtdnUKwv7BVPga/L2K
5v7p2mJytC/wMiDeEaH3g18Y0ul0qM3llEU3QZL+6L8To0nmf6JLxcFKLzz53a8e
oh8KGOGtV13WWQlrMi7KhieO67KesMPRzNz88Mww/RM7Omby71sGKXO3GYQxu5+v
5uzNmjGtYSW/GwPyBQrBggBFELIzF7r0l9AROK3b62pdZAKfKDkTj3Dpg3qBHm5u
i2qSxiwmSSlW2Y40vakI/Jcmp6KvkBphVUYnRiWOJxJcpyTUhVx/n8ia2GCJF6f9
BkHNUvwM674IbNDkbIdpoBQO/dT3hDu7woQ8tvW13pkQDYApce3WLqKsiaJ5S5Q9
zqDJaOF0SzEDPWVJTapaS2QC1nK3j2Vs1u8y2GdFTgxKKTqFzQ7QPtXP2L/0zl5i
bsg97AfvY6XyasXwIkB3GkVccZJaBIO3VS4sPdUzVNv0wMsli16V+hnbioYJIzN+
zaSF3uo96b1jYE2+KRM3P+8Kl2iwC1qTpe/dQAhneLvluOPki30y9MytACFJo9//
7ExCgfPqMa0j65CxhlTCxAZcOgSTJTGFGDQSWf0GrvTZeYizA/Fi7wzYr4GHA6nw
E8rDzeYAV2HJtwcj4zv9XR/bFC9KSJ3+AYT9TX4xPL5DbL4QfrwbVATrDGkqZ5Ju
iOp8bZgReRAJqs8c2wjc3OKFiGnibRr8HM2N6MiHvMNzIuRWxpvpFp9X2hfXm+S6
ypeNBw8VwP2kOQA98MGoRqU7MhKa3FQXph7PsFrdVMF5ow7ZJdVGf6IlmdGlSkGO
Is4eUP5ftd8OE4pTx5JLGKP35hmJmddJRteQtVdEPHnK7EExJbUgl7LJlLgS/H25
kjOKt4pKdVKW36KAlpAajcaNjJ9SNVTkSYgv8oe6suSufDnswewaGh8/rN1FHnDV
2MZESXT7VLSJJ1n/BejTE0p2d/2trIK70w8X2XWRCRzP5XW5WJZpil6ErqzrKT9T
T/JVPJ8Fwl2E0MjK/ypNanndYJ8osrCVUni3hBH0cWUyTChh8mcIlbxeQ8fkc/Sn
coZ1caZHaTUQJDYqRD8FDXUiaL8aEW4KhZ02Sr+D4/NWUt0y3KqZMPNz8NogAfgw
crBccQTQEO23EwOHeY+FCI5h4LWWOow2ry4RY4xw+ZArUqgXLg3gNUz5QTGMhthY
XIVzNMpS3TR0YPK8wrbn9ioYfs3k6Gy5Gfh7tYjCKQowuPjGQVLCUt3ZGxUR2wUO
bIBnZIi9SKBwCRh2KMLWC+0CP1TSNyqol+SOqWjKke3EkEB+XrgQZP9Nzk6sk/Nt
ar0QFxBG+9n/NKE+6mlHJ5nBdpuZ9SvzcLAMtpecAev36ZlyVwBDKoWHE3A8Usna
kbgRXNapso8Ckg+ibuBoX1+HffyJ3vi6oivM9BpDM75A2falF+V4muBm2NL6Ps2D
X7Dm2Ie7U8nEeo4EMFX9wVYEQq3Og9nB2/c7HW7Huh8i1FokzQGUwUF3InqM07ay
/tXAQVeS122PqPjMbIX1PJSQ+W2A9/Aq6SdDGY2g2VF0V79SsHDwEF5Mz2Co1iSZ
kDSm1YL+HjDZvQaElMLt2BUNoazQ+9kR2+4dP8tz1EgxuDms3l/riJJ9Q/FznFm+
SL5wwB34p6n09WJ7n+B94D68TNDQXrloR4BAMV+e+inNzTq251b2ZfIrIUDXrVe/
oiidXGhqUjdK+jp+We36jonNvzuN/x7M6M9dD19RC+fV7IUh77AeB0Gxeg9aRuHe
uIN89dRwWZZyA3B9ggIIdkuL6tvjdgZ0O2lrK+mImuFI16mFy116I7Rz3PTMk5+5
OPj2BS0bKTHelG9O2ldJnfvdS+3cy3H6fvxQMIIMJOWpDYPqe69JZqfEekoxJtjF
QL0FtS36toLe4iDSlgq0nbGN14qljoQetA0ynR5+6uvb69R+3ISMGQutJv6Oih5a
90szFbEUrkWY21I+CQRW2f2JEXKDlcuDGMGbf9ruGkO1pugqaySLsZsZCKaC+B16
8AlBf9+9cB7Tx2ddlUXEQ4x0nI3VD1/BOrpQT9XcMnN20mxwJlNCiOrocX/xNAik
6w1Tpv09v/p6e0hWi1Qkblr4MWa7AClMd/51X+oxduHVZaFVrLiipUFy+e/NDU1f
rC3IEtynjFXk9FOt9g9phiIY+XVMZmDZ+XdK0EmvfXu3e6dLhVpQ0Wf7GgDSdTSW
Vv33FBxRjv3AKxhpy0//bnAjmF9jk38D6A2ff6sAySDTdiwjfbJIYLAMudGpNzuk
29N4kgTizQn53sU1SXZypc6Ncx/c0DwpY1FGjXlDiaMEbtonlY/rMe4LZgCQ11Bt
rrfLfAGpgC+M1qn4phak6+amWYOjuAh0krXxwYY/2H4wdpmpxAl+Oc9u6PofCNsC
GhemPRMAw1qr+CgMBstRv2ekH8tuBO3zIZcEQrrq0TmbOUsj/4hX5BsDP0NGTX7h
fzw99FTiQ/BsPRUOLyyksaMrN/o/MwzVdiq995OFFFgpxgjRrvi1QfLoiviubcF8
ClSsq1da2kiNEtrZpoh0QJ+OGiVq6FDWL3psBRb5W9GJCME9bZK6F5Q4rRmrGUFg
4vkToR1BhdAeVM5FY/VhkE5DL6zu/f5ls0bR2BGfD5RL6CWtuxOB9dsykupjTqkR
zWpBUlzo7g7pWGewQPq75WKLGp0nXrYyWEfAwiglTop15gDSeq6GwopptVI1qF7k
zdF9TaSqV8eHwLcHRUGrDsX3U+s0DiDM4dPP/FceabsG5+bZnm9TVgM2V881CcZ3
yc/pkPro0gEr1fnvLhsYiDaRZgcJWmZfDnv3NadP1QWDZytg3+8Rl5Y10TvOfynk
7ccjqWGJU5K5JEZIyHQIRln+/kICsN81I8cpveaDoGt577UJqGPtOTQdxN7MafN0
7uL5LpYvKRUn4OCC3/oJO6I8SddoEhcZ35Hs+t+88QxTYOYYcuznRd81pyQiVfWA
xNTqBH+2+kigQjQWjxk6LWIE4yhNVkdsXNZxEbhBF1XaPoerMlVXlshSU1Pqqw27
pRZDqnsqu7fSjSYusRb8zLLz4qimnp368Et/7SClmQVuyVP4XitBrLrEW7vIThQK
2JDMyPiXDWooeoWw+V42CpvCtPXiupyRypbD/yYH6CY7MUT+eExCTQmNIAm6ctL5
134KtvnK/inqB0021Y2cFwYFxjYyP+GDScExEw31ckDlX34QDMVDq4Y+J6HPJkXg
fDrvk4u8U7isHwVeCDz5O17Ey6rUCmfxq9L5ylWeAFCuW9xmnLJ3v6HJKOwzuoWv
broDCVBXVgsrf0LJVol6Z+wRZShMrnj3id9e8vXdEUVkMw2iM/cMUd8622yWabvx
5gDneAyEW9sUoEX9S0srKmcfJBkFGwuao+QUHaxw7yiMmTurYgE4MlifsbhFfrJp
aIDKL2d9jkRpEPHHn55saYcuGccKlGnwGKmVFvSgzwuoC52ZlgvYbD//pbz0Y5Sa
aPIuViy8nnQjHVDnrGbsUTXhpJjiZyUQa8Jn++z6fLiHipL/Il4ZoEI3t7RomMB9
f37veuqsonNp36gEDf8kPNckL5s0eJw1CdAzibaOJg1AebIVri3NlJX6DjWeYYLd
4djVN101R1YxgKLnXRrvUHZjcLsuxLR6F32ip0VNucZrsc4yJQ3NcaWDuiBaxwkD
/2UVVQbnG2f82Y/PRwsGyc3abUV4XTQpsCnxMqz00GJb6p74RUqbF3DjgxUEh9ad
pYWGaBVM66eFMbXGAnYkR/Ed5RvCHYHaXK9iJUIzjpe+FEby0AOhcl30gGGDwz/7
VrOW0fiVbxg/dVPCv/+QJNOxOq1QHQvu2eAuzBm3gMEwtuPRj72RGCH5NrbOEjz8
ABRnVEdG6Yh83HNn+1OXIkI3yGcARL8clmS5+iEAi++Vns5/uTeBPhquvoUC8T7l
U6GnNe9tuwd2lNo2GzQCCa361/YO4Kog5KcBWCpTowkM2JgJ05tWfJ1rCltBUplI
nrso8s6cCzKAzpeyFTIrOc+n18zga1juppSteV9d6L8i8U2fdF306O19vb3DgsJ0
NNp72fOAozjWiGi3wkAtpLRRow5SA1+/SNU3WvPyceFm/26feYnOW8wcZXh8GkF6
dEH64Rvl9cSc/PdtzX2o4o4io27j/dvTowyrqkyDBahvyP0RfBqWBVerKPsU6iDm
3vC9ZpWsq3L+FrQowVtXsSlMfqj9Eq7Cpl9GVwFZ8gWbXSRqlbvOMyEYe9vgDhXL
W552D5jwsWa0TTzgKjiKKS6+UcBDCZdvHsuKeCnBdN67QXPrD3zu3+8JLtR69ZrG
dwH1GxRmNDLA8xVHq1O/7V17bhp3i9Qz20FudRY+5tH6x6Up57TmCviZ8VgCXPas
c1YOz/61YjmYP5yix4CLbElz0z4sjh3m1VoU4C/JK3t/EbPWJMLhDFEM1h/Hc+vE
tQARUF2K3RH6Y2GQwpChW7WS39EFUlTScccsBnXgd+g17UWXLOj8sO76mzrbeQRU
nZ+fU8FDthII71e5cizNcTdMZxy9ntseCyHRA82k1+nlHGtccFQIzuv0+T7TyTR5
N/p8bucSj32siliKQ/ftPe7lm7lzL3xwgYlqUMhSrSaPVOPBZvfrqW5dVbjqE1c0
ie7n1mj/+QMmGnllXNuwnHeXKEFYCPquuKGECl0f+PrykPq/WUtFtXhzn6qWQTCK
8viWCnm+qcJSjLch3Z+vJeFrltDROKTeHUUjYERXb4e3FeZj1OSkOJekx1doyC8Y
icjmtNx5CmRji1u7fZeaxaftlvLpLYg2jDEjSwtH4eAzr1YBvWwbDymdC0vwpKb3
ZdOjuH5PfHFOebDsXnxmGkt0HCAZcZP2aZM3OrDol1QxDdUNpVVxp1UGWldzaFWm
8Fr4jNbXXgKmARdWoksqvMW8XjjtHfji0RmZzlN+xRzOchadgPPSOeiNNyXusp5Y
FBE0BwBjwYnLgCVBKDhw5MSdBfGf7hTg9FIYyNtHuQj7qPUqONbNna/Bcx4bg4Gn
m7J6iW5HAtMu4w29lDP9/FOG/JtQN1Zj/bV3pXzVZyvwl48Fyevpzycu1heaFr56
wzQhBkqEbvjPUJDxNL8fvveXJLhqaJtVJI1mkl+fk/ORkk569hX1tj8M74twwhn2
cKVLk0jVjrOxgaoPwvysliJ/tVnHVXCgWvPUytuThx1QFVigFo6rPH9h09wRB4F5
9VruBGtEePT+eRqnlcV1k3lCdc/eiNwzfgSc9e4WkjravO68pFQMrou6K8I6Eohy
Mk9JoTv1g/949SUBk2nfnZLWWahsPco4ZBIFW+q5kX0XGeosgKwwZt/n+ay6F+zg
5kstX/IGC5B5z5mM7Amz/u2G8jGdDbbBOuJ20O6yGAT8I8BG0SSabcKsYeunF5kw
Y1PdWLP9/Bs18t2abXWcOXNzadWKu8N7MzFsOSYeCmQBWJEWUgfwfsHoHVqSTeTw
ropXLIha7/EJhsLU/s5pVXFZTdC9SWsSwpEtVV4F27XnQuFiaUmdgPMdgQ/ITRCy
mYRBOzs0C9OTr/FaEtFGdGxoXtc7JecmP8Jote1eVSk8XB1gl5kyGvVfZlVuUzsL
uO5sLQf48JUnSwaJM+cjLsmUfZAArNtyH0qOBKrtfShp0h+suXV5+Ur42TmZbvif
QEE6LweM+d4MtMi7k2E4hSIuUEctNlfRLtjYYyCEIZhclyOC+R3grM7eHSZrkbot
NQMGuYmMJ4mrNBJwjMUVjw4/POqjBiJBrmZctEgIWSq6FGdwnJ5Fb+DHEtdruCqC
3hUJrmlSL8kT3kLMdX6GNsI0sRzmaIZ2orw4KDFQm9SXhlvAPhN+f7Idp2YJTTV0
A5c8d3EoKfeT4sesQuU/opVjBV5LXTjuM87k+g/20F2J56AvfoBr42txvux4/Cq9
cXwuFFp0Tlcs/4my0G2q43ocrHPh/yZPSx0z4sv02sQsr6erUzlBa9l0xfHf2vaW
rpunKpcttbWaWKEfyQS2IBLz7vvEwa4zs41Vyt8qV3htS2bE/fQ00FzCZFDqReSH
IVrUSWiGS6miVBw4t6W2a7AmS3N35HMxM+O+6huUUr16c9jtiSJIdXmNkk2PinBq
FSxPKRP53thXBC2lnGUdKYvAkY/1d5xYhgfEPr5Cymo9nMHfX0ke8JDEGfPAfV+7
MZ8W3cxdJT3m+oIyrRopBQnLe0iTv7pCpfcunB64pU1zqgbwd+0w6OLrLsaS8wWU
hxdnAXXkYr13mRCpkO1EMkwFh/0wSehvNZaJ+tvEYqQR0opSxNjJ5eD9OufcO1zr
Mo6J+SQMsUwpiajS7gFQxGzJGhjXH+Dd+v6avgUF/Lw/yDHcl2jssXnXGFSiaDzi
efDv17GmH66Uztw3cIov9ChdNKpQVq4SUvm0pCyhf1xPFeGik+cUx2QtOkTpZake
Z7z5Tnm6tC2vl371o1bBk982o7dkUtq1liPy31egRtrlval98Cg5gK5iaA89obTT
9cgVw1m3wQ6kAnVwFm9PLffGhc4WAhYXbwl0h1GT8otV23YvM/KFDlH4KDos4K8O
vnKO/QRGb1XQB/duRidxxwQVoH57bXwe7M4xchr7yFXHysva67iT8vB4Jg+El0hu
XoJixfsIrsiqHlbsln2EZVYaJ4FKkPKHdPwDT2U9W699WExON19T0qLvfTMD+Jfp
lmo/u8gW4ZOFaoh24aGgTvyHC/99HDE3fWR5LYLfe6QnFqLhvauFmcy6iwDC48i7
Mbq8PuA/YacfbuH1gIE5rJ6yR95sZKS7ujGzbJ9YvL55jovwhY3bpAYKbPUsU3k6
KrTHwNnLbva8aQbpDZ3VfGJirdLhClFXDv624IGm05jimYDb0AnxvsKbqxq67zRM
JweGjNSMQiEHGn7qQ/XgpknY/Vrxc0baIqYiyxErnb465QIdV/zdxjD2xA3VF7z6
j0JnTZf1BXkbp5OzmYgaimTVUnXH4D7qjEdAnrakeXrtZELUsbQjyq54QcyAXZDK
eAnmI0CXqLmji0VYpOSJZoCvkddkKLaRvBdK/NVHFHBHauMclMo9lywwKrRLjCXM
H8CUu5P/ITYYqXSa2t6du95B+E2Lt8MAIuQ6ZFEx7F39UB/7EPTjcQooMsKLF5IT
F8kZTEi3wG74VNvIDxOPf+IamesgkwFtC2X9PD3V1QPclljJjpM8lz3pwEHcgfCA
DofmZ4eVLSKnGylQhRFJCGRD4Yu4Ceo6+MjKTFkW4RNLpGcijxD6bA3vr9jP+t74
TqmmkoRwzzzSeRFZaPapqW4fuzZcJ8Z8Npiq5BKwB1CF9tvKj/R9f2/9zFSTGuWp
PyRmK5RTW6O1kv4jD8uPfTNbDUCZiORv8152uoZkjQu3lqja2lLYyPC5QrWQLBwW
Rlk++omFilsI7dOxOMNAoYzfFZneexRXpdCjMpk8hXBFB1yoXB59b9PYWICanc4H
QO5XmmpzKs74I3/ZmGlYNB86wS9DxQf2HCJ0+FBCLfyM/dGTIEBTY7u0nIfoKntA
LOl/XDs59lqIk3ECJprM10FWbZf5l89m8q1t3BEjHtp/rrpHbGR0gnmqgQdgIKJF
krzohbqVpWzZkzDdRN1p+8QIN3L9aaABcEOwyyF8SOxzYaOKMi/hfmOGqTMCr+a+
QHHezX9OE0+ATJFR2Xj7j4mN+gpwDK3OmIUN36AG6h9eGSclqkR0k/qx8Cbnbcfk
TZ6KiwUK073omandkae22IJPHscMr0OazNspmKm4xHNAMWpeK4DLTVuhhsVDeYFL
LStm4C2/c4uZ7jmdEoGOY5mgGKQQgypgKf1YicAZAiwtaOBWyStXvAmurJJwXZBK
ZfebFMmDJfW+Kd7RoI7ZdiNCNK5BKTIBlsCugkQBFZ8Nnzf1ldP0GknPNk4M94HQ
izHS8xdSa7v5Cd1k+jpdU42LBfSkRoe+w0URrLdeUEUfROJ6F52iBm4XR47iI1mb
hdIU8nHAL7mI2eGZrKuuNUdMRkc4YjQBXX7s92lPkjO08LO+c63+qSZgV6dHH4pv
D8h/4cvaf/DUXGN80zd51UNDMuvbKq0Mf5ZQ9MVq2YDydy/eHD85UrEE0gqFEdhd
CemXH0faWubFhc+DrvuKuxvFF/aI8rPeyRIdqOK/Y2AETA49YLM988nptV2NMKSh
4QaFlBYAdB7Zm3kloAHe7KDGzSnvWuPdzhXBpW128ZyRf8fS9h8HHpCkyDC/uTas
DiSayfj+PT/pKEMrBqhI4VLQjuL9Jca65GAaXwd1ee6HeYi0GKkwPGcn/N3mgKQ8
QbJKUxOEweT+h1X0gu+19PU8Faq5UMCL64CYfWXJBFQuaFI+RcQdqg0opm67B0TT
35Ox1sBwkeSZwRuAwpIM14+sPjgfrJCFyxQdsPGK1mL3mi184aUx4eU54BvtFfNc
H+70QrHovytGyVZk/U9zOqWIqgCgCPIAAqTklEjzCHFeibSuqGORyPn+uSepfEdj
/qifNiTARk4w8pgotKtINn4LRAQvQJm3aRtf3qFwVhz90ZKDeBraBI5ty5NCePkO
yeKPakd2NeDcfDg48t/fvV85D4ExBZWDZFHzoFn9Ikkd69GG+NZvjzRfmRcvMM7F
1FjmwwzruSNhLKa/HEurJU4UzlfVtR6BXv3qxLs1AK7AUAdshQ74KU8Pu6W1xO8F
BzHrS68JnYTiyKdMRucakHFyAbDgm50TD3fQYELtVrHfm0U5k3H4XQwJEpKfigJp
KbhRosDobu/EhnSamNO8FHdvNW4iqrxgLLjhl9Up9zPsS2l2fGghhYrydhvQTFCg
taFi6eb7MDuZUcBtSXakYULEtkLxha0aVazorV3bq4Fg+U9iRN207lBxT7Z519tz
rcvboYc1AFe3fRV7Va4srLIIXbqo1I2rQkzsMaUDMbkdoCfuE7exx7sjA9ivyWjk
xtCPxQI9HycOpS5puFlEbjYaHqYWzivn2inmk17jpLU20xeCzf7u2JsZw+CZ0c2T
RHNSpjBKs4gfKnu0CcHsnWUZZiT9LKpIcC09wkaQTKM3KF8JUXs6YidvxLKNi4NJ
XOG25jyx2UWqKpMIlrR3th3AFB2HG0N4j0t/MO41SUkdmYj6YBqJUVADXt/VWXbI
4IkOk/nuJf0Unk+Yhp9Wd52Iof2lHyqjCmHkzm7xyCCc4nXV6lp6y+dg3NamWUYa
JxC2Kz8m5a1JOyA2uFzytGN6uAqBxNeGL2/cSLsOnJX/7ZO8Mkh7xwjA9v2E2snW
TeY14TglBXPKjiTkPcYt2MIGrw30ypUm+z+1EIpTnr/wBMSCvrza28z31ZBOrYdW
VHgB8SmUUPw+kkJZQ8OK8cP8JiB97dZXwY+uJTwHYIa+J8jcdd8BpQz/Id2H9n63
5PFpJu69mAxm0SgtFXMVge4m2feTP+ZmzBAaJeFi024vGIWjd86e1adVHsj0uptZ
dZNNUMrLMqQNp+eJgTP6B871CEgMHRwyPCcIrQtSRUhay2MkDKhecm3To9IgpRmx
OqlxyyY8MOCpTIHNZ6l1xuFDWaWydSrGx4BFmoK7Nppwe8ZvTcYaVE6VNwnpSVUo
82RhX3T4QkKIRm1JD1FNvv3aONjAQ1SlTI961E/jrF1J6Swx84s9qcxvUNRlDwrk
jkeVBXfER/w8secy+N+PYuZM6sgNCXtzRlSgIPX8sTpR32y8dtK1GBlyiIyvjlbB
0K9Taaqmz3wsHYGf7v2to2vaWVpC+P9X9ALldWSCiN9ZORkUrlsS9KmJg6iLqKtk
/koCeoN3496qQvUwJGfFyukbiIZPJ03IxffMOig/EFNAPhoMF5lgEZCygJBZgWLb
J0N2Drkcv86InyxqU3TXsoTEcMWXOpdSFtEd6g2yQhI90mfYMP28htLSCl1xu2ni
2Ko+xfvkekbCUUqPRFv/rJ3lkNEVKckEMA2yXRTzj5wQNzwjAxplH6I3vyp7WUz5
hUmnZi81YCaEC9Ske2jr60RqUgywsaCCU786KVKHoEFNALQywsT6rC3NDLuUtedI
6CNgOcc511bvFkiosBB9cbTYml3JM67iqwbZOS4mQYSyMVe6sQnUrvWW44Edttgz
yA1TWBzSEl7QhKkNd1OMgyvHBOoh2XfOhZRi73RzSZlhfSmUwsdvUs/OiaS5pvnU
lZE96oFad8npysZYFlBASlh7aYcQZ0GbWekuSW75mLb/01YaAXNmrQFAv0Apg8oM
0z7z0j/PeS7dhPUyjZVHnuPokFTkdB/WS3FK/ZleHvYXTTxxyViw6lVYPxfxCoZ5
YCqAO2Il93rUN3fQq2+YRDDdOQluS21ALqxfRzaw53FuX7YUNjlZqde6jRzsL2st
eyXRIQsvY0TARiOOhm50XTTHxJUv4SZL4PgC9JTWApBWiDAZoQp7MQS+QX3bzHkR
Cwba4R+xrGGztWVmC3sGOfGnbw0M+8nYqlS7mgPiL/5Lv6NKi5KP24WdanxCHMXe
7rSmSF1qXpf9zfhjrDDFJMjP/htbYGBwfBHFAOdLXS7yH2HskutjrZ6+0F8hcxRh
yxz/uDRFcMyB0geOgF/C3zV+t9bCNPVNrBuc+AR14PXyaIIjsPwYdDAi9baNUA7o
kBfHIj4DbNPzft2wEEvczkVTqjV0/fao9CwImQqHmyEj87z8x7ZVMw8DykLyF6mM
VZdKbjZdIq54WwoA9jm2VGENfYXh+VLPboF5/Ej5XWVa6R4jPr5faaSUUPxjqhfR
hijzHW+kWPeOsVcam5HQy3c0Gb1KtA+DqnsTl7ANF5PN6Lhp0PycTHRJ2XOnDqqv
MkX5qFGKSjVUaNO3m+VnPFgzdILxOVJnFeqMeeoWgFkGwp2aBiPohSfVhlzj3Mln
m4aazsRgEP0KSDMoCbSKHNfwmGNIXfyTFmIpkO3+R1RqGyRZA+gGi1KTUByvXCer
/6nBf5H2c7MJSRyjDLYnvp5MR6INyDnHy4Lqn4I1QWuYtqvddaJEQ85FSWgdz6GI
JkOVZFOBx6UHqZV48lFYz02t0hdA+8aAAJT9PrTb6CWVsUiODXe75MvRDyCBXrt0
eV2zY1vMal7kV5ClJiHafJmiL4HA/uL9KS8WWVuV1PAObzTEs01+UXEi+yatyFLG
dXTzEpPVD73F8UMmP0myKjvVtRQ2OFis7V3KNSkPt/8MdSjmjVevNOfb0dSJmVhR
9j2CZvbWGVFud/mXvy6JqZRkMqQmLUTAfNPepJKMnYHyLeGqldZ7EEXuzRpLUi6+
oeQxgtd1gZwmQcNtl5paUDnwA5CAegCrUfAR2CaGeI1qW9qYGo0wsX5fhuo/e5Lg
vRc4jvJ1K2zVu+i908329b9ifcQyrMbPWFtdkvOdn/lzPnr3tD1wyvc9VWWrtcPE
J1JVCff3+QFVANdKOeNrACiOU4GouPxiaezCC+sF4PKrPaRM2Qo02p3UuwYuN1dQ
BYcLPV2kBTuLQwVfqMHhOnoTZLGzo0o4NqinjlGR6fQzn1h8AFrkN4I+Yeqkksyf
aox6de1S7Xef5NZdTndYvClCv+HxpH1PKigZ/gkqmqcpkLAO2yBTW0KQ2MkGqe8K
wYjgQr6q4ONyZb1yZhNQZNkfDquXMy14WXiiRUoBDc/P0OaeV0T50ckn0oy8uLiV
+XiIspj9KSuAYRa8wWkoexcq1/lYuJNmlNqU2Jd2LYhHw6NQSzWkzdpYaB7QCY3j
iXEBrloWfrCuxiQ5sjXylhbMv6Thmn2E3TtYmSdEblo1EuV/4ckr6b+pnc+jvsG2
oapmwRBLxDy4EKTCNp69xToIZJdqJl/jzEJOjrSx3jKDQYeY2mVHfJoZntcIOEHB
VTVK59qC3C/mJtY31YPZUb3ZmCYn0UDr5V6o/8X2zTmRlidXRAhTU1xEtUBmLgo8
4PROjA7jscYUjBZcjPiCE2RxgLLhXQ6MUD0HdPkPLhcaFWz39FGtfWLrhd8qMIVJ
k6f/zHWT0GDdPh8SzWWxpPwHH2j8KKoLnvjDnrRUpo8Iy7BXtY2nEY73ULJRGQ4m
vOpbwxgdq969UluIbsnOsbOJViCcNRTE+y/DGWvIUZCg6KJVy22UAY7YqucUN0wH
5DMLKKHNGitRuPXa4BAabZbcg8wUnWt9WHNSkXKAoBvRlQ+Yw6mfET+cT2ewmwW6
3f1ASF8IkYqeIcWcjg175T95glRftIDqtdGZOWqy441LRw9ZJAe0rI6X3/k61rzx
X4SgQtl4zjxUYjBjIBNrhFoa2scTtInKCBK6i1VKxQvLtALgWrBxjM/FWGnJQz1p
tNyCqS29X78Q1ikKFYxMaEEDePG+m0IGXwF2A5eK4mduUm8D6ZKrX0ZBY5udiPMq
DYdxP2Z7theMGsRBJcCj8gpoTMR/PBoaSWkA+6wcXrXwKoIXufBTKSTO70c7lzDh
34iwWR353Ff5rTzKPm+FBIfdluA7HUq4wrCbleufz7PZK/5wlEf3uUjZNgHP3EiS
op/YUXSOkLelL+w6WbTggVb4VtMG7vUXXNZXZzc6wkggCanhGcCI0Wozjxg2IILN
BosFIbcUqgOXIFLhtjch4FJQwqlGCBr+wSpLEx0BjPB4aMFQAa2iPw3JV4EkUhS6
95k6iwAwXinTGNikUbLaHGsq6DY4xNp5qugE2oZ0kuVohEp4sao1rsCYtdhpHJGQ
7Q8uXdGv8SvRg+cyN1jMB+zilB7PzKaLPWhB0tMycXFQXpcgEl/jcE0xKMfxXeRL
eVPMpWUrR2xRmDRA92HcOdqznQYYhdQz2Ark40eHmD7MS2xOOK9mC1//jKoPaL1F
qDrFPeR84WdxcVF9nrAHTFJdquAazHe5iDbQRKmB9c+bVxf5JjnF3Tz7R0Tnuq9K
RvYXT9YR2ta/ITHu7426lSOrCWA0PPIVD0a+dsUXBSMGUL1gn/F4DrSWqkJaveeQ
egAyRclM11OtXciMFbEDUCul1ScWsmLT8AV8JOvovsuXqiFz7pGGXmIh6vT2XaB+
iSuJSQF6aDdP2NoReoIpJMez320iQhqIIS9F0kwNUYo2eYRKEgrtaKKIQ/WUJ306
FonrD4diN6lhfHxci1nmCWgUyRZP60mZFi6srua7OM/cWU1lhrDDgVNzjvfNAr60
xh1wFCz3agzGgPdTBHgXMOF2pnzLjlo6W5nXXGjbZr9AckE4xy0sIuCC80ravNlc
KGKPxiDVTFC0UJCIch33QKU/8U30eeAh4xqwqs1WzUehbH4qyPWfZxEZsTrkLIY+
d7JavZwHJfAoHcdg9z5cnu2Jhhei/1Zd6AwuL8jF9fQLFp9IdqaSGpqUsRVjIoZe
NrYibehAuZ/QD7ayqG0dEzPDnKr98C+E/W5fT1NGgrKDHIK6w0ckZmLiL6S2WrlW
uIS6i3WbfYmFPpwxgqvTG9ytCXHvvxqiY87S+XGT6lW0BFr1+9DkDyVPcOESa/Z1
YLrKoxtsRbRxpOfF/1+YLzCoVxGKT0m55sh/ZJbu9CPFpe7pSnURCtVCbEV10Jb2
+BdwavGaNyaxGU69/NJPNAexQNYLdkBao1UU+espU2bpCnNpX4cFIQGNOrqz3tPH
iitjicarftRoSs90BF4mm9STLxUlc37JNHS0u1YN/OOJUWyaeJiLN1rjQqUD7ilx
lsYm510figJXOuHK10B8LKnAI0G7JhQPlnU05Ec7nEGdy2Lfj82BpPGOG9XbSnGf
cRfsB+D11dQNamMYxjDRs6D0W1kAglSxNkN+OEJ7RSw7fAjrnV9d9cc3Pi07d9ag
zz0qX51mXJlTQjQZKLvIHcE9DR8HhVqpqFTlDbj1B5PnXoJL/KGO7i3MxgsVVAnO
VPjLQhMAYbTuMCrm9Www8Y7Qh1vyk49QIPmjykxfkIpRIs1HTAd8WLSjs12pQgXT
u2hx4QI538KReIRaFINgoDAY9jyeI/eTrtSkGYjHGErozuWkOUw1XZGJrYb7B+5G
VUMO4lE5PMu9WjzagqnUsgAs6+Td+FDfWIBClDmiDhNFOLBvg5Li/DGGXTN42HV2
uQkV2JQV0DkPqLYix+oDkNNRFRtCRSNmInZ/3RZvuWRAX586WahOJeJ1eVVF2Hj0
tPRRFmIBndDpDKMVhda1KM/JF5nbGVCutSTTmFd+6CcF5DKPPRcrafksdRaqVi9c
nPFupVIC+ZQlowJ5OtVSrKlAznGDySWa6tJPhMkQNPmYWm1kF+387e4Qc2Bpmsi/
kni7w+3MJAPWIlkDO2/i7+d19pKl1lRJyuv/2Ugoy7VEyXam8hn88vsiQw7QNLFD
RZsc0hW8vXjkbRhl8FwlL0D1/n6qAif1y5YUgntrPQohuFeUC/OQNCDzAxhL1Xf4
UwnRLlrrolBvGK4v+yegg4Rkl9008nFyadYN1hsnTIGKkcwwWlnpp4ckI7XWc67Z
zvO0MFwLVNk5cNHt0BvEMH8VlOMKoYte9vuHgJJkLj+2wX+O+bN8eFk1ZDNGFUFF
hlhVjQbHyt7nt0IwlTk/QLZcNb6x7gcoX+QDfFaMUENKbVRqi2PtbYk9qFEnpkjS
RShh6BeCYrChE4nnp90iZew+V4fMN14Q5tVazv31HC9pvsimH4je0ImS9xZ7si4a
njebTunW8YsIx5qG8LVCF1QWKNn4CUZmjWmUlbpNU7vQrn5ZSFN11ZCJE4iJqK8y
lrpiwLeEFQDRVwhTF2Qg2mq66lVnU0eK4jU4NTyI3oh1tKOYEk4800hxo/WN5ABi
32XouGNRVeAd1YtgHOenWMpb9nAPs+1N7cTVU65NNYz6kGcakoXz4ABGV28qK2ju
LEJntwJPygTwVez83JhVZwDYxKFC8KmAKva/18j40JapwbW7xSukZqq/i9HIwKyE
Vn8Z50slo+ECKp3dYC0njB4gzl8nNNKRREGiKqXLzRxlmdIt3lhFUH27Q3c+mcCt
Bubva0nJppBd2exf7TUUIFLb5+ON3Gss7GbzJ3GEUyG2Q2iRc5GC1k7Uw86vJgM2
lby7pFMX8DI91gXtwhZh6zkewHYcNK1ojwI1Q2qM/Frzwy1WnVZum2wSQjPKhrvr
bq5g0B8XdGTaMwmkHbWgWaZzMfdcr4d/aApVLtVe+nIBxOhfQRpJ0F12SGAMI9no
rrrqjKl1yyQMT3BziLCCxSJ9dta5PXF/7f+kIfXw0/Az/A+cNemCIhTPRDmOE2RA
/wny0MTyj3Zo0nnEGnARx/D7dERnxQPVNMdz8vlcasms/LMouPbp7n0zRSh7hgbx
QOaEDGvz2pYFCUMVsle/2iPNvZigBw3Tu/bVjbYx6O7inwymWZyG7CytYpKCPsYT
utZkA6i21XPSjsRpBpYFebC5cfw7UXnPulClFnkEuKjRWGBS+q2W+wQXTQTDGf/M
C1AGabSmwYi/l0bY52KQsI9cSGbydWbebVxuQvHEA/8Ru3H1hb//ofjIEQDowlji
Oob9RNpd0udfmsNf5GYJ4Wy51uacmA2K63apZpE6RsoP8gGd/3OTAG/iaUMwH12/
p7LQcuvbBtSLNqEDJZbDOCceENKx9ZAl9L9WNYo6TY8RKMOJtHOUoB+AAj/Bkfj+
d3RonFEFKVTmMy0//AjEGQuKAdOnw3jmpCapG/fOYK8fyJAaNQMrqzAqWCTVo1tA
W0C7mjbn5vWn/t5Oa66I5g==
`protect end_protected