`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3824 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTMxKdsgGXJg7FTY8fitmuVSWO3GiSp4yzqeEu3xDpDfU
Hg2NTTZIua0+CQIAVJrJuFmzUc01RA2Zyyno0q5N6TL8XG/wXjzn+xnHPIvlVkFX
1AqVU3n1a1kARkKsPWs5zpKy2yb5Xndadkg3ZT3lPMQbQf+ZAaBy/LvbY8WTNduI
Y5HL0tNe/yovLgIK6yZLoc8V9ZYqgxhJLCcaEeVys+aZGMTYTa8Vc2EpgvWMT0Ae
EIsYRVZ+8hpLhdp/iOlPClN15Jb7llYPT1ILutwuVEu/gjSpKe4+YRGA+5m7AinW
Sk0Pti4AtgDtKaiANmNLcX5xsyhX9ONICSsj3bptHfSShY7ygvdHXO6Whc4603Om
/rJ+bTLMnD/VGFECXa4Tiu/bzdTT6UxRWoMFB3ndsipvWH/r4SxTfBj/G4Gm+H0q
S7YTWwxGrKKHZIW4CNPLY/qfy0dzBkYk1cgXZ+VqSbdUCfbhNgASlGa5yBHufOSR
CSg+NcVf1Stj7a4yt9tiUDzg+9T0u+2mLhMOncGt+vuVij0jCFSapSU2QiJ1J49V
X8PmDMzH7QthYS9899JZl2ir2nklqHd5FpNZAryllTcoh/A//JWF5972YkIm3ZIK
CZCjeQG0FaC2rr8vyhG/SNN3Hn0mTzLQCsPICQUvlBGKfqDrc+hITjBngz4wd4eT
qMgRTBe7BpiDnU9nLGcz5cltVf/KApkFf3gDGVdnXjKvA/rkwo52CId7vqCMfGlY
tJVxayR3OfJZL0M329LIryPOAQUAxPAFONUYgASiGHL1DpOTkYX2FlgDP+z/ShvT
i6AFgstINwCIoyMRFyiBegmP9k4LwcGBoyEjOWHAUrEjHQhqUoEU/PvxP96F1VM7
cPoBSOdrFax7HWP/v+rdcS/gRGpCsjcDCDEMozAEoWrMm/NihuQ8XI7r6F8H/gLq
zcJ9N8DdvzJACA0WFg4dZGmlvDTHIrfwoXQSK6Txhp0YrDtf2uXNEkycJfhq1OZz
WkYXCk/Fp8T7fAw0WGiiNz5d7B72yrTE8S1IjX5hEIblE88nvCnq8eAJiNvn7KgW
UgK6Tng9FZZiBTKSDDrdV0ggV1VRLJ8G5guq5pf6iH9BOiaHL4IzFysc025HQqcb
Hwt2gCJFLhdEHu1rg2T+jpnb8F3mduEk1Zqqe3Sqj48p3rL8d26evTLN5798jIbn
hpaM0ACAmgW1YZ2m2ACQXJTQXk2C4pUyLv/QQKSwwpHYnH1YidyCmmJuYWK2GIhN
8bpm/2AdeEHPvT22g3ptbmqMLVSOKb43++RHlZuCJmSHooTyWl+eSENFF2WV+Pmf
hiElF9b6pBaVY/2ZHMpBi3WxdilFZ1zxPUoNXnVUudyg9MW/U2M2Jay4Ii8X+PK9
LBEyjHZl6/XzwnCV2FKWBneLQgGbcUA/LNYTaDiuBg+hYtPNMZgAcrhVfQyHpLOY
rk8aD+x0r4MsBROVyvLjpK1hDDzgK5W+iDZfMPFgZgVCzvR3Vcu/cxpQWYzLL1hb
PWZOXlfQ6Dk8xrv69S493wgbOl/n4OgLMEGo4v/QHuSRl6BmVikbaWUH8rmTyxWc
C5kkXpKp9mGwmoStvhnm+N2NbweCPSTClXI9YrbyeCi7KuQQZijXXu4fzl5EMsL3
9LFVuHiRVtdw2LJrtqn6kgc+8S0aKZXeasu0A+Np245o4Dws2iIaQcUceCaNdORG
q8AUGZ5zQnDrOtNrBcoq/pjkSIFFe4cRC2aDS320Mt8F8qF5CKK2LYFlsfKg9RAB
W6oYscEeUSEbRaDD6VLg7poyHX6OVMA5viKWt2POTjPFumcTnlXlEEPbwCxYcY9k
k08+dE5a7SAVjfSazXqW3EU8IAWPXaecj73CaWtoRVHxOdsukfmeb9uuWpsMuHV9
lcnw5lACgQ7cAbaf7OlkMRmcVBYoYyK7AXsfjTKwQMYLehSZc4b+k1FOeKHq/ryF
a1luFHsNbncy4wkKqx0q7USUUCqubuGypUMdUUdJjTkkZT2sBqkmtdQf80X2UO9e
kfgTWRkWFcMD2WqQBiDpOWoP0b1qLjT7jpPp1u38nkBVjZfHtdsvcAIOjRQAwwCR
n8CCbbjyXQO1Nc3Fw3XMwRBUFqVwV3eQEsW4k8nhHq9yTEY95GlA07vIHU9JiQkU
Vv4rpdxb9Yxsqjs9R2dV1DCxXHDMNfXJ4q+kC/Yy6Likj420FQvsXA2qhwyUQcAL
yJhpG7viue77bIAMxPwYHIzHVoUdKBGMDtwUc+TbD9617THUWoNU/mSn5m9QhzfE
T70QRkmwqBQmmrAbfADDBzVDqspfT2UXj1UOoyF2d1caueMl6l9V2+eVPKwJMiu4
ZlzOFh0HU4nf9Yy8p29W/y0vn7MPgk2Mmkydz1RT7/7NYBPYIELixdWJd9sGrjIO
zK0wwc1Z8FKah2FBQbnk/4NIGp5V2G0rZ32KhiwuBEsbLKl7+MppQYQhX+8DFMSQ
zoke0EqzRmFvthz4PRGOSj9B+/59XyNeOloWdVnmaFHQwf1O3biMZY4WrkRs4zW9
ZhDIdeTiiom+i5teCxuZxEZV9flHE8Bdmlpyd/9Ah9KdTpqoJE3QHZzkH3cp4yGH
QfiC5uusns50xz2D+SFSZFYuMLqqflDvk+Z2+Vjt3J3kpjpOQaQ+3N0fehpxeKpC
KRLC2QSIJ8SZEvHagZ7dkW4yaRRzYslY4K2WZHXQJ/8hq1sbYFJzA+y7bZ69kY/k
zOFQEM9S8XujBvi/IGiznqLQ1PvVOp8Qq7A1ndzo8GJ9dtJhPWTNXMZz45wG3l/f
c+8wm/kU2Vk4tMd2FIG7xvqGhhEa/X2T0DUMM8zd+omEW3Yv+ZHpkjxApMiC81zp
rruPrtyvFhT3fVffpmaUyrE0/ORI47Vn3cfZupl1aDx/kK4NAZQo7yp3bl8dpGBx
U02f5OyfoB+ZEgVZaUF+ddhTywbKCuZVnMTgHqObKBr1kwSG/S0duxaimNlI1rtb
OTdb71b1sii+kGT9CmiYNteJft2zNNe0m+1A0i7IGQQkYnH8RQFa5HkMZo/y+nul
qPzfP0WskqIrf7iNnEiBzJMKWMhUVpL2i1FvnfJ8aY4JVPmoKhoN6WnklZvnNRan
L2iN1qr5EkCECHXhg9NpDWPIxQcv98hB+EUAd/SP4m2cpeGs+HXassT1sw13E90m
nEuGa8pYiY3YM/8AbH30HGgf74aM9nP/8TZQXIceMPlqnBS0Cn4l2DHgJEPwRvzG
tWKk3yRix7wX1meeA8YOuk7EAtucZfsPorIwh79bPQtdhEUcFyhvexrgxERN4fgU
+O3x0nnnlKd09/nzRF7eohUmYLdJjsra4bzkyBTeMEuy9cBv5PMW6a395oZ95kWV
XJsrobz9QBEY8+SSP4Dpq4KB7d+mgRjj4ev2O2yXhC2v+d2fIfHTUj8sZ4VDBKSy
PkHZhaxKyYBHIH+i0o3F81sRxla1RODoFxcxrLfnpdEG45ov9TCjbEEggdS9EF5b
WI38Re/6b6aKBatZppjlDrR98hp29zFWqN2x37T7HRqId9nxZIRAP+oREy4xb6T0
/c0DZi+A4256ZKPDzecLO7QpViOQUNdS4RX0Pnc5vHdmeJeB4SkoZvKCn4QpkFWV
bpPVq9hjqBatdfuv2Dpup6mT1XkD+S4M0rbMGX0J1t9teiZtfgt1nr2FajksOkUX
MUPgf5E7MvxkMVT2kpVcJhvvvTcuXMcBap5U87/4vyMwrRcsOGWpqfzhU0SGub9o
P2wcJH1KP75oV/SC4lkKeGQGBJbp+3yD93euCyoOZpbeXEnptlxE1z4ZcEssj2qc
8kd8KuLHWmrJYyEob/NoqfyNwAm3GAK3bFEH/gJTSbzRYW/PbcC/47FUrhCb6410
32KPPM7RRZKT9PTf8jslvtFyVG/yVZMUGnB/V1BmJqatwyNtlcupaD5LMME+5icN
kcrfdlQf9BLD8KvsFCh3VOy6MKtLV3SQ482HH2sedMjhfgQEk/u8L5/JzPDpCcRw
eZuqZPuB7P/KbswRoJ8ab+ECMBQivwYbjggmkqO7xpav6lUxiswrHDdKTv9epkvH
uc4vL/rZKETJrsUTsVEXam1seYXwmZfPMsGMlGHUF0vUATJilp06ApQ+MKl2iLri
0P+SF2Ybqc6Mh8WvO7FilFOdiNyfNovl9K9wTcD6z4+DlQSCVdOlb5i2NvCfjz7L
GR/aW7f2xntZ+7gNsPaSN8i8I7qNhC7RhnDWF/sivmXoOdpal4ydH1yaHNSv8IAt
eV2vmtAOOFGWIBsaZdCpED40TdQMdPLoTn6keBSdJVD9lDkwjfJtz1p/3eMKF49q
OSo/4WszZC7ujTGRZ3yUdigbi7Z4x/65Tlh5DPM8ISMFQEE2Wca6AXYWcjS3J/oy
NCiZNqrRPf+/6CLsWcXlSWfxJ4DryUPVN6UffKrcujKX6E6jbPILROu8Rrr4TglU
BZlFgegBC7osI1x/cJd/wi7B7LHNcg2yap4gCtEeqq7U7GNdX0Tf38jRTIiRWjg2
3wT/uQovgfYEX3L8ynKmFLugBqy3O/Inq52UZyNwj00DyzHYhCvFkrUVryQay6Hi
WYO4cqH2GQew1ZtXktaVM5YGuZQZF9F6qr6SRMroNKTegb5VPh2spqhXq0FWZoke
P65sjzLEQnNkGWxPKNZs/s2cmXpwjaQjnN8AJ1Jk+/tsWjhfhbzjhVD/5FPoLaXq
Zsw8gp1JKzm3xbgxWODlRTdp/hJluGmRxKSlg8BD+T3ECNOQOdJCFXw8C0GYmJJn
qNcpKMWM0QJ+5YRczc8/T5ur81odaoFAEx6qNwAdZAlnuzymqvVwPjJGzwjmJCAs
4+tlqcwiMryvVLzX+DBvN9Zof5curzYsQ/u1NWpiCuh8BCUnCi4KMAxBLqWWlxWt
IYPFL5wGr41LRkPFHP2Zyjy6hUoD5KEB8sQ2pRr96ic=
`protect end_protected