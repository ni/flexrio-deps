`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
j9eMmSPGcKCWAR9PvkqZ1R001FU8QKTyJzFqNLn+qur6INyYDE1AI8LWcxAzfnTc
IpZG7ua3uuk5/kQKKQx8ZIPLfmv6H3t3eWjki8YIAtY/d5E7Gq8Z5mNxMYRzGGTg
TCMm6oOrOTVYlCXHE0X9AW696Z7UGfWirVibl8hs19hrFdeZKGiGht4r09vHR+Gl
FQQmSObM5aSK5wu5KOrK5ZUKGHyBhjnIQO5NnittDjOwxV/57nHVg0pdG6JUqyvm
tEgmCY36RCMRGWN7sekPtNHjqpZkmYrVX1T9QF3h73+8ZekZYd2xY2hpHHGYYeWA
t3+Fmb/6NUmoP8+Pt2hI6g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="wX+NBVcG/A5ruHK3pkDqG8ZVPdOz9TJPJ5saXZYSeQ4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
j/hqWUoxjK88VtH4QmjIrexFOSwtsLKOZ/LCP4cmrqgzmR/e71apdtoL+o8nlfy6
eZxDZMmrZmJGoazz2oK6kz7xJU85UCwNc4cxAsVxNdCP19vZxph/nCYZQ9lUFkLH
uLBkOeFP15CD3jG5/dp945fHP13J9SzB/L9PWvDC/gY=
`protect rights_digest_method = "sha256"
`protect end_toolblock="sqDZkaglKf+bDjC7VKm3lOELrT2Jlynh4UhPg2J0Q70="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
f9kZDbPp4NLiAOFOgATj9W35i3s4a7wbt9jeHjHVcJxMoXY8rb8laqS5bNUhXGW/
MOc7UNc1VwolqhkS7G27SLamkGClZZtXSbRcN1N+5kZpEaBEj1343vVznnU2Dre/
9Q117ZaagFa1275muC7rLkspAEMhJ4fd4dFMkgfYZ69bTJvWveFaKRF+D5uvoKRG
NCuyV14PM4y8rwvPAOJFJv03DUqCR9RswlLmby0zufOTJ5UbzZwO9wR9ByotUIRn
JfeEs5UtOmU57OWzYSkAdXFaMoowx3F0LqXQU4wR3aRHQ+vaAFcRmTN+qvRvFa7v
A5NfsbQLub5pbJr1A7slxwlq3fZ1qo6sJvjpvGr7xOh9xtDWkuEqHuCVyFc9o9Us
+bJpSO9RkQw4aSluTqI9nbSjg8ohnoQOv35T1+/9ZuRx2WbFc4+OS0L+N2B5gVgK
92UsizcglFjTLpHnJyQ6BaEOUrs0Iadld6SI5uNaf9wzgUak6n0sj5lgND6s6YxE
yfrnlJ5FxYMbINfDUbfGP3l9Svd05upnax+SgU9C/yD5RPwBWL1Kh23mnfr14Y/n
+XXiNdLVTFV0G335hzwoI9iRvd/eVc4YFOK4/ugsHS9xErJNUHdl/9cj43AWFDcx
F92Kb3fWpMYAbFxX5DkN+o1euBoYkDraHICqPsRS39NenPM5c5WnqqJeRd0//+di
RB0xIOnmx36x49mzOdkwKa0uCUFbj1CbFfolBoVZ4mIpnTlk0uw7vzTP4x1RS8ZW
62Ta30e1au2+JmgyPFNEiDkqnQhlE9fAXeifn3y142id5gxVXbxnwu7ePnwbhQ2x
ugpRPWMMTTc4Bs0ytCZS3gfTE5K4Yx2UaA4CN4b6oa0OC/WDDgKyL/kbkcqGSJlS
WDCN6cCwZOtv6MLoVqFQsvA4K/be3TTVq5wrJ7NunwtdVQplUVuZxfGoaZNWjcPF
nFBsb7vVCHsmELbzyQAEIGSDIbJiUfhMCwVIbbYBzB1bsLHy1WkoYWkTvvZVZLXt
7SyhZ8YxFddJuDUGHdhqUg4wTl2e1cuQk7rSxAx+k3hYWK5ikApS6NXX2KrRy/Op
nC+qQ5ostpwp7cASCstOZYA3wXHRH60MJPTf/VnLJtT8CUzGFbmR4hdvoS2gVbLS
8HpwlJPjtJ18XtrM4s03H3eE2f0ptZS7uL9aNFEo5qy9SBHX7yxpibChACQingJI
44tb6Ci5d+lJ8B8IYb0p3UMvFqpcu1Id/peSbUATtRYWClSYEg+j3ZJs2V+dl0lB
IA9+1gupCS6ugz0Mb7DFWZEUWrzIcDfBP0+y+y9wUg3pXUlHv3q6+CpAnwLnds1n
k1qxuZ36kz+fiIkHps9Qhyh9zsOegIrJTyJQENpAz6oVNhzuPao7ZuaCZcOXBl5J
rXDzyTC9EgLXYe6J8yAYJWI5YgNY+KHk3ZVRpd6pdlWD15/oyFYjalZYsDMreGXr
g3/DBt0pS6ekOVA/1RyVWEU/zphyhSKvM5k0v2QcolN9mwK2YwjgB0o4zygLN+bK
Fzhn775x5aWYmXbZAlgXQqe0yfG8f6MoQNj1Xk0aSRLMruyFv4n7gQww+ghS4LBO
JEDQwOTCIGkZ/GMqylSQjqnoaCgYra0nT6DByZp/7WsxN2/IP3yFIM7OxRzvF203
5sgrSYR96QIDGURbtvapoJBe3oFUqpJqLERr1QbzkGxM1HTI+LUnK91j2Okb4Xk3
nsTwUVdj83y2oVcUCA/+SdAZdbHzSYiE/J3HJSGz9LvyyXqhRtxJzOrjlsdZJ7yD
8ZSqUKS3HA57uiOdT0l6fmp0pbYbh+/FEQjmHTLNvJCNAXIr5ZYrDvbkFydGqM2m
P3/800w/PgQhrErJBZo6EBhnJltfxfKNbqF0CB7+2NRu5/eBZjKis/Ov5UauItJr
nNMTkHTS50ZRndVvPOy4DRk7feZ60McD9PiGOkyhUuTrPobduPnmRz92QVn0mOh3
4uZY2jg39/WGKGocfAymT56esLD5wWFA8aYTdmrwM8RgiCoaajAg3KOntim3nObF
N0xboRESDTVqxDsKrO34qy6BP0jWF3qUyCxNBwaLecGmSD9nyUVMysmmDyYISoj3
Ck/p6q6OGKSfmzy9Wk1Vl/6Cb+UIvK0BWVsxrqBvXHnsuiE6pMecCC7PJ5fcuT+6
TACku6sOgbjeqmu5Q4r+PrsYg+lj29na3sDV66WLiwp4FjnPu+lUV6jFucNkE6y0
f4tP/eb6pQBtYXpVopELIR+fmBRS44L6ki7Q9xbVgCfzq8TdkNg7qF3xBVG13mJw
7Je4h9yOfL3zuOsKRlTq+o5uUdOJ1ETm3BhMYNvDsWIG3XMmSHWnZI9rvkQCLord
BN3sXkBplGRvF8Sx6j/5aLevZz8SDOKYfY+BQTCFnvbEXLUmSLT+vD/dxGuGZ7vh
uS6G2FNE34i3iG/ca44YSzzzFSr8v7aSfwlQCxF/cjaDANHOHcI8fFv84KMjN9jA
7ND8sl8MtOCKbWBmUoxHfmAfM4W1wTTbq3AnHpEpjd+YUJwe4AW3yQrYbKcrDgeK
MQNzB6akS7r5i3bazZOu2oB275Ixa2qGPH+uhxuKOYPPwAJ31TgjdfYkEC4MKmgu
ic3x5p9USiJ/Y4becWwMpiFaxWn+y+XnuIxzv4debHTHGdLfsSPb6CUHPY0whCOf
X2qlh3q1FtX0ANTID/lFoJbYEdi9NWRq6+9sxNWdKRtZspb12K9fXmiWeNtPhgDw
IxR5mNysPIGMhD4Dl8P+MsssxmQrsuyLmNoN+Nr0aKsxgOd9VxaCNDlg7S+L6or/
s0vsTsgr3pR8TSCXmced9+UjNrhpQPf2qYo9qGpKt6bMIEf0nZDk/lyKjiStR9oo
vFEBQdOQrOZfszdFbLCM917mP5+3vZ6Xx7Aw1ewXzTyqrOaMytXAXdT+fDWG7p90
TEO29x/GasKo8JI8379L73kbV1I4Cjqbd5QtS5c4KB1JCwBJ5om5RIRWCDBz72Gu
nq14N5Ho+JppuwrMPqEpk52RM4QeqLd8D4Z6AlL11Rr/QL3BKkMIkx+YeA8k7Ahi
OHqUticZ0x9wkv9YSCevhD+L9wW7BtPh1hcD24yLty+ENR3nwJNaPEuiw+AlaOAK
UkQxVijNggtSSDzLMLwBSHc5bjXSK23TYm/mOL2FBtc0YtZSPR458/ZytJBSz2Mc
UpK5jcpB5TTXaNeBSrKx2LdL1FPrnqmGeUnW1EebRL5aaHQrwLApNvYX8ALl91DE
myCNFfRHfG4/S3vk3wEf2TMPqmcgSzQ6IcUSBf/vwDp7tNfb0H/K7qgNmIDZ/Ljq
Kd/UAKJULaPNuYhKGnOjiMiPv6gScvkOyw3GRqNMEuIZnFjVh6DaLQE9c+J8K1HI
eKj3kUfYN1BzAg5jkhrWzetYWhjUIRzSOOzEfqj2OWew3VVZdtSMmC68Ji8bnniG
JV1t4xdjRu28EeTeKy+M7evTwlYcB7ylD+l00gmy87nMHSwwyb72qLhFjD8y/Bql
zKqFepdUHMwAriHVWn559SPDYC5awJP4qVjsf9h9vut6h38HzVQhGj5Y6IUzGoeM
xdJFEDm/ql3cTq193KVbvGIPD19oNVaUxS8j6Klaxxt4YFl/wLTx5e1wBk1nLSRq
CM0Wu0ppsp6HghJyj8kXngfpGEzl2yzZtFK5HcJIFbfM8Rfyu8ioAO1Syg3pxw3O
m7sGtwgDkoqf0VemBOIotZIGszJtDYgZ9/axc3B/A8wse1kgzYKrFaud/n6W/eL3
IElfhOjwcPwkDzv4kVuzJ01xQI26/ohwvfiG5LOJh7kEakR/bs1y5+tRakbhpoes
qabvjH73CbCdEkwTJvY5TJ0dUCLxY8tZYncBWwteYqffaEy41ymiYNEfwAajZ/fQ
Z0egprZoWDcoLB7RZ8YrbCy7ySYDYabQq2HVev7gGbfBE1hEvE9Hu4wGO11L5KWy
Bn3/hXDESLJoWiq7gkTxE8Zl0Zb1WHmmlayTP/i/xLBtbdrGMw8aYSF5TnIaC9cU
5NMBX1Czji3+9x09O+eQ5J2VXUc6I+eYM9PoGblb0ZeVd+aqjocpj71XEbIXNOQm
LdFgNtOIZ+5cz89zI22N3omA9FchWJmXtzA5WNRFOXRxFpOzFR9TW28Ym1LG6c7Y
jlaIj3oD/x3/oYxu0o/ctft3BhWN3td3S+HvfZaowGis0PZwN3pu8OZ8uLnRBtfq
JhGPaoYf2X3nYvrgHvo6WEru3Usmb//Y/MqFjplfDteD5XLH4t9fVTsGxMi4774o
Wz/Fekc+Nku67EHroha5V/tBu1jqL8Elw0mO8J4N7nTKrQOppjG479APOsYTuGuX
jWJKdL7SFPuhLZkcY0WZICMyF9KIxsiNal7ICtY+vY7UNOHWDGYZ2MUimtQcOkuL
C2fZEoyA2zQQREFNToESgmTVsfUNjk/dpkoan9WR8pELw0Fhgz252xyaHEgapn8F
oYU8217wLGIVGzQblB8Koy9knGz+ny+sHqxFDZYRo9wL995MPDlu1H4oZu/Vel4d
I32sMUJHOeqXsJwNBBFK+tBfqybAoXxOoLfZNk3t5VoXlNqyJMPIg8q6YXwrQJfJ
FBvVP1+WxMrkgvaBU0ppZEU0wJjZRZ/KoZcX0d7VKfUc6p/X1noUB6M2uLlr+hA7
BrKtBW6Z7MiA9/4Lx5bb/x1df8/TE1vC4SYJIg7YVQeHlluTAnS06wTjOJIAVimR
1n6MVU6LUmFeHXKbzzbjyXI2TtAow4hLZM9VvsFFby9WLC/VYT6XvbzBdYyC6A1p
Cn78ohdZcmulI4ob5QXT3fE2PEJNNQT6Ju00QaIxsE3KXpnxrBVMxr1hdSNVzVor
GBB7GO5B30u0q4T8AIS6jjCUKC/X2RKH6wKv16/5BYbTynDoJHrOmlQ4CVkAwQkW
GTIzmeoCPSYPNh9MB8Fa/cybbe59N9nl7shZppEPyD741ub8B+8zvao+7RuEorHq
JYALRvHQ3pJzUh6HlEqhNly9vbSeseT/Ei1vKhjeiaR0nVCwfM1eCZSKrxuLDvod
5o5iRCAeJ6ysHVBzepK6oXZapJBfKrvILX1bQPdgbmTDsUhwgOFLZ+WMQhzWvolR
E7TfpjTlR6W6voBbuBt21wvbtDiNjf2ErqNhp6RjEOZZTc+lA3r0/Qs+FeSSUonS
a2Wwk93mYzhgSCu4psaOR2co/gwkx1Xf7ZmKM1rAEfjiuAdIma8HOe8m69EyZi4p
Dsn5xWYySOUKm0dAkNT2faGzTZ5r/WEnfP1WLx83b/Kpd3VM9oTW1aJYMwCk0Nly
xPOh3YAJuW+3Qf6u7n1oh8twdiohyhjJzz/kdt/EoEzzV08tF3dWZKjw7l3Yegze
GnHnIUSWyxy1QBFhKPlH0PsOmn2QgUFADLnzFGGIurHaMmogicLUSpfLdwQbul6x
gXneKOy5IMzxxiQxvhT1WgKLrPe34+TUAWHND4PU42p/BMMUYkqTaRus0LtXvV/O
TPahpLFKRw+r5nyEmZ7iLCODdYwm4q21pOrB7yuH+wzE4HoDevAA10v8p7i/TEb+
j7BWwcgt564ufox9XGuRaCGbVCMdi+ng/GAaHTtG8SrK88OPokjrLAmmbYnUM81O
ptPwIYQSf4CRmZP5jL0KFO2Ud5hXHGaX+SFCsb/waFbshyxPYpjrGL0ruTAw/v2P
D2Vf4R+ZAgEoofbJhdiqxImRxbOe+OOcJ3L+3zk2bcEiRYDyIXtTuRJq92Dk8jQq
Qibn0x5KppJs8KOMr3oHMAZaTaKymdD92Djb1NSeCUpB8TG9Fr4cPL/dvWw67kLK
ywXAf1KTtBFTrFgvDq8MxF0Uk2YsybOS/k2r4mH/bwCg468JVF1CJkUagid9/Vl3
L3b+rNZlcPAfygIegbV+0h9c30+hzwwjdrz554gqx92NCxwA+BR7NyLD22OopCTg
oAdOJYszLXsFIvG1VgNagj0w2rg+Ul2F6ahe53VB0tMr8D/SY1aCIqoHcBrH1sfS
UjIG8fDjSEd4dSw867MSF5aCq2JZ8UA0xGAdAOSsO/l/jvhBZXAIOxDGVNM4U74E
mId9x7s/qAZLtjLyOFrdI7VJ3CrxNVWa0iFfeC3aU7QGjp3tzjIohqJ3N0KF3SYH
oB2F9FpXFmRYJlwW5DaFaDYXrl8LZeQiz8dxm9j4VqAtAOJIi59tYnQsOL+g5gpg
oxslkN4E5p8DVooMqyhs9bdIl6jph3P3gYN6nGY2Zo8ISaFaTXsMmeVqsxBnkkC/
2ynENevvMgoXKYlwIjP7imJe9tDJE0HGP7+QtPrfyukQXR0508WJDEPjds8Cc0ze
ktVbOJP/j2f6XUip1fwIr4m/e8fAJWqhZuBeMw+q3IUvBl32KEIQ0P1W3ejPunc5
e4wc+DRGJOTGRu+eJv/OKyx680CXz9IIRUl7Nbm19AHszoXmaugDh9/VWFf6TSHA
V5Kr/gMuEhxnHNPzbzeaDqrxQORsc++J3hdVu8nNlWGEHVW1DduWjRg1Qma63ZVk
CkG3a4yf+W7y9F4rQsn8v8/Ew0YDAAHmtG230Rb+QprMlKw29eOTiT4Q8VBbBHQJ
iKJKOEunFefZHasvtEBWJQqraoviLVJ9c9UBSPa7jYNQHnCWl9RJdouisUJ0O5ac
5NoHUARV+wZW5OYXzJR+0UVtpcKXAwfX6WTZBz8TjJ37AR4zfcwnVSHH8jd69V/F
EqEfJAFB9VBcj6B4P6ZYfBjuzTPJfxEBpXLqKRPx8fl4NXFHblaHTGiXvXcxGkGF
lgiExgaXBYZ8cete8xYE3SVEUPubZkd2SfheBOAMqZZGTGhx8x9wii1vqpMwPgbQ
HrqovsFRF9kwak5sNyn5hNFpr2E7ys0i/Jwg0S05LVTK7LnOGWJWRVpzBim9Q1v7
1Vk2inON+b+DLKjF9UhwN6wKs2k7eseZ0xgTe4CjHYTS5V2ZDh3i/dY0squFrR+S
DDK9fpHEMbUKNnbJQ9Zdt4cvq/vgem5VXg7hfzOUGtYOaYlIzA+3LntSqaHVv+6e
6W6eeSqm0qFHWCMlssMet+0eYISARpxYHbLyKu+wbcFd8Aok6mIqjb3UE0cJnPkN
UyWA7Aa7bT/xHzCyeMmzTQk03REFUsn4OOGXb4NWFWn/i94IktNdh7NOyu+5HM9O
K4WRPZWeQTCzotBxWMBz2NypQuUX8a2bdzI5wt9AgEq4MxJwNyA+6spNaqiQahXm
SDwUc/7NJbksw7k4L+48NtzH+EPsahg4vxo5aQbLmOeX6H/45+DI4FB2MGHTgr/m
Y4XjDXMC+H/bqVyC+8BBDX8CuZWR2xmllCbxYmR3Rh4gMulStba1P6/C9Rv4h04H
kCVXdudb5ssg00zd2DWogaBytf7A/I7Y30IQI/br2QjMNpPtmjSjR4jUAw7CG8E4
3Asbn3L33+FiIXHnHhovg29FwLXZ5nVgrpGwgKI5H3LCjhq+dX7hI6DvNAWdntcT
qNHFKZv/SylE5ORfOE90MeFlzgjyUjbTxk8bEajsvVS6M3Ja7UHmlvfUH36dQxpL
AvRS7U7GZC1LortZ21Zgzj0X1h552slUYyTPkAr1Hp4YZmpLNlzu/ApFe3kbc5Hs
2U9cI3Hr6bONhA5J86metOfk9cuhFGrJkIRPY2jMYmog+xkIDqutBR8+cETg0O0T
fwuTjnaG6qnsrtWLgifPfBHNvatOPnC7uxUhofwYMFE3gk3eGF4fhELmjRY6hv7C
hOIzWGCVPgPgR663lJkZL6r5Gz6q/i5LCQDmiD6Flq/mgly22beDNCycECIrzc4e
GtLhJj5XWj7m6NlxnpQYdoKJu6b2e3ufVckODhhsxjSr9dQzJVDfQ58BQyHpKddb
2k2ptMnPpApSYgLYPsQJ8udPQYyxBAVgWpAqIVT28i33syTTep0CTocYqxfrMUlN
7YcBYL3Fdpsv45vfBZ1vLwM85H3p5JUfyFVgIjpIXYwfvQ4UXoBFTiADR1Kj+LHw
kAi++1MaqQ7AeVRcFSic5JjfMGdakIx9s2X/hjBL6U7MAARXx1txP4XXyLGz25Hm
oNp6nhAAHbjciCwllelWz/iJQysV/IpNSc7WwdFGXPaIvydzVYianlPo5woWCPdz
N1AkPHYDEOpk0sVdlzpdHiQe0e2kGQmemofNWAXb3TKJmjG9tx4TAL6uixCb6Rn6
5ghywVxOWqYKSG9v+ZGxKuj+0jydbgiG8zixQz9INipOdWCBegSXCE+Ax66fJp+s
WdjVdF0MF1vw6RlPrbDjHZttbms/TOrdhqcr/GIIN5tO5N2Le+15iZg92BxmI/+N
uuwkaDvSV+KqbCCbq1cs/bnHJVlOPx15O+zobK7bVJRS9U4WSf6mVuEOOWKL22vc
fDA/kEMicVapW+L5QE+Qeo+JWbejAear5GQaoLLoaHDz15kDoYOC/caxLMi2q9Ms
8sndMe8FZCv4cn3omyGOLXHkNB/0CTmvSvODmm/xv7mFhbNWVdhARdaHrhh7DL+H
mm6z436NuXL7B2PBA+41rq6Y4Yodf3aOY85S/yEqTvms/WoKpfIhZOWnyk2GrmU3
Zn8mDru3KSq6oGA0Ji7SHpUYx5oMFAoAlWixI9RKXhys/meWpX3jp3ynGyqVpDcD
iwP6UZt0p/eixRxpxmEzQnL4wjjV+UaDW20ZegjOT0mgFl2sBtmVKCq+1Vec5l6w
i7ihNCu3ieAJJ+9g8sxpInZ1b6eq5ARqNvYF7ScImGSAzwqywPm5MTGQ4/lyYZNI
TmiWtZCBnkgh3F000xXnfRHwJpR/yCBbb2cZ+feuxMhw6fVFkz7CN/egQBgX3APy
yT5eS9XmPWcN3TxlLCQ6WCuaxO9s5kjNQNT9PQn9ECxC/vupIRTOR6apf+0+1FJT
3B8HrQF6Lp40IVGLU9wb06jKBG3NSsiwKK719kA9C1fsD2VBEgaaUK+RvVnZjEa2
MUUC+87bcSMzgDhbtTP8yyBEXsMU/C5ZlfMZqvJnRHskrAqrmmqdldGFoRnCu26e
rV1bxPcuSJPlC6RaFfIVYtQAlRgDGPEXJg+nhrpVE+KQL3EiNlrEBti3tOoedvPD
TzLmQp3gdPxBCohZ779FI2W4+EDUkQJkzkSplUbGzBLswaOWjOj/mtJO+wzBnE/v
y5yQMABaN4sukmTNELQpSbigog4QJlbXiDXkDygSvHxoAyelBjleQkZ/FgTgKmvw
7mcUTNsNLIKg/62PMpqpgmzRDAYHiqAjS8fjVdqxLzePAj8x09g7R9/pfoci39oc
Md3w4KBZCbzAzW9LbylGG9Qse422Lln6ZwYiYuu2ixF73CtgG+BdiVI6/3YgjmPs
apBsXcNUhwzgSEMt5UDdc2mc5C3mITGhPiSNF7T6cE7+ZWPsij/lwqvRGfjomsis
8elvRjP6wcKXw3ajRZ9F+bSUkWWFyK1C0GiL4Hdmd8GQ9RC6Z64h/VRgiYgjUnA5
0/YUdy5IKqFzWQkEW1lo5S0zP+7U4k2XZQRAQYnAUIYzgzSiUXpBiJv712pVYNuQ
jBxfuDqdWFmH7lcrUNFo/IrD7q2wZtEEbiUBuI498uEozmwpL0RSNlhGzfapdqlC
6oxoxKrdKbeA4yyFlE0UvjlseYIm281wG6kzsekUn/J6yuf+QXyop39YQGWT2AEw
oTaxdU70luevsuAy5rgDLRcffa3XirJVN/rTTcHzXsIY9iCls7ql4qYxTtITcaZ8
8okGuExQojS7lG4/o6etbbGzQn811c5xtV448H6qwml93kem5efaKhSrz1GuUAR7
hSU7vkZdyjRsgzz/tR42jENNnijAc/eazFFO8mX+YbB8Sx6PfZ/isNJaZaGJcb0L
UgdutorpA6k7pwiA9Ig2VTURHQTMuLqKwqd4pWbT+kedAV2VkVeTlSWRSfLhceGL
O/o6F2F1Ix052u2QE1zhYIjZYCsPIUyC8h+K/am0Gy9yJ6unNc+0WqZxuyST4ywb
aCsXz7WNuWp4t2Rpyn5gaEG0EQ9VtKc1QoV8SnshbV0reUz9FLljsctnyBEnTYoC
ZxvoH3XHJqofdrpaIkQh+afWPAGFg2941NV4JVbTiFPlDrWTtLNv7mw1iJ3XjckJ
wdqNFrKgNUma/l3+i9u0rBj88NCIpNRrNoQMBhLIbY0uMkyKvf62BniVupp9kCD4
h3jk/h+HhEclt1fD5Wx53ENJPWkWr1G0CzokAvjJy5zM8LB4BFkGou/2gQY0Fkll
78REjfNFpLQxI2SHVEAybbzhnYhWyfmil0LNDlCyrzaFlo9j5Y+SVgHz2oJJsow/
Y2gCjdY/+NiXEYVQwQ+Hv5C0HNi7VEICb3qZyEdl7Nw0HvcJ9gJ/wwhyLeqn4p/Y
gR13lXxLwz56nqXFSJGOxS2nRAWx4MCGQ/VXskFzuiQncUpXm+8vnsbIC5TAaYAe
XQKGPrZvOXQ1udU4wBQEsRyrV8Z/RPMKJtIs90ynxhrQaN4XCLSuhqKmV5s0exPj
Npomeq2izOcDZkYQXudbX2WCN3463DVkIpzchW4/6SOnKy1Rs6G/2EAqN9zoAVLQ
rsljgPLYEVoiu2dTPcPcnzxDgp6IQ5fFngod8LkmEq8TjK1B/f3hw6KdYwxxxJ38
8YS9U9G5vDzTVLZfnmRNcXuUNHI0XDPkpp9ouV0tA0SsmCGhlLTDhSdFv9jLwECA
CD5xXRcDIexgCnsAqkVeQjPp/ROvqetDNYrU7R505tM1iiZvArc+UeEQgf7voO2V
Pmqe95lfOMKIMNLWSTWV4Datc5eNGB9BXXfSTvk3yA22/RkCEIF7+8qYJ2+dDZ5g
dU4CDhpMYT127+mNwoFzdJxycYSe9qh6Pu+/4xeR+dk/OblIO88bcUCI5ZeF30W7
/svybUof4DnR0SppMlZhTX88DeA2Etu7NOySCfc8Lt5Ie5wj9DX70f01blCCkexS
OqRs+H11gI/d2RWxjd8K06kzuJvvENNpRJXBMS4yCZpckVIpkF3lnYq59tA+PmjX
EuguTSZgCLnn2LukO1bywMGK4hyFY/30l+LC18gEAZurq8szRS0jyRLK3Z2005YB
gsK/7KItDRcJiQN16IV3csru59S+ImME+tONbaD0cA/HusXhwKDkuCCrvLwDR5wo
zhcDw7FyGE/R4GfEGsvkSW2T4+UZP04wbqwmodR087js6QeImFEPxbzhYk2tTx4d
xa7qnDgTRNTiehQ7vYrhX8NRMQFWzECSSOjgxu3YutCb2ewJYF6Pz2F6+RtHri4F
fQMy7inGa9YPtH7diiNHaWYv4K8xwqx03ukbxtUS2ho6NLLNOZG9hEMcSNbBt9dt
n47pxfkBuxEaikdrmMaNXUbsbwVE/VD6RR+9RthMKOiyaIsLwMC5aCeOnDwclR4o
BQ+M0s3x0XaNGXZeFVCeyRNMWCF9FXmPY9IjjbcgnPelCcDbKQ/XUwYaGHx5V91j
gT6/1f1YxJbWEbY3Va5epC2esWGTq7dZVz6P68MqelLVX4ma4vMU/1qeBLNhf/6Q
iLLEhjVgp8Nn8sW+FtebPYGC8J02qEA/xnOTZRipZdwVnhbEtxYi+g/z691/O3Sv
uV13FFWIAv44pItt9iIcQqF0aNzHzrxFn9pgbblrcBgMqK+IvEePJGUMJ+PM6I9T
E9sThXYlKJKReJs+Ho0AVenRaogw0avN1dCU4yX7S9CytbFbPdD34KK1c/zRnTtc
QNw8Pl6GTNbGt3TYKR+Uc7z5JmFS1pnRLUqzJDMIHOIRlrKD+px0ax13Fx5Zqfr0
Jhaoy6ptqGrLedrOo0xuOVgkZJuazhVQQuYWc6lX1iGlXaqu+UaquTtKi1/9Xuow
1ikYDuak1JvaN/GNC/9nV9cGuBixuAIRObyCwFUpabUZmg6XTgsvCKthH38ih+Tf
8TakQlT9+wxGOZhDshXyj1Ks+BiZoa0ApVMda5d+W7lF9Ml6BBqvug47QZctjCi1
GHtSiPIk/6wu6gWJ9+R0bzaslrA3pFJHHCAhjhtcE6Xcj5zhFwGfj7+PxTIovnH+
mQrZD6A+svFiU4PZzr8cwikXP3BxCBIcUFgDCqDj0vCqwK9/LyDgvxNmcbgz3xJy
waPH3HXOSJAH9vMyTKvZuoHfWK3M7CFGFv89c0PKfKRFrtlKmRbMJnp7z9LtEQw1
boT7Gt37vmiz+cRFLxfQbZCnLEmONij+i3hj4pUSE0IzX7xWUmmFLRKreTioD507
hI7ZCVzjzeQbB7IRm6X4V544ryJKE6Q1in7ETdRv985cVVsZQHOKdt0uW4uyBTTq
s9saCSr6/V1wnTGAzV3Bo1le7qkQvsnhAsKnQIK7R9J4UmDw7Zbvy77Z+KtzcfAe
XlHyjr2GL2Hz43dnAXkWML5dELaS79rF4I1FwEaRJ4cic3Ynxoa+94AeiULKMmxw
hFk4YIRtR7QkpERB0zmhItlvNaOistmJ9f8g1PQ3uQAgK2BRNuF4uIlSKVmWRw8h
BtrPXLz5dXTcIb7oJ776RmY5oR8DqIiosgqf7KxtFGTyw8q4aXl9udSa9AKS+r00
/mGrx3DHDUaGujBn2dro9JPF4a17vLcp1R7XQmI2xiqg4uoAMiQotajfzb6FOjDI
eC8Ag6ssxUQaWXeSzDedYJDQRaRs3L7aG6VBiDViASsQbKw0+X6+Tr3KLhm6Kimp
/Z/sZDlgX3Bo0f2wZFkFam0M3Q7nlZokMXTYkFVS4uW+ZU7aPdOKdC9eQuSNrq5I
DWmipdmcqeUQKwnTJrwduSFFM5vJ7BAMz+WXsS1Nr5J+JRw4fQVPJV+Q3BbqZJ03
mDbxU01/4R77xsC5Vi8+Zhdl65DAcZG5UKgh/j+3iGZeLqOCgT3vtZ+BNT7DAWgp
o+E1rMAR8dls+AE9N7kFBEnSjwAHT9Sdewxe9uS1ZBHWwIPuSb8zl1R6t4XGmYRu
50fzLK1Z5jakMW/WXcULhEjIfCOTtpWYkwFpk3EeTMVEwW25ernRjXK+EsQPdOkm
981m97/tNhtU0ILmFUlERLPsmFPmAM7eNTHEU+gGS1HHhisjUIhmvgXdP37qi9Zm
qjA4m5svg4NP/L55OTdDJTywbZgb+W35pu8B7BbEejmLVJhJmzCGminDUyURQa2S
kbplwK2mxxYkGjI9WqyUZF3PRm9sU/KaQto0DobaWN/zPkhAOg5Ahxd6i15s8MAs
qXM7KyWunU7yNL+9qY/SJ8VzuJpJZIwdJVVozdB/TYx+M4DgroB11pXh1D7bBHzT
1vI96pLVMQKVrfdMH0F0gIk2N3wFzSscKotvwDa5pihuT8fsIM274koO1vsY9GgO
CH4ZH0csOTYZJgnqiOeswizuoWdDhM0tkahrs1fubVKNIxWFThEYmDvEvKPCxJhY
nEPTjXt2LGKVY0O4DRsP8w1hAvxGzR+irpmmY0StFa0NIu68SstFB97ncufDux7M
frF4/2We5OVdbxVkfZ4D9WXA1nP5FeAy7DxFaa1cdZqGEw8BNG0/l0gvhQLH6mb5
ry093N/Tlo9X3s632z/aKVg0fJHIfVH+ew+g7HL/jOcj8aV+ca8ehIdZBoOZ4+hC
tGlducE0G3XoaMgm9YumLQ07RjkF7PzhO0+Z5E23hDHvXYqX4XXyx+u3s4RxiQ2/
lD9kAPkLe4zTeQE5LyFNi7zSMNf4ZeH4logjTpIMteRIhXs5bPrlCJZA0tTZDlZK
YFBlfj+CR9rriNG3HONu6jUjqhoS88XnadOtwRyxdlttQdSVxzaUuMlS92t2hKCq
zucNFQCPgxNGVoWKleahPCMPb4O1hVd1kDZlFRA939dstNZUZpgY/9BlIxDJvDtN
uXkyMnzKYa7SHtO8CH3f08yAPbOIllevIkfp1uJ1boNkvEYVZjCpI7s1ebYd2iFt
E4XJvoGMb8L/3aAnOWkEYIWMOOn74amxWRUeLkDPQqqSqQPtMgOv3ecZZFVv6UO1
aOr8laDtPY18RV3PhlBcYqbLvuAelSH3zra2yd2H/v2IljbKMbhAgHBJWPA18Pos
LiBhdDnIPvM/RmUUBRymAiw0zw0fVkEvKreUtJkLBAut63r4QNKyCHZOCFM0wV4j
0GLC0JxqvPKdaJAP5zMxZ+DKppo03i/I/jhk+xUniFfO9ANpoNx0EBTeTBe3fP4l
UywsiKyYRjiu405GprFOHxArDyLseGQfhoYT7OFn3EGMHoyp0zATSiIiSxJOpG4W
NlF1pYd+pUgQ0/R+afQZIG2WM/odrbDU30Ngo1rMfsE8luw0tlnK90iyQuMUwANm
o9b4mym/yafh6aXwfolkoPC4FTQaBB3BbsyXc79oGrOhfItoIcQrk7pgzLf0uhia
8oFsJoDXmiqIVyGeC/6TZkypEupD/R8DsFHh6GErcOXqDMlCSVnZlbLfLKrSBX3a
Wtr2szLMaCg2idlNAsTrjx9C9mnwmJDFcQ+zU9c9uKWQmp+/LHVIKTesCnerDVbS
E3a+a23dvXryOkMUnHigYoYpf8lcjgk5Dn175rZTXzcU+MbFf2O1HtKyd355k0fk
WBYcZTSR3I7LR+ae4+LZFTzvUaXX7NTym2uT1jvRKSxAgm/THZBlSxsGMd2aU8KH
vpsa1zJVqHJ5dtuhQsg3rayIpl7+UUhpgLkF2uMyP2w77ZVfxokcFBBck2f1kFpU
GG8QCECHHq+4lfccvU2b3511J2edyFNYGLGsoFTZr4mCSv7loO3Rxl/xjU1nm7sd
6FxaAMFSUf3vIZCZmH/3XVZKCQOFLD06HdAQwBJfBzGfSy6Josv9/51FaCALEk2T
91kPomSmmSnp5S11jYmur4KD9z5EgsnYotH1SRMBh7aHeCPfFwsV2v/jZEvCyxXX
SYcDG3jnDfZcivqIMSDH6MYVJUt2Ovo+CLpi/XVM/A6KjW4WE2iZXW2eptvsx4PF
ZxnBzgxa4OwFSPZPg8hUqiS0G8hyQsubDueTr/iJ9ioDLFxkXqBWzr2q/hA5AJfp
j2Z0viJVjE9SBqrDrF77njP9yFuWF5NQLo9VXht3a8MA4yTBtG8L9xHBtBhbjNbC
isHbbdM7sDwg9IYjwRwOF3UkLlDrqrO4p5CUePNK7O2qjPCvkMBnBIErPe6QJ5mJ
sgvAxW1GLO3F3pT8vLI1mYDKtJ9APjD4UUtgq6z5nfkQrLnqqLU7XIdZVTA5hYtv
xPV3aLWErmpqFw4TIQVHq8GPhMGORYSs2A8A2OthXtoxjc5qzJ44USsRVdc4Rzs1
QG431Ww3fnSsJXobez4Si5+FrItetFG6K1pyAUfaOKG8dTgc2IBNvDxssdS8gfkr
m+My8z4NLJ3R0Jbc/xmk/IVzAz5SABLMvX5PUCdEv697FGfGA5f7RSSJnyBDjq7q
VLn85thrkKpNlH/N8Dv0A7AM8nI5P77ye7+lG23gfpoMra1V9nyk8cJqlA8HUAJl
kBCNmM+8ovzdqSKrmN1EsVDFgr6WU9GyTGrPYhj6YszCS3y87LA4Sfyut6Rhkg6W
hUxmFbRFMyCIW5QjPqYIYhWarn3zlMq0z3nUgb/+HKLTJ1eCnsXkGYozNU8tua6e
pBNC/gr7EO6LTAelA0rcmm2DAZ9Sxswxc2ZgXgDd3k1FpoqDVZnsrmEcWImskY2A
b9J0KV5vVUsLfnLntBnbXMlkhk/tjVr+jUOHm8Vwf7z9agvIJcUZSPTMUKtjFxY0
PErJrHQhF82iWiX1e2FeTDudG44mvIaQohkcZqDvC9gt1ycaFJWWxj13PlYG+2Y3
41ZCYerp/L7a8va7b5Dk2Lz3D/3vTFgSAwaI1yxKIjrJFtzYo4aGusfRKY0rrCtC
n8NWX1ZAz7tAsEHfaimUUTomuASOPnprBnCztEG+n7DPR3WxyoLCxrO/vD/jy9Xf
ALEe3C1WgfbzrFpco7XCh56ce6qe6zfSY0811sfZ6q4/ZOsUdFpjQEXQ0qykZNmq
mwYeAWA9tOUsn5hwONU0Es/SpZsjTSaegJHNKbGN07NMHqyiGAj06ievpf16h3VX
3V+1c6U5mFfEt6IZeG+o4QVfqbdEmd4GrLhhCg4kLDFMEl6vtfXNfUEQ93HkxB1k
ecvhfMRGqzd7JJZiRO8w05e1nB4reR7HE9pXAkO7OsTz1jgZARyJc9oEkMlOQQCy
r7f6T5AXUzDGos520ij5l5K1kbnyjMeL+3Mwv50v2SQYy+29NstCdPr3JuTIHOq8
XzdE5dmGyvM82HE1k6+ECOWVCDjL300vZ6HGxt6w009XZlh/RvzKrfQWX7LVGc+j
mha9YcM+tpKhJSS0Kznztlfs8fXJae1hA07F7h83oMZYY40d7gehS+bwB2xxjlJt
gJN65JoUP722oysONwXxMl6NgL2KWi3rBFt3ZkdHAY7bsGwALpC6kTjTmGbXe0yu
tltsjeOhlxjf/oDIZltcELZ4i5FyNNUpW5oyTcgTA9tBRqr7Sdibi5kpXhXm+Yac
pjKVzpgNbQQwAPn5vNX4KMqgtNB5PCNh1Zxd2Qdf9/nZH/rsXwCLnlEl4JxC0Tk1
VzNcJra/R5TtHl45ZQ9gq+zDNP/c8P74RnbowKpWcjYMAI6gUapoo5HvJ1Uyqjqo
zIWizdOICoe8+bjAEhFbZjA18RWlBR9NY4cGe1Eb1iHcBMxoxRMI7wMtN3NyOcyz
+3/yvs3w7RItq2QZ+lUklYa9areNVPbyHP/hZWMVaD5BIguGNVfFqs6eT048AiAh
SG3m3I/lNfbo4io79FrckitTJqKbt8zFKTv7Gx0UAsSgzt9W+yB/lrBvYJD006Il
Xpjh+ze4EZV5q9iBQyaq+avD6wAicy1ixrIqLiHQP2hPn3HM3sLlttKSDFCHR9gT
ZukbuVfBxn7+rI1YF71Z/a/d5udLgehTGqh8EO06rDeIngSAeLhK/UEJVicHEy48
jYyvF20fpz14MmawYrVvJ2jjt2/YBAJfUqgbLeYmUEQTyYNbuiz8CM2mNibYYiXX
99tzKzKp+j70+v1MYnMSR0TcB290C1JavTxjFdHC0Tj0PcT5kGDz6xDaxw7mg1BN
p81ZVC3e35Sd+MNoTMFAUNiW4LdB8E+jYe2VAPYinbwWCS1MWoDjjMRSbleWAdzd
RIoOYx/d6ttMCBdZSNsn/CE7h+4STcuUvbsVzoJa/byXxExg9L0eWYP28khd6eqW
WxdeNNNmjSWcxELzRxg/jzYCEduQSViLK32yt37aKXSlj3u8YWsmTXnQEl+V7b/Z
XVTZZKuIs8j+585pGx9wM9XU7ry8GRrNyuroKYdRSNwi4Ru00wvE7fBWHbcKj0C1
WP6THt20iQ1HAXXff1J2GlHKdnNrpAltmE8yRQASpkHtMkoZuEWJdXa6IvTb2GT7
6H8cqr3Srz3v/UnDXVIyNXtPtN0fzHuvm3L0K+W30lDx9A6HXip4AHknlwLOG/LT
wXDfbGRjSI+bpoayCotElLKRvakJ1anNE5ch68KVZjMbnbrJOwacYJHHNSRecKQf
HGxtQScm7OPNJAZnhC/NrxBR50dSYYmMpyma03TQZDNHrCJDUcj8AM+NN7qmIuA9
4eKGqPciy1SoSpo3hVsKaGiNFG8WNroVBwhq7RkcWRiCJFBqEDGzklT4qw8ypxTG
ZwKmhjl7kYFyl9sXQyQJJwYDO8cw+3qfPda+L1bq+zn4SCx5aijafJDSODzrrAoP
mnHrvRfJH/b9n6lgj1ZeFU3txmozrIHQcl5HssSD87PNIS7C5TuiC/TIOan/D18l
deGWqak1QBKjPIFMuChL8Lv7MF07aPpWIEry94E3pZr2tBHT1a2TYk8kUzG4usdq
RidUNATjJTDHMdxMrHflM/DJMO64OCja589o2HYb59rqL4N4NRVdGS68uvEqiuWH
IeUZDOTP+MOWhQYjbrS07Xw69Ij2Jhamwj0MMIjvOx7LFNjKPVkVA/cjRJwUNWXX
mycWKXT1X5YGrZuVkrnEgyUj/73EebsqO2qzwS9onKBrjTlARo1jM32V4cqw0YGI
eeh3RdWztPU32703g0zOxgZhPORF8UZV6QD4vwON1Ih6oiSno28VQIf/T8u9My1F
jcwONj4GqTEbJWIAJx2i4FY5veQ3prcavJuNo+Z5uFnr3ysOpjc4IxKf4wkYTZzd
1moC4Vx8BSX2DmUAIfxUNpQVss39aSGPV7L/qkOVr5wkzKGViOl2kdYwCF7QY2kD
OFO70Cois91zxLB6PolWrZJPUwzEvFefypKCK4/IzKlDSHpUWwoe5NVS+XuNvqmD
kXOpVhmrT9eTrDl2q3fbTBbOgf35z9ilEFva4u4uTbMu2+0cgA6WgbJqrIRkxfS+
IOVQ4nmmOLbxx4YX7qWSn5tX+8/V/kmU4H2a1goskxImdqSX7asyUCkzk09slSCH
37htSMLjOVjzobMHs5hBLjhO801M28E+egaJh7TsRdgKlNG0VkL6zjiLr0LYjR++
3LP2PeJgpAtsuQqsuC6AquUtbwkPix7Jue8Hir7qR9gbZWhT1DUmPMS77iuXjixi
hRAVpXMO7SLQKm3vtDRii7TkW+cICiBbURB4v34v3+XGJurxiGCTb1V5ojSIvn9w
elEWF0QAcyEkzfzuthZFvrEaMAH8R0q7OWBcx049q348A/zzI7BMQkrvR1vCMMfo
z2fS380YzKVEHrhxCrcCSdrXEdV4/GpwVUOiGkVn88ltJhVFo0WcG9KpCFucGe54
bEJrFk0xZ1tlDTJmGFCnDtscedXSKPRRs6Jf4xq0zgiT3uceUHZGEUARkLYR/J84
EYkFgQOw0zuhUxrMy8pnEUYVZuhUQimuxSZF5iQpvEL+Yy2nL7iY4QXk2nZACNJE
y9sRxILqlRzds7hjLsja/fIKPRMlrWfBrIr8+BcZYOkvjJnG4rmdYaHV8r76x9EK
PN+hE1DyJOneYfmXBV2/w9NOreKjDPkrZ9A+UsO+23JivhiqFHDVVA0nHK2r5aAs
9bjJbM6galM3qrRWo94O2FrlO4vAaIPNgnCFZE2y7lFvUe4x7cGgIsaOi9g97I6N
dimCpzEd+UIHWhgPJ/Pp4D/WBBxKuaG2QdKqKJG14Zyqwb6FGB5Mp+mSh7+chPZH
gbYAxOHXh9SUfjaJfzWmCbMiyj3wtCaSbIrNJmXyEnmmm0nD71x4DBb//bN8FVlx
EMEnMfPhnFqtu/ZVEOFZft7HnzcNDAniCsWY17dtV0WSVaiNy0440UigE5S+mq2n
BoUrprGuit9sEjp+djHHzxmfVUN80LThK/ywIYSQUJNqSEgzPwRD+u9yNZltSzFv
ygitJp+gIdF1XKS2JjBvYzveQ9/yA5+j9rE4X+nUwLNL4U2FzgBJut9KGpQqXytG
gioNfYqErkZPJzfKfpr4ftROEldTf82Ua8I4Ue9AS1jbuDVa3N7NLotR0CFwAAxr
MsPal6Mh2ZeApMFUrotTEcn7viQNSz1Ujpas4DnvaEI+VaE1p/6TIvtu9v94If4T
YX7SqEiVYKXw7ZgdRzrXYbfIyHgLaaCEDLmLjdNtjVM/jMe3xseZAOmJ7PMMz2l5
PIOVQGiPf875EAEeDHr2+WigQOiJn4yR3HcOWJbRcQAzNEET1DLi+elDLmPbLrhc
VArbsKhKevUU0dK2wel8nu143de5KQiTzI02toDcjvJWiWNdIoibRzWSS7mZXaSf
hwbr8DMNiB7Z+/jgXDC7vYpHkQIe80LddMCBnsc39ca3Pjs5LzK9LJ/H/zzpFy1p
fVcpvpIRTiRA83ijRx3Z8k257u7DAjv3Qn1I6yiyMqLPyq3xXhij8zuhS+580bAB
Cxj+GsbJBu4sryYVVh99LQn+Ba4C1gUW4cKC/7CGr1GuByRzg6d8pJavix41r40z
C4taQg5PcOdGe0+HM9A0gRpMiWuidC4rli5M0rU0Z3OEV4/LvyGe0laEJ/N6QMCc
d9rUqj8wyegERgfRbbjDtrEcDsv8AC47/zCJxb/G04a/8hK2f5nffTLN2U9bEtU9
zVAkvzHjrCDKxAfh37XBy2FCaQVcvomzjZ7HfymzfJVtEcQLKWRkqZ/M3i6FZomn
qhgSWRQQFmCCzJiWkrNnsoIwLmV0Shtmh3o9TvXyTv7MqpDV0MWAjM3dxt9zv2lS
jPAvqcWhCRhJCcvCRQqs/Jc7WX7WHclHLGYFNzBaeaC7TokjXshIsi9cWFkO1yVI
vhKrQ8/QdSQYGTsdXRB7ZvzncRY8ETT3w8ObBPXPk16wYSzE3i3lwK1edx1WcJLO
zFT1i8xkDN3UH4a5eutSYTm8WrVxbC4SXqMGAqNc+6bqDsbL2/Lrkj9GbzRSFleK
Wzsc8ZzoQFaDhzH3/ErPLVrziQrNxBi3gW5Q+r/7MQCGX5U/r3FlSMF8P+ugGoeP
HqlAB9jQdXAV+XgC/oL78lhODeD1jseiLuiTKpMabE5A8ldh4iHasWuv/+PB6hxd
qhjjmpuSHLh5AAGyRvOLTLo8v2cCAGRlL4AcQL1YK8mDMoXcUP7L3IvtmfmP1pr4
Hs5NxfQ46CWdgBZWJPaG4L/lMCPtWD3VOELNCgtnJyrq2GuJ+n9hhCRUS2eSRT+A
4K9708WMgIZyLRdJz6T++Ue+NOdEeiOU+cvORV4gzxZN3Jkajm0M2F7hCYO7hEGk
yFbvsYWmhV6wQf5s7O0zb5Z7Xxr/2Pgs4EJ8kqZagpmeidIobDkVCRa0VwEw+fOg
sgCZTpK/H28sLoXMV8MRaPghcVorVW+lKZFc2IG+qbrB6xj2uTq2tEUtoxr/Hsd6
ZDSm7tYGzBFi03eFMI/Qtep0na5Dz7e3Z/RkWiQOox/b/eNvAJSXxtYOhw1MRJzv
zTaqXsrLEqh9m27ToOeMFtEsyShKTG2zd+Cgka0fP8uY0bWVWWaxfRjIfkPtcXf3
G20MwZ1BHQgzJu/dpd8DCBqucak5WhKB06qN6dJijPGBlS3dsypa1EuhUfNihZML
KOJArG/VncnD33QdYyaNAxN4xnthUMx+j/AUu1Iv0jKdUP/qssLggeP3wv4hPqhM
aZN3eYNK5zn5FScJbWoGWKZHG6mlXINJezGnOCmve2vLlcd56zYjlRIaBmR9StCp
cicAa2ZlFxMdt8NhtHX/g7n7X8yuzkTK6hBZlU+8XvceTuYthp7fBuGlxyp8kphi
hB1/2JB7Ii+VUBHU+cMWKTnqgjSSXcXJ65uC034JUZ5818qjqpcjEQb8rC2ffkWT
I0ZtPHo7FQBrNufJp5lsxTGFSVQEgSL5vHiYEHQVHrdBG+wyd1Vw3+LDH7f6OvYR
DBwT7TYRuAu5mG+aIOjko5VnQsqr5TuYS7bo5ws5H73acxdlDrKIVpnSfC7hKshb
TwDxjC335Bm3eE61iY7p2mryQFYF9tshlzPKnO2928sLHM0HGVSpMMTJN/wXBmav
NCeUL06PppJkP2OYlytbqgkt+29eyZ9d0BphC7+1UXGobENYCacGGZqPjSl/Qv/h
eFXukywfbswy/ZWGD9KWdUdqSR+vcHjkg4K8osoSpK6ApkBKIfn7FOfqaKWqtLmP
eJmVJL1ZYc8MOMoPbmBSWifM2HvziM4stR2wfbCA5vJGlVNguAvxDzJfcIi2o0SB
+PGCnMC7z3d65D9xH9dJWksv9YKUSKbO9pMBXXwWq2OUdm5WWOu/vindXXQ9NMcq
TiZRWDdDiy5Bz65b4WZ4aQbJ5cyw+XmMSMnszUF2EhdpCxaz1WHnDI/IFfz77zpz
S6impURqXWKsYKk1kF8OWqJUxI3uWTJUatHMLbz3Iqs62TV9cGAUDzqGny+99WfJ
960LsZmANDA1+5ylUWUBBF69xBTmnojUjX2+9b+S4gU4yp/eN/XBnWpowFW1CIM/
6yOLrHPYA9SqW9AOW6E552RduSoBE7Bwd40okq8i/7RlXAiDkDLOu7YEu9PMYiWr
y67tO3newhx1yq+1JyDWbRn/ccfG/5z2huRwchshrlHzn6W1CxF0bDpt7rVeTZTN
CZmtxUrY5fCAYmGP8xfvLNqkj2BH9GNK/eT2Vz0t4uDFgUmPIcShWmZyhlig0AI4
d3NmEp6e8AHriJ4Pg3ZC0dgONpHiIdIBRG/jx46UwJNPqYY+OAeI05tZv8VdhJuV
s/PLoEcFDGGCEpAaSJiITJ2kLZBFzasf5dtQOpW1iCmEAAEHvnM7XvfuiyxJg/X5
73QL30JeoYMl9VL0Lqd0coD2om0Lv0gPF0YmW7K25VXiv8l2l0xw8KqNseJqOYIH
2rKBiy9vSAXvgw8NgAKiRSv/VAEIVIO7WX7p6UanpKrLJ1j/Y5QxNjeRICZNfea5
avv0SYH6MMQacDP5hI6kRxiQ570M1F5MZs7bzVJp8ppDmIemgQ2AR8UcU4CICz0G
KZ7l8a8f+qYt+4mTw8E7NWiJKreCLx09V7vO4EhobkRKGP4cYVi6N11uc6lY0XmP
OiF/tHj7gVf8A4rKTYBs7BAaMn5YSZMIZ1uC3InZFkR8yu437r3sX5knLgqwlcp1
sjjfdfL9rIQp6SeRUyEsLu/B/s3m0csnAIdvk2AlwRVv5ezJzaKUyBS3CJvScsjn
PFNqvg4ADX2nX6eyLG3fEK2wJIyxYjvNQw1yJ8vo5Bk4a4KjEL5BnhaeHSoV27JP
n97zSNlcdHdxsu2lG81FlH1rFFxtMzIDfUkXgd9C1EC6nvftuywfLnSwmWiaxM0A
V0CA6oYoEvg9uTm75dOV3dPS6aWGyboczrHd1ZuDcUs0ygQr2rpI4/23coKGKfEw
Z1GtssKsMjWGJEFEQBzZob8I0W3lZkXoLj6JG8tXvv5VZaWgsQz4JOV5kJlAwpxi
SYGi6HBqQc+Ika/CW8GoQdzgmp0NVQVXJF/ot/NNdqZCz5vat74u+uZqQELhiKxF
QQv44nsKTQPwsiGL4WrdL7TubdzeseUsLU14ek29ubiZ+Yw+NyXq4H8aoS5qwDj5
NxYrUEiaQ8db9H8Wgins2MmKnbTRP/O+ll/Ch59Z9Z5NN7NW66qO6QhEcLA9PBm1
qr2NOo66RYUOHHtDcGdWfqBIeUPCA3yC06BWDrVqd82m5njir/aRGJVOYYQbh5pU
Lo+I6VHDT0PGm3HYKzMkK1oMg30DyrC+6OXSFe5OPww+zstmiya8ZtOjJFa4OCz6
W41g7Bo7buSSlPtF5FN0cozAJDXU2nvuIRtJSAK3SqwNn6YqDw/8gIKMzXZyf3KC
8/tJavnSlPLG+c8/LTlZxJQ6b7CiVvooZUOZ4m3xzmUGI4nVaHgDAgBWJMKL3FmH
E9qxw7R+hTsgmVf5Eu4+nBYmcrhSWLKpgNZjbYCCcbibRYGZtwcDUcWMroLG/dlj
Bh32tx8PhMYyWiwYNzhCrbTVKcvhB836XoO3KZ4RzAKrN92c6OMQBV+fvXil/UiN
ykiB4hBsZQz+9CO3oqDHxJ27etp2HWVoEj7yOmFx+6WhQ5t+fMdMP0285ArCwwxI
SlM6bWhzyprSvk4EVKnQKNeb/hq2HJ5/D79VA0zqGuUdys/uVxtFD0x1xKz2K/0R
AywKmrmRnW7bKKVsieD8lZnlf0qOW0xFlL9P8Wx8gxB8qNyd2X9JMqzWjwxWZNF/
pyJXIWa3QOQf77ATIpgWZ5vmP0AMxGicyXpjbp4I+Q4QbX26yiID9EAlhNN5Q4Id
B9sgAIDSWLkSKZ+USNiLYm+EFWS9jNWPKm6+wDEUfl4/FpyQwmkiQZupCeHBRMNs
IwUnFyxGJD5QRhVS5ZEJG4nK7j8rdKZHifmSBkxh6ffH//OxVaBxSIkOo3yu/9O4
s8u2vJZgT6Y9kToOQabRvYerqSCKMdI/ABjpZ1jWm/Ptec9gs/G5rSOOXxPmppsH
SdMCnHuVI0oUOHY6O0iY3sQO2LVWrd1RQ6jdGjuFJ8WSWAuQ8ygQ6aCce5Mk11zA
I45m1D2MpbHtoE89OQ1h/AVtlpIw4znmUZuqsEVoNfIXIsm06iYedvtR+mPMWMZ6
UFdwebPS/By6GkJBX35c4Zr7RUjU8ymxJ21jt+twXxNQtIYOtHmkKrKQ9EbE5zh9
ETcBeZ0BSibmT50U249rUS+MGlSj3nT+3LjDC/aiImNsff+1fMRQTqA2XPo8iqK4
hCDauw4nvOFAD8AcdpJAXovvZNWjZ4qMcCPOCkr5Uk5D3zxYK5KOFCjWNQMFAQvh
YvHXa5d1+DE/dBwde1FR4+PrrYGoKIS9CMbEt6LGXI6TWI+0RBpNLdhgEsX9A3LA
gWa7/RPfJOJPzl0WuEdR4G+VXGQ/BSUKXwl3AedSbSSvICxZMHjKFn2zRTKV1/Ln
oF6VIvhLWUaG2NZIxYKlWgHdtkxCNNdL1EJ79FJHRqeqyHGoqcycY7yV24YHISJx
3e1AaatmD5VmAkebDCW7T8In6n429n2SyaZhVUNVfJBUmATp56FOU/j0BV+E8QfV
uRA0cslSiaOQhK0ePqXauEExj+MMaylkq1R9VzMFD3FfUAG6SIL5qmczoFMVjmis
mjXy1ukWoctVj1ZgarxklZh270SyOqGvREC7HBJFC5leurSkcT2IrM3Hqy57gE3Z
GzVqhqoa8lzOuL9qsTwgksP5KOpmmZGZ8spC9KrAt5inNErnTEiHVYrc95sovVLn
9iMxHyN4Lah99mNPI3u28Etypu+RDnxE2kKdRLS04b3j3U/u/WhxQCfFJ6SdwuST
TfBc8fONCAxBHIe2YsNN0wU49llQ7v1YF2V352A1WIFGlXHabagnDjOluflxBZCJ
Sumj1fz+lVwFoWqxB1PLisMymkURoGMdzxxmF4EFYumOKv1Z6KEFOtN3TOQIYY+b
6qmho99ih9DCnh68Ix8/e3y+MYT6Wup2Je3ewVBzpfkgdL7QCwQiSAlQ+bQW842o
/FQE6a2CCCH/GD73RkK6Rd4nKzC1r7Kv+IrjDQLzxzXQGYNgeoqOkrP0vSBVkQOV
qel5xNWJsvDynVc3KimvydVoP0RMTq7v8V3tnaYdJk+FVzi5fGM5eqzS/fRs7j5o
5Pn0nP5EPCj/cJ404PlPicbU0aqb6PugooyWkJyTkXZlxOckBjkCbXpuy0tEoX8k
tUlKXCz9YFpg9OC/dwmhQXGqF05n5leWwLbGyMgiOjuYN2VnuZvzJ9mC63uAivuR
aZwaheYo/ZRc2DmmJYEJkiiBowiDfYQ+EC6jejbrvd80Ml5/7yadHlnTUoWZfCGK
GOQqeYS5NtxvNFEJ/O5etyG4weUsHy0q5HNpqFYTRGR+6/szetNuqf8FR2cPiGFe
YVtShXCnI/TKCTfDylKGe6Bki300BlmnGNwi67C+uhV7CQNnhRAfnOAFJBpHfZFC
v5NjAdIepQojm/S2aNFzHPSB+h2Uz5kLGDQusw7Px+bD578J8S4pKVCjyXtjho98
ddLduIJUBAlL5sLzgFvHCrWL+X2uBQG68F4OT0oNRKgs3tSMnZR9r/XHVrKLukab
sPOwlTrO/P+rP1Ro2aTJxNc8OTTPoWzN8HktWTodPNpK24tiMCuDtH6atUG3O6/e
GLK2noqpEO7uRp20Jj4Gva9kF9rQ4SSmwx9F4SQwXIn+SIgNvt4Ekfh5QAiQbg/T
KgT9XurOmnjDaKYI14fXWL+S3WXnS1PtbiHNTP6QX+h7yXzz8L7XiZRqP6LnyODk
J/XEvDDwgZXk8tw6HCBxlNQy0iucMyGuDXE0TBzCYHSw39bcPwjmCwkGxtSSTsyl
+yTGO/PDCHiIMqY8SMeIDPT7AtyK3NXjhEYPN7EDmoNaLJGZQyZQ7R/9bq/KMjbE
ZWzKoxCMYgJ88R402OXAyrzzNuQLSRetpkiEiVj/J6Vu0XgreXTlnoj9Zx5wR9Hl
zE1bTrBRM2ZkMuFCQofy56BIxqHoIt5tHHXR/ywQsUcMmejqyZDhdaB5WYdD8cvh
CCxazr2kpZo+B6Ba5Rg50o2GzFFVKR91RZs/iIgReQp6mBrSf7sU//38qq0QMVne
yZI8hXz4JlKpjxMzrL8bFyXuNBtGkXCa0UaJmlKA8hNuaxzRaQ+BP0ndPfgr7Zdk
zYFFTkeduIN3I63Ajcxsn/i+OQVydM5JZI+EMFpXWrCc9LGsSmu348T5ptOQZXUs
tcswXPk3aG0Zbos5/oQ9aLIT2JIwKZNVeTLupoX3B7bBvHkoX/CJTAhsrl2A+Bbc
5xYf+fLrGGSIsasPl12alHqTFq/aNoPyQVkU2zbQCzYvvHFmF/xbvC888jHMW42C
xsy4dzvpPNGv+3ZBzMdMaUe6Mc3/0eB7oyl/337rbD/xSCUYSIIXH338zEuvOOGR
Dor27wEFnORAQl8EzHOgZ7nFumg50fb20BbvrUW6xgG7qljxnzORKgY8o/Hf+n1B
2rbHdGZztXFfPeqMOzQ0IHyRiX8osqoAGnRxkT95HU11j0e6PTK+/92/lDmPrWBb
YuX8txH94gY84XlDF5H0VbBmL7VZLLIC7F+KmKn/V7dO1IISmXbs7+oD/pdhL//5
HK0flARns5I5AYHrAtMuLOl7kpBGccb3GP4Q7M5iNhGMPJ+RDnmOWgmB842B1gE4
AurSdkPUprs2L+mw3X+IQfGA5f3lKKwu7kVuXbTwgXjj/CNXtpwsZwXXyOZYbzBS
YQ5CICMirNEVVgyhyviLxk5YuwKz7KahRSvGVIl9JRtwFec5mJBMUUo6ntLJdFwA
t/OL2PdzSB49RhNQPjNHDGoTg4dVINFkkKIU1tG4jhl+ACHxA3Pt9AJmxUS+RaKn
Hy3RN/b0HU5NJfEPac2E7gdqqWoHsbRES247wHyQuOQkYX0dESCNEM41kb6jWF2F
qyt0DE0ZP+pUmrKM7Gz1RXl3ssk905CX2qSEPfu/fMMTBc1Aypdsu17bSmtdzbR6
U4yWocORldkjTVHh1AO3L9nFXwQ1J5rUYOGSS7JZYdZlgAtJMJphS8BsswqBcDm+
uhpgvQJNg34mmMs/bj7qYmZ34VXK/6OBLNl1CugXvXlgTBHGFGRFma8CTwM9me29
z9Ghvjf/x95z5uTraGOAWDfBd2nQxihsqVZ0Wv0Y53e0rsCqh9misZ4G6RX/NX28
VDtRR7p2X5OLz3BSP9Eu01Pk4/xY6bWqjzmrQUl29kaBpT3SAKKDQRqEF0nNiAoR
HalXzfQOYrgp5lJJzxiieM0yb6f/iwDk/6rq94/69I3+7amJwneYlACPOAuO6TID
ZesFRn5L9aJmd3dXmoxoKi8kV4EhhSJMk4phb4qVcKBsDTGoxB0ZCd4mo335gvfy
dXtOF5HM4hpUzW+AHA4Ei6H2SOPWnwIv42BzUgMkf2Y+bN8zSlZBoqdZzHAFAm/3
3nkoaqyweEBVjNeObTyIPrz2scaAeA0RKdSDiPHRtMlCWXL/BDThO4dufCoXJML0
QKroLHPwJqyYryTrKOnEiaJh9/1eYyn8uGfIoWrOCUhgj8QAHjBBhQN27G99+rS8
p+rF8fbl955VM86926LsLGJWdccuGKjl4rLoNi+A0DARHFXA5LBsW/l0A9dbu1/l
2iMIBbmvui2/DIbU6hSH8BZgnyF3qhdCYEB/yhLftDd5AIntP0Nm4kmH8iCp+42T
LbJyzfdExo9TGBtsOEnU7ZXZltVts6rSUpgITr47J3z5AEI6jK7llAya/lYMPgCo
nUweX5tDqrRuxg/80vHh0/UOshG5GKNpENdnQUf84fVZm3XFm//8Gaa6UK1BAd0U
1gDF4CUl2KAxa0sKZP3tjMp0ETgVc8N6OdofNiNFIOzFeOx5o1Q8MEhf58WwVvja
sWrhl8dN94R5+ckYkb25az2rrM/x6JtVBdbcR+O+2A8ucE08j/gL9irJaEtW1CLS
nNxXpUN/BeWnHHezXMkm7fyHrMZE/bn0GGXdlOa4BrOrQi5Hbu1bQxVXhDL/U7Zi
PzJJ255C77xdVEdL6p8Cmz3cocRUIiPqAcp9oeFXu99gQlkBB5OXSeiNxZBhFhwo
S1eBfmbO4UwlEi98IZ+UAuczDhizcZacxSOvtrKqKv4UPjDjkk19Wu7H9LP7hiee
upVW+KxY8ZeqC3jQ3r+yj0ka4b3y2F+7rBYSSjdlsMUl0UIEx7IrbQEvd2jr+lAC
Fp1912IATSNOpWbgjEdmFLZ+7InvidyEb3sWnvrljCkM1IHnbPq5bA9mo73Q5nl+
9xzlrZkmLZdKjhREu9PTBFSHguyZFKqwj5pnY23fH3FOO+8uf8Z/xBUxyRBomT3f
yLNCURKKArxeQNYwIe1Tnv+T1aj+JHDMnRW9a8O5agLsE7esQZNxqIdJOSqvDYw9
WZA4ccZLZKuh//uhmvWWqNP77rf3M9SJprjftZXxkLwxYyD+ep7ObdKVFsi3b7pV
ftmy3+rBlmAhPLO4NPNiX0rcIvo0bzcPiahYpxz2J/wm4pw1nIVDcpm/G5WkN+S+
rLejAFhKhv8egT6/NnS64S60TqipQt5D8d8u0Z5qB2gzCwlirGJ11KDri4EO3f7V
ohFBuDKQTpAsZuLeHRxAm/K9M8GzTJxR4nmkF3xNzWVxGTsxM8UzQRjt6pBXIuST
Bjl9Yue4BCV0gc5RrQns0kDY17K24yPsVUX94/sZR7mxkFYEj8S5mWHU8hnNCiKr
Ss+9WwKdf6Hvmc58NjQEeBVtj1WVUuWY+UUX4T4ufhRK93OovZRbpDq23vl+W+9Z
A5MSg80kcAXKKwWRUNlYe7JS1tdcHkMyWkIY1FhfIm3/YUFbxEoTOPpvhdI1JsOA
KMS7kmB0CxNB/s8HLC8CSdJyznsG/K+uPmHo5j/vwl2gTyi4mNzhCYhx52l4ZPH4
xRdWIiaeSwJqZfSw+cR4qBjlCH12WYXBq96we1egQrNvCErp6Mvxpyf4h2AwkvqY
Pj6hiIkDtBr+CeLGirTPQi0sgMyRc7zmOEcjTa3CmuJKxkERzNvxWFrdRqEA/Q0T
5E8NSVuF3LxYe0uPWDEUpU63DUJOK78GiP5lJhuc8DWfyrr+5t9VK6Djo7WMG9FE
bwKDW+7nhW8gMuMngAl8IouwUc8c6rRS8LD6aQXyH3Gpsew+Ht2FEpCOvCM/JcU8
geGqCPDDklCUnDIi+NiRR8g9cojyrKVsocsba9UjFmZ4bFwFckrY1p8YmZ83Pv8x
dsTQvIcnFQNYhbCGTOGHiMN7oltzbAwAL9l47FjMB2wCSJZ/eqX2sNnOsGO7Stwb
MA26/zmX6OrNANksaLHrSugIr601qCZl8tHfyrQuXnqcBuFW8KnQn2ye9fPWsnJL
vpVlzK/4yrdqiosC+ww9A2IYds1c1X2MJAjlt9obdfZjq0aEEF13mKVUS56nQSr5
+pBrHPMbrd5WCFWtKMKvua8fll0G7k6ZKYbwt7ccMT0H4H+UsrOwznGbAlZ7OB3u
sD8u7SfnNdZB2xOGEqnOtL8b8ERFXjbHmW0ux6+UYOugf/H7n5Jy4NvDutRNdspc
BZZc3Co8TrCO1KdzXhI7sBEybu9v1RLjR7IRRKJmZNLbKQ90hrekymuF6PGSaVge
XvDDr8lHC85vXBWW91uHJz+IE8bTYP8iG6xNlh2YpTjRcAy9KC3MKHkVhpr95uPj
U/4fyyJjAd+0ga2rPc5Hvimp6PKn0vGHEfX5SGuYS5BaedHu1HxKkti4gRm2NP48
eQo8mQBrLEsDiG/MZA2QBF21uZgdoApsueJ900nL1dtX4krrcTB9MktpS0GsI10E
cHLUvLYE2A7SLFeo6Ek4uddixI1liVzjr0pFYpsr1Pj4O44TzlEckH0RIuoKB3Hi
98KYlSAdBHDuFvx61vnzqr+JYUCOq/ltMJ3rVlPvKz7DhAnJ0sFq/QGOoGlgXYQs
PO1tkIA5YT+G7CWD5UxxnYedIZju0WD+/JR1rsgjK66addZMhuqchsJ7iKCeVeyR
8UHESLrDqU9L+/3oJRJzNNuH4SjhoYz/igf763rPXml8zJNoA6NlYO1KFC5ieKth
APfQtDgj3qrW8uVw3a6/G9mbqVb0VKqibbhmJzyM/r/eBHVWUAG5KPdPbFxOFP5R
T+FfAwgel/D1bh9y+OeTPkHhuqdxwM2ubnWcB1kzppdEsrORO9ha981eSNUSqoHU
Y++63Joy6UBpiohaDzVRpG9my9s6y0li94ZpGBm0JfMKeWLjZTpm5xyIkZQsyCvQ
RkCTTCzQmnsEoEYtU22Zc7SqCpWVt/0tEzDqLG+hWbTG3KaIFf/xDFc+/+apRdVT
Pb3zoWidThvd+x9szM1mmbtDjqSbgxTL3T35mUcOkRyWiSNpMbUDQ7TxdKXYbwyn
LsIyRcuBGA2eNEAJZftoD7DJonYnj/tqhTXAD/LNxLg6K/XKVG6p5NregyQeLphp
7U/5BPoiA+MxAylgofx901XBVk44f1+k8HLj0UFbeKDXXg0nOVjmi4+y1IwqA1P0
tdDApjYFv6/tJX63hjA//hFoperEbBHEx1jCwRpW1pjLBZ3HquO+F4acC0+us6Zu
RAEUMcDHEKZOouESTGX/TabGkCFSDxGn8yLpgi7lBK3QCxSKz7pz/NLUxyrkH64e
tvtGuOYcpYrbRm4vk/koI19gcLwjxZ78IDIQ83Sfagk2qTRvhvH/3hZAk6NM9uEK
HS3e5vMrBt8tQJ9ozDiKUTNhH7PycxmGGl96a5fXP/lMjcI0Gh9enRi0tTyiZxYW
AcmqmA3FQHywi2OhIaYFRR4HSFvh5NDoJBfE/M9ATcb6vNiMGLxgdjFjC1d9nWXB
mFCWEAkaVC+nSwuTSEsk4R+E5urq2xls1W27n9GqpDlahrlCAhdL5eZpaLg9sey/
u2VYmyzYVrtW90sTmd2OUs3raHgT0EhB/uXRK7rFg+QfXrBg2IZhX7ElJLWxaT3J
+5b2D2+g7CKU1McPE6GiWTOJObFCPNtDLoPceEOJa8Me911+yTFa8uvY7anWhcpB
aNQlx6DYl2IwGivRYY/PpKRAQp/nzUne9mUsps4lkoAsK+L38MjxLwcjM0py1WUC
gZWHvcmtj1MArQ++D8Bj+7rqZCDn87lRc6RbUsDcSGyN6VmUyBawnYPFnY2QKQJ6
R9TjzLn5M3U/WP7ax4tH9QsUF4C+56rEl2FW8XCgrwn6upvslI9qCkIjmVqoXREd
X+jVjBAiXHTkbqzKOp0BFGZCnE5mOTcqQcx8EJ6UDM7WINFj2jBw9SiHMUcChvqZ
fff8mtb6am07gNYq1Tc4VExcn3grOQYhE+D88HWIKbMHGv16zLl/Vs/PUYebgEFG
rpGr8jKjWOdk+8066aniQLwg41EPK+SFQqK1D5ay3tSbePgjhwgUFD6aBiFuL/VP
Etog+44FP6vu1+L61P5gJIo8nak94Vs0g/H6CD1SdlNwSKCECY2ESKn6/amoU3Pp
2zylNjnxeG/pYAftFbXRioTEEQUIEnz/woKTjbQ3GOYGf8aIH61MU+gt1keAHyGb
j8i4kJ1BYfTBG2Yhn7u+bfwAZVHXhSZVmXx45hIFgs3G1ljoFOSPbf2StOLwKgaL
9zkfZuEmdSQXD7lFCVrjv3SLqNjxelFSP6K291nWP6Zwgxpqb+ViI/RsyfS5YGjV
mqJuUmW7aU6jboxKKuFNnUpAKc5iUMQH1n46BdTjyoS+CWq4BrDkJDnUd2wkBZuV
Okyu+3G4xFjviRFnIrD+jDYr444j+uySdPJ7UjC4299ySWQ5oyfdpKd9w8fx7PbI
nACSe95eeBPNBQYnAjcn4A1lEvJ4ZguvFRcLlPYoSWxKbczNYlCzc3JHvF48dRks
rByQfTE6R8x5Ghi9RoVrhhdmweEEAz+zlhz+D3FK2pYXt6s0DxlwuYnP4vPDvxqO
MsjxwHnjDAEwKrUPjR/pvRoZ6r6/DO9iN/+exIBp+dS6INTXOnTXzviMFHTGcNY0
HubQtB/WN/3ucY+rdxMXaxPW1s6aSuWC8Q60dOQJha+/CmCOA4UPcA3Am/8h5+29
SnUjki95VrPlC+NvEmO4J+inH1rZRoCCNw/hjX0T6GX/pfHoj4eymaQmdRXF+LPC
/7rwBGrLoIpqCNnrUII3xP3Ftiynu+Xo2rlXbRBPQrAghwmYXVwbuxMfumSX28z/
yw36DIh5vD3hrfat1wU5FJ0gRQckyno4vPILO7t42UluR6rtkgsbyv6Jk/LGAeGT
r/AVOYcYkmhrOZh37Dx3LNAjBvfYVLcmCQnqvc7l9IzfwKoOrBSLBEz/Z/1/2Xg4
yqIQFF98LX8GR9cyvgyge2gZ++WH6ieV2gZpeh6CrhZhvkRlR1SFCpUjrzls6hX5
5s8F+/sqnsIDIln9s+CwzBKsClHz8ycD4VxOx5XsHn43ZmYxENPk+VQb4das06SI
FA+EMFmACr7WZEl4GK8116mtAKJOI7Ai1LAPmV5zA3g=
`protect end_protected