`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1744 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
BD0Uso4m3HP4S9U6YYcCvZ1t1QHw5Ulm1VC10/sO9Eeg3o7OLsIC89tbJ5x5zbjU
a6PqdPTRx5RWyZp/5hDoUeCVprd6Thp866kljw9NUz+Jt0cPjIyoFiAc2Ao5c0Rd
lFGerWKbVpHOc7+O8uaqGtmR8RrJYbGB3gD+q1qWbKFg9+7r5q5aYM2l68Y317BB
E451Hy2RDoiZBFxVTxqCVSU82umcbUYdoP6lMge+LuY/K+dVo+pn4GZG8owxm2ua
+TQt78a8PHkAI1l0/f1IHGcOGp41HG/CkYFJAZ60L6yt96m4SGOstBNPL4l3xaeM
JslqiWBw0UOl/csGGOR+HN8Ik3U7thsW6M0FPjvOJgPRJfQsS8/TK96NsgtlzGp8
zCZqhpkmVFvqxytoZEN8cs7nMcxV6XbnrV1r/GVRAGFd4I+jSaZhsqLUL8UjN+oO
1QYRwJbUz4x48YucwtAEBbvn//y1ktD+UuoCRYA2K9MEKBxOsFMdcZ8qzYTKwiDh
48YDnDC+D34acDycuQYhfsuTZuCuaVBLXaxxjLqPwSW2SEMBpjBIPSD8jKNpWKFY
XYKF3aokdnfcdhB2SQG3/GbhfhwuhKmOt5MLgQf97/Qc7kRfwRg7G3r4zEGhKyUx
LnMx0iVr3E+wJqqleRybezeo9TWFpC5FC6iKH5suFNgJEHdYJGaveMlQFOO5BFXw
miPN4ajhp0hdTso2Klxv7ElnXnK2aTGrkXsscIXypi6MD6pY6OedutzMNaXZnAPc
kOwyqva4rzPzVYzqI0AH+I2iqsTGud0xy94kkFS/hkRUaDq8ZJEn4kEH7HCqRrK8
7ya1Nnnkizx7m3055HAr6haiT3Z8QNRVxNBRNl38gVIOQPFhcpS/JibUPABBo6t9
znKoCZ/ENCK2swkXAeWByS8T48Cl/sFiTYMJh24r+tK225evrr4UTB1h5o0MKqsK
6f50urHxcqM+SJ89mC1bQPNJorYIy+nwIryyXh5vQsPUqqbWLV65Z75QWFQhyT9L
+4F/OVH/j6Y/qis91OAFWjkZD6Yk6UzTd4MKV83dCsxu8RpNOHUsK1Y2Pk7a49vo
sFcchyKfRybrxfiSKC6oCsm3p5zIN7JZ8lUZpJu34SnHr7Yce0+c5DasQHM8Qo4R
Ohx052bmKy2DOPdcY696gCXjpL+/QwxKRd/YFmXi/jCmLuJH3e6q6I67LxwVGUCU
aGbnLorBSjAgSMM9s6BjWg3w29EC8YbXYr43xYde53Di6jsikFHP6+2VetwWn2Tw
YB9rFpdrpubjD3LqICcu/VyaJ6q7XveftpnVL050N0zv7FUy2gpCUTU1e+ROpBGo
Z4N/1hfzNOdOgBp9d48aj/v2t96ou/qyi60T2yDD38m5FC0DLWsqzWbTQQT15M4H
Z87os98+sYRM3QTdq5wW3jL8evjoZIO4XoR7nv3NPHDzXWEyB6pqlfybqCHHLWfW
/wpgtbrxaZTRGKZfLrGe0uXV4MXtksnkd0C0hotJXr7gF2Gre2I2eA9fnpoL8vgt
x0933j5eynWnUAThAL9OJ6sL/4xwfBeqxCmuM4TmbWUinbc+vPPl4PR786daFxpz
7hGxy4zn1N2V0vbfgpOjvJ4XJpgdBRvs4hn5CYRfyUYqtUaKnM25cP6vcu2zD192
hmU8WGJ0Brc48s4a0Gju4CmGI/CIKJdSIcy1D3AOCoe8pNk57aaB+pXUUvKTOFxH
ykjLpoqzU92JCTmfZz2P3bSORiUpKpuontrMYC+ZFK4YtCntUvOkrVnPciqqpZd0
c62gSIBZ4P3oCotBeLj6jn0lqG2woTc1YgPqCIktv9muRmUofCm7q+A6mUKY3TRC
1SbVZrF8jN69HTaig3HGmvafWd9anGIXG2cIsPz1c5HDer3vomcWwtc0SyzSJHgf
3DOw8v0IaUxm5+Ol0gN28cwYQz1UwBKHAgJzcVlQvQd9xUa6cLsPiUROo4fdBTrb
R9rD7P0JxvtuWlAmwST4PtGcpjKDzVhWHpxaVk2P54kN7gwwCC0LFLqarCjqoXlQ
E8D8OGg/GPHjxmp4Pbd6duiZc3k8S+ATyp8QFBcF0KYwdEe34pTSG+accFU4E5jV
4GumCCbtpL4DJfHyEewgJ7J83dQA8i3Gy1vxBgubyniPUC1zVaS+PjeHw3hG3MlZ
kCCWknWHkAyQuRyckyK5IQ==
`protect end_protected