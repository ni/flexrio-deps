`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4320 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
/vEkqJfyK/81z5lf9X8oFX0gGUErK4NkzKp+wSHlyAyYhErhFejxzkc+tmbNpwzk
gqzWnspf7D2Q5vBzurpcwWcLabCsnu0fL15puoXp7H75bOHljiMmx3LHwKxGQsti
UoPrEdG05eE5RXydS+amByUBead8aBJ5WdKynjpN4X33yCt+GsUM3Bx1wBtBJPwY
fWkXwcejZpOrIvilLXj4e4rHU1KfLrVJIVfbMEMMS3II1g22fwf//pTTyFn+J4vj
2Lx+OBV3fql2BWFK23LSgprpk7kLjx9kLTSarVV3Q/6f+HXLgezjPV7SXUYAVtVv
nS35kK3OxFcrFGpP2ERNZPa0/jWc0sYXkvhyTLNa9DctInINIRlwFMIc1qGfizdu
JqZHdzBMR2kcJVbjGvrg6S1XJzG3fzC0HwngkwrmeuWcBXXqvvnkxnz2MSH58AV1
cCR5/A9dMV3GbHzPMZxtKJoUqpecwoJYH1NW95CXo4HcS+My+E4MZW+0ccCygp77
/aaVmyboeLRupddeLs7cI9g+mjWi859vLZRQ1bATzinEWDL4DAMSYJoKdZvaW2Td
95Ng/U5mDP0QxtslWXFb9JNeZtlAdIQuTHZvZPgza/w82IMRzYC+jAXGT9G/uyiM
Mt8iYCjVak9UeFkxKphZUybpRLTixA2xEZsmZBWEOxMgHxJ38E0hS3eog6jjpvM1
/HkIkrm9/r4aIikiSu4L7TB9LFPYkdI96ufvpufT0Hd/UnMvvDx9FLDyIN/jgy0Z
RgGpW+Ct36ETGVgbg8G30uZ3g8cg0/jHH/c9/ygXAJgLJRytDAyoyFxLM2jNPj7+
NaL19MJlpmO17fHs0cpItuzGwmV8+jhIF3Jx6q/G/k9POnFtKE3BUGl6ydq6i1Zp
P9BlDbp0TfSayLsOYZfPLJxrUVrLa8Upg6YgxUGvfjsLYWrq9DcBXC5Pc18eYEWD
qy7e9Nuli54JnCCReeLBGULHPDiarGx7d8XnTpyrYyqYUxbY409kJNf0bmwftgsV
tG01vb3MkqANG4gp5AO3vYpXOmYnO6/NgFtczIKPDRdbnQcvuT5r43LmQwzKraiO
ZGYhLm+PLrz53a+xuaKgeDrUYT5Z6O8cijnWElBhJbfBVgefdb6LwNgDMlUjBAfN
lAH5wGIsekeDFG3kLm7LmZ8D0Jsaqnteh2iKlvo6T/7ayABhutLsM0KJa/jDoJBd
O3IMvu9t1XKEDm/m0mXE9Gyanhg+Imkqpog48gSv9vc7v/4ysokb7pF9UHWMmT1W
LywKbjS1zbIB7HN3myCqLPML6YTrhMG7zbkGMovS3X3QOyl/ZM6j7eltN8oZjjqI
0HRcgSF7fSWC4r03H3oAdxvWQnyk2377NaP61Gi0h5RWXZM5Un6sv2gxzgYSCBLe
pVV4qTK8JgLa6Vh/uH6VxmQfiiYNFtsFi7iwA2Bbc7ZrxxlEHP5LGKYPJFwdC8pf
F7nM6G4iLvv+SGaPlLjnlvewey9yuo303om4bKWxDKlfoPEuVzw2ZNEUw77PQ55G
zURbQbgI8LUQLpLpKajk8YedvVeJFRbY5GMCyMB9ES8RBX6dB97wgWF/9tzkFFVw
p4fLPNRFY06/YoqKcyf/cX2wcnfWOsYSb9LooLaSKmWD71lrZM0+M/Bt5cudGaGl
ci7z73t1uSIET84Lv1UGgwU6Jb6ZaE0L3G7SKDyakd+2o/uLIvYkGIt3wmj4E+tY
c/YWex7XhpgVW7FLlJQyiPUe4EiZrSifBrGhCGpWkPrVMZxr/1CygxuDPxWMOqNL
++dcc6Kbmcuwkb1BtHjBYLWhYaI2t6RWAkfofSrpRhOcAnSWOX3VNYI8+Rwr7JQP
yXxkCUGfu7yvn/Tx4K0NEHdVtQ03kYNvuY9yFGKkf3HPehTou0g6kauO67ML//vG
3WCMtcT44ZQBwxlRVtGB6OHE/uPkqxX8IT+tbs7OLsBzqk6pRw41QBN90PV5L7nK
LUFT6F0czemWecx1wk/0yhJo73Ykus+ugP8pVh4vbXF6WW1CGvJGCHS3Nekfb5o9
+akVbb4VJzl8uB12ZyX87kCzJ18ajhO5lSU4jLt8FRJvOBW/ABMY2YScfELrCySr
+cpokH4EfOwQba//h8sklNXbxQpI2V0O2C0zEnTNWUIeVFKrhRFd+76CwEd63t0H
nGRdsJzje6rDs+uW4abf8ZpGtfDFvdSvQNOO8uDIf3/mi+ZHxfg9oYn7j2ol/oLZ
ZPclXCvBt83IRblnaD0y9BqoNzUfTEcQ5G3rIBuEiGi5Thu6mcWDXiOAY/iWH3G/
3gyTcBsutRpZwBee2n9rnQ+WVe0BylgaclOztvlVRIMZjYzIz5nV0p1feJcuwLSN
MFCa+YHfqEU3SL2b6/uRJJwBX3McoMxYHJa3kbb+MIzAFzJqB3SY5GS4DFjyRcDQ
flJThLLgRSxUBf6yFzF6rPEamehOMy6G3L6YTGfNRAPxzKj6YDp6q+LfcMsrqZUI
RCr4Dmlhb82ZbJWnRMa/zzBrJxqt5dj5lqOX9entlZP6wJ6aZ9vMTYOnHVA+m5Ro
vWUrgQxtcl149iQ1NkSWMDs+5n+M+mtc84MPIIi9ty48zH0Jn5zqnt57h6cAGbZf
P3CzBoW/I0pyq3n1gsa1pjx3m6xSpuW2XnKr/j8B1sGiey6cQ5faQlYrjEAH07p2
yk/8DaqAWjhETUXknEiBmpVZYOgk3u1QXb7W21WqQuwm5xpQ8PD/SpNtrKt2OKSD
pmXL7ez1Ob2AFj7jTbLdGkRIAvrJbXg8eLGaFOodlyrJC9BgLpcW/ZoGo0kY078v
NsfT6+jzZsXZEs5STdnvDzTa9PZmzEGBp81eaneoaGPTpbQZZCDg+Z2ijRGvLmOJ
hWWnGIChonmHXkwajr5D6E2Vvleoq71onhAj7rJH6gL58ZHBY5unRbriPRjyeROk
SPmcL+s6LbKmFyy4nLLP2pBy9ZZCkWUUyjxs9CUj9OX1ZbPfENwXKcyGeeHKcY2K
bwbQRCGvjA40cw+0BadmhAgZsO80/TlAzKKQHlhCxATHF3l28RWpj2j2HmapKT0G
/zTwzH780YvEIIDlCd+47hFfn1iao/0/3+TOEydcVbYl9Udw9INJdgiDFxkwi0Ui
YwNVABy9U3tIlNXIkV/t2394h5QDwz/zqX1qLXd9J3QcmhjSvBBj9Ro10WVV+ET8
+CJWk7mOVteRvK6BjxB3jwaxUTDoBVAEY+tKKpLnMZwunljnfs5bn3cdXuRCGxsd
RRCR7t5meNkIGDqFul0/n7f50p1ta2bX5Rs0++L4XZajHG1MPHFBqu8IlfBja3vO
bC9vMqWgu/hpl32Kx2MhogzP6gdXmrw6c9Fryq8GhOIhsiVx2xJXoBma+QSY63Hb
ToUBDr6LJyjaVsyAVjfWZKMyxAsCdL7V5EHb1qC8v7lGBgdmeaJXWAlp7gsufuuu
nC6VEPsmU+AA/l6ZqoCNtMt9H38ZSuNlhElfXPv+Ym8GV2kYtO/hnM7mV2LDL4X7
hYSdwWbYYVmTbvnrmHpJA24mQQk3tgx9AZDw9uYzKmrBs74TcuAXKDL6k1cN5TFv
ZRyrtFNCpRJN2au6HkZwqVYJtmhneuJDGRQYMhFsggrnfsVBgC+IF3pgeQNcbTIL
vMi4EnVJc9zt5u+LW48GqPBAi7EKpUIbOM+43hguSIXupGoagv1Z2QBiTRjvRx51
YEr3Q1CrS7xtxv667gihSRu3Yimka1tU+Q43NVc6wEy7Jss6imlUlQ+nDXi4fUxX
0d8o0c3xN/F6e2PkIIOkhzNr2XWaVeUUWdsitf6zzvvaFXI8S0hgE/aN8Hr0MAZj
mFmuERjBLOPCdPJvvLrDL02EOFYjRtUwY3YtXmP9OhX1kc+uO6BMRPNJy9y9Qkw7
Kk7q0YOrWHDHComCK/D2So8YRFDy0PDEONzxG6oUc/Nq9O/sLrtBuPoYJEEpuikj
0g1YyclWCfkDLXhhY+AD99YhQm1m5csif4FgOiTLv1u+6Es+1Y15zDhMCTi7LBhA
m01JMme7ZIxl3dugcEIgiu6pjSXLRaabYpieqTlCLWSdG8bDkfPQZFpnTUBPiIS0
SbR7kDqkDp32Se/LegssyYf3LN1oHgUolvvBui58647GA4zydbHzKzKtBv69h5Ee
cnqt7e9rQp2zVOhKd1hbiS0tjFZwePdVcmF8nlMr2f7yKKY3lJU09OW44AbRW49h
diSmyxl2weDTDlM7az/fjrx2A7K3Vy2Gg7tGmKq7uvVV7b8KwbtroGDZiO+M1rWx
d7ozKucLDyybPliXnkJbPerAWGEug+SJyh89wlliA4gYGI5GrG727TT3uevaRP7V
tqvX4axArg+5GpTYRSSyAg7TWBOHslwxae4Zj474VnRfP1lvITPXWfjP4iXxMoVa
9NaKIi9dF3QUKjk6nMQTQJVuO09peRkT7G2O06dFjJLqcuS8viANdr8yEGs1xf37
p1KmpjWM0XTVQA/+Iju4vISgXKHxffRpeL+6om7WWuFV1VhMRCm9pG7xj9d7I1K/
eM77l1iR4thmBFYFxzLj+KBlpPAWCozVcjdABrVUoYPACUIYHrSv6wPBjB1ouLF2
kKBFUcti2CO/6cS8ri21DXPY3ShRKpi3DGBgorVrTWjXBgvsPtAWwn7wGelQ4m5h
GdQWmtcAeadVi018K24ndC9kfAxtB+RqkO9cKQulUCA35+GDWdTscsEuJNWVLx5n
VL7amQY9anqYz1MfLmEHQTXBu6QaTOGT1rWl1rsUwsb2RzzrWpLxmPdK/zrA7qTF
n/2vz562yamtiX3GPNdPuLCt55yPQX34qN9Wy8KCQpWvZoJ6trd8m1jV4U/6iHqZ
CVfEu2LUYRlsi7iqtHeDyPv1ZFrUEoJ6TS8h2mlTZ65S2/nF5scNhDS/UPv6teuO
cMWELoQYHm1eP24TKKAj9azXwittvj9M7R5idISR75u64QkKmGv3hCQGKT2uDPSR
A/9L7zAkGCcvhMXmUmJqIB+AudvFIFx9Jp2w5J+sAyeu4m967maWqfCYrC9e0c+X
5zd7gZV7Z+L7Izb6s4k8jLU3ldHmIscEQoUJxurQx3yOlPOY3riU7bbJ7EpfhGYV
OeCC5jGMT0xi+krUUgpqcFhV8X676Hx4m2KuvfqUJOE6sKrwJ5dALq5o1eKUhisi
PJANMIhd/btCWMUcdHPoi+E3110UWPnjf4qUOp1hNFg0IVBczS9NJShyhRJeb3+I
G6y7mQ0dbjW0AfZEhKGQ4+5j++0wde1bfaNnBwRExv6Cq895NTHYH+7x8q6O0T8+
oOB/q6c+qk0wbnzleyouta6LWSq0oLk0bEcQHIzSlraUGEsm76ofxToRp2Q8FW7f
xmEGE12x8SvRZ1WT53OH8ggoRJE9jH6vcdqFP1tgqriErzXFshijcUqLv1vNxV35
Ny8LhbMUMArHQVbJrBoBhCqX0loQF61RYAFYzCBW9gZAOw2LIYc69dRPtM2hUqW3
BIDlLBRMXqGHhH/q0edC7stpfx9GlfmVtqN0UHhcBrOGnAIuqrv2fZPEtWCnKn4o
1dMfYHzFCMb4uVHuNGa+ZCuvt9xtek5z2zo6kkg4chBABJKGd8Fc4hh1qmfJLk7z
`protect end_protected