`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1952 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
kGRKN8lkTEn3oWsX7TUV1XpmSjS/9k/OMYX/10kxWTn4A5C8eMqmwbvBBA8CQA0s
rv7ivDjMLpi9iNK0nIxgjoKB3Z6DALW/nP07yplASk6y8veTuG9o06paE9NDyXES
MOiz+naINvIQbTvQOjT8nyWRFanDpWQnqOkIX3ikIV6ABXp/E8vtPmFVe2s4Cno2
ifZL1cwIWhBdd4F3fsOsAMjztfpoKBYPJGx+fzUSUQS6LwFJpsVbuiBWH/11kuUk
eVJjAUap9SJwiC3EEvgAwH4oRtyxeW9mMEIeGSCrMDbV0IgS/APa+7Tp0ZikotUy
MP/us+oduyysam9TR44pWQnn5ur7vmslDDM70Fv6E1jQSET+Amy33Iek2rj9Q/el
ttta/o4HmBfSjcDmrGvyPhYROXzQVeRM8nh1Cu+r6kT2+C3FC9Cdsb4r2gbmKMWQ
b7fscMTHRzB7XJ2xJpOpVDfZJobjXysl4H7bMsdoGBXwLJh/CNiHHvsCel6UrQsx
8ezpXtjHIVbJrO0U5boLcr8TyMyfUNJPzBeUyG/J0ljVm/rmutCvlCGpf7pBxhMe
AUpyWAiUvYTGRGuqywJSvUbHELYfvMRIMqfC4oEIwxVQfCir3mge9jpVHGgDKgKk
+Oj0dVB1hWdhNfUxhVLQC8P6K9ZOf+UiEcvaqkJrod9WOsxfNufMH9xNhC77UbpI
ojmUhB2seppPwpIp7rLFTxwUhCa2JgzWCpzrS+g2+x1j/0KzzM2/vcnithoM8zw5
Q5NHR42e3W9321Y8+q07AHj5kygIe6dYe5z/vE3HzLTeG2otjqY6xvWmSNCgJEYA
jKlFVUredIkm4ZSDnhaJo5dBlfKMKI4ZSnwrv6wBohbrYSSknriSH7A4WdOAh+RJ
V7s/aCKNLipWd94NwIuZ4D8r/sQTHw3rFS8z8qqkEME8Le6RQsUKOtIZIgIAVowr
lFwuLJUc9LXW8EWVP8O9ts5sMiGRBDfVciKlP9r/M4sU+14UUmumAT7keJQLrEHe
XGRZK3RxIM0fRuLWjYx1btl171XZk6u+PyJgZm9zU5i1WXHBjRfaRBFyAHJE+Mx5
csX9Wq+eySOdrIO/JZITOTQRs7An4Wk4uD638Uq6QFTm0QjfB5K6G7rvq6Hr51oS
MouOTRe7LWX8f7KnFND642LBICDczfW3LKoaBXtjJF3DXogsGYI+ITt5kTPDPXbN
qAm2HW22/Nu4jYY63Z1/14m9NICmRDl11DQcYKVJiCuO+JQtoT5bHmPzPJBJIwfE
8ztXYqb0bJdU9QFbc55lFUERV1hz+j7c4jcU/czukE60qcuI0kOg7AUh+LcnYPoS
gIsyjSzBOGPE8fVE+T3DaJQ4whVSXsbcq7Qcb5JH0raxE1YYWZsCWUrLrRn77LyP
oyupwdRjB6u39PD6DB/VftefEHQILutny3b54VXISO04SZBIM4B0jSpYEevnUVBK
01TifZ6d5y7vN+bCBd0IvDPS9KR0F/LhRNQSBOZ4OZE9t6UaFeyT4GltW4rOIkFd
nuLti74SZO2J9xyCMXNfqaFEACpEhNqtbmjDpUV/bI2xSserdaJBsuwHb9tXYzXl
gjZUR89IbTHSPXiigBlDJq6Bge4LVXXOqlXrqTlIU1/WcMLaZN26rzuGbmpThowd
xInKQmOuVLHUTSK3pVTh1By1gkALuanSWomnCrg/x9X5rfjswCS6FaKylitfTtbh
kZeK22Fh89TPzpkPysfLWy81TKozUQkdpV+QGkWNzdIQ+jzzubgAPcx12Ow+wh7e
ATnuwsWBgst6WNhiusF938huIqvVq1YsaGxXTrmqMXeNijsyd5cPWViY3WkPzZ4v
4D9Y/5z+c1R5iKLVApiwYLPbt+IwgEjjR+huWJSNfo4UNhfjF9Sh6wvNCnXxHWsf
vp/ZpvE+XChvywAVYBGzUUseo/eJt28pZ9pdu9WXL+ZO/9Y1BEzHGw6hFYWaw2is
JpJdu7eeeSwZ7ETKz32sTdsdsg0CFOHL4q7+0zaf72IMoHGzjMQbSfWLL/yWnQ3g
uRVbU51m9w4jLs7ED7Vpgsj0iWU6Wm35ARqOFyu64eb3hcUH7sQyrAc6CZMW9Kd7
CI+Td1u2jguybs7VWal9KNVmenXFpLg9xZdOmofgxmCFzvRmnI2AkqaD97i3Zmhu
KHi6W48lFxsCmPauZQWGtlNqO/EIj9eZqE63dqRud8HZ0056r66KgvyyACYMB2TS
sjDpeHaEPitetVWkMA1tytH0Nt0sBj2F4NclLRISOs2vOK7pzil5Pl74WqqvCEsb
VJ3wVw0BUeK5D9r86GBQk9tNPX5/oRXgG4jYK1GEW59/grPyjZPG0UwZuWtbiaCd
o7MJoQQIMU4uTxgR/77nZSB2+i6A3GYmO9qFOmEIkBqz9V7cKkKy2dW0YqLOvHOy
ca7NW8H4uxcW/UTjAqFNKeQ8s/q/kwFVEMilOmUZqwQ=
`protect end_protected