`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
hVdJHWSfELCmA4ds+csnOQAALbB3ps7EiTSHEDd//nts1r+JQrRE4d3bDPRJpiX2
Sl8d+xAK9BIi4i+3ruAzYvB6kuD7r+gs02Jsvd/1kn7JYK4xBxCjtdDFjVHOTEl1
sSh1oNiYUwLuwR1yKfP+xBhqxD2Dv6pCKhH1NdGilpJQ6cvivGkSunAu0tzP76T0
4x1pB179E7uIeRplfHWX03KzEBF+eVtfgXVp2W1BGjfAe43y1pCvNYZOh1+TY62g
EgAFgbo7pAujZxZy/YSiZjUr2mGp7o83qMXyusx8+rQ41D3X6rxfuP0RiId2pOpC
6oq5Dfkx04a1dk4s8w8cVg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="Sm9DkM+kBxuxXCFA+l3fFkxuSWV4xqRc4Nn7Ji3ukao="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
m2emGBqRy4AuduN4dffN8194qYvc9UXRqiQc56IrQYMiIVQPyh59I8SYabcDdspI
7AFHnvKD5YaF6tQfxWm+mlcmMEk2Y//aUjxeiGGs+RkKgbHitJF/K7nqg1dmKvDg
a/GaBCq4Bqh0EehlN4ntP5HxM4qcvSfh5m/Coe3drc4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uG91daMWA1mGkhgP3oZKMYye3UAomMWgG80HuuXg2E0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 35344 )
`protect data_block
c9NqBF2D1wSep1rW7utzHsk2j40aow1MnrccxUTvKej2Q1cyeDDbgAml4eTSXI8z
QYgCADtWi7S8BeChdv4B2VxKcS7CMq/DaQrOy1MKTfQzfAlK0iubmlTkljLy0Rwd
Xim13c6uwpYSg2ONMAUgYX4pBA41tSrlInTA32zpf+gCLG1G4KSCZtXsIPawHjjP
/EVoOAhUXfFH1cuSULdMwLX/IGyFnMi3XTH3uOYKIoCkUe3/1FGpw+Wk9sUNv6LD
lEL5I5INbsPAjPeyAMORX6YmjA4lk5EDcKkTh8aFSETxnOkAQ0FvGcatbhck/F2b
DjqmtXZs0oPnqNK7BwVju78TxaJ0i5ZVs6Qc814fgAKoAAyS4yUONMXZqwWr1xHI
lBynSOFuylqLD4bTTlpRf+LDAJDCDWlXU44KAUS4TFZa4lYUGoZllrA4s1ulcdjR
mKjTqJrz8TZ36MKFuf3k4+GtanF5Y0kJCwlLq+8SUy3eyr5wgWdnJzfWhucPM4XI
HHZB7K6KjIu/kVvFC/33k4BHbxPeALEmAQNVYGLvooNr8q7ivmkrfRxNUAyxGaMx
k1MtkAc8VIVOIt1T6S4/jLINMLPQjCn8PSm6lie1G67WWAYMZbEbtB8WF1GBZ5AJ
0564zkmTucSEmlnzw+ThcIWQDi95aO6HxZ5/aJwaDd4IJXFMLml7Oaukyr7395/y
L/K/VOMezT6A4AQT7CjB3M48stek2i11yOzeEOsMPapAHzln6rrDMM17lk6Jdnwa
rrbJ1+9POIBKLJGHvPYajqNDG1b25zDOzovjE+EXDUNzfgAS0dTu/tLqL/qIWXkG
Dkf44h1wJ3Xwiyufh5F+u9l8cwnl9imHpxt+ymxZVPtYvFlczFgGS/7vJQMwTkOZ
WeFhi3qUGKhXXIS8TH+POSdUbCKzYJhNfGchImWPDWpPqr4guNQhDIb9DjJNsFnK
B9nsInjoxVUHfMAD6HZsEfpSqATUefBLyotJ8/nWyOY68MzTLWZExBYk9MRmNZ7i
sE2icPkll6lO09zMpkdUqIAmXt0+NbXw3uFXuU7/SOO4YkwfREn8Y1Tgg1qoQvyS
NDBdlGzKWWciXOdvF9XyC4XKbzwrWoJQXqeM1mrcxTra6ieAUy8QoezZx/gdZD2t
n0Arw0JX2kzuwG4N7NHno7lPojP+FtZG1T0HI1BuchBBKKzbHojX500qpuvZ+0zT
pEoHE6ZHAI4atX+Ec8AhSNp5QzX+V0wzoHvr4d+NXzsv9FFJH7J8sT6lOcmXpX4t
Y64IPR5NFDpowWvy7D+6ZAMwtiTBc+lZJiAlMwifB13pkrrR42QofwxgE0oKoVNs
3vbgLSCASkQYoi7oQO+u72W47YYECgmuJc7pCOM5theTtfSeAiBcHbPdz9tLpL/5
WvamGhgnFsQhquOapNInzIQekB49MjK58cs06UVL4DME/w6GWAQgPR38Lv1BxDqd
M77rabCrYWE14ujblMioAXs8GY1vGklnF7W9vOQHPfmU7LlpueXLUFpjttZheeK2
w9corGpFmtEOLOF+a3RvIFCwxxiAkmXjWXY976fHI3s84H0fyENua385jQgAlzEr
0Nqc3kgBOgXxtOzMw5K0F48XKXvPM25fPFHOBVvDjyGdfIhbNmdo3ilRoV4AXkLF
7MzJZUlJlYDNgqoCE+S4KSj7QmHwxb2k/vOmSSmJw7byhZem/Nq9kLbqFadkREi+
5YsKq1rs4nuhQ3xH6rnnttux+oRErF2tK6MW/TUj8qqS/7e/S5iXNYMh4KI5f994
BJ4VGQ+r3TOOpA78T3ITgEFdrt+/HCIeeDEz8jjD1A37bRfQmZ1CqNAHKUSdkA73
j7G3Psuq6/FrWxtjCcpiTR3tuG8kdoFN1nq8Hqf34CYqDfxQ6d4XghR6tsmNL+Km
nP+srmD3oRF2q20pOtqg3zagN/2CeGePjVeVaqZxr76QEgW5rgpzEKegMmPKi91S
lrmXHe5Vfp9xID2cI0yoFYiUX0OV7+9xlBw9wmI9yDGON2EIIzShk9cLbi7PcPk+
+oJ/8ZhGrviLxl1IGTEuUkapvoXAupvEHbJrJZ3/4XG/akIKos9mUkNCGN49/8LK
gp+AOYz+izjiQ0EqgmpMzU9ay3zuZCPkTPzWP0WKw5pT6qRE1lK2upvCbI1M7zeT
GwUGjcjqymVOSBl+VIWSM09oe91xbVWsNZI3onI5d8ob44caxzbCrOiJWw99A3ty
1s3DOIo79mGQlUNMuz79dJAOhbHFp2WmOiwsPGavsuk5MwU2AqCZlNO85Asxk8Uw
t6juisOMRdFOqz1i8Lg7yUSBv6UTeqyreXPN0t6p+m+nayrzBk1XyHccrD2vdXCC
fGM9Ts197uEZ9KiOavnjZsf7A0fWths3cb/O6D31zQg71hCziMkf3z1euCxAyO9i
UKV044MVpw0KfA+gz5YVQQznLM1Oi/Y80Vg0iY2vdK7lDsOZNJPnWDxvi5UGBBoY
PNNh119lcd9V4cWS102AghWGrLLcEVQdFqOhiizvrQPX4yH/x4zc0uZFiu6Y3509
+8TOlo2vXLVHuDj7lk23U/LpqIrxIDF8Aaun7yNaDrQXUyto/22xChvaxYj8IfAZ
CejsDKbXY65bi3dVrhL7bOya6MVN4MfQlKuVxDEyC1zQY2czUKE4+fPliLfaVDmd
bgngfwvMtWsWnzwKG/lCwSgeO6oylhvnW8sjt5T0NBAWypBSmoYhaoBQgJxr76kx
xIB0e3blUsaTCwAz/S7U7cys4oliRI+GghkG1MxFgJIUSMJWBxMnHWTflkfKrVsi
IusSAlVs6vsaf+4BbfQ99/RLmaRhF/aF6VoRXVWaPMKem266nHzZyr91eIdByzSe
YKGinXR0F30oFIkEFjQS/aCl6rUTm1R3EKZoyzpBrtN3VD3Ogoh0OEdqJuu7jIMF
DnWV4gXQimoR60v8OJnxANnTC7osO5QGkJRju7D5hYJUxU2+cuKxdkZz0i4b1ejH
h/QLAwyGFnO5zwutD4fYKbXoGzzJWtC6ZIjHP7xGX7HcZ6o+QyMNuDYVAT+qNQCF
+UHyeVwb3cG22fCkIQ9fA6JRoyGW3F98Bqvrofr6G35rZ3phAsCnJfzg8yUWz4lV
6dTbsTwHa5uf+Te2dSqZyAoYx7dgSYAcr0anPfF0/Ru02JYXrCsIvduJq/cXl8mQ
5RQufsVATV3G7p3Yw/KAzEDT24pwsBW3cwyAMFhS4Ih/cnNj+Hh38tIQnJMSdSdf
BUqhHc09wmIMnNprS1z9qwZ760sqJnYU35sbxm7d5Md9nH4cTWOZyvkd1qFlqn0V
tIcpAs1sirWygrkcos8+MB4cj/zJcX7ALXDvgFKXaH6fIWPlRhFANovbziTl62Tb
WeczEJcNJdaoy6F7y+JB6OvZ6C6QY2cUgKG6KXiR6SSoK+776skJOlwxcXHbqOEe
yTVwb96TWBzEx2TP2aaHrIlPNfGibsoyetb1cL/M9kwOXbRkN2ggqDGtQmZY0SHG
L0pZKb4o/HYWmoiI8AKbXYsg0s3hfEGaM/t7ho1HmNQ//JcFLJ76XNqoXczf/zd3
5nZmRHmw8SpjmDl6lPIm3B7YNToff7TpR96/0mFHnDqOWhasQZ/4yqesmIoLOixF
XmclQLJKHaW72Tc+JXs68nnXh8YukwEGVOWHrUuWgHwqR2GvOqTpOyd5MVMGUQy9
HyhfRtbUerxnRgW55eQwlhztVUsUnU5OYb/Y+tyc39eeAY2CP1qa1vhy1Bf94Ay6
VhvXFTwWCx2ec0Wlf86Zw8CHOw92PBhno7T816nKP0qbJolXsBRpYG5J3Q4zSJQY
dgHGGhl5CVXZWIqSYArlF9Mk3m6wBIQ2de/kMzPWJxv9pVwPQ7MflMkU3IVj5UA8
UnG1IFpZLVZvj9vD9MT/gSAhjjG+hQsmkShbasLWWuIJfpbfd0wIG+Dlm9Py8+Vi
4y+aH7lwmRTf5v80FRso0abpYT1w3mWtOSdp4/tGUA3mAP8imvTBc2qYftqquVdO
516h7pmVv0McSvFjnb8EDhQK1npwa+ZVzbTjF78MQ4GTkbIDlVAHvna12I0nTChP
VfeUSuZhjRHkJsgyyzsNO6lVT+yivxFL7N6uYJq070jVZlWlApcIrP+E1TbfQg2T
xCQDZybHKRKOgvOLmFU3FHaPWle0BaCpgny2R9U9OX3zlaxpRZjLpMPHysHAA9wx
l+uzq6DckTebT1oEoMJRGFMfIPit9+Ru3VFIbQJvKM7D/fcWrohlMXoDiUNAtM6e
yZ/kMNPh401u4a0s/GHcpixQyCYqgpETZv03qjhf0RwsXbwbJK5yvM3tfLOcRriy
G6+wBeasphjAWqK3ykJFii93Spqf5GqRMJ4UAhYEuDXNTqci2FQAQF4UfcgsqZyQ
a1luUtsw2/wf1SzBN/vTQn4wRPmtYx2Re5T3xp3+FG973s5p8+ldvr3pn2RsaliK
giTNTtqWqev3l10ukpPquyyYxF6rr7mxqESo+E+KlSSRAdj9xpqv1N4LFfHQaUE+
D0gWNyF2gCM4pfkvNW5hqmy33kiBUz13l8EbFdNWxQ2zlDXtfwl7JXJaS9uSvP5l
gcKbfNOhyiwUzfiHwARVAOdv3d3x1YQWJVWDh96XLMkh4g71K7m3iudVE4qIWlq8
Qv+YL0NXnLZjKOh5odZIkkKiEHsf1ixWJqs3mL38Jgw4OzhYhiEVRhw7VUSPMSAN
G5M0g45gxueRQJfoSTssQyMlI4DztCRhE6uVoSrySKSFU9YA3mW7C7KzvSn4ciju
HCiLqYFS65rQygP2g/hnFk7ZZrNLsBYn/W1JzES9LFDukPnn/mOtOA4jpa+i98In
9uann2RcaVz/c221eAWndRc25LBvZ5gEMgsm3nneaNEXemtlQ8eJvRwchE3pC+2n
yxXmy7xQ/HwUxWV0nV077axaT/NEeIsjAQCmKk6PI7tRP6B1LSx2SMaaHqH8SUpi
L5Gp6ygkizgDRz3HEQRXv67Htak1DseMja3D67dGw6M1HYExydbbqjWhndz9sgZ/
aMvpgxtGY7c9X1zc39ThxjpumkZzd+9Kxw+dpK1nNb95G748A0fOD7WcR55W6Z6I
mpwqb07nnVyknJTPJM4kBtKkOjbpWnW981fjzRTaPa19EeVuc6yU0XG3QXxeMOxa
LkCVtg+7PEOUEHfOQaUSpCIwbWguWP0dKG6bqhdrBKCTb3ZDfIpkmpiqyNpuD1YM
OvaRHvEIjVxAYOd8aGVGgSd0FcHp5sZ205hyrHw1KX/57T7vF0JbuGwOx80tjlqp
V2r4BoOeXPU4M8o9qjgypDwYBAYsJrb8QQKEIcMZ+fIsKJfd/m97Jf9yPUpTh9XU
ekvK4pJfrqPjTIlkX7ju+H9yQLa00AzkqfrxIjE/Zj4UcKPbXgBaep+Xip+QAiZu
w3UgPCh69dwaI0G36675YcwscqMdTW3drIH0C7c2T/m7UNmXT0pDqaTX4WButUb0
FjNJI8G0eDvW/hak9fOVTah/l3W8PV0T6Rm6zJ7Sn1LDsBL/CVoCCxPNYaaoOOMt
DEpG/traEX61xitw828yn/rED4+Phf328jzQBDC9PqbQv5Uy9NNEpEMg3FK7Vxa1
9ZbJSgHJeuK45Ve5qQrqHAr3vBN3fLiU5sm519BommvcVZqLdNVtsGisI0AlU3Qi
YXMaCfTPorHrN23jz81Z5qnWAvKsoecn/D3bnPjQj3Ip4z1ehOSI+JdsZDsrdQam
+dkA6zpBLYpWRop5ahQOWrRsuL6swkUluNb+9N6BydnId7I7o4piXRsUX2mNoI77
B2TBakdlpcF6KJ4pIjm0+RqKM5efn6Zbu+96/30WWnH1nmoruvUxnhhCCAjTQkSZ
gOio74POLiKfpFgpOsAMXuCFLp8rBm0W6oiF9Ph2zGuqCwISQAEDjgJneq58CrXT
O4sZlU0W2tLZLBM9PjlgB804QGdqoJH5snAOBcgRDUX8BGHCGRxJbBQGPwaDGzGh
uCOIszLjmtV4eA1m3JhPr4F36wFNLjEYOjt2JCQSz+zVCVlmZZBaVSJIjNDiO/Lp
nkXM23KrAEB8uXlMPXXYMbm4FjZdxREGZ2MWbOjl4lNXqzdxIy+YWZUP/RGPu3fx
kbdFhTgCK2R8G5yY390BG9itwQEjEVMGaskhPGGilr+jxw4ZFpCkcEtoQcq+BBJz
vL7wyUGI/ZIL4wx2yLOIOqpbFG/fy2EWiBpaYd5N71k/KcE/8c1WEiEGiscIzFTQ
GhWgm/2bJvhaLKjZffK4gvKafRUg4Tka0Uzv0H2+APUan9+ywp8stFFUao2PCYiM
QPi6ZqLt2QFTIwS3ZpcSLHAWu7fnqIa2Yvwpdkc2q8MRjOFjuIvhkQ1DcG1JR4p6
YdcAsuzeW3wCZ/rKDfmEAMvbs2XUHrrq/Zd6Pd/7ycxzrLV1kAm0IyGsP9/d0KD/
crtJKG1Awqj97yerHIcUpbOg1rU/Fy7W/zUSq2QPvIk8Q4VSh0SjzV0Wk6cdjIzH
yTdsDodRj7YAStJSO99nPeD7z8simy6gSExel6TMQwb0R/DktIHTzfkmpKWbeZDo
DBxEz/6PYreY0lrhfr/cptcJtOCoy4KdnWzyGasdPZZth14cTvDYkDLmhGWYFKjv
ADIOtLmczh7DizzEK0gOuAAWyxI2aebNVwDaKGwZhqrroRWuDUgV4j+zY+K6QsTY
DiwhYQr0oskLH17llW/o+LqncnnVysfOB1h1pqwwMoQ0Rp7AUTR/VqYyFz6hcsGJ
cnZEaAuWsqD2JOu6vylEpr0IOI6hu86ZwDYkv0XzrYRlEjKwkWcaMz+jrl6/GXZ1
DvgrjAS9ho2vMBtV7tz79d3T+Crbf9vQHAk5a8AwSlVtV/E/8X0Du7Gw2/cEeNz2
dNlZlBEY9W1d3alJ7Pbby3kZgNFMWPvlFDD+MqXQrHU1Fsvd5pEQSE3SS8AmovCv
mZenxYgXJ04T/cOLYe0NHUgNw2iocjsR3GMwIsAQnDJT+Fkvj56JK5V7UHrQnih7
QbxRTua7ILxtF0UwBzD8q6umMm/SlH+c1Sf52pjv5+EyfhXPE79zEYL5I063A5Lj
7djaNiJoh+/X7OogRg39LVBAEJ+3E2P7cCn+5kMwCyOaSQ+BgQwGFNJS3axSZofm
h4sypG3e05zBG/YjvKHmI5ShxlOJoK/T/fgVYty3QwjZKDFqm4BULgxl5Z0qX67j
eEq0qnViRe/D+1b8bNb8no8a6xgdQbanOCwM1ukXA0ZtQqKn+mvxjZTz24sGHu66
IVO5GiLiMnoYuZphkkQXu7xMETLTMO8pxYj5ZCRjuqMfmT1kzgdQJXTxvfVPoeXI
eQZ4I2AfXyYQyu731e6SNBLxcRZ8VsUd486/taQlSZXwzK5sf0QUuZSyHksZt+jh
mEZOeCSV9NrY05C216ncnMUkw5lCXWwKtQj3iEuFF3HRrk3meu3zOTpsw1iRb1/4
leXRhu+UBhFL0DI6Ga+DNBBNYmZ68pC/5t5t00cjaKCwaHI6/TLE1alqxVgQlFjK
RrvsCcRgsSbkyDptN4aEWFZCajtsAvyoSeqi/IW0XHywcJz0XL6x12oDLS+DZWFE
qpRGHy3UDMDncFUA+PX4dhl1ZaEt7HYrTNmKXXdFa/q8p6z6/wej6d8NEWib0vB+
+NIp+8WQwujxgGGk2v3HNzaDMbygWpjHwhCCvHnHMydqz47+Dt4TnlDeuBy1pCzW
8vitqck5HogfPFKNwn7EJlQ0Jt0KjfAX6SXCuysBtSsbJxKA/5PyVGsICcrYkxkM
4F5B3IYBCUpWRvVFjhJHhJeQXG6FpKwsj5G8TwrfGx0Xoz7knSHqOYRMxG3Po+Eh
I5N1SHEkVlfwVIuxQaVHbyWmj/FIJTv1AL2bl/MmQJyiEYEC3Q/lr5S2e1IkDd6e
+CZYaDzV34DJITW5qIdpVmclFjbl3tKOSyz5rQ5G0RnwloFFbw/4LmqiUKFphITH
wpHM8PeRqlxt6xigch6zXs5W7AndA58NMrLWCAYVj/NDV3NdAu6D59CGXMMfwa4X
Fnr/RjK45j52vTEWH+VYrAfm2UfVBgzB91boLw01t0I7JgcOstQCutNthAwh6PNA
ePtwFUiYcBgvYXw+xO9wWnvx2hD3VcqKUAYxft5dbyTl78pyGuVJWStU0KX9TzYL
9FNu/NGFfJmUVoaYjw/G96eV4hnD2gsgRGA+M17ZaKgHWNwtNh6JbsQBbsSSejJU
9o1R9JaQrxATeSQ2DFEMTMVX/3TiXHJ7MBI45wgeu4fWznGI+Ut+DJYGBgMXA7bB
AxhTh6dlmStxH8QGUzFlJJFHQlRZorrMGKbAOXaWAgQlDWNCdX+7qt4YWUDOrNSw
HBtJoXLYUZFEWBy7YdwI0pLk56idq/3MauvEDGyuup9hqPLyruslb+w9pPvdxr+Z
rFUumQQXUgJCDf8o6WoXG2a6ZZLj65uTcJLp/rpwJeuAKqKq7flOziBpwYX/tuD8
SDJTI5I7+FCBTadDmwzS2aeN+cGqWL9v+Ul6yoMqavaNl1zRzjyorgONISvp3S+l
Yya32bgSLc12Ehs34mrFyFdFxeBWjKY8TLp3gHeP9e4akzsepZVpBPhk3OE2PAPC
iJIA2sfua0N0D0P7vM/nGZQmH+VK4lLTB+b4PqfbY+7dDiBAgI98v1IFRz6/NacM
RJz83GFnLRAhKiDqHeHtCDGDQucYshP+zyD/e6wwlt06KMrFw6qhMDXaGEBI/jZ2
7y+01WLeCDvetJChtGCvVpDnwW+aUYSbkT4M9hICjB0ggKqrtLweEx0l7qhyNZ3k
hgQ3s+z/BBUqvI80HGipfyVWbhRIZvsKPH4n3vfIa32KvYJfnrSxS65Bn09HH9p4
UIGCAAEhZvy9TVVJXXoDY8bsQxh8QFOVW2eMtAPzz/h6pCbkvxNRUjzYLihxxX8d
43KOd0qlJrrL1gv6lNacc8eirskl09h2W6XOWJ3hb1F+IoQhVmCxnjic4vXw4FeN
ItF1JCGmBQKTG4kdC2Kfh7HGI/2Q38obEam0jumSrE0h28rh8zsn1CTfLK7WfHD8
yNWKyCB/3WIqk2UgclO8gUNsbYpniaK3zcJTBA74mIUTnX9M99UYhYdqVb+V7U7g
Pw3lMrzjv/e1EPLdYtFyfkb+9qFH0GoOerrh/dNuMJv2XKkdLiLnkYqxj8vy0QFE
JMUVLXnm9COwCHnRGOorOJ4UUIJk/xnaSp3CJAEFkeyiARJ1eIAqYrKa8du3nG2p
vsXuK19rGcK6zMbvfuOcKKoBT1/JlX0Mtaf6HMllYvDjcroc8yiEYNwnWQdJG/CI
gCFJtytkTyZcDCDPyzkJBkSu04TAbGehlHJsuCo10FdMiivuYfgJuSfOD7jL37bu
quduURpx++I8ozWjjRsjfPdWuEsK9yw0yg3jbmuzGo8uKZBV/9Kmu3Rq1tXKOpLA
nQKjDd/Qf8CE8qf0q2EJl6hGCAEcZ6IM8B+T8p9o0y1mwOcYA2SDhyXJuiSzeW23
riZhD1alsGWsT7n2yzuzoGjUjtZ4pQ0vpSWbIxnUs8NtyJ65E6soGc41tDtDsbRb
2yNiATDnCWMsL/8PErF3MO/7231fdJ+3v7b+MhNQ2lLEhRc3vMi0bftr13U6S3nJ
1CIKvIB6Dx14LaESy2W+M9NiAknj+SljfCc8yN4URHbZ6kkbJfvOD/MM8CSH3UD+
/rfcbriEni0WC3Ruk0nVDkFDlD8EaJ0yXPhL/TU3K54b3vY9MR7zqWvpOLwUDSKL
Z/pY2K+Q2ywrE3a/KJRXpNqr2OmTRSsCmnRxt0bNZHbAtKJfK5LNzJYTrWXAscg3
EjLmeZMPn4tQeUyAVY1pEFi3019dFh7W11ENBPKeirfftE9pt5boxDcfX6oqFRDK
bGLS+gGwnwzF7rTehfFUiHs2MFdmscNA/BkrjsAvBNS1BZR3kWv34ySZk5vuTBGA
5mcotFcjSA689DV8XQ+COQXHf3ZPa50nRA8ExGexSYiBEdS/KEzjTUGMZFejTjzy
xeMk2Dc+//mrLoJutqkttQ+Z7/VKAx5oR5mB+zBJNRi75ei/ZxPxt/iAvgWJpJ0D
MRXQmWvBEX9voI/g8W/S6G/Jy9L2c97onPmk2HjqMXQu4bWyze3kRmxR6XBBZIFZ
XCu8i8yClYtsiHj2aPodnMMRv4OpFFLhOz/ebJwt5sHRqCNMDqi9r9LE1IAMlniN
IMUEUL4YsaReVqVKAEHqjdFQF+5olDquv93Nt13deAFWIy22zlU1SMwZ933LH/CB
93Ey0wXcLKR/r6xHGKMYWFTM8UEucUYXO4QjHMPmzutZSLRAFjKSnH95Az2aR30D
9z76+ijSS1+//Y4kdMuq46oRvJM1aIWRUdR8kQMzd1RUhvtJmnweKxsUUSr65Tcv
C9EvPeYOVrv0BrKjrBhSVcfbGHX4HwSWTILTqkPaG8GLli8YIE1qTAXeXmBvmGDt
rnniUrpvNaDjC1eCAyY3qAQtqnzM+Ctc5SyEVXuDGrhTbcK7ZIEiIDLnFottCOJr
WjZBeTYEK7wMgYoYrKlfOOLPH6JcimxgvaTBHNz6sHLe2kgcepzf7lg5Gqjwt2DD
1bZCqEeiBS1bd8Tq3e2ulPrfoOWehWz5BhWdGKJVMc0hmzkmyNeHkz0PNM0QL3aO
455IUHckZSIZ9Aw1/AP/wXUbsUAExkeGGmW/dORuChf28SopWTz8Q40RytGTHR+I
P2Q2MuErfaStV0gdXO9dajPZUejzEIDNfPVzrSTIEkWkRbflT5Q4V8LBPG/gJ43Y
o3CJRZvGWMtp2Zv99UIQGk3p17PG0ddC3KBLqsZOWW76UI0iH0e1X7ujhSWeA0S/
6q2rRF3VPksT/Jci2eJUtDUEPd8OJvPKfXF/w1eSKCbEE2yKAHIiM2AmAzGw+23S
eIUgBz1H3nnMdV1LWWobOYuvHdLSHfzKWJ0R6tFG2uJ7XZXfRpextW6K+dfWinLQ
yss0tWxAlxzeGXX3mPBe/NyEZwxB2meqQK6aPQfkYSg8I/lH5JXKOozucx55Yd8B
k5RjYgxSM2YtzilOWJwCo7D29ql3HLCcGkxDOeh6gZ3A+jzmWI6FMLYj3iqMbBKf
PGgv+TpsBgY54cKLxUbxnL4EgAiqhvWK7+R+f6ASICm4//92bbGT62aRgBA6FaTs
I9i+PpY0Fq5vExA6MWUD8E30m15r8OwbJeusnbJCRoHm774uZqc/5Rwzy2aPpG10
4ZXDLau3OYk84fNuM+DR9UGoBw69Ux9orlG9unXCN+R3LCkUHrCloVfzEWMMBCoz
XL6XdvKFEkRNSx2eM745UDTY8kcVCcSMv6j/P2Db6ccPtomdooTrBQnZfIhNDeJ1
9HtAlMJP7vGk1ZBjpVUpE2k/ULsbPQF5UUHtz0gadkpys7wWa9CmAAULAIewJ9kT
sXM9vIfdCrdw5/NqU4h5nUcOKVlfW0UWpRYdpSXBxposhM2SPzpHSyciKaf3PkcS
kQq/09xGdw4ODgDPiR7qaI1cJJJ+HX0f3momFKRLCdj5fe7opoeCgOtk0olVJSso
/feeOfo+E+JK/MeAZ6UXEacSjPj4OBRC79SPzQqS1D2kCuGeMLuXJ9+nalERhoyQ
yUP/wWWNOoDW8Tj6xdK3yfIj06RaAwT4vODMTACzuTNlE0BiYafSyk2JRdoYluSM
knDPTWzFsG+m42DNGL3Flsv/TBKhc3p2zKq55TR1PNYsn300SdNrIxwavuyZsMpg
fNmM3U9P6N8JyEfFnCpmfYu+OxcwXGLs6RK6tAUNT2eZIzzvBXdmJIrtFkSEf60D
eNaZfg+HehxCW5Ya34LsASkXChPhFq5dPJOOx3jZIAW0gjT/663qPSU6llHoNBBr
v6O82MPiNcTTRTDe3roJ4CvkrYS7TSht5aOdIzq6TzlW+HDZeMexrWzAze+11KlT
Zl9Z2AHnpKP2wp61Uh+EPYKtEx1YNp31sfRlyRiat30oP4qdYtKhi9yS74oQdHUt
8zZ4W0NaN5DEnwVybkHVe0YYANqTFUKqUzs+IskwizlKTS5JEIz6R4pl1Cm5bQej
94fSsEvdJDkc+IjsNrWHN4oMXrZAhpakuu5drKLUgbZO5sVi06GKReEKB8eh9Z+0
24htAC1jlijlT7cLW+q6+JXtoRVebXMY0wdNbnYLpKtnikBKJBvFp7egTKdZmADu
BxLjCgcmKdZNYgAkagWp54bB3Y4h+j4rMr48pGJob1mtfgAXgwXDhpRGSHiEbdXM
m/bPoknOeDA7dH2JhlhwvsVwKgCp9YK3+WIjBZiX2DXEcmhAASJ6Cgbm2jSwUEW3
myqrDUBn4jRCWNtuCq6sIbqqv2igL0G7l2/TE3abUcUSJahW1Q2foZLknmuh7bAJ
qLYTmLneeYnlnXHXjLBfu0FIEEj3TUY6b/AxG6UvnrrZc4slp+KyO+Pb8wpdDkth
BsRnzyYS94WSBuNZwcZOQ7bpP/0FDWwHaNCbhKA4Wjacj0XvHH5DboYlUoWQ6gGw
tI83IF8Z2pBos+IwxUWse/WgpcVhMF/LSd+9Pw/dtWhq3CgPASjD7Hx+Xw5Pwzv+
wYD0SpQxLN/L/V26wXh4O4B7iPsAfiWgPz+Ya9x9fmHhmVXSl1tMkZ91wkJxKImB
h/vdVLw8Lr8iE5eixuxh/Byvxlblzrz7Fv6P2rGAO3ytqws7pjXA7qPGZyioZ5fp
1ZrtkLibk8XdnFZIR80H15u5M6kRdlMOfBRdRcDTfmZv4DnE4oDPcRZnCElfpS+A
UUGrCBVFKAWrBpvUAFirKpHL9OFuAXEt+M+/2L4aOujCdMaCoBcsM/6WJUHnzgmN
1F7wndkM2Co7firAPewt/Vjf1a7EVuExZcdBd+kBwgekbOZ3ym5R6oI0aTAvcmDm
DJr3DP+0Ju9gxfCmWuAejtJDfNIRUgfSiaXk+75SxgIoAgRmUse5ySCHM/N834xy
EHex7nBrHQAAREJVApyrH31rsFI498bi6LQVzGxOl9rFafM1OrrICSGi1Uxl3C1V
XBXiwRrmjxeF7TUoh0YByJxRMgYZ1T9C8weWYxIq8JQUb6PH3uMGW8No4tj4VYis
qtrf+Ub44jL4rskxupYx7k0jUErOCbTC/Id9sRf5/SDxJq/yDuAnXxQneWNgWBH8
Vxie134iQD2QUO9sp0S2tNX0fzWaIaXb/w4erCdYgvclpGkYO2a2DKQMoP2gaazX
8s6gbdV+qI7jE+vYGs5aicXtgVK7qq/gE1tZWBwaN5p47o9PpPH5Q4qsA5r+2sbk
ShooewMp3meqNGwiJYDWGOBAJQp7bLT0F5bEmoZkVdMN07bYrXxvsZY4HLKlRC5E
/sFFIxh01RrnKwOwiltPM8Zq/Bxy3iq5gmSK/HvugtwvzKKpsIgfw6Fsekna+YU3
ZYIlsWZhyWCN0WOXMezN8aRP5711mUv6N+BWPtDIAT0S0HLpW/QY3IutmqidPKqB
ikHcLe0OSqp6hSCGmCECZCLl7BVEch7KGNWkuqE4/lAWEOlIeoV8px11vrPs0d6U
aSnBxuUnaTe7RIy/yY5vjyzyNwxjC9EOcOOaKZ7JNGdSFQsElo/H14IYJ9282fhZ
gme4mHIfw4kuH2m5UrUoMeX3TBLQckMcgJrjpiCP86MuCzoaAt5wzh9nlWcqFCrR
xhg16GrqSgtrRyiTBr2bgeYSIvZDkxGGaGxBRBlzpggPWDQjpYIB1w+iV8gKFz2k
4Ob/zyFh1ApN3L2a52Z/VmC8gDnnfNlHrWP9akd/p2CKAmLHgSZiL1qCGbjRdgx5
T6LYI0zVj5EyR4O97BMCFDP+4whbMLb4I84xrijW/Pc7tNEX/iHlJOQgaqgGN7w0
6S0m4pPCq9RTePfmukks/skaGZjul5jRy4tbwGejQgtkOf9Fhsz3Ynz4CeQJxSaQ
bFgA90Tyu48fa4aG0CPvDrdrD+eVTLYXBUewqk7bb5ewuzNqreQH+GzhLI3Fc4uL
9/l4jdZZmP/bP1Ulwvw14xero/zl5Ch5pZWYjRyxbkCapMewzucDZcM0IWCiyQkQ
TWHKGXTmByUnR1ypzU7lCb8OVOpOzrsFMxBKWwCJnjesZaWPca1fUNEyLHIxvfaJ
mlanw1NimGT2J8s/PPqgpktveUmpy0e80OTEMkTugmfzh402Oh5GUppK7KfxtLjC
xnNNckYKk0e8vcYEevsJULW5AEFGMpvNBFrBZFRKD32XtfDp2xg+W3wQ/K2P/PJ7
kapXHa/4C7wpvjWwm0/EJYQGOvMHjddo20uIDNdZx01ahAWRIotEWwLVoO1IqTSG
nEJCVdVEFLgNcWJQuVFrJGzwbYVZ/mXsNzgAREsnbqCrnbZvlzlX/PFwuCih1gH0
7sv2zCp4QAaDnVMlFcbDzAjkrLcEYTm1dCEDNwHk5EUk4j4R9cGP36+vC9sJGPMS
pvR/DzMZQ16mK/6b86DaDsKfB1H49kc0f07dC7cjdY4CHFSiybCuQu30pCeE1bzq
jOWvRTH5x+jY1GUcdQGtnaG2W+7Q3+RYgfOlhYZE3M/ef33oyRN73aeqOQzta4h/
hgIM9WxgVFZbgZSEvBXN3sP9r54hfnnO/Ryp4EDJSt93Eg3o3N9e+QRwcw5OqOLA
TXXQ+C/HlowQXH7j2rCS/t9QvcKDeUJSk/jVnhw/3qMk3dWKaZML5l71iI0MCQeS
eEh0OLth3UTD/6pw43I9x2Z8+xwak7dg/jgMV6OVQJcD47hkKinhXEXk/NlKmVmV
SsDmmxRGfufPBejcL+zp3VBEmWMFeXvR1Qje8NEzkyoNLk7aJQeocQEa3eBGUppk
QyfjI2SuMU8yl76RaOY8AehP/dlzWdubqVVvKlhvYViCK0AC0fyRTy+cOwhpmkFp
T8/sTGn1zrqPXhs2eSYrSKoZTlSt4YQnTjnfqlwRnffFwSNDbxj0jEGJXX8gDMOO
NHS1+yauRmySu7icuiO/THN6EzGFO1lULLFZn3JJy+7ROu5w08GKOdjDsa/9rqOe
rfNXJ1hVFF2FPhky5CDDIOJ3LbVUVBOkPDiELNFymOoO4OochEnFXpS99Hms8MpO
q4F8zUwZYpeGdtU2TpN0SNXGU45N8JthLbydNJnrLoQPXY6sX1UeN78KscJUyO1x
oF8yLXggAEHwSCj4wopQ0/OzxXC5hL0UUYg8O9XaGlvZrxuxHCDzkQ+eT4qF2VpR
xMwWOfDih65gvbXs7WDRUGF2WvZP4BkYzJCXshbluIxq6WG+VkSkFQa1HYmRc+ji
Tzisv/+IyDe1kuZgPK9rZ7EQzzxpVgoawExU6WOqJm1lADiDtVw+otf7r6r+CBpX
NYFQhay3hQrH/CPKkUjvkkW1aNxtv5aMjYBDvXmtCcKaiJvgsYmSEFk27cZxSllT
5E6KGQPmn+KiJBAFsb+pq5ucDbA4MfLrseHeZr5+s7G9S/dxXqVVeXqlyU7ELTlR
yIVXtEx/uoJgMlrEBt5NxyRQ9PbH8+WI1c9dVEqecnNzCuIAKx14UK+raClcWrbw
awOg2aQsj1hUKrGQX7mqrFzvv5Qd+UZYv2WvHp+H8bAKpfu9WvRbkngpgwRJ2Zwb
mbXQD5xrw3FHyPfULK+VhwLQTLrXi/bbK2tCDe2vmA+FMt5AAHDZMLAlhugmq9QK
qDj2KTHq9X1GkC523OSJlPuxKRkx1fz7G6+KmGASaEPi/uZL5Oma0ryZc6bk0RvS
q3YbTH+/M3ChNB1hbKwMvV/9ttl06D9J5oL8A4GH/q+I4ZJXsb+2rww1ZlLxG0Jf
mCLXDbykozzUlSv9kyqHfWtY8gumymHENc9qhT4e5uUZg8NoB+SGQiqiu1cZhrUq
M7qichFDY1jutFIDpqKyRFvpRzXPj0qCOe4kKuGYL7PNj06g97GaIYAM7rGlbHao
0aoxHgI8exwFsJvjsLpiPwesjCA8MilGWxf+M3Rq5P3YvDFe+1h/DAyugD5AuKrM
MBbDhYWeCF+tnuczVivl0Cea0v1flVNSSg9MD+7rQeAt9K/zpWzq65ianlpuotC3
21uDzoSiRSQcu156ZzGS5K8f36yBLq1AU3Vo9AQ0E/Oskh89ew2ijSWcHD7tBhU9
9932AjHtg2J9WsVXa0qvWlDEGzBYxo8hMZCuc+KZAA9N/40mKiqa4T4N2hrPm7Aa
ia89Rsk7YduzIJZCLa9IVPDhO2dELtMTZcsJxldvqslWC40MgRpiiJ5D26ohoLTQ
Kqg+d4KvB6TuN9DDNMnCxlz+u0Tn1jTrCAsBZQfX4O1vnZlm5ecXwT3c59ERVPTg
3wDzZdraMyRdzDK7L3AkCXam6nLQbhToKhqHlbCLTbi68Uk8pBmRAPbeJ5jCoHb4
PWKKYIf6/rxFa3rSRBCCzWLSEzGLE5RkKKFzQrZtyjO/jzMLGCGfK8hIiZoLlQSt
tlA8VB+61z1LYdhGBCbMr4EC1dDbWVj3Ca9nxPKrAIX6CfoGrcgP4uEEmgzJVicn
kUoYV1WFQ1DowgQbps65sy1WYA7LKXKC6DPRgMoFZ817VNL7Oq10mnXWRodBpk6a
Cqdmk4A0vw1FarOwCBkFQEEvzvvXMRWsgMwvfEn/pLI8Uxl4BX2BnyfGyWLAxyKN
7ekv0DS6WaqzttyTCs/1LwSH3c3+5SJBANoW0uvHnAkEOAX7Aar9lReCoTZvKfx4
c3Sj7wXA1yK83/8Wd3HceObxOJ2c7GqhnF5mFxm5ZirYOm8RVAIYOCV9N8YCXiu6
t3eyCydjUmophpVKiK1I5tcHKYco+bkRHksMNWFRUWpurElI96Fdp4kgPbAbRYUn
Btanz/EvMwSc25e0nrFRSUmdMrN1dE8IHcbwqadz5M3RcuB4Yfd2KRi4fGOvsdY+
KVRN6Jllj81JRjJkAq85I70MLIK59rHvhSrcXD+rvAgjBD90IF0z60RpqbSJWhm4
dj93stJphg3rvOtJVQDz2xyZV/72omeIY00xCtmKP+DtIdTThd3M4GbpdLVVJV7D
18aznABfUkcXUs0ZKsb5VdnPHYn6ZcZlRdpOIAdQgTzEa1Zp3HrJbQQ8h5GKAU7R
MTKL5ImgiwDDG6Mxi0DjKpLv0OlMlxx7aChBrbcIr0393oRMwS9+ddbgWyD2E4m6
jFIIlbyTu5yZZHralkIB5GtjVNbVMqCfUMHGXEElQWEb+HSgYh+mpo0n1cwnJPp7
JCrbKJxTniCTNdSbRdwsrkZfsKpvMPTdsLipJeKwM6JqOXMGqLAs004Z13RJwmCV
sUfrO/QSmhf/xv/YgrfTyWEOJTfCRrvuEetPpr21a6+TMlTFdCZ8TrQHb2sSuvO9
unqAQqRYqQHtUPc1ohWg1NIPbSX8zT+li6EFEhtvMm6ed5bGw80+Q+ULGDZ90WiS
rG+h/T/zBS19M/KwdJS214BRbKXFg+8Cry+RcuyDqT0I9zqXKFxRW+7JW4rU4rEB
508bPPYPvKnMPVdgAnVqS03GabEEFZALiZKRwW9q2V6Z3/E0zFOi2oQHZG/0VvTl
MAgARABOj3r6L3O5PJGBW1/uHUQVf7zX5G+KHMdzUcmPcFBT03zxUIxpBAqZNrdt
F/Zkzh3SDkQjjqV9nw6wYQo1GGpypVoJJbWgHSNA2/sQ3kJJeoh/UljDPWBj6UHH
KGp3HfH/T7mFCiZonq4g0ds73V9Omp1hxZAATi7h7PbrYIZVcf8MhNUzmHg5c2pX
jfjsbAU/k95gFEw5l3I6xuxTuTFiUEmGC0QhRvCfybLZ2sgGMdqR13Ft3DpdZKPw
4UTVnXQ64W8pSu/XPv9SGWtd2sQOWjwPov9PaZZtDnD5l4a1b1sm0+RKwhr4oJSB
8eMow5D265mU6ciyAbR2wr0SZzmLjLRwWw2RpRSjoTRREySA+ySDbaPITpg6DWiR
MUHwEAeK8f0JND+pPmjTAzL2n702pc7PoaZciU3S53aHcMLWu/SRqvzOR7rSxGgk
+liCjFV+Un2XwbFUXL287Eq41pIpLV5E3HCAR4UIqeTDXX9GSy0wTdHypeaXtJDs
Fntuvrg2Gv+K9Fx/8TbhsR79b2eBIi7GartHAJ0ZTadlXgaDdIbQzHoj2QmbOEae
iFvqMMlgCM+oupD/OAQ7ym1oyt/hz+DLnTgGCROXWRu6XI9gC2uhMPS3CnPw8PiW
I+Kjpaepk0vYDtklqP06Ck8RfEhme+modbO+HHzaKQAtzYTM5AMY3C6Xp7picCRv
TrbjL2hnP5PzI2aqJDi3ygWZXNjTHin3wuZi8uCMhGfmTuVp9uqxcN1qWJwi0p+n
NZfkYnhp8LUHWDAJuHrAgeR+6qXj6jMYr/FlGH4g1qBZMYQ6jNMuKttf9XQfgh55
fIdFz4z9r3mUGgn3tL3axkzxQc38AZrXQq0lEAZ7jDceLITbs2OpbwET9pidKo+n
8QDqEZTUFCN7K8rjjb5mJRNbcd3ZjDGBzYzIbR5wFzt4wpzcSyF1CBfxP1tJFX05
fCRGasYzdwJPlAN3WY76gNkGbAtdT6Dmiz+ufX6waYU8uyCESzpz7VazuUO8x3Bp
S+/PXuQPqsipA6mMHW5RTASzZJQW3ghKIJ53TbeIGXJqTroNhnAXfO+O0GCPWOxU
vuziLinf4Z2U8LitxUHCl2pEw/KxBn1pjpexJb1LgIovozVHRPR+Lg+He55bpn+f
iweTb9QN+TA4RPQfDFc3ZsFPw9JjHprV/+nTgM5GYJeOIiak53uF6TeDnmIxHDcn
juz+l4NTKU3thDZM4i/v7gt/M9Vv174NEwpia/UkYCUneItq1jDE7RhI3acHolWj
quSPzCTNOfHD47oFoxz4r54/H9wnJg086HKPBMgnxXhSQt9/MecFpsYSiPSK3FcN
i149HZVi+hT/MyyLCEAokiZLRuxJptONCQ/HXTyWUi4vMG0G0F4s1/c/zexYVsZQ
K7aCkNe7KFoqdTU203drccqLJHKNcsf+5sIvgTunzU6ywM0xIe/f9IKcWPzwk+kf
G0PVJR9vWvYSmQfBMps2KClh13o2YGutHYwzRVEKqz067k3JtxPennwxWuiu+CnZ
o/BcEyqPJOnANDZXgIAkxYrGvkvSyZEi6flrKboP402snT6WUzuT6NXvgoqJoZPg
KicdRIYJOk7BU5G4lE7IGdMQsijPVoDsesRbvHBESs6svbiezu0uSO55+4GTH2Fo
16iE8umcylfE6umlEHAdIYQ59ocXiXGtYiKrs/Mr3uHqwH8t+8sP09AN+sY7Csnp
A4yxNwC46HxLREBZ3G8yLhBNmRKkvmps66Rm7ze1Wotng+WI7temGvMXcBOBX5sr
SQwTMCeHIX2U/FxDMvGSDKjp29xldZ6qbyp11l6pCKIgb6X3FRwClrwvukmq+O6E
4+WWsJ4ahcl1MhPX0r+RPFTGAdqZJ5PKAKJNoyGzyS5OOxM+bNA3WeJvgb+nnnuk
IH6qPYbr6Ka4CD2sBlmIRjW8bXO6dknjIa+E3y9YOnfxWXb35U6VIM2v+UGB+C9/
AncFDCDD6dGIJXSzbE4wA//zDhSiW17XsLjxQMZs2kgXYNHuZPneTuxOH13GjQWT
cu83tgscoqxEGsVlJpADEZ3JJqK8WzP7hIROpc8GqzdNO1wT8wTZShJ4/g0acWBi
2q1Rb9LNRrO9NVXj8lk1Zb3qCnQPGE0BpNiWdUjzl5qGpc3JaMRkcL0unpmTSSaL
Y0F9Tx2BjjkgZFGfUAL6sB0KbcVVJ21oJYfrNMYoLNdnbYuUlDpFGYPKCZeGnxis
YoLmqfaYo5R3pr2FLfag7a5U13ZhzkNviFXly7AAKLBZVIPytlxkOKOp84ir/KSb
iisP8RGQB+IcqmddfgbI+QvQyf3OVKkscJ/+FDFMFb3nYbwJ8ZfE/WCdDo5jLrOs
6SZruwt+GN3Z1DbgBdYpMKkS5iwV9FEeqw7HcPXFWa/cYbaOPU/ga1B35tg6edhg
AhLXIu4yh9TNfCXDiYla298KF+t5kIU+ZW9j0Edp+BDoPRxSTIPeWYyKywKzeOBA
ArVMKqz/2iyKvQ6DIfyP+81LCX8xA7FhGC5Wi1fbT3949lGNYXyGb9xDjtKVuvEM
MeKcVC4HqkK1hNsXHOsA8zKunT42A/vQhir3oW97iguxlphJwKuskkP7rA7XU/oy
oyDk8QUIqJ5yGx561+UJ8QZiDR/mG9J3GErOib+j9emylom9IFs6M+0fJeXCh3Px
sDgXh7cMbAxznm1pf6eoReNOxcxMU7br9EPzdZl2iFVe3eCF73r1fPFGELvqwssA
tmy821HbgA+DmgLM6x2J9QKhAmMbaOdU+LybVmUzNFeO8nhM9gUCLH+u2r1BXR4N
UoTQ+L02bUyMXImCUmJAG8wdsUJm16LRxixVNEauBXXAi+DLkSR9Df5/ph487IbW
pYrSM3rf6s6uSRu1I5d3JZMtbm4wOJee9yRe1FjY96P7vtCalfDazNsRVu+ad7FE
uCOAAmkgyULUyURXVMy6nPG4WUNNtGUWy/xSu1Ox3kSrhgr/GgzZegMVDXJPlZZa
X8csG6n/6sqlGiBLQtQgkoCTRr1nVdrTuRBLwZuKQTpi7KQmuV2X7uy54tg5qjoU
U9jEAtUaGSPVy2B9cXCzWWQeFcMGKJBnSsEB59Y21n/mmwynmVRr5NirIVlTWwiQ
XGKbLl2wZ9iz1UhJMrFwMkF3gZ94IxRspZAZ5lCHUCA+4m557AEBt5HjvLxXdhWM
6LLMusTH43xUewz2OY7Fw6DenbNRqUvEXug/0/mOs0P8hPxNdB07Y3UIt4/kpfWR
jTVcx8VDnXIbQWqqcPIaG/lW440fPbPqR3T2QsFBdr4xUbYQUkykxejhyy6J6aHH
+TtwOBaM7iorHAmO48vwYZgIdEgBejlSmFyISia0Bn86j6iS1lfgAx6PyqONiXBG
qcZEJckteMiQiPuZftygP1vcZf4bDEeu62Hz2rabi2NCMre/L+jcmCQ1zDAdcx9n
zlKyl2bXTsZ0hXL4zH72ecA1sStcDytrlVdulxMsaGimQ9iFgpH7WYBShU7e98Jd
DR1vBuH9dj/ktYfRErtiMh1h/Ca+ojitE1lhEs+tAaBOe5eVqtmDfyBe0FZdrSBf
rsPPnvGmYWUyPZIxVAlyja2TnNp+CB8RYH12LWUoR4Gd+iMvb9g75jUlLdtKYEF0
lXWidtJMvbxEKOgsuUnJSC+/k5dutKjG1mgjacXmWX9BILOcM7QsOmxgyQBtiTbu
mBM8nxdbpImPR9KUESWQLrslGj+3e065WeOG38pjOi5Kh/agZeCwMdS2X0d/Jsm1
UnZVqbq4ZKrM23PjCO0+IkrDyjKVuciwGerSUslTOxi6cgzD6pekpalG+4HMk4ex
uFezzfaxCDRhTEEIHFQCvFyMJwm8m09sIhguYhCSzIcRwWDny480eIYZsu7/EB60
KBl+ebI4I/w5frm74bVm9YEnCHiRzvaPW//WqMRHQbQ99tPzaB9CF98wt0R+WMBe
XrVDHXrSQo6b6E1MxoRG4+ffqhvhJug9Mj58ckRnFisg6SA7w0up7uopKs17vhrD
LNgxacXXyire4tUZs3F+Bv//JqTS0q7nS2OM8IBHenbFUv9EH6sPArtyV4mgX9h3
MzmR1lmkRMNJBTI0ktvAK5xMBYs4sSXp5xPeYMTCrLNXf/o1LBD2R3TZ3JvnD8//
7eM8p69hqAxDEmtLlUIUCzuxdkSjJtIXtnRyaYRUr0RbGFKdep8bSz8/w4za6EvU
Hh019DNLjYo8zQqrnd9pCrVG9yg9iyd8KVnH6tDY84SR19t+9Em4CfS/Bxqo9MBd
7/CDD680vZdkdSBYYEInEdakXJH9lap35S7FzCFMqUuKWhW/l77XQiUHpWCGSex1
BW3Hn8kAuv0294jdu8OduOJzfVkoH5Fc9xIE6nS1DnfhnoQrmZ5Rph4scItZYrWf
EOHnfWOfBvbi/aOmo4M1QSWEJBEmOtAWqSBCUE7D3BNhrVkkJmkSHYIRLq+oM7k4
jCq7lEDTN6qilhHUGxcq53QuRoSrhMiVojDWTsJodipeEdXMAzj8O0iiFvIj0DsW
e9RexqUUo4AHXVVk533SPGvqclb5hGUlxMiLaQ2AaKuUoGxksmKOqE3sKrObJwin
J/BHIhJplrNa8EZN9qEoluWko/YW7/0Uizrvnyy5mu4Hko9NCL/WJ8SFs63/xkea
xXeuOG1XZ4SXK3sPztqCq5aDJompZZADR3avaJaSHg6s7rVbto/J9JhNjzqJ7vl2
qsN3r2vRFEDfYsnCZw6OWp73djw9BUsdbqVdbZe08UwWJRAyKqsYqRaGO3wQkcsv
eHSV8hYWkbsRSc3xu8JVhXMN8bxwcil6P/y+B72WVpWs5ecMA9gYmUkNGUvfARpi
KKgLVDSA9iyOGOIQCpOIQdXDgTiBlSnfUMFTi1TOUQvveDul9XOJqvwWWe6RxfgX
lBt4HR+5IH1Hn45z8MO+Fwvln0wYGWw5jSYDfC6Xv4ZDi3JhCdpXjwh4paeDftH6
5eEz+0GPCz+BKNc79IPtBC3bmVSxLCoG4lo3KKnaDUQYIUTuwPjJn8LtG9OfAfVx
iFPjCNbtndQi6fq8JXCWOgeI5m/clVeKFMMhKZsV126OngzJXx3VIkzNN6klCvhR
xchAzL8ubUuQ3npvCZhfTEpL1bRqHtiyAPFOnIBkz5uRDtrDX3xd9zPdUIiGKy0y
BrMl1vaZSBZ+ZEXI+MlGacTodgaDjj2pOEdN4Y499dGD28lHGirDTYm42IaUsQWZ
yneI4rInX43HaDSQjgxg0OoCxVoxBLnS6YlGTyl9GEZy5gkQJ/amLSgMxn2jdmYJ
4oKRucegUWzjK6YSKKI/aVs0KZf/Yc1goa1l0p/z7r1cZqYjJPrQCkpMb30dIrTl
MmSODQRgwGpJejbtYDmUHHVPPCpX8Q/XoCCM9SDcUmMnZHfUlTWgn5Cw7TmY+jqA
ZEY7xUtZKLw38ENJOIA5EXgexa0UIAKe0/ZiG99Nnjm8Vbdtl6Jnst10T8Tg71si
iqi2EWpEAeo1UoifFgMtkOX/lhgcqYSeX0nMKYX0RzS2GFFNw04JEiEUJxqTQQmK
25bVLFsk2I63Obt58LUC/we5mdzSu6YapdGrDldloRqtuask7b537spEweKandhj
GFSeMdz9YXeh7qroXpXG3RJjmw6OILlKnWYkSf77AczMzjwH99aVUwDJ0v45WjcG
Cg1Zdn7/V9xXYQZc/DyDitIvGEfYZQGiQikQLW+6PD2jVHHDIVaagq5w3AoWYHCF
ICmoK9Rq6dxJ13uUKklh+Z9RYg2lyIPIbl1alpyIf5ztq2t0ZiyD2tIfP5bbfiKW
SGbKwAH1AEkLz5GpUmf9UTlIHMHgBJgs48P+Cdldq5XziwX+YbAAw0W08hEUQvGH
t+tJC5JPewppYJCyfbXCscXaR1uGGvA/tv6jplWoPFg+w7ThSLIlRkpKkQ8REfS0
Tz9xSVytLaVxtLgP/G2pluchJVoHFh/8MNHBskoyRxsIfme1Yb7TfrzP21Xv5+dz
pgWbAYBWGpGXiGDz4c2mToBBRXM63vkCIET5AXptynkYxNabFwIDiBOSn3egAcOw
1m90EoQYQi1+8ZGkoZL7lKtPwL9e5vsKs7QMhk386Ku+mBfGWiauggzkqeYfWHp2
IJ6lxj2m+PHW89iyWFBOFo+KJRMUzj/BbxZ4EBDivAV7KYGrRw/USQqWV3YuU2bB
0h7r1nnvfPUMhhunYm3rckHBRl16TNGZJAZhD5C1RFkW0K+yw9Q+gTo9t1WoT8ju
fXR5DMDeuJEhd4t9xdErjLYh+d78do0AsIh17uPWDdf3t6HdnbklPeetH28jNsRR
FVZavhwCKrF2Ei6waipY4++Nhakaksffyq1Evw79QxphJH+xOppDc76egZMIqNAp
68wq15gCrD5mE7Gb8zOxv4QDhwA4t2eca3zz9wMRw4V4N2Eih+ntE53VnrsZZ2jI
OWtHkcOxXv4lfrRclczqRrt10x7jXAlPDxt7APNNVjzt3T6G4b6ephwXcGgn91J3
4REGwqTQ71cmK42JCfzJDhnTh4q9WmUJ0z0O2akBlU1xFEq1PkYrsIj+3hBuCQ+7
hgwS5ZzLaVG4dp3Ybsf9m22dBDasE0O0IcC3+UxaoQDAS2LAE8eLYvZEu/jya6XK
bR03iuySiRja07YNyIU0hZX5J+Ig5soIZ6vmr13UGPQf+4ZynW6WxSYA2lv367G2
cKAJ67URbQdr+s6rYS2LiQwkeol/KajK6C7zgpz51fXmb4gExfewgaMHTGSdj6V+
4ymrYM4gtj4hKzTwsfx/Sk1zQ3To5yZ+uXfyXIMDZ/y/APuVZJVtX4lR9GSYUpan
t1HrhQDZB41qNNFUvxD57KaWW6cO5H/dDskHWfU4MexPHwZzuNc/6qCLcb2KEYTL
fI4nRr0NM5ss9R7SsDC3mtCSplBOMTUfbVzVdmUXNPVwT1ylM9KdqDHdRPntFoyO
o1Iwpd2KtmZ2qVSS14NCSpNWfEmYw/QcEl3poY7Oo32jWnkpQNUU43rC+JdQuyEc
Ot3P2SVbkbzM3x+CeazHJgQiUIa6ExjoPrNUSbsY33zJU4u3n2HZzzxKZsxOQLq9
2WOwGozx2fSjvkcDG98iWcTjevVL2ek/lZkO8KG9mXcrnvcvYGJyFpugccH4SPyE
voeqY62SHg7mUNkcUUbMVCP/KdQ7S6gUFX//n5KKGPe1eZbhY2h2PHcAoIqRF0Ox
Dmx8yYDUzP1UXdQTNtj8uM/cGYBXYXZvckaCMrsJQcreUaEEEPtFT3pgL0hWajud
tnorrgW1u++WLbsn/Cgj5MnfRDA1YT4a2bxrFpne2l2lgxA8oXLFWEuXRHhrPKvx
lZsGuKY9ZRgbRLkfSuX05vten6d9TZsc0YnTnH4sWXBEnFZTY7p6c6O9hSIHwEFG
RfIPCbyzbnmUtMLeV+GOBivN2AMhbFYKvQy7mh5pV1i2V6iJDA2rvHOTS81PNFsM
2TJeFzTw795scs/zRbGJxqTm+S3p8nmNMW36nSJR4OEEBStm/e2gJ1GeXflygRqE
c5NiSo5ire/1+oH/tvT4fw64lJFv9274bhVaXaJnZpXpKVdTtjkZu9ZnAyYBH/Rf
PHVMFYkaYqJG76eF0oxybeyfZ59TMhi3TM+JsmlTgaTmhgE34XLTo+97SAZTr+zL
fls6QzG9ANWuhnM+wJbVUhoMNi0bI2QT5OCQ3zlPa7W426VsYvnLik9l0UR3msWo
rUKXECCdr8uBTZZAcvGsGx4swIgtm3cI4EXK049j5F0w97ihdp20xa8s4ZJidybM
mALe4BQF91fHe8ys4I4zXbXFPECGmiXfup0AeDxX5NQogCb/z77rSRDnd+fdWLzH
U3dTgojvl528C+7gCrUqBeByLIzxa/sSvuv1+uvH9yvE9uoCrVDDC3FG0Abu56zZ
VvEIJVXgL7Hwr7juxBJoJvnJxO6r91mQpiktTGRiTpaK6OL3AXrLXlU1ah4IqoMu
iWPSVKHk5JtC0szwSxVeM7/o6BMqrQ+/RXBOf0kETEFOvORjaxlWQ6K+rQUjnAXr
50WXNOiUBd76wwjQOujR+K3G3Fdg8BRW1n9BNcQ4XGakfwjz3asGkqT4hxF6GMzb
IQRm6/kVF41OlqaRmtmWHgX6iSeOyDKS5rm7dEqbm0miJxhRGdM5AlwnI8Rr9RnL
lp2V6pvG6Hjpzdf8cpgrlnmFqm8aApujyvToM7oxye/XpZIJGdFaUMW1tm+XRbWw
XlKYCI60Eoz0E8tAXWtRQPNDzBEkl2iRGwzJMcspLZxpa6G/EYY/2NzED/xnlt/7
e1tLqmWjUCpeytOs5SDjzICEaZWC/oHZbmI+rxQq8j/4OQom0UpfGRnj1V1vcEz7
lYo5C1RQnG+YVo3B6yvuMuIelqT/oT0OapSvQgI36cfz8T6Q4S53w5bWMZIT26Id
7/BJ40pikNytMjCo8CdhMyEFm1FLYZRjNqfhybRyeCcRDrFAh1883d4Hg9kgWyDx
fzBnVV2isOmwdmbEKO+HkSIghFCxJjHP2zx/Sup3ezHqLMF4YpsPlSJ1rYJwAUuB
ZF1Jb+wPy/07vS7qT7OhzqQE8xcW/4mi43ZmZJAetMfllJ5EVs+Fs4OvtAS+lORg
lTSzK7l61y+rlBxtobXY/nMRbmVybCNegHqcUACEt5Kriq2eckfOccMYnqqaqrBa
R7O7h0aQAj7/OT3CLhjnBVXZSeh12gfeNi5/YmpoL69LS23bsPD5Nmf3rx+BmIuO
ZFzJJPmJw6ZU5TjH6NK3KC5G9Z9rdnfYsBJIkmIps5S0vfUMpPKwEteHXpK21yxj
Vy/VjWFGPd5VqgjiqE41edaV2GPn2XuqAl6ir7q4V504X0GWD2JJbuxm47Z+GEOE
TefGQDqTtiByB9rpeChMX/rDLln6dY8U0T4FWwmivH8Rsbv6xKGMN0Wx7l8CPyO1
BOEifZUJogkO51ke1Bgh5ZY8hKuUY+P9C70IPAn5q08S3X5VWqNTGMsEDb/3Nf6l
FiBRuwwQXw9RsRQMLUOgliSVJpnMJmwAjHHaLhScxRH3V6IuX6aunFi3/kpyXXF+
CguNAlAYUT5jVLyPY9r7pHf5sdIx882mrRCwtPg9GRPPzcr/qAlPBzHLri4VTnkz
5QSlEYgfBB1rNUzlK9I7Y1OzWY1tPzBwfAalbSCMXapg1QLnKVhWHv8/SvycgWJx
PkqimCRwbyHjRm4SMASgd5X/oCGeMrpYCO8bue1aWgJVkGu2jGUZr8JY8kZdjAvG
/U+mS4V6v1BANEAiYhm3bElKIqvg0CTFFMdzuUynV4bDFoM00Wg1XWiY67PGsTL4
tKBGI8rt7sqtC26eleMsNZF4aLVfEKpdJgUQb/CyXPWHVdp2j1dJmNWeAlMBlEdO
86dxrfUZWCImg7T06NdW6VdXqS9PHVur7t6UHX1c+ieaXA6csO2FJPfKaDLZ6FXb
OpOkJdn4Zark4f2eoWYl19TfxskQfy0dqwtnEwSK99YzTZS6aZ281qZfoQZ/xR3a
NPO15w2Q7z/HXIpv47UXjG1kt7YzD1m47isBFF1n8mxgryeiMHwVtMX2VgVAmKzt
cEQ+ZdLVhyc7w0hUF7SXfVHqR/9SxC6qiVACxN9yI1ip3yPLwvEHreEKC31t8Mqe
NDsEGwqPgGGhjzvUNt3b82X8Ue7fZMluiJC7vHHTUUJ3rihTt+t7Xy+dpd/JdzFx
HCZBDtzEoL88tLTsMpLK60wRwliXKiW4vFvZ0MTaxNYRj15DcQdDIiMq3ByG6uZQ
XpLAYxzYw1j3e8cvhAuUjxEB/0LwCVyE5Aj9LnRQlIARvYd6Ob0xTky8tvmYlALg
dHgUBpbb0J10SIcZNpvoYZwttonOb4KaArdATKLqCG7EneaQ/st/VMOd7I0t0umG
4PmGL9fSK5MJsF5gy3IKUG/nBhV9Dks5zed8eWKbyH9SzIZZlJHaqFKBqem9Cy0H
IoAIg+Xi9+VQQcy1zjBNZS1GlfEL/svFSKlUDU8sLvoBaVx71TPXuINwBVhkM52D
og0+hzeGiU8l07yoIv+ohAyRTaYD2EJT8I4yx0ofYcaOAxIzTaXAr44z0R2yM+Hf
/96NXszGpdu5r+OYVbpGBA77uDXX+DimBkm7Vb8e/BX5DgK28oek9+SzZABdH66w
iUmlEJCVVNIPBMkKJraKjFR4BcizLe0Vm+7YpylpIytuLq0hAdeALF7PiWgFqZfa
x0CmQvYgbR+aFbrZ5qaHeMrxa7I8nhux4ow0wK2h2072I+MTtsr3BocwMdoIkcZD
n7+oVF8zHm7za9BhZcgBxneYfcvz3BW+CfHeYhvBJ8CK+umdclyTUlAUiKIPratM
bGiyOfXjf+MPQaJ1gDBDnYFnrcODcgOiyFlc8WwMNOJFkluvcbG9SDRqNvCxZZx/
as+QwOTbQxx0zTc+5L4BYhhea5KsaKKXuHsRFoETmA7jSPHwulRFjyizz3It0N9x
f4wQsCGhhDEM2BFmOv5EZOyDocw0HYCasF/1mXlLWsHhaz0uDvQwX9YbTECVhhnQ
s4U6UrkPcVvx6d4Sxz5CUvTGLlg+uxbNGatokSbpQtuu7cpbUhpUaITi6VaY7an3
hzF0wvQCBEVhRZtokMqPJBylSlWa+Ljhk4jqafbJVcBsty0qsOIYa2FR2pmiliNF
NXY2MWrEXntKDmA9iUAqAy7lHS4YQl0IbIAyKSqLHEwMBpG0b6LLfVgkbhm8h1Bq
cOwLJotCaTr0Pcb9vpgeQWHZRxDJoofIOEsX9LHmrkARqTpUvjbt/zMaRc5pEMVG
JbVm/3ywGR5PY/+1iVBX6Cn+qluBM7ozqTglggUVPoSuDkbbqPiV3uQcrETzJMbh
Oog3ockwztIEl5phvSgUiHWUzVvVEyN5Ibdn68bmd4tXL34amAiZVbJHpjlDn+Ow
kj9Rzxg5I4GWomPADSpWeuE0S/dkIZlbRGCZt7TbEQFYZBaLLa5hOj6o/5ueKamN
+u2uOV8/OHLiEcjQxy1S9X95mDCiTRYOId2G3X9p/2kjJh78QzzodcBmhZuEfnst
1Ety3m3ytP188WKOLtBaorxXeT8HjDO/P7CbrimoxeET0h8DqeA7xuhfeaUpgmeS
k/bILAHUcdAtuU7tk0PQaDgCu3CLcHhHnfmnYfVKYuXBZdkukve6OjHLj2pzDOuJ
760zkZb4cZDegMuWQ/KMuJqHs5ZwTSYCEwYhX8AIPBC/OHvbcnDdPbwIH7mJzyNN
QcvToxN9Sc3XzFfaRkSEaC63RPGw0o9tVwEroLj6kpfGzYPITjT/o6pwDelnccku
nxLbSOXOfS+e7HY+d2Oqx7FUEDvyqswBGLubd3LxdC6gEaVQR4okBP6q16zO4DkN
sN3Pdx8Z4Q1di3UMcVtMuX07QOMryxpZ3+Gz4WA0m04uf3WWX/T+YUwHoTAOcghc
tu7hf7EQmyvlqFr1K6MtomMoB3GSjEm6tbv4EMLB/claxzSoOpVfz4xbFT5HK8EF
HssJVtkup73J8PkSfOoWYQmSNDGuPHOyxS/Uauu8A08DKgUgYP9t7+ukM2Aodf41
w3QGwGXOq0blwNA27krMpPN193jNPbySxtUaNOfBkRNdW4alS/LRbOxFqqImwSc7
uAWpONeQqxapg8k1xXjUXAcLBn0P7I+gYe/yTZEh/0NAz8yIUlY/ia2hhi3UbOd9
dds6WfNOeX3/AN1gDiTqFxSWS3D7k8Xv4PUAAI487ZtG5l0hUm3wadoD1IxVVSge
OAvGmREn78se3eXh4OvbYQ2NtHF1FS0/NZDs2gKB3g1AzusLPgeJ0o0M65c/kaZi
T2pLDQpi184jSYMjHZyEIpZYC0eZ7duoAHVsgtV8OVfyDNHG3cyRy4tc6/mpcj04
N4q0up/t0gJYrdTo1c7HPo+lZ3aqgiXyHldFxyceSneo1Pkti47dTulRw80BS4tz
C5/lymkfJ7K3G5+WLMKuij27qfQMKVGfZPirEwd4dUhcFQzlAX85zs2C//xKHcfz
6gaFG7E9RZUlUyagmtONqXPL5SSKHO3HC40hepvx2Wgzs+6dsGTqUbp/ptODGrE1
/hnlYqy2HQowM/ZWRbu31W8bDP6iBw5HtE1kpEq/xB2Yl/4EAuNxa9J3v1qRRtVt
i/GkXOS1B7ojiM7rMhWXE7+q6i/wqmlzbo8vofVU+WZg0WzpfsbVnxuqYKfa6uTb
OEUte85VdBDX0nji1EdH2fiMHnxwR8acdB23OS07KmaNLwigSCsNL/AzrOmqyUO1
OOPJ+EJ9cWPmWM3YHLDV+uOD4VT+w4oULVH8G26j1s6Bytk/9vosDxmM1wqiiNaC
mseee3WiAfacDmbZ0DO21QJEwCqMihKAY83YZEjiwnOP6uZ16m7zCz2ChcD/IIK4
A/X99bNh9gf2/oO0rmPoxeqPGKkSrxkwSHXsGxuE8nAlqysUKpnmIemP8GWXMwWe
E+wxQbmtlxeax+85u19eXVZiYUuegwCPwTJOwnfe5p0Erre5HDxBo6wcteuS4Ca+
P7TYywKarIxdAoPynevCj60pz45oNCZvWS3GLH+d6wQJwktUgV+A8R+ce92l0Q7S
IVzH1kUxdrp4RmoGjtIn29cBWdJQskvpNz/ISo9Y7NfRyi/mgh4RmCv5eNhdk7VC
W1X21yLygRwPxcUY4LRKyIJbwOhp5hjOKNbpExYc+UYsMTrXG8UYZi03dHaphWi3
A7qVdlLH6uqaIAyWMPCZ58YV45oNL4yv8+7vZ3JoiHZfVqQKP/DYYpzSE/ag11eU
8C37GNu/Y0C1f/bDXk2elEZc0Xv2IAj0NmE3GdHH2V/dpeKWttv+7fzxyQH6i2np
WrVOlPkiJV8DyRwzR2M5JT+0yBYLhXTX1IE8lJDTVS6LZwEBd6IV1biQEe46IerB
0KzDGO+cUbvcrNEfoHqvsmBEAeZCrC0RARHQGN4OANz9wbB7mF9xKxmSXrECBSJf
9saTwuQWphYG3H3RDup6qpWql1y4axg/sTriltW5nQU1qYXUNhQ9sNIAnNv7IiNy
yfYWEbZQQq/BqpWUB7h36QjURziF7p/5y+RIJqjQxi+8Txg9FtucB7N8wi5YCFg1
fdKYC0DMQS/E+6xQEtyRzMEP/IgU5ByJ/I+b3WlHcaOAdFTDCTs4KLHwds6GhDaV
4O/A5Bdh02yQi+MQdKN2S9ICAqSsPqLRRbt2R7WBmccB/FdpE05uwCBySZIUsxBy
ROSMcDTPLajNWTsfn3Fdac0fyhMFYBWe8xDfzbYsELhvNKxiJc5AVMno/aEcSKOW
ErLNHwL3TAT/veX5TPM5rcBh40W9CYrDxAGo5GzIF3QprCOucay2K5Q6pr/8ToJr
gPwTs6sXsor3tAdI1os5/qtwMSvyA3cvREIvT9drhOsRCMnaOaMUlkjJjzd4Tzci
RMZv5xs0S5DaFPcz+Rsq2WzDqa+A8F59xThXOY8RgxQNTlGPXl37lCvOVc0oRHVJ
3zoG8qoRZ2G7LxEAyl6eok7mNQr+DJ8PoTjmx0baLxWgN44izLCdp4viF1noPLay
Cr2i/mSWyeObqQVsg8GfLlgUrkxJwBVNemTbElqAVVZ7bf4iOjI8M1Nx5tORf5PI
Y3frjydOR/oFUnK2M0W1qBER6LaA/MfH3FC2D0JOaL2Zjn0x1A0XpcCXEQmm53uq
AFkm8aUw9T6h+4qh2iQtRk2aFzzZGuYPcwbCXRUm/ebc8TIJYxIentTgsVuKg95h
4J+MgMT+TDfWOknXXw8zQWrfkp9ZsEbK590Uom8qdQfUcd9sxMXFWhg45KlxwMCT
Au34bs5d4p2BcxelofN0U5H5/3xhnD2Tk2Mnrs0tjRrrM9ZShD1waK9UPwFt9TF5
n+5ZFW4C10yBKw4MuXiHkg3sh35tp9KHdZNjuf3gSKey0zm7sSYJ0hf0PL91ZSuu
jpjMMNY32BDosHYxBVVzzN1ygszx/4KOqWrKvj9f/d8DKN/AvcnSDP3i/c+wHdrr
onay9Cr0RICef5/2FbEnQ7Y/CpI65PaD89YcKRpx717VOiZYcCN7/HYyxSAOfQMW
xxGwaOQMcMV4rpaqdTtW8AD2jPnWu8KvLlGrOL5ILexk0zWdwEhs+zA/daPy8tkz
iUXVt8o2cvkr8OvpkRnARnRhR8q6zyn51RkX4nT4N1c6xw1rE2+I040Bje6IoXSp
oijMQbQ7bdsmVLchZ5Y5Cj7qT82anmjzOmKTJP7ADsWs3kkAcLgQKxhqE+adCXSH
VT2dZWVnYynhax0s4NKfIKOvERyWU29CkmSve5c/kMmVoXGzwv/ctGe594Kk87m4
18mLQc3wTqDaYKorSRfos5btu3k4jn+wwGLWl3nmX6AQWxUuprtmIOpfnMTBJi/2
8KV2aeDSwx13WnpyPbSZ+icrod6BPP4+WUKjCNr058HoJTGgge9FTMY0PByVq5Y9
so8fKuNF8W/ATnbOyCE3PgBKYzNtovLo6WmWLk3qYOahWpWG44C8670YflcQOxC7
Imqha6G4gbz9h+t4FGa58zx871pW+OT6X7pIEUTDBt1RrqoaXNogFMVPhIf4PASJ
0xOCRujN0R7mcApK4g9sp+FsfkEkfkQesq0Yzo+nKCEtL3JQrArj/4L/ZuyZFiRg
7L5mjcQv5SwSz6AUm/kQ4oBbvs3Hyysk7LzCmarKjRjVrSdaUBbm7ewjNI6D6Ma9
oJkcNdfyo61c8QyCTcb8XH0etUvrYvo0AGagIb7E3whrqX/sisdvt0ipfB668sRb
s1CkpxHmq0uDtw7C0MajjRLw1BA3cdSqUZQlETrUn+wxCLDrgJLWf67nAAW76HT4
NGbdQvh/Sij2eLk1lFwdLlnKtECLpoGo8GKhdQu+ekP+jZfZHXXf7YoKbPM/DCGr
kHRcrgUJM+ylJom3YWo98+flEQ2zOZGNv3CJ+JupmpV69mWg0FeQL8YR+qGvKaso
WFhSmLWmFdhXiSQuPI9iuTdvQJSsJTKMc37rkuOMesGKEaaH+CSwVWNkWTeHHzol
QSkyX+TbhEzF8RCeMKn55fQcuCM7WT1nEPn+oq83HoLJtDcIkbV2zmBNvjkELS5A
nUeIookb+wTLirr+wenRYyQYuTX62r2OkpzQxssEd6CmUB0OFYCiAnJWzK6ArJdF
kKInFzSe+qbR20ZXx0gA5jZfHGDSDp9OYBGHjB9PLNToxLdY/50x6KxSjtake1rD
qLu4Aq+nYuNkSvDNusEM/bqh8QQWmtrjzUnC/RXHIGnyK7fIi12INYrY8bT2FvSC
/O2nidvy7xQeX8uxtLPMUmKFUBx/uk9QehGEPgodStNja1qTgNKRWZmSJ+MJQYD5
WSIj2FWQ/HqbJjiTrLDHE7N9zQYgdORa1wzTeZlYFmAfsmYTI+GmQ+uxUuDTlLsk
npsi21ABpiURek+CLm4tOYGPY8vLNhN0aa4qiHRX9XQiCGMGlTf9m/AHY0TIxZnm
8tXqzZ0R4jWcJ/VDKhX0IyQxTuU3UGjxVDa62p78UWxw96w0wSbUWJk01Ln4HdDn
v4R/Bsbjc/cIV3fJYT9J1zZifnmyuq/Fse7l8N6qYQsZhHvtNRbL8w6YP4lBIGUZ
gH1SSrPZdLkrRjhsmuHpYgRIv9zZmB4vt3q/DcYXjD871dqgQx5fS//7+KUqnRDe
YP3lreyhKEpFXfiv0atBdG6bd5cm0A/Xh3dRCGb8k7vHXOCeDCy3sZ3zk5B1KvVs
Xb1G4rvXxt32nI/0o08FhFCbSBgKWVJUGOvYyQ4KGWsx8BWYtIzP9XeSyq7o7CBi
lqDuIeT9dhFoV3FjBHH0/MxjJRH3soRBwRFgRb30gZ8WaJfwEVHHf12JVLDsaqc2
e6F2zHEh9m3tNAjv7DXrTO7f31MTn41zrbZxjmRT/NsBCLhhHuMV4i7iskvCW7ka
N2vSx5s6f11nNoLuhDfNG209f0WDjLsi2qPlYoQT2lAOrxvYcYyNJxb3bRZwZjPm
jxuJFpQakj6XCmcgHFv1VJkMeJbyL6NVHgvRt9OKF9ITeZKcP8SWtM7xtYbMucam
fc0cli9X+r4+P/UDRb4lbpZwZfMu447M2ck8BIJdKZHn1BMYFNr7Qy/pYRASamM2
6r43V7YOX5cvCx3MSULAipqQWthRPccAWI97iW6lMDCsrb8h/bxUfOJVJXM0wGON
G2JYUiE44pLNppXGu4Fjx3gqOElEKh/DVyU+vU83cT1LzOTkWNe8MY1NQN0GG+qK
RbntyQDXLJauUOVBedZeEvbrn9Q11BZidA8dPx+OcJJJKlAnm2dtkKXCQ6l/mhku
Yv3qZtzWsK1VTXeWvzQ5ssKTJiswA+iy0R31G+EOsMWOQygQuCaw/AZYytaBkjj6
WcuxRaRRM1qTgOG1dBuHhTMIj5rVNfM+H1cphXEZd0mYCVf3Svm6+e1d9WVWWJ7F
O3+ZD7BNTfpU0Oo/mRRLjMevyjtQTbx95PEO73QulP8DomvJdDV2n2osoHCZmQxY
BkpDEsY8SlKi3+kjYftF8/zn9Q+g2CuLQDEh8G4tLgTunqqc6mWedsZh/0tclaQU
+B4EtqOFoLrxXPrEtNfy0u9MMADx494ufhR3lQ1Tzufns/nDMekvfwXbAQNFmUI8
6VAkUbdvoXPhssavHLQRxeG1Fp0Qyvcw9/knrJQsFTeLDlsc7Y9XCtOvwiLAns3r
567z7TBk7w0ZuRHYMHIPCeGba/DicBpdmoXbcRCtAaGVlWCOsq1OQRH51r/sawGX
1ZZ2JiZ0WDnzyvxmBIny31MTf8hmaw4Uy04AmdbkWIR7hwgngEJ1/oMYBOo6cZMr
srwz0uyGFH/dEpEg5LMCICjaNg128wdam/dLNnHLyoUL1tHmEHbUrpl8Js3aOUgj
3Aqav96CoYeCPtdfkio4kNEVMb/7YeHJ65PirGBKMKtSSRL63+gvPmL70yPCKUdn
DMdF1kogE8JadOPoxhQ18FSeRHaLoRdz/X6IrWsviMc3EpWeYGNc97r7Us6SOhCX
mXCNkdIKyKqGaI5xvzjyKWeYZNRZIczW79+A841fYSR7dUX7NMKj43MBfIB9IIXf
J0yDIE8WOX6o34sJ43y60LJX90ykz+nBZZEH//r2PwACtKCIm5J3oeeSvyNC/bwr
m4iqhsKVCQn7NcBCCGUmnUZj4O8pfvNZJ03PcTxQA02Tp4NKb5tOlrYhvPqBVGWl
oPCBcPUhfiL6XlJuLiyMQFdYNAUiSOCkXM1TXXaZdk0TwqcqC1l8y9jyc2gLtA8f
/6lAdLWFGBj/usFOPYNdQkqVZG8zYSkWlZ9EkCdzo3UQnJfFldRLll90MOs2Ukol
jhLiy9QDLfX81WfQ5qYhlDRU9Myn/9ER/gv3I9hsdmJCCruYvaSBXgwY9dEWlxhd
HQuYLtPTO1f3oTQyrZk96Nq+8zAIcKC+I9BKimQPfKiO61QgtIckDSc3xCLNmgIr
SeQsTacKtNtl2HCf+YiuFktOIUIXBLvVqkpHRo3hVjQR0JN5zOmfYKhkEN3GMbHn
US1SThTNBkdsXdwArszcQWGIfimXdrK/gj0KfVs9xZ+mQ+1nV5GMfb9GYYWOpHLS
7ZOtG8uOH4ix3gjZngTnwYH7FYy2Zx5c3qNrzPh9hsR/joMXVQwftv6+7Ww3oQ+k
jTkXcmVWLCbhZChgtnlZG9JZjYW1sBFZXKnh8yOLVSfhsM2GYERtRVGrgF1UJ3ll
ylP8Ookc2a6z0XVEXxpN3aySXUN2lsc6P0SPGkcNofML6B7cdLHUxvoLYU9M6K0j
7K7bxVlT6fyBvZ3L+wZsTmmYOKS2DZTnSmOL5v/akFVfW31ikLopA0rYaHQARhJr
WW5sCBIFeoARSPsBWNvuUcK3jEGY1yUoKaLfRYEAbTHiNQD5b+Q2Id/UsB+50Cud
Wx0+MXkxY18R21QCxcJRTwgtXubKYBy9cN7OFfY2XPEv8eyfOjZljsfMnWEO23//
aYL4Ab7r0VwWJFiEb9hz6q6YPc22foG1Arfy6afErLkTsBQolLiq6P7XScJlfTFm
Dysw8qOS0+0sGZdMAvWNmOlsd0larl4v42TvJ0lpX/Z4Vq7WKG0K0P37Vd9X7nmt
Cb665geWu8iX+mnJmQgwvLODjNjOyFy1zZkxGnqO/n44ZWof6VfW1R/ONKjCOqVy
d7JM1LmM8STq7IOyg3Cg1ZCtyHSF7bJY/XYo/t7FjAZh1VMM+KAbxp00aDWA+PmV
dRVRTwLjn4ntwOdiIkbS2bMdEXUxJPqqcDAjkaIt1f7fXI/4K/WcANsjJHZSd4qS
F2AxljH1sI3Z8CSPv4KihV4K4JGZOWvgZteLoc1RBbWaaduo7BQjmB19/nTaK97O
SK96yQgTHxaxUquaHEs9uLJ2ZJYA8XEgIeiDTgesZYFIFiDw7CM8HLDck1R2ZLPX
q6GB5i5GXW5FgP6RzBnplh8g2DAt+jSSuO+IvytRc1UC5aVp77FZrUqjEpTdGI9f
W8Hsm7AeXJJtHUYvitK1toF/a8rQit6dxyNQtxoBWDjwA3f6h7YJRwZ1FVe6OqzW
7lQsZZseZLv118fKuKkTCGifO3tjAimbNFJDBLYtr+18mHfNqJBcoNgUFIitloiD
S/I01YU83xJyy7TUELEa9o6GriB5uGWm4dUHZ06dcJE6Jze5vBSqDXDqlSZxNafi
QiEJU9afmZbCZ4fUJoImB8vf5ZPoGyjwmM/tVYbw1ITsTWNpgNiXGam1xSn0ynzE
K3E3gOA2UfwUk5lDaIUHOPxDK6wJiN9eF5y4HlXnLUclDvMuHsIGCcK2VLqxw0bC
eo3sa37OFwSVlA2zC9wQHcbu9zr8WHCiCDOxKz/UKAw+QauOtVn92qTe1e20GI7h
9TkvSekLhewrhV1XLAN7jTOTAJaxPfcPExuOhuCJ46H5bLEkrZZ1LkjBKhWGUZ+q
pCeba53LAl9tVlDKAa/pf0A16NeZBMxnXIqHSghH0UcTcP1h7PTPortHHwcsHjtG
quUrJIvi3tBUR/ael4sq3jr6VGYhrHELwPheECq0hq1CdKskucazB23PVqgkZ2YA
VIukyGfKEhmp/JPILFt9MIfIADpTQajz/OsJpxoxv4hmbWPQvLO1ZZSwgSCE5p9n
UE8llMOJipro9i7+swkdScAu1OqSX/mk+0DNIu1L/VNnPLJLc4JmY5pC7caXwIew
p1uKrjhUxtg+1BgT0vtj3WoQ1ELDW9/QJaIoALj225evxDGjlse+kYqLj2IMgvDX
20svAgEdaZqW9ErgfGIpm5zl1+pCeSvM46vsacrSAzl8cQZXL6HVtRY0vW0wB4nL
iU+VcJmBkybfYNSmqWZQ6PW+uKzXEUSIEPqlxtrdlCpF+tWjGqYekEfkgvdFI0tW
HgyOIxJAaWlPYBENIHhT/lxcy9DAS+VEXjcSovNQBmUbEbZnTFGYJb7GK2f79Cdz
kdVCyWiSyu2lltS3ouc3A/DeiYDscoUq9CQ7G/qVyGHSgMeaPJdI7t9DWmXgZdd9
jTgH0HaeDDRmEsXC8LPNtzQHXpuE3nS/SHyxMm9/UpK85loYGseFQXldC71y3Obx
QOTfzaVv0Dkcwi6XUio3VtipDx1LEnFJApuhw4B7nI2Dezq6AgkV/WHV7Dg61Jgu
kVVcpVtqKGsZD0SoXtisB9/1Qv8F/dLrPQcRbTSnTrN8jeUFvhvl0WwDPqarnggC
Ym+L2OZWK251LqTRXzX8HayBDCLbG94X6H9Vp8W+RcI4ZDeqOH63QfZg0BrUIvcB
r00bTnViCiei3yQustvxjDuu+9i1WZR2U38+xFHCBfLeDeYPlPA+UrrF4SuHySqB
rPkZi5GVI1WaJ89tD/UR4tkLZHaBZjouRacIMGkMaGUEMb4lpuUQF+Ua8WihTvSB
hkbcVu2If8uIs6Z4Rz2nl3BHDjXcoI/vq7ZwpQsIZ69Sgpgiblnfa4RKG/NR3Lq3
rCNZF4lqFcaWpuRPEyBVxJY8enBv7suLVi9+mkv9egxarOVfQQaqYTMINsQLf3Zl
MddprwKPahYigLDlvgYGWBDQd/A5Z9kQuDK0KYw/LxUnrKEqPPfdGcGzMDr3bS3G
h0lNx9OtStA5mMqS0EFAujJYPDiAPPCBciGxOPt7sU9nRF7ykMqrl7S8AjW92RpS
Hhxm4++jf/vTjwYScrf0tY441G9uqp8MN7izBaxovdavnrjoRGnRm5zyhsxzwa2R
FufwrAPYXoXXWQvT78l74IMVMc20IryKK/UTXLjTkf/rDXQ/OTbLeX5C57IPEcmc
o7Zmo7JEhBiOspxQGMLPjBxmbSMUDBYfvI5ulGUNYicTqf9matHrlpxHl93kZmk7
wikQOhMBVEINRlVJ5GCLOJai1JPQ5pMN7F5Z2KAT11tQOh2hpHOIphwAgVldMZv/
NMSplJYFePnbXT2wJ4L7jxEMo6w0ZrothuDnK9cZefmq1uqKnPFBd+k9Z7E5yvEY
zjx8OSuxz6nxUtLjl6lMVF0IDgtacH5ad821wSvZHjzklS8nkXePnHuhieob/QuI
z9Fv1nLRxX26ijtiOQX4RlA1kIeD7qmKjQP+HychN++f/m4Tz9Iw9sYEwAsNNPHo
wMB2arWq0AKl4pM27noie6YNl0x31+7csJALSYWDiWEOuzNzN9hTzi6l11ROJxCL
NVkPvqdxHDxtSGN7XWa00YCjUraZSLt6Uec5JUBoHsYv4YRoKg+Ge5O2NAmNzT60
UmZ39NEoQczyZ2sl9+fsDSx4sWU+t17OG6mr1ibj+HM0291hjL750hx6i0V/M01w
WkGQMnU0RE9sj8O3f0Vn1Yc8V8BptN3ZFI5rqbH0YrqfLaHM+M2SF8RVN+NcvRYy
dMWF6Xl/WZZy30hTn1hG1An9eoYAx0tidiALujPAgsfn0jFLoy/0eY+SHP6CTEnG
MAhL2n1W0SmFPC0Ax/LzlKVAop9AGIHsZ0LRHw8HJwUz/ShJJlcI3P4aHqlV8udk
/XRRoepXmv6TG1w/wGy8fv5Yk15i1GbP+dfIA9mUgCMDRvWbnpzHCshMqADVpPHp
qBnG7PKtQ27vXSyugx1ff7SIOWTz/T5AdGYgGDwIZgb6KOZFSgYiMVeqENSrfbN1
+ZXPCPZh5xrwPzU6lRzgy1/bncvZWMX1kSeuVjI54y1q0Q0XaqBHKr2bYdRDjDoA
kXD/m73wBqJUJFn05W/6Xwk8NCpRGAv84VmnuR1Ft9fphwavzvxa7MSMiIe1lTB+
UaMfygbeudDKEtP17h9Ko44vjSPRIvB5AhWGZhB+IVvtlN0Hdrc1GE9Gp+pwDqY/
H+k6OGDDa+aDpJ8H97UjOIVwaTG2q5wntbiZocUvLcc/H/wCj9LWZSb2qwY7/WY7
zRaj5y2GgI2J2+wqw+5e1K9X78x9ktMV19eTQQOWq9gzgsoFeCSTAI4jPZVR0xch
f/VJtRPimDecdOiPd+1RIVPJ6Z1gj8ncux3hMgHqc9Sjq6IOnyoT6sOk1NaGg2H/
8y3TKBDtpTWG+5H13lmGIFLbYfFCeEpOu1LgG4HNFPujtyX2ZN+9r7BhlshjbkMA
E0Cm4eSBuhNt/biZo3nxh05ZoLAg1+kXgGTtVBVriYISDtJ17Sr0aDR/nrNw9Ina
qLg/5ZjV1w3qfK+sPqsYfQ4QJ8r1igQ7toYtd3KUyj5aeQw2XS+q4KSyUKyNSOif
01ViszAtI/qCAWUuu/T1L6TYvpAR3nTu8UbI4EPJZSbReQXdTGlXAnHvmN3m6GOy
Yt/hNmz0NUH83+1W6y2DTw+84xEjIV07lR/NEGU+9Fw21dafBUiWygIcVVNwa0Cz
c70gfF0WViQeD3qeca/VfCQ+ch44nj2BbBvmDkVnZATfWAQGKRJQw2BQbnafds4J
pqH38xg9DsFBEhTXFP9y2M4QfE/xTWdiE+2kfb7jgyvHO6po9TDHY6YK4KLRYfvt
kPkK7k2xdmiqlhgWGAkjx+yySuVNo/Bfd6t+h+HuVwse9OO29vGlGCCkP6nHMeLq
7dDeFZRdK5GhyEJl5OQ7Uk5MnvEJ4XIZ7n1fhFt0eYAB/vVC7pXvYuboFY4BoUYY
Y++tLq/xvAIyX7wKA6wswPPE3qAGltN89GBfr3pZTzgTtAr5Vd+Vv+8CwKp+sc6o
pTzq6RXhHMIgJMH+3IhMNgFHwzsUBklrOmN/QGdxM520jhsg4EsK/AN6Lh0Qkrlj
oQG95BZoAy5ZKOHFyH8EplWYB5dzx/qDO0myovXpsbOL9nGoq6G76tZhb5skTQ0/
Fp0YPz77m7aY2pF4Wcuy8etIitqERR6ykhMvXNvi2jtuYkoycj6A3aaUZyYLqP+W
rUzw2AJiI9HwgsXXh3iKuzNsU1F7g6VhYSk70J3Jr0iEkgUnTj+sauP38JI/iqX1
5JKuXkA3+GzbzY3yxnMGNyA1tfeclbX0h7ZJc5XcqdzRKTsjuc9hTeDqQJSFvTCc
SLeLs22TCT1QPEkB1/czXMJsViEUSMouP8Koo0MgZTKmfCKa9SZmskfjzgvPFLiT
9WVo+VpCpUOUdjmVOIQZmOFybiGICOqJRTGdQUOhc8QL/3vGzFCpSYHpHnMO0CJc
0e2ZwAYKvjEDbZzYXKhwTgdYY3JqELzT2WQXrcsyQatNI2ANi9q7yMagN/F1xS8y
I/aG5ENxCQWXazoGw7b79a8AnK233Z5clu6dwn6XoFZZUlXlIRnfw2PRlzLrsNkC
aJMkEhf+KjFf3dQ3053nLmtt0N5XAJYyZpEEBD3YFvjAhlgsHbqIGsorPbCU3dt5
iAdP9gB1xj1bdKcPqq0GmAH+yP6hSGRfGkqxXEemVVBXdtGhH2uvdxh2GQ8CsVmv
vY4yEADefHV6EX5kdZSlOoSmvNLpRS8OlZPYE1fs+vnYnbQLSsirBoXcXcPPYte9
2SS04MtWdjfLnkN5kol3FevkfBCzlhUk1+K3xz8MRn8whvscXIDSyCbz8pJd+bqP
Kjk9JSwWrRxrrCplTz+fMpkFSb9E47wD867REinrbf2pT9TuyBYwYWv3XgSqo7A/
xCNeaZg7Q5nD4weSDIyW9PX8TXbaRC0Oi/haJV9dxecBzti8RKigc3wG1xfWWe5Q
VHpKErL+WMfLLvuIxVgMgfWjCbKm9xiYBIbOtGp24rg+Ami/TrW2W2PTf2bInDcY
i0x26EnXiwqLo9Op6ajl/wwDzWJD1tOmaegRlRK9rHT4LNSAA+S7zTxPIItmIHj+
bTLunL4tl9jOTjc5y2cq5Gfpp6l2LjLzP4uL/Z65zLJ61XIva6dG+uLAWIeownv1
jmX3lEntZ4b+4YHF6emWXfh/MQ77XDF63S0ftb+7kiMKqjUUHCn+hIoQFwHK7gFy
khlPP+d0XvDTaaBjf5BfeqJ16pTUVS9EVNFrYPpKycrzSGgKThdJyxkoZHTp4Ysn
6xBsBkbJ4+xDgKsZAoG9QvmtT4O2MVgV3gugpUR2HDVV+Rju0hvIz8bjaqWZYcHJ
R5R+pIROMx/x0ozUi0BtjDueNLd47Kl/KFY3VRoDiWUaztPs2BBJTHFKM+bMjxei
OvxvFoPo8l5kqrp/vdwbKKAO9AEd5vjoqCwLnBUaw6y1GQmMwwXR2w/ab/VHWkw9
ENlvfUnMQHkGtcwSg909eRJBJO7UnkARMeTxpwncOwjJpDb00rVztLyPcLU5OcLo
OMZbhN+481IRyVMGwT3nwfHp2zLzHoLX+c9a+XvegKf3ILYEtGKVYQetG91nGcQW
xL2kLvG5UAHWMISycOnaBtvQYZlhEaH++VCQC5OFFGplHFxiddmwoYbE560fuVm6
5FLfVgunO9I6rHNgxnNsJmxRA68Afm6rrX2en1k78QAj+W5+L5dRqRzViq6El5eI
kHy5l2Sts+A5SENu5NBOxNts3/fqlfCVRFUi3jJLhZ4+7lv4njWN3D/na0Hn/hd2
IRqROBlA9rMcXxQmF81X/uJUo6UG6kIFJ8JovpQ0GPoS/pKdUn84Uc7XvkRaj4Nj
MlRRe8X0NF1SgT69nBZjTgLZvti0yowrBVJJVgUbz5iV8pcfz9lch0R7BnS28dBy
IH+TiwuCxX2r+iT0MmGawJuB+94VwH9IF3KgIFXEZftkgQakjSQ7JN4L1PCQLryO
p7AJw95bQdfbEAH+SX2/yyairHM7mXZ1NyjP5Gr+cudGor+h0rCRRnmSqKIrRdvN
cJZC53zc3IgUassJ2eTdc7grsI95bKT7Hiod0D5tc9/K5z1MHQ117tRUS1fQ9zLm
F8AyjsMhD4ywMAOuQjfKn4XTFdEakiqRD68GiD3vDd7dLxvmfEB9+tyWj3mWzCjF
DR6rzr45dMewHrZFoRkKzu4XxWUvBZNpa0GtTmCmOufLAp4IBiZBy/OpA9mkSDt+
stbP26el1MRwOvRJgzvoDKhd/x+E0Q30yDgwYtV1RmJOL3pA8bMipu4eGG8Pjejt
LRTsHqZbjqLx3HXl3X8WvISdvXztkUE+FokwHhH3nTWONc20l3C04EKDC+H4XGeA
bZQHtXh46bXndcYke/bM9BZ0sE8kfmOzUTAdCWX9ruVhyNSUQko87YMGSj4+QAW2
6JoKwlF0ZlZ2TCFUWDO1gKs4JCOKZjkHo5sqF1TFNss1RCPHTfINc4EY7wNrFE/a
Clz/I69GufZs7YJUJqliVKX9LBX/OGumUtjipq/IGnPIZGuZjIYMxE2TQD1KO+f5
tO3xVz5Fh5Ggo0nNaPoEg238icaptkyQsCr0rNP+KlHRMFMnwh5otc5bQrcChesz
KeN0Z633e5jSR68UqFW9SmEYx3z5XwVEhSpHqJnzAY+bsGYS8s3WlSbLGOul13Cz
4IRMBbSbVM9BAJnTJKyhKDakiKF9bhREJpfYMWtUW5q5gzUyrOBIlV3bpxJfxpuX
iv2UhBpB7D2uhcsuvcCMoaScy3d/zlK6sIqkqMtSN+AmQ2Qmid+1TDLgkDGomdTJ
Fu/8B4wK0diBvoY/ONLHx+Ve/6H5G00BiXWKm/bp/KGWMLiZ05sAgYcj4yfYhiWo
h0Vl81QB3fWBvAL+fkpZChhHpCKnY8aNmGDHUb5wSGgC+KZQY+yI5ExoCHHs4Zvw
xc+vhxhTIEZ3ZxdgHMChp+42DmgqjS3UR2E40uySbSf5YVzOCjLUimlT/EU8uHo6
QCxYrVICw67lghK792MoYh2g6uWO/5xTXYyFNfmdqYn2ImeDeqoWbrSmtfknTT/o
VH0sY75I3gpJUvtQqH6j0ZT+OSQHX92ZvhoqNeWPhRZ4Sgpp9eklSuxTlbuHQ536
WTWcaQAzELLXfFCRgudKzTVWOCRS5oOQtMuMOWEFpiKDmtz0avSCaPhUaSaeH5rP
bSpVZucG4i7nA9F83wpxgTM6KzycGB8cl9qUmXvkr3vJBSlcABAcgT/ojK3zLi+4
P5wrzjpSGTVqVEeohAhX1foeMqYcFWC00dOzAXIQXAFHqqTgMusWYHsSCR/Lq9r1
ZCd5VaLv5lTAYEIsivCmCir3+ZMqhRXvej0PleVZy0df0nBwZDntZG3HCoGxLb/A
Fu2IFcw+U7q+CwJQ0v5GOy/0QZNT02V2oPfbCOIwZNqdBhO2NG3BZFSCJXm7RP5X
RDRENSHxmuqdq1LqmfKadKsW/FXgk0DwYQuPRIXmPYit7lXi2s71UfckcP1PXGks
a6OEnvsp8P4w7+YDAHLfEa6wWbpElTLzMyVZEQV+bO77gnoWeSgENqNnCzUQihIO
vg2KY2TY01ToLDeCHQOD0Ht51ZH0Q1WeTL84yvpoRAoJhtWW7NPYcUjPR2kTiXE1
dHGtj5nMAOuqPiRPKE/Y6Wi7NsORqYKnxMzWXpqjy9svMIPaJUzx5a+H039FvB+y
s6p3Z46v1clW3ydtXEA0uNFR1VPD2LEm6znyoNLr47sc9Bx4NuRC+qeRdgIad+l7
3scCBAz+zVVThN89S7Sa+N7QktBuGb5iGryZEBg8PxvDKIDpsmCLxOfrwRCIPG8S
WByRBGaDaBsm8AW8kpIw/Ip75qe6ol5lpKm0CyIQC6oi99nNJOS3ErGk2E/X7DQx
tlg9ZgqN9V4Bkd1Ne/j8kd/8pIpgfPh4AcMVUs4rY+YVGWUc7YhA8pz+dkcO0LvX
A6ae0AzuHhQ0ZSHb8CqiQKP2c4LSJWMc3fD6MtsX6HSs4ilF8QEA/dwxw7HOGpqS
NkUEl9qSAGJ4JiakmqSogqBGh6dNbsD0TjQrKfy8Doi9cLZpKhQlDkDsyKz5heCt
k+6y4jaOOLCMPkwX2Di6h8ZWmTZHG7GArhSXH226khDBu9wHJ1TACS8zR0rlxdFI
mZAxp7c/zVXhYiKqpQDPQPgVKgJQNXO/FEoEJdRlZFxgDsUhyW+zGnVHoVwhVpwm
IfuYMXK9XvBZlsLDm2Ri4DFertXziTwHF518xZ/0bVzXk+rM1sY2Qj52kqXQDFdZ
Q1GlTwAALdtyUXYN722bb4GkjSzYy4t2OEa0gkfkeqxKW32azGlrGOi2XELOWZzM
y2ctjv8niGQxi8uOAC7z3b141FMQruGt/UfWg6JW7+rK5vitYma22MtlJsNCDnDw
6Pn/fhfQBSthnAwMOkkPVLll6wqm1FjIIdEDtQQzKe/7J6PukJCqlQv7w3nxIsg8
rsxwe7ksVh0u+ZuFnkbfms3oFdYDpXnY9qZxWwULFd1scOivz91nopEjF4AelqJ7
1gQn4+rN3dbhmrRV8InNH/0Y+eroYC1vifEH+cWSsNPWRHQ+0VFpWFkwCQuDTYps
WRx48UYcAwjfiJTXnPeaNkD9tx2xsbd4TdUa/RNeyCcIakAEbrKT2iwxuHzzrVKA
pv30s3nEXhe/aKQUk8+0TUkO5lmDZWqgZDcAOQ4XAt52elvTnjRto/Z+Jiiea5+T
339yKLpOO9S5Nwc5vCUs1hWdA2rEiO18DL2I1j40HdGF9oIpAZpfUCEqsKsSJKsT
Gp7P6zDzAm3AC6UKsfqnTXouQFxaDZEqYBxIwegOcQjRUoKjwZrPnN+7ebeDnUQc
7wrMmHzrT7UNcFECRRysfRrJurEhlk1nbpPswvuTjxwEcu19wQn5AI1vjgNVk/ri
rdzWQ5g5OV7q3KV+167f683XfUnmOIiiBaZRcEKbU3Kiezn+IUrDymWAmsyEo6CL
nN/M3Ayj2lSWbIPAAEMKX9SrWwWsu0qDjdNnAvVs5ZCPEqsSFWBIanglzkUJr8IV
bavt3hqbKYDhb4s+e7lFbDG3lfPeg30Bo5czZf1EHi6upkHYof8IlhQCOwunpgY3
lumoSZPnY7kWutPwluyAiCNVfLYS+Tk89xmtHuzB+Q6RqM/8aHFR5R9mmSOzykyj
Gffxp+zxn/QTg8Ygn3ZdS9DNGLVokHlxBrX4f2koXuOJ+8+akrllHbw7HXzW0uFQ
cn6YNaOia06Mp51qlXbKbKHYfd2vVhi64rQiEzP0kt9RuKVQ676eMJnc/dvaxJl5
tkg/9BplZfkeu+8UpfzjXiFe6JrqGu/CkKO2UJrLosNPzs2v9yFqss5uQ96PQ6gA
11/zW6PWHCdtTXqzlqY/CrxYpERfNSfEQ3OhvZIEc60zHAAvMqBiNPhnihD/Y3Ye
06cgsMuVgN3uXnCExOLoiwvNx7w86xEeeH6JTUrYyW1m/DHUWhZx82UYe3pIL0sB
BO1qsAhtqhKj4c4Qj80iHtM+9zZSwm5NxXvuFuoz46DIqEaWo1QpQwN3n9UVQCrY
22jMDnz7LD6iUcYEjeGCsH7TnqlUuL4kGki+T07KCa9nHsOCkhwkcpi0e4/yQY+4
JGLQJ1/v9sbtOFaoJe8rqtqbK6Me0DqG0xfkCDVZ/rcmGYctUdRCk/DoFj1yfTW9
lxA/ONR4+pz9dqCiFxrt4L69AIQouOoFeU/NKQwV7cvVTILeDDpZr0VZqOBSB3PC
xs1nV/xhUqPAVOMG2EPGrzTg2Kc4eF4gPsfAWRKRGRxz137eS30WtcbptceL3ljC
TCKrp79rGvTBEmtP/qDHbf5T+evCq5b+K6KA3X0mvNKOtBjI3tM5iDgMUt6yzULK
8gs3BGE+2enqI1xvRaFDpFSJDOmLvLwBvm3Q/kdh/sMexSBy61lpOrsCeXSRm6of
pYcI1UJh4KRGZxMtNDvPJKqMU9aDJ0ZzmIrCMCm2sXBLd3fr+lLO40evpHWd7vT3
s2wu7w2pDwZvWRr8jxZbulViOyqcubuVFZbe8wGJzsxLIbd0xlVy/fkZP0txhOG4
k6b/YEvtQGpeatuRIJwBiIxwNoawMK9CorzAZwE/LSKAl+f03pykKAC+5IA7iFVs
gcFBURyPEiro0ayJ/WDNV3wcC3eMdfahYle6RwKnLPDXATNAhAyjWc0d3oRKYJCw
j9tt2anflMm3erJjeGKG78fTLqToMPdXIo1XmFcMIfxr6Ju0VSCaTXCEUt/Tp5V7
dlLTCgROl/YOoWDJI/58k8Lu3e9iD6PtFOKOPcYbs4TJsPcZ36YvTt1pjOx2XVhB
rkyU+QDbljjsoErmTyXELmDaDGBwPk+aHfVKfuONsPpVYVbCdW0sSXzIHYF9cpK+
DP2lWcjMCKJNLaGaI5b53DkX3dYVskbqkMm+cmCEpFQ1PjRXSHxU616bmg38HV8h
Ydy7ET57reARcfPHGkOOZASn6cDh/SXm25B5c6dnd7uZIoHNPcpGhc0G8zkMvG2i
0uuBr5ThiZno/yT0+0WJ8ns4gAqPixYck63Pw0Ko8aoDJdE9y+NwDZTJVWCAzHt3
SGADrLACea4ZbxEDU7kVDYGo8r5EIJ8/Cgs6n+PhEU2wz7HvopVd/ssuRW/yPQ3O
ZlPLjsOKzlQSyMhRDDn4SpSKkCNUuRgu5s/lVpKa4xAY5lhzKx3eKEZFolbRHyI/
lkVqlTs2lz97zpAWY/KVYzgeIVhnnnWDdghw017kN77g5yekWsbBWXagDWfGAmDw
0OD3/rP68zN5vda8EyypFGutcoLEo/2G7F7OmcVFMpP7rJIpNDItSmTHycStUc2r
2V2FVfnFKZOb0kekWcabXKM4SSbaX0twgu59RbIlDWAjUpb0BDNXqZth6cWjfMI5
62VXLoLSlHSqORtaROba0pRVLIJx4UzERnzaE2vthzva0KCbvAD7CxCXC9zr2z65
MxXZfhaweZE6BF7+ml6BpK+F2/6vprEGJSHek7GO1WI+0Oi1GT5SlutCU1jtinrV
YVtZb5Zoxm+sG8B1w0IZDJ5C70hL8pOiIqdcPtzicCit2I0dhTAJOOo3BDu6Ctpb
bKN7h3TIUghLpH4mP0kmCYKa/TQEE/VX3EL8ktHQrfBGs5rnXd8jhhxGzHeUJ+SE
K5LkH9Dgc3Y5y5w022eJVgnXF0z7tejcP79rD6lgeCnvoWNs0OQiCtpLT5M6Xs6g
+whA/tDdc0Yhl6RgvxBQUgl89Vszci7ggkTuRmoOeEmr7MYzB1JXjPfPHxAm7pv7
V9LEGdle6qvE5qmKHCSOCMLu7/eEvuMzrNNXIO2E2GAd7cl0wO2k8BkjxHRbvkaN
1LP/nD1PROEzRHMOPu9tI1DY/Sf2by3wQ2a6OgOpPTksc6DGDxEOiMMaKCbt4FNA
dYBle2QqM43YEyh4RHFr5Q==
`protect end_protected