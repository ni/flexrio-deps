`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3824 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
HdytKcppDjja7VfYQkCqvHqziOeatjVyccN5ahnpdkbuCY+icUbachxiwtZ6rqqA
QF1xd8OeCAhzBF6TA1pF/zeHBfeGn2c6tdrd8zSme+mClamLJVFA5saO1qbqihro
FMZB/RgOYuHJVqoQ1kCbfGAIviFEyces2ZRum66p1X1zUQaBjrTdX5wQ6N9maDK+
Xv9U7YRGrsP+96/2jvIpR1VfwXQuneU95dKr+9eLZwiwZA/lX4KTJ+2giylQq7gG
huuefTJAn237pZ0mo8mwZlZYPgFWwODNeRmxmkyM4EiovklKf1AMcsc1b0URT9eB
7j0WRm++WYrXkwWHsNXEbbnT4HKBoTBfYnaygyWI7xESVsLVaZEHMg3fSca/3git
902tycvocNBwJlWmJPUdm5P4PasEx1XTmxKHDmBrByN4vJ88BFfu4C3kmGfW74gP
Vq3JzfQh0GXxck9wXZ2bfc4PBebTEavVaLrofoEIwYLzLYuSjfn2me58aHwOhMLZ
fIlcGfi5KEd2w7ycsiAX9XVbo/aDRUwduWPoD3V2csoNVAhNef5WXvk+SPCwFprR
kmdTPt3bx1ghwIdbt9fl9oUpIhBoZuBLWdO+GsLxg5r4jNGzsDKOgrWKqQnmComN
THHPALsf9yVwQ7KDBR4hCYikSh0CxZ6lypdpN0r7f6mVvpfbHewLLYYV4Sr80bOv
z2Uk4EEPhF6e0w7C1x9L9e6kHHz/T+8kUAjg+nRGgjCVgUAsIfas1fwC1sgolT+O
TI6bOLu9fIvMrn3GdskOJ83kRQr0d1bSNc7RbEnRkJeYpxjIXXlBHIBNakK72XnG
ozkm7SrNY9mG+ADV73xlBitMTYtGfAho5r15u6XJzsWCVmCOkfGs5eHpglFeoSOY
dTYJLdhOMK8Gzr00JnY03G3T20QJ9zWPU+50eSqj3tMIF5bCVGW6XYzbTI8ATdSG
VXnRMDStVXp7I9AMmcSk6FBrpuQtrv1Rsj4ygo/AdlSUp3heapOtavqbfaHKTDK+
XLNA2EkeVbb03+PKJaP82IU0ROwD+c2EJKvzJmq6gUzNoNDSmmyh3RatAPl0wDLo
p8+2cjInt1bOBQF0G05kR7cxhLwOppov1l00eBnxbO+g/rFPBiUqt1dfgLG9peN1
UA+IhPXUDb7SQuce1pxObjw+bkX5x/JWTWs52xesT7wkAe8D7Jl6IT79EBNfza3G
QMGFFSUU7sLqH3/lUuoV4FPUT2b7J+LWkThtEXvEMKWbJ+QE/pWumy8dNLmzqx4B
SgnzRCRThS4w3AG6o6ssTWK3uioHNtVz0z9nd67u9YRJD81Mn9qL8Op5uXiXm4cG
quKhTkuTk+VkZ5eOnPE5FLlss6rSQVwtlCZGU2lhZuIlUYztFfU4BKGQyzmvT6+j
V4hnpyB7tvSQ7FhFEclSbhajesIli/590P1ZdgfvtwOH9zEOYoRLWaFl4R9w7LSI
dCSpAy7nJyh+N5VfV+itZomjbbDfM3rO31K4cR0Fnz4jTTeMJW3DGwkwySsYBaLX
IG2a4LV5Azx19puo9DvKBFTTqE1YLRNP3YFtGrzqFwXQt+IDKECkcubSDEun4FoM
9T2DW0f5Z52k2U0pRH2UnN+zJ6+W89cJyPEQlCJwOJURIXA76xj7CNBDdLJ1istj
ACyFs8Vos2KHNBpdy7e+iOoMcxjFAo6LdPUfmzDtaD6zd2V1780ozW2KqXJSHaI/
MeUcr8VY2DcIZBHSupx4daQKtIDbQAFHQ2nM2jcK39/wt0FA0xV2KvARzFKQUtKN
Jm1LXpnxered8Ggw1WLy+iOP97Di36WzNGfukwhwED3ksRaCceHw6rgoLLSj1qlm
383xvcXvVvmNAhFwMFQtltboY+SwvYAqShqvVo15wqh9tP78D+vTJHNtXLofx55w
sacxXRoYvrSb5hIa4UUiYNSDP+FB+TmlcDeIhWn3t7Q11mIvXxKYroGw6ntsA3hk
HNnkqc6ohrx1pQvYnhShPeCh/xiUTmJzri4UuY84LVTcnGCRMLtItEnBiZJjx2Y7
Si1/tstMl0edaFTSG5m5O4wo4SlsS+KPkGEBDh2NYDjBsH5JgjTGiyUTv47Wc7IB
CxXFpCD8UqJahGyAOXXimC0S9PTTPyz4sFzuZ7R1FM/xcWABpYZIBzDJGhFxKNfF
0KqcsN5U43G8hShXtQgj1SIVW/mcqR/EVVdcmu402ApA7QVAquwQjbmN05MbZlLS
iMYpsuvXRc+aCBbjcVxGOHkzH02iHotMqGz5V4qN230aciuEOUnBAgADjDoIcmm9
kMui7StCOp366DMclaeLkQAcY6s4WFAiTEYmK+kIQuT8XdBA158mWythY6tbRZ/R
hwg+/RIpQFqshR5nXtnRWIw0NJoHePMgh4p79kIIslcysyAi4Ys+T8jaovW2zcpF
WgxZF0lsBTzbI4xkspjytpNmfc036PbiZyHiG62I8c3qsM0uqU+8PsX8CVMcau66
vhLnl8zYarxfSG09nOn1AwTK4x71+c6/R8pt4xyxnBgflX24ht+QhYYB9oimm7vr
J9ytWVXQkXqqmFSOKQa1UuuZcLI30QeS4nhi4eC6z0XD/EGrvrVfvdwWKVBwQH8p
t+RUmf7K1jEaYicYheCWTbJn/WnXaJtBjJ+/6izok6QWNmjr21kFrCFeJ7zhdCey
5j0J1TBYjM6Lcns58HUWMXl5yHG8MKNwRhYB9vXTeIx9Oprkz+pSNBDQ+jgvj59X
/N7BOOiOqu9Tp7vZkgD8kpyVzYI+s+TFWYABt91a/tWyLWQKJHYzEomiCeSJv13X
jaKBiltXI2aVOoEq/TxxuNwmRSfD+mFRaOpkaKbkp1v1vyHhsScfmPcOWca4ocUf
sNgqF/vVKtso4N6ApuO2WuKy8SddRCqMz/ohdsRvmTL+FomOhoNmlRh+1xYMLG3i
fDJdP/ecfo1r3CqqI+zjjmx8nMIESuooXiw6BtCnR+gDi2pKXE139jUD2LVFwzVV
rAvx7U39TWJ68rtS/GLDB5z0erymZbNwGPFhepKfjDjDkuyD0rqOqlKm38aBeLs1
LD2Ug8/GkJgg8r11LvcuVJgNDVZH7LSXov+ZZ346PcAxdEC6WOfxQZ/gXAlc3VTq
swsiOuOEQh8iKkorH7xVZQWd54Gtt3iDaY6s69oD7NtjWhvNEglI+W0IDFBaVtHF
5/dNrBdCoLyu9MpLN3jzQ7YuENVkLYPJbqOedrXiWfwreylzoOgx+D/wTJaykjUN
DExu+mqeA/zemgMrYB/mc6Yx51qvzK3lKjRID+VxNu9qXGWHKAN3pVrl22RgCF7B
YyD6vxSEX61DUUu8bjKKlLJAiVjci0wu4Hsqyi7lOzumAWGcOYVrqBvFvTocVl9F
FUDauvP2zU+NTi5pxsxPTZUjxZf59WZA4hqPWfP+MRRiXDTacz4atqffuHCzHKDT
miDm11PF7XpUqaYAscc2ChLGmaanYVjyD+j66ET4hPkWhmQQ1nK8KW9qKOJYqeqm
VIyIqX5bn2IYfAPnuhmbYdAjsQ/iR3ZHopdXF57kRQSTEJR9ojzBfeMNFc9v42P0
9PUk30Q/4rqB5frX0A29nO8PhbHVVH0m7GE1/Si29V/d1dixiuMwPyTnaOsuCmYq
Oss1WFsu6G78R9lIKYZ0EVSA1oGyGAh1A1NRYJ4OoVNww7CiLq7mkBs9v2hMrLAj
QeETtSvdwpbBWICcftHc5oJhVEktMxBJqmNd7agsxLe2RQgpEp+yi19YRj3Y/Jno
AklE2wgGWmdcz6HwNoAqKwYwjFHwUVuQ1ukJxnUn2CQzwhYoKPsEiY/rTecb8xQp
EM5ltNBicvR7TUKl1hRxa6oWnPySx8tjQIsLTqmAbY/HkgHYsch8ghmKvyNkwzd+
8zVvm8F2IujwFi7YOWTOWE3qTEA8PtW+JaIl+w6nP10YJBs9fQ8ob4WmSdirbdyj
rJ2+9FNo25jJyFNV5V3z3C6NVaTfRpyJ9W5jL73i/bmIrhCjS1BFCVnBDmYnobWp
O3syrjvhiyxDn6D7d3fTtSKS/eoNr0qNAing9bjS0ZQWoitUvG4UJRmI2hVby5yz
f/CKVC81hYg+2SEzxW9t+qXrnn7kiNWJa/jsUJSElgPLYv9RyqLmvjHImXBxChhP
mUYiwFh8M1ZufKi9P0oqw9zUEO4UXLyYp1uaNJbPt6A6m3vPdZ040WGffBGXKw50
5kOtd+47M2MevBP9jIsa9EqEiDhC3ZDumv7sSaDYEqJapK7V9VQH/mNsl4fsAuX+
7iiOfiPyWJM+jaizOJ6tvECYAfwzXlyahiLtCgU8XcuP8p4+n5gcRe/EBONGWMPX
a+9boyoQGbEuqNtBYBUBuoGuROTKXY6qHmzwfAFcH7rKvZav34F1Srli0d0dqVR2
7Ds5rvimUsQtYvYiSCYgJhZ0ho50PYz7i9MGlylXi4e7L3bIfPDgV9Gsdm2UjKHy
3emMCLqsnSlF4N8BbTJBBRzqWLtpFR+dMG295veAYHHoMwwbNlsZA/G8vpHI6yKX
A5LxSKlmAGszV+RCnbfeKiwC1cv/NtqQo7X3tWX2JqsYq+Ziq346zH1ZTsFQ6xy6
3GXIpOymBjLdjzbEr2a8AelPNue6YCMZXpRvADKl3qUyVITTLcnvufbq9e6jB0ZB
jZYzdKkc5vZRxEDcSHhuo4XEhCeZevb7B1qanLmkWQ857ykeH6s4EoSjo2Iqf/09
Z+JMC2sb0WzVpaIRCbRpSJz7yI+T+06kljuNTGs1G6mSSB0E5CvQ9ZEfK6mqbi5I
H8aCama1ao4ENv+abHZ7/d3K8ALeQ8zUM160g9wh6qnuPybv5+J2IfbacWZHntXT
gLmkH0PvXoB3JZwnEu22CySZHKjpTwW9YFvQjpVIuFcaNsMXy/8EHwFj1xfXLtS4
3GdF3kr3LusZVHjRXGVRMBoRjGs0heG49Gl1wTUaCQM=
`protect end_protected