`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
gMcHP74wBZczB0bB0IzoP2xg5wC5NPjD/GsvSQ6VQgzYAsanETMwwsWi4yhFtJwv
5kY07u0WerSDf8woJ0stqW5xF501W3JLIS8KMiCOd55RHBOnavjYiaaLeu7oUCmB
TtTS1R4sO325rP2zOn9YwRbyyS5Ljn+PzFZZUmkt5xMca3p5NGqKtZW2dV6Babni
5HlLuF20Au601B75m2nv+ZRoGSrpkNElxoTibONmX8gBflpIVE7BehhHwaKSucEF
pp4QQ5zZAZjEC6aplZepouGVggAulz5AahlX5bf4opOVlB1J7IrgyjENtw6ysQ/q
DzybQ+ipztSXBGhmcCVU3A==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="jAI3OJE9Sh00Sic4PtM/KZ4WjwT98XM8AMZrZsQkxWQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hyw9IrFLPQsjvXplweG8O0lkaSLBN9Ijv4B5VdTRt6ipKJT9Kzsb5LxCKvkQyF9n
sGPOd5i74hRHnkHfYISGkfxGJCa55ieOyFShOsqTKRLxclm4oja9vTIey6yFm1BZ
54IDCG9h3PqfDiTD847UCSMRvFssyycwv+BRHQMQlFs=
`protect rights_digest_method = "sha256"
`protect end_toolblock="BnLuc3jxknmZOyxfJK70E5kp9u9O8IQ8cgkXv26kHA8="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2688 )
`protect data_block
xABArkLxBOK6xG+7CdOOiGu0zbCbHMrEntFfAZEE/xRFxZaAZl1QLkuFI77OC2KL
XxG/mrHJzO3taVHgwRXNLDdc8ePbxbAiQfzV3NJLBO+gsBjmIymaCa480cPNpHLx
5QrNkvfaeGZ/VRaPiTSh5EVH8M1I6okjx0gQrcfscnz/ZKUC5meyAV3q0pvI8QUP
yZnqpcw36FdLPG62YKuL1y2e2CA1+mg+FCdILSkz0r8QmJv3VKFA3qx7Bp26p9t0
RbV4q0q8bAL3COvMSodjL+1zTVO3ea5K1Tr7y+mBsrBxBwBAFxkPSIcLtBEsGL7g
o+Ly6izfQ2d+hz2hma/iqjYLrI0Z+DeyombIEg3dkR4zOYXkQWXYXz5IDe4NV4lf
5TC+0uo74ztKhQTdomW66gxN5ly1KcYH2F/a1ab79DDbRLoV6GOQQx86SsZ4OhUY
XdPSUKRcxovCw0OtzwGJlixq4aX2v83J1aJByGG9uR6Vyw0MrSQh82L5/N+NvLIl
nLaITqgmuE9bJ+80ZtwgkV/S/rfR1WcsOumLlA91OutaVpL+vyh4kD+6aKcFXyzC
bunKH+iPk4/+wd2/za9TWseulAQ8Iy5Jsb+P/ocUWqf7LE7FcEh+u3qexiHdz1yt
C+UcTHn1Wc2pao0nDN6g8tKMQtSjxT4fJvIQND1cpuGQXk2yuemNfaIlCyXuIhRO
+gGggoWc7aU5Djcld/2fLmb6ovF9iwlKdhLuh9uIVehobTpHcvqwoXuDhvu6d9ly
pWUT2Qw3MDkdF/EvNMFU15U8z+b13i9lmyq5lkPrbvfIRKsHC0HRG9An8OGoHNcs
1HKLekhU/sRdT681YJKDO0hJtDN65wTPS6/GQEMw34w4MYe4vpEbJDmoOKWsr1tl
J3j6wINzYHaKVDUw3DJZE/9L2EPaDVDKEtwTxI0NBpm38F9Ec/byKAs4Rew1CG+r
oYTuw9GwqbLrTqH2+nh+NkVRneJgO8qXA9lWDfKf3JK42mQSbWk4dOpoxyHTWvcd
9nAgqmhOvHjBG2O3az0jn4xphITZr+9merIgyKJ7WXYFam1khpdwQ4c7uf7PcLXH
WeyZzt9sFRQYQo3H6Ku/OGcoaWA07oyM7F4iwFMEU6SQLfwiOcI2Xkp4eGkvDO/f
MCZQNFkIMuK2wvIC+jKHltVuPWmxzZ7MxmNltt0k8+n9Tha3Ewefwwc52jY37HC/
5edQmpi/NzNZMwtoOHCm5U5FwdDzZP9pwUL8uKgjn4tE3mdC/6p4SA2/t/EL3mPr
JTDTo8dcbZgHBY+aJz3pFGx4Qkz2wzvR5Gvz+fMV9nUFsqnr4vT3RSh1eUzVxE4U
k2xjyQkSOOwcC8HrnE7oB0+Dy58KMJgIPjsjhw0e4GKjnOIRUV3wRZhKpw1sV9+W
GYnyQJkjGdC5vpVwPNPDNx6i0U4bPdjFlhEX3lhepNBPInvXQekQasuYddRco/qc
gOZVdKPH/Lk/V5j7SCsPH1DrkO2BwgwyN1dRWXezfqHfT/7fv/ttjXcMJxTVpP74
uooCf8wafiWMF0QT7oZN7hu9dY1+8lClLUXKXXAWmxbLaRCCfdU0FHuJqEjVVGXZ
DUbq4kLLixhnCrWBZ73uwC9itFK18AKK0njHD9yCURJkD4GuKgs62bcZgPRsEfjk
L2M+wVyY28dVOifHMBAcQH6dfa35RnXLBMo91/TxN3DZ84UkDt5r20fB/RtXHSXH
AoGd8ItUPr+SH25A5ontEWSyqy95mtckQwtK9uNbjmxN2F5cUG/PNGVsUm8YSyKh
VMmGIZVIqX5JiGnX3MmIQX+NNvAFBM05f/atdEXC9glwXMeDNNaKaAzp3BA8b/ys
e8KGwhpzjLpr0S6X6JLNkRJ4SJJU2P2jxjkSvd9LCGt8uVGCiXRtSXDqJlYhedcV
bHgJQVpaIAcvIjRuv54uGtH43+ek7Gf4xC8h3WJ8RJwEycQEhmZIeLJg8O+ba1qe
VGtZVCkPJY0fefzzU6w6ca3bCQjBI4dX4pVDsge9yNKvgDjmqh6NXzdoKv2eiMKz
jYEOe5F5W+Y+ZZQNPzx2TH3m/mDKxqJYZjdnB9MeOHkRmhVLOm/56P3ey7JH3I6D
X+F4/7Ftxda3RU5Q0dRon5zdmHMRU1x2Erfv+1UJGxWA089xPLqJcA+0Q2oAPspU
CU9bGu9v33jGL0S49ElyIZGK9X5FFAp6uYiJG+FpqJuxRwx741Kc/uUuNu7P/KP3
p4faISF+t/LCpRPJ+Zf9cEtTzgkbUqFLgGLg7RMuaXLZnefMlPiKdZfbT1Sg6T67
aZn97J22GtB+tKpQl6lO3NdMzq8dMqGyPFJmBXQ8905WumDYzw15zN99CCah3wL3
0htlGnZoEtdm3FrDsdgGdQrf8btjRuEij+wAdorImzXoLCYbtPYzSxnDbpFziQar
zXwWz0FxY7XVQdaAhYz7L8+B7zJ96VjHpP0AfCDgMgK7ubl564VL8BqsV7RKGb/C
cLRoHjtX224uGclX/4miLd7T+AmZXhunBYNW6rZUWR4f87XGhCKk3KYLboXFUrer
zEQWo0QzjdyaJr5pHVJlKCt6fkz+Zk6JZmvYNceN9mqMUdEX6Vk9xv74zbOVPxrO
OtiCSCCNvZJ0I+RiUx9kM62hfl/hoHJuV9UNLxuxBPfgD8ad+KD9bvbs/ODZcxYW
TQSydjUUEfINKxnlEAxJNDgHTaFKP3xJeoW5KeNKM0wUFe3uoSuW8xJjYbZMoFCM
P7nZbjm14A5aJqy1o5Gn+zBtK/DapK5H0HC4d/qWjBa8X7gpgRgSVZEh80Tp/sXK
M2cg9k9urpGNJD1dJqYHsgU2jQhrjt+YLJW46Gdo3TqWhXqt2grMugK+d/uKOuNx
BgSkg0ISqqy5NHbYtqmdUWh38TYGoBB/p2pSWBecnFCCPw6afUt4yuF/K+ThnqGL
EVJvwEexAMPUXO0ygqffpc6lbiw1MNoqRyYEVZglQsu55j3T+UYfmXzb5ZEfAw94
cu2r7Mmu7jblPmvNhg3sdaf4K3/yuP+HVMB7LFcjVPDXZ5XV1YTjY2vyvtLDWWLU
dQNnFw/ZqwYp6CaoMslteD4PV2uF1caEY4Rcq5dFq3K4EVyWA5quRaBC46JY+N5U
EolxE87AuhOy3B2FlQfhohULCfrzUDrVjU5Vyf+GjW1vvQ+65KlblWxc9W2ZxI/B
KYMm4C9y/rm076lv7ZGrmMojosq1i8Gn7Gvh0iCrFeC9zNYroJUZSpuf773wyMJ0
dathLJdh3yk+h++DXtgNXp6rmLqyhTh1MiPBnAoZfggRbDMRrpicpyTxZ99lFgQE
UG5Wq46nTiVTw6Gl3semmcrCvSOXpbRKNZjpq/W7C4F6Jlg9U1ro2jtErt40hCLw
8VYT4r0PU7UvLJwK3ycU8vVf2Dfs10RUNzzhlYZbUVRTyxT0ahjsoPK6yn/Q1bW4
YdlnwXhCnpqWFMgm3Ui/8zl4IoJsFuhM3/Vlbn+C/aJq7NN9MxWpscgzZUE77rqQ
fjqFonGqm2Q3MIR4xdFl/Y8k3G4Cene3vROf0Qg2ZZir+ZITuVrWEnsXZWaQjRkE
`protect end_protected