`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15664 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzpmO8K0c/7WUi9nFCtYiO0+b2qEX180RzXnq33fhvvtL
/LEZjuYmWzm55ouoj8QRUA0Kr7KP3/FrB901oUa3MO2qmA1hIrIwqcWqPder37/F
vgToDFlZbW+delulpPiibb/1+UqBvdUG/ok4hHURBo6CsPSc05iG9CpY3JNSXM02
DTpl5Z8J8a/zyOnaCO6XT5RleG1ALRs+yqPPNX4mavu2qB2PfL95sedZckK3WWxz
pY5oTpeSFALifx6++bX5+IelP58Zjhl9zpknSZmn1MHtzquAysgcSmV3/LA1MgQq
uicUIV/KQffgDkT8OYn0yAGVF9HXG7S5VAr99/M/rxS8kEv8Izc6lq1lcDeM4F6z
vwa8Orjo4NDc+kpVuxZz2HJtt2D6sgkdASlmYB4YQ/+pEPruObgtKuOGjO1ecwmI
Dw6UD0cGJnT/nvZ9+0+WHVYQ+9xKPNqjk8VviDWLjU1YMQ/bk0m350BqJHz8Bb43
Wq/dKIis7ZtD4TQbnFGfm8/U9mzWYlZ/VgqLA526iKUIHJhPV+5Engn59Lq9G8PY
8uTyZvxBqh//+tQaEwDVsovjLvOc/HdT1XaPIyhUlOza9LZNe/c9HVD0JW6wWQ2t
SYesQFRqtSBPnXI0h0LbojX0XkCYdfq6Zt3p3l8xkfSibnPTIISJ8XM+58gS4dlA
8SFmRQdRAU6Mb9CruCDrxhivffUqPESytmcFzpq4UfK5Om1Q1XFKxXKa9oYxJxW1
8eDOirh8HJagWJK6VSuk2RCvRXVgMQPb9LWfH+KVqzpH8Fz3aLrjXXGeZTldKmGq
zcT1lnrPg3jA0R4ivSGjG/gXGbvFcTpksMg2BFixXcsbDBok8+fpTLVW4pEAL7sO
hmUugbFrOZWdjODtOZ7CN/XuDXuRF1WzJBlMNIww/hPPGBJh6tlJ6pZgyWPt1KsK
yOPuX/rx3MxCefeDt0o8xrF21/aL5eIJPU3f927aenTlBP0kJYrFbM6Ewh1bN1VW
F+U4ttHJCxiQOWPUdagEBYZamcJ6avX9hFoyLbhw7LVQgwGdWo8fMk6+Pc/nybb7
5kQqc03h1z+troMBss2CfLza8/kpxV5Smr8+DAL5OZbt0ypzVSk0rkwcOs5niDsO
OvINzCMXcuxqBEZrUFPH313WYwl0sh/AlxGFjwCmlnO8E0qN9gm52M8o0QvcdMPG
zSvG8Tl3GUHMG18Qn6SHlb6KKi8pwvKlp1vXKyvvypYbx/4Qfro4e/XIeGww43yB
WNz+moZQQ9lwJJ0YoSEM+Caie6aF2gRnb5vZPgamOA8TasCBSkd1alJc/UsBz6CI
PBvDTceKhdtWITjrL0Wo4OzoihzsK6vUONTq+vE5zGI+g7nYVsdGbtFLpJbllRAe
uFRzKDDXysfDCZTlFan7zi9s8vpCkuB/UZ3WTfQgV31mcRExkJUHFswBjzI5zo1O
M8hn3cZM+BzZTnlQsH2KWNUFiUSiBDpu9/1oSMrZUQTTgQ4SWrSlUPubyvJtQoLm
E54PYrM5uwW4GVzJpZpll6tgJ6GLfkW8PPeEcXMrrIxsHcsV2MlZgX+UgGP6WITk
gfi83Vy7QBGiFgW2kcTMqZd4dcjK55K6Rt2XxTR2F5kbyUi/83Ym4CpbUgKReFEY
YJ9kikD5RIH5uD64sr6Ljrl8r1uLEKXjZr+RlIYLu3lcelINwcy7LabcI03bezFA
gUNCjelXNpaISCSsYfD8gQJ4CiDqHri6acap6MqvwblFj53zhxajR+diI24qsp2T
gOdD+1C88LY0JjP4eilXWpLXD1hGsett18MBx+wBIzt8ckkf9+pEfTH5+M5MBirk
igXtauP/YBd6QQAZdXI2zgQNiSmbDhEanYecrrdv4FJVe6PF3sdKX6yKvJUYHaH4
CswXaLIEslYKd83LbukyCbDFxjjghkXWhfjg097xM/bHWKzSzyplPHrddtOo/4Fw
58kMzzl+XAZzy+e5qd4YCQZFlB4/5Be+0/8CuKBfEZZJHvqIB/nA2FwpnOOpdD/R
seDSLafimw4BnnoyWLkparGTo+g1NuuePfF7zYt7MLHyR1kvtaFGOVTc/b5bcyfr
7jcRRmmmqNARA9aGYWHaKSt8MYdrGpToFbfuwAiD44S/YeI5w/c5U4HH+dyWPdF5
9A5YarGZTrN7ozpzWN9fSvpN5LXt4w71az0Z9dj7y4Q51uUupp5Kaz5Bmi9wAfFF
xlHL6xdYByq2A5b6brCHXvyluD10VL4/8huAF3J+xPXk/fptRCPqNhoWbgxqG1jJ
37T5ASXGJEMpJ+GEhEx9Kcms4SRKPFjHhZGhdD79hAXxgjMqEbJ4oQPuKBrwQ1Tk
qxeLMBiDV8HaIa1TptBpj0nXxb4HHG3LFJucfzVNljWCQZ0F1q7DTq1q2ZM6YQ4K
fos+d19N8cipy6VCru1VSQHsT2jYwLJqU0Bx+h48pnM0lmP/ZEWZZP1OcF6tmc6f
Af8MKOTOjdnjw+ADpmkDasnWGUTeEPMBy3665PWwwWE6wlU0WXQ2Uzx1XOlX0Zwv
zQhbift63B1jYV02+vfNQImpwDVxvDNL4XdXy2xsvl01BzZBky1dHwb44NSsL/SX
h5QvZ40dzYyeJWaH5u3y0XZMfvdEMC+LQz3ReikI3tSY9OMqOSQpAILmWh4cL05e
yO3Zdl6fTLEXp5knH4U6W99jySW1M8ppxJzIiYvNqMYlkbtwuVQHQC/v0OaXsuCs
Zz2dJifY81eqYl0Dc43tOhCEyqWnl9z+moDYInTQM9VBXVOX/wem+EsJOCyyMjfy
G3SxrD0NeO6fSF2eh8icgU3Gmw2jkoBr1Mjl1Xm8eqDRpJgX50eGtAW/s6kp35ru
sDyrXl51ZoUQ5c2S8gibzr29N1vDm7ZD+LczI1kebDfsTLubnDnlV0LKkNyWBPan
XaSQeWkjLSKt2EGjodxoyrcnaQib09elTVjbnQDYmsvlt1Cu3WEuk2Cqw7cpTx+9
LFMxbho8ypUyW9gXpDx72x1HLM0IPkmpOppR5Nfmy81KCm0P5WtO8WEGL+cp45ly
zjf6rjJ7IMmEyX2tK7f0L8pjPmDnms//Yiav0fCs+7PFDCBhUwgWIOAs7oEY/UEp
50r26Bis1huibMS7FU5VGcrHA/mbQajDs2v10ksyBmh/N2kPEDChTPs+bcV8jmSJ
yRvPUC+BRyXVpSqCqLNtSdQr+aqA5SXnTT8X38wOWGAgK38IAejdOlK962kSeSXP
s7G1wNMDVmcZaLNwR35NrBQQ3JDWsflonL/gZydfR+j8QT/1uq8zWyDRRmOc1hge
xKpEzuFXVYG6r0DAajGTDhUaaX1/tW4+obCY0vDj+6e8uULT/3pTXX69XJ4JqGW1
X4vC5mcYXP6DvqhZOkBb+JIrPE3nvGcczU5cPAS9EGvCfEptf73V4oMrQf6tIpE7
ssfufgtkcN63gIG4EWKp7ODkq/kM5zmMSp5CqrAq2nvoa7dDeVEAlKnulI01PMsA
kiCxZIHqpWU37Pqz4uqYzCJHw/8RneBgX7NnhnmfuiWM1b1Vzm8m+v7fvihxO87i
xT/cL1Y1GswNW+9naWN1tGTcCg02mxIRNyjQ6Egn64Yezr2slTx+PVzuSr9C+ebg
PUOz9i06H/gDG3IudJgKUazduglwKTUmlO/KtLewEkuY6jMQ6eM0cXuLsNH0lhwN
kWtTST3Zh71Ptqj8JgMw1KSx45/9jZeErRqm0u81g7rmqVXyxSqV6OI6Ba50HcbL
2fm/rfpGHj0C3AbnW41t+pqxmwV/9Cbaimfpl6mndYUsKc3M8w+02SDp7o+8Y70p
fkcKvzKa+9C0UOPE5/sIVor+6WZ8/QNT9QvQxKTUFL5y8NAHel2xd04o34PQahJr
Qr9RD0I57Xc26VXlDrBNpuPVT89lO9g75Xa8Kc/GHJsu5QIT9Jf0Suye+iyVTf0T
mE9g4tCuSV/kG4k7WLPcnNRS71WcunR7pnOugE7NfLO4o5GieyKlq1LngZnYBAph
Y5rSrvZKLi7SAGVFJT9J+jp2sLWMYdkxkqLOBBT/W2HKDiKR4ZG2OVedsjo42Qhr
KI3qiwMXpsONYMJ7ToVQGm3eD0TV0tGqEVc5qkY14jKAPjgpcnyRM5cbvz8/5oQk
43+4Y7mEmjdPZHG1mU8FE04xU/Q61ibuVd9BnY07Zwu7QlJAnLfHWK/aYHNL0Wh8
Hy0tic7VxDstjBW/dt1yMZ++5/oKt6u9wBQXjlyPAUztGbAfGda2kiiYdQttCk12
jsa5xKK9YWdeuOW3nqaeE7bgjLAxbb1EwFXIl2DCHOXElxUSRdfRwEAzR3I4JTQf
9tDG2u+JIEZAiWhkYxMVjUoI2EToYxzW0zDs+WMKbkyGCIdNtMu6uD+ImsNpAfxB
tUn7r+qffLMcYviDpJFj57h5FdCSClJ07Y0p0sYGkkMToa/k8ftJStz4MH+1UsjN
Axaz9IM48NEn3nr8ghzlb5m4on9zo/ajb2dl487LXUt4AEHGy1IENYq6dy7j8FPL
RAkqgntBVmSK//ckgxgIetTE+pjo/yA8WVs439FSg2YMSTCd3elefESSqh8sATqL
US4Qt0tQESD+UG1h64m2EgL2fIRZKwwqd1bB4hpltkewBZFgHf+a3mjFgclo2uhj
+VqtoEWqrRpBriglf/9zUWjnV/xTkmHvTKmnxR4pQqYGD+Zm0yMh9dXpUP/+frQ5
NIFsiqvTBqrSuM/z5OvfPKbtrPljMrpRsNjf55oBeAOqE2xOxkS5MpURpFQzNuuB
NJaVoiwlIhu13Y2SCzCoGhiIXTTopDfplWHilPUC7ptGPsE33VAa0v7iMvAwCaNo
gQOZ8MS1amudwi0KxCVyA86jD3A24ELZiDUyof5cw3LpDOQe3ukfi9iC9bqM7UDc
DZ/noP7vxHghYesUKvHrxDYWyBtT01/oPT+UR3rgV6MiKziNM80QcTbnDqrTTZ3a
1u8FUna21oH0QzUOH0HqwsOWHdiVziDxwOiOoYQ9CNNdDZHR/uLd6N5nn9IhsRzY
bdi5ea5rfEQVbTrz9oRHQ66/Az8S5RHd31uVWgMaS5hh1RY5wExbaEgdQaAjVMME
ao32OG8juCQY/Q9UYolfWInhrmPDZ01Aml4UwkUcbQbLy8YTFR5JEH9E2nm6vnAL
1EGiApwxcLOPk++tZvTi0aGqoWEFvfU8OoWdPNP2niZBf9+rj4GR88y0gWJhwRHr
MTS+MrY5HltZMd+CghMc0cP7Vxu108prQyTv3MzMIfUkD2QPfRDrd5pnhGQFVXye
iDDeoOS7pHePq9ZOjoSaJyN+aEdhCWSQwaedckD4lk4k+72ES1Pv+qVwjZPKPoTM
y7m6g0B/Zho0z4Sedj9QDfA2YN2YNRtOj+rUB1W1yKJfD3Nv25plBhdBg3FqkYnl
QCYCdSJrBTxT+aGWQs8iFDvFg1Z5XCm9V4wi0YEGEbMQ2gskg+vO3lnDyafqS8O9
V7n2Yg7epifAtAJYLmYKpywCB5j12DuxYfIQqQpKevNtjDHCq1b+YdiK2qsJXZDq
EcCiW7/UbxH1vg6j+tNIbwDEG3nIcaTewovCFQpTpjN+7lswQglcvNFFXcwGOksi
pmWXDslOf52M96/M82N/uy8IChyjpoOcCnbCiZeIDua4aGK9xZZ35JySfM8MlZQP
gy0ayD4R18tBZ6qZOVjWCZkiaCNnoWSRO5Zn9Qg7VGt3RMGe0oHnPehcZRhm/Loo
lJzDtouHPyVrM0jvU+g3yQdEj0hf1hCLwbrKMDc6KMRgdVWfGEDP2cOAifU3IJt0
lZOyV/ZW4xXcF1G9R+MtaII4VuZqu1WTweG5AK5ndNdOxqScrD1wAUuklCgRC+J2
Oa828VWWkP6pM9Jrqm2cuLL4+NN8V/D9LATTsJInoa0fFonZYGHPRHoHHSqjrIGn
EkAlKPBmzw2RRsEix2KBEdClko7AI/pHDma8P3MB07Rz71IZOzRzCTAf3LdroHxb
6z45A5tacxNbBOT+RNF+iIVxm+hd3BY97Ir8FFqygBd2ZEL6CAtJr2Ow7CymkEEH
Q7GnHDoxWVJt2quchf6lPLzeZtuIg92TtZTD44VCvr8fhmxbkHvn2Jk9crVS/ijY
qXOnaFAfO6Gsww69YKkZVmApJ1xJgi9US0mycwVwSRgEb3Gh/QvKfNzJ12wjHvGL
FlfwkyvxtizT82n5Ik8a28x4EAxxCdQI8BCppQjJzz4Xv08HTwTrMxsd0BvtcSEJ
snvlQek2vXjTPcfWaaKXzarwt9LdcFN9fUfUtHBnSFR6pMiiwEQ5dxg9eLXcKdIN
mwlmPvmhWPbJeNNi0uhhDlXH2k2K1rO7JLEF1Dogd7kaB/H+xd164+E37DDsqx1F
fmuxvTrvd8FLMxKqQD+iw4uuMhfxU+LnIm/juDGls1/d5ibjYyRFSIqYY0Dpcu0Y
AJ8vE+LdrLz4GdNiBMQy+Fsc1v431B/cQZ3YQyF99rD7SGAuTPxKoQp1gJW3+FW0
jWJO2+8LatpBPsN/k56x13/7qivUTN3yxOzE8Z5ZC74YKEmSW0rXgNepNC7RQykc
bUpavQ9qPIxfhwzxOdQ5ubhBgZw67yT9GhuK4fvFprrO17/F80pEsUjxpBdg0ksO
5EKXOTshBSlIsZRZPIXcTj10WN9mOOgaCqmP1TBM7KfhhZOCKfO1AOVwtwsfsJo5
q9VEwk53CgmmGJm++voqp0d2dAziSfg32eV8/mQHKMl0wTTxGIpPan8Wt3KHdD6V
MDrYYLY0L4HUX+iz5Qms+VhGobPd1qvsRQ2k5yoB9aJgshrMPcflwXGQFg7EkHAw
mQ7E+HUurHLOGoLsVG8SjwanIc9qv+o8Ppk+BNrmMWcIVS7QILvSK7gf6UypoL8O
O0DjmrcfIDXenc+byP4I8YGWPwNQv2iPF9JO7iSgcNsxvdOi7tmUnW/QOXo6pj22
wQEA3sXbUf7QhjQYKtsaezOKXW9FyZkw+JSGZ4Y8MNkUhDtEDKsKWygH4ppY2p0B
6UKUy4QmD0X2CvwlWX+8rxhAGY6HzWYKW5CtepPMkizUQILk2Ouw+k4pKkBSPJbr
QvH0GZNgfPxO2x2CYLKX2xbPuEfoMpYzHJ/KHxfQ7Iz2+uOCJOJ/R6e36F92uJT9
yV2yjAimDxIC5WXDFvBM6aV1mYzCjs7iuZHIRBp7V88xbiBTPwS1HafpOpgjm6tp
twEEOpIeuXl89OLn2Hz/bPaJIaJZz2ypDSntj12oFVFAAw8RLmLS9wVpnwhaLl3k
1xUKYhzEPQAc7kqBRthMZ4MW1Lrtmf0O2hlQvGwxl1w1cJgqwpOcDvza+rsywpdi
v++o6LRKY4DEnIzqf4/m5KDjzTyPOnhCDZ5aI/RMDIdI+s9/CnJm/LqEp/dFVu+P
Ca9eOHuYdZNpwqlDbchEm4v8uVIZg9x9+7q+Jqxtmrx4tdM0CoAah7DB2OmKZ16d
61bB222Fmz38+KR9yYpuwqPpPtj8j0NgBWNKN3ArCXtbyeTBmsI2ciBZA29ht8yK
cseDtib/4Xwm8vW3h3P2SbBd232ADat/5ETjf/JfUaxDIEGi/ezCMKC9Y0koHs3T
NmWMhO2BuzfqCrJnRCLhD9UCtaawUKQVjKKY7pMz+y88Vob6PsfMhR22YeHXjVkp
69o4X9o6OZwQ52m9rwAQn9sNLBuZCM0Z6ltfDMlX5AzC4xlTS+yiKmzYOxtrJOI7
mkaZnVDDU+GMiPm6f2Hnc6n5ZGbcoVJa5+et65WHMIL2YalFL9uecRwoffTPvnRa
rYbZ2foiLx0JVeI01tSspe0o6yxULip+w1H6PwB68x3I9juDUqEjp30uU1pcwTrh
F07MzT0bDTtqRo6JPSYAgCg4EeDmJjYd/RlE0ulHGQAz8aKX/TFVUw6tQ5dnNsoB
RRsMJatK8eco/7OS7TrPo+Rvmh81SC0OE/nTfq2FnuZBvzYNYHXvx9WkOtPJZo5s
SoxYo7JoangyRB/OIRpwXlKv00v7U/HthGP6qLF7c0kmvjO5kf24EwfK3p4HiECI
tQHI25bWcCnuOVffGs5JGwZAQgitKJZAVCjdxWv/qBSp8Ecowpo7HLV1XvRMqRs9
bPNmhO+xmzHHqxExfB6rhHD21DPdsT3jfCx5IKNJj5XK3q9uWNXQp5hdw95FqzcJ
tvFuX25AXNFpzbYGSN+DYfcrBToDwyRnKBL1kqvdXxtTi0FJJ9Ca8RHd3PH2HoLn
BU9nPHNYoZlmSK4CGcdK31AWSi5fogib3eVftybru5lV0BHeMlzqjHFrRqtfZXsE
5jjvYwV4hYbSHuzB5X0LWmuF8CZeNeL4cawDRYOYkVgaT/5oW1PyIFWhfHHp/lVB
Hg41XJWWVdBXl2tI4AM3KfVYY4CWazPDMc0UGEElnvjVPa/g2FmYBfRDF2cSpTfP
VdBltk9NPRXSF07JIL7CMW8yaDUaEcP5bjTDOZ8ORsdWmrsjIFQZE1++6Mo/Awh0
0YaG+UkfbMh8IOtTviDXa9qlT1rzkFrN7uQNJTxzoTACxbSJYTeMwEoUilA5XYut
1S6cMcWIcntcYj0F1yTSY7FH/GUoHy4CkP9IUsGex2q0MtCBjWU/N3VN/RshUFNy
7KBbTNmhVZ0jOk7FJSU4mmQsFyYg6a+RW6RUWDQ3/gsa3n0ffdiqQHt5X2ajM/tK
nOwvxIRdeObVSrSbRfshDn+HeSNGg+vJSpuIuUK/4UywiBfKcxXREZEImC2TJCTl
O4nf0AP0hLAMNXb+kMdOBpe2ZIcbdowRSkX3xB0dwAdtPryAMVqk6beqVqyuw3tD
kdvYJnN+091Qt6NGk2aWeT3xX+j/oUYy34kzEW/kI7kQuTrHOAdxLWCpyH30/zLf
bvAdoCUUslQ2vt8DaWY0+7zQtXd8Segap6Z3fc7K/qgecRSG4KN7xIDX8csSJybF
EAiUcstaQncY+FIe7yOTXN7N21ySIAziSwGtJ+4FBwektPKTC4O9lLF8FLbFKNVj
smt/R2f4Gl4Rteaz5xnKP0gfnLwh7fttKTFVTgAPHN2U7lyQQ9YAT8Mpfzcni5U5
wSOVI47dv3NlIGXt4W1XmYPdUJN5FhNdB7trpNToHL1sx85d19Z8Ct6pq7FpFGsq
zXhg0GZWP4PPvlym9LIMVaHcrEpAK0AnBDbvf6k+z7YM7cY6dFwlxFiexviE24aC
HbZ5wBtS49UdANF999kocGIWPk2N+TAkmir9KXi/2WOPhKbfTjQ2UrTV5HOYCiRR
NI8gjCle+1Zn/f6zvqmgJx+CEU2Xm5ob9TeyQtIkGKlj0/Zc7LSmhIPSSaEqm1Zq
QjR14HfF+QxMGK8lJPpJP/vNLm95ViWpbIwV644F0DvN4lUUjIqdxS2PkpiIHEMD
4xCvuViSO4LSohshwDrG66iC9w2r4VkhufeiU9pmN+ki4kM5AP87o1rhQFPlephw
PaYKQdKQ8RYYPUGEtjSWrQGQR4h6UkCuT3JHbPKjML+MkMFYuQCiy5uLG/vtXzQD
K3I4Nis07HKb52hSnL4Wwj0I6butF30tgIRAreHXxG2xnPDhs5YaFxjgd//0nc7c
Xwp0mAwvwPPdaWEZ8G0a49XJtiagxMY9BClbWTqNVf2pkOS87d6HRIp4M3A9UhKi
A+EapKFX75kIJQAQMjmKZPFd2YGihGxd5DtII/Yp2HMgiUYs8SRawSfxK3KNyyhE
1CMeVKAqGpTMKTTK/Y9INykRuQ376bnkgnvmG191OtI4YvfAr7JXBX4u50ZqWxAm
7Xln4Sn/8lvw6Gmyuy4tvXDjzr4t0iziubzi27ooyPmNFysvUeBb1S7I2FVAfAwl
5uX29TzoJ93HhXeNWrkcmoz491Jakycy62EXPnPj+UU8GJlt+H7hkmxgXA8ZQ9fT
RKqTimMmIe7p78MVR21/9BLcJ9AvUVcz4XvQjd4PEbsAACLxU496PCtc9KYjGZEB
+dTtpkBUtmUq8pV95vWaAdr5TE5USBCGJPAyPmUlIVMlrWJRxWA2zML+q8CDJ4AK
v6oTz4eXyEKpNgl3MbqmIb5jqJc3ClUeskSeTkbFLajbb/gkXNLKuhemx+8E3SPb
p270VQYENlZZgokMGiQc2ZrMy2zEghHhjfU70pq8pOGfu8J/evA9CxJGjvH/bKPC
hr7OXOxKCo0sdzMfV09Kq5aYK1/iqGeHEd/0+YkjWUtj5BX2DwDazuqTZuI1sWOm
30BzU2y1vYFAkwuf41L2CJvDoQy0tICQ6IBWx//8NYa0vXRNbLddbVpQyrYEJnh+
2dBndkzwzRvm8wX2+PFZoI+d/1NaZhinMf1zvzVj6EI9nEd4+pIvuSChbr9+bTy0
tIigCt2pB92DI6BtEUugwyyNhnTY7jBcdaJRcG7PbcQFYmbxQVMySiWyka6HMfnf
ybx4RdSfhmpapmb5bdJrONBLZi75GALtaZtfnjsIwpvNifXGfEQoj+qc+aRE2MhV
DOE1rf5sjc/y8dPhkSI4ABetnhPir51dfOEBT0yZf3zPRIXQnRSZHngYZRgM5IQP
rtxif+VsFkYWTi4/Kj3DclzS6lIckhwuS3mdWMWWPgnTXqCOBQrVAFdnslEPTbWf
b7uNkQF66Rm50gG9gFU3ORdfw6Ar8o3hZ4g7m2NgwXJAGOPAI0k/W4r9vWN9RZPx
s6+G6KDCDI252hu6mNjXoxwfzA+8M/XueaZoRHzdsHITtDmiacl0HkNQSH+wciti
MVc95brKun0JrS4cYIkPvlrFclsv34vV7Bne6LSorlidyv+A201N50tX6WfbYNiZ
7o/E5vhK9t43qwPyJiQlv+EX2CHhR82MSCP6hNJXu4Gs75UADl1iItUfKmnVKYMS
/C10fHAdIdGGjWBlGRZrQYVOtvMgrP/lj76FJnX8t+DEB58rycqY9LCa18XsXbSX
a3yO7Cy4jQ7/Pf1YJ/4f4zznh39fijTuZU3LPFtNRVt57MUCes7q1C1PYzWXjRRu
j/ha1g2x6Wt04T6qwVQkL1ShrCAWpAyf2vLtb9bMU2QYpc4nabSt/q/yE2ML3D7n
xWZgKoV2VHWw0igDXv1HIucZ0pS49lO7bMJItroSfDRjKca3/kxdw9/hFDaTVV1/
kFBNBinnZQ/dbToNKDE88hHrg0/F7H3cBA4Y/y1S9ID+LS99DRJeCJmLxIFrcIdA
CiSsBkwCgx3qUunmBk642fMc+tOtydOPkFr79HjnKwyeFctf3pmeHWqbjgXMMS7i
mxiQg8WGBV/en6xtqKR7RUYRqRTB850wGr2f3lW1nXK6kgSgp3VHFDCA9gysVJu2
TGtBnGXpfPydqp1eG3hhK8jnNCPfsT1AEU9FANos32XjwqHlJTRQHuN22rgToEH/
3Kj+IzpQak++W02Cmm8LV9Oo3X67ByMJvmN+hEiyQVc8hF4aX6OWrxH2CZRbIBl8
OIfQP8tmFRpuv8ByFAGZFveKntNfRHtHHxPYWN0vMxEnmmLCSsKxdnKt1fq1Miz1
pfqHts1xvZjJVGNzr0ZP8qp9DTCYr+vSiVhYbUjxosyWFd6Q3ufHHic77LTIjvTY
mnCftADvxJbXUNs/0aUe/bx3hrWfpDt8m2OIcTCtHZcK/MjJjUqC36zkvTkiXMgC
Zbo1bJ6koWTh9BwzdOt7rzvB1gAD9RS9bTY7hP1DIazFTYbRSL71rMvuTaqC4Jlf
zaU3GnTCb0Uaond7GcdCltVkRlKR0Xxitdjzb9kYmXiUjuFJ/zZnLV/Z3YBhn249
SU3rJUsYXhE8A5rlAhYpvB3wC69pXNtAd5oDX2I1bQZ4xkr6KbCFAyyianiq4Eec
0SEC4dX7Eyp5kydiTvH+5TaDBRwVJJeO06XHx1QWrQGVUABVxkJ3XSAn5kVkv6t8
s17Wk88sM0xLIGP3f4UnClBXahweadfCbr+aHRnmp5dnD+vpl8iTjPLam8sLsjGJ
iTJP+weVPWk6KnxIZNyfelHJSC+HG5kBx4+eaGKEpU9XsUpuGHHbxMKyj55nLOXZ
vxlhVMcFDNaCfghi1Vz6cYlz6SgU6HzpODE2PSj1FIjcb/sHPZUETDFfZrY6GaOc
0UrgBKbGeINd6rZjLP6P1YJmVsuJFoXoSydNhYHrT/3zUh2jgLL9xDEJ593+888/
MiwogpaYWLnZfDc8sf0ZTl63xbauqsgZdWKvrT4ww/YpThrOL1gC+KH+4BDoRnSW
jmt+talX+Jzxwd+Pq6nOMcqSXImVgmqhjh8f7GmE1j3SoDJZcESocW1HmvLhh3aU
emeWXfOUuE9APAAmS3+bkxoSweg8a3+XE+n6K2ZOF3/Tvqdk6NaB3e4mcXigYORM
pYix8CDlTYCnz67o4fKB0kKfdUhKG5/lFhx8ivon7YKSFLYPSr9xPjR6GgkgTeVc
Fmz+aT0zZpum6tlgu+oGAdfEd21iAqpAt4GMB1iBmVcky93/5zWH6f9G8BgGaLIe
8uRg7zZox/pHthl2RIvVA8ZsdAGOTG4SbG1unmVJ1jECPY+tERoCOlzFbyO9f4LH
dlT4UPI92yqXw5MA5sB46jOrjOy0v9aw/xfH/dP/VT8naQDRH5e2shVs33dK0ver
pn7tOayyEps3EJrUVdeyQpgReCcuuqCMhk53ownjcSZtkFCwgB9kfMDvDHF5Nq4t
80KQmn40tih/dVBvEFKH1QxyOA0KLizi8DHhFejISE3jqdord7Rtcmr4/x+vPFAA
hWrb3WdvOssro3+ZGvPx8KgQcsZrjw35xNIWBvjntSscjbV/RrnLW4nmR+0bd7AC
sMeAmg08ootK81CUB5ZDUg17z7p95RBLrHPBJ07wNNOT4RzE/oM4/MLYAmy6iYg+
xZyvWWRFdR9DhuTrgEXVPj3CtD2fzPd7b9CAxm8fwll0x9mYhho8JdCMEVDpKpbk
fl+SEzrWnaKE0JNFYlrblmLpJ3B9CSaP7HeBd0hjJr4Fu+kgREK3UEjn1h/qdSTF
g+ULUtvxhbSQad76VvKgfBDz+nIfMaKMYXPwhO8PEEaiMEpsqRjebK3qA7Q/nymD
DTBGrRGj4EaG5dcODtYQgI/jpcrNl2DuWhMoFDLj1kMAxaRf+ReS004Z0sk87OtY
52OzNiT5qFL/fXR5lgNI9swczzZkE5GU8ScIBofl9CocDIsQcAIRbWpQLM+8sjwf
6DvNXBz2aJwOC3b1v/kkb1Squlj5+yrvLEhnuFgbb7i4HYC+7Nt+1olNHg/LZ3jt
1hmM8/bWuL9oODe8MePCHaGelun2hqB5NgfCXHojjpwiomHJklcywl8wOHXZjSSh
HnIfnWPSxcjmbCRX9rh8V1XndmOaBvaFTaZlcuvavawaeaTEUuTdkmiEwphR+QzM
smD9hJqN0GkYFixYXAnp0hqx3PV/eGi7BiopiGmQaubu9MhYNUl+KNl2R3aaBycy
b8oOSuuGZvKDyL5yOunISmLzQCowDSVE9qvoerOKtOKFakede4Wu3kSV4FRKYaso
L5gNANYOvsM1Qwr2cZWEbTWoH+nm0sddBd1yev9bSyT9IIjZHrRzl0tnYew2yXDu
ZQd9H+aYgqmTpoWOCdxwo0wfZA8TCFmBHrrmch3MklFic/NtSVOk72PosFxn0AEy
ZqrnCif7u+YJ+wfD3CsphXa22I6L6NJ58l/NuhHNSbf1Wzkoz6kMJJZuvNHWdbsJ
o0HUm8y2MeDDInBLj7D9L5pRR3V9RWvCgMFN9huG6YluGIH+oMrNw8Tus8Z3KNfs
tZtaj/z5bH0V7RJnO5GGlpWc4y+FAhT8blvsYJhu04e8yQIMECw35DIErQ78X0Vk
jueIjD4s/h45nVta4V7tYGOtY8DOCTwtn1NEg2cuA4oukDQ1JkI85+zteMqLVDdO
OeCRd4WHMwWS5yO0z56cqveXgh5heJzVMXpLN78x1CC9WBACBowchkXFojxVVYe1
OqJdS3dw7bO5Cw/W6W7XsieKPaCnKYa4yuxQqxtOu/gK9TKYhhv4RF8JfybJ1+Di
Va8tQslEryVrSX4zn9zxgq/TcAPWD1akxlAAhqX3v4e1VkWnYNbXbVzJaAoUsmyo
bHiWAQTKwiwTUdq393/NciZ0IBpx7VItrHIsAn7Os+ipT3t9K7sPgPU8av6TVHM8
qe9XsWL3+yQY7EgxLfg0rW15Pms/2yA8fx+LsU6NV0+LC5nSsPdUyMShqegWNOPU
JRT9pWQepot7CIc9B6g5eM5qHfN6bwNxE9nl1NWpb6H/wBHozz1N06q6VSdBVwLz
+AO58+AHw57+QFP5laLccX++fNYy2twjuvWVrh4/N9clHBsYWfOPPg+PLuOh0onj
o+a/eldmxAWDZVQIDv9mYl5rubL0WTxsDEwogD4togvV5B1OYet0jMx6FAkG7kbR
EpLtNFHYrJJKrAb/c3U6MEd7h/g0uhCsbKyAhjDkMvLM5oEaAdsS9DAQjPWApZFf
E/Jea+HLFaxZ5gs2MiHZCtUHrzqvHHZSbnhFrJm2FnmSao1cDy1D8ESB0b0FWlxH
BV7Kzt7FavELLchbDLd7UUBxmjEUf0yh5pXOcs2P6q8PO12jw+C1VDtaCURH9+F3
z76Ug8dfjhV0uavqilTf4YvoAHpbhAxhvnDhe+jGWH4ucqtBfiP4ztaAUiPBL/St
qZhNlm4+NDiwJCUwktkQDpHkK2veDqWDQ82Pcw2qdnn0LLy+5ho23DN7MwRUtdGd
ZES0F+iSTAfmmkO2GFqpzgINDT7FFH/nwlqgU1/YFrwti5Z0OMutYMKXMw0OuQ8A
m6Kv9C9hcmEFaY2sKJoO/q/pnEKvWqVQxautgsfAL1/k/28Uq/VQyYt6cImW7jpv
ZWWxVB8mTy7R+KpYOkKy1HwT980PYwqcCQFNnPQta67VA+LCj7DTx4U5XsDvf6xQ
wmUvZWGQSZKCXWVlDhZAhcwykdilb+PLS/NJ9CJelaTQKmuruXhdNVqGNlyyVKIG
bN3qPdTbEg4afoj+8h2mmo2t68aaqk/OUmiT7wqdhzR9jjpfahF/a3NjT9jFXrOU
1nqPOapYgYtfiSfBtY8M8b7jefwF741HDZwBY99doveJb+OPC/PbWqaYAmT0LPj5
PjmK6OUZcPlTISWM0cObKhbDiViWbqpICRLuoklKtwwQnEW4g+tzt5MKYJagZG6D
5eehxIu2TAQFv/dLd0ZdWuBiEk+EMOr7200OKcPaVfBj6u8ux/PHdeBMieMN2CiM
QoqYpwpAtKPJgFBnjNZxWATkNbHIROsCfjwCov0mM+489UyQJWeuqQ34rhoYDunv
takD3JunTgxKH2eiLsUAkDaovEq8uh365WUL268QZ/IDhAUu5Tfd2QOegR9lktSI
0r3uuE5NU3XPncb/LAGqzrMOj4UOoW3qgDJl24Q26/0xRK59oJsg2UBxWnHxmCHW
zHAVVkFfHlGqPsSCwman7VF/gri34IP+6C8GgF2nBN8VR369lvQT0DaaTCu1ua3C
Xg4sAFxWE/43ivfs+Y2H8dtOebRD98QWIB9kHS6PBjGCdgTfdwsD5E04rrqgia2t
YEVE4jG1lwATSRyswlgO4Vxd9Do1+7ilgUxTlPm0jB3OkG3gLkefIJc4EFCwL48r
oH+Csv3U/Dn3KcKBBTKI3DAaaqYZDgw/YpZKMyHkAcTZHxQMcUkGqZw2yiuxgvfL
34gPvNOS+q95T6P1GIl0hMxFeEn5W+klRMXB9AG9qobr+YEpiSKNm/zzMCxgISb3
SSZCUG2c1RNk4LSB8xzlJgc5Gw1O5F1bK65UK5ChHDqcXBEncDGfoszoLYD8b4C7
kl0+S3CY2VFE5qtDa7HMPIBdN0kE8BM01szrDTUHINolyzXpYbuzT+o+9uRqONxX
MmO1UaxjagbBG3n40bshMfjZyR0hq7VvLI7htVQ5/pn5UmTk2ExCrLHb1cAu86vF
GpVrbmUIgc/lPlsOZvyFy5MJYvIQbOJ5BvZuMzQk68mxhh97F27YV3giR6sAOQbH
jLoJNcszqfh/8hzVKJRMQDbqNKQyVJWs0v1Ux0aSHBvnX23LWXAA4QmokjULDwFA
+m3y0hq95hXryOQSHj3hORCPuBVYTFY2mDVDnommG84r2wbR7GrlTVTF9knp7I9X
SxPBZZZFiL2XfOO5zL4EwqqY/Ko1FqEYIUhiyl9gNM/4l4tyCvFts9ZmsmewOB9R
nSGw5nps2CoGaVRCgQcYX1cqZMNxDLZg9gwMfawkrcYxEhksTklAvGhpNPd5RPUS
4OZxU9djdntGGZQhBi1oQ4sLfmQcii1f/nKzBM2X+6wQm6lZR/TPnc+oQAsTBdpI
m2NsA+++wBIXBYrdokIHfHk4vw94ajT3lyR5mdHCDqP7U0TBWv2BVF/+faqcW8qi
GQyd8jTTs/hLCzvcQw4Uo5f7EF2TJ2vKUClK37jexFyWNmWfwXkY+wHivwo44Qjy
aVzPgQafT63vkMWuPbUF/LurcED2fCajTevey5bhEHCwZRUTN8eboBWU0itQEXGB
wuTz7GL8qW9n+v1+A2w63hQ2G/rbrYmoz+lE2s1JRm3J3BghtqJpfd27so/40V9d
+N+hCR6RSmejVlCPTnP1qcwJ/3D0dNrJRK+6fCjR/m3lqECyXd1//Z7ODYaKU+dP
8Mgg945HLn9C15N/8Iqa3qvP/Cpj0SkbDue3iWyvebKjFxuyh/QAlDBvWHQ2NNBr
dQKpKcgnIVx/ei4BlloesPiT4QFcD9bQFaDhAhmNM8VI3mDADxohG/Ifk8NhUcCq
xkIAw4/KrHOPaMYvtnAAlcDJOkC4Zz0xpHEVABsr9QAon/wlfFCCNZM4SqK+TQbD
gkWoINEeMlQZVwIp8XaWauKH90xp35o8FL/Tq1Jps5EtEw7x+Od+c5VvWWOOVMt4
fOf5gQFEEC7HydikE6fDziv2r/ziwOaheMv++ZS/DcHBzZJADycBYgogBzZAw3A4
EAfswVV31uxYCvZ2XiVv32irZCQfpia9Oa2gtMt64mNdpShNVNtbzyk/LkXY4s0I
FHW5hAZso3TwYh+V93NK0tDzNi04U8gmyL9eFvjuEqyFinSCVILTZyp81oUpD1d3
Ix5f55ieY8PfgK2WOPdV55+TzIokE/QgxzY+hJ9O2kcHM2uRxXwBtoxo1hkwG3yK
YrrcdKeO9m8Q+JAgIZtAXkzdlwbB8c3Tjxz7DP1ECEFUotBNFYcdAEkh9VBohDDM
80B3zUcf67/fI9uuwA5gMh5MjhrxJv3ocbTAjdx/MwbqpDjk7EuLYJ01Ai0Lu57Y
nb+VRNVU8M7zEkNewmMB4d+z914VPe9xSDwVR9x9GtB/yyAlMlPWWzYpdMbeN8JR
xYuuqWAaXvOnxcgpja+ekkrqEefZjdGXUCVFAbwTiMcz4spUcWQYLgolw6JaU/3d
FmZHTGTEM4fySd7eOYQLViFp4fUbSJnUuE0Ttn6PKNZYFUVHNgHFCuDhWes+Ew3a
qGhV1jODORDNPx7xnJci4DtpoNvVMlqQRgoBtCTWNeGhqJCnt5j+HnD8i0gypIGq
B8ZB/ckyQ7AoIGU0FjW1dYWIMDsYm49MYXXImKXMyuMoQDUCDE61c1C6buDVWNjk
C2SRsdqJ27Nr5Jf04KM6hk4WWroGa+139fYJaJWFaBJUpQoYWAE9Q4BP39s6hc56
d9+MmEC6nGBn1hKjvZEZWM6zMHqEyA5jH16euXQJxVU+bjh2AqOl3USUPCgZfli2
1fgjcELWoIjA37FtYRKQyXyOw1JtqKHORYL0igSXFxTyha5oRjpNKPdfSG0R1nhh
BndPPCm3PVsdwPugph+mP/zdzHba4WmbDBlRKOKoTmR/L9Ml0nvTPxvSDVfvVFFL
j1CPmFLIIqSgjSCCXlkBI4Ij/yu+U5OU6dynhNgPSqgriRHLLC5HKFRLpz5KrVXT
uqXvmFy5FarzrZUT8zAE59Rv28/23cI5yh+Zb64zz98BEyp3ULcjiueW2GS7n4Bg
d0/Z4pumEOrZCqr0UPZ+q3U4HHINkjsBIELqnD/gbIdhecsKHH4k2QcpbzUVl1rU
XdCmdOPpPIDNRnsWLdOrNzIRVC2fxqD6rHGmHQkE2s8voCFzOx//P1h2cnVvQ4T+
atPwoMBR4PBmKRW0HaL31JZE5JS/AFq9VEQqiKwGJm9YwuP6ozGh6ytPdWnDWLwR
MZ47ossWFZ33N0pPE4F2tk7+ODpgsCfq9WaH7quZ1kFiGCoU8KncZFxnfmLHKIK8
Y4UjhhzkDcaX8cgy9Gw72Hpno5y5lmmiRG1jRRGJQUlEm8LcoQ0Atu8ss0zn5L+D
BXVdWtJQjTayuJirYt5OTgnCRJB9zVf6z/4PsPdn9mT/HVebD22w6ZGu4cDgKzlz
pVsuQULhQrlA4Qb4Mf9lFf7ye3pukfPDRAnMfmQc2qfjERy+9HliPMB+aRymv4hn
JNFd250ORAKmpikNgSTAU+g6Oe89ZYbQYh7gduoyIYFECJPzATfTulRK0rEq52DB
stKneF3DGbc7bE91MmwQ/AtAUcOvYFWimdNimk2B3zf8rpEj+F71oyODRCzzf9PH
JLJIOyN3Eek28cjktzigfv4i6HkJG2RwzcLFby0r1gYy3uT+LxJdD0CEZ/98z8DV
2Bn8TR4KuvnKh+fMKN0bx83Ews9WQGZrY2sY7kFwUMyCGEWLO18DgFWbOZinbgpb
bd4DnaqGrNpmsr5/O+zy1Ovdarbq6R1yAwIYYWXYGXdJer5xS6QQYvWdSRPg2czL
iMZiktlbANLO4qDZkhbaQYaA3+QqBiQbfXSxTXHlBXBgxCddmXzKiRImnNI4BigL
pOq9Z5g5SpF2Ea8NCJ2vw6u1I2ujtLC/hQhBXJguOyjzWY+gQGZuzvaLrFUQDN5s
khzBpvZyJ20BtyuAzZ1Oln6ZURDAgiXDhyJmh7QQEtRoTaQv2U1ldvtkoGd8qIip
dhTf4uUJxSLPAvEUalS16LGuXMxfixIeXICCS/XOasY3vzmaQ3jUJYWfzAo6tfDJ
T2OKPOT9Od4XIainpkDd6CeRr+C1ZqLBiXqdBWo9pn59LvSy8HkCY8Erm72/nPNG
pXwW6mH5IVZgR6PeFVqk5BegNQGbqsxeASHstg0MaQWlDwNgGWGNQmmxmFDaQUKA
tUhsypSdcOjAJ4XzFropq4YO+zld4kq700SKdD0xerf73xjEp0Xofnwr1Yo6lbvA
2y5yRRX2WFN1KGYAH/QhH0Oga4wfI7+QPH/l9mGAmSr/RXfzVxeXFRrqP3+Yd9X+
e5ygFuOTazaEy/VVVFjYxK9dmU5hEO86FdGlAohm96QLCZFqibWcAxR/Bc3kLWTm
5jMH16N5DEAS2YFSSpFgV5/p2phlbajN62GtiAMx7bzAbBdku36GQ70iMoLbOYyw
GpkZn5m1a5IJdeElL3OtZk6xRX/1tzGhYWjQ4i9ZWI+RbVUr1xt8Qz3xfyHw3Thv
31WZrI+vHdX5kHPL++4vbuWbvz8u56I4f6cO2bHMhaDZE/SSU6ymWQIJj9mz8UEO
rqHUwIfsXhGy4XuUPy/XdKcTJSq2cCCdduh/ryzKVbsWDeZ7V2f31dPIQJMVhtv4
m6r1JLaHbgwmmnxMYF/7ZdSuhvmi1rEgpJxSnlY2FNtNWU8QQFRppQj5tAeCz8oe
OWoqdFzvg3QYGyCXmddyPrdVDpbYb7Uj2dK6a0JcxrcObtoU9ATGH+/VOJ+LrqNP
DOXMIknoQQsgmhM+AZjSSUFuDe4CsFwMZu9qg29nGfYPgrmssviunC1jXpo2nmqd
FidRSyp+wsLtbsle0TSZwztldmBzSieXQ1uXpaNHlgXy3GE2hvoYhpHk1HAbPrVI
cFavQewOpjnrY1MdLnfI9gXUqfJuMN6rKy21GeBfDLaCw/UPEISb7b6dPpSUl1YY
0B7UYnq0FWbP51WJyOg+JTT5gEVUpi2rlrruhChC8PezLcYheoz8UGkZJpA+C7cX
XTQzaLs5H5xrf4ywvb9aQNMlfz/m7XrUj0WGgC293ye0c9/ST5APsrFq2kdhEB/x
E4Sp5fGt80zYQEj+SDPYM6BfF1iBE35t1/QkayRx5EgBCLvsKVtJVG/1oelhtw3S
mlHFBTHFu0oYFgGcA/CmnKcwFDd40pmkJQxL5x/1jfXFucjC9JlD775FpuSFZVLC
3p/x6u0ff5dDddAo9AFrHmLSnwFrELREeR8OS0kK8T1dzSlHyXip23U8eZRW5It/
nwgLCmHTMRGzybxz6Mi3lvy1D2uHqjaUbhPhlHhfqX+4yv+IIP8f7VoPEeqahP/f
iEwkgzjojijI9Dw/VaewcJvhK9mm2+tNMQTjrVQId5KhXgFRUJc7SEhrvgCpMm4m
rvW1s3jDjXAFWLNZ7LYUqYXb7oH1iF1UlWCf6sc9kbgEGNfaYhJ0m7xv31LwZEv0
xIoKZQlOTNzrDHbbwe0g+kqAqbyPByQaSmX8DAiH1kDWrFGHHb81ze6XBFKL8VOK
F9h27Rzh1+9qR4snz/Cs86RBa8rFz0qmdvfZl4TpJeIrHYvTrQUGvFqkz5vRSH5e
219XwMnH5/fICmAJtG3ipalG/4BA0Unv0kDRij5ZJVGRX9dKT8ArlcRAFLOav0hF
0PTDI9wk+J8qU/ggKtIih0EULJ3JG2sUpZIOJo9mHdSahR6iLpVzr34if48soH5l
h+wN0mrYKaOv18Q7cU2CJGdRecRUSz6nGolr/gLojFo0QUxT7bkYJ+HaoIxZR7pN
P6bhkPU5IhmhzhJ07B0+LA==
`protect end_protected