`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3952 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhDB3ruPjBpbjY7601ZaNdHSs618xFF3kDHo/c+eTTl/4
vhEAmXo5tmy0l2ak+2z3Y/avO2YDsiz6jSBGXe0865xkfjDwft6EslxCsp8i39qT
mdQzwHoHQTncbszDxdRMGKW3zdnCk0lN/gmkuOwL/4wp9QS/L3vhv3tz+7wQIgl7
HaQOidshJjqrHuBv0TlFMpCP7tQMpt/cFEdyP/L4WJ2PSe4CP9ZyhCNkqE+0Cbgj
Ywiht2XAT8MbOnluJlo2GjTom8JMNlculisLqr0pk0DeaXSg6oxDXR4S+JMMdbsZ
OBPhkIlvt+T34IFRC5cBLihvXIACRySHenuaov6mmZdJwfl+rwCpVzxi2jFwI58r
7icPcwziZezwuCm5neAD5Zr665AHv/QQAJRLtCxJh+jTw2PqoPO8nYJWNcr/7KuQ
PHhU6FyNnQmt/xgD9MxEjpB9P2h3iw0za63MC7teqwqP3E0Dt5YKhzpqN9Hz1mqB
4AnoWMNysaUEIlSIdxKC9W9ge2FdwGItZVTdbp/TMV7IPzGSiKRDAAv6mO5cI90+
Ig1KnSLG2v8mLBLWyBLDjILUlXq/DjhdfBOZo1LSVeBY42oCj1b4Kghc4fMxGwe2
izGd31MOwSHXljL+bUm4QGJv1zJmL3/FLWyvOaldSbKMK2zApxiVqEU/HcmGEn+R
N1CJEfytqi+oPbf7Feaou7n0na6veTe5BWx8ymZyf173Bh91Op/FcF0ln/MbXYZG
9BtW61OXkfo1jcxxCNNq/+9kCG8GM0tmXIH0GP0VWtNHrWUSGOxvQKa6gWjMY/Kp
nZNOd68WAuxvFiOiJ110iOqrT4IkMQkEHRL0VJ7RhFI6YORGGKmBgyJP8S3N7zQL
MMZAIuBj74MDpNmPrbR9Co/nJ4uLuiLIJCVR+ocW2LKK1TiK+nLP6B4axz7Ri1yl
FSD8iR1yB9ZeB6sG8MN2nHpkITpFI0ktG97DLEWOaYaYajStom3KkopYzeAa/uBQ
5GERi0tuRqJCBZQYdgDC0RP8WyXpKYHd5XC4WxqMawH4M1fFjFPXLxh+Yad2yvl/
db9VmvEfsAYo82Mcp4YjqLPz06M0Tfr+hNQgVT4LzsNSl9nF8nXOQsz80/PLE6F+
r2KzDHNv/bcb+pSzHPZHdPDYF/uZqTJrYe/nh/G4MfYQDTfkUidi3vSqpukYXCaI
4FI7DgbX9f+bCn9OmkT2P4jeeg61297iH5SDNEFbvsEW5QTc7wEDmwsvoU4RRXvS
VbHv1yR23y+tENgElynMJLvP8ihq0zP77QiOfhh8YffO1XJxipjUWId46eXEOyAX
paUoV4mhEkCLIMGiLXmWSMFCf8++6mxsmUfade40+/43o2zUV1shPdte9oMY9BAy
bq7dfXyZjzYC1g8e0j/9CuU7jolMsQM7FmDpf8A+hHe8wQ6qE3WIMSxHWLD7Qawx
FsEu1YQh7g46ErMGrv30b4SI2ptOKE2CwW5p4slwpxYxMFLgYfW7qGUbnFjLiwoO
GHGBmm/H7sy8um0J0I7tFwibMW2peSlppQinT3fqWfEurjc8axo6QnL/gDHu2rNf
v5ERPH4cI4Lkpx1QdfppOJhNaBpY5GYAUFrqzbsPpYqjRDt81hRb96CTIy/I+65u
ko6kP7C2Qg/J9Kq7IQ98a/1Rk8bC37IjhEb72pEKSyHQ+hlanzCU5IIP8+PmsUuU
jFMQT9l74zSwDJe49qoNIE+Y5gk9nTrLJF0/o9yrWRTficyFawu87mOJkQmS0VxM
sUxiRPSxxnrEd4wVqvnOHRYyKXCc6eTaZhKhFVL9IF5+YTExsKt5YayfExeQchew
I/jrJUFiVeLSSJPBNljj1Be3d1nMdc4Clj/66SEHHgrWQ/oNjeoGJB/zFRGGmObO
fgGTGvYNFJtWOItD8VcIMG3LlvYEExX92JqZJ9mlTFEMOZRaI+cR+SVYczdkKSFx
c2BH4A+OmsaZWQmaKkjQa7yZ9evr5Wmp4tCD08dP6Fbbr5jWifQxr2l2xonuj7zo
4ajbYYIDLe0pqAE3owxl2G1BMWk/FGvT4K9Xl2MpQbzyz09jUDm+UhRMZAKvpJIV
hJitH0AjYlVMMYRyOqz7pLc1nMApzFWSHvuanN4sR+ARl+T9mFKLJ7SalaMcB+kJ
YQeCLz1tlnOdD2DfVvFOs4VvVoIR8ty6jv7I5+ylXMn/EuTwzHdwrKp6VS0+xrHY
Xz9V3QQ/K8sJ6yGfeyFWD+yZi21IfgBXMeJzI/INRCxgwDtcNkr1qRqgdWagNhx2
7CBAaIkPKBhk37UNueU9q1NQZL8fB0XLCxoe0efohIe009Bg8cj3e4jFI9AGkMNQ
ZSskZB8oD616bjfcN+qpfEffkZEoQdXz6INVpiwhaPPt7rzjUN2tUihqA8RbS55f
4YU2bBsXucT0IbRyMsMmeeiLCUaGSIFFj9mzifayDQr7mYCJvtGmC4UNEtvEg2r+
o4IJxtxOYI2AbGUgPxM899/8fIG3CKfwslDBmBjOT01sTX6s8EAGEGYnsegrWYhQ
bt6pVZvEmV+4ka/ky3R96FJlV885h03G4IKZT/VZSpo1M7g44cMg7ZWYVDPWjMK9
zENmP4xpEWGKNxbCGZQ2OwG1RKNCKHstZP4kLHAlshFGeicCInVfCOpPViOx2JBT
AeeebtJylR+iZZoFDQZnp2J1YTvQlHwQ6KnYoJ38rHKmBx102lVi3Kwg8QECzBk6
+LsHATx1TpLm4H0krspW9RrsqPC+wQMAlD+BeYxFMabDPy1v0lT2vA3LBbukeJXc
9zyra0siz8owQkOojTme6+0UazpRlpMR2k+CVaUDMv6irXbtAdC5ituxmw48np6u
lbHbJEGhPqi+PaKnt738tyclaT1j+/K6JdikXoLhIKilVtAnwQjVB9kKRyX+8nV2
Sw4z4AJ445Ucx6Gr/xh38JXjmYR4ApOk9/7jnaNYjUkOuDUB3ZgqKE4K9/6W7NTc
jkM/jxeebVMI0L3ByTqcOLdt52BGcOgC+GEh715+uoCIMk7jHrkGqfFQpRQflglv
5yJNEdSrHclJ2vK0jDPHjiVjHB/V2mvxar8uwcJ+f+iIq7xL9wkLi6inVvwIZWyl
jxym1Lbnni+UZEE6zBBptcABv301pkV8BkchqrslVDRm9Xg+6WjUaQn/c6Lbql5D
SSmXW7dNxQzNyJY2bcLsTtjlttuKBHm87bI9/2BgZu+gqdIgYdkPjjHbDUdiH9sf
rEdjnHXYDDtFf7it88m9cILPTg6Oh0+qPQK6VA5Cm9TgCg0x2VyPNElHi3OBxt4b
YT7TBeK5IfI67m0Lz6sHmCsfedRadihqfAXVFK7B6Q4FF2F/oBa6TXk+pxHSdx/E
vTcOc+dJb0TLE6A89dQJP4SVf9cH0QnJyfs7Ewi90R09KlM6rvrY2hlSXxmu3yVA
ebIQNbgVXX9Rfagewo4OcHuoD7EpYRrn1HtMQLZDbByZnYImwgjxfscpCuCU3lCZ
x3CFYNf/5iVfbn3bJJ5elzk2kdNEAjujnc+SweZ1oTuB/uXKh1dJfHbMxIzEAzkL
CASOqCEFqEgO9xbSfQRpJJUC4mtpU2yaaHzUqSSeKmZ8P3Sy9NVBGQH3tRd01sRR
Ce0cMBI6+bJk/y3E6inu+zKapYjLCfo87CpP7Q/h+O2yxtp51+Oyw3s4P++W4S+d
EoS9Lybg3kWIQnDSO32qifeeHgU6XG3di7Y0OvBJOT390i4BeWlen52fRnXyfCh1
LSrPPd9ELoIXHG2hJIpzEu1eoKaC9JCdAWrGwkMVZIlWPaKP6rKu/il+Xy/6tgLx
YILNoASXxIKfKrCTkLzzDDso56xW8u+7RpyITofknIsml6u4lQkhWAiGwtRVsN2D
hUFyPzBLaBu4ZZDoKNuUeWi8IOlMXzj3RkVWn1rSdoNXecfljLT5jifX4F42eigJ
7LkvV9G6B25/zO7yNIKFhQI96I1LvyxPb/9NcYkzkAwhLCU/UOp7TWsV/fmcJiAM
YHdd3BiEVsEgrNJ+5hUySYcgn5bwqbrVT6cSh3wUFZBYNR77KZuIQ+2A5fY+Cymy
ugylADHMnWOss3RqfPkTOq2Ix0ZTg/np7rY+Kjs+xeRFgtqFZ6HEqDBvkFSu6aFQ
X4uBM8dnWe9z1LmLnz9ZuT9fW6mimmEdtde474jgfkiK/n4CHzMULg2VFlexx1MF
3Ld/cj/Ytd6GFQXMwBwY6FopUgAFqWub3T0jLBkNduyLkKNOBCXJ4BbNEXS+23gK
2jNtSD4i+LSx9TsBxHe1J7k5bDokQwsVuYSNeIviCcKK4QFnbXgnErYMslcEURlE
ARC0kUfrV8dcF5ewVuW1CowJio8yCZYu7lQoS630scrGDQ/D4RYKn7+EdKtk+e1I
fYZ6VFlZOq7IsDQrH8chPvnjSQ+ubgcILSH+W+rfm6WiJJlwVOgSDh0NCm4fk020
jnzEK9Ggabr8feFu1eDDQOTqMZFe9GSnMcSKBwDgn/8LPcat63JpSxDuInDW2H+t
D+yBt8k1lRLNIjEMfpJKZ2qcgbv3zb0c3MsnO7aQI3Z/Rc3f9OccTxSHgDDzl3rO
xRzpEoOhg4lQwPz2FPJXyBr6ORyeuzea8/vDRe3vKauU4/Ks1T7dwEcRPzxG2IHL
75ROIxMJ/w9W3PCrEGbV0Z4ojxTS+mgAoimmkyjlOB+5e1nB+9TeNyMVEqFJypxW
lNSlEG0H1QV/yo7nl51UBLTmvE9SMtUzWL98D0aJWdqkKIA/ovP5XxsWX4Y9TfDx
b4KSOgNzJh1CCUHS9MH8wsIBFb2irkhKFR+7QOPEtNMyhwcLHvlvF/LeEQwA5yGv
lCQ1dOoZuY5VbKbN/yPWcc5k8rkqtvIvoCsoesQPc/mUrSUBuDNgPc/4AEnJzoKe
kdYy5A2U6PPCmI/Ohf7VjxRvUA15+1Z6V75tYp0D8pCoEPb6DK3XSANNHtSTv3F0
8BAfTayxfeyh3Od+9P4C9OPUX6tU4M0+Cr+aWGcu2uKr2Mi1Xx+UTkGoNIzpoOAz
rY6x0kDzjoORBDjKWkbFrhKFAgwpdry9lnPXRZ6+Kh9Q9wSL4DOP5yxlkN6h9PA+
ZQh408uEp2egTX6JHczjZA==
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3952 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl/FaAgkiOwC2yHsDwDNDyf0r+Ya2F/3+Yw2/2nC6rDIx
XPlbBbGDs7kNhvs1Jpp7LrCidZ17O8/Gqq2v9YmumGcvgsEAHpZ8UlwA58HOgZa6
E5UA0A+WSxmFcIg+xov4b+pu4fA2IBSpQjffPmvbAf5SfvbSNWtJX2G697k6u3aF
Yf/KRg4GHtT7643PQuQTCpHTVPa8hClg7m0h0EhNvWIjhYTqKdkaLsW66WyXUvxg
KJJxtknWOczXrqCTbcbxSMZkkKefVBSn18EeX0k3MdUtIuE65Ihb6SmCCtnCwapU
V+j5UA7lB+61P1tK5J+sxi4OggpmUJxg/9q0JwrgpEuEtIEo0q4dmHO9hTM3fDIa
MtkPtOhiC7cOt+8HQ8J0K/zl5uN/yMcy0Q6noRzN0S0tolcNQjLghuPPon6F/k8u
mm4iS3tmEGqdoPkC2k1thlxYzX8/y/mPvTPFIWHMaViimD6By/itNJdX+mj1Wdh3
PP3u/GWmA0gFw2Lir0IlP0fU52tJbG/17nlOM5f4c5eq+otd8ZvTek8MwND4hZNK
ZaCZGPHTP3eHYWZ67fGpu7oSVW/8TFcrnp+5lG69tRsQraoDIKq8Ezn1385kFDjP
CxJACoEsEgIFmOlEpTTP0PHzMKr1SfUjo5aMGkD0267OBxFrJV5a6bKaR0BhamPP
+AUDbPHTcZqusSikvCxOH8n4Lurw/9wFpDTSQXCikdH0b92yqfAGp0FHZGfYIcWz
NqVPgyV5afsDgeLzm1M/siSPvqSpoE5jm0R7Ulq3Q24/bqZhWrjcM2koiM0HO57t
p2sc3FLVJEfY5tvEcZ3q/7Pi72IkeBGzqq5/EBq+9nuzKwzFnLHoJUU5Qg7a1asK
70wTzBi6RKHsu8FbsY65BoQ8tknM9t912H2N0yHbdUFtriAoA9kQ/N7LCcMI8QPS
SFLU1hcpVd6SbuxDxAYcKSHV50PaaLQv2ggkQXthPdfy0rlpJ0qu9asx6NQZ7YV2
hySr+jxUemirjkPnTUMXqb/BGra7iPYFc2hsWxmNeBfET8Rj4xWo1Zc8mTrGaDFK
p74hUc7H09FrovzT06wVDg0IenCTUsMV6bqLEYJFRbuRGqE2YyORZZKXowbvpBRk
fM7EAMEnRJeQhJE+LYesiArDR8n9cb3jkCJAUlkZobcHnfPqZrQrLYbosQH3p+1B
txpwiZu+6EtPqjhMbp2hBSoaQrliSQvSbdEVSDv3kUCyooCEs4Z/LNtbnHKI69T1
1lHEY0ggA2FBuVmngAC2mXuQUbhkeSWD1tRgA2drpKcSCQb7ivAnYmqHt0Z3MAdT
33hUffka6oVbqoHLuxMy+0ISFX1QA/tg5fGkTo2K4T0uOvb9s8Ux0+cP3xhLXI8T
/9rTAWOCjr1WVMCDwlphziHEVbjPy0aoGXE3pbk5JjZ8nlYaqVe8rhodBEfWdWW4
SLFAP85mzxoYdlYTjpSaM39r2vOD/P1WlZKtfcnOxcpHatrd63gvTi39DYxLpo63
eBGnR11IVuts0fBtPljO8r/pvUqwJnwgMBlVgm98m0mlVgKhsyv8JV78Qwfx7JxJ
FTN/FklDqjzWLIeX2D0ATAatk8SI8mkYWJsuUvULVV3kBz2P6Lv5W16rtjv5d3Sa
N5Fga4f8YE+Wq/zGkRGjQqgjh10UejrqKz8ulYcMXOX7jrHNodSzmPi/q/y8GXzk
HuwtCFFgtYq3taYdINIRDmAt3+oZGgaSO2A90kz3BjcyGP8nWqG0WnutrGP2UOmt
zflIihboKZaaKMkBw7oYZMoRbGgZWJJHGlIqDOHN6j+xy0v6F9fJns4i53hOQ+pq
aKY+mi74//VGjKEF5Bf0Yy9K2oUj9HoIQWdmS6j0IUH6ufOew/0LuEUaQHXZv93A
x824bRnZG+ZEaBEC0W/KDzM0A58Wjm+7RSbuc4Z3r7j1L/oqt09x1bIjB3AMAtOj
K7qIYRl/955ufpoe5T3IotWlN1UAE8AK6b7sr+d2A782x3FslhidTC/ZsIXYyJdU
e4Y2vDb3Len90RqIqoPtgzoTCgjE45KzViOVxFRwSQsgUURDRbaE6zQSzSZbbqEs
2M2jEjOA2PYb2q+NfZHQBDICRncTa6d438+pbYcwukyOMdClXZFnz7TsnplbXbjF
GkV9pM3WT0lLyNHIaGK6TKSvBqHQBAOl2FB2I70CxCq4V5+DTqW125JRSWroMRgi
Ar6tRFEH00ciBGmBcYkZ8l3ftXWDc18QDck4pE+nymlqldAbIJW/wIBKp/8lpbBp
u7+Y17QnnyBciuhadsokJZuMAo8L9gRyYhZXtkKLZlNHAMBqD4SihCfP/SoxH/O+
/fVgV2SP9n1Ka2VEhMW1ynODUJMhGKUTQkgbik4tUM7GaSFM+y6Hjrh6gHwEuOmX
j0EUQulnDorkdEFJhUv64hpFvL7j56n3k4vLw4hQf36KVu+E+XdXQOb0cbJx2Z32
mZ7e9lXt6u9vIRpT0goZ0ro8kOibHhwZrx8pEJbZwDtM6KmvqFV0lz8lsV1DWFEC
mQ/eOdNJVueWNKwqKB1CuxKrbb4bgFFGenzH+IKA/osuWbAyRUDFO1h0XgBA0M4U
zvQp52EySZXIhNRZUEPHhafnjNPLu7iIq7tUy4u7E9q4pFzYD0iCGfe6BwGXaADi
EbjQ4kRHRDE5sy37dO0SLhmnkAB8icblZ72aEDd4ADn1vThD/sUwTQaDqzi8ZyeA
zAKAFeYWwW6az8HUo2rgXI9/A5xzX6YlEpz/Cg7ocApY/kU9uCEOkm+K8y8Fl9zs
qTZ0b404gsFAkZQWjZfmEsfqp2M0x7r3I8SfWcS0MrzGA/4SzjYIvRjQxQZDvgHY
XdaNaeZzWUcLizHvB7KlzyrcL3v6laqqe9qrOakkfmjaO8UykYhWuZRCyowy6UpJ
urpemeJdmmpEm/yD0qb9gj5OYwmrWaagU4JBtsFAMTfWWrlZwMcrfccde2OYmQ1r
irVlLfk1QPFLYB9r7/rqcxvR7gAOBDa+gdDusFXY+14DpV81ieQ43SJuK34kM1Qw
sLrLPiE4GVrp3uEo0mDWpIyqgACfhZ9FCXVtsaWKSlZCI4ftQYZHlEXzb8kLeAnz
DQpStvzczrNMAWq8qwT/E+CLkGOgg9T6+dqkPOVr8Vw4JpUwo7O/5y8VLs1SzXlW
2OPi1PsYFaQWNJof3UKYpqEjdHsHBEdtVLiOdquHY6gFo/6/ZlMb5ZZCvrw8iRYK
3TrAu0EwJ9Wcj5vau+8rrhHz3ROr49c5Mvcrgb6LPf5SbFc1GcYpzMlqySIqKhot
NgA6JPlIXZGSqXwCVGwethd4od/iWD2BTK1nhQWEQ717BagEHJdGf2kFDPadofGS
Lm9KN+Bmuy7jel+v2Jnya5C0cLqPuew9WmKsHrJvsXlzsLoWE8Ufsn0o/cafdBHL
R3jMJLRQ1CozDIfJFj8gVJkSRMEkQgMYEIiV8xKAwpGwDAUWbjcHM4/WnX9rbfuS
l8SJQAXWmtrRK9LdY3aMnjpGjXpYgZ8n3Vip7VKX6L6p/sFCt0SpRZX9jkNO6HnH
5zrJp4G6Gw64dtb8mlu8WneEpsQiEzQPnSbzCUAasSqDtOojOB8yd8O9mnJlS7bf
bP6QnUgiYYnMKz29XoexXfhwCe1LBydF+2TsorSUcl2UgBIStpdJeo61CL7qCVCI
RAn4P85J8zwIaMdjzwRiE3tsjz+M/5jniGtpE9WqH8LGxLC5XxYGdFTfsWVel5m3
oldbdrFPiMWE2LBO0ADfKVZW8T6k0VGghpCfthXqwxxNt/DphfogBFmxzJaKOami
/hN1hJB/uLvvirRxwJfWQkA5iK9cW5H/WVB2VuDWnecXmy+gPyUuTGMs3P0wBMay
EmgFBhiIOVrEst4aPl5gFsnZj+575dAvRRHgP2KMZ7vkWzxpKhrXuQO49rymOkpf
4381A0Q1Rfs1/uH28tRgduwUBIlMMFwFKNDpNHrisaHzkEE9QzBZ7e/7Mar0csHI
9hJp8xBTSaLf7DsN1tMTArmLWZCF73kxiRK4GCQourPTWjQ/BSmOZVoKSzA0DI4X
/19ZY9CA/joEYupmmT2YqdhNg6dWZzpBSuLs0IEiUDdPrcGHGdQcaeKppVfuIgVF
cYOTedRdFBqs9BdTjt/HlPxA2YYHkqqx4rwGjxOwE7itcBUqWOXhqJoeTJdu5wdP
dCQ7jF3AHFqWyrOzX8l98gVmCPDDPujEXt8vJAH4l0rM8kIRLQlQGNiol3OxMTqi
TNOPQDbA78XA8oK66K27oQNc9v5wM2Q0O4LCFTMuaH/qkrDHqliv2Npul2T8GQhn
may7FfE6svutqofOxp8I7G6RevdSuSi34C9u40HDENeFlbfwzVpc+vgvVnIxmbYT
3oVktOD+6LuvGMXVY1MkoJ97pT7pq06d1bRb70IFtadEtgauT/dObzB3ozYUiVWm
BQbVQnSS1wRmVxAaXvH5Ai89CdvYDIEMSFVBy22L4fdn8vnQJQSJQl40OTIe3W7B
lG5BhfaPlWpGLJxt4DsVrCu0vVVjEc5CPu13gL1EO28bczdxUAUf3+dl/7hNCLSO
zWebCtQm3pc4i/5vFWeoqxRqlPmk9o+zr9AxbPT7mAo/XLNCzXjp+/opzPr5akiG
ZeKiFzoLv2ezC9uex1akDhDrUrOeM9yl13mf8nQPI7oopr3qnHAbg15ZVxK7IjI+
7Inphh+vvzVv8vBaPuiN1dGYWP7bNRlMgzbYx4Evt+Nw4wxX+thlxl9joKdZJvsC
R8B4R5noJGDVjZbt61kqvI86fnyGsDuUW5ecayJw7PVyW2DdurVAOB9aTG/KeO0g
0p+MnvYF967Fkdm8NtMYG6HPe+HxdEW18mnbNkWgVmSwI9jLxIJF5X3dksigL55q
O+XM8xPLo3/+cVvugxbsN0Gs4Lr/on/0JjigGqO/PEVMAe23mzo76bXToYK8SSrx
YAPDUqi/iKGNmcBFlcnAbdzt0R5s9Y2v9uUclw605bqMi9UgYnjeK2aXaXJ17LeI
wJUjiEpdRW1kLnuI4Zddl6+1z3L409eV/u1N0i87gU8C4QNhdyfNsCQ/f2zSTfnm
39xhI3jsJ+aV3gqgMVCC/A==
>>>>>>> main
`protect end_protected