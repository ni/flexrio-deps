`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
a4neElH2SodzYSxeJ5dQUieARoD/OX61rJ8OpYFMFM8q6OISKMaxgfDDExlmIsgB
Xh621YVmFDLAfbDxQSSM43cPLah+jYLk4fuog86vR4wbjEWwGOxuUDWP0Y9d9yc3
rgx0un4r1KxmkFGsZiYf7A7HxMcEa9HnqwnhW9kurZpn8M+KEhIxyRV+sG476sFC
RYGYADOrivU3QGv64jgPWdK2ucP6Tw2bDzcCRXR3cEUhduvGBltD6SnunQGgSKID
/HdUHgypdnlwAgA2keuvwILwgXE7PZQZyPynyrIcJjRekLfRa2MfiRnSbjYjhyij
60v6hDxw79Enz4tSYc4ZR4frIP1qxW0LxPSgWyBVlZuB2Gw5RNuN3Kuw+rJjo38o
Y0QQnpPUT1fi9NLesef9Awh25cn12iR2Vyrlst/eiBxTW2Fav7WftulZFEi9BEvv
8vhfHtCm+rTUPU8kjx4XsLZtU8D7vNmCXhAahEizfXV3r3ubcmq84eY6l7QGzjiG
WUxoawyb7o0VG6Jcl1MTGABuKkMRuuak9pIs9txmTkybL0EGDnWbcEWUlH0S+ERI
jCaOw1pM0C//km2zHy1thYosfcOGrHD7qpCSOA/mGo50q/2CcRf9j14QhCdu2hi8
RCRYr4xw7QMNtfq6RnBjrrZWZ8PtDmrA8qw0TP3MXiEeTt5AxmNHxA04TvsTueHG
fYHbSNT+IuuDh/VcvzazXkR15QnugITKVeY7bNI3tmIEO8XQ+ekHfCD42dW5uh8b
ZEptOxGg7pI6HR3dIRdkm1xkqtDTcvhZEuBU0n/EUt9wzzJcbP9/MHSYk86e5WVp
6PCY0YTiWKDhihpNigQ7g1KhH+UgEJRHiXXwmT85dgaLju/GPlwbwe3GwQhteebv
7wEz8Q8W4u3X97r7/KDev5T3A/WkI+mFpopRw/hKv5C1I4PhkqIcvZQeQ7t10um1
C3wFq1iEyKJqGpuvs4Bl2EwauJbxCXeeOUHSZTvTdRWHartHbPTIazRDyreBZI8x
WiuK2GdC0Gl8SfIeUAZJigLJD8VeIXEJPr4g8CuAbbmbRxJG+yI8pKEvCNckh6Gr
fNzrWXFy/9f142XakcdzJqnC/j7XMoKeBeYt6rGvDR4pIFp6lP8ubvsbbYcnzW1S
fRIXNc7dMNxcHrZBLOED5+sT1klr3LvOYds2rUChM1HKEhM49Fd7PRCVbtuNp8Gx
Kk30QAdHXOyYAr+2DGg/eGTIM5LKSsBsiZzTl4UTNPCPSAhTmh/c+H/IrKsbKv4Y
7LzYPAXKnsmVJpa2ASz+3IWvl+dtFQpvymMXhmfKPxC85pKoVcn4VG7yuDLMm/BW
WGWHqramzQQC4F/l+iPheShDHqYtgVfud4/yEVJIrn4uAm5TtZv9HBNnx1EtvByr
EPeG4Om5Rtelh+7CMvcwoyWOjDKz3uBpeRGa/nuPYA9bqH9aVa2x1mRzbcB9EKPE
HHeaylH/hJwXxdhxJmt7QMcJD3oNsTb5/n87sk4skgeb8PQlj8F7GHMd7cCUKrOn
/R7KZBuiljjMsQehUkD5yUdjvisb6/bGwVRwbTDy+rKMwmX+fD92Hp79w8bWvA2S
owv87PBQWc/4Agy8oeDunNK4abVZaXc5D6nefbd6/vFrccsPN11PBBeN1aWza6VN
VP7oGS2mdc8jKo/L6Op0uhKXBca/FuVS2fCeA61WcfdHSylhMKWnKu8gfYcJZ4K3
emqIj5gXj6D1KneTRyaiP/LZopbqf8e0ff3YBKcMpaNmLWO/CKiN8GIMSqySh+nZ
Do87+nU/XMbEAqK45Z17ATDnIT7gEnFwfmSNZbdN7gKRt48B2h4QE27g4V+M2Gz5
ATtS9WsXmqlX4hFKg0SnEOOklahvNkOeDj8arcYPvZz+7tocdFr8cqmVUE7YSn51
6II/fsWquzLxk2gH+9IwfespS6wm2E73Qh8Xn3bNMkYN1cmcfKc8Y7o1Rja4e9ej
JjOqL0X/A8JzuwqAwGz+/Ro0O4x5FyoLAMLF48e6Iyf2aSJiH7WWg1OqOsgdVRI4
c85kqWvaDHmrdEWuzySW6Wnbb0Sl0/m3/rHkW76U1xgN/Ko9d61H352Jo/2EU27i
QJ9Sy9qnbo0bnssYSt3sjLpSu1+ssUk8o3YqODiwfwQyAYLFUkxZc4CoKC9CJRk3
upPiETijV4CmL5l/HBZP1LZkeqg8/kmzv/W9DTtoTx6ZfdlJDT9kT3hGodhvIL3n
xf5U0hJrwwtKGhr1R98lKU5V/dajo02fH6WFkWX4EbxGJyUcNi0SH8yEvU0khYDq
ixC8qKSLGXNFO6W6oezZdKCMdGX6zZSGYJkUHZ8KqOePUtPB/5i5z8zqAGbEF+kl
8aI9FC0EZspmKS7okJ8Ydg12k7BWYgt26IDfMl57CXrcrgwaAL9rj3AHHMIKyDrR
X8S3lgzv3PylLE+AQaTqC+h8YqHlhciQHLs8Dt2By+N4D/NU4s8RhlPTE/Nq8WzD
+g2KaaRcKSpkVf/HYKghMhtWA7i1YlDREjWJFuTSkrd7DUXDrWi2NS4tT57DAl52
`protect end_protected