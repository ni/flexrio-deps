`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5744 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
DBGZtUPdvgnvgIFp6VMrQTYaaEDbI8KTaIT0EwA16xWzOYNh4DejC+KZDnUzBa12
Y/Gb1HFbO1EHiO4GOookoiYrS+wCC/mc4mtaIK+sIPLiFoCrCtLOGHKcvFHeZ9dn
qT3U8L6b6DYnFt0OVUc0karyxcvtP/w+GpASv7KQ6pN5La3kxRjnI84qUbUcRhHT
v/JV+srn6/KImpIkPlRz9eCgfzjXaDzU4/FbtGumg9MlU1dUHOZ9EgsZnnzMfpgH
LnjC+nHJEnt8nZylpQgaJfRXWEeBvUL0n23ark1WTWNpfnVQ1bL+QOzNPpRZDSxr
CWftp6VpX2S3/cqsYhihSQEnOpzDk7k7G9SoL3RHW5qnTSzG5StGWOZMQFQ535uw
TKIaNWYgMbJAwR5CZFUupAC4QDuJpg3r0OqLZgf0HKMYo9SrScY223SF31ssSONo
BQPMasxsVcn0UsA1l/DA9pBLG4RWfMIcrWbWT3brauJbTJmL3WTRuKEABlEFxRa2
WApyiYgCTEzHSJC8W9W1wKEzjEz6q9epQqKCIOkUSAGR6jamaUocyL1Gj0f46f01
qWDo0T4ndZsv6/pjDNMOS50a85uYanhj0211x3+5U+NqG0wxsdrX6bWQblL/Qb8g
WO5xx5o58U12fbd508nCWantAKOfBUwtqPbC0UfwKW1bN9jsVyfWiK/sCAyMeg94
ZVMPb32Lk69yNXTZ64pnSItAfUJ8q1SVHE/StSLhwm4LSm4ZpqeYY0H+KiVfohPA
hYcayval/71yYMLQu5ByI3Y4G9MZLDVT/KIs5AO0NldmFAN4SHrTiW0EfbM9ccTs
l/4nWofPnn06OHBnMrLsIYX+MxFCMUJC+SZ1rWSYcVHgf5z384k8oSPo9xN4uV8i
GQdDS8LN9zWNWh1sGwMPgt97YW1bHuYKO5DoBI10zxbx0mBTuPKJPr290rdWatwE
xfM/6rGg3sJkw54L62LXs/SnfaT4gy9F5fK7m8eUNLB7YDO0KWPFTAevpgGSplTs
3EfjJhW9Gjz18KmcOUGcS91+kw/6nO4GD1eAGBN0QLZzVgSsrmrdJ2JLzyA2R9P1
MTjA6yOuRwWdqaqQcDRp39Pdfw3O2vHhSkQ+BLbrJiYfIGZ16OrC4LOK26P07nhz
GDyuaJmSfCijlQpO53rqgCqq62RC+BM9cXAAM4uI4BRNHr8s/R6IMqyKwD4v9A5n
Wq3NovRhERVii6EzxTiElJ+JVSmuxCxAOS8qgMs9RStou8TgYJADbqn1XDzMj6GH
lpfasdWZ5Mqwv50EaWK5OOjrpk9LYtqXJ6pyBePp8oabhvJHZXQshiBCo4l3SzuM
v7LxwPQRer45mKq6oOqjjFnN3ISll/DOK5WOG+JxX3wxvrvvOzx+kI9Ht1H0E1DE
it67Mg+GurdutJTRh+0b+YK2p88pVw0E5euBjc3ufsD+bPIaXk3bSy6PkW+vcadN
7W/oM9VFdIBKoCrPZXMLt5o3FPAs2v2+RWFuHqGEU1AhAAMh82tKWiOV5o2o+UcL
0KQerSdhis54N4oaPe/4zlhj0usO9DCBusTpc1OhKwlOIc1YPr+gSMwD7EJwVbPv
bXEU46IP2ILanHP4LSKRO+ktzN6ZAXUNtge1KHv0phRP+eO8OrkVPhFGDkfglJpf
leTzafI+l/rdZG32C/e7dgL1B4Ji2WaxMJfdkraJtucJ2oX6aZA5qa9KbXArCJir
Jh4QYABy62JI3Spj65LVKnO16w4jfsFbIS4bRshWsEdsQ+QK4gwKN+qF+HORfrY5
gx8Z7CgiBQpvRA7L/v5xXgK1XTTzl7bMpNlVw3Gnd9klPptWVrQNXzW5fFl1cGA8
phufjYzZpQBpw0utuDinYtWDlOuqW0VJk+GJyD8nyuVmX+447wpfh8mLfKKuz9Bt
ESBKnFjqqSvECK34GUN30gQ/pEHpku6U7bei63bvjUDqJU/VcKJGhnB7BuNQej+v
bKLqZwWBpQXV6Duj+r8cwFizzRwJsxQLISwEUZs8ww0qKJfYA7Jp1dtU0twxNFwI
ZzlhXC/qIeKA7FUU4o6CAoghN3E6z29bJqQAcSC6ztag5mfjA/OdzMlA2sOLsRTz
8UHIyquDW5STXeWcJSMflvuy3TZLyVzIL0U8p3UKH+vaoCR+nn+LdFenyjyqytye
EE5NnL/rrgS2fv+Kp5vqXWP8/mn/h2TSbXBXHDMtd1Pa33ccaf+leiV1cqMOYuHB
hUP/18yjTIANb/BPg+SDnDIHHnu5wkAJd5OUERbqBvnxFdlorDJgeTMUtOaD7n3q
yeizlgxpu0amaH+d9Ihxv+iZn9ePhyOgQI5zWctgzT8BJpwG/KZ+8jGGI1kPgeCU
ZlyqCQx1UtJPzGUcQ7FM6cpPp9klFbEOrUJUoQHXFt4FdvpuoV1Wyk169e9q94x8
RoKtM1vO+tkYhycnhOWTsE6wVNf0i9YgDti3XNMkKm/FZdpCgUsj3Y+TSXFDnbga
edlKZsGzgQe0tXAms1UeRwMZDKDgkNZ5cDLFExRjemAtrD/tOXmtaF1YIsAVl9V6
E4rGR0gQjB3jV3URUUnIonaR8WITQW0P2Pca1US7lky4OB6zPIQId5kc1ASvm1ZX
9DcV0PaC2reydmsejzQzWchDAmuKyPqTDbafF96sQK5bMgeJYvmJrpLukBi7FDLd
avD9YG3EA5MEOCDi0WUlVM3zOVB8kGTznYNxiR4CCUsmKBOY2jVGxMB1LdYBu2lg
DEehTX0j8zWYYD94ouk5E+RW5brhjBYJURiBYCgC9cLrQhJCjx8x2fqlpYjyJ5wI
8/F9ciHCNNKLIL/sx332kjDZX6AnDGLOfEogZtP5XH+AUEiLU0xVmI0rLNZYMCZg
brrM72XnEypJ/KdNVGGCaY04opNgcDYYa9rX9x82TbUqBikkMWFB2Kn3hsurHPMn
kl+p8ZEmNOC4vmlux90YlEAJu5+E9H7C76XTTRtSpKG+7w6lrhYr/CYcLqgNKhQY
yMxLDzPGscCBK/m/aMjHewir2xdPIrZdQ4H5Oa4FyLZ7PVzieGQMLrxbiJbrV/3K
8G84megfbnhsSQDQmb1C0g3wGCbHRH0YA2pTIaV0iUE4FY9MFaPgzkS/UB/j0nC5
fRFr2c16amb5LtdqOjAgp/wJC5/HtigzxSixT5CUW4ZcyxS/uhQL2OEw46EhUarb
kqoOzR8CJvJzeUpXThpOjj6F9NO5l5lqoaLfScKdtwLmdsbDzsV6poPpJ0L9kuOR
i9MVk/m+OyJO/DktgoOhr/jraXQo2JslFz7tRqPdrEU6e/+k7qsdR7jMhRMwO+/5
qDP9tRK4fiS4kFypIk+bDDYhyNak+ughLzag9jzZN+f85nF8YIkUTyXm9TeGw15a
sTnOu+IVH4tBMV6sf+jIYlJcNv+8ofa2iUSbOfFpZhRvKtNFlG9rZlFhs0SlyC+P
1pXf9BstvY0msBeOcFFaaCo7qrNAnx1OGu9SjBl3HfaxK76z4WQ2mg876ubub1HS
Ye0VWIn1ej+4Qz+D52Gj67omm4qacMni4O7sxA+o+waNeYyop2YbPwqSe98bDCQN
rpEmqF2FguUSZhcYUbDwiSxUPrQcxtRcZ0nlVquClGK6FUDWFoZSg5asEFz3BNFX
SeRzX04beIg/xZgo1oBEqUMWZfW067HwhzK0LG3BhFpK6f+SAOVXskFUK+FA7s92
MwKzpPB7K0+ZukVJ7U7V1/m+ZrxW95TBB3Zu8lKtldg3XVsIlSeGzFV+8ap7K1pk
amGW7tlw7CEYuaGV+F6bLj1jilsP/jwI9Ln0H0m6xdnH75hOvmEV4vR+iQmEh7A7
R89kah38EJ6c9q0w1OLo9OVnZthUAcoyID3FMUHAOwT6AGuE4y5P5P7kuYMHFIsg
SukEL1VyvjvoM5JpjqzzIj6VPU4QO2OY81nTRiS/v4FAKQfN+B8vX9DSsQ+yMPoo
yuM/WzRZ2Ei+NPIc/ki0jjs0jASoMvn7pdrdJKt2nE/Fi77USoDgazcaSV7c0AB5
xPfOPA7hcomxGIp4qMmUkgOZZ1Ax4QpUln8fnQVGt1y5Ua8vQdTfuuAqJ9rsFXvq
URT6CDyd/00MuZIDScLV5sQkqbu9sBdn6ZOsEE7g1Ed4m4xwnoyBXmw7gieFsvic
xKnLsKRhm7T1VaaIU+cVW08wvn9gpxUlrtJ47wGg+hNkbFWhnQO8y+TbIJ2hD0hN
cdi/XOCgaLqkFXn3vHT7GOtEtS/9Feqx66m9KIJlLeB82BXFejhWiw1iXzjfztXh
BqiyGwUwi4W2ddgZdGUwXzZGVxSs0qAws6ipQ4U9VOmDGHO3wEAAiXElzZ7iGBJ4
qaqigXQ9kz6sNVUEefheBxhVBpm+H1EHoBRCC1k2X0uv+Ov1vLTiA/PLSIahHeuw
Iuxk1UMKoFoY+pdelMUvu1+YnSF07Tjir7GTVHyfko8kOv9rh9o5YyKR+bfrDQOi
O5Gymu7DdRWJKxtAzzxbGxxijPE8Nvxo5eYO7mX2Q6qM4992V7yKvoRMeroSLTvy
rdrMFwd+ImZvYjI1Es9utQsvb+xjFMROUsDCeEUxKzGmKYPp0+HCJn5z3cGKGQlA
/RAtARAPylIqZx26b6b/mGXoQQiBNC1dzTZGtw5a0tHtZQGUctsoL+vjipL3/m3w
xlzgBzLZRFSZeiKvLQitzaSnQ3mRCWTi5plIehsKnuVmxepoZpVyU3ctkyJyShkX
qmNP+BQRr5a6F12ivZgSHbaBj8+B7AVyHZ9aMxEAYbqXnsgSdtjdVp27eitmuE+D
qrDUW7LdXMR7Rt9dJVo4UCn1ra0r6FE/6AQKG5V/H0lH877xnsSxm7BPMAQ6gpOi
SKksvKbbn+wjdNWgLYV0wRSJNaFqtQXlFbLgSUZCCaDiS3TzM5i63IYJFte1KfzB
QW6hEO8aEwsFrjkSNj8m7ThXeqmpO/JV1zNtCrcKa/g/BcIn6VKRBBVpkRvyI8Kz
WMsepG2JHKpsoPIAjIgVPHdETwVsNkkgns+6w/9gD9rOgmk0bTofxvUbjRcAPlEY
TRfGQBsQZGZQ29eBV5khya3EDRcYwIrkH7ZfslYwUXq1RRPiVIjUZNyl3JbdxJ29
01nPkjUjQkdEJGRlIDUMQz0Pw3t33y+4OHQaQJ2YCsJ8TixR+2xG6YHdYpZ8JQ1+
Vwt3BUJgjN1yU3aAhJupicFBXSwDfP3hrF0y3T4587Jkkcpy1yNjzau9DyewbkgN
NPdJ5xqhgxHFQ5ikKS2mnqo9Lv5WquyUwyz+mu9AV8CDaBUVOqqShDQkyYJZx/4t
M5JeTMPrn1tKHVrmvwTusAAWsN3xzV33dkdWjcpS2W50Cf8wuZ+QNKQX87p+Q9wB
x30eO3DcUEhU035yZBIcmgpkJgopK9qJ3env5WPhKDFVrj1/Rg4H5Za1TjFL/yo9
/FnZMgObJOwdDg6iLw30J9a/9awbXvxhsT9nhnzVvbn4GYJLimaKeEQaeZ6TDj0w
k+zsf3V+9NTpadNS15ZoOGJesbNhiNkz71x13N96YCZTko2M9f2R9U5DhwXnUem2
URPV1KkEsH6UXfA6TbF+oAboNlgL/kWntOv3mdX32S3eXPNKKvHsBa+fe/546lc1
kAeUCTDo5PYkWzXvM7D4DETeq7BUO9zG66wXpGsH6eX5cdNvQixxLVFEMzmszfkD
PWB4E7pTqFQwrfb9xtA0k/DTAJqbLyJxYLrKV/n3bYtLUKfrj00txQ2UtGY22aCZ
SE3x2Wxda1GCJnCwbnycm3sD0pgQYhiIlUztov/x1uEGUlnAqz5ZeiLy1TQFdNMP
vdIst0GkE0oRb9yjEDyQDA4XSsGExhSeXlQRDTWWAko7kzLQPkfu9rbr0OjLYnXQ
jet3dfCP7iVI484B5tX2wdCyf+wXpN0gFg8HZ0gHv+fh7Uj2TD2/LXoPSHBakAdb
xr9smzMdC56oqVhFs+UzZKNw5kAtIDGUCUeKZlPgozvbI7PnBLl1kET8A28LTRk/
HXzUJaH1dOEH3EsWxiBcUMTnTZNoQBKO6+J6vKXt3LM7DO+AseO2sTpvOMgzSq7B
qKh1v4wROf8thBaEy5/OLv5vt/Fw0yUge9Cq+rDTGDuhoyVRlIv0bJGYfZnONLhQ
PP2Pj35seijhXTF+qKL8puWHWeUrORlMhF+6T56rk+qFcUYz2HzWRJ3B8uHBzK8f
v3ZfQwO7QhKIdZKCbDXdQC52uZAr/Sbw3ytUuboM+A+ovwAVtYis8e0JthXQGNKF
XBiz0cCk5gRIBZD+PAJPafCvCTsCKqqSqGemk3/8L1GrCkoLvDp/gkuKNZT0YKsu
ywmT3ZeKTmbTRngvsJUwvoYvZhnMmzrB8FFgohfYxe9JngXymhD2jIihA4fX0bUT
R9WU1dkrEKpctTWEVgvY0mXz9DerRSXI3WwJDw8uqn2nifU9gKR/X1SK/dqinz0/
bMYVw9xK0173olbnyJQpCKKQ9ASmyGKQgodUIBiAEXlEA8LreU9JHjAOLk6sJOe2
ahJRL3EIiBs94YZp2SepOYfYZs85HF59Sj4ApRb+fbqs2LgDmWpkpuc2LaV16Zhx
r2vbBZ9hTVfo/YhJYPZch7jyxxjYfi/5e8Q3du6pr8XGf1XV3WHjCot3BD5TzQwn
MmF6cpj0xOa00kxUd+I4th9yczUAl7mGzvULC6nYBfOHyxiB9HnQHXfmuInbTPy9
vRxvS1punRT32aIXDLGqGeI4x4GLNYHAx9VtdgiProQMNUD2rZlMAQONh3dGPCyU
y05f3qmP+OQZDRRIPV8lAGCL6tvO96vagEVwUYH8ZG2xa3mO9cYwjQI6fowX+i38
XCF3/CzJVAv9/rU9CsFN+84qHpjKIU4SRU5DGL1313XWp4q/SZXmlNCLGw5cyZZ7
4VRfhki7GLdcAYGsKFrpe01IuHK0t0P3Nst/dQqIzKbovMMwzyTY5no5pZ1MW43P
qtmHUAsB5kdczRM4WwS7VQVIxKPbuJwsixjuaU5VwdTMwO4JErIo7/64Swik7fAr
KfbjgDcArYKk8nTQdWScjnWm69ibG4+kqtmoOMfCSKWrV6RytiUY6Vzukq2Pu+lh
Glv2iNhD4HYnEOeTgIhUV+Lv1Q1KNOcHs5BI7LPzTODu2NrAVLBUq2uvd+AZtFiu
MfZj+mP6Iu37Kj1reuFgIIVEWSaMbtSaZkgLXXgyDZLMyyB696NJtIIOEj9IMZg4
DrkGdb3KzriWSgqU8QKVBPwvqJfFubI6Zq+Hdfu3pmro0uoKcToDajY22bh8JDrg
F76PxGDlk/2r0YegvbNZVAk2sbYMec+KsbwY8hJyMsDCEg/Jz2GhtV88/kEEjYDu
f00tJYIkNyq4ngnURAPM3gBXgCQnT/WlWhdzfFwGLXn/dWoj6qYgXSdoNIsYU+Xk
jRBWzhug4EQgiEcm9OuF4NdLm6DX9xmdkOG7z/mKP98TJxDtXAY4jIGstoDcLETZ
tBuD5xWFb9CcYAMlj4/xylMVOFFhX9M78MD6p2eq4mg=
`protect end_protected