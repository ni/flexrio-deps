`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Jm2uGAVYfY7w9Y5qKstopObZuZAEY3b/Io3MSEcWLhjjnKulVhCBBYAEQrAzzGsT
vMbffkdZgjdXQUg8jOLJXSHZ0Dgbnob2vlppjZs3bgyHCF7MoJ35E+LOsaLimUA7
hlqStcK49hR1hdeBPr/OwfT3UeVrRtQyq0eJXQ1UksinX1G9Pz3/CmcGfTZ/C72x
p9icpt0bkY4/1I4GBvNCsA6FFKH947JqH27OPACiQQRW/K7JToQn+1uhWr3LA1od
lbVrWu8PdZi7zW9gK3jiW5GaPjwbYQGqeGFs3bTKBILjb7sYHxfxw7eDLVMAIu5D
W+OTIN4JiHiE1gCnNEvkSQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="pm+c2fYA/4JT1uhlJGVUubML8hZi8lME4xPobg/m8uM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
nBaXksR//iZ9fraC7WMJWWSrjqRXHxmM1Y0+KKN3b10NElDzVNMlR76DLrcnamFd
2n7uzsxWqhhJR5LBl98SXO3Y90J6BMbw+OBG/MFM/zUulxh2Si5YK5G9GCrG9gvZ
5JomxuZFDu9CzlWGTuRUt6FsE4Lr6sOL1P+hraQDpMk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="M8TXDiNa0BVMX1P60yIvW2WA9jKGGy8GtbuPknDnC9I="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
/5TNZvs8Nu0G+mfp7M8H+iVAGG3Mh5DYZ0Gn3rRNhV8b5CcJKgjQajrRoGl/gSxp
rBAhtT8Vd5eelHgtvBjpvFBA/EBUrRH6CG6pqRt9r2qUDt4UernbZbxC3BC14KYF
4VK7XUges/yZxT12vZRIRVVUYa0D/Anv1IFrBGyIk59Gcd4HQ+79R7gMrw+mKVc+
xaGF7TgoHIoi+eXMnFcbV2kTZNz8lDpoPB+tqaMAiTw89lQbDA35Rf4TatF4JVyB
coUAbkge+4TEukWELWei3IuK96LLcsLJHrO60V9ZFqscBTKY1MDtXwLPAuRiGxAq
BzpPX4/ErD1nvBbX0aM17VZ8QX4xYoBlDd+9+p/NzjpP+lUIhUvQq3t2CqTB7N9R
nllPAN07hstfdefz371Td+yEm0dz5xOoYaYx2hdyQYH1CfdrETUOUdOG+n6LbEU/
CVOrkoXxf8pBM0qOGO6UgrI0bJD7op/qVANz4lqEJlQ+L1wFVj05cNhkGKnPFgbm
iqS4Sjp2IR6dVmBK8yAtJb0HlebPJuVlSTUola3k83DH7hrCZ7ywkhBgq5vb+QkZ
nuLTVWLjbR7y8PpXrc6HSoIZMUTfGqirrATY78ywyCEX2WtPkSkVvijX7wOiCsSS
4VBE7jIu+mrHwhy9S1nPmcpWmy584zz/b85t8q+Ei8czhjVwAxh8y0FJuNQYi3vK
6ZxtH+jXNWZUDrOXClwnSRbgePPufQn74VueoObJjXaVzG5A07OBGWyWq2xm4I4B
E8R8OFTYj1bIEL2AzGNKitjhuW1YthengZPEQNXWm2pLsAMaRb0uCF3WKSxFdG40
B7tE+OFz24yextOIdp4WmhJ5yjjCXmWISdnAl1ulZD7kPiEguiJyqjdflIwN+Dv9
pfIAS3Jlh4EmlEfoKbBE0zj5vu+IbvQaqXKrbo0OjV3RbEdhc9k6x8s+yGPm7AZW
ooPNX0ZcJlMXhP1Xz9appFDdYEZ55eu/aZIZFEUAc+wL5gh9f4zbSXFJ9k27LcrT
d4Ou4/G/2nDyuKVEzUn2qDXjosNLKmMH6q2O6lCwquKF0G2AoBcJm/rF7PWBJqYZ
lISA+e9QswCzHcWi4SjmZ1JlS/bQIrLPEAtZIakaXKEIXb61uUAGm7zrfEnRZJ36
J+Ybcisn0lcXh+TERYG9vN6rznTPheDnfUo0tlCbMf8OyHvf12ESDpteHYbvsmBa
AfHnZtHPe1PwqmOhttYeJyZeiCbrllhN3MfL8PGtgAAlE/qqcfmA0vQqaApSGdAv
+Ex4gZLAtHLXDhX0pOX1oon1mQpeY5cbTNsFXjLVpjl7G+REiRtFuHVnQnQMbiQ3
zFv/0JlOFJKuwnLcsYGRTl+98PwjXXc9+o0QfAGkKjur/NxNujbhJHQSCFblpkCO
EDHqXxIMse2Dh9F9uauodgIZOm83zbpixqxj/G5AWkhK/17HxWIQIbqPSCqM5Rpw
Od+TtF1q28SvEWQdMEIMM/II+rknVgVWTUvz1UHpmce60FW0x6DJAHfAXJfeNp2I
9Tm59u1YKfiTolnsOY32gNr8f+Ij2k0yrB7f/oBgZkWzWs+rgsUTOaSXWramLL7J
onLjZgbpqVrYbyvFz9LSraQz+Uw/+PqsvfEtzFUOh71MItr910H19x5mtVngLR0z
ETLyKSYOWjh8OpigaERxm5w4GEXNnoUxXxovlIukCV2u1u3aDK3uxzqCuzTZ9lNF
e7iVcfsLSh6eoXQX3HAkRA+40lwYZLdw3wzGrr/3lfNNwajGbv4g8nNMFvgm6Les
vMfm9eduPLgHfPHoKS6K+GanBVwNN8Iq+6vBngT+UNAxBo9kyPgruv//akmpPqC9
4DymXhmAm+4RA3MBsgyfyKzthV2N1DM2pis0putMrzrO7n4V2+YpEPA3yikETGIG
SKVIjqvKdyCeMkC1MEcgFfRN75BZkva5tQLr06vFLhvwhXfC0npzOyT1ay7PDqB/
23YWvN4d2jZisryeKeyEqrPj6If0jwXoTosPGDz0XuRi3STgt/07DWxR4Kwogg5g
fvVOpLgaBbLlPW569CR5ClLyVkbglLmUZ4OA+b2ypYjltxPNTezd0a5tFpusYaq9
WF0SMG53l4UR+Cd+hVEM/tGw8SB8/rfEWvhmQ3SIb13dcuQ5jQK02xNysd9HinvW
y6VdDcasJFk88HZpSk0oYPorSRrXhQguNl+7mlSfCndp+tQGQ8llAyNnFYuH+TQp
HgN/0qIWggjlP6TDciAEU7+ADb4ik5rsa1Kn7DKqHms=
`protect end_protected