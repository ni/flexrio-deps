`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1744 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
ki93Foj5FzFLQL1TyB6Fq4btZII2OlXNzt2uZXnpl60L4stEuz4um3m9ECeW5Ia0
n05EKn0i496OKhv+iVmynIgA+ElCGlO8obSUjYP1p3jCrFELKfJhndwWOHUzaBs5
oOQWGfQaiZLau9QGu1nR8gj201Uh1YbaB3TSfu8mC9PbZATdWbk1YW08aucHJfoj
+mOedgA4idUzQt5PgiuhitnWIvAST2fVxPz4xAobMmBIsqHOQ/myUI2wje7Mj/7f
mQaJNB4F7SED/A+3uB5pov+L13abh8OWvd9dUp/RdxSBGvHvkgkR29y9fJk3Nf/7
VZm8WRFAac6ts0aDhjFFp2TwLH08S9dRNyhu+OfCQKfP4msttdxl/uridizJs+oQ
lyXE5swwrFPJRK4efBeoAS3Fp5CaUNUF1NHDCS6BtqqwttLY1zyuXh1ZXrGop1oX
srV1EjI4tUg5GMqanq/Id+GuX2ARwED/1/25GnrYNw997YBP+fkvDPnTdMtMxhm+
oLgWmfpfCmR1Gx8VK+YnDkqEIJEds1C3iGjinTtOHTA71LqiBaw02Q3ePkQYcs29
/zvwWJIhGS4rMx0iZx1+Xmf2ZPnsuLeB+3Ddu20LvgmGopdF71iyHz+cHSuOKHbq
J9ht92sbQ/qwFJcvCpX/8P8YrADYu0t+AUiv0ux2DBdIGemB9xlHW78/LpDm1UVf
R4F8SV/lGsv6F0iwbWAJGpE9rZibRLEeW07oZ+Z7dCrkoD4Wug3LAC3+tI09hOkq
N229YUZaMMBuiezLqxNemtScjYPvpShwS+aJW1xwz7+9zyqf6gtOJWBpSbh2ZE+2
4byEY+WZcUUqdBDaAXVqtuV4I2YvTEUeMm1A95fGZKatENSdm9dwTTohRn1itTMJ
f3f9e3q4iIOVoiXXaFKpUs2ybL51Iy2S4ksFAHMHOU4xtXwz0SHWSz/PfbWt783l
jnfNnfUo1VOkA6hg0zfoe+11CkgeGGacRi3o0VVUPfY5+Q2rc71DNmfBeKgwdeZp
rW6VE3LERSnfmEnrv6xvlQIyIkS5q5rLdfH3W3sn5aemUyG8T++W9jRz+Bbn49dT
Wq/gA42RtosR0lDhS6F7Z/RuIR1BnkmOTeeEWxG4EEpqDahcS/avqbhuN3L8hWZZ
ov5gc2CaFxnwwUef21z2a9pllW09Y77kn0QuVD+yjrl6SZ2jQU27539VmPYFecti
WUF2yAM8BvCIJvrVrLvLbB8QQApfz2grDYJlyRZaIBpZ1JbHWzLxf/5e54aojD9n
PT8PtjUKTlButE1Lm5DLJCzoV9r5VRRrgeJBTrT/TauUVdhgs+YTxLP8AITLcJTD
VE4R0GQ1HMrjBobi+RxRztnx+qvOrhORK9PBPMbXyl0meSkn/uYuRS4F3XLwJ9x8
uvRD/5UA+qi3Tjn8vZjny8U7VihB9eJyXOPHa403bifPT0HgHkdCHHST7/Xd3ekw
v+cIXGQJCF24oyd6eE/sHP8/e77GYa4fUbi/eatrxUvuHUY9HKxaPYMgoRGNPDGn
XoCUISPzzaV0h162IxDKZfK/CsL+T1pUnLxrlJadnWXxznyUu0kfw9aF7Ulto22U
Kj0KTdFzSv8wFTsVHQ8nWRXE338RkG4zxEdJTggb7+COYD3u5Dh920KhxpIsy44s
wZHyqEaujUS+GHoVZBVjtDPa9Iv+ubpCAdoWAiZyJSIcP5oLBXTLE6yAzYE9Ob4V
3RipNRU6IysfO5J6CZxLAiu+DGwv5yjpoGukutpqT+Xn/SjQ3fg185MMLL3/2UIN
04e6KHpCQOnzpWGhE8tr3QcAV8xQKDrMpi0PyMADt7Dk1j2kgaE+R30Ab0f/iPqx
LwKUL5A5CvA2o51XsrxJMKNugP3OLt7t4niDGREQ4qkdx/lkGzt6tVjvhwTHwmrc
J7e/8csqIdXH6cmHjquhCvbsE7qgYhYtpDg5RrSkTxxfTbc4uy58xsJnKgIgUd7L
qJC7FMfUbCjN92c9+4g/7cZSVN9USU/JTtVa62x3YCUdTJYRl9SS2AnDisCB3FAE
GnpCUPTjSQsjXC3wxdcc3JbgN1V+/0HMMfP/F0XXldimdy8AHzsU5Yl2o99Q6ynJ
SMmCTJsRf/IorWmetXlmxAe4uQD8n9fMx6SKVX4upNVzC/KQ+2EAeFVIdHVExMtn
AXAoDUS9FNiSAO4OaVMTZA==
`protect end_protected