`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15696 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
QVoh6/ZMejDNAJddTaZkN43b/0p314vzIUwVMFuDfSyDq9D5wSvlNAfw5fBgnd1d
xwiyVoLMtAzEAwvhT48OYb5ZdAGf+J6f56XvH95Z5jpd+IEqMwSrWe4p3UTpwuN5
2rwavKJH/1kozuhrcNzBSDbS/4EKFGdpdEsgFj+B9DfZHn3Ew/UJFDH+BAAzDZqf
8nG2CCktrM0E6PCygMKQDhzlOaFtGkDehrZS3UbYnsNZboXPvJmv8TWfKCLGPxAG
j2cvY8GYz13QYuksveU5wJv7DTQqx0ufVwttE6fD59T8iOpVyn4+13d7GjS+roY9
MOk8YS2j7N23ImFIaHujpat3IT3wLs3SLMiT5xeSe/Py01MN2DGKP6ebB02dWr0L
6OMk5oWHupNJVCLATKBvbBHAfOcA0ZVgJH0h1cWUG/hIFv+J4APDKT8yOoKmRUOj
J8mBznBwPQ1Ha53idMa5eRfbR/hUqVdyLNuTxRPZvtg8QKuG9O9KAYq0uwCcWKc1
yY+ngklt6rJPQCxmBQFtMjCycX7kb3IxG97gFnomTMsl5mhck2sGWAZMjIQIJF/f
NFf68dLGsOXyR3clcEyWuyn68Hg/Bv1OHqojyfgdfrc3lKPuqcA41B2hf2eQWJkI
SK0RzG4ZD1ll7+ZDie5fimRa6IeA+Bc8XO/Xa/5F2Fts6XTr7R7jBUftG5FVJ0h/
mqIyyzEs704ukCp4cSQIc+ZbbF8xkznox5smjvBM05048HNT2m1FPQJRVIOY+fUI
QGaxYdRUl6qTaqbvlQMZiCzrrbnomiwzKV0oTu4DtMM0O3VeHIWaoPIQCIkTy/R2
icEMA/r7m9uiQ0h29nvRHxQZ5jfy3LqLZqc4RWRXb8d2s63IxIehvg2HJCLW0GbW
pCsGMXU1JW/Cc29CSrPjII/B1VkPHWg6oAppiPDqIjvZDdceOW9CdTbJIG/3eAyK
d0DAQyHM3QdLJ2AwA9A13h1kkvrT8OIJ/UdSJvPrx1NOA74cndeP2RmveBfCAV+g
LDzXt9fJL4qTovgFCO4YhE0Y2Tixktxx7xAo9vTKbemgr8WRacXtlTGVFdeXRgVs
eZEoF7TX4X3djyVoTX6fC8YNw7goPU4+yx0URN7t2KlN6fEwscfPyQLntNJj1kXa
AwJ7gU1dZrPE3SrCIvOj+TsPqAeRN9/Ky/zl6iC1VtssXDtP7hTs2dNljd7mVgp/
MAXM9XXZS8HxBiWQnDWNibivvNj5GknOO3e0gSwr9m1cdN844W+9304fupIVBnRI
s0pIuhqX+r4Sz2GOSaV1XQ8FFXOl+ygusn9KYFWP/lMI8XMRfTROeL3pgkI5TVqs
LSPFeL2H/QuF61xzdSH+Fkp4g/gpHJqYy/ZObwr6JXHD5sEMTtEjTayLiDSqacb/
D061fO+N2zLNL3IUT43lIkDZSs4M01PnrVlfMrNgD73jEYa3LU88w/W3HT6/IXDR
I5inDOyFnm5rJt8yCKqGa82Z3latJiRg7+1uficQQZwnlvQomNtWeUFEQbMhSKyx
zroGDM8kbfWaLCEvsrRRLyAyjrDb7vOTJV3VVoOMGECsAcXOiaqHnJv0z4UvnwS4
g5Twn0cv3tzEtbqmpl1zlEN7bPOyOwqBd18doFwkKPeReFawDJs4ojvnSlooZcRy
AKidSgKsz7DTqI9R+OAad9JpfV4HHmv6bqn25wl65r9vqU57QXMexHvb6ltXjkZX
zkxfytnB++WO85qq0DD3L/8o8s4wpObW1CSh/mc6MxI8DZfziVxiBPoQdz7EWKGq
5AK4i8e1cUxC4hcu9SDhS/z3W/w/1W6rC/cuoAJToWVWE4K6OWSqw89apcUgV/7p
toe7hvV8PjfJOMFtsdd5F/g4eUYmW8f7b2+23uiraGHUSYQ0vfJxNQUsZycK7tcI
Oprr4VSCruyqSWE2N17zK7wnRjMeMt3c+s4LVqmZXhL4YCcOXWiF+Dg+q5OC5kdP
T7mX9YqKCHBGcFE5MaRZq73iFqNN1W1d7hO8ZS1y/185yTOQlm2IwOfDKA0+Tq8W
Zq8W0I2pvZRbgqBLU6jeTuM7r26gzrQn78BUOZOPa/vTwqdDWf2nX2Z78aD8kBd6
WQxCX7mwisedwpt3nHM9uwVv8L/6vq84xc8YC8cDkQvr4QH9RNseZppEjQdsgztM
y+g6f78YYwZ+OqTp0KB1tfKG+L4OPCj/D4P4hoOuKeMKdkdG7kMjwTjmfOfznNSg
zwcVfU3XOOswOq6c+h2b5DsHskRUv1HM/MZZjHGbcpZ6lmspTZNI3V93IMx9H2eF
RctpgkrX9y1x26x2GZrRrRQuc0eSRY9jMoSbe7Eda9ktsAVGfibggoSZmME8U0/n
haJfNx93gYuYHC6l5WlIO8DmRN90dBuLvCCm/j5S74AkOwb9zBQsQ6g1OMobKY1H
0XzdD8lJsXhe0Sf+Kakt9e5ve8IeAND9l6pwMbBY5vbO90XeXdgu2UwuUXAfqmlZ
LsySrz4eVOJHNr7m/bCHBzHFHi/aD9FUD/YCO+XuOkxAGVS0oCxtLq191fnVcT/K
kcuedchpvgtPTKccMUdSzhKWCGPvKUo8UYJfhw0eEOfcrKrlKEJsVSStlTtkbZmL
35lNH5oV45WLIaBxfJStG6JIaX0TBEsIel7oiwyVi7AmOEKMx4IMXs/WLZ1dHzd0
VxtwXcC/tsZFxgAQV43zPz+U19Xq9QtAixf2BGm8hO5idcB59LfyWCQWvtvupq3R
ce4SmtSRznywJkHoXJ5Pw3Zz0aH+DzrgJLQ6oCTkZeFShjhBywC6dBBpUuH/2f3i
S60BNn18jLEwX7UG26kPGcpqNCpVqx5fQlJQPBx1Vj3ZfoJotRFWIT1sZ8PZA05w
7ToJjmMmhdqkzj4xOY9DSottdCcAbVVcQZSygpEi4KZ3DZcBJHQtlyH1F1fu5QXk
GTkOHS6xdLGY1LT4R/eLGuMfEVrfehL34SvZOF211R3cEvC/2E0JQqhkzXhxee6w
rDmcQcfNPcbpsmkv5ict9LTCX5ZbZkNfpPhL3nO8NnGTadFiZ4d98s4pjtNdO+Uc
JclFqoGI3LDZuz5uFkkX0lv2H7Ifx94SJyAzknjMFf36OTBYgro3Im6DuZi/5UNk
Ct6k74cOgf26VPnJ+3RYEju+ekbunnp1UuPbeFtolQluIgfey/dc1pnNt/gDhb+r
xJAyLHG/dhKz67SwyrZqgpb4ljizCAwSMnIS707tQhhxbkpcBu4UwuT5M9zQ0iMu
zEr9nBHfaBgmuWpWrmgvnzOLSV5rBWqkfMqpfeenLCGSDzup0soamgEVzFhTngx7
l1o6Nqgv23BxjC76Pxe9iegiGJkPNJNU1mRVtmS5ESjyHwZxcpa8ken3L+Fcf9Ht
+dMI29RcXSnhdc5UZxwMXkQlx9eIqjKXAYcHydxEwSm/jliEKhjP0DoUYHrOGUJz
MmHh8kwWgxDzq56CWCQRIgL/8QvclIcfiylooB++qIf9GEnRNehj/gQQEo1o6IJw
lPcWdpAJTFYQtwineJUb9K+pnyc16JNike5f/c5nyWfRPqoe3u0kzo1hlJtgohcp
hoAmhChfUgvtGlrsvonojOITjiEq52L5QBfr1osmVUw+5J+/KkHZICKh8JN4ktPc
wVwKMxqGcHn9ebECkW6HGsyN97Z1PBksL4wPrbGgaPf7BVCzs9tlOZM1jwuc3Fhm
JLXKnzGF3RLtM6y9y2SpcoqnWRG/URLpgt2P1EVy9JWzD8om0hV8UhVJ4fCE+8u/
aRUJlrKzbUziZ+mWhHgkSenCu98uOKOb+DbfT4bp7ky9vD0zquUkVnndVa7ldIgi
CgVZ5wPJq+R2cZBrGJlZxQ3PYY2Aw2Z9wiHo1/ZufqkX0DjL+oWcrXdOhE5yYYaA
xBc4UETDI0X26n5E95me/WSnq5/LKvm6OHW3GrgUgolmOsbo3yw8wZKUHeQIWzEW
OaYTSabllJwAg1rSXTSZZvoJl2wu5U51Eyzvo9TapIWQlRG/b2xo2PtkxbQdwSHZ
8ER+httYYHahFh58mmLEuw8APGDN4ojPOLChwJBCbEd/trO1r0yFIXwvAlkgZVbm
6sK5B/oPN3t+LzrKf9Fpqb0BY4afRI5cwUo/OsN00vTjV1XPatSmHs+wtChg+yTT
YWhW9H+xWAAhqQCDrMdE6Ac1XeQREYj1i/LgrFZD5VGig4pSLotJA6T9pAh4LrG4
wSeFyL4UlN0zdpeHAp2XLWSuwA1JOoAxfzyxEc1cwin9ljk6RCtGOWnf4FGtdFAm
XGxuwvXuttfRTGaQhE98XP8FHcVCEF6Nq6DiZeWG9Ho84//pCv/8wSvoVQ76fPJ1
tOWku6erfZLBVtd7GTFCEn6tmxKWi8N1EWtm4KoLMAbStWGfkSEzUQReHZauwKnF
4ml0TCVB5GraD4b6dMG/PX4oqz42HhKGO1+daEpU5fco4LiP6iFTqr8NbHY7IZZE
7kspDuhRlu42wJa3ct8FK53LGUvjGj/pBc5S1VR9Z4u518rAhY+soV5ybe5gdyLu
byQNCr3WStMT2TvTUI3INhepiiJkg+wUmc6w0Ul7c4dGY/h13dB2k8K/Q+XG6K83
Yvp6sAW77oMvCsLH7+HKClCMpTgXTetXkvdbOAsM/8ENL3j/MMn3Vx/RkNYFf9/g
ylHLoNsaJXrAw8TjMeiA+7eIdwb8X2WHFmh1bcN/2HmlFIaescfM7law+3wWL8If
ZjCSHSYdcgqwjna251MneGY0OupCh2N9RnVpLNmiDqyNq4RFscsqaiYGBccYyEtT
ySCB4VDBYQ9GzaY89H7QghqsUj7ATUFJoVh8LhPvhMV9MqSsOChREiYhxil7+W3Z
jVOndCtoXib7l52v2XytUOn6BSR709exszjFkZdvD8CSIX1JfceHKMbWXPAqAt5+
HJJFH8IUgVKNiWWKyQqFJRKN5N/mp/ujU9EsWfCIu+LPBTZHx9OPsRhZbre7Ndfl
B7bwHgtJ+ImyqOUWxji3n6yZB4zecgCykhOoPjuNLx/9i6E6q9AC8IhwhK//lkAj
eyG+boOvlGec8FChAANuP+WpEDbhsbRxXwzYJxhOy0n3M5T4Fmtn/g4g+6xPOKVU
UWTXkkG2B23x6GxiMJxHXEbvvFIrj6NNYOPTYGJIpgP7oYiLNkCKMrJp/dwPd0nl
kf+UzP4FB0n5Wp/Rhxdt3oHrKn1p0R01OOoj0uPeVVfrddy5Rbf+aW0jPkxpAsCb
GrpPkOB4j+7ulJMb8Zf8gFxCOzt+5SQinDynBEWZ6NX8IRdJJCVzz3oUqaE6sWxo
3Xx0v0pUq493pWSA9ioKDMinAmHkiZbVuY/oN7KWCcej25wXAP1epzDgw8nqubAL
Z9W1xqqAuToSR/YuuHZwkD6DBODw2V6Gxw+e5ElopbudZpKfwHHJMM3UE1ev5QnW
Vq49Irc53OAPVtPQLkWZqxCGcEjMJpeS5pmKj677oXfroyVKUKCiQKPWFXxuYMSu
QdOyP/edF/waYEKXHaUK3kz51zjd8s19in5c02OA9yn6hOIkuUChvR1rW11SYz6F
USx119rWWWi3lTnnGjw4KJaQ7uiWub4lwfnuFmYQSYr9n1NUWY42Bn1tQxTCKhkW
V/3kbvvdweHsbVUhjqM1H5tXo3Y9fXWYpoX9AQkA+trZIrWZ5V6IasAEgFgJEww4
ms4WHzn6H0ic9QrLl98gUMaQAYAsHYZHf9ZaGUBb6zMcxP6wn54WsF9cUlFMAgJX
nACxcgkg8uUwNuKz8BeU4cCAiylNig5NjRImPh1gIKafIjXA+KMoSOIFPz2LNv7J
8g0PoPu+I4yF2WRM10yTQTYusKxhV+Rio2iGA7n2/CUzxBgkVcIIVnTazmwhkctQ
POAxJEdL2Zw/MkZDtq1l6aZOfpySUAzYzCEEJF9Sevu+DA85248Y7WIi6oDzCGvj
cldPNWtMSHZDC0Qjy/l/aAtFVoCmXcqyoviRpqJx8tWstzplFuIiCywueJ4y4+ap
d8AsINMsR2hTD+3ak4laoq/imFLYNzIyYvi3m1fnqeJ5z8YRvhHQ6RDWbmNNZPiW
K8x5FgmiisZlJesEt3gdyozSfg2uN+NC8fOL41vr4NlroP/yiC8e1vrt6X6gUnuK
pcd9eQx3R516MzuOKW9uOIYcamboUOQ9OmIe4c7r4k11tTuorYz2ddY51p3gxtcB
uCZPRCSmWaAbMO5JQtVp4PGyWkwzm7V/hte5GdpVUxZ15sxiIIxvt2G4NnSloShB
YVDPkoR7XENVblwaohek5wkSFUmmL0srHY12+FH9Nsq8nVeu2NtHUaZor/5Qjv6K
qiJ3KgihlJWFP+P/1+xSQVE/mdNu8+HoAzGqcCgQV8iphHS9a3zQOoqjftUIpZlR
ZtRRd4YFoPgpKgXTihVyegWP7/b7oDBAHpiGfogZOv4nt4/fcTpP1n8fPiXqCNmc
HmHGCr6nBXDTqtcNGtI6GoCQFWCy8bNNf8dCRkI8B2G+WunaBIA4pe6NFtj5V/R1
PjQU25TECnAe7iM1GU4XG/5Z0UEUvzUFXMgtFWJt2hsMVzL2Pu+wLeYhsdVIRqjF
JLKI/6L24KhJGItpwDYmJB9mHlwOt2EdfDdXx9Ztt87NkuFKApBc2yQkdAPEQxQe
wruG27wS0vsvRq7kUOJHiAaFhPvIOBabTuHXtloxmFmE0Japg1mRi5xW8M60ClPV
y1XocCJ+WmLf9huRolaPFo3yEOC4Bztk3v9FoW85UGP0dMSu77tkyxmiiUIQPtjo
pB68s2F3edFdFh9572rdghNjSZctXEMQhGpBJPEZhXAum5a/5PTKe3NnTOFkh1Yb
jK3N+MS85aJPcnnG4xBTt88gge1lz2QpU806u/Vht8cBjeAe7tUK5GMlpdSomHD8
m9aj+xvy0nqzwLhtNMU8N5QF72SM11zBqhlFZEoYusYiMDBEtFxMGNAal7FJM11o
Wq3Lwu0xWIxWXKaFVSwTMbWRMuTNZmeNIU16OySoyxlICeH1Q3c7nUXUa9EuN8UB
Ef51BnqhjOSK+KCN2/tsoGpIhQz5e6HyFljYzfTfxEo5iHVPAsRUIjHLcxN7I5nI
FuMFMtg4RuAWBnmJsotvvuv72tQC2DHSweclyDvgGtjwZzzviutnhowrVVHJ3b50
r4C8w6Nkvk2tJetlaZyGykT3dAWKIx+G3YR7R91Uer0eBz4WogItLNy51dlEzHVX
h4KBXhljrO1+ooYZIZBeiai2dcxywJMm77+3jeyQ50oYZSPBMkmGlSAGdBAWtgKE
H7UzLWzAlx3eNsSP/6c7ru1PryGGfqwPk9N40r84Ipz2DHzpuaj5Fqk2LxLXPmuD
A149XCx1xoBiHocm2BB5RIrHcukkvTwQcqgSN4/JGsHfHuxFHlKCtBWInyONQe+n
qp5I69Ei6u5yHURdXUCtKEbxWwfEgHcJ03Hp2c4zUxZ24rbcDpL47vWuhSPQiCuh
LzjeipLdm1ikSMSRxAYMgt9MKuljkQoqS1Is+FqlOSegxqL8jWD0LekuFCTdBf7Y
S8NOpQ0hJdr56gbJ7kPlEpiYFEEnFdDuTl/l842BIoEfP3l0kz67vYhOyBQIxGcN
hdzfwnw6WuNugKGwMbL2Uh3+I2Hnl9fWVAYzymBp818j/wtgYbXCSyhUm55J4yEU
nEtV8AVuXsZXhrIKDm6nYCPd1Hp+R8JVWBHow4LQqkGM3unLG7ghc+5dHzrZmy9D
9d7Tt+uKDbZ+yf7dDVXy5s8cAph2h+kcAbBvS9ylmPmDq/zXdgN1CYcIUpIQvZIb
vLIguu6ZFt1rkRGfwd4FIHLcfvWlp7ZCrbaM0DD+7MzF5Uv734IEuPuet0zK7gBX
iCAA64MqoKtEc0jE1s0fXpDbv3xq+DBFV/B3GZ+i4Uy6kUqOOT1rtLB0QxcUV+Rt
YCJJzO9XIv7cGXapvmh7B59ezNZwQdTTzeBObjgCGxaMeGoEO+ZoYkHsQpOQ+UGP
jxmuTTylqJNXfOCPZzbTWMr45fTmsZTq3wOI2xa2cJQNJOwSK8BCY/Yzhs88kHTZ
60MR5Te6snYC7kmL4Q/JQbSUsvf9v+FQFEC13rXbbA4DsFscZ1NnGFJQlZrMgzxm
kj2F8lAWYckTr+JFnYmresq/iRp6laAahOyZLtngOrmxsQcNkc6VjYQIJ1OZTdef
O/Zg4WXkM+2BQpCpFu5bFOSfXMI5NPzMTmofwIYxi8EBBXe43J5p9TyuxDOMUgWJ
KA6oiO1RymBxJy0bWtUaLrUzqOSNk6VgJGDee+zRRGXmaKxxVZZLGGyBCs7wGLTO
fJFuNVRk8zI6yWdg7dUKqM44YA8S66gVb9Hixx15nrJdhrxv5C7ZVwSESpDLFGpV
jLCudaBSb29UXJYF3HUTY0lCxIv2wAH2o8g4gvpSWCScEX3nNsKx0469Phq1x/2P
yyh/5Q8CQm0eAq2L5QggYX7mXcDWXBRt9W+I/oE6mrOtnBvGBmXdyFV+hrBv8T2r
ODiCp7ywMkc0hPFwewzsybyRVW0WCPeZN3rHYBBmq5ZH62a2cdNRIomBjnSSHIzr
ukRNLMX820rfOpJWGSj4ZSAYGeWVLHkJq2i6kDhmpXtMptb00TpMalXRIq+rNUbM
fqf0ye3WuI90Qv1LQVeyh5DQUR85pCLv++pdsWAy6ABGS+yjGMVgE0F/iAqrJXF1
nFloDlpsl5ZNKMDwQekuJBWvNWFaRilxGn+l9EapEmS9Qa5bEVYCWv/6Pcx1w4bV
1WZb9lxsDUxorsonA5nEfuErXthfpfYTYvR5QUjKybV8mbYj3FiCxLloL87tx0Yt
76m4Za7agLrd2TffefugxFd2nHB6EkxRGtYx+w92NuFydnt1rNIWkz2TQg2wZSja
QKmv3WRxajOhwE9Wx6Q2jlLVDC3O24RfgaroNHFl+EXwjgTof+wF56ssZKY4ZYCa
yRaAI/CGtnUYZSWjC6xcGS4fSadUqvVZeE7XFm6x6e/SJggsBDPmHFtz2KVojqBR
xTjEv5e/4uP+plhwLqdToGF5ayL7DDlh9pVHJvUDgNGLej/xh8iq8DV/SJCOo2Fo
6OJ5YpNz6++aP9k0389o42dnwHawgGMDCLwFbcsfpFXyB6pkermXhWzjlyxhDw58
/pYX5aOFkQmrcdAFZ05G4hRTmSz3pCrXAIXaj0SkaBe0INufBUzZzJa6SL/RN1vR
prTB2LniIhhpN6xmkBuvR37Ao8OD1oT8emY55bc6Qxl0AXOwMV9u1WBrpRwTRslV
kht5e045c7HzKn5zW1ot5px1iCJlGC7N5324wUTFxvUgOp08DVwZN1zwE+uwH+VJ
/GrZnM1ncFSTMRzVMACM3SPzLTh0ZxeLB3OuBflN3RNIvRXZ1SJGgEqZeHDGbO7H
EQPccV6Q9Vr3F3qkXcgkrPgkK/2p7pnA62sgjvmmiWxvHeqiuFIgUQh2OGm2r+5Z
nDTjcURbgneNZMi6ejB7Q4NHDC/bjSFUaQhSl6Ku7Kkz8Bp2Gw/yEhGKnbLyPVAW
TIRe66TLufDvuZsk6DxCvjJWAmOlYPhxpMFVy22OXZZqWqH7gsLs7eIA8Btk0Njr
N1B8curZKLke8jIRlNaYdHfNGKd+TUaSPQbILgmEftJe4JmrXSrGbFJsEA2+3tc6
Z0IXa16y0sHiGxQLmChz1b1On6s+e3fltKm6JF5OT2u9Jw1loQROfZ3Ia+qCc6xf
LTuWcZgnl6xtfWZp7Ttalq/qF7d3FGdGBT6+4pRmzTPVRXDVkJLBfdTPkDzE4Nsw
imym4WJmngZXiIwvQZ/0AWallXKaCW/u2hIvZWOg8zdEKTzu19iP0Q0pgEr9jOJ2
E7/v5iLhIx4QMm9CtjiZeccsyNjs1RnJ6oR+jkYbW49Nthuy1N1Al1DkVtasq1Sp
riDyus0TwqacsWffFz8umiJe6zez1AmoHR3nUs8VWPk+YaMmpdKo4huQj2E9pbWq
oj41PkI1pR16kQcxtq8ncSjEu7m603oAGapMDGtdML61334BipvHCYxrN/KABceN
QdUaqukq+RXgR5b471zgHkr9jDFN/IV0iPAIhqeBPJD4OYy7pUvKvLitSU1PnKjV
6Vq1M5PIvJH68FOMKnSl4FhkIoI1psWxLiavY6eiDeITzqFFZdTFwgIooFJrO/yP
yGxXvShH9RQSzQQI1A7DtNsvQHvLBiS8lcGqCgHji+aq/OBr5sK1Azmk8LVkGZ+z
nS89PcKfti0SeWGOj/504YgGiTSprH5k8/FzUdk2wCNh4IphAXD1fRiUqtXWoc5A
Pj9KTv0Kx+G+bWoWl0hcPR2FNCA3JH41IxHbSx/Tr6bTxIbJiBHN4JVfWwCWjf8i
3nO+zoMX53OOyn0gdBpvO2kRNqd9xB7Pegtgq0wZD6on7Lb3w0CkK+hMBCaEDQzT
wBVVB6/6szYnp0saQl1xD0rhuANiDWLG4PgpnGRlyXey7Lzno4wfMOhFO4DWSYtN
hYmMssRrzHife7bxk6xsawBvqrlSuY36fpkDLO9/+rtJjxm3PtF9cgNkTKuv6Ce/
HUjuIPpid3NFWpfLXc2TKu+3oeakuf4GpnMHcKxtjJtF3Q0sJmRaW52f/YtzVpUS
p4I3wz0uCS5TFt18iefgpaJYbo29Y4MMbuIHLsglecR6QV7FAN3FSP9E2iBbkUgs
AaCW6BevGrYsnxTH5fAuJeW3/wCHWZmMCDAeMOyRm28bcuLVflVVaXRzxpA0782Y
aqWPWnmc4QDMJdIBs3n+qzkaWVwsI1d6R2c1jCvvHzcud1j8oUqGsFa7xu9wcVxy
GzNqD5a8jTP1C0QAD3g4WvE/OlMFMELOCZ6lfrL+xHA2ze0yRnPg58oViQCa86KR
dMi5skZ2CVolJdg/oEewDIfe5Ne2ovO/RA1C0xYVNl1AfATQegY9xjKfaaZPZ4MU
6Gf10qm4odElUL+uEPOgbz7CuMxY2afCCUiSy8TesUHXsePyPsCYEE3zOg+69uVg
v98dWzFP7/VbjD2wvcn3a0Rbka/7lYHa0w4cnXPkf19zzrRaFIlRPs0b4djIuNKt
ycUpSuj1ztYP+ihBKCeK2wStH98YK6OldECsdi2FqMCIoRs8caiYR5kj0gGw/QKH
qZqr/9q5FJ837az/+NgjTvewTcSqUXiE2L/BfsWhVn1B/8KakSitvlOaTeEZ5JMF
H2/gMVQ10m6kWdMiyJrw4C+EfPr/rhCTMM6rRA1PF6qYEPkilT5fU02GqrkJZhIU
0zTs3cmiqQBIQDoUGYmHU7W+d0/V3DdoBX3h8O1yJl0s7Uqti9PVbNFSUo10jyaO
iZC9ciQyfT1CEaiaSPtIM27B9z6qeMnSEcJ04Ujmgu22uT19Sex9vb00ymfdHFjd
k1boBK04RBpp0mRqj0c6GIWY4xiLC00IKvmRHdApnvYUQavBmG9B8cGZ/G2sZCxp
YV+2jjj3QWPzxZ6vX9nIwmjrekOIcZ+52osjU6YWNhsITwmp05fZzh0wa908aeiR
9lqGYQT6IzweXRiA95ziTXa05fRnnYKSwhEbO10PBGjrOflvbFo5KvNmUmIYNK7u
+NaNc4j/L34vNPxoxxea083YHDoCe1tli2a8Ye/RXV20iLPTbhZz9j1I6Q/2S0WQ
OoRboGoGqToFXNj1L8opvxaYdbXZmSmtLFT9P6uDlcY5A/ffWx6a12u42oQaVBmV
t6Usd3LX4YJ8jI1tLzZHO1Z2oyiO4aHJvgHi/hUbZqpVjpi1zzv2boc2RjAPow3I
AsmiAtT3trGHGjkR0/Hz+a+fxwfE6VwRWgNNnYe5Cj3d3CuH/xBFQeKU2qZvAHFR
eT2cq9vVS4uiXjm2lWbBtD4VTjEjyOqWkIHq74PSiNJf+V2tL87hJHvljpn7X4Z3
cNhMj3RE0yhMLX+OPkLlytZA4ghfWXXvoPBZ7dSt+gIKpZ+voYVxrjmEiiTtPPev
VcW4i3Xx5HtAIoRQbZJLkk6Ixo5k6u5v2SqdUEz2+GmY4N2lEmUwi4zJcNCL78RC
8ESbG9QJs4tPD/AtYHCPaIP1Xt1Iug6rwt7MJk7fVnFvWji2gTViYDa0b6Ez8AiT
uSUPtkOeNtS/BzfEmdb9FXi1ch3VVVlu7UUd7mGSJ17rrqTpqMm2lhUP/K6OumIf
wtfFDmz7aA0j5RlEZQUhB4GgGPTWrYXNpc30Z4IihBguDUz6w3F+kbyxhpiexwQV
rNe2WT7TWWEIcHFKYGp4bTg9wTYE72OqRWw9ZgAHJVTO4vIpOM/LX/rEHvylNRAC
e2Rtz+vrCZHqqzJN68cWIcRxiANC0IS/UR3/jb07WuOYX47UVa7vMIp4uSA6hnx0
J5EGpUeN11pnysCxEftpf9z1oTqXePBSlpe/Tj0rAlIPtBCTQiKwZ0dLo30rbQoX
Mx7db3SYtEyLl36CwpE0AJB2ki/iza02q1Ob9z8wh6Y9rPQVyJSh53slkVE/Mqlo
ZNJ+6lGWE4JyVT1mcyDsbzkk7sIyNg9LWp8Cp9TPIAbdHycQSHVkuyZ4XNw7pdhz
qJT4toVW0RJrypaxaC1WD6C6yvWS3LKH0kImbaePqIdp5FC04SbOT/yVwoGAwHJ2
d0Av3+OkaPONiYaAAm2P15613YSfVpzXQ8Wdga/5JRs3XWnm5vw6i4o+vKcrbBbS
oP1PmdzybuPQztE9n6qG8JCQogBjS8aBQ9Jw8CMXxd+PbSFgP+LKtwzu6lhepDjO
Cqz5U2gprTVfd+f2ZqRDH1nT+TzUzTe2UXBVAK6a7b0RHa2V1CsoojFg+iRgkzJO
9WNvlIWK59BZKJQyrEz1TGvr/90yXJdLwnF7+VpoefdVbTVMlR1MMa4nWr50tM/q
Y/fDqCLQe9SaCHdpW9yl5w8oKVDts48JG11aRz3y8dU+yw73dvXFLghT+Rg+zv3e
ovQqCHn71yzeKjeyZ9kIkhD/z1hUNUWgSMsibN7Klpeh9JF6Y+tAg4MsdKmQ7eVZ
cqjviRlO61dtlpviR4jnJDpzemnUfyZU9fdU7qGFTJLcgUZIfJY7kAN9Pe8yrb7i
XF+o4cLWXqCUDVrVsXYqpQa++1chZpEku2ivsKfovd4oN16vEIZLMvm4RQyzSCIg
HlpWkzdo4eciNSc2Bpg9jtn3D4zfI1gzzMWsjQXG+h8BxOou3AllgXE2B4DM3mnY
eQrnFrheBiZj5znLPCpl5ZFNb8yzD0TnjdtrXadJf0jjzztt2rfueCPKgTlF7zil
51dibjXcC6CHEMtftKfBtEUtft0VJcsXyfe8aYqIr2xFdTW/4pXfNsOi8yA43NOw
U865oz5GezwHX0hF23AJn+pL4HfNcmSC72ZZrjLW25DyE+cdlelUYJLWcQ9oJfan
L+PGSZyJICLKjtRDauozgcYjAx6B4gIE8Ij6SukoJJyCCTASyt+jASWkytWZnFEj
+QAMJG6Vz0qIF9fot6aHE26XhGNe3ylQaA2j1xQcoTX+ti4mpg/ogXccLBIvNW2O
kIokNOSxBSkUkfRQmBYPg3NLsRlTB3A4N2xB6G64rySWZQ0SeE1TgRr47J+0ddix
pd3MHapzi7N/O+q/sahbgk76Doq/SIlOO4h1yVw2a5hGIZM2lBkcLiLT42q4oJNs
lIk8Tfguq+MTWkmKnaNE7DSzvIgRbxntF//KfNqQBdd0XOv1TRQBXxT2YdeSEYRl
g9NxqXNFtfBzfMj7G7gge2aozbYT/ojLlOkunQUY5IkdudMQK/lHofNosZiaK8y+
YvRtULqjYbKeiCaLOre8akyG0rWmskp3iPKtXK+Hr8Nf9PGMgqrbeBqtWZSz+Bfp
jyPKtR9fDsRDJIQMcsfEvvdpWHkiexL+EF6VuObNNw5R+xS4gT7YZWqyc3iy23Dl
msuJS8NldWc+EaoQeT/KkvRJDgKeRf9Wcy0hlJiXICHNgPvahm0SNaTYrSMuLZZ5
SvHQX0MQuhwqbIqKqkPu7Igx14I+TMtR3KzOcx1dEWcku+VHDSu9vEd4AcoUGuEE
rvb+7At042p4YhCYUTT093c6AIhxMOqiCidUBIZquGjVe3TmXe4JkW857xjEYyaP
4ngF2+479kAe3zmUohY+Qg+HnYKGPgWYJUjwPTDl/RWvhvxd0NfAO5sEXxLjmUN5
iZhlMsxuQl/tpFM+hhroljIB1ffvnr/HxXD1SbvZg3uybbCkfr6lBndXqPEM21Zb
NMwyqq2UKhz9VnRGXsF0qgg4bsI1RokcbJg3J5CzZpva2UifN/zYIdLereNRaP/1
GhGW8onNZNPcC8aCHlYyeMlI/kOObHir3qawp/Yu0aRTs68Pgwj++5gq03qcDavr
wqoYBPGTY0SHqIV3bzggTvlx9tWV3xOSTL251Doimq/zXR4adUVBEwSTn/H8H/6r
8xKA0pHEpyQ8+p/XYFkADI39QPjr5uDLCRTZlaAdju3Z89ptu4TZyW2htiR/G77d
SJ82Q2KT//5I2M8db9PgYB7mhjyUjQK2wBIaAapPAA70Li4/P0wuEScR67xleveJ
uDyyAhyPJ9RlF/ybO7+4B9ApZu+uu1zPwPlVelPrbZ+MX7nSaAvBkm5pGKEkpKDm
63pJiWxosMbLs1EJ5MR2OQxZtNUl9MDO1rZwiCanvKJYiRRE311mur4xETQW22zw
xm7hsfJu8M3VX2qqu3Q+MM/auFmdmqqejRbxXTxazK4TxxyLGnhtZ2d8N9tjgzeD
2rmkFTBIvywvpwHAGKBezcxBGlW3nt4UdEvtmxd+5yAbhqVeUJ7KbJWcE6XJZkHo
ewShNcdVLAS/TA1Hm79quMcQ49w4jFc/pcoAlh3il7scrN1R3e/W6veiiTAkC+a5
VEYQ36uKPPcohlJJl/se9WW4K3bJeG4lTeFFEjBWEV/NeC+xwHFsCGmxhHz3Uanx
l7pmhcDMYPyQSXhjoXKDwEG48Y3fncH3nFTEhKwgHZ0MEdfOwF+oaJp2AoPAcnMB
k/guR5I81BbwWenSsR3yGby3to+wl3A1AQt+TiWmVIz8Q5rbGbh2/MkF38Actcn4
TwzbWT7smE0MOnWaYfhc5/QNi7/GAMB5ajWSnmVh87SXDUxV6JcGcVFOl6MeqsHP
KHC5qLNbZDdP+lax+xNmhD/P1ZcnNGDiySioTuzPT1D2bMa/9N1L2D2QZnPBxisQ
yT99eqNCTd7n1si8RaHh+sxCamMG3mgV5PaHoPAlFRSRNGvpmW1PvM1EjD4gzDY9
spveDr2zdco2n/qp/1GdIoZ6cEIQ0qUemkFmAAsr+C36HVPpWNHDet5KQHQyFWck
RfTYfhJI5m5enKd4lWwPgMgPs4dlwQB6L4xc0snOVdmpd3cCCoDyooY+3Nyd05Dw
DHHg19Y2F5qQh0A8nwLDlmFHktDDLodkGDwyK4dNfxgYp0TQnXTVO0QxsHufH9wD
1ragrnGKteVPoDLJlyRBpwPoeee+X91welHe0NpQNXADFuAn+BD8Utgnv1pL6pQA
Gh2hY6L2NcmLc7P9SvwjZIwVBH8Em0UxfJngJqfGZW2kXvHjTvnvzf/E9WNjA/9E
Nu6MYcG8zOHpF/2IVtQYCVgKQ0Y+6OTTUpbse7J+YJU26iFQlZZY52kSR//LnnPJ
odorQ93N1Jxr7efnzfaJYDMs5FnzCq3186+Oct+EjvAM6TrqapLeG1vFWIpTv7z0
j88ZCRrCDW/ZjIDQV3UOtdNq82EFmJFxm52AGlLa/Y1Kprbx6umzsvZ283fB6CK3
KCAZ1BBgGHOolqs+ppIL/SJ5rnj6Gn1r5X6Cntw0PwYSMlN77r7BRB4ltt6ssT/S
/m0GoANmSmMWUwXBMquD7VPB8P8X7YvpARkU/Hmg/6u+u5FOTn902TwaoR5zmzbP
oFrG1riaZfnL/qHAq1euBTfVOFx5p/gCmKOoECHrIT1yb3LjIgEqYof55lMP3al0
oBFyCmy1yAq5uE6GINikG4A5989k61oykp42AsDho8Kx21eG3bw5Oa6ftEHfYlTP
bjl/NoQzlUHEhVPH5GzaA+WYcCiE+AzUdjHNtDQQk4iub23VWKvAN3CPouCqKKSR
nORSo0KeQxi7u0dgob2sRFss1WEssK7cd0UTTYjmB2RFJ1/zMPEFpl9As7tsQJLn
HH4WTkONRYyLG4ui7sF2f7HZSvFRkOnEyGlM9I9GtVwuiSOESEdJ2swPbgxoHg3d
y7rs9F0THDs6TPHFBh8Sf1MPfDsf+ZSznG12JtsO5gqHCquaOATjU0A2CgpoQ3Io
01/z2AFiiGjLJAIIdYJ0RBPPjRHeBSHcMNQxNNLVGNdUGIDgG6abmoPqAtm9PLbH
rYJRMFuRxyjCJlDo8g96DGe4vJlP3GA87MWrfEbz0kWmViNrAz4S4cKxph1jeWDU
c8eAGEvYsPDSpMiH5nY1RfBUI1diwTE3/ybnXmXEpXcmLulTreoBSYAtr6bU9ary
9Bq69Ph2u3i+d1AMijg4T5kSAqdScNuCB0m7wnWCEbGQljsRqTLYb0L7lUMMwj6X
38ASKoAuvwrL49P6PRia2IAEt5c3plE8XSXs9iF5b5Vvcf/OIT+zhFSh0RuYZYLD
4hp+luAt8rIUzxvIB1AA2gU6XA3xvEEgl02k3Q9gQQoQ48l+0jfIJlEFSmW1krYm
cI3muPqbwtCpt3VCjUZurakox0j+M3yqT0ZROZGqHsluxfgQe1sEAQF8F7hVLiOv
bUjggu/F+0DPYeIZrCk8t3Z4lirz33JwBS08H+Xqi4UJZy49g4wLdSyQt/YxdDbY
uwXPTm278rOpi4M9eZShODPIo99XaHZ7tNgaoM+P1d5mYs8rUHFra7QRRntxFF90
7gqKLvNslAsHKK2bPTjpr8mymVzoDp64jrZXhtLego1+XoBcLFRHTs1d7n848kTR
v/U1JtwmDg6ggXbfeCncsf7TCwUFz3FV/BjQ5vo7HECayJ5J0j7On5/X9xeXyjO0
TiMmmwHHi59LeG4srvWpZkoESo1FiqYEAya5qUmbtMPRFqEQS2xIPm4ji+jcjWtM
qJrwiNeFddmRiTnO7VypAqoHJR3Nu4jsEcQXrOogK/0WpDRunjtqvh4+VTtaIV4J
YJolWKi275LxD1gHdT76+koVfTJeSgKTSmF65pwl5FPNc19G3bDl2CYqJLInTjpS
cZzZEV00PlGeXfXuzwc6Zyo9YQUbiRInXsbMFl8TKEJQR+SMPgk9xSaTXqpUeFok
USE3W9mSsOapQn+PqWdySPoyQ/vKvaZh8GGAVFgADvtye/VwMnGQL6Udz9zlideh
ymJYwYadWCAh+J8lynK+4tb2ZKQ1KgJFSnqs0TLf0zsTHZTMedmE6mmalbY2kL4b
06frow8Ui9uvNYSrrjeAB1wQs5cKBw/VmHxQLuYG6ZEO08DrbRRkocuctaXI8RSu
bVIkogjyNsSVv4j22g6sUtEUMDobGL1XG0z2hTo1dIfuKnpSqKbye+G8o9LmDndG
aT24pNeuuXfN3L/dKYrGRcDFddT/gc7J+bmK10qc1r+aVMh5dMF7UOTEBo4sVwYz
SQdDVSJGblc8TfHtuwTWckr/Yi8FK/KbhfzdId9lur3m3kg1m6Tr4WHUkT2AV/Oi
mZfCqVY8K4O6ul7YfsriPrP6A466l/LmiR+sl+2v5lq/VmRPYkz4BjsJUHSYePnk
s2LoVieGe6xXV+r0aI/AsLqi+QLjZrCrzZYk5y/ipvzvtvXgJ8el1f7c3/fRBzfl
rbL4dm/KhQ4WT7ZaBmM4xbmiYEu2LlAzkEbxjAFKjf2x0zZ3ILEWwpm+Sxt5vF2r
5CG6CKMP4ZEf89IkMDpeWaiTWY4HU0+2Lb2SfEwJZt/2ccZAzRkWys6GAT/XfnW7
IogKJMJuzDO8iKxbceCuqXf9E7YZeWgCXoki0PGZ/xfJFBdU8+XZ4KR0GxchwUN+
hk3Wz0Bbf4e8aFFjNv444VcDpEnZPoz58z4B/8S0pEoNaKrYFPT3jcMYYfSPPSqB
3xk/iMeMUyn+N7N8FHuqwQTAnt0SUSeX5+hx3Ky73fAOKINOJUzK+stYnhFMzVCe
VeFBvRPn8CdYctAS+TGR3EZJV+LA3RqCUbfAsneXKcIFz0w6ALxXR1RfvwX+AWau
k0de8TWC6pJ/m9xqeE37Ih9LfI3g63FhnjaTpUw+3560EP8cSp0Ct2rsY7OREeyW
0oPicsBYQwlmFrUCSYANMej/V59zfjsbUAi2nXDRnFR+6SAIvBgkpI8PkXFH3xqb
4rIxUZD6DYQx7g+54Ks5LeLJ9dYYBkQeDGqWSQOsbg/gI52feRLQb8JxWLMa4tyz
KN9fZXNXLK0wOHMDifb1Y5m6IExeDNtIs8qWH3f6C/3q5bdwT1Nj9Hz9JbY0+RH2
lNyr9WCc3yY5+eoQHbYTCrBAN1ULci03ZwG9dnSB0e3pEQgMu9pwyQrGJaYQYmHG
OvIDxsDuXfE7J8PzlMhCByphChEZvcmjepqrH4ZheOiv6FeSXBOCjzyQdUWxbbpE
8UNuRut2+xkmMSY/V33GSKbBkCI6LN9BbcsWLQlUxuofr3aTecH9uV26DdgYlZ9c
iH1jCMhGR/ZbbXtGkV5eZQCjFL+ouW1CRrTxw9Y1MsUMEKYR78HbL+FiIlg9U/ly
TdpP9ZZ/V5GSV1Ud+gTI5jvqZhSi9SjmTaiElJ/PcMIRGaw2GPijExnTHhPLTRol
6DPBA6EY5bAsV7mMqYUSII3TwIah4qOC7+Kqyb/dzLDjdN+ejhisXH+n3vUPdu/1
21BBB+8X19VeVUKgY+yLKpAgHFSdL36FJhLOvlNYLAMxXCteYKSHMQRMRHSk4XW8
BGH6OkAK7hwcIgPPRsggllhuzx/Qk1mIpr++UmfrlE9k74GunjYF3dJopmzzEL3e
q4etJNWC0+aTkOOtRVeWqakcyljyZ9DamFm3xiNECEpLz3KBLpEDDVOXJ8+VVC6D
av3wRguB6LE7nPYVpDQqxw+69xLjGngnxIAxuSAbICEfR5DnlHWYMFuYf7oMl6QY
e8nH+kYNMhuUi6vjvD75TsMQl27PIvW5n1JxznEqZwXk4i0jP7JxEdwukH/lgjcu
p1r+K0q+c+EDUKws8KCz7uC4kM2Zd59R5lbwe14Zp4iX39AKG0BbPKN9vp+0avN0
YooKDJzLMhQ84X2xP+Cfx4MuLm8y0XctaB7bCL8Vl/9hIFz64sFNB96ZR9zmn+fH
zW9uG7ui/ypCYLhEDcUQkd0BCoD4yxVfD15G178m2xvzhg2YOMXBhLDXWb1gbUUC
C3ht21tUTCFtVxZgDs8bhceOQe6knjDHZGqPQ6T4Ub0JTgepYlNLyj6OBHRkRi2N
K6HJPNZV5/nSVO4yMwW/b+fHcuwFSR5LtdcCvYRira80v7FGavOJLYmvITspKeLn
WuaT8zV04kQJsixfIWb9IJ3kTmSM0BdLqzkb3ZanmJu+EJ+VjDAfTiI3KTmuvxw+
KswJ2bI7Qs+N95Sv3GnZewP91xO7JvxYkhu/dvI7xNxpF6yZWuXqfPjcShGiZNJI
78sGdNNd4wT1J3mcKQNQy7QG/3EVVuVJ1EO3xYm2vDxyubuAaYx+43AAGGPvoK2I
aWfr0eYIKUmzn4SzsibwZFsKiPn+uSpfgE0Mz1YGBW2S2U4OJldT0k3QirVuIlso
OrVn6CVk5WrNAX3QQTlUztD0FTFd0TeNVMmsKKVkw+XKAuk9kPsXbjfJjv9Tfx8S
g807P4I6kJLyGYS2gYxIEvSG79DcN237Sf6R3Zbtw2RUGEcgKPHBBJaRbWxb9Sqn
AAOhZAcwoYOjRPGOKnbcHVRRZx5fgTgWqi0nAjVQmDR1WLyDirEWuvci9XAUM46d
0RxzR3mhZ+z/4MFFMSg1A7RcK1KYaFP98recJwyq5DHR5wTR5ITeiUtre+GSBlwI
VnGt/xryVH+2DkJWMlvFanuGLYy0v5whiIZ/hptyX1Eljqf8o7LU/bQNQC7e7H+G
DE4XLbv64NNur5ds+UKK3MXeKib7CHV0+pWr3obX5eH0ofXZf7luwN58s6D9AjYS
AM+KW5bEOFS57nmpwORzzdkjycmcy5jqYk3DRPF0i4CAGhMaI5hw39K290D3V63x
Y1q3Tbml9l1Gm6g7N8FBXtEZf+vaxoTC1E9+2eDNP5sdI0pyUgoWAaMw3xMLgZTf
efjD00lRe3W1Nm8v80YshXpslKBrKdNtkR0BMjSMt0PZ6GVw2Z59OycdrySx3x2l
E6Ozw35fs9DJgVQ5ljvWX1cZTylt84nvuVOmbu3aT1lIcmbR9gn/eiXZ1H+v1MIp
S7Dij/+5Ddo4YsHCOp6y3qZ5fKx5GGhlJYo+CRFmxocX1dfIff+kW6eddzTDDgBV
fgKGmoVreTYw7ev5LXAYaAww6lvKVPZ8LD76iG2CH7XHBYed01Z/cjBgQrIJ4r33
JK1guX/KTCgLygIhyFzcPdGr/ZpBLaNlmV670Yq3wtBckDgcaS7/TnTM161H3Ls9
nWuCuXUGeWL6DFf3nMKasUCcfuCsvnx9XqrpA28tToh76TS9cYGanWw6DdOdSAxp
3qLT+rdndif5ZIVHrlgyNAxlGAmRhvtJ7eZ3662wLl+Cma6AAS2V+hJ0dDxfcv3k
Yfv5nUo713NYrJ5PluU91D1mf/xH/wOoIz8+aXFamsyE0bShMgDR9Ro+38oHNhxN
Zgiypn0GJp/2fg5hMNbXodZhbT6m/5qw8cUPbVSjeERsZOEmhP2nDJdkHB0hmmVW
oADyY+xF1qjeDcCKNDhiJ0/D9SM1aL0xQ2QBvSSmPhpCINLmbkRKBNap3kXlAw3h
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15696 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
8LkC9eTW69XSSgB7cGeNoDWUfDqjLirpw46YWYY159wLxRHst6VNNdZb1q17TtcV
TtwM+aRxDfw46OHAW4oVUTLjm+cyYfP/Dms/6laJ9el5NYviFxBakXeev1VtAohf
50YF9+fIOol9UvWPS7sGiAMOIA3L4/gppUweVFOmugbzY68MUnticguGUfZQId32
XeLbjh6FNPK0BotpHkD8vVRv+c2JQnNv/PHKbP82fq5RP42l39HzjJ8BLNI+0vLf
1unJ6Ypn6+jBl5gS8OO/ePPYb75qDOgmsKKLzfV8cpwkweYo26gZ+2N3AVTmwy0s
Wng7T/18sR+S7wStoCyDY5rkFE87sdvagudL10BYOAHLdJOQcy9yJNvetYU/LLoT
RQCohHTw5x+P9QdBdOfUhf2mFQ/+hJ+r1/FU7DVbHdIT5pj8Kb+I0FKQKEP2qgph
aewx5lEn12BYF0YZSQv3iJfQQpQrbBM1xDnmrTCeAbxhZ7vXUOKULUDB3Y4TY+nO
y+LW98xAysKZmMUMvF+S1g63c1L3lMNWS8P9wEBsCxQoDT8zZXoL6u0y7BE0Kv51
p1/4mgnLc/wFmipeBbhvnGm+mtO1GLaYHcl086NPDgefeRXwRiGXFXz8ol8td4zL
HMbbfoTiAYcBpUQQrzQfNHlEUTbaLP2rT+xEkO6Yz5GhEzOc88yrwbjesEBnqxLH
QZNCjBU/PDHHX39BrLJjogNc8mDhmZoi7VTGMPoPjODZmzn9EYu+vzUPSh0jIPMi
VRDqLbvmTFIiD80p/x4vCiATQ7cmxVv7edvZ2mv4Xk2fNFhOMU3o1JRomJfK7YU7
YjDz+/bWcpvXFmnJ3za476F3sZAzr+ELQnkrlO90ajZ7cOI5j1fk9Lr5kboMl4v8
F2xKtAnmgQXQtkf+0gpRApPJDJ0UX9gZWtPEeCmneF4HGnPgmyU2MXxNRA2H4Vlz
OVZQJN6XA3T9qONBNtIJr6oNrJfmNP200SsUMjhs5CC2FLmmNOO9kOIqBe5/tKNR
TBY0BAsZ3dmVojWxdYJ4mvwDV52a7LYGmMxzAJadzbYRpAlQH31IizHkBLkUSOF3
aMd7NuQCztKgkYp+BAhyv/kEXxwp9lqXl21JBLWpcLOh/8leNTGwQCXINTd9ZKSa
NaWFjWmF0rbYZ+dim+qP5TjdRMaNEDbDJLX7llD5K5eMrSLnePrYgYtBmLPmoirI
Z5H/2DHA/euR4PjRpbY82igXNdSSCyOQW8d2JnUGE3gkVKPU+ojmk5DK0RRZKSEq
rZams7D1kbidi6NYRX9XC+nWJDRKWV5AIclo+peCWqE1BMaonqYoHCT1UN5BagMt
aQQPna4ngFl7IyF9uIG4NOQzS8gsXCK/OEh5gRtCzXi09TvVV0FsnR2s6MMLlpmY
ZQxwwKDDU38QPd1DqwHL3/M4JXEJZsrxUW+wG0150Z5aibxy+k9JLwjN+j8SE9PG
w+27VyUhJeHLCegGqxG1RDYPFRvTG1v6zoawIZCIpThuHkhwk/7luNIQKgwbvcKg
J4BJjDhVGguOlCoI2LMGqlHce5eAHeOMSlCEuenp1kj73PyetD8f0O8bb/mysjcR
VDTMmatbUlUOmQNmF2bNgp/HotRoaL8QvJyD/ASe64MQCL2eJCmZy9Thorg6zSqz
fbal/3sjzOsdjpe+xT0vP4xPCSkE7toyhnTael2goDl7WdqQF8PNEC1q1KzAvJXb
zbRRa6dMbOUnDSL4aYZKMxDaK2sYRRZZr9s26KxR8TZqgzxed6ySQeYWsVvzYj06
7xDBQteScgcZ68q6LGQL9f+VTCmMfiBUrj2trnbcySWPi1pT9OEiD60XCmlotb0l
OzvvnKBqLKt1A9qAusaVAFsGUUd0d11voDniQr8ltvH4Fh7wxiParMFLPAu2u5ZT
QcLog4SP2QwFX+Qbk6AlCxDOxnBzrZ6NUNv1JB33M1ypLtf1wYNdC4NZasjJP5qV
U7iv3LIl1oZ+pDLtAItyZPi04nh9w5faLV6OmSUK9WsSfeeJ+tn0Fkf7p8dEuw8a
fVSHRQ1JLhVxZ7dDZjvBIZhj7pgKFfvNeBn0SZi6uMwUVIwiXXG59Nf1Zl296URb
3pJ/YI6ie/ZwID1gtZnl1FmJ76V6ex1vzWpP1q+yasW3v/upjazfEAUhPnfZUQu4
Fwj/aSgl5eTVrgjUHkPuqRfivLQPw5Glkt8ltbaUWQobOl7MOznipaQfDEGFxJTQ
vCv7IV8f8SMsbua4S1DRrTjEljwmLKt2J/uOH/NkOrvjGf7FnkHq8IgET3UFLRBb
5DBvDluEWy9wsV1LT0SS7foUR7WKagSGvH1jewgc4XNBu6BpOx2TZgH98lgddFaG
4B8ANRKo4VhZE+mQ5pDda9Yp24Z10KKgFSw3t21DB9SAGSrfl9O/WF37EIXdeqLv
rCfdqW+XfM769WdcMfY6MAF2DC69pVyex5L+z0TDHtTq1Cv+KW2V7eFX/n/6B3S4
/aaogPXNFhk6xfMaVOgs8UVj7KCBog4RxYm8QDjpiGvJEF5RuZKONIEUdm5/aTof
oA6bLYKHiuolxipbNqSPwDdra1JCkBAf9KGOn6FNesxkM3CgLA085vbGlkG8ZrLw
9o9FqMWenCQSdffO8KHmfFPYgWubjF+EjgnWFVXO/r9zDzBgEM9XSzQNRCY2rrAw
1f9KfEqa8wwm6/AIU50dxIsmWuh6uWpgRJudBPiBZt5ExZhijjVTve6ber20xJ1L
45mT1TSQbbJm3Yg7Vxe7wZPVs+mTqQVcb3Rk3/MZFKUmxOtoCAgaVBKRa1+ffUhV
A2bZ+F5LuYIE3zvbxYn/BqLX2OSMmkAApNLSHEmLkZLWUcLecRMAM1/KSlFmZewU
a15SQ6FXvqqGIasALT2o0+nLh+idyqd7vEUi80HU49AqQfeMAd/Qez3CDtSfZliM
a3eUnUzIa1rfzQOw5SlNNyHuKj43I/EJLVAYmm9wayHrLKWxCtUTtxs5ADWWxfXO
FsvDJ22t6h0Tx2Pc5ie9TWj2p/q5HQoGnAjFE+kbLOPjgAxR7nYaHZibVRszLZQQ
TnmBCqe+H3JSGwEjtGbbXPuZrPJbTzt4pTkgs9nMsNiFsP1UvOQTLOSKk+hc4f0E
2JBkTEgV6cMT1RfO4N6NrFazOHk1LvAD2ZAB5Ae4VUgELOL18ryU0xANnpZP3PhZ
Bc2yUoIockhXTM6VAdpqf7yLMAMeDCAsQHbRi0XEBr0fXlg4FYU+HqFY7l4nBh6M
ZTPb/5+LC3lGb+3NYHsKMGW3O3awJnAE/c+3UavtXndqYl1HwNBCXqgPMroDxdff
dwpn+dLiaqwZoIMBGNv6v8zXQWxcMWMPfkUh43E40rmmboudy10/Iq/bG1/yawkT
MpB5gn3M/ubSMh+A2iXH0n5wBSAQKpfhJJCnuXkBMAw99UMX+Xdh1Srz8NcneD5b
3MRxfleNF7UJICDyc+xREMSLuGdbMXoICTMVObpxfujGjt38GJLf34ZzLMWkIef0
huuIFx3e9m83iuNZ9GsGEClu6SxOXl5N8Pd20ngip+uRN/EdZR+92rWbmaARw6G8
RifyyflHjq7XvDzJ5uJIcacHKhyYGPKpzOO0LqhsNo6DM5Vr6p+ZzL9iHSADo9gv
WhPJsjO41ZFeSnwnajrbEhYOWPnhQ2v9IL7VKtCnU9G2jldkGlB0iobxdb45NAyC
IxMaHo55gRctI9Cep+Mu9sEqFhONFMRHYhBVAlUhA1ONOFtePwmvWRS2q0V9P7hB
Cz3LgtQzs4opblZ4dS7eNGk9Kt3KxjXKfIwRxMT2/CV7KLanUHfASYli0b3Pav+8
Kq0ULQJWYhpteFXy79R4OXbp6g7uWb8wSa1q8vYGa0dFAXh76HOhZXq/BtXgPRST
ucO9R4gB8CWa7uDQM0LFl4asUTFctT9+x5KM/wQvwNsSObCBZSjyHZN5inyHPSmE
RgndtLKR+dUqSi/GNivlTsQyH5LMXuAvXRP+60iXqq73cawzxwRluagCAvovuFiw
iMZuOY/zex6hqRjyZbSlBAMsik/HATFW5RSgTNEY+mwxgucEcoCg9hBiEspakLp4
9SAQ9rPkZgb1PgL/qBUzzUShElOX8Hlsgyp3Bh07ZhTofheEPKLZV+yIPOk9pucI
h9F+793uP5XQ1ztGLkI3ngIP+6odGrKqqn8MMO4XXGoiARm4f9OSoza1MG0Oe868
jEHz2bxEKHkP7CkMg+xrwyMGeQcPEcGcLI6vQ78y8JazeHWewTM0md4wrQiyy/Mg
86d65GsYKFYrqLrvkZ2AJ8XBGFvTljMLLyKoCEZ2hTP5/JUXZ5Fgn4x4LxOn6/C9
oMxgHF8p1YoeaS4gTzkXzQgfjw90VBbAmWLj062BECP1qmao1LNPxQ/RynpFymQO
w7KIRCXbGI1WdJA3lR+OVhgAxVivzSledLKddOqGTiPXxxROdch/TjPkdiTvP3nH
727DiEXt1U7rCHL0/3rXrCuoK3u7x/gg6G05nWON79nknVm/Uye7b5286XAcSXx7
3MaDu/DJV4OTCw2WlXrBL2ZujxjhaU9HewixxmUJKyMpYL4Eb6xPpsCdn+5U3iOG
hPfo/y4AwvUFdNW/NosKcqLaoyewTzpqz8iJ6TRwsuvfT/EcCRc3ryAJHkNPkjaq
YjlxWAgT2JIlTJx9tEjCWsIa02M0OTz0yRkZbxolek4CtX/2QZRr+f73LGcpyDrl
NAbeF/BFMQHnQNH1v+z9eHJa9Ty3bHXf7K8YFpTA25nlgItv9KZqhqnHZFWKf80N
4vkcKfGKfMkBdJVv524q/FR7KM2JrTXQg8qnwtrw29uUDYdqEb7wSE/jgUEqqeQh
7DiB/SXHZMc7Fd1YTFeJxxRhOyeuVWg5hK36MP6anOuY8FiH/huLrlYBdx5H6BGv
X7ipoKKe0sJgmiVxpmcI9t4lRGkE3XK2SB3FdJGmh//4nfxVrqxiDlLSyRuJ0pnQ
Xr5XI2aQeyCkM/SxA8BII2uOMKEFyyFRFphkIMoFh5zpy2RlmGgYezvDIQB8Rlp0
Ydm1mhub2u4H8sh/3vWEyWhVzyZU8LvNZvJ/gp41IDS48NDhCn0cBE4+4hh7++yV
Y8/YVvKmb+4hx4b1RTmHMfGKdEb7HRK8JJLXQJ2s6FUG/E85icNDlQz/y5vuhJzq
kWRT/ljjNRGUVib/hFuWUj7DqprI27F79Q9RUq/MWg5x+eFrelDxhumQKzW4rp6E
QQ3l6gmuxNGD6w+Z9E6/tIwGwV+ZJIyBTWoiVvhOl9b3rC1N0CTxlMMxoQfG1rwr
3DB2XjR9CgjR6k9Xgvr/crEmokyvYHDl2faAK8rP8sUrjnuuhw8P0YS4Pn4vDyVA
wX7eU7iM+D8jcEh15WJ9OG1/svVvWrrzRHPLLjwGWRRsfzqsY3fhSpnQvVRZ1tE+
s52LjaenlGUEUDYFBw1blqwh0jKBLWXjtUhodPndwokbFDvDl1z0va2FPXwySkFN
bYUAPRXMm/qB3Hq9LNpvic84GRjXxNyuLPQniVTCvHoZoVO90bV7qv7UFKtp93VS
gP/PIg4a57Z/MyxcOaQTrSGntxwiVfAUEvJBna1sFlU34kO8qkyrmPb7Dubal6N/
Z6X08XF8j0utAloJLuwh9ezPRJkJgJCPs/od29UUSJ/vHj/6L7ZspOB2r7IfNho1
NtGwJ8KRc/uM5b4Fcv/0v7Qzf1aWo60TQt1Hve8lwn1NJPL2e5GVkVADACDQfHpB
TQUC5INPC02KDsM0F0jgBO7df4TdRgErFH1QANgpzIVFfaDqjQ9Bkrvfv/MeI+V5
kXJSdqoU2GsoC0n9zP9qWuTNBzzW/ZoPK3II+zalCYr+qCGr6RfxVGHvtqr9pX9w
ORgMriofCcCti8gHAvD49UiWu3SjhB5iZDuja2eBEouxGfPtz0Ww+B7cEFNEttjF
F1cTA3a2jCi0rcnqnCJclLcmzj06KEK5FMiheAdWNrOMmG5ev0iT1G4zc10MZk1u
XkAnpNCMSBqwyX5zb0QDnR3XpzeStSOrklk4jpDamfXyeKlqSFh/gEaGrF1tWqrk
qMLIQdK69lMjWhnyBK2c+mqkiPix4L8X9Fmi3JMgFAf/YJ1C/CYuGk39qbf6FPR4
/vAvZuB/QP3nN6roOi/Ly/GLlkyA7d7dA9SiqRmMkk+X7NLwyMHe9wOoFEbPi7Uc
tBEAPc3nQ1MSjcz24WYpZuvLKBvcoJYWM6mkfllBDn2ntyNtEgOJsuDeP53ayS8R
Y2WyjkjFKk1OD3/1WM0AIQ9NnKjT+HKNJQ6HtePB7gzMe12npmHHA0eCrbSWv5ZF
mAnMstqJtG70n/7eejc7E85lt1qSJ5laR79O1SREW3A53S87YOryBz0095OJnemu
RuZnoddOan7RQ70iQrmF32Ewzci3lqpX9dALioOnRgTbV/EGUxpI+SU0aFChO/sq
0GdJNYZaHlrK4zbzkKnX06r6ct6Y8PfKJSNoe+WDz9fgd3HaVUHBcmyM20UDO2om
I+BPTI++Or/pq4+wD4suxXpkSHC9Z9EAfFGxU1Hy9ySYpMh0WqRmt/vc9D0UzhoT
gUTmeR9v/sW09XcDQPDgSlDRYuwlhILvWZSNC4LawWiR5ozUZIGirDJPp2dt75Nv
Kagl93rpRjgGIZApPHA7pFqKaGQAjdFisO8iAyJPZcAwgZy5HQe5IubwUt7CUXHG
9Z8TsVhfxF8QHDfEt073eWWzZsJqIth2M3OmXk6TWisd0IWeZndF2LcMQmj8vdes
6op+c6UpsRHUYgvTBtgBkNRpLsFv09tndUhHgLPEMFH624tqFDcBxKinwimJ1T8x
pMOXihYPQ1IagBFC1sgL+H9wfaDsihkSl/Ouj/0j7r7yRdjzB2r64+aiz+RNyXy/
6x+M08qhCaXWinxxbChU9Hb/T6BPH5H+RnIG0wPKuk0B+SCS0ALAzeMu4m/lTvu0
bgEW+1RxY2J1uFlJKZyCSgDdvQBMxKMCPQKfzWjjb+ELF2uGYwKhkHFMyBCPJSIG
1JjbqUnpvST38v0OEi+DQznCUIypNo9WeneQ7DnuHP1PLIHN+TCHE85axhhRNh+v
PbzGomr6kBDuxAfewZVoGxhqe3EbpjdtelXDk/Dtrm6Xy1qUfGDZvPg2EwzBOYUO
Tl03db/dxYQCTnn5hp7LeU9gMGFJItaNbhRIZguQLx5TmvpRtrfpJM6M9OOivV7k
KlRo9mKeVupW791T02W0Y+azAU6uJrQ8D8EiDIcY7e7cyiOKngQQlXfnQwbQHQ6d
H9RSFCjyWjPe8egmpw8XZb57Km78cebP8NtdyUYgAYvItF78cd+DumseuNfXDnz/
Jl4+VjFIkjqpZwFLhfuFXPI5n3LQJXfl338tPsXxmf5Atk3FBYMjRmxQunVWkiOD
5HmIKJ/OhzyfH4rY48X9mQWqU0r2AS3pUA/ER7vfMaS5wv2yb9e6xYc0GWBZlDBi
vJP8PzXqJMbPBAnKVVNTRRgb0I9ppzfAiLJQwCrPiTQ+sHOe/7qBwYBDaq25Ksgd
FAo69XI0OiIAG8BSJPe7mKRMPFIYiAhRl5+7oaJW2rV31Nm3JIbHzNV7t+CdA1Mn
e0TKyrj//P4RcMpU8GdHSSnPRjgAupQPlHOhB+1CHuA2MK0ZwUc135TMu9v4+esS
RU+liWIdxv7apJAsingj0+GtJTybLlg1ieOhAQe37tyK8zpA/SXIszu3Y8CsG90I
BJNgT4eBMhiq3BOqxH3HZ+mPhXqfioXn07okfarwYXFUv3W5ZNmU3hCL8Pr4+rgA
DHgWtWaWyg7TlVJFsY55+se+9AIudOWCtqdPIbT4YgBC06mBv844xqY/uQNdK7dx
iGN6IOMPdmHq26TV5c/aFYEHvQvPqyaHua6QnpsrXiiralx0FdiKTMJjVjsTnXQv
Ovg5JH1AUGQ2lMN4aGNyEYRu0/IhcwDshBl91E17A7XzwrS9oL3SzvB/n8hFhAps
0FkkPx8j0DAIs/QaPPHcvUeDIFlJTlLFYWUquBnrNuAxTOOYkJ916v5amGwIyzQh
15NDquBc5tbhVUk3BE4aQdxNNySqYUttOAWgKa7hcbTDuXVvu2m9yPJb0EeEBFE8
nsROjMokNBUHzhg2erYZornr4NmwCIjCO029KbRfZiSgG9jrcXIeIIdCLrSJRWGv
TnJgX0ZTkbbVcgg3rnh4jyeWYcq1g6ekVcPyEnPhi5sVw4cd/Bt9tR0RLuCBeohK
wioNcaErdd4qdlPT4QQq4RMz7YPzfYSfYKfJzN0F5mBXdaql166LZL3nz5/PicBr
S+Ad8jZyFnzqih+NVZtmhayBXPti3Z4Z5tj4x8I9vSWe5aNT3f0xAlVJ25gkBqMG
mRyAWF6ziP09H6VaFswX/ztredC6uKBsG6g7gXa2aQhFUTGnmBAcexetiOu5bhGn
ZoY0u60UF3huRlyXjydp7KCMyzZLstsDp+PhQhkMMvTy20ejfm9EYBpEI/45WwT9
sZX/1sI9b77epgRlupH0OwKf32O7FZCLxX/OL4FhhamwcgZDaZsffQJIbgDpSIJz
8SIhCb8AqVb+ZO+2Cm6BM9Od/Vj/uiybqy/QYuEhMwrrOgkleB52WKF/u1gDv2Fw
VfX0qoEXsyRhweu5tABm+MhB1Aqn5+W8kwkhxSJV/3ozt2I5ByQceGU/zM4om2XA
n6r6jyofqB0fVKzp3l8DVn3RAayrMx9frMXlTQsI6QUXhMSMiarSdllVOLObyZkO
qcVG1NHzeIA+YN4WqunMoGVAFZcuaG7l1HNUm0nEbgjlUV2bXcUDkxCEl4d4xIGF
lL+iee5D/YbxYZiY07H7a3LQsoxozcvR8nnxAWsk655W7rX124FKiQiQdcMdfU0/
fYEJYPqaD7318dj4qTmGokbFOXo6dByqiWNu+wuhgefcnceFXCoGf/XiJO7uNZ02
awQ3zN1H1hgu9NgUHXYwUoOAyHMM9E7alUHetcuYojxy3jqjMllpuakDMqJ1TeMs
Ru/HgPAYiau9yLFZ4f8hI48+TFvTAZ0GpdbVnvR2GqGG50bSO7FaKK7stiYYxa0S
Hj2Q6GOwLC9TmAR6fO4qb+cfcEQhO5rXecj16dllOsZpoaPHk25HFoCTYZalD5+n
x0sLArshX6SRWWv4PQLzfxi2AQojp3kTEi0b0cl34XyRe4qwcdwntolbIWO74VyU
Uj/OJExKLsuNomd4cMD76Bg2WBUumBb+ZDg096kYxTm4T/0Kj2V52DiicrBUhpw0
tusdckHQtqyb8U6e8HaDhOIbuzmAzCHZ7rX4IAQYvQHXywjm0t9s4FeTdWFlmo61
28bZzI4HQrJR9CQIUyBoL+q3/oYcG90D73CRqQu5naPJ6o9UJAUrYsK2b1uG5ANk
q1Ezq+K2k9a+hsqM56R8mAUp3rzmfcS9cy6vsuxhfu8Vn1jly6Bz86H7AvnFb1EP
QwBi+j//q63enWVwL2JupBoJSY8nrzjHqbwo43W12+qcaEoHua1yQKB0cHNNQvwZ
3q1vM3EGZ5XUAphKOctMFWCWRve1YBI1nl3o+/bOwqsAxhbJRHaxQWcVUMCPBF+l
RqIeC7jn9bzGGE72E/Paism5isirotVEMat9delZco+uKZojd2wBC7Q1l7eC81kt
Pj3+16pM3XKwMP54z7vs4uN1P6HtVGKYNCDS48lGRmx356K5N0R+nyP15HyC7A6c
CFk3cK2MuVFHF9xI08kpqmLzNFTURraZuLxAR3rNc/6OMmf+VlVe9UaG1Ycq7J1R
5WDu0TpMI0AHHHsby6SK57ugbfvrh/+sWvb9/Vm1foSxvWHd+LwmndBgIaDwvS5i
SKMbytUzO/3JQqfq+08KH0HwXYCZ23s08XonnumcHLkfI8mLbBj3dz4qEOhEnpkD
n9fTXdmmR7HEv1oLQDSf0c8ZdLqnPoPzZ9xew4q8j9ucn1E3/sdHcb8shD3jlpzu
3fVsc0xrnU7bcZX3qkyvdV9B+Nq172m0Dz2KMS+pZfZcyOOmltPUkZ09uetwtMHb
9sRgM0KYmApU8Gul7coasCJScaT5+3hNrwYX54/Sh3emR7V3/vjdnOLaYslsPJ5T
rXJUAs6aFBi1dzt52jxw6U4USY9VAw+Bp+0OjlVThHrAKZBVnbo27f9einoIO6kB
bRdlVTguqGl9j3S7Vc4e4+ehkNqOPIrCR1mQOP6QVTy+2n/10+i8gVYLuTR/CJYc
Kt8t3GgxGbxVBgLERbAZgAH923tyN4ZhCb+WopwKVbpzOQz2RHBm91kxP/vCqbRI
uWbQ7sKWDos8r3W7Ii11E04p2Y0M7ucwCFlivqwi5Qp0FQj7Or9hqdpXsFTs0c/d
yuHtUzT++XHWykvdyrZl9RXFly8cZyuQDxe2n+p/WGJhEfe/6zy8jrLwOGZ1kCvf
9eNSAWgdjqvv/hzBjuJh0dRpMvh9nbok7g4M0wrX9k3IsP5qBl7xW5r3e1i82euJ
IpTUz8oHY9JFecP27UDfQ1PKv1wCgHJesrbgedqA3YDmB0NczxgavmCrfiSbyhLd
xyOKpo3JJavwCiS+uOXiEfMmTwMFhh+DrXjCYvgtvWC7478LRjlqoS0gH5dlY5H/
prT6goFA+31xFwoTRP+siQzXNaua7aYNIi5fPULmvey4KAORhwNvgnwpUY0QH/qd
qu/DJ4TFtTmaLlK0U4Ft4r8acG8Mk/fkvGz6IogokimPsNUbh12FXB9HsT/Grq5Z
dt1Us2s7SvQPxfgqHXG2oZCxSN7w6+I/Ks2rXhWmG+oZIWvBcBULJzcsTBTceeOC
JGyAZ1FNHwl4nUGV7iFSUob3PeKR+FtZuR8bYE+idwD94fjCrZZx1jEKsmUjWMo2
jVO8FiE5RYDGXJevTmp8EKsEUtHld+emFd5yCu6a2rrjmpNEQmiyDLuzNHt+3VjR
cLOna+N1hBcFilf/XNSDklZ8ntG+MayelSWlObTPlqjA/OU0SCvKp3WQn9UUT6R6
GV2pKKXv4bPdjCGBzI476+b79gbSu08Z0L3LyneGexRwpYZ+8FzQMW0kFb3yO8v6
A2QHpxwOKZzJ+PuLXqANBbsMy4Fkjrw2g9Ed9QUgM3uoazONtV5Vt34nXclngGwF
1gTCOzLLm04wHEoQpolDT5ChTAHcWJYs63DH3Xkyp2FtUzbviXU3wNebczrimjDO
8mwUwaRrgRAUnfcsM6yhkYKZNMg6UVMd4CUeQ0DZ/WOcuvui9x11NaEf3IbExFE+
kKMj6hA7f3LueHYesvwM2MLui9o7hGZ/aaOxhxnXau2cmfaybflIVpR5x9qeZ/sc
BnAK9ytPUiC9DlVTqYG0y83R6yIQwXXljvsEvROXEqspvAafC5ZMwbcdFDKnLgyV
E0aERBeNodPIkWPg4GKuOSK7oTm0PZAMWkPNJubWpqp/9bhqaEXucUVibt+2gIku
SOgT2BTKNrl2P0n9m+AbWGJhyTGE9KXyZFmdNY7CRpAVznxIf1WM8PxHtMh8iD0o
UQk4LehaQ57N/933H7iRAcKGHJBvQ5U0Ajw4ZpYBRvCy9Bq0sas4MAwcqc5k1ez4
zWumLUNOvG16UqHN5NgiQlxRMmsDeGO/Dl/H73TnnOgx7OirxR7qoyICPTS4Er0q
O7YzhF7hFSbGcTzLFAAC+3btoQu5hA9LUTB6WkStdh5bdX0NtXyZ0M3oPBb8HqYy
HRpeudJUFYEKGWawk9yZS1/HfE2O5PixSsNeriYc8jzf+HKFjoN82KaHLdUQ8ajP
HVt9zPXsxK6xc7k401xX3PiRQEetbyZBFoDOwmcOV1GhGgW3L9rdK/uR45JlGeIC
vaPu6euSizGfE/JEoyNxFDCdaWfBEZGXK8xbfMi00LSTQ5J75MtB3e91CkOp18dQ
cPe558XKjVc3rD85Cr7lpcove0tFO42epoN6YSzA0cJU9lKG62oEMr442AX9QCw2
Lyzbhjp2RO15blfO2rR/6NytdSb0AG17toNgZjl1xengOXh5dKVHQTWCp4HfId3i
Mgd1Q3YScpRmkvk7me1F22tUthGfg9mJuWT0HGt58fFBLtI6mo219P6TlnFZ7SOL
UYXD9/JYfVgpC4fIqlgjS2JAo4vo/PyO7zJTw2rl8kwj3BOBXbMa+3ASf1Opf4BE
JDRrisVgVp3Z3oG15bqCTlBnEniaMwRmOQKiiBvV/8m8KjJx+U3T+sts4mUmLAML
Fa7DNFui81cC/6JkWYo0LW1fIldi2D5TWPIqnKP9HQ1nAXgk4Pb1Fe3t57hZmDxw
uyH2JRoAHG71Q0iz4gfzxs+2ouWOzFQQxv3FGxsUdqjZ9aspBVAAu6V5Mk08HA2Z
YjynBTqKHDTo1wT1QSWBDvO09gxiZGd2iZG29vXoAA2oedbhRHk98TH873bDtAxj
+4b3al4Ww27QmIXqOu2dmbZReVieuRemCNtS/NYPsKw91lyOjhPOqaniFXDSqOFd
xvlWcwZFs4gwJbatlC3qJHWwasg1ked1eB8W9y4RJ2pXh/MLCD4LWXPdMS6dQh8t
wqJsAOsor39IQY3901zum6ah7PufqYuweq7DWTOIvWBe+UMbyfjZs4hmjjOkZ/wQ
YUmbw4A2zmSRgEvoGILmkXkrr/nZuw8FCBMT7BXYjpz/1JSlKEtZ7YNserAo1d8J
SNN3RFJpXVYcMQc5fPIFeaMeJU0iyFKQiSbFGhNVlpZgMKzOOCvhcEKCgxYCHe4D
tyPbpWsWg+84i+dbA7MTIHzWQyMUyk9fTWRCJIRNrs9BXQ/ZMWSvPY3t0++ZHflF
MrKOoZe8dNGx5bzzm86Y24UvtTWVol7ftG/dfznBsJKN+SMzLR9mnl+hkGwoFnYd
hGjhqbzL+u2woFaX5UBUgo10xdG2VXabT18Ah9rWZHm5YvbbtUQYecy8qLFv2fAD
Gn2msvoQusr8YHMwhVrdbKTJX6qurwlWGZxAfuHm7v/8X28t6PBkEjgmZ2bfnvl4
WR9Rg7KLeWwUawmznbQ/GhuHa8IOGa4BJaAmKxkMUpV/TWRE1nsIDvHfEshYQK0d
JByCUlIcIzCtOZ89SbRfdNfROIcS2DIgNL5GzFfbdw80kzWnHLKC5uUKx/EF2FGh
oiGJswPesUaZJzWh6J+5C+kKHW/lj2jrelvR5qHB/X/Mf0AHkGOr6wDWE7oArpxu
XDEfD5M5YsamI7OH9i4KCgix0P6MUmBoBBULtjBqVgMqpmRdy4GmbGH/BWBjMT0q
FYZXNbVeyTYSYba7wPNEMd0o2JXT/p6KvMXdP1STPguAoDyWN14OBq+fCZQO550i
j4Fh/HyHcSz5PrqjprxnV8gfZ8WT/rK/K7euL1eHGyVGhqGg4aFlXgRlp1c6L0QO
7BSVtScgnJruyRTj3yojwKoZVk6nf2ksMrdmYETQo/oOByM82m0wi/8UWoXiZnHt
Al7J3pK0z8xhhrSJMSWGj8Zv16LCm7Hgvu9Zw0gd858RF8dfi5yZU0IctswbiGNL
ph7R1Q11zFXx/uwcj8n9wByQM7y3NctBFYKkx6rCmnp6KqZZEkhdqJKYvIBaOOLy
WPcq/xPlmKCjDkhkgk9MaaZO04xenC4p2QQ6H0hP89AtoD+B1/pyBx4aGuC31slm
+MfilC9nnuF2SVOxn6ChxAQMXypxqonvApm6SYJ/e8RsXDAXXq4YyBsXz0ehMsft
94tTI4j1bhTYA3JtkXwwng7Bf89BJNnDLc5Ei7ssAEp7zfx4Wh0ShAGTy2kVlL/D
w0u4dQ8o5z28Gg1wuiAMEhPBMvmi+Kv1I/smrdF+KprxitQv2u/IcyOwT7hTbILa
sy6K1ZEt7T1Zpu8BiMNPCJD8dLbZaylCqcK10nr4rDJihFzn4qjh6VEcdtvXo9V2
Vqv4s3IeOOYkU5LnvRMXnhunr1Wo1VmlVBcSpE4Ebz46tvO6ZZsQvd+5GAVJIsC2
uEnkpAY5Kjl3s8n15dC2CssMlzZRUkJ1atngcDvXCOxd8FFxIXo7zMSXi6i8Y1TD
FDATtADTEny0NZV83/IVHY2T0DTb4jWE2qyIfAANPVQCDz0tFVWSgF2rmhQEsIdc
vb0/yo7fXkRsdy369F/u4J5YXppjh8VNQWmPdFrgP6lSxyZlhLRQm6zoZzIzuzf8
76F78tfXMUAQbDWQM0YOdOmh82ZdoynVIlg/gXKVPOwyiBfwMSTz/s9Ld96mqpRh
rai1UQnzKr7xWii4nuxD/B+UsDd3hQrzCESXd0cUhMBufBUvaRCNbs3lQasWy9wI
k7AKph74C0J3PFymcIxaWbUw3qTCJHCLizjvn+fKMmWBHIA5HzuhCVkluPh2iaDT
Z6SxaB07R1pxX/vbK9Puj93Yx/zTXmEoQSGuusMwuoj7EIYrk3M3W06Z1ijTZyBo
AutNzSc13I7koITxE+CZaa/rE7rYvMz+Qt12Sz4wykJpS1SSh8XQQUW184UWBU6n
mVkOSPOtt8yZoxlrFPTokLHfTZDM/Xgwv8eE6QEooKZdDwHssN6fRicmpKJenxZF
65IxCinG1RnsPA/0TN3OASeIGyAElawhPU6q3tU4NkFs0bNmpPWER7bIqilw7OCx
SxB2q22NwI/NziIKJWaUhQ68fN8m38KkEq67TSjgXP0w+XdE2rPo4MHggFhrE9CW
caqz2JZaDTndTSWLVw3tS7ANdBzm1NSl0HaNMBIJ+rtlzDv8DBvYeB1Tzsli9s/S
T4BHY38DO9nmigdJKaBI7nh7DLlzQlmFShO/p2DMVujbTkLzImy6sOAz35EDqveS
50pcFCEQDXjMyJy5AvjG4/USBn5jSnyk9JDulXEUoP1+5zAf3dQ7DBNOCU24aGIF
hRJOJm6M9QUCa4qd6NvjsQigCN+xK0CXgQrK9ToAxjeIJowiaMmLec0SRc0zBg7p
OTP+bsdm6ukEzPwixYHov5cxAfaJnpzDEDpfo+69tirgM7Jvaot8f2q6cXGFJz/K
HgIIWMNQg+MpOlAnrdAjcA/Ih+A5Go/dnFJhFRng40KD7vdP1U5BoeZUwTV67c9Y
rJA27/o88R/DDAFm1L4XcCt5KHPJ2xlx7LTzygvYdxdlh1T0zowDAt6TT3Eiv1gV
6Vd/8VEKDgOufJRRLuIhOL0DJD07Uj9Y2A46XtAyeBCmxKn1kBGmT9yvXJDqwNr2
TQSQ9qZe1LhFlwZkhZKDtfgaRXZh0KhmTPXhZouRPq609HU9MvGM12DZ5dzCo4Dv
EpRAZnSD7RW/3JBzPRaxjMzPmCq125VqOlaQ2ga+qjq0O9kXg41NiSJVZOZeAEVG
svRULSt26f75flgw4IPBJNNmM3Suxz4JlI8b7HYLi3KfPfJEpWl4M9VcgGIx4vJ8
R01n6CdtRjTLqHXVtVtk8XSrvV6JErALwVjfP1zDzd7vmXcMJV/zxV7oSPEx4eMQ
TqsU4MVOPsjfic36lXNbaQQLb5IakFhXaygP0jaOm6HjZH9eBYi+HuWjz8AFI5yk
USvYAMfGxGXft61uQ/AgjwWQ15SVXfVnlE2z433miKyKLfLBDDWBpl31fBlOjoF6
MKAhw+1RK7C/uKveKcrY3vZOPTr2fTEc6RdbQ1pXMK1VHqfmWofbpDVxIhAP2Agg
IbIc/ypMSeCl24KVRyZ89k1i3rpxN1gb3KhbXPxQluzBmpU1g1/sl32GhA4WoLAZ
0S63roFt538Is+ThbndTbQ4G91R9qFP+td5803SuLIJYb06h+JSpeDTVO/O9tMuO
twrheKygGeIYbtF07y7TZWG+y3Jo/jY3QWGP8B1K+YE5w3tD6kS6ve2YxOEIM7uJ
JfZIDSCrzjNLyuSDvgmNg8aMo0t/qRlffuSSxk+rg7L6fQdY8b1eyoBdFZoPbcZ1
oWhsky8fYKiuDvaaAIzogvCjpZxJRZsQK7vGm7q0byQZl3S9U/1ujOpEvAK5gF+l
C6dPc/5MBStgTtGMCcLn9ELZmtpBdals91xRcHLHqWOiyOXIu4hIPpT7yJWTjigf
pHmXKasdZwoXRoFNLzf4+HpxVqNlAibvrK3te28QcjhD8J9FHuDpY/qRcDqg0wG3
4J1HjHYdPGLe8rS4HQYkBhPOtzkHTBuZ8Mkps1vd1kiiFmrrzBcpIs0grcQHxoFG
23bQ0eF3WkZzlqE5UViBsS00z1hY4/725bWyplXPm+nuPAiPFc3FE/iwRisUkekX
OfReRRAGjglXhc0dPhh41mN4FsE4guTqief+rzYZHRv2OymqaAUV0rmfAt+Y0UMV
DdHrcQJUmEN3nqqlg5Rrib9pkVAI+xttvMSIhzAjrRymqz+4MYMrZ7gNsrYpOdn2
Zw+izapjlO8DeDqWBJUGpE4JJ0cWKj0/HMZmmJQwOLMNTzV8XDvi9nUgOSy4hTFw
HLV7wQnKNK8hra1jwQIGrwEu8e8Dr+ervmOMH9Swa3qsdzl4eMGg8dmS+XtGiZ/q
RP1jogUn/YdlGVOmpVoO+TNmfDXFdCJTM+ytW+rESfSpxCGh06NCJly6i3wXdERS
E8IdNsJtHmyqTryM4BVKfhLqj+DzQ9JSlQbqiaTPJb+GnU3h9SmX7We9jo7xuzYo
rxrO2qUGkkwvYtctrKYgpSVVj4L8y2Mpcd3VTHp7t47e6hIsIla5VWzYAM4/k3Pb
5Ogr3PCPFdVRYIHSHjYP3MMFo4uq11oKl/emBegH2TZQqJuIFg7THjSdg/6wReRR
cJxzbZrxfUSi+If+dhsTCfw08umJnDjHkPzV53rNIzji6o32qhrqN3zGerGTPRbR
0zb2dNdNp0JQJyg0pez50RWz7wcJFrRWoMKBkCHhe2WPppE5NL2D6pQ6svPKDJBx
pfoushJG05/wdvazri16miL7sSsrIvB2ES/bhmL/BigWzhf0xGzdht2ZmknfKOOq
b+dpma1ef6BvMTjhBrxqIWiCbGBgs/Ei89wfcxt/H7gQXc/rU87rBeJcZy98xhy3
7bcfsMte5WoGYdzE8FHdRS4arGswSB/2CAYnxP4bLhfHZXz1+eRXSg5szFvLDTkJ
619rttNeyifvR/jVBjqA5zSEK358U84V5fpTHL9BlALf+WGcxNY3kkWRAlGejLCD
XeH+IK2TlIXhN4qBdWtIi+KwYePCN08dj6FPlwa7IWGJ99htNXQqfJW+vIgYayhE
HjFMoGkSEA2efXDJib/I+26+gGrO7OEURujEYIwDGamj09ycp5seVkrwDbIVI40z
bqnpBSSDtaDuL0rOiv1qnEZ9GwHpb8ZX0ZsbztbDyUPLDpRNuRYVllzcsr1PLslZ
dcLeEY/wQklfxlLRW+ez8sXFtXqlQsUSZ1WADa/IZjbPuyP9D6PKJB+cUMmGXP7d
N4nQQhNOj0iKQT0XwIJnq96cLPYXw1IY72Um6XPve177QDDbFjBM++ApgnQArNAZ
aMIDiWAMnnC0DHo4DZV/zDqG5M1lt+DVKiIzRYtdJeY0etgVMWi55w7EQfGK/7hi
FE7r++rLqHkcnGNT8SfRwmYVrIyXDNZXJLXnmCrH330Xh5neqrDWS3zkeAWHtkAi
vHSaZ47bCBwL5d4/FiAI8jEaft2VlG/1kUocpIAYiu0gtGEF5Jja3vbO0oUqKu8/
rSbL7LUH1q+7Eo883UnngT/RGr0/kvZVwIxdB6rBB3exT4e3mgeTDy8bVaWE/j3D
f4Hwnr+kN2wv/1UH3U3Bdra8DlKh9RTj/4KJczUleRZOKhDZBp82as2GCwsGwP+M
ZfuEgHgqDRrqVvMm1HQhLae7CGXhZKkhIoMzAoQGCgfdAyLPvoQuTyn4NvccwbMa
s50LvVZ1+bB31cqh+yVpgAiUx1r8lMk2Hh7LCI+XIyVpzw84OY6VH+1Z2FMTkIfA
8FiwewTvvQ7Yoh1wQinnxh2G9pKsUYzEUpFPmpMehiTwuc96E5vyXePym1JzbxzK
K6GtBEZTGdvt+Zg5okjHcbiF4QmYjYI5CDuUP2OzditZHvH6dfEJ8aG24c2vk6GS
RjCX1BA0i8R1/+hp443G4Ucz/8gaC7yFTLrv/HsN6XX6MNNYODkBBi4khsPmzm2q
0HlueTl89lidmbKvSpJ3ITZ+A/5LEF+mi8hsM+Ww0R1bm71Sbwmy5POk7xUuJJwe
7DEntFuy5CavGICG8CNgfFr1EYH4DWIXa+ChaeoiLOxhkIiuLGFu70i4WyaUYbME
TWJtCHAMTBKAwTeLqMraVxIYdI/gcUqMbvFbxqZwSqmwofkhYWZeH/AEJDybjNsX
ha6qgrn+da/qre5IJsHOqET2aE+ohjgYt+rjiFlpTvXl+7f5PyY6CQrpKKHnUktY
pbgI1aZe6k6zHMDFDroBqyu+ACAsK4ATH9fecj6QqUIaHn1gSQSE1PA+MTx6Ltdj
W8cu35p3peR8W0kKrOkxz3Ikl8OU1MTue3lwN0K0LH5CuGkkYTjc7LA6LZyh/lxm
8YUe6w0EqGzqn1z3t6wBNXXjQqaqsjbjxgja7HwElNdAcwvup9HIWLKMMk7CIUbu
CyohFywzW5ERZsUKIsoK97fE8AS8QHOwAzQg391E8jz76qLm2mPXj7TMwIF8yuCO
MONch+me9Oh33EqZI4pucTtlmalrOovq3x/newiLzdRdYxoF0KeaE039iKNtrYFU
MLhhPmNh6Gws2Q1ifIWu+YxT9BIBnXhjWIL5uSox5KSdakSFkfdeuRShCrvrBGeF
+VW/X96IyFPGuG7YtLqf8W4jyM4cFxzgSLmuXAepJfQ5oiTkyJi/ct30k6l6he0J
P4TTIKL6lKgOeAMbpWN6Us4oHAD/SFGwMVUrWnXkzAJl8U4J87CwatvsWcvcp+Jd
pQ1t3MarjoO2HzfYuJ1S3MlWVC11j3h+/k7LPgN3U/ISAJdsMGiF43pGORrlIS1n
T2hhhznfCyy0XVFa8PH+l9Ek5DnwtECtwupUkCY5RJ8FiMifYEFqRJ/h8IF5upIi
LSVZd+TbHZpvT2xcMFv72A/pLfZl62dk5NbYJUC/9mhePSMliUcFFmhuekKK6+7n
9jRQ2XN8CSNGSfl3CdJM0ZjtBzJEtPnRnRvQ4quvFYUC5fk+TdsW9+wImed1xfF7
SzW88YZ8rAFp7UBw4CIG/iLYXKoid1bPBgV8rvlrtCRFTTW54H/aomCfLY8IM52h
jdkZ0eoOwXk2HfcDYqBGligN8N4vn5RfLwozf+wH0+QL+lRNBbHYGtVi5XYAC8SW
tC3IaAXW5kcMyHfTx0OKHEcMU9bn4g+O5hjfYdr/+qugsqFO8sRKcn9lmAo0CbCL
n+pmFhVYVQ/vL+O1pyBcGM9stO/ybkuCCL0vD05GM85LKWg75pgBN9repRR6vEdl
t+MfLJvthnaiV1jhgiiptkQ4htXyyPMZWnAn8UHyjAF/klb/fTP95hug4zJCF3hT
hK7x4l72WSAZ7LYwH5nTTIkUggliZvuzajm1l2fFCSH7IAQjwKj1tmhe1jHxGAye
RqlcR2ACz7w6pfxc5srvig3xvBeEiJw+T1GU9rc2umPfEVhH/Gu16aO5Y5bpWLNq
I9yIv4W2wi7arBPRHKEp1LmaB4PxRV1aX9aweC0Y9l148M3RGYc/xycE689dwLEk
W//x3S9EiSCjfIMNEqjIwhJ9AD3oLfVwW57J4F2MBvDAPRRVAhIf48d8QWwNCYT/
Dnk3s2Tj0Y2KsdRcpmQo3moptzw4WlW+QQ8WIfChpTeO8D3Z4RCf8Bi3yB6DON62
C91+8KTGLfJT3d+DC9209RQXE4CDwTL07A3lyH7KwJLxqY0iAN5FgUc/pyKO/ngc
O7Qc8BiJI2YyN3umRwYFaWLxuxfV/X+f0gJ95TlGRMv9WbmUT79U4pze4rjHRfaq
Xzp5fhBjVc9MgrZEbKjDW5mIeL3bMCDOxL5iUliXJwu+frsFRHNAREZPqZqVNhPY
RB5mx52BZYXutjnG2k+cL8+MdRINevAH/dQKYePEdJhq95uHRqEgwKza/T78Uy6H
aCkpLe6riDvNIMHm0K/1JzuTzvfUFKas8X8TCSC0hFlu8pwvblpjVVgyIRuZhEbX
b5q/dGNHmKUP9X8kDajr8Sl9GEzvPxkeIE4aSBLshG3UYE3ZSwqE2uZq6VjuZxIB
dyoLdRfV9HFmKofHBaue3g15s7Ll/iG/YIviwdN6M73dOA6l5vzseacvMBmxkauu
dfUG7cNXCkkdStiHLIZ5lA++di6bHfO55eL6LbR8zta0Gt5SPaLVNn0CTiab4pN1
QC/87AeUFfRMpMaNVTGAvz09Z7B04C9DPpVJLHtmVZGGdBF54bb7Wve8y+ZC6o45
E6F+S5YeTY7CVYIdgvepwL/bIB9O6vgBdxxtsyxWja2FidP9mRu6rCxIPZ+0MtnN
mruHsBuXFdh++UgOmsyIRi6WPr+2b1h6qWulc+wxCOkfWMJz8Ry9JdDq6fFFBL6D
GNyvw+5lzOqILBmymlKXbceZH7OskdoY4qSJMlEPHQGIq++hG3yxbyA1+hRpMUVm
oXh/P62eCopIggs24DPIaCUHfHKyG2+RwCjzj3cMr+OU6CH7sf8r9+wwtjaPcQW3
rqq9VmvivZyyMxaVBOIm7vUX9+cuJH+UrCeEgDmJAaI2SQMB/pIMgXt+q0rJK4UY
TnDzlUjUArJdmlO8Tj5tL2pO+5ihjrI3gSUYrmzfJk4gw5l3qpa5c37zvQt5X05f
5RLHVXeeQTl0EaNVqVcZ8MmNJtRQE0+opZDZHJLjJw4sCMr7KPTdRGdzq/UeITcH
XPFgIqGM+V2iH8L4Zoz33MMz4guRb+Ccg9sYTRaXh0ywcaPgvCcigMAGrVFVINzp
>>>>>>> main
`protect end_protected