`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36368 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
a4neElH2SodzYSxeJ5dQUo+X/z0wtiTXizGgXCYrISbIgmQyiZTSaYaA1SSEbI/m
tsKGVKrUUFHs/RVjjAh45euL41CvUz2mLS5b5h4KGsDn21toi2/+CWoH+LWZy4mK
ajJ/SCkglzuYIcJ8Y+6Lg+BXzBi9LwdIx/tyYk5y6vNMX6KcXxLn9UaqxD5njKn6
FyNohp7Q1Xtr+nRRRzNXj5zJ2sCSfpUhC/FU6bLNY1LEWzJePG/ymOdBLCijpmeD
hekQ5zGl4GUy9QXXJnyq58wd13cMFiUXUQP6W35SPQv6+tq2nEqi4+rXIAAkL7ZA
reaIDC7i80Fakgvcndk+PhWlYEYYWywd9w8T8D23FJaS3ZSUAhBMPHJrP1QAigOx
LxeT0glzGs78e64JE3A6R70dnGy9YM+BcytO1cBoFyCTSp+oRuKppKG+ECNf+S/V
+3eBgV2ssN7+DqBMeNV9F2gx0I7QTauvsg11QoswMrKANyRIR48Al7ywKuVHJxkH
viobKiacXBNbMtUlQ15cUkg9dq6wkeU5iOe5KPfXMzQ+t6n6yylu/qXk/WQHvfcP
j0xr3YX4qrErPLKbe5bRTyRwEmoi8NFbB4tWpgzACu0wqH1PdfTfCDQtG3vbSHQJ
+QBaCpelV/b0VqohkkUUzhm5tQX7llmukh1cD1+AlzwzKzIW0NpRJt5kVMM2KSES
z3J1W9k/BhEtpXaX5G3KUPBdLmz18+X4jRVpbgDg//0InF6F01GEIG/FHV7giBFe
SfG1XwWW0//zl9mer5+Shsc6TSYH9e/GNL/L/fVDjPBSvJdBtn3WGtSAqfYrdnu4
uJ++mT8kgV1x7r/RLS7oHF+Qxj7/nizKzxolTX+XiL+mU6a8daY0LrRvcFCZfZeG
VnZWfCgqe1XZ3xAwZ5Wg3n7qhlpal06KowC8OJD6+CDi84y8eYwoHQZeNTIceNp9
WhKOLEsoYSgbdXBIsPgprceocixz9+PncWUiz4F+/PoMer8v2mVXJsizY+k6fQD/
H/OO2Z3vLfvjRVt9q15A3zm3M0edo1zbeQA1fwiSepDgwUwkGbCO6qGX197fmmYr
KmVcZHYRtvwh2Egc8DKH5v6sSG4V5xIAkQsaRTjLyo5noxT9Sg3Ms4wEqzv2MHPv
zMQh7WnOetRROuCKXfa+qtsZ3nTud4oHa/0Vfgdj/bIO9iH+jMg4EqLV4tddb0VM
VoZvOEmLc2eXAq+20nPM8OYoXbH+iQQdlS300PGZOkF121zjPAffaEANTPFP4ddS
vTQKNhkQ1kdukCp8DB+CQ8l69bbeN8mMIhQS6jjVjIx0QdeKsUQmipcstY35LHWI
LQL2WUyZQGnHaCNOMUZoNZgwe8gPwC13lPl81+bRBmLn8iwwcsv8qtTQg2vGDYFF
OeC4eS5ZetG2Ebh4KMEZiWrqRffepLqb4onzOe23fsxq59dXDJhXI7nDlzbblc8F
CUvqnAsKhNYaXGzeDM9n/QpKoD8sXIOqYzz9WsHZxHIpwDUHEVAC3hbzmmQHJ+WA
Aw5qk7XLzKsG4Fj+5s3Onf6O+P0aGZRkiY5GCIxK0gtZitr+cvPvQ3XiHSgpQJZv
8efX93JcnSPuw8cTf8jYxP5Y2I+jXq/AKJ95jU1BrfKGgu8Bj8xeUhe/b30SThbv
ozrjoB19cMqILSxLoSefe03Jc+NyGQE6s9TfhOPKrnkvvVvVP6FnZ00XIwWHR8l7
XkDAUr3ed26ycYhBXg9tp1xlNUraUcWIjGOGMThVqsmhEwhFERmJnHjdvgSKNDHR
WdzdKBcFlJIgYhRwyNNa2RAd/qRewf3R3g1fea+qioLmt+naMPlteCFF1jmEqSya
KDHvQ2paRDrvok4md8VfCBQMiYKAry/euSeGKDGt2np34R6t6Qr5oTly2l1SItKg
dSk08Vhzz5DV4Ta8seHmjNOtCZK6H63nWlZCLr6PyaoKcTVX6Mp8xs+gHilyuXS8
SnxjVvG0G/8IGMOHJAPCtJq7KdQnrjcckngHPc4A93AenQGRGaHlUeBh/DxjOMH1
ZXM7+0na7cQ3htJzeiYvwf2qjZmZUVm19acMhbI7GWYs4dZq2LRSNTTdFeQ4B0Lt
N+F2P9qBHMttWksq5ZScfjSOrJrzmvqPhTGCfpOBFaZ6M8NbQTPxoeOMGA187UEL
7/T/Dg41yiZ2SNg3SdVScb1DyFW3AXYrEqcBW/vJXokhHKw4RyijebEt7dQ9gvZH
ypIbVJkzWhEO7cJcU103tlJuxOXfLDsc/eJIR51y/+ogpbWhmPNrXGVqeI46bgJC
yzUaGfD891VkFT8UdM0DJj4+OZ1Ttldg4BFUSx5F7V1RY0FGoBOs6PeUQK+npgdg
F6xjdLwGUHeiXN5OK+PBOFeffIyg4BlXw3ZbcgUWeu27ikTw0nEdH0Ct9xUfFS5O
jr4+u7Wc2wSJRQ0FbabXndxzYzt/oC44ossbW+10E1WojPGncpPUWSKf8tYaAt/m
Fj+j+dBz/oIa5eLzuFnWuHSkt7uJfAgYz6CaiDlei+NS+tLP8eDDb3Ms9LPDS8bU
5RgF5WjArwAKFgCgh4iMmlWt5RzHttvC8fU7as3AYCs4T6oNKP3KCpsFJ2wZR/V2
PhQVAkJOuaLF+nVxe00GM+ufloULytVGii8JDbaZhvU58n/3mE4XJyXxdYIHjhhU
mISbfj22P2XhDOO//Lk8XDRb0qCc+Eyz8bAXZvhJKdrvzgOWZb393atvVLjxIX4v
LZPnKogMS2oz/UnqmSku2saUyvEWnR0BP48Tf/vmfuKg3fAkO5ywluYZ8epfgUXd
qVJFLTF2aFv278pPeYSn6W3mdD3Uv/nAOnIqEVm0ZXn4lGuZdH8qvtt04oPj13Cb
ugaMQhAwM+xaMc+gZlJQiPu/TjnL5s8iukTPlz8aHjPP+ICqCV68XuSMy9YylRp5
xw/jJjUb34izaYPXIsCQfuV0z/nLxvb9yb1mOfAyCtcoTg6EA8Cllyf1TU13Ez+g
uDdbKrL5AUupsCWNK0GtHGZlEscn6styZYAkRXb+ZcHOjCPlmVvjS3j2OuaGeN/h
2F2Btlt3d1+HBN2A1lkCplxY5hj4tx/Jpn1AMwocy65yGYDIsPULXktQ9W+KPSN4
s5x9jdJN7QazZ7MbNcPb2JR/rc/uYCjvv/RQybhlEZhADl30BWOlN9IXjBtOXwwo
QBaV3RL4eBYzI7iKc13o0QQRvzYKWKXXvmCizhJUsnIyBdInXnE7bGJw+7BNumB/
95kCD3aTMA6LG+C0FKh2JT0eN9cYLwMku526QzSP1WuUpy0LEO1Rj5K3lepbEOGc
JpbJNjJOpnyMSng6uBZ9CdG0ykBp/HU9Mj+TwAG4hU8AXHv0QuBjCr+gAnPT/GVi
3JdeN3VPEdt4xBSGHDOogVilKqpqs8100aO/22KO0v3+jHuyoDijDpWpKMY/54l5
BrVRFhSyvFr9pSJnwm28dF4d8dY+oS/jUKid4BIo6Tn55sh15q6eWP5fddt5eQO7
DAvjdfol5niTccWiNKpRHDvg52jsdzX15E2dA8uIdIQlVqG0fslFlYOxyrLfmido
kYweq549VtgnxQrfyENsEY8IS/5vmVDoLB9M4BIOIcOQRpnaXSEa1PuKfWvBPeAv
XY7Yzgvsl4grRRmjNafj5fXT7Dk1H6HoHu10iR8rpBSsv1hlchgP4MR5107WGLgX
nWUEZB+L8ewP2EvtKJqMoTmivFlyxO3iYNbN9nqW2NaBbOtG5t4FUCc1dgw694ZL
83rhjVGdYPM4pn829Gx7QEuaR4XfHlCf3GTkwP5LEyWGjKtDBL/rZboRGkNXrGdj
l0cBEm4xHr2Wu+Gj9+cxDWNq1hzk6z0VR+Ym5amcoqgdda8oKjUhck80W4YgVHpZ
GyzuQk8+vTpL4viBPCniEKVZvIXsTu/jxLllYZuMoARaRH2naktx4dFk6oduTEyT
J3VMeAZzagnq/3pif2cMM9VEcyZVIB+gpmmJ/j45bD+LMnyxneJ8PUPtYoIFb7Gx
uuONh503fvJiHHML1h04uh5iLDUCpzlatoLtgrT+B3c0kPoRnkH0j0F3nongA6dl
3Jb9lyXyBVxalrU4JyUAEUNgdfzbe9Y5Ncm9+M6iROrfvaM5lQyKkriaHkNzmHOm
4P2s2OjFIwC9iHJTH0aljnlK2ip7boZayVI3J7e/RZCQuwank0Z0Un/TG//VGx/p
87Ws7dv2cgthe4qQyqIRRDlV9IjtvkiOHC838tLpoR+MX/jfY/nQ+//LukyyDXPD
e9QP3YT1sfXZ/9YilRsJOjym7MVezXAlOJnjLyjtaP7mnXp5hsQtKj+CGl+RWeHj
RYsT/iWQRcyOjoXr7PM6zZcYw7N99jUIQayiFIzLakId/WzJOF5c4VzdB4LxDC88
JmqDeuxJXf9SgnVANZBI8UduPxXYXS/PgDq8YHrx9KO9CRfy3RTXelZp4dCGAHPT
ESY9STn7S7Z9O/VXi6c3kwd5dbMLXOreuiqXVA14LR2keuIM3xQr3REnyZY2YZc7
j5uuJ1CloovcBGNsg6/952YkDmYacoKGDzAQ12izlJpSXN1ZeoPjBaWiqaoPtbh9
NoE92bkhpYiKBuPtig789+liaLXSzYq7cy6Ga3xc+prBpKVjljt0WpLNwYbtr8Ze
BskO3aQHGrR6DVLTQdTUVbCpCmlrJlGOEdrT3obEhpPVZF7FAtfom7YeTRYAivUB
M5XnZHaQ/P301UBM88okZUeeXkvoniUSdD24hpnIFPouyIO8chsRGJwEafGpg9U9
QH2tt+o4OaIQXlhPxWJQLCjIwLPwGcCDrga9BKR/uS5V1vA3HzZO1fDK5Oh3uBfy
wkXnpsLru26CWV5Ej3Zfoxaz62PiOFWIR10/6kfSBJUbaUp5vx9dcuQKP0inFIYi
apPBw56UHpUXk024gm/f0f4ysYuFsy3ZsA2Shi6hjZCe/aHfJz1YvuEaboBfRFxv
hX94VCJQh/yIWCHXMcvS8bq2wgSvGdWFRIgB99eZx3CcjFbdFdzX+OfmxPP356Da
jn/4/xnni4uScR2u+I1TgEDIe5IEyASzAR6e4HusGiFL+PQbFpKTxVPcHubknBJP
q+Vngfrck/RUxu2idouzNC0A/HyQQtRSD+vN0l54NR6a8QiVyQQ5JawrV0rDay4O
+rephrkaAdkIZADVkAud2BL85ND3tciiNb0q7uso19NoFCZOaIFtJeoMUyOKThyX
exSmZ3Ec5/hFNhyQsBijCkQWn9RSEfcIt6p7dojGdx02THEe0A0hwF/sBLjckIB8
N0vMPIrPv3cbxr4XsOAYqoarcTPBcdtgI58aUoSmEdXG+HbZREAKnuUKQ302Vt3b
2iNDWHJO3zRJFCdYxEzo5q3A250qpVpdJRAYk8EJ1Xg0BsR5OraphCgsFSfi4Itv
YYRO5fyhAf+SzN1wEWCpcRhHAvTKsfrUfePUxF7nzKep2fw0wJLG6MjOPSDgcR/O
r+YFz9964CeedR6y0ARweYi4P7y83LVYgyvyFLRARP+Yiz5C3uc0d+8jSnnxZpoa
Y2vDvaIQZygligiUqvJ/uuMQVGJon1CKhdvm5sVgTC9+onn3eSLFGbvNlV9AhQSB
c0Bf1SAcRugTFqYb1YVPEZ01KQx+w7qEz55QL/y232bw/NTcHHvAJzXyjPxMYPIF
6OV0raGbCW6rKM74mOgh28D8H2E+OJ8kqy/axfLYo4TNoS/KFe9ovqftctwEyicZ
tpXLK2PIxfdJSzpb2mOHZx7RV1A1Liq8zo0IAHMZ/x24HLbYzEbTmNVsSwNyP4RE
yOVIYKv2M6pZU3lcYAooBnAs1WxBFF8DCFMEJ8MibtXfrq8C9pb6J7DP69Irqjo0
L3m3c1++2BtMW+ufk2yMXisvDBHEe50OEFX8t6wNg8s9KlxXfwqNIbwGVtJbl2KF
zEjSd8P6lXS78KpfY9v5vk4Q44+2DLbKhgrIV8r5eiIyYxG6DBgJ+s55AnqPzKdd
hxcQYaVfY/L2GLpuoZabvh9E8QCYuqAnSVv260CtT/qD6rAWssi7bpr2cp0UqdSA
D3oESaCU/gtqJTK53pvAK0Np7XPPCGm1+OK6jMVbkkI5jPtQCILDCGpsJfP+mPJp
d+kJVYNu0cm4esaxJJO8DseDRbvhS5bCqGVuSYskEAcrFQ2BdgQZ5Jn1NtvbFzzy
FDYJ4Eoru4ppA8OUXHWWZ4KMQdIu1zbMdshAdPh26AYL96DXUtMYYa1EHgd6QLOQ
cHWn8zluiQIa7O7ERgiy2s2FMpWd6s/3QLOEBHenvH1mWxAHzHvtd5V6Fc350f1u
XuAhIFdS9MY5QZAgXN3qRZyRyEXQtCLC1WJ0yzEf5NGz7RfUxRTkBPhbU6ngqATL
+X6nJw3pj4JeoPLFPLlOgxoT3unFLq4sd1WFrgZFkjfqLQZvtNtBHT7COiY1wB3C
X6d3Sa0ehVArIASUv+I5ZVyXCkKGb3ivg+Buhp/RbnX5Xe7f5C8j1r6SsthwacbN
9Vd7jHUdcwgKI/sLbs10rh1+cPoQWuJ9SB9ENmO8EeTNEuwkdsEFCgDjqsGhbbW4
UBbBbL6HCP5K5tc4lTVQrlmTnpq6FSGnRJi5igSYMGCRyNMVKi3Nk5cD2OBEexLj
/VsJAs6IuYUbtu4S80EP/JalTfu1DxFMPvyKD0m0K5f4mFfZNpGBiGQ8B8VQBy1X
6CioeToIqUv715dVMW9htBaOlyPOSLeHp1xGXUEVRUbjJgt7Ndg/dzaHJiPmdt/+
VYCHUWr+J4Z9yF5BODMgtuxi8nsJ0WLNYKWouHJNPmhZXmNW45O68q5uCCFq9moC
1d6+g3IXN5Sp8sUJHsowvmNbX2rTaMBnZvPytJ4ko67NizjERT7seUhGeBOu8NG/
H9wOZ/4vjtfPz9o1JGLXcU2aPc81wMij6oE4PyGXtvDKRcNSoKn5H0nb68ANWQlc
by4dn/OHEp4G6gzktmkCs2OiQKk5DJZ2zIh+CTWm9vjaeFnLrtYvUZgCLGVwwYOm
FXkS8hFKKIv1hCGeSL215yug84RXfhJ0LZT8FKH+h0ncJ4KDyTirRy8A+bDBDYRR
VsFjV5s5ZpOXmCNmZPTlvfJYA0FSOuqan/Qh5COZjh+R0EzRXB1m/Jm1j5dcrH/9
03ep/qQak/QJO2E3mj7CgPa41ibtr8EDHsHuyw01w81XWIuRP+2KRwTVgud02uwg
AWvLXMXTGWFtZuL8dHpbAindgCXKeDbWktYk3ebivHfZm68lBnzUTzuD+ApEkvz2
TyusQ8PMGDfocdNW7toowBq0fnx6C1QsyA/TKqUbzlz2AvpJzWAzDryd3R0wg4uT
qC+UQEESvp/nlJpMMzPZZeXL+zXJ+7EM2RWAYwlHUiutq9+hckCaRZjc8C/sz9A1
HWhnDFVM55f5saenxR45vt+KZbtu5c1ImA1H0UY8MIGnIAtdmbqD9i3KCuNPdhnr
PXrvelOcNzmoTlchPWXLvz6STlaBja1MZGWJYHv1D3mWiQeniGjB2j86EQDP783a
GaTbsXffFAEX7y36707FSQZV11hEvacLqI3kiiUmMctj2ee+stXmqyc6+P30UE0J
VIzgNFxNxqQFsqjJa5C/UdwuKH6q48uYI/lIbocK01Ha6kAQuVIinbO7a18ErEUx
mCtDI18H6jvEMuXnEXOgR1sw77yzPmp4LRedWvlZcYlojQWMXw8WkpDNHP2+NHD2
T9mVt7Rss2xqIj3omYUiDwY4K/lLD2TfErmOt5Ir5sxM1LmGGrSq2MfSyH0BYSOr
hYv5y2F9IDn0oK4/2doRjH1NqV1dVe+afGvEGp/js+L1/YDewlf4Y7s/rK6AJ801
uMxSNQ27F4tZuEVc+br3Hk39fJZTpF8C37/5/RLedfFKh27xfjRWlk0xXXwpBRU0
Py4+1//N029PDZ1d/lVQ0ntU4xmoFKLq1JUSvqSoH65TTcwNeo8Fq24SxPdWXL3T
Py1GPJixo3zFpZlxP08ei6kjA+vAPDPKbBpazJeI+0L0y7PNh0m0WfjKIwrn/Vkd
OLzJSBqibnzIpw7KXvB4u5RzZY7wjz9KarYzcDQbkWeYMrD/Eu35bM3faDnrFRBc
wmcJ0TtJVIpsRbAdsfRH8lT6Y3ArpKwxfSkTCxnOa+aOClSh+v+R6BgjN4R0xcYO
Oz6u2xP6D+H/JRUEVpSizAeOjV0LdRQMEAwJh0ig9VB/7QkFB6XaYRsjresNKbp1
SK2jbDCr47Yg1+UIZIJ0eZqkspSEiPp0yQ31rcQcQGdsrR6vQr+TNcqpqCX4hTgU
ZZKp1n+9JYbdCV+vz+UBWXS48dS1YXuodGunan8OAyLlHw34SpCkPyqpCji1a0hX
KvbGV1KV5+0gklUkB7gOJ13mA6G9UGygM9kjD2nJTB+fTIlGEkWTtVMoWnnjUf9D
2gg8XsslRRG09Q2pp5gzP8duDMzSmf2iYW3hUWAYkHzK7DehJwzGUVeAJlhV9FG6
vzOi/Ac3QwpDyMiUQXt+XL3QOLW6qe0P8p6K7KrSSbC2DoS6uwQGkKDpaDtnO9M5
2o17i/Jg4YAO8+B082KbtnQpMd/FCC3C+/eslMrO2yaDnCRi89DuaOCpd21DVF25
gebsoOTCCzwXlYcKT+PLpalx9NsmTIrqgCr/zjODJWah3TFoK2FJR4oiT8loQWKF
kGplH9TKYfr4mgYBGmUiOoickn55MserQdM5U84aNYNZigUJ02xDG4VtaBi65uAz
7Kbw5u4+CFFapPSCIB0Afx0FV+rc/Z/oskf72CRCnwsLMaxzpQxdeSKBAa9r0FrT
fwtp85LrU1v0Ab7Tgs0Dw854kYHPXmzVHoqbkRKHVxrPYP1Vw3sYJa4pK1tOVS4F
5570SlmB82TMIisjvDShL4EBh3HMtHdwhBkEKo0sEzJChe5/+JmgEG84NF8thKzT
pcsCMIPUexJ+A7gYIDSNpLe147A8RPGQY/Bfszoz7X8+R8PJ/xvQK58hb14rl/pJ
daQoPeOjDzmICZ/KpogPJGufBSKD1ozU8elq6/EH6G9whOsEonoyqEHcFm1iNchS
2BTkjnY5QIjcZker9r0UnmJGL7sg222PLQvtCQiN7/sBN5LvPqzMs6CkdLeVrODu
wQGp4ehY2aFlMIqYZwAL8rk24GHbn6kTCcyNuQ9ZqShEkYjj/999iCyHCqgTaWNe
AXyGpRTE0mgS1NyMBkdiuI2pDOoPWkxkM+ZQEeMm0O8ZOKeAbjlRUqPja3jvDU19
4/+73S7HGCr4YnkoPKEgqtD65WtBoRUBASwHn4PUUrslGtNUMgHU3UXmn/mTebo+
dGqbXGE+2Sg8Lm+qGce1QBFgX8Xa4eIW5l8xjmDrYb6oXSCCw0Qi2gwWPkrCJkXq
W3UHeNImoIuWfA8Kl2JKPQ0+fXxXmYVMk/GT/wuefFmoN+rCYSlOTFHAjb3+vmxM
QdPCOi3Qur+4dmcxufkYTBXaJECmoVxqTMXqU/PL+Xrk8V7PUQB0tNdhl0c5Us7q
cpprDs38PIFZw84FyYVu4RKHCzPF8jTqB4K5MzauGkmF6TM+kPM85+g44bG8kPLk
XqqRBjzntZ9VVWqZKurjdH/YmfHVNyNZ75ihhovqLQwz/6kPr6QkiUSnbU18lq8R
Fetd9fdXfByF5iIBi0ociVxeliWogGkNITB8ulY/lZ/PDP1uNASQXgwdzL9hPBGH
MtVnnVXtGTmPB6k0vdGvp3g4HXmDmJCT0zEQzZwv7p30NnNUPRmNcDT5LOBiiu8W
hL8Na5fkJyfzDV97BhEJ54ird7miUdiiZE1sioT2DoU2GsGxqaJDkF1UVaxscOEr
psm5DEZoJ/U94imA0JLaHuaLPz9HmM8KkayldT7GlHtja/PSADeYxBW09UyeUjX1
P4lYMUsm+wVlndWd/F6latjgl59V9MHtWdrvt2NukLZxkp+1TZJiCKYz+VEtkANX
kMMOKDrLWNXbi34EpXY1wEhYfT5OXYLo8AoY0t5uyj9UmQjokTDph0ekRjkpgF5s
NQZBG4EpRKmj56DTGyuOjBk1E+i98VQbaU4dP2o2nuhAJiHJEwkc1yTGDqVRdxCd
vmGy7v+lJAzFFcoyxhl+X0ULZ6QkNdxgywMXbKdtk0HecC4RudpvBeZbLK+qgst6
11LDQdauRNxKzmqaXNlcJOHSTWRkJ1bHrvdLTDFXtNVPWtNYhB+IDqlNJ2jtPb9q
uTxaJbH7clXlJa/tYzBMGyHOKETBE1BSZlPZJwnkCTXbgxxC6g0/3xeQVPtF0oPW
8SbW9OIQBAsmcUxhrKfRfGb0DqT2AiGZuIdhO+xJ4g5TsYcDlwzp6o9cBU4jwM4c
t2YU5dCu97pi92b8nXDznn3b95ALxqjGKqTn/JmVvkizNQfxY8Uo0cjtqk2wVQid
5a+HtV55tI2va7fw0VTc4ASa2s1Sq8hYdiijoqGsruivP3Mw/STm4/rKOWi78Hah
gG7hSLPmrVgmICDDYvtzPZDSZerCElH/3G5YM+/k1aup0EMRGIa8ePEYH4u85K4A
qn3fEGa4/ZykgDQhBwdTph5TfZ9TJngw5QIu1fUTyL6vHLGWRa5L2AMN99azBUO3
rGLQvQghLEMQ6HhJrwkPIa0jeBOVn+rXBhhb/bJn91q7UJ7GES0DUS3C7LwqzjTs
htiND3gzQKmBfME6IeKYfFW01LisrnqbJAtek67dye8s8h0EZFz/egGYlhOIdBqW
SVYrio/VaQyKVGeB+m4uGEOAhp72u+bSEUloRwRe2ZRzptk+6FK/H58qpS0g7a9H
yBZTT5br3PhR/huZwFB39ULoF/hcqCuSuNi0ZkcxE0+8zR7RK31aeMAMVltnlFBt
XjK/OWl38qY4gXXYvQpOzbmsvKc+a1kUpKtad1uEbJR1nPLUA5cGcnlQ0/RNqw0D
NJBVSk1vfomUsimzaVfE3yzdk6SiuHp373BYamzxwCMr3jppQPQynVIvafgGbD8M
fKpt5vyvYIcYtBW0jQap1OzrRprA3O8MXLg8PfAKFXbzErCXFHdx1yncZgES1NaH
6LZRNrTnJLMvVbd5UVAo+IcBUvcUDCth5OdpfYGLRITEtC1vj2VWdJgPFrsT4rfp
3TGSjkaXpUliafX5676On65wsMygMZ0BsAtT0wO9OTS9OaSHqPevnlrH2sbge3Nk
kHBYNLCL8p/mS4mMfWrJccb70sj5ht36eXt5MYNPzDB6KSEbYdcrcDuHJMz4w+qg
VWKValxSE1QzjQT6oQnwvAoIrhmLA5nVc/IFk+gOissuFlhTumG4UiXah3A284kX
1khdZzJ8s4RjntZkbXDDB064vwqlyI/Kdr5h4/auHBLcYcNC+QpHra+dU5Uk+Rk0
bqN51bE6cjmCGprOH2sKM8tO3DNO/0dFrGv8RjKmtxQrdHZtZUpWF+mAM/AhpnxC
gU4gC+JhPWivgWqblwjSHt83QNHI/5rEhffUUaqJ8dpSjFu98cJ8P489l8+sFvYj
tSXOkH3H+si6fgBUnzOYLfBtyU9sBTLTXpIc8WvEV7y3sWI89I5sG3OI+R3tfkk0
k5cTsbSKanS5W+uZ9Sl7hmx4NZ92e1b1H9+/kQgdEt+GmwMpjNycwYvhqPDRzFaZ
0auRc2Nxgm2cQlOyE4Z7DazzXqjsDcVRvUsj0JmF/Pw99Bw8z6/XckcWxrH4eeHh
XNwzDGMtE6mYvYZHZSEs+squgOg3ipXohML8g6HKfdtrDObkzP9vVjv7mXoxflKg
HxGgVIDJWME4YpStcUBbnRYLQ1BmWA1TvALmgjZeL3iJAldbdAoLFJZnB4bs9qoR
9BDO+agTei4fGJFjt0zZlbFJyw5nJxMgjsgSfnxBv6A4soba38IvTgRznNB9pk/B
cFBmaaIfZDkI9DBdMCUyeE2N1oHZLn7eYvQUQV7ip4fL2UNKNvk5lQtXufN3SICX
8v/QEDZH0FeRts46yg7gguezpfxmCsmCZgCSKuQaoJzs4LJGG7k7SeiAnxeJwZBP
/zjQD31oBOCTgjbFHY1YmuPMBBa0whxq9jijtFyHmhDWR5yCzdRQaZEBk9SSF2uM
qZtKZZRUY+h/nV7vjEnFT/eP0AADbv+Spo418A3iouheq2esFYwU6aip/CwmWHlj
TCExS6EFoO4hYr21OPvXIOJPciGPAvtHqBwqFqZ8pRvUKoGzPyi6sbpzuWQe8Udr
X+7WaqvtAkkwXdSpFnyOxnrJJnC2J/mdMuqYY5tufN/V5RgIgeaygIjOKX4EuFnW
1w1/LTx6xZjDlTZS0eNRLfS68dbWFgbfRC0FiHqeR3kJtJ5neyvLLU0irisFTxtV
DKXrCuh9Lulk8P2Pmf30K+IAriINyOk5Yyr+yvwJsNhTf2gQ8mBzQv5zRp82tRCq
6p22m1IU/n4MurL9HzlT2OESKTqbHT6dOtNzrpGno7jYP85/kgEig72xuMJmYlOn
bJdbTxl0CEa7lJpGMYFyAt3f+h1jYCVPFYw2uMJGBiPPl+1JJBpL5IGIYBS856Ez
EtCDXSY6DFbTwfUmUkH4fH6EMb+bJE0qTYgsPole3Fu0Wj0yI84qvZB6zhXRWRCE
TKZx6A+Bs/9rh99fIWaaxH9jpaeVrJjYs45EjWgqx66OJvscj5zuHurBLsXVcJVR
payWiJKwU09E+aH3rbSAIXTLVlkyaJT+HLHi+DuE9mMO93/Sl8Ntz5GcKWc6TGkn
OGOa0Ad/BZLAUlZa6AXRbuagFBJoJ6krcEdxy5y3HBNERCO+TT51Iprzfs4jhZ9r
aNpfppG5s3RBUco8UB5/gJiDSdtmczEKvAKLFlZc3RGGANnyM17yBmPkBLd2RPpF
WrRbhpGy/hKx1TBzANu6IgKMYj+qOe4YE73oVmAYjxT35fdfWqrAC33JEEzo7GIK
xqcn5CJ/kPiwl50IV9rh08ytWgcgOLNi53gas6FotOGCamiO4WxFwWLwrwQyRpWW
yobEFMqAITSxVOxNZdZZZO7UcU4cOY7NmpvCCOuOEYuxUp2kcwfnOc+jRfTCAwXQ
VGrAeD7FDqiT1RXCdpARtG27jkdd2JZY/KE8nX8iCKptLix+9o20cyGkOIXfTNw3
kQ5jgj/PC/+h36CvfnELWFnsyyj6gyFc2z9P60m4CtqNQpLYZPA1j1XQDZrPCSvY
67MrKBJQhd6McKj8K22mHf9eUI+89k3esHRTP3IaQudeK0Z4sIrAbcXJGrEyFCzX
WgLSmd0AmeGdR4o6bzYSc+VWkZSMRc46aIdCgjli5nM/0GpQdmAV6TuRk5ZqF15R
cpjBZFpmx014mo+VJ18fG8vfoF5+V32CNjkBd+i41lZWAGt9LOr4F9HTHb7wnIAG
HCgiURBKGHHs05lLEyaRND159E4msbf5qJUxDkU5qiFyscDzh/FrxLaYw9/JY2jV
crHgRzD9N3TxfLeg2w+uOcYiEMG2fdQQ+azVe5GqNWiKDI/svquZXuQi59lWqRh9
zAtBuOtnTwV2hb5SPFtStXPBytIWP758lmh7VYEPnESURAeKzEqzAmuLvOc5tg4t
qRz0C8zCKSVycii2mTUznkRgb7Zmyor0c+0uZ/OdyHb+Tc3G4fbuJaR3nOXQ4Qt3
AhhkzEJPUIeBb+i0juFWobCZESupnoCajyNr27ebCRUyAcY3KM29PZ5lX5Jv/tkM
dIEpv5XIZfHm1SGQkhUkBP2mjg1/fyFngGeXc40FM7mkvzi4aFuZ7izHN9S9Ob1F
78pNs0cqQX1DpqAN5MwZve0RW1KWnAYhUmNbwBgKG8p8sxmyjsjGFjOQ3TYlpS/C
GPkWovDdaJgEn5IDZb+Q4Zn7PFCJwz+FnQassRWCVyoqmS7SrwV9iht9u+GyDIPa
AqDi8ixDknnqppXHPkoLbshqthNAkm5iCoaDEpjLdE/OFbdhbFlZvZnZTFVh/wcb
akZUMaXECv+uaE/gGGxfWbAc6Meq+zWaFT+hj0YZoFE581N12710GhlScmeyNDlt
nU5OXK1kzSiD3CLV5O3eQAiJ8qcaL98+VDnflYc9AJAUKbFP4uErE2Mk3o9ox16m
yWHGRAEG1ir2x4jFisaVUorF3tytIgeEKP4WieuWC2LN09b4e6WGc/w59z0kWKJx
U8QD9OvtJMYtwJhavvmQ/emU1o4nRb0q0QKSB6R3vc5IC+Or6b4A2WTT4i7iHPE9
AbkSUBF1a4OkO+w9K1Vo4vMQjCnTX4NtZQ4dby1FQ+7BSZ/obc7mFKPckE4ffAvg
s4MLxeysQbP7tCMXoXB37rekJV8hxxzUwqgZnr+0NwsFGZI8wVImEVXgiDjnsvYq
Y9uoAqRnic36kMJaHkl0ZWfEl4Lo/XJqkpJbbTlt8iu+mnhdOcUk66Q4fNKXhN/N
wKYOvSxWANDIIPOkjsSwvrjoe2pyWui0GATCw9ZZTpOyymKzMC8H+BuEGog+wjy+
n7VHL77alm7odTxfQMU6Qddx+0QQ22Pn6FMppMoIwBVsiv2Prbx6j3HBzzmJvLbx
tUj3zJ+fm+ugUO30KYZSyzI5wNbD/zf2f8+xVB4iU073sFzLra7uqCyKEokScZiJ
r/93TGii6e0zqXrK/y7LY+aM79ohWUnZb8RY0F6/oRuq7i4Jkc6Ux657J3WDCIjQ
pAwhd/BqQgUGSZ5Njb3gw9zzpFD/5R+xSOtFnS+W0Q7AuuwkWdUrlHNem8Y5e3RE
gVFja/IU7gLJNxx5JB7c4RPGwoGGhaUoFVX7IjB703xkuIHFtvF/n0CaOaav8gBm
z7m2Mhe/S0qUZi1GioSVLUDVY1qIIe9XL01Aw4V09azwDdSGdmHSmUTaOUPX1OCh
+c61UQTMimj/u43KT1zV6P9XXa1lCKz6fqVWTCZf+tctzegnMDYtewZL3UrpK3PI
4UZvIbuuk+30UIG6LPK2VSDXtQUsuKjB5ux0v0Jh+TKRqDsSWgZlup+aJfk9CoqD
9uiZrOHUCTcPPFCENPxC0sF0Xn0h6jZc5OPJbOgNzYaR8PullgVi0h+BAcbKDzM7
XTZmlvzMr6rm3kJWIjbQq/ATuJNpNfD7jAt8beF00OVbKEMwI0D+38YJEiT3a20t
1chYtLihR3yxY5DHd50eUqPZHEM0LlH8TSNAbAyFy35Lx0m6lvWJOVHW6d3BduL7
DeLhI6kF4nCy4ZPFhlVf2j8+WUwFTEc8BdYeh9UQ7UQH+UHr3dhkhrZ1F20fXl3b
x990O47hKniotRVXrjwIfeu/Gt695scSg3LsFBGorjpYWUEKV7bm1XMeMFf43OMA
O4DfdhvNVxFOIRzqQXQj1I98wArxxnyRa7gBB2hJCNQmu5FNxTlewBiuvM98gNdx
nUBugv10fDfmfSwkVKTTELdXrprksjSbDVSeamKUTvlmyu+sZrjNnOVF/9sausHP
2TlwplSxYwiWlRPCsPFsq5HVu7G8oqY44yHAl4OgKqebd2vSen4wUb8Hq8AuZQSM
FTmIayTy+ntiE8mQm2MW/ldy5IcwBqTY/qzOrzO7esHNUII6j4nvBjOGaYWnLg9P
RfvE9ReQEZud3memxVBJr8/j1TRryERcu2I6uEKsixZUxFdNMc4qBmhdBrYNL+cB
AZ4hWjGkPz7GjhuvW8Euoo0np+J9RkCi/9RhOKAI8XAHgZP+TpS1CkvNaRfjh20M
WV1ZaQYDq3HXq9BCJc5L+1q6wmPruV+2XWRQucdXL60ARhiDOuKDVCHEeS//YEdR
Ix3RX+DZPDG7uKI9WlU689FYlCNHzTD64a1kLVTGxv0E+nzqm2jO33sDrA8x0EiL
gwBq7ETBoxVcsfrjoekxVboATzgMMZPuV/vsdgcSmfArcEbIyfRWNCNxxrMhyD2s
OhgUKJAuMsqa7mbPK9mVJ2HUL1SxNmsWNxh/nNyWMVJ7932ux+iPytGUug+U62By
O0zV4qmzUNKUp4Yd/dkxQEFzox4ixemJFKB6XD+cKEs79fKluaVjT/QoCFcm9/xz
9eqKWfGLYVARVg+5M7cprIIf+kUfCczq9PLgNQgSaBOQqGHKOVgI3Qo6g9tF8wco
+YIJlYT0wvC2F3E5+4g15fOGhP2Qb2qa/l0UzDR/O7jTvaVG6C7GNhGmvLbAt2lN
FCAkZgTji8nZq99nuwBrRNCToM+K819Ukd2UECPre0Xgo6P48fv2k9WdrTqLkLoh
kxjoBEf+wTk4v548dnLGFiqazUsZ9IuRfEK2hrjKcOdVZbLXaAxJJ0wufWsLhAri
NU++KxP3aJZJI8XGKNs29yjqKtFj0uPM35juKOzCuLtjl+sFb1xstEZbw4poj+Me
omCfGGOwkmTXohnpYV5hjFmm96NcR0BuLNgdQtfTMzEE3KkG7xqO1YqRfyyx5Acv
r+Um09phQYTM1Yui6H9B5jP5xQkM2RDeew1RPT3EYkARPkhM/VYLESfDg9PKwf4/
xjBZne2c5YeFrqPtwaUyjqR5aJPsZsNfDjvPnYWtgbRHha1zQzEoKgfjlHXHYcuO
3aHXMcQrEPkGwamcwoz+/h4v1ApCYc+B+cWOzLU4qO4zEtQKjNj4zc6R6sS2Wfra
KbWjHS1NZmJ2NPcVwxokpCNbb5qzr1hFkWg+S6hE7gHkkFNEH8pmKhTOY/Tbjdfo
80+LQn3auhncgoSnIm83NprpXkPrd3MXmcPgE1nWpw9ZGJBCNhDyGizn30lAA2fG
6PzgoTlArLuF1+LyR6EcA3oS74xDTU4LCjS1+NoQIPSgTEi0nBzkVTM2sH1av3ps
ePo1hZG5gpMMQMHVjou6FvPoTjfWzoDlZwk4xlkPd/gW6976q8HKx51/91nrl7mZ
kUQkG4OpRztSFw18eZpReu1F5uxV/askOp+W8FvjVePb2ngJYJjEcSDRAbY2Iwcy
rop0LMR8RmeTY2JHqoOmf9n0DkYu/94h4eyt7vDhFGYvd8aLP5Cd+LL3+5G+qSst
1DdU2xO+C8+nNPJKH6504qPrXYszfagy1h0McYWdl3b5S+8YfZgSc3G5gNk/eC8F
L2Su2j8cmWTf0zFVgsx3qonIqbP1OFqxO5QkGs1czA+qekZztFUfOKLVP6vyhV+c
tGUGucvKhsd0t9JfABPhzPsaa2XhBx4nekgIaJY4Vi8bgQVwIlALSRcuNofjJ5XT
K1dj2Mv6aAsrWzkMR7+KeArcj605hc05bJGYQMyKQVK1oDbGeLLnYaSmScooqCw0
5E8bZHfP9CP3t2M/ROoCNPb0EY4BY2ENUIot+Ncub1MzYn+RLFqCx8NKBXmN1TiL
aPSbwKix7uPtkICaV4OONnxsLzEcb58/xRIdsrU86L0jKyh6z7hO8OjnlWg7DwS+
a9rR93f8rjZcD5ubf2ckN+0OJ03riE/bBaUxV9Kx9IEgqUM7ukueWXQCL2XrghDw
tUZEBgHh6sEcX1SRlhukGvdq0jtqa3qwwaHlLc8mv5/81VTPcvlozWENC1Jrgrv8
hoejtgyWpgsXC6GWC3Q10YyZHHTnQj+nBeMmBBoX4e7pfJms+poQc2TCGIuATu0P
hkeGM9buaEKWho96wHVAdmzJE/0oGQdl7rse4+xOpsIVo7mMkD1NVJVxVawW+7Ie
ReFCdA2RrBcrYa7Lq7ZbmPScHt5N/pHYFgXkaozyIGbNeY4Zqw+mDLqei3V7nPnC
lKj15mkWPb/9WJsGjZMd0ZoDFgwwPiC9D3Ol1hSSRlsAhtZkPPDyyNu3XwfJLnGz
ilygKhAB66YzwpAdRFAKGXrDPd1wizyF5WR49N9qgl7JC/6rOe0IP5GYP7G+9eq1
RFu7UYPbBwuN+F2VhNKw2KPcNIJiLNqu3UG3bhvkNr+pJGg6cxq8vwGWBgnBQ1Px
RYttvfH/Ug5BUO8tb4Cdvj0nTfaw6CUtMs0IPfB3EjvYdruZ4PcP9+V/xqnQFXKB
YKzoEnseDIFRg3pQVvWfCBvWPNXc+omMXkVXO5U2qLfnhtTxWdInv6pTAriz7Tr3
MUYrK5e4xDtIyOcMM9hoo2sco4BIMdfHQ1QUBy56chFJhmkyDceCaM0CpOG2yREz
hvolvxVfX9XLur7f89gCUlvJ04NniVxVqRGr1UKSRcCUsVdQTZ84RRFpC72iUSEP
pN7XM6jIcBBFQj9znrV+BgzUSzHSafwleDCMbWA2jkk6U+v45Q5j1RH07ECTyeEW
9jdrbPQt5mUtE6KlwmfYrnK6mU6YHXVgQYtWbJfeOwdvg7K0j3+xtz1XOCq9HuqY
PY+8P1k4H4XlySbk8hgUGVHYP5yAJZJX1tOnd1D7c1p2cnabIRpYSXuLj8+Ga75U
JXjxrhGEyQYo+760wThjKHxXwLryT4umlddGarhqiQK+AKljRNDqbUcIsKebbt75
nBXgsJ7bEtcf9O1y0jPg0fGrAre7tLMdwOUW2skS9Imcd4XmvK1Haof10FsY/QmV
KKALfaXQZxp3tApD6bmMJBiQRptbcbu12U7tLsr9l1Vkaktol5axUXxOojnmVDft
XKrAsR8Ic59v+JHRl04rUdgGRim7EI8CEmJn5gdeknuBzt1x2NuxlGW8s91CLNeW
PPPPlVUmj/UiFi7CJFJN8v4rH+AE6mpomCDwVzNzajZFif2se3dAk9SleVa4l0eu
CgsVsHgBKluxiKIA+EF+/CuMeV/Fla+Y1Dq0BkwA55HIXLUk4V6kfofgBKfYDW6A
PgXnFzNmywbvdga7wEZZXrh4O6jdV9EOaj+bxHExCALHFC1GGMnOXpkF0si5ZKaK
2UJl0+7S7aNYEUr/ML9x0wwfyDE3QH+NRmb9Fiwra8RdIGRcsXaK7rF6Eu6Xwi1I
a14GoqXOx7P5C1YTulycihiKST17TOi4SYGYrEIzPjLhedkaEYFW3ykocaJXNZiy
X4bkG5NJF83ZwRigQZqIWjm/3aHDVOgzDL7HltCpJjaMUhpSlcrzsacyuioyPWZE
dCRQHDxm1FIUoMQAjtoVqLQ2TmeWPhJchNbDTNWjhPzK8Cz4palzDWU06P0gIPyB
wAyrwDdkwODCH7Pnmdbj6WPzdvEqT0AcZGKF0M/RcHH3QBOM0HhydKgtHmbIC9Pr
Q1zbXWRKshN6CzPS02ivtbIeHuz4hQ5kpfq7PQap/Lh7kwTKs/KnQ76UiBwK+cDj
EoqsBKCvGVXLiBDqQKUtpQf0DCi9dELj7kAs/xAN//1rmvFRDvn1V6ZV9qWb4h83
QAoDQdKX4eH45EFLNtJTlvO0AEK2pAmsfaOGOy17v6GHuHYej4tmetVn497bp1U6
AP2QUTPMqe8jDthIyr5z5+P0f0NiRM2wJLjm230Sjb27+ABrXnpYBaDfHbVdpWsr
8KTYDZqd4PolxO2qQ+jBY4OHBFRq8Nmtdu8cCUFO88OWjtaKzhUZCFuZYDEX0iBV
ty4xkdnZZ355UxDKqd4nSNuv/6xhxwOcDSgGPEZCY1nAryYHQtyCAaS8c5jx5naO
U4XAssfj8lgvU5dtQcJI8wD2xoB6sklKVGlJfsdDNrgMV9vzpE//Z+fk/MhNGXpN
6p4pYVN1xm7z/FJtabvtuBR9o7cuMX+o+UHopqpLv3mC4y2WvOyt+Op2w8q9xBRY
66VdkuDjslffXCCRv+6JhjMQHjhEG82y0SjZMX/fKgIkLQ79rNON+grBY+r29lRE
Cjs8IRjfPFdPqN6ac9NANMfIrb+aUzpIgL6QNTZQW7ySo25CojPadjDo7piVKoC5
IkuT1QLJE0Xhb9GZsTQdFa9QtXBeeUENVV365O/M0pkODV4XYdqo8YEbIZ5286GK
fgbLcq++Htq2LEksyVVpSriAIOjjWwgMf2oIOB3D/jWj3RM5aR5KlHuavM3n30Aw
h4ifuxo1ZjDPfwRPi+4nOf2TWmJ9BZ44ZiWr6GHGoaY+/GsMkcmgsmaIJJs2E8HR
4OZrboLkHnMl3Pmgfo/oIjkQfOYQniLCX+o0YgwrH0JYTT3oFY7GU42GFX304d+W
PjegEtFW7BW1GHvE3Z3i/tXQAmm/QTkRjoyBfeF6PJk0EztcCLpWuGr74jln8Mpe
ncIJ/Lu662/zJLVTgK4bPd3kmx5VSLWoDLzcB3eZ/UFMFGjRav+Hd06g6GKl2nNe
4iRDn1Ae1mHW12HT5pk3EucEO5C+8ia/ws+JkilwYXUYP29YaJVkuDBHH9zUSduj
7HERBQEi4nJpvhRYWkyLyi0nSZawqijNqR2FSKRQrv3A22h17OTSKertWuoX2tFb
5iyzXjUdczl289HXalnCIPFjvZq5ufojgQc8RAs9i2Z4y9AGtir4Enwo0iCc7Bhl
gKaq52jSU7+bvKJWStTgbeIEdJNUHbqab10zydIJZE+P4qEm29U87V3TSuJ9Mzg2
v8nwohEx9IrAvYPDTxFlNDos3QZNJAc1HHV5DJJK0/YyPibZFSjVc83QzOEXUhRy
09sitZ75Cw+4+aaQ/OANaRjjKxieqYC8vP7VNUdLF2zsNekK8IMwfFIEqL85Nl5J
xCRdjoWr6CKizUXPffXdQ/1MyGqpLS7vZYvOQCyckINRo5aV3BYTHESe1bwJNjaw
i1AjKJXy+O62Is1xMb2JInZv4Etfi5Q+si/Gp/e88oG1Thyme4PyVdnERIPVgYfo
LDj+bhzhaXCVJ3v830uVwNSe7zf7fxVUhqnOr3sySQi6ZSGArS/Sx6oXsitEmnPy
7kvMYkUkT7DTj2DC06M89YFNdtoCMgR5DPqO36DAszQalIPe6qLCiHmSpoYemx2B
CGGcyqmQudgFGYzJ2V5tWZp+9tUZkTjHLUnsBBB6UWKV6pCdWoIhkyq/wp3DCFIJ
LMSIsWG1nlDtmJxojIItVv4Fg6hMgJzqTrjX5cgGcgg+dy6j2saeEhh+nHapNXy4
rDSLJInt9Sgo1lXUyTqtlLywoVCzhHhPOh99N3vz3Xn0ohLmyUsqLe5oCayB6Px3
aFS5gRj73EKtdT+D4Cb0t2nXF5UrOPfVzh8tIENgl/VPWbI7IRbYGumlIfj49YqH
bjp4KOJ3XFryaCWo19f4zFCxKoY5lQSNKNPvVse+tnCpznbzFvZDDrOVQeNDVKOX
7ppsdvfY87BjbTjdR4szBlMLjbpkJUBXtbjMK9JirLcgStrPcHvDOrZNtothehUQ
eKvQIWlNApdtFwI4YR8Qk2XYCUyxCYKrphcyC8d78PMQalujvTDt3tEZ7FJWkm6z
r4++7+M8ClvpcWLbyfWJKJr9N9Dlx1FjACRuIp7XU4rD3YrG3DgRg5bKCEA15NMi
DFQOofst42CIPsrnVAPu4hXaDfnOF0+smUNLFCJrfMea+XWSMvBOcqGx5jfD3cIG
JOk56rch6iqNWecUQg4CxH75A7/ETN3x/AUALjH1OwFv0okpkjwbfsWA5Y30V1uK
qTF32v4ET0xef2vLVASBLIbBy4DXX5WLqvuF4PY92T9jzV1fdYxKrWvT3JXiN0PM
o/xafBrn9+VCdqXFNdFZ2lNZNpD2l50N+EvgSDBhYYKrpHoD8YqKVHXp6M6xiKd/
igA48SpySoI/z3HkJqj+YG4XjpjSjf4Zp0dY4svOoJf08BYyg9xIqSog116O/Z3w
lSXFXIebp/bKRXGtUZOJBPeV9V5i6YvKYCI+BsB6KRIp+MB2MxKljgAgBXuMCeyJ
RTDgomONoP6REEPWoBWyAezn+YvLs31iGWPD2Q3wW2bWBNvyENtnGF/T3oipKHxv
xfHRuTTTbbUGLHPc2PAhlPpTmH8ywmjebDz0R6hQnp7/Ilcd5oD0qIshJ7aFxsvp
G5f6NCmbzeLeJeSW7sDyzKIbpgX7pYMW4oZVDN2Xt6KYwAAKOwZLHskNNhynOOdG
QQ3F6oS0eKfd461TlWCS4y6b4/VtaNoFtPZ9uOk3tL8jrEDc63R8ozUiOUsuXSBd
HP3hmRcNGJM7rdXKlri+bGMQSpJjZbVmAH2bcF6/iDA//2xj0qKZ7IjUtLJZ9Wnr
V1hSKlxKUqLa5Lsddmk4i0hY+JtTBDm/MmRjU9zSn0fh1c4pP4DiQ4YOq/bqGgo3
cnyNgSXF3rgYn/ODQTuGQwc3ATh43zK9zgx399OLMm+egSvCYOIQNKuyPqaQitr0
ecjieYacI0caZk+YZ6mHyvW3Eo3McxUZVGYJDvrmu2ft9i0UA8ThmXgCKaPfs6D4
Y/7USlr3NVX5sj6GX5TUCfYLGeaVqQEsGwN0TEQWqIsbkxA9fkNP3eMADNyz1kwR
+Pqf2364b2AiKHEB4zqealAyuLTI6BTT4iyyAGkCT8vMSPbNC2OkpWWsvxUnSeFE
Q/Fv7p1fO7TpNHwVf670CQZ6ivOW4aO0PJbBlCvTDJGhOSTxCYrc834pAtNYQvH+
WBsT/23gXuWUFoDJnaz3UCAxpVQupbZvkxXteQgm0qpD3AbKKNeI3eyEDiLLOAC7
te1vlReSyOATLNRNUuy4Hx8XdqYyngHU+6Ph4xQpwjh6TYgxjl7JR7PbIjYYB2Fh
/YKrJMbgr2AY60Jd8H6cLb4Pzg9FTuQiNVJ+KIswHAYdWMpygEVJgBqeDYrKmlR9
4VU3SnbbpHo5XVpJg5j+FymOdjxcNKM10KMsOw2w+/f1kcFCCIWpCBA7vT27Ktyh
XPaVOUfcC/KQxzNUyfKKARbIvPhuYM8II5ODcZOAAvSnb7Uphy1MnrIFvJja7xnQ
4Lxj3Iku2HYHlM8umt7pmOtqSi5kpVjI8edlcB32BrJNjPxxdoH944eYTcovb5j2
7w0BJMWWr5RTZ/dSN556jho7qRt+CYgn7ePkPhCrp/fPwimGilXup2GTlPYZlaLp
fTKnM2/Bk575VGH4vTClmMNapkjEHtyaiSQQtGUkg1s5nPLS1F+xRweAuCuxhaSj
ZWpdx+5CQ79zwDxupFV5EKT5x0D0H6BQ+UWdHcCKS8E0K+9MFrsr/eTJbm4lkeY/
r6BnZMyzFwIJHERc7nE3W5kz3zoHHF/LNpcZGqhfw1ajSk5bFP5iGut6Xwgn3dDy
XgSOdWS6ADhT2uv77EzM0jDOqaQOWueUwCmbZyEde2Zgs20mU8ggf9L3K8CPO4Qc
PRHz+ulzIOQHeP93Q+z2viCck9dQSuAgkHYcRw3hq/VfHpl712B0+LDY7b+nM5Ix
bX4F15v0jau3o/vkD0W5UGWnB7hWL3s/z+aa1cjlmvbhLQxVMVOHkKh2Oer5K3G7
cjO/sjghp2OwVNxpBS+XUUG3A4zqzIrbCEjMpv1z+tWTDDRIOWpVN+Qwy+J1oi+o
Y9bRltq/5vJEQvNfCraGzhhAHE+AgO4bEAFZYLI2Vk8WCHyKsiYOgxqctHR5YOYh
S3ooP7G72pVhzNbyDASX38t8CU5hnjn+x1nOGzTCVOlBb3vLGCIVYbtouk0Lp6YJ
XKjeCMoYxgjs1FpGsSZJF4K1yqVD1XBPHEyX3d5wHgixFO9bIC2Dpkk2bjVVF6bR
6Zs4DHES5ITcYI9d72X11htZqAk7fatwTosPiYVAm4VDRtRl5shMC8o/9XrWL02L
MTJnUQz+vY9gkHw/LmXCVgzB1FbpOKxh5a60czBxGq06U2zGD1EtUCNNAOTror/g
ZUAxGSObcp9I/JxgKuFLSLxmP1YUikyf9OYSHatr9MMLuZhI80Ahn7JWpOrlJrpf
5IXS7nsXDw7vEtV4WurOd9n7HooUQjEG20EUfC22Ec2ONO4C61/DfZuMXkEqB7iR
58bx4C9fsoOKI/OYHn+aQ7DwlLwOOt8PT3GlgYNUE0DWdAjqXQFk4z0dIdmXuzQ6
oBlfYCl37CPELmcaz1cBkpS24/MVwz/y+SXgB5ju1x/k+Q2E728PkVdv8WdzGISz
tXN/tOksfUY7Qe1+q2LBrrohfc6ya1PX4F7eeunp3JO5ZrGqvq++gGrDnF1uRKKE
476TgBbHUBHH3333H9ZLVPlSHIxwk4hAsaa3c+tn5y6XXLue29lJPZF0noH+rmKP
jWX9BiTJflsfNiWV7anVVkaNm1j8eURIXU58boUF0x1I7w4g6Z0aykK9q8Ya403W
Uly1tPXNSnJtaTCLaOnNLBuZXsYebEq+VtY0xOfSMBiNwSaWPk/TryGRv3COIYEY
cGnvvLjccz08VB3lN3MuW2HOsukr+IJ4HRQqI0lrtrXcfWcCvYOs8lqs0H32XcIL
dvivipkdRl30WoVMorsXGBBRhKEk1j7ZD1ylSpLvh2wEElYkT56jwSSUNySHrosj
Gi3jp2sYamW5N2ninlx6yguSCmFQI+rh+rzXxEqu44ywKB4WiCkGm+rD/0vl99Lo
u/WZn/6oxtjdvvcEjDKULmOqtvMKz7kmdudgTxSAFe9sP+jxVKhSouIrllsbK1Vo
KctIiFkfBYyKUFLYq5xkIHRcVpkOjBSglQHqVD5hAVEQuqwMsxO01FICxq1wN0an
RcBYDcvItoVV3doFa9imRg55sSu4+9m7BUneZZXMNO4wTEf/was7PCJsXo64GnSr
L5MaZ1kV6GCRUPqQl2v/IBBjWSwFF+P1/lEdhHhG5V1xBXgCKCQspc+ON7YRguKz
ra7NoqBcVD4StF5JSq64jQWUR07g8VXQhGceL/zZiOq92Gm+AGHBcIeLYkE+wbKw
ZaEzXumqWLpcwygFiN/e3pAibICa3/J3VUNKaYUH7tWeIeJP0ZAo392N5K6rVBZl
zyiHMGoDPIXR4Wxal8G8pa/0YICLA813PQk9wcz3UhTgaLrT7Rieq8chxRPBXUEX
+NZHsJAou6L1YeNKkvnja4E82ulYWOzRmkxIvMpJ+l1S27D0UFUjvPyTk1InE9yD
bTdsHK8+jRJMwCzxUCWLC0d/SifoIEYuhsLoG8aW8HMlBCBjDLGvKFr7zsDCW6aS
//Ib3dWRdi9tTLMXD8Z80DHp7G5QIxS0nafvbJoQypF70DhGbvEwi15eT0KxIy2J
JomuZQDS4gQSGXhimIRp8XN08n82xEE0sOdPbcvbXYA4IHgFdETE5GaVXTgShMV6
wTeMOidgNwUWi4VQhTULhLwhL5U/yAYFUlKxz7K0BxBFGwb5EN5JCekhgRnExjqu
H3ZCXM5TnhE063Xqb/9L0XF2yTVn1mzVsxJx0kz1AnN76Mo54CCsATutPWl8cHoX
h/o4mwtJdhOz93tJupeevmsXUK39tOlQtfPTctZQ05Tkk72AnA9J5rWGFvXiU13u
EGfINasBKDEGLJz0qcqWTYxbjP63zTk8uH9JjuWfwVP6HUtUl2Wys3xGc3pDeS8A
w2FzO+yfNrA1A636rRCYiDbGQ5JFM5I7sytbcmmRvCiyjSBX3jNHXoa89aI8pI18
XkRiu0dDg0fDyI29WIQavFIzWdQoVaw+y/2Iu+vlhFa7c2y/LqM5J0OX2k22zGJU
3GlaUABrX0prIFrNrPJyKldh+V46k7+Z4oB1IVwTQ95tHplMarnyzmiZXNRgKd+/
8m96lz1PPn7XyzWsafF1ct+YXNjb/5aOEgEsiqjEyZcu2NbmTJFsRNgW/c7z3FDM
Qy+4TLKBlePad6G4NM6WKaE32HU6ojUB5YWDLlgZDlunzeNaOre2t3vzsRHZfunL
Ltf+NrxDweWTRjnevdjnhn7+dyNnff8VoXpYQaFJNXujieGLL8oZvMbTCKrdeFvb
cFVwkuaLPimijb514S88JwdMdumxE4c074BBCwEjYFvRbqjrJmaKpbnCu96P+GVH
o3qV6gxZzNOdZ63JHddWwu2gZ321vr8OZ4WiO9sq1Yn+nkNJvsSTlYaJvC1rypOG
iEgwMLSwg1FUxWNFta2VpS3e/W6zNKSDlxX3WPnooOYoHnU5iuJUJgXrJfgZ2w1p
35vnvyPdtUPIGBY90h2UBSDh96kkOnnY2FLMnj6lBodJISRv6x/+osWnqSXziGed
k9aFi+09c/3M1QQxCqMOnfe4u2vRwhasDYm+xuNdnPxemYtudlHfkvQRf8HIjFyg
QVk9yZE7dt6JS1BULNy0Ufh68ve6//ZlwNWNJ7h3AZHQlGwafCv1sjrggCLu5bGB
bE0gLtVBUrsyGiEhzO21r7eMW0BjdwhvUwcmjw+8mPSmhAkzNa9KvYqDHZ5HxLpZ
ZMeM/w/JO4neW3rHb9pgDD8yLgs8m0GCp72+lv1cZ7fWrIrpiaTxuYRVV1Y+5nrK
gJLBDQaIHu+IG2uLtHYPEu9yE0VUx6qbyi9Hwxbw+UziNKqeJ8tAzAmTOF0DA6F9
M+1nOKkG4yhKN8G7CrO84AehvA4UEEmvJzfnRaZqhLhxPRYweXRtw7cGJkggBMx5
mwCZ1Aeh1xRm6Fznjr2SaTpGp07XMvwBqxVl2IaqOZNr+8lqvCo2/3AiGX0aOe2s
OLQ55/VFXg2+MrrSQu2cPGdEKA0S+0hOlRRWf0qiEZ+lJk0NOwzMPWHWpeXlTmKl
YxjT7A35xiWDxn72Jq84ul02uuQIVTpUWCUDVVCYWjOuu4P5c+x8lL5M6JlPz9b3
JH6XMfupn8eJ6CwoJYMPMPZvsw1iwXp1rC9abtA1JRSGDsxqHqKD5YEY/K8TA/Ud
9SO49IoWzVsw+Lzn3wGRPKjJXfImbNjWvfRNomyxN0W3DoCDrTQ0T8c7/B6YMR1P
3gdc5h0+yhovMFZCHy45DmdgwRElskczoJOrmF/JF/6Rn12+aUB3uWJV9VpR2JbM
UmtnOJTUWzebX7cnPdkRosCHEL9dw8e0Wj2lHBsTGFmD9NYoYF+3HSCTXwjNjXCU
J62AhBj0D6atzqWgNeJIJgq6TBfsxiO+r034JdfO57B2DcfdPNJZjzb47bgO3NE1
mDKahIeAh1t86H7TPXgk6UUaM6iOT84jfxk95h6qoGCveVcWF23Zy4dwmeFyN/SR
d9xmDHS1KkHPIsiV0px/d+juRPLkDwabL00orJBP4kcsJ6TWhHrJjNdO/YhtrOa+
36M+pKIQzV/64nSPB1NpiR0BMYNVL05RmV0ZTs+bAYGMgVkRFQDRByXnVG18u3Gn
OLdWGU6pjk7xLizSSRvrJe0XZ3beQ+DBdndKQKZni9Q5qY3Cko3d3fMvzSXnBlfT
8JnBziDthqIvG/2DlJgOp+INA+9kD5iBEO6cjxVFm0J3MBvfT/L4QgM5mXMGcpK3
3j6uJ4xxUz+D8IWUSj3B8qcvE0jdq4LYXfMBYyjOInj8ugfVPPt2WyhQxxTjLWrq
MwW5Ex1dGu+3ogUQw70xMaG+iAvmOAeufQchfzW7OXFnyGZL4hhUUS0F0YGOLqWT
3uokJHPTFwg1C8nc9RYCclyJYo/6o+QmYuH1RgoyWDZHal4grUwAjPevgUgp7ajY
oO3ULdvXgVFBhiwvU4q5FNVejKM7qUJrYlkkWLaJgQwDGOZFrFs2pYHwHHr7Kuhn
ZxEHqlQ/Od/XCXXOjnukvQXWkWY7fk5hyksaiL/aNMyA/ZWHflc4/1XE4Qi9yBq/
OvzKHfWyNRjEDLLp0elPskd6TRWMwB3DnmnzWhS+YaegejkI3mLNt2s0KTrrq5/T
KzBsmSGGSGZkx4hKDxf3YZ2IE7y7KuVuxG57qXoo9x/+f7MLyzIRcCeA5pRiIcvO
3bHoxPZbJPNAsgK6IwilPawZm8rHT7nfdmy7M9CoqHIwculOUMseGIawBG1wxCXd
yeHaLBB6FEf/9pjoqpkV6IGP3VsIXc7wVRP09B5mbbpJlqiIvzd35hLleerT9TTP
I4PSl752bNMtiyfl/TSBXUSp+S+Pmcw0hKYGCKpxrwNFBkILcEOX9vNuuMzQleYY
n92Nk+sKncSzxHg88hMZbtxf1ezxLpbavGNcHTZfxxfzpuEvrJzk85GV/QBVBiCR
KQY8rhtJCKVwuu0/KWusOXb2+2+3YKXBHWejeJ+Uelq15MCw1TXahCbgOjNVxK6f
XzIPjluAtIeNbeGvgdGMkRaoNbcwoA/TQpYPHLO3KEbYGn8NZz+CLeYi2ZRSxcZP
Rvhhl5H42A+DX01Yn3eyy0t7ysw6+7V2NDpnNJzKziCZgPn5r0OvTabUX4JSYsRZ
7YNdfDvFOYiKOpzQlI2l30A8AQL4rIEAMekDUTUgNiIDJvaSDWSBmL2G4lOMbSCh
SNiHtJ6Nb9UQsL49VpTFVm5cqSrPflNdOK4SiRznirRHmGqoIs2ZzQvaG3NRLlYP
AldeumrceG+JpxG5BqVBvWCHciDnhc0lfWVdPqpREi8KT04IwGLakME4aX6uqd5F
dTg6U/sDBT7SDU5rdqaBq/HC9gbbK51fRWufpTvAnT9jw/kKpzDa9bbubUegbLV7
uTZWRw3Y74JEM4b1zI7sys7f8QcIPfepD9qhbEI1KQ3zw09+J8GSWiOdxcZ24CLb
Ds/jvYsgTTHUJl863irIxbP9F7ny+1PUArFn9vRAy/J1pcE0buAIHrHlUyupy1A3
iqaDOvWsdteOUmqW6a10mShWb3Ci4HeOvEN8Pw2phRA+2i6Px2Jks6oq9Vg2F220
cABEqT2Ulr/b07hlo7En3d1fFMbTvfZcjjSyGDYY1jf4whqa2kCkUrkCfYHbbexJ
ZxEu4tDDVD9lQf098tAYo+3kyYpCXVwMX3XnG/wA9sGTi8zgbaz80tQ0AZJ6/Xzi
p/Y8QsxWqeHk5DVqKqU7wJRUa8i49xZQg/Wd1G/fwfR8bQBwQFpO9OtqAkJBaghD
9rdhCkrL8zvL3RUVQ2YC8TjCdGhhsa5JhUiv/KIfzwrj5dg1Z43VJGRw/DbfP0oq
WqfPoW0A0EolywoZAv4sakUR/sc00jjnJfNOkequ7e6PpTCZGpTDnBTlvGAQSnxV
0YEaO8LWkCfuW1PiCjLCMgRtohRwTfCkuC8sPCzuMBRQL3XOKt21m+ziDQht+Gom
BE4ZQRZwRkVqHm4JIFdCn/yFJxapalZoBnidOJ9tKrVWz1vUF079j3xvyMQS9txR
7dUOv6z00yLoiwxpaRa4foiSWb+GLNk2Za15ILRCGYt2kVaw+kF084lxWbWMKyG+
FHi0Zq+q+0IYfscAyksiixwq6fmE8vKgN4p8ubnbRLYMhc23drzS4Kys99kd+zpQ
3oy72bNSmdNBGLB/5ejkMHgoygLBENl4yWAl1wmnoU052PZXnnFa1i5eMwXlsiS4
bkm+vs2je3lx9h3yet85qRwkWdQwMUf+TIBkODYPpLgN2xiyLKGSFj+h+p2MZB7W
6HvVutuU68DTsLs2z7rDA28NdNqdA/nLLK/Y0AgWOX8xVb7VkqTiWWVwPorzbpmd
6894AKs5e3fYvJRyxXvsyPydIa9Sjm1LUzr4JInLpy6zz/ab5hD+GCsJRFha6aHR
yEZ58a3egtmaz20zmBN/0FOhF36o6D1S01AzdJ2TXWe0PeWuUjxxfnRy1oiKs4mH
9tkseYNjAHP5BurQ+PyZrd59v8bSVmSPwEohEd7gBhaNOKyXx3NwiWavlphrD1QJ
6dgWOAwvNcP/eMOnjSQ2EISDaeUqVvQLeBjdzTDt608vNOjVWyCPFSMVgR7C4e5c
DpusQY6E9cd6JKyZebmtBu2TC2wRbi+mdHjiVu8YZzfwmoKw5IbFCyzRXJLoTFX4
XOeASPt45aGS29mKlbUWtejpzXz58BBILZLc7QaD1hSOPsytOzW/9Q90KVSYNlGL
WLN/LrX3uhHgc1NsljdespwtmnapI0AZxUSt0mwEJD9JBEyR+lXg1heL9S+ALfGd
vHMdbIxfwOj40nzVaMTVZaAR6q1wvt807H7mDz2mTjVMLSz3BQm+yGLV/21pJR1G
9digitDi835Ukc1vr+0F8R9W8SUqfwiADUqO9nLnsdR/joXK+aCekmSGCXA+HkHW
Q0KenVibgDKYgjO3ngmtfmNNnFmhaze4bf/vqlnuFFj/pyIBTqVc4MvU4nrtfZ+Q
8CRIWkwUU+4xmlL0GNfOjSzo0jXpA4HHy3Kw72njxOmMRE0w5yvBuE+cRD4PPizs
oDS+rjdUFlSf14/8dNvCvYDALd9TyZhN7c1pZ9xNHgXLnhr6WxlOmnwVaNWleIm9
wPbb4PBec3Pg5SPCNz0Zc+M8uOFfSlqwCESLCgPQ1BGujFavWNqfMie1M5j8ibA0
5uagUip7+b+2n7M3ImKrWXte9WM5f6HS6NY6hzXSsZRCZhN0r+2L8MwdJ7amFG5i
RcuxWKtyZIZGxug5AY3eFkI7IH9okxzCOJojmImS8FplItTsqaXM2oGEkTExpYaC
7M7PvDIxmCLKTgKC/aPzyuKPfb3B4qQBDtyCdyK9fvKJFzi4gGjbirD6p9HGl8/y
sK6feissW1Nmv15c+hbol5ZT0e5axotHFnS7KvgFZokfXJPXolv76kVhZ/hrwT0k
04ws+Wz+6Gx2CAeQJhGBsTMrUaV2N8jxYjzohPC7dpDcsqlrUFXP2lzZbc5mJBzh
HZEbBJkfUJ38MOo9GbLGAe/ZrH5/cT+N2rcAcucQ4OacOXWkKYUWESze9WKb56eB
CJZjMG17MYeCdtltZkB0J7REMawvm8AAdySyNdBIEagPyICpjMM2AY2fj+LBlE0Z
BDJ5CWhJcuDMDoqCgIL79m14TT2ofI/rBSs3PQrweQ3jXOFzAjpc78MkDN+xpeBW
29aiElTa3BwZ2Uw/lAhhd+8pe0tu7yPcDQAS0fqgWPnTEDLpZi0idbPEMmA8XpOI
X3YH5kb1DqlCMqRUPh3XETTbzZ3jMdVFuCt8bBHLXW9aHyFcmXOpZMHBDRK3trpk
Y6Xpz7oL3oHI01SzV5DrEz1J2bfgCySekm7jppU9D8VB7cD3EMnvb8IgUxK2rVMJ
UhLiMIql/RNdw4pI6N6Vk6YpmR405TLFeGqVogZdaf/WP1ZE+/Ju5EFEyZDj1zRm
c+nS6FNGv8NGgQNEOJ98Qdzedss+dLovyQBt6nBP8l4VDz/0U8pLv2+6rbQMruqR
YodOYQq/1DoENhH/Tfr+tAP3cPGoDWIOTodWeWoLdoR70s+e3U43OrnoiS37U2FE
ilLtAueoVbyoDOf2+b+2kaTs3ih5YvcQ/zXOTeNOZsJnKP9TMBHJzsyGRBOC1Lq/
vDGXJsp+FWvsReaGArTK7GZp+qKBx2SvSh3E4WL+NcmdHTF0Yu2S2iYQ56H3PdjQ
EkgBODqTluCdK6tzGuaR/GNa4oO9eHOyfeV2HvVAC771zMISYPgwy8a4V5I6hpq8
52lBamYvOdS3ymdmzRaCVFWQVAbZRUTNqfB4gSEfhfs4iyp8FpHEopi4hmBjpwGN
2jwqwFz7iLV9AV1jd8sp8gY7LEmLPFhoq8GdiWZ10HxNlUY9/XyMx7gvm3Mc3wjo
28/V+t0AR5m+wJTS9xMPjAu8u4hqCqWXVC3oLPmgs8OfWuozdf/VJyDVRkfooxKy
xHge99FYJWZonTarOn4hWS6wWRKx3W/IWe/uyJMC5o9vEVXpphj1JCNWXpPXejsX
nSvthfDg0JDVHpNjvZzcYU6e+Vji3BpvXYYZlKqr6F1mD7Dwn4pkwVzwW7/38Glx
vU+Qxy6o7VFjZIEEEgGgKYM2azR2j2lTWWfCWJboz/wuI0R7CF6Tip4q+URy6FeK
nkQZC4Q/2I79Po8C8JX64ExXXYJgM/oE3G6zNZEr6PTcFr1pWJq8ikbaxIZmoao7
vsttS+nA/hNHWKKfwOB9PhXQxD5hysVKvdZEIDEHExePMgw6DQXoH+3831+/rVOS
TvChF8d/nj7iZ1bv8j9JdSsRscpFTRktN0aXHLt2iTfbaxtKLBFIpO3kIzjuV7Pc
y1NmS/8ai4Wno5KJR2nYHiba93oh/2Bh8YgbFsn9q/+Es89T/+tCGtv7TC+DU8eE
HPBhieRyv5YpRsTI6EiPqrx9YytsbgNFvLK+UjSCYUE/yW/NXiFKZ+DiqlRJgmdE
n1PHlqyb8/0UUlfrRKAyXvxGLo0MzVdHx2FvDH9r7WvKDZn4X6pWDBm6zj3Ahe6d
a33axCkXbq9OS0Vo+ozL3PTY/udsu3rOJIN7s0GrByEKse50t/BjQbQ0hBhpr2y4
SprUt713iUF/hq6aIfrxoXkn45igOBmReo8lorkJ9QLjze89lHNTCOdPtJMPdHtE
6qj6bwLiIbrCHJ1HuryFHoLCrKhcPoSlXDbz3oh463hJOxxYyTM/ZEuhuJOW5RjY
bVeWIQ3It3k5k0JNtaEKO0h+oHTbmxOFxgHdeH1Pl3RJoUhc5jwamO1SAr3QUngA
j6c61EuXsXzsmXadkzqA7VIAcrPeZel/a20f5jDO9qtxGNW170Z3iC2V+TsuLtFj
gAXcYtSyU2vCqgc1fuW+odd1FQNklfRoxHToP01sNeSWCqLrQ4y4oidIZdK+VP4H
E/FtGk+i0wKSgmcyT5kET8wFqse1M8SQLM3ZpjqC35ZCuakPgwJ/3AFF4/3YTE72
Qhd3q3Pg3QIIpgFU/bB6OIUO0L22cbVA+SqKL8HHTAKN2yMeEMfT70ybz9LhSKys
oqjeY3apVc54YnZAi80Z6fVvka5oItSh+dmkEQhUVvcRqlyVpVLkb/rrFTLKPpYT
neWRggtM+0mPb9zHic2QD9qfcYuGoU8bBFarh0Hm5xGHRXtP7hj//oeEOpFpexkC
CoTBGguAfT/RmOfI18XU1iKNvEQTzA8fmU/3R9cc8ZplCtvmXi3vYdCrIABfRe1F
aoj0oW+1IMnACwSjPB6XrxShX5kscpWW/Q7kWfMa3hKZkQv4vZ2KVS5JTqj+8tW4
xpU16gUheuOzfW1pQaohLQWAkpKRkprklGd423xuzUTLC6As+hvnxDL2PRkQBICZ
+KTmEJqX0PSvC6qpZykHJm0EyD2owROiDh/bAWs5Fsgm7mik8U+WYAYBLorKs1ez
sx2ACvqW9vkKlo+NJ4KbnM3SE3piTCzg9XcqozpaZV60dT0CrhU5mep7IkBBNVVJ
27m4iXWXdecww637dkl5A3q99m3TjVAi3Y0LZ9RYQPhFI6ccexPSM975v97dEMZ8
FefoHXR0Cnv5xJlS1wZsYPUukyeC0FDpilgHGAyewdr1sFRXcZIoBKLXJeXzXxVZ
1v39yz1xVKHwlGo45ViEe0uZVePMHwtWkWF54r9THsgQ5fAASN0iNZyz7HX79GSq
7/Y1/zMi1dY95SPGk5K4rOcZo3yrXsMHFGLJyeqiL1vK0b19aoTMXQ2cDJXK47DT
DmqnZc4r5yZItReWIaWzBb5OAPe2G/R4K4ynLs9e2TFPm7Q3S7cjLNv0d+S8rnp5
ZIFQjzQ+BNBvHhllv1hiWLYSS/NM1wKXodc598Tn+4I8wyQUzfpqpSyJdRNuyXYy
WAeb9l1BfIBhAZ7enRZMeoRu2sZLOeLfzG8s6hLrZRnc85VWh+nUqAm9B5GYlhLg
hKrDE94NxnebdLHlfz7yLEHXvCxAa1ksWcq/8tuAL4U8iqQi64iH0aj/f7sh5zd9
RXabM+ahe2q+s7IT+18XiKxXYR3etefLP/srfAWhzgNeilymzrmBeTk+uHs6rgEL
f4txm5DTsA6fowHBxh1VsndL9R45Ywgc02re5HiaAJ3OTNQPcWclzAC4Fuv9KXzm
ze81H3QGaTyUmWqlqn0Y4VtiT+SiyJXMLZbNKssmZ5bMfuWdvtVtBd1LKBefFIaY
rLc83HO/2DjSDRhRcJoOGpqT0FwioH0AROQVnwOIyUf9wL0Z+lm1b8uoK13K/iyY
s86FPP9DDp760xuoUvnUr0vHGqXphvdqE0Cf8qTKnzUEqAebhCuBnn+JU92pbAPX
JsHpxBa6mGt54cBNCQHQyV4ulE8wgIiJeQUtaPKxe4GxSPFKnK39iHaB92b6rmnK
e0Xqg6JbYE+S8szkf9xHlXIrukwKOt/RTrgod6GxV4IhnoYsGitKLH1mSYrTx/SK
7fzBpfLS1Y6BAp1S82xLOpNGiid4yE20S5X4t/6FvxIgxTHJtwN8F2SnrxzTEg7T
ZZc1ikKQyQMBMg4R5m7MHx+fe9JYhY6AvBrOvTQf/59P8MwwOfJy7n4vafhmBoon
v9KWc/omO6glZgLaDHyBMxfwmCZ4P2iWEArp/ZNLs5zhaLn7cj8Fr9/BAC2u3MzV
wx2Dybwq6JjfOTVVr5CFL1R5BO373o/skE3z9yt30xQRQYdG3wodjLklWVu067u8
xk68K7Waj23wleWUWifpZiR9Egl1150wM/NJl8wha8msE0Xci+jSNyvVft5MScXH
XG6FNKXuUnnmuPiYR2rSQzhQJKvpWw5L14naJ64frx+TZ/Q6laePo+xyROoM/UQT
FDVIZBN5W2xQP7Ojwj6Yra2Gsl/uSCVY1RpU1+lqOZhUukMrlWT1um39nNUJAbuH
XaeYzoBmTZY/ff6cY8deJs3T9JEHxciz2DivubummUFq5xNLcX7ppPOKZ6rMPAzJ
njLfzEusnpZBR+kExAukN9NjPNBURCkfntdcJnLBZ+c+ZFL+9XuYOCy/CQBP4h30
h8/c82oEsxYP/87ArjyNyWOd7pFwElKEodfiRdq2abb1/VwgAAapZg9wPWArUctp
UrLT4tOSftIkxLy/x1RIlfj63zJEomrgfQX+XIdxtKwq2VajbSSzDO3gXSYtNGmg
okKiD0+KzQqG5jvtAl5Oicbdy3V+NoicrKg3CSGd6sSc3D1wGriYhajXlhspXEYe
Zvcle2zdOWvsSB3L7pGtzH496txJ8YIXG1IVRbsFtLDDaszaK4YFzm1mULO+GIRi
4g3h5Poz21MfpqWDFLn3u3nE+aDsQtmWEu35Bl+zEkEtaFhB7rgfEVuadi9ERNqb
nWYf/vsdtYOjABAVe06G/b5/vKzZCVrSBeB6DsC9Aae6LKW1lE/a924U3nFqqmuU
z/E20pA0pjFSnfDA8VNjRGwGlvi1fvtdaFRa1eYmDRQQIFnSdOmYMJg9qCE3j9sX
BDGS1tLxcc7DuN2gy6UFp0iFLyj18fckukYFtZ6CxsV3/jlpCl9PP6JU6ssgaq+s
ACaamkeDsk9TLzU/MXBXi2KkUht1hUvxrVaq4v1YEXff2goMV1Xxt5G+3BsWpXr0
EJqucg5Byqli7mEmmGegoSasmLWka5HrW+6XEZB29O+2r8BqqgwR0MBsylVNZ5/f
TZsFha6VP0jYbAGFZSgLvQT5j34ABRsxlGBPVtbAO9eeTWLh3OfQ393ZN73ovn0A
3/+DEttIAsfRCsNYA1G1hXeV/LG0elD5raI44Npay5Xr+SOfCodJ76/KpaNhUyjW
sDhNveZrfki0511f4uLd1/MBQNjmvMy2Z/brGInw5N9Ud3dtAXGg1K/m7NVAC3o4
Va7dfwsNlvofbpl+qUnlkX5KQSULohUh74jL2TNwvJaq/WncQXyMUDgIbN8IJSSn
3Bin2JobgRWIwzmQc0UbDhCuhjQ2tQaGJ6h4moJMFjrox4pbqvb8erPRb+1VeikN
d6kencTer0QI3e2Gnen/ocnasgBX3dUlvuaMvlv0qooCKAu5ZPZ/dem6L2SzInyb
ZXJaxYaOJ1YypNg8BCK6I8eDkKpuxiCGlAAyhBbe61HRIjKlKVRdx8oVNHmkAsT1
W0j3kPx12+cUA4iqnHwZiwVeBMOq9vLUdhAPs4b9EhFb3iBQ8cBpzzVIsbbn1Zzt
OuJjmFTCi/u/3hbklaB1N/sivOpPMs3mK0kRC7YpGOQp4IAjobf+aXCUcE0j7ZPy
Ebd1wDaWq+At+Zhd2BNBWFEbQ+88xqsDYZVNE5zfEcd1u9aMiapbQ+3omG2B9gJq
uutufW1DQ6hNUCMOnhPjZqp0goTJK/uu40uhpt0lfetPJ5xxjiB9oFATkXmajfDo
loMeSp1CYu1RZdyrLxGJ7XGCa3flBUfWw9X5feG/kWu0sAi7Rv/g7nUUODIoGNKa
EhBCmRNx/b+K169/JPbpZ2YcSpfXwqzqGd5HGCHEw5tTnx/+YL2l9uQK5Y/cLut1
wG7Ctl8OGfRx9aeGnyJUIgx3bAvs1X0/yoM1zvXhZxFGSmffW7XgZ6NTGVZkQRqF
6pURSQWM5RRb95R9GJ8AgzUUIQiXw/3bHd6klwaBORI2u9vv0Ok39JsRaV443v7U
kjTky8Y36lmm5H07Ct4VzlBUsVkBGxGiyx6vltrcRNlTiJQmSFvoJzuxVpui1tfq
QpLonqqfTUcLGwLUsB4wq6i/Vqy6TxSIh7nk/mvE/ljqPfFk+2tnWVThaGjOfhk2
dIHNXT2GPyqbXqBiPE9dKHODEPgDwsgFM+NO/y1ADDdM6/shUsn1d4dU0lfBfb2G
Z0F7bKrjPQBTLKmcGkYHQ9qSTItFYy5xzMUbkLBuVaaIJv3anORN1bCueSH2NV2U
+uyZdaZ8+rXCIPB18ySmuhKlmUPcWY6lUBJFPsDHLRXcE1kPhcojAFpUSkKpd2CF
zOjUkzzwQstZoFzQEg5wFE2GNMCVZv9oRQlPOO6mCPv+1+vd+VIasUqOa3rFV9vi
U12XIze9kmy0O1JwVxmoJz/GgJWJR/QUyGFULkBsTlSpaKVAnJcByh4k8greFqE2
sferxWBCMLhKcS6w4bufPT2yco5lvSTK6dyA6iP0kWzS4lsgM6vwXNHKPNz1NiM6
c/SNYktdrOIKQaHVDKub8D0BMpTG7HOjB6CCC8QC3w3rGuWUEBul3aVALP5XdmmZ
JvPZScNDjipVX1biqOstNFj6kU7Mo9wLv27fsmSBr1KdnCTZUy4oHFp7agfSCoC0
jHJhmxZYDWWbbCGyEGvdL5wuVMeKV9Et31s3hz5pv28nH52qhAUfiKtJq08VyQjD
3OTwpUw0unmoneaKOzVkvD4nS+NH3SKdOdRsGWCymANinoKTOm3AwoUd0FVvqDB+
9lKVJ3Y0UL4eavJyi4VAmcZQdASdMId0KA9W31UlxyK+0uy2lpY3A+OhPVW1Q0B+
RoTh6N241Cl0p6OLzkXarUn4DtObUlkjkMuN5QkdDUi69clFmVAeb1VP/C2RB7V4
Y3YaE85JMNi7nCS1LLIyyU1iDeWcL2nFiCpTe7CfiBcSk+Kd1gu/3pD+rGcySmYf
UlKOgyz7N9eJoc49/3XEfd2fBbUXQsK1FRMEwXAug7EG0JNGMBk+DCSjJSoSxXdp
dq1t1Ki8oWzeK20bp9R5kk5yqe8z5qDj1rt29q5TDYZBg7wJ6+c0iC6pAgjREShU
D85+JpPNwopPmOpyI/sc+bApb9Di7JtMAHrJC7iIatf6txZAp3E1jtZLD8jLyggT
zgYE9aGE1Y8hdQj3sZ8Pp9rIski5/QSN6kChIC3wLQSmddE655omToKR8y0u7TIN
RKHJDL0NQTVOyurCQgdZjilRTkOVn8/xJqDkFr3UT1fuXwRKe0N6tlDqFmu9uWGK
oYXMsqVFO6x11kX3gss6PqRMd23PPoqVZVYTr3gzJcEYqCR5bp/PKhysyoTit5tP
CTg7DxyeomcOugP5sWw1beuxZDc6NdBdvpHbKf7+hxNArgSBSAFTdz3z+37TyC48
WxrvdV4HrdxCvYegGKKDJhNicsumM1F1agK6hLnLe4kyvZgYnhqHh+Bj77/R0DX6
IQJjiyk2LV78RGJ6Ifc9fgG5QQy1T3FhdR7Iti92Ghbx0NxNyUThX5QIHtYXZtCh
HnAfJ0H+ML6YV9pO2JazlQ3OjaPWCz+emJMFf9qkfDuAK1/3kuPVwM80i2UKrrqu
0pQoDgzZsQ2CKuqM+qx5+vE8X34O3H/N97rQgBJwZxthxBK4WezjAYO13L9K6qQ4
YND4i9UbxtnCRD2t8lCRqiz7itKWBDyEA4dYdVCN9+nVy3JPtUarAVGeY+7NwEQw
NBb7B5QgtXFH1Wiugajo4QuHqfxbL7GhInC0r+AbFWF+T9KFB4q9+H3dlKPGeEHi
L5K1tT5buG572XVZpDlAiOr3xDamerKb8xmObDMirM2RvDIXHffzOfTqCPUTypjb
Jcu1TLZZeb2ak+fCme8j64MmhPjLxvsxzrgK968vghRLST3KJlp+14DS9qYpLSXH
jlruPrVLWNbHLkmSq6lEYybby2ODptFvYdVzOzOlTYBym/vAQZbE+mT+s8QqhL3l
+fjIfLSXblQr9QR4NSjtdu9sFhuzoXyjkPiGyQlQcU599o3xKpm14ePYSPABtsv3
B+pWn2S0UZenuJeRdmunRxCRW6EdOu1aN89AtB9a9Y2HCJRSye4tQTo+YJn/XEjc
x8ctvyffEdFBnYDtCk50rN1BMQW/SxZNZzDNym1xF3Vc90z/25DOJ01moy6rkDw0
Klw9mQr/mfEPHHwyasRiwRvZYUMvn7/SPLZ1jZDkuZ7cTg1jFf07BkeMNZ1MCusL
nktiB7BQQLaUPFdYqG2x6VVr01BUtOzMi9xs/4Oxnv+TJfd98GRNKIo3xTc1ZTnx
g3erk1ENoLqPzXjIL1KEpttHOL4ApHshzW6DqfG1VQEfLIlacaDl4vRgXrx0JMAI
razG2qrT1XCiqEn3r7IrG7TjTjbnz04Gnq7q0Rilvxkuq5cv9+i0M5sgB5jbogXe
mjqZlK8iOk8Sj9jywlnvm2n1MxZg8ClxrhyUXSo6Rj3w9LA0AiPSIYGl8Cpafmjx
JGzOVRk3DYBaP9W8of9J98DfYxQWKk0X8T8V8qyn32oQkfWaRjxdHE9FnbRdCcro
OFiiNRjx4Rz5fPzkAxQGZY8JXrZbPP122bNfacFl0c7c9GLsT3P8248H5NhU8z/T
xbM6qftWUUCIIVjTa+zBOl4q1zuIbzbNvZeK+yjeI2d+qFQBkjdR4aGAPWeOW7cd
r3PLauTRLNOg7TyHVeIQJX41d45C2z5gWlfyuiMB97+Rf0lLQGoG8+9pGOBXIJm/
vVv5Y1hrps5jBLB7QgE4QInQ7T/v/xhKeAFOJgZba5gSSIormYDr9vTy2j7nlXuB
p6k0LoyeO4m/UWkQFDuNfZz1G1frhs6myIlCJbKYv0HH86gXnjg0w89ZxlFzes/k
+Q28YxtEyUPTzK1knPLkcdkLXUbpio886pICmGyoL61DAB/YNhnOnhwaZ9Q/swQl
q91cyt+R5ZOUwER5ia35wUlGi+q1ri1laUml2AGAqFntJDTAF1HBUtEeRjO7U77j
kp5Ax1fE4f42bPwatDiqulfh260jWym7v/uyHOF60G1ZndEnX9vhIKkRGILVo5Qb
DDrSbUpVk9c7O4dwu6GZvfStWSvCTHLWUh5Tr0T2nJvlbzCGz3t4n/lvZ7l68pBj
PAOvrq5GKaVZ8zJ8UuEukZRW21YNBFMMyOwWfvLKVyhax4w+oiGjyAb4uws7yfI3
yIS1cmlj5SAi6zqG7tDJPM3v12SWTBaAnNlr1VbAOvRMY/rpUhpGC5X2cT3ERRSR
9+MUTZhpfkMxyUWFJRBpzBs4IybgaimPeQZ1Ql2R9d05zDNXHcd626bo28Z63IE4
+mE4c11J4Ijcv7ykeXHuDXA+k/jM+xyYZxnh2NHqE5ZG5ZtjVjLfEdNYIH6SUcwg
7RdG3dWLLLeOa/PKCdrNILP7udO5446iqSHjoDm5M1JpDTOzOQqHAuP6CPwroYBM
Cg9d3CSNSK4XkQW/xLrbEiauJID44m0mBqGIpSQUQv6KgSu6vo87Quxk9gjM6+UN
gfb9HuCdBgbnNjMuxMrPDe4WLs8npKHOMF1rHLaAfzre80Ob1bZYMUtmln9G+2xN
LfBkpX6Hsq7l1HIgmO3M+KjawTksCdYJB2k69JgZWayeEzOvk5EYTLOK/KXxyoRK
leK9ni7mBOCZnxqFXbMoeMNbvn0oA5qPAjywNLWaXWlzS9gnftjVu+dTIP5ZhKgu
DLUuMJwsLOoL6I3/ELCGJzJfHOh14RT1QXTFDJqWrzIcMuLq0AHATFi7/8SmnEWj
gbD9/znr+D8Y07vzK5rwKS0VqRmgt6JJiLsbV7jbTDjjPPqgYF2dOSov4IyVUUXc
lUqM3TK2clbYLEQcE+iXKkEiknEhQY3IURTwMFrTTr5AIWl50qgYhaXsTYx7y+8m
V7cuEXcFpclwe8/hP5kp1BiYCEKXuuuNYGIW1soT0ovoczzjUnIsFx0XWG5wewMb
rutcUqMn8aRsrsQHZuIvxd/3Ft/4eFPcQd0RCoadQuGeT96Jjqq4V1xGnLwdohns
gP1GNIYJM39TUUclTo/2ClAfcRKP1TePsB3LGZMvj5T4fmNa7NG1mX/OLeUFcuoc
7WRkQ0iGJtz7NF54RDZUle5EbX7dNwNhXlTDwh+gwen1STJeQzFgramqLsKqSz0y
En9cndGtzUAApiTdBZJ7IQ6VMHQg6YtykQDQCS3enmZ9oGnwP6tGPDYVoWPzhkXp
GrGXROxJuSZ7bRc9K2XQcNS2+MV1EtwPVBIFWPr8FoaCmSJPb43kf9snOng/SuGU
4jqadVT5j4rMoDM54PQGal+fEa8YwSkoMO/Rj+hshL4sIpM0vyoAG3NehP0rSg7E
cowEQF+aORD91wx6T86h7CKR2iDjhOo38ztcS9LKHME1qqJ9Z2M52RLpvR46hHkU
zRtS4BUjqDts36jg4PTX3BTmt+FIWZylcLGjRw3ZBQqChf3g4QqRc2lC1jCX6Ove
hQdZebzQe7deThiJPRf5/CBpxxK6MkPcHLwskLPfXGejDu/vY5UYxOjO7+X64vns
09dsXpjLSYyrD7XnhTB06ddC7byY26YVgKtPewyLCosKCovVd4B/TXcRsgGRCN/b
3NK0KnQs1PVPpiMtfbvuEXHYctUpNFeiV+x39NGCCtyKNgFqkuWIsADkDKTA26Rl
BwygbLC4QlC/IGIGI94hDdYiT8144p+u4nllD2hh6p4zW/thXpm3NNznJj8HE03h
siqxS9QyU4j4xtIwjKgIC4TKbJd8NvFgC85l++UOmDDhTIN3VZ2NEFwCe/xkchkr
Ebahp6H+jEfbKVeCQNmuc29q+JT57rPpnvvigC6lMngbdcVIE+vIlWa24ncErBMi
DXxw/PRY1XS/W1FMvKevoOReSWqBG5JiYNIUosCh1sVx0FRupgVldpOatu8YIXgH
d2iEOQ5CjqfwZjosCLFAvO9UbGVJM2gtYLSGPHKSIygCxUQMg0A9C/R0rEQVL6rd
wJOLaDxkyKkAqo8D0e+gANW+R9PEIxyqSzKPEvoxEH7wmj18Cu1tQq2otPAmMSj+
XsRhHwmiEjxRqPTIbrMWve9gBQhxjnSPRGNOHL5M9KCv0QEnJAfGzw0wV+9sTKlF
glaDKcRhXQXic4Y3lPDHMnXI/UNOAoNXQXCT2B58BlJT+IRwmw5hehozBGmcBOyZ
8kf5yA/KAlOl/fu1kXeiYV3AGCiqNmcbKFrLvCQnoKgTe1kPOcDYqzbJQg3i8+5q
+sCptpANwXwUlDx1YFWJBTt1Zv4++IeWIamI3RB2XptL37HXJuGXwYfuusXUY6/x
on01Ut03IYP5zzygQ/WXCR4fQ4B1Mo0yghcXV9qhhUkX1d//ZpyirNo4sON1uaZN
4YO0SWDQKGBhMy70RZBS5hMhih0TqIgc1u77VrJs+H9Mez5dA3VD/6zB6ZZED+v4
SuibZo6QFlXkuaepcnoendWPDDKjN3dnQjkUuGDbwfTCwNdbtAP3MqIIcv/2Yixj
trd3pnhWLn2nvdqcr1YtCPl9IZZl86YyC7VBK7HWVwfdfe/UXv1CqST9Bn64rYRU
5y4u9JeUfOru/dO5BReuCh/SnNbyHax6JzmtfFON4ZkH4CqWem6DHmyOiuGSyqDM
9XB44XQ5cSNvjI4ftaLBtdN8uiF471VOfPb/O8y7oioVl5jUq7G5Wx7E8n+5mgQq
9O6wSnJuNN0ifyVfAXO2LJPxcyQneUNUVxLkPjtZoOzArreOrkZMRMLhDjwQWYA/
RafScR+BGY5zC8jMfuKPkxrDQs36VflPVoJ6j/hPPHnXv76bTTFjZP8wtsQW+TIP
wGgF0JfdUGzeBJX1bDCYlo2ComBdcj1W43nr5YP567iMY9oH29PuUEzyRqtPkSEo
4fU3EWtHEyDol+7HDgsdkG862ixYDCeHB600wDpEwDa9iHsw/7GJQeeJAMwwldXU
BB0BCOt/1ODB5fP3Vwd2YwhwQseBt1eZ768aKzCdXURTQsqYKrUrghTPE/OPW7jK
Gm/NZi5Ujcm6Yb6azidG7R/P8hY12kkAwHnZHgm4K1yW37bCWPnhbV0X3STsfXEh
zgf+QgzrD4ClVW3uIZZGgXycI3ApTwPXN37MV+VxocHNDlyTJYDnD9YcA+ZbOcfx
DZ8WVLQrDobqDuY47ss4W7Rha4+lMgIc/zdhvO+aNUBsxRmO5KIBBx23HDGtyPnE
uWQJLPYMD6cvCrb6QJ3ggr9MFTMcJbmFPaBfK7trVr9X3GI8lutcXl8ifau0qk8X
sV/3HPP9h3jYtm9IQGrAE7kmFdgW3yHjwjYPXPjNLZ9Bxpsc3VMSsoIzbtQ/9OT+
xRR9wxeXJNMfgKv3eEq+f1VlguEBBIFjMu/3UJu2zmXEtoLw5m19GblvA3ZgJ7nM
1rGSX09tG/abzgJ7l7Ly6dEkq2qDuUjHJZTzPJs0kh5D6JqV3xZKa4Xg6L9mP1nK
iqNP3UUDfImT45gwB/fKLs2DnhnpZipwHfrNXIm4EPD/2TCRmMDPsTC1HGe7TsbZ
NGEdgYmo2OKla8RJOyGGj0dXjtl2fcY5p8bIRQnDUbCSzFZ7kjUtmMudX7znV93r
3hun2nhcRQOO6pN3kg7d53KomRblnLHTakbZcR6xbxjApWh7WEaExyH7vUFh9UeI
HQD5Dvzu+xjOnCaVYfXxXLHxS5mTG6dv7NGQHgdg4yEUJUGQRGPXdFSp1CgDhXnz
1wGxAAV3C8SVd76S60TDSSqGMa0FcBVuuqZT1b1sIiDPSWSdm3K/p/N+ZVlVyJXj
1P/ueMG9air43b1nPt+kJPMnqZQJlAzDB2OMnSADMZksvsF+5Xd9JmpIBmrhkHcH
5XTGOPdS//fTld3AEKGGILyUKbOkffLXBx49q0id6BjanVIkFkgRF+BOV3r0b6g9
oEASu21W0ebarYGCXIQoi24XsnVTVcKJDCIOSjbTn3wF1qldbwC8uE8ZA9wMGFFC
KoEaaiJt30InxeKbJV9H8JAPVZ0ZrSOkf/bQsO60vBeQueW/t55aemGaYMmSS9tu
du9ZkoAK0FpamObx/0fxFwYRaY90LN+is0GgpPYSwAISVV9BdNGEAvIT8RlRLamS
NEt3Tv4et+249VQnJkTOAvoj/uk79lh0vwbCGt96s/RxOmQV6rGC9Tqw6n4jKLvK
dKiIBQpTmPmZqDVafZGbiytdDRa1ZKa0JUfXbsSEhKokOxJvWbTD3RYlgmN5MoPO
lwv33i77e59PeYr8D77mQvu6z6vwGtPVk0smmtcpVkO3pERGI/nFX4CKZBD6CcCw
4iuTLpx9Lg2aNb6m/20jikcHXMhx87RnFzHsttSrtoes5DTS0sOuFHFbSYBLNKhu
Qof4ITo18J6U0ydvgzlnI+RnLN9YGLLk1ZiUMHgIK33hDVyl8dUqzzF83LG1J+T0
iJQciQ7LvUVJF+SA+/R8w53FNKmUm3CiENk5y0z/epLGW71SDyr3qbf4hmmv7Y6k
HXrwn4PWUaF4ZVAaGM/gVelXV0uzpf30GAW4DRSxqQdPiyRGkGOQEDVoVbhxyfOc
pF2U5a5RII+MV9avM0DJcf/VTtw67ls5OXo3pywKcog3e7bK/RxtJlFAaKQaeLeX
udikoH+R9KyHp+iNctUZvkWDHmTY5+JVWR2qCbC4O3Ylp0ZUb0sqhQvyLLmgF2fR
+1WSkOYJdGzECAek1ZGekyyVnfYeXZOc1gwVV3P2HRkS/L7gXPpkR8+Wfn161dbX
9k5+VL11hWzglftlcJRVYIuBgi795EIRch5rzcqHa+WchlX65EqZXxt6/afoYM1q
2C2vJXSNrKDAXdfipwvh4Rm6OoiXpfIJ+45G50etMaCF5om08ZSsYA9QxLfAwAGr
LiIfFh+Opl/B+/ppsrMdVK977/KqJ8ZdZ+MePkv4TcJ/TIeRftQaDGu+ZabvxDNA
r7+xbYJcpp+y2IpoXidyj0ThX2NSxnhDwKflFxnczaPyPPtGtTN00jax3izZ0GeZ
cGhA/MvkiiVor0OLEibp3m0HOp9AoBz4uKJO2R+2wONAn67feFHGLVhodkKk2wQ7
mfQH0gI60xZqRy2+zmdm6uQZS7Ohi2Joypv7Sw3T1giMl5W6IW6X2tGxrGTCa09B
zYmI6swe9ZidbTx1QeNKzFlvnd8be66y8YeDvao6OPy51lk4JUuyF3seJyYrxRlO
ptBL/htr6U7NAUFCMTv18ccABTuaNajnI1DPZmRtRveGzNmJ2zUFseODwTmACp3+
r0tb073J+f0H92Y5rOrZAAr4quPk15iBB9sJYxqQVfvquihpjSdyNYI49AI8kESD
iEFX1dQdZeXSLY1v10EVBcl2nagUpEl4Qhlz/BAW3iQvl3ooITQPX1ZSpon+5NoY
DD6jPy2D4yke3BijswnBHvjogDnt32xMS3aF/N8SA6mn+7Bo+a21UPSvP089P6WL
51hzjCz1W3enp4RnZo6ylcwK1X/r7Kruxn8Q38BXmIa19xJ9m9dnarrIEX+KHQi+
+ktyUVq+S81GVp/Z25kHJG76DwG+s1BMy8xjCI59v/rQIPhUhA2WxpbQWR5+WI74
d/FYM9LJd4wmZRNMZLa7NPRprv3vgUkOPOEQgrgxr7y2e6wmz2f/kqGdf+nvpIRx
1SSUO9h3+Fbbf2r6H12a+SLHYZ7O8qVrnWRuoqF4jkx3v/Ppi7Xexg/aUAFv7LFr
e5zg9G4+1N0T9Ei3ZyNhVXF81pUfnLrDPKKOo+tEM6UGB++8SWzPUZW4XKknekoE
dMl7BIml+er28u0WLRheWQLb3DAfq1uJ8+uDytf9LNBoiW8QhO7MhcVju1VsWwzW
RzBOqEF9jyqmDk/hmJcG0ET8CWNbx1mOPIkw8ilzqOGUBuYIgD1wHOYqePIilgSI
hLoeWcAl9S6JTP2l3OykEy5KLoI6McbaZaupnpkEKO2056xvEhz5TZ9AK+N0MZEB
YHdal+aTwlorbHWTFHp5vfYRcg7/7rGxVvQTkjLw/ZQ90XLaa5FE5Nc0RilUj0n1
kzLKFnXJpbwg5sM+S/BS+p5rMJKSFgzZyiU3FqQUVwiMc19BxxCClcJcaZZrIKZ6
vMnfJ8z7Md6PRdYlNvsSGlr58xTpxV+CKidLtdn6pFN2T+m/Dk5WrQUrSrDug2Yz
bnODXv+oSE9/43233Cle4ycxz3HE1y4lqUgF1iQeXm1Pb8Up5CQ3mA5NXq8vI/B/
+yuKrlvnpmBnu15K/TbHi+zigOacq4/nlsFOLlN53VpFeFdbei0Q3sK/eZyPzvcX
rpmzLhfTGdg9HmJxiSPyqw5wOTQTZuvtJ9jk7EMVE66wpJdCXaaroMAcSLtL2lul
djTHTNLRrn5TnZsTsxaK1oMC+8ly3FCkjDdFQRd4sfDy5FuDsyAVEV2M5ejNCtjj
yR76rYCi5Go5ZApN1eBuNiWcaMF3sngM+6L0wX6dTcGuDk4TsfzB1QarmqOSASyz
0O4tiqGOLjgRDTlXTSK+Ld+FN8Qt0JDdUfRhCM1HCpGqCqLHGZPi6WKNwIqzFKkn
e71BUMp5teWRhCXXiZaYIKRzLP1IEMT76mQZIHlMPvnDDu8U7Doh4Fm/V40jkP20
/sLTePrt+HgGawtj0uR0Qy/YKoQF0YiINfrfK6KpBJCOkx5QrtPBvw+4z4Ulruxd
P+E8w5YbeT1o2kjY2nKDiYM0ZW5GqP9xTnJS986VgkKYpCZgKM+/qo8JJrT6eoTV
jlBCzVoN81qaUJA7PKpnxY2voSyoc5mRoa+256MoJgAauRnvs23zrfPO7dK2e3sh
fmBNWjEAe2KHPgzxv//jZ5nWb3mZF1zmNLL52gmhVQyw5W9dLp7whwEPPNg0o9LB
iYpTDu9UIXlopCXIFFbAYO/eKoPKuSzmaZUjCDKUAba/3eIn3LJ4RFA95brtyzQJ
8Mww8FPwZmBmkmjBdbFsIuOh3bUCyieDUe+RKKg3KMpDMs6RNmZQKhWcffeQVh4L
VQqa2aO47yI9/6gseNjTEW/XQI939DE6VK4Ve4/s23mjC+MyMAuvaraHICv30yOf
r6fQBTy4MrzgzPZsDrzbWEp9kA6W+2fHfG7wlErJ+CM2Fo5c5b5vzuHttDERcURL
Mdcmt+AOZbddR8H3ySy6YWRTUJqxQEiHl9fZ6UqE+Pdc0q5N6j2EFPeCCIxzVMXJ
aALvHzEbiZo3/AhO0E1yUn5J6laeLctaDHgS/a/gXUENYYP6/Ox+abju2XHFEeml
NGvvvn5Jr2hDNKi+AzdtsOfIQ5ZU1HeA3nHe9CLMP03kYyh8fKn343petHMlSEAp
ZZcTve9ur8FjKjJs6AEjFFcn0keREc+YxnTHTkKryl489uSvg1hc8RcvPQInvxwF
LehvGf0JIFZkb7Cgpti1UMWPxDrYfD34RgkDcHEhOG+CAveHyt4W85HU+8mIywJT
zrnk0inAdRCfhDY9kKgo7/2JxlTxFrW0fNWDhUSlsmYNwp6IcCWXRzB4+38JUe8n
yjaoDxvRNSg7IZemCUqyHrUiWM6PooWu/ur4NsRJep/fdYOrq+9xwybuljdMNeqM
ZOk9n0ibmidI/jjrYEDQVvZ/B+sVt4psV07kiqskS6z/9JtfHqWW4X5XJMBBuPmT
T7jAMttXHCgxopIlO5x6wFh6VUWEHmc+kVqf5cb8dGpvjZR1CG9CnAMA8Q4asZo3
JiKuBWaV0tEmbwMeq3WepWLe15ElxmyBJQdoTI9KMjy1g3kGHs0JK4AHol2/E7Xx
Tpz98JyjSmwZ7GZAaXeXwLOAh7J3FpcK9dsfboaUZnlHZRB768iNhvsrPDY11jz5
GQVhhXvsuMul16Qu16dnIGAuOD1Q5n8IWS+RJioGQKH9sqJfagnDY+3NiuIlbGNT
Ce+/0rGYvA4jjGXVHtnGZDF3/QX3dOWUbBXAiVlcfCk7ijgw+NLhVhaf/wcyG7O6
9rjuytaZPEaWwRD3M9S0U/Q6nJ8VcLi2siDWWeBMXACCzNfzDM+DmgznyDRWb5tn
wUUh84p4eqSWJWtyJBgut/OKrnRLU5s4ide4M/ZAPh8jJwrFZpEpMO3Q5ojeGGth
KuV3uqZ5k1UGAkJof4DvvurF3I0CcrgLgNFfdccGoFwkNXLeFXddNhM7847vygec
eiSgF/s62n4bBMxf2HCODFndJX/48j84KQH8VaCYrNXJzsg7pW7xONDp0PgAogTN
0tewmOau2ruhJFZhaxjTe9EBusukfGnpS4FlhkkZi3P9tfHCd8m5f7dPEN0THY/Y
Ud0IdsfFxIQlvDs4xkK40d6Jx3WiOHUTR9hIKF1WJopb5o/7zBRZLmM6TD+GGA5S
M1eVNWAbH22i7OgtrcNLBUK/V7F7vVLcDjpEYOyJvBkOSGZeOAY5vDTleKmdudWe
0kbw0hVTcBU82rNMMGc6nv8rlEkCk5apjIYxOC6kdEu7Z9p9OxYImcM8GtK2LEtQ
BBscZydsfBW/UE5HwlrlVh2dULfOD4HyxfAwmQNhmCRNn4W6ZQyjP5jIG2bhImxU
UZJdavbNqQ6spC9ybODp08J9Dzsld4TXJR9iecTJ0xVyXWTpdbC4nKEoZWRfiaE+
JNZS9ACLKFAYwgb1HB05uN0mcEd+1BPeBMgp3VVNQkITH/IcxAZzb3Jb3TSX3+Uc
ZXuD+GRoVbqkffMlHdxCt4BmMMkAvHDabjSDLMc7W+z71T04PcPqc5ybT6kt5G8H
KbuN+jlqGljMEhPoRlz+2Pjc+bT2CYzKXsgdbY1QH7emDVex2XFwgd8a+4n3RHfT
7zsXCxMoFa677+7JdSyfeX8RtfdLK6kquQkUQFPrawMIzKJpXgSeQ0AFOfCS6dvw
OGsGq7CwZ0RLEDZ62RbYtLZ5oOaiv7yr+NAXQiNeA6OFOaXNqM4fyn3RCDfX/N7C
/RFnLi1ajXdN2kgPcCeIj6tDwMG4SWqSqXLNyuHx83tOn8UjaONmgaHvkNmbKI/S
QrmvTzI+bA7srUfy4iltKPHMgyPubTnmAWTXYEgb0L59SHKowcjt4c5khy/rBdJM
5QEVGqlqQL8mmsnX6DqL/K2y7RR5bQy0gHGczSq1Dd+HW8TUroCRwEVZp/iHZBVH
5PDk8jUrJ0Nt3X5vNUfK3hwMw9ve4WBxPEQktCEnKggeMOnKxWYPjpbk8+GW+hJV
p1PveDJbtLO1dFcK3YusnPDP0lhZ/FePzKYGefxt2U5k2s0R5PyzG46T9fUMBAbm
1TidZB9FntOr6vuuiMVBhqgI7nDErJeVgdlfNW0XfvzZYRhWX32DYYcpjj+0TtVI
RPglPpqr2RalhtyGPMwPyyRI0KXg8P0nYSDWhWme69BjuPSHMUjt2qQltD+bU3Gu
+rzhVgiIIQDbzx5XIg0wxdUmcl+54StZOvh8LxLZ3A4=
`protect end_protected