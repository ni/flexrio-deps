`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Jm2uGAVYfY7w9Y5qKstopObZuZAEY3b/Io3MSEcWLhjjnKulVhCBBYAEQrAzzGsT
vMbffkdZgjdXQUg8jOLJXSHZ0Dgbnob2vlppjZs3bgyHCF7MoJ35E+LOsaLimUA7
hlqStcK49hR1hdeBPr/OwfT3UeVrRtQyq0eJXQ1UksinX1G9Pz3/CmcGfTZ/C72x
p9icpt0bkY4/1I4GBvNCsA6FFKH947JqH27OPACiQQRW/K7JToQn+1uhWr3LA1od
lbVrWu8PdZi7zW9gK3jiW5GaPjwbYQGqeGFs3bTKBILjb7sYHxfxw7eDLVMAIu5D
W+OTIN4JiHiE1gCnNEvkSQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="pm+c2fYA/4JT1uhlJGVUubML8hZi8lME4xPobg/m8uM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
nBaXksR//iZ9fraC7WMJWWSrjqRXHxmM1Y0+KKN3b10NElDzVNMlR76DLrcnamFd
2n7uzsxWqhhJR5LBl98SXO3Y90J6BMbw+OBG/MFM/zUulxh2Si5YK5G9GCrG9gvZ
5JomxuZFDu9CzlWGTuRUt6FsE4Lr6sOL1P+hraQDpMk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="M8TXDiNa0BVMX1P60yIvW2WA9jKGGy8GtbuPknDnC9I="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 29664 )
`protect data_block
/5TNZvs8Nu0G+mfp7M8H+iVAGG3Mh5DYZ0Gn3rRNhV8b5CcJKgjQajrRoGl/gSxp
rBAhtT8Vd5eelHgtvBjpvFBA/EBUrRH6CG6pqRt9r2qUDt4UernbZbxC3BC14KYF
gLiaAkKLdB6NWFZG4rx6avxlMuuYaRQarBkB0XRSDjNtiDKQ8hd7iFgaI2XLpX+G
p+dqrrErN5tFljZYpMK4YWpbApEOhHXDt/DtgMQRLauxi+Ig9iPYdvhAJUSl7wNm
OBeD9TH6U9wRs10Q2Ckqxns83xXYWrUt2o9ha2CIHHlqs60q49prTaRZ02rKYWWn
hQANZGuhloE5puLMQBVi/2ctOs6AsFoahxB6VKG6k7oNtr/9aNCgCpq0mYG2aq4e
z8iULwWAnkjGjbSHFEbuykEaAR1FqcnWr1lCe1xguqME+v3GeEB+bVd1yhICijBc
Ks5EWvjYmylOKcwzpa1v9g2VV1A4RnojHMjLat8qjD2SoLUMD3a4Dsz/OAxnWoWA
8C5+/TsMcZmpOUhlI1UJKGl7vDyR03YkmzKb5tE/r7dHOQv1a+ZMnjQQGj0DSxG6
u5I0c/AkL8KY6KFR+1tEJwTAUbiuAtgM4Mp77WPLGNWYS1zfgzJcX0qF+zOvqypR
FxGULKBtnQesPYK4fdY34VYkobQCk4guQDd91iYDx6KaONytSq2c2Nk6KXvFxG9J
S4/AfQxsHn273HzF+1gKZ08VbU/5ZmGuY5AKJdtzeiHLoDbMtUYVusMc32wGZHRf
MaVwhtuHj3mIGHg1qc7fjdOet1p5/NMDm+duAHViH/Y0DMlmtSctdIT5oNK45QfO
owoujA3xfCTYv4zWmsjjhWlCoeylP2EQV1zqKihjpqlejIipBDm4u0mYOYTaTO84
i+mnsw0RDnPI8kMLJjHIO2ClqyGQ0TplJs2Ux1o+Q1vfNF/NHSGPxxx8lU07hlx3
sJ8LEMW8gyDLkA3ocSckHxL7Naw9BHpbbnkLSgoQkq6cE6viLwVvtL9nfhVz/UXV
fpBOT+6SJRBEAEpFk2ntQGSgJBSRcuw6aGtxsD9J0Dtiq5eqLeGdIM5+gwjFYtOt
eckEG/prk0f1HMxg9qATcN27vc5VIJ5oxR3IaS8s/VntRlECeLm/C6AWBqmX2zqb
Tb66leeXxGAS6pL2OvOOVxetRwOJQeU5XaCYb/ykTwHuumPIAZtZQlIfu1QgC+Nm
+jZngkSSbbYU8h0nOCY9ML5vc17PXurDy/yNUmLklsOEwAw+9R28Xo/15XjuO5mh
1HdSpXLYQgs59KH4Z5juB/z2x4CWbQySyELyrNl6M2lpelwl3I9DHZ2TpRahD9qy
wyZMel8RtGiHdceDA5asxEQ5kNIr+A4uLJT//ivmnMQ6iBEiPgAbRLPGuWbmqwfS
Pvqn183pgJqAW0PnPvgv9L++H5bn3nbJVXqOtNg+A8ekp0ob6N3zvWvgtmEuRv3f
qkITeXJuSZJfu13NTpJz9FnHAMAEBEoV/1qre626QDogKGU12pDodKER+YCNx2eI
FNQmhH7GEd3yOmQoXt11vskD3/xjQDMXu4zGBA4L9iPhokayfJtDM5l1j75QrP6h
Jd38/mJlanhZ1h6IfeAiSCh1mimeuy0RCi3hEKW8utKzu+EU9W4wxQbLXD2h2iEy
xdjD8zM95MaYGIcpzZxab7uFmSoelY05BKsXqcvwYqOHqrojD2OAl6DnZuKVFsJT
GBQwh+avheEpvpq8V7Z7pTQeSwzVxzmlGGXPzFzpppyVU7Thiezwkn1bQ3WHQ3eg
RwxNq1isOV+IXsMpvMFVV3aYfvzQSqc/1rXDQzPz9tOUSjogIDjVIFx14Q4EvSQF
0Q5GsIoQ0sest+Vrh4xfkN4iG0N7fjdQt3b2GE5I2A+CrgWYdcVYZ5971wT3dzcu
FUjawN3dwsA1i1CrSCJzAly3DSUCgaGZs2tej4FZVdGPn89pWQuS9h42PfubMVPv
JAdIk5dO8I74WpzkUpMTPanBYUiJ8Pr4bdQY5054qroDFX7bbmFWo5HiKe1k8UQt
i4MBnQcNaKeNLON4tOdXBqjDNyO1dP1217COqglYOUo84aKIpqWesj2KNjlJpqVR
ghAgnLtct/UcGGknL8VKV17tzVfy5tSUc+Tmr5qWr/e/IZLpMw5BTarKW+oDQ1M5
qkrL6Ocuy3BKdegVYc6aCOJA24BImfu/mBQkdTSFpqWEh55YkLMn8Ym1weZA2Nux
QRB/60j3XkqtkydZuampCmJlkXgnOYTn3GmqL9V9+nkb4ZqhnXPM3RY0twvVBvct
5hHTNkbwyD8f/c8yRf+/jfjxopIYoQf4XJTH1YU9+rFo9TlXsr4WWAD/hlRr2aH9
hXIdb+YktaaSjaNbN6y3AgFdaRj1tdX9z9rI/9FwITzs6zNrMd4ONxxTH52GLaUl
MQyDvUH0a+9kKzg4y08I+otNtW6bJ2VQLrS7MvrZ5pC1aMF8bHAXL5rrPgQ8IDsB
LfVmad2Jw5iNMXogk2Yf8KF0z2m0FsKKf71NBoEHRY6mWKKj351/Mj7fDJEcf6x5
cflRCNVNgs+CVaG15vVsBqqaGXpdGrx1NCqn6S9CqyRLQSVzCtrj0yF3cODFGH1v
IEDJDKI/01AZZIv2kmU/eqrSMQDScmOvHHVnwIBJo09irnGG8Mh3x0V7P9KaRl4p
69ID8aQykKBREdl17T35mf9JF8kH0RuApbvDD2moZmX7i8C4mPkEAxrhdFCQDezx
u6Os9g30r6t1Hgha1llDXJ4BWNRT66RkbHuH27W17aV4an0u1AgdJM83VeHMNt+/
2VJmczTO1Y8vBxZufB9o5ZbMU3W5CYxb/NboqsE0K4C0N0qLPKKkJqPJlHSJcDC1
GSEAullkUk/OzOA7i2WkrjereL7cTW5Lax9lF8UKiUJILQ5VcEjYwroYCeO1eFMH
y2FqodEis8sF9YL+XtsCg4QRL7X2n+Gb9IVwsS3CrPwMaqtWz678r6yuoIzys5Gf
oSlJBKVWgqSMkRzP9TSwb04d6TalHjBQs46K9MrbOd1lo4yGVPawUV9YMzEBtteG
ToXpSm0ly6kLpgYE4Xs8Up3CI8bQlY9TYhE7+T/DC9l73pCsYX+6xG8q/3g0njWw
0cId6d7+Uh/a2kutWXWJAJ8Cd38piGBdi0Fa9OYkirTNnJzQj3g5tbfFBJWS/V0v
9txItRzcaOKlUTHvRKk6m/vuoJ2O2c3RkFa8J8JGypRTiMFRN2jLdMug3D1RIVJC
eOS/P1B34c3tePDNCzix9pNrVWu/FprWpLNicqzkSk8xp0MiSZ4xbife2LFxw4pO
kDPkBMuSMW33rtPDkyIiIOqi5m3CdUFfEybwa7BAoF2gjSbAFnUNV90jnvTKBC5L
5cxF012QDe/MJcz80ow+32BTCSs/pRoSdtQfGnlcgpvfdxJ3iLgYlKqh1PuwzzO4
kaZoqwhReqd0IPbt6VZRYsxjgXF0RR41eS93J9hP+9TzBdZdvhdhaHmNwGwlFt/R
3Hq/RJNXtBGIqYlLXnJYFTgY00j/XWO7i0jd3q09ikgKQrhDdzlK0iBwZi5KrrRM
0eFCCP7s4/cVoVZhzeYGQXCzDCbu/MOuXGHb7Z3TpfE1up0qKSfR/o2GihKB9BD+
U6TkeW9zFT625Y6J61I/S0G7mCiI7T6KtU3wZEmOHTdeVPa0qmr8G6of1XdaWDKr
bnh6hUt1zQK0cL9AUG3M22X+o1a+eGlMg8YSGYcdFfCCeVYhqodvIRH6pSDChh2Y
FnabT+HKdwpPEA/r+2fc5H5Rv6XNShYNwJ3Iei6Wxv5F5WxqkTS0PunGTVvbj00s
DiEcdmbeFgRDiGKcv5xNXDcql6M5FXYWoGNuvFzeBvBdqRu4qAqfSO3eJhi8Z6tG
e5RviifMZVqV7NSxJyKEbYMzJ8H27bB2WoXJAlxQ1o5GfM8Y0SEtE4Kv4QNAc/kt
xJlC/BRbCEcJwBeKFxNaMy1WQb3aNrGTL5hg5bGukha2fqwSAv84j23y3xDb01WJ
YmIlm+K2IjDMWu9sOPQs4N35WNyJLhg/xDSPzR1wv63TzCvcdSR4ACzbXPtJoYXi
byPw5TXYBlu2HcKYls7vx/NKhUs8bwdgLpIAMlMLTtSxnqLNV5vDCYfThwLib0bt
F6SGsU9vpAtoWfJr+aYU9P8aDjVY6tvc2G9i5NdQKZouyY3N0okqxhsFsZuotqL0
/OP9to4tO60FOIUtyfxqUN2odxSDrJD5sHdptcAskidH8zk1HFUzdBZV+Cirz6Ia
7ORgVaVRariFvK3THMzMsBsu0mDEWo82IHbG/pwTrFOYChRkvxqICixeloXOe2Rg
qXba9zNO2jB3zPTyjpnnyIk4eBHQd0SltsKlRjkjKp9LE0ksA0AUVxZwxtZu82uI
v6V+/kCTdPMdsi9LkjZkpiyXFdg9K7yauLxLKoRfleVIM9Oa+l7kQURdARbve1yb
+ixS2gq1IKVC5/ssvZlsSJxRELdGX27DG88J5gQuzFqcKoBV3OWTujB1v2zE1M2U
+W+fkpmhxpieuNmeA/qUgeck9PWvDW9PTxx7T8kaguZeRxMQ3UvQOlsV+KYCnZ7r
82hZCFopfMBJnZcaVpqkbL1ZBKRDDY3CLuZHuOMqwLfFz5zGMJyZwkNSw/sgdbl6
fS9iOp2sFJmlKG6DS10oBW4Fnk4PqKT0sKDh2rGgsb53LMyIfo0iAo6JInDPxRqh
Mut+6GEfRMRdbcaBpSKkCQwg29b4huTkrCBS5+NvYFjUY9xQoc9zLJ74CKkr9nLX
bIbxo0y5fIAcIkiec+PBTqjj4JXbhbyO17E+0oRmgCnGUhBWeWA3h8PMF3VPyWQ/
v8zlgOYiZXeEIpZqMCEML1HwZvTdMSM7AMuv1wmNDL/zhfCZk6HotGuzsq7tUs3z
cB4M6J6ATlMFbUSKz1VgHBAbHWbd+CZMQbS9fRhm0fKF9ps5o1FxDqIqyweLdsnO
BTiWc4ZBWepoHOwDZzoj4TkiXL0OWMJO2iB86lbAlbSNzMZpxt6sbNhkfYqVGg7I
r9CDU5UmWuoR9yAcCMHHRhpYDMLUphG7l3h0LHFfcijunkDbs2/wfzIu/vtIlEMh
bCHQgEs9XaXWuGRl1k4fzQZSKmQYocfXeruGcLqZ54xh/G5Lqb8nQThYhTiEF5es
PRIrtFPbpsSo5d7sM6GApCBCYW8UUQp0/HOOzZY5GY9z70RYprxbuREMhmasIi5z
51SNZW7KI75xzxjt1TQUb4fL/RU9nasbtFQVHW7FrufhoCiXL0jw4HwmnC/Pnfpq
hdscEE9VHmZkwn52OBUUyNNLC7HB9HHgQkwAyr9TVMwSUkP5/SzbzOAbMPDPPhoQ
67+2nbcEDh1AIERxzmedkPUpLw0+iK5QyvoKxuDqTwDGPLpU0SKoAUc+8EDsNoI3
rCVUu/WOlcaIs2w/7YUAYrIjRDQwz0m+QzIVAmupoi0uzPVZmdRxYnVh4CbFVGmt
vBDOgEe4AD50m6PTCYzltIcIb1ulTsl8qfJdRpWIAeCxIs1c787/1mCcZphbUhLn
cAuA37c2EZ/DvaSMYbA3P4QKy2MU3SgrqoEZ06AfgJ1pEBd9U67FmK/UHC+Cpu5l
+EH419/DEBE/jK1afliTVOTuoXrW2gaQbp4tAaweOSTWOglEN46AzZYQHSuZ/2hC
FR+DPMdtYn4qbNF374niUZIkOM32DJ9Fa2UMo5FnaryZgU4Fqr3fCzX/KxEHwhxb
pWc34zGjw0gqbf3qXLAzvF22UulOHorf5iAwBXVQXKEyVmwAKkpteCi2DgZM9JYU
MBBm2rg4jnGh/gIB0NN3r9WZTmxEykV5PP36MoBd+Dqv+urdWO28No0xJwKnHsxG
5bhBF/L4qrKi4TysjLGOJe3s4ybUxPUTPxQ8dCxXmIsH9sEJUUqxOkab3ztNYfSi
N52UDe3r9bs9SSVLkkyJygxmCpOhZ0QxlwXmJuitEfpbmjv02IYO6DEvibl46TZR
YNoBC7s5lV8IykRao/I1Q+YPCxgYQs0xzAiZ2lmtUKybX3yYwvLqzeae+bpv0qs5
fwRvZUoSFbpKZv0TFDkrANkEvrB7ysCWfuEq/jUEGLb94+SafgtIVFwS4ivPFCHQ
XF4URf8r1KSrfiF9Eaf0yFcPgf4fPOsvYdgBPAFPCHpTfm6qApSh6mSJshkXd2F6
I887HikHWtth/ccOJ+PBh/Kl4fZEQjkB74QC/GDl3iqRBuL2NQgTgwLPjar8qiUP
AeQ63syFhJKwdMuXzwaxIACqKyhKXekiHOgnp+YpyKsWKXt+rABMwM1W9rtXEJe4
1m8Y50+M7I/Pd38rfg9cUuV6hsNtmjirz5zB973XkT1TM2URn1/5j+G4TaDyGjAF
54ZyVcjhxZjskMwSD7nUUBpJOG3req56edr93LIei0NEywy1UZjoqjxy6BrIzE/8
kyCfWcgrqGDlfm7j5Q5NWzUA+KTmA+O+afVYMe1K1vhntAjemE2IyxiGL8ms7HSp
8t3UQSS59LukEvW6mwioBatSrbOh2EKEejNKkk7bU3oiTmjOV+7mZgivRKdZuSpP
t6DnspXol+Lb/r9mw5RDBFOSVtoA0jpYWfMkCDbSil6leW0oMG+oiDcwKI2493Fv
JpKLWGh116I3rMgEo67KFUBKYZR31/mKzHqVWye7ja4H66wJFzg/KCP+G8iq22dk
ZlHuDZcHrsf/rNgG+7ymYJyT1u3ol77I7eoyHv8A2sAxLHHh+sMLXo3u/4AgyG4l
CawM75Oe2NwnL98aKONs1V7iBJBjiKP731fC3qSlgrSpErVu8QOve9AY7tFHdFqw
4dR5JtU5veTjfBZQT2EJYUumr1UYWzVyJI5qrdiXqwRPJscJZ/UXKjJue/qCMOBs
DPuYSy6RnYUgaX0t40oPiHwiuznp3QvRrtQhKXhRJu+wRVWcCCUqhSyI5lKNNlZ+
jrGyvjh/6hSa6aYlUHgo6rzCF8f0vy8Kx/PkVCLpyz+yL8hEWf1l3N7wbeCcaKDi
SNKdA7AN1N0Rs6AZTo2FxhPzqZLjv+x6mYAOuY2rIDL7c7RcklSZcXENP9bZJLLT
TXN8PYwK3+8Xfux+VlksyW5tIf+FJ1o/eDTOttnEHS3tAJOG1Ogyr1Q5Nb7ZjB+p
1vWVrTqecXJ0aR7yxtAunIG6q2bcJA+5qU64AlAfNpzuangCZqvHVbpITCfmPc40
+edfibY0ZvT3P/eP62NKctbsmFQf81W4ZFT54hutQF5q4bVsKm6WZMASoEfNBHDJ
5V1FoUw/2CHQi+hmjTBlSqB0QPZ8utzV6p+u1GyqA4K7TjaEhpWs6CtsdLHOwVdP
YjlzhUAQIfViu4brPCvH62JmFIfKd4BHhkUD4cRikujRoCe26+Of7NWrt+M7DsT4
xb54VqQ+cQ+/C/2WEvxjAHUUC6ESm0TgLcppteuWqwmjYTZWJiCYBXFaBK8rRdyV
0/KU7ydMcq8FWFH1m6PgBUjygxs9SyXOrdSvkqfXWKdelxjQv9TX0uMuUrdaDey4
+aJ0hBo4prGiQLL6p4wDcAaRHa9Ir6Z7hRGb8GvSejouAmcVuvz+EfKF4sbfkNpF
qr0BelCif27nGibpzN/UXt0gktVn9FCeZnGvCl/IdiCkDe003MXqozOOqkpRlFuF
pqsZ5G/NRCzgUOd1o/GANSQFk+ZsFGKkgecmO5unonsHtT+TMXALQuhcFQyvCZLs
J8pLN5c0uetIOjZIkLD3uNU4oQ6d5m+FLN8Nx6z0rqJQvybUU9AD0t9vrqgxo378
dAXj1/A5DaYli9JblBzSHMAKGq3sYLH5VG4cRjfw6RgtRhtjrByQbLQ9PfqCcZja
YHQRS/KBXoLB/9Fp07n1p2/+EwzTweG3Br2W2UpavS4HXHqMomKItZbRs0bl+KX4
Pv/pV2VDX/NcmckZJPzXkFYgmLD6OfYibKf+ByHXfO6xQu+6APPtQorrd2fox4KM
I98Jw+NI5SjSf85D+yM4SiT+4uDp8Ew/D/u2FNGuokxpIYc0vraPgP0LQl0Lf3FB
YcWgvdp+UPIe4o9SOpHoQzQVZSVt9pMk7Dq8SfMsLzJ1noJ5YWCQU/sUruvkjKrA
TD4O7CSjyU/mHER/S/cBLqmjogWeZ4zK67Tx1r0Djd82vKwkYVMH9k25UlIuFlst
AX8yfU7nKVGuyrv6cfyUrSTaDpxlD9wLQrrStOahxeTz4b+QtelsyfqO/xJ0HIO9
OiMcUSRIm38tIwlSJT2zdzoexlwzpfQk3tK73SRii6T58KkZNpyBYyouRRqzLVO7
FEVYH3d5j8sT5ryuTcyV3k3t56Dez3nCvQVwcuNwbqgaQ4xYk7GJqM1fCefx33B5
DnRuUWbYOvfU2mMKHEQOKrVAf5HBkl7mjF/rLhzJ3nhaeBtXxo69QEjzraVGQ/Nn
l3JCyCjbj0+8qgM4ugrnJ/qN2WCFk2+08X10E7b9PuL/Pu1w/LwVM96m2LCIgUwL
3u4jME6hq0I9uuS0JAskm4qcmt61F96DwYIf5JSEMCAtiLjpjUpyhegC4W32otes
Mm2LjlUS4LJsmOPEA6mx4W3V1EaVr2UPWAkRPKRARvW30FgLYU+bHMyU+kcYVpaz
JGsSdJ1vx3kPi11ROYAhPlRLBMVW47bTStD8I9NUbHKKALnHHCfCNUdoL2tNasgK
22IAlMTo8HDPE5XC8ediIRlptJUTEJxlcL0iWpCxpnlHfHzAR38l42Iie/KPqpDF
20xUwCLatl2vf4FsVB233YSxNUxLOMoisAQ/hpgybz/oQZD51tHqsz9A4YLJlbXv
mNYR86fy9+0kajECUtc0AQZO/JLqnx6fGowKwLYwuKamLEi601uZuEg6RmwgpBx+
e6f5whZpkC0TSNbP4A5mEzwCDJ4AWN+fn6Qk3hCzl5viNxvKQL0YZRU3FQSfO1pJ
XisBnL0xVgKZipqfCriD2CK3nVfwesctNrDQF3JlWqVvHm1ghh9eLjvuaXHJEOE9
YvJaJogd5ugwgzgbevAhY/mIAId3nW//J6OIXSRi136dl1drSgWpPVj7rqyqaBvq
sLX/D13I/vO3LotqksiqMf7fOYY/tr2GF/4Behhf9fQnpvnhZBFEUnVD8gnz6orW
Mnn7wIDhpjXdd9h+8Q2kR+46X1QhH1+ZKW/lBASJSPloJX7X4xQr6FcAZaXEazZR
MseQKanO8EJSpTjI/vBmcolYYf0wtTNo7ux3TADBhpa8RjcJZGBK+L4YnIqHvW2u
fffyiLV1HeFn3mqy/PiEymtmRXMKqp5g+eP1BUgvq+O1GQGtIwhKrapUpT8d07Ce
I+EXn2pytXCRFmX9yZDE6k6qu5pmd4zNufTmEoAxvwRVxYoDSqj8A1nN8ml5DvfI
/9c9hbsJ7PmK6jqgR1KZ70xK4j9oBHs9gvRjcIPlTO+b7eg1hrX5QbBI81RaPQ4Z
Va7iB+dBgIFGfYE2D7kKPHdgzOTSKMt60Xue2GckppAmxgAM6pDudjujr35ZaQ3G
e3FuqwkcvLRAqa51+xWBTbziPkA9JBBT3NIUF/4oeN0dioFYWOZknn75uSWG4lnY
PJGZdpSMACdzgz94BADMnlyTIHdKQR8TQVZlOjaShIxduxO4f2voydBgLb+w0MCL
jVfoEh8SLplxL2m95To7pGTFKC0qgFVFc3pg4riQILeO79uUHqCIxQOVCTb2x1zX
0gfR/LslAZdi39O9zJAh4TCv5WkAavtpWHdpa9mqxfU/GKTPIl9CXsMVC9LDkyot
RbLBb4osv2BQNnkM+nXGf4nMmQ2wKAiLhIOiq1yDwWK3epKae7R9sTJkl2fADGiD
gze3sudPbbtO05dNTA67LMF8kH0euP7Y3QAbtOXct5aEFEIh24GK+uqsT9ZKBruE
Dligzc5w0CY3WrgeazflKa2jMEtIpF77lwAvFMGxsWa7gR+w8cdG3DEOdtaJfu+Z
/mr/Oycn2YjPoxffPfPVWttBIRfl47t4RNv5ZdMNmBKZL8H7oEyaBpRVCDd9uIvy
8qbF0iMy0dBAzQ0voue+1cp0nXA8hs+1xSzwZp9bguEcMC7ktDwmPLIq4MMA4FJq
PlKpwJULbTTLQDyG3b6jGFG+LosXG5dWBz+JuS1xjaDc2NyYVSY76L4d/VY4X5RE
sN0ORGUT/PzdS7FIDLPVqc7sqsf2BaLnjAVRZAlM3owMucBN+OOs8mhZq5lOwhXO
iA8fEE3HM0mnpqfK3bbZa8Lip/gd/wo6tanQkVHiHfGfFZphcOBSRLHWx0LO+It4
f79P0xsUAUF311WEWYScRA9fzMQUOH+yKe+OqnGvEb0qE5JbTD/xIV0j1Jzm8iN/
jyDfXH+ABYTADvm8j2VRi7+tj0gHYPjC38szIgO+IrbnFuBNKR4ydzDYW3R7tSPi
6Bc5jQe4WGaeRDVT0F/Sg2vMEq2/sz0vLqId/mPZq1+MREPSKrLPJ+ClOeduavYV
Ta4HhEsxt9M/oRb4OleeO6feSqyZjkLmurfk6jYs+SwVVPikzUobFpm/cL/wSTGf
M0aBLtyTNsJHMhwm4BtyxyZBD8MzEd3rgfihIyTfg1tlhaUmcGeWCOLKAuxcm0p/
sg3JOayJtphtlPq6pn974N+Oi8W4w29WiTOGG/Wgitk5CrNM+NYapq3ixwtUSA6r
oFJp6mDXmA6JB14p8tuypbyKRtkUhOZazNbnHyvf18CN4SvHSM5VewlcYbfGZBSq
e2NhAa1t3W4g2/MtceV+cQACSges6WyeRUtA5bESpfC0TDEzlhqtB53Xm4TZx+SX
kOGQwLCbvWFLMwBNLiVcplDnYSkTlBUHQT5N4SqFpeNuhsyVpD9OLOeUAJR+cWzr
FHr5zG34PpcyKs05wNcLO3O0YDRF2Rtdy1YSqYeEjOt+znagJORX2RaDMLwPvNXd
zWLaJPypqmcfTVsobK5nn/cRzDh+bN4DX+VGdjNz8308xLtpB5DzwhX7HyuCoxug
zbdH3iZgSXfa8LjT9bUuOJUHoXClqwApw/RtbGLdl0W9y2s+YzSoYByr1O19sA8k
YHebdgzh+J3ed/QQIDGp0Cb0tr/BxBXcPREme1EY7XgI8H8vPAHB4Pinbu12BYwV
xhsC9uN0+bmUshQZ+O1JDzQQFaO34+6L0bF5K1Y4H/KRz53sf35QzkQvRGvVYTW9
SWioFoD7pl6AiSEo1vJqdIP03xb3o2pt3tmdqt2p/R1B2TeYRWft4rYcp1dRHOFb
pahOHaACAyOX3rvWse70tk3HSjwjIWxd249HDJdezhML4w0i5z1YVohV9FIHPd9f
H+ImvbsQm+VVpaAtpvBhsfYRSl4zBUTYz5715ZlBLAzyTsCAX4pDw9jKjDhfnG3f
rcrvlL8NW6slEqD1QdfWokCwNWfDHQYO/o6R/8h6hrBziHA03YGdduhC1wrKY07c
Y1PplxMScK+7GewGfTo9u6BbHYmuP9D1lkyT4S1luew9gWbu2iGrFlGMhYiOMoU4
ZyAj0w2WWAIu+Vjtc0oOOtXzsdOqhJpIMF6ikF98ZXIcxV+LFUGUbeYiGNmDG323
RzJloc5VaR3NFZUc2C9q7oBysFxbZbGqSpnzWMzUb+9mtaTtW5eIDJuFo7wbWcTb
ViqESyF9MsNd5sktShHo9SU3RsiKoH4KeaPLNLcu2CgKoZ2AgRAjhoXfOVwPEz5w
oJUGSVG+IfPxFdU191nMX3sFgomE75mMMSzoMNaa4WyfYVWmnm1ldgb/H9FkCvXT
3U4Dcb0SZCSr60IX1/oqJbEKImZ1MPyJXKe/SkpETcivknQV0JpkwGvj3piGHx8P
E3q9OpE+4hY3Ldp+tiweOTgIO26Fi8TsncavXScBz3tvQp4WzoJUNa/5mozS2V8S
90ZMue+MlTJk0vu/ur9HhIJY85zIODU9QgQ5ut9XwklOHmKz44a3GKd2CLxGmw2O
KGuMK4DcgFSv/HQrkr0taC++YFnugo5SzbwfiCE73zzglaFHOO0sJZR6Bp9x0uyt
IzKRMcHn7DU1Z7iix3NZyiGdVF/jC/nNDUjo01mWU50qH0bbElj32/TuJyvndGH1
Zc1k6lzXetBySdnu0t8kxh3xt2muwnVg9+sCpN2Hp+9F/MGROqLSJlClq/48BSQs
wOBNOqDvPttZu30OqSVTTkvFfh6nh/PCrVxmvqRKxZ/5B2Um1XBZRTEScgt7qMde
i/e2l6iMiuj/k93k95CHFpSN0ozm4Xe8MW8XAa8eVlVSydXNoVVB4DH2pQPqIlws
Lbo96Pxaw/CzFRVL+E7Vfv9nyrhQ3puAqqDFvW4YoChfNYcIHZaVFRVsduVYLalk
yEXd3D4gddcU96B/A2ehImXS8X5W/1DlRnrSpuE04G7xGNmxFLw8gC7h324lCEgQ
NpK/JV1VchcAnPIvR5G/tr/Jq0Nxa1E8VPjOeogQgr4aPqEHDsRlUVbVwrVQm+lA
K3yNa20ImkBWC8BedrqgmS+RioWFY0L8gkW8/1ex/jDVQ9wXi9li7opYxR6JFL4u
BmOuXeJYwW3PU96w6GeQbkVGWhj0QfQtf/OrNEPrzi5+7p+S68WhDmKfc5+GnWnR
ksNMui1LagXLCmjB9kNS+3uyQRDtbQWjab7K4AtzhF2n5asYWlh80y/kNOnT60oc
rpFUymXMZsGyc4sy7Nd243WaB+sDOIEqBn/qrE33LKE3Jv0D5YvdxUOpK1qJPH2H
tHyOAkgnCXQ2L53O/tNpY+sGD7vPxONbiYYyOoAbjWNArdjNj4UDKamWOYhIX2o2
2+KYQBE/JaW7nNEvA2zAGba1wa0VwhApFVsb0lu6s7o8SSCgS4viAHfXu0Q7lFtD
yWkgaGjOaol8qADwTJcIdBnWOX/QN4MJD1fInz2fojjCZvDsQrzmiX02sU6ahO8S
7wQGobMFJIR1LqnvkZi8jvAsnrz2g5wg9dAvj87OMStEkc88MJ86QcjsSAojYIlw
Qd+0qkHrNqHVbphfmuHBqNiBjT7GnWXt0p09AprdZD2bVxEjo9jvBBE4KTw+5hIp
74/c/okAy6/aYkD0g9t2xNkI46TE5H1Zn/fSlbxLjWoETw6rX1qrwOmB2GSSQ+ag
ECLLXjQxAlLAfdDAEGmCiM2rq8ixDXNkcAOy1QNTDKuc2PP7hGakUlHwNfiZNKgR
6bhDxrOxrZnQpdEESb5XG9DixzZMe9WXuVw1Bp6YK7YTx0agxQnEgE2Wa8TwxrsR
icEoCimQnN8/LY0kjyzOMGpQ2oZP6UZx2CS744X4ZYhPUde8do8UTr1h1bmz/FC4
k1IOZKJ8+eSlLpGKzwR4+iMRC9Rmlkd161SUy5VE7zvz2hc8RPbO9bSrA8/nuVGl
wNX54EpR30QdyzBn4555TKilEX4Vn2lDjQcbCBrMEtdOnRSftVkY93w8tS4uf8HA
SUCVJC9X1y5Yreb9ki4PjyG1YHBavQOM5rmL5u9UXhT/LCBfNOXzn8dXg68m+llA
s39ymU/MXzhd24Xx2nPR8L+l59inFsv5cKRX6B151OONkfqldtuRuQqpQw8I4Ktq
i6AnrkH2Vv+VjvUZxbKCGJJ18QK4YZvPTSBND+eSfM5f6FUwpRd6lz7Pgi38CGz0
JGoKJdQU1yco7K7j0zV2t5fW1Il5VJyn6iJxsgPmLD2a7zOAI+yrgdSLRO9cIcK1
g3MujP9J1WND/1gYdc1mo65/Daddk8fG5+RbiUId5Z55WnlF/w1ix6UP97bvsCr8
CrZGx2MtQaOcrhLWS3t1lzPhP5jC6FEEBBC77ItlxfRBIhE+3p/WN3K5g/K50JPi
3tOgF/wX4nnv8g409XgJaYrJprFNLfOA4huXvItyf07dw2D6DMjxuOO3y1RVUnEq
fZv7WGdKLFrjun/VcGJq/Sl2YxDrNUUaeC2lQSkZr/FA87dq9LhI6AZl0q0bBEIj
dNq1281p52l0MkbMpcZHYQSMAEnV6AJR0V7txJl/2gHha755J9A9yJJPKunlIiJR
8qiPJKH/sdDDnO8XgXQvPTmkvuuouCq2MO+7R0RKg32RJ0vSYOIN9rz0m0fXht/q
nU8xiA4yTDHp66WJ2HWIDW9lpoZJQ+OlINQxQV52Or2V1BqCvSU0QU3PN1MuCToi
HXjOXex/c+jem/RrCzRg15IpTdxNbcZL5yoNBrEIzcXW/a6Pyav4U2CGJZkKI75Z
CNcE98CEV4X6OOX+vWCAdZRcq0E60T0gbvLRsnkwlLDkpX8maWeiuFkQ1hjwuwx9
PdVtpWMbk60suGO0zyIsyrdzoXELB1z1rxJFvKDCPrHOxVOjshvEQFvUiOCPfXnF
m3SFZkVldwkczwI/eyrwrQszfS8RONCB5IqvqatJLdyEF7oDzbMdxbabrWqb6Bfi
eqlyQWXFupUPhhWRe2VzXNRS47rrrNrKxZhaZeOgiNo1WNTdnVC2AHXB0GB9gtj7
VPy72e1502okRxzyrRB254PoRKH+ZapwkvSmqxkqsEjPJ+HlIOzFU6KKM5S5HT5m
anUj9t7ygS9Iim7iHaiUpOZZUSWQFZQ0JE9Gp5nzd3QoZkGUmWjKpPRXNhnXdQ+T
a6u5JvlzFzdVRmgR9MSU9aLaV1+AyrlSTf6JySzTW54eljgUC+/j3Le7on0NZlXa
M2b72hdcaSYSHaYIefYC22M6jwnFV1+M1Y1i8A3dBt7cz3ku5rYB3RwuM/Gi0rkO
nw6LEnJjjZ7HkSpNQuQ8Ilqf4QIxMyjp/FXTpRaRcp43HN5rhTQJnCyNPwWjoJiv
JuEPzFKyQvZzXBCyr1wpIc9rs1fqdM/r9pARCqaV/IfzFHBvHUu3kratQvoo7eI5
tFeCKFioOXvJ9hebWhFKwec+bFnqIK0LzStRt+dPdFzqtijUPj1LSg+fWONsQSl3
JKBC6Hii7w5qOilL7usPxul1XCFfdTjeId1xVbNNgOYJMHYY4nuHiUclLyJ25MwU
KSEJJDXLrO1LzpMSWIGrMFDsJS+Y5eZAsgp6fAJ2PQsGoinROa7kj6gktQQYUFTJ
vBfmmAd12iGvfwKJJ/Edz2Wd1Z53ACLg++KeabWmBy9UBUj/rs2e38LYZAi86JuV
ps2pyNKvxvUANflUBdHKIoHOotc71cjtjBUbF3TNu3oFGrP2CsuPeMCifSpxUinZ
svWhhsdNCzyHJiU0vxmB5+uLV0EbwenCku9Six0mY7+CVhhudNgKT6tWAKyit6Dr
nWZkUmRiPLMzcnxSD5zW6Rvg50NKhSsF8m1hculi9zeQwkLALYCUA3zEQwaUVN9G
6owGc6UnLPf8/2MwmcPaWb+P8Pl07lokvuXSLpAEzv4HzZv0oL5DVOvWXcTSqmXM
aUmc4dGSyfNr6bjH4VKkPny2dKEAIe3Hde+Ph5mF6/2yljbowYkfRKEcIX1cmC88
0X7zDx4Ju+s1jLQgjYd8aIDBbGOp48eADruzOGblqAz8jaaMwmYaaMTLbPkNxpdy
HIGDW1TT7LlRX5Y9ZIA5+gu5Gme4gAv5WhTxD84sdIj//im2/0mQce1xNJHruCsf
FJGkMS/A/poi3pJnbHYwy4O9G6vhDD+Q7TsHW8oCanQqFtm0yWbbymyYAJkR3QQn
m0D90r8vKFtRc/1If5qmzQd+Q+72YGfG6xlzNfAoxjctDJuisX2XVJtWC+DeR0kt
g/FmcitamQwhboACg9ikpUS14YanljQ+xVp2aF2lUkJ/gTHpWHCtRUDAJb2Wot66
LUKVw6WVcIQFDor7ZX4UuXm9gPKqRY+1o9jLvO0wS3kGB6pWYSrUxPIE7HXsQsIb
ktALUsEQtwvoF71S3k4SGsmzdHuUvER6hKWXio+iY1Bk5eU8TZS9phwYkuJNVZDJ
RiH031dVq4/T8j/VK85BMwCSU4dtSGxAIWrf/pqlQ5s7nLRUyGGb3INE3mxL4gHU
w1FNTfLSpyU2xgqC5fhGA38G9Sv5hNNYFZ5zU81oeEUDTYU2hAl3nwOBgTPkCm4v
CNlAsL5iIHWK5SQlY5YCSdZPh9On2i8yzqFKmSsctKyHvx2iylxEl3l9hib45ypT
WsvijotfIu+2WdxXJGHFZi2G84JxQ1bktMPInDF2KAiPx9WpW334O9NKuwicmUNU
vXXCOwyKzuIw+6TXSsdZtj4Ug6HRDpcWNKtG7LucJ+5jSOlb2hO1g4mOTYCch1G4
p9UAoOs7Mxzm3MIbYDv14zp6v32TvBTOcixquPIsCOibQRUm/qB3iQGNL+9VMGzZ
2Oyrq4ugUEpbLP3t8T5FGxW4Sao8w/GRaH8WU65y5jeAXcHBTabVMd9wCB5xVsS4
hiIf2vlRDPXvizrP9DzILLbid2QI+jSZEASqnnYMLvQkU5ZtjQsDDtbeUPhYSyY6
Tvvizi0pmQzDSHRl4H6i9SyFb6xOaw/yVN105650XUKPTmH7cMqvG9oQA0bc74sD
J8aa6etTC2GDzfZgD9u2WmmInos+EfHVJINMYMbRUJQcvom6JZcGBQWhB62ynF/U
r7PrGfoYEgw0jXJ+93M2uRNgCNRHIPMHuH3VXi67J08ntaL1mHFDhDEix7cZrtEO
/GS2whMpcSuqOQTjDMdRw7lW65y6oKuz+wNC4O/U+n8glatyGkNOPSF0J4JxcaL6
WOA7ERQXkhK3mqim0lI8YEbxSWmjh2PUqj4AQBH46D1qCMV+q+UpZZcBzT9u/Nsk
5pZggrDK3lOPRxwDKVs0iP6YPGLOF64xKQvl3dzw6XpV8EnFvu3IlWi43tCE41oK
L559KoomhC7m+cIy8D73BmZ7ERfqypvBT00X+9lrnNkRbqwIdxsI68kDtZK/5Nab
lu37LdMGpstOgKq4z37IFjbcMYe17Mo71skorFeoqB/yiUdoOrpqMvlGLi2blsqR
NuQ/6maROH7e92HhOUPByOANb6YrfBkYj4LSLbBLNmNeb/E3v6OGI3FXBZn92O0y
lytM0TlqCYCb78IcJONckOl8sSUA9iGt8IhB76eHgPta4zWlSS8USSc5L9aYq5lJ
mOwTYrFbuUveyDSD3uW8rZJe+J77T/W0tDwobV+ipo664d840urEewb2tOjPwfgC
gJ1FR4ixGASHq77WYfjDJFZvkR1S3AUGqutzlo0PsMuZIPGPFUDwGNELFnhI/v+W
dmxlRiFW/8tLrv3Be8z5/Muq3kX4jqYM4PZFytTQcD8/qvsA5s8Pxq8kYy/k5XgY
AxuVD+XZkEdMBQ2F9049Pnk4Bvn8NYAyCOn5kHI9TdjgG6eyroypx63bHMCXV3CD
t/+6LfvvebdFBkti7Bh/ZRpsF/idQSIGu6gX+ba/IkzWFUN0Y5tVF+bb+gvGV0fd
jzCNR4i+0jppsn6O5Bc+baapyrUuD0GVFuy8vv4/H2d0DI6dKA2YVJZFWtQ+FhPh
OJxDtBU6wNAKrOEeMr88jvUz9clKpMEC8twQzwTuXyoy30Gr9n9UHD5wm8uGNphJ
EzpI9PYgy6zPW+atcT4Wp2X673XTijQOnjNPBgfna3aOMQrh1M3s3+umrTrqrjRn
Gd9JyAWOqcj3Qnz8IJyZXnhcUtTJzO2MNHNEnBfxlXND3nLP8PxPgWFCEqwG1AGB
QS30RNNjQnb791RFUKyDCEpLu+NS3v+A/AbdV60rYlM+1CH4F6t3VOPMH+VQJSUc
Of6Porj6xrTMc982c6Kio0Qxkh8frm7Xl68E4aJ8uaZEWCNXf17G9hGlbfHqw+bF
jaAaBy1pMkHigoW6Jf2GAV9oyNmr3yGYABF5ybMDRIXi6GesB5kp+MlKWO+RcmGf
C7Za/YzsKCLkIcvOYvsd1b1CqnsdZWuuU8DR3Mk7MeYiu/cx/6R5HDTwfVWGzrDM
ptM7B4nJyiMaswwiacUVJl5htjbHu1wrWkGaiQYwOrEXsrHbT3vnargAoQzNLqPD
Fs8wiXIMJe+HJOkzT1YgFZAwgAFWmVnIi9tR5Gm0c22gspZjbnQByrFPN5J1N5Rk
OxyNhRQ0vEjstNulXwsxkMFdnRm5/8KZlInho0VafnFySc8CFvB0U8C17vCZKz42
tlgNmTLUqpgCfgd+kH/RtSkawjUyTTS5wio8UN3eITtgj4uQwobYzc/XDbH8OpVL
VHq5I/Bs8gqM4L1BbsVRLvQlfzMq13QlhC9PisHTT6IzH0vlkqU293Bgzcf3HG00
nh6tySVrMqtjHnUO+OEFyDupm5ncjOrdQDVtUVq8RLsQeRC/c+oeTZdhAasLzJ4P
NMtq4edG2Hcrvnj4M/9mUr6e/Be/J9a7FotBRAnvAgBe/hvb5RZE6SrNK/45zbRe
TUokyWqcO0Uq+yfnZWN7XVc0UjuXJS6KDvmv0F+SEBc/5MNn/jAUZ82I4KBVzEl5
s1pd1qDNYDNB52Q6B9tHUHzTaF6cOo+TJuKtVLW7RgKQvNbte2V3iA5h9gKVzpmk
JIsdnWF6Big2t4cPUK3GZke1ICI3B2mc2os0zprA2uhh8b94NZlpSP1FOjIQqJdN
iqbRPbe6cdDVcFk8wIUr8zGiqsa4wJ9JqQW78XeJE3025dxerzKYm16lIH+l06PA
eg6Nz5hbyya2Y55DwbN8AmARyjgXxj3n02+PDqYDyfDM0b7/uQ1upbgQQzWJeIMQ
aKHatzJlW7jJ9f9hy9J21qOM61sDBcn1KEfwKfUQ9vc9yDFaexupLu6EiYuGXmHF
svtG1M6+22oupUC7e4CTUA4Y7LVDDIWvVr+I8Q72AfRdfa4nvSLaWe6wN0zGfUAR
yXHHcfa96H+qr+Rv/0WeRseAItxPBcX8VTVEJbsMVjtDqeM4Ehna2hfgJABTZlO7
R2ZUdyU49JgrJs6jQFVU61dP8tNL2Z64Ji2wYA8Ws15WI2qdSgSzhALRkGT9VKI0
p9Wn/iPRQqkVjW2g4STTIaeVi8bV6ChR1z7h9GtE0zKd37+XAjJXljV4tPc/YHba
ESWhGI/2/kZ/B/jHnflUl4S3ISSKJ6p6zN9amYh5aXp0j0A44EKn/hyazImquK1y
tEOIlAMI2X0TQPvJ9upoiTxNFwf18HnzFZv1p7b3sAqT/8IZfrk2CjpD2haOFRvj
H+fs1qAVqVxTb/cDj1gU/HBicMeVLxBEZTQb/7oHFvmUi+UIEUuzK9J+MFtDAVc8
7SwKnUfsgh/iKM8LBuRqL7fqRPu4iEDjmlc4eRAR/pijrpDYQqfnKPWYmmlFWW0Z
vqwaKKvpnwm9wWWr2rZQqB/J3Sx1lpptYn4nLiC+jqjdA/vhiR0gaVB/E7VftGax
9GZMNoYWBG+UnAgcSP4Uygt2Oy4CJdZYR4rggQBLqLqzotxqdEP9Zhys5h7LQxNc
IVPvOTOCqT5wfEWvE12aRgnk6rN+pAmaGXzDEXC5xWtZCp2nykCLt5XEPt9Fv3Mz
T76mbVwEyDCQx+2SEj9YSzm+AVJRs9Odeo0MSDDVe+Bb/NN993o7p3Xkm1ng4/0n
kbK1+6O9edRWkhszYfo3pG7FHQV+rC/XqafYXqyMxEJUN8nzgxLN0J0zT1a8qaWI
2mKV5k0PUHkmwAsOcBRhXdeKOiPt5Oacokgq8HaXPeYRpJV4XZnBmXo16I8ae+P0
FEkfl00/RIvjGNDXW6RiUNNynyRLiXRf8x9X/+b8VzekBGAcAYdZBMlhafYhdMbo
rUn96GQCtimjhzYo7ctV0Dw70Vsfg0BRZnHFa24f6D0HgKLEW4/PTiez9uXqMx+y
JVfTGCNvAa6Jsb/Sr5jo81JOVuHSxYgJQomDtmY3EZZVeWC9+viqWVUmIgSnRftE
q58Ry79WJu1XF4z+aZkGod0VuZ8YecG4tN1wGRVgyJjAYvHzs/BWBu6vtrJgziol
7as6CtepeW9PVknqA+38hPjiOI4NjoKgmTiym1FQJSGmJsQ5tI15cXJsww07LP/q
LdJW1V4d206x6vkwUrF5M2JJsh8eDKhl2n8S1VOGkOriMIb+Xk9knXDrdgZ90ce7
ai51uOZKrVid7qDqFFVXXRsrYtjBcfBznp6s5ZBHfExVij4OsUiRmYWBvRu/5lE9
t0uhayCij+hdmPHYbNHs5xamBPi46q/Z1cwJkGRIaibIA52q2Tk+gXWPt695U8MW
vbuDggrmqfV0PgzbUBz93cbCTVtH+d1tNyxagqmZVSPZ+09b6GGg1GOkBkhbMPJb
5NsuuB//AKuLNoeyAyQsp8ml8sybDfKXxd2k1jnHhBMam4akprJX7yimuL+GtYyV
6cE5F653OXd0d4siY5WzRgCFEiF4gPtaJyWMnNI8760HhHpwsGymsKL+BMeocjdb
n+nRMQzGeh8aL7xsK6pTuJpjKOvhkvNJ+OOAEzVoMEGDIG7ZfKuS0x33GDsDvfGn
JMJ8Ho3DvDS3isd/jLu9Gt8Hv5kyEdaY6+8n6r6Ip20VsmQn7qNEEeRR+0vh1q3Z
fR0uGWRQCgzU/nc9BGUvzVemq5iEhXfvSIu1YxUCKEl8M6624tKmuHC/Yku7Q2Ti
EkFaTzFhFe1LlSUaDTEJvXXVKppit8xaoelV7zk1bnRA4fLFfKTGAuHLXMNsffbq
8G1xaZ7+f3gisHqQW0xJkfbWHR+k6vc21ewhSOWe+xQ2mBysxA9NJIkAoo+ZHJRP
J1Szt4gDOCYmngyBbX6MOaUc0RVTcRvTV7cculdVIx9rt9+Z6+gqw+z/ERbZigLX
o+NdUm8YiAwS3oyptfi8cjStvrHqrlixy0TS8zExAb2sDQPKMibzp+qn7QhTRPGp
bgKwurBzkUxjQnK6BcnFBRPjZfXLkuUKa8E6/tXYixdiU+SjVASnq5QY0iCJJn7l
i3fOqK8Vh1PkIaRDTeSSNk4rTKQbMug0ns9QSpBPJe8iqFK8y+ncpotYwATEvr5w
HTziOuul4Ot/v2nM3FImegC/dRsag4wEhKN2VWIMI6MjfjMmPeIGIrFHkFU/2psQ
l/q/iylc9ppByXdi6/TRToax8WXTHsfcn8XzR5FZuPb376Z4afoOSbbFt2Bchc8I
MAY4uMPxYuXRZ92mgQpyXAmod94jK0y4C9H9bMOatEFFILrCD11EXIdT2Ozu3nR5
UzrJb4GbI2uSi5zuL2maMnwrX0VdlzYYg1rFMFjrCB9F1vo8kC33jpzPB/gxDiTc
DanOYpCxs1z3F03eN9rbBh8bjadLHwjPNX8uYnYzf1A1uSbZr6VPyedzVfwrCy9f
zu6n9rmHsoaRwT23fe26MyWOMlyjxfKgWcgx0pJYtOvn7bhs7L8MaEGcLgZSsPjL
rxHPRUmaIEaCBgYObospa+aWwFpHs5JU1HcNmIiCigVpKnFnbzEDA9Aa8Ted5Ycg
MsxLxXk+yZJxCtqBXA518kk2R2Pbs9ojlS144NCRLiAkC7Xhrf/Vw0JHFiyi9m2v
RGsWJnUSKCg1QmIzM1HKWsvfxDsWvT/oh0FHVagztgfD4hT2NTsPfnzRr79K9kCX
/1D47nMXegLOVcOIRWzH/njoIDsWDMOQppOgguA2JvRUBOjTXaiC/KRGpXESXJjt
ufftlFX82AOoJsCwGzcfV3/yLDvmZ8INvhb9gQl9Aliq5Q7SL6Tdzy5TWLUXiezH
Y0baew2pCCuejw12AtcvFPzmr2EV1/Mf/WgfH7p85QGQar4YB1pbPV2ZnwgTLCXj
7DlrtGGHs1ijo7HZT78hw9rMt/cOS0tExMCzEbPHjK1ixM5ThZDcXCHgSQ8j7KAP
PWOebiMf3Tlqotu+nzTRb5s9cqWczXmV34jDMGVUOBMfTvX0gkHSXk7zO02lghc+
cQ3eSkVxmKqwJ53OSOu0ZnaFHR7r8rlcXrNGm3Gv45DDoBu7uI0oL+5WKLHtHUou
vzSWwpumw+JSahgziX7lxRxFYihrmjunK9nx4SY/uCrKHxdqEPPCgktpHj3iSrPZ
KD0em/VGm8FrknN4z7idRs59GHFfjZRDqPd5sww+iXHlE3o4iXU9yhlNRWirKe/g
zu4LqFPOC2gR8qgXUynQPwm/4VWZc5NCeo8FI2Tv6djLUD3RpgzwVhQvvlLQRTMS
vfMdS81KRb82GOY+VCAosqvD4QD/cEBz+UeL4szljDfM+hUMQ9o5UBKgdVObXmLD
c24aWXzzlA009BUoliKN4gr3hy1GsQz7Gvdg9/G0IjNoyRNFhNxKoyfGu++vhfbb
6mGLH9VtsULQADBZwIywTpPxaY+RmpizDaHKamD186bvqpR7NhRjlH/lEsxigK/4
kVFFQyUmP9+giEqw5h/3CfCTACiCi+YFL8CliTGfdrILGls9aedmP2+5WjoN8DEa
lFcOiWv196bZJSTxLhbN9iyky+xisc6G8a2lnHYZXuA/QzMpYiMFUoCugFZ2uMBY
7LTxSaz9k45AoiDLvroOq41OxfEA+/MVdhqIg7km9qzUVg+NdsqdcAl5WY4ofavq
PzqXv5MSzdyKJAUawIcltWJ11r5pFGvzad9SaKgcVJTzpdxSk8JEPABbBMa348xi
9U/4m8sLYTtKACSm+7KyuIiYMxkVNyK/aCZUle+hjdQ/OIjBiwXg1O6JgpJKnRjn
N13KHA3czKLinwO1aRJIV4TUXPA2vbokO3BCQYF/+jj7z39d2TqjLtZEFLu/TEPR
TlZVB0Rxtz3v9RfHcmSYu6YSct93HOWg4zUwSLSDjuCVe1bBQMHiGzeXcPzVmikQ
jsxMrFeNA1msrW/MSdXlyG6255k8ghHj/rX4VSQTMrNJwxX+g2sLOax1IiWQFDho
L/XEnoLRu8UYeaoFtI7QAX2IHgQaYm/55GqYbQnsi6tS2aEL6R30uklOE3nDpDKT
iMA4joAm4g8PMwJge4eb0zsVOwM0jZDKAmO3/QIcTQmJxP3WoQKancVa99qazBqk
Ufp1xvzYEVHR4qmSLuDNVZqyMM5EmIOL2U+Jc6HJ6+BzXMCCn34wINz3RBDFvUqm
J/hVQggDudMAbzRn7LALMK5yUpgmhe17mKcRJPIAjOVrgluea85mwTh5279lTGiG
Krz3X4EJD1Pn1jsH8WfwaAyEGZQug2UIXt6FQTsg/LP8TPr/BY/8K2JwZk3roKqf
JHu44THP1wyEE9IXjjVRCC/ZN/sJA5e6QEwS0i4xlTwIH8xS6J38Nzbw6SpZDW4d
/Bp4iNxj5pUBYmxEmPHJ0sZBjBCQSNiy6iozEik/TcnNjLHbKRBPzfEJqYhi/q1S
xd4MzNXAILVipHaRAmm9E0YWvQJJfeXs2DB3run0lB0EQZq9NkTFqFGlLhpgfSRR
z5BtXcx1H9G174XROMV5IGJzvYC7FlD9IYcPLf3fjzVGCjbzrw4okaZtl2kOPAQw
li+OCveANFfFIzQmr1PhsueZ2RhmN48mdUrT1orP/s6IiaZS0ef7ZGkkw/cQHkP4
Xmyx4HVcOnJFTgjFbXGA91W3NkE+9ROvEuQx9MwYZxitECwDvUleKdqERq7Sv8gx
cdsbIS7znPlcWv+mzr6hm/IrgWXtTTjPEA+ljWgbuAUHkEfj4e+QCcMaU9k8/yh7
ZYDNU0Xm8vyjdpysNtQzKHqkRgjg2+ltQ5KxdVHVQSlRelOGEMN9a5oERMipWq9N
VfV6z2LIzkE16DEIHSb6hhrbKL/8ua+UwmaOGMSq4SerLQwpBojgPIQlWKg2x5jO
C4MEG9nK728TEe+vNkL+mKvD69kqFeO1gC/djnPzNfkDLBngcSYs9wS4jFPrOlbA
BTZc1/mALknL8gEF2VCXZtOLoir56scH/zK5IvKBtqs5CL78G33LLUSeFrexob5D
WNqnSXlO+njNp6/akAoyE+edJVFQ2zl8lKTpLYIZzcqSB10ZAQuozlmtIL1OG1HQ
8DZb/lsZQK5cZNLNb1gM98tmJ4L3iZrwKZqfe+NPPoSN8wBx8uaW9eBRQb5df5nd
prZsBbEBZ3f8Gl0nF6qrZggUvEzno4Bj7L2zanVENIovXRwPH8RTMF1wPizo4szy
dsFF+d70onsCLYnP/2K+7CSyHk6mzV84k4CrTxzHBLqLbDMrgZ+WX32Cg/6Kx6Tu
GEduf/z+KZCwgj2aK7OluIP4debLlhgh2TASG6r05xkLAsLvsRYmDUfpegssBkSX
XXpc4qkA+hEU39N/V/VGNKcYmXjFIeDNOp/zvFwJXcM2nAvfxLi1B5IBJAx+XLUK
oU+yA1WKG9IGWceJFAC7G6d7uHayGhQilHfYIkmOvGWAjs63bBpOrArAFPLsfFue
ZNfVIwnHsbH0niopO6UKnXGqXmvAs08zoXXJBgzjjis4tN6VGV+5CTGZlRxBHrqH
VV/7yU9YDSo41n0Lgug35DPWhYEyfIm8b0luOfUrOOdvOhbk4o4gNS7/nm/Ik0yM
LfnYcEn2lG7/9XMQHj2wfXhFK2gm7SDr7fdk+jIkJ7YTj+39G1Spu94DN/r5siw+
HpsxdzoiuoJIzDna5cmWSuBSFkX+7RZZHECT3sdFlhOnW1fyobViUWLz6oPRvHv1
c6CAhI2q7LF7G7gRojRm7kkmpS8WqcdEXvlARYRXILmy1XcTVgkfdraPpOU4kK7+
VZf6YwN5gQl1O4rg5VPEgxdWvs+MqlXvabwgBHJYnonvyrnTrsvpLmSjrV4STryk
RlTAXAeSTHj7KHTeElYSWQwT3XUygCKsz47qxAPMGn28k4uyjNF0BE7TTtciLFJY
3MwfutmKgQLN1yqy1Yl1/h5BBL54WVqpO62/vp3ep2GeK7mzuts8NVifQ29zqilP
eECZMD6IRaNO67bvZ8epFLh6kfClHuwaUsUI03fZTKofBWUa8rLJ4YY/zdmlxrKG
IOZFejr8mHfQ7pbMI6UNrKaVOWKiCvptJrlt35LDCkBKR6TcFQnEUHWf3rAtkGzH
xNYDUqBnYlopylADVDKj5Ar0FGMTdZoJ8wTijXeYi1GVc6rvhY/tHzI7Mk6eb+IE
5L5SQXo7Dx2ZI8ZgoE72jYih/v2msCneIXfbo2Wu7GLJKr9Vc/nIepRM4mEQRhSe
uwj1IQtks/iqeD4AnL9XSnkJY9t2ue8kl4VQCGgR585BDSzOT61qQDqVfkiSmf2W
1FXj4CIGsVIy4OC+qtATBlmTKMh5cCyXZ863mneMZQ3uOibjphJZqAHaJcbq3HQD
YlzBurICqGpuL5YUOEsQJpnm352EGQ/1QS4YIX177mpfPbZ0bOCRXhqmnCAHQJ9s
Sp9N9g07AQrZSr2l6FxWU/s5BcxbBfDKDjgT+3zXCrzcpP6LTB9BgnAB3UmXjijU
0uil6CUhwyrDuQMM8ukS6+e4KpmQeX21+dw/Q/DtURp6tENMi3e5yB/22RHK2Ujw
H5SWzdz4KwzVfff6OE8iSKfaT5bgzSTcrYwZhNhLrPmyf7pVxIN5h9IodKPouuOn
ZxLdSH1uSdBbO9qKcpF9aYZT2HmMfNnql0fcuij8CaggYOYchtsd7/b58XHmxzay
UE/G7qc4hvp9u8CzgyzX9pYMCxUs0FVR9MQYCZL0/n+/b4TOlwUSbI+yW61uWpJl
/zE7HF8Vzd+c34QkVf/SeElWZZlDbBPO4Jr/nqUXHS79bO3HwpW5qBU6ySVy2xD4
S5IMpdaz3DYNPLCPqvTfIBGiuoERpsUcZRrvqFlyKlZohaCV9xmCdwaXkwtXfsec
enoqwMG0LTXQTbbBZ5xi6TfzY+qXedPaE3K8R6VA3lOo/Iy5xySFKyKgEf1aJsQm
O0hzjYn1F4VUqSx+TOVvl0uzn9hTutGPalsC6mNKcCmwj853upZyiV5txAqG1tpd
A8VkPJFRg26FhnSSxY+Qk/xlVE0Pzsrqgu7obQ8js9QekIYe51CfI7lEDDc8Xlql
kyoVgXV342A3lgDLwyxnyFx0cUnMeqxIDkKUkMWopCiy0wfhLevR1xFqYJ5CQI9e
m8SCvC68OngZbEWoGBznFqR9X8PhW+w142Vhx4kG3OZ+QeM1RzfMHvhXhW9OMq2j
XhPzVNCUsvT4IyziHv789tM/Q5upkg+byT4Svo9xZZxZTR8EmksPd47T6/gZaIo2
skPNWDfCRburVvLcoBZ5j1r31xfim7aQCNx9KvIRQm7aJhaSmNJLz8AxXRpQXC+5
KfHC+7UU8H0r4KwGjcv0WjX0k6/gQaDY81Ooo34Dr9cGZjGqJEx5tWWzEm3uBeJ5
jRktTvS/Ldl3ycDddq7diFqADbO0HL95EmcV0W1VAc0cOshQI4RqiHY6qt1Dpzz1
aiyyRxDewzAAar4pqGQE8dKGgoo4E3WmTKgP+vKATPfM5ArcUOhGlI3MyS1sPOnM
GJRC8qqlYH4ouJSKZVHIub2qHkomKE82zYVdMx2354P5jgtLDJjfPA9V4aaL9tWh
nhObv3LN4EP3n4jur1WS2jeIgXEUAz8OXdAs05S0U9RBt5RHMRoub8nq9KVnGp1c
GZG177xFVR94wlLq3QOeiNun+JqiLZg74EoCh4Eic5uEFoc/IRea44+g3ku79FkM
I2c7usGgO1ovGHXZo4tkJjNf9Z7pcOKDGlxWCNHbx/+t4gjWYX4FppzTzOFG56V9
7n5XFlhZwH0yE9UlVSE4uCcJBkU2+/WqD3LIcpSvWrlfdQPbwy6p2/lqqbLPpFQr
HTbcfWhnvcnRdbBI/N5/ZZLVJZwgqvu8kB0e5qJkSdBBPyt1UEZS371l2GIsW8Ob
eDUyztisj9T5xJcLcBNgyKDc0mt6ygB9Bo/6msf0wJ92q8XlvoXeOBQqyb8YLa1V
I8FIx8lzhh/2XU7ZjQX+a3ZB1PNXyTJMp0aJ185fqgJ31I3wHviz6scc+qp3CmRj
ml5kSaNC9Kzw15Zqna1D538/hrcdGM8QT+siwzC0X04bGT0phqAJKd+ROgeOSWsR
0cc7teqI33SZcEolIz6APTkEgz2QSC/sSBa8CHuX1HdU6x6a2swt75GKmfQMh3h8
PmowP+QmIfXj9LM987meI/V7SOGTfQBK9crmmon36gsjQfG5s/BTH7TovXd1PYJP
iQStzQbhZCHgauSIdWs/rkh3GQtXHUVenZi0Ae2Dwopmw9wj8XWN8FJ9fB7napf4
CmW7Epb3IYoBVTSMVR++u9TiUJfQJwFA1H2DM87ySekvenUD3nijHEHo0iafwJXK
xEk5+JsimSaXL5tmG/HHv+s/j331JO9Dt6RSLvCHPu19DMyPrc0r12VSO/0YoE32
y5U0fqNg1VUNzi6wV5+H5OrpRW/OcJqnFnFUyqhKUJK7ylLUow3oI6lG6heClb2t
nv3OAKvnhywwP+Fqs7NvNfz1ts8xx7opImd/LTaGrJxe+lqr8u86nhnVYjTQ5R0q
TljdHEeyznp3MjT8QjKNeDZ9AbpZ3p5+0L2W5uUl1Vu6OEdF7zSIZhHQYl2yOQUC
h02FNry8BKk5hK4mOGOM/E1P98vxHEXOfY6j1Vi4Ow+nwCuQXG9p/6GbE1ycBL+F
dQ7z0RmULk14RVP8qEUe2bbRWNGSisxOl2MbWRvUIk5XGmkymvRyHqG9kPimZHKb
nhZscpIV+D9Rho7Hb3Oa/t/0ziSh01nCuaz39HIPHTyMrstUT/jQl4I9RcDYPRbW
Fy4mPXsHfFahPHyocaqZL3qCyT8QM242zqOckQ+ZSXSRMlp07zidc76ib9VYPOcF
lKQKUpLNLPnmwgZzhDd21cVqHyDrh2FVlY2N/R7MvgyOlzz7gidhyCBH6rAlZHub
aQSgxrbj11kQm/IupKLpq+HnkWXSjA3PmDfZm4uTKyNGYk62MC8UPKDO/UT5dEMa
QjzRpJEf5u7Z2L9PuhqV5nvWUHAq2Bay1hQg/plPKv1Gk9W+etfWipEaa5uxxHYB
ba8KQi3sR8fOO9YiNWvrJJUwvtTXIe82Yab0BuWsh6K/rHtCrQeW5+ntimq3xo8j
T7E06FIGVxq5ok2s7LxbbJMdI/4cMRzjCqB16jcRY+qYfb1PTLL28l7twdze4/P3
b0pUpl818cjbkeystepMN+gzPM6qzvNmE9YHqcJ06mc4PRz4e4nCDhl4jL2PB5Lv
a4pntpXGQH1uhH/n8j3WYGLX/GtAPuqgAbq6EwpOzECWd6uIskUiEBCVXOID8gRA
yd+jvHGdVrjnQxuYWmIPW5kbu0+gGRt1HcyH7P51sGBEUO5ehziL+2NdPzxXjYeh
ruOiJivBijaYKFZWVvtSxbFYqEb4MslGsaCdzkKAqypUewhjj5ljdlIt0Y/9KINx
3Yjl3mOCQ7TXgyOvjUs+XUOywdq1rBEH3j1cVF0SzbkkStd6Vztt2pv1CuUlHpS6
ZWhX+bD9v7WYjzxPRG07Fv9nEOxDo+BMVXv2snlVlQ4OqvWzDAfBOvwJ8jH+e3Cr
BJdEII/54orsIqps++g2SC9IBxYy7W4/LDckntLATXurL/sjdvts4XBTw7qpL6Ow
SZ7rY/iPAinLWJ3/7Ty6UO99/7pJl2aexbtimgQXFqFIxQ3ruN0bqsHcejXEH8lA
Du2x1Hz2y6Q1XMj/1DXOPoPVZW1Pren1NrXvR5KuUw49reoTMpqpOHu4M1XkH2oc
Qh7YG0b0SuaCDGKmYUdq49Tb9dfFeGmUcMrLkbbxsGGjtw9eU+fz9nQFH8C9zCqc
aHRFgTLWEFTBoAHKLnDmym3I0SgvMFr3YociEm9dcZxkstml0dWZ46VBbUSGbCUs
6YO1Dwy61RqJe9jZvN63HS9U+nrut5TwWXA5oX//SpzewPz6iqCIp97kz2KygVHU
Xb+fbC38sAh/GBhtrcQ4EgIVWuV0H4u+Jo9iTsp2Mb9jS+rmDORNQAFzwO5+p2Ld
MrmR0qHIqYvYOxA09r80aieGPe4yd0ZjBigaP8o4hQ6je9yyOFEFWkmt57fG2VCP
7GfpMVtjbeXSC9eZdQ4WajlChm7jvtIyxJruW6GRKHdH8mKzc+y9ypZlq16eU06C
bH4146dR2GA0EdKJuCObFQwnZtlndzkL/okg5jLqaetzzhtPpBOytRtho1dnbYS7
fkluQGjeQOmjYkLdNMmtNqYaHk9epWA1C+s4qQ4ijyQwvtB7bTJpNqZMq4muNxby
G+31FONMnjQYMfKuOYuCIoNHR5+7qi8RM55RiMzk+xEAEBWCQWJQRD/XeX/6jAz4
QoTzWVC9dz7uWCyoV/6u/uFxwlxOT8M4oTfFY7wudLvOamZJ7SttOqUQmL5mbrQo
7ZiDMjFHruEjfJVbmMAozgyKyrwSgQBc7aDM5zIUQStF5afDspvtDRIDuKrI7iws
lnW+6hmA+CIO3QFSC+p+TsElNCcFpZb3iki87mRGR0LTU8yuJLSKK+6Hbh72nnhK
zIHaI0Py0q9bkbc4OL29VpT1H6ep2QHeP9Jf0l2k0jmk17QglGezdzf1d0ZqETw4
0h7X/BiVtXRfMX6U2npP2FN0FZ0j+rMHbjXKhad/PghxjwGXHRDhykfBLbCgxB1F
FIZuLeocNNfST9YHv9nJxStDD4dGmi2as2QS2azeti5JBCB0IzJjyjM8yCMcEM5V
QIfI3pPKhuYnSX6WBdfN43hgoRH07TCKYnhee/yLzgEY8hKeCtDkcN6PoPH1xPzi
A3tTrv/r6rPP1TBP3PxUGy1biC2EBCeGs40AHbx/P5sSTqLmitOIymS6CfgYF3zm
QWdG4d+Jg/h3Iwq0hD2TgC6SaaDHGs+aomjFpGvbK6Rmb8f9+Wr80A2M6lR6YAG4
tSkWV8WhlTdqmUaJtlG7sVfBXG+xusIxwb8AehKq6bkiIrLqS+CEFOB4trcuFBjQ
+GKSYDWoR7nFpqSQQMOnFhKHZyYBKtOwcmyrj+bRApoZ+j6E8TGJX/8NlRlvuc1R
RCd2rtSb800VX+IpV3c+lFB8bpGSIcW0mCjfzRwRueAE2UWvGxF9+my4HZoR/Vxf
x8U6is47PV2EqnvXPYwu5IB2HAXFUDfwNlgbJuLn5QgHcO0qa+2HQq49nZvo6UQK
Uz0X9eLW+/3fdnADGuiIG6SR83GG/6MRhkqOWVOyM1LXL7/Ald9cMMjOomrIS7m2
i4HBuzz9teQivhG4KrIDkJF+3hJeuE3Qn2FUBvEjYoKhndXvqzO72AyyQN6s1JGg
PvmoO9PFxzUULTeouIBRDXNf4303JBTxhShmW+jkxx75Ck44iBvr4bg32NzewxCk
6eqrELPSkWddJMtK7CBBD42AdISV++uPxcraXOEQZ1JNwjfHoReol2i2C2sJ/s1i
OPhDSQ99ff7eqt3lNHPJRLlui8wsrbzY2HLQTLSFkwb3k19m3Wx2V3f9SN3QzqQX
h9/Mf2Yf0J4NMmRJ+Rm+X4d6TSaqDnFBt8ujUqlSUwLwDN/4WgTiA/6H8tex2Qv7
q7lkVK9vegVKGaxMfUzWRpWXWgaaShwAQvEuNyNZIRzwOQO6RTRRaoKhDl8VWfwm
0spLx3qGPr9kuusPl5+40qrF4KzIJxIOxJTPWolvOUACxtqd2+3Z+1smcKEpiJLM
Pe/K3DaS/vrq5Z6MDFl574Ham8zT+62xvsjgK4BBl2gJsaGTROcjH2/TyFs1XlGr
RzTvJgVZKoM4JxQnska6RCdV1VAShZPBPUJSsX23eBl6Z4TW1hWDTFzJ6n2xLx/5
L1WFtfgViGXFgtmWg193T/aCuc/X9LpUYr5G9uDxi0e14EXHUC0n40eMp/dd1hXX
on23vjZohSvA7f4YljlUCJbo/jz4phf4BI1YBeZxdzF57qmg14i/p/+jqlD8O7j+
XZXdfWQ8juxcYDvPAefmO8tPIa0xtNTRaXYTIvlbIVwmW4K8QxoTDwOQqbPtVfIH
u0lydqC8XFqekYp/g1kU+bV73bcWmfF5jGvsGpNTrQ8HVD1MUgXIWSCT1yLnceo6
swQgBzvuOSbzT32d7TqRmKYJeSl/7zVS/TzujkXZB99JA4+KJuOh32xMi4U6I2qJ
XY/PgVv6c7MOHwrnVAQkGoFaxmlgeraSGkS+5Vyz+yeXMlKukMmEFq/OrUT2lgSI
7OlyfdMUgfNe/eJPki1ymG8nuJnAluqdk/H+kb5UDpHcEax0WIBYG5YDISAGdw9T
Atezu7jP/aJXaBu/40mW7H0zp/lHThqanDdVO7BNS7chpQuhXFMurXU0WZQDsn1/
MDQsZ2N1qIBYHEnDInSUXXlIQvdf6DcEFR+fCNr/al8ZeGK65H/QgXW5jY42QuuZ
nel6+L9dElhrKOHUA/Qbxz9bpIlc4QXMp56aIeFXdJNYZnQmO9Kh73R0h3KmTgIW
hTC5tlq9yqtaYCQQ1R7f9/lyZEYjtqEVdrCACbNIRKrlwwPEG3IOlaX29IAjD0rG
fSg1MpEz00bdL3L5TU7i1zqeAfVtyaG3xLWhumCEXa10MivF4gZPmosU7fqRo6Dm
MPg1JimpqAZiW8NXqEyzYE8ko3AeSqcsoPeOHBCMtEhvbKoLFyNNG42aNFDW/VWE
ibELFaN3+RIvo8mGcwAj9GDhas4QolG9WKozwNb7VVMZovkCBBdiVpEsCjHo3S6r
jXAqUGNM9GVzz4Vp0gzol88PLCpNlhCTeYrFNwFXhgC/3g4PhxAWncKs4OGwMQp2
k5Q0/5eqTGUJ35Dco7OQpPl/kdo+dAsSS671GimB16F4TGmkjc2PT6XX92OSyAqS
wXo73HCtMjutAxEVYQj/d1THy6V+HXa4pgLshjAKxb+tXrkyEgy4cMG+vHgjdIvb
JnuWdg7JFhugenq+bgQwbVXs9UyUqWObbyhTbwnU3dh7JMU1+OyPCUD8w3IknkKq
twVzoDU6UarkM57XdjviqCvIz5FzgQAhn4j69gQQJ9F/wCwp+0oqV8e86kTLExXd
MeXDefKI0OfMtyK7B6qGaLhGQlP8krCf0Pm03ZtPSQYAvbgGshmgm67LWAKnPfmV
l0lwoXQBm7eqGBSN+dcgU68aDdtwPLIoUYyx+f5xwUUPb5vxjLsCzFwlIsM86Hu1
3bsg/57i59wjz8FwyXxOfqXBu+qgDsauKxb6bitytUdI6qOTm4VrC5SLAhHX4TVL
izMMzhZTpTF3uT6OW4itDwbDRJgriy+IOWbfsPTYZ1iBOA7RvbB/JZ6erY7xqFeY
Xttr+lTpMYxrXZ64tfMIizJykRdQgg5Kt+Tw4AcxQvxQ4P+yGu9YsWTXkuLpK9sw
Dcy2Cv56jcpTEhpoQ/2ZNwO5YhLfpsqzQor6u7dbDYrm8p64inuwNcBirdLwT8Qu
9p6npbr4THZBSVqXzilaYtGjHH7c7LFHHAzk3n6oZ16PLFxzTMiSPbD3j3FAhNZz
3rg0lmUfDLYH0s0ZYqjcJdlrn/MYF9qB7jwaJmJYcPtbZcnE2ZF2M61qhngWcTWC
Yh3PNZIIrN59Fd35cGTmiQn6j1Z36JTAkbNne3n6OmGhC2A8lmmEbnHahPg66WO8
18R8aykfStsD8yVWQxIg3tVv0NT7B/6e6spOSKhvBWKLLt/IDDmAYOnIRAKQl8TO
e6AlRlDaoY8lzRfBRRmbApqZEamK8lKZFgzaj1L+c5KYq2C7HaYShuj573msOQ2T
o6r+x2GfzJ/AtsbUBqpNSlyNQtm3a2fZYjHSl8QUCYA0QoiyoElwikFsE0khsaeq
nwJ6+fgrsajD+NJDNqZpPbZQTz4dOYXaEiIiUk9g0Ajvu+BaB1sy3GhqX4M7XHb0
4Bhk9cSmnp1GBjkA8cF27jSBsshCrphI3QTsZxC+wKkyvc+OHYhI3iFqrARNweVo
m1aKxN7vvXv7zosJuvTSUuFBWjjYzhyckz2y54JA74cJSKplgw48LMKf/cZVtzXO
AB19ErFHXqJ4h01SHqC65ziY7NNyDSkKbpTMFj7IEpGfDAuvB5odMprWoHRvhQZP
RSh8lKKxpTMseaZG3R6seITqrQUvKu23u+JqHVwESFxEaKJJHAMZTkuvKjActSlJ
D8Qi9EwVIWQl5GC2iXVVGzR1gfRoqDcDr9gRK540Kkf8F6fmUvanmE75U3VRj8Uf
VJhc0o63SUOCObTFiFOZZEh6Buxldh/taeRHQQDWnKW6Y2iL0ieb6kni9i9tynAt
+TPoc1D57GxP7hry4oZZQfVvCx6ZbD8GBVogqzjL6QhyEOECgegXcH2Rwfu4NKuk
PxE+LF/TuCIc2er8sTUvD1kva4bauLT8D2p8obcE7ft/e3oQFW1SH/ErHAdmQwU5
FmP/QeVOKYy54CUe2+ELUNFdFCkwfwZKYfr6PstRH6tpNFyEhMIMCp1WMOVag2MN
3N0yXa4Egk01AVjKt1bsIQmkSRpJdIW8nWr7O+mJ9pyLa7FRRz43rrlx/GckKM/n
8vsI0Uk/2GkR8IbYe3cMSiAvzpmwH11OEfSdh3qFu3wl/XTvysxr1rbMliQCBG7A
UzPMIu0f5+LhF4kEvYZpbdRQLHMVHEv0pQAfmq0No12/mC00FAsFne0r1MAAj/PJ
3KpAGIUhMExN3xFUcc10S+BWRiAY6R3pLd0DfAA/KWiviD1pXZXnFNZoHqixIDwv
3I36w2pJnGnjds9YCMIEciNL4Y/q43IxollwbHgJgj6hr+lwsC5lB7i1wEdrmhWh
AlHoJR34pmvvara3OHXLM9jxIRenrGjW0tPre3lQVWcdfQhvx1dlKGvqJDf25bac
V1znMsTcv1h0EcQkA86RMwM7V/QuEvG3imDnNg67UmGByupO11LYJY/9ZpPFYL/l
bLgzShRQDMXyKPJ4EDSEd4lSg91Clh7Ip7+jPhR2UfNT8MrP2t23yhJHiWjDbw7L
m8MVrPyJOu2xcbAuXyIwVjhnRBLtLFsjdY1h3q3JNlmyxVFBj0JCy06FUNpFLMeb
UPbOSn/a/qwcdBl76DpXsNrXq8x/2MnbuXKAJ6ReIf7pjakw8QndnD7kZAgVuurJ
PotUh35DzzJH36pAt2tH4eEdJ4KNEqTEjxmU+408PsdGiN9ee1u7VdZt7hL1xu9x
k/1nfMEFcNL4IlncI+XaETEt15UOq01AYGtzX45j1wJNzYrlUHI19T/SUdw+wzyK
/AcGsCXsSGM3CcXS3gnDDi7X5aPZc5phdaaGZFfEecNaprqQEaZMwfAi5ksUbaRa
uRaPkrVhHFtmkcYxsJ21hRLjdBEy+C0ZR1gIllizNrJOs46u86VvGPAovQQoRRco
T3Fc0oSt5DD9F1eeLbfjMC+jw3dYYpxjB0PUyP+341LrMFsSrKjcrTwwOBf/ccoO
pDHnP/Br2tgqa2jeD/zeC01seaHxo93v1OcGDhClGEgNN+5fKHIMjEd5165xdx74
6VtsIvxAkpvgg+K4gwTFUXxawd4lQIMj1fMbo8CieteBgsg1zOkhknRAoqSYJQjM
tWhP8LOZtViEz2saNuuPedggkIK4auEowrbi7Fh4uWN2gwMKjC2BKIu5GI57dCDh
8tvRxtvOvFCkNykQReq9AkUVDkW52x2x0i1l5qH23gP5uNniCPzwHG34a6EY8RzI
0tEfwanwlAFNpe4i6L+md8hEt3SYFNPsm6UoRzRyRoAaAKjZTkXBidAHVh0956TK
Z4naZM1JCQ7CUidzn22VgwP2ckt6tZHFM4F1q8+oZP99gtsyWFKB/6dLSU+nXPd0
9Z6/Om6vxM/loMap2fXA253mF8huuWsOhg2PbvuRGKltsIDKIRy43RISpxluMXJA
yfs2GYzoE2mR/UKKTmwV5SvMHcE03tFjTpiwV5w3U+V89k3FZqVhO96/vZerfK+v
ytz9sSwF87/atK74XWPrkpdPysVtM7fWzMybIhoGoeqMpP36T0Ha/i00B3KPl67s
JMWUo6UtSXdRKorfRW+iMSy9RWtE1EGxngL1rLpIInj2Eid1lDZqDyzABC2PPrZ5
k3pRA8TLwQezVcK1cFwiqIorsgJa2L9ifXnw/lImMtSKBtwg57Vd1hulfiZxswGO
q5nku8qIQOn6YcOZ5Lqof4C8GcUuttMkosHAn+X+JaSDMeyRh4Ie82a+lIiXMHOo
MXSlzKuM33h9cAfIjqK7WRlgF1DnqRUcRKvFrACkpvV3fNbho2LjB/WLpmFFe9nG
YV2eJrSGVJeApzWUOF9R7b1dLnu5vDYfZGhp68Xj3596iwFAgSCibeKvYyNxDo/j
Ik3WiBnto4AJPxZ5fN3T6xKESQa0XtwEb278FMny6mef756+kai4xI8lZhBRDHSl
5WOdSR3EXwPp8va7e4oDyCw3M9doQBgGQ1P/LIYEFHPK0EQ3kOYwOzOUPjXF+crA
e2nF65nUop1kvhBI0FGJlv6qqO/gdeNzXR18m58Edu9zqHR76MeotI0lbUn20BXU
KyM9rIaqjvQ6Uygp/CnuRIqFH0e8JFgy9aQ9UnsaVnaUWY00VXx3AOMCD0C7uIs5
55YnAFpwWgr3p+ae5Dji4VBFdNdgZ+V401cm84nCIXmukfqFU6JzcBNm53IPZ8zV
bXdQ9sa0dcrBzSvV7TeJqbJNDC3rrPrTJ+IEZIhlNMLsQftFR05g2a+Ss51Es19m
vh8A+5SrlwvQy1/YNiXwRmUk28HveuuE6SyEmtqbgpijSD/uvX2vRpTxY0chliMK
spEbusLDlTLJvxZXohoCOExAdGhhPmJlFIxj+uqPDYw7s5KBWXnO+yqqRLsMTc3g
ejf+i3BcS3VYfGPEpzIsSzXbzPAiKbrwdqOTG3KDZeVp104iIpZhlvqgxsHebMaK
SH8Gc1HpAXoAUh+4VSqRybZ2uwUUFDDUB8ZKuUA7SieGqS/YipDshOGep6Qe0RHa
baqOtlt5AqeNb0YjRE08LpejTut2xF/DYLQONY5LpfCtmaN9B/hSuTJ7sftRoMQx
Z5VmVXpCAD59CzwhXjnuEBDLv0TBy9KF9rkCi5xEUYBWE4LJg5OgL2X3wLckM4/4
ld2NMHXCfQemyGSPSh3Zwaqm5/Xb15SlHEQV8xd9gHtHbRzIWL1t22QmSiqMTcHG
2/o5brLzIILmkNa5+X1Y0j7VnxRs8HJttBVmSLiIQVAN9B3/l58cOLlHYRpA0o38
UPomXO6DS3HCKvczVuRddgXxCK9ski+tW9VdnFShEGuRSlzu5pniRzYQVWLUZMGO
TnqssMUAl6/IJ21t8RN1ggnsbbHkXFNor/8NQuK3PoF78sE9iFq2d8I7u3km19x+
nB1Ch/EPUMy0qPXtafSYvYLXnla+gevi+rTLos1s/wz8WzCQFybT24APuC5QChOc
/TRFHecmHynj5dKQN5KRKWtbUX8i410UZSq86X1K5+/kLyoxxXLC4vTxImkbdR5G
L4/AOmNCSaC7r5URwWmYldbWBTIT0+i9Anccz0cXrdAmfCNAt21MYSZMuY9U8V91
uGcBnZAf2wpgDMMB5pCMj+2OmDOQ3fHAymwu2vDsh+O8PrAQbz0/vomRXSHQD4Zv
tZ1dPdqKhDIVtV1+zZCoNr3tQpQnnLdCDvlnA+4YjsWwMThdtCGoACTzNrM9MNhF
r1lYjXagNWOFy3zvQQB2wIIoi9FPga+EkCS5U6yRD5YasuyktYCk8kzs/l2UWGwn
OEUhWr7x/DcqXQ/1mONt0e52LUvgQmuKNH51B1DpzoNs1GKebd5geUlRAhCGlqSY
VIWt/Y6/75sigks+Pmu5E5Jdf6aN+pH24WVKhibW6EmX61coXikkRStgsNiz8AUz
F2fIKJI2UbmdnVyGx4Not94eopI7xmfm+iMKzZYdcMM+A1TKgnpzD77pHyPQnib5
l7KhZjuOKjOYMkOEj2JzR58SOgzqeVkgG57aVZUfU30DtWZTihKqf60xuoBbDhrv
WdXtykTJq9sQH9n+XrzLfOlukbd8XW89XrkIpVEW1bgYxcfFl7f9Z/4C378qw7O/
IveGCDeQ4RoJWt5+y23dSgHE4ht2PkusumJqS9CmX6QkGyGwPHbaX0SsM4tSHpHg
2qxJCa4lljU/3qWnvUKJLH3omizfSWRPXCvoHIchSd9BkwDFkVHmtPLA+0oy4bHe
vHgAMtGds5Z9QG68sezBrjhojTBJEwqmDFZWx8HVq9Oa4lfHaW38PCxKbfRMG4KN
gDiJG1dvxo0agEZxeR9ma1ykmarxNM72jjqCZ7ZgS3WlZe4M9CunXHbTNVmLJhbr
WWDqO2gye7PEswwehZZrbiAfpzAhI+evwPfrx9BH0tuoJfocaHN+KiGpXF+PqsIK
Q5MWnpTI+Nm/qc9AurPJQjEaHdiJr5OmQWBL++qulakySbLLpZKlqFRzYJ/+ybfS
d71rWIAHHf29XTDHikdC+qG9Whpv9C1ROksTzhyXcn2otw+R3eKHt6AJutlI0LWd
Ze9xKMQzGrozzSTxakRqjjoIkmEySQdBBBJdQdiZazXKzI0biH13nw7QiHVi2ys9
k9xJl2fK5tnWto5uBg1aNw/IKcRl3iNv2/2cCg0oCMcY6BYc9ko4AaRVVnH96iH0
1WvLwQZnnq4s4ZVvbZUd9BcImZXOFI7UlskngA81A7HTGM5yIa6EC9ayOU9rFv0O
TRBAMz04yy88C2Is75/iwy3rGIkV4BKZ+MR2QUq4WYATJH6rjW6odPViY1x/gWrx
Tb8CtWll6wxYd+xGSNdKCs3rS9tHf3pcP1OrSUjYu9mJ+r5bQRssfsG+92pqXvZr
d3RGIr+GmHNAgqdbCdPfCar6v9sMjqRBxTcU86ncHjzASd2XveHrPRc0pMw8/xmL
axXl4NgMy7la+DDPQckSaxLKfhQoFW5QCwwsDcZlS2jBtGuOCBM5WIO7l+o8pDIr
Jfc6l6ddjnFP75R1n7v9cIhNBNy0fmABZMTnUB84dnVzNUXY1qj2OVd0LQplCwG/
L30iKz1d4dkcUgz8tbtSi05djHjIEXwn6eEl6rG5V5C+rdCew1ZEZKlbTIql4F6V
X7/3qsPVaES6IxkX7Rk7BUG1STAz6QK4Xux9gHJ/OgyTEkiaHuPAwibUGBJUVtz9
zMTv/x2Lv13Oqq6aFpMG/DoewYrPqEK9m7D4nlLxvh9Bj4bkMDaLO9a7Fpm/8XCe
AKTudG0VZX621HpLotOWcoCEw8kFHExA3hZ/5oq7XUajGsy/i3ADLzTYrAXS/3BA
dVDdSaSdItIiwO4Caf5+hM73HB0xp66cEDDl33jZgbdndHT2Ek3Unz4nnD2/o8Sn
wQHLEyEbH0N8JMvc0YksL8yud7pZw7MdYmrLQRgc1/jZj/+1zu+uwGdnV0dPCllm
1rVWciqSnVio073+OCqopYR5CyGSMs7SkoJyoJsNX+Atm2NB0JMIYEotKhik1GnB
KrBAZth27v79VgWlRfpQGeNYnGqvTYB+wYHT/NLvnYvxRRf1RLjTZvG/f3cBhAqy
OhP7zuBq9oVciXeCS7hbIft2nHRDr1Xa5SybAIOnaEvwyxIyjDDiZ04IxMfhCKec
PfexwQ3HMcw4oCFXhYm/34wZK2rItpd33RKPCUr0ppGYSQQc6GVrRBxTYEfBumjg
G+APb28eO1t6b0UX+m10EN7A9LoTmJ5UYXTAq6uNcjm7bBse25HP4v+ULFehR7Ak
oMk5MLbGNGphi8re8wtkNlBeQVFkUAhTolBEk5dj1PotddkmRQb3KZn+Q/itvrHR
rAT4orn3g8WXJ+0/HRwIjAdyswAEYDJbclI/zkmWzMZaK1/NW1PcbCBuI1kRXTDF
ID05Zlro3LNpiBgn1jpWtUgcQ36/8eA+60ZOJW2xMD4sciBnIGnymZUfhfZyiZZB
zx+y98UfCnSKjT7vLc5mVduDJUeA4Pj2vkeNqNToauhcPy4SU3vLhsqwo8+7uNVx
7OKgw1mZsInO8QVQBCbWpJdZPdX9uJuB4IBXlbEfQIlSWoOqoqsIiOmYFoGpGOvW
ajtYu+0Vd4y/TICoWqs/b9jYA8SDWg9QaW/WmWVdNK0P+iSYAsSWNOK+JXvMdOrb
aM0CckfUVQl4DJNph7EZgbxnrTAB/EDhh+AxMPtz9LpdArQAbTvCk7fvAQOqszAr
3VD+PTLczO3erTDbrdYIDQQhIA89Tu9JLd9TyvyXZW/sa1jeLC2OKnC7kcV4QWjn
N2309GNY+zU6WhhxuO6DiK0s0WNZ+mk/fdXxGNWebEnIFFW0kJ2XPvrCBEw8sNqC
lk1Mmu+UHsvWs5BNhvWTAnadadIz0H0lqw40ycputWrARcTc4S+55eKm8HICRd9n
UYx8otSDF9biWIf4QCGXN4bGckBqboG5U/EwXUJ7nFkdB1UgX/1FlFQyLGIElg4p
8Jyyx9+Ro2RXjoGRJRzOWIWGbRLu/rWIPxI3dsrVJlOoqbOuuZGYIfN0qmtTZzY8
yFgaibIAouNyJc/T39FGIVuYY5WryeKN6CNz+DrBMup+ovhCwI0oGSSOWhYTJomS
7iX22MA0X/wtLMoXoj3KPNJ//D7nWBweNrJvI1iA0mAWECxw995ZAqoyhPYRPtxP
HBR3oOSpN1+tykEM2xk9qdoqMXS3jDhHZ1H15Iv/0U0sX3QKmYRe/Zeuc38dd2m5
zOZIWHUDXHAxnlomCvQVmUFLvEnSaZ567NkphTJhgb8jp1m6TmxgDBQ+Pr20J1Dt
oYEZ+3QJK9iuPsV3GfRspKmlHyVVCQIFLkisy8WEU5gs1Lenadr0K8ntFM3QEC5g
pJq2K/gjGWzkKrIsnzGqMujLBTj7noCkY5aToAy3262liNZx7BhpGUYFwOkXpO5E
`protect end_protected