`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4064 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/aJDh3f4QA2IJbr41pURffse09DeXuMIN3Pwj+x2n282
fdjyCuuuL/QhgyKwZ1vXpShPLxOKJZZClk5LmYnG2epfLifTUQlynHuidUzP/xiH
pJPDUdlrcvA2EkiEgmF1WZxBEXRKvGaA/XRX35v0ocS/e4mFoLJUnwXNHRW8hrI5
pVQt2vBUoPADX0iPEKwbjthoSHVPz3/H1p4oCD+jtXTQUqIHEDfQgGhMcNuMgaIe
eYQNCkis7Nn+b29W+jGKQJtv9qr674n3oYt6TdwnNV51kRnaq/rE7TxHCjAeZD13
9tUPee/nFSOQ6G2Wq1QrklIVwR3wz7+eodQyb3zv8uWai3Ws7Vh43cS6b/dfSPyZ
NtloQoxz6mQaAcgUKHcUvQFdKoC932+lmFCVwZERZakmmOHo71cOJJ3K6hnTkAv2
IlPraHfS99p+1A0n2KdfxuieQvvCW7BPvKkuOh3iLwhmwgIQPA0eAMljYOlytYCg
xIlUlACFAAt7EYpodZ597T291V/aKh0FTd6k6k1HFAIPSg/8LHXiDf2Pu5MHC5mc
uUIbWSTDPonGXscKXDsoP70XGQgAvWFzhoqCLaEccmtDjR0Xu8JSx09vrJcgDxlc
5ICQ6tQ2SpAi+eWRSILrvCWxYUz8tc7+Jd04F8L1h/9JRtxEKmIr5rMjE2fBcmzE
bHi3M0HHfXfN8s+8uWn9dInxawGWxEOv4n/YxvGVfMH5xHsVCo37WmAAdlGfSjax
JikHlRCisWTNnatrbXNCVmOVEQBV7BeGpEHVRrb4GKn4qATwJhhGuQEo0+0p9OXP
+1E3VR8W/rlCC1G8tZpJYOy1O9hABt7LCLiuzbh9eA/7CMdkz3zXfHoLrLi2EQR3
fnymAGXuZywjxnGXo6xU2wX4jVYt6tSu4Il86pKFK+teB9Jda3dHQrHT4oYSzU8H
jbHt5CPMT+GD+A/f8TRBP0mQIsRVeo2d55sJtryF/6cgoM1zAdeBvb+n0IcGA7Wg
l8fr9mt8bf79BLO2iHVuKs6k2aHp6IlFO9Qo0sPoDACI9GwMjOZm4y/9fQSkJZw5
PHYBcooyf+SnC/153SUldyQNabt+t/07Xk0VvKh75W2nylS+IBdCAxyWMakuM02K
kN/SADS68+M96igrf+1ePOBhl9B/PH4yeU3TUv6x2OZL/SW0JS4EaFI+Q/tVgA9Q
8W30+hSjhzS3T7blu+zhNdHib7AKINOqfN2oZMkqxLIAgYinYQyGWlJByLqtUvpk
ZZG+9acZjwaUQ821XnL2/TIx7FwUqaoB+0aswA1HDD6rnOstEEVKeGLFzme3ekwD
DO+c13hlfpFzbtYrhFgHZuHUWqqvZabEwCp7AiLw1DC1A6u7R6ZFqOL28odMY3bO
Xc9Gg6SL+9gt0efUe8h5809Ix1O0aue604EUnMm40o4Vq9u9Fs7dlMv0cQs/Qzat
ww5ZjT10SxuTRZ+e7RgkvhkACKjFi+g1eLqWVsok5hCXat8RKm+XtOELT8TI2H6/
sDOo+rlCKCEGQUmgQpC4W3dZM7ZEe0Q4xdekiFGgOwHBlJwNmtpl9hZ+NEb8i4BW
KaI1NRp77GMiVT58X15+jvkgkOGCNon1Gf+m0vXOjl3GWRRaILf34WOJfW4bSvG8
ktEzq9N7qnj04y4Cue9mkNKXv1ahysXA3osQPbuDlKkTBbWQN2uKZXK8Je6h1ALZ
ucW4Ok5ufnQvaKUzKj+AeqK94T81klji2q7/Bf79qF4cqHrsyxUa5BRZ1CKmOiu6
ngPEAOMLkG4OBBcGIC55VOxSpHky1wo91mUuA+3njeMEcAbOn6nVTx5PD+LxikWr
rvSYivFhn2NpVOjd1/HgMfK0U/Ew7JX23RheVxp7Ha+rqOFE7w8tR4adt/M5tjgh
vHM69W44W6LHcWGa60qM00xDqWOaxnI5cS4cwLaojlq8QRAvqYESIecJ8puvtaPS
OAk49wfoV74yxiEG2VPfkxlKDgXiwoMj7KhVsYjipxAMJ6HUyRVFAvLcyv0vTWFq
kbJJe563AbnDqO+M5926olQVST13CKqNAd0AfMQbK8nn30S4cE4jcfEe0kJ5f0mh
kSKZWiXcvx1pjZufNfAeb5BlPCMPv9KVofFuKE+u9Aql1ZUfVU4RpzzptSenLCYD
Jatzl7K8mGqOGrU+l4rLcWGHHrtR0ibM5fT4aACec9bEfU+uXhAAd8+NLsz7UOGz
oax6clYC/zh5vaBotBvJj9dGiUvaYBFQvgBfO0WCrKM2bYIr3WQ4omiluxBksJLF
ifV0E+uIHjqDRLsfEJPXVFHduVgxns7u+fqhlhDqJjxoXPFHIm49l0obMmJjyOj4
HzX/eXuurTCZY9Gjq8daGk86RJNSJlF2EhQvO+6vHFHbM9qQXK90SGoRQ635tC22
kYRYVdfxfCvVf1rfkO9GKj7Wb2f4JSju1ncrL84s71XM5mNygy5Y9rzM41lqM5MQ
VV4DvZjWS6y1kVdnuF4pURlKNSurJxwKlpzp1cRqE5ah0hNlhL9aSOoHIVAKm9I/
BPpusP1Y3NJWTf+XcpWeiOE7Y3FI1sllYCp+J+3ATEEj42RNT+fMWI7CRuqKC6i+
Utk8Jf82/2kv5FB9+3NWjjfwsZGr/lrq6VJLCmzLz6ZSQdoiQf8CGe0sEYAaW1MQ
RGBSM4COaSlVndxfz+CyxJ/Qs3luZ8LKWIrfNlNXV/bR97CeAdunlLfskGlOI5YC
MYp5x6msxePr5Oy4fUyYkNOz40LG90SsepL9swjpX8VDDSo6LX4tctafoW0rvTrt
LHVOQ5FP8oleWQQ5T6jYdiZ/QfGqqJxgxVzESF0MiWfYYxEMNmqjhUNtwkk3lQ3F
Qc2ZbbS4VKaOXULxXZ3HoEc3zy71uyxluxsdpYcgbw601rxv/RqC036nVc+RF0P8
5BU9UV0C4DbpX36G/qzjRYS3NpL8UIO7b3LuDQdn9ncoWtr+LWdU4VzaLxTHQ4My
sTrKzgTSJ7qqYQaBhaTbpKgQESuu4lNGN8Dg1CXpEoWoNrFh1egC22gOBeeSTvEL
bLXv4EI5e7lBjPjNeFyyE8Q9bayF3MCi1w8ofvg/MzeBn94AL5V64Ggs4Gt5nkUQ
6PQNtYajFKtZOtsZ1OETZxqaWmWKno2ARRwuF2nVnItmUcQpkRg1/+7SYyQPMHc9
rOcyauUIef95r2Q/IY1WH1t1zdzXLTNQK4RwZUziOcuoal56LBMWw5zeSEPO1AiB
ovC4Vuf3JVrFpkR/+gl549zsnk26/QfQBX3nHGBY/Pkt0Uxg9cRe1IaTEyfdnkRg
xUdGPylOisma6rSU3qwf0+USrMAmbFg3DxyHHgn6KwjFT+p0GogkVoL7w+jmplyR
tai1Bo4/V20dCc1MnM8NnfLyvxRmIPgIAyg8u2NHv0f2VOAzNfbOSl4E8h1w/HfG
TUd6Ijj64H2V26cULdx6ghI0gDqyH9ZlO0WAhcGUcgmDgpVaa1N5eO03utYfHLVe
PptbZ4BxhUghZiD9wYbM7vFs+h/QTkHbtvbNBhvZxLuCXPjhF9YSEdvNFOb84cqj
ZdiSoGJ3zd4v3gZsu9KEzO5tfb+jPOYphXI7j04FE9LiTEHvf4NQ+qHk007TxtyR
nSn9Yg2mwFcok5IIYPP3ima2Zgd+O3iKgie9cgiOB6qyZV4YVHa6QVPFkKP84EuJ
/x1beGxxga8wzvbgio02Zk9dEXKF14vPgZyA5alXpITjMS5Zj/tE60asB2/aQJ8z
NzvHzh63PmeWEJVjpTv1Ytp/y9AIe5rFok2PDCQ+A7nfCfqRqjHpcnDxmr70Mdgd
QEl1NPtbKCmVVuy5/DHm1EeMuI3WHZH3o3WoyGCGoSQ6HV1kWcR8IfeJIXLjZqut
dXvJI5xuB0UO1sJeKWuGADRhSMElRTetnVxO9szmtd2h9MkGtgLrocNKDHlDJ7pg
HoCOkJuC8dptol4pGcLiZpbPUe4I8HHLBhR8Pa8MMvJDMRCSG1SfiV6RDhma5Ku6
gWt5N2McJxBKrbE+A636jCvVCPY1Y5r3QzRhrVx2hDrOf6aFNY7wR4rwzJUYKVab
ZELzP67skOFhqSi54zeVvU5tK1kmiNaIirXwwQuL/uBxeJSUWvVSV863XQ6aILLa
0JaKYazDpbyWX4qwrtfICLG6dgEz65nSJvL2iitV4ECCoeq95SAZylMF/fCb56du
vIklqZ/Gq6SH3HdCRsfGKjegH20iR2JM8K3h3xSEZMxHl09dNPBJXBNNGoo9Mmv8
8t9SRPgnShblKMcZ8iqq437jhwOAp2EX+ByPL/xBJZCVd8IAADUcpnTFrhIKhK0E
ExJawX+knXthduMSoNV1ZXrr7taOi92Ya9elPbV7rOKnishxobirOq3fRXz6uqXY
SENE6VdFGTWxDQNwJDPEp24Gd5VdxiTNihDj2bphcjlxqzVcsioFA/rSjwJkt0VX
LzAB+ZqAGn1Y91xroCeQLnvvHFn4bR1chqXqXK6HqUESy2gzbVCuvjH5emQMwsta
5Gu1rJW3ZswqzvGs1RstFH36xe0QRusJBzbGiQ/LT/NMlSn6rfPvrmi2AGE+3/jv
QCK6FtFAQJH2GbDPbrsDcBOLXtE14/wy78Az6k5l4EALxcYl8rPBwOY8Zoykcp4n
tXKv1XuK6vZvaf0d+K08E1fdbU2nM6uiGP1Q1+OzwOpnoIo3weY5XQAWZKzPpNAO
YQBTbImRn3RPGVVGRY0TlmZr6kpycbCrwq3gfljTwosPo8DMrE6pwu3s1eZrn1WF
Thg1bvS/q0GKCMsCXAFImq4JLq+3nv+xyYTeskZgNQZmDOXVDe934770SROXwViZ
zF5wMFUtkKRRwjGlYowDJgSk8oNi15Ld43jZOjARPdt6fKrlYyAkU0QP2QSYLGKM
/L0h6fAOH3/39IOe3DB1poXFBEnClbO5wlzaJxWXpzRu195r9CxDI+vgxE85KriQ
FCdvOmMorM+VSzxty07bG88Eg90YVn7kARUFuE0w8yHkOvTKJ8SROb8nJYxAurz/
8PLM5lxlKfmRIfOUAVwWn/ka8P15U4XvjsdFvckcM+RYktAOhMZrcOffrjkim23y
+1kclvtzP1k6w5ZiJXv+8IyU6QmOn39Y0AXaNQb02WiPBGPVkdHbspNVuSO/QURD
6/8qu4dvWY31C3opHm16+vRGyVsP0Pr6JCRLuI+4RxaOaVn93Dj0wWtO9rtXMxqY
ksVgPkjvL+8WrPHIoPNjLbv3ZfYHCDmCS8n3ZE22+hw=
`protect end_protected