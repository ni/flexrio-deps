`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20320 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
L2bRNdr1lLBT0eERw3vGlKx/bxs7J7VtkJsS5dvu1IABJ6w/3td5OcfyyIltmWIL
KG75ycV86p94HIFNCcdupmmGLP5U554nI8QuU/AeW/TFnom7QjyPTcbTvSMOsZ+i
K4P23X7esP6qUJEFITIWWDHLIWocwmMbhGWVlk8X82kkTJL9ehiVNglbt/PkGEUZ
jxNaRon5mLtnWo67xJpOoO0lg5ejqfpp455X+g/M2OvhMKRcHCnDpUbIgBieB+IH
srlXRJ9P2Z5o3qVrXlMYCWAnYTjO5ymHmlRkrYtre2Y0uB7r2J0M/3yYfwMM5GFD
mtdxVV8Od937+In7eQ2EoDObcH0aJrvmn83ooBElAmcukdPbKkcA7rbz5xjyyTL0
04kL5PQamf6U2EoVswF15z7Mpq1XfSI600asQxzsDaI/acpIBgQ5KAa8VAcWwLmB
BNIhi+8bo+zYkuljyfpBIK6TLmyN7ZNnaUpabX3gqwmIM/Hlee3Feb4HMqmG2cJM
wlikBn/m95hCpo+XZoVUxX2F7NSpFW3hw8wq/mafC4zi0Uue4UnxtbmJCmCDOuoB
HeCW8IjKq7nbK0+zVRlxybFhXHgy4jGeCKlUKT7BzKxJDp56iRQcVbqeLSlD9s17
+mxEWwuJxm00AEYF4Uuk6Kxn1g4YBmWyoOBr4m0iDeSi+CFR7Ryfi+QROiJZpJst
l9qabzWnsGzDzRnuhwBhzL0ooHj8fpPqnPfqVN/rvufRMzxaxq4UO7DqJoebE+Wi
G8vOJE6pXADRPCQ3N9ER1RJUidgPIKlTvxP94KJJxBoJUDwClyjTkH5UAGLi4w5y
l1IQ2v1hoejM/18dGI+oXbfdxv12y0Jzw7VtgLXs9Pz8jDvx0A9atRhlyu8xBQlK
oitRbEmL7VTGXbPw4GDccl3SD5IcNnZl8nGLuDvHPg9BFOr5ymxxLJBVvwNC5wWU
vmtBVnt44PGod4suhH742UytmagTihlWi54xxbXQP/kCS2ndt694Qr5hBnLGSeJM
GW1ckCWcJd3T8Oo25iiHun0eGxRdpuwmGjdh8tp6hc8LQ7+S+TF1mVtHin07kDSO
w2lfHA8vMGQwf5YkOpGjz9DQB76DD6JYW7GswmysAxvxMVZveidbUlZLBfe/M+sJ
e8U3Kcd4b2Fi6jc5lXG2TDuBKp4DWE+4TajplAj2qaHuNT3CBUf3cN9CaWcnyrwL
DgDrrCjBgd+4rIwNh1iyu058N+uyVrhtkwAOdhDOqAMFiO9idWJorphPmjVhzWOa
Ec3nRffnAEkHmK2yhV+hW2HFEIpU8mJ2tPyB6HZ+B70Su6G2ikB+Z4QmRd0Iacwq
R+doUMEL0igADJxirYkuzcmoK7JgUBhMVz0/p8DeC8qG74aRZCCUr37UU9RLZunK
gO9Bj7+XQKC7pmzUvcIvGA1+ahNteCX8hEXBnIzXuZ7g1sGXwZixoS+s2SnvPYSz
cJ4Cs0bkMTIHLcYju+9caWGB55geG44nQVNtahPmZ8nUAFDRoi1JZxFl6XIqN5Bj
ygns2/E8LBr2YMFpmD/HVmFeSF2oP9ghaMe2gVRVkK8YYiXcC1tjnCGGV8qssO6G
PnsTZXbZMVrYU9EoIKzT66NyjfShigxOhdBgGkRQaDbrOOkb+MabEza9Iqhertg3
P0YAR6AC7ImTbHU523d1AP6qNajaANCDXS477/wiBgSI4wdnAeU8m7FW596fB98Q
Y6mhX3WatazDHaQGhj81HC1+r9yH1yTfOGbSSgDw7YyoNfU72OJndUigCLa5raLh
wdGh9O6RDjUuXi7I5ktvPLOBnw6fi0ppObE9PXQMrGOZYxRinUFDyO2iBDHZecXM
QCQK/PUWVWGa2gPceXEGUljeRFdc/pBMcswg1TZrdd4lGjv/1z8ukVySVVTTEv7k
ADDGUjCMjde6sh8zpvv6i6oqKm0pga2i/5dsqwd+sYJ05zouKYYiRRRb2db19kv8
CnTZk+cuptmwv1aRRUqZcG1H0NfIXxJ0RSZcotfAoRykoQCyopU0SuPYyTwlGalj
omwt8u5AloM9e8g0XfYT/oGvQZTsH/D+W9utgy2988inVuLBhLiYVJsqXcTFSkQ6
6NSz+uUa8Qsfi2EMpV71f/BIGwovi4DqGrv56LWcgRTCNdZTWTtimxxRjaVkAkXp
6nV00Zs+FYyAUuxAOAxfGavMwKsOeWLFMFYuDWzJAU2MEY9abREYPpGWoPgEzcdz
tDZkw10YiVKAS9d7Cxnab6roLWHSi63zyUXef9GnQM90uzoV3k9ExXC9k723sY5I
chE40p71pRiSA8ASxxycEDuhXIH7iTPQ/vw+1sEkXRNP1te6NdXtzUhd5kAznSyB
77+oeNnAUhGcjxnesgBAWTFGQDO4YNqGl+v1Fc4LVALgH0HfTwSrBScCvO2CL7nB
0/Y28MSAnhnSU7EhnNpk9LvwYeriFacnlEyzsdpHS0NubuOvHWKmBfqUhwGuREgX
Z0TtbTB5WCkLM/63SpTKogT7o9V4J8Zh5tjyIoBVg3A2yu/vSlsOZC6pLyivyjna
fCLPQPWc0AVGYqvNauVb/bl45zzcCVRrFygvS6zolUeg+B0pTUKP1IwfEZnw6CJG
Ed4DhQydtg5BLJ+xYMNk7m+P1xWM4zj0ORDp8kdLKaV6HVw7up5nJF5ftRYmsndp
c5GFA+Jdire6zq0HU1Os5MI333MhY0mQjCOLUFLrzoK9cK9qXUj3RrwpiWnJDZoZ
IuIJACtInESUfim99dPjGz5I/LehZYA1RZ4epUHuZx2+i9BuAMzvpAKSxUdr/ARb
v0jYRncQsSs2QB+vDHrvB9RC/apJtNCct7RLL/vcIgApS2Q6EQkOp2RmoNm5uaw1
UfX1kP3wLSuM9+Uka2jmGe9heTRU8rol5cQISreHBbh3wmXCBBCex4r3B6ukM0Wt
bhwFh1D8vlCQpgD6fSED+4tMvSPSEWJ/J0q7/hdSCoZw4qLdGLmexr8Rk8qYhy1g
Y1YuVaNQMuwcG20RVCb4ucZbTPTVttm+Qk5kGwWolZoQxXK5003K1xQZzyvYV2zZ
48oc8w8CWEOlYVlIvVjfqFq9ajQtK0fyATKx7jcS78Vc6dyweDWEJvZk437RCp+N
QietaVejPaf+3AV1b3M9lUcHdkT04LIDxgFKP9gRWCHg+9yng2N1GJH0QYyxX2mH
M6vqseUglM3SlkLHEo6pgLNUi2PfKXQUJ6zLpHttN65tdb6Eaif2PA/pqwgFbIAh
s5RqeL5D/0JyfI8FLWGX0F5vWHP04Gy+vuHAG2Pj61RmYQKjFLScxSF4TYtItE9m
+PC7iogpd9Is55hCkgVXU1al8yj4A6oJmXUNu0KBl4UFAtIn11gWdleMOwQlZ/Qa
Xisdu5xG6T3hNnF7cRzD3GDWT4IUyHPIdHKY6SJhJnp9QXAGWb/9154hsJ4FPDuU
o61Cln8Qi8M3LxNX0AaPf2kL01QTABlcsZpcNz/p89iOL/Kl5RihKvZsndmuCl61
KpCsrFZCOAPbwLpO1y6a79G6mhOh2sAEYMFju/fYcGTRq94an/PBoPW+/bu0dZcP
5v4T/LmNaKs1hjxehFCQMQE0D3ckELFFISvFH0wONEACfnhdGUd3xy8fno14lFDN
xTB2crRI4zOFiHFC4ukz+lOImI/YwikdiaJJWD5QjPnIDPxXDWRG4fFFGrT3R2CW
VXGe90l1aAZ5rslTlRIqjKMBTmEGY5xs3iZJDicsy6gfAlh0pddPDqAapNMnzVBo
nmqfhisv/6ddCC1oWHnmZgUG4LDuz8h+Rb+HINhJVAYePPBUkZMsXy3Bjz28eEsr
pF2oqj3zeXQzUvJ5g1x7o+lhWPC4xHihjJ3/gGQBkltwy0JMSPVykrfAfU+lywoS
nmvesNSTs9oPyCH9vIhZKuBLCCq0uzfm8DstSGODPOJRHHwbgeg86zFC8xIXfsQM
JYi9MFF0IywQLP0dSw8aIqGhd4VYzYpUEDEBJjmc/o1sp7GTfQijKl1e85BHpdsk
lzQ+j0fWpEjITa/spV+clr/x1nHZVABeF0EJyQ0w0tHDkUhoRMni32OutwstHIL0
SyLozrIUpM/EHpBELEhB4nWxBuPN6+n1rPkpAfJ3vz56vN90pOI52Jpo39C8Chfq
R8g87Gt/ernM6Hi0tMMVMY8+gHXU0L8X+l8H7xF703xwTpjumtXo0f3bsgQwK7et
RnChi3pndC0J5cclA6RcsikeIOI8sNcai/DlGpDdOK1BbNByJjHVaBws8s0pHO4n
qaSjlSKCzphRA7+I/D77CXwJ9N9g6FbURsxQWJCk3XGylzvOXEedYuMFCJrhkoPp
jabZdWktxcmK2N1Lajk4KSwXrqmGrv5O6sJlixdtsx7Q6w3K+mhV1nemcl3XGO/8
0+5TbxSTNd3XOUn0tUN91H9yuG7xYVKd6ZPAVV/mFz0JB5KGigeAojr4PlqMgBUp
4fgpqkzYSWjBzlWHy0Xf95Yw44sRVHR4p9MlVJJubsoT16y4gsiIikORzlZfbsmP
YkbLnQcntrmieGGc9N6q/udn0z9UiyWASF727zG7VaW85YjyX+bKkiApuAYwilEn
Yr+4fjxXqbyO0hR+gSaR08ypVC/R9neebZoegA0FgQIMKfuG9j94fHslNTabwsB8
A+9Dyh6tsMmSWuhLFcy8V+mrk1bg1YySO58LjhF1EU6Z5MlgvKoEoE5HOWEca8Dh
d7FF6Dcb9SJeHAlui5MK2IsaqNmGom6F4plCJ1LnLjCEtOfoqGXbOesAavUfHFK6
dlVRJvOKthGoMQI6KZOCAjr/qJqT2UIKqDzHAgkZfVwiKdciMana9HwkY3qUoXGx
g1ArGGw+vVAQUDcXvB2Qq9NdD7bQsHDylflvYi5iC84yvzRJeaKeWY5hGOejKErr
TwZauzWmfpIBcgkUGx9yUhQpWsT4w86o9IhEB4m4MeMUVrJSETTbQKq4KXPC/4Oj
pIBeXI3yDtOPlQ+C3i9xTBigD/si8l4wIJm/4TbaMPGYrdHgJuox4u/lAeX+xMMR
ilShmxEpUh6qFGQzhRUJEF/BrfZz/izsYH07cuR3XsDmEy1jLEgfSRnrqwWjIYLQ
rJIuKWfc9UF/C4n/FWd8f4eO2r45MJGzj/BrQdvB0lP7uXIEG4c6/MKED5J2jtsh
dnUfiMcmrh3sC7kOxhuahdWVcfk5vRJuD/I0+/qwgMgdMwVFYxUPoAga+1d+Orb/
VZ41yoGkeWsUNi7/1rMexcJVgoAfbQQPIoAXk76aVlcFk5Hj8A8aK+8s8Kkspfqh
TT4hVPOJSTQacgntb4BuaibgpMqo82v6fbnQis031tiRPHshxC87un7DQsyJYLa0
a2KrKVV0Bv8QGDQla07hKaxHwKz5juM24F94EfScI7SEZhW1PdDC+Ps90AyE4k7Y
XvX3nziN0BZIZJHUrwMdvnh3atE2D04LFwQB/XV77VhBL3PsG3H4YRxDXDCZsZMz
ELMWUbd0vqFdJ3cmI4BFr9O8HKRaGPXLfIwy5SMVsAzmL4Lc4NU/jTvyop61mat3
ROTtWs9+p0+5cFjaoryU0xrBiI7Zv51cwq+CVKuUdPCrYUNsIp6U/6kdGvMi5iNJ
7LblVd8m4EKEP32mTD4ZE+6oJpEg5mKrcgtobZYquBTPuZ2zxqpUiktLchf6Jivr
uuSwW0NslvfhUItn2sdcVQzBWswq00RWr+V3siuSXtSk3xBOcgqbtWpxmqVbww2V
+byyGoX8KutRKMI0dF/AvAtDh1nk8+UQXcRO3Hg4AWYj8PmexeBjyk6w26L/hikC
bcaF4NRzSG/f5WRI+ipV0n2r+cj0F5Z9TpYjbUEVStVK376IBwflNWdgxjkeprRW
BBmW1U5FOsTEoCSGKAZLLW1w+aQ5XStboD3y/HC901svfyMSXow3fWLE90pSF6/6
25B0oR9g/Rv4jh+g3RrsO/1OOKRhWPfzb2yGurVd+t6DYjR/wSpMYBgKDlX2qr0U
NBiVCouTTT7I957ZBQ+AOjGS4M/hfWqT9yMdW5VSiDn6zgTmU+FFvw9NUpqR1f6d
hIvR+btoQFyjNuwTIvhaPSlm+4hXn0/AFZtNhT0C4Ht0bxfIHZwLSW+4sTpXE5t7
TnEbd+xtFowYkuuedwgoo4u12xO7cClTApDiVj4SWicVXhUjhKZyXntjjQauLFkC
XKOGU46UhOv7EZ099pTHqpweZ3cqvfeUP6riuU5G+49bFzJ9YIkUE4Oz42wE0HE5
K33QjpJrSpp4D5QXw8fZUB8COQoKHxY73jHgRXjqy+qoaESjcPSRChGz/4pgQhGD
S2/38e1Ct3Qgxr+JgHCx2+UzIU4smmOvTTLjSC/Ual0hKDvvxs/WsCckNKdOrV4W
2TgsnQ6FsIoEOtjN/E4Tb+NzrrhOnc8gwZbYW+dp2trRdjd2TuH6+coQG+Fw8uSG
Hrvvs6pPL2OlKIPTwvt88RJCzj0iDcMOTN+5yh9SJwTx1MMbcUn9/NbFZUPAm1pj
nu7nRBVis49E2zlK3yMq64xkGfa8g7bdZcYZ31SO9s5jMIIUuM3YfIRm7UEL6HO7
Z+yjbfSspCpfnEtVp04AkFx2zi1dZFB1CLeLOzRH5R/iDP78kIi2iMvdz5g9jnDy
0KGSwDaMLQP2Sx8i7qtaEvUtPWoo4HCOVQdRZNu6uqH1BExrpdsTst9G4Wq4tZKY
gloUFyQylsk/9Z3x9DEEX2eiUxK1nRFivnG5yLcxGtNJkmkySSaoCxqGueUH/bV+
7JIA8SicphT6Vm1o3uJtMDpEGcWxjjbKUxadkb+wC67bOe6usJxzM0FuCP0xR8mH
p5IuvcEnxmr6FyS9lVQweCRdTC68sey2+pLha0V8VquyqgiRQ7jJ18tf4IEDTHgm
IYgQslWuaeVXlHhQI5CzdLEaRJ9Ycgxfl9Lu/Q8EA/qFR8lr0DLpRe5ESkVhu0VB
RNIb1ec2g1qpH0DoFpTjmR8azGKnTsIne3DjH0rBW1Da3cqvi4gRbYlcuVl/I0zp
CWZj7cTRCbGEh7g7Xnz0bsm7xKHsetilhRzQSSecC5WYMB5+cULi1ol0K0jEx1x8
YMB/JOadUTcPMtYSLlmWekXv6krpc7gARAqKikxjylXNKsgMJO5J0jLK2/Kmdfg/
XzNtnVhMT2ZjqHDPAMaONKGL1XQO81epCaFQ43T60BOIZmAJOtcfes/1+o3F3l+j
AjeULn1cfSSXvOUFBdyc2V0Hbk9VDaHKMqMwMuLm74/33dP0pQTWQnIIlDIgPBIM
17LS47fXfpp/Mx0Q6uJ7imO6Bx6mOhwDK460G6xDWi5XgJemsav8foJJGe9Viybz
YwoujEQ6WiGyBMieEoZqbHt/+QaRlUFVcrgoJBOhjGLmxoj9uFyYud7puZj+ep1Y
MQu9smhL4CS3pHGDxjLZPP+pTufaf09kN1/HTd0evDB6IiQiTLoLl5rVwB7+lwZG
NCrSMG2bA2M+5Q4tX9jJ5oiISaUoCZbnC8urQwtrvmeexOentvfgnWKHtSJ1zWAY
8pPPbv7iKXdzORpfrVfIvVmlCEuZ3zxxqjq/965xzYSj2i/GNqL25EWi7lSjzKC0
yTDYpH/LYtnf+X8bPLB839sWEqeiNBOfQEOosoTlHEmWrk89T+m2wHMf84K5Phth
qNe7yAknqlnztCuuZ9cxIcS9em2a8OyBFwJ01DD0RNn2WmGqP4U0ogsr8wXo4K6K
0HbjXq+61yOckNRMpsuFjLoX20ok1tEho80KGJf2Er37jZVj8tQ8YcAWEDqQ3Mns
V2P6WjcKvbuVDVOHTROFpDtHlkzNFuJYIqAqH9dS/9yaayGJPD6kA07RNM2gho5V
Vxp/36fCSBjm8P8dazxMUs0aFWsC9kIsNjV96UAeBvcsMzS712SsxETjrfaVt53P
hvGZt/2mp4AYzPbJrSMo4jr7MD5XJdkx6tAAXik53pEmS+C/hagDe/6UM32OlnEZ
XvyzkCpsaL4B+pk3JJx7t14of1nf0T+jqQj5WKRbToE0dbbOVUOwMJyKel/na0uy
6YQfu1880eZGUDqto30A+TJcSZItmKnxOwc7nGxKX4qybXZExGj0O7j5iR95oVmM
9KhLnUYZoyAtVjiYbXGuXjLFhUi3loOwNwDeF5v3N2ORGRuVC+29Mus4IknA9Prq
D5LARPQdWwNiLY0JLrl4DCMih0prEMFne8pgzoRGqk0dixrRuP/a2SVUM40/Wcll
jl9bv0lTmW5eG3CfKk0esKicELNrcwnOkxtmyzLciBUw4QOryjq79X5pfTMEzElj
5fgvepJXrsLeEEk5biz4T5ak835gR/saXIyXwcJe/6nVDvhnbqC8qhRcHAxKsO9n
bQXf+KGjOQKflnrqv3vh3l5OWkzEl6nAKEPWh84LYGcGQvgIQVp8a62NcwkFMLw0
1S2cvMEWP2eNicadL5anezr/+HxwqqVmoyAAgUGySqRMIAIfenLOKXw7ipZS5C5M
IB6AJO0NPqy6pMm4yQRYiNUC89Dp0t2qX4FbT1i4d8qESAH7FeHdY4qLcYF5e2lv
Ilo1u30pvNBPt4o5wGXONsjZe3zgx4dgYakaLKa1PgJ7YMkOyhxKmuytGdeCzp7C
kFfnBXKqZHgZWlmMfQzqdsI6KkFVgTFOhajBr0+m5KKZs4PjM1UbT2eKHQavXQXu
DC0u7pKD3n5ukQQ/oEiRGrSyigTCoUPeHluZzIdxXxBE1QsIqF63N/qLV6Xg6kXq
jqb5xf0gP3oLmIZowyaWvtmkVmo9a31T7VJu0K62Zl0a+rZ0NS/ReX/2OnXY1WZo
y44gB4a4FEL6GgrcF2Zies9CbBCyLo1CSu2/V73y9nTHowBzNbWCuRiYXE5AQ/5X
roSB8Acm+Nm52bNMnWe/dm1Mcd6S2J0m+hz/NjRjLfZCp/avB5zVJZzm9FTiPFzm
7P92PKkc0cs6YZVQdRTL+47r90MBGpIJI5LCJ6IB2p7KnW7M+K+qAcNCEmRF1olT
euF5JfXCYVDu7Eo44+p7fDy9v9oDXO3hY0/pRlal2JIy5pzzpffSIbBFM0dPzLJB
4kmZd5h7kLaNGY5Ynk1T4AYhio6sGijBf5a8fDDok3ABj8LqHkX1NS3NQLzcGikF
1vWdK7ZbuccX5XjLUTnSoutYJY163/iNmgTHdh+wz3nXxtImFORoFbsP+BD6eQLw
ux8qqdYot4LzSaFVwKjihh+pQKj1pYYPMctr3I7tVtOxkmCxAjALXyP5Ldz73iJs
ZpWhK+37RQoAHlDprTI0iiVzn1w7h4GgtEp7ypo0g2cIw0pH6uOXN90arh1Skw/J
NxQZ2z4xJCBDXWyu/IZSIHDUUpPCDuxVuNA9PfepAMUiy7TIavB8vlstzJDnFF7Z
Kl0G2OdKSU8zJubxBoBjcYNffVuU70mkmYqUa7kLNrP3ERXMhbDDcC4VVGBShInK
QN/qjXf1WjleR05TxeD1GzUXRgkmX9FON7LDUJayQaElsA1uQJQz8oleGkvtntVQ
CcIwOkHae50As1SO2MqHq2X3vFRhD4hmZbO5idTwW5Iez8eUpAGeB25wSRwkyukA
aEfdI5JR5Q+q43mY6r4wBkNd3Y+tdEkIT/LxEqST+2PA1+dKCXuvkJUmew6Nc5O+
lRLacOEQRxSzy7inFYJ+Q/NC98KbSW9GTeZRhbNLPdB+KcSk81rRUPgOchfP2Xec
7C34yd2dW+De/Bu9+R786O+aGOPmb4mkPTF94P2z/B7aAXHQR0E5EAiuzxY/9bxm
c+2MmRXtfSQBJYe5pmrjAwQnJvxguW8nJXUvtkW+mcxz54eJ3zFUJgjLx2D3Kt43
1ZvAWEgIDcoTnrSkQiS+JB7GsW9boQZg7Qnx6CKzmQm1GrlHd9j/Fl3rUUYu4AD6
+qvteRvmLV+HcAKtValD6T5xCE/Gn8ulOOMf+QEZ7910USKLLTe1LXWv08+syJ7k
k/TLyskWV6c3MIePE0o0jHad2xuwB1OPgBIJz7BY87LnPOydrploZAIX3SJOtGvD
/V9eCARfMLwSYgK+24aAxX2sejD+zw2DoJ24Lixq+3CiIeEYldlD2+IN7Jxmmj/1
2eYNc+yBRkniB4WIBG5gb5S/jLfUYNLhyX6n4ZkrUWENXGv5k0iedF/uXLec6df7
KmerXF+yfIlzyXKriTuIE4rJkmh1AXlf2HWjVmIK8hmXgHs1pUTAvHwURpiaKxWv
FXTMrXpGzMbvdgKT6z2LkxOmV6Wixs9vYSxzbr9V8atMHvCpmM8t0wHQH1Q3MLsK
me8MLe4fSqaa1W3OUcgTqyOKBSoG0/QtcnkYZB0nRlQiKyG7R7BoEhMT6gODki++
KQp3ZAIUSh7cEfYR6OwQGVNgygVV9fx7B8P1trSbTGZPaqldkeVyGLDm4uqFi1j6
Mn/8eBnmkIeXJeVa9XW/bOT08mNUqrloRMehOHOqmwMC5SpyeFur6vTw9O/8Pv1s
fOsd7nWI554xsjgHf36KTmvNrS9zxTOad3nKE5eS/EVO/P9UaeaUyPBybwqorf1v
Axr9kF7wC00lsYvd2MznzMXhW88b1Lm1PsHEJtelZdZ88dAJKBoY5OLusat79Wsp
CUbUVVkQANjQKQ1cwUP0ORKY/FQ3jNSimE53tsVpiBsfO5xZxtWQ0rdQC+tRqhh+
juTI7CzasWy2tVMP7UAdzYOcElPQ/q+7RI7FkMaE5WvgTCBjps0Kx7mmQ80VdVXF
O5d0+cRIog/2f8KEeyX0tZqSOYQCZM4Bzjm4csp+QGcMauFdLCE6VZznFNc9WNtH
gqpgxd5Mjwv0CabjRFG1InjfCyQi+7tIQnT8CHn2vpBA38AKfjot2AOwQOOMZ+Jv
7hGHeymOcJzW2/tytwEqUoKA2XxSU4B7VPXuqeFTrYHCIyHfS8pgYqmb4m9GbAsJ
8gmVRF/KNkbTIYubHZdGgQ1I0i7IX8a0mJBb5+O/I8gKkbdgaVGPyGPrHlFV4WjD
UnY6oJCk3Hku/aytAjrm/WNJuq1OuZ3DvmaeRRbmh/QoIMKuX3y26tp5WolwMyhk
5uW71veTtGyiTwZv5CcYotNmUycE0sAYPCASzPc+260vywF4HQvhgoYLmehAMImL
3Gtn93gzn10xwT9NLhEcK0b6ZmUKfY0RhKCjdjhdbI+KV3UojuAkEr82omtjMbcw
LX1iwZG10JMrc+Wz0WypZ5COM3El42VSAtBNHgLGo24+LRfDukZH3r7Tj5MBppbk
1DZdZ9D2ssyRkRE3QOhcI60QsrXdvZWcpqloFGKi9eG5bM/OmM2SI76+3TB50L7k
GkBpjVhUbwOk5h4vEqeJGRocZkCBlPhe3JX15oy0jBwRVsLUj74xiJgC9WLSSiYF
HOnwbgNOj21ZbhgcR6R67ZCcHYBGoc7zIcLzcpTLvfimEcaAQCF1NJmeJk9ihFeW
yQbIuwNrEn07mDsPQhorx/3Nw+8dmPnhgWNbbAHjA2lh73JF57f3MgGn+h881lTC
ld822gnhZZiewSxs2fpa8qz6c5c/aZbGD9FD99udJHn5lQlZ/a7BwVIBBJmPD1uq
suRSzzVjIG4869JhJZIlVcPpHk118V2/RylEI/vxfHmnn4/duyuy69+Zdniq0gBG
KUfDQca/F9JruZOLcnmNCQ7HIWrSSprEsBI0ort6YqRJTw/V3tChD/nHKWORQzex
2vdhuYBx1T/Ln8+40anYMGQqgzoH12CeAC/H3NDZVoh2hMH1+D4LXPi6b93ITOmX
FSkcRoO/R+sjZeUvBexatx5nSVCvX3g6TzIhRBd1Alur0Hrtako7/fAZ8Y+ReTih
gY+2oZgQjcAV1WDtP5wqCoOCwm7xLZE8hINPLZ47iwjkiZT2cdbTiFeqbj6Zh9wm
lTe2//E2QkHeNIx4kwKLfDpHN2U9jIhdNim81qcBpX40adk/ITL1qR1uabHdjEft
8WzsKYIt4FhE9nw5VN/CYgEZ1SSa+z32Q3HQvklwoE805lH6OHJF+ulX402desDj
sEPjGEg95S3PXiPUFe7Irxh0+exTF4u6dbIypSCUpG0XsMCUz+0TNab4yKe03m+Z
vih02vWyK0vfNS3kKg70nr1uKLlGlApSwWJ8mBjE6i9HtxQ9OhLpl1qsfDsctY2Q
/gcoR3u2imKxlmHeqjtfMga6UbgN4I2v5m9mn9vrzfoGg2hsrWbtprDsxRcPEqXZ
XPkYqsAbD5gdRmBBdq0x2pc6LDCiGHicTjAfDNAK38ITcMtLgAdAjcOgkE3wecED
A/0IPB+ODYBGG9UaRRXyLS1aZLGVSzM5rQY8Dej1/H2x/TSHsU3GELACgpVY4n1g
4cNkKOspxlqaHIQxE6feiQsMq6KsOztkBjEgfhyojZBleonXjGqsjC2RSsM2R53p
aFUk5SsWpWUZb4VMTEU9ZDTwmubIn60hEArqld+FKph6JNgTVZlDnRvwvKKgSGVb
nmXwEzn3aGZbaCTP32LRtaC5He10osPhL3xhNP2tC94ly3lt4WQWb+0mAoCzMdQF
uf9EkO3G2zhvvdBYx0qLVuLeFhPr0sLy67AzKkT29sozr7P7OV4nzmv3+Vhw00XL
J1Tdb1+la818RPHztQgT+8hEPP4h0axNsLN1WMctD/ZuCvzad8MHF0U9n0wsPgAl
rzIx3gBdXOMUVmU9x+osKjfAiIkZVlEFrzNeuoa8m09WHzmS4gjVRZH9Zg2pR3Xk
xCFmWRBzOOxTAuEVVzDGfSkdmuJcIi9y4a16uK4rH10cms20ey+kZ4o8ENvCcZhi
wTiRArUt7FteoWlE2KliNMGRbHCFvI9jXywjG7jx9RmWPuxIePGQTnIXK9upZTY/
2ZNZoK/Hp4Tk8uBBCMu/w6lmOjpyBSBX8Bue3E/orIS8DEsE13KvJKdMAdbZOYoI
ZqN++I7BT0bK9wo00fnSopcqAb8DHdc9V4iZJI6LWWMnxiHxrf2P9eI06TS81tv2
J/NOFFtoUwRUIsVXjvbhXKfODQbpRFaRpRFcaH3x6omf+CJl/bCaGIQWnoRvQU2+
uSuzN+YwR8FulSEaPLBeYHCm44dYDtO7QlH9gSDVWzQDiUprr1Pxh/qtyqDVLVp1
gfSO6mxpaTFEnrbYXXoEM7npC4YDRGWuMZyj4G0wzkIfrre7XjKK/Sfc2+C+V4xW
vTxlXOS2u5W8ndsgwCuwEsRw3j9+1N1wUg5SGW3JJseoXgXDbxR0+wiTzgwkieah
DkOBe4YKb02ZdmlVzmaVDbGq4eUEFXeqmP/pdBDRh25PT/38lxfHcxXOSmWirxP0
7QLmFdm1Wpa40St8UZKSQ8KPf+bZh77ii77ABiCLJpES9SFVBEC51mHmlxCqqRIP
xNoyZqxLBpRNidm5POGRKyHssIQQr3gnqgMkaoW8td6maBzoZ8IOvushFic+dqDQ
mo20YlcqNyKhaBJ6rcJlvRTwQIxTty7JsWWQmjfwsb8Uicmi6N4R+yGQRv0BZFtU
XoMwvABKh8mdDPhCXDBLSO89P5FUcd0VGjjl2cr8eucPfNNXv5Wli+mdUqKV5caP
dc5sUof8E/sxZZB+y6Xo2iQe94BvX6L8UsPKjw8cCvjJrb8yZQulSe+orikZAali
t8vPnAb2EySUsQ6ODwAGMUYRY2E0Uf9/PNEcIJK4MzY059dKRnJU2yq4Vw/04aX+
9dwfZNe5JYn+NV6Oi+7OHOzmdsXPScx6lv8U5+faYxwcZ3ourzxdtdGegS72RSWF
HNYUR5o+mC+oSoMVUa4k+gqpz9TpKb4lPlVDhy+dewzszolpc2X3ZZm5tgVw93bi
mcvhNkaZDIcEMlQFWpoMvuijzgBgiTIaaAWm/50zhxTVTrAbZQ1JWrzB1U5yTPsz
JNlR+SQNci6s4HW9/+fS5NoxwjrVhw4vjGNLWEhWkuPM3Uhkmm29nGxq5yX2dvDN
ipPnl93/5IXS18gooGGHQKrIF7lVMVajW2I0Mdr+Omgb3FW+WvJEHp2OySWEoWTy
pflqEEc+9pb0UxxzyXHKGX+HWon2OVR6vuli9iSQqSxFt0SH3+6BXrtF1p3Ez7ow
z68BbfRPEEWafmvmu6Klu5pLQkv8mBpTNSPyBLshBCN5Y53/Ku26lnO6meZuPA5I
WNZjH6BE6xW9zrBaOI0oP4Gbv1dWqIHSjHkfyupewMnWFkGC7L/bt8TvnjBAcIN4
qjluWXpg6FIJZGsKihNfhoIoeHJZpgXvEaVPNT2/fMBdeJwReG8vXbRPmD7X5i5S
++M8OkfFpw4TiMMAKl72r8CUMsbLqL3DjWgi5RaDyuYcRjLAH3XtQxU+vJQfljU5
eMUvjbF7OAc9oDCd18/8EZvxXbOgWJ8RcZv6XEEm1rbBi0GX9YK7YiX3q2GttXRA
jHV1F7c3W/uD4Z/QD4p/af1I2mGY3kZGwZJaxt7rMrKLS41MLMqQerIgpKEhtbmR
0ianrtuEfxsM+IXR5YmOkblwVl6f+4cX2gU6ykNnIwAnksDgmtnfWQa8N6qAQseQ
ctq2nsqJJt4xvn6/8mMPP7BwGiOlPxnKaX9x6K3gW8Ldp7uUOA8FRszkPc7MfnJX
ixbmcTzyGkK20LiErdPyPUgwD5B6wQPbQgj346bCANeKZvHOLMEKhqTpWUgi5+wz
kp32w/lt44qD14po2TwstTKJ1KHPfrglJ5307OUS2rz4wBJzawViyrnAuIUtCgWh
0y4kB7kYHNgk0TAq01SCwlmmSs4D6WqNq5rKhVF5j0o/FQ5Ein2B0ATpuf1iT/Xx
Jc96lREGxrC54Qtq6ZJoFs3r7VwIvM5ZQELZE+GzLZ8uWN1J151Ac17wGfRdExcJ
bSY5PdjMyAeibOFdy+TQOEF7d26UKcCl7SGdMyhiW/krTohVDOnQc0C9oZ5p+aUw
pNXAfABYF50miKC451Ekc8KJR9zG0puVSSAT/5EsAU8W9QgB1ogsuV6J62s/vbuj
n51ZKu8+ZRW/g1nHmeuqyQAqQRFGqk9eJ/ESd4Vi7DqnnE8sGFniG1kMc7v56RtG
35PWUU5wC9qttmL/0YMtxFBfTp19UTtkiOZfdC+tdBlqMTkMWC52VPlL+KQszViF
lfYRXFQIa+tNetSlnTpTvsDAuh4a7713x6dGnulaXl0VoYpISm/OhcrsgIUY7clH
Usd6gfTspj+XZcS4QEWn/mlLipXIUM9w5QDX5K1UCB/KnUfqRX+yNV1KNdxCC/jm
npeN3QggYFHRWNq0Z6tD2GKaGwCApQiRo36UxS8ETXEaGZ40yxCzqYz7pPsOx9AS
pgsArC7VpZPg+UmNhpgsy7C7HXVcNhU9dhlwIM/jYcEx9jACu/R4/c4X6NS7ZKoB
l22lStRX+cq7bWEYLlcO8BCFdboEe+5j382YWW2k8UUeiD8Sv3TvBV9P+5vt9Ggf
FitoxNUfBRE0LAczaQIRl82fUAWw43HuWWVjuYZyONRgqcwdz6evbt2DD68wq5XB
miFOPSC9WrwhSRpb0sEP+75rUkhkcBBuQop1Y7IJ/vMAnfYPFqB7pI/V9uH1qZPe
7TVOf2uker1VwsrZefUMXAv5KLFTwoFQJXAoo9Fho8pfAs1rKzFHA1Y+OTARJvDL
EuBCGZJ7bU4KOxSECmScfmpr6IdMxhVcx8++E/eKFxoZdkH7feQAwjWmAQCTnxmy
SQTpW7tr+M7iCk6I5qsFEHcV/HhmLib/sjGqN12Fzk3sPjMFgx/dh+oJMTuJ7GsV
AiHeN40byM7USkUGAKYJEZFIF+B8zZQ4CdmyWOOEjZqnQ7Eal+TRDNV039RNozE0
g5DxzZP7z93f9QHgoXLxGprJu1XWYmPvWgOYy6F173LV95ZGJ1CFEQcZ+BqQGGQ/
MrVF4X6SjI6VaQCNodoDapdmjBqMEspeq4fg7AfdI8CwO0Kr0jQJVisVxMfy5m8T
uFUWS8ai7ji93bJGFDljfrkl/wdUiMFzqnbGlg9OfCWzU4fVdlhM0nu5Pf6w4r2v
y/p2kljud74FZKozS/KOwZP/K5yaRxVX95c6f4GcTV4WhPfSeAA1V6F9dUED1kuE
xU/hzp0xiiqTnwIwgxcK5HXdv7lnh/E/YZBrijsLj1mr66CBFFsiIX5Z0QlIM7xp
f6T1sJA31r12jDcNNTa0XfZWf3H+N0L1Pjw9nxaBQCa5j6AIll2pQOXf4PxdudhP
szhseRbUhlvXhe4t7rvVvd//qjBXcKdwrmYJRspv3uHnlgHmkxvYojNjAN9larkv
Dhg6tSxRQDausoT0Y3knigauTEOQrOgxzG3PR5dB07L7IOe8bNmWXXdXvOloFhPN
uchYnTwxEeqGpJVERIRr4QCQA/qsrmfrsJ9SX8gDNMZ7FdJAEHpOdPH2PUiXxUHu
GAMlqzlVzYIj+wL24NaHYOUgGH8GXcmaKZYuT0PzPnvTln6TTzmEZ+n4Ze0r/oMM
nynnkKmo5nnJ/Nomenu/juvHrmY+kfYrOCSitxn+G2bfEM63CuRWQiUA23aL0S2g
hR1gCYPASmDDQadImN5R14wA89+pGx4JSMAGzkj27aEOw4K5O0AdLnracnjVYJ8l
c8SyCQjseIg/g2qNYy8nZA1Fvyx46SgH7458pVAZb1GCHwLEFC7VnQPMZKnbU8fO
NmIVO/7KjUwoN6vuleuyEv7JaQdl1UpAtjI8lQHBRRid3aWOuoWUbgKVX0Spx653
szHsrvs5bKbm2ZSaXYMQZl1Wxd0NS3JZ0mAESeO9mCPqdsB7s+iEDT81Evsx3IAZ
f5If7y6SkNdu6MmTqSqr0whum93wzSf12cQ0sq4R2szCQhnQBTvRTOz2Ic0ODKl8
/cWfCaPtGSf4d4O9Uz5bTsBH8uEHY98F61PsumGt0P7m/XUMDcCAH9QC+DyrPDLc
UFkjVNa4VxgLNAB6+EhHhdb5knAgJoRu7Zp6F/V7J+FSmqxzfh5aWkR+fdnNzprN
zusfkggpShOwziyv+XzRsGC98e5f8owJR8Sk73X5poGKpe1F3ZiD/ADJNXy2az4W
ElTRDXMVUXspSjOgjJssuVA3K9OKGWG26/R8qytF1+7TQlris4HNMFo6zvZiqZFw
mGozzFAU9lDjm4dm2m3ihGiCb0MCeRhNQ0yN7/Pqch2ECej6xnSB5NuSPuTAZtQ1
/0u5t+7iPDnTZ8geJbsCep4HsmlBh0Sw16Wu7Gerb85ISjyW5mBGIIT+qlgEZgqE
OiyVu9nK1bB9VBaiZ0zvspQJwdyKHI5H/WtPz7v5NfNwu8B7aiv/Qgyq1k1Is5jZ
w6Jub2I3RRc5tSeEU4cf5V5lymre1G1L1Kt1uahiDgX7W5GdtFQbBqMk4QIuLrc6
nZY+FFlmKc7e0RbHji9/vg0z1KQxw3ysMUNL2EBz9JxI4qEq9NQEaV/cp2oj02vg
39ndaMXwxWDqg2qS6Nzh9R4U8WS7eR2LEyt8JNcl1TsW9sILo/UJw+KCS2CaSQLm
Oweuva8aydGPCi4cwgqIs8FcdUzB8htpqn7RcUDQtD+9twI3/o/DVzpDZC7r8+3H
1RbHbpOEFCeq6Amjix31N6VdTMOoV95lhcgl6M7eDFbxZeYuxlzjC5i03WILqleu
93epuH+jqJRaYmpFni9VLuCZrJF+fSwwoTDCivPPONgjh7lA0YwH/Epwxa2XokUA
uOrPXqxUYVuePRDY3rQ4OlO48Fmh0O3J07lJJ6iM670tKte49jXkom6aK6UVMkkE
4IvNheyh5B/CaNmTJZOgc5WhJ990SRf48Ule619J3GA10tghwwIudaUWnz/fgPt0
Bz5bSB6HGgrJI0PWgF/HCExQgMziL+ntPqeJsPoYR1A8qYRaU/iFMI/9b9gvurqH
aeCKoLQTvunkypL9aAsj0BHvKeypm8GQPWqAGSr+OYghR/YBWvbz3P3mVM6vPD9m
y64A9IeZ/NSPSd8J5KrbpCOwnqCUzMI9+4g2JedV29qfdmccVXxgPOyTmGVYuW1J
P9SkT4Kant6/TRXgR1lr0nTBuLKrFZA71pYVPCCPv0eXHlrXyXlWYvz/HWczex5B
FEfsHtrgzBfyx/nLEMvc8KbUs8yXMtqZgm42lIxkp7LU3niBjP2HZFFRTEBYzCcb
rEXP+8gVj++Z224bHRb32LQdb7/Q2m5T0NkcCWO3Wfitbc3+t/ljzhkogdMJy3RU
hsUHxk+QKsCpN0OQ6tEULxxkPW5i6DICwKC8Nvl2UrV4AJcSzuew5tm6HRNtR0Ci
OmumhWxBmoeeP1CJCD0kCOrL+ip/dBNjUXgAW1HaSfJpvwJ67bWcjBXk9lXThCXu
YX9748ikdxXrTk67mgQic3Fkc1Oy6dZNmB2EVopl+BZCwtJ07rec4GzJZCzFRCSb
jqInJcUkKIznMrHziT4fSC2ThleZ/1aprqqiA2FdxdShEYayyQ5haUqAOIeNiyFA
Tnh1gJA7SDKtijzjCBa4F4H7O/gr4mw29YAf7o7vCnrJ67z6+QR4bbpTs0bocexv
qOV4hEl8iL0iK1LotXpoN0aOnGbS2m16tlcYPB0cHnRQxVuA3kcLaYJkoMqZy1sC
OBq2P8COM7ptgw1N10vbAhA8pZ6nhsZAuU+5I3ZDUdsfTudVzz8GrUxp46vGOyff
+Dm9I2TS+04DTB78Hy867h7JagUqu6KuSpVD8o9y3dpY7Tf5bXYI4WZ/mi+bMzBh
GH8gVbwJjRqkQfpjPzbTSzkXGbT+Yr4wDAnSmrK01/H3HB2gJK3RmJZBDEENlFl+
8IUxJtdPXPgzM0j9YlHQpXFNcC6mGyb4tHTAKN9UC74xtQUWxIypGidqdqcSSuFR
FqibhwAJJuOEMZCK5Jp6d1hFs2FyFpfCCd1ebPZQ9TAfsYY9rfap16NGeE1FMVS0
v4rO66Bn3qRpJvnvc+IG8MhPnSUMtWEBH6o8aMjOJ2tae6IF1VTYr3nHRC1oPAOS
IFKuU+pQCiUiW/SDuG22yP+6muxn7QcPVSRUtTuIIX04VBwIgCgx59Zu7Ef3ws0B
8nbgMfIcoaf1QrF/PnM2w8VHfC5oZW/al57GrVkAM3TSsMHNamn7YtR1sQAY5+bb
SGZ3iAtkhwg0ATfCJMwsOh7svUCtoU3nKDusA2RFwpr1sppJ9JcgbME6eu3BOlqP
iyGp4/pB00qRFZaUjYbi1igcM5Pa4Cr6PCKu5pVVM3AevuM0XdosGIVuhUBMPixi
O+Iq1Wu23m/R2Hdt7kmS3oZesWL3630VUFoMRgsmY83zn0ILnEJIKESExPtu/ey6
GiMufu0NXn1JD9WX79+ZOho8bEhJbbRhQj9wNsUWfvF29DLakS7LgL1c2IqCyskE
DXh7FcgyYAmb8mkPisW2gL3J90o80mM2hbdfXCfG8jBk0FVGw+D8YGEB/HzyjAsw
TakY94BFK9akjMZ+fOhYf9oo/3cJFi29yVggo6BOM01bw9oNNwn9N/akTjYGUnsW
a+xYERa2sy719MeKlE+59miBZOoAtoKUfgsKnh4V2EI0C66jyC859sSyC3YfeBw7
PbMYyjZ6HdA3zUY+3EX1ELbcYY/rgoU3e7/2Z1GDu3G+/F91VJWLLBmuLaWdJwCP
O0XLNXYdGoKd/MlZc4VYnY00fep7u/e5QrK6xJ9r9+MxQ/zf7Y38c2JOtYUSVH7e
Y4iZ55fiVvPCOpzdgfRFiOE3O9B4dxs9DACCiLMQNs/YjOUgLrG+ybVuVxW4ZfXH
4UKc6hlKx9RW5dsfRPJJsG5CIN26tyfSB7DiSY/MDXxL0n6ZiVvNSRzZd5n043OM
KmH2VETIPWVlhVLRgajRhwCHnniYFuEkmXh6N45eegQJvgT0KK11xQ4ufDdpsLfZ
9XIBxmXu8PX9zRXXApEkrGsk704VfA/Rw4YNOcHqe1Eglbcmm3BJGB7G7YKKGMn8
wxUWv1ECWIvzBwvnbh5egVlDvpM7i5Y7uabz6Dxoc7PRtiCTgTwvLMc0xTQKL7Ho
2EG5xsn228MfIBkGwxBup/iXQfa1eqzILACDRHn/sOeJgPnMVf9EM7J4fQojdy8d
6UhuMewufO2WuTZ2f0Sm+k2/p1W0DrJYCmd2riJXdMh0dSF0eaENwwMSoOUrNTaA
MXNu1PvtbXkWDsNyHnxDXGVu8oKnEUJT3ic96kSqd6bAzCqCH9/e+5TmI8hVW0F6
Gmi7qUzsPKrjCBNiF+Y7JsdHHPZ/0cATMJXHdkfWTXlixWmA/mHh4kChjrv35UNw
HE3F2aDdJBNgeEa8eh+RO/05q/rdikTA4nyyrBxplxyuXmASyCr6e8Yg2oaRkbFL
PwgnlS9VuBc3XnAn9uAM9vXMqKEnQh65mXgSuae0/25m6zD/fg1gKWAb+AgW7tUM
nYXaiAM/cNt6KqJdIl0xqDkXYjoKGf9ZwNTfUrlVQ7nIZJMiwHPV3o7KoKq7rnRl
D5tN4NRwYHef7K2zXh4AoLg9DfD0yRSfNzXNOx8ohQcvTN+RTt8A3eYgz3em48eG
oQwS6a+teXomUBI1MfiYKKpJZgy6R82dN5a4FbHu7tXUJM2n71PSY4IFhVCaOtgk
abkE6AsAEPN4pZ0S32r6KXQI90Pbu9tT3WEtEcF9UdbZtcBv5f/PtUQcQKi73nyA
bklpaUI9p1jHDDIIIdH7fA5iBX/ndLgS3Ncd4u8uIpKEUcQfuqrfy1Y3m1O/9xf7
S+2nr3Q2p94G6f0zjRxS7vtAXLdWchjC+MRHcuoW417Vy4nrdW5vvNDgjmVQc0kP
69BZIhH6hMcJ2vrW4hofYyeA8lk/5jl85WFK0Lbho+Q71F5yBNKWWnDJcpGbR7XU
8/vMlcECC8OQnd23nIkyth8kqCimmYe3otKS4W4IF6dnliv/1SlIZ2CSAVwaijkp
i+P4SrlBFhpe6TZTLjbcCE8r3rSPVIvihIBvSnXDKJOmYJxNmxTiuad46Bt8n9HI
4fhYnKm2m5FTx8LQcYD5K+T9LJiFMGF1Ar8Vvbcq9AZwYhAK4H9TqOzRg4mTBkxx
y/txrYus7Y+qeXOJWP2S/PuUFbsflEyMQZN15VBVkuT/VHr91XVqkkOuoVa3LRFX
NyAiG4g6KoxqWWIRsbm0THl8dE5xY256ZZwWipEVxgMv3oOhK6d9aCdUaQfjIkAF
3EzqKMl2RcOOT1jEo6t1Mk6934ljAJFHVXG+ChGG8FVXL1fTy5YPoybbxTTJl5HE
zRwwIzpR+NT6VWkTPjG3lEPZ++8TSPXuf870i7sCJjqeGQa+oUSAjc4nZRpDWySN
yXQ0imYqBP3JKYKCT6Mvo4ZCaTrh7p2osed4+4YZIDRX6VSrVCmZGVkF3L7FUskV
mwWeBgqywCQjfSZ5tsHylevjIFRYF6nITEDvcaIdJibMWYfF4lJ7UF0y2Lg7YQDC
JjmiGV7BFRB+2dn22qju/lHrpLgdmNdjfbo4atJqOJm9fqQj3NdywijAtGwQKUIU
Ek4qDSn+vau9E8Fgc34tdnDsoRcE+xIlU5e/aNJEkikeP9XFhQvh2eWtQzAEQz0t
YJ2O2i5/h8bXcSx87XD/S6VVBEKD0P8Lg4lnhcn0Y3Do66Jef6K1j0F/4V1xpgVS
8GyclgJx0MDpUXmLwAfd9JBpuHOKKxmp/qZGK+07ECeJj0OTkkZLU6DOML9m3m1z
jpbbpcx8fWQ3/ab3vYmpkDv1wd9PgnD1PsL5d4KcW06dzaUSW3rI2wKC0NiYO8j+
FuTtlHEb/Zi6tyJ01fZzQozQBdNrGzFD9iAlNGgOFAJ49gtR37ls6esPNS6b1HZQ
R7hetCvZUyYo2+3Qt5ibgzJnJcwgqfI29Fb8Uqg3zWOXbvfy222sv+aSCw7nploj
oQfKwU9xh8H398cHHQIckvvzbUcFgSERFE4ow/WmnyjUA2sDBbW+R3rRRhYFKEDI
e6uLyjTgEe7bkvQjGdoNKlvDOI4eWVLYohU10dzhtH9df6G5nLWcWv/9DjoqS2EC
Kj9iTNuHWWj89b+oYuCzc2CopjLrjU+RvtzlV2Jqa3sc5AXx1MCJT7usohPjFuS0
a/EDcGVRPEeKUy+B1+xIt4r5ZkERKw2mApLY0awDTawsIrrf0Nfi1J8rP1WSsnkB
5ghaIZ1CVuJSsYBe+JYt0Y1fFI/6BREt9n/75BE2sskIam+w+R7+oUbSdwjMSeai
9/RBoNltad46ayzvQgFaJLYj8OiXjQwxNfswx24rGNxXG4VS+T0X4s7CleQ69dmQ
IC2bt8CT6xSYa1KMAsSNjDYQnCTzUr7qnBKxcrsPq/OrHMgNtx1IBMOLoHyIIRut
Ws6Ta6ZZlAFYnYfrfnJxw7OunnmloJXxz83o5OjOSu3U9HjuEJqKk2Q3CwttygZx
EmFax26RiWe3mV0jfDAlv2A1RZt5JOw8mnI8WxMUc8TSiRFILemkl20Mw/81xQ2i
BltesZ7OxRohryXz+prlJJYHBQBCnDn3zZ/uvXCksd/kZr4fj49FNuv7SyOeyiGl
Ruf0NvpQYlfo049JXiIBfU0vHgH3m2yUZuQC/UhfKdISnc9hIWMiMrljBFc+Sd4a
1E6yD26GeLe72xyzSSE7Ak+FWLPWQ5WLdRsVpMiyBnlluIfAxFHuQBox2c1z4rE/
lM3erQ0hOvovjNO2+H4j1Qo8lNxDIC5g8eWO1x6uJlekzhJKHFY/aTWWTpG/qiFI
1CVsxHoeFGtWTuOwhF1bMR1Bhwy0TSsCuVo9qxs1XTj6Ypj2FT85r6KSXcRUyUQ3
XCaLSTor176TGP1R6X8bk15Z+qhKcCt381xZ0NkkFkdUKTy2ty0xHztKQOK3qcCy
eopPrC6OoAlZiKULOeJz9dvrepFMJkE71LpG0LF+JIdOSynzPyFk7DLug1i735Cm
4U0r9VxVGnLIIwamffRzIJT+Jq8mN6yRpzjDtajzEvVmXWjNzOFrC7eIShy3bnaX
lOkgW0LLk55epqRvCAoFIvp4+kMtsbVOnO7OpDGuaIxQx9a7SoDcQA1pK+fP3Sz6
Benzmy1RBsPhP/74lERA38VpPzGeeVeC4I8yZ77xvIDdtP+oYHF/zUOZmPrHhDcl
MoaJL2TOiMouXwToCMd57mPeimjibQDSWncX1NPMuHSRPbz+rtDw0g+iPAPBpnMm
eNUj+jcOLvFoUaktk4YW+xIwC0T6omCiQ2ApwQOJxm1mwOhzf/rqKOY+RKQ4Cbw3
zLqzTqfAXNgea6Fs1Cwb5aEqRlyAPeBsrUAnFipDW4PwgUeNEvQgcBgTpFRD9H/i
ifF1mGJKTA3Wtv+u03mhcz70S/QXN5wtWVjUHmnsl7yqtnUQGvSphFiKkIVHYTit
VxBIInq4fjC7IK7vRMOvUPMV8yafGDcqba54de3Pv+oWFP1InBcyYSbPKMw1K+1I
EUJ3ANPT9EtF+RAhA1kkfZwxfLr2sHcfvvULfKkxeyZWS+FSwl8n5g9+1i4ufdI7
GN/MDs1F/SR7pL+8dKLIx10HpcL4xNehFMHmZ6Ee6ek8+wpvKIQ0uVJIk4HGSD/f
V4zbbOcuAXggc1sG0B1ibuA3mqkFwnI9uzfm8+i4Ie411MwMUKCQ8dLcYSByi16E
ZkXoE45d7KviTLOzJmd9mn82ulHWcn9RudXkSnjEmZJfzsZXXc9yoWrKYYsNaf0u
FhnaH1Mv158ZDYKjBPZTA0ChSWyzYslPd8cWI0Acwo93IgIk2z6sZYcfGIRbYn4k
lv/WljuR2dcQ14lPCXRkg7vNCW2XJ43rA1E+Kf/nxYDj7qNd7e5pu1ZbfyihLDNt
x9XI4VmTXI8wn/YkFcA6gNG67NQESwCIOH4K3uLlnPVQjRM5kPLc2/jiHVPjtZt9
AMdFw09IPCyv6uLr4k/aCzT4+n2Rk6taghbZ6J2DfZAJJITp36fv4NY8sfoB3oVC
gYf6mb0/jGa8bZmxuczuw3AbL8B1iCIuKeFNQIDnVGG4vsXGcJJrPNFRA20zqLSF
l6UdC05GYnwpPGbeYwceLu2+lpbZy9OWlERKLZT6w1fKTP4bAb6fx0dGJk7uhulw
Lmetm4fM2F9mV5bz+k0NtErAShmG+pn1XYHpLOl0wD1lpi6EOfeZPCW9yvfSliyV
KqnCYHs+PPtOi9yVceynR1KnSqUmO/ui2dIp2xrVX3sp355Q73FkwGd9T0EJRe1T
CSRrVA1b9YWN1YOoboYgOAs9sK+/pqR7/bUhpXvjHLw8qhkVE0V5XiNf683lZMaz
ffCYIhQtn3JUP13i7epAvc7zwBhiLNoxksOdTJYRFDCE96jHuEQEnBWdq4YUVMb5
pjHd3jpDEmj5A5y7dkqWQn+4DqIruqqY2c5MVsHLA4qtQdFau0nG28qys1gPyDNh
a53YtBkEN0aZ5B3gkpGkHYj2TvWUJcKmybQmLIOS+LDrP6fXm8UVaC0e1qZJFDsT
/fjVf46tzNm3ZQVubpXyXE58pKLScR10Z6C6IQ7J8KuLxrF6v9jvLuMRR+R9GXzs
Aha7p0audXEnJtYswF51lrhuibaeL4zxej/8hDKYESDi8fcSBPz2UDB10iOdvO0N
QjVxLQds5Ul9EVHLFDndhcMol4SBhK5ip7GZ4YkBXW4/vdaKNNjOqY9lrDx9tlql
7UqeFoHoo0Z8dsbUh0mOqwhF8GoaHzm4raZPDSo8JlBpbW8iD7mDS9ffqwEF6ALM
q4A0+hlxsLbPHC8U7DYGFLHSMtevJnR6vv2bfg8m5fZO9CiDOfCjXT1W04awtmIA
9TV/XqJqKpnAh86JAIZ2k/wcIIqQROa0xQthdEMrXscSXFaVZlbrBWyTlKQIn5Ks
KOCE3me7RpRr0htvA48AuV5Q5yTW/h8hh0+YZtkzWFHYw3C9js+bZJGOP+/3Hbwe
O4O6L/6x8JYYc1Kz4nhC2nLnPXB9L28ATG6XRcJPPD9G3yQXvFQC5OikvsZCi4//
ByLkAm7rvUJaHBgINaUt+lbB+mY7KhQ3dUR/mN7Hphmg356z7dKDlgIaHKrZ1TQk
xLCG8SynbahradesWFPRIqfDKdwkME8pLtYmX/wMiB62cTLyqgVAUsT7IIYZ1hQp
NLu++y78UmrAoWPxeUUSkJtkN1aca6Pj6W9TgN+R3NzR9MkO9XhD3NmcOsLrnH4P
qxMOnCD9Q6Q6H2xKFuZbpPLuXpULO++Mfv6T+H9C5ZvCFXQdPKjkGJgLF1HXe95O
ddKvxFjAi0ybCvgoDoMkz3t75WcH0QSUhLxjhLdplAY09FujmnblVELHThUhr2+1
GZjhJTsXlICQC8T0hvzy2hUF3jnNk7HMCDRwch1XA/LEL7Dfp30bQC1TQtxwOlgm
1QbpcVdSF10vWTvADMy8WGE73nN8i81bZgJSAx0TYxMJMiJUKAL6KI+VrmO/Lwk4
emSx1SSb0tIWQ2BrFvlIOvtPu5ARY9R0O4BbI6f/oE13X/KHE3bGZXG0UwiBc7gg
1jGCyd46obsfJfjuoc1nB5tG+3NiNfoRLInG4xN0wd81SnW/PBhAbrRY+rWbTHMT
UOSWIZKc5rXytGy7EqQl7hp/9aZJ+CUCOilcXer4Aw8JxhtdMfa6kwmoBl7n+fYZ
Z4ZSi5N+0FP6tuSpocAZc8HthXl2mE0ZFm7Ml1VyQ/WSWwgsRFmorcH3qFUHYXd+
anvz5fHdUxdYfBv9K6NoNtiU+BuFeN+ijoOkY5j4dTRwA3+YGE42ygsF7LgAu3hA
e+aglC6W8QQieRUmKLzhYSoHuiQeUevWKlFQ7y/LGdQCiywqhMizD82fCZL74uZY
FsA/+t0ZszPHjV8PqvhSy7gfoLcbRbo53+Tr71zXu/JPSOjRxN587qui/V/XkC/E
TIt7M1mtEjdRPSszdxiB8oaLCSLJsbISUvvYEDv6avB6Ld3d+lcuHE9arvZQYV6B
9NScrTEMAqJLP2JMrtigdf7ZNZ0vyAiskG8gQx1Tlh795m22PKH2npZnC2r2pehB
6QSlXMX00nrgnGp0odHfG4FQl0bdOIisto80bRTbsvKnABUjTD8w9nmuYrrG013T
yd0+m4OR0WORFcJlA2+pfz2WmA9gmmAxlMdQugxaEtaP2aAT0II/tl8ilDlSCDyn
wuJr/kebYK4I8cdjLz9mWuZhzZl9fWFKXK6FkHhVDolzT6Lkdx5O9fJFJrQTbHVV
+SieVEbJ4vxrIMy19rFh/GJZFCMSjLfFEkTnXbFWDIyUsDjY6mVvYJPvjaHO6n0s
GbE25Dz2nyQfUVMHdGox/httiqLyVjAAd75MbCcINihQVwIo+JSNZizmPCOXFJYN
0LQu32oui9kEf08/evWkG0lkdJvjd+UT8HiI9ND9FQX1HUHS1MTjHLmg7WdxGWAh
wWY8n7IKdjGpq6oTXsUkeZUPMmDesgGCC/E/og7cvPbQzUDngjrT+EQ0i31q1gp3
a/dkPnN4i4AQEP8gjkZREQ2EwHzfbFxn2ceDljIYEH9zTeL9284mLGbjJPpYyR7a
x0h0sLjTQ/pcWLhffYg0J6EiY58RuXXe0p4kFB3Sv5r0HfubfBciudkBPXPlVVFW
oMH07KH0ELmHB5jXSfOlDG9vGufS9e4PnSE3wISQbXGq78hzCeq2tSG44sXfmE+f
eoQNvweQSXEYvf11zyAWUxKqmKDKm0BR3kot00jLxBBgG48ytluw43fImUYsb5ZQ
RlufW7h+OIya7Bs0bCe9wXJwyWPcQOklFWtcYu4f78p2jLP/Dv8klZQdM4Mimy4L
3dyEqHX01mnNficajkMZ/JGVQ5XOXjBY+JcBTX4VETWpgY82P+LrPIbm6Vi9AI2w
3JPtUm51a+BA+r/ORWswllxRorQ1w4To1hYDDa6lPWl0RJD9fc1Ws1orGKHIYHN+
FgakWgK++ndn9W+2VwF6i48fTKKCv5rZiwBVEx8iSKLqv7dOcLqJ18THXZJLzmP9
D8IbbCN1qNWtFO8eImhqW1MD2NvRQrD85hS2G1ZwWvxzPJkrmLfzqX5+7PKscAFt
a8YAg2yRaQ6JZySkCbAW4g==
`protect end_protected