`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11040 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/fb5NMnNt7XXpoSdQ33FnbLsMlBTL82lxNEJ8GkskxV1
BQjF9SeGunvVps3in368btKY4HsNin4ZBtE34InWbl12UjzEoLJHSExVHrgVhtNA
0TVYlFpwp70vfcwjPX6UAAJ6vny3cxfFsc7jQSGk1us6onVMOE77dUQseJKh/jio
HgJ0Vsg/lGpTwJxlvYJH4eq9otrid7nBvh0YtSoW6pFdKSr5Liy4cnyvMj5BBG7B
3u4aEKtzZqXloJXdb+071nQLwYLjNn6Bj19pD6e+aqwUI7H+CaM1COxkWqZ13e6F
AYXJsi4dX5i9nybv70ZTCZrX+rUYsP2UXWouysTRDI9kQES8x1xBuht34dfcJnPy
Bl6mCRorfoflRqkgO8W4IMsmWo+OXfEj3bPr1PzkMrDW1UQbMLovF1kJpTYzXHFS
aIJI6HAzj1l+sy5s7wfmATgqjjgQouDCEwFfUBCJoNY4bbekkKpkpIKXJAJO9tUT
ENkYBDwqxxM/G2FWdpzzxLDIkKk/qw4dlyUv53/779URpNC0zleWLzjjMkPqteWs
d6qKnjbdWYSNjqyDDDK97zyezQ6qbEO4HW3/n/24aJLHVsecZ3vSbYbrP+6d+kCJ
Y0sokimHDi8fWsnoSwA1nEHmGtGVKq0kZ64iv6dW29sYoX0F4KiUNZvFg/flsras
Bcwuy5Ue5v96PWbTxRFWJlASNMFLohefn++Y7/7B+adihLn7sCWSkjtLOgUowQl1
6e7u8ScTGWJcTj2OROltqzZio/s/j7l2f/Ew6ErD9370SF3cXKcpJyWj4dM8xmWW
gqjyyFvDt0EExxTXbgHQg453ZG9qOA+lcFuHYwVRg2mr76zCZILlo8t5zqcBhjFY
fiQAZ1L9anyYcdnHq+blp6+gA8hYUUXWAEH3OlNhdFxO5IC942LVvFm/4TQGrEKS
eJE+tEdz2mYEidxcRXzm7nvBZpqAmx53gq305iFME+ZGqAAjuHZ+1vSgYUXxepR/
zZm6AK+eTAMhzH+cmQlV1i3xDYK8LdJ0AnVn9RTSPhdsB9nDTDtvhgqgLGHMzGZ+
Ewipx088x5w92QNdlbF46a8toIL4qPukPOi1LAc56h0Oyt+vX+WuMx4J0TQ0bdIF
y+EwDOGj8820uRr7n0wMg1l8VLKcuAr67PHgIJx0bT3JF81LFtUMaZ233Xl0diYp
ZrdEkBG9OaPYR3GwWnq49UWxjprF7H7I4R28yHlZGO2S0hw4TFbqRgRliTDTYVG2
k5aDXmi9C75OUz4pfdPy/dHB6D/nHotOou6OXZ5zIPdLZXGuN2dp2gg2SPXwBDBQ
eaM2oAFbSvQBXW+8RMjjJViJuYx5fv/TgRtix04b4aUgDaImon3qVulE9K5VlKLf
+ttwtSCZmQqmM93BwJ4czs1QGAVQ9GkIHzH/5MeFCJvojGs3pZ0gCZHOhab/sLO/
+OdX7oym8rqNQIx+/qRs5P5u7WeYhQJHNTkV/cF9OKTJIpu6LJmD0POmkZJiT75a
f/Meit+1HMYK26rMFBp8RDF9bzS1XsvGizbh5+SvZZoKCX1p+yAg0PwZPs/z1vb1
m8+FHst4W23nChqjHEV4JQmo1yGVHoKOO+FTeukP5p45XE+C7WWyNC8a1lW7dAne
CH3XpWgdJhnHDGoV1gg07DlRpuX8MYZn4vtpVgXzy7M6wGzLQG6Npa+wn6hNg4Ci
k+6/QNo1YLAydMinzkyy2EIO0IjxAGwE58aPMoZ1Hu6I0939GiwFYKsnSNqVESVU
PQk8JQi/DLbxT7Vt2Swu6c8JXu2HoY3Femr94NjaJotgWWRiUpB3XQwpvYBH61v4
L3nEYKemc8eIyHVJRl+UqhJCgXhOj4K26LBNWeIKE7fpdDpdu5nG1xaR9v75ioY7
LCS+s5OpLTVL4H2vAJUQ3Bt6y30wYaThZfGD6Tpvydas3Kiie8JlBpFBb0ZFJXwU
2/VN/WPsVPT1ct47DiE3nj0l9jZWz+LqgZIkAUI7yKHbEla80c08MJylTdCyZSPl
g9DjBK7C8AT7xigGBBJk6jJwnv5lj4VvUSAEpCWI8Ho4bIAlOqLBT+dYtqRn3+SO
MVjOxyGGXBN+kZJ5e5MGvnkbzqhTv/SCD1Iuxz3BckZqA3nnCpmmthUB400mpz47
0pVK4isrGlgTA8IMQ3+g6md3GvZsM+eNuJm+b5Pa+SNTHb1YneD4JBBAREw/PT/k
mCn7a1gVi3rI5QAwy313oOl0BBtnnVL0d1sCIx2hnrU95O9Hwwp1YYFboSXOdoSK
OpBxHSSm/5rFeiOpntlfb7KhRiyXM9AK6fyatmfNcbmVEmnGK4n3Zja5dRA8aawM
skjzdfYfh1GHxGKkSkdUfJrCEAzHCE1B+W9GpKL0Zd15nTt08kwq608SPVgHmq0m
I+QhFNee6jIG9ZjQKllmKXZVLfVLsCZSOC4AzXDuVELNn4Ad7CMuTwV3Gyxil/FB
uaH3umLpUrHCGXAKpJqvRWyNs6mb4DEFXSvLKJ7idOq61OY/17aaHMBYXLjmn5VJ
0hfpS/zqJf5Eoq0ksy+nqQCIDd2V9x/YblDJ2IOaFqPuUHrnOOu1xfVA99Qo0VI7
i2jSFqmfTdQTrCmjRkk83D31VdAt73wiYJp3uw5qoJY7yfPC29oNNkv+6GmtFCQF
AJf1rllWnDoupXcvuMuXH6Pj5NevAJJ6nG7eMm5/5ZmXJP5tPOgUBsn1UC99HK3o
F90aX7by6HxDfBq0yAYQJaXrFjYghQtwz5k831JD/1Y0IV9nHFoe/NR1lH8SlKfq
aDNmP1pC5I+ATh/8rT34/lvl7F9/LN2I1hIpRubqrayhscOybKam6eNMkGJK1Ts9
0LV2uElPiXTf+00NNCZUNZzN8W1tvNz7nxpsnBRNDJ2aomoxjiqwpLXHE/gfRIlm
NcGgdf1iARJiSszwToCStMP2OvxOmtUAnxyVmNO6TZwdbEBDleAsT+pnZrWi4Mjr
pFiNYbQQyA9S5rD9IWHIypidlnENalV+tYWQwhhjNZjmYX224aFZSgc+NmQje8ja
NbF9XsmR/4qt+/j6tOJUn0WN3Aj8fMct/7XUnxaaIYOyoQQzotTNlXTSX+Hzu8Xb
JiCrdcKR4ZJu7Xq13ocP3WoqDwLOXB3PF1nPtEqzNIcFp8IxqtrpE0yV0Ta6d4JS
Wx5yKhtg541/GF0zVxWLi7bibCsFM1/M8WJfFcQmpMqpFx0fWxhJzEbrdHu5pMHR
GIJ6fGpZeaYSXZoJnf6CnN4n9e7c1M+IAKklNXwwkzcoL2o4d2HJTx53/k5XKTXC
2qLP5Okccb2jJmQ1vss0UksKZ4cYQZlsJl1dBngAmm8vSmsN0EL633WcEJ7kRy37
4I0Q7FufjJhZyxzloFsT+ylOSXunHcfca2imwsG5NuHWjCDiVG7Fr+fl5YOEPzoh
SMlRbzDH9l2+bnWrU6zmyvk/P+WblEDxEI6MtW6QXD1KI4Au1Ku6aRLON4yPz2Wo
BvXVo+QBLFqG5Cz0Vl551tqEo6rwMnVwYuXDzDLqU0I4tl1mdM27uiLIVRYhYFpf
d33xnvpTel8u6637eSYhcOnUKSGIKlicDtSMQnVwIrhL813pXB0IrG8PMA1GkHcM
6Wffvfklf7QivxrixkLfLxR378/ow+3YQe15vA8Eqx9DDILoTaho7GQfE+uxCajU
ic9G8d6zeJ03Kwg3XXDlWXiT9pLJpT0RolrDHczK31jyu0X1gmqBA9QKeFf1/Eqj
UkgmvOlatgzh6QgnkVAruabR5Ib64iOGmiA8ZG5G/2R/P578lojbVwYwFZ0r7Ugq
Q8qQkibFcjKmzMNdF8FEjJhzejCEf3KI8M2o5lLA+QoP9D9YlhbowpvziEkbpkIU
voyQdTKwdoxuS2eoy2Sj7L9cnaE3wC0tQIXMKHOINu18Lrsq/B1wbPu6m7kr52IZ
vHjLgnQ0eduqU8SeBom1vYxW0/xo2APRI45/rR4s0qQRPmORW+bc9r8J5tNNS91s
zCFTx/IHWBpcp1AtkF9NiSQTgz1EqtFl8YRVprxJyuzF0a4ltv5tULssk/PRoswy
K+3hVndAS2Cl21/rz3ecKYj5eWDME5d8FwsgXB20/lkl8jrhWz6TCIFEDNp6Q5P0
eSfBG/qeiOzEBIb82Gyq9rc1KGk9JY7o1exRBklf1k63pGv02+v89oX078o/LQFU
QotqJWSZ5AfI+VWJW/E/jHUBdVCyvRko7XmQ96Gh4DYMLx8iTylJoUJBxERAH9MN
52jsYumdB90G2Nlq5EBI0NlQnUkfKrJ53nkm1v2oD7xQI870gGT2eyV9H3VYvJdg
o5bAKC+sEmBl7ceA+hSG079STzKkvFoNGGMiCmuvaxXV7k9/QDTLEG+gjEtS5auy
CbNJv7JTn9A7EV7Og07WgbxbGDwgr6QmFwhXIAbTyteTmMqlmBkRGNZNBwxyNYct
mtGEvIxMjgZq2xCpI+yA749Z3XXPCfGnJffMGQN3Cr+RkQmfneEDOcM+qeoeOCOw
gLPyII5sAjFuMl1uYtfj1y+Ce7D+wSm5mUmjKTkdsXW9F9xqkGVK2V7Ao33OjE0h
vjveCivr98yUnPhLMpvQHUSIIcnW2QIErSiDwVt/UYMM2503dVxg8epGJBTApgsv
iXrLUgydINyyqD2oWjB+ydtdnd5mai9xOLecIFWM5c8OFgJhtxdsyL2Y+u8Q2VC0
5IMScFjDkqq1xiV2W3PgGx43r6E6DKR5HLwVzcuO3RN7ur2z6OHF9+OSG2s7Q+IA
SNsmopetozYba1G9w/K7pWuvHO8FPRadRcHXmJWJpH/ltFgS5DhZqGO1OQ88gWq/
8EBRqxRQN94nfkw48Z6o2NFFVs3Cq6k2f5AAjgEJqF8snQ5ZjV2tkdO5kQuCaWLc
/LDmXTC+His6ce+xrZFdEDEiQYgNlAYMLeqQBtntfY8hy6Z2Wn9zFraeRcoiqKHl
78SO0GMa0Ylmm0NdQVh+7U3fkSEOqDh38FUGpyuMRQtA5ZI4jt5Rb/Ocz8/UfCPr
XC4AlqPkn4cGuwfldLjyYXxn4qrkZrrg0wg7QDHdio3ksqwF8nE47nWHLIGvc+zv
GQKDr3OeI794W5WTacMAxLlv5vj+q8A4rtx3fYh9t0QBUMlWbrQoofW6K+bwofGf
Zf7CND8FOh9lunETK496K+LgaMI8eomOKtfmDJ2GJHIdZni3Vlb6qzGcX0XpDPAi
mXEDJE+FIza8JGmyfmaYLnOOxSJyHb8q2Xvd/rITrGVv5sJlnx9kjM2VkDiteR7K
A5j9if7Oq92HeuWXA75z4VtrScFQcthG4o/EyxsCnt+bXOOt8VC9Av1Viisynpu5
KThY9lshe3r1lsF/Ln3W4Ce6c/FbvOnma8r7CC1NjdrJD1HupVneRMIvJiCB0JgQ
KT1EkRLFXjX8C5wRAIVM1c6AUwq7MKJ5mkVhWpeSZsQvdp8P2HYHu0rdFRsQSEQ6
/StpM21g6TQePECHBg6IxW+bXzqoNcR2nocE8plWLICG0voU9vihyHT/fm7wVUhl
2ad+RHPR3qk7j3/eR75aTsnjnD9JK858W3LJihSZW/uHBOVyW0Jch0nEI7FAqIwg
zupf6X0JxhicmOIa9rKb2tBdrPK4p3ELxB0eYaOnQjgM/K7cVtdrvRXg6MFFNlrf
TfrocfRtwjwHuroFGoUSPl9+Kv+XN4KOEYV7Bh0iCU/da1lyMARIw6+f7Ibc3OxK
Fskj954fB6lxb4t89TLbRnNsY4Ti00eFx+1Te9PAnPu9xxksIiU00a0HBy9rI0x8
Uogo+C5EE/Wq+AZWza/VNQc3KlJaNLYksunH9aijsGk0mT4siwTSd08Nt1MRgj++
5tKidIfuKyKWEa8BYo51OPfdwOszsEOEZ/jgmwoHWeijuIXxXmpZkynE2P27SyJ7
le5exB9g4/5O5QYBO8f395OhQm5e1mkqSm30AAeaL2ekShqjmPcURSebW0s4+k6o
hS6AobvF6EuTo0sjR/w181XWLcir2mNqjtkbyZZ708G/xhjDOHB/xMN4BnQLddRu
bxNGKjJPfjTxvQ29nl9xAUjv4tlKhkbFcIJ/E/a7Vku1eKauV1kNfpAcgt1j2MYy
ECi0h75KHMt3ecuLOhNHg+X66Oi15Xd+IMcKkMHd6sfqg6d6dtykcbz/ezL7rgph
DGbDsEGGguIXv1gSMWpsrnb62s0bcTZT43GqSzbdj6lsEFqwqH8a0xK+iuHnEGrC
FMUl/b+SYnfzQGe0OyiBGinf43T2/oTcEtRZ3sGvxyMwQQ10/8t9m698y8r8SJEs
QUAflYcqkyqGp53KtDWtGT7lb2H7wmXsS2P5R0rIRN7lDyk2QVgvhPS8QzDsBCga
tGSJvQhPKi/zgfmqihNG9ZjAQKl9hFHX+P1CVEURalsZwxPhxKUT0cTFTusKgrGs
D/5s6vE0VbuVuGtIW3brrL354gwGpRyxt0G1Z0Sd71ZIeZA9ovzsCsZRCzLsVLMI
bUKXr+q8tfVbz2o4hcLoQlIuBso4Rqnbo0i6KTTP3MqSWni9CjZLNo81SVOS2zSc
gSZuEXamz47gEeKHeBaflFJbqXn3q0W5F5iPrWrkPEgnSyy8aw0q2fm3Naj3TIgK
Ea9u9rpDEyKjN+B++qLMEZyK30LnvWNh4gB87vFw/eFIhYd+nCgPEfVznFXNpiO5
q6NQcUZbpgVbQfw03B2xgkY7KrJ0pLgBDN5aus2vwAvmSpnftwBELO6zVnaG3/rm
llp5NNOC1PVBme2e6FWI5Mx427MV3PNOoHhBw+LdmaP6oJ9MGOQ1/qVVeh1Uz+hj
4MMnZwim3Z7Vm4sT/TsktWBRV0MBL0RL7qeFXVLajJrryisEnRalX6D520IatC3f
hMAM0clBgCKRSaPvPDTGuD44jvswxJN9GsbBucPeFCDuAdx0lxYv22/gmGaH7axp
SKRo3fzJeNLT5clDo9B+C0kmrWGiiQy9dJaOYp7eXinMDnKxNjOjTBvacdKzHVyR
xE7YsAtlMGHMoGJJdw1HBuzU57EGZovJfTpULcPYnskRJrXomGsEznK9qQ6bQ6gA
h+64ivIFDAK50dqJXSR2+OTvSvDC2hVJ2nktJOLkLC7qDxQPKprtQq8Mw1QzdzFJ
if978DPdM/vt6T4YXY0OWVmOTugf+spvsrh4FfeKKE0UVOZX8vSvHekBiegH7cQv
KVUBwaIqh8AboZdL+G0pr8wtLrG9sQcXu4ulSELJY7fq8i3NpEEWL2xfIOcBk+1L
oCfmtqPMMRsrwhudc81jLfEcE4mN8b7foemwEBunisU/bwI9FWPiMgGNYIEderAi
BKWvsKZO8WO4+DWTsW35MbbtDU6cVPkrKq6IBx1pEvKhmugh/VtrCHXRnT9IbATX
GOpXV5fEV1mooBpfLtCuOU9Ebhag/xa3PDODabk3fi8imUm/9Qlcv9LUXd4Axk9q
VY1KCX85CfIrHkOTa7bqcD9Ug2G1sxwyq7FFGvkBgMDrtMHFcRFjgqCuIKeZdPrV
zYCZKZDsanqaNTuocdQ6vQO5rlz2vRpfjIXsZMnXq22C6CyrpreFguXMVoYRMmnR
tfahlJtd0ZEZzG9kmAru4HHEEgP0TwylRP/5gnWtpQJwa05FqSOKm/B3Vr5/6G1k
oddvNmQFO1+BXBmGtiqS7aQ/fwSbEWje2ka0jNOa/BRDuOkNI4KSQ4wlfglDKqLT
QlYmG3PRzip/RX+WBovDdxj1dmt8THQ0feJygkR2OrOfcXsIah8uy0vWFYaCw17m
1wP16JdhbZUjyU5twyUxJyjjhNLBO+2hyEnquFvfdp17npQGNHsO5n7eW07KKAeC
ubhOvstigILDGfcsfcCZTuCw8FU/QV0KhaEJZCnAknu4jT3Mvyh0RwcXAerysy+r
z5nxRZTbQwab6ba3uJ/e+hoDQAlIjbgzv7GdqRujCZ5/XO8pF5YmJN42UquT3ExJ
bUR8HdlhYulufe5Xgn/kzMM7WdG0ajKNmQGhgz4KTYwF2kbZC86S7T/Z9kjY1RAj
NvNeRcXyEX6nGRDkoFxhbeBFkot2dCjgv45fVpV5s7+yn1sJUPZa/ZyL8lf5Oa1D
oukxxZRLXucTnp7iu9qNUoxDh/4veFsIQs89fSetoaCV4LAcoDTuIlaGTRhry03P
u0rDow4RZCfLwNl5PRSGY5+JcqSkqNvhh48jk71bj9bttboz9zoxV3SpIV8MtQWc
yW7Ic5l3/GhDyJaEJuA/E3JiuhIZoKOfZ6GofiC7Uqo9L1DZh44f03Ed+Vwn4sfE
FexS5CqmJM6UXH6+fIjkJHyaYaZ04bccBUHxfNxIun0Wb3ge3OmJOf/3EOgxY/nA
DruoPQIOqbkcNFSWeYV9Zh+zNWJ/PPBXyYkizhPJyF8ommarn8KTDO9l4JHl/u79
KUqYWB4GYoKEKeJrunVHjrsf2S0xOx/5DvCNbhYPprOp/qzGl/71rClCCi5Olpdu
4HlG7kPcyHftJ52APSQxb4/JihRURp3Hpoak1GkB8MohaQtm7wp0lzAFNljz8DKq
mBwzvNAL4zhZR2OU+iIjZ514VaIddnnbU2WJM3gpcqQ5cCrmCyK1GGrNRp12Yku4
oGif7arcqf+c5PFi4o5NCCc7onNkUT5wNbzQk8NNGKq8PbHRXPwwC6BQDsJLGTpz
kD0r0Ly1u6qn8B9c3AaxYieD5EpAhoOmvFDt70VdcvFW4hYdnB5RoaoY46BlPOBB
QW/cFu3HhGA01mniSvW4tUYWwOdyI75bN80pGYG0qvalzH99GpQF2utV1/vFGW0V
jH+i3KvNiBvqTBi8HNVRESSEBZ23kxyvck5WNAmjEfxNfweXaVWiCy2a3WCAoDCE
6pkuQkm7SyuT/5WMYdPcOXwH/krB3eXZuslUoJl70k+eI/SWVkuMeblNGPXOzzTY
sZ+OEFixEnKt8UamkPYDL3TykjRKojmnM9FR+go9slm49mAG/FMJ+b+SqgtILDn8
swBMYfCEwNsXegCTmILDO4xdDQpr/yTs0nFj4DHPfZvVfGMMFA6CKntwJtD/vV8+
WCrN2dz0jNU6sxcqcWWdrcIezAdklTslsq7Y+Wv0gh29cuRVwcLq28FojMOYC+Jy
P3epbbg6WHy3Lpg5xKFkYwc9nhSy7ofmARVVSPNZV+HLoexcjqpRjhPJPCkdDzVJ
lfuLVu1PqXOgPWA/H1v6SY6oTgNkRTk+vmYeoi/6icJKYztleyijAmzQgf2sNl9p
Pga/A6ItLCgkmqeKhRoOUpVHImA6zk5vSSKizBbQqxmSuIlj5jB+4Inmxa7QaRie
7WahtViD8OFpL+2jS143gk2fJjYX+VC358n3mypGYfCEquHlv8a1ogjDcZAAG9OX
O6LdU+FXGoAur3CsKajvx81a6am0WZ4CmueMTQojakWchmRv455u/a5cL3JIOG4X
AKDYQhRDxjz4E18AnKNtg8H55k51repy04iK3aMeR/0mjPgM2QWj9MU4cgKVpuZY
AFhEb6pawY5sunfRTWcB5PpC1laqV5CKIx6xIkrZvng0nw6PSzFd84OBwv4NNhNU
qw1S6aSRcDd5fK/Mjg/z1LQh0aWEr7D4Ywi/IWFLSWQV6LHDDYp2ebEonS/VZCiJ
WZ+IecX0ftYsoOqhqpQ7Aa/TrKXCTkPCreB4pNHBRv30DIJYXvIM0RVVR1Q/Uw69
V/GXoqF4/WZtZgRqJrmp7TNOqIvJ+5fnEPCaT79/XHw3XErP2GNSe7r1KfurUo8L
uooW2CH+M+0XG5XMAXh1pMxPF6553qaRtF8C/UkHXWpeQy8TUAQQvfwuumhLjVF8
kwdEZXs+2P2DfDxV8PBPWcf19b2PG355wIwa6t+OZntmjYSUYLaJ9Ilns8e2Jib5
nffV+m0Z3OqB4rYgQVwlDiAc0kk//wHcUM+uoUtIPs2nstT9ArY2LYL3iOGZ1D4g
iEik3cN+NTc7X2tlmAX1DkTlC0JlHl7AhBb5zIVQ/G4wogHJWnYeCpqdWuhZJark
5H53grU1wg3N2+S8Ot0+kA1hGKpoFhtNDDSecxc94Cg6XVhwBFkaJM8L42R9LkzU
wvquyGYkoMwC5wZXz2gNGGmDezs3tYM6QCUW7uV52ms9a0eJjQ92UtUsULB4nYIN
lMyOOjBvTFun43pXAj3BXR9KfWwDzRo/bbep/12nk8ZGJ5L5GRD0ZFlBnyzlVuFK
JR49XyhMtRBuhRTr+fhVpeppLhfQUbYs61Q7QJ1bfW94wBkN6V5nbXclCG6MH4Ia
RdO1RwOP1yXbYi+UEZ3XLUmK2RDxouQGVajB4Q8pdQTFbyBXbRydgWLnliDEQGKX
WMAje+g8KXFGfFr+z8NbMQCHTVYfIS7vdc00WnzSimNCQBtbXjZcRUX8fiJcMw44
nqZVWaq3esQOi3DrZSB3wq4CEAZGcskWKUI+fr6GQasLLhORLXT520lvMsYQVsTD
RrO0Jn0jm2uoazYNlhqw7nbLzahAT3JYus6EmxuCgugK7PQX6ndzyKtoOqd4s+A4
98GvkXdF/CgVYwc9rPBOVvfgXCIJRokSC604J/JZXAhS/dqCeKvCER/IPIlAhqEE
DeVDWqA7vOIUEcZu9iuFyq33NwgQHOSflQSxFQ2nHSm/R3q3XG/W3OEdu/x3C41E
qox6Hcq6DkVgTBnH+uCC3HDRymbewlflfUSONgc3ptTBreM2F+4t9hSkhsng3NxB
uDR/zJ1jCdsXJ+QfwrZis0ZjpGN5lJXEk/EWl+13jhRVhnsHXhX4ZaemJaS+69hE
S1pO6wUoA58sVAsQlGR0idbE50AatZUXjO/4GsSeC4UT0ekB02I4ongy2kvztJt6
fQpvgEThA13GYEilD14gQ/CLWKmWbjksfZRYscrUCWUIw43xkk5929Tcurf5IpVm
CaB5eH7+0dCpeCaKhQRhzJQHXbUxQygaHzJ21g3QcOA/s8R+nNIbEsT0UbK+1Ahg
1/NNbXxGkMx4I50s7a5zqVyXDN6FovsN7n/o+lnrsMRAmXOYlbz9ef64F+CAHKeQ
Ts2/XZ25sMqnKYPULKCAc14czyzmq8t7TbV5zn9JOL8qkf6QRJen1F5I7TQkJe4T
BJ229cJDEAEjj6wsPDaAgMGqBqQiCDJ5S3guHI/HqL64pU9KQwREgV595TXGKitT
0ufAODzYkVQUw9H9ghKAlUgAhufHVHhXnrZuXnFGsIm+de/05UP/lAaSuJJ1Jy4W
0g5Fy4p1ONP1HLePxO9uqjYLqPAj8skU6YZ0kbEmwaKAI+lrpJEwM7c+1Rcij7wV
MrUv1W49Hg3gzpSid7vltk6BYYWbqXrTCyXroFJbzWcCXwn2npiScLRVmzYBvNwD
1guFQacB6jsTtJqL64hjeQUXfLw2OKhX0voO+kLHZvIbtzbPNPp1MK35TsKWtemK
FXGr0o9jARpUw/5cxNMtRkyqKv7xjJ2SiUBKu4euCNrVoap6P0CSVf2LEWH8i/4L
LUosqSrZnMby+JkekQZviFcFuiPee2OZpL8t2R9v/FgQZI8ejLsZjuNXDe+lMozE
bQ1BT9nkbIoZ0Z+MO/bwSDBxA6w7b1CSs0l2gYO9WecQmkVtkDgLz0Q6ka5mmNSX
Ce8T2BrxK71nY5myjsDklZ07F6ABySlzqbSSFgpGuN86IOIvHK7BW+XcNUZYh+EI
E7Xi9JbMXJl5n6MAKUVsZVVIA3jRw+kpyx6w7D/3Bksg4YPIzTSJVQGsdTHVj9Nf
9fY1GwMkv5o66wm2XJc31qLOIlvddRIn2QuY98V9A3mFXgMtVYtt8d3kZ/m1MkTc
ZeR+ArdgkRtZ1ZP/QqsgRzxdi7Ro8lmtVijT67oJLq+Ejhn4TiPG1161jdwJF44T
63x39cDMBL8UvGYKrH2g9kiLyjyL7BgM5GCETTxNzVGFeVJvHi3U670SKIAsYlfU
kWnZbXB9s0t0hF9bvnMiREZ8O3Vb9Vi/zC+fDb1cPeno3z6KRv2dnSYKOXZpQvle
XCD9QmqQueg6Jh+tcyvV5ioJB2YOaAI4fiXD6C5EpmwSI96HLHfMATKuUJbPiwhm
JUr1W8x8moy/VPrgAcG2jQhuDNCPdQLih2mxqqpfCg8VOXlB3+R7FYt+pO7fMdi9
FZEZonKy238NRsCsY95WAThAgW7q9IGtWU7W0I+7Df4+fwU72ynoA1SE0rTDfya6
mzqmVu4xcYUQC+g9f2UkD/dHnEgYsoB8i1B7sc7jfHBPNk04MRnHvfv30kJQWE3L
HVsvN17/1CvRcB/4VysuPYBuIRmZuFTSaxc6OU5Ke9mfsWSOYaSoMuhfBxz8Eenx
98z+3rK95rajc1RE0EY0t4KJmw3BxKgv6W/1+dZbZkmCUyQogd0dJH4xetCpchug
QmnjJGvY7gokiNi8zQQjYkTYAOH+BTKHTHoQxAPd4qnXnMa7VSbxSMaDgUX/fyKt
SZVWXhZ3AEFOurYfeqfzbghgrKOPft5qRF34AixRmVhsERuHsmC/cOj81llLfnss
K1yx2F/p5NREO/S12P7Q+AxEo4IKMSUSvbhKhRMi61vaMKaDaCDX8RCj/dhSZbkD
jK09oeduP4QmWaY5nFC8V1rzbn9AjxdYIH5uwkwvMrE0SGbaXsxDVFl3XXhOitTn
ujpUxZLwJs0oMfTIktAYz4RvGb/QLVvUnNRpfaqqAMSVM1KPYem51YrCW0WgZmpp
8I7L5+JZytr3Cbs/719X+igo2y4toiLSZI82SDC9OJBX4FimcGNhnPZnYgyeV9xm
9ffsb/nZaT7YtmBS5P26/7TXsnDTlklENVPmLW7OaKvLY0x0bYegAm4jUVuuxRMb
p/BK/agJ++nJxJVJIOrIt/uXlxsLgXx/EVrOzoVwpvDB2igKJFCpfEyLVy49AnQu
gg2TOp0yxGNGmTRyh5NkDm/HK4CxzWaEMaEzanjOidEZiVOkC/vHPj8v2gM954QD
Ag3c0B9Z3uvGx1HAzg2pVL1GeUGIsQpd8g1VZyvcb6JWTFwarcbKQUMYzAfhfN5h
1SE0fhUl3JGfcdI9emIAG9FyZ/cRZwNV3VUioLMjkUYQnpUU8e7lPORbfNB5UxC8
27Ce9lkIhdPVK82Mj1mEqGk2Wj8lZXd1Gx3Mmaz1OtC2eQyKn9zg30efkIxGOBdh
7GU8Kra1jnChG0pouf7Kwrb7RRJnm+QmbCHgbhIeZjDTy+X52sucVkNFdMBJY+wG
XH6CtCtf8t1cTWrS/wng/8oNcrmYtM6HP09QJ4VoyUZb6bCCkLHCBqUtt8H8etkG
58Xx4uHpOyxk0BVKirhGfw6OSFl49xPQJOioAMe8oD3RYXC/k8aHEPXTcduRMiM7
VeGNGkWNipHNX4un0C/nAiwdQiUd5KZmIBa8+ln6dvBydwZIAVY08JJqC5yLEn2e
R7MtUV3E5wopl9rDIQlOTmMrT0yw9iw6H+rjixcEojbeh/7svtmSbadUby8nCQYB
6Exp+S1CBYR9+ps5hMc9WVJ3p0t71fpjqL5ibfjuWZj3N3XRnJ/9kBjk1Q1C3URm
MzmF9AErqVJaDwGyTluMaDClaVQaT1HU5wNCSOZsELroMqYmv2TqtV5RlzDQKC7c
Npf7TVzUvJ6zIvB7SW6guJRVcu0JEiartbAnJbox4wTBl0DO/NBe+4ocGXdTrbEu
j93KCw0i8dwr7b15s5XDHPUfOw8bpS9dPMXK1h3wdvYC31qrIqWFG90H+41rOgtA
LE1+PzasVPT1AaDEbGAOept7Eo5XIMfvRH4wdGBixGfT83M1DpWV9RMeCE+nwxjA
w38DWUUVQqwIlR1bB5RG2oPMSKzs5jXtn0X5CJLv8ixRi0EAVcbUkJbW+p3bJWvF
2ioT8S8Uyw+J9pVF2RwxYdZ6o/6KA0VDoW/dGWnd/P9+B1K9894zrdZlnYZhvdTz
TEFn7mUsLGaqYnG/MJR8D3pD41HE8fnGRwlAiplkarTS39q/+wZEYNqjyZavbB8m
l6UD5ft9UiPXGsto3il8DY0QZMuPBWioDsjaXPQH9H5XPOi9xYaVYH+FzMrTjzDf
MfXQ90jU4Uz4QoUljbvqlwv0caprM24cf9J0BsU9JKgU/MUaD7sNC1gvIOZiC/Zm
qlUc5mreSAJeh4wA+sGvkICf21xNbXJbim6Cfd9oWpSzG/gJMF+bkv6/hYj6NRTD
bshRXbQUeC8tlUXqrWT58podoTG4h2GE6ZQBaArKsUN1QF/m8XKpuJGh2fXpCBDN
NCw+btI0UAw1SdxSaYOiMBIkEzDFG/WMFZwmkU3KKMiY9t21W1J7hNprL/Pu+eMt
VFTyzGpNGBbMrm++q6KyiYdGbcxu+JAt9/241fGhkP0nWxXTsKkWi77dhC1yhLuB
GdnunUQGpYdM43Ao1NWzcFbMkkYsCoYUhkC86EKnLHqyv/3AfRaGoJLRa9y8pL4D
l7d7tb0XaZ+LOjQpwSLQSN/RUeGGrEeeNBaB3UVJ6fqe1ywHVQsejUaGO9rRkQTY
J4iy/YGM+AeroLUDN8VyVb8lrUH5iRCIj8uz7DiZ2dnHAXDM9/iiWE99wLaJlIb9
`protect end_protected