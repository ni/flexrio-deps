`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
oDqealYugrOC+OIsTtIIFBa3FpZNdTPDcZPFr9k4k90DxkwM0YyGY9+lLCoUE62a
4aLTri8PN/6c3ewf8yrEy+VDys0aELXCE5RvD+i3ruFtL6xvGKiubKtcycRnTP9n
vBaNBFwYCDsF7FZdWMYcLDJa8I6yA/8DtZFgpfbTLxwo6ekPSpjZNcdqTpGUt7IU
W3dcxPQylxSw+RgqH/zVQjlQkcJ0W7tMh+4hT1JXQOw6hfrSQDiN5mddv1BdEY26
o9kPdC/4/+V+7treDOuVvL1Rmbz7LOFu/PTIKahAouIowmKMtG30LxC3NXUggVu6
C0HK2Lf1UsmPoKzn2lfI2Zzin0qE6wjFPbdSqf6hNg0fsDG9l6mBk6Sdz7bTMlvl
nWfp9dR70XdAdn16zYBbb8o6Dh+EwW8BZT/ib6YAtcwMSBMUvyIq3o2V57pKT1Vg
kAeMuCF8ToNbZVgdBr0kO5k/5lotcQtOhOLRkdVPd86YiD8JHWt5eAdJYmr94Iom
tprVawHclHo/7IvcAwjGMbJTCYtMbuw4i3cmI8MkhkAWz9XReVgGyqiCFrAEE8bG
BjHw6Nfd+FBzeEMZthjMqNi9pbKnAHsBbz+wAZrQG11xIKkHZovR+5RODrmYajAt
UOFY6zt7/RkakESU5aDGtpcXk4vYlJYNZDqrEs6/hU1vGeyc3KgnjntXmo2+QJHd
nSfm5jvP3xWEAu/9bf8YEdYHsMh98SJwxJmr4uyop8+mgg7gH9Dv5ZHzcYUlnUW9
OF0LLXNOh9/KWJ0ritGv6SslfPttUHoa5elHylZx+3WtgkEUNP1lO7PnDTQI5km/
4UV9hLzyTsLrXK2XdUetBtT0waZ8bWRJXLvNWNdrKg4dY9C1VCQr/ftnEczG3iKH
5WGj3XjpAhwLNWphl3RE7KllWNiI8+Jdh36ml9jtlX8h6gnT8IAJ5sehh3iQU8fw
jhEooRV716yPuzxGXNqv0WrHTAvynfwgUyggCk7j8YCyn7oJwl6eMBu4Iv+ZUO22
/P1g8qQwLT67M9MM4ZsqcmKGBzZv/t/Zi6Z08OzUjSfAuqUnPhHVSr3DD48X+pvw
FfwTA6SCvfiWTIvzxRcW4TwPcYKSFfSMNBw7IWkcXeQSn9KMgYUmnDcc4yJWu/sT
31Fz1fq6EvQZsnHtVhWjZI3xqx2qzihy4W/2Qz2Q/RCGlhBCVIEcv1aqTcNCBimI
OrPm1aEZidx0+Sqz/KICLuLH30YuUXwzdPXcLgjklidWTAfvuNjmLup1v4p8VEWu
3ehgpkiaZCrkq2w0VuH21ZdOSXkWjtlZowgsiq9Bh+pPFF2++V3eAH8scN6vNATA
o3k7wBxWSO+oUOF9snjGiBhu04Hcor1kLSKvHBpxCuiLBpXWlFhxAlyol8AiQy+G
8t1cMJ1Ou21r6gYAceThRyEMJvPNVKphUNKulvdmKu+/cWzTIVkmygKmF/hEWzAD
Q7l2tQQN4gdHGo0+OmTPSzdeJs0ifN0UToOWfx8OoNnjMxz0Cf/KUX9n3fq6KdJf
7T/LMLWpEM0vWEBhECrnp25cKcUkhcfDP+Gi6xtZOIA9YIR+bn6ijLdwNuCKgxJe
yUb9DzG/FejlrBY3CaGOdwycXcG7RaP3xlM0AAhlxW680gymicUxaqaG3HczXz/9
PCVxwxmXRrWBQa5CS84rUFWhJ/RxI7X9Bgc29oEGMi1GbnoIq7xLVkV2GbWO7F8v
LRdHW4AAABRDDYzO4AONhxTMcg6U7nzztVh9PDx0zqt7JvqvscbW+cHUV3ob5tdN
r4zQA5psidMuCi1WLvtvujh5J0lNWXDT1ntbftuOcHHkDT6/0W7AlbJzIUtuYwsF
TynY+jXMKll6H3U2FkRMch1s1rTAmDXnDgO+hEkGNtXuQnkMByVBbvMm1SnEJlEd
lRlH3fEf0MSlYb+2VlPw+yVMO7pO5oH9jHINFgXilp1TMR/DMoG0rdL4Y1ZjcjL4
ertgBLdw0Ia7PmN2LlKJhcaNaQDyk2UACOY/aHWqI3p3i4JuRb78u3g7/2Y4u7AH
bTS2AnNRC3Aa0XQ7BwlQF7n9+4RIOv8F2XqmLi4nAHpnpkizczgyve6z8A8mGPvP
qycEDqdaC6A0w1/0YyT80VbnYrOZRNO44LFW2uWJ2TbW5/630JHQAbqt+92eqD1f
XXLe+mK+JNQQtusSGFJ0j866FwU9u04KPkUkeYjLBu1+uqUjGk8knbuAjMdB97Xr
9nlV4nT1yrVEtD1QPndOwqtXR+EMP+mLDWbaESNkEI4qlBpkmWn7mIeXCNOedlrk
oS6nuPvbjWDU3W4GabX+yhe0ouoH2oNhGv/K2hNQF3zQZRSmOjvRO7c5411FokB1
Z4ULXguv16g5BQRohOPdqyhFPCeT4DIfIY8WrAf148qmxqot7V1tLFkpozY/oBj9
OuymfBzYQB2Gxbpz6QoSL4ICuQ4NrzGEXyfMiTOyuUssiYbX+p/NgL0VTJ6LNTDr
qu+Mb+EdrVKh6VnFobAKScbeeobLnKYDsk4lzcz5nhl4Pd2OsCQxrRMo/AZ32sk2
`protect end_protected