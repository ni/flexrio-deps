`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
L2bRNdr1lLBT0eERw3vGlGkoZyuoLDUOvCJ2jqvihXpX+RBhV2lPuZk6ALHQ/ugO
hwzbok8EP4PfZc+0VtMrKzMMwEEp8DVGMXKFPGPbNdOnZuFLwc61FXOyUq/pOgqy
bVfhOHjiEgSvBjLfcU6uOaqrq+m+svFkitDToaQ0gdM/7Wzt169sCvbAhsauROsk
3GlJZdFT7A6aQoWO87AMWBF/9QMR5gReie3N9Nm1esCwCnCjsZ1k2zfsaqvqqNGH
9BbFfOC2nUnySO0CTlqz/U+LDx7FJCq1fg3fhKPX/Dcdqfsa/jdKV0NS5tkB1tJk
vULQPFIbEA0Lsb4Ti9lLgJw7QQBuV3NuUqwBvIJSlAEeHnpQenDfEmNT8ABwLbJL
DmPykzxj9w+FVAf924w0HyeXYv/cGBFbk5vm3BI03exisT+1ETNXH1Zf04f7tqZS
aZmk1Qu1nq4CBhHC48hZl8xKz4Jrgtz3YQwMqf2z5/gSqlnQUhJsv+8hS1aY5chy
Swks5jmT0Abj775N1cbU8/IfFKUuonRcEL79+79Ge05unKK7BhOQ5Vx9hKmnw4a0
VGgOo9FTLMkMiSElDpgKyhvCUoHdz2l0d7GbMLrjXtqef4qjmcZUi2EitrRNC9Qb
SdTgXw5rBIt3gt0wByMd0a2mo7fxU+Ifk6062S1LmWFLp8HjjvnJS4rzTECkMRYL
M/xsoRljYcN7VCJhUksDhEhzYIt3MefzPRL02yHATqX93vGzCNfN/GdyYeV6/Qdh
OJk0rzCxJhmesakdWiFKQO2zo4TJdgP1yO5vtCI//MNs9yf6+nNqbS1qV5noMRfp
Izm9bKLZzmxH+esqzdGhAcVy5NehBYrw6Wh1Ck/shoHAvLm/9BFAlBPUyi6WOr4T
vyURgUarRHTUYrmbX5mJ+oL5J7I6+6j73ShwXk0hZ0Ripy72P6Bla4oE0RcpeoLu
Ev0UcMDg4Sezo5s579f3ixzscGb9hxH+ne0iONxJAntDfp1BBO+CX8l31b7igOJa
K9D+uGbWqsa8/r9eyvfH4JwonO/wh5P69K+WZ3JiXaD1+GajS3BGPFnTMZ4NL40E
DcdWH56xiF0WUVxn0vF55Jy/cuPhp6aiZx8172JkpyKTkOii2h5jJbQ4f4/b45Y7
XbPiyrnusfNgTsukXNgGnaP9N1TBAR/6CqFDbsA8y6a5vhAaWAS/lkM/XXLA6weL
2gYbJOEHM3xD+Iza134s95McO+KTH3BYNA3nPDHL8poS0TfuspwgRV5KCY80fd7i
46L7bRx0XHGMbKx7z4BoKug2zK26UfgN6IrLNNpPHojKFSAadX3SKFy0JfGGJCHS
hP2Lgdx2l55TuUOIlA64Ve6O/p0zOAbtq5ddg9IFFxmmruNliW+ZFyGvSG0xr5Ld
yWM4Kg9mVeEvbiyL145WGC9E7ZkbpMUzqkkpUXKINwWDhxvup/CIG4YJGyGFN+yl
fr+VI58GrhazQFAV9QJUx5KILo4KQo7s8hNHcWB2DAxaHfERLnpwWYFsAV2StQQc
u33jpshcDIWxTnsxdkAfOLMLN7L0Fo/fvna0gQD5lOTCb2mZh8/HiAt+HCaRCwBl
oNdPln+oi/nrMsYiQHXEHHSUnpiFhdta/kCU2/YLeynWWO8bOZJBoSqjbETEbaX9
F91s2UF5NV7r96KL20huN2ykD2R0Btf/zqarCmohFwQff0pniENRWd9aI2pu93rQ
jqZQ5udqs4ekM9hv9+ueeTSsuvdnwzpLCFaMARmIu6c0IMv6VewHxqARViuy+n8j
YEncjsANLCJeaKFU6KGi0pIjTTkFbhk/L/g4POSvhXaj6emlhcLYxsL28pkIj4TW
Iid0WD9TQHZLlcUwuvIsgyzkOjb9Y8DcGPyGNGE7kbpU5BaHBetBHxM+5l2OMhYo
uTdih7DK2CFFewcDy/ZbrwwbaiTA63TTPjsOyH69kA6zP5/Vxncgo5/H4GZjRtBT
g1vEH57IzfWwFw1b6oyxjsGGKLx4zJzRKKp4SSeUtV7kmFC9nXwfZQWSsdLI+GMt
RsRAwt8huOA/VRk4MmpHDkP87jqUMG2QfIcIJ84eRwUR+o5Kf48NnYEmBbOv8A6i
kNbacZ4wrWJIfyVVcMHZ75sHt4aaJoMVbp4Nza4OhZ8BTEBS/Q9FqkgSE3fuKMYa
9LvkEmshomXXPbdhbhMkB1rGA7vswD0awL0WAxXx1avQX5FOOJtKw8u9DI9bo/kk
0dOD3kdWtkoxtYLfhqZOa0WidOW2RexTNwq3aK+1YR+cRkj+s5t3LSd25tIg4Jxg
L672SJ20Jhp+IXaaVsboU9yNoZCV50bfL24084ZJR2Lb2lbKhVL/Sg8nV3CCPZ7M
DYePT61lDy/ZkxEa1GEnt3P8PcECkkTvOmhiOW+9j28iYQYsoB0lr8Ft3Lf16rDb
7Gcb3QYIHxp9twysIrC6VDMeuMucLUOP7DKWlaD5iMiOdb9YiMr3+Q9pNQ3dNzZG
9lGa700CT/V2F+chmDUHY5cA7a4bkfsIBKvIMlSCbUzqxRMDK82qPFlg7k7L9uG9
OGlagHwCJogRgS86hhrf2q0h8EzNxRlxS5ooOhH4oxKFonjqvJKb+8PQ84omBOoX
8/aTZFqlsdVcH+r6FB1B+m4y+3J5Nskqq8jt5PVhAQ+4RFIyYqoexB/yh5TpKJyt
4eJwx9Y1Ssi8fd9qA8nveuiQ5IqLY3T/3qKcQLLd5rqdM6X4VI6R3IM9z6NB0urX
MR9vyPuSGl46NQtIb8sqAMZG4EGHpfxMNkNn1PqMTZ19BRx8ArvW+CXH0lo3YjwK
LJBf8m8/RXDLl5yQf2nCXo2XVce3nypievuVguU35Ly5lXrAdqwzSJB7997YmYbT
ZWM+FEvg8NWmDT/uzcAquFGMOgSlqQKnp/MDNzGs4VZbxMpKV4N9q8ZVeBDe965S
UJjbjInAwMlW+pR8fYvQGmI8qhmnVvkAu5CasndOW+OD6ua0y629rzSsbNPFlw6b
UdY6ZilUTuYruVS+En10u3rjXUA6DXyk40XekWq0841WTotcxbVwKEumCzbDpUdq
OFEVWmE3piGD/7jxZT0yMyJz5YG7tvpsBmxXvXl/YtI8s8slSKFYQ3iuaHhxVISh
aeOKXYc9XH6/6mTvUDRaCICA1zIxgViFhZAySdo/n8jTJB8uied9951z1BPBQEjq
nY8Rt9G6GxaokAK+nD6Ie1WKZHGTECa3KmEjdvZeQiWBCJn+H0tC3HrHoDz4quzg
h7iTjq55wRYyHsvFc1WihjfRPUrCco+NAcu09Wc2ky1EwMcC+dlvJ9GLs51h7AYu
qqugQPsiNN8gboF8x7bFUbDLPdtPFwJrjhv2/GPJlbGZZ8Mun/bz8jf5++127A2E
mftmQCgSAU0nQdumhduR5P3ts1YIbusj4aOK0BJ0WQu3kZsZEYYeOsCPonreklFp
ZdR3SeF0RN4PLKHRIvO4/XKzjv38BgbMa4STGeYX7DcSED2o+xjbkFnypz9YuWXM
cPRCeBd+U9HAQYV9kFFC0vEQqsHoVJHj4GfcY62VuMxZB9bW9cuKTDR//aW686ZK
7KWv+DpXqXgp4ZDzbTUPFdDctHuFOsVw7PSHFsMYVKOJivFbRTZRVBW3BI3SlIv6
FUz37bh3zjcMDVasj9zGGmZyvIi2LGuQfJdnUgOQdM1/sDnx/78jGowjpi0oJAS3
2zGRbKimr5dJOlykQihtYJ2USGSj61agjaqGDd93XKnADOWphga1sv/f0nfIg3GJ
RS6x/4LbzB8KA8sI1IuCM5EResKTMkA6BRIkCsYosUQQ7oMKYyjvFBikGfEHQfEK
91fQRFQJ5VcBaggUusltVNiiCr5QpCIZgPtIiXqAiHgDH1XLNxWuGjvNmeD1F9WU
WBaYUPBTLYMkKWOyeYqRkQOtYEHYPRCjl0paq2gmhszqNboAYzkhfv3Vei6Qr3fA
joL7T3xmqpQpZCPFWbs+nie/RqXphhjY9bldAM4GjLtCprfUQJGdB3vIdSXfahn5
73EVrNTVLFHqbxXrqWwbfJri1SgVeAlNX/FzWJj1/11v19QeY/yJDoCkbQdLM7NA
th4I96p+SG7b78Gx3VzaPIN3RxJQhnOO8uoSJhHNy6XuErRfpNaeojTJICRD+GKQ
su6dMJ2z+gGE/goZrT4yHiXWB+XZPfRnd+VdXvckXQpx6cAwuU4ddJMVJG8xizTl
LOJ2DO4tFdfCDBvbpqVtPg7wtvVaj/ABGAk42M68XnsKqv8M1y1X33DwMaARkPUs
Mu4NN5dgt34/ZHOGR+/xDCk0t2dZZ2OjWRuj1htt/0ULuE6gnaB70nxXTJsWZdIg
3skexzsAZCrhPJmBTsMYweVcrxFae7dx8VawlykaEAof66rv6L6SdMCnLcDe1wun
TST4n/2glAhn/orH3FtEMIMsJkh2HGLVgHZsvH2Varls0ak5kUczvwIcmaUfDlAM
Xj3d905e59UOw+RTR3ePCB9QoMd2kAzowMVrK80Kb/e3knBUV+RT94xdeKPD1L53
bDggiB9IJemuiGidMJrlT5HjvfDu1C/80Mdrj2P5tAR3kYU5y6QZgcyBYkEZ7uTv
avz0jFyWKVtGyYNQdIEkDqHBmW8Crv/kIl9jR3oo4CIdK2hVYftA3wpJQnwEIwkZ
h7ONuG0A2XxVqcDBRdbrJ1ovBEYCRyGlc9HaU7vnP5PcVkz0YCiibSh5ywuoHrwm
cMqNzw25Zez0b2fqQ65b0MmYEz93xgP729JP2iVEMcP9qS12CuLLS4HSUEX6T2Zk
Y5l4FYNKKV8YTwm4jChy7KCbn6hP+sHrJ0vZ/tdZRXJYt3ro5ViP13BLwm6kktOD
Qv3XcFtdevoO37SgEBpd+SGD6KV+86N0ZAJG3jsx2bP3ZOtNwR9DR5TerOzaOzIo
0Fuz/MoVk9dSJxqlu2nUGlVe8ievYYMFe0kSqDpvbNf8D6eKDXfygX4NqhM/CDZa
ahcOSdiILcbhuP7Itz4n2kMvNGhQoXe/DFZ0Tz6J0vGo8nutI0a0KN2Bbpv9vgpg
UVwT3cZiDNXDzWDUyh10Zw8nXOYzF/TLMTBR+9PSsAWkWWHMwEVrHvQl9SAldsxK
k8JwPp5tVOFEYBvQgEuxKkzeP0DfBwjE6baeQX2s7vU8u8R1L8sqNMG+gsUD6bvs
adMQ//404kO4tyGo51+drzR/DF2Sd1S1YIxf6U3RJK5ClkGjKVFXdWNZ0Y5Vj7gC
uSvk5pt4VgT10NV37uub0UKZu4oaF/IMWTST2QB6bd+Ngbxkrh0y+KIZ3tqumPmV
cwzMKvNUlv6jAAM5YgOVOeuXcBagPt+ynGUOsHJ5J4S9Yxk1QcKfczJMoKHIMvP3
VU1GFdIshNMbcJVopeNH1F5Kg4xOFtFr103m3bB8dNMQ1F18JFqGbfNuiXQIfvjB
3Sx4VFkWWATQARv4Zxr2rmwGLP5yckXbKNcxeBfMtPaG7Uqt7ny/A1kCm9zmiF+i
wfdDSLziD7508AozAuxj88rnLxD+mf81jGLsYg3TJRm8buMSDLCCYylhxtIhnf9Q
gDgpS7CzV7WxzsmioqdMnstfKqMbyesJO8nmMgFlYpRf1ZI5ENttQMR0CaGJrFy7
8WjX8gDl4fmK1bcrQc4w6DclEkp9X3g8Bz3COOZFQ8u04+Kv15zUujUR2C/Yh1UM
XXqFJGB8z82hZvec4JjeifzpgDIruiIGAllpi8j1l/qS691oonhjvt95pxX5lwhD
pGvtT8Qn0z71cAzasAghWWfUx7M56qC4JcZISY4Odb98i1L2+/nBv8+7mT34ZGyX
Ke7+u1gND9Sou1wuY1RluF8LAUlrzIz2uwSlGIieAHHfP1E1PFMzcPuB2VSnnnDC
LHOfx3txL98C8IpMXaYubL1XwNUL9rdOjmQGxV2HigfmahYFJWLbo8IoDaWOM+70
z7tcnG4F7NX5w5AED1XcopDv7UHWzIJ0CkTh8+lGUdYrkU9MwzjdjU02WMPtJr2s
pdtPUMLlZxqiFG0vW6IyzMxmshL6zPt+KxUOw/eEVwMG1NNEMQosRewKp4s1ld8d
lqjXgDoL1Zy2j7SlJgUScDlrCndpeG5hdX5pu+8UjoubUp537tthngy56576tTlp
iGia8fBrHja07pJoiqxSrOhc1Pvub9wY9xughLsqF9YFOjtVq6Kn2DTvLo0TtLa5
+F6ZtDSrA9oLOtLYUKlkwlaHBXpySCNHD95G1rbyqjBDRF+z94JhqPFp8pfcBKJo
wwdGrI7SDLUDK3iXnuhV/6ig2g0GWr62xRWpODF0vNj0HssVIyX7eozEg5QQC3AY
+X2xbao3miPImWEBw91G8sJWL98zF+OgbVHat+uLO7fQGf0TeqoHRlyphoIeOjPz
0z34IIsgnhAkkyEjabAoI7fcJwbdzY2Ew91CCS973FHcCe6xXSF1xnKG1RJZP5UC
vw+6+8x1SAdE6UlHw/qZo4GsgvJEBmsHepoU1b7nxlzhyfjrMPa91IPGEBoh06bI
W7HAQyr4M4tThHkKNGkxo2cLBW7dJUDoc3EVvJibOHhpBrzTqS0Xe/7ETlR4Ficx
QiVYjbaivfXAJNfRQIofDO5EdTTkk0T0xo63i4RWy8n0wOQXFQDpQohhZ1hs6mhr
WxSURJLqE6eUnPeNrZDFaF3/a366dMum+gVsicyOxbdeDJeg62NxWwKaXDx39MFB
BLjKSzmMRoYrBL+QAjdFscCBZ7QjzGFyK77jFbpMFQmeYxN5xT9joKmZEaFVSpE5
ECQqz1m/vhKcdS+mWVLnw96SEkcLsYZMcClhtBtp63Rll6EvlrL4Oxh7KKo/oblx
2cSs0wTQBfHgeoKgfZVaMJBDe3+yClhGCH+8bIAF+d1U2VZCSTJG8YkFh3vwPo7c
dDkjQef/yaxFZhXkXsSjVNgahZFWe4RyzJuDlIkAA/oAnHUEwm+JStxNW4stZMmY
ska0MKY3LD89kkwwXUUE5pYgH9lYfacHtdkrbeufQdkM/IoDyP3aOYEF6hGE8tns
YBRKk4PQmBgJ0qpnebw+BvsMwtkld/+loW5NJyLCOlozMIjxjhDc39AnGZByUedm
P9Syale176k65E7bIFd4LpNiA17tClWOp2x8piI3nAyVHltrsV2TjdQquSuyIvS2
1+CUfTk540BNwux0EbhQSoRE3jvZ2GXMjNEueAukqMUEatKfOnSEfFvMSi95ZARZ
mm+ofY5s0IQnr7AziB1bOVWyZmfibvcY91JBvK93V2RSB9AaTVDMgifGdeI7Uewj
NXNtkewg5AgSZCeSyF4xqsCSZhwbi/ezNOpsK0+Wri8zuSwqG/zYamidyDqRetEs
PV0H6vAQpME/nv95N7D0+Ih/1wkfCHUbBSUD+MjTVZ9T5hM4ETXMwx+a1rUHh6xN
/E5iWRgqpqsQmFligiBNoqddpuJQfyxrp/uWswT3fjvtGr62P9VJ7al/5hDQfhZ6
P/DfHGs3GUY2q8W0NlCPn+66vBZh/0Zg0mhn7G+qd0uymxBPb4Q80d13LPPAIvc9
pqF6I3nT+VRKhdIMp0z09TG24Y8Olj3mgGSA2Yx+wuWe5/TqXXGhLVf8QrZuCIom
KWeYV1XEIdMUssCSeQg9FYLEiTCm2oWRlTnxbPoKtBeoJAbazFGGdlSVPmZY2f5p
4V/TgS3YjWy9T1OblaUpa5fQWx9z4zOus2uv3N2MN7SZzmrS15rwyEpfWg8Vn6Rs
pg/Pyv/ClElUeoifRRUPBSu6+6BcMescEEDW/A6FouLYy8ALGJT1ZubMBA+AsIkT
HdpcA4UHjL6MfTtzmA9kTJRWO91OBQPKOX/hMt0mRxfZFzyBaKUw2mUk2C3bYcj4
Oa6PdMB6dAVfjpieh97H+c/pzu7YhhB62wcH4tok4YAT/CgyjYCQUIRwJmeP44sp
nicnSQU029zNCCq8LSCKRHDagH/9H08lblzrS0eBFncp5Wq8aGqBpLleHHuEP+aw
M/26krGkbjYpb2EaXz7n6/Nu+pQPSux2Pw/egO4k/7flSDMPao5OfLx/kQGgCxQZ
B/jysOGOuzwHt3cOpgrl5y9T22iy2WBzX9zzSk47sJE8tI1ue7LhZ/wPLdaELuzO
R3pdg+7Uvy17uFucve8QAHnBQiAhmRI/WHGNtgNuX8kGh0PeIxz/0BoR4/7fauXF
iDdUwlHxbcEQr3/t/3yl3/CShMVHGiR2eFjU/FsThwNpt3yiCpINqrg0kM+ciZS4
YIycaXZGsxzwoGVLgRnhmTKBRZ+cpfflX8MA6Qf/lmGqhu3GtftO4ThcVxhvFI+z
OBbIlLk3p1H8oShbpsZVpozkvmpJJlCvYa89i6Al7le4e764OyEyYe6CbQiexU7L
MpG95GImItwo+NO4Hzu/uSr8MfQg4QTHBA5l173AnZ29uffeBJFI3fTl8ojIcSbp
GvW7Y6XaBPa9h6RynqehhEtdmg1Ijmr7/ikLDAgya72N+xjiGBWnO/rp6swaDQMo
LXOsOiOkmOKbv6iXV1rmzEgqFgx1DLL5QitRBhcgynfQwRnry0hdtq9IGklDW/1N
yIXU4wFGrMLYhQu8TEqsL42s7F4/5t1a5FuzME/ogG23UOfHcwNUTZEFEbnRMiB1
MS4ZOMlz89icK4cfI7j63cQ6xBrpfG9LLJflWIwXzAMMmOdGFk30+YYyJMgSU5eS
l/GrSQdPZL22zWsI5aGGPnxiXLM0Y8E3Bo9LTo5mF+uaH+R4vV2cwihxGYrf5gIo
WUU902KUEiXT0atfdc/RtOqr5wuX35PB+eyfkul97egYAUXm9Gip1dMEuyrQDSsq
YVAqzETGeVPFHKW+5hUfOLTWZB7QmRjzlZ3ouoEg8QdgHx8jmIQhX+E2TKGUmlxv
aDatI49asK1h4Fouze2Ikzmptc7UAwC2rwf8VHDdi2QA8SSwWFY8qRvB3VundU2G
jVMkMfRTMjo8TgmLGsnHHKAvJ3bKFE6ZiA4Eeqqeyt3JMLjRZmWGquApZbODiPv6
pT4HHJ2Q/bE7nVC53giplwAnGDBODkDvTmtOOv5jZFQH7RvttCmx8UYzsIGxp6pj
oEhXV+7RWLiDAzRpnI8IUjrYNdkEJHlxarBcB4U+h8QQ93jsAmTvSJIOL/W9JDZV
l4LddeuQhfMmXck2D3b7g4Lyt14WL7z9GVybeXhy88mzJvyr4MNicMAGcktm/U0f
cCges1ei0gAIFAVT2E25PTaicpmoxjdV0OGEBOgAUkCKigJIPJO1qdGAoH4P6hKm
DLt3iUJtST5H1iN7mIBXzjKkCtJ+oCncbYbLV6JyKj3baV0tCeORZkAmZaNpQZ2p
pbWq5nVlpbSa3Vp9lsFetEm55/3irmMFoogKpoHcJXjuVrUTNPoNCwDr0ye9jiXF
SKjvL5+fsy/BHEhyJ52D3Ne8HonaFstYQxQHbCxMPITR1HY2Z3CuPQ0CnnxXc3Q2
kFEQIDwLUQOSRPancPRjX8wWgRkoJj3uf4XPfkw0YYGgTuDxAX2ldjRv7LbvWMqv
3EpBQlU1UizMO5co6tYpVfbqQ2k0IsWeRfKHEZlDDNztd8mYjJNRc+6n/Hxm2rUq
r1Ti8W2fMNtWWVtA/uuuKaXuyZsZXhJt/vh3XPoJrYtbshy729kvpho35OJhaMou
XXROeuHmWwTFgOGcrVSh33OX9QUTTFA2bCHx6yHoq7f5bKO9RBx1SuU0+UDjnhhN
19KX91CyNePgw5V0VPVVWV/y4kXTvoYjjl31afdZ83VIKaHseqMvs0Ayu9AT6LSE
m3Oih9Epl/c6s0QJfnVQS0jQbco64ntCuSRPHBetMVaCJ2q04JqHz+mdmFXnkLu3
ujDZEDWOcQrmpLDiOLK1FKkOx6r8O1b6VnWFIBZnzlDFbKJGuSVnc7F4BLPhFByx
Nhk4wDBEp6H9y/pdqbj3DLT/8hgcL4q13vNFiX4kUwfD+fJ1MA1BMpH/YzD037U+
mSEtmf0T3CFgo64kp9ofWsYbE5PY54xonagxGlzXFf3nz46n0BMe1S1higab5t0/
Xy2CzsmFL4OXDldm9+8Xnqecsl7iWEJqOYtUiTiNDtlzgEP4Cxx7Gp2YPbkjMNYf
Z8IlwqSsGU3zrwARuYMbG0eW32+vZHwQiPxYihLIe812JJ27cJbUFdXmAFvrWNue
u/HzuI3v33C/VL8IGpnQLicOjnMxk57BTedq4YCadiZ+A2ySWpCQoGH2FBGRXPQv
b0HblKEcFiPp3nYaQV95b+vAgp9e21sJiWUWVfKnqQXQJffsM556qQES6wno9yhP
ItWIFTahu7/IU+LVORuenmV9Pd6HS3zPaizG3yz9OPSR+w3sQsB74yz8KrVKoZe7
rfgYQ3ChjJcyW2SXxsCPLLBEj8RCzCAG/3+GlUkjCC9BuHBMrDhlzunnr3vgExwm
Q1241clddwxlo8aJkvpB5XThJN5tTjFHF7ryiHIpC6mGUngb7kiIgG5Bmq2itpIM
BtQKUzEQuC9AXcxuUPTKzBig0KAUTxEelNE2lh+z0WgUc4dd/YcCV3vHsf0951Yx
eIsD0sUAMhjNi48nX2ySx4pEu0In2Xub5OBy5dOWp6YVKAPga01qOAmwEmJqR5pQ
VbfRmloRyOlNVZcnOKDFj+Bffo/yvHQ/OYYNFRo38pQ3dAJXPSchRziuCrzIMG8i
eFgvKJlbQaLaXTaCUeJpal+mwH3Q+hKUxlktiuoJ/rT7TkzXctXPvbuJ8unro0PV
HJS0g7o/6OSpkEVI92jh/9Uht2LFXPmRbxQAwlvaU20XpGL13RtMqjG46sS22Edr
wEBHIGvuXlAHW81VJp//dkrRaMqXOw35T9Qt49GOcEPY04oowwo4Rb52TdLU4usV
idZ7nNGsIxkuKBekB7yz5p/PsQi/+ukhiOR8n15xmgj7i2rHXUbp8sSkOpCmAKCm
Lqvlk/H9kx7THM7bcARrETM5mubgptVFaYyUkIoJr2JyiQpgxfbfMSAAhNpyIkpN
XSaqY6ZydzDwQZL8BSQtM1AYvyXvLAksUdcLEtgKgGyEDpCIuvaVO4qOgFperuDO
x7T8bJ/ePjCI7dDXPF03oHmIfU1mU8yUIrqHPdR9WuFOgfNAMB+MV9U86VqmkgwO
ylMMxqyTZFtIouErqliITmE1jaHbcDYEvjve9J+Xv5pKFL4j4BBPr9N2rIGFdKPp
NBvTh+g0QTrv6y2TIlNuR6YQikgW3zzGSitsTegHNR0iaukniasb5AJ9zCfmqiYC
6bN0NP2dei50/Fwn2sSS78VeuRoLCebiNezQPsg6aRM9Qy2Wp2yVVDOfwX5/XVSx
7ET+ygUyVF6UiQFOTOrxBXW8GRoc7Vq1nFqA2IlOzm0UEJ4cVqz3vuYlTncRPLPy
fq5J0Wto1N6E13MniPa6hLE02EjJNqWCQiBMncAklxDOWWi56kCchqJlA2cvpYE+
Ob2zsuHuwtfhEEwdA6ohfQ3xeza1fWwRtc0Wa8FrQpY6PFTK30WaE8CARyA+DHUI
U7ViMj4JyqVj9QQ2KX8ljFVXZ+qkyVOnIpGh297S74pPO2f9JXk4l94ICkpKwy4V
zJ1YTXXlTrXqUouhG4l6veVhvTYCbrJ/buLnF4zHC1RQYblNRmtlX7emPBSDH2ha
xcjXf4JS27HSQLWCv7ucFZ638zm+W21N5V67pdp23/NacYVkdnjI+9kdKpSK5GPq
tgy0328o3/Cyt/ubaa8VEXO6BYe9P2p+STXsF3NSB4YOni65uly4FLIFiSsFZ0Eb
RCOwu+a/Qh1e6Vd1WgWaC/dOsLpQaJnloZElDd1Jft4iwIrkjRv/Ukx8TDdp93tT
V0f41rDAKCi9e71LkMy1/z/r5QnwWxhMAspFVBSM6ZnQa4ZMMNMyHsGF8LToJBhd
D/tC9Dl2uNcWsaKtxwktKOhT7uv4zmx3ZPO4icQmTPWh6OLMFFZAlJEKXgGhX+Ft
+13zDS8s2Fs+yictV0VTzyT/qsgHwBESzwG+xe6x8TrJAw0QMc7aZ1/CvH2cXr+u
aUax3ngbh5y1TWaM4HzpmVK0a1k7f+npRZRZ0oqqXpd+Znrhslb9YKpF6XC/hK4l
xMVH9jJS58qmF8FbsUkzhQDuIdY9hfPAMvZ5S7Bre7wcUGqO/pD5gBmaXyzeWX71
CVpz6HOHRHJTMpU/UYktfn4WcZqMhu7gIQGAZt+RLaXjoMiHZPdemzYK05nzeRRo
EXEMvnQuZFPpQd1NvRZG/VHSulQ95S299vIYk2JpxyLKICQOY/v26M3bvDzpaR38
abYSUtuy5T/etbfSUgaZQg9bE4LMUxWx0HsAxyKjbnX3CpmtqxxcLm6eonU8mRVR
Kx8FYBjGVQB7e9NKWnR7nt55M344RXQ1jQpD0maJhDaqejuV8xFmffippKcai0yA
IO/Q3jD6XVxoCqPfn6l7hSU/d0Kpcq3H6GUk+hMIMryNZ8q0wm0IDU0SQQBnMlGZ
CS/9Dn1gnJ9iwT/jsbU1zFH/PEwCMKKp9G5mEHVoxyJlShQCJyeQSkhMcXhN/JTZ
oQuSlMu5vrsflo8tLm+TlSGJKEC5WH2iBn1nqBc9RLEQIt1FiwkD4n4NDBCcRTvB
15o06UB9td1j/H6Qh+8qGdJB6pMMfXXYLdpupNTiiBW/7mlSnXHZDPIKAjfMkDl4
sE5TQ5o7MGo0HCbT248aeqG1G2Ebh3SSYM9HjYNxqVDzsaN1mD1nXutWfHN0J3he
BtCGERTAFxp7mfOZU+gw+RTRwIV73drQEu6720v1BVNe5X+GsmhQWQNQw0ppDZ4Z
G4YBMvlld+mVMBOUnHOZwAtaYUSTAmqefsONpihgXJ+GkWs24vI6U43iFgkXBSTP
uMR2Gk49Uud9/NTVwUOlBP6WCZ0TRjdo/0DJw69LY9IoDfem4eSNcah1tw/UXrV3
xGfK1c3J/1wCsOAozbuiXiutzH8bSV3M4vR+EgVqsSzcTewAB+5CYd8HiAZTdruF
cCJYh+UU4vEnEh62J7rb/YcM75IGxW8dMma5ev+v9qn3fvO+8wNIuZ2/ga5zVcu5
xeI8YdZu3n+PJZ4tFrpTtyCeeFQFSpYhsQrnsd3vET88HtF/8P4ljtTQ4O8MfYw8
VODmkjO+IIJMhsyVLfD1G8Fu7yfEeM94VxXNXdXl+zIAFRPH2yFsL7blDJH44K3C
4X5B54R6P6xaoXcrqJyjSp8nj50qR0PGWCThQvGUTDUHyeQw5N3z5hSXZ7x5m150
Di6S0+K9lfK9wa2dJkx34zS4uBOnu5GkAd/XleruRxPWKwTFUlrl4UXQeRqNPauX
JyTcXF8TRnHAyRUU/YE5GiVVivYhHcVdTmufaJgQLUiK+XlM2fTwfF8YAh8TzgqU
KKAKJxvf710KGKhJMuQGVq49h7Qyvjc9h3NAa7AFJPBCo1gc0Vg97M+8EaN6wM0j
ep52yJr2x4MjIIMNudgX+OrQcg7PlEx0/xg8iKV0XjIhcsNN/OfechKXVC45CdOI
SvTy8tl0sU5aJLB6k7DkYjt0anHf9DFt+Lqni5/DOYRA83g/iO60ZASfb6M6YNx0
4NM+Li0KosZjpOINhuifXZatj5Emp1rS05ZU+YX3U9v7tEsKA5bT4JojsPvd+wH6
tO2sVuV5uGkf8dRcT/HNGGxqCzEZKfbLZvSIpmr+We/bnVgs/LHHcItslf3qmgUm
Ng8UMuCkV/6TFBRN4hS5miFc49toOPOxswYZhFDAvBOsVp+xayEls8CCE9p0IVMQ
GnuwUQA9E9FHDwOOjHGul/L/NcOyJYO9uRHH7oxWxEtBQY/kl9587YdzwvpNiy9I
zI/uvsduy/Sq0tuHQPE4l9Vesdt3zQTWcMPK/fvBMnqwsV/P1uw2MonmAMOhLCE1
gyDcSeHk6buPy7VVsNdG3Jrt0CSyN0MN3jpr+toMDUzfsq7Dd6jMkgFDHE2Zw1P0
fKsq/kKe23cIU0nFJNcgk3U8NxOitQddSLnHGphS/bBrRK3CW1UhYW2V+/F5/eSI
vt/1++nBKIILfc5nZrkq5JHzFwUQBjsGrUtgeWKi/Uv5SxLvRk3NtQ8mt/v1O5wb
mUsJN9jLknerYV6myN7xhH+KxJQLdDF7pWT3Vvnwii6v4fJdVIQeVLRodJ5RtWph
dC8JV4mzo5igoYC7pkL/Is1qr7rnqGqRKuTicnVFggU3P6aCFhTI1mFBAJNir92t
SRaPb1KoTpuREJoP0ORTHkj50v1mc6ytUPaW62bfolv81fL0+nhzxN54x+aN6qoy
xdmJSkauwj9zhk0N+O6u7jUclJYsEHZe0q/IQWsa4TUY7yZTzxgwW/mviLgdfFuO
FQX9FGUno1sMYG6kD5K/z0qR6WImfJhXi8oLbVKZVMiysEbhwwiPEg0eGziARHVj
hRVqDHJztWc6rZHu1Xbf+7Tg21pGd6KvRtMhfyd48vmrkToU7j05TjSWCpUiJQgb
zwWvbtVYut9vag9byKw8z3KTeV5PwR7cLXb/UrX5yYn3lmbh7qsBs9cazqLAB8og
jA6bIh1+zFwyIhpF6rY2GlqykrrqQHz/FCGCMX2EprW27TonLdvgWQD4smsMdD4l
65t36hSZVva8BOAqo75AnhMCdHHu9CjJp2JKIioc9vx/jDSb6cdk0p4zdsOMaxGy
epMMLMNYT/VXoV/R9JQxjys7nbNb6L/Aot9mI288OEUg4/pD4WvA59Cq+jIBlHe0
R/muntF1djhzKhyleZ+oehpcmLu8j8Visbn+t6686NqwfKjj7xJUuLPMRSTXkru0
Ma/u+tn2hafWHaNnaUWTZ/GN6jTuJChOGo3mwzLTsQyixPI0jQGcJ3yGjd6FRsew
Eb/tatS3dK468lVsWgdD0812TB9xrJt4dlpjoa3ODlW+9o6av3s6VSYz8FkTYTz2
eKfYQ3eBSgrW48nikyUBI4wmi0j2YLKBoy06W1/ewVXSBFzTHp9Q1hiBhRYfGa+s
JqbIv4gZUd8lMLhg1lrjIzujfpZiBOvv19jUm3iyoVpSj7XegKTWphHTQPBAm9kl
Ane1RWFNMxLZ8z4ih6fY8n60MmOww0EVKGYVsowEeLm30Nlp7/JIZZBhn9gfDJqO
TqzfZpHCVbV5mvlcNejTRBx+wZHuicmIxNwN42gNR0hcd91V4vSJeBo9VebMMZyH
KtPW5nVkkzTTdlDH5IG/lWIGA1y6ugK9/hq6nNrv99xRtPFJ4D6cQgMmvzoNnsHm
YlCn/J92CGVJZI4YDtfxeB2ApzHszm1xATMh0slvZ+NadPeZxE0xEa6usUqKH7i+
zT1jACIaQ3aP0jg61/Lr6014lIlSYO6EQN2XcpnpuKzYetUDZlGlEOO72o/pqwYH
A1fpmJpqLVIFQgnF+DOPOWRwbP/T1J1ls0hYY7j5F/Pwx1UcYeAATonKMxKKLWcK
oH6eQhFU12KuTHMvmKLF+fiuMvryrB34k75Q6VOAVO4XjXSmeuwZkSfYebS+56mC
mVM9UvSglRk+igxlgZIsT4BNfdqQbG4rn8eQDgutP+jrJE0flv7rHQvPELX7CIEK
1FGKMdD3C5vCNsJCzOM36po/yr/2TyS4mT3rlyzvaul9ccx/P5DGy75ZFDsgGuu1
QO8JZjc8DL0plvzcddlJbHyBAd6iECja9qLvx6haDMD/1/feIM4oLYqX1HFXFX07
tncodXR7PFkkXSrMwz5qg3aYWmDrRGOEFBzQmpoD/fmvxqTFybYGUfuf3GDIZBGb
mlGHhgLx8+T0op5bbeeY7/cPjC2lB2LsKNM/p4a1xflHrzIuqyep9aih78yKYN3x
ug+7U1bHFhE2wPERlfQqELxkBsmviG6+0SZdXBdkbL4CXPDEFqM89v0PJFXsRgJc
b0+dd9sKejIiRU3vMwJoMrFjzxN+oX2sjcNtsX6X/BB2Zt8fb51SCGz6wi6GRCRC
LuJDflql/aHEEJLQTulYX6sJSS4w5WCSJz6v6sPSsKvHaXjSJmaewDLfY5pWvEUv
/M5omVeotjlEIWK1KY/fWyPKmgd3bfvEsgqvpzQzydEXdpadZaNuRXJ4MnRMwbcv
cL6IqFnBKUHEVcIpN4JqZdXjoqGZzQBHHAKYIofTU8K3JH3xfyQnRTfj9v7PcZLM
+E/pQdC2+HT/UZ1KjYPBas+8pBoDXQJ8jYFvdl8dqfflNnMZXz9u4kRxHUQ0JDgi
dYQenJcIqoGknC3g4Cx0GEb07EMUoSRlRtjX2DyQBnyH8mJ276m8bHJufZFKq4nq
igqYrGLmB2OOzlm7+mjttpwKLYqwVmE1JOR+9Ga8Nm7u/kticFqACKEGgXJRiAxG
8LWC3OXOLOiAAlMSq60hL0D2EN/ENnxj5jtJEQzGRz+6FSecmy8Ch0787luradpu
NxaXRkY9R8/kHdYqJcDbDFl1+ELsPsD3kjZrf7vnDri0X8R8I5yw29JkAFPp2hXF
jlY6n692s8mJsboFDQKCSaFlNtunVRExwCVPPSUPYZU/UhYsf9NHR16PbWh81/Y4
2byqAEk6QgvR+fFBBsk/U7j0C7sIBDDVNv7zL0F1x60JQOnvLSPBl7UG1efqPgnr
khLo3mecDLvWGgRoykZn9hPL83vO2lXaB+j11WUthu+UWqrqIEhF2L3Sv0aQ058i
mzRWkk6LEUKck0dhO7rw3lpaOYHt41/dQUI8dGc+ljiPKGEMO9I5nAj8+vzSvjBD
ue35Ak7yDmN19zct4eTiC+sXTeq5xxrVkBe0BzaDKeTPzlRNLgGCEoiVfLQ4/TiE
HmL0U8MIMg7clepcVhrxaNUZ5rSMnD6AtAjfEo7A3Jnan5ROwaZQ4z90GzQlHiBP
UE3/V9TCnoZexR57Ia2KXjZ5stNNZ3tXaVt2b/6iDHLdvFZwtZ02lajQPyIJ1Z59
3iWK+Lf/Ual4KTMK4Ls7uZUeWjnR+CUN5CBF1p4hauVz9b6wGZrO2QLBTiQaLHjc
uMDcqBF2/OSYiyqkhjnqVu/Lx/zKPv2LtbuyRQybzhAYO42rJH9yczOfrhNSzobv
nzlyQbQZEs6u2DwtZCN25mC7LaOKhweSSLOSiU0ifMuuPxHc+LyYRvwRc1SdWIN1
LNpipk8uWlFvcaSrkh/Put1cQE/Gc1A2S1061B4LIOzZ3V9WU50hOQXVXzM4J3Ar
PxQLiJDghZ7vNtGhqS5dr1Sh+JpVLCQvUYQ1YNDW4Cupu57fbuXSAcuXJrhuPWxP
zNRxdv4rmOhkG2f89p5wOu+t4nD8AolUxvJQGwOo1Z+ub5rAij552Fbr9bSIpiie
yp/iyNKBcqg3qwSIo9enmS4O1GNFPK6/twLXCBNxYI7LXb2NTA2o97QOOscW1JuV
f9VXOfFdjMf4bKEmCpmJz+NYCYBbySll91Tgjyne1ggXhgsyiXNW/wey4fKdtV33
g1RD3cU+Us5kDza2HCSL4edWk64kk9BJB414kEQOIsedFmlXEbxumTJmCH+1ofWa
Jv8UXv27EnGOXptXxl3/bK0g7v6YL2kR7/6Wis/zY3Pj0IdERKgtI89cgCZHHE7F
JrMMwfsk4wehQtF2Eo6yDpSIXCT4uf37rM1s//pnESQGSxnx21X+JF4NB8E2UEef
a/2eyehTrvp3Nl89sjyoYoU1/YybV9RNZUR1XlEBydQoCdwCkTSIRAGIuZf9ZCEL
F8W5Y6upaxUN92i6iWLsyaadO6UVZubo1jxIDENRwA6f/5e5DQXQSd3bozxKJgTp
QYzqMmMVZQmD2wcIIN8Liq8C0LLZkY0uhNdUyleVvaAT0U2idvS3+OM5cMEMRBzJ
7x5BPLoTsjbQdx3NmFLW8NS9UMj9Kly862zl9A2rLnaQzm7J/odAftUpbGwIQhUj
t2XwG4hojxGoTGJsIBQB3yxpKgZCzwTMc6hl+EtbXwcdk8QEnycttFVg8MgPKkzS
3hhMUt7MigPNAfjclWnGL6TDGP5UzagEACRV14WZVwh2pthHs/vhPyWj3cPMA2/C
Jk/iDgGDUgLvX+LT3E4uOBRWqRW4WyGCTWd8c0p28BYOVN+5YhawgUJ1w+3n3tRa
CRxfU7ca/AarAWh6RNChenf+oBozQFTzxvyNCHHRMmqQ2dV9XBY6ldg/0ppb4MQV
6FENb7H2qLjzTymLy9E4qPQHanKCC4FtobdfaIwaLQuipTV1KzGPpWl+yiEWjiVK
eUkABNx/wf1iRk1hkgMEAd9Obladkl8btaMLbeb949o6ulxtRExzlbLyuD77uVGT
drrqNZnOG5I2b19IWwfWWk1Sg4+aNKJrsXHryzgs6Q+Lg49DdV/d48r4XdvCQn5Z
k4cSzj5B+sd2ox6s8LmsgCJZJKT5X85LJxzK1TYY8BraupqVrS2UcwViL/6lFEra
jtN5hMbfFC7kEJ4VFieE7UFkSnmfFVq4A14yEwZvyJjtt8USNDX3w71YI4XB8Ek8
gF4U2/O9SO0KZb/PMJ/r0VthRWXE2BPGzH8yUFLX2w7WM2xEuDDTTtINlQqub0EI
F7B+o62IDbVQL4jiuWzodhFT7PhQ8q4veLqxrYuKgs7tMXLeIL/KHkAK596W7/EJ
+VY+3/gPz6d3ofas+uYadMYHAaHRznuxEozJ4/ukWykAU0qhriUtAeNabTJvGYRx
wFxwjQGZzHwMd5SdRRpn9EyBGnV61hR2/yrGQm59faq1GNfWP3HLYFlcCBZ1bA9h
HipfA/rIZZkoHxGWmeYudA04IlDFe8JMgaX1BliJJVFIEiBMUDzChOaz476SpO2A
wi9qsxo/Wg7+GNuzBjmK15xqJvt/edPZGW+qyExW7ZypNj9/p5rNcpFk0bfL2sUT
lIB+sCdzkXecpiO3AWe2NKpqjwPkYK9tGUJbe8lBhKTKUz1KGUyvnoIl9mFUdSzQ
Osww515xXoBFijSQedSfyIlW5kjmLUySJCWzUV3wxUSdL69Fc+Ie1Y0k2Tdok0Hg
9L7x0NQ9wlMwUN5HhY7fWb11QUTL7CDJVfuLbVl6SkPzFBsOpEBTnPJ36bL6eiNW
flxXmCQrAO7rkMnf0AcsxOugrbdcZzSLC/8BzFVM7Rw9BvV+mRuFuPhPtytPd1dN
e+HiGW7Lww7swcUMsisb1iBi2JbtdxSeVCBX6y0ntk3NkRkMaP/2cH6Vtdyr1kr9
H76u+Abvnl387SFH0AwPjWJ/lNG4uaMuaWpl0yhjqTmKfUya2WZr8qwkjRxsv2qQ
MlMvQ0pwSsRgICmr2N2EO4IdHUWspYQY/gcBZJSP2JjfSltaIzphinXaoJzi4KFe
ucz1cDRpuWfTtaHQMvAYRzArbOKyD5ybwmGLzk3J5OKh7NLt0UEdCK0IZe9mXFZm
6DA5fgN0l9rrgJMM9C5Y4M79j9F4a2m+MnWegVHfaieU/iOpQL2s07tcoZT8C+oU
RBh8/ZgyV/Rlkg/oNlOpUqnCALZNzEir835BwAx6pLx8XbHAnWylTB0Frwm8e+9D
kL/lohiZfEXgK4nT+x8k5OSPOu0ag7LsA/SL5uJBUlackGpBwVkUEePI+dG6ZM5Q
Q+X7Mw5aH1Nxgf1VvGzMuVaT9uo9MlmJueRCchycWHCCCFXn733Iyx05xAl4la5u
WnEylh5DQQCUS6ijjGsk+aE3cIcJxNziBm9tv9uPxddVdGiiVzHA2xojAH+Kewf3
ZqR/4bIcZgkcXNLTzXdiX1VuXk5OFxi7KMpNzeeG5QiyKl+paLpu/3knefACzVol
JEFQm9OeL9CUbCAEtijGQDc9940ESpg5OQ+HKxytl9zKSDrUsgtvw2XA6h6oXX6T
+EigWFFuohdU+opYbnunJUIDHGLYpgtbKwKRkdiirKjq4FHGwTXute06tAS3ePEW
ZvcJzgkSrWeMos9Q9t3qAKNLIZOUUZrhux79EL1jtiyKSS3h4gY1VImOmsFxZOXA
bDNjMdGLemZg3zGJYyG17zHQWdcnsYwpAZsiYbgfsmI8OUhLPdt/BXnFqPFqCj2A
mb3oLLtn38+c+sX0jCg3FFcGdEGbtPZNCQ8L8kZHEV5w+JzHuWdlpijGAbD8fqAx
rtvUvzfwZTQj3hhll/jrKU3gNvhfOAULkJmQcBKpnNOnAB5q3N9eZyZJ7z7OUmMh
s0VZhv+SjBrTEKSw8IS/jDo7Zhsa66QoJeox3DdML4sFNywaWbojjhqVw8Po969Z
9Rv6t9USLNjOi+Xv/LINbyoCFRKjOJjoQOGS+e3xKofmdzV17lQKartwgPGNkGNS
5VFBKXn9E3Kilat382wlEIXo4Vdw68L+Ec9bxPzS4uOn/xncPewpwFYH6bIzpk2v
4PhS8f6j5WpTLL30Jvrge2+99OVGhFQy5cm0itRrzUDVIWRLGzj1DQ9YGhr+LWEt
cxNhSoSMBzkSz9g1BGJnBA1tBVwWtwV6eJz+jzn35gWpgkLKzbCpyGje6GEonHbP
hFjtgQYTAObPOP6v3h16W9viOEBZ/VgGHMGM4P7IPzoOdW3A/2vED8outMkTevh5
OVVkH4up7mZcikP84kZ+S9uIxb9IqDWKnUhU+7usrclU/YdwignbpX0lF9kHkz8Q
sSNdUEe+bEwxhoPYti9TQZXHCdVk9P5AFqXn5GDs+6ngE85lL2vQPKc41fCEi0l3
ztR28spFejY86URwzEIvwFQHlPCJ7H461wQfK026HIvHFTARPP63wTRCqe8+biUT
eipj+c/T2enceye5/NxBLsI/5ByJx81QM4fqQC+hcQ7p37fffjmnQRMJmtwgg1FD
tDCEqWjagm67IrvJfUDymuDpAS1ak36Q1kHzXAEt/0FyLmFgCVs6ocJzbeP8NuMH
tUiTWbUX0jPk+yJ+w4Mbvyr7WTNKx6Rz9dkCwD7IoBvJxRnLUutf95rZijzkP8Y1
+lLFcxHt1+G4pkSIOARGwwpGfzy69GDsAU4hQlOFE3Jw64YdFjVGER2qPFuKTaRC
D6ehmp5Jmua2HyLeitVm5ARrMSIGgoTvr+hCJGOGCYSqsJHbcWYP/aJ8uGM/ZUDp
0YUbhAOu4VZytlpVxE0prmWTQqM6eIfqXE1iJmOOf4CeZvdlu2y9sZSn+FBZw3nS
BF5INFkn8QAHCNtsv1XdrmcY7Ke01TL2EMGUr+HJjastVXXdEynqeyK7gd4l7Gs7
h/QK82GwQqzGbSbU8GoA1Hj0U/EW45Fi6NN+JaVOWh4m1cbfi4EgHfKet89at2V2
TytsOAAEA0N432EqtbgzxlzrDTVH3OB3TSyNUFynS8ZgObcFrU2loX6eRsVJFA8s
mWzKl13fsKdXb/fWo1Sxz63uc6dnj7BU/xq8KDVO7bI+LRn0f6LbA64FEcX4j3Er
/xgqQyaitoQmq2GktBIl1EUZrJa/I/MW4N9H2h66XxNA05SPE7omaR2uTXy9raob
lEn9gDfoJ5zmmAAAI4Rm2fw02cU4xM+P38SctBCIHl3dcLAHkixxsyS4UQmL5ABz
nE8dxqZwyglntAxUNGTn+OKW2ZLMx9ewQMOjOuR+kJBVtJYSf0UHGgnDk5eU95jn
gNu4wRPw6F/k8CDbtKEnrr1O8NvxDswuWL8N6F2qQenOYABI8At6Pnzfp1YWfZEq
Tfhb/TVRyO4QK+3QJTrQnaWk/TjhkPQZHMRC6TFEnUp8fWxK9wX6yGfeBq0/LCal
OrhWq3hudvHzMhGh5R7vEziWei0fKvfkzGS02s60js/zGQQILsudZYKTySDxLHd+
J1yejEAmy700GJUuWZ/J2bfIBIThrxu6wbt857gfsbKsHdAnzDi6nIkBBCJf5UkU
+DRVfZXusygsA4KlI6Mw51XADRm5F40a0p5MRxonZlgyXXXtjj/FRQhbv/+MWuSL
DPIzA8K/g1qC6EnaOaIGKnbdRYEAG9eOpe+BP1GTnshGkuixAd1LT00Ypu4+f8fA
LEdK1C/vdfKxBLprnGcloADrcuh6OPGhgCyYyVsWc8wKd+jhNEwmswNliV81dicC
KIO7m8NGC/dtQXwxqZbi49YKJd9w3mD9NnjoUAi03NgwU9uqo3o3BeCXjacBi5T3
CYXSQ4zUGL8F65FJ0eb30FJvcjZ17wjgW3S8g3sIjpUCdzBbZgHRoxSJFTQe6c/g
N7nI3gPnVrwK87yKZWVEY3IZx0zAYU35i7J6bjCo7VO4tcPbcFXpG3PrGAJDy8wG
l/a/yG8PeU7pNJNNvTY96Gs5crG05RNWX2xJyWmlC2Y4FaNp7zwK6YEP8SwtzBVf
phCx94cdGpMoJokV2dDPU/kxyuTmQil0fr4+WeoDpkufZ0G6fuaFB5DKI33yKKmX
lovkgr8BOm7LC3S+aAUHJSLl1YmArr3Q02UsxTylpOK4lfOqbFXMMtXldi4GSVXv
m474nthaHHm7hlyO1IhRWIld4zr2c/qzcwkWoFt8ArnP9T2eEbjdF0SimviMa6ks
ru8NKKL+Wp7TKz+yfNgY04ZFN+6hcmr3JtzB9Pzoshcik4C7tLHCO80XCV3Yq3lt
fHHzD+o/uY752WFSoiJZ/gNZj4CwFWy5v5oaxaStcNBe6zRj+k4fzVtqdjMYHv5V
yfGBM7fQsimzABw5MzAFnwzJdOpLTKm20RidIeWr1o8EJR1FoAoyEPQTc0JH1Mv7
aR8ZlNiPMnu6lUZTDEtg5GxYSfdHcvrk5izBPGygWyay0WSODGgSUei4mCx2HcJX
xocZr0moFSLxPozXjZgWEOJX4yh0W6c7vz7UeMUBxdUbmfsC7kiDKFIDdI0+yG8M
vudO9d40Ai9BqtT6kIC3WyVCA97nXWsoYc3QCT+nL1HNe1ikJc7hXlRWa4Q9JF3T
RSnlBva4nkRIhB78nC5xTUScvAetQm1HTaKbgIAhf5GUlVm/lAyumXJobUZIrQKz
25h9/VkCNpTv+K1Od/CrXxze+1o8C3ggzboxhyDAnqCNLez2IJFxHOaLuIMLdaml
adB+s0dRSyXCWleshzX1UJGvwiwY8sqdy+vfBaEH8VF7tq6U4ozXm6uXvliT50KH
QOA+CVVbiyPv3ZvIcUcQoJzXrosUm8vFAAwcMqWnlNdXMvoV/UTzoxYmaIgdM3j6
ih8k1nqT14y9ToihPukg4GdHHArUrdq5hLIp/mp36L2IsHzVMCFvOZSnOzY4qssw
Z2EP4Prabdd3COCSOEbnmeo3/WG5UJtQv0sGRnuydve76kgiv2xbMlTHttW3Ee+q
mZtSPexxiElmENuSI+bXVnQwjiO4X7flSSVdZs/Yv2qS6IMoBUAFTW7BYOkN6hsK
eWVS4C9KagdhDahp6ZntI554aS0sk5zcgUIj3u+MftBpQ1Q2ibmTGlg7MQNpS3LL
wykuxIQkT6PpnGgQb1GB/mfIMvcktjSZWoF1dAcwYhXgXchTQNDoCKEkhCx0kfGO
6/elvUpvqHnFHJUJy4iGpBuTA8H8ajvS20zXQrC9kdpJqMir9kQUetYyHo9zJPAz
TApMRtq4a55ApljJhmEc2OjeD0queoXl+mez+vW8tPyEk2fA9k7ELhMKiYs5/YKb
ZTtkbFnaxsgtOR0R0GgM5ftKwlmrfxxhX+mGcg5TNsFOcC6S7Fo4+KUA2ZGRc873
4hEYkQGvJmGeOL3/PLvqqK5VwQ2tSa8yMJxX/gmMSiqTVTht8rfl77d6gHkhtY82
72Mmyv7FEGckWGKPvpJ4yFAsM6o2uTffTjjj9YDmrRGpI1jVl38rweXHbXm6PEJN
hv5/BHyLac2srAKDV6W/mZnQ5JIkWmtsI095zWEgz2yIFLH34Bur2dqdhcTfol1K
GGF+wjfZIFA0jm5uNz/hDIx7i4Wp9NzRZp2l40lbfc1kWApAgQo9a3wiC8r+9Z8T
rqKWMM/hyB+tMJDSzD29sphUvH5lC6S5e7eRsJs1fbbw0qu7HTdQK4A/89FDClnL
od+OqzhVENnH2AbouXzHOJEJYIqooqnGTVjaPAtJ0Z6pCfXs+zIbGYM+Upv9OV/S
IpNKjDKI4U3r/iMfKEvnSdc1jaaGRyQVUnZvnCiqzrA/DOjDGvO0j45zq7+f57Au
MQSv44OaE72bQ8Qg3FFePhfpbD1f1pD/xfaNs4vxunXoZRZ4LS1gG/O5s7G+41+b
OYX0WvQWufOVjiyvGK7/F7l2IGaE+fcYpG9X27+leEqjQmVKhbG6F+g++04+UUQv
tdq+5S5lQcsr2RvMo3dXvj+sEc8JyrKBqC0CfR/idWPAG+Wu30bzEh8G6nWbcMob
RU6bVhBio8inQyUjRw53CNssppTLOXTZONnPeOLN0NA+M3cd9Y1u9Kgycko/M0Js
3Jj8tUXuaKMbqUGFYm4AGb/ay46cK1sJgIj6zHultvAPqz+U/qVwwG+sqqNqtbwE
/zDUK53ulIvCZUV++d7AhEm0iNlaINy9vcPTAt3ys3oegYJ7KP5WLobveoGaZEyf
rHvuOO9RteGX9EMQPHZxtPn51rxEMenvPvWIZxWteRNfxoLxl5FA3JLr3R2m3jAM
QZHWCfRSY/Tc8xHUlG3uG4fPGJ+TU4UZGbQ4UsKTTsxAG03YVdAoZ72qyt3Nvr8c
Atuj/kALsj3cXVFDo6bRYnDmYuAFtXnOV/1lhVTbnu0URnu4Bc6KPmTND6Qb+vGa
nqaasBT8CGqaA6W/m7sd9sUT7GjmmG4S/gU16V3O9Dlp40MDZMTVGspEGZlc3TPL
T/jZv27GuBqmOFTbQsMQIcf8AEBYlMr4Rd90vxfe0sbYE+U8N/oyxidknvYwDPAh
Fup+BL3vVXDFYW3jh5WhzAugmPO0XH+01sFSVj2W+Adeoe3vCpj/9Y0daFYWeKJI
z7BIjRaehy11ag55a+debkro7WQaaLlLS2dbraV2aS72O+1+DsBZ2jG7efFG4xr+
IxIq5vkuEdH9v/xbIWg7XQKkBgLx33Gwj7mcM705y6EIvA+K33sm5dGEvtjNjhre
PlsT9LjrIVjG2yc+sc25RGmc6EzB4PdMU62MV3g/lujLAgt7ifmN5dI3fWv8utgw
9i+obM80dea+FumDbSd3Kz1pN3p1TtesTLhIQ+3DTMaosbZFVUxUaDiUwj9otTgn
eQrj3rMV0ES5gx8t+zDkXLNGlHWXWrIhKy+vAyJzfUJbEC1Yzxb79J8ada6cw4v/
QftyR5XpoVvkKPNFrxq59JaS+VxBJ5LPz+YqUbfCv+f53jTsV8Ir2LsXokxj7nQH
ExbJ4dzWnCApdv0J2tZ3CCNSgHUsfLrplZXPMrlJ0/oM+A8zptEAF6ETPxFEDwhm
9O0HM2PbM++85wxi25fH3lrfWce6HcsVSEs06xjh1lIpJa7lD3tD5WbNFcjb/K1L
3f9VsAvQ2yfhM/enxI8VPt/OGY6eIu7xATtpSNeRuz7MEQgIGX95anelVdqH7ayx
ow67h3KCyVs27ZfLwRS5gXtNNJGDgnBhg4sOcUgxd09BHXXRqfIPzrpxHivBPZbn
RRD9cIZMnoOkfw3c86mTNdL48dSxV46CcQHiD8jummxsrQfrSoU1NZI2tBnA4zhW
NxrEQow5Qe39OGDaCM2kcX8IadAqBlYtb6Ay7bVVPUTdZn1vLNmEJDi3mOaGqXl1
Cey3nmhzJ//G+Vzr5Oouw1O8JbMrBsdoH3JpCOEH8fuFYSOTfE5YBT0M/zKRL5rN
4VuP4BJj8LGxM1LqXsCligdsRea/iYDet1Y7a7VzihwU7G/okbDomO+cz8q+fWo8
DeRaSDmw9Jxk5ZPUVr058Po/6h0cmjsjDqrDgdblQ18ie1ALgpmQ7TbHJ9y2vJuB
KS/MMRX6KmQspcwEiNlzep9eKwwmzHnuagPPpF5lqWi+pqXe5chiPSZq9NojSp2m
H0Tko8TMGF+g5J00y2N9zoBqqbxfzyW2wfUJW9BOAbZ7kApYg5JVrIQPpcf092VZ
hNV28fSnHi67uhgT1bkLu2inkC9TytEv7UdVC3rzccbsWsosM89S6nfDni230lnR
Bj0zRUvKIKyMOsghB6qM3YgaYSepoSY4L78dBs9J9Nv3lMcKk/H3A4YIFYx8uTLE
cx8deV9o9CKuyXyAV1SUvg+FEpoCq0679ihIIoTEgPZaUmVyDTlGAOlChvLRibM7
i8jospbAQmLGO6426J81YeX+F+t17lkgFOoKQoYlVMHlAMsXN7hBv6aIq5jitRmn
ralraIVDZ6rCYD7m8ebLkxznGwcHnU9utf77DJrJEE8LPoSr3bKIpZpkEVOkjBrE
N7FXlp9aNN6BA+2s5SUYqiBVYHZdKlW7cE6t+2MkBxjnKNibYz47Tw7/3WCh92UK
3xhw0WKb70iC8h3n9Hm+URW4ujqHlvNrtKB2h76TjWETdPfli1wEgQ/O2QMa2hvg
MnsL+jJC7MNaXbPr5kGwjFoJBGIyBlXa+o7+f3GTb3HDJNZvMMZ463btsd36Vqop
DcnQYBtnQRxJm7CYHGNt7YZjDzrVQyzIgiGSjFyxn871PkExPIsclai5BnSEmvOY
+qvQq9mTsxNllz0Fzo0Yq+KpwvmAc+G8ra1Zv3gy/SEMNW1I5iN3j0QtGLDrya2x
ZYBVWiiDFqcFXacv0aDprR+X4hRScCIGz5qhGHBgs/3iFNkBgnKUkO0YzcUp5R4f
eUGWCVmXqPJynPZHb2SovDhoHw6jVecwRVEhLeCGoy9fSzgZr46saw33hHPjH9kb
1pI0dop5lN5g0PpoqqyXztQtObS5Xd9OsFL+RK4QT0pRxDFpEydPX5u6WB0aK3G/
17lWN6+k7sZQouEJTx9M9rjsAl+xHkUuC4XluujTNBhVTwGnDqAA98CfaB/687j2
nYL0uLdTH8be+POBlafMsorsim1cRsMfPoao3RmxfzwzOrK2dFmdxg/Xy3uLwAoH
eOgvIbLx1E/+SvkzsxVRFGsvqmf2TPqhcvleIeXNuELnjR7KGbUKP1C2/aJ1VPP+
qpivy9Uz2G7qt2BWpBwhZDvjf6QoddislSeYji6oiMI5oAgRuNjS7Oso15TgIV2i
8YO8/B/fnoiV/ctHbmPxSf0bs/sVyz+M0ESxjF3rBVEldc0bFL2JW5T98p9cUMnP
PCavrdMNW8xOrAfbCPBpRiolL6a7Qwj5NrEa9i05oDu5SutgHTadIqPHDj9YeGN5
qDeAK5E2Pxoxn93VjyCrUUkwQJVnhqz1WVyOTMjvvUdsISnkQsJ+7lOxavMxNgka
cRk0bJxHamMn5NyVp2xEziVxkCdseM/y0MbxYn9rewjJkeB/WlFU6kdE6UhT1iRf
s/hA5CrcMtdLuiUijFyLACBA/uraDIxZq9mNWEoBUltzui7Aq1HQ7RlDbbD2pSvp
JsmnI/PgxgHXSq9f7CZdbgXBWM+vgl+aAeU3aFdsvE9sHhiKSQ4G70c5mYN55iQA
lF0KzYnxx4ZbG/9MFMVDq6llVAPj2vs3TQPuXN7/nsBYqZSXebfuIAoUj8ZeFTFF
0dSb/is3I45teJAG1iB2tLox8UBC1a5BypwJ1bDf7f/Yk9artw0eSjVig8NAGsoH
5milCt8RhWPYsoR7ia6pAsZIZus2CjqJM+M3G6E+A0saoV465VnUzt3z/07aXwpS
jboa7bszEJrhiPUyvT6apSBH77H6vk+dQL97pQGYGCaZ6iZZFi8DRkE+yZj4/PtA
1gJztZoxVdAGT4PBz7lpe1MLEs3Hw42gDfJKAK+c+dN/8PzmikpWjr7dLea9cYmv
Fg7SpJ8TvP9t1qSyi6BNLrsfNGLLNNDYa07fposBYyqGchEeO9Cp5CiI8f+vasjh
GSzeJRfaZ3QHvw6qPB45fNXWJrM2JJkSWeN458/oN7ZjijcjafjW4+tWn7Oo5PwT
7mYElprMuQvVJyzIPqhH1uuu2wjBEtDGQUdVPvt2E/vS30deSz+mey+JcfYQs7Fm
b02/NbT4A4nurRgRZ+bdrnXOg/sDx58MosfWyGOd5DcosyLgqQn3ySfhKgCvhRdI
oAzkYGBvo9yiPtzn2EAAWOOrX4CTWdS9GRX1lcKr4K8KGcfVUbhFWhePEZpSZvD2
MsZ40y3qMLpDhaWhS6rtsT4DfFjUn7DsSHL+KkqO8b4JccO7nas4YfYT2IH+tsyL
cJTM/EWdDVa951mojDiPsp2Kw8mUcLXdpEvMm11Wdim5N1PIimolHt3i7ATVkYuP
ojujl6NK5xNNM1In88hIxO6WBLbB6D0AiXOAj0UCZrH/JA4YDMXEazc3ep/zfhcK
MQc1IJwBu9rJEAbLFSUIcAeetANzKz6FSRkiXmG2AhDVx0by+kmMwUFc7mBWB230
7tt+X9SfzYEd5tmWeNmqk+PIHwZPvzhn+X66eK1umO+FINmvlSxaercjIk48bObz
T2P6WYKlwhrvFKIsEF4KsaOWz13LSNbQMigkYI9PhkFphcGaKsB+DkXRfg7Olvuo
m4gol5+ZZL3V9r4nckGiaDO0ZpyDbAeAo1ghmbsbFzgc53baVwjC1m7ah6jBUgkl
Itb66idRNa4odrajEjwAQlz7i+H5lG2GulIAqz/Ud5ENMItSMq7YOxDPoN3Y8/LT
dL5xJlldZAez9Mwyt6v5RdMdQswSvsfWpK9cji56J6pfW3ujuueNuE9TJIhBcimD
WcGtJsJjSTq/vW3mk+5z2cW9PoGMkSZsx4aT57OspphDIgQqxB5JVnAjRWt6M77j
dUCvsjfvDmGqwJUbkzRb5wqLaxXEK7QTmQZ1qhd0CS8txtpeQp9MF/98X6rTbOc1
/dG355eRBWqWTIVii015cLx8HqRcaOoT4YenV4AHV+sJWArmvRItSUWtb4n1PJ2A
IjxPsaVHiRZe54xfVU2fWFP8X0IYZstYh5DoiEroG0wOeNH75io+BrS+bodRCS0z
CpPUqq0i8FmAtTpaLMGxxrAcUeRmb8GGW8Ym5f4Lsg6Fl/9juWR7PvsdZQyODOgc
TzI3tuQOdn05+JkBZBe0pEMflwNnweRRlX3CVDN72d6j8/24pxLxRkG0hbcvr40/
xg/v9/IOg4dZuONbvIXKEBLMvAHH0j3Ofq4ZH+BAA2RdnhbEgzEB39+1nd50Sq6p
WgUu7UOWZzU0hmNmZPKCDj2mppC0xi2pZEzCPmUPE7yOhUJnHzh+cCEscoBsymGR
UHGSnQDW8BLZKP3g3OkD06hhweZSH06doiNUiJOu1uxzKYIaQVXlxxATgNtm/lUs
y7IPahamX9B6aO2u5k3tYxQ84xZNpraxXLaSpQQyLha0OYs8fWNOJuZE2Bfhybml
3EbyxxQLTsT+IeZOyB1iTGvDUDWxxhxhMBfjltW7sKsuyQVb1Hzv597yfqAmSVei
WkWqaJPmgAXCqJ01p4pF2pNpEWRpOFBp1gEs5CI42c8UTI0iLQRSYiTl7exgG2mW
KN9ansxOg52YB0rMrQTEzYzrJvumfTWenleb95TuwX2UjAY/QCl+qRLS/ph+/Xee
p2QVoa9yYUHhbwpVvCF7wSEPImk1vzgeqZRD8rpxJNYF5DhwLKVjqO+kKyrrFfwt
TshzJkFfwJAGRc4kBnIYQASa5V2enH7DKIxwhB0bMcoyJoYZIZrrL8f+voS0VzGB
qQSLfcEzWLRI7wjgi5JFwOrfHl+4Jjg0ODDiAcP0sECxyzev1vI7VQzOawB2nCuq
Cm7pJJYcxOpixKu7BUd2vixi+FyrOhT+FsKudeLCAcfKnbVbjn1Qjijn8RXRHWcR
e+jWM9pAmz8L9uRHJpZSLHoW6RW3cigdZXx0sRNLAtbaes2NiAlyZDHhhxV3WWEF
0omO8t6Kh7+OZPJEZOi/wN0nj+Wye9Ar6nEzMTqmrtXib1Bw8aDQKS+2bzqZq8s4
KWwYjlITe/WSnf7SUrReigSoniPSey3BUSbOn1lwYVWjbZ77WHiGNX/bCSpJeseF
WCk3mnaD6l5Uw7gq7Uh+rGcBiu8YR/DhCqo1SZQBBZX83+5Le/wfGebrhkZl1q98
fpFz3pMkwFOIDpKZIKNkkJYXTYIf9ldcK71h3DbiuEEZLLVKAaNnK99URR76xe7I
pKvHoNU0KkYOWAXI3pOL+QPOzPsl7jKbOj88ASFNxYh8by5bLK5/6X8CIpFokj+r
WkUPw9HRupEfEjZ6seyXMWA8u1NsjSzUFLlpq1w2snLc/al7+q9/iL221e7d8JGu
R7vy/7zPBVe24HEPLcKbeCNF4JsRoqOlCKc0lsHECmGVT/+85LCrkQANSWMZXz69
wKpRCfHDR1VeSLNrx2pW4snkUkD0vWlZVqdxxUUS0Bt+S5OIxH2dI0CG0nryp5fm
czqHwBx6WkXuzE5PeATLUdU4YvkCjCOgVnPCP6ChUfs5K8moSB/yQixcchU4cOpt
hvQykk5VV057giZcizBN8cz1gEswFbLvG9N+I+S4y5T7gubQ+eX1Nhyo0+DGCJ74
Si4ObvQQePhCRN5IwleHin6k80byhAq+CA8vmovJSXngC3lTH8gszy4ZYDwtkc6U
Szc0T2FQ7E3308JfCllBNTDFdhW8lai37xZm/Y3Sl4Bdj3yVUEFEae2XDCj7jbmw
UJv5stetSEzsK+mNVfeOECQPuELffFwKCDOFby808TEYGf8lIpsdL4Smfk5gkIvb
Ry+JRRHMOQVGp6TOk25EPmEWJwNohI+DkZqYoQ6fGTPvYc7wi9d/PFC2X8CxWJPO
OZfPniI52Ws+qGaqCygPQTNwovDj/DVM8BhZ9UdBzBCgkL/ctl1OiMyrKcQXNP9l
Dl4dtH+b3oJDG+bmOkBzsle2nX2nPJBb8CvN77XmhR1qOdBrEQWIjE9rUfKJhYZo
3ge/VKvN+A2uHo6DLY0gpO3jmHjKkhJORiqmXPcLZ/ROgq9FmcFuLiWnRe9trpcA
7D7Fy0hilUghm3EVSwRtUIZovCyhLtMwIx/rxxHN7GeWOqAhgpUlyQyfzhIoMbeN
ZPHvcXSZfuwfd9DB/Z/s2zBEmz21CuGfH6kG1N6KMMCRm7ePdZx+kwJY1mMA/CNi
Yx0zesE1TIhmgEfj+wAYyqsr7oEroQvag5Lh3vbAQnef1YMdmjbQdGXXLJ6XxATW
w22SwAj4O9VK8+AgvL3EwBInXhdAsIkavChQevM+IuovqahZYd+ekoy44hfpCArj
aH1GexrHuiyb5k65rmM7oJPiM+UDbBnxCmyhHHPqHGmFrQVG7YyTC0Pro4aXffze
mW1HrfJwD4rmDA36OEzjEsCsXaYdLuu31wsc/5J6e+O7y5ys9ergGJwmSuXpxEgS
EP38+E0gNgbk00vMZjbAtWkb0Cs3eWq1qQ4NRXNvAblhrowWdJhfxS419wyl81tr
3GfNKTgXQeA1Iw3aH+d2xx7U0mOULYEl9DCt8Pch10wDS5/ggMcsQ4WgNUraNDWJ
H1SWMPoBDRUSjCGDuyH050p6EFvrx5GJtVmCrQslihfzBP1AG65lolX3NAR6TXFv
5LgvOA3RjwcXARPEHmsoej4Mtk1XUOIIIxk98+WXRA+1Ahb+IBpq5A9nuPE+Fty1
c4zmSKqlG0WY0sxx/BCgZOj7X3tOJ7gG+QhNxN2I1Y1aYQZYI9GpZ0bY+MS1Z2pQ
l6l9c3U7VWq3qf6uzMLB1DaXLTwDFmJtMVXfzMY0U+WrnBc7Y0Eb5P9/Un86CTkX
dsVCnAAnABBoTLLkwPrHWNKIK1VsmbBiVmOSpJvtpcFeMDkAKp7UpQckgtd4kswp
kOSRoGcuA+qyy4oREreLCNpbtfJ/4HToL3ybGJIMgHBwp75q2xlTEQmFiBDfdJOv
kA/TynPWCMlYbtRZBniQIvb5wUuq3thMVQGLTTdf/5KN8eD0Q7zPbQUOV48GhePn
Xcv7MyNxhh9KQT9ydlcFdDqK0NGSQAsQw16pEM49JHn+qSWl2O+6ohj/tPSNum+V
n3A9OIm8jSbkc93F4QzeAjxqih4xWqffB5UVEriel1cikRFI/CDZRXc8F9f6QtiZ
A3uxZ24AB0POuwrJc8D5lw9gs0kxGvh/MMgDxYK1syRmNjcsfW/fwzUSHxUQH0a5
Y4DFlJSo2TU5MkeQ1Y7VN9WDjwfBsP/7TYWTfUN/tZbXfws/MFb5LH1CGZ2O6qtU
CRyuXNT3kS3kpZLgBQnTILiDZXNwI6gaDpSVwyhcA2ViOCooxqxc3o7XveuiYxiz
0vEfLMztNbRt7RGiFeFZx9UpdScggkw2z9SYQ2UJ2VjmUc+CwykwkemPdnnOWZYp
mD5NWME8UXIP4PRNeYTzT7NNjQovpjFqJso+m65HqETR6u4sBU7KRRxdzcQ3OmeQ
C9BXkpUVbSftvpNiW7rn57bMxkr8pL4kKeCh6ESaI4+GNw/Gg9sPWtAx99+BIMuA
wFRtM0IIU5dcv+6JCiS1H/CTUcBaLeSENl5wkeR5YjZS2tWuKF0/LsQGKZ1C0H/A
yCPrzD4jVlxg2XtI/YMCibWxyIemvznlFGHqKEGlHb1+5RXI6a9LVv9TfKK2auc0
01JdyF4+Q37go84pgrHRr7yvEO0yLyy3anmARZSCx5NXoFFkFV4wWromrUVzeDP9
gino86CGp4wswf2QBN8cOJrKh0aSj2ey7m6SKB3BXEOhpjnM+a4mLCWKKIN+g9Ka
pMb0NmF2ZVkfAMDePXEy6xsatN8kGwxtBnpYrD7m7BlWOJm6CH7CMb1Mlh2peRj7
RQnvZaeU2b4HpuEICVhu4iHx+aYYsOc4Rj9rB7D7ySE4AzCTkueIl6nwMq/PNIBF
zEhKSaUQIam9ihuSMBStLlHM1h5xitRJrMoRn5NDX6OuvxB7tTqkOb5+KTPJi7jO
YS2EiVEtJEz/+BYMEgsu7vap6mFcFcxfjxfydLwQjkSuSaHMiCYHXfHGyaK5Htul
ryZtcg/qHXWknje3Sv6bTMFSHEySlOjyBUzR1CxY7TxbZWNPFfjoPv2rNBjWEv3t
nIztypySgBlUlmyE8ASwLWJtN8WG3QX7UkRy5UgC7tGOP1MVaP1d+QFxFCO9P43m
G7+B4BACxj1h6FwRSgFOtMkVIiBL1AAddYYRWv18Kk2FzhVywNwDPKMl3v1kbmXS
0Uc9K8hn6Ef4Co5Nan4bIHJ850iMI3C6Q+7fta3qsPyesv5M2AwFOV2p+1PbD/GV
hJqmnBhAwYlljdI2URIbrvj7yGZ2DqiEyifIhjKMRG3CpmPRFCYwxDlzCimBX9xW
+Me+xng4cHCx8tO0Y5YPiytOT22nm/f5JJ1Qygi2On2gamLqVj2zqKj+7ya72KOx
af/dBdQY9b3mgfcxTbqNW18GTpyZOy2xildVRV81WhhrBsIo5TQFOTScBOeKXBmo
7a0qZQD8g1mJNKsq3GPytBOeboKbEjyh7+9UPg2/jYCMNcIYEM4V83nt63K7nyhe
HyBRkLgE9iPPDVv3O7HCXMVcsVqY+MgV1OMIj0k/ydqXn7jSXyWXj99ewEFOdJp9
scrHh2wUTzSgLU/kwyxtwiLgfZ5Fz9h3qsnJugw4y9FGCC+GRdEcZkd+Z7JFTZoy
ZmyZ/ji+YhuSIpFRd3s1ua7+nNXTjOXMyQpUmORDACKZM7opXW/o3MHZoGHOMnxU
jt+h7SJLfFBr4v6wNuPWnDuxIDO2xc4AnWPHO3M7mhr8d5SvxftmkGhtj1HB9TBX
i64RPNfxZpRWTKbkn143aNE/bWsE0OTXHoGEVnmR+DIVtH8vLsGZJdf4g8xk7KRW
PV6rXANcmZs4gnRkhSN1Ul5fgv0Uh3ss1xNB2X+SEPwsxX5XiVIxQAL/hm+UDOva
zAMgyhmXc0VZ8DnHSAf1/RBulxUTb9UzvMf0vQnejKkiSKxrPErxKmJw5S9Fa+OK
Jw0ZgHhTPkwBvSKbiupW0Irw1szplW11ukk377CjwSKwCisvWidY3YVJhiwzUy36
JYRrJ+GiJcqcaWEqXOhOVIZNbgZDzZKgYJNH1XRU1cY4sPC2qydDI8wdzU4uHuFv
ZDinNJWG2Erx9qJRIkwKbFaAFFGG60FlfqBwGxRgM8T/1Cj/8iQVxge0z88eiTx+
tm+Q7so0fF9d5lni40xCitz+pJx+e1ODpxBwVgvwUOrzRzDJ2pfLd2r4FxtbQfDr
0Qpr9mJ3AR1WF7FakHgp8Wn3zYWuB3TG/c/VSAI0vCsmyW/WIfKLter5FL9cJgVM
0XfaW3R+ZihgTjYLVbjX7acSfMTvrn9zBkeGeV2EjyzG93fvPuj8X6NBg6Fg5+RE
nEEwQwElHLLIYTlRORl1lFyG6aZWyPMnF958gQkvlTmQ4D2i/rffdMgeMx85hZWR
Sm+WdI7xfOXgYofcjvjq7UmT+JMCHbj9Xda1rqNCiXUf5dVMgyZQ21wtRIoqFAnM
9hrbctLohWx5j9WJ/7aB7UDpb3AjS59KnVzeOb+gvAh+ktyXuSEV7mZWrgB7KkCo
rvBy0xZPCLkWEOh5yrZ2aEd+4VaGzGcK4zhFsl8DZOxbiGz0hHVHD51ORGRi7ZPb
jOPXiF3ArwXJS7H2XfnSJ4k0PBKejdjUBk37j9rBqWIdF1kXg4KIKwLM9ByCs0TM
M4bdZoPHGrLOaIn0MAqFNT/jM0iI/4gwJTMGoqTNYD88wj4UxCRIQXdQOVUjfr7R
19OYXbpBVWOrTezy/Gs5WjaIpv6zGPex0D6kUY97D5kjAbyeSigkSpbC/EifNqJw
Brk54V0nu88IRhVZSpOtCO7cjZvy48plk8HyGIrwhYxNN6f3fT12sI6CsD/w3H+M
TizbMLeBNjdAhR1b9DY13F1/l9CyuUVacW1iynIQZUCUELbeuW/ReTeVFtlggVgV
QzB+pNOPKKXhInEJXm1U+Vg5kMsAK+XqOgcKmi8HppMGUFA9wYp20IVJVtqrMGqE
7NE0LveowH/Wh69QdSUhQlMNPrSNv6y8ST0nxP2zgdPZ0H4Nv2tDIRt1YZqozR11
K0pDqA3CpIAwbcUx8cTknAmBM0LnRWWOD79lf0wHrqxgPQblYkD2VPniWj25IKYS
BsSh8NxFS+IH/zBcHXxV8DujBK8mXlzWOA8XN4oyVUi48AAibL82uQlnCn3ErrKy
rx9DYP0cRSgk50dphx4T/qFpvpBE6UwxkC9ZPLYyms4NlwEto9T3G5a9uZly8NJg
POn1u881ZfNDrKmYu/I5atfTh1FGiAU918PrXgbpqKiYYoE2Ipoobfxufk6CK6u7
Z8YsF+XYI3CGtpj3NNOxLAGNrThpwNSUxn2phcjNxzfQ6Iz1UZqbujQFQJrU5D9A
Ksw6kCYN4y0SNvbcF/OgdXo1mKTo5qjs+Lk2E5cFuHqkWl7iAYOMhOshCHo/0hEw
52tyAu6TwubTj8xoDpht9MrTVqScGgbAo3GykXhv9NIX3V+xxM0/gV0bPK6v+edI
56mNX9RkzmkhySC+MWWwuKYqyICqP+WBzqLc4BZ0URBQLxEzxbwiGGuKdDvP1Xdc
Qd5DKqdBfgBNS3NEUNPi4nH6NC1+YmIQI63N19QT8ygp0PCXEBCLaPl/MiybXqqX
9Bk82R3GvWVUen+qRvN9ohWAiRFsQFwCZrc+4gGFezLCIIcujmPz/jSj/m7kYzcx
MTPZv5rWFORG2ZpvIFEyqL+qc4Zkja8rcr7QHJO6mVF7f/unQgDDj+sW/5Odt+f2
3pQ0BcqFk26zfkAdF+cZxjUUyHNzIS5sSRSF0C+ycD9HttaoYqPjZMtwJFihhyBm
KNXPaNUjoclGWbFrCSDD4bpbsLxMcPA86Ewl4ttc2RFCVGiUH2Cd8xLfLG6tA1ww
bsSxA++gn4GJJzJrBdHRtaApK0Rgy+SQDCwcJnoNnCcvAslAqPbYcE0r0wA3JK7V
T6xP40agVRCJoMi62cxf7wliINNWci2Rgg4XXmkwWtnlNUfaSCieOPfGef5fZMv6
a5hgneHbT+84I7YSXg+WeqPCaN12eQhrLrBge29cFjdBsPNNWOg2Gr7+ZBkDy2K4
HPjHk4djmd56RtsVSo/PpUQDiJIX0sdsvjs9a+FLmf9zOFRha/6EKXTHN4xWft3T
jPj1EMoLTg6uMORQ0Y3l6GAYk9mrq8WPL5b1Dd/WMKSuhkRSpVXl36e/NuKfWedY
iERMFt0xkZbfFyA36s9mzB7zggiTmYQNfBHFAWhViSQz0f3HhW1SFyz+5yVMHMwT
rUzNOpq4LRW6Grc2XRVK3JPlFtTiVuGLDBBOwc0jfzVYSg92a3L/mr19mv7+a6fw
7W7SL7khK4pBz3eu5YMB2f1OLHmp63Nq4VhF2jnG2/dD7ns+xTWJamTKVp8n8oGh
Sh5qAckmxA4eGSHFTDyEaJtoy7rn4OWYPP+wnhcOm1Mc76woxGPOy82LAowY0zvd
o3z43tSRjXovgh8dAtSBc/sKL/YjLEy2f4rHKMct90va4EDu6aDbm0/LwVstDmGR
U5VQBcU9TizCvMH3t5HBij6+6cBFll1UkhgCZ4gdbYZrzB/wdQYWIO8NCd5PkxU9
bkW7G7lZPNZcvWoWRK0QCF5KZw/STsUbwoxaYlxasbp9gtkkjcwDMiCNjtmHFHkR
oBSA4DGOhQneJRC2Yoj8MM6XYVEhQo8Qb2Ipzw4C2/okk8aj+S4CvTq8/LtZoi98
mMFGXmJa2MuE1d5J5E7idqTHNOm95tHFTYQJ8phrldWpwa+0VHtKc/RUuPNwP78A
yHyY+YXV5r6ilF/ucvtrFie5GXC/SZw7IhkFlJrndV55jZB4ZSvdcMjsH1nbTSlc
/+9FWbKCzP81yNb4m5Ag3JQJT0mM5mAIZ6s1GJ0B2bFPuvROUcoPvBnrle8owb2G
jsrwa9GxKBE8bcHIz2O/hJu1ZTgNjmFfeZ1qGmJPQ0dp5r3eqXjzZcRoksY1s8jJ
cIV3iOlrYxoLkerJe0P4NvfTPsTYrws++L7xNrDxu6GoC8R8doenq9g36ma+vrpb
yrxwGH6ixtqPxYq+Rgzqg7bR7nLxI2NNz5tMIpJthbaK1i58k/JcdN6m8OTVgOag
Iwph2POk1gRs+Yop1535HaquQ/ozaIO2EpCukVDw+jdrJcjqD3NOb1zFbnwmnzbt
MUNYyMaAlvI2u1piUJczs2cGi5I6nCoR+MIVM6NRO34r+QbIlLN7EvWTQJgFzuj/
Xjcw58hmZiiiiIrd9fsZS830hA/VEt9uUWz2SeRqNUfRKGxIxnelnQZFQDa9fkxN
G5l+isUTyYIMRP6OGcFPQfF/IwcETA78iJgjrfCZhfjXzACCdhtQk098SwZwbtWN
pmwWIqZJHYCIQGQX9gvaEvlkyhPDmB2CQX1MTYMHBZ0T4wQV393CNmrShKZa1r4j
T+bgysDf7k5NZoIwb4DrT5fXuf0W5wkXDUQtthXf4okPDZV+4WdZTephMHyxMrXr
YyehTS43Buyzi3J2w2VFrClJrqWpHlxagFS/fQ5YUJOV3o2qgZ1CjdvRZfYlzMA7
9eW0STPGcrbyaU1PZTtdWSsj4XExQzzuoW28DVJbJqEOwaZ2c2ehQVSjtMcg+yet
QpXwVH7XtxygOJTiu+tmrmdsG8emItU046GPdrfNeEOQn6Y0OZk06qgd9XRtyoHt
xvEe2+XLJrlyZA5+dPlJAidLSYaECdSEmUgDzK17K31h39JVxe26SuiPE4Wq/+5u
owFjcshH0PWEohh0Gzuqw4OLhDyXKxppZle4aTnhJbb8FdtCdbeW4VtWuILQa5RO
XYq9Rd8aT3/mNlxJbLfX/n6FZ0AyFmAEom6gSFe7xNW9bjWHu0uVlQU82yi+Pdzo
4pwgqKUzQbf8t9gCz4lL3t0L+JCwbKAU+JXihwo+n/bO3GgMFi+59/Bj9gwCvOKi
SPFsGj9uiOvufrnAzcrqhyb2beSt0W0pFOrKkJp+2N/yjIYa0Qiwk8J9T9cJUhVX
YzifBA2CNtnXdK9bMzSKdnXnIeRFMf3jYBhEQTRQ0q0vlkt00W6/GJWzPCmwCI5h
rMOWOaUqyBKfHp6Ps2PPB8Buhe/PrARzg6yMkQ9iPBPZgXP5yxTkwxdg9VZkgCJv
cYxLKDpYKoyLI7qJK5cyV1Tm0FE2EldWpwZZen04YUoCDAx0eAFu+mCCQTBhJSax
btPX8bLAu2n0EiYvXAg214ilpsxZv48nfm2pHem/w6xXlttiuWAHrRU0aubwr75f
ttVL9c9trEWSBAyGiwp5dTArGg5o774rorHv1hjDB6EdrN1ZRlYUmckJ8QfyeoEZ
yL7lPNvxbeuJDxrOGgxsYqP59NFMBfjyGvFmlDpk4mseHKhw/eyUDDuFXyna2Mef
dFBc5XHRfSf66RC6SH63wKhm1+AkjsxgHJJSpXXvtLti1S0JO5E6bUbzaFZap0Vi
fgKWWt/ZdztIk4uHUpko26UyFjvmAWfMTxVIhUsTLRytDfTVhMD9Xf0l2RvCabMP
VSckixJVr4zVOUuQycmNWZkDzct/4OncWYOl5lVFZFPWqxpIv29xeQxA0PbO+Bir
0KGSw2eRU/nSXou7cjGnxqPyjUBj/p8Gofy6omt/zuEl4Yq4Dt8qc5FBFOAMo112
xndv8I4U9oE5AOo6jG4KhVHdRMPceInohtMISq2M0rMDpVTZm9guhef7MOfBLTcO
7EpL3cF6c6H8PJiNr5khiHiii7ZSo2jCVxxszCjxbY4Eppwlvpi2r0cQsCLwne/X
mySIT7nxLnjzE3EM9UlokHGQvlEHuFtoohEOKv58Q5mNerMu62HH4IChu7Q1HHYu
1g1gFdCnriXMsTSVXSPKp700/eHMzgD8FZyf9oZoQiVkY6Ml/pp2SckBVUXvfuWg
NSzQ+LpGp11W7b/GTnhUd4v3NWx6T8BPBRWADwag44A7HVbUMYOdUSL1SAaBDnGC
KvZNv3YyV2uG6nEtn4g2rj1zhCFz/28sqCb9MILSR06VWPpgsFaUhjr1Ce96w+Jn
LFElwM50PnBhUVO2qSntDSuluUeTDYVQ/JDsVTeBg7ZoL+nqkTSPxqfUktXjIg9A
V4diDijNct1d3FPYbd4RCHgHg00MwzjQR2jSiq+nNbmUIGsFuclhy+dNV1SQ3US0
8sGUSprJBHBXp4SEM1oHtGRokUSWucRqTsN/LnLM0W7nOVt9RBkJsho7ypqgoci2
PowO7Z8dDYzrJHHh+UEYcjtriK3B6LGQQwzoamrj8zor1EAKeQ1HF7Qsejw9doXF
zGMjUJsaaLjEbQTdAfHcXVpNmYBXXa6JT03SfpuGD+g3fbAhsdaJ2BVC1SvPVUL9
3HStrNwdF6vetMzX3cugzmD1THvtsXW9jU3t90Kyh5nlNgZ3T2yICN1iOIHRNx+m
HyB2YT3M615xAVhPx+mhcYCsuYF+qjP7Q2MYMCcqZ5ZVy45V7QioyCkSdwsv/cZ2
zmIspfu5Ngzw3iQftn9yEiIPfpPDnOAT3HEBtJmEkJn8yHnATwcdmQ3O89FdzDU+
NTLmmbkVnxM2vVH0t+pi2P5j2P+wWG5ryoB5v3pBrcH3yrHAUGQyeEG/Xzh2Pp8X
9Xqref43NGhz9+Ooa9QgcSlbhtvJAXuYXdMD47m0EFbvBGosRXQgjWAbPc0xnIL9
ArjjC2toxqVLmHuljHN77P7uGeqUS3M1uBhhg1c/GfPG4AaSxjwXyhSVyo3AwwTc
QVWiq6BZeXH8BrmXlFz+jAZW/3TKGzG+eS0xpTlsPlVfIdqL/XFuBpEpPG0L30fK
SaflZpUxBwk+HkdGNKoYAJoXpprZ0yp1RKagOwyCR7Yvez7GZPYOoIqCiOtUcL5R
1Nbi5/aihBEIfvxfg1cFJZM/gVZVPfTuTgjtWTbqV6qYA+VtwCp2CjFlZWqZbpT1
ikznciFoIn+4RKTfVFNYfkWk0OdjZob5NBlDb2SKVGkKVAG4BDPjnbR92Fa4NddE
myv/MJ8l0gzX3ysfVYhsOFbdshe61oBqfHqMERuD7vxX9rAgE7BP3cx83SZAi0/j
rax3hdtlvN8YgbDU23QTcAvJSkUv8xeFMUOUFBtDh48uj86CVTrNvx6oReCk34ch
DMYTYHZgxNOxMAv1sAw4WORwb0lqeqB/LmcFZ6t/c5ljxC+r9cbSXGSMKzKlO4n/
KE53GS/+Y2cEm35fycG56h7VCUUtqjNNZmnKJriJGimBSV4Wwdz9aj3apREVZDSq
Vi7/JkKGcQ2OD1lqOsudzaeToLce+PzHdyNzd6AUQe6BQQOXZZOBPPE1wBk/mzLY
FFecOhhwJsirNyF02jpyut2eHM4puefaJyLSkwFLTinvWQbKpjHcpVp1E4p+SgRj
vo61giSl66QXiFHYsnCvz7te7gYyiPqCAiArP/V3GzsU1AWTpajsWQolvC1T1Pt3
umBRIInJ3t13mGGgNHboW8GLLtx1Fbp6Lt4bkOcJCpn5qeS4aOb32saMObZEbkuZ
el1XyRr05jn3rAVlMiSEMs/8jJQhEftRbwzeMHbGWHZ5GggSIol6MwzT0ymbtM51
aqJ7GLaCfkw2pzTtWBriux+21do+4+PJ2XljtjI1fRmvMAzvO0MgqJ680CdXHq6b
jMGA005VXkzldlX7Xi8frIESWqECNBcmg9zA2Yv9OJ+gP9yf05PmonEibH7f9G/t
329oyvSXHgvkXkSMxIyX9NGT/VZbLhgMkSVJmRcrPn0FYXjkLv2C/c0aMeVYvBn4
iAa7mtd0AX49NXDcfuEp/bkm63LN3XiEthgm4sxPcRVzG4PEmAuprgftSJ7TAygv
Myep0LjLRErE1eXxZif+jkvMN+g6wfff8N5t+oa53WiI1iITGK+FUGQ8+ysgqvS9
nlXUkunqWh5C5n/gBg3SRz+VFNxPh/Rtx0HTpEJhiexUZ4ta2lFpYbuKk+uwcSlj
uDCnrpJXhqYCGcsCUCGAhN4ihXPnNgVODWwuDRR91BlQK71oVTrAZ3sateZdp+K3
v0g91ULdvw74VFA3wNYhZ7cXDDzjDh7gW0JvsCCBSB10SCSTPano4/j2Sqa0m3cd
x4zmsDAv5/9aJSY5amtIhruaZuHSOvY6ksgwcNxk47wjj8IBnIhbnZtoHys1ZmTO
wl3xjD+lq+/KF1uScvGNYPIyGtdmhkA+9FwZN7B3MIbjeKWk6WazrvILQIJPja7x
XqsA7dh9sAdwddAv8B86lLBZ2OgXdORlo0MVP3+5tnvK6aSOoEGCCSVFEn+pMCuF
PSYb3plhUbfTi3xqU3mBI+9mF/j8w7qRRzMx4op6nkCXLOsSihfap8EjqRu5/FVa
WUgJlUm8kdbmu+myzpY2V2C60boW7ids4kTgUez+PgRtjbjVbQEYpDRr902Mffrq
njPpcwCoMtj6ugguQGfNEr8uvZ5JdFFU724HQqYNcAR9fErp2rjYS3y8jyiDAa+D
sxdpD6gCI/dJR10HEyq4shNz591yG8r3u8l4KlgLhwvCmC64+BlsSELDmBGYam3u
a/t06wKVNUwag+pPW1E4HNsQupRfKwaQlf+d3nUWKkvoiMCEWQA3o4HSRGp/GU1F
bSQDteReTHZAqC3tlhajqrIOLftSu5/0ys8Wvc/q5Rj2Q+/w9gFD2Kew01aieISb
00iX6gR/AfsjUxOQIP/4+RlUDfmu1XE7STZqkg2/ylD3lIvaBlGfImzAUtAuh9s0
o0/I+07WV4mw7A16/dNRtjvRHA0XEFwkU5OZ5VZoVAbgAapW9nDiI8YwtdtNkJkI
beFs3XJvc0n0Nz9wXCfbgcpA2QaA2fX4jMnks9otp4JxFdHbkZL4I0oDD9p1kid+
wNdtQIxp2fSNGcyzKMMOxqYlfvrz7Fsn7hhqk1UqxQJFa++3oL0PP0n3mmowt1kL
PDypAuOaXoOIApT+Q4zdx6I0Xeb6gMg6i58MuVz+d6finGSHwMIgqJmZVMJtriOb
3+Q2cEg4ANUkAGvubOJeprikgKHuJCqsEcpw94cL0Bf2jV9csRPhBKGXkPGSJRnb
MoRuFSBXX99balxTs0snaji8+bdbU9IRnCF2jG583Fm+bzjQCGZ3U8RwQ7bOzrzQ
llE46D5GHU7rORYtz9sLF9txjP2WFCCeqpEDFz7qaIiz5VPa5o7KsaXi9jINAEKB
MNAfFuvC9D/WWxh/do7yVVO5/8PTxk06mPnxl6IR+0VPpavisYIGf0U2xRjMczrq
mAq8+BywFatlkXVEAua+bToXqxzLyQ1sL4x1fu8itRdfcI/v2NpPYELtAz7OsLET
P1IDQ0EBKRo74kcgWN5YPlKEidWLqxRYH2jDIKyl48c7dhbEZ+SfyFES7X0FcHYf
lYTIXgeCCJZUrDlVjyygOshL/hbhsGuTm+DqmX9FmZ0MZLHjv5D8rf1T96tMQX4I
Tuobw7LA+kgWkK1k5RD4y74FzyInVhePNoOrlNkeKD/b/PexbQcuM0Fe626+pUhc
M8JPs6qzc8Gy1zfEGMWa/e1tb3WKiu7lf48Z7utzC1tdPMElj9p/r308JJRneJ6A
0Oy9M7Afcxn6rLpLQZbtIntbvT2VpdEw7pQ5B2Z2EciPJ0PN4Aws+G+OsBWGSOfA
qEd5pQ9KDxjJRS/kyMuX4kMPbsl/ELCUMJLLRxoqQXohZpGmoVObEsS/FA4cBWCM
Rw8PqmyQtDl+JqT95InFv8jJHPAk2erAbKJjMSi35NqNxo4FW1fqEZsTtr2MNLw1
2beSs6VzAVtW0H0oQdzy1+qnz1ajmOOYmP0IEy/hXQVKMpNsYDNaSPQ4A3SXkRSE
WgziFCdCv6Wxi+yqX8k0NtpULfg/Bz1ZVUYVrBhT9xNMYbPOB9+HhMkbbJf7/4fS
1WR0SLGHo58anSdQ09TKthp74kLJB3YUnORxskqPENq5oRnMAjFy+qHdB4B6L6TW
PYGiCb8APoxEw+pvV7IxX3d8U1OCcfmLZ/jbiHpBKUC2N1cVJQYILZqq7ctbqANI
NKSxxDjvBPmS8vcrPG3ZkYsA2kplwvHmdX4fLWlDZS4+SmYG64+FQSZKKCcaM366
hYNhJ06oYigM2ihMh6SOevxUhbsDC9OkfHA5r7vczL21vEDZA+QtXbRk+iLI85RX
ZhzbIDGaf90BCBgcUsvUe9cWgTN9Yj4OakXMoGU6YjBFlWXlQXZMX65CP6Ml8FCE
wQESyt7LrNF2R/I3SAyzpw/RIstcm1Qnh6rvm2vJgc+/NYtHvcfoGwe6Pk/xY9GF
I6xT5lFGT2yIJHbexaKVcmAY9l/rq4YvIllFhtkY2muJyfZfHgEzy/ompUQDJyNs
ZDKg5gNoDvfFTFb2aRmVP/dv/iJf2wskz7s0jOpvtReIZKMdqlPUfkK5oyWqJ14i
MdsOijlbDN+Wr1dMeYo0vB3fSAP3sP/vz/AHEuKyw0qWh6/z0e53Ss59DkYOgKt5
bqKpglMI+xshxacZtYzBK0FJKixPUI4WbMGQE7w0N7X1794LKIBNmTzFbaHrQFde
kGPMg7hx1dG1WMdnHiLGrCR0EfMOd0JRs6xxnp54FD80+1jwgviFgmu8Q8Mxx2/1
pf0l4u+oXPXh6W7zGocTVHjsc7XjItZ21CAXLqMMvHnPZJi/RY3LH8VTMVfrv9Dv
dOE6wbEej60U6XgqLzZ2+2Sb6PvqzTB8IVZ5EljYDmKPwSXaG3GhpNfju0smfHVx
3waRi5pfUD2MFsja9epyQw/pg/k0zJwJYAN3zHz/U7Q/zbUuJxbE1pXwO/xby38m
rjXgyvKAJQRvWRKQ+VodOcWZjT8DlFvzw9l8zipYD2Jv1uxpQqXY102vUR2S/AoX
Q09mIq32IcIOWuzh4cX8FRFjMZ+7RyYXaWh7UBkNBRQiHJtWnffOBEdxaO/IYLOO
lWKhBW4pe3LNBIZMIaaYM8xgBHX1CWLLVPFuxvmN1VCZegMzCVq/+rEj4QirNoYl
yN1Qj9TjlZfwENitCSzEgg5BaRq2BXUWnv1R0eDCdWQ2vu9xBk03Vl5nglagCa6s
lXSfBzHR05mBBVzB//Bo5eLEbD+Qg7E96TbvpE6yZigdol8U3TP7bgZ19rRxiuuu
PUMlFwp2Mi/mTlDLEupg2i1NEGs6fTI6hX9OsfsNev4TufFO3qYVagZB6SopN3No
RYKgt3M8BxYLViSQ0GMeQB+1sE9dmpIWpTYrDRq4LRvin4seKjongiU5FAZ+Nj/w
Vd1pNGtOkYTOAh8edSloVPg8M9Dw2Td89XaneR+GZWhSeNHT/4tl0fPOH0FoXaMj
I/SSlNSka0ZbM4X8t/Wyl2Up48qEgmsV5HYYLkNTS2T2R29e81/epS+DI6OCaLE0
ITIK55oCyb/Ep8H4Yy3VEsnltKNehx/qbiGW7P48aJA+4tSTqt/wF8TuCeCqogFm
kIegyh1eQq38QpLc1F+54bfx05s/5t9B5E3EtWqxUQCB6tFkqCUrrnM++OxyN+Ya
2Txm7XFzumjZPUkicOEgEGDm7X0GHMUAAm2jwmF7s5LFRO7H6WkxgAmkpq/14ApW
cf4v/I65pOaXEuEv/YOWdUvUdWhPHmc39I0aqkxrtblxcFZ9VJSGrsrCCZgHUaDY
lKtYzL2L2NjNQ1WXgLVNWp7rvMiwGaJ4c2LMteHDObkJ8g0sKRiYdaKCmEt/Nc5y
zcEW7dAWjrA1fx1eicORqGe8V0d09JrDKEYprVAWlUTQeUlWvapbO87xt0adhyRh
QCgOraVmT5EjoGaY3q5/Bg0fbaZLfgwQY+ATsfa3GUxdPHQh0lWgq/s7FJGouj2L
uAKXzflNs836oJUwFTV1hwzlY9aJyPGXldz8DfsiLTLadAkLP6/euKYuc3bFHAAF
IRAMRqdsAVl0fFcUcW8FchREjvXx2z5C9LA8gCprTv0bXhQMxdcRcvnGyN3BJ8ix
pJ/uQIvWz7tKW+EXmuUSd9uYt9WpXS/uHNVXkLnIYIMkdg5FSvzVzFzt3WyRAbv2
e9ZkAuVBBNCErx0rd+6KeFPOUNnFbXVci4CyS+JX/iThifJuEGsdL2WfTq4GuVUo
0uUyo5Uv83GwqXpX2xQOpQ0LvzjJynH2vmVI89eNnbhZKfOoenbd1YFxDB2FCh9y
n3SHOyDEvcm0ev6/yCTws1mEfBWlGCIU2RGhHWAD3N5g7cUjQPdWrSeeEN1R9J7D
kRtIQqYb06zqFK/lNKuhBqBU3Aplp3+jjYI8GGKtIQOBOb9hOiblh/dVPWZudjSq
LtV8FYsxGcO+ltpedXfeeQJnVcVzXI1HOg2Avin+kr+pC6vpYNxQbXStT2j4CSiU
f5GeTP/mMbAWCKPuR0aidZjU+1L9qQHStsZCCTH6t34Co7m0Nv11huFcowZeHN+G
2+Szh4Dx1aiQ5wQtJEJ26jLBhJj8mjkmkiAaXrFo/WykxOyoN9vHc5h/5m/TtTzd
Ejwj0bBxwGXfg3AEj76IgH4uyCj3A64MBQPuQToydzhV2UahRavRUepfBRgXX7jN
P5JvrQio5Y7Y+t+OMTBvSG4TcDLPrAwle6ovoh3CBAjoCSU5v7WWewHIiMGEpaX2
c0MUckWklCUCvLxkeoyQ7TphlmpWhbRZFFCuATE7cgRbfOlmpM38gbmlvCawibeg
bshkGQFO1acB4b0Vwa+QVKmHUTOH/PpQ/rrhWVh0hqWd2v/5vj1wmWG+R1F4/NEr
VEntJfwSjKBLRHjQjzr6H+NSYshi9++/eMu10/x/o4Oh3HY8WptimN1LS0ldoX/e
LnIFASGjyAeFlRPVfLw7BRuq0BRW0WgkdgIQ8BYItU44eTr7F0VWBZy6dxUIiqk/
CGQVpOFUpr+FikaYd4R8Ixe/jNevHgctH166fXkPdjO3EdQ3/Fhu+zDcvEEAcN2N
+JGbZo4yeSCKjWqkdxPpx9dHvn+2YmEH5RCu+rkiq4MFsT4gm1B14DIcuBnuQPDN
FFN5KWfTVoYuiuitbjEDL8xBp9xa07NAKUYVVWZrHjZeknZS5M+dRFwTCCbdGGPC
smdvYdnlDwhzAvfyeHyuQQePbySQYGkLJcmKBaNFf0ylO5++N2b9kwXFugjdwF2y
mHsPmIPLS3tmH/CclY6IbbtvCMmH7jcJuhXw/Ulyz5bcy/gTqluORMk/rShs6fTG
hVJMhYW/5RXa+CyA3ajaPktel+CyF1Eq4gB6zcUGTCu7jsZop74mzqj5FJea7ANJ
Rk1KvNAVP2eUsw+cHFUO/GxAQf+RxlxRzIhI+TF89FLVS31sKmuBqBZcN9CTsc6Q
PwtmVV1iZj/O7XP4F5ju3vIpT1FIteeDpBNuxhZHAL7UqsycIc+7o/lUVFopXxQR
Vur5q2ZQAocGTLWpmoAv79ifhazz4szH/zAvHbfCYT6lu+EWqJsUYN2yfYrd1/5j
4tuC5c7PXxogtNTqBwL9nuKQaKA/ehiMGQAxrqw1tAr8/gKUzXAvAN5IIBoL/J2a
gGQ7+Yynw1/L4096GtpK3omxDdD3ElWTRPzvQJNSQixXX1kw1Owv5/P98ErYizFG
FSsy1yADiw1sBd2fzVzbCFjCPdHQn3Kf/QBG5W6VzhajiIR4ZLTz9XzopSdUh5F/
pBc3NHQPL3Dh9IPexO3rzEN0SxiYTzUscdircMFQKhTWdIwKbhbNRgPercKQye5M
X244QzRsVYNTcn0k4J2ejAVoolhykpnHXdJgeP8E9P4ACRi/U6p1hg1GclXTGNME
PvFYsHAuiSzcffkOFO8l/sH6Mhb6GcMd+PZl4dEbZ4CB7GGbYp/E+U9KFKezDPPR
aiIk9c3wcLCWP27ATVR/4oQYTIwCq37Qe0JytmnOfUXFEAU4KMJhxMGKi1ZjkwYz
4hbobyVTQUVWOsWb7C6ljZJa+2BWL8x6YZwdN4qjO8Dl60KT/rmBCP+dXg1/y89U
/OSciqmSgbkj8rJ1MFHnkuFNvZPK2UUnQ2Xw29DnyuC6GBGtXuP1T8MkCTKG3xlx
xyKHNDIugdlnlcoOX/Nk523ez/WmXPWJU5kCHUqo7CktPHH742iz1xqG+6tN9tpS
jzij4qRDvmUehuge23DAWt8gmKFLMpyY5rwDKqeSbHd5nJlUrX5W6rxBZMhiFDS9
cxVxRaLu5hjCiXZgJXcWF7JNyYRm1Rrmcr6UJTK1j+zVgumSNXNOEE7qN5YQsYhl
tOGQ1RsSzPaFdJl5JeLcEcElhvY3rnN9L//s+58czCFIRn/Jj+IdWkpnmefdb6SD
XYaQDmMMqy2NIkXx4sJTGw1OSijZOWwPsBCz7ew9LKIm8ObHXu8wABrZ52PbYOdQ
gypdH9yrX/u1iZltJskFCwIWRe1zZ5I7kK8PiE9MBzslU615FHvVcZAeZKNZogB1
yRlphl0zTdHKluyymjqeB0O7g9qhEI3k0VdlVkniE/5wYIXXo0LdaeC/CljocmoK
SMODjjEgkFFgFcp8vxLVTFpKBZUP+vwKVkyJOOVXUUA460fW6P2Rb4Nwz4nzsjoO
PIqk72g/9azOo5PjUanM/0QPsQIvJOafv8z5g0jSkws1GulboQY3F+1amErlKJZ0
XDOLlzNpw7/lwgCPzeXCSeYAopjMBgRp5iiHwbbiGorv/4YLbI5Dx7GDGUws6gso
BhY4eyZdBbtR98O3py8DtcwAa/L+M7+1ywt7rx+R6uxqQH2ymPjdx5Ju2PO4LW6A
1KTfujG5w+a6PAMITYSf3gufIX8A9/8fFoxfPzTGyfVI0O1pFi95fZU9igXXoJ9o
XEQWa5cVuLnr5KVZZ5G9fySbG6ME4Tunz/h2W8M08vnRo5bnl6u7a540duWNfAnr
UlMuncEt+JpMSNs1JpdQ2fXUcFgneHMNe6+g9gxAlE9H07VWssAzXKcsBxFnMmjM
xoA1HBRwI9VhG0jvNmuQx+dVoxubZ+3pzGgsQeQb1ZROQ8+/w17DGQMSMdqzeWB+
JlnWqoIsXu2Rs4GFIE7LJHKvJ0MPOZoIQ7gWyCOsaXXRsoydKzfoi4iqKRr7DWwi
s3ZBqoV65y8dWHu2X42a6Zw+YnvvdGoBO91HZxchkFHZcnGQmTTPF9im74ECgNre
ofPbRHq/cKHB8B3xVnVaaVe7O8RT0jj6bhNOqluBh+B196f+ONP4sqFu+p2MGuJd
PU2dA4B3eOFTT1YT/A15UJJe1VlYBKqTfvPhx9+8iqkZj6Z3ccFK1RH38r+MBcv4
AyVGR6/ZDXliQ3CfU/Gnqi0tPZeis4MGQZN4WhtWnsZCDswsrdhDsS9HoNI47PGO
lfKWOnRcPUdKFgUu52DrXvSN2uzpebHMQKo0rAYUG67FzLsUZJecSsV7IcnFKNEm
MUz80dboNA5CZklaSe0YpkxSZT8urrMGyK4Tke5pR26cIWcogw5j915mfxYzN3eG
p7W/7i8rMaEzsZiUVDFVDvy3FgTKZbDwipuUfSWqobHOJo6o3+vb/cQwC+zZn/Zk
dUqYkUuNgV3FRF9xh0FhLOGy+UjE2K8NR+uPpuERIeX978w9RK/Se2IO1WXz8ufU
7VzHe4Uy6JPv4cTDv5bRPSgiKr7DNDJh8wInlMpFyDcXK4RV5ef1e1I7CJX/jbTR
wlav1hRrSdkwf+G681tp3mfzjngKsruD7VJRVE3iYwg4Oj52s72KoZh9v7PL8Stp
SGHSgeLILpDRCL6Mvb7igEglotYtbwAId07zWHbUwMwviT/aOKJFsYjBA0K19TBU
kZMxWCJtz5rBpppvpNYeGBLU4JLMBbcTP0s4SYdo+3mgW7uTS/wIdZXyiMI7cfkA
TKKFgdAtmEJt54nKV9xlPFDRzyFnydBXf6gnuVnsAb6V3U3nSdU6jvIsISEOsyBQ
cFEXvnGhbQfgicRceGvfY93+XeSrdvL8YOnNBjLgyLed3ffEIcskMsj491gUwpz9
V+nAAtrRPQKoEKzraWOtfQoUFDNKlhMdT7W+cmyS44QR3Xc14YSLIXW5F901mDnV
dLm6MA2f8ZtdXSzCeVS24EQdvt7YqaEgskEaogI1J0dXaLRpYtD+x300Y41wAc62
ZfOp/LR6GNWy/sMmM+x9ss2M4Z5DgWEkTNVmhwaZPMzREDeeAuE/4q+iGt6tAIoz
P7yPMvlQE1fH3wjuqtQ0AUbznHTTTx6ZkuftIEWD8xwbOZ7DUplJtkiRAqKiKtXc
uVErJERtsju3tY1gCI+ZxlcRk1w01qREW+yTOnU9GCluhCmJwpjr7Las+2MqR5Yq
VwTfFabIoRg+TZNy9EVLTne1yTuTgvuDIKkjA/rPxpZfrYIzMlPh4JtbLGvtdUxW
qSZHnaGimHunbd5wf2ISCRpJOE4T1sNhs9vICh63wWxYIkJRuj7fcvRBZMBcJQxf
V9UMHwn/oajthaDhjKPZgDa0wz91wvDFRK1EaqZ8kj39e08S+kKgL1j83ec+PqWe
zCJPpVTa3v5fQ5Krn+RIRgAf5QmU0ViyjJ4Vf36WVbHB/YmQHiNRpFDCGlXmhWHZ
/z8il/Vix9Jw7SE0iA3pWuwo1DZk4Bw4ultdvC/5ajXn+j8qEAhC4kln2J74E9H+
87cnHrglP9UTALCfT58gJ9+UG9Kvelm+UgHssTqY2/pfvooopVg9xZTuTb0MBkRw
PhduPMlGJGSaLfFLwbUJfEVFyh0y+GaA/m44IMn5llXcYWROdeQT0AEThSLCzA/n
49zecnuSTryEi1T/TlRw8gSZ/3+uWsAV8GpFKVG9TZJ9SHp5CTBbxoh86+wf+PBV
mINUtlheycEVv9ILLfd3u7a/myuD9AcRZ4YLpm+4r0mFkOjNYgDPM24XqYhwp/3e
WDPTwOem/iRqJ4UPXHeh/O/RBZ6Yb3Dt32wv7Lu941zIKy93Fz8YT3Inzdnu91sG
VC9c0yQIRKkNwEgeW49MaE0jS3KWakuuGrFM2pWiavPZvdsynXjxle9BDDX75ZPy
2TMGAeMdiD0adn5fuO+dqKeE1rBSWjZdP5GPZJl6XLLZGuFtfhkQWhz0PPIl/2tw
849YZy8TebBcfqup4zNJPHE8rHvx7TbAxvRzwFHRiybclY5JSBOrQkJONpXUz6K+
BtZalwLQVqc4ckKa/3BcmFQGkohRBj302ExPlEXAtTIVR8ni7JQ1mPViurNrNEZI
4lTVwPxcCVas4ESa5b/CUsCrz5Sq8dE6l39gpOGcKkqZ22UkyarHGLWQ+BeKrtTm
5umpr9VhL9zYnPt0g51881il7QCUeNZsMLY6656j2RcpVhgoKt7JHnF9wInAUwze
Igm1mD4S3O6Dl/3iJ72ocE9T7DUV6cX+s3PlIURj3cA4k1CA6a0/5K96rcsvWadM
kvzP04zO1a0GYZ9GpQPNmdEt9pJ1tQb+lVxukRPLGBsmiofZgbRnkAfacaU21Wgx
AH8ECAy2CLXtGxYxDohzZjT4CuVo8p4seOcQ2Dr+Lz7UiwLPOh8u1yxb8+ejgYd6
NIEOdPxFgkAS55/fO1cWdXlnxbe6tu17NtZWWE50twRm6DyP+UGYHAHvcdQA75S4
qEfQYmWwpMpktYdEE/6WMEP3UZ48x107qdUEHS9s4M3CIWZlSywx88jET5TTg8PU
qvZCgGY2DPFTTB8J525WTuowG6m8BTpe3uW/ia7fiF/xDxhgYzjKRWBkqTAUN+1d
yY/IfiKpQx8No3HLyc434Pnn/F8SfuZFhuiNmZw1mPR3KxH1eunGUgtvPfFhHf8U
5/1vo9Rbw7yx7q+kmwV2CGXxll2ucBw7o8B2ca92vFkZYsTu9X6WBrroHpoxE2Yv
uPaS1tX4nBC2RkMqYKkmfymU4MwSikKKD+UEKTzU74Hbd1Np97LdSdb9scrTznFk
G4ovH/tp0gTezkqTiSgz055r4flGJHMl9xIEMY4+qwgdG+TjHB+Mg3tFEyklv/th
22u0Hx+h2r813HANLMW9xjxsYrKRAgpc6G1CgaCgupfstBQY3rynAUABha1wJbOI
A8LMIfscHTu9IbUOhY/WDdT2eq7+E5t2YmNIuc735aZE7RERLR3LQkwRheDrkWhn
od1I3YKAi95EKdvFLq9XEuTDpGFs+xrM6k5Pj5JKSiHu9A/iyHfWcHN7lbNq9Wej
ZQFwwplWC6Bet8frVsndN8Nim6FRUVwyHrjL3lgWQppqhFpkxzPV6cYi9145lOrX
FRfAN58a7XYQkF6mFqs5Hkdr+unN8ZsphLwluH49sAgLdanZoGITAtJDSDE4k+Zb
A111+0RD3OkjLhOnHGGu2hOtqqXBzXGyxj5b9M/W0XN9fVD9ySDyBM2Vq0o1c5XV
LwIhaCVZY4HgRCezDuLshVSdN0ZeoDI5mBRe0IC015oeA3J2LDJ7HCPBofmdh2YD
zsAQRod2Kgiab/FioVceQaEWKQdRjUJ8ntbHA6+L5JLUT7GunJO5XXTqUM5k9Pp6
E+AEUXP33hTij52JDIiYBmt0Ts807SoE2f4ohKA0mN4eZRtkpvKLZbxCwfjmxLet
EBJtuM4duDRaSZyW/S43/3HaZos5/DjUwKYOjJCb11ibidMc5z3TSJMIsoLQv1Us
I0oqHlLT3AAgbBRx9VajYHb0XfXDj1qbgS4H25oTOSolIKMPQyn1ukyjsYALjv2P
MkBmwZL9nDJARbQJUcFyW4m2K5gVpqTJvSmIwl48YyHsrKWQfGsjcw6JxODEcIXD
DExGJwxhPwQWG4mgd/x1npLn3xz3m80e0w2SJqkcKa9XJrGNp/rpeiS539WIoQOd
GAc1HI81ZrSQWQ2g5F5nxVPExttdHNDIPS3M5RdfrGUnsv06T9i6wL+9+wgRix0G
EU4gWe5Cg2uaEg/k8OI/518iSNv1ifh59AeS4UJ3zbf8D1VX3RstteAx7nF0Minh
IQ7TF19W2L1LludBcT+MhZDrv/Xb+eiRIKVqmRt76+PZHyouahG9nIgUv5W4Q5N4
6W/GZsJ5QNI4+xqyQ8C2ktJPkWxD6YP3wwtAwWG4fLqVwmPD2jSyGwtT96zzTcgb
RZQuL5grTClLKjj7vmkL6ynkZOiDFK1qe2NfqK66edrt6zVdN1HJFdeeYABoBH1n
UpUZaMGVfcoxSiQqgW5bAsZSIF8aVYyQSD2uTDDZqS/DhS9Zz9LOgNXKc2qAPrrs
ugtxuhXSyUF3nZOfogxBfhuRAmOBjUAOc5PvR3XEa6AR0CkQY0RFXdz9N5F8fvWn
0CiMlcudd2eVex9Ap8TtZk7yxiHrUtcO1pArE+edtEGcyqM2yYn23Y+3dbT/4KyZ
YK4wwLE8t/EDpXNVf4bL30mn7nPXVkRug3WJpn4T2J1ZLA3A5BxbEMIwPOPfQJHx
V1u/MHcTzngU4BmvpFZDea/Me4uan4mgBlGbYiRdu2r6NTqXpSlq5UjMcqtNqZNm
CXeb5SjW+4m0Ye8KAAOL2NPD6qsn/nh0MieoOT0nd9lakuefqqXwAVb4AjPaV61Q
FPVKM9rrMur8QF9lHn4zw+xkWGJ3F7YjnwG8RwiPW1wzDg/YmURhTJ2kpLo64BTK
E/lxbloynNIza0NQQRqz7hqVteTlJ6JJsrLu84n1umuS4BFJe8QrdhLJ9UtaEnTv
SNyZg64o6wGJXurSL9DFeCRmx/7lniSU0VumYHW8BWQRsbRV4SrNolCXyGZCB9z/
Eia5vTNpq11qBAn2v3lXNXn3WXpPcg2ShuLEFKxS3khFIeQg8omR8AdJwHdVUP4u
CnhFZLLe0JRh8WD1h+8IsIanJ+ziHhUjQC99oTfPYLh4HCAcOJYCywTGUj4aRtYc
NEhsUum9Sd42jDDRm6AuxXm8Oxa2NqzJquPJlHu4EQ2o0NQffw9yHF3gDBso1PaR
OacLrstiWJW2k2u9//vGF0v+R0tMSmeuyH7OThsjEgOn//LrZiJWm9HJX55/Db40
drd7I2VIPXsVWglAqB9v9ZomJVQeUW4Jw4KulyT21/zb+0aiQ4XvYdNAFWP2+Lrm
Lpmo0UqvfDgI/ZHdxP+8hkQI+RexqXSttjVX5Cm2e60OvJJEP+zmsKprJLTZQ9mD
uYa70vRiEQpGGRr/D1n6uxD7xLoga8E3Zi7NfzgNC3vk+imVMBym4w42thkXfC0h
96CnKevBTX1ECIjYBt5qmn5vuey2wilZJq5KWG30jXjaoYmIv7HzyijCwYFtkOva
ui/lzYwQyh/D4VmEg938LefwiprEA/baqwrLi8m009Ch3npJ+kQxu4CNjioUS1Hw
2jdAv5o8ZTSxjau1i5swZsUxCyI89mG7/qZsatGyTZXsEkHRzNZMYu90++nRXSYy
T7dF9jqFHAlhietdKa88u8d981HkZ3ZQOz67SwTzjIFoGmS2dQ7F7+DulUjSQLKk
LkJv2HQD72JrmgMFysvhkbdk2+wNKYQsTse4MLccdxWK5p7IiIoAGjjAguu/RYRi
Bjgvkt8BpOm3A57WoD+5ajIG+CkwUDdc0oLAXmfCsCNXUssd7ZBGvrTdw1o1Q9Mn
pT9nYFRgX0NeiulubJkWEIb2j+tP1eXenKTqUViq+JyMgpekaAkatA5E46q7T6jN
fpPnYH5cuLt9mXurWl9GKqXlprbp8HfmNNab2Bzfd6aIxSejuWgKnAASgr1PmsKs
n4tjxRjGd+yx6mVgtjQLQiqAHBaIsHG0CHIymPJc3Ndir15bkSL9QpuTl8G+DaZq
6n2w10fZgapJ1hYWMP5h2rEKqc0AXLwRzNuSxYxb9/pahCR353V+Kx61i+Sw67Cd
u0mJpwdne6sDwZw3ygOVRce+dZqx0hgzRawjMxawnjZe5ZfzFykhlCdceb6V5/5Q
DttzzSXpmyosuY/lVPSZWk3MCxJ8tMNOBICHXKjp4+lKo5gi8syHVw+l7D27Mo43
zXVuh1R1hDBcs6cJjmUwY8OX3zE9JhE3gOmAG9tsjN0oKM/P2hXBSJGB+CD1jKxo
aWxwGAS7+jF1USPYQfOMG21ZpopL011qLHbuanB9zkOcojfGPOJ0A4EQsQ/+NWzJ
Lx/aLLuI6OIo7Y950MHqOSpPyP5gtwARQAAKiQkr0l0RodyIqlObE2sjlfP3a6T7
R1A34VPomVY+dwAYci3fMHGAFDNTfixl84MA6NrvtXSxstOYPxSZIuC1arALCkUZ
IvBGZ65A9xv/uHPNPvpYY+fCBnpcomoyCIy8GfKaL6+nKdhGFMJyxcFiT/z/9lX1
2TwuL8edvcD6aHjAnEYL8QrsZdkapZdz0oY8UGiZEljte6Wkbso0nWaiJn/k1pnh
F2TH+g+cKri4sUmsziCyLsA9p8lLyOY/FMW5NgKVtBbeDyAKX5anes8udIpAbJ2z
QCmxDXGW/SuISq0CVjHmtEwR6I5XpHyCi+Sv1aTpD4CtlAFGYjWKd7qfQ1IzLqpr
HhkYk6/XFKqK/9DB3cDI2woLnhdTdScNU8PNDl4paK9mS8cjnTdPv9bP3SFwzgXy
Prpu03DJUBQwVR5TaNV8TEH3x4FW0M+O8AWLujvYuxjtse/CK3emjY2dH3JxOSv/
Gv8w3OaSe9/ai4WPT50IHewM14K0O/84KRRpkzTGP4SsOkDzVuyWiTKbliu7+VgI
KdqT/tKKZC2T0XJXSyhYD6abF0dDh+6C6LOH0RbH6o4rDhn/a5xYl+BmW0GI+RW6
jCTsQ0IWiSgqklrmW3pgYBBk27MEeziNcwymiceY/ffICuog6KMfAP4Dsdy68+7L
Yv5q9i+kxStDSRjeyywMVFxeorl05NaP+djZl9WQMBBdJZ5CLVbodx8gq546dyKm
eZ41PVpUZygA+Kvr/Qo3rh8JhB6UFvmMs+aac64dlUM556jeR7q10xOGquPDCmxl
HcI4fYn7bBSVIh58qiAfNuteZ6ZUuJqDOwN56zQk8Q9AfD+4mztiNJu0fGpXxqeq
55lIkXfFzrMGfklA5msaCRUKMMkdw5RptQ1B9XHm6YOKQ80nVndbdYtsNX5ncGcN
5d3MZfve/Sd8jSJH4cDX3U+w/lV8bgyiBGnradTgHt3eKZO2C3Pe6ds1feBm6wZF
j0C30qaYckYQYNIvzLAxOwAMdPb57djgZfabAM8ICGxGOtylUZATwEWft7SOorS3
N4l6WEAU9i/kAm5LTg28cmvGaOl/NPE1hZvVGyu/YIWBJgADnHDFtIP5nRZMfGAD
YNvt91TIbsdWJsxnZVjIEK5CZ8kHDZfaZMoogiAWqnQu+aIysU8Wuc6ynG8ZRm0B
6JdNoKQlCxAWseU5xj5P4JZNSo4WQsr4CUHp1IA30K5FJ3ghwQFtrNW7gg/ykeD/
f/lriab6vbsNkkKCdBnRpyAKAYrtUpID5gINu4A2Sv4IwDMAPxy2jCWmvG2Fb567
UIM6tTd05++n6/gkDwQrWlnUy5RZf5RI1EGAIoqU5EbjJ5TYvP2z6sL+4PL5EcBs
v9sg1EUI82dvf2WxckASP5cWhFh1zrLFV6M0ZaAKvqvxsbBUUYTvOhKN2CDAMsjc
+O4/yCR6Fjur1nz0xdUHBy+yZGucVLm1WQhU1ClhA+znIk5/Ho/F3VvNMZkBzrW0
2C1nVFVxs2j0PLBR2hvCvPPpESQtQM5Ou92aRcyJAVh37AFBSvT5EeeivxDLqN8i
A/YmQXJ5yMLMdhRSyhYZp55PoCx4ygtsKU1Hs7Gcsz4AS+x5sxSRBwZk3gCG/ROq
ZCgOSIq58EPD8/2S/pk3u8pxOSqrTbrLOrUcmpqStPZqHwGqEQBPjCINrF6Knt0r
eRxjh2Z8dPyFX5B13mDIwGp/xn/hoi5NmVwKTF2XWlVJ/eZJuT+tqBlIHlldAVEn
jFDYXeKGZZD7k3yLYs4VTwMqnIBadUoU8wvU+t4kgJ7LKF2naq59pDU25AprRT4i
YNUH2wQlY20YKgjFYPhgCDu1NnwMbEkOHe8i7GtmpVwtf3oAxI5KxHpJSWGHlW0k
n92DxmcnT/OHIqG9jAMz6R/q5Ze+AxN2MSb5OQnPP2NigxEpS/47hknvGynnD+kp
kJQblUGYNZgYbvpYF8cgHAbkKZfqZpSQrzKkZtdl5Vs0QawYNYoriEe6+yLPjVdS
IZDZfS3I+u/20WohMC0ox0A4nGLQbq1BKQjGFGjnyRPbPiRgWyABIx3kYpF3/tuT
uptDJQhuPqzNBzPeyxNwBaH/d33lPZ9E9J45w40QTUnXpUc2fkyGrmDm6KeKlDnO
np4295j2ZqHL9bpl7mOrtDd1Nr3APpsd7bR1D1V9bzELe+pYZv5QZzqTm//4DYAt
x6wa8tPh6eNTnK8nMhtZispTwCJPGHC4E8QIZTLxgJsMf6knpLVlDms0Ggig/65I
cykla6reg5AvLGhd8AEeHMWXEMDDJLZaqh3+rqQOLwCaD+b9muy8GMB8q6cxydDr
kgbN6egssD27hYwgxBUb0BrTTbUeqrM23YgOqymIbxR7CxhdRRuRj1NqLghnwFcm
9k9SQY4FHupLZk3NrUCxiOuBzd2U3t53oOMdIEPcT3W9ho4cj0UPXK8t685vEGCe
jm3Yi4SSOEPqffexufOMfaYBGPKGT53muOaOnEcZzR4w+a/TyJTanoL+swmzCafy
9p/ZwgP4zWqGuUBfO1TifFd+bwEnaS5nKmeCFlyewyet+dxNnp8X6N0DPUOxDJ+z
YHnFMhjkUccHIV/Mof0mhlDVayxwtABLRyoLeJmUcsgWhOMGpr1jdJg5Wvs0NPC9
ZkqBQbjm28YhbZisy46vaXl5G+Zp6tS+QEO40DPesYJCR6+NRsHytGQS2eTmV7Oh
FuDaVr7VLqnzueT+Eh52gQm4PggH0C60o0Zj0b91f4lX8Y0UF+1tAwZiXlNJjZE4
ObHn5/Zq5MIpmlbe0gX0H3aZL0OvxmXQolK4mLysHfHf5srNYk5Vuqz6g27Gm+6o
BBapcuXYxVh9Tunl9/6RYo9dP2xuaEaCJomGuiWeRH4LHdwVQ2bz+EhgR7fIm/V3
p3cXOiMy5DhE88zrKK0zj7uGoo8HkEkexaC2g850TXk0aFKh3QGcGj9ysqmPgiFY
qoiAFHbzOhI4UldwD839Rq7biCmDihqKSoTT0FZkciBmCoEa0GyFWqZwn1G0EHPF
R5xg+BIGfyBFSySIC7heA0myAqYMpH6Le/uNUq/5MNL3Wb5aniredd5YToD0v/6j
qOMAC4HCe2kNib+kbuQAyCHM95TIbT1RGJ08dJtyIkb5coqMjIsQ0DN4ylBTFk/e
pc0sA+12YsBqkjLlAsW7hjdatGVPqKRUKjfgaXZMHLjaduN03Omh+zsARjT6uHzN
+X4HQqT4X/Y3H7oXz2Iw53LJtYQsKWra9tFx1xa0Mfmuzy3vYm5/Gu0lZn7anedc
ZwSzRUglobV9sRINAZ/YAytFshl05u5yKgZcJHB74aXWaoKabEutt/KoA8upA2hI
xNOSbpob1G50TE6LQDE0D48oCQVWJmAzkLhy+TAMPv3dINHAWlhub3pc4WpZI+g8
gzFYC5UZmqcKN+slIjQaY4ez9fLjTiKLrfyQICiZ+o9CBgVZSIBtRhjpqo9uYYKM
XhdYmsdJYuZ+JqoBTABdgfIGoc7zZFGSyyx0O9zEy5qswinttXegSsA2FgbDkbtr
RW2aC9bl7Mgep1NmicyG07ERXRnW7fwlG2edE7VnJZu/m6L0S9+lo60ZiVVgFz3f
MbWfKUpd/HrnpQABTcVUVH+S/pBmtzk1cMqzpg4DdphUei6Bd7E+Bgcr56N9HB7M
SMSan5/h6jGRPs4a9AR3wXNAwvV3v45X5N1UAFQuUGAta/r/E9Fg1vZ6Jgmhtxs3
fs4iCf0s9Uaet+2WHUUwD8fHy6wTavS+ll6KthWuIWC812DxoUbU/Ulo/aSP3KQu
ZL+ZDkUH8DfucWucWjOCVCSUgGbSxnHwpVa3olCOQSb6hEwJ9Jjy/CgNb4P8WJVv
lhqaycLnGkR3l+qxF6Y+RL+ym8l4O4dYrE3XkluT5ZxOaMAobG/YAIxcGI8qg+4Z
foLgaA8defO5odnZUs6oQUs1estPRs1BcWl8eNSF0yBQI71++ZnXHCT4KDGdwYJ4
dl1tsgRa/KpUkfqr0tPsI2mQYd3M2r7TnTAGuooWob5azoNvosmeDNveZqUVKbPQ
/5Sr+oVJK0nqLVc9D1AI39j0M78r/WGnoTyq1lMuROXQ4rg/EurVaY1L3nC3HwUq
DEMiQhku9Q4fjb69bLzKj0rr8POSgc2M5Vk5ncoisWETzysqoS81AUD0tG2V9+9O
5FXlJc/xFNcxABq8kysGJfJ70XKODRy1Wt54p2bLurx5tgomoSBG1t9ENJNk8AUh
fyXmhF12G/6XddOwcEBoc49iTnKrcSRUfmyK7xTQUoqj0mBq7uf8NhO9HgUxrKfk
uEAYWO8f7nr06TMuSSu6v1QpCIV9Mk34oRAxPYwlt6mTgdM6apKD4LPJ0buwfwo9
woq6OaKvC5GbFxpjh1MV7xxULau7+w8/DfUmP1ZyUC5UQa+9wrO8kgs3TGUQ+ZBl
J6ueEHWWoSTeVnsNbl2t6bgDKAPtOkI8vNyvexLxOCO8XSewUE2BwY9GkriqEzE8
YjGG6cxLOIvQLBoGLCS+OHPZcMa2UzbHkqxVJ3xVikuBcMYzFbv4BGTEHlPPB3Ug
uuoVrdyFX4UikoxJU0vr8TaZ68GpkpSlGybhIVVOP11nUnI3o2QWX60H/JhUWm3j
8ONdAUT02VIwyuhD6vRRhyOz1kjbD++1c9CJ0tH+UftrSk0fEJJMTzucoymrnKf8
Ya7696XxG7WuM1e7n22fUwxhvTW+b145RhplG76I4Q0VIZsXJL2qQmphJiGeomcj
PzUbxfdbOKPfNdaUNDFWhyITh8l/sPGayS2eQ82l0U3xc+3WyeEzc7QFc76qpF4E
wYjxBwBqGge5IcLz2+AnMpN/rON2YwDYbS2CY16T93Ntf7FlkQdIpMhzJXQ1ROqD
xsLUUrxFE+z4iTxOi7n78iUG3DfwiLlTsuRMnvBHTQZ9hH2tGxFT+h1xdXb85qEX
SFqK8BjM9LAp9nwd9v8hCxHGrSpS4VOPNECbIxNvFs42Ynn3cT57TGQ/5amybgtc
AlJKLbO1U+S5htEOMfOAHaJcqYY1qT/YyiqLewr7/CYHArtXPSVOFcaIyISZkiyv
fjMmqkhE2fCi0nq4Mw5PxoJ6RmeZdMxyfPlQit7MnBlZ/OxFJ3UcoY4NufqHmbaK
0PaHDYCx//O594Srf7bF39wpzBwV2YC3AVZDKpvYZDDuX4ZL5C5K+MCfU0XacHT6
qOCRyIYKh2GHGZIFvZ/l6lLyugBi0yCdx1brGzTN8q0Gdf6P9nsLR8m1MBURkjG9
HHpCdT9Dfws+dWQKmfRpXiRp0rV7oV/s6LeR/DNvDkIn1090X+lgS6pF1VlzErIb
4NXIdDPN/v6Xpowp4XHm6gbg+QutJ1cpEfViFbWTkIHkIetaLesXy7ybZae9URXv
p1cvxp3eQ6LsPaKfAxnMrJtBxkV5xhb9cbDtOzQ1EVQ7ZHcGPEo8B2CHylHdAdnj
UgAZHWbKGuQhrAljuCAA3sPXbY+H7QC0Da+n+Ep8QaWicEZuyjS9zSQhukQxaeqh
zEUy94PhZfqx79I9Cam9pC9+zPt8Hz89amY08BnwcoxY7AYEgr0j8Kma/rQXoMpl
S5abTJlYFlJosYkkNDPuZQLp8QLTQnK6KnKwPC8r79hoBaqmrmCf/O4C6OxpZ+3l
2DlPb5eGm4hyiMdatWZ06QArz+txMXJw3xD/PXNIgPTlD++tK1+s0PnryMiqh7hO
cV+9FTsON9Vt/pnKjcljnnf1WnD0adbpXr7At756iySQDck/iL5fJAQQj8YoprZp
5gg9zbCAzP7gLJm1gXVCwg0/dxuGM+px+uFg7FdIzWy8jMgYKBtshjJYoGHtkBdg
Wh9IuNLuL42dXqG1o2XZE26NfhiK+pd32tGtpa2iBatoDsh7HBd4/S8i+C0pWl7n
Rv167kbNEkmrzCL7TEsY+VHi8zJ4TrpgtwuOITexXwaX33xl1xd9CIS1l53ZII4S
13a/h4T6zDisMM0OYHLOpY5gin2ODnxHvVVg3K5OM053i2izSuHqnyaA7ho4TORZ
JJre7r4JUPe2IpbXGRfk4g+xlus4gtJKYqPIDYe2i55tLP11pLQ1Y0TQHNQSK77t
V4Kdzh6d/bKitwU5VOL25VRp/x/1bRcaWyt7roxK1Jr4UOBLIuC5tdFSdHWC5DoX
yE3PBG58gy6T4X9i6bt3STAe+j8iBoLofgI5Y7mRrhCYB8L8vdCptjnEvZEqeVHt
4rilPcvL5pPyHv2rZoFerdQhynLpTOwJODooxz3NrHu+3aHMiG7IZQVpHXL42ZLq
xTg2Le1BKrQX/91VkLREz9HhntvCKf/vlKL8MjgG/C/OXC/4geia19cYKE1mj0SU
fIbjuVY73SESoygzWpYb13V0QTi/pNE8Mt5FgV/iGpEUfriFaEIN8dLcIzeJT7Vg
KHbKChYLVjAvBEKEbWdT8jBfXYQWOLtgy0kcaYvuLt7/OIiPjo/uLEhlteVXLle0
uJw0FWRDp2rb8Q3y8h5gsU4VMtEUFnT8soquFpgnDLKkdJcVXDuqlyCenmfsgxL1
dCoB3adnj9wifR4TqVxwCw9dS/tRKsQUxSk8eC8drbI5wsxgi8p3PbQVu6SwXQWt
yxLmZIwr2s7V8PHVM1zJqwPf4j++4ZPa/+P9SzA7CpZwzvCi/3UvpxfjzemEFbJI
T/MY/X2dvdBPF0c77ho9MkGwbNUCmIb8e/8rsOQnpXwg/VqQqunCcYhHHjGD68YK
2oa43PkJO498UZ/0KvT/9v2yyB8dCiBz9xwABK2dTVhhcl1svw2rDmucpLUm3UT+
TNzotxATJm7By4zBpVApYYq5ZLxsQkbnVx+9FK6s78BQL19deh/HkgCh0y7M6KjH
xdDtdf53ij8WsZJQOtfO6oWiCsWIKby0Pm7qQ7+UPyXcjJFwdq0xfjjX6iVPuvzi
HNyiKAS5+YecvskxyGGN6NBn4eOFzawTaV6h0XT4eLtelZU5MKgcIO4XJu2wOuDi
eV/hzLsECZv4Xpq8zJdXbW+RqEj8iWTusLKTsqSK+xjZ5CWZqGvZ9igjxo6n0ulg
7hOqwWoM6yz0yXXhv+6m59s5obMyQfspDsDqg1X8rEjrs3HVTYmVt1V+QTkdMY/m
R9FLrMorF9OXFSt2OsXcSRlqzkVCHEOYTAws6fAo9kMRWPlMEPslJEet9Z2hIpcw
1ELWBB0sWBdM2WBIG5GALU9OrCOM8ybbGXukQdTvkC7Gx/adPWcW4Tn8BD0+Wn2U
b/sXWBoWCr44BbD5x536X2qVpmACzfyjmCkbOrpDUV8gpQgkFlx2aTtdzZSfqrhH
o2xpjPbl+tlKA71zG6FjB9Of/meH+DuFq8hMacC5iiVjMiC7EXgiVkZBW38fJpI7
2MQ7ZPAva5rIbxmCoKR/GDz4Yj/tu7c8uX6fYypCoAxvzjtOPFx+mOspsRhemNld
x8oO+euwUQii8wBa84xXkjbaUER7cB+JZMvMnDg9BmoBLRqL7v7m+JJ6k176+tJ+
IUFZdrozTX5iRd/p3+0jmMf0VpK1Hs3gDLV4zwQ9uHLEC9kbAQm/QMhrYTUxx0HJ
N4u0cZsuyVB5qj/kOADnqzvrUmglsebCwJDgIBt0dtNJYHctW66MG2YRbOGWpWzr
VjaE/wSrH76Quu6e9E55vb43xjSFhta763EPks6HVLJJgxJWFD/0F39JhiK2xqGu
yL4tlw9ujz6CRGg24Ecuf1Xt4zA2zRsOOuPEfddy8CIKSKgsBZl+kM+/Hx9S0/a8
qQ8q7wL5Fn45Acx19aBY/zjAB/1HrOvnq+hDm5LaedBx1fjgWLg6oio9JllAM5+m
OVvYLAUPLlAhmvhE6p15bsO8/HGbxX4GBetY6SFe72u29kHUSiqoNS49dTRWLou6
goTWihFTnY3irRUXo+K1Vf1YlynRAywto2dNt4mg49D8LN9SXY4RKRu1oY5IYCl+
recXd2cPJA8L5ulgpX2M+wv2FfTwfcoGVsz0WHO5D4S0LdPyKfGinzeE0wfLSW+7
OKa9eyLLL9m59p2JuL4+fpP5K1D1eN5Z6YzNqASHAHvwgMk2eMT6Y/EGp0Fo/5wh
ORdX+X6KkIyUjTl6p+fUN4DQOd/z02ri0tk+Rxig+BTtZt+r7k3qQ80zRfd8YxoV
ozvC7jRC1yNTEMN/JXKSGMfAMvk1MIsh1ggy9ETLAoi4rrN5IGaGUAjdtZ73oKEZ
5V1qaMLOuDyZTlvGAPRCXdBh1FPE1SVLV+hEU2JZ/I1dY4KuschJ9HqfNWkNyFcT
HqKd/6FyaKf0tLgxaKEsWPxJ8ARhn8rdHRB5tHXdOjpsG+mLdVqptd1s/2ILgCJD
VxNToYhfLISjqDEHYMFYmbq/ZQPsaGi0aQV4f2DDcyyPMzpErh2Tpi9lHJxF2a31
ZlB/TR+kZll1bDxMwd7c+jAZP3ZuGR+bhmzbIgN9fGmrcGWHYRW+3+sdLCmwWnpu
x/1ppiT8fWwRF9gHaPkO41DwrbId7ussoBcb2ftAvGKIKkhLT7ltGdmUGb40DZ5P
YQ/Umv2bZ2VYqQltVdwGSGluD6HKcZ5doTP0Ldp/Fxw83lES7z5WYWD9FnRl8sgJ
hP8lfpoyS9JXmoMx05KmFxBWlAwt4xArWJ88zsoxe9ZBy1O+1gduFCcURD7pKe3X
4y8oO6CellwIm9l9yyBgLTfwFB8wq/NMnzVICa8kCQNtC0qPEzZf0eXp/SbhfJXR
cVU2oAUdDJLMXc6OMGV2c8uoju0+fAoaREQBk0f8lm0u50GK+pEmvTnIn8F9NOP/
DYgOGWSadc9OokCDRuIZAcCxz9D+PkUUsLayw7DpBFY+AWuzjDXaOt//mEv9XP34
zOXcmqe4PxBUOJUlIuE2wIpEnGx2RNtnRXje8MGDFDp1XkU8riwtCFuZTg9KUxoN
T6goD5dKHDJ5sN+UBVW2SduY/lnv+yV0RX4ro5+t5myMtfcyjNjbnjDpWhww12jW
M9MoDOYCS4uAmhXp/vLB9mhPLodebh+Xlmj7BGGCGF8wj+EOoK73E3YsFS4ulqUX
EKH/xbTdIZWA1Vh3MOUD3zT60OZEGgFlsVvN7zsxC/NqR8oWJ86tDVORiwwYBtbg
jaNxE/d502MXQnF7Rtrb1KPR4koI0iJExxT6bl+qF/GHh5w+w1hsrgrT2xf/Mnib
EBIubDzPx9CTcBnutQYqUbXIPyfxlov++PakFXul/i/dQ9pdq9BFgVuCbK0RWa3F
wC+XYYVKhMQJx1ypWAtbj4fSViT5Lv0AHTN9G45d0I4f+KT8oTsc2Ks1JJSdzVBV
LXysgXXa2w8MkGEpdc+24av0t7R6SA1Ryq/rPhWSA2uNS22E4POchEDOmoofE6Xk
+LMLewHgvXsjgsjrmxdGykYb7+S/pyWtM/phWwdAtxazwfA8WstlNrlCIQATk7lS
V+2HOXOKlBqCHNzMH4xrNAtnH+MNelEtPFoIHh4iW+Ys7X+zkzqiKtS1e1curY0n
7Hzmo0UV4jtYnOaZVvTLQSYhozFOxNkkB3WAAk5oH37nuvCAWYYEtU42Oa/hXGJo
yH7tzCsRl87QoJAtHrpo7tqenXsNv6251QS+liVZiNvy0lJvMd2IRQOGj6nEL+9C
VzTgXP5mJFuU3lIJlScPgfNTA7RVd+KgCQ14Kg7QalJQagdDP67RfLPzUf8r5I5A
U9pJbFOhXQNfIpvLDQX3vH947XHiglOODqMb+RG2aqq55YGI2uyI8Y7mUMrIOI9t
991PyvTDBe4YS+vlcLwo7rElKgiJFgPeuzkJP6jutaZSd9xuLG6fDWWsAt5lr1I1
kN+zNAQRRg4qCNPK7cJRXE5mlJLwRkiwqLPOXzYS5pBg/y17n7/mmfOli0K8lJzF
z3S47Bj+Yq+zqOw24eg1NJhzNlL4GnQ0DKNoFm1QJZeXG4VP5v7EzdDh0KNCsj/n
sAu4WW4JmozoWiENOuzYMcT6KaA/1Ga4vqu2bWXYW7q9ETfuNWCRGI6SqGgfPAOw
aFJ2prF6M6d2NXA8K5bA9eYhPWXQF5n8Eic5gUXDBMUHWK+6hZxlKiZ73bywfyyd
n43qCbB/KNJzjCCRo+32EmuFt5Sv+6KQfEisSrFHeJFqQiQopT+3Nrag3FXo11Nq
9jgKYbzwGudCA8CcYu796vE6yTqRIF543zffDcM/LzRih2POu3l4d/V8VjAykVV/
67RHvOFDOD+aDLFj7djmefnxuO1NlxmNOAsGwwoG46Ou1VRa4AnbMTQV6ggnDO4q
WtLP4GxIcmd1E+4Ij4jek4jGCtWmGClPAdc6u7nIoKnTbdh3U5WNs/IpqkaQaxLJ
VOnkKdFa5uKWak5ppIES3fey7W7m06ktBB+E4hBdRb7XBXr+EBGScgLnO54lGELn
gincx3inO60TEoGjTVUlF9kugAycoKG5F9dHnQ2FnEbx2QE2EZ9XNPilw+9IE5No
MX8h//nzayYeg3PFUetnPeQ+WhnFOQnypnaaPoyM8oR1shlM+McTatpdB77BK5oj
rK+FnsxoxWx/wqmqb66T4Sj2mPD59E9z1FiyLCxfHnoI0x3CwNThFdhnbNf68MFK
AiiRdyRW1FTwnGpN6qekPXjuATLoX9yN1/2lwkhFBgIROieC4g+bDWZ5whFdYhqK
Z8es1QVYjdvClve1WADOl8qT6YztRAC0QVDMwfdlI3q0BzTikgs0e+AGep1TQJ1G
qpJK/uwf8ZKplsIUWXjdA6LpjHTCWoufQ/MhHDj/ycgZWVhaoZ8Sx/m0ZZ/2t/t9
Z4qQfS6WN6lUXVB03pOUooxLq9J1ag3Pvdz0/+L0Sg1S05R5mrHpwrVA1ezAHVcP
VzhJM1ZhtKt2MFdGPPfk4sXXotLGLhZplTFjzeifjL5jDor0Kc0/R4HZj9hjXqYl
NF/Sijxhhfp/L4a2zwvx3vx+2oKSItbW9dG36dJsUerEIWmKGnpY3wIPPK4wbGks
CKmnxgnwdZ3SRijE03MaiMRgZigDaxMUIM+7NwI2ikxfpUmBKUGHyK4Mz0Unu+0p
F99Xk+Nbz/RXHFUkthBAHR4F2EbulQI+xIsM6dfHSabRlpWikBEtG9LPH2mTwaSx
MSSe6rgATTmt+aG9yVrv/55+5Q6ncBFjaH3H5JRj9ax6HL2nVi2JoAW2Wy1ZGeWA
z6Wx8x9l/TrAsASegyarrHmncxPFeAH3uBkyC9//4fwAL/9eZRkg1e3r0xULq2ti
44JjdRIAy145EyXwVyelwqbQGu0njnZ/n6IOwQGkgxFF61iG5z3PAux1FjxSwq3r
pU7/keBykSSrrYvlovGLMnEdPuP1xfGktxKc2yjMxFtcrTMGfylhO5ss7nXVrz92
igyxU9lsrKi+004u7p0OBOEjBz7fVYI8hQ+UmTb2M6Mjm7rs040YQEtP33/22sXU
oU9wJAMqJ4vMJxuq7gPq1iDwOcWiOMVA5gwmSHBDK+3B9uS1pTxw9MXEpCr72PJO
Mcz2JtsHWBaAWGvTV8icAX/QMjs9IsBqlrqr8KXzBZizMIZDwyvmy//ua8XBfVHx
1bIAHrALxcqbtHqM46kQMRAX+4A3U7ECEJvXbOAOjg/g4B6hEOeXC0Lj8VwXEnp4
T0Tb2Iax6zdSxQwc7IAANoi/kwdPBSOqGl8CyMif9Ia9pCcp7RfpsUzVfRHLLXNJ
YxoixIwWPU7cDHcAMEYUZml5afJcX20B4oCW54uPZLaAnMKcTPsprwniMGlgSplJ
2lIvvF49vjXfAS6cVEFiA7px4RjVTwr6UEBnk9C+7iDxZKc+Lw2XNe9OrApZp5eg
yxRkbxAZTFtTcmrFvGK/dujPWPyIfiDtNRXdGncjPYS9BpYnvSgp299tEr478K6G
lB2C2+OikHQ4ebSpGY+e6XzAdZ5nd3s4EWpjd5EpRZYC4rCaFv+qAWh60VcY2+ev
JobQRY7SRPA8pEs4uW0vlOH/4W1pDejeUQMTHscYoS7jSwoCDDj8vbLlmHh6FlsW
MhFBcfW6YjSr/l+fHgTcbvAeCgoEpAIQ3K85I40i7uFsrf2pk2HjXwJKB4uQpYEC
Hq9NiHw4Gz4JkZ3rxR3Cj2ngokE1EAIjE2VruHOXxykoCjHBEf17tI2KJSAY97rf
qeg0SHQP3Lf3UR4X7zmKuWnMfC47Oy6y5XGGLS9KFgubM6HFca0AWpxyCrf2F8BK
rU3/SpHlMTex7xf6CxNEKlyMKHQ/r9vNTVdAJ0xcZih0xDhEXNtVFhZwo2C3qoND
35bL5CVqu9zz5IIoTteUzN4bRVTDSHzyFciWWyAfY9l9aIP6sy6A7FUnSwp4gIuY
kT1nxVSeIwg7OJNrbcEgGka8FrfS25MGVBzAyayQ0NkTvdSyyZemTXv3n97FZoee
Y5560ZEaIrnxpjw84jAyQM//usNUt73gf/iM/uUd+nKkrTOIaNXkY55/gAspWQLN
GtJ/7LhgHMmjtk/qVJ+EmoywpV1JBq0cb6W9T9p71KnG94kaVCg3oVWcYsRmg/x0
JX6TFXBHzeYzkKLE1saGkDMfsQ9tzOhGoPfE9aagW8dK/fGG/jifEPGx4RuwuC5m
4Xi7hmkizAPWIciwu+yA1C6ntONCkD+CT9v9LXdYYxzWRpSG0bHxsAoR92gfY7++
59rbBTJrHWAiVnuG12ykjm900P0oO/x3SuOmdA+op04nBYPX8OJ71hmUJgMCAWrM
sP6LUBthx7JuBbZGbgu1pBHB1fBILqD4BkvdkgcaC5pLH1Qiv+8NCPl+bfwmeRlp
gUD7qzQS4JnZNu+BBcxWwtbKNq1sHUlWwtU92dBtw88pjX7+kUOFyukdTye0NXIe
GQxV7vvsuvT9D/CFEkTRtAB+gDJ7mzeBOaHHIrJ3rgbUb4Cp739vOQQ1uKpUiRY0
9LWje+QDCouX+tFjtnksRrsxpebaSd3ejXr4cV1sW2sZB07aAxBch8DYUqf5umys
0QHPLwUyqbk7zXiNUh0Dh6llOcNfAd7KwseneLsY2/8CrYN31JszH3LscaNqpdcI
X9bMoL0oz9CgDsKIy+c0diLPGaEDT1y7o0cYXGs6cQt17U421SUxXcZd5VPd2B2f
yH9s2ccJ3/E+KjcCkv/UiPYlfAf4s7rebZMtt6rT19/HXTQHlqB/qS+/HIJkP7uB
6HSHrvwUmdxKVbd/UEkTRDQv7aIkM3SSy/exn2XkPc7sDqTDIGSQcbHaDzNUmuCr
XUQTVopU0N/vjZ81FNG4pMmCZbPy19FTOpla+din8UzifyBedGB74eltG7JQimVP
G79PiEbH9TyushlrpI9OS1heZW9dtNQNHlm1kAmrB/feudxxyGOwzbCKCk9Uv9hY
Q4j4gzvE0Y7RuuENWJDCDDKlJRG4tX807vuFTu+QCdlIknfQvsMSzblleZhOSiaC
Zz1Su58qLB+AhXYk1pl18ZFloqqcQ5yjKx3BZsmqw8sqeW7ReNQ+2Shai7WuHP93
BQlPd759Kj3AmUKDx0AmAmh/2jvCOxReMqIxzL/P8e3m7Nuq5BzsgbH70bhqeg7o
vYPIs7NPI+ZWkunsL+GUGg==
`protect end_protected