`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 43504 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
DyHOD2/rTb7/t7SYdpMeYslxXGtdIr11gw2Q/b1cwtUG92paD0rQkWcqdc3f3Bs4
g3BS1Hwn47//22/R9a/vPHplycucfYQ1gXxH/gmV9PWXpPFm9d6tWi8B11Ac2Ybr
vPfKvrlE+zb/smlYoMLTgDCatg5RubMPhFTbKr7tVvOFsbFA2YfMx0s4Gg5L90Ql
KtZLDCvIEhlplFK+E31ZmdFEp4ZymqOWZe0YG3qqrUUsMck9OCWhMR8aZ4Fj2sCF
wS0i1S7Yz+ONN0Qr8AvayuDuItJ9mtJn2kT2pc9bV9yIQBe+ISPAipmKRLcT0O09
VF4eFYX0ZDxmWdosq6u+Aa5c4gKUWnk+8O5ayCmlLeu+U+TSOv6Jou3rj5ZitMn1
E2ZtT1AhoC7B/0jjQnSBWv9+voGprPrDx8SHrkNVOE5UjY2Jr+jCc8fF/8kVgt1z
fWWHvqWAjaNyfTNgdVDf04Sg5rrUfPGAtbahRXPb5kSX3TDavnwRyai9yktcIso3
ArHImodRIP/V7sOqW+5+rqqvKI+orObMYTZH1Qye0oAF1XxEazFa5Bbg8FIC3e9C
YhU2TmR23mH3ILwe0xmOlb7r7isF6B5FWjUXOqZ6qoMKLWqhNkh1iwxt0/YGluK3
ca9rxVKR52FIqwKrSfthohtDzERSdK++zsE5rR8K9SziC0xw40Zh3mmIFAbsBXh8
0x25uaN80HjURynF4tQRMtG8QYUFwEXkqrJTu89btIOa29Q5XSSSuZUUaRU76fUg
z8X4OfnHr34MSqBMyYkmDnRmWmWvaooIk1SWQjeUthUOYnBDPfRIbzNkp60w+1+9
INYfBAeK874Q3Q2qR6hd3C9lJP6WsuYU+q7rsB0oRMjxPL8KpcA9OaiOepBvptlr
KTmcTWvqPdF5fHAHotz7zjpgTLfBJ3UlqOlGt7vXbG0JL3ualU1x8kmqI3L0cQbh
8X+4uVu5iLuCv3dTZ36Ut0QYyYTYfr4JBbBN0YzvhOufI+7HdjC6VgokpCvgx4oe
+lBVyIzKl/u+pJWoVnAzvFiczOkTvVJZSqQsrpgQ/j53nZHk0w2AGVHzMqgfZT+X
lZGqzucaNyAlqWaQTXRyz1Mk/xQc9x7440/qNb3Zcn34tA1OLwY4qGPWX6Nj2G+2
FZvTvYFFrQwCAwFnm70xiWhJZiiuR4iIDPTxPW9fIWrRzvpqnG3FuJKS1RQnDEXl
C0/AXTNwFVn40+WKgq4HRXihX6x+WevgNMUqCUPWTjv2iqvfGFC0qwl/GYeGK2hQ
xMDUw4f9f7Mw64b+Vq8u7ZAH8r7Tm1FeX4P5Vd0upj7XW3E+Ac+PUJQXFvb6XIou
U0il+yB4EmHvbg1xWgpWTW/dWUcNcCMXRzzvt2Uk9RTY0AeGj88Y95Buf/ISv3ow
mX5Cw4PqOKSDmNlbqoLPo99Ltom3VSs80zVLJ937zCqf3A2WnNUDR0hKQZyexA/7
m9I0W8s/Qpg0A7p3q0bT/zHoFcJaOwUme3/JGqR9zbXpQ58uqHG2ak0PlQW+GZsB
XURFxetTB8+Fn696fxXOQYlhxJRsRflHy7t9BmzHNIEEBk3B/Ua0xjoHgASCQcSG
PJHeVwQXwihSoUixL3wLc9CpEIwIKKzxrAQGDtJYsxU03QJ2ajgdVEjj4HQ5UZhh
gm+4vCXjMJKeY3M9Mn3Oe6myufkfET5KxcF5vfeXdevKYUV4gp2DNAvpnCM8zHdf
K0LIgLMhRSvzgwt9S4uobCb6687yFFCOZYIeF4K2IAyWdTZQ45Kfh2QUjDmZHRQA
4MXf3bZXVPWxJAbqqaZF7WJqM5kzuUZvR4D/HJgxIomQCTrYs8HB2vS4V5xXV9eh
JtZdzo1msuhhtsYDW0TagtXFzLdl34bOYTmizG7Ni3U3xeUYTVJyL+o+SJrhGSlY
wAWzsfGsB4gdSv8T0NQHP3tHXhljz/6Isn9sg6sawkngumK3sn1kYZrQI98ix/fD
zV95JT694oE6Qr0jGgzMVhYx/KUlss4uNEDYmesr0sJ6nV5RCJkoodgxG+fxzu6X
IRz3+6Maa3NRtYFHE7nsbOFQpnqEa4ONdtfKDZfWVZCfDNgxH6Bbj1IrTBbTJkyq
0KXnm3hvTycD433HzIN2toOuG3A3oQ4b4NKRdGTB4boGPNp02TfgQUViWVdsLHlV
BZbqjNcNbfyWWR3GyHMWsT1TlqCfZhqyHldzbU28FwMNzi74nkNjp8+Uu9C7wUPI
fze23WFHdMMPZh+gZH/DPM8FYozZcnE+Hva2WSy/JQk3uo2oDascIUyl5aIPOUQy
Z9dHNtLe24ze/Lc8dzPlWPIT6QVj1vY6mUlqh2tRnXGyTKiKz9MUi8BybIuHSX7j
GKXvG4plwfr2Hv0vcua05M75dZ7cw5fWaHRot/pApu/4OSYqMdCvka4Hzv50PADc
NeXVfroaYbXAcFJUE4zLYLqJtvW4/EsvOXw91+T+OyoRonmbS4tZIrGVEI0scrUF
EFJFveXZabWQMfhhrIX8GeNzbaq3OP2Qqg3cDV+NxqswpB0ekpuTErMbmFUc6FQM
FCANFm2pwsLcaIQ5tUsqnw7pfqKc2mkk40pn916YL88SEiq93pV4T69wgvei8Uum
VcN91PVhFY36cO4867EdSeiYx+9gnYCmJ70AIcVbS7i65EEzWvW0CGBGVX8TFtqr
AEh+FwvhNxXWhBHvQ8AyYnaCq5aJw5r1GZ7NMLBgw2f+ZZCu0JTRQpR7pSUoNAnr
nQQp+Oa1A4ItZIX+xWuvoUBv8J/JcP1WbiZi8hzanu5OdvEPkWvt+Rp38ymGj9gt
iNdBshfeAy9Gl9Jyz9EKIrOfQ8hCoJU2NKx8QdIWElOQId+EYelhlAQhv6it8JDq
ZBaKqPt2zWLtJAirndLZQ16IN8oJR0hDLfOWmA+MLRcAqFlypvYRMd57ch+hVvGF
YQPsFpGoMeq1lACCvd9WK0fbV+BdEgGXuT+VvxEtxUcR35W9OsBKlatj0U6exBW5
CBvmuP6dj4wYfml1tRajjKNQHpWiMNofpnPdduRb4AI1UKnmTORBbCAyqcEbB/99
wnuJeUtGyuTI3y48XqvB36nC7BAIZoa33Pj8C3DxFY7zRlwYqYrwm/Ca6QnxPAvy
TukQXjtRiSEdXgXqNjyNwCKmjTspakhr/vHB2++pZv+qyPeui6RwiA/S2U0OdRvU
hKykduQM7rudS5pnlg32gRo02+/6V6s7WrkHxVBQ7LYk6iJEPWgg7GOfL0qpJj1/
YadnYebvpYkLjFbt9xKMQq/rTFUAETtv4/p07GZktaAm7tc5Tyq8H74Lm8GHmC4A
Qvmz+HFKW9vbRTYBeuEg6rOJrwhFXvLtPmf+37IxWv/mQ+VKDn+UULea5fUoV1Ad
H4wfnOQczfg5jdJxmczmzkKIu5G7ImDVWp8rF9t+kIDsn/NizLQC8JGthP+6M0Xd
pVpA1d+o2oItkCveE3MaX/7ZqfGPgOv5yUN/zatdeUPC4njs1bYruc/d/pDkGrAk
OpsLtSP3zVmatwi1lTuwPYZ017fu77YZxODekaFDcwHlA9CvIIRu6bkJa4vmmt+M
Y+OcEqQG9C83jA9J0gbxyrMJufHn4rP/AguxUfykAJUHiONdnz2QxZTNQkPFFOcF
VX2HqU7u/kyLX+Z0f6y8K8DCr4wk4gVxTAkDQYfP/pkyjEHNhdT/BasIaaE0FSGl
fS+AL2UUIbhQivi17xEsBUKEE68+CISylz0Q1DybaoLd8oYKIBm0ui2msfrY11rh
PXO1JUpFgeukZ8tnanpQqEH73ltu/mWFbVe7TSPTVHleXX2ytrBD0NPrhAGn3NP2
75xwnHzhcEelcdeQjdVOwco8CN/k5oB+dgIvYmo2OBivR/8ykPh5P4aITqtDvVyB
MfnNgOlU4fNpAV3aWl1NtyKnzkrLiYz6whCmTCk1QDyMFW0om7i/AlVgXoYiqdho
PsexlA0fkxvtR55Gu2zpbWtPskaCDqnanGA+zjCR8KDDrJ24iDpd3L2W8EUw38CT
Uig1jinSWH5rerHPgmcrp521DCdbkSXWKZWmf+lmp22/4UFOFnYWRH7scNENkMaL
Okq5TXCIjWGgDlm/v4a/7bvbtsmFn7Sj0T82Tqnc1YN8OHkoBEI72Ekx73pyZ+gP
d4FVI72Ve8nkeDLZpnirPl40hihKTdN0tVTgAanm0/gNg0hIvAgArP3lRjqN/ufY
/JT1uZhUbelNdWi+ykzXyRNXw92sakKXDpXVYWiIZJ298rglKjXvbVVMPSILjrXS
SFm3d3TsSH94DAQWXoV4b2uv3j4kfg9ceyaYcNBO7X49WjickYnZix7ANnfONreM
hh1BkhvbTOnuk+/ryus6DvWIiDA2oLTlL79Z8MSEX0VLXJ25jjUwNq/63RcUHtcB
Ux7WAJ/rLKZdSZeesHnVREMLVBvAIu9BUrkXDbAx4IeW5gTHKK4Xp+S9I8NnsI9a
FSPyqHFXn328qnrabyIgs50XB6DsRAIeOXldr3KIc+VK+ibskETQss8E0VsjtM3O
D8PsNMtAKfoyrdaXFIwpKkcVi3P4hIaHtvMVc6rojbZF6vGkm6PtSrf0Z2GqfvfM
MWufoMpyOEWOxGh7mnjud6LY+oVnfOIsHnlmjfNZW74sunC+8VAS2xAp3idndXl8
aMlIuZ51BLZ1dhNoHnQhK4mZbRdj+RnbC+eu6nQpDdm+9fiXw/eq/JSzEJvqCaiS
1FNctArbiri/RmCXcQC1c35MXXeBwoPWuPrG8i3bUWHCgn7Sxgqkl6he5DTsYsqW
8l6bHORY2ssW6299W218jr0MsXY91+Tx3I9K6+dqkdbFrf5ot+fCyYD1MvzYoumy
NDiYt9EeZP0s4dHLgpox6YtwZt79PAtvONk7Yj/opes+EY1/Ah0J2JUEKr5mz/NY
hKSmJRpwx13jtsxUi8RTogvGtb8oebbm3GLNtOoXgkZEPTQ6myMxorDRlRWMfF32
7G7a98It4hbvklN3SlasWhCPmd0m8hb0P+kozIYdSjYDy0mJ5SYJRg+SNekWA0TC
/fQtwjbF6UEjw6p9bf2CaR2BxRFn++1EppU/VGjtT9Zg5kmw6rhdLvc2C7I/Y21c
V6lqkv1Dun08f7oSgYf1zNFIDHOvDMTjyw57b1lkNCvkULKz8JinKz6vepHZwj9l
xv7IMsmq2QZpgZfM1kCzGOrTCCVTbkaO6ZXw2BReKhOqYeI7+33uPxBp/pEGpyUV
9dvcW3BPskfYAEhfz7icznYJLz/Ht3smj3T4EsBAxPZSspkeK82ejdBmFFloriPw
XvZRx0CfpWId5KicY9rQvQ5pU1ECchV04dXiFAo8LCmMsTn72M1LLtgV2mnrpPif
wsU08Bhq1nXfGplbHb8dANbqIXYi4tmXaUn3Ud87iZbTllYCp4YlqnpfF+qV8lju
aqxpCfgZlUOXdomdlb8X573NipT+cQhGjXWo6kVXdgDqg/ZQZ6mae5iDsKYnh/9o
eYvvVzhzdhurkVNIuL+xdHviY5gTEJG8rKYadz5OfSDC8FuHe1AcPgR2n27/FR+G
QjYkN31g9QDZgYpwU/3lbTmzejJy8fBlsZZRNnjm7ZLdosJc78KqFO5qbk6jTz90
JJpIn1fA5GOw5tI+7GDY/T4L2p4I7sUA2lX591TkchcsXTPG2mRV59oGAhDCCBR+
h8BDyl7rs2Ru5h0oCuBWXLSnNvrgFJIIa8Qp4eiCxJPi8s+R8LNvqlqnyrDjayor
++WKIoRifpdWEZyEsyn9KqWRGCTlJUAo1PzZcD6Ep86gi+bPq5FPaABBeUL22KJR
CfoS7/pjWkk6eHcjlE7l2XBq3ud8IdfkF83KqESGvBTvc+1jqo/+GdaIIKT/cDmr
VCv64ghWQIIprZ+1glIso8c0KiNvn7hGP3DTYwD7NzW6VtuoJ0tEGwYpBtjSDke/
UkJtSWrYZL4b+oodDVwXj11nE5fXVrUnqOBEUJ4Lyd80Gtt+NbHQwz/iBmfdY5o6
a7ynLva/UHMqt5710+zIyEzF6xOPfTnlNfS7pS/N47U3EuFH17Xgs6CebPDhxxDw
glCw8WUuvD/Tqk5j35YcFjrxcdEx7ZSpJqwLQBgbel8rwwAyHjAkeyCqa7Wwhk/E
lkJt5GxBCSsBtCBPKeJfhuudb23u9tqwc6K6pbTYB1hzRuUECEcc+K0lcECgVmwj
TWALvqCuhzrglZwJELA6g2GEsf0b2tfi8s7NJA41lcgqsA0X3qrSdmbvtRndTKTG
a/7ID6p2k7Is7mYwDIP+Q9p6AtAOxcfCK9QOdapGKUmisGJacaj66+5DZ68x615Z
5JznTWOVMSg7zISKMqAuMcHsoGJ/bigurSJQ+6sUjGId+C7yotp0J1IXvHj6BoQD
fJq59/fxgOS2kWGxiZ2sPj4sXG/ivzXLMES1A6OuoNp5NEGZ/tHILtuTZV0+/7o0
8ZHDgoHljxM1IHWbTGZtXBDYbaQ/LqBCQjmijfdB8ldNgM2l6dAdsXdI9nMr9nyI
Of28vb9/CQ+WoFRQ+nZ2jfAYTqMQCmslgfIC64PUczsY752QQHyuoC+DNoSY4Y5p
MQR5vfHBFos/ltt4o2o9R33QbdfVfb8pdGQIaaW+M1M6/QRbmXW38W7oHC/bL6Ck
/djMp6brzP6pm+oWutTVhZknV6TQ43XaFSXOvTHsj7X0EvCF8wJcbeR+xSd8kbb3
cyKszAq24vrAoXMltYn19Vjyj/Q1sEoCtiFAZ7/BFxXolCUEnEh6sOU+BrV5Jsal
/YxaWNcCjpW/Hk8rFRrWcdNmHBUOiDi25kQoukGqP3R4mURkdsZv+gjZie/37K8I
+RO0a+7mW7EbYhlfOfbfzi8J1nF/zFMmB1i2BuRfwItU1pWf7CufxxumCPcpcRXL
Ruqn80e8rwrxpZxUYTSUPd+7nEgcOxE2PuA+AXRfNOUmK5vH5yJ6IyCsh3nODNKf
B8oXZ/Vr63BFZlQOW29j4nXPG3j+edAhnaczLyb3of5y7EJuWd5nZWnh5HbE1bL5
S7bwnC0cR/zxmGf1JwtnIlj9FkgGHJkv+xZvo1r8FjuY7VF4wQOwY8VJugzIgaJM
bU2j1Vo/ZqlavNNcbXGy++CdkmDt+SQarvA09oAYbYkL7gHhRcQtM3CmyMOXhtvH
OC3inW+LqtFsXOuSSTnSE6WTaxIS0LYKtb7D5WDwmwTxHrqlzhQSBxU767ZKkJ5u
z+we9HIgY3Oclg/ZsjXEmCRMwh1nsIZ3xeMP3+BczgtTHMj1chm/sMp/5tRQgLoP
wPTjkCttusSyi4OvhKAStPg57ACjdo8gai3m5slzeEpqJn7O3kwkDbMfiOPkDITJ
yNsAFQ2NVOmbRK6oNVHw1I6e9wAqpiPZIlJbfLIAxPN6XKJCSUxbl3qFHS6eM8nn
o80UCRoJOkiKfZk+bjbHKl1qMponn9YRiYypazHZ2Pdf6MiSK4ehkxOyfx4LQovz
shBIQUrpo/srapjK4b7a8Py65RlSGF7DO8QvQX7FkCc/qOZN5vReGHgFz6cApaMv
Dv+UZNU9m3R/NMpep2mtvScjWVtRaGWo/m9erkAMJYpJY5kw3RWeYiToEP2OmPGS
HwPAyUqJ95HpKLAUdVB94xfd7a8UBvfp9+tEB20nLmOv6ViC00eAs31qbeMU3OOL
ga+H4SjeYUEnZO+Ph5jherq6IlJOQenZw0NBJL4N11NnOGUxKbI87vzbM+P+JR13
GFJuXLVzW5R+3cXpwcl1aAgstz/0TpitaHmtrtdhcUMaygNBdXQkUFBV0mCK02DE
GYgvPg7+RFV5Lt4DG2wkJmw0P21+5b9ZzWiXLshZsn5aGyczhqu0HhycYhjWQlPT
7xLmBRMINzuWEAYOYHwDAHDuNiIxgbv98AFdEFEdR5EGE6avfJCq9jG7lKKDBDNM
AzY58ztiltiyxiDnZhXee8HzKkFI6I5wudDmvjQVnkrvZ2B20b6Lo5vgfCZStYdn
F0vhPQbx4MwcD/9QjIgdshR5cdN+gFpcjvrqE8xuK3PBjCrqVJlh1JBlhrePrM3W
jFOZ3a8XqRIsiq/ZrhpjlMS5dcTneh9d9DRNwq0ZoMEwy0+zm7PMg/SQpkOTCgHU
QElEm3M+gneE/uPG5X59+ZUE0zJRvizN/vTSVmBJ5lpRyxzqkG6fNPz5+rIS1Hpb
PD3lChBQysEyyLjHLKChGNX8zG2bxlPiSno8J/MRx6qb0Sh0fsd64gBAMAaw0rGR
j+8GDKBQ7+N21M3JF1+2djn3Tw7iIXz01mbotkZYMvK2QOeLFcOYh0BMDRMbqvEA
D8f2e8A0N2tO61IHkXhRLg4xfyFVq2GfltUD/uVNWytIbQMNnFvyRpKRFjPQkV/g
rpQKzi3/UBiP48LO6WZz2Ck8o8iM6HYKsSzkXjCUWwrF5E4YNKAJtm5gHuPCc0A0
lSWuf3XViId9IrsNU8a+6KuZ2Be4c6XdEEoIGWSdt+uk4XLtCC1lvQMP/c3NgHYv
IdyQFMVtwk2+yRVYw3fOUmlINIBzc1GitTq2YKt9EpolXsSU1gvgZ3/Bh1CFkjar
iyg4ZDUZHNCt20rxT5LPNa0vjrzCGZKrU4teQoX/h85rYVfHcupDkdQwvKdOv1h1
v+S+sGAm5GLh5G6hGAuBoXsW7FWk3XVzk842/SDi97awme9zf9ZTYlJJhADG3acz
fyCN7n53Vi+f8hwP4AeVdAbQx7xtX3znPb7a6L/FceHZWIdAdsP995AbBaRAykBs
nJOE3Li73kXiFhDF930qaqJqzGF76SWAIzVdOuZwaYhpc20fPOjxP+ad5ns7go8L
KRSASXHvfTeNExocrs/Vm80Rttxne06/VWqGO/aUgkm126GOArp7DjU6XjyyIuRi
08oX6HquqtjaV7G+4QJQVQSkEVY7a/TKQx3p60v58Uw3Spcqqpx5TjuosUQ4+U0k
DP8OzwQo7qNoXAKRgNH7lYp5+aNKg3g5+UCoOzcsqYO7ySawrl1FgD/0HvGHm/Bd
0OUIRI+aFNyb/mMJ5eaaqzoZpvzWmMSzoenAhKim56gcB1S4KGx3NqvKoHSR28Vs
Tnqbnvrku93WmFQTZWKNTyUcKCrPyr4BMN6TY3X+tLl6BfCHMYtYg34Vf65L9Omu
8AQ5h23V29JRNoTtOOUcgj1M+Jj5CIFxL4CkvbATCEJjfYmHvmexruDXdq3JkrEN
2LwGQbPescTiN5fVexwGRgo41mYOQWrHY/J6Z/oF0dRSpyQCRVUKMnDQPm7MeVhD
recKiBbpfoUTRf/Atz56NPJp8kpkBVc+aE0JquGfDxY/YNDU167mO1mlT90ZLqd3
3HdpVP03qRxr81KjMCFxLiFt0MICgn8D0DvlF0HFL4SfeXL0CyuNgOjBR+gDaM4B
DYpcEaIvpkMQp2+Z78EJoD8cUKi1HNaTBa3vnI6WRvTrRDMnBm88+/Iq1+mnBnw5
5TzOEfEdVjccyhFKjvfoiy3XPTBi7VT68K2Hp4LNPYtsfDyRZ10JDuYrIQv9JaEU
RQLxNUHDEYe+SwrfUyNIXFUprUep10RFdcjpA7XDUacgEwek0Gj6u5NhVlteXICF
0rijSE46R8zEStKIYQQKCmAxBI1sy9EKT0FfNK5Y1SseNxw+u1TLuMZD7epYW35Y
vdeGXvHq+S3U+CgsLGRmg1OKENQDgVJSca+Gx/xNg7RmUT1l6zdv3e+UJa9JgOEB
zeypZyPX/EtKLftYUHM3yygl93OTO+4xiGm8Dp3QqLVfJkXDDdcotZm3HY+TTcjp
YWh20+29V6aSQWp5WyeMXHFvuUan+xQdTVHYFGVkFXTqsceBWLMfLDvHocXflsfu
uvSnXdWAxn15/TGCVP416OYZ3wVwGvFK/WQe92bFOEhMXzJJOaMWsskFDSl8A1Oa
0qJM7/LOsqq6GnZeZiXRWMKE1pPw9E4k52WhIh8utbJetxLetHFSlZdjMKSBTDke
87N8okVgFze4pBB/HKF4PvqF218t+3YLjJioArC5jTv3pwldKWUWXuLeVDKKv8EO
Sl5a0WlnwoGzZKkntTbmRi/DBvpH90TKwiCMz8Wddujfxtxev/68sJfOUiF2hF2x
eu1RTbfjZ2bmeKGdRJGXKjqX0ZZB9GQ7brnr1LeWgUqEfTBLb+mrIGSm5j/ECZvU
3RqNILqQbj7O1CQh0zorhJ7GI7KMmSokP6LBWfb0p2PShE5zzOhbQTu2IwItSLa7
8qR6GyfAk2NTIi5GxBK7yC8uPx+PqIfCd1yZTT/33UcefLJuhW+5ZVc6K27GrZMe
+dU+q+3/ljjg6/JgzHS5ALIuBAG4euIPEMf6grnxaMwtafNMZsDCMQPQqzw+/0Ng
Q21Ug54g/vZXyUa6f5ePkv7V0UhDdjvhd4fZnj38usjPxdJnTX1cleZQLYBNvFO1
wFZSORXZxRm7dz+WytMc+kW9HPjKU06bm2A2EOi3fslfz8DlbYkmciYtzzwwlgl1
58ipnJJR3DHE/VWm5/Kyc3VttPxmpyH4pmPwi46SDMOrr4kWbi42MCLYdcTH2S8g
xeyWbuCL3qpr+U3oqzbrGQYylivzwDcoUqMwW9qE0/KKVkwC8REtFEb37QylJ572
It1zOqBd3milsF1b3Bqbd/0WJqOAaqXO+zT8qmQHjNLr9PxtJtDDng8/7CtIyF1y
i2t5KqL+gcH5U4askmLra24xiGxshaQOkB6J4L+VZGU9FheJyKZhvt1udxqIhiNY
+G5l/Mij38uUi7VURXq1qUQYqOvxoX+cUSivhODs81d3E/hP45BWL+onczhgB4be
2Grphx7m9PSVPVKsIYzqWsqvTgokKulXXGNsRmaFwMKDiuEpFBRDrhKQ9B620scz
8N4suYyGIgZ9eg3tUE05q6VsuoODkGSP6RCzQHF3xgaj34owb7Gz3s0Rlm4mPg2A
voesRCtMekasdpYwNk8vAiV+qYv5eDS/YG2saC/fAxsdlVkWLp0jaQT/xvIyj0tC
dcLzSlURQ56BGAOOGRO635bBXOyGmJO18PntXNyrF3zw4J8sBEC+YK3TRYLEMENd
7lBFBSg8kbyDjzdSocUh3a0512guo7/spQOA1dvE6UQTKk7I0ti9gRons8Os6f06
CJxTtE16WV95L7J+MV71l0oOs2PIHa85N1u6dT4g8WalaXcCxbKogdETchycog4N
qF5lbCCWksckFl7weTVYBapU7Z4L1IidBO3Jv88CKm4xRBHUu8ZYZq6a1vt4N+nw
Y+QRGQW5YnMrf78uyHCkAdnl3Lwl+HagkXza///hbFPLXOyagd7yXZvBbOpi0uHY
wXM4PwAgXD6STPYFTTta14LZZUp80aw/VqjHndq3dj1AV+6yrzT2+S54mE1yemue
fna379cavzU5mMyUKewsoLgELAWjg/8h0EUUUMmc899ws55OdXXiSWwfJJsJB9Ke
EvhstzgUZUrpEsZNo2yhZH6rZc+KlhuGl+x4jxx9Ec6OC1kHqrXOYd7tqGdlO37S
VaM0lTug4KL2atHUZ1SVB2b2TZ5ZCpnYPaWUDiHr7Mm2P0ROhn4ti8z2LqeeOTKr
+93AaCGi9QRu9p9zwFwuBexktEvrX+X8H07OUv0fAn8c8MyU2+oS6pH46H6GxEu/
q3OdSrdOEMuBEhozkm+wB93bH2CPu3/Y5+jAFUhprg8fuQN0u9doEarUvFgwoLSf
oadH5LzNyWoqWRK62ApOfY///NNpli3f0f/ggyf3qQgYiSLk8Oqps+eIRmJYPpie
a+8M3/ub6w7470VV9QdXiANpCn0C48L4wtHhqsB0rNM70iWNBLpDb5KENDtqmrtx
l926Spi1vP7sod2uAMrbsJv1YI13oisJ/tuhb5Gz+lVoOQ71f7615ET2SoD+aTQ4
2nOkM7ttYcef08te+BUEnHT10KwBa5HTCVV1I+GSboZGD5in+UUtHFY+fRwEUFBx
zNZphbQMR+Z4rxs8X80Ak1aHq0QSibDaqpMGjp+n2C5+veNRn81KsSm1QxytBYOw
L8cRdQNd5L/43mbGE9LR3eXQd7jOpKXD/22pmItwDPb4FCKZ2G+zXMe8u36JHHIC
jH0X01vlKUBRyEGKynU6jcj11pVEpY+Z8UG0Sa4P0C4WOFus/RXUmvXWO9U4vMu/
VZqqokaNoJhra966aY6CLp6fyhGcr9c6/pk7h/NFJA91eL84gG3iPpYd7k3EVCy3
g31B+I7Sl2muPS/Ocuo1OLamsuurKtGrH7RyRo8Ou2zgO89j962YrRH6K4gI1YQ5
wozDTc5hUtb+yPMOrCO4+SDvSPAu+rTsD4u3U7/zO7XqgstpgXEfkKWS0FWk/lX9
tgrEy8U+KJ8kBOSU1WKcEd40uYKEEpWvvg8Gymbf3UJ9V3BZwiuEm3nC91uynX5Z
fv/UD67Ilcnp3PaP7FvRr0CP/DcqNFgI0akjzRhqfctbnjIlxaIXPKgSqNF9kxwX
MINpsQoqJV8uqDova4UQPVgAarX1k8WhQeuMH3NJVLtaYQQRc4y2RjkG1kNozrbx
pHUE20x/LbnRN7Bs+NJ9Igk3FBifhC3Ne+P760ywMP4NmJQvwfnk/zGdUfJUwKvl
ygHzI9xohAI4qw8h5Qbg8O2DPG+iv8K4etswm/H+rN7DTU2dzWRMNRp7GcW2n7dd
3DFZkDNlIHqi6VpOAFWyCGYvlvSzF5rcNe/pKoq4bAnSKBwQiJz1ilaPKColEL/j
g9fQ0ATn/INfF9vahBbvaWkW+qFGJfHwJA/6OW9owsrpG+4bLzooqMhM1XYLJrs6
Go21c05n/hSGmwOQtCqNP3UwTGEan4HpyFCqGwnA3lMyUoSsNsFHSRPPt/8gCp4S
BYPZdbgD05r67JOBQN9vV/iyvhUdhun6+MlArjs4mKpCnBWOfR/aWmRLe26eJ2XS
+BDx0XYm1ikGIZxAT3HRRhEHpuK7DEZT7v5Rsh5SGYlhnhRTBIO8xZNWnWcLSiun
iH6Fy9JgwCdS/z8wlY7O4aHUZqM8FGVBLtrKHzSZBSAw7/Ozi+buBGsHyfR2CTAQ
ROFoYp908F2OhO5PhmPGFpPINQq75ct+eRKbJNE55TZK8tFmSkv1fbDJl+ahnAd8
46eZp5aSj70wD8kffJQ6iZ1VGhelRtYYDUvOkLGMPmeIb6IbQVV/TXjduWLaiTrK
8YCtJYN7dWcVs8ekH0DViR6ljaPZ2gmd+tn0W0IJ53W5DpoXSfav829OlkaV5nY1
q7odGNqHLGxJY4JT4ZSa+3NbVvght2NlM+nDKPjCT0/Oh6xx1Qr/md8sRLL0zCZw
seEXWkMYI1tKwh2mJzC+8JVlkwcg+mAak1s02az+AKmmLQ8t7CGzXV87uSvqgCjy
8aTFph1Ux0ztoSxf+5ckLY3173y/XEzmGdlBmVKzNMESeadAKSwYjY+pC1XjwvIM
WnPkVzd25B5nOlx1TfYKlJC5sl6cHhfz7dIhYec+dqqFDhjpHe1WRSZ4P9FnIMTf
dzmVoNOMIDGSl+/7PSikdSXdQnOJbmxFuAOhuoW9mRrkNCFxhnPJ7mo7yIs49kMU
CJ4D28+fJR6KWywPE2yxXGQrYUWUoMHGjzJcGOhP9kAUMgFzQVhBMIFsvvsnFKc4
+5qR7zrebFM6FGo10TabZTbJLfQBoRT+D32w5tVUqYfu8yDmObBYfBPEMfrtSuty
r8lqxoae/Ahb7Z5ajw1CNtJEjTFndx9HmkwMvtyV2qhmEil9qsRP+N9onQ6bsP0c
3ROj7T7Car64lPOORbbv3DA9ycrT+K2hA1n9Z9QGzaszjVRX/u1YJjJBSXIbVXuG
2X2wUfe5P+4u6U1p6Mnicgd6ZV0y82W5liGF+b7csimyZh8mWA6HlxXT8vmOY5FD
J0bDX03VETGpfRbk2bRB0ERlR8qSVrTm076IdbRHGYbYkJA1cIyT5PAQxeYr9NqI
+bjOJpoqcntHtst/FGWc63tFWSW84eKMmLNJ9tCaxFgemYucVDZw9udtKBfrFTk8
djjgu1+e5vRMu08Kb+XlgonxNJdvLCJZNUKmnwzEozk3wP1hsNAooEXziNlEKD+8
73c8LPcQdPqUFdUSoS7t8QIBjnwX+O8XWjo8AFhIrMQbk2dbiHssRO0ZqVkqTfpL
Anvm8iHJ5mtDZ9op2PO80cySdmqkzHyVL2EPxCJKBHj+bVk0QIrg/aF+aYTbmh+P
5+D1ghcBAA/3tuDXWOJQ45LCJcgWTSDdPYAWAzLuFUQ7C+CgqOcHF8j6aRfKpI61
axwO/DcJ4CUCeCe1+rI1MrZjEmmWQfxYWEGv0xmblnW6wO4JIwEyBkILC1/jGcea
vc4rk6FwUdLnAjInplKdbUpJH6+3NUExGWZWYqanPBp2BUnKPFZcJCCBuA1O/TDP
W5UiiOPAt2KVOr8UM+DGJBZdYudzzk6RtQdZL/3QdQp99KA9524JcucAQpEEeG/7
7z/j0ENZPL+0sxPOxFA8sorurKkClKH18H1we15MO6uqvpI1ZKQebvYHOhtXYdpm
b+KbvTU0yCPxwIQQHMlCkJMyMoIOCH6wZoyA+XyXOfZDr1PDU46ma/cwtkbqMcjq
eV+Vuy2+ptsV1kzqEQSmIj9eRDOcWv3HJBMXokVD5pf9O/oFkieZ5fQVpILuXFFx
QfMXjD8Nd7s6sVcH01BRDTwgwuDwof0DxbB5YDE4miMMjs4/Fwz1pPXwH9a2V2CR
bOvs44yiKiOs+Hy6FNmgNMDe8tacr6nlyiu9OX+jJZ6w7AS3rG1AQ1Mx2lt8uaFb
3nx7wBygKK1U8k6qb4sztAPsKES9CuSJ+J+cBcoy9LlhP4w5PHMCc/XylyjDmqVV
n2bZVfDZB1fW0ySVDJYCzHMNryfqdADkaH0Ps9IrruJtobnEuU2sSW1bk458j89n
XrfgEgHUiLKEA1gH9iYUnta9wdlYGI1XrzrAvOfC0HinHvk5gxhc4O/y3pUrKmF9
HxU9A74rKOxVO00G7sOOnMWxIDsY57pgt8tVhDMeD6uG/HHRR9Ks1I+SyAFL7Drf
C47BL7kn6Tcj+O2vXvqHI8qyLiyAM+7qD5tfecUgibCcu7cRqXawDFkY+h4W5Tb0
oVZLWCxDbXjHvm0QzHiL7yix3s1UDAvm5qJg8c1LUwxanXh22tNqO8lmezJPl6Hi
EnHxNcgLKQp65L5y2VMuLY/Hh//oxRMxcYSnjWL6pAZ7AGB10fiE5cGT+evrVd0R
5ql40y2CCFUCbCq+qgJyD9ZjpFHgqA0GihWZS6AGSpWLnWnh9gbO2mpupCnFsdkv
jDeP0JYKcJDsjs8zRe932NWcf7QH/XtSVW76GRkdAnN+frq/1OQYkmfqAU7y7C8+
kA2Q8H55H2kHaJOuQdbqnTY9ni1AdUdjdL4XYohCKAE15xSfwW44AG6bg2lPHH91
AGr6Ahz5sVDiiY5TjDKx2gKy5UNqgzp3+9JUoF+tbgUnuXuXMDtZCgfb0shVFXq5
kXzsT1GRtVAPFOupgIlKQKI2yq2AtnJ9ig5yd2lGAW2WS1ocKTdqhx/8VSSEpqVI
yd2JECxh4Ih2RrlmtXrh9hr3/uAlVj4NoDY3sbLu78sqX5q/BzVuj1RBCy4AMGEq
q9uAMe5de/lb866uxbZ0upZ0JI1xDWu9pzWFqocJ+TwMn7XaBXVLV1nkQvgTTyLE
j8dmTKfpi5o1Ubvl9/60AA5tYTX35/VKfX/xqKDHIS6YIA+jvEEeMwjbxFPowfdb
PGuRYi/l/zHFlGDBnzjlMyoosj5XuVg5KtwM3gYxKjhu8pqvvql5IPMGA0r/xYR5
yAxZDGLunhDeuauvbfjv6Q2LztwWlBohrDp0I+58sX4vFpj+4ItktEXyFo4r7ISt
gAe0YvnKPh832E3u2i0XquMqG/ACoDq0vgTPKTlfTSoo+ZZ4rSQLeq4KRSsZDXO9
fgjpR9GOgNYvLE7CJI0xrRXopbbIEPMr5Zhb9OSk7qZSFc5stsoNMj938NAoxzUm
YD1xVibUG9yrSbOt1u8cEQUfyzuSeHx/ij6jID2sx0KiHkcfU5afWe53mBNmpPXd
unh5wYRGYfpCns2+S1+ze+QqRiKPtbakLBcUTgSwxJnc3McCwkaq1/u9sJ0B/qb2
lHzbVCOiDafwOFenGOj7a53XfXQifcMoxEZgkgvPvaZzJ5/A2eyqBqQqEBmDcB3F
cy/OqrMLhewalB2+adS7lutJh6Uu4d0ZIT4ZEnTafpl0IVie3qRiaCinjuFHG4hn
Ze751+dbvq0dwyYjwjNHlUPVRxeE2rHT89N7epB0mxXMPjO52hELjO86mq4OKVP3
VDae8MZ+cEWZxcnWIkWUlFX3e8JwX1oETS+8OaSjAE67uxwPkm32lUQoTz5orRKD
vf9As0INzuzJbuWd4FEZwjOVz1ipRex5DiygrVAxauCaAjDELOzRfAIAK55zV9rK
nbOwfOv7Dk6BBlB60UdF3gwT4N7dx2RAu9dFDM+rN6KWTpJ7G3QVOXrmrc9vJIW+
TE33BK/XZj4CpFHyCBab68ITmR1UUF0JVYVg+zNGhhM3FK5TR24HG+TMcx8PKE6C
KEDXvq/ZP9J4aKsTNR1PwkwdfSFK/wcoeTw0z2Tt6eNsOtasHhJBXkDfpjzjJQnz
HMEhzvJt/ddxqP6LWjlWJoMU5nprT11r6Z6UIMkQQBWcwScvg6x9JbKc50AOvEWn
j/w7QpCkQsmpDQssFvrPKrAODurVSAGZm9+JxDjOsoZLjVO1BS8IDUnAwHYkrUq1
6EeDdINDiFwmfZAeHouKPbpGyk2aB+VWFY9v8Er8Z7FsqOgbVo/PsrT8st9plhvf
NTNnHqcebluZ9IQy5GLYrFNcfs46IZY0TwMxJENtNGN9OURi8nJj+KAipbr0MGbP
ihjjamxVGbVEz94Pea9PungACA2Yx67lg5g6/jhuupSSrM4acJ9zkWdlky5YJmAj
pGTISkVn9JRA//2OTl7HfjbHDeBSn3Lup8oSD95d8n8uLLnSkLeJdVCNhSd7pD+m
nwiKU5wGMhDHdpmIvzYScnfldIptLVq92W3OcxL1J3S+PSPQn3G5Bzkzx6hVyAO6
BmMgvf4X/H+r3xr1i+YnqWd5OSi592MPt5aTsqWJdywaKQpcq/Zyr5QhdBJRj/2b
Gap+ZCjt3cYQxWtUIXYfAgXY7GWwqybcLSVzeZZ+AJrZfXbKTa6crfmqScr2VWYn
FqTmoHx0loym4KUeBOXlQOgJRbSqJBBm+vcNnmOirUzqDMAh3zToyLR3ClPZrDKE
pvY/DcmMV4BpTR2rGo+5P3jKq63wShD34Lhl2ieOik85Jsi/iUyoLwJfPMWqUy/S
vRBME7K0S+djlXfssnTSV29V2NpyXf1QtZN//0hlMEJsMihzihL16bRO4MuL57vn
gr4B2KJsawgZvlDXOtQ1KyotsUwRIbaecjdcGvfxyOPZvskum4HV4snAflOeaOjB
QZwC8R0uzl7g1BcVnlRmSEkYxdk6IUcbpvGXIi0VmsxnIjqjenFSc8gJVt3ff4NP
835Rp23dirdO/pEy+pNjNIUO/3Mn30j+kDixeWXt0I5w25ROSJt6wfvgjyx5nRjg
0xeoO319sf5si41AywBH9WvLudhbH3D9Q5ce6JWb32jlgXDwGkImHIbIkHdtkaa7
SJ4V4QQnjIaJWXbx80i3UAKAdBaK7n/VQhaXjf5DlJadnWGG2ODLXDjjJF3zA1GU
PVK3JnYwYSgRkyNBsO1vui/awIp3CXKwezYgEMQh3TPVslSsN1+Kg7tqkKHZw8JL
K4daXs0jyXtnLHd1kfl0p3MOJZx8AFngOoeLDGpGCxIu4HHigG3ZG2aKFNFKPbBP
R0B9PoIsbiHn0Qyel+jluyVloJRqm5kPgz3pV9PGxCSyEjE92A8AjT5bRq3XI2gj
fCIgRz2T6rOtQAseYIxrX/A6EDV9aV+xADHJnWO98fWQ/EWIhjVn7uVD4sXUcP+j
oXyJR0d6ojeYfPm9a2qLNNdIjnyJUAmQpf9RVKw/ITnfd35CeSGYg6/wpEt6ygJg
9TswlEDE2VWSb2kq0Sw4+PKS8XuAHLP52nrWNuBFry5Iq7MF4GqYrAaf2nXjSEY3
QKl3lAxjk4giVLHQq6If827ThiuBC6jMdulzFfOw+Mt2DanyR7AINTonPq3zQ9ZR
uEvWokW7t0QdcRT2UQFK6+KDMegKs7/tPavLdu0+A7/B3ofNoPKaBV81GHpSgIDE
e8eSmzpaHUVybuylGOoI9lQPd2m0gE9AAesTQl+ybUPGfWn0wsFYCmTD+HAw7JyU
z4r9fAVjcSatwxNfG6raVdvCy5MbQaWsL+ll2qdF8zLVtjMhW9lIa/oS9Ooasoyz
/SutRAdb/i+J4Pv2X/ACE5FIc4jYKbHtjbCDIxb93wG8xEjOKmpTQ31yHsKsTWt+
dS9Y88PUY1UVJhKlY1Sz9Vq7Gb8IIMA/ibxsyax8iAjN0NK+PyRbq4HvziyKLX8b
L6IcGO52jSXok2K0Mpy35vIQg/r+UAT/wZvKp7gym53n4M20nU6M+LYfiXPzLVZj
1FiBlMg92XJyzH9Dqm7+GMw7A1KKO1769wEZ/nWifTfk8VTLGnYKts+saWDrYmV3
oZfjpCLJeq3RUOo/xUklkMh+6BRK+JH43bYHC2OGVQ77iQZfHm0vdYbHpLqrDNZh
pJ8qqC7OddcpeiQFBeenFQmJ9y8vsbjddJ+qyMJDPrJKDV/pJO8uRe/7SRotrUGd
AnVXj90jUiNAHvVO+tnpoFwH58hpFfZHt+Ab6lnilmzjD9xLQE2Yg/cyxPoqh1mI
lnaHioZuNUoiELQ9ytwthaxlBO9RhcyBvWxRBVIpTZSjt/D+p3ebb0Oh89lxuc0I
FDCMZyN5Uc3uKJFBRGK35hxbRFEB3uu+uPsoPPvbSspUPyAd5byvFHsGACOlFVV8
1bdH/aMn7LUQ8Gl4Rd3LO613MFzuHhRyj2IvSNuksrFX0GBt5T+4hgLyCR1wRTWC
jjdOBNH2QguFfJj6LSWZd59XAkhuaz4DQvA4euSRQPLf+einR3vpNyoTtETD6KP7
gxZfykVz+kJN3QocOiEsncJJBnK6vLu847TzvgYBb3cK0ieBhRj0cS2Wx2XemwEf
U0O9XflKnYT+CAW84Y0dqJDe3lFSMDL6O0f48Wupuaqoy0wR4sI+BOL9sm+oheA/
7fnfr1QJQWz4bidF14P7bvaeBRVXstgrBCOE9UFwsfqWEOqguCynywZzImQYk8zl
pnCiB6kWY0UVzUjIaxwsRb56Xl/3tLeRhGvjFtstwu03x4+wmj86xz98k9dUPN9+
QWdTJk0Bupy9HcHZ6QIKsVFePQLy4BgySfspEAblYWJA/jPirol/ohuAcMSTNKLb
qbkYERKlttNwrNi69GBCbjuvfBpDzZ2+pTUVra2fpL14NjqMc8gGKLjhEjQnRg/q
8VgsHOBlPh7age9qkAgw/51r+5auYI9N2kGjOiqfIC6SV29OcRcjE46g4FZOWZTL
y4tGjIV8cQZwOl5ZZ4eFdp/3GPqzrevxfWu4KXFPq80DBFu9ALIEkZe0+R5KJAF2
8VMe9Twa2gvq17w8yge/3/gu6yxphNJBUfBByIJ7EgSr3CHNTwAfjfZGoG2x0Odo
fFrHgxk9I931s6o1sffE2FF8cm6KLuZl1ErGYj3xMqEajaf1hmTrGN86lnxFgqKB
QAg2Z8mwaWbBZMp7FKklKQCUAVW9f6q623hkRPi3f8kU1nZuob2DZ4c2MoIDOPFJ
cJqm9s8IxX1+Sq6/5/Nta022yG+6FjQjLbkLtkuVhaSTvrs+CdjL/SVKeSgmvnGY
3ARSRR8oYnH0H0s6ZEl8Opa5sv5HVy6kThxfXbhsQJjM73s8Js7JTxtNdu25O5Q0
6rRjEskxKZ9hFh4YORUM9GdodOts87hysUVQoIgy1P7qu7w1Juv+/jKq71AFNnKW
QsCONHVSUS8uSku/lIix7ZJhcyHiELXTz6TVWzUXVkp8fq++AUWSiYe0BfqdEJKn
xrCy2JFMKjIKz/RCc30JAOz9uCXC6J41UmD4tiSNpqrplWoDVq7cnCuktYHRklV/
dwCaiYRnpNwp1kChMUokyFLmNF0r9GM16DjuNVKNmJrzwjiIExJORrHjW0rK23t8
GQk9HcuXyO9lD15mZULvwKB3WGIkRQSMcg0+mBQh7ftuHv6pkyyFeyB3QcxZsGLj
KVsULTulaFHpXWdZ3XTxLrszUR2+5Z/KbpLdHIrhg4kat3MPXd49fvtC6ZM8aApb
HM//swUdZuD04lBVsUMGv9B4JqhLEzB+dJHy/9MzP9ZHoDO1wtfgY5P5WduPrkjw
DRvmNguv9FUXWcjUEgqCaSTcwcZTWGO8Oo/xz2j/ie0xArFUjC4kuSabazPxgBNH
r/VpknGeb1iuW8mpgI4PNSpCcjlq288s6ANYUkCSVEKlYjM+tsa1VIeOoiOEPeJq
cGtQpBAJIgShBM2aiiwPPe09UtqjXUZeit3Mf6dSSLi3TCOJjj9GQci4cxglvmvl
QJ39lsHEee5PqCo4CNrjwka2gRGOhxpx7fxucw/NF+y8+CRukNQVoVFuKq19A+Ke
nIQrvho/EB/BE/mnApmOmKGFdkIRFM33VXZ/XPXimdcMGKBm55jCOIK1rcJE3YzY
/Rknacy6gJe1xYoQFrfhU99U61BvcGfAXfoIIoyyqfrPWo7e9QauARq7HpMRxFCD
093qBB9I4XQNrs3p7e1TL6Jj1ES0Iz95fzux34e4WycuzdNESRq08IzT0HjZSBqy
pkLGORzYAEEa238ZBHsaN4Lqu0cg2rarJ1eVX9ZSaCW77tLZwH2vPA4/s5SYOYs/
lukYZ/Xh5QGaWRf7kqt/Pd4atw4fE6wzGKUKUmOx4arPE9d1oFy0wURzIXTRVA+1
9yUW7QfMTlLlU0dLkKJR6Gcl5roUQMJ9wbXnxLw7DGHBf3WbMrmvabzYo80L45T3
ixsoSjxFVImayI2NvDaZoC2zeuZeqBw9Lgvxmga2Na+cljsSPy2qxUMCx1w9Ex5I
3UnVHclx6tfB7VCIsxUKFZxXxI4LTSKzygCvU8bY+nDNOWT1v1rv7yBdPNZrtbxE
Nfy2OmyKWLrDoZTVE7TVGOKs1tkMNUrHn8dQXnZHr1nY35A9N5aLYq75z0oRsfkX
f0ZSE7Yvxba/OlGFeEUedMWzJYOFYXwrj2tBwCSC6zipXkfRtk/PDFq1OtpJIMsp
bEVoAZGAMZ5aMbPGu5JnkLoFlSwzi+IJia45IA2P4YOQ67PHD62TNxEk2gK5BHsp
yz6c1bJs48UzU4c/G8EIYRYscxc0mKwCgFo9P3kZVROi1dB2/ifSLPbErmyJtXnE
j9JNtkhqqMlAW3OWiM7pPaI3oKPRbeYLTh8avE/PZpUdgMQRKTGlwkQcV1/PO5bG
bjpH4CVufcumMmOcpM7LNNyPF8LLTXWMSjQHs0ORQoOHVShlnJPuNlZ/XXGUYBLu
6t9IskxrxNVqJ2DTG+cYpMuec9qj3z3RJd1ZXn1QoCZOigwxQNwltHlCAovrNu5I
NB/KlIgdoaduNh5jXBAyfOb4UT5jGLXWa9Crz9rIWpdUJ8GoH2kvAsp4ubwLDE8s
SY02ewHfBsrJ9CPxDBkiDWBCLWOyR6v5AmTn3IO1xpa5iGgYDMMhRME4sCMJ/+AL
umSh2Qw4vky92wBMAZxlekQYapotJELtpbVLBgyLAcjbcKr6adhLMj7LdxHBQ3it
TLJm5zlBiKiMzdK93GFq+EgoMfkm938HpoOsc9oRbgLmdfAu65ni3zEwgg0bwGE4
BRHf1LQXR4nLn2MOw2ckLltwmx0VDUr9skFUNB71tJR1Dme3zVo94rW6rhielEUU
6IGmub22mwkZjBwJR0Mhf4lOAgS2Y/SFQ2PxP2XW71E/hKBTaueVt0jhwYqT5Rld
0X/MYSYd3EXWAImW3AckCTPl7IWcXRZOTSGFkYpf71OX94im1VYJ58jBa2Roap31
1KvXdjztGbNmZHkjzb0mOSwzpLybCe2WsHXmVkoS0qqyOEA7gU1n3iyZ772l/1bH
C7P9XNjYyfqy72A3L6DPqu+OqExDMyCXjZPUh2FbqpCWNtuOa4fzFohnV5Penq0c
9SgJ8NhsBqOz+VVa7GU8sax41YH2Oq7hkQRrZd6g1R1txJc8qDW0epxwSr5a/1v9
zhmlEW7kCzoV+KMRGdlQRo3XbVH6QfsnbZXqOsGzdOr+UFpMzUdovGgMi8gWWFmX
kg4d2poHYE5/rwZqytYLVXcDbOmEL1WiD8SQfEGnjzBjqt6Nm/imbK/P4g0b/tEn
eL6OdwhgdB0hL/wvAgPkWi3RjAx8JEv457FXIlCXlMr5lOUCVf8rm8HqAz0CSpcx
637/N7Yn2+bZ7/yEt/G9JRMB90KTUhlJsOL9rD0kRhMQ5D4kruqngj05tbNpbTZo
CiycEe/RL8D11Uf/zQBCKG6/HGj8Uy5qq5gOx27Wlnq6HAPZH2vDV4DsMYaH4GjK
ZBG/nkfadb+Qo6g6wYG8OByKsdRquO/A3WHEX1ycAwlrCQXOlBg1vM4caryYr7yy
laQzdsWT//wotGkW05MDi0NOhy9Pn9b507tIHmBPWkf9PliDFgIVwcjI4txFMplX
5R4xRjUrorOK37Pd2PYY1AwJCDFc3AAv/8pv26rM10XkRJaQS8rEzvrJ1JnERHpd
vSbxuBQPPw5dPoA1L07wuKA0SKd+Xjp1lDl6+S+fB9gTx0VjlJkxl7tM6aQLH3qy
HSIxS8ohCTweauCg+7bpA2QW99UuVcFNlOpGIPwGEE6z+xoe+vqIzPx+w5f3rQfb
MjDuR7E+NtaLVLeOpJgoAM1HPhsHRfSAyWJ3/1Bu74z2xtJRqTu728mIRLhcUm0/
VOdK++Yvo/XvaIY/ThXslzFyuOITQ3WTCcO/dId+G1VpQUo8LvxJAPLeY+cqrzks
fFz00zpj148/IJCCnEvESf5L6hb7u+AcAC4deYm2Tf6nhKVcV81r9E1/HJKNTGia
1MqqKpmk1WCf0iySRfUsv1jSAzQyyNdl4pmDNMtMMg81GKL2V3Lm94hxT7wapXB6
RK0Q3VPlC9MqAFM1ipBl3uN1ufNv+q5w0SVWYn+lz5d1Y71ajjpb9DjS+UfYIKha
KY3ee6rX8rnRSZf2urXkTQYa3AiYat0MfiSy/Dd0YWs+me0DJ4j33rL3BRAf+KsR
CkOBeFlPpu6vCMGX9RprwBfqYAIHmTilZpV9YAc9adNYHll5hRSLshhFNGXBzSwN
V2Ow1H8nhIbMbVu+3+q1xCmZK/v+JbmvP3efscaw74RakGlV4ZQJuI8Gf70yydKc
Ii0ZdcXdnr/4Gym6plmhIq6X9HxWms02jPJJ2RmPDXa3i0uoInVB3prJmf5MVr1D
MxUXO+Cn6lTDQL7Y1eP+y+ak3YbHQGAD+gp7AWltNDzQYzp/tLgmpVgaODZSBwN4
SnkbCUUx0gSlFB8Wvotyir44oPLFI3VFZo5j0exmCctq/ozZsoUwaJwFQPKUWltU
U147h7pVXXmwtobuSP7H0LuyYvJsA2tLmeiVqNq7QD/pmlqW/fAgnX7QUmvGH/WR
aubZmc+ZYr2EKztrBt3SiOc/DMgnuMk88khyGXXFjealsu7ZdZro554QTufcvNBu
7KlqIZgLLCgZpq+1E48yzGhRxdCx1Wcd/jf0KOh6Wpvqpd/XbnB9wHh7JDJDtFTo
+hMkB1/WSHogE1LvFaQT4twQoLrSwqNMC3n3Mtik0VZdoY2wt+SFc4Ol9qqORulJ
N9/yUY4ExqB/OI9QndBXuga7UYlj3rP0iNSP6AWSsIFlj2VUwIfLXJhwLdyLSbKX
1/nSKJeNPh4jm3q3YBLG//UBdHRrUKlO58QmU0AGk5MUCAhbNLO708B0lxCLcAi6
+gs4AXcMkoacrNgkf8Y1qGNQSV+K/XrQ7UXbafk3HlkCZd+PJnX9uvLd9zZplqwq
HZP4YeIh/by5bAO38GC3c6g5LwIKNE+iDy2yefnm0FvFWUeQlt2rd49RQ81C5SNd
MQk0RoDL8fQpGAxQ61elnRTYQkbBotpAWAO49fFdvWaLu4xbdyISsSIWm4N4Uog2
MZf5oQ35W38J2gkLiooqY7Z0NQlNcmcu9tw/SdBs0s3L078BHH/evbVsnW8AHJvN
clbEQlh3+TtICZuE8iSYgBZnIkdtJ3sBdISwq2iKsybcYrYmlHPmjFQmZNWHfnNk
hDtzzlrw5BcpKuCAhCWgJM678TCLm9lbewl98FmyXon5VK40DSHxcsovHAV2E6Eg
Jg2KnBQJ4wrZKatFysXxw8UNG/cz9QPUqPspG3ERwr/IhgHKqmiL7/g4Urb0HrTk
siuR8cEsxxPdlDuyMASoM7+ufAtpJxNqqYEJhSLfEgBAdyDbFtQWKa9Nap0BfOiQ
DdvYVnSXgiqIRTT7Kv1Xo9QMigKEkMxQRdqedXLmqK5y8OG1LLMdAgMGaUIan/Av
DY9IYiOTlo5SSHQvZE7fCTHt3PLr3sTd4D4Jy5LAZuGilUX+sA5CZ/3yRweEd3kz
c0JDC77VMG5/Nq2fKv7DUowI2PxyZ4aDf7RwYP1oiFSShCibg0yVITdZKBN1+Jtt
ZRTjl6UVO2PW2NXrwtz4JWSMSOqCer0A3b5Tsu3X5Q1C1ApdFMBtXKxSrM0+cByG
TZ6j0bahuccihn9ZOB+VSkyE/5u42QrjUjeTim9eCeerVsFvqum/gC9vdvbF1qCu
1a2o8kdULUS13oXd9G/Ow3cf5ME6IF7AwUDt0AFeRH2lmpiyWO2uyPi52XxkRrIf
QRaAuwhSeKZn0sFDtz0Dy51Sawg/2OfhEN3whvIIA2Ti8z4pQpJanW3sH8qJW/RU
vlAZJwkrmYahT9hownhnJosLs0JfWZLyABUlUXy3fY4twrEEUBIcQdBapMpogVYM
SlTJ1JrgkGmIp5VrMXGYYy6n2IooVyFfYYBZ/6hL6m6xSWSp80VwaCjmJ6Q48fu8
SvApLWlUFWxCQmWRZmTYMJZAvfr3RKScw/V2NYFKyWU6wvqISlrSXZXLUTILBd9Z
71u0nfbKyf25hmhqxAhwcOMZaetoMcIUkmGx8CSujMfDEDmelrtbjQGUDbEDiYC/
AuOXxWoRYXeXAVMb37f96th/r3gr8BMyRUPoSAMdwGppgOLPF+Gi/UGb8ZC2qPVh
GCG3601U1BjouEjQdr/mtRsMSk6PnjkEptLxSOXAQgIO5OfkBRZp27C+j6Znak1v
ZCEQi7BtOYukfdfnCZJRJ1N4ah0kcf85EkGxQtKx9JAYXW7TF5pkOjyRoZ4tDhHF
AS++2X8muOP+oAORx0jY5J4RIjn7ys66BzKEpp/r5fWjVstH1yMovkKj6eiXot2n
3nu7Wp/zufKJFB+dxvDVBd7TzSIXGPg81bAfIr+0pkj9RqpsF7+bmJGcBbDktqZI
B5XVug9VMFcGFzBVhmoj7sdJLo3BXvXmjyzkwVRKyX0TU/ZRF7j8LBXEOJn6r3Df
ZA0+L+vpD0v++7vSgWBb5vUk8oYvpPpxfjaWNb/6XI8nl+P2dHx3Zkeo/WMgnxnY
3b4PbuflgCCuh+KwI4VC8UyL1gKxjnHWHCBD7iDrRqgwUhFcWATZTS3Vq3uh3xkb
Y+nx1VV/WSeUJwrj8X7EZJCoMdq9sq58ulj39pm/C/lNqm3p3v2DsfCm42jrvx5M
9Lhw0FmXpwGL8Fy2CXP1O4/FK9B1dOisejBqRLg9+6vcDa7v6bhtIgE9jTEF5T5+
t+MVAIhnF4/CRBLVWDdGIqRH9GHqoTM0W46yfuGNF1NcjV6zZrXSSQUJn6RR++xk
ykfPC1GdVh1EmiFSBljwNes8x0I3BCw19yzfiVAovEvaupdMJSEdcBDHSV2VpvJc
D67NAlMHBuvSdDGs2APk6PdygjjNmayNZGtNF6B8nDgLry6b7WcJU8q0RnScAMFy
nuawRxu+Xx0hQ0Iq+mYQFkY7fbBw8YMa38HolsIgmlXSwJbzT/BKiwSfJpzsBnMw
sUDzkAFZ9yw/BEsBgAEutc6FUMxgHOTXwkI5l0xfCjKywm7sCqotmXFVJoBZUBwY
gb5VxjYH929rRJT3Ry1Lu3lXyZz59SCxONTRuqMy/NdtQ2MvdUafJAtseex/N9zK
LU3HQ4Msai5NQrv4MBl2yVj+0JFLomaZ5nmGxiSUJGuwF4R6Ohup7Ozs7TegYAyZ
0BoaFJP4ZBOmBEnTnrjPcaEeY1v2pdlj2lKofK+okQoOjEJZwp/22lOaf/L/91TA
RH/AO8yMSxB2MaNKnDS98jtFLh3IJT6+BQp824VsTJO1ag3ak8WdHsvIdhzQHFnp
nOOutj41N1o7uHpYjWBbnvcK/Z1RliaH2/eDpdsFjOAj4myoj+btXuPBTfNqe2pF
utYTCN1/gn3zdC+rESKi2cz+l+HER4hKU2cUn+cc7RoXUKt/V6uq+6nkxxfG7cFX
96V0cXRaTNGi/tY4Z4peofV3/ET7rfDYZZ2lgr5QCiXTCUfp+QMAlNp5png00FgR
/dJ2lPjpMBn5eikXs7hBULcBdrPtbjcTdgYXyR2chjQzt8fTNKoOvoGdAES4v875
fCuZaMZL3FnnIZYYY34L7/vYy/aXtWs94VJK8q2r/I8FWm8ND48AR5pJ4pNPQXPj
YeJTTTkFmhQvxBM1osERzdjo5bCw9Xl3BaPV3XHaXQclHeGybafKjVxe/FjWMU7z
73qAT6gcvRA0cFdbtrRKZfzAavqOs1Nmg2sBJJ1HQ+OcORHkz6zx1ay0Cl5rKaQ6
X5wlpDJtt6T4KwpbelWNPc45dWyU6Rr60DdvX3Aj64lklE08viTONR+51zKGho6t
bXXhSx1MEQgFfUDG70qPsFtQxhDp8TvyEm6QA+25oBLa44f7XlCBDnXgixdb5T3s
o91wgkxOvGVeukk95HUx6erG8MeripNkYklRm+ESVvObjVsdiT7HP7lNClVi2BZX
J7erQlCz21E98Qtp+yRhG0Lt069NAPb5WAlZGGgZiOR57+tn5f4OtfdzoUXH7OdX
JT16hECO8jYQj9qCvzL+Q4C3sEZhwD1eymW9gl4dybx5Bok2ciYyAU+FO4TR4PWV
eWWT9OQ3AUdBIj7te3Cjqvd3ntx6ck0SWWvkmAu80l4Clt2jaf78+o5GFkN/omHH
6bQv2TQjwWOwoeSl+nCwks9ldqbzUOTZsYI6cmgkuSP8jt4yEDnwPt8VTu6URXc7
q6Lsw+ZN3hCMn4lRzWQNTL8iRLSDygJnqYnq+mrc3+YEWX7srJtabPBOqZoILKa8
2sVLJGjyTbQ3dKHz9iHgOFr7wZzexJFdJnkM/s9JylQp6cVM21vqtyUrQOUe8zfT
ZSjei0UfnU8u4HmP3o23HchV1TkXCdAeFUy3fsV0BrN7xHqURTffNhlXASas1Iw8
7MSyaKqGyYrBCWhxHL6+olhDGNnlzuMQ2pd+kl3o0GqIwGFPIUp8mSq5UVXApIDJ
aiwpLR0WQmKFGBmY2FAXmpq/gUp4tMm57kjVwmwbex2EBuEGZ6v+oEFyVfeVMO1x
UNZpP4+g+YzM8rdtechV0+hIyZT2aDWaAFcRg3zT670VeWjzS3J4snuEGqxU6gt8
ZXj1SBpPNJZdL8hUO0s1lW8uqtXdkmbsdCZ101OlcO5J8gJdzUP6WB4hwSSAriMO
lZPe/+0Tlf0Lsn74WWVrbv631QROQz6mTbCkQUJr3i3jeRikCr37jXpE7l5JXmAf
G6JQdfblzUUDHjGQJJgpRtmQ9yEtliRkq6wLcMF8zxWZBdRBgxFgOXNRB0Qm/j9q
Xyz4lMgyRDf6rek09moiGPYcJosCd8q2fKc3rJnvpg5gVjaKHYGWIhaC58sWqDEo
SddHk/XfychHRacbhMkDQW1T+UWkWwMPIOcJRAEsYN0GaCavQ4fs9eJAAk/qWqcB
0h+dLXF+ItvNtikO/RqIKqY7RxZXFb4VjkxuH8ts4NNv2iRsWpn0BvF6q9VCRZ2F
GTbs/zJjnWbA3c8Zsm74Spim1Wznr0Od/JgOMS2y4coWD2bBULP16cApIQX4PKsA
XQ9jYffBtVBwfiG/bPcbQ/S5w01IPG/bA+1eGf/epKnxqeG8Naui7nwJcTA3Sars
3weBY4zEDnZZXsXg/gBIdG6u4Cc6GghptlbFbQieJKYW+svGhPW5I/LBZ4h8WU/l
OGXFEkA9bdROc9RLSJZLMc1NgTMBH5L3yIt9+Q2sHQDVdM439m1UpAA+WwKAKOoA
QfL//c7oHFqpdUst9ogfCO9lWigUC0QYZToTG3eAah3SYs+kL0y+gaRkowxgJC5S
7QeS/clRS+tvTVCE7g+BG/mAfLrEWTPFbWHWrJ7rwdM7NtBOCatllO0RPmcWQtZD
an7T/Jd8kxNa/7BVgRYKLbNNaQV503CqXJmdrAcejTMTAXFgE6+gxbmdnsaX+mQf
wrRtmaB7ItmwUVptN0Z0FlE9stEzU8xl57piRSRBK68ml+UrNHovE4oloncLX4AG
4sZnjELC0QyhSSXuRvyYBCqn1f9ouuZjWtHrJ4ka9fxONdMLzG041WhCCLZIkoXb
celZeRlX6rdy3Idwz2IT5/ahgHenhkUfWZ8UrKfciR73DI1MCpcopX6v+Vw72EDG
7Wo1AHAWnix0sgiAptVw0LernXnuslrsjTv7qQoF8iew+YL5hap5cbxRMLjtrnXQ
Sk8iuYx1xQVLTTIVbitYZq1QE05S80D1horgm80ELBo39Habq/N/7C4nGUfwoXrC
+wQQyvQJMhYMGUHcnRZhhzLvDlmK2C+zhW3PGlef4ybjJz8WpEPxfYbhvxpP2OMv
uMb7evMZO9C37ZwGDorscCNVwvsgx8Meq8+Lpvki2SFe8S7KcXzS+1lgPR47GfK0
V6SGNA1DzPftwwwz/Czw1d5cas6G9qq9hJR8l9sYofyEv7gy6ACwytue9zzM+NBz
dqJh1wOk3GRyk7c8ACuY4rvYagQzRYO1bIACQEuqummKzq/+5Yq2CTqbhuh9AzKL
I7fTdYCGh9/8v54gQK1dpGU/UANncf53k8/6BFItOmxcenqr+vr0r7N6K2CMzd81
sJIxjY6hHhsJOQz2ri1Qhj+4heJvVR0sekDBZQ/cwqglCsxnRszt0rYF4iptVGh0
44r4gtbS5yu40iuUndqN7jeRmVr4Wyy/cet5QgzOm22tePNfQXKAm9dp1B4BKxIF
WiJ4FWyV4Jo8ELL6OIXUBNLNLu92Jo3tqz984vp2Yc7adbSRHZzfChZsvRkASFCn
36SclvKacDnN7QcZ3lex1wuOcYLqkLgdzT97AnJAisB5PUeKpUvyQ0U1tOU8ylgn
QYwpdLls+hjNNUIZX371Y43NgBxSrwX/PoblG0cQmyoC3bWI5XCflxMN79C3+AkR
8Yj4/U6BcabSeEViEdlua3asLsFn8LKZjozhIH0YjO2IsT/p0s117xB/wQ6Pmt/9
5UHb2ELsRtBkibH9Fdqq7Zyfwu3VHtf/QlXMPfcBz4YJQksSNzDBk+FY4xkNYzcC
ghYWidH0i3huB1dlBr028IEkSwfYF79cN8ZNYhcZXmuz5LOsvBADBhBhM/ppoKD7
C/89Mi3q0tMnDZdHNDuDEflqdR8kSlBI9BoIH6lbONeeF4f+2GALr86L+/oGHURI
jlu/LD/oRuFL/niA2oDhPCdtBmeyQBf7YNjgY6F5JU0/KADypjlLRBdZ4KNFqlPq
p5EUaaU3Mp+3zGe0PxqmMmNsoe+gEdualruulghPzSbEEW3yn/ohYAz7dq1Z60+o
/AwzlNe6aJJG0DVnQ1pAN1QhnQvBrNlYTkvC7sYmzvsDtnqxHqfLU5yB2E6PAhM5
lNS/o1H9GzH2orhOD25JbivZTTo49mQQxUJgdAEj3ow0CWxahqFd0JQWJQd8S/7Z
Ixpffd53FlXBLngKkLSls27YSWrjQiJiGQG2UUblhbO83n5B21vxWhK0uKjpPCHI
Phlmj526YPUf81IqlBRoryQQOQHSzAm0EiSvYFEREWeQQsXSxWT3clzlIWP9lMY6
/fXBCyRtI/dw4kszcJ1R2ReqNinJGwFYLkiR5su23wA/L8IY1rtEPEmpRy2/OevU
fwf6Iz1/swKf8GJT9FARXj0NqPBe87k/enEbw5EhvH+4EqRNN4uVRKiCybKNrAcL
v+xwMtArhlZCrTnD3W0xZvpPCdYD1u0Ot4f2+zF9Ec4JwLNYseaztz48mrqYPgX6
x4b4+L8AILV0WsMcuEx5dHlgYP8Co8fYKDDLl2uz2VJ0IpvjeN53sdc5WyLdN84j
6i6cNWSChoSvCO2pMW6zLGYRnFWLz+CUkRx5wpfsMKtwJxInatU9qrezIuJSkh/C
UF4C0IJV3lUottMPDZwkwsYz2eoCdetU+4KLqK915SRlDBAz1YyeNaSk7V+TNC1+
eLaWqXfecWDHptL0kfI1hLE0+zzKcE8rR9s0SAiA9X0vizhK5LlAYsK2khsupC4Q
3nWwqhs/P7AdKHMOlPZjApwKb7N0RaDQqx0hYfYn72frZg5nuG6CyS5UjtguX96e
/AHc6A3eEjGGS9K0r0uGOHMWLu/gXE8TOlPWYokvi+BQ8DBGY9eDNJhvb+yDvRWd
ywFdSmzHTUpMQni3xEseaCVPxa2VozqcpE6qLAbH5bDK4hOgIFdE+uLKNRAoyrBH
MTjaCcwVHMXlfrbbEE5YqebGad4DbYmC0yrm3/FOY4Oys3q+8Cfvy6wMNmVAiPkd
r6hiLEJpTcjhTWuEWv59UNiALRVRofonSAa6Kh8yv14fK8q0HWemyYMSBlh43nH4
602Y8TsmigCxqCRemlgtlm8UvWj7vh1jK9r+mHVB9Q1tGQtCK3zCGqixH9Cd8LoC
OUZNsOrG8iV9CTGshP2/093aJIcjfUk0FBBe5SL+bYiao2umXXbJvj8ve7G1uWJw
Mrhk3xd/8I7Gk1v6xVns8y+3sdFnFs1xBO8Kg5Sv6h3JrGiun2WqBOaASdSzkpzp
KgeCx29AHj7rUEYlaPrGRSrHulGmcmJIclQ4iiTbD0fMOexkJgLmfQBq+1R/lqvp
tttsCcIC5b7+7MDVt1uEbkyHSJJ7IbUA2ew7AP7mjX3BYJgqikQUSl8vId63ap/5
S+Sjb/Rwv9tL9tZZyuDyUiqchAf/Pi2x017R6xCZ+ZEvRThExYCiixkqdVFLoGRg
/gd6jxAgQoIy+HNwujilU0C9fROMCktLa3jrY2A+9MmisOokiV/+oLTMhJJQghbY
MV5H+NUs87y+wi4Vun9zEegdFquYSQJN77SfrcTzTbi/dGBv8YmRsHeCw9IFPpQl
Uq9KE9Limma+Rsu8yseyQc3os18mzUp4V2EvJfB9fL+T5Wbpdpn7Bf5LiwEGXZrN
QykAYRBs7PWdcXz8pbSrwDi7c8m/whQCZCNppxRAa8Hznq3RRhsAe/AGmChJtFXS
3uAn7DK2xwl5ZzkS0EL2YPJX6mAi3e3R5/gbUfSjrcIMgChkXLOa5g+VrTMi94Tv
sNZoNBohXrJ+xz05FKlmoXYz3a61bXGriMhCQAgIB5QsdYZ7A26Ud9CVKMndCY62
nCzZ81ydstgQ3q7HRicgpE+Fi3fAw7jEHqnnJPJmygNju9ojn99XiD9bckBfbHeD
rhbZQz0qDLI/7WnFiv8eoThXVB7G6XQYKPXHj8NukBSwXmdFvemHR2uVY2UaXTfv
vAf6lPMqOjt9eXQ2kce6juL9twOghyjmjQq2Yr3YiQkdlKjgKdi7XXTDVCczJC8d
JFwaforlVJg+VtFVH2NHoWVOEghDFT4eGq8k46AQ4g5IX2LE/EC+ABkFEUi97Eza
NHBBgo0/HYM9eB3OH4L1fChMO8wBGaJxPEyGPe0un2ze5AE5BJYvT0OxvzDr/TWQ
fvinUtEzj2dib6j6dOdf8iUTKiVnZ1Vv3+/Xk8zV6OAxQSaoiIe1/B/tW0JCbLUZ
izFulJQG9XKEFjIMsJYgtO4YXqWXAoSbJDO1XHOBo7Va4mwonFo2ZCR71+Zqjyxw
IDq/vUJzHbNAeTevHBViTh2z786/Z9OKqXNnXj3t2GVSFXlc7uEtNV0zGLI1c01X
bECi25gHbrHon9ix4DY1JHTXPnJvqROPOobbuDhS43m4nDij8E6lw3BrxBU/Xwl5
gNCZbgyLZU83Dt6FAozP58QZjk0E6ggoSEvVB8RRjM2fTNAlGF9uuAKa5M/AGcDb
MuY8CLJX/dB5e4W6QrE/NgGCfTsGtBmHST2uWbpu0qk6oLoIGkp3/aU+u324vtn6
J9s+8eimqDch5ZKx6ZeNq+3+cLVa24c4VGqTM79RJe7fCCZwzQPi7ElGpkfkjQFl
EcBNpCoDpoWw9GFYOKrdXZBxBUSGwS9ZB2fleZ2KO/bhCXJODTlA8/YhvPIm+Flu
jhVX+99K4eOMWDXErfC9dntLTqkifUKI5MImMAt215MEJXJkBPdl0iCx3dF4z7ML
5TSdPYNcVocvp5sV8s4v1mDg//JLK/9rK+hcQqEbx+T7qHrZJnzeRwFsInugfggp
PS1jK2FP7G6qqJVYQTXoZADGzOIXU7d8vujPnQqu+D6Zi8JGeZZGBwXsVlvdWzSW
LDWE75X0jmmSiHWIPi3HDRe5tMBGzbmscd512VTdgn3Vv2WPMX/iiVZ8T4kNlxiS
UHDAVBrW97UEY5iVCueDkVWJUwVQ9G6qtUmIF8A6qQlsX7vKE8NZhsqQsHX3x0Rv
Q5ysSHzIgy1ZYJVxrdfzB/pBFA0F91+Xvykztq2ULCcKBmx4TF1CktohRyRoG87U
O9K0r72FSUhXtnwylVfvx2u69w0tU+RRSkaVF9cKbfUDWZSwLN54xYeK3QjV9W61
Ri9tasZtbV5h8EaM/9/k4C38GH3lwDsXt32nlJH8G9GCZGfVE9TemFYV1/RhORg3
Eiid0tDCSxnvoqfwzn+8GMn3DKdWc0j6XJj1R48m2p2EoB4ZNWc/6K+Gc1PTIjBv
Php/Ewhw+kNGeFN1IzoQts+COg1L5nODp+qm7JY0g4jAfPrGCeO/Atvs7sk/5fk+
XP7phfzakwuathFZpqgRAXobptTRq/DRwY9GNOiJV/b0ir4zctGuz9lcaVd+Yvsf
sSmVq1HZooJPd2OO/8gOdJ1iG9uoAlO+5+kks8o+XVt9ETFBNZ0PDGx631kRGTli
usv1gdwFoiq91n2Yh2XMmxPQFlB63LB8cAoM6Tyvv9DknN+RqlzO6o7Y5LBERSIG
+8oQOPEnLgwWPErIMEczIr8Qaq6bLrfoJKOoiO4G1tkN30QReCv1DNQWCjnMxZib
rKLKcBcllpOojlJuvo16kHLAafVwYfs+PKvis5p4m9Jpgl3q56gLwu7d1tQjFPor
cQLLA+HzqWqme1CTKTf4a4XTAtt7Ji1SKSJmF+zduAf7vzwQrzkJjQJmWLDG8TiS
TQNSSDLQHRrMieliUiXEl/SqGvEYNcuLHLUErmydjfLJWmzd/Gfmt++NXtpVr86f
gQm8ygIPEyhcDVVZjtuO7Vu+n7pXm6bTZprZLLoGukV9coxQDu9qCrAKo6tZJJeu
fGcqw4G4fyjiJ/XVV4I3zVcZKNyyAP6m0DZcZreml5nVje0ggFbCONtRv4c3OhlL
ENqeTJznfsv2xwa3j2geVWBbzszSu5j3E2f4AFZahcdLWTlAgMHGQBn7momvof2A
6h5Aay0ii3yjw/MzEb8oVYw1msU7RhM4n2qa9QeklppzSQHb/S5K55Vg9dUoHRZv
YoAjRe/VoGkpfAoLcZM9fqX8mFItQc0QSWDPp2mO74C/GINRWMAU0QjcdkaDRCdS
i6ebyF9c+D7M5enrPfDWrvuMmYMU0OfwMSIhPSL8ivxnkZD9/HVJZJaF8uu+sw6t
sMcezlpzKRgYy/qrJ2ODgA/aZ8gsZwRT78ZVROb70s2LiMdl6+iSny429nwKv5Oe
msG1g+DAjTLKWfATQ9gC+LJkrrxWqvA22rw36dey83fJXf2k3XO/fkwVTx1DAlt3
BAZRGYW15qkS6CxvSJvCacRbQZhv7W8lER1kLRNaxphucMoqZQ1kuTP9L5jjmbZn
D/sMDd3+KDamn4smiIrmfAP7y1kTDnTmV1+sUiQa6RaFYzhS6pPFu8Fv0kBXzcOi
nmTmNYSZ67WUTVP4EtwGm59ncZB5HchSj/w7OACpiW1zFyLycmT6oxZStDRqfsns
zUukN9atbP8gR7jIMR5HAXLNmaRxjMiXzYYu5DXi1syolAiTTEZFNjAj+1vjbChJ
7qzbSSQmF0SL+It7V7zFiu3NZ88Wgv08QAQFgF1+peGWjqZHbu1QMzXzWBmMDnLM
O9wAJrjv9xprw6RkvE/3dC1jKQIyUunlCrTT40+G2y1m8hJJ9G0bGlBaWCfrp+hC
SIwF2KWEBVRY9VZVkYQ837qmSoXKlg8GQVLaLOfgAear2IO2IL1p9do5ByhuZI+Q
r4673UCYZ+Jo8vOGeJ9kuARCpwxnvID45O/5HugUCjieOeVgkd7huel7D5nvYp/a
5NC34Pic9hUlG5H0riY/eebUXVmb4+9Xas0+ix/CreFSh9TnDzUxU/9jSbTKfftI
F0LCx6/AXUVXqQddtRqvj3CTWCv33V4ZJHrlQ+OMhf7y0ZEeo8iGf0QVuV6sgXwe
dNI71XjgIziSXT39DwbbEdfc8OZtguo1iCwclhXReV3jNJELrNEvspPcQY0n9Psc
lR1ZEuvlKG8efwVvdwFk7+MPQIRgdNxbkS/La25U8cuC5AmhRXipQ+819p8aitKT
Mjtl67bdTzMYj2Pk4MH/6t5iifaLbmJ4z6Oksa84+qhfyma/Won/bm/acneEcxJu
ZmUYJcsEXqHR9O0KRaaNHgreNncIaoz//GlmQy6R+YZazbKh7udrY/F0bPDxs2dR
3hfRlv/xDFlZr3rzX1OGvd6z2aesNJlUQ6wf04XTnFYDLxQ0jNejSZbGB8xxHZLD
eKASgLytw4Pxj/d4MW7fFQqRj6EjKrojemvL6y3CwsMo+xUnbPJTTFKHyVDyy4Dn
uO6OBxcACL9IR8eNb+IDAu7hICncCKvy7E1GDM80HEcS5Ah7Y41TvCv69wp6jUFF
YJKANNVtGXaQOXXC3oJd+Naz4uaXsAVt/+XONczTa+7J1yIh+n8jhieWmZoIpidM
PaimJ7jddNnxWBoF8QN0qYTQ5spamVx3ibwLdRdieJcpdjQkFnCknsnZ1PWl4iSV
OmPhmDQqdrnjV021kLadBxdBgFGZpGnG8Tbl5+bHIBiFke/xQ1dDZHb97oGmCh0J
ssrNQ1NXZeptUkIilAWGWbveeOKDEQiSantV/a46OmjGEZwje5NgZcwSvjJtc+JV
QyimTOBBB4KJVRtr2Td+GvTlUP6OW9/K0bVELv2uZrwDnB0LZS7OfItNqAMK2One
gZph0byb0LMsLkIvCy9yJs8/o3f3c7A4OWhrPs9iOTpDMNKJaAw9nK1CJAvbq32K
peEknlzm75VBSBItHhGiyq2fGlx51ajEo+1Mz91rN/Qgq9lUAh2lg/Oh1YSqWoD5
BOJf86eY0XYUyjXSjZ63Bo8KlCJC1dstuphL3dIrS+RLYVLZqhGar9AVz1DH5S5+
jJzYhOUZf8tJ6tDG1DHHeu1S05Z4W4xqj2vxJHSV1Yr0yCvdaO5jmnMNbUmQnnV8
VJL9WlS9UU3BnzxrlQF8ojaxkkXT2kc5OFQ63aD0bFtJnw4hXzfLgF9dCFBm96Pj
zt65n7I9xLBLDAOLcHenKycKgJGphNzD09y2H6L+sp8VHP/EvQoRyjjIof3p7xbk
CPU3Q3f4aLA2WtMJK4uSYQvoiyojKIE6eHLIMrWkOo29ICErjkzWn+feEKT++GF8
YVXjkh9HPFDYvnVHKF2s3rvQVEuRDATqSsMLlX+dDSjQlsc+6XIxBogZdggRCPSZ
W+1fqzZxjxW0/bvBax3EqbNwGTSqagQRwzZ7ysnNLCGzipXVP40FZ9WM5nfid3BO
qbLKGnC1cKBbD7o1CG1x3eKjahNtx+Ek56clCvza5lmkR+s6iICBdQloiwi3LnZp
V3/QwqcqkNd92JUMkIL5GVc68cqijm8nrHAOeRzf+e4BxSNKrvd0OIIvwWPK00Rb
QG6rV7oxzRrRNEq/WetCggHR5o1oLfyrQkIt6ggodUgcDSii3C7Qq1+qiIpSQGSJ
fbN5JK5Rlsfd/GcP6aLCdU8vbyro8PSF8v+Arwg+gGOQQALsxGpuWcO7+5Px7IW4
ETZvnxrRzyFjEgi+x8Z3b8ZC77pWLOGb0eiJgCDGeTTAc/3ln0hXJx79C+KkJE6+
0C0H4Ds6Qc2xhYfjdJ3cNivGw2qhF7W+rEkd+FP9hTVYXkUrYHS2HWudMBawKFqw
VQBgR5LiLVrGSfgot9MmoQRkYvocQMhwor1XG5bewUc/QctYMAgh37ukS7cUtcwE
LWRSA2RAA7jR/dgTSxXMEn4yC3lIXf1P8MM0WbQNyWR58Gv+fHEngduX8CxMTYDJ
Jd0hWnFESu8siJVM9zIqNFaffzTVSiPonawy+EQ4hTKmEdJMiP69fE2GhNLSt0Ye
Kz9uXW+aJ+uNr5MTKR0SIa2/HYXlToW3U6ljNh9jO4ePuoASqYXrOX0e5stiRvhK
QOwD+w0j2nOcvLz7Sov+1gj74sQXe0G9+sAbxSv/KYOQ++H77rS4y3OxDtjY0PNK
CAxgiX00DIgozVStc7bemaIZalDdC/WvUDM8OsS9f5IHje3555CneV3HTtnOf1ED
gy7LIub6RpTOrUfn/yLVyvGpaFFw/z5mYrTbMPX6tJZfZ1pNyL4EyU/0J+d6vGFt
RRIwA0SpSwd5tZkGWigiw6vWPIW0oacmVXhy+i5Zn9IP6KRlz+eIaM/KV4Py7d1g
Jc7MMHomWYxEdTWbHpw/tgeD0t2XdYz0uCOjipbAlzZPSPrDBentj+6aMmm+iHBH
hJL1kD9hSBzvUNry5uWlR1Vjcxw2D8vzKbXvAAo1V2/pCXou2X7+OYN/1wAmoBaq
duvt3OQc0gqLGuLkqdVljy06VXXe+Adq+nb8VxuFv4AJasjIDfL1+3ysSCfIc2US
E3zf0OvLKdQ1R1mg6cgcBzeecbcnX0m0+2ZRn4DuRMjZun/TVsHH4XLNM10mKmw9
ME50BuDtPPuWc2+glk1GAXZyugokwohQwDEX2xLnzGI7e6vmQwx4LugDllbUbNXt
urvIsCSYAfMDtILpTgzYSuCUN28A4644PeXtAGdTozpbvfqfKX5vWlpDbbhyrvyO
zDO2hLvyFbwKtR7J8HUxbkUl8jBWlBREluBQE5fRoK5c9Jh1iDdISBOVk0wkgmIv
nb7LqQXEZiG3cV0xT7TRSg0XSxTDPylP2tO95MIAN88dp39ia8BhJmOmBjpNJrnl
uWTuOdpmWChNFJW7YdCAGSUrBZLkmpGRIU3D2+4HmsZTC4YoR3b4IKC4cr40GrDb
OkbW7jOh72v8a+sezqPR0ocTfdbyWtl8QE5JVSfKswvh/SM3ZNLaBrER59K5mKWD
7t9TbUzICwD9tZaGSbtEADrfLxcT9ASn/3WaB3Uu9hctsUYPR83JOhM1WkS0SMFa
47vZPSiKQFhlY1KhOrKJrW/qXuq3BfTcvl8RhYj8MITQyEFTXuGA6if10+vAvpsr
Q/F9A0kJZ4iOhD/U7t5OL0M8Qf7DQrERszx3pA7A5t5jL961urqyqozZ1L+OGIVU
E+nonv2lII8ke9R+U5sgY+6xQRGoEc6uyPu+e37T5P73/0kvPdkr4Fh0nlgtiU4P
gNK51gxbVcVR9TbDcEGYZ6bU0rgQp6biWNJWV8SgW3Lrb17p0aaGEzu11188Upmc
eFYEAnRePi+9fHlWCXh1VXsUruB0tHncEthJJ/o8aCXgiGPBKj5fmcVEx3rnbvut
JJ+Hz+lWrnfZ6claSJgCAOqynZNdEpzv3tYQ9+Nx0NZEmPoCja44Xs/V3EDE5ph8
n6sGP4mmAqmaylw+gxwpjWGbnR1NlMliGzWqLsphpitnnArznpPSoGbnRpYolMZ5
gSBNvY/qOixJokE51Lsc7TrXHbn1U0GqURJUPFv6VZmeOOzw7soj/RcknfPxh6aP
Bqf+RWPnp5PajMIhs+9oya5Xi50D0LvMAyLij61ZRKq2r0gAjxFyteeEstqKlZRJ
EKQ+9RlPxdCK4RpMWIuYy+a3aNrrzd4psnd5GE3coe6Z1anJSVq/9WXjO+gNOFFo
xXCob4D2ZAUT7UySDxyvDBgMuYX/CoQWeB6Yis5dvtPoKeeEqOJPUHJQNEQrWbCf
A64ZkB8+9CbkGF9+zGnN2wfSYtU9Bo6MU0rKLqxnWVDuSFR3WRARhh9fr0w9oF4c
/8yM7Mcke+eFWCqmfrabOqM8s7uEIB0uSJ6bkXbKR9cghX1BEac4Xc0KW3Xecp3M
u4TaDSPqTnfNZA0SRVu/Zj8Z5MNKYd7cd5bOuGcW0sv/hEsB3I3zXXJvdk7t1yxJ
FMaPSmRbpm6OY0dqqTRWyIM5w3mm4D23RbYvMQLR5sRLDi67jADhdUAgrt7nYR9Y
zWzXHCtjhkRCBuC9aTN8r6CC/VMQ6I+GUnrGWIJ0waqsbDcunPLQ9xXxnczj65o/
LaEZcre6nffuagUk1Rx+I3KXZ3c2+EGzJhDl+Rvb6IcFAuolFuPW5uN0pfeXyVq1
mhjur8Z4AQ5U71Dvc/Mx05tw283sirtGZ9RlnZb814WvTeoMxosGDL0eMfvxeWJN
OXT3pzwJShae5ck3rIXTCBm999qhMUQynqCK5WGLuaAVfkwdplEBM8hbFTym+vhs
Wc8ci+fUjE9TyFlgTrgGz/gxQe19SY76fzKqbP2JDUJAIpRWzCBqvzKhennasZsF
bsD1WRN9zWIsUFTwHQBnlIE2eDV5FSJWPzub+pXMMi+nzZOe1JBlx/ZcF7dfk4nM
orACPnXUf0L6u/+VUO5B1nmsz1ktKmpvbCli3Lay+s+AeYXX30u7wnOSpyW4UfQ5
nJANEauViAxglF/odGmKSgbiqEiZW4zf7/ai1HWMNuodaeQbYfl6gHm7HQV/GRSN
CY29DRkZ+A58MiUzutQhfo/FinqPn6O2CJ1pDuxQHtKDKCkE0XHzUzaDqJjTgBIE
4zw+zzlkMdJHzFPjVzgDtkjifvX1A2E4JlRi09cZFzYC/Ourw50eXAFzZwmJFQSZ
eHvLAZcmFgYeAZdptKsJ/deRhTzrPxGwUA1Z5xeJwf4rj+eyAxxNpA5uOO7EXffx
YxkMAiViaqRE8ZoQLStaKys+VeiZ/iLJVRJaYUAc7kr/UKuIstPFl3gOdGv34bUf
WlCDPtfmb96bhjCH7z87CdagDKJOnf97cs2Wqn9v1JqjtZhBefz1vCgUgOjQeA2Y
pgiboKWpEVnLHuak1XD4rYeip6oVD9zncnKxpdPeCrKfxA74swjKc3fXTkX8z68r
citAe7hJhO0HLt+1zPvgnr6qo3DAye5smKOmA09PPZj8tfsaPqgE7r2KJPEE8uiV
ft0DjgyE8OY2k9vqsfUrzvRaMuxUA7Jnhwo/MWgoF7+sHUqbEdkIwhSKI5qlhIHQ
+XGR/qbnucKxVLhFOB68FiuW49Ko32XcryQQCPiHP6I2/3JD4tuZdPpZfoTT5ane
HNF3xG0RCY4UQx8xw+tTLm4j4xCm2DdNm7lFl+O0njDjk65AoF7HwuGLrPFZqKam
VXqCY71hE+d67Uc3SQ8inrHQHvNxA1jQ5KzD9nisNLibDZZR75zBE2LuMA3UdCHi
PV2Rmn0TydB7E4VmhXfeG4Gzq4p3QvTSeJkDduzKWiMaFgxrx2HvLrSxTtYQOnaw
P5jiS44YqM1AcF45knvQZSW8TmnJbxa2QMijrCErwS+fw2/8a0Wkn2uUINOpzCzK
Llr6S+5j1zpVZJ6bCpi0RBaWmyKbliwzy7cG5mdZJDUyqz5v8erTnV7Wmx6X/Vkr
gEG49IY2CBKXSRu16ab7Z0xV0vR5BUVhm3z2w8DED06S676OGxtw9O/ahB2t8XkN
4xUDRfiSiiRI+wZswrYtRs2UNpQFvahKvktLsnxUhpnGmpwMP/AWb6EkFExR7yXJ
0HJZyEv4Jdzf7Ouhmf1fsxoXA2v3wsBbna//RXsCpxLZ5hu3GozoUpNmTTgiiO1M
capk70AN6aDBoI5doaJKSyFApcPkRx5exF4k8zqFX9IVX6e6VoP0PFIxR4h12m09
Tl8ObPUT/qMlvaaRyPgZ9c7Fet5P3/3wRhCGVIwVTUqAX0qPNQdJRpahp+G+9NDr
/MrtMBMK5Y0E57MmY9LQ3foI3QujN3oddtHYJtiDeK7GdI4dMutWOLT4kJWwFwua
4atwY/EgCEBpgqAg0dKogIHasybl6ckdhqDv0lf5zYW6frmeV9wiYkfh2W7FyvHa
yXCQV/qTrX1NZDsEgph+WM31evqgmYZgZkmJfpMJBHNdnMA4oxFEMDrWhvGzDSZN
eNl5PlO5N93cXuacLwsLBHlKqAeTRbq4D1+Obp8AFIAmHsfAQnEJfZQSBbLHMt+J
BG+tqKFf7leway7Keiftz6Dd3x2BmTd/q+K3mzhqWhy4HmaMsoRm3GADtbiK1ofc
4WcwUt/jUUtgEr8fi4jZD/wJcJBLXDvoUdclo6+FwsmKgIun+bHtgPciXL2amCcN
3r/fBsLJRfyCqCzloxBk9uorkSPKaha9O7B/euMTsysyZx5OrCrzELGRY0kxwOn2
Y15cWBVR0lF/99Re4+yhtR+gq6VNdfqF2PU4cqzo/k/slPu7vYtf/7UjbNSxnPUo
dPTtJe0aoSORsTBSm52GHwnipU4AKdtTFKya0wdXk8WGZ4bcnjgUn8e1HVmcabQc
fxLTb+TRR0PYxG4gcSmU7GKbs9GgboOmzJUJ66cpj2J7l8uAyhnYbxZm6tbJ9hu6
wECX6ekagUa63OZEZrrJJnwQbBC1euHbsiFJGp7k1hXMVL+XmLGZEk02lWLMHQWm
6dLY1sM2QYX1c44KrGuB4lJAb8UWaeR2bmqyCTeg89xE8QjxqdHekQQSVU3o6DPz
zpxf1BmmwBl0W0QxMShFPFolCKCRf1Jj27SLa5akZ6jihW52UB2/Cfj327fiRrew
M0f3FDDoMKhLmNYIGusclXeHM0xpj5UnTOk41ZQ2dIw5h9th0LUsdlEWkl2spgKm
CofFSJkDCtva64EHFoCuNwzgUKEUoLXbVfl2g8vXn865Nk7stknLRatsEg5uqcZP
mirQHtlSG6uTUkC7Sqln7vIr1i3qQgE0taOydOb5SFgU40d5FeiNN5taZe2mrmlj
3VZW0LdFe/9J02cT/JKKZhg3BY3B0tOqD69pIZK3xzKUro/2cbP35ko2iOn4wd+t
iVfzXSTW5Oc2A8s+pUtWbTiwLLLUCrRp8hmWbUK/eJjqFAMiAS48zpo8EBkwVZjT
7p9ZBDWoWqYbWSdkvSZgUzKamSX79t94zFfQ0qn8TlnsZA9wNubiEcpiykBFgukS
V44LseNtspIY0c0J9ecoNOEYU7v59h9tvlw+sTOByYKAo/k22uXPq8RJYcvL65FQ
86Fo/DW1g/bme4/VR037lnX88xdG9bPGtW9gBgurk8s0Xsg32xu2QQykyGj2MyI0
LZsGQieiny4IrWMzGCLU3rPqukxpP/5JfzrKi1GP3UwwXg3SEfAI5yUEIQIIHwaX
yHqs0lWZfa58y0kY2UiVSsMgeV0E9qwXLBl9stBtCYKgKqjzWDB+zmg/BT+y2uI9
EZFNt0BKv4FrwZtgKHEgZLdscmWCknZwqqubbkr3omtp1MlqrfU1boowjSUc6WKg
02rdiYXDxcffLh/d1pSQtQG0WaF7sLOHUDkwKGggttyknvx2Hkt/sp0IvuRFC1w7
vYNWpiUzHTYJVCjvU8SDPIzTmSiM2fQNS9PemcF0uzL2yN7RR+M7s7W7lTL/g8xy
Q0StJCX30aVBwaHtEj2kZoIGVOf8kW3Dd3TejlAOiy+XMS68UE+46wMsJITwPYUK
yRIwaKPqisLAw4lWGBmWgHwYQOtFxEGFA1HFYK33WWfvbfyMO4DU8Y5jZYHqW1Ch
vX0Caqdv7L+82tA21XCczif3f0ZAfe51BNlcZypUWy8v4EPaP9oy10pX93UzFwHd
29RP8RJpUpTl+go7jWtw/58xCg+UWR6k6TeNMlKTlmqjKi4zoF3Kz0//xeA+oJjD
dqjnOTzP/IkoBKd+g65gTOWYr908XCOSRHpN+/+IvSguCU0Opq0ODvVxU+5hz+8g
aVmUNgTuaC29GX+XRk+Ep+ffTm5qp8Bc5s5CamOEMl13xF2TkysXA9/OIQ2KAZ7l
iCAn+UWU9anpRK3hVsZ7teePwBoAWrUb2s+nSZk5hplrV+BwV9xdR/6xuLLqrj2H
z9koVmPrkimJsq8bcODr0ofRQ/ppkXvRzseW8IZqUwpw/Ie1/koVluibvIijGEU5
/nuXMPUtW5Z+DZ/mNDUjgv12RjV8Z4On/elKqKqSp8ytln1dZezX/My81yHlsVnK
u9Oi54kLkhMrNcL8VgCtVP1AGnQSnrtfYKkZ0akgYRjl6oIee4HlhPijTy7ezWVe
f28MITGNVmY/S30oDREtBgJMhvglvbzCysDZqibbVp39HUpb6DSCec2e/9j9FXCZ
aWOH2YaHY2qYSedQVF4Jt3nrnz1/SI8l4UVG/VvuUFdsWxV/sQQTHMhMMujnAWeY
Mldy6DYN7Bf318IqHrIkhZgymNMkaLWbhk9Y50Vyz4jYl6Rr7nugCK2Vaob/e64W
RmEzKaJcno/7nPweFeLYa5Vda2DugJFDaHZ1WHZuwBAz3gDAoW9ePtwhQY88DruF
5vBDMj8hHWRph7iUXU83r6ht7XqaIsoZUPHjp9RBvMFOMETbkk1jRpiH92v61fos
P86nf4SMkZ6AoMp+sE8BOsqZO6Zcooe6kUlsaN9vsENMMTa7yul3GE25whG7kJ1w
P/NwENfSTCwiLRtxq6gbSeKtqwUuLJ1oyrSJaH23gD4eAo7VnSF6VWJK+kTPM0dZ
BIeYyzbGzmjerfZ9OFIp7L0TvcumdW3dxUDIlpw/V3V4T3q49P2SKQyvddDxFD6N
SqvSKmMSnC1Wbve1v1Me/aUmS5vv3Aqlnt7/kcSDF9VACqDO2zy98OdVh7vIU3tY
d1qZQ6pSk7R0DRCl61IqheP/Ul09IcNKro9Z6PZ6213r+8Jron8PrY9VoXjEck9d
329b9gnQkVwjomjjZY+TwznJspqKFByuFpHOIX2a8Obb54QTf8NLiFIpiX9A53hY
k0z9Ptjrl7e5AKVgVREr3j4u5oRViZDJTzgvTcOeNyh1qzOlMvchSelJsNmX6/oS
1QMLU6n8UE7iLELP/33ugmngEUzkUUEyQFDaeUWOxnLAZSv5xfT3jpdi0I6iD5kI
RXYsn+Ga+uIhSw3r1I/yeBC/c3h3N52BRjI+xy2KknYN6uATR8qolmxLJIEnEfPM
On7NeEOwcp6iMSzya/epItfAP5PfzDE69bBkoPhcirmNuYidaSWnTBXyrlKN2di9
LZI2hCJJbybAZFE7G30c5PO9sHfDbMV5M+ON1DOEyDR7rKV1+PICOfMAA363MiNH
mARCoukNODroCujfSUvKVYtarh5d95Lv6RSXI0u/MvDxz7d126ZHWOAJlk2dg9xA
xJBMPmi2petYve6We8ONMaHV0HO/i8PnTq4aWtcJENTMLEh2G20aInTRSawbJ2Gp
OVOfomJyXkpKv+nml7tu+ctMpFBG+LT3eF7Ia/f4D6iLVzWFkubTv5Stevl6UhXy
ifewLsXMQs5z1sJhp83m8dj95N1+RaPght57lLi1/T2Z7VYxB3WwmdMgBEaq3le6
wpTenWVB/KfpFQLjNw2Sioaw6hR/r5DjDHtSyhEKVx18xnOaCXaGN/ZHYQ9A8KY8
i4BlnP5CXGvFkmxVwox2PtGqqEiR3qxbsAehTT15Nah7JBdIvO4uK9brEvNt+qw4
q4/oxxH40VOSD2JHNrYdLdphhCKFnV2wAXtOU5eGavdchSUnz9knN96u4ASIRF2U
ft3K9lwPr3rNcwmQ9CrrcTQ9Q3GyVtoe9ogVn4tyRkoi+M7Lkam4tBDs6Ejb0wUl
WAuAaHUBkiHAnIgsC5BzuDnyKUn3+Em1+yQVxKnQppi8lfoPJPuR2BSo0jJRUEjW
W3eHg//WxeFPb0p7cvL+gyBk1rlJ08SI7gppqk+ADaDpxZZV2d4xPs5ylxs/sobO
r6QyR4SDsIUSIng6n4TIhsNpB4wweLZBkUINGyf7ISbwDzXQH7sCDUfK0U7GmFSK
aIWPZw95jYw8VALvVCetO+oUb5xxS9y2Dx87wvSAvy/J0inp4y2eu5W060vtMcXr
vnhQTLqmqWNnqNFFtd8ltkt1F4vmATAioMk5dSxdO9r4q0QRZvr3mhQ830v+GrfO
9F3XpFMxxqpdCTwjs4qefnBQX8sBNoiRiQFskMW6VoXeZSdKtIEQEUm85jrxTUH+
TpkBGa04Z86U7aXJg9qBK0IpEhjTcDN4BLJKWx0ihTSVMmamVD6/XK3TAKsAam6B
g2N52HyItMKH8sAq5HqLlSDEX2tOwyRNU3cSxtk/NK2w/0hVtGuh4DowbXyMuKkU
v07GD7uEvRsQWPmpi/7Gumin/IvUbNL7K49JkZpFHSZs+nU6kcHOl9uU9tWsJTNs
diKzJgJam6XCZ9RhDwvsyN6HzzEBVjA+73+gxeDF8nJb/uFoDloMRvOPcOU2UZD9
6/S7f/fN9M2G3Hz0hm3Z9ZYoEew/3t9EOV6QAvIb2iQK1IHBewdkZzqXLnKCNRTb
k9poE3oQKmJWO5p4OU8UPxw2JuzAY0atglBdIWaO2HTM/IzB02necWBwkcf1rifF
TL7a09WttA1LNlm9x1ANcAfRbmjm8B5Hu01zaJkt6I5ikrkWmIQAEW+/wxRZKaso
JGUzFQLNkv5b9rbdTHc1UJv6ooOy4wCYLjR+UYKzq+heDGGusiSc8UmsqLG3aUmc
qQ6ZK6sEKRs1RGPgdC45Fy4mVbYx6S74leyI6Z53FVycAZpqaI2VlxQ1spEdAfsV
ge8WsxJDRjLddGk+vBJu5sb0aW8TMYYddx6xwqLHUNH96fuL4GSPTfGnq6Ai2kLY
G0ZLDQGqWRoLS+1/0o2zogjvTx6Es8mLSbTeEY8tC0FlD8nYXaT+jJm4tWaWkW0W
rjzDlPiZGNykt3bWgKhTtMm1sQMFwKoxkuUnpsxy2XKewJU28z91lgzNIPKXsoc2
lBTEcUGbxZTx7hy562i/kj4qUvspNIzOUMcMd7vtc+AMpiaL80D2EvybBZsuK4tD
wYVRUamt5zKpE1Bz98f1AlAEziqIaio3WUs3S0wsBHloVW/45hMAtNPW4gXwtuJA
03VWYRFurhPjKkBWtd4XRrRqfFfdhrHhs+AnTuc8pcb4cEEj70mJKR6Xm2rB02th
5vVVn5MTnArmetdpzqAcuxXbJmLemtaAkmMU9AWUryXpUd6kpIclIu2lbBbH4JvM
1gaopDKUHIIAXG7L+crj9sssMk+S16hDaZ6/kbJZcFuE3Wc3NE5wlFGz8Xaqexys
+MCuqIkEauvQz3In+xivrjJ8U4zsB435IrVnliHR3enLBfI8/nmkZH9fzNOAncH6
uInhxG//v9W7oZDyIc7C4h0Vgru3j/bg1Ovb50KAcy5VaKwK6MeOCJbukGJq9TG6
L6Y14u1km7Jmiw8PkgVsptXn9wBDKn7B7tGIxADj5zGRhLkK7/PsbLNnv/Dhpsv6
TH7PiUmS0GtbYNTjV2pVGny6LDNuaTPAZ2edo6e1eILk9cvyxGiHQG/6tsDNidvz
g9FGHD12PmVEtxl5tVZKLjxo9YB2aVOgAmGbN8Ddx5kVczrLlfw5ZlIVegHbekxQ
nEvVtNlh26Lekc1FxONLuE+sbT8mOZAYK71azty57QJHOodjMz6gW8SJJT07MWOf
fkbUC8HMhPIWPeibNOhFsF6yBHdGZmWpiLcg6kfHz5JkxHETluEFm4j+5tc5tDgs
0T2tmOUA2jNmCJOuWFCNIjNTMSpvLvpDIegJvA5a889vy93JCxz4vx5QEqalthQA
l0v+sXbHO+ETbDzCGAqn2qxApQQTxCbJiL6542vtwuaVMwPIQxD6Bu5ywzzUtDWp
JXM1qFpa5B5PiF/sF9jzh9So+hfVUo3V5k6M1sY7mD/yZ+vxKkBuQFz/I+hyleQc
y0EHVbwl18uwRvBh4L628aJdWDit3fdpDegrqXEyXFGgwBeAWDszYNxi7Ek3b48r
1lgzc5ugHhPXAewIwCNW544ml4BWYohJRNQZH0pxYeJGVgJ4ZOXwugp5/G/ovRx7
yKDgCWsxoUoMYBvWTcHWFLWcWDFIdnOCq8gZGRa0YyV/hnMmlWqyCY06ash2HaXO
mwePOmQAn/00zL9WndnfeQ30d04Ipxlimk3SKs5uykj8rcwAY9zc6+Cw3LHM0V+c
tAmxQws2mjJL/rVVwMXfLGVFmn6HaYpXsU9pTT0jmOTZSrvpATUBQJWQ5OQ8mE5n
62gv3tQ92Qq75caexwxFwHgyZ3XkoiOJaRI7Y5mdKoAUosmEeuwfDzH7RRrqeJgo
0mA8A30uGpRSMgABau+XRT1RruVOP7GoIyfDq1a61KjpK/iwNss6oUKlcooNE5GZ
bZjUetNTHzynYDvyBJNDzb6JFOp+HaR8RVi1dtSLXms27/I/P4URV26puJhuBK6J
IzAyUMJ4lIJ7MHyHtRmWYZ6we1n0RwnvoNPJ1ebjtvsl3L3jA7FNEc3WT64OiTmY
SyrgA8GoqQ4Op2Hlfb2Y6QoGlTTBSgfBZcJibzUiE4sMGlIxoaSupi1nVNTp5ILT
0m2PqXpULtqLLeKbkKp6e81jpXQuyVtWxKsLDZUE9NMpBHBhdVvGpraIO35YEQyx
/gE3gCGuMWdvxcPvfFN1AOmLgbqadUjhcU3TcDgLrMdKk50oP0JbQuZ/igV/7/OM
5/ZwW/iac4saa5980/uS6fHdPk/y5SZd7/ie4AP5sBTpMtUWZhxIoptTfmpZv+cn
Bepy3X/ZUlnG4AF36PnXnxwP5peWty5CjbDNPbjZ9Wt6D0LeWRQCjqiwctnws7gV
OHWxqroHqZUt1OHx6S7v9L4Jqw8uql3Mqy2vgEd1NNw/OUFEhGCzViEzF/BzOZCT
b3/kcH7Ia0yd5MRCN4pK9EVFzRXbpMg84ZJuYXfuNA26cDwvOK5KV0HIL1z2SbNQ
gW1NJwe8uJoyOaAVyZRD0nwD1KGVnh2v3tIKr7YjFSRgS6/4JKrBwvW1gMsxLNq5
3Xp1Te2Z7FCSsfu4+bth9j8/xpsbGOeOMpGcwpt7D47Ft+x2L/A1db8SBkNnSWrQ
bQN3XmHcYBJJHPKtryBb6hiWVV95SvhUgqmdC+F2BnLIBMMPeU8XT5fRsLUa52H2
rRdad/N/oItE66vzG49ww0wydq0pjGoJww+BS2abY2IsSMullnyMEMOctz1d6/Hp
DrkEW8xIb54M2Q8XngzWhNVjJ67kERiY/vPr+rkrYAREj6Pb1I5cPSSuFBfhY0ww
4xZmINhi/tooWFWIEIY2lADVtQAS9RdmY1E6LaDNyBjXjPuyTGTtZBIq0EMCYjVP
J8E47/yXuYG3FSl9QCkvwOq06AR/rI8qFb2wDwdLOaAudXF8lk2b1r/TQ0x24i0G
AfRSID1mkBG546YhyvKJn6QB+ONKh3ZwL0C1w6zhtdg2OtQ/EbXUWG/eZagntn2M
E5ZLIRjc3YM3MDLyTChf2DjwUVYQUqWJxxjtXXnDJ8z4Fcf7OV6sJkuLmjG3luYt
7iajAVDdpOPkn4JM6fznz1vlLhAtPrdcA5WIEujRS2P/0t9FBuFNrgYkbyyVn0RH
8PnYdpgE84PU8VlicIA3nBGaIGYJasgDbdXCqLsBjLnhKq+4ceLwCEz87ojs9Cc6
EZNyZHUW3RHNgu6vrL7uX4TBF9MPvzv789gGJ8EAT0glclHoTnpvJluLW9oEvgn2
b/oKYj+MoH5uj31qK2YxxqxD7++szslzD1N1dypnGzCVWIMxgKLns7QCmPdKSgj4
W3yEnwBfapA69+7WcrSHUBTiqGnoweCqiZdBvNihWN3lDwdhpfXnNVYSq+bXkZ8P
hvx3EzhI3+K7FRNzfTBaHrok1aKag5biFcPNh5CcOPSSt71ioTYg3mxY/8PBjsQk
N5NsLgkG3Rt1sj2o/hJqNkaQ3uceiYSjaFB016VaYd94xlkKPmW//tYyuLRqbKwX
xTsJIN/E4UTPzKSx4xZheLq/7bcEvS8JBNCfilrns5PTAN/YtqD+mI3qj1QgKiqP
e62yOoWPrKcTXQP4qwBfmrZG8biLxo/AB4lbHkFonE6PpF8dKLl+9f8shKEvtuut
FgemySPX8xdd7uolOYHGcts/MkN65grUv/0cEiDXR+kjm9TH1q/oCG70AeHUGVQK
rPtjqEhC6mflehBtipgz8pscqJ7++61tKWIonpPsidEEEeo7dmK5eXao4w/4Wk6W
4Y7NamXY/JBqB9axY4cHP5cxgVMuSRqHrAXNXbZzTCX6U/3rqKmf5z0d0oFYEYlb
LS7BIEYGcxsumH7VBJ/b9GZPGlhe9PZ51ygEhEluVL6go5sfXLxtmEfmswuCCJWM
5VmDLTOxT0TbjSWIMW0bNJNvHMacPD6CSGTEnawFc0krOHYy9bOsTMdvpyL5zHUm
VwBqOXIW18pG4V/6V6zzBYkh5EBJwaxiItJTSc7KTYAslyn3kF8vk42CdF4IE4Dt
hkQ/BioaniJcmi+mPf4uS7d5+o3ks9krAwme/lr1b9RklpEIQB7iWoACqxCmczli
/8sedbPiPYH7lHIZeHOcJEBNNDtg/Nk8IwabwtkxgGvgjIXu5Jb2xhfRw4Fjmxuq
bHeoglwoHeuxsMJdbSIvVRTaj4FTkxi6DjhoC+Qo58uxE/qBhAO3b5Mn2pToqrZy
tFEiybMkmLoHTiYUTXg1pQtbvGQ6QjDQ9O9+J8P29K1DPueEllZeLVwylvpR2uNE
xamQWjKSpEx1A3MoZuOErN8W6wGcp9kNA0Rk7ljAuFkybIaC0vmS1g3PK4TmnXus
RfCIA/+1ntDrvDkTblRAQIP9JnibPyBfuPLAnqNnvTDKnkr7ieicupEJfM9RIgMs
qMuzXSf7ypHgvt+Lpdw+0YGXs79cUdx7wNDrrYy8WvB4f3ZCCgwB0gafFDqqpDK8
ubYGDdCJSVuJnI2V0qhg61gxY1DgV96QtMCIqCJC061t0tIGIG6Xj4klH7DVOMd+
PNGWLOH1Sm+nwYxXVOXi4DmDDjaoXZtmapi95HiU+UzbxnFE1zd5kCXz7WCm7a7t
hAjJeZVQPzCd0qSnUHiy7+CsfcG350QrOCi9IHEwNoBRUEuulnUedEynMPROpCEO
/Whmga9kJeOMlk/skZo6BwyYnR/dSvSG9+BaJPKUKvyVeyq8UhKW0nj86Pn/fmw8
2hB01A+sH14PQvbT+B6jPvqX8VFliEat8sBW9U7DrPT5DAxxfgjU11jXECgLrhR6
s2q3+i2Wn+gN4wqD91Ey8+aqwP2O28B08wP33+9MlnOK/wmWY3m6yLcwaWEXTJxb
rCkCgLKkNQ14XLGHdSUw4aP/eCq1iz4WNsQLPFexLWWG5odD42Dd9SM32gK8DodR
NCm28j+PUNz37ztK0bdaIEAb4WW6O18UndPBaCMXqJkXCZqwhYPfcd5LQFCxFBf9
HFdinsS4j964TKjinwdeTdk3o60xmDPmQUiXsUBA7aleEwS9pcj6HfsabL3v9sWx
wDnA+1MzbHVw4NCSClK80/N1Wqe1cYCzWa/LtZrsZJ3XbyZNKg64/tT/63GEGSHz
New/UBIwqr6brA939XitpFwu9TJ2DUUZQ+GslvnMv3DBu+7OcbFDk0yGj5anmdTg
kYKv/XP161DKn4Fyb9J5BprwwF3BpXpplAXmhA1Nrjg1eoHpLI05X/E9S+UpzDWE
kCxqhyvFBove9UTy9Ryw2FEz4T57oY+45nINV8vSn9mF6ohtEcf5OLrZ2aLK97Hd
JzNmzaJjnWj48U7FyV0+jeshFp7sORY+L0wYH8A/dWW1nVFtWjWlCJk5on2jDvrW
f7TMMLJpjgEowEWueS0Bdd+0ggQGnU10iydaX1I5SPjiOMJstt/3Ck8D+QtTMEkk
e/hHwU3B9w6skLS8Mlp/5CrtAK3tredDogGCYplRmeJnDSQdAHKzT1RjaiQy9X7L
pqeNgVuxLH4pAErDN8SQtU7BZUh2GPH3WwlAptHkykChBtWBAomqLUYIzXQRdp3G
zOYIiLC5fXK7pwZQpwIeyt9J183TsW7NRTvNRKn17TSA9eKiWfK0HrBKLhec2acu
5v8GfINxMCo2nP0vCuH4UYhxJY17ZlWbaltp1NX7bleU+Px1miOzYZ5+KFkJ29k3
8wBsS62XYB0XB91e0zQE4Np+qsCp3HjGxqo3IheYr3dQRKnYge05tVgtA9fQywQr
1RTJWUsku6/xgfzWmXY8bRx+4mHmSR+5RVQ9i0i6zNYkfPy1e6ctvsCCaqGWLDsG
VsJhSvTxduU8a/zKxnKA2JnJDe2AVUlgY6vQ7LTKELTHQcNJNTQaqIPIkrm4PCqI
cP6boUmJ0HN8eAjVWM31AYcdCZHPq3+XipPLg1cvtP+ITLuUYOM/+iEtLNvc8ccw
vy8jyq/FqBoGeoD3eY+0kTzf1aONXYLG2tUUYdhSP4czQVMDpcwD87zhLyVhUurr
fG/rwoIJI3DQjP/b6kDph+Uj1sCXJ7kLIDONblFZDorL0XPnkDHwy6O7aD7Wydon
rVoecuXF0li3stKWbaZmkHKp5JRKl42GCBdDjHX2J5aMg7ZwFkgF7gRF6qI5pfNc
RwSLA3Y/5KehO6UE6/xbccf9NQqmLFek5lCi8VU3Uo4R6YIChI6xsILpiM5PLEC6
Mqsb3EOM7Dw2VHJva/bcVMnW8sz+xYltdfm/+K5BNk67d6ISyJaemNQBZZMJON8N
iTqFpz59RpXJRIjZ/9KoLpze3PLvkqohg2Yc8n/1k6+pwpTACjWiw4VieiSeFmxL
On4ogjEulnWeoQtjKLalpEzWj8b1nu9Cw5ECcsHiBCOJuEXwFj1vwkDvJt6bLGf+
DKCIX1NZ5OcvE7XkpTjJRMHcXQXlTdjXsswxyuO3KrBrjn1Oivv/qhhxaORBjmNg
8mFPR7QoBJWzkErP9EoROGAJZ8qkDfoGSD/7T3tD38v1AA0kyMn9wViMhp7sAdHy
tIRKRvJHomsyTQ5ntj5t5UTc/gEVF2/aKdKgGEAIZ2xdoqqqXqreLjeC5+lNjzhB
BbQOz6Pr1x6NjhoFe6F8C1rkrE3mdLNyzmTxntzoY+dNyobvxBVZi3Q9YikUxHyj
hRDTyEaiZWz64BKoW8sRuDK8Gfp8SU+T93Tv8BRHZtSh3iYntgtyxqFUA2jSMoV3
kU+oiR1FreUl+7N8R6+TkAgFiBKYGmFGzz5F4VvuW9CBv7R0Z8penXaM4cz/faHz
6uuAGgtviZr+SVvrxhijtesQzw0ChRy/FrgIp0qIc89k/rhEh2M0Tz5VRtza/gu8
yrxzs5rqC2WrO7ZT8QUmoLLR/l5aoBXb3GTGCRFl/9QbAZH2AYx3xvvJ2d58hOs0
BBSbOyWCinLF+eOgP3vcHXY2uFYbQB54uZZbW3YGUACho2EKpdIKjFWBILNHYtX/
0goQOobjTELBEky/DQ4OyAYsnET5UrTOVvduZNLnUuZG8w0ha7Yl1Pp18KzOOs3P
wda2nhaIQSx7PndL3DPGY9rg9eLeATAi2FVGq40S6LqywaFQpfQdnTFLqTcAD/oa
/FZzhYOAmBlFCusvcgpjOjN21SsQ/yNRjUBX04faYa33K2pwqNrhDpqBwHd/aedV
UmPLRMoq3BPyyMV8crtZh4vqbR94pAm1pde1ufPeEEVN13xeiiBUt/qvCe9gwXgb
xbANN3MPZBEfXXQCaF4UXDM5keZO2QAuEjLo9SVNxDMHSs+CAox3mFPxJlX4+Xgv
LFFdQJx1v2ZZzB8VBq64C0ZAqauPoAWL/28TnJr44BPgc4SxxsikZ+HYtqgRqI3D
4bVcKHdbHhiJNyXKYg1Wc+4Ohea3BjBsf4FAHVSw0QhM39fd0l2CKpSi1POfL0/C
prB9sjyHfowf7aNod8e7I9tQ9+MgzwzsXNQ/rgt5ba+H5iaX+/VwUuU0UAn1p209
ZkLgHg0V2ZVN+tQ6vAWyOO9juDREfCiMvCj5MCYGwmeBK59WBAodckF2rSrKXMNX
4UFTX3lvwqClXoXYwiUx3bZ3TbMVIdAKCE5EBjeqovefZt/RwKabKK21cVm7E3ki
MIJlHG62AdHCIFlgBEfvR9FkJjvCOvR0eY4Yz2943H4EGPlCcHblP5s+IXbs1++Y
bemheEv37jSp4wO9QZOlJS0gEanN0JAYDA5yLYo/vVUWhjLWzT3549duV07m1jp+
kgokZt3mFlkwXlHQhsGd+Nhv3DJjkU4hHIcp5ERJuvTqM/9LPutiEXw01OaGbW/O
ohKcrXGTAoHoLbI9ywuOW6A2z0O6CPPH0S9ESTr4d3uas5cIWGl+6rpgclX2Nx1W
h5dok3GI8stOtu50qOJ0dE6WKPr6nSvQrKa9QF2SrbiDg5jWV6oxeGAK+bQKQ0uW
zH7N8q1/W9HpfdsHYthT1C6vNCfeoQk936cMtrwqxF6yeQJXdshuV6dZIUU7LPVZ
XYKxcghwJopv3zMnAFjc+/3dri86Q4Fvu/HlAixMYdSYEdePgdm2YMPO4LvUANx+
oot+Qp5uDsHSxgYbOnLuJI8IZbReFw5RHzT0856qQw0UflNfZbcALHPV59QDdaWY
B51ToUw08Aj8FtgGBucEeS7Jc86oA30I1IzNJ4GOZwsEcqu6kvQlU3KHcvt+LKkE
38OSt4CvIeBI7ag2QjU7eBoXlim/w6qs23V2J3sa9V+YqQZdciO41VEvbO60jjCo
CxNWW3/FNM33ys5xTKCkTVRGNB6lTiY7KGv1xktgIBdAW9CTC9flWKXdvNSxw+GW
/bLjwbGHYg+x1Pr3ZVfRGVXLk2XQZ9C8AHHpGg0E9K6+eVIPbXVwXvV7CILJq7ST
5AaQ5YmrSD1FuE+ViftzIKH9LOSIONXSKemOXj5tM+KrQbt81ZoYLf8BL1L+9bUV
ldjSiOL2x9i6wXHNUyS3L16eZLc+qsMU4WklVWpA/ZRX7s3j4CObNK/gpXQPMGW7
0fa5/2ILJ2xGhMd6N2svDF2BE45t/ofsFfxQ3dj/qBBQc3cCAxy6xnjQAHY2fMi0
Yc8Iptg2Lm0hwqRW4iaPh+6pR6mOJB0AVy1T5txjUggMA97Z6LIjnK4og7HwYGhX
FRpgXwZKm1eDQGIJFarztZOUp7VWRIcT+s8SM5yIrC1seuXnZpLVW1ikdNPnX6bZ
9KzAQPGlq/JjMT6WMjBvU2jYg6WY9x4yAKVCltUr8SZJh5OSjNk/Jg+ozVPOX/tj
k+8CYQHVL2nYi2os+LMhx1apfEDFlmEyDW5Or0FHYKZ7NkOR8fkFdM5gCEpSs5ON
68NYtTbV1B4L0oHIXeoqZ6hVgtjX7RX9Q6HIQ8JJUC/T9tATYqddFBNdQh3xahD0
fNWH5lallBfVtOC53shSptc5U5g2uwqKGXBGQ2opFeKmVVT8o3YhxqHq+AxJDG9P
jL7Db23T4I3WUFAlILC/P4jZqQ8Nxxk3/tLG+Ngs4kArIn8Mf5tgB5H2rqlcwvcG
qSVaTdGGPrLslr8+aWMoXmkPJOpL7dr31ec49wn3GUvLnXnjn+CPjvl0kPWCZwtt
CcYQndSz4j+mCnFMjaWQhu+sN1a5zUMpqiA1109dUZeoslja2/B5FWocBTBPaaxD
fYuYV+SNZctiNrFLvPC+qBceWXye34pFlDYqYFxqpBnjFZ3NM214rPgawjKy6G1z
yYG9Vd75eO16Ljlb/kRiMTxS3N2MmOLKwLz0FHM4h7xlVVY3Zy8LfeWdF5q9IpDO
/ZLTT579hGf5EMgMNdvk+9VFVPMHJaeIxWRUG9X4IVJmDhAA6fHUORBK0xIQDm/N
6oH2+zKrBo0wtSulbide9I+kN0kebDNCn89XGxg048E+eDqGfR2/maukV1Am+5ZA
rq1osbUpigrt05g0k9XMOPs0+Ujol4R2bhiWUD5Gz2exdVItVqR9x6d4WfD43YfD
7z7mgMfarwHkxB7Z6IRb9g4QRjIJUAM0RFIfbt3EIJSC8Vo8fhAFPPzLY80qS+4s
SH/7KrrjBeMuerDKG5eiblNef0Fmb/AL3UkUxXw6owqmnAkbIAf47erFazQR75zN
Ik0d4yhjFqXwCtaA2XtD8WSEYFkSz3uQLmi+U4gKLxOwjzAG6zAao5/rjnD8XdjG
y5X/h+c24RQkRoLlPdW/mudU53U3+tEgBBQeFrg3QicCTsrHS5NvjOktbddKsHSP
9rDdG4TpdF9LCyDNwiIpUkrhhhCdYxVyVaRYwdVjfKX4MSYxXkpkHlVFX0qpR6qQ
C4DNxPOXYbDYc1HY+DQv5VDjgWG4JZ/uH5NGG3j05ZVlDrP8WUKX/acJ+4lBo7Lj
TqLsmMUu+uoc3f3+3N1jwA7H2D/k4R6vI0wCLrrFq2XMx0aaRNUxNY3DKYB09F8n
JKSBIfeEvGszqsfKHNCJ2aZdiu+8jw37eXH49HZgbUcE3xrIOzq/pAnK2wEEJsmI
6a49BGb3XxXL27LyVol8q+1A7kG90Wi/R664agevsPq40AabkYvNDH1tkvJny+KS
TLDf4gj01/MmQqZwBrKgkDPUuxNg6nrW0bOM+ntApH0b0c0rNX/x1EB6yWOkPblj
E8uHVsczZnolGgI/Vykf/37zrjNTbgb5VFLhv3Ek3gb0+bjAU824wgk6MtP83gHh
A/Q/cE4QE5ySHZhu1rKcWezPKL46pM1NV8IbYurYupAII6S7FskkGfiqBikksrii
GVkCiFpKvyoIncq3d805HMrvM5RxXT2Rs1B/tDC+glTnRhiJM81jfqfZaHu9VuH0
tXI6z9RYDyiOnbafy+bQCQITlp8dvhU+09qtlGSustqRXyqaUjAOKguiFnce8ZM+
H6qkZ7FuLQ/rNeUtnJg3KyAwH/C0r4Zot6Fn3uda9rDcvTnYdN0aiIHE3wW2CNrR
5JAzY+PRRNv3iNJh6YRrCPc4vhWZLFGCB2egs4MoRFHxm3/k2qw6BRJ1ad26efSI
Ox3B5HtCPz8/0HHIZyue68gfh47NMBakybgsCECYnWMEo0ZacfeyNt5JG4JbExsp
qjncxFinBTsrp4snbhpOSRyhe5S8c2Nz8AuHEH+JBc1w+jKf8kPTjaz7DhsG/78c
PdpIIPS+O+tS+nYi1NN9pw5Kyu7xzoPghMP9TSDWc59ASH2fLVOizs3PEW77t8fa
CpVWWw6pvJ5xeTaAAYtU7WXzXMjUAh2ztPNTfN4jpbf3ksoQunavM7TygeZpnb0H
kiP1oUmuBBiZFvckiP0fkJCPiLrX8M+0dqEX8SCVOG2YE3C+zxqDOsqXdZ8uiE2R
bZ3fCQj4tcDslKU3tCNGJjfFU3HpZRHr1Ilo4/hyDRqE7Ett4kvOY/E6uMmTnjbc
3Lnndjq+pnTzy2i9SXnC6pebw4FMDcdSL8kedMWoXqXLzYfj/YsKhABLhR5YpNBm
asOw6HpOocgA0DfCFBtt1yGSrQJ/imMvaLig3iULUbImg77pVqXfT5vQ+xSR4UVs
xzcPCONyp+4Vqm9x2DrulcV8FYZ8n1Pnen4jV/TYdubQRxH6rzJdTFOonfmHM6kb
IpSaBHcZYtiEQaJiWzS1NiSsI4lVVIEQVgDZ/ypYF/lXP1aYbh0Nr6a926fIgLDT
SLHG8e2ZeaUcDM489OS9U2YaOlCh5vgSooKLlSC9lCotOgFXjP9dmwMGEyJzAKBn
mmG0bF6KkWPyvDhLWV6/nHrkPEK2+3WBWFfL6e3lYmcTdHK8bq94MDLF/7ttCPb2
TPCbB8yg9TY8KVUM7jNT4VX/eBcUx79jpJFbk4Q0F6FkMhheLp34r8eSxjVEre6S
LJjH9vu0gxvGBWREIPgCMUUFSLN75AOmzkO0RReexASfB5wtt+SBWieMQ6ccyiQ9
QJqqbqRMD3QJUpaGSS4rccQ69ZfutldrRbJPV3UnB2p7gU+BmWH4L1bTxORLz6rx
Z7fxkBPkL4QOUuVq7gHO0MNTdGBefPWGR2Hv2cMUxMQbOWKFDN+BOO66O03MVRzq
EAGsoD7yGvntYBTAa2AhEQZbWOMeoSLscvj8n/Lm+ttXC+x0o3suhRfP0IvofOy4
299X4jmhfebdBrh/nTeLpiV/DR8NT8hjCY9TJIIW/UMiHXfv59RLgFNxhfaRmH4c
5oSVZhmcTG8vkciWZS10YGoIO+FcZoLEt06fmeDkVuxZ+w19qNrl6gSq11MQsOzL
gDnrOBWvVin2x7OP+aFxmpwwWfdn+et9wB5pN3+e6CFrIp5wn21cRK2FbOzv66HH
0o9NXeLmlpRxAx3XuEvZHsQy1VDS6SXT/pYw1kQrTWZ1Fp9nGj1CtsgQdWGo6Ruc
WmGiqgq1kP+6NN9z02TtNrbyQEJJHSA1sINxwduNUGq7kfFphFzFI31ry/+HMrX4
R3k8ZfYsQcZunwF7x0pobiHRiDAoAceGm0mTszZTt0kvZZW0lFp5HeMqd+D2c8Yb
0fcIYPZqFwPM4dsWaywG+XfN16N6FFyueQezTxSsRMcqT4TZJyCIBN0sBfAYHIS1
YNxzFREL2rjNLaNY97J4KuziXG522iiPI23ZVDOVZWEhmaL3JTb71JqdXfJN8o+a
g9UtWmUk1/fUpFQpDMpwPL8NopU70mUKvSPejHE+VrbghdZEiHEwpfzRdULjQOLg
22wXBxo9h3fy3mI5MEkZi0dPv8CpRwIBBJgJ7y7c/QR3KC36VpzMZOPNccywpoJ8
7+f4OQnKLPEaTpPUPYy9sObP7XvECkSRgdpa5eZkQkEh0QiNtNX9aYdWGEAped7r
hw/4y7RtulDzkhklv808yjsEC7YjbGpg2kg0BU9dhaJ93SdyEgVZ/SNQckLlExvX
TkVAkDN1xwhLFRNPyFNxP/7z+MOpodo4Tt+9ITH9moJKz/Z094VOxYFdRLZWmjY1
5RRiHN21uiaoVQYK3Bh8issDTaGiZsKkEKXA1VJwoHSQukZiRwdXMYJ/mzS19AsE
ZhkdQX6kJpX/L9cBfElKjOVrebG1Kqomm8X1Jeqi0A3eiP3KQP+KYkUCUql1Y/k+
NP3rAOxO4ZinMBxnPp1gr5UjxmyF95NGgGg4hxvl1spu9+MwfOASBwaKEOZ3eYfP
hwoFnsTm3Foa4p2bnq9EY7Kc5jQd3I+LvAsUqdjP2QwkSy5dyKsGu2uKGERBvscO
tsb3ff/0e3LXw3P/0YmlhSX9fSKGY8YMk3PWeLLIZ+lSfxgb71A3KRFwWQnuy5/g
SSJ2O4M18I4bej/es5R+MzFeR3m1gM4Cev4JuhEZduJ7GiH8FoXd4r6yT8gVaQf9
IuNlm1/HPpIJkH7kW+tHkI1wwptQFl/rWwn+W9SiLrA4k4CjlCtWtlxyhyauqWQR
BP2RNQyO8JwNliSvpV/huFfvPQQpGXxYuWN0CfeIQdRObfx7laF+rnsPTQ54GwUO
+724CNfa3LswoHmmyfyTjjJfY7IWzNAkJG2ZEe0bqduwgZKxkFrt+gwODxX+TJiO
j2N2qUzpbsAOCaWlLGlR34tDngEvkLz4wkVZEIOFpVxjxWEJ/Zn1WF/G1BE0rUxt
rjJHcdH3YXmqk7M6BYtESw==
`protect end_protected