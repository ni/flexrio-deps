`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2688 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
eqFSpb+CvMuY5DmKJBrN+h/GgGEjTlt8UIqe+HyUAP4Q/D/UpHx0jBpEd6VKbPLZ
cqQh9ZSJzdjyXOTSWLBPWv2nkTnWus9+mlt4qgy1p8fg9rKYKIOLVveCIsVsKTA6
f7RWyaTGa4G35WbQmfkDzgeiUw60aoR8sj67VwEeGQ4ODbsRHusE9NZO1cPjulQv
1NnWKIr6asbUk3nWHI1Zw8XlLFJMy4RC7YdoK3nmdcFZZvgA++ZGtwD9mz2pmPZC
O3PAvBBJaJ0jzNe9YVEHfm8JnbKLYzdiX3eGKEjmNSwOFgRibrK4HznrMXR+TBsv
skB8YAr/LOCnXauu+wUtytsOj5M/kowsvW3qGCmY3NvNgQ7oAo6rMEE/HTenz3k2
9Z5AYzMA58/NphcDYsIZRff/YkZNCkriim7Z3q9M+h3Y/rIqeBaUwnYhVVvZvX8p
DpOhej50dxo/mtGjHE+467GiA4b45jtCxjGI2xDXRSUxVronBrvFfBQRxmmh1vEx
2HXkQvJEWdVrZdo3AsK3qW4qQqYUphisdhquf7oVNy9dKa1RArqp/ighJFsmS95O
KSazhMXbSGL56fA/4Fb/fHtektOmkximH39SPmgooxQqpZs5iTpIIxhnzOmSEY5f
mQdW5I5Dx4xKr43sdFU1NDOzZ6tfz8b4v2qTNuc1us9Zt6UnCBez6Z9MBQlTzozq
k4bzwW13zpgXl1E7YO+n3ppWtBHyvIz70k32K8uflcl48MbDOBKXSeckEe8T5zws
jvrxWM29eIbWm4bGDb4Vxa44AaV0bUKO3USnjeulhk5jl7uCe5kwQLAI5CQoxVny
vzK3e2RIk0iY1I6sdkms+cDrdY45zPlUIU30f90JQsmnSbon3SitqxCrgLADQok4
PvBuyN2IXld+BMlBoims23gC165KnkFkbhcWt2VxTlfSKOpMB0lO1adQwj/fbRgI
eibWhrjL4L9bYWbQWrXnHm/l0kl/+K54egLanruvAqfDOpxvLcnVr8nrYL+rwWMr
ELZ4cQJUqEhMFwH5/ytWBl/4haPIF+TxWDm7S3hhzdgwlWy4/TuFUp0C9tR5mJ6C
zF92+aYp0LwkQZsEnUPJJf5ibH8Qug0bwFQ6uTJyFDSYrSijvfTkEb2NRkmsrluT
rIWxE9dhmh+2xJw27K6QY0menwkhsMbRJ7EUwdcO6OB5qRGrVmf2/D5NdPKoBcbS
UpLYGr6nVmR2Av7ct8K9cs4QREdnFahLDf4t2b4esAZVZFfa66OBbIRuzQeqkyAy
yWcS9XX0wWMm5X3ZLuIqseiY8Voot70s+eK9Lxf65N24B1O0rvVqGJJmk0+MPJMy
jkMqE2s6MS90ZSM1cWq8O21Sb+PoOFi4/+oFFKG6GEFMrQkYKSEpQqR2oHKG6+Em
NKridFcXJXDaUTEy8oLzCqxvr4FFuuCE3hXNZ3S61uE6c6CrajEyl7U1kF8BFfVZ
47EqDnCQweWYe4aHWKNPYzJPCUquBx684G8XyccsA/1ZhlMF1+lQsMwAm2tOjELM
f38tme891qFEPR3wh0117KNCH4dASvp8he/J5bq1JBS2/b/ndBL1itmA2IGZDB8J
U7keEQ3imyYyhD8KKbEVXtgj2Lr6N5seDMyE5pLo/5DZd4MEXEbdnVNQ2us38LeC
lDdSLXC/fawKGZORNtqxDfDt68K98iwpeOi4o7/1T+ZrCl2frAtFnSacMBLcg4J/
7F93kUy22yww8UK2w2ejF4GK51LlnhD1qKtSHI381E3wYMvG99MkTRky2eRxWRGU
3mbruDuF5iRUeyp/Usbm74Cm7t3vZp8KBZUwtPDy243q/DsfGnUZK0NXuddPaSTG
5OwnG8NLV9TZt9laH6gYfp2iWnr9HpZDubxFIQT4RL738PUQGqxwP5mxwjz5aw/h
Qo0+gh9A4Aan9FlEVFsBcEqTW3jFZDvElxgNS6uqgciz0hzVUGfpr44udQDZ3pA4
agrNilxEaet+l2z0X54/2ZuuYxp9m217MTLns4J7Ju3hUiD0WUWA6HONFJyAJiWq
utWQc4lEmYmUsTrkEeFmos0N4pyVpcjH8nXmO6qXrn1szQnOfi8MhL/3R/QnSPOk
ZQrpejqoMWChnDh0b6KbW/C79wB8ST1cm/cZdB9Q3zmtgcDH5wwFiLSDU++k3KmI
uAHFhAaxYZgA9dk558VrnA802fWY1BTJkWfP6WVAJwXxR6mLRllTw4np7TOEWKkV
/cwPvelYwD5W9uILsmRPO03Jm5kydTUNWUMelWNgN+BUtQ8fgMGW36VC5j5V4e4F
0ekxHdXAjtLKEkD7F8nE5i+gRaUwwxb4CXi7QXlfDFQWW9DLvURgYsgEQ6b4hw8u
+Tlo3rsS0N763Xdpy805+jiOY5OeG2G+hNYhcqxLZR/Qk6hcCRyvBfNArN8tSDf3
B5riQSuSNmrlCp4zIDHdfbOKC7570NsOLKdwG+2REQavH7POpde9bLf/gNAoTT9H
eHOK1U0ToSvv6uOxRkVKTFhLo+u9nhGS5a8QbcA8rO3whOfkBkmo8jj3eFU90sKF
Y4iS1srWg1WEfvpTbV3ws2d6KuZfLTh/WPM49EDuTW4eJmQ9MqqsjW2VgfC+Euz4
r3luBh3i6LojvZyzqUgu64PIyMT4NPsSTbTN6g6zpPJmU1KPmI3PqHX4sSFUnNTZ
yrGoGeTVx5OJDjoSQ2+8TKLQ4SIXgBrSmc0MoesYymE/gIFiOmd5qfjoHYK9MJn2
uZm5HF41BCRFa2dW3m4T0etmfRvSgQIDqkQ8WMq+paXD7JutDVocDQ66u2bQ6NfR
ClU2ZAFqYa25HBF7av7ZxV6YO/8TabC8tbvg/ftiyr1Z6MdKGKjte3TmIoYsrQmg
ylQK3/ZtCsb5mZwaUN2BOuho6zVOTbcUhj6vcnORomIaV84mXxoI3c2wW0MTXr4S
nqgJvezrMuR7X70V6f189bZmIzl7ZhNjTvYwvMYpafxhGVSyqL6BtV8Sh39paHkC
B4emAuzY5NSvHA+brr497CZ0m1bVN/rPJo8RBNyDMX4wu4UzfNLwIrLeQZKX5ajq
2DR62dpo746EKQ2H1OW5pczhSWCAskn06c7OG8CKoG63tDzKvrfajIDofL4wtcSk
zZN3BHwMkDG5b2fQbblEVX3Qtr2KGb6ecMtHNgtllE5dKB4GoHawK3S43diXZC9a
dX0PL/pTXuaFNQRchztzC4Db1rjeegtdG7GVGM+jjcFC0T3JC/Nmc1rEGOoz26tz
qLuTh5cRZxm83uYp1vNlsHy5GWDkZ8zWw8UV+8zyMl0LJ1JQe53cRu/SmsHAXumW
tqzCy58uWvY8TyoBQ19DQEsaVeQWVabFrNdqjGD8NBT1+q8/EGy/vjJNop3VDZbG
O+rwWze0uT6YTvUDpfGhrkOUiST77RgfePAcM/vIBGcUa19Mq47ERBNAGuxYKr0V
`protect end_protected