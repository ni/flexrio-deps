`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
YATj3kULTF7Ty4ORuRfFpnT6YIk4rUPRrM74bVTnc4GjdV8oSnW5PtQkMCLOi558
1V+/wvDfc3y0Z8//ksX8sZm3JZWtrxUppw8c14g9Y7owiwp+JumRtO1zuk5xFbe3
0MMnIxxoTKLhyRJtAxElG8sbx8N21OWDGiOk0Xyd5CqAmk9dcOIbxzMjW/wndBXi
maijUdqS+5KiRCM9+Gsp6k/iEAa2LnYTt4WtjkmDD1P5jZKsiMgFck8WOqLymplZ
ml3TTfn1UlLNm/+zD3SFGP0kABAiUT8NK2xBPQ5UzQ6sMFPd/np8iUZ5u4QLTWOZ
hTrU9OSX7lOvRUo8pJ9vPg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="BzW6NOo8eyBw+CxsNNo4wIDxODIsVe0ft0K5tGuSUZw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
DhjJh9S2BY18dG77XPz3hsiSQ73+w0XqfJhD+f+lIDHHVjOB7CfC8ieNRTexgzn1
5W+qoqOEwenoVQtit9u3XViXJSRJ0wfUC5a9axblRNyD2mUbyfH9+f59nWqGkVOh
ieHxkA/DPprM70F3APxk51m7/gNSLICSvbONgLGndWc=
`protect rights_digest_method = "sha256"
`protect end_toolblock="L7NTNW/5Dqy+2kJZXKczEa3js87UJ8H00YWI+92sDHA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 26864 )
`protect data_block
6eHODtGLmq6ccbB074dgNWpdzW45i5jL0Nzx5wwM+RA0eeOHXxEV143NNyQGmZjT
bzHAi/6AyRCB4X9z0c4MjyrZE8GF4crbMH4T59xFHqVrQ4zXCea5w0kG5yvHgpKo
rwIIbW7Xn0p+GsC0S8TZEmVtFJ25Dp0bWrmdXjXTdmbvKT330FfOOWETejx3Q2lu
1W6Whto5XWcxtPbO1mr2gKF/F8UrWVsl/3KrxXrNlX7lE/XIrVwXnEAOgyx8hShp
NopfSq39o1sbMv5YZnfJGs3VqopML/kx9XHRz50K9Jxly5iwGyWd/OxaDoLINSA0
7m7Oq9hNhEKX0s6aKSD9bf+YC694BqEj932ZlYm80ikJOcObEhnf9Rwkx5Weqheh
nu+mPJkCL19r/anHTZk82zq/cs6nildWMQpi8iJx5v9gC/7KEbYyzcvpLlWSCetu
zWMvF5bQbwwD2Wy7XrKwhoU3WB9O3B2NBWaFY0Kr8CpDV/2NUYgochDP60RpudkJ
dmH2i2B4vyi+DnCt4IkYWE8aHfXxDhoyi5uvCpobGFTXh/HCFBSTTBKZbzmiOgBz
75ONr+KNkf4EGRfuP2x2FBwCMsLS29IqclkpnBZ4U1d0/rm51vgCvYeWbVuE4Afp
+HLVcmgyBSCog2ql7X4UlOjbzyFX7KHcUmj1BkKDamaND3fz9z2Vix7A3nsYxH0Y
LCXuzgvYzGTiN+hzVFMgH6u/8ZVLhuaavX+xKdN2AJlb8vB/QEcrxUx4QGbUWvTD
ZUmBN58fPxsTJ+0juBK+WNLYjjj19A87wdL9IGIpaBysGV4BMVeCJQiKzXA+ZR8E
giuNq/9B9S2Q1Wqd3cr7GI4KGI8u8/0b+vOQgj7bUFKOQ4tNMbTnNLtCvcqHadJ1
kpHZtQtWqQk1ok+Oyedv/2RMFfvaPrIqah7DRXzg4+x2iNDGl9615z3XmisuZAC+
TqiXsGssJrWSyDSVhyoNuGIbslXbd4zi6wsKfpiWyTjCMf2pSjk8whdQStLBYU3a
QGu9iO+wcpkAlrE6v+6is18oHfPGzMPx8hRgf3TjzFKOlB8OmKjZM3VIGiN4qWPU
Uu/coaRJwXh/249dwbtxvBbJKcsDfcp0qg1aPyV3uRBBGorLiScJcVcUeHPas4jv
td8t8PTR6BkqhVEXmT6PhJtQZI7rj9LDlpUkGeaP0lEYGaYm+yhTGCwUA+beJOOU
9d0CtlpuIVb4H7JwOVEHxu8D9FIhdzflKiyqmkKL+RJXUYVxStjrsKHC4hCrj6Xj
V6yUvxmL7mr6zI4GU2jFUTu6l13b3BUNxmtMWuHE1P1gu00EgQyUFQcoE2+o0+bL
WXr+uRYYmFZI8Znh7emA53SEF+EMi7Ct9WUV2H7IKPKQgt2YADbloj0moUq+zSH8
RgwAcopSqG6t+sFNqncDGP+MXqOkFYdKObKOjD+jeTCLIlKKOYvO3zQAzr3nJQ7B
UY7MLuQANutx1G5b/3uhxN5Le6gKlJi+uVtp4TEkNHGxw8jYMhLmdmaTKP0Z4OrR
I0flAZhoOpQ9RF8yxp+eG657vcqXH2SxV3zOcXfbTGqk/XldZ+T3Q0acowzPxjNo
wyfm1PPNwGUFrtnSPicmBtg7KIWruF4IPPim79crCt9fJvwZyQXQK1RQQP6gRJYy
nLM/3VlFp29xYwrdecCxRLN4annuFoSd66/9tyLS88irGrqjl7yNrnqqo4/f4i76
QD7bU7CvT0jaxcU5Fk2tHb61vPuW8vBlgx/JRtSSm7AF92Twqs/XHDKrpxlgSMES
VacruJQmizDfy8NpNt88ah4GO7o2vHg/ZlALHxZUFslTyd1f499hOu5oU4KlTJoe
b88Bu+PkaCoIXYVojglAbE91UN+fTpF3TGkWutpBqiHdBNSLdN4CE/bBLf7H0n9V
dMdiaygoengJ2kcWHeY74Twzlc30mVD43gUHpsMrmE3RaGG+K0rAXfHe+Qpf2KD9
diLU/RRD7qn7HU8jwz3nxmHUIlVTouQ6/5clWj3mJ1/bqfAYyJ8oOg5i3pM37bkK
Nm91pklOvPhu6/go7eimqa0rxLYGXIoNOdL08mxFT8y8ATIfna4IQ6qxuRXgIKD7
0ELA9lTzjyNkJQ8N2eTIt+83pxOsPTkoylWt1Zue/wWhqTqkBGluf/ivqONT8qCR
PEwSHWts5Gn58R2mrfjeX4q6pYarqsL8VTDifR5Y9D0XOPgYLnUidZhD46JPxSZB
SN+PPZMYth72liswrzq6q/0NZqsGBcopUOLzM2vwiJT9zbdse6/4RTHEo+KX/Ejf
Sgn65C7AANLkRSR+4HCltgPhKEdE4bQ1MJLA+J7IxbEXlv0LW6BfDAeP42B85ng3
hv8kygcBHA4Bg6yq3X93KDjDkR3gTstw1apWeait89jFXBbWJSmuyKT9xgTWcjzQ
cr9lj4aylSEykzYJJNdn1ACah/wbG+YqUzjCGpLiF9DAHBkGPicYwyvmxmeBf1vl
SvjnE23Iudm95oebUAV3CySJ5cSwgBeOPg++IM9tTx4PcV2lYrxSfbW/HdGimCt4
K/R8psllYiomXTh6bp+SheXQfOSD7NmkQHQ4hFR0VLylLQ0nOPS32CrqxS0rWZs5
4vzPoyiMa2p3gqyLbwy50tUM4hG30ZGdTT/sZGCcL6P2r4/piQVOu8zSDT+RV0cd
zenbXp4FsbNbqaudmA0AFZGqBlmJ6oaCSZjbvtvYSnHb1++QfjEle+54zwBOSmIS
Lp5aJynpVblE7eH3Sz6/etzHAXDKv4kXyN+y8mro3EBLubSxwrgictyoXqXKlaMd
Yd0Ne7r3NkUIf5hHvCtubgMzpiBNFang3dguQBPwAK4syyeeF3Y1sq6JEB7oQ34B
iAymCnXDKz1OiPCC1a5VbWrKJEdzHnd/QlDTB1kLlL/b4p1WIvMLPaZi5fYbJXyK
hmIBeTrIjXQmJK7Un5W4ak06ObanpmsCB7CSeoD3LwkAW/RSDgtxj9m+99lLhw3i
APxDEmlTir4QJMcno4BViREu5TX+9qnzYbgGwgKlQL5o1bRdTKTcm3P0xGeBxgMx
wEnMeOBBdJRotMf8/R9/eSvG11ZzE/IDYfrggccfKIhNPE1S/0pr4bN+TwWsGeoP
8yP6OYfSsae7yy4h9yQGPfpldbRb6KVI12SR/r0wS59fOwuiwnrBlWUvMQ9puGzG
G5IkLNLzMzrzYJDCCYfnZ8V7TBRzB0rC8hmr99CAdBX+65yyZvBmI1+uekqaFT8k
xBYD3Fwb6jSEqkYWZi0wZZGvQQfHzlcEAKOzNqztGJbTKUNLb6xc51MvNJv/DD8y
dUOYldlC+CeOlKLCD4qWwTEoQ5rh3Ig25N219qpbboR6kSiXppubDX9D/V1V8T9y
n9xGEJDaUHmPSGCVtuCx6yPlVXrPsFSw2DeeKoAwOnN8nqyLU+36EkNz1RtKEDZ6
1vF47znR4BQ0FGFI7JLweyGlaaxOulk67EfYHdmN/0cbs2dK0pSYwVW45CDOzliz
RoLDKsYYybKOhGwcecUS5YClE8ndi4PQifErODcESACOfxAjehKKFQir2vvWq50C
QRRMm6STYm35Tm16aQFVpGdl529pMjmyyUXaQPsZlfU7zFxnyw6HhBRuvXWBiTrX
PLqHu5yKpbQCdFndzCyupcBCBAne5FNUuO86+MOYQIXPKvA/l0R/8j1GevDLco5W
JBEG+tCe7XdcQBFrX+YciC4Kmngu/YxjcbKfapXnAqI2wND3pdkyQz76J+xmPesL
yvqeiCccz3bCZzPmxYmmEQIQFBxvL7Rn8f3sXj+L4EzZB+ly+VvNL1MRNJPsr/9x
PEuNmCNsm8EfIalZdjgUBantEZ1fXXvyIL+TbD9/OTqV+aR3ejlu9kcT6/O8aMP0
owCC3vx4hqn6pPwFj04l6LrPHvVfSS5ChWP7otdb/rF/elA2G64F5RbarNndO4sG
zGM0U2U05gYE/d5kmjyZKdGtJMk/fot1KAO0ojLFku5BJLvqGh4V750yYt+75f+r
1Mm6fW9JfffUlQmHGXsKZ36vSUdmB3ocNsFMpHbV6bLa4W3MvdJIDJgsXPDD/4eu
O2PodfyYvGdQvlhEstGqi8S973kanKjOfq/U39QjBvphE/+mfqd0pnDOMXWU1eXu
55AXbsXNuJtxccn6BJgbZQNSSWvYtyNPQ3iEqIy21/FTctL/gfNuja8Sa3Gzuom8
pua6SWZMM95J2YXgoiqHPLa3GIQSRkn6JVGBEY+GdFuLn/RG1lLXMNaF5uKv/S1e
f81cb+LdIurUtkjmDJhqZhhiIUki/yTyFt/lkIbF7O7hjGe2522QxgvG1v5dNNWI
w5YJaQOY1RnAVBWm7UTvZ+CgwudQl9fU5mLv0eA9H7YeSXfu45BFmsEznLonpwC9
2zPEpORYdoZreurfZMXr8p+2p8cqKoBFsm93RlC4jTeVtCZMGNHd6QMcF64SD+U5
CRb2nAQ8uc/4ZDU6fGlSG5gX4rncV0h4VCw5FaM88cq0yWZjWv6rUXI5q4wrEhuL
mvyguNqHx0EeAiET2/7t/I1pKFqOgdU5g+jpU+PxEtu4Pz+rBVI+LIeEnOZrA+FX
QOfD1mPR60G38PbC/4M6OVkfSjAaelPFF2z9F8jO3QBm1/bt4z+mrb93lvuV1SGB
nh+4zwi9YVJJliNCalzT8hIguMPRbhe1Y80MjvWcrAXufgXBFRiDBIHaj6JRNlbF
VblVeXBgBMoBZntxI/gXZZ+JOg/0gv9u5VkinXTXepKdX5RBkA6bf/OTAnmtx9Zx
M6LKtEpRfvdh9sI33KDmGAhBcZepzDQYav+BZ71avIF1m8q6cHz63Jk/tuz8y5Nc
1Pp+HOkyhtc8fY2V+teAuY72olfgFf/p0mppFrWqFrvCmohcnYhPZT+gUlyN5Cct
aeBPojjkzUHt0Zy5IvPNSRL1go/F2KqwvALUcCvEsPDp8fiD+ndFCofp7flMU4u9
PPKXrfmrpea34lUsez2m5tnDbtrLjUZaheTh+t8ZYPEzfSOH06B/ynhOlhDNhd46
aM0z20HW0NxuHDBSf9PxnnDZsPQ7ntQQrQ0TGhG9DYYhVAKLQ1iTuymKaJpWey8t
kudGHxrcFr1Qu9zVBb2ZV6RnApiSss6KvFMDR+wHbhrIeAo53NwdVSDKzb8dWyzy
SA6AZiNbqb5q2T9eIb1/2ZmG44LigeeXtYcM8vYDAQ3QdPPFqEUpJ3R/gss29Lh3
S9WP2BEHcFZU3PU3vVqM28nQKOjs8LegXFxoNehKTA6ySGadbQ/rwIcZvk/XwBpj
MSH3n7WnnUa7DChYw//nf6inCR/StPdDt5vkoAN6p/o0aKtuGZjR0vjTa/e9w62i
GVdaltz+1kXMPBENoUvDR/qN8XIEgdxHu1Reb97Lvk44+D2UcDY2p4HyBAYQJFuz
2VQbz8gwZ0RgnG/bY7ruGuOKmx0R6WvOMnUrfgj1oqKVU8wxYPW8kBBNDyixPB2B
N4kZTuwMxbgwCGJndqVMN3tWi8FJmQV2RM/81OVymQMCiyrlXcwiyHURoeNvubaq
BlwXixdPc421OMGZzxlh2JwNz4xe+6Zce8SxSmBA50cetLoWl4XfltZ44RR6YTBi
v5+sVLE/sPcBGT8LD68MDMWd+Vpmq0z5oKDGZDdoiPJobT82wJf2AeB1+XPcfV2X
jslSLleUn571D2BmEPrKify0w2TeMKNE0vyfNzTWl7/0vUbWC/URbpQH51SR3n3p
CD/KdrqnymxdgiKFkriX36wWyQIXzCaMfqgLW6eObwmRI6Uniu1b63BUPoQOTk5A
7xoDnfrtgtH/Ussvhw+8iCK6T1drmH/ktnpjyx2PwSjy7pI+1Iqy5/NtRLElD1Cp
shxYh5YsYW4UjOOluYmqHIe2/owTZG4UzbrZu9XAIWqy3vHvZjEKQqpiRocyU2Jz
ZhADD4ch8FH0P8uRXN+1MtmXG4TbCif7rUajLsuNs3olnfl1JxVxK15pBcn9h+i6
VhTkz+GWEAB+d6m3jljKzjrIadbtdOOlyQTKjwDlknFoQguGhlZ1/Nn5/yn8eSKp
VBYTOfR5yq+wafEsWsA78459t4/yOPwPIFDVUrB4zn2A43+Qi/Ma7y3TaXADkhl3
1XLf7E1agKD+slZi9kz9QeHv28fkxoL0mWzlVWHIIhZst/HDurpW6rnBP7ijnIKA
Fho1809ylJOTXp/s23KuD5rW1Bc7P3z0HIIMeZSD8ws6pLJP2P9TbTLaOUqPh/qO
VYdb+C1CNOTCtx23EXBpeeUKjzx9tm1HQJR6y8WM47100YMrPh8rygCAFD+AZIY8
5gut2c/PbCdj7tHx4U2VQo22ld0ryOu7Sy/O7rAEr/e9y3jivzW/ttU45bKpCkVE
HNrr2S/7fPlf8AbVOUze9qUVhWlI7d8YCD8R12vEIfoVPHRgsn9x8dymOpbxD73o
UkGdsAMyuozgb+c78Kpt+G/QIeLvA/lVnhRyPF3bu6Z/l7QVrhEt1aEe76ZWOdR7
fTc8NmWw/+tYPdOANZ9tQ5yOhgOhyjZ4DZkvOYcwstFr7Ufuot3sPCf8OT8gp3T2
gYLL4JcGGm/DBVvnWeIgsK2qPTk7uentW7/HQ7osrigh8z1bAWQeVUVh2r6ogRVM
wesHjb5A0H2pqRVPjhALI1taStZH7AXFOJ4IIHCfAU/Hb6Hph58wsq+Dl1d2K/vB
yxPVkGdlYOupRwuHnI+kbNv5oL7doQ3AVDZzHyYJ+XzPDkLptDd8fIW3WQB4y1Co
iAm6h/Hm/gWQuRBMLv+Tkl1a6WSf87N7hzDv0QKcqk8AeOdCfNwite1XMwtWffSf
nQJas5D+wLLigPk5Ptub8e8wxmWqbyIsa9vWZUppVh3V/PKmFOXyNFoixHPlW38X
ks4F0sqOHgwrRmQUrs1xlZ5tfDM4V/1u5f3UQ82bKKVg/DDAudH7WHbjAZiHOJ0D
kjoJdU6rDxDczRUpnahATWWt2oBofjxcPi/qHA/mydXC+sECpPWO2jyiTZRzGk9l
MYOSLzZ8+4gNt/8Z8yXxOymqyaxVUnLMIt5ney7D2aW3j6DzzgS/8WQFwYvl2jyI
FQRGC1T9vNINqfkInikED4C5VTuBxi4SlTdkgvIki9oboJ0gMtKLF8SO6/r8Y+o6
JlVmhtbsaT0H7eSOPhodx+ouKKcm/2FnGr+Ig8lSSssq0d6F+ZV+/KTP3bc4v1iV
fD8HVRE5kTsFWq4sNSgNRATaffZ8hoEI5L8RDcpbAZkmtkknExTbilEe/Hbjb1UF
s73RDHgq1nHgMjoJrtRIrElHcl4YDqUM+flGbpJox2QVFW9SDmvqeAcjlaDpQC7O
wRKaHEvAcKHir1vJJIK0SULdKSZq3eUrp0XTokMil8/B+c93XgU/aQZze1QS8oZJ
v5AtkIpvAh5hgz00G4y3Egswt5ePjWvDuQCDkvtZ/VYybdImBWiziTjyGWFKL7+v
6ucfHjhJ40klQ+kbCJS1QQC9cfE1zOs+Sl4ZXwiz80Jcjbi0uCeSjH6wxTr3PF3R
BmDROi8fSKbGbDLySScX8swU2DP5ad0TGOX79Znz7vNm2uGjasfK2srVG4fBx4tU
bCZGgM0t0o58ZmlRa63UdlJlTFVAAUP1By/JnvBje4zUZcwlaP8u4F7IcUhFJSr0
HbNxKiUGorHcILo7Fi2xAOLG3mXou6T032neUChx9288mg5+Ma/er8w11nZIxFYs
TRrjbRhuBF5bUMR3PISItGnIQ1v1bOQ5Rj3c9/BVMUp2x07xLs/aPn7hn2un2yF9
qUcOsDuq53rxtTcO3Pxhr3HGDTvgr7Yh5dbtUETXGTLew5Wm4aPUMRoQ9/gKV9my
4OBXRiNgsyp8h8aON+SGHZoLBQMxuwfBJKxeplnJ7ME7xNeieZN1hETMg69EjzgE
UHvTBqK5vtV1agq9tuyFbVVB0JaGtZGi+O1/Dm7ZDEfCaCljEeu4e4NCSZFF1pvb
KgIMBngnyQCBQtlvu5Zdd5JvN94E0+CYXCEP7EK79mdNHHbg17jXywtr+L9xbMCn
euQq25XlDTaUtp6B5iFMND7Mvxo/KH59VQcKZphiVUP9eUTDZDyp20r9/YCyFfJ/
Jz8t1C+m16tI0WFPA3MTbv/WXnXqIR4r8uDOe0mnsg1lWmSIFz4F0iwLUgZBiXqG
7SaRZJ2ky22PDUQA1PcPRyYbaxwBQTYJmKj3C5hAswh2wdbhDY8ihAZvFRDQJn2C
lsXNSwE13JNxqx9pfNxevgJS0WIcDRY52JuFt2cXlqsrFPs7c0L6gFVM8sKquJ6C
SihwnzJ7yMXHmORdxZr3CXNSkJX2a6cNlEua5Va42hqQlnEgGAbOncrHpG4XoRmS
y6iSoaDoYFUUGHE1m3aKji9vDE/E9K79bGVEuWblWmoVXcFRZ1RW/qBTBApo41S/
JAn1hpSaja7w0jjqeZKh6k0Tw1lH1aCsrDCmNzkgvzri3YWLKl1agLv4mhJuymlE
iikKedEaXtKkJmoOwubdU3Fz885+LCNS8hx9QeFFA/7oCKB5sPRHvWCThVTqk+mS
fuiRgAON9M1gUcvo31l46dOmASpJOoaxKksHpxQODJW8+KSVL3Gzry42fAic25Tu
MgSSygv0I70zul4AqZbNSwV8jYeChYNDVUQSVurB7J5f100zagGSGE8mHH3i1LD0
nJkRvXEZp51o68wuarwb2HT63el/2CLBMHLF9S+r5yGfPtLDJyzHdE4rfcyfHXG7
1rtgcdDwTX1dIy41akOiuAtvJfkS1DIputeSJFY/2RpfY6lPQB1LSo+eblC4Wbb5
R/Nw1kIDnWltozwcI6736LNUyiuMuKyeV6JiB0k4pgjPfK6nMIpu9bzi+/WyGTKx
bo1DK+gSIeMb0hW/QE4M7MlSEQTJoAD/rPJ5gk8Q9OBtPkV+nkCcNNNcxrqbphBd
z7t81F3L9AG2ammm8Be3TfG4xDhZqbRpLUIKuOTrM1SKVxfNlCxh8nVmBcGWyCp3
70va+u5ziQgLeyBoHOr3HKozMXFt0XvIZHJGAiIqJniYiqZBSEAikyT0xu+6rUnp
b6ncf2doC+K1hHHBc58iEXqOjowaTBPRRUjGKU0UMSgoeFSOaRlm5lUCP9l7C8Sp
fBx/8ZMgWkrGKxPLjfeCVehABVU7EjWcusB8V4piK33f5fe0qwPHzFpBRFaxYLAk
k64xcvGfG8VFth6Go8B5C3U49+wOoxa2Vx5hFO9bDJ8AlBfynExSfrAhcY1uXNrL
O1i0a7xe0x09jJ8OVSTHLoQmxujG3JiIm09RDaGqYsmLU69rxkkKkvHvrwtuRIZO
NwGZtEtIyYyA87yjNmBfCUMKSeGNHOJc+3xj9j1JnU6D8lExJQNzsuWxnBJdZPHv
OwXaUUGexoOjAJ/KFf7KylYRmy3hPPr+g+l9sNBF3JwYFCjE1AAuDG9XSouUuluV
OrxRNvqUAjL2dv/RlyZpwy71cBa/i/0LY21kikK5QJi0gcEjdz1uoRJp+79FxEE+
4l8TXtAv/RXeoEz2S6kKOiZsFJU+P1HZ2Zj8HfHOuwnOTfIX8Nycz3kmiISp48Gs
oyNCvr6gm3/lbd5/j314QVlLGf4cyb6DQVTtuLTB76bim4ZxfIAprIi1XtfNbzEk
I7lS20VttAmJ7dn5FBSsg67KzWtHtNYDN3j7z/W6MJU/yoUZYTfTDQCW4G+GX+T5
jbDi0/PRWXtYLcmH6D37vhZFyeyNHWGU7+UCgDoT1bp3yNuY003nJndPRp0imuTo
Y+cb+MQHPbiATZCVLl+uY/01krKtoR67OEn4SWa9rOkk0+oF5mlXVUOBX6ouIfT8
8thg6wLpmaWf2cR0BCfWAsnT6deskQlQaeXRVjvvb7TS8MWRQZvOdp+RSfb6cSwG
/q2vTVpz4TyFzNIVGprT/ar+qzfTDcDVKcJrUg0UsPj+KzsRpKmBazdYVkwEW8LI
Li9FEkbEl7SJlNEa3GFsO5ixR7Pnqp77sNLenaNZQ52OanVrbRbczy9VasxU8wms
R+iL/qcC/KJD2/eujvdzZyFjNWUMndWSXX+6eKZk+Q5/SE4U05/VKLa9P/fmNsOa
iq4sfjoni8aHu4IBFw+qibXRNWZCeFuW/S9JwZ2gDBfI1HGrZ5t9t/e0AhK9F47m
iLu2sgmKQNuLIsXSPoPd2SEwXxAgv2aRjU5oxrNqe6GtTq6OLdXlZZv38AUeaV0J
5Nf49q5M37M9KyVN/58vy9oqgMAZsMwn/tPoTpkgjWL52F5De6jnVCQUN9wGpLyQ
KEMVL5zljISUnRmjFUyXjaClUl2rWy1SqfmFguvpOOIVyI7wmHvxYEJ7fdgGHCr4
2cg0pjVb4kuK2VJ/D6tePeDr9EF91Ajj6sGqqVyvtoBiPKZSp87b52BawdZjSuim
pWDkOLBfylPyAZgH9CoSAFsTy2DB38Db3OvjDMR4wOc6iudRyxLn2BJPbB5iVkIm
9TXKii7gmMYvWWCZ1IjPm+3m+Scxrm31eNSTHRZI7EmpTTcKIB6yGsVQp9+j2X0p
Kqtr9fKhkZ6jiXloBTcg12Vg0CrpOTz7fFxJJJBfZONCO+vUP2O4fTgGcJ1dnPWS
KwWLJfxX0WjM7c/KRowQIfi0itIAdNqm2ixFR9znrVywVki/HCnAcAHjdcl3PSy2
4hJ+zmVtVSFQBUECEGO/gPqTcFo5uNGpNK5xIOBW6vYs9G6BCa7BuuWn/9BOVklL
wgzQlx+EFhSFngoc2DOE98HO4e2hZS1S/GiS1r8yk9zaghQ/VpCSgBwBqU5g3bpO
Q2EQcPaLL+38Q0uDPhqXbKRw4Y1np+fNoqd5nJJbQv+Tjt9o7NMa17SXSmZeQ1xH
+zEl0SG8yGyTZS1ID9aXXDACgbWy22aYDFMblPgWa1COOsu6U0aF4pBWJ6Bx3TE0
JhqV5cHHdKOLiZvKCXmekhZSVpVOQdc9AJdP/4MnBQPP2hNWe3O6P4oO8joycBfY
ii+qY1t7vAhe0C6mv/+3QuLB+bpbUHklIUKmPMZAiAGF/G1gRzfKZCoYdJtvs6eW
e8k/oYO74HoDlDZVV3zuKYTLuBB+jSCT1rJ/ic3e8XMLEIJBJlvWdTH1ODksJs0c
6UZNrKMztKYpT+iXkS4DuHs/AX6CULPlMGQ11GZBt9jsjEIQgHjPy6NEq4AHwTXp
KiYP/mi3XeyCAhyQL0pyOoJB4cbAx1vQdDOt183zZHGBbZfWV29ThWiNQHFQsOMS
+dxHKXo3BVdKXUxFNY0EaRios6C0TkfeKjrilmRibLmuOACUVIsSiSAYB/JKKjx7
cV/9hnoqNLr093dghina/ZDBWdI/eaoqQuDP0CvNCXLE7oCU739qZw+3eD+7ycpi
C8cyafpc0C6W6/UB/SVVkQW3+o87MffVXlyGOXpEvczCjiNYuu4hv0FXUPeNlFNc
U2xFBW1vQBkkxYytov1vl14theYke3fE5Wqsx7uYzCttLd8QcrAuKQ6BvL6pnY7a
S4BhB2ckB1pnp2yQQGMpVtFNu0PYVcOrWnc7bWfVnWYgZRDdf5dYc8fGZ8RTpIM7
pUN4CJkA1FF9gpso1LQ16dU0+oy8yILcNVQxrsys8PqJ+OvENNwQadmyN7m+4mOl
zPm0+0gayaHRntPQT7cWB9EpoXUs3RG+Qcw05ee9HSkVltL7W/lFkXPBdS7W4xTg
L5I5U0nQWYIuvTTaVVreXP9gzPA/FyJ43BXU7SEiO3b8uO3JTiWVc3Tysjf3w02p
tbZhSvN80qcOqzTu9J1QKH1MiJEyrvo6h3zZcCgJBIdGShM4SGJIrnNVNOyFKc/D
ElcMBff7BwdfeROrzGZ+wMXmWXRLcf2LpXtCiwzf4JPNo5LR7DE28QLuZwlK1z0k
MmskDPgfFgyBXuqwpRp+uxxAGN9VFZoY2Qw9Faq2LHYOhzSl9hbVZxmP68/m++bb
lfxnedx3o3ynnP7sRIHu1y/15L0Ntea08Aq81kdxmmmzUpJWZJlk2VGAsJVvwyy3
Py+CIrlAyqV9noneSvj/S7j7VBmrSKhNhHBTr7P0ZguwlNbLpV2MAI9YrcesTy8M
X5ZqihSpywBp1wCQzX4GLn2Ymvoumfd0CBZKel4zTHensmHvZZHInyi4u1GMn0ks
uBj7jOeL2DI5g7e2VfcWZfgemzx0sHRJhpzTzwrUmoLMJfHf6s/Fce41L8unPHB3
tEw0Ko7Lzpo504vuQUX9t+FI/ZfK+tuVzlq8rEiCfFCV+XbSv0f+Szk3UanD3GHY
pZ6x8liufrmoZnUV69YHAq8R+dgTBNmlqqsyH/eLklplWFN1vboEE5/bE0mzU6A0
Cc2+3kc8hn+iUqE+iP6YsQ0NK0bBd5AsOmvtty0lASeUA1VdSI2j6EBPCk7kf75f
uj+mxKA+f4y2RdWUPCbuivlYSZJ2N329B63yOvmtw/wREykfK8kL2oCO5VSLAfhd
sj7BnY0pzMVLKbSb867dOgXVT5Brl7GTlTIJhsy2ZX6gKOJ0alNKdf7rOuwm6WTc
kMY6jB6Fd2hbp127RWjXEGr21rUNK2omkJ/ajb5HdR0i96zHiTQNzHEJ/9saeXe5
NNBFKU8ego76+iVLbGx6WMewFuoOF1ooSRzPIIQkVOf0E/M/pplfN9wbYrhfaxsO
PNVMUEueCcx15y33wlBhtVZfUax673yNm7PtarY+cp7POQHZEOWVyy4NQ1BxFZu4
A/eoi4EVyYjSFdy7XhbcIJBkWxEASQrbeSqGLDPz8R5jWX9SWYHKvKuhAmbWgGtq
xKak34pt+axmF4eWwWcsSlsE7AnomaOm6zcUTtihwwLS52D05ECxDVB/w1U79mGw
w+EGS/NcKpcOnqfInNKfxraDmdIolBQYtE3srnz2DsJVv5oLOmeZRT5B+YRw/iWD
WO8MCvs/SdyZpkcvgJlnElYwjIchEfSo+X0XIAeZq52zgU3FyQBeACMdXcgFDucq
QsB/y3Erkk3a+db9yoESZqs/R+z670BVjYSnajGqcx7Tn4+el0uzvc1YG+9NaGoW
e0kRFihZzOgpa3VYBmO5T2cSKkpU73cp3tookE5QzHko+g0t8XAYfaIZdzi5BHZu
/FIvItsvUTV4me+WxPCsUbd7yT/0zgIzp51m2AbkZg42nRMdCbk21n46PSwdeARq
vIflokQRUSYqI2/JEyMMXlDHlBCtsNcBvxFWBoSqCUTxD6WzmZxolDtBpZFvChxe
XNriG/UCGKJ1PqPRPWqgwal8scWagOvZqPFbERyjniuYpDFjh8BxNGa6ooAge5WV
TsBOL6o2o4rAC4C0lR7uHEQGohC+NhkvyDuCT8FXTTPaZmtvpiAB7cZocYslfHWH
4WLX0S5EPDHwMxILvhkb5tgeq2Vm67yz58JqlNTCHCgYzCQpJb/zm3FfP5/+WaB8
TnQu7r7Q1+fUqekCT9g6um38ZNE/P596+yro3cuctYW6UwIBfWo+T2RP8FQ/KiVP
GEr9ZsBzSWB4+YjuW0HH12HgKRgXoTr9u3eak0Y2Li5h7ZYdPyKtB8q3nI2u8r+K
vRod2HCD2bKC4fzjMUHD0k4PSslQ+RhbajNBNpV0g4S6fCMpTYh+VccOZUUb3OU2
+RY7CiwuMPxnr7vZkfXZXXJ8wyL8x0rrcEDPfIOcxI2hYqjJAcaTkzu7eHmayspd
92LZe6e8thCxAEE7+xB5oYDQ+dRDHrT8qSxP24auQuAFNI0jIIu37+g0YHYyBz2X
1o8gfSfnoeXp4TgZjPfmTHvi/nESTjoIfLReGbakIb/pnFIJTpVjaV7imZw3Gbge
I7kSM3L1NXQuuIAyOoqNoO7BVap+jAwg9NlperheCkJ77NXm0evH88DxbD+kDjAA
tSJyWeezfd+hJyPqSZZ+Q87KYP+Zar5zApdLvTqFc3cR32BTzBtVLj6XhW31qt8s
JGRgqC6HaLl2/Tcb7k1/jVT/pN/wzQkhcUsWGr9dbMLfLr4MeWWw16o4nccGP54M
+A2DAaOeBLbqTr9VUZsd4aqDp885MO+3qwFrH6pk2S8i/gmbNxIGsyl+yHbbs8KF
uIEruIKUyhDQImKcpyOrZxuw/CYpXLW2voP1IjH5GtaVnRqmHuHuTYEFIALconGG
D+5qsxkFeNun8K4WzYh3eVlKKzmNXp6uSwJ4o7YXDpNaK0Bc81rEv4iUTIxtypQM
H1jMtmrUPBxxrTQKRi5SwWOllOaF1taHeaLfAv3wf9Fpv3qnqfW9uhEOC2gi7AQc
F9jtNyg/wZCdBwqCuDOku+IPc/KIx/OMj4yQ5/LPybMPuj/UvcgPl8fcseQ2NbiI
ioL0Oke/Ahs0/5wCvL2P+w9UpiHC4KgsjMmEiX89NvlXEg0CyNsz3I0hIobX+6iK
tTvbvv3SYxipNXlLbI9AiqJ2il2cl57oVoJXEIiOOcr8lrruXzWgMmKLSLzKHl2A
+kPx780JRn+zttCr9ZvTbOaWqhzM7nVyUw/OatSSSjhLPA3Z+rqSwdcWzPNmAbnN
Pm5q4lxlifNRnaXsi7jLdTQmSnv7cEFb70XrkiXgIqjoVCY5/rrlh2cV+N46UC1U
j2RtgBxPXGZQmHmsysiPJhImO20TLJRlViCtHq/LEap4IZL4zb5tnfU8JhY61cxv
O4RTewyWatpCcEmUQqzxT0+6+vxTRjnRJBSP1zHUTzNCAsDGatYjwZZgPiU5eiHU
5IFy/63JGm8sRsfXnzr1ljUcTYhkSEtal5Cb+jym/FqFERl5+TH10yUUdaXb/9el
N81XrOtpt3+0f89Cb3lQThFulRagcWq1Eyq0il+377nsGPnJ/Z9PBcEpztHFLGlZ
6TYMP2oige50pSYKm3STXrHGmCCD1MmN9qeZVQ/v9ymY7sxAjQ869c9eOLU2yWZf
q3wVeZ5K8uGr0t0+Ll9/YACrvTAF5wvB2aQ5JQrP6bkwP8HRVx9z4bD5/iaqApMY
sZcDrOpwwSODTcc47rHWe5s7vzyhiHQ7DAgr+/O7QpesbXC87WlUbb2YfQFM8f44
JC8tv/dwnEAZvi7ezR9Fp1N1mdDF56W8HZyTeZaG1vUJKxEhI+1FQnPS0xgBTdp4
zMB/koo/8MNekftwVfanQAqTNQHPNYegh8J6GVIVWGRuKV/JHic+ikecm6gHan9g
4x4N/EYJcsOQTFsG6jKmhpek58jUBuUjtPI4C9+kaIn/o8MlL2GbQWW/2l8sjGvB
2kwLvrUqkGt2EjU8V0iBXyOqOVpHEbtlQeP9jsQz4E24O7thb8kX5cTEw6NyoUZS
nR7zpEv/TwW+fTajxdedCleNOE81/0cWZv7LLq9bmrW6GCepuHvU/p9v4wDjkHFj
7MiTZuJhPN+nDGIYXU2+jwk3g0Hm4Dt36oprWMJ8uUNBV2wdxGy/km2boSjN7rVO
NGLLJ43wKmm1OzHMzlQ22a3xBN92DL03QkFYI0Vg6kaqRvAgkPj31NtNBiXYo8va
HjrzjsTqH0aEghdlWREYQ+RYa3nTaZl2+zz38wXTB6klYxcjoUB1is+qMtrAgjev
/+ReysHUdvk4ZcAYcwxcoRuXNa/AZDmX8YU11LXbcaZN8c7I7ue05D0rrJ76rtdF
MV9O1skY9kLzfy3mkdOxGF8G6MVylQslr/twb1LrQg+HVrIHYkzugBnVfAxekQEJ
xkcUVSB5SbWv9LQNRTs9VCLGTG+cLuOnl/XxSf9HbknqpqCIT/+AUZ6anRBThMmi
PFfQMyjSpLY4g25oB98/GafO9gGaktN1iNlqlqRa9lqyWsUQfz1WHh9/ELr18tHc
2oNGJoX9cgVcNFWqkOhDRtfHBLWHtDFLtvRGiyKwx9Lq5PPED4NXFCMScCKNpOzL
D625ZYxFT9ZTWywV+HlDnDyNGB6SfH1SjJfdt/BF7FZh0uGWCejTZ7l0jSLykEP9
wxokIrEln5RHLZIhS0/GArvOgxsCwWT2IliWsLqRM8j0H28J5f9rT5tuwrUx0Vb4
XmxSUQDhr9B/1ply1ySBLAT2AYfEpSfUoHviGYcZHYkvLBy0n5+YHO5+tJ4ADQrB
LgkbLZtHhAkPCZTTjB7QUWfxTVgMbDP8nR6Xat6ZKsixH9y04GeYMijG/FsO6q/t
mV7mrqflKfv+z4kNI9kYlt9EEVX7jTHG/h1S+q3QYwNCG9mbm3XJRPeysqmBVm6s
t9kFw6uiIVvmzR90sdZ9pmnvo/HEqwUy+5+VCWAplQMtsh9VOfuJwV+295UvxDCT
+lbccFheFmtuGitxmKYULAgM0F/zQGnWu8Fhj/OYbXvlNmELIw9TX9EjT4NUABqB
PpOEayRm0m37+tgoRtPfZoXfPPxAroGCvJAO2t+M7hxzcLk7I0WGAW1aQ80wP2CC
YMYUdR3Rez3/49iDSpDBckzldOhI7YEXuYcFm6X6kBlMvr/JvPy2MIFmkvQdx+c/
wrLb2v8pUPveMLlgAQwWz9ALEvG51mhMJjoMRBCVNblFFpJg2z2IM/aI9lE0MXqW
7zW+JWeU/SEF8KzN9IzOJBa4GZIfcNheKtp9GHtxySyBb3AMYx7UlPU42p126KuF
nG+uWEC7UV/iysT1515rTnyZxC1lf4kaazpwczzfYznp2G1994zFUcKiKroNSjvj
wtTjjWbK3fnBY/w2Kz5p7WEFSXG35tCE555c7FqWZks/E6uGs/bWOiBuqnllIwwP
NbmrbUhEXNzGguw5qHtr0ebWbocX57YA9vXQjODIqDV1OIKw7NFUMVVSg2yZriRS
+xjWybqknezz6ietT35qlSpF6Ev5KIqHCnid0vs+OxzKWJgSOdWrW7aEzV95OyYo
HJz/GxJeoZFu0/vGKoFqgY34jYjlyT1340mFf/GxywM+7duinQ8WRBgZkKX5xjwT
GvYP9t0dnoPZJh4GIOW3OIKucpnUjw+VrLyHU5Tgz05jSXhyE19sKR67tnP28yAt
bh+0wsbxSoCSTV4dM7mneGDqlxQhG41nHNZCqCZ5jWRb3jLAXNTOGdwBtiCe1Izj
6EPFAOhbyINnAewcacOJ2cgCVwz/jOh1dPjekvHWt2dWFZILDWqysyBFbCrte1Ch
Ozt3tRNk06RrzXcHCjoFUzJ6qi+jmsyscVpjVpuTP9DJKyWjPAkeXnqeXIKvWs/U
BXD4UrMS5k5rUMNhfkDG6ivOKsP8yinZbr7fKCz9ZjicnT0EDFv400YU7S3w2diS
MkKcS3XQjk5BX39tehJQN5g0Re7rQPfRedDdGRxnLZnv/Fs0uj0+iPtSsgkQCi8G
X83wGSDf5zyo9qyAp5egmkqlAKX5KrlPUJUEHQAgQzhxf5CrfU6GFfmiuylV1zPf
S74oSsexxe3APZBu5NTcko7qoOAcm8j+Dl+H0WqgCKShwTuMxhQchv+pn+6qRUj7
FVZjvqicBeikPkNZchK0etsG3fldBuXrRLFLHdY330rPsTa24I2YqcdSpT4eu1uP
HO6WoatS5wwZULaJIyzy51Df4jUSEY0V2sMt5COdf9xs1bMU0l0vFRPbYLUPhufM
zi5mHXaXLVsm31vS7lQ7owJJabDLn1TxAXvdRoB9H4n1EG2tQewFr/QGivL4xKE5
s9dY3Wbl0vDoWNR/SKrxj2NgFZ3DTo/dCCatrDKgGR1HZvgQRHFk+wftJazsDJzT
/DbE75zSIXI9GBBIPUkmNcOf1kqHw5qILC0dCJeMk/uNLXSHJNaG+ZwmoXS/CiKF
mdOgjgl5HQeg6JlCoBqfukrj4ZVSbV1JA/hdsmqjQi+T6xKgyryU6xUocTap70CI
ko/Uh+6D5Wrg+OsAJtPIl+mjCcHsf6TFEMkDZQqnDnii5UZazNO50d0Eae/K6hUk
YcAFIB5UUkgESWONiLH3nwzYiiMwI6j9az4wIVzy18xULcH7L46IU/bWltYHcW/G
+Vb6uMCAMHgabHschBR/TuKWeYI5+soRA9sQkVDh6KG0gGXTo0QN+NYVGfdn3tp0
HGc+EvsbTS1i5IBbJaVyBjVidPu8b8F1EMrrhfuux/bebjpkL9o/pEGk1Kn8a1zI
4vbWgedrpfLq5+Sv7zdtuzo7N59Y/ErnrETwTgx0urT+PaLOalDTTpHqtFkTDqWV
tadgklDhAmS/Ry7M9rtvS52JTdqWJKvda/ClbkCsKlnieJssWnY+PhB7ys38b79g
vJPEokyxtO5pMjLwNIEairXJzaFNeGH0M4uIgVXWS/M8qAiNGNMnkf7Mf3v8AYzJ
vEI5vt/T8AZGwiy0hKX4UpybuAYXErbdt8uZarvea0NeykvDug1rq2x8X+B5MsSn
E54vToguduA5EHVo0MdWwkoZSIN4uz+zdY4/YQFy3THc62feZlpwvF26Cv/TUmxN
DF/yHDZYG+38bgEbonUcSoVruugU1nIqtyp+rK0Cb+rXnljy+B4f2Z8iDiztclLJ
m08c9frhAalxJHuZ4qlhlgEbjLcEqHPYBR1j/sS44Z8b499n8A97PzsdRXb3b60p
mzEFjkb6uD1x3fEmVBk5+E/r8F57EUQBuM4BpaR6/qVKJOYdt/KeZw+z2CWVG7Bu
QIJlFVMek1OeWRKc2E1U0hxQoX5c4Vl+AznLGHm/OdgwvCfyNmPMAT/yBDm7RzYt
4BvqfBs1oGcS1erwaN2fFzLiOPFhOs5KXfSfhpFlwi+YUib5lQ95vTXafo6OIpjx
ztITo2ksdd+qhMQgO9V86jH4VxEEjMrXhmnS/pBBisdvelM1l6CiB5pZdNmyd1Lu
bhvDCwxXnxYshogeFLiQ/PN0BJdRbc5Amek5+e5i31AaQTO8w5kP25bK+ua87q+r
6gkCC55QPiAfu6eXN57MFRHQMzxPIGDCxiDQL+yb019Cjifvyc1byOF/f0NGDwpf
GiRjpfyMzbLdshJtd0vun6hZxz6d34/vtZAfvQtaCS9h3zvHr+/g+km6oldiUtoF
A7YkLiZ86ZiYSXn/s/UBWTrrnpix8vTgQBp/B3gwIQ4BwKM1E7C3f/UQ0sADYKF7
uBKWBgVuolDqyIFT157Tsa6xS0VpdLiytBG/xG7tz8ByJqmpBvv09ZGGXjMpyhEH
StNpqcqdvmkmBkfoxANQ/doND2KSWPfkyKVDS2eDipa9SnqxSKhyoAOFgKg5RorU
9HMEZQBUT6Xs+knz9WuhWzYjz8wMIVvORJWn72f/WCsHKJ0xC+Qogk5sgR/NMhpZ
Xlglh+D954jFfJFxJFwpTy5Cj6alwNiGjtjP5IRcOrpKSAp31Vd6F+pJ/kQtavXL
9PSUFdsvYeMfVYTH9Llqf4top+nV6XeSdo4ea0GP1FHVJXz/tk/7O9WNpVxPeMFg
kOy10OdLWHHkmSGIfpvtuNFrVCJHCmRwhPkE0RJwdGEPka3tZIc0F3jdNCuqbNAZ
4YvfrC4wUw44M3qVXsggeDXywOMRtk5dNRQHQbmvJJ6qaLDQ81qU6Gpy0tuNvtns
e/SE5NvcZfzAeRs5EHyTNSaTW/8Jt2ICpym/QApCKKEl/15DuovmIqspN+JFLpw3
jdYhN0q2JieSjFGp7eretZqniWxOp4xHLuWszYHYm+YDRS+2JOgJrV9VHDZZ4p97
YKMv7Yo/QgwvFY35Omfrtzax3vIc4Lf6LEBHSJWZ9VyPb9ULWIjWwxAyysmcy/wS
kjnZEgSTb34QpR+Ccb825unwfumV7eRRWH49nkpxxnBjm2jsxAYOjTCHHCAGW2bc
cQKXTrE4R2awl9woIYe/w7R1u41H9P35PuDASkOdCVmq9tsTwOXdgLb8iACC3F4V
vVNFVbgp6f8gisK9TmElNycifCjQtY0uspNP2Qe7bn9nm2gCmKAX/Q6JARZ9HZGD
IXXe9lEVYMLjYokHM90fYJuC5RV65TOVuCWwo/6xZziYptmQesZFB8lrzLDjAk3y
t8pqzX6Z57kHyACBP0b400coWuSHR+sZGcuMtD0kO4f2DYJm0wgotVwDZ8Qv2679
Ig3yCO3ixbHchFAvpETFCaBW4dTfbC+hSr/9gGSpWSWPT0p1F2Sn4e9++/YRA21+
3Oe3O6kDxC+OR6Q5xrNWRs3iejlLsuyhcI4ypXrkD6TOBgEBbMjvw7KRuHZLap55
qa7uWgJjefC1TQmokD9IaDSW/LrPDRUuz53uhEbF5qeBy9f/NdpQSYqudfHTuv2G
EuGq7S7uEH0/vOYylgG/oSBxup+uoDCDquyYfKvDcKjp7VqptJ81+SyptYXjGAK2
JUQRljUcp8M5VCfo2nWOlh5nszchMQNdqNx8BIhdK+CdmT31Gu5gv1TzoAWwKU+F
ykvN4JDXDUVTH1gsRWMQaVyUJ8d7yTCwFY3cwwcRcbp8IrYtYPgRjbFY3dvwD/fz
7cBuJUFC6Db1zDJlT5o2ZRd9I6xlAW0zh0WWYQwOsPVwWQUt406WxDC41Dvl6NTV
lwPBc2N3x+NymdKfKOXfPT8fHcqMrFLlcqEvVvjHVpm61X3mvDMVvffoq4uyGuGv
ZzDGA9DQ1BzXVUngbVczuiU+jzFqv+rb2lnnod19zA5hWIE/PW/fTiBLQv2JaFpD
fOhnBMaIiUOLCJg+sDNV7aYY23MRnhWNIZKGhi8RgsuVmCHnE4hJWxbL9kaWUTyf
lvD+6awLmTtxka36j+DCO7F3q8qtKAMHPDZmjtwEHhI7WKufODv6D0uHrKg5zTEX
g/9JRc71X9HkC7rCCOsONddjnRZFAH48VuD8vYfyVzPNIQgPFitcnNCHbduwp85e
cvdWKPXdS1L+7jGrrP2vPFyt0z3ok63XZGWlBvVVhOq5pJaFTD8M+SBZLYvH48o7
NMLaXl4Bw0XlPRp69nRPSIaaYAjvb70W2LwLnrhRDRDJVFNhgsGuAFl+nHNem1HU
ODDEOKrstv/L/s9vU8bXx5M8+KtguRKbPaABqrcpBdWl7VolnlWTqTffLNnS73gQ
CB3MwkPMtfkmz9dDw4HQFrTbW24Pd+WVozhrXzDXZDyJiRmPuOamYACfX3HxJoh9
sfY3Oh8yclbLYg35fpQwXsSJx/C4z68BK4BF7/vv/fxZI3HQtUeAthnmVOj9/zXt
wMpLJaljJcaUlqQVnwpqNAu4PeXsZmikFT3jZcs8XeptP6HgJP4KB2iPG9I+ysF8
gS1YohQyWMkfAF66aBlj4o54v3C8JGwAOpvrp/rhZEyoTZxi4AFqIUibrlzYrlNj
NtlZnlJcVVqQAevj0OjrEJaDG71viaEDHpt8rvxtzPpyq6Gvy/41tZrDtatky6Ds
/Y0CCWwiS//K/6MMtFrerm6km/YYxP/V60picu8bwHnbwFjd4Azgu5NNiHRjOt5Q
lazU3p+60BZnw2X+jIvcAsN9rROAyw6cHVCyL8znDqBA4e+ZRGWlJeKTt3nwCniL
tZC00ahaac4bvhqxCn5FxmwUqD67ETykb2hiwp+uoKi2y/jL5QjqvkegI2JWOEwX
dygp+qP4VLtDk/29oz07g4Lx4cgu3dURCJssNgBKvrGeIlCiqBD922glY/b8NgHc
QFrKcU6KIFB/s0H2sTIsdzSnTpA5ZS4nS2Y2WETMkpqwceNw1UH+y7s74r3VSvW6
MmduNWr28rcPoFM80Ghh5gvpGQ2wnTLIlmin4bwqkCa8C044JApIHGe4LPWrFhVe
qNJ07f+BuDk4JDJTvTF2Y7wMdm6AMWKC3wp+5+tY+oOoPROZHxy2eWXil+W/3ZfW
Oj4qjN7VOs92sgSK6cvBNko0JGG8pCwue0Wbam08ZV1s9bziIaKeg7v5o0Gg9FG7
A/GrAa8IxHesfQwAvvlc4JAfRbkPt/Vsef+iR0B1IV3P3+CnQjyrYDi9YgysoAvo
m0GqD+aWOLGjzinUFMIldmUnpQlIyvWyNRn5euI5kFy1xKh23CWEyMaSEJ27Bp8R
kBIpflWfV2xFv2XP3+hpqCVnyFVbBusasss0CvKHL0s4AI9eWDPJRUhAaafgw4MS
ljCqluzkzk5oGA7WC55aQd7K56ES21zFtfZMDygmScLLQuRJegNN0N32YsZktmGz
Y6xdJg70osCx7rTT4CDBdItNLJK4QzmCKz4L/U1a7Ys5lbtEP+slCGmZV5dWqYyZ
J91O91TC9yjuXIkTfZsycEU3UU7wfs+ONTEf/5T979ecs/n+JpHlVjAhHGhUG8Uv
PsyDLjl9hTpjZ7HU2gH/9N0JsmK+aaoOqk9oAZSyQkKpKg1TAHQnSQuooiWdukZH
E2XZadgHO8tk542t8qNJ824sjshubNASGxVr1qJTju+Imj0kLgDEQ43eyMXSdD2R
6g9koQeLHr+tRpm8+z9LhlIHP4+z003Ilx6LAQPabDL9vSz1KjyTM+xGIIoamC2i
OqrezAElHfK6FzyzMA9uCazhC/ktavbJpx96NBTxSL4v+4moP7OEMJUV/4jutQN9
EjN5d/TrCmtKze6UBcyo7QoE49C17YQ93bF2MRJjHM1dy1ofXOAMNsAxKFFO4u0H
dc2fbzPwNkAPiNDJPiCleR5UnCL7LeEc8rJ0q8rSGJSY44X+9cNO3LCbNkhk9DEW
fWg59FvmDMNIWjr+rPdwIxx58m1POiBvoyM7l3SpjB+TWJA5gKzI1zrv5ZztVrNi
xu2CRHwzkIAiWPZ1pcgJ67hRDT9OymKWoDOqmGqtMXOjCg5ydV2L9GlZKykImq8O
pp9dCFTzcf1mDGMset0cqrsFoeTBgXGKO4IamfwbpB2WQEQuQ9f+DhbQqkg2d3N9
xn5/kpMIqYzocd320rQPGIAPRI07i/XTzacWJZPP5ueYPUnzZ2OQIb+Q9G8UJPPQ
+Ls8fL7OB4fCW+T6ZfQP9Pibi5C42ojB/fy/aqj5Rv2GXYivb3SbmYIfj8Ge+Vmn
JVTSD4ojgGG0FDgw1qH6Oa8l8/e0V9dXNmeWmrYn2G0oEBQ1ZQDKvoys//UMZSoE
9yBarFX4MBU8XT+Rg1ono7YML/6sohbUe/RytJGZDkxxMvWtkfzqK1osJuhsR5Pl
ptNUH+pUUv0kLfC72RwcrX9iuEmyqaaMj7yPuleb6XQ9HQYHM2vUFk29a24isd1Y
9fBQc+3mocg6zoRH2iHnuXf6Lie1ZXQdzKjsnOnNBjlrDq2v0ZMFneXY4b7R+NEY
29a4Gt7wFHC4TuSVC8JhSCBtrH7Y0RCZ/39Z3AfYR36AIhzG1cvRl0y1YOLet2sJ
p14Ur75n6OIHQRHY6BFbFHlJICOkRhAi5gp30tbWa7x4qREWWkQYfgFpPDkIlR5d
8wyYmuR/p7Pbjm08ubNZb54wyRmCa/5Mv8HKpxbN72wm5r9IY7Hkl/uxk199tK8v
uwuOHdiwiX2W67DSNDD9fJEKdOdayIZEI+DylyzttbGYRGmu6hcRgKvzk1MLEUXZ
sFS4fmGRR/nbPFwDQ7ndtXxTZgLzfCfBVao8StJSiTKSSwe+kNh7WcZbRqvfArDq
ny45CEmEUyb8GZiGN0vQoa7KYRJQHEtN2G4X8Lijym9j2rMr2k3mfFzwFaT68lkm
oNjyuPlG6QkF5z4l/dh4LBlQIytetGbUoU1yIIW0AdpvuoDvtCUVSo12pxSADVVB
1qY2wOJ/INfrkGbO9v+/lkKIQ77tunPl0L/XSmPoKtc51WljLCy1INVnAkQLBUYQ
WLXRDCz30UsOLmf3+8qJ0CJVOfM6SmkpCzkqDfCMHuX9Vz5Fl1hdQp0evPcb/uVD
5JERzGlKM8mQ8pj9jSTUfu7x1FGS6gL9NXZadEAb17053BK6EZCKbRj3kOYOILIp
t2+tRc0I79c/diX6sE1l7sX+HqxZstJPf/gpFqjfhLMLrKP6oireY1B+3e07+pKk
mWw0pZmPpQ/oVwYYvtDwFXoNDiiwloFqlJu+w/jlc0xAY3ZsydCSiiLcpxCozii6
U8VmpdUNBO6rfF7/8R7kqfgl8mh6mxM9Y+MaxD9NeMXleIIyuNhBUToWbZahBXDw
/TAQ4hRt6lnw3Wb4oiYs1QxdYSq8ylrTKLbDFG8jP1Fyi2wZCGEfOkmvpcdDz8eb
kAzx0NK9OiH4mUl9NNI2XzI7X8X+cfDK525ZTrx5lU+SrIF6h8VSaPJ/RXWORl1O
3DsxwclaZVTFIS8ktyi0VzA1jPcmlbh6+hLwtUGduOMtI7rcoZ0rQU9LXk78n1E4
h/VpTCVmAz8uyCeYdBWBvRk3VEJhQSW6JPxP9p1z+cbx2u41+8E2q4dECWACTBoz
2wrDhdY1x8+qvoimZbEYMEizY1ThsF9OdlY4SJ0GDkr0CKLIPIYdOE/wkBfCSy9C
SZEOMYGlMzQZ5kV+JM00G3h3+DRdT9d6sk7yTtdvIiu6M/K0bzBwrv1BVUgklDPN
pBH6JgBWuu2suUPNyUYyT61ufOYuKhV77tJpUB1xVfS4GZiQvzvqT+UF8wMowISY
5eh9IhRRUHPzs0y4eNefhh0DX6kyjFX06g1t+qPMPqoY8tMxerCVaF0B01cUMrKc
crzOtDl/ZqFXT87x3u1meWk84AHGDaN23eJO6VXUdkoAEXLRpsHS3X1GHT0+T5Wc
c814bliOO1QQQLbyTRTE4fmAqybM/SeuSbCgBl1VtRK6VNCmJsfqaAch4rAfb4Wo
GU2dhb2PodVjO5lM5Eb11mKqAteRzwxfXTQTO6JfF6q6SMdCBCvF0RdFw5zDV69i
Q2WBBG3YNNw9VD1KCTXjCn89c4QlpMz9Qf8smbX9Z7BgffNK+h10nQOxDe7IpXme
J7rZ/+celf2UFhzvctrC5DFmwHgLBRfQKDfMVkjHPbXUJ/I79Lxqx2ybXHMTF3XS
0Ll3u9znaQqdR8KNoGlE75Nh71/mFmAlGK59vVbQewNxL3E3Wsa6ETR4b05kO9Kj
wVxYjgy44nHWHiir6VQ43nIWRZJz15tvLoR8Jvzyob7azwzWNxNSnNLBvpm7l6QI
7/FJSHM0gihABZjsfK7niMl6CUDTDZDh8gj7mQtxtImctQX+6dXcTZ73PA/aUPeI
pdj7JFHHhOfbGx+7SfrEN0y8Io9Kny++8W3IqJotjkXTkIAMXJCPPlPhYBEKMxj9
K0/UWFykERvc1ZxWx8BbG5tpJovd5NuiiN2ulKOKfO7zowgiZMk/K5J9oxPlHF5Z
iuCo59f9VFQ/J0Nt0ozB9xq620lrqpH37NLUUf9yDGNIqenhoYgDn5LpI0Vqd76c
bH0EXGBPQiy9/5dbNtmuE7/qA1HSGxzmq6AOQm9SXywis6z9BvecDH2Ooyq8bkAL
zvUbIdtATt8BZpMImHXrg9SjZ1KAgX5PyiQy6RuPLrl9BSTelEsCW6cGc6a1uMZW
FGDPVALNBInNU0r/BjbjTjb6vhDzNk1Ej4rAMMQHzsmJgezNF1/QSH2AV6Kx/69j
cjPN+bksLC68sJbCCTp8DqJLCJHyFijBL4vDz/qg+ksCMQDfuSOFpa23bbh2Kv8O
1Byn7jdpq77nbFKg+Jz/wJ3FhOcbyDnfTBiU4rayFcIpt5iNAX6ihfjRUjlGQw4E
sEYavLmIDeJ/cg/ZsN8H5Efga6WKqh3zQdOt4XpR4lS0YAiVhIfih36ItqJ2Db3S
Wn/XuFa2H+NeurdhU7tlacFVQ9ZPV9WlA1lUJ1RRBYRkjO4dGmnsm+dn7ZlwItqv
GwAvX3LQyyqdRCXjOnOpYntnLVBA5yRGreICbW7kFO6wBqMa2kTobgc5Jc7bLqkc
8LqPUnidoIA3qX3v7phqw2UEhWzN7F3Nx3u0Uh2XA89kYF8aky3jU1WYGJV/Pq/+
ELH3L5FTeakArEEx/1TlbVtUTkJx01wIhKew1n/IoTGCQ2JNXZx3clAyJOZe3+pW
bx/sHzeQmG/2EdiImpPc9m0bCWUvFgxstbElb/uBVvgitdKAzLz5VQyJ/I/TTush
8eA4K4Zud0hQ+dYf60eDSN8QwlimPoIgQ6rEGbxZNC+T+SQU8j1C5bgiA1IR1Wbl
U/RzU5tJAO6s8+FkecE26GUjSJV/gQHj3h3bDWY2oJe91xj4Xf0dCpl7pAl1OJTD
boO2XdLPawomMxqQtKngmqUQWVxrdUMGWMfFwWdiO0GuWVsuTbEjjmGNsWGpgipY
mYcOiTyknuGmcU5io2Ih6UOk4M/2MGpMaE/dxi7Ku5I7wO6n9BQjkiDiQclqT58f
usydOCxcH19EXQ3R/CeeSrmRrxLuoGo7sjICWIpApChxGlff+ldfils4bX6ur026
iGemhrv//dS0goJYBSrwJ38x7ipy61NUbaiO7SlJ24Eli8NkUH/sHbCnhVmh2N0Y
UgCxd7J395hYvjsC7t+97xecLGdcjqr7L08aTmlr+7GH1UcpvRmNC8V9U772UtSc
pUiZMb+v+7moivA2KihMVL+vXt+r3GC5jnfWnFwg22yMAY4/tx6tM3IcX9oC0BEx
8LUWMAHqCAOb0K7EThW+WUvNU9h7zDdTHLyFxp/jiFitnQTNDkYqTzNGcyGnA/eO
6FVSJvPpgKEA976fVzxRwuhfSTlJBW/nv3vBqsYpj13yEsrTb2vf9tfJ1nQJs6/u
fJ1RELvNKjZTm/F3Z0xnYVzKCNN9AeSNNd5DHw9+Z1Dvw89CblT43nba398WxOCn
XgeaI2h1cAZJgCdjI1NvYFkbBiduYKnY3yzfzwd+2SqdIqJtXft6huGh6tJqvdvN
OnYFIH6fYQHniCDFSW/EyexlJaNIp3ZFIxkY/IaZsiTkRpAzxca6pjrf2HrcgoPU
RgfpaPnjEJg7NDYc6PUk51LxHswFr3M6cnJehJxXAjxosYYFf1bWLNfctwNnTWpU
vo0KjB0g+xswcmeR6LaYG5VIxFOZm/bx2+qy6FsHIPVoipOj2S5EjUAeHwp0jJ+U
Dgpv+Z08C9R6o9baybT1hVXrtxy3l2oZAewPyE0A4uTJ7f51XeMtJeDwWeTwFgTh
rz0SzV1YIkxFb0XLZpDxCC/bPMQEh/dFrZjti82TefKvALtvxtPHuOuJCMqtSvzc
6GhdKhlJzB33HKT5QJvSQTNHZP+O3/8c1d1H3+UFjH1GW1J8rvzO1j1F/aFXoHdN
kFLmFB8EKti9AixlsmVV4xybAqnr1UltKbq09tR6g8UBr/dSYvm3xfFltN/JiCNA
l5XCq1NJPmxsQexjdw53a45/DzOqb+lJp+VlouKbElBWxDxhRxP6nAqAb1eBCkDD
f6hB5dksDzACRiu7TcAmQ/D/9ewvPwMllC/RUEw/u+JYaEp4ki2F6v4FAqH9iqvt
3xb9097R4yijvV9AB+d9SLGy52q0HI0IT8luM1bT/wfOzuYJx2Ns8aS5umvKZcNk
vTv+j+mtHqchIa82qze99EVStS2wkcIOz6UmqeZe4S2DyE6upZTM5C9OwLSY/w7J
7ezBLfsv1jT7GrjOUe3X5KrzC7b2Cq83eLfpKdarvJkomvVbOusbVOXUpXzIpWr2
gIJhxlSZs67bF07waSwmZfr6tArpYCftYD6FHYztM/F6QqxU44eqQhb1F4brkvqt
uCQbKBjHUOm8CgayqPkuDsEAnY+DfvMPt3GM6UoftknfJIqCsbKcDPBkMZidYOBq
fxhn0+0krAH6aG5dKkZMFlJwE34zzvMWiAOqS9J/lGc/xc+5sJqCFBRWH2rA5AOj
lwpYPe5jtfydpVlLKGWfmA/2ThlhoknINrFbjseZ2+Qk17vCj1EKWfkRNaUdRaIh
uFsHKxJ5ehIYYsZTo49mf4QCS6mFH+8MNADCYkOFAaZ+u4MNQAt9ZtrjAG6QoAU9
9j1V7sMrIa5U1sLN7hH7vucQALq18Ya9OcD3rvq9MtBtv8TBBPjXBGkz3lcT3K0p
1tSufVqdkvp2jIZhvsm3JSKDP//a5lIAY6s1HJKPgUzG5lZCPnYoRz4F84gfeFln
SyUinjF9aFgDhQEF0Fpr5cCu8MBGUhS+/JxTtk2bJDeeU5jg1XgIoimowlAB7XKd
AlNNPtqLQmc/4Gr80z3OQgq/uA7ng8qtLN0SnR6WUvYNlFigKCwoI9yvVCo6DVSw
I5zDuoMIykqsQcQbh/IrBqCFIp0Jyn6AIe1OcXuB0SOyDWaFHBxTr9LJIiU28MFP
IZVRkMWC2ABATfjeEv0sPpwMUUClLR/FgpwcGLk+F/pMZWLLHnL5llBFr6zW2wRP
dLS7HRl8zMKaBSsn9jnFMfvB/TBe43M8hT8MoUEjb0j1Xh9sIdS7Sy7jZbObYvDp
fC0oUtA/zs/l3LM8utjbA1WEcWmTD/nHDK15Pt+liZjNP+xNtU0zElf+LadLMVl6
V1vpUjT4VYYFhoFT2AJoyw/a4XcDNkq06YT86ib/SYaArg8BvA7TvJbDXTPo9c5S
udvGstUq8v2AD0NQP6A/5uMb+qMLirlrv6QNVMLsej2bBrNBjN3YQXAVI5by8dB+
HDc6EXy4UdPADoyYELTlGuleDwN0fNpvOvwFWMfPvInKRZxanVeokI8swv1dSpS1
QBpGwAA0EMO69OKn/eCJ0aT8XxQ2aEQAjdFMOGKUBSz1tfaRqTyLumDSPTCoZuYN
k43dSzWYvX+2JApY0R1ItzFs+YaRABByaFGvtoAd5Oc+UFutJR9QsRGEJv6zxhzf
SDWq4CKg1VctmYTVvheN1ttcGTpocne5FMfKw23a69aBRATnCFuWXGdA63o+Knl5
V/gagASt0kFoLzBJGppTltXCP/bdIndVbZQF0y5d3deIOH4Ljfr2m1vdMYbp1rqh
Hkg3ehSx3WzUkAs/2Lwt4RYC1s/OcrSXLnh2l4xdxDreLXaD1PW4VGYzESYrXwKa
BoYtnMlqEbqPRnA4CALx7ZCwnvixKRird50CKppnKKfvmvRCkswkNqKwo1znP5P7
or/sVYdBfbMGE2BsC+KtXACnKSIjBfR+po+uk2uk04WazO+B75tQ7+6ZCGqRbgXc
F4jS2SyqxJmNxbWCtaowBDRBhEvEEFuMjSHvetcopPq+v+WFbr+neZK9cISfF+DX
BlsdyIokfcYVg/Z+JK0koaJcr9kOEYQ3ql+kt/cBEwKWnvvC58rCpNK0yDhi4piU
VjNTE0CBlaGwqGILf1oaIx1AFiH2I1SaXaUUHQopFcMKZK/vlslXu9HX51qoxKk4
FOKZ40GlB7nysOMLr08QtptnJ4q3vay7ge4n7Wn3Uz5NwhGf7q8HJVJAeqCbYwbx
Wk3IL+MhDYMgEGCiGalpmohDR8kbPjqiPEzl8ZMdfhgrJNPSAMBVnvdz1qVZdW+H
ygH84furgvtpnxNIo9dfKMAtjHaDMbB9eHwsMBBCAZUMr77Hl4IOFZQUc2dxplqy
dzu+YfJKBm2e9YSFF+0nRbRo8iK3Y8gIG6aDE+9hL8rW06HSHAi3EYpb/QbEzKm3
wmtvcUPrQRatfeH3aRXIfWP1AQ7RJ9eRjdI65IrHLeoH4uFZtj3Si3wgeGwxWijP
oOcLmBEEv7zoPCOR2+0J8mioTrRA8hdI1P/qonWmSg5KJsEIbp2thJa5htxEYkF0
bDEj1oaReGJ6lv0yIfSyIT7iNhyUBGPv+V0oVuS22JBQjxcZWbhqwVUwqAgfvciq
jRCnEgvg9n7LU16hq8QVdllanc3jwmAD75rO3HUUpxkB8WaLLgQRdLLO0XaBxPvc
agYFqr4+8x+FW28IL0YnveYUtezM06XVJizVqTh1nC51aErugk1LQgv8ff9ZLIoH
Ldh7WkWtmF5MLfudatgoBzaVHxi7w7R8pfK/LeS4Qk81EIwD1FtiARiEMsDGiBVY
x2fnbiUuAuH484IQUwJDS9ZLNlxUk9yjavUBQlGx8CcQBlB/5IknLWp06WrahXoQ
1nVwES7CSHD/2n0LK7xJ3/O1N5GldjPI7p46E0oU8GSRLgC2pCzNbrP6OLm7XkPu
wRCdCWCqDjc1fu68Hff8tBvJnTZ6YyK5x1Wz2Nt3Qmnvm65E485KQpwuVJcPhDVD
xTd+nrlsBKfe+GnMnUHUfXBPsv+rQ6ICwSBg8STfMb2svE6z/KBFbVDaz6WuFmV5
SzbjxTUtCM3AXx26JPRwDXaomPhKFsAT7Rn+rYmgPQ0CoXHRjKWiFoGKoccXu1Xh
JO136pkJffzpJeTdNfusV5k0i32FabkV/L8w+gfFW7QfbAmbh0Wlk2PIBZ3s2eGy
6PdXeewT+BvnjC980u9ZFumS12mR5BQQKLYBLl8cAKt1YDocO8NzNXvF/KkB4PqR
Ci1klPXhx7y5R359rXgvvhbP8h5foSkJT3RH/W7zhhcEfQyP1VI11Sj+/n/vAg+v
WrQJ5LepJvFqn1Gvn0CWQprFdPOWLg0N6R05orldyDmf6faXsYuZP0JQ/vsGrq56
YI6EHje/3jluKjOUbloozNFaFUP1CqkrqYs3r+pMiSu8PVIwH+NZwItSak2zKWLH
/3hFpxYhHPf1UkiI2enKCCFQorIaZ2mlyEgDt0yWYW7MI5KUvHa8uGIUD7fsTB/8
Ei/+pg4eBfvfcFIvaHZmrDJVxAdG+Kb89Ji1CY5yNIbQGriIwVKZZvYMEr+M3HMr
7QP1G10dx0pmSb1XTz8tlQu+ck6MsCuswcvkv7IsPoNlZAQUfsJTu6VlWQi4rC+s
al9uAA0VrthzP9FVq92/2iUGGHiJx+dftWcsy9uIg4jiTysp/8Bqdne/7yVo5WFm
Ltxn2bV49tI96xLL964+HccOsbYSra2aA5Xv9YoA44zKrC6CdtES4QMDcO2N262A
HrSE5ZtsPyjj0UtxEhJg96zmbgUrElLiFMRgSLPjTj1lQvbRIXfwcWwhzMqfXrKT
K3MpufOppvtOqZQZTOVgXPqiXs+PZ11pbPanzj4VhBYk6XNOIMnl+UYxrZqZy+17
hw/bOtbwj3jaLk96aPdAkTxKl1n86DfhX24AmJqt1gXMjCFMZLQ0UMo7zEYcLP4L
hGcskGdD91I6/PHfr3Ry8Ez8DAzWoeIQOao9pLOD9BihYuJ9s/HJO3Rv6WcwvrY1
A5tVvuB3F5hApk8t88OQo/fz6UDM3bwboF1xNILeHy62B1z8rKEfhGQvdQRFUfBs
BkVevBPIWx8FXVvaUQ5XD5q1VpoS1qMdK6dcVKexFrQ+QNtS7xJlOL0GwhY54tuD
gxHpXLb9RZCEru7Ys2gC9U1PgM0uykNgWxt3r3WfhvlG7wLmAgy/MtQ4qFKDIbvr
MTmc8QuvmdR3jTE8FtFWRR2bleu6VEWQoc2DbVBGUp6tswX0ycC2JeVZCmEJJWhw
/b1Cebfb2Lnbf+p8eTC+HDLcAH/aBuNQu3eOy3d2AGpaM13wU95pQ5M2XW5D4n/5
BqzSWp6/EgOTCVjfez1ToOZRSiNakPrzLdjwphw0ns8glcLUu+y4IcyC7rfTUtzW
sS/ptr627FRIAYVcD89VIWEbXnI3ky2pKSM4AOLRHcBeVS3YhPuekG+h0gvzZ3dC
4ZTxvZWbwK+xI5uRE0heQttVvIg62mTiXoMQrXSjCMoKsfjHuPSMA9l0BCZV9J82
uYdVDGNZZiraVEM8iFG8sUOd3HYPFUGVVpFvcVVelrCxEfiOxa+oOXqog3E+Tpos
dtUD/hUWYjSgASKwxH0EBxYRFIw75OHTnOu740zpdBsc+/wNig5zhrbw2r451hjE
oRPtfLgqV/4ghteoNDxrgZBMhC4pUkF58U29jgcEWoeVtGOZf9bEUmWQMdjxpNs1
aCiHfPnd4aIHX9NlWTSNFPi4na4H9exfAVcE/a1kXqQXxuecqpzBrqfqrVNvIQR5
KTQc6syRU82YdK/ioMtXZeFgJ9TFuxH1cL/wyobK2NKH3WVT4ikBgTpY61TU0wv7
rWrvE+BrRxmPlDK3WbVnfLv3XsEAYISCGHqR19dqUOZ8tk1VZA6D67gHWy9NGHts
eFO2JtcsHxrUXqas3CZSEBg0Gi2RA4zJHPedK2XJ31f4LG/AIjt2wpi9Xi/x3H+f
F7GOlZOM9RBwlMmbPeOxXEAUERpwWTAEig9pe7mppHIsTXDnYl/19kCgYw+d9yir
32j18nysMczTHZocU6wE3G7gmqv/uUXZhjrPVZgnfVdPmx2Yf7wCuO00WRdPnGZn
cglDCAUokP6WKK1jaY9b3+E5MBIhF449NQROBgLj3xkC9W3d2+qkqpF/LMpu8NBE
1pHw1rXgz4f7HMZqGWiDZRmysId1sGzyT/qAkFe75iOh/tujg/xkk3toGuWKPR+o
koMe/+BuLfD0IFL55a6I+855FR2HiPz0Adbi2WUsWh79xgNMYJY9yvJvKeWI5ULy
m5BrjJg1bRlZdjgeN0ZkW1NMFysPRFI3xpMcwFvdfwMDGIiklYQT8ttnmQER35m9
5A1Q5AUgf18pcbEfvxOvVWPeXnmHmHqucCx3IHLIIXjli9aaj2U5/9A6zqKDnIaK
R84yxmKtcxkg/PnQYNsBY2J9iB38dsces1ibDsAT/GmoBZzubsmyh7MmhHhfQxUT
4DO8tG7w+vCBW7YwS+ri9FSew2dH0dNxb3TxN27uAAJG0IQ0MPx2Tmyj6UI0g6FO
9hohrHwFb8x7ix9D6Bzk2WuKQB9e6pOAEYEl/RwcMOnT23VZWAZQvsHof6WA63TR
G5sUWjUMSDEGT/WRXk8Hr7FZFqCFW04oq3yLnhSnaVosIxKqDV+BRpUUWD3LgCEP
2QezinTAwm7tZlViBh3mFVUhKsLzb4e0YFsUPs9koJtoHjfgvw8XzCSu859c+5jT
EBO5judr/Vhxc2fJq9OOQzdWxOwK1XD1NyHuyg0nRLcYfrKbwKxkWRraRiyibuA4
wI3fXPUzn5RWfpmRel960+6brY/3npXvpRpK89ERjA9nA3u9DeMZteVjI4LrO/EM
ilWkwtrGklA9PbvnQ/+evuwTgkmoZav4UGbgmgH406yUIWD0fog3SwZSod/ULwdd
yRQlPyWmQkrJpinvXl7LnR4gtwihpFvwLvAPR3I1R7me4lrgyNxqDCwODcivsZnp
hLkpa4MVPP7ReUUDhSLoUneZXTPzgB1BX4cyx92ZcTY0DQh8Az532AhKnMWh9gej
kIi+JNtfljXYZ6h7JG9oK8fcxPNOP2xKxA2rTmeEq54pmH2i3G8oSV4WRq5CNJ9e
g1hqlqfu6ggmfH5S1cCXZNA8n7xBEgMLzUVmBbeXOa9foWLK3ENWxgMiWFfCnJm5
SIyYfmJ5tEzssxgINxKZdVhcJXYaO0GmeGf8ccWqhla+rgMGagdMnp9a2/YCSkX5
fRetlr+kfqnt5tIMNlfqm5deU0En0dQ06inJcC7dklC1CbM0ML/amRaNeq7FgWXr
HxPpCgco2eYU9R9wYET6PHdq1nSHFCZNsT88zSn/fbekziNFPicGirQwCkm1+8Ih
R6oAJyPmUyU/HnjP/gthf91MEmxPFfPxaRLzGvPRdvF34AH7crubmpAMvGqDSCA7
cYKFGOmxYQc/sO+xhT/EcUZxYCKdjmQ+K/axAQsVlHx3nUpwPkogZHC3AOOlWgrX
6QUyJJMd09oDSwgUykc4Z9t/F4dcLTiTuw20rAfbvDBuDYnQBtzWAMiqS63s+YT/
gGs6Xe+VdlCrf3toO7zAmin9CjoZMJhaT9aFSt8MfLfUUASGM1YKU23TshzFuoqf
6B3ZHRqsAgZStruee7NQ+5e6oK15gAKjMfagbv8xCwViCWWyd7W3+mHOQ4xmgj/2
u+t/DcCsctgZEIf/LZLA9HnMdDfoPNpAR81euj8xiwxBOofp2PyVmVB2OgGjDa1T
cA04U82/ZTtJJR3B28Uh+dBNUSyVcovkO+vtdlYRHM010ovXDFWG+z+jwBExEuKa
vFW3Z15A8eu2fgU6G9ag2KPXgkr0j1XfqDSOej6BWZ/aEBCCGL2NuvMVaXhJASLE
8QVCxvIsMM3XYL14jLR/8jXgMGZc32KCvnJO0ja6qltm/TrrB2WgwzGmAa0A6dKr
+0ls0w025NAjRx7CTTimGac6simV2BYXL0qdBAgKADVC4FEeGmQ1HymVnUM4X/hb
bdz6fsggIzuUyGs09I/IwJ9ALzx2+S1+3IgButBQnVDBFGSG+RKft19rxXfP2LGM
FIJXLpbpvhIAz2rtjuQWqXV2p+RQOEqP26PsHJFb7+2Ufzzb4pPndBNWAYobP1d1
YoKsvZ/QcdchEiaL/y6j34SXrJRq4uSCDtpTOBEkQ6gmk5mE2OSpchwnlnECtgtp
mdFaur80Uw5t0gaXSj/SxUQs0emE06x7HcurGf+yaP6dKk3ex2sMlr+6Wg2HnyHS
nqCRPd7PLtf87yQkEUm1X8M92odf6m/hcQiVdq/1jwbDKhXooBiLzrOCTwYK6jfj
CIExuRPMYWfgTw77h/DgXsNmqG2uA7SWv4KA6d9mcF43M9PvCwFD75gcggJNNCIN
DIUM3wH0lyjUjaMVO5er4Qr17c2lad5Yo10FobZhFKAl6YiK1NzwVLDnqwcG3R5Y
UfwHZhGPL3+qmQWOR9oShfdKpBh7kjjG84lV1LiyjqZ92NiXqLIUQr8TURJVEiIo
P2OJ2kAsVFVwn8dhbtme4y5lXjdt/Y5TRUhOFEFmVpA0SmSfUjyX+sMTMcvBH3tS
AqCJ/mWEgvwgDwvXZQVXG9WANAVJGWR9XmTJDL6c44R9pPBF2CtQEutQwphcGvqL
YdqUyF9aG3i/C05KBMLpapqCdy1/nOOCPS13n20qQ9wYE8ZQEyXFwEQf8xjPS6Je
qBO6/17n0LRqdCe8LJzmmlHHd2+jQStdZQaktOn3jgdreEfGBT/W7Nxgdga/X9Yh
syt2Dc/hMb7zv8M5q2O0LtrUBiM44XBEyGWXi4m7dN396WqzZIvUxqjxJq+6K+5i
nvJt3lL2al87nzBCAMwSufQxC2v0uR7b5/oI+IS1NQwiAhj+0MPDkJZ+iF/RhfOs
akb4yRulqML6UXc1ltbl+UIVmSpJ65S3OOAtTAV3+ahbYhNlZBx+VQwFZaCOR7F4
a77MgSDw3MFLPm8ua190STW/52e3WKUbk2DGb5clLz8LBGLCwO51lmF80nzUHRxq
/v6oZi10t0WpS+Y9gygpymfgrJXqGmA0KLwdrSphvFGIUKj0s52GjvqizzY+FfqD
gLnTZu96psPImHRNqSkn1nbeFtCk7FNwAg5soetGcHo4+1A7vf7hmIt7lxnf0ool
X5hwnK7JaR68hXPOPM6/LkQQ79IfBBvAwq/BN/Qx2ttxk5h8qEOwdP2Wgw3iH3B9
vaGdMJSeqC33D16HO12d7Y9aMk2bOMAJwHQEj+A6ind7203cMih4iiGJSw86otMY
Tjq90zBdcF1CkwJ2KJi6H8qeYXFltILWok5z79p1avU3+6/TSZkxdNCefCmebO8/
KLYXqslusF+YZpdAz3Q0X0h6YGShNAi0GEKOQ+kZL10lZlyrM49FQERpqLBmv+ya
mTtLHOrE7DfE2HfCth+5HlLOSnWE+XdVJdiKEAwuuZdHCPAwDI3qL7Fj/KrDwjya
0cE6mQQN7dbXiYa8OuasD6ztXwx09uk9JRmWDfVMDDSR1KI1YM2zTxy9qVRTRSIF
Ds1iY7JubtwkQI+164/nbCXXrkOb117LSKTA1GeYYK90+kEE/hTcPEkdN98dzrnn
+Wv3W4VkDHOx6HqAV8jZJ0zJGCt0YqK5akSmpWwNsLd4TEBgrnvkphx6EwYGL9Bs
nHYo+vNU92tLNgn/RuysAAZxAWxsoDKJ2nGyNWoPHuELfD5/CIBymw/mFAiW29Jg
EvbDflk5ovR9DtA72PSjWRBls7Ce4Wal5iVX33+KcUI1hQOFUYIXcF7YTGXlxfVR
eAQMHQazT1CtBhztK/a9y8jhJ88GMhXmecFujuvlsgb2lV9lvDFPIm4jXZEnLwab
29iXf+l3WUBwzWEVMp1jvZjtbn24bJNu2T7/CBNyy9g=
`protect end_protected