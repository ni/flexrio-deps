`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aMReDmrPskJscpWYThVKVItA5gecPPZO1R595p0GoIq1TSTG+UxXhmmUXc+VYHJ3
u/C3EW5qePLufxmXxmhmDnr9U8/cYC1zLfk44v/2OPb1TBrTsludEDQZdGNWeV9l
cPUMSIfZ0dHXN7L1M1E2XtgoTWQxf3VDHs7B7lU2y9Rdm/ibz0fWMow7op2nWdD8
gJ4QlNl3f9Oiotp1p8vz9RFzzZOF5gBBslZxcTF5+z4qO2W7+xLByngthWm+exIr
3Pzy8qyUo/m2DDwOz3VJSvSNm7RUq+0/yJNOOz3jr3j7ZyCj5OqT/jDAWjJSMH+i
2402Un+wDMOQxi21JLo3cA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="5R6K2aWI3OdbT2A+sz4o9+2XAInTqB1/cSw5W16RnA4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
Gm/2BIZF5/H5qen8uQizPH9RftTuEE9mgEOF0SqeOKegtP64CfvEUnIxj/ahmIpA
6xUR2v2l7E5duaLZh39Mc1GYsfqE91NCPU5whLaBPg0UuX4cgTkO4cYbW/7yvcrd
4wavUfwXEp2VSiN7EVxL8RcZTSMSI0Jr/aojiilFqVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="TEmQtJ1Dsm7TOzpJk/CeTSSFx/zKExk04H6I8sT4Meg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36704 )
`protect data_block
nvPqn26PC4XWLLQG0Fq8XsMTlhB4evbpiwGjZroFFLgtNlE6bBjdtwWsB89WW4j7
jNfYbKN4sBv0hDeMH0AAR+8g+TCqoX7yLdIUd7aGwBUZJr6FdDs2wTUxRkXFYNTL
Di/FaDEab+b2U6o3pOQ8Z/wb7+AGx2vIVDuOvNk2eKGpz5VWi0wBtyZj3mBUn20G
kLheJqwmcwmJQrBlBeY0xlsK43NS6ZZxkI94P62ELsSWkAqTZWA70cb+2TXDoahb
1gHkN2GjC80MpT433TD0ibn3Fpl5GPlzywv2CPdEKRD4Eb8tUVDy/uO+twoknPnq
v46CKLpdNi6NUQlUNy+UGFISKlLqbuYdziD3Wqdh4ZZgrNJ2+81N+pg9OIq0e5P/
ptvemdEbmNxVRp1gXDy7IDOE/yWafGfUJidbucuIXHwgwgdJb+z8uGwLDkyaItRT
74cQB/3OL531wZsnzIn6aqC8Wx2zbMaE3tLj1SW1vFKAUioqKWGkRGw2T3PUNs5e
zIobICUec/A9B8MMHZj04RL8y4iwxsEgWVO6SbjDxQ/ttD/IPk0jdhzpQnSi51FR
daqlo3MPROF+Lfxexn6bS39V6Sv2llH3BVGTiRPh1cv8Ip0hiTDZOafPnZhUFKu3
FqKoWIWtQj9zv3CMkLxSA3dROmP9bEUcXUmysVZLnQc6CyzvFUD2InE2UMYsdgmn
49eQEVGJKWvpJAzPUFr1OYiCBdyF3SSKc7ki2B5ItJWHD5gwSYSGDvIwd9gILfY7
GsChVsNnfNjkI4oEfjjkNYH2TtwvQxHXCQkKYSmrV9PfJYBdv63nUzmDO4gdDbdH
hA/QvnXMiRMcon2pNx7mGE+A2n1zZXUOnbCX3wAVxThHEV/nHS+GClMwu1OKrj5p
X7YOkDDhNlbYQCJ8NBVfw3Lw2yFwIS5KFRXSOObjHndw+5qF5FkUmoRHpZL7Nu0e
PosJ4OhTUHlCg+fOAdlhGNWPHz/30B7USCiU5HDlaRWIIcssp83cgYkBvpDaTUIE
rpdS8j8PjkB0aSZKi4MNsYhKk4IEFuSQr6nnVYfPo45jofqenE+bbnH+3PKrXfaL
0E+i2mXdYOSgJs1TYHkKZuT9ggWOnCJeQxdRHVQz57kkIdCqy5H5jRufH0Xuq3XQ
Q+kjv//eLunMD/PXPCPUTQDtbNkBmR6FuJnQabdRr7ip3HE7NQaKOd7o8aUXnFCa
SJcDMqyv8E1AH1CbShBiaSJLRDqgHVpvczfl0B+JwB0R+7cH+GH2tClCEEAQnk6Z
dhObxAzDCbNj9iI/Xw6sDaa+5SZgnCmhoAwNs6BTRH4cN+3vKmQG98PlaEVA6iDC
t2/H94ie4RkLONqOeTxIlVWml8BDeSd7YTLP+E5MhRvDXqzcQyMKkfWMDe7cLJYC
lcl2Yqcgk6b5r9PfpR1KCS2kMQjL5h+Nw9gcEaZnGmgHRGgLXI7qysbcZhPhQ7CY
Vw9c/S4OgHLjBBdIzo+jQhiQZTkBwRD/UEPYO2G6HkUWFfQaOkn9x+uVj2LDYZq4
qWDUmxYhz7C6ppceGhRR65h2cP/KrIVXkmozAWObzmH9bG+T1gSOF4r9YOyNHRS1
K65fgHM7EeQyy+T7blXkvoHv5ZyhonqoUmRs7yv5/rx3BD4juFuht/h9BB3mXCjk
dK/koXlXudrIQrhlUDp+6sgejoPzMwTKRxuycF/RrEhRwGMaPvohuS8O06f+WvR5
wHhCjMDGSE5WYCHFlk9Hkqe/kqXf/i0N6wtsSkNJInBkASroYRyxr+KAIEXFmGri
W0+f4B4T6h480VpkJM9v/eKvfxp63KdA3twiTOrXDOwlQ67tFpVv28GaENMF7iEJ
41oScqf2p3OifIaNlMqfSav9MJ4tF73DZzrSVEGTieywIHjnSBJjYz4ZQwhBPOQG
QO0uK93eGAn5bPf97MYJqgZrK3BTfuyhLn0sCEjyaxN70yAW9vrLSEdTYAVcjm2t
H55hiFVMdcZrg46x7PDWz744c+tAFJV1N7cSgv7Sx+3z9IJTcsOx1NVBbIZAj0jc
A8hdiD9x+t2otCSNt4IKmZjpqDqQZqv6BbYGGNtsTwwqBZFvU3bBAc9oKQLn05XL
NesDNBewGRd5oWwUq8tGnDQjEN7Xw1Q8UfdqhK8ea6xj5ARPHFmZRmyGCK1K7e5E
0hxPu33sqt5UtRm7O4pZqT7FPkZJhnoXiHdDS4oG/P993Wl84DXW+LJY5eAosFxQ
1/EML2aWAjq7kh38bJxZ3GpqwSjq+OHYkO17DTqitit3GLgiXoaERjU2VcGgO4WI
jxeJ8+QHaWuFh8p3DEmkv62JdC15e/4KM2aAYKPhenJocsBGH3xhd/Ei9ZIvFZGW
zTUeRlYCFbNuABjNuD8izStyvSk4K3WXePHBmHOEISSv4yvnYcUDBxDKTrXwwbRF
MSBTKl9PJTKUzBz4SYUgY7Zs7OqCisrPL4UK1xX/2k9StbKPlX9HkzETjJf7SmG/
AJKboAg1BKu4TMBCA92zjfJdgcMMd1x7s45iWP3hKb86qDoQ7jKM9zURobctshHD
SJtdy/t3rEp7qzxK2kvWQDtTKbU2uPhRlULmqb1+p5UeBGejmZIg3hwLbMKrskSF
Jp3arVN9O/Ku7wCw8lxguDW5hDkekvOFAq9seaPTMGYLku0RGR7qRJQeuIWz9uIJ
PtphBDefbiVwMo0tw93LGwmTPp/kZsOtsEvyrBXYEPH68bBRJMdrfJgbo4mSqKng
F/4iMFhLFW+qFNkeUmzodhlT34QaPbg6n9mL+o1K3dXNy/Q6e55Qmt96Tw9Anwl5
TYBGqFdxBo6/Ml+GJP1v2ECnyyDBO9h76k7voZpqEDpcsoaJrZLDwz2JicHBYbjj
kvMjDx+HkDOFTqz6hV+bzfR2NzsEsw+F6nertllrNs3Sn7Gb9JU99AvYj7WtJYh9
wgrQp4K+li4MbWcSlHO+J0sgrjzr8wpvGLUokNpsjouD2ZtCNg2T7eQUBLdfq2k3
PT/togERMvUE0vqsbLharMpK8j5e6OXq5FE5oL88RW6ay6nW7041ldeBc/GmA7pW
FgySK1DTDjJPTEUI0ACRCS0CzS0lZWFGB2STLuULZWTc8r7qVdgWn5fABUleJnvs
J+L7I7tCuAaPVp5fIta8kOeclQQW13rg4+zvYK7DGpgkumXwOcgdDzXu+hZMO96o
jHqbRyskO0H6pi0GRC8v86N+VcfkFudMIuM5xYn2S4W8+mZafiRU0sr/bN4L4TC4
rrLv21OGeUBpv/I4w9NPk2ETY55bxdedpn0Q3Yl6ALAYTMGjnH9JByDVYlwqObo/
g27VuW5TlHejBsK9PnQ3WJAvGLH6h5lP45Z0/hxj+o7ffSPOyHSbuzgRO7uWeFOW
PHiRC3tMa8IJtt0ux6wS83Rh1GUIcJGD7Qy9pbApQQ2j+wfKyC6n3KmtoI0UmpAl
tirufnYbyUloxdBIdkVznj5rIu2E2IXkQdXVX+pnDikOq2F1yZg3wIcEfWKsmrTQ
VH8y2we0awpDOJ5DO+At5ofTZGhYwp1qFF3CaFQCgXctVIMO8682RjsOcONoc3e3
jP3NxOn+BFeT4bblXZfecTbaiG3+jjpP4WDGpDcQVv3EyCkAofQFEdXqtddHZxlU
csYz1bySi4X68OMr038048BIV0Hbg7FLcASpH5lZNdpShyILMQ4xKgVL9HB49p6n
x3HdaDw6jRiNATXLXvvSrprbQpJl3Cd5A74g+76vT7xajBi1yKdf4/UaNt/3I6Ti
pSVq+WDLzfyjDMPnuAd7xapoeZSzhdFEpp4m30n6ckmUOTXtzJS4DLH8ddpASLrK
cN4CIyTdcPdSo9/LowWsp3DMD8KwuOAVom/sDbiV4UVCb0jTeCieuy2qTVx95wN+
CZA2uYmWdNoKgVJ2QtsIK6jtqKJHWmX8nkPcrpRUNoVapmO/VVN3P9GRcNNGKYMV
8/oXPtPOuKcAq907p22NapV25X+NFQCuaqnLirMezA8U2mLGdblCQjiJNOFcCr9G
SAnVrZebMC6CRtl970rC42BeMRpRaieZdpBGjW22lS8djEfPAc8GL2K3OcQu7e0H
99+eAfLsee+wTPgPp1GkQQWpQxx3d6X9JQO4j34Hcl4Bm7X6ZzaqJV4w+KUJVjZe
M38ZdAuzspvmnxIO1KIbGPuHB8hInpR0UEd4dILPJDvKM+uaBiDwCEW2Esvblz90
ZsBod/wf9NyycQdvInXOyRmu7P2HKRaQx63XKRWcvgqw+5WizS+eBLMazp1XLKky
nO/aGSElM3ZmTqtmRHpddRm/qo8xBE0PTQubf+fDl+d3oFhngb1TUbfJBhwvlNlC
8NV2MUNRCVwXBo6b1gjnJ2tWdWQDuBi+CJnXewrvoS3kgKEdwFmS3FKcvdQ+Wq1K
qKubQAix3khzQ+gM95FVyIsW9refvzgjXWOVIaanDCK7mD9w4SlYkvQrfAkyWFTL
YnwH/sU1xhS8f312IfJjuagxUnn7LUZI98Cy196wl+nj7m2ERsJ9pPwUgvgozc87
7X0pWKRYYzkQrAd9HwJlo/PQ5UHJ7NPlaAK3zBBt6OdBn/tfMYrpeh3q93Nz3B6r
xRz36dSiswu33hc+N55X54v4uac1Dmw+B/dOZoc/wYhgXTd2VMkBJ1a6kHuSrZMa
E6203YXcVHy786xlF/0m2zsYf8Ir8UTsa4EgT6h82REXSa6VyiWfhHQkqcpqGWrt
PAxx8A2g0ov4ENX3+FaSFt2YOu17hzUptbd1NjVFUW1bnN2+99I4BCfjUwvfRQUG
6VmzMULXmK2zQr/vyisNNvBHzQ++AgRVtnSxvTzcnxIHAtQ4s6m392xxK4JpCRDQ
hporQ+hImuincifIogkk0/ff3WQ/UBOGbkFYGcgSQyY3osvD8bqwhhEqodYnEI+E
KLP9N41iw6+oKpeahC4HYDAkKXSz6845EDHvzLfzYhM8+7MQHAwbJp5GO7Q8+T2+
+VrgLu2WuyVovFPS/fPdY2GngiG43tMaVZv50kplMqqgO+Sje8cFuJ3bRUkLSXNW
cMJUGuc/yHByOnPzPgFruT9b1JQAxlU5d2+qMd+nxGHJWYPyJMEBhF3S1mdx3Z3Q
i2sIwyl8ut4MtR967Zb0+9t9SXglN+UJRk3rNfWh2/jfW/neTZBIzseN8VE9SWts
4JA4IUyYCOo3tEIAsrIE6vluQ0F/RMcnfrqi5+WHIbTmfAfT0vGR1f1rB+RODHJP
Q0lX2fRE4viUxMMzdfSmrW7kgie6IdMipSNnT/1QCEdt1fWXAE8/3Y79HVLNxMnY
NvrXTTn3FslSu/xX+CUo2n0catjyTGYT3yxr/6fjW0oKfNvRE7Ha6Y3piywFDEZT
VBgL9JjIZn9SzA2+oZXTc7hUPx+lLjW6YfmAPLLMT3f8I3dDFlJmvtGbUhWw0XbZ
ShGHn4YwGoK3UL5N9lWI2UG7QUhfkU4tE/RbfKAb31IuQ3Lmef4tV3TzkZHBRZMh
wxK6YzvY8CpnKtg2yY5vJsicq5wGt7tq+VNWG+4ojbeZXtLsIiOQin7wIILAN2Ta
FIWDWLkHqDvD6ekTYFWIBx7Mv7mkuxlfOCNj1aUtn0O5O57NYjKr8srT8m043Nnk
bpJSIfFhNYPjDIiWQ2XuSBrwZc1IBGpv+T0Ky2zygAeCogJ8seB27oiRW4MhE16X
pWaWvqfyANawEfB/CsUvnvimpg30zjWP7hi+vXiG6j5ZM6xwE231JY2MotUzlRYD
Kyzi0XjBVDklWi4tx74af8vhofTvuMU+gXHfeXbNLjl13BFC0pPxCSeoBt1jgz3Y
Gc0hOoFYEn1VC8D7uBEo6vLJz4YXcJMAkpaBBlomh2NgEDZcreHsS2c/rEzFmO5Y
68KGMyR1fiPcqNiIekxJe2MGr8F5hYNrMgMMdFv1SxOELsoZUv4GHO1yvWNKlxPL
ffodbWI4zdpdH74gq0lJAkCmdzC0wSiEXBVC3/S/TXfRlUSuEuvaKHv7wtQKLmDv
uJ250rYLSD8WhQ+bRhAlf4oy9tv1II/Li9x5CO1Ax17jT+PIp2i638o2kPfSMCsw
k819NjdXZowtrHhopTaY7mzSG+3DmxmdthodR3PydtlpOjBEe2ffHEPEZFOvvO8g
lh8qT7HJZW+qjcYwQMKr0n2BrZyALar4jWZ0P2U/4b94dXI6h8ryCiiG5F8bTuEN
/WPvIo3I4ZyR8Uiyqn0nGmXNeMjwwxpjZvlsTeEfx8pZiQiehLlJNWsKP1vRl05N
1y7C9QaS2Tni/HrWoBREKz4VWN4c/31gvHiMqcKABDCwGpPAABJ23Jw7uAGImzAN
H6FuD8Ade/q998hyIVlFrAy1m5MQE9422yaiqBnMgfunYslMy//qgWL1dUOgWZ6X
7+Th8oZsuoWX2UlY5p1NmAJeu0E0vq17EN3DJCceTXzGuZsACOC3zG0jvNVyX0Av
JXmdZeoXFCIs3JXWHS5zSmSgXD+vesHHdF5adBQ0L6DcTolggUbDaqdJSt3PSgjV
IFDbnvyRsOmLc2AKVROxi0Qn2LoTNeIZijwJQ5bLEjV5698/t2Q/UhmFce3kT4P1
YHD6VNQD/jO67Ja7QuLjaoaH6wIAZfaGtEldHH4reoaYsA1f0mwZDsDD6nfOpZVA
l1urjDLoh4ctaPt2eIhTzRL9TzSFrq8cWWlZ2vTzGojJGCfaHU/Z1Uv+KuZtMkLM
5MaboQEUF7XaOjLjz61pUzDFaRHays4CLDGBPvWnS8uE73uE6oVn223DSGYDhX9X
Pw+uI/Q91z3/gM4sHokbwUtuZBTPw7yzT8brt1e+JF2/lSeEN5PU7rCJgE5cPXQy
Fci9vZAfYG96ji8nYC0MNB04CdCIAG2kTmy/w6WMu9fQNo+/f9A4RiL0xc+uYA5v
m6nTZf8NQIqCcTp/1T+RVAl4UAIAyzGqQF1UZwn9m63tSZYgFj3vk790kIC4CF+r
B3w07QNQquMnfMPkG2f+jTSQD3UNy8YzTZepJWfF0jUxyQFucbhv/PLdbkP1vO8X
NM/rcoAStJra5c87E+99Ot/AZ59tGZJEML/Lp/urIMxQD7HXFpnezT3snLfrBD8Z
psXDyMYT7e7HBkxPHhKY8/XxZcYxOO59cVeIFLuqwW+NmPIBPsGYTaGMhoI3xZ1g
iJGrzNGzoIXMEBQuWE/kGUJnzr3E2pMIJHb8xk44HVVWAif+wG98MbMJIYI58CUT
gB7mHj4CVV6iUnnJRN1zkExtsYeLgRJkfEur/4Ea+mAQbtdxHnvSr3tZSovuvTCs
6nY1Tm/G9Kk13Gma0D8+j5eGOaw64GfN5bFr6EBkUIJRrW02auJIjtnUEGOgzt9e
HrH7jX9rtMnx2WW+27h3eGmtmiIUIuoiQhnBKoTOyvBLzjgVTL3/f5eoH1/R6WTC
+vhkhmO8zBORzJzUlE1elHyUTN1LVEJZ46DCaFhLvi8XTiIIIx6XtDvWUIFCntzB
hWErPukXoV/ydbsrBnzNx7K7JY9F6ONtSYxdxzvf9zZ3O7RBG2NpDJlY5mwqoIsD
fQEMQASgRVn/jVX3qXOkcLN19IbaasLKR1b7jl4Uu8x58hgy+HFsEqdbmR+HoKgL
0SEGg3yWGlo8YTFK0PN5fORXFBrC8DtuHJoOghv5I6pL7RfOaoPgXaCvb2939ZYq
SIa1aZa4jVn9XYwbbA7mcaB4EKLQMYi/bq5HqdvH8Zfxr55/ejDJLD7df6Emct6G
iPOOlx/DupoV8ioEn9kNnZqscKMZzGlkE5Aq6Us+a3m8w1DI6pN15fZ+cBRjJ7rN
J1H/tqmjx67OUiqcE3K2Z5ICAt3BJfMLdCnDcMMR+dgUITG+dxDWNu5HPdn7mQt+
ySnEuZTA5M4iS6XX21vPoTvU8s1PPkuvZgIOxYsZPy7A+rtPPn6nXianetXBmFY9
MgybSKYbrK93tRnzx+Ods2Mc+RcP1hkVblVxX+xVhI4ZLAGqiKXzkWmuVWSossFB
8xgSOFlgLuuOFNhMbbNH5/UnFAKe1CDkwz/AA9aE8HbE7ViPoWUqwsQBjBoqPhhd
TKObcnXUsJTR5mCGDgd/KSINEjEtEvAdZNcy0Npyz+U/ahDcN4MSF6tK8U4bLbVr
YNfAvftg+UTyB/9jermCDmUR5ejjhMa47gt57xrLCXyOS5iPIuq+1rc97NpRBYuv
7n+AdWyiO73tneGpH0F9kr6vJDvIs1l6Zd61+cR89kkX/S1mKvy2Yc+pDL0FBzyY
/37bFcoeIGKLmm9djuUdEl/z1RmkHxp/SkqTFHk0Ozdn7xY4bRYVA7vwjJd6hIIS
AJ88uS4pa+SSVjmn6Obd5r1RyMfG5Ujk1Oi6KdboXp8NDxvuqIpPCWDTnHYMKbi4
Jt1roPe/mM1YlkzvO3gQkisup7Kwyl7sah8gzmk+9qvEaceBRBREHt0+jDMhKrvC
j7gDHIiU1mrJfEEpbNq4ZP9Ig/We3AYlgBCoJix1jUQRI9TY0s2dWCLnIcN1Tmr+
kjjW/JlNwe6/6rozKq/4NImYqhRqTzUpHlrwuP2p6JfGLGek8RgVnKFs47Eoub0a
Kipt5NBsh1o5AIHXNa4fu1QcL8Oi6XvCIhPCoEQvS15VDQLaoJ8HoTdJSPcDhWA4
DYyuFtNJpEdRJtpTqeKEkGCdU4O3LpQVvGvQsH+N8XqOm4mwCea+QVTcWFhjXTM7
tTu5nrTYGo7D4L1GTjVCvTKF84VUiBQYoPMJFEkT48JwG0SgJop3/H2Fl5ItvzHF
4TohID3Rz8r0EQIJVCkIfF8WcvVPMcYp+3vbrHWC6d9HiPmnxcK2QNmkG1Hcm5Fx
qgC8UGm4Co2k1DSJ9znYhdclzanu5qbQp8Dsj1In/atkk4XD6v16fMcwFYY/NUKq
X9t+DpV3gj6nMnH4iJM6IYMBYGgJJKQyPcxT3c+CXmR1Q0cbJB1+AuQOVUBXDNnD
/VVZ0c2BuZ08iwyZ7TuuSD7DlvVUbA19Uo7lICJGUIDPbj9gjkOg21266x20a2Lc
kKiCkJSQMLu/rKmJCnaqPPNvRJwYmJ3AvHoI6PcbNfpDoYgnLLC5BhQTK5inFaeA
69rWlEIiodkCyh/S4MAaBSHPIGdq0LCBXlBTUwN852MMPC5kxtcQiOerg8546IWu
uQtncN++C3Nzsv3stuFKdV0bRzPOsG/dAWUTVV8GWzUC0aGV4YvkkGfSHy8QKiAL
J/u/ynol2pEKGHIGSoakgkKEsJloAd0Poo9PgcNVHKjKY519g/q96uDDT4oqor3Q
S8xvR8f9bsf5T32KQ39bYrQ1T3Y1WUxncKYcMMjWr1gygyPViCm33YUfTKKQGnDo
7fL72IVRXAhXsgyD/v1rJe1iR2kpdT7qXXwLIsRSgLM8CHYzkPxM9kjTxGSMJQCr
RbJb17vNW7EHY3sQfg/55xH7ocZgfARhkz/pFk+IyKCyg6KHro1iEjsH8xJ/og0O
urnvbg/ZnkWwV+AwAdFrGgewRH6oOi6k8swq1uxkkcYRxYMe2kZCSnUOOTQsDqJ3
PadifeoHw0/rLn2Hhh3Ciq39WEkU4qrk+0tmSetCYofs8cpPl+6RAZunbFO8eQf5
JYMrxd2STPMrPjZIbi8bmKWu9TP4BU+os+uiqF9s2ZYUs8vwLUiMOpVopc6bapnC
OmWtBnUVcdOmPKBRMBW8Ve7DMRPwLVyhG2j2ojPW6xwAZSROPC72EdzyzyKAHbYK
GFJuTlmPqs5GdFuUurRC4ViKI0vyNuTNgoQk513HQrB4Gfijo39kvXFXrMtOAc8u
F+8Z47DjGdrSI3qoCxWQ++8peC4fT05JQqFVIK7Qpo7WfD02+bkaQsUyNiqN5G0O
xmWjA/OTf/8cAraJV4/nE4xrsgm3mh8KqKNjwezNDBc3p4OHeyl7dRtEIAkFt58H
5opdDjSn9x3d69ytjZSLeB9QGLr2bT1TBbXAhRfrRijeiFU1P2qiQ4lIQV6YJBZO
1DMq7wIYK+K78G3hX9qClBtHM54SBoVAX9hMvcJypBkbf1ThNbeGMVWFkpuRK/Fx
kFWGKJvjMQ/jzdrm83niWo3ZBxNqGk6kTNf6/NvCSJW+7dNER6yo7Im0BfsNh3Qz
5gtefb2r2qQN4sUQB1qYBMudeZ6JNHArMHV3kTK7KI/H3BqIEPWN+NTcRPxbVe+j
lffFXWXdGBhEHQ6IIihNJRwCwpLAATvBKh4swFaV84EzZE+p0VKChjMzsoKvle3h
QF+iQx+lFOdUrc4KRhVSSyHtjKEOJOnbNtzCwg+vq428ZIWpJJNoOxaXTCZMhv9k
LOMBnTVNqR83msSZwkO/TxHu0NuZBcedinTQcvxXc1NbovhlTS8IfyBX//utWjb3
QDaH//xvlWFrwDpgssLlvd5JWSNRxEIEvjanh2/gBb6X3TkOQ85MSo4+ythxUZGX
zdTwJ7IhjUEwxEuvyMRMLndxlX0TdTJ4SBKf/Q2Y6Ye0yMFOxkIoyU2gp4iE5VeH
+kOTdcOYilHoHPU6ZC7HDJMqVo1e4CBhv0LbhAW8uhuFzXCQfWpTJ1xsQnMbqeeN
axSezy26WnHheB7ET3S8D3FWHU23c9mA/hPCFeR7vlaH6ovFJN+AFDTfNTEnQBuQ
W5uR+2WyIWkkJl9h2+AKy/wgDeE/wbL/iSqhqQ51bIgOLaAXBde16dIPPH6WcRL5
CNnjAR201hdlJqYRwf/WL1sDFcjIBm8XGvK8bxf6gl5rDG45ni9IYmKvFMnnxvpB
gMSYO0zveTSgyvTG9Uf+rXBcmhs4mOJ/XB+IdvW+UWsxLAozcUiasr2mJwl87HaH
1kMDo9okQmoNxNKCMdQ9gzE+fDXEgZirWux3orwC2+5Oz62zjmygJBZB2aRlIsHh
/P+ffbaj4mzpKTvgeM+OQKFaQHpS8Ft43ZCTY/BUjMjAs6Q+jKxiMxbRfpytWhKp
nAXtMAl4sK8g+SmTCid4rbqkqmPsJAidTVlZoUnxCQbYiXeoOJ83L0Jr80QX3ujo
DHyyucYYBUxAVgRDLmVyEZFwDTVtvpdQ9QVFunUc/RvNYgxqQI0T3/ehP/60rJCh
pKyvdiFDGTxg7/1QbCL575z5SDyA0z8e8w4NN3c5fwVF/ssJytafVEDaaWji3mEB
+4KCa5jzZFw3GQ6Oc3MqAfNNOdWP+BwVZY+d9sXX2KdvZG1LqLnUgLINmKmEqOGr
RmdMjiGweyLU2yhal+mwhB7FuBxoxGUlYnfII7R83izZI8mYYmVI/3I5n8iQq1I8
8HCwq8FTaq2zTcYlK1GdwK/pRN7/VqtEhutIbosxZXoGJuEGj8iMCko3w5frEhQD
vZgKfhZvF69gbgkemOJUJ9ctXIFe9gw0TRq0dDOXsn/lYhIHcJKI7CxYM3MBoZ7G
9tQaz0LzoDdKp0viBRKPR4Qr5QEz/ozV6JV+q3LipL7hNtwtp156psBihc61ZGi/
soXZeCdXtRYifVHSaEeroce53EBSxUDZ+tdN1RgH2yTn+wzSFalPzFuwZVSqkktE
j01/VHrzDhTu8Ur9yMcaXqK6IJO8cC3uQlWcXN5oHyBU9lfoFpJWlYJoMZ7QfBt1
Nva3BB3miWBBj7qyHvhbZ+4hMeak+SvFIfNQ4nJpV35ZsTAueKdHJ/t3rL5ihk/S
BlToQdwfhIyUH3eIbSxOv96DZ2Z+X3clWiG0QyXErTXzsx4SkkXxvGdnPFUzEw0a
Ei2HMhOODqFmrhO2Ha/k/BWJwCpTXXJTiwpAlbUw8N6nBThhv3+CsB/m7Wkm6iH3
evtrfIxZZ+tOlgORm7+Y8OuA83fUod18eA98KoS05j0P3iCx/ZKpY/dEsYvUW7FE
7jwgkD37xwDnJSuimkQSQbiNdr/66FUZUpFrUJ9a0vUSRq0MZNRpRGAxwIk83PKE
XO6a39m5dtZ2O3QqdTBqkrFvsJ3ue2WcaBGrIof1natnbUZzrXdE2kf65SlZ1IfZ
aVIQv+OyKzUmKfEFGVT0YZvf+zQ+GIVnPVGQykRiQqcjdW+f4Rd/U4XJbH3RCofw
QXGp3eDaJxsN+skpAAVsc1kaYrczyVFTdO0dq0Q79uchydu8FG9BXHePk6pygOWF
bUkrXO6AHgQlmAbYbbotYAgVi+pezYDkFnWgDzxTTvCaUF8VledbZouO8yrOt5Wz
KGaO8QMtsA0Atj98eFy/wvjTCZG8v0L8YPR2nnF5tXkTIRn+MK6pdlTB3DgIqCWY
7rhc4tH/GzM+gPZEYhJZJt2dQYVFelLiit4DLG1AeQfctionRv6glWj+cARQaajz
1uImHtsGoSYubbFG2CoxmJ+3Q/0NcLuF3umOTOXRl85ZKgihg8ns1PUCxQRRHtBt
fdB89T06jOb5ILjaQ8xbpMJjBfPB2pyRbPOyhLb8hjg5ofB6tI0LDV3dz/R0Aab2
VAMPoBJqnHxhLsYCf08im2n70xOgfOPoMbUav85hxXNMSO8q3DBF2EK4p+y4UlA0
XbpsHo1cu4G6Xk9FGr7H4t8Q/qHOkRYRXKgBjv/dZybz2ldKSnsCcvFsGAwOfxvD
ddil5KMU/WlENvmrKu76Pn5AdJdRSkLZWGuoMZ8VgCyb38KXp/dyufD6/0l8SWVy
WVXi30U/nfhbeS2TIvW7/hMZ9TGg02FJTxf7zWe8N4HciMkGMFvsTzFso6KdGTKl
ORMX38OvfHARF4cQmzCehEidAHRmbXO/wnev5BIGVzmA6VQBiP2U4UGtuD7HYjNm
NgldiMxP5P3Qux2vWUP5NR0abUIYvJuI5WrwPBonN2+d/HlqqST4SrMdAAMYtVHT
mvyaL6jhlJ09N5fCi1H8VgXDjc59/siWPBVoWlBJfVUkSkUSbQWByETY5tIwE26v
J55WRjP2akITVD50pxPrQCyOvM2VQ3zrMjh3/k8q4rtr9z2KWf8a4XAJn5+Iyeb2
ph0e96xgeRVaDWB6RtBYXjk19xhr5FlXWR+i8sYp6hK2swYrNAUalKuDoJhDAKHt
zDUyCjaykZyks/tHzEg1xbvgY7Kp4Kt/Dw6qt33aGxx6TlakeQLMKUZhAxFIpsFp
HeJ/rfidhhp3nvXBiBqvK6SgIy6g/ZZKGM1o+JudMiNYa0CZ+wdqa/7J88PnBMQi
xEir9P5cAzCGUm3ZkB20TLTojICdo5Pob6KxHhE4koDjaEPKU9GLCrHEKxFKfG/m
rKx90alhmxHhcOzYtjhZh0iLz63mFxdC6H+JLq8/cbB0xZ5rzK3KUvhw/H37PJ1v
K1fEH5Y3cH2UJY0ZmlC2VFxQ+I/j0yI5vo4L0ovhcl4WaFKhU+EFLXsG3I1ROV5D
rjOKpf8EaLFZdmVsoM8l5s3g2Hb1YM22nDqhwR8M6u+RP3sAVvKkrZjz2Ecufvi4
8LN1ZjvIGMQs0Qyg046iwQA1cT2lPvbgqJNKie5eFdJbIC5xSBAMdEIQJGwBA+up
9Gflh9m92do9j1n0GsRSTo1lWPj3+mzrEuc8zmM7ja6U856pvUamh8vyAvEspvLj
O1oq1lxGkTrkVGPDcxnYSUHsvCN94T2HQrsH1ExsfB7FHPQuZh2GYHahCYSDFfur
XajHG4mB2B3LxWINRnfQy8Ysndvhh4vuiWE8lTiZBwR5f0wssL5UROM/ZzPV1yVs
r/9N16JaLOz0wTfnEjNkrhrylchcZOp5gl6KXXt6AGeVRwYRKiMVvLkSDtXV59Jz
mVyNydVaxA87VusCSicGHXeOgIs1p6H3t3tsAFp+eYMaK5zqRgljqQ/HX5kYmZu6
my8xOvB0XbeHq18MuPhWRo79Y95TrJVxHLARSJsxLEs0HF2q0RePdm2qJHHwj58W
PokGJlsMQTPO+f6y6YMU9q9qjVkRSIMgfLFrgMxe/7DYcTS56YeHa3vjwaeyhT4W
ZBgp3j/m9xIjYdo3BeVl//hwHeEiTC2IPA0lYRpTVw68uwMFLNKwjdNXHbU5CeSE
v6UlOEv7bBubR5SbAWuRtiTCvpAgIMwFuSd6BcirE1wpTjf4REvSIJ8lp2L+XCWs
IyslhzBUNfHk/1v8/JNcJ9QqCQC1YwtSoBga7LfchBOEAbjerLVhvmfoecd6Wjkk
xS8UOJ6KKfGirNyVbMFKaH5wxnJyxg/IDFXjBfct65rTFxyps+Phy4+uGS/3Wjh3
7Fiotj5zEHGgTtI/c0d77aN8jO0nQG6n2H7dmP5QI1kqxghCbeWqTBjEcGMD671e
aTpVKIeom/vx8AWnJ+5GBkIgHvXM8dWS0cMfc2Nt8DXdE3W8uSBmj10vhhIlsg+y
v/GvWvDXvZpZR0p0GlfhER+oAVasD/sJYGtye4uLTe/7I2KB9oN0Omoc3AI6po+h
TPT726nuvLYFbhUFG8eWP7bCayHc7uIx9wR9mdRr+HLFVEpP6mk75bp5vzoUuuLe
AMCbn4C7xFnxwxnELspjSVx2/FsLa2+diZWWJY6YXIMzZxl/1Ov1UyZacFfe/055
NZMyHFEhpBSMu1Q1OrzgvGGTpsg6L26gwcgyKyjaxc9Z4wNFPV3IDmDZzPZmV+dr
uVsabCMW7y/pf4MOzrI26jf2/Xi6/eDHG19VKBXCxRCrp/iIxszOMcau0kSZSK/5
PwwJS/FrczGKCqt3eASPJ54StrYrEtkvxTTi9iL8SEPRUngddKT2XmeiFbKnU3s7
ioxIO34QxeG59siJpMJPF0JG5Q/qWRcSN45ca5PM6B05zAtK186/0bUWDHH0Y6zp
YDd//6BpK9JpUrMuMQDibIS4PKFO+ODL0X5KZlyW+mdEIHLqlPVjlc/zrUn4nTGS
s95425LaVcNFfnVFtxwkNyorKOKRzHRUvfB95ADXIdz8Eslyu823YDv6/FuMSltj
G5HLnCtKLGWIpV8hp1E1kZ86enlJJA2pN8h3ffC24qBH/ewD/cjaTrDTriGSxAsV
psziPqtTD75731Fcr96UL9OF0GIbz1jxfdECAX7bDfa+74hDmA1FreWQdAn6eFgV
gk4MxhxucGqomdz3i9FJTqfal0jGbcXgoGZav4kfSsmh8Rms82wCCApyHOo7SDSs
YHEM9T1HxP0MbHS9KNIVLHRWe0XWeUkMU7NrpehXin5E3IDXZeaPC8H7EBaBC9XV
K8pzlyEHVBCcvqHI7K/ZtzWZk7l7peoQdxG4AagYdFh5dUCe2lbhjpMlS9Pkocmf
ImksjYb3H5uA5qv5WOaI7TTrJ77//25vAz80CziqZWdepy8hOPX3X+YZMLuB2Z8F
1HwE0D4FbYbzKLL+GkeYH3f2qBruPs/r8mjReKTX2UPZvZzF02A1MQXZE+Owv6tY
7wqFKUqlBxFyzP61p9YHiaNw28FGomN4HRsFeYqdSq7hGTtqHolzu+YHjjYRLZqp
7jz6MSKfAdYopd81igUvEFTOlXqeeLmnTKp0p3zW15nmMR2lKsCgJSmgLadcIbZx
iE/5nlm6KOzDbZCNKYZwX+IRDbxaoYllL5A3RXhC6O45gE7/ZpvgTJ3CVE79ZAsc
Ogry/6rDbipm/4+fLJ9+i6oei2vY+3J/1FPD3GpmHIPuA9En63/q6noqZx8PHbBi
mh6KNIodGf0tq6Z6iMEVPi3xuVCNb2/GdP9eWI6fDRG4uurUwvhddLeyE3UBvSva
pFrEkye9Q4JNQ3+PU+oRYaali3sI8+VyZPmkifa/KKQaaaCugc2mPkvaUHnIWJOE
ZyrqbUosL0qWOW+R4zoWb6flfnQBcWZUU/y0dVlDTt4eJCHY67w+wS7Gen7K+ZRS
RrRu4w+htOi/pe9p8BMfYhooAVN8cP4ROAWlvIm0QnVjr7dMHXZGIsVMfd0WWRY+
Tn1JCiiuR9hbDKKXJeXbHYhSSk03BXA7Whc7gMzbwiOBK+i0nFBr8wFiI+iQbTO2
nQ4irrX7nAPfrmrZuZRRGE4hieezTyl1eh8AwG2qS0zY6kK/iXyltA0TQGAyLUCC
75B+7WgE/SkLvDTryJ7Rnjv+ZDRRZZ+O6REnRO9HFfmTnxbN2rbq4mU7vwALVbIp
96uXE3W7/3zwP9jyYwOkNoDgxJ2pJ5rdoG6ZtR2PKG0fMxWLZaeDsBsh9m2w4Olo
Svxjd7lQEKPaJhfAiA3gYiCDFHeGi22Xfzdg/HzK2PBJKrYMqeyuBb0eZJQ9Ro34
NBOMZvINx0lSOC0iMx94FZ6FSnZRaPoteK2S4XE5TEcUjG07KMI3RS1NSR+i15WW
bcV01oTY5MkNnp4e6SAO6yWWDBnkkK8RzbFzB8PWZ6XocPIIJyq2mos8BeiFRE6Y
vSGCr9jxar4FIP7Iby3YBppOBw8Oyc4UcFtSRlZKi1BZIa58DO44T7CSqYbPNms2
25JZix3O3YVrCIk56VrvE/4PYrcCQKgWYup92ZUh1LMB1c/2FbK4o6ESIQ00+VYp
HNi8JK3/4MTlp7i99aCqYKz3x8dfMPSFz7tuQkO9Uwvj4RLkrxd/SKkMJOpN6sM2
wC/MBeFrLcEHvmWIej9BQIXxheGPQRvrYF7JVZsLyD+gLOrRjP0vcgQ9wcZsnig1
cG/fYr8UUMyoMh3crFYwqNXMNVcK9LIeIob6fIWQOHnLJ6orJPgDexnk1tfoaUDC
yqA9pVLZ29b+cDsQ78eEkwDJKeTWulOQuysdctvFhoLa8ORp6uGechHt0orxiuyc
BzvLcbr9SbuFjI5Vxfj+8kLImuuDFY3GFpQxEn1xbrYZCZLyFiqxxifBZQOohupi
SGQTfT8m+FdIt5GlGIsNjqtHm8aBuklHKpBgRdrJjmy5r85AnJC4VykY3S+yZ/qD
sk+qW5vfeDYSj4oN7xivwgepNUVul0zlWYcK0do8hTzgp+v8TYhRFCfM3xxpKVqK
crv0HPNrAMCarrsCRFNxzmvLU5SdjP3RQ/nYniJIb0dx+1y6QsOCovy2i1G6qbCk
XH7vKcTHuZ17ssca/45ml+VT7cJdK2g11JLa4+20DoW6yW7ENiZcz0Xgkff+dDLB
po1TmpJXubPvnkQ3CcUQkCpSh5ceEz5bwmvUUapQlGikQlH0B2MZfACWZ5OHl0Qi
kcGUGHFOgNrFPYjn6os2ZyokfameUXitdVhsR80w4+cWQ1+OoDe6OQODhbLkHyP2
iUs8vNe6xDZMXLAs1e2qprQ9LuE7K+1X0glT5y163xZyguTy9hW3aQcFaKJ2NlHa
Et++hXLeGS55LJBGmEhMNOD75Vh58dpnWpTjHjrfJlAdpnjX2TzNIU72TOay3hA0
M1JTNsMAxAB3jclztcmZyRW9hSyj9kHertmHD0eWpdhkFErB0T7YAsrsr6RA9kSz
kH4l+edm8nDMDYJqN/uvRKjk+jMAVwjLOLBJ70ayf6hdLp6+17BL3+ZZob1K9Mj3
erKO3cebv/GTIy8BZukANnmAWzqjNrLHEyWq3H/Tiu3uaaPucBGClt51kYgJ/0gL
EUeEkj6CcTTpPHWbo51iMJO6m3ezhXGS2XypP5ToY+j/Gtt5VkmHs6ZGWF9djbaQ
rlZZLUFSTKZQ7tikylx5y8+5J/EHZ6eVZI+u2F7yyCiRbH2YEyV52cPOjRqXl4C/
k7orlYR5Qf8/ivYiiV2ixc4FdpMbaNYgWiAT/ndse23exbwXtuHzHvq59/Mw73+t
tHZyxVkHcWW87R5Nvzudi9IAv+oYWK/MR5PM8fJ4h9tTooy1Eq+P8vZBCGywKNIs
I1moO5HvbvuUvReRJX7PqJ/hGWg7jgqOuLYo3fzSHWMRvwcGrqG/obdAxu73qkht
O61mDP2CxnAGQlk/HPaiD/VzNxvRLT/qMWIf34RiAiMOod0oV0fnqz+PkpUH0w0s
F9r1ImYtclYbJd5rBOCQoU3MhoodBpOyPzRz3I5UrD1ThxTb10zlm0VAl4JrFuxA
aay06CsNJVqOfee9dREJn89HOEknySKyL9V6Yn9hanv0p8uMMkYCfDWCyz13mn+O
7CHy2JwDM2sV/xIK8yuPfglztRO+8FSpeSp/bCQtNTmk5A8LWTqx5k2h4nQODeNk
hFUgOHP6qoeEdKyGu8E2t6vZY/rs/noH7U49QmjsRrjJRWBNsV5OCtwnIrrTZKIq
YiIORRWtcVogS99y+T94/UR/NJp2ehtbPq4gH9dfXygEJt9ioUc0OJky81opLKHK
KgPtrM/V00+8U9GgnjH/cqjGVvfUSWlp8CkHSFZFosmNChODrOe6jglgLjYlXi74
HNky9o9GfWKv86Oo5rxaK44XylwVcP1NKivi2HRbzWyWLNYwIWRO63L99XckY8+e
OTEMpUKKy2n5tI0nMPU7kLkhcR/lzZmkNJsHz39dnkWUpfMWmu1iRY3Verx/pJK9
IEKsaWr6aAJVMp8dGVlU9zQ/5s9t8bt8I8jsne17SLGssURr9vX+zW3I+u4uEtWx
1RIoDYUvlIEiZaTih9pKtZ88ki+BG7SsnZW9Un5ImV+eoXdC7D3kgbWRfIDixJuE
M8/faB9vzYiU3LKtLhV0MzsZPwz1ZIr4g2AK60xOxOKLlsBUzCvtBa7ys7KF9nbB
Zew/TKyxueANNMRba6b0lWToLq744cCwpiJcCvuNd+8ltGYqd1IAxzd/OoIjLZ7u
WbqzBfKFA6V1rpjxaLc5FM2SL681tY0m3HHACPJ3areU+ZfMsEaM6MYg4Vfdmw9K
vhn4HgeSUJpquO/7SLhhICBC0eupdBIQHackt9pgEIy1ZL/3KteK/g3705WEpMCz
ufkHo6IXeoHMuAs6CCtUGJDBUIZkmyAosv+an0bQmJ5n3GyqWZwheZgaWJfIfZ32
FehOaLhjhJ5S02rXNygTb2Ifm8gZy/b97LSDSKRV8Oiqinh00muRFl1OCDhyRwsW
9un7CaPy7U7SPgROe5WW3JLPIH2cl98MvtTNtTf6pLiIy16Hdlzq4myv+wR2fNyE
8QrGAYb34ZtUsPBohXxLnAIAWzN5yfzESJf+4MZ04gBV7/M9Z3WId40lgwgofCOt
yXvem4gXrhOZAHBDDEMH+dFlzRTkrHjzbB+kCz8yqkEZp6j3VtREX9HDJQAVxwd6
2osExoLE+qWKFLudeEGBs2b72hO9w+OTPr4J9BSJ3tpTcdSS2K/nP4aYCOSV9mJ1
mJ/1rFdxmSsAWeh3n5v9iy/QCebqWnCsidMT6jw88AErV3yoaipvGrqVCP5WAAoD
ieuNMDNvnV5oVaJpEQHOwYi8x1ZWA54Fr1r9sFB7eXDvY51f8Flvdn2rjh/blyPz
4YSDcLpXETzkXKORScULy1SMl52dlhaaB5GLqTZYDRvU6hcS5TTZSVlcIB9N5tFU
tCNDEpn8LKW5875mCcPCPK9wr86qSWb6ONy7gcC8aNsJvZmjbck0DcdKYYj21vTC
QjNkEzhrTtBlmi/My3p2evIK4DJkQmIKtK9/revs9pLI2Cbq9SowRQu3tTCCspaV
vPyRF7btbEL9UKa6tryYU6IPjEQgfsHGTG0K41D+tMiVSrb2Q7+5pjK/IxZCOgWo
55xNg9CcC99V6Jek0zeaP9bXuui6Bk+bkjJkZcqGexV2lU49bIkGZc2hAvoK6mix
h9JNH48nf+88JYruLzmayK/kePJEQZURLX6ejlPzkowvBewRvgpndSDV47ULhhGG
W4czHAyvqSe7preBlbIP35zz/hVnngzLzH8ImC1YyE/LbZI2haoL7oozKeCgQ1Bl
Onkuoebxz+0vEDxa5dZj9mmX2U+NJmFMmHdvrQmg1x11UQncf2fm25mvx8TIrnxO
s1b3eUXzYIQy/7VFGGOF2kbw6mJr11DcvuEm8D1DOn4QxhQN+DGvVu/rcjP3Ycc/
LBLa2l8U8z1qKgu42lX63aNTYNLJbI4tiXigzt+4eOeK7brNDZZWGWu7xB2lxdNX
8SY+ACXJ8sXLDQYvXraa+hyQ/R/K8r0F4xs72AXB5p1iLKNwCR34xeZEBIclEve9
2qHYoZi2CleWY2xTt9cRA5oRxYbvhFOz9P8hzx22Ma46uJGBqBbbB55TkpTYGWy9
c7bj9haVwDOU4k7NGvBQgZE5VAlugrJvXh/DozExugUrhQe1qj2ni+SKWV2ROEPh
Y8tkwmMrMMQvynPHkVumkPWoMlavOi7yV1mibqXzeAbU5snEM+gfZV5mTS/ueIVK
SaJTC7Z2DFG3OjDTSgHiAZ11IlCVqrNL/i6ZUz1vs9iQJkj8QlkkoD4tmsNMAb3V
UHAMfqzko41AhnweVx/n6XKkKQVXb+zqGjeIq1GHuvTtmmQHVHf8OdzInWvSQ24L
syJvomrqy5N5gA1beISBlxuiy/XZ0AGJ6synqDY4i+uOYYkYdD+QzHTCxFJxXIKK
2gcqAeDW6wLsWIwILOwjRb8rHkQyck4hN4MJ5c57xhA+59p+qezFMZjZbE7lV06D
i77U5ibBOJ1b5u6P9P0VpFYheLqbaQrC1FF1O+WTgCKuOXUjJcYHHdVNm/LvZ9L9
jk5CCCqy9XFq4cGNHkDL9Ye1mhFGRg5e19Y0Wz4LXVLQucgd6yowkAN/eiwRyITD
cI5ygGXttVGxAoRTrUJimNQG94lhzvzIlJbODNnkOT16yaVp97TukZZAP7ObCMck
S3HC9XGkEv7IIAttJmg2RXjqHnA+YKG/eCzHGQDVVJXfgm992ku4txbZLfRh4K1b
uERS731vhRJAoLkcWDI91FwgWxfSxDUbL7yq84OU4nuvbJtqNOrZonwig/08FKJO
i/UsKZereTPNLbZ5vUZ/S/C6q3wLIzqKjSly+LzYwomE8lPzbgV10jOmSDHdZvfw
3PO0fzwRQLuli5T7of8KvYDWMhX/aN55xgNB5D3zAREPJcAO/3JNnCaeP/Vqw+wc
cvRhWEQLEcyMLX6WCm8C19NMsQ/vFhSum7i3lIYWYN8tlwKIRzqvshLzfXBazg9a
dRfK/wqQDxK8PACi+u2V2CgmtncGzY0VHKrXJf4tViUAmNYe4PbYHZPO27Tb4A9A
40Yh6VQffe5dd5KPR+vtdg3bAN1DGgj1sTIsdjp0SJ/bx7PGj/C/4UIMZsD9YEZY
04+8hGTRBg7IhHIVXb1RtsSegCDaOBr7CW4cTeiqfLzNxr7UvBGsx7xIibwENB2T
8O+Mynm4ZzB0GuWN1f0CDfxzCcUTtC4EGDlF8ktLpVuAMWHkKVkSL/tzDGfItXoo
ZrrZCB2p9TQC6b81yu+vgVrj3skXGn5mPgSlX/mkKzKlUDO/YJDRAStRSL43eCN7
K4Du4PF5MQ9Q3OQ7uh51QBeT5pTaMxnE4KrtAbX0U71+J2IV+4YgU3tP27Brp12S
UWyb1usKOCTMv4T5AcT9jtNUej+0xFjt1AFrvlcnMwS/S+nLKw759eXKTp8sz7BT
2X9vQn+G7fL10+ACVr0XTX+m1i955viGt7pW0NpwEYxTDALEYBQzAlRAqt9Or4Sw
HCVuz6jgZGPuOjlFpR+pH0H7I1P83ZjZfiM/LSFkcp9nbECPeb738IoLsfZZ5qIQ
HMW4YqQlAfPBM7y+GvH1TmTYSAykN79uzXVHvKIuGrXUrShJjBePyH+bzlRQM0xe
IVjnNjYdY3AesQEUEenQYnjZRoAFI6ASBuBXvbdIlJNWvVKUOmryOhJSDx1R6OBP
lNoJWGDGpm324Q3nN9JdB60/oWnJQb4us5wOKOm/j2M4+vwzmZZsIvV9t+KdL8bX
U7dK3kWg2kgHt4WhfTAzbzsUfW6bh7no+w+pwUZeSaaiDxWURQCHaisIcUiIv2N7
wbqLNZIVlSOi7iBquqizxB+GwhNFheBzUba9m9YHLQ5tgCxVTS2zOTy4Jskh905c
741vAa9II2XT/wczhDEpc+8a+6G/dEkNV7VOAb4CHT2fnV85hKNQ3P1mizJ5Y2+d
IXo8c09KdgNeQSkTG/C95j6rdujxBbRxk8XX0uBg5L6RB71dtQLcKfGZRXi8zBQo
407dEiWv9lx6XAbMX8p+ic804RTqxoOKNYZAUCRT7Nia6OkbusRTUfUDgn0MYbYN
rFrjBrtIAQCxtRuO0C6vbkU2KD4A6kwW1TO/hDZjWtWGT78FgxuUw6N10eJCSsFW
Ns869HZMhmEFNWmpk3PFqsCFYqHPyaiFzeRwlYpNcPWcPW1eZ98GGqleL1xXxbpL
vphIDdWbA/aIH2hrYPo+bE6N5D2iN81AewGfLjObEk8Xa2CPYmtp3QMtmc1tN3pC
SaMaaMD59NuirLGlskwdXKBtwcTudKoqDNoJF4IDPSOJIoazqQjmTh+dXUfgm3iE
xWppgz0CG9qJPFBXsBEuwu0bCPuF6TaipRnqZ8kk3UXyqeAL3IuDlVUe8VTiifOe
wgflw7mk/mI6sNiUoBeNqwdWbLVAYuXND/pp7lbWrRXgkd2nMuGVmeAeB5CKAETY
SMeYQeAbfoGaNbI9D3y3+Fc3+Vp9RUwiITeqinOTl2u+vWlI8ds7io9zwlTLwO6T
Mf8sw3PVhhP/Tb1219DQdJoeTEvRFxngGpoDbjFjNqoMnCmlksyRd41/0vUj6yzu
ay2oOKHDQJRKkURn+Hvb8vbtxuEd3DIClCn8SWIGy+LP8X2syOsoTfq4T56kt0jq
jKnh/9updgLQDCGPxpTKd2lizYFK1mAWdiv6AxGY9eGmFmDIHN75Li92hu/ads5t
vQ23iBKw4He2LNeDnG5ekQHvkw/1sxHwt0+kn0YSWgEp8lElGM38czkdBxAlQWSP
JhQ0+cvLpG8PcWczlc8eZcPquG7hYXl3rNoCyE6DfM8akicpAQSh4TYLlyXh7ok6
+TnkHnhDMDtKhfR1aRh4AHrniyY253+lQC1oe8o4ZmstLeFyyVNa0cVpFrpjwqD1
tmcSz9cp8hDxI/xAB4ZmoR2gJ/DCbeWQAnutZOE91QkXvv7Au22PSUHWI1faIOiA
gZ3B+KIhi9EWbQlSf0WjmwJC97CEh4QYmJK0q/Tb0AMzWpelxdaptbXVV/og0ZWO
mdYFP/FIS2zi7l2+r5RKJindbTsNOd4DiNbfc9OPWsbtAQ6AN7fci7NcO3pPisBm
df6qt7aIIdOrWTTAwsTqCvtBfRqdiyrFzpOC8TQmLssmUzgkiJ2k6sDzfl+5W3GZ
y103iWXVhzHuIOV1KU+JEmUGam9aoTXuXwI9IVYCzgxwSKUNkoUbTJi4YJ4oBKHs
zqk5OyOVyinu762cDrfDkWK4hyom5NCBpZXCUs8MpOtVVJH8Nucjlg6PDrBJE8nr
91+A9RfIkqKm32RLSh4nkgRz8sfO7ehAcGHHgJYztJASLZI+etL8/HEmor+VXGee
DIqtam1wpbSKR044dTy74WC4v9b1D1cYCvrvvk1aciooQpWYqxm6XSuS4Wp0blJI
lxn2jNkKxuh8RmFEdEYHNNpUmjXJfrWpdeP3zvZDP4+qprifFsrjYYLwNBWofec6
fP2HOfGDz84fo/uDUDX7AurGWFOMsnk/yUD2Yurl4LGaPR1kdsj5c08ue3eOJ3br
kIqrMdNX+21vG+JLy4iYZwCTx2w6MI5xAy1XEl/C3Hy9t+C7nPf1QJR+EiPfDqwb
bHX3M40qBLp8MjhJAhjWZ6RBf86dLsIJ9laQzchUg/Sna0xC/ndkyajXEtGyuyZm
2Ik8WdrhPUEPk24kyldw5sp9UQBsTm4SPRWhOlrQPqBG5LzKMyZEt0P7oNqVMIcK
fWTKXAKPJXvIN+fQ2BRKrnpBvNH8d/AmI85d02hVNSepzbPVImCZlMnM2gzjoO/L
WFvZGGTu/jr5n3tu+ZmxC/FtPGRBeD2uwtdYTEKEBTp/PBszV70j297pRFSgVJ4w
G2tVtDdYif8u7UUH8SR6t0Ty2da6UxTCME1WDLPOrcicdvbqlHuR+vPubfXW9Tgd
0FBBDKToWJ9vnZGvceDwNzSVJ3R02YJrHhhVCH3nisRujl65urv2EIZUULetOPGE
E8vhdUCKRw/iumJpTrlXQyOstpPb6CFpaXxINed5uIvmkEWxWjK/M/PE2ItGDRia
MC7uOIa65+5D2XgWUAC1+z0Xa4BvSgBAZWKRuBxfhXCwjUTDDdVnKceMW1mRsDcB
7R/M25OpfuOH+d+aqimv6hp/hSv8AhIMdiGX5fK9uXLu4cfaTRKSayRX81rLlxvU
Rd0802BwRCUvrojf2sz5hD4jZOWLzP6ld61Dw0L3gpx9LRAYzcpwCKSrqb4lHWTL
055AwjpCHXUfnwFzS6b0bPnhPGRE+RR/voUgXiXidPRiAqY/1fwpJyqMeqDZ16eR
wQ7wtueauZhDKzlGwLJe4OXEH0F19rMaILbIYpuNHjkz1VSAB5YV+Ji1J/HVHoED
FDcqI6k1guUS4YiomC+7FUM8h0p2A8MOXylpQNEahT5SnGymAvSb2oJ6eri2ycLs
xioFDuQhrn9wHVQ9REinxxPGCeJCrECVRMeHLdt4k0IEJTZ0+/70UV/GGht5xts/
AXbSFULE+QLKfgeFWGm99BIINJFRM4/3AyCbA9HNIh2yVV5frW/wC7oYIF386B+7
KppPvofg8S+Hi9ikfou9Etwttth23kk2xtCvXnaujkntmJYua9CCQ3+dF+NSh8DC
E8OrCPwbtqKhpDtMQq8dcdMTZjbryLhI9HVDhGYRUpMACXZsVGjYmU0Sk0cUvMvL
H+KSwjnCOZozKgSU3vdwfmVoNUHtj7W6hf7UdSk0uAdS3ePNxEy6oTx1ju4KMtdR
keyD+x+FBuWGQFw00GwkzICbfmw4RRZwTcNomLElzVkxK0ZH12uDlSq8h/7UTRl3
E9b9DYT0E5hu87/UQJfaMGdPJ1jS6dLgAd7+JMF7/PDsMaV73LGCSKnhpyQlldRW
9IhScb752j2vD/CMm13ld9VhQugp7B1uIUGvSyYNX61ZeSBgXuYUVAD5pJjX/OX1
3jxcjBIiUDIp4QgrHDlPpLnJPJ5EzjObbroxT2J6rOMVeNseH7Aosr3UBpE8KeiW
rf23+Me+ugnbQDUFPnnbG95UTHLfG8OfQPcVjlfC8nlwbz63EP+tS4hKR+3cEb0x
g7ru9nBBe0gtpKNbwrlTbGta5MVVQ2FR2CEPT0kVbGYEtRmYeWywG/MqZ+L962P7
AHnAp8zhHTeaGSYgdaF2XvqBd+foK/Lg/B19IK9BEVYRIL3lQn4WWFso2OcCcASQ
+w26qVJTjwWfedCs3m+/WWaczqsO0cAA76c+/LFIgzVha8BYTbtahSAPbHe3iOpm
lSD0cql67Fx4QDI+S4Flouuk0uwe+VCGROL05R8fJFV8uSrD229IXHtOKbLpmFJk
PRNRQGemX1OLyUGfrapF33FdhMk80QwcHdvIQJCPgdNQzjFILOl6xLaVTMOMtL4X
6y0EiuBO4DQeors9Nldz9d6gMyKYCQuWvae2MNaX8Y1dw/9lvWkn6u0uYpZJsnkj
+1BCT1SMHd4DD1YPkdt93+8tILSOivT1tWm71mOOkMbZB9qtJ6qE9A3YfAX9feRO
j+MjbX2LpvM9i2LDhwqZBzLxk6uG11iofX8sp6seoVYpUsx4APupOsG2qXTVBtz3
2MZ58vBE81u5fJuEZ9Cx7oc9SFo+691B4+AFNC/mvxe4Rl7nrsop0bOxYlX1vFua
W2E/ME2iAP4uMTi2nH7lIIwrJ9O4I9xv/pMS4x5yAdoQGq/Y/YGL3u8XRi9/IMmJ
42UrtfAYbGYop2vsFSBrHrkjxcP6EndD7c8gNvl818QXpWjKGuRynJH5gKmGP4eV
EUKNw3aPqt6O0NHf0P6IiW96GNjpJS8LHTtm93VomZkBQxJAD7HBvwg+lit3bZcs
dt/8NFpIAPmfrXtVuLh2iv6XQ5fciBdSNZrrsGXEW+FwuZNsZ8SegxSMkltURF+t
jhtCtkHHdkrK0mbAbDVhjj1T6+yj0B6SCc4QRn9wfAiejbDtKOGyn/FVi43dmI2y
ko1ZWdD5OkEYQIA83CLvINrCZKyd9IzHANma3LLURs+h+tRlC8uvQrg2iqQEvP5c
fzCXCIAE2xbYJytrn7uopv59BSihjtCvt+vn0B8LnxNTy/Thc0v8uLHDd5Uhe2jk
W/LmksbeBiLTKoVyRzE0zUl4qLLCRIxpMy3uaXe39BlaWd4rEk+OmSM1VDmPXwws
gqO0QLLnZ9mNTU25EMR+AjxAbOHBBpC6foB9aui+DtuMxjxikqkedRke/Top/cVH
jBA1T7aQmuAkSSdRUQ9x9sCL9g4bR+EFLd5YdjsQI2iWmAVZbnnRs6Nvd5qgu6xc
nNsxBxZ+XuIwfWQe1nustS37vtAW53cSAWs2YnjVZ1c3G9a+BRSikhC7XSZ/lneY
aVcwGMsJC4j0g091GwjDDE8wuc5Nu4sCQy7jGOSs0ozJG2F7cZAfzKRULg56KG6+
uoPp8QFTpHa1oQBUkrYWxzqN/Kp5LroQPMiUL/KK88eOHiDI+vMzNXOGDorONnhX
JdVz4hs3th0ao9icQFM7bQ/ohIxz8YOahNJU/skKdLwg4Qm7MHamOAZzFkDYtaDF
neuR/ksCKOdfIcrQ0FZNP64sLUyeooqPsFAkwSTBfG3XfaN1oH9ZzTuXmKjbeYTp
tWqcA0A0NNiHdRnZDg2evt+AdBX4T6yZbfk9k2wkTMSY0ERW0f4wuWM3EXZcjN5L
T7WaoWU6c+JBGU2byp/A5EGy0R7m+JdajZ5pOmVsNc/KPosV5eRgydXh7zz7ko+A
3dwnccAHOJiCSk1G2Hn2HrT09waK4i0GB90HRrPpZ0/iZNLMTNmUzmDfUp4VSZCP
h7NY6FnHCYSy7lu7XB/Ag4acQC/wllIMfnrbxqVKKOH7N1aTNgC/ksGCrt5A2fDt
xr/jSatP6W4tYC0PRImE4gVwKGVC9zPN5ImSWRA0LLTV/buXRXjhxfk0TJXDb8h/
uxvMD7ZjRAOAX9bXvLg6Rd85FUCSCyT/F6Q3O5dXaTwJie9PjFNvlu5RMUPaDHdG
71YuYgoF6vRn/l0pzCKR1HcUzkoCxHqitcvjtmj+k0PzLX4zhwPLtk0RJGInrzfl
2xmqFQ46JSbcDtis82pIvOPDZx8VFRKub1UZGbn8vffou8opwwAyu1/jtWcjTHl8
JxOVP2pWMtyvE4KhVjEZXxUAZ1ZgwKeKD8VukDQVswqdhEdBQA2RFRhp3i7lY8S2
E6sY8dxNBnsfDHJH+p47HTHShQEqJnZW17ttVocsPH11PElwdQdK6tEU5gp9k6CM
mH87ZRxoQJaG1GlOwxQbYbL270gDU8s4OjRZI9ue/S4tmnOo77ZeIgxks+VY2xqn
/D7lCoYCgpXdwO15P5y3B9c/dDzMicxtbOphq+vcGhmUS16UBNwXVrPsdlsK+nro
vaDC61/sAkL1qD5tYHLm2RLzT2ywe2LASZv74DGlDoR00O4kiFYccwAEO48PBZmL
7I0JZ/Xo6QxP5ADLq1YI7Krwj4TvtlwEfUhSiyCUNO0FJDX3ZfvXqIAGzOgZBpXq
2yifhEKZi78OQlmkDy1eC4dLOfuNWQ5j/Xgc3DLe3LrnLCGogQsyAzDNS+xsBJwa
NknwKuvJw4sVgK3aTYFYewkvRp+/IL8j8rwoMIGCJuV76u7fAdXLe8mwaUraYtBp
OFWtW0Hu8Cft62119M+JLCGDV6gwECeF4Iv2g4bGm8CwmYGd9S1Aru2IAdG5qwX1
fY2NX9KCj/FukQmxRHhucRANZ3T9uU3ZJ5Kr2OXUVYfzL0GUWZzP+98P/BI8EEKR
ZsM5MDrKhY/hpq3vcrUEbE055rdrG87zEGuncEU6CZhXJ5JPjfjdgpuJBjqJE32e
GdOu/VLy5+yRtjKGm1Bd5jpLs0FlZo0HL2RdLj7gR76m+V5Uteoz/GdWpilEXTXz
k9B1An04RSH7hCYnwM2RQ3e42OH7rIiyU8W7bTwWCp9Aocjw7KbOnrNKAB465kof
mBAfdoCsZEKBpD9B5gWHeUNNJYO+yMnCm6k007sJ02nN8UvoFmUeoHeBQg0tOE0s
Z1F7HJBhrVin58jiba0SVFxM+sNt0gB/W57luzi0OGGwJ7hEL6uIsIwl2GyFIknk
KQxpeyBR5nIfXWtO9GSKQK/e3wJjv3MoJ5DEAVoyRwxa5MWmHZSUJU3PjtOCfhUu
lbgeLBRrImvH2E4kaSk1GORb1k7XeZh0rI/DJVnZxYFF0EbNIbIpYtcr6nlNfaq3
qt91nWZJAIXzzuIZWIDFa87RU7EPGDnd0/rrcX2CfdDCWfB4PV440UTtxFJ/0L62
7y5lzVNSwWeI9NhU0My3iHT3Tcc+1XAmWnxx5nPMHimdC1ufh+6pnnmEgKrrE6Tf
2bRQ67CRcAav4efo5q9G3SuAv4N6lOOriBzrRzj9WW0s3Uvl8KgPYWTPFkgxtJqh
SPu2KN1UQ2Lv3HtgMMZs565ZpgsDtftsyKtsJgvIjV5bydOXfoLKtjeftijCGO8P
cN5DZKKPCPgj9we2vLX799vBuuj8oX0Wi+ta5IukdLYEV0FaIqpz01WfkD7Jo0WU
1j9iZXOc3tVoY+5+mW9NDcxMxGseDZw/giHMOLqQCfgtB84sQ5vboFYoJXE0fCZ/
XHqilWjO2V4LJeOtmL+ZN3mu8WhpeOiEqsx3kd0wX27e0J7FzRiUUKi1eGZvM09l
OGNO1s5LsxE650jXmbW9h585ZFljY8fXWo+J1WjH97WcEvCfTS0X+KnEJtXGRKpX
9NV2MK+mducUNc1HhPha2F725xdu3ULKqiQxDhltGyOBgz/U2Z61tQD/4agIw4Kt
yv9aM4MDNdj2UjCvsoRMgzRWobnn6QpB7hG5OC3sFTNQsN2dRowcpBpRvjosQNFf
7XU5M9pxxKV3TSajdVgLxWKmFg8qcZuhQJhODlKSrBWLzSu9OLUZ/1qPGXhj69IK
VSZrJD9VnkaMqlmFJHlgK1iVM8tLpJNlPZ+pD5/6nbQlEy/XLDhZiRxWVIiGDdWQ
TOrB/gPAPqjRtxLXIqhvwqchjXJzX7Px5+Vhsvv+jZbqBvoCx2Ppq3kRrNJzCtar
Hv36uQPENSvIXJroqMHkYxmNt/nkcAigHTLaoHk0xH+RkKfgvXks+ZTORA4/qf+r
2MVJ4Bwq8UZlLwQXd+9ykodU6V3mUeoqCQgc8Gs4kiwiowQTCKV4XlXU+s7MU/QT
M8+KUrRwlmHZvuIOaZjIDu/Xs0MVyMSiRht2oAjvH/DHLz1dlhwnHfu8+QaFhFa3
v5yh/UtDfIj2CrswRANMBUKTsi2N1EMarJd9qGM6F3SagcnlcRUhISdN8wG8MLQd
hM2V4Mgte2pM+MHOZFubOPkGE0CiNehz7NaApiD97aKkbTgVE0NMaFGPgp/0klRu
rhvKFF3Lk6N7jJNfBYW9pREm4Kev+WtTpjcNVA7p34VKNyFvIeay52U+IB/2QwHP
QBKScneAQamA44oG56sAkpfbwJDQnaszjy7WRtrhv7PkLamx331CPEJqbPtLWTm4
bzq3TP3y4CVYzt24MRMhUVWoBkas3Wzf+LGjPxX3qO/UGy4A7mXDifYbQ5GjAr6Q
TcwlN0xxecM5vE6ROZUNnL5caJmBuud+zDL5TPfWMba4Omrq/VGI2Qi39WsVUIDM
xnHbvWSHXs/WYRyGDCGI2dEUrAJtvk3L2Z0ME5M9zKAYFaYXA8hrpg6DibQZf5GW
DKF9s9S0rOrkXyW+q/orjsDRYtbTytqykcnrKHbtQXq0IXjuXmSaWu40uDko9oPf
+Z4Q5curggKnISB3wMs3vnvdt5jQdaL11siwMLwPg6DU5P0dEQKVnH0Rwl9uRVOo
rA3V9KU70iUPyNJVham33+pusioDyEJX/XZWWyM6gfio7djlx9aCI7UvSGw5muJS
tGibjQi8dVBGJlcoKwtO6TTL9Ya05ezwzOZlOCM5HwzeY1YJcp4yHZtRDdVvBY2v
d3LrVTR4WkE5OteAaloDjijvU6xeavn6EjZQ9NcLQAHbxSQREEPwbyOdqEtOSAd+
gqduJKtId7cYMDaM3pcOClWwKnf5zl49eT/PGQU30BQGB4IyeiVCQcHZ35UMx73v
Ys6c8yP5B6/urLUI63obbydfqYrQi9pw8sq6yqH7gJRj94eMIKzyx/kqFw7BdQTk
CRTsi9dxebzao8LfywnxHlr4LsSiCExqQIuoIogmn+dn1G7E88S2G83gvy+pe/sz
ansaoT54oJRlEIv7GgS32wfo2i4wDxVtI3t/+sd12PB3TmqKEu0DVglBjD1Ldtgr
O+lLfwtUlGM67wacjpDlVbLLRfxgh1ToQxa0ERyNzyQeeFFGgQxOBGjRL8x1YwVE
ohftc9RBXZxtCbwXEm5LVMxqBeAC66z02mJqWFRjv7GeKtbdTe7ff2+KStrXxRfA
iIANprN9DxHVKfOTFcNisWkCx5pxRmFQ0fERQ3WRqFUyObYbiRdV5PS3GZ6stxE6
Bt75e32VTv2cwoGktVIA7lWWiuiZ2jLsrX8cG4XK0S9060bCa34KqZRDa4+RkQeL
iwxJ+ZdzIYH8YGAp0pxzuC5C4Qu6ljzM0uYzZO9mZRUCcaknaM4RdD9c57nU1Dng
OZMUISmByrP5tueY15cmix4bSUX9GFla/kiVijNk0ILTeZcg+DsCSzTGZJRBXjat
+z37zCOODUwqUrHbWlOjMROHAeEUqt6q0SneDg35bE+bnX5b4/xU4OfHa6whRdCB
xgKS/JDrYlyao37835B8/+PdRTUmK9vXq45tlxtDoHNWWqBhFx5vLVyrhkDMOrbi
MN39zwjnyg72nrilcg395ioy3QYi5L+mDP0iVK20mHaKUwIBnUSBQyxNpANt3o6g
7CLzclw7BWdo4FbJkwh/hG5N8J/aDRZ0CtKknwshu2Ww26Om+RxLcAlRQxI3J5vt
iegd1qqtOcVHw+/HuJunbi0Mf1UXzdS9op6epVB3v4ABR+gflSMQXPcLoARJLvXa
J2NS+fw8X1N6UqQ2gEj3sc10qxxXWPfChWUU9xSxrdeD1hnItMwLmxApegzn1oZR
hz6iW4qGwDDTTkgCSmuKry+NKyzUqA0t4zRGMmn8nXaZiHDkSM8Y/NtB9tbh5ptb
b5iCPSqhTt/i54IZk/OJcwqtP3I6A5slIQqE4FYDG31/mGWKECsqhIoh5j7jJXo5
c/FZixmKdCs+CTO4GR19Vd9G1/QOSZEhIOOrPOSpXL/7hQTOH6xiLW4SFNXf54qp
1hme3Rvljkq/lbZtQSE5JpCzAAvZnigeFn3VU7LOIxB3QjVW8oStQttI16DAMpK8
7slOj+8c/Ubnp07upjdNdEMxvCx2SdETLh+b5Dttdq3mv8HTdTXsRpZb9Zhd184f
Eb8NjGbUMn4AC2anJf+SnVGItxfSSZVTCWaH5LAR24YNOPwMK5VtsOyolKRbpxZY
mt7twO59AblJIQ42i9Mq/9NjGl/LUl1eWePOJt9KFd6W8wjxT14XvyU4Ty3jZ9TZ
4zNpjPqxVgZFUPmK8VjhTJm79EEuVfnG8XHiToZV5+y6U+I8Mlzqz9t8u9CTsyCe
DAGJmkWz3ZQnydl5F+h4RPgbkDMA6Rcf1nLOiiqlk+nJpZMbxpeS7STL5ZJnwdak
KQryBbiatyrINAmRk3D8YhEPcN5iA1UPZZqZvEZJR6aGa6WMIF1FaihAaXJX+WDK
WmxZrJK6XiFq+e6lmBdj41hkQ/OjIykDoA826xFt6ph+9FVWjLDORl/snKQs4ihL
p9IOcTBcAfAIbWb/q6+hKS9+n1N+7eJvtZWYbtF1bUM5x59Hv6skF4xBj3lKQ3gE
8Jm9+052F/hNucuncVVy/GCVsiFHpvCzJgcOPzxF7pzxFclZwxxDODubeHAp47uZ
Ba5T6Qx9E653Ztl86HAvS0Py9tRJKUeAHGktmIPSmssf5z5bUZggkLEgAkfLv/++
/y4OTKJDp44mnzGjrQ+VXRBY/d0LlhPHeSr/WXvjdTuBW+u0Uq8ox6xXL+QDJggv
Y2+nuO7nDGDz9NJvJ9Y06oIb0E+RW/3nBV9v1MdEPdfGcpUgA97Fb3bz2wORmJWt
MGp4boNdOgLvnM4THK41/TO8wpLWe+OC5YVH6tXiSsp6eFMS28zsGcsS/Gs/JzL/
j30bqJlNIKvy8yqtZLdajZip+lgnj6biJ/bHddIcdYENRAQDDtnQ9AstvCqNoQVm
8uwd5mU9KR/oIKA82ezmodcFKPQFvli2NOetKkSxU2ZlFSrAMotmPiE7obCYwG1T
Dm8o56u1b9xaCJEv7YKND/iUMKHLlkdvLKzSPyZd/16ii+MMoLFNwlscAm6m+uFW
yQiJY7n8iIJKYHmp7suh8zbedoV/82NZ8IoFCFBmyhPg6Q+psrejrBsFf3sGRA2O
hwD+9/2KtTWbHmHu24/T3iwCHeerroe4Jz47KtuUe+tr81OnT8ewE5pUY6qH8UI5
GNTPEPlr4iN7aYv2zbBYHmyB1QlM0/IOjLo8eUjMEgKqc1/p3ovTU9YiK04jgZgJ
DLN9dQFDxVxrMsWV7KT8LJ90/kq4CwGyfHaqdQ2UVJQh71qo51VjRS2nnMlzOqar
+gXiAlE653ZP7RXVQaV+lkJPSrLugOX0F3oZAsq046Zh3CBtqjGnJYYjaBPa92S1
8N5OK+OLcu0Xvxlmfm+Fe07Lm9Pmva1AURw7myJrw/HigsoR0IemWX9+RqELidN5
kmzHA5KoKRk5AfBOwynuxSAFxA3MpMGKsY+zmDcg0RxL/+Z7BxI8a5Fa7zPGn7YX
hpcgScbO8Be30+c6di4SPsozPLEX6mKwCEfkjcFEZ1h1Dz+p5MleGiDVknOWviCf
TtyJ6ocfKHAgvhHLJPf1rVelLdUYjkspRhogQ2US1qBSAXTNSbTwgWhmXdUo1mtw
F+f8HGoPuSUYxRaF+CdnULX5CmjMjQ6R8TBCMdB+K404P6hKDDdwgvOxuHnk6BDZ
n/tw3ZVM6ovtQI04GKK0VuaFHewKGjSzY2ly5ZPEAH5lAdFN2U9ah611me4nk/+Y
XBvnqfe/RLDlGk4yp1HdJVKzxiJwS+OfowW7wTKreIeo7WIYZUJ5bpRHvOOcmle6
YPskEpJK17ZhitPwdhpne6+X8rvSaYNycOVGLfGgkUYxL/PHc5pMAZpCTiHSJJ/Z
Fm6E5Hs6G4Zg31Xizk2QEzv88S9WJ+kM4xBGrA3KNYoljidosuTNuCM+nIXBycSn
kGnZJrcWwmje3x8+TR064wywkFdoY9LqneQTtW3NPwyu2wbwhkfasIUJKUYr9ub4
+bF+uFtvJLDaEHh/33++W9Vx0Ox9TaZqyC62Nnzds9r6Mz4kkqE8yn/pkXAfnz+T
wRZjimBFf7y9a9jiX6L4MoeiSj4K6ad4AgnsFw3/6fvi2+10z+Qo59/0KqVLnC6U
9gmiqh3BWyBvbEarUN3Hxtmwq913QVVRNGGfmwRc/qd1gK4+BOqkDTvA3wzesAHL
sGKm6gFhDFQqI7Jr8vqicpTJiIvd0xuV4AjXhcDkbBiH8aflyQ9GIh3aww9CFTzM
6wYe/aRowW+esMC5jSh+SXyT17djoYjulxXTxKyuL4bsUGjqEUT+u3hKgqQ9cAex
b8ElCUbpBkExvRLq1v/dhO8/aZSbGAdp5w9eca9fTc76n9SmGtfdWJH5fsLlKLL4
MYWvyEaStGW2WNujPlszSW527exKN5D1ArRk6CmJir9FN+hHx+aagcOxigW2x0lZ
GIszkz62GEjSH8KmtcDqO5OUPuVqFYISNGrH7YO0qA6bdm2yinyml3kgB2UGK4uU
gEVmsqncGGh58Bsd278phuxZXAdgrQS3a0dgDm05fqN35QZWKPIoyd4W+7Z1XiUt
HLECCaCrlSQDZ5fmUC3OMkKmCqMP4PZReIS0PNUCDdRz0gKuLTjQ6qiceJZDN+a1
l8Zjvvctt0DXF3M8dUk0Zf+YQz6Ac3kZigpVDEdxQ9P+6MIXO+t3dWba7fAwpcW6
JgxSmKFjkOXmu0GVQR0X6uCDSE97od8Pul6kqmHiZcjFXyPyvHOQUklL1zZpAgd4
LSRWYZWaSlzqvGVKgxCJ2n99tlkjPxYWlI2nND+t3abdNS5uguOdekyRtUdHocse
IgLLJIPlQkm4uX0JbJ2+64YtTP8f5R7CEsr4ODycBw9pT+rXD5mvwd7wZ3B8ZyHT
BVpBr9RBT/5V0kNJ7mrhbFb0vPK+109icPNGHGDmeHHn5QxoKzZjjlJ4zEZ/fcQi
aIbG/Fk3fpG//hZgs2RzcfwddT5aGoXDZ7VeNfrlDcgo9B2k4Ucn5FTe9ZHN4akU
Ha3oGSD0Fy/v3X5eWt0x9wi8NQfZTfzvXG5LOn+Xdy4eETZnRMKl867NzqT44GnB
EwZf6iFnBSCwldXdOIglx/EdNZBfdmzW6Ifh+EFldAALjP+qF6pbCa+43JZil9ra
RoJVDThfwyyd/ruiRBIcp4vlOJxewhtBk4g9mVA+/TljGSyZZTzrQcCN//XHFeq+
lrqiduEM9vi71mL2FZMfIjX2HT1+CHkfxeek/HxvqjaaSjoDFqJKrG1hLgNp+8aJ
5GcWNdrCeASCwUU+eQcFZFY9S+EO7LSqYy57wNYGIa+icUpqbC4Heseg/kkg3j6q
FPG264S5zuSsVGT3JH3BFNCXctGzo2Lag2vFGUjDEFUD9cVFAqOA8gSj/xrdVIr+
YPuyIIVueJC8FKZUr4GAHIpBeifygAYS1YK8NJ6+V5/hbqkI2VpPXMLMttcAXkXG
zD+eL1c/ojsk08c7MFvRXTcHx0+yF4KVzpw/0EuKVERQJ6/KxjZqWZLQw4qsjTrq
RqxGcyR+hokanRr7pr/FFfX9tzEtOkxMKtXkNDtEV3mx9dBsDV3OFEQl09NObO56
2P7fNbtiui/Ff1WXupnKErGGC52wjDIJiUTlgPnUM1CPm37uTnVU2h9vVdZuregc
1iAvSxnaR84+m6nBUKIgwITPZv1W5bGxRhTubxnXc9hNQAyNjPnF5ndGmWF0pwU0
fJaeRn6KTAgHh4GgQM2k1seZjXvG/MJmDFSx64SZ5EykrFijOYx9ztHhG4ra2n7S
JgUr6vjp+snrBcXxSS0KplH7W9Bmt11GGGsI2I+ER2CgAtITHsMC8dkJJzsSeeAr
xi1JsDVn+aZBWUZQEr3GtuL4Xsp1ZFJ0o0+cjJih00Eu5hWMzDTiGDrdH8qtKt/J
7oyUoJmtZuo7gDO044tQzKu7isJvFJJr/rZ/ZrXEHdU26GPbtW57+WlqgK8wFujU
f3QGmrbGMIejGcvDwpypJAjG/08m3fTYD/ewrsGYcEF/h2nItQDWDtsJ1+GZZOzX
o6ll1xL41dBrtvhKXPfDP3WSppBQGDs9daal6KnHNNbz4uH2Pca60cLlBVAta21c
2II3rRKGggLbMIDR9XAdJ//fB2aDgDFOcqTyS5n+2rchaUjnxUxMR0M2hsNQUftX
2Av0aw5z5xk8cFkFypIm+yHfNbI4cwU6GSgWwrP75Dc4eznuQL7mzj+RZxZ8OZky
AAfTjSGLk7ZljSG3x0qEa9EWmZc3KhgeTKW3bFQlSJo3Jr/bIMfUVhKYE03LFs1A
9vbcDyvsS76X62REmbbCF1lOw1n3LvnEIuCesRiQRUPxJujNzaD2qwk4qMj23Kk5
kV8BaiFIKrorAq4q3Fc49hFZsAJ6xwirtsklbIOHkW6SyN8BC5QZBPcphdxht364
b3MzC3jdyIE7bqMHDVOE74q02vyM1Pxe50ubMr6lU5ikEsaJRvChc1vkne+nEjH3
MjHwTrW+AGmtfoKFfv2J2Gh5VSFBYBXSoyzShpzKtNrwr61OSUJHHjE6B4kiRxV5
QF/TRJ2Q10QztHcBFRnTV8S9Qu4xKKq/zFCCyttPQVTOL0iFxsGNwBRSQe4GMXQT
XpjvAVXm2lKku4aVowjnkQuhexPpzEcQ+F1LvR8cOYWHwJVyAb5EIftXidUOvtEf
M3tx+FroywTZQ6QH0nc0gxmmKoCkY5GcPeq9cdfy/6SoCbBB5UdvkkWI9lTTLC7Y
fFTLeE+/D3GBpgwuIcG6cGQw2Ee6b4dtDmRcCNo1++rUJTSFwaeKT6BcXwOBuRd3
VIUoGRSiJyfG3an3EbrE/lb8s4m6GMWbTN72o4HH5iypW4ok/K3yi68eaqPx6qcz
zCiUIuSW1taPZygsJvPb1cyJS2SsyzGqkP20Mindrf7R2/o0SVBvcb1ZoGcCZbgB
38LgI3BUl8248plD83aoqEYp0PPovF05C66pBHfDFSFPf+FoWgRJGXpWUHZ3d/nC
d8Wg52Hc9/9wcMDHFgC7/ID475v+7LFs8+sfvh51RWi2vcJRse6qY3i3Di1mXy+Q
VI/75EIuEfPYX8IM49GdId0UVa6gM6vzsuiu0eIA1fAktxiDhI8Yyu2+0ZVwU4YK
8sJF5JNASgmi5Ryb35kMzGjMQCJDb7MmeEciJJ6h3LtkSdDFcLmETP2SNZ7/thwR
xrGHc+NSzQaybr6izf3sWtnfnxL3ivis3Ysjvgd4gLiNIx974zIndm9DZzuNoVhc
TyPkL8rv7TZ8sPwoOIzaARJ/uF84kdUy4ZezNq/EXkEQ6ftJOndSbsD6Ecm9R1o0
dM76PeOP2l9+lufs9W8ZI5gyF62qURVvPkvnN58KBEfBpBzk73O31sm4PrZcxnlb
RCp5+vsg7BTIS24HnCK1T/Wb9m/yl0K8Rg/rwEitbx1C8JtiiHixH3FhKN8om21e
uSmQglPVj6Twm26Q58jubQVhTPYttLdWUFXogJX008+aWbE+JIrV8kmoBKMWBGVw
meFARx5bKNaHlK8YEMBiIJdWZUuaHPdH+uJVPZX9DLNsFO88xshOQs1gDuv6nbsW
jNEwdUAZtk0dHd3xvwU7oAxDCg0XE1gwoZvuapWKKHqnkNkR35utBSgxq/xrBM0P
SYPXsQEHPJCY0DSJ79ZbxTjUHGKf7Qznp+VOziYyh9yK1RuoOAFKq1DKLO3VjXQy
Ja15f7jnddLBIe9Z/HhuTE+BFagPdTYUUFTbTfRnb1IxQGUyFdAOE84wFptvyDtd
GX1LZAfnCal7xxD7psRDX00ZFPIBH9UGo9Be0TEKM2M2tw7GWwwqWWZauyr/pB5x
uwjvSL270noDCHwjxbAaXUnjRDjTlrS/eeAWtKPSDmS9SQU5wKstQZ5BVwfxRG87
iwSiftF9OKbtajbWdZ42o70p7wPkg52RtRAKmposOwT1i8tI+40+8G3GcDHmklZq
N3Jwnw8oWEZBIpa6pOwgpPS7J/UGp0v4SlDZmUK1W8XLGNEkGj6hntJVaMkHWo8l
lwkGAVp4NVH2u9B6vyNMp2gIFDR4yIaKBgXt3/4GGYPXdK6DRfLc51cpy7e6tYW8
18MPpi+TOQ4jCUPM7GaOmcHtD1dngy16qc2nwS9HTi27ghrbO5lO8CsicxmVVUy4
yFgXBu5knxsG5ylmOT8B13MruMGTvCY7I/LjJC0hezYVUP9gu294VTzkLALXAYF/
D5RmnoH2FcQvNK+O1eYJwu1LxCCqJ+ePLfa6T3lLYshsSbjsD3JxWQ4f4RDr1VPX
nyTQ0pQLlj6wPOBa11KDH3w02vYQUQdkuEImSL0l7laq5RV+ke9KEFSXd8kbQ/5u
wfjSkEibMQbAcxA5yyaeTuQOncgS3VnL9Mkw1sTHfBXlZoOSe6UvVkrApZwwPFnL
DuFhPQdyvm43xLeq8Q82NbQT5+v5bef9zL2Jq7p2aJ+0j/OQSsZnaRI2qgqpPK54
Q1ctycWb99CB+h1Of2qX+YtmN0Du0JFEYMpyzUkYPa+GJw8KQhq9CmHgYcwGBnsq
AdMhaQxuNo1434fRk0qJdVbT63MUVkjFqZdAWTQByrtC6lieR3kmXrVGLsJZpqbQ
nI+UOvsLcqvMMgHEhhyjqu5lUIiuv2J9fm/Nd73o8lHhehrFJbgW3a5ttQpr0bhQ
6P+nZFmXzMcGtsT0Qf5ox0rvYkBpG1MV2+sVX/NGQgJrxweB3PWEYyA2lrRzwXj1
iIARqGu2wTaD2u2oVKqSPR2EkkqNhf6oWJWsvCGQtqYAYYnsSIl1T0nqB8KxZvQu
+2jsoix0pblryGF0kkhtg6w7V9FRTwqtsiovLw++YVyUkQYtSiG2sDPOyD4seE7L
H7Gu2I+G86hAFqhxvCtiLlLdCjXvHjw/MLjxJ1VJhAMo1xZ/I5MVY9vB/K2cZLVu
y/xIbXwH/4GLUYIBZfXCENpqo0ngyaf2hPvGHwWkE96/NFajjL+Lad+KQ+WQOIIZ
fSX4YyQzkleqmV65t1BRxdiRRVJxz5b/5n7j6pQp9wro6VDBI5qzgA3+63xsctnJ
0HKI7UgRVEnUKKlSjBrTU3By9dtqhYM4g/4waSU5PFvXGN/NVpdvZ9jErNN3vTxq
elacXf9P5Mmx2aiCYMqyMitM0TJvowyUnqdY1SHv+mCC4mn5e5q+kkhEp7RVd3JL
TSBfH8TjZ9Jp+AZwzCWjgn+VIItoADlX9vhBgj6pnDw/21n8IZAoEPlhjAGu/3Zy
Xp4SsVV7VrNMfsZWwErBk7qdAEz1Bi0rvaZfxmwVKwMNlXYEv3WznqI9lwrdhZbH
TucP3Szjs1JIyg1KPH30HzEUyPu+t4L9/ao3sn+xHpPhASzAbM+RYEShQbBq9Krs
rkbzp9kPDG01k2OsL0NQAS64lwNgliH6NHA2KG8ar1Aj9HG++3c/9Jkxb8tKIwqV
OSi+YemI3MaiiYO6Zv8PBuuPavd+1tChVxl+adGbXLw9auXyeBux620ezLt6NFEw
N/yxxd2gm6rRJDcWyKPSD3NzirgXL1IrnKFDmLGkvcq+K+PlKZ3ZijBUukTpZEN9
vCutI+sNwl44iF7q4CkLg0gt4vqOVEuwrVFB3ME/hBLp5aQSyb3z21IKm6T+ej9X
DGKekhR9b2CvnOIL9/RwKakZv8qRNOlsYJZzeoQrk97HFGamcjTxP4ma2EmX5Qw4
MlirDh6Uxrxt1og3bH837WbunF0LCwIkOB+WKTEgm71vSMiUAo1YdOPOl0UqTrkZ
TiJYewkdMW6zad4IcfjLeD+seY6V4Y8I4kxt9x8Ma4vm5giIuiZ8XCA7wIiG1tqR
YJHK9XHTTdBompD6sN2v9GozfhE4MvQRhUiSmct7NCj+vSRJn7FlXV59a4UvUbkf
ZGVor86/GaTh86eDOE5MA/gBUILxrl/1Ep5S3dp5zA9CZLLBkOBWM9UFY8I9w595
6xcEiNn3xk4ZMT1vYTYCIrISoA4caMq+TqrdE7M4ovfW+UTbAfsNYuFQ4vjKEzWo
nIZpPxvkiIq2p7HjGcBnZtxr7SNOSX5UqETQ/MMW/ovb0Z5mI0Xli4akJhP9FslC
Mq5yxc8/qF0Nne0XT3KvCJixxbdidJ9UydRIg5R6cJlITrHGHTkKYNE24F7Q+vYg
yniyBhICkL0u/8JrZcWPDWt0hzKPsA8zBnimB+QEkOHIpA0m+eaH1V0imeksV8sv
D7ZTNffClvL32V9IJgC/dCahO7CUvahVnfhVQ6bIJYHel+KWOCEbEKp8wW7nM8o/
M9hgx6PUfTD4WNDSzZ5+K5EzZd27ZV8aHdw3bH6TJekEl0K+UL5uqjaZ3C1vsTuC
krgWv20rEsVT1i4uVdE38Nv0awm8+REObiuSq5QiDbdulSlYFXTDjM7+p9NRcZG/
iUbvlDntSrxg2ZEbHCgwNyxOA7vsN2j+YERWrlcE3X2Ij8JTtHq2Ie9bczSBCGGW
qgOp79fSybv0VlaXwRzChFNXFQ0xfqAkMnQmZ4+8Zu4yTkgFEximYqLJkdly06qv
EMQR8q+syNQ8glguPqf4ISyzkP0awrDRhRZbH87TXK/f6UWdb5vzEiERvz2CjaeH
fbIqEkl5GZ5yVub/CaXs/BKaNWgmA/R7LO9lSBz0UVEUIHdnwX8yFOLeePlTCA/Y
z4VZafQSS8bd7lKDa3ytms9mpiEScx1vvpEVwtPGmxEp9oIMTU9xc2riSMXflFSg
EcAKA5F1wy1aqolTKN2uYBrV0o7PMc+hdtlL1SSPVlQu10/MggcdhLUr8PKte9k3
8aAeGez1T2BGXFv5se0xUo7S1nSqOww/9nWni/3rYd1BSBLDKu7kyqQOq/qIsDG+
JFKcwJV0HKUJcwWr7cSVDVbwBgYFyedBrjy4CzKbjXXdrFYaawDp37Fedv+Yxldp
7hQ4rfr0lqUD5QMrv0tRX8ZdP9ghIiwqD4tY8E4/jleyhxOrj8KOM5OW2Sa/3si5
PkGIHaDbxZmZgqfQTAP1JS7tGLnyHOmXyG+XRJJNz6Wr5CS0/9qge6dXDyAMV3bN
8RK3ZpExqr7tb3djgIeeN3Sur+InJD+AioScrjeJ5a77H5IUh2hlnLVLGqXLYM4Y
91q1W7TgNka4dR9CxI3ekudryJrQUVTIihZ/3+qmMJ4PzLnTzpS/d/qYcQ5VY42c
2q8POx9VD1gdpx9gJkA29t/ThVeOC9aYnHxe10hoaRAUrSyvgX/CMiMpgZsxK+e+
PIZ0GXHg7lEuG+c7EzZA8Ah6TdKB+30FVBBnr0LpYzutmr3cSkXq6+neB+5SeI2v
9JFyN5ZFMrfilcUiYZyQaVHCyTeEyywizGK3ciznv27Fu++nnafpdRBXFgKPjD7Y
0FHvUADSa9i7DVqplODzvK1yriRxP+rQurnAhnT2WiN+I2G1RU5FyvKlEW1xy1wn
aC43KtsMBDh/ACnQ7N3TphIGbGcHNO5Npw4hy6g/qvKhLl5LiIiCjG5jAAbHUNM9
Gnyp3hk+TkcZkDyHdth0yILORZ9EXhtuiz4lG6cicDinIqr0c0niWGjIhKmNDUH8
keI3qrF3wJcSbrckWcfSYa8WsQNEC3Z0wLnx8axMzVRBndLkKWizZvA1kAH1C8mz
OLpoMfIZbeT/82Ex9wY8u395fWBpubW0TK4LwAK1jb6kcjQF0IRiTPUtSSaPD+cc
yxqAGQLEFnJGLS55V6TbC2r4/NtDgwn754gZEqun91F22lzKjnGDGSoEJAc44Cis
ZEFe7lTw06cT8J5RhPYUVXJXJ6bGi+Z+r5TAI5I86cwsWNWQm4jyhuRhwv1OWkot
vvWtz/GXND0F3iW9LkRtQKmxdH4Hj5jvi8TduJokHHUEkcocppNw4wGfvaxKatKe
J0057UzsKNw9trDhGnWTK9hSmpIIjCk8palBJdtch+2pYkOhz8XXvvhU9JUjit3+
OH6cc5gbzrQMvhK7yssYEup+7J83mGlrxpYwwU+iDnEws86IjiytwItgHTszQkRK
kQsG8D3qFoa6TE9jmGOWNJRbeMVlkR4cHAwm8bGB8CBq9scxO6jegp8eSLC6wcxj
mznuGCLsHF3Vc+J3pWxrTB5zZQ9uBr4ML7NHHzavrmzHzLcMx12jmNrGu7c8YY4d
1mlOcOP8Roq1wpZoaMglNuA5k7XXGeLodL1zbB/UBEszZ14cVfP5j24VsuYh2OY9
yWNxwoqQj7xehKmqgWtO8dZ/D9MNmJEGK5LICnJan0U4k+SxMELBDkpLmSUuXZ5Q
9bqEb6L+vK5JRd7IB/zOEo3p3UZiB/OVOBKUo33we1iA++mdxLqiZKkXMPI4AcXu
PJ2SdBg+DC46H5FnoKUJwaYUloovggOyQJFPt2fjkgIrAvxioJiOUEZhkdacrfOK
venh59NsGbFqujYwhzv19UDcMIcDsArmFzHx17uMVFaPazs3yJ8WkNwJlH3jxeQa
/njerZkeNhirdrv/PX3i5jDflW+GoKJ/fkMj0ovDIMAKdwUpsceEUP18hNd1rEm6
LJgBK/2L+DkF2x88JfF5XCTgskJrTgtVioPdgk9vQDdy3+q+ziwxxXIQTQlkazEj
5eEwbEuJ/IElSlSNjoOBBir+MvdK59vbwt/x0BKJExURuMhgf38D33WJa6ClUAwY
1C+K9WuO4KT+5lxqnlgRKNYNni3EX2H25jrbeOS+18A8ASLmEjiz+9LC2MbqFvBx
yOyxSX6hdFal6uhnBkFcB7125d+VU3ZFtYkUaDIWHroDczRopIwjXUVa4huEsZR9
lKQbr9N/09IescVom4Jhw/2RRa270s6KjdCGH2Hj8Pk2sIqKK9Lwu45BVnwDOeF0
v5vQ2ew4NmJLsBQJoueMdL/DNxzqIlRQPp0JnYSeh0acmI0QRO1KAbZ1cX4NLUXS
SOFYRP/F0OW6twre0y3pkBiceHx04lzHqo+qC80jcDVOE/81jqv1y1iVWyLX1v3M
bXPW0PfM+gk3wGYVtT4Br54+NO/gE4Ta7VIb5QkHwUwpVr3JL03H+UHszL74vzkY
vQ9TJW0A/+XVU6JHUNTVWHWzK4ElsGVq5zFUoymwfXOrbUWNJd7b4mPjGtLoUAsq
tea+WKqU4zH+OtNFraXMVwW6MJBVvNu1lkxJOtCYUwoV+w6YkPOfVwl96uwSOIg+
SFsbu3MALJ7e7KaXL7VA1pi20qii9rQuvDJj6BfLh9zq2296e4zxcvOw0+qyMj4k
5BADmuWYAKFIiqdn7BU+sloKRdmLIhPv/29P7voTTIzeJ55zQ+1srFcFZUem7V9B
8wsSY8j969e15TWJL2eIuelZVgUDGOBGtLtSKKc/75AFVMSSS3THF8gh30Rl21P+
1Az3B9YmPeYvfUhM8ucguPwJRv6yaWN7UFuVt8nTDqzqvRH46eQGmQOhuYz9cSBm
HZAqKEceWIbAMRAcCaR6cTP5hyr3qlN4bcal9BXl4C2ik5KBseWrJra3Sx+l4mgL
LuasTCk0t0ZERpbTxcd41Jcp/To0Z6fZt/nMjRHRi1uMDGWq2YdtezAukjptPhPI
itQQeubZslbprIMnlwHKx9tvvc9hqXNeE8v6Sq7p5H0cmBB+Ae5LHtDdI5AZxfNZ
5Wxkp25tR16zMIksZcOQtOaJWINj0YfAklrMW6RlWd5O3X9kjdNpbMPQ7PJMmWq5
Y5QWd3oGaF+oXuX+j7ly6zng2pl/rdGUg2TrnBfghsSPbK9lnPOm9WQoTJ5LUPk8
Wv8Bbn5XiNRwxGgh2aucCOdsRXrHEoElywerDUdqB25NJDsmrLQbsnacx+m0bhLW
CAhVvF2mihKAltImlCztx906ifh3J+WKB7FctculXBFCAvhrsosxlJwIcS9wvzJR
fkTrpmZ76B+GgFhG7WC1ndGJv961wmKdMAA3kkGOaWTj2qAqA6w6R6I8BlFuyi5I
xOz0xzBBdDnUkhmrpJVAmDc6wkfBnblfac0YN3cyl99CRLw3Sc46yFHIuHsz1oZd
oDaWF3k4HG1GLagNuSqwDVas8Semri3e9TYTvyyOXgsrhLA9QK268r5PmYtrELIq
fZjjuieFeuDAqvX00E5P/96vCrFlKgX50owSgoonw9t9bQde4LZstsvcTaXqPr+I
0AejVSyqnvPXWdlZoMwwYiRhxkGvtJASrerx9WbzPm1PA17hJVWtO6XKLdXZ2t3L
HxY/wmM++qMgfgQ+KSixPqkxQp/LbBaA4Iha0qOcSmMthUhC745utLa5vXtMtcDz
JUP7OZmoxEd9JpOixGj0rFn/UFJvFE6GDNXt9ZJcrM6FkRHqJfJKlc2Tey2VOsjj
4EBF4Wnv3oQXZ1e/TF+gWVwW+C5+5QsoibC9a2rDan5DwHNyCXwgU/ZZ5nIdicBn
oP0ONUulsyhxAj7Lz0R/DD7j8MdIz35fRJpcbPaOn4XRd/tgqVsT2fqeMTD7kTPA
MvvXagZDqg5yukmNNXnHA22BlsOERWDN/vp8CKcKWmtCwdHstSBIcybzx1iJyr0v
heyAg7Z6E60M2S3Q+iax05QZaFhxTGq8t1JF4idgCQ92gLj9XgXmhMTWRKeYr6n6
sg/uQbmVOs1LDWlCzLfAZr+S8z3z/ij02ksLEk6ziJ7Pe7oPV+eJgiawoWlaoSQf
PmhIy8xY9vZ9wdnkQPRoV/HD4BUtnsnZwPL0r6F9XHCg0nYAJArnnKPUdhGZJ7cD
dGHPlbM2P9DR6GgnYTuigSxEsRMtORTtYtKPNSf+CuhM2v2+gOQiB9hkppaGy5QH
CsBq31CmefdMSWYzmDt01CH3bK1eiGHP3pGn0ZPRPBSOy7uYmPgrvvLQsMQcERXJ
GooYYncV68StficTDGy78DxlBMkN0XZ+gM2bQOVQJ0gTTciZ8o6I1tVWyXu4j0Ib
U7+6/k5uZ/1oXSEpHnJx60ZIvHWidoMVuNOhG+qZTifEaPw6Rz7kt8wUas4uXZcO
fKNfqRk0H81wgus3at+rw0O70oNm+Fg6c8g+noZyv9KfBrhqKuB/IEWURtjYV5qz
7d65uK28OZLCJuL4imVHMjv4RXUwcJf96Qy93T7653mph09y8s/hkDkTOfEQacs3
ydzgnKetrmZKA3PjJOd5q1K72XHQYOX3waCRlH3uG0YPvaTFUwZDotZS0kYPVf8i
9h3SDVkjwDbdTidlzg7xUkdf3Q5YOskzKK/0EfBGQbVYuZ1CzAt1Wb5XMKAYz/fJ
8XuCQ9X8umm3AtPqy5CD9/0tww2RTdxiyuRJWNY5kyJFZJxd2zc7aG2W+0fqM80x
lEu1gYaHbLz6qrUBORiZKKgeMKFMcYdOCVtFUdvILvYFcnk/4ugu4d1Sh5eWcSdH
zpWONpYccIME2oKPV6KMsFCCn0ipHXyqnzJB4q1zXdo+9Wa1aLyWZKPcGYrSkzdl
JrHoBvv4SPucnl0vdIvkvWJ4HEii2RkdCEn9PHnEoaqE/vkNouR664/+P+o2UMwb
z+J6objavkoBe/jj8fAuiOZL4+2bFuDNEPA/sYa12Qu5STtTEiWdNgaogohxPfRF
PlvuNA0Ye2jlr2xgvaxOp7bmx3rJx3ZcSIbNJU36TlDXUB6n9TptkuIFVQsUr4em
UIm1mMa+t6ybbirqdXT+OzkP42fkfbZ+PRXSWdFffiUpvw2WufueBUrzPJWRkVFq
drJUMVmIKAShSUALU1WLFUU4doC2uabM61gLCLSW1Gj5bBe50F1lLkKweAiZ83ZK
lrpFrNenQeyjeY64m0+2mZHAPpf5uAVyKT9pp9vITBS7QJX7PQ/Dp6VIOSWZ7MOk
V11D/BCiVATxeW8eIUulYid/VUQot61TQaEY1w/CXpqpnLgJUPso9bfLaqLnngLx
uiNiohIhFV70mVDfYnaSJfAhjwNNnaTMDXOhvoNSI4b8ECcWmhL3l0yeRWR+voXw
1lsoZYXJ32vhflLbCyrTBcB+vx2/3sYj9OzznaJlRCZpO9uT2tATZovHvDgjCr2K
OB1JKele9xbzNeIIdOH+ohWLbzHbVmpvBCBCESBbQe/nw1Q9nMeN2yoSVNBYa6L8
1m6GfvuNOSf0MyfAKM/ClVn8LsKErFQcJpHVzMmYCGt/f2dmX7foKXSescvcDpaD
QrKUPsUHZnVBshj0S0bTNQbYOXyOt+JkEx3JRJCqDg0e+mFTBcHWRh0XYECJI5+q
whP6bPbm+MmAqcxBHI0XNfpQI0RuixzOdJwPwFq6lysNsGmKd9zWHClJ+344KSlP
5XOF+jlrpuIR51/mSLjrRrJafwIXwuAiZsn2eisqsCcuK9xTt88wGJNNp27clmMO
WWdPYQHIIR5o2dFQ+ZSn0uGV3N76oVcFy+T/Q5w+sH70+MTLFvf0eqZdnL0mPD4N
AGsEkcmtcUshcZ7SlUfcntH+k5DPJra8dRRj1nhNi+MtaYcAvRq7H662LgBkDVRN
wbihKqYGlba+K+LAJiNdbpAa66SLaMJTXM61JpjdDLFR78hAUFYmLRpWnwyySGWL
PL4h9v5NCOKUdJdjLBg+agcsn4ROgKxv1o5BlRkLT9Nw6jtrm1121NTMcqzQQLzO
3il7U7tf7eIpn3VWc6NAF6/zXpHtAcJpAR2oXXiXx29IOlIIyEk0WESOdpAN0ZrU
iNovt0sgMPzwZOnIF1BL6CPFUDK4NQKJ9fFJ3yrKlydQInJHtIA9qRjeu8ZqiW4L
AIGA6NJmKMDgTE6OBPP5X0jh9mI1nw1HV26blJNvsncOV1IjgGeH6dL8urVNCa2b
p22Jn7scKe2h3/4Lw8xA1BjGat1VmzHJ/dSuCuh9VCsoUhFfGWwa08RwLeJ/VV/J
64cQXaw1vchk5aXS6V2fKcyP5MPp3/C4fIFfhkBZu+voVAUNVMKo539QTeBVHZt9
Xs8rqWoYJETngeqeVwhNzAddkN3pLO6Ai3Isbb0BfLsdKBizIBdxLSbXE//W6fYA
9pdsjqKt0JdCr98k8Ahxz8ZO2HB5qiE/qaC0FI62RebNShQkJg2g7U7OHDbrBhZe
rQ3ByIdxxZtjX+NY1Mfot64TbPKbGgzpijCpjW1vNQO1MMVia1fp8FCBqwoNv2qp
Iw8gPHm+hgQEBdqcyCEjFh1AoZTKCHYIW0G0JGVgrQErDAk7CwoWPt6f0U68l0/B
RzNBErtqdczqQFsgL5k0uO50/2av6XXqr9taeBVx/2W9WHoDMxe+fsbaRXc5K/po
hVX/JyM3kz4DeL8hVILAvyW9Ktd+8MOmpXpSYc9NmuVjeY9Ivi/mqQG00PZP4nTl
OeG/iZ7HqveSNEELZGtmJry0V6T5VHdI9FQLJFxXzB0wqg8Lk1lf6r2g8rA3paNJ
16aV/RPH5r8RefMju5z186DEEVcIvg/XlbLu5S20zTBi1GVgnB9ceMbgAPMibNKi
NBgC1cXzuzGAV+oymeRVpXXs31M+07kssBI+liFY4UODSDlKW337naNmrUnUhLTG
aA9Hv2S1o1omQKJY5LUE20jkbc3rBq6qtoiU1x85ZUXI4mRP9RtXB6uvD6u0mwzv
3htumRitXde7BTl4FuVDCdtBvTnVqcNJxAUKWNq1/89Ct69SmMLE84q0OGGrgWQo
DhGuVyRiUufK+qCdqwUtPAMbihEIq1K7qfJoKZKpU2ki8800cAKuWzcCaxhA74/a
CZin6T7fqU92nqrRqS2Vsy1vUNV0Hfhh1cagmnp2j7cVfeUxsbZiiQZvkwNjoTXN
k5pK2B9Ft8KvvvoSMCWffdmCIzlBZC2KeK8H0/ee0doXdWEnTiDsPdnE0MFlq7+m
l1qyxzKLwwEBBI1ceJJx1t4xzHTwdR+pNn1yQ7EUTQ4FseCozv8fr9sRAFDEfIz2
Ea5Da2WhdPS5jpLg6UH0zUvE5ImiAlelItb8Xp/S2kn9WrQDf2pUeMSDK8A/+Tuv
NbVEeNDG7wi+XtlctuS7xpg1yI/LMOv+1ibJyWXMunGQmDFRpYmBeYqp+0eHVaNj
ov18NoYGS5JFtzqBEXHZJoYk/JpyfQ46p4PV79NM8tkUwqvzFRqjoapO0izFIQGd
Seow4rTXUzQAvcqIFD9V+RxBX5TxosPwL9QNeig4SztYuAyoeNe5K+oSiO9ncHVl
jSuFzTwcdtdx2xAtPuG5zhDuBh9ERJQ2OdvQ4ncV/nXZX7I3sS2GUq2PVcAYzYyW
0+JzaHBuK8p23CA1se1mtGJl+7VWprd2W9JeqtLuMnMs0+EUXjANTRkK0jsIci5P
MEgyNNyO9zAb09aNElMW1VSYkcCtLSi9Vq5TbV33bpI/Evw6wfgWOEG31uDm5Omc
B9zdTGJk9Q4OyOLuXDINyUK+jSrM0v5kHiAvpjur3sjq9TuekFVPLpudZ4y1Yt4+
9nJbyvGXJMeUK3Sao0+mO8N6rLHvEbGRjRT7pFrI/21zMQtcxewIQZd+OW8jQsW1
Juo31aXssHmSYO6XCivLm8IwdK1f2ympISl0UGF3BMnQ6UFvoWawEnxscLqMvsYN
O5FJI/de0ZRWWVjnzNaQ7gyzFTuSAu2CdZmV3bXk0r4dV9J4ILtNDalYHk0qmgxb
736q6J8jfcmr24WsbRClQVvWkfkAwPfKl8FfuSYO/EKs25bpYoS6/Dqxcyj/Hm4G
mf4VB1t7vD9I2jNYvYpaTrDYAvqCEgeVAzz7d4YHt6gmLyNGmQs0JHkGld4mRSIy
4kMP/jX+CErVkUnk2lycaof1vO5YxhWwbGJozKyv7IyREVjda20Iyo53mlawT19v
TGr6N4DwI4xlKABC3ddQRamYrP73CkHTdg1UmM+FJ73uTy1wWMwWVACLM+QPs1eH
4k9Zue7Ex3qmFX++z4jYJG+Iw2pMvF5zi4ffMs5nn3sSCuU9KCF1B3dK2EvxaYGN
Xr/u9FpKAf7R4B7Ne4Yr1zxDptVLObffFs/YYamHknnLnopyl1dsKDjADxPzgc7R
ak6ghr3QNQjHzwbrzmjulpwMI6PjTIqBSedvfphUIA59x2FCpBWVgnjT7nd1Dtj/
YlRlo7wjwZ9OcVkxE+ODyFEZEOREUp9HZvm1/UioTvoJJlBZ6vU4PHKWwuzHFxNd
dof4JwCo+kDvrUlEam7rn2bo9hmmzWeyQ3DSuAVydI3khbNeBTtd5MYUvkkQb6wZ
aHD5BvDWkes4SUP7iFqVCXZ/0SHvc9PfS6teyaaI43lrB2eRSKhhArTlWd06gRB+
J1t3Ay6C42/htZmNjxMhoEFpua/64nID+As3gHYg23HbfIud3S5KRo3dTyXmGWNj
96NssGemp+FGZinDtEWykvoQ09uJX0UPXciRmJ/x7i0WC4BY+hncG2bKGPcmjfG9
e1nWKSE8zheexLI75Fy79OXDOhC+2n2Rz5knyRnrtUQTwcRFx9E9uIYKfVv7ze7Y
smuU3WmeAcaZUp8dxqNUxRyKeU272JlWlQC16SWpwlz8Q9XOZwiOKKW+L2Takcyo
1b505+d3ITs+7st6Z6lgWOS0oelecTcn4Ndboh9R0/OdgwKAskIYvOsfaC+VZHJk
czZEgT2v7fWwTTU+RrNWvsW9o46FHVXczkm0rVC404jHGVg9WG31nrePIxOXI+Mt
heCxcx4hVP1ymYdbVzWwNty6mH141ZFXAxCbhkFlWrZi+ZSqvmAsxTOxhnZOrOzY
BAEPFk7tSBRzy0w0km7tSD4XDFxzHIMQLEl92yLjGaRFvzebDAXaX9/YFSfMAXJq
jwMyJS9Pk7+QjDvcxYUBIzt4IYe7SlNhC/MbuuF+aMjbvSWNodLNHMQwP6I7bWeX
koSVrnnSp38RCYfQZIwJ8vxWRw/zUvcs610GDyXtjgA=
`protect end_protected