`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6048 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
zZW+FE3QJbCmBLU2wwffRnlYEYVztmeRpkSZxl+yiIgPVffup23DucIZk7x2bqmh
7K3s5Parbj0+cHBAjlN0tRUhX/D13ixaYo1DvlHudxEleGC84jcQ0BfyJvycjMBT
KUaehqF/V0rCc5ked01HE5ukBhosA9Ofq+OW6STy97EIYGu/6/H+FIiwQmuKMd3+
vAo2DYoYSmxr3MVM1JE9zXtb1wH2LrY5saRfWYCVCZphIFgvjLF4RF2pQ69itg0m
rLJDVtze4bn37AGPssOf2g80rtf6UJuB1oZ31Upcifd4pRecphm5iifSLqtxwkXE
Z3ijgiadTAvKpgJ6vMQ3nd6QnCYSp7IqdzVcmfGFMU8DX1yIdmVnatIA7QmWWzAk
8e+l/gnFPCdAe2p81rKNhr9PLURkJQTZ7vtvX9+j7MjFyHn0aNY0BgROr00BIT1e
ijJPM0WY8man0ntFeZjyEgcvmVVedqRzML5IkxvgDPIyOH5qT8deaDnxIrA+VprW
giAxzbypsBU05Upp13P9WXZuhKC+6FddbGJAisa/L45LQfWzDMFmFVivXEF6uvUR
pf5dZLGh9H2mz12ZoIzPAT0ewC8i7/GRkkvbXt7BEKxqVpjbJ53W0idrz9M+mB/X
6LavpnIVUT/kUqk+BbnQn5Nhh6Mu3TSSATWhxUYOsyKm8NWnZwo6D7/QCsYosueN
J1CKUZ1AbE7SDjeJe8AGEGwYKY/VZ3cs/MOUF3k6CPBEicSr6mo9AxlpdLgtMxj5
aZAevR+WLLInKNLh+DNGSs5Fd3HMb7Vn1s6GJKRmB5bIrdSIgRNla5UuPbYaENd7
joPHJHzpg6iw20LHVLVxiMVXLlWQMlhlXSPkk7HVbkJBsXCjgpZBTPkw56V+RA+s
V4kvvPdnitUrE4nFJVPL1sDeHhHb5MDCkNLmJRxjdFMQOXO3NBgaCs3wpwp/J1UA
nQjW0acb2tDhOUkg25IfKRfuG5B/IPkvo1pei8rFHqkxKilU1IYVxTt40U5reqXf
NwapvPlifQqLLOnHGVHvR73QY4DdKIquVNdj0xOb0v6SZZ3E8inCI4ykL/XTjn8d
StIjAehFygYDgjg5N2HAAZWJzqLKQpSi2IDqLFx5d9kLFwf8B1OjXTqyeWQqQeGv
Zk37sXJXOL+T0UOQ4zvBBCZzswimyYlE6jHszZsqZBnBB0j97sFM/X3/l41Vr+DP
hPVdrtQinxMN3p4C5aInrnmZQlfzb3V9A+V2O2CSP/h+Jf0207IOPhnPvlEoMcD1
Li6E7oHDQXSwCBwLrKQPVZBZIXFE8L3NMhYYP/D7jvkAhkgyCz4iZka/IyW33Oqu
rGo6gXyqUkEUksNiIedhomLX+mtC0Q95nOKv4L3Iog00DC+XDJxm4Me8NW4Kd5W7
6djMLaG84tVAmct9bIVzWP56TIip0rBf+6piX5gbp3xtmnza0zGoG/JpUYD34eQK
69pd9tx/rK4ZClty3NtdDdBz+LoLDKQxOpo9PNc67PsboGf1jUw4E1A1/iG2DvEm
YHFQbyE3djVNB5trlhowtpSvWEL69k1s2fFU6osuawqnpOk83cb7cXIAaQzoXHVA
cecRyfJeK1Wks6NXJRRa342IZKdfJvXOa8af+vwpIqIqZDKJtXvjvjMsUOlMgffM
jVHfIKqhAfB1xMWTzPREoAu5/M4N0SaTVFe3y5Y0q/KzW8IbNVn6/awK5piGFfXk
m9Sx8iw6T1kcSBw4SF7FgkbtGx7zTsAveXHKuODrBEq82ec0M4GN18mYHIbQLMn2
+Tvo/k/VD2qF4O0wxOMi4ezw/nY4BghL3ZeKfEtnERGQJ53XiIhUxxmZnWLYpyLb
kyAfK+Rjbzn14BqXN4+qcseuaoNxY2Qv2Piik23LVQGbRXIKkPHx8PGEBoStQ1lj
XexW7Iuwq1K3paLPF7YgNhzSFPXTNkyeWzYwoIQ5B2VYoFzvL68QjRa28bPo1h7C
vrFP0VIGLEViNUnrnoQM/RC4EQ7siH56XwQifWxd7Cn90uBe46T1HIw6Sq42NYVj
dZKKhyrgp895DrNQaSbBOGiP9hfNCGvyFmNePfnhyKP6WSvlYpxtdiE2xjyYynkU
hf7k2r+ONDyeLFvg6L4zGlUgHwskAvbCOtwXFZ30QQLFVvNVskXM8MYaST1Kj/Lo
OLL/HoXRqz5YeLxYKfdvx36IA3Oivx72ccL0F7MiCdTyFDMtsswQokrnyAstyRDu
mjYqCW/r+3BsgY2D7amXBhFRfl0zznxJPab/fWS4ett9XcgYGmz74Xrrc2SW0vPt
pvwyAbAcczpBk4Uuy7BXrNRd9Rp4MgsjzEWJDAOAF+ikuRqu/kfpLnJwZrHs7c+8
RdHNKNFPCluq9+LI7VL0rtQz9hvSkq7edqTQKnRQZpgQKFwQJsySlPyUHpn7yKpl
4EB7ciz7tIx0EuAMjVmqT0Qb8ubpUZeYiiGDBWtZadXvktRkRUwk6k2lqP7J7Wsh
D8ozwuYeLZU31nfoFEdW0PPeNiTwte0HxiNTUTRvj6X+xdbH/nRRTolWo1gEucYJ
ylxAtp5WvdAw4yYf62FYAbBXpI2Ecm8Pmn3JsIoVppZYz4q5Fn81hfjs+Q6S9e1l
eH4Opmaewo7c3PqkuKCzCylnUPstlGz5EnVePhIREsYcVK96Ej9j1dXO8dFQ8Z5d
goq0W71wZaRXIZjsVmY9yxLemNmvCVToMrwIuPC771td44vcI+n2NKL0VpTxsZkK
4sgzI61hgD7N4p8gg7hRkLZjn8XdIQTDw3Tslj+OqoXPlCaoGxHNRmtJ1GZpOrq2
dhU/7K57AsYhiu9WRE6EuArBtAn5PbzJN1b5DAZD2i0siJB8kpu6UDH3IABntFMe
eTvP0deKdsoM3CEwwrA4TzoYfoU2/v09fZQK3QY1s3r5dcxbBwE3wUDh+avrhsj0
ceNl+DVcfgN/nSDEuYvj0jISeiP6tapmwJGIV39S/Uraxx53l342UR8m8if8N5kF
MksQfkMu4YjO3kzVl++8+d0ES46jG6X7QPPyq6bn0e/PvpJP7bw2RNWx8NzCvfLC
3kAbeMdDTiLsjFG1Cjn8pk0jqFdnqEfw7uUhHMzPkIg1Qr8gaxb/FqGL2D/hJTOy
pY19IOi/rMDoBVDmKwbUJ9n+BrLWg9r9U9u0hX2jyGVmrnP4Traf25MytR8FcOs2
h2+SqLNLhO8gEgFebvUBIyx/+jkYNpUJCr9h843YjZLcVuHWtUZiDhdOZN/Ien5X
kyZSOyao7KMJiJc9V6QzTQTyeVKst4/Pa/hUqevjSW8OSkUcYq/8Ld3wfNXehtFo
8sSGbJzyzZ5Wzogycboilgeo/XGFQcZE4wcp0L0LkoAIMBKMgm5AN0dZDHTKE6AI
hSAKhemxkxK4q8bZ1yhCm5tuLAfcReCMo39MiCOiSGgLfsbaIKxnDggalyGphME+
1eujqVeuOSE3FeACsLIsO86MHKSq2/BFy3jyfvCBA3LWRM/PT1ZjK4g6410REF5E
VQJrDI/JiO2DyT+ULJYc9X/mzlqXT/mQqAEKuWmIVrNVFNkYgrj2uDsS80eMa7ec
TF3vuJ8EDTGlIJpFXG80Bx8p1AyGtU7wObhJqtSc65+0NeikP876cJaj9/mfdKHE
rcYD57ZAS64sOR/dagz0pzjANPwu7abngg5VxNtwf4AriGPUrwDOyRvZpY4TCX8u
x0Q106O7tlQdbvV9hjg9wGQNReKO6bhMjusk68G5zeZlquLrypMShzEGbhOHBQMd
b8v29v5aEtfYeuVWtLwwDOSWyNomlMyv/OVaFv0bTK2hvY4mOyCRkRjide2SnNR3
7DOEXNvJVRavXWMX2WIeHkjv6j5yLBSqvwq7Zyk+89hMyda2QXL+Im8+CmFTAzi5
nAKAlTmm2GFMj0nGQTyAvjT8pv8BKtyXRXpF0ktwuqwJcSlJg1RjoqGlcftpSBUm
MjpU8LZq4rfNsN7JDk6gzGuR3M6JugiFIvnmeOPu0A1fDe25r21TD5VO4iBQj0c+
aAtjUQ8hefZLbFfkFUkzPCu8igRcdusJ2XqLK8qLeIXKdxp8WtLOjW/xiUKA+mp0
HBTtkRxLqbazXY+xMa0Inl2lA8Xe8dshFYzKHAdCDXuwWZ8ZVFICJox7TWGx218G
Gxd8YzY0PrmN+70nyXIwVKrFuMQ+/wbWV1LTQvY11rH/iSL+7kFhj2qXWag8bqaB
71uNlb4hkIIVfCO9/Ht7sE97/gikKV3YCE31V3w+KBX/s3WabKHTU5KS7M1p/F6q
YprMbCTI5pq8b2eIMEDpFnI8SWwOBQ4DO5ZEdl86W50FpsqOyvCjxJPCbqojiPdJ
VX2UTZJxUtSHJ5/jQwvXZasB/2NTl5vdzV/i7tb8pVCh9XAIWoToqUFeoenQhzHs
3DqlObqhXdP2TVykwk+ktYIcjD2bZqgc8iMChr2yKxwyKVn9kUEnBjXQIB6tpLoi
fK8pFKxqkoZHNNrm+wm0UXtykRdMJfQwymetF0t2gvFFSas2/n+YAEcrvAcvAC6C
w10AIUJjqjzlwqniED8JoOTCQ7s3nDyMWVmPgHiZ3oIibSA70wznRh7jJXDtgH+j
MgGJOtGuSub+lJfMFzL3+zzp7j4Z3h/DyPaCVEZ3DRNmObKNS4kA6i9oEX4N25LS
cXj1A9Vd8uwMJvF7UoLFgWcQmJBHg0oYSyocdqyEtEDrJklURNQSVrcgiSk+zX6c
nf8JX5eUgkBIS6yv7b9a8ejta0O7Pu0LFP85yJPhehZ3Att2eYpPkNohjEMQXflz
1Hf/bOMam0tCwfrFW9wXfiR3+/PJFzE4fwTUDjyIMDp0tR/asJigWW13o2ljNcrg
kuO+CQ2dimIMeRqByqNOk64Z8X5BU82KK/6al4yZ22DnRuUigWyLbp2y88A9ziOr
J/rczRWCqYM4oXYyy7YAwF1LzNqGfGXBI3qhiK4EGJ8wLcVFyjXxrGNYy9BfR+3e
ZwYrdynPXia+lT9ONtHUXkFUPh+j1yfaxCsNyetDctyih19oqPrL4txd+8c4mE50
usWO/+dZS5vlQJ2MwbLu009Qklxwpi91fGO8vy9gxP68KiBRllBUWr5bGd1QUPjt
Zw50ZmHpihJSzep9kqiu4b+WBFTobxRmM4DjpQ2xxYKGRm04TFsfYddIAB3gvN0y
lBp3CDstmRyUGzpql5/J+hIpgKbpCWNaVBgvcWjiuWuaDaTfJLjdjWFLeDX+UR0S
vvy+ty1+R+29+OMwqa4YJm73VEhLf1YS/7znCkEZZPEEH6w63ntTWGYykEjtkiQL
1eDcEZhMpeKqkUt4vmSrZqhU3rDFJUxfxCO5rQ5yJ2UdWwVSeCBtOtUJYHSdKwvR
2yNwlDIpFFLynZ3kPI8hA0XK3gwsUANydAaO6HGpiVMtHapC8tdPz7aM0d1OSJ8/
cfG8qX8a+tT4J+THtoNAVkHJUAx/L2OctO68KMjR0Swjo0ZCBoGHEf/qkAikjU89
AzddK8otr0mh4f0gIbzaGW9YXOof/LfQqj7pvmvU2MRfQ0dYOO5o3StnW1Nl3J8Q
AAq9a+47MeRNu4vXeH6phV7RRpKCEGeiXXRp2BBZBb+vffsGI2ikESQEese+WC/u
KkT4zE2CuYX3tSAxWvnTb4ayyrl/LYCHRkt5b1+5hoXN9dYBmCI6f6GKM7eWu9+4
0J/ZjNgfyxMkXTCcRRwlfsq8m59KTKJikhl8webkOZwoGufTRbQszx6y2KD0+sFY
FtcLylGuvAYvVTnQz2o59vNQQS/CeMDoh1f9Z3KYogTh6U6MFo5wHb/88I8lGkup
wFjQqmDuf15GJ2sCsKT8wz/8RIS0CFWmgSULH6lUgVLUyE03wuY7JD8Uf6bhGuxJ
OvohcxiU6EPbtcb8qFLGmU4ZKka6WvXN0AbMp/lCyVVDntFR0j1PwuQM3VemvJD6
cJWfvctFaPU/lAUXvW0MI5Vr64MVcncOyFSIQgaZq+qZszNEqlxxU1F1Ye9bjLi+
/6hXqzP27M4FiXlWFMqffd3WW8WtjWGub+jHYJT3yO1Ov62zZi8eBa+oYkauKy9v
1sTif+cNCthbf8kqBCiMq0tvXsN19sSGCAqIkV02jMC+7nz6pdG7F8Hf9xejod6G
YNGSWSemyCIRB/dX4GuOCrt81VTuidhg28asKv69z8hJXpf2P96M2ZLCdcbA3fk0
ms+B40YLyASD2nKsaphvhJ16F3O7Y0i/8yROHdkhXtmkbQmdOI3/koCI49QQrXC+
mV1IOqNL4960L5Z7rg9KQRgo5jyJ9/2aMxIdqFjGbyJnokj5koJpJzmfMc7Vybs9
qcO5y5KwyJ6Jx2P2CSXGb74CnDz4nI7eBoTMDds9g/lhV5rJ6BV7jil9Ofh3ekRv
BKknSEUB2U3ZK1DvOlig8/jsfg3DiV9xTnJvZ5VVyxCoGVxPblcKBHVxmDSLWOR7
6OoDUSghJEHJ49n5Snv0XBN1QqTRFfabtYdTYEq5uz0ikxHktkG6jP2D/IVe1LZD
smnwWEbjR/2YTMURjoOvx7nyLwl5PhxddTk/x0b8Bmbq7/ZJnZb8Agb60L1NeHn8
/EKLEoz5uakCyuo7l4ilrnWUfuJLAVnLPARvOCSrZWUBaVwa3xr7psQTBeFs2k+V
XrsvJPNyYtz5ENFFq5WK7txOAW1c12OeTceq+NrxDZvuN1pNwZwMwP3q7yu5zS1J
b+4ZySwFTyUecI6AYmv0R+MsaqmLQJkEkbZ1DC53gAf+HJ6GG0g1kqGSyLvS9h8e
D/z6kb0f7K/eFtbdOJIYPFbgrmfxn1m9xanMKNAJv+p4ijeZELEzGG32HnFOZiBb
inPDEZpYpl7tbbWU8pzx0EQDOvrnZYJxU1fvm8g45omIsDM6wg7UnOilElNTZsCL
Ay6dZVvvlC3NGjuVMdLcGMu2L9wXabfownXYVBwFJKKn2hBGU5Wh+zsgXIqvbqYT
9IvDpB9vOGEFaUc/VjZbbg37ud4KS1BuSCQdAVUrOC0FlIBqnHC9h7Q74+BuDMQp
0lRnE09a1Li0vIgxoMk2I5pht6GlrpQ2NoprU0hZQTcN36K0nVv3zgHpuIh89cd/
sJGDoqjzdg2FkPQgsD2QQxuZE4x+ibyrG3HYLlU48lzNMVifyGdBFk+wFG3ypyTO
XAbPLsxsh+ixErGifLqB34hdmJDqGloAV+pZHNVoo+MS/PljQ6o/TSkkwP17wuNx
c0/Tj5dF7XfB7tjJ05zXfvoDZs9khWUYsdqOB77sx0PNPOu8ZmnDvBnk2n6cBWYr
3CDOXpcQpcsUEEzqw+7/66NFJzl/pLaAT9owfjbUL+YFf6V/EfOo/bANvJbWa6TJ
y0wHX95HsKKsNeBTrcCyTmBBnvC7FB1fYi2B0rikElF6+dGGAfnNkPWckSNdjNA8
UxFRZ2O9PIWdBbpBoL8De13IWdHkKBcRyFYpQn/1enxswBvMChapKzsl+1eTgTEq
g8e5ECxtr7o6XCEZPgufMlKYxy+8OipKCVp+wRfKxBYqEDu7pVc0mxlIW+tTQjfF
lu8H4ZlOk0MZJLWU7LyLfCHQ/rTxyJ0m53wcFEt9epaTRU1fJZx+VDwJzvRBuLdH
x+LuMP1vkb55xzWHdjotrn5RgGHkhYJ+khpfDnB3D6bAapRmt4jStXudSJ1zglZM
gFGLtwET9npErSVE+iYKdA9EOBG32NljVxDZiS7a0GpGuAbZ9RD9z3LmSJ+PrOC+
dW2/Eyy6+xCYpkM4JaBwz7YqgUu+1C7YpjhLBmGtG4FgdHw6rSVItTqW1UWmYZee
Fl3Gi+GSiRj7FvE9AyL2oj1xOUtQn+yUfmgH8zakmJS7dR7HjMH0ldzW8zrJCDph
KtJYGHIplD+lSqJ5I7hYKpGdj6lNUa/pZbS9tyf9XHEqsqz4iCLRN950Nj5h+z39
`protect end_protected