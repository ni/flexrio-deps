<<<<<<< HEAD:flexrio_deps/PkgNiDmaConfig.vhd
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11488 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
gjQxfoUVC1+c91Q8h6upBlWXS3x+ITA9lKmGVxpdDEVLC5pmmikpTd9jQCKFTfWH
oQjHG5qQ6+lmA4r2GwdXHVU1md2u0Mu+olI56A/jW+gd/voZSeAlTN6wtWwE4eHY
FIbFhdt9orARX46RyfQKTbsHsWvWNFTayyYjCedQtL8id2ocmZKD7tD74gg/tW0D
H28Nj1O4LK6TDOwUeiPnN1Ad4TbJsGQsEK9Flh9Co7Hv6nZVRBCGhbO0rJIKJbgd
F4+KlZUlaHoDnmCZlRJizc8eQds4UDMGbzBolqOZEPh/6MxPfdvoaIGVNHvSPqFb
eDsgRphR/rjHRnZPuVIipZiycLwyvAaVQFRnhCxPETuc5PCcALR//W1jH7juYfCQ
EB2KCJdhFdud0J1Lon1rZdCGZKaEjEDJbPV8eVToLkdQiSb3L1YpGaZzeA99Dp1Y
Lu5mnWeC/gpZyxWFB87vO1MhdkbIy9ovZa1DbCmyj3wEAs/M2VjzVKg3Ctt4bzWo
DyYT6DpV+n/kWFWxgZEIZvE8EF73gDhJz9jIa+Zk3IbmPu3kQjTw0XIETHT42E8r
Q7rvWfajRYQISleoUziqlMtWJt4YqWGgkzLtf48Rzlax0u8LuAEzTzXDJwsQO6gu
Cs2AthnDUbtlaTH/jcXMoJ2i+5bNvh/quKW3U6itJasTBdfTOjkQI60AaB6GeNJj
SYEdri0GscHaeGNqbFK+ZdRWQF6er1WkodR0kx+NDOwDQjDhAGY1g4r8kD/U7uZh
RkxNmK83zjI3NZLiPcrFMZFAmgNWSh1Vv9g7YQDyfWSyp30qEzfFgJtKwS3tcW8S
B9n5M/bHXvCGvuKkTpFYdK1EA1w44Zpd+gVbJr+3LQIYmxKvmuwVOJSUrWJyPBP7
VXv15vbAIbZIgL4Vldcft4KEtaukhS8khXM5fdo0RlBBQQMH66eVZiga+jNKTmlt
VR3LTHJrJbH/XHcDpqQpLswwdxnW6ZxpC/YStwbGcaaMP98BfjOkpfBeaPLzCj4c
Nvkm7e8IHf9qgfwI+0wep7FZjvyt/dd5nhWeWZ6bnGBa4fdyRRMGtzKjQv9MU08T
ufcKkRackd5dqfEdiNQOgqlr0LJTnr7F+viKOUag2lEsaeLKd90eyxfe8ntu0q22
IRsExfACID9hyuVBBXc+IaKBDAr4StYXQGbbWAg6afLVF4GR1cUmHJU5vmFlmzDw
dFDSou6WKPAwcxISU9GmHM+g/JQihjAiLWfnnBMJ+wYANxOSc9BcgGK3WQPl23tk
SAqM8JvcTcQSRvtVbuUFnl8Uslf/HE/GyD2jMv8r+ilm+FgxfjVtapeMxz/GrTI5
A08qM6fX7Du7T0IFqiYKfkXl3u9aPo/h85vpHvKUVixReOdGSAzVpoL/ueAvwx1U
m9qHuafuncLbYRY5ErSOr3NaD6FpNVT//dZHcA/JUnCbbelqD9ifiVyA1ZcsHi08
MXzpVDDiKzPmEms7HZ3nfODIvXFht4ww7uNfLFL2vmkAM8pz7aCgUAqmdY2Yzwrb
tsV1QWTzmxt/aBBTIlhkG/MhIvGW/Ee69OKYuutlvf3mrirwF+X3GlBBvc5D4Rso
bNd3VjGzOIt3cifFMD5FR4AQKLnPP9xDACVLmUvFolaBZJ6XbIdm8CvOj5MDMNZU
nJRyiNHwsxRR1U/+HvmgMIQ3cJDU50SQ64yfYXp9vvdBrr5q9CCeBimeeiaJ9GdO
8qy1sUHm7kiKyLfmVx94yORnwpUYs9Sv/2dr5F42zofNvqTgXyBOnY/D1SQzZpar
qy+Ml0xEBfIv8rVKQgz3JmnTu9BwZVLkQsbZ8gr28gu6UkZevQLADBXPMMmmq978
sJWCWTrGzI+9C9bs5aw1brI14vUB7crfwmNCyCnC+zSAnisEvR+Ta9kjAWCdOnrN
Idvhm1s9K56naQBr6MMqIKdx8UlXN6sVL4ywt40dLSp1Q37mgsdsgUAv9QsQJsQl
sTQcYVbppxPudkD3IisndYd0+lQkqhXlIVzyVCVNKXqoveFwYBAJ1qqF5xL1RDbW
ssKSTk3uRu9XkEzAn98GjFc/dIeHn4SWXACZiCZjki0gy+NLX0o28K+dhjY1D8kn
0AFFtEoCVlWZlP+/HvkFfU3m1CcsRH9aPnllk9HV6eM0VWoRVRW+HSL5+xgPxHUa
jZ3Y31B0iC79b79GW3FEtIiBMpSYwAaVh+3N4HcY9+PfarUuCEFo4o7Dh5GFavt1
Q/U5uReESNRJUtkyo5Lyf49bEfGPD6JnOIaJRok7rxuLGVr9xfcdcbWHzmNM/Dfe
pjvDAeT7jEszaJxguoSngOFQN0CDa4F6I33kCe91IHeLR69BXBadq5v7Sij9zHbo
dPEQzPXtik0K7jGyf3P8ayd0BNnUJXpZM1zbJtBTLwFLXGw+guch+lKLmxgk5hVm
Lsb2GjGIqnPmBsmWXhhLMTCN2h1YK5vlDQ7I/aUb+372iqD9qMzf0UMOTNp/p01r
4OQrt+Ilgxlckh/u9HcBUCG/GpB7wOaPWhqUqGgf11sX1090fKAsNQ9zpBphtdYA
r0eFIgVnGAkIwP17VXURLMZh5cKOPuLT/IquRYM7gBPdwxPOOpSE5xqNxA+WUM9z
+Yb0+3HRonH5yf+VjVLUXTQYUtbE9hJFsZq9LgxdYw8cPHtS4FA92UFkjoeEMntt
hr9WmGHb9/D/juWYILq/0v+MFu9K7GWMHNR173NUPk8b4b3lifhLcv1SnSTQEMlQ
q+w3KQp5wXzquJ5ZMyAricOGSphMykLOV815i9Vw3Y/nHfMDMLqCH0fgSObOW5Xh
p6hzX/g6h2x76AaX//svX/8BzgLz1SDFcJDINYeGljSL0Yz4xbmVwPYKOkJO018j
NA4Zq2IUOAuoZSFsY4L7C9QxQ5j7pq6IUOIttPIwfGdfXhHCwcSogH9wZPWBPt4+
EjHaEF9cbvsmk4HaMgAXaXi2Kj2qCojyUBZV6y00ijEZVMA12bfGpBEQ1xKcDLec
IyRwN1IcULsj8BqhbiGDfIcZxGWduOCcSHYjc2mx9/Q0ROdYxqBCd1pr16OjEQPF
EvE9BUEJQVoM0BkhSisc4Af6SOnE5uk+N6U/kWcm5+YBhDvyhgxll43Oiy+Yk41x
Bh8RBzovsc/6sopYUubrL5+JUtLdvaOgFckpAhZCn1r08jNbMVIuEgaGSOc75Qrr
5acEPlpVuJBv/8d5a6IXGVBnjm2/I3dbCLO2suTmN69NUbO66shEY+0stkB3/tTp
CHeYaWvji67PEvlcKGgIRbfSLyR2yJuBFVAzpfBDE8IGIKrS0lXr4KigC6b0stzf
X/UyJh+XjeX18BNQ6xhQi8oX7NAX6jGdEpXftCze5cSLfDaYSFeD/Gcqzi7lbEIx
0L5ETK2BcwMZ0zBD7Bqf+99NInGdtD89c81SQxjnvTYMfSaU1NtN72J1Rk5pR3i3
K8NecSNsQ/4DHcXHInBLGwFW8XyU8AX7GOGD3PoRpur71tLcpGass+W8Wz78wIwV
Hd6pbxpBQ3D4kTgs1ywfSKJlAD2QpsB3+T7LBUORzMu60X+TL992f2ZRzW6YG+hd
XseZnidB3cChWX+xrsA87FIvMkVCbLoRl34+iJqHrLZ5TfoghEYLV3BVwWgvq2D0
bWR3DcMhi402bnMAPzyBI/LJVwdotbCK/B5gR+Gsa8LsbXaK+I2qzcceGWXLT2Id
0KtInDmXiVyOHvsjjWA4JD0WoF86LYiLCeFEJGneOngRP5Sc1CrzEZOebnKi5iNk
1Q1B0aZdJgMQ059jLeihPQ5vWXC+7HXKsfCJddcKmTE8nAWJnejGUcvHiymQV/3z
C9DIHq0p4xhegXIKOsLXbD5e0dHFmNr/UfbYZYbACnPsCv8XoEpoy+xEGdg/Snf/
59eoYcpwYCe+4g25z5GC72I2N4+3ulcxujmLsnUuDLyTw3mLRzMg0NBClL9tYLkw
r+2F9vtK0VnslDQ2lmsnF7i6VSqMCIlhSE4UjpHqZdKQLlXg891N2UOYIJMjrOHg
5zDwVgoS+VkqeafOKvl4O/+I0DbS8KFGJOny07LicZj4P2Z1PtTxg3gfaWjk/KrP
ufHs6HfCFxS7tzCcB/Ucl7NZCu4w8JBqjfzNA10C1IoXB/0SYv3vv8f9RsBxmLpb
0EVQ8/1FbIVCDysqa+i4qadT0G4Ry1wuyjLJ2c2S2/fT5m33v4RwNo0B2HMPIcx4
zv1aErBw2T7Eel4Gk8p976vLTq7gOuAfK/ZhHXYgYFv5Fi8b3jxhTimZLT5FvjiX
ovfqTrneIrGw3MjLgV3+wNfGzdYT8N0RN5NOxQHMy+rwdJq7VL+t8eIhn14NYDEx
k9cGNFRManhcOW4BHTFb/t7kARFKBCe0PRn3U80lr+l+hGZAzs6PFEchvG8eMjoy
JF0G6/0htTFk+0NS+Z/adGEHMXQ7edAtdRCKaiPmGLhFV26jrTnK5Wb5nN9/0aoE
97IVJC8BgVxmJObF6Z0tKVKn5NgLuBPrjK7BEzJfRlClBmiSpuELa0EV/eS5ezn3
bm+ZLr0D4p7c07kJMrpJIk1FD6dludBHOvV2PRxZ4XmxDI79Yby4lm5RrU4ZCJHl
57Bgja2nayVXOkZ40nc6Z2n/jG23/rBp8oEy8p3UzHJMBIbttn1wzzflXeMTEzuQ
xd05xqVe/fdJ4sdqiUmtljgiztOPKVNiYrs4yAQ4H70FTYhTWbBH+hHCUlYvEXZ9
FIJgSUxKTHStH55ld/Z4m0syzJhBOpczI5e0xeMhlTo3AzGexMcVHJ9LC9UAkE8H
YspSgH96ck5f9bYbL93Jrj+es3zs1MpoQ6mBa8awDSGNqiG6DLQHRzIOflJv9TI0
GGZ/G3gblP65nTDDSFL26zz6EBEc2m0mdBFQqmFxE906XqCV9NZWCYz56y1HbBiZ
T1YZaSxW9nmPfCf/C58UcBFsJqcpXhYUgjckRfhWbErMPwHg77VZuzt/HHGdF+ZX
gm3hAp+kruE03JiuycwFQcUIQMsxhkJa9AE/5M6ma43fzKlwYq/eFfgvhF+OyYmX
onWGhvqkx4tGG/TLCMPPKswSsoUXv13CIfTBRT1uR+g+KBX5DdwcvOhk6qi+b0R/
j098oXSDSZckOxQPs/sfyFAc0B7orxK/tnRA1XBUupE+qHgONig6xmvhl6UA+L/v
ysuIeUhkJKv7PFxfG0Wy5OoKEQuLiHMPPya4QEaa2Vy3TKFGqVxzP+H+bPWu/0Xs
ken92CMWdNLyUrZct3uhk7gfXJxnBqDT4fLi1/3ww7qfbf9kRuArg/ClcF42tIgk
gzrlaIg7FZ9PvLkXXCc3hGcJwXedsuyQ5AqEM4ErQ6EuV9K6CrPTmDppsVI2QdiQ
Sm0wKzeyismjHF2cijNnFSL4l1qcbYjFFP/YYb9SRBx9ybHyqG5zkJC+kP3XGerl
azO4/JmfbMGaRaWWu7BYlmcR7SXjyRgcHk3Nl2xmk4ieUWm41LTetDVyh2uKMKe9
CuKGyKOiX7TixUs9Bl66qoEKhBiocria5DH80G+M46noRaRwk0HU5WfoP/pUbAqM
/20rapKNvQmYmOyUbrmg1jFlVVMGEO2ZKcWPoLL5S8HiWTVZfMOF8H0lBdETXWVd
eS6YjfO536vQcXrQ2x/BrQBp9wOEfEybA/8Oxd5DUjwTpbvihPba0hF4QgHx0OSW
u6brq+j3KDzdJ4hRfUJrssG4LxntmjKCVAT+LHdvnpQHNaCHxT2zan/7EWDObjhO
zwfPYkV4h6FQdQVnRKrP1jTdxdB022n1wyJPQ0lFsMqxcb9suvxf9fhC3kQLRtlZ
KffYyq/4BZMRAYL9ckHggdUOdNqxEVy8d1PAwPSPXZVT5DwAzm6jUYuIKVqb9Crw
H2cuTcp080B2hG1F+p6Yt4S9Y/H8qpz8UFoRHk6pNoESj0laCqZAL6CPihH5JI9x
cNCMiq4LhsXhEkwN4pJYongwAFhVuGXBWmJvcBeeb7mRJ62GV4X7wPYCZ9eMrVcQ
aLGv/rjvXCUvWIjfe0F76QZxfdcSu8wypYySLiQP90YJCbaVtuFn7oIGQpKuzNfW
oAw53s+zEGHIPuPW3YCY21T/5xDTlxgcG+Pw5haf3r4MkTxgb16MHwIJ2fFz1IdO
FweldqP1QOPqX0XjspidTJnvT5ObNrLbVS9MLSWTv47aJ6CHLzLlH3IhF6Bblspo
H62SyiBga2n64MjqXBIF3QCCjKw3iVmghavbcXEkgSJleCwCyCt+3Y2TavobNm8p
1g3qQPJLzSSZNDOkT22xG1Aj1o49yeq08K4Eplxz/zbDGoi7m8rt1NpNeS38eODp
k6twpRdEdy0igMMVdHnlW4ronDy37/014Aba+O9eZOyWXz7koRHfv0tz4kq0Ko7E
sF3+8CU8C53etjc48OxlPAx0H3S3v5S8FtmSSV/8WV4T8kx8ygC5KdeoPHmIgvl5
Z0GpguKN3nJpVivByUtrkDeE7+km17meyZwzIZJ9YHUQX36FiOQkxHMDQ3oAWsRa
JsVLmQoZoEypL8/AF9u1NliTs0T5caWF/8LeTp8eAj83ORYCK9TYgJdZOnsK6ACb
4xgoX9VZ/aU7yN4O+6hZcGpGEldoAWxIh0FKJ8GV7ExcjqJkBpOqGHDqFrNIWVyO
kARRTq9Ng0o59KbwyYKvodzQfXrqs+HAAOY3TBOnFrztSwrKtD/Ke6TDi/CgHxpo
XC1TaW40QnxveYoWDdhmKMcSM4z5YjakaWto8K15XBev4b/pXSsXxi0bGeuY4PpD
/FF2xLlfiRQm8u7FLFgFDsa9pVFiI5hESEq7yOqM1AQtqiujgrSfAcUAPncuu52z
4cNoK1MxHFmlTqZrb745N31zS4vRmS7IzvLyX3Rj3VV3ynVCJMSK6dYxHJhHH1Pg
OtKhM74UI0sshedlUa/SSslNmfWK+lYc/WEbA9L9z0obeJJfeGnRYGergJxslVA3
TUazFv4QdkVqPo5vrBQLk4E4D+EfivSGBSreg5AX6JhCk5ZBbQ77bFO0LjbdOqa2
7Pk2iiMV5bza8IaUt2IeJrnnV0cC1X0rCHpiDZQLBkJyxx4rZ9pYiwIvEuU4gAEx
P/EKjdFDzJ8PztyMDVSjNOsbceC2SUtu1351c1YngCFtG+oJ864RuSjePVljEKNm
2zUOpFvM8hJ9fjr9qshRKGzxEZEpyY99t6Owmlzw+Op2glg9b6m5YofCHY7NnDis
dLC/ZxDMjDV2D7KBGC8rOZCKw5xu3VQvXBqhU8AWtSCA9HcRcZAMgwPH5ur4lAK0
JaCKAn4sMOzfwXHLKJoxO6ujUXQXfXlWfe7FnL7TMiSn+rQDbAthkm+QxRDZAE48
Q+bkv+7vxQpmiLSysMKODPp8sZfw2Pt+dPIYoeYCfys+vImUhiLONI5283nk2L1s
jBpWeT8E0hNvdsXzhX/6or/tHldTIv3l5cLHnDpL8jk/Yn4umqA80I5Ykps+tali
/82NZzLlFAS2iTWjXJMB5NkM9oe00H/jfQE1FpVUplB79I6b/yUWTzGw7rsolohs
ZJESxfn7rXMN6k17WZxtjddw/yFuYDhzSXFjPuogxtu7rDifwSUjVmBcDMnYg1xL
o6VoBqBlGbfEdx0+QvQAsShe34IxM4dxbNjO5xmyNJQzIt56XvJBXBiPUisKx4iD
7dXIdoPpxe9Bpm+AwvXAMXXiZ1VEnsbBp5KTMF4VD2ePYe0qFYFDT6RqaDx/7AXm
SBXTveubJwPURV85B+RANlP2xdXuHHa9sI4yLZHiglNuS+ieT88DnUrrtbHWigME
k/6UB1z2ZiYuAEs07+nDzyNbF5koLsdUAf/B8Jyff9QVvUHDnWkx6+D8Izl+ulQt
sfYQZkHnZw3ZYKRVbs92EwfcfdTfgCEBDNxMhxXQjiReriLP8ttme5pFd0VYUHLP
F4fMr7yblpixRiNG1iJKrCg4PB0rLyMPdykFkFTeljN240zm1B3b6fQuE4ABQdIN
SK3ygaqlBRFcNuwTBTzhbgXhrhTSMNAwiTqFQfCluzlAYrAnHBeo9/We/0jwgaKv
/lOP++1D6Pv0GO3lVxY3ex71CvMJtuwXP/0JhJ9WmD0X5hCCT5HghwwJcp0QjuFU
UAVoLlTdUcVff0Okmf3ZdO59yMpa4HuLHhHWAgBCsoFWr14hA745jKjCExnV/zPw
A3dkBptTD6bHCDGgE780++MF4IUCfj6I62l7N34m5glpp9/JOlTZx+M9MJdkzwWM
vmYEuGXN+2SBEydJlcI2EyY7bavNdvr9q6yZmXSzOAWfMs7Tg1npBRX871e/RwF3
ht41H7s8gsq0qUGEks5xb5Ync4CkR6CkVRb90BU+aKSSh+VFiX3RFrdKjEiB4MYR
XpwIAVC+9EQjOGJaQFWrQ78zpGIeInQadi5odOshvGdzWFd9wafO+e6uE6QMKGuH
gOf+iN6ykH7vdOEHfAwHdK4tjkArzX8+dajw5p2SYNsqWEq4DbqemrtW7EWs00EV
xfJfdyZDggtz1fbQlUczzek2U1S6W+dyl4BA6DEiA7jFrFQfMvYF78kSzx/zHLEr
Qo8EfIjSmV5GuQAOw4Fh1h2e3QY1cgDZxZT7z6Ufm6LgitMRxB3dlw7djEVt9x60
RGaUm9GI49Z8XT36DhWMa8fkxWb6+2IU+nazdrVQB4Ne5g9Jb67aD5c8RbbIqDom
dkstkHb4Sa+EcZEhPuCZxp4g8/ddYx/paBs6GBgey/IRLjbaFa+jWTAqNkQqsoQg
6E+fm2Nbd2XmHvVJb0nVZw1m7C1zrErvvPZ3IgByYgJHGFRV5qVViTmj7ws9TLyt
LnjY8rox9AGdXCTskc5uNJL3oIJbIyOyFU4RSITZlP+dyp2vuT2D05/gxlTHA92z
yJ5sEwfrhDfQ0FkwyFLS85yiRJ1fLL617WF90tNkzzRopL/0oRMW3fBjOMmNDz32
1yqJOe2GXiVZo2Dl7YyrbNhgqjBn0AkSjDmwe23iHbW7B3ZAh54WOJuB4YXfLEKP
mAjFaaRc9HVzSDPALLLOJwd2Y8bm9NsPBG7+sL4xVLMZ2xrYSYw+9N1PqBX0waGx
Ek7F6OePh9LKDBRf1ZSOAprfxPYn5kHdsfj/ENzYpIsikAuzugk951lps3zhw5hz
+GcrUIuzg2DbnIbap0JecVD+o8gu4NyJ9rRDOdRLO8XCPzjn+67+4txWvtEp5R/k
9Gy3tHnQ/n448YfR16qAFm8wXU5gcW/sdEPjRMpiyB/fE9+SG0qYQxwL/YoZi+rI
RzmcZB4c0sXDEagBhdpS77O4IX1pCt9A0GcTyLe+tgmivZK1lPNVipVXl1nukrdg
9qUwNGdx/BYm20uF/lxud40Mn7U/yrpjiuMDkSHBH/3pBSU8UbhL0Aq/5I8rNW22
fhk2QJrFFyEnD+x9i0jiisXE9K1O5e1LVSJjDcpTiEllvKillBK0JWw0GjRTaUyI
b1Gow2y2bM0ve+h19Qg7F98A/KdcJ0pNvrOTedo0Ue4sI7IAILUWigj5OMjyGZB0
AluCuF81/n4PvOBAhhYcy67U1AsSAhWjBtDThAMGy+Iq9sJDa+EpvSPfhwcuqB/B
bEmZvTkn/Bwe+LqX0sEKAa/gN6z1dVAbtScWv9jPIusV0k4ni3Ydu6ViDdaKvvp7
IEybQ15652zWRIOc0l/R1RjbKmkQ6oF26YIFMPfGS0rQramWhcAvq073HgRxSYfp
MZ1QgvGyLdgEGnMPP2PoSopKjwKbCnhjvuHw7BtG9HoF7mdWcE9lhvtmZN4F79jL
9Nk71ma5Sx+o3VyfBskZHjy8/uTYKYWyY5mCRR6v0wAgl3jYIq1TK6ERlYsvpMzQ
dopzLojFx40fzutTqAyG+GYDlaA2XuJTY1ODH2edXJdQskvM0geLp/GPQt2DFnor
QR/vAcptUo20M0LMRONSQawqDzBKX1q3ZlFf6s7NQ48yTWI9muPIxygnhze1CY/Z
YMRbcKnG5NZe9P43ZfuNTGJIDANfYs541FGndMSpXn1dUj4XOEfTn/XqCKohEWdt
R7qb4UWj28+glaYmb8MAA/EVRER7trUhFWsvAa96qEC1msmUUMYYIJMYclI/29Sg
gL1nWBEuvYVPy6GKXSPy7cXU0tB8TiHvhJq1Tl5KG8oVRQy+a7PDwRiadyV5fCPp
q6EzCWvIbmZIWVgiay1f5BtTNYDh38Y2qmKJqb5F/3sImlf2znq6QWfesGqr0S6r
ClEcj9SC1C6Sgps9eEmEj9ODvR49bveVTGLwr66LwTDCZ0gvXijIa3kxX4jziTqH
njUr+IPYnDu6F5tskeCZ6znpFEAV18VRRbBDO2O7p4i/5DVa6II9eNUUM0rWuCQ/
ila1OLaOF3aCj3uaRw70yqWBZreNPvJ1APBIhPBHkQ8J5Mi8+YmCym93Br8jZRVl
qI2MWgf6X1+GjryBN7YXz9w7C48EA3Dn3XaD3cjJLUN9R+zEENpU4hc5ze6iceOx
ExJgMbZoe6BChykdVYTMEtIrcjcPktTkmajKJVj0O6Iq++NT9Kjkp8kkulbIqQ28
Qf+Qy+R/kEXbSPEAtwKQ+HHEtOzi0MiEHdCQO/cFCNuIZW7QLktUXIHova9o/Mp8
MGJRL5l9Oj24EdbWpUMxIHddrNADHzaR+dONR9TioN18qEHfRr1vlTUyUjUBG8h2
RzOc6iXaWg66Ood8YwvQ3Tzb7T2k6/WeQ5o9csaCIvPG0DfkOXT29EiBvmWp68aQ
7ohJZWvbhWnrrWzDKgjoAmX8f1UKomNA0L4TyslpS/t2PDjypEkmMxUFYhGsvMyw
YDyyhY6OcgCxNpd0n4qLTsUSQ2BJMGADh+KN2av20S/dyQ2p5wPGRGttD3UytfFt
LoCXHhS1aHubBmCNwbNyzFEo8kbC5KqJN3tc0RgP2jrhHygqTjQzbSdlt54w1ajn
S9IWjnmatc/hGi1ImHxADi2X8GPI9MjOfrQf3b1HQxFpJeZrOxqj7Xi87ws9MqAN
kEKCS+R7Y0634tqyIc5J1rv62UYJ4hyYOsnKo1qDvMyyKeMNZs5sdVgayiCaSZbc
PoSkSFRI7AaNAjRDxd3GWm6a/PDuXrv5AHJzeBR/Q7Im5UqVKedUi7+TBibTaXzA
DepoHJmwD+5kcl7KEfZ0SdO4g6FvtCn8uyNG4sAquDDRAAgRXyQS+z9Pnysqiqbu
vp07MjwaS/aLfpkU4/IHi82F7U4CBMTad6+z4r8v56BvOt+9ynGmElOUwK5jBKQc
U+hDLMSdIUUIQbA/R0qJZam/e25ofE5tI/aAn9/HvWswkHPC8yfjAim16jyTERdQ
GQ78TNaHfuQ3anurKGsPRd84aPQswoDIVakL4dVSuRtcB+x8ucjXEKS9oAz/W9KQ
gGyrKvW6C8LfmvO0KUve17mYVwKlkDcZqX1ltC/WmmsJNisisGnscrknwfYnbWQB
eqQNJu9iBxZx4evYaNY+a+a4SY/NWNUbnHPDue5kNfrupyWknKRSNqcRndZ8G6Ti
uXrZL1hweXuxXTNpKdDGjJi9HFwErAMnSRC9OFDFohwCD0k5oc10Lt74uiXNKG9+
2tO0sXJg9tn8NoWy6UVv9qUQXm9iBfOlZ3GtXVqK6Y/ucaEZprgKygs7Hp2NQlEh
zqnUdeOZDAlM/G8xDniTfzxT0lKye5DboGnS8wNify88wQM/r+5o/PMkUZnrcUGL
KB0m2k31Nc08Ykr65MhCPzPOmSThvNmwff/56saMQgjV376FhFSz4JuhesVvXuZ1
xAhvQXF2TKzQJnNfqn4v5197HCfg4V70nnN7l6UteXMcUpyUL53wqQfZy75HpHTp
ffMtr+9hhyLVs7xMBY7f7SvKrhRwuZkVXpsVvHQwFIEfJMHNftYZTByeo2BGe/ke
aC6EFO7mmvie4ntPHW5dzJm5kRRNUclX89umaGsKcDt6aKykAsnRH+ArZACPGPfL
5J4uYHaF65e3ctnjijGUaUjSH1UJOGwnbcIpc2Vo0pgFHD4twSl/DjpvO5HfzyhW
eTbqFWILPD1+MGhkX68pPwZluLCm93fv6cIo3LIICAOisfzUvwR1wDUhtPFWrDXo
Ej6cV2/l8YiMsY5EuNfu0MryCJDQN6nNF3SW4AY8jJgPBmYrjoTxF/cJOmEXFaUK
XihZjGNqm0UxbzVKkGxHoxpG6mtxPbJ52F5nTb//zwWhd+Ww4YDqAaEFjsWjjunx
UBXClNPmtTpzokgTuBEj33LNAgR8YPY/VcImHqHOTuLFGSByFQdzH4Rz6CDVUV8m
48UjilxTnV4Xqrivsobehne43hQm8bfJWAKYNRLekcF9X0/9DiUVOeiQxyQXIFqK
lxMtMje614RyvgQ63814NpanKG8sUe+m0nnC5W1Cp/40cuFjP6dYMo5kEjWsnTbV
2Q6mpg99KPiXIMmvcxeyfn18WD46MiQreP+aApM3MDjAg1gujka5sGJYvery8vAH
WCa+ZoKf/IYLGeLLV2bw230MdmyOJ8lvXjs5Arfzqwh/PuevQHTHxCmH36ylgsCT
GKfAGSlMSQxhmiuZ6HvS2e1ivLlFQbPOgtaWg2ZJN2bKsnTrBmShHBH2a8uWiMqN
U3Xbrk/UJMqk7p2c/nop5q4rRTUp4vlx5579gDe9d5AEz/taR5a8oy+kvEhXMucH
WW8gNNqB4PBf5KGCInYhYcjmedOb+R8NzMzx3dgYR91rqrjDVyatp7z8uzn82cNX
xXt8hJ1bOenjVF65nc2WKdkkn5/vwQYwTHYAN+VHLH8sBwUrPhLjiCVpyqcRHZyO
VYPFtu51CpsK7M4Fg82NxMyFVHFUuGsGOIDyVH1nMLEqIviRN7vaDpf7AOu9J0B9
V7T09ZzlH40lxjSKFsgdKEQGsDJ5HNMB0FUgdSaFDnU2uDfIbw64oA9O4VM/kXdl
qGK9D500hZX8kA/IvQ/gN4HSykCos0JnlYgL82Rya2SVFy/O/n+gMcZw+ze9agW6
2FL8R5SW+LOe/5Rmu/Rq9fCX8C61/KZnRUP8Hc5rOE4UpTfU975j3hMGkVRgoW22
3JxIT8TPEEn1rz1mgnc9w1sM8RBG87wb/rwyyKqkY3GDUfSBw5OGcRvtBir/fEAO
M5EYjQ6CygdMYFhjqG5KLzXjYxZb+RSUrRn8/yXz4eVVk4McbU4U9ixnjaB3RxnX
94sCXcJqxXR7INxJfg3GBwR6Re8B6rrOByMzC21ADZ/8ZgiqhtONQEgHjyCwbO3Z
KB72sB+KiLCvWN0DyUPPRKvTt3MX948JJfbyYmNy2h7F1pXHaH5LbynaiuhSit8m
RgCGLCYLpFrMEExAbl9TxBW8adDp25x7qbf5kAaVWnnLdR05g6GVUhB1l3sFVrLM
QjB91acNpzmMr8zd/EKzrazy2reBvXQSRH7ZKUCunYX0Ao7eX0ygemb6jxPMGjJT
bV9Cld4gMrCd7ZufWDwUw7tKK585qVuJg8I0H/7hN6lX7YfnjoQgZjIFnyfPlfdz
tqW1e0mUbPFLmT5SIdiqM4QOuknn6M6Y/7RoXDvUCwrY+K0tnmXg7CqEL5/u9v+5
mu78tIJZKLsWJ3uytZbAwl1Y8KPt3kkuOoqQBYf/ubpWrW2x9Je6G3CFWrLbFM7Q
wzxKIsUmOH1piy38N2+lTC1I/aUW991G8ZQOMn1XFbDCKMrsMZo31By+5/va/uyf
jG1knu7vQyDPgX0OfGxV7KK8k9S1Wyfde5bH9N2zEE9aah29nz9fDYRZJAfPLGq7
Ctj0Cm10FdRKONP+5r9tJxLXka8LML30TYBoNmE5DhNA00gmir51k2wAHCS8d0Mr
sV4AST37X+TyMGESx9mwyfgoKgWAI+ugAyp3jVvz63Thf3wLhzktffNT8Y/oR9B/
Lta3IwFFw7FDH6V9MCJjXNV4z7jM6XDsFXuRQNlEc1GgqGPx3Uwb6vPlfaOJcpy7
scCMk9tie/Fwv0lrze2ANx1quJBbaL/Hp0UZu2A8ehx1tOIgCzOudU6wuyM1F3J1
q5Wh49Am/Ibt1ElJ28NRYKzs3BelpH6EXBX2+syE8T8c+IAXo9OSSh5NifvpMb5S
gpXxwTN7qFl9o0DapaqfvJ8WEF/8jScClBPm1lNTcwWiYmacRSocAQ7jZ4PXcnBK
ZTtIXkLUHRKEKYP4Ro95+PpMUgocUCc2FMqmTq7onpVMQuqBKJxzNOBruPN2Ia0R
nlfj0yPDgWW0ktbZxX7wNg8Yv4jlUxYajUO+D6nBe6dV+jqmG3fTuEhfqCH+tNPO
5fTjITy4oHx9qyhBV7ov3IVtS/6V3XNuwG6w+/hnZHH0UBmwCyMMJJz4+3BcnNML
DUXOEEkBkNks7DRJxhj1CDO+biAugtn9c1jDovfm9L1y3k6j0HmZx/uM1npxMP2l
4PVeFy8Dc0GqWRLICNO1WXqaIPR9EPpW6wCuga1MnmrpcxgCPZ0qNBGJewK5+Lhc
WuFCsPOlkBFrR5QlcMcop+2Qhg7+yJSXbfNtRteQY/aYS3AYVfPEyyRx8omysJdE
kUN2NteLaZiMjhMvk5idtOFFVfMXZr2ywAPwl03Pa2TTXi2tj3ZXIc8NCmRoRHsH
RGAKIavHh+tRGHEzcTgFELaf3TrK25XzGNisog+9HMyse/uaJWsso9bz4t4LvTMw
aiUZWFxb1VuR5COcAcz4cSfIajvOIigUQ4oXb4xXnjLfhAZvjAbpHE32HpUrtX1y
thM4tBqSG86o7Nt2pqH7uLNKfv8W56JD1rhX6rTuw3wFecEmoQYgHGeHn7sD0K4v
bwpU29qql7/yGp4jnI3n7JREtbW1WoXOE2kJZXg90dj7YrfhqlsrGL+HfSP5Fbma
+cbUYpO/Jc8qhWkW7uWQzm+vcm/j+LGXRwWavQWeQ/nC0ckw7+pvyJcXQgVlbV/z
+zLalHtgNYwYEXksSkNfARYpXX15thct6qL58aL8x8uc/qh7olRRRS3bC+qH8VZf
yoG7KhtBUHJHx4Y3/AVofxYg7Nl/WDC0A/9bfNWnZRg/nxValou7vIVN51JT2luX
ndGUPHej48z3C5htuSNplAIc+KXtCRFMIIljMHt6uG0ze2T4i0T/UeFBzj0GQuNL
duRgjZWtBQXsBLjrDa1rG0KxZ3PiFPfnnrBN6oXlOyRdKQ1CpsFMRGgtxP7xoESs
9OhB5JxvkrGqnPOiWsCIpQ==
=======
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11488 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
DyUmSSJKy9uR92lovAin2mUFTEE5dUNHM4ZRttnZt3FBywxZK5A0V73xSonUxiGg
NFFl7sHYrwRQ7TyGPFUKYk1vqTK7Dpke/d1gvxx3ARzUziY3r3/5iSN0KzkwK+z1
bIG4VvU5H7ADjUEra9BFBVtGNpZuv06HI38fEGC0jZV11twp5CBRBJJl2MPYMqb7
TsI++HaACM/DzxK9duyzlB3tlS4fAdzaVePvsWibyC6IqPAPFFHFh0BN5gWWSvUl
zMSNOl/dYzXSwpi/dF+5TWFbCTzzvoR/0KFSvYGbzyULfwOU1KFnn6GK0J6nuW3q
qMjLiYQbk16Yd4L+RG7PinLcEZP3TANOAXaiJngvLnBkIYMohkeRTa+WnYBO+1TV
Q7Xp2y8t0g8Y+6tO+SNLwhKSccbl2ocK10e3P9rjUCmTVZ/pnozrWdGx6JQP/SeA
LNmwwQfAjED6Uhs8IxNKhmtlxhNgxiwf+qsZcGT3Ru0YNE/PpUV7ettSOnEbuYwf
Q18v7LbmLmBQVezse514Q++8rvRG0TtiBq++m6CcdO25dUA+bu7e6Sat0iufrERN
Jb2OITrJIOZihsnxhMSWgmQB3Dk6G+qPLPQpfxOGsPL2/lZXQBrjhpsuVKxbSuTS
8+SWCwhXXLZhWtSIwdjg/hvbOz+D8FiT5bjceEWVrQrUcJ05frazznapgqpfyrS/
dNQVD2Wv8XxXX4FKfSchMTM217nrG7AEq4SqDKOQ3/n/gP5BSr0CfoUkRrssdxTm
z+s3m7g8IH5GCqH39LGwqSnSQK1cbh5nN43bYVUJ9rzGs0stXDxWOigJd/nzOMqW
3MsGM0k/ZALfzCL2OiPOn9R0M68L+xOnp/aJobCLddeAcUr0OGztS+Jj5NRVmEVC
ADgjL4C+z0XhPA1lHIZnyCTWi1R5eTnrQCa/vqAUjXLZBXFSNEoFa68DRFBln1Nh
OgTzh7yaA8P5jslZqeT7GjKgjNPduGr0xlPdJmmq6T9TUkbdW5erFWfWxhsGTf/4
Uvf/dzLsboBQM5DPKXN4iv4xBLBiMa4wa4gMpJumShbfKi4FPJf271TwcyS+RjZi
STneIt4ToWLE0Q/5Uil0Gnz9BuwMK0Z7py1xC62erWhPb6Z6lmzrl2ruLz80Gcm/
tXe40nkATEWifXjrn8sittVdxjMsDSssDq30ioc/jezJtn2hvYCf1Aa7IuBPKnRm
BNbjyEsmAISTy5hkUlXAEw1ypXjT7W0c8CMGd30UW3w6Wiv3sbVK/PBxalhOyOy1
ROCCzBaoLxN0nhzo2BHi/sH9zfHwFCIGFqmk/W30006MPndHVhhWVWxLQ7h2I8D7
RoXRVb4SeTyO+mSdJND73GtMZxo/JgRNxrJ46oxwYqmu9sOS1PwlQc/eG7YJpZ4Y
/lKEtZfUL3BpY4id20tnWkRUulF3LSC2GdcJ0uXTJrCefFrIvNCiytdjCLd6OGpC
BeQFE9Vny3VHVtMaMHacawuWOVUx8BaTeVLJ7qsRGSnS9Msi7/StUA9CBb+a/79w
8CluD0Awf4wsBtzt+/z3s9O6rRakVwgIjKYT2+kkWljetBzf/9Xp1496/YXMIa78
3/3j6jMPkR8AbLf+5P262wTadAA1Dz2meua9cTC2FSM9qaP9aNNInKki+TwbyN68
xtGUcUTrgG5cKYa5m7JauEV4t4X09QQgiCoWgkBLDgnwyX0LH7DcI6S/n+VoSSz3
GunzjZip+02Jy7MBvPM4pNQ6Hch1NItZh4mF0HHYzrf5UmtOCKUcjoXP05cY7nyZ
0O6arUZJkGaAS1wZEAY0bIL4tlxaiCnPrsxhoceWjGoUVjPdBWrBYa/WClusNOBz
HRDr7k8RMTAbh7j0F5ndPOEUXOlKp3M01FeSfivNxY2i2XnYsjK1xWezdtjtk6QW
gH8yOK9Cpm2iaUjj6YH8M4pe37RAcMIygSHkfzhyUMfAgiVqg94UPNUtclF17n0H
QoZht5JOLDHCaWpdpFitIVtvF0KvH33SC/wmlxIJkl2FU6lJqLwyeVkDUOH6/fHu
6oy/hlv0ZzmHb2/YYb0MHvXuSCTPCk+UYZhlr9WYFTbfw+M9IUDSEKRwB7Y/AsQD
SJmLEBmDhIlMexIXoIu/fLf/DG+ZrYiGdhNLuSuT4qGVJzDLN6ST99L8kPtrtz33
3XBFjpMLrwj7QBigoK6tBhI+f7mrHgs+MNyUVQ6oMy0AIjC9rtnk5ZaA64FjzqeW
SM0PXPcSbRWGVxUREsMnuTFrjMMTvADOi+OBFrlJSlLkar1NaFUTBkumjSl2pWDt
fb+kKTVFBtar6bzHXjYu8+Kk1OUEyOlVJ7ZGb3VspG00E1SZK3TGKgMm/BzYDEUh
qPhfvGC5jc6bGUir5UCJ4qnXozFBYTmOtZdkarEHJVJYyfRbN0o77wFWZPG95wt3
WXLkfubOjhHQMS/Ka0F6TmbQWjkjI+IoBjyuOTTZx5S19xCxqYZiqo2xLBsJIppT
+4H/ugj6rrjAtlEJxzOhE7OkM9uUosXh6S4jVuIUSjW7AOHvieMcJtGBS9bJ5AGV
QxVUSKDOuZDhRU3jibeSnNxmRJ4stJM/mip9ZiKxUEndzA2FNmcJWsabELl+6Z5U
sRXPZf/Fwr+ULzx0wo4hf5cJdH4G6QtpEsOjObzoU33LPc7ECQRk/nz0jOa4pTQB
Vdn+eYo6GmhWjC9VFmSqHMrYkEy+hP1CS8ONDXj+VtLfRJicgAb3nYxzJlvqZXu5
KsouJyIhtrmnyHE/MeJ3BQep30JBeFwsrBlnRjJCdidbcv3KdUmBMub8BXBMfaFL
smpUU9JOSOS96ycaJ+AgfzUbKrKxn+oQgt+7GNK7/CI2sAaw+Tvt/cgpQnkQZGST
3x0F0jyc8TJ2VwXPBmjVkqqZJmLJAY5QtmrIaFQDFdmSfdfh4pN6RPafce2qj/4i
v0O+rPhhP9zQz+k89jSLSeSGahQsTvgXe/W0V/DCVZLDdCngI6LYNM+EVkNy5Ra0
oKoLc0B9cm6pdAROzNpBMgtCjwoLcOf3HnkKm3o5HK8ooky8reprwI/4tlnwwJt1
1Ey5ZLrgAPWORLxSUKFBMaA9QveznPLjwdBrqxIJfKgFINLkoMNMCFq7yHmLiB5h
YA1vH6FTcUOuT1+Vg3Lh624gaMWbEWVFczZbtn0S7aA+MduZYDtJIoM/LVVsNYT+
pFIt2StyQoxGZq6YURkbnDMcGBf8y2lKZdqYEs6OXgbWKCR6SeZTb+B0TehkJv2k
+PRFc1fIjoVKzzeDtefaoAeNv5/6TvAD2E53PsyR0L7UYAS3cY++IiROHCbnvt8q
bpXfVLDvN5I+sE3BEOGt8SqursK3D3Qf53PPWYlgJXxFQ8UgluJtSXMFbiMMFW6a
9xW8lLN8Z8M03srTY0CuuhuC2TL1O6ciRttgLtM9gLVdkUh3SQeQR3rC7yrAaTdE
dGZ+9bYfGfX3SIMxdcfNpfF30SekHnZzv1QWGh8WYUQ9kHavzv8EovK1+eqKlwgo
gg8FfDGGcvorQMjPR+CVjC+ALLXVB8AVTCSD71EAktV1UBdR2CPbgvMi3t44IYho
VHxEMwe3Y7GUHUOEWlyb1VbzR15pXV6q/JX2DaaY1ln9qg/zykZHBdpaPQ3BWEqH
OIV2ehCTcs/vNE5Cp4T+EHjMM7+Z48aX8rLBqTtOX8nWcfEl82aYpJLuzKKYxf08
sdukRulYkLuZeWO/pIVlPLF23lfS/YwXBpKfkxOBF0R4Txm8Kt5TMkAC3jVhx4My
FuuQWkfixt7Ii7pjRRjaUEfM4j+k8jGaVe0gD583zgv3wf1h8+Q6KYNk4fYHUXWF
YgwcQF9E+QDFv/VP1RvB0PZitVsSy9Q83fphz11Iu05rzRawq0fKprhUViFJptpm
5tYcTC7XMvqR+hQKg5R/8CDGEAgTshFTDHVrPSOH9rA2XXhgTq3GNxVCM44qG/CK
Fc6son0KAKTYaYbytirN9F4d0yuJoPlFt+0Ga8vOrTx6ofJTDkFOf4Hi8lu4O+Zw
Uh1IU9Qe3gus6AhZsERlztcZt2O8VvKq+O8Jmk7N+mX6vZP42eAZ+4mJB5ssPpyX
ZTQsRKsJXpTZ70ztFzXewQbWB/RJ5grYOeGvG+99HFPaau8iLHs2VGjNjS63TXh3
OkaaxM0whZjqRUH3lKp+mfS39yfo6AyLdX3FHeEuDi9Baem/V5zSLns1VSyhdgqc
AGfrN2cvQUOA7GxHPSSALus/V9Do3HeGtSznKpzQEoIjg41Tcenkj4VgVNgkStKy
MicN/vFV/SsQ5Locx8Hvi3V0m9CwCqAUP6wHAOmlRec3aRFNuGmjeffUtQ7FaNBl
hYPAFey0cp8ZtFa/cXhWhC7bOAvapJ8u6Xw1gk6rkiDdtEE8WI537piYrOG0WLe7
GdFttmi0PtthodLHFq4mzTAGIhcMHTpYcYIonsyutxFdT3xuhh9f/B4vgt2rXD3u
iELOZLbEwVn27uFs9tulJ82C8nyNUD/Qz62q8lyJemmlExmejMxFxHMwOSYcjvkS
ZeE7vV9C3tu1eJtHQLoZPZ7iomDIYbqbS7XdGARn+LsS63YbTE/iElXDoN3BRmVZ
WIoBwhkYywtO2j50f8uAbkdv4qby2A+StVW7LbjgNuNx49PUJp/XmyxtEU0qgvmM
va276VsQMMp6dphDyciHHiTkdANTKedNQscRqrBWkacmy2zUqlopLW8H/auU/9Cv
40nsxKG8hSIyYwCktQWq+a4dJKkYqgvEBw6vBPSvnr2ch6HubA9GT1p2r7gLyG+d
v9kvZe4LO1EguulGI3myLENVVyavilQakSWLzX9R0qdVDQGbQULUAxSnd8RJRgDX
0n9uYtt7X/dEz6hVohGhSCsTHlxH65aPZ7DHvr1GNALlfXkzMWIU16bz1/qKIG6u
rB2NFAvP1b0lhFI0R81QqLi0J1nfeVbKx/r3n1cTjNQG7sNg0PTQFPUwLLj20856
MP5QMlX8p/zO6PJ8wR9aPU4roI7vvdzU8jaro3X4lU8AMUm6iX1o3AZ8+aVxq3FN
U8Cnq0IAgkeQuoMBWEsxsd/6SON4YxB+N1yY7idzXEm0n9asDAMmOM1aoHs7m2rL
E2HOlhS72xjQyrhHFjCx+VyGk6MIvMOTS1WSd+fZVBbZ2vc3LX0R6IppGdCt/9lu
Lasx1JTOi0PC87BkHSYN2Cjq5hD4xcm/rcRc314eU9cb+ocfXh3/8kXknf455NOx
NQWUG7jbxNUs4Wcuy0CJ3zFETg+2vEZ1WSPvoQPb19r5qvWXyBghPjtF6Jc13hQj
YMnvDnJ4DxTB/A6sQlGkqRSihvXdR3ZgAss3bHKJk172yJr9a7uchHhuwd0Lh3IZ
f9vySZn/k+Ahnh7zzb7on6AnVnwFG4EB6uq6R+d8og6y46YIyPfhNOOpsu7b6rO6
OKWNIXZNFiGpiOZe1oN+pjAs40n7Zu9bkvAkq6+aYAbJyVWB0DPYPNyeKFM53k8M
gYJSWnnQpLc3/rKt09ESCp4e/3r9oiAV0T9cHbOpjwCw4gIUkTFFvlLyXvkDYMt5
F1Y3aSH3UZuhk6Z/4s83GHYzBguMWJKiuOFmIYuwnFHGcAapsRBW7gEEmz0N27U9
iffRcmnmXRWw+P4wspD0gT+KJ+k5oTF18v60JEduaJzdgFEhrqSiwg+rJ/zlXAhK
/zU09TVvkgIYCUYkIQBdnebuHUJhHFs8clXHqa9BEYEyEemW8WGltOdw5isJbTrO
3K1mFUAivUrKhrxrUe/3+rtCjE8RhgfVHYqc1+Yk9Yxy3YyUx1pncue5jGm9za1I
PzsfApioCwO/9lIjue1h0nJM+3icZpg/UrH9nGrw5Cz6CNQsu1OLb5Bkush1VDl7
zjM5aol0WMy0v/r76l9L5TEmibu2WZqshTz4lPqkIRvqSxUcwtcpBKDKf+C9pKE/
t8M9NZ5cBlK7Lohg352urXOnshhZLtr/qVQq575RYiRPutM+1DQWcseYM8RFoj3B
ZJQrUY9PmcYsazQ3PmQJls8ZZHv93pj9MOxxhHzltMtv23YX0Fex76SPxKgjiqnj
pXzC3GOseuk5EA/M4NOmoXY+Lldz5ODNSLmHdf1tV8paq5YOU0sVBkZ0JvL1JERL
HKC5W9Iyvv6NSoZZgeIUsLn/JBejktLYZChq6Qk+sB4nIZVBVil4RrJJAMjBWuY9
fkhBBUFwmhauakJKRnPDZYy8NFxGlPaIiDZhSIno5i9Yk4165Yfkh5nPFqy/5ATw
zIwG7AVb3/wmw10DYyoOQydvlJkg13AWUvtuKTMotPEZsqNp/crek2DaL275lPP+
kfx4DCZdB+n2w7MB93o7j6I63/IJgz45+t/3vLCKr+n5oC7/o+PNrRjB7D8D9zsu
z4pbf02hGWLW/GYE0lF4mRQTSUVZpwawNnHjwx6BpGa6FF/ovstA83hfJ+lu/Y5v
OAJ2sYrhPbk3LUzcwvrK+A1/eVzD7W6RwP3MjgQRQ2wHVApzI0A9QvE/4JXb9xrR
UcxjhU39VVAp6DhP+C6cuur0A6tc1dHwEGKT/5LSUHSeP0kt/Vsyuz0y5A3weXfH
Inppvj5ZjqmNUoiLRn56kd8p1d+AXNO70qM2c1fiCDQgNy+N/atVUug+pmXuQWmk
7rMTTUpaLYOssHseIghpXhz3Wh2p61wEyRqY++/Mx5oN4EVJvYYePVLZQJT4zouK
GOqDDh+gBTe3IgeVtKnTHKkBmaCHhxgXb+uCj74hqivnUcIt8VmJStAJDEfwCyHE
zqkaEIhvmvacEP3Qc33a6GBVhaF6AgQ9WSG7f6fLPH8W5VxTsnUw4cLXwgvUyO0K
GMEXKTX0aM1Le8yZwsoQNTddwuvzL20CrASAr1FFmvGtX4N57/4oOU44FacyuabU
TvHDlsLIAXP9aUXyaHBcfImTmINrWFtpdAEHi1J1IKpJ7TQFA4CQXfWnD8EdycgH
5VZcureoKyRdzCMTS+1975ivpRjI7IKtsvnDM8G1Brx8/4bHPlE1giM01fBxe3Lx
vr7+79iHEKekJ5LaCn8pprPlk3ImLykCLgIy25IaMpMo22T3ykK7zPv3J58MEGxS
qmvcQIp1MwFJnTBneLmwcWQJCDvGnnxyq2wUrv1JVwvhIiJHGxMjnWmER8ellgM4
5TT2wB52Bk7i99lm/qcSRnMPiFASBYpdgnl5Z480N5fniaRm9UH79NctMfm3la4i
q5IYP2LdtZTdBzbTVp9rS6hyoMeeJ/B+A8BvL11Pcjtou+oOmrsPkBRGscHaE9bL
QHlUcTHpo3Uq8SK9VYVRTf4ZCcxHcFLWV/XLai0HWh0VSwnjHiQ/ZUWloMbspr71
UMzlQVpqPdBsKrnzsFeyqB7h8Q6VsJJ8tIB5ck6XMBvRPDdb2xKazlFPjMeJsU41
u82WnPSE2iNlPwUchHfLTQG/4FvVCwRWNXA/+0dbIL+AYVzVGeKTFcLwuYWL0XkN
mfeGVoE/eS51GMHwgiwI7XutS4DcKwKjY3fskk3nKZR0hJ4i6z64OKtznqBp/2NB
s2AyOtTednwtA9bWTVOaVl9+0u2mQXQMGB8wP+wWknJ4dX9A1SAFETPaTrZcRFzS
yjCCtubi8w+PLvZhG1hU3y5HLCJlxl4tJpa5JN5HBe3YH+Z1/31c460XhRefZn3I
OcOO+KCk/wwm2Scea357kO7EFPd5eP5rRRAEeNy36juSGgEKUsIabkGr9xS050iX
nyhBcmCPRWykhnpSsxnplnRO7YLQM/4QR50868rag/Cs85/+tQa1t4CxwE76ezpn
m9Jh02QBcCriKfSn0vKNiYxnxamohILD8mYU++GdpdWMMdNOH783jozFUngVM11Q
+reMpc1dlfCnUq8pM9mBBywQHUHbzMe37oobKLFePSf851fPArtOYRBdHVtUnoOQ
mzL/uUZJ7gAmFJAVTjKzKwqRlnFBHkGk48M8UJmoaFuC7ahHFnE5Z4IPIiUKJOQV
2erEpM3gFDDdWHtNhD2AaOv7IlPRX17kpeWZ0XrrezCtcRjAMrcXCN78bFwzNklW
JTBMclYxRdWBidTQO9mEq8Xu8L5dVMHSKM9eX8QxPify2UNFpTBKa1MPsG+iX+Hc
+MzenuyEmX8xmyVfNRZ8z8QspXClsmstucIQDP0ggQ92y4Nb0Ly8pjTt+mF9cbPK
pHCcXqgqNqGjI2Fiuj6rgd36qwydpVWc5mX81q8S0sHk0TDaoNhtlnShfEtNdAoC
4Pk/63CvG4sQYrGxFx/qI+Zow7KXRe/mY/N0jLxsTV9CGg4MCxwwLyKdaH/gYntn
uf0RydjsHTCAHWB6OabfTj1Ng5JjRk8/hhEwdXuZUN1VnA/tzP5dksPN0ILm7Ret
MWYeryWu86E5KOrvtAH7MF41OR8UkB2z3aCuNwMTqWT/XLMTFD7vqwxRzINKzgmD
t27XbUtmfFb4tyXVqkLm79igcebcV8gFbwDVZ/HiV5X6/+b056Hg4xuCOTviMydY
Z0sOfpgWpkMXTlec21Qde+GEzkcIdPlBiWFng3RsFnA64ShivDyH/Gch63XkYJOw
SV6alMxwX5A5NVxnWFMvaKBGZLjqux8/cOQbjEe1tCnGqORmFdTJpBZ9HjUVXUGc
NvLHW+U11vlReL9ncHvp+ccsAv6WoOjl9bDEferyDfL0YARqeHP4PoF1pbuTFgu2
OHMWZf0NLO2LAJm2cGy5jCwHVcaI8FDmBH4649Jgg1pOBDOKP6ybWiACdL5QaHvu
H3NIYpKsPsWu8oCLYNJsGAzGMRCRyJE5F4zLSRltzcnwgrbeVXO4MjBKX+4uJtGk
M4lmWOpyzIyK5fjX3Zw1l2t9g8cGsIikV9lzdy7b2lenvG38/VPcx/cVz1OSU79c
VZY87B2Ldt6kdJKQe7vffF8w1Z5UNS4yA6r9zPSh90pbVbAY2mbwjLNQopptQQDk
afeBwwdhKflnA9Ywqk6YFQGJjRWhSujfAgQH3KY6jfNdJjOm+ZcFGXOWJM/HUzpi
HmsBYAENGMiwRQvBGX3wQkvDRecKahZejfCWL6yDPVNO1JqvA7Fkp3zeueAqRLH0
fMK9L3TOpG9bedvdg/85Dh/QZ9yxopE+113rosD+YAURwZpFydOuY0/B+SYAj8bA
JF6CJWgPQMcDqepreThZygqxgBwT847YWeJgaITKwiU9PuJam+wo9/B0j2YKCKuc
IP3cYzFQQv0vBVVLK7klzSKAEEAUlNA+F2FShuMLfKzj3m+s+ir2SG9YpU7HXUAU
G5CDyJSNBlF06GR4Cg77kc0PxAJ6Zsll5c82UsGs8fub30s5XDYS0/p8o161OJCU
W3Yf256AD/yeHLvzWMt5wD1hm/3Y1sWmWDTtAgyPrPQXuJUW4PU8uQVLKC92vXqp
jhDGpcr46LRJXDT+BeTEMz26eI5SAOIMjK/ei18ef8PDkgqyZXxtbF+gFo5RCRkb
YBVlfZ6oQM4JxQ8Efs720ra8j9asQTvAj/CRprOC0lvYRtqFG34/t5xG8+pyfhuX
/fTSv2NSaOnoW7VkQbn51ZWKow+ZiAnF4UMNyxF2gMM3M8pEAR3E3HtK23lc0hM2
5lqzvFicJeNY8fvmQFmnkB6MxkY7mohFRl+iCOg9DreYBn5kJLSe6LwnQ0uXV2Tx
TV1NpN6kp7NsmmlXHYJtNLqiqa2ivapyHPonypzxjXswSubrwMSKlOBzVSwV1jzP
j8sdMUDnafK30j/5MLpxYcNPm6Yt5obOt5+vl3hROzpftF5SUFVj20L4SqbuyLAs
Fcyq/dVaLsfzOwAachZhy11dVLQJPtp769a64/cqeUK01s8pQN5ejtIOrcJABpIp
AVuAtms/HGkQlXhVeYzuSYVV4Acq74IFfoYrF8xc3yg0PGUdgwPQMEmig6GaW2DD
BCMxL0wkap4d6achpQQBTm+Ty19jT7FUHGlaKSlzCNfUsUQFBMRzjdwdmCg+5pSN
8MOvfhQ2rmZjObgL48DteFRcjmMJDB+SqPInStcD80MnBxw15ABbyafLxDCxokah
BAKabc1d+ZlJS//Ot+3NnCQ75JY/6bzr3zM6fpfq/GdKOf6L1FW5fmA25baxraXf
oIcK4RKtjlQ2Ptj60WpY1aj8pI2FBukeVrNCkyyD1VsuT0tSLRd8t3aHhOSH6iLX
iH0nRTjInngj2mtfLnNxs+rlHyvD/hKT8sfjBSvsEoTwIxl7hlFkdOk315hqLMVQ
yesjzDx0EsC/e3cMtbHaco4V0fYmqYeXOs7p/PfT/5E/xB0c15jyAISCbcfCLkO/
Y9IHJBzxNXpJwI1EjyGjdX9ghqPbi+k0AnstTrfwy3PLIePMttG0RdzbDk+MXdHJ
y/9SluFAnLHIazE7soSajbpiDMnbuUkLYzbI5XRcXplSXKXXZWSdE4SBkXaWosbF
P9FyEbz0cv3yD+ldHRq7O+wBDerA/I2rLOkMBtMinPp6AmycUZYrO+5CN6P7Ncyc
ZgRvX79jF+tA9zgeC0azKAVH7IZe+wcBBzCNwhzEhcDUP0tqHOJ4XXc6KhI2to0W
LRzRw+bYg7+z4kWy9uvMCJrGYXMcgQb+t7RsPPggUCmWfOOq4amvtPZWxTZUbmIi
JGX9EvCvNgIJaSePn9iKfZaS59cPfONkiO+3W4Or9tRH8yXnCoxaYmrhz+jSz9d4
fQxEg+t6lFB9OVhkvcA0sD8f/mg3UCU44SNBpMBb7WbwXjNgopsa8dp3utWnIUmo
tn3CIz3Ge1uR1A2LVuCEEmo4STbI0OIdz66uzWaSNKFsQvH5artQC/SzXeCebXWE
CbT7qryC344adIduu8AJqTjXRDNyQFxxumsen2JFv5QKySL8B2yx4sGPlW7AFBvs
Ph3XvE+ulRuk1xO3zeTwYTC42TXoiKd7vdqE+QxqQPx1QXe27Ie8/DeoRUJlIdj4
4C7nTB5GL0Rn8IB28ZqO6izgmfiZhzOEHC+FVimtt09l5ZbrZnFs/CmzPvAIvBC6
VNC1imEATacDnPE0qWSrq+UDF25S2cqs4oezmxfX5AkeEezatIgBipcckAg/1nRI
1NnobUgjbcz322AdYK4IF53czPUr+ADY2fKdP7XtWWQMEvtqMFoZRQtOE3sOYevN
0QvZzlEIGR9MTpqR+OalxmMrPQeCWIip4JhiVxInALlb8+qAM8FF73GmNCF1INdJ
trQvt/A6VrVCeNmRZxMzlJ2dwn7gD4wVAYNRDaHxdQf1KxJvKFoUQAoP0FdIiPyk
CjcWgmc5QhP+ZomT9s8bNDyyJxk48n0O3aeMyaGr7n3Seerexd3TAOgRnjpJFDQN
DlTnDcmdXuB5FwrdnGDlJr1v49D5zkOABJ/e9wYJr1svcazZWCDbfcfSeErMdPzk
1+YrE/8S87rywTafF4MTbYYQh0s/g4kY7Tjgb7ywMZchKAy2Fk8x2rIaFAS4Xmfm
mgq2frsnuFo5/czfDzrF5Sgci5/u4i2mp3/0HiXctzs42zqScRB6MstJ4Boitd1Z
MJGd9JVS8eCIHIsdSp5oFQLTu8N/FqZZbMyQAv2tlDxUn/vGBDVXA704ig7SE2NY
MwwTH+Ev/J6eYwk+AlBXzQsby7BFyxH4epD/3pJA7Pw5cDdqeaVU57qPe1c3Tpp4
U8+4vVYYs/U6oLx/KxpCBLYzcLO9NhVmu5vwykWB5Ko9xGj2SxLitecNFSAk5GNi
rVO5ejvlAmnaP/jb76qTJEYY1hj1O/K060AmGEQmheEqDUvYPlUh+wj/YnVo5kXz
JEeZWhc1p9imBA4VNwOM/eAV/lvAFkB86kEJ8YM/cpzBH1+OYgKkg8ddkH5tN95X
BX6C9JMkvCCiZVUc1/KHy7e3WlQ+jlKJaBStErHXSvCAatqhRjw0fjKa/pfi/ME0
gxn8mrFuq2/wkGDqV81xPWUi1aMTWyJaiQ15lhdYlJhZ/uaHbc1oKdEvaMxgQLQe
OS3ryE90WTwLjjvKxEXTJSKCitL1V0oprjzqJitIuBmQzZv3MyD4UW5gi1MTCaxz
393CYL5rdtNGqlvUFw32Lj8M5t6Jd0YFf+S4mm4iWx7KHL4uxxS9YtpdyJUVJWK7
dlEDxpMVL7RZ9WCw/VKxoNmcaHe8gydpW8RtfClbj5BU83svaIOuj9EOfrZVKuHn
Z3xwARi1MI08Vzv4mc+8jJSOBiL15dYmx03BdLING+n2i8jZu8kRfLdMpjCelHnU
H77gvWepZKg803q0hvemPdLxKlewKl/bpMRpVRu65FGBO0FH/kt0Udre37vlhiH/
VXB4ApHDt+voul+Cpa5Hii5faznH3/f7Ef5s+zDAFFHcELMX0v/jRZXmbuCsG+YU
KdiWow4+ldKhG4OHc6aJBGG5xeCcplp+LY2+EZaaAtIRBugMEQd59hWp0NHwT8Z0
cSAAxBRgma60itQOLZmNz8n6dnn6QU/3AYDZrAPCHQ3yyz1bHMiKao7HhNLpdx67
cjBzLFdjQ1IZyYO0cu0He/lBQB6UBOLz2TsDcCJ3Sqmz99aEYTH9lEAF0KOIS1TP
4APzqqIu0drXegfxiOmByF8ah4dSwMN54LqSn8ya/d5YfvSeqYFbPsBQA5lg2Qg1
U4Khu9OF7yXpSRR98GOEMxBVKY+gZVJwb6eK/gF9kBdARwk39Dc4R3lfsQBsC9JS
3RhCeMulQeoaQ5VRp9JAs1iDd8GN+seSMXygI2EH7YADBg5P3nsUHS2JU+TURl/d
WW1RN6XgMTZsIUc6ZM1OE43iVOeeQr18vn0uZGG0nT2CXLs+76KqELqNpX6UWHcc
gc6KBjqjp/jw9GmitNrsn55vp5B2k2YOegNn3zVS6Qsv59qEzSqNX7whBrY8IWeL
xOvMkj1QAVgR8lSJbdyHkKS/oMJgcsdPocyjmykLuAQT5DF+8AWriRe1zuKrycrO
WrjikeO/ACPN1hhJebQYbQ/nTxNgj6J8+ELBhgMAKl1Q8VjZrspODAk3AtXb1uW3
DAYfZ4aNvCh69SMslJSGv0Ksc7R2NqfwL+ZDAO8A4bCmdUJt8aoI0/uYaoFuH759
UkhgaEZS5io54AXpR0DZhrmgLVKR7WNFQuzTHalNWatNN04ye/hje4o5XKSL0/4D
y0wBqlPzQfhKHZ0Y7A/r85EVtZLNzS6MAofNsw96VL9pqmr/4bbCBXQthg2xCqlb
BTQmXPmkuuo3BI71bkXd04d369rU2sAtd7xlVnfSk+CeT0Qt49/63LRXvCGYOBNZ
ssuge2n5gkZ9N8CV9695FwK2Bvi3gRARZoQPZRrlObShZeTAao5+ngWB+KTsaW8D
GAmVVfs98paaKECKDR65MKQQMDb8YxdGk6jyiZ6a3NLxJdKyJ1xWyz8iKGXFAXFf
AtvFRxDFBY/mSETmx22QjOLA+cLv78Q4DIdyNoe/1VHPsk5HuamNSsnFEpC+5c6j
u3LFfaUwtjdWrXvz/pPYmib7fzbbj0NnseRV+CDjySZkX54iRC2CB9Jf9J8Str2/
zZs1BgpDF9MtoQBlWrZDOmYqvbRY4QUBGFnrXAo7hZ878yx3VGF7ZJCdPQ46+Nn8
zpsSS5ce28N6Ry4fb2ham5OfHc+H0tlBcxObAPiArLXaUIIKBZnT0SoXiW9iig2L
wXCudAmOU73PMFRd2wY12BE9Uyozw24K633PbrPl/L6yXMS4pUReeFKah04jqo2B
y8UTOUIDcgxaEXX8jLv9aYkgACH3vVLuw8Hw68nWXs3ROH0raspRvms0kz3DozVs
2x7N3Rz0pVMMe+HkJwuw3ttwUCok/oNnwh9VGbhr+uC8IIHrRuGyehYQU8SrqH9p
hciqSz9El4QanS0Tf/cJcP+TgTYj1BhIFvSm7/OLUS80t3RkruX3t2pj2CCSUuWV
EithMQ7XiG7wZPgHD4WoJJRL7R2VnhAqT1nUoqxhk7/d4INilZZt/yX8pOfkJuPF
mro25wufgAwSJbUKphkmmJQYn493G9rApGepVB9TL04HiUkg+wrTApsv7GQB6Yw3
Ggs0DT4802MPgRL9CCHIB2uxA3x1tEloJjnWhkpXkIcn9I5tWnRkIFAoV2eZ9zTV
BmrIhRIjbYwBgTlv1iT+ay1ssv+5d3arvRs8Yg9kCZ56Y0IRhA0iWmCdRvi3r2I9
jr7qCz2zjMZruAhFpIdbVYnjNX1L/k52UWLG513vkPVvK/0I3JtbByAbBnkem2TV
2Hwrr1amcp2qjRxnCfPjYNXHWFnOz5dgg7XGIBssbcWHs/wv6c7vcPaXjNiFKemx
x4GZEb1pzBJuxHzZfagSbaqP4R+CwjsNRp3qNfjZll3rICj4TZFLXF/tTYUga50g
rrY39fkHvw/alw9gJaoddNV/qCrlNAfmeBvzEm22QN5VdXuSoHhsHyjDP9ZlInDq
7c1LUt4GOgrjDjnR3o1viYZcAx1zuABRUtF9nULHZJtSp3EUurD1Rp3WtajS+oRf
BTCzKdcWt6uNYlpfdCdmZJZfb66X1BW2RtDNCpmPc3jSZjYHu9RSnsDTZLTF6j/J
bUrcgT4mPDikKXhP2yDxLtGG3m1TgK4YSEMupNoIuQfHlfJY6a57v2c5XmBr1hj9
9WSZK2x+rWVpVhsL0KFpZdMqtYjfHeN/lQSzH1nq6esDPCq6CukS02KWjWTglxs0
YYj9aK++doCCMIlWxwTcTXSIQ/t1/K0ry39+V5zzwiP2+v6nthZQZ5cnrSexdtvY
tusoXqUll1YrZOU6AbpgKw8uLQtiP6m9L9aFXKQKI8+5C1DMN/4kiKNT5DNertH8
BL5SyeLGgp3nUZJlU/MQskP/Hc9Wp25H/XEzAVdQQvDTXzak5RBzojnem2ddn9SQ
WzvMQMTQWc4so3+oXGpf5q2rJk5sah7JElB0Q8RAgRJbFRBFej68TKmx3DdXFxMi
hK/Pi+GRYBbQrF23+0klhPfW2TxjmBpzu+5AEsrtFK49Po/jti7CGOJs3+C9qwMq
jzhaokLWE2E98MSpCuTmaMRCHaQMcNUbVw+V5bE/2fYSQE9B3fST81jDNw6QWqiV
+zbs7/zgWRbXSiISRzjzkosSznMa7Vq0NlflTGaGv5fWtEwYYOjeRk32AWy7ZXux
yRTwXQWkVPquCTjYVw1oqG3c32a0LBum692+YLQmTOMtwOB7BIwK0sGpiQdH78qQ
jOAa0sa7II4DNaqNIOLrKQ==
>>>>>>> 426889eb8ce467b9c9a9f74dd4af433c5046285c:deps/flexrio_deps/PkgNiDmaConfig.vhd
`protect end_protected