`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6848 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
TDkIdcJUWDKCGvmrQYRemJx7xghVDyeQPUm/6J/zmY13lHOkosGaGGX1sEPT0xxu
0opLqpYNZELzew1/8RQgGTEZTl5S6hLxxhH21m5EfijA5TZXSThKP7IVpP5ficKJ
AB8SehSELBKgRm8jwwrEtjCciWKTusiURxA3kEjof+3hmcpzAQclQYlRXgHfAIx+
boUUZm6e4OCJ3mLv39DkdZDMvEITeGgC47kjlIPFyiuLglsrYEcbBK0mzzjGak9k
F/6pZxFVJ8HZD5R4yGI1n1uG/9tgrs5dozG8wqc+l6pAH2yT6heqGED+5/H3jI7V
FycncjLIrIR4V+jvgEYTpMj75X7nSaaaYN80l9Zyocw7t3W5OSlHrdeu4q314FJE
LvpIQDwlqnEBL4YVcZMlQgMcCN+r20QYKERAeEgX3rFco8uqGDZTKeNmjKTCJeWn
H79nijz3PCzFAkuSS6YhE99nCw8pE1flBc8+xjzJG1I321J53XOM/ZOUyHalfFvw
iXdJ08+IJuu23woReeezKJzSWpk0bcomaZvvYVAj6piPF4SqcOV8fv9ohOaF2f3p
9rdQ+PX1psbjwTZlq/UBxs+MnjNqdGHVbD+g4ydsffAt+CknDSRAbyfuT4s3t0fF
oT7ww1wOUOeOZejhxOchfAiaxOEIS0dMRpSBTeK/Z+eNeBABPe8w28J7ssUdjEr4
ImVn0EHp4pQDIiMJ3vxpAWZgEOVZlszU7ciABfYJqxqiSzFndyHiiELc6mDGsweW
QNl12COV0GP1GrCnUPQcJKa5B+MBLAvu+pOnfLLi4leNd7HneRy4Z7f2hqMB9m1B
CryOEG3PWkPFuFElf6f4bhX/QRLXLpiFF0SVdj8kSppSklN+VMVWeQIHAcD023/4
TNPPk+upm4FE8SXpzBK/lG5mHIovZE+KunYr104p1G1l9QelcLHwsRlzRZggoDqe
3ss2Bfj/8Te1pfPve6Nzevp1a9hz+3985D9acwFFvqVjmiqfH37LruYBYO1Hoiea
bOgo1Efnc1aSv6TRMR3TKYuAo6udj8bAA+lfTbLbnuFStK8WdBJebsMGkUThUQXA
69PzY/rswjyrsUcAO+emYjyv+/58tyJDy+l9toqmbsLB91bR2mrWnMEj9QWoXEXP
AiRb07FqEKmq3jj2hkBuaKiR4IlDTiQ13fEnKwqiF538R4S5WWPSPOpDqn6SwFqO
6IqjXFWZ1KoWdYvk8Sb2Lz2EeZvVL5ryhNZL5TBudzJdvCT29ldHVhvE5p7NFqR4
4KhNROK8yPqp5otd2ev0TTUQMnBkmHi76/kSP3G0iUVwvLG/GS2lkx2gW1z2l3lf
+qL/prgWgJTGhSq9P244R08vZWuKKCgWrCQlOQ2PIPSCO+uLKQNSyrgo3gT5H+Gd
S3yr6fI05sgH2is0GYnfItDpxByUOX49LNW7/U96T/tHA/QwfcOhei/KJhoVJ35r
dO4XezOWtrPkHdxETc94W/HGIO0rI/ahtK7TR5JT7P6w+yHxdKYOKIVZhE6A++qI
qluQoGmnW1pq6gIh6T+4XWp06Hg1Vu4nzpAN58aMa01KSesFjDLHhoN5zGL5wuPb
6L1PrtCKxbybstA/EmUuO9ZBKcEKT/62ETOZypEGWIhVKfiWkqaIDXPdJoflZyXb
afmg85n2iAh7NPNTSctA+hUEpCoYPfuOtaQFofYEa6UgdfeyzvUGYIeUIjXNdPKV
mWO3NMD6doDkK4g9iMX1Rmz4BLiYhhuDiKYa43rQeE35evwSJqZ7X/3FFauCT+zV
Cv8AOidWMV5Hh7vz/rIYmj+bIa0qtJN/+S/D5EkAdM5PWU8QrG+dsoM4i6ZS9jH2
eOWcKakz07bbDPkMkqVQrtvgN9l+gZ5zBYAdU7a+j3CHBXDwPK/yJgC0EJd799Ci
o5nHPttWPG06UYIdw7dAs2crFS+2o+vtDUDRMLrw/1CGzns1YuB1aT99/n7D2ld7
89i0oLpuDs/OAoHEVVQ3wjhUAhuXb+EERogBSDjnhIoQDQSnBty6XlzYfBAJ+sXO
zp7GfFEChBWfos+jZE2osEMoJMUaOvpCYEJKzPfS7gwlIkaXWEVpoB5/zUp84usR
umsTMSwm4C3x7xZvVA8TDpa3ltzH0SeYvzT15BdUI794Cet8Iezu6Smr+xP7n169
xQGNn/Np1cesSMQAgrVdXdDVA/Xa4wT85ty7cyYisjmMIlCl59YTWUIRxtMCeaCm
cVeMeNYVU0foGoOUrUINzWHnehugnFVBDGz52ob03PXxx9TjzDRU6Rsr+c4g9KGi
g9DkV93QFXyqoaXWZS+YJpfMb+3Yz7+y9smPW4+FBJWkRQHC1RTTqQ5tb60jqPXL
YR8oA3X3ALvEzIy8ZYD1tNrI3s4JgRnB/Z8tXyVuXbguS9KQkIoUQHtTqDqEGrTG
gUJr1OTMQgM6A2tj7Hla9AGQ4stcIKMcy/js+KJroJSc01WV5BIxupKoiPg+Jrqa
SR7b8YO2+6sRFYwHs/oOJ0U3tkKzuS9gSnFpX72pBpGCsECrnpz0cqPxNMU5mlZV
UuA1X6HGPRbKESLP1qgHyqEzTgCNdZvzr6bH7KkSjZbnbWztYFY5MnI/6P8kIhZc
EPDz07DDTM6pDtYbtP0rFgKA7vKtgqVuuKgHH3xNoma7oBGfGxzVmj43TPAV9hm0
v6ezZca0JyGYv2FEO2uv3OhU5olEE6HQry5x3G4gLjMMV4O+C96y2wHfU/NNeltU
Nb2BYE/R8V1r/3mFsARFV3F40lugnm6PZqxhLkAzY1n7opDusPMK5bnGQdp3kFUk
uVglyyR6cSdMFdfasRtpxRregeo6jUY6GYJi/eWeVPK5O9qCP+tWcYdRO2+ZFw+/
u6OmeddknAquFH4XEnIWve6pLeByWG9QSbeKkYJh8DXzEzefO1ceYzWj8sCu3/aA
nB5xLdFvgdjhxwRJ3MInFS4LDI+H7RshRgWjeM2DB+Keq/8HvdSDyXMyNAO5qMlK
hR8fRem3AjdkEewUbA6n36OHAtt30Vtwz44Lp1OPXy6sRSa9gPKBP0/gv/eqGXCo
7o/HEVHKHcCAS0c3OsLOOV3Qr0onPA1t33qjbsrlwf0BopCd19svT79mRVCci5IQ
Q+BnI9kWL0EEkhbx+y3c/eR707a5zZ/fSBSaBSmSO/s7fwk2v5436c4EhTeAjG8v
xFLI+C+iIH2Veh8NBwxB2U7s0uQ5iJrSALpfNINDx3g0b2fTkeryWsrjAU7MAAXh
79ew+EzyfdHP6uMsjN61pSCe+I16fcK9n29Tyi8h/bsKnRuoXx6RqA2hi3V0Rd9U
Ok7OhOWk63UVfsLN8PHNfIRsbZEhyYuSNRJ5kdiwMRbgcZKQcP120bmPpxjNAPiB
UTqVc1K3YYUEJZ93xm+fpiAwYCuaE2jheqp9A/ZJdMDyALOPowQikR/QZs7/chh+
kC8TJSbpWiXJwVNnv5cdl7xcUe6h1zc6Na5jPpV47HtPx3Wc+J79swOTkMtS0pEu
nkP0CipXu0/cpYa3mXYireVYWE0wuJbNX8Qu6Ud6bx7RIygWGuCqH9bHZLmt9s/M
Im07Czg6jq0xOn3pChWzZKrp6wumBv2FncBH+1y0ohr4D0S3TZT3ftyaLd/ucgXJ
KCnn89MPbB8ZcJ92iOV2Lzjqqil3C5q3x1nHUgXmsTFI0V13VneuBQXgViAMBsR0
w3nHS1OlAnmBTx7LrZQEQNEIIYEkAmJbGkdXpvOoGTwYWmFANIuze2ef7PUkgFvE
VQ5XdOYJH8iVFJP9atpKvw0ryocM2IZ92noacA22HwajIyuyP0ZawLdMvTuzfab2
zp68pmhu2shn41PyaFg760dRm+uBjBq+LlOcASknrZCsfzGfV1JNe2r3xq45ckfs
oBcCx07QQXXWALMPfSHbittaPZnmnJ25nTQ21/S6L39IjeA8uwBvTT9gH9tKsat4
ncMSD8o20Gwzjk21ZCv8KADB1XHiIXbLx+OrmGB+C7d4RuWo967gqz6uPri/fYJR
uR4mEXMG4yZL11alMHUpJhlTCkVQUkDzUaGY9/ipJWXdb38QNXasX2DlWNqhVsm+
0CO2XdkobOdmeNBXd8XJeFQez0cYObL9DN9W/bd7eTANDugJpYhrN9ddVvZfFNVS
KHipID1f1a7gRTap3lsl0pCrZM2HjE89ie37neN9rBJlqg2Ne1K7Yq5uiRfIEvNW
6L9fE184L+RE11VwiNJHVKGhSQP9oA3f9WYNizsI83c4ZHeZnIFvKjyrxx8W847A
VQGJDMx9Q4hC4oxM3w/TJ+A+0+z5+fAALnKzEa4M7fkkvXw51uIYc+wsiOHydesO
V/Oi1VzNxZVqBDAqI/PRiIbcghAF/58lI1d7Nrq1K4gvKTkMZKzoUL+h8DLyKzqG
EeUDlFabvl2rVidrPwYqPO+SXbrpzkoEIL6/HHmCGJ0RdTE4K6qbDbQStp6LYHZC
q8y69UNJ35pdGkTnIOkRBd7HKePKWZCJ/S373swknqSsz7iFd60D9U+AjgJX7Scl
Zry0KP9DYJSHLWXbyE3S9prqaCovJW8o8F5O7lM3pWfUL3Rw3LBcXhma3wmmQF9F
Xng8G4GpV35W7E7KbdJvx+mFrUTpmp4Yn7jgzbiadeOmQRd2cHDgT4Z+JXwpItC5
i2ux1H3zM1QvAZFeZojbkM9CSkGEvDB+RYf6HgoCXZwsKbOHPMFYh4ghO2jBBZt4
uyIUiLzOHIrBn8WR+IkLwhZnxeMDYjgdpLbU5D1I9DxxntymuEqvkyF1h6Tf/IrP
4tAUaHG8/7P5QWN0Ymr3AsGgwn9uScojSgdJUH8s5uS1Bo0nkLh0pbBvPg4pzmkG
Q067pSiWclDYk5YlZs/qpLQnTa7KzVYhbAMoKzLNzMzNN7IXJQurZmRi8O9zHA7h
C+vjRcAZQ/0D12mlFIw1MRcriI9fR8iw0y3bMSEEWQMcry3OIUxZfqDsmhsEQy2n
RG9u6npM+M01YO4qtzTR/6gRgnYFYhNIn79yc9aTWlv8JNie8omXvEekVv9X2mSX
+qCAwD2LpF/MMlIPjmFAICBfktfwBBr5UZP8qQ45W6CJNTFtWgRIRtcZ4Fd8Qb5N
v+hp9+eVweT+wfiCuSzvaJ56ovm/n83HWOhrhTk1tJel/28HlwdeJdAg4lJMjZja
hSvjnQRI3pHt0m4FlSP85NAsGNwu8y7OzqM1+JlNZLbGGkgYWEJoHvJKokJSoR5Q
aDOrN+vuzxBcAngyEDvcdenn/5lGrgydBVUHBBIqpGbRmOQmKN6QnXsp+tUkxb5H
V6w3n7uYSWLWdzLiRH6Nk/w0Me4AnpzSjhaTh2BSd/1USBIGFNon+KlWpNqS1BgV
yPCKoDagNHg94+PD3ZZrdAtihn0UbUqQb/GITk0ipRG+bn5eXezi2+5Ra0D6SF3p
/zSFq59fEk2E6nh5rRn2xH4ix7hux4W+0OSMOpq+YARxO5ojFxYB+yNyY7nswT0H
j2SlqMmP3iGAHDjeAuZ1lDq6D9aY1UYQoE2qhTQ1Mzm/8ceavgv5iti2PIp6MxrC
0UURZvbTbSqpVT4QlWFK8mS6Puwx9jrVnS1IevYESKW1AJSvvdEYL03N+O/5/TEc
g0uS52/NN6e1L93uticQaVOjFeL97XJNEKq/Gll16sZgnp9IVoVunRcTOXYsGuck
80h3GFIv5pmN1YmP/AKks93U/g0+Gjl7bwwuNpddF3cahXberLmNSU7C55Bo23oP
jakYlVzaoXPSb9W+xgxQ7A9xE5XgirWfsBDtuzuaVC+wEzED0JlaR5dDjRXwO+g/
3WW9/xtGGcdsvsEPoOt8A9FxhbCKRYUlq5NlGQFZY4MrVp6jzhKTOglCfnmaCkVc
3haO+y6x0jUBCHYvtHcaRHwQ9My/cz/Lj8+2ib2lVNmoxsMdN4rhCy24ggo0OkIh
Iszjd+kMJh1t7texaUgitQt+i8Sh5yn7YKNUrsW1ORsEeX3oZL/DLLlcBvFmpzIS
ir+ZaThzoqCT0d01ZR4Js+q3aE/+HQKYzYiRN0PrAComJcYJVdkRSOYIMz9KsXu+
9HHSpk3gQGCZIeI8Jr5cnK/FusXEdD0fylVaMGb6Nd7e2H7+6QBneitNZE/sluKO
2lnKHF9Mh2L1gtNuDZwQVu4nfKFSfZTxiFhOlEdwM0xoi2v2czouCOuOSTKBg7DN
C9EYsuYXVih8zoJcR0mQIGqV9X4Hs/y2Oi1hw09+8+v9k5chjIS3AF0CELYvSNMe
7TpW4dj6g0IO2d3oYjbGQHHLGbLMeDwlmRx/10+7YV4+a5jrbUMcNLRL9ZV6kGGL
IXTYzN5T2DSQyDbxKhUFb96DqGVF/rsv3c1C4T/bo/b84gElh2yMePI2Y/Mv5nhj
7kOXFtxewrF67JtWbinaplh2QpKnYiv+daRsuJ2OC99P+W2StTHr6BIwnb2kTkZ/
gbbeSzlREeN6FMA1NtJNcvp2aMJZLqlrmI7ljWPmCkZc18EePatqYmo7EtkSYTRY
w2p2MM+ptFapTwJd+/BDTjegQwjdf3kgPOnG0lSHb4XHQ3M73vHzMLNYxgX+DV9I
XYt2WZ2ct4UIEOCvw9j7xJKroVW5T7X2zgYq5prc0tEko9AFrAUr2FF+Ct8Pf0AY
15PfKVtOrhZd+J/KvznxUT+8AyU830aRjo/gUkjQBlzIRaEcB6zFVTcqfLrTR22M
4/OAcbfSQDGRIw3/WWAk8+N/G234wfNWRrIujbHylFJ1scrdJQNkVMM1o99Srx7B
T5VR6Kc3eYoX0Zcsh3jyaC2lx1cMLCkDu+U/DRb961VqHJQFKigIOoE2C7RiB5Ry
dewt2gWl4Nkwu2AySJVevxV5QPu5Su6m3NLI5MIrL5nTd5OcRzdtoNQGbP99Vedf
YnysGmGtjUf9n/cEsIF1JPwrfpuR414Ar6OUfI2EDsdV1gxTjYJV0CTw+9KGQbSD
AnSJcgtbqAmdsCVSaM3Kzdes5/f26SltK7EXhpumvcF9Wv9oyQy+O/IFBf3UL9/C
FAQLqcWYNQmjoZeTIAzk+dLYLiIvMu4EhJHB0oB/tWt9bZgfW7kp5ETjc8CBMWSd
auJ9PQi0TCAnFEGJlCFNQ5qJgPL56iPdXmWgcznl/KMOFlYU79xcsQlHHPkSKTPw
5/mBJ6MTd+A8bgPosALQsty/JcNd99zz5kkBxaXM+1QkudYqdNLy3tDRV7NHn2aV
En3sMQ2pm1Gg3cAfohm5Ql+QZLy6bZGMdiCUbUmlhcj5CHhSFQNwrO3X1yHZ4TO+
fW5Ppkwef5syjs4JX5R3JEFs7a4iJZMPZ+d2SAY0iQOei0XWUNNqnimmTZXjm1nl
NLzUN+XJH1igz3PceXJ2OYFWufn/FYiEMuvUGd3YdvRRQnFxJpJNixeFPTauE8Q4
cZRHRCGhGK21wp6DTh4zDiwdBCuy3ghdRj1QRn0Bq6bRlKP97t3jEC33Irr7QkiM
P99tdKiTY4fkf+mHPMKJma6Lp+paxWstM50+Q5J0tLm8w0oglfYdVZF+QOz3/rMj
0062LFuY9+5GAw+K5dVSEyCcv/mh1AIobcaXmA2pvgCnQTTgytxjQLCIG3V/fWVC
qnE6h+32tQVnPDxz9EY/QfDa9HDpor6AMKSU7Ut0E/zo/4BTW1Ki4cdNDD826PFZ
SP/1VRJUa6bG7tBEn9XtD8PNEou1DTcfG3ibGOti5h9kj5ApvMheyh8IV6aA5t7g
lWfylV4BUMsv+F4RGWoIFg4okuQ/qFwaFU7ZjMGaPy/RNARGHsQkwx9ihINKofrF
MO8EuMtl8q9Lb9cDICnBy6ko9s/3xXo6WCh7Ma9e7v8G4F3uP7eppaxoUz8V3irk
BM89yzhF4+WD2840ptJ71ecaj7u4F2dz/ieqWMkaTm7zCaDBasDTv6GabtTIiNMX
V0G09QiuIRtuelNXXKO+jC3Nayp5J1RlQHaXErbUyyO+Cr8coDbGN574KCuo3+MD
ZpCZMgU1z3c7/VysXXgaXpqQR/ZpiucrMfm8iqiXdnqgRocD774RPle/2iiOFmfV
7sIjCS0/FYFWVUAJs16Ci+qTKX2pw5lG7Sy+qnt6YTH7Vynz3iJjxA8SLvTGI68z
wuhMSabZPH+4Bm+79e4HlA9GpRiJr61oW/ZqPpQLUTaxWsXoD41bxKjgjhvzdPhY
81rHUu5MqYRAt4dhLAzUv8US79JCNUHGLTo3BL+Zwn1ab1fAm2i1aTg/VTtYltwn
yUz9cioXfEWOze0LQkiIf67x6hZ+/Y9EsApFgf7+ZzzqpjmmRmNMQMYTGuzsJNUS
Tq1q/TvdQqfXevaKUIqAthy9hywHnwxfSIVTdUy4dCifoLq4kkNSmEqLPxgV3ecZ
hceB4JQx7rM153CiTJTAMlJMH6MjSJaGVBmM6FkxNag7hbtiThOw3RhbKHgcqjmG
y+srgmmATNLSidWq1Ou8axerIO6RNml8PmSGfRoXjY8+is/4nX+r60Opy8pZDv7B
XjPEKPYSuOiwDlb+33gODa8dhJIOTUdb/c4vQxiVSLxMvTvRJXha9Czfi0rQT7dm
F4MRGrkYxJcTnELL1Rtr/KuqK9CbYY5ykMdcN7G+jZ9DHLYgneo1f70DfbLvD3uS
/2OuM/QrGs0pL2bNDIm03qUChpAerXiGVs8cWtDx7NA94Ty7TyiGiD8SH7uu2pCe
DAA6pUGpVYtxI0Jkid2E+8dF5tacGERRspDg6xp9USqcFXI6Ectr1ngiUuoTHZqG
ThdihjGjlm4K6JpD+QZ6SiPRG7Zb3UP59eg/O8G7l75EiYuwMWwv0Qa9rE4AJ2JX
enSQMyLLdeT8fbuu56hxUD9r6x5NTycYziyBlT1y7n5g1lSSlbUfWE6Es186E5Nr
bjZkcUIi4BiHx3jlewK8NA/Enbwry4q3o5xp5euSca4OjcgfPjrpVfD8pLYnz9UT
k7fEJsuSEzr87077NmI79lRgHXelenwUIGGlYSK2/Gw=
`protect end_protected