`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2128 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
kzbjNko0QODHQexvxafFnbMOjkLlKfcI2gbR9IFP8JktXDIo2Iyp/i9kNufz9jwZ
ZjtVPbEecnom8Lhoz1asaveSraRvN0jYogfi6usAikqaIkTHE8eW5MOgxK4L1VqQ
IDIlMLlofU8GH33/useC8cojHaC4EcJzpTsvxAjdC3ld3FyT6NQgFhGpCQXKUx6r
Ry+aDILx28jUkb+BS6dQYs9Ex0o61Gls5aK/JzBkeuAZNvNcLahT6W5H1nFHujPT
Wd8nU0G/5RtnGG5wtj+ZXW+fEWjpq46icCBPLGfN6CHfZo/VCjs9zvfJZqy8Rz4h
ol6lrIovplzRSBM+wRMPZlzrXwYSVsbPm5Tzo+heLdyxYAZSF7H4LMmngZElHz0F
iU+Y2GumHIFbKQ3oX3RbdhIMq/lyd24UUSCc2hsZRQkNCSpdUqSgBddqZD32ECAH
eErShlZSM468V/1YXCzn65wWJgL5oe2bZcnRIaTi9VwByJ1tDSqw+D+uh0ShEuju
G+L7uBYzePXUYhZuSQu7+RYA7dxE8gOopbzKyiQtslbs4m2EvWxFQFqhctkhHKuJ
kvL9fgVRc+rsx3XsSJGITVXRz7NYQsoc1wKVUu2LDV6uur/ob6jWzdA+arxF8vyr
Zp1foRfP6Ac/czzsFXNDAwuJMYZdCOUXLPQPHnPvmaELeU9Idbt9A5jcgYOBzePj
AtSEyxLSV6fSJ7dgSLIdcQCZGj9D70THtVWlnxL8o+DMuh1kssmavTBZls9sBlJR
g96AvL2BR6Md1Vfq8APQVdRcLWuKbboeW7xVqHtLs9wppYBJ04Wmwk7ltQ6lccwt
C5f6yw8iqqHZQrSQm70QY9fE4CA7EwQuywQDudYh35mrlKH2U9vwzyBtqeBcYPbK
1hYt5pQsEW99ODkSLr415I8amsVmSfR43CBFlKFzIExC8WuuHEMV6w6C8FTR8glr
kIeNu4EU3FzfF+l2xtdSwToFgNC+nfBLP5+/gzheYsr8AIz16lUd1T2u99gpbJgs
G9GYCJ5m510+s4nHt8dl6zBmpqMPyjeriud+nuah07wdwPoKDU3OubtFvDf5CErN
uoT/FG7cp2aktOagDMvfJi2VxwCMR+KIPRf7rbEwOtuEo0B+tnqXceQW/G/eEQtE
n2A/IXwYVgX/RW6KdOKevvEwhZdeVeWNpqF0JjZnbJJj2eY+rTZZmPxSYPf3jjlQ
IaKNfJegdYvgAXXGeC3/6kACISXmWjhGU913Ko3bYOWwlMAoKr3Ply1qvCt44YEN
ePoX5HnQ7MVhqpRF+bEtdvyfUijS4j6TWdr2lkbaGMYyYrV8KX8xXZcsgQq4zw5z
UTwj0GmLQTS0Q0wjOGzYbAU1+S0CFa7iNQkAzGr5ghrYisXKzQFU4kBSBegEQE+Z
uvBy+/N6a/DSQqape6B0OZ+mGHausRMnWDgTH5CWN/ozeBdYj+Fjr0nLWDCJZDQK
LP1Yu3y5KbTSdzP/THHvZwTiiBYF9G75UuBYQk4QcQiFOoXk291zAyTw61F54OxD
P/jANS1Rhnz/at3LoypQFcObIn85SLHBZfd9IhaibGlHVWkBeAkBph9vW6V7fjQ2
7h6HT8fEp5UZeQMziy0rxJvuRRpEMfHSzGqJOByreqyzxKIFFjXzyfxctdvgK/D6
VKiAnD9cnY5A8QipZtSUjfSyBeIZNKGfmEkN5UzvRcftH2NXXP3vqVfVnTq+ml1Z
PzO3pkYL12BsVmfnyQYwCOzM1V3N+bKp/NbKQArW3o0AnR2tka8ZTpEe6Es1+RMQ
JczAb6Fq5OJfsjCvYF29mU+tZUagi15FsMtuc5mrhRllkN9UJQ7looUFWAPx9VQw
zjkMNqslBlp3EER4F4ilmUJoxS1he3f3325ioe+IR7G1bNzFGJA+Q8YQIzofzgyN
n6Ks5MrgIU0VRlbQwM9zBY67lMjkwU7h6Vg3micHCdjvaEwvdXqxF7IDmPC1NwSu
FmqOG53JwQR3mYUPHIjlH2JZfHAchnIkF8DUiBvHE9XKFvJAF78ejLZ9t0QyFOsH
D2LhJfytlYbf0XyExdp5tQnHa04Q6+WR+G9uosPThuxFGJEW8pfrPoiHLWnRZRxA
bD3YEB+4liP5xIAcK9e39NuxPh2L5rnZmbGx34PJ88MYJP6iblzHxczWF/SCyHxN
d8bpIGQZNQaj5ap1JHPGU6nob5JMNOyOYPw2crb25Xy5o5uAYQKysagM9s+rhwYU
GXRDWU2Q6YnEgBC4X+MPh8VEHCohJL5mmlgVdV/FVRvPyH1XZkstu0g7zUQMT/ZM
T5gOliDQyldNgxpRr4U1kiznOUQyzLggiB1fbkZUBBbGwhtnzI/sATfLpKNn7yvM
F5bHZZ4HKbc7zMms1TYnsE5nDUIRkdCuRHN6PKuJzI4657tKual5moWjOTfFGVEu
fLYHHu8ZQ5ofn/pghPqyrJ4jiew7+wDhWo27m+OmqzGbPSmDkTxbcFJh1vkbbaDZ
sWpP5sNaoSk++BoXsHi+iUpzYf99/5O6PQihJXAjo1HHhZv+e2Ir48J2tf3vaquF
gy50V6L7lLf8a+MHkHbEvQnMjOIh6+YEMdsGCOy9qyjwFVCFP52U7TkDzycoJpW6
cnC+ZxHtDzkb/BkB4Ryh7oF6zL+srYoWbRY65tGx8zI0w4L77RjtewqtDmpVJD9N
KOlYysBIpeRVErjnIz1zbA==
`protect end_protected