`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13312 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
3urUxeojDObSx2NGJ45J6z9agCSGYA1utAsXA1ZCiJE/xOby0E0VGU+qySMUFwAB
tb5mVtxoswTqVUSUvk1fzjmGDQyYgsQGjc1EQbHIVxMn7S+VGIyvDCBgPms3wT0w
42k1Z4kgjnSAWGDFiJrSRwhjNZEmyHNcNu9niK7540/slcYMx/YwD6rmHTXFlADo
EqrUYLphdTw4KsyoHYeEBoS6fXkHERxdER2ShLCarc9iYEA5D0YjRL2vRvsWE3qT
u8R34X5QYVxp/NOkjO8MVe9VTBPK/oVUr1BR2kdAfbCKPD1f9ySY3MUZET2LyX94
w0gDnd2UaGTU6eCde77OLE+P6v9Z8mOoHnkvryzH32chDVnRFK33KWppS9B0MVw+
So6+s1d9+ch4wAik5P/8IIDWt7KNYuvAWJQ4xgemj/ytvsi2EUUDK4Sx960sh8ff
+4HfZY1qbzzSzJfNeZDo5iFaWrut2B+YuLIt9ZsCstpGcAp+/H2j0SnjZE/5BFU4
Z4C6brcUuZCfgEYRXH/1Bo2Zmit37vLPbhQx8ryylQYoc3RF0fZKfh1O3am+L8n9
aYr1ZxDkZOQ1GCzy8bw+HejrXjX8CJhoYxO5liheIRVPbvecgPkUe/3VNmb/Befq
G8Ur/a7tT3dJkky9gINi0x3/Lpax4jEjTOtgohbveJ0610pd2sKvtk0dYvsgFxkQ
7H5GIiYi80/OlN3BpszKHvvqyzoI+QQd4D44/0ntfh7DvI0hbp0ou+/Wu2YwXAQt
52xkYZ0yIc4X33SZSRyTpO1KxL82BIEfvbA1fxETtJN+ffCuwaAdaoo0kZNuDDIr
El6WoYcnimVjeJgV15hLd5MIjlJFKmuS3Mvltj+uTHacBKDloje/yCNUDZqynmTi
LSJKuiH8ISCsxsSRySoMJZNbwFVTYIVeli0z9+OaKWB695hHgGZTKw4TiqQocEgf
E9UhomZQp8La2rbvllmSeQjT7ynIJpY7BAvSyiRHvGGV7v1f29TsUXlpGwv9QxUE
Odv9QIulUz7aNMNgjzW+ycGGt6UucouLdzlmPtLNwwNoIUwZzd1lsEeofsxH+n0+
sH7a/9b+RPyD/Z1R5aLRYdMme0lb16gWWPu2Nk55Emg31WUOOHQw93wr7j+rw40T
gLkgigA8kRsqr9mV3Dn3i50yfTv6Ifzjvgcy5wH3OAhhhm4C1iiPpXbxW0Fr2ed4
+o5jH7UIZk020T/nktdMkAK6Eotn3L5NB29gsmuGGYPa0zE6eFQ1i+CngF2z1lmx
cMSdYYZyobTNH/6RYavdUWdRQdFFDeNHCQCZl2sza7WGUx6M16qZLeF7lqX3ex9o
/tjBq0p/kK7fsnZS5h+Q0n1UAtsjtTRWx+iPoEB8x/ejQ6oKBOgIAEX7HMtTeXKm
cLLRasusPQE6lQexze2W0xQn4UPeo0bgYNDidl1IIvTH4dRgC1GfvLBpi/KmB3NC
249tM5zgs/hpzpNtxA1+KiOy+wZRH/RF457C4jgY73BNmf468ZTAeg+rLcX9Hf6m
A44SCqQSy7kIWaih1iI/db4LyuD7ZD3dvD7IvbxVJZINXmbtzTJQqVX4EeTiYsAi
YY5Kqa7xVB8fmJjjVxlNshQxt4rFgirDHQYDeL8OzPsLipnR6YWO07qp7nZHtnUV
PcaKOEdzpgPdSh0vawEap7DEtk42ET9rSpmHd/2/VNw6aYzG7UGGLQ16DlxqVCtE
3wO6n3OMTNDTRLmtqWOAN1jRLwBcIIXQ6Jd/hD7kbv0vVp8UTZUW7YBhQ3Xb/PDF
g9mDUl+soF5AxfocnxCoXkFfYMsVsXjtPNe92srEKrWS+nyt0Dea3WD8wh7bV1fF
hJs0PdthbPQflUc3lv8yVjgES0MX9uH47NMnJjE96D1ztk1TGC67zPofzuI8vT4q
CoLyRmOPaROT0mn8GEjA5N/8J+NOmp/0MLTnV7QaCnj1TcJOAa9uz/JJWmXYkPc5
wpLA1904x+p29gulo0TWQiHpMJohvgEYaKsIt3/xV9cKOsT2AWbvdO8h8/bvoTxj
azbYvdM9Pr17vNGvfXDkrcLv4QOgOEBqSqVn/58waGCcOOpjcfB8RNgoiDciKr8e
Av26y/Wai1cqUmlRs/6qF1AVYt3sIEtUgj+g2KIoC35K1lFcmTUEjZztJtd8kTBd
VRrdlvFgGCDjkmhg3IBRPwnQwA1KfIO9qFirHrFqXo6TZmlEdQpGA2cZrmNa1JIJ
LdmJsWH78GEXaSZEG0fs4Nw7PuWdD9jUvJw99wUmAxwuNeXGFWhSk1irBA7UCI5U
UAZR+vubY36lww6oQ9A9MjUp1AtXjw7cn/207CGTbfq2tNEzI+QfC3jV1t+i+SSl
Ms9jaPbqJvFYt3LLTN61JqFFTAoKPAI2FsGBHHGznZYyO3kZ1iRmIWHB3L+XPTd8
PCaKrnhnXO77mDWfH7muw0NS2Hb+nq+edJNhQKyPSIUkh3QR9suO9vYNg+kVHjKE
5hDHKEYCc8aAmhieisQ2ZqMuT8ZG3TNGqszuUKyL9CSMNfDX+DIlLWuYu4ajCrYI
ObpNCRfwmz3DAcJYGj45NGZGoo/hXdKmJfZ/I0NozFTjVV4yl9TXxrKvSKaTP97j
Aha6aD6AjZPcic+2drnqLykA2eWbBjwXVBNUovqnXCTUZBrTh9s7JrTz5kIFULdC
7SnAosLEV7rezUa3BiY5tE9Y+G2YO/5Mm8pCb27QrhJJLrdDjh5snbEXv+c0PqhW
yQR99R4nXwpiIRSiDzkU9tDVIUl2hf/41nYgS3NxOGa6LxajeCDs6x2jlhsgvWlY
t0pnD1o276E2PVA1LZAH6NLE3Fy9DhN7WWQvTXhyvbjICCAuWGlf6O6rGvWXB3uU
lwvTeVhh/kwwCTnZXIiS8Lepgbbl2+NDx70otDwN1/RFaet44S0ykj3VbiqNMWu1
FRdZwwEEUxNBkawuiuVsTiC34qE9l6i2Eu4eVrkzoaOXBC3/Ntj28ODd6bZGM4CX
wSbYj+l3g886F0KO8r5nSpaFhe+W6jMazj6b3at8hTu3X7asqm1j/uxjSC0iUTm5
OVfppAvDgb1tzTAPcldVopTSRtsKYbnX6Er5Oc8gIUkQgVbXwOIxOAQWkbsz88ld
5BP2SMDJ38rpmZZTTZobIX9UXJ765XcCVxwe92GT43oRBtTAZqPVhLQ3FbcNxdgL
fHgcGBAh5mBhBZHB9WSsjyL30PRUHU7sV+6KhBtti8h6GFmw/G95gNsV44fnJEKp
nDLSt4Eid/hhU51pJWfNeuBH5WFqvPQ3o7e8r9QO8FU5A9BQ0XF+UnzV2QaQBVT5
FEAwPbEQ377VJBYuSOs3AMJ33HhmVRFMJY8U7lU5mc0onM/AJZSNGuzwDeEb6FBc
DFj2RmkEgav3DQ+MOWv7CsWkOP0SK2YHeLlwhfYiwy0SYLGWgkNyvkt6xRluuN5u
N+GQY1myWAk6+fdCHSeAbC91cyg3im8S/4sOqDjCBJfc5gZMY4GvndBWTvFVTqmM
lOfOmTq+YyoceWq000MgUYgHKDF2nDxsgU/Hto+cQgLLQtasPrZ+d9kFGUvYvYwz
rDMbzK3Xg0cJdzEBbRz7KfeMiMbatEBPDX0ZXd3aZKIOPZnLkTLrfDaLLB7hv0+J
lnhLilPkByozp3TDEXUAvjB/UW8qPALYpvh++q06SqzjZzICVlYgT2X7LDkbqap3
hufhTrioSuHMXfUUyR/455o6JwiNDTzus3PtCdQzIvvBpq3p/3+p0FBO93Yz8glU
bDJE0ecoHRyzEolU4Ed2SIgW1ttf7KRZ1brc9JtKb7GabS390uxl2vrufxYhn1Zu
bD/gmkZvjrcsdvknoij9VaeKeAIzYJyUv99nXMhnuQWr5tR82T9a8BJ5+m4K8SNC
Fe89E3dy8I6cVG3ROnHWtD89bumwRnfF1lcVCyYOyOwGLgADzReup7iUEoHSMYzm
fKXbgAnRIpszJjKGk8wAlqeqd8C228K+M1r8qsZSeIQaIrOW3yP5DvihvIzzHnwr
9/wyftzGjYUuEhIgK1olKsOzforcsfxhfjgrbXLIrZH1chkuxdkPO2wi8K30of6g
up9OInHJ9xOe9FMLVK94jIjc/BbYZhjpbe3vmHkn7rkZr0/ntvaqaU4T+++z6wvS
NdhKOzMz/LeqEjF/3opdJqoJLceOwwZ1ti56h6ydxWPs1AMnvPppYcXHqSH5deOI
t6uNc1yIHdWVOYiXkm2aPX35DrCuWlmQizML77R1nmp0tVEtMoxo9C+MJ4Nw6N0R
exobf4xYsBw31HivIZ/hivGUBpxC2xIfjq7dnSnFegBp6FRhQr0XmDZ1AKDw/VT7
M+rct1k3a4mIdSUDWGqZrslI2P0ji0Eif167u7n0DiDgBJDn3+0cZgT9ILw7dV/6
KL9ZPctJFgk2FUrr3x9hx6uMcUHB/Swc8W5e3jpdD/H+f0GcStLW0WlH6oPoImlm
LqcEky52f349leUlfRLw5z8liraqeD/AXZ0kcO/D3Tja3wY7j5e0zfd+AjEPCuI1
NLN2cscrUU3guYkg7qgtnQnoEbu3uqjSMTbUG0yEhES7097jRPRF/kkmlmxTI770
scWkr+vRefs80EZ5+MYgqDMBGo09ZzUfaCIpyi1EzN/i1QE2OShItP+HOVTqmUTQ
MHpPjhiALX/Jv2eBED0v/YjTwXmFdOvRhwTVIJk6MbtUcvZNzQZcimj8RODV/nA0
kscyy1zMGhRGa5th/cGaB5qY2BTFLmqVcactO2mNjAu8v6H7oH3Z01dDzJDjN2xW
HmiFKjlHRp/vXo7KKP7kadkk0+C0pKvO4iEgyba3z0wUGqlgvLHW4JtM5ly0wvZ/
a+UXZYrlZgOx3HwgXISfRgHKkeXK67UHjJnTCR4ze31GqQQjlJBGchanhGpbCajk
jKPxC7YHm92XKnAb+YAShbnyAFjjuw19Pr5/nFzDzTXCaOp0VlLfvyRPUPEt9jiA
smwyMflBSFuK2xVw5amUch05fu88Oo59MgcwFrAT7s6y+KFh9TdqqURyDPH4gTX1
NP7dgqOFMfy1SjPrqtsiAYTppMcn1d/ssvJMVqep8w1gM383wgdXog8G8Ab4ndj4
PdQReJ3SiubAiaD/A1XoLe4pLHarGNEWbYgnYHWLsNEP4Vm4RxyT08Nu5xe6d7Kd
PbhYIX94QZMFrcS5xA5adflhZE5MpoivhHPFXts7EbOM7j/eFPsBqWwMQxYkeU+V
enJcQ1Y6PHVHoxEYXwFmG5Zp2TLhEcTutLVmmgEz/IwiWoWhmHtzXjEKKqnjq6aE
93Zssf3VHrxd4DUIr21ER65HJqBk+rfTaVxWes/5Q6CAcnm3M7R8l+e3kdaSKFgl
InautLYWAHYXM57b6+rDwSV40m4Kx/JhTfvIFLLcNO8GP7fOPhQEW7Jant3u5SZ5
lWWrQtotB5lxnkxqKg/gfepevyzTK6c0pkj/uZlHyRo+eOH4+G6hcPCUxsil5v10
KS6+zM9yk82hZy3Kfz9gvjOA0a38Zbh8j2RGQS0dE/Yl8yNUp5bORrcyzz8gtyDb
6+zldy4Ki7t8kbRfOzowMKXbW2X4xgpgsQajKLCbhaqpwF0faFbeRs3K+xTWRUwN
zBGx43qypaYY3Xf/bj7DKP4+ubZGdCIhiaDmVRCCtPxeVf0gCVXs3nALLyiQHZcG
9MBjMll01Yz/I2h+sYT/2YN8/Ju8qO68wGLh9ity1QoLJbECDzflP8PvOTHopuiH
zFOtKhDLs6QM2MVDzk6YmDLGUw9aYkGT7lka87T2Ypx3N5yGaGZFL667Chw6cTnh
TLuN18evAVzo/sndrl4HXqXElroD+wdHAWrJptH+G/O7wW/hfPycH1osdDcxieKa
HIOYR7A64ILd0/j6cvSOELzjAkjVPyXe7gS0Az7duMMbf9eE8lx9ovpVI/Dei3Ye
9HSuGHY+pUcVJkmi6DK2+mpf482EspDm+JupgOJee7hWoBZR4ImNheyoxbTI2GhW
1Bj23nPUW32AodZodfPsTgN2Y4Rgm2JJDOYggAjjT/jrVPwmAapNLLDKntlBJcpJ
kZtHKomlpnIPw0MKaHalxACMHGXhf//nlKVrJC8vVYWVC7+FS6ConRKyLkgg/1ET
u3sbM0/CQcILNFAJfJb6dJJF2G7ZSxvpHx14S71eaB/LGGGTkwvykfEetGjimnjY
ogvdWUSHrPtf3ehXWaMwC/gUAb4rXoMOlI3nhTQclmW08VazDza3OwpaYuAV/65D
6i6JgNMPPs7SvKswdbUfGJF/pDzgZ9VYywl8mwym446JAJZI2m0/jGzXs8v/zsYN
I43hyA8NRPLS7zyabqa5y1Aon2BDSTgAA2B8FJ/I5Fyc3KKWoWqlXnHPHaknflqH
vK05wNYS+17FSDuv7ypjhmE3qO91bOIBxWkEIJuUbT+aniTbJZPcr5zKR0mEZavO
5AF9sP2LWISorH/pF04XYa5kxPJbypaLIG66e7dsv4MNv1E+iNruIyJ/qSQ4Fvvn
lAZ6hlundHsYJex7siVXwik+iDbLB8WpvbCn10z/MhkjfkEmrb457iCC2PBVoL2b
4kvLPF4+sR1iv1msgsW+vn4X/1OolyXEZTD2Gcot+Ebjc8jyxymoEoAROTke059L
H34gWlnnZ7lCbzOfEBN6E4seCo873ykaO9Bn5hm4lFDwZt2wLMqR0ygmtlWFKKJK
WCN9GugAkbdw/JPu/8iYj8sg7Uba1+UVxpFTWFF+YxU6A1S38fIFBfrjt93aoDpt
0EvyMucFQ7pYfadEYPjAGMxjbgAVBAtwNjfuZeTQBpiPx3MzPlOP3QPgsgXYK9Gg
Rs0/OlFSPiBTFopdsj3tkWA1Dqnm5737Tga6MBVvQGwx0XUPaUTh8J1RFcsEEFW4
hg7Z63O5N+p1XgMWDr2jdzKFn0p9eMOAsEEjDrjTop9NsxVft1MFHy0l4vgd+ylq
0tAdyiXQT7TRWgCvqWcVCcu/yuPFqWlRL82WkJzx2CbiUkpN6mTbRPR4zJTYnVhp
QmVkFmtaLx9Emwk9MlOF1GcRpRyN7glRDvvR1wKWvLQkUdM9waONiJOW5NKv4mDG
zTMxwZewOyDhhMTM57BiG9rIv853lx8/mlr4GIiMOt1cdALyba0mcg5wgPT++gCc
nVJz136nfeMuI661AgdZwF0ZoCg3KjlVF5Vlsmz7s88z72xB6HnDDPlF5j9AYeAu
euTExWz/ijQdAGzJKQieioScvimy1IO9Hk9+dKD+EEdl/TtNrnHdlD1iD+vMYu06
a+IIOaI/QlxsSSU9VWTJ/CzCFuGHVSg7LSaW+rXl6GIRluSVdFgt1yhPHTrKH/Df
k6LggE2/lVmmfpbAEybEZhb2SinlEAiC112yaZU1DgE1v46al+iXXF+lHNHK95se
Qt3wR6EH77VwVh4aOFGtfO9YO3o7Slx74A5oLCB2UyYjDssoEZ/1cvsiN51U2vmt
/YSxZTGEfkUY8TW8IMZGXAZzfqEqJ+xlFE1eDFflmZnSYRtkTZabbMQRVL1IbDK5
LsccCypL6mE4UGH9Lu4ycTGb2OLYQj3Rh08LlnEDynunsdhrQADV/TP9ACwjFl3M
UnAOI0vYgl6/VRlu/zJ8ubZRnAYUyffF9z5D6XKwSJH+vRk8RNc7lxT1rSn0lZLa
s/DvTHN+aGB9y7WL4y8RFnRbDl11git5Z7qBsMHkXOmig+cY+6iCxB1uMIEVgl0P
tPtRE6kYeJ5mjBtLGxz1FNJtGQWTeUm9B395huKHOEWajvudawAJHO/HvU7c4+hj
8bRsSP9b8zTX5bkKj6K0ADqkLlusEXaHTuTgXRMJo8NbNKV+4QWOK80nnGAPASHK
dqVNCVE1I0wo84DKyfk2xC4HEAHxnafV6PluXwZBvyeYIjk3KY+2gSR9aFvIrgRm
EPqhVDf6FE32b0P3dxhSVgcZcI3al8L3Y7z2P0JTU71XkEuXpST/HiEvWn6YiCv0
gddf7LT9SfmLFZ7Dp12RRhqdIrCeWvxN9w+SCw72T3uYEgmoFcrYXdaXJkn3f9Dr
1XDOdekDfl9Z6BlEFoD8b+iBO+l/3YC9GWCUYt/wtnJP0j2jmWWnPj6hJvuG3w1+
PwjYgvgHo/yod+0LeC/1IXGpF8DuJzoxjSuqr0AWYRoMAmwxiSWzwrUWlLAl7gix
4GNE/U9K3n76iZT8SjVraRvzZMDqdIlrfnCrUe0UBAyMNaROa1vBqPl28FONZOdU
2Hc3SnuwKvhrxAJha90fiXyUhws8vLomflOngFWwQUoRpobITuQ60MJpHoYAHGGo
BW0j4hIbyjH5YADITdgMlzWe5VygMFBjVmvTpTZu7R5KBy6FcQVCsR9KJuijA9j/
YoslVJM6/isdWennKo6QJMiRvZS2+1NeDg/7CaRHkBeAuo7ML7rzE7DS60DpnOQ6
vEqkASo6/ch2tC48mkxm/v1Q7QLBLQ0Y4rPeY5ENqnqBa2UAzZieGEbKzmzIiBl6
5WilxpmlHQIdsye3KtwifZftgPv/UUCwzvcr8OPcLKHg0ds5ijHmJ8USwemXhfGQ
TTxVe25IK/VRcPlXfcXtrkYhxWd39hA/MTC+re8K53r0G/oeJFT2Plx0ETK/IvwU
KDDy1BgwtKvzbZjJyykbsRRkxDd9US6fdUclhWQc/HHXQBkDarfOmmgOiGKKeCLA
vxXtXOjn1tBVpf6sNQx4P6e8MM+5bNG8OCVC/3+hKApD6yAelBgHaxk4tYQJd1eW
irBxA/6uOAxNFBKK+tGoKSxIEr2bSDJGW2Y/Minx461bnBxW47B/H0zOi1zOnuKy
3FR4cuvwNmuZt6XupXEMXyooztwbzB3uWcDJgWog9hhOp4qvjpvshfkugWtca5lc
yTASZonc548Hd6WZhg5xJzYzFdg0chzQz37CAk0bQv38btwjSSaakBCku+GL7SQD
x9QwO58XnZhX0VUJ7JvAyvuby0llrAu626YAMTq1i0T2EqQPQNj2exJXOoMHR8Fn
/oJtfblKB+uCvL3QOv1buoBvdi5odis6yYBm9Ldu0HLqC7tBF+nWyIz9AeO5apm3
Q5wFag6S46hXNaNBWO8xcWFp3XMUKKcAXjCZcOhGYIEWltS3PoHcJlKxdaLgIES6
p/bnNYbyBWouohSLc93/USn1Wy7echa4mM6Baa0LS1UgBvEvNjgqNX+M9qUTAXeJ
OHzsFv0arVJFzTyg0nRs5faxMKSsTwchyO8WWL3b9+mq0608OmR66KjAsDsncvUk
4CTxU5H2o6cUC/FJ0UT7nvMpojiXmTM3Bjvn7+sp6ZVmDn5Fwgjl3ABTR8sF4n/0
+Blg+LKeE7Dj4I4DHvwhUdObb6UDdFvsxEdsfmltiNomqyLF9PIFlcfnOngm4etd
qcQdEH5g3FVr+JAhWEHNbgTiaz3NV2ajMrRdryzh3SJINcBvHi8hgTwwm3/kA16w
+bzx+jSnxLag0Xi29/rhp9vxu7r8NXEVV+HTVbKPIibTCNNPLvAeeKnMGdLZMVj3
rZC/srkRagGI7TskGUGYPDDpdMct1djfooe7WhcoU75MJzh4kXR10jJE+JolJrzP
TQNOv0PuelD1Hs+c3OROs/HQNBD5KX0pyWc7oKaPGTCSFgePqURJABYbGSG6xkdl
hWU873xGlAYLhPozs+OG4GUScRpRIHWz5mAWcN51XC08MDRvy/FUPD8ZqfmWUXl8
ToZ0Auu+YB+xodZ1L3shK0KO+2FNMKpyW7Ij24+uYsw1wNgUDnqqnKYnB3fxOMsk
seybegdlAVTu9MyYeUOi01MwXMo3L4O/GBnLWEiU0Agipvspzb8mVyAK63oy5kB7
W8MMzCZrCEVRXvB38NGmmhrfyC5/XYg+D2Ax4H1B99NyyrlyEIGD2m9afq1MUr2p
gbLt5spg7osXENkBu++f59wATBQKvpY+BuOOPX4jIJniSrAaCp+Lp4+rKrv5EVg8
JBJapbgsPe9qVME29/RNxy0jK73WykxMB4FuH3DYQ3EwfKmYhJs8fQOpo+5A8mwr
HUOrYehb/L+AWuO2xnqAqy9FQN+poY3Ggx6yxBH3ytVVJsZ1sVbyBM7brohWEtMa
7BoskP5K7Nm2/Se0K/ZXBoaypv1UxlvhVWFz0rrfAWuCRgG+34VT2O0RU/9wQlnJ
psT29agY3JI6LwLrCqf+R28DCrKA6yPQzuYf1LUCgOVv73bSU3AmKxM09/jH6yUP
a7gx8REZPPQUxk7/vCmpMo24fUuqmqPnsm76pkMVRSJUsFzsKpCEASIKFVKNIm8z
x9WuZhqm+u8xKEmX74Zw4vsdkbdX24p1Jg0+8OmRmyHCbVQA/wv2thqdyP/BLKzG
KJ3um4vxhcepBDcp7wuBbfXbvRrFdcYulGgG2bFJ3Ok1Z0jM4PBJNcgLoKImRo6A
6FE4cFIx2QkSGtM8k0PUxs1RXkFF/uhw95r1/mocJvCHPPER3MgUVuoeITuf7AxS
4fK9aE7vO9VD/puueRW6iL4SIt58zi1vVGPnIohQpQ1fovCWCcXNwuo2UG6BvWCf
LCQP2bVRZiscYo1T5GHBob+cvvltKASnHzEvEiO1Z3RwhscS7q+ZQpqSJV6Wrqfl
0dmVh2g1Efn7U1qb4W+HjQU8GCPtB1Jh9Gwu1GUm7r4XGt+jBDjN2384RFBAuiZf
uIRij0nxhzNX6otdd1WIZ59ejmKFqp8lWaCUq7YpMTRNjOk4gRWSX/zVLF8zgL4w
JrlKetNII62OUWSoUm0jJMa5QvITFfyidz4UUg+di6dGDMyZWUc2JP5C1vjTUNSH
9Snmx73ZBiA9e3gaalukabRZLGFY+y7DI64RN3I/fK1ow8XFj2FexcLsyxGkZTCN
L+dgvPJDLai314O2rqGo3JBfhca9YRcOrPCb/MU7dKZ7vT98fs5dOTALbvemVVmA
LQ+nfsrKMZctl02lHEmzuzwU6PWXYUCh08WHqvv5npMHTCrn6MdJpkqMiA9ZkxIh
0N62kDIE18w0o0DxOxrObQDGB3UYo6ii8jgfmRUywNYUisXl/hMm6mhNYpQBiZSH
zbUfZQoniAVjptI6/zBs6sganPlZLwA6y7Z5kgEd+4NzMUfkfnQ0NPef96gtZ32a
EgFsJSaZ4MF4p6PbYC1KlOJEVam9WkJHQnrWf+eljnNEmfCf4n1US6gGJ4VEuYZl
spfEMIdI5M3l7vhCAJw6cTkaeDUhQiML1gmiOzIDIZR4vihR82PXF2qwAu2E6LTO
QGVu9j1HHvZOnDLv6uW4Y79DTpVCHoTf9MhesLc/Burhk4/tyearSPZoRwQCc/2X
aIkSPrQTzflFxy5RPY3wCoixRdkykZiMf7KneYZVHR23oGWaiAYjgrVfKB45k+if
NkeCuKwnE7xDxndk+96w77kF7iwolOvsjgV5R9zaNS02cIZTuiperIDdgcpfvw6z
7uE6EWuF4NgndcXiMldOHkg9vEl4l7GR4uiPksZjW7xwwrOTz4eq1yyfdOPzwTVg
Le1acEgg5MF6VoYoGF3eKvdHBTPeHPum0S9gRAhtYb2evGojisMl3wB0LFsHLs/b
PS/4BKzbNCpqwnZGsi3r+YeSp4afztYXmdc6zogVPiLc9sXK+Rjwa1o0ZraPb3bQ
Ch9TLFQzx2q7O6yEXCaek5YOHRExlet6iPadp0GiQ8uREkgVWodDhar3JE53CwMZ
s05IY4BBKAx0U+TVwK1enDVCITQudFCHu8e9DUpEjesLI/y6GS+Yx+KpJ6lCq+II
nljIr+7/9e0GscsGD1q7ZteugN97XdFIUjVXOBxkGRq+bF6mYQ1iIj4oa6oOUq+t
d1Wv7f8SZVhlUVGR/CKto5Jh+ZIDOA9PC51l1MmsOVn1nhR7aOeh8BtAY3xQYPVc
zRIYeIwTtHpD3+VB0XAphW0o1vxbhXPTXZClm/aKO7TykGj6DJT4Yal2+NF9WPbC
+NSPyziTIGvB7PEs7QNh/IMYkbpuCMUama7MrKY5QLCtmPO5igIQvgUpoRTOH/hq
IJb2i3tZHPP7jYye9GeD2q9XvVtrRjHoBhknQB/KJ8bjoA2f5cRF51U6Ho+6vaKa
11dPrDVKV9h1/elphDbBPJiPoSmwMwRJemm4e05lYu1JVLSx3aWo/AGyGMH7hTSv
6BrHj2xIR53DA+rAOpPtgawzUCUFLD+Xh6sMXC6fapVm2xdnta1Fp+Sq6rWa0MZz
6OvJ55Va3OhRTXfhWqaoCaKMasujcqptSe8vUSLeALRZS6DWVb9N9tC+3iP0Z526
y7EAgKqxI15kA0LjNrvzjqWdTrh5Xqs2rUww3G/W4Uffz3MDoPkHmfrQJHmtvVPd
y64rnaJBQzEiHUbjQbJcl9T6tESw18CtdPRiaQENajIWGLJ67g96zyJ/7G86UbHc
PY9fphmMHVDBa3zfsLDLOH1RK1X3P+rjfmM17New6sgWZR0tZTY9XneIWhGiMfG/
vc03G8xh6J39uB51AULXnofrX0u6W3tvSfM3UT/x4ouJnbYtKimGnuD79ygmMrCf
BuFNV7iGXCXGKzCErju4abeUdZJH21DpC1diNJzKKlFUTMcwoOyh5Srik+HtF+yg
6s+dQPbTmdorxSil4kMUhh3o44FFjpL+wt3T4X7ufOQGRG1ySCufwUoWq1IC3BGQ
wegUioepuK4gvJ6oeG1l2BFsCOkoq5jePoUAe0wefDLATGNSqO85Gy9Y1IQLIAHH
9aa18kPbWtNTX12eGKrMhT9h99OTLQxp4vnN1uRGYFpHaiLh0iLukw/GQkva6c77
Z1swdUHlW2OPmOI1yks+KEZe0VV9whJvG6N3np8TIqyooTOEtw3q1oDwvw3WRMzP
lyd5cOR/HNJH5W4dcmF9wOf25gSNmm9dNGS4/LFpMu+tUZvCMHDGKRj2w1YMxZmZ
46fgmS2CsQWPwbuDc6+zaw0/Q7kowJDAlkbW/TEP0pEyMhWJXVvewzpckx+3S/bj
ZrcZ8dUQKGZjbIMf+BRuZsXqntsz98FUYaOHke7Qdj43Qeie3OgH/Rm99kpvYUAu
J4mEtd+i+kLIifJTlKKYgHOwn92QW5hpAbrLAavi82kKbVZ+RN0uL39Fy1E1y+gn
3huYHI0HkXrzVWxTDjQORKZoDt1mEmxBTdMSu79Ei5bK4wxsku3mW1hgryQsfM6E
1yb36FMqj3tFnSmK/Q6IVLI3Z/RlsAEeVXsD6ZoPl0c2AdO8XD+Hi3uVkoIvFV9C
0ywpI/UEMOUZtZWqbNEJnQfUGjkPTjWJ6hymEBc/RDHb6e9EG1dOID5vwUG1lFTI
kG4jyKzVF4cp+YszyjzuKtfsO3NSQjlsnJ7UHwREFOwsllouGfNrogC98vA9cPgE
lMi9NqmnApg+O70tvQlem8p6LrGvWjZyynWpg8aIdLeAq0en5dqWivU210NqokVF
AlNECYXYlql1pBE52A4XAB5NjfPhK7nkBzfEOJKj8Js2mkkonEpEr7wW0faPAVNm
d/nHPwwCtVDEqg3o4UKlJKYf/VhQDZ0N149WmH4iSAqyr6hiRZL6uUaWbIt4dgM3
NhPnACGvwo3brzm6FNUm/njAcQW4rUNepJe2XrKroe8PO1bjtUqucIntY3L2i6MI
6dtJTEsIrRXHiH5yAkJFGscRyEmj50oiaC2U7Dy6swPiXgRtDiPXDtuYULj95mB4
aZ1n1F19YGOodmmqiS/KYTRh2TkPfINn1qJdUZ9ukA8RpfRxnMT//MT6RIE+Bhab
QHR3KXY8npOguGzEkY/n4AWjgZev051kx+D6nC9mDgogrdyXvOY3keNt3D21awY9
2xYjI/oy41nss0Z5NoOovHabPy8ExdA6cIM1xrzrJEkzetX6hy+EY3jeepaicc+6
tihOth1Ol1Vp+gQQ2Bl9nKE6rq3qz1/zFnGgGz+iyoqK4AJ8ChcAgCuVh1pvXVFB
6DQ5PJOgiy23sgPGjncFvf9EnOk5K0XCxR0rziCREqhXJZS6OGDUJOl8IyXabIRw
9y0H4Yx2vlvcB45y+Bh0+SDJt6SUUg1bM0E8aEH6jvarZP3r78rOfC1Ui4fcKp/Y
lko4ab7IWr8Dz5ZmVCi9xJCXC1vkB9KHMB1/HdSqg1bt6r590HEN3oLsCgf7ylyE
cSXndinY/pwWDoP8XtZtr7Hj21SylGs2M8MA5/SBZnrhbyUOYo4airmiVaGSAqMa
Ib7l3MEVDS1qn837a/6nv4ElBQVJWh7YqygCIjb+QG7k4I7n5oKTfKLLU98cDKcT
waNDINAVbbxb415uiPXrSC3AGWBDftZD6kmG79KuMwxZf10kB5swl9HEyIGSR4mw
BcGxlmDQCiV/YqdvKjvJsmM9mFZkrT8ThqHO39cclO+FFzG07RDg76lfbOliuKE9
raHBhacIzcOVjePbl66ZqgCOPDHcsbf1cNosVfJZ6hDt8A6JkwqiWGCyZeFTYUhq
0xDgsUJRnyBUsIut0kvkQibQjlX6r8dcPfv06E4DONSJFau9JCpqtHirj21MmB4/
8mkESLGmqYi+WFc8uXBtgrrnBli9MHMO4VBtW2UA5atuXVU0fDF4Plzeu+z9rhCa
XC3VDYzLDCOb+1PqUH7lpywfvPFYZTvzAtPygFKJa7zymh80rOpwla9a6ipO6zPM
HnWlqJkzrCuFMpuXxMuMa3Ls4nwTFvm7jEcfJXbXey6ONO9QlNoD6Y8og5sJhOiP
qQz/VG4K5wT33ZLq6bLGv3Gt+UPxcpf67nu9eSlGwC85T1tknoizXSDiqqMsIrGS
3L9Rad9ND+BmzFhcDLEoryatEegrAoHxZeOF1EtTpkzQiQUz/tZ5mm/puVyccrY7
wCkeGb4imRpKoelXoX9/nvwhGTH7WZzecLb+a8l+AEJmngq++rXxQ6jBYrtUnfFP
hH5Nxlkza3c2H8zszPDzkwAM2y8ohsNuARBXtobWYo/R+3RhYb4o9yltbnKw7hng
QOus6qYk24+k9C0PdNTi/cUJpJ8TDAe4Z20ee8lNs+NiKBNC9FxFKwHGlA03RpPK
iUsDW5k2zamotG0W9D6bnNv7+h313oa6e32Jn/6THujeoQK8Suu/s+tNGYtYgnTC
+QYtyK+060JPRa3zPSMYXALWUFiiwuqr+eebrYx8uYqkir+cAN6kVTKqFoHo+Kzp
Ag7iOIN2S6oYSp4MsVrpZUmp5ozKLhxBuj5w6c6uqn8+2UamyfFhTBNcEkn7SCoG
LC0eB0BLZps3LqJXC5vrsMato7PS9WuPFTs2ih5d4qr3pns/VwthummE7QrLz02q
+fyx/BN0I5VvJO0oKvPk/JRfWus5SbIaV5+xwiN/0U035YHo02Tw7pW8O0zeUefT
Fg7yP5iYGCJSc7POBYLNStxxqmvnpl2v0NkArAns5draNgQlUCsfWB+1Kkn1csFK
QChvD4T0Ee6hFmgGrHJV4Nwn+Cap4PDGUEOSOXFO1wjcG3nPhPhfGtahyONO/kIY
tjouphwagUqan4zUuRfZURCmevJwUJLsN+g1TiuGN/gD0iay4Difert1dhkz8lT3
J1EWGmjCr0qcmCkiKs1TRdeYTdkvaiziK0EjN5prFVTmPD5cQCcHYO5a+DcagCEE
hyXnGO4kxzUjMILHlP9zu4AeGzaKmOsCC3cOKRthqJff402ZpPeH6ndcwfaSIITO
oJTur7ywH3qEkVe53MrfFPYVUSynsM4MgSrfzpcM0elyJKg6ch+dadYlRB0yaLPR
9Ym3oIrvBbNTfvWHz/eFXJWZZ3XyjgG6q6Et+taVp60a6Bqx91hQT4Fop0cGr7d4
MScYdGKS84U6KLVNcUEFsz4CDamoR31enwj0kAk0xssxdjz+pyy27EzSPleU1LVv
hLREoLSrYuCrjsLsaEtJqdgfyO39xvygG2vdr1l1Kz+biQVXD5m4SRKNwRS9NkSt
Zv3HBDGCx+Dezs1gqeScV8rvXmZiGFj6Kofa7oYSpUTf0F92FccSpbWCb3yIxWia
lAu1P2PmcHuhJ+qdsYhhW5vA4C3y9tBJyZQgH0eVJ5GfmSAdiX/EQCHHTmzYRe9c
eP375gj/sEAPCNaQcFJApYGdzHpbXankowBqOSALVz+T6u8SdBJbHOH95sEEAgBI
mdStAAiCdEKiKssQnMC1NQdX+pB2L8we2tUhJ+E27bx23Eks069ACdGSC71vmXOJ
jS/NsQvfKRJvOGst340/TmG8WptdHxP6JeWEifJHLsHtfRrjYs3RpAOHyd9vX2gC
5U1tpkRLaLs/WqoGTl2AiIUW80nOrIcTwMDSml1v6f8GWziD/gvdLRiS5UaOGaZb
eQ6c67tPtCZWHsJWsjuq1PdxyUD9uSgaMn4zm901xJQ7VKf1tXC60GOkw32Nw8D5
jrsgPkdVngMUzBG0gkvLGohD+0KbACNhMMvCek5xVPKw62C36OoPue4/fU2HHa7h
97Lb/J28/5JDw/Fg5aY3upecEPJnRqtgD5XIpt/L95fxq4fL/FfuLvTl7zzbnWvw
5XkJ3UnYfAEvZK9urQKvBX1buUUQxfI9GuLh6Lv5OLzh6qMAZeMgvGg1sHKz2KCQ
403ukZpuW562NaifL7bj1LVQImCsSQ1x3W4hYJd9jQvyHklLBqfZERHEE0aXbb6E
Jpq1K+gIeCr776U6BjM81s6PJNX8xPTiBEDrDH2Bdgvc4E52qQPZ62Yu3miVYv+X
K8NRNT0N7hC/p0qGApyoUzzG/1rhpp6576d0lyD3wGZnlLcVbTkrfeXo9WhMWi+X
620T7fObAPN2Ub0Rr9xVkjuGEgRcSuHxEvlH3ur4D05BPHewyEzK1Nxt/mRjsR6r
VEmdzpMwEphhbxrWeFz25VXDhZtaM1QsrC8Q5inACQYAYcOqZDOP2Mt43ICHgqLw
6SrqW3X59R+eboe5XO86Q7jel0yfLxixZm+7U09vbqEIMDq+hGxSuan78qAZoO1M
KXc9QVODKogZQwrHEhi4DMIfEbp0x13wQmqjAspavcStaq3jbrpGQAOYBA0McqaK
MzUYhlRovYJ2XtiO/MDq/OFLUyoGVfYfF+aFdDBs5L0Y+sRKZB+iYzsTKDmq7ET5
PhQG29TUH2hsJU49veQ37LbLm2PTLAMbji17TYvxWGn3R/m/xXGTotrT7Ksk30rL
3Zzd0Y42xa72YeukyHVO1wjVQRSHf75q9Ld2Yphq/Z4BlCUX2BkIYfr9fJJoHqLX
CTDlBZZZCZwaKivy8Bk3cgTdTUHzSplMbMTjsQGaWdT9ImmS2f74CMtUqm4OYJ7D
37Wy4YiL8h2JYtEmfXrs1YVdckZC6XNUOECASIRXo6lPtgT3H+2APooIX0DOT0HD
5GOzsqm/AIvv8hPGA3QlA1EGX1Sl5f6jZSAt44u6k7nW+p2xuLvHI/lXHiQlpbFj
aAry3zoDET0cZlBniVF9BILNofBLR4OYVJvGGwwBIK2cU6CSBkj43g7Eee4TZmrk
1PLgcbyEW14emRcsNRTo0Os7vnSjmUAPiEekdXCx5CXrozuUOOFTDuoGchPmAdTp
3DFOYaosFNj9ReQzpUrjbeYRQRAXmh2p9J3Yrgl9KgBiNo9cW8EFIfbiZKeeqW9D
tBjpgjDH6WCf1+hL/YTAvQ==
`protect end_protected