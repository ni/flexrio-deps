`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24384 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzowYN4Gvm9xQvwMwZ34lM6H5hMwl0KNDDyvyI1nwdTjp
Al7axkYtXA3Bhc1GIWgxuLR0j87lYXDxgeZVzJixaDDa+yp5NU97CytpT4xHwoIY
YzSKE1b1R+sZutITit4vWSZI+rznlrfHJv6FNxVvwhMelP3LTA5hqZWchSPhGDst
swk6jykIH+L0UHDwTv6sqpQmrqvt2q79i3tdFGi8jx9g8jCNz9Fzd30tNsbVYkX5
WlY7DdFYVZpxolXwyXVV+MzUN0dxT8PZND1cJd/O9P037HI+M2nY5WYm7T5ylE9u
uv6DCp7yaUIp1dsNmdIFTjO1fPPf4YdWtPvQy12TFk2xp/Tq8F6YTHD5MgxMuVJC
jfKKv2zWSwFym+cMPSRfhU2u0OuA4WBZdGMKymqwbGAMWgKexFR+xe7Nx/FWMAqd
Y85v0g/LdZoN8tJnnIMZwakrzp3QpQNSJvZEcmppkP01Zg8D0xUzRssYKoiaPn+f
NTiNaTxART/VUUfZzIa9bEIbBh7N/LETCeAdQLRjyIOFSdg6Eq2Qz5CnUQESsF9s
rFkEjzQo8nRyYK/uFduXrHhK4li+4ZaZsp/Y2nktYC8RW6a+y5ROgvlKtvBMvdUz
A17REbiYyofYQgzwYzUQsU71MgKeRTpH39iSvFWm7DH0Cv2Wyo/8vnBlsowJqBsD
ZxvmA8KASCdCZEgSRn86nf/mtuc7yJx2jZwm9xLUeo5JtUy67ehc0mm8kpNunwyr
A+hhDysGP52O2iFqE2K/2Ubf6KKN2c5UYssRkx1gnial6aqI8v5BVrIUriCfi+07
mTbbT2t71Ml4Bcc2+tWbBlYP9J7sJ26V/NS4LtoIQYhBoH8pUWPrFMaREgWKmyWi
RxK5mdHVN3q0ojKUMYjKP1/TqFwS0b+7bRGDPJMgptlUYOSqC1NtrX2XdAY46TS9
gN07IdQH+keHIMrNkDz+kFTZxICQp/49IUnYQkYdWvzd22XFSa1E+mEOjrJhID7u
H9BQGqUuQktGFNQ7hKi/5jPSTygag4+HNXQlyrEaHAHjeFQ6CabFp009wh/jQC5R
AejNJZk9KeWqCbrZyqzjmgOOO5YzjVz6LtaKXIgCDFraUMJ5LyGH7XbiC9+/2pka
8Su5GfaKRdmomI40RlIp6JlnlOHo/l3ROcHAT46CIbbWscB46rfvyFTnh8g3x2Kg
pyrkoPEV/lwgU9B0TkC0HPuEyqvKWGKUi1h8jzmmfShvx4/g/w45b74kZ9lwdS3z
PfY7mQHAv92x+QDr0zHZrhFqU3SJyal5ZmaltVAM1VYOL7rhQrGVUz6qCalXeV+v
5XM3/4zYHRJTsMbb8r9KlLkogT68kfbR8H5+m2+wkQwjLsEAJQuM2jWZb3Jj7yjj
Chx4I6GJuzuEzrBEF2iTL1EnYCYUrokQ3Hlc8Js4M94jN58laZ7zcLJ7RW57QAZp
f4UIJYB4/R90puI/apZcrjQVX7+1S2sFZBHj4v9ZfjmjXPDc7p0htpFwhdRoRtPh
DaNpXnU/ijOqdjY808u26OxkbHRg4TS28RNW2A1z3K/wS28quB805P8MQTJ5A3Vv
mPLCd4jP5I/4BYQF1zhZtbDRnKHzARE6FVrIE/Zk2/H0rLQ/tOBoE1NRKzGBAvnr
T+tEDr+Qy2sJtvSbkcf+df+cXNiMJ8BkIF5X7Sok+aDqMl8fz1Sz6wMTzYYqADQE
QXpIvuusu9+j3JOUisarrBbJgTaxBnzusNkXNaVBQEa5hH4XSgoWgnXNRGZMdaej
n4K17CW6/yhUr+WGOeMWuxXL2vdfx29tjJMkhn3OhPCUP4HeKD7R6hz0oGT7LcMa
9HSnTllV+M08r2i+82uK9wA+nZWLNaAz0LfpIoJf9R1oZqRsnLaeGsjoUEkthFcW
7obb/mSNGrOQUK78EeIJ6ovjzUjucOxEowjNCnXuyzz4m1nnJE8Gy5VxoOlk08Fp
dbvnf8ciu9m/DzrYfBK50Ol3HyKr4rpy+TCSHHjhFUU1/3tM/m/rgSZw1Pe187sA
zL3LsQ54Q/sgHf97OAFycyNtehvuwIuFyIRZGPC5oOxcIkAsc5PmqJXrVhWciUbv
yDRZrz00zmOAQMtmvkrB8j+eFxGpLFiweNwvBLlLJGXcVFlGWBhL+UOMkIOzC+qi
JzMZyJo568UtjUsW30l22mForZ8DVi+cXjar/f1a6huL5XZvqKm6ePAch0U7IqhC
ciE/fu8jLBFFc2JeAcZBOpb2sJ7yrHvjxBovsDUkxnyuQFxHExY6vw488P5TCeu5
tbJHCRPttH9OCZAGDWIZYIeCpxcS4C8tkgRKcx6eqSCf4gjc2C1+5CIE2LJHK63e
LbVHOKVk6pDBzksuP2eIBzAy0g4IWmSiTzc8SKBporo+P2kpX9r5TGpsZ+rxCQPU
jxmwDyevs6Pm+ROF2ACfNXQ7XfaALE/NuRlBgPdcMRD4rbVzZnczIYOACbPRG520
YYX5gCvBg76Nn74qTnobaghuthCpStGjwjVMJ+bpiK8LKFs4TG7ef3UBaPWDtgC0
4lmHTDVpSUSgjTuQ+knNSWOQeJXC6GeHGXGuOtuO8VUn3cEkuUODnBgDRKCH2OL+
VlZ/suPODMr/RmY17DvJcMe6O5tjq2F9P7TiKxRj4y4c5+O5+zGk3XLlUhwkqnzq
fxqp0OaxwRZFFIx3aED0L6ScLUicZmNDseZbb7wMOff7joCqmtCnRMisDKIj3sI4
XWNeDJ/f/excgHkUSyqSJzSsDiTGlejGwQOdf0H2bASoyGff4I53dR/Ewobc5CM2
YoAB8Ha4Ek4ESwMR04NGajw4pH7oQbd4n/Sx61nCLzJaHzmWbMDEYOVp+cH5SHXb
QFEKlgVsayBE+YNCOUvvTJNnM80SWT0+FEZrYEyvYU2Soq57SUvOoETWTp14sO6E
asu0rQzXpsuAvw/qjPk0yrW5o/G4QLptkQUSrD40DBjmvLBuhyoWomLSUEbgMHWQ
f8Ynfnp8KKpWmh76hy7VSyHPGsXcpdicjcP98HxhJo32EgtyoD7v4Eud019jhSnb
LtEZHSlkSFrxlVFAbk5cAE5nPhQZ10qZjtiJzegjhc74Ih9fO+lpgWfD8N5bVKs/
o3urgzf0xp9r4ZGIesT2ktvfDuYaJfQRik11K+2N6XAFI1Uwejn46cYZLqw6nZqH
CUu70Cgz/lUXywZevGVbfbVPDbQpuQn5NxDcyDk6EB0LnkpM5P3zu1p9/N1UyPEW
59ZN0Q4KpTPYN6jxD+u+5wawjbJN7i4hzinjDoIQFzExLX0/9VtKXVkmr2JAJXSb
x6We1tbrgozLtMjqxfsfn1sntN5cIQ0uxU53wLzZNu8INQNXCHxDFxWQuvTRixLH
czf4tm3cPCBPozw40YaJxGXyHiwhk91iUwZVkAOo7XSh4lKMREFl1EJhviW4l7S1
UnFGK26nSIcpr9D9x/+gwHv4Oe5YGNCt2DZ+pshGVoT8U5MOA+ONk6eJyBPbbyiR
wnRuMbdwWR+O1++EkGKiNKXD1YI+urImJc0DDg6t9HWsEW42ZjI8FcdCZbLXp+8+
1kLOP8YjC81wzDaEcUEj0m699yxUd5rDeJrpphzJjzsd4DU+VtG2wd0QfdLfJ69N
HmSWyei0d1qJ4B3pZZgN3ZVpZHKRwd6IUC0xBF3P3E5A4yXCei3d70RIWll5guqC
+yJEvV3LaCCmGdFA0zJbe6rpVXPzOX9P2HT/AEbC3JADfqKYul3ZY17HC8P/eiN+
j22jdrw+CA2SC6zIlsk7UEC0UIAZyO6lm8bs6Q9G5jC5qx31R2yG9NKu8AM4+DMD
SriR6q88dwr23/NI2Czi65G+kMBanDTTW7SYMnP29rft5QKWtgVxIGt9mZ0MNwIY
8FiWhr5EHoeupwutieDIIgdoBdz6xRSHsZXVwK58kDm28Y0zikscNjZEZ246NdVP
cr1owZrxn+kCPrYwPUfFHByPBQj0XTonAFY5SYbBNPRRJSsoZMGGcELw7I03DlQt
e2cTOtaSp6CR+hcYQXbcPjTyt2QIelf/Ve+OSRtvb0A7cEmGoM28mA/HiT4mR8EQ
Wzbz0QbBuQHCe/qccd1417TK+qusWTsQp4oTEsPsMGNwbPPuTo4KufOJSg4hojQm
3X/PZW2OXO6U78EoybFNy3TQhlGQxMyc55/2k1Gs+TWQWVqHbDKMeBTxxSHaXJyH
CsXSuv0K6XnZPduWHYrlJ4UB1mxkZ3BO0bPUxj6cvjo2kvolOi5eRRttEG6dUM/g
W9YtOSFIWoeEFYr7M9lW55nTDJnz/y95GinMTiboRrFQQlPsrIsZN4vbkhuyOnXm
Lkf1RN4L3Omjn+MQMxOr3VyTnlaNX9L7IX03x4PMuBj0un+kmJr9C8UZEDY4vNxH
yPRucyoZQDuANdU+z7hFeUryaTMz3hUmyTPDG7wNxljWr/PD9QoGZMZKW74yJwqn
maNIsfFYlsaVF0sN/mYvtCRsVXdARaS1sOJqx/6oWOAGSHvSvJkdcLwI9GvjBlsK
vNNAZfmO3XnadctFlPHRzdP6GgcynzNQTH9om9JULd5mn3GE6Bm2z3jtH6EZ37Yv
41zwHLcyULYi/zfBAtVjkJzU/WR+flR7EX/H56BIrd0yDtZWVGrMXLKn5ERs8yVb
CjxjE65jBtt0CZI/EtrXDcIJYT7lUMRb1UsG8ldGz1EihUlZrkAf80lLCuONT6cS
OTAoa7BsIbFMgvJL+NkUr49xr9hv9PqQBl9F2di3CekSICYzdBqF/bifFlo/It5s
5vsUb1z8ZepLs3eft8h7JHBxMzmcvTWD+eIRINjq8Xi/7Zh57d2mXd7l0olOMsd0
tkqGTAE0zP8ChX9O0Oq44E0Q0+X0zmRU1ca0GwTrP8dcDFqjc3UPSmPlp9mqRL/y
yna/j5lOjWkZsAP4CcssiCW9rMXUoLI5nvKq9p+Ff/Lv6m94nXqNbmw+hXos8dS2
WK+pMdXPB/1Zt+ueKgzdNIFI6SVDfnbeIU6m7Wnk9uk4bWBeYxA7gADRMU2/qO44
LzL1QF9PIH2C8rWa+dH/XBZW7mCEQ1xo6qV57ujgXUcfBbtutwJLb/W5UJiQpJrg
vGKtwEluJP5B2KJvN3hdrSlxMio3PwQ0BWNSjynl4ixpypY64zvCBvhRR5qkLtdl
Q9PO0fVMYKH7Qc/xUHhOem4ulvkn4T/PJaVlrOUkU1h+yfPX/8qCs53x36lymdum
tOTVLIogUb7ujxBfxt037naXH9xg3qWzCm5GjP5Ca2fPjDU/a9UOsTfpWJAW6tUp
F5i2SCp84P7Sg+KCfcGqQU7FMQjH9MmjDbE7et1hrD7iSu+YGqMSGPRwDbb1O9XN
r/vXX1Wruzm2FLi5tXul9xi2hI8Ggjdy676BNMtTRmwMCh7ujKFstH1ONUXOD82N
qEjdXKw20YvmN+h2Oj2UXEXNVw/Uwf+TyRreGMWMtRhZE5ec8PD9P3tk2GZU3Kc5
UsArfUkVo3FCXE89LJlNuCadrm9AOj+LIamabtwf8xpjhhrfW7tcuBtb05xTv0P9
J1PcSFm5Lj2ADWN2Y2soelGorr3w34TocO1JGU6JscWDruF1FyrqJ1DDUUcVRCTB
1XWk9ZEWamQGbZVQyraeKUXI5ku/qkDKpm6yrr2PbL+FyvN1HBV32PDHnjPMJsEn
vqGkAh4fyLPMFkXhNWBYaaeLqa089uGAmEEglPMqY/GLl+CQOES3Ebdh/biuJAGI
PyNIBH6FgULg3QK9xONgPPwqXUIWAqVSh1U1q+Reej+0TIew7H7INnWZ1C3CqyXy
G+5MhxEM2yF+wL6jTG7CM5fZvwEy6PUqqewfzoIXuycKrHAx0ZZQraMiG310Pns8
kFF309JkttqwcSmBQz+KHiZ1zw6FqdQFKl9RflnW+OXOKh35aQkk4YOUnCD3T7DP
TqUsuxi1iER8OEO0JJEWNZxZ41KN378vXDaYruIAmFHYF8qT+FvTd9PQ3inc5OAx
sDbnfUtkoE0bMVofqBHzgA3DbV4MiDcN6NHUxB7ZCHq5XBrfnIfTpOn02XAbzpis
576XfL2GrlEUkzTQcxzKgf8F1A20Hr0WjmE9WZpADoi6xmn08OA0Nah37IbHHwZP
WEO5mpVDJddPaYaQuBOvVltkK2zJWcoZn2BoBi/e2XKsjlELYHdCOrzOom8gDJHO
lEsT3JbvVIS/cqXTX5jvl9PExd8x5l8eMC3V09+RjFY0hz1HldOO+QTMsOSPd+MA
qI+m4QkWBP4bR0WnOD6v/mBMkWjD+GNoSfJVRd54IgAfk3Cee1SNYeP2rh0BjyK3
gdznNmIPXn77C6QCmPR7JvJvrjUUUxAXh1oyBJTNkeU+tQdiZZfcJFljTf7tdgXt
u6PKqUZbYr1h1XLguF2LBDIdFlPGCjalfWQx0+rXS9/QZpjWHjLDH7MXfQ4+cAhD
ke4hF2Rcl8SnjqAU74c+fJYFhVpE9A73Apetzgsvx2reZltRuG9y8erx9fsv1h/r
8oROVVxKEgbWUhqds1OnF5slIItpqn8/bPKYgcbS7x7GuSIuOC/x5TkkAxKdtQis
TGhzNMj5n2GBaZgIVC7AndamnFuSWFMejwBy3D04LUA3KXJb56PWSi0bnya/virJ
SMj4+57fVfD8EWrCetwpx+p56WQInaaHhVRxvw6iumwuXpXurtX3CHZGnvGV+/q5
BNub9aOymmGp5YRMprhkzwepZaLKgrY+o37EZ6B3WWXgnwTtwtDFQFX9CZzyLcFt
Jx563GMGBtrgicfAXC9PRihuQPyszZuBPSUkdzCKOm9txXuysck8BOAJGinfmqfR
lyclHz/mV1bI86GMD9/nJ1m/eF5e8pHMnU2SjQVI4t36LfW5b49bK9WdQ5vbvsng
miqsNkOMFFO/jIVTLysUNWLvv6M7po/LJa1DVtK8ocm7gsYmk5Dt2eBQtKK1yJBr
5UG5a/+1FclntSbi2qbdOfLNHlrDaLccr3Raoey5JJNuXNe5ZRc7YxVL9cmlsJxl
DLKrK/ISI/V+SUsT7MYWWeIRl11K8VPhWGlLGuiDB8P+KRjnBM05b+3YlBvRm+Qh
vKxXXdrAGrIi18t4phHLY54aYJ5qLq+P9cs+YFIhKOE1xjLV5EN1h3U54xiMj1tQ
kaKKNcaL5IedEyv171zUBhph3ZYLnpQaC5bSQnLVqInEWtGh0hl5Gvs2KeV/zeSN
iXYhiteyXYbthSvnRWMzIBlZWj2XM2LSOWfIRMwTKkzVkWkOq54/5H9pt/rC75QD
IgepcIBziJnwwwtlDv20YXpBK4/uDVGRTFmkVBpng2xNTNB+r0BqWtRJFCVgJL+z
f50XYm1oytcbyd0OAKn8vAdLz0Rtz/RdDqmBS8frx6cDCBaf5PcgfhutsjzIE7Ek
UazrD69FkTwNROEf1FlviwfZLTk2oi7rjvaPW1lx/Y5MiaM+9lbisnbbW7G+whnN
v7nFBscvrBNGl4BCWskDfBV0DFcjz03NkJyeS6AuMkWKOa4eg4A/PQBAuR1pA8Rz
RrTFmlfhDWAhMy0HnMAr7jqMlNM9Nnqbz8WcpyPMkia+HkkWbGBsw9uhd01QUgwO
l41ci1hE2ATbStKN5XMpTow0OG0Ity2tgU2R9rpPgxyl9jtHoM+Uu+3SzYAK42FR
h4V5R04ozPrvGiTOa3JIK+3FP9HZ5QX5P5G1RnCa5r0803yTltZskSgeNl3u7Jqc
NpGwbcoTYQ0dwAqJSUPOuAsnkDVvHuPC1P/eD3sBQtr+CZvmUnjJJjssClpSJLxT
YI/LL/s5RV0i8+w/v+PdpGMXOmZ3tRd2tMri3q0xF3zKZpFm1Qv9jbqhgf8a8IqK
/G/7kyp8OmZFM7hj0UCknjjDI5TYxePhXRyYELNNT2X2W+tgABLHx/f9wGQhcmrX
TWOBku0b95nNV7O5/XzLcq6JTqDH57lhW32X40ea9dGyhPA7iaGU4K4fejPVAvnW
Itl0Y8E2vl9VnsMXF9ognYeZbAU3JTXEf31gIi5mZBAE1efmqKDrShkmwUAmse5l
HbHGR44PT4tkV2MYiRClNzwU82ZrdwR2HVjAvZz5fkzspkgjjXPfug7fcPgD162F
FSyelcNUW+RUlHuasWigvJ9FkJV+RA4PDb1MJjD4yEXOt3rTR/HhMi/2DJ8kNCUX
bFSz8769rx985u8QzYRzzidwnM0hTDDaq7R7dOhGWp495TesQjxywSfsXL/vwy4F
EnpHL4V+zpuJljaN5kfs5v3QvDOLVlb/nVAEmR0S5vP/zVEmk9v323XMbBkgCRTn
7+CXljMF1ZgXasgTi8u0WBFSilLPeFWR1DB69sv8e6tPM7rg+P4E3DSj7kCjv/Ze
WMYf5srhOIAdyBVRdb0qk0EOZkdvZ6gjp4PnpUgWAiya5phFcjbRQ3OJl2uZNvUd
waA5pbebECPcL4qwissipbCnj/J+/hpo8pcK8fN+bo80U8ueURPkIcy20A1j3ztY
lX+uejQQqcAnUPbu5bMyDYoMDglQW0JTXCm8N8AieD3u/zfuIGb4csGc6qEzsbTn
e0lpxHNoN5Tid5b3zpQubSCsGb+t7htSCE8TenSwXiFZstAifaWBzoUN8DiwkSDF
rVbyXoacBcLRgDAMMh1S99q1IV2HP6bcjt7hVcEab6qK1MR8q8YukcYfd2RA3yzM
5ZQ9njEr50ipp2CPTOzZ8o5LwN8dqtC2lEcGAvCmtEfFT/JQ2M8QbakHcUMRFTHj
MVBz56dH5kFnHkyd4VukS5TwykNu9ZFOKYlA62r68pg270+qZYhxtYawzljQWk/+
//eo5owJg0eSyTj+j8rU3BV4+I7vfiPDngSSmkOj/PhDAxX9C5uCV53qe0ge1fsB
Zd8E4cjyRcEZo/Lx4GUL77HagSbVj3NYbxGJQUMJpXmzb/TcKu5EVWWD+SWnZDc4
LDYWKNRA/Q4Ce0ETapt93udJUIMnjW6EmGLRG/4hn1cMaKjT8nBkdbqdYrf5Q2XR
WMVX9PirHGyp2H9cnIKTPhWvotHy0eKhXJpxPzxtjNeQAVoIBXuERIG9kUMmK0o7
YcIKmx2OpvR7nciQ+IS0A/HKpgCMdKopj2LcoTxNpZk4X2qct4H9xP2by3ztp7UA
0JcCixYp21O/nUuAAP/xiWtT9iEan2Xdv3Er8BrX/vjI1UzykNamMkJAWN/hYXGE
Se9qZyQ2V7QfeP3zO06gb2zXPLMGa5QRZlygkwROog5+BJQJo1ebCdmLX228/5In
sq3v/H32QDglEMCExh9PeOxEiOtc+7lcqdF7jshN6dB3FDsFE3Uhi0B/5ROlQotf
FUCVdbcvtBRXwaX/Zf8xl8v0AwlcJOsnALoY5xWClK69YS0b/WLBGoLd/3Gh7WLi
zkJz98HTfYWtZQtN944eOv5d/JbGT9mmb7/SaJlYdVYq+SSEhKxrepk/t0RlFckA
KqQr0eSWOe433YNDVNBNGwdTprBYmeMxII/6JvBfYrnJQtc1V5sw7KghxU2xWlRJ
iqbGpvVTZ9lyzzuf3WgnEIb6qJ5bDaaRsPhbH1a82uTftBwnYNR83jWEqWaQd1vV
AbbiuyQvdJFMUx2steIyhsL68Ony4T80xIyMkL5etvsF/oIDM+WLV5g2yjtVmO7U
b6PwW5MwxfceTyxaK7RoG3zTjipJUTjcgdreJpqVc2EvdgS4fQwLmIXYJj1tXkeJ
kd/zgIvINg4j8rspbLP/kaMYLg2hyRg+UENq02k2D7m67qDRXKtWPuRPe1wGbrWv
8Oj+dHgzq48NpwGBu00iXv3Mrp+gmDiJcNiaHsjrjQVMnGZRCrSW71duq4eoft41
8ub1vnADHu2bmbwMcdWuBbXVG4EwtntbXcTHXzMtgFJlir26tZ0wgdEmvmPb3Hp1
GhDjPVs/QpS6HRSHF0woZmT5piWwWAwIs0Y6ya/05fWXAbpBzI92Zui33WLgF/Ld
TbcuLS8uqw8Oztyy/7xnbRCdRuWSHaiJWUltV2k06f0ovAlJUrfl6l3LWvoavXnw
5x7vJ/fW4HB9Cf3fWQ59clBFGStGGqZXXa+oxfQeKAKSw5NTpDpPYnnVlgK9o/Ih
o5hu+BXOUDpY7lZJSQqOyN+kgy7ptEhGoH8rnalwLvNoj/w3sV/Z4w/lG9o5Jn8U
qcCSnhui+ep6VxA9XZ3nQezbJyfb02aBN/fHDScAnmxU9VTPNKBDoL4Y1ZEzYE2+
an/d6wHls/vCWmM/Nmn/1ifMUU8dDRZBXZUaBLfM8nuft9P5tldVakbDA7N9NyK7
b0BUBjumL4yXiMp4/EWJdFxWD3Q06uyPtZNkzsjB6S3V5Ax6h3PiOqFi+2C9+XuH
23L9Yf6RWXblQBkZ/CAy152/QbHbuTcHCpn1pKDP6HcCGVgXIoA9x/pawhge7Et3
aOx5kxFwhutDkEklz4SxdYABgYFizmMZSCLDgY5QaVEMN1Y9QnuraJAtmZiVWRnm
jusRVwjyz9m8Sifh+JLujH3vQAEWafpd1VF56T2U9qyoaK8B5FX/V3UzvxVIxN8K
67TrZFK5W6eidouzH90MaLgkHI9+usfflDb8tAng1jSgrKM5lN3rzmvYaRfxQygL
5YO1T6H1aJq+Kr+TLGG3mqL4SJAJngKXlbyTI8Mjht0EBZFaclYuVjIoDFvJRDGW
vHVhNyJx3YQFAXgfZaVtTcWVnXrbUXs9pKiWGpYFaVFGcZtlmtNrA+cgIRye+pFU
tHp8qM8j73i/S70YUb8VWIwWRf6OFKMsbcWNLLMcqE1dKzGbtU+np6nylRFbBuEH
M4NoDoTjHFETtJt9PO4impwF0eIca19BBSfsd6Eur4gYOC7sp5bVAP2qN6n5Ir78
5k/mXTwR3yAk/+sfV7Cd0T3SXfBOyUEZnhq/gg7st7qOkLrTvrlhZdreOo0adOfZ
fxqEaM2BDuDz0ieDqIUX/QRjEEYDtFtEYjCrwUYBuhn2NIdcEhRbVDlGPV93PLG9
nGDZsQLwVGR/4tpdpJD21DIgmKHwmc0SNJap3CurmrmdHkfepobzkKI7F8C3FAtA
euhRKFxiiqi+56M5W/trdhFyjKQq67Dk4yBh4LKpXov/XjYcajb6YA1PbYbq0i5M
KkDBOOmig8HGn72PliaKFfE9e9q5NXeunIfSxTYFMJXgQ9ONKXD8tsDDJ+HWHuJH
j+KEdFhhn3Y1UGy3lnoHzB9dpK7puvN8JpQq2e/MV0pZeEejChTfwhiUAD7OYNSY
VTgpuOKBzCGbRdwSD5qPPjI4ceanowofRz84/Vibfkt11L4J6pZV1rNUhH7DzcEZ
6/gv5ZaUOu+vNyMMQ3d+7AyichBrEdQdhmK/40i0Vxu0knCiWn4w7NkriiR2Vxiw
APVTqCz3uhGE/L4DfSP/opPE9Pb1+FtF1wHeUq3BYOaVYysuiYhfpyOxbymH7q6v
ZBUbq9/OsFyF5wMtBsHNb2nJXsXG18iJ1sOmQR+LccaEoqLxvNByPh8VfsOnMxL4
evSc1LRgbmyBTaE37SsyWDS7dfb6lacD6Vc4kMolY8gD3+Zq+TX5BXZ+/jbK3v+C
h1BR9vZ6L+rPRNJH8SLksTLan1/2zt3KY6vsRiJz3Z9J5cgZnZhRGk7p/f9QT8dW
i3UWLflyGdf4AIIQpgKfMWi0JAwsZ7ADDdZUrjr97phkGHZRc4P5vE2jteiWqkZq
PxV/hBx7B6QHGhj+EHIlvzY9/8iu7apy/giU78hnBvhp3LlKwDYEcsNVTAWZPx3k
gnh0jhWbiWuvEL6XMiw2l+LzaCH/IcOTTkt17Pl2Vk+85I7Hxa9Isp0pKikwtWgJ
D9dhPAAEl3EXjjbhWHleagcxIstuWXQ2j9eVqWOenxEl7jwrRrw40Bkbp6H4HW/I
Cr3JMoKYyedGLt+0fPYMNgqIkmCFiIeH1JxBi2Ag8rfd1HA6hrGnq6I0UbWIylin
isiVDKHOxNfhbiG7/X6WLGVWIsPlGUJRoaBJZai8LlxOpYEG0GOXrIpOdPhQtNsZ
n6jqzLFeJlnH7eM6Nt3q2CNMQb2xWvqoEXRWEdbALRYFwvjl1Hk0NBeQgPFcwg1k
RHgxwZwmrSH10RzOC8lf9eW8Vc9DOvnEWqJ6A+wTOXN6WFwETL7WKna7xf2zWaTn
XHs3JScR2PaUOpnxZ8QniDv7hoRxPkP4+fcbXd/f9YwIpb1FJK7VZjg0c9Qwq4Db
MCeuDDHYb5xUK8eB580xf6PZYvTuUhbqE5IsR4S+HgMoj/K/XALlgzIzVx50hgWQ
ClPg/ynp4uwZJRCaBSgQKrnIwT5TJlmyCknWaRBOUqDIVWvqP+XsvRsxbi80FSLC
ikEYfWmPsKqVPkYhRlahkH954bp/yRQTO6DOIkDWKPz+ImK7hRwR1EHIYi+euZ8m
MVqoEUOkiu8ubyGaPM5ANtVcxBcqivZK5ypmBL1l784sX/O1/d0+RvZJacYAbUiL
rR/f4w7viXMYnbomZaze91AF76e9OxGkGbJz7SiPpAiAgLCksBg2qpgSVTL5OFnm
sodYyn4OMFeg4MqsZN9tfmkr+n1XhnpQEeD39w2YE+li9dkGvFsSv0YXjvjAyw5x
GiKtx0Ve/jp6ZmC0eYBMXZRCS4jPCql2Ijw+8yvWHV8eIYxhGx32721Ws+kIVisP
Q8AS1QqXno273iQ18CQdWRlhWbvini62fgsHIZFxYpb+SNtIecXoUuhqoxYw+O6o
TDr8O3G/q/f+IKiAOJs4afSOyqwU5hvV0K9zUTD5QRg/qKuGfoz1eHxknT7wM5kW
hqDE+mmml5SqDMixLcj7t/ZDRrMFLXLOxeF7GyWR9vwHY3Lu29rzzm8xfg01Jd4B
/5q7ZyL+W4pcDBTf7p5F6qoxBMCZ81aZj44Y642H8g+cHEOYmISYpoZhO6aMT2CS
qItmYEoX10wQWd+QvGqj2MZvAHfgXYxgOyYO+8m61GycNSYMlz2S8MjJwQGyFEpA
7pFXT1yRm0qTTZflIrKHTtoqSl4y4Fg0ZGaQJjfUhJtNZwGMnb4QlinC4epxY7QE
9slkAyYcUhncn9XWXk0YxJ+j/0YH4t4CKsC3p+Zr6X65nFGqxMS7RAvKU2zqzLCA
qYZNyQiEWIFABUF6k3YdPbW+uAERZuW8A23KkF4p3uMbQbJwqlcRvaP8ewJCB8qM
J4FCh0SSrVrvV13R0y82kHPvqzttvOrh0k+o+wjMn5IHhRMJ7MQzTC2eKQxAPelx
oZVw2jS89+xa7ROPdUgRRi0suegaZjhLnXG+59Xd5vtOwXVyWqPn5sYjY3IcKGbg
b+R4VlVg5MnxJ1OfziPFGNMNo4F5i1XpxmkfHxeJ8rhC3pZaMQqVfUPo/yuRPkOZ
ZsFdH78dnLUxiUoDoH4gq/ZO5BHGZzuHPR6Uih8PtwK+8fOoThgEHskw4TM523XV
CA2HF1Dpw7S31Cg7MZR7rTgkfQ9S4Ttu+zIwBS2giHFtaOdwgTZBXSsYRUytMlyI
1wbaImQSU/JYjRpyCSQiHEGArlpg9dDNhTmnW/aB/mhYJNsfPFTwhSNvIiRauDgZ
e+eAH1FXof9e+W0W68DBRoqLkC3MUZOjmu2HPIzvyLPy4NqYVj9yEFMG9yUlo8K+
ICUd/7hN5mKQjhGAbAk7zgaHBkupJqUw7sWHzMP1OmnQJpQp6ZzPNWI4hT+JcKPI
BLC27h3otk8M5Rr8XO2yJC/onK6QnFh/5DJHELuQfRdxBxKiUYN0hQt2IXKRrB6S
1fI5mZo7woIql0ZpoeF3e+EPerreZ7QQq8vQGSW5VIbT7xXWl+Nn4pJCw3bBErWw
xppbkpuxZkb4I6SBDRAprDgcj4cayW8gSO3EveWWYJiuHwjyqQuSaSbttEyVdmMl
fIxoAGNeiNifn7SpTAvvSl7OwhVdckrnA1uWyH2uBEZvZNrVuDZVK4Vt2dUoH7yy
plOp5UrpKlEGILoXd1CTWa8mI9ejONylYlBbaQOr2AIKs3ZGXoAVwHq4wbxkdYgG
LO+ra4JEB0H+yY+l5M/yTw4tKe73ZCrNOsDHlgHnlyMM6rRiG506xiFeVy2E9akJ
TOTlvl67x497Jv7/mpTbNQnJszHbMuZS3JdXT/5bNEn8fwxHbu+vVlCcchMmLS4i
/I3qaBy16ToI0Adw0kX/FT+Iaso8XEcb9v2grcwEUZuJHSK+usQEyHbpWHzrkJp1
smHXXOPLhr6OY/0yQWaUfiS7vQc01+KrmEkv0ebhzFAU9PSoC6LYcf2/gJ/yT3ou
hvHk62hRdlrhtgxo7cfg50Bk6oDN0q4OlBrQzxaTATfk5DpoyfbYmExFm0+j/AhY
yE94vre46eDSlAXJ3Xfmt9i/c4KwUZF6zZBEeEP1sIq2Xl/dUekgbsyeCjc6C7pA
+KT2bY7DtJsepB2ptL03tDp3RAjbxEsZZNwRi/h6J+ZWtiqiX3M4Y5h4g0UJj0SA
l94NO56fnsYMSzs+Ig8HlZ63vmcDutIMcNKnMvODlj+ZYJg5H2H1VkhR6rRlS08P
Vo2CDA37A9slk86ec1VM2HesHW1s2LrPdK2OQ51Mb4SN3bKjrKZqKlFTVSPt8tbX
OeJ/YIcQ3jhBP9hOH8NbaptSj1KPeHZ/OAj0QCsQHStFg5Mko9bPZpq5zKsN7QhF
NPbzPYKpt+fvfdKsD2mpohKVQ2fimei0yEkoq88/vuSPTyvZITvhYHuggt7a1JYW
svyf5ze6bPx0BX8+F5z0MWPwhl1YRXuzdu8M1I4qjleO/OJXhJa3Ogt1F9wrugzj
TAxyXjvdiymVo0qchGfQXRqBs5jeRgWKwhkxgRc8n1dm29a5snenen04CDnu5+B8
4ZJew7q3hmr47+3Z4TbgV3ubia2xQU98P0A3lMLXL3gDDjqKdoSPA4gT2U/jXhF8
+Z9izwC+HyN7T/kOXSo50Ho7mUW7KR/nbV67eQ8HrSdRLFbs3NfV5NNWBGaTnslG
9mNfb3nmV9LrUjHCjh/i1uiNx2xnmqOpFNIKJ9YCYc56elsniXb5vepOhundn07G
YgvqHArhhhA/spcH6lgZLMpyMhGZPCR1Q9KoL8VGCS6byK3y4BPLV67w97v8QFSt
B162cRBUt8f6jekXHNDH1yNWSOZaNtdwH0T04svf5e3Fq6N+7SVQ/F3ecVJU0mzU
XN0t60lwOw1wtWX+Gg1bR8L/SgWK4XI1xgy9h/+7tnUwuR/qk8I6ANAWgdew+k17
asze7RJo39E3Pf6gkVNiBm6wtnMTomDp7N3r2Eo9z51LCRW2xeG60RMqJ2rtzS9v
1U81V7+yu7QhOQIc5aHtf8Xw6NSzdFEcpSsuXjTI8jiGfhTA/ROW4kTpRup/yZKJ
wMWV8VOLoWjDRaUQGqfGHtGMxlxnUGguIhbZA6WXRjO1SZJNPZzsAbVNq2IWF4Zx
pRKGX5KqqgB2IExcKHZ60PjGjR6Crkt2+zW5cQss/zc1bpp1TuavoSWFtCPiHRxW
sPc2JqGTSV1Osm6QX0ferHIV1fIS93XksZu62xfDsMMqVyFC2DikZ/OTv2E/KjHY
4Db+5/lxZTqy0pRGNuX79Czn3bAlKWvKjHT2gVd7CJMW1V60Krpd/FO5y3LfLQA6
kOv/a+qXorbn/0B+YniuY1J3BwDRWu/JnjC7sM3OmkanxmUtw22TPQVwFf0l+ov4
XlaHTImMGb4kwY3o+IJTxx+S3xW6yEPOC8j1EuXNQlhBI5cOOqgZzLV5g2a4e/J2
5weyI9icnNCIl4owfflWJByWDUNQHjczlJdA9HcMD/GuKqCv6l2BqcKgNYqcd2nN
nSO1BhLAQ4TCW/oTWTy4PG8T5LBGeuDGLDWvJL5/j4z9u+eoGqcYs3XWNpZOWMMS
XBmMbURtPMknqzm6PaQ+q8lxGupHhZJjYzrJ8zK9tO2ZW6vzSozWMtORdI33SChD
5S8CroNeWFWwoT1hF2S2uuWUly+ThEPzT5J+lputI4CxMHcNeX5rxlgLJFnzJjEz
08XQud52/e11wwnSuuDS65i+Bc6yO9/oPRJilQ9VRtgcB5m5GgazCt+zfgRlmw/7
fwMCbTw3gONE81Ck0ImFMoPEAkgSaZDuD/tQ5SBQfoGCL/aPz5bbjxK6fHIkdvad
qtg/TqoD0U0ofJmtAcnWHPzMmuWOokRco77IEcDxT1bXgXq1Hynz3M7n9zHU1MVl
4p3pwaXSvMb1RbiWWAQCTGaN9mwyOPgmGP9caYdbttaVIFItFgbnLqAoprSk9Esu
ihMUMS6HhM/maKjf4iMwZvbMtx3p3rPHzGChDf9KD6Bzsv+t5hwrvm4i8g38D/s9
LsRaAYMwaw2tC89uSaQ0wSi/j8e/hgSweVCGWHRzP2H+iKOg2GXM8yLyxvwnYGh3
/Y4WUajcv/7yVSEC5gmq48S81i+8Bc5jRRdybsaEIvNsYEb/cbGWLJldloSjNUWJ
t8DUEVehKVWkNBSU+Pt3aIQc3+1bIMG1iI+J4lP3ay5VXKbCftuU7Lw7hG2XXap2
V4UDCy8KSlmZzn3LH0FqB8B1GfZAQqSrmn0cJ3d2H11XrRzp1ZxIrqbQs2Kwuq00
UAhJehuaNpRQr8JSo+d5PDvv9T/ZUpLej3OhekkMLboA1H2jNIIJ055qtI2TCJsp
+OSnXd5DvF1P2kGrCUcB1txpVuAeyELYA6S0UcB+r6fAK4YpxSXujJCkfWPHRblR
dPDz/GpvNi7tqRPfNRyYvf1H4/AyzM9coTPrby3MXHc6pZ/k0iGYv+qlwUpi7bsW
bWY83ouUURjgnJu2ccvVkN9vLtRvTJmvuqbvzGsthQ3D8pGoBq7zXaLTof3U3gJe
iaREcK8c6F+8enOYgt7a63AtjCMHRP4Srm7wdUtOuDbBlPS0/eWXBpw1uDh23b40
ATBRBvK53a0f2BKmshftMvqH5z8/+G0dcgj6Hx7uwGfA9q38UHREp5QaIGp4rS8l
xyog9t27GLZu1mul2rUPFZrr3F9YcuDHisPdhVt7tmuPCih/01DwpbLL4bJdwyOx
4t4eO9AfIHLgZqQEp0rSIzJPGC5HsXdm95Y0QdrqcWw8ulGOUwgUYpeDuxjTWayy
9W7B2QSZARkuMRKoFoGFJVK/muZPwL05EbKy7uiB+nP4RpygOplJa50NRTlyvOTu
maM6ZOgZGZEWCO21wHCIW008jak/6FkOYZ3JfqK+s1hZ7gTu+BKFFF2fUNnm2fne
PgXKZ+jgkCmYTIiZSaKKxxSjWoFpKJlK5b3rsIbmSeos2qOydwbvNAFyly8VrwWr
PA0m53bAcrG0U+6x83zCcolLv/KqCL5pB128RW13u/Nq6YZmrbl8y6i/nHvWO89U
r4+b+2NtmsoDMRm/GYSn0b3r1BKJE4VZ8o+HHFLkXegGQ3rKrAqjnNf7XpALqnds
88z+RG10MhCM8CTth92Sdrz9H9dykFvIBZC8yyq1+YyDk/9fDtc9Ajcbx6XdbbSq
lfvTWoP6ifHN6uaNX4CeYMXuqJcyieFHOzVz1YGQQW0laYZMSbyJWyleDGP2W+s9
ZnqdeO3C+aUulQpnoEKvguXAM21nm3+wQDdYfV3JMaan30+WkQySwoGjwINjssPE
c/C1q1BEF4ASLHvHbE/7aK1GmtJJlalihJ5M0qdl5h/WZXVNZ1Qa6Q5wdrq1WPqW
IDrQ3N74DrATfbB6yU5qUzubIRd/pvSEQZagbfhj556kRVDDgJYbBKv6Tus/CgzS
a/B30a3e075p4oe0uZ4bTHiM1+AkK8shrUxbYTt1ue2FKEietsngOVhxsq2EDvfz
rE5/uTIhzenvhS5Z7WYJ/g82SbQ2Ip/chjgMKq6HkywGbmpIBZ7dkQzAlBD9a86n
MHUz3D44Ooy8Ppy4bKnnOihWrohHY96TgbdA3JSyWX7dS+LqTI0bxH+wjYZ6fclH
V19gM7uvTqq8PPzxdFSXILBUgkfHHNRlBxbG096jTe29Vk+ylwCHR+RnQm21EI+o
v3iLqz7c9bF3Me1hBSW4LWaxZVHqY91fx090seDsJvkrUf1TOjtqoD6BQioICBuK
dvybmwXlQ2dEy2Tn0NSrObLqjzDuyS59fUsILvEKUu+pMw2ZvVBEgBfDNtqSDd18
Z8FhwuyHmjpZH5tOyO3aOrzSeXxC+nvnQQ4IlOrb9QWHBDpqQdHtTXd+nB/7uUIO
qiPKRjcVYsEJkWh2/4rCcRMqXCd7HdhQDmxpBiS1ECLuIBrhgwtKaKrJac/scCKM
EIZ/NKDLTtYp0QdGGwO/BGZCbM7DVbrUpVwGCozXUc8ltfLTNW4gDejjv0vKpEJd
wPDe2h1YBNbXNhA5mHaS6U+75lNAXoEiebplqhScbB2WsRPwdKujgyOZjSbCr/v+
GHznOWUmwEwNdHmlnUonFhyoetJsT2e3KmCVmskGyjuT1RRB/W0DeJ7/tllHq398
aany8hstmvivhszEjH9EDveyarlf0wJ3bbYE7WLLfH3fQRayqMaRaHy42fFkl0qt
TA80nHJzsL56q4lgQxsnNupHZKpI87GTY189880XxkTZl97cqsM4D3YM4aSXQEsp
K92NA09/42w6r02asrQGUqoqkVZmwMz4FumNypoYYH+ZAy34lJCA4wSOBM+NYX6L
xhlOGrUYWDahr4PC64m4i6tcWDoIGZwSU2ltC2qgBTLi86vMApPMdE53tFTRVxNh
yuP8EII0R0GNhec3dMfNB/sEuhiNo0rzZXw8m0Bp5V1fyKrTwGYchAPGxNWtaQ4h
ajOylm6UxE6zf573P1dEto4+jeloqzsI4YjH9Mio5XdYBYHhOLrwfBBdhWsQD+ZS
CbsaMTncrz+Aw03Cu3fgjWAyshwguSJ11OuiJhB3Q0/iDax8bDc7SeMwDzZcaiyk
B46ePZt9agaEWuche2NaGR2XKpgoPPOTU/lxqK8ItocCTf9Q3aTv3soPbET644GD
40DBHgXGTTeakcOKFxbs1IoHPRQgbfUcfDUEZspXAuEYRp6jhSlnee0USYl8/rUt
Z1tt7ZCgDu8LS18ZA5f+xgh/LUKhE+L0Ud0bhPgidmS6tmXSi8X9NVBaZQxkVvce
pWxEX7BEIEKTiTYQ7Iy2pqTVYEvoydBWdzYa1Nc7Krdrz9u76zJjSSwNvMCWUpOR
D3oZR0yF2+fwE9Bx2473frEiASM37FucUbE9GeChNi+kY2KDgdkUPTU/+rQbVYZl
oLRxmYdY1pJ87rmdBq7RUV5DSoNwMm9JPB4uhAvNmx2h7b/CiEMaIFzBjdeREyOj
yQoYYIqlo23xge75yyAMMWranwYwTaz9EVPZ4snpir9DJcKVNRQ5GwPoxvF9rt0f
k4rEwkE59Gs1BJnC1rj0VaRtkqujnN0G14hYD/pd4zOcM1vqaEpsuf9A4sxUQKhF
0m2ZRCnVVPB70fNRiCQqhvA6sBBERaiT0Qr0YVp7GRURszb/07XktbedZrxyu8ye
KxCrtSI9SZgl7kcLn+u7FFqlR7ZTNKHP4iGSBBy582nJl89SiekCeV/jhzubgVIm
cADskRFiCIdFRXcW7qO6h3fe055UOdw/TyQCyDUSXt2eLTzH5aIkfDRSKTJ/NjtI
C6CmzF+v5EIXYvRIIQT8FBNhiliEqY1U3DVk8K5eTiRvQVXOSua2SiRX6S5q+BA6
EWQ8nXFchururXDwkJSQqQISKAN0AHxNxk/BQ4kFBehEh/xxj6Cn6bC/Ir4pNDGc
8RbO9UW7ZoMBlDEf5KYdiqjIQSvlOxXe2YdgXYCavLE4LLt7e6nSH7yNKbyMCAJP
lq9WY/10AC9ofKW+UMcRFamSbaawbbQd3F9GI96HJURs5uBUhiwVYWwIeAaXt3Ye
Zz16sVWVh3q1WLngw58YQ8Uc1nApFTq5ZR7oJeEfBE5MeMqmMhS8xuAV/cDQp4G4
ITKzFMrOMwD8WnR8fyalXBXt4yBaDjAccBDh53FbdXpOsC5ZJq3z9QYMX0bQccTq
UP68kilIi0+7Tjh13h8/fq7WFIBUFugSUvrKIhOCt6lCp6cII2GFJc3CA5ITVY2l
7WipACcAAgI8w8IKdTRMAq0z9BdKLS5nCPuj8W1OFcWYWGZN92478Y4ipNzyrNLv
qykEZ4Dah9cjgIopf7aMgZE+bLt61vum567DzpfJlrhw76m6ZxAyDiEWDuVjNFER
8gPre/MOFoKBGIB3ryVogvYL9KTX4KiN1DDiC7gQP0Vuh2YLYOGCcxHfpEisEF3L
++qOPtv8MM4XF1hD8Flo+eyjFTyDfGm+YZ3QpTAED86mxureqzv0vR/d5Psh7poj
5K7GJsN0PujIBbSilQxij4ObPai54DdCwuIkiq5pH0/eE1DO3289XN4vs94fE7cY
x1+mK4jL7caTJqIZgdmtxf6fmSPxwcebYphc09ZyLkCZMA4Ot6z8k6IEZmDEb9yq
NHJ8o6nDHVtd6ed8c1FbEtrxopvjbrW6IW9kEQOldSJRiNUm6209qoxH+YIPWIJZ
kgpCAx350l1CNHXa1tiFAEUGt1/IY/nvhpD78UDSLISWE8HqaIYGFf2Tb8Q9xDDi
OSK3AUFqJn8XUdcQcpX+VVKeqn2KOVbs0KoKkYZ4Vwd0yvwdnJpEYMI0pk2FPuHi
PmrypMkTst4d6MVHI4xuyNuKJ/DdKJmB+7dDDiiH/mPIZEujKuv3TDvhlp5Qku1I
blkKWbbl9oqp94YRdqw5YB7zjfUqU5pVEkQ8T/d+C9h4R3ZmLgy1mGAucDAxgx0T
3Wgxc5Pzm9kPVy7Ny0Bm1mcN2zoEULd595573xlasMUHi+3YGIxqKBFvoo3vXrOb
ortOLnCziWMPOGLAlP7CdarYIHot7O69IfocwsYfLqj3JjtRBo/vWZEoIKmSgDM5
7qvnpfSKt/FkZdZe5OqzdAwskJEGabiqXqRC+JNOrCvpOdiijGbU2tv4UcrBzCNY
gmgHdDDjToE11njEQ2wQXTtqy7D6fVef3qH1e/uBvsHXBTN4PVmv8crvlfGl8LwG
v8Iq2NcnSHW6ztuawXKZ9hYgcNyTOr7QkXfkpfM1kh85ehOCbcLyDEw3M58PMppJ
kh4wjSUSutc40/NkOmid4BtLRcuQP5WtE3SvwvaApl89Vo9dmkc1AsnE2kzhpIZT
N/XUjm4wkZkNFfXXcrqHxD47vInpdMHGTJV956YdvGVRXYM+TOJJN65iLaSJF/iK
UAwZHOv0UiQkQhpNZU39AxpIg1rzsbCCl10uruH6JWa9vTKMdmXv6PsZr00rGlOr
XmxYtGXc/12kMi1qzmljYrwYj6iyxgKl0PAAHS2qgqKUXrunYUrFXAVehKsVZGhb
zllllMoP7YbL/HSkF6vCXNuH7CJ3a6/1gXwZADkHyYWHLrtH7mp0gNlFRROSl3u+
nw+nKR9EcLfrBBf/OWtbUXiqV5PC9LlCwndE6ngsZcOakcc1gGeJ+o7CFQmLc/xT
x/SM8Fbuq5+x32RUbLRQTSv87+5doK3VDYliHSpqNi8K6BII+vOnLJrNYMX5kPKz
Rfq4T2BRhoHSDUlSdqRtxH038nWgM/nHGCHuR7HZBly/c5B/JSVUMH8doqJcnKmZ
0bvYr3LMMzyKF9s8T4uHhWbWJDEWfpk3dClKdsl1nykkDUk4Gi59fd8xbD6w3g0Y
p045yrZ0ElYgFbiUkkbZguP5aGxfrHJJrjxGLry0BXAvGlMO7YB4cIBODUINotiJ
fD8wZp7L5i0tb7U/+gRiyXmW7AZ1yo63x3715klaopPBhU5KoLYU2kJmzj22JM2i
KVnKAUlldnWi9eQkh5UGAAh02jNwi+RlIISOvecNw1nQ0HiVw6Z77Rmi9Suj39nf
n8HeP3EjTcqwmTOHdZXy98KDLv52SqWg3ZNmipPWDKX4QXBAZwU8t1vlQjcnL7aj
UyL7oXVveNIhZcXwUu9QBR1QyChd9MoAoX/0ty29gXekvbL4uxmtrY5tUgs6XsBI
l+OZaVM5mvIE5dOExmHtHGKn3ZZVZXidLI7QyB8BSMH+iv6aYtuDiB2uYjjaCfUh
K1sj+e/p1lu31JogWpJeEZs3hXEnIkb4XqB80X3B8Qs0ddCwQrEcU1NkNv6nb5D7
L84YWlIAEWbRYX5izhKcJ1uSdLYjcRCAUL6/XSWJuQGj4rpckS7etKAWhJuZmqRi
uOTP5naMTFakC6cRYxCyzfVA39OR907CpMG21fBloinaUXDde1YTtqcJGzap6sei
78KVEff7YXOxKfzpnup/ttQnTVbb7Nn4AU/PdCj26NkeR6yEZkB9ocVG6FprJCa5
FDpyZca6k8t9FCjU5zFbxy2l3bAL1o6dLfAYLogWTQ4AHnR5YqMrpy+KSDK2/4sz
2fxv3dy+0N+2Xbb4l3LC1nvNyomTJ7HigheYXQB7VQDpuh9SsGTPlNxP0iZ8DU+4
N9oRMJs0zw+/jQWArkSc9SpZMQxqEH4f0zAYgXTXsgmCo0MKEkFb5f9p5hXLyYuZ
syZ1q6srXoBEtqS6En63MByd6hTXjlUATVy1nKNxtIY0DOkP0z6uJ78Dr4re9ngV
Nm5dWUkbB9SX8dLm5+q/4t3laG3rA244uQZLgTwphXX9zDO1zuu4NzmFaoGOs9w7
ghPNw0kYHykqpcfToDY/rwg8yUKjELxVdIRs+SSkmJ/Jjd/lTyWuOyP+pTbJPgkN
SWkFtMbqYqCFkbErAt9DJptlxUJAqKjDmhlpwOmbh9CV5M3hlG5E6BY6hnpOfLZZ
B5/x4q+VO+oFhWeVIH5+lIIrPL3ISeTlO49Y7FaoopjMfcYS8N4wQDNBhC64IzU+
6wlDinnbG/39eIAFfijG2PsCt/1YK8josyZjrhsSkVpj+GDAqD7ycxXAxNPnoeRR
umB/VLIRyovElppx3RtpmMFTIRuwUESA1qlxHKSw3FsbrJx+brOQe1S+r2cBlgCb
OpqBuCTkJsb36hlNsENaG7jriW3mGaAQhwAly/Rqncz1hWj3fpXXr+ynrL4CIGSq
LEB0DhSLPnb08i6kylrFEpifYDqAPlptJ8XSC22K6K8BjNuUqKONGdrhpkTqdB06
ReXVQgMV0SuGrEE6yZBajnFoLS/W+V0sbVl+ict/0LcJG2hSTxrdCWxMQYVWvQZG
U8UqwttyEGW/aVUj3ICF69Jz13ooL10BCWeuh6S31qHGOEmtuAxNhga6KOf239g2
VhRexvetgXOf0gox/+n12ilpYiliCdWS2oe33++ohUSsiD5hS94mUQCo1Z7SjEZa
4ZfAE5E8voAE6Tpi0gS/9Ued4YUOrsZFV5hiKapwht0WbfpBum1UIQ8epfxw3MOC
DBm9g86BvZnXv+EvMf5/qrmpagzmy1KItMPT6bA077kPKIAi559RoZbIqtwHqRU/
CO5dDfy/SMsX5Si6Cf5BHfo1K4lCrOZxkNIK/zhiopbuOPM0WaePViCjsJlwxKEG
o4780Yw9vtnjDlA+5W9K/1bz0RfhDOSdQ4Xo8CZ6J1LgyW+iWmGNu7MTUR/fEuV0
g4n4IVP99N4lz9LsrDfBt1PelRhLeR89Nx2PVaDX121jAxxpCPVj3z7slevW0L3d
2fDqj0Y0CID1vvnljxapMDHG+8XOauQCeju8bM0EasrPXW4h0IFu8ohz4vIaY/BD
nuq32LNv+JKemAvwai4EGOuD4P4tRL8lXgny+jt243nVs4zQzq+lOB98OXUUAe74
23vhJLKBfndr+Enu09+QLWMUi4X1aMYA2OAzHxbsbEuNlXCQAJ9OE1NGE7ibYEII
jDEjzF4edXl5mPn3XG3F/esXzIPDKKky0RHyc84ayCl1oJbrDkmCk2DlTMXkOLaM
o8Ym8LQbw2WSLcY9ZdVt+Huw85PoWUrKnFL1dOGmPEGKIy4RjoYW30Cs+/3jfqRl
pVi1QHIIPLv0af0R9iKQ/L9M1J18BsD7rMqRIqx4xmOTE6GlKH1vrHi3mG4eX0dV
ANNnHFpLtrGE2FeCsWvwl7Y4rPQpWg3YCePl0DXubva5KXQ/y0gAb7amjIwUGBjz
Oc0VkUfpdsUtwEMUSE0SCd3vkqbhbZut2gXFYGVwfXUCHnfZ7cHu3/Avu9V17F9h
9c6i4w1zy62bLKxjlDcuq7zLI4Fjfj2eztralul2GMLscX2n6Pa3gUlJ24/PqlBC
cfjiXSvutIl6fTzoxl+9ITeevdCAwTkSqJ0S186lK+gQxr288SSMIHyE0YZn6+B5
zIpPcoYBOP+Eewb2UuX0zI0hQ8bI0tnFNuSbuLkzn/AxlQlca1INyRREKmhdwTgC
hSKS2RbMAJUgTeVqkIrAKr0ToVtJnje74An6aVHpdN25sTQ5QZNiYdRoI575iYK9
VvUSblME2oAbiwpdJTqTVVnUx0GvNuGm4/eqR/zKdVFHEdCXzlmEdbfhgVIowdpa
ZrsMbF7TWWflcDPoB5HoeKfxW4nAz9SoNGqhAeLXYy0EEMfsNfvbLqhW+LqAN2yj
/T7+35av2cBWPgom1UYYsjXbwtfOIgKaVbRIt7pveHVImhkI0XotHngehY18pLrt
xwTeND70i2rPKayBims3Xf5WYV/gigiuo1N00XEMbkVdVrhlAEQtm+7tJF5mmH8l
ZP9jNAm5oiN5sPgqoKqj/RUxXFIvJ3J0cpdMndBYtDDKT2x+5fXlVEmIG3YBEAGd
FxnguCMEzb8LZV31ZkBnFr4f53AaYKSgs8hV/3FacKmeFwd5vGH0X6A+dOFwqYHf
SrombOEhjj1xj6LI4Et+hNz7BDILPd3bTyTT8UfaWpMPD1s2cStjaYiFyJmdg1bT
Bb4GwzONlSGfwQBXmr4U9hTpdatqYG+CiRiqerEiXgOsfMeS9KIvTU95EtzyacCm
k7slw9Rv4Z+tihOKX8/ftSo8FuZQ1IFSSoBM6xb2YiyA1VrXw8PqLqov+WARtQMB
4aA0CFDpgDI+G2RQJ8urTh0Um2BhqabhIFpPvf40pPs9Vkr22zxnQtGR1oScoYfQ
9WAfSdhzN9cGaU1RHbw1YdfYzAeL30GvIxJLodtPnS/oP2jO4SAx4IrABFy9c4bu
jpfQcbl78aCnKp9SnjpJp88UIl5EzNj18T7Rp1JN4+KxIs7/d7aWJRbhl9i1fFdZ
V4Y6T4OySwzbk1bbI8g73FiqriAMIq5uLVVZWGIcB+hxXfT6IYcvsloZwY+fu+Jg
JDZUWxIKnsMi+ERHZlzxaju4QBi9iAzm3BQtWculzKCKsn8VMgK02wt4B5gedUYu
NfCZmkYO57ED9cAnFNjgvb8dvIorcwtZO6hhIDeSNEk1wWSyeK99QnEtCGcixNF3
nfqhhUcC0yOnkkssFGd8FBgd7ZgMMcuQ1/drrK0EOSAPaPjpUeoKCTb/OTcIqhk3
vN0cJ41ckaovSxfTfR5I8AYM6i40Zmmneh4SSHLV03iyTPva2B9Vl5ak6+s1GuVD
P/JKqmHuDwZhgRXxrJAkiPZ02+m7gG+9CsDJGcluJPvkCBGERgFCzJjLnTFtdklu
LXXilR0hcJP/cy8ikoI20xCCnY+f7U5dvKcF2a6oCeIlTlP9cFDzRcvO1DQRcN1H
FeuV41ITzdEulXn0v6moMfpftjGzpUrcjcQPVaX8O7oSCueBpHRzFvtbnnru6k8a
nBaDza6i67T3aovAWzJtLoJ6r091VtyaPB0xHfKCUIEwdnARgmT46dFeBcDmkyeP
ca3oCk/WckvE/Tyw48W/1bWTOql1HPfW4vidHuwUXx4fopcg1eMTLW8y0hD/vbay
aKcXCNyaj7w72ZcHi+7rWVW0mOJqh+CpbPVsC3BFg6jB0IpwkRBeDqMK9FalwYIS
bzPv785LXI7GNc7f2YPMKF0roI3sxZH5v9IwF00tFRyZWmOzNi9KF8KyxOQZeEiD
E2ETEIBtdgw7yztCI3LvMNslCZHvg4THnE+LKBdItZgjVlzFYymAMvN+8dmpYIQG
OmDyFJ6zZ4dxrMwK+2xUasQMmNkX9VW+ef2uFpCmQ0sFSq7gc7CHSqvuUaOHxHm2
HM6Lmxp0Rrxxh704fMlhwGH2zngBlqX/ejYwIsQi8HQ785N32Cshov69sLpCT5TD
KsY/3LIHzWbvvwBHFBfKkKeTJ5tmcW9upNCYHXv2dFN5GMSgmWRgMcGmbQJ6v004
eaCArkIn6BUKbwAScupRSGEM56trUViidzbPBAD05QlTTEKCIBlk5bN7W6MlTAO8
fn9zMkjkKFj6ZVy/6sLAPu1b8fSY+HSkrT6faWBb+Z4QAi0Vxkza2tqRHsJtoOND
TrZZEnRveHTjgByiZcEiovxWIPYU/ApZ5BU2h6drmqiMDIxIhI6/GLZTgdHgaKta
V78hqvUJkuKC9uYbzX/UHPvBFYlDtGlZ2sCGJMdpcjHZzGO1ZnQDpttx/beaMmJS
szBkJIQ9Sh/sfJQFsxJPMdj9ZUAdSKX2h1b033U47VP9lKEF5bX+lH89yAuc9+G8
1SLPXtes1EfCqgAmfP4VFR3X2YYaFKBz4pbHaAY8kobFeSxC1LS2DP2Pk4c2d1ce
CPndMfWMbV+wOoG4M6SVS33qEtutSQs1scPsfPKCD7Ay+DtB0Eo4u9BCV145NY1I
dj/QloKiYmdif40kU2AIrtyPSOt1LJ6siw9vR+zzFhUD2rM/oOV5y5zZMQsymoYQ
uEFroF3AIrYq1FiO2r65JErifG7Vznu9SP+iF3kIbWuZG0MEYRSud4NrTmOCAhDa
HRL9uFRUxaF5CNy7LBrmcTTKR+Wlypt0+jLzz5DDBJchtpcffcAgWwE7fJ/DcL4C
iJl2a5jtfTeEKdudEdgMuZW6ccBtgD6dAHgogjnVeZNCUJt3IPAauH9V93x9g6Zi
ygOPPP7e0tJqhbdVrm2SjvvncuFgBpwo5Za/mXDV9UT+dLQ2NKckhoVkbzTgUC4K
/QZ1vkBibhkaCuBXhWFcmDgSjRre8JAMGg/wfu+WpXjzY7aS1lij66rqG8q68XSj
lF0aqTq7fc55pb+ncUvHH8LcKwuRL/dChwBfW8xEMmyH6YEvS0iZDJtwPt4BF8vX
F9Ci6iJ/SRCVzGLWXvbwNj2Uww/KhpMe/nhOmP7Ne4rqmH4q1pMQfZ0d6EEvAdGb
l1V8MxPjq/r9zsKp3RgQPAXeHt2VdgPRV9X0rxZcCn+P1XOtM2rh45mQz4r6xt1D
NJjFx8iIw3zVrfGLdXvkKSt5wNNAlGSl879Jt/6Gn+RxFd3erBMDvohlXMllsIX0
Nbal1XYE3+mjeXRctciTGeOYyJL3HIqdgPyqUDbYeRTQmpE1y8bXdrH32o+Y6c45
7+PCo+Ba5erbpmvFDPa+9sv9veMGLGz7zthYmgJuQZW21OeG5O+iPizs8VRnUZG8
20FtNUOtpnTQtEHSTnrZdhMIJr8siV/+r7Bmj6CKMzAtR5fdgNld3vCn1XZIfCvg
JSqzISbJ8a5PRHDleksmbhvRr/gNVPa1RcpT0pxJ5+RIrS2SyHtFc+rsHf6kLG6x
gCSsk1jpMiH5uDUkDMdU1mUmASNf27apz4ZmmFcQCvUcKNa3L53Oyx1ZwcF69y8d
PvrkxDWlNxMLKGolRwF69ZRPSld6A7v0r9KCm90RzcvtC65mOl+YFeWbrAcvwrxd
IoVHZHTXSj6eFZo848L/tcwRJr7FAGOASf1r26+BmmOh5Yaou8eqY8G24rSDsHrf
MS/d9d4UMkc8u2yhlLskx29tMWnw9t3qmu4Ng3DMrjBa1wcJddEC6xJu3PwJpa+U
vTSmkgIW5IvxdDawQylfexnlNzK5p54y/+s2fP+aJzFun8gNMGN23mK/zdhEd7DW
93HbLzIUkuOSIXDii3JcWSNCLLXeQhlCsmshdJDorUTP1aLWBdSXfWRcMHhX3pZY
RKvpJacnpckuzuISXTOPMIsNB9jKIPIFiiWBEw24Cn8WHw5k08m62Eb4Dz+Pz6Tk
QuzCCLyIBPav+zhjliizVwTGOqQYzSEnFWjxxMNfmv4H++BiZB+kMtBRxM6t5ANo
TJUH9t0irm6njcC7DcwQuuueVcKyztAU7J8E1SslPHTQMxcJE4KbwbOn2gcEqv2V
wSasS8Sns5ZjPrQ9X4TOyIG5EyojtV3FfRFp8KMtuehS/J71UgPvgNoLgFFwkwpE
vCC/2tSrYr2WLsS6QhnSIID8DQAKhEIZPm2hDv5RKm7kg4839S+uMM0Q77I2NLKP
rfhwn+id5uq9BaaEn3ZmX4Q7k15USHGu2OEr+oNAszuqjoBc9U0z4OXHxMpFP3qU
irmjTfLijnoz4YBU/N5ub7LYnAYOo1D/0UCT5CAP4evaKvj3mkmsDdgAdQ6Pslfr
g7sYk+cY3iY9TvW94WtYDf/p7bg2pKkiIIo1+UekbhK9pdFswSvhJe/TY36+PRkd
FKBTZtPfIFCEsKpJwfs4SVBeJWAM69jXi0NLGcHoVpJsJ+N5F7/HnFBrvqv5/+xw
yIfGB5BmxmkreS21772vSq+UFqkMu1eXL5x/js82hgBfeVNf3yOdgP72wPw04mFu
z6WDIZxHh38JiwA3pFa1m5KoUh6hf6+dMvhScr/BV67sIHffFAoD1yaBRS0Dat4l
lw29B0ox3e7Rxb2sliMu3UUDyMG7oQ1/CqJlXL4lw9mNLy/6MDmknpAXKz5xJiNV
psfy3zOYnOXNqKegxZTn8iP+i3BEQd9wT9QU5KKiWe6moGCJTPufad+bIxcCWj1d
eeZ1XtlWM9RTMu33FHElo/ogfaCZ1dYkcrBIPredjld8/lGxsJgWSHdvClyHYWwo
N4COGrD5eATWs63vqKVeGvxj5sdn91+UpRMDJH/KxJ9+W/bctmsFnvp5c/WEgmeq
/hCcxsqjkwzoTlkjnoRa8pyMkkh1pyC6bdHQtsgvZDScFqxxSH2pTHw2cyN0SfXV
IHT6tPYSIyF+nbTa8RHt0rq2QJALFNS5QgcgL6UOrvk5ZQt/wB7WaqjGVdz8pzeU
/ekGm2qx6PT9nR748WAEppVJ5RyoNVKezZCQTQQf7TxTzwjEEGWuvkSHebCOSakA
ApYt6CGHG+X2rJTkwKfOIe6pAKy8TrVcSFgSzsl9uFOLZcYhFyGYY7BZ+FCNUmch
cFdZHblXQi6vhZPsLBk7vnOEOxNavjaMd7mv/ei+Q9m/fVzq04MO/hpP3cVeYA1c
QGQnSY0z2Sy6FAVp0jmSKPizpeJWigKcfCosAGLIkQcPTpBVb9RDVytWYXSWwgEa
3SfiqmIprizl4OvsnykdyFXMukIoKJcl7l3Jpea95ef6Lzc09IIDLdQIHjstc2eo
opQoAERtlaKNZ9iHmOyi9aYL+P0GxEc3r2b5MiQ4Vm/s4BjHHIYvtUj7GTeJl6ei
kJvee9kXOSJiYxn5/tEsPXlTZa+y+4OUocpAcB+aAIwTXbhT6Sr95qYcqw/31yxa
8aF9Ni5mCUy+c5PBQWBdHwoC+nSL5eMh+yn2ZhfFmilhVDR5w3eiaHRSaofnhnpq
UE1djVGg6LwgJ+pH4TslyRxtJW4zpTwwTRqGZQIoxL2hPlUti/UC2mFd11y2yeMb
bxOsXOrK//NFl8xhWlg/0WeJ1K2QTo3de81uhj9UWSvmWXVlKisuOuF2D92JHmE9
jAhePnj+8nv+abO6yCscBi9wdNhcTfUJhQaPKK8FZALXGHk5Flg9JDrKg5sHux5A
NjGKg50vLYrUd3/Jk0IH8qy57SVmE7ri/PNZ2vAT/Wy3iAZ9StrBVvDpPwxMt1+A
3dKB3g6qEYv6zeUDt02NK/a8J6jsdVyD3mqDcu/hxSCliPjJPrI39kJZgpQv80Ga
qcwLr7qnK7AWkBspj6unsC+aaivNWxJt+6tIO2UYg4ZIZ7PP9ELAyDq/r3bDPX96
JhylmQOonIvhGvO0tI+5tkAPEr0rfK/wLsEl6tNaOHoQqa1mwWtI0LJhAcb+e+uz
AHTMngexFQ02qdtjQBGRubaYLP9dRoI021AhaKSjVuB4JwpMgWZMDQArZlI6rDO5
qZRvrF63+galL+4gzzgfR1j3DzQZzwjybVYa/VHp7XmKmluIi/onLFginqgflVuq
Y/Bl54PBSJjgjFaEdGudMSyEqlG44VL5aIiwBb5mgvNTCkOgX5PHsZHRnRWFq1fr
dnEKWuGY38rV7MPe4T8QTtF71+q7y9MLvHwFY2L8Mk3FEHDJlakmyQ3pmRvNTRni
RYWb1b1pi7rpTEE41z+yFssipUM38hdsW3qp7bYfiqAmcS3BEEGbznN2bZVSm6LQ
H1y4Q1vmkGk4n8zCRrTPbPr/FxC4XDfdHl5Rh60nfYZH2Y2IX2v0i1QgdyS108ts
EbPXzgyh8667uEhK+Frswz4Nc/n9u41lsVFAY9POuPJdsmACtMbY1FuNXSKp3GeO
Wdr/lGCiU/bFXC2igpNrJ9f//MFUx+sKPh1jqQtNU6MsVt5NuV9rJOkjZLXqoE3d
51lf3xDWScNe8+IamwP32DV9Ku69XiSLAzotcxp682zOKNm1tcffgKe/q4XvydFw
Ym6ZEYT2MPCeW2DC+wDnJRv9TUgfgUEZJqRRkhS6RPk48BBAClOiWNjRCLZuvj2H
GbUIOp7vdv+qJjdBZn7CqFoKyY96NHtss9vDWo/ThFjbQlJUeYFH+mMhqOTdItQS
dsUsM9r5MMUvD7L9KSqkVbLxx+XBQOBb0apFtdeN6s6dWmD6puRBRu6N1IfPrkOm
ZRiRDs6XvxALX0kseM7NZrnUXt4pGkt1Fnbp1T49/Qfq1tO0NtM3fsHZwObtRcs7
oZ3zc69Wq/rPwr/rKzWAUmix4P3fByBpx3eY6Zg5x/hAuV9W3V1bjZu1azAoF/qU
1h9R61V8rZPOkuPY6kiU66xE0KCWxs0mNRmftc0CAQSyonihXQA3YWsV6aDaRnG1
oocXpQMLiWCK4+oxyRl3TI7y8r45LGma+PlyhvK7zl9IxqxtTmKVMZbFUm7T0fS1
DZKtbQwd4TWWkKMudvd0ZtAgANe4fCWSO4bq4KL+AX7l7gm5mQNPDc4jfpzWe8vX
Vmpf9z7334TTZQuYAJZZyOv/xW1JMv1MZCJ+gGYlwxVhRuueHLWv6IL8tBvFSBNV
WikzyFP1Ec2iRiRwH9H+ARybqAc/z+BGNjojJWcCzDXD3QIosWthJ1+AAK2f1ST1
afKvd6LDi8vwQmOVw9bWxPMaVSKU7OimvJ2auS26S3uRxoPKfWaWCXG8LS/8zBig
agWXyur4KL+TWcvsMyvEbrcpjq223hnm+gToaUYd48cIpgKA5c5nUAn6Ub7clsjd
VwhiLrB+55tRgP+P3vVBAHSddBa5RGc7cTX9WOSa+kRvAg/c55IN8mUFDlvzSeYB
K1JYcAEhoUdA8h3dwZ5PYgBnCp2zs3ZX9lOMYfRdiuL58PkesrsYRj3bQCU3pBs/
+lN+GCtsb9RBMERx0shLWJfDwIRnMJwSuPFqgRU9Na2G4qQ/iHM/7x3NyxrMmYcR
tcdwR81aPBsU4K+OTpJ+9ZjV8bhwKPT8zhQulBM6D0cSHgzUdhFH6QJtNsi1hQkF
HlC11/4tHZL6XMcrw2qQSrG6HtismPYDoRpVNqz6+SjZ6USRBCiyVm+DAeRvtXnq
M4cPhClUsv0v/qqLIiO1TYhKffqpUVoqxu4LS77+jdfUodYJk3L8BSBOqbB+KHC8
x7LMR+aGtl0b6w+0Q+/r/QXdKHj6rCaYucFGnCZyvQ+rSyW6Z6bNX+DKkAM12JKm
TIxbvR+M6YUIndxf/64yesukFHi3RiaXT8DgtmMg6E7+tgb3F09hPHstHsI+LNZ0
6XdJ00ksZEz7xKrueMePKJQ4pFGneqcemFitr6SBhvoNXaNpgpHIq0LYZAfH07on
ja6/iPbiGr2JvQSJGe4P32CYWQu3y5htFF1Zdum7p9slfJJ95OwObGrZ1kuSIv4D
2VeNe3S75szs4O+X7tKA9m5m/pslx4ie5Z9S8UGaS+akVghsOB7M1dvg5kE85XEb
Z2Y48fOVOPK3YnrQDEwnLB4Akb7RngR3CAwfogz5rNJAoiUqNaBFFwL4zd4WRg5J
vq0Cv4/beBbn4ZUaA1sG8BRYAOOuv+/rNINVQy6iNGPPkehu4WvPU9741LBFk9ZF
A95RNQ8igQy3oWLE235CuV2JxB3PkXQ7TIqOeBOTo59vhQYHrXcRehRQ6nEZwWEg
Pojx3csEOntawztYxhKQp9DJeqoShBc1sV32Vx6IFQfq+erV1DoA6TySuJDY5s4q
kJkEBazZgwYiFWyMAp4wenb2Z7zwoRlP4qYAbbFZE4ockltXo+bqdSuybG2i2Km3
gUz0hDnjsq8TsgcEr17XzRddqi4Hr8U8GgyVQ7NgNwQYbDqNuPhe+k8fH0eArUJm
vXo8pbd/JLG70Hsaan1sCg/QFj/Xmpg2ou/9kTUqCGZ3QUsFURjPOPt67FeQSiUv
`protect end_protected