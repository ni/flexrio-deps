`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
gMcHP74wBZczB0bB0IzoP2xg5wC5NPjD/GsvSQ6VQgzYAsanETMwwsWi4yhFtJwv
5kY07u0WerSDf8woJ0stqW5xF501W3JLIS8KMiCOd55RHBOnavjYiaaLeu7oUCmB
TtTS1R4sO325rP2zOn9YwRbyyS5Ljn+PzFZZUmkt5xMca3p5NGqKtZW2dV6Babni
5HlLuF20Au601B75m2nv+ZRoGSrpkNElxoTibONmX8gBflpIVE7BehhHwaKSucEF
pp4QQ5zZAZjEC6aplZepouGVggAulz5AahlX5bf4opOVlB1J7IrgyjENtw6ysQ/q
DzybQ+ipztSXBGhmcCVU3A==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="jAI3OJE9Sh00Sic4PtM/KZ4WjwT98XM8AMZrZsQkxWQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hyw9IrFLPQsjvXplweG8O0lkaSLBN9Ijv4B5VdTRt6ipKJT9Kzsb5LxCKvkQyF9n
sGPOd5i74hRHnkHfYISGkfxGJCa55ieOyFShOsqTKRLxclm4oja9vTIey6yFm1BZ
54IDCG9h3PqfDiTD847UCSMRvFssyycwv+BRHQMQlFs=
`protect rights_digest_method = "sha256"
`protect end_toolblock="BnLuc3jxknmZOyxfJK70E5kp9u9O8IQ8cgkXv26kHA8="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
xABArkLxBOK6xG+7CdOOiGu0zbCbHMrEntFfAZEE/xRFxZaAZl1QLkuFI77OC2KL
XxG/mrHJzO3taVHgwRXNLDdc8ePbxbAiQfzV3NJLBO+gsBjmIymaCa480cPNpHLx
OODJjficJi5nZJCxFgjaduaCEVuhi6xstyfYa8WAaKoggUvzhYl23TQRwreiuVxF
ENzWqc7FVa3y1Cs3c2RHAWy7Y+hZwgRQEAZ1KzylG8Vs/oJ9lMkltz2QsF2fqqE2
+BwfrZYl6OwNHCui6HvQg1XjDj5B7fAie5BZ2S3azrPntXwcT/daFgymZflo4np0
EdNtFCC/BsO8cSfL3Gc6wA5dZ5qOAZ8EgJDMYDbdUTgz5CngGT2qqXhB+uDmJp2B
/EOiDiPAtCCcj6BpPk5e4uvMR6AFq7bQ0jQomiuuyjmOXL06erqc9lKW9iJwCU6i
MAdjRog69avh3NNSqjkOw3IpkRyUdFbZUcBuH5D663/MpUMLydclPp/vtHvAJeFS
eikMfRcRfqw6187KJuB1G7A2reAtNkdp7HpaK545kNxcI257sDYJelWCdyOTv06h
ZdoAfL2Pghdzp4Jdn5a3As5aH5c5lf/svdl/XZ8YUh5yaKh4MJ7/s9wQ2cjAfmkT
OYNgex1bLcfA2P9NeRV8sJycOAmpjgg7dK0yV5KH5CtTVArAzaauvZ/AgbA8qEcu
gchSzz25pbcdv1h48pflWaJJAA/SIIGxZ22mjPg6r/bsR1s+U3LrxI3jGbyYEhU8
6bLimCC3B8IMUVEjIBFDq+YD7VPa6tEkeJsM7SCkuTgfQ+sPxE/3JxiY1LLfkuqR
RmZ/2F9gqasulHIM741+r9mBR5Z0zn7Ih5Hfh0gUJFnRsXSZ6NrZM1Fzt+fcJiy3
rXmlw2YeXCcJSJmvnPNT6GNYfBkV49hqJT1gqCgWWHVIEFuA/G5CKogaYdX7B9C2
trHQ33wPZchaLQSzO3ReG1k4xD7nKsWI/E83WGakiDH2yvCK16d6GeztRx4BzRJI
lhzqP4NeVudGbNGw1Au7aDndWhouwuj6yOS9kS2+dfDQobhmyIqh3k601QnvGg/X
rF/Bkw/eV2anUCwBL41lsdTc4OxydB10UXDelcZwJNrYCvF+Jf2cfL44TP7RK1qX
GE+OKiOVBwtmY77JTV1PZPga+YwmwGoLxTKKtu7d2amV+oOFQBFFNuCNT+tMjcaP
U3Nxp4dN2QOatUQ5aBnrhaShQaDoE5C2fKrMbzHx3l6wHnh1UMJ5n9W+Q+lzc08P
WgVqbbQ3xQQacRYKJ36b/8KylLs3ths2Hf63lfug3l4YKkLc+54zbsmkG1CqnN05
Lzrh95USNYzgQXx4+WB31Ofc7tm+17klQCA0XbZV/vg5H0DFo6ZocFBS2r9BpFTQ
3jEN4D26vuAL0lIN1mSRMC4MJWmZGiMhuV01sVN2A3cT9Qv6pKSvb1m3DsPrp3Q+
FlAEQXwhlGp1jC9t9qU5eMbaQNHNinG86lJmyZm/KcW+luKrnTrOgs432iFKKp5m
jA0fkQKlbpAJb2RwKLogIo0FbKBt14BAQ25TetA+yZNIm9rdwrxVb73fTvSZBbaF
cP6p1Uq9guwly2H1YEmhM1+COTOL4fYfmLqamLS5VK8uvnr7PHzq61Tn3dHo/eP6
vnK56RaPfS29E/hTzyFzUT3PavZ5MuKecpjNNNWquGDjIhNioaHjlNeVvG382BIl
3BF7Sz74Rc+GFWGMn/vKmANFe/IsAJYxvNryzEUoV0dAYekBa2o8Al1Q/Xh363dT
1qKxPGFBRB220VrLfjWPtL1779AYIx0G3XfTDGHsbnP6S7MDwrz7WPaMJ0BG+Bqd
ZhHG0zYy117oU36DyShJH7Q7XovMoU1BeSS1VETn598a40QaOHeZpam2o5qyp5dV
VLxe0VivVLmdGX1lqucf1iTEQ+Cnxkoe66d04tUnCoYvGiiTapeNZi//ycopMpg1
uo+Zl/zGS3U52qN9jxTM+9HQfkAA3WEFMkdxZ/WBPiZVAtNKaqnWn4Y4AO5WURk3
J4cNqbNzr9XPsiaqQX19KM4754DS826KzQOMDE49DBE6pskaArMn8iJmFREO5hW7
E08BY5OkwqlgvibH823VImNBBO5bAWHv+pJMQSnVTpErl9o5ku0oyxiR7fxzWG0b
eYm5nbNYdN1qQ5tj4oDA5+BUDbUKIxDf/YeFt6fKff28HHwHJo6GQlThQP5O/Ie3
jMXBkeOpQSafKwpxgrWnrDh115hT6wQDuGrcfmyhJtk7QnrUnIOps9g3DvnqPytM
rSQZzt1xpPkgYJ7VssBZvvxyXqOgbOuEDUj6S9QAm76POgC+n3r4MNP0Q5zNcMCl
vrWnbA2LfEmL+BvDWHMi+G/ZQq6A37lSGBLXCXx+2ZljiqEsDPCS0ZIaLJ+bboxl
Byt0DKwKhEoCN6bKnqJ6Jj83czZk9mGXjaHxnU4qNNZ38R2VZXuZZSvcIZ1qYF7s
PiSGMwUEnzXhhhTYOpTDOfN25Q68N1K3MA2YgsQDeRiQKqRAhYIYDKEw8j3CWGz6
MgFe4p01XoDiWx+B9Cq+w3ncQRcjbVdVEt+RQ7fJuKwCzMDMAYSV3z/nXwNheiDe
vBjim2jL2BwOdEje+OejNRKXknbw4MsT/hsGq8YvK8qnISKCZsEmEw+7+oN3O0ep
/ghh0iF2yYPOy3rVwqu39qknjyd3ljSf3+LZgAcBixLH6ClL6AWNQN6mkM9CncC5
XfBmTXz3h6nilq59nu2smnmXq9QguE7jfeuPQ16sEEN/HBdVIr5n4ry/n9oiIC+M
slB2q5LVSsYTMGrVOBHHcOvYHQ2OQbOEP2I7UFwOAddVgDAPQOqa+PL+5PAWo1yg
8gWye7bjf3FGOWhso77Avl+gQuTgkrJ80EiaWuz7Cktq+NAhg4F3jZ4+vtCDdw1J
nGzQrpJ3rpmKLzIqQEPRbqnyku2U5gGrIQ+sN21rFi1p/CV6DVsA4v72OIwZufRJ
MgXVZHSihAWr++4oIYgylcF4OlzzyKqWON6VN2B47U9c/ozoDV+6GuJ9eh+NKaCw
hfeDrgT7s0UPmntdYFFxFeAyq2dYBSI+TcqwlFAlPAh2nrBBt8lkCBEEGBH3Wmrh
cid1lEX8CJQnEQBXQ9hEEqoGCh2zoWKaD6tHt4XHNL1tDxQSbz3CD6OdmRwieMyp
3yNfykrefcdm/RxrjXBDeQ5UbmKeoqoXV3EQWUUZOC34+0wlQnQJyaE4OJt9vlwW
Rei41ikyJ0vQE4eGjyqjh21yCXq+PyvHU62Slpny4/C/u95AHjjNE+tPbVQqy0/w
IZFzzxxkCjqUml+pDB4tAPocNu6AgYgjmahc3mjUMEnz4W+4iQyJ2FK2mjUQzJe/
u9W7Ins80dZeLvMPuqmDXfzPwbBPxMG3GbCPP22w2+5W8LOfSQaFakf1lIUrywmA
JMlmjAxS/vvQJglbltoOGQ7K0cuL2Ok+glOUx880pzOkojxeonSkCwswk9XoTMNh
jjZDEgfRusnRxI+0UYBj2s3TVLsCsWIQTyESb46wwKJC7VgATVLiZV41bTwhv0Y/
SJoxPIKluzivYfV9DJAaycDJT88ZJXWLbn2rFf842wOfLceoo7Ais9ivEbzy8u/C
LmVn7LAkoIClQxzJPZUCSR2st8ZX1tvByLfnQpUrAIsfrqSs8S7zYnB7M7BvzyXc
ia4p6BYxTEHFMr1JDCRVJLlx4ijUd6ZG+dTk1LUxeNoHNJbQSN2FtNhWfKclCodk
xuTy22MJHWVVNMIXuZy1CuKGu3vlXyzGdLv9l2JwPOx7++otBnYHSuzf5VfL7AkO
I8iUxw+yeRuDTHE0/FnVcQgTTE9q3ofYF1zA555Sq98bUrhDXxoY1Vl2sByxk5Og
vj2APeOvTHfrMZTh9YS9HgCjulS20anZ8VoV4HTmaVlbJ7oyIwlWi96dquWoCE9G
vBwPhTOBMKaOMuZ5Pc7SAVfaNgd61SaPlXu/HPQtki+0EMfdfS4K5b6qWDQEEFS1
6Qel/pbYrMS69uCxFp189pOAj5garD5KGzk9cwut0dS9TtOCSIIxCaoKScwiZc3e
YjBL3n0PeMuPeCngHn3nNxvC5kdMAr5ZfsA/F2XI743lTOZljx3lgRLXJE5CKaMd
hx/J/ux0lRDEGJkAvYM3tIj4/mI2Q1P2lGnOlhx9IRchmjudj9+91j9eccSWWUSE
4p1UfaCwTIs8qV/3oKHaxvUGkcymo3SWXYzPWGQ9NZ60IErPA8DRraaI2it2B13W
ih+HGB/8pHKEDlRZ0+LoEYrSPAy/ny+C7sl3+apOPutk2bF4eyzc01wrrs9G0/It
HX1izg2reft2Th/zwfexWv3OW3HVJLLftE42Cy/9uOKr5XaEBYaBMvXwHkn7Wehf
kNVIjNsLcoT3J+aWp3qK4tYutJ2uSlVGZM5FfhhoiQLgOZARELNZaOOsvYRZADCT
YqCb/w+6dYk2KdqpzdgY7Iw8N8djfSildyhX/F9D9xZGV5xErxv3TxBN0OM+QaF4
KT/V3FAZ0TWzSmjP/aMmWmYwaUB+JLgdBy07rMFlBTkKqkRCkObbEYtbulaaZ7mR
8TY2lXEs9HMo1w2dZAQ2Vfz5HLsuyNquM9cNZbx2V2hvh0PcvAu39do0YRhWDSdA
JbFjRjJMSlQemgJX0KN5dUAtB47gNxe/9gu0zz4AygOG3vxD3/rHMkXLbPd+QusR
gdfNvniE7bPYzz7UiBavYRRV7085trBtWT/gRTj5B3vNLXMaLVpO0RLVXA8yp16l
56/M71/UE8mXr0qGFjzNuEgZlnmkMQDTmMZvGaj4rtWw1obdGytx+8QYhN3PhxwF
/v4qq+liozqgBaAMSqu1UH/MNpNv61gfqGt5MAYDzGFjxDJDgEfiNe3c69TXCZ0O
sX40da/wvoHSj2Kdm1/zirUsLDQzo34hWYjB1N7NtLFaB6lXgZ5AqfgOcNau3G7j
ZhcRwI+HO4hp3LZ3UWVKgQxbXEVwPctaaArGSGsNTLdF10HVlvltPFcCQm5GUBMu
B5O0gjSQAjHsYQLjZpDaGaMiBbF4NvqQSEwAP33x3IBWacYg3mHDjZjz9yoSOonE
Z+mVn1DNXj9jRKG0XVtabe6hjHLk/4reLttYXgfAUjAHRw7Dz+D/zvfRfZauKH2Y
TNrinN/RkSS7e0O7Q/arEHf7R6JpoTA5lbcI4nzg0pD636E+ZUHPNibO+o4wfjcL
hoq+woNLNa0p1wTcFOG+wAYwBGbYjqw+ParzGcWlKjkmV2uX9hmAsRrwchpFG0qv
H3b5ZnPDWneMKeFo/X8hWkIJX01O/Eis1RsVD9Ao+Lm03asc/jrOVjp0iTFTBUCl
eAewCnrHOEWFgXh6noKDonB68+PorC9I8qOMEUYAOVkQlhfB63eq9qU1wZRUT9kr
kanEF1O2PBg8+xxF3n7wvyciRf35lBzbmZsvpwGp7jOx+vGnXq82MU6oYXlaLQx0
mOLl4hVKJ7LUMxENW2yG76NhdPdpRoDtijM9z34mBd6cJfhjatIn8rsPGrt+CeLn
8CSBt6tSNM2LOzolY20h/206fjjQtdvIYSkYzFNgDwL560xEb+0wLXm2Tnk/0ROF
FC9nZWBULvjFaD9tYDvJkNZwgA0DZWvSX03KRBvQW6ffx+lDu9UyThUsgGT3MQQK
j7Blfg9CCINkaU3dstkqNhI3sPLawH7NUf7R5Std+2pcv3xO3rzNhOXLO3R2LA5o
BjNRYqOT9xBvtKwcH/TV9IahQbUJbMsaiEe0rs0kbd+eOvk4kmC4Fwag/Pgv3RE2
VRJSwPGiKWkM/0bSnBGxpN3xrJxmLUnZHz0AGAo2SLwz/NNqCgQdT+YGG7XvRXoK
/uK0iRb0KtADdRkvuXqdovo3lbUJXqyP5xiK0mtEpR9geEvuw/V8kfA7gXQPDeXa
k6lqZFPKo/kKSB2D4sr69AQZTO55gxpTBAHeWIvvrrTxacgDPfzivv+UDRv55eVP
w2Ng9g5ISNhX5OEiG7ShHmKCNwW0s6uYkJBzofcuPzEjZTmD6HMfRlx/AoFpZH64
S3FHxXI1pFuScYLMkYRSI6Y2BNmqFtz1KFgAeGk/PUzEwgfNViGS9ISASzqljowd
2IjmnsLCp3wvL+Mf0CF6/+vJmzIIjYObrQpNqiCH7SzTyVd0RAhZKp1B4dMDVgR6
+NHjNWz3NMEl9tvNrx1jSUnPVebhGpoVgSzI5gn1k3+tiICOn20yTnvJ+UOI4zGK
01ZoUVxqDj4i949IKxvJw1lu+GyMWk7ncBpcqiXdKxXvutnDL7sMB+Uf7JlfyPIX
kMYuKkrRuBX1FFPSv2CNoelGAVtAlZ+9YoBh0WxtFtzMfPytQFJc9cMWzk04gAeo
xo84m6JeU8Ofdw+DeetxlZUHsnWAG6iyyDx8MdI5T0djHG0MN5F5aUZs6jqIYCpS
kY3zv4FvS68dP8l+hckC8C9tBNpc+ZYfYRIyOsk7oO36CqfklqqC4m3IvlXrGY0s
+mJcf66ElRlshujT5ictqyE7mDSCU5WxoVW2MX6akOlft8BuTUpFvuT01WKiXvpN
DDhbwWmoprOahwd4h16n84jOMqZTQwtk864zowt1hy3guHqNN+ykdZUCi+YMjXFr
DqQdxMfmV8y18CLgHAFEc3SMn/v7aaszGjgh1dgcuA7TYRxROungqcES6qGpeQnL
w8NYiEr93s1wEOouxwIgTFxeO7YSIlnRYDkXpY/NIYj4i6JpZR40QK4G3OjYW/HJ
5biO1odwGZKD8EWU51YsCAr3O1JaIg9sPdiAMPv0urRTIbAeMPaRFmUh9n/2oZjc
u14Wqh4h8ugObdVmQ93lh2nD8kbi6vT7NVeqdjYAVJfEtAhCLtvwiuyPY7Dyr8FM
ywktDRfzEsDJawkxuhSm9nG0MKdDelGtV15w4yBRG7l2ATkxfOXcgYJ5F9GUH8xP
eydMSYLGJC0sxWUWnblXCbRCf0kR+pG0tIn2dBom3QKkJykXfR4uQvqD4hjx6lKY
sPTtEjDqIPnQmEUKQWxyrcXa5RINFlaYMNWruSzVtxpSOoCNucr0mnJY3kCkre2E
rtkiiWFEhCqBlx5USHG0cPbGsu6phLzMkRFCqh2y3bkP1q9nBl8v71drCWlWne0U
/C8UXwlmsBzoHE3NtrtwlJgfs+S7D5vH5DrH/K+FLXulQpFh1IpgTsYJpbph7ZWb
cJWKCP3ML8iufN9oHCmsyBbjAVglqW5Hl8R7TMsT/Y4ydD3DU6m/Kwl0RJUyoblX
SuPkRU86tSqjxvYJ69vzKmlsPmwtKt8Tt0j6qvDWU/hdKjCQHtDQLWCKzIYOugW6
9X1d5LNZRhJcY4MC76Qq2Dm3K+0GM6Zeh8+Sj+VbWkvLWzavGSMawtJZwzugghIZ
rTm266/DRe7X+C1VpyxFKTk6RiNVVOlxG3XLI9QXlC9Jborgm51ylWfUGt4H8Ail
5J/64nM6aa59yym0xo6IPXbcNSlqVmsi3eWxLCNqlTMq+8T8kJDjgggvMB+igGab
sHrZYNoFM070/3BsBQRZUVL3bwSfg5w6TMis/ywJCh0I5Kp53o4/MsCm2w2RuwSZ
H6bHoQpAGE73CYSwyFttByhCAvgikoGB4Dt/uOn2pqy2Wa4YPUE7QxqriRo+GYC3
1qiTK4Uiy9VFF7h/00Yc0XuSOdxTvS2omtN4gmJrq3DnZZNzZswWj2x6nEkV2G8J
y41IDCoMTX+A2Wo8F00k7YBjDBmNZsoDtChVBdapWVCndT6BmULPstjCBFI4VQQi
fxyZeIsJU9zWA5tbKQAdNUieSwt+iG7nJz9A9bsYCgbO8bo1zaxQTThzKzhz9qxE
WXkt+jceeVRaAsxdwPucbySahkAxtWhXtrzUpjfEbyyMVzeWKfYhNWxHi70JQ/dX
0mkbSxGGb3f8AhoGhDUDsrZgvfFtcnDTcTAcpW886zZ57RMNIcb+mLthR/Xwdl3/
S2flP1M6uFSf3i6bmryqBXFSfRdNGx+4Y+rACP6H3R7amogSga8YFbxk6H309UAH
E1L4iv14adkw9j8WgZfiRNLDnvNoa0GBUfNP1iOFMY+7w2W1ER9ie94JrX1A6d4d
KqkvJxFtYylHxkREaJW6f1IDmkXS0GuGGtCl4olUCmU59WFSm6m4EDGLxAISWXF9
yfx5g+Lecg5Xi+aUKyZN0VNe4DMiA8XM0gde8QP0hiEpJOzuWfHcmJihHf15N9GD
k+VAGGJo8U60LX+BED5YfKjrg2frqOiO/Ml4eOYCMkQJN6e4rnpbugsItBzDz/ex
30UR9E9SPGxvs8w7NwYqfLiPvzuBRmT3mZg08LBISmwLXgAjs5zLFBIH2NOsT+4Z
SNkJhDCSt5jlOT7NZZx9uXGyhBiM5Qzom+Sqq/157P2AEnhHmkAxGOSYruDs/vY7
5CUgLc0PfLK7iu0iechMhWjbBtjs2XEZZwa9YEyQ08pKvgcfQaA1Jvi79Z/zHkUt
cltITqLhKluoFkCEZyRUFLmzc7Mgu1Ul+afvT6bIL2GSTYNjSqvdE64G5V/ZKhH/
XoX2weGWovLB1fhimsuduwHlS1nizIK6xza5XEBu0n9aJkuVW0Hrgv+2eUPhCUZj
Di0dZ05sivcMzyap424W2sBvbKVxwI02syvL2Ow91KqRZ4CnBOJQ0i6Osi5+SCLu
O67mwkdBTAvK/K5XBtU4lIiW2Q0o37hdVdeaMgpa9hwy16vIr6/yKTbXhNkCZczP
9pBSOLpFgSb1wP1+402E1j6A0kJkdAPfwu2nOPTSodOtURgpK0HoQxML1pbg9Qai
IyOxZojKzRsILhjjtlHSHJcW6R1Je3GpOjKflWniEvs2fa6O1Blfzun9RfCwxLlB
dRtos27fwlLvWauhy9sglor78OsjyTUqONE2u+nyBwZiJNMsuLCwe9HDtKXcu9t4
II4qOAJ6EK7MBZyp1R1BDoSqblQBNvdVaM41KBIYV/sZhmr6SXxYNsFz9aQ6LzWV
WCZObQxEw9ILbtpdA3IOvrvKiiEFoclDIck0qYSQTl2/cjUq1HMBccGq5p6pm1JF
BNHXktxPPg0ZrrRSVTQ5QepZk0JyoDjqO/UhZHjy6ehpJzd56jEWPgl8/sRTfiYK
Sip4e2b9JSKROsDar3mY74vNARQSuSxE2NOhlD1AHZH/9Qj6tldRWtAoznP/oMiv
YbhARgtZcAfiq4qC83+mbzyUTsaw/811zhxQnb03ZHnlG3WLNvRNQBx9mh/qkMGj
rkcFthcDIC7pc9ApneaOmURot0nF9ySptw5KLUCMx9g/ohovCw1t+hkWVJmkj9cR
Vuo1slksNK1OmpBl6u2tV/T92aFtgdwHm5OFffaXjCak7Er0mKbSzy6sT9NTJmWE
zKHGJfVBJUAuEmo3kC30EqA9RYzRzMbWKXhh1Hpu9gEOMfuCn44/51S5QQt5LdJM
LDZnCKBtVqVPdGoWWInc+Rj1awF84av6scCcaCnJ1Y8MFKdMX5GYJHwiVutG01HF
zk9fGQ7Lmqwgm/5Xcbaxfi0vTNO6n304FN/bdxeRvkxbcTr//+KLLh85ubRY9VHu
Jqww9uV/Gd33J2xLuYAcz0ZQDvqmuifo9Q+3yKr8leCaF+KuSHx3SpbP/nZpGNuo
Mkii+LOAaoH8gOUxdpciKQHPN5ru6MOUxYdpFYT5+JA92UVn6Oamzvsqt7ybKdGy
arm4P5Xkp5Qd/yT1WWfk1FUW2jL3BXjYD/HCybrN8lOHLhhe3ixihtWmS7KAPM+t
t7H7Mlc4KLszzdYlX1P3mYzhZRP7EKk6Mt/5ZRe+TExx1fRG0HKg6N0d/3d6tZVZ
NEWZf143SH2swWSfpkhR0nn81MlKNL4+2LmbKtFiadfYKa1+p95OJD/cCqRvhFJk
N9tPD1xhUCPuLnPq/p2s6fWBxh4gg404g9rirBysyGwNwFCzO/oikw3Uz8OABEsT
+Gf5dZjUoq6xZnSSj3zaeLlKGK+KgcHYWEC+5zpR9TvjjOP7KKiJuIwhprrB3i8a
1GpOaSN8+n9Oef2dcobucqeAZiGVfCNzgs49Z+cpZXZfaypGQxP+sh4osOAkAtXY
ZqnuFQxO5qLZcohpMpmcrFcHX5IWNextS2crlvlxWv7Zq4H9GSdcoFxXCj+Vt3EO
nPClvBwg8eD+iE2BslSPjZZdIuOw+YPmRmHiPHmFsCJaUtOuHeTvsyELx73WaKNZ
2HWDnk4m/VQkoE04/HMRW9kz9mpI9LaFd4ZNlHbAHBGdtq1dkMFghKxxni8HGQhu
Z1OX2jzbVoYkNy4HwYcCiaL+1WD5AFvIo2A9ivFANzKskPuVQAE3onQ88rfDn54v
dVqiR/p1BmFxfNL5F0U+pnuogGAMQxMGq4+z+Kp7pufndVjWcI3XNGU313xg5GxY
xAAE/T/S5Gnt1nBWMWKadepRtbj/3x8nODwY5DzWF1uPaQRzzGM8axAPvr/u3osD
Sa0tDkMJh+Yh6zN6HIcGNsYx6Te2x0sVBXSl1CMBxfKTXQ1IMZRMJ//l3MjHAbD6
VdhiT5NmRdelUEc9Oi9Ofog2BPbo8FW08u1aun3BI54MPR0FG3Ms6iCdu6FpAugY
hn9t5i037cOpYaw8Wx8SZrrJZy8BVDrtO/9PlKHjrvAHaSgnPbhD7tu9bJQQtb0n
aTmqMtRqYkw38Vsi3Ln+v/SDnGnnLlrdFU8MGgyJ+cf8krOBHSHLhv+JGTnS5rKP
IfUEn60PgvB+B4fkaGoeOk+p9zw0c7BhKvJahQs5/HLheeH1Q+RIrr8JmjG6P6ba
NbWtQm5uoSJWESVjECjQGOyzfDeaDMIRIMDpYtrj60xnADwXl85qxkdzPYuj5zP+
fWPX5qdR3W1bIWAxuf1Jfg46riSxriVc/aYLHDrLYyqNZ50tw7S9Q63gslOX2NHB
kzT7WJLocfjnh+jtO3rKXB/Q+ao3td6MPqxrrupPwO7C6aMjI+4GFN6cVKj5Bt17
0+ofuOHGfqW43fpQ+GzcgYN0lGsUOHxLn4qJRzRE62amaZtMMH7LpiTvHpPm9f7x
tqVH+B0pDF+kXrXSC/hdwt58JJO4FrOXNRILs37nTH27pYWLci5gddrxoTk7mYXC
PCeOy4xIl0zamjYuSj0ciNV99G80fh3oFHG5uUfws2aRL6ozpCX6DertIO9gMPuJ
nADzr57vldnAblRUfA1ht4SnUnkS0lmOHjO/iLHOTaOcvaGp/wI924XmRDL9A5GJ
23L/bVtkh4bGqjCa6SPqmPqmm5ReFzNIALtK4/sgwArviqliT4I/IqyFoGozTE3Q
VO3a2rOV5CuZq2bnTYSW5jH3uU0rguqvai6p3TkdGIS/FSucTM+GyCt/wOXLQ/qB
c2SWcIFZlr1btoa8yScvFfDCBGYoHJpt/I6rE8+/cF3uC9RhdItd5OzjWTTRTVFN
52EJ9XgHJCl8Q2c9se8JZyUd8CxVDBebhE3abWhizPJE1mYN1a4gngVkl42y+MPz
Mi/HsVIl1Wu7pJJXQqYANbtCzCPgaghga96yFETzt3By4Khhd2g1zSDO4NNwuOeI
Mh3tkETDSdc2JsInofgG5tMmvycbmqsn0XlJz8yiYuFFqYvQUu78LgKuRV6sv02O
P8jviSttg3OOG+MqhfVzIZcrgTs/tJU8bCDtMVzyXdRXG4+lAQsymqKmodkG6Gle
Yb3hBsrp7EHxMABoJKi7CcUB59RDqjNVYwsANjlTKBFF1v3zO6qv2xf81Pk8ePxZ
rL0K0Hw+inFUjO8v5Z81rV/HxvdOv1E3QV4OWzQsi9r9U3naIB3V+gOuz+y1yeFz
2/hbvSIxNvbBwZXm+QV+XtWePBwz0ZCYzG324uLHjh2no2bVRvi39GEnWlcu2XmU
DG7TWm7MMp3S2LRga0Z88b3l1RnmSRwgsz9q5bg0Y30msZGadaNKKIo8IbeKjEv0
PWESBq7BmOKgjYASYCWykrE0Jm9IGVa15GxHMFUbEovgOY0EhvToidBIx28vD5lm
2nisPQ2OyVH3REnWTlDRMVPX5vd+ujx+oVZnCHHTk99NWU6n97/n2R+7mxAPPh/R
aaVnpiegSP7tfmoPf/z01FaWwTZIvAj+OEYwvYPSHSl1FLp/hUIdjxbCNxmeRY79
s91WLItW81bL9T3Y4uSxD9tPLS4BLAP9ThNVtd5+XkFXEpUGe9alluWg5fagpGYN
vk9jhU9dLsT5Or4A7+j8amQXOtR2iLYkeg3afVbS1fog3dYqBd2kQ4ikjDK5gEWB
8QyL9TvfzEIWMDgks489Tuzjyl4V03jub7x9Yr4Yxin2IJqGqaJeetRwnI5+s0bE
R/tp5CuGoBGHdXFd5YdIBYSn2xMadzyii/szcdwHi2YCAXhy7CJHSjHtdJeWeabR
RDHNsY8JR4rACOmwnHDxoTjoq00ydquqj4jYon2VLIEmVF7lwm7F7uPI1dj67O+N
fEAhgIPUeOyKq0ZKhzqvlzKFGA1y1ZTpsBPrM1BkzRy8FA6slKIqxzupZN00Sf2R
QW0RkGeZ1GWe3Unx7Au0ghhLsmP1MoPp7d8xB1iHLpBycMUIbdtxw4wLF91Gmx3e
gwX2sa9fIlpaAEqHTzwKQwmC0RI79DIctti5dMU7Z2Lnh1EBjAy64JIoMq5AUz8k
lV1PvoYY8ZKLwlf+booomUXZ/5gsk/w5MRP19VXBbIoyrKoIll8Sh++4zcB9uxGz
3/r5iOhxshO4Us4HemIHMOjaDsBXD/UzAEOS59BY05xooaTuI+YF1GPV0qCuYJ0/
k3IE4tYWijy0CtGhkyvKWttU1T1Zz51HJiWUXEzklQn9nlfpqs2mTMAhqpawdBLi
zVT3D4931HxHHWBSJCL1VjB5GrCjx02BK4JOBpLiYs43yq8oeH7WLT/CrcNKoSkx
BhIJzGeXAg9vlYVu2dgL5xKWluQhkmbPFodCyuIDZE0RE/F0HHWRx9L+9Yc/LxSR
xVjscVrHF9/bHeKl1S/B9e581aG+RxzO/5alP8DtjuzHt7l0foKZ5Wwm/QlM72t8
gRPbsF2WIV7VzDvzmhP4AFFVUlEUN5iAOP9r9s5Laq3ekL9YnmXHZLI94Fs4GPY9
K+9oYEYVjeki8v5M4HOExJuLoYm/7lKHRz26B2v5zz+1kTCPgAqHLlaRuUsnQjmW
G/CCE9V6QmOR7KkDk2OooRKtriirnhcY4fvZ4Yk4FZeS8gN5pieRP7JW5rHLLomi
MLJshZFmku1iYMFYAyG/RAk7E5Pc28IV+AdkEwNXKrEZiyZDTFUSc36AcEFZH6JQ
RikaCSF3w0szEJKldmXiRYt6koaoevBmpXmCbIosFodPiRnZmSG2hhCy+Bizlham
9So8VmTXePmHnJ2bcYZvdh6krWWdbkw1BsA7k5VbUGfhTTkGyWJiyLpMgIESdqcO
PUFW8Mui3fk2iXZVAslZwGbXBLHZNj8+Gi8HfxsYb+vUMMA8xYikcVOvL1RAvEZp
a9yptUvc5LdjGvyCGGt/0FQoqqJc2pKiNehZkfgfWXYnnxvgLR8TajItg9wjxMTW
gYV/4r0i6rpOoW13g51cC0WSlXYerKcv/fv/VPNP8TK+gRU+or1x6pdkrbpyTQUY
lPdiCPPx0SBhtFp9iFDPv/nZKIoVh7lCk1IEWOwX2B2TbveRdxP+yA6FCjHONWCg
zPf85F46PLpCbEj/W3Ioa9dwUKouv8mrYFYC4Kvw1KjkPyvt40vpd9IWAe01BZdc
qo4+lT/fx//T2dNuqoC7pV42mLZKgE3EfuI0DblTc0qMXyk+m2x6Rylg5ldQyEpD
dtVIfYI6S4uoIl1M5upFZ4dcBmnL6RKxLRmsct1tlu3JSFFaFK6fzLE0EnG3q8ga
NJzTKPoiRs+ntqP2XVLAISJAnR/GJ2vRlLzLxrCBl3N8RWQ0RtQ016tSJ0xeIXsw
5gfIqlI1rvAZBTGjd/pARZj62vQqbPF8eCHO+w41SMvAJHmGA6vOgjMmRdWcQxXN
LjAUHfdsbv8UP5UA0y5JJvCuDhY06xPW5eslH4pQCuTqdoRhD5vKQETd9Uy13MVO
IDLHYf0ZLR25pAao67RsqUmSXEmIjnLR4vrBgvAtTq6QNP7z6PPk3W9df+ZCVskx
NqAclOeIb7g2T7joCheOSXx2a00y3uZt65NfWpK5o/Aepyl4/KeLScnx8TraN31r
12rgJEIvN2/zj9NmP8OeP5yyz2Orjvn//v6A5d4naRRaejRSIZ+fL8SP1pKqyc0E
i8LW8PjB6zBumXepRTiUsw7TObzNayEpdMW1nIZMpiU6nw5nQXAdywpqy9NBDYkz
7aPIfVSAheKEBiUK+JcEcp0e7lLdMhy4Ka0Aa8q4bVA7p19IRdfnv86iSQvoogtR
rdEHpM57opmfp8CoPMCX4qjzZaHV97n1D8eBY1IdKeGdgMaJmi1AjpXE9/t3zKNX
SGuybgBPz4FBAnctKiJ2uKcd7Lbwsci4GUkAyvMqmMhOBPrXId28kkqq7nO3STWq
yHZsKvWdysDM6+gkOmNGDMMv5UzSwztSI5sY2psmCY/Q0KgQkIhp7e+s5mQh3r49
EXSH+NAehlUUelgvy7zrc7edOnGT5boyVODvdvsQ9HTjsSy0ge/Zdr/C0DfDHGlx
1BXhSckoKmM1k1YkaWTW5v7pRPvznvooujKXmiM2zGkB/a/xIK/mQgFDcloLPvfh
qMw3Bq/Ykfpf2h8MfHQmxVUfNg4EwQj2zfEL0pKufAgHupESh78XmBQFgMHa9xY5
9ax8fFpM/L1rCKH2t+9rV0chjrsWH5up0XnxvX5lZiHDECrHXJLYsxXEyEmpTI0l
eegn9DVwCpa0KNauOBsDytwzmKRThNs45GaBV8o+gxFyBSvzNJj+aUQV2SLCfAos
ru58hTa5sAfw0wf5OUJAoPuBQBlgzJnaghoXBOXHDU4Tpuc8HJneKJ5pYK1OnAbX
crSCluhSHhFjet1jmvx38CgsnPTR2pN7DQbvcW/7u9TFk8zMJ2sfEzDkFav4zUNa
Cfdk/E5/l7bM6xpQzirr+4KlWtTCcPGvjcUFdb5QkvtJ/EQ+/su/DPkkq05RPcPs
+9UIhAKY1LgkqGUjeaaNc5w8VFlXta2tU9iGwJcY/+MlqVILbYdI36WioV9HOXVa
WZxVsXKoK57CWCeml0GEVxER0kqODrjsr2l1jrkO3il1YA+NkWsjtjWbQd7jelzz
4lZRGN40Drker5T5YTPSDlDluEw0wpK9RpiwPH2uX2jgOa6P9kjF8VowZmqMIvH1
Cnuu4+7LIVORmCu+UD487cZaYHKKDWsNuB9f+6RUI1VZn/s6TRtR7U2kUli6cvUK
QccReGDeGbIsS3KuOQGTbzGNvdCo7fhN2Qmh5uFHsbDdy0ircB9TY7Os6zpjSLyT
0t7tgNshRXW1oYNamOX5aP1YGn4FEC3cAexUMFQ4GTILP44CsXdmpG97D/Q7tvan
dT2+I3VRIoZCmoW6zAWfC2HNHVWPgNcmNW80zFr4N4rqGymrBeVHdNeErSS/ZsT7
vpkwdCyKGeNl2FsYEzGK27u5Jw/KFfhP6zFLt/pJWuiy+ycL7cH2nuWYSWEUX1eW
hZUdAdOzBrWbm85kca27BpcQzabkCefOP/2jUBHli4rwTHj4fMueHSJcoRiHJf7s
y/05ZwJkHuetwpPuSV313P55/yD0kyRVcoDsKgtszdPJCo5HTgmHV4DNrUqxkPXg
MOCGYcW76EulMwsuoYodBi8nne6t7xAXJGOP35OHZRrIr2kbiU7VLbL4JW32vHcM
WMGU+o2xWjeSE1USvrUmEXiZq84M03RkxcRd7jsrj9lP3pvu93cAdYjLh6+3HEsL
S0qYXYmwFM9bOexwlUeU+NcZq6OD7pIccVxrtZwD83ieSgkoocHgmccixLbzk5wm
2zRwtCYKJwll+Jj9OkKLUfVPbEycl+SiVFFdzlOLazsHlA1/ZZvm1zlDsq9w7ptm
uL9LjERZ/1FTEtlWOtegi4W4grjhWVHfsrHSTIFXgsZAqBLsWdpNKf9LfRfnC/YD
om29dta/Ug/ZWWD+PkTn3fsa7x/kW47FF8QgXeplPPPfhk3g5Q2Wp9RtUH05OJ0O
/Gwh3Ql9ggsje1Mh2a2J1oi5jjLUj2Fnko74piR1Zd9axNbRVBdTpFPVh9IfkVk9
bMTJY2a/Sy6DzwhKdGEqj4yzejs0vQoaxovPhbi1IQveQwBosmr0BRDtsAEiF0nL
4dIz/RQKDCI6Vm9Xa/m43OC+1Dm8mcj/dzAYH6YoMrI9kvbCzSAH+/BmgCiea7gn
uI0jOnwqRoHyyEt6Jfetl3ix31O16urnDZd/MuA61r2U48rXfKj1SMaAUN1iEhI7
4K0rrI0AvhRECEIj6PeAwAvLIp3rpBgWJh7Iv2VEN3N2MVkvnERTFZEcxVZEGizu
trIUfn02/ZckWo0519y42C6QwKcRsYDJV8ik8W5FJEBuohpvQ2Yj9vZbhPQkUREN
QqBhyxQ0+iYu8s4T/zh0c/0mIX2BC/VMW/tOFm6Cp7YFC9TqqcwPI2+3ESK+iWDF
A71EcJ05szNRU8Jr/N5rS997nIRpmZoI9KzX7N52TrKp8eeRjp8jhdpny4qLcqzj
m4AO0bTiwsrPueM9NZVTv8yqbOnug48cVWYyvf4mlnno2lyg5l9dVt5G/hCZFwcK
aVU8UacsfIax9KP18wpSuQ5qAZAf0QzOC926haBscJlBV6T16PT96m9b6SCLqIT9
F2zWmdyO/4sb2LozXXUMdj0zxhMWftUTlaXliboQWAEJjYzRw4qp/wZcnccvASwZ
KV9nLpyGFF7ZrQdeRjyWhGp/r+TPgsyrDrPCjLg+VmEM+PqDvpiWcwRKrqTMURFz
WIjaqYtSLC5WJ7zpRWfMuuyVgu9vwz89S2dEetb6gIuOkz9U411Mwk/5+yKa29tZ
gfHRcJFeBsb/euvyvTqyNluagNN2MupIteHJEaKeRwAbHXgco7La1zP8cRkkLv+t
9wVj5jhX897J8AK+gt0lzr4UbXaJnR+9IhpOXE980gbqbONBERIMbnRGnJ9Vtzie
b8xNqNaopImMDqYwHxj4eoH0clhqZkUYlaAltdNr3uRigiPJfDzyLuViBKf38Tw2
MCyfnKeF2O54rJ/mYP5XAu7jOkab0lQbp9zHwDGBYZwemZVmeBKXVrDP38Mb5bo1
7wYdYlhVFBsvHOkMYUrrLvVqWhp10WbeXBZFo6nLC2xp1USXsk8wY0XkDO+vF1RE
dJmN1bATkbVv2usHxn1+dy28VonzgiEKJNYN6ehpGgbvSCEUs9oPIcRcmOEj7EuX
UXOq/qfozx+qRYeovb4YeHpGtiONv8ikcWkTWorctfXY03aRAGY+91WngjbaRIaO
ExOoFCbvCGz441Odizh7X5C5s+08vRgkwv909MBG9P6t1zxUI85r1+FYaZSYIKwg
HG0HcxI2z81XxLHe5TO/26X5Tu0PyKS9oAdUE5oNQ96LPVExz8qG0Qb3YHklU/s+
gj7Ef/CeZiP1wmaoXu83Ya0MNKyXA+PNn/IqT0HBh6JvQkJIcvTsD8pZCXcicrxg
FqulQTNk9Qs4lQpAkAEiWhxY9M1L44Ovyph1bsr7sMbudZP54VVuQPrRzlfrGB3F
2S3aaqkykjvhF/G169MIB3l5eQsJfyf3CmrpvtPCT0vIHBZJrpnuXG+IyAm/cE99
GU1SPpHB7TH2aQWY7DXr0QVM1vjrCkcDUitlHe8AbLFyPws3XUjepKfEONeH2Noz
9KPh0HBKWSjdWNWSTZgbxixUT6M5Oa3Ns6v4QhbmS4imG9R4AXvKfAQx8r6cqdGa
knsBO3dp/iiY5yNJ5U0q3lgEuiLOGF2xyUmYpLVdF2iCh6g/UOjouyimWIcwACJI
wKMl7wdfyo+TkDlCbgwvvL7xD0WLlRSL7HKfUnr82Se4oJxrrKSKegaiH70UpDnB
zNA7TjPwbQdSmc5J6KmQCsyiCRsm4pZzwFlb/r7Gmg8kl4puXjT0Z/+hymbIZZuT
JFrBfHYXtAUBbYfckot9aPbGF12QYD+t2czn/IdzyCoYtOExuu9470OzwUorU4lt
FyIo7ID4Uk0jZQElP+qWB+1ZL2TQPiNH3teleKcDFTOzFAeXquzfev5OJrwhtXgB
hZG79SMhFNWE5LerxWIX9+uENBwigBuROCTY5i0c0w7R5tH9iWBSJDHn9fUiafc2
oYkvZmoOh9Z9ylWjx0nL3QD5feldoGMHnGTpqq7nWYLq8dLbWYigCV3JF9NhAr42
kX4fz87RMHe2S6zdLZx/3wnUSRDlGGgQvDEF3gfqQW/1BdCmKkHmjsB6ijH4/aQI
qCjpJ/veYMdvzyX8Br8YosPlbbHLGOC5GbiQ+jJioFWczpcDBB4KirEAuX8hBuJG
P3X2hDTEADwFF5T81M1s0DMfQWJifbYNTRVa61yAfoPKNp52S96bkUoctdsDXlzM
Q6lbb+5+rUam/sfOmL3xIipZgrytrapgQuoF0Rpr71/0RXt2ZTo7Q1bXhS++4Dnt
s0WmrslDTt56iwhJJrPDczXE2DRWsw5pbpkqKmwbFBEyR7E7J3nWWQN41ywwGg9J
lzZQeQDea1b7OnaszWe+5+7in2vaKMYLvkoOCs5JKM9NBGun5Pdjaj0fqIh1IGuY
OTXPYjelrMumuCuLNNV1jSPGvHWvLEhImy4VvH3MBpacZMc+RpRIWouLuknBDDkM
85YmZuSGJVdWxEfJSTcpN9K8HYQu3Mqhx5Tad/00GzYKTIOctWUn33f22edUbEFD
jhKL+1hcLiPzCvr7REeDsSwxPE7hxLptCGXlv7ohiR68XU9yCMKpTxFhh3W6Fp5D
/gLru2VLchWuGowTuNn0KuxhjE68PV2gsFCOYalW20IcVTJqN6zXvhKu2rl3Qgiw
RrZrkpF74FpvDDnBPHeHdjaA/YxElMN7Znx4N59ptA4S1dUQhFj1BwsflA89owD+
1g9FrpJrxBpPILg8zoX9mKimDnxMiTyLi2FIQXi9To+CAYdGh3J6d93wsrtmYPly
aJsFxiljZpdGzpGQGy+NPeWSASp5ob44jbzWNka65PAbNQijJZnk1/y3yGBJrlVI
JoubW+vdyy+6gDYMG5k4sWYuGVuX7tSJzxsJYbeiPDBJ4Q8QEVxJ/JgZWmngsn0Y
T8AmQeDgcOtI+RdEvEGLBfryqKUpch1KhIgF9wWSfmVJUInCnqCL3yzYlaTpCB5c
Z2g3KE1TnYSIjgnO5QBYrR1vSJSyylBy/L6Q46vKXTkttp3sMpy49gTZXUEHncxO
MPMuXF0hTO49QRoATbB1lRNy/jgBmAFhEstAoqy4VJwoqwKYNp3Gq453qg2Xxoz1
1FzXzxF1MaBdmBqu/94Gl/9KDp/8QgPE5fjGsHR9/mLTdVMi1IcjD8qJgKmwCBol
/1q6uuRV51MY8X2DBD1ZoyOyxx3ckE/FOpr/aYopE4psqvn3m+Iu1jqtj0Fmp3WL
+XlfD+Lfi9OB5U3LLrReRuZTz2ppwcwERnUI6sl9bGksyxtOAsOMUEoOnZVfAK9n
Ipvb+O5EiKzErkWGZXrf91XkvaNX9QFmzhzu7YAEfe9qDdioIaK30UZjXYg90rqY
ArX4hgv39snwLp7/Ea45IarzLERc58ANJkzEgNn2mZW6wpvMWsbYThmD4MqpoFus
xDyFBkY9jJs6t3ScxAGJtfuOsVHPCzDokjm/VfU2iDaXEW4UfnqVZjtX3lJ0p92N
phXPft8zHDMOENpsafEQGMLSOZ8ldL3G0a7TGFW+SWRQFNv7I+ahWbqB1p+dm2BS
Vpg7muG4Zsuxj5BskpygeQbbyO02SrNDJ/LE0YFrief4WKSCc80ISE7SAdx77jr/
rWEWd7qsXowpmr1ipjNAUaQJs0h8U0it89J3Wf02Y4syzjLVkgTMYxks0BzzJnkY
2FJ9DYUtaJSEizgzb67oDfg3Pp5pjgAsvNAHf3P61kpmSb4gVY/t+UyGppcvQ3lb
C56v6Yes/zDv2IT4UlPL+kRf0RvUQuSwC85Lwj3SESBlGq9q7JxUsq76McQ5Z7Kr
TZaqHBbXIkdrqLv7NVUcwVWWFpBf844ZXngpCrXE+GWq9rNL/tr5RZRuIm07SN2I
+MZ0Xv9dHV7DF8Ob1s4nRazgnl0okKLxfHTKdf7ECu3Cq11sXweNjjAM6CLTnfrJ
RZ8uCcEOG9sjpjs6+HJAEdqgz63TUaU7fM3YOBd9ux0STY8oeFQKSYf9Ay28ROav
NuLWZyW1RMrHZt+4IzQWpG4MSJCRFLbrtVi+nphrUVtZijM24/OYQ5NmRKAoLp2e
wB4RMeDR3AtseuLI2UN/2KBEZzHf+QDRHnjnw0yhpDwh7OoYzMJMUlDENRIdA+Ht
UZcZoUrnHYDyI/whD+H6+JFXwiTlOpooCEtFR3fBB2phPsxZSGy2tqBWsrEPuuIY
Bfy9/yj25kA+yyGBcOzwXXknlZAjP2+ecT/F+etASxgcu3lQlR+nVNJRtkYF3YXI
Cd3lGeKyRyp0/E5j0zqWJ2ePdjCgyuop7OKYq5GKJrwETESZu6y+JqvZaOIPFhCj
Nczo4s5scSwJSvJKWQN9fBZTAnCC2wl4/6PiUGxp2/bBqfIC34Mnzl5SYddkj/2o
z/KXTIesDadGXVz7+zeLg2Rhz8izeNzYDIGg9KNVvqE554oIgGD5ueAk/r539OhC
ENkANJAtJDRW0xixyHqbAWJVBdj66xQgOTzg29Gn9HoGJWt/m0zlhzdN0P1dSlG9
1RHO/68r8evivrx+xFEgbUrGDOkAF8aPCbhyeu4x6ToB6nVitKhd6IXopndImrXf
9jOdS5I/kHDbvEOvfJE9pqMQ2dnLFlQ9102OtmPrrc1aFhr1SEHtQn+DATey/Oq3
fpUXc2yoWZYxP0bxbyXFY68VoJftHoCiOI/p1I34Pu/H8d+GFD5ycNhLC4trYspP
BXbQWL+KTzL7DEeNATd0kGeMu1eofbBdwQgt1XFkh+YI1gNSn2QcXezIzecEr48x
/G72F95aOpJ3xqkU5zJYVnD5SPIY6a2k8oItpNwPe92K9ppwI8D7Ieuwe9Rd5CPa
gRChucnVK8eK7PDZaZ8UCDgxXJVN0v4AEPB+JZcpNnmMmScWs5V4B7fEkuHkcL/w
K1nJNUpV5GCv0pR8pUfhKEA49ZU9r7ctVw4iV7nUfev4dgKZGlMieMU18kyuEDcF
/HYmBRFWz9JQgdj/14QOKQFi9K6NtxIPt/zsJ9mI1xOaL+rxkdHQ+JXYjj/hrSJV
2ZkuX47+ZQEB3g3zSv2zswglfCcO/hlS2oeKb9rSGIHp87RXGCt2orNwXEIwobjr
8dYHLn3HJ2i0XTIONOCQ6Bf47nq3835ObGkxf3tOSlz4uAM1iFdeJ/qX/0rX/ero
HDZe8GMafHXi71KlAUB2gbOsP20qls0IH5mgNzKTexwL5siSkVG6EzoRGEfbwZ0S
Y758Qrccj3QAE15mB2ziAHrOrdDrvh8t1qBZBf9Wp6flEdKZDMSqej1le+95ZDWY
RU098gCFp8umepN0Of8I6Qvt/l91mR8T0pyaYPSaEUeewwzT1fQczTGrx9gmcMvr
vBhunUXFKDuUR45/ZVXpwPNlM8I0IekSsAaJWMb+++Op7M6Roext56QYTpvSvksb
FtnuIvRT7C4Z6cPgdIfix0fvfSzveK6EYy3+qDggiwJH8twSS6Z34tgLUb37MkSE
C5ppl9Q5WQoDT9f3my7GlpYiJ5h+dpo/lmG1D5g6anuuUJXSp8y6Duncj6YTCeWK
ZDaIyPcy5UuK5qq8mbnm+BzdAd56y2rEF9MV9/piiz1pYew1cY3h7y+7O1U+eaJ+
3I1W6Mck2fTNPCCAurHtuxX5y/cn3wh3UoxOgVWF39Ic4xNtdIGWBZGkc8lgkkgp
6t2ur/PY6FMYnGHrqWxQ7nTfXt/nm2pJuoe14Ba7GTyfNXdZ+HDL8IeUP1kaOlg2
fvV5nYOYj68BNXGp1ltTCF3Wjl6CcU+OgjeXowuxyIIKKigr62FYSwU8iu4WZgL1
AViNA1fO+aUUvLZHsTC61xYt/bj/X2t26Ujjg6Dj1zGay/gQzlJZ1YzAgAHJ4O4P
eIqMHq6HtSuW/Y/VoeagF6xYXNMCwJcbujrzAo1y3osnMl5QDtnfJ93TNPGK+VSW
8wYbfnhfbNqO7rbS0pwHgnbgGvJmhm2sfoQOztuHtuPrbQfTeIUj63tDKd2nIsyn
lvqadnIK+dMaLXimVYNJIpHkovuKB+rNwJS4PGHII+8Csf+62KxKHdFl9S2HPhZ5
mG5HvdimMv9zoaVOjZaKSgMGOKfvfUvAoJ+s6Xjksp2vfWbZt2s4qellp8MxdFcz
sL6uQPpWl3iOKyQwWfV8FghtkxrsWsHaxCY35dyxznBAdSZgVqwrHKMJmTTdz4Iy
dlz4W0qFDF9blVqbgYKD+LScdtQfOLnI0LviUlfqZRn//MM1ptlFdQoIOOXoQ2xg
Ub/GrFNi6L/aT1NPDtVoOcmLW21Ezrv/KLXl5VRpPkvrdzZt/1Aems+LfkEDif/I
97+PNfFhNua9U7K15snmnrQDFDK9h3cuOa4xajzopvVq8h4cHVLREzNllNS81Nvb
VzSb1W31xt6MJkllzbbj95icxjujtMvjAi9WuF6FC0+LSWuaeE4G2gNUKf5RoIrb
x4EFFAfJjKLQG8+iFiGIMLipOMiSNj4fZXwjFowjBDshyelBrpyzdcaSEPyQM/ns
YV4wo3W0Gi9USAa0VjiFXmVc+95Wzvnux2/C9k6Mk80JB6HKzQBLoN7pQtf4nyI3
yOBUnBeMOt9CT1cOd6b9JOPcbIoczOmU+3sOeJtBdSDEsjamMEdwj6tIPmlZIBnB
B3LZgcWdXtEcnoTXY9pd4qXyFGbBTRZzyLL1e38IGpqLpAhsCoMhuoQPvEHjTtna
Wxfdht+PJ3FrnGfTCB6uTY/vpDItbYIWZZGnACORbJBCD9AJgj+/3z8BGsJ36eIU
3m5573GxOIj6vcWBxry63savujpw2G2xEMBRgVzv/kuHatiI0/l2GjJ4PmlWlqC5
fIR/KzXmOCR8lKb/TuP1MvyraPHKoq0mIPyI1nkIwPjwppm1/Cnm0kUcT5ihoPYe
lQbLTe+6d0lyFF0VD1XhN0x21WhM/KVJa8CDt+pDKVDVVmQxhJVlCleHbHYmuXvY
BsOzOTX/4dMaQ322OHDCTe06t89xwjYzmNBTS5UXc2g6XL++1SenD42Be96H+lq3
QXueH5LOxSoIhI55Nc1cgMu5hbHASY4/zbgxrH1DVNQPAPqGGzHuEMWyC7Y9eVEc
MlizzYIUDutGC6LR4f5npQKz8UbP1BGjJTuNfY5QoIhzk6q7uhNU9JUy7CAeFQBy
x3pjloGenM/VD7ewrf/d5S8nrKNQbULXe+3nQo+OvTqd2S6S1v+drtrbVLyU61/x
IDpUz86CZ1NM6d1mirI29Y4B51DQ0UAsfuyhIqqKOgWl524fCmehMaf/Jr9g2+Oc
6lvpNJvM4GQrbLFONNu1K8GAk3B+As6Rj+P5y4xtkXuIKpOcFpZwWX99Bkhpqn/a
jy4DxBCvlWNE4XIrz89e6ezwuws6YgqdPozeRSz5AzXztDC07K+BL3e2iRW2HO/b
xM09lZJzRtALhP0Llyx6yeqaIQpwkpJCsOyBuAa0/a64vL8Aw+gEWEofgEEDiDz0
9Ts80Tc8LrkwVNHP0YzH5iNPSy/jj9mpyd/EiNmIHWwIQLf4eMke/hVQ6ZegH6Fx
iNjkT+rwLcSiOF9qmov0uwrd6nd9uT95dr+IlFN+GZRK2qb464fqLzlvuNbjjR0Z
fkcFSveYy+zYlNBpX3W9trj1ISzPno/q4PQcUDWh9j+MvVjD/9HHBdViXWKLVK3x
5uQOQWVWVwAfgMJdwmUO1v7TWAe9fsEzENyA+d5A22UZ9JFVl5kJP0yCtAFx7mPi
Z0oSg7guU/t6joHFM1F2APqJkDtygYnpTtBh9i65lwX6SomvB2L9IBCb/HbNhDA8
gx32uNVCgBriLTgCnkpFkoJkt/G/ICjBo1bD7/yZYw9AOGZeuZ3RNhktWwbqpO0R
q7WhcKOeJG8HGyRbwt2bKZ+xqE9ihmgJtNFr7qRIa8nVywdpi8CwHp2baXhtHMXx
0rR3tPKo/4Yla2c2JFpVG8KV3jBWbxPVIwbnLEZG8oaKsZneEYHAyIuJwLUIfrYE
Fdxd18cQysJCTuEUKM5SG0dBEzXF7h9LyygZakiXRoVHoEwj2CiaimHAsiJ414QZ
EMVH+rPzOxqelhmvpfWWbK5qvFKkD2zbkwP504xozSpwy+xSDk3Bua+UVlI+4Jl1
JJwvyK3lYNUW9H/ys/zHTzFp+8eAsRmi9dQTsR/wP0giUEUncz+i6dLkQ9QWN1+t
JovW6wnS7RUXEKVFuaiY7QfXCJ0MX21rXIgLPGpJifKq85Xlma/Ji80Y505GnMa3
zWka85vElm88LypWKelPJW4qazuZGpY1pkQLmP+GZ/MIOmVL3yUwG59wBZ9DQQ9z
o8UBGQBI1YFxPYsaFuwctYMUl2HGldWpaoGJszkVTz8K/ya/37Rv6sBlWpzcuk32
48EuU1cliwnji4MmvC7LWOX6pmEocxi8tlkQ+enx0iewJAYUzC736EIpMbg0uK5a
JJuiejMEiVVzo1Rkeayy+5i7MXG4WM//rw3MQCfIoHcFmYSCju0K7AFK+8WbRB76
vPdNnzd2cxo3ztDzuS8ITno0l34mmPxialwE6HWxZJrKnj5VipIoaiRPI0yFEM07
sWjFG0iN7LewbKth/2hUk3ka05T+ofY6G6A9RsYq9JBLYuLT3fEULPD1Z/GWkUP5
f4omiDlH36OPDreM7vFua+4LpPaoDZ5+SLh/VqYnn00nvRqlgtAi6r3fimYeHNS6
ugWb7LgsIm1jfjUQRnXRuus3VjaQE+VuBw0PQRV+0T6xI7HwEzK4K/s6VLL6OAly
h43kkgDu7Gxb8MjDebzirfXuy9EmOWESVapejAPEkCjKpAvPFDmScOYUe1xz+0Ed
4/JaIDqkQxjokwKLZ9ka6P0zihae3ftQAQildPCZm6sXTpcyanJDd5ZVWUfUTFAE
jEM7trHkzeW2QBq2FRZEPyGm9i5zZfaNn7MxZWfVNrO3iUimkiIt1Vfn2bGXgH1G
D7fBTTirjxblORQHKxVZUEu8k4mlNPzNC2M8ufzSpwG9m1Few8uBtPWSx0GXATHb
GU8K/B6X2eEklXiiKRNaL8qGh2B2GLZIOO0N9g2up9m7KFqnk/hhAts/lWV3J9Xe
2i7sQp0j/drj/qaQV4CRFbsZ3Ja6lj2RH5MbR6Gr8SPiP2Hq+AIKwbu9+2791vDI
Tavc5MNlSJftrXbl8poYppxjrp3t1CeoVmcap8ZbmXtF2jaG5WkP4gP6dJhT6T3u
dgEQo8Snamq/7eB9M2VQSAfVAa8x8X75W1dBlhWNlv7yinTpJMJ4fxPv4tq1gY+r
k9tu3nv0cA+PGo3vVqdMUgTc/vwSOTrf5Cozh0pWdxIaG7BVFRViFEB3b8LdznGH
sXJDCA7UeluwZprItE9Tzyt/zTWNwHqh7KuCd6bYBMaxzMD97nDID1PZMG2ftwGW
2mfbLFKqq1x//gYGH9L9eI6CGncLWxweg4MyltNMbA8OQZQrisf9j/z2ScsuOopO
DwMAfW7pMYFdVjilOYLsujSDuhE9e1Pxcu5DEyO0ePO+sw8xay1sH7xfhqjJRC+L
dnDlzfsE555ruway9wPjhThoO/ibVgF6gSxxPS+bURPDdW/TIqy6Jie8xsM78Lfc
+iawqixFP2t0VD2v//7hmPP6dl4fP1cIHAOXTivIQc5WZqMzjl8hfX/hrE5jtSUV
AT1U6V42Y5jDXqDI0ZRe8y2xvndYRzEB0OvQQbUmjNa9HhlOU8I49QXpiM8o1NSg
h2hoTWpzfHdWQeC6h2cb/yNulCe+de+g8t8u9XzcXR+rnuGMtL7LY7/Lo73RuvVt
H5ULaEDPWxqLsi9O7W5hEAYj9AXXpElaEoOb/9vc6+2x0g6gQvmsjtJn0X8uHZ8d
4zmJLJDj4GIZFCp6lpXNVa7s6EZLPRK+kf78vtWMTUKPlS4IwwpFbrX6bvIafKjp
JLrPs+AbIk7oIFJ86qjEwQ5iPz4/OI3A1fzT3W4pAnEDtRdjqy8VrJq2SHilL5aS
x1/zQCQ/bBVeMAxFmUocxVQTbzg3G7kHBIxCQtaQ9d9IZk5LE1m3W47htVXX5iAG
5NXPXetDB1tkwX8UX/OBhUMlZq5NUFyWGVdi3uPpjzCW6CjwfcxxsB9PnvzFtzKe
+7byvPbye36K7B0mXQN1exmmun6yvuTVZPl4EaC+mZrAE1QVzCT+OKmNYIH9Q0YE
0x7/EN+AaR1F7ZCbUPzsh5I0vqcjDIX7jq1ZXGtWTPPYu5F0cmMCkegR9Ktdc+KM
vKS7uQ9/Nq7jb8PYpcD4xa7iM7/u9lAJkXIRGxngHGAEo1x8ocwURaiMNlmUlscK
qxS6zYfmEoBPtLnY4qb95LCaLo016M3xhq95eBnYTQTRSIWEWLHkX1yUXhhwOTAg
U0tEPwMJjXzxD1EYqVLnblOBqvrkDTj80XkIjHmao+jDVjfYIMvDpCmu5fEeS/QS
aPTSdSINYwEZWDZHhC16iBh5wtgMaCJBKPUa1V3Tsq1OCIbj/dSCHubT5Rh8+uUi
cS6EdvTo79Ddd9s3TbY4oBaT9EWqJG2WR6Ua8H/LugiFq0R2iZKFF+bydhzu0QDg
RCVotYF5vjsdL9iwMZkxIhL8jcRZHdIqlSJq3m1Lp1MRs+ii9TUA9j7bAXj4NI54
5KVrQ191vjT0Vsm58uK00LEoMRp+ojiqtYh57rRvIC+iYQm0KNcK23PWPGlvdKtg
KDkJDJsdU+0XdGq3IOeBsUjHoPgAiAWuTagC+gRjwnOa2/TiZUuLvmDrEa30gOZI
UBICRg3WufdJQseZ2fQmAThiGhMmlKgKNpb9dm5yTttjo6IZyW2lyWvgvHEA10Vu
jdGDkZFGTAFq1tEkvY8DbvlC+2MZFFSZBDM65cQxwzl7m030Zq9KrYKQSKf+8NuS
IRFk2esneqXhmK9Ce4eTIHieQ4S79ue0nHI4qkt/pi5gyT7Py+RDDyvtJugKax5Q
SFxaWFGjxDiBRCjb5Qmd//8rm/3UjhwYL0u7RZBIRk6QvSjWBU2xp1HGlGY8G8Mx
A2q/lls1KQdvEDXQHRcljJVLqmEtJmabBRcq/Edai8w2VpexMe+JW5CKC4SVw2G7
5R6PhuJDpcp0V3mdKhBtbrXpPaf1u4NGEZKA22NhQN5Te0JqJ1Jo0/LWVgGloiTE
oySITifI0n+rAASYxt4fcWvQQ+H+eTrjZoEmtUDtSWtfmGzq9qJXck1TzHioutkk
OoclUU4VEiqeoV2cCmONHUzgUig8qPyvRhaO3sEzameSQDw3CFCY6+I69NkANrOZ
se2iTJgYFaIr3aq6vviP4uQS4RLDm5AHMcyneGsdZALcaGUXJlDhpM3XfquwSmxw
vS51dIy/WsZm+yQyGHC9MN4urZPewosWIgIZ68TDKr+UzbSobS9dVoNj+QVvonGP
XrUyd8pdLSDJWZ2cy3W16JWatqopHPQaA8tvQ1pjTkWHWLm8BpIi9gWaxTPgRbQ1
qX2nzk4YospfOJfEnKVKZDDGuy3hmkHYKcXZRPMDZv5IgL1RGiyInyROmm/dAx7W
LZFNVdU1T73Y/tsQ0+LqUHL6qdgnC9kM0oVvJG0f+qik6ADvjOLH/n51vnGR+10z
8S9g2+kqoGUdbJnkzzaL2MCMyzx/JJS8iIsfC0sxvWFoGjmaLaw70FDMYzWVkPjN
IaWq/y+h/tR/q5Pg2U88pM/c8rAb0uiHt0klYyTWsWP6p+2rJ6G3x4GKhl6UMasr
o4NM3azAEXcW/SoZ/in5v/cjNlap9b54Ovxt6hHGZ/Rx6ts3nnKSzwV8uudelYD/
UtDDEdWAFZXx/i/uhBEqT5RIHeTwBMkOrw1FlV+Ql9nTaZQqWdz8tkeUR54DanY8
Ro1IYgh5G3HGVtn2W92GmMIn4+8ad2TxglVk+QzwHDb05mhC0My6a/nu/3sGCkfC
YvDOq3q9/t6xwiQM8xeDBLt3erhhbjDQa7Y8qFoXiwThafC7DjM6fln0bcl6oggm
pXtcA9M/pGGxpYGaKVMUa3wGRdJTK2EEE7aI8c3e8jMcI/ePlVZssEfsjutiJGks
UCohnAsPo6KhogRw5DD7YJtqhTha0pnNEgFNPrK63qGQYOhKKTHVkUPC+NJzBlxu
7ZLv77FHraIu4gHI4Q5lve9OeSeRBLuHhkgzrKe3aCd5BdT36h6gjuOaqz8JS6KI
0eH/PWd677IB149PWaGMkP2uz2KNm2U0bKhc5vq7MZYPEjO9fcq1ZcXywxuyqo/t
ZqigJE3am8+6Di1VSUZD7LA9uyxjXjMQI37tofsBnJh0uRwpLMz8m3QWtr+DZQ22
3lVKCZKAlH5RM7YtCfQRxORKTQpLeKLMb9ZfJeeHO8HBtnO2sB71KLCiCX36E4P5
JSuNVzUo21tOB6Kk1uGT4+pL8qOCYxA2Iail4Y61BsfVN/INgMiYGtG/zF/zCp80
SXFC7oh1mKIZ4Xt60DHSAoENrANq6zvggFKcBY4p8hF8+ip9j0/yY9acBu/YaZB4
IiiMXZk3lq5sU5wdLfXy3j0xMJx4vN5jlNrF6aUu+3R9t+V2MUTol/1sVF4P2hlm
RbCwRlXQOOSE2/y8l2nDfDjaURqhpSRq8CM2YQOj0H+mIyYv8LeeNLP6FQb9Yv/V
uiHrThefvo6w2KSORsWZHb1H/5qwPb1jDyNxhNh6XJGQLvnX/rJCz3UZ9iJydg1w
gI4+NCV+tcxAgIbC3WXmulwuLdlxlJ398p/9PDGKSjjdd7VhkXpGMsrb+QsB8+c1
yVe5+V7KgeNt2zB3bA3qUWTQKGccIGCGOHW64ouqng6OyPX2tvloH6Ds7z3FX9HF
fpStV0twaSNBK5XWSB5s94XMdqpt+vs/gjOY65amkaPHaDuRHegJqWOIA+2K/01v
fq+9YIILNFhm+nSTnOl9pR2xlbmgb9E+DPS5M5U88b8UQdicikgAIVkJcPtix4SP
h3w0OxxmXihdYKs1U8F11Eaqq8PZKGzAy9M0JjN9wpDBG6YKZXPDq5YZaeg+fAkH
Zm2YXZUJ3mYD32bDzfm0ap2ikoE0zFSV/jBBiW6+fq67/rCe2JJPL3+yM3EN7nJH
xQY92iGI8p7teAJ7A/gQ8BHXKl4aOrN+tslDnZU0zGcCgc96TW16Ec+aKsGa5k9J
+qncXsoaSzMleHLCf/NlZpI7OL767Q7du036LLkNtcvY+BSpdqakVB6unx8MjTCF
vReHAwlMnxpYbZNLkDcD/0zy7bcM603SzUF1jqWzL7CW85btDC0CGgvI7YbS53rD
YwyXq1WcRodwNFDRRvaNweIhUpqMKAuqbiG1yxBcsstdeC9Gv03TI2prGy0oEsV7
mim59BZtwvP0arHxQP0vF7Ba6BB2VD5kZgLntRdXBOxOPNAH4hXB18+JfoBj8SoU
OsOp3hrNZcNHeje2GC4NPL4rccmYH0dQQbYi0A3njX3Qgq1r7XKb1ms/swbdEg/U
Kq1md+gtxZxUabst56pfswGilqZEX8WQH3yhnump2HLJGc06Jh3obZqGtGeYyiXB
EDrEmJWr3KtLsybksfWMMvSGqOy/aj+nPbZK0kY7yDAh3YQdL4QRCRBoh2/RrFkC
s2Iqk8N/wvmBjqT6pE4naohhl4CdB62vXKLUbTAb7Hu1bCa7qoiVbRz53HP15fyq
F7FrItt7As0J5rSBGJCoor7rCkQl4qhkTFPEuLRxXkJGl/XDJ9wGaOwetFyg6co/
0Ktx6cvu23E63wqPfqEwPqrg6ZTHvibileGORdZw386WhkZtJzIBQSgVaQEWQcd9
up1c9tu4wf4+D0j2foVkqcEAjtGJFmHCFdjJ5g7koT9PiK63Y0PXqWLda7NC2FtA
6pYSG8c3LpgZ6VJPhADjdGt+s8QvUurlYA1HFLlu/NkbBSl5EuutYrgY24e/Yb6B
qm8bhhkJyb+1ChsocwnMj/elB9ZtKqgcOipN+xSv/Fw4oGhHyfmURINq0fjv15yr
v0IKVgOO8UNOGyvDXYqAmlguHIj0TsPTPzcO8uwpvuu+sX1TVcA0+jAuZutZ5bD9
F90WkwmK6cqbrGow0E5imJ7lzwSo5QeFFZIm72CNSTPQ12oG3Jm2nlGPMUdBq7Zt
B0CkcpM2NtOSVbRDO8tw21jTmQpJ5VMKHuLgfaRXMBHoHNyoUqTNqs0xbW5U8MG6
4q5Chhf+PC7Pkkcqdhb5K8L6bdz0o3mrBZT0tejL5fGrzLogydf1h5YXbEiPihY4
gKYZ41ULx6zIYMq4KWw15QE9vXlaBNbMveSf3m/nBWyNvFPYE9E8UtuQYPFFmjzI
N9+leApu7ceQcx1Fg9Ue88P/qXQZG7f+EOcgNLZNcBrBz8EVys9xloKiL555Df7Z
L8C9O+CQS7qnBvRNq+Be3AhE8To7vbCtxPHjtsIel8DlrXBqu+ahYQ2zF62JxnRr
moCU+zHH/myBPfEdCXwmcbCtD7pvupDt/aYpbD6p1oaeeas9/2cm6Yj0nBWtOq0t
n2DqNM3jpwD9wq4IR8liqFrvrL6JdxjMTpWZVmF9Ml8/IU/m8EGMu5j4ph273nrT
RBeoNyqmvUw3ff03GrhIA00Fofb0KLJVmfTOrcTv6lfdcF+IjYrK6+0c4D8XL5Kh
AxPd1UzTl+sIvLf4wUYS8NUFQQ++EF6JaYNphN/6kkxTj/c1UGKdCfl0PsHtapmI
6z4S5RK6yQrzSxSPPUxCT5ry7d5rYSYa14nJ2CSAGltC+btksgAelLEGLTFW3rCe
S2sKms9CaC+TUuRCLRYrXTHj3oHvJBILMrZFmuWujEiI2cst6PXAnP9q0BQI+EO0
HQY0U/NJiitiRp9/wutdDOTkGRvL4XppEOYX10wW34wQewF9XwCPY8J6Wxb1TVki
Iju2CMZzkmbcB1cLHAGLVtBoIVdzCQJqQIN9W/BkjsHPz1ygo2XXATSZpwTZPfng
rUQtqiRZM9rOSX8/ocM1JpHRNB6MFa3Zs66NqMd/HBlYqVsSFr5JfnPsE4NV9LNh
h88lmWrd+vkF+TzbbwNA2snV7KaY0VuE6PsYTLrcfweBj1+FHG0LwywsxAKG6bFo
hhRof+A2E+HEcCo4RvRSXSTM0ve7OFG0fZeDw9t4+Rn09xNyuSKA2c6sbeSQ7Xg3
BZM/ovlU80+3L6vn3cfcn1qO6yqWWP1T5x4Jxj1wgAHdgdQ2AwsM8i5Dtf42EHpV
AWbD5xmm2QV91dBWLNXSnRKKRvvoyFPAcy6H1khbSaGI7zo56sIXJm9g2X4q2gcV
R/Mzeu164cyXO/DyJI04Vz9jhvYTQ8Zy78iKEB+qQVcMRAme81L8kBkxgh+TsqR7
RF0ZzzyfTPPXpg8DxPkt/JctQfA7lTLC6hSyKBEcPGfSuGNQonZ9RrCCwlR6qQ/E
YAaJZcFWGBAmA5EGFfwXuDAxzQ0WK8VVy6r76gdvGzhj2z3G3VnoKN1OwHcv4aWR
neKB+KTjJOPpydnErPgkOeqo1yAfhD6HtB2Hxm7tZV0X+VRqpL0JC0bb71SUFsh9
RniojH9YXieHcBrCANd501uYCRO95usJlMONG0FtRO8MZrE9votRWge0EHU3YqCJ
pwVvrw4oki0/Y3EYt+C+CAarf/MKQy//pYDDHXNrpz4ZuCgPIdR8cVlGHjd+iXbZ
d/siFWc7PFudPWvzRGVLWxkPmQCG2/xAdhNoiJDdTNmZ5Hkv+RPzaMU9untRP4tJ
RqFJSBBIEXB9jdEoKvgoPOq93egosTDCWQhaV9KEsIJ72rUoKL0gbUKNAKAca26S
1k3hyKGHp1h0pyJcpSVhLwnxa/8QQW7A3HNY8eMESChn+XoTl2MAat/nS/kugyph
WP9YkLxv6kfw7dVFN8LBlfaSfOWV/YtDv0zSWkd7moE+lkekMC94rxDYX0+AeGDY
eyfLiV+3GW4HKewEZMKvRwzgycDCf5aAFslqj1NUIV5GJvko9ld21INcX4AD7mgt
s8mLDRdMM1ZOLqHToBR5m829fSSxEkQhMoWRH0ogfwkUTtrR1wGccU856gu/bm5D
JRqKT9yKxS6UeURYi85gxDCvXoIxpjQVl6jnXTLmHd3tuOgo62hArDhK+3hvgd62
tElQcHqQZbalfZt/cGLmeD5DxhVJtZ0g8PRkNjdO6Uua2Ro4NogUV3hzrmmijXzx
WyoI+ixGxAEOn6/e9dif0cFScfNn371EevkDBT/ZXNzDjOYmuilRiV4AVkqUg2ck
Waq017YJ4tnZ3n1iBUNv1TZbUa8IQMPEkGPUgL2CPPzV1lUQBL+ZT8VUCtG7efkV
7HWf51knjW8leXij40bBfrQl5tWIQDhfwpNwkzHTQVmjOSClA2KTtZkdj9tS4LG2
Ix9Qoi5eWISocfFbUAV4DYFXAkQCxgPDQWdYfxdAfa2ghWho6SaTfzZ6xpg4qrpf
sE3hgMpDnqXe0S5aCx0X/Nte5dYiIHhJxtvdII+tX4NkBiWIeG1TF0C6uaGSyxf/
dVr8vTBB4lJm5atOVvgN6+r6KOyycwh4y0Y5nRc20g6BOucoXjdhskOQ7ObVcpTF
vBUutx/A9vyKoAzNKBYxgCAZxdPoRttFbtFxCwjZ/JJvLe82X75OJ6Ynxjlx7prH
DIbRHLwkmsELE6ltS1KrvKp6jOx2up2NcuBL/mYDLnCEBnMq++u+ja6WFwXKmR1Z
LCdsaSq+Rf5iYr5Z2mYmTQtxq3QjuDSmQ81EMAFxUXKMdJ40j6TUPkbYRWbYU4Ly
uRaZFvIr4kaGb4m0wWRfC8+PjNX8uVJjOoDa10I8Wfp8t9ZQ726T2L9w+nk01V7t
crN78hyrDgESxinTbnaqfKupm1TmeLQzIVcUnlRvyRTdBNttE2OQIjwpJphNY6st
IQJJA2/D2pMoVjXafdHi1va/2wTfw9h+LfSJo6hKamfqV2bqBkO38ZVK8imVs0T4
+34uu6kK8VeAxBdbsMDmGEs7utOwkIVm+Om0LPd9ihgrM4F9PxSRzJ4VKa+u4/VV
OYISp1rAa0RtNmU0tSfxBSYD1a+hsT6i0los+K3xp+Cs3+OoRmazzfUe2BBSG36+
pdqPQVoLHEf54uPTKIaDx0HWd13LlswfbSngyEMV88MHcfyxuANV7mWRI6gAz6Gh
OeDf8DfesYU0PeRfbMtpIpiOegXqXkfn7Y88BgRhFBQpinn5X6uOEu1ScPqtw7bv
OPxmHwiUFoyMUDC4hwILNsDOFJKq28ycGTqleomb73zTIj+X7GGzQZWDYGan248g
2hjaJKzzpyLsR+RC+F1R6Mf00OuLXM79j5BWRBcgs+0CrPoU2S8C5U6G0757sMG9
eSLeDFYO/FWgms0OvmzIZe0Yk4OVDrfE83pzriylkVQ4IdD5V4CJ455VwQwsGilq
e6iFtVY2iqz6jhQwHPrnP4RlpSdJxwps7MTM9HqyLWfXyPCT6gp1VjGkU6cVO8HK
0g9gYZFMzoYeCOV0YlXVNdUDhDnaNqulOEdLRpnqhBV96L2G9Y0Sv7MRf6RgH4np
JinIsAJ9O+rgn4WuNYnOu3TzMpfvYcgUT0ezdfc7HE1Nj5WuOAcZ9azqPtya6odo
EXvgJzjEK/k+YRoqmR7zU+/ZM9jIP0GB5GQEeyW7y8HSvA3DjU5FlMWThWYIfQTt
rTyrQ9SsHMCBCjZvewCVI+EzFn7AzrXD2B4MWwLaySGqHgUI14ti0LEheAREwHkN
V76K40htzV6rGkT+FVYfl2V6CFaOfcUSeYf4HiSewXLE20YVOXY/Vvnr4RjYfMfx
RVLbsUyaEko5WtRHbHnUMTST7LLLj0vu3B+bD6TkeUZ3xxeWRiR/0d0mkq+X9QnQ
FrKnYzbz3LLPeR0ygvxvPSZdO36Hu5zuSnDJCwh+BM2JyQPFZ8xcnijQ5r1IRrZb
XTyJRJ26/mNik9M5jMi/jYrOTjye2b5zOUTu3WgNoNxWrVdFITJZK9qu8KQiq500
3xuLUiKVGR35YhdakPuvhKWWflbwmI092bJdOcqohAiQQ5m9iLUctEH8lAucT4CG
h3WWoOKtLW8R+MdGiGfUVwEyrHNYN7Vyh2aVaelwKeRwDYD+ofqrGq1nSDIB67wJ
55dEkN7laaUfTXm3pWRcrYybnHZcbcDRLm6KNMfI70q1cN4FTffrlYI7EECmI2ly
KalYm5L8x+cOgZav6cH6uGj5RkL+J/PDWM34VOf3h0eL18njVStQcF/OlWbZlBsL
VXbitZ75sy7LAms9z7PkDTUIdPb763Iv/yIwNwmuyPN5DP7ehfNrZ1d23xQ79x8v
vrPCboeijfryYjmNKJSjwIheQ0Ya3zAHOYzAoENybmF1figb9K0+h6/ODsK3d2ZC
CcpH2IAizLyX5QZbtKh4PAPJ497I8UXA8WONm7uwf1dqnsD1h0TLTlUZYeY7iY68
V1uEjgy/zNHXC+zeuioENsgtvkJKo9/iKPGXu2wx0E3EcpIbkuPTtzy4mNVBsLjz
095LB51bkFiAlmaNC5JEn7fqK50XhdTxCwXlL4K01hjIvIAzpdeBgrfS99SZXtyJ
u9wHVfw0j2kn5bNX6et274c+r8HwvEjCcn1Jqle9DQ8PFGfnsGDlAk0K1nnM5srG
U/sSjnFubvKory/EnwCr8kKHKwZRh31PkEAQjSqS57EGEz+WbO8ydFZKwgOeJUkK
J8EZbgqTKqBWSSqKDnWfESZFqE0/sZHDu54upT//Z3+KG/AcWvgC66bHocZW4yOk
yt9aK+k15IBzWW6QF5ADS1VH3Lxpl+XPhZZ41dWGb3E5nse8ixY8/IsLY0y/zKVn
v1sKdPKursvpSr707s6PtPs8IENzgdeqTabkvgF8pnW/cC3bHdvt3iAjKXDRQOjp
WgdY0n59ldkJ2mpv4elYE/QLJmdnaYtRNxXnOhJrIcK+ufpP4wygT4bT4vbSPFeD
iB9dJec6ZuWWCcNVIkLFoI1Wzr8vkuIXEkB2qzbV+qPPZZcPyPdPnBveTB/9D7R0
UtL6J7bySFJel8oHQAlhcAWqHg0S7a/XpkQ3lG3Lq40gi/+6YC9jUFlm2PmIeRDy
+DOaPqZ7VUvwLTmya6PAfavGnKcW0yv/FyI5rYLfHN3A4YRqG6loyuJ7pFcmI0LM
7bHOgtw9Nihn4B1Q3z26hn7Q+YBdEO/5iFzE8wKQjHujyVchnqVRuilXbiX71blr
A6l2YOSZctmCYY3LdL9WYL+NUARFTtv+EzFubT2ege7fCjjFrlZjzjeVMCt7g4PS
3Br1T74DEywMtKbs6iE0ff6uhga8+Tjp2C7wP8ozmCI9rWwsTAIIwJr3diPTi96A
Uz+lGDO+kPrhwPVZifKv0JVBMoMtuiF5JEDZ+1kvZ/PB3rfVA7cyvVLJD1ALtxzz
YOoDVMjr6YChUeaFa4y0zvPK5k4F7I0I8wbNTmjmw5x8BJeF0LPYxOxH3e9RHI5U
CK4Mdoerd1VvJijR0F/1JJWvtCKvlyDE7bpNniUW33/r9fUmQyNuUNqrbIDIiMIw
aXe7Pvm/HTzJYutK56oRjw8i+vaSh64yZjkeNTuGQ3mKvOD1G/dfEVCT+5rV4apM
Xy+iHfeT93SN3+j75b0p3ezPwCJwTA4bFZe4zH9+e1aso6vD6lY1lEAXc9jb5Mpx
tEqNAV5C92KUNjwwyZjZBmANPkvktZl9Oeyk997RQNGeNfXSotWm2fpT+aA5O7Ki
+6Xs2M+/CqNNpOobHtq+t6AEJxEJWwCTB5c7ZP8HmqtnW/07awqO/J4Q9qKNadHv
EW/K1KwWM6Rcaeul9FRRxBGHVNCXSuO+LZwyQQRUZRSxB/oYkw7BadH5cPp9Ewqr
u0Jg6fExXOYXRswDcZJvONd0Bxmi1aS2ir3CcQIUF1BGbKPf7vpbx6JWsTpX4LBw
+vdKi4P9y6rk0glzLltxnH2+dtbW+jr0dhcskzq9eQ1wR66ebPT8jayL96+FChak
6E9GHc2yHH5qg7FbmfgFPhFVSx9Y3DwdLnh2tqW5S91I+iz1gMzJrPTmV8NCeF84
UD8Rarf36RH/QWOP/9ac90bkkefqyjgGEKA1ensmBy7OaQoQPuLRUNpceGPfEv4j
msfPJnopWqIvCFaBz63g3IehrTVQbfJnlKBsBpcohjGrHHIH8odMVxJF9uO2n5ck
M97yQ6ZZVGOjfXUPqn3AVBKZ/RD/v7CQMNOXyNd/ph5YAdqFlsuibHcSuxtGVoYS
d2qFctD8xAAQbdq7y4ueFqZ1q/WIVf9JWU1yLY1hpquvGg5SZ2y0ldnvJnd0PfML
oTA/m2p3oSfUVe484OozwOnkas/npVT+IjVgCam4SVRR1cFqXfLySIX2ZVWiQ873
xjqgJQ2JvaePHp+0ctGfoUV+y139hoXQ30QTgSyYi9/C/9c42ainPq+wDhjqXOaQ
mT4LOhuoLMz7fLihqTYpI05f/ApY/67fpycrSkqhJKQ15oyS8vfd1A555CP1Fnr4
WbmGOg260xrTKS7O/8EbM7daDaDFuFG32fz1vC5EsWyF5U64n73aNrbzMEUFUEYi
dhJn2I0UvIyXRH1wh01J56Qp5xs+MVE0B395zINTqRKENTc5tASm7ketMVJ5NnNe
zO9XpYLgOEnvYp/n3LeAJS+WCDdHKqW3qpmlT2OGZAd1DKiuIR6OMiosGcoD+LHQ
SjxODA+jU6Iana7eF5P1W/FKNKwJBNmHf20XTKJmBwWpStRcacFkZAljnN8eQw9w
L6KUkQhjpk865tygHg2s0NYHMGFE8kTmYzrnW7gealLef4uY6GNsQSyAscYKXtdy
+qOntexf9w6XSre9seeQYBU8FbLqqdrVce3q8QTq2HnkGnF9ak+Yh33YHJL7DVzB
O1MduV3uy3RnLR2O6xuAI0TAL+PURKeOyqVBt3bMohljqjF2nl/JZ1YTgC9lFI3z
YImzwNRXqszMsCFJmZdCQ8Ly1YcOdtUul/1iD681kSEn/A96ANpb5VNvVVo0bb+f
aUgB0IVcpbXlA4peqz93nbc5vsJwhpFuJtIWt3v0Q44anVfuzvE/EouI6NnM8cjz
TbLlztpsvnNoltIGCPzlDBUiBAFZwXjZToVc4rfe3ZRbshTbK6X4narQG8bULkk7
Cx2QDOqCiNoJnV004X+gC1ftAHLy0ezf2I5+rFgrX34oiddvHR4WLeX2TPDgb06D
MMD0DkfSKlmxonTP/JCF5OSRjHhntMJ+ECBoLuQxpnHU8iXNzXX3mbGhNpfzWqCY
qv5dgh76d3KefbyfbUpN72Z70h8vyvBqwbuPtON+CSP/CxlgfXpoKZxwXN41JjiQ
XTyWIK/xOD869fdtmsnllfr8j/XtO4Gd13EggZPaRPfpN+emKhwgGUmCyx3Ilkm6
uGG7iSQzoGvg5+6VA8siIcAL0cqLbo+vxDCwHvKnBF84JiOWcVQ5kRjt4RTImrBQ
HDwmjIOsH87sbNkngg/57gJJ8hSdbIV+3Tii+f5BmIE0Zc6F+zDPGExeRVLhQesS
lOlP5/cIhcK6RMaE7o2/+n5/V56QCb+4L4nDsd1Ay7BcBvwIB1NwaQUV+0iFJI/E
VxO2PfFobngSvaIkkf0ni0ko00/0S6bqRuv1W48X/joUMWDWO7tDnDSMy9hDlXK/
NttJOjhYhK3ZoXzT4QOWcmh6FuTL8fprbbZHhGRE3Oc3wYaOcXfpWzVflNf1Fe6z
0RJw7Wi5+in5Ow+fzT6yG8wQ4jIAanWKn11oxVjZ/E2Jijg+Eab7SDqt2b+H2GDU
d0Lgd7kx3oGT378z/nG+Gj9bcLBKSbKtkR5X65tqQ2h0OMF7PpZM/A2kgq4CAuhH
GUiJ/HQb3C2594kRT7rgmCN6JNsu2H11uan23y2OkmFjw349lPc3vpwOI02CUoAi
BMgq+sTt3guqGuWsvseK0tGeLSkxOwQpnJml9h2ZIA+naUwBFC9vhJyUIRxcUJZz
2dSpFZRyU5BNsBofzYvdJU/dwODutrpiCuNE8jU+hhs+Xbz34ZHDDJPuuUqh8Ux5
yp+x4aVhhW3MHMWW9pkIgpSlIY12QyuvwudF97YlRBmAdFZTeWeupX99NJGr04Xi
Hx5ZsIfOj9y2GggEgjRpTTsQVG4wH697w4ojkGaxot8/qKJ+41Ro81bw5NiNUzUk
whGF3NrMdCv7sDqzEQM9pkWO7VkRHkdSWsIX4bozBKWYe4fKF8Er/S+Ae2ki+gqR
unAUfHGK/r4yV5fjOM7IeRHEH5+S6sDwECNi1A2nYDkyDtmanLN3JOwhGhvTsrWg
5WayKQghidmx3VDUeCVIzUcXX51EA59SV/Ju/Pv9LHqbNwTdfkg5GhPMVoRqD73B
8sZhVGeokwb/XGtDa5AAYztL38Q9m+574q2GoisZD4Q78mJYt0StMeDqPU7Fztzv
ndkITRCj6PHnsz02I8z8WzoFkZYqVUNmB2Wq8KQdna9V0334XnJek/Z/U89ldkql
o1xl4rB9qpporYaOIALm4CFc1Wdu+dUeIOEfjDQeWZKK+VHe7cH8JWp4NGT3JbJx
SlhInfQboMlRKZRYxQTYKYM71nKb3Ta52j7NJR+9bmWBOOtW+PctTdnzE/Ob2FXN
pkP4sh6rbN2iz2PY0D43R6xgFf1yFlCHgZciPjVErvr58iJdR4Opms7uk1Z1CvCh
lM+6Evqt9dj1RqsF3XMHnF/PVVOt9cz49h7E00wvywFyC2kMn/RyrB9+TqTdmdt2
suDk9531SdJI0mAWypXwgiX2zW8o5eKZ1XimsRjHK6+gKe1LzR6uNEIGtzYa9Nkx
NjtrPVlk/kx4ypJB7Hi9Kwv1SrnbJUMDIRhAvQxbA5b2viBsAuzfoahTY7vrQPwR
Kt8dMCJ12iQXjzWNPrE5SVL+C/S4dW9LOe9XNkynDt5RtmjeVrWigNFCnpvMhENE
NrLeo8g8Q7OSCVQWm19o8t8dZ7TFhXQXH3ClUvqRc6hWNRgp1JLfrdiIGwMjRDNF
L2aGslOtIKjG/43PoQC4yftdZ3KJW28tjIm87khttjFBAGxyMUS3cw2/AGQ4dwTl
YegmVp2U2RKGoSz5eLId71m5T1aj95ZNV8GUEyS2LukoQ8aHQUa12aB6C+oDqR85
o8wRbVH7hBBde8YBDU2vcLBaFgNDsRvwBfnYtYf652B/9Yu9NMiPm/Eoi23XPmq5
v9/tgsfj+pkysbte73tHeF0y3cwf5sqDTVJmlaXYi3FQN3MYjNINQE4+GnVjZPFJ
t2zb1CUVU9T85MMmmA6yCJa8MPQJ11Ik34zZoTuj/vzmZpzyLu4dj7OBPF7VHrRw
zMBiU1H0njOkNk1sonVqJvbFFSv7o64XcKImqOqvCNu9OPV13k0qdnTtauL+aiU5
iT1dLwKQ8/HvSU3ega7CgP4dWIvlXSBetKcEqySqme01oU5T8C0p76cBzswa5KVh
nfAbLxNk8G3xbcRoL/hfvM6O3qBbetf9RGalmNHltY5dCwxEGIRcunKOKaKT3Bk2
zTUoDmKlXux8j/Y4qA8v/jS94LaK/z2ZFqac7o6VkUF0lTg7kBISva9/r282G7oX
Cz8QWbewclvEthMtqsBk3tqG8xXqx5PwX+8WYVUVQb98CtfDAdhh5ZjI595Oe2IN
THrhg7ja6gTQ4Alu9Dfkwua4JhfTn3DfOWWvynHM24cc42IBqdVoHHOpATxCUK/K
5W998FPgLZU8PSKMxfv9pjhTb//tzWkncfEOu3wGAF9L7pUx9LXR+yZvQfN2syKB
ps9ldg7RL7Y0c5VwPuhpHCd0zoLJecC8y6RiKmiQvUjjlHlLYcvNzfLrJR5GMqUs
MW3MFgFM+yaXoUQjDUAdfOO3YJy4st1AsRCi3MmSmHMBSyASyLg80EW1YkRwOvtd
r88e5e+NnroKONyD7OACWgAoIipwx/eKDJsKN/pRmt11g7PDfaHATSiTYmWmjp8E
dTSYDOPc+bc3mHTQbxd9APilcA0xyGqjeVmKCMQOTXr45IYoRVVQRabHlBX/bn+u
ja3Fzu+tE0RxQv2j/t3gE0U8NlbLEpNCkb+VnTaav2Pde/Qe49fKUHz0OhOsrYy7
BVmDFki3qMxleBvL6ewitWKTAHDAkTif2ldCf4jMWZIWcIa7kTK2dZ6HQDFz9zM6
C8v7QRTb45DuEq6lsuC7yIM+OS6O0GuUjNBvBiKL1WhNH9HT7NbZ1Fj+P33P/JoG
Y6F77VIl3foUyNXzUcvWd/ylLCclI5e25GdfKPYaraIuPEiAV/E8u6f8ayFoeX9J
150h0WwehZnvFKa2vlw5VFyWhQ0/2YI07pLwgAt2UvrI/y0OhkvQxtSDqpC7HC0F
p/PWG94D24A9MZfz2AVQ2UrzD0K7ensp5MGEf+yQmjJkBMiMbto8l098N9rbTE2Z
Qg5KIHYnob/8SmH0mf9eTeQkNdeaj5NpOgrRzMp8SP8xLa/iX7lXlhRg7rvxObxe
pPlw687PGUbORSStDBPryv9YMHQnpz6f1wuF0gbg+0uN+iZnO9BSSrUEkE1T/2EG
GChktgcBY4XuB0nDRDvfvdauaEHJFzY4Id8qgRlXuH3lLUZJxCB0GQipsEKYW/1C
7B//nTa3JyMf2EenHs3oJ3i5+iwvQZnmcdNqyFWoqaJEAUFAUsDOMPHB9kP9sZTn
5mhr8BRLyIV2cLkvL28b6DixHqU3oPVwQoyST10FGezRSTlNvvOcc5Ftwqvhk/2I
AmBBG46pShVkPqFMisZ2ilekhiDPDAbKjVBkzbSnHoGjmhYJz8AwQ7i4fS0AzC8v
vdRFskrwoXYGFRbrPMHkHUSygvSrnhkL0JJmiY+A170L1APD2o1KSapzPjBlP+Me
NNJnfLESUhKNmfb9fha2EwR1agQHgTBsFxsZORorBlYwKB+DplMdn9GN8Lf0Nbpz
H/bYfgVvTNh7ldTA65/YDQMlDFeCYGIvx1FaRy+1OPla3W6fP5NFEMSOIDrQemG/
gw7sINR7Ncg/brMAB3VhLwezCDgLtzj7p/jBeqsjHaC+unGyC9sjQcYgNAE/DkxF
VM2lpJFxcPCDaDdREPIMGDKAy9S/izE53tZJ4L3L4rbTkNFFXMiI5H3e845YTSt9
UqdbyIBmRQxe+ITg5raXuemPKtrbyBfzFjit1DMSktSQ+I/tvc1PxDPyD/W2CB6V
z5U2/S0hI1mJzE6gogqEzbsXLX66DpYHaVyOZOl/5QsZwGFw+SpbcRwkaLEmFWlr
jbfaHKPk5aOINLoqhGgiyvMphyLpYYBdoLaE/d3o3IhF1lIORFyPvZEs6olBa8OS
quUiLXIw2ViPAAAN6UpF/OjvDHu0oba+4JMgZN6jW/Hc7u1BVctM4mPK497aTjAh
LGqn13xLwowIAYNGxwKcoJrNN5Ss5FIYb/mGKRPAeOJ+M9ELipIrHiHIiukcN7VR
k0KJq5EDHVHZloG1wgN019n+/LPSIzIaqQc4Tzoa4q610/DxXDkZfOVST2nootK2
MeCxJyDnSj7HYiUusQ238iK9ciDnF3eQpsHSNhC1cLvNDNLHcs7wwBJ4CTh19po8
iMJ4YN/a5RI9oHFkpxlDtA6/oWOd11XrqXjWcgB3/z/8GvlwYOjwnIfrhcW3xROa
IBhQ9GRLRQaGH8Lf8zsjKouV4CvNDrBbdESlktWTYKbxDr8oGEY2SP1vgOG+8SXy
aXWSdUQKF7dBzND8nZ4X9uh/B8UmIPTGRlQCxHiQILeiClUZzSDxRgGOMQhqOZHQ
ovoKDyOu2bO6YnEPGdDrtk/ToIgUsY/xMD9qhN48kRzw0JjEk6ob0RO8w+Xig2Fv
vRDtQTdZFkapXVR+L/LpsGWZWu9nXpu96LPks3pD1gxRffQY3yNnnL19i6ChuZXL
mls0aCm0XBPQHIS13xjBvl7b9P/Cq3JTRbscjJcfHMGWhRfxgMuKPCJN6svHoNJt
Y1BbE+1LxJKav/+r7Fvna1Jg7jXngpYBTKnekZQAXBYzBU/737rRRQjFY9I+N3mg
xE+muYvsEYkcqTihDGVKtYjxF/QVQTOBGHaxZTGSL3SY6rbzkR5vWy5qS2596JOl
GK6oGNYGYoRDcj09hH2tLutZAk5l6Q0gAKj90/WCDCicmaCl2DcDJx50OwAf4Fwt
toCCkI+tJwzxxJqQNBniTCf6p6T1OqlgBi9GxHGIQZ+rTA79vGcUa8isbMFeoR6M
KWEL2H2Gh0uF3KyLreuOdyzjqqYDG4jCTUSE9CikrT7012JG/GYbL0DXuN3Wl7KY
wr9alIKezi8Yx1Vp+VqwEsTvf4lnOw3SQVCL3aRMdlsgXAY9tERL+2r2EAcDfbd6
lt4t3S6AE+BJaqmmPq+mUmzgzVp2wu+dTceXqPwB/ZHzDiSu0XtBbtLJuRSjeG0q
absCRuLqqevFftEEunFy+MYZ9L6ZKZXRjvi4ct32mzCCE7SfYMuYqkbL1qizhwgA
bUTx7sp3BftLW6ylt0zhHdsxbz7R6hv8CC2MUqZuhc5A6qPIB3m1jyfiH9ZJ2xlZ
0HYL/ZRj8PVWbhVfSxggihw36dr/grd3SghcTbX1UvtjrfzotP2wY7yCOf0VOna3
B/HXtDE3LmUWMSWjHRjCQHfb08MxZsXooeQhT+j7gn+ncIrGyb8KAEPmUoJDJfD3
qvUPC+lqFy9Yn2FUeDhwqAPjH4JPhp6MEN7Yu2MnpUfzQR0V4GSwAcwn2YbF+tQ/
gIjkTb2FZ0p5bQR8srPki0vVDQyiMrQkr9O2377OgnUcAfNXBoCmU1v8epw2gvmo
bB93D7N9v/M05Y4n42kWKwjniwWFikufdHs2MRC8b2o612rmkHjwy5yrs9tUMY+e
xZG5SEZFVWoF8Pgk5Gi5nh+Zz1qqL4mphysUV6VsfyTJfSi6MGKc14WyaihyYERS
ADgrnGhPkBdKpG+WwfUJ88sh18KmJUCJW2nvYO3GTzR0YiqgO2BBkf+hqkogB3v1
RzTJZ6+fXwGYXh8zjE61pizrTHqxGBYg1kh5IDayEeSqCdS1f36VyvTJxksl0yii
XTYBZrK3lY4/yQx5bQvftfRYSBvMT2nnm/VRfSt/yCb+RkHu08F1WHPhBpFPCSQy
rQc+FlFj3HOY973PiQ7A0PJ1R55R/I1Yr08bS/tQr9W8rfsqsPnxy+hlMhBRihxh
yc9IZ7TeZMo0Z/Nf7LLWYP1H2mylfn1bkmkQYd2mA91rHvkES3lc2y9qg9PgGyRl
YEbP+IApzJ122e09ZKiIeeAI7odhmews+1R0+MFf8Lo/bW1xo6vEwWkBs2IEKtN8
If0ud1I1DWt0lS0NLAuBuzdx2DHOi6wIr84b9t9xBhEhmB9isbL5QJeyDTKO4ObG
LchRSDVWWbiKZ0IcA19NcHjT683/XJpdkHoKJ+m+uwz6T4VrD/G6O+NZpChseEiJ
LTr2wYHM0sCFQoiJbOOPEijpq4jT1BK1LGGRZkHq9rCBS5QRN8bU95m8Ax9Oqyyf
DRQMv+mpzuIDUF7qaUc0EQbTxuCeUVXYNIj08ELvPnV2kkQTH0s5BT1TDH8ne6eK
YBI7g/jGMuG2IAYlOeXVDy1ZdhogxBePUjC1hRJ3Gh2SPodnYBcEd4ewOLgMTVgK
WLZdrgGMd6fOVSPQ0C+SaiLyeMk+0H0WTSXnIS+j0DFag//KhQbRFmD2TPXDRRQQ
kfhcbJhXtTb6IFIO0lOrUZMdHgmm7ebWZJ3pjRIDwVpS3Zt06acM/d2VAXhY8Plr
RnvUf7V6a96On7AxXtK75xpCxEvfsFCQ0et1WijBIc6pVPfPssAJlCl3vFzSiviQ
X53Bi2EmWqrvrpMRt1/edacnQLf3h1+Hb6TuJv/aXOqpgduO1nPyMXMkujoliD5u
JTP3HGIDQa/h0ooJVxzU++AhoNsWHaFjpFe1Rw7tt9R1FJNVttcYYSiyE0O6gPld
8BaPJNXnEHLEK1ciLtFUXX4M0ns6n611Dp/qA946FJ5hovEeh0Azr//VpUswlaSs
WLnbMgmjoFjQmkmY3gXvqVe8u7AQmzrtxp/Dnb/FkdZj3Nzt8GQU/t6MrrMvz+lH
9yGNJty6Zxpg1mTNvwqHNyteqge9nBpUrmQUE0ZuYBV1gpSGKiD3nS/2+iFs/N4E
3CyXbnew6xwrJNRVm2Lawb4sBHBVaKfkckzD8TUNZybl+vF7ZCJmIqGwt/j3tQvs
iZ7I9WsnlVKjYSygUVUhCe4roA2oWLYqB7QoA0ZH5Wlk8KyN27+JWAnhX1qmWAWz
6BKEMu6q8Cz6l7bJAQY1uqjGDZEySpmD7OH1er5EewdgZuNBkDtB/aUfA+C5T1T5
PuUsyVwEDhe07malvq4k4oBMJE5xnpClA1thp4RCxiqU1WYHslyOWncwW7YYBNTV
9/C+qpQZH7CbZcNcpNJEXoh2pz9MtAYjZzLSMv29XWoURQv6JzbxrFO0fiFImxRE
+9xMn7B+jXSyxI7qeXETEn4BQTH4slkbZl9huzht5yYaneP7gki4+I8REX72w3qa
2EkzdCEofC7R3Oj9whAnwoi4WEISeab9EUs6VayPtocfxdHF4OS2ORnRGAkd2xG3
xxNPcgNykoOEEUxwSrJCnGXXG4E6rhGmKbkZdJ6ONlsDt++sznwiab28avZDA/3F
WfAShLXkMBlixiMvTJFw+BUNvGrSX+vQMTz8rm77vjaXMcrIjoabjG4MLfWdwdhu
Bqf1mFimAJi4iQdx250Q4zC1bMZpXrPf4XoE3OYPh+wkMgki1FfGAUGO1ahaDUpr
Iyk62WVNg6j1nBTwD60NR7fGXIHDNrpeQGqNz4iPRo0JH5I4mfsVOaBHhRPdZGgj
1LqOw2+wwiC3rRVMfJP4RJUm8x3NZOu65x8Xbvqxc60eTzta4paZdr5kV5TkEDNM
CdwdT0CeDckXFF4G1LDmyEkE6vtBSXDwNOcnggte61jucLsAGoznwOX83bUIG53M
hcct8bfjlEyykfDLclTkhg+nvz5jGlilYSu6Tj3Pm/qobzEmSlR33ObtFlwweEhU
JKWNFEhXA/nZsoQexzRnWPlpHPdATMlzhViW4yCjGuk5irtRd4+m3SuQAebTsF97
xOYjn82yUWBhABUBS9fecWIg69WujK7Mmpeb4hfrcN/V7TNJJxeNmmA6mNEdaybH
OeK/pI0qtlYA/5W/NcegoVKN2NWHHAinI7bkzFyckncN6l362Ty5Pn8E5R7toPNK
KWlcgfNVkDhkjwG+AV4nSt0KrbvrlykoDhNPr77UOQJT2G7ZX+5rZtTrtUEY05wn
7zJptxCOiO8yZ8NNkPFR0ICHAt6iV/E/oeUo+M0mqCE6rcDlChhTRcp2fUTA9rzN
nunG8gU0PZ1b06n4zFuBDbwWMNiuQcI9hgQGWkc5tPYHBG2n0xE3MJn7QeMvdhMa
hEw1RidZaqRr/oTS8N/jsHhXU4BgNTbXkqi+9rJmeayv/LkmCdL6cCUkYMtH1BqY
NpY5U4TVabD/A7FV1pdkb26H/QZ6QeJLMDttgY5N6a+TueRjJh2JipULglHBCbxf
OWrlUQ1tTh0dWiWxYhDbijUkb6vJ5W/an7wZBXwmoNZhpjfEWEHi/4GqaCV9es9+
9pN4LWpEWBL+QmJ+J2/rkiU6dtySrirGnlAkxcCnviG/NLcu7ENF/eqGeeLDvMBw
VdnTuewzHuiF0OOC6abN96BuSM2i++AEt2cWkpcuzYbL/PY2+qe3jIaIipyZMBQf
lh5xobw4ItafaarLavU8wFVlEzJ4MkKLtDiKfKK9IsNxJ7ScZ3NZ23WUp5DSC638
0AwhWS1gD+AtFIKTzVOjMB14OaRgPL8sy8FZFfZYiI4TE7ft8W8eebGg169SHgcr
35MMpdR3IiuXVnbsx7hvTFyCtzby9hb4sumrIdbzV9Pkj8c15jjz6L+UhrLPysVe
ObSJi+ghEUHTMuo4pR3o8ayNqP23cjeU+ey1tLQrMA1vIgn4+CC0IZH7jzdh1YMk
vBe7jlQUx8xPgOlEhbkSEbBR+1SndYL84Cgdk5NccMG5BzMxQpSl9LCfGVG5zrfp
8Fm/XTX+h0Dv3XD1ABcx5UI4zMyH9adbi2LRCt5ratC3IqsZeINYI5BDJVklbfyp
4kJN9bcLWWodzI3KaPio6TEcSjduRx4TH2ZzZ1hwhZonGvQh9VUUcKdbuk8ZJTDv
`protect end_protected