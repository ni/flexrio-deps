<<<<<<< HEAD:flexrio_deps/MacallanIFifo.vhd
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11328 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3b6eMZvf+eQ8z14wALfTJHs
q3E8aWgVMNpEXpVH8GIRPzdig6RQTDao0E7IF050lcnDGBUuo8smSU3lxCVMCwZI
D73pqLhh3mNnD2tU8PLH6Hxw73vdtpUi9EfNfbSppKm/b1TIE1ZEKeCsC+1f8ii8
O+BDX+JaR2Um3PrP2AL1EgUIxQ8WX4+kuZDtp5uJdYwYy7VJFYjH4x84Mebx89wB
hNIEbVZO8f3CETn78Wc/r1Qnqh/1eH7C93gMFkHIPyYbhlXSCGOH8gz/DMeD52PO
VOMq8qYu6d+UO23xAzxD3kw7MV5ip3XIX6YQMdsi8MSeYJqtdhW9CovkLAVAlE2f
mnPCxZHKjQ5zFU/TA6ucs2gnxGm6MDwy85fu1Pi/vADchelvq2TIZgXfDKvos6KF
pppsM0n6koQ1bB1btgX6PB2T/myRs9sMIQkG0GQ+TjQJ1Fr/DQ7PNjqlFgofgWyp
L0ZT3cKKApjdPlvZ/LaAjJMZG4wzhsIqx4s/dtw7BiyYWSsXnASpiEE5iMBSrZ45
fI7Yk6XYkG4VGbrFWrPQ2LCwO1nwTZGGuycTarHaX5/FghFDerFW0qVbZmpMpPid
gLeyZjObsOxkoig/bJTqqkWz5McC5pFHhDiS7kToeMef76CMge1H6JskVDeOGUNm
dJDffDeJyqcnTTc0Ix++6iLiM4VffZgem/i8EPqMcB2Z3zHMC6eTRtDdQEeoWKMa
gaHImrAPMkF5hWWqepdOM1wVKGIkWIA6j3Rq15wpVqHz8MAAtk4ffdMSVaHmn5wf
LahXeuLZXnaiPqkeV/NHtYg466aIfXFJvzpJlKNzbit24Wpp7H7aBk3TkwDqO0eg
xS3Ywec+GfXUsetnx6bTI5A+RaabgewGNo3H514Mr7VlIr0vusyMAHfBDe4hY30E
kMR6CnQlF4vXL7Hs3p5gcwzigd97u+GI00924utek3iaRO9tY5POXgkzmD/FH1ot
NZQjnf7xfyzfbP8UI8necNI9rXYbt+2Uu8Kla1OZZG+JE+uJSotbnIUfmZaxXTWY
xvmXhnQmDinzwGc2kYX2VuBShIQXwJNqVaue1S3QCBqiMgxNkmfnm656ibNl3+aH
MMM/M7ejzR7sajhv6TRtQ/3KasPmU5Ez30A0LW2E3wCTACPEfG+zPLgeLRh3FV72
PTy825wPK2hNgS5vOA7ehyGl/1oxaUkK54RQtjJYwQ8FjR7C/8jxU/wIxw2VlPON
8ZkcTDM1ddQpvynj4xn28d/1v8gH28FgnoDSjl34K0RGZcyAQCVs0BNj9CDLg/p2
OMrnZ3mKiHM6nq5kaZ2kvPggE64ryUkHNyQ3LkXQBy70O8zM753VK3K3rdmsXSIO
RiUbyS7PmyBJwn3Ko/rGC7nuAr85ySZ26sb7JP2gO957Z/YeBmvVlw+/pkY+RLRT
P/R5DPosq40eeJSEQO3n8FhdOGTuS8w0i563QK66y+2U9uTAMRXDBU/jpZT5U20O
LkHH8Mw+mdnwhAp+6G4fEXOqEGJecVWg1RygY4L+B5nXOpmbpNlObpIJkx5BMVKr
jAhk6IFVPmFSSlyI1kVOHwypSwLTNfBGvUBtcKwZ6c97ZOVukL5z14kIhlKJCDws
9GoMcaKUWs776cDxu0LfvcO9lylXGBHbtOcRLFLVGJaX+QC4fTcgFX2XJL3Sy9zz
dBG1LSitxiUDPw1ncw2NP/F9Jv0zegL3vKdSCQhBkDaGI0IB9k8zhRsmP4QaDGrQ
3hMhv8aVnpP57YVVuRsnumkxuCeXa6XNC/JzGFZ8vqvG2RMIFMbg4dQxvMcnGtEL
3crF4/25iTH5M0v/aeO9XAnXUMvsg3q3/ieQ8FaIAQCLBTi8A2NKJxgJIANC070n
ZpyAXMxRqHC/Vomz5aeYcuMqXZisC93+Cf7h3k5c+PcBvoCLs8QVWl46EH6eF8rL
ztAhdo0X7xM1qcfL9JzmpJH270pmxTY+eXRfmsrBcmxzZseQNPZkVJVAXST77I3w
0P09S812cOxRjPEpo2L9KmzQzM2NRifJ7ka4qNBk2GzMXJiPukQDdhU83dPRLUzp
ukGBnrJnyhSRtJglalfoMGIlaN/mlYkRfn5+E7Ip0P1l5Q0sXak9bE5EQxfko7sw
T3LlZjo4rOANrxGJAh6IF2oR0XNFlLhQIYIlOVMkZjUX5xITyc1otFJpd4IB5CJ4
MfMNOvxfCLivD+SlZGBvnkDfP07CV7NUC7dbFTjhcfn/ORRrCsG3EjhmmatZgkSo
t7Mtk+/tM8fvV/nLwSloo+OcoBnfcgCkBlrneWSboaG+SOQ+AtSPEvwyeqQZc/3y
8thFFsEzKwlSVCQqwGqpMkL2Xhd3xVaLBuZzOudz5Jp7ae70gJavxeYEhVPdShWw
lfG1CaLnHDYRBs+HFkJKn/mXjGjeopsYvE9fGuf0yIWoM0NrEzBXUlgXxfGWWgnu
399Un1kjjdmbBuc99uHKF61r6/P369G1kKEGU+mGyjXWKryrykdHsayH69fO9g4u
tthMnfiQQl4NFrRtcZdTvNwbrHPBNHoMJeMFyV3CfmU1ModMzhYdND0pCBLBEfNt
uC8fhIF4efLch+WeOz88MEES73x++gzqZlE0s2475w2aAIZIwiVRFitdZyuZAWzo
OUz5cuOLk70o8CDBuQY7a/BmE3ufxy7lcQyjdby84RQO66rFvU7aR37wedDM8PC2
yDwQDyxVtoNfBhAg4JPQqu2vrsVFW6Zmju9AHBrSr+PxVNPwn+pQ8JzLU6ekgZcl
sho/MOJ93WvzKc4gOJVLw77ZDyRihXlIdiPthdUr6mCHjKeOZ4XfFIoJ8citekMI
IZwlczzRaA/OqrVvm6HlJzhIiUyREWPg+2+EfsWTbxAjvUg9b5QLcHQIC2lnl9/I
nge6uIPC6N/n47KbPV7rJcD00ZZgxjtKKswNAKWpy4DpQxXpiZnwOeIgeChoowaN
P7r9Xar7DWuP2ACikkPbyBMBQHed1glpJv8dNN9d6YkbAV3MPztbhecYLjw3yfci
EKgsD11rdwVlL07LXvwyHBZlqFBZw4ld6OwObulVHujwZhj4e051CQkBo75vPOAV
e1TUDe/1Js3NxPXNVRHY2nNkdYNqx6KUXa5ExvYQVq3SD6DKNwcMDFxNgNTjMJyn
wMdqTaoQV8jeNvYUMg8cxud8MXZyk6qLcYOBFosu9R0OC/qzrKPRkOkw4WdXzEUx
NRMMlnroC9/R78w30pe0jd1fQOcE9fSFgEleQajVHPwMZgrcHdWfALJhFUuwCtD8
6RzVpaOCCrGt0BYg++PaZ2eSvrLnqYDV17aKQS/+lQF1fp78al3ME7367OWs/1PG
qSn5MOwclcU7Pr67NKh3Y+cLiPpeVJ3/fvC3rvb5IddCalayenVZhMmBnZvQ73su
EjVYeIdWi0KnJhCixDi5RFqF6K7iNrI3Kr5vAHHu9fikw+fM7xmzwArQj3k6TAQZ
tWQbY7QUuwMrsK4nkSvfk82u/LHjch4O5UOWN2b9XFp2L3HS6zcBJKCT6lJhAt0g
1qj12Lo1S1AcIihOTFm04BFkfkIpUHjgaGTL9CT9/rZ/EUvVWhvPIjgf48kOQGxL
isPo574P5yz7fMJB1nCip2dGKJkUrK91/1rdhoiPSHzAnjZX91x2A0qACF+x1QPa
suTVUwZPAZ2x5gls/kCMFzEPqScnHmyrsUGXzD0d3x7RgZ8HGzgUK0mTAS00f9fT
PDVS9nMXkcJ0ecz8BPHOpRk2cfLAcpE+LeiRhoi7G9OHUslu6V14JQaC5CGS0TSI
G/tge3L8pzUgo0ghwOuqifRRzNcjmIhdNHwedp7dWLVmDMgCVjCtS1O39C949QZw
pB804D9jhGJB+bqESEAjGKnPZSnVTMCIg+QnV5hwnfPudWAl6wFSn6dp9/dDlxX3
SnKFqHJE56PxDuTT/A96fkj2rK9aTEvavGsLm+BRnOIx2So8anPAfcY8TV8xTZ0g
CN10qOvmq/U8gF951DTDH0s2xEZgi9wG3SpfL9cTqvA6fElnEcPxiY/dJsFT27sn
RgVshTwU82BVX+4gKI4pMguveQIkB+k8OL6CUpdWakHs9mCz9MRFzvUq0JiInRXp
aSzdFFH/nzgEJn8jvjRZva0hCRAEmOHOhBubunhwsZekenvARQTpp77fJL/V/ypm
3GhlCCTOyxtv34f5XwUwiiyn1bLhrIBZxBQuye23gKbIaIEptjinaQcNpHVOTDMO
COgRT6tpSTUgPVVIclAeDtwUxJdQiqJE/IMbkptY4u4jO/slyzAFYfUNzYUgOn5B
/yo2QegW/q8K8P9ilvMw67MScL1e2EWBxm7cG3BQlXV3Gqtb3Q2jZ5wzrRplSMSl
8MMYg2YOUOI5orr1q8cvsNeB0hHj1mWXCfdXl7UzXSkrCraWDjLmsG78Rc+M/Brs
Ph2rcnOd2q+e/CqwXwIck9ll5s+MmPDO9KMRBCh8msuKFmAJ4YAbFTDYMuNJUwfJ
7giHQ+IlacUGOp+VR1BNINd/3GEcAf/9pg+sLZVsQj7g/sBWjzFCU8e/LlTYHkLK
vLYaJdM88Pw3+R9xIsw3V3qp/9owwVOxbisZyGT1LdK+cb9y2GLfJ72/n4Lep7tN
O1kaRj3jJUF9KsCU2Kf79N/oT+NihVkenOf01d1Xztaos3AG918dFv5txGuCNh1k
KRX6W9eSIDFz/tqFEbDjWlFdVH0ewzOleHLBgsumDmid2tZhhu/43AELrpuCr4bb
5P/XNOXDMVQQrXwrEmJe0jL+xcI0aKRkkaYSzKjbp/w8ZoQbTI7WF0a7QkSCRuo+
f7LPfpaVxuxHiRJzqZXjalc9Mjdac4icIKUj7DPpPfZT+nc+pHEjsGCTfToQBcST
zSldE27vCxs4DOe+5L11U2GDi2V0TF1jwkD9WoTDfS0a0manGxkn173fdEt1+etF
4JWuIoqm41pea2jq8U3wrsrYIS4lp5ct2TMlwVqFRzq8Nud0vNftcI/Ak4Jy3Ak0
8n8evMAcpqcvRjA2wEqcCOhWNXrW1jKlPynTgRu4jwyvEHuLiO3Gp7nXddoKMI+s
mSSzq5K+jzsIWsGqLes1ubmnehnIQKx2kBdJlg6ldTrufl5+EYrqv+bN6hjXr4H7
Bc8yKjaZmhBxqtGBU258vthoE6JUJBHnF0cd9T8J4gs5cHzxl2MytFRcCmjDvGpJ
6hM4GZU+rbVYSI9mDAceHCMSo/2hACAh+Vyenb+yXyYe6xIsguwhbN1y8NYM+NZk
4ZdxxPDZPrYA/LzwKwW4TfAdAROTuPIsyIK20L61/HiIb8HPlrDLlusB+T5KI7sV
FPH52CefiZQm28d0wsInN16lGooE7VRxwUhGLVkHxFvxQ+1/SlVhUVWL+QtIbBE1
Qc7Kf/xzJw96Z+o1O2cXXLseqk/MIKTEMejorgXrxY6oEs9u1pW/OdP58TohG1dD
BLSCibnm6uK1HdMWUWI7jKfTpaVMzuOokOO0ytctpUS6zHjf10WZzpu6pFSeNwC5
2+C6HY/E7vU/ARAySfO2DCWNGBd31vX738FQnUe00IAYfC8xGAoSPiTl5H3EVoMF
35CoBg+yAPUta2X12SzBJvGkoqEkYTZBU5NK3mEGgCijgoTpaZ65LP7CWYRYsf7R
2WEGegkLqmCbOh5AWEOMUdyIlPyxp94ODsvlJHGhUCOcX5GTbRPr16HJhCcIy6NG
tx3PkjRnv1NB9cLb46Q/3d4PCFOnLicLK7NZ/CCwzfgYPSFV/28GM610nNPDwrN0
XjyZf6vZm139BT7RCoIJBlhuWx72VKDKZHI9wOO+XsLb3MOdBnkcP7C1hJqHb9hU
XWMnbweemzpzohCWa9e/F2GrHTp4xmSB84kkrQQP+qYeuc5H6Mi4514pG1mZQ4XA
kcN7UB8DTCtCzuJViKtgcHXtxiaWXLY9loNeZ/I5+XkwcEpCPu0usmw/lwiMMUu5
XubJib+o6TVX+sso/wnRLyo/v80nNamMd59kAjat+aByE/zYd2wcKSFHqmQ+SmeP
c5v3jZyCg2iBjYFobjFTeVDZ03BckSerLRVBWSNMisKU2HIoGK6p2I1b0M14oiS+
1S+S+77GTILW5ECeWxTVVHZK7Z2/9Yis11kyGi7aD2B7oXEpa35GGVIn80q715pC
iRwCc3HRukBvwRv6Wfmjs6t6AtIyXClyM15q//rlckiktmD6jWNPthGcFiqbP9WA
gIvFkSmM4+A5UCXp7rHn9ePnq7DdPkhFqBsg2ttBoXTjmNFHbrA0/xnbPfaJGsH4
xG0VJoH/IVv2YianOM3X0haPNANTwC0sSLL87t/Vq6yRgqABtiP6V4Xc17zBZff4
RHNgXUHERkqkmdRlsmwhCZtFMwaThmgorKrmBykhe1ZvMDydDOm5n7W28WfmulJM
bX2tO3ahuZIhkNzUP59oAgsCiqZiQJooB8z6ysdlO7ZinSGsDXosR40dSGPPkp9G
Od4PQgTN8rAMzol1/hpk5pCEVcoJZ2sKdOTjwVUmGc0bDAoCDAqrZE4zwXY8SOt1
wXvO4eogSvam1zqIY2HfVh0nh28xs7yqMDPWwG4q1AHLnt4g9EWuAVd5tnsWsqtX
NP8pV1IxgfqjipNeFnn/SMJimNsng6aURTIbkUgsSPYM7aTKr1FppIYnlazUQOhx
OYkFeJXg54wDxwpZIdkeGNMQKBDmEtvv+U8St3D/9WKKZAXP83loEgP37ZSeozs4
x8BwxSh9HXC+MGjZAxyLsjVKkRJ4dmhmM+ncYSc9kWBs3IAnngWYgpbf2ySzM6x5
4nFnYsZdTe4DfyKE/ZOFmkDYkMElpFIp70JuQ1XV72CWBXk7OYbTip7muI2qghTg
FdQ2GlASd0ClY7deFTbjfKkrsiczDdgJiaO0+O55/tUNl3+zem7RZ4Vx/xRncuJA
cA7PCMZ1MNl81yo3jSwaDNzpfYDUFwN7UFKsbcNSw/66Hj2Arh5eXsYeGcYE5Voo
QpRTe17qUzcefdTGt4FSbBe+lmpJ8seRzNvbdIXxIbaqvLKUg9OjcmMqWs6tHqgm
qVvzwBah1iOdSPHRw9D/xxGjTBH5/NA2BfMPyEXaR4wQ7QSjGZHuqStQiSPiousX
hSJ5BdtS+t6ia0Sr1K1UeUm/M6/gDNBp9caQ0miW2tS/Vi2yqUkEIjmUa2BhAUjc
FZDI5GZuOIt9oK34g0ZsJXD7MJeMVgG0xwxjOXk8cEIiR2QGwa6JE0MoalW3ID0f
E58Qo8GKMCJRGY2dwGQzCFRg0fUY0Qvq9Nat1d2I8qXO2rjJ9/jCi5Y3xdFLjtkk
QwVEal1ttbJOr9tZ+QTsQ28Zc5UjUTL5NRcb7uU+SfzAB5UCeyOFjPAuzDbDRSpe
1gT5SKVFFUcr9KqaEnVT16qt1ThdXw6pEQHTXcGm4pYv+C1G3cs6JP1LEo75B+Wu
VChaFS62TwhN4Yxx13PIkgrJzxntF7t74QrF6l6RZwd//oZzYafMthy88fHPAYc+
Wmmm0DgBuZibPdkXhH4nUfdJ8iPg5184R/ce4nKeiz+u48JdNqD+w1bjqwH7OBBl
65cih1oYObpr3EvI6dFeWyecOwuoC3ymkQFUqWBIyOCSrYxPJscWvXOj0YrCEGfQ
6QxZgDCJbo7gHj09B0SP/ZjbpjW/QqLZp6WRuXlNCANOp4AtwbXMQUcbT/AKbX2a
jmKheix8IVWcxLv5GlxUiWZbM1tfCq31WDKs2K3Oe17IXbDv3JG5LtXhp23Hr0h1
31+MA1jIV/POv3E0EilqthrJXikOLVxPJTS1/XHnrBMim+Nnq+M2iGa4LD4JluE9
m+moXhcjwgASHtPJAWj28Lvu6bivggO7+StAD/WDL2mmKcWazTAZQ5ldx1hw0R9e
sYdIHPkNCr8My1oJF7nff/Vdl28nb/whlyrRJTLgPfz80M0V1sZJdCJDnNYm+TwI
CPgV5sB+9OITYroU9i+Mtzp9/+WIXJ4zFixHasu176RlSuAxHQWoxLGWpa6kuJrL
ygO571isNlu9jDbt+GBi8l3Wz/j0XxEpGrLU0C5ltaLTtVO4kVrDAEQ9dpwJ27cC
YUwGaMp+6o4ncXHqEpulteG7zxKYIDTlllPbvycURoBiYmCD9CpRgADnAKGiADMK
XQvmSsL0zKNiAhqjtkfSRjevchPZBo3RVGk1dzvQUJT/FxAUShD6/RGO/jDJ2qz8
u5qkEwdJkjmOvyvdr/0H837bfxLBBH6LxPxivQGbeDABmzVBxYU+6CB8acvdDS75
SdmKFDUVGn80aJAxo16hJJJxL6bVyor1eRgwBQ8/rLC3ruRTrsjYb+utUAK+atRZ
SvZdDZ5r6waxW2Fna9o3zLuaQvFE5O0Ox7R+CnIT+oZoGBiS3Ni1fFxXwPsItsmn
ftv7KLrc7W9u2aiQouG7tiEFEgToyBSt//NJrsc9HACJ55suAgBnj2DWr2MB1JoP
EOpF7gV2IK/c2sgTuruejKAJuEct6ItOc3Jj1vl4n0dVoEScfLywUW2gD1j4Eqy7
DsvRRVG1WufEDaPgUYcLwonCMFZ0FsxnEJ7R2kM0dNEj2n07hcX0vIHhU2sDxxyv
TOrU4WBvxap2Aw48VM/mS+/+F+07S/yy/tL0BWaAjG34oGhXkY0Cbbwpxa+T947J
Dq87IX/4fNPQTlYKd1/ZhYNqzkZxpi33jGoRri1g0alO5lrKZS26eCqnPGzyzn9p
loo0Hka4bvY075RjIvAV91u1sc/7Ttr9NNqvy46SKMdoZ90FCFEAOm8HsHWys7Lw
FneXNQRjAkxUmK92xvKibGei2PBviTDWzHjxxavHEZYzrNCBleALpXaM+KhS1t4D
XF2OEkQAX5QeUU+cvraFWZZrJGUBXFsm0AFCpLh3rJidowyz5JKcSQ5Cg1YluvqU
RENagG6/jmxlOXUEUNTjvjjF99KGmyEJW1ZDFnYrumLgK5NCrw7K9OP8kbkg/SFj
k6sUiHiQVsgLPuhY4SogUQdoH+/QZ2hg2b8R2Bte1HByT2p9+FtGNRBDDruUfrGP
7UKxAb4DJApVhq0qe782AYs/NhRQgIAdKwLxxQLD/CesksJyi+3KUFSUvUMswsqC
ct0wLuBNJ0KJ5+5oomtJaTlENUAtmpHouhR5yLjrJrd3mIFAH7ib3PCWCpfkyfVA
nM+lvZ/6aUZ9dLbT7pYVjxZrIM9xliFPUy9KiPvHxMsr4epe8cgC6+xSgKemhWYT
CYO0uxh220AqomDQjkD6/eaEpgyikjWwasBPelFwKX7JH/Z65yt2USTcJY3kSxdY
UGJSvwGxKl/uKMgiygP20TYojlgICNOqXtroRfHUEktaKsipOQa+WGBsy/y85VT4
kQdUWQ2hH9M+FmrvMBRR7yGEshDqC2DeSBDskLIJ4aerswh16k+yud0zPCxq/ajA
Xld7B9l7MHuHs21eUFkfg0DJ1lWiBRoj+stb3vKoSiigdrT0z5m42wPIg5GRPIqJ
TI/UgipcobZwfoORYGNplD/wgJGlNX12soj4z28zb1pdIeivXV/E45Vi1r+xjLXX
OP7ozKp+ug/aZMGCVbvSYilkUsF2an10gacQS7aPcUiTpN5qyUnG78mIEkoC7SJr
aH9VGNNl/VTopaZS1IZnSD2aNFj1uVk4DWhn//R/Qvu5PdN/ZsFFGv6OEzftgjy0
nM7j+IPSxzELlA+Tow0qTIX9od9zKixcRHsyR2AeEIJSxR0iKLwE2XbaQzJyqsdf
RsRdJE5Q69pJfrRYcTrjYgVURX2uBoIUjavvQs/mGfgQauiYwbRIHaJkEDE0ctDv
P+KmQUty4OmZdrzlV6E0brgcm/scCOrCBvEqv7PoS6yH8W1hKy1L9aDArTC4RlVz
DTV8jPC2uaITvBw1/VPCv+S5YipBA5qEjfWRJakIBUoxBOzZY6qQdEV5bwy7rqVW
Xb8q1UkjYaFw1/uOzAmy4rVwZisa5BWyivcd5g1qvnYIBnJoc1PPC43r0+13lBCl
aRi6yp260xC4B5uwar1ReE260GtEFmf++p7ZcPBH0o7uKgKGwHk7TQYhTUIz1OFR
JVVb5cO04hVVEwbNNNIQhmQrVXxzt/91m4UxYk06RHa8C6JGlH/rO6PY5XRYySkV
WcIqke7jr3ozUZsdHed4FxCidHhA2OoblVWMD4AX71Gm+AR29LjdPrXKc01hiW3z
oVsN/g+AseeIUCo7sUzHSEATi5aydcHrzLQ+R2ObgV5Hd3SaLAqvAjHg+b0waQVn
yNI+1lSdEtUtjjv4eWGy8IesJ+5+r1Q2vr1lpM75U+osrJomDMvIJy3OgB/ICn8C
w99BPtgHdDaNV5+GDs8IAhI+Z9FvEVHrgR587T63WXxdmvyOC4VxP5opeVkA/cNJ
gFGw1pCrPIJz4EIr1EW4cTssl4vyZ/U0JYATTNxn7bJsszDdICGJ4Z8DviRhiHHo
t1c537xTDQp0PsdRi53ds9R8StosKWCSAoFY23IAzhhvsqnAFzJ0zqIm7oGYURSf
w6BpZAaa/9ludceyUP5CRo+vPNp8DmwweGAX7ukMT428eke9Fca6jChY/27ssTZI
+n+dlzI7fWZyeo/YgfEdSAicJXXsrQ6530Wm504dL6ErDgxkmDTt7HUsUJ8F1jW8
JjC547OiQa4hKeuswJ78h5uSasUUstKUMuM8I1vJAorBNVdiYO/DNvfkfhJscx62
1ittup11UgWnQebaLwg/spc4j8B5wJPMtnocZMRvg1QuPDDAHRcHUhfwKbSTs4ol
niRCoLxM3GbocOFxi5H5d4kgFSceIv0LEYUCR5q6dzaR+0xfK50r/H+luwGRAzX4
55yXWRDwnwoHApl/py2YqvCW2tobsLVnHGpV/6XNFLw5R3htkw/WEFmtnMVTfr5C
9zEHc6y13ZL/an6VpaqghhIHtsP6sClnrSYuXOQTPvaB6dL/ZpvlYSDo/ne0jWv/
dOaqDt/M24oKCn1wVOvMbB3YBg3jUrNfxINyEkUO6RREboFvxjLp+aqcgymJgVle
OnDylXZalArjIpwcSi6nQrnF9maR/TBR2Ftb14MMzjnrQshObYoM68Ew7lWajgAp
etYkKsJt0rmziVYM76fm8SRFT5WpTyAcdX3tesbj6PPFjyygZyPMbsP3R+zhUSEU
lASWq6JXxw/q63BFKfycM0LV3UbvMfgad6GMvxMu4buXTbLDRJs2R+GWCxgOZ6yd
jxYbC9Mc8Yvj0uMQwrEqbCINcwm9HUnt5B8YuEysGJTh4cAU/JfpjJeU4xO79gKq
zy8vCUyG5EDHdXEuQc4T3rD066yZvC0AGizyZ3EHKDvv2HpTmISQPcijVJwu92Kg
oeonxZahKRfJ6JV03uuprpch1MgfXut4OGzgc5pJDYjQs4nXh71H5YRpJZGdJjUl
slHycWBkv0pCSsdHrMIKLDY28s+96wqQNOXW9ho4UWxJ/ld5aYvy5PMSFRnHsrea
jAtJC+x9El2jO1r1HoICe/Y5GzDDDV8pa8Yk0hw+kgYHWClKekEjc8RbzA1ikBHe
/qZkwju1lcPERvzYcnAjUjBDnNUWPegNE91lrQEFVCq19Ika1Lvdi0E663hzRlcx
Duu1+nNMJdZM2MkadDO5ib1+/nfIFcIg9KvgoFJnPuED/DbZ9rfXu6FbhUSDkhL2
e1kVPeHB8nnIML8Y6vNj+5WXR9JSqRKh8gWdugskqnvTgbTMVuwbeOZ/FsVbaJSR
ivYpb72XzWXdLcdNMzu3Ll1ZZ6XZioLhhMQ698bxcY0H+L22WTAa66RUb8njCBEC
4DyNlsDaMcWqiXPlXSyfWeKFU2d0A1Mc3K9542pjHmBHSV8Zs7TzGAw7TZnBD8u+
5xKPgGhFYqJaGHZ4mDOyARClrJT2376Fv7q1n8tkcx/04RBUvjCK3hBX8qLUrs3D
4EGCupXT8zcWFr+DCOCrBqzSkThEz7m4T3tsJoj0siu70bCEZKUVEGRivlBnS1Rg
qfBOouXoHTjOIlSYihmq4kVRdOqngjdveeOLX+n5mfyAscnyt4RhHoU0iZxGlA7S
SIAbuDAtr7vLhUnPJASMrmswyAtotmIhYQu2Fy98pHsUa9cZyTMkp8C6m2DR5kVK
um4urYRQ7kenXZLCU4bPvUMcr8pyeT/bn5MtBaS1yMJdw7shspuvFonaTlC22TDn
1P3aaDN0M3iA16J2tBrQbhrXqtxi0/3hGDgh8xA0alxA4s6Jurq4kGPTHvjz4JTU
Yt4sx2KcHBks5ORUMMuMBFDyPIZagiZIW1nmjMglzKzLbtsD+xzP/9A28XNhIUlA
YZYYotAobWjxUbcHTCnwBKlND/p2qq0Jm89z6z2R/jpm7I79nU0ckis+T4amDCUO
91Hr/zWmDFDqA7lWoMoPsWcO9S7D3AFCharjZPlYzmJpGlkA39G406lJsITwK/zH
RyDupXIRd5Gv4hVuQ8fL7IuQ8ehYaGgPyZnDPIrsR3bHX8Dvyxl+tojVygex16uy
O6gIA9Ur54J2E61iwATHUgr4Od/D3IRW+XPkjbv958ueM3NUK9SUw/SccgUgJG7o
wUf02HdCmozO5x4ZDjWbSkOGmda0PJ/s8iUL5dYc+dEoR52XC19SECIPaEhOgLab
Y/H4YsWJoLYDqK65/KPvTvaW1hSDtyDS5+8t+8Z1JqwFmG/hRZb2QAEY/TPK9MzC
KA3H8zCtHMlAjYdpRkEI4grm6L9MXBJMgBQYhxQ4AZL3HWzZSzD8fOfCttLXfy/l
Z8vRTHjyvko378+RUUTdgrhXK47ZzO6GH1dFE/bm2/KmocAMZkeTL7Osc17R87vk
DlFsQChRM7AQaZcEHrPxBvjr+wEAhk0jLyv2c5pB/5ENCuDv3tg6nfDAt1ZeLGCu
29u0+FXg19yQ2H/Lb17LjcCUYUXaMjfAw2gmjJiVwR5+4Op2DLW2TnqPfPqHSTx+
lng3yotrYHTNaNyWam6nVdXD5Twc5A4+x4KMDZyKitfStp5oEtEYjEXps7d7ieIU
YrzZp8UAOm7mlpnLEI4cXaUH43VfUx6MjdRu28Jg/+vPVEicN9uG+Xbu8aFhTeOw
PYige+S5fhdggvFtQadT2SmTcpivNEU+khzlTFHH30MNXt9/Yddqv1R8FkxLJ00I
T7tU+5q4L/e+sSRyAMlEippaNSVRX4IKEpyV01OC104wXFJ5EQnU5HYjIaefiqff
EzYwbq8t8Q83tsD8b3kea0kOkL9VAy3WNlpomcNH8Kim5alVuEzQ8QZBoYqFLfU0
VHYry8zvXY6ckvAQL+EWI5BKF+5+3WODze4eS31jQz4ratzXrbslgH4O5wFKoKkC
fNNNEVIlsCwz29r+QyaPz2JeHZ59vlvWqg+md9pEZg4rbLzCjS3xU+Dok43SbKoO
F+3jJFSey6P8O0myjAFsQuzM00oyOdgqXSjK1yUjNeJT3wENyolio5EK+8LnQrrb
rdMUeRdBzkvcwLRgauFtkP40/oVZyKL0HSrLh0DVPgA1AxaGjgxBr9eVti/q5x/U
GCg08WPbKs87vpjmYgsbWZPTJgtqs84pmsKskGV/dP/OmF92LQFezXo8PIQdGa7D
o3KM8E5gNT786AuoS5gVpXLqOvjDp2ejdZMKwVzHruHKxcsqL8Cfd6g6VNzue/Je
U6QIhvoQw1KuAGOYIJEFjscKBQGtVENs8HOyAaQPmAMsoU2+/vxAR+i0Nk3SpniW
wj0BZmLhUmrPy+EvwI+1fCXLvRhDWZ8XTwW1us0ArsTe+Od9der1DAbg4Qncx6S2
fBA9gXl2/W5SAJ8Cwf/AncucqKIH+0G6R5rkeAmsKY3/TdP+YU8E/TDtZHePY5zH
rP6DJXkPK1VmZTOygfXTO9wef1LnUnZla6fNdaA51nAaLDKS43FXvmFhM/cTPmyE
6LD2TgNyu4eveA1AQNac2tufGSph4DhVOD6xq95CglAN6ifEXo8e1uEC3oFYBjLq
/I5CYs1hOFznTg6wnnCXntPbUm5kXjFP/pp/CyFj4viQXdTQPhYkWn7nh29mv+5j
nBH4cXOlGMpPtBqZef9no4sWXGNYEWkcdBARbNSxM/KEzoJD2lYP0eJfBQ+5KziB
2uCsDiJf6GrUtzOwg72XbTS+bZJSJ4OBfJlBF69Dz+fLVBCEdSmbwSg7rrO0c3kr
dw572DGm63Wh95KisN8lo+3M9jtpmcNIkxDZAFkrqjcDqZdA52u12uLVEmI7yD7u
G+NQqLI59oqm6iu+8ycS9nE0vVN8olXbog0idj6cVXVtO2MQwjtojTAtNeBRowIE
ZLKbq9u6azLUqvDF/dVESQn+usu3WapG93CYEpGh2wCM0G369Qcbdx0CbwuzOZWq
LUVozpBqD0JP5HGeVbYKpLOCPViJXVmwczecykxR441rzbEmHkQchZrx+UinpUjr
BOvqkDunrbbZTxXdmyTeUsHs6RU7Qg1i+8LLuBJFBeU5/X8bNGSjRiHwtSg880hk
Gl+955y4mZs4aiu+jnnQih/9y/6rv9bmwogFgy6JlqbGVnOOYckL6cxKG/fz1fKp
ipBtuvTNxtXFOBAXTro8CACiUuFytnca7cIdFqpS6kB9ZuLk6Sn/r7NaSN3XSn0d
Tl5ME3R87JJOVW9Ub2iK1KBzQ8+9Owg0IPDwXQmRA+M4WlFnRk/pd5QbF4xJhZQA
QSF3e8s+8+K+4FbS7GP73GuO38YcHFTrJa8g4B73xABhrLoGLysxM6hqfIqNxMqi
MYpvB3jiUmLkVNrcwiYi+2t+ZVojDQLG6K1oIiRadp3xe6IzrSkxFBVvW8w2Xq9d
XjKCT+ldWX3kVOIJYpL4U5Vjs8ooL/tMFfSNYpp50wIuhcfpPSCcaeQGAMfKEcBm
iqAkNYnoEhhf4l2t8QyziArTPKWyw/J3/Vy0x7CBY20l0Vsxi/Iu8AFI7aYEuz2V
2U2F9OrFMn68mcMrY7/3wUhcJ6nHKWkb9knMx9vNDdigvcyDPoexF0Q3Y9i9vhcU
=======
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11328 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JXz1+zHgF4n2s6TEZD4KtuQ
ATkS0e5WlIVeyjNZ91Ns34qy+0bb/YiNerGVxnowI0oeIz+VnS18aWL1l9+hLlc8
0B5WG9yjxV87BZmdnC8jBDQRqixpiULvuJYUq74hGxUVwsljUzqTHZ8CDj28xmM7
kwDwrCSh24GkA3q5IwGMzkMXXMhw6mZKB7j2JMy9nHvKj1ahMnTB62FF7bsQ5O9Y
mxIbDiZPL+fqMDrgxXTpKoqyHXqo7auZcy4jrY09k6eQ4PaiVtOXoBMXD5EleOmK
47LSE2xBOiVbqZQgUbZCdqxxOF5rKo7mzspqsZlOtOX9d1m8ktx/da+vK+VbFBN4
IYX2XybSbJCYREzR2OKm7lk8nuWV1zszHNG/bLHveIrxDsMv2pMZQW0ptJrxHQzm
VUTGb7t9Zh7QhOXT0eChvWnFv8l38cQVGKU/QUxYH1TVSPDuUkPpx3hjNGX6gYM1
WM1k+BHuts9skZhurEU0ScoSQmGRnYJpfjM9tP58BFPwiyupvUHWMRbZ2OyzuW64
DS8HKhiiD07jb6lq47UjnFfETHfE7zYSUH2b1lHziCLaaw8sfjKJdQQw0qE5DNFF
IgtkufCHdKGtSUMgzjcquG/3BBMHFgzAlppD8AMuh+avM9n7XfhVZ9p++GAlqbf5
Gm3pfl6XNl1bNE/HMMJ7SRy9ntEoz1yoQ74+ScZHbyceCeZEp/WnatamPBHF5pDp
TIc27wUsw2Q79XHLFDKd82iinNd5JOYUKQ+9Pt9mzLOwKFdnkm6mDyzBlvMKs1sM
zrz8WYvgk3NM4aFflGEgiKZDjoEeuUhtdN1Bzkdj1exWAnqkv4CHMVr0Dz12Otcz
98KVZRzKhmsjnKSdZsErlfGRFnNq8tSja/rcKBUHkr/tGAv5yrnPRt/9uyrSGQ/W
tzTQwOcFMi5rVX6PU2jjPbpVopt5Ro3cLkSXXR6W+EZzFfpGqNsmRVY54s4BV4HE
tkuWuzkV1VWEPvoDGB3J5MfUKII0FY+66fmE0jl3iuxRjG+zVqVJNHY5PfllHrlg
nIoDT5G3ViIkLA4FkFTgcuHre10O9xAa6Ho+PlsdzrEA9TQsKUgSW83DiVysI4NS
ljEf8QnKVnEA+MeQeUm6JKoAl3xCL8Uk/SpRZHfeiApeKI4TJBL+ElbmyYPPEhwY
qkcLM7ZP8F1jZ7psWbLqgC0BTD/qsWgEQwWbeW2sITEz3RYJ5H1Z3PwNW4hMDuSS
v0rTIRrs552Av2oOyTV6j64nGrYY286PKoSs/kyIFl0sktuFGPx2bUiSpzBhJpXo
OO01IjbsTspMh1Bm+aQvbnYoIiG4sdwnnIno2gA63gJZBTKbC71uFaEw3IQMk0pD
EFDvUFD///Xn+iugR2A//wATnfBBI4npTKxJqWawXB7D13Pd9jAw9ZcMkwZdCrJo
JgaBRx2zex/92TK8ULtQRIVrnezjInYZ1EytGcO6e73SEK55GBIJtN2Ds4ZNgDDw
KZ5+lPkbP20pdZ33zIRgfqJY6jT+S9osclbHtD3mAKwBDloNwdcRoPH7MWqz04aY
jWuSqvvmdTAgrakZnsuoYgS0JTmlWkKhtsKrQj8bq7c6jVkTiD82OykRsdLnG2+O
vgcYgO0H2aGyNnl37180IEfAmzdxvw5a6vsjZurykIn7kCh0QP8VUw5nXP4riNpd
zOQfkzHnezFN6sn9FrIw4hWpgHPPx/QB92ICOvNRpvSST4sIT0EqoL8QVrl1tQFd
eJ8t/I2+8GRMz8X2vzv0kZpA+a5SoGh14Uk2p5WviRHuhroHYwFyXGG+Kf7eOWHb
jJ7YUO5PnqcHXkGtSBOFBprGk1oo0wxSL/YYcskJMKCJWZNVdTLq21NX4jB6rw1n
1Xdcx7Pfpa/mEgz5/BXi/QoRgqaA5lkp5WApIe5icFS194Lde9MP9nJoGV3oKv84
Ex2K1JOkn4j68ks4AvsXyzj/n8pgmOU0kAVVB1O3zFK85VED7njFuXb4HWPk7voP
1azvagEEp0zqOIKAybSeiV7AF83qShT8CVgwSYMkP6numDZ4yEx1SHZCtkShWJDl
rXZqp3S9h/lpD9qge7RpzdaIJvFlPJ1vlDV73iDFCxFHeCjnim5LfREum5pxb7FY
V8UTP40kOM3lJ4J7B97MtZcZPsck+f2AMu4BQklWDx26HEHq4CFsAs1fRIICYJCV
z2wxLfIDvQAXy1iCPHVjryCIAkFYhW1wcalvqJKYM3r1vmNlQ4upzKuuH6ExFiVc
KotI9/9tK3sTK30zcXHFmqRod5TfQZbABLnABapiCIUE8o5F2WBVa91DhY5TVJxl
xLKwvXvUpP9JnoMS1MQfnr6lQD8SlrFKy+qZ64UKrSd/zqFcaIrwwGcMcBfgcXjp
prce3yZQa5PQfgoF/08etZtU2om5yeCvlv3Mo2VWK4gXHSeohPAs1lA5txbtqxME
AOY265OslRiNKAeA01S3CTC/ULONdQMNIIuO6NJCKonAps/y9SOkl+bU+GNsqtZh
EFzu7C6gcqfBSsgT/kc0kxvMVRJUwis/HfUUxFANunUJlO0c3iy8C97Ep9n8a2+i
n5J3NNgxsGVvq6Kv+zKXIz2ZqkJs3UZP7phSaO+0mdrWnPhN+k4K4RnUy4wuqHf+
AvaCqOf0Q/zC5pB42MVDGmRcp14+vCzOd0UsiES4wj6tlJBgLUhd3d5ZElvoaQeO
m01Zl7wIk+S+u/xdeZVZnjRfm+TqFEtu/jZQ1bkqLMXumR61WvbbSG21M8heM0KP
GvL+PJ+YGyII+jJN73Jt/FqsC5tcAHnKfzBJWWKrp3K/fWrijFgq2Sczzka5GRLm
1rxOm57TP2eaTuE7YaW+z0IxjHNKrmYtzzeujZs1JtFd1tFLLzXE391URFasrDFp
myOoZlWGUUjwV3lbbW9dn23YtdWLZ7ep3Yjry071wi36CTPEEeQewmA7Q+eZ9VQp
XFa1Q9KGkiDDERYOnEiWfgxysa6U2aT72YPvXAMfu+pyavzcqwDEhASN+bYc2cor
YKsJyUaAbzfR2A4Es1ndrM6ga48lHYmcpKelvpjZ3OwjB8aS+UFxs9ETBznx1dMO
xceu1oIhSQuurWNIKNSqq2SYhjKqNxz6EZ52u7FrsAgjirtx+ypqv8LVboID3Q/C
O48Wmui0XiQdQmilM2WX47aW1SGNWs6oJUOEAKg5kXk73bkHdMMilxSDuV0kBaWy
UwvgNYIfHMi5TMF9TqUmiAkL06oY2aW6cPPS+gm1drsfLi9G7pO5+OmDiZc5M3G+
skT4nsdQaz3ca2OSJbWsoSU6uSzm/rcNUBtkTO3TObo3is2HXuQDWkJwi4Nr2Hnv
CzXsAjKu1c72ctdIBKb5uZUc7jvrrnqWIeKE1S5YQRreZ0soBbmx88IJlwHpLC4k
r/b8GYvowGbQQ4amc/oOe2D3ADdjXlZ5/5z3UVH2OmXsc+YIRdU1J97TLbFT2NSt
t4jNkJdBXV/D83VBMLqL1pKiASxQsWvXIM/h07nDKnu9luVcpGWBf4bopvdvmuOV
zdxFL2uMEo9bM/s74MmH1ff6lcFNjTC88wDu5ofXsugQu7EacQlLK04V7sQIMV8v
gRn/hlvD0pL5xUd9rKOp0ES0U7BtdHy8Y4k+TqZjVqshybD0cDjZ8WgOUiJlZHPJ
mo5uqNbTJGyxuQo794VprmnqigX8p+Fu4/kWH4xgWlfQ1gGhAWPGAFTPzAsq4eT4
d3RLvEqFf1r9m2251uXIXBAENnqnm6UyN0c4OFGdbEVcsW5aL0ZGkas9QheF1hoy
xkkGHY4goUlz3+HCoPn82Ps/bRrdQUCVWfohY51do+V8edql/rQV7RKdRlbzVMqC
5l4M8JWkI3ofX6FxOjBgUAgdZVSzVYeNvv/sTTJc8efzDe9xoSLOgC/Y10/dcOIt
jo6PymYc4ITmFYPOtXFUa/CL7hNemit61S9IsD1vsVEz+AIau40XT+KLAXdwogTx
MfPPBZH3NxYRybo9eTKUM9YHXAFkfWoBoIpW0XXblVmlcdL7DxPFojHe56Wwk/9e
O8cr+aF5aJchM4fGBzDWg/lwvrMblzXb4/5KsiN64teWaPBqItg8+hV5de4rRR1F
vpPLaSIP7/HpCr3GqF2h9OfUStt5lvt0/nfIZzASviKIQFXk1ulwOh4lYXBekSfV
iD5NZph1/GWlWmZVJ6ZaBF1GYqVgILdwWWzO4u6hlrfwpobL/uAGj6axxwrBBm2X
vGaGwxiP1QB6t3rdrJAtbVFLs8lYaRYvSVaIldNzrRQYTkcjnPuZ4Sv+BfqCWSFu
hg98szBHCm8FUqxUMgRfnQ63jQ+U+oU2EQtTWmBuB8ZD54/JIm/xvDiXQ10C8Uvh
PybC6x2I6jIZno3IzO9rSBkJbVEt25jlVfzaqyr1HAPtfe+6Sgcr/h9jJLqNDEUU
Vg4bsSFgXsUL1rA5UrF4FN0Mfzpxbb+0lHkk213hmDKXm3mpW0MideLHx7ksvyqs
KkTEcP+89p6Zz8+1O5wnD5fFjTDgOh20uyrcla+agSv1v8oWqIYTBzRXWybHjlVP
tRXHr1LQ4m8eFTpQiksUH0WDD1Z8/fVM54WjgT3kKy1ZKKyMdHzpvR7eUPt5K+rZ
pPl8YOSTPXwW8XTiGWRdVW+vF4kdx2mumtqqnuR+C6ANKEa07EQSfI1M/r/7xbDB
gkEiWz82NwExt5yCalHQ+GW2WbTkHB2GIChgDKwZlh+EqVjxEJpNk5DiVUg8HMIm
t7U8EEDrF5nS1KkdnyK+JmUr3D6Ot75X19hwkhn4QjqDS8rsLeIgwuUUgAW6MnCi
LGJzYAksHaNaNeq0V3QbKF9XaHeZQi1aIzz+khwnGEhuddpp5kdDMdRVhOAnioZn
U68MBYeKR7W1L8bPWEtTBib3LlzteUtSdpTp/sBFnexvK3g7CoxIVxAhv9rZNxvv
IlEEDnIgDVFASZCsSvg6cc46lS4jDksRSjnTddwqZrEW9MBMYkYvQ1y+5hiIDgk/
ZE1T+sWLIBWnoqQOClKES8fHOc1mhLPMD3jGBl9siEtzizT7/hKx/o3DGpYj5g00
HerGvxCqELqqxRiH7iaCOZ/AsmLwXDLedwr54Uygl8rrOYvX7GqX15hZT8iOBxRh
T53XskQE01ZVEFhcKwTEPuDYY6OnuJtMNMwkKy2W0ScjQpVvxYFqdePRQGydQSIv
XCpOTAUK91d7/ZeTVg9jw/guYm6Q8m+MkY9kg/AacJfNST/V4oEYxk6qIy25zV6l
k43DU8B4rAY984wmC2wyLrGs5qZFrad/HJdvTsLXeEonoMRMgOeQmO9julzWv/Vy
DOdEGEj+BHjfi8shzsPwwa/5iRQjj9BiYoaei76iNpjmRa1xReqao/whUzOu1xjv
9MCIDdvmGJeVOCjlyxdH7CYbI+r0yUEzqS7Qug0LWOcptuESu3ThyzbtqnfLO4aI
FEDVxBhTBRcRnqNDUfdaTZxB97pEYlgDve4sGJ28BNhtJ1t2lM0e43a0QOk08mcG
aiY/0UJh/wqrbAo+bIoHSKI06b9+GpwcOE9ko/5C3tTPxwsDFbC7r+Bq1IgtghFA
KKo2RiVWlapQfM5B/QZtu8S2uniA6ZumOQPz13diLAOYOHvO3/6EyggYpGMGM7+9
RmO5PNH2nq/t3t8kGxlFZEp2F9SUqmiPbaARS596vplWlfaBkOjatljq7Cdo+GXc
RlfnIVGg96Hdce0PBfzUVdyB28q/p8/0W3zv7y7P3gXPPJKMKWdIQcgZ+x7OvuXu
tenjNrWgQFavAti1jxfcun2cE6DQbMSZRqiN/+HNgGX/deqZiRWYiyMjN9910A99
IUDTOgnZG3WPEl3vLSrknaKbBUV/XHz45MmYvhZfiW1cpXqudcd1bo4u/rygR9wV
tV9AN1LhBxEbMdAKlAjtjxsTha0HRIXKuUIhjvTBkK+ly6/c+PwB04/yrVXgJbsY
QH3+sTjb2M4iAzSY/kD/Am+BnHAPKXrmbJtOQSB7sCrpcDkVc/Jj/eXqVdBx0liu
uTBtcIhRruc6KORRx08RlmqTw9k+0S/2AomEvh7fnf2qr6MwafHHbQxbCWRIE4Qr
N5va/ikQWlYtwx9ClWevbTaio3dniuDyjG4IobKtPZ++HUUq/41bKrQDAweJhxOG
5nXmk8+Qh9qdhLmq42gjqtnUMY5/xhC4laFohHTWwj+TUHCIo4BuwQyQp5wBtpnQ
4/C3xwGwP78YwMZiVkSs/kXzu49M/ceEETqsBITFHpQy61XYP5ey9Yss0nWhiwdm
F2zgjTfi4OsoBIo5AJh4QzrLYCfK44yoB1S2vsjBw52sd5V5JIrLzuAJFzZnkHfr
HqvQnOSYxND76pVMK0qUrZ2E96QX5Z2PeUg4TGcWcm2wKG/eGM5Yc3U9+zdk+7a7
8UoW6B73iVANNMq038/xPNPStnJZlO7goZrYjK5+nNJKtmR57Wb4IrjKIeSzPOJ6
uiji2DK+hy1W6AEgVl1c86OTh2XU9lwW696TqjTNewWJoeXS7xJZHaCS6J5/eXK9
ikArkpCdVr2bH3wVJrrzFoF0KBYnyc4fgMcPgHFb2SWlep9Jej/tgyUMpUBRzzcr
q3AsT1RoWkJQZnv3JDWkmRRg4WP6LWw/XIgeIXK8d3Vj8r0G30Aa0jgIdxbrIzko
YkNRFec4R2CM7Rz6csSqAJPo1/CnREYwLiKNpmcVnz0gQMsfsQB2PJQc+PfdbP7v
mTAHTJhlgXYh1gkC8BpVC0Wa4jRLJ9CabSBrUpW4ChZLg8g/cZuVcwKbn0473PK5
MqQJm8YCHoRz/wrf3CMcQe8RW+T8hl6MceR5d1L6G0PaqqOQpfa/ScZZTCKMEo5N
Zs1Oc/u/wstNAb3K7xNTrPUllLlLCZLhB6wJc3rneXDH5pYdqpc1iYtnHUK8c+Te
haxYjP9Q23lA+NHfnmqmmjKLIPY/Z79KQ5+B0dvGchDQMznuf2LmDdkWnTkyWkdH
AZUUgFDNQU2/AMjeqeSrxfr7gE1nHBcYxopjstp9hD3MH49OKV/OYSc+iBxDZvYP
mYf+bylABR8lTrfm0Y4kSAHJrvkD4LL6aKlgynXagv9UnaKFre8IEwnZJlMXr7Nk
FmvwBjsUxiCbFl7F4WwX/jQrKnF/Ps/TPHr3Rq8Mu7cjHiTB105/hePgQcR1Ilpw
qXlmZaexrWbzpH5FGTCUwPS757M8Qm9CF5LG75fJKHHTwxlfahFGTm5W/K4T5iTE
RkMpXjU0Awo87RRUjbqnCZ+onsp/kP1bitYX6BAnVzXSzyikuaZhMz1B5dborQQi
7GeHGQpFHV1aWr0M1Ohi6sH7/M/JOJCwqal8EjkqR3dlVDbqqmTajJxJULu3glEQ
7dVV6j3HhccXC65HBqkGBX48wZAZP+c53Ym3+kb1jRGQ8v1LwqNvWrRNBeWXNgVP
1sbFTDV9Tjn8+oOWrzCh2MZfMrfwv2H95qQTGXVrXuIvgJGoSBoOosAsjNn8CQUT
WTwTKc+fSIRje5dXdvGN/VrveEWlwpQoE/8sQMX2GXjwc7pEcUJOYHyp6oAvoePD
1tlEt2FcO7rvAMggZ/RnheapQndE/PSWnQcPCMPFiRMl9LI84589hJP9M+ssjDcQ
9f3Gtf+7ki2kqwGFojsOG5OY3VdMKruylWuGzt+YsnVMks1Vaxh2GTg+PAD+tmt+
T7wl3jJZWrSueGmZYPTsmmRod6qRahj23jtaNRxrV1CJcDVCL2osNLIAn+gdgMGl
g6afWrTlw9NpYBFHeulmleBgcBNf0YQ3sk3X4d2RiCFbsgzcLvL4GAiPOZDOU+R3
Wv78l9ZBOuXMq7CrIZEJ9WBTueFKobZ61IJC02hbzGyhqe1/V653vcy2bBT/CGC1
9VdhOqrNmc8KqbVT/O8YHS0Vehfm5iuX7V+h223S+d6aPTKAo9DeY22m8bkycBTv
ncdpeH5OcKqXduajZCbTs/WEXdbhn/3/EGccydv7R8nc4vFyxox+rzK1riat6w7u
9197QzohUBRTvD0xlz4QpwUmmVAVyx7taM8OYAvHWcAUfZJeHxNcuEFRpQSyLYBo
r1Se0k5TpO+U3uW2HauG44ITSj3qcdl/bEJodTzpg6sGk50ABAByvgGy8XM4Jart
8H58QLkbF7ykcxguTLn5Frk34w1KiruvELrBwKgjVt1Xzsf7cFTaFa30hKmtsU8o
nRI6GZiLQpN1VxGt8dc7/6A6fhlLCi2GL2WHXTRigyNF474R8sbDjB0B+MpZr7Ee
OSti7WjZUU5eWwHTRB4k+3oYB8FybrXUOCbRfjFr86bMuuEXDuJ+Sz7cHCWXQKTQ
xBXnPcOx0b8vlZtu8A6Jdc+OQWDXmg8Ytdv4hdsIcA20CwE79s4tXBuGd7cg8IuB
NSZQ1ySdNawjbddlPR1URct7YcHBAWDvZISNXGjnonIUSYVUty/SfiJ+nF4TGy1u
WfUBJNVlhBFx/T+2HqTiyBFWcCPgWjKERKn0LJ3rJRB9i75ssKWRqh8ehepmdvCV
l6rxDbshKvm9yvRdixYPo1N1TY/NlC+uQbDH+ZJunOOqG5FGgwKvwxTjyl3HDOcb
8L5yg+AZ6sKU63aknlCw7XIaFy5wI6KK4AcjXbvKENJqh5XQdLBQsLkZqoYZ1Tb0
dF+RKrcl9NlnYhr3mwiCrMbuY0YKaR5isyuvq9yCs69tOL1L3oS+Y1defMUuPtXl
upNTJ+feb9Tn0Ez9RlMcKSIRteRPWCZGi14s5ey5qoPFdPAsq6bqYs7qD+lh+PCs
nHgXyQB6fKe1b6kSwSIGNocBcx0V5PUQdIac9HJXXEO1ZciRim4o3KMzVvroDTy0
zLUDZU0fNRUv3b5DDNzyQ6mra+Nd9Z6GsUah2XyeKbYpO8tEwufyfVSwrTLLvHiU
LsaiC3DmAyjHZpvRaGGVUlfafdyQTlpjVqT2ji2snwzZj7TSdMpzKvTQa8A5OqZd
H+7UY3p96993/L8603uCgIErw4tSjeSSm/SUFnygw46hoBPImDeLhQfwCpV5gpcK
fj9b1tX1M3/HGajcMXhVl3bHsSlJYFUa7suIzhLe3n2Rqr8mbDosS0kg0krl+ihE
u5stvVbTZd5f13FUvB0d/V7OipyF6PIrKrkrXY7JMfhVk9ZMo9gSW5ZMiIpPpvCX
UR8W4nHMv7qCyGm9ZzhQCkx3I4D1kE1h3S74kFr/p1d4HMPJB1i3xwZwjIlDsfER
6+yptYK3Ej4TYCQqUwtypCBfY0Ssv9lJ6zjAN6P1pvhWaj743Df7d0oOgs8Kl1Ep
u447AFeArcsBk4OXT52/TLF2UaN3gOncFJ5yj9LGCQ1fP9Ut04d4wqmoA9pdCbu4
exDK2KWO4JvH3aR+5PgHhIygHHt+K7619zoxQo8ftH7zKujrBJT5CIsRTRZTTj+e
NqCuSh54Rdn+NvIHdVyyiVX4/Vhng3b1ER+/1PSHKJSXU78Oop7sZ/gmb6fkCDtS
6b5Zz/xU21uzlGBzPCDqjua2LyIToks7VQByr4dtxmDcbLjag9QAhWq28CdmeUy6
oisXkpRQikIENTcZanJDqupVF3xUcAYFUuHe7bQlbaC/NpMCAVNrtu+hIIaqJToT
NWd3Peq8gAyftSh41TraN+vC07+GgfJErrrZvVrieXq4Cknv5ezYfpM+MjbhPMUn
P0qS7JuwnFhaIeNX/piktrPzau9HyXGct62fke4FXiEIFLsrDMPmZdKv3eyqt6Nh
zuxnyfqKErLgn7sZbJsHZ2XOgub5f1tfYNgYh9xiB2K9cokWO2RCU+OwvLZtzZTV
s8lUjomWZeXDpZ0/PG+lTC3ubnTjdMsbgq8dC0MSNlcl7eLVaJIVMsMIXc8TNAFP
i8Iozgnazj4IhcysJnQMwdIGB5tRWPT1s7OqvCsevyqV0yev9sbAjOTVevTxkoW8
KMieaBgjlbaVH5+q2zDuBEdK0Vsy+vqVFHW0xfEca6U3vh0Rpry1pNGs9M54EO9O
FNHIA1rhcSa12U/ayoCLbNhWS8WkNeL2YHOWlQ92S/ZEIcM184oZsVuScWhtoCjB
yc021jIbdEcQ36cbG2jUOpEHQkNmO2H4QR9hZaW79HQdPP+uaD7o+5uUR6YRRKE4
lcy20wOilmSwa2SIBSGWZMjQspJxMnX/0dyWo9ZMBR4ZmofTBxfyuhMVz85+2tiV
1tXita3V+vEKr2yP3FCr55aWNIIiIlJZcjmexvt4kHQtprgF8Bg5EN5HHRPRYkxu
PWGVB4rjP4X3A4T3hwYyZD6mQa9eKkCymm6suAPh0sLFMQ9JYMbwkkDn1p/gdn28
SyPFkYjpK2iBjs48MsSG98MZ7me61UFlBAdBUCwZFi1H4cFnqK89CeiDVZaGAIyZ
jopL/Eou9YvRbdSLAjYq3EfdoV+cnZ7blGb3z3szLD5heDlpt+Gaw/QhBeQeK3bH
WqgojOr9pHozqKNbrbsdo7Mg29vNPOOslsFWPS8gT2bDHOZ3OQ2q1075//evroxA
RNJej3e1rcsqVqGr74wACjsenQps9YhpIVS3TTF54MR01u3aDG4AwjOf5HLBJQ1k
VxJ+ifBdnTLgXDAVHwB/aqac4Vo2a/ZkEZzFzVYILWYwNYBML29jausvdwN6lc7J
/iQBEgtbG4ic4pBYxHrtgAbl4r6jvDUr4klTXszTUK9vJIrcRI0V09VTx7f/Tfwd
Xtgx4mmNGfNvCnaFLlUKf3cbXENkYoXcEoSl6Pd2SVEI6CULunmM8KucqEqEVlu1
NQxYXrhaO3gln+64CFlD4YVaLiL9oEPK/+QOJLpnTsuDzP0gmMGxldnPKjrbKrD0
/RdRH4y5gB9tGkVBLnGP8d2aP2Zi3nvP+CDUTg3/k+UTBgvCdsnvnKK3T79LlKRS
UY6rBa4I5jKNsaX/Sj6nalKz4SXN+oSnVfxInLAl4tY7FQUr5liusdFh/SXr2LON
lzdUTZXJ0lzChtelOPhV0hPMdaV3uljtPJQke/E11B1mqn/NK3taMAVdBavLbJ+t
mkSdcdrx15+hT7MI9LDp46Shh1ys7etcY/ghhDpIhho0lmAkZ+8VaDQFj5CndHZ6
FlDYPxOeIFIS6NBNIDZfQidx861J/YrhNuvjo0QVMhR2lxF6kPOco87CHhgHg5aU
I+an2BQ5PNa2IywXPDtUeYqvaojQg/7swy0pon7UyP1JQWELqEjKqkXao58AG7M4
PUZOYojtDQVZ2flA/RrCIhO425Nj0MEoCEPI2kEpDn+MJ01NEzJTfaip4e9vzEXP
/48en3F8Kgg6mEwnmCdvzHb3PcUkUlKEIURdU+s0T2yToFXDnT6MyhMDOjMuNi2/
2nF9VnSRoYqQcVyz82VzPB73xR97U6SrW1yYqHt5HDxop193OrgYe0YHlZLN2yqE
E2RW4e2PufwFP3pt73b9HK7IdarTw8WNFd18gM9D/NgweSwUP6fpgy3+xiqKiFIW
U/moSFeYWXUBn6SJ2fDYnPDeb1V0IvyXqtm0YJdrsjvQwMWmpXnOYDM8nPEAbOhI
VwAKRQ6PtXaM06cJz//LesgqtPHDbS9YvvBIQ9gun4i2fG+x3a5xzG5jMYsKuy6M
KW20IDQ8Q9O7ggurrMhVtwiAy0DjYl0LuPt/Ut0tzRWNASXuUhTLGb44q5S44Pzn
sY5T23LLmDpVFSpPhjLfhkApUuSxkJRepCtjoP4YixhTDvedmc5fz7Ck07bR8C+A
oXPDamR2tP0XHl32KS3cgCZ8mf+tVoVurUTAaRgtP7mtjoz+3mlO47OvC2Lr8kT9
BElW2dj0hnDqQyvrLBTdMlj5z0hKA6HX1nyAy7j0NsAjUMyVK4CtrDMTXyzsKuCy
yZDYbTN5FeG498ChQqtGS2Vkhsz+eLmK2iKpPeoK4cyoUaV9vq59zQZqLjqT1LtL
qZI/GIyTwYyHizIvkUZrYFNe5vtxx5GBnkDeViJ5GyaEgcLpHHRIXbqeH9g0Tho9
+7gGb3jcyUeVPftPg6bvHfAL8885smzgDdAhaswHd9frfUi+5NB8kJR17iEGvUnj
+oPthYGzQS6+GdpuNFgvrxJJI7mYq/Xy1Wf6MFu5va5t0GLmiTy4SXiIiMqUMd5t
QswyAh7jno+mTA5NYGr1e5xX/cPGlG2/+pZPTSI1wYO1JXQXPPIoV4i+2q9i1E2g
8MketDxRIyZ4nujF03MNgrF4jr1eP+be2LAy8K42rLCavGsP1avZDfp0MQ5ca/AM
fwhm2EW3Dk39+A0b5YNb/Yo9LSMMyT9pq79D+Yupehd24d+bG5DyndNgktc7l2qO
OVOz1I0nEBYKp5xRACS6Q4HXGNG7pg9NetIINhxA6/3aCdSz+46MEElDuv6iLDEu
E3qhqUL9Pjr0D9oru2l60NmoAfEw6hBA3haA5IeTe9k6zOGk+Ob88o75emyK8hde
tnlKU91gKkD5Yc1NJ2AT5j+PYwHDrUF9mxBh07Fk3mEarIv2upu3SwRuwMW8GOmF
4FWHnxX2f2icT5eD5nrc25shNtVIEVJf5jzpTmIRMVBlz3wxDfRS94+YNz+ebAdG
ZeN3icZC5xiXxdBpphT1tm1Spf0hye89iDJHKaROMnXQA5jxkT0TesYzcO5ifoCN
3yk464GeOyDuXbgickGIl2ULgpmzhIVsqAVBjk7Ae/AYCZ03U+NOqHN5quhChKi7
3AEoszoDmie6EhFwPGkGddBcr/bCFtidsZ3Gltpw9bQdNv0iTQHh/1O8kJUi4j0D
21Tk/r++S/5yf/Z7GXdWgmXvpJdQcpUrgHjjw47b1gmSoZi9qbjYUckbDZXjPXMY
ph5pHp3iyDe9BpuwI4Jyp6BXtI54WUwslvhT52YPxxz74RLMLgQUZUfbLFf+ssAu
zFLY67sxtxtqkFMYaJ3dcTxBfzKLGm/ysGXcBiGrp7ylHxBQye4vJqPhG/8/xLl/
NENPhr5Em3gM4Zo0U7QgojWaD/qJdn+gWj6d0LmvFKPzOwamY1CspBz0COWU5RDy
eLx4PsOk57PDcr0DtNJHWDYHKm0ivANdj0yYTqHauRk3a6J12ggNEhFpa63T3+BK
ZqkyiG89jAtrAGUXQrHrx/bpybwpSU1VQCHAf7vZt2VKtBiJFMN+3mKXZrjhbFcj
I8I3tanyyp96seQVoYzELYBwWNzSRHCGH5jHpJQlcfhkCwtkayG9zcHboYhz3zsP
z9dRXSuLiOSJ34u+AGh9BUf3BSG9j1OWuADClzG2N3437a6nWOaAjrI+n0r2IG9c
9jDk+17+99NJ/xJbs/VmbgLrhcXWF46/Pl94du9XARq11hxyqEU8Pc6OkelaO4CM
VG0/mwapTBVI9vHf8UQznbQ/frYPUXl/cX/NdA8DQgDmf/CPB9mGqEol178P4Us/
7O/X1K8eDCkkc+aEPuClMFHptHqH3c2SmfYBECANJp8ssWnMZM2bqI9B3Mj7gKZt
gnKwXXJia93guZ31q0Cwsf3qFWabaYGRSolAe64gM2Lkb0jyWTt4DDy7W0LQF+wc
BTK770YKtVpsuo/9A1WqkaBgISk5HkrOGWJIk7rA7bq/n5mL8apWJcVyKGpOfT1O
EDy1nVkFc2/vl3PoJhMcSB2hTsrQH/o4WiFcDilCCa7k6nNFZsDi32z+4Wq5smUc
Sj2xm1pnwKR6y6KRT56fGYtmAsCLmavXroDEWAvvTlraT1e6q8gWEhfPI9aYOPnl
S70Iu72ZR9xRnWB59N4GWHzuPswCFWo9yQzMOaWwDVCTXbHMLwRB0dhJnk+hByYJ
ZKag1IJutW7DFsk2lmi+KQgmbRZFMYBTOh6w3rhhoN+o+moDzas0SXz+vMHnI7Gt
k/tgjHRZC7ISvREsm9BJHtlWH7P8RIoNZ71sIbP1zA9JvAEb3KovFxzS+gUAZ3Zq
0TgxDZ0V2SvRMsV52VG0+0kSNvQnQj7VWdQIc+Pjy/KwGztsURxRIiXE9hryJ7J3
ZN6H7FG9u8600/RSfPakO6K+lHl6+7boeMNpDuQv83pi/YbuprEkPvhNpUDjiIee
PnPfBJRk/Wzcba6jVzM4m6aFLLE5EO6WYECILzfWXrFQTSWslXZZyWCdhuiDBJMI
cYiq2CAaXGcz1/mMBjtQdRuJ7gHDJ5Ng5StFTcdo5yrSWI3wW6u0KRrZKDE6GqHM
3ixIYIC5I4fQo3Z05tRKidDiF9IZ0d8UoJJj7JST16Hd4m7bk1mBK8OLG8Y7e+2J
ltJcG7w/WCgBdWSejPKHqZDzBOziMNuSofR0cpiRuMWDklS9JrE3/hwifJhVZ0tR
IPsrjdF6LseAXbvquTFnGy+oRNu+UpSWnWWrpxhq3pl4/+BbCXrnNmq72vV+gVHT
ZXP1mDtsk1D5s5QemsntaX7tOdCCaD6dv/HFuN+bOgA6VV1S+wn1Gs7EFkklyCOH
EXXWFFNr9/zBQF7EQh8Wx0nDb90DzmtVMCmM+T6qwhmkKYqyo5L3SzrDhBOferrl
I/assA3rTpWg2BDS2VaX7qdisCD1LGHd90um18TS7fKIJbGBCBZbbvYmksI6YEzQ
oHIPH4lnxoY7NVTv+Qsm2GcaYRHPkkmVw6PAAwGc86s5u2zyn4EfEcL9SsiL3wwf
L2IusRQmGv/uj2x4MvjVrC6dE9C6GRHk075GfT+wC7Xo8pT7z66vfX5wfdKpBRIW
vqPrjrGXAeu3J65v6Cag/HC2edotxxzaTdRb03O81yNgsjqxVbIpl4LpkTk2Rtfe
D543YsnSg3a7zf/h/dVZsVvwT2E8EY7v+hlRqc1CTpehN85IulIVXr2azTlMgtc+
VMEkMJHNv20s0WaOaN1Z2rOTWvXwuzisWsvRl3IzVgIxif3xpCJ94/SJ2sSmJ3Hw
pTOLVt0G4RGflJwH0wtYixsu5MA7gsGWV7t6iYhnOK8hQIuT5MjPljc4OimqUr1m
N5nsUxyGJydXX0/6vc66jyKJmryLjbEfKIhFh1WOGb8GWXuecP1zTfrqZsJvPyJ9
>>>>>>> 426889eb8ce467b9c9a9f74dd4af433c5046285c:deps/flexrio_deps/MacallanIFifo.vhd
`protect end_protected