`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8432 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIblwOHrDC/GFb3kYl7b/cVSSbDnwT140FXlEGhIZq8kxR
HBK+Phh4snuAqhXxBdl8dEA/bCJ0NIINixNE0ZT+lKL/z2qgDlx6jtn0+yeSRYDL
1JT4cGAkF0Qh1fVN9YRcd4otv3l2al50JobWaKbpmvIPFZB8PsshQiyavCgysxud
ohW2BM0OLkciUxGZh5LJubQctASnxNKKGPHFwD8GFeOwhuwmT6b+uD5TRaba3KQU
qC9F5sL1QSs3Y3yV96MIFpD87YlkJIhmzg5yJ7yAfuJAkwdz2yAD03mLpDBC749z
dInlKKRk/6iu+JvALQjSRM9XmGtmr+ZmRBFYmTin3jWljIpovZubx+uEvK5S/sFs
UejlczKKyrA7XijyG0SHclxnVPXV/7ud4uIufL+zwNwIsB1HnuBWc7id4IUdtZdt
G941CWuGCwPNPKZuqn0HaI7KE57pJv2YkcsYtSLZxiFME10hEQNgl2eaJCKbz97E
iHpx4MQg3/qHVnNHw0GIA2VHarfYB+zoZQEbPXQKe8KlC6WRfeUwZukW8CSZimiZ
7gEvWAFtiVS/4Q6PKR4ygsjKAEGTOfLLd+Vz6GBn4+5opDfJYYoVDFjf6aos5mCe
RD1OUHtk9swQmbbajAcPSk5OlOZvpYEmI4JGFSxawWXuLk6EMlmR7kfqS6Mjr8x4
wG/blznepdwTVdvurFZ9tUC+Ga9D6gN3fSRepwtON+SKaBOGByhH/nBZg392qP7l
HEzxntcuAtFB+KeVFIBX+pGo+viWkJ5AExs7jrJJignbepYGQVkFQjC1kc72mc6G
ZjtLNaMiJab+AjMNdcg/hSmlBlR+UsstizIsJ659inZalOePTxlvKMwYE0hWFjoV
jRf7nseTZHATnIlKYw/x+EgeyXO3JsMrvm5dhC35QrLTZkMuOa88wcvMIbTBNHhV
JVthUBUpRUQUsKjCLpQ6MAdQA1LBpW9TQh0bo1W3VZV0UJEqosruWMOW5INxj+ym
MKmVpbSeLbwqBwyhHRFSnPYaxlqQQWlHOjP3yLb2H+puZcYaoHuLWFY5kayhns1H
X8b4Jp0DY/uZvJsJnGbCol4Z/XWmuh/loqgrqxSUyJAOL/97HxlduNkAnl3EELH1
get0EgcHZNerGKz3mgsI7b7fDSjQ7ho1aTRMqKzz42Jte6QRoBql74gncLrwTCOw
W00UYhKHhkH71Rtd4nfJEEILwalp24yhg+7cfV3TERmWut16C6egwzB3LSZQxwgu
G4Cz24VxRMxD5xYNBRYowNHKTJkuqnZPwtdtADHjo6J/T0feZ9q0PLgNXQJEuY9+
5VFE1ASX09jjqC1p6iLD3VjKg8Rv20y2a+5kR1eeF6kKCTlHn4gVnFVw+xJ/oVi3
c9GRYLabNgwX9eT4igh0Vn9uo68PydUNpXYcDRx5JXW4hfvVQfX5AqBTy2Q/D+P8
4+CxWr1DmEbyCdyZztpjDoABhLSzQJULbCt3wR8VxBpsPw+854v7h2k1W5iszWxQ
5nMo3qAE5IVvGrQhM/aXWbiKrSO/RP5otVtcKylOL3nyZZMygTKCJwuSiumPVL5h
zFDMFotiIx3JT7ap3HHYj7ucLDlwveapC390YF+x6GC9URbUfwLZznUZ+a/qQ3DS
BNwtM04nXAeZaV1JzXOqpGphvAZkff8+HsxRkEo51c3p3evspQ1jnHQ0IhD/HGuO
zseeUBQp2UmJ6Tv9IDRHnWIA7WSR7tgcTpMsWw/KhljEaMvbp2VJdlRtgW+nPAcZ
l6lnhVDS06oUVD4pF7+5io0/QTnRHNhEyTqQx8kzpTpG6cTmYD4c3htPJxiNY1jr
aXPlTR/wGLPyMn7V/QDsc1PFjdRiPcxrsm3E1JSGxnF/Wn5JZSxFrqxIYwwDcqIm
YaYzTF/1im9hqsZD8FVREFnJW2f0zv20NE9VEhPktCzSEyvUqKgrxj52eNYGpYg+
GzX1+6EMJ99Q5NA4RGXq0ux2rFBzW0vVG0CixAOl5a9w/fkKiRnZBcwdpqtoDMNK
LM+9q29vYDLQoeLJ4lKAim0mPNbIXgQmqkW+zV/d4iUbXOlTOUrHrNIaFtj0lJeU
IS4roRV9KZYCJHtqZ7f6/pboDQqt4uQiE1OLTky1HK8gBVGX87L/y4Q8vEixZaj/
gToLNdezOSelUAPc5xJc7JfBeAL+GLsvFxq8tw7CU5RjStHdqR1PigSGWd0LaWpe
GlUjdfLMjNz9EIUXa6SDlbVfv+PRWXfpPi9mxKbWdGa1kAowl6uHnlogVSs1ReWi
lrOg4uZsN2bdUUW23sAn6EJSuc1f3M+SEI8BTlYKvR/gMhvbu48d9WNV6Ue8mdnz
++6a1iNQrOspiMAiUfeuLT4IjzVKfo1SOwvkwC4S/mHS1XciUMlWUZLaY03J/3Zs
6ccaRUFthnzFqboFZLz5a3RLUO1I45sYVQ46CgTOOIhhXPNPSgBjGUeJELAB8AiR
1C1sfyDrsdR14nR98CsqK+qOBVHDk/L7RSqzjdMehr8JKFMk87LJPNXBXEtsepHp
WEFq0Kh51LPBSBHWrkUbW/XDDXIuV/C35XZwOiJzYtinGCxpBoxMPxlnm7nLQ3h/
uS1XDNJGPDSMJK+MCLFfYaTUwx+jbkuiso2T2FntK2fWzgutcY5N//o+IABisDAg
uHwLh4OwlfbMU3fZdohia2L/uP+/EO6rThcQS+U3+V8MzucZODIMvXKP6ZTjaaS3
/CMN9nqqbiIzbxYii7yyx7v2UUefe1Ye6IHadFpf5bnaV/yXUUry04dgA4+o7Ww7
dONLaph9G8qMXdX+w40w2w/QlkEjpDvokMXxHcZ20j+17nxVV0/N7+j+fBXM/7yy
C06rC1ZrWZy882EM7V5/CiWsfMmFHCz5cnjB5rt1dsSXfgWxkTMTGLenSOZojoGx
Lyyl9c3K8ZBSIjUimYbJP5ihhWItDKPtTA5DqLfoB2mzo97IIfWqSTc4gufkIyZP
WsuqiHCm3LQCXlwCVcC8TPVwpNOqJGWREXL5F3Di+AvJD1zWvosk6ULMdu1GiX2u
KyU7HcGWNV0itCNyCsYvcMQI5bmJDOjlKEVD7pdm6EA5TFowkthKGK4jTUFlpCVu
L1FjFiaAwi2j2yQrLmVohFOULN64PsnfG3igI8baLbwkyZac6eaquKGPRzuT0C4t
XGkC7cgRBDvcQWgkmEVhzJtPOvKB/EXZVHGyMqsXL+9s6EhqXixtn7fIwvA+WHxw
m2VNFTfl5OrQbqxwnnGn9vZdydMR5NLOous0P96MRe6tfozOKaq6oN8xzJAhdE0H
AUnPAfp11XfGFVt40JzDxhjb3bOI4ye6F4k2mXG0YQbUG/M9yeTIGITnk433nYp8
cL4mVxgJzdmiMAWXlRPIXcpM3wUehw19egilTNRExaflkjmq1eLAXVR9bsoapM8a
XlSeOUfUcUTdR1xENoTfQr05bArF8zU9ODrbX2ihE4OYrb01VaqNWcljBrWP5hf2
h3+eGzCvnJ9w94PUpdqUiJ7sUusVpNYvp4k/9Nj9fTcKxZj+wBUZgiRt7B5xQ4XR
UnAwGquIPdEHAAGd1/2+KS41z4SoT8Mdc2czrDmpxr5RvmXiy5K0O2SiRv12qlC9
xd3iAaRUuok4N4KbjyXkom/Q1a41vnUxtNspMmagYDIblSi+rYHfmHUBVVG7vVAD
SK/ch6zUGkeH/gvVWWpBkg/NtCSnw9Q6wG08mZtipLQj3q70cFd7IbTtbRFcF9FN
QbAlEl5slbQ5297kGNUKhYsVsN7JhsYnpYcX/Ic7JmAUwjPS7o336z8eRBaTQRVv
L3SLokVBvSjnZ/xzNXxK68Bcf+Ik1+gV0v9PqHJIHoYOKRcJ/6Hyx+Z/sauYjEwJ
ShpmdE/VlN9dKdEjoqu4pnDFLlNHEvtvbBF9+psCRJ1E6hVVzRSS+eP3HQJKVCK+
PwHdQRmFGUTeZO4S8cddWu/Qtad79BMYTUnSU9wsGFCuxzgfnaBfPJixZHTtQrPv
JbgMdjRwCJhfYIm1tqEs8lZKTM8rzj6UGSLnm1P162Hez+7VVG61+ZkIxpD/XfH4
tToxTdU2RdvLW0rJQRnY//Nu3X+CsMzMXQuOd2D3UkmLIw0bGjNvxdxYp478JPrs
qpcb/eH+gMF7YvQY6pnCQ74XjgJFhDJy3XfuZ7hHsdrEFUt1br/BH0YB16u4ZTht
Yh3DjL0SOrdZ71mR3p8+0X8F0FI6KxE8WeJ2CiyCgcFn3dyLXoNYvvnpjOW8H5dV
Yn9/2lK+8YopAEEzTJC+Ec7Gviw2XD0YRfQKFoOQiQdxSoEB9XIK1Qq7P70qrKhs
KyD3C6VBQu91cnODM39FgBBVGI/5JnksfTo6aj9AVBKN0Jd1srepIgNwNCxfnb6R
wyVkLQlbTuGjEpO0W+WrdoFGfg8insbRQIj4mVPFBuYhgWSy3R77AwZxDVsC8ORS
OnNZuj1zU7SWLhgAQA8tg11G+VS1nW+foOQFGKlhpIDl/ZnsBg/5QsaIPrguH7Fu
c40F2ldQlfgJ2NtKu8pfMWYDuUqzjZ+hvmiKDbX04KBigUgLlmhlxAi5RJI3QRMZ
7lnbaNvH0CMZ13S9wYggqE6ATxEhzM4ya2biyaif8Oz75L6IlUK5WIUoOayx6J8d
RcMQIFHwupZA40vdt8PMcrevMbz1ZulL+sefoAC9wo1eHccsYVi+1RDoNQtdCRl+
d5JJLbZzhbx/P8yYkYGdL5VXqiE/D3ojITVP5pDTGAWpAiMTh314IAo9RkdansbE
GiM9pkkxbvy/okQDIMWIXQACGvATsKuONBIzoowBg18NKr7Qg5Zkx34/d1KzY9a+
mjW4Gsw95k+AThlJKfkXXOhf1Xgw4MqV/u/7Z1tG48vhU6gMowMmx9eUGKviGVg0
XHaBoJfoUsSJX08YChlpbre9XfGMRqiMZxMSZ35nPzTEe3UJZ1IkH96eWbWkgKST
dRzF3mepJ9+H0Ja58MnXhNNvALO8Z4sn5sVgcn9/3DnNiXskNSKvLzPYMbNGOIjk
YD/v3N0Wf2PuccjlLIM4uk8EINr4cHHT+HU94+vlwnxYIS0GtMAuzPttDKpGiRye
C3m3zsDBXdzogfb7D7cnM+TIveWPmAV4ZkbUmq2FkZyB3Ry5b6nxXqETamobnmO2
/WmKgcZ9EM7LMt+89w9PsnMH5ycwAmy3llb4c3CHOazN0lpJ7803qZ/IF90cyoux
xgjqMhd0bSlY13k6WiQ5AbYzGQT0R9Sm4umoNihwiLnAZylvmKD7NtM8IyFFBzM1
NClMz+2TBh/NFxl49HPNBf6oWplvb1DXZhqjDSncSCapopc/DbRknFg3LFzyn0Rs
1GroVFNcm3h2ZU0MyTz9sV2L9x/dmTVOsTGEQDhH2HGNopCb9rsahj+EWFefWcJf
gSBVXpByj/VbLAYM1w7wbQfRLPoHod3l/F8F8+wnhcRqeRKFmYUwW0EZZ5+YaIuK
jAy3zOJhyfFKLkjdK0O5g0xAvET4W5bM64BkHDffN1B67BhdXOTITNDPU9ScGj4I
w96ioGlTwYbUOGDEr+KBBgj2D0CRU3+MvxGTWmVgOlW6xltDp7RDV1EcKr/8ABPE
QfETnxmiNQTVEDO8XWRU8fWlXdL5YZtNVCQzUzAXSSKg38GqUTAdGlkljOJgb46e
gvt4uAXlGJxkgRiB6+P1PSEa/vGVweYSKsYeRBolpDR/dhKgLMQE5z6kvT3R4N1a
rJFZk8hJ4hoFUuti4Z/5WRlu46yotoh1TKvAdK9rqV/LaaXSDQcq7SZRi/MBl8ob
8ka6xvgNOA7LGka49faCEMYOo+U8lfI3ITfy9IuwgeQBrACIKPk+j6QOhmNeX6vh
g/MADrXTQfUW9m6Bn5ELERxE6OGF9EuNtoM9GQ9YHd0dRjABEOMzbT0JSLMINUeU
8qgx9DTZhL3ghXX22In3IPbqZpMa8aVTrLQYLmcmDVnESUGfOu8u2IpE0runk6V5
ieQSosqFn/UVN53jEtefHXH6jM1u+ZLY0sf+mZOK8rdA2jWjo1x7Ytgo+a2Jp+b1
F5RenAzPJgivcOJJj6g5MPvDGvvuuzLoxJGgfMmHpTd+oyL+ZcRCwf3gzQbEK4Cb
U66dIE17jfkIbelIcDSATovQKtu2yX+/ubs4qgsNcOhn9lmYQSVdLY/Ckpws91Ak
ZRpQzV2pHjWq8jUQfcglsajvDdy0GC+Q2FQ6eBduNYKhdSpvgohsIKacj8t+xcuI
RRu94hMC4YHUZUlSFGfow6+IPMLE5qgnJUoqW1IXETNVQUXijr7sqMLaHkzBvqDV
X48U5HGmkOpZ2kbNFL4HzjCiyMhpyyeGtCzAwdQtI/7TC2JTNR5dMdtIg6SPwAVQ
q2xsVYXLa99VxOoJ6iHf2c4Ze6/AEiOLbnUQ8Vcqf+Dh6eiBGHSSoyqEch8gaFna
oPN6zjlTsuVrcdQOuCkUbnMUFGsFM/8afoZ1+fvV6wApcD3OalhE4D5hJQxIpvBq
PL93nBoI0G5UXzU6uQOPaAX9DD9pOi2tsTM/0U19mLPov0Uqarg+VF3aqYAZNdyw
lTw3WAm6q+hsiR8l8VK0Xno1lLZlIK02FWT/vjD6HbGR3jGYyZFCd53gfOau8hMv
QWoGyt0PZdNXtvNcoxtUmJ3dwOUe57Yp3KJ8YOEy3JhJPb0XFj/XgCIwkruk7V/O
ozwZx4ngRDvxw+N6/A/kfd/SZxObi8bJ/rpDPUzMsjCOSGOKEWd+dRUNWKD9NVRY
LtF3jktI63LQukGRfT/RPyakrXCmLZ8Y1vx5rZMWYTpEuSHg7ZVRLvl3jQ9qqqFe
PKF2ZFpStB9mFP9xz5sr7Gg2hsgNuBKyJim6lCwxjyXeASZXHHSEM8DC3fcOGVYV
6ffI+J/EidncI//jzMhVJYvc2o2N9gYYtM0PkHUykFMwZy5pyuG57wKUp6BAyDlL
0p8VOPrMn6B9lYljLLxZozWqXFLzXUaJ73A29GKUFyYGRZsFychKbtuvwWak1eHu
J9K5vy254Z1XN5BTF/0rriUZchZeiQ9+mmLHGbsuZ7Ysxwnjdguz8coK/C69u/S+
BtvFVXCJ3bFFN4xahCR/XtWevVS4Rdw5N0YOV2CfztT26dsInMZtmDZWINX9c72f
HcS1R+9MVzIKGVXZ4hHhZhqpLiYeFAyeZxCp0TKv3O5+vCKXBuUSKLBcebm9t2DT
hnX9POFJ4jDGM61Z6wk6AlnzCjdps5JBBPpQoSGq3m4g9SK5RIPEnwW3UlWKBif4
oqcQK3SLZ+H3gQxUEYjNsalLIPUITDjyMM7aYd8ieu0udXSkbTp06YN5bQwyK0CF
K1foIacRlcuGkmBJ+THcyXlKJtkLS035J3EmlK74MEMpx70xa2e5mpvlrp92MRdL
E/tbZdP294WKt2AH8qOcLP5I5FQwBl4350aATH4ozvClDwuNPbQNH4R2GCfmh4Wz
akESkM4KON+CnZjUAgSH1o+IXXGOIofJ7GhnHPs5q7YbwlOtdJyc+vr7sWKWZBWo
YwEAeJly/M5QL2suKpRQzI+d+4MFYMAjjq/uhVm3OQtxlNOVdVlYAlciR4hjDmWT
wH1HOc+FUrFBB7BNw+1toEF7+38z94CxSOVOoO8H2T/RVFQe13J+F4uu26Buoqy9
grz+06plvf1J1PR+LZeiZwtxYeWJIbIMNhYuHHLnxLOFWjek7kbLPKHrFIP2UKeQ
cuAZg161uGu0Oi8i66+4O11Y3Kqfk+iSg65ST5uPCFuEhHo7tDTKXYcz2ROeJ+xH
dUd3NtRyKe8RS37iJCpH03NsXhWaL++mwOMyo4BEdTfrzM8JhSiNIBzZao03vMGN
8SIGvD360e0bZn2+vJ/PQeS4pUu4jEKCi3iDhuhihDoBI+r8Zwg/29CmQqdJaDIy
kBAAXw0PtfYZwL+dIl09ewcTeMZbU8WuRAkGdnkJAbGGciiRd2VMZIoOfyK22rNK
Twkq1olru3fCpl8EO86Olpd1JxQH7W1/FNtgAdGBvsmruvcNQcJTCr311v4L1i1O
fxCEHJBkGPIohuB5hTcVUTDSRHbOMfGwbf8eYqSUrNOdgTUPbhIbHgE2nYl1+U1T
sjX1fiP+FNkEZ1C5HAb9t0GCtbLdzss+1kd62SFQwRRrLl1c8Zut+g5Yqv9Na2t9
MME+84IQYGrYrCTNOzDu/9nWC3DuaMSoAQKtr8YJ62Uh+Jd9hwIYC1KN2B+typc2
3+fQ2lz/aEOvrpqq7FuhSXsiyUaGCtrkc4cFuToXLwv/5vUdjJKd62R0xjZNC7So
IIvLdyRMSOTvTTtnqlYty7OYPrftPSnQK1En7Omh32y1NgBs49YblR8Lu2M/pc3A
mzS4JVxo4rpoTnJq/UwUVuINapTMhKLy4B+1G3KSlxJIjKQylptENFjY5/EZWBzL
4ODlni12t6BGQLZLR3oIGT4Ufy/nPneB2FaZcxLJdZG6I8SWRMzt/YlIeO+MTelw
SyKIx1M/6G6ZN4orjPB3ENqkko71VTv1voyQcyoZd9nVTGhWV65YTw61djyjyRP5
Z7v7VBQgGr0J64fosnYlLLmIj7+nWjUR+sBje5vRlzGzK8/j5hsZd/okqBKqbo06
hkBTNDZwKjCN3skOXSyRaJtWrRvC+I2wJhkYWK2LnixaJb1w4ry1tLSqYVRXVkYT
YVZ4uzzA4cYjNI8h7B2vwPytzRWGcNeIjn9jNAcJu9UYKJjb0X/DesTgbwXf89U0
uX34oat7E2NTkU5tuxNVk/wg6oo9gp3z973Ac277k++isRah6+2fB+G3TE1AbLqJ
ES8OAPZ99wy9+se5Orli+LhTBgvzRwBadcUWy1bPHSxS4d95GjljNP7wmXrwlTJv
9Mm0Np1EEXgbBlVYGVyNsgPM0FOTsCbPWOCL2Q5EKJoZ4cGC4i75UUwt5huMvSMX
2vPA4OjGX7+SY19HSyejtia+GVFhhNrKJKQSg8bA+VBRLPDwEmVmE+A+wmmwezDO
lkeZTPHgV7GelBQi3joaQLlyvnO/FjzDBsNTxyKCaz39apNRDOiED2m6VQUA3lUK
MphkXVH1mRBplJipr6I9ilBcU6+uq76zAsTflp8iyn6+cMS4YYfSzzG/dCPsgLig
tq5Eu5AXexn8CKxr9scsLB/ku3IB9D7vlp/U4mw+fb3j24/Xr9f12h7IqyDDir8+
3J8wpYarEXnufyz2ATECDQD4ExowY3fcn1g6Nnv5/T9pZPu25RGx/gNkfjhohT12
KmGVjVGjuWEKFCIWqwnSs7aQwNQBBGgFSoyQX2tfktuTPA+6bjAX6SMYx90VRGG/
z6QhPHj6t98/MNei75d45Ry4RvDDLQsJKXnfl4cLMLdxdFR7GIxTctQvEYLPKm3L
mYtpHnrmiVal/IrRBumkKoVIbBk1elERSXyw+dfvTuXANHrHSjwB7fx9TEtLUzOc
VxJG38zx3DwXEeJJisUjeBqWXKWMmXsE399YsmDayj5uA3n8HY/00EVQKXLuwXTD
uA5/cOwi9m6wROhTEWsQuAF8xpmfX7WgeXDgFaXD5UwAfX146TkxJKrazgUB+C3D
ws8q9Mc3H2DoLISHp1l0hLXuHIBP1vTRjIkxV4BqsItsrR3mEGwCwy+2HiMHDdsM
QZiMUopMUjWPr/gNuOn49FB3NHPvI66FvMbSKt99dUjZGmjfHdWs0HE11NFvbfQD
AFIZ6Lide7szhxmVJ+civwyyrbq0q3ldhhuxCMNfE2oVmbisayfxHuODVKu9oxrw
YZ0BUd60guH//ht08O/l/cSA2fkYnaTAUJ7ZC4hoWgh+hU9wifnevZsYkFG0BqgN
0ZZ7ckMR+qZ6JP6CdBhfMvr1VBcXxR+a2dVYnZPJK6LRQs8OBluHUPol7sTKIjuw
6Ci6kqwCF4rSPqH1ASuMtUsY4WNX2FlYg/mtIhAKMMwHvxqnRLYmY3gKa4v9aVsq
mUWkvkx8QKIoQeMHxcE2WuCrM/igrk+O9rP/63D9GnpGv9bsXh9vFKjwqwqMqgcx
QfaTnyLnqoyRxh6XGzq1P6c7V/BU00e5W3SZgna1qF1SZFZXviCUdXsfEjM9K7Ud
62JDiMZ3AyBB5nGMc4kYqgNOSjKZIkzVdGxtOo/KxQW8f5xMqF8pXBBSQPu1wfLp
l7FHEatylj/rBzDKQ40xCtJ8kbu7uFKzKPGN/7Q59ZU/OardutmRjNddQdunOvYE
RCClkxkMFaOqaIdiCYDs/sDv7bq4K5HfsB6JCxOkX1Xi2jU+CpiU9YNqe0MTREG+
Z9b7TOdYfNf1cGK1Eo68JOmoHfCVdDvCD0k2hgB/eSOFk32e0nnqxaDtf/desp4r
4RUsDbBfoEL1wphgEFTE8riMRqTmOkXYWTsAVanR2o2kgze+tvrtLwVmcWIvlJSj
wxpwo0fhWU4Jbo8Ec+iUK0p3zw4UgofPc7sSdzeWcw8oH6XqMHw8JLCM5seRxQ+Z
ZFgRrX2gokgZiAV01Cg9B8gdLhiDKSyUI4edYyfZTs4mY+CCREA2rBogBb0YBXGQ
r4+xoskrNrM1wypHF//itv0acLiwGO3Pxd1Gs9r99lMOyv9lXWskJ7NWmfesePjK
DyzusdnCIpzk/N3jNgIKihutYC6eQhAmJI/YSsOZdTWbA3TSKEhY4TWap3HVrtAs
Iczooy2XybA3+awamI6MdZBxkVptyhJ0scmz6rZ6+2AxWkDCWrfF9MhcCNBhnO0j
2P3nXJrmztP6MeDxMBQ5wiSvtsYgfT9HmxfasX+jzSRzlav594/DKLB7CkYUbTQi
1nO5FRj9H7m1IlHkidqQzAPH6ffETfUVRLvx7A4aDpwlTpmk643nLa+wS+dW5kQs
ehhyEWcX2BsOcJSGznroYJMJkoarE9w/B4Yi5rLgmUolkzLgyz+kJwgzAcjwOL/d
C+6efKYjylHJvWvAHf6ZsT6ByZfQ8mOqpbqQfUlicd3Zn0xvVLEvfkSha/JbLt0R
Z8RMU1qjQq8N6UMFd1y0T8wD5D2AjSCqa6pv1Ah6t8jBZ31FIHgl30Psxn0muXLS
1d90nESCnGPZLUn3Hksf4bW1rlKsJfSqTiU3DgFxbU8=
`protect end_protected