`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1952 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
JqcB4Dlx24+2+JyzNOorx+I6w5eVeZLbUdsauWuiuAbdk1fsNdTSu1N+iOZyqzyd
TyiZDfhkc32zFmwPlBcpWwXjRd6bMzq8J5xoSn6eqoZ0r11SqIoqoJFr2Vs9ksOS
JIbby7iYJn+2nhfgfpLxVU/sPUepM5C/sp/f8K6ZwyFbV9rSvvcS5YUIkkrfqtOZ
gCEqRIh3XiO+ep06KQ5obBBCwF/ZpdyWXvNHiEpGZskq+N7vPja4ro/k0qgaxE5Z
SjZewnHeZM9KYtjsiBTAcfGaPwDVUunjV9CFHecoEwlbt8dS9L4vT7UcZHBk5w45
bbFBmpqVG7TpHCWCXz3j20CdAKePdcw6r1P9AGMQsOn9h3MKM72I9l//48fjqb7e
b+jg+8kZFj/AYdQneUuQYsS1gk1PQGZQRO24VOj8RR0yrsad1Xd8Vgz03g3I4zQ6
Eh5wgAX8S8RFOIp7BMKBDf7U0xLArbQJj78z5WSUzFoGuCgN42vp2YaDVa1+wZsZ
wGNCSdCBZuMESvprG+Qlux8l9FwIxdeJbG1YBJhQSHh2Q64QW8i6JGcUljuagxGG
BfdIZzRobvoYwarDEHQvUcT0az/XzslhPwBsN/k/JizcfeVBaOdYitrRSo6YPpAp
EqMaARvzdWVz/EW3UU4upis19FD/S4d5xRQvKD6YmRobU50tuSZ46QINnukyIUay
W1buxtzBxVnflyO6vW5bVZefN/q7spMMbDqzHgv6fPtLmHHwNkbHGFrt+QPnSBJy
niHCDHczYl13U+c+B0jyKI/VVDqD8DA0hfC2RqUZLFeT42NKjnNnBWxR0fMfHoKd
jrkVr7S0/dDefE4/Wpv2mAscJh2c4e/D+AZDeeOI+9s0ag8Lvicy7vdL7CEClULp
aAeVVb5NTtRlvwcnkyvx3v3jrs293Bdaa+ZJYsQ55etM++qpwDwnHaAOR/fhGdBr
ZZM+yahuHks7f7DQhUWCkizR4eC3zTascTN7MtfUicBI0RKBFlvsaRh5H+Bq36hC
BrUGoI6If4inwqNC9nxZNWuXO/PoaIUe0FK4KxugVxRixG86g+bSfPTOgUsX1RH2
eClQkzmpS8jW+xkjR2lE/J34lBrlf6Lv8k9A+YiUIoUNRcm7mUxoRcngU5ff3lmt
jXU14ywVwRMHW+DxrSYEyycEhzO4VbIzqIHsBgySlveEsy+Iht1BQNG1cYHPvxxF
5BwUE3CWWlXQhk3KDCUHaebN7yj6NVviv16I30wwzKIXDOMkPzzMwEgtHHAbCGxx
O/g6qprSCUdT7CQS3unekEjZWQwYM0vVviu5YAA10h1+Ov+4cEpyaY2hZ0gAIQ2G
+7c1BAXQPM9ncJzAjBBR3sGf7hWX4TziJL+XeY43ksUJuSEmJ/3Yw0HiqYNeDdWF
tM1SVOFRfU1Vqkh19abjVnsMVO0WMSZVq8yizCiYQwR9o7aaKJQ51S+lci3Z59m4
by57uRtbZQSAMyDVm5sLvbsE8AftaZJoFOHE1kyBtOg5k0PuUtzFGx/1HYUfonT+
dYW7RoAX9klUapfHJM/UamRw7I1By45fXisva+FdRFbalZgZn5XTSSvK5BOu+15M
4y5BLs1F1zLqzMcAarmkjYdy7YRzNWW/ImibNK7yHwWNylL1+w3YUnE4sn5EoqIl
y1h1zZkDVq/jcOdgftnnQac8625SvgzjyKQ2j7WJrRaoAhp/XZ7i/3TP2hCl8lLU
H48mUDXBXUZrRhervjSlXsI4H9wa5HdcNMrPPR0R/uJ5jmnh7Y9Y07BOP8ioo3DC
XmxXMN02zUii5UdVgwyjuK9sIGqV3+bAKhIViL1P2N4OlrGSmo5I5A05HzPbb6F1
EPzgx4kb7huapJUWzBM2qh0Y+HcWZ9FkBcWVXPIs06rWoP4whPUkqa1fUNK2GWCc
h0k+ysSTPaVekE/Qe1f7HJirR16TcWrlxxUTts8a3iVpTtYZmZmxKI8ht/q10/Qj
jGiO3C8BdIFG9FSjE9ia6flohrPEODQcVIf4lZ0m5G/cKPqhN0d5ZFtymJURQrGU
e/NpbFANPy1JX6t3jG52Ib/cV/o9xCBVHjZdCD8gnboUrpZjr+igAGF3mvBM9+dR
w6Xv7NBGPCReMglIZErsTTQgo620JYX2seHWnGfVOZid7CAV09gtlaV7/nhkruWZ
YlD9XHgTIlLMXxb1yCztIFvXWRjjm/+LZ2BQE3KOY604PvNBQdc+USD+HJNEFUxl
ldFCcgWYXEexhz0OTUsb1IMhsYFMfVU+deB6hrMJLJBZ7/fNGANL+U1hvNXI67Oz
LrzLzHJaRRSFRNbC65frHm5iEhWrc9IsXggtRX00BRCMqiwfU8VlO5WkG4ZDxBfs
jHHj5ZL5OTnqaV12unMDDbZFRNCOF801qLRf2d4FYwYYL/tG0DdWBSm5O6/3jRaR
2oM8NzQB0m8Y4+m5vWsYt725OFXj8m1Hn+g7cufv/OU=
`protect end_protected