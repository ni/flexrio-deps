`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7824 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JXz1+zHgF4n2s6TEZD4KtuQ
ATkS0e5WlIVeyjNZ91Ns3zPqH8XsHq5wEswhDHC+TXnLRWt0zvL7d1Sg+MVoKhNN
2dAVF4V37ZEJiU/hX3YYDWxYi452CjC+DORbTcfR4+VIic5Utg7Lh5MYfXqptvnH
ixZ61chzq9egcqRvdkxxYv5jD+8wveqFqHCEQRW4VhnLYVsSYuzTjfmVqpZgLv8r
GAhQIJOLgWZeWK8T+Hc4ctWvOYpgnGAuX0UlPNePYDPhbmxwx8ufNJZpYQtVKiNL
JHYF4XQsmIMKbqRC7Hj0LSX01mo6tPKimm7uN5HjwYbOiqNTPg5S6iDNvpGNSfUP
u4F63uc+cDYebGpFxXEb282GdIdoy1hDl2DxZ/Acp+Xs5e0v635Uz0V6u8RW7fBZ
v0yWjtcKDKFznV6LoeuBl7zlQUMtnp2Bd3WdeZEL/9bhGFcHiS/72/fomCxLKqn5
Y+tyWSx9cwZPSxZZCSDzJXgHoNUvwDFvhVSLjm3ieuR3QmMgLbji7joJZK7k1a+f
GuPjC9eCLRG0G0LcqNNJ03Pq1IKBVicpW89TLEs6H7ZW3MUeqrImzWJ9IGY8RXsX
uzzBKc81Q4MGtp5i2fr5jtNCC0GEP8Fda0Jvz5nrxIf7w3J7yMaKSrQR1g3rmipt
mpGok/agJiWCi06ufSO/VSf+9vwyGlcfd1/NRwbijNSJEgfE6CcJlgmYHXEgUtK+
8FIjwii+uPvMaC7kHD6JLE+uJJGuyCgIrtAqBB6XUHkJmx+W7ATlP0IyGZiUlAAJ
zuZUuJHJAo9FPmYhtfUFOcMO3LnK8Fh2WjMZhx9dBm0oC2r4Ca2H3KPKn0UwLwzs
Hf246/LwWJIh0cwDxhQ+V3kKD/A+yWn+MDTbNQ5LcOgbrzYbiB1NRDK627lYc9hl
5RZ41sBCqrHoA/K+go8Q21hAhku9S4xuv7upoUHMbA3HHBUIpnAW3Y5x+dMMM5mD
V6yCxpPnVP24QeJDaHEfF+lKlf1DdkAZgjWhkEvUBsTSC5luPn5Vro+K7s2JB1Et
EX4dMnAzErsEtKjsG6B8p/9EqafZCXgm39dYb2+qfczsN8FuWG4mGdiw++nkpnX6
YflyGr0WqBiUaLf34vLNDIzIypvOqVthUNw903J9OpFLE+2jjtC9KFmH+4PYuT5E
1uW0XvWnlQr8qimUvl8wdZdg38pT/z2xVhFvGTvkbEDlBUBsmSWnGQ5GKK6Cshfe
9/EvuJK7WSm+/v6aRseiw87kAaXO8R3vv49saqKHDxf2FY+8/BItUOXUJJSGVA5O
PlNiI0yDRuIsXxRn1mlOjvdxWhxP2OTCEa+okCszUs8w62IiXQJEM8HgSacPLvI9
fQjm6VXlXBIOaq9SbAcpZKS78ygfF1iDp036kp4t29lClL+hVVMrmFashfOdyAbc
6h9qtbbC9QeTA8a8nX4T2GZPIW5kccszkClcKoE1XEO1xlTsoB5QtZNwXb/llnyr
tGy26fiMqLR/rlsQ1FesTZ6elEpQZEGbEQ8kD1u+wT10fcVO8EK7TU5a6hxIwzvq
C5UFDoc16kaa6MwUBOuI6GQvbDCLv+pIWEcHGLAa0JQPOPHOsQeGPu9LiGyvWKT+
PSEGGzwDEpCrbcUdim/d2/Zh5Sybj2cxqejnH/Ltd0lUbVoIN4eyQ9d1BY2GqqdZ
0LtLAEMDd7WfrqarA9iy+wghs7a37BUViaiVaCsOnHydfSBfs23csRaZ6fjzlE+y
bQ/FPvZiJlE7ZMDCO9An6DdDWPY1k7FIOJs75COM6OMVFBTo6oHPl1Lc+f1/lhA2
7BpVdDq3hzXJ0O+XKJKTBFOSVt2t3ALjdQ4eZgPksveaR5gLCr9SBb08E+8Iyd7C
RPSTyu+SJ8wCeRsel5Chzcvav8ETHkr6XiHhqI1dISYPobkmVU9300PMKcYqeEMl
Qhhv2+jAba6SOENGe4Yxy7vFXGJfN0My2IfkS3LZgC7/0KvTT0bcg0zx+4TAqeEs
vLURlmEwxRVCsPAFNGPHLBenqr47y9KKRl8RaeJllLoXCdMRh14x3zzM4nFTg9yW
qng9PcdfuAiClEO1qmDj0I7At4vELtAI8EiJMZ+kuSBJTNxlujndvbq+pNiJUjVW
Mqw3Q+KHWX5N346kfLGxZ7aQ0+kFgIeYHfNBSkFHNK96s2mqjSaeJEMoJ8GYv+EQ
+rOi2qsqhfCx7R+8Meinf/z+jmJSeE03KaFoNjtFkW3mt8vzHASWw8eP3RM8p10H
oLlPHEXDeFDcTULp9/n9ESuX2rdW7/2cIwI75unC8WYRG6ixbrWC/Kkugh4NPZnM
UtJIxzhiaXRJYNl3BNOW7oAgPXyVXa/KaIIGvzHgY/IIj+UV2MwpCDyfp+ocPmB8
u7L/rTjUKIPfpHSdKCYXwszH4u7o+wazeyNiSzRsF8q9HjoVJzT93nKGmOqKn+eL
3+dxnV1zTmfXcV9p+Mko9eNozmKAWmf0pbiLFBdylLacsg7le+A8E33hvXMojt7A
gO/nICrLY+QtvsqvUoxfuQTrh7WZVuOZQ/lA5tAzAE0sRHxnWiEtrkX/rBLWTGy6
QQyPt8h20Euq2ea2JLaJEVjxq836yMlK5byO9vApQZQea1rSsJDY8mTlIkQemDNB
hAsawgXnuQxmXE0VB6Kn7XZVnEHhhwW2/qysO1O4wGMKz6waKaut079UAaddv+o1
ahXLOS4yZMOfk15IV/OFwp+vUE+3mUa2T2q6lzBOyaAr/TjmKVyPkElFaAbCreM7
mSFqYjoXGJnTyRN3RObjXsrDnTxYPW/Ey7ju45WyKrz0XNKkPYvc+ChunjAvNCjz
p7WrH64Vb+X43w4UFR9UQF3E5IK4R7Dg5fFDlpkL6jnbVpi27UHSzfwzA0ePsrgE
QTu6ei2RotjV4ZA+TxcUeLeVvHg5uOjTN0e/4WYEO6u88qkHjgHe4HKO/+A9pjVm
8MmCiLkhjJfu/bmDMUiBfVBQWGK6mssL/nN/RJhWBA1nOnZa5Z1EY4Cqk6ZL0e/D
Kk/n/1nBnfIHC97+oO28zhMBCdsDYs2CtVgkEz7CYxKUP0RA27S+RRo6ye0H30Tv
Aihr7sSzKSRFv4/HOb1xLIFZzI5PSTxsTbWxsONeyIavX4Y6FNhOT45ZGFPCijgS
02yJR0BrX/+0wyxE0qE3CAERwWGonZGOGswrrEZH+BtNEegJ8TokbSOzjAI/i4A8
iSHzyHRc2SmqfHz5hg7qgMSr1aTGpVrQmGUi1R8cnelsE4fYgPHDUf2T+ZyVZrMY
UQCyqcaNkZcuZPT7vzY0aBbG+ZAJV+QtBxLrE7iMzNuUkNwYl+CPOQh5Urg++b6/
z7GwnTOHuLfmZvnNTr0lewQ1goaOKGUm1xORTNe0sZP8fkVcfyIXGmIAkCUD7ZuN
8wQMXzd/TTjDLDM749WeFXLcvqWXm5AkYLrRSh2kGX1wF+sKvrz2bHjtTz2OsVy+
t1JMMl19tyeS40ogQwj7k9sTYy+HY7brtnUhmYQ1UUFRgTkP1MFwx9sKEWx+PzMi
/soR6e4jrX16TBwMHSXM6ikagchmRRhhAbjWWP9YO5fLG/3dX7H/wn1U1UYtKpiQ
tbIW4Gc/5+tNU2LuIX6eWUbgm1Ybjv+PjVAWZtBhev0LtXykSQIjkwGP1GTRMXzP
SuzGpvwwoDXppgN+p0HmCQKeGiXx6lcaptuXAHtY0HvWkmpDg3ZCSPlu5irlbI6H
aDxSv8Lml+2m/6nKTJkMO1vb/y3Q5Ib63ieu8AHejrBe7wVseF9J4lqu6oC5oJKf
lEBOuZZ6gEdvJrhqSml/x4Mp5X+WRi7pn7NOmzPsXgNsdnQvX3UFmdmJU2chnqJd
o0aAdY1new9rCiNeu/ZbRFS59cqBQoa4gb/Q9iPZV1tmqZfDEd2auIqPC/s7iLgO
8rFCuxadxD7UfzXQLQMGlrtdP7V0xgyHe+weC5hKh3eQ5uKz0IiqiN1RZpkqWuy7
uW1WxXR2eM6es4mS67Y7Fzlzw0Ynk5ud6zLaUqt/Du0GHyksRsvq0zFs0jJ/zEkE
fl36oVzvr+nTQJECKpneNspADxzkDVBuF4LUBLBJCzyG+2kmV74O/BTAP0yj3/dX
pTcVYCmsr3uPuedTVcWCtmBpyVX8w5ykv10i/1jYDYcgdMOge6/s+soRm+hXkGDh
mmq2fwRK+fo0YHNuEDfcYMVzQhBHTq1D1cHxkhuzqguo9Gcs1xJySCCANbQk3qcp
rgp5Iq/8Xzp8uBWOHcbrnVwPdj5wFfZJlpu2mGpeRz+zcPJV2L7mf5lcS/+ryRqM
D+XI+OxOGj5a+sdGRENNUWDS71v3c19UPZfYQQt1gUxvVXssVWCYgjQn4DTfChXe
TXdb2EEaQ0kOfUczELhTobAW/0jBGMAkkDB4QMCsHWcwR9ehnIzWH86uuZizKnNJ
Sl51Ov/6gFZDac2lbINHZFYcI8fl2DwFyrsGpNg2rP/W13F6f8sIk0xHMRNjEp5h
kYHbSaiN1haO8OJliXvRya5cpMLhj5QXa55PjWtGixtdt276loagY0D0z/iQftbf
jv1rMgl/IUnbBaVE2Hil84Uznwp78B7ZJ4hkoqTwgBpE6ZPtUR0b2l6N7L8i8GVE
SjEtuWYHt2kZUiQKIZSZs5Z3OQpfib5ju/HtwD6PQ4eGtIe0+lsnvLYraJM+lMTE
CWirIV517aiUpF95Ysk5fgY4erfJ0kS59Ie2SJj/Arm+mRQMdeNJsqw7d5d5GQPq
+OI8BZGn2xP+endc7pX20FfYvbI3B7LesnlX+r5y7On5uAyobySRYNcEMrZFa5Oa
J1+zb7ICAMxcgfKMSYZ5FXqZQzttaM8707hinLw8HEhGC+OqzaVYzQ3wncQMacXV
VMloEbiI9yaDthAk+e6sPSCBPYk2NoxxKu6IqaIUp2d286390pym7E4JIs7ZfVmt
Z3f4rj/JCt7gwumoXZmyabXEIJNkzP0+SpFY85O6qRsM9R6v7cM/JzptsxOmg0NV
pfc12YsI3+OyINjGNg4ilBt7E7RgZNX/bQJReqj3vu8pkUY8nAoay71esos0+l7p
6x7lSDCP/FkQql0opnLKoAWOkiaoWFuxDGvoKt0LX2JiWiVBoJMDay+T64BDtUXa
HlM11YaoK6vQYlqvkCy2yeaSSyagNOzs+4vC+bib3WEVOV8ftI7swtqZxzeK7EJh
nF5A4vjRSqKuhjZWPiGu3Q88kC7St2o6rTv5h2Fpr6mItuHXKwkQb20f+a0uMy6A
VptPVhPxlR37ZznU2IusJTMe3+d9cBO3iRgPWpp5EVHYAqOovxv5RW5m9qN8uZxt
6G4kxPxPdTGmtq+4+hoftP/yFTrArtBKIfPFrGiR5VFCTG6zS4YkdTTYshvYuRCb
yU+ONOQSXV0Psngq0lvFzKiZC0obS9FoDm2ElK+Qi5QRcV5rFP8M8xaVNrwJdtVP
W127CzcRZ092Ll2JvEPQ3EiJ28srxSaKdxfyvNJXGtBxh6eSVtSfeZeVGRqu3udD
qbc1Nwa6PIyvlOsnSk5cLCLmYXenqRkHDIKNMTbGXmBJtDkj7sEveIxp5K9y5ydc
fSBnLu++hzA2OMiQcIYk6qXMJW3SGSfdTxeH1mi72qV34o2je0LKJNuQyZIwD26y
SQGtJNhrBf0y1cC7yLGembQs+BdnUWQDRcNr/kXf5AdJKY8xld9mQQkS3DZWzzVL
YGT4GRuVjTxIEvBgoHBg/eXjSRaSzkye4+PMgmuuopTS8WD7Skeew19TTlgsQjYQ
RyhyH+vZTJaKoNtdrovlDt8KEKptuB40hDWSTmeV6+gBALWDdfTUIAbYJLjHqP8L
aUqDptoIARE6vNKOdCVZO1PkE8X2tA4HUpYfs4ueDFnaQmblogEcZfP5ZSKYaPwD
84p4i7jf1hPUw43OKes34fF3aMibc7c2pmnu0NQ0EzpzWtCiGZjyG72/pPaL90QE
gXdEHBYM/eKF172+l48mA6T9LqAZaymbdM0oB2HiOROR8T5NPbDLx1LTETRCGZso
m++RNY1pzZsYtuAjU7J1YTpY3L2H5Z0EJ6KTML8hApFSolyGH6Te/J9WQ9xhCbQU
vgt+pyrBJd7MAGmcUvqxsPxgRkCvJBszyP/tvoO8dDr16/RjQ0VH05VErU0ly8K9
wcSWta1hNspek1UsYh3zvQoZWzBEf99acrbVNM+q+5zaM5WKApV1FrFRVFq4TPFi
YntvJdhdTB/PpyNvLkrDVAkrNzkfLn1ComC1FXPJO+8Mnb7WdStlmmWB+OkJoJyV
jLfq3AIf9JuHgcxoFWeYktVBie9+5RPJkbkEa9DQk0KBWj/s7GzRJSmRjebG6gbZ
G2SF9lFFkngmOw0Rw+Y9NrlcfNLsmKpLXf1vFB9jtkup7u5Sk7U4VeZakeqCJ/6O
spZZVYsUhSwlLVIVPzy2N9ucmMbnQ0VByJl2P4WrwlfYwRV0N4nD78m8Xhgzt1Kp
3qiYTfQntAVIaJ2w4XziV7VyhyAYdnhB4HkXUeXV8QTZnnec7Zp+zuNwGgcXy995
H7Go59jopvUhucKsPkLCCIqOZgkPtL5xhaewpU+5sF6vw1pBMazW/a5OWVlvVQ4H
JyIzHIVTtYCgtRbafmMx3wmNCA5lVeeXq9Jn9iU4XbFO+SfujCK4htLssnfTVLxK
vC7RDA3mGX5FXreHKUYG4E+a1P/68VGRO56Q38tyJVS4QVtOiEGMOexNuCz7V2uI
xXEwT5qOKzT08GiKx/ZCF7jrRrJ2drPdJ9mDEOAmITncZQwEg8trKq3CoX7/pGGW
H+N/kuR5ED7qK4UpiiwxTckfHHvtEMc8VELwz9AWPa7vAT+GJcEvue2Sszuws7kA
mVGoj4QJFEa2vY7GtfSYU7MlX+gDW7Pq09dZ08QN2YcRZH+onim8BmQ4bE27NV4/
SzvWTNykN0tGiDg5bgaKs3oY+PtXfTKatCucuzD9oU7s601UeUtOuJtplT9HhOrP
aQ5mvmbSnPntXoMOuYhAHOiJXTV1I6d+xE4UQI8SF36wVgBtvf9/WXxKvm7D2xCy
74YaLRmaXod5h6Bp4g8Lg6pOodjZpfrIokS/9sD5hwfNKIDGCWCtbhD2jh5F+azi
QdZJ5RuTDNtLxs1DaQVAVX39QbXC//9Fd2nvbl/F71vjmkMX99hiPLFo2CmtK6+9
7x8cSyw27gBso8B0986o55eKwjFivSggjXAIBi9jQ+yH3V/v8fmg2dR91ZLONkee
oc8PdYOwrHdV8/nvhcOTuW2a1PPKWHl4R8cBGEpOowvLBHrmAcwdj7nVBIXFdXXl
y9Y6E7wT8sfbmsgnsCnJvD4m3PioA/LEJHJvHRG3QUBJhqwiwbbOW4GiZRUw7MvS
mnuBxljhSBzQhGUL6E6RaIRX0hn3o2989ri6A1YvHWTa8tYM6aYwOWV0AvZ/f/gb
NKIO3m3fLM+hfykyamp9OaaFCyeAwnoh+oqbSbwzk968+Oe6N93Fir/VIobtrsKZ
xVaq0w7UCTXoVN6EFhB9SxYqZfQy8OgUhV1VG7rnORgDLwPDrXacNZXXIqHG8jmA
9pV6ikx+MCJCobHJsLwGRspfVIy3dtfTm3EKk35ka0EeRDONHx4sCUY9kFkrDNXN
wzWqTZ4WkpZUOBohmyN0vv78jAuXDc32/ckuh5tlY0K4QQy2zZcnwHDvK7tEYplc
MX/tIlY2FO4NekrWPA8gMp7Vfiv4XiPJn/Kk1neRXmb5k5NQqf8CCCy8aghb+tlD
tcdYiaKs/XDRLGuBPcj6bZD9RTxcaNVl4RVfAjWuxiHWo+Xpo940FkZH20Oalu77
WoYp6bYipbozAl5ZAhdiLxTrcfM/6hdQ5JHXHlX7EinTSISd1U3p4+KfIyOkndhl
1xIc1mQNnKWcuVuCQXr2OVzMnS2gDnvsu8QLELnLEW5pYcfGrEl0yyAb/YMeaUq0
ustJSxF2O4Z0BJjELDVJhApbfTGgqzYjtQ5zljRh/yUG4GwzYoQf1ZIZbqWZQWfN
obQ1Z5gioj1btIJn1m6ATobc8QceQHzNPyBGYc2jf7QCKCgLgd6vz2De9FZBH0Cd
HqsSxUWSxQo+amufcN4ozZ1vEPZkpkYXPbg1pfMTSrAglbGR99h2r+yxgWeJKZvF
8ovcLIrBAdB3d8TTdRxLJvSehXc/2Dyv/2UwmpaxdR3u6Ezr7O+Oz96iwWhV67rg
lc2hq2Mk0atSuF8YY1vQiD/q9+x+EJhESnemd3B2MThA5Rm5xZGPG0KH0AOa2FuF
3JE9/IDs98I/16JVebK3RON64LWWq3VwEfHF4gl6AcGvP5JTseSw6jY+Y9eEW/m6
2/g78czAsAUWDx2NIlVmWYlDfzFXuMMc3ImzMys9bz9VwMClomzIKP1/iZ5/7d9l
KQcAXRvTfDeTgz/FFLYUkdKaquF+jiqjGkN6VQQSBmcpi3e/zSIlMpcTNnvam897
Rrxiv69Bp/UcD7U1ow+D8sf/fz9Ab3KIJ7qvtXW1V1Pov6YQqECoS70kbRHHp+rz
zR4vdthwdW1XY9kKnhhnXJj0n2GTvwnbGF3+DeDrCKjOT2mqn+TF0MAEPRei2DVm
fg/wsMuSXGEewqqGvlUZZ0nRyHGXQxrXggbMOAWJd+Y/XWs4w7URi4jdsQ+slaeX
i+rETEeiPaO6LHgp8s8TwaaouF4tIBrUb7Fh0gvF1uojDeYYeSqDKnrb9IYPAIFi
gaUH3/wDl5uiBsitkLS+54sry88ylRYEV0HnR+NaqVvLlUvfN8+nDZmzY9MKBsa4
F6YQ0zoiZFDLJuUtwWSCdwRXtw2acN0ULvzRpG/Z6F4fvdgDm3Q8egNuQVoIgFzQ
sDx6HPJGORd45TkuCcVWLGaZMnYpK6FCXpu2m91aruy0PK+omSMZtpN9Au1UZu72
APqMslhU2hj/RDc4qKBHtD5oGyW0QnTvFkFvkeVL4EYTMjGs2m6MS0IwuhL/xegR
6uKNIvvcJtE224zw2eKeKqXaoRquAm+VTlCdyLvQ0FxVfF/GUR2ixXo+Wm5ze9Oe
nbi9LzhP9sZFUAhviQnCahdQvJJ69GVcyDrpGtOnk3fXTYyNiw7tCEbTgOzfzVC8
hyAZwePIFtXqEiAN7glBa+gRjX8+1HrF5oXpa6HTJypQYueu6BS5Do+Rv7Tes5e9
GTtBFYThzO+0DoJhqBJYvVKZaBOsoP4tOTprpKFRnkXgO3PutTi9nuzMQ8GHRSi6
dVAWxjczV/bEoPJejDBYOx+mQ9P3eLepilnyzipHjYAUcheaPzM6c7nS5R46A4PL
ZykSLF0zJ7u1mebcFDM0LKqAK4DGWqpFAeOLwhL/0VPdMyNr1OjXYUx2UY1qOByx
N5LYRx9/SGvIgki6pEOwTGEcWZ1ZiANG0yRlgwaxXtvVSK9Q/8rTJ3eToJ/Yt/rm
3bWTmCgQq0wdiELmG76ZbDhIaJPHjQxNTWL2YVNYqN9gl7mbrk363wRqebNRuw2f
h2wAw7bUuJqUqoyDfMxWPMtqapebije6EtRsh/qzxP4tnxgwuEGnpWoZBj2kq72H
k81/S4RqJJrKD39hq3DLrwhPH/TbmRpjm7rz71zurj6x+jlK4ak/k9PB3ZFJ/fo3
KGAZ0/zRfUhAczozr1kTVsvI9M4lT4QVHmm9Ud50Pm3l/rCIkcLdfboGVFPA/7M1
J5DrX4qGlgPGESxKKPzqdIO+5M1GaG0wIiwnb8W6sQNfoZOFP+yNYEZAjbsEmudV
OyAvsUDya7i+ceGwP/4r6CzNjf9tznqL4ZIl3IvwtKBOdxmnFhWgZs4CBN+fccu0
3IUVffnHSvsV8oqR1TKhAhVPAw5K0ThsiBM05OTWCU3ImLZgDDaWmpznfUuPISYq
/FPFqAx5A+yp65x9QrOZ1BzXbpG05aUUHqMVENEJZjH/JV3gr+O96Gpc1KbMcnRF
9pwZA9n4NYmik0N8PvH9Us+YnXN3NHwZ9XFehOnKKiPhVExDDocZg6kPGsg/lgBN
nfYAeEZXpSrUR7PWXOSKKvJkATkxaey5Ww4mYNjjACL/LeFOj7IBZA7MoCZFoZkm
ubE2vRFdOAcvGZ0lvtHJ57upsG976zKxA3TCvVNpZdsE7hZMS2RJ80voeFExKkM0
DcyU4ohUzuPwZsvqVx8BcjRp/bE+5q4WBDFOgUiwG756Er4yss/xBqMewJf98Pc6
QwN081X43G8P9cK8RO3jnCCWQDozS8aSIBWhLRKGhbFQvgraIVbanpzbFhwr3CeC
5pazga1fwmNe6PrtaWOvUfR+Rcfx1IahG/fVgt93iCgA0Uz1vYbIrXEQhq5kj0Bn
`protect end_protected