`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20320 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
HdytKcppDjja7VfYQkCqvCGAQ64T8VPWTcWCKCzyUfMNjktbC/3EutwfYD5goeRp
K21w/RCO6zvHCId0v8sxFIvPHxbCTvIb7WFMi/92b44kbX6byKwM7V6y0RngllLD
d31+v3rjAxdo2qC/Tv122oKaZ53FaCfjQpvXkoKStX5ZUxzGOzL4hBS0VtkSpKOu
1WBOU99fo84f+iV1awdoy1tc9ZiB7VsflhE+iKLYz2zriUKiRv+1/p0s52C94AzC
iZoUqfOBkXhPklo0tbvCUFwVtp8bo83v9aqoM/bOlQLS6OTvZFSu4LspYpcO0N4Y
4RxIUv5cM+VGYUWeg7hfkYa5dsf6ZTTU50M1gbuAJUIVDbB/uPv25Og6Qix3Nn8y
V0aWgJloNs9Q/3LiTo2HGxSV5SwZ1+ilopIG+gbsRdzKOaI1MKsFDVCZLxlABO1P
SILeOnV+/hk7qir+Mv30dZDzYMIYaNRFsMZGO190m8Eg9oKIPONI1m3X3E/rpzJu
61Qx3qpj2PLYBtzaS4LVRESIOS3hnj0DBkydkjPp+VyoufPDeVUGGsG7jSoZr9IE
TQg4EeEkEqu6nkXdcZYGNQ4UjflqIRQcsJvXz80gz4E8/NaIgUuI74jM3cCW2+z8
JvA7INU19ILHFlin8CfUQjXPaV2x1ldmhpISKmtvwlfsNJipvWz8qGJuoZkJyEuh
LTPYNNJ98oKGCMiR16OQoxyMLoUaRTqc495pGwgt0qHRLOGVGbkKkKn7E4S2vmpd
c8StISojbPMVUElR7quqZqQPfb5PYqQFzz6cmJOATUgzCSmj6XqcFnt7pxUwxP5M
mDAJCtaHpygR8T/Hle0zyAVidMjJHUVncn9sA/H5F+y0kXkftR8Ax4PxqcVo+S6/
jsI+2XW4N5G+GtpQEVCmYjfsmeLo+TxJTus6Yj70Qmcj1W+ddLJnpSAUmT0P1X16
VLq7YFD8GPZyaZl8E8tx/DhFNm6CpAkaTX+Qhz2LFsTzweJ+3ECElxsyuvebSmG0
KoNzfPkCgljAq/hFdSwqW1bznuowdynWgQx13PS+JJdQccQiE4VlqSUoxj0sf2yw
W0eVzcEzoJ4lNfKx/cem99S2MR+LLOVahtxXwPcv8j5E5XiZHf2Ulpf6zgdEL2OY
clNMma7eJhpe2Es7yPlIVnBX6zb+XmNZWCWBmzmybzwILDhgXg68RtSUTnBOMvId
+lupIhyA6ppRzGPtsSiawIKt5ahABPblXKtqcrln4qritcI2R7ocYwBXqqhj6DnG
T+EO9WXHbFhP13kEmBxv7udOG9zfI9bxD557aHb21mDB92JwDJhBEI2klohiKXRw
DRnfyznXnDVo7Uzd35mj9EVG95vlhuOlZ+z8/dPqDSUvQlFT842CxvY66hsMzjX9
JnwZyFVfYlCa+N6FKZAwIRWE1vherjYlSu5yKJ9gBn1uYNSXOBStPP6l9KsanlOU
0CvHk1FEJoorQ8Quk3FVR6wGXzbswepfaTuGyYAjYFvQby/qxSbwFF8pBxDcvphh
fxHdtvWXg08SbD46ycoHjd5aO27QS4TgpbSYStK0te81QNhMuRyc+cl3Hmy859iQ
5KMTUYbidUV1XQLwtBgh+k4FQI5fiIqFFJeTxrBUx4gAcFXgnw46XLYmjJamyAdg
is+3J5YeOVydBfcWKkQjHSkvKCUKLJyIx9uT2PqoChfkXZcDL+qDFM/jzqoHj7em
3U1FeYqaN8wN011EX0/mDEOqzhSJeCyVCfOZy3iTbEdQnW6BoBnAMGohtOBtkbed
MR1xW/YmB8zj8O9XJ9Kr0NNsQjfyCyjW+/76WTwZqj2iwFamEWutzZ3fLTzvmzDM
twUqWN3HlOfTCKlfG0BGvn6xxhNo/1/aD/UoxNAU3YUHyoRfyJ4LR/MBhdcz1X/U
vosoetBm6Pd2lwpTm1c9AP7UJ9ZT03zq2eKEQbLYIWNOvXM58tIlOCX3yTlloFrC
xlnR8kJ2qmIK9SlAtoumfWqXOW4jkVJv+3d0BaUsZ4K7V9Sy3Ps9vPp3+YX0/07s
pqrTxX4SXhYvlSwLdt3AUmtHPSSOncINtfM58SSmVaAs2GnMjjAVWVyaVs1gZumd
80X51r3Am14hvUXRn9rhPkDUFSxVT9UpH65sbYUngHWkmVvJBcH5bGfD/PkdxhrM
B/u4khTPSWCHwzQ7CDEujR9ZXk+WhAelaWhGgX5rq2SZg+y4gN/0sY4cssjTyEt0
YN5s8Hv9mf3N79tair0TulXk4evhrIq7Hj3Fu6DNJlZr7W/Rk1+gkBDtPIgcBmLu
AykLngPPN8Vfy6rqOsJA6MWr5RFLkL6jrdVM1H+wJ7/ZgkvR8fmiJcGIBMZVgUrr
C3sJEnq8b1oekphxFm/sgaQD1rxqTzvDb58CYUMgrtDODd9hfhtWkYcjlDrmESQO
p2n1+j+fnWdNWtAyyvmMhw+hrjw9m/mwSUwkZco1qrWR6GHUUja00rwcstVscj9E
j7BB6RGI9iXSuUQgZ0rpwY3bnNJgYHJTbeeuarvmoh00ThLzsWsUrVeHjArajQhR
U+us2L4aFI1mOuolNwOVs6CudnZLfBqPYEPZq36y1wxsMq/Kl3zEKrEEJX0Wbw9Z
xduI699/GAXcFdG5j79XbsUt6Q7IQ0L9Og1D2q+7LFLLmT332lciP6juGOSshPCR
+P0iQUiC8qYdwjCPTI+SVGF+CkNg+ib2cyAMW/uYKrTDlphmqRF+j9UkkSynz13n
OTffyM+rg+p2uvSUr0UrLzVE6Bvo0AaMSPdu862CNKeLbJKJj5qZxeMBoCOLgcuO
16FtOzuDOLen/TAUhtHq345lTbh72kHmT+WS5UDPmK2fM9HkElU6h59PGogOLVif
27SznJyJPVYRVLEOvLgPTehFnH/l6ds6Qw6xVMkV8LLPkvR9eXwX4FMP2i4rjiqb
qZDxIamhni1ezQhvIwPhV7w//B04POoUTLlNR6lOhWIw+1NdxQOoAreIN8xlRBHT
d7Sb9NR1D72mNIA1w0ieHgJ3LTeIAiCF+Up8BmZH8VxSev6Bcnd180npuZFUS60x
oRaksIhPhW7dPNvvQRT5gufzo3i5vdcc7vD/k4nQK5whxSqVKZyWiUKxjr9JaMqj
kTXYEcryMJuoopXUROC6qgPjbniFksz8wNBODM6xyCFTfo1oMmWtLJ9JlObuKIsK
CbR6dSk5p7WLWp/QV36pKn2wQV0NqCV05xFsEYt1WgvAq+0XF3Aw8yx5SgRUPm3T
8YwcBHlThgbKOd36DcCNcXByJeCAscw6qsdo3XMpnRToo9aC7YNYlZsLCW4vGLCN
Eh2q9MN5XiXGFaxRnNxrqW0DeT2C6oC1YEcjVcs9oZJVH242kWrRmZ0EjDK55QXj
aJa2VpuDn2ChEvk5zhhDDj55/fRZ286nwx+/pmCLeylCRb83qrwpt2dVrW29Hju7
4Xxzh0M5/I2VqWNiBxd+0NPOe8oTh4EpLtwcrp4DSt+fOEVRYyuf0U+91jkZj3Qu
5+VWKX30qsg+bJwgp7vv49jkS4cUi/5iCQQ7+jxw+8D7JQYFYONsQQjxB8WlUhpR
WwfxmTDl0V6UfHk3jEl/RfFsTCRwU84tML1ibK1gKgQiVsv4kdkkh5mhHA4wAcIE
3WNK7cxeptZTTKACAogvhi8uBBeclXrZvaprNkNX0/mvHIySPdTyU/v7FGxEKToR
FHXfTpx+FwaCWs8NvJx6enLpDFgcg9vDOQ4bdW98rX4yQX7Ltf/eGjmXOieq5Dp+
hiC3YShW2z6AAg87Jb0hiPo8j/F020F9vT29i6NNrL623VUjCtRR1jqNn866FeOt
ngfsT0y4UQ69kGySD1in7SHXhOES1/a5MD6/XpZ85XtIFYee4yVdQYZzbfpxfi3L
E2/iza1NJbWn8dFL7xVrX7Rjdgh19F3/FTSDQ0kPAq7JYRY9et/izdSSV09WtvnT
7e/NMUv5wqRp66M6d9NlKU/stWkfvwgZ5FuqO+JHK05qcu398BCm5fMziKI8ZW02
VziJk4xol2EqWZE+w2oT5wV2hYhTZ/ViLUHPG4IPh366c8XLMOuf44RydlgqQfj1
K4vmWOhNj8eIUBux8z12KoCr+dGOr2tLQJOhQ/Yec4vJ6tZNAATVT/i8K2KXUwZe
RpukXt8GnYXcDWT0kvPLeAQeXkzEQFsW1WsjLBamjAajAN8GQogeF1YLboJPpShw
H3/L1eW92MCW2yIuygFo7vT52HqnN0eR6Ok7bDTURb+oS62WuCjpIAmTl7eeqWS7
6HGWNZj12jH+vs9RImQD2NCx2u2S0yolGcdkW1BRGwukg6p+JbPDQp50nz7BlI3/
tA3xOIN9Es5CqaTMjpJtBTgUezm8hqVtiwPCSmZxsNsiqCOpuWzVmIA8HNrUoSVm
mMjOTPjRAJPOIfUpAG7UUsEw7Fm7jXbaI3Vo894znJMrXb5tn42VtgYfjGi8hPov
NhEJuXpXEoG6zBO4x08hX/8YlevQus45otWyTuH5C7leOGAai4CnIXUqmQ/P1nwP
+azIxrbX8W4epaUg+enSDxUFDTcG/Lu8vDZgxNHQA+Is4wkcjI9q0k7AnJR0AJdQ
CYr77bLaPaemtkHGipk/+BrBma8Wo+m06zK+885+icI55wlgEQX++y1KQqA7VunS
VwjBSi5IDoe2VDXlch5H8Z+zNjJIHZSmm0QAwYEfkJy7HUXgW2r/osaiD1RtRKw8
greBGW7xQNIspGAe1f71xfQZj7nMdeCuMi16OWt7isFQ81SRMP6gX3S+QgDjz9CW
OS7OVBHtHKb/vf3+/80maPOR4mINS+nXX8EzFRDMGEon+shApMJNmxHSV0G42b0C
UZ2qdJoJYTZjpt4EhUg7z8OYq3oqKc6vIoOEMIjzrEB9eDu6m/eXLviJXT22Du0O
Q6sGup5hcjOELBRcCMJv/s76OcKKlCm9BLG+kftguyD7c1rbl67yv+NekLZMKVSo
YLu83+qArsmxvGiVUxYFMHg0LvWzpgxA+txxjIbR5nXvJ//3ec8gs88qDZxuzpgh
2yfnCaXbMozZrwibIJag4Dap5nLLPZ4Tq1tjcikIYSLbbAon3UKP1c3iji1je2sC
YlSqmlu/fSJlQFRAQFEZR27ELu26LoSkWF3Ybmg49ZQg2CCVoxjDXJGJBxGIB4Xt
InHVIsn2xOH3icHThhxperb8pyrTrbk4SGD62BKL0N94CwmkobTda+6MHWjaeCOX
gjQRmb4ellSpSn3QvvznA9OnA6Oc49jOJdlGyVZTQn9S36p8CiKeQJcLTfcxyLmB
3pVo177yUruV0Ua1JKUKx6QkQHBQAvV3vBml9yyjCYzASzkGCs5+4nWa/yR1RZbB
ItZYAppnfXyXKOc5kGZUchZFY8mBC4o0DhjsW2pl/janlSRbgGuSJNeW32+DkVO7
Uxcx7fIP1EHS/ERKhQmMfBKDQ/IAGUv2hRuQD7K8LxxtOzMO1/+RrVSzZXyg5TDV
OX2F0HC+BKXQtttNUZhVpcKLUZE0ORrJTWKIC7JrJJlM4OwwaTTuXwpsYtiCyqqu
rAm5T5FPAXbNUiK3hDlTvQo5n09OW5vI/NC6UUmd9kfkqqEIY5tC2Kkht+w/jNni
xra8jxIrYbaWycNZ7roNJndZBWjJHVrenX8ocZ3zNa0Hxy14P+HcMgumUm0yEXXe
2wbkakEvdB8n9r2qqDVdUJWSMywj7mTlMju4RRlx/CNvLj9hnUrZDZbRhxK1UPmV
egEnnO9HhfJnkJDFG4ul2rzF3YPPFLaEPmJK29m1tOzshPOshQnGWg5COyPb7Dz2
eFfMP6GiB2Rf/CfPQS8QX56oPx9mE+SaMsq7gAFQZZ+GefId7OpyxkC3CaRZ1sd+
5e+KrJc0qLVBOwPTe3DhQ9tppI5/Tx7GDmKBruWM+xi5hDZXEfvvs1GjqXlm8lNF
QZ0a+j9+I84357j8pH7V3+fW9LBzvTczfT5xva8JqpeJb6rAeIP75hgNWJbwgsgw
Y7+7R9vRiXGEJtlsDQPG1fCMHXEb1zZkI5zQQ59bJmeVsuUaLFmzsNFCOI5DILla
pKleO0OhfOPRhjIEVXTLFOd3lD+Ba7N9CSntvSsNfC/v6w/0Ivo9Eon232XC68ON
L1PYJtn/V5C2lfoJXDqu/i0AuXv5E41c0FShp9JCs8+yi7rfHA9mAw130SzseChh
jBUwo/EXWLvrMDgNbpAlmVuPQBkHlJ0TL6uFfOsk1wBWqs4NAc34q7oHrD5flVFy
RIE6QFhyy1fO0e9alxkMzlSEchjP0VoSjZASV9s/74N0YTw4ML/diskFrzeYIx+j
tSHJrCXayrnnT2krLSD1aU7X7DdeS0nCixVIyhOpfIacBPzMtl4WF2UP6Uv/g6YL
CU1Z0jtjbnYTU7XnE3mA8TQNaRpERRwJXkNMJmut1NZMYAhRRb2FZJj2jqn+/m1w
OkzCOIZadkLFku7E7z1Nqc0il6SQjvIFp71WbPtKUDNKIlOXhxVvri8z5Ab0Yepf
ayZwEgpnlzPuEI0U0yFYbdDg4S2OGnaubBJVQkk9soQLB//tqZg/H11voWIUwz+k
mX89xyR0ezjLTyXra43/sS11RwPLZJ57pPCaDv5LYosyteI2cJtxBICVQjB/kule
GMqmzye2mZXwRZO3d2TVHVpJZUPaof10wBEUG9crn1MSPKTdmYU4Ug7yZM2geL3t
6jUDpyaZHlRIDvfdx6HHKBY2mfirsdfCAddVD0beEiMOBtLCf0jU/eQYg3AD+axq
LIxjtqyoVSuTgFMvltEfDH+/+093sHZ7OahwTS/ibPPzTYjDwAW2WB6MsA60ujcO
Y7jgzfcozbdxPJj5Zi0ZbL3VBSytgGMVzncXIrlmFz3avhPwUQT537l5JxQJxRre
ve5mkQaXiQKl2/euQwfc4wQUl+6qjNyFZIc/0HR3PtpUMLQ32aCUZeuyd1iBIxgG
yn0cehaI9BbJ8pU1euTYtnbft6ISGR7vUHnixKcGHTIatybcjhT17/96WaD+OFnY
S7/yGRbhjDl1JlChQRYJNuJ0xVrIH4mNFsVF7TP6+G+F8IX11DI8dgY07jDWdUxV
Qp0gwLc4K7MMvp85BnBBFU1cmCHWTAZax3nj/tUlxbRVJB1Y5IgnV4YCRt6m+Xj5
3mf3zvSFKc/Gus/VJrKgLO2mCwC6cpv+mlNCzzOpSARhVfKQ6O0tnC7+ZBcfsz4a
jF8NSGJ3ev0tlVc4lJ8+WjtnusIfiLa/QXrj9zWAt5ulJCeAXqpXT3SpzLcBbfvh
9gWbv20QfN/Nbj1DDPDxoPFrfWVNlOKFFF9gw4EwXqDJipHLsX5LpljtpdhA6/l+
2dUYWqb2zKrUYSrCRktEg/gczDWK32VeLeqjr54xOgT5/BUqbbwDVc2dLIQYL7tr
uJNNiuJQWc5LqMa1mb9k96zXbQjFuKmYSZ6m3+JmAZ/K8vgFp4QRGARrZmDCSo1p
1YTK8c2KwOQ94kc0yHRXWZBZsfQAAKmPxqaf08fsB3k4bg6+eRvUNWawrOzPPG9G
YSJhl83aPNd0nTmcjGTJqmW+JCM924YPo36aQuux2mrDIS1MUFtxR1rV1OrgkEAN
0/eOAdTJCklsiI/qrMc03Aar83BUXO4wYExY98yDn6Cc27LWH+HSh0BAZnYl5beA
qfCEh2LZEook6ZSiNNRDtR92eoVl6yISBm5hFnSZvlc6uOHSRw3vrhv04LPB8yiR
7/tstWEC0s4k09rZ+rF+N+jUCADIcHwpAag0Ilwr3LJzdLc9Fq/JbLcQ2sRAL9bB
jqNV7G66nB4aJ/Zxza80SvJOhvj8idh8RofpeTfJkZxvWRvoriPXzi+nnTieVNh5
pqODb1ah5wWmeoLcXT6fMJVduARV7+bAhpKu+KUX1rXq630LpNzGhKAt7qDgfoAh
BuvNmIopNyyoC3W4wItTjqROZzU5FETxG0MrlAxtf35tcQNV19pv9LbAGKsq5TQ7
HnYIXQ/ca7u1L4hwGbwa+1rZBRxsuOKZPJwBpgKenergc2+twl98k/LeGz43rJTJ
5kEFSlJc7yptSM8bz6sqYQlYtHRsCO9ZcgWH4pVJmwgFaQuprysHoA1Gz9fxtKmR
5VziWLUBDgg/liZdNqwszfj7V6tJfuR60C/AoU5QAxi68DbyiLAQawcttL8/HpR5
gk4EGh9Spj3ScdscE7R4aeaLsmWF54r4HTxgNgYLOkP12mkG9s/Zho0FoJps149F
lspgh1O67/DRIKyYZ4aZa56EmkoEul1kzyFEXO0aw7PWlNRliRZNGQY2KX24kdsM
tFmCblNWaSe7ISbT8naJZor82C68cqmxU1d4ZFv51CsUu7LFZVALpKZ3bFSgCav8
SQymViDIH/9J+GPH+10jkP2G1ztDlmGPt7gvgju2ywLc8HHGHQqOZAPPk0zNMjWP
Cwx3VppYXPKErltGQi01sQ6Wi6BYwcD9hRJ11gBecd2T//iShWrpGIcEUS6raeh3
fLUJON27ys8/DYvp7cbHFe/AW08T+G/A+XP3Nt9UJ7b+isej1JD8UFQPZwo2JAlm
sPd34oNh5Y/9yZi2h0jgQg0XjxQC98cuWfRPWhFogsS6KBlby44jnCv36HL4humW
0mPexyJqbHVyyUpDFwBGn6d4eTjI4xWuFx9lKrID95A0LstqINhT6Q0Q+mNsOmGH
UjwkBqohiuIEkiEuAix0tZzk8IVJP/+SamxfHuWOJy4+JfADg/etqTu9wIo4bNQJ
2Sq3igAhXIBiAPvC+jIrdjtMrpmEKvmZ1+KFBx76R/KDRTZZ1F800smQUUXwA1FN
XR3udKLCWSQ+afAMefbBiEDsoFbRburkhonvPbPsWZQ5Ac6QEZIvvzTIlydBmvi6
JEFrc/hhOg8snqNTHqU32J2vVoH+5z8PBBMZHTDRbPCAtIVnHz8P9ZB4aizc+UU0
9BZGb8hwI7yILSNFlWwhQPGgvJ3t+KfA8C/R/Xv+IyTL02+GELNjQYatsrBt82+v
befvyRKZhNpn0WTgGjKCT0D/OX7aS6F6IU5IzYboGS9yy1kg4gGBAr1iK0od/QZq
o2noFgvToamLqfV7JoKZfsm1I9TNiALCsTmOMl28n7b1Tznzmk9O5oC/m7WLEEfk
ebtvSoovfRxjzXo2Lsiq/5oiQdQPhVEkTWkbTBUHr9gdRJ0uDeHcvZzDZHXrI+vk
2rUTfuobdKj1lm+FnvXBqvOjJSPeYlrm0+Y3xT4suJ4sPaPQboHXbqgdTxuUogcM
rvF/u8ObKi0iG9A+smO7r1EmdDDCm8+adv7HXDq5qNSizKl+0ygqqc2sja5yz9O7
3/WnT8cP1AnsW+Y3lb2LqVhaveyJJuevE7oNwwULsvRR0SbohM2X9vkhuH3QNlzN
tn24S1PguqhGyUZd+cvS/kwNjiXZUoR8Keot+cCy1JLNjuDKR1/2DAr/GiSOHenJ
/n8pFGsCXjGDd7XYeUYLOiV263sBa+fNr7V5zB9gELefMJAqzalX3u4ZHsTta/n0
nUTQdaE3rt1LxUmxAdKez9SG9feuLEN9Ho4abAy4KczyeOA77q9MFl3yVwfIGdzP
l8hDV8MNbSVZoFv223Wn1WP51gfb/zbkp4ZIvf9YqP9jEHtddV/brkXsaY/7qjWm
xZuz6ONEB7RY4gCr11HushhvziLk/SKHOZXbWyz9+7SijzPuXdeGBZC3mphpulud
mUc7girqof24ui4S/rvUcSKSSB/qCQUBzJi0R0Moy/f/Fs7ghDbh/qHCMtD4twHs
UiwIRnVciGuirp0TNf3b6ezE4Sak1dyrP/xSfQGzX7pg+GbCIvg2dAd+KryXfNB1
nlLd5wS07AccjzoD5OdZmsXIvQRBhuVXqqP8MwxPaDHxGCYAxr/dLteGhkM+Sjxg
F7cbqTTSnt3OlGgURHkLKnXbyDuiF8Qf754diqQN76v0OXf2upCa1jo1TQDllffQ
vZXJsWY+IG3KA2S3Xq7+0aLFinghOTZCx/Isewmlgw+8L7fuCcQ/RAdhZCKVvKAr
JZ9Cciuda2R3nCyFXrc/Jl45M1bZsAIez6DPcq4eDvykUoJk3NbreQIwxlyDS6hv
L+IettP3SJ/2isn+mi86gJteubhclJnjQAW15ztuob+75dhp5IVQBIWAyO4c2yWe
FjwZ2MkhtdElpKkDMadKIkQi1Fa2CiL5V+vtEoYl/QI4ZlyLONrtqRSp/4k72UuC
C5fdNSIwuailWa7GiEDu/t0769TBUWpu2XVtSvl5kIOluDlocwyI7GluNixzmk/J
zn+GMQc9aXwwBmdQjZh/+uIOpTyN1rQCrSTrX1MM8vNPy65nVwJ76ZXQKxO2rkWb
Rn8u3phY7FY6mU+s3evRMfXv0D+biASNk/It3r97WPnHbiUCe7b5X0Wna5SVnR9x
09/lmJjcShqCCNssuhqJWLhUHQ5aKTz63Z7y7fJn1gkARliYxw8g9laReoTT1caD
GObEgdRgKXbn4j14igoTANQNdmoNfkJlFq4R4Nz97eOPQABpIgC7igzIHTBpNtk2
0kajH1k05Yw9YNCSpdAZ/fT2nJmuA5crrIecsGiPpBjbnDVQXm4mabFZAlw7a/8B
eNPA8y3lgON+5L3ZKOJOmvPKrCsXWbIG8qquZ8vOI/zSrFfKwoKo3pjaDuGbmSdP
RZDPRHm+3LoYtvWydqKYN/Pq21BpRYvfZtxByVM9517xR3kbDnG084eg1nZOB8gr
KHmQyNtlkY3Lt1dW8wHh4GpVjv1stzdWgrjZr6AinqnGfn5ID8/BbNDjaWaoaZwq
ttTUI9i+FdOpre+UMErt6Ty8n+YRU9urRTXpAyFRdtiZAXnH+Ywk7yYUPzrVtgp+
lYNqGtuySo+xMfQeb5MDu2Y1ITUt4kKi4cw/londhTUTWvm5aHM/JnfoYUJi0f2U
CuH5qSqIPrMpHnEAyQ0Ciw8/GD29wQXriNvmezc6D/5+qK3lawwvHUx8ky7dBn8M
DU9iCtVH7mOooQKAETftJ5JRnTWCshiXT1zhelHSw8yRUBmiG49U1Pyh30XokIAC
tRcw/auvSkOIoXEj9J6p8lDnCuMhLch2DQnLznWBgPm8qaKM0kQSTm6F64GPIYCD
hj7oJX87D4FDvxkkQCqSgDnLT1b0TGEtLOrDQNONXZmUYWPgTmFz66mjvV9TDIuu
fZ+kEz8XScOrwIQDm/BhGfCOT1g0jbU1NJ30WVgEFT7fMfDBA4JN/nTupelofT9j
aFtOb9miVvyO8NqJBhNiLBtaGKEMv0e/3ylJ/aVvcTcXC/m0pfzgJNlWJ2olNXkD
0buM7itSlE76Z/05+oikpeM+/uuHVNWQsCwXia5mwRowFhRhpYkNRF/RYASiYlgl
gAUkxmnRPjYI/fYGAlv8z0W1N1oqKzbunxh/h/Ul0Is/vuaTPzMPhSMZpgaOZNsD
iyrgRzlA+RUU26FP3bhJ4W+4W6RHThpdIFHMBvAR7OrCtPR01D3gCmcuHMtYun2A
McHAMwtuS1L/R/YeTGZuDS0Vh15CyibCEkx2wzqJWdc40tWi+fWdrfNpTTu8tQfB
9WT94DgZhHlGUcOZCKITai5x8iNAcG+oroV3G9yYq7kFc58d4JZ1qC3KzQ3cV9Ix
NrUs84A4S/gi0Xn54IjW6DM3CzVdzNDQlpY+AkxybtYKVxh8+TILNLoIUmTwxG94
ig5K5Czs437PyyDWVD9O2369dm1lsSrJ92xXk9lpgXvWIC2BWM2ZnAa1aCx+gwrf
Dfx+tncUtmjhP4ZDtIY62PdOWpHNyodvKaSnecEOpq3wXMLKgzNcREHSTYN1awvt
7z5lbVy7/yO7tXkvcY5Wt3QTH57w+QlemQCwMW7vrUE8C6Fv4tlsSvZuz/jTjZl7
AADMcTRaNFxfdiBGab65TttOsv3CZQmbR/uGDdJdSowMGLTEAqyNYLO9NDJLH6Tm
DamwxjsCV6gVHeXSZ7NLPUmoq0EG19hbUapDISsdFRp9jaq1B2E5/1/bn9NFq9S7
ooOEzEybXzsPAcSBUpQsjCoBJVTdoprWjFlsF7ndU/ocv3piyILjYH8OMpIjENQo
LDygD8L4lnfL6X4N60pcqEAcrDK345jhLPPo2ay6VmHCMVCLpyUbDEXrxTjg+4ba
0kI/Ni8Z5BrZypVcjiE7KKl8IUNvWz0Nug2a/kG895GNeFo7bZYxREnYINRBn2rk
UdqYOMROkUqp0L8n6z3rxm6EOCwqbOQP3Lr8tR/HouJayCOJcwDp5mBXBsSQS07R
uZYqcogQ+XxPSB3DU18laOwtpxU/EfHSByIMnGdqf1JONhOqntEF9b2IHhjUCyLf
+U/Cz7juIWJvyzBCgZTa9pKy7jbEYPg1Lqai7XuOHqwyC4TWeg3a20KvtCXlQOyx
ekhjTXd3+lY/b7ePRxN44cm9rHNwwpWJ2VFGIWiwCHcvQWvwPK4ugq64cQ1HjjNt
QvADBHYG/D1J3aW+J4cJjxtcgrBh7cUi2ns2WBxKhyFbfkCC1nmJ9OkyWRXdTv/f
+YecHNzkNlgsz4oVoZwcGI7Ft6mimnZvrC9JdmQbBKchhvIT5UW7AnR9xsumzyia
X/tTCzfu6M4ThCoISYh9XrJk+V9Caegab7H0JSBhdQ7XkeWtO3lEg721OzcrVu2X
GEnKHqimyLbiBkNI0KWwM9IrdKtBuo3ffWUb5KB6cxQJ0gDEbyCdmTGeBSaX7SCb
rh5+bRduXHQgnyxAbLxauEnVtTKPMQnPw72lIcoCPzMdmJKY9lp8A35LpDp1w1Ob
2j6+1aVlE+hQPxyIBJT3HCiqF7xnhSeydegihwWq2B3zzVkAlT3OAggF5sOueOh5
armDzD2F9m+CA4wJnEgIkVBVV55O0XvMqSHE/BB8HpBrnNlcvX5BodCsnYcCo7N3
meIeqTWWTPjzOExr+VnGNOqTs0OzJkV3pkJkOjU0nqL3jyf9tRBR6Kszsj+sV069
upTNcYy61bL7tg/aKPvHFziDv4Rm5TzE3gVC9YeOL7cNJz2XnyE8CKGK/gBBV1ht
VsBfbjGWh/SrE1PNBOwG9BFTukgFGuyI0PUUfKXvTsmBbrirZ00jcoAYPrQqfrLo
Ca/AVCi6TdZEJhFmEa02GMQL7TUH5TfiEQjN84mvSFQTK9sd/diX5dkjNZk81Za3
nrEChdf+vYLrq5LQMcIrCAvcDtrrxjvKXOebXED17mg9rvM+LL+bM5TSC1arANzx
RnYu0PQOz600Vc4OW/pHSNPZVpOENFQqfZnR6bdU2HVSSJnsTA9R/RJX49gT+F40
xquoBZvrbscjSeIWN1VA2xp9IY6l2AAT003eg0QnwgqVoIYhYoD1qmeaNKpZMd/T
jclW3ZwDKLqlwmrvlFJj9SwopNF15fB0xpdutjeOR+T1b/N7KavmyXYzI0YEziyv
cssHWHLH37sStgYEf6ph7u3k3F38BRaNefFi/di3fYq8ihfJl/0rBGh5sgnC87xa
1CoQaECfpKO071aWA6VXdfvPzDKihIr91wRH2TW9ygxyzs3qZP8mJJkGSC4cjxZk
bPU6y4wGyAgnfS8lpfZVj6dBINrtm+EQ1Z1QwHhRjPY6UMrpTIcgv1AcRoU3cBhe
5VF85gEioC7SEmhrY4YRNBsot4IrmGzsYhqxEtNd+b3EJlQ2GBN41ukEgxyUrF82
ZhsvNQSLMIZ9ugexgJ2LPHZjSHR5Bgj6GsLmHVZS0NzmZ3/M+4FRIvnWQBj+p5h/
n4AimtnpSUnDB0DkAC3e1YSkMyNXsYYXKTSWvKEFEXCgM6UngUOSYvG10WLK7mcQ
X/0ts3RATyr/jTZMBZVKYHg11O55V9cVFVV1n8t/S6KhCYe4JjAEjcHkO11ahFOf
x3wntrYHx+4C6qxWkFk6r5pq7HybAhhjxoFVhedvZO6D1VkRqzIlC1A6CqQ/qHG1
gfYBtYkrgEJoK/eHj9l7qVyzBVYj7fout/CPS4ZY6y6exDDhITwKG/4wf6eXXtcQ
QbseUzb7wntsZP6CzOT6/PcP2JJyaQ9F9hqHTBQweBSwZuz9Tyls/QDGRQ8nVpwI
BGU81TfFfFQmVCSwzHES53odj1HOL6LrIplqMycd1psjGQgKqC5GG600kL+i9DFz
XoY0KacF5gjT1nKrgj3SimmjicAhRDStydlf1ILgQXmniZxqiyacP8Lqka/be1oE
x6TrE+n4Vyq1XPA8P5zTb2OjqNOGbnv4E+RS9ZRYTdbU4XZgNlfoVvjEfQ13/e9r
emiYpdG708s4HapLBOE0vRDtUPwk2/HYpG5/MV7FjWAVuXOtkuec2g1Fj0qrAw6v
9sBG8xYGhx25ZmtAgwwqICXYduuztlr7NC9r1Pe+iPNpY/P6HymQG4zAuQ9SeoXg
j+iGBmpuccTML1W7duKK4vh2LXMiYeyqHuhcbm6WBVJObkoxAUFrBdyw4dbsg56Z
g9zZaE7COvtubzyL9YBqSjRQqS4WDfs2V9TSb1BwPTkclNG2xSO3eIAOw9/gSQYt
j/c1kzDFPBQHK/7BS9OYQqeMyt5Z7x3Mq4nXPpgpeXU7EjOsJ47mVIDS4GZ+ydis
ntQrlH1PlGXyspvt14v2LvBsquAeUqOb//eRasCS0dRUQai3y1Z43Nac0dcgo1wD
NGFfHfO42p8PVqYjrlOfeDhdSOLWBixbRblYSWmEyT2DjYeKLvqo/xB7FsWUsqCL
KsCYQZvgb7rlCBas1KxIPP8DgA/SB02KCQukcWF+klaG+VRi9g7V5JJnKr7nm/FX
YSaKs0Mj2f4rBNq8SDm+4SzGZfwUgwF+fqzu7o8quvO+19789TZk0EnNg1Edmin2
BsOzENDM0TCrwkesmcTVe2/B/m5B6Ui+cimRthiAzjB2g5wmkS/+JaZEj7A/jEeC
1CEuRV8iBXOkmvPVGdVw7k9CeNmGlg72YIbt/6ZXMPyE4HXTW5SBBulsBiTAXiaE
pLdF3GixFXgI5oULJbGP1yZfXtiIN5xb0hpJr+Zl0fGmIP9uiwy5ABvduxN9K3jJ
JBEmpZNTCFe/uOU5Sh7Is5+wUMhrj5JtIsvd+YmVDmbgN1i37Lbiti6TapHy4H5M
EM8SzuZqjPCts5TwAlaR3i5jZ8VLqpUl/hue0JBTQxjvbH2QizCZ+LhYyfz0Au4D
ddtTtm9Hz8R/Q1nW5BMp2Qk5y7e7EMIy6DkknpqeIAjJ1Ep/LCZmDwGBMG5rxMEN
DSbJ94s+CNW18Hvk22grsY8JfFY7bhQm9P4WreluRTDuX1u4X2e0CuTjJF8HdnQT
fqBNKM+TQUWFx1PMjN5HoVK18JInK6XU4hNnn+3tLXNwMJYtQ3if90svbxYhCpas
NFQU6PmWTIuTYOQPZYX6+EiNRlEF+/h/i7ddLzBfzC4f9ABWGLvY6ShY7tHrV4qm
VrPHYXIESJUnBkDshbBcjFGWVyw5/iXQlZr0Xz88BCYHP+YdOROJS708gsrdXb+v
lePeeYWnsQdqtxfk4+sRLoeDUz7ABpTpIpPDo0M7bxBUgG6XxKkwMBaUx21v9v/s
JxBOS4f4EBvPkxonzQqpqaWIJVOXA/IMlQszWsEPO7wkzU7apYBUqjlNwmdyNolq
C/pYzS2mpf1Ez1LPpVwr2aS/YKVmtY4uquRjx+xEDPEP499v0Cmj+UEZEboMgZgi
KNrm2ugo/VcDAEHhIGDimaRv3IUFNyGfW9Y37tFfdM/y6mJqkRuw0LZCluwkRogH
zrFZlwCmq7o1tu1zHjltT/ZqAzJGMsvOUQT3roHUOfLSgQrobjsezwKwxDfPLikn
YZQffj4bFLcUcFQ5W0mNKN5cDajobZSHnRrJq/3uJMFsGrV2z4AGAYkGtDwwD2LG
+hSwvah24iOjOu9e1p2VC9AFfv4YgF4VKwDZ6B1uCqUIaOL27ncK2U0PDDvUQL74
pmTYOru7pnS/jO047xxt9s8wsjamZomShdIyLXmTokq38aNQIAVlX/uD8v1AUt1d
Zfe/vMgxlrpVoUoGjL687RVrr8WPr5L/zocrzuXu+hwpi+K0a28a8GczE9lYHKa4
2ze9vMXgLSceC5V7fIvEWwgP8hZMCIvwWk9Sr5cDjS9Q+EblASahTSPSo6L5uEmW
bKqH/DTBfZgPj/XEMRqJ5qCk+uNfJ8vVdT4wl+zkCZgb9UPBGD9Dav/rL+Mjq2bo
PSntgpY6pEidO/Ki9PZgh0GiIaprglsB7iOEPjyUU1E6ZWFzcoMTHLep0Z4vY7w5
Y6YkXHMiLolN5uo+sNCuPzu+G2VzO5f9SB0RL7kx0+pGmZh4ctP/xX/tAlpXCOCe
Q3WAhQFjzTHu/JFmzwkYef1UVn6lWiCmyIh8qLrOOU9MtvRPAzxa0p6uz4eBah1i
t/X8/oo6B7iEftdTa0SY5JItmSyjchLmZpHMryZqD8DVR0LSRSR+fRFgSK3csof/
/6LzL20imPD/B3CzZ2kVt2SFrZiY23oWs19E4EJJRFG6bxADTlHS3meIdWFz++1n
DoMXzSYaXDBY2ood+oSSZAEZWFzjkIO1f2WxHNlzczXmR5aeIAwbi7+PY0cre3W/
VYFhgxUZ1U7sjkzB9kfyb1VPB3UXhX7X85mdZGkmwU+qA8DGAkzEznzmhvzr2/yG
8m0wffQ4GSgRXUMd99CHot8MSQsK+AZl221qYvFYivzWHlyZJPWY7pQR5MJifu+j
CtTbM8PriseYGrR0Piv7wCvhjUaGiTGMasxYKW3hc9gGsG/xIGYCakY0QvBnoTcr
gnQ6jBXeuIJyGP1KjrXFOASRhV7HrJqaBL7U4LEKC0JXXzlROMpL55VLHlp/lAsx
FX2ZjEJPvBjfeTQPG/XQ9DoKclH1j3hTUupmXgWcb/v2TO8b54Y5uCqht+3BJo6A
HSQP0bm9C/Mj79b/p1asgKleSS9p+MEz8jnxnQdUL49uOytQ1xW22qXXQeImR9FL
tPY4IHRzoEcCwrjZ0+GG9vcH3jVFpPPL/G3YYR7XW5/I/Ykelacxu/So/+EJRQU4
7N3q9BVlLWF4zcW5fBw/Nx6tNpDSrUQU0dO64RGsU/LQQEjq0uXczINmSR8qxDQF
VFNOgdmT7mHz+nB3vP4RSwQNlo/bmRz+E41feHGnpskMUIuO3O9Rv/MPp6IK2vVG
jkDI7HwwyoW+DMYoNgDMAfqOgwDrhny5Nj2hwQ7UToU4zooUDsXTarN1z7HVL0Wk
asT8kgnFoeARosBmd8W0XjNkX4MxgEmUK9U0eCjSIAY7pYJqKlK3TpBGWLhjQ23s
VrVm8v10vZfErzYU4YOUWJV8jGhkLE2AuBDZbxDnelK7xwdDm3C33Z4CZAUP4vpk
ImyqbBdRpIhnEdojbC6I5XaZ9u+khSPY3GyDmCykunfdBCBXupb4/01CahdUG/4d
jG9dg/zFvSSGJqizmPDf9E+qPPXNSeJ5DdQuPTs9QdVnULLPPo9b+PadeLGA/QlA
aANnHa6GcKiOzHH0v2+pFAhe6thBeczLe0LmUQffxvBFUxDv+Di073SLSQMFq/hT
IhYeNriHUq/2vNtTOs1rBR5ZUJ9W/G9JF9uybrgx1S9ZqN2k/7PL7wMN13yj3ZSW
DMLo1+DpQWr0oXt0hngVA1UDzblhFfP4iupBHMSprmXXHjMfRT7ZrONdLCAqhg8Q
FgTNeuC8HR2Ve8xdMUZUGLLAaxUf8vt43waP4dCYLWdTAJRFbIQTp20WZ3Phbrrp
HhCSD5iw52iqDn0dru9WJAXgIPQNh93AcL3voU1suTfvG70P93IhCHVPPZS69IZD
qnkIneEF3CYJvmncu1EhcisLFfZOdtO84IPaBpSsp9sdN+0yGdR5eQd/BRbaY6Gw
GR5qMQXQsj6Rj6JOU7DWL5rpOFDjq5DofRWge+hKc6U0D1UWPs9Z3gmG7pjfRYmH
3OwwzXqoZeFoz28efTDfDzybHZbxYjZeJ8uLOa17c8sTCvf5HUDdDbDXBBa/nrlx
uwZ1Q76gIl3b1yGxqHZUhgoz39yiJoaOIC/CgV9ZBsL/B/F6mqTS7wnsihq6GLAQ
ns3uJtITc2cryABUaG2FtQRwukzcQvVhZg8+g3Wn5D8bFJDoAZP2FktGuhuNad4b
wRHwtVNdz49VlQUr9m5qtgUg/gcn2Ufm1KmcjoL7x1MWOipdzIYldG9J35z2/SSf
M50hJkPv9llR/9y7H+QCcOZtxcfM4YzndUr/egoZv8LvVs76id8A4/hl/3IKJtzd
AesmAna+Ba/GJQ8w/oLKed15ffa47Qe45G+Fn/GVf7O0iq9P8QdzcKo+O20tM/x3
VQCaAGJ2vX05qzPviE+8F6VzK+16ZBWG2bQTJGpb7+VQKQhsNDDNPsz5oYbc+zXz
v11FPtZloVeP9zo7qY6NWdD2t6Y31OKhcg+8aNIblwYReHbINl9WPV71P4PblGKy
FmYylrZipZAoZi8/zyqFf32w1pZk8kX4Gliag4zZMipjEid1vAkPe4NL4k6LAwcz
e2oX+qB4/pIdWGHBQU2gblqumijqZzBGwvHuuczwZaDGbyxl3qoaUBynq2rGzOFX
g2EQQ1V5nhRF2Z+1/3t/NJhNdwaqDUh/trc3ishqb+8vFcWlGLA5z+DqWGSJJd0X
jrju7sHjNBNhACGd54w7hc2HyKwAEvKFV47gqVNYtp+ETWkA7wm2cnMGWveIYCyl
p0t9k5Wruug2/FkBcyUwHBJJK9r5cZFZzDnmGHtUN+Ws6/QGLlowN2Rl/FT5vu5P
GjRIBL2CKfrvXEfVGggAMvEvdtAF1XFDZ0x84NaiiTvMXz7K+acR3DWsc6q1TCjo
XiDi8U5o8EL3Rannpd2+jnNEDHn9lysD2EE3q9jWRnzTWVBvgoo4HkglpeNtDrkY
X9ZLE8/D8bWBjUyhFrYi9MCSDRezwkMysjaKf7Hp2D878dReSX9Ha55CMo0anC7E
BdqW3R4//SNBqDXHb+oD2fXFCAaBvAcuWhzWyRjSG/B8XnnVBsVQHwrGNGgj860f
ehdDxZHsVHb5ZdanZh8NcyCkdS6cULWjSjPpNg6n7nct9R3Vxc/JuF+rne8MGpEm
JMso/woN7b5qkp1c0YkWX482TstV/KFQcOsuUEZ9/hKq6GnvKA1ojUV5D0wNcYqa
3lVpcxeEtCZ7Shk4YbHnLlmcFtg1OSgFMfy4QGXnwgQI6C4yxMpwUU8q4SMfEfbG
z0E0a/a3QNeXzMdhIQGQwu3cjX76mIpKWsNyQl5Oc8YlpKNfytkfm2RCuv1lzeEj
zxjfcORX4AitTWf9PXek/QN9hfwIuT6C1AaUeh3YxIKxAmTvciaGSpAfiMnwGbeK
lrIDN56OE/o8dmXwUWt8pdjkEeRTLJmdRwf+2qgoB9krIyo19hIkigRbgZ0rOMud
sW8MOh9pajAN1w6rQM/M22sVMx2HkffLFxiWH0QxS/TFsA9yiiyPr+/cJ1fmFKid
evDvfuM9SOvg2ivjKo3kZgEXeoYKDlsKrt2g90E5ra8QlPz5MtJtWKfBOjF1ve4E
iWOwtklgWTCRcdQWYxZSvDWkJqPS4LoRtbLH2eRGrq2YkrfamM3aAN+7GdCG1Dmh
wGsB9evJb7y/XfjQZwWtR5Bas/irC0VAcvXL/a/auDp2n47fWaTIada8hpIJBHnl
vJA2qDiVi1fBi4KhASVSSMo0Et2rhBRshKoodxxKXOOKpQH97IRXOMVjdyTlVXYB
tFoelqMXZrXvuOygQ7SJ1q2eNjxvyXJMwrrpsa8A52z8UYrOFQ361fuea2T20uuk
Jntr0bwTYJCquNcgAjmEWXUrBEV2ICgMaIHE4NaH3nJG8buVmqrgBbh4sFEyrlLD
QboL5iSz+vyo0CKmx3l53Nt1B9jdgU6Zq93r9oH2N3eDAxcGn5uyL1TYGzY6LZjW
Da/7rdQHM3n+R/eNZAok/Fd9dF1oRigKvOmMYHjyJ8D34dCr89Tqqle8KXDhb0F8
KoSDuOLoQUWFvK/FBsWulpIqw5wLMcD4uUmSFJZjOpAWMmhdbniwE+Tjsg4SXi2N
6Shc8icgYg167iZh/u5YQA+IAseAn7xj+CHwjwPatl7VN/Be6h8q6oRJtcySwIns
Zik2ndn4x8f8YufsOZKKud3kNPxzVV3QB1fE6cXOkkD04HDe4XE/zb7Y/4CV18kI
wpWhLAnDnDksT+IMJCZIA+twYA7Yk+h6z6XaCP35cyNvpgaFG2Bucw7M4oLHYROU
63Cdpl+axdp9hZH3AS3nfXcyTLWTb16REOYMk6RHuJwpiBs2/31BW022j3J+XkhY
p5vVlLQZx1Ra3K0ZBCWfK1NXuNIGYGzmXkBRomXPdQHHR9AUGDwd6e4QMdb7IxpJ
QmUC/q0+qigy0orKveX1TNyxcxhQMzBXCibT/xOLB2yclsI57FIaDjuZQgKycWcX
u2RZF8wPQOUkw7N3t1OSqx0mKryeHhQD8eiLmMp/ZMuKWJK8I9CW2xMm1ftn2M8x
yIKd3pw6gpt5ZEGFAxcP231juHVa6Ap78F+lk2a8FCGSZlelvIG6sjCeuEEaTeg3
o4aNCes7mqxcHajWZviseOmWiHmLw4avgbQi6xnH95YGBXBu6j9weyGat7zhNEf+
tXBbYW1YWl/CTklAMRC4qYw01iqAIvZm7ws6wwd+jB6KkUKmqqU5fTGZnifeq4YM
49dPZJgP+LjX3voC5srmxwdy3/cNbq4hv98AY5R07FO5yz/85r8FcvEJL5lXWtSR
TAb+GbLQiK3HqrwU3FFWDP2AsEnRkf4LbXZNRCOu1KmxhTfwH+NIvdJFxvhRFLyZ
J3oCF5YLm634lI0kutahQ3cnIhQ70l+F0imAa04wWifLWZB5P7FgJn4KSY+9Xg1m
aLZxzE5cHQ7gZSpIcSvn446H2R5nl5MAczEhz9gUlGU+5egDIjFA3cp2MU1p1TAC
GrrOcLSk6eahiMszGSgL9JoDffA5WyXeBwfiOck0dT+rZIvLn35VKuuSx6JzNTgY
yrxhyzjult0MTTohxJXrXesHXaKap281U64dfCNMLsWcM9lG2YSdLimJbxEg0QQL
h+ckoS6LPAeGptDi0YVgzhGB/ZOlwRRuQAKOg6FagnJP0Czn/Ba0MgjOOsHq1pYx
/wXaenMp34ftUWRCXREN+ddzfcAZkqeHFez1wnFu6tgyAb+T1ROkbCL8LkdgeB3a
XGaditTYkXQQnd+PZxoCDipm17j/clRqVf6r/jnuLzgPPGfQrR3otS71LRHTZ0uQ
j7qNfgU144Yd1M5gw+b/Lh+PHeI0HRpGwg6Yv/yeS4RFrJRdTB4x+2EvQsw/Jv7B
ITuU2cUcVktb70qAIZLHH0DR7aG/3BM6rhhrJBCNOVd+xPvNpIUzSEy0Uvfu9IpJ
jHjM3FRmwPHT6Vs+4DJ++HlW/n0dfhj8wcoNAYLbWBThqi669dFKsb9VnMTwBTRm
uh3T4IsdphPUSTr19z7t3UMo9dpVoeXUcb2QCjVk86NweyacwPF2dI41iELYOTSw
87hxqkMleHR5KaBBow4jZD2UIUnP0lg/QOVlpn1KUzkdpY0NLboiHC8Fez9DksrI
kebTR6SHUudkgfopQXt0TCDtRs/DKE6l4KKJKZCCSWwZDFfBcnKWvnXrlX+1SM+0
65x58prLxzK+G+oOclDFjfzjOKacHmtJKS/Dxu4ZEl2qM0FXtoQlQip8ghW/htLT
sWIIb5yd0sfoUOlPDbIJTtqDM4xP1JFIu1CICosoZuIyUlSx53WsARNW7aK9JjEs
3cxJZOT2UNCGFvXQ8ZgInO7ZXlcaCpJv7TxZjmu+ssmVrWjC0d/tAN0quInVTGya
Ivp4z1CMiQljcVhX61LD2xYAbRae88xkh1adKwKJR4cJqi4W12gOAdDqiLHg12qb
V18jeJk7T45lRxJ5qvPIHMcF5EwRPfRhtclmbOZUYT7Key7Pk8CUCs5CUhp/QcWt
VfCaOyYuc8fZeXJ1HrkRSyQD3DC35I6RkbakGvB4mYXrw4+FeSkTvuYZzAGUdYbb
e0KV7t7OwOJeOViuiyhW3RzK+n/yKCwMCxDoQt/I47Q6Fb2SDjrknPUHqLKs3Gi+
/7LN06e6jM+wjiZKKF9o5ScAuykmHcoTIVnWf63ZLtC/E5IDFjs3y6lGHvxZudLW
/bV6jrBRP8doUdCxabWzkHLyjeL5NBQaHxNJhbLCscrzn7++Q9PKUjNuXVxPZmrc
GBmhKD5NsivhbjMJSd67G6Hdd+yqGiQYxSzI5S/gz7fbVoOVxqsivH/cFX7cvg0v
1iVa9oxpLBcK0IhpmwySUsvz4Eox8qiCJOLXmvgQC7RWaQnIWsl02pqpAxy/tEmI
MQ3oeiwTaIpc9w6m5WUAE17f45RgXb3utNiZMrBxuYX7LZB1a/nV40qJq5DqwQzD
PpI2Cz0jycrzLeLaReZj85fT9B/1vLCIhkGEmwH6Utxfd0dPVrciXVjQFQNBKHh4
GqfMajIK4MjeiZIdTHTztOTmP3d1mvnNu9mAzIiHdZFMCx9ReYq/lO4Az4qy9jtt
PkYVS9C7kJNgd+obvwWOIWFsMiNave9gwQ6YuB+lMuyJxQyQdsW31k0vbRwKgfPK
soQq6f0+T46WCE/Od+hF7U7dhwpziFfLwOcTahQwXyiQNqYye39RwdGv5hOYB/Qp
UdBqEGMT79MgaXtjESivxBq1gRUJICLq6oIOEZIcte0i16omaP9EXKgi4G9MgkUr
oqp2INRLNxrRPaK/v+fSc1Cvmws/gRNMqijc3h63Xuth4P9aNlC2IA4UV1NqZfF/
fpmFnEHrgtOlIZ4Wu+H+AS5LlVHahyvxf81u4O93Jzg2AKSo4aCPQ1zyoSUu0vM0
ECDJ/U8M66D1svKp2WBZ7Fr9ArEHP1gNhxKFQwsHiLRLs0v2KpNe0G+tBRkaLSYN
Gp5VfW844cE8gK2Mj4OrqV8gRRSVg+Bnb12Epk5wZOv12miIn9M5h5f9vfzWyJlH
SMUiCFXM7AI/r6/jXCQ4pSVuTWdu+C9WxNTp/e/KPHqCCwe9IQg99C9PpaWPMGd1
X8Y5K6uxY41bsCEc2ZOBxSuIodvKFa6jnW7JD2ZCk/8pykKLCLGOpoiWkCyzg3/X
IsEXz3xgaOyIdDg0ztbfxPZzrSPrPayxMdik7fy4MUFViQJDPR/5Kycdxj/2OJMh
zou84ITbbb0FfjFKb19ORaezl+8y90KZSFigMY6CmAhXq59rR4kwz6A4weePmkqC
ZM0i1uukTIso+3eIPPvoqcmXo1BH3PEo9RPWJrdDRoS7tFIDQBVKrNFGB9MPUKnI
DNCfTOezWFV9nKnro5gPVF4jsL84pKknIhDUFjbeQxPJ18tBqd1oWfnywvFV6N16
w0wJCovMhrDY1QRRB+rsQMs+7KxY9Wy2viEqQgQHyqO0ZTVX3HOa8iaf2gts80Az
PmrZz/YD42FtsjEvOS4HX0FUf/cB9KSYLpX5mr6tQfZgexsNu5greuHOSbq57UJ2
X7AwMj7uUT7oGs1XigtVpaYsi4e4oxYfqCG1lDzMP4MFKh6PzQ0+6/TueJmUStwf
EFkhNS9TDepYwILj7/AAC3qTo6bLL8WiIP+8HGFbT5NMjCXTpPzZ/mtOl62uPOIX
CAUkx/SYmYUXQgRbUKdTHpEgiEOH3hfl7QduJ8PDJ8vx+Am1O2BRbO3+9S72oXt3
Zr+3U3FkkkwIGLSsy5QNRP30BN50ZS22TSR3CSYZXTITrimKaumjugRcVoWkOhfn
9v3NHpf8hsu8tTzMBc20TSVBvvw41i76I6cfa4e13T0sD1e9PRlG8rswHKBe7tx+
dMdKIGjridWEXJh7xZGMgcSYvYlKAHn7ckno8gjS0CCEmbE7/Tj8OyAAB+4fOn63
KVXuCLjbQC6ULTkBFUsLhaH8LbaLX8O0l6Mf+jmDTR4ougMXcyg44IoLmFhVHAL1
E7ptRvLbJWyA8hcOXqifqEzuXRrTS+QYTMzPxqi33Ju2qGeFmsByZMWuLarU4pFd
rswG72ckyKq8EZm18gmrU91PvsYiuG8ZQqxWN3kGr/Oo0CihXTB1on/xUmgZQXbA
F221ox+/s9WnHlGbM7y7x71Rxp/oVC7ViH/G41aDg2TjPRUUmKEEkIP8UytIO8Zf
F3DFUyp2JiQKzJTZpN46Tnt+Tv0qL7OOussKS1Tf3hzpsOqd2+qy3uLgGz0K9mDT
QX+ptzLU2gEQr1495IH7kLdWSdDA/9Pkcqe0Yk6mWPkH0WPkKHTS6Aar66QcOSFu
Yb/ObdEhKxX4yedVjM0pXHPsvAzA9cuwAhZFGzp5HOjrxiTd43C7xoJ/a7+LSbCN
WEF/edW3pM/dvpfLa78OODi4Xe2VsbQfoqpB/4/XQ7rXecfN/6rhPw6yQQ9e1ILz
PZFmRPHaQva38aWNpFPn3OnsiEiAWL48vymV3q8QuXayWcwNyrL7HqeZ0K/BbPxc
hKu4/yFtgFXFy2nMBAVjgdU207zwyKDAPNszE0RKM3xMwy3N3t66nZmjra9qvRDE
dppT1WSsTiv3/fsa3A7kO4KC8+xUrExuyCLZJ88O201oWFb8RI3QLckWv8boFYZ6
BkvrTjkNPJzyc8qh33wNcgndksd5vZ2juqlVnWipH42D2DnyZyEu+caAF8iSZRdF
625WWbWP9+4RPE07qPVCM+hvusiu9gV4GBJJ2H88gsMMWCzhkSykCN5QZhCet07R
BUbDIIdAcu3cOewoHNdvfeSZad56oXr7pAF0nMp+PMc6a7ojiTpmBsGfoBh4mPjy
SR4TpIki0Pm6jf/mGdtVRxxe3k30agqoajRPUSXAy2n+CxwYY1K40FgN2qjfB/ZY
k4QgCd5RtoYzsbNgQ+sM6J3WIxPvV/6fe7yDvjw94ZVzFl6jbiD/cWCMp27MwcNb
/2ZgGDtW2Qnk9tweboGhkczmBaivPnwJVWANLEzRwzFEGLTz5xud9AiDIxF7IRAU
H5r2bJVFSKZ+ksnOyC4M/IgO97Gk4tNhYew5wjN7SoSyJmPH/lmhpNRhJusaruOE
4rMl3YgXKZbL5NX65YTm/VcL0JINSukeoAiNjCi6xQB2KhZ9h6nAVDR6oDmu75Jd
FSimukmC5YXWqYXUxaXMpHPP73OR64VVAtdS3+U2cxzZvN1ityZTjAwlsLyglhZN
q6Tji2SfxklutbK4bJi2c0FzKNa9UXos+PLbrUHk4SqtCBmAnbSq+EQZBsd5Wg/o
WhPu5T19pTwpBJGVZnqxHpinxM0BoqRP/i+SNt2Wma5Si1nxjWXWIb6XeXIYjr2o
YNc8aZZRLDG4rPoleyry0HwwFiVRMqxFiFfdZaFhbAMY2ZlJjbaDiwYQvsl6xH0I
eELRaPR0bIW6JxMZ91l7N/6lYoP1eJzyBr+uyzFeq6KoPBuUEoHqRbENsdUC1iNG
tCGA9jdDzR3o06T4GFWFuHXYynEE+JLeDMb3PhYbvKJNUM1lh1FKbl62ia/0S06G
2So9l7XkdEfUMDeLVcirWAzvZxo84wo3j/OSQs1usAzaO2ig17Sca+xglxiIZmDH
GDSVScPdnU++dujexMldY5JM11REAXZwOdMgN9MfkUj4reDqWhaLHQmAqiB5e82j
3t7H+0CbdUg9E2b1uAcOaEwogZPRrVuEvR1Getod70kCwlUbrhmQh8kDUeFrxHgS
wme9rCd5uZhX7JBGVduOjhBoZMWn/1bKvUzV3L4suSLwtVrImfIlaZoCohXpG5LI
VZMfH03EGtDp3HFEIms7SnWqxxRuiK/kIb1djlHBuR6P8NpRWXr9M3hneeNXVfth
tF3j1L6gUm3HK6eOity22bOuG0KUYgHj2BzxPAtZh+OKkTAwMgGww2y3SiRpbM+l
uOquQNSo9d4wwKcnz2DGE/2k575AvpHdpshyB6Baxt2fiWN1UAUO5xDGXHsqxJ48
QblVcEyn5uyiBY6bmekYzl+aalWv1HDM8aM8yg83hWglVWU4rEFXsOmznMfhWpc6
/k0NTZJHnHjblJcrueKzruwbpe8k7v0pyaPbXynXJyiiG31cxWaAMbyovQXbJs4F
SPQuB2wzAXDJ9c4CRWrWC6CMZvRGqjGvTax4mkqU2La2CiAcmC0SgThKMxH6Uu1G
L3DXaigJbdBPZnqS+oby7KwmhTcDigTRIpCrnaiCooQvjZQ8KliOY4GeBaSUjPIJ
BG1Xbi13+TCb34GyNedPXxjkBLdMBOq/1mqENaN/hY4QzoflIoKo+H3/QfTg36Fk
83+qM+RILB16bVaMYNT0bPDuoDLeWubHXyMzbmqld3zuGo6Ow7gOhryENMn0JBhy
jo85u/3zjsrt92txjRiRBOqgXplmbebQwzG0hVsBeCj9Wnda3ArY6SopP3h6QxLX
RuHzTB6TLueN4YNV22HRmrfpZJmR+KMnBRdEOwKLa9HEFvrXXUuNTQvcFgIwTsc1
YH7elQI1Xc0/7Kfbqz5A3KZtQD9PpKtMMe9fgjqdRfji8i6JJviL9FC4efcl3UMV
t6SNGUVN006LP3Mscd3yWFj2ra+7FwiwB+bXcGe0no/FbYYgOjs2PZO61zYvzhbE
NTpjyS4ue9RWF/iklsEGd7YWX8nXilNgPUDCSSBs3ALbgNUxuiVSYqPuGxNG49pF
FqsqTXx4rJl3xOvC+l2iZXsj+kRPAVq8GYMOw/7/mMFb2q/G/4T/jLS/rpkKk612
w6ZrCyLGt+p7v7N4LRfVGA8me8N5hhsxA13eQ/ea+3gh80GVHIH6w3mFAgYY+uVh
6Plry1roWRsejbC2wlE2VTIwsEzhYC08u7Tks+5yc6mYn71acA59xhvloM4yXuVQ
UC++QAuOinmwWNbQBdEaiMp2XQHIxUaYuy+S7+cF+/GvL0KYufjeAVcCjBxgCzpN
FTggR8gqGissfiER7+Ai26Nv05XJNeID3A06gG/mr+85LQDGyNlIuGejKu5Fohn0
BZdOigOBK7KrR7o2tkjGsw==
`protect end_protected