`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11328 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhNy6VWIb/c231w6GZGaUgwhUZXi7j8zUEO1Z7E9J3zs+
n5pb+7+qRdKaLN9hjD4guFRFg+no5bkBYlHATkQA/fp24EelXluh8psnF6ekBxtx
Ek0yCIlq1rzLmlDK7vfgVl1YeExulRE5vh+T+KJ3vBHFx6XtfnsMGOVXokqffOKC
SHwkUSqitTjoV0x76ZsTau5yepw0CHH+MZZwSk+uYNcUhrbzK9S2k3Ju3m8NERRr
uFC2Qz8V3c0y2PaqkrNA+QU1qO6hhX/B4x7J+aBsZXG4avJVTG6fFx1Dx20MW85q
Wj6rUTUZvVzcS/ZfvPMnjjeBdnqRos6MuYIx4v4NrY/Lt73xqUIWXfElBfL18aa6
KdImwWv3wHiaU47/1tsM+/CZbu54iTuU2fZLqQVGdYWryHssDAz3U5RJwe6+NBew
SQiSrR7URD2hdmDTeWo8kGGYe7vtbg1eJCbX7+Muyjf2v2G01BKpp8Uzn+xsosvs
KgqSzm02ZOOQ2C6AgaiDt+4EeZY7JrJWrVjJN2kBplZJV+wv+eEJV5Eb6LEmXsMw
IwL1+IUB+I4+9+zHqMAzCnHReHV6uYUNlQX5FMjPxQm2QBmSCgmLdt9ay6CdlUj5
2a5rP/Rzy6BQsfpRgPwU27lFOMgwjGkebUkOZOuIAeAJtYtQDZEv2lGBPhBBowL9
kYQw1VvVrk+MKhOKsYz+QZLG8ik3gebxHgwk5e9PWBPTlT4Dw6hryvhoNde+iBlo
Y53KdRwtlZnQr+imwm4bwx1LST5CK2qejOzh/x98xNEgF7+ddGfbaZ0YbKro1SMA
3EMGKUruWsskYMMr6c2ZZjv+IH9OSe2fPVdPYfHm1yeX2hN4qn6DfJbHAXB7TDa7
/LQ2oEIk2ezfkoj2aHBJRme77UfMgnoRhSb+sCvh/1q6oucaO47H2BAbVHbzPOyI
egucxNsdxgSDSusEj+dVOmux1bhBKjrqZU0fs+lMavo2u0VHvj7yCeMu9VEdCVNG
gAlIICBRO8XsOmpR32S52+IOZMvnbkI3DX6yC+KgpL18byUz7SfzL8bD6d3TtiQh
4yK3P34PHDHxweY2cljnmGZFNUOcqQitcks744CjX+L6tr0yiDjU+RI+xLk5t7mW
gY93Tn8userPhztXlOPY/gzqXy/XkFEYbrSW7XAfigvHL3wgAIdcCXDTJ2cfyPgl
km9NNwxxtOwjSwyV4raM6ABce4eh5YTa9qHc4khnGMESKP9HujRDlztZLc3mR2kj
oiH/aAYhCWxxEmAPH7IO4/TuKDcFow9nqxLLvcPKsZ+WK+f2OXhesSyaq9ifenPl
+BU74AQh1JQMXYKDGvocdk2Lw/9BNsnlfwNO19qL6PP4kqn1SIaskTH3ht87qvGh
5GCM3EVfjhGl5xOxtSUcaOZPQe+kcO9m7QJpiwPoSp5NiGhCaFL8aq0P23DU12j/
A/EjA1JYvkSUWGN2rGf8Tdf304eTNIpX9dF78ANnOLgD3kOLEsHqquDT8/fOoXo0
Wd9rxHpD0D2qupURod21SzlRswgfNJBFbnj+nWIIvNt/ErMeELIcQNT3JExh1L3z
PmMtRwYXVAbJK23gTUaCqdPcEmzsxiOGwYE+MUa/pLUdU2QiTOc8AYSnApAhvWgY
lSiHS6sJflBdJdDgL6C8zru7QTbcHdRX7ofTtLx+GrZJ/9QvvnfgKraY0k+IRnLM
6WOwT4ioMx9nN8fEvBmqwuO1TlKy6jmicqEWZ1q7RcW8i4xlOBBQRbZcOSUQ2m6c
T0HQL77/f8duAaHOkdCrhago4/0RXEn22F146Z67XwdF2WuFUgOh7NRMm5fvyXdX
N/RwBL3Qlo/3hxdjgOoQh3UozXPyL1GwTQdytbTbwt6TkIt1IocuznFIYa174aoq
llapI/dJ2hfn1RaOq2qfrsc/Vpu+4P20HXgttFJg0wDicwnxlhKw1fedWYWAdR67
0OIFQ99U1UQnJTU36xkIYHdVivZv9DHz32ML72M7vp7mTLbTmnwI6bN7kWGalt8/
rTYafTIZBhPj1NOrwyAONjeBds3fqsPz4ynDa30sYSOoipga6CCR9zCCUgkczh1a
WKZfKHfnNlJmzPELXpycvObOh0B8FJE9U3/xF8meP1sgiM2rw20veOR+8vRv0IxC
0XT23N4r3QOhUPS8WYwreJAZnhR4OyXVnhzC75UZ/y5EQKAQXk+qfV6usNvTFQRP
2ANzHcKWjmMUITeYIOK5toekVxPUFuT/+KHGmszvVUigwS92tvNZlcTXNfxGVDH/
NjLYvcb//Q/0FpUiMxeAxqf3fJiRDitU7upJsyHWqjSCFLT9hOoc8q4xk9f2AeVr
rJEgA/xApylwZJLX783DuhRtMdbzhe3a11Zfi17QJu0dbYGyYsTx+2GwBoMl6sph
TxMagB+oWQCoOFqTqQIn/1aoWCPlnhwBmxXPKz3QdoDHiHlbIIXSYZCNsm4DjL/6
Xees/ToYVZ1JsvmVVR2yt9utS4rJFXoDjVhK3IRWpFJWiOagAIVLXjYWPfAwb/Ge
LGuSHBt5UzHane+WTCcKCl5KReitYwdCc+1VqUzPdTcjD2cBLJW4sGQLKSPGL4+6
Aphf+q4xWeqp7V2ZACDxEIeYgWqUWQTOxNrw11p5oVops0rsK/6xwRbeYRVoXu7H
wc3XA4kHHM7JwVqLdVf7/iZFKTQx02GGYwUWKHn9ibw9f3wJdzPqyPQdUBjvCJLD
QDXOe4r1nMuL6nmTAZ3oIJI+rU4/StboahD9H0YB5iqjqBu8PJPl+NZHCSMJmiHL
dnrQB5mXnOPCGOI0CGWpLJXJChzpOKHJT/tus0z9oVUvuWf1UcEhaLzXDmSlPq1z
bTul0Ju73Fizvk69ZqkK+R0D1QWa8GYo7KstlCo25yTZd17yliXu/ih0Lk6E2rJS
VXgl0nKE7IqU6Lx+G7PveAgeA5xtFRfCOBPnBFUkM5wLrSw6PP1kVuP1fNMc3pEt
iwU+YUWmlgA1QsZ8v0us2HHbmjGmGhIcuo8qndn+aI7Zpf9F5GnwRc7cZQ8hmd1J
aRlFES9jdrkGwZrzduVm+gGo8h1ICOg3vhn48UAk0Kv/n1Ts202badCjI0WAs1M5
6OEVcx1UWY2/5DJecpWEiWt81Z7T2A3wZPSdxnkXRs24uv7tNMTQikwNSu2ioj7o
uTmRoAtP3USRqsNbUKdbMVZJImU3LNMZ0qR/8pinuqUTPZGLJAh221sUizDnCPQl
pL80eBQcKrcU/by2DobmKmMwT46P9zEQMNKRRKxp6skm8c9CbVobDooQQr2K3uMu
JRDIdaubZXdjMzsVYUhxjg0GgHddH4IqJ/A6o9GJteVqUkYBOxjXNeP3+5DEpT8s
ZUBmVU3isoQPDS467xMl+bCbdW9U/FgMMWMmSU73ue8YqXmDT/OEk9yj891mrLTB
PcENmHNSFTU8pt/PRa8AeU4wpLNuiE9jFIA4m6l1fBx0S/r9mTm0tIyV75fbYJVv
F3mCcXpguuuhUjO5JMmr8NzhlShZdg1FnmvCiRRNnQo/CvfjpIuuUtADdZZB2xET
y1PTkih2ZW57ngbboPCmtxYsjhxMD0nbojAL39MUzY9h3gJgeS/f7z7tVx6mg4sh
ghowz2Y0qLHswARttblUbiGQz3Row95zu47mBYuufV8Q14qa1lOolLxiQlOEcP9G
/1LpCDv1oUGASy9yJaLt88Cvwn6gX5tWaStEvPbsBqQPONXeAP1vyOxPdkbuImKF
w08x9u1vaJSF/zbIlfSijyQty5SaIf3v1hr2c8C7hRwKqVmTHu0bfxoGPdVGfGG/
pnZHKvCh0geOuCfQrBA5AvTN16f6xm1ciRvAzbxnUjZuTWqD/AjvJhvK5wSKV3EU
x/TsYyiMMkMLpS7VTQeEo54oTuOCJS2cBVdfplNIQ3r2blQ07DuMkhgHb8QTlu/O
Hcef02mWGpLAdgkyGPzRty3a8D5GOYqO7+VcnKQwNkxWNEuhm0ba6vDhsSAlJYKX
qg3Z1FT1Ff+RNjXXc1WdpAifWPV/8fblnm1iE6ESBLBZKo1Q/OmAU7tYRaytUAns
eY9ottDXY+yspyJ89VPf0KvWpFVf1ffsZ2Cw8MPAYyXDWnGA58kQ5vM8M9jppL0X
vr1elfR3PmLb2O+nAu9qrjLu7dshFN9OeBkh4NJzX2+v2eTa/G1x4RPHVuB3pflk
mJH2CXe9ZJl2cdoLsrMvYg+c0nZ/uvZBi90Mz0aXP0p7hb80QiXCx3eKrAlmFhLi
IF5YI8oo7R+3t0cilm98+fCClm5Eyi10xlmh3pjl6Do4n2r6cVAHfEE4KiJeguX1
DSWUcwSSG1cxp4tIQ6C2ELn0YOawY3vlnV22h0mlTD4lFnuT7iZPWUn1v9qiwwcP
OJfI7j17gznH+1znMEs7NQRifIsrgFfypaqeZkgWR02WLsNrbbpcJOANoVihoJ80
NxN0ZXPKgflgHnnb6Jik1ALlt5en71Dw62qwgA4G5aC/EqvbSl3gKAAaSnCjwLg/
+4D0Yhb9ROOH8ujNo6ncTEyjDSWmn7gNSP8aa7gpzoxg87nXsImX8MgBZxWh+NF9
xN2BXYZTOoX4cBvuGiZinrNnOrXOpv+RkxqFV6vi7iu/qR5itAHArFhF+bQxydTJ
sedabSbLwbwho+Q3d7dWiUqknRJ3lZbgM78aHzwIUzOUPoarL8SoWldwbfWPaM/L
PDgTU3TFel9rfpA6iiqZhpzeDq/dDyyFKIiEtA7NYUsGwQhta8i7yyFzOpmSUDTR
IjiGvxakUlK9k23PMywR+eAUdVRdpR49wNL0WBs6K9GDmAdTIgrp81OpHKWxfNg+
9EIaflQRzYeYxHzeaWI7guW49T2CqBlsDImFM2XquXNBO7DrUzgi32uVvnPcrtUK
7nVCfsju60ELpJZoPkWQX6WkY1DaA18BWI4GL02z3Gyn18KrhDy7NSKRYajKtt8u
hdXMK41auzjdScRyKzvtwU7B5MDOwV0IXpWKBytIcYfnpS8WXetRPrhtxSZaC6ll
WWMrUaRUxwCNDNrmiG2dS30bxd3Si2LxEjfLGw3k3BcPxsJxC3AFWYeWyfdNLrvd
M30psiiOSaTPkPjH0GYvUHaUJp4r8mYGHDO2P8ibU3DVn1gHsauB023igtI+vFtY
6u6w5m8d/hlOyop5HqTRAeXg/xOJZlbS5jFIDuPkw1EJmKqbMlnZHONVMqi/8wib
NPCCIIIf+G6JdH/UfGm7QU4u/5rg/bTb/q9OeKzhFY6UoSwA2rHXgpie7W9x5a1y
kFYTXvYCCFC3ItyrUE0Kwnlz9/nKn9ogxDKhcsnK3Ci5KJ56u807OdrJao0xCCHy
ooGjNRkSIMK0wlAyW9zEDtYDpyiccoTPdLwwSgCPvmC6Ypf7HbwqcjXAzw9k1Nvd
vC2JUr+Un93sIY7ekTAjKFbW6mVAZj7gh7zAAnDQxgMQrlgJE6cd1YKgXwDysX+J
BDe1n/Gap7PJaYM95T6nx/AjiLOMlK6XyhNbBvI0/td4kMXhrr8Y95cCQVJuZhsP
bXGVnXypdgan3M0dlh2XIDtk+bfVPzW7c8G3uFM5+6YWmT3PkxQaBWd7SxQKJWwQ
RGW5yF6JjJAy+9n2KqgiutwFZDT+C4i/nbPI4JOkBElA/A2y+rE1M/cyw6/CnyEK
BSEVI0mBzJefDixQ5zNZRAAPLN01aBTEq+t7G5y2HtU364l6Pkp8Y0Daf93Y0Z3m
wWZnpJA6XpNN1AMUc8Oqh73368RUASl8IiBbUdJe48NSFp+GIz25wk+zjobv9k7a
Zfax129Whb8mh2yk/pgNbcPgoZofyALJaapvr16ClJH/tAjD4sL++T9MxJUo6amZ
QhFQD3nWL9/dfBeN2VFtfOb+V8iQtGfZgUDnGFjm1r0TQ5aJC2vFinfqTaf52sbr
ueN8skBCvPfEvgMy+SYoeqS765XH4GVwphbsxz1cWyX/ebniVqNJ2AqtLV05ocs5
X20hEixu/IpGGUShZUrUKPDvbc/xwxa7cMN67Y9wTdgeLzzxgmOnhHkJv2Lgyvp5
FoJZLlcuV77YVLqHzlzQjJMVuOYTJSYnxjwNaxxNrNxOAysFNIiVC7eH6mdVUttc
6t1qKJPoYE6CR6B9rm3ZucdlYRyGfwv/OEGzZQxr1TNOu070k9Dmmb82aqSwOWm0
A3cNREV7CqAZ5dCd3+JLrPmrpxMGnUv+qyo1K/S24UiVdj4dXYai6oejwevpqiL4
sKaDqHveUJ9TnGswTStKerliiH3l/OEgEddjfetKbpUqdcsAl/KnsFXR+Cggomaz
KDBnwS4Jbemd9+WEuapBA3Koy2LrFKQAO+oOpk1uwRzXlF63IwxpPmPcPukY/d98
0htGKhbAZmtwo9ezZ3+3CVKT3fSbzDo3XeTGChQqhBFfr2I7N8GYf0Fxflte8M9w
ihEB3348zPLMYh/WPoALkeL7DyQFgfDPH4/wru8jElFtXOIIYvGRQoEHIOVKD9Lm
dPRQxcQ0EXN8+hsNozlgTQBoJHt+2G1xk9mFeDXe8Op7GwMmpUCuqGJ7U+DHAFw4
d9bF2dZQ7+Eu+XfECZ7CSxORpqO7WxxFGIcs9K4FIS/EUBQqe7BidWPsaSZZLVC2
G+QtN4p/7fjz++mWO3HK7uKQzhNaa1vM50MO7PBRKv7CaY20DAr+utCdZ7one4I/
VkaeFOMnzcV22IO3VY77ICgUDtYHxKZL241vTobpaNsZJwaJwrW0NTT76XtuBQS0
guhU5dRie7VxzJxo6Vx5vpk8KbzKPF4CEUOFCCpIkhwcGJMJX0FCEOm40WYa+IhG
zkuNQ7+LLHz2qWzcFrhdj0WXVsU2ToFmdPI3i3I6y83Z24S/DjRd9UMuwMUTVjF3
Z6NcbGfJdZhe/T6P1yDqJPAzYpIKztfPamtzWFH64N8DuU2CCpvVgYuGMjBS9GSq
0IlD5KW8BVxXqfycyX0YdMZ0lEaEOsZKxfDPAXuPAW30RWzIFR7gyQmGVzE7UMOP
eF1wM+zydF5o7zllbeXVil28cI04HighmLBBvV8q/tgwPi+ncvbOpeK0ttNsNyTX
GaZEu1rlUzHpnRkA1CwB8t2GR65rIIMzcYhn3I3XTPC3+Z24yGufP2i4GAS9Tceg
mYkviTv2AFRESp+1pdijudKnCsZKyPDj1I3Tnfu2gHXwJb7jI8qWhYSohNRZfS/G
JujYQg8cmjTboSQD5xeeuoBrXaqENVqiA13sjTIsUuQV2/6SfcXsfvLE4taVhY+j
7Ng2xaaIIIoT9PCA7YEoY9tac+jJ0n85b8yC6A/+3Lo35JNJXajF83E2K4XcTrzl
C5nlaiLoiYX4XkaTnwIPpUpUt4zV6HJSY0n13HcF3BLN9YSunzFayUVjve7dK5eD
z43kdhQx0G6wygwaH5VGAxNb7L23nmV08FMdizX7W4F9ncKYEln+5eYxMF3MZjwe
2HYbimVd5l/d57wukcBzFmlCztx+WLbMAv1zjBGSf9j+fIGy77WfOiTqjITczTh6
LmCzkVWvf7dIa8Gk+q5Y/fnuKAUWCiAkAHc8oV73sNCYxDCT3C8pIL2k/nX8o8mV
+bhZeQTeDljF1HKc6TgqnFEk38cToelNBBlywCGMeO/kxH8Oios8M/ieqtl0tGYY
mrY9lu+wkDGCJisHP+QaDhTKZX6PeuIaOL0lfuoDcjhcVAjUwQnVCbkdxodQyDHF
V7M+mNyXInJ5xmNSInq7dQS8PU9BGjA5N8oltyWbJrjCVzJrf8iYSh938dDLb4uX
i/XBk3RlBWOfXS2yd/lSgmzY8dM0tthupSoyt9Xf/1f/RxHv4cLeOvLLUCTJcWcA
o7KqQUZPWF42vEB6pAGGzQYEJQ/Bk/o11uKGFSICfxszsny0epKRo3SrL8c3u4mU
Kdd9GERdb8rV1sOLXPv4ZbTJMUHnRK7WpQSzC05ysMHgLhmkDdKEjW3s64Enmrqg
MOXhqRyLNIMOjJx1nuAomCkKtKWVsBa55JLnxOsDcC/XTlQP63Wm7/fwpuWHxtvq
2OX8gRF2vn0pJPYZWGPfCfdT8LAvKNeWMBUVeo0nG9d0FRqek/08dcB6zrLMgAht
0QpmfMImZ/cAvfUNAHndy/nmRzIEC+yjA7DRCJjTh3Ri60hOJ1puxZ2uC4ENa9CQ
0RiFLPUvlH2G1cLkA+NwbTDU27uwUvCH/BoND9SwQIO/SUbkEn9PZQgZVkHvbt+b
FnF8lHZWuX/u2w20CmX2lbmm+N8liQkSvhPIhAbOxzZpGXXZKHWVLk18yOhLaB9M
vNXMs9tT/qLcLGXjOB2c8crCCRbAr8vidF0Pwo8KSXD+vnTFKDlNP2VpuRc8TY4Q
imdnVONNfAcIGxtmiu2esj9bW6mzN/oiuIrzHh0uK7NFdAixNKAuaA75VvbjdSAB
H1BoUkPKU28NXtMxFijN3U72+P95EKT/8GoKn0sZy9/6XVxf0losnGCmDmCr/4v0
GD0avSrHyjIl72WxdWbsL9x9lwsPDaMw5zaN2HhHknuIQt/GjoGD5+tlHUcO8vjy
tT3KmSWtK7UPlQKEIR1Y+dsW+bs+t8ZQi22l5lVlxyDmqAZMVu1ZK7z+nxAfnOZO
Xpo/M/4+WqTUHB9fIfRqErIjCJQ8u4boygRyg+4PGs22YMhGBsfUqZcx/dc6MVCP
v7m3dJ9noPjCFxZ7lqdCTSTrL01D1igsWBimYa/2xyo3xxDTLxHAKYuZPvYmtyDG
vIUDte25ZpzFgiotxHPJIdJgYI0bwE+VCiz2nVE1Ttn2Y+q+327jbXUomoekB3uI
GUTWIV/xmyS+M1lyj7pjw4jsmYWX/rQpp+8yILICFgCGdX+C23uCtZQv4DTxe1IG
LWOqa5Y8HXciufHO9Mt4ufzcS3N7iYZar9lbT6RD/ook8zvhU0shnrgOpu8wBsAR
P19pkqRuorfWvwgf+E/OUD4xDGyNOhnMjs0qbF/yOXEM9HROtMLy8/wuy40/ae83
S7CEk25i1KC9Rp9yDv0iS2wr/jr7fE9o7+AAnIJ3Xxh9T93gr36vMEVg/ahw35xi
ZVnVCcRpcOdDyu/T68X9eaKJUAoH3DeZ19kSIJDCVYRpauR9OmTj2+LZxXpZJHnL
XAvo23ehF/NiEAVUmpS9+x8TGpZM9CtKRnyvxGpalrtFhHs1gysZpkZNlF4Z0SJR
UoqAkjeDOy+o1JLhiiRBZ/P58cOl1Bkl0fcWyxa0S8jMPzl4KJZ9PysagrzSjfkG
caGwwH7tDrg2s9LB/FZhkuSPEcalWkWzfpmr97kC3Z1a3TP6Y3AOOolQrI/HXg7s
iFTWOEFGtPJsJZxzBY3aFabtw5y7kWjeWo6he7RJyYdW+ax7LU/b6X87xxE33FnV
/8TDozz3DnsdM4jhQlTf1WOA3Be7XQcdzHwZy+KgQ9ZQH5zlsm2hOtIdok9A9RTH
9y6LlvhP6e/f5pBpZaKahKoyzr/OuMVTMRYLKQG18KQx4PkLanl3TqeRWmj7Turw
Y8DvKzNKEzxknHNyAcpv+SoFFchhVoJMTNQb8rpdw7AuzNE26VXql1wq/Vj7bJhr
mr9PQ1RVnbpXy7/698lTSB18E2danFPiFs7RBGSfURn5EVplfTU9zvxIHaehVcRm
/k9ZQdLXw9E07pa+Y7DpvLh17FCYjkO4ydTcjZW6W96zU5pu2ZRmIUdI1KrqY92M
px2NG1/xFMSAguZG8RjfAXti5uB+u1bsy+gLF5XC5sxCaralEnUAL73X9iQtvk0r
gW4MWoia6BFImqVnahuRMoFiMw8EYmoyjPbsVeG6pq5V6Dab/O8UqjxbP41Wcmjj
f02UUHPkQCA/zaigS0F6Y6AKcEbUES3NBO6j33/N8nFnxFlAC+m9Iy3sUD/kwvGf
VQXv1GNwjUUJqKWdss1Pbhgg8nIPqQWtL7G7SaRn6iUJiZbrasVifJeDGw+l2hmQ
Dg7K7Rp8KW1K0kKjXVOU0F1vREIBk4lWiwPTZFs0qVjU2HdKAsYMPoRikVq13t8j
S8mEg4kUrOX3vXwnE9ZnS/RtTXLcvykgbUSorM05QU/BDrMKLjANogYb5aFZ6gsZ
4OmxGUPCVhnVXTOiz+cG0rPWWKUvMCqO6fqf3yMGQX0qys8vvoK4+YI6FGPQBhNT
+WGlmQyEt69+eAoReZASVYxLoENumpbrHzAZGmVXDTpAjJvQxOyGIWgeaIhebWJz
lnVzRzWNgUBYKEHDdSmz2YgPG2J8XrcGF+OAnuUxNhgwMmGW5jcuhXac7Po/SGf9
RqccK6h1TYETN9yihPGKSboEvGNPfhWvQ8GimLLJ/qn0Mpr/QUdezJZKafCJAUBE
xqKSIvWbQ5478jpc88YwE0F+gUCONecndxUkEryz7qtIIKdyodpy6qW6m4tfuCou
ePlbPVOj3cB9jlkO/LHxPuxRvgyW6FTD3wXRzmd9NtyiYk7fwvlYiV63F1MuOfR/
u9qFnTSgZkaI1UYuMGW14m8tJgweh6zW6Xn7MQ82ljmTQ9tfey6AzZ47FpPlsJ0L
mqvbfJr/tFe7NmbzSc94CMjicIPFbo7VSKwn4rOOCVmxncs9RxfNYEUdDw3L3O+c
wGZYrQgzBsEwt03uRSKm7oj4f9povLyEgOgBgX/NzXhER4ATLn2Zexid3CVF3W5g
407KIqhNAAZ7wfKDWlcQfhI58OpzZRf/3KRNrkUOqfGPT4Nad3qG8/KxWrliH1am
Vwk5tu3q61UT7aVJNH0GYfZWguXjbA5W35ISn0Ilk8PbDe5Bi9+XZkVII/pQOFrP
F0Lg+KdQwL5nGbLr4N6ZuoIbm6pce20qsrCzJhlaotgX7iLXaqZSVqzrOzWWa3cc
2YTMxRuxSYjYnTXpeXc5vff7kl2bCpf64O6LJJc346U0wyah0g4QDv8ZoOLX2sFF
26Oh+LDCGnfDRWU12fWRph90HvGtcwkm09K6BiMy19XWcu5XSF7ZyLP/JvBhHtfB
Jvo6FNXnGgzKJ+YZXRBiXVGsqnbGEn2Zw/Cv/j3UWLL4tp4IDnZIqTlDByM6LNEW
sMjATCpKwxyhAGjHU42Ub1+Dk0KlEVlY23u6qUtUCb+zWnNCWH4cZtaK1BT3cLXD
Zn8Vvg76vRixACP4XXsOnoMIcOzW6Ye0FH3wn59yJEQv24BFtKFZ2NY9rpbsseAc
K5+leyozSTNVwqmnXfHbxaK/8o5Ut+d2M6kHw/XTem9z5s7/1vj/2Dg5JOyvS5Dd
VgT1VjcQyg+YcObRKGlfhMTxXoInm63duukZvVNuTzDdesTOz2csJaH9Xp3IUUb8
fhjziqorPwi3NbDL2X2H3qIDbzEuKgc5wUyBcsPOp43tHFyJOwvP29g0lGbHIe+m
Hs6crGoIuUTEsj2el2XvPmKBHN5bXH8V1tnoJbtDG98aj1K1tYkaBmi7qTRtLx1I
9WBLKiQgzirwGMcDfvuf+itA/EKpRfHe23W5qa0fTeVqDAc/As+Fh+B1ZV9A4+Wj
TPC40zE4f8jKRzNBfLzxcAjRbufgpyUEUDmJUe83lTW/0MzE9jgfBmZlzx0fgQJi
1BACGnul/xjwvI7sXoGK0odsaAuwG8Oc+NIuljJr3BpSLtRHR/fo+SxUqXwfdF2U
UX/OMvm5We/+p6BxLgZ181AeoUTdrKIj+RfRItkzaFvGOwKMtmS2rfv4vUrKlXUy
W7TtHw68t1PyfYeHMBL+tH6qfqiRKO8IW1UPyLs6PvJOuS4BuaPpJ+mFjWG8uKgZ
z4I0mUwbE5tsCs6qbbj4D0n0DP+lxZ+fE8U7ekITohuoPvKvygk9iMFseyXYPSSd
CtImZFcDKVIWuIBPq7ed9IHmJ4hMbUCDp3RIhzMMD/pUCSw3lh9Ikji4lZFj7df1
kKKVUvM2N4pcg1RiNHwlKgurefHzFwytz5uQJZ/qfN3QvLWAG3H0SiMOHfamOEJ0
Ns+vDBkR+hpfkyaGuBDYKbP8adjTxYpvDsFV1nbnK8wmLdWrrmMeeQGRuWrAZKvp
QkqoVLOgnq/Mg0nhJT4mE3k89bkUyQUtzb7t/IJKwI+bfrvqxY4TVV3KuYnOOM0Z
ecle7jPx8oWXD1r7g1sWlf6++gVq2XJdcUvf1IBNVOc8K/kbLP96L4kd6qpqbxax
wPpjr29wyJEdNSyIZkFmefIhb2scxHsq10I09QN6PFs3VVmIVC1DH86RXWsv8fs5
TaX+nOvVse/MILxWX2cKNHXFG6x8Xq92ZtCdG2pklm46iqHSnL9truYt6uf2lMM0
4Kuaw3EYK5NKVZCsiMIU9XCzWVpO9Rq/d3lkanIY6ECBRVxg//q2VomXPNN+/5qD
w+iGho4RV7faZKmodAeOO+T/P61efQotk7rQdTMtU2ePG5LN5qaldZYG/x7kN9jH
oZa/H0/TVZkDD8pc7c5XOgOtSt9kGkDMrZzOh2Wqn1xWZNKA0kWPRhtca3L1jdjm
heTyqspFHqV1+gOE62rbgle+VGyx6kdCk3GaTl0/iUmEVCZR87fovpkyJL5PC1XC
Y22PTp68HPYta4ZhrPJKgO5wPKtX+ROoG60iG6OL5GAHiL3F+QHuw2mEql+biRR4
nP32VE9dwmI8VV5yGkxVU+c1frIDcQXfaesaaHLfsAoQxF4wKEdcoXS3pI2BMcQL
JRn6SwWovBXN4ZIGiwM7MoGy6xsVv8dEKwp4SzLNQMw4Uk1KQ6WG616DTz+GqVSX
QZj5QSaiBfLnAlx8KmudDNCRSvuOrZbmFNDLvLspXwkqtF57dNJ5mmtTjUKuCQl/
NkUCKtPGBNZLD+QKdm3OcOgH/iRMn4piab8FAIBqw3uNgxgVlln6mn1FOSdKTAm6
2NFEZSjAIQfPbP/qeJa/2aArf0K9dne/Gae2rfiubkc9VQ94LwwsyOKQh6EE9JZ6
90AoYg8pDKSAYH+2vmfdW26si99iqHOHEdOuwmCgo6C1hgkdCXod7X2jpcu5UV9G
uE2CU359445CM0mzZl/oMaVXi8KgZg7xxRhX5hOq6g2zbLSXr97W3qkJNN6bbuh7
4aRPcZAq4KeCAZ7Zsr1HDAC1sC9WrzeugZ1tUADF9hFKiV6S3hcIQFEJxV8epY7n
4xRKZBUZu30Mzn6fsgyT7EPmu2b43D4BS04LeJM4PLfNWA1lLyNLRNI1OUc61Xdz
M3kdjfumZ2a5TAT4PaEMxNKtsNevBvDel03fmRVQ6VAF0UR4ELczt9JghzIgphPL
AjZS6LNGMc6Ki5M07NbNJnnx5UJGnkIAT2K9txvFF4MmtJuIklgpXGDhTMNowp6V
5GYhhy3epgzqcBSMux1hq8riYJL+x8zbQkLWAbeKGiUWSidNSQWEdLXujJoWqV7m
A0vE9u6HuLaXIC9qEayPKF3jlXH7Zqti8Jiz6cwF/iekyipf7Jmk1v1SQ+W4hmV9
JMDZQnAFL2H7bk1fpUwMztDD4Gs7loQm33LH2X2qtQMbMkEjNJGCDwhmVi/An6cN
c6epFIqy7D6bmssMIAh+ALVbcjkQ/ssPEaLGzsVgvk337cABpdAyImkeQt/9tbct
WTk5iP6D3r7cNwSGAyYm6g1XIoANIDfetyYxi+5EOJ55WyCq/70V8ItGQRYWR8a7
Ozc0hWuuDv/hOfQawdsPLxlPnjp+3HecCWO9KuDKOSDPoWWD4Y1m0B61Ncc8zYBy
6lrZ+K3pa9rGOOleq26Ayp6wGtZVYH3E4+4UYM+s1fssdoCV9XUHvC88ctIjI8IT
SoUuDHmR7Skhds6ma2VBxGjIN91K2r8i42XZV6dew7d5sJoZErYvGfHWcsTAyhIa
jFJ7yuG04pN1eKmkMeHg7L4F2q7VNWEGI2am0gHNdTuYYZSRYxeGsVIbSTinS+5t
9nuxpuMt9hlx1GGf0iBft00KU55OxVVa/RIrzLPQaMFW3+ws2w5HhbsKChwqxu+m
dVWa1DePZx3aLMsFF2rKl6HVNvQ+5dYu/HFkRES4zo7XtwMx2tDK00s48pLcPfQk
42ZmF+rtiRynKwlJURGBBz2cH/I9F7/fXh1ZOy2u+rU7ZVvsanowE0TUK0e2EjYL
YPrdKO+J7Qdl3M6gWW6aIbJyEJjABj9Kimi82i1g5dDXddXnvUGS6pwFAWruz9Z+
tMVegNJ8yZq+ECux7FMciGH1AYB/XO+oH13Kp29usTnUpfG24mMg7LlNmgSC/oXZ
oHBItp7h9pz6PaG9WbYMjeM1FSDecdlgyva60iMoNwNcj12H94ZBd5z609csblWf
Zf1mz2kr7OW0ZAucEeVBIMjTqAT1QcmgQOE7MA6LZqjfOPbFcpdD1I2J4OpQ2DRn
gUjSpat21kXhIZfS8B8yer7gaboB/nIvmjGpIsI9EYI9pkNL1ZLXhMGF1LlHtZY6
lUCgMOKm6mxutr/InKIG/hHBC3gDP7BWnHLMoOZo2bcjRX/LaPLX2B4mUtULQz+l
9nBjim8ROlnoHfdMGDZXOUpwSUBQhlACh+T9JLqhjp4EwC4r5nT7Wxws5ttjdpix
Uka/vm9q4pRW5TfIRcKQJdncSrS72ofZ1ZMWRwZZ/UoNrrt7Nb0U8M0222Nt0QjQ
924VXFV5by0P0a56t4KrPsZD3iMnmMD+AJ1Mg0EjeQIFuIMLWE+DOk1nkggJNO0J
N+qsJoKmXQInmgXqAuH/lD5RoZGk+Fr8l0kKSoKjMF9D3U9cN5nUUcGFo00bPsub
Yrr8UBs9zfJqGXHTtIQ1un6tU2CElMU4X43Y79fQfCt2MHCB6jT+4ih2N3yeHuBW
2aOzDpJDsQp+emEaUCZ2A3R6GN3ePMTffI3CMKsbgBrrGoSwBzz9lIU+U0LYw4J6
BXqeXzIMX2N/njW0VLngOAVyI9c/tsXmIRD/fBLF8/x5KYjwSvzU/17LKT6dY2ZL
c3nJThhCAcJ4DdYtfTiheP6uJll6fhauQCBI8A17N3ic9a2KfXSZkJZekYCP4gGi
`protect end_protected