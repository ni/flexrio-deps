`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8224 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhBNVMbsl6PTB5/ApNH6uD+AxODPuZxQZYuFjLlj17wTl
A7UTN3AZY/Be5WwXqD4f2k0FG4yjoJUmHJYp5diUDJbaNMtYHJFEqhvU/hHd6huA
W0/1EbF2pQ2I7mITqVVzxySeUNq9jd5QFQ3t/IDWS5qElAZzc4EVk1WcDqZ8KC3w
74k4kLJwi2WO2IKnSlVldogFfaP4da53f9FGoKdtmwoweTTgDzP/cby4GigqVi1q
yjky/qnsI2vtrvAI7wflhHmfQozGn8QmCzDGDyjBKW7NAlATvsWZCWKR0wwetPsi
For6m0qCJix3WmYYD5675+K6YayBH1xe2oM1cVg8/PtwLnXQkbQTYWMc0b7keGQ3
hDGRJ3jQqK+QaBlOw4gE6ylNnS6b24X5AU1TsnD8MMACxsrLtbifq0/oov3zSpr4
PpQp75ieDveNb5IqmCI/EG6qHLABryDY3fZcvSJeTt+97VaJK16+/akQ+ug/4IyX
GAHL/YN4yIEWHSCCDcKvEoJWBQxhSAh7g03cm3BOWf38/Qo+pl7A0ZhMTiPhoWIa
x918joa5wTUpNr1NbDZQdXffFOKpquCr5qz25Mc+XF7AYCXugssH2p0IkzUVWGkO
wT71KsmgZHcU1r6iRVeQfpPUcG5MO4I1QsKpW7k3Vg3vZhifPO5mtgyWGyOh7b8E
4F2fgm8FyfStAo20KGMzd5ZQ5LYC7dZPiBSquZ/J9aD8KMiuK0OT1cjiVYkzHRah
zs8G0Ib1FpsEL9pI2S04Gw7Vm5fqXlkvUrENAkcZ5fSOiLgVWqQaSa+5wojuJ9DS
1Pt6sVpFBT6KcTk3GkCxI4Op0ZLMuwpkerq1c+i8wWlm7XAGwZjc3qbUTHzYMM2V
5QCDAPcfYtExP/tPRYPkyLJ1fFU4pjf1ZM7t5FCtWjoTdV83Hp1TlNVYDPuOxOyL
UdLqhzr3pI9bUTe5j31oRQj6DqC5po9eH0DIfqoaNiV5qC0Surkrfque1WtPjw3t
qkn7gQJa1J1AeOoK53AIK8QPJhcX4XiEchBruFR3dB/QQiEgA5U7tXL5ifQzx5jY
zJcfbmGHJR9oA7z+DGu5tP1YKYf3QrvkVEiQEVum+FvQYRWOHYAJNYQ8cL8KU+Sw
MAf01MOkkcwTVHAW60kZE7+aCREYOqnz5YpFjI6GCtxHJmjafdJiSLeB+3HEqsOA
hZQzR1hRVcGvPvdS2I4AN3Tk7E2HtL1RxUMyuIbCXJ+csHotsVe9xT3ZiMgN5Q23
LQQRtcGRvEYjkMivxDCMzUIx7fz400b303gEHp/vxjY9tAUoBPwmySRyIGuQWims
Qngt4CNUNiSxXmkBNluKBwPpRLFy0yU7TIEFfTPB7v9uLT8eEKqqUSi8A0jNsxMG
L3EtXwMAdtyVFgcnZKweONRL7wdcMRp9CgL9MNin/sUjVgzIhiOCv0AUiEGXyRZZ
iI3SRx6Q804MAGahk1IXwUZAFjQnxIG/WusgziHfHsIVrSwXwjo6uSf3ikiCYoqN
6CakD9hK9J7pqxQLcWkN5mAJEq7B7ybwmEj7N8ay5WKU0MEDEp4+JmcPpYLzodL0
RQxSWytenjI86MNLzf5aYotm8rEITA0i0bnTljAAQvEFgecZiQdkknfL+cH5MJqa
aNrfTuCu5Mouvf3aaFKSCFsrCMIm1fOuQL1blPdYdftmOID0EjVG5rmdcXRl0jG2
+gCZg5NvRfll0r6pHSPgCM7CVyXp7fYRLiPnpAvkRMrk2HnObn9P7OPpISNqKSgF
Xlzak6pkvfoGxnCLQ98zaidK6aCd+LmAmNkB/QrUyrzvyZpfHRe6vyTONCbLQAZZ
83wx/TV+cAybJIntNgZpxZ2lom2yp+Bl3x0dFfTvMY4VPiSiNnHOUexS5cU8AmUf
QBPGU9Hdze2km0Cu+m/98cRuOoU85sCS9VH6oeejoJR+on5SNqvpn1fP86e4oGlC
WpkCQMRtCFDxJbNmnShOhVfwrxsZwfmO0xThqK4F16b0JRM8dwNFbTIhwaGLV5X6
dEiohjbF+ZAEfOxyGA0Skpb4jOGVxern/+WN1JsT02VN7HxRsTOk/aPCLlIGDbbZ
kuD+otryho9fvXN6gjYYsXByBSjB/5X1qoGRFIF6kCZvAmjoTL3FoONWMW9ydm08
mb2uGb6UugJZZaHNp4L4fI36JmaYjVpf3Wd7fxNk3Cb/ga91ibBuYRPlLSH2i4Ok
MzUpAJcBi5Mb9M570VNfNeKWZ70mp5n5aoszxzFomUVhyz+hOT9KbHxYdSv4Ff3Y
159Oa9tGWEx+K5i7JEbfK5RkpfG/6STMJ9mNqMVKi50Pk0EBXMPJwIFUBHxYWG+k
AW+WSc/huRP1ZrBdpdQJby/RzxMx0m4gVZWpQ2UHL3+YunfB8xCPkxDLEDpQk2jX
8ZYa4AQhILcpaJV4z3mHg5z2IPbZAq7RKtk1nEL6j1g/avj7JeKLMOW2dm4btUPy
P8tsLT7Kj1LPNqPWWNAvXQFA+6shWdvl4bOKOQ3i2HUr55gJiiQEyyZvY2ohWXLg
XK1wuucw8S91fuG/Svts9Pf4WoMkogKYhjMFgQbbuUbzwXfQiESBz8NGfgrAkhoO
hf74QtGwQ6ES2l9eLbXZUDLWqe7ptoFaSktrxUU8ftGv4B83FdkWBPrZj024A4Kd
ZqlLKl5KqQWRYjEHWnVOBydWmaPPf119M7UvPiuOXxGLHZ7MZMQtsuZmXsRkkLH7
EtbPzamB11vfl5AV+tKoiHgXazlQCTAGeReHKEk8KVxRy9WxpuHf0AO4Ej0kAjRV
d/vQzZ7cqY0XV0SDsqV75mrGrpzrcVAnZCkAAkjTPXmm2MaWJbRxulFZxAr+gZrU
3v3BQV8m+vgbA0+JtZ/7Fo+kp9ceaTfR8eKrnuM2rK6ras803NOuIQM6JCwrCqCD
XWNfv7uQjFga8gxX7JLkeLmaCNlcoKGGZ0unajtTEOg5Z7nX1OHmPssELuGckI0a
8RSIL2k0599bOFXcXcV/TBlwz1POH1NM5qZRX8JxSHpk24gOa6405ukikEAAd1Xg
o3UPJN/qzbjgb0o5vKu8HjHHhI3Nmr52Y9+MSww2yeb2xQd0OYC8MzjCygmAyAUG
zYZxnNcr1Yf4YAJL4Wxi53Q9QaeGPnr9j+1bdUNEQH+iW2AkZw9yAYWv9ooD/qYd
XX1hSSjzpBUPQ473UFrJ95YaIIKLKmc9lmmJZPZHUzLEBLynhM8ZouSFaWUFxbdt
0fsmSTxQNTtES2b/bG41tcF6e1Z3GJsArtNYl6qrd9dGVxTYyRF1Ffp5KJuI25wm
8XPVmnl/D5t6WTLCKH2loUUhCQD8cp8/T7/svpYo92wU9gRKdRzVxkGia2WDKMiy
Srl06emPq6c1LXRSuKlkrq2I2cqBPvR6adq5BZS/LK7XkMYfpwlWx1xWhvJZofwd
/rx8FdmenkcZzUCdAnaNZVaCTQfS3C/7l4NOqU4g1+59gpyneFtrdzQl+QN0jsy/
D60IGYQod/BBqDS8ZpTpneAfaw0O7ir0A7/6BWpmj9KnHXfD+LvqOtP2fAflbH8s
KnkqTvz3TZYElFbkwCKaDI7wK/43m+RbdzYsIoym2NZ4upz8/VQxHSIT+rhODfds
7eHBD3dmAFWxyWo6FnfyUCEPZRd8559d+v9pVDVXSD+w0tP7UkkxoYzQ32H37ZXF
dwvTheDVz2r+QOgwKnMKUe4HF84oXqw0oVoQsMJ1MLhW4K45u6JCZQM/cirZDwBS
IUV1mgp+NTEVXtkRfoxWxUA4ymcR/ZeLCGZZUongJW1fLO3jdgAQzzVN+0ccDUyW
W33SB2mJKqRDfF6Psd2ygC2toO1i620G30IddiqhCkE3O3OAg9gMZGW7koWp6/z+
01YpM1X9/zYVBI8lzoDBHzqyzP6YYHTBRkfHNu7IF2WaDf2eqvjWOyxNZl0/DKbp
eJ/rQLHJuS5WYM7EREhCeNNZmBno3IFy6JA17MzIA1S8edNDHoTFj+KRW1UwJec7
NIPHRglfHJcMNk2o+vZiGL7zsLdzPcOjwlHOBYUEtobTPFDOQbo7FOAFsRhsoWqj
M4KJOkpSrjsUiihHkJ2Q/89hIzmohzyGhH12ilLyDJ4Zu2JbMXvb2HY78znqGuxk
dWnTQSPkekp3AFwWcVHYcQ3fecep+ZZu1IaFmDFw0coJEicQjA0vsZpHVpTRu3/o
yDvn1afqdq0fBDjmwDZohb0RR96TCtqaarnbCqQ6xTQi4z/UmqqfBWn31ySUCPug
qEn5XOERalfgXtJNg8ZOuGWYK2+sbR2PEYwE/9fufYIBe1xfEraO9ImKKbnDdsRe
vQGsT75zcz6NcQFDmkO+NADe4pb171r1Tn2c7if+Z9VRAheNm+DBxB0F39gBlbF/
AjziZEYMBYVuijhIPtXgqKxPd0Q3g/MCZhkONfQg6OR1rIQ+/ugfUdGS6z4duDc8
bNj8N8zSTRwfEbHdDVMhM0Zm4gYR9gYU+pKA59T7d+QpsGXUDSNcaIKOlrxsAYeN
VxfUnVoKsdBiQwGfqhV8z45BqqmjbByHuw1Yfx1vIFia84LfLApY39pZ91KfZ3HB
SmCTYa05cXpoL9e8zM95hPT/H2yDPmZ8EqglFLgu+UXlNrAn5y3xScx2rYZo2LQ3
wH5ARsmzGvsxCZFjQaVR3OTDjyLxh4Ggh3olXLteYm+x7jSBmeRD1csCQCeQGFUl
rzX3hXiAZqr7HAGXIXiCS2mPoYRuvcni7OTaJ8Mr8h5E62AjQrbqdqSoioVFDOOv
B83Rfm77XEOKYBGQof4+qggn/aJF4k7QoFJw2LhEyFCu8y4UmE61uW9NElBggWcA
vhwj7W6PyWud/sK7pURLVJtFFzaQTYwwXhTeToTjV1zlOcJYzzG83+N67JS1N/WY
59J2iS/wUcMB1s3o3yv9sT4H9hLG6QVeX+ggSyVgNT/RKlNGKVfL9FEmUH77RT+K
jIZoRCc1Rzc3XI+N+UECzBvmnteBageN7bjBq/1knJcz04312PxjXECLONST5F3E
I/G8HND/t16Gyv8jWDDlmaiK5EbZPYermCKo7i3Dawifz6KrocG9mNpZgHuRVJZ/
5iS1WCG2mxc+UQqZeubnxzmgKu2T/p6Si2gB01zfaCD72O81vYOQ4i/Go1CT3236
dpsMOAXP1wPwHkU2OvVOkpTIQlG92uqmLyCya7UlVrtEcmrJgDetE8vePNU0XHbf
0L0hQE3WfPi0QxW8KnlX7k/Uc1Lc5AurwwANvXfrywM4rmHXD5PRoaBH/1mALbMs
pG9Wx3LZeI/cbQtJs6yRYQh13zGAWhUi2IROB8ADCicWnS+13+qv0Sn0IXx3RiPe
NZu9IXAUBQlP9AlBFEF5MXSv6IzZ5KJQij14tVbe9mmmKcyuRVO3pIGClqWdybsq
tZmPsPC2PKQW/u5hnCKfTR+sBFhb4wkierTi6qOpvQvjjpv1SmoDzMG0WCkJbXiv
ADnlIMP8hmE+jGyuT8QcCaKdqV9KUrvpqb6uSBcTsiPFdTH+N9AM5UCD3ED/diUn
o1fTqd1RECcmvbur5eCXvU+kkvTj21sNC6cwuhGu2HRzZoWEZszROZSIVVdRlkhO
gN400Nd0iiLMITWVuwwasK05cWmQFDwJWN5nOeYMaAeSdcL8uQbNGTNgMeXp9N6l
pumk0wuGSDxvb5FNMrHhrwrqkw1A2ivEfzUJz6aXSDln5aKhc2cKBDok7sj/PTVf
TTeDKNfnZfhxNnLH6XoH1vUP/8Fkp/uR/VEkvTZsDLPYcKyFaVnfT8KIsQEz2jv7
xzCU8hMkkAzrNq10Icp+KOzex8Ek4l/MlcEYLa27yTslqdUsCQgMp95kJ2wyJ85b
3KXWW6trt2hecCR2ShOccu7A77toj+Bk3+3tf6gWOMRz33NC5kCbZrM4tUE6FImc
bplUloVvS+ojcFjpg4H50N8Aj4MYHT08ycGD3SSLeC9aeDeHDxclNJISsJ5Yzyzo
EBCDI/sFRNiutz/41BKUpbzvATdYuU3OXZYqC52KTywKHUXiBG+mGNuJsiUQDjCZ
VS7NDv6VF9hryOARzqrYtLPyi5cw7DATCJa6t9Pt+PEaIfKrzqOFHn93y08ZNqTo
+dIBKzACB7lC4Nk+Aur2109HO/xex7YpUdHdtJbgGq3awk2dyuz54/sqN9ZFoxmO
bEadlo04DwhoUJ3fqyz0FB6mkgG2pf9VgXUbZ7ZjCLiNf2pjx/JUaDt5wUm/sM9M
D89QrmlDbPaWReCcChm4W7ufP4thQO7cgDEtrOyMLwRghovsoeSyHuB/G/7mEiOS
e42SkUT+pip4wX1Ht7UwJIU1F5rW/nBRGX5rslp3a66yW7mDm/E3tzfsDFxLGwLV
1oKgAyzzpbXIp52Ng2OGMuPHzkDssNQScKHItPaSklnPFix0TrjSJw+oq3t19Li4
wCF/ZBEEkRHXe53Yjpz9NDq4qteBlNRRlzijyIoVXqs5UhA2TvcYrJdJ/9T4S7Gy
lnCYIC/x3TYIH7F9sXTSyNvoC6If3GWLPzDk8NwSP+htZIjhgokCQrYacSJ4NOHJ
/yAdxi6NNRpxNj8NfFtuP8+sW9Xh2u/wDqlHDMnltpTArZf9uoidCznF1+0kpwLp
ALh3wnDwgTZzkoFOIxYDYxu0ol1bNlZSFXWB6vVKu0jPaGxYkUZFMIcqPT7X9v2x
GbOfiXg7J2waD/Jco7J0KRXaWttbm59Pxamuu7H9ppsgg3f1yWWVaC9HDtTM9FU4
quZFtQorEpgYIyahtFOoRm5wJyXTG2G6+PdM7GYBy4ztWDvOcMxmp3ewmiuMiEIn
PyiKkYWvpEXxUEssRQ1Iin4ytAEm1upLrEM7ccbOC3iY76fSubrnNPb/I+iHubDo
D/PRu0zRDHVU4+SYb9VPIKrGr6+ZoL83VZZ4b2XJG6sNBRgLwe/+zGaI4PqXDbuD
zHbRfS8VjkcaN72rjh4PGiXSo80i/nqrgki8hKUITU7UPuPs1CbTzzUCuW0wqnmU
09hoYYZh95V9M9Mk8mcrH9y6TpKzT5gCry5J/5xQmFSLFZ1NwPtPPxnPl6/gyKcE
RBJEM1Yno4Ot+n740CuWQJ+M1NZCRHPysSfVeWqSbdTfw522Myvbvs0ulkqRsYmw
c/kSQLcuXBHYQpX1kOoaSD+BQF3KkFYePqVnRWftCYR4PYYL8vftp7esUCBcEbmH
95q34ZSuuoM9BVQ0nVFfc0D1OeWIua9zBQhvp8ZCtGu6K/erUGDQw4zcp//trTzl
uRqvhWKnKfCpKQ6Q7tkPla3AKYzEJNebee7PJX6kg1sxI/kxkycNMCSTzyyVgN2Q
IE211kwhj/x+tzIYzBz8OJTkqjx03i2WPITXQV/9U0jD2neBiirTcB49tVE8xkFZ
doVgtApGElts/gMQaOwrhvuCzTDmR2uYUj3kPH0PcXNBm7ZhT1F8OIACVTTOz4sF
kIet2x7LbUGbufeeopJvqAkFqDD1YqmgcmAtve4hU5S0uhl9fTJzEPB/pEj8G34f
9nA2hhFN2birK+2k8qc63e96y1gduAMq4s55gU8SQvxUT5e2qJ30Op2JE2do5VZo
yITpw8zb60FBo/uTFLaMvdL3JVPhfjBUkV1hW60Z8Co0ctw6bfvDL1T9cUF54xBF
Ybt4cgROiRamp002Jg5VGtsec2oCT8QUy896UkoPlHNYRJWTA3o3CQqtXTp8nGvv
nKdc4lO0a1w5ILz93H73X9gn8Na5tkZpfJ47ecZsG8X+hk3ZrEn/60hSaOYpIQux
tvcs9cNK7HuBLiRCmv0mWikaq6pJcswKD9wG8sEa5sa2fTwYZKEoYOAM5mwdZytA
/oZ5FIBu9gZW7Rvam4BYi+MUjSipfN68ejakWS1oLU0YHtXTSL/PW2Ls7dlQtrb1
qvRlklwDZkERI0V8Z6ILFKzeyWqLBFKV78hhx7ic2j7zcQTS4X6cy/id45xLSnn7
Gse8pqL7xxvXUk04L+FMj0LK2GSYytQ78Fp5iofEmUoUqZoD+rEaQe/mdW0e1i62
CpGdf46sP4dBHZwaeSGFXJLg/4kfh7yz3Qg2bP/eaI/aqKXSrrEm+bmzxFvheF/0
hJW31OfO0hNY1ay35ZmSEC5jZoEMU6RbR0aBfMF1VHYK+IJmMTud8epoEBDjQXkI
k+dE1FTTr47VhP6wpXDLqvmJuF7XVEYt9jXid9QKkp3w3VvxbwfzP2O40KmvCz/p
siBm9LweDpu+5T0NnDvjFAEqTFxxCoJ0LeyQajzkRFJfn6X9gMZ0EoI39xLbWjby
H9tuYsUwN3WosUZOp34Zq5+u9zVbPu0BqT+Wy6smGdgLRPS+BtE2crFrmbai05j7
y1HUo8mcfaMY5K7sFADzmiORLRnp+FfB0XCo7zfL772IKh1glUxgdGYmF19PidHc
h/GxemT8z1wUDjmi4wOMwnG3WMT72HiZZPYaqCKbNZGeb1EZ3vdlSafTlOv0mw0z
ReuWb2ZHwJQ5wu3LLHx/sEldD5eF5HsxqGF2iFgRdIaUfM7BOoyQj2JQrdHTuWTB
/ckjxsRzqWLNRfjX/3pTjAf+y1cIDFN8THLeRgl90taG96blntGhXRuc2h3h6NvA
efHc6qNPNRRMXjXsRGV3r8aEjSxzUI+dpcdJ+rsX0uplgDJkwsolI2J9ENN4uh5r
cUMgAyDLlh2tnzgpIR18uKcW0eh/PLL5jsqr4H+2AOBvtRj4uB4B6CzLTnwvGwYY
lfjyaMKo7K6myg7AvO/qiAxDLZdhHln1bRw00SbSEBQ4PKZz8hEGpy+mJaMhPYW1
35K2Q1rnZOeh5+9JMOqjR+z/o0BaXV/tMTuZIV0NnIjgEa8YQrQcwLTaxdcptxxn
+8I/oMJ0Y+3MPqBJgjQiXVf+CozQacYUcCCb8Xhd2lcszN2bctW5q5ye8tV4b/Zb
+LGvs5qq6KznHAUWuJIII82KtjAoEXBGRO01SiOz/P2XJ0woGAltrJDREEYTU2dV
eKCYgkdE8sXeE9sguwQaGQb5f45LVQudc8Kyi3wMmjZTb2GKazIVxW0KT6NSGzWf
i94LCZLJ8xZDAkLK72YrT63QPe29OMZ43WTNfzzhC29V1w4S+LoAYn7VtSOH/fDp
IJJZN2mXY1qGs1YedrSETk/1W0aUsETCrGZH2b20ip8zAwOiAFfsmNu3oZ/FauU2
NRWil6/Roz8QtbzvajZ8cIqlEwSZW+N1mgP70YoAehDLZGCY1RHiytg5HYe3qFHV
YYxwq4wnnWJkzm8k04EzOGaZKhnlUWrm00Wa8WGk6/aL5KSynKbTVTa9Vkfqwcxa
xPK59ZhFPtzhQnSeCw8h+2sYNMgfdPv8LAlLQBwfDKYp1n97S6QB5VxOmIRf+RFc
yb4cV58m3L38lkwsEoJPqA8shUOerL6Hcov4DyxjVXbpXksmOHAo1bGqSr8x8Za9
F+fQ+1/E1r/mdNd00s72kpUV+tz+pC8rSJ/lzi+XKSbjZXskpzWHPFjDjEWemyNx
wlEfAGbhEoOEZCSp87dvhTgnnbQq+cHlrq2iMa1iYrwBQEqGA4N8ikT3Cu4Mb1gG
lth0Yx/b9T90LlhMtUKIdVh5ou2XwWKoqvHyreZDD8g/dkvPbGU1d7EmRiWu/28l
cZHWhOTlTAb8Z1vPW+q5ojDsfnpZL/9IgYFh6f5WnZP34cN6CqIkQBfe9hRlitU5
f13MENqpVRJbRFLR6Qz5TEodrDk18d51mnw6x3LIUAaOXlU8LbxuaRVkBhZlDD/0
aO8itMvdDBWwMuhchEQlu9bmT2D+RX0/w3073yz1jZ31UQWVmYED4UY6qMDktbVV
ftPXPN59hynj2ypgmuxIyRD7yBrXvWotqhs3vmF+jU+HtI9vunw6bBoqyiL//KBS
gPHxrkNseNMQZ/tmdC+0DowXMG72WNZ9gsIhM3hXDmyjjgHR43Wo1COU5aU3vMCx
wS+4VIKaEE2i4JA5/WmoGaoz8ZWWl6Ttw6lm7CPSqsKIaz1uEN6eqSZ94ALeWHzP
EaYcZ4IWmREZPWoMIR3u2VbD3wSA6idmUoueEuKtnusi+ed5Du4qh1TQPsSYO2pC
pi+Rts6biE7E8nabpNnsGg+WtC1asdL67+cqKXsynBym53M8sADdG5LbuwnozpNN
XOp/KDUdEDPHzZipUaTdQXaUOe3CBjzHlp75HCVcDeeJ0mKQHI6rNblDvEMfzdyH
WWacBdfLuJxpmEfEhhajf+yVr/V55XzxusexWrNmgPPxoMFhkHb0Sgqn6v3/63WP
chvOcKHcQxcS+Ri3A5cYzrn1lyntcfYAeSyJWFOWO+7J/5+zpNJabgxVB/C3PnXm
+B4txEYevMQs06dSqFUgEQ09qYeIRMbSnGcAP0+dh2QKwq9imNo9Ts95hGFzBAyk
CNwyQfx9hUT4OuRB54kCbuXNZBNijMCwc+wqck549vebxhPpGwOIbW05hFvEvV26
Mmsg5mdDF7gF328TW+zuAPl1L4Ms/bguonHXVXEEzyZ8jT4FcpNcrJHyujgmOJLh
sX7vBGzbkkNf/9sYbq9I+j2WFKHgH6EMQMZP3khld36utpO2OU0ZfQRqIZAK/LnR
YE19GWoiMIKTfBgfrY4KerAvnMdM7XsBz5mTwQpzQ7/fb4fW2iFE0sTbsYPeYeFa
KB20r/ZV/2jfG9DdPLOdWp5nB5Nn4KjJlbkUgKEOK7G1EWFeCUBgAFwe5lF+W27t
fkzxFeOgg/KwN3SsaCTU8KntoVjYyeEm4Gwb3wiNEEhSEJRNPPUiJKOmUyC5a6sP
JBVW/E1yAalciXNyH1Zdcw==
`protect end_protected