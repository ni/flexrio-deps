`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2992 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
wcmpwSk7Xh2DEFViwcIwocn+IsGqsYMDVY/nyA0zXDqKMAGlPiXBLpMDMJP7gi4D
fpTyVlnAuqQ8Hz6T9RzaH/1lCSG7Ml61WEuaUhsB1F8u5A66s4dwoQZM5i0Q1gWZ
DtD1/ngt7+BCNBETUMq7OdG8Ejl2J+Kd95I1u8hHXeERUQ0yUjH6K7Xs70S+8nPW
xIBwZUTCGLyfpxlR/MAJDuTeumxaC0fz0iaXUSB4IC3Mg6HF/Juc5jRUus9ABIzK
g/RJp/38XsBKZjSCxFdWhDOXCn2UKn/7gVVNOrJeIi4LLGJ8YVl5QQzjw3ZFrO31
n1EdHOPnKgoBjQZa7PgZ5fiNe4ZIAF9vT91Wzav097iBiYxx0WEzb2dL8Wl3QtXK
BG156v5a8o6uhRzGBow3leil7mYyz+CdVMQyNJ7hLjjhgGeSF3OLDF0psT5RniXq
/tonvKhYcONRJPtiF3EpEynkJcxnCbjsxdp15qvXvt0qDRt4YuyngOstekrPnhvO
9B9N9Y7VZKJvxmLVHhUcuLHTMO9jww24nh6dwaluaS6R3S4Aw1BjZ52qA2tcOEDo
d5c9t4F6/XQb5ZHaBWrPZ2pCxeOM9LG00MfD+br5DOUTUiZvyzFiQMEUsxg0AHUa
2AvVgUSJIOdGyfS74KDYkHlLi1RLnwxVGQzf0nVvMQQkY3WfmtGvTrmPRjas+YGQ
Tu/rzduB6At/GWMczgcFO5O1UGUiQ6ZgsbodnNCviT329OBd/9gP9jMitz1XHc+h
7HVAJHVsjF+4jf19LGeiE5cnb3T0ChLNDhL50tq7a0pP+uv7ov+QJRNOLAZ1goqu
ZsWz0jUHn5MnX3YflCCQjZWi2Og+VWttmo4MPg6t01HGnEhEC6PK6eg7JHbLhXWs
LJQxzfE/kYhYza8skqCE+JhnqRPgNcOKzhjZ6Mqv/JHr3XTqT/IZzDGKZXx20yUJ
1VrquIC6sVM4HfsY9LzL0MXXGED/I+swN7zdMQSzOH9uUMOYlaoeqwRurJaGA7i6
ST3L1QS3Li1vit8MgpmK1t1Qq7fjqw6FjzWLmYCu4bB7qRCUBcYjPIV0ocoERPmj
0p8PIBBqk/aQphxyv8PJEKV5uQZ1lh+d8qrqTVaXUjV9jZcvF4MLklK0Qncrba4a
9zACmNqJ/j3ftvdONpztrfCBOcT5I/cm8f5kTXeUv3EVEXMmE+OU6FneIjQlcBuI
WH36rxKK07RlZcOkotEM1jvRA5b0rUaCkSji7gRY1QHrAoSPoXGOhjG+zw0upMTv
EgkTJjsKSpUZqTi5MdcFG+LGnx4YgFTWm29KdJW90anJwJ0+LGary5CuTZJdlfe3
krTYeLbyRS2f2QCzM11LVCRvieaPGHk2+uldq4gw1BBTCgEvAKRzvOfgsr0yA+WD
FLU8IRgW25GfoJuckrWWcqtI9sda24AdPZfVRKgn6s0SaMqJN09aalcEV0qijGg+
AGtTD58Diw668Z2++PbYw2IQstK9j3uDnwPPizqnUA7NZ0bj06iRs7P+kKSA+oFe
zq5IApPZOXRitZ1JL148yvAg4Xaj0bYqg887f8OzAmOU/2uLLxukpK1gViu4g48x
mjC9VePTpxf2KVAje+ophk8g0vLmxTh0MeGPsBFN3NqZgb6hwATl4Vu0oV6xL8qu
OnDniE5RqeOjxVAc9uVdh/g3qg6eNgAu1zABzVN8LDsgplybtVLM5nI13EVvlw5S
St0jFMUFuNjjHn8vvZv+JE8HsXbfkYywL9sOiAcKGMWUB6kDwydFRRfXY9SJiC0f
nwnp3rDhTyITP+EAphlNe27TFKNvUlwS++tlD3weES9yzj2Q0T9N9yahtl1KrIHj
614tnzhqRKZsHrhfBLthyIa+FxBnC3gka4ns1Ln3nAERlhsQ08OGgJSWKGtI2RZK
PNt2GFYoRZpYc1uBQm4NPIwAKEr/P0ve6uBlEmqRbQ4CZiMGgsd1FQZvejBEcxtx
2jeXyu/N0iXIZ7YA5HGUoxgOcL0ZCNYkxXzjzIZWtkCqj7wYhP+6WHP2h+zuc3xy
Flk8HNhRY/8ODeHuHdSrudrH5zIt0bZSRIjlmMS+rlVmKi31Bl1PuuYmteKyNsG2
73uvgHV0tkVeN7MN4lfXeTLUhYJBqXrIGWSEWuHGf7HzolRfp1V5nDDZH5sOC+Te
XpALQyFfHCGtrpdg6vBOuyTYujBAYrjixuH+bO0qQIdw/a0NRBOCtRrReLPYv5xM
zXMKWlkCb+VamI9OOvRp8NRWGv93wuLZlR5SaFdXgLEgptK/kwAV1VtNELFAxSAv
TdcnjebFC8z9V6mGhBMRAjGs17hjiO02OIp4SUeD80LG/ENl1PQC06RgMACi+6FC
BSIvXkIhqPB/vTCkTGRNuuBapFi843Tczt7VOUgZB1o17RuB1tVY361yr0L+Wb2I
fsDDO9000kSdHZe3j9lgI92Dr8e7GFxXgzxgKevq3Ln9FDtynRPzKfY/XwdEoD1P
avTOUaYsZiWTuuPnJ6PRWd9HMe6TwvxYur8jWHoKXsPTGsO4enboMlaQABrdebCD
I42wd14r78paPNNqVhDAP/tguSB3IgQeRcDZnJzNVKlu64BVAZ4OERs84oaTxk0/
e7lNxwRGvVcAS22D/JDQfbV13wf+vjm8UhPs+jzSPCEQydw6tkQgVXTXx8mHSh8H
jHheUQ81Opr6u6lFdJYt0YW1m5zkBtsl8L6SJgbSA3674JvqOiqQK6q7D+pPtwkI
pVLoPp92t+gFNCb6bfSvU2dW0jSeTgmFcMQwZPMY44B3cbJSqYmNVu6o8SiwziFe
qa+WIDlTrIKGIEJ0GwgOdCYqYiKU1avvUSXin2tibQMoLabb5YAc2nAoEN5KFedv
ERKmpeJfUYSj+ITrJU4S3R/sSCTaAEK9Hs9QFw/3X76nnENXXRWyU1KeyvLqnBMs
Ot7YAn64gJXReFKqLUH6QnNehxcI4WqBpFDcok50IfUDL3ZCAkwX5ExT8jRwzWsb
rlpCyDyCaA6RzO4jqOFD+G5xhEXTXbEtGCAeceO13F+YAHR9QVpqsb+xeLlgyePT
q7A+zDrVeCIz4tm4r5qcWryuWIDADMR8K/f6rEWdv0WH+Awi0qIKFWLEYctBswju
XauRlW11b5Rm6pnPbRbcT+gue52/qoGbvOclfLbI4QK8/CO9R2YfGEBFUG7hbkbe
6RuJgu622ENyT6ouelUV6etIsWQHPJMtTSitCHrhcMYHw34BrIVxTnGCfDuIyVso
9224S57Nmkeh7kOPZBoV3YbD+2xwL0vITpANTtYln/Yfx0eHqM2YJiGnXspZVU4R
MtFlrKanwleCWQx36H4eoEiibBtUFoW4cwS9zJRy8ufSlwxij08Glq4BgDrjZjwQ
/+4elArRywOfk6ABVBlm5QLSFWg7/pnbEaJUkw5ReRjRtu208IlvDgTtMay4JK45
Chi3IYTMYRyiyTJ1KuVCk/e2xjtpT6iv1uK+UOWxZeRDmQ4XKgAio1cLxaQNqeD3
Ps0lgFf+l6SoSrvOnBc9FkPEedhU+yuuGrBbOwwrrbpdQqmfyzOTpX55xN51Wy0J
Kq8ltkLdNbK0kntovnI9F+dE8HQlrbQaXhunuPEtCar/tMIeT4U+51CMA4cl2kn1
h6idHrvlf+9VoVRt3QDWNtXcIAOMF5+L/Ce1pgxBU/eW/hoTlfpOvyln2zdf9nlw
LouetGGB0BlzAungtCW54mTbWQIG00Sdgwky0Eo+Bfq5psRHhbh0UrMyXcGo6rXB
sfftM/6SnhbjowJU72eBXSMIoQ363F1nZnTpkYyTtxQlu8G9FMR3p8zdF3Lmp9Sg
bPMjU03bp47+lExxBCDubg==
`protect end_protected