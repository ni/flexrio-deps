`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aMReDmrPskJscpWYThVKVItA5gecPPZO1R595p0GoIq1TSTG+UxXhmmUXc+VYHJ3
u/C3EW5qePLufxmXxmhmDnr9U8/cYC1zLfk44v/2OPb1TBrTsludEDQZdGNWeV9l
cPUMSIfZ0dHXN7L1M1E2XtgoTWQxf3VDHs7B7lU2y9Rdm/ibz0fWMow7op2nWdD8
gJ4QlNl3f9Oiotp1p8vz9RFzzZOF5gBBslZxcTF5+z4qO2W7+xLByngthWm+exIr
3Pzy8qyUo/m2DDwOz3VJSvSNm7RUq+0/yJNOOz3jr3j7ZyCj5OqT/jDAWjJSMH+i
2402Un+wDMOQxi21JLo3cA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="5R6K2aWI3OdbT2A+sz4o9+2XAInTqB1/cSw5W16RnA4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
Gm/2BIZF5/H5qen8uQizPH9RftTuEE9mgEOF0SqeOKegtP64CfvEUnIxj/ahmIpA
6xUR2v2l7E5duaLZh39Mc1GYsfqE91NCPU5whLaBPg0UuX4cgTkO4cYbW/7yvcrd
4wavUfwXEp2VSiN7EVxL8RcZTSMSI0Jr/aojiilFqVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="TEmQtJ1Dsm7TOzpJk/CeTSSFx/zKExk04H6I8sT4Meg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
nvPqn26PC4XWLLQG0Fq8XsMTlhB4evbpiwGjZroFFLgtNlE6bBjdtwWsB89WW4j7
jNfYbKN4sBv0hDeMH0AAR+8g+TCqoX7yLdIUd7aGwBUZJr6FdDs2wTUxRkXFYNTL
V2foUCw8RCp/PMc5/qua/j3tB2/nhJYhWJDy9TTbv0mtQqxzNWgU3ex4nhw4hHTT
PWJa1MbcgkhmdSmqpPRo6o2TUNzhKwknUggV2JB+y+sOZSX5swWnp35tKsrs429Y
jM3yqRzBtRkTHXdR1mW/5M0VcMHGbsWdCeiLBJ+8NeYB4OGbHRHbaRqJ7ZBIPw67
mFNqXa4F9Zkyj+cMFTSYz3yXIPrRhIHfjKtflZheaxTcdmHF61A6mGzq76GIgdY2
wCuMJi6rvw4AE8jT5ot4Lb97EazLKq29pf4M67Jn/V91ef2Vg1c9t7etSBZe2zGB
5+N3sKhgDm3YRIwEoFsIGAIJedVs/L1o9EN64prpKwvr81UIMSMLFscvZv2z9WGW
5Hs1ubt7nEBiY73K29q6jV1znhCw7IsSwOwJHLuHWCq7JmCB0AqcIdo9OzMAaKIY
Hnv3n6jaCiWPz+L+QFgR3KS3yiY5/vjSoJIJbc7a1CEXdmeiWta1oJaK0y8OIjH/
vxNqo3xCplo4BtWmN/4FrKLSemARg+eDvJtT2SiP7cHPWb2aZU8NNEdb7U+M7mEn
85dozun7AgOCtFshwuU7yoqrb/LmaODJPvcxIwrwqgXM1KpuVPCB9Y3EXkLkuFhl
JpQZsZwVLfz4wgnOHXjhoC2A+WPGRqiBTdqOZVZCUEg3ij1Ez4LLdGrLhBiOvF4Z
2saxHfOYnmNplrgmAvGHdIVwjYAPCOKo/9tXIKztlpZc5qzPGF8vjrvZOLonnbEI
e0nYu7btBfeIETaksrNJ+y4CRgNI6xmOPGheRvU0z9h0zpvrq7keHr4z+shOVECd
dpPqVDVTmH4AF+g4QrQKjGgDlV+WLBTti103hJhPPuyeZWCkHQqC4u6KEzACSC+f
18u1bFxJGXwyDjFqNfYQh18zeptfJKRe2gd6BC1snxl4Q6oXXFdGtu9u8jIyeiEs
WjQfZ75keudJXSby+jszoRrDVswjiK7uBr9YgqaPtfEVdhi3Gg6bDoEHK5PhE+6l
1W49LyXBQVjU122GLvs1gd0VtGrpr41cto+2/GaMy0zln778XGDTwW7FEnRMWaFE
6H8VG+WgpJVjV+31WYGl02Fr6HaktexvMDxPMv1EMquFs6OlQ2n8hMu8x95+AauQ
0QhI224dDSfyWNyxUD0FxfE1a1AzG7Xhc9P13XzJnUzAgPRnyN0kKYUqaq6SdLGd
6TEhSssbjdWpy09pOLQDhnWMLzAwVeGLPvcK4NmaBM/KVFrcaV08Twtt9LH8xOqm
Je0rMJojGzdj1tG75tkw+4WIdT3rIPQv4Mfm9Qh6UAKdchakLWpPiAWUTRnBHtah
8YfcWg4JIAuPkbRI5MMCbT03n+oAstNyBQM5oQqyjO4xvgGQEKPeKvtJso+ZgMCE
kBiAz7EsjAopMVaF+TZWvR1cnZ/xZsweUAJUtkloDYpob977ih3D7BUtXXfdyQY7
iqAsfMcriwhifeDGNfuLliOi3pn+SLPHhMecF2hDyRAAaaXWhSA4BMAgKTV40T7d
w0/BOn8DPXZ29EZ/uS4XdHtquhwiNsA1apmeHIuVptM3Sc+EyRw01qFeY/DpajAt
yvTTFEPKsYSry4oUBXNYsJxCOrIjdWm3P/v+9lVmLPihr/WO3dG1WjBMUAPq5piB
jc5JeYXpulZ/zcg5hqGRtDAqccZyKz2Bw9nnbDyXZ2ALyyh5BIhhey0DyY+b2717
meH+D11WvcyFHCf4eP/sMBa1m98KCHbJfusNItyqcCBDjZMiORNRLwq8JdWx4IAk
QFgCPWeTFBGioCZuoFGKeJiuevrRNb85CApAtCZG7/rTy9UP0nLbcCq9AmKEEQao
Geu9MDqG2wIp9FiJBhyPR/QjmzD3l0Syz5qPpDvZBd0Kha7PKpGJ2xNd1sgbaK1h
wZI4M2H/eWBTaPNSTbiP4G203Enhv9Y8WKyaeXX7zXNtJY6OF3rAggWHnXj30JIG
xGnYIYpMbcb46uhRD0ZHsu3iWnGnzazbBsQm9nakLxWJRVNlrMC138lpj21/QWI5
yXYR6oyDe9CrwvQjlhCIdr61r9u/vngPyrdGedxWJbMf29GHTGH27tDoO3SCxuoW
FxuIPBPi4SOVS15L1ZJEK+GUxnTexItvIu/UHAHESCAnRG5cMhfO2x6KCrBVh1oA
jd281Y1m1/KzpvF1SGL0EiEAead12Wu6RkFW3VvHZm3OvjNIx5Y/Cvqbyq1AC8iw
YslIdqfIaWeB6exKaQ7eDoX5Uc5rahzYt5gyvhJcXfG0nkWweS4jClOpDl+Eg2cJ
aQZoy9Rl42fUPHRxKR+RcGO8E0W7c4Fs9S113+qoP4p4lukqSjKX0tWtXIC3lhIB
uqDHA4R7sB7PzAL0PcwBOGXjMXcZtNy5dlI1OujRFZryxGDzGl79SvDpMWoTY0y6
nk0yh/zeoGV/Ew1Udys/bVx80ncB0FsJIq/YToFH2i08PMQ11hXJoduI9n5waHSf
mCok8YuVzw3WwT4TlIPpiSei0nlHzlFgeEaXlYHrixgXlfKA7D4nZJJOsd/tJNuV
`protect end_protected