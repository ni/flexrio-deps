`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
rC6KPz1bEhpOMfeLdNDaqFWs22wvhtVsPMaLmxfCFPgk3fk0DvFSGCUF0a87ceer
E57jVQ8s9FWnCZiHv7LMsu+kGBUm695j66mHRxrNzB7Am3pHg+Hgj/glROGquQgI
+23Qa1oLAuy1Q++3zXgolhKBuUhWa6G5HxtcARBk6M7dy05HkUbjibHUjCEep+jq
xxaMzhJXgx73yKhQ7YQPWyiQNu/bvI5VqqfL8He6FiblNNej1Qo4D/yKu5znsU5E
ZXRCVJ+dx45fH9J6Wt/zUiFHQ4X9lw7eDzK9tmSzdssz50Xkh3GS7r+reDEUaMVC
g3m6gIskgGnadle9SyrWaOP2jy/J/7qjeYKrAT2PS57PnEFj1JyEiv26rsSW1KEV
l3wa3lkXjevZktFXfxHtYn/CHQCYd60UeWLiBN1Mv3jm+XRWwiFHYPjlO/NpIDwr
XNB/IF4c+8H2PIQooN2cYkW3r/gxLBA9KU01fM6WW/P94Vhcbn/4h6tOlXBpnfc+
Wt8AsV4EVDY9TS7YTNgOs7l80ccHEMCZHCveQqRxp0P++T0EduDXydnSkR70825h
YvGzyo/GAlO6NfbvpOTBUCVFXbBGkRQDbHp6NYg/yKYWW+Sg+66N8slIpFaRDqUz
CmSyUrobortEGKpkydG+xdt+HTla5K91NjgL3YHEgksujCREGnIbPi6i2G3Ui4jc
Jg9Q6mf92jmX1PlH1Wxyd2fMrDxx42nB7OnAqlCdJQHa807Ex3eWOHDsaMYNdkUY
g4MpBNtX+ve8sD6+RPs7Ru9S5MQkL4Vqsp3Z9KRjc2A42mYF7XLjgJozrKJ7GnNu
1KNdsDrG79ihckbK4jHQY0cku5a5sRf1OKg5hR2sck60/4hyJv4ATxgPXh/rlNNo
2s4DoYp1vRjt3Sw25deAyibbfZ4K5KNk4TzqtV0LFKmyWoanwRp/vfkZW3YWflmV
K68NAekMi7gRG5fF2/AZaCGcKgo6CP6kNv7hv1IryAWcv+RyXU3N4mK9UvNmtRMp
TIpffqJ3og9RkNdidy2143cwNzvCdgZ8i6xO+MnUvf5BsTaJzfkfMM/ebM0o360m
ksvO9Jx59ITk05wbY8cC4U7kLOoYbsHV+eE41yukU8qLY6QWYcuOg8zcX1bZotrf
Z+kIp535heTtyRPMm40C87hBnvpXcUM65MEp0xyoV9ZblCZhBVfn/MTziYSdCcCB
cH00c9HXLBGAV5m6ilRvpU23kbr261U2aBorYdJnI0Fb4xFoz5pr/aqPLbRFBJ2X
r84jcolLOOMUDz7pRfGh88oO5lxxcNqatSDAjhErU+z9Eb07angOqUx02fyPFR9T
Fm/TyWPLKJtcMaUHPLBWn2aQ15i3aP8xqLiHgoHDCMwT6A3x8HQLmWVCjBn0E4xL
/8oGzhNuzmy83WiOo0C50Z3/xjixs1Nq72/Hc46eITsQtrTxjILdYkHXjP79slbF
97nE9YxWVOgjriMqYDjuLNxP8pX1SWVlk34DRoBMalMYP4ZBZmcxYSFESeaL2MUM
xnu24QiJCUcUBPi6WYk/3P3NZ9E7A06oxOJtRmKa5oqX3OkNKGqKmLxIjUwHXIoO
UnvNRbe6o9TK+rx4VSr86KS6dcyLMVqdNWA4xqF7MVQcTeQzJ8T4TXI/4+T/BhOF
A7x7Fe7bLojD/ZvRU4VmVIGR/x+ZZRRYWXILsiluhZ1pAK/Dk/yGfrXBs8E3jRbS
q873kaXkjiHc7iA+TvxVuatQ9ScLuqrTOS+NUHGRQwB7fARm5bFw8ypGvJH9uNhL
QfLM7ZnJdwyuZn9ZOWPT0gzf0dvR3nkR8VBXZ9tGWQla/yJMfZZY3QbGH56FMF1k
bA+6AATgih7jA8BaFsNObiIMBUe/CXdX2jj1ZUmzLnMokIgxGkwfmRw/QoEiTSkm
NaQmR67QnibRJ8GOewYpCRxwp6q3VcXjAvRiAOMMP2NHnipd3s0Q1iG5Apn0JYKO
4gFzMLD01azjnUSWHKpZnAfIVYxpCbT/mw0Yzpy5y28xHEkP24TIo4V/v7TCakdX
rWqM9AAPoNu+MGchY04UuErTx/EDtc7BkJ0RgoHx+epxLfB/BHu3HUs7B3Hgy4Sq
w063mcObGN810vVbjv6rc55ufpZENipODYaMpqG51bERt3y9dvowXpn0g1Jes4WK
btBkqtivbKYTYtU3Bk3Y9AWNZJp2JUOQOibKmXG47LSdyykMvCU+MMeBXULUZUQb
fuQ9DDCSX5ww7STW/RaK3QhTmJdDLoGswQYOCDxE63QD4pnG+8E1VMmCk1FCdZ/1
Cwxf9/S59808BY6uazmwGTOFityN0Zsl1V/vOygqrcSx+H2ziZYLHMiZx0aMogjp
lqAvrWXCC98uBrvvIzhhrhwWC5q0djQq+Eh3RbJURKliiBLMcepQp4UnHC9IW3Ic
nB7yrCdv1y9FJFRBn2vt37+Ty9xTDr+oa0uu3sBQMqsHDYLPeYCipoQt/ZFgYSL2
G1+7svTPOfGy5GHpm5OsQTSGfH8Zy/v1ncdNUw2HX0HiKSYcDkB2ICGWFM8dbReG
sTkj/rGZ09FHW0YnJ8KEvkT2iiQDcMqubQPrN2/xHfgMAQs2UFYU02keOQJhUWfQ
9R1EHT645qHz8hirSvOmeqQo8YoALfwfxNEyB2ywhfg1LJxoZbBAadIh1FajY3Zt
ARU4wTWYj6EuNwDLHHEu01XOhMLGPX0OoxHhZupEUEnpsj3JBnkd1HBcP6rayFyv
o456TVvz2IbBh0pd4AzFQFcLQz8hN/uUgYdu0Ldm/OPg4TMSkKdkH7Sb3u02PfgX
TcjLWsTazpX3lOC/gnSNvtYetNtcYwgsKpt/g2QFq19NEoAYqFkt5X4p9ZtgdCV2
C8b4tEcB+FyE4Z+Sj6M6ZTg+dGz81WRPK2lX3pcNbMnPk6QOFdcBeQQAylkrOeBC
oNsdBt3sjzOJwQnwCDlS7URE/KlmvJYQIdEXHBP0BXX0m4TY5y+J0bZOD6mDLj38
axIhvob3s0JIBXRa3i6dX12N6b3XOvv3jxDCzZf3NFlnanTmSdkFXpApZUGHdR5F
6IX7yok3dfHfIz8gkok3lOK78L6Xgd78gtNH7qyFQVnP3QvXDhhqTPbncB8BgUMk
G2Zz7AsCA7preCMWbdccwTMEPk0RCct/WvP0bUKUsvx5dG4rMYjQe3TWr/SIdE6/
ToIwKZ9qCGEvd88VJBiscZt8JD2NfLXy9898yVjRIOslnlufBl9SNJIJWXBSgodA
b0p5ggFYA0x1iQIAOEtlKfFl3EYouaDg2fqrFFIpTV94f3uCq6k5j2nYk0eSdF/N
PpzycE1OMFg7WHm0sm6WGqqAKw7PyMCcIgIGQmOIilxjUv5k8fzDEFFQHAEakL/W
dDp2kNZsaVH/j6f+oY1Wzu0zKpR1R+3is9axi4XNPok/SSo8gvOuGfGIuKvT4dI3
kaa/LnB2S5PQU0lSv1mVl+YeWQm/mnZuCqi8Yhl3QHHeWmgFaCnOdGZAbCw8Gqdx
HrYkT93yVhvHobUe9WqIH3Q6aQNRH5A3LEoktZ9ZB+v1tLPU9fG6aZ0LijuO8cbL
XesGARpqufvd3MdOQiLrqlflNcEzvWNoMUe2QA1Ci0L7atxI93zP73srk67Dw3jz
+QSYJXzMJSQpRgZSOtoz2jnz4ZF2Qqijjl7+3FoVXv05nepQ5Gf0KLzciLte/o3c
v3gmbtPaB9wW/rmX/VrLkPZN8C3FCIenytBMrQGc4inpLTP/rX9P7uLb7oQhg5CF
qQu1CJvLJ68l0CtV4r9CxdkbSqdmZivGg0YVtPTcdqUa2g32wPcPcX8jklg4hxPQ
cdXEKS10NfN6ZVZvlGhizXsvDOXHmHrdvp5lOt0yS2i/mROyqJ57SjIeGUKTmZNR
KGTtsHfQOLEFgtV8JtnCPhSg4lzTRob1c6igZtabv1wIPFJ+t7x6CkfW0s9UT6jG
MN1Hgg9hSxI4IN09tLXECenuefJf3UBfbhBxmbTryAr69Rc7FJfiTsp2Y+4TTU4o
imdcWA8ojnVPrZnEvRow7taMrmVm8BTF5EJ0KOoBviSUjcDwQx/Z4npMsW2Q53DV
kRyoRt1HfRTyucMuHJm16T5vtCZzVXGilCPID5+luOMR94Lh/ohlNPozBGl0D57Q
7CEOSuAXrbKf9yngiFdMk3tO2v2G7CAFFV+1JemYyUiim/CNeOZg5kZwtuY+XzIe
JFJq/yc3c9HIPqzeREzVCqqS+SwtQkgg8BpfxvuwQkBXGKc9WfjVfJAyO0uQn6du
S+x8bemwK2uIWbDCYnKFgvuiuYMV0CEMwRfZHhDKaMfNS31Hjo2e0F/gkQ7Jj9sa
C6ADnRdU76/A6tJUFh3ye6hhHusXq6qgyO3ojoZuQT7Rn+v4ZYKonh2HWQLtaTgX
5Wdq+nQd43OSMKB9njtymevaMTi3gsRRdffclTbyAVSkynX7+lbRhz6DqXwBL7t3
tcTjkW8WsC01j0XF522adxXHtvaZ0cR96/GfK3ygsT5+vrf3BQKmurE8xhHhUvfT
NWPcsMuQW8gCXbIiKK5zL+IuNiMqySk/mvH8E8kWr19/w3lgNZKg77ymnsxr76fo
vhKa0aWTE6GhUugU/phMDQnOb96y/x76YWIx8NS/jds4opMOc64ReunWES/RNlSW
bhYwQwWtpBoYF7suDQR3amuLhSdjOUH+ONWx+0dMiq88h1J4pD7lBw+73g84Qjy5
6raK3fYAdHaNtjXwPsLLx9qx+xcey/R58fR5HNfsv02HrZ1LLtRT5QYsdOCfXETx
EsUn/tJHUo3z58YZNelhLnlEVE7Wr5mLzugZiE0ml8bKDjCJQ8fNCl04ebGgyRIo
9DYRmWAPAx1NtF9Sa9i4jlgY3s4n17XSIIUWbSo0tztNR60Qdb4Tv5xttItGl1RW
zdw/0zmUs3aLSOlMOJNScMGkXFz5xbEmmla156VFVnXxbnh1ziZOu/r4iMmZdPfZ
xKwQO4I/9vqNA9hOm9cadbfYD2NZ4zqOMAoPcIwVD+pDLwmW9pAri3y9JUBnBcbc
r6lvcHu86A9pdIckLMSVsi4RGWE0Pg5mYGjxaEFmVYcG+02431DJS6k6EMfGaU+k
AENq/nSA0tF88PqtNRHqJ6rL3Y6xTvVFPQbpyMlC+/FyCz+EPqVMUg96WjUXoGAK
9ySRIbpuSUK53QDZJJKjUcpUdf42zenw8eTVgpp/hGIzaHxxqKyy3c6qf65p2Hj6
rn7eoTBxNvdcWyPYUYVZmG07CIHMLiGR0tnaYupSMfwLjzZjsYsU6bbOe3Sg7hUv
LjyrBBpkPaSuXUZBiHFWjRRWLtE4DAGMdphQUAKn21AZ/bB1ysmqCPE0V4FjKwLr
Gwj4f1tv8VoKzI84q41+5I+0nJGLVTCta7SKo830xp6CIbUWw/2Lc55Zqkm5tp4y
HM2HI/QLpuna2iCZbXREhMfnmp/Q05hH6JTiCWHR36hJDZ91g0a4Euz80pTNO+ur
5eJCnL3QhsZJJqG+cdz9D2z4xqGJf3zYJ3SuGJIiPKJxZ3ET0rqKZzNnpHhEL095
DjNJllc0cOpDexCE5cR+38y6U+6o8lBCE14XkIWTmSuK2heLQrFcGztCLsO+b72C
jbgl8/upWluaz0w6ivrERL6dNHIhXjacG3fVzn4Fi50PHwcIh09iI+9YVZNfGRsv
1mYGgVKiZm2jHtNwaQEFtT508BZyScP+R8qEqLZDnvA3PbKQgL+2/rvH/B64nMgx
iX/Kod/2m5hGOS3ZyovV5Dp9d1MpF9pyPiSDG+pkrTnFi+cjdoKR2+MHc0T5OZ46
3LL8httR35ym+BIpr3w8tvzSu52CvBgsd9nfynAEFrAlBAYB3hPyhJEJqSfcFBQa
0/q4SUBHZhxnQMMFcsEQVTFYo4IOnw+bYz/5AwIz9XgcHMT3MF5agZ15bw+hZigY
UJdKnp+4mIrAv81d0RWeMWuTPswdubIuQ1H6JNanIgYuAB5LBXxxaSoeJSr0NVWq
GZ9aeUwgnlu5/QCavHubRZXkCnd9c4nGycqjnVWBSjK2rPB2cKlgRY6TWjVxA7H/
MMs6Zt/WWY8RnsuN69I00qPJua5HCe7nnMWGdw/tN9OPwU/KoM9ik52+CECwU731
9Y4nZmkiD7WF3OzVkbXRrx8HJjJFwXbru0Dva9IAFh5paOZp5LIKIAVky3Dub7Jl
zO9iT0yMuIP8syAPoq/gEWAbj2JVYY01fvTuQO+m3o8jp7LyjmUj8I9oIj1WnN3K
Gbq8Yh2wL29+0dvN/47tmwCoQie3y85z7Z/vA6m2ctM+TgAxjvH8kIURLmMaNKxh
6dq1VH85IEdCYlZNqatRzrrcTVwkkHWqNfIgbkmo23TcGfrkHYKyMws0veoy8Nbn
DQpjFHf4O+S3IWVEFNHZtyvvOwRL6GFBiCGvg9Y7zIeWN7NR8cUbkamWfZy+zGQT
iA9EB4vIDMQ6ipb1vLOsBXnqXb0g2UjumZaVCbIBkw5TR8hx3nVSFRVa/EwPNN3a
i4I0aW4kXGM2hsl6pZd7W4lQjJWj/JsXPVeXHfLsBpWKcWTqT6bbCyWQpeIaohtO
KbJZphD9gryeA7RZ7/TprRH5qa4aUJCyOGfr8kcvM+VJbOBEE2gZy59hwbHuyr7r
H5dhV0Lc329eaj6NplR/QO8c2OW9/sKwkoMIru9TOeGjhu1O65+c8/2kfK+w7mIA
mXUODtx5T24BCPiHtZvzsezxrtMQ0F3a1c0WXVCREoETF2fenNePYeZsTKlXETg1
OcqbrsIgRdNPiu2u/FkjxiOhVGbrFJ6aMo1wWYZhLuBXRk6JLhcMtnb3Mrg+KU9w
QUx1Cap+SIUHKcAZPs2Q73PhLfiwOm9XDDq72vEneZTRixAuv3iwljw4wi7ju1rt
2T1oNZAyEXZ7y46YKVPmwgvsGFGUaWUy+pxvjgHHDCSs1dlkCXh1yLL71XE8U2x1
JHg4+LrLWiqQz/3d7kHrvbBHnSBlA70UoTaAOc6mgh6rRO1Rj4m26virYTXbcocj
xTJJwmMZfAGQYaTnatedXuyBet7rCM5tPD+LBY6gjiay4VBVV9Y+JkbHzDNJpgh3
WnjQV9IMXRSw9gz9nFEoIe/bjFtgw12IJ0d9xlbxkM/k3LwNAHMnaI0kLwKw2Ild
usAbTE2E9YDeNGCfzbOUBGm6G0AHKykv86ryKeIOv15fD77qVRZymWhSFFV2nKzj
T6alnFIGCHSQRJqhOTS7InGTUPT5fKUU0Z+OG88Yg8uUPeQTuXgVJ67e/Iv06tlu
nL+0m8nG+62aFvq519BXL1MVGwh+3fjPalHEptGCJ0Xz4ey6FoH4lwa+LmBRIWeS
KIreR/smzOrdCBaoBle/tRgn1QtMYnI2n03/QSwLfhijFPObqxNtyxMFViDWH8ud
/g6KD1Y20IAOBhddZ6O4R36rUzLXXsa3XMv12pmUKjYAuWTbX9s7qQdfhqFvy1u6
whiK4D489OYFtsZMvF0mnvEsVK6khrmKLp+qWsSMYsfTyFS7pewv3zLyRCYTjnB+
jGn3qi+9CRxAZ/tV9qh4IDFkrG5lFLgFlSbiS9sSHS7kfpSenOz4UGOJYOZkVY7n
UVgpCL8WwJtPaqiJe59Pg1FDLI6s66pcAuuOmzfuGSBmtfz/UJdBJT2N4xY59lZg
3lWArpm9wkTX/F569reVyp4Fg6NAy/7yLqtcHqdd28+KKp8aHprikxB5fJ0ZTL9m
gfEAWdfKLucgWG7p0PtEaQJju96XD5Dc0+fHGKXrvSuNfy1maNJ5N0mz92OrVsCH
i7dGMQIyZ+LGMsnyRuiblRsHMvdtDN6E0pKjQsHKK91VY9lqPJ6/Atc7f32l5A6q
gK/1hkwtjiZKhsRci8EZitQUNp7sLe8ggJCKaBIOtjUvqifZoeRbKWLRrhDNFhy2
Pw6v9c8vL9llyz2gYHOZLKNBMpmFcvijUCaGlBEKzWNsv838Bm0QajLbX1wNU02M
xL8C+TFUG7yNfpV+ROolXRQYiISQEcoDZlHU0XbZdb+OG8vouSUWA1u8xeUfr95s
zFZuManHB3OYCEfT7HhiSLVa1ij94j+ugz9KFibylLFPGNIbdTKCO0a2KO90VZ1l
yonKHyA98+CbL7yvQg5mtZwJMHggAanmJzYWJi4QWZO1qm7paKxPk++FQ+sXaEwR
viTRI/shcPUgNxHPRGPCNKjSkZgKhz8fUbzFs7zqKakzd7ynnDyN2nlYhtfOPbq9
Hu+KY/jmrHw7Ie71zro9wAC999scb7C7T6/K2KfyLRQ3PHQUvs5Bfi8/7YIn2BJN
8M73ayntV6PDZC0ywXO/RL276M0nLr/8C/wxOvlS1tbG1hzcsgbNJMX9HC7oJvYK
STGI++QxxZbgqitbNlOjcQs+/QUtIX8SQJAXeHd601QQfdXBynWBIxkBKEvydfPG
fF15N7ndjuJel7OdzZGhaq7LSIgptBsSWOjix9dSigJ83nV8QpaRUqq47BbM88W4
+XP0j3utYfK4SnyE83K/x0L+HqE4C91JCqCSLgiZakj28oYDs6V7yV63bEIssae4
SmOo0Yo1JFArWQl0oZCDpzem8bSGMSW/1WwLKwhkNPa/tvL3Lfijc+/p3xGs61YC
b2XnMNvUBWDodPjYxHtG7sHYrx3H3PvJtbn+3Gztq8oEdpsCYqNS8E8x5TnQDRvA
O5czoZ50SCdCGMhMVrsay6fRxTbVg0yVZFyo1jj8Rwje2bAVyPj2eckFO8HoTGxd
cWVbEW7VTyChPbY9xScD5g6zLmNN2cEAfdSlivZdBhRP+Vyj3UMks0joMULM9EMu
HweB6Gs9MCWL7nVldjwGOVmngC1c6p4AvCGHpKwi0IpvcKqfhBnpFoHCvFWN3dWO
eibCXPdJu6pvpcF5z/7ViOpOJWM2bDvWdpYfSAlemLyOXHsrynl5G84gXOc29RM4
BL2gfXhniGgLDoS//PSTAqzXI1sVB+3SEg0K1nRwy3ZDESnI2ba+zAd3yvLfYpkj
bluQCNfRpHrzKVLUTyqD+Bi3Jgy5rhYKxEHMNFjajNJIcQ5BmnuxfLYGqYNaDdgw
ZV74wmHa5hbHH7zXq1UeiSx30GzUFWchMkA7+G7njY2sAWBCa/JoB5TKKjaWzeYB
BNSdZFIHaI9LyJIhsV51QN+W5q9G9aqW1TQaxP5jOcAck+mIp9ZvTCchcCVmeiQ6
xccf2gDYRSwyWy6Bp7eQG13nAWlwGaXZ02NQ+kWpWt+M5D4um8pdRYNUYaC+6tI9
eDUsjgqemSxIHPQbOwO8qvz8eB/dv1l8JDcJuGOnm7a87Ll+VwxBlbLSXiQk9iHU
bZZIxsgdN0j/qe9dUnrO5ua1PqXnI6901TtAVlrgC/BwaNxGtly+jcS4T2WR4iXM
OH/G8RvcoILZAgl74qWGjcD88LncBdv6ARfz3esfdCayYjTqfP0dG6oH8CZyPNG4
Xqt/DzBamws71J5tCdwQgPTCs8TxL7KTOegfLe6Q2U3kVmLYLKpB14gSHqsmOSDu
YVo3UjyXw4ABQ3tb2jNa6SnF/VxL2zWTDomjygMBRtyRYES41LBzNENh6FW13BHr
AtV+RVW3QG2R0t/tLx8ENU8FfkGTsDBCByyOqxfaHqE2qbW1Q09PMd9UKUG3xajf
rfg+i/xHXQbLP9DYQQzrNLeAlfXeC7XPx1apMeEZTkcn7tWbg6QHbO8pBS1Y2Ac5
R+8RQ927DGiO+PJ65V3I77QhG3O3NdC4wtcMR4lra8Dp8a8D/6wEBZBT12AjesXM
EI9RCBwT4sRmn5u2HThQ/9FRe2VRAO3eg3k1cfXXGg73/DH/xAVbA/YnBenpKoXc
6mXZUFfdBIKiOsjwxiH6TufuztDYadUMnqNQZgiaxwnmOxi7IQ3M3MWwHfEp4KUe
3mypVPSMFM8GA0J2oDhevrUW+oSO5inb8tclfiClt032GGq1ZZI2MMhNBIJihJXN
ZYG4BpAM0e7jN2FGccH+FsZHU0Yll1sUEkItwJcNsOwrzBq8JL/+D+eSRrphFC6n
UvRpjryBLjNNS7z7BQG8SbEMhEqQLr5qoTI4MmaWPqroX52Ov73GmOBASoVprMD2
dPUGJ/JJ3pXbjWMcN3TDnXFLsq+o/y18UOvJBcKwb+06UVtPPKFerREN6/EpKNMI
FqM+CEcwvkpQd4ZkL6YR3bUVZK9+VG0yL3AujsKN9y4TY1q2eBq81HTUI2C4ZKhh
VMoKZJGVWJSxVfZ38KQTV/xK4ch5faRoHes7TatQh2rAunfrPqDBThrxK8/uDlch
qZmGczLJJ1/6vCZuBzU9eLbefC46MqAkolIm1br4E4eFzdHWGuvgxT7tpb2d4X2l
ME8M12A+Tl2gXD7+ozqgi7BJ/FpzmLak1qhu7JMoL/i82A0Buhse67n9Str5KbUG
iNZw6EwNge267b0LvKnHK3ae1/2YZOOSMW29hK/skP/Qts/DughH8mmqTEthunXo
UGO/8iMkw6JteJ+7EceCRU3SLbl/lj005BGTA4UIvhceC6Zs1Gl4Zs0VCtPLFCxd
zE8XExJqGgArvh4XfwU/ELiOlXxq28p22bJ6A0cdQrWryFBNXIeWtay+DsivxofT
e6pwKnYkSSmQ8ONje+Fd9PB5e3ObQhg6SjSrrY6XbjizKEPYEja2AOUPjkCkcGNH
daeciJjxElzzT5AjJO+H4Rz2msOekgqhLc6bDTlPoH/+/PtYeTGk9azLwuz5/KNy
fqOmL7mw7VkcLzNmb+ygSX81xOMtxnv6LMuFobTin/570yGE2Mrq6kz8kC+JyVsX
ghAFVzCNkSchLyLVdOVabqWnicbEVKctbBGN/sg4QWiAYRoT050SFMbbNYeui3DM
sRSZMMCxnOHK+5xAXNouZ8h5EfKArS7qXBYwz2dWMenJHunVTgyXEO/+O1k4LpuO
h88YMFbA/2TUpe8t0YizctPy4OV2qvSrtN3WfphaP0nEgjzgUx+nmgcabMMQZWfl
TKcEf/IOi/7HRdvxoL2sqwJ9Yfwe+o2+cBNaqFM4q3CxQbIelFtCXjfdIHyzbcrZ
RsjDJu1kfjsSPn/o/tWCwveefCpEyZ+7VNPMZIu6LpHFfflDYPQUBVTSZ8YtrXDs
K31fvIBZDgw2LMRlwGuCKh4/9CppJU7Pa0q1M3uXG5TgMijZkoy/K6sn7rx/lL+x
55fatlhda+ZXLEB+TQXUPOaVMAM0FoFPHEE4M4aiPPZIeHvOe93d8kwAiqgUsFv2
UFjWdALbUctbWspcZ8QjoeuU+TS4yD85Ujid2RNrtl9CSR0cWR4xLL4DfUvseeiu
es7cQio7hEMdBHrf70Cda01HwUmBdRvF+Z3lqsfGjx3eaxXeR56q3GzI8Bf178Vy
v/O7BC94zHwW+2jVH70RB5S5hLEnXMWxi9g41lumDJ5iZ/ngFgkjkgDPH8VLFwi6
XHX39kHTnd+j6erlmhusprMvKZtZedBh/7QPvnLkS3Bjkj5wP50oin0ZhJ/R2qmM
didH0GVs75ev5slt5VnpIPilSMJWihaFCC9m/jn+4ZUyevFKMrjoJBI1y+a2XcWy
ieDkha/t0eeJtIQFBe4ZWZQUq7teWqovW8od/slQqBfGXcKLlkc5hj1NU3+d0tJ4
wfQrEZfPHGm7oJSjSCJqt4HyWTsXZQQ3PFyEQeHjM7yMgsNp/eXjnepp+jQaHINx
dTwRkQO5PEJhfcAPqb7FZaELmgoemh2bVicTrmyvIWXx0DB6MemXZHu0PfRFfQZ1
kp6OF+LqOvowfGzumA7CyD9RFOp/A/pe8MaBMcPM2dnedwoEwrgEuFqpyrWctspS
ExgZDKqQ3rKQBMZm6wwzwmmu/C1zTDyXDOJ8nXRRy/KViCIFP8cgTkuooMsDytpU
pFNY/NU7Bw59RH9YfP1QhekOMp3nbf1yFvWDeM4dpTjVc08bqGcde4p2JbG2OqP9
m/JFBYALdgybqOEbD6v7Ku6Khc0JSvwEWheo3lo0ViNHKLEbyQ3K8Nq0gytudylW
eRUoTDzuNumNt4LXzvHfewBNl+GkWIi1qQUluoQtIJLmujLfDtI3e1R/m+iye8Gw
LAGT/C5HMvEMGVBpaPwYcgLWOZTOiYtfVhrlkNKAFVZ+7bpXMW6wMyrxX+qcKIPf
utjfj1XeWRjzztrJMrNAP7s1GZ2XPN+HoVALwr+WQ12D9dhlv0kGhi6KyGP4/M+U
1eKKpVKlaojgw5sUG+VW/iXr0Ior/3o5mBX6H37FQM+3XJKCgkrXFCQ0y97PNbUV
nk1yGVbuPR2jqiHfxA4h+3cZRjck9+czBQTeKg3mjGEvq3ht4R5jUaMNITxKpdUE
8+MFD9tYjDSwAN7JRm99sml2N2sE67quMm87TpgewaeXzROU701dwJ7TozJoHbZ2
hAqDVnn2RplzrK5ssd6n8e9AJ7bVlM6n1NfdS+BzwFvFStBw6IMVbvQDlBsZrYc8
si+QYVhsDL8ibT40REWpvYImCe3m8aAYwRvT9tYnr99bRu5tqrv5u4IHMLW5QLTd
5WFU3jeIdC7lbO5nU55VE2WmfPjeYxp/VbwofbTXfVkKBBpX/tZhrXTyQemrpEVi
48BcLFb+Ccbodom4Hmt5tNPdkbfsrXyr/ZTAths4KShXJSjroqkJLZJLCchNYhri
96LPV/AxhHzucu1TEgV3p53g3ewOTrbjjFVKiwH/bnOOBt46ZXfMMLWYP+VGbqy6
BAJtu8wWNiOrgI2cN5ejs9dx6r8J/JtgLUJVBUH4hzW7YTET7DUH1LSPJZGL0ZhT
twLpXQSP8K0YhKhw6pEGVqnncqF52teuxfbi+3RAU+fMyQQSI8A+n4drkKbmv1Tk
gD4Nr/RLmM6SKaYWhHjGB9GNgk6FocQFwUvm6m9gvKB/x8OV4uypcFb4PbAyXZpu
Imf9WZQgLA2JOt9nRKyMPuG2rZ4bZoCE0MpEsCrXMouir01weylLZKMBnyxCVlaE
GZ7TrTD+l/N+qQc8YaZVCXjtWFKknj7kK5fnrdZcJrXLsyHwZ2cxVKrKEc4mBKTy
x3tHmYID4ugqtBLknB+sUml33kxPe7MlnHg7ArimCZL7Syzla9L8X5a2zJusDJnk
yLxMM32p4o99tozAf3yar5PqUuJXFJuZIekSAqhGQzayUXqAaycFsjClJTVjejYW
9e/VBr49rBjqGqmk49CIrTnY3pA978o04M5tQSYWn8xuIzMIUbk6mCL0PFJFcM9G
7SWF7SvAOQNuTViN91yc1QLXQID5bAKKlcPkCh+wruV74LHHaJ7yuq93nf3l49W7
uDvriN00sQKpDlcxMAIRArSB7gv8C+1RWlYvP8404QFcRc7TYLfQWEzVTtHp2GhC
hV3dvcUhO5mUh3LnTKwSq0plMSll+hQuIG5ZR1bFPIuEQD7ybtbvqcqa5tpGWR3O
fDJ41NmhOue441ix04cmzmX3kpbWELYsJz7WXG8le35XJJYirg6v5xE4Ok2mN/Ph
YjAPCHKXSDCxuj68ZNvY+Ez5g4IRT7myO9l9WLldklTmAMznSjZYH2htfBASa+OL
RDrDN5iopEizOXt4noW+QWn7SeP9IFLUMBrZBgV6tov6UrfNy8KBWnHtM8fMPya5
ki+lfWkhlcUoE9n5vDY+IomVPr5iMuf+dg3QJsgC1wZHP73RoiYpfntWf2/9KnTN
Nx2eOv16w1t1e8eUTt0VbnPq1RNvfLEukxwYAjm84ncXbvvx2Df2EZUBy0X2JWlk
LKJjWZsbFW6RX699C2qujDfP0rwn+1oDbYw1kulnQC8DufEiGZrF2+cIogFkbbBP
e4wwB6zSf0K4xEx+olg0l2EeVHUG27CcGPrnBSe6Irgl92auptJw64g0tNc2l+pC
iDiHV1o/0F8/cCqlxB1WBpEVXAjrdlI1xzHd2KljWVViRmfy8O6QS0mSRgpHWQsI
hdxvIk2p9VlyTkzpAII3qOiSxuE+tUXtIpsVLL82nsVBTq7OLwitpETQMJu5T2mU
K9Wk2NMMyLpKPvZjOZRTNOEWCGJCpv2Imbp61R3qWxhSwCSa+gyhWLzwWu5d0mza
NFSkRkoB/IByk2aTStdiDBKcTh5gGi8E342Nvr3/SE6I2DHBjL/W6dwkWvU9EYRP
71o0lYwAh3ON5ljvZu1oOfr+9vCWY8OIEzIK51EdIxvsx35D/Yap+j0AQ3nllsg7
+DClDK4eX1AZNhaPaGi4vn1+gNzWsuvTw7TdgM3wWT1KRAK6E01NX+yN7l0UWOVm
nJLVA1fDcvxyli7MgexZUS8seyv1EukG6TUBz8lTPl9k/LKwp+FjFT3J9tEMCB4b
DGYJ32d7q5G+6dcbTeup54+x0nXgkKR5YLyKaZtJuyzioVMStu8KofxXqlE1lgem
A6fUYzuuoO/lPNxJcN/BOCLQJuQwKj1QZdphYGVk2xjvC83RI/7HqIDcPiTbgFjn
orKQ5NIGJUwzdeR1dDTUViAYGdrpnpxJmmQUmA8x7nSB0nqBod+WhHZm7uBP0D1b
PYdHFaDU/4j1mv5DVRt38g/q/Yxf/1MFfmbCGRuTGbBkxYG/S1j43IBycN+7+FPN
UopJ/fewWPwNieHCeGv1ppkWiP2I5NaVNboKy+UWU6tJ09SWKAMpoFQaDGvu1ULt
Gdp/O/sZ8UG8BYD2Q3WK7EMaUHsEYqwO//Tl+ehJ8t0AYn7Nt/rSH7ijQP6U32l8
SWb8j+JM8mNM9E534+ab3h1V3MOk0mn5NhZ3adct5iNv8l6UuPAVaOTMenh0XdpE
voneSN9c3mR1Rbd8G6eEZehHUl7jVhrXbSI0Wks5f4fA37eNSUGU8343sAMefToY
6gjKs3eDnpWljcoxBme/VSBUhIEHRHACdHLeH1vPELVuUFYmZmvq6DMOZ3g+UAWP
zRawKURyzkTBTbuP5u/itW8eg/1+gb07yqlmXtM9HJtfcOghAXK2l/SqZo6L4g9Y
Zy4yZbp8UI913u6uSHvTiQ9b+bnmK2a5IHxaycd0VIOms4f039Ri+ZScx79WckS4
gazDkMOGZJgt93Z8Rs77u1U6/AwJVBylPxmkWKGAIkoH6UcBsi9zk1EyldlxFLlN
Z2TDmmDO46CpfASpZyfQ4MQGi6aDmC2aBEcpuI4G99zWNIDCn9xEwNbumJWd+dgU
upJwc2EXxDBbu+Ldc/Oj9whDPIQXtPcoPPN/wnuIEcROYJQ3IivEyzcPIWSXVDap
tRMopM0Zvow4hnN24BD1fgvc6V8F25AjsTQxQEk6v7MoaZksLd51fbxRtqtRWu20
PLjc20eFV3VBTsiIAznxzRIcWYFMLHsXhmuMK+lJNr8jWXtRdNQPVPVrm17CSH7s
XVhRfzjMD6iaKIcZlJ5GQAH3P+z9mDllQgN1rzSbDM9ER7msQgtSb6T9yAcnbd8+
WMKZD/h5iJFesh+Jn0dFxgu6h7s5ilf0aYDpsRDlRUBodzn5CzkdBovNY+gmv5Cp
xc9yd6+28PIhMl7WOZIXwiEmQhO2ZhfxmKD9WEWVoDhj7Of8spZNiCf08+QLUjaq
xbdoce5Y0upvpH7pDeElDpiRQrROKE4lEFb6lLOtqSEVovWwJTjoYrEf0RZlFQGH
oW1r3zb76C6AzyD+fRwsl+BQCuzyvu+/GX02OTuQ9zZX8WxPKmWV+R8yPgAW7lJ6
E8Tzs7kqj2dd5PjJ5XBOGVvSr1q3Tic80E/4qZ4V/tWpzz4RtM1HEexhLi8GAw/5
uh6t8CAE5DbXXJfznfRWMrysOw67lj/fJlerM+16Iva5XvnksWiTsp9KUoQklX6H
jevu1Ows2yTu1ZOKqcC9VSLQZzBKvayw/iWsrP3iXYRucGicyrak4wf2cEG67i3D
LA/V0dpCWY5S9wS98SXyevnakYNJDQYj3heYE/Osc6Giocln+PMnfd7dxCxtDq5V
jrdM2lBWP4CjZjsNl9jjnc3rch2EJdjwz+00ch8P0jAhkqZaJ8Nc5cQ3K2cVGPT6
biNvSx+K3LT+en1mNZIWChIUwQw6nGXHzl+RpjuNMe/9pAEBpB9Xk9uJZ97opqvZ
0JPKeabwNcxxqY1VceO5Zs7Hr+2oxxBgB+meWOcUJaWv4/0Now7BbobZMFifFJ7g
pC5j4qaeWGbSg0usM3V1a0REUU8WGYkhtsqNI6f14lEx/tyQF68tVj8VahH6/ZAi
cB/7cPHqeYEMdDreE/BYFDrycJXOAXQyDotjxf5B6YSXLW0+q5hklRENlWoExNui
m0eUHZNCx80lnBUxm7XXOlqvhwhP/URJuO25PgXZUxRfhVRpUtBqGaKIRBG5vKiA
fFzQLmY9bm1XNH3uvoEULuJFz4dlGwLfj/az7QQ36Hro8LQelOBAwR7GVz49+xei
Wbo+0HSZJV150ZtdRhElWTRSesgx/ZvZhSEQohNoh5OPRGjHi79lSVJS+kgnkR0y
Y5/azjp6U7o/yBL/ka3AFTnv8OKY37VqOWqfOFVmE7z7WJGxiBY/praR12owRFao
FC0eJl3dLY63HJOfXG4sTi+fGuUqxsaesMX5yrg0xOFdkD3bjn40V95p20cD09nk
XTE2kyHmt2EahoSNMKdvAk2HIeNhUzFMm/srBIc7TTMWc3fNFUM4sq68S0oJDlQh
pQg54wOvJvtjCvNzVYuEQTTpCkxViFjrvoGzPpT2vOuYZflLgHPEliShIBACDR4q
UhqL32DN/MnVuVKgvp1/2Hkx4Z6EI21/NMe5vNtTZliW0FUdqkEXl0KJpniZBVw2
J9RlxxEDGPgUqdjWtyzPudIRU9ZYYIUgUfEpnsSVWSRPM/VRbIsPN65Ld2l9GIjh
tC+L9rWtzdzIJMaL4gwRtRkItkyt0glxAYgGpHh60BxWXxlQpTv0XyUZOmtc7wSl
5a59UenXBa8S3BqFBm8eLnksInUqtxJ4xYyTC9pZLdOuO0AThM6yTLamZYW6vyEt
BAPfd1BRf8RMTbZZT3Fg25Wpg6tocWl9bHHj5xj8p2DJ4lt/Sr2VcXgKXhsmZmPE
/Ckr9//Z3EHtpC2sF26w/FCt6yqPByRgG3tDESvyf45Tq04BG0hpXjOxomy0OGtm
ngTn8wImQGW7cTupgeyyCja8neRrEVlYveDreq719UkQ/fOmYGQHzK/jjyJQo9yl
3bY7sHKDQT1kbYo9e+F0kr8eIBpS0oMkbLyXdYgsoTU6KpTClTOipqG89xN+2ZQL
4cKxjHZt7lwpLvfoPixgfS6kgnL1QOy8PLM0Y3zWJdN4ZUNOpD2ds0wjaMZKwRz0
zq96lgseh2mKDSaNFnA8oXy+XhyHd9ZJvuWqSv2Gpg8IXfcnT1PF7q+eTu1qZ0xX
YylRhRYUcd1l7qtlydcjy9wsCpmaRvsXhs11s6qEw5ECnUUbrZEspwx3PW+h0SKi
94q31LIoXi5oEp7Cy2mNU7k8BVPJhXDUx/qYDa1zwsBy+C0n/zShEinNqSzuiruz
3WHtWFhuZtmP5yNSU/a5CmnyWGgw2YFGKnm4mIa/aRTJruoNDQ/dPpoqz0ZQMukR
Y6/MBMT4Y1wdOS18k+gJFGQN/4J1V7sZlu2kYZBlXB3Vm2wqSiis4QbGM+t4cbYV
rHlESoZF0Y4/X3yxpTruIJNjFy+tOcXf6oG7cmQW+WytKM+DCp5yyElnUKJES4vK
9e4TQh3LDoLWQYu9z3RHvtviMzGZ+L6XeG2ba/mZdy8LrL/WzepCMobO+cFCn5CD
dC/wZauP1oHZa7LGOA4YmLUH10JjIw1j8WTby+R0bgmDtaeO/FR1LPu2TJTM5irD
w9XCcphrORN97QYY0Qr7h2pS0fRChinZiifJsEe3iaYFnj1RR4fy8EezUyluwvw2
T/6a9i4KwB8O9Pz98E9u1eHLHMXJ3zW/3Mezn9WrFYiga46AkjhGsus4pSV7/zj+
I+ku9qk1nlu1YSzKN8lF6x3rQRcY0Vi8+AMR5sXHcbRa8Dt9nnB3A+hDsObtsZzF
kzG7wCMX0KfisjejLd4DMthuRpaEU1M9PGnz6anoLSGd9jjXTorsaMOEPO+TbBSK
OFLBcrELqM12bIri7UTHAr3U3ytIotgL4Qm8kjpOx/6YNtAzK1h3hD9zOC5IvWno
abPjqU7RD+yPAgthnHPJV6JeXiI1arkF7XrnTG+RmCWvfNlg6NPhD6B0gpi2sMeE
m4wgUDe6+yQoOmWs4HkKSaqt0yPlkYfq8cfCK4xW1sn34KJCl4iLCeBODF+1qAh4
GxW4Yo0VoUNEhDthrbA29EN9MiB1MnFVE0C6+YYcQA/gIo/BpU7UQvLNcAChYb6C
7d3F4eS2htAeXSFbthP6UlDSjbj84VjBzAR+MO8SS7CCCdplo2wGXWYvcm97/wuO
znarW647LsuNA0Yhp5CNC0uLT1LgvM/WPokZuRMt+c/MZ8HqBsTaXj4IIjpgbcSV
JkCU1HOdlHOygsPGJGhlhR+it+7pztsHatf1VktJwOl0ikgar1RQNJOmsfBQyh7K
UWI5vXmJjeRWsDExizdlt4z+Z79UZh097FCne8xXpgBEMmodsSiCvV8Ol29MNfNh
93Pth+Xap9XSmGWBFoBl4hEhq+SV6dHLAe5hzI6iSkBM2r9jiyjFBG/Sht7WuZ/t
NtacflRzGNHYbrYPwqdEBA44N99CLvwCV1ZCGRqwMixPiuU6nLdxG2gqgXSNFirn
QuDhtb9OF1zma9dh2vvTR+XLr43lYN1xIEGvt5PIldIt9Z3qP9pZWxknX06hv10s
VoG4Pz7OAZg30R0UBL9rBLN3MRH3+Rz3Tpwn8tfxDx90Da9/nvgrFSzYHQwOdFvq
njcLklCW1B3SODgPaCthJIHPHTKcA3dmNVa7CsnZlUNB6++R7ui58TSy3vzYpDMj
m5Zt0EsZtViEU8E+KYHU2pchfr1FcJqJzsBFyxf0RpFcgoUIqAgwY6/OFtuvKPMc
MxRoBsTJNzmSRfsO2n6U/0+aRkhdGKWUVgEFOgmqs16q04L50dMJv8Zs+c1bhOPy
G8zF0HHR4rqkkh32egTZZjSA1G+65JkUjlfIsdDnry/XVI+Gp6YUezOlj/ttAtGR
HJGBl7SEibxDFEZ79IK9x4V112wo5r1o9ZCePJWBzlAMCohwq/YZpYT6ajKO3lQu
bOoHl8eq65C6zxPZ5pbfErHOTv37J/9wlrphD1L48NFo2hJWG7A9WSomsxSaMdrR
3BNPUo9Ac1jt/vxoE3XXB6M+1jvUQQyEC/+ZN4JXoAnJ6udBB0uGKt/U6j3Qkbn4
9aW2OuDFG3tUMA+5gS2yrVrPqyWBuRIMXH2vyNMgfIN5At+uQKEy+zrCCrAn2A5w
FyoOfQiSxuLhe+pe+nD9hh7CDVRjaOAocUmdHj7zX5gmyi0gfErC5HkIIerH6oKu
IE/JthmH4QU0Bx0cAag2yd28EfsOz9AfhPOy769UF3wpq4SogGkHK7xEiwrucsMY
IR2uRjqfq9sK9JaRTQC7MV3WTv2zMnh1nztDTqj+N2gmRasgcb1NZkFmUsbflATk
7UTcRAAP9QbbiEJkj82iPGW4Bq/943tLbP/sY0E6ykTW5D6fD5Aqe3t/GxrHX572
SEor8HKIUsvJPUog9fwY9KmPYyM2L7bUF6aTZfWhB+S0UPmChA7NvPHQnoj7pWd5
+q94BC3j78UNqUeXqrXiIVpvNiWtx4Vv1IVoJ/fIpZLoND3P0a160xSCEslboXzp
vySFYZbsEDOYEI9okMFPSSqBtfN3Ahr74z2FLu7eWe3b5IP+W1NBNdKLPXPqcAlz
WYRWmq+oGSyb05CeE3Fe1HyP67315tY/c63xgYCZIf/JA9VcMr2Lz7r6U+xFIWQC
Z30CFg0tUX68WwJgiP0gQ7PMETkqcZKySMa8qMOkUWTQDBZj6Iu25S5jq1EV3HAF
jhjtBDoTw20J2qiu98VOKkUTqa2d9/WAblvDQMR2P4RIzxGDc8i/qeR13Ko5l+18
RXo2VPXcOqtSqAJRGRe9Y4jaT39mbKfb0ndmV75RbMAfmShe0yX7qcTb4X34l8zg
AkKlm888DcVPiynxgbG6WLIrakA3Yag+MTMCtjvroQBxdd6IHdO7yv0dmzNrtLI6
8Q/wSe9N7Jp+mQGde5/8oc9+GpRF8KOIj56ev0R6e0M2IcpJsFPk+VsqPUZK4fE3
Duy9ZT2B7powDfp03b6esgTXIHxf1+EP3SRITDQpDUn9pqkMZACghe6M1/Dh7/+i
ifUEpEOHChEPyW3ZHYLansbVMlwcIvMidMZrdg4vVwNECUOlOjCnO69v7sKhN7HJ
7dgIip6n4RXCgvDLPjDz4nmXV1MwDZdJvG1iBvl5ZzbDEjUDA1B6L8Czub5czuRN
xagUpZ81/ykG7Z/lgp9qZxuIPpBWJNSiCj4xbU/W0Wy4HnVw3WP6P/ytqIhFb9ho
iGgbTvDy/2BtB16juJMC3mXU0KkntzyXnhzH1cuimBXd0TRUck0UbnrrnTyq1Gnn
JkAxw0M+Vy7sITUKizKZSWbKxdC0psxwPlfRsNZSPJdDnuVSVcEL/4HYyW0KvMlk
A+benK3eINtPUqM4wX5Zo5SUg3k+go1bvRx3kT3YgEoR8Fwwa89+5Vt1sTiqlOWM
RYU0m0xc7glb7IhG7dugx+iCTPUts68WXA7gXXRnZoAWvFBHlZ33DgBp7L1DufJe
K2WeonqUPfjX0s2tCuEO/9oW+7n4u2ieC5ZT2t11GM3ErQtginWD9QGT8qBUrw1n
Nepin3rf+zqavVWxbaf56eTTVOYHz/VDn+lMO/2NeVzVUfE+CiwAj2ssmyS1c8jz
1puGSY2bT66UovFkaED9lsyV7H5Bs2sb3LHVPpED0zxYxI2BwE5QUMGGQo0W2th3
xvHrS8W+0BuoRFgdHivW6DFqjq/kJSFeCY7keXQtLkWTpOsVSsm5lQXWHkSN2Ihs
a1kjuaFyQK+11Zcl0LM0z8knGzEiZVqSl47f5r8wWGRDAuMOUn2LtRG5Rcy/txET
Scn1EMkmTjOF94mAdjypRMFEPRYB6iuo00ZfA47MhtuPgAe1CarxWUlwznx4WnHD
xj1U0umtb812HFOXGl7pZ0WufaScIYig4ud7es5Jf2ho4KYM+1KZ7GzwLO2z791U
rEwGZnSfhBpgcNCrZynKLdbfqQS5F2xZr3nFmffe58w+VAS4FrEJKjdFM9OVGs0u
saDMyHuc1aW1MrYVMzdADoB0CTjBYrzZebsTWT8kbGMdZ4N+QGXn+9Rj8ok3gFYf
mUJNE/rS3SoOYYmlMDheSvGmdJbgA5erFEUIGHE/HSjmr9VLfI94epbCEYuLbD2T
Wq5t0wj9fYOfrAc1dyNB/fPwv3GtGXE+AI4lT1yRZYOTY4Mf1MZ+DbOUjs5rc79B
VDDMaB8uIlkXQxXCwuNT1wKBh0KvChDRNa53jwjfR5TYhj7SMPvPWUQmNJd+2nCu
idNLK/AGI1c0pu1CGWJsBFAIwEWj3/6XwtBCC52Fs8qvHH0maTxE4A3AjAOnnUMB
HYjS1Vhqt6axagrhvpEjwbmHDckhd1HRjlJifFylhAXN8uk9LBzI4KiCRShA+CPk
XdwvN+t8PaN170L/a9YS3uw9/W7wKZkl56CRj7DFOBht77kEJjdaejPXf4XHQ6rJ
RdLO1n0bNCHSbBSeDx6JZAPNJIGAKENbsyOaojfy/FqsD/4OD+WpcSekjiBd1ujI
l7DDIChQXdcbr2LOKz9/4JnSiTwk2V9ovN/8oEVo/l75EMK3460a+GUsrvACrqY1
RimbOOct8NE185YFNPpxm1i1nR4UN0lHGkZ5W7N7mvNKWdQ2f8U0jZGwwUEIZD3N
Ox4mYpldDi661MnaRUwLdUee4koSlVhjuTcviADdRb/PfpcqYZotUwaaqz6tZMO2
c8KuxzPDiAjy13Ll71fZANHRmEEtAkYCJW3k+OCi1e1F9EdJAgpGELJZnolv3iT8
jeN2i47a5lwM1/ssxAw7/kxay4Labd02WE/W5F9/j89zLMpShAPm1UFOscc7MPuc
GeELTs9Nvgn865N33tjWrjE9acY5oKyAvrT83DWMv0eeehT0ts8MiKPR+8scgubH
4vokXAYlTCcUAUlBBtMSHf/djVjBEJej5L4M0VaWaPGCW7j9sgEYxpFPRrViYbWb
VoRa81BEQX/8S/hra5WL/vzBvQEmiEph9KFE8Bb0nAhmAbcve9N59Hze2/J/tZQe
Sn2u1+X6hikFYjlWFRmRaFq4fT/4Kd9iWiSUeKCURIFPL/KIcd/4OSo22BzwrBvu
sLB+nTTQjPs5P4NWEoK8a+kOeHYZlkxQ9bnYND1JHjVuhcNs6nazAXEwARpUfDBr
wtiH8Q3C3a15QCDxpbp6NeT424sqZg8jQUV7YxgieSWJ6iWptEDM6l4A6b6wnzh4
G1awYEf9BVG8K+vDfxMvByCApGMEmMO9icKNrruwCYBtqu2jGgqKemvu4k+DAwlA
v8AuuGiOZ0mZD+PGT+2xBxutmVjRM/qRLOsGwBt5ndf2FvH2d0NdmRhWCWRtTAMG
v+cT7ZMUAkdJyGfrALV0oSiYJDvDY8xFtbu9/4DfkpAICFZpKEhHgL7C5fnRYXi/
5ZTk1OlSEJui1EPOAKxhUvCrTPYbJBeXj4zVZg3qWMm9r9ubSuJzzDR5WoE+cryw
9CcRAn8h20+5SjlqAl03gGUASN6DBlxpAvRiHwt8qCpdA9+gR3uK5FmtPAtNu53D
ie/bGLjVjHSQCMt7himpFBH7ymQ2DOlOZEIuH22KLbzlvlo8jrQxgJSQ/7y91r22
C3EFZ6c1/WZKIQrSOn5wlWaf0gEoSkdNUhU+OriZf6JMs7jsSDkRBshF3d9K+OZt
BCWWXGYZY6zVatV/AiKccptDpaXsWi+RALrER9tIIFW/k/XTjP02fZbADTDNUA2y
aBH14MJ+vYL2vusp8AG5L+Dvkcj9VhQwD12kPgHHv84LlQWw1wq7+4x77eZImoUN
TalIhlAMlECowkhZ984T4DyLeAwfKAH7uWDTn8NNMTqPPwijEDki9rOCNGiHYKOW
+hVKSddmnxwy2K+Riob/woBqDqDWs5DyTA2Rx3igUpPsK4pnf/XhnwFw/ykPXX0d
3am+YTgR2TeHn60Qvgfu6xLObG6sIvi2e73TjzrCpY2EpuczlTXnJVr1RUtvylrD
pc+vkFe6GQOI5TqSUZ/OgV62K3t2MuJvoJ2cLIgh15xYnBmejJ+DBWJ/KtkjghMX
1vTTlvLcmxTaic11dZCf762jIpK1J4TJ9zJ1x7Eo9qGeBYCFw8izp3IRbvAyuGyO
Y7s+4F1Nqbbui6L98qPH8SLuON+RPu8jBBw1NScn//Ot/UsvDqcKmDLNMU3oJlsy
hmYDNv4N1CF4OjihCRaeCRNyk42KyrEL11v2Bio0u0EkK9nnjq2O+5yq+9GWC4g2
2MzkBzJ/gpPbEaKwCP57RjhmJfXhVUQIZcZehWp6Y7HD9qoTfjmhLiEvEwkPDW9w
vrHvnS+rip4aY3CUel+ln4elU7qutnYWEu6mBPAawxuQJeD+RkqgmV24rTENgijP
bfQWRXmlymN8brEvfsL2u57H70Bw3xhHWfuZW21OFCbibInFBs9H7CZcnughr/PA
UFaZRRtGxvLGtQ3odAeZSWn35pTr8IpywUuN1keA2EQ/B1qyVfO0Hk+XzRoJcihL
7U9g14JtZjA8pmDPMJDR4I2t9bJcmVhC9uyn6EcqNuj/JZ9A/k+Xab652sYNqAXq
TlRi+Zk9FgCq2RSZLZoA9PiqrXzN3Yny9kFTLE4i1U8FX/rKKe6a+qyKlxB18R9y
FXZUKe+9JKL6dg1blI0bouSQWMClyoqg/eIFUzoMK4tZUIFSDEzOICEx91bsHlSW
tDvgNmyrXYUfeA5B0wQdp5jorKZmyhwPJruRjsebrhom/3eLQ6NSID8eZZZODvex
ieDQWzJ3VPPFt1Vt6ui7PP0oHFMthJUswuxEKffrGLPKLAhnbr2EACMpt03Eh9BN
x0SFqYsgou1A+6lqxRiV5NkaXjkZ7EkPjNVMSY4bSgbkWZxXEIvPtXWdptqu+uxc
ERgwCIzdquMCjrDuz4qUVb4Cy+0CX7Jn89Vf+CBi2kKAh1VYnNm6T44EMV7pzOoP
hJR9F+8UO6G3TLV4FxfjiPAQmGMGFZQzcr9EPsH2M8kBE+IHUmItjKXqbRkIhyie
zvDKan53FYXMBmV/LCXGUe4UaGVSbUhg4FC3THJR5zJYmS1q9hgULqUcgacJXkpn
U6imuoFmdIczVS/DjJpjnlq1PgPLnTjXZZIFMNzcNHVdgq8gBmjVAmNxyW2eAcRW
IOiTeQTEJuiLElykaNepmelEGOgG5zTBTZzC9aKn/4tfraEyMuYvaLvd7QY1mALw
7R56x0yLu4KFV7jPrasnwfvhQGGIp2IA0PvoWYW03ufb4EuHHGDNgwAJwRhiQglz
IxUBsrDz5Pf6MuG6cm/dkbfkyQee6nfIKkP5ioSi0G42qW4fk2MEbBWdU3FxXZMF
PZBKdCMLALednvxqBNVGdIzkuPWxRgw7wrVC1BD/y/qnFOdNMCc9P8m4bih+EyRl
52/mTFWvf8tXNeuA8TKD7u+WjeOl28Njcm8NRlcpF4/z9QEGjrTVqB6J55tP7wUD
W0+gh07W+jkIC1W0zhtvaKUCIa8arsQcS/Da8GD4BGFjcOrzGCxGNaEZUHf8SciI
e3faONvrCUGUcBRaLnpVetS7OMlW3O+MHc8mk7nVI5UUHaDBHby+Y6g+TdLNPq5v
kN1a3VArWyvlfMtKNkDxBMWeRsjfiYC7ukPG+skK+Ae+mqFU2mK9wchsS7c/0a0f
z30Fu2zKPb6r2GNZUJShA6AG7XMlmGBvxHQSP/VgjnksRqdHal7UF5BZ40eC8xKV
zbmpJFKcE58ZKglICqz0rRiUVHvCYymCLe5e5Px8qDO1r1vtii4FEMLNbdhF+lxc
6oRZK5c3Xv8fnpN7QQz0z/A64ZIhFgefe3biCmUWILNyLY3ndEOPMhkQva20HXKG
ay/cSXVTZFKbnKMovLHIAXOZ/QL7MrW0+TJre1O2/ESHCR6tD1+y9FhDPKyOzPfZ
xM1h97BPQI74yx81hvyYPS52vp94V8WR7RcO2/vf6V6l2efKmFs81HTHyjTsWtkR
zIc4Z+Po98bBqcFwLDYgDs6WEhfGddv2WlenrFL3KEScIywZTu1OH9MDWDTp5Bme
W6XcUu/nlb9BdnA3JorWAUKsxqPNceb648jxaBVBVgC8GCgOrQfMeRpFxAEidwOu
IHz8dbfI90x3t/MlfWf01K5+KFJD74tTG4bSoX/2jj0u2iiS4VkfWXeqSVltbD1F
I9nnyxNEu+c8XXb1dRiwijT3nLJIzPu6RQMaQXJrZGCaoxVkOaKGvyERw6TgBMwm
5SNPw3u0KekhhcIlf5Z816tQZyFD4l/5a4qdfEvMT77V5lzHz9Exd8aoHluCvQGj
TAkLEHwfI7G5W1EibpW8y23zOflo7wrmr3PLzMrKostq0wE0pjfPaov89AzSw+5Y
De1aRR3v6mbwpd73UVVCkp+6M+G7c09oVWI7FBgI8V+bU/d3yC/ycDmIqH98PKl3
BcnqFWAcWluihijh1rQsTU8sBnPtNd9MuWWjRt7Gby43sLXEfIIxkwYxw1W89Mq4
eMLaxTCKYPzoiNGXzTBtLfZi3lrshltjr/oIN0E+cwT0aW9C+GKxrNtH9IFP0/Rj
TB9DAOBg9H3If29882HhK64F4wxz6Qys9a5muJ8430QXGigzyBhtH5lGlWZi4t82
T0GW1S2Wo5gUywGJD0EUYvpTl7mS0U9WTBNMcRl4zqZTxKULNfT+1KO79R3m8oUb
lB47dOmuPuzG1ZtV21h5yaQ5yOR3wtGtxI3zm8lq81jNreHOnLig3fQhkhYFv12Z
TK26QcrafaV8delo2LqFVJnFhhPrPHXQ8i1TZuQ4FEqo3T54NJYnhvLWmOSuIl8C
sgpew9pwWdPVdDd+s/cy1sGNIDi67VJf+tHOiXoQBGqn7BRIliNeMc05YIjH/YrV
hfInKCy65osPmGl3wFo3VHxrqOTJYg0rNjJN1iJfW0e599vbgNfdej5rafcEdh5Z
vNPOM1kaojqlkTMUs0aD6cSCuc3YjVC9oia5XebReEWh6A/aNKN24L8h/CeY6v3M
BMslCC27Wlkraqhv/UncfwEhu6uTP9H2KhMfFAxKFjEfZ5XdWOZSIN7/H6STWxTv
WGoJkzSsNnb8yzK6gaeujgkRxXVxgeqsd54DwMtuKgQNGP93dAIW8vMv79Wx1IAc
7+9sDW0X0xwF9dffBFyQmnvN+DgpxNzbBNmvnVUE2v0HduNDY3YU0nTFLAnl9gLV
zishB6If6AF/B+Fk2E1RJgft5x92A/RCcw9RDTi2eodE8ziGpkxQBy7qSfibTwEh
74XW6ST8wnIN0P58sXi5KHEXd0/LhlWCGUHli5MEYkQqBBy0z6I5RAI5A1tji5hn
EMstu9nz3HiawYq3/huMnLBrv54CYv6Fy4hxYpNqh+sK222Swumuc3bu0BDSV6p9
Ahu9MGFeFyeKmLFWwxk7qUt26tShJ1mxm1th7a3CC21NyBMfbS3LxH0PFtNqXRLL
/Za2f4o7uZZ2mCshtsShMmqG5CVDasQccYScbkp7gtR7ZfnUv7urHkQ6OWGdcVMt
5jOICJasZ47AHAZfTZuxo7pDxWQMvX7gBQL6OckhyYbtN/sM27wtndG5ryl//Kf1
ZA4ya8xRFyAraXGxcwtHRnC1nav5FCRA+LPH8f0DiiFyy1UOu+hkf03nSSXUBqST
ECIPa5EXl8lF/sCmYV86TipglrcATihnlmcue+qlQS56HSfC9cciI0wFX/lq+M7H
g9E7oq6Hn1RdZZIbXKXSkNYFh06qjO7a8Yr60PbFUG5cP2pQeTWzk+F9PM0TEi4P
3JczV1sSBnGsxGjkk2yi20uTpOaizdbm0RtChrrgYVjzB1WfMBj68VhmU0ovDqMR
vnFFrvoxLQ0OE6+wuo+DVMURoATQSeMUlEkUFMlICekbCQ1uGThz8n6Si9uJuiIz
+nbizOU9BDalDNlbLp/otP5YP2Phv9ZTKLygctqrPpiwv+0oPeNpIXnNESVeM4GZ
k5u7jFD2Vya+0clWdqtwBYbK/3O7SfNejScbwAT2KkH7l2UIyy4TJhJRwJJtUTBI
KjcXDBYWrnlY5pNsDm7p3uvUPWbqscQkuHKlw/dTqX+EuSpYNhTRsZLpkd+j2x0p
9n4iFqKPBuQaAp4pXm2MLhA7HI4km4mgafIgV8TkZX8dUkRD58+zRlfP/qXJ8ott
fS23ntfiSgGLCBPsh67YeOIjFpBF67U0/Nv+qfNG1BRuJGtvEfmXdIMRBDs5RPR8
tWKY74CtnsLPZ19DfBiidkisPNGeEmAbG2gWG78PXvakxExk3qAPkSHtZ8YMDLMm
aPdGyxU15/SexcfuGa7baK+z8Dq1BtzayJcCtJ+DjjNK8oc0xNIRVt0/ZJlxsDFf
keBSVQYa6lhnv5HJfOHaoSNL3ygDpfpaQwjyG2vgUhmzNoXwWmSzCF3IgTMx9TRo
g2yfShHH1dTE0UESrkhgyfZGlJ0/mwhOc1oDhixIbqdBbNerUVO5ig1UC0x18eUm
jhm+qzfILjyU+WcKJuaiOcZzaTyt5qOkN8Jfivjr3k4h3KJGJeLZ+198GNk3os2C
PRcIzGevJzkU7Xtb+M9nZKQiYdEM2LDLghWizySV2joqn8RB3LrH1NpnoaJ0GtRS
NDyHx9RXmnmQXON2DBfL67gVK/nC3F6Awwe/9eVq7+nolj5K4LVWI2P03OhBE6WP
OAc3WLeJEb149f2ijxBzNadR2+eXtHOsu0BrkJN7THqFCkBU/CsaXD/sAOgMf+18
IZN78/maBtTxXr7B9A/IvG2/7DqPsjqXatkM5AUNSS0872i9YL5MXCRnIk9pUYoc
YFQo4sMN0mzNAFkxO9F2fOWIMSXtjZnEEaiZf64WtKAG9HIYNSmDiEZYBv4Zks63
Htff8KuW94TDeTqv2Wm8z4KGk28Pe44wUnEIa7EzTekttJaq2MjWMBCSrYChIQ9t
bn2e62bHtZJe3nEYRFPOHLm+fbGFN+W4kE1RPRymMBw9WZ2TZYv1Dv/5IP6ZOMAL
RG1MOIUfSY54xuLMVFEIU398xmiWO1d5IgzHtWh3AMoKeXo0Ths3OQMc5mot0EoT
zPPD/ZHghrcAU7rIbaWM3qWAklR8RvUWzzRaMzUdKSfI3BTvC7Y0tsglkUtJxDmo
ehjIT4oRjVbutI9yIMMu1lPE+rzlBtTbnSDANyNhrrzAOzm5vAwoxogitcYA5DVP
DliHZMyY6t8qq/DCmwgRPFbfiiqJ9qfjzg9K3bMwpoFJLInEOIso8NE+qnIJy8ip
sIr55Y6oOT7b/T7ALc+MC7a7UON1dYZGeTg6f9nIrPgHL2MMrK4K6or8dBPgtLpN
n0eB6vhfnqYNWmPwjimJZwIdDQznGNAjAN58PLfUwwBspz5+ey4r8sU+HZCFW2lM
zB7mX8o9oiUX4cK7Ou7Y929NsgFbDu9OHH42W85/vG5JwYbgc8Fd7CbIHA/CRr4J
FtUm91X3T42XB/xhKoQMwOq0lJbPjICdaKQwtKU/Yf5MuprIfqBL3VriUCOeOAaz
AuTWmOSdb7ZVqkDrO7yB1nZP3BBONBMQc5R5x//bSwq241nYoU5ZwGMm9myVwjHP
mRRLHqB3rtRaexoZVb4OwGo5JcbHl99cBhJ0xXx154jnFR7FoPDzSqqR7ydr0etm
IQpAt7HQpU+HtbZiikXWyL77UMAJWYsD4Lqk+070C9gGGqzXz4fI1GpjOmE5wws4
xwxLt07hW9grDL5unjkfDsuzXJMJe/avf/zksUSK8Kfmw85MoZlW41RjNP9aHhlv
lBhKeioYoYjMTgql3lEn8xR+LgCNH5uSwFXQMxF5rQ0/Zh4PrFbTwtEq0CdIW91s
7l5DgffgPgvQagssgG4LrTuOw6TvI68+qGUOx0NB7Hb60RZrwa30Lf7IbqumGE2J
6pWwytSj7hDOtSlnzKyKeJ1vjLbPG0FJfJBKn9ym19FwAEIOUNL6/v4qEoojfjF4
hxn8D/QngPPCcT2W6yKXNDvyDIwBJDmRH8aoBE0nUuERgb30/zBkn5JSLuIRLuPI
tBSVkzKDpo4aFlA16nfAVmYN8biuNdJbVKb0RrLpTgJN6pc/EAUmoVR+hrKn2Aao
9QfYF7rk/9UC7NDbvcg2L7dV6/YoDj01JWunUW72bul5HybRGMtc+7NhHLEKN7dc
oIV8Iwl7wC66KkE+npW1hA1BDcM6n53gSjXveG+rVjiSaYVJeUe6p491GLKR0Xu5
glOCReR8TcTEyqcZIi/k5N1ucMEL7or7rJGjEz6Ph5ncMTx3/1Ll3PbC9VQ2Nb/9
/YrwYsMTtsCcH4kthLoCQxuCgR3OYrtqgXSxsBlcMAjDwwSCBQBlqChUJeL/ht4S
r2eGcQjgvwJPZtBxuIWAJEfb6z2nYl28A7xfDBoGu+WgPUNX6NMlmqOt8ySJJqAZ
zSRoGZAxtZYlwaqDTRiIFxBX30tE11BfajSOEEL462pjCDSWj7Rbv1NsBOg6QuvD
jvAPlmf8e3SvjXWg6kig/6C5E7TxvqbksxJxYw0wA36WKwpoVd3cc1OVyOUjJvER
XOr9D++FkxxDtE/HiZwsIjt1wKPJNvCi9ACO6p0vtY7gW5uCTqO1Ng1Gbb+Icu+Q
YaNzykjpQCvYszR266GKfv9p1ezZtXS8WzSd0MtUhCHBMvI3/QLApw2aebodjOrh
sYPuZnxLj1xkQAbI7CeYsFqaijFXq1B2TD+32MWOLVeUXOAP742gfSQdhd/oHy53
bYLWqF8UY4inaLeh75x2tDZb8T8uEQENP2kpVHElEOq910BkJRvfIj4k9Fyq1Lt8
W4bh5q5bTRL08lp29nzrDDxuPJh0Vu4EB6lkBgMQPMhG62O0IIj2DS1fxCUKZBou
gQBFBchqlpG5IkdRJn78hLM1kF8NHYUaXmlg7g/Z5ALKhuhnBxjX89Hj4tfCJK16
3QJwfc+f1CM41GqZNMBrUtQm6VBdsndnTlORuULBpXUEmZ2xduIRuPx/J3gelpnP
ekbYX/5LLIPL34b/aXvsZFw0NSA24jXJnh7/uDDFJ5pkGIhwDSwedaREihDUh4Lo
wAym/eK0+dYwJGNy7zc9aQRGNuVqCdCEBxPM6Uib9VX4hl8dMpqctPSVF6b6k6Q6
79jBiAj90HVH3ci73BETkPUoZXxlGLHL2mpfC7yWPy2oBiF66n/nrZmn699wZXNo
33aZQhSCCdDNZ3WjNQkzZPRiTg9lvB6OFrDbNYzcXLBnB7DW3SC6WUVvenh97ilw
1qtwWdbNnIsl9WsU/ehhlTXJ404IipbakRa25Q/UcnxEsrk7QwjLy3rxbex4TMM4
IXSZxquyTYdA8smqhR/4pu2dufM2fgmSY84xrWZAGp1+EqDpOcN8IZfOFjuhxJdi
XtM354puuFohZW7xzi0hzmUjXb731OtUBq4AIRePMvLhdRQ8hvxnq5hRMOpCYPlL
WQauVai5MKPBBE5WNdZt0q2fkJmRjrdvZmUpdd0mKtNY4nj/ffVqvpwnFrKSqWFF
e206kDwmwYDjhMnyEFxLuhlSNMwP5cKI3Xl9XnyJ6y5nZqrinxA7xPa0CUHNIkSf
1UUduCCBA9GTex+viWPPLjLZlG35zJvpnU5mMdmg/HlO/rXKwbeeRay7MxtM9IC9
P1wFkpHlKvrriY2s5rq0ZFCR26YDXFil+pu3DPVkhPLRV/mA2HV9lyvz1wo5EZp2
YOx925x9rEj6sOTsV625y2jqnAM4Sl1flIQ2B+8A0qavuy468bPAl0GYfYZJfI3l
SZn9tJCQlZbmnafkZ7ZOGGXsdPAzuqmURj3ymp9r/7o2Kf2mfgI83vFmpBo4Te2f
s71hBTsdRSeu5cCZJaKWdNIJRlMwMqCyOqWFPMBYmw726XU/pNrLYswN7VmdGKwh
pgG1KtyTlQAVeZBeL1HCKsewG7GP9QqRN0mDx46nQOWqn7V1Bx18pe2xH4D7RUJm
t60LGaXulJyIi3/zp60SzUohLdHspP+InrB8P0LCOn/zP7azxfrb4a6mhypasH0O
Gw2fiDddDeQhZHH9oaA3cFhk/DNF2d8FQ8NQyRq5gpRGzT0GrPSVzqw0tVb2KwDr
ZvqroxK3LCoyrzS6UqEM7ZPlfzcmmrdo+eiAQFkYY4btCaqzlH7gN3avA1djTn0V
duLDywP9Jv8IIw83MRLN79rk0Oayc1Gq0zNw7PfsYSp7u5jefeK7dOLtOqwp/whl
GFjTbel/o+mHG/uzsuUC4Iaxz82h8hH2JLEP4rz0rlYL7t2fG65oO8pJWgBaz/Aa
6fqtS2HhhFmr0AyiKEaedH+8PseqWltQoohplfmo+aPq+hG3HrfMf93CCkN1p3fH
PiJ5gAar/kM81gvAEFrAxdo9aOh5zB8Ahp1pDhXkCTupbQAQQt+pbm11spF9QF+b
Xqxj1biYaEYSHtRuhSvR1bNfyNCkqQkLGn4fkDdsjAeRmckbHAgrPyBeXLV/beup
Le1x3kbVpdAGrBKBbmXyYvMGA3o6vAKNI9OEq2O2qkvRWPp5wB5XfwhYMtoQKXXP
N/xsOgzf6dMvnmT6TbXugsGghSenPPZ3L/Fo5U+NZ9CnlPrMxtuU8fybVg29DuFR
OS/Tk6o+u5gFdJgsU5eO+UDu1k5vMQOZWD1r7DucieM6MzCiLDvKvS2ecVwxQVx2
ADFvAdVVBEZkqk3qMkb/QC0w/PNd3BdWz7zTIGwj2xKPQEOomO4ZryMg+IejGD8B
BkNkV5Xwta69svT1Q2iWA6zx2oMwlscpwixzhHJlDcrjd5XZUAohHK3sli69zBbz
hEsKlp/reFoZPWd1Nq+9fM5RAiIJx+tinr+vAkkupYpKUhuGL7kY1eSI3R5DKshz
0dU5yV7yvzHPyvjxq8Wr///oXTpRh9ouZrAn9Wfl3Y2Yp8M0INho5JtsoeY2+Lsv
k8ucT1bl0wY3Rr1KE4dI1LH1nD1DeJtm+WF78LipHiDmy0ZKdDsvUVXIpN4BWVof
e3ZwHsDXhVWC/sUbVhrshMCfjLG80rNyorV6QUXstA7h/A3WVluclaf2giHP1fqe
IVHBIQSa/eljKDS4RXWW5vVmM7YBMVjxpRcZ4+UbKSNeFcBXv2DX08th11hgIfUJ
Vxb9/fzeFPOxQM6MVIzDEm2I8AYuhgs3zAO7h8ag2J8hRLymoX4wXmXFtUT/uRy+
RC3xlpM1Z070hPwKIGda6IYkLN06EqOQfRccdpLwhos1aY+77LRJ+fwKEMJqDWFa
tB7VAofAe4rYOA613IxpJQqaGdnZ/odQRCR9FHTQGlZhu9viE9rgd5rz2V0+F0vK
UELk+JZ6UfA8aP3C/4flD7RbKDIdtOUSR1A6FGWfpx7HF8To11ZRDpbq0Lf4OEFe
0b7ly8EmZg68e5Xzwm92ttPoy5oUJNPJhZjY1qvPEh/5Iw5dpNwKc/dGMO3ysEeI
sNFsWWC1Yb0OX2s+YHZNpUYxKRtAAItLYTTUuHQagntanPO4V8t9TaG6xjRx3jvN
Ua4c68XKOy9fYIHhQtmlt32tTDHnoB9VMiCvLxTmS3V/mbJ0vDjz5GmXTjb3VLxU
kjQ4lNaOVCALkrUG2UBZq0ctVeJMqR6VEYydP34nPk7MEXEepxfJHZgBxaGSRpJn
i+AiMVauoi9tOpbQ7eKVdvc59s8ebwg1hFVNjBb6WwCDw/cHG9AuxjGCAYqRGYSd
Cjk5QC2boxC9OmxzY1MtzD+dtdm8K3EMyUmXYVdDXcD0EBxWG6Lvs9kD+FYKQwCD
E4y4TTob8BBDG9wpah2/jBISc4VH0rGVuvXreuRl3ipQPakSPZ40sKzdlslhTFgL
VNGvdw4hqgYuHhdHqCQwdBqVHKy75c2t++Rwv4fErk/dEbpph/iJn1ZITyd4cTIK
l5ZGimMigAlsbpDXomrX2CEcWN6qtUeVBTxdy2KlnenJkVs9NDakY9rFWq891Xgx
FwzGKMq9XwFF5z6LnTlfwIjMWJmbJeHGx+jK1xrDBGNjxMkF468mmzdZZi18/a/x
k0DfL3sv0dIE0xoEgiDN7im/ez8IZUk2+KME3xHuui05NGVOiwqtyw+NbcvRlTcx
VNOvvsZ+axOtJVC82acbr06Orb6bFH6/Ilt1WqJnj4uGSNrhvbDtTQijt/OS7xoz
x1oLOVVBHOJKiEsVLWYus3zE/8iHu/bhAEdcF+C5Y1IKYKjXY0hO/Ao0JTKuRQI8
qivQLlf3Tk/PcSBUaxOq79Z8h5oMm8DymcNjTUkz7+e5r5XmosQu4vm+JCKpZJW/
Uwy+ya7Xt7nDNOCa3IliIbix8k7mOMnrD6E5QbFzSGIy33NzuBPFiEKOnweOLrUj
DIx0CdUW2/CfbfmvuqdwWNi8dnCWS5dZjM1F2aldAaNQUFF5085pOSgdizPQug+M
e7ouXPe8F9cWsdphbCMm8/cIwnlw0OOEOnJdOnagZqDsugTYN70pdAwCEldf/92o
WQvzznLtz/GLHGEZCzuJaUCS5CcX/gBPtyP6YlDOXqtFmrMt/1YdYCobN1LxR8nY
tEN3Sgqe9B8UffXVoZSb8kqfRs7u+VMgrLW7PJ+C0aol5e7u5kNyCtfUm2nF6Fls
nfvXdDJbXsvkI+KIEJ5uNlkzOyzUL1hM/R2ape/ngw0Th4Uk5N8Qv9ywhovLh0QP
Kqesmqn/KRUBx6g9MVb0tQq0lxlkWGcMMHsFwBMZi3C2+X8SLnSwdpNLtkeW4XkH
rWU/TlZJswekMWoGlXw2rUaDEOmS2eCMHdxupo3ugRp7Lp6BbiCSkeyt7Zxzmjv7
wr3vKEFxqCp53E8JZUjLjf1w3ESdnLAo50athUc9lLp6hekGdj4BujEyOrnqQKm/
MmyWlaIj3UnIPvxV5j8hT6NE1prEMKs/6CTiz4vxD7SkX5sEOQzAI0ozSmDTJl/K
zNR5tuXZ8NdAEOBYf9Xq4EAy3dDNHpZQ2/p4WuOsLvKqfpUOQLzR/6zhhurbi84e
e6uhI1ANH2UenlfvYqf8aPSrx5hFjyaMotTljRCkT7PowIsuzHKJsG8YeYoj/tG9
tVli3F+IF8acs7sqIiWbbwlPf4YR9WIJTL1QxKjwXdTqOKKSXKz9Xc4XvFLJTbgy
avG93Rw8QAtb7hdW6MNCWPfI8UaCl4ylk+M3dv6u+JaR8lSHKuHByijf1RUsyqLH
mDWUgQThzNcKZ9ID5oeCEn5/Fb7kM7k/D577JlzW2PZhAUR4mqlSWOYSQIDMiNna
r+t7j9/U+2CHMsOB5oMWThotjTpLbsniC2SITPQn984yvYEQGybdjOaHeUXqi8YH
S0UYPdIUlbdnWimat/jZ7eeXDMBuIDsHuhcozV039ffcQm+7kf4Dc16HaRD02oGq
rB21CJjD+VnlSwOYIAh3XgBMeBf1ZnwUeBtPkGVvHpg8uSooekHNxEnTV2hRGfmt
QZsrYwUpALJM/xJdN5wSrsKHlxJiAuyUi6lhu7azw3RjPbgHqmkhxkwJIkjyhe47
fv6h6BpnhzUx6dvTqFH67WEwe3l+4/MrfzvmdIxMgjzrdsSH5T+8e2tBTQr2TM5n
xgCJXZNu7dJnmD59iweYyMo6YeSS54fnjAWydmMS/D6lyC5Iq/5Oa44NLFj8VzfQ
eff/IUgsqC2TB6fztD5qmSVxvh+3u8t3xAhyrSRVi+aZc7k1IfAQ7Sg0JytOP+7L
5n5dVbl60gpw1aomAewdO3/3WMsH7DJp505C6PIi6b8og/JwQu1D3WgcC2yRBsQW
SofSD077/hFJ9DulLYU/rhpSqmuiDTQRT3czh/HBGV5ltMzyDYC6d9dqiLny6YHL
sNDZgOJvq6oE6lXKeSMC0Q11josgYn9oSohdPP1evFnksMEhfZVTkK2aiW/ooKuh
nQU5+QR6ZXqZvdhtlu7BTub6NT3wqr5d2BkAmpMpC0rWwchMn2bt5WoEK1u5lpZW
GW/xH70lleeLA87RTTeO3ufDrc8BTZbR6vHw1aNl56/l5axbXlqC1kcZJqhcvWLn
Bk2zE98/PL/DuYjwBguBGsiax+Dg1fg/n4sxm4ekdQpaHO5/jcIRtP0Z9CawwQ7C
KsXEbOcznfpnvAx6cuHvBKwMnUAiJtYB3dWTJFf/KcfZfmCBjEDp7mBM1e/hq+TC
izbdh72DSmpchZjZMRI0yLHloVnVHAiiyFCoumH+UYQ95//MVcZwa4cjizvSkAKA
yHE7IquZPNUUBixkbYnztXOQYrEC07VFCiC1sRCwUuLdF4Y4WxGVMXJ8j3lHylEB
hLsTL10e10bVC42uxCCr3Y4d3iNO3950PDcHZdT9tS/LMSb+RDLY/mUFGa75NYRA
gSlDst5N8EW/wJkxYFeizZOBalLdouVKP/1PAbu+2QdLtexP8WoE6bN9nSy1zKgD
WBe6Kma3ci/VzWP1zj96bEZwCPCd5H5wNaR4OgL8f5sHysr7VwNEK3LRvBOA7KuD
iSGGmiTya1HQGYAWQzIjrpFTZTz8YXP6kgbgfu+Ey8jU6xprior8HgjcJ35Kw4Dp
xn5I/MTaFFsvaDfzE+wixM23qKhemYMqgHprwEuShnrZiC62Z8rMFfILJxp8mw9W
Fyiflt9E9xsgAYc/qStsKGXbrpsYv2aTUkmwfFgOSvinv5LPpVvrzS/bpnSbaEMJ
62PAK01EGwUVS8vAv4INobopV+rnVTlEebqVJKmAey43VddF0eg73UQYwd+KTb9V
PKK3TVT7tHefdXWLyqGjseb68GK8gUVJI1bnw+LEUL/b6QSClv6NAsHDSHDtTH7y
1J3aQITlhYRfVA/WJd5o79dKVmwLGe56vAbdeDocKFXQqNnCOe7B2vxis30355R6
1LbLivQgyLAkEozoFkuT6hgcutSiR0o5penVpGg1e7Q+MnILQq6JNtW57JSG9/kR
sqd4HIfk7aWpJyX5Gb7DM4RiO7Z+HxkqP+itVWbwlnet36n2sUCYpQX1HutJo7Ky
xtRVbpaT8g+PzXyXw/EP5CvMLtTPhkaWvlUmNYEJcM3VHLPl+NJ0bS2Xtgr44OZq
FrHSLtpB5Ff3JOfxN8IQVNBDPwD3EgkEzo/b7HXYUWGcsxMrTiBvqhQuuLkUfWb4
Ob/7BXK3mbPUwvMr5+isWTFWAxA07/NE7W+uU8I2uWDTQ5fbhVyG3EWTkWozGxW3
zv3NY/MVxkyYhR1ip8I6l07x7JqAsuYmqhCd4XDLLNhYPEkSocMHK5yXYayp0+u5
qt/se3YOWcA2tD0vvb8gVMTsPKF/I4kYdYi7Zu9Bnmzh+3Sn4DePHL+2IBvFwgHe
tvRgUjHQje8J+Q3/lu3vfVd7DOF2wtfJGH7SeTh07pCr4391zCYJqb7q4IXfqoUG
NuuvAJhHTFVeZ68JJn56JMK+D8SSEv+lnCcrpHAsbEWCA6YKtqIX2UEIdGJuWNMa
D11GpQdkz1JhCPZHmA482eN0a0JL587SRzGRRYmMqvdjh2ECMxBCL9B1nMeYLstp
C4Xb1S9E3Z85WA5CFR+sFhREdDUmUttrJsZBqq5Pvc0s1xz9iYU/ydquekBf9YQH
znjzAxG5DIoOko77zEj2vG4o6kIiyBUJqXADjWF7TyGLkW2jcv04+J9fXCe8t3kS
27zlR9eFZNcFYpxDRdJ198/cqZBjtPCXdH8zic2h7KBPM4etz1fPhcekLSKZBz3u
Lh5V9THyhokblCYUKAgXbWTZr2f0RdjMEg6jVfcnBhYM0sGLlO1fhgix0ZLOFEnr
h6imHd7r0U5NNNH1EH0hodc1guXzMIrhs7/+BJJ9LfdJcpobR00oWj+Gsx4DLqNf
Qyqpt8eGjr8s7yLjc788pLg1GVMP7hYkiwBevcKNOgFwqdOzyqOxYS6B2v3dQz03
nskVzDTZPivHY3TsmtSfZPivkoO1rWpPkXFhD2xOYR0GubLoycSZ7gYKywOzemxP
MEU8FR0MOuABiLvTXj+qHL9+QRo5aNKTdrA3vNJ+Si0UpgusT36ucF/7BCWHHIP0
8eA9qv3RuNSGVj58i3jCe179z93lSIiAcE0IcVHSkeeJA+Uq5vVHBQOFY4ndjhcL
PLSe+3prmdHnomlJCLyOM8GoUcYGjBeLaxzL0AXLP9ktbaINAIZztLjed4H7OnQw
krOOyOH0GZVfXhVr4So7NNGGYXJAdul36TRxXLEBqk0SYEqQAoGl+x4lw79Vu9xD
X4KOPiWBlw0pgrAMnaaaD0lWZmtGmc4br2l5e66SukpQIoaoGYkplxBz3wPMNh2C
v8CWYMtRYFAbWTtK0zaARkdLtTA7K+dD1YoZfchrHmqa0WKY59pTvDNCgBec8iO6
lf/Y+GIvdTcnAE48peOwdoBfNIq9ouLkjjq0oZh8mo9RmoxHaVFx75y6o4mPlsi8
eGuSaictykZZV1iPuuVfhjf3km9WAP0THVAkqJP+Zs1s9w0Y19MABzNrO/2XXdbr
RISzO496geexSp1EdnJH7GfZqrfyqcXVF9l/Oqm0s3C6YEn9e5kfnOFBEow+GksV
v6zcZGrg9g830MZH3sj3bBgJyT4xhRo8nJKjAegoLQshGi6l1P98JxkjDPl04lU5
CrOld9G2TuZ1XX1E26B0tTBLm8+MkPz+MRCvlpURu0cGW89GjoYqFUFFto6Y2XRz
Ez9CItSv+sPIQRhFmeCeNKClwerS2byjGoHINwLoazwfyA19wsp2mcpfHwZhvcE4
WCLqLeBo5H12fSvYulqRV5xxXMrrlZsG6lqjk6BseMvMXXQ6t18EddALf2TDWHSW
7kvK0Ty1VxU3hnlfvD579lnrGYPIZutR/BT0KxiytXDeksumyEHPz7Uba6EkRLp0
+4MiUCU17FT9p5jvmxZifRxpgAagICBqilxMv9tiwztjb7JYpPZRa+GmWBKrCpWi
Eb/TpsmWk2ZCzx91c0c+jIoi1WUKOgpOY+AmmXe8WveX2AvPCMgglBetzR17DUuy
2Y3EsLlveRhZIJ2f4VM/R/g2WzfgQI3JKioq++HIm9y3JOfe4IX3AYdiXeVvOpdt
lfy5lyRxZL/jeQZqrenNdiegQRk3UIsJTzXBsRQzsc7Oy1/XytbQXy1rIKyBCmlE
yuZ9JcxqnNyWSuugx7KGFQVnYhAwDaGurlGi4MiAxa+qcw7jQywwFNrQxoykFq7N
rnWPyns/0Eo+6t8CYga6PPlX20AiHjtIZMLmHEFv2y5skNKGrtMaaP0ePwkgZP2N
l3JfWezOEtRZaxlPKYnrv/4N+RRqx3AAYNBG46qtu9iAUho6gzU+fXrRJ9UEsOIH
a1DwZvmqxb/HWLnBObBMZ/LMxXlHBnue583s73XY/GNiv/p7/lor5SPdqmEcnibN
uUyi5O1jBa9aBx5jwaMyW61LGUrFDgH1RUXDPNfD2w2Ts49oO+D85OvwV2wRLWLm
VUZgTlSCXkiVFmMT8Lrw/nvefBLKhzGmSgiD2OG3xmcwxVIKIvjmRoHo9Wo8uaw3
4w4j+oxmYMUYeBCE6M74eFhpDtlXorxAbMzjbt1H01KCV0fIaSOr6gmVZLOSbu9U
io3bJ/jLx0+OOQl4hQXRgwvcWkKiP8/twtOecUP2G6AMULI4ZvBABrWAew5+N/TB
Zp8381Qe2owHx67lXiFVJ1CbcO8Lnchcfpv+TxQfVvStGyrFCDzUqfq5sFqKIWur
xwnBaeefdQ8BIeGa5sadkk0Eqxef7zSEzJcrNrdB4feQYS5gRY3ZNqL0+B35991R
hjyCCQF4/M7vuknbADNI9kdOWJvMkVbex945z55cdy4IYhYMW/5pi6olDaYCZ1xS
Z86aM+sOoIYJ6x9Y/0hVCqw+1L+z0iR7JFhmVg2ApnkKdW1yoIyXrWBbjQWHFWOW
8KOiZrfaI47xD7kQS+IEvkXMy9/zJnHB9bXNFW4rpbfV0dLlWhCM/KWXw1No6lBY
jIuwd3TaR1pVtcREw5s6b6v5bY5MFsJDNpioaUqEx7wjTAYB5d837VsB/StW2by/
BgSpe5ViUaOh2RSR2vY+vPmu/4scAAllH5U9dQySO5XYrZ6vkLMc8ErM814dbymX
kyYz4d5x5ZsITaJZvyEmUFrNxXtNyC6wcHLt36pE7ypGIsZvlXBKSMfXbr5sZ7XD
rW2v9Hhc+IvvX9X0ke9iCmmBt6E8/SnhXZBOUQ8tK5ozC3btzCgGOjN//ipqFsJN
5MxIMdh4ZzGvZng36H9QbstjSWxOyIohSzgfrNdpn/xRgyNQIQYJhW+EuyAbYICY
5cG2uXgD/tu+fsCKQ2uRaPRUnRqDY9gWljgtW6CpzRgn+ieezc3Y/uUYerDz8g4S
iTsIjHT6YfxuhXeIBxsS2ZXeXwVPajSMFF6B6B4wWcatgoy83KMw6SrVdyXxBdVw
EQsV0Huk1q8h8ai2bjEv5BkvzSSEPviznDKDASe8kvkelTvKcnG67bklMlw8EAz5
LONwf+ZrVuqwweFmV8kNcR20yX3V+ILhnxpV+uONQnr/RA6npojeL9MjEiZFw4IS
zx9Qg7+5r6uLXlKis42LGpBhcZk7jyTAphOvo4oglR8DvcJ2MPGAx/tDW1wb8n0R
AWT8FnVMScKTJ4+p41DzXhlf6tHrlTasTKN6wTuY+p8X/1eW42wXaMcZdABc8tjj
hXjsM08RiwdVqRh9H65vitOGh+VhqY2hIh8/u4+p7IPQ/loDcDuvM3nWAg5vAeDd
oHrSmjAbSpcP5OxKL3LlaxGYVDwgX4IhqLJDNhDLSUVLHpP1BVR6+ESsUiwlQFsP
4kY+RNJ3dUCDN/7xmTbZjtioxX2C2tnhowETo3zzgdPGbcZejRjrZmmbnJh9XQa8
8wMwLsK0+7May9QyzE+lih56H6Nsichvb/OR+opgHpzM9WMjaik4/AayjrOAElDU
/0qgJ0YWc5T5HpkjRKSXWMlGJqA+z9eiy99AqW4E7fwD00whfT6GSyv9BkczI72A
4q7F0t4Q6rsPbiRqMXlBKHg133eCUvY7LcDmaEJMeCEy2U85cCKkBcWa1Q2cWskQ
ZpV1pWF7qJA9V7/agLEonFDGeZc676TlTFzECtqfeLsV6QZAm1KeKy+jMb1/N3KF
AS8DDbi2021VFdSpOXte/vRu/n8QQSFwJQMcBEMy6by6zZj8ReiPuiKvKzNxgL/V
BsuRouA5oVH370pGydzMYy/MVy5c6Gz2G3YJMoZUqZWfEGjd4fYcNMDNdB51Svq8
uZ01WzbQgEMvkDFNYfcUZArYpoWf08cAb8Fc5pKdtKYVKSg1LSg+5Rp3+eUgq3Aj
k5PdoqznjHMfrdEPNqJ6t3NZnEWa3jgWSGZSaKIJ2jH9ACvw/M0knzn4MtzkWm6b
rgngO1uHJj+/zhbPYv7ywxZJD+ozmaUh3GmT2M1yeBlEB26v+zpYloBI8G4cCuAW
WdUbY2VHdPWiRaTIitynVfpbG9s6HMfX3beLesQb6MYstYtf8QEEH2IoHSP1orjM
BK03mgf0VmDo/WkUzUyUQffa9Zm0FfJN+ulrUfTPZVH4+w8wXrVMJ4RQHpDcuTiI
rzP43Cw8K2Ol9dH+cmEIPIxD/8za9H9MHYQWHaB79emdVQKPZ0wnRZx+iM+jKm3x
nk4p3lFLjEhV5mN1v7r2ETkTUHjxQmE5fbMHNr3/lOoKCTvD+EkqtLOplAXmWea+
a5rSqSAAx0kVpjhUk0m5ZGE7g3Oud0oeFfvPgBJbJaxDSmrqmo/2R/SsaUBWmLxO
J1/IuXuYGOfaUhqhrZbfTR+rdEehrJYFt5KSRPC2YMrPsFBdyP1U0fAAf4UcKpN0
2UEhSw7onSFlOqaG3NqSAnMhPU7wL345xy7nzL7nsZJ0ewos7Y+1oylVYH217cWz
xUW9LS2nscVYMObyW0QObWfx35JcFyuaWiZ0970Q2tL40CsidS8/tzamwa6bseXv
rWmnwGgBAocvrU0N+VHJhtuNk4xhs2lw+TKbRWemmB8ONBCdXbIYOXpWp36ZYwpM
p5uUGxmPNKzxjzW3b7ehv70tH/HSTrqJo66acRdm7KaovsP0SagOmyKJVij/0uAF
diBbX8Gf7SlXqNrS45qPgltFyx6rXFyEx3Owi5uqbbqdTuX5vMkOaca1hZ4FKF1j
ZmZsJVnJfVwNjFfW/O+BHLMaR1NoHT7+iFopjttvy0m/6kxPuj+32BYX01dBWlOY
n+s2zKf4S1rcpUdCtisCUvbehXBxGcezU/qpmtkgpEw/5Gk82e/GPBa/Mrr/7MS9
RPhTXN02S8CmS2RyXJBKn5Bh+q/AhvjLURlgv56zFyjK68hGhNXhXgNS12TB9hhm
DfPB9ENxzq40e86p+DVQ5mlzjlzpyf3xPVu1vr1wNhJZVhMhXRmUDTndQPILUIjd
8lZGBcFSZoxN2wcgoBR20I3krXjkEqfnPSEJ023I4dalogXWORNO+5zrmoB8r1iC
qaHtVDU39lEdZoPa6ekpJa8pUSU/SDVgBk7aQ5WMYKMJor1/3J4B2RloOWPu1PYO
Xyhgxw6U1SVV+22o1H8ZNl24kZ8V+0CkWbEmqMVkepf0Xowvi5reQwfcUImFkA+F
OyfcuWSRxtSp7pmQF70e8Zylxs/SChvtIfKRxtmKC7JI8QGjAT8e3HEfGTUFGBZD
aoBIHLrx9BUcdyZFP5/Q/51AsG0ct4lboRpJQFRxM9MPcqCSx2VuUwbEgd9RTeHR
MamoAV5VG8OYq4ZLNef+RceUH6lL+fGk9ZEjS81KGDVKKBj9UjAb4Os0aW0OVe9x
dn2yccKFRu4TOWCJ5rnTJmXFSZVuV+1Oq6Lm/nfKbg/lapIzWdrF14C95I+le2Qd
P43wMqCjVWASGV0QIHNZZuv/h0886T5tUlBYaeAZZ0VjWthrlHmhtb34ZFtg6n11
U2Qft1UV+4xIdOn1Z/hLj5b09naLmblqrgZxiOpw61IoNlAnCRCAEhzFYFTDtuf1
F/mnjkVgWg6VzJyda93JuRfh3CKAWCpt2jdcAfPY4IuBU/zBYxs4HnCEo2ef0GCS
ElvzyvUPY6NJwIRm7ZjWTrR2qo9Kl3HH055/4AAzZslzY541Qmc2XaA/FxlEmAYv
eKJmJo7/z5DmsVtQZ4AY/LbchwZobTG75jdIKL9Q5lYxvupbyGx+TOejzbwK2Qtc
M99g1sV1aiJaDtbFdqCyJXrVam3YEwyq3++PhqUC4rAs+Ny8KPFob92HnMLl13Fs
PYjpI7r1Bt66VwMahv+lrvb1f6XgwB5kHvKGm5ChssPTFOUj9/UCB+Yeunkog6EU
KzPaM2dU6LcdsEr1o4rPFO1vYRnl3ntxmF/ULkxJiNmUpKKkFb4gKRGQGHT/EUBx
5J52gx+hsJkIxD2fdpOHjYQgjKDwYELXyrplUdqThMmtKtumuykKQZumnS25uWvc
lvUICCi5iaTMjAqquQWlvTjaMo9O8SrOSl3XdnO+0XWJ0n6FQ9VlFkKpZrqIFOY7
dRRvFRoUbyyzjytZuPofs0IFbS5WohO6efvskY529+ht+6BeZzororLD/U10GyA3
5n5Q6TpbycFUrOpY8wM2ibT4kBWmyJUhHU7Ov5DvkfaYmE4to0VYheJUjiNEExJ1
5ytM+BKH3yBdIUcjmO+DYh2pqnmCmSJDmifdfrMTzAp3JhF5516Q9GpEfjiQslYX
R+es8F9w3T3kxVBXlK/PzTXBwmpzIdQoGddEG7AsLBAMRg/WLrThir8zLc8RCqQ4
ggOdB0dOYiXUKLANX99GeHFM+LVmvFkRMCU18s0S4TwBSW/9KFggoAVGSBjwnia3
4vmCFEl+iWDt7Wyx8Myn0qhWoBzhujGf1iUa3d5jQQbyGbc7GK5GmFvS2ffKtjBo
uMBX3jXBjej6iK5aLpGIF2dbv1bvS8Cq1IptEKLshURwC0ve+VYpzrNdDvd1f/Ny
pTSVpCHmyh0dQK30OpK7q+V+jePtZ40YtFrYpuS/kwdOitSzmyaJ5F2vDaPDzTli
6KcRs0wzOkMK0GnzBhKw/KIGVREpFGhdGmEIuKhZJ9GoCOtZ6DdNa5ToG77RgNmp
JYUgDrfvLhFTjLYZtR0dow6rJBorEiMjxBSCVicpRzWo+1P68w4UfX+GY6wCBdTA
9t+mqdtt+0FH/jfYvNPnd1EUJQ3WI3XHM5JOq11I6G2y+7NkgnwSgZ4FMkzzdX+0
VhZBnPfCZlJUs/fwNeqm+Y+k+JxMc2eZsvt8e03N5rssNjMYIx02PTIH7Xtl95hl
FGV0iW0UD5JUsYvDg2PkagjIqxoZFngSu4g4Qi9WCUBA26xRZ/9rsV4qvXdpoaVk
l0cIgDc2SVYn+R5mMv9bKfHUFfxTtceRVT5mLFLM7gqmQARBTqT4J1gZSCPIfD71
g72mTdkeUYjdlwrQFjhO3UGhDQ2U28eKa8reJcpwFEbQ2egcaSwu3eWY1OZlhagA
H2S68kqZB8Qo6DNItzjL07HNAgxsZ6Z8GbFTGfi+0hZbmBXrud/HgABAwLQYJQbI
KDtF75zbapY6ALiaZ1VIa0oZCTEtgLsUwVLc2Ez/FC696tFje8CVyUDvQb+LkgIS
ZYiuKGz+L2jKTuFWc04eeM/Wn3wYoVpmCXQnXSIj5pI6hVjsLC3OOBCZ7h24YQc6
hO6FdtpKHL5FFK7Pf7mkFBODjSNHQxVFWAWcaXOiMm+KYuvqMUJom4rDvrGeAQTZ
u/AUTWgM8eLilJQKvKH4JyEQsXnqDNE6mLHiZkWeSzK5TC+B88GFX9E3f0bprpCM
Q6o1jICINEHe714tozGdHjmlvxnsz9LfCPUAgvR6YQ4aTgACC9JYLdqWa3mTZodO
WD6MAUKdVygYKJlKdMTVgQO4PsIASTRfnuB/HxlaY0bTrHpkB5sxEoqaD03idVuU
9e4eckNpEusFybiXdRAhoHN7i2fmhdiYlHyVTTxgWbweg2hZoA2yurTb4CtokCxz
nTakoelJ37THyN6nwu5Of+QfOzm+MWZDab/qLKSx8FGKod9MEX+D1nu08WBMYHLt
fZPPj4BbNfudIYW36ul2Bka3TXyEp7kToJeLbZx+grA7ZOOMYhEgW0gCBQoy1Ydz
/QbnNet+YfkkwgThK1i/Lb/aM0IthCm/WfJXG/ok3lVOIm8g7NokfmaDfz5z627f
ljKkFOecnSSgTvVBIQFdCRvLUgGxb5mGurmDxNHM1d0QOFa9Zc/pA2NrtdxbHqmn
haF7PvT97jC88SrTHeoU0vSiYODCVLWkInUnpcr8fNxPQIzIY5lgwLsqcIjlBeak
Nj3LX565tx5M71xCkjPQltKk18BEzorb48i122F16RkQGgBXVzl8JNUDNRU/F3iF
JEZjjEJteOnC1R5XnlKI5vLed/yI5Dj6Nu1Q7l5EaibV2VBNlXG8+AI30BSsIzj3
+qFswU5HjTrvQwE5bQe1zyRvc5ugel8fG70PC2mFGGfVh6vIPOo8vrN1Ml6HdRxe
u5JpjcujBDn+wLm3k2J+CpZVwycV+aNAnp7D5HBT/gjRdAS3XXsK8HRdicztw2Mh
bG8g4IyTBxuLworvpfVwBfm4JC1NNbRlpDpk8VxsxRhDCmwXK/mY6Wk4LOWpf0cL
1Hu1bJSnZN0wOjxJkT3Y90+ICltzmVxWmqP4ORgwkcvBFl8zrZM2h9XekGvRBHoC
Og7kyk6pff0uvCbpkhx8hGtMjQyDcOFZO9wZIQPGC5BnIeLT7RXorhEbGhFbuCp6
O+y+CcR2MLBJlXP48t4p6xzZqfHtBbM7QAwERobhGgEdap2H4C5D7UyHmp3tQk9p
HfrYNROJLUPEzPflna8r37fFUssia4Hf3DOSHFgiBmsrmhlBLxEDs90CSnedP2he
KHyRhWH9JElMXwpMLzUGHJJC8x+l+APqdHyx9loNII9uGchEVxSf3OYeeUvAjPZA
v8SjUotA8bKL37gjC2Jyy2FDTDLF31m8pt9oXW9z5qkPynTopTOeEMrNT8hA6xi1
DDrdz3KSAHq/RXrxEey3Cm1zWAL5499nb6DKnWc8UjiSd4+qkz+1azhv6fRPf2z8
98r+lkPXaa+iMEziqLmTdQpsGr8VCioahUO0N3cvI112E23gFVmPia922gSuHE0W
742G5zFOJ2h67uNX7tUp9Ame9QG7+QSZ/vyJUCQNs8QGx+NGxBPR5SMTSV92/lF0
s7SYyVrPrXiVOy88vp+IqCHp/qK8wWUKsXw6GYFKiPSD8pw5qR9uczU9dDkxE5Fu
pdVRdI9VhR44LyozX0iFKC9EILykIB7ExpcCy0NO684NY5iRLBlgWNBRg8TmvjkP
4WwhKRhokf6d3Q4Rg7TzolY9Sq/WUyICm0ZdTvgmVNN8bi3nuFcbxo9h/8Jyslwn
/Eu6/a4T0/K5mYzrYsP3qGii97A6FeW+jovW+smBVBSExsI7q5AN3A/rc5PE3cBI
CxNSSYL8kd6iP/ZLVjLpzBKAqL4c6swpjMCf7eCXAhsPIfFUFoxjXkiAfk8THsgB
5lIIpiL4uOZFXcACE+XLFNMzhaS7TxfbvL5y81uPN3ir91F8KEcclPV7uiqtueX7
lP43HgKyGLRzdgpPIixTpGug9gO1pbtFg2wuUFfiISJUZL5KjvY/Qud66eXOqY8Z
RCIAY5P0SbZEp4GbMFuRyX4M61fRyCbNlI21STIlqKiRzYtDDvsTdxVINfwlVK/c
P3qABGp/FDAlaIu4BRH/lUP/ORNBgbtRXfj5HR21Yv4s36HwuqEQCqsHTVyY8uSc
GuWeYsl+0KgyPBBMlmUQkpucapEc//ZhIFYHWym4rw91dttwb78EdBp+wprOLjEt
As3N27i1/eSr//bmHmZ5G0E0LxT5l9dZ/J95DOMKP3FCGM2ID80myniNia4MysAd
PjOIaduf5nBfgoNlNVnqCYkSjJ3QrPj7Meh9/aogoXesydqAs3CROE2HwP0jZSf0
trkZJXsEAM1cTUW7QVKazuho89t4dXxh9o+rHByKR52DYwzzrplL+pQuFTqI/KBF
EX1spqHGPQCzJGnxn4+Ep9FkR4zWoMWsaerRze2jJ1TjDxE6xBDrHpN6DXZXp5h2
mH3XdAaYsL9xU7DOH91dl21oh47O8rap0F/l1rDkcjh7F6Ss2IilzThMg8wfTRXZ
`protect end_protected