`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
j9eMmSPGcKCWAR9PvkqZ1R001FU8QKTyJzFqNLn+qur6INyYDE1AI8LWcxAzfnTc
IpZG7ua3uuk5/kQKKQx8ZIPLfmv6H3t3eWjki8YIAtY/d5E7Gq8Z5mNxMYRzGGTg
TCMm6oOrOTVYlCXHE0X9AW696Z7UGfWirVibl8hs19hrFdeZKGiGht4r09vHR+Gl
FQQmSObM5aSK5wu5KOrK5ZUKGHyBhjnIQO5NnittDjOwxV/57nHVg0pdG6JUqyvm
tEgmCY36RCMRGWN7sekPtNHjqpZkmYrVX1T9QF3h73+8ZekZYd2xY2hpHHGYYeWA
t3+Fmb/6NUmoP8+Pt2hI6g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="wX+NBVcG/A5ruHK3pkDqG8ZVPdOz9TJPJ5saXZYSeQ4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
j/hqWUoxjK88VtH4QmjIrexFOSwtsLKOZ/LCP4cmrqgzmR/e71apdtoL+o8nlfy6
eZxDZMmrZmJGoazz2oK6kz7xJU85UCwNc4cxAsVxNdCP19vZxph/nCYZQ9lUFkLH
uLBkOeFP15CD3jG5/dp945fHP13J9SzB/L9PWvDC/gY=
`protect rights_digest_method = "sha256"
`protect end_toolblock="sqDZkaglKf+bDjC7VKm3lOELrT2Jlynh4UhPg2J0Q70="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61520 )
`protect data_block
f9kZDbPp4NLiAOFOgATj9W35i3s4a7wbt9jeHjHVcJxMoXY8rb8laqS5bNUhXGW/
MOc7UNc1VwolqhkS7G27SLamkGClZZtXSbRcN1N+5kZpEaBEj1343vVznnU2Dre/
WS9HsWPXe5g0wH0AJA0FuKjPl9J/xf2fBf8sDxx6VWCRRugEK5N5v4vmUIrmwFin
sWlkRgjqGZyFXum/ADIu1FJZrjXRd7YMMdMSGWqTJmksGeNsSZXyFTAuRVt2fnjT
8fm+4E7NlIFcWDiTaPEe3ranwJCsXE+EZYQSuHJ8NLwwNaXtD9zPJdGQInHIZpwA
gs8DfKfKCp6aavsWD1EAA+dBVH/uwjXb7WvQPu7w4qwGgqVe1YWRmm10bomXRWBs
TrDydPlWOoRsLezMCVWGZGm3OaS3l/3sK7IoAMInr+0OrCkCTX1nqDYvSpmYKmMQ
F/j5akWZ9qW7LhIFcL8MaaMPL154BLfW38owzYxHdLdSEFd+fe9bdWw2Ky9B6Npq
eT+FMWliqYly8vh91LgHspLiZV+HRPqYkWhyOjc8CYiLRofv3jYVnxpttJ4EXavt
qPmgWkpgjqtZ6szgZAOVgkk1I56lsDWhuKyucyaJJ97JHWZbF7OkXNFI45nPpYvx
0rh79mbKqxXVGM1miHW1kISZ4wMHM5vsRcbeznjJtCFBI2TbMQrkwo/809OW4uPY
oLH0XsDXPKiGcR0aQ3nFC1xtj2hyvcul8GkfgLUcxQInhv+mc4wwh1GRzUbryXd5
zyezy//+7B4JgSP8yy5f0qCXgrNr6CIALmqRFUr6gF14CAooevfQ0JdB2LFFZwSw
F8/VBktDkU4S22TyZ8x48dHxLS5glGAtLVn4uiUv6KU0D27IE1NVea4ogPdpv4E7
QPcZpbt3/FElMLPzY839Yc3CVnh/9RuaQ+u2JQtQrFjPriOM8Zrg1Qa+UHDFKHb7
p3Amc+3oUNeqGUrwRl2zrxQgzG+tuIJMe29ionED3XlzL14QgwuWBGSzRApL73Ow
UKVUnJDPw5R3vtfnuwe7VQ+TVs8jTWfN/lW9RLqfS7mAI0yqMk2cFkvJb/r+yL4b
fU9VuaeF8c61lAhF7BGSh58BWVzxPtrnSpucm+ieKsQQ1LU/7M3OI3NZGxh34fv6
tzWKDjEayWYXk22R7X65knjUTcGdwGYFPP7cn8qX9lZw6vzV74n96t2/fJFnXYeI
esad+lp/8ibcRB22WeHYoh2JVZyjtnOEv2uat4McOJwi1m1td1+pH/cSP7qMmsXM
NrJiz/j/FpOGAEwl2kEYoqERnc6k9Hth0MzBOUFPgafYUwidSpbVzlHGHV9GJUso
vNyDrl1OSxkK1R+fd+eewCaX4KqcB4rKi1TcsJVrEuKGDkoQvK1JFT/ar6ciLoAF
raqqwX+6/de6aYBFD+/Vw8w6ld5uyst8FSy34IjYHU/ytknkjbfkqusrvbaBC0LV
PpL/YnkNY582mCfMKAnZOd9G53gxquTHJ1vL2eeFQw9f4olc00ngPtNzSXxkhQxW
0U5Ztiub6u3T6zB9cdZaLMzAI/7UcuL4Gv3kstnx6PiWXt9q1SgBKj8NLFkC4YiD
VpsBJsqobbA5jirb2aH5S+yGQeLfIq9Mv2YsDe6ZHT2/RS6NCoQIIIKSoXDprWL/
9zt4eFNQ6vBae/fmKo/uK5ZaA8IHrWFBpBHh41XkgHUdyFOHf75U4VYEFrO5xqg2
4sm135P9aZHnJNH30avMCAFGJZ02eZCFxp4Pr7ySelrvbojdvVgS8SG99YbnM368
KsEHGaf/YEKqy8RzloJPGiPENRXAaNRS86Pu1Gv51HrJAekO7ovLfxUr1h3fAhIy
ZSVuIgM/CO9ek2Z8bfgeru/OkpzItyMuhgKIjjzRQejiEwZ2+etJN6J04J2WuAS5
z9AGDjR5ht9jPJZMApQ0gWHFzYytz8Kr4QV2PQldgCFjdfxAxfn5PBSzPoWVsLp9
t5+DTklmnHqGJEA2N8bKY4RB3E8D4OGFJ/Fp7ab5nTKB9MtOtzq+OMH7m4dP5J6M
jIW3+NF/orffkyvUgj/miHQpDpmfFwVg4t2WC52XL7hSJl007fuXF7ntwJEahfkj
U/KXv7Wd2TQDtQfrrpNrL3R32WgQ42lRbUQ1AHDxwwJ1nJ46k58I84+jIMA39I/s
ebWr3NGqeoCJqn83gjZNxDHkgjE1jHCaTPPKYDJk9pLcA3o70OE6SsQ02fKfXF4p
Lb4l0ylYhzOWNHwE1n2/jJutFu8Acq1EMlPRkSp9xNz+1dklsjWmHWakNzEfL+xg
CGTausNIrEsAhWeL2RP1MFS6hxj/5tbT3nXwrfTtL3JbMToEPCXsP4kh+9/zOmwE
GtE0Y1Jo6YZpTKmjSo10tjtU8oX1k3GLbedrfZI9uxHWiHN4kdZXk9y8miJbr4pc
Ro2UUr30FP+G/EabvuvapJ2Ms9+wymzcwNhwAKPifDtC+/A65HjgPRtmAjwdlA1b
wnr9dd75lnZNjrGfRMvkc8ChvWalVumg0U4vou7CuDfwgJ5p3c09RXCozD5L1+Xh
oQV2DBKNblIlHMj9oi7huFkOMDliPNWsKUz/nTjBTuRoZfJ1lliVF5zjtFbiMjh1
kATssMlgjqOgUO6bkDZGQy27uL3Ad4jW9ZWYtZvjt2+VOHtgoouc737jFJZE8qeX
/md5fDZg5WQW3PYtQmCDboNRuPMSXcbsZ3nEmpPD/V3tVBJznJjfxmnC9CQA0mKp
hvVEGvvZW1fddW4UDzrFwVlT7BWcY+3n/gooovzeVimv/7ryPLDclPbIGWRYBvx7
THCj1SEcKliebXGN6jE4RwP6d2PSpvzoaq2y8Nxwxne5/DhQYUE8T7yYdJ90rIwC
tUlBCK3/zkSk1eECOEPSBzMDTYEDiEoUNG/PetizWL1W67XcjSXzfED5WMYGGJ7n
gfO/UUGk7aruJiEa4KKBVUwJlijAwBGlnKQ1ShwwRyU5BqSfOLQQ966154qR5NPd
DCymET8FML0qC+I2uzK37A1j8wllP1ijuNG7iOEJ4ADWwJPbHYvd84nRImFNxKyS
468jG9eJW/+c3K5cGLyzfIDtMKdLrCS5Ruko8itQLqrlTHtT+5IReK6pVocpx1ER
DuQ/qy8GQaqU7wdPlmEbcXt7NvXeDYPpAo6uxSHn5YEm1eVwizSOkpgLwzvWZ7Bk
AZyTPwlfkZgWYD9mbFp49T6FSTO5oiJcYVPQExdeZ8FrpmgTR6Det5XLsSvYqlO8
lyIfMzriNwC2VrLL6ioNH4eb3V2CoXJW4J2pABoOS7KvWNQuy3PG++ogoCeIaqWw
MmUuAKTFYm3tXDpsGMMpVVfQ8h0bT0xR0Ghe+IzVsD7OXLYIvLsnVGtLfdb9sfLD
992PUCr9mRhAqsJ02YwVp/km7Y1W62aPELDEzl8y6Z5ryrn1CFTn0qEGqFLnFsjU
B7RKCUbnnJNEGS8ZPjplUiNKjCMV4RWRkcatFQDUKpqguT88ECCXkLTUn0PGilku
maiPEEkXuYKmw+qoT2SxhDKj8RptSMUb+tf+ARAl9UIxhY4WrEbaYnPnzXfO0WHx
sEwYt2xPhrMEB7o6Ci+zAgkzTG9+dgUehcz8gB3YhHFrwiJaCYlEbkAzy88NqiVZ
ebSejrHonZyt4pcxpfennSqeIoXc/6yt8dZ5MEUWkNPEf/+qdz1a3nNGGQVoKR6Y
l4b74mlWnNYPMz4PiDeXYcVm8zjdoztdUuUEZzGkPUyMH1rMEMdH5nDihaCAtlRn
ppZ9HC8cPlKz0dJ1ZIgzePV/YYgGfKIztt4/jaadL7AFejx+V5NJ9t43iUv1jMgf
4FMaX9xXpEc/7z7V87kkORuN2OJ3L1Sl9l57SHktPEY8fD2qx7l+bJx3O+CB1O/O
mlE4gaD9KwcQNP9QNiGu+jwTFqU2MpuNTGoafEGKPQmpPWzmhLyCKbK2xhXk/rcj
NTlplaCNolJ03GPcqCocBGxFAYwwxELuMQeQKsMAgq0dIrqykgy4HkHbY3PEQckg
/Yvj7R2QQAUlgrEpkScju8ucw1g13xH4gXCLZVbticjOwpKrFJFKCfLVqO3+m2Ys
SUelogNxvq/2dCf+t2OzNm3Y5WcIC0hLAvxddh7KLA6dsC30+In2uLukR96c8sH8
3tGHoOiYJWhIzZmBQ7obHgKk/A0S/QgHXbXxhKFuqlSgYEqIT2WwQIKN16dYo4Z4
1Oc2GEDMqVOQKKdOl4sbRpnqlKMw9WsLx9zCDJHmEw/pDcNwMXb1Q+WNmxblq5Lo
6eS88J94WcYKi1oMFKIfFkYRkBmd+9eXO3YlNWy4w/g/u7Z9HWktqQN9IngyUBIH
gm49/YF4A7Mbo0r1LU/ab2YR7VCWqk701SrcNcKtVqbrsX9CidadEH4xEeRt4w8P
/298fzaBnkd3DKdr7odrjibcXfmaK10e1ZupxU3DUiH+TYvqol/VxvULiStsNAHF
rM9mnRX/MxtGGBwJVfa3y4L9RBp7OFEt9nS8DYcoPuLfHkXU9uraK5pMCSALhpSv
NVKD3SqyQ/KV0iwIuUPRM7cPzIT/crEAuYJQmxSCJwfjNNLW67ADYU5/duA20nGQ
33rw7asEOpsL4GCcjUW1RhAcv+mgQlzgB55jxqMFyRhawcZccNccePQTjvEkIz7n
/u5He9gADJlmyX33N2q4Rqn02yA0XygQBf1MxNLsZEJfC5fxm3px1NPfMVUxgOdT
qi3Whg0mB9nbbGGgHGiQi/MpeZs8cdOglblQwLz52m/J4alenRDjjQczyiX4aC1+
iqWLbfpIAomAk3iBiiQGb2+c3oToJAAT6Lux9su4hPSq8UlfofElrLddbD38jQxe
6YUFZEsCu4xMAjmMXt0bXchHFxzT1oGaU5ayoDXOgZdF+6+lExLfBf/aLs28ZiYi
AUJbxSdheUfXMiAcIOmS91LKIOyW2JcW50Xje29sDFdPABJ5dZnQ6r1itehK+iic
VTUseV8gNafkBnKfPpVuGSul5vCkZ88E85/RMN7njBEu7K/8jx70MqHCyQYGrSOQ
t+kxyI811EhqGT75Y8ptq+d5Mz5XuGHcBPt3a183MvUjqh9/OFeRGeqZXUz+6ytp
wkg+94lafPnNas0M4XvX91Mer8ZCYagfUr2FB4ArMwgEEhEc6CnSjjDNqsZAcLFt
gjcpatlfy+/kxhyPEBuDguPDYReyzY1oHuPVu2hn3apxpLYVbAKNDPFFVTbe9Tgb
7gzrbwE4CU+p8FFzBiJRpMaqnKk6WdufO+fWiKS6Qx9TNF5UwexZTC/m9wPHjReZ
GPnJVWicK5yidmm3HU416DxTZf+dgi7t5zakD5NclO0FY73F2xKCnHgQ9W/QBznC
xZoWTukamRr4cvi+fpL76un/sdT/MZjLahmUfJBg0UaibR5LAOR93m3SbBIAnL10
tfnQS2HWeTIgeVZ4yewUcbC3EFu2h0dbXtNKxM7r+3FbQHZb4jUtdMXDNQgy0K+e
3AGwmzuRiROWgXX5j/Gr2HULfZvabArcJo5Dzt0t2BPe2xojYynBvNJo7ohpJnIC
5U2z7cWuIPQUa+yYa54YukhgQlTSoppUAA72kNE3DjtbZ9Mn+A4Bw9G+BPKTipu4
QEo/bYxmxNyTg0AJL0chBkxGt55fYG1qyXUmW8R/SPCxYFlSwbk5CgA/Tn7GKZMU
8YEniqi9/YecnuNYDzemVRneTeGM3HqtHDe+1nNTgLzdVQmjEI/DftzkJlz+MIQH
TEraVAxauQF/QsWORIKoDo2xXUSGkdi+3cz+NTeC0nZvcXn+vDLwz+uAibiJkmIg
nV68LQ3man+X5z/gbJuz2k+sOEvPGVOq2wzR3h5Edc1QqFqizTXa5OcsYeAnF6iN
0O3faHfJpVbshUv4cqjSX8JjKmd67QkS2BNStyARFgHDB2BfjySMhIsOm3HqCI7u
5f+W1mhTuDMe/AakOLElcPWKUmgtD5EZzyaAJd0B34diNCR1npRAiKgVuSwHXITQ
8QFLPkdfm3pLXdnB6ey98/7eTHl0fHCXKpnUDBIP8T8tBglnJNkfrNo6ooM+ozJU
gzZWZMlnwNTplnCr44Bz6Pgn1giAmfchsvtrM/9OI73cTCWAQfFbrXXX5egJJjd8
QhR+F7fbkiwogPZQk336nfdc59sry6lcYOQR2W2PRz2ErfmCpo7JR7A7tTfLu2yn
R/Zj5PVmGc4j5tm9ohyazppGzFaUge/pozsEAA2sUhMAHIiU9u38gMKgM5ngllFg
qxWqGg/jqrO4T5Z9VuwzK9SY8b5Wp3yZ9qU5QgyrTOYmhZdbCHIOHQuStxun5eP1
7/RXXi1FkUXpCM/lM3wLJaaI7M+KuIyJIbkUTTC3OiDO0v0H3Jngz0Dbnq/+uKl/
7Iymk1Ba8B2sZj+THt3UQRjNiPGHiyFH7WZ9m5an9cZLlwGQYm+oOu5ZyYXWBXOs
ekkUoOvtJFYsL3oRu/q7jPnXINDiARozGkP9xj2TOv63/G6Z3CKja/mYYWP4nJER
dwjHOS25XQSXm4E8hJvBlIWYStvmnNaRUY1Dx2STpiJ/nxAHsdVgaLFDP+xGWkIq
RN6fibH/l8alxZoLRzrJlzQZLGYukB30XKg5vqg4BSnGPsFzoWwp2uPRTu3shOTu
43waBj+IhJfvp+7c9SeCKEvxEDvxe5Lo1UMUWdUSpWy1fltjdVd/kU7MrvZcmFHE
RKWFfDRu9Qp5njRxFPEuhjhbgafc6olH+3QgqZYHM1rpGvjZRnct0HwhbcdxADmP
Wl/1anF45RKxiQ2lpFIfyAOgwDFH6VrAMlZPbVEjKyr2Ut5CjT2YCEsZo8X+A7SH
jPLaDHL+xh/CYr/DZd+hQX1PhMLmduccxPzCVeweH21Yu2BhE30yZ7gH7K40cT9S
TMsD2ohpQXm6LhNlPMsb9OfQFNqrwPm0a4mscvCVS2O56CvXfWw+4GPWdXCWKEz9
3sdnucpd6aKD/dHQuM7WywPMw08nfO79+gQ1qlzc8bE250WD7/gDeiwDlF1HXMkv
coJcI/ENA2HnXU2fdEqnE7G2aSOnf5qMEqJHNB97oAlCvH2eTep/RrrbTBUXlJPG
7VNxrHEStDxTYsNCR2b3gj+nxS3b8p6hCKhEK4u9e9CHLJr4KFJMfNQD/MSnbWVA
kmnt58yFpLjisxxibQTEUWEaJv9lX2lVodw3DVbnM9mnk/okOV/8iP8OH+NCFdMi
h5RWZbDBi82qDGuGS5fQXSX+ihlXNkgCfSZmajpqSIScphvrFLIwgf17bzFAI0sG
9X79zmjewbQcullMjBkNFMQwW3Cy5NfH5V8dmQVGrn59J+vdX86wN054F7lgJK1G
hSsQNmAso12cqkmhNurh4PZGVv1765b/6/p84HIB3IcynU8ZRO0Ipxfv7tXVNmzm
Rl7Wbwl5x2xGcdwbGEodWsuaU4M1iYcbMgPB4Gu//Y+OQsO81EzB+1i9NtU3UcwZ
NJd1VDX1WvWsRmGk8yHu3aVu50mCpHfZx5TubArEt2WhncIalPBtaZpf57IpLiFL
O4tT6IsP/+fNEuy1m69LAiq6lSIv1JEmtDsItEx0geD2psvLutyLHnPvsQ3AdcUw
WF76i3LCrzNat9h6Aj4vFYQK04Jjr3vWGUuuE+wvBpSyCDOAW7NDgKT35u7+ogg6
wsj436kyMGcPv31Pf6c6pSyB2oDCpVVMHuO6ES6/uSnnKkt3NMMB4Zh+92PKK7Uh
UOnh7tQ9Ge2QKdRdIqc5Y9Ciwj4Cm08ZJARSEiYU5p1JlfP9DSMkCounvjlzA8YX
XaAFquZ5CtPdPpwts1gFP57c0MzZeMM7usMYxBwNTRpI+hIh4wbSvpnqjA4HqH2f
MBKPM/EFnffdc1QOabNMAk0mX2Dbke0GmwsGjz7tp9eNvmXr/AjHdx5GMb4yyA3V
MyBgU2OVV64xXMtt6MurozHyFHJOfxrGEleZUdeKkK7xlnhHQa8XrD4c6KQib5Eq
cS/lGq2lpo93ail7E2XyhVPmmhz+ea8tOyarZyLVDrAX2wadioSziyVrEgEBiBlD
MmOHmFLCItAVbQ/rTdyUFdZmSU7zLuhi0l9ev+FXbmhB1N/SV3GRXnVjcU/ipv+y
l0ePWiyKyhLkAmgwT6++oLJ8KvnhviNFTl5JXy4B14i9P3/nl+DL4HP+qXESrdqK
2RC4Ip8bq/stq/KBqgpbnGuWZ3tGu/G/uEAXGaOPVEcCBsCOSnuFBMV+5dC1L5ak
pRXAQGPdN3RCHpfaMj0CUl8hG/OlAXCRT3U7B/nj5FQH5M1yRB3EB/PPgvjPdMc1
UjMZ+RaRDDMV8y4yRNa83x6l9MbA6WlMsfaRK0PkduhHol27feSouEVIrcVt8iVC
ahD+teb29tTVPeuLyMDMJ3FQlbaSNOTxvl556/hitIWVUX09+5B9A7l+7qmTHo7l
kPEv5JDRbeIJ7AwUY+xyvE+5xXreWGuosMQvOI29mOzRYcpmIMiNVDcgpSqzzqDU
6pxThG/vRIrrY/P9Yx17ZN+Q8TPIRojL+l8UtmEpUHqbHfaMAunzqJLPeOPlns5J
tVcNgXdIoyDXXTHINGLBLQ5WO4ho0KTf+I8sXgnEVwIUjUm6j1vLN2Ve41EEKegT
K3XKAfAUHFhgaU42iDrwNuYvToFK7bE/EyeUIxMpQhcCRwXh8A1KWePEy3QbL4Ul
V75BQ4/M/2Q+DTZ78c0wumh2bOU/Ys8pM5sYleCqBLjs0lj139rogeMQwCZwc3aP
T6xy9eyN4Qv4E0R/oZ1PbpegDOUFJz3YpgUubGKm26veh5PQL1I9v6K/qMpIlBhM
eDX+Tipbi9WzyPfmqGGLeBs7D38b5fi0Dcz9piz/Am8rlqsNO8mAACZYTAUXDcpz
dOEbjCd+QgQ+nbSSGPV79gKemv1tbvFmPTw5T4eb/LrSXMo4dVZKxoS8iHeUTA+p
bhbv2jcakcxkzcOMn8HVN26Rh2xY6u8E5Jg7XAcVSJNoVXKbgQvHfUKjx1Tn4CD9
OmBUE0GfBuLrEu+nuxAYCYQtC64caipYv7p9JdyPc1yaTRv5sOTfm5XoZnWjNQGF
99hiIakfd30lj4q6cyqpEY8vbwq/4FJ2PoQBtMC0uUhSfVejLjBNWG6r+jnsONpR
Txjz3BadB8dBo3Uehrs3UQTKjCk2u6Bh96N3yB9FeC42qPohvDPT/GXWFq0rmw2d
GZoBjmyObexk24eRKCWv5M5Jvk9hxGYdfFxJibhzGIck6FoLQ7J8p6STS8H0ni5K
1/STOFtoRbrU1MBHBAn5r/cBldJHeN0hhoBJQ4z4QDOCR1bCDTIIz5qqR41/D/un
wV+CCT1l4IOI3L6dQBT68Qv5nanHDwKTjs+mccqrpYvqz1bNCXBk5LtzJ3SLs4D2
3x80X9gv4/Pb49FS2JjpXC0YJf84al8UdGe68bl1aGkoXIBF1O+Y5kZHaLa4Kqu2
M5/FAeOyF0SmKb9jIswgUbGvCmDvBSTti7RQt3SbF7JB2aZ+LmmCoTTv+V/T2Vu3
rWXoSBwGOe9zi7lzasmnCYnnsS+epuOIEkFE1g23ajcxT4mBmncpoidi44SGdetU
pFznupHBFRxQiefsnloftV6RlJGfW12mQhyszDfvAcB4jNaXw1wHSnZNg6kxGy8p
qJW7VU8CQdrovtjrZ2BswtYkv03ni9Q1KegTZQI6Bnx1bnkwoYceU1TFrkYoTJ2G
6go6klm7/YpFRQhdL2ToIRjlVZ9QJ2i3vywfsi71lfJ41nFcAsrHSIxQFiExILY2
ajtbWfV4eaBMOd4FoP/0stg6Sfd/2yGjkv8j3bvjV/gmTv2c+gvynVXF4+NOZ14l
XGf1JCxBJ51MkmUiJpt4eJJG/QZBNnr0BkVaAS5YA2bC176NqhHom0bcCN1WXrwp
gLEAO0T7YQyCgZ797V8Z5ozAGynh8GIjGSB+J+ae5YDXVyHWU4qFF1A0S4pt9VfU
H5VxHgaV/477QhmjE1skbiFLtwnGBzCyVChl8LItvfRxcLi7r9Viv5AQE/pUlaf5
hv43Fr9FNbnkgJx4ccYgMkcNhZ+oXXAUGd2u/+09axbyN1//ny0jq9Gd/ixA3GXF
zeiv9npWHj8xdJ9WssOOCSNYxVoJtTbDn4XZrF/6izvRaG+EEd38gS36dNg37vWN
BPv2EM2bTtdKjrBgYP2OwhgccqB6wSfD6rRdx8vCG5y/jJZX66nw+L0YF/RtCOOF
ogh2lchTWA/n9bbhuM3gz1fiPBFV+dwr30sTLfDanUwliw1kaqTBTNmYTqImmQON
FkKsHKWYx7gZv+vHkkl5/GBcxs1F+vRYMm2DRxCdmx8XKBkq3rHWI4vUzgOt39HJ
50EAtkTrZpaL8CddECK60UrZ/SyM+yap2Y8D8bljdyBMmtIJZ7CrPE46//VD/1UL
sVL3Ve4NI+AgJZZIM6XCxlyYKJEwI6pIrY14NvBfAvLlkrtST2Jo6Qr09AaL0//S
3ICmYQSUx5DSSEgi36r2yrnF5bWshOmrU31O4haOyg5KkfuxfycBP60fXH+P19Uq
ltbKy0wNmHXZMDeV24+a/U1+NKTk8KG/wI2rrwMhG/929HZPJqcSg5mQFlQJMJ+W
dgp4FNRZlz/v8oz8Xe7jCyOigrDsWXUrob1qvIIXwOOzlYQJiblcICbRXxnYIC5F
0f/kNAVoXs1dCgNfq9LZpCqoTWwV8gN6ynV7q/Q/ONsSlnFMpThfsWrE2BTiWBms
WeYQivYAxmNu0z8Rp1jF11Rdj+HDOYx+huF8TluUMEXecn26Qt+FQC+5d74jbOHf
t8b542z1WTEK/4H16ndVtbn8Sma7er4qBDc5RNvYMB7vAHdovSaamv67s5/8QysG
iO0HAZsAf5XgWbv8T89ym9NThHy0UdfzKoUlcKTj67cPBG60kDj4xDxDEP1FAUEJ
UX6Wueq4dU5XnZvB9JFiAoUu/opyIDGL50MkNwkJsYCW2BFk4FwjxSSdB1TK4dgW
f3XXgFJ6tqLk6j101N2UhPtjvCt59ODxpLrLBmOHSy3s33BXg6uP75lxYoZZjWAu
zfyDUmZWg0W+T6tQFs3pniSNaRPJmsg8oTPqM0IdjNAgjyU9Si3lAbfTJGNW4APE
OKfvQDApiO5fyXS6ZtomnPEWzlglxG6exdMPl6E48u45zj6oTflZeVsFZ5UoFprE
OzvK8vyIfhKFtW9zS8CGMTXVpKlnxoiVYEnQPyvh1embvGYsfA2+0dG0SjcbnWrN
a14PTphkn9c+2hFOogWzoEzofpQS18YJCPwn6Un2V0N4cyw9U4PWe2QWPMdjG15r
a9zX9D1EX3EAsa2UsRXORBAMq7Phc4slYET1tCqDRvpjoED9EwUv2tn8cde+Lr4X
IpnBgwlU25dJT2Gc+p2XmtXWEVWSww7aLbslCzgOF+/NAgL5ezaN8zr66R4Nt2Ix
5L0SzFSYR85Vf2h8UgQPjcuvgTzaDn26AZWP6G1e2s0+YftU6jYjQx6awtZAldmG
uiEBMNk09K3Jv/8dz2RF6I2ldziXRn8nwuTsSlTCiyqCBpanJt8XyADFET7DZzpY
I7DidDod0Srpa718pYY+pkH5qcMTNEUMe1OP17+ybXzRRzm2epHMX0lCn3UneEh5
FFz1EKJtkWa11y3WjcYmXcILaVyfdOeAA0d68dNzXtyrzPLrsvCl8VaLIxu/LeQ9
n8bs8OrBzUEVJhLWDEmfJlDMRHmJhqLzHA0exYYruDrZSLj56hygFWQpyouw1Ja4
s020sZ5IA2xXNFkQEg9Zvt05A9PYAI0eVjoDR/ilhq0JhJOm71DKOhd+BfnwB1VX
dPEcOP01DqeACfCtluZrp6mUJMDPPY9XR3T1jJ63vR92UgnHqRdXd0+vcDiuX9Ms
8pn3i1KbDYSCs/R/KYoY1ebLPyla1eqh8UWZLovgcGMAEdQOEwy1oGGM5FXq0pGw
JAkPxH7RHbC+dKl9fXzQRLslQm86/HdhDYi/rWO1IKq25uA6u+EMx0Ccf6oGkPjb
7mwRL/eMrVKEqWlxi704wZElwFUdTF9sgGaUSTZRG3qtC0ELCA3e6xsc+uGEuKLS
5+IsiWK3FAlLoW+vpsTDyH2d1Cehek/uAiVVFaN+mXCQTLu9f8QkPFwUpyWIcyqm
YjOSWl65xYubKrWnE0xtsxe/cq61na12amReihdyIgkxoYjUdjbSliDG4SsQKGJR
0XaThA7028trXUE19Xv6IDv6CbfOtjfIx9ljEwhBxwTwa6p3VOWEqxRDs3ucr2Dr
XpcN+ghpwqsYGZCwJXHthWaoNN5djvdNsrd/ldiuK9LgBdU5Kxbmt5FOdV72b9sq
/dZtPHtgngfR1f04JtBGdxknsNijQLBCM6yAXdggVwK5w9lueFNdVp0/3H162D2o
WvXmE5oEJLa5U6xj96zcV2kLU5X60kkPO4P24xFWuTLUSicWXwNIVBVWzlvWxbeY
wx+Fsw4H+s0jDQuKRQW87DAOccJNfxJfDJmpjk3+vTOW6PcGAd5NK3aXhlSOpPjF
MeKaJ9hkMRd3Z1q39u13QB/Pj6ljbqEEmZQ+TDyMYyOM3hWCSG02b7hNscv2ylFU
Rp/VB4oWTXi/7O2fSbgys5VDEOcYWop1mI+vljSy2KCkGjy2A6DozWuvyIT+Kupp
MWWM42Lr74AKCT9PBNwgyLrXxOeSQW6K5hF2xQTNGbPYFf6C65iFMHOVNvdvR+sA
RFC6CUD88BP3MNN5/q/4Khvj3IEX5VCjtBKqp6MjwhdQ8aE1+QVM6Ke2Lsamlc6X
tAVbjd+Pc+vhONjTDkntktds+eHviOzRtfqTmTrhZqQ72W0b+xNabe+j25egaVb1
9G/VL9PyCM4bm98blelhXajvXsYDYAhZCLL7T6vTzjoGuZWoIIjnOAzWozw6L6DV
gR3owfzlN7vQYT5H8evJa+27HAsUFacP7ra/cCsS0taiFYsLDApihOe6NwiqlFft
BYvxdARk/TfWivHGrT0ijwJEga+/APeQvP64SPfXrRmX7V/XHDltWaL0LvLDZvK9
fgbPq594xJ1exT+QwHFgq7bxuCOENBnW1GM/bnJgvQIqRSDJMPtxHfetKFGfUgrF
v4N0wF/EHSwEhH9ObroqRY1SfpnXWoa32sCzlI5j+hpC4h167ddO2sf9loDk56h4
B/8R4077hepfptXZOdGYr7y+UgmJ5KbMJgYH5cGskEhnVSCyGEz3mo9OcgAnif8s
hpVq8H9zFJknILOJXE5ldJlgpNJ6glytoOZgGPgXYaDLZ+zU2DFQREiC9nr0l3Hu
M86H9Ss8hX+G0oWVXv5f1SDzYwEkpQYtsMLwDt+mSFqRcu32AlmRg/uq/Xes+zSb
dJQQ7NVq7812QoAaVl2xVPYHTiDRDNZmRpJpMfBDYmWDPFXux+zf8Prierf+R8yO
lPA+ZQWn+tEg+kiMhD87lfuYVlhBwH3VCBCD+VKebcmFy58cEQkURxVBRPsBN1Vj
gdwidBcJY3GALWTESHvgczypy8NvT6jhjVVJpzPu/r9gpLx2ShSWCcHMmcZp4jVw
hfS/n+y2exzJzMj4x/mVJ31NSWUDymYdnW2V6dnMW1apHLsIll09do8cZFfwDGBn
gBRdYA1MV9XdPQyihE89BSbTJxo1sVFTmcdh9Dn2WsAVLrwR4fJVT/zRrYAIfqxe
pH6BFPOWuqQV/RNkzk14bhoVeQrVB0zOTsCHU5sVctVYewcwpSGTpDFmnLyA7Bse
dUDfJrbwmDbyZhNX81oJ01RCDbpwHkRgKSTP5CG6YS3LQR0uHfNFoBjn8KsQzs7g
sRVdNiljche1Mb/WxnBkXQS0UXA6+imK9rGW99Opnm1LOPJ7Xm+mrAFAFVpC5yLB
0NdsKFpPj047T1Z21WaTFw2fUlzu4rq6Miw9HnKyet6zx5WDvXi/J+9W+92BEcpu
sIitRHliuy2Z90b3HPeopl4di91zjHGqdyNhKF+N2cyrHTk/eK1q6/GWjHJ1Z3Ag
Xl16WLQ1CLEFlUvXrtcETaoDt3BcKni5UhgawNdw85M/2cukxJ2AtUXu2JVaf0hD
VVANcgeVkfVbQmzrOIlChPCbuKX2irz88s+90cWtowXh0aLTl3xBrQleCiMEpaUI
J5SkXNa4Bk6i8y++0YF5z+zquC4mKhuPoFTQAQOXxtPmzPb9Bk/TTnndY8tLrbPh
DLe7M559KwYuKWi55YaBdm9IxjO6S90FvQhk6Z9qweHiyEu7Fyv1QsStRMai0R6S
OOcRl6W0uVB3Xia393CRPbJeV5mB7LcdPDCqGp0XQW3QP0OE283ZTpSaVdSgUwws
trk+flJNNMsoZuU9eJquZcgNt46I8X0/0+ULZgY8kLaC10vgWMQQoz5Ld6Mg8YfJ
w8251lsf9dDA0rAsalKwM3HiFTUW0lxFLKxUdCdO6XHisSB5+1JxZSBMsi8eZWKS
UJ7GApSq53zFGZsjL48qbOeXkLU2o9j1J4bu7Hw+UiR0Y5VF+45FYvPSAqInmjex
xbjCRm2VZRnQfPz2sLYmkVPolxZhge835oe9XhYRQPyW+8aDYAHa049/8kZ3rMXK
BWJRIrXsyoiDLChSx6S/ZK9AqRAfl/qSgzvjEvlaLYgLVTmmjFYk4A2KjU46jUQj
qGkCY8VHGqY8VCRU9phRA0HGJr45VzMU7JmE3qqh/VJzbHPL5FHMu3cJ2Jsozy0E
L1ap0Ix0lDzVXcA0/qZzHgxuVf9U+uuUSUjluj/pmPTl8+bZ2qmgvalEZ/yzIw8M
Wic71IviPzLBvGalwU6uPzSm+qeAm35XbPLUFOq5TvSRCNxtLcMJq82ejlucRxKX
IoqA0kufte9oCEzzCXlf1cADjx3HW5zvCY1cRqYu8LD6Po26OuhbipnJCt4uGoDX
IwLJS5aWjeGD/pI1Gb4brFjWITcmQnuHbIZTdcpQ9SpOlf0RiIRpMHppmGAnkYdk
t7c8PiVxjqpJJnuHNCt+VeBnVs74kP5JL0AWmNQ/Z9Kb+3Egl1hH3NTXb9FMvQsL
oCiHfaN1fNszilKWkKzBA0S1SfJCDmuw8+tJ1UP3mJrPVcqfeZisMCoDfdgGZs+F
uRWdOM7RU+1QNOLIeoiMSMbNedmCpUdCMhZC9RYTy/peGOEHz7Ktth3145GnErIs
95lq/pIZgZaVwXbpzhI4WfdtyHblp8TQSt2b7aGBYqvpGlyA/mbYmluEP00233O+
UbwlnI6Jk5mqztuKkUkmKQJ48K8GI0tarLU/F56+9UTPnX8UF4aiPH6biLa5Iz8b
fWVH5SUV8vtAJNZx7+5orUMmpY1UNS3VPCD9RXZzEdLO1otAU6ON0J1buKuJFzgo
H+6X8321udq91AH895UMEE4+1vSvAbI5EskRqGc2wI5yA68F/dZ1lW/F2YO/8UMQ
JG2v6EuS1f7JpX/saL9XLubUYigsBqjzBpOw0rR3VAwscGI2jNx7xQQMRk/ulf0s
aLA/Tcq2yhYRJ3PyTZ+tD/xWlFSkOqlZb8yuTd0464K/LhDlr1L4rLMDi/1fS+WM
V7RqP1ZHxUHRslDsak+rKQjOhhlazTjFASMLFT4Ubh081qgMNcltuBk79OCmixat
ToLf1peBR7OPTtk74G4ngFjS0N+eQPBJZJtDtBWnbRxMf6bCEX6upqqNqqIuN+Q3
zxXWsEhXR70SiWMVtXKP1lMezsgrZFYu1SPpvIoY0Hx+yEJg2gQI1bGmt/p/xFml
jWAlsAyvPATYF+Gf+AuipD+AUaDddp+hw0+H5GJtlPMV6QgTmvo6zi0jwBhkV3/v
Zw8jfHPcfLPS60LnDzEjsoALjnU1m2Fjy4v+mgwpPemnQK4MdriZGIURcBEGBKwj
G/W51JiF+t6PUCp20q/5CYG6SG8YYx+E6xIeNpNjw6pOHiLPwgH0mtv75mbwBAsh
DB/sIc5ZNxmSyHv9yTJ9wXW8B9Rh+Ws8Wiqe/hsKU3nZx1N8HSUfep8BzErD0qB8
HyMrH1F1GDpJ+H9Dxgze6dRwAfv1RAx2iIi/DEGfFKvTku6EBKDspYYZ4rz+CblO
IwTG3gzzNn0jVi+OkSc7XSn9sblBT93AbjLYl9kxZQHOK1uzRBmLA5rEwy3CQxBK
2fvhuo10uHq+wwuOe2mEQXp1r7/Fjuve+fiRYfhFZGpGIJtrMb+1xds89dSGAnpm
2wsdyqOA25t65MPXdwQr//BUp21SR+rEs0dvrqFKBP+Hl0Gpfdd7IPEjIccjSNcV
bz0JI3xU2x3XYemSRDZAQwsHzjlYHxx1XjGbGBtgKy8Hmra/JlEL3/WkjnwGRqPv
LH16xHK7IQzkXcdarDNAa3hyCL+XIgKzEeeqcMYYQk+7PFi5WPvztbJRa9lB0H6X
WHv/RxqZvgCCHl+6+z2H/Cn1j5AI4fdVRA48y20d0AqEng9m4waCXSWWQzDsZuv9
x273SrP7sXvxmechieNHBW87nGFCOG0wu8VWo/4djACrybVp+OH88909Uxs+C0o/
ZUXKF4LR4fm1O7GdJVz7RTOWwt6P2kC6wtDi7cZFZklJzvrFKbdDwPcj5sVvSWi1
hf5dVXLDsW4NIYCP+FxmLWJVv2z2GtsXNQtIRFnEETKINXXy6tKJYonzQZ/PAZKj
YLHdHFe3iZ9tSXrM/1CckWA2P676+71mv8ZUwYDswAK9fGTgQ1SgnWHzdFERKHx4
AmiA1hVewJxj6Lk3u1P6+E9MpcyfI8v1ie9/4FLDgiwPFL9pD/UwhLBAJeIwI38L
sTXKAhUXduBqF4ixPVFogsmqghAI8sPG2oxDZWQpgfUSrPBuYAy1d6OqOMYrCpi7
Y/XHJF7w3jCzR4+P+IGomkQhFJqLqgK/9QvwwMD0UcaIjNNu6qY+KUxQk/JcqwMi
wDRCetRmdJ+r1YKM64PjxPgYs+aBB8Y11xf43f1HhISkYeGhK/CpnUwvCtsuHLw+
F/j2ABZRleWLqUKj4m7ddN7lNl9K0g3CD2Z4T0pdXg9zbxCk+PXPClQTnejpHC8z
eCS9CWwC/1maKVP/JJqVTZ1iqnsJTvbuggdYCn0XhqB/cRV6OL0SY+223+KEdwwv
tf/MrK4XLlwZUvokVBZAsldyXoqCFm3gRuIavcXTE6JMM0HtJVjM4TrPlZGrqHlp
ilpFRjeFP/T+zRXGJfFbCiHwZItJmnqOazPc1MSA4Ckn5ebphUoJr0pkyWaVUVN+
MVcJ5SI8bKNhn3OZrwaLpt5pNa5rB1Rq0ke5EUN1GbS/GfHBeRkGNFeAcJpTxUxY
NmOTJSqKaC5M7ao+b60B2u1BMkv3Rdu0XIPmmOS4Z3WOUxcai30JqGQoowQzn6qG
jvnUCp2m11hxligYskfpakcpteeR7P5cOUj21Cl4yfJ85oCqxpzeCpkir/LGS47U
4u9HxIjRVWUrrRoHAQiiW5kWvWxCidpDfcO759h/JdMfViSPvjfVHMJ0JOH9Lr4a
xEjviT27aupP+TownV+z1SmcYnhtV9TLu6MZfAZ+rhghKR+1vSAF+NQJItiuAu4Q
VB+uNg6a2J9sV0CvlYo8LJ+W7RtCHV75x1AphCsY0KDkc9CI7h0U4PqCMmw0xUpI
6cjYleaPe8wVfKb3XjFs7iXpt3oM9PJtb9P12k24ULxgs9AqqdTF+EHIwYaJYc0S
1EwXYYYBkTUg/DpHhkghuWg2hcgzDdcZf8b0YAiWt4T+dDoQyN6KL07Y75zCeakA
08w+Qj3KOoB5BTBN9xg/tAwTzi1tQel1X40GPaFkT+u5YAlRdd9VdcL6nzT8VzHQ
6G2+Sz75yrq3ytHXL/8gPig7upXcSW/vkn8BAd4F+uLVuSUe4pDb956vpXiwxGqo
1epV0r38dIGzA3HWKTmo1YWPr9nPrGN1AHn/7YIBuclGBGAC+MLSOt+gQ6cNtRgl
JaYm1oBZEJ9MRLjSXFyzcVxQ5Jy7LnEj+pedkgXBW1PvbPF0uUJmfL7a7qXuxSc1
/qCePvAEdNLaCNcsHmynJKSp4A+dsLrGMvXtXfGmaLVncz8vD6tvewTeVN3Igwjj
AsS71f3SKMjTjOJJFMTGsNNpunIoRgfkeXLvNOjhJWkSWhgN4YZ8DwBQiFvjtUbO
BNq8J2wQhvcVBw1I//oGnnll1TWEVp0qzfAt4JnRiCcgg3Sjt0ZgeqEm4hsaQyp+
/jEWi4xfRa6IHSrah/aHSjiiargMIBZSQVKUZRGVvLYYA9nr5tqrAx4sjINLslq/
X5GGttGG80flXRzkgmHASwh3B+O4iI7nWBl4D3QM4QSC4PapLApJ2LYQrSfCOumU
VlAZdrqS+FgcXQBZ310Nl797f46xRmgarodCorVo3yfBUbbsRr40bTqBIhk7oLWg
xkK4V8pQu8FFThWjL5VE++vp6uF7q0IOAyxv9DCLZByof/uC0rgp5H/eIg12+4Wt
uGPzvBMA2mDx99JgjhJv7soVqoYUWks4l+R4JgU3Cxr64zQXXqXZN2UHgDu5mGqB
7qqhJhKaHWVBeMrxZ1hm9xGphFTznpnRcowPYeyEntMzNkAKeCENtJh/9RzLhCma
V2MZ3kwQkgEa8Jq+nJbBlaOPUFd33Svq3CcSKrPKLgePh4699tPI04P9HnoHmpVV
6O0aanuuBl24+B2DHdzX5eYuRJC1+b9+9KM8JyUA/8NgoE//7aeBG6nYRf9JDvNq
lkNotGriLgezGhoo+8mhcminIfcq8pu+5NgqxVROw1kSMjVgRN4A0Gy5Ylr999Gy
500YaIhjayqn9nvpUIT1ToBBY5FlGa4MFJDvP08MzXTrzesqO17K0dFS7hQGAIXc
eR7OyyNZnABY/yRCc4MdKNvd/loYyjBmVAR0qCvJnk7zWIClaATcDHTl4xmi8zsl
YhJwMNZk5ai4X957VBuc8wANAE5i7zKwDlkbHqZkJZv/yoVeqyZwNHCpm7yJMs7J
mP04W/7djkJ95HGLsvdwGUrZq1MFldbsTQPPSoDpw36whVTFk0kAExWKOehYhIOf
9cOXIY+3Rek/7kSVVzFhL/gr1DWbGHHHv6KaGbO7uuly8i73ih5V/9+IjkkdkkZx
83OFbLemPs2J8gpiglz3DaNpwRFqIcUAgFMPZFDOhYVrLv1LZLFGlaaHlHiGt1KC
gfUZsjsyGZocuY9ikBH3yRpA3IeBBrAJmRAig0Cn0tu1zdGdDVaLhdPxe7qpltDF
1qKXsarThuBBtnm+TiHrDgZ7TExYXz/q3YzlBfO7J2RBxyiX/s5vTjm0/j1gCn8u
OCxT9srbol3xISRuJ4EG5Y6pybKgg79TbEyjz+LQ9Sj9qk1eMjMjr2P2Mm9w/+L7
fgma6Hftqwf0931pVhHfRCbpeT/jx0F4/rrX+IyCTF1uK8SevJ8ZU87mA4KL17Vr
wVAF8Rk1m9O6JPuImkTyUgnAaRafpxZWJS2UDAkyEVjY4A0TfAHjm3q0QuEAgx3A
mIyvOs/IfgnZO+PKgr0AclrR8CwAvFIP/fvqD1tWZtXh3QRvpea21avRwpe0/WiH
2tuCEacK//RMFUcqrJfY4TjJ2qXGzhSFvMaDYC5lzqIHCmjOL+tjBAKlBA4YzlcV
qlMJ4Z9VCwWkFDghX2QFF7UZmgR7nkiYdZR0jbAUwB62jLiTDSFvrOW2nMIrGWCP
r4LCyBs1IcQIhwbrPgXsmHUsc927Jkiy9zIGx5QJWxAnZyMlShtdVLFg1eoLcgku
jcVbeB/FBG02hXEWvsdypjkfczZLQDUAJzumowL9IC5DvkR202wFC0+SKWOZLBm1
WzbvrvbMd/21OawFsoU42K9vqVGaqhBwTapulUY5qCqLhsmBL0nULaQwohRqEpUa
urfSDSQrzt/V0Rn1NqrKA0QJbUF6oNgjpR7kiXcHoVsbeKizH6wjODSiO6S6cumk
s2ZIWJpOSerlABUXS1qmPM4fDn23UVgb//9gcEuylksCeszzBPTS1HPmvd7J8QHs
00mxngBo1M1RmsIrJImR5JNLSYFusbjZvGgQbYOJza9B+c9dPy2SuUxUSAzv/CHP
ROBPEVUHYleqKW1jvM9lqJ2go0Ge3ZrGL/vIuhmeZ3V0vCx1vGa5QFmNy5HqjNnG
4l2th046qJPeUVuQWe1NdLu4TfaWSW1GrX9xmAo2EVUtad0e7I+U/N4iUmcQUVit
gvxP74stiPW4yQuzaZhtv+b8nkuqYuTEZ+Vyi6oViAwbyBC49JQqxMLFvdHrWN0v
8Y+mFFXz+JJ57fj+qANkc949Jl4ykrFDityJ70R7GkL8SMmAvkpzNGmvnnExYcRW
bqJSmGvBCL/KmSscCDuT+ETLpik6WfK0YaxgmW/9vJIcOV3faU9PEWf925UaPRxi
yOwTdZLcajk6Z8OliCpGuF3uZ+55pGpZwYjYFl+f27o8OiH+fR8OFuAzAPG6dlUR
M+PpspcwUTgS1HUx1DbWhWxrzWi+qHCijKGwSjtJkQ/+Jo3zafWffkpVNssSoUv4
KZVL/9Afluiw8jwiRtenDqJ6kzfrYyc4La9mG7iruDQW18C7N66oBkaFaxKx6N59
KkAtxUSrU2g5c35vFgGGJc8GWmGkfIJ/ERDI+v5ovhRcdxx3hvx3I4fEqXKnSCsb
NHQgp4uwsnPaPiE2nNofyNIEgmmfXxsYMvba+D4ZabfQ5yOP9CXYnPKsGIol+xdG
WCtggWWsh3z/GVt+W7CYdwxXete93gO0CrO7IpWVNqJ9oMAQGR0B/9Q7yvRKBQqW
gcpHCYdQQ3LA5m3R889UMJFTSy/xO2bglcrnamo4vDBE8RIJos64908WEnKwRL7F
VoARtNFPBcyIcW3UP4qI1bqCOFq6mlNG5wDKF1J86PUCZkBjbUt2Utk/2HOJCqnB
bBe/zTlW59wQu51tfbTEFC0ZAodIs/CQ/jwDPbL4DAVmRR6rlg9hnCG0xSjsnJTK
tBU8uCdYvf1p+cyPtpAQA+fHatcoQR6Ut5EOqoyftdxflty5fk7oU2B7rf0VotI9
7i0Ef65di/3IDYfy0w61wGwHnGKDNgy5Aep3O2rzs4sddbevjDbzMcd3g/diuPUl
C+uvNTZ3gsYUwDaMl/8v5hKccwwEICGDNEnurwnrlJ2Ay2uglrvWbEyyfZG91HhY
OU/XIh3BYW+mhJeeF9DAsu2A1hibJBDLxa+8pP9pVJSyGrQSSP06RkkRE6UZYx0S
4VgNMquoqF36ThO4j/FJcbFiMarXCuo0EdPkdQwkuuQyfE6MEcrGRDJGHOToqzAH
Is8fYQeDYh/KDfJvUcWPWyqU24JOjrAZp6uJonOzG7q/ukKfFAQsjwJUeCB01goz
16sVl89hK0CTdl3bRmxlM+t44/92RBreS6Y+gO3JHFPio2g66gxx5fHfC3KlJ5MY
y89w4aMJMq2SjX/jQWK0jL6mt//bhZQ9Bh9kJgXenuee9nioPW8eEcLE7RxM8jzs
v9iY/oakPAY40FVX5ceulhnHCp1L6oiObRVvD23FBrjlRyWySdSBOUygyQi5uM2k
Xtofm+t8I57CzgP2KIB7yHX0E0CV5SZn5sdeAHml6Uh0VjfuWl+7ZX/vRZIef33S
nyHOO5Xpw4d9GfmHtV9SqomK9PBJhY0ZDj0KAXz09qZ7j/uDuAeLznKcFbe6Us1z
V/ZgZHZbNJOWNk16OSt1VF1vHfcVYPk6ilthsmDlLi9KMRFfQocQKdJ7qO+nDmKZ
H180iv37KAbnvN7K/mW5eijJ8DEvL4JcsfUGGfEL+9r/nCijCzWEBrgn4hUpIQyq
0dvAw331VSJcp6u3SjOv6gWHiVWTazEVnXTxBrTkqULBWF2JZZww7HHL4CYAHgKn
wooqzrxrhNKPqnT6w9rIuyg1wtNGmDEK9QzI7vDwZM4j/wDJ5wC8OgLSd1spa/fh
ZGipOfY3n88UGcsoevnUU7K3Ng68jA9qCBlWsG8d/HY3iKd4YlV3bgupYRZ3DwxM
FJZ2MPr+tr6NJp97RxmTn3nI0gPYFBHXsIZgBW5R1ajl1u2aQ6uXT3CRPMT+jVMO
gALUpCYOJmOH7ScfnbioR3rqc8guCoCtdjbsvv8Xb6G4knR5ognB/9gnD1xXwiWD
veChk82qI5Ld59UB9fkZp1p+Ji6QnRfSl9GJ22rEfDD5IOUJ+f0oOcilIh+Dxl7x
ESfoFs/2lbRYZxeYegTYVYAh0D1u9roF1mlrB30Ik7PNtuibrSvbP3blh0aolfUH
CxQiEyhCHvf9LWb2vA1kdykZMXkpNfVPBpR2i8gqpnaJXzDw4b/H1hc1R526xzDj
+mWQu5+3+FLKmprtPytS+Y/m7Lqo2G5gex1fdc9SPGN/yfgWOJUL2N/mezKYg+6R
ZD7SlkYfaK2InRWayc90GB6yfcOzg+jy/tNTCO3BxqGOte5/udu5sb8h8l+ln2uo
GbOwX99jDz8kKG40aJhI6jX1U8O1M07VgNdw3ecEIJqBM7/p+hGGyjSunvEh3zkE
KGj2P+9sFbhUQTuGVlK6MCKQlPuMqZp2VnpNJRpnYwN5prilXDnx9L91egEvoZRN
bgTHYWPFpHlHRz+yoNZJW0wXiK/BJpVHkwh/8HxhKH/WAdc+hyvPCTZyv3USxj/h
87Q72pd3/rnHl5szIR2roBEdJEg4Hhtn0BhB2+2G9/sdK2mf3HhCKdJNzfBYqHeC
bE60VmXtX+8eQntuK0/7mVI8y6689bq/kTDtxY3B8OdgMP8kSi69PS+T7sKu0lnV
zHnsWm5TTrw+E2ykNcPQDOE+UeftV00VmV2oAlFdzQ+aXktlL/XOXdDFoRVrxnGQ
DvNh8255y0MYONGLNvU9q8vxKbi5GxBn42maoyeXhXX+mXHQawa5422doe2236o9
DWkoCJX49CCv8NLEj0nj5fDUKqlP2u1CBap5tlqZ10w6B93YfaFBNc+TEsXlCsXZ
xycS7Z4pSuAT1OIYGk3gCGkyYfTUTI6aIucrtdoXNW3j5s6j1/7xc3owDQTyOplQ
S1l+bUZFpUaeam7dvAspwtAYA1Te1v4caXvIu8rl6LSQPHFj0Ss9Dlc12g1gF741
mclclnXskLbZwc2R+Tu86v5/n4ZcZ/9iUUtz32GiVEvkCGSY5Uw6A6cwNHqhuAzP
tfVjVuGcRhmkybEEJRhRUMktvdwjeqvvIk06w5c6TVS7yBFrp1b3+ap4TcRemXw9
GUAxZO6dwbxG6D50eEAUhddyEeC3x+kKZihZh2R6SmV0k9D03z/xObY8ON2+rQCW
2YmtmVXEkrqRq/T2lDBA3UDBFoxpTKV/eIMrkMubaUHTbJpjdNIE6syX2tmIegyu
jXsKcb54fF7YH74uEzKROL1XvC3TVdMnOcnB2ZAmOvD1nHS1NXIE4JNwzQbSYpPX
ILKTApXzDJqyMDJPNJ3FHM+GP4ptLridbL/3+QIWhlZgN6sPpTUYJEZzJS5dwJfU
ZuK/1B2VmOa2ghTQOKa30eakmsPZDoMDXkk7dtD3UYnaKWS4YqwKFxRxC7K0hdzp
B47NnQ/vQBFV0Ay0nZQ1haE8FOAAp+Cvc9adK4e3WamoZ2VVlyOCZ3MnTjspagJm
87EKyTwFibuI/rEJH0cn5suA0U6zDqO10U/Gudmnh08Vfau0CoxXFIe9KYOxdHKt
d0PhP1QYVuM6xh077RkUqqVP+Y3ioCpFX8slhmA0a+MhL26TO3GxFyG5b72LAMrn
d5fcdr7lPo8OAkOYg9ZhGgN88pFYtCbBcAOy79VwhZVocfaef52osAPVyLTz5wiF
zO6AbQSh01jUCP5oDhJhweA7yHQhd7lIff0YHO/zCefoFO7Zg56IcPR9sfKhrF74
5iqbNMqmqTWajaCu0Z/E1t6gD3qzDpNfI54EPGjJD4ovIdaLx7VXjsm4E7YMmlmm
8JcTEQZlFu8/CAg52TFTgEpyP3XyB3P+pts/56mXX4250v7H+u2Pvcm+UzT3PyAH
eishx570eJ6oZoQyYma/x/pl8DEHxH6g+5D5ESqBi5WjKaTVGzXCleNMb8y6b8Ie
98yF858TJpOeBilFTfvnTDJ69KzO7THsmvpMjZSygeJ5X4Vf9Cdsm5tGsiBraBQI
cDAfKvL5FWedPSRIrX9b5P9bMaE5reDZuJIp/hB9IabF61lZMB0xj96dvAULNOuu
CQOTDBIan0HKuaj+gxNkcET83iQMxIih7alj0GyG6K4089CZ7y/1OY1oSlOS5xGo
MB+La70AE42D+Nfd3gN3M32MFX5XKjTSgofChksspJ8a2snikB8ysfKxZVOJy6DX
EeNWuQw497abvQnHWImMqDtN1xePkI/DHwUDUHVUHzWBwTf/l9avxRZc5CaJdTuL
HIGsY+ivrCe0csmWEvw272/49nlS8oagYo7vvp7fKaOSaJOTKA4Ehd8C40zof5G/
OoXHbzXw7NgiEzawnAyM6B7isGZdHql9oPeJGPXckxPXCmiJ2C9ldfRD6hrk0h06
c/AIiCJeNWrtDA7YcxethB2AiKFYjye+yJRgEteIHRei84dFkmmS/m3Qoxrif44l
hnuOUrxd3SrYvf1cua56vHjnStim1rE0c/zLPNq0DDoVay9Q/sRST/wKCp2jiGJ5
14NRYoICPSFUIIQXF4vE4jXC4hL2sxP+RoErfm4qIfJHl8FhgZWbGMVXvatZV66L
Hb2vh5XZyJFTNJDxS5VQY8hMpFC2+oIiS/eXyiXEB0xExQnhGhXDtXdH+lherHxV
lOeG2xlx5JZ5KVZbwoR5xpfxy+C+r+WY1S+6v8DgTdswMMhis8ufrIn+S49iPS8u
SWh3/U1kWLUo14O0gUYtF1qIRgjK2h46N7Lh7Mo5HsRtF9cdfPIZE1/YtzHfjeKm
8HTG5x5eQAkmBwQCc99h8g3TOuQy3MuP11trOmcy5OqhTCrTZG69OdL30oIWxIfj
g1kpyIO/Cgez03leizN4U9xx49ovD1tl0nTqUmHYLWdO6Jl0vug36wK2W+cpIhXV
TWuzln/C57EQDH4jPgubdzDaEm0Fxy4tz8qVKZTxdPCf+5QLiEIWGG1nnyDqVt1Y
p1tg3ExeoV7aVfOLQ8Cu61NBiIBTHsgkz5iRmoLJX1gF66e1OfjnCgFjQ+k6TeEp
NvQtaH+VBNarbGMI+D2AWFL2/KILQ9OUBKGKwSxDBWgmIZgMqa3k+o3ocJSYdLl4
dr1UGwiSbMhkzVnGBnozeHbC6EXfT62mJbuD9YohHh/AZhYFdakIdMVXddvKJDR4
y2GjWwPWR1BxR5PIiwtSK8DgwfpmXGqNDOlkPSOo68ECKD4VpJuz/QeUdvFjnuPG
2I19lgUTSZHZQ/VyIn/tGDhsrqoFR+zla6TQ6BwSgkHA7TK0ZCLTplG72yDs27ni
o764io6+YA8+vOtDkB2HDVJE2UwpCMkF9w9vLjXEK/orfT627gV8JA2PuyBF0wMq
tRcGGzxIOnNe7kFB3Yilp+V1rkzy7bb3u5TrswGGnMTrmbz9MqLk57CrF2oDatM8
t9RspLAk3xLsDq7jSOwzfYpYUSX+y+DH5EIiTUyhm1PUUkWVFMxSSDC2a5rLe6wJ
b/c4AIfspKL33WtzJFyvFfEgkOpOfs6MVgv0X23Jvcp2M/JhDbvcCMw3dBzNI+FH
nEbH/1TsZrGfYPULrsyH3Mo1Y6saIl4EXJW10wQYk6Cjt21ehw9wrI/SaV55nft7
VzGnI5HygBpmvPbAGKPpp7ihWpW+wV6/Z86DZBVmOoOZBf8b6GDJDPNZhkT4xCvu
h92Ia617tvIToQ9Wkp7kKt+0bsPOqm/jFgcJUnMcdSW9owGi+rATr2rcfOYLmGe0
w+JY6/8+Gf8TkwAJoHKQyzvn1QBOn1J3p4EYZyCOfSlhjxdWXMG9LQn1egjYJmJ3
lOV+UH13r3OCSfwWU5gG7kgGFaZwCjclCIqIWYj1c0TJiXq1oocjGgItp3pWfxfp
oXBmpjvC+VbshbilUjjqf0o5QXrrpxG5jhcQ5ojQef/XK0oE8Yy1iUc8pWLK7urn
OPtD/SpPN0jN7wbFKkCkcTVGZ8JgvTPz1MPe8y3Qr4jZHzD45ydLpOwLHwq50nAJ
6P//RdAOiAiDJFv9xDED29WwpqCkmt96J4Eo+L22ogDgUfcy1FNyf3kf4FRCLxb8
7beU67uqn3jtZCdVd7P5fLc9FHift6Soe/hyw82tns4Rg/6zbXtcghiWsX5Jeh73
AUB9QUkJSeN4+4Y+oXyhLPKRI/BipIQcPNCN8W3yea/Wk/KGm9cdkWZiZ24GT0wF
fa7RaWVLoDLaNVh8KNaj53vT+prlu8uFKzCGbYVVtAaHQpqlJ+6Vw/SR48Ln3Bbf
KMLQJ+cYkyGYiO1p4RVLw4r+Dp9UWpIr+f5bs2bmfErdwMDMWEr0tQb+gAYT+r6M
ilkH4QnrPbreqLUQ9hY/m16ZRUY9ErcqzXT8Sxm2V11j36xpgjuM/eiVu5Olpn4P
KvgkFoJ0mAq++HzjdV0N/hRaJ8HdMro+hQFcjwIRB3fH8JibsYJRlYuXa/AEMBFD
yWYYJT1WJK2NdZkbvPCJVfnt+vkl1mASLH2903CtgnDSBvrzorTtPHpSZ6DEbf56
7lfP2VRZjMN2Y1d4AanKNVx7ymiH/XtpwhZFPypGG6axHY6ZxXZyTGKVou4X02MY
Jpp9OUXyRQqcUEcbJQgJW2Z3lNzD194Fuseey73BPPneXKJCagaVfMgNP5Tf7KSy
b69X1aAWMLI+p7yuSmS3H/DFpHWWfT9Ndhx1Ue78YmSonZepMRiEUujskSIDea5B
2WqlohpnrBybEOnk+yM+POoQ/S/VSFcjv+cARbETraelLyGg0gYfxUD+Qspr9kxH
UlOlx7mPpjw4h1fFxEw+ElsY6+IPxLDE9Z3vQJJUeZSnJunZ9jebWchEVWyAl/9n
YSN8KOdNTp6cC/pfMDd1m6h6/0ixiKngWjiEKJK4Pcm5BmmNyvLFwGdGP+125mmR
CVo7fRNuB+ASMw5pXsaydSaUbxasEx3TG2NW65QYnMLD6SY40xTWZhiJ3s0BLQqe
Vgi3n5lkHOhAp+XE5pMlr4MeTd7VDIgRp01zHjvPsKnJon9x4rBSFvppQAK/zHVY
+tJQLOcCbUmh0EajKoEI6SeuxaqAoWUdmy4l5AiuNHrDDAnZVriaLNcKuZG0LORn
X9Ay7DGOUA/Yzyq/AQzxj/edFO8/IhEg70foBgwI0VaL36I0HlpB6p6le9rn4c43
M5TEhkdtVLXFAytSxf8olKORRMKZMrkkG5jzm8VcJ77ETv8l/sMDucDJ075nW/Wf
jtIWE579toyCeGIw2aedskzPNZrvs0vyFiePBJ8Z1E6QQNdPbYPsobNEUc7QGFAn
oqPgZtLAnWnTiv/lksqFF442Hha+YaDiqUoG+zmRNQL7bf73ZAM0GM06zQ7idjSa
SozMGrtB6Wb24esyI0SLXy3CY7mbDm8KSaazKR0dpNM3/vqsx81UFxHJdx8+/uba
mFbXievbKzkUrWqL4ePghR+ru14Vcvi7ah2JjecCTLQjLDqykqCovIpbW+83Uxbi
9W41PyH8ooWsqSKItk8E+4G5KHxH2OLloUTRXsixcmMX0Nw5j9D+thhQQ/0xIcgE
rcV+TaQXnth1AdLK3wi95shWFInOXpWHsK5Tym2MwHgvaCJMuDaKOwtTe75j/GOC
SsVQsHWg4fsmIOJg87uV4WNmiUW9xurEqAFqOwJlZTeZ99tODyEt27P0j1+VaQX6
hPvuzeFwkwMHMDMDSRnUAP4Oq7A8YPTsfA8SmYrsBFjY+nrTHD96TBTbW363PtsD
6JrZyf/nL35YHmOucxf8+jcDhXnDs14ZwvMNaZhdeX+gOKUwTV3LoYuJFfvY6j0a
Kl2HzROBRKHGMam99oAIlzW69ynmzTn88shi/nqn9r7o/ONSIP/Qaq0Z0NCMwra2
yud1MB5t88m/QRrHtJpBl3NsQJCUNwO35FqhA6XB/8v5hNP1BDg4amsrwx0XzIsx
s762JRR8wDqUf1IKgOI7tzcvH/EUP33gA1J1mASFKlKNLpmzO/26THmRIQ7iHhIl
ude2L+gt2GvSCc9CDShwk1lup/sm3zrjxuA7PwutjeEu0qjp3trTnhWZ86wud0vZ
komcuYjYOOEw9PxzUrN3E6Wm7pFl43nNzDmXwUJeXeBkQoUZzgkUEyM4I4MW1/Ik
la8T7e8ZTG6NwwBXP8wniBiqFDOovKs5Ou3cJX3ssTCDsKnIr92c08iSUmWjQcru
JcYXic9amNcppp2JP8E8TlM8S5REj+vIY1QKCNrme1qOdogJ2Rc2F4/5fyeFl/pD
dOtYhMkQuAs1h0S8XeZdWTsMwXUzc6+1jaUgvG2Gl4MKEa65+CHdE9HJqXOTUzMc
RGzOfyggzz0XnreAt7Be5NawvcPyGBjYNemv0hkHjxmltg2D2VS2Byr+CxgFxok0
aMqSL+rLP+w0l8h2D7t7Y2zzSNiBNtyMuMm+jNHbvxbqBvwNk8OP4uiSQ+ldE95A
vcRQDIahyArUi5jPABTP+h3oBKLOsSim2ybkvfmdR0vKmc3Gvcs8jR2RmtH5Dzut
z56x/YrZkLJHKuBP/gWkEB4+qMpg+6ltMASeyEuBvxKWhTJegtdMPL+WthV8ghAm
ml9PXwcbuu0nUseYMGIHab65In1+5HBiSIJipDXVXkymjbGNs9wUUNtEuw/+e9KU
kKUoIGsQ0nTRwPL+ekWv3PYbpxbiU/iCjtRIGKhVaL+nQUVvUPA2aib8ouzSFtig
TMdVW/jc/YAOttPKpDKnjBFbT2J4e9F9Yf5KFmhQn/xLExAiHdIgAmiCGRDvUtsS
LIhDzAbPsSu2nhmy1p3CLvuoQboCnmsbuWeDP+NnWgoyt+h1JCUZw15KtabiOMgt
/0lZCABfWQJ248W+Drw6+bx0QyR13qdEjiawo3R5TcoG+SWqT0YQ6vgNiw1+uNVs
dRRecvezGJoEGwAhjQ5Ni7t/mZc5d4AwjGwzLSqDnzzBkRbcQRRXPjXspzJ/1Qch
mTfdcVYMgIICnHx0AumAXZNwFGGsdGZ/QAYWyC+JiHo1/+odOXLqsK10h22OmbIt
ertwE+3Bb8yHQBZFZl3E4PsFg0fjcFYesCG1AH+IrJnz9AwDMjFyeERGDQan/DB8
ypxDsT6XXbqWWl2zp3XztTGUq3tJm2fO1Drl2k/HdjVVWc15UtMKK6ktBwu6ywZa
WMghNSvDDLkLNBeE8C75ygle415y7mVP/Bi26aPknleZ/DQ6kkFkENPpsbfpYTIV
yUBsK9M+RehhE/dpL3aZqepSSi5C8Fr0vtNaEv3FY4/2QawhMdcVOWLpE2veh39z
Q6EJdHwMi9S2UpEmuhk1RuZuCYZoZFKxveSj+4n/NRVjP+XkXB7TI1mEo4xl9/i9
87xPEAMpIneOxlfpYEat8SZfcvG0mpxJcU6mlQokYgfCLiyFQGcTbvOLYC93yISr
mIphP+jrOLR5Z5SPs+Ua+FkG04Hh/SL7nl/ybjIJSHHVTTZulgqKp1kek0Yf9Koj
vnOzWDINPFMqs4mxP2wx7+KvifxSq8pO2aBGyxeBziRFeaAmTFJj9fE/+FEqqep+
OtNMwDhKReBan1kriNj2C6jalLPjk9EjssPUXHAtQvHUxFJHfeV+6kG8bHsRmtMh
smnvWZoAqixHawiGtEEwQEOblurbqGcy5S3BtOqpNyy9r0cDJ0LAdxjg6dOYI3h5
PQzc4fiIXPB3nTEZFpw2IPjeTm7hECBbM7lamtRwcFYZn1RfdkYaqdtBcQY0btbN
7wIgTBav/cB0pF0VJ0bjJOYuhZdSg2/+NODgPOcbGhAwctXwnHspCr4KEcr8fLtq
B7MkVVQp9MjMjeUx0WiDgZnM9EnqH/LC+xmMHuXyDTEH4rEzPQFzb91vy7jWzyaR
ePW5CS3enJ/tPiTdEMMJQ53FpMz7cmxIlQYoQaPgpJwF+99d/KHy1F5IsHKkRKT8
K3wUD5CWCDiuz7JhBIABxAN/YriaUsgzgXNL+Z3cOiyGCsb/AoPJoPnOmYRwJUNo
sHV+j8zBJG9wQWzYd7r+oZ7wkbuFToXqDWUwMhtRyo9sV0HOHtS/j/4I8KpkpPaQ
70IT5XbI0g77a1QLnDIcnqRuILY6BDT+lKQNMlqQ8jwDK1jhrMlLeqjc8KyBrAJN
TYPwtzThP4Gr8iemtW7wxxAboQGCglSs9itGvA+R110FP/CD8zKkE+G5MCgo2a/P
QjMgXDqffZvor12z6oJlnU3kyRUUo5X/unk02rWo0MZZ6muJSKsUBsp6B4uDCFby
t0GWmUcdwPAYJyGupoIEOxc7cMofhHUi5reDaCSNiJj5bRLe64fbNEgBqnlbUDpM
7B/u4JZY01OkHWsKeGxalam+Rzvtb1L9SPc1HRjoVo4V4xmqxIQs+kIwlQyrxN59
UQWqlLTX8sCoGF0RBkr3njyTMdQ07TxDBmj5zHKIZSKkpi0blLBUt6F67zgndtPa
Hm4FAxm/BXn+Latx38QRhWCUgWZBDpIUgoAkbA/d+P8TST+NtuJRlpDSeAyJnVKT
JEDOL4/s35NS0OtKV57vBkNEtQMZPsMhN7bv1vH4JiO1O428oY+KI/GDQ1eibpYB
hrMZkZVwQE9cyaAen+lc5NUOWEkDc0J7YGz//7RmxXRcSWzO5fFrCrcEBrJURXgM
V4ykl/2lhFlMnhObN6PrgtPXwaIWI8QJRPpmOVRZQz/5ROl9D91Ha0pAeGoKTE0x
50PJc2qi54s5mG05vy5u6xcGhldM5C7HH9Cddp2ARwNpNLyazQdxmihdwAD0RtcQ
p7YvRCdOCLD0Om46KEidN63ZrMWLH3avWrQJgX5c44gFU7CSWfblpRbHKrPUiYix
lHUWoP+STr3NkiwTZepbt9FeE7tcCgsQMC1kGJbncotm331KiXsR6G3KsnJGs+t4
9rsVWVGblx8qiQ7/wxwwYTk4Xt3vktXZHn5/Lsx6bX8wcv3BFwaO2ZlzAoF8SXZm
I3RLQMMLqnvgontQQclWEBlq3vN8NXocfq3cOezoB2QcCw7TGvx+qVgxxh23xy6U
zxz9LwWmV7OaYjBvhyPW6j8wyKxO709pueCGUpPzBGcMkWiuTlCqpOF+Ymk/UT+0
oLAt32/dT4jWD4I6c7Lcnud4+1jxy9alx6nvf9jfJLqG9yHUkIHdotWZhcxeQNkR
KCWnp0g9cSR8Scpil6k8OUvCQx9lu61ntDmlk6BMqz2UVVDgJLcUhmg+bo7OW22r
WvKvmQndQ51KCV+ESZGYbnc0HBkKfBau01X6OPcY8Kj0chND5e0si2AD2mcbZoxI
iIuOtcd2hIXFdF5fu5wU53CE7X4yMx6/uTeISmgFwaAFJw2fGQEiR6kGZDpru3dn
KVNdloAxh50bN9ztOBW9/k5tinMed30ZWy93VhmTlFNyygkbY0XLI/BOcfLE5QRa
BkENlMRXQklQmlOz19DrsRgwNRWfVwxOrcAVqkawinw2qBw9+aKAZVlAAMQ6xv8+
Ixx+2eJ7Beub46rXzUomZEB2Bm59iKSVcrt/AhrJp2mg/q/I1wVmZ17mZVFwS+VG
MXnCqeWD73M4+rBfu6GrlQqxwcBBMGRiBPFehUu5pbYwg08G9VOXlSs3jHCmZDPa
dBxz08pAzOYnsTg0dW78CYt0jzKzoPUFghzV7xdcJeNCHxdJ+dLHC+HBA8eDw3v5
KvBV6/uwLjlZ59vztyUESfbIW5Ux615uQQQRhJdAevO9WzQdiXDsYczHufzfsis6
bB1/7zl1kfpSYpH2xzxW+/EdgwK11osJHrlAfiiAb3NhH77PAIRTOh/OoH9QFLVK
7xs11Jmtfql/X3wRYy4q0vBS0YgNEx6W+RF3lOZ/PKVdfQ2CpBdi1K/S+uCd8Noh
tFdlERLDOH3TMobPeqUwD3j9tZcy5uCRUQ26CVc8SAhKFHmO2xnSg8G68fft/FoD
seE4ltbI9wWeeGqQ33r64vIaFz+v1/VyI0uGq8CxSEgeumeY6tueYxqa50uyH32y
JVo3n+8F49jrkPK9PIpjEA0/92cS1xOMhlYrivuC6+YbeeBuOrr/KjMxM9yiaxp7
ARBQKCQMO5Q6cpnCGq7oAOlkas0BsPHYCoNcz00Cd81/TIv3tA5QVVTlEG/h/UKU
NlfudJGhziis6kM5rFzv1+yjkOTxVqAfF7pX/eNWsZMZm4FCaF1rAUpu2q13SkUz
sYH7BpCrlXcZAo75Ayb74QEYi/69CP/FHbA0+mJsx/lB+0dLQ47PhHQg6Uqqb7ZV
RGuDnxXrBE4slGGjDc0O4kkUu8mZS6PKNwXkAZB54D58D+h5cSYrRHObHqvXab/3
zFDXXBk0CWQsBJpeq4C0s8gO9ap5PZE80++cSc0wIiYn9kP6OPOffm5+zGziaPyA
f/sOYhZV9HVOCWGNKZEWozwDDcy1Vh0Wqpel2vitDJGPIzde9/M/9Tli2+hHiQJw
kEIebScaC0VFkDunPEhMHBkitN/v1j+Ud/Eqm4WPmZAAajxhdEEGAAVb8eLc0dms
f2sgOC3aENLNp85ifmIk2jQtoq+l/YFPofT/sUH7R0u1BrvLLm37U+3h7rNEG4sy
Zz5Tfwlp6mGwU88nHEZWLqzHaZJhdxymlmrazfkB3E6ILFkgBzUS+YAKrywx8T4C
X+mPI1l0+rwz5UcmbJrNLAFlCIlbh8Z6lb/HbBKSke3czc8maxvh65oGXRgRuGip
PYtsnfJ7LjAZ/2ztjz3olaNuqv/PeuRJ+AP7KeyPjyIhR/PKCAkOWB3ZcM1Zunza
1Cw/BRZOYGlUnupL5Xw0s2Or0qySjjCJhl2dhpDcV0TvZggM4m17nhFeLVjA50h8
yjMUdZCG56W1Rh/SG2/OTeK6kMTBcu1mghWIkE01HjKzvT8BhnrdSiQEFy2uP3hH
pdeM49Zs6RT+9X1RhvF4fqSFXFCfKk6dLnRv4EJRiHQsc/zhzsDCp6VbELT5AurG
c+pObcouJM+/PjFoecjpyFUcr74Pg5WQ1rNwp0MyV3TTj0sxj4/jECDaI7s99U02
4UJwQX9iZM6oD/XYKFXax2guD2KeF/aAjolgNbdncVB8Xk/qxpFROwZuUnikCZBk
CjLqR1yqGj2e8+I4IOYLVADK3TS8CuPUuUwcTbiAVnH/MlZd7pV+nJMq9P+RFap7
miBnzdsknyoZCYyxIaXwKEFysZvojwFGUxfq/ya2Xblc4MpziJCp1YVi1uSVBkVi
vGA2pg6Zn3xxXOnDsM9mPX7je0LMshFcNiANrYlmk0To6wO71UpQ0Z/GW1uUslmb
CJpKAZWxVQDzo1rNvj8us3teJhdzWPsqIwJF3/BlhSe1/kkiAayAMKwKI+nx61R6
/UVGDkr7WS2Vk61DMf4AjpfjTRZGkmgBtzV5os/LoSjKpDS1O5jlr4aiCCIOulPi
KnzmlC7w/hhxLgPUQdxUd0v5aW5vjaIEqUuGMUeY5WiwUjbBOlUsN4OBqg4jvrwe
10kFj+gTn73ecQyk/fQYVsTT62lgpixlkuEA6JNoLrzhDBwafBLJZ6wDZcxEmLlK
tcnlxbQV/VGUxIx93ti2eqqFYAxyK9LwRemjcy2HE2UT2M5qVqPLaCEhKL2Lwv4a
7g5e9dwdevbkkWCbbEhTXidsGyg5dbpfDlmFFZDP1fe8vpjciRK9MGhgbV9gVO6B
x2SUe/aEJ6WS/cZxbh+gWTo6s0oSsJH3MwLZLr9tZfstgrOOYXY6JA+SCJZyjMCB
VnGizxrEm5wxRPzSASjInpTiVyApMhkXquqPCXVsbiDD9XQTzNDr/f24HvmNPVoy
MmoQ66oO/MiHRiUIYxUdEHEWrcJOTUboDPKL44nhW55hSAHCegYGrl9Vv7zNmXdU
ooahQt5GOuwqePRi5VW0IoYMZKGy115YHqi8FdJIniodufnE+aOGzQda6f4+5frH
gX6h1PxTmOjoYcuASlItGraYcWWkZGjiZy+OygWdRXpFIxJdhsxcND9fjqYEMwsu
R1nzVXRYBbc58hQXEFaJU+lEEojjtJfDTxP8eiuAYKUmaMS7cf9XeBxXDpnQwXzm
G8Gg2XH9Pq+WwvkfA8xDtJjRQawFLcvBUafv40kOWzoQzfivtgYAxF722iT07gBe
AtnCXpO2o5WthHOCzMML5zq1CqQOWk3HumZgsu8An2wU0Xt37W7LZ442ZEY8jF1k
5nUEEUTZwUU37bz9/XukOTHzVeMwWvhpyh6A7qfETRn/UCvZBrfxDSDRSZ6O0Hxh
ygIUO11/dpoVlbXAeJ9jwAUcOc33BMtkxaNFjKGijyFWf5MqGnoiyJaygjpXfJ2Q
WS8GflyCBXT2r7uXYZ4BRcdzpkFP6VFR1nTfG642wO3eGAgIbj3f/n2JhY+IcVzC
JYYeGkMkLCvjn9yUtCAl08EREzEHyDEU61yXj0dRSXuBc2rDHYuqebYKN7ncT13F
VRgtUbdjvGn9tyyV7XMACzky3Qro+M/O5oeXBdG/GWqsfH5NSBbjy9c3dBJv0viz
9kOI+tQkbwzigrIsdCxH6cS8+Xqq9ekDpvxj2zXqDlGd3wIxUUdNiuU2JGfNi70D
yCNqkX1fZ+Ovi2EDAAIoTZ4q4FhJaQiCqysW1+uWsq5YtEDjybataVe9ySaaDF99
VtXOtSgAt3w1wJeQANB/QrABzGJvvyz2ojA37wPio7IQyjzCDSGTa6UfciF07p3N
1RWMlaA9VyZyS3lBeKqtTvTUgBB5u6rVFFqW/meQ1x2Sl6DqqupVd9pKLa8+vEXq
0fqPLsMvhOuRchgPUJsFLnY/LMcwSzHM64z6HxqeQ6GXsBrhpLNrHHh04c+F+5sc
3fFHobrZn5eB6vZWiYFhvBV8r9FH/JpcwZ9g4gE76TwsING3p0JhcPcBDO1YVS6R
sbkCy+pmCJ9dvvEv4m57vfL2GVtg6rHI05LeRhgqV4dE0+TblW5M/hrawQTYyhm6
3qWUEI3WL+Et2VH9NZPcnOrkss66puIgcOAOPKOPPXDWwIukyXV9OsHnXuuA/uMu
8ZXZnQgmerk9/Vwo9PZMiaE6n/BitHenHq/vnS7RM64XUka3gKWPow+PUvd+3SWd
U/j8kbndB7Koeeed/bZ/iGKf5/VvteWZ4ie5J62fQ2Pp3U2wczxK2jsikKRVGDKV
GsWmoKs4Vxk4Pjf6WkTmmiiuIUdnS8+umYfAKfMHSL8BfM9WTpxDrmalBVZ7a08m
heUyF1/CnHqYZT7xCFLvUDochp8MZdNtmxFl8M53AFyYJ8m63o0f9kyGyG7CXfEU
6mMLEG+meDfdpibDbwQgCeHZ5+loEQyVxwqInadDP809vRbDaiDjmh6tPoyXw04a
tz4R1h+6hkHDjAB+JF1F/7PLlUTewG4ae0kFY4D8PwF8tqdskAKFxmJYUkY8KdxR
eaAVKSLyFylZJzHH84N2MnzPA/LPljiVQyRGb4acgmn8JeeBuOmCzNikv7fTEVh0
oxlTuscjtbgaFEfWFoRGDOcqi11Bi2aZR/73om4AvsevjpTa687nYeIqUY4crqJd
+DnUz/ID+5kiX3mcKCL2WMErz/+Q5pFXAH3isbvymj0ix9uZaaRiOXzHfS8Ge7MG
H6701UlCxhEoolSEVmmtKJjmZP4GHCGV4WFaHYBoqTLPdezMfg1/gccWsLQlorKE
FHWtF7xmz8FhNZtpfQA+Od/aDVbZLUVRirESeF9HwnWMZSETLx4KiALMil2KKuN+
ED/DCj5EKdGGAZXCAKoqN25MDk7T7kx2rOa4I8fRXWjRcBPelDLth7nk1bAVJHFM
hEBbqJs7nlxSIF2HQn5qsxv+/logSxOw4603CeYlmQ+3XsKsRlEJmDVOHEpK9aYi
ET+xwEu6+gpEtS1vB5YeEl2g/INQNDzwpL+87DjALj8Xsoq+oZNI0J9jeq8xb+PU
oXfwbqIzd0G6k6SU3/dly5dURV5nq0xrgd8zvYG1GoHkegBgZX8zFW9IBdw5SKZP
heaxDCODQPGTu5ZAX/b8m/qjGbV/nlW7/qnPL48Hd90iwAJWgJD4qEDsal5Dq4wi
GgSbj7m47OWXZfm6+fjpJC+uxmed0aArQAyGGn5eJaVEBHlX59HdMiiNyFeuK8uF
16AfiieJqkIm0UnHBgnrtD3Y5Lx8cX4Od69y5Oa1QTL1Ns+6E5wYFU3UnHhNNG9a
MiOsucO4hCtPbImUqkGCg7LHOaamRWZ+Q+6cu2uNjrpVzY0TonSM2cvfnCD0EO22
+EVidczjra+UIQJEf7Fckdn3sEuuci5wWKUuoZzY3Qx9qlH6DBfgBu/td2DHQ021
lnYf82fY4I7mPKm83apt/SD2GgdHy2UNtJfFDkShoZmeV2usf3gILAn1QyxCt3zz
/7V87gGQi9HOJH2q968ZYaduIVDk4FqT5yN6wAzaf57VI1/nURObuzBkr3PNIX7u
513ZUJNHvGnr6LVfWdojna7SxwslddnS/RZSE/OJeP31Js8PWdZWdGReV/Qz6vHG
IuqeeEr65QUWIfIBOUaIMA1r/fVmUy+pPpkn1MPjlwjpSpPTjF8c+ags7e3/Rcf7
cg3zUVaFCkSXlXTZBbzbSPYuWxwvL48lpWMGr5XJhwCzm+QtdmboPsbSHMt1xh/p
ndbVz/h4l/wIMhfOLfpDG8fSQ6q4HUPmkcoB6Foau/tAZkk2Cbmr93FpoVr0arKl
k7qiG5kWgdBnzA6BaxYAL0Ov6nGhschAW+avGwGzSzb+j/hg4z6XAs2crK5P23Z+
rU8dgM7uqnET0i9mNPGowuXft8GMh15zpeltVI0gRIlzE60xUW2f0f5af9S+ZeIA
KWHZglLMk+SpOoUxBqntPI6ILuooXgzYgU1MnlkFOqyl+zZbNDZZI0Iu51JCBo1Q
6I8XauIBkoYjh1BDPNYR1sJninhpGtflfW/j61gGEf5t0zUfLQMf8W3IaJ4Y14A8
jGkjVAbvGeMxt2tWxAIV4SirRrsHlcvjWqcwCY+KZLCqdlJir3gfIVfdei1C7hLr
bS1+qGoRXwaxc4xmok/v+Pu3FgNVia0PKqLFbgDfYsIwOr2pkh53nAJanvxrfVfZ
Io8uX2Lh15RK/vsCdQJdoBWNmUKI+1BnaoA4LQxlvElNxNEkwCVGNQ2eqMD+9aGL
g6v+pf/sx2pVWg0Qc3unrUSYkaRmUiCpu4BphQDTOShLdY1mYgMZTZzptNSBsWZK
1Rtscu0M/eRUqoKCfedVA6xRFxJ8Dlyh2E/vOr4LEdPHKu+lTbPl+N+RsaKCOCq2
EEFHvOH4lPhUrVmt0NqUovcnczYRJ22eF0eMyFLyDTPFH0KHroDoVIsOljjqvtxs
euJa3jSeky6hYIRvfaLRNTRPboq5Sv6d14UHv6+nwS4Wvi7izJkfVUgBmgbyLKgy
0ayXFo+XlbvittRN7ALPBpJAslmOtaVdGPKomRoEobcXyBgtex9djgedWcjZ2rLv
I04MCz4yCG1i6RM6oidwE+KDXF856EGbEPL+3ylveHeRkQo/pFPn9TbAxtIAXPHB
MyeJHAscvPhaPuS3zBdASRt0IZgl5U2xaWjJNWc+QQdwvNEq2XqK3OGPcFpil5gM
GDLLMb5YykFF/Z08APg8AETyQCbtuttH6+uUwu2HQHlCSrX9de+Hi7qO1Gpt8L+w
pJAxQrNiSApcn2GdWo4Ucowq6B2srX24j9WNm+xLpTY9L46UKLZrHRZhK+aQBqh9
9A7FySfmt3tX5MUFLhqGOXfIWeWwrrinp3aht9AeL4lxpBBD1ovxmdmckozRxVFT
PTBOuU8AwpoebR9FTY8q8TX5j98HscU63+veywJ+vkxZ2IKtibDDqN/oxVJeG0aE
x2SPoSpKXDmI5CNmXKPsD3vjSOFmwWVlBPhKtSbC5PQN355D+TfnMEG7wYSuxoH/
jjPJFMgQ2936i4O5iIV13xykKcTd9ahYYyqwul87CzoD7PaaS5CM6swcWOZQLE8m
NseseGyaEaWDhIvT00B+tUayVXc08WviP5ph9c59INYS0QRCgaW7fqvkhIXyItDS
SQZTs+HvaJshkmyU6zWtCjNumvI4wUtFqUbLbV6k6VP2WB6N+0Vdlihb60/wb4TN
NPWXaS7E1i00J+q1NxtuGUlqVWeSCljfTyziL76sPdY2KF+jOzzzFUUOUtlgwQ/M
acC2qWx3y3zxDHM8FprnfweAnlxybMQHV3ZzmCIocjIH6YqeUB3nmyiclDdjh8NX
NZ+IGAcIDqTpGqiiSAncFkafVwoMkqOtUEvluuSta25OLZskz9g4cdC4pqYYWPpp
PC+uyPwqDsnhFk0jPRY6byhtIa0AyhadxS7GpT7wXbJUOsejcwp2/ZoMDbpedOLV
be9KfA6KyFD9H4ppV8B9bhFmLT0qsCf5YdKscJb9INLqH5Z/5SFNNF2gzHDo6ofq
g2ElEGisTP73Stwlms+ZQWQ9fYhOAg3d5iTZ/ScKFE5GlkBin8o7WBmTsJt7RqGj
97mEdS5FZ9IUDmYPisShqvREyCbFXSV/7FlA3RWKWUpjMt+8gqj+2YM4rZaaPJYJ
JIn37BSZsvU6ThPigNvLqs7yEQYo0goYKJYKDGCoL0NwT+FtCp3Sn0R/3lfFT2wI
pXvIayhS5YOy9xX4QvYSG23mwmnzQYZCOv540b34LY8st2vGLaroClcv6bUDx4rc
nlgNWJ3pvwcfyw+k38YhoDS1eXTG4ItEp3dN2ynlDjc9kQNizQ2Zmo3ncYJH4XG2
rmflEE3ON+/NPrZYXuog9ym4Qw0u14cWgGFbmhtokAM1RPFOB3xlTB/Xlph/QPHC
2rJT4d2+PzvbDjvHCGYBNjWTaepCUm9esx4WRo2OXN08YRULEHpPxFJvkqpKb1RW
rtmhAAIkuf8uxShBCTaEdf99+iSkdsCAWFdVH3U9Yr8WIIW223joeTHU6j1WLUJn
FQi/J3e8eDCoCG2Hq16ElZ9wiEcruIt33tGIpy5yGkVTB/BiBs7vV0bIYVIFlwdn
mk/4cvDth2YYWo2jmMn+pcSE4ALC9Qsh/g123D4o2CWxyhlotLrpupV0jdqJKDNl
csWAFAVRoGVGO7W+tg2q29p+eXZTZzD2MxlfS8a+r0WnVDdK7tMRWA+yODLSi8Kg
tXGtSm2bW2+vGPt65vLbd3tCnyWKdbfEV+clW6UmR5mKXpGTg1UpNRBEth2TGCAk
XnvtJo7JcAtiJNE26GkG+L73UxvS94E4XhL1r8R+nE5PDIsDDRSRYHOPhee68g/A
PLZ3tkGuJoNAP+D4dWlFy113QbQBJrhIuIUErezbQMr5mDkd8QYZU95uJ/qAJPnF
CPI3H1rc9j8U2L6qk3gdlQgxDEr1lGisB7PlXUKT33TkUkrpdeVOudA16Zpwilkc
rYcRsHqsNs+OBaLahNCFFEmsZ6eYsH6gh/7nytjiDEHfVsBM30xcPg709c6TpU3/
iDSDN6BSi/6aaPQj8+fg3AKbvD9YOLJtIkJI5xsYe0iHz6kwdixXoGdyUiqVk+by
XB6BOSAvL476NJCoN7REBAAyqpGvBcWeupJeQpOuDKb3i7Cl4ysLHWLX+Jd+0wXi
jAKt0L4gyopAEKCqriFFoH7mkkZ4zEq/gkBAPGfk5Za4hRiA9TWciOpwEwltEVii
NAbAeELLxez3tBBpZZ5dOpiY9wjtcAIYz2hZunRTKi0yo6t0xj3HIHTkBbAaTdeL
3IK6I+1IJ5KwVBAYvo5jEUVxWX/WubQBg23euwB938H90VZ6wvy3YA1R44o6f+5N
4TXkV6dwZfmOqsGMUqtn+jB6k3FaDP80q/8+brwoTu3DdaHwnqSc/OEtBOyFzsXu
1llxa3kgm0yAWEf5df30vMVyazWs0YmlTK+bwQYisOqBTxLPdmcY7enDxDUidmn9
yjCGX/MI+oiTWuo4Bn7wIStD/XV9UZyjixlxndjk5llLTNQqNuBJtLxBTR9NEXbr
FD8+oQRjLKelhOindVtIfUI4JnIdXlH9h4ysxC0XRWbSNmV9a9YrOPW6ZGlRaMnf
WrbK3outIM/S5SS5BcQMvmlA1ELBG5P9fNT9dXVPZzsRulPk7oSRv5ndjgpwTl2D
LVrYHOnqEiV2Y4C3/FiDbiHV2xMwLv8G3RCENmTnM35jtnttnJOVBkTCWPhBImgT
0q6aq5sdN6uvRLCxuBq8PyeX+wrOOwLEl6J6wEt7w3DgDVoXDwqtRe+cFe7fdBvX
DP3dON/JugZQRAQ6wTPV1uJA6LK2HLad6loORgXqmLzKwNh/sPvKiBV+BAg1qSt/
V5w4k+lWvnt5BJwuseS3GDlPNb2BPvHsu+jnNrGBzs56tBBguQnQk8HKk6oByjFc
6uwW9b0Ni9xUOxqEuKTumQk1QiMi9O9quPcsGOe2atghHkCvAXYpYKSOJ58lyg/t
04k/vbs5SKabJXt01P+Kym1eXsqmOuqm2dQZkRs97wxGu3Wp0Rid7UDyZAWsDouY
dwCssc4E5XfhQ4vtdJ6SOC17aJoNpJo2MnIaTb5asBx17J6QRa3np3gHXOuqFG7t
t4GmjeSsibJbLRwzsjByIAISZeUB5DT16XQXucRn6t3v+WcxRRpQB/voJY8Nj0tp
MDZS9A3uPWDPa0hOxrfs76IKm0SNDSufBrWwye567/MfBtWPytJsDbuaClhbmehG
d5y8lQxkdtvMqWuDuknaLWGEkU0dM8STHmX0O7ufYV/9vynGL26vjh9CbEP0eGLX
cRBhsqVRmsVDgIuw8p4YNLyuaWdIGLOx+rweSzz1DMwWOlcOKjgd5LD3JnSQNvaT
88wB3+o5hAIZqf8J8q59OJwSceX9X1jXSUZyYLl8HaLW3nMJDnxiz5sbw0Ct3yQ0
53RGyvYFLuRKPAfkFBfkJgb6UpjrWAI4lZXS8kXh4Ydv2X7cXRjY6no3KmKaSHY8
s72jpPJtVAoAYBvsl4te6gh7bVM9rSlpoo2xBaMUSLkFKnHkon7nIGUZ3O885c1x
HN+RnMvU97cRcoUvUnnWIOcnYVnWhVriPmP/tdka8/vPAOMoWFLq0/Po8JPdpMK7
cbgmsijUyUWtUmEQ5VA+fuMvihDjjPu4eny3DnPf1LonNGzqaPGy0IlO1WHE1p6r
gtTJ6jkgysFtNo8Ma8tXGDbMQsKBMo5jIIj/SoTVfSBwOr0MSH+uEXzMz20N2QhT
/twXcQeORKhZxY0iT6+RvKeLDto+x7733e6nnSDSZxhBNmK9+20qzh+cF2CNZ9as
8r3LKrx+aDhUeaJbDVCsmNICTYXgx6Ivaw0r5GyH9zvTE5cErjaeEvHX96BChJQZ
NegB+1PW/okXx9MVAJXlMG22tc3ML7ScSKiILIfDhun1MFp+3L8oGia6xLmwQAlZ
uZFWfHdS9elKPPa4lMDTplMP6jp33+LjsyvSyD/zFkZFd9lAOQV9qUrN77S45y+4
f0yM89ukCxQZszf7UxOCDl+K4GbD+o4DxPn1t/xa33Fsy/qmmFQ9LCna411oAUmr
CswhluogoKtylkjSprGAiViz7VqutFOJzvRKk0Mq5eA2NYaSFtV/U8cXcfcRQ/Db
LUeBKhOfU5QrD+pwPtojx91+bj4z/MBZePtNJWYVthv+Q5JTCzM862Fpt8+vYwxy
QDEH6WQMZaCRCK3ZuLl1mF24TURh95ov6uUlzY9mX6ON8Rbqb7YtCqMWeTW2zsv/
slUuGb96FPKzRDeEu+UhPsrze92XD5OM9vhGQgeO4rAARvaIxnEPMy9SPTcMMsko
G/juSAvrNDJD3GwCLZS4lnAnXtHiQ+HRE2pK3sqecYXU15WWbZUqyTUMhJOG9xF3
V0Hv4rJnrtl8Avcwel7AFwwaHIkTjQ22OH/V2lGFJReUmFTvoFDgCme9mlsCIFMO
7FQuYtECTNLrQn+gKCcvI/2TZ/AbeXrW5YBKxupiGBf+2ZvinrzzkbK1qmoVTNUf
Iq/nj7KnmIBvO5OeEXGS1G0GJXlUHASAxSNdc9ay/Qi4H3INtBu/2gotPKxtVONH
BfH62pE5KU5CACs4GURRcPs6XHSbs13f+a4a6hDNQxlUqJxNldDNDtffhE1jGtrP
tGeSCCZQWlRTwx+WL3+gP3nsYcObQjnMoiWiDwUasnYHJbnEVK0MEsiqSJzTm2b8
YvFbid+uZ6elK8cem/FQ29a1EwwvCzlPqB+bjNROJkmbfn/MCUR+wtl1O2+/5O5Q
cVozwg6POnYT55Ez0xyG7xbaVRc5AbrksnmqKZXcYSm9XURp4fCI03/XsLcEaSi1
HnYryHJ34bR2cabvl6V7y3UHHMk3vSylY2kdaAHk3XXYorMidq/bebUYXY/HQ/qw
6y0b33qxfKxbmdU/UVv1vyFiu4VkC1G/GonHQu2OlqosnAiXQok+niX3+FL2ubOB
AryY1k6Q7I/tL7N+7PwGL9XI1yzEKdtRKqGiXMZy6HEgysNxIMLVUs8jb7TEMcP+
8lQW8PyB6UxX64tWgq3PjVjfQOmlNN97LNzEjrP/KuaK/YuHVix25ge0BVzWFSHp
Q0zi1/fKEw+gLSU9UOV5EMr2w1GDTo3a9GdYAVkWtyBMIxzt3EGErwncf8+ZN8j4
6MhrKMjyRvRN8aXwlckePv365F6V8Vr8A2+8O6leVXKhtBRLEJCFd0cbFHT1tWSv
gU5JzeAr8yDnwcXOGzlIMuhd0nXSaQ4pPrM+KOVGAzQM/d63wTpe6aCGSN9utzX/
lB7P8pKI9JOGkV5IgoULOi/a5NiXV/EOvXz6HUxnV+e5vtZRNJKI6PFHg9mPEuS4
KRSYfqpxZvrbEaH0J58pjlEajgILt6sFya3FjYRhOiLWo2GkLjUF2u75762+ClAo
uIzG1b5nVWcuaZJeQg3cJr6YjQjMMnq1UksmW3EvqjBtSm4xitcbP+/dMoEmER26
MTACzqAGZwj7iapd41ZSOD8t0vbkG5eEHmKz/1ZK65+BEcSvKhqT+3ysS4PUKfZW
tP1zy6Z/46gWzQPNpzstx3ZM2r6VWJxNBaP5dg7dS9vw/q51MnWyYD3k3JMlr96D
Y/YQc95CgTGffAc+CnTqnfCB2WSV4xf/cv1Ehs7unpr1RH3NjwM41pto3lMemo3N
IMtFssjHwziQ+A53ocdhIve5Mt4ujUGjlPRHQKjw8O5hBvV+KisM/9VEi5iBfoxS
eN9IsylaqEGsgTennusRqBenL7RYpEcgBh3B5pfTqqEY92uBpaHXrgHQiAzA6tMU
h/zOkgXojd+KAZDPoQbrmtZtv4LsAGiBfxK4K96NH2ESFumQNkcApvw70DBSOjX0
wexLSdaMS7Pn779fbmjK5qwDs9nAkD0xKiB4lk6lfBoxeC2+nljlw73YI2/VC1Sz
YCo9yTv8turLtO/t9bn8REsVW6XVUAkHvmJ5Sfbx6BJ1TA3LBw8xoDLR5/gFG8BY
DshkNiXjRzc1iU7KgAHQu2boudku/wiTmIe8s4cWl6Damig9zYC3KYLyeErUkLA9
iy6cC6VPMUlrC3+7tS+Osa7mVYXokNrj1ay+AIeHq0W4zTfT566PyvTiHcD5PSxe
rQhyI9KGNg0CvTG31VdKwUbnsjKpQk8WF0QlYOu00M/+M2s3fWowtYnlLzmYRUvQ
fexTQmgaAoVnoNjOHUgd4Bk1xKrItlp/xzgkwgfCgEzV5BBWacBhW/4JLrD+Uya8
H00sppxa70KxDS+IJ7z51etHtI9wHQ0J1i1EDSZ3xeW1/vPHUSxr4lZmMzKiP+ur
VkikEGqafBjyEm6mo2dWZz5MR8HVZsGrn888pQcvljV2Q2Spiyuf6uu+piyeWFS/
SoikdR6zgPouf2XRb41rXDMtNaNTvG5Z/TgblVleCXdL3aVfCJoelY36FNmhUcMx
oeWhNJtd8RV2tCduXgEQhYLXEymDg9QwR99EOvCYj5OYtX2wGT4FZ4CQVp7MBNHj
PtLCRxL48iduAuwdIinmnjtEaHDU3Dw09ivFm4bUl4ZEypk2GVSv4oGeuhhCutpi
qA/a2jhHHGMzuUSOCluSsNUSlg6e7bfigtp0k0LDHzCyuNyVwvn5N1aPILLwcshU
VavhXFW9/Cpi+S1lzQdbtptfYzqA2IPolQZQlB3iioboZ0nNx1Jurv5vuizK4QoV
Jn/xg7WcBTIz6Nisjv/j+Wn9APS2nBYjmhSW6b7bdTqLDvfeCBZp2ZdN001kE+YP
eFMuBA/WPeRWn1bFK+Rx5KLxOku563VVhCAPVrHBMIdAk6L/9e39OkXUHYi1+brR
3zLDkCAX+QAdri1DAmNVeyRsNSojlNg4RTCn2fqZvcIiMDQBa1cMXNMvmTK8xUIN
tgwRt+L06jDjmGQR4b6a0rRTNzrsQjPOnX1M64IUtM5YDNfDCjcX8pleL2GKWbcR
dmG5cVNV8TW1Cp2qOOP3NNVTUpP8j9Ji8J4mXcma6VkKr4U3bGs+fFvKtnov/FEo
06z0NPDkqEphmSDgWuJWIOff+/fuYn3oVW2y0w3dwlMTg+kIK8m9BpQ1G+HuCTHO
g++mXiLE3IU7W46V0hNLF4pridFai+fkGw9pzdMT5eFP15hkPlpLAi5O0HhcmxGl
3AlnBYXXyO3rt5GbQ2KvHVnC49tQbTsTlwrj1XAgsTCFZBjLdyBssgH4/X5jevZu
d+p+gTZmm8HVZycaMhMkmfoxAnLiFTLVT/PDpf7PRYTEmd9NKQvmPCLEuEIq9n+E
P0Kh9KHDZjKV/vuBuXd+j2Xg4WfhA0MIYqBi6H41rONRT2zkXQ4MiRucsGMdNFUN
dB/2z4TkA1dG8VzFRPPw39qNFXYGtayNlWLWgICOTWDquC1ZGks7KiKOLt2uat3F
bvTIct8Taw8Ztq5eA9jlq0f+BjOrb4d4tKv0f/KayLKg8I77ROWqF3XWXnEATlF1
JxkiU/ESPd0JzzlH0QDUYIYMBVLapIVB2Z3wIqH6/taTutsrW7ydkDG9QT60enVo
dSlhNWuXaDzCG5BY420qgWd+YYRO0yRONxR8lnEhH7Z54hGu9VFo3mzXnjBLYnnm
apm29jG9lc0XOqJchNzOMbriG4/fXv9EmIjqM+28EXl2aOvme6bBaMpcggcL2Kxi
Xz4A7vnVgMt7Ig+qgsiUVzKTCdP23LwZVMAae+Nr9hnWcAIocSDv/zWAjf/NCRVA
elFItBmDQFedga/vYrLMetDeJCdxeS4zId5G82STYEIrmTf0q486fEng9ok2QbdH
2Q5DEAYxhnxiDO65+2k3zVB5wmXBvCG6DZtrqEh9GhHmqYu+mOhU0mbdCOVN4jhx
wml/bNJGEDy+SvF5KQmBZEpBb8jsimCDZVftRYghNIeBuCUharNwUL4r6r8GewcD
3OOQ3Wu82KW8zkBRXcfYalSH7CEdDPjgaoSxTqsxfsgT2pRnJAKDmq8G+y+phjaE
FcAMP6AdxQd/om8inbcSB0fYbHbfMZkWfM3H0z+X5feTHKVr6S9HUXPA/oe+Evzo
dSsrKfmGwVECjoqmIIU9HsnCeI/kwvDuQMhhoepwiQX9BXDRYAXh5khJHw/VRy+7
RAb7CbU+6bLXcU2TN1HXdBFbJfESuWgEYiJoZgK6CaIUmjMXTWtEjYdegWcV7a5r
yRmFtxurAvECsfew3jTbbeOPM52oqLUenWQ48SVDB+wWqsCaYP+2Si7kplBfYT/B
wWjY6p2amrYAXwH7NSNJ4Y1zneFyBPPT0Q2C+4fVFAc8tLROxBCY5W5Vaeg5aAr1
702FaBQlxEIE12nUpY++3k/pgdjbXCexpZvrX5iz3hdficsA3+erxDBP5PnRkxSF
nkpN2lGi6ajeCD1EDTxz7rrUtT610YxKeu9FztbskRHAcSLCRLQ0e4ULIkncwyup
4kBEUU8yaNddtpgUyeNsXUvw/l0qT24gYy/rMttgftsLy3rd6cWPN3Pmofpr85W5
MzZ9rfIaRUJvLcKmOiheIG81a17pRU/80e+J3hfysc8ay7I1vVa29L+aKc+fmAys
9MZkAIA7ehxajBnjp7XrQqSMHklD/oCjXEkPeLMvxqb25t+vJmDrurPPz7Iml1Ta
F+P7Ko53h8HwrhBxDRC3s1qhgqDCvJwrhmAd9Hvuh77FUHVjSphJ2Nqel5K359qN
f1T2znbqvPCFFTiSb3nDwUHKGFFLR076BuYwyQxUxq9DIUr0zjnrgsraaL0B5Se5
rwwT0V6Bu7AAT1MnpMC7MsFdzd6EPHVrSk9hgIuOai2nuetzDTPzGnap6bCj08Mp
XAGXSCPbawMUCxl2uU6B4B36KQ63xU8a/2PQ4vi4dkjsyl4dsBHPNAGSoffOetYe
GqOTiurJSmOLKYdhzkMznc5NGLGO79wLH5xuLusxS5/WoJbpLg2cvWuGhEwpnduW
qM1NQjhWOd3TXtPqm/ZHplAWYcgeAkMKK4x+m5YGJEWEqEMmatT8BK4E+egAEV/7
kGuviTOWdAzfJIx0BseQW4fzvsx7YuH25MYCt/YOjMPTSZG2MOBUjcScCP1weffw
H/AwxPctzR2ngC8WLIzhZru05JMQonLaYzXwe/eIZYngLXpM/Z9/rktj58Z5ZLqB
2LpNrC9ktJLI4uLICXn0mCDXDPSGqgorX/sGqmA77C6PAzwUj0YWmPuC152uFeF2
+FBZFuN91+6bruZgAgDH2/RkcEB8kitPiF8Wlc7BWRCuBUSP0Bvr5P0nL2We2R1a
Q13sFlX4ERb+2b70ReMXmtBuPSPxRyzRcoY7hc0XMBWgGmhFXjGtyaDmsq1MUywq
A2Cg9CZpdkrp/ITWzw/l/gE0+RTwN5wnydMEq+cwo4RmRoSEGgqo+8mCg+1Y/g/y
N6vpqf/45Y/oNSGelB/OKhmSzbKPnBRIrPHMsFbrfqUAF3Z4JYM2t71F7w6JD8Pg
3vThqKaLfxBWP8ATI5acKFPWKAT9z7hmqsp1P6njqUV3gt2iLBJCaEP7jqGmBRyg
giY58gbZdfhNryffJIwbrXpz3IPbK30vmpElPqkbSNI7zrAJEkDQ2rEkxpzlzxgB
LIIJe2ImQJu3DyK7nzQhiiJAMGbEvpWqfCJPsd0KjUYI6WC3fpkpeLlbpMy4sVBJ
TkSlizWOp5rYV1zv6DVEHWkqayvCIK0gzLia44g1rrLZqY3S9m4Hce4orY3mXuD6
bK3tWUMQKlrCcpoK6qvSSCH5Z3l7m9Log1FZR7lQWkvMypDbj/jpYnBQu65P8NR/
Nq8LfptLOZjFDGyZ6CvsTtQox8ufmGvRWY0rSyky6BRvKYydXgdGEUZTfNHkGmlp
tphVE772UOuo0nsMf8/UBPnIbD+qcqeLfk7QiSe40PuV/jCd+Vv0TSBAeVzGQwdu
p3SPq/8dSEKyD/CiT2KZ0Pn2jNfW+98q025s/aecZsYXdqUCjD+Pux3mnAnXZi6W
+EnozeHCII+fktMisycSBpb5/8g4acLWqyOpc/oNTMJiHDbV1GPfcX+CyQifJ3B4
hwRuVfM7AgEUHTUCD8Z24si+j0uc4/xYKUZtWLU9V7gCKUjBgHqIJptWTZ+yaHxZ
okprjIt06Cxgs0kNvSVmbT6JqVZTFMLeHHbA0dSKLnXiUylY+hGqzTsOW6ZJZQNa
zNlMhJYtncgAVhxkpw1CkR6f0sYB5puXhk/lS63zsShNmgDY3XM7/sDWoZsIvkfM
ZUH/yiWzs56C17KFKNmaHCRRGuzFKfYQG9WBn6OX5wkGXuvwli/ySsFSRVcYjNnL
qjsbTK2cpLSCnE5iYt8cZUWVAOGxucZ0DBcROCQu3z3uJeCEO2lLCR5Obnl+DOlf
eaCQ48SzCEsmyGk26I5/nLrCIE6Di/8gQLLdS2WyXaVbF9YYWEUyViXMl12IPDv2
Yo/zY7BZDacPN3FFb/POCAVlB+OfUzIpkOI21EEbPrA2Uk2h/wev5ZqJqpPXMJIU
renscL64kkSNWNpag63xWeDRyDWIhx5xvF1m0nhF3QRvsTu7MePaj7aAjPmsAizK
ZmlhzSTaw83r5WHrtV0cwAx1QY84J1ktBFsP3jaG571lCU7l5M6oGdW+9XmcUS5f
MA1Cg2b5cwlmkFlOLT06jqUFfnArtc/llqbXG1ig9qPa4x/OMZ2K3Yt+o+Udwgjr
wa9jUeD226LEldra00M21WDZKXnG2qGHhu0xYa5CEYZWM2l9Ba+7+hvBkz53uxtE
LqqvDoeca2rZXxfsj8k213mcVccsWIyvbdTrgfSErWx2Ee7kLOHtF7iibxVZ+/c2
DPr24KrU/Tkr45BtTP2PVAnWtuauYi0MGe5qQJEkyks/tuOuS/L4cONQ3hvmhsju
n2ZeWPh6QzY3NMaO3on1W0SDT/RwY5sfxue3wRXltjE0NsaVq37j73WySjech1Qv
yfJ4qlH1ZUqhzy2pJQ9W6GXjHLIg4buWGBhT1X5AmDEtOIghQBAJZ3VxNyIFUGLI
qmkKyR5fmyRdMHG8wIODyR0Xjt5+BqNMEN6yHhyisOi1OPzb6XqanPfytGiVArZR
36VNoXZ9nkhdI2RsUdVJ7cH0uRKB8qXxIPMFaqSEy++ilbKLb8bINdiwyeQBBcaF
meFAgvbTfNjrKPcll4n1kF7rD6nt/nUbISEA+CXc5YQb6dXDpszRVeJkAZz/mEVU
xfuQAQqyPl3Q2xYqkPwerBpv5kOj31n0CVLxkxTrWcWxA2gRS0aWMhmhhyqQjaPm
vxhkx0+gmlsxg0RAZU0lcXCMiCh9jySWZAK0HJl/Q/AJZ+xlPMCH52ui4xUzBMlu
fb/1dklH1ICs1MORFrRdnht/mahsyQjfoH7oBYXY6N3v8ntXqamNUtf1KZ1PbX3n
O2kJXY98YqIusCkaehdW3fkCqr1Kq4S5LAwMS9XDZK5QT9IZYQ/fE+18FAAzjKrY
TtnpBLO9W9h5MW3SGTMaYPe2e567OGsl6YwEUwCa/uCTfvA2lgN8RHP0E455POz3
Z1o+0dUfbmCdEo5lI0LR6Yb7w6sdc99F0+UNfAZJCohfukIlXYzxAsHeBJmXJnhW
wFc1GU6MRIt7b+XdNOrX7JOj7n0rGEpDXBdqHUHwCOip6QEuVf3EFFZlr/oDvA1i
sopBCF0gpX6uFeuHP9MmVQjw0dQRTwQk944xgl5o7E0h7cF+ZLStTlU33KVVPK3T
J6JAk1JYkD/SdJpSLxEStSYWV/Hx2ed5ZoeP6cbE/aAZmmlmCE2B3vAJEZ43Fi3p
uVAFEkqjv3m/tn+H4WJohCnzz2TSlw6PALFEKiWFettZ2mUvU75qocteLEVdM3ZU
ryvLhBtjsvyOE/sqxRSknCvZ3hJoiD0P90ZmqV7V1tWGsu+pwbGxVt38NB8+CYsJ
Cc33O+wIc4r+6/0no9aFf0yfY0Jr0aiC8ooUvXNF4qIE/AWy9IzwlhLJqbtJA7qC
4wlkwWfxUUYKwzDcygovFtAqeuaF787eXdnDkjFDpr4ppBWl0baARxgyQpTM1Wco
wxGT+CdHDBM9W0yezlYBZaSpoK2SPNcPBcdjH/8OHGsBQXsgU89PmopgGB2qEobP
k3T2ovxGMnnA8lgTnMngpK9LcKfAHkmPDaEchgqqavkRVEvkiFr2TWCV6hI5S3io
LV9agrlPFKz9UWmcoxw7IiJf4gKre9/T3AFRJ9szy8lhOy8BA6Y7RUBhL/3vl6fe
NQ3B39CMcuKWgE1mnC7qP9v1fuQIKXe6yuvt5rPo+gKZtlHmaSBtbNtZtueN8tis
Vz86WCdiovNj8e+m61QG8o6G6yBrbzOXyChAlNm4StPzXZ0M3GRI8vgMx55j1zaQ
vIesJk5+XogXijfVL7uJa12PIadvPcZgsspsHLooweQoVlBzO1EJ9Sj8yLLHn7po
qFXgqSLaNkx4x+MEUBbvVEEioKoydSOX3oPoTqz34kbMgCyyN1/fksHIY7gNgpk+
2Y2fwaDJ2NnO7WdN9PgyTy88XSX93oTPDGWHJyxWZOD2ilLBM+erDw9LGHkabveN
dMRG+tRJ2/Hrwpzv1JgJrDHqY8DYc0HNgZPKmShd4VDSh5LMmoqZhZLivxSIEXpd
uraSfyo1PVVFMBDEwPcMVe4aFghcgAsMdBJQ7HFhLFvWqxMP2lEzrAuaxB6QTk32
Ivp5vCVlM4KsGNbg6c3yM6/F98tu4VnmpETTJ5a6RTI6gFb6Eph12nc1eDpIwuTQ
qX3iNOJpLvgPPTzhctGmLNgYtRvbf5FFXIiwVX9b+cdcXqvdoKXa81dUFmV68K61
Hkrf86v/sOK8wg+cEGtMuCgQZ/gqFWdPwdN0eievCUlK1oNi/fWxUvx0S72BWEyv
ruQXqkqaFLyjzRCPSkaZ8s0FR4K8sxAk82kOiXE1ZDJWynimBOLVyNjDktmefM6e
+SNLhREVpiQnOWJH8EOhnXMDzaCS93szw6wtyc8VNnOQ642a+seouq7GNFTATYtl
upMHkMpnSMNrmdnKfTovYavkXLaXOasOvEyugI+9TeQMVn6Ue90lAHnXWX19iwf6
qOsE/55Y+3gUTe4RHZhg4oHlPiNodP81c21dqikZS6ehADnkWHX+8iySigh+vsAc
5b1NBXcYDoY921bDSnjrSFTo1LNcOyJqgxvzckKy1IKFmUMeuEz1lxCcPXh9OKPw
QbVlRkfu3e4wMJF8XT6X4SMUVGxHjEnNEp/0XhBAHDKXIDjgSV3eeJgwmGm/iJL2
dniAA/bKxDnDrsemWI1SKXqKLHicOp3rxR7g3+KWLxzFVM4Toyvo+fOQVS8/u4hT
kBIoo5J7C89ImkzIcd2YEAoi00KrWpUuaJT7q3u/AUh5tzQtI5c+SgmT6oXnKazA
jcaSu/kX6v4Z2BlZ00JXRzMrGThsR8w+x0XeUpp9xve9BhwSTl29tPgbPvqkJ7XU
O+Qj2JxdAl3DFWC9Uf6YB22Ts+uhWblVnJx0yz21NjmaonvOHTT6xlsSuKi66WSP
uiiLoeDX17A0g9eXL9HaL6RQTINFwQaD1RPfzJW8PKHZK+0tg7yJ23tZ671kdd1Q
phJhffGbIiOnr0EGzZHvKvohYyFG8REBj+HtNb7lISZOvpwUcJHp85+HjmUuznnH
6Fd2+nQ5GKE8J5pV/EVQmK1D/iJ9mMs4o4nQN2qVAN3TLoGXWatrYf2dkPiLCvu8
otJ3KH9+VhLTbJyAbENFUs0zqcgYDO7IPWisovkVuJ8ADDTFsFirkx+hkkxgTTg0
Ovae4S5QQYeWyQE1WujvGtg5mFEPdWGvsO7VcYSJF4dEddGxa+4tnCxK8EjQHWTZ
wU/kuSatDmDvyGgL7Qj8WJ6GAXojWQAm2irGQJj5j2XTbXbLODWR2rjzWZ/e89XP
EnKrG4upwi/i5TSHkbnY4VHbvAwSCMRa016iCP/EKRnC2BsIZDcJLvLD4wfccWPL
+K1S0C+ZxnNkd0FLPsxm+U9fBrTPCcJsjTZCVQRi7HY10atnshiAXT/Kb1JYpqmz
jBgwxok2jogWrE2xZY3d/dA4eue9/XqkL9aKxdXlhSRKKMO34iSEOLXSvs0v4AXW
L/2wdAGEcgDU8d2u08NH1USObl16z5UQcy2uVbHNzJ2BvdNR3BflAKEfMOEqD2NM
4och9YOrdtxcHgSdP1AXBCDcLjmU4jGUfw+eLVKX5kwQU2fqGaO6qpU0yONWg2PR
B26cVHPkU/A4AZn3hH7iQdIveuFnFArKdO3sDboNAIrQXbLOdkUEHucTRpLtdzMx
QnFBNDL5wzwe5af+ExPIHtNRcoFXlEc3Bn+FQKG2IBJWQPduzowAq8dfYqFO2kki
rFhtWokiPew34cWgCKovGhJSF0QSISWhADza7AduVvT17MC1vMvwbAorP1fo1OcE
I6vK7OKtO79x/QaXg8CZMcr0sguoOOGer9D6ZAoIPa9A+TQnpXeRLHKLodMuT3s/
6V9hCKeWrTtbSNWePgV4h37N7tV6CIJD+8hHsoVZNTlndWTg4w3lTq6SXMo/Zjs0
FvAvXWkFEqmRhSrufEwHaBnEiIOJJmk5Iw7zctlo/PMxNUC8UVNVKz4VWzi0Nf7i
bq67bB1fB87UNKzLTZPTOtoDljK0ZGPyDaNddZqFn9lRQclKSmS351Rk17hIkPt6
pc7WoPM/WfwaSBWigY32B60DrdW4Fo93U7jJps/H0KNxRBfCFt8QQ9AJxSrfJc66
obpS5IQtGwp2/jQgHTLOKpNXzte1GXBpaNUTCsqNVCBMx+IFGcBwIuvstLnGDMw3
Ix64gOrLc8J5JJmS+Zbzg7v7sxfmEt37besV2ob1QhqlGnLhVHCRPUjfN9zrKeJh
rxwCyU25hg5cAatfhHXmJO9cg19lS8ttAJBqAS21mpb8GUWJlb6n3IDjHj5oD0YL
NcihU0OaI3DNXpHAVIzi8giOiLJEk2m1+iZf3ptbfosjdr87EHE/oYejop63/lnz
76wxb7sZHYfzOoscXZ0+5ruq1qd8x/BQcVWfsyxiLVnZ4ARrLBUJUhtYJbJpJi8j
Pxi2w1LQGvZd2Kv8U4sLVztrIqccMPEAWCkzzk6JUC7bSkaZe6ZgetOPok5HD2oU
fOuGG9zlfmkO1pacFI+wUdMZ9XoI9DEMp+2XTqgLrM3Mb2CvVsVxTtnPzuswQlim
pIi2iwQdzZT3pD1nhxs7WSBUzx9A+gSSyLsH8/KN4W5yK+/+0Gp/7KEJZE13FY1Q
JlVB5n6SOtwDB49hza3Ks7NeJYHCbh7owTCgPtOv22r4lYOsumbIUZpbZOJ3iCkb
MJXDk0JOEj1MtBbt2wZ/iEpxuaAphr8C4UHx5pGFgai90cXb60wDbrJycLNqWot0
LZOS64cYGleg7UtUMKCiDKOELOft8tfDVx7E2PDtU8AwXAySb/d7GLhKKkealcX3
+TYyKLwWqGitL9BoFFz0Y1Naf0LO5ZL5F9vqa8/A18YHiC/AnXEE5AwuVb9L9qzA
XyC49ygLCd6SFm0+Aj19v/o8oHlooM0JgygxhG7tzDorjniveMO4OWC/jSoujl6t
idbyPbk31diF/4moDV534DLNMX1x8d2S2DpnbG+UVkx5W0E/eBOm2HmMsQlBQ9rJ
dutEKJ2HN2SdCh/YZfkH4AbIErAGrDniTXRzqdeMg9dp0fucRkB9dX9PTXqRHZkS
Xgn+PAr3PXjULxNJdyvVmHU7Y3MvBGYoM+7AEVm7aGrdI1bg6rwk3490CmmXHe8X
wQOObbYZ4SACBc2yN7EFCXBkugeCwdxyNpYN5miIw6CWV6sSixgmnJIopbLC98GM
ML2Y4QfiMaqHfcFNHyvwsbSPAIKGlFggxAtGIKMQqDTigd+FensSlNAenjzPCw3c
8grzoAKJaRNUv8N4SB2jqvxr3Y5L5ldaPZ2xq6nPzQkmx9BS/6suhVbHz0JE+QD1
zuBLpjOF2AZ5wuvzeY5jm1t9LaBdWTNw/1cpxeEf+4TEiyivT3qYbSBs/4tL6xJr
PTKL2OUk+kaMJ0Tylv7Occngs2xFyP96uAr65b+6NeTmld2cuEaYEIrNb7syGKyC
voSDs/msXs5eY7sxv0AXNgqjpIAcTdvrxrRYMwz1fnDWTc7uXJ3Ltedw7WX0d5yc
VksG4JrAWUD1HeU1/HsTjBbGdy+2Z5VS2uUXHm/APuesvQ6i92YNApdZBse8Y3Yq
eyLVOPdjkBfxTwi8H24wy95dIWXVvi7Jfl/fW+LjQtdD+FVef1WOo8w6QpY+RYoC
wLXdOhhw3k9I9w4opLlJeriNqfpNaI4k8/19TOOhoUmqLwznL5sM2d/MIWxrDRCm
MxvWinWW8Ybqx1qewXH92qeAeeDjwjTyxwT3xhcp+WPny4vvZUwK2giDKBrUPAlQ
G9NkLE8mnPevqok188YaKnCBIV3lBt58HtRATSHB3nGHIb6cTNHBMQCOn0VjrIyn
VTiBfTCyIsIccLOoVq3TfnECwaMlypaRC/4Wsh1hu+sCTFE0SVtnuNFutvt3jqrM
AyxO5OJFdrqvxfEN0kyYV7upQjcy+0f2/BPWRVeR35LpGPao3oRh1u0H8RyCfo+0
/61u3yBMv/GvNEu0JZM5eHyBDQ7YjrfYO2Qc93hqdEfEJq1PyUhQLRhx0sa/Dr2b
wZ/lc7l6fmYyV2WtLCpdwDCyzV8uhhp4ugONCt0MNqoHKsZmbzUmu3T+FpUmNJKR
IyX+XtKqoyfxZ03EGYLbrFBhfT2i+YOnOtHQmhaSi+BT1Wm81+Yx7ADrpm8Wym6i
tkyTgGqAsjOCF9j09nJQT/3zPhJV+S6DlL1PQ0765tIaFVe+rpgdo6AhApWZ5tz+
vxhQk5ZDr9jEUiuf6ZfBsWiyUsX6ikhCRfgFYlKKHpHdicUHdcv0r5NpA1hbBcHs
F9hg/UdcslIRvtoaIDu96mq6V0WuOooy6vvE4CItq673jKRgTUWbWmqncb4tCcGQ
bSnfd8s1IdvTlhED7IAPUxSLqGjI0HSlageQ0V1A6FiOEX6alNuFsRK8TEqfMmOr
XFRqfPia1KZHUEXLo2FWhhMSLqjpLmmOiABuaoi+YmXKxAIp7OAuA2h2Xm/PdKxS
rSXjmOlUC+ejDRPhbgudNUqPwmOatnanJhXx0Dq//DiPavAYBVjX7rRQua7a6gLo
qnOhnfdBrOXftxIdm06c8r2Tja7vu+Sw73fBFF/76t8jHH6VhoGTR1ZHPF22hxaH
jYRMaMFV1Xy/LxRBDvEEvOqRv2e1ZTxZVHiuzPEkXgWTbqCLdcodwe18vsRgVZ7q
dDZ+2cRt2sBZoZJzHBWQnIXqPdJKAlvkRMZbnfknnxUAZ3zImxZKKkf19WZ3lftY
c6hw9L9wyz4u8bfBf84tPKjGfS6BIUBOnIM4WKzcOqLgCCgaTm+QSifGStqE//RD
HhfRUreNt4APACDImJEJV4+v1C/dWloZa17Pv2WIDGYN4xamgd3RHoClC9TDJbRJ
EBpMlNKm05y/m9+A+glC3wq+NDsE3PLCaXklW/09FcozUQmp8j8z8wS4HQf3Pf7S
olXpZqjgazl9lIfFiJXNGLBqAmEf7RwtpVJZhNU6uPeQe1POQuMqMxbulYqzKptp
CBIDCu+fyJqdOdnKFuqzaVC3ii2+NyOQQwelalWfkfAYBdHCF8ACby3EaVBH4V47
Bk0ypMm+c/0nC7DQqMq/vQY+OnlfkFVAOGqO4/roPHhUenlCTPp5exIxjW0IZ6kz
jXIlACxmozSyj8AdTeMWEWsDm9X4qnGEjXJnPSLU4DHFCl1HCmu/Q6E+eIlNDWZE
IeN4eClQhjRXvxjlKB9Us/li04ykL2K0XECO+8C+NKip2uekFa/9DoZ0AOQ0NH6G
+62ybjsFaYI4Jv09eYZtoQuJ3nXfY6bJ+jEPNSZ1WydzfK0whbzMXRLSy+m51Ckb
fJSrdAxSTGDRVPbOwM2UwOlpRNWVgC6kQc4/k261EkGX79aiTGOy7o/xCOFDDGjF
vbznE27/kRzP6FiY2RjJqHPujKXSV8c0VfccuhzO69Z5MCku0mkFKB6VKuvmbDY/
BCql40o6LZERFpoSI2G4WnnIH+JhbKhbL3VMT1hiaJbmd0rOwZLFBVU5FBFzGXVa
wSZM9r31MhTozHV1jtCIxYIKsVUK4aPbV6Pu25fY6DsqKbCB49PVWzKtRklRVgQS
kqFN5ZV7Dfv3CyDCOJG3rMRiU/56YQhc3a4uViVObJMMsrwazhDxuRZYs/GsoY9F
RutUz/+xuF3xKSMmx4YbXS4KXRxRUlj9fxEjECyGcEhChfgEaeuMih0xqJ1rj1Rl
FqkkxE73W/dQuhx4ng2MD8+qfklsjUPVv8pDUwRBluuWqOJpeXxOEUbOEUTPVZWq
f+O/1HGvvUgaZ9NBC2z3YJg62vJgAFsqatnxY0FhGqnLYTZ1WWgzlW0+jfgYHFCc
7ikmi3206Z3FVMponIIxG1ASX5kCNw4sKd5cv5IwIloWbdRmSW9jn8HdjZ/hk0KE
iaoDpzWzwVN6RI+stvoqcXCqVlQ6cX2AFySBRzkPUfZXoddFXl2LM7DZEKOiHroi
OJU8IweQy/yexCsGgh66ZDkSPXC1a8FqnZ6cWds2Jgs6mYgoQryrdW2IWZuGX/dS
aAa7NHBzmFRvuoUkvgP24z2QIzPVxxRWEqoxQmty+95q3QwBmxYqRPrH84ZWnjg+
kiFV7nJ6nxo21KwAu15hRcvzxMKbQVJk1E390wSapuwM3Jl10Amds0GpBYhTFFpn
ddzAZhKcWlr4xoU9bzDkeGZDsRolJhIlHzD/IQ5kv62/GOAM3wqsdfL9x7c2+9dx
Awg7ASGqLFj+XS+qcuJNTD84JonyRLCrsRV2AJfPYk+LD7s/onReMHmmYR8e5gnI
OtjVVE3kqoRtP/M6T9eyTKoTWXcgSC5sSG13uHUKoaQHCHRP6vHKjpAGWow2BFj/
blsZfXCUmNEICci2kibTuIh8BESrlBd5mX/h/ooTKLScnNIDREEpitiimrxS0zKh
d3RFZvPuTZ7p98NvGUDifuOgBJ/zevVisaBeLD7aZbuForG9cgc1uJYaFdStLNk0
n2LNyRpy2qRgsXM5rdVjBVWPGu8Y2sC20JXDrdproeEPKOXpCoVDNCwhYggW1a9l
E8yTlg8YUgjFJIZoGrTrSfvAgvrXxA2Ju9PhIvtEfexrdGINRS0AIwTPOwEC7QJU
A6Vz2OLUS4qP7UzpE796Cy/FXmLn0Htkl+yzHzXSEAFG5OpkwB7YZhh5fostza7l
aIm72RsCFZhu7V5zGMANTzryRepH7u7ArcwumhE1fbK/yGBRzh7bV16p8K+FM6BJ
ZDWkkjnh67zKxGe0tGia/qhWLOhaORSXjiPjob9TDv8884R3To/vMoC+sLsP2p4P
4vpj0RvTzJBeNPmEv3WoyQ3vFEsGPc8kGz2gdw7g/Ob2jb2xWTdIkl56iZ5QIdYc
o6oiCb7jLDLpjFRtTZKx/ZArxhi865++IXZlm2VQn0gDarE4QOZhkZCC7s2+ufCm
x4OdY38u7KLDIjwXRGqW+PCGm+inJVHYCVY8oGMRNbJWmvKsd4t7aGPPVav+DMmf
7jPTdRtEBeJ6ddAwIzBloVDC/RJLVe4TkBvYNl0TP8mmplv1ykxQ2qpD14ND6niz
/woxalJhg364Tbc5GfKIw4e2HBYMpGkNvTph+O13YSgt66auwKwnOuRfCGYQY61u
EFZzm16buvnSWop49hSTpKN6a/z+rg6POLuiTlb1WwOVc/m84lH0JQ0/L4Cd5ZVg
Ty2TwmTVC9Edxy+kyV2Z5uEyKLp5tK669K55C8UIGEUvE32U3bEwySMO641YoVj8
h0pTlRM749E9Bx10ZXW1Yy7L7JyQF+GL2NgAgjQSnlXdQntPNDE1qzWqNh1qVFcz
GflE2XXvKVooAnW96RxM85d9AZ9/9gXvc6dCqnG/rPqi+4OBnVWFf+i4d6ZebgL8
O2wImgFzVA3trcYldjFC63MuO0kbcbeozZoodTm0JB51tX248nBmK2iIUJ1Ohgvk
8ixkGSOuayxB4+tOy6Fw8z6c2LDULzwvHO1mulOHUCas9+97jF8ZSc/G4d12Vths
qnMzFFs7Oxd3NnaBOUrd2HiKxmgJyNPSkDAGtEJzmMuQe/N5DnYUlhNpjiRbnebn
32UA4r0QVKzwqRop/G5XfHx4vNRqNtrNIvV7X6kOCENmiVoo1KQHqBpbWHh2XzQS
192aYBhj6e2Oq/vNDZoM0auH86CPsAydioM3jvrwzd8yoph3de80NzIB7oWgqNWz
V/KBKUQJRD34EMF4IrSiR8rrvVjiYty9OlXY6bNn3OUmPt57pE29xMqjGR2v6Sgc
8Y/OwuhObCW7sRkib3zHL1y9uie75YSuLF19ZNbJH7q244BVtc2QwORsu6IUsj5e
PvbIYMroNRo4R9GyETmNAASIRDXXCBnlh9lH9a2LqBFkTVaiR6bJkb4ZqwY/7JxM
jnmqEK+x9aiVfLzDDq//wVbNPvvRe6y638SycoQdzFB3wyVuUtvAylzaJua6BKY5
FgKgQNtGIjnqiiQ0g4yyAktpTZJPQpnfEgtc15WMnKkhdbcIxDBXnHh0uSBMHwW3
4yy9RnNSRaolsTVgIPh9XkYCnsRc2UU38XblrC7cFlCpnrIdy0Ai25Oa+uoTY5Nw
Djp1ss6ndnE08sSX00FH0Y6ygD4TzmxVYeO0V1sR+fR9vBaeh6MoTCsoaU1h1NVT
cM39IH+Uj9GnA1DVsQo92bCOwTvyNzxdXFC0Q6OkiLcPFx7DtxuEjuwuzvFfX3Ps
5P3b2Kp+9yYKwAH1mzjhaNo1opIWCKtjx7eHxXyuZ7PwZ50FNuV0gmJQUiyO/90p
r5ZQKA3GE694r2T2ur89NVXqSLmtPZ4UX24dSOFnyAx3e/v5T3g7OL9K4X6yxkhP
F2ptz+FJXzep+mqs6upGHxEjk5/a86JcfiVr0r083fhIA7DmeYcqZ3SrYp3lq4OY
TCm+jocFHqgs12jiQYnqD5qKXAdQcSmwA198f8SgSvCmf9Y5vqfKwn4uKm8yko02
ozx9VyMAtz6Vtoi2YqJC+2Wb9FUHkfBexoNTGjqtqStiiUsrPP+o90e0vc5wPweZ
j1mqZYRcDFuhS3TLNFzRUwU8JotUvncrHeoanhmGH8/AX66MQChk5qQuJARzpWD+
3xk5omiBNCex3aYvgliI2VC0kdbEEHBrKEmKJyjUfMvmFlJIYY9P4od44+H6JBJH
+OLRI7SRlr/VHfZv2arPu0Sj2nyIU/eyA1x8LhsmX3XvxFXzg+Sdy+j44ZXWkmvP
hRDFgW/isqaHuoWzq6kRPflnc6oZ9iw4SVK9pP6BdUgBq6C26BHpSX2VRP8zs9a4
HLq868km2eorgGmkSDhrvn5K5jbAyN1HkNdypTXbPMvKfOsso5Z1mitZT7/styo8
nGJJ1bSe3UtwitcpZp47M1WKHvL9Goqpsha6NGwZphR9yefeMBtpPt8cfRrm3Ix5
KXUR6fL9vNz/SnftzgicGbtKI5DG+S+rnop2sNBtWe3fjYFjj9G9M/qfBKVOzVUA
ABMS4nqEXJmY9OkzNOTCwHk/8qfBK++hnli9pL6+M8fnULdaS41FRZdVDdg7HkaT
Z6R7VGZR4Fbumu3SUKXx5JUXJ2aEzAtl8fnv0pxzW3gUPIDPGTPKEuniMUU28ZgW
7bp5AHyoduWMFFsWAIlrG8SMjU7/iqAGTpXvnhJmW90f5WseOt3nw9tLGYE+w4RC
UkpU03KT7+nfxW97B6gWv3B/P+nYSHMlQ4Glz4p8baDf6ypBfDPNE3jn4KTly5q1
vC28Y+4Hnc3PHdQNgGKsgJe1vY0D0hCLjnNEunXeSm0OShgA5OW7HwfOyumEn8ui
vX8+AzcYn2RknO/NK6aR3zHqDpjJD0qYfoSgA2dhyCehID4bi++IZEJVEm0caDVw
3fE2oovWOEqaHbVeJ/m22J9/SZQCD7s6V6/C3okOaczUAFZJDnsH9Bcu6n0dHY3u
cDpZvLLjXo0lYnUyyQOffKcW6Yzv4i20UVHMlPh1FsXmiOi4FVfil8FnnLWUVTiQ
siAbCEovN8AjRnQX4R2qaASE7/bZZBfWqrTD3KdJwD2a6knYKdKSW5mRC4c95KCT
16bE0s8JM0PLN03wBQWr68WGUlThq5d1EXe1FE8Mg0wyCkvUeDtCHU+eJ9BRaMlc
2XzPaiHTlJfVgr/duOyo+21HWT3OkboGtWpK93YIwlW8tNqel7HWPt9P+V6zSvyk
cyK3YRW2EAwvajso6YU1bz/GUxSM5cIWTyiA9Ismzi1qIT6pXMfBWgq1iEwzXpZI
K+QvXsJOpBLW41eX9l4hTp/Gl7Jdu6l4wOh5dmOmm52tMkafGNFPKwjoHYHIQwnq
HvMn95GudCzCQhAkqOZc1Rrzi4blkc31sMDW30KcMSNV9FeegKzpIw8bzg/gUWEs
UrqDMqme60mkirt6Ph379o9wtNyklz1jW2Cb+u62v7RCOKime7KCMHP0x7TMGBK5
8Ka52pUtis2Eiv5d6KVORSd31Wl3l//M7NGvFemGzGd0ur7cByHRi/0d5wlwbNQm
Z9ZzOKr0R1jE6WaGXvDXg8xR6yH8d07s1m50qus6vhbJX8FL9KeKyBVqgnBKhFdi
tI4GW4ysTkuHJAMrE3B61vCmjLmUlEncFaWn7USmjgIn9l2GskUSkfr9B7aMmo1X
+QyxCPF2UIyeK1AnovBXeEgzkZJ68xgiLdb14rp0u3MhlEBgSZfSDqajpgjZ6vUR
QiPtWxRZttEOu6+x/5feGbijSiD7HfiON2ooOrP85fi0+vHH4WiNdXuYL5h/+Thh
ro6RoQByeyuQ5HmPSE9pcEY7iXYj1GYl+tkXwkUBC7ofRpd98XQwWHMAq0uGSmmQ
o+akxN6Nd9G9YGytOUt0p4I9R9SzTgM4PRM4zN2nz0IomqEhtD/y/KfPx+ZklYSJ
G12pjyQnNURnwGRLGaj56nHTIDxMHWM2J6V0lD48zKIg+HduqhYDzv5mnJt7OUmp
HvdsVGY26H3XcIaO2LL/H22rSh88AIhBzYJTEY/o86WUI7efCXx8mTBoYYYPGBKz
bEETGxhh+o/tjecsgIJul0H/GHXBUhQzdFpUcULLWzhKcN4tFFaYK8NiIJVDtXHu
YkL6uwg8CpIOJkzBj46yy90Lhk3nclvadsUDWG3xMLoFwOU/7fU6aMHNmL6l8wkW
6HfWLHtbJ+47mplxyJ8HV9ePfCWfh0mwquta726gNKe7NUgz5c87xTs+TCG2zhJn
W8kKYYmhZ7WDlKzIAIfRCT5vajTSBGgYdEZXR8Fd6jl3Idyz+5Wvrow0CcSbBUj1
LlCKb+AMQb4yzEhGvAX7DyVp+U2tE1AM0I/YcPx1xD+OxA8YkogNhk0ijrhpqV6G
zIyJQBiE0IdshvhsdNpQnK9VKM99yTDjyLBYEITH4lavPHwQsctq/imOhVCLp11v
bCtq/KY4sPEP0QO6LSuqCtdt+NyMvvxdWZMbC9BlO30e5WMLRyjfc3oI1JcnUVPX
njBSFN74TgcUAEBNzOnawvmfQOC0yUcyKYSwQ9EV1eDZma30SwwfZ8AMr8FWD6M+
i103AYAot7rHNIYoUiTQsSjULpkYcZnU5dmMbPmn0HP8zPzLZH+XJjvyxN8L+SAK
LtYfi1h7GPFZMPKd9g4n4AzZ/v5pCjsRB17y8RXBoFA3w4wfAsrdLvNfv/0CQqAZ
LPi74uommVjWhEDqklv/7iNH1EYSr4RLcwqf2xkGhq/+iywiE1nVbWynOKgLDeYF
SK5mXPRxUJl9q4YHwJ7ClIZx9T9MyrloILiaQBF+25BDbPF5NsLVHr9pIX6/Lo9S
hEireJcyXtnwySI1FKwIgOQxj88/+/RmIdZSNukss3eJXrHHvjBhePmSaRnaDcI6
j6Q2URf/Chm9cz+ZS+Cmp2568yZpxk/D9OgODMAnbBkc8Pkknloy6mdmSjkEY9q5
2viX0SbafQBHW8MCImEGw6zkpb0gIhcURf60UavYsj85fOOD+oXwOBNyfiu6HePA
k2r5i9aBY/Exd/ghIxvydcCrPQdkRL+DZYb1lNLUpTACxu/4zo6a6/GEG9hXJiPW
pwB1v3NDRL8daLLSBLL3Ze9aiqP4V3qLDiYOhsGESMIWfV4q9kwz13dYNfrZeBg0
bjbfO8SpPm2WFW8Qm4b4s3+PDhL2bMj+3/G20GqrD44k90DpDFJideQsmd+GhLwS
2L6r6gI4XtzSOt2M7grwc8AV2R5Pyfz6Csnxg3mB/Nn5yNSkk7sf/a12abLtwKDI
FGL4z80F83j/vhwDt7I8O5j7S+tDXhW8LLdHToGRt6Qn30/QR2EPdCJ4uCBuFi+2
zJpGLKAsehEKK+LEwC4Kg5STXN0C6y8lQD+9KR57ANJg1arTQ5PSNWomwUXEC4Wf
zw5SnK7I6VMBlINVVP9fvhbBZzgsHOCp+zZ/yV6WCic/wg+GFMtNLf5fTwxPa6g+
ow5fktlQsklmj3tUuoPZno9AH8YQx+iLaoYo6TIVThyTa/u9a2yTm6nOwNEwJtuq
I78b0g8PQeV9r5sbmkmuCgjlj5ijgXGsb9Oytn+YTQB4NzhfPPDNIb6zGLCyJ4pv
V4tw8ZEiXsvAEiDxkp+1tM1TZHz9cNBALyuB1sjch2mHujZAAIITsoy3MTUodO8C
4W0zCuqfiLhilXwNOsEaFozSW6khGJPL7KVIjcNYgal/O17ANWikRxV/cdVKWAK4
noIjITSJiaZ6gl+Tky8wzoMDEsjWOpeJ7K5Uqvc2ZhnkSxYgmlIZOD6k1lbxj7YS
6se3UJWeEocfO7c6x9F0hMZq8ipJMJzZ1HARS9JQJaOQTfyklrVYNl4NiHWOMZnw
MfAdXItlDCsmuil/G7nSzup/sKyZQN+L/DoPiFCj647kJuMGuXakk40uSYXi9Udw
cZaD8n5+mxdD9fVeupf60GnnmHS6VIAvwxH/Gk/jHdrefWQv8NRAS4Xira9U6/0j
vvT/e43yJu+gRXB+2IsUlRgmU22AdlPUNFRZGYvG8OPTIJKV86gAS7BoiEsUb9xn
etTj/8YoffYVPo7ehgxlei9oopKGntl8UktR2m0kQGweT7uASqEI7osXBwFeJOTt
cvAbl77LTEA2VYJI16fWiH1OwmEVVV0vABavyEHmfdq163ycyG80O4MbHBjQu+D+
Mgia6U72jQmfmicYXZJy6Xqg7lQkkhnfpleS7GqVc13c9KHHulwYfO6NR50jjaxV
nPjMTdmBSIQWR6yvXrIDe4ex0fUfpTAdI4lNzFeNwZlRTIzt2mT1ADPt3M9mEHnx
9lWCHx5wU14vCx3Jg6naKxTyg96q9QpKj63VrPBAFbTd2RQ23t/EKgm18VkK/JIh
dIN6nspsPb8Mk7MBTxnB76WGFLGptaERAKaLxwWiw5yXH93v/zCr3iC6JE+0LDXR
xxz53mXxIkOM3P2tmm6wTTnve17lmRw+rcn+ksUti42r0xVlkN+qP3FqC1DKO6qs
dp51+JzR45QhoukvGHtLXYeK6aeH4uJpaTetjs2u2tyPmSehkiZ1O7xP24ifc9Uq
/KcSa3kzzfIYVkXvAzDlZhMp6Rd6dYf0EXpqnY2bbVdBW5CNZfRKibaZoKPDWNfv
AdKC+ZvkU/dI+aRgmjLiTV8JJ5zekmgVehAkIqDCSmrnpaJajS2fpnDR3d17gZWv
yUooOKIFGwp+91VBWtP13ZTtG+0KxcPbDpxLxg55NAiMi/R3Ab7jfzh7vqj7rLbV
5lIheiWjcFwsYxC2Znz08zNPqGUql7jzT2rWsl3nclA6u5RmRSQpNi2lgLiet/ez
aiHO4g5eyhmWw2abEa3kdM99tA9dSKtyT4EtFc7+MN/or1njAA/yyDQiKx96ve7J
jWQ66JPSe5IYLTj/ekLbd9uFydl9bW3etSNc8RJukgdwydKhp6jss2t7VLgr/oYn
hADgIIzXP0BPORsyEymJmuWuY4mwf6aiF9GXNXO6WVW3DWQMtnv4MVMau5xMGO4q
83cuHjPpvgjnFlaC1xIZyIIlL30m3caFQQMpZFWHZUMwzCGQrLrPdHJ1i6Kqjt06
RCalU9nWSqNbksU4KWglFl5NmdZAJLSYIF8Qo9kFq6+9wbfT6oPEA997G92QCmeC
lQ+lxD/aJFVXazbJpIQTj/zIGqnL0CMaw3Kz9aeCPKde3SnHPlAaGJg8Sk52DpmB
Ts5OOcRX4lSPzythTASeEZB9Q//tCMWNevDWwRWw+nrLxpo91cjBKF31AI0qkzy5
FS5cauTLCW7G4j654LcPL9TqukHnotRIu4UQrpnMXFGYtXnCOP5YBWeIPUWtPe/u
xG5qT8B+pM6XosyFFwGq95hbIcKBe8spsXQ0HqLK/haT3LwnuRhPM9dLg2mtibyB
86oYn0WSluM0CYOnD3Xhv6gQwY7RVny0pAoHgteME43CgHWO0fpbFC4X13c0FY8q
EYYt2wSrSLoPpoUXzGXZgBCGL8YWyJK0o9VdZKZJNqIvmIIaD6Jzer1Qlod/YmRX
lENcUMcMkjg2hmvlbilxn3Y4rDVh0xTIhpG4AkzV6uan4XUz0ejUziVPjk9u+v8V
P07DcqyWGnfUr4434kVUeJzkOfuWgwEnMDZU25EdzRuqmtrjK4dFZaAI6RaeonNK
m6oxUhJkxO54q1H4zL8syy7W6HLFI/ZXfWbGMEIq34n+olyyvfuZJHDhjGvgJfRI
s2IreCLab9EaV2wxmySpobRRGpSE9XtXYODxws8CfHU+6XWhoLnRL3qxxu2bTxLh
CLd55phcIr9sVboSkKXFTHd6I17YZBjksB5kOWQA1VGFoIectHUqP+OiGhc4v7nD
F9Ay8Wlzm5W3LeRypo6NdFOsTWQAM/eiIfM9HiTYK2wQkMvejPS/IuFyNf/AfC90
InMfWDgAZmi82atAcSt3VGWvlIcfy0QaTlhJIuds7YUzgTq+FV2pQkGvXvOEg6e6
1SnHUc4g4f6t3YGg/h1FxNw/hFTnxjw19W2DcJ0n0IDbt42MOZ/d/fPXlUdcvKs+
PnK7dc9b+aWPg94a0o0b0Vno+7HO4Qe4Swcs9skz2wg0fUZasTWhxLUqISacxAXT
4rpidp/uoc/5UcgLJ1FcM3lQ3YVwMT7OhEbCXqyz3hG6at/hcPLBXKnG5KESxqQ3
0PCZ5jBwQjfTQ5NEkZNXdFPeCoqiYK1NnIjv8cAfJbHhKaOjHVEFBk4FZKZgjr6N
NepTuwPW93T5rho6wPDgtgj67Cr/ZX9B8mIlY9xGbz0T2WvjI6rHUBiyfZ9rfotn
sF5I+tXC/iHIiG7xFzg88kKqlG1lKhV2Fm1ZNQcy9WfuYCU7VSfrBph5I34hB6gz
eQjHR2TPTV8cJ7nizpz3IvuHL6hhuc2y7zoWjIwnyIFygkaxhg56p0RL9emZ0AvM
JaGILvLyw+knOsmiTBMzpusnrrPwViWAmfWVUIs3a3y8IZ7sy/QmCayaiWdZama9
AJx2TukLAmnHV6eTAhHsMKyRIgBS6ccZgQhP6+ZNkO+nxWD9uBgG6qYeYWhesUC6
NfvutNa0XhD+zSWf/NOdfraEeX5JeRC+iwPx3FN5tHO4z8a7S+JFVXkSDwVvqORQ
cyuvRCUKfRlMdZsysvpBlbKOqSS98hFNE2NZVye/tY1nLBrCiPf+OYIqxYez2Cqu
y0Dlnb8WBXGp5SC39UDAFYiETGrAVBVwZ7HbIEYmxJBx8LwJjk1RmrTOq1Ml1M0v
6TYhNSTUkBne8duPV1MHy0BLBBJ65CtaFgiD/wVThgqCYVG+aUSUOhPBqO10M0Ge
hMj7Ega65S179M0ECZId7ECfMHypcfHh1vkE1Bu/kXH01baL87nh7gmos8pn7hVw
qpnYVdJvFdoD8IH7rRulqmzN8exgwCgY+S0VJ9BvX0+5T8NgpVYXrNUn3BiaY5dB
BP6wOaSDm+vixmdLTvzlIkII1nR/FWbLSpTIdRpE7DAQ3YI+5kwEw/npNTVz/CCf
/OVi1GCTd6VuJHRYh2VzUmEU2ubT6SLKruzURX5j1en/VKmsTqcR7codrb7+adOn
9+Z3Zk52UGpsY6m12PIOiwGLdfY0g1mLzWgos5wrSNkcdCOjj/H8yxbrQ0pEizlV
Ub1ENAz087WIgW+fs92+4VWMtUAnww+3PU7POYOdpT9irdahu9DcVLshDA9PwO2d
XBBs3/JQGB0015XoxZVfyCtBaJBa7Iep6O8HzJ/8RycH6G/HIdMAq3cLtYzv1xsY
Itp35ibQespOTe2I+2iHyTWNemtMQumlw4/YikXXjalsKRN6UDK79oAIdVpxp77z
DP26a/CBoBECZ+MH4y08YEwHV0MUV6evpKdeZlsdmrA3ShXOZ8+9TDm0I4Fe32Zw
EdN6ElR1jUr1t5xsK1k7CVSWNWRlGo+7RQE1N1l0d15ifRePLeG+cSpagw9aBnbr
mvucxk43CT1rbhQz1s3XVHb0o8Q7erj2D1EnjSOU9eEF35iNu0YqspKydXStc3q1
odbyrVMd7ZjZwNtsSVDBcNCJnq8Mi0znio/NVzeicL/P276fQ4+lZbYDcYuJ1Aoj
zLE5kxGtYO2ZFKua1u1L/3iQbzX6s+qc9K2aek1O5Yb9ZLrp4vjdrniW8phVU6ku
lALR57mL2kW+0S52738aGCpmhfQ4MDxOjpdZwqJGjMs8nB6TWNc4G9F9EYwRSzid
jEYv6jO0yv5MLX5I21wSMCb1WFGbY+A7JTMXvLJEC5X/dFdMnKycBxi5DlnRcuK2
WMXvm18KikuwfkP3++il54kJ1khVCob8cZAibMacGfTbk9zfoLrqkm4pZcD5j/db
tf1ycMlTmqCQ0V91bRi/fFG/vNqFQOoDziHfKYNVdhTfPmxrO6FlD1Ku2zBkf8uU
sjLn8uwJwdcHAJr7zN8A2kcU0m7xMFHa72lgwopgp89l0Cvn96VOKbOMGEaQCCJT
r6sg3o77YJBmot02FaPbdZwVYi8K9/leqkQYhGPCcv0KxGC3UBJOgMRjejNIe0Ms
DRCHgoWqEaAlyKk0p7KhfxZq1mCX2f/wBrqchlcEmYW5+9/rCbaj94yjjHVWc3B5
My3wc5BCWQ9jQh6oGQ0LH1T/h1FCGD3HXqTg19TBfKjMyP13jAFMXfnP4vxYMjBa
KYulsUZhP+dtBJuQUKbs+1fZ1AbufhJ19QO7ExM0mYWRnp79JRlcI4TttH9od+Iy
ArarS+Cwk12jvOj7IerYbh7LWgU9CTaY/GVtQC3sLHcJSS4mmrgrz8zlwahdTo3u
aA+Xcxpk8FovaThnR0XGtSmkL+yyq9VqTypqrDH+fq92DNEtSqlb3o5GlsAWd36G
zkLhGkzUXkhTcbdyOTu/SNWCm/JbwD2MsHCmNbuidrmvtrXFSGvJq+i+3nLEKMUb
B9/s00kDDfIGWoLZlcH656W9/vz9RhAjcJKVBDweO9PWVdjo/7X1a1Rr0LXqm60/
ldCCWxEO61I8IE2hkqRG+UBumFXi0Ar05DYTYhgOPi57nLlOiINx40RAm6AVLNfE
ZUvW/rzwpcu9m/bpoeXslLH0YrNAyFwDXL2t8q2HTcc+EGfxZ6QHtW+NagP8Ep/g
lPM+iBf+SP3kRP6nLlWjHaFcgavwtGKNSTWinqkOx6rGZntYhlOpwNe55kpEZ1kN
44I/Zyi+eTmatIQoXbsONP5KH2Vh0N/PrW7VjqgZUVx/s8HIBCZlSPOTV7YUW7Av
/uOJSR/2xbrMYRuMEcOKxR5YujFbsQFAh0W7aq1XtX36thM8UNOCtKTs7PheeKeN
7BDres9M9/+9xNXGTIGX7X/0fzzwWCScdQHa2FGGoURALcj+FYD8VPNC8I84Frs7
o/pqft85vE2UQbzbDw16xK1DiL+0ENtuGTiFlqYD3MGyXoQMYEVKzUjb829n4MpF
XnyGl4fKhapubdioCzQBnhJMyQ4/tABXflBznzxfvoWdVulqOQXfBZ9cblE8ssL7
/5dg4U2/cRbpMjuYmEXAooDXPK+rfc7kYJupBjQifQBuVgb7T1vrVwRc82bRBkDu
9V4Jr/bfXZhEc580jrfZ71JcdAuxZo33MSYli0NVyonjWNzfY3rTnTQy5zZIHy8m
ib64HV6fBOj3rqLPiZV5HS5xLC9loESYzUE4kAkS0qt05LkSRNxUN4u3KRespx1B
2txWMN4w0E3tGkG4yRSCvfk6WsMSPoCecAWXy1uQ9TrdYcDobbuoL4So0Y74oOxY
xIB/YzwrAn87IymM2F29dNOQZoabT5DEZcbt2FO+IedphNv309TBEbSnX9sJ9hTP
PLMyOHt/l2l/2+Z0fCU5zJG2Tol70urjPZq0YHWxc4osWD/mw5N/+85ZU2vxBXze
NpYr9Ri7hqfcd8pX6chlgQlwMzf8+xAuZEq5/k2xOV0IHhcx2bs21h4Wj2eBxrL9
fbYwdIDK3tcksVYaY+BfXaZI76ztc73G4PvREqc5Ul1zc/CK5XtPAvRb6r8Nw5BH
VoLUBBbSUmDFG+6a1Q/nsoJi4z44eukc6pRYjlPbak+ZVPwBhuAPXrsKiSfqeMPh
XHju1cC2CJBzEbkbX5o3FxZrgP8aS7Ixf0SJo+mbAGiRa3KuHXzzjOBVgo6y3cWN
S1nE1DEdije8RNPvihfdDDOdh6nsn5AQHtY5PrtRg5XXPRR8uXrb79MyWwhH2/6V
1bN8mxH4QWFzIfkiFzyPy9zaKxIc664eEzPo1oYaLqFcg2RpaeggydYaZ9adr4BZ
X90JRWJsksCEhP3Ot8+Fv5e0w6Lz5dA4OPgjdk71sDx+NCpjUuD7Ul80ue/WVgDO
EtHy8BoTQemtKqXCj0ZDSOrXyTQEkhi99pzsCtYT/NymWi2GF2AqgRsvKMLa4Iqg
Wp2l9aokC0L51k/RSqddO4cPMjgyuxqtsFqNh9u9UQxuYkO9A8gTcSIRXXRH8t81
oKxi1oyXLuwcmTE0DRiH9yg2zkq6QvBBmZe4FeBoJchfZIEM/IM65DuGrKK4oGXl
sg6mGz+iDNFSGlfYLLx5zRb8nY3CErWSgNQudaJbbqYVSYePJC1DILD7EL+JUxkE
EPIAuLtyNa9+FuY74yFFR5bt5jgtWS50Bt6PX1vxA+6CDN2HT4Bi3rf3eDcGt3gX
u596MNv3Z0I9lYwhm0rImbQfPumfMsKuD+KR6LOgvk5Fw6OXBip4Q1B1DlbQZ2mq
kl2x94ujrTppudxL/MUMPnwE8gVxVTnbuesXTpj5f6K7BuvJtaYxHDU62Bn+RxDS
88l1++7uxA9TD6p6OiqtA3B5eTVTJAgUJ8gMTmc0/hERsZaoyXDulfe15VkHem47
9wVNvaL5mQpy90wGhRiVpWs8ez+O7XWthPA1pnT0Bhe+PdVuARS10EgtgnXcz3yz
tV2IPmdiVuuq+x2hQPIwajrZDjZni1SOFSRjE2n8yHc6HYiIQPfT6FErmeRLhhX9
5uELUrE8WqdeegVcqZgvP0p6ifMtixeyCuaW4riPwNrIyzRR4qvHadAUhhQNG5eX
1o2o2xKlK4gk5XQyEzCJqWPr0qniw9RXekzffH8X+cuy8Z904+jZw2CYfwnOfsNh
5g/kjm6uKX9UbCL/gToeJyGOTVUv5MBIUiPSoRelmz80KuMoCAfkf4c9mPQuXkY+
RRdPFp40kjfBawGzwyWOS6aLTBJKthLZKnYK3tNWn3fDfu0zihoSmd0iLQ7JF8SV
WMkwFgAKMlbXxiHQFBvCAeR/q0P+eCIxaLv6fuvLp5W/FtqWTNF1whT1Q/B67YnU
g01zSoxiu4xLIIG5edEEsq7OwmDfbYzbwL6dI8BtLNGQAEUiB6ccpDEPgNW3iWv8
HPgx7CiW7ZECek6tq/YRXcSzoLbGn/nO/WasojuMVIVRZbVZiugt1p/ZjLJetVs1
/mF2GzJrxI+jLvWmAXSgbqXEooVtWw8svxZe9Bv1npWCPsarUvlt+ECNBI3ATHyO
IbO0Lf4Gl1kJKOt9tVtl3fYzOs6Qml6eDc7HYK02hP+e4uyyssCbYd7XZ7jb29oh
JNkQJMCh9LU0HYYiOuYInqriUzTg0hyy4oipOBD/waEOVRjRefBZqFpNauc+Z6bZ
mxuNiXJt27mZok9tpc0wSpfsrGT3xH3Z9DOjWSdB3yqCKCAejX0plcsFV0/Kd5Ji
8Aus5HzVeXmNJJ/o4A61ryZhhPZHex4rCA96M7yDa9TBuj9jhnnJ5dTEjwP3ncNd
QzbTug8RWsRgCCMu7MVjHSdO9urZWMf1ZVPd/ppNzKraKuBWFRdgd3vknBU2nrLi
fYTbcwodZHGtDbcyuDD+98EUB3B0hcSv7KTExEbx+Ij3uVzMkQTU+lCq6U9u+Z8M
mwia45hpwFpWX/X2boDCS1KT8/s8ErzJiBObCQss5eXbOmv+DYghIGgNcuZ+G5Yy
g2V4He/oUyq2Wf2rusCPlUCC2wfYjQ3Ra2oCuuSnMdynVELkkWL/PXhkguEJ6d7m
ZM0T+zdiLsove9si43a4xYpDN/X1VrPZfZtF4FsbC06wpmL/6GZf3bL6goJ5ZELf
8ZUfkixy3rVHRouAtGkSmHLhy5BKmZpv79vuMMGXEygKQBC0nxpXkRdzroBSGxZJ
5agiF7luJQ5sAScZILdc2bPvf/vSm5r0rmaFseBoFIFnDhlo7cbi9uanRFh+Z9th
+zFGcuvMKfgkbQtDKlZeXU3r+GGpWuQ4t0pUJZ4u6iyVyuhp6H5y2CwEEKfepv3C
/123dgWMWatBX6eNxM8/47TQw5N2Fw5n5B3MzHjJNLxsiwTzFN7n4eRHNgROlGGR
UjgeMpSwhkS1tKwk8jiQyNM2nMfxYmoB+6o0VznDXrksDcgDnmxIEzCQ9AO9jzVT
UVOsYchcPpAPuAeWJMo7IAsp573wTSsjx7q1UJh7JUZ8oBunO8q+4SIkM1g2SSGC
ukr8VNbIp591Jzroagq8msF1T/2bJBYAybGJPKdSw67TGrFSXHqY2NshVGJxwuU4
qxXPU71Hmk1M+Dgi0V9iguHTO7RmwVkc49pCS7c6WffZelyg+7bRikOU1Dj4g7bI
22NsKlwfB/2g2lBaGb4euhFWZrADJxpCiI+jzmIRUM831YiPYdBwr3XYfpA/4As6
gZZ961B8zFpzJnhag8eOWhYmEKCO9qllxS5BI1mf9XmSFwVd4ilL489Q1dJjwnRn
u1sO3Wmn3KVZ/D2DEUdiSDvHdbLAkP0iv+BTR1ls9qxUQr0JnSK8eCV9OIK7kjsn
+dq6xyYM2xdVxDPkw4N1gloELHbvKiuJ3atSLbJUJoylnshCafhz+Hjcn3tydZaB
y1DWul8NW6ICerXp8vvRGZ+hzxb5A7BwITY4uIAk/VVOXcGBv9AIllJTAePqCmUD
STa7bf1d7meChy5knalpl6GfXR0IROruhH9HefpI3bccQ6jG4sRFwFx+2cf2Qpuu
V9CNFopquej4ohwkFBvE6lhZVgNWYiosVTvS+mR84qILQxsIxQabADwIns9MJMdN
X75hVIa8kzsOIbUuCGN9EwwCJXiTvKVnqkK1ewOksvRkJaX0tmUBTkRFhnZDP+/u
eIc9FyO5t3fpzT+8mdfC0cPXm91fPbEgk7tQnnbyq9ZRfRXjKy1iGcvRL3zhoLo2
DyA8q58Y5Iz7oPkNN1dTqhnSkuu9ze2NoWo90AhijcL1j8rq7vNES144HuhPAAcE
DBuIDVHpo/AnMCP3oZ8PasYS9zPk/8sJ8aiUttplx7XR1R3CMzvN9894ZNbigMgj
awFDx1o5EGAR8cUtYSRZKf59BzIhXoBdCUI0Chjg/zx+JPdosf3mlZK9pyGnI6rQ
H1XvLbqzlcc2DHIzvXn6FRkoKCROM/rjZ2lAQcgnriihpUgEwhA+3HtVNuQ8BAX1
4ilUarrcBZYS/8XyKG5YCOrTW5McLFCdOyWWIhiVnHmA1QCwL40pzWCWo+wZq6b2
hrjxKsGzONXkuF58sCPQOZpF0Z9OzJW6gEBkC1vtF7p9csEV+XoxpAVg2N4TZZNN
oiAxNshsuulhkUjoHlZJ1ULdcpOlOozIdjAZObXskLIRon/NMj0/HOyMYr1GX4ga
MvGH5QSKVPRbfMtmylgW+8ASuc0OswtFDcA5GfRof6Tnqj1oCbkJYpSh/03arBM3
ivsiHAFcqYTpv+g0wwBHOPMazaP6lFWYFuWX8QZ86aIcxxu2o/pCsHJgAy88Kh2k
NKvLoEsnPnDSdQ3RFd5mb8SmCMCJcDkCBrYjf+Xo2dEOu2FzkRIxsjXmW9pMaJor
19/Dbi5rfskA2gj7tEgWyYN5OArti+o0Cxz6sfAOC+4yAQ7QEt5z/ybJ5YBeTfMd
MH73I+cGlp10r2ESUZlfNf7ztsQJApynm1H1ghirZJ1Wz5v13tXHFaoSkraQqOQr
5MI99rJPez7tkMQKF3OS8L93ypTukol2xgf4lVFmgfSuFXvVH6KkF0O4R1tttKX8
XVq/DY9G+9uEFgQoeUoj/Y31nM2f5NC9tKHvqZpbUES1leckfPP7C1EgH5jqiWQd
z5U/FV2dkRoMZrop8F3IDkIMQ/1HgD1iONUFGnPBet+iIMhRG5iGeJzuuBfKP0tK
GUMGIYyoGGKY0gC3cyYs6DYNF8SRlgJrZEL89Vnna6Jokr2whuDvBP662O7hvRgL
De3WydveXp8Mi9LWjd5dtSQuzXz3AEpMG2NqWNOC98BBWWYyco/OAOv4ggWN1hHW
y1N+IcF39useKu8Cgbzb9adYLmWhvzDLBh63F0fYfsCznsWkmTbOyajcDRCMS8/a
MBo/fgvi/tSQBUrFW1ok6mWLTo+b36Jm48h9mS1uYts0GNCk08LVSdBqihZTxyet
HmPcJFyedP2suNC3mEiijavhdUtKAFBkzldnhK3EhKNcks6jHHJKDxnA1C3VCq2K
rMDIJWhvFjv9ktqa7M5iy/Mwq1+M19a0J8eXZezFNmytrc7JIQsvju0pILkx2LRD
IFV0AFXm16BhUkD06cTvdIt8/f1FiLjgMMsIXWEqUlcS/tLdWRPLfoZSlXZuxQ28
s3VcFK84Ri2udsXuY9pVxhnH+99KKY3BAjBuheoyeVqp3U7n+4zEixweYf/OyV0U
QflAPT5JsfpwMAndlceHiZkg9ACgZZ7sTBSO/Z8lqc09C/KoScE2i4gf4XoRlvNH
dT6yT2j5IYEYO1Ic5MUHvyaK+kVaINEWBqGUNY2HXsxBDe12j/mdaOTuPk3QLEu/
hr1wv/tXqjrsN9xxr11LFt29hddrGoI8yBvbG61BYLPMr6yAjEQdA7wEINiI82td
hgHHQpxXBQO7v1OV5YHhT+csSmQ+Sw8+oaRItChfn7ZH43ERnCbSgTVvwpA6pZB9
Hl/AJhyvMzGmsXQ3rHc44+t5JvdoXS8SzAuhmYN82JD331t/hPaH+11jWDemQOrK
IQDhfV7kaZznXamCBogZcMn1IQ5yU6FCFKoikez4U8uMwIpjU33kgju1aF3AO9cB
izGKoovhdHr6hjpJdIvdb3uKyruEdCWr2fe9TP7NNW6QfMwc8/NHvCrUdVdY7Fa7
n93fPMV80ZLJvp/FJgg6gCwcmXpy20urEpw95hzYfNgLzWdSaMFeoppen5z8hbyw
GHUQ6AtWcHcXBBtQ13VjhA3MAsxMom/wU2ulutDlEAnsotPgy2/Bv1VNistl/p7r
d8GPs4CLvX9kTkMJih+rCkIp9XYrn78Pbqkf7ncUIlPakjASTxKt/kFUJqsAlqJI
jKdnq8YGw3x95m7zZQQwN6R73q3qjQb2vPmzmF0pNPivcAPbuRTNlwvWraOriHAJ
UafKe5tVLTbKUBSPg2D/1n3TYJdfw/920/YLfslB455GQI+GmZQQSp4nnKyGE4Cs
l+avKhz7tArN/+/JFqI80cu6+fJ5eA6oJUoDVtYUg90zooTIlcY2t4mUHPnwFxKe
0sPkLp6t3QkHKyQeCvCQ4wZtPme1oAczNxnETWL/757mY/7Kds3tpF7yYWQWW0qO
0iuNfIOmZKqu31OYJ+Y5mxN5jxcMGf0Pn0UJVXmM2W5rANftZ9cmf1tO6i9Asc+C
abAYTGRV/yLF+Z+lknc9G7LhWFyKqHYVemBB+LQkmRfhB5x+I3xjKfguo9C/mnW+
LTcNcbzvjfjqRTbkZA+PjSQlSoD40AdYZBdEqQfuqb1vRqu+Yia2bRvlTsEXCAg8
cd7/CenK8KX/etA54Wp9yZtTtTDW14WQz5TfmN96dwXWfAKPgKb19j/6blsiOhvg
uBFoVkjaN0+REwHsYaE9gYQ4dCGFE/fSYpiCc713QMSj1awnY2Y20e2Swp1Jrt6c
FUZf6ehcZIb7kfypQtfmtak66sac/7ymdsbn/zfqwi4EwMpyTtPBU7t2sax3kN7E
p6VU7KViFeqtljYLs8bcPZ3CJcDdruajFIAAneaA1qc4o+3rWMphT/prrU/U2mNy
DyUbhDWcFLyZjFYbyN/iurdFcHp3IiAZTTW0UkQ3s7E4qSnNpWgJwxHNvNA1xR9F
vmVcRMAxXp74R1oxsMXdyzVFHq3cP5yYP5CCGpv874S6aL4Oy/hIJbjgSJZgywou
rNYhxLlngrMTdaXdyItAi62c0UNkl/pvHX3/UITjrO+Aq+/Z6OT2vJHnEHysP4oq
yhlYya4nNaCyRTuD9c1tSady9W6bbr3HmFYHdQaOwHCoU8OoIMqw4+cJU3pqK33l
7YjgXcY/ilQPzVP5YDT7K/QEQIWK203mSuJrPdF/WuiR5A2JMV6M3kiCWk2UK9p8
dWaoZVAa1sqEcK3ZumdG0fKnHm2+J3vPAgSA/8eZXLiQXyQjyK8OAnskaja1w41k
wPrKYAsZV4Ez5DCrFkZ6hn06l/VHtA1Ng4eeI5m2OkoUzhtdqUUx1XzwWLLQcP96
GWBk6g9OYql50IXx8AIeWXaR3JHQ3UFZbwdVSBySAtq+a2AiLdc8VGg7eGhfNb3I
9W5xj1gB3+plajXj2/kKGuys9y+oS2/Z3kHXrO79N3f3AbWgvzT91jJS5TZOxhVG
3lhZ3uGUpLqtDQbSMjS6a5tTd77WWdF0Pe9MaJq4x7uzKnyFX9DagB5ZYvVtqZRk
K+GAYziRpHTcAGBxCEEPVV9andTLAvKqfnPgeg6GAEwj+8n4GaVLuSveJ7A75htX
uX11bV/rbEWr4WLjDSvnW87WVtRzxwcAXAWjeRAlMVhJ8Nne1NhCmvA3X8Xx2Oim
rTTlCurLkkPULqSfBQvvvarsLh/Ie98k5l1dq0HZbznmJVTe4rnw4rtwOC+q7nNc
UyGC15wiZnw/YOdX5F5jcrBeN0JdfXJRO/hASw5NjOekeZEArHIKbTux207JTVzr
f9mx5IKfxIKBZlDF1m97pj4/hm+jjfKIHLMZW0wY4Tb7WKCwINLSOlIpKKU2cyv1
c+97gRXBLjmQ/UE1ty8sgeXbBy0/6yHoAG/S3HWTFBBBQAZp1m+xcI0LrtPGWMzd
OiPdJri+YbwdniwWNMV69xi9P9Ha81plaeK1YvxFvUDdQXuJMMCK2b/5rdfZWFGa
RgOsKb9DoTnfUjTthcAyxJjNfmB2EiLDnJpb9sIVKZd+yzT4vtByQAJyOU/Yevu7
CYFAwXb56GdN/3Qiq4K0Q7YAS4R7Tc8jc8kdP+S044PaCMDVrvCrdtTXOE2fSYsI
t5OTlphPXIviBUvviaL9mTEmLuG+4rww3aQqWcWyN26sxzSAYsNCHkdW4PHDeDBr
B70i3y8FojxmgjpT/j8mC5+EYCgGeZXt0zJP3gRL8yRrCNextvvwJcnVwfiT3L5n
aIjHAv9G5C2Zs2wBPd93Wqy3T9ceb9pANSloi8u06+xrvM/MMT8QW98IEMlrfjox
S5oJapJbEGn+onTpwbhpSfFKTUJRRPS/SzXH3QyiQplWmhYfDGlDgh3crfKMPlSL
BUSejX+QZL8IER+GJZYzfjQYqJAh8loIE24JKNA/10GiH7vHOwTzH05bNQqFJVOL
UZ8TW5KvxUit+Sx/2w+6RI/1aUPNA5jIwEgt3HwPPpl2IHbsN1KIzFql17sjbYiR
rq1FMixjx0s0rQN2I5M7JwOP4vyy9c4G87QtJ/zCHTBnUQH+IaKgBlT7oKK0XS6c
yoYBEGUAqRlCFuJWYxCXaFm9RvGDOho/0VdhOVksMgdiM2vKUs0EyRj3Pdxow4Sw
pYHbsHElRdRfyeOdy1OQGhg6CqwTwoT/wK/s8l+wARjHXSmyfx2bfnSn6kih6UV3
DUIYaRTByQQZ0RV7fQpWaWBAcA9pcB2NuBZuqvBsDNUZirVX3WzMtITaXpiEjjpT
UOR/ZmICQYL66CP+qNw0huZISLzC8EMPvpIfPvhKssqJ7MKjKAbmKD1kuMWo3rFt
4TdfVD5RoJrQ2WE5lwgssGj0SQCqEqAbRLPifhzJzHYEG7xYlOqjqXmzr/y6phPE
o8iv1qygzo3pttc7n7oKaRMNTJjJJuDck6OrvsaOOX0RlLDC4JJVjY9akdUILl2B
DIohWqm7c7uAv6UrgmvIRXPBcL8sq6WaN0xQdgoVgftHsbHejPBuxOiczDIIWb+O
qjuGSP3l6bPojmHhCCCLNxqDA1DhQXj0jLeMQzrRPM1TY+uF8VGMCY0036JmTY8N
Eo+fXgzu6uyITA9uLjtrhxtm7ukIv+zck0UfCV7TJAIOlSZAXxo6tjetSnIlYwHt
ucnBTJZdtBhL5110x+7F5Zzdev30BvOCl32FrkqG77D8IlCjp6c5qW6C/Vf2cy2p
aN+J3NzRaJ857E1tBfy8pfumrFaDBomWhij9WE+OBhN8WnpBFj5+xVVt1e3Li72h
SIZOIjNCClK6NT45z+jlTHpu3hJ3jEoyO8IGgyRfqubZA+2xKC20khRTcvYdzTgU
DM3xmvGdqWxnOWPWyZBprsQ+TJJQEI/klCkmnPNFjTDHbK0HxpjOg0G6PdoTvJIk
S3qnHr0D3l5S4TeOG6vUaAKdqiSf95Okgs811xbdd3KoOy3kC06E4VQJkZqN+Lr7
PJoQR6aTFUn1eRDht0sICMJwYRYtD1KKVQKtuBuqU1UccfoS762wZDyMplGl4Tnu
8NYmDK7CPAl51r+mpM84zyIcRxBCuJzwS56msMB7LOVwLPz4M/kvbOUnprIWpGqq
nnrA0qTqOXpcWzYDrlyAO9GPsuZEoBWU7iwVOsN0gOk56a2hwtUG9GtBzLtk5uvx
lgBLi5HxzyNW4CrbML1Rb5biG1TUzZIaRMWAbo+cbCUx4vEjoK+dRqyciWRSEf7I
i4o6Jd7/BxurXaBzT0+ytpGkw0XGwhaG6hFqo8FrSaIxonNTN9P2E72WszK2Wd73
lZbtP3xjlRTMhdIE+OKU5Pbo6n5qL2f5tk7pzSK2Kie8ncZItDyezyXpz2JYnQ4E
reznFK8oOQvPgOV6eqTPyLw8o8ficxWjN5zYa6dquhAeD48Pyq5vjM7T+QsMwS7d
yl12DT1s6JZMu5ZxP3zWTqQujYccsRw4YY9Jl5xaDF8E5IAG6Y4FQzLemwvRe8Lo
cww2s9U2mu4zVG6cDqkBYJWEoYUPOzqSxz2F/ER8i97wE7iBsieS/q4jCsvM36cQ
0PMXqtanzVD9x8nL1PmuWwlZmLgUdVQ57L1KUOJuZEWawYQZGCObm0Nip+K+8bjF
Czvt2XLqubble2X1+d9w+Jz+m5iOsyCJ7UBuYURP70bMaBF8OwhMGrV1oJD+Ev+N
tjr6W/TbmMZjiOUbBc9hvaUbTVXENybgETfUIc4zFCVHxPJRvwt4sqy9tnNU4slw
gR9Sh28+qaEJURgLt67XviaWG7cF+64wcyes8WruUAk4xf7083bHYyqnpGhtZGnt
Wkm6QzU03GipIIR7UOJADjkdRaHrcFqA6uj2RRVmEDVQaf2ae/lbY4oAaE/JB3tE
+cB1pgra4C4S+MLXf9CVX+HaAhPr6C/f5+HtOjzf8x7VBXME2NXlL9lDSWM9mDDr
KcczSsg7PrwirSG4onsbVSalK7cwb/HbWhs+TGz+/DR9zro8Iha50QMbPJ/Bf+Hf
Mp+EwtNEbg1Kojr8etaxZqL3HgsdS8QYP4sU6VwyChdO9VlXIzn6wdHvpd+kNhon
PylFOL/9X/udpsX11LNocrZePTCUTHL2cp59N7iRzTwQcQdAChG5NotZhwjN6l10
PB3oarvBvKbwuMtT7lGJ63KTPD1ps52M4POM7PIkPW8JW8InnEBKB62CODxwYYvk
0qcxlnggXphgg+pS8C424Wl/PAA45bDpLpGGw7Ldp4lTLOGprlpQ5ZPcAs0jiq0x
0d3iEJF0lnB2y2V0UNT1qQ/QxfrZA+dkvIA+mWYD9ebuRwTfGfIjuEHULjdbSWEW
NCg65nX/+kUIUTUZwzO5LvfShxFwngaceHmVnf6ZkoDzTDlzNQ5FLjL3VRtCYyvj
PJjKLt3OpDGc/Jix74fRsU0F7ZcyCJrftiapb50nzgbTbLnYNP/5IL9T+nOZMN4L
kTFtXhiPO3RfQmh9RO9NvaPftmppQKEuAk/aDol+T4W92sOG7OZngprcxqsb7375
PyW9/PY9MFPkUkoYgyKJOe9evYj2nFUGjqq11BaKNugGK6DqiqeHpR2lHKkx7Fgn
296RUeGE5EIWii5F+5SYdc3U++6AB7VUIOt4oF4JIk4aL2CAgC0WrzMovjZF8lCl
gM0UpcBPkWukmo9iXgghp7DNmLboJz3snlw+K/bNIrRvqlj1kJWm38t3b+ImSJKC
yNW24z2+YdZny0V4TvY7teb8UGurHRzIwxapoN7q+kqX6sslz18eIl/JnZDk0PHb
AU6Gb1lppQ0NNNL89F2jko/WWXpclKZU4D/3DuJif2vBA9huUx9QV7CjBga+d1n6
p5XEvkxVjOBdWofZggM1tPgAwjCr8r+8i9ItWWC+/Ay4nIrGLDw7YvewTkvKkNBN
ooZEUmDeg16FFc3ZUNQDNoiXc2wGWjbzwdrhOXT92HfiiPVeQJp0dDJKw0sSsMse
U3Ob6l+xJXRzvNuo9QO0kOgkZ4QKne3k5m4nxEgaAqhQbsgILyDdZSebWJ1I4cla
ubNbHZunQhHC0Mtr82R4U6IwhzayfU5Gb+sXL0Do1MG9lcgnXexroZT3R9QQS4tD
WGKpaHoHUEO7u2DYNtFvJciDdGjxoeBqeXlYcad4izY5YwdTIZaB4cCuNM1t5orA
n45via9e/+JUr5lYhhHDxeD3Qont6Gcs0xrzByJb2lhnly28uyv4RarsvOM6OThg
+V3eChJLcbulViDmC7eUef0Hs4a8YBPQrmFWqH4aL0cmd7XniRnqp88fSEr2xiv8
e6gpCmino9WQd4uZvkYNX9dyYQH1QtMXLc0W/Oll8pM4I+STvT4XQC76OMtBWFvQ
uyjutbQqASrUwy9Y1Vh8fd9V03SOuClcFNUdqxAo9ouTdGxNPOaKLviTPvcqIPVk
erEZp0jqKg0QXZtSVqfeXcm2diUCNtucIXxuhkglNAGUxz5+ja/83cxWWZa9cMHy
Q1bWuQY003lsHqoTwrhwUyJR0pV+ba8ctPWvxm3wn61wRO2YWqaCB+sc2CTKrRpB
2HKM2Av3rKaYXKJnOTMxdUdo/rG3o24Z50m0Ba0q0zCM7GGf8gIdWesFt3OAE+wA
E3GNXJiTnJn66qomiDf4GEN0Z29cYzs7+KOxRmwYC4qwiJkrNHDUYLhXK78NwQlz
HAZWDgBYCkh0pkdF+jETdQtBQol5di1WmirlelNiNRPEk5s+xwTSSRW2wr9oUS8A
2R9Kf7LAgxmDBmbQsW5eRRUT4+OhSc7gfJmCfj3kvqPxnf1QBbJKUGn94Tr0Epjl
tqFO1Nvg5eXhNbeJUFsDyEsuV7AJK4XhMGpAARvFQGbVLDomLvYMay9LwAs4nmJU
hbDjhIz4xgxe0+tHQmRGB4fVyt9qqhfhw0iEjzsD/6yodHHW35XdwtVqmOJRDDLY
Ond/qX1KXXNXqCQoSyTj3rAs1oi0eP6VWLM9oa7+GZoR/G/DYbEsDrMvdT84Ztal
ukYK1F1LzN2OyROpj35RXXxGIxL1MpUATP/8m56Tcr6DQncz1tuvyBdnlTlWvS/Z
QNNEV12XArGexzGlwWW13R+YKFHCcU/pqY8PCtcHcUHIcSPXJSmqbkwwM4X8AXHT
ybRlaDyzDr67avFsVXhwY9fSIXb0tZjN5kkNw0kGgnJpm25+kTWEwZZwXAMFkkyH
fH2uTUhpmg94AVte3AlCWrzFKN2p2F67sOxHGPjKI+/zZIZmood/l3bd9nMbC3Lt
SJ3rvcIyElaoquSF+PxOIIR/bCNN8YElC5hej5nYzgh7wqUzcWPsMkPA0GrYpQqp
OrK1IPOsz9wX+u1is53EqYj+7YjjzIDgeYxscAG41/zBXu1DlGV5ra9QXx7Kyyig
JJuURFpBKX4X36RJzqrXVwL7aVM/esIPEgtLHMshQXrchnKYZIXwUsJr8zgo7WsT
HdNlon3Jr3YU3kKXXhkmun1NgBf+MLmt43Uws4lYCx4xPi0pwBiTKB1hP3KeH0Oi
16iEXnAp+FuyfAj8fbQSqgHVZeS2BA3C8YQJ6LNMYI/WgM1nQdXjbhX7pe7Qe3yq
LQCSz8wylh/aYYWx3VynwnlgywRUrxwr6XU+5xKn7+PosTv+BWl82ZfliiGv2lYr
U9ftmuPfoz58LptN1o1N+2/KBYQRCyvad2SL98H3M4lCY+3SH/JJnRe8J1YdI5Bo
5SUf3borcWssV3pWK+h/3IwU9yE3ar1SFg+1Ee8D+C17HJMHMajkV9JmSw55FfKn
Izcz9sd6z3ShJpx8ImjgiWuVKHOZJxzcbw/RDDb34d8sQwXdX7i25g99aI30drex
tNSICWUkJKMUqTwJRadv94asZrYSeQKOIQSQ8pIfn1rFvaD2T5wEVRlR2AeYQvm1
o5QD3a7HP/DC02zNShL8Qd2UKBPK/hc23SHj9BfS42X46wxiQyKDm2wRNsG0E42n
VR74gocB3fxDIJA7KfgKTwDA0IdwzIgQS7RXvaV2QEL4MPmATktiVs8DULhkZ8g/
QV625FufsZvzg39HgD222W1/wnnly+KQsKMtcsFwDpsWFwxcraC6JIRAtcBoqj1J
oHJYInetSXTeEUHeXMbme/HmEv7ZsGuog6EXVwS7HmcUYSLE/5iII636Ol5Ngyoj
cB5fq4Jhg/nIahrd3Qzn0cfDNfJgyV358wevF1qJ2tdZeC6lOBOQSbtLl/FT+x1x
Drs2LJ73thyuCpUoZTlP9kOUKdoZ70qlDtZmBFwXUCoSgqgmOxv7/bqz/xkannBZ
msa3ysmzcC5ZlTVBc1aS4Ynw3zwcO57HNXqZG+plaZ8Plm9xUdfnHZLX0xMd/stO
oS2+v1MZk11adfOfRMieuvYtZJlbFV4rJP7lBCXMVS5++2kq3Urj17a9J/a/4D9k
AxTL/72pU85LtUCi+Blun0tHFm8Q4qo3R8w9e65l6IEDgokoDcTKpfjHCfx398Ya
wJphv+m3h5XYCyqpbs3blqedpUV7yLKtmiExdEuzLUN7wPK6EmzU7GD977XjK2G3
zvZ3Yq0017qFX0UvhcnAxkLESm2TgqJ62arMKX+CTMZMnMGDtQQsEKD/0kkuhH1T
LZfboumX2/ZBYRrAYDlS6YSO+d49Ip0eeB1yPWKuaeN6biMLEwW0ZnDKtnb08ttw
qB9WZYXAtUfEmaJDnwvVl3DXk296ZaK2n3CP4jplC0neh0iIIz+IuBpqjcdw6uM5
bhulQD8Rn3w+uF711RlformaWvTDJGLI2Lnzb+YMlhkrFwcQgbiGrADMlxSFFPzI
eEhBjmYxI0//X1Um/qJLoQEi1ouZ7QUBD67J+jLsrAyRnA7fV2bKgjYlZq1h/XFo
hGahzJ1KnhHw0NmWry7obqSUe+erKAiPwyjRQlHJ4mIzdDxYv4bs7+F0UwvHRzaj
ygBVdLF1J4yO5jYnNjAh6IH8d7slUawN555QK0imTLjLrXoPSzPfgKKNByzFZIoQ
TPuN8lWuimEemIODuOae9kVDwY/H8vz/5DypmeTUxlUDpfHhbYMOS/uexkPvpUxi
stRXV8BL86rqYLNsOVyoJQAaXbPvOzhYmXqBz+lEHCVMICYjXih8g2E2Q9tnW1ma
lBbZxhWgplqcW4zLJ6qkRhuqS0nHxZClhWJlbUoEt3mFIR1r5o9xwZqtajxXFIPg
mby7B5DKj3o/q0J0fHJ0vzYUzXieC0I33IoxA1OA/J9GqJ5kgpRJUvOekhI4xgpM
WeE3epNRRrBOI3/cJefR+e76Kpm8x5RqrSwPydKexNcWPwFZyL2W2yuNW3IODlnn
aG6B/8dPJyf2JWqpUJ3Lm3j4WkTA2z5Wpr5Ip7eV2lJeyXCZ4duRYUtpaVwLQs6j
wOZ4TIlAGqopQUReouCnhe5P8fQKsgkT4P6GAt8r3Suwr9j4Po4ZM6ptViSwFanQ
ZbwmQLZmxvtPbC8lU4kbgEufFDfdL+2ttsBzUFrYAC0TUc5oG7Ce1GMIctITaYXr
qxVP0ADB2XGfU9ieCcPcKQxsE5RXT6Wc7U3sTROlwhv/VVpbMJugy8Eza0x4HYxv
tIbLAJ0RAlJF+HOGYhHimn6PWEQcjaVwD7HqExBv1v4=
`protect end_protected