`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6272 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpBpbsgrlUz60qXw5n7sklfCh4l76WPon6Flp+0+P6aQH
0aKAKrZyFq6+MPb/6YqAFTmbG+u5v3IaZ9ZlJWzrCGfFcJ5U8hx4fsivrk04oj63
h7NyZNRVhDIVP7O0khKwX4diYFdgD7yEUdIPLVwEk6JwROsSnGqyv05sSaLFbTCM
4d4sc8jqRKFPuU2YgcYMq/LIzID/NlNMHdoevY6OmHHYak3sDrjv6rdwVzu/4hId
Ag/TwyWRtxan2HqfqChLZXpTjFcn86BhOvwBNKnXHGz8pTNE98PUmRqGCNTY7haN
8MLJ0TThSPX8IAOmVTVctD3JCqYlZl4I5P4PZg9U7ZvhWF7sAmIzISbQNp2vB0Bn
K/FK6GHfCWDvJoAsoGgItNKPS2xygnpM54e8EkWCiE0VxhZkjb9T2J/8iAZ4zYOo
0HDTU6oiFW7tB0RpbVgwV+L46OU2Fw1Zpy/7pxMZiEpIyN0EeJnM7nXvMrt23+zp
zbQnysOC8RX0rnnDwrINPd3o+EHANOCKK6baPINfQ2A+9ucc05ZfcOi7+mWL01IH
t/xcSqwOTkDjwNDSTU9ieDI2kP9DbndrvlOLOiut0/tVt9/7T7w747tvTwzDOb00
0Ehl4aQ0/B6Bsvl99tOHP2I3ib/I6KKIt9wkwiKbIeNCk2jPJb0FZyRjmEpLdzc3
Qv3FAIhBZ02HEV/0xD4/ytfpk24dW+mgwJxQ2PT3E1O1oxm7ckoLeTIx+ui9ufpq
Qp/t/4NzP+mxIL9Jo5yyMubmMntzsWRrj+E5K4mWbMrHNFglKnjmkO0A4OTcgU0O
1aqKS5b/9jKRr/MjW6G7Mb5Mfu41U9h3jfcBy72L3yGr2WmnIs8/Y60aQYEIfM4B
QD0u90psbuV+E/YksUWHR+vjtOmz0FLtLOzXRzDO2hn+zheaw8ryQYzHZesHOgUV
9tS9dE/nYQYdTFvVy/oGsRp25HN4+Zw+nZs//NoXwm2WfkJLzMIqyk83y+addQwe
b78izE5SysG3K8/tjuvhAfDMzsNZuBxUzdxvN5QqCOP7EM9bUdQS2FWZ0XJpleTY
i+ufUJRgjzqxSktnA1o7bE0jqfmEPhQe9GL+z8T7OfXUrVmbG4d3hLBg92uK2aJ9
CmbxQ0DvnYFVXMUs/FSFmOKbk/sIqbo4LYBR0j/DhhFj555Mz6Ij8KGmLnLii3yV
+9MqjAbK+j/7Ghh41xpMbG9Q4e3uIcLa0yoS9z8jd6F7vmLMeSBKfldKP2HhzO0P
GnUvd16skJAI/613uoVXJZ2wkmBaVQY6uyucsfl/wnxgyWnRbwhHQrPy5aPLClA9
UcfRiIDjn4BxpDJ67fqYkZ7qpfbNI0XP830LQZbAFcvB/T2B1tx1eMrlxesW2yvB
F5+Nl8dmPD5g93HvX3Fv/Td5av+nOkFr1GPOekyYb6mmXYoptODcSQ82eU1Hbfd/
Yqv55hfyOTrEiKhOJDOS7y+VbZE2D6A6r0ev4a0nqa7d1qIcpfDNKbPbr5R7Qa0k
n8ktrBuUQglpV8Ds3zldXM3KNxmH2e9BFN7A4jS8CEt7ANxYTSeKUK/1KnpFX9eR
gCF0dGrMxBLeJWcgx8aEkspr5F+i3MIq9NJ6x+x+VklXChBhKN+xcRCDXSl9slxp
q9nnhv8s1QtTdtkZ19OIGPE4TrmvQwn0jkziOaK66Vjqzw9bCcIBjUxTN/lNNuYi
+vF5AEAe+1bvoPzBkUH3vjgrDuz8T7C/nO6qy61uOxqmQTuA7dDOuiyACwM41rbA
GLxB5q8g+bw/Xc+7rMNlDBU86e4mK92clgVURLQnw9GFyAI13ex58vSIjd/Vk5Gc
g2hABeAWyWajU2/K7FNvCVEENRd1nHAWcE1XnyCQYT02CDKArDBYUFQUoJp0ehf9
UJIO49d5IDh+mlJnd1p23GTV5DYvzLoje027M12f1bjUmDTi2b/R+J1omjFkjX9f
lO5h6KiwqJw2Hb+zFhJDFwY0/aMxN0+vvBBnBiqILSzRhFJ1dlvX8PliDj3nsaE4
giIAbKmVFoAw3ir1cw0+gJ6/LTFqDwi9uuNOfVHZ1Tc5YD2s6OKnpS88Td41R21I
CnUatMoE57UqJiTYZA6ojHOUIOghn08nLC6MjWzeXEAIz9x12fSwLFSMXAkWIkcv
HWrLUGK79VCUgHPz+jt1OY0Lq4YAs9k3YXyOX/1ZJeVl/wHoeRiADOuj5QvgOOux
vCPeMOTK2JxXCdNMvGx5Ik5A68T6rQHx4mLnvR9I16/KLt/56oPfyFAeYrw6nuzl
2OAZF/pSD61qsHdZIlk96P8kDthKZWVI3+zH8c4vRb3qAIfs4kRF+pAVVHJevdes
eHX7NSFp29JZy3NiqzJ0O97EV0MeAFXUUE0KFJyF/cVcMLGWua8cutZ4QSIEs0OY
2YXVEK+EKIdukRjuXCSxpsubHer9LGFCNWE4C4a9U3w89nKzUmbVH6J6YYclXVYa
hygLopf+6BktmmPGInYhr2tNFUHjMuKweCsjsYL8blZ6mAGCeg+B+7r7Pc7LMfKJ
5vSdp5gLH4ipv4HwaVnamY6cACr6Dzb9JrujwP9m9dtnfg3jA0XL0qmVZij+3Y9w
bcqq3oB+V2pjPwKJSL6FLJJtfVPzdIwg5zpE89V6ZaWmuTYMbp17CKwJaGXn/OET
9lnXIbPAB8rSvdcMl4H4PQNVCS1sFxObwqFejJ8aM1AfDo9Frd9CVM0EivuaFDiJ
243suM6IKNtcPz39+IZ4Zi+E1KdgBt5Xt3YdUybmNLgUEbV6vXsOd8Pk7LCdzZf4
6z4zsD5TbRHYHm7jXKWFxPTyfi7B1eXeJiCkU/OvtZWAoYwT0/h8qkyLaJeIjuZ8
oijUEpHKuNRQFBpclji6k8Jx+op9fOyNz/yEQjdNHY3SI1DI4iZIL5z+Xy2Rn10q
MNl953aUyv2c4rwEsC6l2U146lSVB8O69U5r79WFWBwE5Qn1FosUXEH307J0dmZE
M/+i+zU3j8eQ1fyF/Hewvs1PocZ5NT8vbfbbzWJrZ9bxOi3hVP4XnS0QgpXogoja
1uydeu2RrmhHNYPjDxq/sxtx0ynsIUnc2UuIATURxYbqiquQTGV1Q3eBY+Yw+KIf
g+XLGKW2+oMjqKWWOCHWXSrxw/NNSD+cI6dYJHNL0waifxkqN3AKJAaT8uLs+0Z5
wpQXGH3uQSE3/oEmJRsv0sbHm7317Tl4iXHAzC6uP80aYXtDhHDpmYTk7dDIe8j9
bN95LUXWsNweA14vPs3pWMuZrtZ3C8Inz/eEDzgIY9UOuFPz3Vbtnli0lvgMbk9v
P9yJsSPcaQVVDto+yczqIQNIS7LtatxhfoSXBvzdCkvCktuzUjQr/guz6U+9Uvec
4Lmva7N2vRwMbL1ZTuwiZebA5geJO756Yxo08NM06ku1rVZlUQi1TTgXOUGJ3Sqv
HOB+GXCAeUGEn1Vf0ZVGyDghQ2C3cEJ924duHyZD2M6Fh+Y5MUMvakF7MM22ydEZ
DwBc8dKRnXmE4v3l2WXFoMRRDdj2rJvKK9fC6MsGUazYzAvTneqJV2gk2DCOVxWN
H2ixEypgtYF/queNwC3byzrSRmj8gXJioPO1ncyN/BYeGM/okwV+Z4gSXvhjewkX
L4zGvW1ABqR2x9slQyJdrx8vRM20nc8ftkxOcyDNkaX37eCCbMx0BxUtVCgQ/Oq4
AhU1PoTGBRPn7K5oZxtzzS2RNcx0HtAxb16cGNSG9zIlyfh8jab5pIE9lw8jXsGi
65+W61ANQz+fYh5KqmImPAuwHoF7QvIOPrV+RAvS9/ynyd9tWDOcYUGTl8l7B1lC
g1S1yK1TE92BZMDI2NTAXMIH7YtKVC7DdgJe3uGERXL7J83/ATnZjIR3Stk5mW3V
NgQf87gXfEk6MLLvBbbStjSAp6fWfnULzZo67u00BX1thoJqlNEeChmXel1sK8yU
arUxnOkMs4pzUZYUXX/WGpFQB0rxydtqVKNwURmwABh3mWF3MJ118kLbjRHpbfKy
GXWBUSzt08yXmk1MXnHGxe/B5w88aatEdHwdfATtwcKasnSoxoPaIEA3LgtD/ups
qZLHlygE8S4Q1NAjUuXrlxev0npgKioRTK57QDNNqfjut5xqjAUDO8ntDuv0RIn+
iTE7jQyze5j9ByxdFciVKqPbqTS0iRwF7Nqj/vnEH5FpxK0heObg5hIcMYeBrud8
I1fdTspaFjb8fQXzcDcjrczJCTFzvoBw5oApjd82TLdwO88h6DiT79XZwmz0Rowz
MCCdtd/3VRvTAX/1IDi56I53GYrgf6cbhOVWgvNFgR6AX2DJWGDJFABeiGHDwIym
rUIe+OtvKM4IcZAtMG59xBK+Q0zi9J7mgow5yX4v+NrCPHTc5E+ExYn8TbkWgFtE
nwAsPuEhcuCSCjDjz5Isjk1kzcIckfzNoBff1GHP0NYa0txRwVlbtHASL92P9V/C
H4ZPp9VUeQLzafGOFt/LLYGCuLD6Jkjv+Pfngdu1kZyhTWDfgzazSGji72LZbkV4
eRjNmykRHkNmaCZlEDNt+U1mQeQpAq5s+5bhBibI1UEhiq5YCCTonv13rNSFEE6/
t2qnWgMuPJ9LW7LJ1jZxfjP7xtvla3WHubJYkIRx7zP0rPWlr80ucBlt/DVlYEpc
wmL5HGDwKtECbJHFNbWrNa5YJoU4EHNQOBYiSx87zfyp20FMxQ/jy2EZjDP0W7s9
l/lEbIG764iMw+WAir18mxIDEMCTTeiAzg5VHNymPdFhPPXRPi9BtcZT399ZfW9e
OeLgh1lNkNeyr8zetBB2GDVwzciLrumMOEZ2vom/xjc/jif1Hxp/kKrMout4dnNx
DsfTR/1WBNQnHI4Cek/7cHaVfQWZ1KXiCR4BIJveFKUeo5cA9CrKFfLOAUtj1Zpp
nCeTAfKEFRU7Ufq4UJ7ef+QsYaoMhyFm876eLk9+T148qB++wJbF+keGhzCcsqq5
1+MrshSQBsLjk6vBrHil39/fQ6sFHPnN+sY4HCDVwEkSCLLENOgNTQwaSDkAFiWX
LdsLHCH3hAufv52tAsoRNo5PbJ2D1R/g5OYsou2QMkuwMJDNnqaz0MUNiL2HgC3m
lgum8tir3ScsDz13AKJQCu43//1Bl2R1/2T9Hasa3UTT4Xm6wmlA+eLwmutKNZ8M
z1kIRmvUPGNHrIKBFcW0LDNpQmV2A54IZApY4uvhkLiQ16IOHRP1LbFPLcwfv33U
B7z08/FNYiAPjNZ24ubfQ3N1EFjjk1mGyK56n+YhhF7zMt7o8enoE3ApLkqo0sbI
Rf4UJKb8Abaop7jo+YeTc0uI10I+x9grCvDFOZYTF0Br10Wvq4Gs/Th+r6S1xFYs
mp8BeZ1vZdZ3TcmSeOd5POmASeaXbkHKUjtiTi5PBVnw7BUq3qCiAn8GBUyxHBk1
VbOR8/DT73Es4FUAgqW8RRZLw3i8J0i5mpMhEd4RPDR3Eac8KcGgVRv/UcNF5/rn
m60wARpHd2USa9AFPxMWnJxaWyh9sni/8zg6y/Jiw1LA9iqB9xzBnm0eb7k3CNcK
7fJNdScCJGKNpeUFbE96ucdjMe2WhXnBI+68CNcZlcdGnwv8WfuBevt8D6yYT77+
XIgLNjzTla92NbR0ADQb2faiAtN8cJOA6N7NjxcBWfa3nRllZ1m7nJB16paKwh1z
hzw2XVFKUMTL/ZvcyPK1t7tFShhBDfGwRDUZZHO7ZrTKtgmPFWrtuaQ/jP5h4fSi
JLs/KYWaEDWLb88KE6xhM6AWgAWWNKwLRdDbV8k4jWtN1nvnh8VbG76kgRMByDHE
jTNbLYaPLn0WYmukBiuj/HQDeac6U7pw8VVJTOqvRu02+Im/W6/vTiL4E7O4UL0d
Yfz54jW56dBV6bpSd9efmkVJ9q9rUZ8oQuqiNzsfx/thxh/68z33UZDKyxFzMHTy
1eglaZ4lx9SfNdVwgO+b7vV11lkMeQ5foTNjJ7SOhH7i//grXrfE2xSCQthqSeH+
QSm/8m5rkzoY7EJXVJ3Ck0sqfxawIDxLExc7tsYhnpiRj2VfhagB9EVshc431hCC
m7/aC1RWJp6ZgcUQU82PYgz1fclxE1Eo4NRBX4/Fw3m+ZxIyLTQPOwh9R98daHOV
RabaHWIYFtp36lmAo/QNUnCJDAHK921UnUWpEka6K62TlFTls/8Y/PkUr3dVy7jV
JvHxteBi+EgptZQIsmb2WGjSpqwDKklEyLpIKcjq4IjpixS3wVcKREHjnWN6aq07
gl3xkmTstFGGS+ZCIV6z+DFEFFH+rO8QUsIAcTifEptn6oDx8deTk/nLCTzgFYIT
DoleAXqwjtjDNtuTDF173jAugxEbtGLXA9Q36It2zQ/yZoty9KFQCWbBg1tyePnL
dsAXTg1K0mFFCcjRa35/hEvzCC/5L3CkYIFCjYR2TObrujNtOdnM9d4GydbbZJBH
XUgZ2F/+7EEVLgubU5ndYfqx1oev39OYPWEVCFlkxU2LuDNtxui5KR07YL7qvIr/
tzq4l+9ooPxnOsksZKhtiBuC1wG7VGF76XYhC/x7YprEa0QgTBELuB+xi8My9I1C
khYAe+eOHZme6avH6WFsIfIAvJBZk9XwLZ6btu+fl14bSzTe8kToDlTmEgUFvLTa
VU6Bqnt5CghXSuNs4C+pVDUqlXc5RLskUE0AWX3SgVFwT2cjPf84yRLeU7rstXV+
qJRjamRhhHhUBCCG3hHtzkVPr97gaKqTnI2uPXoLfPAdYVu2V91/ZnsWVG84eivo
n0lJugz6joE2bZE/9RkRo0eoVbVshx4GuROq91xvMDuD+CO0Ko7gRZasa9fkenBH
9iVrmZxHSddWh69JyQSeRGUPfbi35vgx1WU/DY0AzcW7IBaGRtUvXwFcBZaCYdbm
NQ43gboGYUWcl5lS4Rx8S3OReHlNBAzBQZDf22Q0qzxW1TIeZq5b8pk8fEWXoWA4
ZqO8cCQky4iafrBtoaEsHqC2boF38uVIlOXaheG0Uh4CZNu8iAd2lIRCBR1+h6BE
itbmqYKohoRCniq3yW7+3BE5jofxOeaNLaLJWzLjWz2y/nzFIKGZlQiU3yZ8EChv
ko+fj+i97SXoNNNbjyGVBlhBoy7X2nbjseOqpeSbE5eOIeh6G4NI8gkPRMLoMYIA
0tX0pYLE1jq7f2QYBn2b+siociPr26jEHfWiAhYDC0VwTGJSV42nsXilrgKQ+OKh
dwvtdkag1AU6lSOdZikB5/hMHYgotpVDzAC6Cs0+cWL+bqnKec/OW/lvFIMkf/Hd
hlgFdtoSl+aLBBj2Y+uho9KBAhC8M+BjirM2y8RuCn0x3LbYQ3YTlV2WPopGKraa
yJIRHuwIKStntKxXEcczxtB2fmypERrvnkHQWOqFG7pRE1ttxrGgNz4o4c+vXcpe
lzx6EUxljclzRhoCigKho2esckzMPFfH6281zNnJdiM7hVPleadEV7FGSCw6Uy3j
pW20Ba5v3Q8VSOAimhqaxoX51vNApuN59VvInoGjoBhrZFX3wWd0ucmXkk9RigJN
AIfZDRcFyfVEDUTzTT2AdsQ1VW9M46BDYkhYsgtX0t4UCdZYrKLH+XnK7RlmpvTN
o/4AoST1pf8/YrBdE2vULVb8chO8DOP25OPxlpHrep5FGCLvUdRIbADsfTNEKXeb
Dx7VncSObaPuHNpNl7ZRMYaW3W3d4D9xohgDSCZv+mxWIB3FjFl2j1sluxaP/XeU
65Pw2engeVfNhYf6NYEUCypTL860GjDPU8wYdAG01pu86MgH/cR+UGFnZKy/kbEX
2aYMRDg9Pz+3BxJxyiL3fXX6K7zWqoVQGuE8de8hRcsLRVYCJURy/s7ydM7YfrNF
fpCI/V+vyFF05HuBM77ChD87qcg97C0gnQvvmZpWC9r7y70Lb3t8mxUNsFf28kJr
zvHjxHgoD1XxrG9nDcelihcKOAoXpwxE04D1pLV/Uudz5zQ9RO7nGS/24PSwGQIX
cTPKsVk6ZSC7MB5Ffu6F3eC1eXEaCwHBlV1D3cJnY/m+YIQ7tuEs2Ih7VEAZ48if
wLAQzDm1X6uhPHR5XqR2OcZWJ9rrjcdOK9cwfvoI16vYrrmuGWtQRzwJrdMg0gd2
OmuWbSgp98Jr5/j8C2HMCb6ThUTLBOucKvyJvAyNEHSfIGhUKPHaOFzpgzwATOH3
EVtpGgX7hLv+J+ljrPFKgw4S9srX2jND2o5BPuWhZUs=
`protect end_protected