`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6912 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
DZr/8BrRXj0KUruQ2Zf/9sOODBm/9HDMbaX+5gKOC78Dpjm6SRMzVUaoQy4UCXr/
/BrwJETlmJpfex45YRdJCsmr9FW4r4K1F7ZOdJmai6+ac5lq39wfL37/so9dVI7D
UDcy32uKv2VuSZTmt+Tkas8P3Kh7sAWD8lbRLhF8G9bfT0zpFjz2ipe2/zcxi8Ma
yThwNnDp5WU9yAUrrRUEP//NwrHuepMFIUhOL52Bx2B6GU8Og6JO3c2JSZWa2gn9
Mrc1bebUo9fGtEva1bZOSjXxNkChkHpPrImMr/iXR/9TR9nMqtMkk6HZo2kl7yyp
kBxFy6ObfbZyVYoxuPptf1xmjOqa7/RHhEJeLHLOJy50kXnnYO2a5cS1r22X9iK1
TXcYVg7Tdd4MrI210TOxVPJQuK5lWhQFamI3homGkUeE+JaHcbgu1Aw7mt+86J5F
NYZypfopzOnk8qJIEoXw+23/r3YleBKheskxu8L3X31MMaT6d4vAC595BWZxYNIe
Ty3CvJaP7T6o1v3yUIpvejDSbvJmVlCd6JxPVT2pI2sJO0ci0/03/3pf53braBb9
FjnuLDtsYJjV+rl9SeVpHU9ho2lNfdZA2o+DADZyv+SzTH8QI+Hz3K/u794Y/Nv2
PYO6P+XRn21wuDoTJfMpxpkD34eT9fdmDu5lL0AbuJmxGhtJs9mhO3uYQUfjb7jd
73QzHFS7kDfVOTy1xC5KDhg5zhFLyoFBXsT6ousTXUWZboQSepbxj74SybEFuZ3e
bd8NJ0n5exhIqFaRuFF6UBNDhRNzxgzjzzcKkEc0766G+/R/Hvst6B4l/+o53AXx
Sik9zEnYDxcbHIibO0HK9pcOKPqE+n7oz8UTgX3KTmiHF2fl63bSE5QuMkt2D8du
iKgTRRXoBMJdUeuuKSs9/FY9MshoNqv5Euz4RLvIOq5t+RP35vwuoAvg7z8GAqU1
X69aLenzZrD67zs/KIikeEHETUQ2XobGMQF9O7Cce0W6DfmqMaGtl+X3egDdfUhm
Zy79P0b3QEkNG2Acl9v4nCoC/rO2Ik43ZrUP/f+NppF38OAXU2Macn/9ua5Pw6ze
qVpvQT4n8MroVIjrLhis2AvPIej49U3MRnorCaAKbV9TICgbKn9sl/uiGAo5LhWT
l231P6uRWdrL0PvmS+oear6pudjXfZNl80qgFFFsrslZHEO3NYzwxN0ue27397xH
vyhGpLvW6+Jy8wUx9M53Wpw53zQ/sr9MqK05Ps5EsmWmyK1/JnjoSomRnIjbZFVp
fvie9m5FLT0VvQ0+3kuVn3t1NR/s1S+DtbvqJNsjYCFbkQncg1I02b/XKar3i0pM
0fyAWksegAoq/YgMZ/sqvutztO5rDlk4QjXzlI2uKJEO3vFT4G8c1Mf5Txc1okBd
UiJ97GXmBKmvAOQD7TqS3zRi8k/fYsdVuq85jipH/XywT3nx7PSpjZHbFM6KNvfN
hLWlsNQvCI0GHMaJS24057Kw7PD2uJJoiBUdMmd3VgYkLUt55BYUUbSAG4b3H+jX
O+r9hCxnU5TQjcHl7f9+dbHGuAznGYDJRJnUELeSwrw3oQs0c0kksauiv1p/rlaz
+hMuut9IUgTcx9EB+8NtU8+QJ9uR61B8/9ZHXcXeDbTR1sSXCxSt2xiaDUFnlSpy
YWeX8PUV+ouRjp7Ui4pww4dYQTJvCGlNs3LPKEHgPObOBZ1+K+iSwbDsMnsaAk9V
yli+IfSt8w2ie+Xfwh2+syHy/gTpewUbQ/nm/yc5Owfwg46mch4Isu2q14uqdxIR
ljLbVl0VKraZwgm87bburyC7OKtjiqVBY4XWtAoY0+BkqSexATGvHrwv/4DS+idU
d9pfdYZZ47/Yn0knXu0aII76PkS1RV553vSjkmawPED2o1Kv0kQhDR/j89BxIbM0
jmQBEPFAVcGji0eli7HFamb2Dj02W7C6xOtSNx33/pW5Du+jybEeR1PfyGLE9srt
afZNdWIoR4e4Asz06b6QsTFuBIhgicxbUF8QuUno8+urVWRpYBEodvhyfDPevb1w
MhH3ZYaTCrSW9JvRP8x08HMZk/24NKGDpsK/IwYDodEqZ4ABNA8j+SROXHehhPrT
yzHVnDuKbYdTJyBhT1pLjJzRN7UFg7L0g9bRJXvtSqDCECX+HmJFEoNrxWxGSJsh
mCiOC+q2Rl9hhiOMm0OAofjN27fxkt2PZh670Oj4pPxGzd84QLoMlPAOmqXfHks1
1OfQcytXKa9yQg0B1kDanc/PmX8gRv7CfzbTkOhc3GNMWPirmLBvSVE2AK88UE7p
G2A4CTsWrHs04IfBtXQsqajWkXJt5I5bIymDtN9qzTC5YVMIC4xWMtVmjvaRGnC8
o8t94gL7acmT91MzNnYx7VEKLlLOJ19Me2wa+whjirnpZv/GjtGcuR6Ud+GGCM+G
jfk64NAJrMDGJY6opkevNPU9uRrdI9ruuShAeCC3VHh71oUnLOFYSxTyx5/he06J
pbthMEhm7FwlwT6cLw271VQ3pK/+BOdFjnijimnthbR6Ca/FN9hzZ16VXKqQ3LTK
JHDY6lYszmVTh/1eRrIKFqLNVynnNYOuxqdyoZiUWgOhL6aZqxpyXGIQTdqQ1EZi
r1IkY8qvS/feOy1YdOzTV2OoCwEyZhydNo84l/CHQyl625pIxB6kYe41jDPLpnf4
ztaG3AWwq9xRm1J0Hfw0D1vqEzKDJfPOvJQvuOzHlyauTAKlhX7gStXTll1FDFms
coFN2cMEbsa3wzU8IAggGmXkGYVZthUNdGBgdPxGZYGgPMlJdzA8BAuy6z8gXc18
dILFSoFuNwy9jJ2/9LA8czUwuDN23Udlpb31q6S6pcUgeQSHqdJh3q2/kZCIGVHw
efluk3lF5UhIOCvBBzFDUz8R/M/tyJq7wink4XGCrlhG6spscXp1win7Ym1AyGp1
5YV4ie5TwUMNPzLvXBLQIRL1yh82MDruylhSD+6jDYWdnFSYLgVY/8E7RCnFXGrK
k2PrEzQiE6KxV4B0F+ci6nvFU8ZJhfDHlySCjtEPxXacOKDzmfR/bbJLEyDKGZgs
Kk2d7wcbbzZ7HO0MXF+k6Q6tNUg40KwZP7EZAc49TLL4cH3JGPwQNg9P5mFXvhf2
/mRHjcIEU1A3dJODsgeL+kuQZRElW+YFnGTmFAzD+Z44DpipLJTfkVvJaUSy96Px
bea98tzWsiCzqne7ekahApR2RZbbZ7ysaFcwSM2/G2Yp7OUfL6BU7HKrBH43Dvye
eIrr57JPCLBfv9E2mTZHqcBtrfSv2IEkWwBuX4DnhVIWT/iFUwIgaz3JOMJhleiD
AO6YdTfXrTAvLK1eXSgSzKXfmbE5SnDBkYvSVMEOtIWz7rbumxErG+suecFF+n3Q
lESWL1aUtgnLWIL3FxmbrtFckcjfijrAi194dzUYh2v7J8wwaBXfRgR4DfkFMg49
+a4VkMeriKZfdr+mzO6ZsQVumx3A5E+qFcQLxVCR/PIDUZI0PJs/vV9l/UvAVDLL
D+umia0Eq/ZyVnnT2VRkHL401R4ZM5mSRNmkOEzDNwfTKX5t9lMDqXdjNlD49BUy
Ps1WFAhWdyCKcwD0ESyBjQ51pC5p0hrXFmrSF3En679/rjl+vii8FEeeqIi/MSa3
iLKyKFroXp70eF4GSdbFrGmRJYJM28FiaIH9fccYiN42efdmB6U6rlH/nLv7PhZb
RdOzsrrEPUwMvB6VK2yh4yNrXLSJLEzmU6v+WyT+q92iEnzxVCD+rVgW6JfFhMt1
kpqrNLoye3K7u+oz2KBac/Ujr7A1fSQFat3W01uRkcXJb9bO14HyreeIbqEM3O8M
pusXD5epI/j+vhoiZ1JmcQ0MdMexIAWZa+Bg8iEGcExHDeZdVXUmEIOqljn+lBXB
yF76Xz/y+/CEsbY930xC8hcs/emjgnlX7rnjhLPM9SZfCzcvJ4UTV9Imh2pde+Lj
MNRdeY92DQQ8gr8//XzSyLEZ1X68J2kgXOM3dgNmRujtw5saFNZ0zW5i/OgzuRek
KX6IQw/ynk9lwGFF5acMMQ8JrF/u56hi8u/IFHe7No3xWsHBkSBzruYYJ77tvBm3
NHagqUilgejZVykW6ZK62LJ1bwb+4nsIaJ21qS9b/gFa2pDW1KFhIycgpB8wnLZt
8rFBFbuB8jHqxXgArQ+kGZSz9vJQENsZdW+UVf1+7tlo7IHUSaAYSKr2ckqM93AU
H1S8zTBC7T9+UkcQH6qwOdHU2+ZtZK2v38Rb/NwlCLqEQ5MVQsqiNM4JZk/zUTxC
rWer9iz8Wwz5teA755tK98p/fZ+xvTLiTAZsAqGV9mDflr/EDTIJkRGW4kav/ZDC
qJQzSSVlHvpPA765tDnO84PYa0gM2vHhM6iMRR1lVzmL1nEU9T6/CUbMfCAF3qRz
2aXHFR79Ff/5NhIcgkkGWd3VQM6SIZ+u0ugiejzfRH2skXJfHhE3bTGBbW6IX2zD
gMDD0mw0UkE9+CPxOb5PeNG6cHjoOjKfs2yVB35S1AvnM64M7Cpw1hnpuucKriIT
kmkjBh7XdidRjAWphZpGGFUbf33M4hSp5Fiu5n3A7UkWDonVK9I/cGQQmchD2PCS
9M37g2LbJngUNJ+knfvVwHLW3dskrrrm0tSmHiC+slBh71ydb4B+k8ihftZ6enCR
2oCxyGhj+21YhPYfl96hWE/jTzNItg5miDgkjxKQMw0gDdlXJ9dreQZBC27m/FdK
akK4ok/u7GKsIZtdy4L0SVnz69LH2StN2ceFSdta676jrUT86U0ERpFOMwx5ZERJ
k3u6G0QRbzAfFr9VgjJ9DyNoCozUq0fqdpbxhrqCKFdYpuewgCsqdiINJvcaD3rY
HhQcOMqzaGg1qdp21eV3XqvxyU57wgpw3P1FLQms67A0Ykek2HCYftc51rU8AJP3
W/XDIEXq9p+TVFRxZaeySjl/tUo68i4KD4DZxTiMbdVVf7/qNQ+onbrf+sYuHOjX
pJ65gJDgyviW27EY9FKUZgfXk1TD6k0kHpTBLS9uUycI3FlwueudtzZHFzGn0dVz
i6cXvPlfgdQyNUvNbW7/p+olQPli4XaRrvqAcQiXBKNteImOe/3eF2xMdb3U9ZdN
y2jua4YMLuVRogOdZheReodPMLgQxroLvHnYnuLcYMYma3xmdv0iPC0ODIXtSYX6
Kc2E6obKculeYAsejTAxarYrcAT9yRtUwYqO8FzURf6MOj62J2xFiwW8LwFeKJj+
/5tbYZCFWBpHEp/UKZqdHj5WEFWQCYNkdgMi+QO9lFvwfv/stLnf0zVkf8qmlVPp
y0eJts3CrT/JqVuNkP1p6QGbEILr0TOqlHpJEkbtqkOouv+DlnlPHh3btCDgX5r1
2nl7Kx+SFyDaNFcPCooxym2jKJdsasFLYgD78jxQRDWIv6VRyrdNrFr/W0L2wn57
V8Pjk/z9SPygVTg7WXU0N/ejqpLsV53wKDk3A+ATJ6hmgikgkekxvdXTMuUGq/rN
HVYEWKPu8tXwVSFU/Z2x6NGIcHpgBxZQMfAvvogT7JxnDXXcdAOasImyk3zP+TC4
TcM3FyT94ENxx34FxUvsXp72n19sauR8WYHMnu3+YMpnj3GZLfCtVb2bhJKjHAkU
CV8JtfsQyplIWAo2BpW8UU6aqe/C8n2SaZo6rbLzqRxAcDq06d3U/423fxcZ5C9f
TMh6/SaKZBaRMxoojd/rrHcN83dEDaXbMPQB5M1vfHcAObgoWvAkGeepIZpQr4K/
4EeQVaodL/y94UsIPWUoFUpGDkFRZ2BTkom8fWdHAG0V6AzJeorOu5Xxs1kOHHG6
uui5W5V/wmPunxUkhm9S8c8BE38IratOmr+Ct9D/peLBRlKDUq/lWinQ4XvLwRB7
tD/EVFnb9M+9QM0cjgVtt/ZGQ8dGybmDJPRRgfjxaRnIK7Cj1ct4uiZhRejYz9iz
/lO1a/lWY97HKMVaeQ+yysjsxYLjA9F/M9pad5WVKm7S6G6JKWWtnoveer85OUL0
3Mqmo95FIVHjcKz0Rx0KMBWAfH3jepXaA18kLChfk6JIW71F9DOfjpPyzHA/KPdX
DqsWcBfMkhzsbxhMgx/4nSh1BCZu+lwsBEMrh5ddDWITZygj9yrLQ9LeFyvyvTXy
v9CeaqFZ4RQWY4nBuJWudEDwv9HyuYHtJm/B/EpzfTl4mxxle4q91L9EapdTFjV0
l7DQWLRIJzbcu0fmac0bdqnYBzfDFFsi2n9YflSEG6jCi9tU1b+C751sNpifCp7G
/oJ1AcHQYbo3qUcZpbBjGoTvIt3CZF3S0zfX39T0bwdIgFjrxZpl/k9bsthhqmnZ
VWM/00M/tE7QIc3LBjAsFJc5VLEYNwWSvWxbzHvBxXgd+RRAfh8ErEDvuAyhb9Hz
1uJRGs8H24HEHB+vMoCefl6MGXXPq0aNcyqCykGcCYFhwOuJqOqvhkJsm7e9x6Mq
yBYG85n9fRtZH9Hq6JOlDDr41ESBYCJZJJdxevHBjJ7OoZuuBgBl5s8oOep/LBfl
qSfiPdjBmvWBg54EbxSKnG6NcpM8U2qGrd/KjpBPWYu/f4F9Yyqzoxnop1GeEMC5
TE/hqBeHNHmWWxmxX1K4rM28rAJJypH8ZDCkDb2ClM2JPauxskefB3dPYkZE57/b
oBQG4n/SKOs4flqufLA69LHAM6hbb8OcAeHL9gb2Ao7mRX/KYGBCmfAn1gMsq6oP
QbgZTpI9JpUTtD+r2v1lyAoe/9wzwbyE/5XaMXtEtAayeY6IzHdT/K1lwYzPaAZz
3nnXG6tYi1dgPQXN/+KV2AXdCQjFi3dPB9qutf8Wwlgi5KJm36FXYfB9x3efWfGW
Pkiok75rsa78r4FqMLhqWUdrnVjr2GuBT6BIvqYBswIALIcVWYsZq/lHSz4oJdLO
CayU9dV5DZe0/zreqJ1ofTAtteB2vYUlYdeohd0IlwKTltjEi55wmvrzN6+DXQ+e
59qPFQtoDDK2G8DkcSvxbNfHStKYhdZmgkJjMiQxH+y1+k59nyI2rBJJpAvC129S
kkjZyJ1S8vHrXUwwU3C5RVNZ5gGfutZ8APnkBmmyPCtXDdLMDyIJUykCgVBorpv1
tFM/oNMSkOKmR7/4Kcq27UcSUskFY0bzsMH1yNZRtsISDYcAZ11U5eKhwWcVaAIa
u8Lf0oFZbvUyt6bgDlm731Nwm02fuBgh7UCSlOSLw6h6SYTx5s5CFcQpIZWNBBbC
IrpCAHaHzXhuQ8fnDXo6plT9yx0emVLjTVSW/yjwv/yC1jXwQq6T7/hw78qG+hJI
hF9HQ88YU/khDIp5ofcCb9VZIOWaQJAkpYEU9wvZQn6PSrDn2lLVM4Wgvhs2f1l0
oovLSkN3oEL0I3whvpmbJcCZ1RNVlvszVMhrTmZhLyP2QOFQ8zgaJtWCKgZGThHK
YOJC0ThK+4PkZdpECKDMdMikdRMztwVO6eWN/fVRiKPUXNXJcgDH8AffKD649eCj
KalYMvmUgZxc4qlooNh5GczJG0NrOtmV7Ldx5eVsh+fewFLgzFh8XaasdDUxv1BS
qRG/yBp3hzJjal341kO3nj75g9wbogAvqcxdeSOxwPyq7xSgX7L3G7e0WHAMmCkm
T3O81LCktarPratSJce4PnsAJJ5byke7wiDPeBH0ddTbMpApquu4PFhovSvSGD35
Yi/f7iPjv2jUJCyhhCuQbM6YSMaSTaXjkkHZVdTvSaBRcTnLfMgM5xDbT6MdYgno
5P5Roxav/+hImeeNFauauMgUnz3bj1LWy0lu1t8uAWGBJcqflNUwETfimXp7P8Qk
iKxQXqgSvaQ2Pk4kau1uqAqDuKvPhN5axfyE3r1WgYGPAnX6B+JoRZ8L0hJAo/L0
6uXiucmnUphFuGCVZJcHTdZ8Xv9MjD4H6OBgIDzBwZg3e81mEPuRGwKLjxcdVwSQ
BZdfQd0u4Y24ro9M3eewvpHy6HqxEj6zH/TMMqYgzNVQgO6DiGO1vdfCS0GcVc6Q
30iMAOLR4awirKVPhfSW0D9C/MpEWfiK4hRrLP8yq6qkAe6547C7oPFzkDm6tzAN
g8ZnASP8+EII3+/zDh0v9A3h5HVFpk1J3vVccbL2W5/gvXMA2UjQ5lOA0YdUPxP/
lY8aQ7XpaXFrPBUegNENxZTmpQTM64Bw3vrB9FPoBkx8RekEaDCbuMDfDzCafMic
sZ/e5YVuc4bhwRulRgS2q2wGyCoA7rRQdXcxn0yOrMIfogYOoVlNYjGTN7i/Oqyf
FILcc9HF8QJQ6CW3SgZMraTTi5CX1qH48dF9EywvvXro7qJjgaXLmCP0jYpS/Cvv
5WB8+23Amf4Zx0O1SV3XZCemokTlkxrCovyFDaqKUxRqdZ9PWF+hgSEmCfcZczP2
06Iw+ZQ9vHbWY+x3xHeky6U0SQEDvwdYk4pbp555AZqHKQISaT9b+yf/Ap7T7Em7
oxadqYfFRkHVCBvWcHQZYb421laq02zu0Gtc0o6S+lYQlRG2bhcENfGyO3nAnwRT
THvSHuXnBgjbLK8IO7huReprK+77t1Q9or4feKE2a48iTyntZXCAF6gGZjtPplSo
mZacJWxM3yeh/WrtVX8ONn1aPjIHpnI8v1iL0BzlHpm1fZCO3OchzuGfvfmxCgEY
zKBg86p4oV8LcQR9uxAI28HN4DUCD9qaP7w8Rz5loqrVOIFzBnxbsd7K78v0VADn
ZpEK7r9K9EsBhBHehGLASmAXq4VfLll/FiUCuf8EvxeyMFHuePszio1FGtKFd7pm
TiSIIbb+FB/hOlSulJSggxeYKMC/rmohbkQhLLq5EMjwCDc/JOEdQk0ycJ6YZzDB
1s8Ie/HOep7+5zZcWV3VRXMiE9vhmamuX/nmfYi1pDD8KjTyvjtKqWht4ayZ/HTc
gfP++PHTGHvuvhL8WD9TIab8NVVNb3P+dJOs+yp+NSer8l43Va7FtAHvUcyZTD/3
GGOedC/YTOq0nMAcXpsAWpKaOXai+bd2DTz/tX1eG55BDy+uGcQzVfnRpzZilPwO
mr6EP0YFJQ4gykjwm0zqXVj06ico76w73UBzsLy3GXq+pLlBgL66bSS66NhcAZ98
`protect end_protected