`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
YATj3kULTF7Ty4ORuRfFpnT6YIk4rUPRrM74bVTnc4GjdV8oSnW5PtQkMCLOi558
1V+/wvDfc3y0Z8//ksX8sZm3JZWtrxUppw8c14g9Y7owiwp+JumRtO1zuk5xFbe3
0MMnIxxoTKLhyRJtAxElG8sbx8N21OWDGiOk0Xyd5CqAmk9dcOIbxzMjW/wndBXi
maijUdqS+5KiRCM9+Gsp6k/iEAa2LnYTt4WtjkmDD1P5jZKsiMgFck8WOqLymplZ
ml3TTfn1UlLNm/+zD3SFGP0kABAiUT8NK2xBPQ5UzQ6sMFPd/np8iUZ5u4QLTWOZ
hTrU9OSX7lOvRUo8pJ9vPg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="BzW6NOo8eyBw+CxsNNo4wIDxODIsVe0ft0K5tGuSUZw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
DhjJh9S2BY18dG77XPz3hsiSQ73+w0XqfJhD+f+lIDHHVjOB7CfC8ieNRTexgzn1
5W+qoqOEwenoVQtit9u3XViXJSRJ0wfUC5a9axblRNyD2mUbyfH9+f59nWqGkVOh
ieHxkA/DPprM70F3APxk51m7/gNSLICSvbONgLGndWc=
`protect rights_digest_method = "sha256"
`protect end_toolblock="L7NTNW/5Dqy+2kJZXKczEa3js87UJ8H00YWI+92sDHA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36368 )
`protect data_block
6eHODtGLmq6ccbB074dgNWpdzW45i5jL0Nzx5wwM+RA0eeOHXxEV143NNyQGmZjT
bzHAi/6AyRCB4X9z0c4MjyrZE8GF4crbMH4T59xFHqVrQ4zXCea5w0kG5yvHgpKo
Er4+TXTXa9FsGlVtYMafKUtwPO9VIsTKYDTht44OjKOlomCRFRKrrSBibdZ8eU1Y
ajDRt/UQi0jjPY62v/f0UNfqxca2FSfXgFhNQEbtJqJLO6IPT/2jKe2mjAxvcLcj
BBsuWvO7QLk2kLrUcmSQBik8zNp4YL1BWMnN2HC4OtTmIUgXxCgt8bKkzOGNZCUh
IVJ4ZeY6F1xzqMxcRi3K9a3G0PP6rWkf8nky9xYSBzyJRQglkPFSVqliEu/5pIEB
UnAxjOFLeyETYncoy8Gus5rMzxrPrm6ydmmTwyLMwYGfGBhPXsqxgme5hMAPS0Ml
C8o5f1LZ2XIvra7SOPoD4QJt3xKTH4m5agTLe7FDwbCetxg50tt1AmVBXmGIiCYI
Eh9s9sSmiRYif0B2Z7vGgd5Zk4XoMZ7dbh/Um5OaFYbG+73fPP6sFuNDPWyUIQiI
86j4pKQl3ZA3tokM0O2acdPe0GeXg2cAi2z4/bF68Dgb0VMge7Sg4oXSNXBetdJz
XGk9mDqhVF3kPKOlCHvVjnnsKOrmaKuGcxAEKEGnhZV+cUrGpuuCGQ94YUHt9SlC
b104uW9lI/rarsG8TDzLz1IFBKiQNqjAh5doR63NHOiRdQaBLwsIEX3SiJwPpDwv
xnwmai4cs7YMQT1XXdH4Pru0ghqfhVn0UsXWvCsp0tUzc9BE6BGln+jL23XPpfX8
9RXXuHvtpMFzoMWtfUYj2xH1zLhujCoYIvbRjevXvhMRbhmubrlNw2qxmBmNsh8B
Q9SNkvuOIFvgXJa91pF4407T+0Q9FLAkWGpgjMIWRyfkb3n1i9suDRs2XDtAujjg
PYbfAFnofigutJYrxLR9juiTWtdbKvQ8OkYk1TftOw4cWnXniUr1khLjhi2ngLR3
WWPJxU6/T18abDT/C1T90wozWBihZ+j42jzdsgY/Wi93JepJ7j/JbXhimr5MFw42
WxB/jmmxnPpkuAG2AbL1EsWMVBeMQW/n7Mz3opNLpwTdSPqCeYzR0ubcN72pNVv8
m5aRd9yG3jPmn+hHN9Y3t52f7j2j5ivHDf+xzWQUY1wcAvG1QB7OMsR3DUyuLaZX
pSw6S8l8DsWw27ncMyAy1ii2QjjJSOOSf/PVN49Q5Ohi3C7sq9ud81B6YdnQ85AA
3DZUjHOkNOHAEYAialA2gckB0zAljW3A5PA0cjd08sK04Erqivbj336EJzpzn+2s
OCWKBOFemdln1HLePw5NxsArMy+NVyiT/n5BwjKnTFFeLat6cp7ipLXabWhaewhN
GcB9V6O4OCr+Lr7kpC+P+i4+2eN0Rd57YfzonphGeYjtr7qD3N0e5IsBbu1BLG7P
Om5cIMDBEXpnjO2NXJd+m/QT6weBQO8VzBEn/yavZsym1G7Az0ji8nvdFq2RRrTb
UuS6Q4vFnuyNhRKHXyoYnaSHFNZyaOHOYaeIbUsKerN/QnesoRpdw97haVgHYZEu
/OS/IrasEIfo0/xBDPXLQxffvGUNdBntQUiT5kcWzn6jHMRgqn6yanszusCCoqBA
s0X+dKHHocgouX0YxBAT3rYJHPalOGa5V1b1aXG+ybOscXogxo79pfE2HBJON5Zj
nR36f0gx3vlkUa1nLwZFuwwTOo//c0ouiJoP56Sgh2I29jPtZV9jhWo6D1YDGGxM
+vwca1TImk9ckmcfqOI4wUE/LJTng7PuqQpj81sidZE7XKCcX3c5g6iwAlFc3e3f
5wkv6nZ7B3+PVsbsxpsOTM0KzbzVQH2y0xdtiOUm73SgNZH+NcGjvQR6aP6uh9Yd
zHxN0l0WdMHprlEOqe2a22wzSammiMh/UbOQ0vO2HAghdgm/5lrIpfIHsz+dnVEc
KeToXs7D9EGLrUwn9tmh8dnLzjxmlB/Y6UV4y+zox6qRMGuBlWuIhUij3NzrW5jj
WDUvgN+VzFelBuAzkUt8+RpoAlrnVj9TS+BYwEaTLT2LxqPAqgchXUs0hn0TUfeQ
lq/AEOJrM8pjGuA1E6Vfnz+xATJsJKTyBSzhM4ezgrbTDVBlAGAu2106ElCEp5sE
IgBmJRMk1MvBp9NRuisEtFq+FQA0bNt3nj0kwle4X6SxSyyc4jNI51AIhTsBlONc
2Xi5xdcEmun5T2gZdPDASkNjnEgQ36wVDYTNRc7kSN5Gg90DppYcrpR36q49VVFw
Pge0cmCsIUbDUIIGzxkfqDggkTDhvgaOQ5y5+BlpqKIH5kBqg/2/+5+l56BBuRCj
rtRe+fMNwNkmtaXAvFC9vPfIYLqO3MXXRQg6BJrIkbC56y0rKMcah4uAuWXfzTTl
8NvWaRHXU+gpPpYuHwkAyUj2ZKFyXLTbYXxR4uj6RULBGuNvOwVsa3RRyrvJGmP1
Qk8dFmlPBa5IcLs/KVZPnRM3Rxh8rn9ur0bJ3AXlKUTA0BD7UTWjxzY2pDAfKT0E
PboH2hqkGyl2gz10fRtAL359rpm/+g5p3O5b/bgyu0TRT348mhHKg7HH7K10kRql
PbtZIVBYQyoAC13jka+TMZgc62SaefMMNXR0mVj3ppsTrOxL7bxgakOSWUptZsSu
07765bDEJkWyoTRrt8DN6wdj6wDEDVVp+tKHQewVbc7Yhn1UXRwv9qUiqgrQqFIj
tdiSaEbv76pgjj6o21fFM3IWaenXd65Lj07ZNs30SWINLdxgToyjccIofzMq5ME1
s+WhDR+82nO9LMI9zlVgJKzfyaOMIfly0xa/SMFsvOg+d0Shs6ZU917tD4feNykH
dU1j/AnJxuIngxdUms6elCcwYoJKaZ+UpfPgP/Wpvp2E8Z9ydMTQIVQhrgmVP8sd
3jMvJ/dhr1YjiL7l8hCgQDX/UEfUAUYhAfiKobCnjIpMiG5oQuvJjRr6quU7E+nb
hIBlz5ecDMXQ9Rt2dvRfGCTZvG+tpuPFDmy9mDnc+oWuRE56Fl4W0asiojUBk3rw
WmIhb91T702SV8rFjDFtefsuyL8lXwUo9jMibQJvfI9+AjPhrugFrXg2smTI2dxk
40TPSvymVocwz/FB9bosvVABgyW41f7rlWn7fOg1AGc23o0/IRoXABCNcq7ZUleQ
+Ni4B9la7N4XNWONDcJSNZ7FVFqrcFDdXDUaoQPwkT6byD9tK974D+u/u6S6oq4l
daOpTk2qLJuNnQTvJnxr0lW14Sp8uWeZtOaHlZBdfNRIvu8s1AbNUKj87aXCbj1k
apfdIrKmi9wUQ0w1HTTs3AJCHSg019q4/DFNzh2BEDGFQfkwdxQoHkWGNNrbswSU
j9DlRvPS7OJD6iMLtudAf82Zp5JxKelI5FBYGlJaLR+gqUmxYiDiGuq+r0rSvf3u
JkAeyY3DfrtYsjzxArYAnxWP5jQbUylYpbXBWIMTkPe+vqIXnGDfZQ0c9jwLDKqD
QR7Vh+z6rXJpdW2/vRH027ClAQ3ynArDF1Pj75XUvQ/zuS1iaDLdafO2QGrIWFpu
icJhEJXZLV2eTsZ6uJovquIoX1xOTdTUsS9Gm/WURAt/zrNJI2yIAq3e7bXRMHKf
VvUo9DnjjXESltyMoaEsKZE8y6RHNzUV5buhqFlkBj61kv4/+O7wPDsRf/IZLcX+
+rP13+uZeGbr8lm/Ysm+0L3xec3ewFDN73PS9217jQXWVdmlJGFYMlgGM3UxPf5H
pLrCUl+1rDH13M5rgArQ/sllaz6utGFjDTzWN346V5zI7O50tcuLqZ3wQoYGubPl
TYbv38FSYP6taBFutiZvCi3hx6aoQh+c3aPe7UbIlH3v//0aFX/61kJLHWP/tJdM
jmBP8mieIgvBDZjwzWRNCyW0icxs+ypmO6HAVTXJX7uNDw0zc6fwWUy/sgJIDzoQ
HvXaYWvRbS+ms6FTW6Xs7MGi75PoZ+FS43+P2GRkxSQm0NbkLHrMS4XwshIA328V
Ej7exAysihJw0X0baZD8pAND6T2Yqtts6f9XjKh9UUzvcKZcx9FP3Nsg1gu8SlHy
fWhxc7Oe/8J45hsIzNwFonNZRhBmb4GW6uiYbXXuNL03A2s+r8mt9GHIRu6mOobl
A6bNWiLCNhlFYx+Xfkwook3SlszJSI+uXOLW/xSuqUJKDaWu64nggiPZlrtaKu22
2qeK4G7DxTjmijHEsECT3kSwgA3rVfD9xGOs2I3iY6vR2cbjESbtYFNTtgkVVU/c
3iJkmowblUPo9n1COtaY+7EK5Fce7XI57ZRq4N461XgsOHpRX03rkHyl39rbZRJN
9nD58c4yRxvyLpL2r55RrXIBY2zolLkFLQ7Ii33BfNE+x2h40tFvpQHKCoQ2TSv+
5rHGtmqVuRBqZrZHuHHsvgyUkMjINqQ67wMGAJEf8NsnnjSaYZnR8gHgtm6JAum8
zvgc8MmeNtBImoNM4/9b+dNkMvMK+zH6g8t9hTlaa/w/jTDvjnbMb5sGmoNwasSA
xHUOVayYSpmBQwHv4og+/rrjFnidL7AT7U/S7HVcJjm1NvLFgKz6sqaM9eY1z9y/
dozwiehDvxOi2GZtVpL8fHPkCzkN0Y7EyZaIS8yiG3z/nJEgf73yfDbbv+bmdbWg
RpaVzzCTWPTQKJpIvyKRF8dwYPzXvh0Fi2Im6cUervUJKtSlf9AoOmEjvMNtSiOO
UB72afsd2x7kuh+owlO7+ttuiGcA+RieV/e0EXPTZVkfoKCco7EeT5NaK48NaKc4
TyPRUf0Zhw8USy5KEsILF3kNiTHfbFZgorrHVSzXGHafgrOmBnY8iYM8trHpXT/+
mux0LDU8VzRK9WGYi/cuTfqUkakPHXMwiJwzwjqPx0LUyfVsV0ip3C7aUfkGwvHI
u5z5ISzKrSFN8CAZSH2IDnAFDMkqWQMANxWJ6X6fh22MHnfw8cb14s/pLt22H86V
HonbQO6Xav7uoEqm8n48YtaEoqfZAt1xjEP1FRmCHKJUyK70vebmbBv5w4z+7zEj
zvWb6MAmdbP1QDFGNW5fRCD6U+p9YIz6lZvgPyaIjJ5bREWOwb18IlF0DZKmaK1e
jxUc7LLYB8ErahfCDcCupOszoDGxX8jyoHsmLIx+jHXN0otSaLAOlKxQjNFTJsD4
MnuCbYnlS0NCSquPRps0Ql2nxxcuAAvsX0Duw5UOA9GWdlm5gU6RmWIDCnWTEG87
S4WfAAxPvA8bGJN9J7nEnbc/pw1jiA9CJdNbmJKUm3ionKQskuhf0OmInxo/P2x2
BANWTeuszlGaNJhz5BTUn7swVvH+fq1caUGTlZfjPYzUV0nxUE64Qfoo+O7Q2TWP
+srK1yqAyf6m+Dseqqil5ZnGJHqHm6sS5qm1xeOwAu0yS5somnkbqbpPUTN+/IPz
4JE1ciFt/SFAKclTgT4HqB7P+7Cm9SlPIq1Ab1QQexnueW3koTmdpqUYIdJJECzI
ybTNe8mngxO4QZ6fuSZOl2kDow4F/vSUi824PpDB2FBfATxBLYdn3z01gOKOb1fn
PufRqV/ZP2UqAtsMTdnsJMtvda71y3TCz2noX7hoa1Q7xQLl86K5OWMmTuCf5wpV
WZhR5Vxa022M2LhZzSA5cHA/qdZEZKWRE7i+C9f1vD6Gg2/a+tUS1SAr+604+lzh
ke0wuUaEOFqA+QSHcLPExfTXXMpi6XhzCHJuM8UQt/AGB5g2DkbHf13aOSOztwuD
4WZYt8phFTbX0j84mqP6IMgYhBo49ONrolO0p/mzP8sBy+ll2QDK8vowda7PwRiJ
d2mhaXuDnidAWnWsyrjXLp5AGSv9oT2zbvc2lJzjpIDiS4HvkKpN9dPnEau1i97G
c8Da0aDkK2nywYKcq52w5xkCdkC7n+Tzu+6RCmCjoMqOYEuUEhyUK1pGY2W02pCx
NXwEVgrrtwdIn14cQ5gkYVr/kifzwvJvpoG++89qBaoeHMw4hKHNV6xWjcR8/UQr
i+wEOY/9WSPf1RaICkNjWmRzO84D1vVCgFr5N1lFfGcrgVT/RAdU9wsqXqvCWm6K
r63Uq8Ch/1PRw8DY9sQU99cgAHFUjBxwNNJ6re4dGbwkx2jC3fhhZWL563iqJW8g
It/oXwDKqunZOW0PHACMYRfSJOTKzXQmFa6Efxu8pe6xC7VyhnCMt8U95FYirXHB
pS6t+P6lUj9/P+1UhgKnvxdf+pchjZ9oUS2OPgwzlSjEmHqvR292IJhYqNZ1OqpH
jKMsc262sWSpdhJGi5SaHQuCIE1lzTQx7XphYBMZDZBosxRmliss/UYbhFVm1KXA
at1iCaJOZJkKS2sGKHixuWB7GlX+plHhrjuij4lydXHu8VMJOuUssnkZk6wnZf+5
wFpQX6kXhpYQ1nUOQTLRXEgLgzoKzWLo4u5Ix4IUqb1LXChEzVJ+zeULldJp/tuf
EkLRd4KeRDvU6zou5/mdXxbae4QDhymqzUs5oVoeEvwBMNOIrhlfLvWbletoZMSR
wpfTa7SgFkR4zG/iuOhHTZ8EKqpPQ6SNOwwn3rjhaKJtF6o4abg+SUT5LoOjynS2
6EisyENXSzd8qmTmq29uVmQDchghUrqzOqAuUEdaXD4h1mLogN/7lgm/S7pKvzIR
sIF3aM0iRJAKoapM9WZbSNXHIGnnQBXXOSpQZ29TC7Kfpom7LtYcweVLTOnoproo
lUIcxjjl0hQqSCedwCiqAVV3SiOPV/NhT88zw4dwzyWPsywkqt9PjCXIaahrnfzM
1zv0i8fwpD2CRqGOGk1OxfckDK+XCExO95yJkthu1krE0yvHo5lKy4v7/sHvyRcT
qAmbESbuHehbcTw4f68/D41eHJoLFerqhV/tlRtlgE3IZYSEQO/CdydXpwlpZdJr
sWyAz6u17NvhNV+SUiCtGNHRA9NHQabY2en7ZEUOEe2MQWAmuT1I/YipOC2Kq0o5
MzeSTo+xQ85kBUZGXVa6SwjqI5c8WNUYjOqWjsbx76KmvhkO0HSVyukvEPDID7VQ
rTx8/DjQB+R2iK86u+TYnBHXplQWyYcoItWnoC0YLnLj56ZAn9MsxEX6zXs7DGNs
fPRFwyIXuJkiVFx3xOeB1mhffOT/DKmq96uRZ7DyW+WpAEFAAIwAf3RZfIqD1rLM
PnPHTy8Iuo3qvo3w4QZs+NgVUVYH9sCR9FwnNLt9Z+7PhS45fHfyWsJe33uL4Dy+
xVJbNsosV58ZpRXlgUeiARtV6EnJ9hdvwjx6TcZvpacb2IuxvTy5tR5E71WFmtJ4
QpCKpIto/xLw2xU9qJ+wfW6wp3lg4zwTPUtIvCm8JhjsS4p0JI4grYBvCeVhyp6R
hF+kzN1WHnnIcspcFwmOjVWknrC7w/HXk1InU+xPG+tp9p9hQp7LWqaqaLJlFhFw
Jv+iXQqf0TMui7cmahAup7jCaf9orB3GQoIRQCioldh2qbIt0umg+PmbsDauLqqt
SJMVAupB0f3bXWnnlR4Co3Agk6/5jYP89eqAF7Ree7aZXQ5FZ9HCrbUOkIfi1Fr0
+OMuMosguiyv7DPh1EYtzxh+YNRArxLxYMyUjtS3G46pqrBaZiOkYk5v4Ulm3lGU
l0pmBzJu4AlXLEa0TXf/9Ae+gjBoPGjrR1OxnOJSX8jzn26SZthcAuBKDQ8vummj
7eeJsEhEU8tvuDof+O30X2YJQVWiOSVl8jyry4h9IXgp7sdecJpYk3zIzswh7/zQ
d3zz3k+c6krC/axSZK+ve8AZd4AmZqwYxRbO3Z13T3LGXmSPQ0WjIIYl7KWebbDI
1kdCjJPsoogNT5Vee6XUI/UK0CGC5V7g1pW1gnqY5sla2dbEsSle1lgHzdo9MDug
YVsa3b9uRV0t9cp7BSB5IFYDS7ir+hD/edoCC20u58b1mxaim5CEZ6FUAVR/KRQc
XDP5s356kW6tvbgUTl0TVpVTvpwag+ogfbzygYuNckNFJs2p7xGed/vUhrRperwz
jD+CxDdsuXyY8vV0U9rpQgSqffvZnq0ej3eNpsf8HR/cNbLXGja1063Hi6LK1urE
1dLXzOgWFSiqgDyoFaT+vUhgMj9Ze0EkXGnoHKERvs8OXobkc24S9VY33CvBDJOW
P1vOi7is8d2+PZdau7H9m1i+8N5wV8UrvfqiHNLjl8FwEd4U9MzgA6wuueE2ic2B
JgTBEYpuuCDC4FFHJjVXkuR0/hnG8SsuIwG/QIHyx5Bs57iIoIJI+AbOcIb73hTa
EDbRnXNXHSbZrT5bOxSHIm70N/6m8Nc4N1qZq03xCIMe+OYOn1k9ljUOOMMM1Rlk
i+QyiGQJYn//a+IAH3lMN/tb/YggGdbR01XKamsaGruC0k6c+DhYnutQmT4YKkVy
anZ/Cqahnj1Kqq/jTCgPfrNCZyNChm6bwZGg9o7LTNLxCnkjC2e2HgmuazyoW7d5
awBouPyhu3fKB1A8wseq9TeW+tLqyZX7ICCY15fAHQc1IkL/Ib5RrgWoalvUU1GN
1KYX6l+r8DxILLeQ+ePbzMIqtKLJeeSSheBOirx2cezNZMOmAoYdHKjbE/4gzhEQ
qAV5Dv9STcm7mR+HvSdIYbOdq2oAjyWwNr1A0KVHViylG0zUxBowaNMi037kVjUK
BIjVzJbxpctElvh0kt21vGQRuveH88bIk0ZZajnvlAPxUOBkAk8jHL79Gl+Y5Px7
LDU+rbyHyBqN1fSIpbxI4lZ9ELW0+5aQKk4IXWYCm+EgjoipMMarbyASvmaIYmfp
fekxjN8/6Cpbf639ohZ1DAnAQrpAaPI8FqnvWgTRjxG1LdZHwAJNvfgC58jNC37F
gD8RbUVP0MdoLMEka81dsDsExvqN0oSm/gNjKY++J5z8UHyMKddK562THCr2LlgC
abWlJu9cq4dcTvbPC74VlzBffT+2XzhIr4ThPevLGutuVj08YLgWGQcs3SknJFMa
uN8jq31kl70h+wKQa6WMyqFMwna5OpoSAVS504QIenQsldNT1D0Be6126zm48rT9
3sKnbReJQBAajTWyc1wLYz88rLGrC23Q+rhy96UR+n2lkUc9K4Q9FKLPLQYH2OSK
bxr99Y0adiD2pPzeGCbXVOfEBS12CIi+ZS+nmrb4NEDXmgKNkcmGEJlwi317ysc/
XTJWeI4GhUurWsta5kpXS7+7k4AK8F1KYCEJ8+0UkmzM+r1L5/c6tApgkPr+pUNG
c3gi7/P7na4i7d3yJtyCgnOhGBrm6xcVNIN0ff1k5qMAedtKQLRBUecF1+gl2E9i
D3LHz4nzUpV4QU1YcTlOmTS8ZHhZoyN9rhEUi8kF18TQGuZSoqh58NOyK2oliGeK
jEA8Zu+OYu1KVmGCUnSct7eG/2B/EpXjBGsX4++AnnQM4QyHSWs4T7U6R4d5FS+5
Nks0a1dRo76lsxPRi+0pgZ9JAA7vqWrWuhXrYG7WfT9yC4jnDQxsPpGMGxJyYvca
IRcDxWikO2rRKlrhom84XdKli82s0e0qK2TO39OqBg1RaonHbQjkSl7RUjBgRJli
jaMmjUOtoKeZCLQVx/wdJLuaDavyGbZm/HENIok13YdJvhYpCzrbMbvexBJVAOO/
3QfEy7GKqvKyEisyqRcH1+NMCKpaCX08bl3zt7B0kVHFVVcFbnEaLuYWQjGHmwOf
oNvoV/IhIoYjdvzTjwiHRARCvuYiXXL2nsNvHo94cxk2kKQsfpj1EdFHwWd93gml
NPFGHZvVBVfbyBSZk4UFc/VkBlxfnIDh2/Ua9kyPWJ9ZpuPgq9siDfU/QWB0C5W7
xmucjryfEXo867ykRTs96ele94kTgesnYF06daakQwpAnVT4nwhboq7MSoV4f6lq
31RRN6UO6U8A29HIQieeovZN7c4tReMUOAW7KffzJWJfc+bRXLd5Ws2+d430wSIR
pUlNrTgedB9whNfgNqhAalyXR738sGLWkUHgN1+zpHYQGDbASPNz+7xeAK6l5HW7
ZLV/iyftVd3MmRGRbcxYN0hadTN3n6LGBT5ghhUduQiQ+tV8it3qhvS9gOfTw/Ub
wJ1Lz1Fgo9DMa1mvb//zjiH1b3j8fLGEIpa3iZ7reRemA/G3sIGVZNaIU1Rnw4px
/KBWiMgVa1ezPJgRpPg7iZUhzU4/HScEnitBFPI1elhBcBjUbROaR8nL6NwywtuD
0L2muNNpEqakGa6Vc8lBi0PdHfqAvwbjzmSmTnOjDu6vxGWnatGdG2hsqkrA5+jc
wJwAhzUwpvswNhDiteIuwRK/GuEXUbNkoKp5qz5KLEDNDZb8F7nwjwJ85GG1WqG3
XfdLzBgZnh2YHDGVbMrociDFwKlg6w1OspTs7dvRvx25STw4f30Oq0M/cEwN/Qtg
ngZdqRpCZf1cb0ZSwGRFcw/Gs7swgX3YsMEqauvHY+rUzwUXFoCCoQ2kKv92ATQu
c3X57ZR+gnK9eWVerVlG3erGTsuMpry/jFlw1TbJp0GR/R7oUQ8V92Ci5QVN7elh
ZbUrFySahFbcIqGk676wGlllA0tQhSXrRjFpHlAe+gmP1oA3MA82qijJgjyAfMJw
9YB1cX8UzE6bUokIzxTeyB63KskQeqsRNN6+GiKpcYez2R20Bry58TpgYrajvkoi
JphFITT1pYY7APdDwPW9QK9aZIDvJtUtRCfDRV/Bac+vL69X0rA4W7BoXqB1jSrW
0ykEdlzIgM91tWuQzT7hXmlCHnKSeSAxSVSYCHkfg3QBhexZ3SdXl/o/J13DvRtb
EQJ5UqZ2wXYmln6BQJWoFedM0+k8dUtDFBzlSzVkG8bCSjGUl4+eutXa1lcDueel
91rUxSTvEP7G46cZGzMQLtb2CFFWmVhUHSotOQ/xrQYGCHnW0HSiOlApOEqTYJwJ
53L9rgiXuFCpHhCOMY2JkCWI4lojoxLQ7o1JkSz/4vm/oK7i8qhiQ8lCLmhbpQLl
qBPqRAgD8Kwe+snMFQ0+pPSWUu51WQ8T1mwUt5PopkIAG63FAZzlR6EEZeCX4izj
fdLV+lFcthlPze0PL5x8iGA7Tnq/2Oo/VVoFI/U1S/ZDltirX4rAstXkRo6G4yw2
rgnpuy2Fz9RUeWC1EMKfsougJjYnkH2NxUltDLCD61lA6q6gQPAz/Dg49usoqaVk
ZRlnhfuscQJyG4O+r9KEd9WP5lSfYeO+0Jj4sLcvxErTrg5VR6jDWrffzFGe/BtO
A9fuSlbFiGaayQrm9+w9q+h6DsuP1cb8MYdS8UWYWz9rknchXwajJ0CtwYsYgdWk
DnUTj5yXPXZORHdE9ViKV421sne4cMUDMrvwkS/9XdwWVtoanfzUsa6S31Cgj7QW
RmWN7yKfRpMHo0sd+04JxSwBEjsawuAQ3zay7NjpYitYD5mgnurvmL7c20myMCVU
2pFNROx9YTtid4IBuBOFuTrWBUNKcvK5OPNvSp49LpZWGdoc3JI41uTwZa+Ck5Fd
4Zg5ZidOtyb28fWerCT5ewLEIve9+3wu8f8lwAIHNMC4gl8lVX3as847wA8z8zAA
okUpcYxmWf04QzEGSaNk2e6rA7QOV/iTLd/ASixCp0vgQNNhWlj5tjSRPbYxqbdR
GS2JRW1WgyEK6iaUHoMSB6YuZH8JhPcNIQZTIUIGDk+xWPALZ3E8vskAi9PK7nm+
GoS4l/gS6ES+yZinal2fGUoOv+C7DjOEN32hKwaM44EVeq6JPwqMVPH7RCX9feoK
ToLEC2ffUZoy1w7FiG6hFL1teHR+CacSHU7PqpnSmiD00xvsBycuP9s6lYcYgewk
lr4w12V94nJR9Xli+T5HDI8XgnEXUlXHIUqDLjOczgfDCEW4TtoYkfZ3Jzotzen9
5uBoIggiG4bKIIL7PZNmSOtgXlwthURED0btRtvavkWTId5ti1PJbuHg3ZjXBF6a
bIDCEah3mHLRVvxnMkRiRg9MlJUkPhb4IIPQIbYhnrJKkGiO7zynQa/SPGGKERW0
2DXIeI8iKCcXbuG8MzjczajIVXtAIZmmfTsXUDuk7Yeftlq+DMPMz3Blf0tcaCGY
zCOpNTAfUDfBIoIhYCn+g/RrTKILRcv/dC6YZfQ9qCfWUHuuyPFRxJbFjbXv3Vrg
+xV+/do8iuR1Ft2J31V7Pk59oscn75/IIzB6gYDEFna/n6kP5ibbi4Ye/zdvX1v8
E44FtzjpjCcgMq3OHMlPk0TfEI4ZXvulhJt8ChdQX+k4h38bi+WLjkub0j0O3JZM
Iqu5Fd9JFzKg+/2j3fcEBhsOtSD9/nBScopSGxT4/b+7xHpzt9QzEiR4ZV9q4FyT
0gF1skRgB5pjm7nW7jS+t6qtCQXExAWGHctS2vmx80n8mhREpVO1t9BnY9UhVuF6
M7JiNSkTM/f2kMfa2UdY5I8QFLmlBV1pY5lYlWz5c8JMBKVZSLZbPQ6GTR4o794R
gu8vjdDRgtIppC1PhnrLTYaL8QgFeDhA2V3ujAZqwMmEKtSPYYjlnCL1sWX4vw0Y
OWP7TJ552e5aHunvCErDaBZC4yG42jBurrgG64eJ4nj4TX2jtq/ynwttrRqTSfNS
XKR4k0ES1l4Jt+ZQ94dQNughluqcUe0dOmwEK7LBVzYG+q8TVRRvr9toxs9Wkh26
wXo4OPenZx1DVnyuzymQGDBwWpMUZVlc7olg1G9ibgBHFm6LV5yLwPTp7ZH/iutN
wAkTqwfhYak3cAT2ugVhJ/Qnh06Ehx0N0pdXjU+N8HBs1gvdqAuaqUVpgLsaVdQ1
rgqssHtlF5qNvwiIzHgCb/kLt2JTmMZH+btpBon6pTSyepF1WHwiOV837stn8Azx
NgxHqIgyucCMeUseR0SadxQBg2r0C4LQ03up0gUS/t/eP7+cv+QlRhLiVKzGOnHi
nO+N4dUO2f26kEvjxILooRP54K7l5CHaGk+hBp6NVRQOUXosGNrHMZA7WgS6REho
XIhdO+BIhNxJjC39ndLggHTY1KFPIvveOAvztV5wgKazpadg6O2pbkub4fN9Dutx
f4EHMW1HNjW2ECaimbhmty2IMz0Hdpal1CVPZUUPOG/TpeEFQzCUKZ06/22PErbC
OPwU99sfbutMA0+YIZz3xq9vn6Atp53/Uk79N1b+wA6AtRsybwcRu1GMFzWrjaKy
AkGm09uv6wsxULxKvuzX+xtUUK/qJrK9CPw85lgiQ38LfycmRuka2q9+RdncRwbi
VIAP1/ZLF+cuiggiqc954fmvVcYXeKFZAe9rhr5OOWuF2vuowF+E9edSkw/Ofd4t
+SSD43E5rat5SUyngilroJN0gmUB6x2IehCVhJpfcKp6KRyHtsDVmUU0ceM3DoeD
biPENIev2NKcBfHUsUyotl9L79cveSiJxgYxihYiIEuIS2pLoesjRLDBQXdK7KoK
Cahps7z75IeWGG2p5sxPTviDiOREpIqBkeD5evcxqqr9M4rg0Avu4BsmFsXXerR+
RVbWkUc7/j8kCZ+SSTz0kBud3DpUX5575WTlGId9mrnfoZ4jD9ORw9Wx8XLU/zSx
OiEP8RP58NNFdn9Mm7mZPnLLe4PB/pMqzD+BiC0YS87xHgYI2Elg5fNVOfHapIVM
rjCy4Qu+0GTUsRz8j4NXcIAefGJgtUiI4jLiaZ4nfvfUyxphN0NLR10jhVDIpJ0t
VfC2cchnvvPUYcLNFn7UfoyfBAPPViBgH3j0GGOd539ruHgnyKfRfA0OvNwx4sBO
f20rV7PSltjmN24rLKhnIRAF2LWPdGm9IJJgROnfhcSZwSwhMg5kAALQVLEJxkBm
mSIgOf2YfU3TPUDeX34aF24cVMFPz4vInLWC0RZYvx9nTC2xRfXaL8BAnNWLIvwo
kdf2rPT8xsRA15CyrQTmrC++qS6DxAaQzy6ePjv9KYRaJolUKIkbmmvSKYXcVLxc
G87g8oozGtowJ+1hjY5MoizudZ6u+onsGVUHPZJOEh06znJkb5NdGJXxJu6GzH3S
G2XataivQOyV7WeHLbn3GnsAoaZyUDoL2DIsnoE/usCoaJ4yCDIo+n12IEyHRlsL
WRAN+oSVWJquneoeA94RNByggJkSDPNbAtdrbzLw5wML7DzUnZUpxaTZ88iIWchI
VE37O2DnFaSYq4zhjSLgRRRPW0Anj5L9Bp39Uo6cQWlfOdtJ3rXpNdpnmd2LgNn6
v32ueAAUDcnTzES+m+AS0CLi6geuspR4vX4OcHId79XFo4XYA4pI8+PSmzlR248G
i8UyGdyz6iVD421xg32NhI2Tdxt/gIJngFlfF9QgroHa+uvh0DNxQq6DFEYTpOsM
vucf1Ui9Lr+xeqwtinW5HVPjYdmTxyhAcmZWzHoCGTX2z/jNjSPjYZKoHGiiUFwM
cHbImJWN+muXK7UiNfC0um881GMf/zbriEcMKDIinbQVytfT0r3QjBpcHCdzr9iw
ZsSxfbrGePCC4SA3MKBogG/0SSKXNT0C1kZ76je6xPBvtGNlMzdbMrtALHKMdpaV
IDy9tlJAAzFOFfZizg4M92OIj0C9Cf+SS5bEjpwJPLu0vIDtMwviCZHDjS3bfnBA
GKOY2bPVOBrNp+sPX66jKdAvj7CNaIrBCQYZ2rXorDowO1BfhrJl4gjFoikwkfdq
D/e+V4qeLErbt/e7cFpXI+Fa4QwNREAgtutNsQC3vJK6Ao6rwvv5gCGa8D5NurUK
tcgwdviu83+9AhCFhIn7FRZnjOLXuWNaTKrSSvBK/1RtMpHQlloCnE2rkrjufrsN
3a+FXRs84VINeOczSuro18ns7mqVV4r4D1d+B/F01cU0o2+d7Chg3JVH8HEkSwkJ
Llc1EMkoWktk6jJHC2S7tDQTTLqwZuThsWZNzG5tbY8d0vnE+40QKC+PC8q6FTVR
oJMH17Rsh3pD9AkYDKDggASm6f8ta43FH8fZQr3rrsH4q/1E46GE7DiT0kUzQ45C
usfr8FFL30n6725VrqolPP4r6Wvwfxe0+gIuKj4/opAqrduiBA0DKDKzbH4itPua
JPS1QnHyrxLxK6mDqme/lvzypeBfoIZIRB7RxQKMIv3iNtfZGZySFYDT4/i49NwW
KtAUvs+Y+tdieCFxGFHcRa124JGaLT6arBnFjQ/hVHXXWXtAmRxahjWsoTBNgJTz
TwuNufStaIScibs37X1rVgFlRMg3r0vk4t8DOKMtnk4rLHW6xKkyAPAPNsBqG4Kt
U7/7tRnYIb9nL+yKtcgTTkXnpy7QOCNNOXOO7ONn7HmZQaCUPWQuaf3T//M2DLAj
KcCwfkA9HXfDDa6OVT32Dqz8zsPnvtlSa3v87tlqCoxFUddB9LMYFn5u0dCA01QD
sPjUDaTRc5y6wSpUcsvX34dfhH/02oClDfpz/HBMMaecGjIyHKlwxGRYv43GLShc
v8/ZYsi/MNC6uMp7Ie0/coXsoraX7WPcq/vzYHbmY8QBsirucdY4k6q5nn6BYDx0
YWt5m/2cdpKcEKdx0TeNGe9gpt4jI89+HOz9gMd2UOp8eUHnX5MTQ9qqMv1N49Fz
VziWwz50OUY2NSZXltljc6KpSa8qYujf6EqTVevTe33bu4KvvwKZPLXBYS4r6rHs
XOgCwiC2P9fWLM3fg8ts9Ue/7bEDa8SLkgPpmliBnS7zuQ8pGZVtVJKk9myftZqz
2bHDW6IpL1Fj/JnzxsNTRFRPSqySjnzZ5O+iqX6uZVbN0aKGG22cVvgyO7SVGAaO
x0GdnFPlZYzp7dOs9HVPw//JaTzBsNRY2erDNOcr7EiQKE3cSrDpf5lsTxitZFVd
avckBS35ZaTeYSqAQAYyvRMN66AGKA+rUtnQBt1q37wr04sy2M4lygvAVLzofudY
Fy9GXDzHIy/lJf1KECa245HuQrpswEva1nVKNNiByRmnTPedE34WeufMzC9X7nGU
CgA8TqbmQmAu3TFdVJlamThAC8F5qjjgpedOYL/RPzYa4JEPKOE6ZszffTokMugE
zgFvIGBPbGN6mj7KlGHwU7VWOyGPQwDHpXFIpuUPOE1t2f9mnI8zzqw9X/UJxO8G
OfgxJvD9RKCP+UVGjvLqXhDlkFTWSb+x0aAS2i/abr1wDEwrr8+l5RGABUlIitqr
bWsIvZE3gcLli0tmO27CtwYg1Em3j/xn1QLvCnXXOpBnOpB4MXSVRz3N8BRuF9I3
D8JSxifFhNfSdTsy7V31Zw/3WNvW5Xxhz1V+hi9JapaODi1ztggG7t1Zp1Qii1rR
9jcmlaCOGLJ0UZOY152VCm6zpr8o20yG5mMGgCwHd4RPSFzE20W+y/cDR11+V3/s
//dgKxqVVVBmb0GMqE2/RSRwEybOcUrvWBXjrsIUMV1B1HatEVnmmCEXvciE240C
hKhevHcfRw8iHeGcbAkwkqJnGEdRhwq8CIGgeU4oI+NnJu/oEzN1Iei4E/NQ1FQ+
fPdK1gZ+mrBehWo87W4xGGPci+uue8cVJk9q4n+P1iiXi1+P3mITNMKAxe/wzl3m
2V1892BuwEaPOJnMALWmOlPDtYLvDMwS/Pp2CYLCmSDwhoYKx8iCpoq62+b6U3ic
YcmX5SmcwVKyeIacCos/IhbAN6gpCGa1vFipdluovd76eVL06jfeAgGA8LF0GCRs
mcl3E/B06yItB7YGY2MyNYbjA7EXGE3VdixkZ3ojaqd2dl2p+IwubL4fVbIZgTpM
538NX5FOC5T46nIIJ4gmQCNm4jmdGHDpbYty5LGmPyEm9ndfqtJY0joYet9Ls2AP
I8NGutCO1kLJnlj7xdINSV/vCBuUvKg9c3Hskfv04ez5q0j0U3OT9sZzu4R0qEA4
U980R9wtPQaot0ZF/PgU2UVCVyNUSRHKgJIYjQvaic88MfRMDSOrYtkxIH6qdSQs
qV2J79PiS18RROAfrrm0K73HcQz0//Bm9BCoGkNet4DJnB7xFUfN3JkCmi5aQtY3
NJ6bcQrXRpz0+kUtJPeue98G1C0PDpf45XWchK8RZUDFZlSl4deuEK+6jk7xa80i
yitr8eKbBSW2CjBRynSGVhtyP0l2Uqaqor6gZ00t3AorG3nZbHpAzt20tEBy6cbw
frFvvINzo7v7xrIet/n9lUqw2ErSdoyHfFU/O9DVXcWNNio71tytURMlqc1J5Q/F
mz/7YQA/LOi+TBG0N/zNdUgDpFZxauTR5sSRyiVDEraaLxUv8rDpA+CuxUZAszyU
7zeWs/psm0WxArwf/e4WjSVO/mG4A834QSp8QjfGjkaCbvcsAkmCDxwHIRaCNkbY
B8SD4oWH+GLyj80Sf5pElS11chO0VgJNas2LaqEf3MYleXBt/AfddiL4dAOdyvJH
m8/ppkf8uH7qGvbthKQgBKwqwyyARej/YnuOpdOqc0VpKXoeMII4pybQ0e/GHza0
CTPK78qegaImLO0zXvnuoxQd16Ekepuq/3MiRAiYdpEJDZHwXHNw6h/ZhtgAGfaQ
+jquSyzXfqXm06SZzTDL995HlKN/AlYt2Sxxicy/zBM4nyTSgxVeXSIOC9kXLUbQ
2rmDKeWZ61r7uXIwtxNkFuVLxxlPSqWfAmzmwK5zSSojwTkyhkrjXOBOB2VWgnkD
3My9P6T1mQwEe8z46TXvshHXwBjApEt/pqccVlSdyGoYwuDxybzsf/S6euczVqpX
PLU+ZHrVGQUKTcChjhk2qrAXK0z3/lNGYZ/yfsofP5pbxZ+Vyhm6B4tEQ6NpDLJd
ZjK13hvMsG4r4B5syygQ0D09P5CBgD6SkpLOeXu6021lBHBUpFmokDmkfg3cKBp9
D3BFhNYikPQKi9Utsl8/uE8eGwcmG80Kzgd2/bUf1kjkJSTxfsRVxHVD2wtoo3hf
DQej5Os/bNjIVXobUNVokdeJ0+tHLigPFMZXQ+GjA6RdC1YYy7x66qQEjAwCmF8A
DAI9oLDZztHB2BK2K94GFa2OaT8xPfc4Sw8yue5GMyGdemrYlfRXNg0Bl6oePU+i
bDh0VGxhfrH7O7brlOBmkc4tKnmLnF/2EQv7Lc3HzH8CUw3MBjrJve1KZFRNPJ78
EEOmhpDauUUMVV4e+PQwn61bXiCzwWcHR+AGrAkAn7LS89OGPXv39WowMpV9gm7f
VdA+W3r5KiOMjxKvTTzFojER3jumgugb02SaOLvXT/KSGAzJClqJBUXHweiy3hQb
/bv1bVDoQzHHRflcOnnt6+eMU0m2reZHoJ4iRwD5YmBFNcCO4H4PTHNMbgD1LnKH
CIGD22AsOroTtsl9gbyxZum0r8HEU1W+xlCK64V9yTMZx9lWx86MtxgHI+w6pnJu
pYxM+BBNpLP+LD9/O7N4HDwmEddVMNDkwcUzKCL5htJAdY4UOIFPjF9H0sGnGCuy
58DhXcUz33v8dwAh24az9YMRcB555kducKKB9GNJ6Jx+gnyuTX/6Wx8fU+tAxqwJ
wSavvfcbeh6pVUxJe8QI2Sdes4kwN4mkq0g6hOqRoASQZbZ8EHXaUFNMy1JKWdvs
wwnNC2rumviZuKhD09LwRhDn7+5EQ78J+X8/n5YsOlm+RoI+vsPf89chyN3JQe3p
Qrjt8OkOziCUxa0n/cAycbGJP9uuhnkhgl6qO/Uq11CN7jZ2Lqw7zXPuKtDxUxxJ
48aoi5AV/0xc0FXygj/CTQwxPgJJ4z8XiKZJom4Yns9XCXArTMa+cR3qj3Fl31WK
GAfkE9mEzi6JqnNggYlvBRPmb/aDkeQPiYZuFNJRbUGdHeHOT26gi/fimbjCwTcA
mifNI9hTLa3DdFe693Vld6JZCBCAGuYNhgcMoNKuk2fnA/YcjtTbRpPEL+FSAlNC
e8m7btAfV2NL1XWRuXRKGgvIrIrrxZhAAoBU98bD5mIc7bLaKknvAZo0mPINynuY
QHfvX3yUruEvNGOS9s1ylGJSB+wnva1cDwX8zFK23lf8MkPZbJtI3WAf/syaPV4l
Ol3y6bU8ZME72AhurzafKqG4BS87Y3+/i0VAuyJx2/xNynqvaM0N0kr8S2Lc12nz
4//QyTHALqw4XT3OI3RqEY2bn1PH93mCgdQXWiU7V2DrnP4EMS6tnc0UdGnmnF+B
8MVzMnb2wMGOM+EGZ9s72vtepM06gbhXiv7AhB3s0fJhr3KDuDHK8XYREbbRmFpp
9ta1wcUE3kLDEk8yMTk6/MB3RkmgXTf98KLDr77D4hRRPxVOLVox48WKOdedqhIp
DhyC7L435nN3pGnc8Otce0QcY/nIMFWwEbJCTk2HyHn6fonM40DODqEBb4+ifqXm
S0c/2AIMPnwgYFozUnqoL17xXWDxGlqXCWG4sZcvtXsuyb1qee/I4PblSXvsNN/j
rACq+pJIvyhB02e8JydOz3htRY79tSyS9TkQZnv6UukPfZOE0Ac45w9KlHEo6bcE
9ckXxIHfevxsZxqlx7Yt6TmECIqYqma4+avSIBsFJDUYijLGrKbUnnd32MYx84bU
oIJMgCtuenpPbKDquDt56u1cu1LI7YTrJDYR7AQRsiJRDpmMfhOAcqQh/Akirsun
lg/E/qMkhg8HFDrkkjWQo6MKg0CbMpz2uqFsQmSJ+2WqU9C/crgbSRmY7JyeBlv5
HNVRiNn+20ch3//b1dmSrVPrrVVN7jS3i23IAj2rjvMkcL5w1XRfseMLYlqJcNEO
0mhyVEusuwCAV1iBgKEUntsvu6/pp0dnS40AVOVV9zzmT3zBToqJCWe5AiIjf3jN
rQjkJ+qNaGWUUEbzD1nKmKja/aj38wUzHqhAUWwoK0WSHP3XpfOhyCdcvN3vGSrz
B6J0QCK55+SLMQaAiy/aGdSV7wVCbiNzyhgaB18G25yteKPbOdkqj7A438S1WZ5M
5I32uMxuO/75yEn5w4Dj6pxd/pDPeItklb1hkqClrZmwHpVcRIwNa98LwB3voalO
NX2kVuSAWC+kKwHMR3fjl5yz6uFeIOZK0C9p/hI3ZnwjRTXt0wrHgu0ynOLvilbU
Cn2F7rq5e0v+eWc9gCdvK/7lXmhP8kZOroehVhtr/D79lfpGL1y4QDrcylbNRCh3
UQ48xRZwZpYutfB92ZeJFmfh3KegIvbpOJdpHgtXEH8GCzpLsqP13ajITSTISP5w
vJ7lJ4CUN4xzxOU2iS0kUvwXMz+2sFWUTwKaJ+l5ozgd48rTQ3opRut+aZRwPwS1
6+s4ZfIp3tf2iftYcn4YjLpqFXedzu6/8gk+0F7ueJKZ/YZxfvcz5DG/NL6Hkqx2
sZ0xnU7SxWbfRi51hiYwmFrXsObaDI2rYeJ/gvPdjOyyzDulvZ/LszBONvpwmEiq
ayDfTbNQu7VRXK9alSxMuvrftctzYlklpJlmK7KHIfVYk0lwQW0drsPxJiyOn8VC
N/nkUXuuF32UN/f0kMIOi+b89+PBl2K8UFk1d1778FySdzk3nYiJMo6ws8Di3UFf
SH0VEe/KDBbQJ4rA69CafjoSAOqwmRmNyCHOpr7wC8B8pBrWTvabqx7gWGU8IlUV
QbADzSl5dbxte2Kjje2bRBRaFp4Ne8sdiuL2/ZkESWl8rz7BYpgY9RzCILoVcoNV
4bvepuAuVFTkKTIGmepLYFyuTtRknpGFOJCWn1KCdNZiVZDDronVbOHOKJbHu9/9
K7fP2CKg4kjlb2r5iE09k7PkEolQkng00DYgJqWiw8WT1HmmrnJdh48akZB+e2rC
DMdl5T4WWML9RLqq7WzOVl3BNzSAkFROrXK0E/G0ZrpLyrqSE3zHPGTN/SIrXF9X
ybLIL+8BTF2SgPTcijL4fWuaXPjBisvv8T2dBbGwhcxqRdzS/veo0mKntTe3nrGY
fgmdP87jJPMe4NaRWy7LnHCZd2aRZE9d2d5pLuIq1laQVcFCIBsyGg95xHOjSwMG
bse67gJJ1c68291goW6M592UwUvPhMEdqpq8HTSMXp1yBBQyztvysNGvHUvKt8w4
GBCad87UVqEPGLab9E6287Ix+/GdgjievG+k8aa+p9uADk8twVg4pkvIsukVuLAu
ZsUG+Txkd+chJ/5TSjTDECNIChokQjPf+dj08u/dBxThAnH9rDY8YZnuyhtKVZmH
tuQF01oqgbbTkWrbG25St0W8M6Dpm2UQbpvRy9WH0gSb6d1hXgtcRzBgYQY4TMRJ
qf/A17pShU0T6HwCs6AjSfBwkxpz7wE5QfUPUjZxf9yySRblqo5la3t8d+PmrTIQ
aks+SDYGg3MU4Q7A2WwDkkE6U4k4uLQshc3yXrI60m0CtdLnJURDuoHb77T1iKFH
sME4OXQRZVf2ZP+uIwkzYzeOD+Y6n1pIVyTxwOzFVQiZS9s7cIdzkyGI57G4IhCl
F11SRp+cE5hyr3nw90hkNq+uFTP4FX6FhZH8D09U8yEuLTsPBCkrbh22GHYK4Okl
kj3QLePV5NpUWH/B7kUSr/Y3Z00DZutyvLGrLKu0n1Yv8075W4ebtMUAj+/vFX5B
odtpj4LMtnGBu2HgdYmqlwnqkzxTLcuxtWb2zUIHjXHQhv48NJVjro9Pch+VM9BT
sCLDY6kHx3/Ma6Z4yL87aBRM6fgyt65owEerM8Y73vSIL7g5057MZK6W/GGjk9sx
mwLnHmHCeqYhdqGzUSkV543paYHgJYsPW4FvSDiGcGx0rb5uJp9pDTT0NFaf9/24
ZAwWKU1A0BpydkmcC2rTUclWwAcy2yjado8LhLUe2JlW2YQ86kbvMYlfd0H61faz
460+w7BA1U6YXvaMtZnlbgY6Jbe9e38QZNtp04W8klkG76ZSnELOjQs56SRg1OW4
Vo80BFZHKD6FapHAC1Dg1w6B5jpvxr7XKv762lvZ4DVw2fIyWh6FIbzG7s+CTbCz
wn+RRATzmXobl05+Otck5tx+TAmf3VrYoABe0EFYtQ0TDt+hOZoBn5e+kJNCZQVz
/IEPFHYAocz6UKzbbCQC6vmj+6/bdn/AaXh1yMdrR6mK/AjOptw0f1ohtG7lQNc9
9lLbVEvO/HEebve0Axp7eF7bSzXgL+ZZtd4Pfcq+A8/8taEgS2uLi/etsD9+tbEY
jpQiyinl+jbvDKaC25FG28B13t27LSmPS8DEop9F9jG4ohHzRqxRyiD/qTiGQu/N
RU3npOHQOg/np/5O3tgsmciU/rW6dkKT24/aUrajSe2kNr4E0P8SSBmQr5+WBFrh
aAk7+U4wYM0Gz76RvHRqrAqfBrnG4FsclPqO9Fnx3MgmFWyqJL7FfEdtPvzydVNG
DpmvflzZ6Jt7TE4vfNIcRbRzYHnDOCk7+zlSNDOeOvawR0lvcWSWC15bDyjt9JA6
H1223I341s/OxZj9ZdI8d6jdwpR29zHPv8vfbwGYoyN7usdcoSKZDA1Ngm9PGuht
zKDLub6iz5+fjgX5KAKxmCk2vc1/GaqL4scHp6ya3rWfDANov1Nyq6zkP9pXoh68
2zj8W4U2sM3p14RtcB00bdQ3yRoF0k9IMQmTheR5J4IfxDjLSIa4TjAaicNDRkRk
jPD+rZ/RxwF12g7V+wsJeSsJFF1G/6d7bKgxtDXDk2l3bFVrwEXZIEDPK7LpfC5m
EUn7fRiGYVANTFCi/G3bzqJIjcEpv3HxYGtAudIgd5ugvB+WenjQitI4XQBFQZ3n
eI8H0WyQEpF86zSujkuZDNVXZWd63HZtShPhYaGKmMwEzT3Db7ozJSttSo412oUk
tiZRthBnySt2mMz72doxjfKjKJGuWxMecEC34CIwpLypAW/6z66ACITbuAjxUa74
NheF1Sh8yRg5p73JsNrdOBGhk/y4q/aBGPANZ5Iedmom5uxKnpa5H7Rr6cOb7XkO
l3uhpAcUXy/HeUhZfT5oFXLgriuPnnIK6aDQeBOK84lymFQ+rd+6tlKWfYKJa6rS
rZtAA8h3Lr1p3KccKXt5TEPoRYbGs+4O3onZaZDyGbBkF7kFje97nMYFZqPm6zyt
tPq4bLQuwV7hLTq+fq7oakcNqWjX4NDQLpjIRMsHdinaJT1KILRfKQCdmUXtqyX+
BP8Yp+XNrkYvrjkk8f2J1hEaa+yO0Gyozrn48Ppb0GhvFekEN5GIy63PqlxOAfHp
1ylqHMrrrcow2tMjIyCgvdER05o5+Cr6vbXqYBSgDIsM5SvwGou0EPTBpEpDvhiE
zz1jVpArgz2pAMZfOdxllScaHCmvKIQLmnve4Wrl6IdnzH+jLH/Pl6blerA5EXik
zAXB6aWACSiFQOMFH2LEaMw/821Zpu8T1BWK4FunlyVDWbK80JzGITfVODsa7DbH
SqrbKaafAlq++tlX4bd7Pf2UlIUVMIkbdic3sU26XCJFnkHKgdx12SJ2HfNLnPS4
LXobz0EfzEQmDCNnixx6mqKNH1WYeE2kkkxXWD+NbFNr/qBQtEeb0fmSz+4x2/XK
GVZc3rBAxi2taaW9Xyp/GfClU7gtLVJMqMFLV0u/EGJfHm/pW57ZNmRvlGSUIbJ6
bbozTlCHWHDNUAVrwcstI9DQloYUknyNX5zoLt2770uUkiCcPBqZFsIN5PJtjDMo
7r/suLaWkttrmTsoBO+n9M0UhUnGIgKmw8jLCy32hWwEgWEdLufGGSG391clWY22
0Pa9QjEoXDmH/SpdxDhOFBxyecvKicTSSahtstcyA2Oz7G56eZYDg/W2OzaIzLK3
qZF+PKTRMMzgxUuTgU2K4GI67ZPkvBfmXiV1Q8hgJ+4vwTkqD1bJszlPZFEHErS6
YBV3mXFTbJ0QR1G8CukEyIqbpQPADtbnrQRP62J1YHD2ofDVF9jduUPDFSqhI8R6
V/YMRQqotmmzbAY5RMsd9zm+xAZGb7sbS1stfTvxsJk9bCpYLnSUGaGq0xeXVH+Q
hDwQq3nxjwrTo95Wv0fGK6MyADnhZ/dIQQbxXGsGigGuPeJunAo64vIJV0XkPyQC
uPFMgf/lQJQOfWMJS7CcTqMdqYE4EjBXt+lMhSKQmXo582AXidIu2wl84nC9G3xO
gSCyATuqkx3NFh6FRuuW35ESAcyHlrwR79d3x2pzU1w8xn9RfpkPTcIG7En8p1L+
1Wj9VVq7s5JmAdSG3WFzEPdrMhv1WatiJuhw16sfnzUScgwwVigY0msRNOoW4nS1
dKXXve4uScnaGt6Uefu8g5ndhdXqdbr2LhfRHjFsN5rHLa67I9+QDFE2z3UFJBcD
PEsO/qIIz1dHULP0blKhoJW1FkmSahOhehH7/+JQn9sWOVlMA3CzJc9063OmyLzE
Wy5jhUk9Ydn4y/F4lUS5ubEu8LlmZdM0QoLTUCGNlVZlr/Usyr1GxqMT5exy5tbm
l8s/WDG1DVGVpjgKHno1MMB8D5YTc4rnpw7lGAbvpfpHBxLvfKyGduJKlx5LtrXP
OsDT4CNAW00v6bULXwdrqjrgSysCD8boQUGbgOdpdVOTS9FFBc2slT8lE7k+JqG2
Q3LRLXt8jWBwRNCJFY1Hq1sOPkeXBzHhlDlHtFnAX7hcRDgr1+PRaBYDO8L/noTe
9fKn48kwL0XUn56jHQ3nVftWpqL3YDEbqQHhYcV9yCjGnSheBUQKusx+ELPBKYmn
muA/tqcv34ogM5FmwuiI31ize+7ATk6i83lON3Z3FjKtuubFiTW/8y2t2yoQzGbm
Um3PW/grzb57Gbpjo2Hu0B3D7n0aLJhL4ue+ZwtAzssc5LS38IKvW9FSp69SVuBD
0HXj/yYqaBIL5cEio2M4yN71U9BKwjb+ulQhWickMsZ7E9R+iA3ww3eUcdRFElBg
ldkl1G2nnixuD90ZXT0Uu6F9ECPscEWq11U4h6wf7xh24wxviBdOs7sWFS83CV8h
YTlr14MHEhrtv1k2eYZdueTs5t/7Ka6BavZdO7NOwe7B0f8UfvJ62M3s3bpa6kV+
3aYig1svfX1ICanC4b6Xe4RCKXFybWx1VlC0wMEZACKrvHNQvTR+hUZ9i06fQBAQ
ywOkC/6vtmQKZu55hlHYqFtywQefM43SAcp/7ozSVoa6Ts2/S9VtMO9FYrtiHB0s
XP6fl3U80AAPsmnXcCSGOW96xeoRZCq0VWT6+vH2UlRAFbJCkyREZq1POHIh1xPP
qiI4XQoMduCq4HrCj3qCGN8qlj1l4+Nl+PlEhsLC1ebESnevevkye7S/BVBkyeAT
2JhXBqmk26lOcMcnVeLOCDndD1KEnznTs4pr2V1hO1lJFGSBz+UCL1ikv7Dzol1D
8/suRj6r4/EzwI296C7NUwbVb4FOuraPs9YsAZDwsRJTsnrwJixgCHGNskUPp75z
D6d6Lr21kzVSGspLSslsOWOaU1A2RZDpVT8weXwrN9sMhpq07WDJrpNwQ8R86ARz
+wfa6txq8kDlyyVeQWsVDm2Wy3RZoXru5Nuhs0Aa0/lG25PKkzD3rGUgUWS/OLl2
N/uxt7SKpAMnaZyo0GCtMX382jzoDZXhmZ+gIl7lgyDUJqsbs4OeTvcX6UA/btiq
jkcs3+6XYUZL+bJlU8FdXIEhRYi5KsdC1sBA4jGhJvokjT0ipP2iaRMYPPsesOtz
mYiQxTGcNXPQTmaYWHWspK5Y68Q9dUGs/MKw2YE7lh7HUoMEPj2AbdTIqZ7acNKe
AZLOFGUyiNN4k28JZA0L+RIfpGeVag0K7N6wn8W7O950UUvNPV1gdpocO2UFuB2U
xUmCDu/kZj9xDYZTx5tq6Ax1wBq4VwBzg5gO6VKZ1QF05dqpSF6ygYmUCz8AEwtx
HP2N0TWQuqdEm8idAyMwyiO90spHK0uqQixoRk4RiZdxNulUdxiFvxuJEm2aQafH
t5DzQjOEFQHfaGhhN0DljQK+wTLdZ/V/ZuLayeeJjazzp6JB7HiyTTKdYI5+jgt/
eCeUwhaBjWLxyRSIIvYwHWM/g+R5UFsVIzPe6O/NKQCedJz/XZYqB3DjtKgRoV06
7gqFG8WU0nOQLaHXcoKxL7TNAsQE2DcWmN8zhnXhUgkdSUAsvUhHd7d714EfWfPv
W07h0NDzjEBs/je3b1giaycnsFBVPgiMPAgBvIsRGYAeB/IV7FH6tSPm7+7liugD
Af7y9lufiCO4Jsu+gcMuVKjR/17yKr0ImLDas3ajgkan7e89Ql/4HqehOzZ2dpMf
PXzHjJ2C5JBDf7prAkAw+7/tj5oDleMsAxrZirXltQg3mWTdJzEiw/YMooiGSTzd
TwXUTaDZG+pefPlNO1RVyHd7JGSsx+EPScXCu22QoUbf9NLConKZi9iJze9g00S6
yOO6TsulXzYbFrzfyTO/y/F9CryCkwLCPguA2+f4IOrIA5cR3i1wWqjpb5R8tkS3
74lzDL9UpDDYNZE2WlQElr44FtewigpPEDSzhCDgd9VXAbe6qEVHPCazlPbzAai4
7xLDRUsPhCzNh5ySWLIiIZi2hy39377gvofFr/+ERdb6KQLhwUIQ8QbFTVdZ2nvF
3dQNW69huM4Ce+RKPGYTedaraL4uqVm0rjRush3vZXf/gMxU9w+ed0Kewd4ViMRW
lq0HVYKnMVdPZMi8vSaObGdo10DVD9Z0OmanFHmvA2kUYiEgVIqGnhMWY0BMJrt4
ILOQIP5/+EE52PojSZM+fMg0OZxA9ovJwDsE62Mlgo4jP5lxR4/cKOZyvalBq2ZE
qEPh/xUl914y3yymEgIr4UjCMgjqqfLCso14fp3UL25zxY0/g5Iz3WL/sGfQ4Vin
2XvIcoEcwTN5aUVYJ395CEd0G21guJCzJ/FmlWCKR9lqUEJiP17DkD/IbFFcwgiM
/1mYC4/8NMHSkaNJz96OukWlsjVbAq6yZmPdrt1sb/Vmv/gDGVZ3dgvVVsis+0l3
WBymea9lcJav4KscmvZkbVjNILW4LekQMgtlW/Ehkl8tr/JuO/OjxTT1Ly8UKCYL
mPa4TP/D4Q6qkkEyspb4MG5jMS44lIlaMFa8qV6K+P9OT7TL7MgbXuVACawf5QiI
/f/eJf5f8D1klVTOraj41DNNiK+DE7ZPxJLUGPoS1MDg1cr/pqccrvf0PMyjLuHi
JEi30g8qx+C7c5lQ9L8ca24Yk6Qf8v2g1UcUxxY19jlxJ/gI97Wo5a8yxNlKyuqw
pZRfP3ZgJSZh02TSZyUFrUoQAO0/vrF1UTih9gemu4VpYNuFqp/48Dya6A0vs0uk
G0YM7wwigJUuGckskquzepeYpmsW3nyAKnHtdlWUyUoVRskWFthspQMTu51KtzEO
eujukz39K+lRzAHCKmuPMf5zgopYfCwzeebDyJm/VF1dKxWalpqJMJGpli7/BoJy
qS6ujGcOZb3vCLrdV4SXQtluMv9RQjco7Ftbm7maTCf5HtqX1C3/pmO9e43fsIsz
fB+JrS8n1uG7FMm/L754xBI6f94rsN200rWT/MS1co1fHDsFTRa+wpQP7HSkgU87
Ex2Zf6hCfBCWsuxQHc1YjmcMot2RwPMEfA/nY35w1aAMwlXRShhgazq96n65QQR7
L5sIEuyrNJXc18CkgB/fucY65RZI2mGipoWOXqUSlDxU/F/bwX/nhaMRTjBQLOy5
iLn5f87ccgp8sZvltgOmEsw3JAuigcpwuapLULCgkPZlxMLEXbl+l3v3YIrqYuNz
5TsgZ4AFZSGB9vSqeMWGbOsdX3vqsq0AdMXS98UTUAOzzMLalrJtGidzNKnGdqwY
MMEryDM0yL/iOiSZmE5uAByFgNvAspnKdVtDTR9O8eTB2q7E4b3LOaZDZh2qlauA
P40s0D5smw0BYxXO5jorLjsuFM9ZYZqsXCQ5G+wN9LiHa1gLjZBp+Q0eV4iC6MzT
Tt7UleKjXna94Jl7RW4djNuFAIhHf3WEXrJLim4DRx/1H6zx4igbPGEj2czEI4f4
kQiFY3AzqSMDd0WEvHd2mmqdkjr9GHToOQntSuujGfUXhIDvU02KKyw3FTk1cBdl
yA4PRRo/9rJo5R6XST4h53Zg09zfCVrXJCa67gbYbl5elst7ByRdgIxrLPeO4G4U
yJ1rh8eeoXDYydsOTcymcwamd8Yqzz8eIgCEGapPJgCHlPR2sxlp1ATD75xt0pYT
ZlGM7DeJTFYN8NpLTdFRBHJ5QiqeGNpEJdAKtjyiXoxtbOTxVO62KB99HfjyNjXJ
CgeAUpii+XjB10p1gzZh00Egi3nEv3DKln2ENZf0KZPH8zvHU9VrY4yiI8TSJR96
vme/w5oEzCuFAEGw56itoertE9behC7Cn0oOZN7jBilBsis1xK3lZdMAsUtFZ86t
iZpYkV6yN5UkimRn5Vk6fcM5bs4T4JO8cTUeIJDxlSOUmAd3Jkvnlp71WauRuJbM
lQ9CKeDdapZ3qIwrb6+Wlzz3fKxy0x/in9DDFZ+C3538tVdoRxclzYTxScruB7Zu
F0toUj0a8d5EomhqFdk+Ojx0yKbuxwnd7f0NArHz0BobwG/vpzSZxAnN4ibdnQzU
w55KVwci2AAwcXHWC9KvoOgK//oZRX0BohfmGT0sOF+r0VEeIbcMSQ4XgPzzlR/5
to5ISzS+VQ9Ast2h/g2Wcjc9Ae8OnyIDqurmhJb+enI2oAJbgj9Xt4cILuT0EAFT
eePxipNPRhbR3GDaRLdy8GcRLgNRKrHOa8Y1UsS2j4tdzg0XcJoIwZzNP5nT1iW4
NP+TWtYjBLhEWS7voOshS3Aar/lLfC3wfxSsOviFUTTZXB6dGXcnETgmWSWUXZKb
S57ezaW0P5famOGg731XsegKGxLz5OdnBFF+TARYjuva6hMIpuUwBaFNPvLT36qZ
qtRBB0m3lgXVjannG1PlBtYeCESNjYGxpkMpMzW355HkSA1muh7U7hvqWdOchN2x
T9t5AKmNcAYYGVF40/tpXke3jMa/0yGgywth0SH5HPyNESgATsbkc2UF7F5jEgb0
fHsiqvA4K+KuEOoKVTQ8956CWVU0gGz9mZIqxmsiNzdTZCVesLgXsnT6PvfYecfq
AS3nir3bjJBd3ABZ+IYeUtaUzHDCVoEOzln9BO0YbeIP5YXnRqgCpPXljLIsTLdq
xdM5paPriHlSQ5OxpJxBXpyFkZ3AwmwajDxvOYYntGbHeMd45uQwoD/NOo18mb+r
k1XPUUn1PVAjbSFSfFzNukK/ym4snDxVhNbpbkCktaP12cIDj5XWZsuAoY5MgJOU
1C/yV+wUORJNDp1L+zZ3MUfG7jjWCEiZJCEEHczTj/znUyS3wNdty72XBb6a94GN
5/bTX+RIEW/5uvnPafwxOD+vCS7WOq8rwRlT8//ebdtFsyIZsZq89Dg6k0aDPzkt
HBIj9cTmpXPMgtKC/6nKdaOl06OAfs3DLGzdPkfqUgx0+sRLbGMQE9XMAuK5WQGG
U3fPSpkTa1kWeQDvICr9M6BcRexfOBCpO8wYSXJBGGaH2CmrpF5Fp3SRCqZ/GEb9
BE5dLaxdOChl7MpDHxss295BJriG1/wwWOsVCeESmLnHPl1o38uYEXVwa3iutrqh
3vrgJMPpE3cA127xOqzyLGu+rMG5PyNAjO44493R+vcBXqhmUG7Xz3RPN9EHvIgM
7tM5R4hpjA4Du0RhiRjAiPr1zVnru2pGSA+nO1Kx2Si/X3jOMVsASbGqspbjzKQx
FXARmDhq4lLHhwM+U7epLIvi0op5s/wiIcy7ZQDWcdv0/e4P0Xv375xfhg0uVZA5
sZu2xxADgmCDD/vLASoV1xx8W7YnjSRUf3SDCWeaNXO8fmfnwNKrqwSgW2MQxCBH
/G7gD1hE30TnKBvEifBxK0EPWM3TGPsXOS4HBzWlXBmKXvrK540IJNPSTTmMLMXr
hieY7mp5lexPpEJ4TJr7n903lrUkMOtAv8m0gDwnIEXojE9Cox1UwfTwQrv0vJkq
WhTgvdN/K5GjzvrE8yFgSgVsu4ONO8Woxt5QvxBkNPGEY3Icy4AaIMZ8EtsXRZ8C
vX4IStzaDzWUKaX2coBErxyAPald2hwY7F+URoEmuhfmPXziLAn/YmuWQyGlm74I
JSwM9tpO8K5GjoSAHqFrEIyTdZyfGE8WCh3hqwK7z5RxwFzRSeapqZ/F1xOLV5mt
/YdzSg+dWw+d36lQt2oqAhk0Zcy0MxlwPrM52DcEqU1gtT29CDuASlfrVjyvESSY
q7uhDKz7b5YKqU4CTdMnwDV4wCmMGW0m2F6S28JrJZB8IjBlAebt8kI1wXhZwFeu
uhMSd3YIQY32xQTm+LCoQ4R1Li8fYvm2DQJYHRIvV9lsoqsG9UdF8B1030CwWkBW
mc5qgiIXNVxCFNgg683gfiKQsQZjTJESydKgdDRGksPamZz0QsJj1xWPzsYrOLvR
RZhyObKoCYeLVLZwGWYV4RhiWGk+DpoFZYP9VEomUDLTc+71JBmieio6TlxOxEk0
NuvQvaZwfn7/GCKSxMJCZqWFo8L8GUEz/JsDpX8EuK6qfnAkdluxAuBbCx/JeOXD
PXyhrAoZh5WkJfvYJABG1zOkRSpKXRSvYjSg5TzHKjjLjB5PiJZlrdO9ZRDbLRCu
womidPdpyvIuIdl0NJ0nDqU0VBYnK1bfCaMyUT9PwqovRAf0ursYjgbxO8kirO4p
qMXVlTS5+g9vAwNQUXUk7n5fq+GVQnYrqz1ZwpUXJAZalU4midoiaKYoRgjhBNFb
n3jYPFsMTUv4cbuwE4x8y9+LJFBcbFtNVSZoI6POYGIDFuvjC7ygcgyeOg0qrdjQ
FAGhBz25Y7/PYYFaWWowL04J2vFImwninvTlcmdfJCCJ2j2r9FFzHn53TRaiCIKB
bGnkvzVLzmR9ZLWWFJpmOSEzflykL7JasyjNubnTq+gZ918qRqeMtz+rilGrGzDO
80Y5FNwvzlia9lfe1EHu0KFkrlaCQHlDDvxbPmCWE4ptNu+9tbdO0WyDIYTBNmm2
VFcXTRHg0LKMvh68RVZ2AK1ZZiVSHPF2HmJTDYCf8ZWeQbvwsM6GLKVHkVSUFgC2
ppDd7SVhuFddzXOXAvuNZw8FgC49u+IeTnNf8or4HWIwHVy3zAyH9eNGAiTIEUw2
dHx4vvumvtgk4eOouy+XDQ2O0W8XCHE64KcoqyByFTQNSyIXdXiIuwlDHtkzpZno
kPla8faXB6WMzm1Fi+30wO3HSPw+RsvOq6eoVzbNkzyWY3UvOhrTY6Vz5DCktT93
BPr7SPbncx2Jp9QNYZa6e4BW4ZiASnERMOQDntkVYJQ4DlJiveRGhqpTjN71CzAs
IbYWwnfdP3n1oGKtrnmPZKhIC4v5QGSk0StIeCNggTi3mrSOU+DJVjnNhm43TUlx
0QdpAPfoF++/TvzuvX2MGWEmvuF/2RUZnPdfAoxqJXzptDb8yx91KhfKqa0d82Wh
vrR/PKeHWQBGcRVU0rMonqQ6F2hIXg8qCm4dsepHbqUvPxzBms+EJUSSm36RSFs4
p6dRDz6GW+t0h08WdNdW9E62D4eDP2Gv3RHMAeY8yZyddKuY79VUm7l1eyT4T4gT
4nUfi5yd2P1F9Gx01mfRio8N3PHdb64qCtB03/4c5dTK8b4fhWOwwfrlXpp4CXrY
WjCWaYqEVeYGE6/geMthaCFfqn49yA60GztV/f3X+XYYga3vIESKDUBIVel5HB6C
q/p3VeCSO+6u6wb42Bq7HPdAV9xw7GG/NsP0i9oKeQzmCSCExaXzeucX5YLF8nGs
DUQLnQENDztglWmEwKrDsMm6s8lT6naU9Az1WPb5Yi44htbFvtTQOVQ2oOr5SNgz
CDAwrdDVYy+259jMj/+XTxieoaM4q4kAsmDZSvuv/25VZeOJln/u571BQxM4T3Rc
Yxze/5MhM300ci7vqTNIumpWgAIv2Oi+82hfhVIoP2QPa/jKyaLm1hDaEVeeXUJp
XobpcfqD0P+zO0xjZmhLjuLW0BEFW00WkoI0C6yBrXurOMVMS4WIsfCzPMZdvat3
L3g1ZWtZtC++S/F5uzPgoJi7HGscE8aVrCFni8O4uOVN1ia1u4GlawJh/I5tElLU
nGVSU24CScC8Hb0GlXxQZsYDPp6wl46AOIhWvit7jYq57NV0IM+zowSpoCpAL/aG
QANXr7yhxidz1z/hO1Qj5RbC0v2m98uvBsht+8/XoSoMoQqMXmTtoESKCQvTWfUb
h76Vv8boD0Ocmy0DDEwzc1BUjMqVCXzbxaGFytKp2LeFTn24HZ5zveErR3FbkODG
T5oOS5c6D9rTYxr2CViPtFN5RIPQvpro2Q+cAwnMVw4qYqSbu4Ej1sTcrEgS081/
AZBayJ43Zsf7fzBfUa6KYl4VqkbekN08ukRTkpSKbD9YOATUHBuHu8sJb8//Lm5Y
R1g/UI+0kz+KF2CsL6+onCM4mBrOPEYpP2xpaN/AmQuEcbxABv6B+zq2SlCK+8be
Astw4P3lim4AOzVhW3W2OLL2heOTrYCfZ1cWf/yWdc88W77HCE25jg6ddOelXT7A
9Y+V1QNqoryPyZcAFSl0ytaoSjUPVgpTqEliC614A6p212+/CN4Rq27IbA7Lo8lJ
u76JAqr5Tx0JpcM4nYcifbuBGLcdQ1UrzBbN3o7USVCmIb4jCsZbkDQ0gXBmjb3e
7Qgs21SqmZJy9JmAYruWlYW+nsFAshA+wPPnFBjGsY0oDY4XWG/wuh7DV7RCl41R
M+NDFR3U74/IbKp5VQeNoUlmBVodAoDnLXpu8whh6rX4GliFTeSeBeIE9VVhQalk
NNWuNEIy6/szDp9Oguzd5wz9BrZf+D79zXSqEME6IHaPUxZ+a0G02DokDEsh1Gms
pLsx8NYkfAKy7DWAxALUu2iyVge+DKnc9mZwE2mixGf9vmE4xrXynVcEFTbjtecf
1QbKZ0QAuet0yOlu3HHxSWKbgNkzkMyWrUmYqvkFnzhomEKh5QEPWsT+u7j7Frwo
mWxRM4EriA6HD5tPGF6vgL0m3rD74G/nF7+nP6Zj2lnje6fAlHiDHXtN6vgr2UP6
O2m/60MkHlXUK+GXXkdjThpqyi2I6QHIYBc9DeyGv76IofMb7C7czRy/tUPEbryp
IBycRoaGLtewshU89ENUqKG6mIC2aUHmx7YMI1Qr7sw+W+gV7JRkdhV2J5Ri1WgI
i55BoqZOA36+7vNZdVC49ZIeVm0JWFoXH+LvynhUk9/Nfa0A7jh5R/pSLV8kSxa8
TUw7adwv7eNPvMKeNL6cBUgL0DpQTqa9n0c0tLcpH8kv5m3fhkh/DWB9tIzRV0tw
sicBozU1s5mzW9S3QUU2p+K5J4tLjgLl4XA/lyqL5/IkBbFaEVwhHD4uZYXkXjiN
Fo81wCSd+ea2fkRpveJod4N1A02mEnlsZS/lSHhKLWyuleGdFP2SGr3nFBvMVZ6r
28/KiO88ARIqwd4vK2JoVMs4UyVgnPASzTXeadc/oloXexpUKgcV5PUEo3tuA9qY
S+Jf4urjsQII38zV1gd/DC6fnWYFI2r6kfTeNfDqZV5DAdA771/gpcHYaZn1ZZi0
QlyUUxLu/wJQxD6Z2F10kx/dRWDN+MUwiorjyrpoiDMJoCPMX4kNvmudIOoGVQa7
wHuCLY/2tzvCrlxzH1TGNDZ9tWT4xfun+lAK2eBp7aTHbq/Hh3owWu2JCwfqb4k+
BcYy72qR594L3MijV987oHv8z7Tm3uObhx1v44bhxempjj6yF1n4hAhXqGJnL1kb
61E+/D1qppfwk8s9lDPMzyw5+4Omiapbmr2bWPrXnbxFuVHl+Vg9uYvVHklhW0R6
3R0J2dsGOBoGWVZbmpbizfBKlCYF/xp2dlRqq3AfobdUrB1v6tlPFPyCqMpgNJf4
Rvo/kxu7t4kyoUTHsywueZi6Bky6yAmj+0MIjvviSLQyg48gTtzdB21SHOQcHRzz
V+Lf7e8q86elE0kmNAz12Z3YE0WyRevDjA2n+EdFUfO0lC3JvJk4ryy9ZwKUJVDX
soktiqu1W9pfWmUoy+qPwoHly3ChZ2jVRfYOh4Iwq7aGP+7cImzrFzoxA+Ziwl/z
czW3C77/89IAoLyAZ62/fjFzr4Ow2TAawOhGGKVHgI9mxevc3k06T66LlG6ugacG
ILDDsu4cYB+vEs4Sm+WVqOkmqhQsCAx5H9S2G8CkEotpfl0jASL04V7YsZ4hv4fh
UolIk4BkT2kGokUgpube/z7XukUSFrXjWtpNMMmRtX1CZTjznheC2xYftvHJnci2
TX9ZyKs/cxBEv+S+nScIfbYKbls6fYMT6ftViR/++F9HfTzDKI0JNY9x1oO0xMf7
+MZDE4Q7mj89V6Vci6edswBkTms2h7ztCZTO++VqQt/pIV76pQKkVqqbLZFMOgtj
8DjFMy3KNF3tTyKVUgFi7tN7qieV7qgr1FCBnvHH2NfwtL3Y2Vd9KVMWKF6WsIuz
9ffW/PZcbTerEMv2K9mc++/42ql0E7+xWqZciuU1L1sm6lY4hDUEVGcaf959Jsyv
ewb7nsA6zf3Vp+8lUPSsoxOhpHnYQ9Kxh1REC4eE5NZ4IdhGjQRaKzdluKI2klbU
IJSl+rsShMhSTDvw8vkmp4EkEmBslsKGopVZf3Rb+2NTjVagmT+6QQSPuo+ocZVr
TJZV8nlIMJNUOjuBFJc98186QHDYAEYAHKmU7Ejn1dvDhRLZLILeXGTYq/j7Qw2/
h0dg1oIHge+GHTxTPovqXckEXyvW/eXUvjrZ1AkpeWNfMMlxBS0aqeQD2IahaYOE
FnKQyZr4HCbZ7yelU0QKtrcdB+nQ8iy4YUMJcSVxNL0UD/yOEOMu+x3CaUqiNgAv
W9VAwAJ/SP3YCYDx9xsBe/NXa1VJEFUudWiWWNAeTSw2Bki9QXHji445QEGCiSFn
kseQ+k/AAgFQqzE0zGoGqYxO20L4jtAC1DPBUje1ADVoUepDHmZq/rzahOlDgRum
Bgmf2cPaKNWBULv9LprENsPZ94gr9zZWJEqhvjg16jOiCLNY+NQsLrwtwl8BfhAb
Bs/1PaBNAQUGi/LvGAX8OqCgT5XocBC6sl5sPY0zP02yYgVsM5EEDHZLAQ5hFCW6
+PvaOUbqHD+W7j/6r3b59pPc4/B5Ff1vp4x6U6yywiu8mDYbZgRiHwuOeRRCvyie
l18jZ0ijslGCSA2IDOnydbFxWyBIk12W0TiZTZSCV+lr3OSV3MFM4NKFuo5VfJyS
oKdQiLIMHlsGxhk6lF1ZFJgCloWPpcFQOqi2JNV3czICa+GeAsUNvh7zmF6Ahb1U
TnDeMPQkaxVsix3JTMKjQYKa6kLrxOp3nKIH6VxB0ox+qryqsqeB57Q1+oE1Z9To
qdVbbACkcdPhCevIi/DXwqsnfz8hCcuyV2U00gOWsMhH/awdgolzqubcYX8vdvy6
Vj8/6U4OWeBp4vt/30ndRmbPvFKJJPXbKdAavhdOqDeIQmiK5BBt4T9H67Dww1Zs
GA4d4aaaBdi5WFpvkD+Tp4TYP9QgxGbuuWgfUxFhZzPIKGjMiG7FH+JjL+JI3Hdm
o7yvjamRll4J7bLDET96x0LBRX5sz0wbMKyIV7lzjLMp6FLSf6S/3QGwcNNrVT1O
A3RvY2QtxThQDDLU0wgyYQmMYi702eoHmqOzC/MvXs+l4r+cYVM2fwEPy/M3kOWh
Hj9lMiJ95bSyiGHtl4H62pbHmuglsVjKtZ6u4JdMHGt6JGNEECjl9jWY7xa3Mwvd
pIE5r9gy+xZRrtXhL1XX0bUTEoMKLaQnfTMAa0r+1QuE69l7kzkQ+lBbxKm2YM/s
irvTK5p9NxmdxCZuskR8X7F4e9N72wCj/myf9QN//EKGv+UM5ciOYcMcHfXHJAEl
1UpxdlBSIE3nqg7MbAhhtSjwKyfhvObKN5xwROtAiADjlh58DiE5/xPSKjO6Rqv+
RWxvadQkT/nzv9nt/9OC2/dgp9/N1/hpLq2Nfk5xgTlmEbsuFSiQoQ2qv6LK/JHr
BoO5jrR2G6ehORB6yQ1uRP/JD+xwbVq4UbZ/wGE3ic+kEB0ESfBD4H7PBX5zGfNr
5othzZ9lovsSfayvnaC8WcERZ0TNZrUIHKmaheSbfTj5bUa+tbvV1LEcBgzLipIQ
6dMMPdjgYBfP9DZIMie5O3/S/xf6VaTsZaFREU9G7l08gqUD47s1OYbs20kGnUgi
vI6AOBEutEMjN7A+S8DZJG+s0b+Y2zRT+b43eG9a8OZ4cfdqqxLazhuSPNX7esVG
EEVX2pIcOeQcJNmumTqjsEGpBtxSdwIWokfr+ZVVlxMB+NbcNKvvNDjSzQ2gzwSX
snWbjLZ6Q8+knmRBr5/elmLlQ7IOdGAJTpSSn4iwcjzAqezldH6GpkAJuw2Xj1f0
imRKalAlDmXXDQm/DAA+xs6VUer9udpixYQKIU3vXZQJ9pI3Q0pYTZ/NAVFEgz92
XwYJH1GoGDg8+3w4psYOw4npMv3cwBZ6kBllEllZNxplFoRLehnI6LY8koRyZTcG
CEMMAP3mP9LHabaHMaal27b6CHMMqqpc12Ik0YpHewdXdEK3HaoyVZ0e00nFU+0Z
3s8uz0p4Fwk8MAbO9ucdFeKzWICAfZW6nVd3vena6RO2qXnbxjO9qRJ5+RjRpk2L
XrGFpbXd2ktQJpJLDRllALazKNcFhTkXiIBRihM4cNGrFFNWE7D5sM5+NFWXOqw1
+d8N6pka2C4MLBxtGMzi/YWtmBbtKeQ7fGmnwN18q0FgpY4sKNtU1fFHhe360HgT
X+gaYTzHkk6g3ymyIcYV44a0o9+wgbRZfJI98CRqTq8o/vj5UPInYV7Ytuj1IBkY
8qClrMplGaGWtIEKt1kFNE7V4kVunrOPcxOlZOqUCNWmhVi1qZ3Tj+owXlZnXgRo
rtKmjoicUQkbtczYUSu3+Zs2woSStSm17GAsGhJu/ld3mxayzgvDx9ZultRUdbze
LWIu13Lz37bov0sF30xjcEd/Co8QD8DGmhs2MK9YGEboaZIC3PEPD9sHmK68SggS
sYxk5jBgbgb7hUQF3PD3ruroigUA4V9kTWf/oVCUZXKHgaDNh8yo4OOoqF1JtEOj
8QpixjY9DbJ8IM53+Ufw5Sb4TQXY3TNX0HUdlbJVB2q6MEBDbYFBk3aL/FtyjbP0
rWYCXIj3nsHi+ElUa3yWN6oDLKZHFQFBFMQAbg2cOu/OSyQGTi6WLQ192fZ3VqMQ
dF9bUk6J9CdZz09v61MYmCltmHNLgs5TNnoP07A/UuPv5jKT4iPcdlMEzbtPfYiy
XXRxbfqxCfTgnpPGH8DXGOc/vOyZxHh+3Et2QyFDBe+VUWrEftB7yKPeUvuT3imh
7iSMy3jE6SC9ltNqQJ12mxHhx2N2i4ATa1Q0Q0yHxfxPKReSfkyiTmkHjuwFA9vI
VmN+irldcBP8eNxKbTMsHlBAIKLvBXCXDzMnBYo1oZWP9pe2DLdpPWPsY+uhueDa
EIHvSynsXkZhIGxjCPG/5nvpviGdmumrrzTlcEMCtgKsaWqwzFjZ1EoacHbzQsw6
p6ZrKyLchAwsRYP810+nCeZ25bivF+7Dowv4n2GoUl21Ac/rNBW+bSLXsD8usM45
WWCPF/9/EjikMZA+gq5Ud/j19yr22MlTlkYklZgRfOPxfMwUU2nm7yAQSCSx5US9
MQBStEr+nRyrmM2qUdQLKcBDvy2Pqq9goJPIgWGm/rI7ggagUK/D4g87Rno+Y3jK
Oul8fjjJP1IqyPa1F5tqVGHVyssNXVi2eKNPR4/wt65dmFXuRpvLLKicU3RbP6y7
YjNGaRCbKfOi+Rgc9vGbxbRg0X9cI+IS/XaYuo7uY03DuCla+Vv+XP2U8E0a0esT
tY3Xtx4sJkL2/uHg5E81ooHebJAN2UKMMB/vWUv27hBqnsA835LVJ+Bj/gJWa6Xp
5zy3VsGj/Y1Tg5kWg6+wMGXg5mYnQRrDRTSrHxnhJ+3WaauCiwfs32yov9eM15I7
KWHpA0pGDcwxnmjmZ5wWby4tuel2wT2v1B2WYSGu9BxRdCnnFX1DXm3NEOsKgzD0
2A1FAMTCjHcCqxGtPBMSsxoNht2BBhHRu8Uhr3/KW8TTvD0AxWcpWxjxLq1eLlU4
FK/kRhsF+87rRIwoXzMe8ZehILqHZgw8uw3xcx9+0ExgXd9TtIToh0uNGY86fVCY
HCJ9GX07e5R+0tHunbQmJe+etOgICi3hsvPqwpt3v/42vvtYNx2MKiSLB6pPJPgp
GyB1wwhI5jD7Z+sWkZEqCRf9Z1T0TrXPAbxV5sg/uKJ4AbgF4Tzi0RWIFHjMiTa4
2yK97FdkC0hpe5Oi8pHlVmZ1rU5RebNYn7YlGIfacyZ566YGi3dpSdaT+B0KPB8X
zB1nqZqI/fLbaf7w935ZNWu+dWE8rKPTxIsUB6c5+NRhAx7Ghw7lAG0JlNyVcyxK
5qIrPSq+73tXod6dcX6emI93Fm1T6+G0Sv0VLzotnFXtvgZYmPan/EBYw+km+9uK
a5nC2k7ev5xLDE6LCFkHdkHCT/TnWT84budZlVxDtaE7cuANoA3oLl2BOEdBxLVR
KPvviASwWc79tfRx/pCk+DQFOey9/Oig0UrmJg+1iUy5KH8k0swSXkq6lVcplWKc
w+vUv5eEKIaxIBXp3mTtVIdQPiR1Y1VjK6KWNbFu86JpI3UXjC+22yJXgOL850KI
g1L54cyujGg2sqhGyrOkPx8imBQ9gMcdpuY00bbwJEmnPiDEcopzArY2vDDDbmE7
NA90kIzAeVyVhOg8MN/j36yEiFE0PVQMIZaIB2pqka3sQPLeg6EOORVl9H9PiYYx
+6B4VfYhlpsZac0MRQB1ALZtRN2hP0X4LxjCEUfl3kMRUHQtiL43DtoKHTpgdE1w
UGrC53EkQ0hXIqYs1B+TDl9pOG2dSeHSGDyfxP60hYrcx+bNbb8LxbUuw8JCXmE+
Amc9kvwQ4NE/CHVr0zG8MtP8QfJuZvNNeAqHtOczhQ+MXyxFZTXZcBNvTbN2wMLs
sPboV7xC+M94m5TnPdIy1IpIv9GlFfc5Q7NIhdpOBi3MiDwvT76R5mMUmBmHhN0n
gIAibA4ruYxRYcS52KuqVqoGITg+RTnR8lYZn0z+in9YACm1t250Id8jNwjjfd9A
Wq60V5OPzqdXEMwpacUbuffWYj0fWrAV3dUR3NwXZ4fQ8bzOj8a/ANdomUo6JzIS
PR0yVulsh3wpvDnGJmGu8tuD0JxPMHLr0MEHZu3AiTip+8493ojXmhPEf8jMsl6A
Jyy8HKTZtuLkcmJR3/Ii4yztgQbdCf9djdpFMLEirgslrPMtDDiWYpNCXaiFGk0E
qvDZXKeAqz2wC2AQ8dDUE3GYCX+ASp31EW8hNCtyC4jHS+3Z8BRvj3IOY3tZecHr
OaEo8TePjWiVzT6YIQQK2aEl4DEZjcTGwQ2THuXnO2BScNjDU4CnqXs+Y7CLEYqj
+Lsc7R0nU8H2d+EmIg6MzbkdlE22Ldzjmsp2jncQ5rlZx6S8ZLs0vH/xDHp3wlyF
0z52UqwJt2L9TjomuphGqrRseVO/ByFSLXrI4KP463NMrrot/Xg8seDEm6m09F7N
3o4bmGyjVSewE9j0cckGeQ8EC83dE3v1wfuiKTio6XDMBNQjCiHxw385eizQFnu0
kux+WHBiTv2WQ2YZl6ydzDHxoUON1iLyx3FLPlkavVrmEHo8vXz65X5t7EYuBbUD
2DZ/nydR4YHOnFmA43TyQvbTdqpy0c/KNLChZnqQxGAFHZnKYFy/MdoFiQ+MoE9K
C5bMk1qpuCV3pE96TzyHIm9yvMB8heu1su3qC6hOHIPALsBaHg1hvhTRQOt5rBna
YZqwG3t3C35MPvWWB6bayRnWWr8upVblSA4qdf5xrnU08QJJqD1zyCry+iooZLAK
5InUYO3r2PBxvaAgfQk2AwVJDEgoZY4xAyQw4mFo3C6Ydlwz8dVNZwn0mzqADXf4
Ml8n20XmQdbNPoq7F/Ke1pthpdHoUvr1KZADNvLPlek7V8lJmQnx/hX8Q2lVqg2q
IcStB/kD1QJu1jUJB+mqBnleF8nxdR+Xd5CcXWcDfHhhowR/e6OQ9umKo/unWcsB
+wQd+Z8UTl72uRxAgpX9YqmLyxJ8/feAekLwr1+zIt7EUm1YQ2JOAH1B+X4qDoRv
YacZRntjkfeQdCr9UfY3WU0kAVk4koKR0E105tdv+gKUW/W20OKnFlQ1sP6tVHeN
88bh4p2s1EsDN98LhC1KY+Bbvd4B2YnVafeCHHy3m5seoV7hwDqR7s4naiiaRsyY
yJTjLgy2UfXjaM9xRsY8j/3DOdKvjBs+tIGIXoMCEJr2K6YX5xgrtXUN8evJcr1k
iB7hTJj75FLXRFO+jrBW4IHUgMLhhCZwJ0XMOnwautV+vmFERIumSwev0Swys0mn
kO1ZwzTairL8/40ayGm8Vyz9MV6yPzOLzDgY5pM/ErWGdppHlBUBqXQpvr9738SY
yuejvh5k8lP42WWpGZ2uw6GBIJZbJZXiqLLMhj2n03hk0aNxbOO3dzgqqy7sFXve
ftLvps1GRy+odN+InJfq+63M+Lvt/yT87uZf+FA3Gh62wr+SLHzKBfgZWyzSN4pK
IzRzb4a4tpQUbuUoLcnERTCnfH5MGWwKXTQHvBer2nvi4/RXUBozT/nm48aWo66S
RTEPyZdNzdf66JDjEdSH2zSRrzUTDqx7OR/7vTydP4b7nx4y1Oh1mKgtOuQSRHyN
Xkcg0pbmnfwyTAICDe7U+tTmdxM38MHlF6HRVook245elMFGR0Faw7gGH2bLLgAW
+6ZAVeBmMShN2SyVwqv3Tt4wgBVa6lAN5Px08k38pR678Zu5n06mXT0NH7pDzyTc
XqV5CcdAKTr87il1oljp5nz8+j8TXzfWEjeRRiVDcXzCEGAjXAci9k7NOOmW/C0D
u1mkgeOFyYeo07WieP7O5r9qQtIbiCn668FzuDDLBe0PpOfO0jaQIE0OG1NfKTIA
pEeLcvEOwvZJ+1wFLUJd3WMoav7d/ySEtbO2pRn3/wCgv+cdF3OnIjVUS8eeHtab
jvVu45Et4gONmwHURVglN/WcQrluuw4RumJrN66aBW475N/IO1QRvUz3AkbS17R5
zJTfC085nUFMuhumL9B5CzyCBa1CalvbcZw5m0zteJWU5+4acB2q+BLsbxfRSAcr
+SSMbI9JvLqbKbC9CuUVNmI9c9s+ZXTQF2dHHOgNcHz20rEgEJGjstjpHSRHsEHM
9CIRkxl0Rps1acSsG21w5w9ZFOsVqw7chNfRMKEFBP6ndMzt4kn1pUq9tpI9abAI
aeBP0tg859xKhzogkmW1hGTay8CBWy9E8ZJYYf9yOkoEjYNhOC07ULSPGitlpajM
561TZpFa/vTs8uo+MYVpVUZIFu6rlmpD0D1ws4uXN3vvLt5jBRPNeV0w4qxoFF39
IuLyskcrTpX5Pf7ql1LXGxHxkgsjDO38zCxVW3Oy1J1+yKvOt5mGPVzEQUSY10O1
/07LTDJq0OK/KmMxwscIDDkCEi8oBFwTnVQA2Ax86q0/dM0aEElxZI/p6ZgHra80
Dhe7tCbPnO+1MPN0s3jaERjpqZKKxa3oyr8WbGNaydHiiPScDlRUlSdLte/H68Zp
dv8ztUY7CU9+9TplzqyuQ4FR4pRk6PRUGh+i4Q1vFQQmS7pfKhoA9uaLTYNhPqIb
VzggO8DUsiHRbZjJF5hsRVoUP3LODFmBLbUxnABRdML0j/jq7aLflxIdCyi7mwBT
7ZUz4Fwy3PNsxVU6nqziw2LKEnAjKRxtt1jeoYr1ltmTmyuEKUKrB9A3STVkneno
z5PAOJEpUCkyuBtNlqYpPKsk2Ud1f2CWeyqUdWfjP/gWTXMhgUqLQGIlBuf4e2ZX
A0CYDtONT6apME7xIDcGvzD67Ge4RKlk7W1KwwqaPmDS9JeKzYmwqOFHeml+V4nY
DHpd9YNdGpQyT7Qcx853omU6hhAe/KllEY0fFz+vENT+usCgdo80zfBSh/Fn/633
cynJX7eFFYBsGsgrxeEIjvk8KQ57V93LY8X50iG/z9gKu7IEN/biUFygdm8vcVRR
Z3pd/RDaQXTTHhu3i6BJzeODOiXy0c/9sxbYSebsrLF1m5y7ORjcprxsxYaoPIxc
VzlFQaqo55pWGnzJeU9cTLu59JHRctY48vgzzKBk3quWEP4kQehIzZfSa5DpCjl3
20wTRIy3QmUqgT1bSVGn9U0YrIqDpbtCTAP82mKfqNK3J8gzx76yUbAUOjcj90r/
urbYbubggcwuqOEawOYNMz2eMMGQdCSWnYf5ckYd35ZzhYHWWSpnHXhfbPNVg+5X
kTlBgYTHCJVD9R2f0BVtkH+j4WF5fItYqp/Xj8HSHvz1QBWFdXb5ms76bKxhs486
xxKhd0VrDUDK5JiYCT4cqo9X41d5891uqR7/TnBIB+2/yvxcmQGA5KMjpfEfudRs
554Ya1ThriLdZrhMi2WgbFw7KZgTfeB/Yv6lZBOy909KcWtuGeMNzv0Yoo09MXL+
MElMuBuHrQfZd2dbHg1NGua5IFlR01rgevYKyAf7R8OvqMNKlCQDQNcysdHbyPNC
jtcG/GFgyJR9ZVOrFwiH7XT8JOfMxATcynrPmoRqYICd1i6bwoZn2o0rzqhGM3Pg
nuqR4djxc2oeH+fXH/H4jf5dtmPZv9Dg8w9iUR9+/sToedgtHPRT5kGmRgXZdrEn
ggYSOerhqB0/GOhwaAtDz6w4YTLwKx54m3aqtrugBh/jSxbR/K8eo1+9DfOP9Pes
VEopmqyi2WiX6Qx1R3NDPGuJTL9JJGL3lvCROIiXFo0EQ9xc0aHZPbVmw9Ry3l7x
kAm0kp1LD3erIcB5/z8pRMukuDeNG4ikVHfWsHXvmAMtSNpGfLSMPXeFclUnuCGt
sjzM4a0ajWlmtnr/CLD7ieA/bNTeIRqUDPi0EKxtd4KhRpLjNuZmL/zGku1Qvlon
1IQcwoJwwvalVnVqBRmPCoUtx9bwNHviZrWeO+LXa53Dyu9r47doJ1TpRGKsQr2p
gwS5tVLt8ZLMddxylG6w2oIXemVpAjaX7nbIG1CHj2Bg26F2mCr8zabn8XNVfMm/
FZ92NXu5BZhroTW6s4ikLIYNd9zI5emglMSU2qyIGRTfoxRUN5RA3Hx8XPJ4YsAh
4PrEpsCfNOT2GBGaulBr873k2B7mz5nvRmX/pfu6EcQjzG+8CnM0Q8s4xY8rrrOJ
LmyIfSvhfpfpZsfmxNUImDqeueNgjVGemEWlSjyXc9+dY9cb3XADqCTopQHI5v0N
dbZe8F9aT8uVsMZ39/N7nmuaQEOGlYv0I7uBh/wv0xc/UXw1n2ybxfyF2I+rA9Gs
UIVnnrUhKA06f5ckavIkbooeJ0YCgc2RlKiOhCzhrGAQSIlIN8wQMPrRiMW2lQqK
1zWnRACC8wPCraNazBx0gU2MEmTArD3k3ZYvmVeNAw2kmS0EHvmnWT0CfhvnX7UR
Cnr8//p90eZhiFOKVI8cxvC6GWdZnTTBKcQHZJ/Ad1/34jzrcXearyNj6M3QkzcX
+FfRGhDZLGseDVIStRQfLxMiiRo0d6GX0TptVzZRJRPLZGom3dLyVF8j6OOyuwDh
i0cQAdMbTmPUXd7S//Jqs2EVGDr9UJRv0NqAkJKDQZjLZ5N6BjgDS77Udpc6RKFi
Z3E1+TrAEOKnq30hFR8LdsrY4t7rpcWlrmm4MNZwGub2HFoRmc7erzcLGgi68wQf
HjiquNLjDB736tyhdSNY/ef1AIjJrxKFdaHZg9W61Ykjmv1OtarE0ZeNnsrsxY8M
hCK/kmdF98kbk18XLUOYeTl4zMzcMTNKNIFoJcAMGHw1G8I+8IrOwPw3R01+nOMi
BMI5e20/3RoQQ9f0HBHAmH8iOlbAu5WcXzyWNx0QraFI50IGf7rt6Erb5Jntks5N
hihoLDDYk/ctJVzr+YZa7qu4Q2xfGOINJVnncXPIUMiB4iTfUf0/PPIqaT/swGHb
azV8GZN6mnqAInUWvlnkTtQD8Bf4qWDl4/65KHxm5djC7jNXqULmO9rQ8e2BsTmt
PmJ3TUda9evM9Clcio80gawDellH1CkqBeanqIGAL6mJwbOg58RLQxEy7Yvdx5hA
EjU2A3/h2nfaj9uae2uf+WvohjkKkssLDYAkc0vJN+SoAX7FYjZABNL3N4fIEyXv
e+Ol8ViQLNL8QuDJ4VngQ3YPBqLckRN1LLeGnvIqua3AJGkMX1TMfLmGcNicchJb
pB6gMKjppKiBbzSMxmjUwwO/+gE6HRpCRRFHKlIiPksRT1ODXiBaphKVj7SscKVs
N6/zt4JBrJBUPJ3LM1Sn65P0TAOw0X+Ler57fxSlZT7aYw/xXspjdhRQuPZz8qNT
ygg/6WjfIVvcVciDNH/pcne70LlunRp33soVdoLWw0kQ8Rhr3E9wuT3kzJrdgIUr
h6Ruh7JrRhcLo1ps/qjXjxoQ3lpXHZTroPcGCArcBRQADwzrizrD/BTzSoQ9mGwi
IUi+INz5NX48rp5vIgAifHGwknYeyId14dV/T865ZeTmp/HCD+KKQfCvxGcCJSaO
24JKppgo75GVuiNzlshmNYAFRDLUxJFb5zlgnaFczsaEMyV4gK3anl+cAJtLRaZa
XsX1ulC3g9+EEIa8pAIBpUNZKDVvYZitdxRcLnbibXR7KP9oK2vSRESL3hJCZPEr
FXOP9D/Wmuhl4YnwCJrgmtmGch6T+jFyC2cXNA3T9y1l9Ceg+Y7Fj+SznbhH5mu8
T0KEJsEFksuq7LdQz+4s/HlqkWDrn4JZg2e5x0mKfAPvNaKgwCkGuYE+ickAWKeZ
7qRvxb9WZjPfvOqq9a1iFao9aggI7Lna0UuXmy0Z0pRAb0QLx4Dp0qdl8azQ8kJw
nEcrbAbZknep5xrqnPu0CUx/SVwbv6JJ/HiWzzLSdI1E0ifMN1qJXFeYB9iyrTMo
jYzugySQ4HhhYmE2heYSb6PNTb2G+1cqiA3T+3nlcSsaobW25pcTlkxZuYJY1/Ww
fm1jwxdSizHhJzCQL1dL8E3Jm2r/erYG0UI39BDpeWmq8zLwbeuZofxzkL+Zu5no
eBLLhhq4N5Y5gKjWDi+jm1xLxm4jBdXmueellVaHcJJRZFwJvke6Y8m3u1vnRxkY
7sWfff2C4YwvwDvdnK3p/YRTlVEu9gzGVMrCOS2cida2NH/6m1We/03MusdvPmYT
BfeOGU6GP+AKhhkumSz7aQrQGPGG9ArtfpMGGWcOMe26yimMJjMuiK5XwIbrYvH5
/Z1RHlGoJAhuwJEADbocTWbK+enRZFx71O7bC0CxNf2oJn6vD9o7Ds4xj2DCUTpS
krnXhrgGxMjvRdiR2QK0jQ2OugHeQ2SQZHTciujsqsejqZiSv2nGrbT8A/VL7Wii
5gPo1cf4h/HBR5BNlk90WG6kbvm8UZDTWyjYLP3fyI1SArEFi+W0CWohQbdLEXQd
B8GVQcIJjdeKI6B6nK2WU69uloESJ5a/mbFVwQv15aOYu2xCKgik+IatT7KK1lVm
bJSp1YrIQWBI32KEhFF38Ted10929q91iei9fpqCvA4aVAkT8+WWY5ukkafM4AgJ
2eSJC0/SayW9i1fgHDQbbaBadA2QwtMlRiBCgTLFtE8Un91LipbTtUe9TH5CViq3
xPHsO+XlU4h4ob7aSjmLQy9Qnl7CzsRCK5/MVmcSwjxWYXl+xk51H9Dy8ly9UWMR
z04Cj9psGCvgyT/IwH5PsNHYviA+6pgpIyr1FnE7JhKRmulD0cUvQa1DnZEZXHVg
AcA8D1KTUJ7lk8d2Zf92R6Umg/BB7fSTF/I5ewKFNquYw7FMJuYxT6JV8u+ZhphC
MnSr81U5NYnEc0xj8U9el8SE4I3HboAtKjRaRr0z9fweVFMaxtQ7qtmLEMp9q72J
zB5tuIQ5Fyif54ihMvd0vSB4iCu+TnTeKon6cJLE7LgnAq5rRTHOnqgKwDTqiW2u
tE+q1V9eUGuvl5AdLRL8VIoA+VqfjKnWz4NTl1eA8FbJqtV/T9Y8V1Id7xfnSeXb
4qGDplSBjujG1ijLqtd1qFWWFgzct1G5t2JLzKdZyIZy+o1/46iolIP+LCYQwJ+8
fujR8FsP9a+ovroFfJJA8wXTf4VvxPia5SV5h68cK7VX3/SkWGWGhOuKMtnbIWBa
fI77ncuHSE6MK/s1xqDyz6JXWWvBPWxiSS7DGww9Q6qGiYR38WazxfCO8CT+050X
5lYmcBmIpebFw1q/OoSuhsL5n3IEMxiG8cb3g5WE7Y+FRfveT9oTh7MMZYUM2ori
k5tdTj2hyvuAVsjicymBNxQrgbnZETp/VxemH54Wr78rwvzY+y4/OSjh4FCNvWur
134lbaB6Niml19maxqSgJT3B3u6y1GiEFm9lXEulLnXxuDwEGKq9Gu3GVBep4mHn
GG9XC2XozeQ6UeZ6AxdftEG3gCKTo7mRVCBddnn7LdS9M52G4oXYvFauxfWMJbOo
wE/dwcgttZPHj9IQnXjn1ouDrTiP1YvHIwCR/M0jBxfjtLSedCMnx2hYmJKtV3ez
qHGapqBWmZky+KbAv8l9916pAaEZ3rpTDG+aihPJaNmlYD+z7bKrZ3ftgYHZRCIJ
WsXlaW1wtw8/TQax3f5ljdbWfBBodaQDiTdiu7Lie8KZ0yF3Uq0ggGGSLbKnFO0U
aiuhSfyBy4K/fmi9bYeCF4G4hmKP3OEGNJLNS0sB2tofDSJHlpWrjwUJEXHuBvAj
NmpnZjhsSL99uvkFRcN8HPVQxIqUvUCaoICJe2QuNis30EzfBhpNGe5hDgJA0ZnU
PkaE4SEm+EmPSky+bttikYJc/0IlX96u5quB7pBxPNMlwrXAfXJ4/LXQawpmLXRB
//RxScBRtF/QNkuJcO6gmz17D8ePG7MNjPou80p+0ovTXnJdS/dRtb9U5ZARwomo
V4Dj4sq6ogrkKbOq8IxpZgP5J42QMazM3p5iK1A3+YIpLMyzFn009s/AZHLyR6ep
62N9LU6omCvaOj/sBtQXCvBJrT+xE2CaQouGinxJcZB5xFScTF/VhZw62lH6re8c
g3LvvAh9WnGfiXRqV0/C0wgFFFccDFnUxYqB9LX9nRzvlT0OMtut2QVcxnRn0Gqd
wOzKwS4DzajTR9fppQCUS7W6F7rwazV4qDDSQsAsCNZ8FY9OHplYZgEaDsm9ASp6
u7mQ4LudpO76OrAXo/NzAHxmgWfGl6SHK0yuUaDg9qIMSha/M/VppFYZzkBeHVpn
jhxFPcXj4EAqgD+pk9TrVhVZwXG/zTcbx7U9Qq/xMghk42K2BS64C3NPsDcoF5qM
T9jxuFFZkmdT6VAouAKjgZU+Qm+XmMKkVkm7dr7cGSPWAd5Zz/Dwav9MrjLB9yy2
oaTgHLejxjEHtXfneiGxY/2Zqnl9px4yEb/VDz3cpgvr9Ii0aSWWXi1IzsdicJiH
tUHle8jQHd1bNGN/bNceNah/MCezL+CApxFp8+rCkoZ/KdUOj0gp85Tg8YEJ3i72
HeFfRb4EGaeKd8RN0E0bnag+GFn4wGVKAi4ntcE4u0wpjhFD7HVwRAbBvLhnUOGC
PwREibZ7mDsozg7kBxXoIslcBs8sZKvS8Zap5SBLriYZ6pPRddQHfy25rSdKGdXx
YrtREbiC58i3IEBV9UeD7uliAyJk7HrCHxGuTKlDty9SM88PKwWc8+auGX1lvdFV
vvxN4N0irFJ8CrKokUXrOJn5QCo7su6Jhphla3OMRFgwKXhz3FUvbyDDRqMIb4/z
yMCIKHe5Nh2Ntb5B8vkh+eAROtjjYlXJCAORqGqKTcFyJxZ8cipsq/00O5Cm+qVZ
24DvdIil9vErWTJFp89h2rKYl8rO6L8ExAlYBkkbMkymuYE2GQ3eJPfigjJwhgED
qGRHhz40+kg45DEObM8aO4VxilL4CO0EBl3Z4+tI2j8wJ6OSDtocjdwyeJBhD7N1
rRxAQ3qoVDPbvVAu0XRCnTlOLF1WXXiM883oabx87+f7Rqr66OgIDYNfNSbn1adV
UTB6ULBMGBgZ68YMwwDkfcC8YeIKo3XBcBov7JjMPkBHiVJnk9eKVsczVsCvQWtN
/QHKI0cZijNg5R6NsTGhlszqk30/rvSfW3uUPt6GZh9QIKPfqf4S8RC3MfyE1669
Wi84Hr227r32djzpWbDyVDIoZS5LQsBgM5RtuG04zjsSEls5C4WlEtWauDDbJzZX
CuhVFXUrNiphGNE9VHd2+fi/t9KPm1SlEsmj/fnzxeir3vfYAgo1OoTGqYOxn9RA
KxaSWgdPaPFFYYw/pGsZsFXymLb+mzSQqiEyY+NDKYWI0VYL6/2KOJmvZaysg7vm
Qwu+mJT5fG0ujoQU3+n3L7T40s2oKqEJfar0xsDir3BTmtNdMkiy2wZGseiALvvM
WjjFkIotqdDytsWa/0wy7GXfY+9szKue7QdOFs34JwRDMC4jwc2Yq2JPF6i+BNov
uSYNfxGZXdIzWY4k2Gib+hRoeYea8/P7VfArQJK23pbBi/oUZ16nl9aiMR5PCBqs
Xqpvfu/HvtPZcgM7QaFEtWo1y3Pm1wirpKFBEen6tu5PG4gsLfiNYK353FISl5Sa
sK6nEGfkWP3wnpMAzESPZJ4p291WbLmpMMA0ULy5gHltoexWFY/drehQwXJQEHoQ
ALiUUNCIA3GrMt+D5tDJ2vHOlV/emi7jW5+NtR7Nys7ky6YHdc7FIWnBZbgntECx
yMYu/RQ2yUTK5f8KwTiZALcUXjLeEDdfAN/Hy6LTjIA=
`protect end_protected