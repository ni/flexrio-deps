`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
j9eMmSPGcKCWAR9PvkqZ1R001FU8QKTyJzFqNLn+qur6INyYDE1AI8LWcxAzfnTc
IpZG7ua3uuk5/kQKKQx8ZIPLfmv6H3t3eWjki8YIAtY/d5E7Gq8Z5mNxMYRzGGTg
TCMm6oOrOTVYlCXHE0X9AW696Z7UGfWirVibl8hs19hrFdeZKGiGht4r09vHR+Gl
FQQmSObM5aSK5wu5KOrK5ZUKGHyBhjnIQO5NnittDjOwxV/57nHVg0pdG6JUqyvm
tEgmCY36RCMRGWN7sekPtNHjqpZkmYrVX1T9QF3h73+8ZekZYd2xY2hpHHGYYeWA
t3+Fmb/6NUmoP8+Pt2hI6g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="wX+NBVcG/A5ruHK3pkDqG8ZVPdOz9TJPJ5saXZYSeQ4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
j/hqWUoxjK88VtH4QmjIrexFOSwtsLKOZ/LCP4cmrqgzmR/e71apdtoL+o8nlfy6
eZxDZMmrZmJGoazz2oK6kz7xJU85UCwNc4cxAsVxNdCP19vZxph/nCYZQ9lUFkLH
uLBkOeFP15CD3jG5/dp945fHP13J9SzB/L9PWvDC/gY=
`protect rights_digest_method = "sha256"
`protect end_toolblock="sqDZkaglKf+bDjC7VKm3lOELrT2Jlynh4UhPg2J0Q70="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 35344 )
`protect data_block
f9kZDbPp4NLiAOFOgATj9W35i3s4a7wbt9jeHjHVcJxMoXY8rb8laqS5bNUhXGW/
MOc7UNc1VwolqhkS7G27SLamkGClZZtXSbRcN1N+5kZpEaBEj1343vVznnU2Dre/
9Q117ZaagFa1275muC7rLrChGUpWgeKPRf/z276lGCu5FD4SMuli6oKTM6AvsKrs
JdWfxKwFnD+wq3aneftmYQ+S1OUaHIYFGgsQYacY73t1QeUT/yqqgO0pqUE00eZ8
cAqGWhQljd+2XCtenMyP6uNw/EXlWX5fb5/TFlOdBkpfIr7NuXX3+3QrRMG7L9R3
vEz2TgysTNTX9By0LG+14iXbotzp3EWHXB+/E0vV3/ckkDkPqmt6nbybQ0J+Xbou
/PGg6e5WCbWubvTUytyQMjY1svEQ27DeTCRdQyTvJl2XpFZ1ddgjdbYGj+Q493OM
yadrQTjrBytdseiJzeqmbQWJ2Xdol+f9vplYCKJoU96hxV1S6fVwNEscSNE/KgWr
BBOjIPxp5/A3meKyuiE5PjCIlvtcEiW/NNBjr2gTc/kgBYKhlXwVTx5domf6ai5d
7JLbitGqzTU+GK4KsFY0sWXWLB6aZVmtPTVJ7OdEKcXfbGDRPYTTYTEoyf4Su8/G
tHWG9FcQiiOEdTBV6QYh0AhjsuhyZ54LnNXbMPHzl/qUxOmLSpVJIBVgwGa+S0GD
/BGpsPIaKwMiknjn/M1IEH6uaYzbiiK3foSGLkq9rmzW7hvN1UxcK81v/AnMKKRm
D6Uhi0iZRwSV622QmUQWN3PSAKr6lWBsKuhEpXTa0BXH2tQ/M89RWwFIeIcILHGz
JNkXGoNbGWUSuTdPhbCB9vJT34TbS4DnuZHhoOsHyJ1tPlmJ122J9usS/6+I6kKn
JQh97yqbgBW0Y5nY2m72ZeJD1B/DnKb9vyyhtkjttNh9C6l+SkirkjWX3eZiM10M
KLzDPoe9mGwE92bPCw1rZPVYjkdyP+HEqaQYh1orZbSExwtduhfgVhXbmr22kcaQ
nv+kwqZpjJoJG9H3bCLOiI1a1bPRC1faP7DH8RFOPV9+SBz1GHWSfkX93iFySONg
JA29dUcBVqDEY5gZ5ERItJAyR1DwzMkJnLb3oeu77/K2vaqeI6IfAn4Jthcy44En
19mofINCPXT+xduHi75IoUAoJK+rRY/hJtCh3NIeRVE/IR0us1fopc+Z66qPG071
1+lmgK9/tcX9i5zmAymJwTVUwU2ImFur4CcScfyXTiUJiX+0vMOZF09tIqIXVD0l
aW+ju+fi+rGxvXRA/PHmbdO6zsA30EKT4pHyLaUF9OZLcHyRli/ia2ze+wawMvf4
LSJ6pfb/lo+sUtVveHgBVr7m7pldHliIVnJsOnQPzRG2eR+VOf99jTBpqrznnIo2
F5sSFH7dCsN0i895XRUFk2lBIBy0h7LpJA37KxqnsBdq8iZC+IAamlz2m8hsr60l
L9NxNPkb7m/zhRtBBJydTp9QbqlozRtxHWrsZrEvbPfOWZZlfhFtd3ldQtcokUP1
a4YymtX6tjZ5tg/VETPG/46kkx5bH2gX9cTn+mniEjWcdUcoM/2srRmJTaFe/1f1
wnplBpQvN4sJ2B/jaAv2SaMqBUhtl5nyLeXh0D7DcZwozhvWun9kBo+vlGNkg5nS
LNwfhgiQ+m31aKYEYOMX2TrPLyasagK9rfpn/1P3fqKhhYfI4DpZ6Yw4s28Swl9l
aC+vqLuk/GuBcmyxKHEX3p+15x4NSb/teRHKIDU7iGWpbgvUCiL0qxF3UgN7b1Zz
gT6KJ2algnftZGAIYpYvXLB/HauRdEEDFQm1XQGVb5UqLAq9nVNy+1G1LpvE25uB
1Fk0Vp56VljS9ICeLCm9C8Wty6URnNziRHYeRiKvVjQ2/8aVOEjgMpUucFI0KMIO
WAc2h1yRxegBDt47ucAozIyAD7YhcXYfRpiZ1Lz5IqK4FgSN5DWPaPEh0iEVPSeJ
OZYj8Q5dNyWmF52nMu2rOF0ch0lbYMdoTNQ7Ykb9j2Av7tlPJ82sLdnC9zQeQz41
3Tn8VgyXwl5M7+XR86qaOYaVbcAb52lrsMpZJ0pIPrBbQ8Gj25OKkYSZhui9B7OZ
BwruaWNw9iyc2GKGsIOM5XPBGVZZSGwFeoYk9jiao7LIB96FpJUyFWWueRDZLYWF
gazS0bqR9SuwDeQwkuCXvqLs1QMCHCwhd0ZEXawx52khp7Z/eAi98PvzFTNgPnoZ
4UUWualcMxQBedW3Q1QVFDe8nCBK7JAVDO250pdD5w38d86o7AOHrWXpNm9c/S38
ByDaTNBDu9iZmmMPpD0BsehgFlp3CnAfcICWjlQzlU6rpbcltQ7s2nGxim4iewe4
G2uNUg28u2wYNZkY5hRYOCh5OkFLPzuWkbQ7vFWP8zr4ofEEf8sMXQSdilFFrptQ
44s2BBMlr8rjEqBZfDuz1pfDbkMv3CcnU8LANFgj+ZvNoMf4q+m4ZQSf55cz5yL5
MBNZSmexz9n6T0dwbSrBKwJwPNKeETtcQcI9Oeo77YSLCN08g3QkH0CH66f6XMFY
jYZs2hZFCLP1mFbbD9lIKXnsIuJx0AX4Jo7BXluMTkEMtW484mSQEmW+iJEdLgU0
sI6HUBADvN5gM3kcpFpK2AG2mXD4Ojf2XGuJJmm8KXEy94qMnxB6ke3I/Kre/fsy
w2ZPPR26eC7RDJyUPAnWHtXqGSw7igHmgi7pZYuZTT/kwldzqCDMr5v/OkrgpDzN
tp6j9AiB0wzwJWOolMexyb0mrXLCBYr0Ka9g/0r6axvbxEgXF6C3LiRaoXFtVFTm
lgkn06WtNCiUUNhnuDXjz+25KKn8dFO5FBv75KBS5tRyYtv5p+H2LWZhxOh0bMdM
N/eTM2HnVC2/baY4HVi3LQXio7zNWEAsVRZu/lLq2dk8XLfCwlDe2ExOP6Vuy8Hq
CajRaIR7hQaKL6VLKy+2kV4VUX3mZgoj3hjAoGZ8/hBaf6GHLh7pMJLCTDolnn+E
cRYtncQqecmTENO/8VU0c81iMPNWVsCqIWdgC5rTELBbJa9HAvjdmhkzTxO60UWk
YDkDbsq2PO4713ENml+QgwmiT1wCGwr/7Fptrv3gDCTqChlXBdL2xyxYEAVXJ3Hn
rnqjZc3YZliZelogy1Cd8AT8PPqbQFaiB3g2iCXTsMiBOErW/v1/lehdwgd+lydo
7r+ZqZC2LiS+JtzHFc7a4ZK7NILOHiJmC58iSCRIkcADBR7YMBNOAo91MK3+NDZk
VZrIdBMSB3oSnzqxdsgb3m3jNBOpYIhf3pNk6zB+r77d11dhrCdxwhfqYA0syiZ6
3orzSfX9qhWY0BVU3t9yoG7UZcLHuyZeEDBJe+mcJu2lG5kdtZ/25C/baqOw6JY4
jUm/P4sCypUz6PPNppNz2fN3WK0s1DHr5sciD3NOtvO63YaRS/tzc89NG3olgHS1
9GmUR+WBklRjLYPeVnZaIm87vMgg7P+R6OTzQ48xsdGZ0bC7iUVJdCxotGOfE+eZ
FO4bWIbco6ujwDKb0mJMP3+e7bHr1fW2XpxgCDWYrv25+UbNjOt+JPEgsc+jDbW3
vEXuQoUtTOtIZCZG9P9luciUynaeg/SDJmPtwKQHskJvhleagQmFL7vDeaM/ipr1
4hmn6uW4aCRv9F1XrnxFnLAVVmINW1Si+rCfQ8mSoOb83/VPWLm80wJI93xS/vZh
LxGUOFMtNTdg8GpXAAZANj/4sI5qQoqz004gAGLOsFob/C26PqoyiUxi28dhbtK3
7ySn8otkISTK2gQ2LdbzzsKlFnPnVV5YepTI30SZ3Kp0DBOQ46/qOv0tTCv60lgY
o2YxZqPqghFJrLONYDh5N/eOgrhS5NAtD35IHlGfQvlD1WhvPR9NhkVHe9MR2gHS
vzoIV6DbCkOp2im4DGg8ogdBbJUDtxpq+JMfk7TDEHVJZzYoLs4YurGU1GPowhP5
Jb+D9AwUlW/gexe0nf1Asiawlq93WzgFjmHKMQ6RSntAnkvNgU9Ebe1bnetbhNkw
2KZwF9/T1Mxr08ci1b62LEkg8Vuu533WGgPacpyimySs+Lz/i6yAXrjeBo2lMfYH
I3ywtyrJC89dw3yKFlBkapuQV6mKFrpfjXFIEI8y4yntE3Ex3ZxmpN6moVcLe6bn
Je3CFQUPDB+5AsR7Yu7VEacKxDyy1Pghlq0TdzCxMyHsrSegX6BrsM8KQLbZUWCC
5SwwjnuvSU+okWEdbXvEHNqMM+ncNrFijg/cBZeF7iUi8BSsG+MYB0YtahjiZtmI
O2aEP+ks9FDwLSeIU0sXka6MXBKW4syFMPgd7S7XhWJk5ceJ89RRs+Vbtf8Lrrn0
00/1viaViEAnZvtnKSQEsPA8q6WnqDnmE98TWzIwTjYlxPtdp2WbcgBCitGXoNZe
gsAp9I3ml0o0/YR4zBvVne27XvRVTbrcoIinLjz293sLh10X9vybFfJVxsYrFQDW
QgL6h0JJJqgFmxw2anRF01lmBEOT8v4jG1oxcHXSBqmvgObLAUl34EZE85gA5FZ9
kAmwDWBFs5u8xoDH19HYF7oQQ2gwwQuS9tsMKRtlDEhLQhoL548YmrLdhPTCi8QM
O7HbBpC4dXTQlGICX++4+FfpkWOjKGokM7nRbCjQjqYfA6xxr7bOT5KDnIyTbVTq
ojvtKJqatIWNmALP3/ZMI47CCREFfpBnhh10E3iLSLUi3lJdNmSERoiePzcvUvWJ
8izhM1h4Zs7EgGctF5ClZuRzSYYglSQ4X6lSi67/PAMcjOqVOCuMj8r8mueCLucH
GNE6dTbTj4p4K6eD9zn2U8mdDNGKDUqqshh777vswLrL3YTWhp3GkEY3YF43i0hG
SJv/k9nwixZBpog9l/44eFw6rAVPRWaUftOIqTXYyeU0TCiwpTtXzjXVd7teo7D5
zMoB0xCtPn/xV6MJ2gBYoWlWluOmaCbD5in0lTrveo2dFi/M1okaPWXw/u7I1FXN
ylDyfc/6lVPb20mIK8WmZzW0SWx/NtILmVTyNxBjBRYtP2exARxtN+xJYwSryVZi
+dSK6kXzDpW8LNdBZIRTyo2w/HdbThMfPLuhWZqGugJAMEn4aTSjEjfkQmGRUJcK
Le0SJRfKkTA34NxacwYGJK/q9wnksePW/Hglu0yW5A0WdROc1f7Mo+SEvfpXBj5c
wYSRGNrL3ISLN97Wdjo07E2n9vrlUbmSRe6t9tG3ImEyZ1BrhvSdltzmC1PGvInd
Gd1IU/qYMeHhI0PkwyTLy0owHi6P/bMYr7fKihiEM/MMkSjsdQ5ETe1FCrJC3931
aPihYItxi9Gt1i+/U8WkmoaE6a7sbgzLKffJDCPqZ3zCgAezy2M9Hsfcm34+qqtl
+sX5oXILABy6AcpZNbJ9nfK8eKCnXyQ4jPRL2YZy/NkASMDOefl8frZiMGhK9uNj
Dh1sc1pNqrgVqCKKtiJ85bSFKAHAzksAmZNK/3DioAd6lBYJZudZ8u6yTsyhDda/
zpcx2M0A+TAkKW9f6b6AsyPE6umonxpBTtUHmod1XIIHDYKtxfr9Fg8mAWe8tY7V
CGz6nsAiHvgCSHB4rY0Djb+/YNmJYWjp2dHqcrDIGs+x28nojtIcytLPUpHsByeN
eNcfdRJHwSdtXSf3SSllHi3YDXroEIs0oMSFyk6iIbJchY1FgpX/EtF3dywkBXaR
6gGHgRZtvmn/WvMvSpxu0xDjvLczDLVwr9OgzV5HBq3+aqinFaENpXEUg+zEBj+z
QOukfl4E4+LfSH6etTor2y6XoKLn9WtDrkMpd2N+BP0hhmVdJPbwzmxSkpvvhtl5
tJ90TqTfpsPtvoxC9oPbrliPQGegFoVRzMvdOz2DNz1zBKFfAy9mSaKnF3ff9D2z
yoFLdwUkGIN/RHyJV9MJ2af1xzOR0aP6MnPRKP68l0hi2GBvJKTikBHy+G2yRNLT
XjKoxx1EGrUGj3GxAp5bEubT2s4C+Pm64Rz2xod5IlMXGwcnbynvGxDrhDTFYMdL
LShZFeCUdCkQvwVOC/50E7iVgml2C7PP4bt/uno4AewUbgXt2O+U+rwhDhVus60f
yeddTAAEAVW44G/429rlnhlpiPZZJQh4zlB1X5n7wyBVqtnzbDEqjynLTLJEyakV
H0D+LhqzxxYey+nJFDNQkw/do+BFAQHd2j34YI2Sx3QyexHFvqOPYZWQ6bXU+LKa
e02GWY8+5z+Z7zcck2lf9YrR8g8FbdMAjzz4hIXMYJBQfoTC5dhDXju0RBGoWx8P
GaDIkiZFLXvvdE7cmBa4gyBPZefjBbfW6o0gvvr0gNFXXCIDVBqODgIS/9MGFg72
pDgRcmNtTGHDNYtNmAbK2pmUa90Dim5J0qCJfKoG9sK0vAX/4GB2/nVf6pRMsaKY
EmAFLbuvirzbCIAtjB68lc9yYMPUdaAXPqkiCDv7amVYLZ7hY9Yf2cPJTamrk2YU
Gfo1BAkbCxvVzjO2NxU0Cgp5K4e5O7q4OrY8VTCu+ZiSkT5lZO1YpNg5Dk32RCOi
RiPN3KKti/lcQVq1bbXb7SCZv1uzmASXzB3vJUXA8pSw8hNd+L0+F5eT92DeljCo
zIHUexuG2n/2USQ9EXAlfGCr3mVRhpUh1cgUzlPBpSCZ3a0QdGeXdBeqgEl3J/vS
QoMjg9/oZx2QB27Ulba0PgyHHlaghLrEs65PoHtOrJvkjRRjjPH4gwVuXxMVD8KO
XiOHSZC0KgzAkgJZjzyZLfTezovpFJUe10LhmHNKBwL/vXGQwzI+H1HPr8lnk2xU
iS/yAqvQRfZFTiT7z3ZVFXerX0evyLtlMces1QMHbiVEoVsTdM9Z8w02XY1Ba5uB
oOtfBJjuZMrd1gkfsSe93CNgdY4Ml36DFyERy9MiwL9fnke9v1cmkCd3PNQgUVsl
9peS0JQ80zeGG4CIxp6QmSY4oP7eAtbK3aJNeIK3T6nFXJrI9HoD86TplyXE6dvR
HpSVYctvQCJ0FF9QtMxRHZDPEpcBp14KQRLenwcso1tjRHe+DxeYBt2Ib4Ww/6kY
69UhMpmg7fgFT7Zdl8/lnB4J8d+wuQWtmO7yDUmdp2b15FmSvXjWt3ZTRVWXkFXp
GCNbzIRsqJ9x32LHkqh+nMfWN/911YhwpeAWMGrJIpknhXGLk8uCztGZhY7U4tA8
nURWSJfRI1QP2diz4VESMuB94EBQnDQ7QGfoEwGE2AFiQ5VsP9lqEjt6jRrQc+f6
YIpXEzIjFjkuI5YTKHucH67Iq+Xl3JpPtHWXu3D5kMpdwGz1UNuLiBDQaOdVbSSC
wTCgCzbMg6f6i0KMTaTU+lqVO85mZqfWQSkUHkBXEAMboneXVI7N46KbXyv22aJt
S+11Rjsfa+xEzDFWdIRP5FiK1EMYqnxlUXHaXc/f1ii18eVMTydWqnq+Cy2o6G+4
CVxyX8NYFds7D9Hiz9xqlXQRGW2TeJR05EguBfom5KoQ1S7TIQxc+kwgfDWFJbZX
OclQCd/njVxxU2b5nDr9ZLwAzI8MTA07jUW0W86ZQDZlz2lrhKuNAv8hOfDoK402
UBujsoPhby6nNbUGxQdaZccZaiDoEA02be0sm7kwGh6VVbhVYO3OAUmrX387DP/R
x/yzN6WcImnGm7ZmVDNeIppA8ePth7LeUK3tUdc7j215lFStGQBI1PD6R/ckIZtx
r31/YDZYJFX1T7oFr9XMh+Pk34GG6sSVx8OytIqVKtbWzTCGJ9xqvfHmAkKqnLX4
rAoLe7u+o3Zl9Yy8YCQX54h9otVYf/Dksewlrt/tbBob9yb3vqi+Hzfgs6CtJaxR
JjAv4JctpptIpKjmHAiGk7LGTcT7mI5Y5LzBpKehxX8C1WFnZoZ4t8rwRRBUFMWE
MpDoFBPvzwMl6WjAdRy8AGINwhJWm5eoMcVZDPzFMMo03+GWZqLOVqA2VMT55PJZ
oJxt1z04GrInKE12HaHumv3ahG2smXStLcMwuEJtjU4sZkY+X4k4xT4KNLirYmKk
dYjYB3RQTAOhYx9NQFiQ3fR+lS0jsp/+oDdlf3qmeCjaP++YJbe237ihaE7faqTg
/ggwZFKcc2Cbm70LG2TrFaA4RUGwnvpd09RF8k/0Bg2jj8e5S22hq8Pv2PwBV760
GU63Yxogtvc5oj8z7Oki+xLZV/Sfpg4LkZ1wC+5bXgns9dXxx02nPWEgQwRMy8ip
B4PRqu9iQEXfmiBKuo90f9qANvUmRIK1yGM+1dMjMMuuPioPqZJLpirYm05u0j5/
/i8femOBUeTjV9rn4+LGXguvtsoR9mzFZOw/LRfIGKZZHSG6HLReVHraUL2goImP
L3fq+GmbQoBSCeIlflAzeXYb94Egm6MdqGRag4OmP0pBrGifdcHFCDFCvYfQCgeN
C5CcV0vzEZOnCZNfOPjokP+leaufUVIcOhnmxa2C0LW13oaL4EBFmyUS7AyZ7sAz
C+33n0N/Ffa6OewekeizljhmmMpNyOp3FEh4vNeu7E5LNEW9XRFObataw0zKjSiv
Ot+xJywCUP/aCyqqqFAzJD/rge5LwhOb4IGUW9ucgvBssLfZmSft4jbLHz3ZxtHx
LZZy+na8t7mQbD8Jcc6kI7yJ76o07/BATuujN5MPuU0yCwUt1dgmbdYI+kv+bzEW
c0KpNW3Bz5+7v2S2EKhIN0JwOhVz2tiSe3lVQ8mR+ahs0fvCG6CMQIxiuYg45+OB
2CJDF3h+1hWBQl8j1rqSxRCjS0FjNNZALOMvo7Brztw/xm4ypMpNQj13UZ68Rb+x
74o1CXngBZyYR/3PfwKy5AT8DQwzQHjTe8x7ELVBSno596Tcd7SBb6W8EX4W559+
SFC28ggpcyNyuMmFLAY608aU/Jf8pexGvr8wNKi5iAvS06kwA0q3FJNM1tdR1Wic
jS3/x73e9TPWUH7wKnJXWwar5JotxZjBTY1+xBvUPonJl9BQ/MfN3SyNgDXeOITS
2rKgiHQbwFuFRI3E0PVw57/ypHEiZRfONPxW+2waGhbjjen2hruh2W+CvY8AhmIb
RleDhby9oIYdcaZqT6MNT6Mz5eE//UC6VidOBGoUcKxRQjC0OdJsPIF6BQb/rn5z
NnVa3ERQCL5KwQuDfXqw9NChoBoB3/av9Y0RYh5T0TZCkJ3INvmMprAUqWvwQn0X
/YPjkjWPfIspjJ384FIxlGlxBwl2vCqDjJwzF/kw2C3T2DIL/eYXW0s/ODzphKhe
6Rthy7fD1h9tXV6lnjeqa2u3HUXlzmwGnz1o5GTyVGF2JbHdfkPGCvfTvcG2v0O+
8JxvwOxBPxr4EHdiUFPgwtloiWM5MHIJ+PzCNXn9cU7BjVPiVdD7hwkmp1JPPo/3
h7ZEh4EsrnzsmvlHjVRCp7RnxgEMoi/tWvTSOT6edskW7ZLVQq+9Vim15RETA2zV
/PwpdjeUOB3Q2FhBgkDtPlWLyQ3dcHA0gb3zpcGI+MlQ9hbgw73ROWHHlxr3JOUW
bS89iboewsnygc411CAcK4AmQ9nDwtuSwM6vg4533p+X8EFgYMI/IGh2oXWWRkSp
WVKQDDTx4OhzPzeBuracqbqfk2JoGl/L8PF6fv0GtryXL42SG9YgTEgKIgvZw4mV
/MWNGgECg67zQrHy/wdxHLfL5jz6844w0qA6+kYhIPFReEZxC5brzqIFuXv4Vkvs
wN4cVqkBSIqygmyRXZHIoEXIz9mo2xeYUGitGuZo38cnXXwZ4nk+qZ46f9XZqc6z
HKhbYQx3gRUZwIQQktxBK72o/NRw9U3ariD9CJ+uaTSbS0jZHk9ZVRg+rcJAhr+V
GgYa8IfolM+Tgh+6K0i2LtKKKr1uXGnlX7/RLjBP/8x7F83ae+08AKIwDsqcz/RJ
Gh4YKJ9c7dypqCYJpWpU+mWJ2UyJCzsemcOOzhz2rrg1K4hGeiojAxVI3+jObQZe
7o5HnNZJ34cDu93vf9tsYfcHtx33VyzeQa18FCl1Y2JP+sXq+xehVfnWJ6zAGuHi
zRIq+Gtm1ZzCiy1/wLOOpnM5+XBw0dX6ccImlwirlm0ajNAoPqX84vQtfOSBeKU1
tLviFHzPmpa2BY+7j39HMusr1AfFUjqF2XPJ1TnHmPLTHJ6vn00oC58ECP8yoI1p
ajtLYRCi2iKozF1VaN/ygmtPPy+8TdxBV7nFUuw+bnpn1Vcoi1JNV3NFhKYTNkbI
h+heJkBXVDjNgGxlQ4W8aqwhDGZju3AYQD6HU0Da8a2EiCeoxS0zx4S+nHRFHMpb
e47SgdF49/WfMlnB62NJq8xxb9EVmK1X57O/A1HwZxbgi6UYcAqlsbK5ojTivKSF
rV6ks7zKaCq2E5mq28Ihb/n22YqD5yoQeeWcuuyG/urmC3REKkW6WbWUfhe8svkT
3cRFe373BYU/gkxTRcFFTag7Khrn/22ptz8nNon+Md/1Jj8l1SN71t7dpupa6mBm
q0e4Iu9laFaIT+I3/V1isOsmwYlVZ+GDWcYQzYjmcZWCiKdexmhZw5Sn3f18+51T
TZWW05CP0uB602JBvgyE9I9OzwZgj784drAIcLeFhIe6LYEESbj2n2CBlUwXJCe7
L9CHC2d8B9mSk9hpR77inHHa+Eh2Bz6iIPg/xacA+4c91F4Za1gYLd16jSohm9jn
lHUPu/bQGlKE9ZsA1Lc1TevThBghp6P+tT8G4mY2HKui/Ds75B6vwIzYFw1gRs/y
qZok2jDpEtUwUaKD7OUp5C4q+IvvFz1X1uU4tB1eY1a30e3LT9WItv4Mva8SkAfO
WBl4ZFcVHBrDFXHEigs5OGrR5xuQj5aOW5NPrTX3TmsK9TZMen20dIuYObN6tfKh
uUf1I72yQ1xHihtl5MngrrjImlU1BXTXG+xqu7+p5VDh83xUAye21nvqedp5aCMj
lkBDTkNSzJiHKiSgqTa3rpeNRF09YD10KmyIfab5rtb1t9WqY+CFjC5CFUFf+wWI
+Un69OVbQQIgbz41A8E+ogNnMvZ+NjclA0bsVRX9omYY9TlkUezVnItCs1uKgoD6
imvwtFUZdpheAK4RBXWe668xk2+S1sE4Yl3YQrodHImHnv3fom2Po9fOQlumlhEJ
ahXA6TE3qTGRdZrLS7CwZqfail/DXiH6+dzzIqmJx1IHp4xHLa+Fq47WD3Mgantp
qYlfP8x4frwJNE2i4bwCnKC8B9UjBy6Q7PTESTMx149b4gqeMLhpgb2q48mf7oIR
VNyZ7+L3V+VbSsCwMFsdZHE1FBQSWgawfMf8B+ziD62YMcwAzcE+T5FJKcuiB4Wr
EZ+SfBdmBX2BV2+MW8hs3D8cfwM6TFtYqOHhfOa7ZPgq39nhs3RZIwEUr4woDrvx
rpiyH1bMvBQSEAhXNabJ/veOzq2giZKCGmf4jrSTpuhyfU7Dmvw77BVIgv3Gxvsd
hLCtdfWmFcz8qWy5bImC2wXvZfjboB5MYQD0S6I8PHVm3r1L3hi1yUO+LRXd0FOM
BSC7sGs30pv1hMTsMST9bw/1Z1sndt8sxyMy/5CoOHUtATf+2Ti1yUYedfIlUZ0o
G6z7q/Zl8X+UjudWQSSCbPPPMPrPcSReudzONc5/Ii0NsR2AKGU9I5a8Uef5OuZ/
P46pZTqqd0pKZeb9L3TyUBspEPdnYxovVEyEJGqyc94+kDVG2yzMe3dYekcTaF1i
WQojXkal3FFzJJJRR56jc2qJUMc0T7qYAJLT5/Efpjluv4MDzot2CNbqiQO614h+
MuJjj+GJITpIvxc8Wb0bXBdRQy5Cl5SdvzLBtt95pd+V6K5WByjmGxw4ExZdbxRQ
Qv87iTDb6ZM9ylrMBgQPhnD4rs5yjs8bWRpW9v0vPVZTlmPct6Ab9/mVMwIP1M7a
nqUXshr1l7ITUm1yq0FCBGZttUOkdPrb5lrH5CSOwAswevpNc7Ax+jijGdd0L5ti
zYbelad2Saht0T/F72sJHhLkhUeoEas0+6y7VrMb8qIXSaqjjWNrxqaG/xd3L4ok
fUaL4RgkqpkBOYTSVfXUHp2nVg7NEJoMgM8s6EAnQCD0AqK437lJJ/usI8yAHvxy
02T6mJriOUBkCLxfjlNJTVSoMQJJoGHrWmo97X4hFk4GgQCKbpAq2RbMKP8UOaPn
d7oOm9TWmkHW8pKufZY+FCrEtx0wco2eiOCDNHNwHEP/UP2SY2Eh0dQbyBJSe+8m
y/KqEAwtCcQSnNaxW5cWigy4FuuIkw+yaSnddZLlzsD/KQxPDktlDx0Mz1G3v6tJ
hE7P2uIKsiuQQKqR1DdcAq0mvr3fugQTISDSAsIRAnTsehCdxYtJojZ2PvEsrcxD
ykzATABPKcPeNl9LY/EbVNyJNhg84gmEeHEYuO9GzCDBRpJTNiAFfb4QQWQmSQ/F
0c7oxqqbic8KTnosFGDmz6QY7o8R8O4+IA1mB/+/Mzlc7BCIWEniWiJp22Fhka5I
HT/YXmN6Xh8+cADhEIN7bO6GHp2aCK4jgcBqsbYl32meS8ZKiPNQuv5BvyDaWljq
E+jy4VHgzHAaz0Er0GHz02di6fcBUxn7AbA04m8mDifoQUzwkk774XPxs+glGwSP
m44Kou9gaKsPOj6WIF4ljBe4d92HmAv9xNosno641telI7v+dmmR9pBzkTObwfPZ
c2z0aWfgT6a9Qy/ztMCzzSViVrTVz2ZrqNIJfjxDn2wx7xB4Wsx7Q2e9iL/mViF5
epeQoswH4X5Bro2ofjBdIV2ST8SO4X4W5ACXK1mbN/hJbCQKykm/G0zNLRZv+O53
Phx/B5fCpXlP2pJh9nuSrm4mDFzdLftdyVE8ppepbyxiDCSMk3t4il4qwdZmDi6O
7WCmZPTuGo+YYzbp0XbBpXno5gJ9HYAeZXewLnMJqyqf5x5ERn/nKsHQaTdk+nKW
ZYZ5k1mFXacevv98iDIvLjnkfnJuf1SjGMi2/aycRO9bD2Er1knmTbCBMw2kqu+G
XYSwwnit0gzWdKF0lJYhnbS9ktqjZZVpBwB98FCoB99VhFOuA+VjHImMK7ePs/Sb
zSKmbrHqdS9p0GY3Hm6mQGO7qV1V+52jWqbQON+2LzV3v1kbmVWpJlB6T9RcqFeu
DGa/tss8aorTQ8Pc+WGdGEGi34qJLE/zTbNmPTrF7XdUDs7rUZgO4u54SteEw28X
IJNyoD6G2/rhhYlrDT/6UbkHQlmJefl6lxriDsoRejyUShzEEt0lHJgyhKFkbo7G
GUpvBPZuOrFBQMcNrmGe9czx1wp9emdhhs2CwqE5yfk6+KCawhZPr/Xb/ZTuu3Y5
G09FPhVvr4nMAoHe2s6dqX7cr94hSQeR8IYoHCF1LdepaSl4E6tvxPMJX4ul9Nyh
Pb5IXZnxPjTqg3q24q6Otlx15xYQSEy9glp/GFgNtzHwG1LOR9xNoiZ/ulLmPD63
WLmEYPJ3PE99kWOkOV9r9SJfclJiXsAnvtDA49/E1slnjodJ99fNYlZZQKsP3PO9
FmZXsAlpShrjD/TaY3CCEERWv1cd6SxZ/U3lrXCJJsJV7hov5buc3ii+AL1rFEuR
oZ9li5gPgDn9NNeu9oEVQQNoORT8KdlgYCXHkw/+MYg8hV6zCfvAv18bb6yeESjx
nozgZqV02NPcIhmzPpz2F+mUVfZvwQ7e0oA1wRluU4Xf5v+Fa8EkjVus9M+01Ivl
btpnUvus6/7uojG7gLCsFlzlDQ0QMoCLk2qe3CR/dqlTC6FvoFfm5CuFl4oBRexv
5bUI5EDrK70iV0ETDWW4QVLStCDs9i4xkAl0NCp2ed/OgYF/vw5XCGy5QPIBJPLW
tMsIRy+Lz6exBHtbxyeCwWpFRo6n1bGz1HrQaEGQeTxMiqDVkdzjq3rJVZdXa/w5
CG4GGi31e7rNmXyXZI9GarWIsXB/vrE5al5RTuGETrGKU5Yx3nPel6ar/k5ciDT4
4WJB7PW3Vm3X40fr6pEoVUAxItZRgq/SQ1bZX5p6GRR6C/mYDYZK4QAk1I35FkiU
x3NoP4y+86K4UVvM/VciAos0LC1g5hntdQ5hR98/TsIGhs1xLv0/7bFDjTj3XMV9
GC6p+hTnc0ytxBVcbgR6HTlMb1WEM3wuPas1UeiZN1lYIIXBqsPJXUO2aSSmOpSp
4rn2KoF0SswmRIJl+UZawwlr4++Oiibxtmlx7qvnzqhr0n7yucHQ4U2Vbrh8AKOq
MnVs6dEKoSd09qjzQ1cB/MGOSBqkIZEAdcgsGprwWd+rNWFoO3iwYamhgq7DQ9mS
8gY6EEtn9HeSB2huMhS4SVcm8JFUWQBcNfrSsSVoq3C24lFQeJ2Vh8WlHcnq++Mv
WmlXbXuNo+GLxW+CXOvROYVzFR/749eny2VHpqQ9RP5ldQABiKauoCsY70RVKUPv
UCBG/TzQb9tPqSzMGIL7jrZoJle5280lD9uFwrKPHn0sE0t2U+a1eECdE3iUjzkL
3rCn6MejQ8Ndr70ER2qgjbJiLT3M5cunlexJ5klvg5q0LRF0ibYqIk9daeXvyAY1
hdvCMSY5t6LYW5g5QiDbVnDLw/iqrpIIXiztod5Gux8s4YJ4eQ97aVmeTyGBaatT
gYdjeMkAcUqSy8Bh/COZ8WRya//udMlEJSPeddqiIDEvRMpqhzQGzWnyKHScA7aq
kQ9ioY9c5s664Y1Q6+MBVXDWPcCntYUEl7GxjPfAxGK9SjXXFStRWK+8ROkcuwhD
fJXKtUKrk2e4bIlITyvDkypGOS2NxBhyoa0SlE6sDK0ElPhn4Nr0m0ynx8H8Nm0J
Jyc99Bv54nBNg6DeBlChZGU5Sib7A7G/SKJ+vz3k/hHGVw4c+dy3GlppsebmiVvf
OBDIms6avuhMfqgFpaYSNPNLvvUSoabz89bZim8yYNWmeGQminTgqex/hgXSjPh0
ZgBeWYkFMlG2ZFlz/OkU7kPBGBycyTwt5RkH8Z6NRqe9b7IOJlX+XN8p+8DAQm0B
tIMT0aGIxW0M9vbrX5dppkcF9JQqL5rxzV+MWXQ0N+Rxkg6k9cZkXjxXcVuXGIoo
zGCoYPdtWCKvwlWHeGDlsYajc8zbusblXIdDallBtGcnFhCLN/YYkpUBctBfhBUL
82PfCe7MjuUKM0pMgGj6cOipP4GDHtboBYvEXSGVpCYabEfvh5mliwL5c9gS1g3l
2eM1YcBvCQkXvToUajvsD0lbfjHwfJUtULVhp1r6Fwlr2JHUsp2X3B3DHmccgBYS
etdl9z8iYmTy1O8nT4BP7MHH7R7q+qyLy/gR3Zu2O0zR2okxA9xHBnHdjvIzDdpa
MVjfsYzkxHFd9ISICsEYYx1a+1rVCsxdspwZaiA5fUI4h9y7FahE4/aN+MWlvVzs
dFp2+vJEJDoov7LtFJpK8auwPPSTBiabXIXNEyY1EukZTTWShqfJkxRRV1AffmL0
zPPH4oKcv+yLM2bhmLPF9a97uJ/winfg3WJkQssV3oehXPlxUF8xSYsUfL4ZT3dh
zVhdP7Rvp2cAUYHPFYzqvuPo7MQ0tco/I7lIIoNdIPcXa7F+vy7SKDUFc2T/fB+/
p0UmyKZjXeYFiih79kAiAIuMxhpQupToP+kYnXA3iBUeOkKK9wzns49ZOateNINv
Al8wOVW9Dgrabh1LfnXw2bqNaBoOEbXle2p+Nh3W9FOfeKP98MQK0HlhTfn6Yj7i
5v+KJhiMtOW+vF7MaLIHZEcydLTvz/e07e2+Fh6fAwz0iL/6UI+LWX4tY/z8ijhs
K8OGO3zg75nD2FKvMB0XHFF1KnT+FcixQclh7oHVeZ7wvMN6Yov9N/n9czD/aL3R
GXRJULuzc5rgUoEYAKS4LgaoZF+l/I6dCJH4Yz4Wt6jQjA7ClPT6oCuHE0Nkxtdy
NWEhTMGclg2cbvw9GAJspUEk7fp0AE23soGTbRfRpMLLHZLa7Af6o76QUqgXopKw
ifVJSEXIlYQxZ+WcxVo5KaZm136sg1eAKxGsVKlX5hHfsXWoBDA6NBxaMtTN1/TD
HnQnpKRJoqk75DPUSvRI3OeMM+G/t/ACzzlQJp1AG+6fO2qvP233+K3aRx4A4iKU
81hH3ga6/jk3G6OovoHLH7yHrbkJS8XdkpsFcPwD+9yW1Y0tRD8EsfTahFUbxfUI
g3UcTYzfR+deZMw+LaM0Lfof9ELxAdYv2WiOA1vL4842VIMbxJguYfnuSaa/soBI
irgFhgP4BTGyXsQaKYZI8S7wxoWDBI7l0xpNc/4f+xsFdATnAljzgU/M5STTK0hP
oeiry1MlSZ61c+7w11v3MXHar6+jf3MuHuttGKNg6aZwveGg0x40vkg8snArstXL
dHuUjqiQh9i4s+hk+4chmT725oJMPAGxWeuUgNSHOtV5NCXavJ+EezhOHA6Lf5HN
fVNndQYNKnZEVk/ges/NDwCsiFYnEamgDgqFu2XCbeCae+rANcjvst+LGO0d96y+
Iv1OUAkGy5zxKiUzym0sXIOehlTr2HbFS1HfgTPocoH90XFyiK+tBIvNcLoY4FzF
PU9/2DpyvJJvQWgVVK9SPkOdXuMlDDhFDWQyTfuxCnLSYzo3574rwm52DDh6OUpZ
eAL6ymyW45ekEuDsoEQ/4qw2y/S3PGMpev14Zens5frojq1FFdNzPTiyMl1s43Za
wsCW9z1SHBAP+1a4dehKetwXJAZhrpFR8v7kXs6vy1mzwMdmNjpNx3aQujRiz1hr
FsFzivfI6fY8s5DCxB1tUuUY2y/q74TDIph6HcBxEDbJQAVnjEmnEXUe6fxNI5IX
iXOP9a+K4RcfruaZ5hxjiyS9NPIdahAK6vkhz8m59QnvVLOraBbnFzXOFHWva87h
57fHwisgLdr1mP7+H9O4Jp0ex17PPznbFRkNy41IiKzuxucd8xh8+Ql8iSIyUjSl
ZBwM1C4a15uM4pVnCpq6NWhYLy/5xmRGWuDBWysxTZDpfXfyYUWy4dIbwsYycBiJ
axeaCUpUxKuKR+HgrXwZN+imQA4n8JiTzuVhbsriopM2WFXz4JnGsHqoBHJfabev
+bCInfzibKuMB8u7Bth3AWim1f2w1dAF8KrAkYLIitTAK6gglRdPFI/fJHDQEwO1
fsppT10l76Q264z5QePMql4LohAXFpHUB5pTjn1qGYtNMyRFtD3VUe02VPDpU0wd
372N5poYw9piePV9yn1sLuehwPfr9guxBAcfc0dtc3W21V5xu7yWRI3SMSlorG90
DZh0/t/b/C59Qa9kFMzloOWdbHbnp7ls9U4yo1uQ4lEMf5hUjT/tDkwWgtcztur+
FekeLPYB7OGa5Fg0/2et0zYTfIjPQjBAPH8h5DWitf+QtYbumByo444vC8vP/SRH
9F+Za9NOlk3sr91QBo88ZTHEDXtdsQXZotCklMLdQJ1YIgTTyPookdqxnGEsfpph
5pqZGCIRGchYsuUXTwGCRvDlEbru2I2O2LtkzSQDPjNiXWmdBqWllafMg7e8od9p
9oaGCXMEbsqNs7hchZwBYfM22Om6ONuuicIh9l8MVGre5LL52J4CzwDFzxCZ4s/P
9qOMoXCQxuqTZZ16qyIW0G9+akvVEp+bWMQhv2FeLXN2tPcrxHe8wtZZvTHezBrL
CVqRyxY5vgBcQU2lsttOzW0ude/9Wv/A2aVluv7v7PrdPaSTvwn57btUANkTFBL0
kToZd5PtGwu69WJYPXdWaEebffoSC/zC8o9vdTDHALE1CNJ7ITTg/sMcCKa9AXtB
g1IeAtAnFXKWlICnXN6VLcX3M7NRFm5QVENU4HTsYiZboc4xLcxxS57jGdiFulq/
7fAlhhxgLF+a5yMJFTX2MfzolmrsZU0zv5aZwTBoV6v/zPydhEm3CPGr5egZHwRN
XFt142w3Na1LXsBAPHBgWHnECPMypxAv4Pp/HYD16tv/bhSkSYrtd/p0rYivT14Z
U6mOr791JW0wxvoJvpm0NpgEbGxCH3h5EcfyhCXGKeYUEu29M5TWFVXVN5e8mRt4
KWVYoIzkD2J8HLrVnT9ZgNt0NYWBsLOi50YEtfQX3SjUwRvyZiPWD13t6TL99vz3
a+42m7+deyIYVIcWyhhYw/cyOwtTd2GRmHf/bV3pVlJip3+HEFtgiAZQiGxUs476
vM22I1LfCt6t/3qwPr3LZBhJ2N3MKuE9wN1ULLY8jqQA/ktJV20wYOFF0gcIi1kR
mBwUi+Qi01adK0VsdReys0+kwk2hpYr+VXHplJwVHvjCLej2JfjUVHkhTchKN95u
xoZ/mSsZsQPfDJWJcJjtSrFRxNt1E33zJ6Dahiw1/4424X06CeKLp9aoUcSNJ69y
7VkCQkJbOBHm/NgubtBoMWhkaJhfGSmiHg9PakceBdsRe1m0+PvsWH9+2I5lFgdH
fmXrd74ViebAkAdQsQvvgZ3tpTSDtjE1beoLbNero7u6U8LOIdl4yvixHJjqnwmJ
0CuNuLwAR832I3FXtUsrEF1KzDDNW0l6pyEeNoXGWzcjJXY5/fMn59SdV66zkc1K
99/QRM/24QpHXYnDyCExpviVwPKkH9NYa4bmAKe8aK2ml7lUDkeywtG9/o9kk+2G
74/WQbZPaWksVMsFEDFh746SSKXiO4vmlFALKD3VB11D3doc/LrXhamcR/c/iGhw
gSJVSKcbu7U/t6xfQJpv8nzvdnG9s9ANBjORe4UDIS5gwSymn7J7HgIzLc1LIszP
rNhh/LMfxIwP0JJa18mN567kolWxKr8EIFCp1nTNlZC3uYXZ/R2Y1rowkF2vRrXU
w9/A7mOhHniyzELle/X+dD8dK4ElaH29p4PzCvvGlJdd9vFuQbji+hGL5X126idm
dvqd2esRsNVkJxyFc+wLn1MDis7C0gpdL6V/bMyX4MUFOuatgj/482XOIaLQKFEy
lS7XvFp29lCskrMH1iPifWSdL7a/HvVl+MfVeU80oXmDaQmAdd44pZ6aI2aifi91
E6Ksl5EE9uZu5ooxlnhSWgtbiW+aIbHY19/Zdt8TMA9oURqJqF51WCCfp84m49qO
c5e5Q5sBvU0ckpyG3zejLvDl9nKqeXuEcqf7mqMiaIZb/ay9bEhghZmXTMrPWnFi
HOjrbXLFghiKrYBxavfLV+IUYVj5cLTzxANdIe0GT8tG2R0qLQCvbk7+XKj3GKiC
N34ACfyR1vYuo7MqUbTM2yQXq096BM7/UNjoXQ6rpl93tS+wgHrwtFf3va0VkCe3
DxdQokWVWoZGyI9hxJqIHaDi2nvkpZ26JAHepgLFSWAVT03Uwa9aTD0n8bVdM65t
4aVaZTJGOfVo8T/zYrR0Ts7mQF7DXBXylh583kxDIccl5dWfElQhFDuG8coQ6wvm
HRoz7RfuC1pGYtMEDPS7jt+2miAZB1M1QoRkwtHfW8DkWsE416HBlFmwB6PbYEQY
sXefjLDXh5+lHhrQazqnZdisLHQokB+mzfFGXDvFUP+LSN6ZyInSubAWte6sqrcp
nIEz3i+FAyTumh/gaPuor/AHeQfySXyZ5CgT7azxcwzn2x+G/gxhy4F7fo5RGteA
Uw9RteftMDfd2sReUUWKYmSzcXHswE0IVK42E1vvgD117vz3EzOQpJuAaphlAMcr
hLAEKargH8Odcet/Drtw3Bh6kG37ZLN6BIRKHt+j5XFYEsBCG1m8iWItb4IVqsIb
1qwDS/6j87V7YSbyT9J13sGlfVSkTltB4kGDISGD9kHgALtoUrKJ8e88Mz17bE4i
M5RBW6opJNtuvivDKB7BC6zC7jIA8m9+fuEG/MkUzebGFy+HURsfjm101XUZADyF
wtJe4uiA3ZsoLn9cGGvsEcEjKtedQZiE+nogzORXRnaBBuk8cXp9etagxAQE7FtW
jD2JZx1qxizq9xdEl9DFB1mtFWfT5Fj+I8+jMQ9AXAZhLFCkkfI7fafZUyzTkcQI
BhlgrDHZbqD+OH680wu7XMHpNqdzDBfcgebznyiU7GhideRBez1vUd1OSa8DjWSG
MTwg0AKYufvJxDjr7V8WioYXBzZNKpSO1mGXGuAoY8DvICJeQAU+UFSBAkqTRwga
+xjJbiMa4X3cqgUHfBwu26HgjiN5EJ/Dpyj27Lraejb7jVYOiGaRPEFgapWA7hw2
a5/xU9WFHLZhHblirFv4YDmi4T0LlCrUFM1duPHVgcXEq+bt+UdyVcbgNXWFYtZ+
8/7UXLwxislFzHtwOhDMmAeY6NhtyN35AmESgRO4YmGNQk6zdzFhF61AWTe5Iio9
FttTIsmVaT0DRjN5c2ipOczuiEWCDH28S56wpLvHX84M/8fLTlVXeDUoTeFw368i
skXEQ/mUuKl1vcbZ/m97kdzTEsQB0Cjvt2VPjwyjbJPYznQ4FlQanhm8JCKli7Y1
ZfLxQTEUd0eepx630MAHbuela6x32X7Kv3wcrAGDjN47ra34yvSB9cRwJh5L3jvn
tz+ivvaIRjaSHKQ1yBHLCzUvyrfwIEeT6APGfQIJsSks05CowG2aq7/tQ5se7ukE
BOi8CSYzm+iuJKd+xTnX1Bk7IU28d7aDpgxKJydBp9xtw/VaiNQrSbfmYb13FuB8
S0HOyDEHncV+66nhz32c96dPMpdV/Cd92CJ/o09OgTo/oyDaXPNwGsTFg4MpcOR8
QAcyOnUVEjwERO3bSvXodsAHTNfs1lmdb0Tw8ReXbJZCQiIEbrvCixZv6o4gRbe/
jl4GKXrAUr0zbr82jswHSHtCwz7R5BXEOkCZEuiIIRNjdBPa6U8syZfx3W4aZhne
pYy8Pqlc7Rp5d/Dl0zVqFLJQq1qh1J4nDVtLSCxP6a2g27Yjtka08tVltoeRueFv
119GiqtHY/o7gpquNHIeaMjrRFB6iR65lQ3oNz5/+AYeDy35I1bYamAjt27uVVh/
LY9+kaKy4i2qzF3F2Xnec6zHjG4lt1OJZ+YCX8RHaIW8+IKRNSEiPPd2W/rNdFNX
Kc5JsRpelv24vBgIsXYf+dW/UykwCuuxgXmenwPz1TbFdPzB/wCds7FiwZ7m0DiH
2jUl5XOiHiXHey4JyXx3Mg7i9N6Lht/9Ulj2zMvI9YdLo5daCZCYTfR58kNoU9jH
0SuRWVJGp7sqowi7jmT7cxKmeqvvAVkTRrg6Rn5jEhGf32ysg/dGNP5W4Yn5rfHh
w8oPgY+4TU7J+/fK5C630Vs+F25oQk3/gnBGDrtkFyS7B6ALCiNTApvon7HGvJ7A
BpMMQhWZrY1h4InfUVPjI3E5GV7tJR8KBbfFpTWnBsjtNbQjUwTkPM1xUsO6tZfi
lQ8czapOtPqTmJE7QELxSgNKS5WmCa5cezdSMiecGqplfapPJanb/aAY0ImwAX5e
cuhZPwNYZqHuKMiaJEV+7vgg4ZXBrG+chyr0ku2AiFd5xq3mNImh3ukeyoSfrdKU
wmNPLTmJ2M2TAz2rx5Pkh7tHkTWscQlpuIH7w4y+tw2TV/XKPjTCQ7CfCs031IX2
/O3P916dvK8g1rwb+sZvckceCuVTFQ4HNjijmnVeHC26kaROObEyIrHW4sh6W7gQ
iXPHSxrUo7ARwmT+5BQAgZhpHfd3QL0SmjVEd7hTZOx08E4OxpmCvQBJQoTRf0XW
tysyLLrjRjMTyOwD6C+eICzaujQrrHkjI8f25WjC1fqTbq4rRJChsIbrLVxzAS+s
HH/L7gDk5A/C5i8k6zB1d1L6zyWMWU91/Y/T1v2zmZZ3ILvcAKUWhoCpwhD7y/vI
O2Q7kQfhRnrTkWgRBiesPJebq8ld+L2pUTB9GGmWaU/Ykbte/e759tFM0ZLxvpYm
/xQ2o66ar8wp49jj+h9Ep1EkA9blZTDMThrPA4I6y9jvbgYRfoMavPKl9Zt8HHVy
3YH/wLbh01tRB9adZ6KmTVmERvFcePlO8+jfC5f6QtLTITf7Z5quj2jO48J6YLuz
Q9EDKy+vkWjrzmfrnoWM1z2YH9Mg2w3+QZbXXHTqVb4BDhOMsKHOKYTwNqSXP2cS
YcYs+9yp/kIHng+AQ6IWqxQWZpvIvxqd2AMI9QVTfN4DdaNgEdoNsj02qx2om+IH
QzheEi+ks0zfj9824FOQ3orEVPBMX1XZ2y4pF5z+NFls3UQJ4Tu+z94ldxSzNShr
NJmhm9hgHpcsQwIxdTPb3o9pqKbxERjXE6chz3wvuMVhN6VOlYq1RH7GRpW7mjc+
WmMZ9OcSCqk0KU1/U6m4k1/bwULQtngt3Qc2vbPJucr6Md6KaFKVz9JP8ycCQGZx
BGeGtDfdtb7ISJTZxPGZZwowJvBRqnVCZMwKWE9SDU2yle342SIZ9liWoBhZQX1W
1DaJIXvckXiyeynjyyV+oyiOCezS2OlXMGVrkgkxZ5/530Ylvg0aGgCcQbvN1Ph5
iaepqCIePvLij5/FHFzngC1W4ciDkfSrXgLp7Cb/8sLIKk6euddgIPCa0kZQpzDs
5rqriMLMfDQkWGS12kIgmcbYTUUJVHom2AtSE5pHeUIMH/O63Gb94CCUNev1VZ7l
7o5xdq6gjXTTSXZcOqaJ8YatayLKTaFicZlssFLtTATZjBtXK5dmI/F73Lf1/koZ
dmQlvPdr7qQOZsx4HFeReWPzB5KrfZXMRz3hX4XqfegMvUWCS7+YNgRQ/zLgj1HX
MezYdb3SH2zreR1aJakW0pCzz7mkTX1yQCBXgQ6C2f1dY8G7eJFBXZJBC8gwZkE1
5ntwreEbXo1ZVuQSQMHkJ5dqq/cNpQdhzdbpfCcw/k7eFXwrk3hPK0BQL0nvTVUu
yx0Mjjn6SDFDYL112JGbDJTwi5UjbYEtHjWS1BNk88lQotxrkBigyz27oFVC9ONO
u210tMiB/ZbPm1ALqXaj2NcEZKsKmuDt2kd2B2L8xZiU3cMVV15FDxhn7YZ+4+zB
9ALvRIyfBGEKtZMI/vqlG2B8OfVxHzP6yxmGdk2PZkbi2TlhK1lck4ndDJ+VHMFQ
LQK3d0qavwNkmq12fmfaOmQnQ3mbXHWL1T26Lt2ABmnVBNWqXbuHwfSfuNTtzHAn
Be/22UO0iMSHhP48YwadQXDhJOREOaGEp/Wt/8p1iu/hj4mZ8OnWpbwZ3Ljqa8FP
GDVXYsoLyLUTv2hHDen+1lQvQRyVv1UYL5qEpgW1JYVoYHIESNtCqjexAj3ofam3
fDFfzmVTDs4nGqq3ozbzPUw2U700/qR817xImxcDP3U7PI15IDLPlFNrfbkOpMAh
40zAejF6AMCOyFDjqbozbQDDKEkKKd8rY6hn9Uye2P1V3wZTQIfuhAq8TbCTZ2Z/
pxfn7RDmD1y/h69JLzb1CHbrkxV4ZUlILeWWf+h7bpjzSp6Es8wwgjLa0eyiJZK8
1GmiPO3dmGhq8vzhgT8IR6rPE29ERU6fsXBsMXePTbLa6L1VSdoORe7Z68X/CTV6
B01cxV4u9Vi+mNERuJ2AXWj3SeD6rDkNIY4hg8YYVxwfOESbxZqjfy7+8wRCncKo
wlr2ma1xgChciT23p16Z30KOsB8YuO7r70z/Y9BMhYJdx/tEumZXfRLc7iZuoNuu
baIQsFHbI4KGfU3TQsSFoWckkZRuxf/DLqVTfg1lGfHHgLwsTdp2lKa4D63MaHMv
UAN0EeOTRXdWX6H+D5zXMX3KP3AQ3lqi2qFoGb6CV1b5i+bD1yfF91g6xNGZjYkG
0ZiXlV7s+jLPbTzO/SGJ48OXdvVGqGmXHWi1cwsdf+8+k8Abg41qQXt32jg7dlqV
bmMjChx5Hh4Q+otLBFpTWxpu5Ci926nNSi9d4CsJUr3LeVKwgZqWiqTEEkvNRGWX
Sx9dCE+QIyoRSem4yLmvcjSv8sLSdqhI98F7QBFY1yxtirvUUMyfD6d5TkQsxPPr
CGcADi+u3XJl1z01BsqM+YD7ux276NhBvU2b2V1uGiKWcJbrnSXeHMcaEdlyXltr
0IzZWwwHIgPKgGGsvNPa5ZXGMtkFIN2gU9CwZAW/vC9+meb2pJA9ZUiF33FYMxa4
PFunm+WWYX3crhr5MBELB22okcbxdUNwza8W7yF3KDO2vNldJwQs5S1yjLUaVX9m
AXtCCh4ZcmstF7MFu9MXRXVCNsQENrVQJa2gp/jwnrgQL0hdJoI5HY7viAMvFO8S
NWwhePG20O2Ym/GYBXdIR1muzHGFxvd6bcGxArHHxMNUO+QDeeZzS4dOjzKgKeG2
snRHLBIHg4IR5j/tCmpgm6QQl9rXWcp6I1oeOg9J7uJhzmc/ZbR1VhhOnTgkmWog
1Nq0bMwhT4wOor/TxYICoE6OuCh2vzgRYWsMjFwt4nGBE0VllshBaHmu4nHFaq9r
dHQBFibFkZ4HdV1R1Ygv0jReIBdxegk48tvnyVzkhgC2SPs1wFcV10Y+qdMJNTXz
/aro+g93itqMHEiMsLfLaavzY/zJP3uffPXTA6yYuea1EHUa/26g7wfmmoHQ409E
jqqJscexZQGTzJjTAJ+y6Ln3x2d3yImi1jDZkM2BaaTCs3X9P6r5bSBfmewP3g/b
QESK20/wLfjubtZfUacT7+d9E/i31VRGVew4OsDM5re9xVVTzpp9llOtm7nvNciZ
2Am7jbQvGKdLlHbdw3rqNKgmufLqb1JfLXr4zAYMDEIrXZVapQRO5FguXjh9bdnq
9JlccmUuTNX/vVxBvM5mtDpR6Sd7f4G+P+2Zrz3+igivZ/hl0xSUVJU5YYq/3/hL
DL+dNy8uCbmDrnZKPDpvJJsyQ90zfzqSmZoZw7oNQDb/gqZqUvkFqIcoTjU5lCMm
q8I+VvBnF6tpJORTXeC7buKhytzvAdSqZC0x2U8M+FavPM9IL3GccHRkwcAYSV7c
xYOCik3O/QbQkx0NrfE2uyIRrFGZWOLLQtiBc4qGD6Lx/9yf19bku5r/ZLMFxzpX
J/FfHY+Rb8RBc7qrGtV7BHsAOIuNlG5lab4ftBWHa4m/6asSnxUIx9/DzN0vNXnj
p8hTb8tqpIlQAQwXKk/Jyi0tXd4A111KZzBOBZNjTjz9T5YOSx4PZmf+1EU91QYu
vdQlLrCklqPlH+HCNpkm8SIJgN5H739u63QiRjKXvQd2itf9Ks+RW/imwvKPFU36
JO0T6zlwLnlsxPEJ0V81ofwWyoqbeW+BKUErrZ5JKvEwyoTDD20JtlGgIh2rA3TA
7gx/hKvuiltY2zhnLOymEo987yatI4LzzoJan87KR9N4M8Gi11cQZMPWpeRdZfsP
qc6QJfkZ0pq3h4TzTp83qtYjhRVzR0I9Cpu/c80mloPf4c6/GaLZwAwu58DVmhQ5
x/ymWGWPCdU4BHd98fM/Aa6cX39dk3Zat3NwmNls1/l8mXcDoNkgPUGqCkpvWcp/
J49ZDkmvaZQeZacqYFvdFr31ZFx769G5SXaaCQSuaSdT9xCBMy5Zn+JsqUks7OUG
mMXsrClUpwW6QFg8LOe7q8M7Ydmk3d/PVATFWFm5zGYHYQwek9cAvuki1jeFg7o+
Qb86ZbEYZqyKZJMsB7711KQ+CAZmz20iUMiBNhmp8+Lev3ttwKrPA/uCqT2K8pXV
6SLb4AFUc+SUijvbGr9eDYwBJAB2cgFzfHqIguQ+cw84ZoPEg4tGt7EP+uSHnYPn
Eh/h9JiGW09VA1awRdP8wArB5A6PINorIA8y/1TMNa2cDYGJSAz3Bp7iW/8/sMRl
2vB4SpHbDl153MC12XC98IdWjXy+2qusRV0w5kARPZ4VpgciL/v+o/hDVrHUR7LL
uV/MVvREj8esdSHn9jV4h2I/ahWARrDDQjcprHTZ5yXkI1PAzLCIDaBlTyk5C4+C
FitXKdT1DaXItVPr16OP9DU8jn17Z1rPoxrBN9DHriqDrRYw5sYhsxoqAmK2d3Lw
zdlQSNaQYvUO8A6O1II6Rq0niHG+DX0m0yRUbTsn/onH2XzZP3BCHaYcPunwjWj3
Cx7n5XV6UYZYbf7uDVjKv7nZYNptWSP9N0bePq/kUQrhbgPHBlwF/uvgAhA504/X
+BQUr+oHxIyQXDGmQd/4/thhL+Y7feilN3s17XjX9mXL15iejPJsgX2mWZ7bFMxd
dXAGlWHymvjLLrIbhk1bwE5ru4ge746YfFjQbn+IkJrXj4w1x2rg0lmTsvVi8XRo
URQgu1YHoRfpciH5L3HZxDuyXBAQdojZQoEuMbx4W3gGujXL5aWq1Vat23L9otKA
4fR6t7bszWfOnKZRY0sXSUkMiQAJaRzK9qtxl78a+upZ6/PdoXJiO6f66MTMS8z+
g4d1tNoZlLjpAiK8Td0PnFU7QA/N5UHlO0HZCtx4ng7WkDkZlllu1Unx6U8sk0dU
w6Apr2eLouOWgD/OoOVfnM+TEzroE6Ck20vUB+sHnDASY7nkr9m/s30Km/1zQ05S
V3YbgDzv3v3NLLzNKiYQMfOwAn/MtWgm5heA480qA/nw6JYby4AsMLDG987ydp1b
uhJOHu/W/be43+WH0M6LXTIIMEAOaIMr+YMAUC5gby1WFbo1+CF0ymV1mZAUPA0F
X/MITIZrI5yF3Trkb8XBI0kWz9MgwfWQftiMAWy7DuaUNEuz4lS1iraVnqsr9TMW
w8i7422spRUjKQtyKOtNsN4frRsMp+5G40LPTYx1TT/hWWdOIwR8qQPnxWULtsrj
ij9m8AduaoI+2jxxG7t7H4oT44ADiyO7t+AzxPkah4nnM/OcZQU0NjFetFVbttaT
qZdysihQjkD54tPmVftm8k+IpyiM3nxPrudp7HfSI2M9YZO/+CRuMdWZT2tzzn65
LB7OpuotzU5S3J1QtGGeFgnBc8fneqc/4z8InWXkMvtcWGXm3YZ78lHsEzFfF2xA
sHiAb1wjMGfQ2g7C5/EKzc+9i7ouc0qAOGTvgeHodycwObNoqxCUTls8xwk9ONU+
M7UKj7BIhZSp+yVi5YhUwDKTX6FFplZ8AAomHIbK/O5X3PbaxlgyTDRVzq2HjQOd
EZc3YjmZfNJRZIKsuRS1aYonsmzikUKdHCEzSpfd8ycMu0kwVLc2Nl1njnoe398I
yB+SeF0qvqbHup9voeK5zfDRDlQGt3jBTeyuweKDHPxUbhJlv+naAelWIAGlbkI3
0mvdJiiQYqzY3itT1WCu7/mbbBj7HsKclpZT7wV8a9r4OQw125f8PxYi5kiFxaxe
DHq9NhslLzI+KhuIqSZK3o6hqWtBMkf9daXkq12bUuldikfaOhKr5tIkwkCPgSPJ
E/o633MSiqJ0I2fP5xGOQahQqsSE8/NtbfX4Cj+kcAtLrRX5eUqum7V5RH5f8uzx
tDC39P6x2sXWfKW0X2PTWZDB8XwPRtrH7MboxIoxSlIeBv3/lFHQA6QRg4RfWqMC
av1p8/ATJNHH7Or99IdKEOpmsCFcS8KyPQpsnDL327t2K+AnxxqQw2bnUQkGhtc1
s9HwrODDlYMovMrfg5E0ISxeqzhFJHqj2aBCWzRO4IOMQGRULCEz7831fzgYKiDM
C1x676NuuhhzFSSz+mwL+DptEvZSwUWBeBTbsPCgEVf/9DUwmEqeoqsIHAUFDarf
SMHMCULTykSQehjVp9OzFILSValiPQ4l3xX//zVQE778W9ZMvU2ehPucd3Zav4TR
vki0O9S068Brb7kitIP6PDz3lYCyZWL5MWWclySfxUMx6KjmjwJIimRNHT6vyrqv
a5kLM2zvX7MJJ8jCPc4V7LgPmf9FdVSIYMQYwNUz/mLLEgPqHa5VVWZZUac0uKnv
yRu7zBBXGEp8TJlXYEQdaYo8nu5y6PkjiZ+iyXocGpaniHPQYr6+EGJy4MZov+jL
DhCOF0mjHqmea7e/epSmr5fRb5jQaRJY0a3KAymYMTkbDA7h4zOuHxA4xDN2BoKF
YOVUn+s5J5Aw4eUIGnavbGKdczr0hAk4tjISFkgH3yaqSXAtjSdwFPKd3GCQCMYS
PhYX+TNOt1AN3YibU6VZJzPEu1cd9Qorvt/Ouw/eJ4boOIv5M+jLOrOfIHC0dM7t
YMmyxNw53+yAGoZEh0xHzNqPO8zBjslHlibKVVaxwHhVejvbLLcst9P0lO0RJR51
GLPpLuDYvth+zoYLpfCF6/u7XLWiORtHoGj1JtRbOmtYcLOzLpvhORNipJRzzBdY
MJqXLIm7Z0ihQlSFxB7yR8lLYAWrU1DCP/ZT90atWdbzwhzJraI1w9eyqIYNKZBr
ZyMd4TGN04CYf79C5rbH9EPxaMo69RDl+Q8Rhfhcy+UZbNtRGffOvKCB+L63u0n+
09EVFr3qcLdLNi4JfBmrrEqyLyJp+3aHtoK9Xo8OHV2PwojkwAG1h530q/OsrMYw
uUKIxvPpTsIumqiFOUTs2rPFOlguxi8uF4Tye+lW5Nw7Nds+OukCHr/OOjnCJXkZ
CtC+VynzUGOzETvnD+IPOmDFjg0okKnspgCu7CXJC57tHFWg00GK4ZAKsOX9KQPf
2LoIYHpbOtoWwGWxQA7gFC3904Y6KpZMO6w9Dj63xu+Slo9ao1tk7g5XTnUQw9/h
eihnoaLNTXS02mSx4gX8/DXmRh7a6fx+BZGIo9Pd1ms1oi4JaTkz+Ar7dbzNQPhN
QmEIM9TcC1+5TPHOh5Xrlm4/Z2N7Z//kpZj+BPcjbCB244hyDofLoi/ZdBx1mUM1
nE0KNlP8c9LyoqdScjArE1qLd3FtB7MQ4+ogCG/ZyD3fFhEkGjzL1US948aGjlTS
NlmnaRvft7UF/UQAFYMrbczIhlwutOnDQFjMb1v0qF80gbGY+Bnd3x/LgX2dQu6B
UNlBcfyhtxphizEhBUzKbn64EMOGOaOeym5knfnxig4nKknanvXSPByZEOGyBeuh
EybogiK+UoqCHIJ75TD4ArTxPZg1D4kjjjpo3E6wblC1/K5BHvu+WQZ3t7iZI0h5
he2HvdaEhzUIGycygBAiofkVBK2wy8xQQfiU4ovO+0KCBD9DF9eFzZk+oAJJouQT
xaYcRABgGa5bKkSZ/beDFYL9Wv5Z+I47zY01P43Srk11d12ZcSiFWot9FTBRgGxz
L90o6o+KAziVqu8Fwiwn1HKVtxzbsXJvqxrSRhwqNuXw+lvyvNvLjGJpwBQMr8Cq
YqnL1Cg3Vw7OKU33xsHcOP4/regnbX1BloDHTZc1WMkGwSR+ctnozvjK6KHzkAkU
JJ9F5Cp5haVZHM/qw2NtHVefI1mJZQTtgqv4sPmhvDiVZns4lp7GIKiEgoAt0GN7
4tAF+MPbTwh1526dF/W41lzq1UR4kYUzfNxGgYcidNHAb+tJRTnERadIhcT67gqb
v62acpexZvtkZyMBl8PQIy8Oz3s2ORIcJwr9PQg5CqAQ/lDAK0dGb3LzfC2TBRMe
WfjFrSScTngG3gQVggLuTFlLLaqZhfbi8Uq9PBD+8aGkEvurhA8O2CDo75H5i0zE
dbrQlMZ56yo9G4XxgUvE/6PaIh0hI0stWpIIsHUF8AH9CvAoceiPBVy6v9SsKREg
on3GluYo7bUtY7kEjQawiKL9asufBTDcFGPf+s3iV6pP6BG35XwKfA0L1qiFQrtW
MVfIfIbT07xRr0pWb1dteeOE08Rj7C6xaJR8ZB2VK0GmLFVoVRffMweUpFy84ylz
8h7Irl34JoUaUWg1AGmXsMmzBKHtpG8EhK+5JT1KbBSnrKw3906tEzPc4rjdMQVA
2OMv4WEI7z6HUijTrxV7W9jj0aboTip5TH6WRPnjj8y7w5nDetnydzuMubBBHFKy
fMSOMu3kbJDyOfCvwFNfEZxjnN3NDdpTJkEQdPvl9onNkLTxn4o5f71K+2lLrfxK
qYZGrvQtZwFEmO5oqtLYzJ+PuMKDKML8Xq9chXIUPc3Wo7wy/s5M13GV5AHg+FyJ
bEfUlWuhf00klLNjCNQ3O2fIsjKy/whBoiLVREc3qFxEYcvbWsQGie3MPGaY+l4U
G/mrwFY9OEKy/ExaMYJDepP/e3hSpuPqdEHZ2R8Wc9yF+hZnyGjtW3WqAN1/kVqn
Khs38kRqNeFo/JKpb+XN+2T2KuQ7884uBihQ6ZQ86XZRWYQp63Ctfuwcz99nv2Bv
N2x47TpOInPSU5tmghb+mE3JW9EOz3rD5wuzecKJ7FjadkvW26c5kxg1FBMSfkLb
XgvtI8/KKKuGeNgYG0iicoid2ewupOXlYb/ns/mPIeXadoehIhUuG5F06BHn7/9p
nkQ1YBaqvSFsJdPHT3Gx0habDy2uYfYt++HoXN/fIr7yp9rhwXZ9GZNTSkLuD7bh
4jDz25sLl8BqdutXbqlX+E95fq6g8AqoiRISusnZ1gf2fvVDnrOX9JDLfDt4kZVt
Pk4nHayQP8LMbEQ++AO71zjqCRFifiKDQUFiGaTe6H3uoev4RIavFaqjUWqCYOe4
gc+TLrbXtVVlxnwMimZcNeS73gE9+0KX8WBH1GjaAwKvWlrsi/36N7Zjd9OmIYVB
pDhl94IhmhsRRbi2E35s0cj8Vk0p9XYDLuI2jHNFtdHa4IPmNu0Of95Pp2Vei9wK
jMDYYJ6emHsw3d3rkCEppm5zzhrT5mPJQzOpjv5Ey+YOCEN/SlsNzgBPEEq2VzuL
mqIIZIAwzWNiCM+vi6HaU7tXbFcIkaFUTa/vEjF8SAu0uJLb1SkCjjB2+fSP2RTa
fuYB0+X0gCXxoin0nsghes3x0CCjy+vXxrEpPYhoGjS64ZXl2/nUxs9s+3ZNXzhu
nhA9W/V7gZWcNwNG4W99nqnpvZx1uaGqSLnwHwAzkuEwztElQsONLeL36WGq+9MK
sPNPL+EvjgMwj0X+k1Ruzx9glu5M8yCVhxju752be7NCgSz/9veCAvSQ7swFVq0x
Kwe95AQG1M6zXoBWMZfqp9PkEEt0L7zKAs4BiLC1jL5NqsO5aplUxna52MjtrC4M
6UY3iIR4FDPjlj80UNkYQGuCMtoO/lzyQvtJ6CHXAj8NSzM1iMMMjIHmY4dupuXu
Lc/5DyNP+nxU7IKG1fmTyeXY+FUhEqT/2pQ7+7u2kgwod2iU875NhLcpFgiApFbi
mSLEYpv0iX4sgDTigSAtukTc3PTdQnnZHLgA/Y+7B9cQBP992eIMG7eGhZJlLxnr
iGVKTaVeMUVpmUeN6Qehd6Y4gNG1EO/+F0AuBpfuyfvQLsZlkpngnjOl1lyNNDKC
7nPzQYxefPAItge28/HS8/CsKTYBhcd5EX4iwC1ssBKggzgch13TEgZykErIaJir
8c/ungcxftOk32e4yvd+7963/whclEL1qeiW2/eRbDjCdkYfd2qTZ7v1eL8jC5Yk
d9hVKZRcZecgEO6V71SjexUSMeWEdjL+dnKdBr4lvih43Du/+4Km0wPDuecj302U
NrKESDxpRsWB670rcAVVnh3vywIZFSx1W/NBKVPr6hdMuQe9K2cBxJxc+qYdJIod
TPvQImM/MEn7tl0a21VQKlRJh3KcpvobvojbhtamGNf8Zfgst+Zo+NMFVp4dyt1v
dCHlW9sM59a/tT08eGWU86ICBngrIUVgnx2nq4DmiE+Y6U2FunAJO1Mk3v0d0U2C
sLkxr0H6wnPW6K/691/C7VXNEAsAbD+t43G9KSfuttlivBAj9zqZrav0kSwQmQM1
f53NKYIEjEdgTqFdKNTzLW/BNiMlT5PBpU1RFMzmfLn3h1s2TsDvmDIfMwy6Oi5C
q++fZqOsdhV/2aZL/WFc/iBq/MZdjA6SPuAAdBXhHdtjqV0B160aE84G06tCZ7UF
0BUiMdBlwaMu0jKfFnUyCWc5bjfQxqaFA4u0Za6wmswz0wQ0+l6pqj8XjMyjtiVG
ZYJz20BX+it6A+BTW9qyyaWr3vBLSOKTUBGBSt0T5WEN26rMvNMqoUZyeW80ktCS
9hC7Jm9zr2gnEz3LO5AZQnDQcB/b/DU4LbmUmjls8LxCEKSYsGgvJXDVgwiEsqQR
bqWwvPhVoYSSQ2fn9RKff4MQBHBv6ABDjlsqbQwpaCI+OfKb36ChRCI8XPWd8urQ
QzZV2JgnXlOEPXsBGAg8AYgcUNGFbguShq5Z8A3qE+m9Oy5u9PvT7ZWD8trISuZn
rPknTrg1o5GwQEAh4Vg4VYQ+xIMdup0rhrGP0He+jx85+23mDs7h5EsOxhjXHa5p
f+cdEq8Hv39T+diCX7W80hGOcOI15rTeLyAJiYM6DZKgX9U2e/cyUVivi+jk+whh
KHaAE9W5XGF5sFk9Szk6LeJOGg0CJFgVLg92eo5ewpXH4WznmFWG7Mn3LuenyIYa
f5t7WYX2YHTG03T+NeF3e8zAJGHtOjEfT4fIpYkwMK0j8rJ3e1VkNxLC+Tfjg0z0
avmJYP1BODIqRkn5IeJg6rNqAbLwSgXDzE209myPtsVrsHQvunFpne89zkBk0w0W
24c6p5ePwLizFGBJVH1zrZ095i3BS7jI+iT3+1zfwqVCK/83djr/Q6K1TX/PD1A8
TGssNDyRwe7dPazR6+6OQtf5Iu2o+pS5QxqcPbKEpoWet7q55hCidFXGOLaPy8XW
bZ99zkPOF4wb0WMKXAGIngjcLfm5Ltf4DKfuwYCCU6TS0rP0E3flfJtVoSKtxxMu
NCUL0P/knm0W2kqHLkfB4lzumJ799J1PNWxPkgSGXbcRYeqwuB8WLToAQP7E8GCF
ZCT9aO+6vmNtXy9Ss3rRXpcEdT8pnI/bxfnRAWbve6Oms1LwVAw9wkaZ9E3NK/TE
jgOPuyhnF0BIBnplfBdi4sMKIlgnjJ1IXKv+ZqVCE3Zy4Vo1lRF/E9x5J73wIf2R
V39CCrlijF9goet3C4fCDyTDPdxH0/iJdkGy9fLLs2ybk2EZ1eU+O9XCqiIIC/OD
a2pjiQmpxq4RXwoIRNCY/7RTtrYJs4k6lUQbBhv7zaHvk+BoKXh1U+Rni41Owxgv
Z9y9QL34ItNHRmyIyWjftLVvfP9UR3eU5pFEItlAqc5Hyql34l+TYpGlA6sZcq6J
XWGC+CCiuZRJbnBJyhB6wKjTvXapxYwQkv1dADOidxLeFvHEhcyo5G16HDC0lLRq
xZ1PMAWmi5qc7cHjih1WgbYP2fvkTdvcj62dlfr++FsXTfSoQ4Klwhy0HY2gjYXC
kjEQU45fuiL/bhOhF+lcSrCcnYy7cvJKG5+KpielMcbGugLgu3/578bwjJybzTQX
c+pR8s5j4LvB7qGk7SDhaiwernX1kVaqa0+i59tscKzwYzwTV3KmQ7WMv1xWNUYA
mp9pWOZvrdDEBHP8njR1heI0vn4jeForkK8keK0ByY6NSz2frlfFvz0Jse/L+4hX
JJWu34QgKlsS1dn3dWwcs/suELoFFpB+UmUYZ4E4Bm5Z9R7hD2rHEpUG2Jpjutrk
bf5CaHIIzseobOs0/XB/T+Lcz0q6RbiVHjFlWc2mqIiRv6wUNvwfNQMvLuZMIMoJ
IMFaVm3by+V8vBooYMNrThom3K6y6jFtAqBRkviq7NKKWWOnqdGrJeQgQ4GaEuxc
/9eT6+v4Csalg8xMQDdr5iAWDSx0kUqpm1lefG/Zpq30LG0XQZ0SQur52McEPG4M
VBe9YcTiMwZUVQevYpamBq/Z9KYGSZG0mGPMVSh13yotR9tZHP+r3UVhm21xnfce
8tjegSfZOv1/cic0ei6buptTX5s4oev/yNbGAS1djEUkKI12QzD8kkqlY84KTTcG
mtLm5fhU396X7Mtdax8PnAx+86GAMHO6zRlnfGg341CRWDeiq4xdaul+/IPrRbnt
v6oiUNDpqrl9qBO5j/+//YF1D8KbAhZJzFB+FMerZXt7oUruQ7/KN+rawNJpDD00
E5IP+DeOYMG1kvxHVDjjookCgFpRIvyKZJDilWlEkn8MLH+JDrCwZtv4mMNfBjun
OJ6h2Gabe65RvnyliJyfYvjpW9m36QPBWmGdq5sPfHKQxBAAYIqpP8e/INNYbAK9
PE5hqgSUg0jrVlQx4F2pqzh01fqfQiOtq/xcJDBRw82skFPVA6oHoLmTOxwq/d4L
Sx4D8kcZC5uWeFkznDtl3Vn915gJk02ErKzorP7dBY9Bhd9pWy2dDEkS2A4qSq+B
ukyLJ3xy7/3JmwccqxAN3+z9GYhp3o8Ky56Lbf/87Ia2QCTVUixZlseHUP54Rtb2
BH4RNeEnS/FAsG+VtQorImBWlt0zFX58wYkvDSMm1McWv6bAasdiqsTQFt7KR6l/
D8UgyaLNzI+zQgpn0fpAJZfnec5Cd+L6ls/1CJgy3G6SAZcoI4Nw3e/1EVP3Bzh9
HYJl/tCB1lPXio/GdR1/pPHPxlVlhpfVmnMDnjnqJi8OCxblTjqtHcVTZruLct4S
GLhY6vbjoj3Sa3xjdNJTaNpi+bU7RssvHJpvpilNXNxtlnqxowMDORh5IK/EUA/X
eg+VC9L6H4dyz/wfuD6l+fulfVbQV7lt8f5SNUiaq+fOgibnSxqe49no+r/hDQmG
NXIU/JdblVfBnINTHUBn9hiKH2wBJy4zolcmKrtEK/Ka+llFBvhPEDsa3Tgxu4oK
VkJ4VrgsBimaSj02yhbDjdBcL85MaAd9BvtyYQ5gBWOvByfJE4d5wTbEB5wwOZQs
K7Okq/B2S35+hKLY0zf/tbYlcUsUmGOln38qz4FnU5oej+4Z/dWGWegSNWHTaBFf
h6RdQ7Qlzh0KpFenfXeRWFGThFrwTrSJrK+EsZRyBVCBEf6BXhmUbZ8I3lCWMUJY
0U8gbM/B4+iaPzZX7fLnfubjmfGyNbh+xeqxTt/cbk8YQjJBcy5BfcPcfsxRoaHc
n9wG9WsIVyNsxO+L99eFoGNWLN6bQUMA8l1IBSX3NXKcxUIUw71tkJ09c3en45GU
wztVxIju/iEn1AdRg5987S5ThU36IZknGmTDzhz8G0bLjTOJxGqO9LOzADDOqStU
bBU+X8bmCL73FribOiFfa85L+EPm9PrPmTYUp/jB7qz0Uazs2mUKTbsJ+WgnWvOq
HzGLNev9CEV+0q40xDNckvnvDmTzKe1WYgu+SU7p5sJt5V84XFq22EchnWTrXIfd
ASVz+TbsJgKSDwKaaMf6/gqqh/TRRrO97SSsL/lj0Ji/UxgizAqsCZ3y9/tCAR7l
/pTRh03T9bjv8vfHHTEYHFjXlSurAaxJNFZ1mits20GhBqHPLwmhqAVQil00E1em
2EHBK7ld5ziQ1YKo6Wgds61OZPZMamJjDtjUHA+M/OBFL+49Y1kYzDYSqtdM56JC
ioC+XCNtbm+Y9qYOF0L/vNX9zaIX3el5SorSd1fnhg9OKAm2j9qlHNXDKmBl6AUT
v4VOtf+yeher9v/4ZJ/5EhFHljjeJixMkIiPY7MjQBC7d4wm3byg3OPcCsbHRqLs
27R528brOAsm1u1M/Qvw9GJNOaVd3hlDhzcn1OrphkUYsYIpzXssF23FGg2LcIO2
GzOX3bgXJ0cV+USJvie75Y0p7aQFL3UiQE6IH3CcaryQc71mI6vfapPZK70Hnznl
W/xlSe3w4q9Gqgwsi9AAnh9szr06v7Lcp9ViiZ9mourv/5/YwrBQYTdq7TgRC/xy
6aYfc5AINNGqSHJDUpuVUQk8n8dm4bGoMRbmenghFtEC17ub6Ld0revgSxT4zA4A
yDIioEpndugxFqzwLPAQQ9HABVWQSktd6XHnA37Qe8BTBnCVa4Wxx0aostD0RJ2k
2Haa2w34bFP4+IKfIRsKqAFZXUogWfLzmiiZvrtevLeVLD0TQkF3fjmZKJ0NhRXf
mo29/oJTR5F7EzvbHUWn9K7hijuvF1Bu13OMddm9Dy2qwqNAN4RbQJxsspcvnGXh
pl9c0dbX8VhHEZmGUU38g7xScFemvxkxOFcy6jA+cGEmZHfQMuFbXyuOdLmwzuGs
zh9qb+8aLzaQQAppMiNT3GgbWWoR6SJVqKTcxShycKGeAa0dZTPHm+CXEGo1bOOI
YDSzdHFVmtkRQxytskU5Zg1JHs6ndPeosvNbLhcArM64EMjSfjmk8T4zTfHQtYqB
OSmJ2IXBxHumlD8ppl4E9vAgbx+w9d3v+Ae4Nht5a631ja3UVea75MpoYXdfhrmk
1o89Xm1lJ4PNUATC5MQ7aYqlNyR6O/eEUNXrQyYxIwFVYpDogem3a0FJ/7cdJO5D
TQl2N0Yy5XcgtiYTNka+q5/ZvqSRHPKaenL9MVXB9P0NHabcOJP+3/XxvjsbuXFp
nGILyygDKLsg3JCwGT/mIgrgliz8lou2DqGSUscZhiWHVPBIO3UF82Pf3/6oUqWs
J5zHbnyrPi7FsLYn0FHcB/9jDRa3QwtCloC4Cw7mi+l4nDQ+w9o1cDXHHr8XwzOI
9E5pojpHl1WEqg6SOC8Puq0qDRr24lE1EluxusKV0XMGNRzDRQpTtHDhcxP4KmgU
+4iKG/Giy3hBqLDmHSDX4OdVqoTk6amLkpA/9Fdcn5n8luJ/dRYcNLpnfZqQPANp
b9b8y4IGtYXCAi17S61gm/slWEryfaXo7H/1cRVm01BDebDo8voEa/SsgLnUS4vt
zHX+nUSmQWeCLNsWF7vp0mCRA+pTyUnq6wkxfHZ7Q6k2J3dRfwXrUuTxilob+lum
itFAgLhxXBaGa/7dmpxVGtUvop0F+WdMS85vI2efxnlMGDH/E1bVk75Zx4Cf+vE0
AGm89ur2PVviqICv3EA8/hT35+9Z7dtUn4ls/DdttdfpkSvg+4JVcwKOxc/NIxjm
KFKXRx2vFFN8fWfWY5nk7g/45PRN7e5y2e+wDImigG6riLhRhrNLD4lyh/g6Nxqi
8T9QjkrSasSAdvRywt8ymt6wEAHi8y1quluzpEPJi9I9lI8z0OXpO5mpDfpUUBB3
/lCk5IsD7n6TdNiLNTL8+ZCGqWDPbrFHummx1PrPGxOUhBMJtF4LhvAFO0xR8IMB
LpEqDIU14uMFqNrRjI0lESLBZdcP/jj9cD8pgOsivVHohAonhN0XCxbuh+OKehhX
wi+D8I4DAzI7lbuDASjIbt95Y/ZW0aR+cGewloZ/mM2tRUdD7Z4g+FIdE09CPgea
CXmMqehzhvwPp4NVlqRIM1Qd8+KmMUhVNaDc2JPFnBYU+BH75h7ClqlDjVr/nNtG
YJQ4vSQ8bF627xr6uWsG/dkkzINGFrQ1EP1Wou0213PfWgrKaDxPQAbf1pnEDgbU
7AdPalxPx9saB/v5g+trE+q164sEmlt6vlsS/NNJxBZbWl7DSF2JTOv77FsdWBAD
1lfSKLmorzt9sgUX5rGpLMrJvrsuubpCMUn0es9I+spk7sycI68LnS9HDAloqlGf
B2jQD2r+ZDrtkefZhKKsylmXK+1PfzIt48TznaFzhdRd0fh/SaLRuQA61SiTHmlD
gZ77ARgQxyi8k923ej7zYo099XjenRf0nWPnRF+VDejFHrURo1L0igdek/YBadvd
u4BSQlzMTLcyYITW1cWKhxg2+hEXGfpxX81wlfUI/+EgoTXkVXWavi7u+1OUcC7x
TddPswnD/kYRWcWPlwXz09QIwop/eM7tloKU4X8spAEHGro9i1fEL5RnJYdpKFP9
7FvNnYT3UMKIgoCPL47Uo40H9mGrJi1kCrcEMjY/B36eMzJpxv3PkScitN6Lqz5V
BTXaYzBrjBg+DLXSJ4ko0cblhRXOv2eHAXLovBphTs9pANZH07m3VUmzHsUra5E0
XrMkRt/ZltN6F+z0nt9pQWg5MJLlwbZCiM6oYujMi/auu6e8185/VA+gu2+8Na8r
XsIZKEzi0fzkzZrMecEK7iqZbKpBywPHOQmVQAlzurDKtBJTqRU6P/+tyQCOuX8P
TwvoGi+YOgmIMLtzUfpGOpHzXXxjAmNDxUpZV4GAcvRtnk0WXIbOJqpJQUxyp+RE
7vFL7itqczLl+4lieDpa58pS782hBRGDNdird9v8w6LfBYYpi6wG1DX0oYTQF5EF
xOos2pV/JU4NxOqlI/I3XdT9MqzyS6lyEIUGJN8GM1wTc134pWOFhwwSOlmp4NBx
yf6UZs8r8NjVOMcQZRdEXuiCPTmuTpxJz2avKXHjluILX5zdvC50lUXBh0TsR31V
jrOTcIEmBhXEJ3MP2pOIRhH95sWgy2klPvc6Jt2NgLvOS/++BaZwGkrzpicqVAJM
OOMn+sTbvlk8iHOZ1PC3UkkoqQb3tqUAMImeoplnicyzSfpKfknpLRzBY5y4J4vi
G3AqJ+N//Wv4Pe4HEAeS93ZV+oXYqrXj1VTWN2pPiKH2jupR54Ck9E8W+vOHh53M
1lbDbfjtt5rlKPx+5iB0+YjyzEIzEnopI01NCpGatXmZZ/nFluyVMTEE1c2+5jGY
5HpPdNzF/G3JUIJaF8XEdLsjC7hpSQeOAnv5Mv8MLMOFaxk0M/c+AxI0zRXSwhD6
txhcrv3/4sTAOaE5z7cm9vrSNtBKaMTf5f6viUEYcTY5hitM91QVszQX+dejdfws
sTLUPmiDjU+1ynP9b2ulwpUTTdf36Xh8nwTAvJbTVgsc7FqCeyshKz4Gb62VGwyX
6KMd42T9XxTVn6cxDq6nMug0FUWHGAVyzL7wJ7+UdoXwqTjWXPNRfeLdwrwHqWMf
RJ+jlrzuQwpTyvzM7ro9SXbXjvdxQW/4Im034JlkUh+tdCBXJWAJDarrSRNijzN/
vscEib2hKIb2PetGZ/L7j+4COYDBbtrOzBAKOXduzDntvnmhL4E0BvdYhbOaq/SN
RP4w7U3xXRwwVd4h494sd9wyt7CEbMk63mEU877TDjymRxBLQdbLsSgCmKigHxNf
xcX7dBqejWVaPo6HT3TgGwP127dFq2RLzbAEMj8oocaiAJSNu7bMBQk48svdcSAo
QGacORBUVlzLklT1faEg83/TJk2wrNy3VucF5F7fmxzmHHgXy0q1ZA+edVGFv8Jy
eLF4NqhDxLPahVuXjlN2j+5x3nWhhj+5JLa7RPInQqZViJmokYgWX9BbQIKTnYNf
ysbdydPVKRA1eOxkUtM+JXVZnSG5aI+SiaqhDAEprb4niCJn50rBmpBSQuuQe+KU
csqkn+2AtjEI6UNr53KOOI2F8c1zIcCuAn1jEaWnw8ye5RqMcEqQg834eu86xL15
TyXZFieGvn51MPRoTM0/RHu7qS4b4CtUn7LlVI+DB88R3AcmETIepRGdmcfkLbdW
RieYV80b1OwRgHmu02zyHA0HOqLXvN8DBoMjCRETdbMjajGkcSuwIkdBnyUu3fdm
6SMPgHx2kL6uAT4/xz9WWFBqnIqfsuIukalCaYEu0z7Qfsdl66WCxPIepWbMlCy8
mvGZ/is1YP/1TXxpXHGdOfAXiV5re0jZlSMoPI9fDaeYu7NyeMermse/dJeNLN/O
c2QU7Qt8yvj4NBO3B0ZfIKrbfPigXozgVdd5orvVkcbTKvjGy3wtgfAsxxZjT3fW
l/xbz4zeGo3c1TbdOfNKSgNZMQ+49p2/GEkrdK2K2pk0K34M4zMWlP5oSQRFJaIV
RJY2xnVv6B3U51vOVNrQENmzkvFeD3bZQ8es1TcXf9/NCp/8tI5kLpjDSAspDIwE
TDmmYvMoPQFo3siCJbtyXhh8ADaMLB+kxRbvSfMIv4mkXlcppRcJXqzrzBYrYmGn
LRBV6rWRP5oXWnN7uSoCyf/VBhTa3lxRWM/OeXNkbO0C5fvu90cimI6v9t4+p2Df
1d6KPuHAo+fPrlG1PgTvD4fETPeAxVffKUx33s0luZj2uE3/y7K/NBNvpXBYvpWc
kbm2xzKVIICGmhkFF15mMMu+kro8F/90yCcOMIhrhkT41KTr3ar2lEO9XS0wC698
cOk5iOx6uTT7ZXG2wQg/f5X4vwXFqbFugy4CYAM7Z3/wM2aiWBwJbNp+BsSW3hvS
VC0IEVBxwIItM/OUQSCHf9rlNR10mcJBO3bNCbb7AbL2hIHADsJYcnSI8cXtfnWe
wExn0QFbBm+Q+00Lfh74Dj711XcqFivaFMw7ONm5zeSKEVZ4IqL3mdAojtRCIAPm
XcB0wzfHtNZSOmHm1hOxH56Sp6iNizM/Km6YS+Q893frrmNDz+7Rf3X7LP44Zlvi
DPA8COGNWgpBP+DVDQfJgpBMjjYTiJcAO8AFBge7rLNZ8mAEOT7DDDkDD6kKJtfo
FV6lYFkkyy9UZkruFiig1dJKxMnx1og3RF0ElScRQK5wB0xD3eP10FJYKB5Liyj7
RKgtKqIgK9FiRWCVdpNzeLaNvw3UkSb+Lf4t6rpjpYXhSYD1R3bJklsK7H3PeUEh
ymNSqXHc3SDi8il9Z4347yBLSf6Gilwco6z8kJf3Xcd7r3yL+BYA2QBdm1rABrGo
yLvMxoevaIpGkNf+tCzrrasubppnbxzsyVeTvEaCo0TzNCZNluNNZLHqVxfeqKUB
LH/5jOyswLaskOOiAJDEcoXwMDtH/wdh9+Pa8CEDm+W3+I0g28JJQwN0bYTbxVSH
AD9feh9wbKltZPnSTmWbFmNlM49VSJIFmra9r5DXYy6jXMWTHwZLkuzRHej0S37V
EqmhEeJC/DUHBcZBlSSXxs1YQutpNtTcEh7tqav83ckaOD3JtTTgoya+ypI2Jd7k
XEse901pDmu/FdjV9RXoUz6MlDBT/2AttqZTYj1FSqBPqFr9iCLFLH+s+64B3gRi
DCo3gSpDlbS62ESNxGvYZExJXo86A1bd3Fw0Cw1lq2hJ6gCZW6X91YKHl7Zu87fQ
AqvPKdUqhS4cFvwj6h9oFijJbYfV7hnKuT4Q8D6BX3nHC9gN9u4d2/xtZlEpf75R
A5OSWY3TUuGxXeOgu6MVIAt7s9Mj/nqqz3BEcP0BzrVfWDlLiaAfWUdODqX/yG2q
EwglOkHpqqZReiWivSQsRfuOsoSiQ+JLJVfG/gcK6nQ79qaK65dFFX1uzZHcl4p5
v3xoKoSUJgIRHhHxqajXmzAYLXPTcaJM+wk3pGakUsTZz8O1pmNkRF5wnArfaJBy
4ZhMXV9HkebGxrdtQN+bqoossTUl6MDaqIHtMuMwlRSTK7dMk3e4RKy/NUpoAFIU
yhDw46Fr7uEEMf5Roqh42h/8mklRjAlcs+JUkijnAEjYIqyrRjWqMWKuolTSoIpX
0X72lahhAeqybBqDEVJLB+v9NCiwIsN1FB4zCm/iKm1RteDXgK/P12eVarIfrDD5
JXE6qCsng/o6y/+5nxNlewizy3MvIjkwPyWTiYf9e42taavgINZkxJcXUrbEys/R
XfL9PZdpLIWS73Rwz2p4LH2T0MgA+3zxXuO0UaXpa8ScGCOZPJbT+Em9OtLdNPXB
Wd1REhvFqjez2LmdcYSJr+07SBhN9uo4Jfj7Tb9IIyrsW+eUytLhETV8Xq6z6P9F
23Slwx20aCu7tqiWPMjXBQiQZvLCd/YVBc/7mnnTB3UGS/qDRLvfh0Zt3+IQK8Oq
+w85yIbNUyHKxPH2eiAWTuusvj3gG1kK6pfE26NYK6ASAZ9OhcGhL4HyrHTwrBWR
vbZKhObEDGOWL9iR10fpFgN/MSrxchVdHpYlDUzVpCXBUFSbPhC2sMirfDiNdXRg
LYh1AyQ0HnzyFd2NuWcDYtR6XCkjwFFoEzEWk2zs6Fsj3+Bbe9wDuFcGbba5BJEW
CN2uCmAFxGXS3cd2P5N+oCsuAgaC6yxnHeTj9Qcb40115PTXVVpdKh2jN1l4Ftep
499kVRaPHtUqDeOIFiF6meQdb8mCNamVzGTrpDcDYeD6udoKK0NYSViGDEa664/H
b30lreiMMaWhhXJ1fkxCofIO4wr3AGOhpHYpStWn9NmtOJxK2fMCiRvFMbmdEYKv
Ranb2X1yYv1xb31rDjqbyDZU+KeaeqD3M+nT82HLRM/LEWop1JqAPh0lqcNe2+GN
FfvK+UieaM13Fd3Pd8Trki9oCeYD5sRBNDpzZo9x7uROEsXd0GZA6PRtROJ/4UOZ
sqQmCGqEDOtcZr2rmnlcmLGURXl1cTNdAvNe/fSZLfLWojXOxiVfr2UgcrAo2z6H
fj7qNGXYK4U+7kaQJ0zyH2uINGem6uJ94IcQH4kFu7SWc0s7vvU6cTL7fWM7bwc4
zaAXdNirh9v2RdnGIX3FcIEGZ3mvO1sh9tgyPAs8/hEp13cL4+4n7n5VyRq52Rw3
UNeOEI2yHP11ikKaDgq4vxDH/O5JJg6ZRUIss9UMtwRugcikNAMU3oP6KnE4Zp1o
u0JiZGjS6ur9sUdys8441Elj77+FowSxBQUd81iCxMKAPZoxT9O+l2vYUhRHbBqZ
3EzQmZQqcmfWeENqCrnSzbg+DGvG2TH2ilF6hYygcKZIbGOfKqHaL3oxd4gt7Mq1
enoX+Vrax9Gv1Jy688scmsu1+e08PfIo0Rlij8+uffVQhQe6zSQkTVMq7lB4NpU3
VTbzyzGSiG99jvvU5E+6M27565upUetTW3VwQ6esz0QBNzeQj4yElAdgnpY+q8HG
xLGy64MjqCdlUN75aIKcX44scce2IK2qbeGbViWXCzVxnK+w+dVNBnQUmw7+RiNy
IXnGz7r0oMgTpK9436zybdT+ZhmcsdxmgfgcIeIaPCPYe+v2U47+aRW2m0gVsV0B
iATSpd8Y7NaqkfqfhSfR/4rWAIUn5an8XhL+70cFF0m3Tp9UeheA91XQLl8WrDCO
Ku6VSGgt7RRzhU8qPEpj3NufGAJwK8tMZsDAJzPPDAyUFkSD4aY6kPpKryUz9zES
fOujZER5R0VC9fpYqkPReDanjn/buA5nPgYGLX1vpR3deXmqQgb7/3P2wc40vWbl
pOVxmYkHP6L1HpekIEETtTZFHhDCHfI2Syx+v+BViXqRn0FnU1fB13cHmYcPUYX4
x+5iP81vyTPLE+cZ2MBXUWzVg1GgqM7rO0pAmXXt28wlAaZpcFa9CcEx04KmlIYm
VYEBfu2nT56tMX9JotenGR+QnhOvgqe3IyVrmv5ChouBOj+IewgM588tlVwJxyA4
HNsvb1+lGotvODCISzdirYfgLrrM7eajRhyWqmMkPTNmpmBAy9YBdmod4PwHIU9t
xwnbAdktnE7tCmcU4t5gkTZqt9fyh6gU8rqQcHvZeyLlzlWrE16jnjJKIlhenZDV
SsajNu5jthDfGEd91tLaC7SL5xDBrQGE1csTOGet8aeHP9NdrU70YaoBI+YGTJ/h
LqS+TGt833eUs+C+W/sHSE5qMkzHja98k7NwJ82WgLOXr/6ZtjLdQ6StMlf0CY9f
WMfLN4GcjLekSHcwHAEz1Dd5+8/LAqJ0bHjbsuEF+c+oq9BLoT0h9qRAzRRm0XDk
8xCxSYHdjX4iMi6KduCB5buZ7sEvyQpPeDIQPtA1aDSILRn6eJVBV0wcYvtOds+z
++9Lml3AVvV5c1YoR2V+qxlLj7hJm94bOfGMXQwqKEfdrVvHJSLhIhFMDw4tRRMN
ymetcVYWsiwuTD5hrXgK5W0guu56Ye/l1d1k+zCp0EOKq2cy9xPOK70VrFQOURhq
8sindyLi7uYQll7qXLJfZd8mWWyht2Ww08+nJ00bdNdJnHvZJBO8/eE6+6WFX0g0
3KTzmoAP5uOUw4zOsrKVzv0NxQs6pp0JW6RtJMGwPonDJy6ivx9oC34ubq8GkF4/
rRswhX7QQuhhHqS1mfcJerNVuGbz8i/2uliIgVQHcXX6ctfVC/JrCoi/JyIsWOQN
L1fP8jj+/nlJSCt14jVCu78s3JnFrkfKPpTlPZbcHCxpEmsvzrS7PypNagGzaFEw
gtoKNyVTzo5vh5+l+yrRihJ/T1wlZ/hZm2MOdLMAeXTyp2cwGuZ0GQCkB5bNcmrB
tQOe9fxJtbjCtd/toL9doc7NxAK9nwb3pFLXR9lNI/N15FCV5MpZ2/QXP2IwMA3m
CracFyyEZCbNH0qqFEezOb8kigQhmAtMY+wlCcXixpw+EpsNoe4fs5lZZpaTGUJT
yw6nubrMnXq376Y/0oY8m+BZS1Fe0vhRFTrpgEh33QVCbPeI73zNZuaUbt4zNqSF
fj55rRW1LlGZRsI6i+YyucYyxNlHj/aGFYbhG4ECEGpRCU6PwEfDWROId/O6Gp7l
c44xghIXS53d9j3naeICzmJgmwZccMIXWps4UnZ7Pk/69UiGaN8VzT+7t4ymf9uS
Fo0hU6sVr4v8hw9cbVzhdcLzHnp8RLfdix0un9FBz+XwvEln9VXUXIXn01PV3uvr
JPVnGMFp+ZgkcRUSyJi1sQuYipq0NYuj+3Ls0K/mREqSxs/P8H/SMFM1W3yR6M/F
T8fYAIhpWMXXIoJtLf8e1HalZRnBH/EWsMiFkNnkKU0aAZsUZDD4AWY+yZw64dsI
waXasgI2MnWKwPCUeVMomUmxwCtq+4gbRTrbuHqvS8x/dDW78yuHTgtowIBUQKbO
GButzz4vBifbWKGXK4QGNRpdHHsgLeeUc7wlGQgrH7Bt4OWZ8YZi7+geJb1yKewS
Y2Wr9naeks7uIm27+uRGnXu5w7D/VuBYW0ab/evPfwgQ+1N2GZb1wMBEy1Got/Ls
oPfB36FQrxTyiWTixLukZh94K4XdBrWfpepgGflDojD9AJU8dJnjvesyjaHuIKBG
SFv1uHO0Zdd6rTZXhtDR0ju3B/h/a4NbfhibP6CnbYVloBeWd92fYg9VavuDL64Y
/6lI3sZFotW21AG0JOamxE46t8rCd6OqK5PJoVA4TktfgkvJD0hEIf7KyRxHs903
rwG9eHMxo/7AWTt7P34TQBGwcxK3aYWCWeqzfl4MBgFLSty+OAfcfUaCU2c4wM//
h5KZ4c4VE9047sONxcTlNeHZWPdqQ7H3aypz6JL/p2Zu+79uL9EO6Mkb5HcPAJIH
lQ8ieZ+kxwnavtkpY7lwY/WaOB4kTqgAtn74K6cm7XRMawhEPhazt00IEx6RJt/v
OFLFFHq7UqHQfL/Q4gMOTuMCcgtSHTdvzaXkO6lKxNBqHkD6F/z8WBIPl4wo80YJ
R/kLiuoT/gghrFoG591dnifonzdW3T1lbvNbYyPfgVIMvzXADv0t5vpbEpagL60+
LtycSSiVk2HY/qPXqCJc9OBMTtDK3fGMeT/tPRfTYw4bU8oXcTmoVddiefh/GuJW
/kOHnBufcOvQ83MuKZZwfNQs5Zw7cPN8TQCAz8I9sPnDVN70AbScm6+IprR+haj8
43hPKgVMOJ672MZG7SdmhnMCw3o3mJY20YNU6p7JTmH/lG6O6ks9ynEITtME09EG
VhOg0+8x3vxBGxNuQ2JUsXF1EJ1wrajoqexUrHISE61jUxCTUu0Cokc2OuA+LoLt
aGIWm+d2AS1pCKot1DGDcjW9ohnG30uXMyP2tdZpdocs+d16txCdlKLsCREbmvUy
UI9CRXy1DwBLpExVo6EWXznL4NlrwxlkTS1m+0hiWtzQ+nEtBqHB/SW3/Jcqu7rV
znmnsfPCPKQZsw/+zq1gQpOxB1g3DkqQxFAtUGgAZGqobQ86QOY3hMnnBInlRGOI
ZsYOMoLlYDO8iDbuU4URL9R35ZMepS7otqVNPQZ/EhyaGZjSMQPoTWaA5isKDKDR
nKdSippZX9ZqehziAY/JJISCeHnLRhRND8abl+cmf65UJbUauYLt2c/rWMRjx85e
VbQEktzA8g5T0ZEWJdc3apbh0npPfpPtu7TCFMc6pZox57NJSX+unMd3Z0fw90V4
Gh01BojOkGiLhPMmuhwaCrRaXbFRH1gv8AHFI+NlVZFvd2Spfc3b5YP2fb3aCjaT
GRT5PB4UbYnVlBr+afRR55SXHqkggtMwzecQUlzwX5AnTBeZgDy6Z3FGAghxXlQi
ZSJzTDZ3a6NJ5j981AG5JXOZD25blruqmkCwTyUr874hVOtuWPbH/SbJcktdnx5w
Z3FirOK2L4slHTTmP/uKdtP0A8MU3t7wHTraNLsRugSPNQwXC+2tV7HbmyyQVJnW
BNVAKUajFHIad9mc3ACZhR5gGbVTZZltqSBP4i2RAU8D+EaUvwURB2KoBvxNlZpo
6d0609tGqTu3cFOOyWjNh93RZnqM1OZFS0erWPSeWEGAOnQI9QD4MgqzA5FUiLZg
ac66v6OvcoogAHJ2Q4MsOuqk6cPZRoBu4j2C55ELWGd/l6p5T7/APZqqJhCnNJSN
65xLwKE5b8maLv6sUvLRKSkMFYYM+HpKMh+xG8Ev+ctBOWXhDm6KfNNfWwuFJVWY
G7GfVnu+dKCwibFmaHiEBVbV3vA4d35+lNERpKUPSoAN+pWlU8wUmi2RF/YxXs+B
J/cGDUKACmk8tR3libEzuQgtSysciPvnmhZOngih/2GcCJqjRfd/ADzaBINcEcFR
Q2PKomE4G3e0UMdCyTtrHH/HDKuOBR1MszCiZL6CzQnefKg/ri1m5E2LHCmKvw45
BJHyV0lSGO5ufwzKxbMezcQ8cHpFWJyNjmJBvkzee8ZncDg08dOeUx3PDGiI1hdl
PNhkstFTlSOZIxGDvyRY13EeT0yPbqbiqHMlQEgXPllaJX8lGGfMm55xtkN04gVo
4PcarGIuHhtPkaAEyOM1rs1OIqC6pIuFUc8on7EFMdZgE/wmxjbGURIeDNJ4kNFY
0xOmTjBYY4MmsW33Tvp+v/d/s7QxKIr3f2ujVMAX1ruvkumeGS3JX+QZARY4Ie79
wxbUkHwC1uNC1xUSU4jGCN7L2HSqfPcvdmfxRiv2T428QocIM+OdaNuPngMoPXkk
Ubtf9IZTJWk05sWSLpU47JPsQy5wsN4ip8ypWDyQgRmc1w3FTip2I5nUA68b70Ip
Rtutnb/SLP06kOcRU8fN0Oyuwd3BsX3mAKO3GZ2aE9C4fgDPEhqit+6T8euw7fHP
VXPjIbWJs+wN+754t2HR/ZN9Vpr6JhDdGIS2UwunQUcDt+hWlSbxP4RL6SNJGEEw
AA0T2aDxwmUYYf43kVZ5JqVkonCdcVYGNQN69GgGnTc8OH3LoeYsK07vjgE5CIe9
KQgDJPk12ttI6dc27orY1xdYisp0JnQMerAD/nPyaYnLYCW6cQgGnhYVdWvSyy2G
hFA5upwOKS7QZe/lSR0zGURchjyFMW6Ubk7FDUglufI8ctrtom+c+fyzCFokzVkv
06aQScwHvIWVO9627yQF7xVYfMmG2cOEJgYjpMxORTEYR7SSNAQgPfFQUTexs1ft
lml7K4TCGi+D/ZBWggZY1GMS6e6BuLrkliaZZLxsrqjWrS9l8+vIigvu2JgbviC2
u/Djb05uaiBFm6RTQq+FdKX7gZumcR4J/Lom6irokbeRTviskQKrZwg+PV4DTs0f
iPBeL+N4UAAbXfuXnuBur7wEQrWrg328x7u839FtraE0pTBTwjSo9sbyPFxyNhqI
iV34nwuZsfkIg6fwsqxt0Ipqz1KuKTVl17H5JP1n3hoFNpieKJkEMvJ2aJUXryhj
4VcmwYRw4za6RVQa+nqfcA==
`protect end_protected