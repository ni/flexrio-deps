`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11488 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
EmxAgecO7UDIr+OXKjjkXFtjHeSATKWy9HzX+uXGJOcWWaHkTcrnCad1vxRvAjUp
TeP1EbamB/hlT5U10rDUsoBENZqDn8xt4Ijrc+mYLckqo4cPjqGt/7oqQPFuWr6K
uCmjil1MHsEytY4eZ57ASDG/jGekFqD3FZc7dKBrvNNpU0GcI1gQYGcZ7ddatcrX
TK4dymws12TxhoxCow68497JGrfC1q0K/FsEjhwBxYoeD82tz6cagyBYiqgcjgWu
+Rr4pONh3p+yCGRUcv3+RP61D4w20RBLpqHV3pUNcfcgi574hqXbF7PKtmtjMtkt
c8uhBT38cIhmzYCzzbw9scizvVhv0fOnyjUmk/lv4AbTI2oIPvnQsPXigAUkvRV+
bsfa4BbCMYMuzHvx5kqckNDCdI6ZVkzXu4U57EZhN6l9JWRqh86I5dvSSU+Tfk1P
7louUYQCQ7rp3cbC8ESh6NHWdqeh3dTTRZzN1bQZzPXKIv3Y8qgCfOMedxboPyWU
RD3vwkzwS5IcaLG8v7pW7zoRMlOHUDDBICnjD1dZ64Omn+b+GQYiKcKUMpJQpl1B
SGemAkg6aB5xIk6ERIXKovf93l2QIIPY+AxxIChrqwdrhDi1OxNRtgV48+6twkCR
s9iwKcF3wzziS3NWWP4cG54TDOXfGM3QUGetbDXIEZLedoBSXY/Tnkza+BTcvW2c
v6ZZNuRDgg5se0neZx74lYpxLHIHuigLNLVUS4ueFfMdmyAjMcJ5HRPmVqUkE+FW
aOEDnnZLM686BN1t6ydVXGbA4umF7sOF2vKS5Zv68iB6YvBvAFF3uFR6k+JhuZHG
freiYWrk+VRhkzQfd2ChLpMrj6Ci4d7DL0Es5+HtDiN/ov8GeyardATFLIOsZncH
fFTiArUhvMM1VpWrWn6GYAuKEMP6WNJq8S3wPkjzkNbznVkIS0LblNUCV+tkJmBB
lVNFmeTAaxYKu66WXsgK8R1hmSFrzPpYNxdbGLt+pjqMnGgMoaEE5H0sA1Usf5n3
PKv3RkBN8l+swI1PT4XXOBaFVzngIzC5xxD5qftyQmpeKjwvvzLXxua9KaZ1FP1n
75XsNOGDbtKy8wxxKUfviQA8AEUG3Ik4qYI5LeYUhs0/FWqOFb4trEdXGT8Lasob
dPtz0CSv3OEGy9SfnglJJi5VBtkLg0LaALtatKmYfyz27jITka4hQ6ZX3nOW3/6n
NHbN7FgGJ6i7Np4AMHdsCrYeQ53DEt+pSN7zWO6YJHH4D5/oIq4Bs4wCck+XwdR6
r8gAuWMHdYgGcKSh4yMRFqQhjcoEhgJqezemIY8dA6zi+7vG17gPxGSfsRV238Y7
hdnalwdXZy79uGxVpN7VweenzFXBfO0HMv7JIWZAVK2ppLlSqK3T2cHn4s8Di+0q
TkVwe79vZjQ46WKX8CYoA81IvSh+BTznM9AzpHAbEWjAcd5xlJWGeOxpaVvsAQQ3
AoND7A2FXi0CzJLoN1teRYO1svoTFqGejWa5NOOLC1I5GhpM7gYifxFizIjMYJdW
zeqpIQ0DAjJjGaorb4WjoPXHo9uleRCuuKKVBhMVk6JMWRMs/SRJb6i191RdBXhZ
FJwoI4SOpLortQEKedI1AhqiTltgJ/RTmx/KZVoo0oeR8fs96DlHmbdkF019rmFP
1VOOXXVULnzivOzleTBNxLWBQlPOUR90V/YG55kt072KrmxfkHkWfAAFy3cNbo/i
X0WYY4H9B2z8IcjZwKZpHLXtDsiMlwzYuchGKwF+LtDK9iiyNbCWREiD8SGlv0m9
dMuBrcC6ZAmQenyUEhbIuiAiv1BeWuNjqAilGasTGZ6zIkblLux9u4l0S5JfOOjH
9P6oVTo465V7xsiLpK6G7FLDQqVLjwYYH58iODWMlFUuIWI/2vdBJ370+2X1K9ww
Ov9G2ErGBH6vLUbAdZQKY0XsMChDseC2qf9JAvjFMu4t0Q/iNKR7pEZVbbNzp2rB
RznJy29Ai5cYKRI6K5NTVzWsBuq76hqmdVFpS2e9K1ZBgHY/MJLg32B4Wi2m155q
ZzpIOLtyrn48+aFLDa1t4lMOQTpuTAvall0HTQevai73j44vCR2/OKKIYC2CBJQc
9r05Wqe2i+YLngdrrf0jcimLNd3Rw//9zmRTD62OvbDFzeGVC/1EgWnfWlRR7o57
z/Uq2pbpQUHvKcuHxVh2tiKMjHTD9xXbT5adkbxV6C0ji2heOpspP0IHfGE/AQoT
OflD6tl7PDiz7EjT5Er2lxB7d76QIYm5VngGC+zpD4jT2f2vM/yPc41y9LY3+TLj
TshMPS6fruraUvMXL0W6RIapem8X0AXgOJK3ES9reJMr5sVfx9TYw+LIZUm+PNOc
EscQtyLCozwmizlQXIr7akQUOGtLPvbBN1gZ9MOcAp4b91dgjn4mwdfCdZ7HCaxn
W5LBWxbNByqB0xk+2Lib8h6H/AKf0j/KNlFnUuM8ErEzjxPvYQoZADSfQH9WVrz9
F8rql+VIySzmnBMktk3rnFbEyDlqMEyAATRoeKUy6MwmzSCgmlfdiGwQjNPexcb1
bsqkmEKVD1LIl1p+yYDTyD+wPT4iI62DZBpeCm+L0CQvEZ+EgBQg68apK2XCGBl2
ojU05bZ7qu25NEtjHNGSwxhi1eNC7eQcjtpZ2NV9JYi/WOtbt5mEnAB3EXWWTCDM
8lfbyGK4UQ2VgO3CF4X8XuqyisPS0uS3hz1ifK4/ks31EGpswdMSffsER5hN/nzc
DqHqBySVKwigiij7upQ3IYoOMksrfDNMbVkPoR1vWm4hinyuSyZs/jXVbqnAGdtC
LQeICjYisWcSV3G64LdUYeAKLbAHsIWGWCwB/ArKf3zxV5O4RGR5AMF1peL14pDb
4GrzlrB68oNdzohxRxKwBn8/vnWLyxhrW75iNK+wr0wNHEnGsbWR7Y0eIog5qbX4
gl0NIVpYKeKPBurNlxwaW2IL8R/amiJ8Pyr86dPLhMycAtffy+IvBX6S1JcKIC9o
bUt7zPTj0iI/sbgEiiO7aGuJ1B5EjEN9W4oemF9PWSPgLFkcjznV1JO48Bz4Bb61
vAPu0Yq1R/DyxvU2j6zNw5Tx0aiRVl7NIcSTY6Vjj/wPi7ZyEvyF9XeHa0zF2FOQ
0Lja2ROHkGK5GvnhQpKVuyAVBgPc/YAyaRDpWycb7ytlyonmpL5/QR9I6CqLBFya
wtxT/2uTj6KdMKSFjcLHbmCkoF4fBq54cOUlBxIBipXQeCIxcAUJ1RjgVDVnmH+M
HttBN60EmNFH35BLERW537h4518bHhiQ5gjkkNSyTOXXK7PX8ng4cXnlR4ZDHXYG
pgMIeVaRvh+wstoqcW6zVINHA4EeGrEzmqmPIAqB4MzkriIfo44EUrULYZYGPQeo
p9FYB/OW9eYGaigm2e8Biw/9YMrDiCGvU6Oij7vlGgAI8O13cPrjTNxyjWEqGQ0y
t8hV5/R0yQ+gLLKKqSFlD8443iXvfe72MDYeOakk1zxraYMrFMw4RxCMyEyKD0JH
MG58/E8kjOTs5s6l/SLQIwpF0IIEPxoqiKwzRPf2/cwr8LaDXBqzWnM4I/VCdeFG
QLKvsofpOequaly8hptJ9xQJhBZvD91OnGKMgGN05Hv9rFxDKdM0/3keZhWvScLW
PeQ8xGqvxtcnpGWIffU7pTtk83kZMI8Mud318sSPachAQubJsFxSc6G2shzcU6JQ
3ee8zV6iE/bAHHmThxWLJhD5Mu2HjYFudd9Kl+P/Q9aPWWwdYkEyhEyzDLGQ5wTV
NyyELTKxdR7A8d6dI58o8UimTdpwPLa64sxC4ogo+l1MLt7Yztl5h4vAfa+ydSxj
iO7cIgcqQbThxBs9RHBi9tFj65d44OkIqoc3bRZy9LjOlVrQXqw3lUzV1fhXeNUo
cYN3+a9CfT6bHhM8A5fgsNiW192k3poL0jw7eK23nqdMfKtiqSYe0VkhcTXmC3oq
nrR6gvJWJkhZNx2GC1UHeo8dvUyuC43tvQVT0ZXaAeaKqQzwfp9hDRZWFzJJl6hs
WttBSOn7R3nA8zyYAhaKuUdYTd+jH3EKonTKT9SX4n1avC4TgBhouqjJHAfLQs3s
FLLOHwDSQ2aRKJCvwka7MlXPqiywES//PU3WzoYCMDo8Drc4vwnE7csUFvXX6Cpw
V+dGM2y7GdXdMjDfmv/c+mcK6sUlNhF+aLkHuA4CW6rW7xZndGgV0ZXw8cdNv0M9
Oj+s2QFX7RiTmWlmHjYdhpg9gaWYgNJLNy02tFh2qZMJOYSNfn8Gh1yA1hvYnKHQ
X6CEUy9z1Zp+K3yJ8RxjygSOPabwpKhZzO7zdLPHBGx8hRSzHIrkaPb2+3KsBKuO
JSuROu5bPZZqh6u8sstkB13YPHDOsE1MbfhcyMCGDAyha3SFglArgD87pybYst0f
CoRizEt7fDxX34DZmi1WWqcnJMm2vEjCVFZ8Wkh5h5ySIklcBlDXqhjsjdGs518I
qFiR96eBYnpoeGDr1u6gQQinZ+UaYb4UiRJoMTiGKkfxI8H8LDBNpAi39ifGXvvl
+LmRWMbD8PZE7RcVqWCvMyMX8n25cxqbCG8A2r02gUGDSoLbEijqgC3gtBqCHOgu
AKPsE+fldp4ocreMZL3CxZPJgHqNGF+cpZkBEZmnU6zl7W9+mhNStzT2UutPh4Et
uPBGaZNBtFCZeQTaB3YoIrx2VCk1HRuUTuAc1IJGyWMHcht+Rlz6JPfzviRxCN6/
n21NL3hE7VlwSJE1V6W1IWiEjyawgNEYdoKBEW4oDIN0QC/pk0URdcuf/UPefBO2
9x4ZB5g0Yq/W+XMr1TyW21kmXn0yV9fuiF2WXTpFZzRu1z397yh8xwyK8d27kWwo
+nz+DDYgh/zlD5/0lWGRj5+BG/4OrL1GtJlNn6F7xHtZG5EfNfdyU1OOLvb2OMd/
M0ORWCyencl9YGghYDw6lgLtYuN5qvJunY3Zaia8lIObmcc2p3OgJZzds+UY37BD
HFpyMIvPa6FZvGgB2gq9a6F963xm8gbE7ejdgragtO6WjQuT3XedUv8RIYQhYHe2
awes1z1eIqNi2rD0Q82CN4AtgcwojlgkYheyB6T3kM4IKdznnwg3lBIwwvqa2Ykn
6u3Qbk87G8pvJTamH/5v1rZCSy1y4tUge+nBmaJMNG8URkeYi4nCyAaKd5T0zje6
Pmlqh5jZBzDq6GU2VRqL1XHz19CiRozMgOzYrlnQkaaVIepbwguv3TGHu4IeZB2L
v6bqbEbfOhodvb1Y9eLrx+td+nQz+8o+7USBMgTqPIgmdHCEKw9IygcfgeHpkfjd
mDdZZyNZSLApFGfRa0lOEotclj5TDIiPf4jUmHXPc94cbiifBqj5jqIgM11LCu5o
BpHJ704A43n7XdQSIVtsRhjIFjnpj5tKKXp2GtNL0Xy4FkruGM5pANgP0RiH20P8
WJPE/KNvhBXrGg/MTyC7ypGMqszZkjA04pQD5VuO3y9C8TRNE/hGd9QkKdeOpjP7
lcuu5bqWHLqzzDlj5zFEgX/7F54YYuonDDl+jdPXsMsQx+Gru3i3mrk77NqHuNAY
KD8o141feEvcSII36cRIJ+55jDMSF28kBw6uW46aVfUBPjxWfJyB7iUE78jln8Xa
cQAf/1xwFUbAbB+HLMfpNMtIj2YfARU7qvvVrHzUZHhbC863fTb1t8GVOczdSdgV
bXm05sN5GiHLGHVIR56NMJQfULXSkxUbQdJw1rXMSYgdLCoIeiStOAJ40+zVAs5n
HwY92+s4f0FseGk2Xw0Eh4mi8rcC5R4r1YcU3CJV+KYXpZAPSFyJwMDsEzYFJiKv
jF2ubaBzMVipVXTmsu1lNa0pIHv37EdhS2GpRP6TDqtfMyOoSFpg9XcjiXxHPRxW
Kan4aOdXpJjuCYWpmnZ/P0YAGTAa+pPvCJE3RnEiebcgJl1NRxEvaNh49k0sCngT
+bzFMwiXoWeiEt65aQU2tVvHWBD7B0WaTFUH9oOh6b4WV0lL8KEx5Wzw1sFCbAOh
GXyIcKbuDW1y15Dnd6/Lg+xEDc5yGQ71DfLuJe+3/HNmIos/tHWZ5tmqjyvsEWal
DUUapOo47i9W0KXIHl4GqQNhM2f+LVT0EMCnqc918PX5wZWZ4llU7xIJ2RnlPAg3
iqurBEYii3GoCs8TKerj/nIcBE68pDweDu5i76+1BqWFNbNybmJNLBtCtBwWfx5L
O5+Lj99FLzPadUnPeaH+WLz9nSJzd4sNLCHkbdiQkU2oq/Y2/Rcnl9/KJ9MN8fGt
Q2PsMOawdUHgPKaNaASqdFkSxcQYt1agQDwmGgfWGxdZJu/84C4iZYjubLsw57zr
c9ee3tB936JRY4JkLW76o6BIGxTM8Z7zKheEjseHRRe1TULGyjROY2b57/VfE+j9
Scxrd76lDO4nVFZjrntwD6V7wx62ufZdM4bQ2v1POjTmWwzOO+RdVRZgqqV+ZOrA
64zIW+zS7pXfledI9WWmXy6plwOE16Y5H17oCxjJvl+ikWhFapHV04z8nDn6aRtZ
19BUMnFxC+BDwQgNlhMNeUu5UpY9DnXA+qkG1XAx90Ln23C3egutldh6RgnQ9WBq
r9n8WYE+PxzbtqkerfJerFiQKY0H2EdtxcLQJPUiamuRkMb9w9Ve8Jhh3QGlTqVM
G2o4Wl370fZcWFVVhUylXSIBDnvHfKZNkub1lHmmfyEwPGf83sk4ZD6RhZfZN/Dx
oVhm0BfOO+6cpsd8bitYexlOukqhTk1Trnb+IKJnOr7UoIulC1GGlJl+DiVlnkVi
EqU5/uqo3P5vXcE2TCjCY9q2uqxx+JWdeXO1c0PJSMmXq0hJXtY6qj7953RUnk/p
TLIeYO7achEfohoAh4Xb6NT0KkK1c8FUSMe+b6c9nX4H809RjljSZQLmy6IMk6yz
mwAhBYerF1VScUpqMwXToE7KVFN1j4XT0tGRI2k3qx8dQOeQyRWMonXWL9QcDGJB
Ta2JzEjeksKwsj6mnk1VIPDvPoeecqVSzBtsj2O10NB6wLmGww98YTjtLV/4/uLL
ViiFZO9IjUdKWhJk1lQ41SyiaBrNdmq90VCrNlOusxxGaTxtjU+t0Zu54aNXOgoK
X1oHp1ETX4Kv93oWipt9p2XptXLSDO3CkHUr92N9BnmJ4bjGF/6rwNr2xQv5owmX
IhWz+SM50QGVfFYlHm5g5WIwzO+8QCcnRtuKUjuyDWbke3+KPicDBQu2UzhF0aR7
9LS0SyGTovb7Zu51HjXx5fqV2uWE3AZ27glXvQDTkAJXi7kMS4+WsQgEzD1NSvc4
OuUBkJ52/tWg6DBLi+87lVeuXF4dr/T3eWeFsIootrP6sa3r+rJKdBywaTf3F6YF
Y3Pr5A59AyBbj7RNps3OJK1P+1MoY6lu64FQrM3Xe1DB8kqGlYK3KWa6db8s+KOC
nzpYzRdu42gkc2kumQThtcbqXPdLp7G9679yyr0F8pMX88dXpKod05OHgpSTmlRQ
3qGKt4RELETahlEFvIhF0mRymhligHcG8LIs42axncTCkBDQoyfkriPMvWZKYhvH
de2W6lDoRFrSiX0TKiqWqwBdA0JSmQjnsd60w7tbGOVaLCS36CHFmg4ZsrQ6gUrz
9Uvpu7wRqtX3YCzHbWpdG2jKWbLhBNwkpeVdvfYrmIM3P+TKwG4v2QZ53Cutt4t8
g1PcP9XRD4VyMqF72sN93Agb8tJ+Nap/RlEZAtv7grqQxT9y/C8sFRMlF5NqGtjy
+Y6g3RbihEnUvzr9hdHykBWf0/VTK389+lEbuFSOcnt1yEF2KBTlq4vWvXzPQTRC
/iUWAzdz6utt1jdbvRBaH9jvbzGUoHPkyxtN3oDIS97C/ZTMj47zcfRseJa6qdGJ
Zb9nf6hp2XWIDfd8qyK05geNRiKVzHGAnLaV0bWn+P7VZ1uWZLXDSsKuGqCbR8dk
ZjLvG/xLbpuufqG34aldXAGCxaB4Xq4HDe9FNNCTP/cyEdTxP3+UdlyTxw79qV3q
6IAEDGKbHrTtN+BKjpHGXRQwev++GN/m1+PDJDgIliTE2NKoIhcrxMuS017YyVaz
9/QZChqxzJhxHG0olY8ZH5VEuQf9AQX1ngTUrJbuL+uPIPJVqEROBc1y/LZ9rJ2X
cmjnetDtKaxmAcMPNMYL5Hp//PxJOQd4C2U6akgXNcldwKY1k7d+Uj/jswq8q1IT
P82FggESAq34zymchX1+7UiCEHCvIdWAtPNkcRrRE04xtz7+Go1beyhiwGWyfHXE
oMPb4AST4MWoso4+A2vakMovCHavUDLMiVeXopLrQb+cArk4IUZePCzVvZHnrpK7
E640aMZaiumfjpENcFgoe6Te9czz7wg71Kj1DEVVAuAT5jr3Xg5qNi9c9Y5fAY+R
3kntUjpbcHpFGcgOJryWcpjSSLp3IQVP2oMhEUl6VYC7fPTte1eFiflmlEv6J8e6
Ngcg98vjHM6CpV8zThbLGoaQHVK6EZph6u+d7to1c/zESkv/1xzNqjsl9o08kMvg
+cApPUxZlWjM6w6dUarbx1e+ahU2ZnV7X8XzqOq5B2Uhbg/dhYGj4jKgxo72+GOU
YT3lcMTOjQ5XpccgskV7wPE91GpJ1Q2+3CzkKhH3jyBlBTaRtHY5Swg2PzOVe3Lw
jNgW2FV20kS8HpDiQ2IC3W8/ftklEKxo44FW3Y7o6xqWx5Hd0CGLhKH+M2p5gjXP
+6Zk2uTNRO/CfOvtL7kQ/vSVXCwmFSmZ4FQxF+95gQdUmk0O/l/UkVbebnNW3UD1
kWbvGoLIhPKxyqcxv7cRo2efkicOMB9k+iXcGcF86uBvLZ48k2uEUdzOLDMxptG1
gz9lpkWcREjn/fDD6k3TbauoW4Q0Icvg3ylthXci+WPCpN3hLG44qEreGUAmupBQ
hu2XgoJC1H+elzCCwe7kSvuplGk0rtpOiKFmhd90F4Cfc1PNhd89ptT3PkU4+F5l
t3M6qda0vj8kE/g2hmKgqgImLuB2C88eU4D4mynOfvfnRzeKN5jY54onGcfcBmKS
OopnZ7iBwRy+xeGMXrudcG/H68/iq4QFo3U2Ryqj6uA2gww0A2iohu0wVFTTEcBv
bKJa34isI9zQKLWQjK8/jXU4f/46NIdhpetcI6xTHIa8QLqyyAFSIq/EHgW9d53A
89Tw9OqXeCmtb9OJ52Txsv4PQrK7+LvRJgFgb0RZpbvMWHh/D/lJV8eRFKDlcmr0
QJziIkIAq+P7O9N/VVghnTV543Oi2IvGd1Yei1JUj9t5jHmbQJOZxOJGUNnsEfK5
YO5t8mTHUbta7OuQAW15H3YDBaqysRe0ZK35UvGxPWDqmpDZJXQx+skrzAxcexmJ
2UUEVdFHkSwv9brDpJE668kBrsSyC8DMoMuwFiUxYG3yR2UJQ9fnw/6VgdmF+5A8
gARLTDtNsKLqDpG0568jH5yDBPkv22tJYRkTXTluTvHC/8of3S1ybWEsFoho4ahk
dQ4hZgVFY/VJdp2O7oUO37qVkdB5ZQOs3PM2j0jO2GzImT1K83S/RIliaVB1kxbY
BrbaYAykcxZRhkN9GAaom3nC4DjvxVy2GZ4dIX5iFDJel4ywi3MtecxzGLj1xvjF
DCHTqyKfENfCSP8DLTNHUJmK5otgtit90wJndeNZhSdmA2cl8p+wOhtVDmyEKKkl
cvywxowt/VtBkyww7ERwEuT0JsaM/06CoGq7RhG6o2jgw8nbrTBgf8W8Bj3n0/VA
1AztJqx+9NRm2WmREQHgRnbP/cvlvTFNmR8k9ujXtRbZ45wh5HeGyiBistHZ2zJN
ehkpLpTPQODeqgmLKekmjDdH2juDpJ9KIKF9hWkfCgLnpMJ8qfwzg7bwn7ntj76T
iXF/0+74wFJC/QukxPcXnS5FV9pEEu50MTA7ZoDPwDDaTszvqvikxQ0I6M4C7HH5
QqB343oAQfCH1VcVqWS+O2j2kHQRN6ge4CRiAtmPe3KZ4FMY90KQgUx4H98vM2dN
vx4aFwmrydXVFYy6fy7tmALbW/+nqoaXi7jH5QUEL+j1w5PHH8azefb58RJUacFy
cbWy8D4OXfAKa77JsoDxbyBfx8EMKWU+tat0RO7FA6IGn2y6IxZ4WNTuiG/8JgGo
Cb7emlyBx2DXJOCp895ZGN8rCH6wkLGBfdVoQO2R5XqDKiK3wOYqJxeuK+jN2TWW
x/s24Y4I3o7UjK6REzRGEh7s3mUEVd3yjdvHHOlm9tNxBCK2Gm/YLZQiSL8CK6+0
P7zmES/JggyT13TE32CEJEi2TVUn5Kz7RDgcBsi02tH+JwrV5kDEQ6plx3WzlV62
nd4F1Np9QreezkY+epD4rv+cmSeAS5yQ2am/r5g7NT7ZImJUQHQnfkQsZw9o1cw5
LQsJuPEng8U08pbmT46AW5AhlMV5jqu5Xryqxwo13Hxb8y+2vCsBFeVo4ZYTSB6z
cvSRDzSLFpbcHwOJ+Na7hYVbqjDJmd4aunI/091kciyCFfd9+TPfocOjZ8FKg8hh
8CtsO5b8bsxaqn28mCdua81gd2HvhWr8Xdu9emsu+iTBpKMLpkFWdMCGvPDUbgGV
GguyuIamjSYfHJAW3Y4xZstSzA/qy18pCckLHZq9T+/WJQ5rWLJ52Gzoadi/lkso
pjDptp41at9YC7S0N8fNAp/VttS7CZHWkI9V6N/6pEk2Q9hGZBKg63zkYWW8iu0p
gcIwc5cBhhW7YS38t5PJcOP7l3ktRIZptLSa/2CE8hULWNMOUvsSGWbimzgj/33e
D1+DmwU4wZDzB3tY14GYPUo1YafAJI7ZSukGmEASeevK316lJ3kldX0cMaw6GdJa
vaobIEpPK2WUSaUgLzZb3NtbNJjP4dAH6t6ZpSbxm24qeq5wDwdyxubTAoVtPuUm
Oq3y3/r950dTQLHa1iMq58ROJzUJkLnSKtNwyg/jJRMaC/WJbnkJ+pghntP5yxSs
NS+/USLNXKumTxqHZRgEBFZ7PwdxAzrX4+J+CHSgTCAREgmTrJ/8koviOkU4bMfk
MeGJ7DgpjiGb3aOrqNxLBC30EBNJAfzWahsrSx6W6CTKPnb+yelRa5d0HxKny7Gb
uHRbifLNn2PjmVvVhyn54G4Lh7hd04UXJccf3s6qi6DhAZBJyxcm64fzhZxEWfED
crXemXI2emMHizCw7n3dp+rLg5tEZv5PZ+25aUSxqApHOkNwFAdIFgAw++W5egj9
7efwZaWqLRApsNt5Pn8S4J7VvyyfllhdEhD2OpHg454qbei2/k3+YyvgZ5HyucyU
wHJMjaYV1n6HwI+/suPpmq/CptgoR46auvTb03x1CDQ3Vkndp9cpddDCRE6fqhmd
wZy7jmj9QBnOU+4BWzPzTbWu7G4HYajUTmjopSG6H5OM6Y9BVi3thTCEU5J4rmDS
z6y54GZU73uuv6+fZiy+T86GyRSdseLM6EG9gYvvNsvNbfNG/6VFXfGXqTVPLu/+
ddSgSPW5b9cirLtlDFzJsQAc2b7xhJnvCJyDweYFk9knRqGhxDj9x8O11NglJ19j
S7yk5AJeQlLEfAGPYwG5og3vkG0caWxrVpeVaK8TEcFay6BIix0YZYoPGzZ7JJiI
X7vbSC9HdEtF2UA2FFAa4WCn0DrNn5WeTByORoFP92HPzuJaGcaPYhOOoGcr+qLp
cgK+r4bvKILmlf/e6UnYhJHu3Z5EZf6LHiyUU9agGnI0jVCL54suqRls7Y1XfGnB
o3aIXkd3pQMWUqC3pw9IfVJO+Y9Jao+3P4BUdpekVIrKc/EB0NGs7WMeyJCMDAjO
oxUfLT22voyWfSlEHYU/Fm0Gub5oxJvsev5EoU2koqo+8+qrjVM9x34kSTdE9jXv
X9CwZMwOJ7VcPHKXGOMKiHLsDnw4Vs/NGEQ9wCPqOQ6pdmsY/zYw1Hl2PyYuz+Z6
jfo0Ln7WlaxMPrzbMPKqzjVBu03EVoUppYyhIyXOISr+Z6WDE9PvJxBf0OXI6E7j
CKkhFwWJwX0Bgmvrz7L7Qtw7YtZcq88p1Ougv2Kr/4DDmrKO6O3qD/sAFUQVOuCZ
EDuf8Mb1XWmK1U6+FmPzFXk3j9D1yOYckgJ6Vyrl4r7dXdqdRqOFOkBfVE4+Czja
mR2D9gPmIPpMzkIo+QMqm19AH8MfnoYBbXAXDdLI2T2GL7Z7fAkYfOYOc6FdKzNx
24v6o0CR5mSE5cnXo4vcZd2TTpqus8RtuhpwY8WUsFrKkFI8e9lEIUXG9ZQMevI9
AsOAmZG+2hKhvwpWfUPW1YPt3nZfbX5efBJ5NWJa+LV/C4Ldx5JFcXN5WYbVBVyC
pSnZTFuJcyFks5dE05TTdHIZbWGfArLGzUt+sSetIgzeab/EcGGywg17rIns+a/S
3aWuIeY72AxrAtvEy6oEPGkQPLi3QAEVuOo6s9J9DVmwpRlJU5r6o/wvGMA//ihq
cwjllKeRsHWQ7QbLM47wZAHYfAhRrDhSFjGj4Olweq7VOGROdo/rBjtNJ0F1UWoB
wrDb7gnCorMK4WDMeygR1IzJJt2sNT/wyUl6Okzdid62UYs/gokkp6qGhffW4Pj4
/6ZQmMdxUCWmL4OxPj1iiigPW1a4ltTgqqvq2Q4M4Ooh/iFHXRGlnvloH7ytJS8q
gHaYml5pSuAWVMjNB6IX8xyg33pCkwlpUrC1ScsmjwFrgAR0qq5xIWi+tFf737DE
FFI2h9FMQOZYO1DEDZTaAksWYbDxAsTN/AoHDlfreIeOUAEu6XsvcKHslxvkmzGQ
vLiLPCrFhiqPgcA2/UDL/DIjk5SupErMXFYrcTYJSkEThMPEFKCEHw114pJgAf0y
NOtNgvg6L2mAFRgUUxzgPP06m+jDSvQJ+T9Hzza92n7M1PPib7OM2l4O1CQ3i8B2
psgsO20ibSKHnRVRhGbhMkeC6YOLuMuABrvn08QIbz6vqi4O5jR1gr6tbAzHuwzG
H1h2av0hsa1uW7rDnS275TOMpkGqJYJ3wyTqfbvvEKX+/EqtwdWvJkKvjmyHQvJi
TdGaQ5kpnUEL2DnsjExdugcZWuInhc6fam6E5l+/PS7n8KIy+neZ3gKOldMyxyQf
SYr3ABi7tUi5ozZv6Mb1FoMSEo2lHOHw8XZispz4mYtC+WIRXpVU2LIJSNfMiBOZ
20VG/6n4queFIgE2Yg5pcFyEC4lP9KxhSiPWVy43yP/8dQhAKQ3Cgy356i9NfvJd
uhPjqJvcb7P75wbgHodT3Ggme/d2RuMLBJwUAS+tf0olOBieMq0yuciBmrdKPhkz
xamwKRRKJLrPCPtqORL44+mfLjr8PzV0FrBdI0zopkf7YQKxXiQBebsUisMguAEV
pHpVP8byHsHXeD/Ga/y1sKq2vrJua5Jo7No4M4S9fnt9HhATHHEcE1aUwp4TQslC
Bh/UkJ2QNCrRn+8bZPU6fs2MeV1F0lVlesT6Fnv97dIkp+pyr22JHk0jxO8u/U3t
iGk0OfZ4ik7A0E4nyZddsS3kX/KzMdWc5gtoiti5n7GkQNZUYaSryTPlGeGdlL5h
aEcbsxzF2lWbythXjJXaax8UkvKVWCxm7YoNyTVWfWJIkwvG399hCNmwuwNPDmv+
/2Iy41st+NL1IB2TSfZobqJSbotBUDmt+qxwE5/D52rprHeRIX7Gievqm823zRfQ
L2zxmyXsVkPaWpQuv1siQMiHf9xDSgKHA9scLxUCs7AgcEbP98VIk/7BQQ1ljqGV
5ijJ0JTW2SyzW7bViQFawD5HAD7a+invjx7EyrKchzdKNrQJX09Lu33nN1zQni2G
j91ThWOp4gKwieFKdQKx1fusNEJQEEIzX5w5FzSkK5Pdo5ooMEfClzibl+6wzGv2
N/PUL253V4MQTRCv/CMPYoB6/hAUdUniidQ1ZJLrW4EGVzxh37a7w/wH3i/41wya
wuw5PiA5rFScWihnfzK0HgM4Rdu9f11LCmGvUt0I1csXIxsdVwYLiaf5lcxYW28S
Eb3/rIGLUniYbdIDsfqQlnRfuJajCtX+9jixWgYxO7QxQV8WVzk93WyYztEsIcGv
Onzs5IgjLYZ3DrF4rCg9XHMl18QzXvCTxzeG1biywgaULHJL3nu8JRkOMajba0K4
pszLkXXJ1BBTdBZXG4svzCOzmB6UFvxhq3LXbm4skU5w7OoqrmllCtte1DVBLJUY
LrgppIA7tcmvxHMNG2x9zdm3zZi8SYzRdzjj2SfLq4mSrNlD3+QxFCqTbraoUeim
IsSkG4aMlensznxJP8LzOmr+IkfoYJJlPLLQT8uUNEf8XTEsKDdXUNQO8r8AFp3P
7W0DVHktKLee9QgApDeerSWzmzV2Jz5wxBn4sXuVVF9M99clKIt364ePH/iv2zIe
yJfFWTX98KpQMfezvdrcqHw9+CbLj7GLOkBejxMd6LkIv/jKY8lorlCOECPmSjvu
+DRqZwcStJ/08WS9PtGs0NMgl6kbXu8Iibse5ACcpyPUcwDOxxS2JlOfRMTyGDrO
OPR4aFeDDcqLYIzdTPOXUSU2vThOZE9ToXbjCu94HlRZjWeVEtbKR0UZYAPbx6GS
fIe36zws9X4KNunUbieqBOS2pPx0mnBx2rbmuWY8DLVlOiLLbWUI2/LwciySidRX
jW+hNUrZaKFWsvLtX+5SfCqsAIefrOpilnG49lu8SVGgZ8j174GwooVM0R9vQUNm
1vVySLNt8so33d/51ITp7xKQ8o+2z9Ntr5KSfrhwJjfRAdLC9bUDjrpRwUH/7JfH
O2zdZZhJgRCYvyOLIGySsbMUTWrX4MXBYYTu9GhpmHY0l74qdAViXXp4b8WnkMys
xUX3r6wSmhvJsgIO82QlKnLlizmURTg/z/I0rSZJGn0yR5l8BaTbHD3/PSXuIl/w
2RJcXBLt1no2RGSY0Hs2RvbQYTBCekvVIVn1jaVDA95EyEuUxEWS7O3JFMFVuMMz
0uE4tCvblzTSGXpI+1FN0uJecLBdrm/teX5IFjCCUTczWEzCN+iRsaAEhxv7qZAW
vr5TjofR9MmvBCLtjewy/klJIla82hVHwT2/sbl40d40wJKCNkOCySqznCzhSR97
6ezBDQycpr/1bysYQd8s567G5jmb4htEfVntff7F9p+Imd5m1jqDr/Hdx3WzeYp2
StvVATCnF5mwCFPCM4GWveryZ3NcFWnE3s6vEdBaaDPGLvg8o4h+hd80vi9Cyi2L
SL3vQprmV9mvGXNvOhHKVQ==
`protect end_protected