`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 22016 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
FPPR7ws3fN+RQyk1V5tkgAzXCgALhKXifvluKTu1nv2lhEtufvs8M6DBuMoaiwkF
AZUnsiix5MJ0ANcZAJnD1qXNGvhPcV3/mmUanadRy9TPBh7XzRzn9U1+hAhZUdpf
3LveEdaYGhKRaXTj6PUS/3g13sqvpr36KTRgTDc8jcY7a/dB5QdzqSe0Hnokm73n
ByfVkMx/L8nTpI2lwM9o8dRRewe2yT438Q+sddaoRnxgWNrPDJ8M+5TqA0DvdEX8
SEaNy3jkW7PY4WG1MfpalpkAnIKb2K1TD1zSTnDdbYi/BwfP5ccDW57bRFdYEHAk
eL0rTRK6m4/hQ62+UV/+CENImF2nJME5kIvcs+mgwrg/z7xCl0b/rAF90wowavJw
PK2tT3z9UlUIGkRDxnlNT1jBEzGRVQB9usgazMluHmElUs8QdMW8VK3aHeg+1omW
z5Qt/rzoSfBya4vI+CXKvK0ifIGjhLFWEUi6y5oFu/Wx+sTcyIcxuzZ4xPY8BLMv
l4qibaITjBzJ8dnadWYFkZW2WdIupsMVtpIkA9iAH0oac/NlF4DhMee6ev+gpUZQ
t2+tM96Ntk4VvSp5mucKPIC3FXDQ5ER89oXdIS9h5LbHiPj2WlPwlHO49Dq5CV0G
wSKYNWJP+yyNQZ5hRPSHb8toCvPMdUmu7GwOajmyuRBGbE9S1CmKDDmVkxonWTpn
XXllhgBkBm8YSexui2cR1lbFSKfXnrkep9ApqL0CqmpQxSIvJ2TY1kZgaPYZtkmP
xzC0Q7j7Bzntd376aKGa3MOvrRWXrqhb7ZFaFUyuUg+zWENVK43lceTcV60gJ+Hp
H3JEj6W+A2ua4F2EQDEkGSt7wUYzcqE1rsKXy/ld/v8cBI81udHqNQJsSvg7YC8b
6b7x78WGeBUuSs+aeUgf4P5TfOHFxxaPfevwzAkCCs3+wxKrHZTUwDSLdQOiI40L
/hEJK/w2ar+J2Dw9hhOJtx0FeZtMLFQU9YwlLJdrbWFP4ugwN6jg+dBKSpod0Fn9
13Ns1mgG+ddRpqySQ2X4h4fFI6OdDY4ea45NLnn3Sfion7yi8DlVKZtAAlmkqKNc
ZfxkUhfS9dqbnXL9Mv+xTyBLIFhGWSCcssm2sCheqx5cR7+i9VVHxZLBJxcYqNbS
OdabiIcEFlcYmaN70UkC90dmgCET11szgMpMNz37EgPsGwGWUAPa/Tv/wQhpc4XT
jvLVuqbc/+pm/1a4YINp3nZoxxum6Ix3/WUlhwaQz0CSy60csuMzApRbAyWotmzd
2zHZKR2dz4O6rk412SF2hW58ARm1Bge4+WK3UpdWQYzuiKetm1LsXVVhIWtA54oG
gmRu07VnT/Ep4TbEnV3mhSHcqxRIaZhSULbCAFJs4vDkSmgwuQSp1HZL16U8/xmH
v9pzInNbDssOUY/Fz6EzyXqmcp5UMB18L0ae4mtxCh/qAY1vaF9CrFYlHhOy4RBn
ed8F7A/6mELH7tXSBXl3bxjycIQQxM9VY/0LrTfqgVLTqqzbHQa80qCyRUTGalzn
qgZp17zj/mtieemwyz+yCTHFvnHYvbqioydI2+OMjYlu6MoqI/6cPUWxZB6dmGsA
6I6bS7+TLHABuFfIHBivcDpDO5zkuXrK6bpYMOjgbqGs+tL1bpJQNMcSa2vZaDep
vACn4hmr5HcZVX/aLYmBafYUq4kfeIcK5yIWPk5dFuWt4dTCO0iZDCN+9Rvz4obr
vJCknPxpTxPyfwB1pqGZFYs08Bk148G1xcGCZhIpR30Fmz0KtovI/93qFbf1ulut
mGDRqjL4Zpd2/tfHmMvV5Zg6aYSUBYhRzzPtfweTPFOZ8j/FAKKYlpamB94qUz99
pWnRhnCoOFkuZPX2UlSXYmT6FxEWMeeWqjND/aw+wpcZRwMna2RNqBwwl/OYd+yB
razsWyJIMUyc3mma97Q7d1Zwy211ceLxZt/nijvlKYfu+6735gsQhnSyfEQJjyf5
bnK230bCmpg2IKx4xq7+Yrn119JoHW8mujVH+C+EHk71IWn1OBwPnq0r+fdVF5mB
CPNaJby0kXlK5ybObXqaLkhMgF7d0ZfnW1ufGpf51Y5wiTLlCKBvUTJ1Z53swfwV
qcsZdUZ0TTpzaMuHKkdQzA1N1WGjVYPKwnMqM7yYawtXlC2Opu4eM6NoS7H0+usx
fQKHj1cbPQnj9vG+VnVT7OMSNZgbFzHMpOycdHbZtF37n3rGbzp0fjBFohxYO7le
I0wylqu5DhO+tzJlOhoilpW4bx/0grfV0E/oDRbR1K4Wo6sEihidyIiwrOWWHLEv
MlJt48OM4FF5/fpHctWZNFmTZSj08POfUS7fLYhPcQaWbzwSNnQNSs3vZ/qU24yT
Y0bZ8xbeSLjUTT3j1l8Mxyti2Aw0AlqtyBUbXK+P4lK1k3AU5ddDMEU5tzJU/o/h
EMLwKqMGKghFfMFpVj3+GF6evZbmH8LDa094vg8tLgSGbCG2Im9DxQxASQVGgX1Z
feuuxHQJGYiZ/woaYvEaLtl/iyI+oIGF9TlfsnH0iuXUmS7McH6lmxP5aLo1IOkI
cjLtzUMn3wbBNzjWmhEZ3SE1FEiK9YPPZe79NPfFdAn6oKiGXdZlbwjAnzVdYqWq
Slii4KtvOlcmHURpqWT2F40CEqaj9rdl1PDu9xRC8DCQevD20ORlB+rzy8URIBAM
fXs/u0J8+hPwr8K324qpjHD1dmdVwHRbsawrt+omwePX3Kb8+negwCk8tSUin1R3
Q6mCEQWAlO1BsppQoUc2gdt3zxGQNyd8L55Z3p8cSln81itfkN0o44sgb4KCLL2f
ZFIfY0oWJXy3k7sbP4oXb5r3NDOFvnn/OIGu9hs5u0Zf026TFj4eYjJLMHvLwlrw
GBt3GGLqcBnEqLBBXpVVAipbDRzFXXFeGpZ68HUBGXAb701hdVJedmZUI5esq5hR
AhffOyRJtenz7MAIU7yL99f9XSQLajOgQR1xQsP3+VSYTVU4v4HprObNktWuiJhX
mgHjsyYgfjhRuwhLAydyTL4fPsWQAf6wjJtUdeuJvuZxRC/By/cx4nn4fhDl0wCq
Q8raK4E0MzY7mPoXMj+QEAlSiRIzCkx/P+Q/yNDnUnTtYWItIITKAwbE1BRPBvyc
d4GIxjV7eCxcAqHfmajeqhOCC37EtCSnXHCL1+rY/J8u83tM9c41ozf1KH2t1j91
0T7rCDLcHD5TNY8lzTuIPMvaeveGzHwSX6lUtA7j0msevT1X4ob1uai7+BsCL4P6
EDVVew8Q3KzqIuS0AX/JRGFqEUiCrGJLg34S/5X2Q1ExPiALFDsP5JSLOE1bpvQh
t5+Psn2OJTi80eA/xgbTsTRkj1GvKmxSfLuz62HYfY2lbkRZ8ySFYOXML+aCGlbO
1Yc/A7oVrGhlbsblI4MHRSZU0jG0LmwnAF5Jom0qH5nmtiASvY/MLiBJQRE5vgcp
O+hHkS0A7HKAvOzdUueuojNjJFccT3+9qZCBS35orz3oVmS9PebtTgbu1o0Tp33M
udrJfEtxICeCdByjhk0dPECAfkkynSPU9jZIqAIX8JgFEiLuAWadEHEOHoZl0DcQ
WiYbjy4gfnHwV981gc4nYe7l9lIcP9MgaCEGdpkTZG8pTK/Jj5G4bxzT9bpnptWu
4trNfJGa0F9Yy3FLKo/f1Yt31ABYdTNKV7aPh/fh5cfyOr5zliFgmVZ5+tHS3Pr5
yf8+wz35poGFFj4qUZqhk7sENQQqAfuGthhkG1DdI9oSYGjBfCu6YJvQF8LdKrCJ
sBps8W5xxXbEOUYXDUuwFObZlJJBX05Cwy1dSBdoQLeQjr8lbBlvFDxzEjx4Fhl2
DLhN0Z33RDzg4ipIvuz/hkgnKuZFtkgQJu66PESpZqf3ojUcEpM2XOQJcUAuHpo6
UM0IhUFRtRdSv/bz3XvGsYYojywd7akD8wkdRbBDP1otP6i8zxtDs5Q2IeFMFxld
+4kP9y9faEhqmZ0JRwztFzT40HJMeDxu9VBCPEeKFhRwhSY5D2F0a+G5qZYVfMvE
7OmIeV6M8z1YQQnWgku0qr8nSNfhXA7+C54RXYrwRwIhO5aSP5lur04k6oTS6vJY
qDDDyroEJUhZbFpspGaJybIAClRPDVQQ1dXoPiQaHw/tEsKX/QQ4qoCSgj1W+U3L
xKqXnWshDer4O6q049EpJwJj8OCezOonE9ZO9cMF+2VO/HHQVjvCleH/6cp+Kn/p
MLsbQbVJEn8Bp+XtmwdBRlWPWB3AAQL4hOWG0cuNSYXcTykw7OyLnjYxQx9rQ7js
Qn/1v/LeyMkceqna34WXVrc/upEJPwd+jRn08WLnUp2L+kGnPY5in9JrZSf5DmQ0
71yOUcG9O7FSVWvmouRf2nOOsde55lsgf1eLQhQKUvjmj+tbppM19rlPJW6+Qwia
1zUJQ8qfOQBmDMMrHeeYhUXDQdf3Q2t8m5UsDOdrNx7KiYhjGTJpQqc0DOybzJhp
llG0O8+cowqIUc5P4oLJZ7rbhxbp5X8sc9wX0oaHeNeD+hCIMaW3GYBecjO5yGsF
NlBz3YLTBTDe0R5IoZDDAAQQ9S6B7DyWk+cEoMI8aHdz06FUl1ZqMELTYxhAWQ0B
uTReGkvHe4vHzqu9tGUncxSf9e47SjCGuqVsw/RE6AOcW+d9Z8QFC4e2jsUUNcYC
r1pvPnL6n23HLNQNx2g+HTJJJPHZ4qIl597Artx+gxbeC+FnSmJSn93Znzw4nvdB
V+vD/x0Ahe9CZ9KW0UEnv0bANmAbl6deviRI/6od/TTI51teZUjaJ0f3iBT370HQ
qj2UDE+DdLGWdIIIW/vxmlek0Tnqa62zG6lhjNuUJFMKlxvgMMrqyz9+2FIFDSrC
tIaZPqsVXwwCII+OS774JgOVzBA6wd7/TKa5xGBRg6KSAhYUU1tufTEE9IBeO0C/
CnXYznCExYF06yZ+kbyg/wcrOZ1pHtuBe4sq/A/iPg46lJPO8qGB4tBEbLK/JTGE
dZ6QX36T6UFf6ifus8LxLy028JgIq0IKg4mpZT7RJwfIVZFG9i++WkEUdgqcQdkg
xVFL4C15SwpekP23gQUhaUAzFUeHx+0/BKO5AoaP7y5lP8YbCbL0fVY+GVMvsA2i
+B2LbrbW2rVhudCXk+XDCRexQLnCo2AHsC5W9VcsishDdycdFL09r5JY1FImVpxc
hROGHkHT0qokhJIESxBvdAW2iNOmgQt/y3991H/hnst51ST2un1mivbbhO26bBdf
49m0HJ/Zuu+26vURwUtWkIss8ySqJ7uLwAf3QL0BKov1mVy3fIkWN6lNuG2OtJpY
stLAzr2d7ahA0mWkvjxxqjD28Z/azkKqXz1rrxsT1puJ8mCzoL30e38ClE60KvlF
JNVOU8xh9mC9zdAyWhyHg0EEKGNmy1YyBP39hRzT/smAT7Td15PGdFIBV5BQ9SkP
BgNoI9WfiDU0Jz7gdJb80ub7z0sgIEgyt3mKw3utY/phdbGPJzln+/GapMWzGpXM
bDRljCNlS62E6u8QT/2coB6UlyXc/4fRMBORYFFyCMgPa3B7KHYEruP77qU3N4uy
nMUBsLQ8wdPXLLHrJQhGuZkjMsj5Cl6TUNDGhOps2nW6R/u+drozRQ9uvifPtb2p
cGASe2OGrirxhc7N2chPZ+fITE5RoKBC6OXZcSPgbn5axHwPtgmUpJhmIm/se9ko
kZPLC26gtl+/Td0QlXP6QNahBJWOgoOyC3X/VxfFXdA19eAtvFIazlZWM1rBgcdc
9pbRRUYAnkrtbCbwp5diM7St1GzyoUTyUlpUBjTJBkgt07fFgCvCSneg0JlIX665
6DP8TKo4yWexsnmnJcwDnIfnTOLrd9jmLTZ/TYW++rr5G1ASzzM3DpD6RWK341LD
O6mLyJIwhwr1XScRGFKK7jX4QNKta/bFJh4gXN9Lb7t9QhNZDHIygplBKt8mgUO0
/yM5hN9Tr8nUEUpyG4SmDYtXjewp/XBWOo6v/lv3RqCswBhFx5h9IIMQJLO8pPN5
2bVy15u64e+tfl2UMkX72BLS57ghIoH4CXR0wpcWA/EAhswBz5fZ0bcb2j4jct7X
X1Nny1xFBqhi0IPWxnv7lp4OU4bXrCfVWK6PSEHw/sDBhiP6/hTSP2n+Ev2prheE
Z5d44wQsmA8lqPx+LDv8g0sqm0pXKSSdz2Dp6cTDeB0DJ3KaGW7XABUbN7W05t6O
2YgrAwzE8IkZw/rytp1W3isRwM60WvNLBmWy2TcrXuDTcF/qCjw/gXH3vuYobwEF
k/9uElzsv9Q1+cvKkRO0VtJSgQpukvVUYZeKvSd+G1whBkgG/AG7aQE7bFG7pkID
kBSPVMbjgJfrgqLMVNpQeFHKPnEghbLbWBEzODnvo+ya4+nVOfhWY5KVIeR35B82
dYnfwdy9TqoP0dJBdqa4Gd1jCwiFgr5PQvAn/UAiPFOkSeoydjcA3rSNshdxqlx8
a4zUghgTxpJj2GZ19HHY4gRHPrnsmOEemBV36jC1gCPgH1hX3y1RH/CL9VGUjlKn
lmNiNZxQOxv2m9C31eIkZg9Ucf/W5bUPK3A7C23vsQ2PNK/KfJWEw0ebexR65kSK
Rh0qR72RmqSCOKHUCp2AvCPdYQgO7FHrHnTOyTY2sdpzdQJ6658XRmk5xMf1Vf6T
ul+BX6P9bCNyDHHLdg+ekl4TRgnlti47h+ZdOq9xK7YCgHzLTTod3K9UbZIAxZtA
Qiu7SA4mlulYcc1To7hjrQAGwa4plq+izhz4Qdu8Dxk8MixHCd0VEXFdYu/tJtvA
DU54O0tB95iVUDvgEf/eeVzlq5LEiuf/pGGG/9XdXol3QDBepLOaJuAGNd/S4aTY
CfTqZUim6MSvCnJTTTvWuYLddG/ipBhotOXBi2mui/P5LjoL0SQVwI061ma47tTb
ANLIAQgCQ/LTR4IbIdWtyMTgkEiB+Fk69qExiYfco7a3QBIrOmYjFf58afXEyQrb
OefRGBSkzbUEpoWEduYS76L0hjlrSPaHF3lhE25KhPkZ3Ws/iv0Wqj0o6E2bexd/
GKq2p3E/YFdrDOptWx5Jhoqq4kTqb6dBIpB/hAv+sIpsGRuRDEP5nV2ajWQZXfid
2nOZ2yj+4OxoK2fDVH71GTy3HWWhzhgLHOBfxaAAVDL/1SH9GlfRtf1qja8pDGNn
KD4pUKkVosSZJk3QrbDy37rIwlW7EAKWS67mGcAYRMu7hQYvjWUQS+GL628BqlQm
FgPI5QYZuygS0qhtq6dhpz1NXwQbH7S4iY/wciQbpn6HHETQCcnoLn+223YflP9r
bvvzCtcmeELEWu/Ss5AFgQNmA+USxgVT6B1kq87I/YmA7rN52/uPnOxXv7H+Zi2p
deGP+tPZYEnGT7RYuDAAYmJikXEew7i2pY3nuHu1HHDf7pisYxBLtQ2o3ryQKdkP
LwtLGf8kP6A1v2/rSm4ZMtUpSk3tbZeUVrSkSvRa9qxyvWT1t8dTlPv7oyEPn7AV
ndt+bjYHUQ1NrUbiI/4tK7ByaMVsaYLqQhndAYZvk3VMPbkQfUWEobtFitrA4yHy
U73uiE4otnqKEPHWtX6c4K5YcDuDk9xLan1x8MNa14/zIZqBzUzmmuFfL5txk4kA
NT3aK9AJVEi6/Wrq0gqy1cub0gq/G0QSKNNt5wJxjG6bM+F9TH15p/DSQZ6D//dW
oJyo01pisgUL04CYZ4zMNKZmJLUb9lH446tLu6fykPo9PXZec5CPtKCJryggbBlX
A43P0wiVYtbITTkL5OJzwgYi3bI7A43QIlilBd5wpVzvAp/CHRy6ZcAYxKCCKRag
N9+yGF34M8rZg6VW+bl1SQWUfjpFtOveArba6AlRP5b0pOPYYAzx4maoDymloqRn
1fYuJ60XlxgREcM4cJ9CbW36HL0SnRyix2UjcKl81p+fQCVzLoczXP3zz5jIsjUT
YP2lJwlMTorCaB4lvQWG+Uo2dFZ4k64y6yBb9AMDfpNYq5FwvEBAuJxc6AE0D2Xd
XglgROcovK/XD6yu0gH8biXX4M05E/MV0ezdiV4CuPoLX49l0RPJi7mIMASB67pl
YbvWeMQ2MrSaSPzcfPpYU8fki1FDmia0ojZ7Mc1O2XGaRdk9SsGGyaJD7pc13X3o
00HHrYHh9WeZVWkIUUp00HIYoI1y4AaSr6WW8zZUYlTaAYhsm5k3/6QhXe1pA/rd
MBhOnnBMwRKbiMmYM8PO77p0JAnvBmM+7K0O/oajrHqpVYJ3OCs9bA3CRxw/SHbu
Mip1l6X3TRTMfESU1eJnv9Ko1bk2iz5bmwbpmmIm0E4DXjMZFcPbHc7sekh1KYbA
81T0ou7vjI7Gmt4LWmGfAp7qEYAL2HIAEnJCZOoimio2/206O5v1aRW2hDWSb0oC
Fk7Ywz4nePWFZX4fKOLXQUBYKg4vXBCaebsnN6VnmmDw+1DHmIkPwYm5fqnEItpY
eIhI9/T60tihFPOJ+nrP8WtWB5d6953kA7YKYRbcX4jN1nLzS6c7bvho0FW9xXdc
aTounAkCaYZOAyHf5c+/I1fpDZoKnf5faIYXTxh3E9TuQF4ApxozX/Rx4wVocQu2
hR1qlSTE6MvBLbttorc/ES9qTCgMFZwqfyRb8lFMucFkxU84VXQ0uTygydcetGSK
c40xT/tijmQbkigBfwm5artBUDliANGWOCwbOlfA4ZF23E2rHO5FV5v+S5JXXPQ7
/GpTM6rDmLqO2LieyUr2Uq2gWbammfN/xxaxc8HyhW5BrZcTz16NXB/ut5xUURNU
btvbkVkh3HYVxGBo2cOjagPBY12yvnmkeugszRIEKIqFxcHZcTplmwdlsd7rTOqH
GGwaoxS/Bo6b5Hm8OxYQFiz7T7rB+IE/4RKY0sJYz0CVxezCiI+tjE8/7mfFEeLa
W72CP4TUHFBtRQsi2vUCMNc91mttjnhafDgQqiNx/a5U01dF2RBfjsdIxlXy0/0O
Q/HcR/haT7bA40IifYPVNVd5VhMH4ld2Tgl9h2zSDEMvTqLg7d8kqsi4WBNyUoTw
RsltLeAs9AVmhQMTxMvFHhCgDxIgHZQuK53xsZ6UT9z0xcPztt6kqf1lVlgMI2bn
BAoYy1Pb6J8tygBGBwk3ysgGigGjfzhJ32IDqRfiXQXJLlH2+FhBDzStSAN6q4m9
F7X70Uq5ysC48JFC76OaFvv9JzW+RQ2pKgv/JC50ffZtHjsFMJ/nAzlbizSe00ku
tDl7EPuoYVqrP1JlADBnT1ctLRNUblYQXKbgKEgK++ELJT9XCWKrYtDzKuaIqxtI
WHK5726m3P4O1jgGAV3x8gAsaYLNwHXzGE++NvyULACyRSLwqaSy3WHgioInBH1e
gnrVlMMDcIApil3D7QkyiOJ/ooL78mnuktMenu8HtYYO6xkM289ks6uZU+KHl3KK
dgX9n0ZI+AuEjd3McjAhewUbgtgohe8tAL9ssoV9issBOUF0Jvff0y8g36faYbqE
SLp7JcudPl31yxEvtxmFj3iEIIuAOPmtCqCe5gphYDvDZHBxLzG/uQJpwsfoShFE
fwmONqt/zwvU2PYoCHv19V8lQ6m/haIJzgiWV63P2h5ksbYMOvgbDhtdS4O3pwzE
3A2/oJb6oNPtWrgRqpmCB4hPRSJ0GzLTy0ZWNhBwzXBxY6vZ5UCsXIlO/Yf0DFGG
9nPKJZy3YZsHrE+OPMsbuqWq4fGs6A57YAsFNfngRYsnxqxNpt6wM71ZtOpNeakv
r68SMnne9dFKKAWbesrA6sXBGJGOhLtbvHZH5l2ziWj6P1/PynQFTcOdz7UB7QC7
WJSx+FKOlzkkXJzUjzCnRK/X2lPHFoqT3bdnHD2p5PoMpr9Y3vwlUyJmx0UdZjLJ
TAs6KxUnmU/yOeIGPDyk/z9aIfQipnRVNGte3L7wfbrQGy+jG/YfCTtbzyNyVX8v
WvrukWiBcYKt9i49vW9cOcx/H8x9AsTrZgfveb4XCFKk25DaoqNfQ+CMLldCJBBI
w7rO7HnkAPiqgfAcxzif+EgrAtSx34oxEe10Vou5Xgsk6PICjzwSoGU7XxfUfJeG
nHabIG26mRPSJHAswOVIS9TzumrBY+MfSjHUJCTU99yih0E8S+lVgJj9xv6Q1n2a
NrQ45n9aYswnXdxJbJ1aEC4M56ZJRqh/GmDmAAbxKvacwwe112Kjq+skdUbNJ+2O
K37y3A7cDGEyOIyX9CqvODJmDU9s7bmkTICbA7TlnZqhgIs/OmyKZjgdUhTLMXGH
WUAFyKRco9N8CpxA/bmKM++6o5qvaiewTLoCER5g360Cxmp7s6M6OzsdXItciCJO
qnvrLfXPZflzHuvY51BGgR1ZyBikKAFvcB1wIwfJw0IGuMIWTTNx6s1oE2CYWH4Y
tTadlqiHbfNce6XkpJoKOTT2pCNRQqo+dNZiG8LT5e8fdto1mTG+gwbLML/kVNLJ
iylsZ/837mjPW4lKTjfeuN45HT4hlrXA0I4x0uDTCmcL6+cgoagfrKJsr4ItClrN
k5fZSEiUsOi84FfaPI56/o2h12GFg3AvMjyV6yx2SPjoMDbreX5AMpMfpNOZbfID
k4oPgdSZeeEbCJ/zMLODW7WzY7EnqlZ+HHkRbVGlFEakyCEwaAGLNSmFPBVgijr4
h+WU8P3VA+fUrVa2EUjw648J6UuZBQen3zEk5MGm3HFcamVaJ8XzeNV3JLi2Vry3
Oe1xWt9G7Zm2AU6K4U+vvZNtJlvxJ6yHu+acuC6lclV34EWdRth2hC87ZEp/eeZW
7Al75fmUii519hikXy2zWVPYHWHEMLbHcmtvfwb1vYdu2oWvh8jrEMUH7cgMH+o1
5Dr6LF6iqYHJJoX3fCmopHYYAoOKprlmFBDM1IZqX6ma0U89H4EtoFBe6SpV15Qm
rHeNVgGbgNLqQFOOZt5mqrF7X8OlEePwIl9SoGC0ALGkh4iCySxhFvCUU6GtORmK
6WNXWNgvrjFWoLyx1E0YhfMYNCzgEVCz4jZoc4fkW9xs/AglDhAVFIWaKcvyRAsA
/+UIhSnmPV/92IXduwnhMNQ8jZQHWIPK3unGGkUZQ4GgjHNF/aX1nT+gbnTzZuN7
J2nbVaAMx2zfmj6ZAnO52msX0282Q2DuorObT0NaSIskUVnWbtsmvpoT3d/9jATf
axOIt/Aas0zdWFAOchOckg0BeQAZoQ9kxUY5xmrTl3hv4/sry8Wmj8eNemZ83A5N
JHl0DPWC4yWMGHZ7ie9/uk7Xrj23FPHPPMozp6EzRZc+GJm5rKqDQUnazmI8x19X
BotGe13qH7MjiDLlqCvAkp+MY6sDT6y/uyHbpCwmAV3mjpxrwLYe+2Sl4d9yhHa6
DAbDRrQvPHuhHXRriGOBGJGKLLu1bG/NzDXhSi/kop9K/wdLm+pNqZXsZ+rzrEsZ
HXWnXb8LlptPsWlbHfgXy0uxT9ZKjoADHi7dRfs4SqMs0d8NmCNK0KY5NRJyCLQY
na3sM2MvtsFHgnhktD/9y7dG9eX9N3Ud/DA3wdsTdu0R6pC9D4AOrVjlE4ikYbA8
LVEQgoI6w4EcGADbydOf9BqX3Fe7mUvvuNFAUkqRqn272wsXfBynpsBvZ+M/7ibt
JhygIk0xBpmMOgUBooxEh9bKVcMUoT76uLqdzuzSQKOFJLsYrjwynO1FIlwO/4jO
bv2OJ4saje9pfzi7L/y7nOFr6nYxKWtzvxFdp1dc6PrBNiwL6eKRdXCkxHwxaKvn
TVQ+x7OUNK9HpTiYqtY5ohzuLNZSlPBmQDq2mM8aQCH+4zEaGvJhEJFo7MIfcFgD
OSgJEDZtihsEMhiD5Nq0elGeViJeS7CKxqsdqZu54lcHCb/bGB+0izf+MP7TiNrc
+xEdaNJg5kN0F3BH+m75vZDcFWXsksVdRyWzL4stXbMD3HHztPe6qvbmC2Gtc/qB
Fu93Nk3UbUHGSzZLXQi4QoXYN/QWEFWdH76FnHUrTP6tp/9UcbI9uRTl9pQY6by9
NYBHtQGhSY0wckFM8JvSAn2W3bByOX0W8NPyi1DmCv6X3ZF772tWFA3p++80AXLn
6mClD6mF2Z3jgl8UxYWZGsyNYW4qb6Ucdyo3oRnqFbY2+NnafbxkSsxCKuqPsI7z
Z/i0fePCVIcOYIZf9QBus/toOj7II3dqsubc+oiGKFR5HJg2nrakeXea3wco8zH2
nLDAOv53et/zfTYoNE42fwt+8ltBTwPrPyGb9ZfIhjJ4al6GuNU5hlQU8Ff6qemW
3lSSRdVt46Ou4ukHkcryQZl7a7e32Y+3OricSKFFRQ+ZktveQXeCznJHs72GAQ7R
IupoDv4IkO+Ljlu7kE9P3I/z4HD0e/vwYaHFY1+5revuUWVfe6BBn5T7pK+I9YiP
pmFLXPJhb7aP5RoFNkVSbmLuSN73rjbUnKfy7oTMQ3APh4vPPp1hAHkLTgl5nrMj
2MBjH2z7MN3S967wzSLv/MBlaE8/yRvc+gCkcNlFj2c/Mpv7Ky/4MXEqMZWpqSzE
Xg7Phz5ZUNxI6XKFbzOfnh4lgB5bT3oyoNW/wzIIXRtgmL0HXl8MU9Ztz3SmuWTu
Q6S+W4lIg2y4GpAw9agW5ch6G2ZWqVjti3x2cLTk5soFiiqTGbP1woelrC6pJI/Q
+d7b8qh7aGNGutaqOFEAbdunGknEQEvAAodr6xM6MC/Cnsrpwlsg03QMewUDGuAK
fKVxCOTGso2owyX2GFZSCG8eZXpZWpYiRn64iQebNS20JR2dJaMVPvcgWsNIEpc9
GoALfefQOgDAz+zpLJTOlZ1SdIbGaFFug1GFR0TLV276Y8XlAYdVl40lhyEqlwO6
/zJTYj4qOg5a6It8tENEn4b/RluokTCibohwl5YhnYN+X+IlyNk/ygnmZQc15G6w
98lXorWVve5NBJNvTvGQ7JSR+VGEx+HGl6H7jbzQFGfasT4ShJgzF+rXXu9VRq1K
zD8jSKkjFJwBFfLYXWMTK7dgtLDCITLuWitVsn/tEJ4xEQbNr1+pMm6CKWPA1LIJ
ugdixpXZoi0M3DEAyCUZN5pZufZqWkOoOKU+9Uf/aG9DmABZNHG2i+OWQ81L350T
Nk6J5X3+4f/FZwMS6xzb1vuA6iDdMbi6WlZLMi8gko3QJ4/idEMpMuUXbANYo/w0
TQNayHN1KEGnPYdawaZ8F+AxpeiN/P/J1801gzqmUzCXRJHLZ50OcH+6xyjkZpTu
8u8iRBiTyGpEcfsjT3jRz3z7NQrbwzCN3pvH7cbwLsoiZ/M5knFKiPBsbvF+ZJtC
0JP1bdHMn5sCl+Wl1HQk6Kx7HLlTMSucSzvuvbTo3wuBj8PiyaNSFGt4ernqTA/T
NJDmxVioF46grxOdGKd5SmCkFJsN4s1SaIicnjq5Bl5mkQ2FVNhzJvD4IA3Vlufv
GG4BwM4Plgw+Mhr8Z9bCX8j8GpikA+Uwes92pQ2CNXaOPd4eYxhPCD0j3Z1zVqIz
KnvsxsncZjFvf/QPQbKwJf1G6frjvSsXX7nSMi2U3Y85MSJvd0KZidgcs6Elmo9B
irvQ4P/zoJ/aILPqFxnpXJ84el9z5g+aAK6r3iaQKk6b3UAPeWLFeqj6txuyw+bT
qzoVRTVVQwoA8dEdytCXXx5723RkD8tU1lBM+R4m7j+03Ol6ygKj+2Z+5v7QdNrj
p4uXhItlJfMa83BzZHZxdwKejHzxoTcxLSMbUiduBFybKqpYkYR7qUT57dcd4fiy
wVoomeiM/6RDLnk2TplCj3k5n2DRpQ2OiPCD3uwKmguzhWyj/mRUq4fm/JWI0bRg
t0VdHUM01gfwTlunu36jUkR8fhtFJLAVK+T5r2yqOzhIvVrX21/NrKwxfpq5UCRW
VVhIyeLCzsrtTjuF2pwp7VUSyLSEoHlkt+aaJ5jBVygMe8w6vlgIOpbBcmNc9xKK
ZMYPPx2oxskX4aYRunKPjDDCy4jSbn9DB+eSyu6lAwAK7eTqhxzY3iDk4NT2kQdR
w2gNUeecvVnqbTSGVFxGEfMkqefgpWf5c4LdtHu/+CUqAdVWU/Cju1S6QYqqa2LR
W9y6BxXlZtsn1rXXsjHvV+5pjXKZDEKTwNxGa9WRk2eX+gL7PHhyi8M5ZM3I2X//
ErGcZHTgtenQ/NkhXYsYq1m+WNO1CV0e0gfeSWrR0HeTP+Ml1neiix7YvV8rIEu3
CZLNV7o+VP526I+F5We5mdJzSmyq5d0Csfz11fxtPdgeNz77gwhRBAaH4xsotm3E
7YxIpDAJPq8JRklcQwcUmNiKdfzZdmc9jruD2jP9wiTmnsbKrziXWK6O2XRcSwFD
60qBHah7j7KXBH8vii1hyKBmcchEML2cxgFVSUPl3mz82uiJlIb7SFyuxbo5FzCS
dK3cKc4MgaJ6AnscSrZ5fEfJLmlol2WdvAeCNOTL35iuq+dfiklQF9f27x12lBqZ
zCCQwk8NCX9pgkrLqwvVGV3JNieYHYrE2hgKB4cVXljGiyGUbjQ6jTD6GU85tqqY
GN6QRG1Jdc3+I5fyyS4Fq9R4jYRuUnHx+B7ImKnlac1yXl7U4OzyptirHaJdbns+
wvR1yZ5mOKuCcnSCbZbosF3kDqbVGCZiwVK06gpOM7sqaBi7jths/LZ4iOeu94JT
UPaiKaOrLeY8CfodeCPzVNmJxlwRXPfVsvLnCuoReabXSP2bt/yO+2IP1mWIIYRP
5UTOHV3OfFuwDyyDnoJqYzSwtgjph/w2Jy3FptZYrgj4ueKw4uWDmGGbTKiply8f
8LYeB6y6rMbVaxjMfMGSyJxMC21Add1Ibr2/5sep/gR5y3xZjbC4y12Z8GIKusXO
YW+c8oZ47doeJ6rRdJRDTQr2G4aoKcGJ15r2YMuOxKl9rmazdjSvBjz2U/sTaFcf
INvqoPcrX88R7vOcsLaYpE7m+BSpno6xjgb8nMMSkMJjUbZcl/rYctVSHfbereqi
SWA18TcAo5gyTrmLPq/JJi5kC6EvX9hDXPAsv1CDOXRs4ZiFJ7Dr5DiS4eZUkeQB
0k60dO1GhzRXNH+0Rp9HQ59etR+4H1xuXSaqMbMyvi6tvwZnDDNqKO9t9NSaDNqM
u4WBPghRdMbrKfNj2mbIxD0qdmpqy52RUoj6j5nQ455PPtk1IT6a96uU2Hd9X3zU
Kdtgk/9cdfpkzuJVtdnf8b6DdCLPhZKpupvav23iVVnKKEhpLuVagRMk3KfpIxCe
4ota5cpeirMNE9LEUbEnWUdMk2b/+H8lBE1iZrGoyYyuoYhQYYHgtOHIiYpkk5Kn
WOdAvy23IHZAoJM/3YAAaKwJhfXlS7Dal5SBZRwR5tAHnDAInfvgqjWfr2svzqYK
nO8qQS80OsX6WxSnTzT5+RDW5YVa/yemFDWzT2St6VZOB6KoWY+1xmJa41wVunW5
Z0lJaRGtogl35VkKxw6AQ71uQe0/p40obh2WFO7D6o22jfv8PtiNmoKawaZO+d8k
VmK5v9zNlbIrrqXnXWHR1TNG7bzo8n42gQKcb+ELk51znTXMZIupqUBxz/kSYycj
bJmUaJGNB19sIoeRquc6RotCtAIQYKu7ElTTa5XrUHKPFMu1FDjF/zds5K+ntFL3
jeo5JVPJqhKErvWpq1gaVwtoIabueCv5+HVd6EkSjzhRIrTRyXHI3gtIKvE6fbTM
BpW9JV/cscWoScM42aESHWK0dOv29h7KCA8HCVhTbnncIrnmPeWT4f1DgOqoyaNW
PzvdvYWfUScFi8ndqNK/zdnZiZ1Zg/eMuKhpsDvo9COXTf0UrllOYExKLkUjBC+t
SD+yj2OM8EWsxGgWcSCMW5Uh6+1BHxCJNk4VxwruXxkAoCBZFgw+YuIigWRHPhGF
EkHiaLfD30JZQcPPo5MoeoBJg6hq0G3WG8EsGonahBSvjnQmCmQFfemBcmPQDdzJ
U+I0evbcYgczLHdo7sq/IvltjdOD0m4w78MGyjgfFigUBgex9WTO4KMxDS3wVnJI
tarEQRLQlVBJrkgwnc3V0msG7Y/jmVfsx8BfQb4hGuFw8wcw86/8AIL4QQWU7UT3
1Z2UV8in3QpAIERrMvytQkEf9UznAkYzt/j5vqmJgPoBFzGlnoExnLn1Q/9F31Ig
Y8TiRTjhKi+k+oedvtJudAlLnmrYh0sBrWp0IFeCgKJJq1h8CDrEKgBO4y6cBvaE
CoTlNfZm585TUt5/SiaTa5GLaC4QJYJFDm6eaqlRfYS3G8B4ycBEGCsYGeLo1GtU
/lZrDwD8SHjZpROcLK/HiYHNpRLehvSOnYVn1gDjMfG2/e/BRKY6WRnBtvCvn8fH
eqBWcRgncIwHcC1VnXZYioBV7HkIaZ7z63N8AAS9LCUo3ArqWudj3EVCBpwsmZvn
e47d1FgUugz0iS+OdUcH49zbXWkwoYR2sMp4v6jtgS/9vaTZGKZ4ljwqr+YOb5sY
K/PCsbPAl9IiOxR/+SlXkcyslYYLGUCajUIgMTISA1i4eoebs/uDT9q6xghwIvRG
dEzeSKGagb0rEujlWUzmYbplo2h6Fcdg341F9Das5g6LbLw8DYF32ZJBTbheeHzu
h+2dmazezW+oDa2krqzJ0vFgf47fuXgzKltTas4O55T1JH6hejIXXrjnHlIESlRo
FkhWrnPvqnhBhpZMn7HVCphPkYZ7ubEQlzC6X29PxHh8W7VzpFTO6Gw1FMbxa27w
XRIdwnsYwoJMvY1wq6INM6RqcWwZizAYpaAaSukg2xKBG/KtOMVyqm7/q1TN7OcA
V45BDrdsXw/RoK9fQsKH1k/gmu5bN652Uz2s+SovmxkUHLjMmSNxGcs/2ls1Tblm
YdCaAC/qTDiOPq+Chm2tchgIurhQ7HyfPTeE/zgtlbZQGPRiB0u1xVWddCRKbZv0
DfoBs07LntM4wluh2p16XvqNI11SXzGVXFvUerVBxqMn6YpH2RbCHEl0t7FdTYcM
Om3XMAKlD4q3vycYjxj9iP1VaQq6x51JA4fHbIoXZvVoKIN2JCam9Kj0opxNtscI
t/c99An7XoSz6GADbPFpdb+qP35oK5BM2RpDCk87BKJhywtPrffimXxGanyswfCa
+zYuSj0PEkFrJWwIWnHsxG5xYRvn6JtcGFCXt9HttttsMiHLaVs+Dr+KljLGxy2r
KdOiGV+tqkj9xxFZtpR3jGp8kbPYXmMv0JS64oWzHubzsyAayXDfg25gZHQsEHca
FrDqGcqXUu8LuA/PJ2nlOfixp4e7f0h40LpeBnYeM+92e25t2+b5bqhf3XAIvTCs
Tk4LNMEN/cxFojpgUtJbXVhUlDuc365/tNRkYRo4XYgLbbKWkz5Gyy6vQCSTsDL+
5QpPNqZJV7801qip9qEylOtOEsd82LpwXpfRg8eUnBcZYU72rLIcJ43qqzEq298Y
ZV+2u/PU0YogLRinrAmeOMvN1S1sASMKoSzo/8/1jezlkqiedvrPB9he1Ed4UcRL
tM1+oNkfCr5XtBfp0a7+3Yz8XYrOWa3jbwMKx8j0NoZiR56Uj9iCf7k3nzH9V0GN
CytLM6Tf8O9go65a0cHYUZTXsohu9l8RZdclU+duuawZyTG62HmCduz4ZgCp5Yc0
mVEBUN3EnCVGa6GTof/5DO5xQHIEMiIJ5V0MKXnh8T0StPbHej2yu8X2W29KoqWC
+mx5lYposGxYCSe7R+rv4+DcNEMSEY3BpVKlh3IlkJ6wCxtxnN2Iu6OeVHMGoNx+
tH/KOOOqdK/hvy342qaejw48MdsLovqcyrFngRPTpk/QXzXdFIBeT6ClHAUbT+YG
9TEKev2+nyBGNlM195RyDUG/4WyBAHLzinTh8Sa6pwjY3E+eqYyb6J4kMm1Teyv7
2irAR86MACH/Jqc9qyj64eiYaJ1weWGlZgNSPigvEcV8IzFgXdtpa6moXAdZyFYI
u7UFsh/cVGoKeFg3c/1JQePW4Ta4p7BdILVjPUVrrqMded2SGakZJoGlBs+j4I9I
p2f/7Lc930SGh1nUa9h7cXnMjhWV7eKj+0J9xVXD2sMq5dBO9VuyWO/jQD8ukFGL
TVrDqakkZidzwGgBcS+G6PRn+CACwM9nOrme2zDkMZNhumBi5emkmdyLVuF2xEhx
RxX5HSwlFoserDmjpZdyEpqwhd4coq00rO5hHegRWflEK74nVmltWhObFulIKxzz
Mxyp17HfIkRCJu7lReQNov7p8nMdioI/7w51t4bD2alTQYUlFQJyAsP69MP0dtPB
KFd2HOZXLzfA//mPdKUFt5+qOmMXvF/n3m9dwDBm5YPdRzN+XCEKeVmGfoAVNgrE
pVLleKll3We5S34gwm9fsqmSSkdM41gsZ85y7dIPk8sQPzZNEJqeFJl8l2utrQ/R
aH+Ji03fLYveKhrh6EVU9hEwWJ1A41a8UQ13mMCErSOn3PdNywZI7oOxld1/tge/
APID68CV6eVsZ4d62uRQlA2qY2zFgJtvPMkI2OWUWmsIF7UDuZbaePQ5KLiKQ4oJ
Owk0LO8W34LMTvyTIX+sXMW+nYbJKwZTIuqvF5SveSVC43C5HpAQP0Jyu4tPvavZ
/zMYaxOYZXlb365Yucx8gy0666s/02UQ0j2LLwH73Bx/+dUKmGLp0AE/wqg7zcXg
3IG9Ksu3oKo2dezryjiP8cYcVIuzy2BJFYN2RCnDo0Eifbk3fmityeRKSR50BQIq
wOTxf/UvxEGkAAgBEhPyFR9RI+HjDOY3Mml9xEJkftPbyZ1GUkvt0mSfxxbC54SC
vDQD/gKzwUW/pXufbBxAv6O2DhxbvCWKGAUiyOZ769LE6SEffVDL339cvFHClPVs
Sr1KyIKaljH6+qEkfGlezZfxMbNksKwB4IyJz4Mo52qJH2xem2pUuGt3pzYhMIRh
VifgfzkPW+FGssqFMSohjOo4F+c2DW7C/Ka+LFYvpVeUEh583vQbveT2czu/eY7D
6EpjR3eT74/CCaaWTFcfMZLdArN3kEHzNpMFd1Qf669EkkeoFd37o8SnHyoO05mt
wI8Osu1SyxqN/bPFK/1CPMgYBS7yUKUxdAxai9Xz3hRp928tcYnVcPEGA2eiofGc
qQrqrBO+XTvbblyrPdAS3SViC7nXJbVJ+Gcd9ktXiUXxa0OgLlQaUIfOdNaJew0v
OjN9Hv4327y8DeZgKwyGRnLGZV142atFDfev8xfYE7revWjkvTMalaCRemK9nbDg
jZqCl6CicExysvVsT5Nj15TPUQmP0kSSFi8+e6VnKo7NdZbtgjm6bvVhUuHe/O79
Eb9pypkx7AHevvcwcvI+qMs4cGW/tS3jEpt3sG+125dbDRwfd8UWUkVG/hNaPLFi
7oWyQ82vz9LpfCARZ6MasEGOJEwfAp/iZP/kCiyesmDK/kgdV5RH+78V5y7PcimJ
/snl+aY8nhYCzDZAhMFY0UuJELtKAUnR/PCnL7uV5iztJnCI8d55vCBdCouNP2dn
0X9DohBSaBvZ6DLjJz5RdbT0VwGGnROCcNqM9g57GmS65PhGACD2AeIFmXUgt/31
L2BR/3dlQJwLaavNeRtQExi0+IhbRIk2SzZCq9tYqNTvdEmUbhELU86VZ+UwOgqz
hSj3Gd7INhGFYkw1hK/0H5IXPR6M71kJj2zWLdTY/J4JJQxikQNh4jJ8KmQoHHkf
U8lqn+P+U+LC++HN6IDwSROWxs+h1eoNDJnTFXbLb+EleTfQn9TqsoUhz+FciSqL
hy1MoC9AZVoaATYcbPyZKwgXeCcxYAO0sXaHZtW8D4uphNcWiwsAkvYjVRzQ9Nt/
q1dvII7eTzv4XRS+9C02SqCaEEstECSVpb42pqw+rJPuNzuGUwRM87u0+rOWVnPU
o+TLkTkhGaD4N/EXVBdRz90/5Twhw4A1PwreZOrw4eQ5AzqF9AqHaW5420fSgSJy
3k6PLT14xHbG1+YoBFohf5tzlNCuzNbMI20rC2btvjySD/y0BphwRVjEMW2hpUOe
87Sl8EDoBmK8n2cSXedg3IUvvhM1CossxYMANTqnFySBAgJg6CvJnnfmtxK/47SP
qOHEEGZ/kLp74SlySlB/kde+mrIB+x7rm9XNJM7mq7E9ik6ApZgsAV27vlMwkiOF
HDkDSUB+0ezCR1GXmr0N5pSUiTAWnH+rsbOkN69TvR13+m27oGM4VLXSXSSmrEDm
SHV+uldoKqstIJFw5yjZovSDrawbMfkL/dy8+k1oPLL9NqsNEi0dOfNFMsQx89on
vAAb6l38W4hnPIfcjzZ+7rUHe1Cc6d4VdE0CYealYwnj0ecZ4UQmmF/PjrwPz4ZQ
cdzyPnG6PQcWPo5Ju2HXnRnzhyLtULwIhg9CbYE8ke4XW5dZRHMeXl/jHKaFLuoT
IOmkAdO5BU9Vu5NjryUoSuGz7UWhPqMXgIivAjQJaSVC4LQwM/bjRMVWcS8JJU0A
8glC/RvsNeCwqAlDqPSepJ/UB7CacSdlW3LzTEHNoqzwD9sYCZsxRRpybs7k29np
XsvY2VwjJ98w50JFVgjqzI3p3/MfTWG92j2+Win+0vMJuJuAXBxJH+cB4oXRsxfc
9+yYWCLBq8cYNqEwkoPTUJ6H8Z7OLrjVnMkmNHuKu6+d2DU3duB5vWs5neddG4Vr
SwMwNaj+2F6H/vtFfkoMhDLLFBC/DDBluzFtYJ/KMYoGE7MwnNsyVc9E3+SsNToD
OopI42Zd9f3QUvojJ+vKj7P2CbhAobQphit6MCwXM/+zbSuLIGxUtGHpSWx78Pr7
kSsGRq0RvQYb/rHlb11vbEGBa5zIIkNJaIF8AfE1KMKZNkl1nx18QOWP9hcj8Lml
RGs10AqhWe4jn4clAbSQvCD2DfCJLc7IfR+tEb2J6f22FpDfL2z+jCI4nVLYLgfW
1KOIADOnnWmCjzOnbFmx8KciZ3pc8vPTlq6As4mNOc0lV/VCejYX0McTmT30YLhk
2CYpAT4Pgmw0dD3DHJVGfOo3CzimK7qPh4CQKQk/AX2g9k5PgXA/LaChL9oCi8j4
Z7ptKHzfPOybhDEuP3SZfdse7f0LZT+/Iw5by8rT/+gODF4Di0IcMVrIPxfhYoqL
e6/9tJc2GGZj4VRzqzT9uH9LdTJWZgrVs20yEbdwil2ZeERYDBFR2e0CVFW2EJjS
+7EI5458VnMgSXVZoc+0Ol07cHcgGFY785/lU8PKtXFxHfif3BAVmm6ovihAsv5W
bvwJTQzW5UXVQp2gidxj2CQRBQiNMOGYEYRfZBKRLIsB+7b4jHWW2AyC0GbgdKVm
+0md0l/zmmUjRSvBqJsEWyXcQx+0gCP3XalW0iyqLzR1WkwGenOZbS9GmyHo6ajP
hVDkXDGTzdJ9T10Nk4Y0Efu9GAWSydQhAriYEW4Jdxiyc/L+BeUKgapc7m0IPmwg
1RBuCYtMWq5yIPgaWjUlxwScYx1OzxvAzgIsqfvGcEctzGdMVyThnv1CKOdbAyJJ
RU0aDMa85BnKnqIdxmBNgg2oGueMo9QI+UKsJhHqov/ZaiI5S98YkOFjzSd2EBag
dWixACW865i0JbqBg2qX90++CMm/NR7gu/Es3bvRixWdLZ52WXKwm+6GJ04ObKxz
KUuN5rS4lRQS9nmFv8LyXNoKJX1qMFJoBLCjntNIFaJNUp0FKVPJRiCfyzj3+8wZ
RBW68rEC31DtjB0yKjIz3ATXO7ddfd4E/NfNvusevRVPfKcfSClD620c/IKxpWop
DGBg/UyBRGwaVonoyLdq+z+fM2IlKj61mkIEIrQ++o6h56mLDmV04s7oRzqhsYk/
fm92i1gcZiQ7AJPFQHZIPT0OIcafb5R1IYJDwALB+hhpPgMobS3i47LZCeGjbd0V
uwUguhkNU51gJOzWVnyOCPBIpVBV1B0NpPO/4yWAYF7tt/KJFwdlAKAY/mHf8Lsd
zDYuOwV2kpf0f590XIzMkeR7w/s+0ra6AH0g+UFw04z63q8zgnw4H8tEeA2ciMfn
jZJonkOfmJGluvWHaZ3NnStzB04SQ0/UPSiGVVZoZ/wGneJnp3uIcjJP98H9RzED
3tQI9KhZm7P4lPHdNGWoVl118a699S928oACunlWvkkdJd9WwpJmQgyH38HvWHVc
mixqAGCnKQwK9yZvcEeLsRFXPik258/4pIzEG9emDuT7FlaRttm8e/n+nf9D9XBe
p9+RV3LLQYf+gN/W696tg0stOf/dVJ84F+A/YInUo7E+Foy7xHi3SqvzDhwJEtGb
/JSGIChvEXVcKSsEM0h6xfVo5yGguQ/tmiMTAL+zP1nrHhwyVIUWgctuxEr2PtNJ
7OVief6Kf6kWyGj9A5FcHtiuApxxkzX4Xa+nRQRlN0o16UskCKXKIdNOYInK7E33
emtkolqiVeHkMVPpGyYztqa3gohOSvXKQvDX8ti+C0gH/rnVEJSSKd71qzfdWI0i
+8JCnl+AK4elGUuES7Hb9FI+uIpLQOMN7QOkOET2hG+1HljY9fFP/1UTqYKUyPfz
Q2atRnLEAkOOUscKCOayCPqjQa1P6sF1TqJrbymCjSuFcfMlTXb8DPj+QYxOwo7c
CVt4+B7zuclb+N61nEdmQ2tzhkXtJ2VI0ZfVKj+PMAO5zb1WfHt2qwVnC1GEsHTZ
odxex8WSgCzcfxbMuTnUFpSojUzP2+6rGBr/8t3bWIAE5MOU2Nx1cw5ulDeCk3LX
8I4ocqwBUtptU3jHWfRuWkMMKwDFccTe+g4MTHZ0viCykbR5wribrhRhkpTeu2E7
+I7bTU+Eh7s3WutHyJVNKGormBJ8KfgLrWHtMNHpx/2rS8Svk1hU8OFyAosrHWDM
b8eClrXX1DXwUVnD3Bo3f0oNPOk01yrm1XYPNoLIyrBjK4SGL5WhYQYtUDqrBDD2
4S1GVGGilkaW6NfSI1gaVabNLKkF3kNIsahuvmDI/qpPikniQZEb8bMNvLfYM73Q
QypqNe2uL/UlUSAXEr4fqV64mK1nAFjORyvQQvVu4MK7OZcmyLkfmsDV6pBl3S1J
6Lp4q1P+3OEtumu7r7t/VVmLimbKRlThnQjzpVWlLJtfA1SBj4vNVyIRygl+9aq7
60bWK+R5FQYqnQmI8HZAYoqq3EInVeCl8KPALENTDSPudumUrZh0be4odyh72Sr0
3Le+i6tX9XsX4Pe4llVuQsswp4T1QX5aDEuBEKHIljzN87TPKxmRH6J/KCe6kYFJ
wfWrdHY8NZ5fywd5lvkVSOCI5xrcPdchJGKuM/HW48VKmjransUwG8YBDIMGJe+t
xWOogXo8E1TVAj7YmQioYmyAbOxPnR5Q1lF2fAdfHMIXmS/BZX0z4JK475yndEO0
ePaPWgOCeyyoYXxv9gjQEfnUwreLYjDUOb1jbGuxvLXw/KJ/Cif+weHmybk9FqHK
8/ZNfHvhO0iwRHKvXFP5qudyMcE9lLSni3FG0LDcff0m2A7TkLS9XbMUf6lnfzZW
QyjhQGZazpyg0EG2rWwYrEZHQhvMpZ797PzwkrScIlDNMP/FV2RPcTarWUaKgIUp
DWaLlVxl5UIb7mOBP3rvSo02rCNgG7uOy5v81sjfs41OhxDw4MxB33UdrkmuZkUy
JboxkIy7tU7hG+7rY9HDZucvFCQwl1xoWb2PwNg80ELZvJZuY9oo93cfKQXK2fnL
LcEUxwKFZ7xTegddP9FZnxaTRfdxYlOin5kNN3sHMCw/0m91lsxCDB4OOYDI/VL+
oJBgOvAe5O1F3g5fQjzNiOW1A5fQqqryuIWx1o1shzPOl0TNllbUUHl/4Hjtcngg
HlhIHcJASOUGGOIJcXraezpfA3QD+GQ9TgpDpRQJkS18YlHwqlT3811CR+V/Fl4k
LEOklJMQ3MmtX86pwBkB0Riu6sSiyYJGA1g2q5MtbDezAbe52R6dUby0OMbmUXGN
s7Bp0671zP2lXSy/uVhgwpULdQiWxjruNYC28epq+2P/9x0G6jfu/lRsszcNQeMf
Ahxgtiql3UsHct5Huk0lHtjqGC29tPJSXUGCjAU/iSRxkC0gg+j5YG1dksTOqhao
jcNj0M4hHxVXz4B7j1/mKNZep4l4IRNcbLW+pf3wz3sPSXtvDmbZzDnEq+ipAY9L
4dfbgTck0mtVg6P+I+1mDuvg0wT9GgE4veepj+l8LgvO98fUDM0Bw7d/r0KtLTbP
YNFP/xtXiklpE5k6DhzaF73k8GSxjPqqyhr0jJSs1wqNFw9SffCUnllSigiVN28J
fqpseUIZtxt5zaq6GCaSdhmguO1+35HhDqgi0rpznSN1PAyrwn4HgPqtEvp/6cOf
rL3dYPi67+XmiE+crTTxNbBnEOC0Iq6bCbxpzPu5uelZLuU1mZHX7EU7i4ndToC7
zUJQzuCyisx1awyfjsXcIDvQn1dGJW5bDUORmT7GoBw0PyOEmqdBb/EWI9l1Gkk8
G7/HxQ4HIL/SR7WJD5JckNb9+vUBkFGJFHHj9zhoT40cnLVbqc+1xzoRLt3jLwnr
J+SfJOGoGmUrIEKQoYNH8LuV9sG9DvWWMLuzmAK40JPEmD2FqLwBmsrARsfBGvsj
8MmtNjyWb916/NFdlamXIVF8V3LYDHoXz/aWPcMzW+yy+k5kw/KKZOYXxJEXjQtW
ddNR+voO85PQ1e3c9nqZwIIew7zZuPRpn+DIcWTte0uYN3nGLrr+8uRbayIfPNrq
k/8PqZxeAm+UAVaBlE972ocj4e9wk94MZTMNh92nCjxEJONjAjf5bIAsKc/IFCcc
zbeWuwE87/YmbekcV2RXOvXwAr75aSfmf5lBvU4L9YZwmyAj7oM8UvNRLnB1BO37
2aeciRBnGSBeGtf4EQVBn+vLttSR+3bEUG/aCSsK86oIlE/mimipEIwF7Ld8a31y
4eZaci6OSjl0C+00TB4/lC2HrxT4cWkDH9+MrVRP10/LaaWdBiHdrBYTdsNGvYKu
woc/2qIU1R6/3AHYCjklMRLmmflaoXnGjrOdeAPyf4ZCXINj6CiSN/8RsEisQRqo
vH3huJezpoCoaWSs8Yfd4SmzWamp3rsew8PIljt52qoyEKrLx96Dp3fRLngHYM7N
dIAOF/ZS2S8mqSZBSxpn6fdj3cXO8QbB/KL9slK3gwU7ZtSSLEp7f6KN+lrzYQtV
iksrF0FSzclfZc+ON7RYJRX2gWjEsp96pi+QT1vcDVojfQedRn5Nfsu4mDrvXHs5
5cabV+Jf6jNZIFrZh0HMN0FMNNS/lCWzqf5/iOu7zeS0Ymt71x+Ts49o84dIzVJH
034hmboGamfDoFkg/vMiHhVwoT6vM/+s8472mOrJX9pZ+YYrmv3YZC50ez5CJyaI
jc5A8ptiOk0rGGmSJCSba5VasVKwnC6L5PFl0kor/FAlW+EJCyqRJTD7D3N6W6Ua
37ymDQZIGsXvJwdubTFkZwN092TMCVToQHVMRL+ByE66V1chod2i15lOAYOhe5DV
lGcuBvA7yRwhUgsG4P9wfVJQrM66ZQJvqOnIdj1XFi0sgssW4tJbm8WdplHfYK35
Ehxy/JewPeS1FwGR4yTSvUbcc9H6RiWiajrI04k0br1z4GcDuv/2FdfIx+jgcQ5W
IeLzO7tpiMJ7cuu6Sf7A22LhJJqk9tZjrOU8p8OYA0VHtfRanevvsBc8tCgmynLB
BBTvHrwLTiGQPGsV1i8ls3NhYlmpFMRlTmYTHBA97qpan1uxRiMQ8g+4gbyntU7s
uARVIg2hH7sm+mwq3zpHQ2xJQkUxwsx9BH1izWXCmdpQFVzvSdRnywVp7w2GKFIg
OW04FIiMibt+vxQM7RnYz4VioIpm8+Xct4k5Mui3esB2yKUzuGDJv7bGpuZQxkkR
M0w2hcMHsb+nHiB2dPmGlm2TBmgN1SCA1rgW/pp1i/K/CX852rDQYAu8HytF9UKI
A1ob8kkFwAEzSI3diDUGW66BY+paw8H+nnO8Nv3l3UdOcGvpxl4QsLna8jS1ADt4
0Gnzkhd1EpYre6D9rDTPO2WfSPCWSNDZ2nyx9xDSVtGF4iX+VW6eXuiCn0VECo26
37JXS3yrIfWk2IKRBjJetT/PQdVlCtvYBP2XnyE0ekzfRyEcbsNuJJLwKciRRdKd
6oNHLDIoaLhM7gXbbfTpCGubkTGvkzHtyh9H1B0B/1dJUURjm9zatC0t4R49sTKU
ZjcDB0VXOXNuavyPSanb1kRRkRdePHEX5OAwe5WuX384SkGmd4GgJKifg+qywiAh
wn0LGYwfsPZv2W8r4hhFuG7W6p9tzXOIf+TJQRXu2Z/WIfW0tMFV/KzKFVTXpoqY
x6CgfJggEZds2y2rsZItJDn0Je0+gGjm9iVJLhX8LNXT3+zod/kYe43OXTd7NcIN
F+iPTB+PI34IEkNc9Goq53+3wWShX2fMJnxcZVFiURkD3KgISehcke9y5ev7VWr+
3MIoJpouXcRcm1ahz0OV5b+r2vurJZuE3N+xmF8sLZz0kzgezMFpgi3zU8XXd8HL
+qdPUcsPENfqNOoUvciOqn0zis4iC32CVx+yvoOcSuHtAREpmGzh/uR5XkC8wC++
a5+KNdR8FGkYfiTNFaytIOudpVp9nVSc4d71qbP0ZpVmzlKrT6EruniXtUm95OVE
w2rmtzOzgaFjD7tNfLqYfxyLhJUrIQmZ+7sbHB7yVljCyO0BuFTfQTbQDq4A1sZj
upv20o4pF83d/LiZTpjqLPUGhyHwxVEhrjW31cGw5lp85d6KbVxCezhfgtsVgt13
rWKvJPhQDUnLRk+tTOhHHDfMnX6GDoW6IdWwqajwwQag6kiDqhn93qi0aH/Uxr9Z
8kUssairKmAzsJKb0L0l5q7HElOad0ihJDRuXkcyqJO4swbYJsX0tyjsOwn/81rT
tofl6xBNzLm7IKNYCabOodSuJ1AXfTpyTHvh/aLDd16/9fJuKgNdlLKmOOxv7evo
ebpp9hHkYCY19wkYlFBYp4vPKsFDRY6KqvxeIUJRfqYf6jH5kckC2mG5JIhVuBYg
DKJD6UWLOVBr+PhokRykzf7u1HwLTWInHZ91VCrn+zCfq/MS5HoEHWtxdfxwssNF
R8wKmjbEqkx2M9lwRHtNgMfTnWET22/ZoUcgcMpRzat5DkxIHzsSTc+YdzsocttX
noWaUsAGMglTARM98K65UxL5XFXTvWQnj9/I79uVa8+G4+sXdO7so/pAlSxyp12Y
/iatyidU7DBEfd6oFd11FFd/mp9AOeDFG3/aRl8n2kWqcJWsSpcmwCbuNa+H9+Ck
4XTvgDMbgBIxZbHrhmfRseAieITyeSneimuDvX0Q0Ii2wwuFfWtC10Qr/sXuPVe5
6B5S5VebnsCi5h3lDLuq85o5NBB7elq9fYpWYlI0c1FnBWhiafUHipAwJvLUE5Lt
Dtny+HI0cb5ISnFqG99D4ZUTPEt7HSEOnjrmXaLX+c1fjMTLW+AGIBBT67J2Q9ub
SBBNyPZqHoByfU4o/oiuB/V8bxdw0rMAmVVASyMit7tKd8cvl4Z0X9D/ta/b02NL
DCe4cAuBM6GMpJN2MQlc2uc0iNqMp7Y9jN8sqex5a9r3jwPwuR3db4ovuywfWf18
aRQh2Of177c6rTfm7LloEWuTxU41VMQVZyH6vrb6xe/M0r7oD0W/+uoMc/GsmqK5
w+1Z15nT57F98obsTNSu3HuYnXd9S1jD4x7GnrP3OJpb2VIW+1I9+TkaqYrkrBkO
Vmo2LqAcjfBnHRMBZg8RCxo4MK4Qkr+qpoye1eWLr0Y7jUYSzIq1ukHsdAVxnORO
jAcCyI3XBjWr1/UxLnO2OQ8YCN3TEAFbdotw4SzQrcA6XQ5nNEO3gee+Ip0MtCuw
qGTsi11CBQN3FFmX4V/htHzmw66NEF9ZiWEc35qSgpItJ2WCHs9QD0ffY9noPWXz
zavB5qvhefKQ0y2yLw1wcF8zO6j4fgX5COjC4hrjTt5WveI0xt9ZLKvoE5mRvhOP
cJbbf50pKoQCl37V97tb+TxgijwS83yyi9gkIGv+Z+y9suIHWQFAvJyNy+d8Jp7E
hbtyfJ+KOiHx5sSluWp/034WRpCoHpQH7mTYO8CtnTNDrzDjx/FUk1MDOcB526uW
h6fjbMlRoS2qiU5Qa9wVJ5nPlWP7d40CNG6ZNCCIFslhlAGEnYCw61ByTLkdl9Mb
K9LuYYH/VJ1WSc/orRnMH544Xrjz2CyepS4XwpFYXxrQ6foCpREL6c0QKZppk6ef
FTUHxhIseefTnlCKFl3k2rgKn6Q/v1rZ51rfd3MKtuGumlozTIWbcGJSl861PS8d
Lb+MQLTcEc35XbQYmcC8/DNK0RZXmnfraF+3qfYR77Z53Rms6cvk/erhUKgwMIk7
VXaneFIrv4xCUMmX+KMDWnYsEAEGSxfv7lNemjcVDxOKC9t3pRxuM851wHZGyfT3
athuvIB7pT1t4HIAEipul1nxqtbYlcgLST6/J9gqsuHZ3hohNNphBGIjdx+fvvoJ
RUCcxVumQBkSOAfDI61FpKsvi+Yo3e10gBVUw9j5NfreaV7uniF/elRMPK6BcRVr
Xh/Q4fqtObd5g2JQk5OLe0R6Gy4L1G2PU2Nth5sug5wRZq9FU8dFTJOjH0UhMfiA
MVSBo8BuPh5Zg8yJZjG81VmHU9PCc1AzV3aie3Jibs88gNP4ZReAYtVnUSGLaMec
qUuh6QjgWRAbMpQqUyyH0JgluSCkaN2EE8BA/wPOBFBeRd3qfxgITrmDDTlkRduG
3deHfCzxLRFxyJDzro0NDHfKMcBiC6rUhZFey0lUrd4wtWEIK04EwmMRmHxiIvjf
hJN918McVbcobQnEgc9yRhyUUvz0VHh3ELaAy/WGe26t9WOFtv3IX0lrwdVPaPVN
fUJ/etU+/bVkuodFE1TJOsODQDGM2kU0yIVWfS96yzdVNg/AfFzQS8eRG8RQ3ws8
p1nG5nR1h0EYwTAvNkRTxMPfzPgvokzsbu5u1lqIhY0Cv2n1y9b6cY7jtvyCuLkp
WUcllM4NCn0PyRZQsmYVYMWJKnk2roQdqqodss45WRJJ/IGvJLs8j5Opshvkg207
M5DISWHToluyZzgOR5VEVZ+WV0IftaoEkcbRrqlGQBynM2xBpUVw2cik7Nq/0fW8
1el2OOektybH7FxCBHfrt9nyZnkC7MC3A1ueE5CbnNq27WkDK/xMLtIHlh2gwaAE
IY3PzxCB4h5kbRAIYO2N4Wh+9kyvU8i1Hk9g0hdmw4t/4vu6z4q+5akv42fNjigm
TIRN72OaqnUennoyVnqslVZO1pEoGWfbbfkhgJSeHMUt1mBPYZBqjvpc8w/YtJBp
TOOq36S6rTHlWSav0OJmhHKDs/RNJVinRO7J63CNeVk=
`protect end_protected