`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15696 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
wGRcZBVOZuvqhRggId9gWb94qUjT59JS66nSXDHJTvw7ZycmSEeL6KUbilBtkBcw
hWqAAlAGlDJA3HbKR3PqQ3lmv1PKLb06ZFHq4/Jzaelv8lxbJWxoijhnAdJN0RAB
J12tC5aEy/dp+XkeKPsAo79srFPzJv6iHkRK7EuEfBHv6HI/pRmH8G/4BI8r7dg6
nHyxd43JvYoqK5PwVsuL6GKMK3HH0UrAWfzZMfQn6Jwqi7BXqAfmU+JGr5JuJWXU
Kt70M9fxVoPHJ4/LUfS+sHMdlNisjX8g0Ich7yVFIs1imBTRGexzDzS+AYQGE4X4
FFPiPNOlxODiEPCzvWfLAnbFC4ma6EpGP9eNSkTlY2I4N0S8m3yUUhsgR2eXaPOW
vw7Ww7U+lq/7e5hd2sG2ni7tOXAiZF+3hQ0k2w9o+xeXI2KWDqapkAbZ/uXiDk0X
7yaQoRZJJftCa51iZ3xh71fQl7/i9sd8TkR8bEcy1BLXKcwy1H9AOc3B9MpYl68z
va2O5QSU2zc6Ae/ukDzki9NZmPRlpraUKDPKvZTJPteZnlPjtsVW5LFlAh8q9dGV
2sXrvj14p27QJlSL0r4M15qIC3c+gS2P2ZouJKaFTyxiXCvFEVVYG54QXnlCx6VH
XOaFoT4rmX0FYgbm5nZqDOMOWS661+xmwjrg5QPNkiFZTnGla0R1EnViG4jVrB4f
ATnYpO57BmL1ZMxmXjtkgPypM/5zPRphbNMk5UBxIFZhOOFXVRTJJjaFCtII1uBl
yxUKv3OstiO1FtxIb8N6hX1ETdK5m6GW3m+cFAvnPusAx+VlHatN3Xk7QZVvzbHN
31TEYcAsBKLS9KdggNkGcIStN8c9HaQhNFaQKjjLBFgQIJPgS8dUh0Te/l/Iur+J
xR5M2OgXfnb7NkUj9hC8n0c6qnYvxgOA9y3IQEV+gTs5PIO2aycuWIQlLND6JVtl
dxFZHrYUDaShHWdUJ3kzGAcF31q3KSv9h27x3+Et2csQY/FpNMzSSuCYhTGQLMiI
MW+SQPWedRDx7n4/9GGxvcErT6qbVbjGdN5htr40epBPh/4kVAVGjSKdy4jod32d
R3WPP3vv4xVEyULSQEqNKq1KqBaLac2yKULwFlgWn6l87rQk+Ck/Fyar09C3HiEP
qct3A3sVpH9IeqJ1WSEWCMuO3FRPZxN/s/oGKwQ3d5ENjPnLPBDgm6oexu4MqbGq
+pwafKGLn0Nq56m06nYaMLO/lgE6fAOe4DXrnzk+raM0bHBtD4YrexUhL4+5tkyb
0G586L5ZBy1lsHvaT8keyESgBD4BI+WfRUjrw2M85bCrOJp+bKPTefJPaYhXMS4H
tdn5KNmKFfiu3P4bRL7QgPwkJ4KdbTCFTO+r+AYIoRxlgqT41C1Qfmwl9GwRZz7s
pZnbf+x395XpUqw5Rjrmeqo2u9ePniDVYmTL/GsymW5VO4CIqi3KoWMv8Tqh0glm
Qw1piGBaXGfLg6mvY3SV3wCQf8VW2JoyGhTD2UmwesUMGSMfbWm5nhZ9BAL0WNT2
ZCkT88uf1R4T/eOUydzsukeFbuwb2E6vji7lj19KYQKinnQlo/HFHr1N16IsgeSF
1ynexpTH6L43TARjfSIoYwMW/XHtDhIgiJZHLmEOUe2I1+GvhFn/ZcUFry5uNmRp
x5zGnT3BGHI5roSplU4gg1Y3WOcnzmS5nDFR7RkxKsUIUEYYDDDfj2gqmKjVsa1C
XKAF7FzzcjSCQQHx2KfzQliBkNfyMW6aKpjlmFheEl5izopECu7bSDpksxDkCrQI
MnhAhxT1Om6XeNQTc6CR7xyL6wWRPdXuzr5zzLA8WwMRXaz+0fKYblLLZchWkxC5
ZHsdkeYcftRnN4ZBed0u6AsU+aQPJ64AS25wYt1MA4XjPIOPOzoZHGHzmFw2Tg9b
kBhlb7e472Z3xmsEut5xoxtvY4UiFnB2yy36GQOhfzpJ8z44Jb1t/x3X43NkVAmi
J3TTLL19/Rq0R+Rmf55CHA6obPD2Y9ibnvWAsVD0ZeJ8hvkPLhYQ/P6FTv5UuD3D
KBiH6ZYQOCZVIHOr3jd+Asf/f9Y+/QgOpWDERFzb8m/K86OFsBtQ+4U3FpnlZhDQ
1+DVgtbXcCn7xoxVA+6dTltTAofO1HnjWqtBjTdQlgPVmPdxACeVzi/YObdl3Lk3
mEl/zeS1shscT2NeDBnWHX10wumwLCrkGvgVVclgi1jaZuZr3a63XnzS8I+rKCgl
/quNWeIHEae/xZ0B1T/voaQvctTspqXDUvUDVHwRjaMs9BUg5dUCxLk4DNz5bpmW
okbv8N2eIlX+TJUcOcexTIlwH8cENyZ+KJwAsNQRflpmrXRGWBUt7iS8NoHTHaIH
PcIFyPel2QJ0QsIfHt0OQXoZNfkKDvkZARyURoC7W8iXDM4xFwVECJ6gOR++zPrX
c9vfLqq0QXZjlR5lgUoGmrWq2at0nIGWl0/piCPD6lG3zHR8gISsH65bJa8EtRov
2LqKP5CBzN2trOuMa6rSdTCSF6gPZUgxrM33CUWkM+wB/yBtjdXPM1fexc+IcC4y
gHg2lfrA+wzYf9IW+cGvggN110Jub/xLhZoDW9UuNSGADyegTckWJvKACjtk2kxZ
CVsroZHdMBTbr6jt02rK8A8vZTKLcICEo1C1zIbpJPGAA1eYbZnR6oodf9ZlSafa
TxSJMa4pwftDNg77uw6H5l42L6NFyhjKqG3GQQs3ny/cX4V95jtjTwXGcIV6K/d/
pjxpH09X2FuQIHG6rv9v89upPfsF/lHSBVPxmXDV/7qkSe+VS+35ojVq1crUnUiB
Ct37x9qcUD7084tXHNn6xLWP1FY2HS+DY+oJk7ovFEm01ZEtczj59l0l0NmTtZZ/
QuVEg2c62IDHWBysBZCpNR4W/7Ho6tlMraY4q87Awj0g/q/DvflEOXuNrrUT8h6c
n79LymSlTZpSEwCybMaimC1uwvmIBdyiNCoE62hZMr/xUVGzHDLPB5h5fc3tICHk
NDtVrosmwmzvq1808OoqUCfGHaA6HodbqnLJnYjQVaO8HH2iEQaLKx5Zqvd7PGfH
1dQXvTnJUsa418ugA+bcIX+U/uyAFr7vlLCjMqn51n5r2K2nTZCROM+a+p93Wv+H
vkEd15u42l9R9mQ8yQBJP6DMb8TJCrhyglq4x1XiGw1KpshFTCrDLv1GT6q1YbEa
KmmPZASydCtLrxYaogLi5/zW0Kn2xnntySQ7q63aU1V8CF0hUZC1+o7zbRQe1bGY
d75G54ZJ8Usgr91n/OnyVWpU0rQLl4A2kjCfjPEeHmOcf48htspWWTJ8n0S+BjBI
ATF8slSedk1Fs5eurGrSlUNDvLU6Hwa8ks6X9buKCttfHYjfVqsU6n3ld50yduG0
u7wlQz94pIByexVfLusZlH5Fh9d+zNMrk3GvLz/tCDlfJM+wfJXtxdqbOPk8FvUL
Vyf8nxM+raBs8d8WrzFAY1V2XlFY9wogOd37fCrvRS/OkcQdYto6kSSzcMTznxso
6XUz6dGWGd2R6grBon/ZLDZyDLkDaqEc4/4fEBvpFTbT9ixtrpwGXSjpe7Im3n2S
7Yqk7xhv8EQu7SeRE2AoEcqN+4P/Dj7lSGx146lOqq/rdg3YAxDYKO1Eb3XuedVV
q6HJw2zbfZ9yGFp2UL7eATgrVoI2hx6+rW4/ztza3xxz0+Z+nYN1hwgfnM0dd96A
n4SDs1Z4TzZcvdKR+YH5rRF76VMJ11gqHezbzC2xH8hi4YPMYDuSHP5WfWGy8L+R
fqcnFSNw9Kj677dw+6SbxJBmmM6aDkvrosGF5BvWDBIgn8hZZAbQ8PBfy4tgntVt
LDfViAko/uM++PqntiPgDD2twVDcOhXkAou6YjaTD5vIQxRiRNAhrRK/YInzI4Jk
AsNVWOPPOpv23A1AcQtVizVt2Q3lokgs+9spjeR2TyhQh/cKbVbhbmpjXfGftHkd
WzqDY6GtuC0DV3NEoh+7fqbLScdU16mKgprvWOnsljeC/00oAgkZYWSg620HyL5E
4uiPYPTEfyZnnjZbRI25RglxEEsQYvAJEWZo2TT3nlNA356khBOpQOsP0U+wH8px
kV8ZJy6O08/Tbih0ya2VVP2nyR1tce9xzINvf6N+gdycB/r0kszlaC7jh4nKbnBT
ProWUx8rL2AAk7WpSWCSaIsS4cAv2XwiHLFO3FDhhr/wMbzDFpD04B1fwkQReZ9f
gEJmbV4jZ3/+jA4jbK0cG7rikCsYdX8mFTKsPrGtxVUf96GecI6RkNE8TJM9uX4x
M45DJwYGqy2+oBMBkBYW9ShBfkVSh7xGL2+8mmZVTJ5DzAVI2ab2RkjvUM5tQ1LA
5YkhNVOBkHVZTqZYVzmGoarWxOP0E6nIqh5nGE037dpmBUeTWcOr8ct5prtzogCj
DEguis+t9dCuxnWn4aDdvGEDtUBgfTM5I2g+FYB3EdG5buHGMKmaAMEBaBxYjcW1
yfnNTfbBWRtvI9FK0dnYCoAhgTQaAivGPhHCy1x3/29TRFzm62KsJyBRAeJIaFLT
lMIQxxyHLu2+6BOtJM2r5SPcgWqwA6Qxrew4QEDL28G1DNKBVmBf9t2OrqM/P0YX
S6xRDiQSNs/sqbSZMGHdoNrp3Wn1XEvKKqvgTTiMlO2nshH5O0dHNDwzg+ROmy27
jw/wqa2KE8sOqpZGGconL+8kXiAAwbJynRcxLeLzyMDx2psTIS+48r7Kq6YNjac6
UIPQzxHmn9XNVSlH138nP2x87z1RwZpwHj1GNogrhxovXu2K4ddcT7MT31K3Ej4u
zBNCifFN7rshLhGHeHuDhBM3MVo96BHKiMcX6sRhhT0d1AtiXlKPTkE0Chd57f6l
TAnTMpGcVNeGWImTZXgnXIjksi/P+zgy7Fm3bwHcKrgRMzQytz9CUUBezFy1l0AA
OQdljlIf3zXIpEL3shqAPseWJtBYCwjtY1bnrYIDbHH37HkQhSsmQ9Zhvia/mVgN
v1hURUVTtJzE7KJl9mXu4u1uQa4x3tqHqlSyMvV1DRvK2cdQshBoAzISSvPEVjS5
Bc9vI3X1VK0eK+cLRYxvfvIZA5hfldAgohjxOkZ6Dhkrakwgka7ZMrpA8WHT/UWB
CV60mI3tbUbHbN94XUu4jmagw1U4xDrP9JBiY4lUBole5WAjykXbFukig7Be5EeH
+NMzWxVdu/l2rexQt0SsZmNsw6W9wMqim+jW/e2CIFPxm5ooJd1OqtSI8BYt8IL2
OXk8EkI8nM6gQyadC9pKi90uWHOElVDTWnGiqUGYsf+47NH3/J7TIF111e5EEbnZ
fskeWUz9LkymbS76LLb3BkF5MeeAMD/tQ1dLOdWhNW1SvS6Ze8mKTmF6KFB1WYxB
hBLI+asG9ncDDiTTAKXNiRxGLWv98ssqqi3HI2hod2LNVrHYBU0JA0jPqa3hvkzx
kKBBoE3EeQgkFaBYtOT95Lm6dcf9esnnC62K6f2bbX0FaA1zqQqE9RdFBtX8L8As
bFrbVGYLHsnN/mF1MbRenHOFjhp8wHZocXjRZGZVs5eICFafAr4NU6u9i9yRxdnj
zktc38o7oWMRFStD6XxiuhJZqoOuSSxo0rqgCZ7NXwb6FFdHzyWzfme8hhQ0wtKy
d+TvoYLWiALLDzusX/Tz9TlyTuCj2XuNbFKiIU4rodzk+yngYf5BpnovyXCx9cld
h0qCAsH55tGpILe5rBFkxfOuWbYkIAUmHJ+l2lGF5gjnEWXAfl7J1HebxTHn0+B4
n1KM9eHy/YE7O8eGGm5MHYVdLWSNhokMNoZZYKVVROl5X5qitU9sTukAD+F25EXv
5ldzUy6eEcRx1iWXFqtbbAMRDWgFfaFs45TFZGNBe0LTASwamlKaqO1ZuLOy12Ek
3Z8sy6pCmmE8Hc1N/4RTW4LHUSCUsinnyPtGC4cA/8hOJOj1Ls8L9hwQCqmFmAW8
FNME/NjoA6kCxLcconKwTqP0kd6pgWSDUa1ldCDNuGUJ3OqHVLE2LwPSYI+Rdo60
svez7tvMI14JQJC0y3RJflR6BZ/g6d64bEIIu1HFL1dF7FTPT19xQb5t6pc8AnLf
tz5YwlvTDRlkwblkq/UZtWlin4RMaNts/8ULLU3Oe/h9lDhWIlaUaFQ2oucbzyoJ
tTDHnS05hDkMFCRA6CJa8mYKTDR7hBzz3nsFUx+8X91mcP224VetNyKTiVAoPIru
Y4jFX8WUiDwnIcxEvLPLTvRUX9Wm7L+VXmz3HK6UK/1Ds7JiLCHnbHSbuesSk+l6
7dzVxszkOVpeDpIw/mtDQXu9HhfIaXXuMJfI9eUp01DMSeTpHWmxqNdhU51R3eVc
5T1aHvJu77WBgYzJ9h1tOHOaRjHDCaaxeqnSm86LoJpcyzIFfJtyO1gP0G5lMpXI
sXLA3u6LVyC8XrF4lMBafFImKB44x1AiF5yPYpY3ItxMjZo1M+U64YZEQmTzTDxh
OmeQGCfZQFfo+eY2tGKskTHhzoEpHYbXca5l+6oxD7eTJ3qLv1DwJ2+2rcOV9KAA
yKgQiY2cLYrTVx9Hg97dgnc7t64y7ibFLL+C+dkN+zYviMLYEk70yqz8ZWhV1AnT
SKG7tNPkR6sNDM+CCyPK/A7ePrv/Cs+RMIpwuBM8+sN9tcxx8xMOg8pMoFyOdHWg
fXtcFoi+1WS42mfgMXu+Ya+kROCcg0ol/Di/Ugj1uMPTKwa0RFRfAC8xVsvx1/bJ
h8FVSzNraVQZm/4DyUnqgpQPALkSSNQdxrhGRbVA1IbymfjoAjzloRdhhPLNry9p
d9OX1idNqC3XzFf6i0tzDejCEm7jg/uVKOAxFZdJDp8GTS7oIzHI9UV66xVr/wAo
N8v14jMbKr1mOqXDMMComNQbyyVU37i2QyAhHwt6Mao47BGpauU/B/iw75DWnL6b
FHFpOG+PqPBl+EIGhE0furm/xCeb3YUHkPwCQ78KK47K+5x1LDHAGy08qSmU3MaD
W3PNjVc6fxiibYFjoCWjGTCM4qOPjx6ZFLbQ9osyqY+kqOmXtAq9dLcfv6iERdfB
ZLv6cNnycfyz+SZrgjSEgTe3x0pshsZ+4h9aBGk2Q7bnvFMDrkCsN4bQNq3cRxzS
ED8gQxlZlaoqvXJnd/N4EztnwT388aDurun/FhqmOjswSVPo4lg6IMQBFy5++EQd
PfBCR69DGG8BqB0rAjFcNaPnRRVEUBZy55YFswPeqB44jotYMBzs3Y7V/6quNNAR
GbzbArFDHxE4Ld+NXcQ5ZgAPoIZOhOErjuwVnPI1r5IgqUn2gySBhhI8jv0+6u9S
oqryLQKjuHAOnj27tINUx+q8AnAXX8zJxDHCKcmY4DgkhbePgSiL6X1ozHAfeOrb
2j1Ypz8CWj/SxZ9Ja0zDGGRAAPzsYl5Ndw7HjFtCc8UX6rdHthG5GNZRM0P/Dil4
MfN81ceZ/cDGbH+XJUGVgClxBc5ACWfrvRCti1wbxB28eE1jfaVDQ7ZKGBdJbSNo
JaBqiEDN+4OXXIDwVJHBY30apFPrCfED0gK79BwzhxA0otTAM1WqPF3gLX8zC25G
u5f69C0ibVRwYR+Fud8zWmp9dizbDYUI+dwezjSGWnBE8TeOLmgUxtKxm49PL0Qt
UZLFqEm0711Qn+uJL9JcrhgdMqDP1iv+lBCVyWZMqZbDhHvU0Zm7+HwYxuD9zVm+
t5XYHqm+ktJ/7CcOGa8lh/h4jf2IQ5KsWGOpPWlh3h0dLauoUg+cEmBAdryx/aXz
+DwwucMQxKoZoldxbdkqXP210f+0gA5UhfSCr+ulxw/3BvmOs8k2mhzGHMskH8yL
dFkoS5aSiHxd28ZaIH+wOm5/Lu29hsYi/ne+g7ehniC+hDuM6wxOgrQcx9NhH6vm
myx0gkbq7gDmTSgAN7AWxRBpVMTbvsUOUq6wV1aygcdLfPpWIVEkFYOVQYfQh5Hw
8VVXmn4JQn92v83uL2OGG4kiRbRrOqXsFypNbRHCx4pjStU7shflHIXLS/V3CXSW
fzak769jRFAYVToKi1iokhVjNTIFCoNEdOzk69TIlYtuKP9XuqaZHQDyYGt8QUXr
1DKG8lbYIFpqZGj3lGZPOnRpZFJNNH/B04J/34i4Bq1iwAFxY5A7q29iGvxWub+5
12j6ZVBG8z/1aU0tP6nY3luugSZftEWssfvNdqqh6gSGIVqOtk68XcQNVHO7c2OI
Urzilyyu4HEDFTqAsv7P7nAYPND8rBu1BBjXnbCNhv9dKoJGu5Vc6Hrk1CGVe+8y
dB6ruFnEPX8z/TYNTW5rtiCIZzYGSXJGUHzTn16B+QgRgy7GdN/0sGmH99B9nlOj
AfLBJA38aMh2UaXwmuL/oAJOaEwA3slRZCRSukGF/dTSZIMSQLjnmOUKbrRDCGWb
jaJwYr0DG+QWwtFNdJ4VpgCur3DpcYc19w1Xf/c0172DCpq4DG9ixzmVXUUYv1iB
MTIsCQ+u3nmr1qEkbNx27dBJv9sLzyMlq2k8iEuxBLhX2t4TENhjOLePtRt7oCUi
GNMUrh8HzvtrgfSakv8cwwA0TgtrYKM1dkK1wAEderAzLu+fD+peeqeYnTIs7RxN
lECVLwXs41YOYQprRZ0K05fz3udd0VrcpdWOOb93Aksjd52B7iEtIWvSVdXjrGUo
vL6sBOGzVCNmJw8xkBf1MfTv4V0yz1OTD1hazdnHKb3/CRFz5kEcjmpGK4XqMS5T
bvjAOKRuP02u5aPxVwMtBD2Czz7pYakDPTyDtAY2wNoA0zx8QP27nSiTnq9E7lyv
dSWAhR1DgQjfjTwfOtMf4qUhic/k1Yy41yKkiULDB1BjCYsRkpFZ1VHlumhBPTv5
/slMZC1DFcw96nu5Mi1UAc3GPy+WHgs+7XyyaPkf0qGEcAS1J46Da2p8DViGLVUg
fPyeHer6Bu25RTPzRLpXd5HTGMkxGdjQV3N5yEOank3D1TNs9v/xWCPf7tIvF0VO
BTUEHfJzSJZNkDu28t28C2yIvQ8FKBJQqaF0FFdhxBgxSyTSCtHB22OV75fg8ofn
NbLphe+AdAN2A+LjzMrS+o0YTi0ahII6ZOPH9eWU0OYjKDqTY28YPn+s8eMrNpqV
TRhLJTywc6bIAUZ0jjWW01nZWZruPvANFi2gJub1Aoxzk0/OycGnEPB0+fuLSpQn
3TAyeqFdvsYJCmHXX9QS+VTeEqadCNQzYbrV58HF9QUIvu44hQXwn2dMX2KO/CxV
ZFtmletPmqyLMUI3FLNUDX21bSttMDZSBfmOQOo6vkU8qcboFb/RGT1CojC+Olto
kcUFweiu+cAplN9i8/5b9nkXrz6vyBCLngWG+LrmHDiWsqfWJHqydxlOFnn/LUgL
7P2KNfte8IRlbfRwnqWHCzXOS1nwbipaOx5mxXB8FTcB9Y/bjLkq11EQm60aTtee
ju4+oo4h72D3A9ZFAKJWsg4wNtQDSy7Y+BT2f3QSJTVGhqxX3eBDSOQjyYt6SHSg
+oJjBtX8QlWXjJ1+YqB/1tKuHz+p/gi5fIn9nb5Q70s6pK0fMGYLd7JD4LRZrcLW
DXPiWTlmMrNakCht5gUD4fovS5L6LGdCmdQdkDRTnuV3mb1ld7SWSNTdAND5uDCO
xATRTMMjBBspdsFABP459WXehMpdnWNvJQNpNTCU1wyUVCwZ59YTrQKO1pVB4yzC
AiM6/nzI4aX8Joul/QPPF7sfzT9IoiYrRC0H52PdT2rJLmFAa3a1IOQbKPx3L1Xb
95v67CBei6oDxcMSZgDNgwHLvZwTyDP7n+lzKwUhLAHuYwH4aj770sZy47vb+mZ8
Sbc61GiC+orujRqYoLT5tNiy5bQq1YXIVQXjm1hFMOWIEw/eKS+npagumF+1x41e
SsR8G+K/saqQF8c75iHMSIuv1jYlkEfqfQG65AMitj5Q1b9nN4wID6B5HeXd6ZSL
c2QyLxtOQ28+sGOXFdW0brK1aqJ6j+PHnm6XEyfVpgO7usBo1et0kGArslOVFSUU
UIjlF2MxSE0CmpUhAid2qMM6up2gELKdQrpybK+e0XXRqx/OGafhkqHTwSsadFS1
QbqRtB2KB/iiu5tEddXgVEVmkE+rp3WsJlOLgZmDY/LGaQddjWmJ8joJnsiad1pZ
yA+nrOGSCu7vOWFEd1COjnrevpNJyPjakdp+1ciNviLdbm7jf2orfthC46aKJaZR
sQ2lpmRr+usT+5MdFYqk/axgsdSCkqRCId9Ns1oveXZTP5CfTuaBBV0LKs3ZCrWl
pC5nB1eQjisSD9FAMTqqFK1UGkNwfZR/ltSk9/erb8pywG/R6zyQ2LBuQ8ap8aYt
txGQfAhhhgjdMucHscF3JIUqm+2ktTVEyI/FMMEc1AkGinvKs2k+XLecMF/L0Cn3
1BAhE5dtRdwxzTxEbnyJddUFWtbMqa60PHybJYqTtSHqyY3il+KQ6HxGmm2dMHAu
tzDQIJwHb7FXZYo09Dn5Udigsag7yR9rJ2fVbJjV6pqfzdlcfkV1/2+j+2VfF96j
XC2e5l/XqsSAiV+m6B77dFjirtn0gjGFvR9lGRPudtEsedHZv10oBUEUTPVlVniq
XXDprZ0SCnIhGiJ7K3knwSsr9KCtlQ87CWfnlyXcVK1SN8VqsxlDkRr/pYFhxa5H
fZywVJmKCRdswJ2bfv7FyS4+ksJW0Nn6uIA9xaNrEP/h0oPqMTDFuFEbGWpFJv1g
JMBVk7sr+R+rsjO3cmx4VAtpYxbPi00bP9vmY+xAtF8u61QgVbeDPtYGgYDqeWAi
aiyIsV5CC3WWNCWPgik/Macep65jsY7UIxhMcjZqsXh8HAWLeUATi9DTSDkFXQ3t
zrMwL+37h8y698vV8CyRv3vRWiOdq3KZGzjLqFgyIBwVweAKc2M+dKncDivnHoHM
oObJZxfux2uA7w4ccU5Bq+lRRaP7yHSIDMXRAsuZDogqLNUH7jV9i93OyhSKvjQx
+eqGQN3+Ru+R4xFo95fLz7loxABVsGYv4ep+kHmTKFagRmLZJAo9arfJyGi8Ws47
t/3ni3eyydg8z5J/M01j9jJHkyRnII88VoeAfN6Ol5MJHBUQEjDXEkdcIZGyI9gx
7vM54NiabyaCNSSZLuACF0fNCdV/dS/sc+bJrJewiCbbdgwzswavT44DBPqyuevu
oXUDFBG/GQfakNj4FjUMAAiMLW00dkN5xTHgTxpU8upY/g05mIwZYyN5zTbq+iGi
hWq0bNL40y2v8cb7W56sP4QTNrXp8N+Ba/aHZw80gHP1Kr6KX/i/bZ+vqKALVQm+
Rs+/g5p7OKQMOYXX2+l/0NwqjH29ct4aj6FlXVp82DSfh60S9Jjx1nO7JfY4RM4a
uYYD8A8WYmIS7RSRYvN+AOxSQwMIbkIBDVlkeCRCjTwPZOznRufeSOVsFuzFw/X6
cO1eycC5Ri6xw8TykOJVgFGTB6sHlp06g79ZmUPDNl8yeR7YDOBSN/B8sWzmrGS8
wR8+xbNv/v+HATOqtEhNVJiWyMRny+B54ncOSI1GCPrgNyPZ7+FwEAhwtqNTKqyO
ZB9HE/gPilB/xgQAkyvSq3scF1ihyOksmGtNN0j8HJgm22ul0twQuYYtgDwqMlmK
pP7jXHlJT4L4mtZ6+wqQ7hbbZRgCkBtkLhN45tAkRMNHITZ2vrI8ZHqjzhFra5lQ
wGJf/6ZdhCgOyZpdS0VLE0Mw5+0vVDHOGYRqK0bLDeiDOcw1CuGDv4W3560EANxB
KGzHyXYF++Jwyr6Ug2ubrrMil05eQ9GwOaayiPHOOe978p42hQfdnr3CeXT0XmsH
nwKOp2rIqd3YwVtc5a/HeHkmt/a+pnOPxZ3/v9KFaYsdds+6cEKjHYFs7pNr/oXA
zhheqkfkjQZyv8H9EvoY5ERIEz7+M/L/lm6DwqcSh5zdi+EAagX6WppaFIoaywI/
Md0xVqO8BZ8amDbkh5fJnk6lJIkQBJpQA5BG241KHTNCEJe3oYsRFlVR9Ue+hw3m
0KfrbJu9y60tWRFvVntv6Jvyf+l65HrVZH9/ysGszUmjLv8qcEcHkpNCQTTpbT/5
lPxam43ru3oTjKsW8s9VAb/BV4PH3ebGlYIHQ+ECb+5Eei3EIECsXwFK7jpnDIWU
yfJdkhmaU9czKMsr97BIak1Temn2x2DqTBaLmSbS2rZBr+fcWJJLfxtQp+5tn7qW
Z8MdF++SwcjJVrkgGqyl4NBO/qCroplehQJYS+SAsi3oc58+LloC3j7R8Jxq2Aq3
MKXvRHS+G476uc6JSGo9ocjTYPu8BxK77k+iFrh539ne1AbAZ1CPPiLsqRnNBnUy
LAP6YDYEcL9PiAQ27+g7VTpTesZ/C1ZXwGV4m1+SBt/fDi4E4K+APGyR1mNYoe+T
6iFQUr94FVIGqlzXwlB13pnq3E4fpjWAFcGho0/uiKNwMdSPWOjGu3i//BOUdtjt
DkINvs7uwG/ydZGi0IOeAnOwHkXXADSRz2mnGCRuwEqxdhyhicZ2Aumx7uzJsk5a
2yjZacz4EVTDc6P5koRdFUaDRnNz6bfNmhmowEte7y5dqNpf4e8ECbsUSr9pUxL4
25hObn+pZJrsW+YKPYN5Q1h+L1//rAcWkr5ih1dpjjBzjqcSB2E3KFiuHjDJdeaO
TCdNGwHirVb5bxc7TMq940pm8xmwu/ZApzqYCQO0UnhuBnI+Ze9UbCd+92/El47R
NGl0d9bUbw/pxo3UGLcd9iHQ8IbB/Tl+Nu9ueGbiuew5I6FgX2+dr/JO94/7v2CG
Fa5yT1cyCLJ61ozpuE3/c4ifmwAwx3G0CSs6sevKYP0dZQ0EyDUL0NZhy7juDqpv
2OtkP95T16IPFEOxbzuJdv68ufGf96vVfvpqOM93lIZkdyeeCqoo8bFs39/3A8XW
m0j5lMCHaPsI1oFTZD5lwWS5/ylS7PIair/7J6RLuBTAOaWd0mFtq80qYdl4zngk
OkFu8prRiDMDdo4QNVeDy5ffFi5yJ1nt8cAc2yRROve/DXzxNn2qqId5dBj3Un1h
PRbhcREWPAqh4mSBY+bwahD/zMqecpOZZUXjmQa0/hSkKdSS0huWe/TmiLBPUipc
gtDaDfwiLZCMDIPf/SYDQo8FpwOf2Wg2M2kH7ImfMjp9K8oqbRAVOve8k6Cl0PEg
GPD58UzTZIngbiSNGdCZ0ofDvEHLevoHTp0wbO1MGR2mWEphDHfZKVY9sAFA0pAy
ty1CyRXQUKRXdgJR9iTQ/tXa9OBn/ES2jKZ9YRbuD9oj9SwOv5b0ZpAAgbO4W/1H
QpT4+7MLLYekKRRSrvgKjra5FDyZEmJY5YmkfwiEf8/eFd47eP8A8yuFlzUO7npJ
WIy/sT+kwXQW49inVHokna9WJff/pcjagHjDqmkjcsPmtrFhTIMbXge2ztRLSn1N
kGsP5yhYy0Z+HXsbRVuC3kYKMwm9g9AF12EhLmeffE2atD2Nd6Y/zlvzvcUa2kht
JD3Lz475lDtLNOKF3gEU7oVoM2CIZ1zy/7EZXs+HZD16HThIHvEYis56pvSXWxO3
ouzFzJgqgWxC16ZeHXiew6ickd7RjZ5AHoQnC5cs5c9xEdpp9l+HjOGg6zq/6cW4
rdQ/jrS3Cl+e+CX6kzh44jc0NOGF0ynhZMleEaIOOeM76qNd5MXIRUEaJlJBOdWK
+qmelZ5PxeuKABx+1xH4k5OS0yMzKAnmAdq3t6e4fM41O9KCPuC3Q9Z5p6jh9aca
XpMPv4HwmHX27tJxFyfV/db4MB4AGbLy9VMsRiMm57O/ZX31hfj44ff74DlL3VpK
OJR8OU2QHPOpB1cnSCZxoX66fCFQ8REIji718Nd+V9nicAVs79uskTJSmz1fyFje
LDI0TEiEzy4ez1fAZTiD53dLkuJmWF2bzedBrBJo0wReJIFvjQZ/K/N27zBg1zGP
4kVbQFe55xZoVaBAiAfEoYxJf4fKdbz/wuz3da7AQ2aUybD/ac/pooY06Z0baPkX
E22qGN2JF8G1ZFdtSDUwmTR/59Ujg6MGkpC3OqSVrwJD0cxb9K3SkHRA+nhKElAG
jk2opSW60V9TkLLePUc1wduhYUCcfd8i2e8QQanG6wtvn19EOzng6jGWmzea1xXa
e/lWLKCaetY8WFAFacXe5YahtfhKlWEshO2dFcKNEa1ORYt0EGSURCFWLnv8UDtn
inQLE5rgUFUAzaQ7UN483YUO+MtCA+1cMORt7agNWMj+PZSpJ9rVuUVNjwW/2LI0
+dk5UzNTQZ8iDo+zgZyQq1+5+mF7Bu3KufaoeheonLxqQrWeh59SHqyYvKjj4NOC
lQ1rp0vb5YzQnNFHfPsntY13iC9d5TLZXepiW0sDQAuB0BxcbTE/9ha3ZyT+aC+C
nlqtSJbjyb6VPsWSx4FNwvu+D4mNs9sMn9by65DZAr/TDvT89LwKhVecOeSqoQ4Z
nL1hgbou9I5zjpXkzitAaKoxHURvKZr3nwjQC1FtuyJKVELzLzeCt1p4QYbxxmpD
AeTFKg/21h33WiI/U/vpHlkTvadb5OglJWX0TG4c1TEfcNsNZKyzhCEFRLFqLFPQ
nZ804kz+843ExqhK5L11DtyflHlfBROePXPK2M2TmuLH+dPtsrMnACa+D0c+hXJw
c07a7W70KeNIf5q1BHo5fTjxCQSdf4t/QPe6fhSdaREn3rvf1yJUj14H0xl2cD4h
+N+GBF75+e+TtHKVK0pzaYmy0/4UEeQ42nq8fo3je+JG96PnQiuUhWGWevAamU4o
Lot/dxFOGFhlUZmCBva1I7Sp00AaBSYx2Lw15G/2kZXg2IO7dmLO/zbp/JmQ71Jy
1oGbd6ZxhppgiN2mXPn5QG2eNFD93nkxqSfFN7HPc3bX0yHsFnUp0v/pLfZJMm93
MumK/RbXaupglvknL3HJ+eWqykMErAG/jIRy6coEew8aAIxkX42CbaxhU2c4TIrR
gHCi+T1bEBeSFD0bwcTWD13NMnQZd6MtgzZdNx/G5fjC4f8BoU3o8eprIci/Lv2z
Lj4dKzInBEpXAVGvnUvM1m0tzqk/9jMnjzs6MjK0LexajFpwkoQ00aS7vn3gW/rk
hx+tLYOAsMZ+kLBLgShHCjYafdt3yz+MMjFwIw0HfZR++eViRc4lUrwwzsdsZf85
cNDI1/VBsdT2MHfw4Mx9CHtC6pEte7gOczCwXLcCMQS8JG34wyeKdzqaGyHoSoFD
E3jmVbup138P0oYjPddvpss9TlnK+MzzdBZZMjn84t9XRhrlSfXpWnlmZh2CyRDM
QQ6Rj8bx5onDF0aCviWbZEDaZIAYwexsDxXfyFNOHw3b9vJ7bOyYRlhMTHkZL3VD
AU1qcOqW8uRKEx7x8BLqVKuVVxfqaSR4bMkBme+bHwzZ0T+xN58/6JNU8ir0ui9Q
1dSuEII7qVSL2pHnuhocN9/gXXftec1MhFvywTCoLhOz2NETOvF3OCUilprsAYmu
g/ObnziQujZeBlWwjo4Wt84kJY45Yuyd0PyneLRQ2DCodU1sfT4jlpmsQPMRjSSr
m4tm6/ZTLibi+4HWGLJufIv3kwyj+6bPE5JSBQOQXeQM+8h1orsxjrEfR0o84mdo
AAO7bqqJ8McxfepDpykaXiEzXJOM39r4VEvvQsSroyVCpmgCQxrehZbv5wVrVoLk
UacuY+9K1bDkMhUxp32Y8X3cA4RktiEvI6QqGwCN0/Zi2XwJ3g7IjrBhgWz6ZAOD
G24I804PSbmpaRPbs3UeqCOpiEfwjBEULS8JdM8E1iZN3unu7GZBDqjX/exM/phR
k3FIxS+pgEk7MNaWw5SnIob5DIfvZzQMRsyYrlJNKUoIx+DTInr6TrFbazGQMLKL
mSJQCSgTMfQHz8oyAE6KeyNK7Bh/SgdHgF5aiYLJMpL44kbc6lY/7rNAXaZLGOqW
IBAikFMSr+h58kQ8x2EEuMplD8IbwPckJ2auNymNtiY8Ie/yX0Z2eEjXgXi7aGji
/5r1ZyQCedOHmrWL+tPmdhyPpr9cg8lxBtHZevdL+qf4M7MpLtOY3eItMcMPZxtq
ApE7kiNFc93OhZqIbDbUhLDkg2HCB63jvWAZKR2U1me/R/IRk+qkIi+oGrAl7exU
mZIey0mgPPRxrkZ/zrWxuOmSshVR6PPEKgET4QOe/fVRWdYCkNmj5t3J2AsAt1xv
zNk7OkXvuIRLj9lE/4M9+iWMjWM6JyiExfDTmdDgUrl1CpzTIxs4F+p3XnFoR26Z
iOp73i41x9fg9hjhaNm+X57qgkwDjAhUr10GJs2F/ie/ynY+VK0qQZdvJMiiqxMw
6KEGBRV8rT+n0fSpxo/Dph1NS7MnTCTeTo1Sk8S7mSYuNGBDn/lvrxX0RuzNMGnx
nauL4JL51PH2R1fK1siEzHmEo2p0UVDU00YWoAsLZUhHvPvpzDGMyp3o6C+/N3KD
xG1xYD4hUpmS/YsYeMeJxEfJwiEq5/OLPEEB5GWLUd7Z6RzuFIvWE3tCORuxjk6H
dJHKjRoH4XZraP7ocnEnjoYnPV0JdcSTIIvsf5pSUGfjS0ahRbBIUYx3UoAiB25i
QYLu+ZkaFc08bsRuQ9RIJkvOYbMX9lHDFiLds4VxhveR4Vy40L0ehAt7UgcNJXJQ
q95opWduqGFBx5ZTtnPRgBoIbEqI7bhpkC+rCdqIIHC6wmc6V3JKBhsUXcTpAcid
EAZLhoNZJxQqsMvZ+IpzZp8F+YXOMBTlMY1yEhwJraKEmBJw0z844QtYwhPFB/Cv
uqtXcg6GCGrme01J9HMUTs6xBVU49j4qe7igaZ+GVwfqJKpxO36VTutBY4TBH7EE
8DplN9LGaSy3ZzYj1hXF9apR34c8rGHcnhpJf9Ac7Kscsp9qAJDnfXzmzofvhq6p
XsB1SZ7mJ/Hzr45W/N0VsKcjkgYXIIqYv6nGoOSRZ6bR+b0KVpEjHf9rdhjaCFrE
6xYcc1bggQ1wU+bMpW45MfkWKDT7iI6wuoxut/N9R/XaDVd66OpsBVbmydX5GvB3
tYAfZNCbjbGY8ZwMEVdxHMDe4kQS8HuLi4ia4NDM0MH3dUy0G05Ax2OFqV5MiyYA
Ca8N1zPyZhZ8PTJjXcdfDnT/KzmacVX3Inn8OXg002030DR6Lt2nJ+pYlxoVysgh
nvwMvOM1aBN03ugbvtBt4XqXdJveGUBxnklEohp6mMBBgMakwv9gVEIchJk/I1qV
CZA+MuX7YC9Cs7Uf4fC9cZkMWIFbKPo9tJlIQJL5/pr7FjMJOW3efhu6WuyksY+L
3lVat65HvKNjJFMrm75UY3ZzGA6rVZgGDk22/FqJeGf32IGozRNNbFZBM2PrtZOI
HtqipJhLkYsIVBObMqNJBSdlQDVQroX1iwk6rdy+moSRQYHeN8uhftpgp9odener
3nnbfY1NrJgM316nJf2W0W5WxjIA02iahSXUttExDHi43D6F2GaN/Nx1BztJ3xTS
gPKIIySmFYtUfiIsRGWArdbL3MFR2nvPKZkAzJrZp5X4SLPSijGjxYZstvI303VE
PeiJPycLn8iSpB9J97uLuQamQ58PYy+C+EfQ7uo3AraNOZxdxZDnGDG7nx1V8oht
5+rUHQRIieV516ClVAfb8EjjnbaHQ4lRcMOFJEiTvklSh6KA4O0nESiU+O/Vk6H3
x8do4/jlu/v+LzDc76ygI+E0oNlfLn9luOLC9Farppn8EJ/x0PoK4l4GaqZ0tjrl
+9xcJAJz2jJwCfzX4tl4QJ42mPZaSU30GmaRImRoqWUeIX0JsCNGpIxu1/YbKA+I
JWbcl3d3568sONdQA3SAzaD4M34hcBPdKUi92lw4klKarHu/3q/Xb/jYeQNjOSZC
/XyvptkYluMdIW7P+biFM7AantJzHQqSTDG7aU6eZX8cML4STOK/LHUvefot6rK+
aSV/JdZudaRcW4F9mRFRfHSRBuZih2fI9gad9WFF09m3bBNC47ryg0bHLzNb+oGn
8G5CAYFxJUWU2GI3pLwPPFMRxZYHDrJ6MqSy/nPF1IEQPSQV14/a6hNgiNI/BjfU
gQntHrwgspwH+X0unyIpT2LMyNphllz7+lCxKAPah/VOEQE+XyaGAHc58mTuFHGl
kX6LJDnmyw/6mJBIaiHHhc07HX3pWNxzkvPoe485xtgD6MnywlB6nzO3X0jtFkmg
FSAf1MPXQpmre6gsxpa+aAHVloG1D2JuThfMZJq9+Z+qd73rNEuf0iSSAxzTedwN
ruVzEdKCemYFNOBsR1mYgu1w7gDmuh48QNI+gY96sCUx8c5QxN4eHubC5zdQDKMO
cxtJ5akii6Nr82SsGF/p2VVU7pEQnrxyvun4R+zH7zbL2koEZ4f3GeB21rNJTcnl
0yB7/CdtAe5ti9DHgf2v4ghtw4Evs2FuVvTV3ZfrY/h6phGAyI9LW5LXSroXujOY
ilggJ+voTeeqqTWTE0c3CqB3wpo552q0JrIHCEfsDP+uiSQgkW08sW81Uozz/Py/
p6HK6J8cYYbR6sqY2aP4vBDqjfaLhkq+fPxOsVKXqIw3yZD9Pk9vseRoiJ5laU8p
OFGxwZN13AZYQJVGp128qapQyHgSzoDqBBJtakVnDp2G+2P1ngJ79pN6BVsA74QG
5PkBGSAtcH9+lLfD95sTPKWDZEMYQc62Ex730TDCLN0h2RqE+OHzUIf7e81dtD3k
qKTkBwgqGQTHWFioyCV5bpZgrBi7Z7wKWAcKDFQ8sLf21V2PfxggDjEXZNeTgUHq
LC3ezTZAnLx51JlHKqa09G1cnTHbKFtvH2dzSHxDOABT66I1eP4RnY6Nm2PqulJu
+iCI2roVjmlhmy6seeeIsFVHOQaSfWZ3mPX2WygSLIMhZJqKyVzKgl/hP/d9NZe5
/GivkQqlj2eIVCMjpuspkIffr9wyKIv1cLrvBV/1G3bSF7z6JQj63Ma/QwZFGsW2
55g3+to+DR9zMHgL/CRu3dAhUWHL9122Z2FOMDrYy5DMMwWYH5UGXLevnWjWxyC6
qjoVr0FrBLUTcJ5s6gpkm03s8jT8kkEkrjwDXFRQQZ7ccflEgiryyVZ3rkQ7hJ6x
1oaBepUyLQRDo6nQ2AoNPI1+UOHXMFMVAML1du6Ra/RNwgsBO+MHhXdy4nnFd42i
3JD4gto34615v/4v9Bn9FNf7NieOD4Zx5N0lJiN1dB3M7fIz4YmrueXj6PF2Jaba
jSKfTsFRrSBhRBZNmZW7A+JADeFHwWyk0wXTgwajaBDqlRVshHXW3vfCFC85y3o7
VVy6dPtKmwMULOOtpUXvLdj82orkCCTSOEe3EhOmLLXuScrw5ac4Y6ssF0HlHvuY
cm8kFtzmdWs3qNI6KBidSvbEgkqltRrN+cxN8II8AaZB+kIb2QCrliNuJl/KOozm
/0piKji8PpIFX1kx/U4N4pFQYodBmivy5OvTTda6zWMEvaRKPhmVQeKbIQafsWNF
WqaXDAbGXD8AlgpRUgfnuurc1IsKjNTjMJwjFfF3k0CMGp6h6v7rBs9bs5e5ppsI
kotWCU6nGq9vRbLHJCwJLvORA56RIdzd54g7KuWERnn98sixcSgmjdqh+dp0o05t
eVxhbvqj2oAnkVvix2a2iqfOt+9Ek5zYBAhOHdlBxcnFT0oXk++md6LWcmPK5aGv
jd+s4GyfoYlfIPvFSD22c9Y+vHEoSCf+DaeyiIkrROzLwgR7JRsTbW/FnTplZnzv
CbwzLJPYfkGXr6CTnU99k7JE8bInOtjW7xgQcz9rZ9UXQqC88qsyTJGpiOmTQh/E
sBK/YuSm1SUBdsBAFjT3bk/gaXOS8vWFqqfVmSNYX0sBp9VxtdrNSKhxeW0Ip10n
qSDkSS/yxN6s1Bue3h7GbPc8wyrG5TF4mlf11VCxAw6/XojMbnRgkljWXv8sFM6+
Uye8EyVSeFxbZCWF691xQD48H3UeIjDoCe0Q8ONjD158mUETyXQyZfPn/Ao71XjP
A00tOdquLRVeCuYeV8fqrxA6waKMAQRh46PMtKSYmQjqUfyLSCD5Idd9hkU5HYaU
m1hlh/YKfiIZdP9nAyBHE6bEzd9hZTrSS8LxNAYhtfoWGmqUmcLh+JPjFsbeiP9s
CqPV5HHAq5yVvR3tzbo/2Jpz0oTMZSFkawGhm54mi+LaOsIw6pl9cCKIcEOcwkpU
ws8q5KzzNV6VeyKOimDknodqmIlYr1mpB0QJfcvif/iZYqhm1tqKjZISJ5bmqoK7
QhcGO053cXaPpKmB+oJtcEPj0602fvXbF0tBBuqV0MlfFkUQEwDkop4cUKhcJUMo
EL9a+cSBhYS4MhgVIcbyQJXRJYGN/rDDFJq+MlUfr4nGetEZcUNK1DR/sBv6ri71
iqlsN2/8md+M2v66gycezI8Rd3+ogYiD+CS833b9yDEfovTLBwAmPX/oIZ292eOT
joM0IwqNZWm0EbetlbnUDjA/38XhMqo6/xoHxNFVlinepdfgs4mqA1GTVnya7a1X
M88tS3DMWJ1HFohWl7cLEIdToMhD6VFEo0geiDp8zuYxDhiUVPHgwcjXPoWd3C1b
ldrUsTK2E8j76AuhCm9YwmC5udlUpTc5+yfjYz8yQ79q9znV1cgcyqba+haJQXAX
8D5VQKqcxUMqJOM586PRBp21EqirFKEEtHsXp8lpYDGSeNg7/q1qhH7sazN0yn4Z
rGV/IHQPjBpFKJLEFhDS9YccmtdSuSQmWRyStGnxhJIW4WJ1uMnN25MfW4u2pO1h
7ZuV9OtZNFs90fyHgGjhfle98KaJ4uXS28m3Elc8HNenSCxqHHiRMEJoJwHIsceP
VJlmhzBXJ1jIH7XAd3Pv7scWn9fWwxyMn6FgZLI/uNdl/4V4eUV/+QsU5m0FxN+6
`protect end_protected