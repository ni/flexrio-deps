`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7152 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhBNVMbsl6PTB5/ApNH6uD+DTAl4yTWHdDqal89lO0QMs
oiUFbXcPSlFGfo4o/eaCazoUlGAb56ydabKrt9PYHeZ0YG/vO+GPFN49lAODzTTP
Sm1ZI2N4qGSTeIq1lCpXFHSkxiQXTjhJIo5EzJfBMGIQyC09moANNYglVYv2yYZ1
2tySVBA2vZe/uGdgOnQgpcHSZkGsu80Ff1jw/+gvPE6fsbWj8k0spAOLseQtr4g5
ewbC+mLZRdD281xTHa5e41Zdpxu4jPcU2v2rzberKzsObuaXSVG4gleL3jTccR+f
QgUV9mQrGziL0XIYoK5sbsImggr6Qg3y2u6CKMnFaNHhjeU5U7SeggzfV4JE6ZnV
KHAbZ8xkDJrAyi+vNQ76hBMwLoNcg0tjC2fuTTRDal0eBph7SIHLl+2wgAlYQhGD
dHQwCtKfET+ZO5ZTftb3xZB8dkQkPMgegvRC+fWJ/V6+3oPA96G8VLOayRq3LeLY
pdAi2G8jLfb0rt2f8qi0LvUbyVyr4/UDCqC9ReMwSQMReBJ05kqrB18Bo6B5Q6Dp
GbjHfjbGhsrNsq2OIONTdevGelk+WWpQmMtWZJfDPZPDDyyx/c9h9TeSWylM9GZy
9T2znaZ3xzE7DQlmBgs7ALUiU3AzRqPj0Dsl/6P4DrC1ripaqRycMz9RSVIC1flw
jfWBWOUYOf5zvRdaVB+uFb4Xwt6IGy+8D3jQoKxt7H/bahC1g+sXHFyHKKO5zkEg
5a8TR32OdsikzJxev5vbyEq3WTaR8XZIcJFljGTU1DA/DLmww6tiwI/F8egkgRdl
zcQploN5XgDuinxNHDA5T6WdFi3xNmonuAYUotyT+bDb0eHiRaeO8cRhjJ24DTXM
EX/DHJ8snnSzuTLryxE7w71+5FgyXQrYCDmrhfIlXf9+X5x0xFzQqjmSAEUtU0ss
rb5cjlvMrLjuB7sTIrYYZH9MDoR2MW2sQvVhsRsZtbpixRGlNTXY/L/Na26gNWpm
2oQv2olfVs6r5pogzLSeGfm6VJsPkGnvQD4N5O4BfDZs/nzqVr0sVGj2H4irpF6X
sf2TSi2JDFAxM0Ya9wUS7kj1rW9NTXPOp0Wqjr6+Pz1F2XesfULP2CwfZIsWqXv5
vKYmj4eN66pvj6NqeaFVvBR/1z2d1KjiquUyq2hh5tatXv1tcO5RPPfV0xJW3tE7
820hsgrygy+jUFuToK0PLKm6+z8MOuytXlYW0vaxAQByNROLI9+PJkc0TabiVzzf
inM5mQC3VrFB93CzoOvOqK/qnkbsOugyfkLfkoTqCOh0aFE6Dm+4Y8YSPDDDezEH
96GQsZ9Yc9I+SMu+AUQ8mno6ZDy02TdWaaJgY+nADG+/9dhcqTLbeM8PG83q91qQ
zh1zll2osWOrN6kL6yRfjLueMKJI4HvmHH9TQbkh4pNDDEoTdAawb9mYG/8k1SQk
8nuQz+Vub/gVulogLbyH13/W0O8cRsN4OJKSy7w1NeJlWuMh3VPyZ1EfBWY9C4jm
NLpVsG0trvOwDl0kNIoIn3CZp5XOUiqnXwC/WKOX5S00e/600qfQKuOWPcUIdlGU
TK3FX/CGLmd40wDUvoUFnUIc3+iYjw3b1Ih/1QvMJya8g7c2/8ySYLPhBPevHeRd
2UediwbJafXUUmZ7AYYSPfc1e7BkfqHCtnmkDvFYNIPXV+YWIZfaVsjoIxxLLguU
MaNI65kcOv4kqmTy4expAdLNK+F81YFQx628hzs8R2qJqUoMffJOLfe6xUeCwkfx
2xhW7yxCWvFrU2WXtCatmSd94287iCOW6r4S/UAE+7UKv+Bc7NaPJPLnS4QigTel
zIpjPCVNmRlleSlwvkVV/MZmfQJdFHKpLcgyewEJJFwb2m0onURRWRzwXOLF4kVj
CpvGOujWxh3fWcsub1eSrMuL/0sLp6fh8NnM6e8HYJBy9v9FZnnqDQQ8jldiCSsU
LfGii3bHJQ/ttYVtalSEgZUIlDIqn5dlOQw4B4cZmrIRCabRXpFW73pWOLJN8YU1
BX41+AGlp2nI0AfetHjp9yhfu6yBHaGYFETHKNuwGC54auKEm7clldlnWmDCt+Aa
TIdSa9jrnccPzX38Cvb2TqMT53MWFejI9enbrPBIdjZsPr3IkHkH9YsrT+zYon3O
2ys1V2vCfnClnUD8Pui62MQlJIBiH0/8fhi2g4e+mt2a55gEBOzwGUi6XWIz0OGv
GGzB6UnTraLwLqJHWgVMbLbQYgba/7dEXTBwnp+3r1cyO9EShi6t/OOnlLkCJ+vD
Q3c0CI7LmcwXlV0TRg/vIGD8GC234CDmc0Ym6CHYDD26IOaG8am8lTEdi4Sxuh6y
3EE660DoCQvTAvgqxmYC8dZqflqKHoSvXDkgKF1fSy9t1AdvyqY4WlG8QOrHwD2n
M7Szt5IzEMz4onKNGutXmv28sw22p7uqo2abKSb41bsYwyTvs2+s2xNOZZrKVMdd
Ilx7XC8jNhWvJZUib47lq04OIbkSuHiji4euxdnUk4ZgtUwGXuntJv4SqaoGb+aS
ddkIPgoNFGlXpMRtotB7sIXDUGw5yp64+rAcnwWL14HeYhpBmsMvMt9Xo7imJXC3
mLO3GB+BsY0lZ6fmE13bx0f3HMUJZANzRdlRB/8oKAlWsfe1s69JosQqHzpwmgVl
C7HsjPrQLhOkN5QW8ONbKnSBtCzrUuoOho+j23nwDFWjZSvfWbXwGFOahupz1ugn
CFdQ3oRurY4WuAN51bYriSfC0ZzcMQOa6HeDCR5PIWvv9oVG+4nR8Ek+arlZzU2K
21P2oF6a6MTLnyEae6Bf/qo5+OIR0qkzRb9Mwy01fm5h5aF4wqEiPBUZyJ58cEaO
CtGQF9WEbP10i5l7h6aRfxM/Mc5VwBF3a2SPyPfk+wV3O94VX+FnXp+tpizsOijB
S78HJyQC0RopI8KTBrACkSsedkRpR7wt/lL8R5n2loplCf2sXXKksj+jGTYAIRVx
K+gywCPewBSBaMZhAtsA9ZHQ4CTHE8ujohmXU5imP5wwb0/uQiQmFlIp2EdeELhV
71BWFtbq7yTl+gQ64cu3fxquJosYEZZEgj3q9V9QwE5C3THuxB4pkRnICjTLJk5u
CD2w8OmFYt2fMCukr9ZVfst4Re+VPebd+mmodSizf80bcwZPz+xrZlvrUye9savF
VjKWQLAl2HohxXXbVLA6Qa5XnexF68NnP37Hc5iU+cGE9ijE6yowJhB+DAk3b46Y
7Kc0ERDEVz4dcZ683H9Nm9z6JAm2qsgysZm4hK+JHvLjtYWlOk8W1+4am8L3T0nv
kFch6XOCA8HNu8L5AkObQjqigToDrMuBrRJUKJWmCWJOguZ7iG8MQL0V2tD5mJ0H
dmOm2mCm/hMc6bYWX/aUPFt68uYPW1JVQfQmOWyozJJ2T330axMz4fYM2A9grPq4
1te+BgWfV/WChhf2ioa6PcV/vuGYKQHhEld2NvMB1P1xGlw4ut9g0rTxDyUNLU7V
0Pho0nUPfOAlLmn0CmC8hoAmU9fQ+yUsawdNDmYBUZJ+yaBOGaXKKvxmYumX+Gpa
DRX2p7mDKzvIqE7XEhIKzYeY6kwhZ6apfWZTuw7KfvUazaT4yI0JxkfALShmNFxH
i8CNwDsYRnKauxFq5IO4TS/+g10fwnNfDglepf2HzsTAiwSW/3RT/dU3b9v71VIq
aNH77cHSy2+zEf1CiiX06Pz5n8Qzh821pJSV3BSIWpkbEfnwwT65XyquagDdgpKe
+0KlNWsTSanPf04CR0pPRkcGyddvG9eWqkAXAAWbJ17BEEos+pwmWz2/s46O9JLT
V1bKNI55OzDttgEqvgHKi2KgSQODkVirusd3OSKDMkn/qMyVXhna2iqJ+UKiQgI3
AZtzHtoeGjytl/ZakvzMQm0hooGoY1wx9+JkNUM8QJv+svue1w5j3l/DHDx1oA12
bWbrFPOclO1N8eOo/JNF64riI0soLsaG+2GJxJr1ldg3j/Rc5C9PWft+U85TJl9r
j2QTGkaFMZsHtQZK+bGuGUJVJX5f0OBlyoXwdS12EjqBoxabzUgNdCRdSOp9VoZB
akpAh/vqhvYe7/OrqyOyOfoicn3D1Zt+ooc64JeHRZOMwH9ZWksdoIKZtAUj5Xwq
bLA2LP92xti56F0E6pREGl7lbro0sUo1iy98PSrtDY5QoUHAqRo2dDmrC/bKu4Q5
LvLfW1UxHc+VJXA9BTDnBhZtkiihluiGN3ueda44HCIHzhaX5Dv0xhhq04qGdLfc
AGP3Q5hV3QrztQQRVQlxKVI6STO22720u0HhAs3pv+FiUSW+FoSIPeB2lc7BytM5
yzIV1lOlDM9as8RfOkJugIHZQvm/O7NH5Wu6Q7Rrucm4AonT776/JScD7OItU/N1
6J/LCSxuhmy3WwaL/l4uP27jBe1iOKEQTIGMtUQljcO/9DtzzRFRXl07MtLejCxR
q05P1SZJR+a1cJfTqNKE5O/YQKc7rmb7bOSAeJOg0a05hZ634YUT6aq6y6UcY6zI
0ecYHTd2fBMZc6e31HYsuwL9usCteCH5eRffRxfvOr3yniFPqJEoR9piG7aB8HhN
xsY1sLd93ZhAlXu6Rm0l7XfX5OBGo/6sK+8ZGNG/Fs6voVUDKIS2bAGXnWDBVmG2
Pp4ph4MsrxZchGdC9PjNFUKJeiSpPR2SdWobodTavCl9DoqezE24jidqexT+q7Wz
UgzgX9I0SRQx5jO8A4oyTUcmHsGXMVa7kIiv+zvXw5fiIt0HaXL1c6VXC9W+0OSX
hgjjnHswh/wv/Fu0Y5SR5cOceR7OBLQkIajOWUhJhvGHsfd+h/KwIsmfgmSeUdrF
EoiapKWFn0nF1+zK+t42Q9zEBcOa5QUHPO4WNJT621ipIvGBynNdWU0j6JnOj9Fw
lysiZkd7614DB0Y1LwOHpfE6X7ud9tcp1QF0fTzutSa1pIOx1YrZ7fOPriqe1HXK
+T3tfcMdSwdkDnYmTFO4jp3iqQbmKGe/iK1Yfe7G/q4PbR7/hXvvLGLqZ4m/2a2k
CD9TPNNBQrxqVCvZ1TN+t8GIzAXYjALFe37zWtvy9mWJ47YtQXPsvLXE1aKyf+Sy
nUfUvn8ESZgzsBrStBI5FiiMzUSFrlYC0DxmdvSgWW2aw6zLdcmce2jydg+VtGLR
SgwoEGKrv9eH0Kk21oQqilSHSSAIAfY5YpJ2E9/qAG9lpUVYWjfYqiw171C10sBG
TX2WrE8sAD6NjvL1PWSiSqVMbfb/FlbZfgiVg2vSBPld7klciJ1QrmsZ8nHPMkM+
VE7o4bmTtKH6SlYBMhsiJ805D62F0USakEicw3/7C710/KspU5JjlDYQQKC65bUv
OQA1/WCpOSMax9XV0uOS9pqZbppdDvHi0zA1Pr5LaaoelnWP5moE79E0XlGD33Ep
92RXLrNDJBkCPAjpQHcxHmTnaM5vI2/7T7ihIi1Yc7pgoJQuRq0ZO4BoaygnsT7F
q3MlTFCXDfUa+u7LHENnXViFIVT2dc8KdMaCgWXN06JO2e2NoroXlOVHhXvYe2wk
DsmFgPvxgErzql/SR4cds1rcv/ljKedlxe9x25+ReqXRJWIqH4qOwfAt/FzXlSjp
gBbNYWyhKDiGJWQUblkttlqd6mGI2Argl2h93pbf0WcWGVeuZNsQ8wRw5s+lfILl
GWPf+kd6cIfSAQ4U/Und8mtowhw/XXyevnwkGBjFZ9lkLe4NqwiLKRpy7659w4n4
UsY+Flz5REEPtqY/ZZmTq79Mk+i47DHwXN/hPOGceSamJRF1WYEM1ctiHc3lHE4v
E8oEEUcQ6Qa7jfwssTjqjWGcNDgnx3b8WAhGosKu7eDL88Y/iOZejU+r6h0KJdkn
bnoQ+lboRUavbowU1iEKbmZu3Bt3eMZ5kQiP32iIs0HNfezwiGx1dhXjk7Ea7EQr
7j/yqKhJRP1DS430tAZbnJq5JmNiOhjvGgEIKQT5HfG7hW7nmgPeh39WcnD8WoGr
Xx2EN4VAFtMsmRBPqbUTEsjZ/AhvDIa4tT4ROzpsQlzZyLVmDMJArpLPPZwKnlCY
92kzRwc5n3Kun/a5ubDd+IThGuAldZqqded7i9Q0jVRiT+SyHxdo3f1pD8W5X1tF
8oVMdJYv9uapCjN5GhujZfw5z5stiOI6vxFGZVi4F3mj8JgAK5atc6QJXz6oTD5v
m7h1tOzxs4JE4dKZxiZFaNzpYoH5eUjoGMOE+mdlfc/iHCOWCRV36pz+KWDk+hwk
t3FWNs9PINKfXiFEuD3uIpAH5cI8dWPBwvAiRClBsZmWg5XgD4Nc8356yM6584JY
QPcKDTei6/kmKoLHH40+AODqMg20eT/lHCiKJBx5ItMVgK9wDSYm3EpY+oJyXyO6
4FyapFp8Sz5ZmdrGQSMtZKinL4jihIbjwQr7H3UiE8XzfcN/R5jcisOKtI8Mzmvi
6g06i9B2tfqoaa3mer6rgxsDADiNhN8mBNBj9iJSlLme/kckkc2v/43aBygVvMtU
kdWopZcnXS9mblhJEl6GvSAO2ovflP7tefeApyusJw+cuuGJ0mh9r9m0uaLTtzWd
/UBgdraFZnYW0Rj4GHxMOYeeh/vSRUQwTrGaBnd9fA20CLEgazowS6J6VHAC5Mok
JpM83OYymHdc+hhWnJVDJZ0tPMX7KIg/ogleoyj8plPgFfLZvcevNs/uKB29dWg9
4Y+0QL5BxagRd004LoNWTPE2v7X8G26P1bQDA6VlxPgrciwCjaUGwzD/mvkmfo28
vDDXpxqeT+oTVqpVOVbXzn/CbwXRK+1fdLT4yq6SGfkP31X3rbkltUoiku5QaIV/
oJXAwb/lGTIBtlxOLTh346h9XX3H+Pnon9glWtYSRqF+ApM0YmohtwjTlNfjITwY
G00udf5Z1IDvv3GEIiRUrilM7CCmmVx4B/qINzrNC5UnqC7GlA0nAQdTiojbEZfr
5cWhrX/C58+NHsvjwcyr/uea/vYFIEZV6TvwBhhxXCr/3V4F/+gkPe4UdFidajak
AEHBrQ9kOf8RjKaCcPdDfUg+9hyJbz+J8+VxR5Sd0v6MYnmNd3ppss5bYhKaiE9s
WYGPC9vbiHKJpi8Mcv+91zeLiBuNosz1zD6ynXMxVZ3IrWKS6VVoPffSBxgNFsrr
53oZeVVmgkqkHdMI6HImfELs8fW1A/lJaYJjeNGLn7qZYnwhS/ojMCNOZf8IVfmg
iTyqAuPaP4MBTLzqkjxe36d6Cuekkp3cWTVUbucHdDZNLTHxZR4rTuygDzE+ZN90
lPit9sHgNthwCohR7LgyQ+LVOimt8oAcruckrh0PiKFXkDzeNTKgYI63kCA7klbL
fmD0GXZ+qAOaNP+OokmwWf6MCLci38tuTyzx91H0mHyDbm9LNRnC2jzA2CkLnIfH
jYooo98yJS2Vx/k8UXEVemkYtsgE/ahW1oAh6VXxWv682EFGnvQLBeGKbm+UsUSE
ZI8ARA4I2wNm7e7ZL2H4FJ0F7Oef2jLVBfF2JuXjdIUj6gNO1PRsK995VHSCia0E
854T7BD3Js+Q6VrQKnKtH7URn3DDtDp+YtF2bCc/BSn96WzqwsDMbj9QcGUv1oqq
wtx+E6obwp/in5kPZLyFgbDF4Gef6ZjnCDvebr5aPDAxmyCmMWqqW0tVVlvfeMOX
a40le2McjIiBq5FMSrmoVAIbWR685v/1552q+Wd5bblUcDnCZzyJupRVCXXLB9g2
v8HbxxyRk737VjMsOgAMBxrn9ohVsn6OpfiGzU5whue+FX0BsoDEipGYDFJxRW6x
OiVIc6JeLQLUkMUgQypxPEFfBufaIjfS/FyLw4UB87E7JswxuYL/B/YycQKnPUPv
pR569n3XNngho7KDQQLfWTGXJQn97ze/ksADkNc3uXhMGh1RDVCZKWWHxmGtVrgS
Z6BG9RtldBdYYKjDZIgqgPXhXqHikL4m4TnmXMsz4oDOuK6WjM8fbg9kMG5JdVvP
E11iUkLP0ZrxkrTCSruE/74gGMNnaUMQ2uk16jL8mOCeGa943tPtQc8tJNxlG/vE
Lr52RX4e6vMezFQ5/BqWXbaNLwe1qPq916kiIu/ZP29cWp9BHkITCD2voViddKrB
dV3UjfaIPbdTjFr7N21zeVWwztzTy1fZHCBbrONsOUn91pxQ7OmdgMwVFCx46QKA
2yI3qRKf4I+EosHvhkCpE5lbaTT7yxY0yFu75+ptuSu/5LZ29+qDNi9N/FzqW77P
buLx4K8MglVLMXc7xDV/fbOJSiVVSruxrg90BXUtowIjdO7Ri20vR889/ISXeE0i
nE4tI06VsazHHkyIBQG3+BhZ+ZKUm4k3Q40ScvOmkj+VKQ8FtMIBZePVAJFJ7TqI
6atYM4/eLgL1BZVI+ZPtiszvf+S42UA9dC5mSElER/3aq+CDFsSzp1hZt3f0/GYR
qbBUKrB9ZRSvZsA+wV5s56bahvJkJKab12RXe4g7tjoynG5z20zUFw1GDrOgX4Aw
ZiJI77awiU/Qwij6y9sdbjWTShsdjXuNOH54WEnhZickUzrF8l9l2B+3BdC6tyAj
f6l+ALttdRle0zDqfv0iN79T9d80x0hZHcaxezMX96EIferB0HLJlHKdH5oDqVKX
NEDidSiYgLUFOS0S+qeo/LNagsMKt5tIdmYepg4kkyE2mN2i85MYsspPJKE1BrIJ
dR+hgDsOdXvmgEWGSftxRR37tmL60YbtMYfE65IFQtW834wxwNgNbSvfHaNfKWIo
xZyjrT2jHofQZc2kgobAx3T9kNvqEebFJ2gXa8lXB3zyj/J+O1Exsz+U8Oq2u5HW
jGrzsRog94W9Z5cGyCoDW/7fH1oPmCwjc2PMFqp89d2P8VGhlxgPXW8nXFtrEjPJ
njhuPe7JHMwIqhyaYAh3kq9O4SwEoC/PBCEdWkfMLyteWe01i1z0O7/GFTHdR2Bc
TmUCkEo1tyiKvUpb4PRyf785X8tao0lOYzZlKCW7S6OPpJUNROlQ//6rQIUfu3Ds
mK1Jjzy6QvNhVBweqKHaKzXdOyExJzejRkm83ItyQ1SHqlJ02o0PSOqYnTLxvKhs
vYguaB2iUTnq+UupiyjGt5Ow0eZI6kbvjRFDV+uJ/J7Je78mvdnWxcF0S/35KPSM
//ek+6LzxDpzt+eZyu6gOo8rN2Arbez0R4Hxu5tcDQYjYbQ51o4v5bsE1PX4JxWQ
JpfBAC+GhxgItwfAXevsuonnVnusCQ89PU/9aSjromAcpAaCMpLV2LYZ6uDvIZ0p
OpE7PSTsgrKdQjYsKGkyIfjs2bwKRvwVsJs1DNZ6XpxXZuQ58XgN3fMqenyYxemZ
NbmfNQ4xbL/hIDfAXpFiyG6w8M3aoVlhbFXn/7Q7+COxOe8P4tzVtM7as5Xk5UfP
`protect end_protected