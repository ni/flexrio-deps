`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
9GNfeu2LhBO1rvG6TqMSwN9DfQJ1HnYmA/jtJYetUEPPvZj7Hlo43NXEQRfOVHCB
DItTg6zV4FlXnCh8U8uYgajGPOQu4Q2Y6a8BeUOmC4CY1iIkK515IdllESVIZvVc
2/fPwCLv3WCwBIYHV9uu0CgoY263HeDKBLRQSSdMBo9kVroW5YeU4BoOwufsDRyX
SNcRNMQDNiA6g6wLHGRXqROWSkEsY4ZQFLPu5WzEdaQD6xyQylRDTHCIOPHNOWMn
nAYhZeUmww4GM2hwShnb8Zv9z21qMn0/a+pouKIv7wENX0vPYnxOyeiy1WEbp9C8
TO7BiQbIbpmhOAu5sAF4sB2QTmRH14m0YRwvzqq5z72tnepTTX+jfXGw4eV/PwH6
Czu6+CFzhGC2Vjy42UAWlAvwD400YW1KJHcHtQCpSU4HrLIri6ysbhBGFosYPZR9
Zwe0owyxwKSrxbOSQbChKTBIKB/5EBjz6rvOSwHm0+yjNxmX4JxVrg53rdYImPqd
6AqpjUi3EnjNt+ZK3et4CvoU2R8LhOnsT0pd2RKYKTBTVLQRMxA3Wv+P3QeWhhKD
Dq4OoYTKyEBA6qTC7zBvuLSyBVfaxM4D6BbQjv9545LXDsq6mBMCNSB/F2hYZNVK
T3ibgl86uVJbG1474nFZK4xUTIk9opNLNndpHR797CkFm9PGbz99Oq6jptCq6COS
Y3qojcSTZJ/gTPQBdmU5uh7b2bar1ktDxagvCEmEhU0OnciodzzcgeQSxILAc3rG
IOaxSc/EG2p47U4RQWVYu1tc+f5pSbWQkYCrSGgzgwYJw6dCxqMGAQlBKeM6Piox
866I//ZVWVS1qxyerCTD0zHNBeqONctXI4n3J+HcNb9llyQsZsDMrQkK15yg7DYp
LagJUsdzwpxvDb/kK0Ug7nwEGBEQf4a0iOolWk1GzGPcd9xJ+W8URJfRZ52zrImZ
X7sN3zFMIqi/g3OlW0Mu0KM3FVIr84g5pf7K9hNYomw8CxFBoEzG5upa7dhDmA7A
xlEixvWKc+qvhpooxxNKp+wnp989a11V4Y8PLXLy9O/FpBRcyT/BZt7JjgOVticT
1xtv25RSjZfwiGPtY+6a5oEZHnz0OAOQytC6/879tm2XAi2xqPkzcK4vWO+sHR4k
xMW1dw1Z1vNO+pYcWdbV5xW6HRQhEeVqqEaGIp1D6Di2li7hY9wAN5Pn0rFLnbWg
+yV04mY4+aOgoB3lQPHKVBGKyxU5i8GSEGlIIHn0uPTJNoEiPiNiBPVe+omj8fKW
WrElxAz33WQz1RCyoOlkCDHqZzaD37Kh0+Y9XvfT4FfgJYIiAtAV+Ua402SkMVaM
4h4ov2WJ9VqLH9gk0eSMn6YlZbBjjhvBC8aWWHbB28LNNVC9bttJErGGx1S+yKpO
jTf0KC9qomD/bY/OOIacHi9hxWgsamN87kWf0dSXOJL+BbTGWCwEJrrcP+otp6t2
Vg/BijXB9T57BTBMFPU4/4QSW5AQDaiZdlA+zJ13VUJJXCOZ6aEx1wOZn3LKEIHf
E0TXr3ELGhEtdBgO54CpTqneM3nRLvq9/fYDpQeHwjCcJDmbPYNhBzSnvSXnUkJE
nKA2LespFUTej3kY9WKEPLKKdJ5pvfMJw1P+AWw1uRbsnczKe9C3XxSMlTKYKcEN
n2TlURw9CGTFbTqpIUOufJ0SfXNKlnfI31WBe3Ui7pOytaH2gzYOdVamUIX55Sol
uf3NDUcWr36lpCA8hfyyVsyiiPDWoKkKcHL3NoqxZzDk6cETSgnMn8oEqNJrnPzA
B0ZaQQUBq752+MVZMKyzjOgZ1gzLOVjlbbx+XX91Htc3WozCvklhB3bJ60Xo2pby
3bHNzhDc5KdYdfeqPg8Ydz3VHsQf1evtipjSjXXG8yoG5pQGheAOsufSuJ2m62ju
BtPk3OT2bicYLh5nBZKERTaMogOhkHlnPlv75SVPpFyCeGuJ+IcZ9KsQlpivhI0p
WXxrInFmxtggkaBbuFtD+Ov5aZMW/8TF0jNe9HBT2ewzZXKWx1L4ssvF6ijtVG1e
WLwKplD6ttLOtOMM54GC338kfwxG019fZdsH4PiLkJOxBgw68vqkP8yPltA1BVFy
iHSS4C4bb9rgrKBIyv+3CKbiFZqTUTj/AfUxMcKvoRYVwwXYkJRQVNDAAeClfoIz
tFPZLFeuMPPQXjvE4pZXm6F1yvs6I74tAEmCUmG3YRfubRljfU7jAD26jUH91XEj
z+j/MwbzfOk0oXDkfeMfBhJFgYGzN+8GfJdJnC7UM3/Dt10HGA6FRLqlrCYfdVF9
/1kFMBYxjyp0SS50wRSkaJkdV4QZOcCLt5BxHBq+JsA/aJyCglKLAv+P5S/EyH5H
QHwzg1GW08DMcyuQ9Nwn6hBWWA7Jj5InSw/h4kJgijxdSZAHnF5QgsZ9k9kqlkAe
UL6YGG0iz6KKkR8cHB2tOLXd9VBOG3A5fVVGto0lFIkGJ879tnnCSDh6G5HAIGKn
wrkNpQGnfld67U9/7w9IUUl5+CTLmtH2+cUHXPv5IxpO4TMLtnt/EYIeSJZ+crua
`protect end_protected