`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3792 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
2n+M/KhW/CoPvt8soGKLVoD89v1NVph8mFe8lvpp5FPMTimESpgtc1VLPu2C1dcu
fQYk8LNsoDlb6zcNF6OxbmC72yBx0vCj8GDKdpd+FchFBxF9J215hSq1Ku2Ait/3
pL+jh+ZqQ8RIuPZBzCzIvhjtvc8COxU3s3bpWck4Wj4hYp/dcO4kgOZcJH4xZMGm
VHkmfSmVKc+5Qss3rZfaHWUOrXT4yRm5THAQYJtvDKp3wv6QY8sUlQNC4fQ/+unp
OMmPMoh1hyCbBDkbrY+clBHwZuW1kAPolzESpGKsu03uIzqTr0DdaevGgovLLgds
oprJYKQD8V+MnmFz6xsKJJd+b/5A1/OQyubF/Pof9jj+0WX12xlgx6AXXsn8f+Tv
ug1l6tm/25pvM0o1ft6gKThJpQQ6qirdqgoJKOch/OO0sOuDUImvSLJhQEbxo1UY
bd0alZDmSmRugLHnMW0c0EoMZ56ILror6klWrVSxKy09PJwT4J7G47BKultjgAsl
Ugs7xqyMGfli3NTeht0IxVijEWgXIonox/6DGRmlmjzfnbbY9d048j37Luvel8O+
1I9o8BlqhoS4DUhfLGxlTmzwxnn0HokJ5NTV9ptIg0Vp3HeYe2trrUe4BpYCDysE
i41X9hSgYqu3A7b55+/QQZbjMsPosyBDx1ZHm6fPrc7+O1w17Fn+T0B4WJ+YrR++
J4O8X2Xmx68zxguvCfXY7l96LgrWGrxIFzQISQxvFXHHrQAW8fT9/t5uj5m3WMHk
P10zDzoL/n7HwQJq05+ZTdcJJlCXe2xO0NUxOeEs4e6oDc1tkXlWMOP5Z4O724IO
bkHGH39iWm4jp+V/nIaeZViK+VB+bqoVRaEVsxyl8U53ZF8GSVf9SQAHFwjF9PP5
/iQ8rbA+VbpbQXckqxaOJM+ofLluZcobnbOniYydF83qpgkpXLENp1MVDtsHTs9s
gq9HABjM4UDIUJSIoHx6EggSdMRYktKPGelZAGnKMdaV/TOP7vhgYINISXzsnXlB
V/UKVG8xS2le5mtp/sioYGtBKst/34OkHvy85ukvKB2ES/3JMGmQD+b4CbMVb6Fm
+seMISGL4wsAxiP3q0BDkrhjzU0i5XWD4k8MP4lv3zlImI7KmnJ0yd9RruyMx66x
/5mLxmmUsKIFVtHqI2h/xIKUXd0JNWSBl2yXCHBGpC7fE8RagmSb76oV26Wsq3iE
fpRcevtFlOKpBVDyWj3jFrJZc0pEWBuq9nlALTkiFjmsKkIsT1pWAz/Ditj2JTcT
1gIyp66dEvorhcYCntvQ9NS1tUrGXjE4tnZcL/FwuN7bw067i92XXDhYurfufWQQ
upVIegkzAqu+KTIl+TlHnEUf2MgoRiI/CiHHbEgoamZ20Y+yHThQNPNR5hvCgQ29
djXRQcWp1aUMm/y0q++/LSc9yZP1T9XSJhHUEwO7YjreHHDJ0rKY0rTJgf9Fg4Cj
i2lu6ivqqHuIcDjq6t9o44YDUxLICvdFGDZ84bJUakKkmMUu84oDPayY6VBuXOPp
mQfdT/ni8kRkUwzPKq3vY6Ni7wZ9RhgZMyu2dFyK3ykh5z99cQVSXAouJFXwcuEn
y/4D+AAWoRYGfxe/JyFFeYjftz01BxncH5Sj49AI5/ltU/J6uWboGchP2RZPRLYG
ywkWM2u0T6xOoEL4UfoB0P6E+ppcepmQFkzdJ+HiVsUVcd7OO1SB2p6/0jTdj2Vi
tVT/Y6KxQDCrswf/isWkqCU8j8Zx+5qXXfzlCPc6ihn4donqXharuJCzRuDj5NEd
BQ9EB/NkbF8cv8Z6EvHih3hK5uBA20SPb2qC6k0oyhw2vsTOJq6pnvT+q6QuuBPA
uaaAo4g/Ar5BmF60JxZjVJ9gR2FtO0xv/bsmV2xggsFVsWaV66boGj/964v69qPO
XvHnSTiTF56rNFqWni/3vb9yvOAAH1MIUc/kuvmDaPYj+ARd5YwurNqqmP6R39PH
QG5rHgAD53xsrnGdQaKD7YQWIb5rBUDkltbKyDRs1+CTy/VxhjB9AHVdwZRQ0OBS
ReBTJ1GpwFkDiWBjt11PN/T7qAm2GZJLM04JCs5XrE/psVveqjFCBcoC2qTB05rS
hf37nVDKL6Lmoq+/KrFy0Sb8Aptm6WprfF39fPcq85hzo8DZJjx+grzdXUnNT4Rd
jGWS9YuOzH74jwPFSSeNZYc2IxIyOKhD+cw8CJbdvoYTAx/yHcVcRUZ1rhMVOZzK
P5l8CR78+6vURUVx2Zs6ZKGxb+KhnidKAU/VRG8tEc3M3ypi6QAQvgSxkQB0nMWB
TtjRYo/dVSlDJURdh6oZo03/Vp0QsLcic76uXr8NKYSz8wcUr2S4fuhU1XT12p5x
8Wy2DCL3LdL4UBUo7imkA7OgD1pWbgxKiH6naEYTffKs/CIH6xOjytK7xtzdnA7I
9DiBtLMEP3H9RU+bgAE2CBFEhhRvgWHvE7Ei0FdWof9qMfdS+6EZTnCorAebUShH
mdV3SrfzmPqFWF2wjTARhtusdhPFEXl388GoA295BFJB2NBJ9oVEeuvkkltiTxJ0
FGtxeFTpAyHGBDWvAN8ftn2uviK8fABpwUX3k1QiPxFpzi3PDDWo9XhmQFZ3Z4St
/ZyboFu/lHqJJ58lf6no6gKaU7EKoTIiK6ecE6m5VQhSdWOY2zBdn5su57Bpd/2M
fmwV5ZU/Jzr2SoJhCSikYLwEqNkpqMPF2Tvr1hCQ8YR/tG5BM2wzfKa9qabM/lNN
2d0wjQ8xdM3KVZSLOOeis9mvTU2f6QLpJNpVHer9ZcpvwZ/dLg0mJlTYm8u1ac9U
8j5TnZUXC3hyjIUwbec7+z/6eBEHgAEEhp7GNFCc2+OyjPdlKz8Dr/hnY7mqp3CU
2YeJAznU4X+4v1ZEzFTC4zwizlBaiM6Ps843N8/+L6EAAsLDlGJcNuOvdk+QYTod
pjFO2sXQsA/XJUjLsYtaJiYpED2GMdd6jlmBQvtD78CWU/KLb0ajEclLQe/65zja
ZMPXy53YBmWjYSZcCin+Ad94ZbgE4J/7pPfV+YWppH0XEviUW05zyjK2V0vDuguY
CMVBz6tNLZhUwWfEUAzrh2geb3KRw51V5nrIeITwPLDZFt5pJf9aL7MX0rNsBpZT
8t0BlocDS5WWDj+z7ghwLTz/GbGNPjAkDlJt9fjNXa9R5L6F9zPPS6+mMBDypn3O
+2AwD3sQWzJm4g3DK3PygKSXyEl5haBZd6IGGbRJHmgI/7fqdBSsHSovxuZ9mODM
NGWyYLuTO9t7ZidgmFl7HZJC4bZUbzYfqIAPz8W4sTnOxyN6OYX0JuH8Mny04inP
7fA6flSvbWSqMFmVfbhfSFSknhGCzWFzpkAqVX3QVkgEkhlMx+r84aZCeQcC6A3t
mc1nFd2582JXJ6/K7ASnydgtxhgmzjfFqyOGZcYa/twfHNXwsU6STmv9vDf15GGb
hiUvGvCoIQRaq+mRIdY2ofVXMbuf9HkimimZCKRqONyFGA0y8taMcNQcEl1E+hG5
mo5hK0IsSHdMiWsRgIAHXQd8UHT94WjCLmhsiWxmdLJ2EhPOQSSNKE5BgN5ZZ0g+
g3p1Qa6J1ql/RL5TDoo7aFoClhlKtORV50nisQPMOxfhCnc4yyNJdgo95+70gaDe
lySLEeA1Qu4ZMlt3ZN1HBL2AnK9+30pU4cIc4FgoNVmNSArkrxaIbHKPS6zdUMVB
kgMhAI/4jhc6ssVr9aJol2ESliBqNScv5gRzaynjQOaDhqxJPVrxT0W8wEza+9vE
Be+4gDs1a1Ki2KPHhM/mzMZ/Jall8TL+TWPjzUtfYJl2mJKbz4ZmJeM8e/76lCSA
s34n/u65kg40B1NnJUtARa3JoebOxqZPcJs5BQ/AU9hopZRLkhYo+bY2R3Idw/LS
mv3IJ+aLOJEupZLzEgvoq8fu4+qDv4fAl6C4C5/8IIp0DNCcbpK2I1YuCWh8Ckg+
y3Ph/lcQ/wVCxls8efZfFBD6SG0XNC2IZJxKvyuk8yPZhZ77J+aA+AjLi1idbwAY
rkx+2fHHvg1n/PDjxTPPkDnBjPz+WFYvpPWcwwE9wu+ApvTIAmCPCKUxxMurUlv6
pzD23yCUSAj7+ypDRns52cqEBi4CGF82E9qCXE+xx+XGFGbJvTduWkzaAU1GfNsS
eSiVmD+7OaE2v8fI4LAWzsXd+vbHa62cDqcwXgdFKbOO5vrbxfqil/0Z4mJjTPfu
yG3imCuaH+mv+HUDFEnuBKqHI8Ggaq3JE3xicMJBxI5xmNVp6NNlgUrIh0hEPDEY
6VQe3xpWODdDlalqVwTfWAigOZv2/e9lCj6751czn03/B7Uxpm86Wzp254HUS6Nn
9Wh70xqDevI7lFbisBUFQG9ko4wkHjKHTC3KobKDDJjzPUXRVJRL6fwhNx4i07lp
pTttpjJWmPtB9czzLA1bxjyTgWNKvDVz4lKeVuQ0GHZ1Z6b/pQFRIxFZBwLjdvrx
1Uyy7vUBfuYnOmFHoT7ieUivjrqDja+Ah2595nOZOzfIa9kSJy2DyWv/ZaW2SfRh
hd+oDyVPqGMd7cFoEyltlQNDSc1g8/mv2kbpjGIigegM+AqCVmwhRy2h9xfzwRhP
1uaA4h/Z4O9sibkYRoglrfwxpMGyq1NLj88ytEqa08gvDxjx4UoKfois1Z8cSjYf
AEbW5mKG3aTcUyF8ydvaxFLoqkN8GP0WvTpiALQb04hdpnb3CeEcasx1Oxye5BOI
e7kWQ24RArHwnjsQwkEFE56rPHaKYq9p/NP4jdSDV7mCEOHpQutUooDovXqACJWk
CKbjIW102zfR3Clwbx0eEyRWzpGdzelOix89Ye58/lW3t2VtFDG2mDqO8X1La8cG
O/HxieR4i3NdfFQTVVZYOwTdf/RYapqWGBFLMm6n66jCIJUgaulPI3jE0+Dx0aeZ
`protect end_protected