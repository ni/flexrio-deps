`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 27696 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4sSkgcOrtFFGmnZEnVbxgx
+l/NC0KUoptgPj67g1Rb63m5dvfkhH6v1K26/83I1fvTrMh6ed2Z7LoWJnzzU1Eg
CpbUSz1900qCk4MmvIt0zID7Jl2UuZP0LpgMhAL72oecVPZ6shGND+Re86CWT0Os
btSEJ7flLp3tm/sSEPVc/kc+xMABl2fytzRzrGUg6azUodGp74kRgB/1KV/AQYSr
ff31JK8tjqY7iJ73/6DwCvouLqNEMlMYbSB+kLhyJC/Trj7XJZdeq7Zu+d1W5bOn
j0SYozJIOkxPv1mKQ2BE6QS4iqhA5KhSx9a7K4uSrgKN7CVX4wUzzteGW1yi/Iw2
ymzrRI2ovKUK6YE/GtimwL+sDKI5VXTFpcZElom6hGlpUFdwNBJdziqVLUEpB0DU
n0zZuXD3HALzvA5cHeXEMXEgwVvBqtOhxrhhv69aY2UzU9M1BJ34z1tOJ0jr/Jr9
/dLaSq/P6As85gzmJDb5KjeawK4jvfgV+AsS2HEEkOYZjahN5R2hdHNXMhGc29/o
bUev9gHzTm/ujs3kX9ASUUs8i8eOArSM2vjfJ+nfRynZNdZpQR5+gtHuxfOlA63U
reWt+31WbONmCbNmEZ58Dx7yRIm4qi9t+r2Ss0hFBzmvaTxvNMg9h2IG4/wzubVE
ZLZHQzjNC+aPqWCxUp2ngfzBdZm5Y/UumpoyXKIvTezadEWIK9Gi1OkBoJhkHPev
C3Ga1RqJi69NtFLZfuWRmYJvU35H1MQRrbriVNBB1wMVyBNGmLn8aFUxhAsg8EbO
7JrUC6jLUHr6CSfh1mJRgx1XjDmBqrS8mw0b/TZDqXQZXTHNC5Z/zm+LW9xPTV0J
pGkZubhmkDk81H8d14yG1YatfdyUeIy8ZaM86l5Lwfp7/gQxr9gqRUv58vbYxNnd
r6UsaKpctTRzF65UKfrfArlUFJxwQeGqZq1DP0EGR9apwSbR7PSvOSFY1OqSXiXD
vf1BHdgamx5INGjzox+u/IDxxP2opTVtSoSnN2jCtt8bxmBNXibuoWyrPkfDt2AX
yhfeh8WahjfqpAxPXY+LLb1EpoBbIDWIX4yA6uk7IU4M4Sc4UsPfg00v7GKMZNz3
ge+m3EuT7om7DTX+ny7zsYtIS65Ax+2p7swOLSl+5tqTLy7DscXoLHo0NaXphI+n
LNRrmhU1vNbU29CNz66rp1QyXqDYB/3STWZrKXC8EZkegrhj4QpQ5xbaF04sR5tC
jzowhMaXKDulfrMZSzi7zPJuWyRUOQQOQlZg2J2tiTurbQjoMAvC/bkESIsWZPSi
Y9mxc2Hznc0JjXvMBqF1fupjAyKZLcKmAyc2iL0rOf9H2CVKUvki7V1BlhgnHoK4
ngxvSHh4R4TtUlTLUOQyiHsn4tX+zWg2jt8UvUtqVWtA+u8VfFDRZqaSwOaHI6hB
WNz4fDAr6/8TMYcOz7DPURHbCvlIt76pKUwVPB4Zda9jWMNWeZWTHSfrQN0Hb5FM
eVsnQN16JBIuupUi24tdaTS395DH/kAyFJI+aVA3t8kOHMxxEahxkWtzz9rM2jrn
pw0iZv8vgNyMuNSPgKJp73AOvvTj1TXrfIoQvphjwEBHdHmn4u5VWTG8JJMHoA/S
aTxZ4D0/n10A6ViLD+nJxmGXMHqyM9m6JCrYcgLftYLWWWKSjS5XqxLEPI2Z4ZYY
pu+zIy3PEqZ69L1uabbpXEiPOaN61oQZ54CY/H+CHLrkUTH+opHaXen2h3eHcSzx
/14YuEbD9Y7p9t/7HdAmWtgPm9m/fOf9UqdgYbBIVsiQaQN+TpnFG2asiL3/5naN
dcds7GtiVteQWGviKrw0cUmZuVohkespUdU98TjTJ1SREJmlTBlsM96D4aemPeK4
bZSrSkZtVRyvo5E7HuSt17vKL4ksYgD44gchcpXeNjCdgoZIK4OLDZQFJcn8IInv
wst1J+n5Jbl3Xe+OtJbGFtTerYh9dm71tYz5bQ6UUDXiz7qKdmzD9LWcHz7sH9gY
dvoeo7m5Q8QKs0opaPgZUZSPxqgU99cEZemvx0s+QYLsfAyfDXu1+f25DW7Zicbp
dK9owJRlnNCN28nGRcMOLTHvi/luM7a/mLShh8fA4IT3dv/gq/QrCfcKeCWcXMzb
GgFEI2aa/aYsTzi0z5KyUZ6F907/C6fD3gja8sCa+PBZiqK0d9Ck3LiByQVQVPSQ
kRiIK68hc1jT2dopIabSXD8zFFzPfUWNqhO7FQlfdyjHUedbEPNcm1PCHKt9vjTt
IHagppFCdtPirO+oqq/pllAtIeCzj+Bd4YlX4nM9U0UGxfLEUgERWPNEXOp6O3rL
fGUcNx/lnma5PoS83Mi6Dv5n6GWT8gni/8Gk+sbu52JNn+bB1TvSCt5DTfrX1THo
S4B30dBMd+SerJwTxGA76fE4Xez88GD5Qt+vDfOV6AG2n4TIPiKvtCl1V5KCSPOd
M+C2t8jT5GTGqWlBZsNF78MOYKa44BfpHK5FENQSziJdE5IFhSTQUojHzuPgmCSg
wiOKEZ00EOJkT1i73vk2FOXLZx55Ec4n80gHAMqa+V1QEvB7ojMEQSWZLwY0XeCi
D+WeIv7S6EmtSvm+jWKy90+zHg9BtCtmLfBdwTiUZACrA1wFAbuNIKMRH2uz9NYZ
zJ/uzSe4RxOW0P2bmSksEb/Wp6RKw1pA9M1cibNqjg8Z72U8n8FzDfQhj2V+IIGL
Ni5OXkHA4kpDMxI+2Z5gBBMW/4BzxW37IqDlAy2TkyL8urq0PSaWa7IENKxRKAPJ
m3Lga6A+vUUzzLWDOR38xR+13f57v/6sNT8VknLZZiK5xR1SFLpbcLzF2EhR9OxW
OEmjPcJv7cn6lThhQMVuPs1lSI2wM8XMnCk0+cQXitz38gIERVbuHIUpc9RN7qAw
nwHlrToJfbgaUMWPqhux0uajCjeX4wO95ftOoecnG8cIPhhK2SYRp+yrtLFxQzI9
v//ksc7F7QtSyw2eVv/gnHefXxDLrl08p4/cjb+jGasqcLftRvpR9HF17H4Xqq16
Kd7kLK1U9TpDDuMlvzab1yK3KdYezGyxp7kBq4GaXvBCw2GLJ9EDyosFbQpznacA
II6ZeHY9QSg9hHpoXP9pFexeC/iI4SVIOU7jlp9TTXUgr8xKWr2G1F3czxr8MhP2
5PRlYRc9NEZ32teFkqc/csd8et/aFz4phw4UmH5yiQzSOzyMsErpKWEoiWBy0rbo
a2bZLBJVTzPJVGT6f9F69Oe3AJAPeKc3SglA3mnvwFWsgFrC3s+clCmzGMqEkV/E
vHgR5RSyswLQrmw7OwbxsY9mGi6/ywEMCMvWCNBsfjvCTru0PGTnsMnwKwPL9+WG
9E0iAwlchl/FwpCOxwWCHcEwurNsWQgkPPZcaBuWxE80nzWCLul7UBouIrw5kMN9
Ze7lgn1Cv1x/DZGbkJcX55Sfix+ss8yLLQqJ470wp4BpiH1o6ByQA1SJHpvWriAa
oT2Y+9s8/CKByQEdgD54j/1Thxh22q13iGsJ9Wy6TNOCZ7vhBM2w5K8W1RsPUhEQ
3CcwuNHBiB+eIa5QfQBHjyNvDoQq8HfBXuGvfpD0RRoLYEcoBNgg0MSBDSqBi73p
pMStUDtHD+tl4Aq/4xYwGeyqV+c9KBQiUhaf4sRybLWbu28opKYfQ5VUSCuiDwSX
V53kprMQ1/m5UCCpHUCUwMS5GhYOSHyzRMON+ASaQujdsRujm78hvyNDXDSQTv5D
hVsonevaY5gPVjbdGWvIH+uV0gVBsfm1rTuWC66hIkvrE7OSQWe5bp3Ee+CrDqDc
6z4LnUw5aZW+IbH3e04zFBuhjsAIXCkt9r9n1CNCa6TTxHuGDrooSuPcvSlfiw5Z
W3KymY/dyzzNdPf1sGyeTkhArXk5QIZBIz0uSeqyY7+6R+Pj2YPQxePQ7EKTwApn
N1aUiZOgOLnYF2DJU2/dglJpqT6rz0CeFDbFp9BIPbJjiPUdmctVOI1lJGqpPK11
peTbkoM1OkMs9R5wlXK92De0+bPrsp+SdhJGMUGokramNggrg4SWfvd7pZvgMmi4
Rp9/zkpm9k9qcF5TffGY7pFusLfj8/vr4jkAwsM15UvcqT2CdUU1xH7znrCyEBV8
YAljzhnvQfWFdp+NaG6fsTtLD3tBQUItGQi4G/syhtIeCcsvhcfndtWFrspMitsI
7Gjz180muKekn0sIe0LF+HcJykgR1wjLD6qQZgeHWXWO7rg1ke1NLQGRuNOoUi1j
ZTfbnyaJ0O67vV69ux8RVfB2EJLozfw6Jit4QvyK9G2MpigjR7z0IqPjVDT72/VF
Yr3sQM7zWmNL6Sj5N8Ib0kyTwUrH/I6vHSybAN1VYJUEyL+03flDYZ2SZbZ0D2f5
tgTc7chhqTx0/9CcLzHetbNqPTR8zAXFdpoN1g9y4iWV1OJKWAUUSwM5SXXVC9+U
QywEo24zwPkTlbXwJr9pDQ9yCj791lEhcuy4dyYP5xEODoKoODNjZ89XULLO+I39
Tb3hpYS0D9qojzSST7PQgBRc6OTLuwIevsLGLtVmLXvZWQzDMSb6gBVDYzcxnHro
UTZGAKB5hEgSku6KOJa4gX4qOAoz/OaLnaK6+hXcobmCB50vRmw8TfmY8BJEpl8f
d4eQfO/qAbESrB5gW6/vJSzT4pILl6ON9it6tn34hwY4/zo8mLXFPR8Jyv/Ekben
0NmJmT5lO6toOby21vWciC7md0AfH2UNJSfSlqHsPmJmgcZCBLIcTLuFo7ZJceEc
/caRkE3uaGNAdaOjRCw3azwNwn46YP1oQcL3cgajrYhrXi9RL1SMe2yGsiR+983z
j3yur7vaGZJNE7QyZG/otV+c55C3bWixheYjQsiCkFyiYlQ8ZZHKx2LDs2VrTjIi
oTn/4xclwNN+5qeDkMy2VG2bxpK9l6nzqsSeMF4LXS1RtWgZ6M4z6l3Z77GvDo4G
vqijjasu1ayO3NUw3kJ6QJzfjj2AbZzYTBD+q2Tgl0raBoKft62aXX9OE2IY33r5
uLhY3eagRiiTgXrjpv8MDC9B6lA3zMvp6inwpYT9KSCLYZRNVMFpS2aY6SN1cokP
7ZDIPrXcqqfjff0FF1v8w7u4ZARCuSwwPLch5q276mYYxuGv2N9Ka9U7F7wjE2uR
NgVVU+rjoXBvSvJ/V4FA27vF3EdaasGw94JCxbwHJHu+vO5c9D2LrHtbtdAilLnw
U0jF2wO2Ud5uDGsmTHbSpPQxyvM3mOKX2y7hV3d3sOy+MJPTOv2wwXkzbK95EAqX
RyTK356sGjamFzpnZykgvQ2Hmf+CjjlOKhumtTMXYABICw83v9cvewaq63x1wIPp
LCzKfQMv6azhTGb4k6DosbLchOHGcaV0W24PMF4UYTSI99qXGl8ZyVSXGIbIZMY1
En12EEw2sxfuouYLlz+3VS6kMGNaJpbCBqZGnYbCoAjXwEHyukoDSW1a+W3m9xG+
DCxxO4AN2VKSYO+FaCSZoCxro1qml3yonSLTfZ9gEud8M97tIN4TN0BE6RIadSt1
hNECdLzTIkAZc/erXWSjBHXVqHO67CmdWSRLZDJdu3XvT+h9riqi9/Rohn+rG8bW
M7a9JHQi0FXa0NyXhSU0Jb7Hcz/Kp04d00GQEbtB9vOYC/puA+7YBN4+9Lh1iG45
2YLyr2b3Gy897gJ9SZjENRkN+YCXUyywbPZ5ATqO/rRVJMS/f2YB8+GLhmgnnQGM
FLG968/h/8lZPYrW2/ZOwl0PXrVww+X1lJuW3c2ouGPduxpaEVOADMyn12nAs1h2
iWdJM3tPMWmBE+q4mxBtybDn3UXQFhlQm+toP+tyQ27sG9ETMSMrM83NZQv5MAQq
kfgFLolKL3UpIY8rV/hhmzMoFmSKqzmEJ/9HMsbQ43OfZT3QvVMdxo0Y4hxL/hyo
DtffQAbginrKoAeU/Evy3RIa7r7sQPXr33nC7J6WKXO6k2sd/eoIr4S7y09taP+l
vibWi0tTeEZ5jAF7IgsoT7zLWh9LDN/2WKdzVYQUNln7VBbDG7IvhhZVu6iN2yLT
e5f595vqdji+kZBTDAXnhiCG2Eqwgd9C+NsQ/5PiKKGBu/tmuLtOpZU47kHiDzT9
sIF7HMtdLnFq7UCaDD+LLrKhMnHpcaRIxKvflkG41HZcRE9C5U9d8/ooHkhS2sq1
s7QgkSZm6ZDA0MQHk1yEpafRqrxRLbi8XfcpDDByAaHDZSjet6gxv4UQc+HH6pI3
Sa9hMuAjEHFvQLVA5Fq320ZTX7/vWWQxa2K/LpJ47O0edIapzwvZXhI7F3/PoNwa
CNfsiBpgxfHeRVQbIawbTiJq/UwAProjV2R6gi0tTImf46cesHUYNPkmBfVc6K4i
R7IixO9VyzwG1A1NMfohP+lZVp3JIOJiw39JqfBWptQuHNMD7SdEZv52YwrfGiNi
yV0fWmum/kLn7mKlMvTfPnQjX6cZZ/eVLQ0jOCskwkheqS7Cnh3EM9m/OGRqZ285
lNej7V9JUpuBR9c0e6NqoeSCBnMgRA+2d5oWUemBlR2NBIBLtaJrTbBjLbPaZ3Rd
7A2Iv9Knf/ml8HcfVqfYgxMN8q6XzKyT4TZtJMVji0NWcNALODOjFGGxLrshUjMr
oD3o7bFLAIf4UjYsCwkUert6RVT0iMJP1RXBBm9DttkT7nKcCit6jW8HMimH56Dx
nJ9rOUZwLNLTtkOl6iW5gRcQx6dwkweZT6Xm0AIBtc3Jv9dkaUAfA9rv2ntTQnYm
/YOsCl/l/G4/CYUkCvwXzTKFNuMBFm9rKwWlRCV9RpPYXY6FwNxJE/fv4ia4S9x0
u1kwCEqY/YF1Iq5CG4MtGnBzStw2rNoiyfSfvz0xUXIopLNoduQaVlE03+n501qX
qnMJo4+TzDBlfPeps5KWdY0ffQfg5C6gm+4d8hJ9Hrw5umI4wp96s3lpV0dBXoeX
0LVLDQMirbiTnP0wnVlc+yMaRS6IFn9t58eTas5/UfiAn4ubrRN6Epaj+8DYqVQX
o9vF99egAmBMN254+FsToqXilXwn3uaAxRPK59/sqgU6pBcz5U+Qp+pH9PyFIwgS
jsqEs/0kyfDp58pBAuB9ct8aMDE0TzUPqOB5Mcjt+B4ZPrM1c3zC6LUuaof62YwX
kGOcarHmlykr5narnU/ehhMVm7tjpc65frX3f9ZQn3RNX1tDvfhqcNmBqNFMsfl2
xm/BKiVYO2OiydZ8EZh3PE4nxaPtyRQ+MUw9RnkY61jV9Kuq5xOTFl8YNBF6czuN
7OWZz9Qg1rwPSVB6YkEZQ76s7hRiX6DkP5wDMLgGAqGV5IMGfJkf05abAEFro29h
v9iBRoB+Inrbqb8lEKt5C6EKxjUmKXcNWWlPHwWr08WP92sgf9A8xnboyF7vhnZy
LK4NT6V0SYVnaKlxqYf9+u5pV5UxaGlKyBBzjDSeEa4SMauhlwKMSDHhdulfTPth
laRwR0bRyu1g/khkBrHHVn2uPj1y0Up18XzRBcd0ijFz1CyzYB3uqGLr+jpoNxeA
ZAw+xy3bY8qtnt4tJD2R8eD0RsqXCS5hN2ZBB2ygXRW8v199UCaGBuzr6sbZ+UbV
S/2V4GI9lgWwFYbpEnpNYLYGS791md67ggOKSL5J3IYFGU5pamv4S2YBm3DMboTZ
Dx3mvFGEzhwhzBLYWT1WoLY6b61udHtx1SkV18Tl7rMFH4Qj5x+31fs1U+251EOM
oBlSiOnPElZG32dCffKaUuyAmOGlBLnv4yHoaCRK/xJHw7mE+GIcu/RrHSt9/0yh
3hWG9E4qjqoT8MVaJEt9zdnCR416ZM1K+V/hml+1jqPS4ml8wTbkCpE3BtgIRZMI
uOS2DzqyxA7XR469FBie9U2GoJskyad0lSNMaUDNmAeHar7nteDloaljpifh3I86
EX9dau0Q9RuLVlXI0AE66K8fOb7JlPoJstz5iE49EfVdioSN6Xw2WE02qLJjgMdY
sQUrdliYZHDzKfJgpAWgIk9MEOM2MpofmFp8W8Smkccmz0mkiHeIyHJUO3h389A3
2kbhl3fQ+LIJKbFxXtNDivx4amJlkAqEHqIlX6KunlZ0AyQfKzSbKY6anhiWIPQR
EDfYf1uYaT0bg2ivYvZulylA57ugGXUEunFOJL47Bh/GIAGBj+VhlTF7RE7lh1hG
d5H4pg2qhjFnmQw9JdiTs+nVENoFwCkOWikx+hxCQ4lIJW9zl5fcbPRQiIEt9J+B
aVdcYJ58ZbpozgmLRXx3kqn1MsXmz8UG4PRM2+fCDE/ey3++Npyb4O3C1c71K0AO
xiUgYIpYprvSCVd2ioHDGKpX5moYPEqcdG9vUm9ssf1bg2lfSNcnu4svqfR8HcA/
Ddb1qegbELEuR1OnWxH3438NoKMBfbT2BDD60yhhjbJe8x8RvpQfxL3aOSJDVLiQ
oDcl/z5fUpH3sNgvT7vNETPGDDecbd80c4XCBXIvN/7LvItMvUSMPz1CYHyI2a1n
vt5laiTuHdmJTJVRhTWecMYFPqcX1lggo8210z4UJJuIfjJz12UH5MFEUu3V5Ydc
ZKiWZqjQP3ga2nEWv/ORhEBobB8T4p5q7Qjq+8w2c5WUBnzUZB36+ddOS5vFQrxc
7QAbpdDujfBAq7cGriWd77ejP3IjAtkX9cghS+YsLa4V2KXW4+E6sxsj+KLVvDrB
7BoxbEARmnoG4SKdL+rrtquffSh9RIXM+hsx+gbqjKI2Lmcc4A7+feZF/nMEcoA7
E0mgSIYBHSd8Di7XD9RpJ7rECmsaDeZCLKM1iZpNVIaOwtuNMRPEpOhVZxgjqLeb
45+hJiuaRSaVAaHr/AxeF5DXf8x4IPJTCnPMKwNj85UiV17ZJRlYu8LagDxw5v1j
8TJIIYqZRb1caw7kvevXnHEsS7fJjCP9Y0x7OgUP5uIMJ/a0hEESKHrhbG4FJBXE
SQfeQUKwd7E6i/7EgQWKxiy2miYaVXMEaWYB7IBzbeJ/EcP3/aCkIxwPg473ONZe
MTWnhx+ZYfFNoT2is3isL6EJ9tNlYOvfM10MjkZSG5ECk8gkEMYEvcziZokswv54
rder3L+ImcNhyXe9RCV9RBcmNcIpbGZzN0ZS7qVyUqbX3igdCwQXS9VbPYFDZAEQ
9JB7IktQQpPBTNbjjNOYbri4T9JLtblUzMm916sG6Db7+3T01Irky6lEigwC1npx
j4HaVbElHi/DebqJvmN7OZHsZvTQwNE+csS+QlyU1n4KWjOC65HjYlwE4xdexd3A
YGF2ZdXCmyvt4XR1wYQInTzbCaugB0DhkDC1hOohEYid2L/MaoHGYBH3UXwKuXEX
aKlWs/d+LrbiztR8FdCE1nlCEJ//pae4QYI2+jSAkb8vh+kpnDwWR5Hs1VX2eyJ9
UM0M42UrMec4gcc1hE5qJfXOT0OXaVsfqlak2VSwBVZ1l6FzAvOsqkhbECenNXBV
HdZGLQdKFRHsRJ2ftVv8VCrdY972otwnXg1GMSosmLRTwt/45yghQvUIIkGsFU+R
/hrFYavz19QKolGYWCOmUOto+8wjHbN9dOz/I5Pimv9VVOU//hmULKA1/BWZfmVc
wFipHx/wClIWT8gAkLy8MrEL5QA/50+fif1XkMlfHR78dfMTvpxnhY1orUKKHzOd
y+mwUsvX2xrmV+q6Nmow4SZXOybqFL7oPQpeBNSqd1nUpqVxVvXNHT5yRpcRb+zs
kBajI5OUqP3jjev1eq+0VL69dkl9T3/me9V/I/gLtD6GHuJbWqgBQiDNC+9LNxi4
gx0fPrTA6j+0SKo/Xdh+EVuX0xzhj5LPBDyu4JMZu4GQ49P7R1J4qE6nfKVjgiBP
QnUpGIap3Bdl3wnZ6vr9kJhQhhnFFiEcdqBmhGQ4BO6dFPqCEvEyGEXrvJMtlcwE
XqVjzdiNH6VlYIedivOGUUxTJvudzT7DcJkVZbwjrD9TudUuIPR5FYgeTlV9k2vf
daOtY2o7jbS3zAuT733uQIuLTli9hqTqE7uXXFJMK/szX/baqB4a19a1x/U0Po36
mqvNYIQl0guA//4QP11z8V01+4PPNq3EnRU7pqdWLIG5kV74bEtj2RrzvaW3QMLN
g15riqN7RU74RM2CgPpts0kSD4ZFUsioH2QmIGttXREbICmXmKUa8ynpzDrVR1BV
Z7jkx2QI04i/e1PMyXGnq50tYH5jcDr2eZ5/sr/k0cBa0MbibnqKbZDDfsms0nPP
gc8n3dNy0SUwAF1iClhEYhkwCuqBgx3QfdPUfhtDIeLpAppfatne8DSk/NY9tZoc
MKtqDR/1/fLwM4E0hAQ+dkhRsC5ipLscqwd3USF7tIbk1wgw+OF1eRqfwfftnmhR
/XMLTCrTk1+v1t8bkssHeh1DVAJ0Mf4wMyV1m5CTUIypQnl2WDcG1M/IkFLsqKUb
YxCr+8i0xqNgaiaYDiNOPYgn5LK/tskVePFUnX/CKHJMbvNwb0Hs3KyUb9v5070a
ZY1OrRV1msoQ1Sqs2/DbXFHXyno7MiQ7IEHHxRRzyLFEq8+aihu/Tna4aP5/9zBG
sh1D8c3F8ALKACC5ksYeC6QF+o7zOeXLnJ9yRytrvIpSlvwZTsYB63YmnvkY7Otq
EDCvbJ07f7JnoH5skWiiSmcNYED1qgILAsjr8sPD6BsfGQ+X0TPMpknp5rTJytUd
w+kgENFl+PZHUhw138lmLArOQOgk+bqn/+KYSP9jUdS6cGl9zt2MyfHvDaYBHKrR
JhgVjP6hOjLPJhCeuN8EdvO634y6GhsJWhMfJTojYq4lXNcdhAxVXCLfYZJ2TtlE
Tl7aU915inOgra0GuR9ftityKpIfX6PPTWGz3k8WfTujAzzU31FuOmoSs8RI+8b9
BdltJ+4aTDPB6mcdqTvU8PWzzy9wiovhVrrG2sXIaPF6wbXLkE2a/pQQxe01vAs4
TC0lFivqMd/FWje7BJ2aaMg+wTxoOiQKyG4UXqscx0B1tv6KLyJQjaS1Uv2fWGq6
CswcWUE+Tej08dWkbjvGxw0sKv4zXHt/I8imX/jLCoS+Eccp9F7nbVa5i9UHtksD
VFTd00D/VAtTPfVv7UpbreIhTVO/hVnLQwa72e1oIe9PPvMprXsm4LX7GMg06nPz
WxZXarCUjxXY4sBnkch3ROeC8Ueyf9GjLgFNYbpZw9Le5V3SRN86+uXCy0nHcOr3
kaVnVFGDMur5UmVxr/Xl0HT6pQgPon/cjcvEoDavbdrcSqWb2tu2xPz6iBiQWATn
kH8o5cO/t9jv0TRMKKBumShZxsO1VdUj4zzTO0aC5Ah4Q0U3hQWPs85DlKUpoM+P
aq8iEMD69tGGjlBsp5P5TPvZSGRO+rQYkfR9BD9dEqBznv9iO1NSjfef8OxqUFia
bwJ0s2iIEwSQ5LEkDbl8jOZ2Mk5CJwbpDUwtjUrL8HPx/iqf07RXCvFHSyAG2tSU
HTze6dtTjZxfeN3fM5Dul2XvPRAhj+VdB3EKep63L5Bl3zOQ2E3FDQyM6zeqBone
GbHr0pOeIYA7JbMsxHYQncn/ENYpnoTMl8qYKRcbHqovWrCLvmyztu4wh70kU2uT
5Hzx8Cd6EhYrajW1LBifJfeMTS2EODQoCN9eGv//Oovs3YaEI9H160r+6svvcnhh
4C337VGlUPAV6CbpBP00DUok8AYZjuYjTps4/gEmSnAJORbvCYaO7iUmzDQ6Xd+e
6sQHh1EQY1fNN3F1CEEHEM+GTjHIPh0SaXapj6ejwygMgRM0GZdJ9MIZWwZRjr38
xRT1YWZvicSrz6bNjDzaGkIqYNMr8/LqL+4ebcX7V7v/SIkvRzxeP1AtnavubYjj
6a95bP5F17vCXS9HjQGuvGw9fCy6DvjjldLBzDs3rbBPhoJxb3UOy+nQfjdokplB
PQSa012kUmBDG4WrcwH1pugIaDj4gnB8Ke8WhWY3sAHdW13/V2VQknDKRK4E4c2s
4SQzYg8BNYWtDMuhwZuJ2RkYljUhDe9Q2N+MnqmeIyDpJVRCptt014nzWF6a4xhG
895+evmp85UeKJW+KQcq/8djfjmxFmnWTNsUtMjHBSPRu4DO2yv0bTU5QnPQ2MI6
Om4iZjnEM2ACHaMu0g+Oc7oImRBzbWuyKGOrH9zQ2D2ty374Nt4q1+WCaRcvVL3a
0v65fJs3gav9HUa7+QWEcfquSvgmvzh+eNrlpCIo15q6xf+cCbe38lHb7DB/YMfE
lGnoBdsuKDpXDu8Jd0YQkRm+dh8ztkl1jvupJgCA4Y7Jl4D8toGNX8KPouN9HKjA
+Np5Lg8D5KGAqJt/A9StHerR51KER4M5NCz664oJ9PU6D//8mUBPz22s/Rj0rGJe
0ldDboisvmMBATUw+29EAAragNuQgf+Jh2bBMK4KsiaRTQj8WJ8j0FWVDSEra5RG
fSTE6BhZjiyijQjAj/Pu4qcFOOb/0r8UwdD5sevpy3zlCoQ9+4ZH22Gx1cefuHPD
a5oUt1Jt0sa3q8//vZieZljFuDK3giy4VI+UfjSboDvJk9YIFrVy2Hk49tBybS4A
1Gvoa85sNHSMpNLJ7vfnNtUTwtiDqWgwNaM+2ZQStmFbi2pL2QTtV5akrXZL3goN
UFuWS3UPbZHjxM0O6BA6tTHg8SGtvyrA7Z2KzSaCZCSGi326MLgSlFLcOvHmZ/Tr
bA6FwBiqD65eQedzzq3rRvQsHN7ZhKjCVP3IeCkngIL9r1G6IM0m2lMVY0zB7hsF
iQ4HgmTZBv50B4/SNXMoxDeyn2fztWMjZaLzfcOgronpWCqARAtTT5UdZ//nyYGV
g344JicZxgLRQFj279vc8ZvCWiSshcKnvxKm5MFo25fXI6F2DgqYLTStVA4pA0FA
EiZml+rUUO+S9mCwy51wv4V4hSwUN+R8INH3ARK4/xdc+vLC1wq0vVTdm8kvkZRo
FuRHSUNiGEU8t/yBh/k0RIAoY2xwbDcKL8mqYZoV+PbOPKcCpWg1JV8FDGNWTQO8
aYU6mBOS/Syz938meu2qDSQ0CvFnzW1afsjtAL43+JNKSqG9ZjD8pnLhl/hXlA1Q
BCiLYOazsjZKlApJcq4vOXxbCAuHavRozliXpBrdsZenpqWpbAmVAxv+Cgtfj1xW
xSIhWwTU9CGtgnuiukxciwM4R5E/uJPpvGp7oearAPxYrKlaKjajCXtl1Y7Em0wJ
43QeHDMGBh9ztZcRiz8BmTkp/MPPBeC6aLC4gL0fi51p4l8nXROJWfu8fD+CHLB6
735bSIgmwoioQRJpOyehETmgEujC3Y+8+EDcx88H2G6MFgToQFFfWSX+kLVwNQu+
9Iw2HpFLgPbb4kyv0jjvbEEJQnDMU/YzeqpvKJoXMqu+CGaXIOG0VOkwAq6FYKws
w76xDvJRRgEsjUk4VnX33BMXeKGVKdd0kv3rtsz68pUBascvl8vaNx/yjid1h3Ol
h9V+AxugHDCHAUxFbNOjE9rxncJ21fMwayueyf0Fd8EvbR4aEtSxZll5FqLdP2L8
QHvJ9ZcmnLrqtV5QUMhtDounv5a36QTy4f8ZyzkppTNHN2faHcOlNWWA7VdlY3+0
wONQ0X5olSKUxYrq7CRHujgn1Pa1BHC8IbBzpLsQcQ6h4ae0esdixOLyeYbQQRG3
w3SHZQo53lsbUzUaqk9hdq2KDi6a7cB3+EwBLjkKeOOaOFRmeg2Umsuw2NLbeDM8
AsozrN4wAbHcEIpZqL2i8w1Da4qOqlSZPRqtuhJGXYVL/GuPLnK1LtIZ0tUBJnq+
G2fvggflpbEpSgY1cD2e2/t0X+0OrHhNchgreYKVdy04I2+xAsFaIF4VIXs46Ox0
tavB1kRL8cojyy6ACNiecWumNAxwlDm2Wd3XGktifQ+NgwnX++dyLwuNEygB3QYN
XiaRN6kCVVXv6SBCf9i0bp2dXNMQdiqhcjIRs2O3c74AHck4nk4hyBDud3+uHD7p
ac+JirRCk6y4BB2uFK/z5YagGm0pkKwukfpKzd+lvrBWlRD4ivqo28O0Q7pK346z
WfXZ8IJaVBYH8KIAdQSWF8TyTJbMSuyGmTaLY8/gpT4ttoO85W7m3vhhHzClt+FU
PRcFchS8hRgwqLaWiPvYNtseUoiXXy7t9u7vdlbvn6HqkgAbgS2khYq3NBVyjbXR
Pxm2vTwkH2rJDnrDrTVUHOxFJp9NbTGji9TCm9JE8q06reR7JNVWiKXGre8ER7F1
J6wez/PTEffcRZxIwsPGq4ebz+F5IegCDEo+tN67Qwb+sBLpHAa5b/nAKtmCCkBj
2iVlKKJ+f22Ia8J+dxuKIX5Rzb1arE3dSnNaatBmBiBgO2pZsicDE6D+Z4j9kPiS
olMQrc/fxwkoDPmcNFbd8wivFhBGdSDEXYdiOqLyhDDf608Fvls7vsbKcRrj3G2T
/b+RN9LueODQex0dS0+7p26Z7eH2/wF4ssgLCHOWdha9lDgIaqphH/BLNp770pm7
RcFlMoGBy/PoVvaGrFgZ3dzWdglXKY+6g2JQnQ3l8GvGtJEIsNkD2JjHFgaBtFMQ
HwXpvwdd+JCdjc7jGkjqt6PtfYHODOMEFwefaNUFcCyMjkZpdl4mQXkN39Ix7KsZ
Da33NfNS4qJ8yNtE6thUisg6VGMdjhUMIhivg+iPOH7y7vnlffTmaB8+3CCV6HeK
LsQFeU0oVceomVaOdNIiGvclFRiv2kjkvfGmQTD1+eG2dI5tdealW0J+f+/6+9Zj
iv/zrRhdb4UW5dDsmp3YuAdWiVkrUT/Jq+HSnXQUoFZDDWBHixuJJFGE2lZC75LN
6gHcOg43ko6zInYWbwW2u94TvrKl8amSEVZTJuBz6a4x9A/s9edd/NcHZ5Bvt0jB
4B1kOyCvl9UrlZBGEXz48A7ZlnyXw/gT8i5BrKmQObRzngMinzPT7StXuFzwUnoy
llZB9fl/VnnrYXS+1WSeHR+5H8w15KUMwDbjV3G+W2ZSdBNznCm74/wEy+rJIABO
xoAcd9nzXp+TmhKNO4ZgAmGuL3Duix1lJkLXui3fKAqXKhJ47lwuo/Jfrj/JCQgT
811USxMFT0iTz4tSMxs7X1IueaON6QTfmi28PX1HdaOai3bzQzcjkYeKmctas3R3
8XixZBoLZPgC6IeRSNYWbLbedokHavpK9iQxLNCdx+nZYro8n5/RkRisibjV4L89
yzSLQ51dSmqPKHZxtN/HfDv0An4T659KeTFidzyPXX4x7JCaTVx2H2PAR4xCzCdx
DBEug4728CJK9BbPIwgFBdotYe26C2bV04ajq/iw8GU51Ujx7KksMyQqpnHhrlKO
kclB3Cnz6vlDk+M6aL43ljEJjLsXikAD+NE33JtZy0RCGjr4GXQVSOhfcVeLes46
+aYraif+EzT/tXC7AXf+q5GgntexiUBJQD3w15/pWp9CLf6DxWEiOt6mGukTfdzs
iF+jyHe5DSk1YFJfon8BrKDvIxgHVwrZpFIVtz+Gm/yxdKE2ncs0WdpN6GgUufC+
T63LxutVqzqGC9y9sT1iYsRMu3O68C86cZMcGVAfmx53rPX3rWm8rVLkOVg4sJ7g
pqDc+WpH3sSil+xJrTwlfm+QbhZvIWNrhuWdj+4+NBScUsYgiBJ3z3LIFIYNWVEp
OvvWjjVYJxNtD1xBVhvbJ3UDhslroOoZ6j7jTbnXkuEMWQQ0Y4aUGrCoXaTc7sd9
koWGSzCdLKd2N9wr1nlJxKsss9l0mxxUs19LgtDFoVCz89PvMgfGCl47RwT4bmUw
tRU1vuX8rIo7Hr5YUGtjnDrNMGCdfPaY7lV/CLLS5bRZFd11TNmUJefBiO+wH5jY
yN6xGdXCPDcMGn4PpK9CjeQcwUQYzAtpKcHgvGCxURobS7kb5dpUXMyOqWGwpgaO
837g28JoF+y6Zhb/Int7/I4toFl6LlbIz/+ud5ePQ9kPQ96gHw/bgGUg0GrS81Ie
rso4VM6YI9Q5H/tsuJKpZdawMXyst2oY6sDwfxdhbuh9NTgL6ttcRpuwHwXRSbsh
ZncKQGDAgZ9qjt+YMqaAe0qfTl3M+vQoA3sD8ianY+OJUnFMxAcHMahaAgUy326A
/VYixUkq2JVvsMg+5RMGAnx8JOJiNJic2Fx38JVX7K8oxXcajmi8Br7OHVXRtfr+
Mr9/lrQ4srhhpe7p4LwdYiHX+mbQ6jWPYvAby3QkN1ZUzQsI0xCCgbZlRs3mgRgf
fjMb+ZP13985Ub+zc5hA8+TB/aSIUr0p8eE6jdutdrAy7Myx1brMm8bVMMEeI7d1
B2MHV/nUysgx64+QnV4cxp9+WyT5hF+ro4JypRyW673RTm9ScT1JNJQlRhKjhoJh
+zo36r2zxkG1+YJxoro3KjOGSmwhXq16Y/PGJzWlnaT5hb01GmSiK1l1bgCR8XCP
erHyVd4xYD3Cwd92AbwFdrTmuN+RqRKBNCsJjibqgRTO8XvfjWvwzfrAWcWMaHGz
LsvFGMGcNG0OUeB2pH3srBjWfLsFQwQRmgAYAldYceLVrT3RyBonLrDx2ZRtYVmP
vjti0rxQUwtFDhFfrL3+Jv60P+YhtdbPSnsAMLjt5WEUm9upEb7scdihjjlek9Ph
wmWdly6HgYVd5grPPKTMlaJ7MqwydODFZvpMnWVpaFBvSe05j2eDB/HAOZ11SLdV
64w5GiO8RYn0DW5vbd4f6KxXZxZci5dBcM9wSBANjPYZF3Qm5pVcv7kgCG3mt1la
E8LE+iS7kP6q4M0nTom9AutRPgMjLDhSZXQfuvbsPCsBZ4zfGgty4J5yMH7tPJI/
HV/yKWYUYexQB1lsySFkHET3xVocWE2IsNvoK/Y+fyKENdR9xxkQiQlXRdSNHp9q
AG0pqXEwamqYuwjQ3UiSYpn5hlYGnLuK1T/f6HZl0u640OQxnz6SP5p567VlvF5g
Yx5BEnfAdXFOwZGp6AIcslfpPAfqdSzOWepf/sta08akmLp69TSM70EQOrpYW744
P8a4PXilLO59N+VCwT2UkkdJcuviRrEq45dLieRSaJ2Xge+V9GaXc91quRiKB8sb
uYYpzZBkwuGLreGK/W4k31oCgokTYRqael9WMScIyqjfUelGscXh3TxqxbHvj+yo
KvxMBdrrFUzpO6qkZc8Jv759Cj2KoP9FO1+rYoM3ifjwc95ESkQC3J41IFAr7WZP
fID4abLjkEW1m6UNcmxWV66SDHy25znbElyXLpFizs8AJA/8NusB2R5iEiFJ/dA2
ba3iIylnnhLo1hc7ukNyXg+UwKLIAeoO+nj+W++R5LKXgkv28/aSa3LOLqUGMyTe
9aehM/LQBRtu3UAKTW71oMs4rRNmt/3nzdGeu7NL3oQzUNaKM+hUIjlQQnNoq/QK
VuPl76Lns40qNTUgEpp4Dk63niIJyBdCimzPpmom2vUmEcEk4TSiGN4KpFxYos8L
Hz0ZaPwUt/mFm0g4e2NPzr5aQrO1+LyoeKYO8reefnTJHiSDUWqNRhi0NY9pBePb
bQD9CRSNRuGSxQ1aln0ODd7eXruGIfKGPX4guK2ZkOsBdr/4ad++ay9PJ0kxf+hL
HjlAJqmaGfYULCIXdvNnMn0gZOepWVoAMDRKFzdhGkMc7vdmDpbIg+mTx2cWSQaL
MAZiJHCWyXF6PXuPPeW9+pTeerZet2VYuwoHDRkyIzIfqJsStxCrVaPwoCuS35QS
n5rupVoY14SnxTI0LPODCbkH/E8euFSBkQW6AwBvNPVx7hHCkB5giUiTLYlhUg1X
9Y9E8DlhabOWoQ7LgcLo4XGu50xkQlka7ZeX1q/1tnodI0Rf0e2FT39wmfgAZ/Q4
wOQVvUkv7HoNBpa+QP9vMTxBvkQrzXJjI6NNUS2tuGmyRxg5f5lt/aCfvRpp8vr1
LrdLra0hK+l06LFLEFIkCz/6AeBPcdbt8SYe/a3fOBfIvQZqhl+PVPx0poOFN+f+
MHu4WMNaZdBWzRFo0+OrSaGGwOxlc+qiEZclM85VuBTO5I0rdg7rnxY6Qww45C51
xG/DAepT0lMZ0/V+TmHfebV8Kllmw7AZChI/6ZOSpqyWgQAXUiM/a5109HEBwInw
Dvnd3mhANaGQR1KZXrcuZWHWqMHyRJQgb3+k6wYJ9rGjdZPa9AQeOg3m4ISVEOrA
mhp9k5854uEPsfdR2TNFMaXgq71ll1Fg7diNYVDk75KWc/23mhLQ9Iv5muqjGmxV
GdjUKkNTsIyY9nxgAfa3gjsn/HSRw18mMnAV4SMegaaaQDqMgPMQHLpIBEshr2yV
8UeU9JPr9Y7me+xwxBrjmgpGj48+aNjGCLA1yun2VBUTNcRbrEH7pP+QFPApq4ht
5K2P9VL4gefhc7QMpQQw5yAS6r5oMFE/XtvHfvCsRAuHQ8ABy28+TJ9tI9/gn3j7
ZdtEEXOAEO1TbuPl/RHf4hL1dV6943B71SJbXzn91Mhutrbh3kM0e/klQSTQkUPj
VOQdz/o/8gX2v1bqJtubzYjVFrJqCEnhibhjAEFzzIlp5IGd3lJGMTANBEHU/8JF
6CWiP6RQbGGUvgsqlD80HYYFA7E7nAr6JqeZABJVQXruFoPu4sDJNfz24V5eDNBJ
vJfwEl2J3EK6htCuzR8rIubiYx9ZU+KY3q2Eqyg6cDnPqArYWqenACGPfERbWUhA
SXw8WIRi+0dC7Cg+XJAsObgRMXib2O+K2J8HYCSe6niA1Ydj/7eIg/pnckNv1xXq
B76xw5lYcn6aQT5Hv4wXpI1w7uz1G2lf22Urm2ZW67LDEu93j/CFChlDjgnAtjWH
m0Lio+VO1xtCBV0a6wPIeYWSIBb0pqJj04VGLyXNDDCnnub6JN6xWTEvvChA6qQr
fUgdvYDnhqVJPdnSwvrIKfbGYldMIl2EbYF3VwIciVD1jJN6S80GKGyVEOsh6VEx
RlphuUZ9f/MbHyRmGZ9bxPVB/fTHRhDyYlji1iXgb6qKAFHsChMQEBDIw3v/luma
6Ap7FOz6vbPYw9WoOVWnJVIInMI59Nl214sHj9Nbwioskrf4A5pe8qWHUA/E5ofA
aV34OV0V8tv3zlzNSnDptiJVo8jo9bkKi4ZevFFZGIDl7QCzL6BuCSHXH+JtdoFJ
4Iy1oKphp39GFZvP/ufxIeAJYTyztJCZR3ROQ1UOVSFouJ0WFqYYiysicmIsbDjR
X07+tVWI2tP9Az4HnadaQn2C+I5QKdDCKH11upR+z9j6QFGOEYChziQH7VYx1qIj
G03yGyNkDtWSsjc5Yyx4l/0s7oscqKrOCEN//+g4gEb5vtd2x1NrmF7iIDEp0LVZ
Ng7qpKPYf/lLkjCqkFX9+PdVQGpLutD4QxRZdk+Utcs97dmmX7flSLaYi8Uutu6Q
70kKlbb21IQgNGWKvgDBGI+ApBdksCkmLgGxVXtvcrbhy7DOwJAlTp9qjaFPvWZF
IKZZGzrw//3M+AQxPvwSLir7uQfRZBsFeYi38OZtnq0UzSr4PCyPy49RzTJiMvhV
ZANXvCR5r1fP2fbrhI/ROUEvR8d/Nt3ETqYFSTpr1PgmKFKhJOQ5vlXMR5ojHiob
9HOuuoXNkzY84p0thYYTXHzFVQzrzIWQ0lSEEQu9Q6kZFtPheyjJqW2h/l/6koja
hTHztTPecplFrBVmDM1UMcZ40h7OQ9L7rhykir8WCKSddqxCpKG7ZJdHOYQOvDmg
bBbcv5KXZO14n08y09QYljP1c5AdmgukS31oMoYCEOpqpnW++a4OXps8u8L+C+Ib
OW03cnbYf5uVBJ2g99xAUzCnhG/NFeSsKc146g6AvPsKpAmeGx/jRGObxSCFX3Ki
2eCoI/UU7aId1AAUsqu5b1b71w+hT7c7yudvTLgtwQ+daMw/m4RcGYkO75pF0C1m
4JDXxLqaTfpXCbD4Bpb+Lw881si5E8f5Fp8JL5s1OjPlLBwSqrVECXK9/4rDlVK6
Yv0bgqtaaIq+lMBgOrPhcfmWu8KN4ahm2RjolWsE0pj6DXSIB/eblMpzGNlVYxIf
ZkPdOI8VvBkv0H7Z8HQjsbeK7SZe0coQPeJLrWaL30w306ZizLtRGhk/ZMRguK/C
4AVhsd+V0/NqwYCtuzbHP+KFjrl4zMpY92hwe7N3y1hJUYTqU9tjtnInumV2RCZe
XnDdaa8hgJMGqJB8WH13HXIIkrI8EInWgUJsR/N13kocISKfF2ceNeCgK0E8Zonw
XrmcTR3QqxhC10SGEppIQImqn+JwER0A6JmtfrswZbY4zYO/gZMiUmdI41JZyIhd
2/DLioS055A2hwBxECUl8Ab1qjgrQcqpijmncnRztFgRjmybmnGSozs74o8mAvMO
AfjDNhxE2ytyTKpd/Coxp7kBivupc+hN+yPnK9bH4Vnqdt5xYTqWRvLWpSxvOpWb
oifvEgb8TH5LClgBKSfNdPot7w0nuNGjtE8AXFff2mSL59N55h86zRzdFFETKoCa
WUNzcSGChT+9/I8MCQZXvGOWSvijtUtizo6Y82T2PL0MD5xJIROloV+1TkE0N3Ux
bqVIoEvOPjRxCX0w73LJJucwwyQ3i22nKMWdKEzo9lNQa82n0rOwSlnBJqoru2eM
G88okuw0wLAXN89rvxm3ZEPBRCxa84YmEWQfz+ztyP1j2Bxlv+k7VrFgjWT8jP6l
TN4qZcZ2S5Au0K4ULxKF7W4d4MSmrdmrDXFDOOxANzF58oW/Jjydbd3pHE4C9ysg
joOBa7+1a48IaDQPupRle1nONVN3VL3qdZ0DVqVvKwpJO8TCM5wxlFsS+s2mbtYS
oBvDYGKnpll/xIKzSlXZFxCP50GtYnk/lM8MKtfq2hIeQ2AL3/J+b42yMFkTd11a
ryzCqOhb9gMNoMuZrIpEZb9peLfjIOdG/8NqdhgGTSJWu8pe567OYe0mvYZnjLmO
Qdmy06ebD5LYERnuTP2FuvfHFW4CYwJyy/4ShZ8TOqp6ILErTIybvMLIUrjEGQ2l
Pa3cBI+qbDFqlkCxUk6gJF0n7SPLrcyvP4+8bsEh/Syiki6d/WESdrsdltclPtwC
aF8cwdKC3MnflHi502ULnlOsCRximPOOknuTpBJxwy2JHHGeO7nWNcSMFbM0QdTm
13PWOj85+b6IacilUtP4p7dgCFCl/fy1NKGo4ekbpogaSXLowgRkt8OdNFoNc8Px
elSLyMdW3e1WWodWEcAfoYq8D4MO9G9eRD8Jt+zTe8+SYvn0+zu2w1wU1fRdLOWn
c2oue+sRBZ2tLLFfH990PcFzHSvTmVJQ4UDhiGqKBZFfabIZOwXwCkBeXBOqeqdo
PloDjwjdqICBxa8WJI9r1siVp0MdWS+KtS1LO+s9ULp2gZRsfkBaR1UnnawNx/NE
BWT0o2KRdyYbqKtBRVdrNCtzjD+PKbcVjRsn69uEEwQRzK2No4rmzx24FAVGeGOP
gEkPi2A3hfHpCfhgGavfInFVMOJrUBppJ2AtDIRzBraKCGvqJVlfO300qxQebeTl
qN+GT90FE0axDypcU3RNj+6ggXNAff8txM0LnPZKlmOvKC5y3F+TtbXbATvnUcY0
DKd/RrN39WjlXRL/hCD3aCDJmNM7Lizh6eTsNzoYv7AnwTF5DJKtEhxY6xn1fape
GbS4lFnzr4uylwajfTMKGmfq7JNPzoSJDJ9lleaA8+4Iy0J69gkXJ8Blk9s4Ft8c
qfK2PjT1Br0ElC7I1AqURQLDrbmOWiUQOdQ6STLEG86dTnjHnio52YfjXo4PZ/NX
YabI8KAeEvnOVQ6o8NVOnPz29HWNiLKpZGyXjSYcZdL5IBtazouhmnB0q9MGhrOe
2igHMP2n0tasxvWAiSdQt6tnltFOyzG2z41KCrGcYfiKSF1JmIBm20gmojQJ2kUS
qjaUs3zc5HBI7oCbckEdZszL4PwmWI92CVE94b6rikDkqlHHt1YhWNQ7bRCRyA7U
Pk4vklNXM+adMErQbETXWZWUr6onXwV0pgDKaZXvqZMYCHzRfS1UD0fWCQhhXpgU
rFulWhLy4Z+Kks4G07syfwHw6Z/iSKQq5gymCRGYyfjcJZIQAfK3R/YbRPkB+nd7
qAr8UZLx/fjpNU5wTYwf+0jqIRlHZl2x4Nu4rxI/XyYlLlIwLvAo1SOXsobIZlx1
yNMhdedRQNe+giRvjmfgpAGp/Xo0ALwXwHXI7LK9hBd3oRpc99DQ4GHZNleyhI5q
w5ObxLJ/jEGJV70Bgb/e94Urv/knrZvElzFqoy/BHStJ97RYNqUH/Z+urrbYEdUb
QA0d2G9DTxDp5wmU/5Cw0s+FstOF3dOirqYkQho4VIzwep3gC8OKRb+4+GNBAjRB
GlSv75nsGxTIVUtwr40hD/NWsby2kAkFvprLH+H0sOCpmhi7T7FKY5BomBYT1Q+/
4s47Sam0QRh5IVqdGAQyxkkP4Y/HB5m8IHwQAPZ6S6teslJYib5gZ8U+bMnPS5AZ
kCmAUyoiBjLoDq3eYvVrRfXgcVm1XKTdsscXpntomyFNa1ZNFmspy96QC+j6mLWq
XQPh5JyC9AS2c5+zq6gBQjqML8XJgXAQI1KdHGJiXHRXKfbnD11D8B8AD2il1Ubf
giAV+KykVSNPmF1sWztInzfg3nKVtz0wccGiLduGFDQrRQWrx5Ld8B3hC+DLxn0B
m9bB4oySs+Ra4nhdEydhoN3uvOCMZ1BvMP/pxsIv6fu/EnYdHxHTAzmeF/qV7OHF
BkfRHsQ/V/zEmrhynjERWDAQiGkt68SS6cymXHTAimgQadZyUNJGTar5FmaJT1w7
pj9gHz5S55Z/IAj+OjW8hNbFqTTa/dWgupSs7M+ZU8Xhv32hAqDXtOpa7I7QsKbb
b6GDFLjGnIqTpBLGmTmrkDczJoD+2v2feoryeXpjF/90yAD52Oc3WqevuQFF5gTO
2Ol4TEtM/SYUqOnRGJE3YQYIYb6TNOGlO6FwhWO/piVlGr4OAdjAzYvifIrJ9CVA
c0+F21+P0iYMaPDjEMP6SXQc7l4d+PQdT+jSAMKegPjQ9O2G8bEeEhcAvpA6hKD/
xGMITZJI5jr57DK2YzWyaDhNVdgxZnegJLf+WkDJGITN7FIAH2S2X/u7SdV1Dj7T
b2xr44AwaGMMLT91cqWdx/IwFZ4QFLwF77BQAZqRuRWex+NesC/5graZd3JcuVS2
fOzzeeibYYc93fv3vWemLm2Ba64Uxz/NKlG4HGBqfJdb8/kTSg6biN3Mm0N/UP6p
SETslFMnialnt/3uU1zRYYuiqMnB9WO5oBCJ6Kk0Wwx8uFqUzoqrzKulQY2MT/+O
tFZ9TKzLng1jWmwjVnbULVBjbQw8oYN0yatw9q5DYA3I3eEFr55qwcGKoatfcwZU
bzlrYDaEGgwOke6Iu7pG5WymD/lxYkqPLqw7tIA5qgGUys89ycUI4nx/892bH99v
Rx96iPqycHL3YOJoRHVdSaiKODLeVbMT8Pp358l6rY1jl0clEZvaucWQF1gEgfrw
IANQC2RTpEIJQ8ysbU+v/P5csmI2QeL9AM+jtTUkbAUjeAuJmIQryq8huw+NFXGC
yij7GPYGxPUNU8YBwVmdjJHljWilJFNLxQV8426Y8j02gNxe0mwQ14aqkB5y7jUK
6JPlUmEkgijHOEx8SwqZNT/weSSEGskrACx9z+0JyHNTbt1SjbLTZm42PAcclAJv
2L3ozigARTjAK4hLJQS6hP61ofszQYB54Ys9p8/guB/suc5QzdsF+QWZ0jUtlN8t
o1qSeaja/TFINLObckWfRP8jZZ8DVWGs71y4HdFZWwEYdElMmbVV/hOBW7prqz6C
b5GcYZ81tOpWbFwEu8pHfr9776PhqEgGDXesQHyurCX9JsNB5taRPtEd6nrLO5pR
MhtH+QgKXC0IS5zHUOYWz5m1q/Ls6kPJpG/HrR5piTTaqmOAMhm4Qp0FhwIWjSPE
NTTGl7Ac7A0NkOpP1EaCu1ew3uzDr1BIkp2lz/esZ85SUCOsf3YopX49hnGtVTUC
wqFbUH5Q0PEqN04T4cf6QMErgfEwxXe+OUdMYz2Y1epVKrRe/P8HaURr372gUePs
RFmlk04haPkHAJchrvKvPInOOHYItogWS8vOo0dI5he0Npj7Ueh4woB64/40pNJE
YQHaSVsqnEqCBK1mpts92SbRgm2QEtKufNFiEa3fi8rstTdPLM+b2J98+mp76ozP
DlPvcH0+hRzLC0QhE65j33u35KpaVIW/+FzgKMAnWHKirRJ2I0lGvRxuRa9B+c/O
dwGYhYqMsLjIJkW4GVmeaRYwlKfm1MEi1ByxvvrfG/4mT+klBwMI53yzS9GnkQqw
K+WQH5GWN7z1MDaG8Bm53g8xgubtuBV3jGqpuvPSzyaXG5fvp0D0NkUFpDWlcYa3
2VWxz/N/ctlKzA12xJa1WtRASlPUTkHd2ZLIqQaLNQGgrEr7J0zaQfJWCsSBOeDM
+0xu0np6vQt40XFrCb3ywbfuInzdOrR4eNGb4pgBV1igzUlYcXxWl8gsJKOChEH+
IMFVK3zv3vcn+jZ0DzJmClqqCpErHXzJ4FOw7RDOnYrFxuDME1wEfirEC8el+j6q
5wYcUQEaNMkDuhSosjauJ/Jy87TlOaruH9dnakVSMx2LQXKvqRLsBkvDuCzVsVIf
LyxayCHO/YgGiVmS/H/RT42G/+JYa/ytFlItIGR76DyXCEQU3Niw2RaDAgWeG8pm
cW2tY68/vWIfcR4L9fUSx63kS+yPXZ0qMdtT3uAIlrpRJqssDeTwFSbTZ2dwBDYn
6OSzsa6jLC4XX+sF7ksFC4sfVexbbAhe+g+eerZNWpRpyGob2+JOh7Oz49rFlyBQ
3+XxtkE7XhJNCClT/CQUndEyCtZ/G9sPP82C+9zqwaHooLNm5YOAK4j9ATgfEHqZ
yQ3n2phEz0CyKYOM3EIl4LWeZ/Rds1Jq8PcDx9u1nnmHekgMqfC9niINBPHAjgOA
541V8Ae+kZb2lbZCf/S4J2GWJe1+T7yX0BXjvQbYkFped3+qQgoEl7lsZg7NqEG1
FdU7aWLbFoQxVFq27a3e5FbkH5sWIolOnGbvmzGCE0vvKeHjzHDd/6hz364SWKbB
fr/mseXyz41H5FJIKVBTNyxDoH8wtWpez0S6Aox1lpINI+5dsWL/FR+RkY0f1TwE
KabFk9fTldnxKAI5zUS3TMuR3dsqKXp9V7t3UqwBRGNbQFgW8BpWx4Phd42+eCV+
sYdFRyZslL0oEEFMlzhSevBen1gZkNj5f/nzY+L9PO1Vgkcekv/IZLyQXDHcY/w8
CsSNYRJB3GqjaWlNybDONn6EIADYWEKX1ZyKxU8gf1Jl8J+TG3al3eZ6zdYToCjT
S0t8GEntGbZes0NNKwUSeesi2gm/5oAg2Zzrl/lJ9X5JbVGg3dSgfzUFny6IbHC9
4KeZIVQMiQa3eNB98j1GLO8HKXlLUzD3dejsiecB4Pob3En7qkJHphf81VtJ3ji4
ev6e6CkCESeNvUngp+J4Bf4yF2vYsUoVnlFpcWE08OyxnYucQZE4IIMct2vLjmkb
oVYpAnV4WMKt8+LuVyxTgvPlt/86UNA5JOHn1SRcfn7wLAq+/PqUgtShCA+yhB9S
3eaUSRXYfYt55qtFRBI3OGxr28i6fEEHvvcwcSHyoNyUL9/5TigG235JRmsOkfSh
4KIcIKzVRpJ/8C4dR/ArIEQSxhzBfP4dKcxZCdBM87uFthoGG5eiaGUmcS2Ou2DQ
9Pwt4TVwjO7zcF4U+kpGDvEVOzMeyaZ7utqGX6amLadmcuXcnBV/AbUcF8XIaBZa
0z/ox82Br/Ru1fKDQp5Gmg1eJ7lfH1nlyY7G7xj+mOxWH19PZSMEWA23fhKWMbhh
qm/XCBGtL7DVtR80VUjdCkkOUhMV0hZd1m1cwfeJmeI5DtTML4zNtTbYJuIiYHWD
YzfVIayU5ZhALClhzErlGNDmaBhKE/Bwcvdi+465rMD6e3vxkr98uqJwPLM+haa2
0CuOwmaLzppW91RyvjHLz9mS5HK/XXdGr8clu9fVaIy1PCozLaQ04ORoygC1iNiP
neZCPI1cL+BAHEFaHyliiFknfj1MIqgW6XuCaFtmi5iAU5XnPM/9kvWQo5Rdaume
fiTA7VdKaJDwXUFyn2mBLwRwjH/rjfklQNbuP3AJZHNUrNzSWtjmqhyrHHDjP9kG
5yg3pL6SyBPVKa+LPwSAAQhHbAyeL42j3CP/PG9R31raoA8BFxkje2TRVRgqXXme
MvkrOectQwEaJE18lUN8LDLeMJ5uVmojXiPFFt2FOPcQ6V3pl9rVuHnXX7wb/Xe0
CzEDYWaTY79/VXTOb4nu50Tko0PRSN6BgGDr/veFCgrC5o/nPqZGfLWlWDw6b/8d
Y5ezq+g5iDDNhRT8SL3uJTo1PGKx/bXkUYQ2s4KpA5A87xh8S607szVHqFzV333Y
NQZ/sPDQhopybccxddlnBadcY0yy6MUqU4eMpIoWacOGBdy0SzQlT963XA4EwNlX
Ub5JnuBlBxxry0Vi0ATVBe7rXkTAvHF+QzolAa5QrPOc/6FIppKMkpRtEmADango
7CxbpQC0UaEOBXbxp3brxfOht3LR2EADtSBAW1Lfp8wAS0fd9RciyPBc4OmjS8xE
3fJ9JEadnQPN23pJ2JdXueQFn65SyvN4oMcjorVah7cD673XYCEOhgfn82/MlSQo
/dRi5+qbJgElv4h4dp2Pg7SkXtssVZfZvLlumaZz94FM7N/rsiVBXfYyD0IWI4GF
1ISSDFP+URk+vLnHHRt0SBBSu/Urw+Vu9+S8HBc7cSYCfqEgk1PV9YTKJAexOW2a
hLjdZ0Dm+WIKHVPJI7CUfC6XF2tK1knO6TJ4QJRAtx71sSMQDelL6cBsm4SEvWM3
Q71We6JyJZR+6voNObySMYqgKZ5VT/TB3nIb6s38Toxc8fHeWa2HcXOQ0/Y77LtO
4ukMSslKUaDzghWn7825JfJ5yjSvmkrhwnzM08ilFvvcJjeIWEXi5bDKAd98c4Ca
gc1swDBwWQSyeti0E4Y5Uh+9r8bzZV9CU2qx99HhNG1LNM+i8ASS+7J7flh23JTy
ygmYpFOjJa0Mqa3WPzikRJ01kAT1w+kGsH5dSnaHI2dUdQO3Copt8RA95/Ah34Om
L40/Ji3DpB74bmNZiMUjmkTUvoSQ21s/iW8ql384l+xSzZceRpYcNrJKE1qewnSS
oKAsenmRGCJ2b/J4ARq9PaKhnJ0L5MtIA011ThorjN8A2U3H4+P10dE+i4KCEX0k
eqcmP298un9BthrE6xQj2/zYxEdP0vh5Lu4UijyanvbFvCo7xCTFGMtXzBSqsr6N
/OlNHI56JVtfzveVbBv9WEJfpLAbivaNklLfFFX9/ys603JIrWHuUTEaeWrkCfG8
jfaqcC7AN1Mj8Y10P5cmz9PHtNOdHiaIHtViwBy4gJac8h/fwwQxyWSB1D839LfN
Vix+s4Pv6VF25DOWd1CEL4/mFj2EPHmggy5i3iD1ZnSriFYqafmtel03D+TD65rl
45FBhn0zdar1DiQ5GIq7JBP4vuYOHtGf9wvyeIWf4g8s0neruLQSH12wFA8GJlCv
J8UwKo0d3YvDx2W802r41HHhBW07pBmyoX5ErWx1FcWKIsKzPTVxd2jOdHiSGBg9
AK09PwGxGMJXJV3H4xM6D1EvVYr4mMYvCJY5M804+e63g6BbywU7GmCQpDP1CLgr
nfDDzqPebzTD8+edMoENAIoUMxkH/Q7cVWQdfebD2sn4yDCvjyHKrV5P9bluFvkM
PhU5TkfjonFO86Idw8mLSUB9J29RQEqjIoiI5CSBzfsehp5NYB/YFdA7Lqoj90t1
wINWwvSrSLrMoaFCQnBUlvu9Lk4pv23Pm20FSkn7StXEmsh8cxFSv7S6mWSHzT3B
GU4A3ZqWNxJCcnI1+Xu9doHL78Bvda6HwzigMPhxMjDKmcTKgdFtQ2i65CYQ5r4P
c67dEosCkztwAbbqPkFfOiLRfcdilvODSdH5uYHe9xYsjOt3kKJU52xKD7RG/JMq
qw+f0Im5m46fb7x2OJ/Btn+0m6ImmMmyrdxtTL6WRkqu4ue70mAfCcng5SxYuesh
nGDQh/eH6UMCEVzUwDFfaJp+hopuHH+nXYsMcHrlorhMlby1V3CHrFoHYnJMGqNa
oMtYGBblj8wteOy2+EXLTSGJ1QI8q32RwOC7J6tuLJ+spK03ec87hHo0oXGkX368
P9WO4K0owZHnCXUHoI1Y8RDIFKuhzkzt4jVafcNwr9Hh+YiQRlXJ2li/JBv0M9W9
viKuPhQ/3TVBut0seoS7NxV+y88S9PzjXX5uVm3nWmflbsae3diDPJn3Z+oSnBsa
q5AKXkCls3LOS1zu0Yv/pzTmLPefD4zIECW5aH5o9hUY9Kv+RUj3R71EHZdurBnb
ZiImxbqHg5YWDeTK6P/w7wHjITRfDpEJ9NLhk+BRQVuk7UC4dQfUC/Zb1L/lUyGD
P8Qq+8wrzsTBSYBa+VK7lFISmSw4gbcM4m0WZNl5kivfsNbmLLdNEoPcm8wnv5KR
ePiVYG52w12aE+J/L9Jn7ehuRaHrbFPUYZ1A9+N/UXdEX5B9fqEL0mu5eTXxrbu/
3jgBa0P1zbs/X/mLNcb/GZwa2HWjCOh9yYsyIIUafmRqcCMZkh2H01nAdw7YUlzA
cAsRE0YcgQlC3Y7Bh24iA4D5kw6S+xJibDyYmgW37iA7Yik3cd4UWkU7H5s2hitt
ZEVpMC431WYefzLEWxBZSppk9WXZe4nWkh/FdH8f+Z8awSXbqRJJeMKjwaBLGeQY
fwbn3E4WOQBKMqNP43LfPgMuziVKNqThicHC0leaCIuid1lOaVpInLS/Eqfc+Gvw
ERAyBSBestvGrmoIxsl8NrtG8fE3EhRxVsDYdZBOIrTB3HMwdVdNB/zrYgZDIbxo
Dn+xPJuQtNbMfpwA6nP+IHAt+wMsjc7tKlHA7iv61/d2uB5obV9eYQQOf4lVTEmf
A8pW56Jx3p7ujh38p4OiAI7RJMYdAFTO36jmhW4vuWt9ISoCWWvUa0+zGFjFDC4K
WFcNlJQC8qXwwJcBKUxcX5y8AdUmh7xzrWFfJ3LqsrfRz2OpE5Q4pJWRqFbtLnua
vwrzrAW6g1rTpDCIgRCDwY6cOBdyy6YleLEKuICO1QqM1DelefEG6sXpta+tyvOc
kORtU+lNXInnjJHC6QrWFaYUNaWkEVREC0bnTFpxDQlAmNQRqlkAhKbAR8+OapiG
OaeuKUnIehfB0ZwQQmjQhDRdS5PgcCLsCx2OmiVNDA2zSQU7Sp3MzH0UVBemhxO0
BS8kGANI+eM6FSHPsQb63n5hc0rq2RRQzWwdw3jQSbCEYNc+VVzM53430p7PbXPM
fA9YVkKXTKNaoQYK2heoPwVhmk1yl0tjfzqp3Zqw0rAwrtnP7MxsionPuyw21aYL
4isArWqkkdFiaS9slw6qdXmoBjQJkk/ctnqX9POF/N7pWBNh4icSjuiB6/9tgnA3
Zt00qlwWXwJutqjDv/I4h/AZygemwf2302S+vzlidYB2/XD0dJ/UNUB1YMKijHA0
2lZSxGuyljuWrr/xxSXJueGc9/35grypo+Dvdr2D6djx8Kd4IAts3jpPGFNIRBn+
/izoIeJWxdl/GfPFWReVzHgLv9mBzSy8zOLDJIDNinmjiIO8WLZKL3m68+D2LgsX
jng/SybF5RHxKlwWEB3Xuj2tZazBA4YyPUZU57hMzntJa1h3BPRbqRMaOETKUMjO
7MFC45pg310ER8NTf+7AxRwDjY0HXYbhhmRqX+hP6W7rnxRi6/B1nJn1yCwysYZV
Lx5J/VRYNNeiuwYbMS0OeD41WiqJM2X4BDqFPvlLDLYxPRAXthyZHrEhTM5LJh/V
OnlLN7Npx9B4aIEbnHftR0gOHdohZEvRs2b/0XC7p3c7apCTSLbqH7cfKo0DiAs8
t0RKheoDwjgR1FvuiNSUEc63XUFvk1xMrXrTVcE9l9cASFGHTucfGvUkka5YINtg
UWOC8Qs4kRNVZCullLom0XLn5bqRxdv+Zgs2+1JMZyobZp+tim5vgUfC8AIe2YyH
OtjJ2WSQ+ImWBdd/5n/2cromz2YB3uq+8Lk+XacB2axbTVJEQIhNA+movzCwRAQl
HVPzcXAlDvr3TE+DdGqIXh9aEUULOeQsqt5Ho+CDnYZdOAX9QkfbFIgC+c1LoqaO
4S1li2Ulfg8izDRN+E8w2wPh/0p1+jg0uwljmzM7vZ6OJtwdLO5/VlL9UOQ1ZeEk
QlvE9ITwxIaPJ5HyD07Z2eVg7fEUv0pIsvBHgvBxsPMohtr2scV3nW22MaYZmBXD
9k7dkVFs0sI2ynSaNxB4mkcg1DnPlK19H6qSShpZjc9RGBmDg9ok3Ta54R0ByHZw
pM5DFcRn7WZvtbR0h9V3nSJlwVCYTGSNw/R2f+6UvG89iXMSLDz3QUwFgsHT+L8p
aG1LUpx4WamZV4vnOtlhgmnRWWPADrPzwjOeDOdGBXWwkDdwgc/fsgT1zmvaPYGO
Yd9KGJCMxNNmTHG4xaAyhadcAqObLKwf0q0gFaRVjGOTF61Jlv/WNlZDFjYl/5Od
Jhs6dLymuld1xYCzNLUM4otxrDhRtttfbs131z2xooj6u3/xaZJqizeFvA92dwzz
/xljuGmky4MhP71YP3gL4f7InFTJ85wVK+kqLLLI5/nL608JLTSOQbPpbSXkexLK
obvHR3t0WSRQkCJqn/LVbdqMsTLVjavQ4UqF2q7LszxnLM14Fuk6DToeJC7OdmR2
7XYRXZAZ643AUzcXUl4eVXLDukEJV4aRa9ULKTmuL8T6FDzRH4II3381A97OYN5e
fNAq0XFc+19KMERXPIUodlaElAP1Qsd0fDKpWWhoCox0yFCQgbIFTjbgbU5n2kmK
pdy5RqfBppChSw/jiFk8rx2PoAgBqSEZW4FJ/bb6fNp8st2VNxe/7RqKShkAp4RR
qc2FcDJobLBLOo8EUZngbt3wpWibvFvvnVHSaPDKALEwQirbv+DbDMnolzCqJk8n
ag/ukPXgmK8LiASDMrJsJ4JWTLw3cJv1o8CuV7iZO892UioDKS0bNDbPkcbEgnmZ
P9fLUc2kLQ0XmsYEnbFtwvUKADEkWB8vO1eGTEYKj061hjfzjT53twd+rWw1nZiA
GWWKAIXqiP7bWfEdsa6NinnTNtdhX72/2ziAPKPvHxrCHpacA/qnkjsLWI0rzOPB
J8hJ9+WKsiOkdtbC42pXcE+FZl5xFCvdoYzfRKMdx2yXzNn5R+ooe4MnPkJcfsG0
FJRY+jUo6YIPkfZ/zHESfP+4HmLZ90v/q/qwp67mHrNIMQkdE493FWxfQKdCrxVG
lYpsDMxGBKhZw0pt8VtqfFJr17kaqv2hOBKG7XptpIVK294L3XdpVkIiGozuUV2/
MVzsLQWimtz3smp8CPnTvYIR+qM6vOZ0aymYBSArNrZxk/e054R0ip3DMbOrjFLx
U4R1OYeXx9knd7fNcylqQv5wnEXcxdHtgkZ6R2J2lZGwzLFdYm5We7CMPSkRoxJn
ZqTta+LrXIviZWJiTstQApSMprUl2vPjkbwNJ14ZaoYAfgSJ5V8HpxeYwDDeoGxK
d/MC/ewOyq/DpdBWp1aNvJsWVv5Z5Nee2xqp4/s1DT10jTmP3aK60a4J5sWZDB0k
+iox/5jNOexYflY1ZwBfQEpWfG0e1xGGxfScWxcO68rSIyxB/9q6+732klrUXjX+
jQDBDDYlY7Vf2gNizUpY5RK25XfO9OOSWbJinH3vEjldozsIFkDS3vnWn2aOtFpv
vD6Gmy9iHTe9OCRnMoWKoS4nWalG6uFz7d6YGPXyIql51QiNzXzjVuQivO6CCPOh
LmzAJAxHFJlhEkTOoSEZGnS8G7GdXiAV0/4HAvmlD6BuTZElg1v7SwJi6n7M8vgz
HN8r7M6JkkUIIwJD51rgzVEX08LRVlzJC5CswuICBVjRk/vR3MRL+bfne2V/ClA1
7RxL6SKsP874bUk1qgfJQkIuW1qbq1EVvSDetNaAMb95kSf8rXyCCDdEk1J+urlt
vjCDk884VM31Iu9WM/EqReHNCSOv9yDPS749Ipbx999W3XELq5s76w7TCPejdGsj
B3iYXmB3uKbIwA/h1XFXS76XUf47t5SnzBqxZC4cz6Gj2j0JCUleu2gKr6KMw4gO
oxVqcavwWx0esj6679Uurgqax1Vdaoo2wWgeDPDwtnUN3RGNprumEn3PMNBN1ro4
/I8VSJ/x2hvJJ9QzP9UWL1hyNLfzfSqp5GEa+qq53R+FG5SschwPeHxB4Mtb13Zx
39z+DKTMmoqaoEXB1mAwqmMNYAM9a+mMOtj+GMOfjGNWSewLolTY92Y5jiPQK8d6
K3xXjeK2sXpwZ2pel5fvyhAJ7tTWyA2NJf1OwjZMT1hzvADr3zc5zDRrFlUKE0wB
/Z1xraRj7nTUXqQ3/jrTH1dn4ED6eVk/3DtxVO2U+BOA944VLtNmoDAuPisN0GkF
YB/6OgOvfLVN76YH65jyyJVvFE6xTdmS7pDN3bOF5PB0iuV2HEn0SN4d70AoZVB2
3CE7YebbfM5M5Pp20/T5M6Rp2cHLa1o4LTJ8Sfrjkb2b+TFgEquiJwZwrbfiWt4y
ghli6dfocbMaknaAuCgKA+dAQP/cfXK5z7m5YTHaRlSGE/SlehPdD4H22+uQ+lyL
McH5jD0/0aKTBKzRqOwVMLD0I1fldSmWWJylmQbDTDEhuimcPc1w5BohIBMCisbh
62znZUnly6HXEf9N5t7UjG7EwBMpmQjEGUGaUHG7sctlT98garPQOseKTj9wkfD4
O+ozFie0bCPI50/qReY8FfFTdrSCt2aVvocG2gAvscDc1AHXdf6U2eW6D70H40bL
9KhmRJYD/XqdSqY0s4WnbTkGjqMYsx1EP4ZtBrgsnZj09fx0xhi3pXa6r44z2B9r
8XLASaETycCUnbOiLUZl0N07PI1+DjtTQg+pVPmNxqxtevQVpPS4X/KMu714LMSj
5Ea7xpAwrU34nFM3/fn2yfh8E9rxF0YAx494FsOo2Qz7PX0aj4P+dsB5P0NsBHNk
TVu0tReYZ03YBUnw7LYsqU/AY5gf1ZSCjihP0F+FuKYJm3HDgAuPY6ypsmBG9gG/
o/KhY8yPPQMdVR/DmVaJRsqRPuetfC51k3Mkm1NwUKSgetlXkUnoj66Ugzy4TOSm
SIQ3xhvFfLcz55anCLhPjdRc8hYDm36DJSRG3HqhrVVoVz/vVRivMr16AfromlrY
agkv/6aAQnx3zeBIJbrzwohBV13CD9oUPFI6IPsjKTzaI/L9YDGbFqUL/w+eAq8v
o33HJMXBfEtsLXqcOCF0h6TJ2mcaipRJX711N8Ef0cubMRlVkH++K8YSE2uBuHif
4LwtfKTrbbx8/OtHyWzjVYVRZasmjp6hiD5nq2Mi6zA7C2VekSlXcINorpN9Zld8
ZTEMzrriusj/of0WGqK7emaqv7w+e8O1bs3cnox4pNzPAJSXcwywru4k3qfDSMS7
exaDtqtHZTCr3mHNnneovSZLR8/ZMiToIKOcaZFDdXUcFMPnSFpzGJxVIU6h6889
M3zvnKoonVgZsrteRFt05rXyQtIcusaeBM6eMDyUV9u2lJOHq69bQ+5rRdvAb5b3
InNGqjtFxnnolLkSf68cR9jgwxwq51v/FXHSHhNrj8J/aJxYMLHUpPsWDsfwm6xn
bN65DmE8li7SRMr50xJ4OsHJS1eBvn31bXpImCAG9/NyaK5jfVsdLr4gI/gaoE3w
AmZwkHEJcsvUXsEL+n9MQI88+BMpywLRkRPM89qsZl2fBML05hMdSypSk8aZ2tT2
TdqaZyHqNYdcK1tYxAt9p7jIr5v9MU7GmF7DsudjFOecQipna7teKsuWgNtgaq39
MmCFB5RN6A3UqXTNv5aX2RiW704POR6E/ICGsaUOndy8NgvyD/sNpTx9jo9CNtMG
lF6DD9dvdoRk4Wo27mTL//heQ1B4m/fCgyEcACDk4X2QxgKu5JVKkqhXBOPGG1bg
KeceSbrGoc52RwZ4pSL9sI+Fw+cW+RHnBGI0rXLpPpbLx3nJGgYZdX9/P3sOcli4
HjiElFWwMrJBVfbHQOSfnGR4LMZvbFjOWULPDlrsJlg9j81LEOGPH5F1tX5IuK/+
rg2XRZItgFdVVoKTUTOiAaRqM/w1huKXCaRUbjnKPgujZVkrv7jM9kAszqTru4Zu
/fwYaPBXo3YuGAAquPGBS0aT1iOqTnpz9VkiF7BvpvPSd/CG1o4fPz43wkeN9p5h
6sBr8FoA7o7KZWRTYjR/D2mw3Lrs6p372fFPXAR2xT6qkgx0gTz6UwR5f/XWmyiD
flM1Kr8fcZTu0sdB1mC6v5euYDwMj4H7cQ5WAnprPQBs20gZ9HR+RSHuhqRN41K6
w72LSBLWQ/rO1746kH6a2fV/WicudDz32BphcOr9W3vbM8Aj/oG/5txJ0bnwBpPa
wNL5nW05SH92nCvFNFLYMkkKKa4TaRoR4EfpHDp2aRWDOVgywlp5GdwOXJ+i0tWP
4L7XRCgQe19SSCj2GfsfcwR/R9r9fo0od3LAAOAzOtJ3UgwKS3ujnnxATrqFGcDk
Q4iW6dXeFl3b3l+H/UAQq1lWgI0m7IH5Utzht/n28ONGd7qMaL8sl2CLJ6/pc4pQ
6YxkoCAwYHABJYwx5LYaz51iudJcJ5h4hydOZWFTIjAmLpAjYn/MoDIyubgRMRfe
8HKT5tVwhz2CL9PfFusR+kVtgnBLXA5AxvXh789m9wbT0YJEGd0pYJ9WuoemsPZn
L+dl/HVHY/uXDOq4lJuLXq4l/RUN9scFMM6xAFz3YAS1ZrQN8ZjGa3X++nkC9TgK
H967Qd7mWs+gHdXVO9LSTuW4KC9i3+j9gsPxCHPy8pLh/hM2Ana2shstfxj0aHo3
OmTsvK3ugUws3fY6DDsXLynKmdcY+qg6COMVk0MwZxomQbHe8rdJzPqcOHSK5vz3
enYsIEdetTpeOhe/ZDwmQQkh2tzBc3s4KKBZ3WawQofHI/btkrSnQUtUe+t5uFfY
VWXQTmA0SezXgUGoO8TWOnV9CS/WOZc+BK7TmB7P4SQLxZ90F8twtNmhRdbH4/cK
P86t/vjZqVH/PpoTaMPM9DdztDRXblJ47aIrX8a5IqIReT/d8fI5sV7YrI9HM/fv
gg4uTPmgsCxy2iXC1UBMDthTKb0xFXjgj508IkBWZ4pATdxDgqe+cp8tOijyeQIj
lB8QbyQMaEliTC8eHXnS2x/F8b8S7cV1lEX9tuZd3IZjMI+IuclaBRtUQQ4ae7AC
yGd4jfGqquW2zXJ97Hog7d3qGzzEQ6qHkNPdTsY5Xk7bXBClUKfZHIwa0FurCHGQ
VfxneIuklRf23794YuU1r46tQrq8Vtmf2+2NWXhLQxyuyb2ySnJJfZ38x0jriTrI
zETJT/QctSgcwvmgtzx7YCT9eGvPsty5jZUpiqcUgmQLvD9gmwR178gDNXAiy26q
2gYD3BJGNxBoWQSV7VFhaFF8Sg1l0Z+iq/Kre+Gd6Dr3jHMFzok+J4ydJmrPgZWg
qsYeCfdwix+ahntwzBEdEw25kkzXOzAgk4JM7o1P2Dz14WjigeiaUfyKW6xaPsy3
s/rb8xLVlCAiFeWEqM+Kma/6ujRNzY+2PbHgbqgyR1J3Q/yMT+Lo0s6ZkMcDC7Bf
W9Q3ghTEbf+seAr5cx8z4fDbV94OpbImjfKxTSumcyYTSvOSMOCzbNvV719Dg0A5
m1bw8Gu5xtOksAAhM+EWl560q5P2gGpxyaQYvGr/z/IP7acFIi8rTkaeC433oNUB
ecsvdm6tyuRZWWxJbEFESJ9B9GlFmnMxds2b6IxZ4vHc3dsgaxHULo0KW7+bTX4x
wLIY225rZ8zcjBDZP0ZNXR/LmadyC2iBuTeANeAzMXBh+g+RpnEN4wbWhalamY/o
5C67mNqwhDCI3EuX492keRFgunJ42GUBDKh2tPOPk91897hgX6RWQWjNmSOeII1U
bljzdgwMFeeX7G+ClibFrs1KfEikr/INt6pBSKVTxITtcLE6izslKUjdo65IUvft
ZmX+T853T6nwJsJNgybKtsDvO3Vn7qTYYhpljjkW2FhJJfabX++oYT55Iz9zwrv/
Ts/TlhIANynwHxxeJFYC77G2UOtGBGt+GvZ0xu1zDNhLwh7+USG7FkOhgozYP3cG
+47lChERRrJljZdQxAW7PUBMEYRiDWi7q7RZ3/+vjoxdocmuFbV5iAPza4pHvESh
/DzD3VJTTcvAyjqakGuulKLezBAdjPYH4j62oY2L5KK81MYSnbX7cfo/H52RGAHw
VEFtCPb0tYcpzXGPKVMUAv08b7r+TcmW9Jiy50IksANtEsoA036QpZXho2yFeAct
sTyStvgcCY0XHe92Vei/1R3Fm+5lAGdLJ79cr7MqNiqBxxh9VOEeBCCRkzG6mM9f
0vu8WITSeUx+QgwG33pFtWPFHX8kGpOmNeU/dxaaiSmQRJB4KT3pwRmkBIAoX8Mj
naNuOnAlTmXpGV03ymIzmIKEIkwfLreppDAHKR7QiCnWeXIPO0vl1jZooqdtnx1O
oo4u9VCJQ+Mipjvnm4kxeV3t540s/LRnUiB4Tni6Ebzib8K4mqhRgaE/6cRVlWat
c63aOUdC1azxS10vN7Fje2KbPiis0JwM85FQpSGEvCSNBmnSTP5OGE6Y8/rtkjbw
gml5V2DeFktxmUnxbFiA7odyqeDbY0SZSvoe0eKke1hp0GBa//YLz9QxHy23Woim
gjnNixHqxuxuTS5cS+Hf4H0/9RiKxrcMoQgMBcJtlwJdCQ/04461EgQj2HGbU3rj
whhuBifspyOPK19rQl+UkglET0TvDtgcn6ObbfT++rdErU72Eq3xATLOrPSf9B1N
`protect end_protected