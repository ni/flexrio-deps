`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4816 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhBNVMbsl6PTB5/ApNH6uD+DikcqmKlY6aIDJdxactegY
AxVO9v0riIv3Q5ik2YxLJOlL0IidSVjGCiQjzimpEG4jKXxzHibLTOKI+N8VHIjP
pTj8N+4qNvzj2hgWhi1h6yJ8Gtkwl2/jjWP1ZTjqutLaJlHJj+4gux7sVmIEqDOA
MhDx/utau0E/i7EHoBbXTvBU7saBdIUbrSe+206wSQCJ7ZCUmH2COtjSEmwIOtEI
wHO/LNSLvY4DlVGY8fmsjewwIGwuWVGHIHZ/eMxnNy1Dl0ttnbI4kGVM83h0XhtG
z3oMf86GyXPUSxe55O6BFPrTRWrmRMLG41JRwLkhhrxO21xgXUQ9FqotZnMmo+k0
ZEje9WKurIE9YqwWFeDpckKq0c9tbZXSxtgu1Jygme9V6oI/Cd2CVRVLhabsGszw
bKhz1kF+xgod8xIfw+vs3lSJbNG2bTw/p68FNcsNGqowDVqkXC0DmW/1jMqCI5qI
re9te2SedgbRVBBmW7oo0mGcxcqTiReSfdoUcqQN217HjSsmpvpyXAjT0CGK+OP5
ifXITMDBZsBuVFO0L1tHBTce6PR2bsGxUAxjKK4lsOmSnYtCU5eme1XfGed55gu1
iO02op5Y9Qg89G7+lhHDzqJPtD/rT3+dTFdBifEm+DqWj0x17smczdEUpXrtrw1D
D5cEy3ZOVhqezUU/qRA3CewTSEaGFXRyaVOXHb07tpBsCbcZmaVCddbUOUamEMF5
0Rzgqpydou7rpFu+k3vZlS4ss6bxcOT+w28unfM+qN8/plNhvUJH8N2JuTO3NiDr
bFntamMSvBTmGn7OkV0Gz7l8DGFO6u3py6vcl/8Y1oPhaf2ML41aJ9e73+KufHCq
SD7DMNfFq9cKoYGgGY1W9EHzBPUhd3SxtxhiKtu5Lt2d7efSY7NTzfXRswzE1h+M
YVMUkO7NeMul281af3kvdy+o7LSwBEm5kvWF6kj5dXr8Cn2gkiY8DyXZLt0wAzj6
uKNL79rUadvGnuZWzgWlwWEZqayZuWc9pxbecfW1AocCMzVBfZ7hFohQE2V04IMS
/2uilrMx1SRm+amQ3lwoXLR3uI5BO5oMEap9Aij/HEoFn59nC/1niRKmtRJH5dLa
f/V+hlgth4Ih27knVjStXMemPHSPhVXeD4ly8PpSeKdQxhW1/68s3FzI2v8gD+Hj
MGO+ZV3NMaEENtAoGwNyYlHSm8Gu2kA4TzaeHwsFhoT4ATysH4rTT6PMK1HfTSjj
B1yMCmDPBf81Xw1sRpj7A5Fh3iAe2YMXSHLh2UP4W2LzA/77VWZUQgBg83srWJep
ou6fhkzdziSI7Qm6gVuK10+Fjbw1EnvpUWLo5uEh7BFrP6bj9WnAMZT0bilCu/lp
n7JOcCfw2OMlJ2+nkjrlTujW+F4LInKJHvWI7iKZw089etx8Nk6qri8FFNZf3M5u
ZQ5HvIvjaHzEJ0gQ4QmO0aq+MIJebZOahY9TM5Yr73QIb/VGpXgYFEZozOtylhHS
x8IUg6H/UNQyxih/EZHOOajsoaSsdyJXR6dLgWC4XWoxokuEc1RTeDnRKuWBIvpy
cZUt3bzwik1ng/UAiuI6RBlIWUS7TC0Adm+OMFBAVi5m1D9NI8xwUSCSeQZn0LYV
lDcynPLLAxADdahihZQh68xg/jviZtUDpRwJAo58zWxWjvriHCxRZYaz1WLvrrIT
Jq7eFDmVN8qUizJRVOfh4BcVufQ26t4bEQpF0hABiyT8TRemZXSw0s+Fi8F7tyni
ezwIFFRTr7P/Xh/bOJ5n5WgegUMxrWGgAjsOLFYiRfFTdchtv57y1N6+doiJ04/L
pZE6+EQZo7RpOzVw7jxsOox9+OGoCdaUpOsg0a58LgWh7gne+nPGABvx5GsxXUoi
aNGfh/Z1DgH4MrRlsIWVVozc40Gxbl6kOk+1cCvQE0qIQhD6GXDNn1xeSQX+ixHh
WWCxveY8489aoyIfhskIDS7P6VgblcItdOS1Jt2FZvIVRmoc86Z62YqZ+/ENBihK
Dw9x1IPAOtUjEFGJySlV/RK/TuuiNfk/L2+e14mx+utBWVcWK96S78JXhCZlx9QS
rE84r/KaJ6hH6oIMV1GJ2GSk2+DD95ohvbZKpLHvnCct13zx+oskFYprEO4sB4f1
07o+d/hOkgtGEzrKaETZZbgK62jqp0ZEoEK89Wx2TuMXbdhTdyixQxo0kEi5k5Is
8S1vpP4gDHPO4VVEhHDQWa/UqWzc1+Bg2B3fJ9Xe1bv/OWgA5z9ZZNmsr0kmxN+X
N3DEsk6jEKi7Auyv9AZGOxWUO5GZrCajWZtGJy5eXgaeJhcCOytXq3MmH6oFxuOX
+yYsbtc9p0N91Qoq/Le5+fBp9LnKQMDIqsPxrySHf3NPuHDP4fQXF+4VzhLB5giT
JCryCdWmPlYIsVckdibahbqVbt3IIqMVsUVUihOwJogr02kU2HUBjG/RHoHbYJnw
BQdc6PZsVIYRcf7+tENQ9BtP9Nwt2Pg9csSdyXRmvEeu4pFsiLv1Xr9aMqWj7vY9
c+aNatjmY+IYMOgnf8UAlITWuyZWE9C6bOqiXCVEg7gPEx3O0wPXYo+PA8r5jvid
YgycwRluTzgCU+49dku47OmzwlITmghZ7zldjTGp18Ns91g7xw3naavzC9bb0Tev
3qrSk245zn5x9fPPKo7R2Oo5hl6ja2AYfkxhdHLJDmSQNw1RvXxC3p6pFctEcyzT
h3RpvL8BhOXfJxXHfWYD7O0vqE8VlT8jk3mSlk+HBe8ZIF1ZJf22AB96PvTDGmW+
U33zm95xKhCIoiEPR96WPaX//ed1oFgDpRkfvFGzwl+CKevkpG1aKRUKLXqr2W0l
Rsd1XxWuXF5rM4d9c3Nfy57xjhWP/za1z9qaYQzTgeptxvTdeA66rxbf69VVskue
v+K0JCy1icF/XdwZkmYgyQ3pw0/UqLz1PM61xBtoddVAXL4AcgLwWblZcJZ3ys6Y
vEChsM0Vl/IGprTekfhROFq91ssC5Pmyyx32xzKoy815TVqzX6wuxZKM9dA21DpN
s0u0bZWw7/QnxI8muLQXjn10brow5OoRyQoTnE0AsmcB+XDD9QGO03uLNW2z2O8P
Am8n2TXjFIKwBya8ZiOQTKBsIj0bk33eu7Em4huCK36NYgPiVu4ZGqNcOB0pNnOn
/mwnFUNNysrQvAg0QxLTc1O+TfjNwKWD8h3gvVBUOLc2Xe/EFSC7/0aUzGBk/wG0
HDPZg0ugcxIxv1YmXPFVJQYG69wBEaFjpTBTG9/VhLsxGU22iE9gA9e2rzjySes6
7zeU12vc7s6WDFRohZHT0AHVN3XhlsUi/WRoKa7JXp7c4TgBfxaXMt1g0mq//OqM
Ud4JYaiMHDzECu1bbSt82EN49Nxppwg5GEHnhK+GoyQfY9lQuxL7QINzRJdlKHHh
Ti+VN2Eh+ZN5UVixD/tYkUcBcPo9HKxj7vmk82+Ta4PXZPe5Cf6zlVv//4SIi8Pl
E0OaiLc4sxaESwPBtY3QJq0fpCXpsIxP0Tcrgrsy7h71TKITNVB0ODEFPJUUCHoT
CIfpK4GCGnNWzYHQT4/pSU7l1iyj/VuK9E7slyUlDyZH78HovCzGPkh2tV0WqVKO
HWSkHsxG2RY7rHf7KPZFZFx66vgb+whJgpANJ84DbjJYOHoOOl/RWoNFTVhiH5q0
7UeEVuOYcd9oNyRYAQnX9pUwzGZIAbijJnWGAJTlhro0y/DU3RHfaRNQxSey2Avu
ZThGcvj/UNVsEzj7BwJVPfgP/eS+AISc/b0e1NF1clG6xNBZkzZanFiKwOzDZYsT
zvLhLldUwZafmrDa9rMleYa6XYuxeJOByoiYA6RwU2lWc8hjQAslZTZYnFIYzqu7
aBNPQZT4JE6Ygbr+hnf3xn4crbIpm89xdOIA8S1lWxeGgFZEYh5poOfC5ObMC6ap
BlteXoAKOXrCvwki/JJeZLsMONw3u/7YO1Qs2o831wAC5wvxBqu492C4TWSCEzU+
Cr8rIY710D4RK3+WzYGqsYmZLv++CI9ZpwkRVGYwIRX9mcTZ1b97pIHXiUd6zFNl
oqrj2PxNHijZQqOvkVZFeJTUjWd3eiYTM+rvJ+JyDgRPHoxKmLr65fuXF/k/QHNa
PV/+Nv1vLoCIYzRRywbtBMJauXMgaVkTAgNI1QpEEHRLeFZ31M1CsF84kLMTHg3P
N7vRv2HA84iJ1LJzuibO08c36QTUi5v/Z+C7eRWSM50SPK+TohYRvrZfyOImYamx
s6SuasFhJdQCOqDZ7+ZPPuNns6Dsk+7By1ZPI5bC088n5+111Yn0L7so8UqnQYXj
8+ELzeZq5mdwcLk7hjIwdgfYAVCSQDIjebzuUpxLZzB25idPsQiw0wboziC8OcCW
DvdkQbJlNbqPS9qt+bLpRLXuHSRellVDDThsIGPBFQ/Su1nJRrYVddAa3O7wU+DJ
AkZPdx0LfWro9lxG9xxVmdAlZweIwocmSro19gLg8ff7l0YlgV2yhvDjwYPOm4Yz
lnGuHdBcGBnpvTaEozTXRQD3mBQSuwlp7ql4NUNJv6ITDpv+bI/WbcdnYddyzBcu
t7Qx8ej/fs5iYNfte8Q5JMKBZiyOIjBvwhvXsblw9uJKyc9VkHtzO28K+EocCQia
AxstXxI//JdiLP6RQNEF3qr1g7zUnHBNeMAYg2EIMAdVSvO6Ywlwv6wAMcLJ5Sb3
sL3isfPkXxaxsrsaO/M6jLT04rD4IlkfLtFadujLgtSBeQiU7enLHqbVxKwvmD7K
cztp9E+qqUbJsdDNYieJJGf44by5Qch6h8JDQ2ACUdf6rUEFRW0e+9ZEp9V0XqD/
C16b5/saclRwObpdywpxIAmMKY46DtBzaYKOPobr1LggT7ELIwogG9YnHhJv0wYi
wOoZiTy6rzigKmNT8pchGMT6k/lUisZ9YqUlK/abeqAg+5V4G6Dw8++g6M+QEMG+
6URGWlUbADFRUMBfyeBMknfJQTy/F5esUspyZtgrFTWxaTk9BIUQWERT7+nWWFav
0pRaW42GyTkD/yULVb+2P63c9/+Sk0rVwKaL6p6ebfoz/PIuT9LYn6bdUtehhi+/
D/RTLIlNECrMIJb19Td4t1X4UJGIfeSx+z+WLElgviTL9jfJJRgCkbiwrtABC3UC
+c/NLdS7mPvXIc2DUwzt/OFa1jLS2+Xc3qbTvUd86aiD357xbxe3pA/UH/mrmGWc
5jXwPyOgEahJ9tlXFa578SE2s3QAiHzTdulyKHsYC4qKR0IAU2p7IjjMHr2nvHWZ
gGbnWi/rarhuWSC2xm+lzxDPMYJkqMlaqN9qyAmtucHInO3PAMTBACTwklZRziX9
Rtln32ZOfR50x0iJ5WOWp3OoYSeiCQkCtgT6ZsRpksEiU21JDQ9YorMhWEbYXLEo
0BZtcl8+O3cNjeSXpE15HhfbEQwVEINKhO+NQPzBX9adjftZFgBIooCrDYHHYusU
U0Bqw6fPUiX21KMMRsTy8OcH0YjaJ5sBWzayN7Z+DC2dOlGslYOtW+8RXsbpehxL
Oc2yTYr2zQoTddN1670YmkmpiSpsfLw5Fzc8Oa4cm+zPOa/0VooLs7/VGtVeqk12
isvT93jS5kmsKCLuvGsLSrOmw+OtnH9lBwXd2mqYxiruoEvfNJFq/R1zWTXLyxwq
5HhYUsD99z0zvVn2bp5YfzZ6nNZu2MvfWs1PAAzYuB5SIohv99cVRUInqEUDCp8R
+ClGZVHS6N2n1b/X6byw5b4GTMpEoeRtSsq/PNnCUf226C8IGQmfRUt4Muzmc9LS
y2II412gf8jkXZ//PyY7Rp1p0cTgKzmEVU8CwePGeA/HUC1I5GJzw0ps9TEQ8z55
uaonP1zjvWktBPquwluaQM8mId/H6EIc7ShDP1Sg/18xv4jbVb30H3fD33Kd9FSu
xhD+l0xs7NnpZg+qlmqsCXoYbwEI5YgP4Wi8xQ30lFvtHnQ4TsXJcVHO/NxR+BvI
P1idoKuHMNK79cED+RG/SIvPy6h+R1LpPd6oQo8pMg0iAWRVz/1CQENNavwFzpvL
ABAlivdFmh6DTuwHczDdlLDhaYcfmJadB31siAWcr9GFfFPdVi1bHyWUCZ3OgWI6
EiV7uMHApoYxykqcw9Un1w2BlBBq9BClmZlhFg/fAyXv7j9HMO87jjtN9XunJIu0
/twj8DT3JWyPwOYqqroJ9f4XTwNP2DCJzObFKWT8d3TnBrKdDB8WDKWmi8ygMx08
q9YPX0JvhcJofIrHBT0NAw==
`protect end_protected