`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
YATj3kULTF7Ty4ORuRfFpnT6YIk4rUPRrM74bVTnc4GjdV8oSnW5PtQkMCLOi558
1V+/wvDfc3y0Z8//ksX8sZm3JZWtrxUppw8c14g9Y7owiwp+JumRtO1zuk5xFbe3
0MMnIxxoTKLhyRJtAxElG8sbx8N21OWDGiOk0Xyd5CqAmk9dcOIbxzMjW/wndBXi
maijUdqS+5KiRCM9+Gsp6k/iEAa2LnYTt4WtjkmDD1P5jZKsiMgFck8WOqLymplZ
ml3TTfn1UlLNm/+zD3SFGP0kABAiUT8NK2xBPQ5UzQ6sMFPd/np8iUZ5u4QLTWOZ
hTrU9OSX7lOvRUo8pJ9vPg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="BzW6NOo8eyBw+CxsNNo4wIDxODIsVe0ft0K5tGuSUZw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
DhjJh9S2BY18dG77XPz3hsiSQ73+w0XqfJhD+f+lIDHHVjOB7CfC8ieNRTexgzn1
5W+qoqOEwenoVQtit9u3XViXJSRJ0wfUC5a9axblRNyD2mUbyfH9+f59nWqGkVOh
ieHxkA/DPprM70F3APxk51m7/gNSLICSvbONgLGndWc=
`protect rights_digest_method = "sha256"
`protect end_toolblock="L7NTNW/5Dqy+2kJZXKczEa3js87UJ8H00YWI+92sDHA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 55056 )
`protect data_block
6eHODtGLmq6ccbB074dgNWpdzW45i5jL0Nzx5wwM+RA0eeOHXxEV143NNyQGmZjT
bzHAi/6AyRCB4X9z0c4MjyrZE8GF4crbMH4T59xFHqVrQ4zXCea5w0kG5yvHgpKo
rwIIbW7Xn0p+GsC0S8TZEs6lC30gMOR044cabk5vhpL1bgF8iZhI83LKRJXvrfT8
7Iolr88V8cBIaCmqp8NnmUzTgu/s9CTe7zcbsA7Me/tVlUYUNGJ/Cw3MkfS9fd4i
ik0zXQJVjxvfAHm6B+ZdcGGUtzbzJ+CCXomEbIGx4T7dELSYZs1Ht4BFQ8Od8Ihr
cvNscWMohhMh/UZzLgA7R0xGyXcHslSfgEkt83SqTldSmw+f0Cqcum9hxeUwR+kr
wSqUrsZsG53j5//8CKLnc+z3OTbtkUg8STFPVqERU2cSzYTCQ3TW92AxZUCk592l
pfSebY52Q3nP7P1+sKqykZzoLkzPg3XX3zoMAnu2X8bWou72D/6eRJGk012p/opq
xpQt6SIoSGaWv7aUoLIv8SCVGirobWWpzUc008l7RHMKuK80mOxZSg9S1XIk6w0p
0gctD+YQh/bnN9xLidlueIW3U9jclBMBtUZRnfD30Nz6uPiMR9ra6FCiXvcMB7iN
NqTEtA/8LRPK8XmF5JtGzoVV73a4VDKaGPNQUHSF4sCsw4UNLY1siXCpjCgQ2XGM
SA4fju04jSKLtKV1Zq7lyHN+zwE37Hbcuy7sIzl3bs7EUaf3sRbb/7t9xhqo2/Cv
1JEcWgtboh5c1vgkCNdt/n+HouK+gg0IwImiVtx2zGInC+R+/WgSNIY3L8ryoiac
sTkd8tJTlB+ThDsDXcBB9I63oxIEFoCIe1S/WQVXuAAH7M4NTlKCKa0Bm0vZNB71
DsK0q6+sAjsAI/bwqxxhKY/6RO9mSQ1K3WIuvkqFfqAphS7DKedRSQJ17x2S4+3C
FHjHBsuXruA7kQrMLWD343IwtOtj5V6xjwPuZMo44mPR8Lz0O/XRJzl4fZ73/8Rg
qlr607lDmMHthE31ZxwMObFI5pyzYA8snm/MtFf40JFDnmeHUVHAUSJYnCLUAQ99
brtbjeP2KhuV+IAIuFKIvvGxM1C9UWXdBJns/US3y2uLND4wbpLNqrs+5I5Yr3Iy
m2Sm24xrvbde6OKvG6FD4jmkwJwI3RjvMaTUv+uJRGzZWhbStJ5WnyJu4+bBfULH
khOP41utOBNQWd9/n8qP6IWRbG8q4cqVoJ5V5EI+WYatP4e8zX9qnJBtYWGxMgSN
CUgPfuzQCrXauCvA3GYzq/CtsizIeoC4i2pRGu2n8appo6w6mAzVNgPttxy5SFcj
ClCqmJf80+IfRdNJrk0tG9BhaWLIwg98YTe8mw++8y5o1L58PVeGasqJkYPdJ59H
ooZIfky5wzjLpvU6p3j7cPAqabKDOJiDsP4JmFGIWoyv0LXWc/0rNWDI/9WBCLQH
QYe7uXVey8qrYIfYEeYfTWwvkeh2hRfIYWhoEqb6RpXomqQEdQk0gUD/K9ILEAEo
fGDwqWXXyK7PB4MAlLnKNhr5Ak8xiccTVtalTRLDj7D0MLLlu97tf5PU2JeFV/o5
0PEjbPWgIY6kR78HPND0i6Wqprd5REP6r7yyd8C4MJQEh78wq4RizeyG7AEuQMSu
mhmeQCuZ8q2DiiWThYvOIXEkofVBdJH2NVyQjtNUqhSwl73auDLgl/z7uCwdiGkR
vorOBJ1u2Yr4rnDESJz/5g6cDiuQCfZCT58mQJLlPGWKEZPLvVfyO9ICXX5fpBbx
XUgBJkrgR+M4PZxPqwetFEurJJCp/ddTbBxNjjTwG5JGdxOriYQSQ3s60REc1ig7
YxXfpP2hLhAcOJwTLXM2+y9dbUzlXAUKwH3+oMCiw8Ob2ldl+iK8valKbw4hpOV8
WKJkFE+BzyfIrE/3PAA/rUMxB++J1YYJhC4pHcFlMSflVMIH4oqu/tvo0hnrI5E4
svGDZIBuTVf4+q3WR5l3MX/kGyhsPzQYqGRV8rO9qb5Sk5WO/j1AZVjfUHsUR7O1
q0oHlO3XlmSGSHY1qgGs+3erDPobQZ4m1Kj8kOGAOX1VS37T5fAN/+HAkknTZQNC
dwMVx3NN9XbfDFETHDUSlwrQlgenoJFfcGlw3tRymKninURc1J2EK+/gEIh+vC8N
gGqM646feFXRNlD5YyYpVsckzUFMU3wc3K9wrtYcY3qLeZcvWo7rhQGo6GRXdeso
FEXQpA6wD/HxEgUlmmfJ5i7SnZSI0taSE6F7QLHDRyAeEbGK3X7PL2q6mtBpUPdA
LhiCEpadwhCZ9F0ll2H8qhUe4HOJzwR8sltywadP4Z5veQFn5eMPw5VQnbemdlqw
m32OEIbcgnHZAyZnSwwAgQ5JuXT5n7/IGQ5gxYZsFRkYxAD+KHDo2LTS89lK25CG
a/OGtGOuiDuc63Tj2u10CB3VfBWB5MvMaE0E8GALksm0Wc/prUc42M51NRtucgwS
KDsEAvdLfBMWOl22xuuluuzu8bm2vLU23y8urqlXEJcEd9t9LmQURBK0FZ+w09NS
gvexIE2Kx8V090QA395qxK7YuccSQ6ILPzgCyjOiyXSLUj7h5OMvc23kXEazZTL9
9rmeGSt7S6ySCRLSNFrPgzOsd/njgEWdpN5DBVKHxS2nujm+SenwlXsbx7aJDo+7
WU/F54WpMqucn8bh2Hr1E7aZvLpkaZghSlpS/G2s1Z7N4vVGUh9qNfBt1oQu7fxX
Rvff1c/S9j4CIatSeeySTZMrzchawTrBZ0gzACWusWZwEh2OOmOBo4NPy0FsjOfG
iAwAV359C2AvaOXiaTCu5RfUBNLeVYRv+9n1AWCvpCJGNJwY46NpJlsCYKzDiFGy
e1qFPxUl6LoYNKiiQVGwMPsXe9I/SNnpt/7xSrRZfeVsC/y3nc4RfPbk6iSB9clc
2lb0ltLJZfCElKWl8QOrpYhoipmKIPnyMuT26HikjxGVOj7NauJcl3y38hGAUODc
PKLakYFUUKjBfFgFo+tjfnexYjT5ROgFfYxwvclSh4xV9JOviG4MurXBvCtmOSF8
DQQqt2TvVtLeHagm0etNjyplZr6NY8UwEeomfxKtgpWiLuTx/yHEDKUFNcdHTid8
GTj8fWpXD3EK6EnuLR+ytEJO0NTJ4zEN7q+wLYrGsub3H0g2419Qd+6RK2GlyCK3
o8LXODAjJyaSjs9SG2YFpUyTAv8e3nbCgT7ybpRque/kTvsHDpmmFt2/a8kJ4LWc
oJQCF/ywWQjZxf1/kmtmGcTNvXH+YV8OK9SxyR8TbueCPLp0XSKZ13z6x+NsUnEI
fhGmw6HwxawdEc7bP058OwcVabM+5hfqa+774r/aH6XEjAAvhFX7FlqogLD4sPyn
nX+XkDppyT60OMxdEHqw2iqNUgvvZhmoAetjeb3WwVlOfR5f6Fw7f94rztdFRPh+
hen1NOsbQ4zgCgb0MUSwCTh5AiPgYk8X22QCQJ/izypHA35Lu1jpp1fwFf6HbNbI
j2qm7T8VzQ+1TYwcL6sM7uuHkvQqq3wKufAk5lo5HdfghV7AssLRnoOn/XX7zYpa
rCX8xAp3/ym+VZrpjOX6/hFB0x2Inc4xsflW+hsl0ijmt798yN7KgN7vrBoQ+17E
Hk+Dz0UaAP/uOIh7ArlgiKCNEJxkilalHMivd9q1Yi3sKAPpSYLwWGETVcVl3T65
iVH/GM3SKshyyOfuQ3E+V1KHWbF67QS1KcsVG8khhH/Gmv9KBLrQP+4Ebq6XhaY4
IhSDWnv3WTYgUMZ+v3oTZz3obfsxVrcFWpMIREdugg5+9Sa9Ue1YkB8PNqQ0ewBT
wJXeu5Mse/tx57wOpyjmt6nmVOhhCXrIO+NDy7NsZnifJN7I8iv2B+3XMgbdDqfJ
djj8nvZ/RYsOrRr8FnXq3OGCCM40H2xahOG0mkFQcQnq+cAJYyX0IUbLt7LTT0Qj
sDUJlwQH5Y9zRvmeGnYE/2kb/jJ4TaiW14z0CtWbA1ujVoYph3BASRelj9lYG4yM
ERsz6y/csAsZ4rSRt4jPbVJwFNMJlukFRe35RZX6FJgDoDMTLhYT0I3ziIpdLT8y
rsHD1UADtRrLNnsnK0MMYUUEV3LlOD1GAbvZ9lFebBSp5OMQuf9g2VWGra4fW3Y1
DjvFaPKcW6o8GblaI++yPLNVUFf9DJh/8/lVzEPJhuItqqrdxyMdGWe1TxDc6q3W
jmnYraOjyPXJO5hVZ2k1YQ5dA/e0siRO5y/9s1TEzjEzt/BZvv5fqduiNpXkET1f
1VempaSCYSc9p71gSiqix/D+2tb6x8ApWvaKGcTsLRs/edw9pXgVccr3tWCKv7Ml
Xqc5U6jSgW7MhfaBygqU/6xbmynMWn4koM6cZ3oAWSN1toPnWSmWwgDCKcm75w26
UCdavJiNQh/94YqaHD9cHpzWmdNC1TCUiD6QnfXM0iqCUHcukcx3dRw0UwtjNB6U
86AaF3oiBtlWEcZKZSoguk2KffLICAC5Kxg2mXiD5jcCB0lohEL0dbLLsdU153ct
gbMNHY5UkCwHsiQjEvNL/ReWl+5ev3BndfoC9tK5sLnU8GsMCfeUZzHbMj0VO27B
DmFv4srinQaW8b1jlmO101vba+hM8U8ucYExwbIUN07tg4Iv6HtP9dMkUaQja91F
EKFEMPwA4jAP5qPh8wTNPbt37+wzStiaM/QQeO90MjwJFS9eQ7S1/nOJilPxcMLK
qYoDWWNZC4inlHkCpAg+mMe567nrqOwusw9g1+zkeGI3KA07pIobtWd4x+PtWHs2
2Ta2H3QpeoKsmcHEDHrA369N2vSmT9cyCWZBh5KfBMEq0hG6Wl32PCojMPsVuufn
YbzJckmywGB8vHgoMuLe6IyClMv47UQWF+m11EYN4i0Hj31D9YZFQXjUp8YDi8qR
P2BBaz0SVTEDI0C68qKDOPVryo1HsoH8KsDaDKdpW5HXahO6mSRaTUqmKNDJ1naZ
zoikyWWeI3xYBnylqrvB7d8D0hV7Ne3hmBlbPl1uXbiWkwrKN+fQl6fV+DYPC7Mp
uKLKxrF6FTk/Z0A/9x/6Cs3cKL8H1loyZtEt9zoWtQJM0hkfA2SCfB8FdTdy8HRn
F/369Er7+txzpJLJ9EkMdsJINPxpKj+2TSpilJzy5RcB29hM85sVbFaDOTj74a2x
xZoYTLDN7BEoP+FD6gq33bdso3LAjW1HRgfHwKTAm8NnzxFliyuLFtKtwjAAZl08
saoie/rO0spjqXtAVyNvYs7PamsxbJoetmTcWVhZJNYjKTEwX+QWU5++wSMwvNxs
HXlyyjZ7ihjuUzQmRYuki3yL6NIG+DsnupWK4WBe2GesFSVxd0BVSjX1KZ3ps/I1
WhtxFtQnuUQPaJ1usIWyRJwynLo/sMkgmJkT3HiNpKc7YiL4HbGzCunkioU5rNWn
D4UzD56+b73qpk7RzI4J5HkBh/WL8lakO46KAThNBJet2SaUFIoEfq2zP2Tyqm6C
AiC9ztgUs4GPFTKWdWj1ABFNUSRBbsVR4Ih+itjr2RRMVfOVtu+exMfQOs//LJfv
gv2JPLvbizNnnIWqBSWmtWy7gm5JTLVpYgGtDoiTbFykyFyDtdtgjJx/GbHd/VDv
4AYedNjUWWcUgyJg5jnhgF9DA5hku190RMv0jErlHz/y1TYEQfrXoCHtXScwmU2+
XbNANZAbG8QPGfbv4j045+sd5ZjxUhR/1h6dJdOgy4m499zLipDE/818LAg1GZtl
NZ3TJb5z+0N9PJkbRUqlKEhzA9VFlxRPxuV+dncOiz0Qt94L/6rsXgciwHyzpx0G
MqHi630LwBK2zAyPHPpaVc74vJiK+FeyNtqFNYliWENnmnMkHRRm5oYmdH4TO1Ig
19lmDTdB4ZNhTbZuJjTXyA8W6A560st7Kfcot/bL9LwOCLbGxastZ4oQ/ortauDu
U+r88l7u18u/CWibDbKQQYDJ9BzhgncoluUumcZSTBPqKoJg+5JSqCmqDMkFUBOz
uyDDOtQQbRW5gMpvlvZWb3QX3XJ3KnJCMBgRtbQ0jYCtUmBNtJNHNntDkL5UTNQw
+QJsWu9pffj8TIOcn33QWrZpuLWTJk61i9BWu1nzAM5DtDaM5Hc2s9LYbQC/7EXA
DpKf/qQvZPZ14RhL+PcbaB/THRlP7r+oZ5V42PIbN53PYqm02Lai8WbMo11dOSxA
wLTorltLF4s44u0ih9sQbevr5PTcQOvEu/i4kSUVQnDfo5YVW1Q9kVbjqNQYLLqt
4RDnfenyHXRNqFXfKdRTwgfbwabpmQdx6A3tNHEkzK6p56vHqDPGuqOSvjka2cZz
twG5Y31UTwNBH+rAX2vDUTWWXNcZGkgcXcK/31g+7HCfEfTAn03O8xLqdWVN8BgD
WevV1RB6I83hs+25QCP+sdmz0R0s3vPacONd4aaw1yl6hRnJ4mzEPHfit5ndS2eG
OJuBdSXXmYjlCn+NdgnrEPdHDjPLoThmEbtbsMby4BvKcpOiK/oiLnroPTfH1QXE
EXsGjAllHA4y58NRjSq+0qqNgLb+7QtNPWVkNLQtr4IqwR0LAduBKnnGbR7Yigot
eCUwMJjiHi5llR0rdzJRfBDPG16ygPCnl/c8eWAYKY3HBALCPZrMFT2/g3HKI+T8
P8mDfCMtncTBoDVpBH8cLO+DXfvq8PMNc8x+OYSj46TH3/Er+ygoW8WYq9QBY3mE
KHFGREPqxVOWRuAP00J8UarjOYFC6AXES8SpAAUJ839BqqudTloAylhnUFgmERj/
C19G1qT2WC9KNtVJsXl+MCpUScGC9v7VyHEswWPchUWoEBQPMMEyCOXuML1BtGDe
QIHK+shB4BOvKWw3eY1l0tPPfVudWAOGh74FLG0+eCRn9QPm8odqX7L69/XJeTwb
5pEZjDdtB22yXFu/EpyPMHhDYne5S8R/JbmLhfQc9CKHMGVaSQaMmislT1/KDuI0
f8P65uhpt/+HSBlIlo1w9BPg/yVEWmiyVoN39CIH8rz4WBSZoNUP3fZblNNa8ieP
zzlHNVBMl+yohq05rniHG68eYHiQkW6g0BX4iGxAoa5GsqkVqYyKqp9c5n8TPyZy
pStyb+fYOnXF0nM/BZnuNKcOdjN+YdKdR0Olsv0x20I/MH62azfbANyB1AX06Q8B
9vlAm81UdXBsasgUPNIxY1GB3kveIFKXEh7ICDNSvZ2mm32/m9AyUHw/OeVovIqO
j7bdgFpuNhCvJBhx7hrxo5ojgo1LqvVk9v/qBLgPxBPyHRNtoNZxI+miAeaYBuqG
wp3RY5HXUQbPaDQYjhwxNbwCce0z/DlVUuJ9L70CT7ACeBzra7Q5qDV1EXICi0eR
7vtBLJ3Tg6317MaGD5AD+vIb0ZjeO7tFJnuSBYrNVI8/oO9M71QdsIjXBBOCZcgD
JJK6NNURrdPq0UUVYfj14JGVyPl0P52d4ZdJhH540QcejfZ7UBn22Uw71BG3Ze7q
mlgv/0WMTdGqqknIPR/uS0gKFteETZBxmaYaK/rlp/XuZlulr5fXbHha311epFq/
NZWtB1OyS7cGmQ5bNIPB3nboqAig1SUKIfJuia3YxGAMgne1PKr1wb7uKJ3Vy+U+
2qysWXctl9d6WWX0JBCm9+T7USzuhPZkqi9RUpAsn/+Zs8bOinQUNIZpRezOeFbC
JT014QPzEnAdCXja4dr8ISh1s7Wwhg1zGELQe40FfgcV/pdgR+XsPO1zC4X884sv
USjRJGvsVlQFIQY5nrmA16dZa2FrzVay8cMcMcH7CRWIj9wlNBIdcfCutDH9wN9d
5ZWD5ybFKac9EL6NlSxTdr6amfxVLBCdfZ/zYiqPZaAvdIMvdhuNjLJJHllrga7g
PqzJmVEW5x+fbLKIR8J22SrERfVy2MVSKFDoHBjpfGrloQwAWZI+S40aX5UvqsW2
vYpK8NNNo3ky+Z4mroUZF72PmzzVryM8dI/JjzzUenZrhJAPPNPRM5V8KPBuhcZv
AYF1LJ2m7tNbKEbPWtZOImekXay7qifjSls2ZF+qPIHkSNOUNHKswCsHNeykrj1e
EyJQHvVmJviPJg01Z2crHBKtOLVACGlz4r2fJWFCpkRRjyqk5uAbhK0hSoIz4rxs
7O/xGerydytPQleA1znNzOswOXxTPEvNpSs50ECTKWOoUUaTG5DyTLO54f6cAltC
DJK0LvLHj0a2WJ0qsjORdnkUgKDAPI3jmgubzeeI0oL542/gq6quRgMNyzWMasaq
WbZmRjcHSAdoprH/d6a51UsC/4VQNm+FRNUFN1QuokeleMrZ/cJCjUKw0pN/CVZl
g6K15zNf3ToPaAXRQVZOcB+Q/qAAJ/LBblz9plHAmQFrGYIoCZk4Og07S4F0ocmm
xePxtyIV58jiDMbav+LCW8fJ2GRFpFyGrQQGRRRJw58K3dRnyKXW3v9k37WwealQ
NZmZvyaHOZov2HdYubI9ertYH9Ml4YmglEVssBKTfCZLNmgB0ehnd3950jqKHAWt
qADv6QiaRkHaxE54zlGn2mYJp0tkbMu7TlFJQ9/V8TL/3llzxf8VT+8K71cMicac
6H56y1yG6MRKpmo5+keeXmuqqzzdHAJQ1/BK3ystKyvK64flHXg3Sd8GNmBkJRqc
egxm+FeMXaSL3RZNJWpW3HkYXO2g/edyePYqpwhsqEZMMgnRlADnH4Bi4uTmJLy1
TH9pfPKmqXx0FPmxKCLdR9S6eSs4VK5GoOTpGcRmQ7XQK9ugoZ1HvqGXTylR4XVt
koLVg7WADGVjVXTERKe2hli3tEtDU54gCIMmXX5OVWsU2jLfUevDDannp3RCFFKE
tAIyrAfqEgkHFWWnLEI5wE6V+516o5z/Dtk/LtQn9WrWEGNXiQZWXF2njLus+4Wv
MYP9WH6D2DvqSJMbm0gljZEo6G7s6yyrQvpBcZ9OJUZB7oyQAyQjVXwgfcj2xVn+
+l6E9fp9qztL/eE2TyF6MInYH9GH5y5+98Xaz2NRyaJ2CTKZKByCjJKvKq7CEREM
tZwgUjbYQS6XI7B5R7BjtClt7njhaUSIDS3xc2bXznOdmOcrlQIAJKdvLXvAxcFu
sH7gx8nyH1Q6+v7EG9VrhouNzZlCMndU6r1et281ogcOD/ZpuXJZ2m8KxS41hQXP
/WL2z8juTn9chUvH349UKw3AIzlOA0WrqzDfnsCdnvKOc3K0CUOOnLPfwtWdxkXA
+jL/Mu6dvUhO2e06W9mtGayE0grLUZI+ghU4A+3H9goeNDZ3WkelJPydLxr/f/Hv
/mv8rzWV2H9jvwNPWvmhK6+muXuRtloIjtH0wd1vELhM2RmcPjCVPL+Q06oiI99f
hnS8j76AW0TzegzNduGo2O+RtC4AAfE8Ugy9vvJrFWldaDVMaXgPg8d9IZrjGV8a
aUTpfKof0pXUVseAhUR8LLqm0cNVZo4oHF774gj7bmAcimALxrf5wG9gG1GMkKL8
Vgzvz/DiMWCp48kMIrTw3ql110s4MVKAt4nQUMsWOeV1uAirici+DtOe+HXI4U4c
tsSfcmP6zqPtGvnSCPPBYeR+j3A4760M/3OAKa7IH/1h4epREEo6D2vpqVwZKwJJ
gB8uqlaHdY8U99zoux7oOGi+u4nKGsLq6ijg51GPPZ57LdDW99s2GgX495N587bf
xkrVQTUJL4oVK3bFxdcxrw1WlCBdLxlwPPre4r2CUN+EtCm6zMebSqTMp5JgPbsH
y7OIZCyf4K6uilP15KOZ6jO7ftSmi0adAbXZWGl+iF0dDKh6VJg0xmdXpsthxh1S
t0Td/89Uv/mFQK1IKWl4UK6D9vqDPD0PVQ556XwKFbtfsDoXnlSdOs6Q52/XDEHx
ju6sYy38GmWwWTH+Kylcca512apU9YaqZztkC0tOGvDYzuSgGiocXdKt6QD8YzkB
ZYMbT103RuG79HngmjbLI0U5RCbJmh/CuqRnAzOAdwPYtMkiUEWH24DreCwdKsVb
BOrmKmGUeFy6n4cisMJn4kUaQSO3xeEkYlL+EzmPQ1HSAAR9AOg3w7MBu8Vcgvzi
Quj9k+PRMduQpFiYYCJOLTIJeXeixaT19DH2KKNxJ1IjeW6lS4NChiGdrVFaOukW
OU/iBYf257Mf+yDTbvAi5PWAnF4b0+c83xZ+dn4Vx22a4uTPX32Vy/ijLthqbkO1
2sx8CtQPMEKAwQ7LYD/Hjnw84O1elbQOJxMMEkwnAHydvAiagVW5VivAgaWn2QWp
WZTYtWlBvXr+UWldzuGOHfnOMHYWd9sKPP7M5q0ODzfUydW1M2xA1/I2fwQOwLc1
RGy6V87b6Uhc0uhJLp91crY9g3o9y16Ydib3l81yZ0BaSfKW30qWy1hD2WHijjYe
7KCTJ2JDUWialEV65741sBhnxJ1NegiOQHF3XZfGhMg9fopWC2+47G2xX+Jkr7pk
O+PI04k/fAasETAYMK/6aOAQTlB2jeili14CD9Id9s5IKzHn5Z/c4rneKnLjoBzi
AOyZwniXDcqD87MRsJvbCCPc+c3bzyqFHBjSbhOIzNWm+vIMKOi5NTHegLvizWBS
e7W8UbjqiEUDSkV3/pCEzVYxQKDmtZ2g7TChJTqi/n30IhRs0nqjGKv/Nsxf5vzc
4cwA+SLvgn9taPgTUAlQ9BM9A0Zu/u448ax5lsp9j/Vq7Es4eNhO2SIM15ubwh7N
o8W13OboatiEsfixPKHq/r1W/Nsvi362AhhgSudAU2sbkn/L4wmvaCqJbuj3OBOK
NXc4H4u2G0t91aCnEhJ2qIC7ZcK2kgXRWNsufcBeb7vXlj8OfXNrTpG10QZJyozw
1QjTjdbZGUuSpqc6jED33tQkzmVzS3kaAu7ZugHXKWeHMY9fpBmtFFzzqC2U3A22
Ey+uF9RgdZyqa4mijgAxppJKVeiT/DjwEinRWDsoi2vuFSvIDQfq3cr4PhrXCbHl
QIvXWh0YPJynkOzMgS5v1u83q15WXizLdgZoMsfibG81l+FWo9qFipM/1HkFFmM4
c3cmyVaY3/EHjpCa0JowZmDdGSSN7rAcpfESukZi/JigDMeTBjOxj0FGVu+kvFXY
s6FSRpokwZHchS1vv+Xp76j8L/D4z1tTxp8pvCI9KmGLYa98e7xMyB8LVTscDwi6
2SAP7SSxaiD0uPBRpaXMD15mmUANOrwYO2oB8CPLGfKxlnmBU1X3OSKtRcZ1Q+zF
Ay0b7kjeFf6wfqOO1SNEC95iBu6WfvBTMDafhLwnFCWjJVchRhsfov7yMWeOTF8+
ql1w5l9neFhT7sL2/QaeXBuNf89osMoiUrAEDVMJHE55XaVk5Kx4QHBMIB+90bqK
LvbOUmNUL0kW0hAsEZz7cX41sUV5deiRfuQTWCoxUwPExzGiouWEGzq7uZt+fLPl
1saORjIb2pajs2YeuOAtwHbOLg+88+geU8VxocizogowDWCmlDYQ7NMDkgEdX5BC
nB2Dd1SA+rDhELUXagLe3JPwGuRaxeX5YXb1mKPuOt5vA2+RtghYRvqG1D/EtlZc
5jOSXoQP6yMDWxU6qHZBdMr+1aSi/SubRNt4xjygCeARJplYdJ3JI7jJaul3r8cJ
JIfbS/RXxWN1LC6boyq5A1EZtSjPZOkdkLL8HYMhVRwCcAKqgcHjQ384zmYQvN/G
fc+yJfUgbhfnv2uCJbgf+LM+QeQOnFwTUzcYt38MabbhVNcKnvpewel8nbS5TFM2
AsMIE52sBIwBhdxPVDPGgs7VslWwkMqjUEmkj4xScbsbFi/hUDN5p6w4fMa05onB
0FsA0BOhKmjx6gv81w4YjfD6jwMnTnfgZFe880w6eVXCIFdo6WQNfa7MlCGJo5YD
ez4YKsDtZdFwkYOuqjyU5WPdvQdtnb2Lwlc7eCHAKP46U6nigKr78o18sgir3cGE
VfzE+A/jtcGjibwcYdWQE1pDfSdlSjdY8MgekE1C86qq2z+Ys3n0/koIMlMxtBs7
AAT06OzXAoggLIo+KC/+Fwco1Q1E2WKAst7KDDxHel3pUKzUUgvZnYR66RPyuT0T
Br6oQ99BLpgf72tvMCTqNPPocxVA1MrWIei7Rn7/NLKOySMhdG/uv/43O4OXFTRa
fuIgmhnTvxnmd7tJ3oLbcB5zAEyZDLNnk4iR7xn3kznHJcpzqDB6LMyduoBjbckL
WW59p0SJEpIfjnwY5dtAkh5Gcyyt5jVpqPaICAiOlvnHajbHpJREudA6JEubxFpB
qtV+jjKSVvToJuYagmWo6tukn+Ro2qpy5R+37RGCttg4333qZZ9vfWTX9miPuh60
NJ3WN+h+AykGaIYb/k1ddwZeMlVMTeYIaBjaUnRIVdmcccXqvlOY6+avh2XgjVTT
+eGS08uQX+k6fs2opT4BmZISpZ5dfM8cwEm8RW0t1IAIhSHoWpBfB8dJaNEcrzDG
JYWvSMquZjGEV/t4GUJ+xABCIGLEolXbuQ8LV7N9GhtSJxAArcOz621WaTjf+Myw
vjQS488KuABA8LGFQIeVT2KVWhmUBHn5iYn1FvZGGfastzXZ8uxbusmcp4zZHPNY
tTgpwzRfAHtHSj90ZT8dob6qSreS8vc1QHwcFp3yYW7YdSNRlABTq6OpmQQvyAjd
4Mv42ht1CRWZindMc79ooQpyvWBchLdJ4AmknFe8Mulv46Uno8Vcg22TgLQ9RY9x
EJkqqKFCT8U+AlsMwwwGrmHxmDsykxyKdES7TuRtPe9X++i1yRl9VhpUi+SMAYV4
1Ak7MLU/ozMTtyBdeqOKq96CESisuDERzRonU9pauXq7A2xrS94XezZf1k9oOMBZ
vWaV8UfJ8QpLsozlpTzEBCm7uoSz0G2SPS9WRHOSYPndnzSqllckzuO11UBPJApw
ek5BwNt4xh3ichjk9uAmhPLUj33nqDd1ZGfsjka5Fe1wB0BB+W7IhRGcmrdZIpDy
O5JU4PDkyBPoGvqDBbiVcHy1mTL4UH2+QKYMCwjBBcimv8P2ixVeqSZH+OofMakj
yaMHOI/HoYYz4opzkt+CRDyNxy+sT7q9thLseSNQDJwk0PKi+OCznGBnsswy3J8x
cH+kn4IiDUU9hCCNC5bK3k1/Fl9wBkOvhsj64WzuUbt5lAGFhFy5fgl52C+ua2Sq
3IELNJ64y+bItaw7bH71XFX88puCCUyoVADzwYyT+AjOnkxTdwQI7EI2tqlmBcjM
kMRPfxtonAzf/v0An2IV5PnjPjj09n3xYAlX807WdqzWbswScPYtCj3yjGlkYOM1
qk8Tt4/IVS5cEKL4LI5bWUYOvNCy9DXjxwdonOiYYF6xNu9d1l6w0ObOlXOD/oth
AoxfGxmXTuYZPVePa1ymJYGnP5jeesUQy9TBBLnmgNOl6/xsM2aQl8N4WWr1pCWt
yrm9THK59XiEml6lF05chXuhDJeST0Woba8rg50ukeL8u3qxL0ITJRBh9qMtEddW
am+rHaH7KVaYJAhVJU7KDUGHQsVrrrDHKnewIYH2tgugxyDeLfmPhGJTT8JdXvYo
LbxhUKMdelSrqMjsX3duk+7wupCgtsvaLqqv7jo3DqnHmOOzS6Y+QWl+MrItXk0a
f9KGawKeLjdDj0acx7kt3LB2eZtJIX0PAl91ROVcns+gqORYsBPJY/EzxFln7Nzj
nyEqpqIz7ne5ivNvida8jBgsB83F5J7lv/djBHuTVr1D7sBq15kR955xi68s+w/B
b74bR6FN7Rxszc7fKtqx3KjlXd2nH16v1tm6PiBPFVxyUa9fGgRWoEonDtErkiia
8bOskI9kTaX23MT0kDFBpsGPXNpfSbLda5ZhaIaZMO7a+4xsC50H1dAFh0PFaIYi
JB30YIwykbEHqZV2oUZ94zdWYTU4cJesDUP8YRqk4ZpZmzDmtAXZtfv/qB5J9jsg
rIlcapIPqaKHPVlS/IaRQJZ1nsH5myaxPoqEZW0CSC3wkJKg3UWBnU42JrC+XuX8
7/SIB4c7L6Br9LVtehRE269efENRgg1US4wxbGCXBITrnzKuqCt4lU/Bav4FXnmO
gqtNkwpx5jhS5hCow+6Z9VjJXGvA/k7Xc/XY2RBmSvYstLTPWc/FFr8BTqmEtnMo
6lRDUY1FjVyTsvEWub/cXO1S47vIByl7wcW8ly7UZPGUA93ANS8qUK5S5TSgxDh9
B3VDd33bFJt4SSzWGkqWFdDgSOy4r212EXNBi737aFhkVPQd+bQhoFU6oGQ5+oCn
I/wK29CA0RV6L1KkuFhbg3KriWHSERA4OytXQVGliwlG71fSyJXVWcpNt9wbEMlT
gPp71PbQ01+0GVnnPWNay7CshuHF6Mif1cABwuLmta+iPdQaNyEhkDdQsVmWSRLk
AJc2KEboqE3bFbsxcKda9rZzBdBEo93tbHlMHElnFvdifAqZVgsxwGKkRdzl4s8o
jAhb2x9jeDxFEH1LX+aLnXgPJ7b4/MCYJhWfi5yNFLt2SGFo7xUGj6ZYkc9uaQBF
n825XGJ2vAm2Q1MJrUotHaZ8scf4/wYCrFUF5KvJ13O5iubVKeuPJgGeoABGsMQ3
tzBbE9r5zUoyenTlqlNzAzRGP7CMXF4SHL+3Cc2Zu6sEDMJQFDtryQFhGBpdsjL4
UqVborgcwGdV0bXz5gFPzARBRu49vi4geI03ferrv4xHDJ79njwriZhJM7lWvQUY
l+8F0nxD6q4nmG/sbeNuZsbQRyw6I1VskijYLfuEVLolT8H5kyqU0r+lVP86p0uN
WHlN5g15OzgBmDu+Befu76nqpREawafi5agRdvB2RtFmx/9ug3i5xsPIk8LB3p8a
FAOYt1vvZTypsO/3egw82UxrKU5LcKSG104V60yP57OzxzJijcRdGEB1ddnznSLW
shWk4JwLEv7eSoz/hgxE4Tmj55MbsO3bxYDga3v5K6JozAFy0We3ZY6ocZM9iw7U
2e4ZtQ/1gtHa9qzL4MuUWNIBLp09SKxDK3o3wyL2bpgydT8d3XwslbvardBstmVY
Qbb6yDfQqlON1VGNMz37BWwrf4OUCzPvKw8zmwUvI08ZbDPm68dR+gRopK93iAiY
CL+4C9qggHGSZgUH0J2LejRqcoOzb3QkbCPXEfrlS1ifL4xIKuNslD9C91WwG/7C
6WZRBW8d5CdP8dtTmIn7eB4ikez4o4F6RqkXp/+B/VJVWs7Ud6BFwM9Gq0RNdmMW
g3L/4Oxx+EYK+asRg+xubye4BDThmoTOLZRMc5UBMHUTKcIoiybqqse60FKy4KOa
aSmZnhHb+OPJ456kF5ZjSqhU0JtNM4gR9CK3d7i88OcnsVc9szi4Bfty0FOjcIGU
dRgQh470vYIqH1SrtQwmQ1hVrekkEVp4gj5vVgMD2EddnKjgD6Yny0jBaZW3CTqt
MaEDzjClbaS7mDCtp9Xj3Uyfu48TE6T67y5gmCQ9Q4517D2mi9z6Tm3/NMx90jBt
60R0IevRpxGRWtzxddmp5I0N8fs/lwA8D6YLS4wrizeWxjKhBbmUeKgLPdjn2MYW
LU75a31vgJyx80utJtPy2Nt/qhyz1F+CAt6+/rF0CqqE1AWkUee+Ucg4q9y3z9+k
ce9fe/1aiYhQZQThcXuDXKk8EI5fWHtkaZv+lCI5Q01C6O4DZEoWRnkHfw6j/Bs3
YAttIlH4l/ktnvbb+F3eIl6/H6w2T47R9YdBecLR23VBu+0LSvTYyFQ2SDSCpf3x
b1rBeeSfrl9ZoqbfaNGp1tyqrpIKABv0mdINrVy7+Aw9dRqypdpc+lGWYSfJd6T0
JaoHEwjn+AHSz98rLvdQlP33PTOqmY5Czp2jA8DRKGaqDxA9ZMMi6C+/9exK9V+C
bSWhzyaVLOuLUd+C/L97ANN8eJP6lp8X+dU+ACyj7z0eIFu71dHUGMknSSRT1kyW
mQ69FpoyWKfu8H5kKdAqdEpeY8K7yMAhGKEggNdacj1b41ryMkPJRg/RIzOnDBpw
RKoLP+XCXpicF1r4t7cYWH73x42Td5Mt6VQ+kqopldXNI9kTsB6t8LW2JovoJNce
DDpy3rcRx7/3aid/TLlr1Tcx2HPj0bQOb7nPTNKpbUiSqDIwv4sONBPFAA2agI2A
ygUFZTYHH7D5ZtSiVV/HCkBHBVFBuNfyhsC7mtVs4Kuk2zx5sY+Tm7UO65pT0B3H
b1MrorevpR+37pHOCcdf3iFWl/7QFGPgBzbtgXj6V3HRYhSbwCoQYiKZ/Ekd6wre
jvxV+Fy9rZJS99+onWrHvZH1fuRJYSUD2UpA5YgLr7SAiO8LnFL7JZ7DcbGJnyI0
TqHBj3xjmdXV30C4oWzl2q1rcSJyJVaC7Xh2iHZLt3Km3dMbwqv+nNkyGE+KIp5C
PM+cnY6NvEr2ss0zUyVhnxh6S/ZrmhlY2ZP+8pAFEIN3r1sfZLnT3Dss9Gx/m9xf
2TaF18m1pt7wK9gqAtpqELeZVrBvg+qG/KcOycaNwIMhbP3xkR6cjCnqx4JuaJyV
d3yyVjO5uoASQEOSghc9ApPDIO8Ype2biB33E2kftxYKZYMQv+KyBvZMYSLWwkZC
CjnqP0Q2FPtoJjMIYPR8TQQiiDq11Y2ZLYdLmMD100NiLBVxu3FHrMwk9IbGrBD+
SkDOdRtwfNvpBXTJE/NZeRrZXpXXyI0m9c/SzXrmpT1gcU6lPGZMp667kynXffQ7
40RziK0xM2c7Dn8tkeHh1on4P9F7mmX2nvT+L59NS+kul/m/S3GQNb72HxBg8qFV
B30FUQp1DOB413XwcCrEFwPdP7vma+2ZCSZmUNJ7Vc2IxxFwQWc3rD7nwGuBfc2C
f3qHDuPwEGMCRZDqWrOKsU9J7gvxLfcumAZot8sWG7JY/21Cyq9px5tf7SeKXrx4
OCBvwU9DYu4jeWHcl4EFZbDF520R1tQKgawiSJyNGPKZ6qRAWDXEPgqCc6cJko+0
zM8nHdT9pvWGtdVzOqQfk5c1mqBBBoq2c6qIzxg8D+AGFXyCMquYPzF8dP9KohCu
BHvX6fYvGtaCOCD58CsGpvvCROspIKxohNUSmP1lbNfKfxmEsXQlqVbD62f9dZBW
WDU2elBMVPWBcBtY2hS3VE0uNo5lxxp73R188bY+1IGoZApAeFJCSzjgs6SQue1c
Oi2SJ/+xaOP2vtsZTSCvRFY9U7lOV1mwHAUnQR0topgJUPGC+a6bTIKSlW+UvwnG
fdNYUqrugN8pdV6DLcKvaXe4AMPLei5It8I5z0oeypgUvynf2QcPLty5YbGaMVYQ
95G+Sw1IC4lTBjgYMsbEr93CO9IgZ7mNXPVAset3BtrSzpERmmI0ddGyFabhjab/
Ml/RBeb61HNqP/Ry2yc7ERU1aHV8ZVjHOQixDr2tijId8lyLl5A7OTCchnt0YZwM
htkyZV9ifraKs9i2x6RhMucPaF5ZpywrdfTW+HXjWj1GOFW8ZkZ/uyGVLQlthTf5
pizK3sepChc8m7rn4i3lKmemD8AMG/BSAVNBIZD8menJGcGI/a9zr7JRrBPp3069
lQ2R79Kt45S1uP+6P3Y1lpAXAaTdDPBO25htf/Thz53ZZ7NUIa2sHrmv0VNfG8Ux
jofQePo0LuA3+y+pYC536+GHb/zTbUvcUFr3XlzTvcoEnhz6Cwefbcsl/BCyAflz
uN1qknvPw/e2g0BWASjhepRUxRyHdqBX7EmZ2mfNzG9VKvCgEk7NfzSq0cly+cMJ
LjIhpzDY0W5OedOffFVDA9JXxUOed/z+DuftoQmc5Cxb5rmrQAeFzX5eA66MAXo3
xoy1/thUT81Nk/MdLkdj15xVTTAsJgiffwVcSce9kZh2CVOHdldGVybfh/GL9ffO
eWzmIZwX6DB4SC/bBktH6f0hKxtnc2glXl6Kn7oN5ouAz0X941j+n0DR53UGTowl
AUG09SYyFiYecLORisDWdVklYhYCiAaO5mOEz8JPc/LAd+GMACCv9N8hjFNXWIzh
d9D4Cj4XJ7dEaEyljA2pITnqWERDEU+NnyD0jBrpcgGJOb9hhbnpTY+CxvkmJEgc
A+zd1gAXzm0CVnp8rztVC55En6YIsgfA75dohSu+DBCTJdsHWzVtizaZLap6sYFA
2kBrbiyfKz29u/4ohwbjPsfwAhaVjuXu7WiFwTUXQ/RnAeojzko7A3hL23/lTd1m
vLi3+AuIu94bVCB6p4F4u9vhamyS8rod/mSY8PYQg/OycKUhCIBxSSBP7ptv4AHI
TkG3D8rats9HqEBaMCYm+41SyNpSFKD8JFkQYWkQuxLzxMm3sdm0o4VKnBTS9I0x
Mapph4RcMt5bzwiifXn0vCt68No3y7uwn0xdeE/AC+eOab3br6J1O9ARGu395bn9
5e80O6mYBN9TuS9e9ikzvjE0GMv7Kcu/LpqLAjSAS9l3x45HJ6caTTHPIucXMeUx
jBfQCwUcmieuXGvugOBBJsB4wH3Ar+DavWw189N70WWYwTaJrY1nN451Uo4cZMEF
Uf1Qeibk7Id4itOC3RGfu7s1ckYv8OSZZ87Qppv4mGnMuNXuKS4YwSd71+RpcDNu
AjZteBmaILEqzYqy7cOEJ9Ro+ZwUy4D3Hj+HtapjrkWYa637ZYl0kIsmUCkTKfXS
N9le/v30/0AldyAxCYJKlcj1MzZn+WsJ46KIdKfgtJDiqvzs/RHUQ3+Q95zKGtpv
3Z9oXJ4fm7uw0YiLkGeOTXuBki+fKhMowKDjR+Hy8wC4xydX+OorQ++gKTVVYoSo
IYJdAFukoNwUtRsW3SAC6UgqsEaL1zNnYcmk7W5nBGf8zAcWcMs06p0nJRPQyNca
haPRQtS01aw0bYCNaNW7RK3bjubYXvsnbGKU3n0kW7cNjabgKEqm/P6SdlBSIALE
h1fdPGR0LQcNwNoTlfvZyphFvVbDhEmUXCfBDDNXG/5oivHJpHEx9QSvJ3GSFuHK
IKcinzyeqqETcs3YAV3Wn3CNnJgvM3zJgIplW5kS17wgPUnTMM23jhBGJ0rGo49X
e7c7I/g0vLkb43bucqtwbd0fsuyml7dXQ36nHoEhwXa9S+Nx5zLilL9JnBYVGrZY
OS+4/8GdokCqlEbvj+WZsb2TPQ29gIDImxVd3zL6BUvRfRxuvYYCYlliBQthgOfx
XgBezVI2vUsJP1xgFzM/TRgRzYqFQDPzP02aod9PoVyqh5JZbQovXTOVhIQy1Wkj
ggswcym27nulHcJGAd75JMAbx1fy3rF72/x3+4LR6NtQBX/qhhqmJiEPpLk+LsKR
J1o0VyrgyipQFDpNgIgUQrqbFFqowL85NvufQ2RAOgux92NXiLVXuDcTukbUTe1A
xBGsTFTTSpybeH1Imvwi8DSbiVgLWnEXQ6kPVvlj+ANkq7U/46p5QJtdoYKqS5I6
2BYFWIEcpyVbkR5la+zs0Hgp+ZpF4Wkk0JTSPZ626sImQcJ2OzuxfqalrlHdILXg
mBcAUwfML/7ebJnuzjAboxm4fRl3o8qsw7nd50aGs1XOHy3nhSf5CwsgoQr4xFEC
aXb23uj0qRj4+3IB8VwgN1Semw2tBQGefRqr/rYT+NF0bX6Ip97UTqAhQBoIGNeh
zVGcJMHS4AjnAOVDfJIKPOvlpDf9yqsTQTBgdlUFLpldeK8VEkLVughOtcaSdNjE
kwZy9sEpH0QW8kXNZ9N0u3beu8LZSqrsr69HAEXMv2JdNdDScx3C7lpzCJUNjE4O
7phPxzYe5U+MwzHUTGAcCiMsIXBmf2pHVT0J3km23DE0Bfm0F2hlgnT4AglSorjX
qOynlEcxr6IrZ5qiF38DKfKsXYizc4EKxdjGlDCiX2I/FsoKVDXPDKb0G2YdkTv9
uj4ZO7GqIIvu4nDXCz6knz3SQm/8M+vilfDvA1tYwZancUHqzZL4CM4lY/fYHiMc
7pqVwDz9MZfYN3pCcsgQK7AtNe0O3J+/ppIbvAMWHqD+zYStNWCXFpcSmaHwQ7hI
vVKnbMFFMtvonzv9+plZaf+lCFmJ/S479E72jUGSlHiaSxpWaPRtRWaBe5nyw6p7
nd5e7kcwjimIqvbvdSX22fvrHqE9+uuN9j2nX+PUNDorrPtlsfiiYSgBYGTzTsO9
AT/Xbw8dGiy5gHKn/DlCjZ32eira9op3KA/LjUsgNPoVVf7NTZ4iiRjKbxTgR+Bs
NL8EF+FeFXpOWEnD4lMAIdTwRqb0n2oBKAjqcFExJzJMleobWan1Ojrh2KmoZFbq
osuqSi+dAYsqE8D5VlMhoirI7nWk5QtCyK9ifN+v5ID7C0PbOiiNBX8UHuBAIa5R
IZwIYljtYY+a+n9UZHPbQQ64OePgtEkwhctS/YWr/gU4+WKODnHiVi3foNrS6ORY
yXXNRdUUVkw/pjaw+ZZRG9EibthykDrlXNC15owjxcnBontrx33nfysT6NNbjnIt
7uGtl/pF4FjWz156kzb5W1SipU67pycg+T0BEr5bMSRf6euNeY4H31WEf+Lb5/u5
6OnL7jLtAFAoNXKK4r+wjSDyCddkGgBEhTE5WM0Ri16ltx8tC71SnNroX05GKJTE
ttHixQiPOK/l88pKVnSubm94OBwckSbKQ3l4FETKvu+8x6Z2RODXRtku4m6hrdyl
/GMPte5OyuYObhsYJ3jM8qtqeDRaGDTlk/rc873D5RDxZGvK3153cOKP71744m98
E98aO+o1MmczbUc4RMwvJxNwzxMYt2iNwHufS8ldF9pENTzXVqGkRorse3vBU4Hg
SCOc0FhuK6uCBlp97IrFPS0JJT9EV7XGFA7EAdCbDMD7hxZJmrJEIdq72puwtvm/
CrfZiJpUuB5a6jLCwWR4w3PW5FG14yoko+WeYEUfDBqgoQAL2b0ClffLbwVUZtaV
jE2cyryPoN6PGJmi5tHg+LcA1+KNL3/bV9AgbteEYJg6w0i7Ksdq4XrWYANdUma+
4Bsm59qZYOVZBErP3G8Dfrt44L4XXhHH3nBQWdAf+TJyqZ2dMCBwfshf7LXsQcj/
8fVhTk0l3qvyLUq2giD4Wcs0L57nzb573+XprgTxRMhfJDsBcQTvnGSxdeuBe1Qz
R5mxMK1vhay/4HPT+2hfpXMhc57L/PALr3xCFOdkg83iRvtKYFlLMw3mgj4XWCys
jTxfqi69Af56f+9kfyse3IC3yymYb0aT7JXUvhTgnizGnCbDl8BTJsAuAl52D6id
cy7tUWyrOg608AxdgTmPtXTo2T3j40LULtxJRu/oVF9I3q8AdbGEvPXZlz4TzGoK
X5lujuGTda0rw8mUKa2U0zsKHmzq51b+jgeH8Kjyms3iZ+WF4de3SF2W5nIvcz7S
f6wVCfPZyu7WIappPP9rBrWd4b/i/UcnULqAdnqpq8p+ikvKD7N0y920/SiNw6rj
qGhd5j+Xh5eoQfu55iI9PBi6Zq++HykUuR59JDd38CKjVw45Z1GGJyW4MFOuytFD
/YG6jyNzBiKqPNiNehYZXGYTLRwHgOcaPFDOd+5A+dK9xhV1IHBsUiGT1KrgSk91
bAz2nEp7tHcpYakX2VHRmUZn9K5H4/yDY5vhm04pO7hgh905l4RAw0PkhsmcYLsq
pV73FkOYnW3nz2g4uE1pVgJnWe55yaFsdSxSnJLVVK9P5PtyManBn4SQG9EKG/sj
WrRzP2Woxv1qGyY6E3QBnV/nRr6NViZ+fQmUGicczY3fFTSt7TRrGxtzrVAs+/DQ
CCVM61Ej65qBYP9nx9mIv1NfynsWw/pIv5eHxEIQM9qm02g25dFxD6pNegD0fFEc
ibBLZcIKhvR96xY4IcgJzKBngEDksnFY4hknTIhlqg1ugyz6nrAk58urZAkuO1Pz
75OU9rHQ86f8gY/9v7gkPIGeqWYM8iuCOgrF6tJKyYcTjtHCI+JC9Fl68imO9viV
zqCGfPi6H7kzrcbPHSHhY74ij+zqblwpTaRgsIoTvx5xr23dw08uZYbmvAJg3R2d
IpqEy9qLg6UGJuNnYJEuMHjkY5njk3Kb941I6JXcpIof5ACBSIjMV/dc7i8CRgmV
DtrBLy+j50m5N7aQhV3NXUoU+4jDE95FxXBTuNM3i8ptlvsKQNnH19HrPkrCeU5+
RL8lrNfXf5UyiQQsVNdIayfSqiw5uNL/SRbiOPVfdkCiX1YTt0rJShKUfZ7evUK3
22oOKF9VrKT96t2R5WUXXtTEj+PirhO2qmu1CiLbLyO8bJSiquvixPdzrRT6VvvO
wWCb2JHv0tQ9HTDfj7RRnBRLCoZjq0Wi6EwSTqN3fsozRApRXDsPJbfTbL7lhzdw
uUOjxtfpANxxkVErcIUQBVSKMTAkyJdP/HM0GJR6gFHUjvW4gQWZoWVzcMBBMfSZ
K3npRlJqV8NHlY/3jP3H2gKFD0qyoDvgyfVPJraYXwt+BRP0N+5Bnj1bkbSu+Xhk
OIb+Rxr1pQMvFNQJ2aXR1XKmGvU9ik9T/sdMM4ilSg32V8Di7nRmU1+E8V6VTZlF
dehXKgpZeNrE6163aBJbmVzDOks5y9yRB3hy8cslVxJ9Tvy0dTnuHtHN7aSq3/tS
x8R3O85Su+zGvnqXzPb9MTP/YywZ8/L14tRKRk+sIjKPSC0QJdrxsU9BUw/8TSMd
+qnGJN3ezDHBUYTTyfjpftlJ+dA8m7TS08Jdlf6doAUXOzvzsa7IHORpnAeXRZM5
PDoPaoIHVcZm5B4KLWZn1vG6XnUGwk/Gv7g7m36HV8h1Q79TZAtzmAQZaQess0Rk
Sg0eS2mnQ6jkO308OqZjKMQYHQh3hfiZa7kw+CxCCfV2tRO0DMB/jxuREIAUEMm1
KIMOtzmLdPZ8542tMghun48k0Tc7K2WjhIBhPh/C7FyWXchjnF7bkb+My4WrEEYf
vkmECc6jvtzhOu+wUZkmHGvFtGetpBQiXtnxLmtYLAy+eSeCvLGYrUbItcHSfdmL
0Jxgth71jIo9j9oq1HU6QsAD5GZLvQI/NrrB9kCKvnl0hoo8XsEmB3ITuaQjWRVn
jxjvY04Azlwz5/QQtnhTW3dXO2or6dSRZMx1mHK1f1OWm6z+345blRJZxRBDjmF0
wxmYqXcJ2WhYez/S2kjV2WUtNgFmaLmkzhObUbgka+hf2qYxL9q67IIk7lJfrQ4n
6aRbSDWNjR/c1OzLasYXfdxcUmRnRXZcTWswIvyypKYXRqUY7v9Z2GYo91MgqaX1
hpx5MqE8D5nMLw3qfVRqCoCsN0/KoKm+3yGzPTbGMGoNcfb64ovqbzko27D4tUrp
8yP9nMGsbEeDg/FfTGIdEnm3d8DRHcCvA5cWFb7OYaHrlF9ssmpvNMpFcR8w/Q5Q
cwnrFsYplj5bR0Q9A6urMwHHC7NDyxu688ZF26nLRGugflPsVSb7E0CPDaGPM56r
Nc6RsNHu5Vf+9lCrC38KtvOm35fQJ/R4yAMDMqKdzEj8K/GSh63V07dXPlczLAl8
7bqBv3rgl0jZsDeu3b/ZMISBr5RRV0dG41d8nzaFTQ5k32ftARykmIzS4rRBBkW7
vc27u+yPP+xmzIXZalqa4tikrAa3Z8uPwvOD1Uw/16kwQVoM0k2VF1f5Ij8MtmY2
yuPDpl9m0qYx5/HGfrgDsKDZpgLQkkI+mei76IvmTsiN5MmXD8+KqtC2BZGHgDwk
zB0Ea2QH9B3Jn/tSNDS9w1mFcW/CGXEYEr8mZ46gHvdfGYzCia0AkGTt4Z+9JQ2S
M+3MdUZuIypu3eEMCmwMNhtcCb8vTPpYIUp8JjCPoJE0VQClRPw74oP/xszvAkXy
cxeZie90mDC8PFfswbbbxxQjqIqvEzQ9Cab4Ute3uabMQtPQG9GvurI61890fxqh
iifQSS2MQ8s6THxPA9q1TeTdWc0B3djJYzJVlOr7MBRTzMxCG7Xh7HQ9cp6aps1y
KFbwye6p34Ti8gVoejpN2fnHV7nhNWF7g807Gr9oUv2tLLeOyZIcwB1Hi4GVh1Q3
Eaorbg+X6P8qgIpNaniQFKLRh2/XBPurVc48biWdHaxosziHFpTvFOk0xkerziVD
6sZ7Mn4U7a51s+++jlu4cRxDuVzN3qevHOplNhch1uaJFXaxe/FFtnOJD9shtJFm
Ucv1tOfqVXUstIl+IAH5k2ugcGoUiAVuD5gDZXc5+6erbOpDXISSJdalRPJ73nN+
u+SBM+BJkWT7OZ18sGwpaKFdy4yJRnQ5X/ODX0WsL9zKt9iKHHeL8eK9X1Eticm0
Pb8pUIzjfxKTzbF4DdK21NGrR28akg24brmYMbjw7SP/vv9cPX6H0F4ABkVwB5Xb
H5timLIKJ2tuT/46ybHATG0pplLTx3nOS2sKaHYX396xOlcj0cJmlGopiHyQC29W
luRT9BWu8ZZjiQXoSgGAzrGxmaO87CDGL62Lq3CaGSE0PodbsDYATciXKCJxqgQr
LmM02WNI+gBlk/Tt4gvF/mLh2nOHEucksX0GS1HBSH2OpKfnNMcP9tIemfEaZEbQ
BCk+jgV6e3VCvZd5ahGNox8HedCqrhrEjxJjufrlXFr28RzkEiLAOi3ffWPuOl0N
u5Nuy/h/SFMI0xuYqvcsxURdUImWQIBKeydD0Zt7zNwLgLscfXTDTr80TrTAys3K
1UJuqNLQsPpUQyV/wkGXRhQk+sPOnuwI2gRiVNzTKDNbO03MsL0PbThHtieJP7+m
TpdbAw8WqJ4J7sQh/o0dE7NclKsmpz89goQBXqUzm1Y+cJCbgS6DqbgDX+PNj7Ds
iMAvLqkJEOinT5Nbz52KhIFe8TQjV496BmcN4kJgnrL/00qlzARsmsme6Whw2PSb
UIAGAiXvlLuNp1TQ+/gbiH/cnvQdbv4n8z1+lkRou8QN3ZHX6XG/R4jzzL04XylQ
n0K/aiE4rAuF6lTGiPYGLvFFOhIGp410AAB4LEdv7e5rAnQExfldDZ8YYGSegZLZ
nciTSce2WhLy0DTf9aKDNs7sJ60/brA00OHpc3uJAtEi5oPIztligNa/rovyLr6W
/HMD2Rbg482pAFNRZwGY3CeLw0t6wPuQlz0R9N1pE3v0il/bsMqY95CHJ/9KpTV6
vi7/SqbcbImtlH9WKbwqLQIVDKKSp8QQm9MWkxboTPXZbjdB1k+sG/ZsSakP8+OU
hT9LRremp1pEvYmxMKIK0NnC0FB9MRx7kY9dSmELZnu2Zml3Ym7T0tsEzsxcLcYY
vIe+dKGDkBhnWToy2hdnl6uVsaaAtBS4lVUWBNrfXVle4oG2scnNfzOk/WP9z+TZ
T61oBZ6ozqXwX0dfPNEnYWRKVRTp8+G/sNKBH96MKVsuzde+UXa5YSdCH7u0Ev8v
bUJx8UTE/wIdh4g8JG6HEvSmxuSJ++Oy49FEF0UGDB2DM82GPAlVyIcf4N6o07KY
UBplQqNi0Q6YuxIP1IzWK0jf6OV0UtPe3KJyiEUGOilTFNtFhAfYeu4JL/HFxzQ9
lsBEEHEo+hPJo74yIyXd8ZIQ1zNkoGvuTOzE8S41qJWD2SID9YLM5bMa4C3H1ffh
HmakK5LU6pFrA7GPvmPIvbilshmY5EaOgIPP6f8DgL03cJEbJ7gz7eSDI/BaPZU2
EHjaUT3UDtkmcisgIpS9z8vO+RsX4GyFdOz7DYcQ89mTmTbh2ZN7u7q/eEiogn32
FXt3gLAEs620DjQnTP53EsT3rx9nPCxcoAiFu+uPR8LU8SvFFF3BR5+HMPW4IVSu
WqKGpGu4UGJ5rRPngc7RTEV5TidSkao/vLgSGsF/L3F5WkJ52BFHV5xfXWiZ+jfs
sek3weg03ITtl3wrtYqgpCdmRI8dkC2akkoeIqJgOTovVo4245Dmt2G+kbqvXFXR
v9RecQj+/CgWzqS/Uea/O1VKBQMrDmuRHUffHbFPJXbwcm5bxKQL1tWxvQ2PRoKw
G6WOYaQ6B785YXOF1JRJhBYotjSMnqkZE99GIOx+pfmjftOJzThRBGUkQBMh+cXp
8HOmUn0D763TpqJP8oHXpH0723p+s8sG6pFB6h+myYyrx9OhVeTgYrp3HcBYa8n5
7XqTW6bYhJ5X50zJMi0zvWC1/EjBN076dtB4bvZAXE3uy/vMzipUu9C9bIWnZ9jS
DUqjlkB/y3fvsSTSOdyDX5p86X0etuqDpKJNC+bdZSUH5gpuIycbDGtTOEksgI8B
czw8o/2JdJ9X4kjQm0qs9tVfPBBuG7tTWf9N/K5ik4DlxwJXD0cZIz5G4kI0gPY/
CAEFLHu95P39Y00KCPWaoxmdn6pj/DSMhRQvoaSd4KcbXjI7HPaa1mr2/N882ILd
rkRO/SUxnqasmBLVWSWHrTAQMkcvFkjIoiaeT/HRAMKh7ZIAva7htCGpB2YHxBmz
4t2nnLJVEjnjP9iA3bdFMyT/1GRbQB1YkuZWbQ87nyCin3yxyo9Rw6gn6SCHxSNl
KG55arKPKBl7TpEWO3GT0ne1MHptqGvMSFBhJ8HJp3vKOnl1Y6zx2mSs4Ei2Cxqv
5AX/fZrN3sdCVdCIN/zmUPwhowPwu+GXidvygbJEdHDtC1Zr9hKyxBN/MYwbSS6W
djuWmjGj5232E+j2hBOoaGBBAtdGRdnnF/JwZsDghBLnkDubKFOepv6gHaDJD/Ku
+XJZtJHf/M6ebolNdDpp2tgRhav84ZTihM5lbFvCOTaZSVrfs+qd43J4r5mBcBrk
4k9VW5fZl0N9b2qMlUe8nz/jPA6i5XGk/BAW9YpgobVd3If+bOoqsO+lJzN3aJKj
ZrJ9BrnIUhCpYmqzECL3B/jWwYnrAXc6Z/QBtRcoHZ+O11HA+Gf4J3JxkjPNhaeV
6NBlq4KPc9xhr0GNRmssdBuGyHozeEJI52Dfm4/VCUy2mc0xSD/llaQPqKiIUo66
C0UVve7JiKezZijP90SWwfmVlaYYISFrG8bvIAd+9jF8Dg94L9mkfMueogsoLr4w
yzsUKJgEcGWi/+0jPzu+l7tCejvjULnvvdnMoFxdbUrKPz3hmTE9QKRe7vKugdCV
Umxx3Ae89c+BCj27nOCdo7wmkazYiIat9xBdT43v1UGYwBjuEu/QPiwcar0387dg
3NIajF2hEpLcXD+nSNF/kT1IacTapC6hrTur42E9cOjgdv4x2xgoqAFodSE6NanO
qUXgvAwrMiOSCmiZSTsb51JZX1UAg0KEbPhaR+Ug4GH5MmxNE6BV4/HNdC8OiAlU
ZG+B7Bf6BaeUCGrjrlqogqU8DTfnIpS5fMucHPr10dg0OOLnk0LiCMmDrAgEV/M4
50RZckgyoOn9O85JJk0ybIhbMpg5Sy+G3e4m4thJ3UFSgy4t+uZRq9l1fBCSefwd
QIa23kKRt5zUafTHWMmLHbzIE1WEkp8EsVKUlxOegXjH+ArNWPVDLS3wW7aH+wJD
B2JoSsIfufH3sh4+yj9aXSnJRe6xqA0Lwm2YD7ZHMn0Kcin447l/jRfcVpLxclPz
0mrd3nbkdfI0GSVpZ16w/Oe+VFVh0izMUeUfhcUeUzfAujG0y+lJBZ6SOI+6iLQk
tNDfkountDCw8wn/eXYhcnyFx/n4p83/bBWkXYGAC6Xs13g+SjzOjPVst+9y8jns
GJ4LT+CNSXO9meg6CQdc27n1bdQpe97TPhlCrdlNKeaS1PC55gJvGQwcIVLhj7Xh
YUi68Gts7UXPZzWMSWoIUCJ7OBXIRoth5zEk9ItErPh5+ZP3GssP/nTBf1Zv4ru+
aZBfB9fzpMqnfvL8vlUKjD1//VV0zl5G62b/8bdeKv8CWtdz8Em3gLk/t3BXDTYX
/E/7vCIdiFUjm1kSF3wjYy1sUITeSRlTawMIWGY1W4mChc3/wCbjO0oEr0fgMgMH
vDQC3NGH7d5gR9OwG4rOdS275MqNxCXZfKWKT3PiMn/3ymg1qBb3R4AAZy3odzEB
xKgadSzJNqXaJQ+KGwqhY0zZ+42W3fjOFpK1x6LSW7gcx5Vkt1AOVzbDHQFDOQym
Yw+1DipehLruQo4p5CQcnmpVlh9lBLGi/cM8V35ZvuFiWjHafLWLbsibcvdgFrat
5uCU992ZW4GMczqMxGTpSK0oNxO8DU8xGYwqr7I2RoHoWXf7DMXT5ghcT6YAfuIM
x0mJIg5+pw0yj2gA28SH/a38Sf0cl/thhzkHNs4WKK4/yLKE3VDao2wbiy9ahZdS
e/TKX385Tfvp23PtvxRpJezRIU7UulsrFdMJMZnWDA1IonkSFzR8IPil7AEJ8jyQ
FcmpSAk6jouT7MvYKcyaKKxxVE0xYUfPprnvXwBvX2FkNc2ZemslpDzJg+L30Ihc
sUCZfiO5p1NXWI6Cl5YS+MyRszKylijvDLySJS3b7B1MEuNfdtgoRjF+Hew5hP2U
GKgr8odkUFMsddPO5LrjzrpT3rheDM6W+3IEyxaqFqKv2o8sTXQNX1YJa7W0jjEX
P3qoUdo2/HY0FKhtnkCkWIkNhL8fqCiieBoOS/xvAzwfRUmcxiW+6SI7PIafe2lZ
CshBefPR5wRnb9cuWhW0aSOJfmL4K7V/eW5kRhfmK/L7E1xWVfZQQZZWYMXcXU01
BhKywb6dazjcg/svz8hPmGCWQPCZoSs8mPuxvrWbB2+7+I1/UVMM4Zpd5XqFnQYU
zZ8mtwDTZmuA4M0iqtZnml3cWzYebeHRWMi5TEqApbeB+5CKoA6etpLr3amPsTwn
1iwQgxYeqtgtZBkQyQXrZ4DfWflYy42QkLQfA6B9CgAawFRLaw6qroXPhPD5lklm
7rx3gsB3aIkSSpNhulVH1amW9//3v0C7UQqOYoSDL6woBdoILekFighz4tTRWOhq
710QJorovCt5YapCCDhnn85TSOrNwbZeh1mHOklIspqaTyTUuQ38tKMufMijnSve
z22WqlZTfUyqxUdQ+xf9zXUONjf7S+jHK6ot7KF1zUfDNowNibjdYiIaV/p654yU
NKJfF9PMbuNk5/3DuUh7Q2S0Jw/pQP0hj/dpVspOxKfVb6qCvVDjlTrcejlE5/Il
4bykkARXxYqXtiLX4hNWTo2uRMZVAnYdgkUSk1Md+UP2ycCUUvmzfeR8JpEsKILj
zltTjl++oSQfeuklUbewYjHunYxw8dFTary8CCO766qLelxGpQ9y/M1wyFr5IlFs
VWMjHQrFulyN51KMuj+7lFvgLWI6grcNQr3+byhooc86kqVsDx7lnS8yUe5X7WUB
yWxSwF94ln6by6q2piWInUywysYltXD/9XHtV6+feNx4L+KrzqoB++dB/s5JPDwq
fq514X0Q+EnBzIhgBSyF0iNQ8uWV8E55IJkQpkGwofcvwXpbATn/tTy9+3WvVk9P
8O2KgrWPsVM8xctgbnk8cPJAFNh3l1HYNC6O7K1EwchnVc8HzKDJfpXtxJUjGP1P
RlOmhQCgBkQliBqWWtt842FxbIplA3ZX86/9v5Xde0F+qfP5eMqG1/Pkug6aqIPk
vbD6h7JGDagtK7/+3SveKVgLWRvAtzADFP5ukHasaqgdABifjeogvqJJ8rplTXlO
bPgMd1XK7dmtdourF0sl5YEIEyYdF/WTP6YcF6nLLZtwEdKTPjbHH/e8H8QWa6sY
a6PlyDYDeA/QB65CcR4s9reDKQFLpk+zEpJK4QiqytJSfpOMvTQVNaGN+JPg7qRP
Eyl9TYjT7zhMTfW+0hOuZPlDeWfEIr6NRI+Vyu3d2KkZ4qIR/SRek81PRZDl04D1
yxgVKEMuNIdc4Wz7p14zm4rwrYBA7D8I0sgGu51MmPSN4qsTd+VaHmsB060pP6bL
EZgbP5m2eqPtckFoubnsFwcUX1y+YnwjrASUzp/gMz2uDdGSUiax5D3F1hqSMWt7
sDWeX79v/2NYtzw7nyiLUo5CsMmIWHnhfWNsS2s94AOy4v2LblL2jzRwAazwA8ae
9gIyFZkwXgsAFvno1fx/Tc8u26/+35nVjzNh5sqBL3wdr/a9ZkKjAIF965ujBQuI
FCDnNTwk3kG2PIdlu7OnTsHxXVwnYCWUcTP3p6KkWtdEK8orf9TRwIBeqA3PTk1B
SfzJHf0MJllFTAzA0i0XOliVPTCxc0RzABOc5Xg1EWUVRguj4vmu/EWQNH7uihIF
I2w6ENyQ6wQTui1p8g+YD2QI42n1M1Y/TOhvYv7nH0N5SN2ksy65k5oA7JHRFgjk
atfVcZhYDy0lPJSx3q/ORzHRRH6UpPU8weRNWQflb2UStvJufTZ1ygBYK6v9/m3x
6F7bgT44TBZhAkAzNJA2WYZxJjxeTvDWO2k02QwUKKBOjClBAD63IJ2r4iioE2NR
GH+9Y+0hOhdZBs/nN8ZoncSn2ZmzuSYM2DHdRw+1gg8l+Y0/fvJboI3O1Jh5dxru
U2ESpVaGOBwAy3y/3IVsTonS9baI0Bru0LM1aakT39LrA2fEwom3WI+/TsY5fCY6
2GFTwX9ml5lkLODIi43n3IxMfuRxVEd7i9C/Mf6po/uOJG6kjxOWGzw2nNWFqMAA
pbRHyDGEFyeUfuNuRLFshI8tWdXdxXm9/4M9o5c4yC5I7/V41pMBZFFipnxfVNP4
6ofUW6//4JsN3Xo88QnCyQMZEUP81S0sujob5IaIqxi5HYpFJm34Eu4GGjcJe67U
eUzYLYU+V8pW37t1nbOF9E/D/qOWnh+Bs1IKY5lzWR9QiRaOTw/rQdoyCy4bxuf2
1JIMnLC+ErXYrVXO04uzEvlpkY1jjmHYzKbuX+a6X9duJlBcuLJoFYYDwQ1KtIdF
nHY4QtyMWG35F863N1IveCu3+K4nT2g+Jww2CBnsBOcX4Li1wC1XxzTwKvB2FI+/
Yx4mUC8yqEa6/g8jaqML9WAoTEgDhqEBdPqUx42vlebxCvJOq+f7FN5sz3FZwJUN
CaGY9ftLi4Lq+ai3wutF5foVDDmU/bEVIUA/ELCW0741JOMzf+KhOuW1V9KRvSDw
DpEqVVvP1CXrnbQFpi/MqcA/jC8WKcQkwyqndVB6n3SrwaAh1ZFcwhotc2D8MHF0
g2WH219kWWD/VSrfFLalxMF8q9hsnBgXMIYlr7h3ADmTCEmg/km2a/8YuxpoTqKG
+B/dfw7vYAWWcf71Xr8gtjz4YOetnotHuOZgCciv7uWSnBt4fg5MGy5stoVda7u3
+zKcgG02S0HFtd+ETJacF1Zhgej2DNLfOE3Bb7l4V398VgFdW7A3TbdtNwRUSAnp
zh6CALBUYolaxG9UAPeX9joqzEASV2gFy/99nZ1qk/f2PePX12x2uRBZsl9Yu32I
FbHNjCCfR/F1Ab5MW3TXrMET6oDbEUqudeaWNQq1Btc/ByKR7wNiXLeaOShoZIee
8Eqn+N6Gv2hAGA+ligWFVWNpIoOfQZIa8VsNsp0stKgxTlNOD/DMReAOLQo/ByVz
MWxN8MPT+M9U8cTjGFtS7eUkW1kbVzoGr33eX/yp4A0NNdqCm4Ny994R6amQS/9D
tDt9hDltGyjFC/OGzg3OF8qaM5BZnNbtf6XP0h2SKVPS/hT/1ZGzFd7Bn0D73IyK
WVh5LxzjK84Bjmig97HDVC+nOKKDJcZBKQ9YUXzN5dHyK1G/GsfOi32vUOhJX/ly
wprDDOKM3qrF5Psi5XMpmXa5snfIXaJdAHllmkwr+6COmJmFLEY/PwDq2k4uA1vw
YGBRQJTOz11b4gmKVhQDUmv3m1MUQKPgt4NKejYfhw2wtDbb3qqNHRzjhbn7G+oz
EGHCXLUx/R6dnTdjOEoeaN5f658uz1u54CyK95eBn16T27sZlSfkSxIOpa2+m5p3
qIvimuYGPcZBR2QRQGzzdIGjsGiTRi0ubLKeLmDLonUDQM73mvhgiQ/PmsLX22pS
qYCxJSd0UHodHY2vJfdNUr2wOdamikhHxww17AV/H/2zxtRjuBfZjjRkkt+mlz1G
H9fIeeLhqYg4HqL3OE+eIAZanvvj8jYfJdyoapQ3vEO3CjToZ7Laia4GvAebDB2I
aPJRQUJuPE4nFiipS6QHMUx5a5W3h+6xpDBpzzhWyErPi1v1EGWf0wL6BFEYLjwZ
06MbPHo2tBGoviWl4sMiIFjFaUkKgZyzEIOQdRwk8SFmkNxJNM/sS1jIX4AC6P0z
d9Zo0JTd6n/ugVVsaHcSjqpcIIubuLnEljb6jXV3BiX54jgpDiY2SgEh2vnZKYgl
0wFlZV6q6+xDN3gAuZ3Uei7bjdIzjDqLlrwqcy7G0FwIXqMf7uN4EEgDwoBQRo1R
sHf6DmFBFhTTs+eEWHTwSaWz036YSmk6KBZZZfBaw+pv5GPfxdJWnIy4dPjTNVin
XNDXGQR0C/v2WDvR6KmbN+pZEA8AFNKTBdwpW0luevfhgko1fEvCAmMZ6h/BCN7B
WW7Yb1NiGDbPYLyxg6RDA+cs6DD9iWoo07PBjEJ5wc65FDh7yeejwvPkXoJ7/QhV
C9u8BVtu7RGe7yJPr1ZrB3vgiB9g7onxhNOtwyfNL+FwQc/wouXUCFyAU3IHRjm3
LreLlcB8zSaKBjAmG2hwlXrWl4trPMelKZG3rxfvQ+ZSODDptEln7BPTUjwfuqeq
rzzqXHmHwg0f3kRM5HkOmvxAHbUYSkasRKdPeOc0UlkEi8tKUKsCll4iNenKqwH/
AClcxrVClkt9nUAZYQAlWH8Q9mULlI9wdny6hYNc0EJ+ogYXNM4R0vPut2rc1lpB
RdrA8j1+XIgQ72EEcJDgx3GU5S4RU3wkFWyUf32AWON/Rv9oa0jK9W045qG1KiwF
KVgAQHGElQ0Hdi6xSNYTXAPaMtt8ISN80cwKiuZ1lBtYS8hwp+I6U8mgxMUVsCJE
TJf3cjOOEapqD2kPUOEuuYTVbx2UlMXG1uYVj8omJC35wAYHvCGgzU5nHQ5yLODv
M2yk8TuYHIr8+PhW5u9dcVFt1l/UA8V2cf8rBZHfVccHsNzXMc16yvr5btNo/hg6
cmMxWNMOfXW8hKkXWqaTbBEFlg7IPoDidTWgeHBSYJMCrIjUsAZBYkEGtCJHin72
dDmJHRX/6pXrpYHYfItRJdIrs2Quj5eDDlwCZJ9jO+uwpcGboEwjbWv7rIuRngFN
tNwrWwHF0gw7acLt0XFEmN9AlaaiLDcekEXQ4Y/cmaHNksER2nHX07+kOypWAWFm
+2Z0N5K25y7Ue4X0tLD29RGeh9ryYpMqADRNZXS9adFsEq+Z7qEdB7pk6v7sgywc
D5Ht51l0rA3d8wLXNZHXIbnIRyQYWHYCYxTM8F1JnrlI53Ub61j+yUcPZ1KRFzQV
s/wX2jVrAxzNKtJWiHCTEnr9XKKGz6N21O1EEnkKShYCsLuq4HKxo4V3ZQ+gwsnU
CWpzC+q/kzVmH2e4WsvMOofaGF56uwP2LrbtI9Uofxj7+s6koRcCOS1okf5Z2UNH
+PuFPHHaCPYyKoKBoUYApC5ft9V30svLZq64Dy8SAnzJpv9p7XtctTUWPWnz/Um7
BfNBSvSgLBHioVq54XiD2G0kdyW2xSQJX2b1tCaMbUxqDE1F0C6tsfYGwNUoUa/4
aDeut7ZV9d2vnVU4T5N7QkSwp5Imsax48zy9b982QJg11eUBOEtWFSg2O5L0xAq+
nRbarQXWT6/1XXF2Y4CA1U7U4TT+uLbuhW80J7lGDCaBOYTAbV5FaGjUlTK0QbX9
QdzH54Ri9MbMUYPoxAS8UNBoOAxHt61gzJTRcWBTLwQndQd2NxzdA5RU3xmPmPar
J6WA6206mTLFqlZ6ECnDSf7OBMBLbDIPCikPvocx8+j4va120zxB+qru4ERDY3UO
4XmUCn9Xog2KKjFdA4vWVOHe4P2GYXSB32pw99LWgWlkz8uRF+/bNVs0bqySdrPe
+9y/L3g7NMzAyTmYjcMYXOPA3YlQs1uQFTqt06O4u9arv0KxnUbBhoaGesUuENuj
3fJULvDrFS5OHmFGkkNZlPsTHhOQFHEZPmwVCSeclDegbR8aJqp5KNGb5wp7oLDL
jmiqnFHnw9vfbGJI6Bqs/yORQwqPK2bLIYCCwUMk0BDMijDL2HEeHZ1R9D6/R2YH
QkswZN/efCRaSgStgyMeQfRIviXiqunE43WatlSBJ5tG+HineMFdeI/Snl/sop6V
W4RURJnp9BvbiPhTf+lvU6sDr7AYF9dawvy2VoanzuqGiwrN9UhJ1uFh88v8i5eA
2wRojC2zpkyvw7EvKtHMCmmWQfrKVo/v4Xi8pWcUdY/FWshrIoV59RcjNnzEg1HO
i9dbv2hYF39Wh8HYOjTMxAP34NJ1kpxnFQ6O09r5d+JN7CK8koqcAQXvKAviFzWa
emGN3OM3VtbS1OGAn/MZ6ZP+o7hiLTH6eQmDkw4ENLglDgGqThgp/R3uihgeM60X
BGBBjT7eZd0xU9ZC0JUCkXK/Kac2F/rNe5SECYj1O7y7uQ4CewmbS4PryQgO0jLz
Er+DPRzGPDpE08R4l8WEPvWgiZw6QQEEqkMi3CUrkWazbz+ugCxNLAMLKoXUONKb
H5wbT07ZDJn1cxqDboRnwIxlXkcbXsO7GWL8V8QuO4mN8WCFg2RrdhL4NpS7Fqrd
jqZSIdwr5cD5KaGB8ggvmyoFx0kH6f/ho7zP0IL0Pwc4sGxFniVHHKWSl13lwid4
OdgCIlw0iC+ftlZQ7AdWhpJ6IsYxyFjLHcIlbIzDS3Op5bnopMrEUTZtuSZ8cd8h
5ytrxHncTdjas0CfVzsMQCcL6yTZnaGnzgwYOBFK1/SEGrhGJzfmk15BxGNE/5Cf
7MkprV+4qe5T3Yud4RC8ZDGe2tBMGyOS995QJrx1g9GJ08CByhi2AMjUJf5mKnWD
Sq+bvp5ztPJ8C48FD+7lb5YHIheGlHD6rQwlKuL5a/srPmF362y2Gx0dRK22o9Qo
AukfuV/gAXO6PSqmIY+lf/QfS/W75AEe798+zuSl0NCcTju1rV89GLhXNTw+hByP
aL9D2BDHwdp50l2NE4Bx1gnfjWgfairxXU4C8X2CuArPKoKG950BcW3bbfYuBAOO
r5l+HZPZ+0ZxWjhlzP652vSEGfad/zPDBmDubfpaosEToJ5sLz627v53qzdEBNLM
8OLdbQQRqR9uyjQpMH+kuTUT1Wd2nl53Mg++KS1ORZ1AqOm6Q4IMyTbR+q9VXe0c
m2UaqIzzoczjpBedBevF62EMA0mZEwaviVvEgb+Jhjkc6133ZLJaKPCGxfvV8qFx
huoL1oySm5eFarRIcmog0FJFbSzmCH6c/mLN/Yd4ZNTOaLpMGmcI6NKMkJ5HYLbc
qnJnd2itq8+/QLZGNG2gQdkaY8DxflSO/bWMKfNzIXqtYdiqsJC/G3AMgfzZ/paO
eSub78dWWjYcj5kLimh36CMzJhI3FwVu0GeX6CJuxxiMvHALCmfH9h3ilmAAkIRs
wpjCI65slEX57xOCMLX1bsdCyTQ5VjaxQ8UPSrAECpMK4+YcanbXdBQwziPIUZ2J
DkOUH3FtT9dgoQmfNnXuzeaXyevqLpVErjF+EZSRQekkhv9AOwIzV0hMYanNWXCx
AaqW97kmnpMkHehZg416RgDYdvrNNmaWq93cxZOBTr62mm/Ojcbjs9HbcqDpx9YZ
vqAVRDEScgSeegvrBEFCnUBnbWHIYxDhDV9+9hB34a7igRyujFYg+l+bUv7RIYh0
VubWizqXlvKXSk+ZgZlRsmf7YkO2htBUD1CfCRCDWvNNyFnbVLwDtAqeDVKxzdbr
DXU+0SpvBH4Q7tI25oWwYyDIoosfnl5HjtEfiiwwTetj+Rsb19S5PPLTIGLVhCd5
ZDiulHFerX6QTr93zVw+64XxmA57RgBhbmV+wvIEudwIUnl9tbhpwFbmGbs374mS
PMe0sd8xkS0vledwNw46/42Oe7cYx4oLzUM4YVLPHRL4Ehommj5EfRJs068xhW65
G8VEPjxK/KL0/mvz1V/YRLRxo/I1SEGVWrPmi6egdRBIWy8AV+W0rUOm1CfhbMBX
hIHWJYkjs268NMchjuOSiGNfd0uyuh3P55bm0OncmnJHSrQz7IdlyBZx5QSPnVBm
jvLnXNf/i7yXC5UXNTMOWxkAbgQg2nLiNIK6nMuliaEUMcImZ8sugjdXVKVdZJuK
wsF+pTcDr0fVDGKStrTDJTOlx/QVeyVTnYjudOtK6OeopY9cuknQdQNhipf0/hwY
4L1Tl0CrV13nS6Aa3u3svOv6TwXHFZM+P3luEtPm+5vMcYJiPbQHV4Qo+9O3R6GL
IdUiRXc1zu6gl7KTLlv22C0zhbjaiEFeDcfzFTHwy+8hfeC2EXls65MHK+CxuhLq
/BJmLr51lrq/D2tlVYpATjc8xqD5pPC6zYZIW24vXj+s/YGSwzgyFolTwKmsIweS
J8/nnAm1o0Y6OXfwB7BEUte5N0VmrWpfR350e75YUcI9fs864TTmUrDfqAtOvvxH
w6PIJ4ZYKvy4sZ854YYZ+ZZ36NXhlcHr8sKqHwWj9fM6BtOazifSB9/RmjzmsAjv
50vnsx+9199x5QFQ8ljey0t5a2/1VZ5939jhYeFx9TwrP6MOsdndhd3STzfAJ7pI
zs5kre3nq3lkp8Bhgzhfdprd9RJk+HucFKzQXPN4p+fmXd7nBinaiKW4wBgP5mE2
48wImtz5hj7D2I3b1q78Qqf11JNz3O+sGfhdm85UeqeHAfFcMMRBCgV4RCHSWJy6
Rh++cUu7hsXh5107f8TSGG/kPzSSG+9emw+MuC96Yj6fbGudsdYtPRQGnIBZThYx
BYf1Rfj6CfQfytp0QWUWuTBdb+QU+WG9f52CGbniyuhpty6pPnP5Um9IUxXbr33n
A5mOepWR3qI2H+mO+ELhdL4BneyiQKg7EoK8RV3bB6H0hDSiA7idN+wTaExtI47j
4hJUkAZ6HmfGn5sK6KLhW4fRVndRW8jDUEouNRXlE+wahdHB5rYmqXuHTPLTDdFn
gs+o4eJf5Tf7hKukTuMdZgKKoxc4jDAlcpabwp90zhAg0F4ZXd+cwPQ5Nv3RFW4b
xmCfu0JZ+wBmQdd0tY/vo52mQUs10yFfVHKmdqLQroadbm180e6OPkk+fcMh8izp
/7l22rzwdEMSuS47k8FeWCqKHCddxNsqMpC6iNlD4qXUtFpE4bV6/jtPPh0Hucdw
9Y4kgLr1V9cEzjtUWLtEaIwJ/v7UoqbrFgt2QMOagIUNkWoZRbX8VM19DyWDlMRP
F8Cf5Hj4C3K92fQAk5tsNpnn1bIFJwmI4Jt9KRsweBK+YP2hF8BcJC1lZjGjz4dV
MRux9BTcLlfrMJxp2krjDni+WOllO+lo0AW0zAr+rkbRNydruNzUZdF6b6ZvsX2D
ms+KjmY8b4kjoavh3jj9/TEXL+UixwBpLZO5aMuzViG4UgVAc30X5833aiHp5y8b
0qIcTxODduJq9hIBS0jtqfVKwWbZunug5dp60aB+HniljpuQV9jTl2nourkpZlaX
M3QwdiRH/E5TR/1KTpJQR/1EU0mvAbmf9REY+MaIWl/FnyPaDkwgjVRtzubjTzQy
Suo7nksO4PfUaq9MFm3SeyBuLrqQo9tPpsLsyYaFgoSQKMDkntDUhH0zoR9dwoQe
0mlox7ccMW2NzP6TAsddna4Se44wqrFpCROMctuWzmC5m8vQRTgqJgfkEbZxOU7H
Ahi3DiAFRvdADTtYS7Is90QvV5VtSaiq1uNoQjVbUfz83OCnY7tnaFwg4EzWzuAp
ThMP7xK6S6zva6gVoTHL01l0KCaE97iUZ7tnkRCJ5u1SXdMV8GBdoswYNyYIuq/Y
XTKfkV1u2Pn9R/T2L/LBG/Nc27xCqJOa8DnXSRsSvlfte9aFtsiln58wEXV6cHAt
evPWmuB+OBuYHsV15Ex3uWb4YLCRBGOfqid//K4LwdgApA2i2W/RDd2O69mx4PUp
AjB9fju4hd1SZEIgitEs+lmb1aGHrmqZs087gbH5CIbzDRJt9OPwmkD0WREzRS6a
/cQAPtsNoBHrhDA7ZQDuVwZel4f2OEYWXnIXYf3Ia/PAD5a82A6Tuxt2jk7KmOZF
hHychDVBK3F2idOD9QW0MrA4LGP9AxE9v7pZp6k+ZG/wsbP+7bctR9Mw47wf1JJR
Xh8Dp9c6iqN4bcg+IWBNdu/HklLiGQBOLPEsg3qGCK0ZBjzkVBlyMKzR4HKlMmuf
Vh+rycVw4PlsQFSk7pVnNGDQdRqYRo7JkLOAM9L95VtQY1MF6JEF3tCPd8fw7b4N
8R20oWSGEd0Pm5fLInfSuVUVMypjEAAgu5pFH179SPRAtcmMF2WbeOTQUg0bHxkq
iQAPr5aYbZbbGEWlf0eVREcOMBTbf1ceUDZBwTlG1+DM9jp7cFh12WPdHPg2p0V4
G4Z1mbNu352leHoOGZHEe3K4x+rV9K6KKjKvC5em2YqmB2Kt3T6Muzbfsk5H0bWK
17xl08Ye1r//eKnlP99PLyN0NnbWKVjYCul/bUdmuzxa+kkrJIxxyWCUuqh4M5rc
c+z2uOEcrUORwdqF/RZEnu593p5RuLR8XvcOoxRM2Dbqisdc1Z5NOnlroaDfasls
st0vvK7dVSJLFIuZvA8Bc+Cu0CqVd/6+tQvlgxayIpR2Ofpjj7qoTCcgm6zh3yfG
Fc0oemC7HSfa/joRkQ0sXx02fXP+2vd3aoKcrbn+GF38jCP2tygZzbVgLdHFf2Nx
mpcIWIMtaTHBR44VMBuJGA+vXu91Fdm7J4iBEDn7O7APtLyC6+7uc5h/LMTOm8vZ
hq0bjfD+UOErCv61Q2L3P+LrsPkg/fgK9SIJLi2LUpF5lI9c1yUGfBMkigozc6bh
jbZVDcUqQYKByCTSSfqwSxl5qbarsQHedQ5KX9ejEBgUOiTTjUTRpQpSS1q4sJ1L
H62ajf6vsD8yqWXQjiaT0JLl7yiqEHB4A2LJ6OKvXuHs3ITciCT1Hr490VL9nYNb
giM0mpMaXetTQLT+LzICV8GQsqlhT3CjsGwAS3Hb3BODIpNJLstS6x/oTNrgiJ88
DRhGNCBASplBrmyd35DegFyjCD8QGlns/TqYli9WMFoVVMj7xTOf83qrKmCkC6uL
Jtbh0emwP+hdEkFuo837GP0GRnAcqHLOyIDoS7VmoGNsVeqskafZ7RabY32pZ5i2
xJFxU4VWe7QP1a8NOM70odj5jhHLQPXvFF+7vYc4cBuTmanrzxP2w1mg0gHGV6Ty
7twqo/knye0XAliLi3jZ0WfUNuPYbJuaI4cteEylXlbsSJndBtKTbc9qJbvvKH8A
ptyC3eYO6ngJHBpQi5Ky0G+RxQn8bmNeCpdDaY8aKj5+UpUVfYjvcN4HSqPbNnO+
p5NJotHZGARANplLvT69umwKHdGPKpzfT3DX1NkpaNAqmWS4ZkweJzdxAvW1Bs0J
bc3m31sQBSCXvfELzZCX4A2CjS3/EQR35C6YOkZtgiPJ19PPg9fnE9ke6FRHu3wn
xRYgmWf3PJDRQRDzwRlT2r1HmztPyPR3LVKwvvWfvtTZvhJ/bLWPaGXtCw64rY8T
Pi94x67ezGNV6Q/KwkP1donGE/c+c8q9USuF7E6g+/RuWzMoq0CBCo1u4bHHa2Z7
pF6sYTX6gIl3aQ6FzFgF1eOvrraGXtJLYpsfhgxhudehHIrR39Yfkpxzvn7AwpCK
BsN3Kjh29rlQ/5qojcfrwQ3eKtFNt/JZhoQIeV2uh7Cfa+tVDEtpAzkyqIeHf11n
TTpHqOiA0eJPEw0O1jBlonpqPP/33p6d2kAfg4m2rVGpig2ZT86wKcX6yiGi1TGm
KLIRuZrThUsVXCBF9qJAogkXP4LN8hi4DtojhhwlXWmzgvJv5HTD2Q0w3z1bJp85
xmPOIZiDMECIQn9wq/pEyiaUv111vU1GY3gck08o9vdPq4Q3mWT3uWmNsfjsMrtA
8JhNFzcW3ey6Rkw8oN7IAlrU79kduf8A1BoANBHL0YL//Ypa+TpIOqchzRySLVI6
jThr+0EEyFn5gjgieRm7gVIR2rsL9IeTf52GAYYyic68c6y9Q6D0biAGkIl/yRu4
4Z/Ib0gQiM8RSo3sRNFOqiEBAAnRy4vLjdd5hM9ixVklTbYQ6rVGpMw6OmsWcsth
obziHxH8zkK0Gkj7vlqqIcTI/D/woToIbQr8PkeCGMqM20YCMXE0R6JBTvNuBLM8
Akgpp3ToTlNqwBedgB2kIKReG+sTG0HCQ3F31o9hW6uC+4MzqvlFg4HroEP5c37C
Snmh98RVxJdPYBl2mmMY867UW1xHBoIXpzJjcPbt9qm0U9ShQ2yXq95u7z5qIhwH
DDG1S5Ij/ZyUoim5Uy9IKetkZVNh5LxrDpCCwMWwIxldLZLDMc/Gaw7YhukGG2cj
BSR8o44rCueRu4IoNiolDslrfNdTF/WdA1IjBZxv1PqrywvMHykRZkbwH7Rb2boO
rQDFlRFNhLa6v2vZB3YTKqJ2/8Lva3wiclbBLkh6HKjQ4VZBusKnAUIY/bKjm+1d
MYduQ9XwZTG5oHkKBJB9U6tQWnlu0t4iBp239XcFVhJ297SuJRkHwBBGaPH/M5Pq
LQRpfh82rsdEabLmica2ZtXph0mhdUmQNDDFZzIBNEYeIZweRrAto2huxsCU/hdm
O5KKRHfbYWgwu2CPJ4JlignAfjCC0iFp0mmwspdpbD6Acg52c59n94iO2bv7Szwq
HM698ES5Mr8ABDcCML3B15vm2k6EzuxXZhqOfuKFmkPcbIkiOyfsz3l/OQmATA5A
IQmQpwFGIntPMbcHaVgDZauFb602F5P/UFoCvLPFgNk7cvPCc4MAALYk120vXSiI
v32cVa8W6sUx2/Qid2rUqPybDQ2AnufJC2MKD6cVWiP+X0TOcm129nArmW9WqZpk
pCEcGfzx+dCp9ZPSJpWMW52OnflkHVpF4GR305qEwiZWu1K5rAVuX8oXGaZqFnfV
kTakDrRWCNGFK8ckQG9Av2h8qYem6D89tb0fR1l391cC8L+ESM6xbFrbGiYgYBjK
uvcd+193GJDPCywKD7LiBWj9XuA2J1Rb3k/KazQlwnwL00NrcTJKtZJnv4cYsRBG
/vw7reJqAi1bnmEGOVpQbPvfSKslTzOfGplES9SGx18sdaCM+AZOSIklkWZ/+go4
eVFFDBW77IPQ2LfRhiBxT5xkMK6+OfwlUWfhqAvdNJ2N8RNQgRIrf6qR6MO9J3iY
ejIDG42D3MC8dcvnBE4u9vUhHopJgZtm+PvJ6KHBJtFVG0FRiMM14BWGvt8FNhu0
qeepyE81LO9PQ4MB5mhnJw5tG//T5XVouRgvO6Bn4doaex0aZVUBKwA2K8OlngMh
x2nWUpx6mNuEW6AtuPr7BEqjGZ78ValN3FNaGOf6F2QwokPddqJPRVztS7AiMuaS
LFovI8MpeRwTec3lSi2DeDsUsFevZG8UsovVODKDC8IvVy/KZCTqerCJtkM1ZS3c
HIkTAwOYQav8aJhYeywkLprjb49D2/ZwdjEVADIahlKlfZ5PIxWTuVFn2UtHgVKd
/xiyJFKubq0mNJchUDr7lgmkG9n9ckc/7ibTa4ofPlZuLoa7PDWo6o8r1gBhd7AP
96qeTqU8NdF54KXd/6b29yiAdmueA7Fpw8jNWYEHfcbKs6ZpeHBHXSx+Yo4CMiCW
Uefu1QzvZt34vQZUATaOYmAL/U5IE5xBiE0aCZ/DajQW/50W4Se/bPw4+LR1XqV5
TYnLAvtfhrVmB58vLic2Joz/hKakEDrGlWGyB2BlrhwWKk+bkuz0gdeVkuuiBOmH
LSgmxPxF5dVRyala3M5050F2Hr5quDtGgjqcerGfG2UyqfZedhYSMDOFVYhtZL0n
UL5maZlaOAtrw1q+042JbLFJkNdqf8UtpSnDMV27k4i3CWt47fFS95Gmza/sdqUw
2dKSnRK9TTbKyVyIFJjAyxrkxaNiZsWXvPgQouqAkz+DM5tpcXYfsu0xgJMibfSW
G43EoExHPLkdiYeld5jzF1c9pyP8AE5cJW+YShmytWNcBdzjAB/mr+4fZIJEeP/Y
xmQICdZ6Qh7DAzfsJTn5swm72N/7QhIZrkHxuJ2qlPLQsHh0dxcLm2Iq9vFnYRvR
gM8B2PFOQ/faX66fi2wE1X6/Ie5Li6Hra/nzq5xIIIsuJEZkBAI/KIXyQFXUOnTL
XsMaI4XYPSQ4f86TLvSZHe1dG8CRemt7xYDkDQbEp1tNgXcc8ao9VDZqje/hC1tf
dAHZNfGlTQgnzv9X8FOqH1y70o107MSzd8Nk2QrYjqmXMnDrNo3OPD5bxZ2Ef90T
dOfy+N734e0jtc0wv5Qops0kw8yhJLJTVRHJ4fG5A53yzL40XMWdcIKFCdogkgmq
deDaQkZKWeuF76ZQGChaor+8ilcppku6uwxqNeGifuq8h1dbHSF0WaTRNxltTmoo
LKvPLoo45SoVTEyxumLJN9oSmKDAcCJtxTHE14jMTcbnnyxatrYdTFnDeQh9rdgK
qexzpMw74/Tt7xzQ+KAJsPx3I95DGS/HB8qOTiZck2IYj88VvjVqVuLmGI5KjB1o
v+5SPvBNCO1y1VMiAbjNymkd5S2fNfvN+n1ifFXhUeLBnVW7EzXjDEtARMBa/lxF
aTyi7UTx2zaR6k+kEHHH8I4jyAduRblpsuhDRY1CTP3cPQSCVZA/stvuay/VurA6
BcSfYCF5eP6efmPf7vIwxmIcrH3j0IPKz7U6afKShkdaYFVcE4i3gioxlC/3G3Wr
QsSPyeKmXUL+U3V9AUIHV2hY/kPWHZzIUMq5wXKzpZpN8lQnLrlKFjRssHOgezBq
VdOwCx+xHWFINw7NyKbCYl5Fy6pFmpWBNZnEYjYK2+g6EUDE5KxKHARgTQ7dwBO8
PoNQ3ZxKgoy9x3hV4pNY/LWUhJ3goxaVABxqBty6MEMeGrb+cML4MgXgrIuN/Dh7
cIwAVW9KYqaWVKVGc/9G+0LZkdZqgxUrPYXIOlrhyZ6W6iLUi0z3Boj9xLdlrbEy
QbXw7nlfNuauLeOfrbT4zIL3tREUnd/NWNQUFKuWm6ubiw+mKpYV6lDY3QACd0BK
/2GSSnNmYPVk7HUrlfJj0//hFcHLfHcQznP942BgdQSFEm5XFs53uUFPtHgBZy2g
aIubCyVNVQ1pUvqHJrxhtlPtGgdXKaXTBYpYjbjSkLYd+ADB+YsVOJyqbybR9xGn
4UUEqETF7UYye7lHzaFWX0a0sQxaWkzwIPDlDFGKAxj0bQW9sDBBFyjU1YIXfQNm
9TFnfbWMKLisG6+ne3oqFPL9bu+k1g2vx/CuF7o4zSTXA/exgTGkYc+eugtJmNKJ
LHIzMiH3n3gYyYMtL97YtLPvhwUeKbvQ+DA+Mr7cdPUiT9+6ix4xlPsHTteEE5j7
Yrr7aKEmXgnytmDoYqGzTsGdOrHcaLsL5Ujku7yXLUG476byeEuIT7HSpLpKPxhn
31roKLqp8oWygH0BVNrSo4HPdyOww+FuR83+2TwIQPkb1P+nIsAny0wlodVsQ39d
XRPjUsNnMT115aZxisW8ZwgM+xyqYmEc/nGKEQcjNtYdhb/IFbS5pNeyG24ERDwq
nY4NUJzuzJ9ujf4I0DiFYy1j2lYIP/g7m4Mzf27GAXuW+CmqSSVfEiO4CiUfHOGP
3Zc4YwVKLAGLbFsROl6HLNaSBNbQccLVpRcRsLF2E3TNhzZrRGQCG6kLNzL5Glar
u6dMY8fX4G4Af4sSWDQpIdhXnHAboJWFCqCrKCtISJFkjAX0SUq+vwTP+NCPUZiz
D2STFh6jyj2x+b1yoWTxOYteyA7c5bnGU5tQAlLsM+S209Jsx6+A0dPgWr8cPdBX
hGf+tbT2G+dPyar9YSFnbecHWoevVCVf3ocs96zmxG+Nj2ICKBYq2gQ99IMzOxFw
SKZNk2iQ1XuuSPNSxe0k37XvNZFWSMBaQ3MAhxW49/T2aXcnaHua13uHa5YJm7ey
7H+XKRrhCvpyMCPm4tkq5Ow0Pai2DsX3Nv9z+9OFumNL0PAppcvSUF5qNJpWUV3H
nLAiqXM7T6kEgj7XegslV2nGEwJnqQ/UQQJ28eim3graJxdnTTdvMhWcRbGGqblR
tyTCZ9q7ASOr0yYk0DHiFNXPEkWHZ+7+TL5UAooPvLOGMGinMSV7Qtvq8R/srdzI
SG7krwIziKF0hofOJqNKhH0K/C+6QQ0ux/xLA/ZhiSieS0T2aG8cFKsG1rzpLlyL
QL/xUt+eEwgJs35EU4wtMWqKt+otSd066Eu8i6jmE0WMNE/8rMRwJgw0nXz8gNHv
BhXb0k6noU2x8/TmPIbURXTJuOiQ3CQlILyth/1Le0rP/wiV5zqK/qH2DNesa/Fb
IqI++fylU5J6w+gB8Bw7eX1ETYkRJor5/y00W3Q4U0k28VK2netFKIPHP/+r8R7j
1cO7uidCh9W26USU1RyfCif2jIoADmnzTTJ+NnISR3Oznsl1g8B8mhJfSvYprsmn
/7JW4oMVksi6iSm8iThrtkFhQyGjl2/F0I93KkurF2Ejvd/gg1Yew5oErxz1HlDq
iEArqhSzsPm2k+vtM+Zisnm99JNykROuBZu4uFeWqyTZxchqpqoH9gBqHduEatt3
47HE9WZrYRH/D9gPSIaWY1P9J0eyiQc4wdYs7ISDeg5UJ0YjVE2cQXQX6kPfLlyC
6D6f7E2eC5gq4VdxDCjIt0+ACFFzEZYzyjv0W/xOf/pKWIomhmDhOm5O3bganXNk
h+8thj42R0GQ12iD/zmnCGx+KHFjry3RVoAvk/XDIi94EiQuPinXbJmAk3LC9iO4
EVJW18RmUbEOnjmkxt+F6hU+XwCB2A4ZJpeaFa40pi5FhnwQBV4lWZrAdstyeLv4
3ZY4/X2MVOAC+64mZJCPM1+YRCQJY3UJw2T/TTI6mkfF+aWGNDTWfYBDCOIKRGrf
uITvFrY4EMTstXEiKhOYs2o0WdwTrSqiqKpSujR17sN2OI+5D8r2xeUSaHqlVkd1
BW5n513TpNEusm6n9BzW7OgSBivqNePQg0vp5wyUKogs4sF0HTOJTGCjAodz03p1
UHBFcfgKlpaenaJt55dIrAxbYRXt2IDN0aOZNe6rKlbt190IdePmijde1BM6Oahg
NGeQpLJdTNdM8epMiqOx+iUETkzD6VsluT4iRtAtA7zxocyshQgKXKv1KuyYfTl/
6uFKwsjwqu+KGAYAPdD35/OJUF02RcUZwlC5N4ta5qe73zs1ok2OKO2g9mZzNhcr
ZUPMSDE4QQjoP3p4JtmHC3HSAxCBxDZDrftCOkzvvpMuuHjGO5FayC3jVA7TCxik
1GrNyCYeURGNq7Ksak0HNVAng2M/V/A1W8LUIkjAfJEWLp4c9L/90/i/RmsBSL4+
FMs6cfjOMFuf7tLOWw+Hp/kBeS091V0DIKGG2g9G3cShxvSZV+VA13X9vKDAWiPQ
Tlk1LjU9oktyEeEWh2hVrcqb8A50MaxyrhFwH9KvS+zVto+Rzue5uapkNm7XrolA
QVjGDoCH+8yNx+XeYaS9+4qWNODR0crprS3AT9Zo/1dejMPlOA5Tikjf+j3SWHiv
6iwYfUmOFI36/oAKyO5bRchBPakEbqodxqxXUQfM2zqHwALUHT8UB/tHqxPzjIRp
TpYe+VoCR+3NO1rQjn5LG38PwkLlUALpcOzwp+aHX9c/8WtsPHFMJ5i2ktWcR0R3
TifLEwrBfkCgUJ8H2QjgdguUkDNyJJNE+5uS61VyJE2+zCZZyKk/y6NJwCzwv1Lw
CNLVDQjgAFkQFTbNZsutBIwQJWmkpgfLgFnFGk9Z9yJSixjbZhWaddV9IeV46FYg
a0khHQu6eVELvxJuVWyYx0UEEVphi7tYlU2Ty00UiXZguO/AIrV6+gT3HoDK3NRU
5YL5GgpenmWg6N7qeoUFyRbhshZ0KguquVf1HNHllkzP5g5pg7eaFnQxKfN95jny
UlWyHvzA8DelcQRVbXm+hVfpX8SPwg2IHr54P5F/5HpM6igh1gmJaW29YymEYSAg
thDTYmEYsSOUCO+oDQOD6cJ2NxTvysVCr/vhlF10WkKlQH8iSkSO6eT/JyradvIh
vfMNZ812G2wyKy9ylhakZSXOzqM6sS/w4Xq1dSyEP67qt+5a282iOVfqc5qHP3No
iF+ovlqlX+0Lo8aI6BI0Ll0Ayx5E/W7H5Y8p6Z3mKewkIJ3f15tAntC35cBvDoSW
VSVtBXf3IK5NeVhYKjayhgfdjmC6DgnAoRYxRdsAHNGMzMv4F633gZQw3/ePMKbk
Ra9WaHFSY6oem7tSvDg5B6ULM7ez2xO7rtKetcNrKak81+gZ+v7vn/lvGJQeq0hr
DuM0magXmFaBcyGFxGKgELB4xAAFvg5aVQFmHIwTUMIbBrD1vWqLUgxChTGN3w0b
1mmzGY6yVtIdE5aKkyKw5q6pIaCVE6yg1uRcDd7MNb+pkH5p0t5ih2+UUzs0g8DP
Ecv6+LnovlMkBNGsdZ3gzkHhr8Yuc42GSr9rAR3dCRdORTiGyFPOygSlY2ekmATc
0NZlpy6U6b+9gYAiD3zKWgijwfDXhsC/kLLv4Z/moJ/W5mC5ZjdrxtlNQjCx7Syg
O8j0o4Jw1se4HW4zmGIv4BX6/MAdQGzlvND6pT8f7SaPApY3bCWkjW/8VKt6/TqQ
pf2WHDkF/OiHS2pmlkFZm23HlCKwOpO420Ve7vJV4wZ2zNu0djpUBHOBE2OiJFhy
tyETtPUISMyp12Jiio4vUlcFZ2wJsgbxCRe8neaBl4Ou+lEU6mcHIpmHFvEFIvWm
0HPGivudF0SkFvN5VmXivzUDqj8mfomMzSHXU9pINSSnNoUgBby0oWslSaSfd4lY
AFwc8v7E66PQKJdKR/L7JqlDxI/lg81Z2I6nNgFzRpbPjCV32PLMJjWPcBEU6ORG
KjPmaMt4dhz5IL6akp9h7thtwnU+mWTrCxywNKxIsmkuKSGMjDPB8i60uJYwRHtI
Xi7A1DVw2mwMm05M/R7wyDi7aP4N/wO65Yy6Y0nalGPU2C7MQv1zFGcAAVCCmRyY
SSAJoeTbF4XJiuWPjbXwigZwghLlnWkWchRg/rrm9YEmOKunodMC4pRMTSSbKVjS
ZRbf0YHyZJ2JGIrMHyw+xHpBFN2/4VoTvP6JxwT2cRWZRc9atZlC8NG7dxWHLaHI
raREHz9Z0M3+rYTOzXjBOKbiNs0o2SeTVuazGb/9LE0ANS8vdDGfH20q8UIJwQUC
lEwqqstBifNbFw5hOJnuSVibK3Q/s5j6q1H/8Z28lks7Ki0jdepBKqi2owAlU0Mf
kYHxQVu1+3agkBC4ULpoKsbfgcECMRuFsSM+A8a8JP/IkCPKkBruksT31SGJgsXv
KkU7d7U0zi/jprQ/DUSdgXED7VJf9esTP5NbBRi+UY1i8dQbkxO/Dwxjaf27lWSN
I56br/d8Ud8noK6YQ9yUDd5DcQvlNSth7CkCxdyUExPFJxCSCDvA4lfIX9PvkPLj
lznE629MUv+SZ/ptg9xxy1XSMRqJBe6WWZvlixElnmQkvL8+MOi3v0kNhm9eXco/
seLTBe8iOtsu6jh6GP0eY/X+Dt8/GftX4IKsjMb5p28MpFmgXbL+Yyj2zlSncXAt
bhmAILDBJg3WqyIe1BpC2y1Ag8AdPWDYiB/cf7k2kCgeSBqt5bxu4fSitkuJR7tH
tWnQSxySDt42LhzwKI99HIQcs1oQRzQTmZFgEWumkRG6IjhmtC+/yqhwGzmeGTxO
toy20Ip9yLtMoySDL+ijLrNRwpygZiUK/wVMsw5MBK0P8cf782uCD6PTgX8XdoSj
HfIYiu6T8xLsjDwwnij3E0WF29FmR9BcVjBJpCc34G0gBObGCkNKtUyrxdY4S3uD
wdbCkK4XTDb0WUsWKj9jR44yx1Ab3ac1ptQ3xMRejfhh4lFjB/5i/c6dr2GKY9aQ
vutRjgofVUOykZvZho0ToMg6Hg0/wVQXJFayOER8kT0IAad2Mgpo4xiR7oFx5B3b
224JHkrOw3coBb/7s3wIRhLCx3Dxf/WQMCJSAuKNFiSTLuWUDnXrqAbMgPCZ4BAu
0t6qU1tUtkTESE+y/t/J48r2YpYTlvaqX3tVULXogFtfmqHHyX1iztGZw1ax8D7t
0lFXzT0OFqOuHAz8YMNRDd2zS87XzI2YjEeVZxhYbEPjd0RkWVZKJEcjrzAa95Sp
3XrmAPngHtp1isLT0Bzgh+A12orMSmseeCIJmEcqZKk1b4Og4WlSPDQ+ERhkNal9
ytcfr+7/vQVbpyEIwNJKS7trXRu8hGfj7kL0bwsSa7zozqMUR1AEEJt2QD7blEY2
/7q5CBdsXvp5HMgt/3UeM6047TiBazyCr0rX3om9N9gdRi+fyX7gCmDf/fIrEA/D
LIsUZQ3TYyV0jKXpwTa1iNuM84KVXoORNp2BDsrX4L5u2BpGA5/CNmyeHI1z7Wfz
3ly9Ctf1BlyDAg/pIybPh61oVj9dcYJ03UwAf2TEK8s+asSirIYPbfLZKE/rlIzh
JCftrXaRSOtCPJy/51XvBf7ci2HHIoZa3udT/PXP86JGsb8gJGoSIx6fRVlXTuf3
1IoBiKdvwmoDW56Exag/GvNIkcNvSv5B3haakHqhnnCpgwYiBGODJ77q3UM4/y4X
Z4YulPD0G0MwyAURRko1swriuje6lgLDua7uiehfS+nwglxWDSLPnttwwRCsx/gj
W3Fyy1mJEEZfY/b6qRla4DxJx4RtstVvnrFKafyuqsBKInMwTS8IGRKpsP0Oc8tB
w9V2GBHlRd9AiYoStf5xnfZ4VYoD9OJaVHRys9tuXztfLdwmfBq+EV8K/ONpGsl9
TJFTUlS3uEE74qA0LM9NeGPCmgPdksyj56jrC5aKuJwOlO4Jg+zf+DdvWm7ggtkH
inu7/N7U9H1u7/NoJLVqCMpGu1N7GNpRO0VpJ/d83ztCo/Gmt374XgAYQbsIOgFB
mUxOQZTpxQuSUnUFxbsq/EryrS/R1qCf1wN8es2ZvKk9UuT290G+Vb5JTBF7fG1y
PBN2EE/BBuUe+JqQVBkxXLLh73rv8lgL82EgNCYMI0dEMJEJzLCOQ0oHM29Gq/yZ
WRw3gQBJUMBFRPUVg5Lji28FKDrVlO3ZDgRiS3OwHPgxZnYa6pKeaRSbZVvikGyC
5tm041CsvozMfFYO1U1AMr0/YzKAmyYO3zSP7xLBNZU8MA/3DeKpiWPSmYp2yLKY
bMCPlI+NyFE4DUMC4by1LewYkh8jOppDNm0nZG9q4EYyJH4RxJJrfsF22M3S0Kvi
Kdb9+p6Hk84V/cGewEeDmLnrQjYf9NMx+9314XfPMkC9HCcwgN50hYhNGNWiATPJ
75bFfahuFr6ltxi2QlYOJrh0jeffwllbqPK3XDF4ZrHl+XnfraNDP//l5mMZD7t1
AmM9jO9RJVOaqBqNPwxHq2yV4yU9MslBSCO086RHsc+7NLkmIwfIDY1ErTQoH/+u
6mo6+g+dLUnN0v2Fc98hdh0L5iRgFfhGJ362rHxdddJZ5t1jYCAxMhy7LimrJe7e
lB9uCvJBRQZwXRNj2vQKbh9ZlEjLhUU2dsc1NFks6rUbKlcAC6WXDPZ/Bbj3uFeu
xhrrVNakNzqWM7IrBznNCxX9Z1rS7TJtocyrNUcoR8idcMQaza3lB2/5+8Nmawv5
3eNSGitXZftEjT4K30JlEGQCFFOd/98mixh1MOE/wFcFk/pqhG4FzFT8ADkreqSg
TdIJqK7R+fcKbJP4jWJCcpnVVCl8h/8QRf4Ff2j22O06xAv0kmsoWcZ2IslcgGba
Xqvx4HAfuY5bxmR3UPzKz9HmsRHqNH4kKdcjpA+syyxnBsxtiK321K0pcBHG4FaG
1coavpjIwCRV4zjcU4oqAt6Yn5a+fpTSG45yDA8ksL2X8CoyeTU+Pt2hy3jGeW9d
HOTeJHalZEkHZV+2H6QnlZSa7OtGgayjqJskyx+FKwSav43OY7kvcEssn+OscVWC
y2qcr5bZABhq6cTEsePM6C3koedzHikxh2VHkjIATE4KgUmJTcrwJGwv86U/joyX
J81y0HJagv405u+dAjrz7vKZYm52s0Z5yhF04jQ14MFMP0Ye+wyOfkiGF1D94QsO
loBpvcdNAug6RFw7KENt2bEDNPXmCEzzrWsLa/CW+FwjdncfGIJLRMAdC8Qb3E8P
MHM+Jx6A+JPQIiup1s3LYG91gdkUpMvH4N3gR+lm/kraPsEtGI2vme4QCHsCjk45
2OXbJWPJUxzgvszqNdKG31Vfk9N+06UaUvd3XxlV5T++8/PcXAas9Fm0eNt63ggc
LL9rtSleM3q8PiOv9+mXcxCsucWjjnSpS8DetwSZy7MJ9dhyuaMakvE9Fw7Jcg68
gJpPq0p1u7pDYzrsJgq13t0ib7q684CrH960LtDK0gAxceVSAosw7wd5g7OwNvMV
toBziQfFdVCfdWSwzCAXiX/e8V8R8AvHAvPN0qkALJ0Bmz/ngEuIKcniHLEuYVEN
tDF/vYm7cJq+Hnb1wiDEjHravW89ViI3ZXLGTY7/vkTA6/5E3sSm+vLJQFMJqt9D
NCz0arg9ufjmaJfxkO9WnXygmKMZNYuct5YLLfxzzshziIv6GAsjXuA5uplwL9jK
GWlJYReQYPedySHnthglSCa+rOf7Ug2cKzovGezFQ8i7Yf1qsoK5/o7tY4+mUgqt
//iSVOlYMCZpgl/Y+kbYPDyLLYjbx9Hd6I2FpCfcox7Fy9f95FRe8ILpAlKn8o+a
Jy7dTAAQABAZO0FLskQ6aTPYYGB1bOaDOfXWy0AWOWm2a2IyndgDRijiKpe9NxOV
piSm3LPTUGHrCB1jIdQiahooxaggfQDJ5hpiMUFAO0ezkR81Ihv3KDXLXPsa2FnS
p822CuztEqa5lajmPeaI59OsuhgVbxy2kUc+KOCPmzfwOPonMrQjXJ51J9UOK+Y/
uW6vukFiMgk8jtAx+k4aLPpEYd6Hn2LWocAdbPfAvF7nsT6IIiB22i7Vw6QlALqw
2TRplo4BQPNDrqZEOEcccXVOzcAkoGdh+gz04A94eund3/0IXfhYisOXZnv88EK8
jOqhLnexx1S/dejkC42b2DHPCHow/NGJXKA4ZqHijgkrj0Koyw6EVWw3RDpV+HGp
L8gGm+kYr+li4lS8OHdlD3gqrFXvZj2bAC6zBvoMDARUx+fL1MIxFq/VEA3mc6iT
/+9KLxzSsKOwavaB6RJpT3DvPfyAbkpB/jmwKh8zXq6XY/SxcAuH0YRck8S2Z8Zr
n7YM3n6+zQooRL7ethXo889B8vXvtpseWmc2VVGy5sFJ8RGVztLUpzMFv7RHLCBe
rjD9QXmyJsvIAttbziQOUWcrokhFQ9NanLrJxGKH2mINRB3+qJOE9EArUlVJWOwC
c8zoIxlIc6nhfk5EsbXtnB3fn+34tvFz5gNYAhHLzDk/U7hfVj8bDugaIKddOWYo
H1AGJm2l3UTt0/GDrDkqxALIpqFQqK9gc8Jt7U6RrL1YMM5OjEttJXCd+3orFAAe
dxNNDSDLfAiyFF4fcxDw0eI/5KMhGjGKL2GVHmXFuQzzIqytt1KzjS5l8dk8Yu6A
iRN9c1cmR9IGqoe5nfdji0xD97eFeX4z4C1SgoGCgvkd/FCg4hBzViBZSk8mUlUN
9hDWycnFUlDLQmSFfC+HSjaV3Q2WT7aRO9JWgnPcqufeQOxy15uDTYE40Gbb37J5
1vT0s0caxhCsRwxo2N3i0Y34nqPa1Z7FzcuuuabeUyOBYHGKx7X+oX80ka/L0MIo
l1S+RziCCk2psev9mPtsjfqroxK2qjugkwg+npuCy/VlE7ZGMnk5ks4pCqiVIchN
nkGyc700F6oQ/LnxirzeiYZ1c6J4+Oxo9Zl85euHTHh5L5EKrKnCuUcRYv7dzHr+
lYbMMgXhxGZJLKwXoT0bjN72JjnWdYrn3Cx6uSKfWP2XfgZkL/LIQhZSoHZYIF29
sVOlmm6/mmuH0RIGhwr92HB/JEvPXhyP6JVC2FzSX9AAUVpvvg7shb7ptgPZuT0P
1YqE0mC5C0ZrhW7iNXWylwsf4aFFbZZmyiZ8E3jRXwPKZtqs9aQ7cxhQGd9/r4fZ
LGsQzAa4DKV61gfvgwBNuJ0D51vPAFTpNFp46yoJakp652q9fbvgI3aXEXCkLyiT
nl+tvE6x8/bQJ6XvYdoA7F8/nKJPsK6tZv22zII7uCa+t2ibibEaKbE5G+6cISmf
aLIrYQo5dhx221PudK2ivm0wL2ZnsyetY+ktqtEgUyTgrJeGtCINxy3yUZ2Gs7R2
YkMjPr2wVSm3OLXu0XBaEjjr2LeaKd64ddeng02z1Rh5uaf7kEWPmOyRcY2wnA9P
qknvAShQoJjFz2OKHFgItCpQMiK6d9f4uJSyURhD2WUo47Bq9LR6LU0tPWORvfEg
pKX6GW4g7lSu5A7Ck0mYN+GLyBUgAYYI72Sl9qCg7LLEO2SVRgjj1szOMAGrx1E8
dxBH7LaDRqfQ4GtFaSoI+gmQ1eZHIqCSQv6ofzAx6bOE4nmK2FAmVQNhgf+U7MXP
AG4D2rIqG4BnwKInaMKh4Jt5U21tsmmCcvKXpZ78qzijvHacVWfjTcFmSSEv/Euf
HzgBFj0tJWBu0p/f02rHl+LZUktUuE4O1fyRWrGgMoTPngEODkyKlmr4knyKBgbS
QPIYfnUYAaFfwXGDLs+/+/uunCoOYT6+ft6MrYdJihljnFH7P85n7PWrCvZ2RCac
S5asbj0xTKHjKHPa6+Z+BX+qye01I1p1inEDPiQj10uIMbmWNyExOa4FppHMnd3+
4Nd17pDofGrPJbm8CzJlxdC8qT5P/atXS5oeo4wgybiRfTo0SS3MjHrooezlP8vz
ahyHtu6M4rcGxHogOQ/QwG1acEe0FamtXldjTJJUDo8uio8LeqR2anhre524nH9f
BZqX5IAD+s9snwT2h/DHTCQsbiMy5GIkD+U7SFGu5Dv2KnWa5636nXJakMAitaXr
YUYiggPTTLeUoK25yyEOy7HaS9Jg+3RVtEE7TX4i2kD2Cim5QJYTZ+1EWd+8vnkq
1zz/4sU+2Uv6rLpeaIik0nvYdpe8i0M3OvBql3rlWGvsV7FbxbvBrq2bsc3viEil
X0w4gpxnzxsK/ljRPbyVnl6SXNMRlgtfNfRWvXWC08VTMqkof7ZcKQQxzB6gIOvK
ZneZuYF5IX9Qo05fO+1VY/uS24kg738w02KTH3cTcwDbmvnCvbu99h9yVBCr7VLJ
On2ZPwNE8CDN4Xe/rx6cveKAvn3YhREtj75eB+XPhUSFq0n2ccAAYZqoZcgXO7Hx
ebDEGNuvWUxOTIU4IX8TgpjSRd8T1Fzu50pDHbWHZLewCJxCkPA4S2tO24bB/6WU
b6AfnTlGWFTsiIa6JBKBSHpb7A2Azt3Nr4h56aYy0P/hdYt1hMLnY3FgjGKQuY3n
83sMgnbeno4OLJgjHg4osGG7T7gljx01zynpysWZE7Hdqve+aU/s5RCX92AV733M
HMfOZCgMOmJ1ohQGJzNdLwWqXUmt72kyg0QfRghrrVtpjFbSdmEMvuN1T/3iYBhI
2JI8Lg5my1CvFav6ZAkqrPPrmJgRO6qBu0p4NKv69v+BtlOoyLeCsfE3UkTqU0Zb
LM8tsoJVAi3n82mOKU6VOB67YSLeR232mrQGlnPg+b3Qx6QHteMkJPjI/hj6ND5m
SvtinuQ8yWccCms1Pccg6qounBVnLbk0boOvxVzhXZaUUPJQiePPO5qkEAg1Yi6t
7lejkpTEBaJbHcEhRVRLLoHXnYSzxbfXcfnC8/Kh6Kp1NQ5dDmu3WsmZUrHzMUEV
6rVTyXsWXIhLB7oW3RWo27pcwCDTgKFUfMbgES64nMlK/mKJnKL4RbBhrelP+f52
DYbOvmbTkk9FelXVXmMgkx/eMnl3mjdEWcPJvyvWpVjtnRqxyAr2rX/WdULlnUhq
TmVI8s+zYSV0ZFksHCXNTS+iTvZkWVaRdVe1AKk2NierX+UUZnlYa+LBJ4fdkiqg
Wip0O5A/iiFdqCdu8CcwdEYR2f1bEV0P3cmKTsLRY2JWg7wOV2MBepMtUX0bLpNN
MHLy/ciD1qP87e2sFE1O4Z1Z9bPhp7X9ww9ZakZ230WNU60/JaRlshpwe3dzzLLT
8vwWfbFhK27kbHnZN9ujvWxnJgDwxBQ7/j5rP1TiMjXmWpclMwYejwuPsVKN/wKj
Vr2zCV0otxp1CDw7irn0ATHNTT3f1m3jbmaNeSie+9SaCGzU8RHm3fNknGXGZxDo
690NuozM5Yi3iRuwz8DaFwXECdDBC2x2N55f910bGgBxCzoPRgyDxF3rLFIJTfNY
1pUZQq4Djf+4ggvKObswBxMcDB7nqEN5e8WnFCroNrwNMUyBGSuGIn2Jf6ksp683
N81lkraEPXGHpsDDObqX41BXWOShqCH+ycqpwDJxbGiHfwYENRBsx80tUjNHXwY0
Lm5669XtsiM3BETTd5I4nWOo3Aa8un/CXQvwhQpTkzwc0eLKEfyEroOVLvs6qzpa
5nH6OopVeDBbDmY9WDprDA8Su8hvtaana9j7zqw1p9921GuqYlYYMCP5po/aHL0h
/jS671p02ye4G7lks5jYM5FSH0PAsHNdFWOeiPkTkLW4RazG0OuJ0QqRCbacLnQ0
l9Do7JtaNF8frcbhklzRHDgGPhZleCxddzUgcJ+VIP5fP+7b3Y/VjSXYTbCuTOZS
UDTQrjW2yINIzqJX6WbGBw73xh1RVpOhtiopBnaKXlDR+Weufazy01ifk0ipZ+Ic
74aYX4cBCGS3cHvDmsZzSwlt6rXEYCmMh0tuPdpp80gFI43LcopvPKpb2tswV78B
Q+4dAvbCx8c2iIr9b3ZYXEg+3Qj9oXNkfEiM4KhMxytWs5cOyEWEo/vcdN8Rby9F
1G+dpFzCDgq1ezF3QMt0t0prvdOfT6de51Kn5RvqqvGfs3mZvmVJZ/aAVNYrL+gS
tr+YUc9UbWSmNyMSNV46V9it8DQ1+YTMGQo+VZijA9+H0secAt3fJItj3TgpiVtS
zKWunc4dDZ577uImLVI4ZoXnevVbO6HhO5SLoYE154uyhRCd0YNtDHzY47KwIA22
u1IYrbb1lf7kyNODf14zZHWnMmIsZosDYQHZYWVZ7QNVUPUJaOgSWpGfDCLkr3ig
ZkCvhZJ3VNlvCk8PusJL2QCC5N3UABD/loDPitZD1JJxvVXBoFhcGxuhHHvZh79G
ampVoheuBQoeaeTbsVH2ZMuaEKiod9pBV7TPyknl3F3aWmQBIUmEXykcMgdvUVwU
uU2bkfwoN7+sfectO/SmMLw+q9pCl2IjbWP/D8qv8hGDfsibET0ATwg5V48sc8Bw
IDAEbgi6wfOOcWJ0X9p/MpiAjpKxmcY+kxnx0o6ekhWcsUYXRjAsGRK5oyx1y7lM
3UGIqnFWt9+zMjz7CvwqIb/5tjIKSqyMuUtWYx92N97GfwuFG9H9lkpPXr9O54Iq
u8V2/hGcBNJk1fBhM9MLuCQn/XdiDbLRgrZbkgxWZS4JmBCgjnD0HZBDc5VBJ1KK
+HzMay1KF/6F4EMIalxMlQJUi6cjE0/W1NB9ELSp/NGj1oV54H21jGwy9BM+Z/a3
HpQqmGXsLzngr1TMFHsShFzXPGubSmN+GcGD/V0NcX9/rxMM8mPoeLiORphC/RZ0
exw4hZe+KC0a7Wp9MNM+0we1yCYVxutxvq3Ib2IFniCfkTU+Veezej7iKnz2KhPM
ZM1n4BfMAAI6eFRkHQOXOU1k7i+V/GRtRRFcSh97wunmWxgry0xzybpDUU6XUked
7mvcJOR7bYumRcV1sBdv/tzH3U8jJbDw5sTCdltJ8W8O4Ev1j3kay0UcLlFS/rsR
4cXpEVMHy30nt14mmFZQ9OmsMeZ+Ptef00DiUEHbDwSdTecUPcT/JlfqTTxj9ort
O+a5uFKsK/PB/mrmPvprHfig+RHSaJlV2+/rfGSAV3ReMiFVqFfxVQf5UB3qoDr7
AMt4ECklHbcMBrs1QKU/cAQjN0VlAQbfGBiaMsYm8COwUb4Bvk8vXWDijwkC9yIZ
rgjggijR/7PNN9LFTAdSehRPVZKxuwVntNAsNkzMRagss54ElDVqtoBfUKW752Oa
XyJKMqBf4BC21I052p8r+9uQVoZDWTnWdZKwiPcXMJb8COJ4476fYbjxx/tuYmTz
EQW4TlEWC/Fvia9EOKjLVA5avuS9KwY/676wedJdELeVGF8JNdvfiQisBnHz2a6G
mXC4LzZYEp4Id/H4ods5zEZ3kTr6tm+S9ZLcNn+6jZfayYKvFyi1EvhBIJbAm+FU
vgM0+moVwJ1EpyjsG3iHO5IjJd7pmIqsG7chjjnE3bcoJEQKqAtfIOTI113TGfJl
MlDZIkN73QrIYIf5iepBr564iJ+4vMwuS2cZy+4XCbLb8kObykZc8DlGYquoFto/
zXnPEPT+RDz2b6lFZJkn+Qpl9RbcCTMM/nX+Xkxo6LlKJlbEdJYbLTp6WkqCmq7h
uKYUVfEHHvnAgs1gjQaZ1lcI9+y+iSNGTFpP6QsuLGXzxlf4Mofhnlw7W3bL/ves
GcmKhvs0JBmnI8DI2nTt2IlDZbqw4txGpVzb+Y5McaMwgy8Is0DKjzzr3oK+bs/M
4YhbVoEhPg7Q18ckH1FfjVPxBKd5cRBY7ZHdS2nFXjqiWLSsS8cnhnshJfawW0QM
a+skguqMF71lzA0OZNdbPOKQW+aWHL+XPxyz5JRloKjkz+vrHhd59/2xXqPrYyy/
R2ci5h5DRysvjLuWKBuo/P7TMasUhbV4sLv8pW/BtnlNZbRU0QkLgC3MsWP6V9Lz
j2Py6oawAvRdNOXlrO8Iu599UkEiuaOVvOI9kMudqXlyiYPd1vVjMSbt8TG1A686
5HsB7R4IJ5rvnCCqTR6PHKE5zj4CAq2mlwgD88jh5PaOmY2KzzurBSIPl5Y1ktRk
05kxLyl36gGy8rbUi46qQFnGZsS2AecONIsEkzjNboR9W+e71YQp8rNUlvBYzjkq
WZgFMNq5uSrdaTaCP4jO43t97zxEytG04qFN9k1efwS6b+GpehD/Gisc9kPAOnhB
e7l0LhWJWzqPPGOE0FEd//GtxRLUmLs6kmGvSBT9+tCMpOGvpDh12W0dFOkEI8vA
7o9K38eZHQ3/dLp1vLGqR5UED5Ys3cwhzLyA2QgycAhfkNQBxjcqpzdY5cOJihqv
pY8mEO2kpEjAvLzNtBw7jvh89j9zoYarIfOFQp0JPtI4BeAaDOE2qLqyyVnvr0j3
Uma0QOlDZFQQq6SxDbTlc8qWYN2bZIBIymqq82+0q0EWtf0SNFG39inNUCBDGTRn
V7estUrnPrz136pNkeHGDLE9sme2QIMJ0RQr/MLE2WMAWjmpFkI45b37PGAZYXXM
tPbWTtBHcZRHiWnp1gdcXG9G4XIhwfouDXMRczp9UbdbF9MXxdYBhKxU8BB1KJ7X
qu0xDbXFhv2tv1RXgWxYyiT8GIVdR08XydQZAF+VUfw2G/kRR5BSHqJmI//8nEjb
2fwDpnLTLsNPGw+xGFj91C/nUEAaaYt/EtfA0ROFd//40NQeibjgYkiIg0lWxLGm
6QfqV1EYy0/C72kqEUjqA5ELuLvT7gtJ/hwHGui8woOyqOuzHmyQnEee7MJYbdVZ
xvuUrgpspTKmFPphoM+x+elbSg0h9GkU2Z40roLYgKXMOPnAI8ndvWtzBL/dFpwR
GPoFh7epXiwDGLpQZK+4WDsidn3Io8UHSCQqF+GH6LDzj3aOrdMiH6ENRZY7tRKe
QsJI/YmoU/j/Uk3kXJz+rhn8fF+FwkpQtL3yU5ifRMjstT3ze8K4M6Vl6cZy8lNs
fnJ0wiJZBFk8CzWmX383uVUYt/LcFdQhfsElAuOZsGHupopkJfbnTpRdZtEpXMAw
YCiYs6UFRhRG569CkmUXxAnsGS4/5tkNwO8rY5wiMtBL9uAyejQSFY4I6Wthjkg0
q/KVm9F2PBzJzod5k7a4akBgiGZ9oHRWWJrGxgkGdaH2TVeKOBMlk92GuZrCsWeA
eFrbOYZeX6HSOfKSi77aemvK9ga4R1dfq0w58xPfH8kLRqTeem6yt++TkR8R0x1V
CJu4/7K57y9twR+u8b8PDXT0fGjdMg9pABcWKFbRMb3rOtR/gafeEonC0SUROAov
m+K5CMBLtfQvjr+RE7VvMp2epgDThYt1nqREA9Xr6q5HnIPQcOpBx2hs4xvMpFfv
uYaairFWaLADBHzfBHvgqphCt2wrP5P2FOBWnfqsvk3Ml/EqE270ILlkoZJZi2NY
QSs5oiG3FzwPnOubA5vupVLPxlmcxxct/cpVpXBPM4ltyKv4IWs1mWoxkcUlyOlL
mjQRGO4CFkBiYsmaO9ngfXOU7atne8di+W7bG706t59woqpnmDq1/+Xsr3tZ2ser
RlDVN76aSEVMPiXXR5hUcbpoBmN/dp6KPFIaBiQvQC6V6B6beZb5zXLKX3pJLGhc
v6FBCstwQZk9FZJjq32eot0fABTZLqoIjEf1zOPHyRKJ0bvJGoOQhywlq/tpEpSY
g8uVIII4PTFveD51Pjeay+b6j3D3ojYjE01RSP7BjQWOuG1lGZui+BrLJAEPxeRX
95eqsHHJQc76dWt8cfzj11fDK8U977PeYIn/+9mC9mayLG/gqT7P8KUN1stJ71sx
EOFs3H7GgDBMOY38S3EXIr2V7GXMAlyjQMAPfByHYLtYIBNmdxAYQ1kUfrZ6d5EU
RwA2BLNKefk+0n24Uh2BX3Gvb4M7gqZUmpZBAaPYgoXGMxkEdk+MI1NOSPo0JRQZ
llDGdSsO1xqY+9a8GABTqEOWxKdGbpTdqrHKiMiIQGC7Rx4atMq7V0c4HkXAU37M
hpaQQ2CEQfNR2He7clFsa3uEbCJRLe1SXui+wd4KsaO1gCxNBJOnFX9ZYQJfNskM
WgApQ66rqEwTdWjMQnEdkLRs4P0yDan9qpyNH514RU1U07yVpf54A8DXuJvK8Acs
PZxo13nc9SVP3daRNwKFQnocwppcubihgDyJILeRU5xcBDp26h7SIj7PYgrlkQ36
bhqrwnwO9xcXEBLsvTWJLbL4MP+mp0y6Ie1iJ3HJbA8x/040T4PRGYH/m30g7drX
0KFqUFOLx4WLmPUPHvTavxX/OTEoLjdCsR3O7/FR3vJTYB1d/OtbytcTO3n1iNHr
7NL1mESG6PcOI7RUndxqP7H3HQA+5BGwi2KLtP1b0UAEZH5U9FbYXhIV3l24hkQb
xFLODQL0BLRSe582pE48oc1WFFphRN9r5mpeMUy0FFsGm/X6BHmmZLffmRlylLcL
5jYmiR+jkuEes1bilwMSJXDPT8/F0QVM+rJYNh0I/Yg4TWMkIrFBIQlX5sDX/nP3
6A6olaVTnQQIX/U0rxzV0OXRDoNHqNc8nAoCP4NhfUKIZVfVpFzEjRXfT+e/FsVI
hwa9KOZ4AKhk+7pxhc3XHsZWhpmmuiTQYTmZHzdctgsoaX53fgb+F92ugj5I3SoQ
XnhAWXnfDkDLlsjcs+RwPFzUXNPIXaQ9bz87D7V4vUA4Y9WSHSvXV93BI8Kj0DHg
HheouZpqkMLTxzh/kVVFSD1b5Ua53hY/OLxVWGuJVJZzj5liZ9FThmI/gZZ4Iq0r
d0BibaxMYR+KFIpy/ruxYEBKzd3zLDzjbJvwalXSoPuQZKudWsg5WAcNexEW3Ofd
6ZE+JluNUhAhOkd7crMcvCfTNy28IpgCobqSbjO4HXTO6T0JYOYt2q6sIDoIJiSk
4Phi60vvARPB6uyHHE4AEc4BK9sXxPKzyLsdhuBqsY/UkcVyXglmIjuC3TgKRcrP
N4GxsFDs0JBAp4tYEBq1YwXxYu6lJDwk3qy+RYt8anMBYsVhrZNUnffbfk6iDFd5
vndWLr7VqnS9gdBg09/darlCjO/WHK6U9L/6k7rf8gVbq98dSJ+pAkXAukkaZhPw
gTQQvgA362MRAXtHF0s197k10+NTUSWzKwbmrLxy/vVPqc+mZqeevYMMkKEJreL/
r8X/A8Kqy+gWJppDdMRA7z94hWE0PeIT8PaRtpHh2OLkIhMH0thH5rW7eZv0zpB+
YYI7vAesQQxQDM2A9jYc25Gy0eSiEhUo9WlvWhZ3o1D0pOJNz/oxcc5faWqyODNq
lZyVEQwiyNQuMQFGJDSMGb0SChOxWNbvVdWV4669ph5YzkHKVhSB1amiwxOwtpDA
jBX45d/VOOv8vIpCrvOFc5M3zZi6jt8Dos5gMYzBK3l3VqaBRei8vfEMD3t2MFji
16OFV0FzbVrluCn8iFiWr3zeGH/exesdEkRN8jUdbIKDwGloDB7K3DzeDhT7Yddr
Vq5S/3Z12JR0U1nigro8N+UX9hIOJieDevwIuj0n9wyKtWvrafwRaTFfoTs0Rj9E
2BgicpAf6XxW6T4ZHB28LVjwXoDNwqQ3pydXVwIGeY++uXf5vd44WO0LzdzryV5m
SUfi3biIsUn8hP3xZ6YhI3qqcNZvqBYbTYy0I52y28gLFwp6C+pIwhmX7fmfKW53
NgoAsOfvz8wTFhzV7LzV9ix2802b2ZWTctzKvp+RrDrUlTbpizyCOp6V7kb/So6q
CScr1eXtYqQ98on7jXjBd3u9YhPu9iRZC89czauIwR3qajrPESGNj3b9zAFG2CvS
r9dyQnQHTt13oAVEM9M/dTS5M0kssExelt+s0nAcP7zxnwMOBgFvQh/2lcj8Zv6z
7/Ptmzj9/lbIBX3cavLQqvvX8ikg7q1sUuTEdMQSEb4HDsunVwWqwnO4tARlQy+r
g7eIyUhZ/7m/+gAEvsJg/j2HOoRfReXKe+oWRWBNYYwEOBWZS7u1OP0OSrMNtBhn
lHGraQwo37p5mM8J+WjYS0uqdo39igDSMiIdKRUbp76dIu8tTt74WfpyE6wEajGD
14oBn7GNaVuOOB9JgX8KHp3EEI8s/herKAMRUK5A8BKT9E6ngA365Zn9F3j5mNDI
4/GeOO/X7OkNj1ZR19ly6/55tL3F3LnocPTZLpjSlsRb9mj3aJ4F88k1lRg7uPPp
v/Sn3FLkWFY8vjsHp7gUn6e7GbegSNdBRKRoHvH0X5qLTmCnfnG8AIGjyLNgYV8u
NeJcpL+AfrF+SLgVoeHjtKP/JONkqsYhne3GtnAwpJIKhPWvLEMo1SC3kcodZZ0A
DgyYS+BUlskAzZyrIuHxwpZfJpKDBKRnnLnJX9om9a71Se4zgQbduPI8RhKoYXNf
jF7i36nO3CbFc6Zz2BddQRML82fskUHaQGAmuDggImOsoSRq3yd/dvCvTHn6wbpg
VaOKEM9GkJG4LTDdGRamkCw2qKEsb1L8KGWJM1Cc1iDidad1z4XeWEpj/qPeysOZ
6/z8OneiPqNxI3yda2zVrPEPia8ZIBqXzgIFLzz58zzd1u/j4/wlFEOH0P0TBKtV
GW3x3WaVJgIUE1ubNovtcsuMT2JyqD+PKDB30UI/ZjUSSeuohBPyUftuOxBeX3Fx
Sgxvoa7OdTLNNRl0JVZ4ISui8c7auRmp1wrxWgTrFV58/J4chTqGqt9yL14NZRK9
Sl/CHwO2yB2QHfQsZ+NAXcxdOMuhArh2wLgHzG799zr7BoIFoLdiQxuROpPvafnj
Yn7LV0sal3ak89OX9D36H2/rgRRi03BFUoCJ7VRWESV7XBPV1d6lbsJmzP7Z0tfC
xKPy2o3KK9mWDfppH1zQTkvknDoRGg2+hP2xG8P2tbOXL+WTIoPDB7iw4E2HzBHO
sZiyGFtfKZLYWjHaTNhkETiYQoeVL77xjQbJHclIaahPu6qx8sH20i2b/5CHXJJK
97uybz2hXmkyWMfJHkJK8qgM36764cSLnLhavG7fXC1BtvCMrL3Ma20HalsYUPDk
/uDRi2ywNGl7RL64L8oG/BWh2X3/hnVXU9OEkO2dlYK+cRiDrdqYYrr9F+K2bd0q
XI7U9M8mqM9u6Pf6lqaha3PzNN8mMylUP7ZgHVWjuAjdPR6KP512VzDXcqj0F5Ho
eDByWzjFlm/Qfyb0f1AXWA5N3mngK4RRKCeDKUHif37244Ry0FVXO1CkgSu4avwe
h/C1UmAmnd9jq26rAowyaKQpuDJLOuEN3RvAYWEMBmHyk3iBULpBMoRngn5sKpVo
QA1aLRdnV7oQkrNZzjFxOpH+pY0j3Ql1ejRCTZ9i4N7blBNbT+Yk9CkBPhd0uTQi
3RmPyGUR2lsawTQlSLrqlMTQiH8wJzdkjB0X2scZW8UsnkdDvBtQxBI4SQo7OwPt
balNGAkqWhxgaXXM+DwdmYmbYVTQd1K0UvK1CfjysMkTmYHFcrGXaizmMT45q6gD
dVw2yQPL9+D8j3uORVStJvGzn8kOUNTafJO5f0D0s9Jw/b672NZsrdpeCgZxFJaO
Ynx+OQlwQZ01kon794ElJ6srOEoYIMnlW9EnpuHuunylh/ZCEki3SCOQY6MlP/vb
L/P9l3uD84xp13SdW/SiR+TWc3kTWu2XbzEOC0SsWYFtFKrNDs4QGgDE+RBMsQg1
fGMks4zvhbGlqEX2pFmySMLHTyx1whCfog+JbulMM5j0QpHcHJTW/NhouP4l4Z8m
BgQhCFY2UrolrTZXaYc2tKYeJyevI5xmMJcC2jUUZHl7vpaqAuKsw7unyaWjzLED
IV1mEeU+hil2pxQqaj0KPrwhOp4/wTSSYZ6IHpzt0KyW6JtkahfEW0mVAJ03XnnJ
DZCJ5BnAOJ1a8xwbWKpUYVG/TwifH7mWlR3FjluYZ5MIHUXzJXFBugRjNjlKzsRo
GrbXX7yMA27lE3gT5eG53WDnQVZP7GXlLEwpHnVmU6WFctKV4n5sS2EqvAdohb0B
bgrEcJ8jdwCk8Lbo1soPo5qtauMazutHXZqwr6IrgGceaHN3tRL1Sx2xJZW+Tq5a
9HkeSZrB5UCBELwr5Hk/MJ7pOjsi+5nqE+wIhRYGMacAn40aBVwKyQxih152MU2e
QYv6vISnJCRlbxYz/wv27MiCMRj7nzxaiyupgJBPM4AR8MlG491fIqckabSEK+VP
nc6+k2NPQW412MHlIfihecrYuySRwFqYW0XlN4AMC5xEjGyaghruxjZSkeRgnDUQ
pH1zrO+sAMGOftKtCbrJV/YMwhh+f1P25BFD6Gp+/000Knr1Flj+14AcsCg3Su/J
WNAL6pL1+basgSXzJW7O5lgylTunxE6f8P/Ku1audA9bpAtHx/fi1oCeiFWlghTd
fVjO28jywbpC60ba3BXrIyoMf7+yQTxjYuyc3jz7/wQT3Ux0El1R0BWHSEL2uQgi
UuMXJ9+bJj+6GT2q5ATYrUy/kHA8VtLez4cvPkf+EAjAEOitVzbIm5DaifKO/FxT
Yj14PjzUib6txN7b54tZDCVQR3jX2DyMxEetI39+zpfo8F6d6GEBkT+r9fhX+7rJ
Y3VbJln3k1GIWKqtbBDfdjikIHtRGdrZ2X8HqKPc6+tB5RFPgNi4ZRpfk7et8zw+
y6tF+Y9RD9j3aLHbJaTv+Rp5FSEhV47jnXH3GTJULE63lkmA3bLRNqawqeE/gNQ0
trf4CONygccvFBgCEdeZuq8evekmiLrGVHZRst1v2bmyNfvZUeHHlzUxln1LVtfM
Ap1lad0lEkGmfIPWmoZkLof71S02WlheYKU1KWojjzgSd4bzb2J+bz5S0ED1p1BH
CdDuhulSpCF9dkrs0emfxAuJSFMuNnStFNNmAWFQEdE1aN+R15nyrfMTUbleN/Q/
m/M5AaxAtmgCZP6VL82cYoBP1J/vvH3PagCC5zZ4BIkiZ+qKshfIS/vyNqUE5dZl
zLIPGnbYfFGg6KUo7mG2HwAjFGGsfue/gEFRkqXSzdyyQ8lTaQfP2cA7WKPP6f6t
zJSORHbNBy4NYy02JGWHWgInGLx1c42HtyYys5eP/rR4cJ0qMry1GbherSPXtimN
myaJZp/JhFpkpbYHtZ+H14CE6KRh87tkB40kroc8MMCSJUJz/GcJdEGRr58teV/I
RIdYdh1iVmliyTyfXP/fEA8XcGnmd2L9qj4zUL4H8WwvzD6PdBnqShN53RbHWD65
nIIVRW79IZ3EIifV5kk6FGHPrzkvlPZL0VJtsi6+FGOPDHTTs63JbORU3E3G5iJ9
GxjDbUAgNMowHUOZu6toMQKgaJmSU4htymqNnef4VqBPbd4OWa+5MINyRcFjcron
wLM8c6yvWz6WuzkzD9rEf8HU3g1bjtz4VlF8uHf4KuR4ROEwbqZxpfsCVKkEfGDm
nYfRqbRiqvba4KXDZdW2UF+INlcax32lCxVLU2lUpNau1gLqQoEmJQBLgX3rOxT2
iXYg8+3Lo4YXLxyGsHyijleoZWgeW0Fj14WgioaYvNNJegxMgdmkhw0Eaa+vdIsf
eB3oblv2OC9+/Fa9jssvwHmIhYUk/yBRNRFGZiQeZZNjWkHxsDmCPU0zN4F/I+X/
u+LdCcZe/5S7YhMdZGs3zPCc9g//aHKcUbKQmP35qagw9qSJQZN4qPB/bdieD3xH
2L3+qES+JLF+iY7BSqiB3W4hKqkSFoFcfkgdgKlr3oGs31ILRUwEtEEmXT05oMr2
keerl5U0RPaAI5Bs437M0fmJtaAct8Wk4jzX5SxRtxhLg5s7IT0F9tZFksMH3PEW
1x1vbaqupL1TLpH5r/rhNY8vIOzbozYgDCEsGolwpkojYbZsYzEXIKmakwFY4tPC
viaNNQn6luZXqClljOheWj0tepQdrwTvrWZ3wzm5vYc9qBHZIXf1SkjVPRHzGA/4
+m2HEt27w1AGQx/Q9MFSjGrxoU+MlqZoeSFDbYLnk1BlYRjImA32EQJnu4xnhJU2
hb6uu/1FMuzhH4CSodLO45lIr7qENHx6b7dw1rn8bvVjhHc0TFeS5PhsbriTosAB
Hl3Pfkn9PzkqCtT6MmgqSBnhMeEk3dILdIE3hSiKg38yiJaXP+jIKWUiaT+AYetD
9dC7uKx0HDDwSsNV1eO2aS4v4q+kl2+igX1hNwVnUwDfs5fDsX+dNfAlt16RnLHI
E8TRCmw4VHDf85balKjRbZOKcWxjLohHLXkRN8SevxzDpk1+EIx7C6SdyrPI6Pc2
lU/GsjJbxgi5MkaxKOLa1Tdy20sTq4OFUcfozmwcq3PlKg04S/ynsuo+YMxPtmo/
k0sE1wVcgDuvLLQ8WRcB0KL4MIFa+tWly2hyFGKtv+m/f5tmyzQcSCjyNx/DENIb
tatD/aAzqasVVbS+E57sxBK/SIMbc4wqtwRjSs/Bm210V4ZRtnxrzmbQDbnmjwh3
5VenW3WDS8eqi6D+5sDXH6E8ksJ8qVD3oxMLg+G2upoTChGQ8ZuIl55JGy8T7ndl
kjMrCStroyARSpBB/hbMTivyHeN2YnCnVNu7PmoOUedTxJOWm3DD0yvyxIr5AICs
bNNbjog7D7s/MU3DZL/9k75xRHTDNhYPRKtQheNyS7C6ftb/FRqTxOIBrq7R9kIf
wIyDmLGPPjKonjcKLnI4vf32daj/QtawZ5n2fPa3g8KKRUZojaL5dEq4TLCAedwR
TPRwHsGY4i/q+1GW/yU5tBkk8RStzdNGg7Fdx37yw5oJ86eeY6vq1ZfTuHSfeAd+
AIgVnbo9V7DUdil96KuYNUxuXzDdBDZCtl3me20BGXTjZ/dn4iBM5Ly0q8USSq7G
Jd85gpleHFxt1cDM2CTKlz+dpen7seLqmwtYjKPNwSOzZx/XLmwUPy0vxL1EHKJG
9ba8QXMnmXZauiVyNF84yTvXSQftgtxIerg6kPu5hBfb8ywmEO7qpFvQjimMc+Ib
BQpnG6I5FsdInfBnqTU3fxkAigXjteruA1n8M/wBqx9D9rPa/iWITg2ynflO8czX
sQpMwwb24WN0k8FZMSaUDxnTrtkKTR8hS9XNWrA2WTGYcKhvBxtAyqV++jejLbMb
rqW4hrmY1MI8sVSdulmyPxVYvsX4Zdnfm945NGnjL103Ma7qUhdvtgfVLEmUmxRc
kJrku955YOKJB7rtnoRll1pU2LaSuTko1o170bDQ4ml0nEbG5a/bnfKBRWeP+ork
Aq1UyFQrUWSpz4do9+f4MvtkvkDUJq3Mp+If4Q40/Y5+WA/OS4OJJ+RPmbocpnkG
SksNxetF3RL3GgvWkaGkbzidsGSUWlGcZy5GcpdzTfe3HQdC+q9Gq7keNjdx8Ola
+Pz3SAxGcOSOnsMWaqewetWbq//V4tWLD3aU4OrD2ACfaY6mlnGq6xbNwg/qSStU
mX1WQpm9pMCcJHhn8MlHAuBkDHKxLRVYBZy/vGa+J/BeoGtsCtjKWwdCxy9KwGD/
IbFbpt/V7zypuJvLIJQgaEHv0+ZN1jv4Q4KnJDFgs67flsXvFVxd8tBwx0X+vtpE
R4GeSy8qjIGNdgYucr5JDMVgAqVOY5bbtodDG748EiX9IQ7ljZ7D384p3Ki+sIvx
gnN+p20+R3fKL0gHrsWMkJB2mEH+IGQPOHY0mChMaLo62F4svHJCOS4fE9dM1OFA
nqAm4LaQdApoFMhnwd83LPrldLXHTSV6MKeD47CEnd/yyp/IYVM7bPbE7kGWmuXm
4q64qQ/NC9sSKfrvxSqMRO7NA8Bz77b14OTBQUsNwGAedERxsA69ijq8LrFv0tPy
j7TPH/NIoFbaCpmp5hbuGGfeipnSyPwpvu0AuOTNrfnuVdCGDbct3mhIKpzlqVjH
fRfdp59OM8p2oNfkSe1huI3VKYDAu+2+PBtaYUpl7hlact/lVpqtH1Oto2Cl4dXu
CU6lw6hp+2ZlKOF6PCC3ppMpTbVy8HidAPgzAO46LqoBzCTCagINVNJeVjOJbHPk
LfrJz2l+Ue/zrEg37vc4+UUcWgz5L986iWFPfHdKTFu3kMncwJSldXnu4RcUHUIV
nqvUHhyjVZ7qjAsji05+BXW1fLNuGwFwehUoVpM8nhrjdDD8puFPENSK1TweQ9hk
8kNFGq6A/GZgfr22zp6VLyVd83iErHoSBsuX3qRu+knLJpJCZOhglbxxDMwVpQer
1ir0YSilk7PxMYhvhEjDv4G8gVrVB5yXCd/Vwon2NTKNAqqGSwmHDshfp8C0TgPh
eP4d3/W1JOAplWqGcrppVmyo+L3nWqzYj4iVbp0KZlyj9FwrnBob2MSGiaY3H9Bl
LwfO71Qj/uuNaL+N955yrYxG/BIPLZU/RhZP/ttklWVur9S6IjBxyhW/qL2t2VYN
a6Xo6J8NMqL7YpHN0mmGkZjHrAIuuFIHsHhYJNfUv5NDju+eGtqCzbAEgCrdGrfr
Yi7GUyPu/wuoCYT8LKsvtmZi7lMoXws2hkVJmbOVQg8i+SQPtgseRvvLNcFQRnc0
2NIl1tXhbiAIuShCg0nudkE996VUL0AITh5OLDktm1rueMZ8CMw4StsRMQZDMvyf
st9cxVcvKOhRDX0cy/uVhnCZbAV9AyfenxGOXltfriHVEoBDKu7wQzudAT0jDyc2
tiL+7qY4cK7jaXgOYgTzwOTP1hr1v3aNkul90NTNYxBcLykD7H0EC/ZHsMzzUChp
pHP8D+KdNgmIWwN2T7Angi/JxE6bIet/wabwg7k9gCCRN7KSW6JAZiYvCs91SlUJ
dSmav5XU2ToVNmpz3mcs3Z+LcA1JcHLBOqHyAMKBQ5HOduN9GMKr6XqHV1cFbpCR
MN4pglvdZtWwbh3bJqbIYj0C2+GzT9LeIZHb+zVHcoUbhJSadw8wcuVG8hv0Obyn
+CrF4vkOrdefMSvFLxYDwmG1/ftj9v9xs2cAezPlXYEmhsdXxTYzKG1oDAVrOh95
WDf//+pCbonZn+nAV5k1CcCU/BxGpb2R3OnrC0Pjq8S7M7EyHR0OBT+GsfUrcWqj
grrc+sslnQB9j+Csu4u5f9DLoqXOXcSmmcCmDipJBNjJE0oYbTgIz38V/I5yjpss
XH65oTvDlhJuUjeucEQSbXoH6sXhSKXUzVp/VPphTLcX58Bq0fCzPzivDcMQ1M1L
KdzWWJzM6XYLjKDGzfQJuxpIY8aApvrbWr9Io+dcq/YhMpLE8ekbDqC0kZpFTbHw
79aAmUW50khaqKyACBD+s1N1fKVG/9W9Ri/AV2D+Z4p0BD8poDJVaPfrSHtILWMw
np2F8IXgl8hq6XOqReM+kRV+clHkeGk6ntCWTnmVhS/xnXOOAJN6eVXAgRURqHrQ
t2YKDHp9+cc2NOomVIlJn9nV4UmyL/kuD/EPCwo49U364YZG25VwZ30SoGNvfuXC
GDD7Fq5ptBEGZfbZGAtf2bTKhLoVKqjfEe5A2tAPc0LAW53pcYb0Qww0uqwpgMdV
nFn3NUU1GVAtKMnENG4Pz20WKV4hdLM7Rbtf9K/pI8O+VxJ044FaxvKa2wOc6U+R
SinZUiJXFk8ppASLjLoRMKeQNYM1th2FURQKHJho2GTVUVAQQu0McRbqYkcTAUX3
Gf3E4Pp34n1MuNQqUDkQPhZMP/8JwJFZ4NgEQkCYv7dpGJBjni6sw4Zl3Vb5nm2a
W0iw4zHm4xWB2G49c2mpmfEcXlkQt2ChJg5Nt1QMW7hzCdRuFjhjbL6N48ZkaAM/
SYIkbpos7xfxjtJLOn6CgCq+tB1fpv5jP2cUugNBcAqqNd9jm/nQ2D+ALzcf9Ya0
XD+selv5/PF/wzzUDgtePYQBz9cnzcByNZTj5kLxRoo/NtMLclQlSsQ0mqGeAzbh
PuSqvP0EOP30nlv68jFZNp6NukyoqC1NL5f6FeWYZLe038uqbVMJZ3AmC9rhBqo6
CXRx4XlMDbDIgYPdNUje5jPQH+n6rzvXVaa6+xGS2vb7hLQAtIlJseRvJjJ1d5jk
pYdZkTCcRER8teuWhvQBnl3cs1QvyaEXaGnVQkAqIfuIH1V2XPoetj/9pnuEtkNq
hKk9VrND43XzfcxI5ZiG5iTj58qO2L9MW+l2qUZlozVFOMhbCdQCp+AkOPEyezmT
30c2xxTa38OToESRHkVsr7m7D/0UtFSVJyPRnijEFFPYCRQDAmGQbKCPB1Ytdkm4
l38Noj0GPKd1RTAfBOHIbyWLnvjLwC/I3qs9FiMqDKbwyNaJYGvMQPRTwi6hTGER
ZVQKIsgDQxaP8cD9T8GiojaZiKg6hVpv1R2abEeACLO/rlm/SWMl7cT97r3RyVgF
LESMaRZZdd0STia/mGyAOhsbcKJEYdanY5VDE1z2YhY6N830iFvTKQwYR7raKvaH
TnWrx9DicnXtPnHLT6eNrIp/c+m2/7KGp5rBmyrh6YXH3RpRno/lTK03FwodgToq
h79pJieTkmMbpC9SUrcBoKfV195EOyxlgvhQAQ/ZR8f1NxJkjvFHX7OC5YR35/5w
GBvhaMxV1oDb1s0N480CrztrZPtpPp42d+aCGu4cn5ko/jUfPKNSqcbm9Czc/EGS
8iGNXvWivAgclDy59oV8T7HzxInTyYmmZ02t/3ORASqPi4b+MfmR10T5WnKb/MZK
/zaf+mn1sadPvQsY8WeM3GINm9s/Cl3ZkfeuPfXmjpl5zUyLMg/z6tAQszubQpdf
K5jsKEodpcptoArG/1ItkTpVxfszjJpbNAgS22wIM6O++YTDbwNxoRXizCk6Ntzp
gpcr/NTIuCrOfmhovbS+3pRBKTBkOzLmV3mo5MF29xv49Z0x4hQ3VS+IZ66fGMFc
GC58XioNJlqMkTZLzELWnx78MyUIr15lzYegjRsXZGjJbna80VXzMQf0oOihS9WJ
pBX0PGxGSXxCg+gz0RUA5ubX/5NzQEn3RX+qw30lc2zx/8IaQaecgXZ5byzPQuj4
gwoXz88Unr1R/Ol3s2RBpsxPk+x5ZeMH32tzW1SiFWzlAaTRSF63vNmtl1A30hne
oiYCwn59bH3PHvVd7ZjqBD7EwkaugVvXUCeTsJiP8wUlHGkoainswq108kkGGLj4
R1jeQvetObBKmCdhNVd38pooEM1vSq7syEJMt2InjDtAAwLSGyM1VydnGA5jocNz
D577vYcg7FEZJdO+CfePz/MQGcACj9TRNvBcg2UQbjKzHgaP8N9QfD09V6Nc0hUp
2lnqqzr6Xt2yUP2C9Oq8Ar6Lh3HECQpmgiGHPaHrVu41s1utasNSwbfMJ8UddmOT
7j8E55FyIrjOPOrqk4coChLhHDDIpslEB5jr0RKGE+uWgPHX3d1hYVqa+OFeh87E
SSgBRYvEzQariMw/eAzYpOUP26mtcc9OKX1SIz3w5diJn+MAEC5yFyx1Uogm3OoW
ODTCtH2hVHUKo+E3ZN1tWj79/wrF6gjutlQPxm5QDRQhFmmvmj0MbcFtfMiuWmfO
vn5UYoObdzduVNPdfKKfZO5DoB67sLmKGFnO39pr7uQqC+vEi9ybu7gqEwFLue3l
HFrS6hTm5CjllT2aD0T46F6c6wXAl2pYMVdtDsNZuyftmIqLGOfCRVAHIIFARAly
vR3RmsHlaNvHTYldiK0BfwSXm1/lAg0tveAG3d/pKS4PnqHYXOxZsIc8CTeEd52Z
FBHTYnQrJZBY9wYBV9TOGOjVPvS3GznwdfFHCTjwFW05+tZGMiGmIHnSxhz8ksr+
M6KVwTzXH0UZXc+qU7IK8fDrbLFeZJnP//rFXVtAG7+oSoyk5GDCkh/3k82/FyuE
65IqUbXi2Rvda22jWS9Lug8mvh8zWulsfJSgNCu1sgkjT7Q9mDiMjWSeO4Y84xms
hFrhu3y0EjKEdzXjbTs1OmRx5ayQCbjLYh3yTzewjloKb1Rqd2y1MVuHhpT1mBoS
M6vM0SWQtJHULKAu8poJ0QurlO3ikzeFimZ2XHwEx8fPAXnKmzSJIGe8OQY/3Yv0
ckT4lSDI0tnaqP6tIiXYmiLmvUoMySB/bRA8ZNbE9K825s6UjD+8Vx32wcsQhBI7
x1yfSvxsQYbfd4h+8XNeMiZvz5EX9TcC8zvTvODolfcMadhE2ZbjjvXEhp76+gPU
GW8l5W4EaP5BTiH/2tAZteBRqo52lZAuh9G1WQaKzwoEGcLXK5SZm/EE2rcnPZEY
dZZsgZwJ0pxUsaBQlebL+xRFi74uRTYjX/xgc7Eu0+jdut4e7WUd/BXOfVwvqive
3i6BQ28iZA2MdY+QjvgM2r1pN2X4mvWXJ/wYAKUqi72xWF4BmQa6WAnk6oTPr96j
AFWea6Fvhnr7vYubaf5PNMDWCdVcuuAB3/rG/h/sOj4xF5kDRFMxQtm29E0PbXA0
KzcI+IuZ5T6exSQWofQcrSASZiJLgKjWffZmM0te0bUpJmJgYuDkSB60bMlCssim
UjG9i8AiYPFq+uSc4IklNfZCCydphjUumYtNIUk6KJ0K5DZuC77NIrM4ojbrRccL
fom6FHCyhG89qQRU4yLkIcTkD29nN2qXwVUOdj3KwwCpGj7wrCg5FlAC7AK9qgEi
EdVWvGhZnBsuZNs3vgCPMp5bUTLmH+xeFPPSh2sqKUPk7geLvyPz0WJsLfS5tT1I
t+jfWTIwREZzI6wrRyYOkCoW53t6JnPGUWBGtNfF5R5tAtkWtTG4HMIBAQG4Uv49
RynD+adXax7Fa1NpEsQPIg+I8oToCgUpHvJg6nz3bDXy/3VqzLPKRAOXBmYCF3vG
QjaqFNbI5CegG1cZ3qJbeOrAUWqGt1bsz6BsLqenFL6zjoZtA0in7e0FtEKkueG2
PHtktmTL8jAArPznd6H/sAuxCCo9yIRq0ZpRLrs4hHHS+Fcc0NVaT7GOSH1CCfqC
UoVn6QGrf15HDJPiKGIv3czWbj6DsQGXXFZ+arc3Y61txIslNoPeRcts8BxC9GzW
rkHhB908ZXx5ZhnzxnN7BWcMInrWiBJ459/wVAiMSZ4MwrOxcRkjnF/eqrZUilI9
bi752FmGD88OEbm/yCYmVNXD3HQV8UsiYTbVL9FL7ZSs0RvwsIFoNaHqxOgCFuLb
FSOCuDebzjKN3dGX8dIElhXcHpSvHuV2Md/YxYKPRZ57OO177WKqAb6P9jDp45r8
oCrwgt9MZH7fpVjvuZrndcMW/cf47ajCFkuK5wGNjc0L8u8CDwmYJu3lP8rXT0oR
E6HSNxuaymJxSXE1LPrEAV/vKf1QbXOC0xFCZs+j9wko1KBHBeDMpwXbQxyBWRIC
Q1RwlTegzrRO+38fixeVK8jWFw2TWCL1FFkI+swrYZv83HtPTnlkq3felt1nJlDM
4G54do0UmWeobZmGfY1a9vnJcXwXUXavGgrmnMMfL+IE8J/0yEennY0mSuegN3ad
8M8fgU5hWaBqGcQt/nWzOc6Bkfh8HEW7uGAY0fvoDrNsogZMC0mcsSIXahQIYwqS
EY2QeOkTykJdxWXC3XT9OH3uMQJGolR8dZYaGK1x7MQu9W+SOxo8ucZuIJuXYn9t
0gAPtamOHJLk+Ie4KgGI3l16ALaytWq+3XPERCqpADKar6L53GdUxXRmQmtnNVGl
92WCuqnEYkkw5zZL+sr/okglV/ZiKbpJ9FQ1kIOv56vPeLnlY7tLoD/MpbGVsS/3
zUL+u3W4eTT3hWbG/yJiIf13TxoHndcezLxYMz4feY5YJ0TX/j8rEoGseRL5JSK4
Wm84M4F/DewYSlYsDkmnBWXwjZlmb7YME49ml0ceEyV8zvsRYcP2DiT/AONjgMH8
EYimLQrXCtfiti8ab+8vBniRExdyi0QpU/ppDNgIqZWwxzHpeQGxGuyikbAgzv7S
IO4IrVfvDSXRRQvXLE3OWPIhaCdNgOHJ3KOQRSs4gBej6t+Vli599pv1FSOsVSVj
iylv+modNbxskP04kRerU5/iYrIKgQMKR1QDx59cedZ8JJ01zgoQrnNnyo01IfDM
02h7IcrVIopkr29MncJoRsIc4gLCiv1rJ9dCylUv3Ix2ZROOGVdH6J4uTHk4xo2V
9TYPjHN2iSDDEAr9ztWDdXqdpXeqz2aJbcDyN6JR1Goys0wN5QpvWQNThxMWyywH
3Prp7OLf7aON8lo03mhOVuwizd5IcpFFqr7UG9tuSzrSPO+wIfkz6D4gF95XxdZ6
o86tcKy0JPE7WaHyOLgk0xY/0HhFD12FA9DeRLFS89Coh3l8EkEkVYNPaCO3IQSk
G29GcqLoc/yt/O+dDLkqGUkR7GR/5cEHIghjG4MXq4NcNc4kfTfDiYiTQ9bGyMJk
96NFHnZRKn30l5suoEbFkhdD/fuSOwQORZHSf3iH4bKEpzY97V/dQZPi7R7Yn8b4
50RjcywdfuvfcYZ15qYnnZki7H1PN7rOrISLH3k0863UHiLs062Nmc47gKpSnr3U
tE7d44lP55oh/SrfHklt0h0+uvJR+VFJvDP6eUWs2Uroiw3WItQD+V+VfoawcJln
PJw18x9Cr0iMcmC3sd40S8uf64V9yxOcntDefeYqfImvUI1Hq81V4TSFybBuT1bH
lafkvqXQJm0uakMZMlSu+CgZeJPtsKLNZEH2X6MjAvYykA0Lkncwsu60OuSJzwf1
VXskaUjZZBBA27DRzalBvJPEBpVUzt64CWWdq63YSxCaigFIZ2advL1W2ymqM+NI
GEd4oVp7NVTGeejpRfRLf6ZvmmxVgOa4oL0HvBsTbftd2W10exdLjPzIcb2SRGzr
SX3ES5HPhgccHkKdkkDvhcSVLm3hBVKlfg8+PYrryL/bEbSEh85awgSu1IS/ni8t
cNsk1Tz6DuIL1CUuRlvcw8hE57FCWd1iA28Vmbr94XLYm6kssZ24Eb9JcPJ22yVr
`protect end_protected