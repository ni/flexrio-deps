`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4064 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpCQkVRCAeB6CX9jncQXLSuAEg33b6Fu5EJ/uOrpq0+Jw
6qso+oSBhkUJQrPAl5O8PIbPAW9C8o5LWrizlMEKt9P5NsA/pmgcbcjRlyVXsIdV
3khW6kr8CmYVecnYACccx4/nmTv3pkkx0Ah+u4rtNzPYzrCHHx9rEKlY83I7nfIF
6SzWZCmddPQFZWD7Mm5MlCA9ztf26YmWYv38+G30IkJje2+h+QivvQ6J794331AV
04V7FheYEsWWQ1LExNYeendI3jFJnRSkGR2u9fFr4CLzshuDy4i9YLstcaDh0Vs7
3MFnT9ywNcsdQIwcZi+3cuV1Z32GhJPbcL5UvvLm2kj1s2WHYIZ8e9CQRMGuch8I
n1bucDCPr9LEfWupyQQ9OFTPDEDmW8gJpOI3g5QAuT+VrcS2c/VOhtyv6G57jiVn
bvmzjkxP+4X/oVOvbph4113a1OSKo4pMfI3HxlSPnk+iBYMvZ6gFCsUf2/1OzWDG
m6jXuQ9Ue82lSZ6IwK8+einMp5VnByEanTqvgdVEntgDYCePDG8n9x2CthGgEZXG
NRVvlGka8PHyiYpgqLhxLFU23taL53JvFeXdXTRppU+uUmpETvgm9aD0OtnjCSLL
aM3pHpXEzZC3J3uj4ypokUagqtCKC6AeMlXo4o3B65tu/+ADGfXzLcJsFkvJ6SwG
JTM+bIlrN1IDpP/b6HjOqfciNHJ8noWykixb8NWYiS8UV1VFFJ15jjesrld5ChGY
nHYv8iwSwmU5hapBSRlEqpVJ8RvJO2Tas15eietiUbI3HFysG2PvZ5PAZJA5m8TA
OZqGrIVbtSgDEt3d1XC/hGHJiMVZanucqIAwAI9h3jDs26F4mYk3G45RdaFpzAz5
ZnHgXLedKepoj3dVAy80gYrRxbpncCHEIEL2XrCYNZev221tBSHibzfgP3gUte7H
jxvhi4ZpKMkHNZotbIXJtaJI2Do9xjBdaLqQMIBprWetbdDLy9wGhVUp+GDCW1rw
x4hDGxEa6wHCqJDsHSFUpZ07riD6wP09qE2ghCb4XEwr0b+ppzydcDt5KeiHvWZc
3lgcBaDWaWd41TpR1J6o/Au+2R34hWS2Jgjyx5VMGTZj+qpdiKRGnec82W/yb8gb
6IvY3ZAScY2hJTU4I/I0ER9/mCEkG2qaM33yUG1ZNXgcZCwjqmV4rCmTYLU9+XFW
q1bbwqxYmi7yAs/kekksPJPqqRaWmIcP8saMhBhNJbsnidsTSV+mU49UsnXKgvhD
QudftBAf4DuOaEBgNyp0K+K8mMHLDGlFDbaNqrKBehwHFGwt6wInGlgxuJQJHUZt
7xbjSDv0IDnf7SXpr+o65PwHMGa93Gyust0s8GGdcq0UsraD/0eyHCOJPiQmSJ/M
QUhbF13R0kGm1//Pvi/3EaCbvzZH9M+lnVQFUwOSL2TJKytct7s2kj9V6lD13Sr+
u0T6P+QNGg1JAfyJBA5Rn+v8Rz0aJ6L9uaU8BEUViFpPwL3gNcyrL/FydFr0W6XK
8ubsr34Mmiz5jL3magZBjboy/A/8OKkfyhm3D96Q3jq51f2nAPEqtMpv/vkCv2Jr
YjspPRPxjFprRGmz4GfZbbRvS51Plq65Ze715VVPOC1nfu5W2/smZ7BMo6Xb6HpB
zuGXYnbtGdp51Bg1w0EK9fR8WuK0OVGTI8e36L7Gr3MeeaYaJElesvhcKoWjUcxR
4542+yXo0/uFgbw9zhIflEkv/0X1t/NPMnNwlh2O98UIwgQA9wB4tJhG5Ah8hZ5Q
Ek7eQNjxj47I4PzTxMp768DcBMn0bAuKoZaOcZm4rnN0rj1trkdGFZDo5+nd/j31
S/OZR0J+8RQq/RhEi388DcxaSnJIebOYA1NOXWyAvfAieEqKuVAV0c2ERny3OjaY
aYKTN4Z/jZlVbU+TYVh+Orw3sut9ay+QLAyei0RH+fvvvRwtyXzHF8nwxC10unXW
LMnquVN5tXpIuX62RX+52dhzbBvt1R12SeWdcpVQ9vSWaewlWfiG0YocFnV2luLc
L/Ks+19KdkjUARaNNCDJUq8ovseDDrkMAL6iReu5eiixkz8kC4RRJT1QO7HInpU0
JA01AyC4PsCvgKJv5hqWHRnz7ZdYKXyZ47v9FuU69kt5asWOsWrna3ki9Uv2ahZg
WEjdm8YxTsEHmlWzAMq1M5rTioVIQmIZAkvHSjeFioHtd5sYfnSQXunLqwPnx7Jt
CtNPqEL8v6/qeW1jfOp5qvdDIzpvP0/pUzcbovicGfgDQwbp0MwrJTecsL3+aW7/
3/C01H03BJqysFwkrIIfwBViVhG17ESVgiXW9j7cZQILHoTk2mSKbBPlIfyBiIQq
BO/ZUI6Qiag1nlyzgQDlMT2KYCbHA/94PLseIxEoemFWRkkFzH6X31B6NRcHMB7R
bq+78vHFAklz//M+T0CJFPZ6f39ujGQ4FOcfQrbaBcmj9A09VEyGMSsuhtwAWQ2/
gN9uT6IrUcqZPYJ7Wo2UMLI2o8Vw+OKk6ett8UCjucZMF1yLw4LuMhu1qJ2Kp+2U
Vx9mPlvJzSYVoBJFzNsRCIb9LYB2aYVqU9IRjR1fI7JIcktrKrw6Ny+kaqAYKdEk
evI1cU4qk3jRfOIvsxmYte88H+c4Dvn/BucCVmJ+kAVZ09vDqkCtL3QImxWu8nHZ
PDXT1vtmSueqEJUJTRe6xE4NYUtMiuA7xo4g3xU0OJXq45VWQnMlV2Yk+lLTvnCR
3bv5etiik2dKxAuThIkZg3MSCkpPzeS15cprbLSDyXaHPVUbFNojjgCZ7KgRqr95
2jBOuB7vWfN1p7dkE8sV4bLqdcHuPZbtsfb281Qlsg98OE6xKtiPNCXv1D24INtQ
lqzsZeaQmEobCXpbqnmK0szYefYpvsHAXvjrWep8hNTCFFGWX81spyQ2TDTcDK7y
cPPMGVdju1dtUXERas/C0HSTJR//qwiLkZQeVWUen3V6h+uN1l1ZVp4Tyj7nsQPm
Ayfr4mHqyxIaZIhRCjLNvDHhnIB20r+xreJQY2yZBX5y1xsEZMwgtdIfPCUH2rZZ
82Wd8Cz5iIRVu/htV33601F1/LW+MlGw2C/y8qL3OjCndFxRBgTxwbAEhomLj/Gp
Rji3+eWhwfu90FM0dl61MUyhBX9sBbL0PviNdMSb5sbCMQXZIw8RkA7k1PNTwiBn
cle4YWPjj/+tLfEjVFnfYHz9DHtWpwmIJe9Y/vLqfS1bZmtJ8hb3lQ3q0DOcUTHy
hrdIh+R+yx0hcPruW4/saaDCLPc0xFliIbmAyrS+Fod8bf+hd8zpuyaD/wtf879K
T+7LWl92nOQX6rLcAk0B/bLh6QJliJa6oXtonFyEQXKvPtgjnBhJXNDjpcsEshAQ
BDPKbrmkudROCLdE+lDtoJ8WfiW+lDeB+rPCTtar1+OjJsFLaKiysqW88GUe2ZQI
J0u9QkWKjfREFGXESPQFna8wzNqwau1Hz+uVud958WtM9/KIVL5CzIJaCD0ELapW
wDVIe6cpcwnCke9AcWFI4otIqtSTsInjfCwOsST5WeZQq5ur8eyXHQyKm4Xn+tuC
AkLrfx2XAWnEL2lDIlU1pzhFBjt1zjLCTiAvRlMHYNBkwPLhXWtHBFudQ+8/wuP1
MRR57xEPYCdUmmRDuaAjpMvLwdiPzVU1xN1cN3weDOiiE8qiQ8v70EviWFpUh69u
xdgUQf1oZgq1DpDa+EKgbAJikL2Bf1Z9/EoClJaZfcR4+Vgm/2F2z6yFgcRvVJ+f
qeBVC0KiWSCS/WTe/Sz6Uv8X1bIH2JQvMuVdEmq0GeAx1/EBNC8vgsDehwQBfDEl
gzo2n+wSSWELwtgVmSk1d4sHxoroH7TBsp1YLp86hqJj6zdbd5J8D39MesZZig8l
eDm2+XKsJTNOCERhtx4ClgS3Q1v7Z2uyCZ+tucH7nY7En0NAJUK8mEo+2ncRYrGz
2sbMe71gFq7llrheBkw5I99N17X09FmS7KDk4tVepfQngrsWF/uBdLunTTGGQGK4
F2lekR4hYU15UeAzE1FWfMUypJeXhr+1k8xE854Ma8e6430V9t2uRw+CatVaSbQH
p+urGY/0A6Ji40mDkgSDkkqQ/on8lvUDxa0DCWo65i9morfWTBnGVPnobesmk9vn
mzrpAdtHtQaUR9+iNuUlfoSnGV1CUHHtFgJcWGp6dL2irfwj7l/g6/d9KFnfqwDF
uooY++D6wy1laWYkITHk7pJoeYhHPVAiAD8vFARkAZ9LkvcWuLclDH451yvsw0fr
SaUeYhZjTg40nr1IFMjTH4Dho1tAJA9JkadJ/ZpihYu2+dDhBSszoo8rBZW7ZqRS
mMdoVKBX/6/Zc7xNFR3uMZEvjdrbQjPn7wzj0saE5GHKw87mx9lVGicu2CbTVvvB
vkk9QVWHx4GHzcebVaOVvFspDjOj7iDcRxG2mnwTcrPLCPa0Qk3WpVbrhORzAWyz
qnYk334XRVVwJy+gIzu78ErEeV9bRSdj7Bcu3kel2OD3s33Fq3YBzTIf7WplnMp7
RkipT5NKcpr8t0K6cD60Ry2O+I1g86ajgsLIsAf3aUP63s8KmHvbalN3uFzlMAS/
4Krwgtb/ZcPKtmYgw9j7aQazszpCGMtvPeCi672ThuKN/fX4/zOFS6Be1fxLwdG2
zxrg/qoJ+7zEdaqgtz90MRO29I5X1dOm2VX7OyMkJ9efNArDoPnSVV5fU8LU5rpk
Seu6cj63DJ3YNtA9gzD7GD2D8nM+YtPH6xUSY2ifC/+a9359BU2Sj8ERddvF27x4
4aaqfEJlYeWifyMofTsQYt87frtTP7XloVHFLTcQcSYB92rdVHsXrI3BOFbryfy9
HDQXu6CkHjDzymSQDr3aSRO55Dp4iXAQNji/uoQYW/cvD2YdG7m+njh6L+l3bXT/
wmwKJMGuCSR0gVynEDxGT+74d+l3kY7DiCfwByTgX7e2pNgkD+EYe3N/fHq3HVVv
mAEWsTKBmQlSjDSScsY/9/TxrGkOt5sc11giWWm0sO2XxdX/YzmYJChpcxotT295
6IAsxkX89rCe6b8e/wNYIjWXlO4jSGewUiXq2S53/zoTCKhLeiLIPTTviRIEOmW2
7p72H/+Pg+r4h9li9QijsZM/YCc9AvK29WMzPAyIH5lyLosGx1L+5LEuIICrkm6f
+/aaEJ8EmIL90OSoiQAV8cTFBkPZ5HzL3QqBa82AJ8jq9uq5zoNXHCnNsGb2LzKD
exyFekbP0i0M7bSxCzZAOeOwwYbeWQyVx+z+VMlbK80=
`protect end_protected