`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1456 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
a4neElH2SodzYSxeJ5dQUhZ+Il4HxCbBem/2yjkx7Cfgigs+EhS9xdirRifbSaaN
ZOLMkEqNMF58GbjE8CR/SqyCTmyp0k5lDkn+9qiqyzO5NoNz3Zd9cfKFXFXjeF6o
PW45uj6Ct+XGgpGj4j9bIY/zEqkW5tZ+bz18Pn7irOY0kJsGsBKFyAkOyMaW2I0H
9SaNArBzOPpv6YSflW7zBuykHLg86F2Sv1+RIy4YbeDUt6ia1mGi3SCJ8RwcGn7r
FnprJy6enWC1Dq2DeXOv+iCbkKZuqkcWBxCKl5n4ZehEKCvQGIAT5VZpyN1GNTOG
t7VlW4SaaTdigi3cSByLvYkbjjMZ2ZwhfDR391IZUlGCpAhNX4jBiAckYTKq2IfA
bzdLt1j8ZFdlUf6XmqV//kOiMsXjeTbAP2mzdtCCksTWKpf8x4eTeQ4g3ZNeqLRS
+M+a8JIa6iWbU5xSJeczlY4r+tPKJYH3q3Zpg2p4sIrYdHPe38oLuOtMhwXbZq6f
r4WG+gTva+YvxyUNKafO5G2rOcCuy2jZ73Zbv3pkQ1bAT+cKszSXJyX7NmHmajn3
NF/+mtjbyQ11zTgbZJOS3VgxXI5Cm4ez272uvVJwzTvBu6fL3PMnF3PJ1E4Mo6F1
NkfW6d441NOx8Mdsk3cAcdm0LThonmzMVQNXAshKYcGtXuPOq+CLiaDwJNsKavrs
Gdo4dYZZSr0+SUqY7Dzt7+0XomSbAQnoa2OF0polE+QaKBFd9+WGwm9UjqKUXZ+A
GZ6LFIVnr9CfFjLAom4jHRutx5Mobvn0Pyt8hqsOpIY0YJNnFTsLxp/e1v2aijZZ
ReOipoqx/2DstH4fKXfQ7Un/3aD1UUr2H+qvKemSW0RfzJSmG9bzGd46j1OiknWi
ZqOgULDd6z69Wsop3MQ9ZbWrSFbx73ucndUqmHGREYBHeGEzFXonlQMKGb3mTC/s
Dw443RBSk2S7/TNii7UMRBtiqejZcxjz5hajUGQ83wfa18oP7SYK8UskiF6QxRxR
dEzgfqp4vzfOPzRGkVFl2DoW3NLisLCOtR7AH4h6xPwFJ1TP/eBwBIYnPVub0bKe
bbzrmzv5ecDlT8yJc3zf+jhIh3YGB7tDyqEvxG8HoiCBTqGFt1N8gBg9FAyBVPUN
Zshf4z4p49jbt1Y3eC2/ju19Wo3CHkPfuLPxCkP0fBw54RXBmpIHb4A7sNjFTOL/
XOwBa0HEf2JnbKykgot0XY2a2CdteV5tdhn/sHKhuiPicZ+yPwjvejeFWp2CutFk
17Jr6ZJRhF7IbDjhz1WZtnG+I8e3taGfU2XhJouRe6whRhzNoAOiR6rZ17wfJQyw
fEpKRxyJcxf5pSYqHLWxDVnTQTtbXWYpxlfCPCa8lbFef6iIkdbLH4d49zujv4Y/
HNJ5I04vAWriDvMtHzfc/dqt+YOO6sRctGv2Jt+Oa7A+EmdTYzySm0frxCujEaRf
sX8B0COT0q7Hlbsr//aBvqFkK/w5elT8hqtP+MNRxERxu1LfsZjtuP/9OymkpY7E
ZEL2/Yg2v2rVlhttj42l+97KVynQHS5i4DBKmTuafZbE9WKxqtcKS207ENlKwXuV
Wrr7RDL8jycKVvQPgbImpj3c202+s0aVt7yp8a5bVIKuM2xumALgMHjSkY6oAB65
5KrLJsw5FcE4wqXe2h7dMvYzwa7WIwfKAoukyUAdHH4Ba+bpLVgvxWrDfQAa2HAW
X3+/dvHSfcbO3XEiwUvmt/PMOrELD8AYyENWIFF8RED5c6nPZJhIkrnwPkrUY90l
o2Vpcy6G2qs2eRcWK+cYCg==
`protect end_protected