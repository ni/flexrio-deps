`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6288 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
BpTGUlWg2cHZljFhnB3CrPQY/YzBZbCewEnDvpvNu2ICJUdYcs/9W/7yZMC/FKyj
EIZwlvcn5FLysjkNcSjCnZOhsK+LVz4OxeEzhQeQSyInsgB1rV0d/pHDqJbw0H0O
dSjErAAiQkANFtcjfytP30SFDmIk7U3aSFig8amzn0mi6XvQLF2QTW+BASJU5Fmc
LJmIb0LOxMSpkA5kPB09nsw8/NS5zNouTFDatI0t767St7is/LKZQlUFZt+HpL5N
rn7LVk6xh4kSPV5t9TEsYLGZp8AbhQLa+bEXH7BLyfeV22OKeKJKXGS1elSXgVzx
jaYxtSTclREfawMsD+BD6nX2i5xgsCzVC3vcCaKzpb1GP04UW6Is/mROGyEeGgEp
isQDJcid1eA2taqLiCCALFR+biHuryh3vFtlC5bfWbw0/pDTTGHaXloF2WDoJcNT
Eu3FOyZcOgHAhlxaHRegffDDh0OXlZJ8AMvVrbrxC1abPRdPnYIkXndP0uiNRd4g
E6C7dtdgE6vjML7jhxWCn9gxe3HuVGy4alWKwE5OnW3A5iVvHK1CY6luVsyNhWGY
eeZIauklQ0GQ82edd7iErDHG+LKf6+oWpLXO4k6Evb6RDkOcsmnEPGsPfx0T9EX+
9ODBaTwzkL23wMuoFMOsCvppSBE30WaOb8+KZB9pPLc/7gLQhzEskfXG4WkPFilw
I27K6PnRNsFXqZvcxd4cPoSByvBFbFTOW4vAU2z4XLIUQ72USaG4hux7xgGr4E6n
bzknPDdy25w2drZZeJcDA9xkG5Z2m5BN7Tf/meLdbRduRepDX/sDMKx+oFcw8hTv
xpNh+MkyUWrLL2ItvER3yZrlNm6Xkr+k+qNF1cFKtHh+7jSs6ki2wjeP+tMhEJmx
g5tHGE6eAINSMrEYiOurW/XomvNwwE+0AobkI3X7+BIUsJun9iyWRoYoBp07s48z
IU0/TnnEp2qkD0MHZ7ikRfq/vokRXMU7pLUF5VJDtCCV0a0/EmDIuAYSnt+t0aB3
bxx16ScmkTMs/lsWnH+JNp6ItQAOpT4A5Yio7eJTNgxIgxPL1UaXE3FKjnIpfAKO
LUOVZDpEjlfGVKimbi02DHxSyP7nIaE4Jg2xOXwrmjNWLc0fUifWaVN9A2vHNEyg
hIMDa6XL1g4mNRwZIN+rBy9fdpOiNvC+jCxa2D9ca7ghvx5SF4s8f+UvuTl5knFf
DDrkd+AR94h2GsgzF30IJTEhbM5uDGrUJbSd43OYHm8wzqsMTTJw99nSWnJIdFAf
6J469bsOhob25ZE34SEDNoxGg3WR1SXHpfAfp2pkZc5GC061yjsj/mCitbEepJER
4QEyeEwWQFEkzZldCGow3h8OU2y5pjjd3zMmWrj4HSMTJ0FbUkbv0inb+vULzw5n
+0VaZ934l48JfBPuxm8rehrWuYu3P7sJjM8do6X/diup92YOOJ51T3N1uqNnDA77
mURs6BmVeW23ZB2y35mp7pMhXvF7SoWnhZC9NqWk+vgc3u1nS2oweis60DYuSbdH
9OFXQdCiMxPo5n4u8pvJFOIJIQt1JaV1u9/nKzHKHgO/MiZgDb2F09nxUporOmD2
heHF8TLn6meZd9vfDG2Pbah/RLEnLtaJERLbYHYlBOaNTbnCGdHic/hoC4LxmSl1
HiFgG+OhyFqF2XpDhvplQQOoYkutNcQNeTC0Wh85jF1MefzaBpadJ1RMUw7J7mE4
fJDr+AOdStvhW7m5AJRj9jCXZE+CnbYxrJHxyGiPNpfdzHlzqyMOHhJijzAb5NXh
C8x7B4rUnrkliqnPkW8bBrFWfIinTqkO65pkh8svKVtAehut6W3m0QGrGgd6cT9g
eF04SDFZniuOwITa25FThRWqZGgt8hFx7Z1ErJLj00gcz3Gw5s/al8GlyMu5sTVU
25ZN5C6/yD99/32EjJrxJPe+JmDq4T79XimpDvfAbb6NqoVB1ZbbUi7cauC2phLC
15wAky2u8nzYY2jHTcR2crOBvnI9TvC+VcdepJnZEsoOmSjbIjsqkVcbBsJj2yys
6E1opVfOxBaVBainhJ1hNCwNgMd0LzbHnDRv6QCEDBKwWLvRhlB55Sz/cpyNzNjj
KNB2dIWBcw4KdPNpqbp5OedssQEaeo8vQtyCCfJJN8dI8jUSEtzeJH6gZE4ChV5q
mQX9zUu9a+3mYuCyeFn1f7TNW/fgbQN0VXqC1GSaqnkWS02AsMenE771wEclwj9A
4GFmzDa/m6QgH2YMYpyEqtbb7K5Fi89NVXVx9eAOLNkq9JXUAnyqYycjtdH2NjTn
OzKvJt1AM4Gb/7mZR7mLC40jBTeneeADttnMfOrT7IaxhvrjYQMt9WVmJww8uzNp
nhp0LWpVe9z8xQu8jYXYuKcSdPvsddkZeN+QipXVsQsqryXbVGN362LF9SO3Ppfn
faAl2/fB4Y5wAAXzSx9M8ef6bSZO8dMRmiJCU8YU6M7TMt3NoMJYmWGUH806ucun
m1fJW0cnkJ2Rl5GMwzX7D/Bxrc6ww+0A9xouhgfSAa4b1wInRYSr5dh9wkpnVuse
nVw6gGqnTRS3526eYT7BY9ogGO04YRgXgtfmjLuNzMaAnPkiKmhsC+Rmgn5CaGNR
rWzzeMs5VUpqMArgD5AK0Jxtv1gBek0VqC5D1JMSNYW0BQAJ/COfsBK1GBQeftlv
IfZXTEXsD6TGsmti60Pe+5Kf0hygWjA0rOFM6kVCSLYqZRXHQXpq0ATcd8AC2ybD
4tlw2Bp8FIHoxGVSnZ2PuLlLCrPtwlhIpxdidUl571K/1mKZi6tjOcrRQ/qqpWId
NHeMDUIo/Ml4u+A+PJjd2tBYQ7P2UggV255XrcapOD/vSbOpmUvRqiNGMzw8FXdz
sgpTsTMIGIgrNg5nihdkGZ5vwJXjK3D9s3U9hlfqJvhhBjfky2Idjk3oepwBRBGr
UCEa6m81i6X233zqM6XzyWUCSkDU/ADEY7CT+wj0uQhktMWvdZdSQsE11+GWVU1q
xo0xPp0yt5WCH1FwCNMEzT449suGHvgeeBcRaIfol2aDo9leKe9c78UOdRbCfxVw
YHKF7xMppjidHBgSce6gBafmgWL9ZzJzZxp0+bxXyeBSwbGOzkLzjg1NDUw0gYHl
PQth35xA65/86n6Ir1yKg+oqd13mHbah5tuOYCaPMWCqooLdeSJSA43yKeFNAjid
Qm+m1Bn5RoTdDmPueSEwz/cL/FngKgFirKsA6ZRUAkmQ1we+J7qHJChLVruD96LB
DBvgaPD2TjIlp7Dym5pNwqAhBU/pGG5l+UE/CPj3fJ5pDlyg7dmjZrgZxLc9RZ/A
CFu7Ct9Bkzjv8xXF4OCCV5sI2XCqFb/XyYNeyZITrwin6kOSt1EYejYjhefVpdwp
SdGisLwegjgfqGrSnH2IJ3RdgYOAPkGSj3g2LuVo3LlLDyAJCxBiWeLR17GTqy2A
nCoFAA4Zl7m7HlY15+K/0H6LMy42g6q+wz4Pi2xcc+Z8TL3V8UpPSRzo2mIUz0yn
LSSHYawMsrjpuxIAOruJMavAjQWOK4DC7jZ508nFJkMROl7ZcB/ssu7fAQ/Ga3Qy
uOHgfjTXAQmZs0mF3VcG85DrQ3gHt1NFf7qWfODL6nrlupCOvjHXHFCWwiO6TTQK
w+0dkgKppjT9lDN4Df/KK2XPeIsLudGI2Z1YlBUTDubGB+7nm0H09I3HFzq9I7Pa
Bx/UaEUdzB67Yc/KptKz86+aoogRyjvcL8bDWOcKwLB/JvyOzTfRCsUZzGyaBtQx
M+y+EmT5JbMpsXHa+7vyTF/TOR/LuKZz++GarMtuc7UMvqIbHLLiOnC2JHblmm79
FcUEWGB1DHAmXmYkdfIXMTkfy/D9BRcGwmwdveFF0Ot5ZIksjl41iVdGmYssPXV5
lso0X3rpQIGsU1i+ex5N79pdqteAWsgiFUFejg1Koo4HEf7W0Vg2kmNSVee1OnI9
0SoIqZ2utJ0spAgM+kX5NXc9i5IWEjzcQmZt7sMrwR9sTQRj1Qu0p2oW0MYKOREp
jILZ+M7SqYiZ+Ic+iWfDmmnm62O8/4+jYzfS5NSzVdEorFTengFvFv9jsLtSSBQZ
SQWQHssJGAZJGX3Q8uwuxOud6fI0A7v7WQPGocWSKeWfEs8RvNHHlYuKpuQUO1YM
H2R5dGYWB75WbwILjJvnS+6xSokgi0M3fogIu180Jzd7mtgyQcmSpGBEntEiyfYK
qQLGPJ3DzOWeW/DLL81Cety6MjrzODb2URz/CrD4zb0pmH303IudnSUoV4GpApR6
hPNa8aQF/GjOARxmMJJlRmry4ROjkz8mw6jlLWRNZHtvfXVnX78l9Vpp3SjlVaEW
3I46PlUnQe87f1TPs0NL3Jyn4RSMJCgiBd8k8MwFS0J3dSzEuBDKjz3PFSypTIW4
4feyw345SzNVRsr8Y4xLVKGTVOgy6vXue2/P9DFCqmYWnSzi8VfqV6ULnsReHbXX
/v8bwcM/D5SbVTKDnrT5FZdYYCwvSgdgTBGW22zrVLG7+BD8oR1qz5UvpakaNlDw
pLhPDNRK48N1yWL1G+sH+TnjCYCsBeaWwH63kt59kOA50GCVpmZVYajTDqLLJrtf
QuEYc/Q2TCD6x1yxEFdU3wB62L3qBTWQkf+EtxM1EI5VdyQJPSDnzlFJpvOmw978
26fMML+4rfDIX05Yug4aDYBbEzJHxUMceL8n9Qq71kf671DKjPbwlWj08LLIAfd3
nz9U5vuDbZpxVo0SH64rLIHLX/eU49gdd+WODTvjkj/d5Q4SxsPvtoU+92kKpqXg
tmLRNhtB4zF9dpyyjmYuynCZ1qtFthHWuraNoihGKveVYX5jdBTsEVYYjXuFxTl2
Yxx9gK665S1aerice0672rMMpg42tr7MnoAw4+wSSdBPJbQxfrdVblQF7ZtjsYLq
D6rZbNHYdOQhdgEjw3LYI1Crb1FtL9TU/FVVrFx4a/srh8Qg1rYRTmScuxPZBsko
hXW6fMzx/+nkvMichWeK3QXkAvu5eC8be+VZ/WbWWDfoqKMA8JPlAfArWwKwYRWo
eBk1fK/Ybng8Wb/vV5MuVTQ0cKVd+iLRn/oVY+NxXWMe4upWWaXlDr+nhzTbAt95
3N9Q3O+CVBtlGH1PzdBKshY1ZKdYb8ImEk/7cWmZUZKlOohF6LIhVIu1ksY89Lli
lofveOH1vGNseGZi4LxdPwBKcG3AYUHth83rC6HLRgdzgg0WIkifHoUlh+LsaD4o
vcuckt9f3L5lEfaN0gKi4tATv/Bdqvw3G8dcWzy3wHPUZHa/857ajlRW1aZm4WI4
mj7lnf6ZfVQq89RCb8FR0KHFxM/lUqh1vvJ2shhLokXYAa2LlBBILL8rlaNEoMRL
2Kn+zvxensBM/T4XfC55vTdC2re3rKcfUpm1DjIesRKZpeMmaEB5xpVzjMWdRHrl
r8SkfALrGPsVZbJ0fcRh0ntk3v4nshxaWQCb6tGugEBWmuHAQsVxMv7t1D7mYqqx
EC7b6MPKjVyMGt5Ai7nMG68u2DdZLxJ6OyGbF7Efx963E4/H1FH1yZ7cQKPqGixN
uUFsCg3GaaifGHW+I2h9pOjanbDsHPgTwP75sUua1BYtKlDwg1z5m1uH5n4dzvCR
CwdYyC4B9oW4dC2VSKLvVKpfYHfQ1TEQA89+9GBfq1HhpddAo0ixQgJDcJfsVCQD
6NifeRY1myv9nfH5t1jp5wmZ1MaGnmXiXK1LjBCujCSIHdyA4SqmFmXpiDEWGBdP
5+5NL2W9oSepdOmJiDhHAnBtaYnSxWFtGt1Q1QPxvDcu4fTB8N0gO/oN791Qo4VC
ZdgRprYH2YsWtl3BseLObZGojFPPV04U+OAiBUzIBUtSBJZNX64IHzI3I26EbTKO
9SJSZTS0auff/h2oQZJ8ORIXEbcvXJlkgR9qlKDa9QA9RlC1X3JtMRmJweXGUBJq
pxi1IzZIWgCrYQ7b0RPwPRbRLu3YO9o4mBA+BbFi9TU9ZRRw7ddn0dWCIxEIOH95
6wrDKTgyemyV4YFBF05KQnjlp58nWyIyRa0MRJhOg5pU2YIwz7dQV2nKTs9ZU5o0
/uBp3YvYbOPSvykKjOJRiYq/jhePLypUclQr/OEJkkCy54zlW+O4W6ClhRBUW6sP
NOHWAPBU23Jj46NvpL4aDIrhksKvOZIEtnC7n00fsgzSds0AI6gfwUlOB8MFTOhX
yHGIzfEfiKsblczEEg4VWbIAdKsLZa7D9pd99XEjFDwewMhShdKNPCYGyooDl0ti
Pk/CLVfpEnCssLgJE2PCW2qOKftKxXgvhsyfuarRas86fbqFT65HzvUC8dDd/CVD
XoJzytZjiqamEcSXTXrOCdhRgPiisP0Z2D+1R71WhlCZLj3G3Cu29BwNOd+m/mIL
sd7WbUxTYycQtLfPdOoLXixAsjV7edlOpJY1AabEaS27b1I8TXCNn/zXq75Kodjl
mRXu0Va7h5EqOuksma3WcTlTpUofwsTlAOPI2ZqDRhUSE8BME1tbFLcvOykP6b5L
wmBghfwbPf8HQ2ze/ekmXue1OW8mjjoLdHzgvmwfEgYSwWZCCEMLVdEij7tQxeCY
c3hlQ6QIpSjhNEtZc4eTUlq5q19OESfvUfqD4WTDkcr3wcBXTJW+ggQ1Wk4n6TKI
ubM/rkbm7kQNezqjCTYBRLkVm9qNmjRGKR89W/Er1Ryi5bZY1BFr2bPeZkjMXShl
JOopqCpOLcmQVe2iKnl+eXqrnex8QMndh6sRw1WLk8YD5mQw/Uoh4DBUX2a4LIvg
6dDrOjtaDyhE3gL3J8Quf0cxMtfAyVzRPAnctqWLGhJBlkzKN4sz3gRGDLM9hjRD
592ho4vh/7YFnGgLyYEqcDoCO40PXbYT2I/GtB+cmBGHDQyGAuZZsPBB70z7dPw4
xfaOaka67984g1lLqBL7lAA8tIH0BJprfutyVnsS2H0VwERN/nL7ZbmyA8AK8mma
jMRw8kKWxQx7s8/StgYuF+FQK27ZccniS7u74rjLbzCC6UO/zUxbqvysJotz9JQ1
oC7bPjB1Wo2QWxWHcxwVgoochC1rBxIlq08keiOSouo4mWibncljXebycF6LL6Hc
vP3CW5z5B2PefiFnqZtOpX5FNtN0nVCfJWaIh319HdInLMZQAOe3fbeTMSmcJIyC
nofxEPLg0wy0XjhjcsgK5vjmXzNADmmqFub1rzXmJxXm0phTMbcruUROj2cBoJWp
wQPW+l0gD9eInHGwY+YEtd+mEqvbR05+mbiWWQn6YNl3RWDrwq823SdSDGOgsH31
1iiIMFJ10H3Q9EvlKShJygUZqgVC9AvHHm+I+GPoA7WGmjz1V+hu5n14tU8ltX7I
5pY9q60rlnuENEXJN+gT+qfhi3pir1YR5YoaH5Pw4mWGYLvDLVUWR4DxWS6RpsHs
KMqlQKQ6GeZhzGF6rbvBPNVnMB8H4c+v0hBVtN22EpiNbQ15q0VxkThHK6zOjfNO
C/wESUc49Ar/jq9JMmMlZ6zc9rDVue7sTLTdzE7evxyiXLJO5GvMEtpZLBxIPjlw
7pl5mKN57NxZjP4NeuM7OpvjUzQtxX6qWim7F6vnfh75YYXXyhibhxUE6gtRJuaZ
LlprNqioJm8s4aV8Bap+Y0KE5dC+lj9sKpxYyAenLMKiUEgKWNEeGlSXoMQY88HU
FM+FRGnaLw9RsP5l9u8VIOPoBvPcdxuKofIQCN7Sv6K2YMFD/fGrsqYHYCB8rXb4
9EQo/gW9pN8lb3p++H6Xns+dREMdoVv3KmLuyEnvJlVoN2cKWxa7V+PNnw93jlcV
UxvN77Om17xXS4E4FNS9YxQsxbuEwKtOE3GCX6ObEqQN7izxgdib97DV157Wauw/
+UR+uG4a/N1eUTQFhCm33U6sm8h7wEr8WJVFu7HhUthkXRYK88pWal2HxZBAcLxq
yvz5CNNWKLWQbxa3eJg6ME2gM8DpjtW4svAef3ifjQtCc9wguWRUHQg78cjFEFQO
lH4u0Uk1Ww5ubddg9D41pDalnHWWtMGYgEM0F0GfDJxAwmOHk/6XN8MzTgLK2/ok
VQtYyNjbyQ2Iz3GIkfdMLm/qzq960M/FTdRODiI0MDri+ROGz2S1YtOhXffOe8Ly
/r2HafZeEIRtGpI48XVIRVHgE8rtFaRmC+wQnWiOQWCTyml1kTSBnEa6wpcaGAMd
3KsU+BEzUWQJiGKQqHcXUTdmjOL+ycv02U4pGXS3e/G9W56ZhseGXRAQu478zWeF
`protect end_protected