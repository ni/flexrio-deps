`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 19632 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
akBpHK9XojjdOyFTP3pOwlqmu3HKDkgfdD3J9PBzA3p3o63GPHdzNoQqMFvwio/K
aSi2W1PkWJcUd8Kg8v63LlFeyZBkRoUn0cAhg3KuF9IaZpbqp6d4aQpWhFYeXABE
81hZEZyEqm8zObFZhNrCmXtUKvJv3EySb828saDJPRliFz6wh41RJa9B9y+sT9WV
ol4JAjviK60/9agmupko3xsbH01BJuJwZLQWfYyGqMf19Cq4uGpIzp6qhQalQtWO
Td7W84/XU2FqUhDVnQ0XTqaOMM0DMIi+qhDFl0Z4o6Ge4Q9d01VKQlaRS4XiGw6U
eG1WwguwiyK5BZ9laktx4OTHSwth8f7PWPcLVYuluEgn5UVTJAuVQJnI7TH6onxb
oKeSZ59dmWhCell7Z76GUjRXmd/qA/Q+qCg2/oamfJDXlNLfJFNgcR8iUcZpp67x
bArkVTRQiORr2od6Zg5uZJH81HT5jIpKObgqtKoDiWLJUFHggRGxMWXtiHPZKnHd
wxW/uri1fBoNywzc3jZdPaoBJ2SwhVi89pGduOg6Mde87JwJZh4GLgS3PigFWOCH
ahmQhjdqgtBC6Cv0Pb/DPCIQnelMzVlG+nlZNQazceBB+xaGiSTWO1E16tcrbOkT
jk3gva0OAJLfxsad4Xze1YXpolsLjh0nWH4CxO9VuhNpfX6yvvN6Ak7eVXEYgm7C
wGH25X1Er0gublAQl7vWiXzQdMKhD0Dx32zQqxn9Cza5itdYIw7NnD7t9REBDZFV
V9imwRxCSYYNVNx96+Gt+TjXW46qN4yeTHqUyQuMJOVeMGtk3hxk3kEhfpGKmD/s
EcU8JfzXGTIV7MH2t1ul3HFNGloZKm/K6XvEKdISfOeeYNr9YHFfCL8NWn34qs3M
ZHn8wJ5SSril7RqLXw6GjXYdFknxA+R6EywBoiG14YgYvBOUrQO1zhMj44R4QDgH
Tm7WKaRt5OotLwgjhTag1rZa2CnDOGX265WRUA+Vvf6UgM5sOQTOwj9GrhX+ZWYi
eiJ7NGt8KD7D0M3DvOFr2IZwKnvqXoquw6zxDVt5BKGxGN2tZpyf5HGNdDz/9EmZ
4wOMZoh8EqhG08y4aNO1SJbHZNPFYUJSyhT8UYvNLrQYfY12VBMTv0gHtsL6TWR8
/ve6wr9s8Ob94NUnME8uT5aaFc7MLbnvZBgQPwf9RXGTY8vyptwyGEJrQHOIIZuL
934kkOuuoJ1LCv8MKji7VCgrOTmlVnoJDVe4KpSijAYxwMKriXAaq9huj7PcnOCt
WnV0h2cHtVnpDHRR9kn6HdavCqjnrflGGKV+zVf7qFcM7WOs1C52NeDU5Vci9aHV
5rfmKqAXLxCc3khS9Gx0WRTr3eigCHfHjN6l5Hdd+sTpDPs7Q6SilSXJj+StY6OF
44wrrEKOElrTaZmAFeXGiv4NksEseCqhQOIejt9pqkCkVAHpixL8xLJgKhvwStn1
w5gL7h0V27Cp0f5L/aDByPPVGsq45/cyUPXHY04XD3aKKRviStkOEV11fFEE1Ixs
nRKfGKUrsPbnud8LYcB8qY2Lfrv/oW05F2jtlGylvDz/TeJCTAPDAAviMriaIQF/
VzAV5m9kDQ66tHK9eQzSyZgCkaKemdcsH40W/xMOMZSNFLFZv8MmZl4hnXYYpbMF
NaF1fM/tilqZSx7h+IZSni8r9h8A1S/vHnM0pCCfjoq8upx2Ilcbg+H1EcG0/iea
8lj+jm1laGXkdnf2iT+8SIX4qeMyU56PDw1dq2qfAEP6CN9W8T/6kEcP4PQ1EbaF
uAK5AK2DejRaSZoUTgaJ6CKEXRiYLsVCjJbtN0Wvcdlgs0CvnoNxN96epgDFdTVO
lPBy0U7RVmq8vCeLkUmFYN0SKmV5P73Pree8D/L8zwHCJ3cNDyHFj8NkZg+5LxGD
S4/ULrffDWbL95Z5kezZemVw+zaecvlL+QTPnS/5cb0vWIxilXH/D7O3ks1Rf7l5
khjfNKDmJnbDK063/SrcwJhntw7C79NcIBIj0kb+FJhpVXfr2NSNIyD7Tc3ezujL
TxW7pMpCOc0bAZyf9MFvB4H0PHSGS2kIvYoo8IdFP649PXBuoWT7dol3iUGWJ3EA
Mb6so4dpxobjNsLO2pskFs1S2Yto6iCjXW96HGRvjtMMuziJCskPW8T6OWwHsW+1
PS2LLEW2yyUNjb8d7TWZ7qUBd9I/TScwaRuOYCnmuLadBChkBTso2e32u5Oq1NlX
sJzS/7sjEDCRZBa7pOsDEgNSdidRbsQEziaCWdNFUeGPp25UuHYVWEp0QdMv+2IH
/kzl7WFR/A9s5jY9jgHRsqxLOdmVbFH9fyheajJp4uAXY0WrBRMCCNN+k0GD8Mlg
6E2YFhkYul8rdOtphI4OA1QzD4w1LOg2i4AYlKgLY3aoRWxccHm43on/+dSh2Rqp
yB8Sfmj/S7+/Bb8WKeyADLepdctm40ZNYDExrANXboZ75VuO4n5FtyQKemCFS1UI
dQ8MUldpR7HoHNFCWcdqTNTOHedEjfT27OLG9vFly96XSsqjpNfdDhFa5au1oxb3
2KW7Omg3yvDITddZ8L9h8QF5xy1Ae8qlScYOsTf2VVhIYQmp4H24J/ZSkOdozfXm
ZHMyN2V3WPVrlMuEi+tCkM7xf+r+6eTwSQ3A2JLvl85e9wIPcYaAga5z2RVQb0wH
wgMedZISGfpR7XIHRs1mjx6dczYa5n8btPIwJ6/N4Td8JSXs5KSJIyv8b7MdTSqK
H17mxQ1N4Lo0ffHruKQF8EaWAR0GCkAbKaZNbDzmirfcSSihQ2Uvyefkal1X8keU
50Tw2NRLYgmImHlPmmUVzdozCfM0DHfJPyaCyrk+JsUetW2J8GjSvmztzp2vkd/c
UhL89WifqNoOtxIhhOZO4fKJ13KH5KKXyIUOuvEOE+rbZ2Y3gCmTczwk2ltgsLeq
iZXY+PtRCEoZjqL78kWefuW3uFJ887P39wJYID8TfKZB2WJ8lYnIq6zA7t1G1gLx
/xY5AhDk6xW9rnmtrq81JSM9qnQ+4NNJ9A1Ai3V93aEa2I+u7wRiHi8ZdpgIyZaQ
Kvefa9r1rC+6SPGsQym6p3lKrhtJvuv4nNg8NZ5AiJbJEQCubRfBLiJViWlJeuaZ
gBbuODqsjYWcMwntSAgMZCDwX84TcztANGRuh7RDA4ocCd/QQWhPfhTW1StYBX1l
tWSHfByKT0AZJn2qxE0cJTwaa/pOqH2esbkCvgYhT7yNDstnZsHWfNdw9vQFLdF9
HLND8yFOy6XZ4mP2j2igMzEaoWNYKN49u4P8XitTeKMwcSTeXYL9aHbyvNvT0cv0
NJKkt1iMO0WZWMpl4MlkrSjsDMHT1XaIUX30/c1BUYX1aAE4HkZu0hOcUjtZBZ1A
B5rtYaW+x82dsURBOKFwgUK7v1n7t4etiHY0F9RyQxuS94bzERCNtx6Tw7Wc9NOq
lbzfJcMg+1EbWQ0gD3LKrYjgRKb7AzAottpYJpxW1NSmbkhI//bTeUqucwTwBYVn
Fk/rWRJBcYQimKQ3UuHYa4C7cBCP/VCLCDhs4MWEiJ6BJonYwszHQgbgRpwM4Pl7
seTuAX6Pudn/yflF5awvGmCZkNh5zbd8tbIEZPPTGpVKbmGIJaHqciysMv7WDIAz
MAXSAJKgcApciZpGSI1HScGe60M8tfPP1aSh3sEdykTtf1KSfTkxfbOhr96j/D94
lJa6JKNGpEZrkVtKNeGQDb7Uwd/ZX5zKT0qR58LQrsZ+8SAKkAdqEkPqRmjg7Uck
Rc5TtUtauen4/Fl8NRVyi1nOGVRpf5UCgRK+8au/HIcJmyrjieFX421cjM5tTe/I
QSfxIqcG9qyF8hdZmr+BogrbW5422C8q+cOwtCwI1kyLTsttzhpgHBl+J83uoHD4
8H3/V4EzizytCJ2lwYDpKcYqKZdCdn0r7ysnMZ68Y1KwgrGgDazZv831xujt5aQ/
j7woteo4VkHyB9/cXXZIj7m27nTodnAfAz41/wXS6zlbwXpHUJCZifg9nMuDRqOF
EWjDuReXstsVaZKr8OeccAmKDB88yWF4x3R6ftqZQ0CEluUJXv/auG6LYspRfBot
z+4ia5bFnEXrRPmd9EggzNlKtTkd+zVx8L/x5wlvg/5/6P3p/lwTXIxqyAFIUMMv
x34umpB6ucdzwGt6Lj2IOO/bYbwcSDcd/HDbrHsZVWTpUT1ejI16UW2+sWYVBJL6
AQ4cwFa70sy9FpmsPgJeQeYvlDkyzFZfbrvfxjXjR1ju+FEhoRDFnYcjm8fFENxT
27Yxft9aUGAddxbeJDA2Lr4d8+D/ddA5jzySijUX0ZyMaVhxzBoOgpMi2IxR9uYK
+Ck2JIi7BGaafKAiRGiUKYJnOR6WqawAioPTMC25oJ3yAuLktK4axvoSWnbwYafL
Flt6X8/Of2WCYzxxqumosvapI7KrfUsQAmZbHSyWwCj8vDl/cxAw8UIgtsZqJ/wh
THjU3nphPezJUv8OKY4INJsyhqpydxmac71RoHyV+Jv1ghuUcDq35zq7CwuxMwKe
cKaA4WgSWQDjanopOz19IpZwP4Dx9mBvz4Mxief9CpzTp5rFirh9xx1TG5g0hm+5
kaZrqLRVsti3HE1++L/9d73H9PL2UIh3x8tMSbE7EblFsS7ZiXb3UaNG4iPwVjLG
OX0ZVCvE8Y0JWU6xmqrxCPvwTuGqZx/J5j9xxc+wUTo6bQNRXPt1Wvgko+LIDRK3
+PEQbVKw+W0Xwjzs1NFIXNWqbqP1Ea75LJneUphQFIGBEjrLuvDutS9LH3zkyYCb
0YbIsnxbvTU/8QZqo4CyA2G73YaeBG/2okhW8ZVEKWprHvOYLUkbA/gy9vST+JIL
bzlklVw5+vKK1LntOiNZR0/2fe523M808gAEtcSOTytlg8/AErBLOknvWWUnVGbx
1nwuaJSOq96SuMTy+Z+RSj6gP9B596VJbYGCzKTy8OcE+KywqAnFf5HVm3jt5MAs
Jl2Tx+w9ujB8wlzMUlHpBlRE7kM7WsvfZ+SLeShUuNa7E0oab8yxEICy/zakhkft
U4Ddg/Flpq10BChlRseidQBJ+9Kue6Nlw4/RGoFoCGtm6PeaUMQ6AXcl+81jzupS
+6NMH67/0L2jDgVPnXMOX+7dqrZHHAKydjxxsDrm9PVobfQYRCpZOD0WKCQMRwMh
VTNlm8+j1+8fugHU1RRPvnz+uHICyJzd+Rg6+dSphrOnl5HgNx9fuT4eUaDuqZeE
e542etf7tIaki6wr3E0OfSCZ7S+qsGPP5hy7L0ql2rAdwGyK6aM88a0eBl2pOkgL
u+bvs+XgUtTZYd2g1Zt+j7Jbn0JsDINYs1y3iY2E2Quvz3WmFbI3m4j5/0mmQUtw
X8kJop9iXkPpGfWadFIWXQwsdI1ppZHm0j0QKVnx2+gqxzc4f0AXVN2M7CA2ztBS
5dXtAvmYRs6XDaOGEz15Aapjk6s1seMCCGynir2c3ZwY8Oq1QYFMwpzeepHvyeo/
mNmRBxSBJdOSyZ/U6QONyEgZhLu7SgK1bKEQ2fMscxpSIb9MYq7yuPXFmE/LdF7u
AB/2rLC9qZBGeKmCdcdLLxCswQpBwlIaE0Jvz9ilBct8NV7ccQotHGGnr5B2w6ul
TgFkTS2Ux9WRzXtmvRqQuJ/e2Zc9WtLk4KevE+DBzzigCRUT0RUNnp+0n+HtP+Lx
3Xocd3wnipuNaJjlph5Pzx1JBl3kjrPFNhielTMdli1Zy8EREO3LlEqNeW7cTmr0
z1PTc6bztR2mm3ZTj6eZp9bfz5/hRAi4YgTAyP/LF2On5fV3hq/k3avBqM2fIp/1
PXUs2ymxsi2/X9Tn0Y4d7OiLeKNXxATMl9/LIkmidFGldz17F0Mogu9sknpxQRjH
T5OAFWBUWljcvS+VFBVvYFcblX1xwyKe/ULl1Ob306bve7Z7R7K4ffCx0Z1W6kRD
nMKMgVp4kRKyoJ3JqZTxahX/aOpe+uZeZtm1enKgUOGIiW5fcb4gZJysZjzq8xJJ
lZZUMkBmZdrFLmV5lI8qguHma4E3/Td89Xy3KQt/xxRswtAew7lLHtpM00RPMFgE
0D3kxHbyp3XIq60BXFgkgjOGDGIzI3nfgiJIJCXvtfohD+bHYPdAjga+g509eydM
xVJpwGUfePed7JX1qGPtgfQTIwhP4piCQssxVFr+zDUW95Fg1lE+i5iCAalbNWzm
6gPC4hDjqsiSteQKWRm5K3lbVwwPoQQlYuYaub6mDe6on0YeelNA9IhHTR+51zac
e1lRMWnTOJom5F8pniSUcu9OWWzli+IQTL0aOEs0DcF4vRxE56Wzuelk+l26Quh4
6eUBvVflUQu3cljt2DXbhnX78BvUXXYk3XueK7MKDz3OQg7j6jyeXfcdqkl32HI6
YT8Gu7cjjSANAa0ggofV1wDUE8zXfbne7WsBA+3jB/2+DdkQ4WRFRH6BjFICm8bY
vm+C1zOVxankaTkstWNGL2YpHwILWcv/ofW3zbILpPIWnsh8nk4qUgJtMGNA34Wu
y/AIDWqa9S3HqLmg9bOdTBEmL2tA4m6hztwAIXjkh24xjUxRu+XbcYxcHN9XC6uI
IbJYo8DQ21LZPOcedzzPJg4YAAnydbTHOThfFvpculQlig8ARBBfXmFULwwEUJ8G
xH+zhajqUQc+IFpDglfrxQSQ85Yqga1DS6wU1Vvyi1kvskF0dZRA0fhxjW64E5be
rC3qHBGZVPU1c5z0rFRulb/pg++PwWn9y2S9SPxPMBDMdUrICVEylutRsEaOp3TY
1oojjY+RS1uUtqlPw+QQZdwQf6uaEsDpyusbd3V0H0SKw3BfPGnNXjyzu1lRZX1V
yrcmVaTIMoDQrCa2nSO5h6O+0r0FwtsC+tD4qo1x/J0axnH3Oo4R44jL3CeT/Crq
C1knrsJ3MfLgFRVWSvTIvLQWd80pxSffzZGsTwGAe7tRpv71f7lo0TK5GcAStuHb
o8mnUZQFu+Ho9BUCQsWeTqinophPIQ6i4VKLBG4+WBPB5G3ZGX2FeRqhby9noLpA
4p+tu/qYnaLJyyQU0srvjVTwG4gM4LngZRLNwJyh1MuAXYiM7kAneuuscXi+DKhC
+tcGzo/7OCYCiqb5dtRwD/Mgqv2qfK8hbhOppM2l0jXxYgKisIrgX3NxSaKovJ/d
hfl07YLxP1tFKIhsibr7tftgLGAndUZPvPFF0BbzE+4JBQEx7z4aLcUxhL+G9cxk
Wj0/DJ32SatBFzjZkb4BMQ2dj5fCV3EUeF+PDOOl+gKssf1mfRxjLp1s7T6d0WEd
2onsqoCJPR/zeW1OJjny8lyC4wlnI5O9LdVIerrrOU8+8rEY8k7cpBM1n7n8cT52
U0M4GntoKgkll7GxIhb9xCzxSJA1f/43mhjBSRln2UWX8xO+DG2y9dWMiHWeC9NM
rSh0zAYeFE845xz332caUfc9uigz9DcZz/5/GcPm//O+ke6q6Ar58CeTaj3I3Psh
cgs4Zd2gMceQMj4jzylSKzMF2r4+UYm/G8f7DZ991U0KWbn5O2wQ8FMW0yT6LS4P
6RGcmwNv5zoX5QqMusJbIyBWOS35bKVCTXyrWRfL58g7vrkTkMbrjxb+nj7xSTwV
w+jJ3wIlC71gXx5lk0KWltbD0WEuHo3BtzCyYFXhyO1w2GOZjb/0UrL1B5jc3pkB
3SRzCiFGOmLnAJcJi/ouXOR7JCNJ5u+Ct9QuB+W9q8nhfgM7Cyq8bmPpZQqNBmob
sJaPLyMfW/9xt4kA8c4lPzjrVNVVSXHZZ7Og5iqtNz7fGHJ4mapulQPJLHmcDedJ
UM+BcY45QWaWdHed4mk7rWhasiRAGQJHxYkMKOcPXkhZViZW7VQeI16bS5ekLAla
orXO918Xft4KN0xojU063uwQJyU9CO5UYGtD7c9Zkdv4KgfcMhDwVHiz6nIEChOJ
NRi6Ec+1RaE/9f0eCxjQF5LlWt8EZmSJVncAbHHJGwvSqiwUNG3LDIGGnRHf02a8
LckUBOFKvC6YSMx8SUZgCOM7ooUrjRx2lW2NQ/9jGl6jPlbSLOmbzZqalvChkAQl
4V2GftolMXJuZ0Wujj9Ss2KBtUPDd1cGY+WHTt4aHmfgq2yynTq9laxMBq+hf7z6
zQpbV9fe5K8WxORymzu6jF0/9AI+ZJ1S1/89lH4xGOaRUrnan8cAaWjNJPNVDsKu
uHX6ZJnRJtbvrnbxPF9DhUYmOz4BZScIoSHc8pjBIyFkPDRRp2U2bZZstspoiKlp
EbW0WVuHf3+5xveofDWJBelcVoyhkMwWjX4WWfR6bG/bXVS1ZatBHdLwW6Fc9GBF
JpXDkLwPXJeJbvjrw+XavwLUsG0hLDdp4OxFE0sjnxij6I6dja7tuwcOr5kIIxu+
T9DhMP3XHAGoH5Jg1n64LgsIourS6tgivWHuDeokT7GFM3K41VE6QPGycMHQ3wj+
HA4bkgcinQvg7a/Na5h22zz3jHReqdky/EhKzmXbeaduuWSrX9xUvqY/6RLi3ZO7
KBWVQvJ88kAxl5pzKZu6WehRAyYJzSGx1FYMBt2kBgd5uUx9qxdaDrowh0+ihR+S
glDJgC5Vw9453+TJH/o7+KAm3+l52MC5ZLZ0z5+1+sA/o8mE/K7CGSylKfevLq+z
8Kyjds8rvbEuWDeZOSBZLKxv8MuDM90Cqbq7mZR3MstFccean8Q9DrJOCoQjQ8Uo
irKHShFYSJch3W6sq37o1e7JrgWkCkm30UMCFXzVTSp76SBE8r9lG4DhLZsvzzu+
S6bHRn2zwTABINoFj4rQR/W2MJ/SbZip0r1SOeTHwtTL4Cva8lpzotGhPzOEeRAX
xvhaDU95GYN4JLsLmIM8GDd71pWi6GKS9lq5QfHjCKh7MyVdDsXieRBFNb87WhdB
p5VCSqrQKVQnbEEzo1HbqmpzAX2Cv48Ws6fUgF0Re6HMR9DoSteGqSRyl1SvPID7
q03mf1U3t/vAROnnV466FSiwv+PRDI9p6kTx/S1+1SC1xKcWAVU9GjO+zI2BoJMR
Hys0tm7Pp5u8jC8VKGOv2x+IyslUnwimu54waoAtmAQJ8eMDn6u55NC+XXTJ1ORv
I68EMxi4mO+CVitPehQRYwh6PFlOWLBElhkpmcf89WZyWC2qCheVDN12VLQYOv20
aqCoW3ggREP64Iw5sptV/Crti8betSAQD+xtr8rE7maIfnguImJXXxdcwNg0Gx98
KWN8K4KsEzoghlaAxICnz71JN9DoEZgAsqvoPMRdBRaQVhNbNjjyQd5TfHvVOrJc
I2WTGzx3SrChXhWOyWyiH/jFWe3y2JOWpQAi7scE0MGw9yZ87PLPDxiEK7vGjwo7
/ke3u24saOVTLyp3dMLQbM6dj9IzlivhQ9yi4+6eTnu+0g+yRRgU9tMSEfeqlgn0
l19NAk2nGtYIpH2jRChgMIxXDJvycRLsxLLWgWO4E0RRkcgzjJQ2GcDrmwFwTbO2
23JrpCc07/82WKdZFkWerqLw+VH4vRm6kS7XWz42D9zNsfZ8KQBxOiPZs6lQbka2
9DIRLDQEsDISGRu+l5G0Q3QgpDuH/LzeGby9cAi42wP1sqlo/pYbYU4pc0Uwwu79
vZf3u+56efUJQfkvjQ/S/gEm+Otj/W31DIDfRmnPr6eHB4gtqvfsJYnJNJi0Owo8
gsA/TKJTubXIU/u24+p3AgfuUaGCS8/85KN8nLdj++9YokjS6yMjt+vfumBe9hbS
hobqONTe2LtHkhcZkbmeZAJyJQtzcMBjKEx35+jMLmuQWOWSj7BRb/1siDho8j79
bHrhNF9hgwjrREAlsrz8DHVYMCDsgkpGdCVVZtw9l3ddkYRu+6JO4y7CJkiyDrMb
b9WpQQodYC/DRFnWeigdZOLVFfGwRv+aL3NAo2Pzr/hSFC56tyAqZvXSrrTU7YMY
+jqbYs7MTebfCXbjuVVHjIymlMIyIe7nc/HDpm+EhFomQ8/do9Tgysm437NWJ5pP
Tw0X5vAh68k5hJGinoKswhXCMy2Kuy/7EtrM4r3Zav5OU3rmnPwidGvNFnLjfSMY
6eEP5v84M9HSbBUgeBsA9dnmHphqTLB9ZnWijT2MWsCpxdKFb/pu+RbhGuw553Z3
Nx7wzn27B7kwtSrBI0iWEQ8aqJEj3jonwLqOpOqAkEtVZuHDjlwZfPaKBKtrpzAR
GIJAEJZKjKo1W6pkfMSsNcuXt5X2WhWc1kAokylAMQrbA/wxoc7iH0CrH4dbOh7u
8vHCAxaLdmIa8eB1GmkRJOx1iK9Z9Prsl0WJT5TZo0CzWnHZNCVp6acpxl5BVbiT
MEk/H5xs9QMH4lb1jGmGBryiFSblee4fSYVObaBiMiLCeQ0LLX1C5MId0P+xVuzj
eGZDJM4BTy4GmOMYRKwp0+qXxz/zJXnIH+MmqjH3pCLhZv0i/lnhmMkNr/ljEtBh
5DinsAASA6+zpDAeZJ/OEnZ6UaZDbKOqnqLKybSyjUe23sbHxIugChWQKKeDZN0B
31bfjyMvYvtTq2y/TV0iygfvW5FTnaYi9mHrNqtWcKJi6kZ5AEWENvAEYrV5t7sG
Wlyl3KBv3glTtZ0ABlRD76ArHJAEymQR61QFnc/o4XMk6WKkQRyDU2CvDBD/hHKH
hZXz6C4BfuW8knsgVrHuL0PI3kAxMrQ9ZG3u4rAu0LfiD4rAjQ84+yljuug2mDah
s6+Sr1BPVCIbhGL+NmtBvTsi9InBZ9cjPgKyS6WJIxRFx5Vs6GDRAFQ9Rz8PVDaP
3bZ+8j4NQBQUgn2XyKBfJQGWO6W1oUzfF7VLdSZfnWgeQRwtqgX/BBlnrWEq0OlJ
RKdgt1RrlrXLjs3cjhT1xeb7OZfsYcK0AycDjjkI4A7gSKhPnvgW1fVL7RfqURHV
o7htowV3Q1nbCfTzVZVYkCeEOTftO//VgruEdU3NAOt4HO5SmL67jbdGwmLL3SZv
iIImDPNokOA1yHQi2oW6g03OhsmdgTpiUcV7aVv2pIfiEbPWSYtaM2fm4ZXrOUTR
+XDIvHn+zEfQ9Jqr7CWDKUKQnGPfI1DbytNgEv7aVQlxXCtVUQkjRVDgEGAOi+Jv
3KNtUHIStwB/nGzsmtjzqSeVMjp9wB2h0sPGpcXuG1IVTmJ4Qc+Reut575wd0ZkS
tVOO3BVgJUzAUcUC2wI2d/Y9+17m6psVcBKJ15JwwSdqtpl2SWQ0c/60F8HKeuQM
k53ik94t1Re+TUKkcITeI30jVZWksd12XQozvopRqPQYwdlOS5LRwG5jRawU4Gix
MvECiMfhvHI7vzzpE4f6qRQEJTp7fLbKFpdaqpnasvFYClCRuFKS9tVZAGpFp2Rd
NJ2LeVEtJcygU2AH0SIu/RDmse6iFuLRkE8zdrv0xX2FOrjZphIp+E6kG9Kr8Q6x
t+kp69dmr0TdOg9F6iqf8TqcXujzVIQXKA/Ig8wFVz1rIeoK/cfvSRHbiYgxrIjT
ZGVlTI0XWh6/ymqnXOHOPDjWzea2G+OOC64Kk/ZkGRrKnr0pTfYfp75Zqey03Mlb
R9QhznxSq/Ny0jx8sVyqXWD8DC+7nZBuYVwLFca0pl8F3SmTqP+eVqClNUEy3G9j
3fGHWpS16M/3ss0ciJ/nS8EBE1poazc/8DK9DS11Ao9IeABVFEw+aeTdfaQeA7Mf
s3nHT/lGUps2TrEwrmvCdBXZX2vUQ6Gki/8yOUELuNreMZKPei0v6mStLst+XUML
O8zZGQ5GTvLuRfDO5MPkqskp2bbn8xy3dloq+d6Atvp/G0NIkztVfZ+iAXbAPiFp
T8DZe18sJFEQhbag0PyvZ1V9PnGkchqCDoF0GjlWB2vorMFj+nLjQzOPWOBcCWpo
JGITBRrBPbDwO4xEA32F8+YqaerkIdq8qskg/8nOw9mNqFyWq8PkXulOvONKmOm8
OAPboSg6RJGD/2CMqVWr4XFaBwygsJExCgY288hDzd74LgGcEVqwiii35p+kptXF
aHLYlXHOUpSMHX4Kxg5/pVIB9BjqSwsdccGpJ2xS3LcINOiXivvS75nEUDXnIwrN
HcE0LDk2a9qMp5jtz1Jfzk1jkJHxSAhVYFvJZiS84yg5pjkzvShSSYefQKEOxC8B
wdTvjyBZhkiSOFMvrCQrkY9n0QOpqnAd2jvNCNVOmf26TCpTZGxtxORHjRZXKi8c
pvCavUBRn/8vIbBPPsdGwdSLBt+j1+mSukihThiiy9jDDJdYQHObe7rPtM1NMWAn
39YtXxgk+G4HH3V6vrqrBduWiiAgsIbvM2jRvtXU9g8cty01o5N976pL0zBt4z98
u8mEgG0TY2IwiD8UmzZtDsu3xXObgbyY3bn+2hypExw9EEWDlw7HMb52m3/RhykV
GkSvx3K3O7xYnptULm7ozSdij6xwNqzRyKbaTJV2HdSJ1rnE2lzWa92MwDeElvy8
u7T97waOpYWMHIIOvTtgVdtwfDophmS7uPOVaw6ZQr+qkbmz+nVGNqm3/TOAicqm
NwmKuNXGK8xmUaxHU0Uvz2KIDjxw2HkyF/Tmzj6o1pRjcKTLIseNM+ezr/V5idIm
6nyK0WmKjzcceWfnXn/9kaP2zRkDJt/dDa3906kh9+6+HwXzNaDkSeYtR+J/brvr
2A77FPaSFaVOJTaIP/N3huRer3xLUq1fQCMzjJAQ6F1L0s/8rHz+lsaEQRth7ihb
dmGd4RxwPLGzPUsjcVRjl1q8Mw8eaIBfN+92wzgc/9aIbUoniMVhN3J/yq/tsZuL
vrKWF9lUrlhFTqb+JfB67abVYn9mBMyNuOWiIpspRCefU41Ko/MlT1Sj08MQNK4/
NGgLOtS/Lc+yNyCRqBTMWw3w1xgnRnnMKlvoLYRAp+USZBJzCt01cp/F36voR0TN
ITZQfzt536JKTmPlfdy8G6CxbR7mfKynW2rQVBYxgFJuRNcUR84mitMgJkjhf+Z7
9kwA+BGLxfJbAwF4BTV42QPQgucqUtTQQ1d+x1nRDTpK4xGUkfxZcetZ08PQyvZg
LpUpwVnrnFLsTG1KnobVD8vXuAL4QXA5Biqfy4+JKHOZ+V/g1956IOB9UfriMHS8
urusPuRLWk83p+0ROhemaVEa6L/fcsr8BzIMjM/XN2DUaRSvYraVSPBGbpxkr+la
SnH4GC7+sgSYK3nSBBi3QqgqvSr3TlyW9tAGv9FYQdj7Z9pdimYAWMLzgvkqg9Eu
FKav7M84ZQjSnbJVP3m81b4nMhuk3euPdCkepU4uy7dFS15xV+3GM6rGTCP8ulVI
WvnX3Jv31EbECftz2HQIOMKyiLzTJMZnfgBQuupTvIyN6OzpoGSIrdK0c1KfrW90
X3mwYPfF4IWX3nZATi7f9WIIgd4k6NNCaxP9wKhYSyPZDWKdR19cP1bt6z+Kye2j
oRM73xCcZRbeqs6vJQXOENdP2OKluyyH2owd2e4AD9R126GIfbF6V2YJv8CnWAjR
w10PkCR7KGDjnb5goqvo9lLqO77OVZ6SfXTqc0J8XZPJrA97f6p6pP1jBR0WQ4Ke
yn5I8GORwpIOOnBR9VquPzctpkbRFgAzkKQe3suf9DYqm7xqm92qnRvrS9CdMXFx
17t0MeBMQ3seEHo8GybmPWZX6Vht17qibpEH3O7Eo9fuXWb4guXkKADl/ikeBGCg
T252pD68Kv1kCTMZ40xVeLfeEULN55en0lk3bMUfiR9KdBaxCIsCN+twbVQRE1dJ
MkqCb0XtnUKrFb/rGnv3Yf/Oa3j47ya5acMGJI4zQ3gUWu2n68wg2T/SPdYvXvht
N8KTVUiz9xi9A4Izvw95H/C0W68nPkHTKH5w3gneo3Az+GM+qnVdCZowcSbVMj67
Cor38rOuuA1+mPNj27BLQofEwOp/Jz3X9eRTsGrD0x3LCrq/UP2n4KkTod4Z0GWz
uHJ47QR9AHgPpxOkP0i3z8q24S0fpwxzrumDJLItmS7UQu90yiD1iNCdBLOWe/jV
9G2wf9xYQMemMex8mebBSitZsQeyD0RbccFaxNuf4+vycKigAc6Lwr/GuzGuXr1A
EkrOusI7b3kMyf2uzZUuPVmeoQUr5Bu3oRIggPiHwR8vbCnwg8A40GfHqAA2jJV1
zltYCiepblyd5AqPbxaWIfbU4NZjPuM2KHgoiSTa5WUKl3uDB4+0oBzCvt49FN+/
0H4JbKPIT6CjUdtgQFNAHRZw7tRzRqYfjboNQMVkargqndmMYiHuiEjeRcBUwpYB
kNYdvUwVMGclupkwW1Ox/M5HgTRYN41k0Jex0V3XyphoNJMylVFbp63iZT9eCft0
wmQhuAvcCXSy9gM0QxEwp9szWi2FdUKKn+Y2hBISO1ucoSMab+4j5gLq9EcVD4i3
84IApZLgxZ1ufXY9HDMNLmbdq7zRqzoNt8hswlGCEMOUK3x2afV2GrccSAIt2fPQ
NupLZap3MNWyHXgf8U0dF4TOLOKKc8/8We8A6We1oCjcBIN8PZQMp5vmW4IuQJbR
jr0M9+I3xr2snEuKw7BNC1Dq/filPee2Db4snX8wGavfL5Lqgh5fd5VGSWnl/x3C
Q5W2ZbWHFh6APfxX40g9p6jF4NBT2OUi23ClSfaSuezpCMxL60Z0hGnepBsS46u6
Qjvjwdljqw+TkLhBoKDim5bnMPyMvMbkndjpYRVg8xfdvhGuXHdNL3Ln38z4d9aa
lRNsc5Mvc1KoI+1U6Pw6g/qne/ddRqXn0+p4GytSXy/UkoA3m+hCgwyzNPoQVgza
3IQ5/l89TCN4GCedJZDxCEF/EiF41j23/rq5jp1mvX5i/Ywr1tKxMxKvsnn8ciBE
jUhw4KPdQCNaAcL5SR2vfISj7re2UJLC0SQ3yRcYhBdFoc5eCjwVQt11js1jlJ/8
ZgR2OBwIkblcTWBqggXZ9PSmAfeixijkRO6y2zhoNPfGC3kEMHtVVwpx8X5vEnie
tQgL+ELrRGmXml8AWHNDJ+Uwp3W/tUbrpPZ8UgymtC32C5dN6bLnCSciROCfOzRQ
dSlYzZtK/EzgeoaVUDjpKQc2iT2UpwFNFl8XcVSevBGEoM8N/zPlbGw/G8pJzDN1
7YXKzwzyTBITp+OjIbFq9J2Jo4y2TzQe7M5zwffZ76zvyqbxI5EVvAQkEde2Ncpm
nhhoZQnBnMZkPPRIfK18ci5efgZRlK42Kx3dActk5DixcGMlNlvom/QBCAcBTeE9
G4eP6n1ETQ6WQU27flCVjUA+k6Wq9/PJNd3mf02K/1D4o0Vz4bo32K+qWj8qbL+c
Fn7puPcbD80AVnurIdUVDDMUex7QLUj9rfa/i1xuWM6EPwIHGJYNrp/IszoRdVTz
MpDI0v0l8iHJo2Jc7+E/cuGN0esve6Gba7AQESJa1QzuFwAcMmSGh6bqaoh9peyr
zJurRs3caVpyCPjM9Jvzu4rHy69ASwTLaOIXP4XnVSWDp99eBUOk/YBmIkHZs33u
0WR+/KepdBZ5si4B2JQjchvMSVIvVpG9e7SyCKGkOhaZ3k6FrbW0bN2nH6drigQC
xOiDtbg+2URa3duOgIYu126lYyDnitG5ebww9g6cxGE6aErZhqB0GO8tR1fpg+Ld
oo0tc2ahsV0WrH+v9l739cUUD780icvMQGAa+PTdyW0YNfHt8bHly4T3cETPb4Xo
5POPfAuAkIfta6GT/+m/o3xv5hmx28kxMaYc2EPU/oJ9gy6kJ4eDaipBZFA86dVu
Cr6RtFYnjsoO4hWwvUGPNhk5pyOaLdu6VoIYGfWt2h3VY1Ig5v0g345fI2gacMnL
pbHY3JlspYf0D37m2XG3sV20M71s+N4/KIDI+mwVobYhM3rY4+kMyP+CwUi5bHdz
xdCHAi/m1k1z2ZgQCxaYC/xVtBFElddiqVp4oLM6DPlQpgt2e1YfrELFQuN/QZd3
+Ie0g1Jz+7DoUnfuLD4stpnHDvtcBiiR2UZTVCBd1KqQP0C9wcnYKNCecZMbJTQx
+rNezbsHnWSAw/V/bevuFpoPp3yCUUAdE/F9TyZ1x6k0CmdFSpT+6qa2/veHQfuH
KzXjF8wO7QwtePeOIFRBOeUvXqeonhYVgTNcFoyqforjBWY/mgOD2qWiMWawBrdZ
EK0YArvrCXizKoLSCdIr6aibr0QTQG1xdVYxi5F2D/lEhxVkPgY4MS8KLfNNeXEH
GXDU4v+rDXJI81ci+TIhIwBremmSDavY8ThJfOhI9ik7nmZLa5JLKMdECLnYCCdC
76A87LftUiVckspdfSElovIRFW8eFJQoaTNxIKXXxh4eHJMJJ2jaja7c5lBLyqav
wdDFHitv0OZ5Ikqiz5fOuMf0DTTIEwGHfzC7hT7iD+oQtoM6gMkce7GrrLx0dIUx
b/SBX282FIbtAHFxdVdJq4a4FkRusiUtYrhURuIjKJ6J3Bg80i6d5+VLHr22RLZG
UJ3PYgKPITShgt3ZhszxQ43BOC646QBenQ9mhllYhfFCD/3MbPDAKPLj4x/pBb1S
YMOIbdX5HaBuB2WXdcpZVh9dfbnIjsKTrihY4AIHRKiNxVqazPGbRSRVbJN6sDJi
sO7h6R6hPTdqKlk9G50nz07CBC9cfVPPwgE/y6mpuwZhwGQhWoXhtx3WWGWH4jT9
fOS2mhEdqmrhO/iV6H1x1gFg7wM+QLUQH7oIWPYigJeod+vm8iDlxr82APC5YE86
K8ki4i4ufwKP/8vMjJK/2vpFCGRhBbivQ45WsWonklDuE1HsnNwj6COanUzGaOqv
py4ZwgpMdMQQyAn1wrZTHezmiEBNxlhyFUsR3H2YZ7vHx9mu4im6MLMuKjhq8veh
9zN6yr+2WUn9XBChugy628kK4ZP0j1ZUw2DgMaAmagnUK8ZO7rtQOe1Fy158VAvO
z208AyCRxkPf0ewJY1N8eTdsdTcJi3SPtx6YuwtVJUGW1U0RPDdZmEHAxhG5jYK8
nsLrBKdlfRGLAhj/a7MmI4+5qJNYR6h6axTDUC7jA9y8V1rXvicci8JpYhnZxVwS
B6cPXheBkidawNchLkZN7ap3PYbvRtcl66g8438d3TcNpZ8trv11uPOy5eLPo7qj
+ltYPGj9rnQ/16eRFGI//4mjLZI2fgNH/yPnFXEtHe/WltgoGiKmxQWP8yP5L6o7
izj2YifGB1bRTfco6/25a+xKmngHSamlGqxsCcc1PA2sXtLgouKdvREHjp/eRYs2
N+x0ZKI65nlr1gt2Va8o8swxpKHmSGtNeCDl/EEPcZB3Qby3HXa2A+B98NdwiJNX
vUPZhWCmxyCo+rE7NmIeqcs6awKGV42OfvPYuYTGgllrufRLcLq/Vaq8H+Sf1coJ
A50NCs6pX8PEFyAFLP4RvxG2xbbjTB07ZReqgcQE3NY+2DRwbSFa67XkVF5vme93
Eqfm+H+C4xG0uU/IK65wqgQVKKpCOxJKug3GhVSUutDoCi8LQ/pz5XJOYOwo2ayH
5gcKplz8VWf11C9Z9S4lbiyWuhA2pQJKaNmBuSqwPrZogzzH0ujtMkQ5jQLrjQ69
WdBkezll9+lTDZJuUuLFvPavXILOM4JsmW5dExmQOkecCHvKrnnVuGpxOmJkc7yJ
loVuL5YABl8WpB2EKyqG7x0G2R8YPgDBRj284Zohud6lNIyQxQbN9cQsdz06ExLq
Z/OKYPI0pW3xS3iD8myvK7wtca32TnIeKLUYnmcWqgVV9UGZ/07EsVcN7rYszCoQ
QT1smlbBw8s5Gl8XBekxwJ1ZLxxhSKedjYSn/JNkLdjZ6LAWFmAjCBUTCTE8XC8f
Ur5KPYMcpHSIiJ/eTJTbeosF4TyyYOWo0ibf6XW8sqoKPbknRiYXXlPwx7B5Y0Bd
tyOLyuXhBwvD4Db1xlqzbpxx0mAFjtbsrF8Vlqq8cRKNAhXR3tVsuH0hEPsZkt9b
KTuRv7lLU5i+SG0cU12GTh7n1cO4McC0k2Bc1W8ywbpQw4YgbAWJE6eCwbwT9ggd
6cBf+aEaE5YbSy3/Ff2vgFMSMbcNibaRTn0Vaf+0Xtdcb4bmoo6faS3JSrScw26Q
gdGYB/K001fe3jyOf5OxLbIg8m1Y+sWONs7A1dShD9dGPrBsmnrLHg3BF6IQwOq+
jRO9itmTINFc8G+XFYiBlu+ZgOi09FfkXvcfl0OyGE5/s0VIGb5gmXMR4AqBubkv
ioozYACUz8laUGWesNq8F9lI+iCfDWDBFJDSjihAuMBDl2P7FE0mepml9m/35zJW
Yy6QtbduvpPxizaO6ceB7McpYshZXvytv/jW2zKlnShbxktpaoDCA/E5qasngfFr
sggt9yOYeBLiQhD+OQ6l5fchpoa8tPlzMTNTfEYVcf5HQjwpm7Mh41JmFmZ6moZj
FwJ78l4XpnRjYTrVnRM/UTlkREXFqkP75SDC0UT2nIrvfkNhLfPr+l81i6Ij8NiU
WvLRk0iW9mBh5RlZF5Nk/a2rtfVsXH+1MvlUo2QrUTNp6iYeR0z59lF6ya/5zyVT
EcOUBUL9Jp0GHL4pCKRopGCMbBY2G6VsjvBoOnvPIvwsRbJH+AJtsSsJCU3KPzGU
K1ZZIovEHEWkrfVVFMAHAW6A9rdxQ/9TGYlVqQT726ACBpaCWDn3WNL7//2qWcme
9Gu7E7UnGPuYinhTpAa/8QcW9gQcFdyHxr3CK2MjK+Reo4dz3cJP1y1KsnfBWbOM
/5ishZOVd6RCyncllaLMbqMwtua9OB4uVhoSo6RVfddLJcbQcuvWxaiiW1SrvAk+
K5Jv78L1Yeerpmzfge9lMR/h0DWS00vh6kxkd4vJgqpfJ96733vkMsApSPY49Ne4
rYc041YUuqnKdgy/FG4mKYq2QnaUe+hjB6OPCZc+0qaFRTaxOe36d9jT2O/pUWWm
opqm2bM49nPOM8qO8gf5f2RUuWw068jO7pP1SE/ZT+ZF4SxJUm0RguHEg1c0aXaz
HZS31pZyY8tXvRjI/YmbqGkLlCk7xeCuVvbuS8mJrWIzjZLUlKZEGYu9tBmkBA7H
NwdwQM/YwYbfu8l1g1JvyM4yIb4WbpqirJFDNoGxjtFxmjxymx13RadW2SSlnsLq
j3OsN0pEh+QtzE/xjpWrgPggCGqdJDWZSVHG84GPLAhY6p28+U7tTY5Vjws9fx8A
CRvFspwoaOwNbTOppa5/yn3YNEBmXxlBKfXEhXnuNtcxtAmTMnf1HjIw7xfagtri
a8csBqzK7qfkTxUYPhFG+bFzPF1vSXJgwDCCctc9+iPoqqTWJrZw0cpSuiVl0bbq
T7d6II5fAfuhjtncdZdk34gdVTd4uE5X6FXbVeVnYJa4vwB7KkX7EhOLAYPrrsvX
LO4VuF5bEbZKNm15p+++775HKhGWXAo5Ec9yF+vbqVUW4M/k/vEfHEkNGRAxsIYK
Y68z0CdzJLOXgIgstgHNaOHntdWEfRtla56DIlC6fIa1IPWhiwIU+HTlMfbvX06J
B+6XJ6EFpzo9czjPrEILx89ET+XFAwinxF14BS2cT7B+p8DtYJrECmYZtGvn4lis
zw9u8fMu8BL88tJxyaYU43oqvZpq8IQSHMpxwxdPVGOiuuMXTMLeub8p0wx4q4Aq
k5oMytzsck1oxi8qf3rD3QuHouNrzjSx234YTwFeuxvOBqmpz24yam3ZKCZM2sEy
jYpC+ucwMV0La53fn0PuUujE3JyLxiRqEt13RHf+UZ+8wEKMR/QzdPfaoXBj77mJ
6UpRISqK9jbeqvhdxWpLEaOnLBu+fgRG8pN8bj/BsRNr1lJO9RkloSoHzFBbDoYE
IG8p7/vl+qNYqxum0KA1wnlewivOFurtrR2MPA8FBgqdaua488OHO9JdMrngOPET
PawzXTPy2NlfK+R7A1hwRMLNTZB2t+4GnKDrfaC0KQpilDsxoUlvxdx3Fw04LnNq
9yF7QAYhvINZGYSs+iGCScQVD2aNBeTX69SKrFBe0xZIpOCOyM47yezWES3Pu293
sVjTbg7gpmAzG2nFbkkxHbIHQRHvqa/5UWzlAFyWm3VRsyArnj8o2zX8rWCTV33K
S6TZZEKpRLs/pyNS6anATEfBTO+MQQZEx6gIlhhyHu2SvJhrU4B4ZVAzf+oknwnn
I63Aq+PQfEcywhHgzr9RWQ5nxWE6kDveXqOnnP1cI+ypP9EVTjIcgswq6Q4xnMYu
Xof3Udp35SwQnsl2qeyTpr4t8D2VRgGvI/FOr+OBXhQB0hYPjcPhMK/G4m8fsQ9N
zSQrXkkTwrBoFviI5oIXAV9j8leF+johzloaDSLg1BFRLje0VwanQnGkz1yZHBld
NhrilSLNuNacAS1dWHqUYi6HBaeqmpZDTnxjW6SRUhpYp/Bp5w5MyLR9gz6GT0Pf
0pFeBsEyXEVO+oUEm22nvwIRR3yEJeSyNzy55yDSo2SE5rOqkybSZZ47eUFoMmPd
FAHvZ/Ir9+1/09Brfyf1ErgqqAD9j+yPABSNinZdsxYcAKlkBBWCUvILKMpWzpsw
dPwulzWCS70jx/2uUG7FqPfUDEr3fOb4bsFqVLravtBF1YdudI2QFKfGBoZ9vfYq
Z8B1QSIoVGGjsl+QoE+87RDRqsSAaEzwFTBL9OZQ/Aon3hA31dCmi1KRctwpX2l4
bMS+Es5wVkYcO6/xeuNozq348Z5rNddWnlt/+ZOl027lBjIdS0hbNH/JZYiLIXnp
4/HAdz81KTCHVb7Pl4Aj/2eV7vFxiM8CaMzvDaJdAG87kiBpbNK3WrkpBd4Z63ow
yIFV9bOc+g2jjTtWKpYKXSSidrPwSYHJ1rZe2+jiKdBUXAWg4ZHEJTpyGtE/CYRz
zbrloMi/kWu32hA/mK07s1x6nxMXwXOcDv9LDsuy2IRIYJpV9Mei/k9tHRGjEJh0
KmOisQ31lGroIKHonf/T2slf1tP0YbvMSMdNbR1K/Msfsv+UrLlgXHPzYzxA2AT0
qpR/foEzjctk9iPPeUYsXoQMc1Ogw6vEmUT4AQ0QztGVcDRF8fRjjK1ruhmojFSH
pkMdCvyEZdNP58CBglsOHfgZcNn0sxphcL2efK9k67ZPUeLCq7e3nxNGFdneYKBE
mXX6XFMvS87hrBDOx8dzqHKctigZv+XeUs+l3PRp/2Y8z9MeG99Qx6UIo3hq8UvN
x9NADLhdah7q0YD0MP/fPWMtamEppminGSHRmJw0a4UZKXOLiybUxS6VxZe7Qspx
jMpj/YRy5yIfUrd3D3kViwK5k/ySEXcNwKnEVUl7iomU6j0JZ3VxSP9RySTWii/j
5uLlT124How8aOEx1J+e6Tj5/BeTOuIhjz518hLq9brRwNd7tu2/0Np4KDvDqK06
rV5KP/vIAkfQHT1an34+Y9QnHGdG3OwAkf6fWpsf16N/H+yQLTcJtmPTnVrfkSfs
urlyDN13X74bsbN/ClITWjF2bkMaqORjdTfSE7JkDwf+4t574Neznk2wTqWUq44A
D/uj/BW3LcVzgt0R6vuLBDzUsarh3f2pNHGx/RpOPKnvH0Ku586qTE7mjSxWKeOZ
Px8JrUlnQe4qbm9w4zgNEqlch57tHn3JIJhBB5gUE23clf19BRHUWmqnK2mixa60
cmsc/9diPzR+K6PfpM+xFKdbZ+k6mRlzNV/8JM/ZtW4EI3V0MqXfq2QiqvwVwPh2
RmsHb7BnBS9ckLVIN095L2RT88XLQyB9SjHfNe0n5ksxQi1RxiS/hPnrJIWaYSwr
mNj2+zOGZK6CgJBFsifiLlZvw6pnisGesSS2RVqNW+xHmUVCyBTptCHFGTvz1mu1
6p3/Mqh4sbldIXlooB1FBjDc8E8mFrGKasQqp18illL//gX6iy0E7/FNbPL0ugRF
W5dCFNYb4DXFRDIQalY26VAMckcAp7tEGOd/W/qyf+Cv3PYsyxSS53VQ/YQTrdys
gyplgsaX8qU/s1mTuh30kaenYYOTGSDfZQkLwEFrVuxBWOa4vhJtMEXNjXeTRnms
FlG6JcY7v7CuQ9H9Ih8Z/bpNXhfBi4mpzVxybh+w+vmjzJqXjyf0Dg53OAcT16vg
6qLsibDjaEUdo6Kg+IRyxy+iWO+fMo3bMGDmWEo2wMVVakOWz4ZOIGkdpS948JqU
LGqbqZvGAWtI2/fYLU4OByso45iG8AvZ4qFcYvA8B3qIzXEMOtRQ5JefBUrttXX/
1IKTXmSbQyI4t1D43g6FwwvEtZfqe0aFVwonDHDEmkPIXQco45YlWXAkBVA2azai
DQzRO00Fjka8WNExeVAAvjnJckNveewlOxwYdAQgaQ9yYbM/DPOF0taP8XARAP6b
SFvJPi6Gr2ca7fmedMZGgX7JRoST/nyJbyH5Vbezq3Xr7M9ZIaDO+jHo5xU6MPKO
w7n3IZyZRTP6JL25O49kC4M0TT0IasDyE5kFnT0u4InTNY12ZgZ3mZon+ZKKZF62
oMJ22/tRFWpVkhieI9MO1Re14aXEZZZHHd8WNfgdE0ESlaBWQMU9GiUz9r0iTKEb
KgALLnnM4OFIy9ERLL5tEXUgravqP2ZJXVM5GFQb1WzAZjQHl1QuxLiyk0L0nIeu
CJ4ojTgtIyRdbPxUURNkF6FIrf+4R/h0edILQ4sPyQsFkeVe+gM2X42mqg0okd5u
K0eu0I6UJ+8dUjk32WJNxwaDfVn6QQ3jNGAOr0Zczml0nsUWsUrgsSdYpODpHgHA
+2BhSgOEYXgjRRusZY0nirxMhVvmxI1cu2h0Kfg7Se6KGJOfZs/VdMFxtC1b1kjC
qO0u1Jn0HVeNzb134Q8ioRrSjljAk85mHfTlcMIluvtEwGyN/UoxIKtq5Xs/dCZ9
1CB9puYH9p17EOWvw0IAGiMr5CeoTc7WrfMCDjttjwa5hgi7MDwfZiA2JxH6R41I
F9vOrbqiI9hXOyBwvoGLUhDThivGXyz4JFVW+//Y7wqIPdw0qS3qx/aJnCVPhVDd
4sl+lYbzqq3+1zwDhdZ2rwmQzJ+szeoCyhTaN5M6ED0zYc0ELDlpChVMFMhEYlUl
R/k+EMP+8HiGn/tjfLmnFPMlPTb8ljM0UW7DKI1LGkv3QcyyYpxQGx4XS4IU0G3K
18G3hG7CzlnoGEo3sAC22Dyzkb11kHPgy0bRKVSu4+P5Z306x5a8dIdI+UnVVYC1
kVBgdMe9PJd7RbvF/vkkxEzkdoL5xEPfxq2BN/AIjw2nxLn7VyXjn1GmRMCWoOFf
mMV1nKPsL5ClsrkHNK+NM+5TRYIPpKQw4HwEK3hDRqRvpxVvIkKXcrphR+CoqO5l
wzvrE2urujHk+H6qq0M1R/18fhUX8OdXJKUFkTvvy/aE4YxL8QQGat53zHaKQ2rO
MacIfIMthZplDSIhZzJXScRfrca75ZklDAmVf/GavS4UBQ8ocNp/vsmU+WSBAAx9
ExNyZqraZUst2NRfKyj+bX9IsJnqPevVDg4KlZEjaZv2/gL50a1jlG5lKQ7hF39G
VZKBJGEL4wFMXrPwPqrT3x59caKxbzxh2VWVuuwBBNRNPjtAP9RKHfdrtESrjKSL
7GzFIR7esv2M+MXzGw9FDKk9SSe1f/FEXHI6ZJlrClkieEbGtej3HLrNZaiBnTrl
XXFq7GJITAddWZ0EqHb0tKmRKiMx9WB6ft17drZ4b0mv+AyDGbNNftoT3ynLAYoz
etPYYTWH8ch2tn6rvlpsSAAodkiPwB99gp/s7nJU9312kha5bsKfaJn5tXN4hs1p
STBy7uKT5Kz3QeR5gIqL5QilrmxklpgHoV8x36H2MTLoRCKcYPEhkxO5PsjaO9LQ
deCazRqh18uDtfa9CaMeNKe7g+scaYIPRO6CWeV2VkT/gKZ+gwDjpQ8iIvGBdl3/
2tR9CDKy+H/pgum5R6zmC4ta9HVhnxDyxKWejBU2W6m6KGeSdUkFHvghJ0QznkUg
4zqrWVWxyFgcl6swXLEbnkIJg3eEbVIpzR2vD+uFx5AgnWyPs+bKE70x1Ra/stle
u5EvJLPcgj3RmeYyEO8a1kgZqQFGP8PHIzr4aBf7x5wfyiL4LDMtpxSYDL4NKkvy
DNl002FBrdp0wQaxoi1FocqNS7nhU5DC68tXSiuEKUkP3WXLckjOXsXFMsk7MA2b
B6rKMBz9F/vlzeHq//oy/Rv8ttwhrbDgSEbd/4q3nFNg6xR25R/5PRs1VdzzLf/v
PcFINyKCM1EviFuAlzSt3dVYrFOPSMozfAANQO5dLmB9moZUV0Z+2ObBh6vrXvaP
XaoHxol1K0+BjiiAYWgqiVC0cuUQS6tN5mIwfYLXxsU6ZrcxkKA1cFLBFyn5RNKP
VhCDUTiYGbRz4lM7vMcRZq3H+x6DZsilc5A/D/DCMRRrtJU3QrKAwI/MLPzDtOoo
ZOPJC/XmcA9CPXhUfDhhOvOU2svABj6BAmPAMF3xxbIdFF1p30ZN6oUpQGpylL2I
akYXaq45jIZ2S3BEcZ+ATp0sDMeVPj7vwDexvyj5SCiuvvYRDtmwV3/UKKEQR+Jb
ejnDGeM9B6hcQuk8TBU8Z2HwYOmZkSSW2D3LPy3uz1ftg8Iu/obqcji+78nD4xka
2oWZvq9yDzKtNoW7fLQwyIaL2rNM4rBgx61e9qSZDrjBGnjDao77ldAGhw06emFT
Qw5FrkBHoF59hVU8wePehpCfw10ZrYIxry1LY4VbdP7YOzZKKzpNkrtQQB/igZKz
pOuSBMbCPuI5YXtB5oBELizr8laG00hB1D92vtnx9Mn8f8PNWCdLV3X+s0yFfPPl
qerBtRv4LHAHfcfn/y4GilPOrzSbARnZ0DX+5k/j9vhWmIg/UrF9/XJTFWb/71u2
oOMb+Acx+LDV6stOc/cH9dGLr6SWT3TuWjWZq8FAmc+0YYLcKjr1HezU5iebd9Zf
obncbsO3WdUmmZ4NbKR3nYbzdf5Fi5EgDGaD/Q6XOk07Ghoq+aiP7cZDMOG4pJ6+
vTMlkf1CE6+0d186/D6SJb29cbwDPB6pAG1NegPaB2fCAszbdbC8NFZuPDFiHCKK
KvSzCEhY8R0XEpCmDSI5+8IGPNXlYagjFuilkVht0mMholRC3FWtLufgQuUI3Nan
mFS4Dc1bIFDbeykY55OfPt94J7CiiDE8yTw7QpBCm6n8Sxsr0+HfaUrXC3wfqKnK
UDSvDp4CiixQy3bsGv3UPp4LIZiV1g3XLQphK83nTLhVJIO4mDDB2jDH79B1IXxv
d11Oz32t2dHCK1v+C/qwhYnpQvNFUdVD5lGZn7kkrfjFK/CwO+bfL1PUrayBbj1a
aTk5BKJiut7IvkT5lZBXItjpAY1XhmI8LZq2uhSlGLQViaIrppoNFVmZfRKLghut
qP0ggKz/aNA/zKfjlH3XTCLwVtXfwD4xmVBkBG0eGWYvpukTYGcISSb8INXdT3QJ
zrXB9uV3NV1xgy6rcy0yPIGxk/v8PjcCje6NKFBWOidoLh2zJvm1juQW/ZUrOC4q
fFAPaPuX9nLB22R88WF2LxWXl+ncgrMpxWxxHxLwJVyFw+VlaPmwhfKqBT2LWkH2
7rH0+I2Akq8Uw35W1AmtjCzIxemQpKnBQc6xecSx2cqtlu6O71o2nbo6nZiq57MS
/v58N+zA4d5y4TtNCyf0wX5fCfabFKGnHa9EwoJdkvPorCy80X9Ybco9YxA5TTXX
/4eowqiNPLsM016mxYDczQ4nZBQdIUt9LbSO3UFz0Pk7R+S64mKIs1ezX6sF/XFS
a3wop1UKBj26n5CDzqstdXVLA94LUnM7sKR/KUctdR9gAnMZnXzLE66Aoh16WZfe
fqtMICXpBH0wH5oV+zY5v+K6X58jBlDKrQ77sk6CdzAAALPac5bHxaCXrvK4PWFs
3Jvq8X+Z73hJT7lcvbzAPBazk+2cyPyumNf77WCDiAbKIWpq6JycFzg9D6smCmNp
USrnqBTxmtV9SXBDstXPLoT1kkXdYoyxAHIbXHws15YVE74dH9QC5plMoAFJg7UT
dy69bSDfAwQU8oDrJC2kU3SNAwNfXru0BghFnsXsuIq/ixj54as25XdaWtE4fdRJ
UPaWwanwEXVwQHsqzYM83PQiEFegTPK9wL7WLv5mSWup88jmT+ve+bCh+N2vYUym
Cn0Guuasii3zDMwtIDD0Jmx2JXiTCyEO5STw1uazi23xr3Uo9T+7dnc1frZ3pp+v
`protect end_protected