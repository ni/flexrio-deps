`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 29664 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
Z6yALt3nnSw9nTnZfQBUNdesazEaaWTJnKlG8RTtxZV2xCbiQadQf+9Z8lCidq6y
kOxhVCZKhX8hx0cAWk55hTWrV6XAvARxAMxvZFb/kI443QZ5xNcNGaA/DJuu04iM
4HQahy4o5vO5R2SbNLCWFZlhD0MPR5EoIpxiveU2lT+1fqniWBHGVQaHdeS4UYDK
faL/MiYF9u/o42WCMX5JFV2Gsi/3Mt5YUixC6s4PiqaVmNkU7ly8qrAhexRQ6j5t
6Q/GkkzkrJbFInB+DD1fUFBH/tVAGaN8fdWhVV2dKXlothQJoSWeWM1KOdA8n2eJ
dGG1H9FcUu1ACp043kpKYkmQRYADANLiiCcQ1egnrVzNtCX03ZZT/wEoaxsi8QgS
iarfsIejPjLArNy/NABBzSkTjj24FCC+2yx9G24bYG4TjpIrNcZ3di4AQRPzcGq7
p4QcbpM9JZEOyWGFQ3ZvRWcYKnkBXkBhB5hM29C8RZ9WxYKcGpf8rbH4nURza/lH
IEwgcarVW6YQFPB9LBowBzdzkZBa7cbBUp1grwZv9NO0k9oYci+cR+qKOCuwfpXe
Bv+ioUAY0gcR/9vWxe8w5ajBiwiUnJEhhxNuoaGV6G9AcITVwEM+eOxB1FVTXnbC
ViGhAdk59YGFows4+3rWxZu0X1JXNjfts6UtujxZrFmIivGrQ/r53se1twHfBl18
T3pD6ncl3y+06wpvvsNrjKpsuS7L9XVf8ysQCvpAoChCxWXYct5OgpRgVuWZQ9HY
bVsjBGyVZDGgQmBYUD3a9tChZaaSGY2FCy5U2azW52JZdq/olRn4D0MtLAuVTdki
RiFge39g4Sc1H5T4POXCnTCogpEJOlBXocDNEQLto8+1eVf0WO0xZPN9C+ZMp8Fe
p/kAPSQm9PMOD+7BJefJQBYkQ33L8sq1JfTlOFUqUgX4yfPMaZyV1EKkjlOjpYlq
3WzbvlufuKKztRS+uzP6v5ICis8gsHUsAgLfE6ROZTdosSTjdbQOgsqO7nAancjD
kdbOKPhkm5yu+jSJZ+zGxihSgybGvGfqjx0aqyDAfFFALy1U9mYbJsVlfg0KLDD4
nq5PYGJJ1n+iGsVsoKT0hcgGKEIv58J4hXESLHBxz9AW2hE4BDyoQHlhhRsjVxES
+jTA/katRguiEUo38k6vf8FYyOgiajP/UjkQ6+79ZZUOiukqb4IkjdQ0xQ4kHZSE
SbQ4HNztZXe4MasuKcfJT8AU0NEX4/QeuI8vUBYJkmg53MnzQkA1YIcLwJAFEaut
OSC8/vBHdRDeIrU+GDtxtPFT+ii46YIaBHYSkblLEIPw+oLHEw17PnwoDGAd5S0R
dH405KrKUqdxyMgQfZxRyi4uZQvT85tCcga7rw2TKkK6Hax7Q15fgiUzftT0sttp
FgtOQEiXpACbuX95Df7F3dfKVY/Gq6BAEzt9eXcqwFxitweyV5g9sjSiOavE+m4f
9+uENiaL6i1EvjBHwQ+f6gx+2L2B1pvyT6S6601PHi+pCRj18pRBRQZ2epH62cYE
HhNt47q1eOxekvkCtnfHqQ3G62054huXNIXvUwR7bSUVUzRRc6FXDqsrbqXy8ML1
EVRgqEBcTef6rdUm260yRdI8LJ1TeEff5JRbrQCng3FW9LXUsNk1JrUKM25hf3PK
VNuQVyh88U8QfKHYuX8cSMeAzSs/vV4Cuf6tTIAYsvQ9VGXaWFVAikP3RQs64ldz
F7bnQm4HPwZwd8TMMEy14Z05Pn1nwSfKN5Kl1zMvxwQdCZtKU16WZmO45Ozqr0sQ
t54M7oe+B+xNaNg8sxOpgvr2SSO3fxBcZZryML7fJmSCjdCdwmzLNw9nH0zJ6XAH
TmH4N+hZYo7nqtYA4VXv8F/NhYoQeUiNC+Rt3rSeyX0bE4gDbxlre4ba+iiYIopY
gOTFCazHP3L1PTLKoJZ3jL/PetsN9qKMBXce1MFTVMh/JSepA43naxfJs5KFk7ix
lFYn1X5QVYEXgtAdA84uJbke032DxR/MBvjTDj856HNJ5Y54BKb4FmDkVIaOy5aO
qvoZ7Y3FHBjztL3+0atSKViM7IoraEUQ7Re56Y26F5r3nmaamLkBC9D9TNPE/umq
QCfEnOh66ZUxTqbpPztC6k/CaRvCI6jjn07+86Hc1NQFwZxaU3ef866+fZ5+zb+m
mLIpBwIvrwurCblzcY8t6/zi2WbIkr0e1tW14EPzxKi98eC1XjcqJ6eHxEZJF1Uh
/49Q6CzwNZ0YjyS9tgabpHtDj+4m3ltduCTRGU/MFIoZ6CgQ0L7+lC2gEhINCHKm
oVB5bJ8QF7Y+/iehNdbNxW7oq7WVnyEOmP4LnLp4s4JkN/ykuFaFeDFjsldWxyrB
o1XdylsP8W3zXQsBU5MljtAOzVVvOlXiJ0dvJX1Z/BQOhq5hMYs/YJu5PTixINY1
jSoZp0YyDcscqTOPgIjWva5vSzNIMbYwa7niWyoZgitfNRFrG6c6KuDUzxiDpnuU
TUBEcAhcyOPwsRAHKUHUFyYcT3MPOj1hOOrUEb7k1daOiRWrr7eMXgZ3vcxWDcdj
p3noQYMauEYks7BRkjpeKvHN8cG5+766sCLAtA3GJqNkHvR8isRPGg+4kZNJnh2b
yIwk8n2JT6joJ09mcNX/5ww0qEDDQ08DLd0EWOCDOQnsIYL4OAcyPQK7kuW+knHV
L4+jZOkjNSoV8FIP2GO72kD8+PtRkt2UUwFTA3fr/M4XCc4x0EEgElLOPcHnD7+l
GQf2X21+dphLuOEE83fnLimK0TD0YHtfCjXQDNTvIUK5WpI7JaEceDDDo6PthG1Z
GEGYPf0oAADCnM25JFgW6eK039LQMY0MuxKv8gtAfGTqsEVsAsLUnoXi00HWZEOl
L4A5fF8pouKMmP3wvAd84TlIni+J1QOxqclqE2FPcfiuZmo4z2so2UHvUHMHWcPo
OKGW7+Jddxbd3VDOgkTwDwIqFWDSt8rrx2MkBg1pm3EM6231/SWY1700eb4E2bVf
ygykQa6P0k7RNQv3K7VBsG8sCRGUulaR1H3Xlqwe+YuK6H8ys/Cly//DmRKGex7m
r58tOOTLUUuxppxaJ2DyPHVT1gfvo7rkLh+nga7Luv7qxAiB0ZAMes1btVWzudtm
FZCJhAfR+iuujAybNPMaXohxnP1jsrRS3TKD6L+fcm2dLsInW5NuneAQyyCJyQXd
fUkLKNisWl+SHGFbVboo5tSbUFpanOwsKSK0zuHCN/z/aoSE7lATLzHlvdpDexMW
K2zQwfweIGOvglqntOxY9pipOz3kZF2sril6p48SrcoVNXmHiTIcAX/4UsSakNxr
u4+hhiHV23CDxt6Efuc/+KWCAst1Osl+shJ6PhcJG8LvtyG8t+ZeLBEE6CvXhkVS
/avi8poiBuFPcfuoklltrvim4yCBFPxr1fpg9lZlAs/I8Wqytza8l0o8ADhWAq68
TBzsH4Ffx4JWnI+MXsuAi9/YmvBVwIJsT/ZV4NBUOdzB74RbL6lkbc7mLEy8U77N
7P2dd3fi3V5U/bSgaKZ6CYzdFRUaueI94u383m9IWnAl0sJCRh7S/PVOFBpkfl+Q
rpgkgPXhKO2t7djz4fYS9z4mriHMtvGzrPfitnPLDsPTENjg/5rZNnWcsdEYy258
Pt5xqy11t0k7gPwgXQ4OalQOlJaVXkuyHGMDVGeG9MS+RqYQnAh/mwjwF4FvfKEr
zyAQOgMisc7W8q6wkzSB8stk7Q/b2M6hJtuYrfGlGzN98AxFwU1UdrulW44cXpZL
IX+ltc7Xw1aC8sncuIVsjOJLtKQkWgiVljnnUkU47S+EuQExCKJyxm0D9QyaQsUr
pllGzTLk1OYJU/DT6E9Q75Jt2FrN+uemiRLScN12thLTDsexfE60UTp9cNlhzTZ6
+iCA2rtAWGamH7SsGz0+n8QJ1r/LetCmcYmC/k+HHpcrkZmD5kUv7LSpikYyVoFV
1wk3IZWEbNHpGrjiHvA0TO+/TZ0zBceKlehHfQUNZu2L/WGkZ5nduw+MuAtKK2I/
2NvzV6Hr8rpnDVU2rnlZWHtIaXaAvAF/1mZmAccjwFgo4sV+SAA3mECQU8gjDNj4
90Sa+9P0XwtjJzpjY4kH/NXKFmhmxj3IuGSiHkJQ9LMoJBze11+XerF5ZC8wuetG
LNRR51u0WlHQS9tDH34ijPOi6+EtUrBG5ncnd+kw+31idAmZqWkx8c6WlWUI1IqM
tAW5Mf889dK4Bey8TI2wG6HpY6Qp4Oer5XZaE7wT/FY+nwXiz1hZfDU78+ibGxOD
YoUtLTK4KKfqrTN59B83roflzLp2saIdR8DfWCDZXUaoUHRtq61jAny6NQGm5VLu
vFMUzE30Rt/g9DhGkpMQ2qaBPdBT2T8VSSyhZMbkdmfoYVMsDxaEw7BcmO36qqcO
UEFi8BteRQdz3UU2MnZGV83c+9UvK+CVAVu6/669wQaTv4GH/P9fl/yNiQ2zuwV4
ahGFRdlAo+b4EOVRNLievF5tabNwV88681bixlUgqGYkN2A1nAT8SBjQsYDmoNoe
Brb80Hwgvc5UUAbmde7SrQyQu8QpWTYLrFLvMpu2L82u6xtXeQJXCdItaarS5erg
86PUBVNtGW23gJOubsIPQnUr1GhjogNjUtSIWA3MwsBoM3Hy5H0UgUjPHdzk+vOy
W1YAV2/h+SE3CnHsdNJqwdnybmtSXi/h/ydGjRTtdbQBm7v1cENI6GxoTvMoOGkG
oxiTvP4Vg6NGzh/NovTq43NWKCe2Di8pxMe/j/sMTpkxKMEdVrDGhr0E1IJNqfBF
3hQbDdCJShd/Ij6Pud0AR5G6RMyU0d9G6kvf79aTcZhp/i9qbmMvGGvx+b9BSQBq
hadPQ713OBuPdpSYHwfZ/WpwfPSs4N7ImBX29YBCzAgfydRVu2FKovWkzYigm7Wt
CHdF7Bco3MmaTFSdWd7EkQvHOz6dLP5e7dxWatdhHrpVo/OxO+9jTbacm/flR3NW
lmZzwuIYgoxxd1B661d9VMvFV86EXgzNPUiXzXvR1PPUbf3/IilNzhFLPj4Obp6e
f/1wlMf1whdchUKhnb1/Fz0GsL+rD6gY/qHh/dDpiCNpdVwllnA6dCZoXjsOWgIE
8PLhykZ4Ab4u3l3Fw4YvH7P6KtfBVRH3rUNPpsNmy7dWRinedW7oCtiVL9Tr9m2C
6gx5ZtdVtN2D+Q+2nchYNHm3HjjgtzuI9z5FIZbduD1FpnJwuEC+whxh+1i4tPfd
aqsnAC0G258v7VtfcnxzGtfZ2yjZ7+Fb6YZOwpJNXPWAu+fXkt0hMVpp9S9WvVfg
CAVfDbnsNwtIQ333F8GxbYWrPKrzV2BrJL4UxUG6AqXqNeMwBBa+rXHZ7oUiygvQ
f8ewr2QUq+Eqs7TwwCXuPmaW1sLSUtdoKZ8uv/qGVh1lGiNRW+ws04BW4eyqoovM
ZlxCB3Gikrt5Tg23AFRxhbgE/v6k8dfdUh59rA91oBSCAzdIRrzpdrZiykefQrmx
CJSg+6QSQHA7Fdhr0rPrUsMFX/FyIM2BczfHOYsJDV7YdsFwlNBZNyYXGf6JQFKt
TXRZYNAvl8tovBsdi+AETalpim+FYvyiQlbTh5sapU9IiDsxFWY1Z553ME6zT1cB
sPzKyo1/NKP3t3uk7/IE+lfljIi0UVw7HfdF8xH4cyJG/57sCTIDdrEccyRMLiAM
c3Tjnan83K3+2BN+mE70qlorLVkrhePeWrK4kBQPjlPpS3VRG4iRYkoS2I/Nf0qt
alVqtUfFPTn8X8sDoTv2zHVov/kvjaKKXR0bZCNuuCTTz6hK4nPahByqk2wy74T+
04vFFxwpPTC2nxP/q/sP0qj4obi+E2QglW535NYITK3FfXqCi7B+8MJ1IMPvvNLD
ieiOF5q8FXcPMC90th9K1vjtkqEwrc0AvLgvbku/16q3g6D9qzT8T1rxqQ9rWvb+
NWCEQqaEUlNG5nDd1JDvS7Y2Av4dx5/VoUkWzWszkotsrjoTPsQZAzWL8Csyxl8y
CUFjncFd+RnhoqvLbgtFkfivF4fxzOlM6SWilNfoEqEYKLObZMhvRfE9x4K1qWG1
0kUZ3PX2TaIgaCLBoH/wPqs32pcnZl8tNxDPwTP7HUDjadUdCzUYOXKy9JMxWCC3
pVlLj7a6k/67UvPeLK/2aplwCPd6ZMEhg1kzSwLM8ljdrB7raS2TMQpB5VJ9MJQp
IFJ0P166IKLdNZG3sNAMvQw8Uks29unoSykVD/DeJ01NAbmSXa+EEh5XsUsE7utc
w9KiJcN3yKnl/Y1JgiBlXKWKHCNZjrN2bcXoEE/8vPEwHoNbMChgCFXeDi1vn2VK
0WRL6EH39CrnMEq6g8qnNaahNlJEyu0IcEAFc8kPj+h3yt1VgHnAwLz88B5zruDb
AzjAFVhwAgOUc89fwygA92BARGt5j9onWzkdUEobQiJKV4cFp2xPu8BI6Krye4Pq
J5MCfTmw7Evg4w+CS2LBA3HhGLE1BmpFqHxc8QpK7d7VsurcEOA+6GJcsqNugyRw
+GQJHb5mAkEld6MU4Ubl/BGoh8ENzZnRCddFg3dAJLGc1yvwN6pfDPCQJrwlE5/u
kyH+mu5z3tlcnwvK1fO8CDtzs0b6xirwFiCzNv4uo2WTogRx93QwoP1Nze8B1fXp
dz0XjuVe5g/YALLMcm7ZjWNgVNhByxni+3FMZuA7W0Xleqgy/q0jGUy0YG92M+eR
jacjw12qCUQvaf36toAbiZYKGIAleEYfckPYN9FzLSLtgQDliRav6xyob69fVzq9
7QlBwwdc3DmIewjjWk5/WMv9JffknRkYT+kOrnnuUsEv1zcTon8GExnRX+bVYboN
r7uaglcxXk3vQdo5GzgaipnDI6J29pIDch7aGA/APcFNVOeet791G/Di2ojIhf7D
PC4iosOaTcq4VVstTwXB3xlBW/O8Zw/vUadHqD5YV2sR6n2ExQGACGLBch/OqweL
fdG71rWOHXXaQdH30m7ewC+h4DBcqG8ZA1mqpJoeormcqeaSEq7CXd8pJMxAZlV9
7rVvlAL5+/RsiNxBeb4l3TgYoXXRrBuwBvDiJRLJzqZ5Op0/MuR6oW4pzsy77YwV
rczZO6ggeg3d0/jOb+vnMxZhRj65xTPy6UFGN1oGc3jdMM+mHSv99F0IR+hHypXX
e6Akl3Mb8i67dswmENPRVupqSifrCjPppnwMyPqrabalM9IY3Dfs7619PNNqBlg6
32SNHDW/9CJ6Se4oDc9Emdnfo+q+P6XJIY1ZjSaii60AlXphxWRanQ+W8U0xtCt8
dkPH/1aVgZNEyVfc48ko0ljDvaukmr8xDLiLUpKB0KVXFpkco7K0o1z0Dd2UdhUF
cd5CJJWB4Yf0LRvynXF+RQ5hfZaNRfSoeq0HP0RB9MdD3Xrv8OBsDsdaUIcWzUxS
gv/tO2mbvLobCXdckfVgQCBRPSuqW8MGEEl4yqnlNtilqW1g6CORZZs7OwqINg4i
LvL/NXe7QB23/TgHYdQ4KJ7jA/KTSNVHvBTladBs47pZKUxpXNP654kLtrInk1bb
4m8y2ds8c/yBzWeLzv1A72lYG7F3/97QcjIFGD4+nUSrhKT97uYfTPP+yKji2X4M
5a3pshy65/Kc4d6rT0h4VXWAMom7AUtcl1YfC0A/HLi2z9iEMG1YpvibY0Exn1a1
i1R5oytAcuhE3oNr9vau4FaxCvEnji58BTS6wam6AFbsDZfWWu86+YgxcbV4hJxD
KmlBdrZm0zbmOQkb8Ml42yNeih69HUIHojJ/EesbilmBx6FwvjwOY6sq3pmPzDd2
PW47X1by5NJkGQOu2LPjNaLevK848Bk+CHutGphj25qvfQLxtpnuv9CpkYWsKxFL
atUURH+roOwsIRkTmM3PIcUnQku4a8L8XeOvSoyak7q3nvYXNRg8nOehn2wPt7dB
XkVMA3a+a76SG+6cbYPnuDju47VObs+7gEEyL1NDvzA6uERFldMot+Hcnd5LacBB
bwigyu5oVRzOT0nBrtrNWGLcISIaxe1QtwlcTICy2AZiLVt+H7qFVXfFwzUEu6xt
CuM2XXzDwvKNYVi8UK9rNhnRmYzSkvFWJZJrPLsiqm/pSJBwcKihVec3u1MaVl4d
X2wfQcYMIVcQqy9hhGzpX/Nd3rxvtoEe/PIDR141hi/7dWso3SnbFZiDV6QnI+8v
yXjsF3oWxgjCJHx5RUunFgZiSvaIdclt2SZgM88s88tJP6izPs3NoMfYQlAVhvyS
6od6dXsLQQziR+EgpEwNXMTVnM8v0APu3sbXjEmUsiBEtFmQGVsiec82rJhCDvHP
ttaVHHhoXWI5PlCeXovdQYLt3kjj/f2FS26gCxmY/po8s3nT9OfHbKe7Dra2sac8
GS7Tm60FlSTGEfyyZG9g1it/xMKAWYRyX4ByKkKJJctejWLWDxRj4fvnQvJ4NFmg
PhgPTCJcNiSs64UKTFDVzAId5ecutzyb3VlkI2Dtd2z1GY8PLA7fw12S+UaEF7HN
q4bu6hvoeNlvP72580a6AA/2m/uFzzTXegvplv3yo4Wu0a+p7L6+459HUMLEsD5s
Ki8cn+QvMzUYt/LAp+xXXfVPf7oNXY/rWdFk0ZuA2fb4Gd9E17mjvFL9Sm3C9fGK
aO7ZcXdkp/3Kcu8TfICqOvqJUVga9AB6TeClYrJUn6NX2UUQUzZrSlMErtaINABT
ZSBqMEKuSkEmacczsbOEs47oUtznZ68ntevmd7HdVCUR58jwtgxV7UwKc/6+iSF2
n1DyzkT3CeHJNSEAc2MT4GCTnW7UXJep3O2W1E8eyBOM4h5J7Mox73UC3QJiF8WI
B8inmKe2KjOb+zQZNCPD9r/MDbuTXlGzImLDtGb6RJaCUaD+eIuSFwzY1jJCOdLo
h+sG4bwXEWBYT751ZinRro5hn/iTj+Y5prRmt5uT0rkmFjrUklfUaUrQBR26UCnM
xYTtK8/GXeapEFt6ZDbZNY/1T0LZlGd8hIZx+q760PtY3L1irt5lsTuFvqp0QMH9
IEhQ7wsbkdtfXNQKZtJfBzexBBZNObCeU40oN7hHogXiaXVxi9rwWpBybyFILvuv
xmqQgD6z0FuGrOH0lLBttnqDcD+H0qAiQkfBfxsfmmKxZz/+aIddnDMizdPDnw6B
es8Jb6gGbFFHm2BhocdIeN537EMLZ2KxFo8sUve12/7sVXll0BEkp8BH1Tl11rcb
DFXKHPlpVRgPw42dWOhZND3vuK6d6Mq9EJ8HY3/+nN8kB+r5AXO+fEvbXlCUymrG
Ecep+VlFFR6GxD3MsnFsjZV8/2OKMVd+paHzLJPJRn7cMqVhbISSKAgtkztjV9tC
RErJSCa/9SHwYHY6HB3u9DcD4igbs0YLorgoVaLUOQzImqSYbbU91URvC+tzdU07
KyDWrwwvYhl9AJ+kjSL90OgBMyDPYF6WgtCHxqyJUMYml1BiCzKDJbxvoL6pgw8L
983ZeldYoXP5NJxYPwvwCWDT65MnGMyx2PvjrtPBt1ZaetH2bwln+BKV0i27O8P+
pQq67Ls6hoxkQrTJWBUb9DkqQzREc3nwsaiN1gVgRUb3D+RJqhjhBUDdtV1LWeE6
9Hvhg1vAs5TydF34hdpnLYV2RdLanygOSfKpGcVRudO70TWjCpIIFDnhzIocBZsE
V0Oy5LJ5uQ5p4+tzO/Equs1fXlRRk3DgvB6aKgjAKesVFsQNRNjOQ9fLNEcSt4lz
qdPe+SJ+CbLjlvcr0FPgLnH0s9z9JpJW5Xs/Z/A1YCs4H0pvnpuHCPkxL644hvV9
qgy5K9tqegNO1JoitkfMULTZzRZ8u4BJHukCUPQ1JM9inddDUy2IOiu7AwhWgn5J
UP2UFbXBfPwaVF/Bn7+K5lqws0xrGHyw+ETH0n+xEx29kUjPISHMJtjH3eScn7Qb
nk3lXKOyrbQDhS3FH1ecspl2naNfeUfKYoiPXomVyC+/3Ki6kCp7/uiVQht8+HX9
SvHcsmebppHsUNR3x5Xs+J0gnoU4i4nAlNGwZzVB4oA6pceua3CheztutPSE9vyN
gyM7kOEvFKOSQ8hmUd6hVCr6DP2h6qLudCGDpjSl9xcRS8yizaT2xv0oJwLSbdy/
Ph/0vmy3C7yxI48Cie3DJVpvVwozZc0ELBxIcg5icNV2gNgwZkmhO9TGrZ4yP/G6
YMgOyx06Lwh9haNG08fQfu6eltrVfdXQ7hBlT3rUHgw4imGbUQyYI1yvkPF+lBMb
Q4j979kd2RK9HKPLpFs0oe++9wv5bXQOf/p/9AS7PYV/ilbSJTqqc6s/Y6D2EwOG
Vqrmqa5e9/DVSWCKyfqK1rmkQM8THm22KUs/X3PPkzWkztjrYbxlNu5ZO+amdnXp
n1+NkblVXpIx1M5egms4VslXJSroaq+a4/J3N5iN8z+V7mVaoXnMmT6Y+iNkyk3g
ZjZPS/41Qg6Lrit+WE0H3KQRykazytdR9kc3t8j7Lh67tLjrY2/eCz9krO/tYUjj
u83MPRtwuDBUCQmnPjCTusoYd/Y6RFduNJ+MInvYw/JMmiSDB4Ps3sa1Gu8kptA2
F9UqNg/m+CbqwhxPqrG/4mPDoCVkaPtwm5ae5o3ltyPkqKoJ5dqiNRvebjx+t9OX
2/C3ksJFNBh/e9sBtWHbpwp1lWfhRhLGiZc7ur1+P/sGmxBEzbigARSm1yw4IEqQ
AAzio1omyZvbopOY59r++G+AnPF0tJVLZPkpNc5OBQ/BAHPi9dQsxak/MNE1Sanp
BZ4D5Y1tPmzkh4ObJTQnehHIEQF8hEsUx7kzzcy6WopQ6DMkAWjEuRz3AAdpsr6I
Co7csF3OTebDv/Dfs0cdg68MBimJR0qWeJPFoX9hZ+N8fGgeH/Ep7OlpOvWilTg7
3HmlhC/nlM4Kj3ohQFSH69fsbGdhChYktOXdbHv5yYmCJF2NqO78WSKl87jSkcQ8
yJfNyDCHel032S0GJHkDjNwQDnWd3wtvih6/7Wd/E0r34jNsMk++VaHJbheRE4xU
05xE2oZmG0o6mGsA/bRwC0Jass2vTYpnNo0lh1975tQUttJPn7qoWrl5/CL91Uc8
oVX0YAmz60cz1WMRHgf7pP6/8W0JBjjHL6wObhKs2Fgg9/zAoHDvDz3wUyC3Qh82
L0/EUbqWy5hpoWHfco2Fu4CB93vmj2v+/B1gDVeebTyFuOA7oa/wEqFE0sMqKIpQ
3AmPkCXxVLgRXYo02TbNL11vbwViloSbMWe2UYdVODB+8h7wcZuy5Z5dN0/d3uCd
vqeSNo7OZtcAwE4v3+dIvA70qoUUB8vjIpnlku5Ad63QIEVKPAg5sdVHERTcLBPe
tlUjCeU4+bNXmO4BBgyo1vBSAAd6b4E1AsZd809qy4QIur3t1vD6+whnzZzajFAn
XXDUvpqkwUBTPbiRMkrWwTUFk/8GRSbpxONrsbNjHRA1rsUrp/WOz8pK3CFm3bNP
tbSwZrxu9nkghH0zuBGzqi4bvU9NuCkXB5CqnD5m718VSpTJ1RMf2nUzWU10VimT
H+e4DFtmUwwoDZ+H4VmhaTRC9HXI+6G23fEyRkTkiCGVcmKQP03QC/h++dg7G6ir
Szpo5ge/0hWemtzYpNllq9OfQOo7mi5rZUu2tcBOv4/5MJhe1ut0lQB/v/bH79Vv
BKDMQJzJ35Sy0sEbfsQa8hQOsspKYHXRUxT/vueMYy/Y4wzSWf/4rUdMGc9MPJYZ
opgTMLlCfVeg0Ggc064CYGei0PXdSDqaOO/XgIfdAQ6WbapOV0AmvaJQYZZwXAog
us23CXjk60W6D8H4JAfp+5Mz2JjEuEUfs+KibVk8rff59dCfSgGAu9WBc8KQD5nG
jJa9AY0p59lkVS+1WLK8y/Pt8LD0If11ONHgf/qMVTZSsY2/0Bq3njSmgBTyU/8y
uEXtgfg7+gQi2+mmVfMO2MsxlBj+QFDpA7aWlJ3Imhv2r16cN+jt5GT4as8yhVrj
wsRpufeCM/fi2v+3w9NQgdxwnIRyijuGsthIDfEW+gJfTHhzyr6vZ3m343BACLoU
e2D2nPEbdokQSSgSyAKo50Bc0E7Iw6Ko61fk+PxZi0cZzc4F5+14cc0dZL8ClGAi
rX28WEemol0+10dUeQ1Bg3ZrTJAf1e4zvOa8JqaD8Yl5smDPN3jLejWShs6Ae7WB
wOmBiO7yqzLd0S2gl8D1LGiuP/oEAQD0rdJ9xTTv7nY/dfNpW70Hik2KUndsaIQp
vg40F9+qTDseqD6QHgiSXaEPte58KuHYTTN7nNxZ3dlhPEgSLBHZx5AkSwBju7VC
6T6jx0SeOitCs6jswRTu2EEw17sj9DqxsN3GgQjOUeU4BCc9As5Rs+iFUQj9zIa5
1XnleL8BdLoAx8zIWl5XwvCdUxHKw47FOSdRvXsf+3Vs68XS2X3suxYfA27M8aiR
nhGCoz+7OAZtiTHHyL6NUWcRlNLDJMN7lsVK4UooGYEoOU5L4idmfff8cmBuA+I6
0NEsIQkSXKIERKj5dk4IqbzVogx/dgl+83ftHgroYsrjNew/NwXWfy1dimIDIhmV
aldt0VM4AInX+yC0c6LSPSYnqFh6MmemtiIJyEMM8dyaOJiUJ7SLT0NcI/j+A6MT
hlmnxtWy23xDC6jow/Inv8MwG0FNMq3D3BJfsOcVNslWOEre41WDyfUw0HATpW23
91xi6xVfELFNoIeCKgmDjoF1AVp2jBxnxmtPC9XD6u1FobM/Pa5Gi41zZlNjsvhl
fqa8bWXgu135iOQ3Y8nnOnEcWXUrcL82DPy7+rn9zeeNtPJdkqh2SmojmAfu2gS6
NJc+ibAkYTQ0+cWkQITW9jxIF1JBoStcVYEByt2efiOHC1lP5TkdodCatGX4NvEf
Y2gqweUi+ie4H0Wz8gSXo/jyiEFhYd3pG/WeT2G0w8eTWkK080kgFA0ANCJi/eeK
xG90+p3xh6CHsDD1cu1XY/fSN0emJk8WuEVHasH3dA3VG8KOv1yNdb/DYLaifeOr
otKFvNlswB1RiwwKIUIEeMZb4mU+JuLmDAWqSTgT4l0vZRPqELzO29Op9TrTeiLf
HczWbT6/J5zCjiJ0KY4cw2kwYc8CMNSGAyRI6+J5v8gkAzBRb0/osmdcKZ5XcIdt
SUbLM25sizpiibjb3WObLLx5oE4cRXvBZzOYQeI3wEuzKkUMTvBe5KVD0Lh6Xy6I
iLpfSFVH1ORvyHTAMNFzb7oTZZaMTXhLzTrAO6BhZRBRUQIgdQNvXgCDLssdQt6L
Gpvx/TaJsliKG+Lu7KwgZ5JdbfbhQPKVpulzphV5S0v+YF1xNzztvIhsVC3+ZA+G
ADGPUcVH9xs6YAes9waX6x89KuLO2DtDfyUBRrQST/xkB5zcVCM2dxVMn6aOXNv2
6nIGQfP0t1tAUIlWxh0Qr9cKNKIuhjYpUABQga4FOjipoesnFPvNCvAW+5LMpqlq
QubL3Ql2C3kVUde312fG/T8quvg4c8DXiS+Cp/B/pdCUgatCWIkrpCjQloqVHUGb
hBhBwdRMGWaVwdAum8HZCgLdLoo0TidHLgDQZMVo8t5aSpjNa3qW28WvtMiXvhQk
tjiMIlJSNR7snDVOTwrgxqS79kpOSysiGzXa1qFouAgcM1V9OwiJLviEWJe9QcOv
P8HNMCDCSMmaj64SkC75DGF2gFVuv+cW9bF5V+igj7MByzfc8Oo3SC0ck0LfgLQ1
7tVFjIrJB+qzXfcf7k0DJZWnb4DDuQKj9HMO+VbzcOZcwtNa0+5h80N2KBTHnL+A
3Znrz9Q2mO25QsxKJU4Du1myTzIFrEWdp5xVthivOpfNyJWONgpvV8POvOTzGnIr
1iZ+th5/YNFM7u9+mDILxTpMQaMlaR9ZAwItJPp+4VdCm6KrKvji28Y17iWWZeGJ
y2YfEOfHeQ+fTDK667avPywWnQGPwfRxjveLFIRX/fowIvHqvVepih5Un4zLiGNb
RADsIdTH1xidG79HO85xDqEXlgSzbPXEzB47vokReiPpAJMw1oYuMk7zC4djsHQ/
n4YsTUCWji5zzADVk14Pije2cgpEnRbDRyraxJfeoF+CbiOwKcN2KtWtfiFx3bpg
HycJwAneh/eeRAzSxV5OIzBpkjXFT+N1eIMV3A9kjBD2ECPJoU4M+3IbiIpNAhs/
mnMnBaWUNOrHP0oBXfsi0RPoj5Q2+H458gGmGgIcJQhD6H49tGv2V864/vHtc8yk
DWE+PjvSz9jOp7mlbeD5OlxDhZZtLhH3m/z7KaXnPPIaXSoekta07tyZAfBLHGqy
mhfAOyJ06uAR07v23BMSE+/+rq/s+Y2nqsJXcUNOiSpW9WUA43syz9utkWoDS8ry
XAnezQTOUcPuclKrpT6ot5Jbe/b/ek9nbbzS/5PRiH26TzIU/suPSVlBRWM2Ma5I
gbXapd6nQQt7EIne3c2YitkINUMnn3M+lx2RanomtQxP25E2pgKfonndI2MCl66M
i41FzlFTjaJm6t/ydvWKW8RG3+0h9aUVBHsRfPR0GrJsXs0eTyZj7TgEuICoqfYg
hxjIvPvDLYQFVaxjpBTrOqjtzsxkD47qmap5goOmxggFjwTG54B3oiGoCNPm3oJR
8iRAfqhPIaP+lu3MeTQC3PrbpofUSBrsaL4VLEH5b7FNCSTTV52HWYeVXR9VH4Gh
I/k/SM1Osf9v55/tPwd6awMCzq646kVIuvHluorNXcQJZLiXJIBuANjXIg0Cz8l4
lJPUFtOaGNUn+XLQPFdFZKT71faMDi9o5ZsnP/n8jcKsuD40jSXR0TMAfoXJuiq3
ZUicx55vmjrelYgPhjr7vW+0z48Hf4jPW1gCyFSTgC7ZohO3EezqXzhRlgWiSV26
TOFUEY4qtIjxIv6P4jb1P5lVz8rxxgMk6xR+Gy1xt/xFlJLgSyJPkcjQ0n3O/OQ0
qIk9W1aEIKLhj3wg5weFFHjE+jlGygeRs9dNSm1Vg5YNskO6mZ0GMKU0UfV2nJlJ
jGxmmLvarNENjwL/iD6iX4vtKrx3kgliXSXrE4vNTnGwpbRbvdMiFVOMd5Sv7D+9
C/wcMmkwY7VD0HZSFY2RGmPaPU19QBq3X/bJySaMb2baWZJPLE24kOHl13sb4NDR
cFAXGhMLMwx8rn0H1si148XDH1dN5VBQJUlOjsvstBao5ni67P1k0+xD3NMFysFf
QlMhv+zVFS0sVy4FV54yrYWMG9ij8v4tKvpctiJd5ZKQTcIY/T2AhHLQ1Cy4JKWG
fzlVUTqHruf0x2gCwYINdDrFR/M6cafEWVd+Ej1QM39ADTqOk1PLvvNt/owGGjww
k6Dviw1o/9V8KHgynC2EWVlZaB5StiJ6D1/8cGjgFF8xdqz/05oGkcAy6v9LxtG2
SIHIN0kKWSFPc4TyDUNK06gkuN77drEkpuqzcBo2RrZLUoFM9pfcHMOXwW0LUVLN
ABoZQmXpHQtD3OnzyvTmTyPEmmVDtuV7nW6ZhA3TGlou/+htlDu8PJEqjAvyTFgt
xQjNONYIUCSC2cwoJHNfS+NkJVHCfyNs4To1Pw6t3tvttO4rl9iMkfnsq0URa/lp
uQeUZ2tO6fjp9KAK2hItVeWgSihrbryumKeBqUoRwyNMdSWZ1GlUy4s/ajgVjbP/
17sU0rMrPjjYL8hqkkDV+UGiBs5/heCQ54QeMVDKwpoOeyidx6LpuTOKJ8+iQzTJ
70Sise+ct6x1l4VooHrs3RUvC3Vi/g5kzs5Kj+zyWZcPuHo1R0ovoy8rpwMBkuKV
uvA3gt9RqB2dyJGheZjeus4h4MmsKmzAfXKhu/9HocNAAmVhhbVPG182ZinWzngV
nlM3oQVfcO5ASFqYzpjvzEV5oW94YQ4Sr4kcfWZxMwP7KPF67fSzYSNpxgtqDHf5
sz0QmDkBNGSVJoVBmBmh+onAVhBP/D2V5cMv5qk3bx0fzHmKjBFuNxCMiGXjLMup
OxoQvLb+mN4O87yLEECZLtggLrVCmJnF/zvaO+hY+2dTbHHJFSxQlQ84EB79Zfoi
LynetNZs5H+qutZoKnxbCPHugfDHQ63wA0Cxt1mMWXSxzxLfYI6xPJTUa74MBI8z
fY4mDonjEfXPGoQfO6PyTf1EDvp0IaJhNd9GqcJHRxuPoz8DHt74tZFqxhTz1Yzs
928S6KxTrrnuqA0XA6eZvl7rHj5qOknjLepZkYjgqQFM4aq9sxHmhZwLpJVFes51
1sGNT6j47dm8Z5ERRVwQzUsbGlpmB3xJ4/Jra87rZ3D/WxPMLagWBlkc4QizMfio
JJN4vzLlLup8obWyxtAFY895+UK7XOy3U3rZjKM3FgYMVlXxMf2u0dAqC6Buqp+y
viuj+UlE9EoIiHTa02aZ/Msgo06cUZXFgvEjbyQFz/uv5Kdk1oRL/JXBTwKh90j2
eT1HbqVoEwZrRfnPmHILpxUtGnDxRDr7+jG5LKpuMLQJtj1e3+m8oZsm4LleZ1Un
QT2XX44gPBmaohR9Up2FwQ3nvic4K6RnT5EAJu8nrMBRUpwXYAXXCN3VTALhYe5y
o5dOMpih5ff/TQ/iTXHNsZoGTsUL7t9YbvKayYeUpvkn2rRVqq6uWNNqdVDo+EHP
KVYRsAcQvAuXZ/eGlfLFmXjtFm7Kds4ymPPObNKujp5MfGkpsfoHAJLY6my34vdv
20C+ywoIQtwS2BeHJSJDWayw5Xi5WKet83rx8RLRt0wz+lL1kF5ipFj5afEww5iG
EYLBUDOr8LaLIkhClDCCB68lt6ogyhNhBo/Cnb/54QfMTMHYjnDAoIh4eTbCDsWv
IO20NXqvc5+kFCOwH0FxbSm6hH4xv7Rq1VtDwY21wT+tEgJ3LdJjZMb+ETnUDFxJ
068HLw1vdJBJiagCckguibqseNWp2SloFXWPmyrgbe1+codA23VFntS+74VBlWvh
EvFQbqGwe8i5HuftWIK+1xeadYoWIHziM02xqA73a11RrBg6z/3GWBUIQYyF+/dm
S928eKLrVzVUeFk06vYHKsEaYCbS0qOGojmcqX0Lzu+gKQ1jFLlkn6Yw30QXvwMJ
M60fQrkCyd3Z2b9wHEW2hFNv9FZywInOSe6AzLYIIGKdb/qVAXbEwvhbvpeUHvuf
QEkkWXnd/MMlyaPPQ2/Wz3XfTKG79Cuagf5twpfy7cTMf0UtaYDoeLW+H9soR1Qg
Vbm4Zq+CVc4RIxGTRSregZeWoSZrpO17KPBPUje5vi34OL+oWbSr8kHIfd+8LNI2
Lv6vq6vSmv+aBalcmWpEYA93+E/HIIJTT8BUk2wadShrfaBISUfQF+7v0mC0JJEm
FSRZvbxMcwMx76m68sMpUARMZgVtlE9b4VHQLU9169tZRTVHIHT6lAXlY9ajP6ZV
q0b15fE2uJ/17PagSfcadOiVUQhhXhuLCi4LJaRjpPaLttoslVEa2khp0GEceVkS
lGSC+pkwo0uG+h+kMnRcic47xVF/oZjREC86fSskLTKxb9uXamKxFgDwWVRpMpoX
sgHHBsOG40FuFVMljocC3npXmaqoTMH4ZbIOC/NoQIM7lsaFVMk8Fm7UPjlmH+Gp
pGwnwOuZckewXd9bIpNoTESX+WKav7YzQJ2SYyvxnb8HTuNdDwyM2XY2V3hryhzI
wAIvIoTO3HL6+HmHlOUIYGQk2j6jLxfChStbcLODcDzvsG1LRRrmiT0Uttz1yo8Y
NIPqJds4evNij1A+4svRZidP7qHsy0WTlDw+DTfmhO9Bv6zhxFt2+p4tAxmFpSmG
/dNxpa2ApOsfYF2gQ1++BEI0lNtoXjcdnWMtxzfQNtk7uyFBYZ1aFQgtJZOnoEZv
CP7o3y4m6Y2KNtSVqldxMDF6W1LmQJm/IFiC6ww6+MOixjRyMOl2UK5BhqFKM4T2
ktp+6VR5Awao7Gkdo7pyub5oALQEy+yCcSdS7Ux8IWmYfsnneuzxWis7SCvXIDeh
GnGb2nvc6ex9PLZ3CALyVhp+crnm6A0X8frepu5Wk2QRGkjwaa/IE4KpdyIOWfAR
6fwWjE6pzx0Cdp7TJDQsw7txNSTSFTIp/xtfeJkDpk9aLKCxVg4rc5tT+AT4Cpcw
g5BiiW7lAEsV1zTRZRmmFbVKUGBHmooAG4uF+G4V6yxA5HexKd0L3N+XUY9KJAno
iw3rPv18WIB4WoBXS2rkTIOkGk5stgEvlBNAtgb2HLQ+q7L9w/rulvFvVRWbJIv1
5eggkD4PlInj5C9jJUnaVRfFtg16snEIk1xJPuyJpBXD9FEQunX9xbcjrc0DIbEX
AF2zuryarlGrP6G9wa+5cpJywS4F0Fak7JwU4YFict6vR2UhESa76MCHWxdH0Dr+
Aweo1ZXbvvHHVXymeMByfqA5PtwF9MQ2yyJA/lI+GpV0ynAm/ZA2lunoSydmJKcg
YSAjcOkYkJlVci+Wqfwtv5b6bIqpDVn6pErGCYTVxH/u4jlVagPkNqaIfpGBj0dw
BRUCJHJ5/zqjesT9nujxzX+9Y4MDNGYR/to5oKr/kycZ2o52Qkh97b16VQjqfMpz
dudM8Kw/Xh6lComZtqeeV+p9+y3o3CMZHDnJKKW1uodn4/y8Tg1c7mHvGt70NX1O
6fUsB4CIIW/UrTzeOq1oKmeaaql4DN1fhnQ5e62nQL/oX1U29kIFi0UlGlQ0B3r9
BAvpOeNjWldVBDpI5CurP/5avMfOH51n/5Z4s3ydZhgv1rbAC2pJJ1Iqy4pn5fIE
w4kJjJ11LJJm3//yuFIfNFrZLNT7DydnSu056x2agw6YtrRQ79sI6D1e9DbDN9xO
jnBbeDSdh/u/C6Ehn20lxG0ayCm5u94bPKE4Mdgag5yyMkxv+x/2NHAID8ez8T+V
vpQUMWjPqukQr2X9wNqhFsVEB9nzsyCiPMjZAywdG8WZV/GY1hxaX5akIfu8WIKE
g1s1wsNnquVyqs2rTU3+UoZuHASW3PHfgcEzav4kR99KRsZ/jtIG4pw+NkpgqVRu
D/XZ1GTJ5As5ryo7FfNGgTE0r0jyfOupHqG9NRzQk3I0gq0ZNtSvYJMdpkk3MMWj
C8JJHWDyJ/Dj/tuuBiFsuXBf4ePZ+63u4hMuypbMb/r8et9PknyywPVD/W08g2Kg
PLTw9/NSqQocez3kxLOPxbqbfKkUrSupcwfRJALRjB+QtyKn4vutIvTzSIq0AYG1
zIbIvFLFoyrF3I7OH2oOpswXLTJC/i0EEKgnIl7FgGrbyRwauGeWXIAla2TaKly0
WJNabJw93Ri4vnltclPMVObDXFY3SnZMK885NGkfJ/NKXLWdHDgoT9JHuIL7tdkZ
hyIYo2faWQR9Oa5je8DRfk+wRgH3Z3x7Ls8okn4flP6XEP9GHUQLLKM7snO4a660
EiUuXZTRNMWHqLq8LiV+CewPTSpC6ZnVV8aFn4aDv3soYSLuWAumwLk9RvtHXZWy
lCyyOgBJUEIIVHTsYTbTRBRhzWsrtw774hznbz1bZZXXHvV121+2Irofn+Q94SRB
uj0L6GhMVU3xCWc2ROOY74CwVcOUwDklsZKk+oa1V/qWh6mnr8d46LI5KZKDuf0D
6ZOi7zR92fvbzV7yQpB/xs4i/L8pEO5CUh/ihjE3ypMao+im0VZbKEVkQfMjSO+X
fl4pQIr5fpRjmwmf8DYGeymDiCviD7XB/MFvVPw7SH+x55G3tWI38sQcqy5Z2p4P
WIyw7aw7Cpr3lKbvWAb4QHWY/C0cT7iBkfMOgwJH4/z7vf4Lo2Q8k9jZGRI5OkKS
6p7vnfnAbqRm8tUB0hg8tZYpwR0OZZ3nca+yQSx1Dgyr+bBAmLVBJW1cMv0Dg+5L
e3W2J88phG83fW3yCgKREAMqSxR6QyupkjPNcR6/Y0IO7x/4CeuBkNr4g8faV0xh
tVeEeNzGITgwSLpSrwaE6+OrqaRNFOtra0UEPqDKV6Q7IQAT/xy4wqtHgW9P931j
YMg4rfamGyWOPJkc6kYimb/PGiXjLMstCz6vHgJ44+r04fcXka0RCM70cBs6w+MB
gSfC8MZqU3Ajb9KoBhL4EXMJpWNB2uG2Nh2BM2vPpQ1g6Au4aNsIpEYQKv08ZP4Q
utl2qqVjoAvUsN9iJXY/zK3fxaI9yJcnb36A8kUV/bDd0P2fIq/GzOhpH41tmxOC
2DyXpRFol/1nULkXj1PriXPKv1categgC7cNVrZ7ow9k6+ihC/Ss3nCfU6mUhxod
VQ7prywQgPucqhqaJX/mN+sQNnLArL9HJIi+aQigFQjF/63BKoYWgY9xxirYiMRg
ovgzWUB8AqN86X/DtxaXYJrJyZOcXhcYGbRytJQhDyUbNmrUhSyTWe4ErtvLvAp9
oEdILLhBpEFWtHM4cv+18asP0G8RuNB70drM8ZvBpqKDdlRo17f8d3a6CPk2T+aO
shqHqLRlR61HKJpNSbfoDjNMfrG2CUwt9ZnWB+zumXMe7IvZ6L7ia8EC65NozjEe
KUXstq7d13adGFPkTg5af3QSjXurDJH8EDfzULopV4WmEwt2DiT3Z3ulsvaegAoS
27QKFUKIgZMH0hHpuMm2iInl3GXbS8oBQrGr+4gnShzNzN8F4okMS/Wg/M3s1bbF
ZwNKHLBrIGNVgEIbYGWX8g7zEinvTk4ayYUE0/D1WJY8W/r2f0xAna2C9c5OCAXW
5i3vxlOSuO5eN5z8D1l3BL9ZbsHgDxVcY7+LJXNBjqiS3uZmkWC6oKCORF2XWsb8
lNhaBDgRMaaIQ5KQn2wJaysM1Y78cUVrpdime5JkTGIIM3P+TfzQbDN76E/4ZaxE
C65jL01VOE6Tny2KH2JXu26Sfn32bPegSmqiw538pTEof15jQTlvv+uHKMRrPZug
yXwXGlUHmmbkYGFwCmK7pvjhZsUHqVvsPcDOFVIjD0A+bqHdbyAnueCa2qLOAxKc
4XCEO+mG2E5G04bcCs1F2eZfFlGeBouvgObWV3n605Q6ZRT7ydQxI6WKaEGMZ31O
58FWGz/JDAH49CnfjbxBFsFNZQNS376+pKxLv1DLHXV3c0qPI7aNfI1m9BmHD+aa
eml7iuPMBm06J/15TdErTxIbPQTFjDnB4ir0POnkI44hbynn5/VNjuzFww4vrqEm
MmAUo0iSpnvvGJKmxJdKC5txKbCCAlFuFaLiP7cf7AyVxYOC68/N4g/rbD40O91u
CjvEhmYXuYr+efg+LzTdpdRXNX9wCJ/h0hXg6dKQ9EZYCYfVMUAmTy3cs28ZVCjw
BIQ99EIyU4zkaRvSFLLceBsyhG5zx0YvqATNJnyoDRqChLv3x7zSdC89BM2RX0Ox
vUek7Zj24mafoBysO0YtRt2jM+piNWF4ruaBI355PPHv9Me0bXpaZmPeA8pWDNEM
Aag5eIDvmX+IPo1i6Zw+qijhJjjmAgarr5FfFPjevQKswIXDZCC1GFbDiX+AxiIg
sy9CT5/vS9wx1ZUEeE6mOPIHhrERmtTdwNikvRWYpu9318vzWONSOk8xp0uolWN8
5WNn49lwJpRXweL4TS/b1mWMTNhfi1sJ6avHj0F2FxGAFS0vs9J6nXXQDuZrF378
ribsE5PQuNH70PWiXFBApt/KZ5ClQneyB77Mqhnwy+97T46XWK6kC9od4mB4n5w4
zRuG2A1+n5PGc5WVbNJkJJV8PUK6BhaJixp0pQc2GYoB5wLHxk0JarQLhvq1A5jP
RoFmwWeHo3ceH4lhmRyJ+njBJmX9YJ6H4wjmjIZccktSnDDO03huY5+gHXQmZRPw
8aA8SPiOm+WqrNW7Yv2om7ZnvfsouWIjhNPNpq4qQOOh47MAmH5oFGg/6gmrLQ27
Hjeh75UcPcIVgD3Bci2k6RY7Mo+ZaKxI84tURNRaPcLZQmw87tuaEqO16B0o5UDa
SdlSlLnxp5Y5yAV0tssl8I4MiG5BJgQgzk2XI2uh/P4xBZocrK0PzqCVUlBanz95
Ly/bZSKipw+6Fw9ZUpdh9RvezDDf0+h6v8TUBKAHe6o3xvRz8KrTQbxsIlI1/4yG
LZJHUuZWl8GkMdp1NzuimRsy/Z23D2k6A6HikFn51kbk77ZsHkzqqgZ7g2TpXcHP
C9r4XszHQSlHc+pP3lql2qzAfMIlYUweKYch2MTBFomShPvagqirCNckPfm5wB9y
1ru50qfw6Y6nViq9E21pqlY7maC6X5rcAuDZ4qv/1zNgn1J1hqHI5NrZn/9XCVAt
tPmn3J20/Hg0LlzB+fdI+4Gmb6CIZA4DzA3OQKV9RRaWWDVB8KlnCG8K0oKNn/Jr
XB3Lj+iW/kHrvG4P8DBhoNEHm5cpx4XWoc16tgD14F3o7xr49IagQnUsBcWkKVno
X5OGukOV+aWOyqfIzFM/88zzke7THP2N1TG/CwvKdxIbHHpOUPYL8OF8VSzJFrv0
OcOGllWBsXgbep62/8752TLBwswovAVPp4r4h/rwN4MNIBdXyd4JmQcmMBtQ7G35
Wl5EzIJt8/uv0C6+DTm3Y73nHXAvEtBhMNWob/KO1szORM1l7u46r+Ar7XaWXZ2M
VBVbn4jVbqBoxXxTCKCkMEn2Tp21NXv1M2NAm/veaqOcDWhK+jd0Ru5OiVKxq50A
k+syoJSD1yWfXsbbF+fiTBf0Vg/OnDMOQsvvaPBQUpiI42ElDaC4/x64DeTND40G
fy+MIquCaQCt5Wo/Or9LcBlSjLqwc7vjlM2kjv8oxB35oRRXwTMsywS/HmE9kQ29
UXKa5Kbiz8SpIxYGutDPIgvUIbuRvCL+dqACQoQ2Q+T3N6Aw4T/m0ihmdV08K7X0
0Hp0/r7GaP3ECjX3MbEpQAyC0wiihJ2EDnhheDjVKeLwEKwmhUL/P6gbw1ud4V3j
LoPPk/EwpcOBqkVYc6hPcMUKVC7tHeiV4vKBiuB5kcD3p2opMgUJT3C2qQS1rt8m
dPk523oVykvckQZydQgUXlDDsr35djB+F5CyKoY0b7mlC4Ism5UeVnChrfgk07ho
rJk7DAra8LEOJID8r/UAhuVedvkbSma27P72YbwgT9zBRC/cSolHYKUlGiTpebTU
velHEW9R3y11duKmscBuJKUkPk9BSOg4DcfSR7qtCqh6ePgZL3UWnSC/mL6oxGM5
0F0bEzLXLQXo5v7VOHWvGmpuN3FOHBKMc5ZoX5368qDS9JJZktCaQPFLUbvDNk9d
nGbSaAyzu46iLheeJZAvmA9ZbKJxYJjtqWv3vMmx2xa0Sc/dUW6isAiFnEEcIGjE
UJiUv/iLZL86W7abmqvQnoaoerK3/Woqbhjqtz/vySGb2I+1p7eXNrh34oFVcZ4w
9dMDHsbn1jmcDJ9v+ci3tVQEUcZuwcEsUDXLR73UDfnd+OPZKL4aAkoixOWdNTFq
i/a0SqF6lHPl/vsl3ti3qaB6yWDAlSw0zGUBVQ4lMpqNzTHEGXiTkojJDhyMMhdy
U0J20/u5xu8+JRR6tlSheX4bAShJVgYWO3d6qz+w0TLFIBuLxmvR3/VWCo/EYgHP
VenILJq7XLLZcmgqVdVmwlkAhprGW+XPz4myxNFxfFfsSOxcVi82L6L7X1eCEKB6
i8aR5gZRkysk4+sAgqYKZXoaBjWQikmxGqBaS37C9voO3DhFDP83tJvAJbozrPUj
4dhzWwXO2oNg+mH3q0omgcFaM2kQSPOxLBMWZ1lZNYhCSWcF+o7jRUCMv7vrdnoQ
1Hl2rDGhxrkGhfByC671terAXvgu8HbIkXyzG45geysQ5HJXqUcuIeKnWo16LbAG
aru7khXZ3hWhaJQPu5RyAs2hRX1VUo9uDgGnoysFrwnf/WFlz6ftT/2QAe0qHwop
oLJ42DmVHSvlEnNzOkSTOh3v7m0ee0UjItFJnGyFbK3aV6L34FtOZvC2PCBkyBDd
Nw5JhmV5tD0N/9GJ3B6sc9vmBMbtjrPtc3Cx++2sCMC4nFcDx1E4wxvURoTV3FPC
vTjJoFLh5163eLiRrmt+3UY4uKneECCXOecwG51IGzQXTx6P8DcwZ5Gp0Zstnnnr
vYD4ymsz/so2Tv68LysAqL9gfYnXYPVW/Ga3/NU++hwQHKgHLYrMbl5iWIpyjsJG
VVm0bBcybbZ64+wnBWoaRpaoo/wqJqp97nF8VsmKBdmTXbdflBTiy3jw4HSUzWXE
xtUIlfSLV5MKAZqssxKpYcWr+Gd1+ohfXttCEUbNvlRsZXxkdpEVRi8YH7Es6om3
ESz2r5oiJpIZG5Y6bAqj32T62nSw8UtRrat2hZEUi6drwTZK6AQB8jj5fB+BdilQ
g877+ZeRldWSwfTLtvYMh6bnyIfI1zDf6zamw/gCxOT8QWc2hhtA/y9n20jz1P9I
38/ieGcfVeaNbipURwjRo86vYvZc2WdCLicpPpTawqWFnNS3NOR7lLIS00Ll/3pH
G2aEdSCUtpUafUtLe/r80xEsAJGiEdKViEI6i9y0ZSiNzlQdB9CWV0Ps4A6s6YUZ
CZEEFwSltyHGmNt72yZCxrgMY3SG9hrLLe/Ho5j5SP8xpSAPImABbHplJP7oZMn4
3N4YeOpC9WO1ycwY6ljA0JS2YggbSWb31MYCOnw1aYZKa9m1I24aGAqq1aWsKGQF
2q9z5TjU4OxgdPfrNlHpKNTO9JhfBJDnPCYjRDiUgB01uQMeoVQqzMyH1+VHIjaI
euAafhixG6mW12cYJpEjdVZ91fhEPzHdeJh2srZ+ucTu4OukFVhRWdS/nnbpklH9
P4q8ZhFij4AqLq46TFCRDVlDsqH/rfhUxu6IDh6fCTfXv/juq6Gyw9y4jlrDi6Ti
si+6Fj2kid0V6EUcxsyNypIrawQs8P6JYqPq/HzfI923natUqQ0KRYodd8CnC4Fj
ybaSKkNKgnc3hiYZb7JijDuCD8Nbg3yCYgd7NER++V3JQbyd4Cheflr6AqOT9lQq
C4mqR9OKf9bPFEQZKoi6MRyjnyhDotkYStBDEA7bAIZ6iDXoFejZarD2q2u07bwT
1UenOibcyKHHfx9cTmay3SMYD/WqHAxM0f5B9s95a6xfEzKDhELuAJZlcXSdof3X
8es/szji01H5RnGwFmnkVpxu5V5P9qDQlKDvOP1H7W79Hl7B7LKjXrj2zdMUaPAW
ZdByIjuIJqO1d98S/+ZZeQTZO7IhVd6H+Id5q8RaxInV7Shj4cKLmhYr0cD51AoT
nbBMtUCQbcBLXha71BJU20azaB/cqRaFK3A/pYgMMGZr4qbbhmDMtQ3IzJy4UILy
oc/dUmDh+MkKdzemeGQsxAdUcIQg+wY9YYFJe56NQ++g+FFNbOXy055VV1Hq0JEY
52pWOFnzFlnpbs7DYj0jqHSjNVgOg4kbdUu+JziEQBKujX95zRJTspPnuT8DyaUu
WirvJSeGnj06SvkD4XBIjXT3cu4cE3PMojDrzmxzTDU2sU9ZCMFOxanDZB9J5Cxs
+KfOzw6+ScH+/oxZ8JUXkY66yLhyW7oATtY1eiV/mr2kcBVozOpMjiTUGqY3SkKE
oQAezIaUa+L/G20k81yD7DI9fhwCnwVWfEbiyrqMGmOLtyGSYum50YKcpVGxqgGC
kPkA3ZN3Nl02CGKUcW0uYu+Fzjp6clj6ZTQOha5VktLHF5J+LIJRN2yIQvr8QiVF
H35z1pnuTqet+U3xcRKbj4Of67ADeXTB3u4xCovnoQ3ehEt/dU9Nsag77/dTuB9x
r8Atc5cB6qtKDFWVEZOy5abhsq66CiV64/eig/EShdgxoRTabsUNYTqtONcpoHGW
D6IruLUpDaTcGXZispOWoCzI3vwierahwBhKIyzIBtnrRDKk5h47+ZsiM9y4QJy5
qzBiDUb90Bn9GHqOzW3pY2jhwm2jDhQWZluaSqxnbhCw9R+4KTMAB1TPyPcruk0r
uDcv6A/MJ1j0dRn4YD9Th3Ib4qqhJnpxTZQyxGttCF+piZEh4ec8lKG00hBuAP9G
ATl/ZUrf2hmC5Qh/fCP2O+oIJaALFroCW3UDcfi95dPd3mN2PiOK1WswntIOalsV
zlbe29bfhx+siBFXsgvbgOv6DdAI9wfHAAu/ZdFMA/gDveb9g0gjKh6PoR0ZzxUg
OyJFN2+tpH3YmUsdTqG3zrsWqJsPGMA54X0NmHnoMiBavgs+7P/kik1m7PaEm3Yh
Er79zIRnqwNKhflUZBuWdkKFFM7L9UGtP3NkEE97cYMKEfNdDiFE/mZu1l5C927E
MPMOLdGoyxDB6t55G5juJQt/RZqd17Krv/s6UbsaUJPMHy9vXHpo/Dl0ldOpqObX
8V6NJX04IpxbtIDxOUIz0hgqm+FB2nZAlWLMy1J0gVWGskIiWHfzJBIka6F4Cw66
8NNJqy9OO9brzYHp4dBRpnW/Y4yklZ9nfpwZ8mzdszCtGAHvUOY8+/HXhHf60j+M
YvRkkOWV5mpeXf7WKg7YaF5tRvyFkAcR6tIiggCYQRzJktPfFO1nKggOg4tau4hZ
t92zPjAJl5rII3atz30LQjENrunzRDbKAF8H6wtRIMgPIN45Ru42zfigQgrwr4ih
Q/CubQ0Qhjns4oT7cuqkhtKMGrwH2V08+z1HSItbcIZBDrhneP9/L4PW6Q5AeGaD
FVvgY4EAp2f0VqgB7yugqtx9LfGx+mZxTXg6XUgPIUqKKvURyFSgAVcHtRI9iX6F
eeC5EtScRtapNgDjVn6kbbDTlOjLUf6FMJ+vp5UGMrpXwMAH/9E/3zZlHJdk1Ijo
Da1r7iNds+HgS7cgatY+FrUgva43MTna+NzO7Gif7EM2AblAyaEiC6q3kUO3ePCt
yGpp5/knszrXtDtVL59YigyPvK8cmrB62JTcsUE34qC8Lltte0HJJ4NhjlCcsUTx
X6gP7sszr+RcovHnT6KIH+hE8QC/ZeECGlqcH8cE2SL0KOWaPGEyewMcdztkbWld
gmUDzGBDFmRX0mMIyEy4MpV4GkzpID8edPVOJBET+wX4C9kT+MvxOGnCLdePCqXA
5nGp0QGJ3hzLBK7CQjJ0Pd22icPtaEZmpXVjCCMlHIIaycUW1QVJwDy7HcJ4S9y9
bQN7adYr9gm3dupSM9Sk0v3JbNaV5rrdTO3VigxpRTXtVdf8eT9x2vgc19gfGMCN
cQicZBUL5sTAuNuUd8dyFPvSwhhSeNj732pNdeFXbQhDG0khunjUgzlYfjenr0jY
XWm5z3RkahzNjkDLoR1q7/CMbIJ39kLnqr+yMwptWg+5TzTlOpnN5HhN3IjYCg2J
+caSHvl/i2AoNmd0BP5uUIk7YiJbczv0JtRVBv1G8dH/Mr60cUGqHuW45bYD2l4c
JVtBStsuUo0hQgoiSBRz/H1NHYxl6beN2Wh//waPLUuOjxTS9TyNgvEB4YRrcL6R
0gbkk7/wfQqWcMGyCy3XLhbJWjchSG+YqPu6G7n3bH1Xry/YGLYQD07Y+d8VxjDb
2pDAWhLv0Yy7jQT2z78jZs8hwL0Fm27Dzud6Hr99rtUBj7+lnSYn/jAW/RkjI+rk
aGJkGmgotbeilYndaEg2aFGUx7NtwIUZlhF17m5TxUL4+1QB1psYwQxQPsySWpjP
2D6/FrQX5FGwEUUE7LpODoeaqAXQ2Guup4O30fAQnndfcpxdNJxL0/8R0hqulgRX
+0FanQlWb7kOYqKgi1/HedjWMP1/qj/TPKQ6aiUpbIGfxx29SZeSlOPr+xQaWEZP
Ijt0O1VEFxbYckYLCQCeKcmZ+qlc6fyKC8TRcN53nzORvE3WamAMdEpTEJN6O85G
9bu7wGWaRxokNslDYdPds/T0enWThoFCVP4AjB77V08Mw/FzbVqEO68dw4D/CHIR
p9eZU3M7iCT8GxRvEUSpHyxAwfCvTWXpgu8/0RVi6HkmuTYTtN+zxz3tc0eX0vMP
I3EeOSQKuhpuymsbgHpVZz73Me3hYJvSPNu5mbuS0/+TiyR2PWYZKdcH34v3H45G
fWsl2to9F5Q/zFU5DnapWB5u/QBpWVlz1mo6TnQai44meSzgc2uAKEFsOTt9cV/O
7mp3xDctLuRYNx0HCS+R+rYACWpS5V/S2OWfncEhJOMD1DctT5lmhQ29jSM9YKAT
3XML8R/4WsqdZJGmTbz4IF4W1ojCZLhMVDou+uaPuZ9QuWmY+/NT61KpnsrJYNsA
8si9vtCB2OFIIUebPnBX/ACrPTeWXrvGTmxanvrnDhBxpd9oCPwRIdRHm6XsVjl7
nYrETVOPc/m4S0iWybyUPQUlrOX1aIoFax/8ZBN1WbWBwSujRHhYSQFbh3lo8ezR
wMLZiEPaRMEl+T7Q1b3XGDz5d3IEr+TdF6Ihp1Z22uJ1e2nYf30q2RwRsTzOTiFe
ajKLdDL6kg34yktMGjjGCMUG4tf+DCsDxFe1O9s60kWGPrGY/QEJpNHB3w3naFJQ
Fbzlq6lD5fPP3cJznRVqCfRX5p+KeHjY4/n2TQxHOLj4d7dUZw2NZ53sWkedw+eh
p4GGPYUEHcUV7g1PRfJefj3RDFiENFrp46wQ/3PIgVbT+tjc3mM+KJowMjf1vX7W
KHmlPmjrpnWzYEAY+HL6IXlGsCRgkDCUoRb/2xv0ZDb4fXBTjIzHrQ7lwVKYTI08
ck//T3FsrlPatRVy3jQ/TZNSEZlPlhtRIyUnv/8fQob5ovO/UzzR44UKaONIULQm
J9cwOibKs6mC1XzexOiyWIdn92Re+85pSY4kFH0PfzasMa3sR6v7eaARXJ6s5aY+
c97d98bw8yjSkJus6XHeVXnSrQV98DdRmSTj7/jHXcJpEOLogHBIaKbLodpIAYeT
C0cCU0gwFuTWCrv0MgWkfQ0k9n6AfU8EUKW6WAVBfFH1vmk6szV6bkhXAYsi9BIz
2utr28RIhXAF4jBdh5Ws5Ub/l/aq34xK/zQw/N8EiNJYoEdz0qfKFfo8BfOXvQBX
Iph08iPkn5PYMTpyKluIqc/oXYOoPez686dYPvooYG61QfUqeOQNKrlgKyISsduR
1rdzw4GwpL3wIwddjC1IwU1i146hlAIJuqeTHfUmkAU/4gJGNDMv1XmMPf285gku
0708pf2moPXbPz1TEb47TJs7jhUG2ihmzlZG7U4SzokzxolfE8BoQ3yvxtTFDLbi
N/JazAFdk1ww7YficbkpWPL7TJSoWKwpYPWFKa9ujVcmtLzU6I6DRg6OY1t/94jV
8RXxLnfcpjmGP86BlzpWA3E+JD+BCOlu5UpM/+6YiJfMhOLxhhdtoY/WLxomFoxE
HLRWkHdw2k0Jt2+wM1Ow+PZ/K4lycj9FXwONh1e7VvPhjk8jvHtfmVuhuReSqtQM
jbwAVlmaP1GbuSBY3yfFSoaIA0i5j+lOpadmycrDnXPFcIBw6ln8bOSPlpPptsud
h7IqpaHFerMfrgD9DIW4/D81OKC0BYh1uoVDdXqTVrjcDB2uHhuiFxk+3ZLCo3Ry
Iz0OBq8AUbcfFQoII1TnnU2rxbgIWoxStIb/H0uLMExsfNHgD9DJeDI5YSM5Uu6O
RpNFbX5OehDYu7Er0YExNTkZpGArNDL29+EnyHFRhFh0v0C0IVtQG/jq+UTaL+K5
OecWPd+U2oC3phDr4YhvXAjK0cigMd/zgCFyADs0mKW5TkSDM97qhrMcudbni7zQ
QZWp/CgMzfXrbWatLi61KavG6A3BtwRg8F2A51hdS/Rbq3D/Zu+ps7eIn+p6r1bs
5kg30e84bP+5dTy7E5NlX4Mcxi5NcAyMEB8AiRa7H6vo1o6HFD3Z2+ec3pbldcMI
MxVanktQQlF4EZU3+9JAgSNNUk0xNzmwcZhYWe0XBOKdPOZTEIwTFcVSTZMQxdrX
dBlLXLoXwXqG9tsyiZfSifjKBG1Mrhqyf2BhxFqZ749m4XbSItU6W+wh0EnjX43j
oDVWxzECViBFAASGH7fkxz6MBN2SHOQxYCUYlYALPabftTYfIxR/jReRAEgc9u0V
SaYyVAz9ftKxEB2NTmHtlagJTsInH7CyWbCkwpm+alChCoNc/WrqTOeHJwc4pmi6
Abhv9XSuE1DttRfN7AiuXuRG7C56M504OOmVzCTIiRwlWJPT97wqQjsk+Ch6LXZA
4C4U/v7bUIAD1zxvPW8hUvnwTu66J8AHfDzSnL8OWwAXbvC1n79DfERz5n5AvlFq
BKLqZpXMYPXV3n+FUIZFM4KVZEdDuKBlbu7sY+aJq/NtMtxPcBwbjs6pww0P7RSl
EUzNo7vKsXWGk4IF8km/C8EEyIw/cV6uJEeX3ub+kEZM/YwLVpmvNniVNxANSAOI
8bEtWNNQz8mYeYLqsZBqUGGEgbP9SYc/W+Qyx6zVkRK6mMrUZwEdyobx9VqZj0Al
WQmRBJWFxHPikkQDVcWwvMrYy6+Mmbb5XTV0lP95/Xh5QN9qfEm2QiluhEF8Usss
EpknT9mk/WQlclNwvtLrTERq7NyD0rj/Xa0Ab74GoiMqLXjKd/MzFEiBZSzG7slM
7ZD5aJ7ATSZ9u4Na4yXMb+HAsfI1GtbAItxM22VURl82qrghzvz6YhyD+regyN+t
IzTXptWFFGs6SWGPUNm9/ZGrrDnr9ihcW9Yb8cqaqzycWlZhubBHyCyOFwGzc7sG
INPf3eYZHBZdpPkR1COAQEh59uxrj1JgTwOputBukSHKJsDzJ6CgB3Hhe+bZPv21
aK2MxpJMw1yVQA9pLxf72/Wz42FvwMZEtC+2+ZobKT+22s4HksIhoVhf2lIARBff
hHz39Pph52nBdPzDB6GgnQSZw5Rt3Z4BUjaA+pzo0BBSag8pyf5c2lRtf7gxbLQl
AkGe+u77P5GbxEMEv2XP3TVdFTpTJe6XobLKG01v0JRLIru1Ui40xLQZ8C8rJSUP
4IalHRyhm/VuxLkRt4z+cjko84XTmC124REFkqpg9w8tZvOdL7Sh5SwEFjgvlkX0
Ui4FFtrMYmG2jDu2qWJx2Qs9F+Ha1vWxUR1f0ss0twQBrcTXonLjlnkRQG2Cz8Uy
U4jzPE1XVGZxhuyve7LWNIEycdVoIZn2wIKRNM87KVIY3eR8xN7f4E30MdaSz4Pd
0aRxVKfhO/GTMl6tL5Wc1ALmpAixQwraN47z8BAEwSX9/H9RH/Ge+C8OL1SVtDDQ
9KRU9Mi1KHGqmhvTiVYJ9MG3CMp3knkL5nDNxQOHucS7KAAekP7iULUlK3yvCqtG
O87lkqANcXbdF4wqGQye5DwnsIZXSlS+va2VwqlorxL8wAMSmsqA1WLIKLfSDzyi
+oQoPGTMErvICumAY+xaVqjpS1nv3pucvEqFa66ER6PMovIEusGls8pr0X8T5hG0
H7Ew0330VUTdkNqN1SHrehoGRPTSBep+mzVColS/F5XyBFZGYTmV6Wt/IQlqUO6D
u7ijfn0Z029nWj6YQuZm/yUA62VzUSXqszwqNHAs7LI5uB5i9qlyv7xlb1QlyAvi
73K+Ro9Q6jB8jNAe253EO55YW1H175z3zqcj9ZozKKcG70bWhlBg/K2Gdrfw9aRE
07TZ0qMAXy0jezP8peFa/Fb4aPpaWtgqtdSHajt5HE1rQSETSCNCDh6jTJ0DGGlN
fBUUG01SK/H/gannpR/+kv6VatWpGLuCrE2R26AM6+YhwR4/2qcDg22AUIIky1vj
YbV5RDZNDJD8jGakvUbJpb3nwvjekcGVrmnHhghDW3L8O9U8rgs/7v45SNwpdJSM
j5S7Qcu/LONk0Syr52z9FaMNOnkRPn82Q0hmFthxsM8rqdORnuH26xeykXjQebv8
0LZ5mZxYOEeYEKF3edLtG6b9SCANh66Cd8U7sA5D2f9NRzN3As7P0kBn6rgt8aYf
3E9tBB8pbSVvflMJ7LwXKpHPXX/zguqDvHmkvRREIYf4hmp/dFsFU0D5o6p487Rb
D3SJPtsE/HiJuW5XSBlDUkdpvHe7zSGzAKnnNINi+yMRnoV3rlw/8iM36dPeaIqK
7MNtGy4wnxx0ifOxV++yXCCmPBtA9OwrP34Xbf4avQ6wsolsI3iwFoc1O2rBBD4E
5hA3WLv+vMhxwppT1gpNBW0fN9XznM/2LHWZThkQSG5A8m2kj3UX6aRnI7WZD2tH
MD7+KCU7ryByPF3xm1odz+cH4YgwuoGyLvV8/ChSdgrh8WZZGyclANYHCXW93jK6
pSz472mG3TNolmyvcckFOhlyb/uFsVIqN98hNaCTixgVVpJw2cTHo3di+Aw3o1ee
L0JJxxchsJZFK77ZjDVidMUWdr/dOJnjnmOtzQK93ZjnUSy8uICjOjP/GCeSPjCp
mLgP7/53NlCgMm7ZcQJ2xOIP/3JELc5k7rss56YRP0nsN2QONvg4QielbQ9dNfvp
9Z4R7A98Chb39Mw3jaPXxipmzDwwKxQFK5XJnpZG6IWcedlRrImZDxyre0LNG/cg
/7jvHLzfE7jehYIrPXr8w3ssJY3a8OygspN7VBzX+FeIYbt9HOLC7eQMNnmbWWGF
mFA4V0Y8OU7etk2wBbPvPshPcqpVTL47hb+o5kEu5BbZgglWbso6vLp6K7Wmz4QK
PO7NjRaTqumJ0VvGvP6Adq/j25cPoNWaxGkHkbypLtwbsD/59wd6eyCwUVXNeEjz
5zWnmcuuoGe1MC9uMltTfkUguP+YSkWs+hPxbqqnGijJav7OduGfP1+ckLzmVBhP
UrdiPRGfyhsDkNZ9LT6C6WBrpC+BeDIp90pBkH3jN0ebZP1dWmFk8YC2BaMUH0E/
ooJNGdQETVwaPFaSgv3KTmbouX8JsIuc7m0uEQ+8GGER6xucHWWavyAE8YA7a9aB
HSCE6s9PjK3dvtTgPKNmmR2VYKTbKbKTHPu27XKlr1Bg5rrxbS0/mE8GwWRQwvTO
0WDS4PSkGXh+YVGpM6GR7Ac44ovaeRNlE6rrk6yFLsrETCr5HW2WSTIg4KZQ9Dr3
BKBkbJEOcbEjRYhtUtCqp7bixQBEkcHwJRVHxfFn0vkv78nEIUTSqHE/es6FIQyo
rXUtn1K5AvKI2X+t/DtdzFlCz75seInQE3u4c5gQd/jDvHbUDVg38apJveG9Rsc5
yZoLlxhGqIbdc3w2rO/5d2EBU0zvpGaT/Wrq39KlwuLEznAjlhQ3EbBBxu4GDPLD
Mpjssvhzt/w2A+55vHvnnZDiSbJ14RgFb057AryJOiG23L7FSlNMJ4YUz208esSb
xiZXvRwkzfnYWdaZ8gFwtOOSf6IIZRh4eibQLIn2pk7rAnFJuyf2fCB3+Sp09G0b
0dtK4mZWrGJZxy2qYT6WDPHX8kx93yd7CeF9TXvtEcKDgIrdE/EGBWEPdW8ryfFt
imHuLGXdRPtpmjzbKYPjxz+Ycyx1dwzjeS6Wl8Bv61qu9rrtzCPB7y71Myj/2V0q
XJIt/deY/F4HerLxfjUVvGHEa97lThN5u1gq6oA1Mz8171YCWIklTtAvJsFHs0CS
cNzFRhrz2yYIEGZY4u8K+F34qHQbcK60OqKSGH76qnE91KSwBH23H6QacOpYLY2T
J42xZA5ol7P7nOJOSa6LXjwUzU+JX9J4Kcj209ViBjrP/oKpWPMIRRbAz+4J7mnv
xQUi2ha9BcQJlSSvozQAF+hAskKXCrIPeSxSd4xxPvwrdiG+b+d1Ma1PCTfN5Io6
WW0yYKuz5jZJ0z4SUsg2uMrZ0qyX7MExre1V8A5edztqkOQOrLs3l67xcTMTjSJL
nutBvy5eeOmL7sHb36Gsg8DUGWf3ijDGW1BQRpxKGXRmZv2NIuYDpcrjPx8nD7nD
Xldlwhw+O8/NIAtJtAHp7FCueyO9LqiWoARCg9Sn1DvufJdHeEfWhz5+aKSAkK+j
8yAuAbraBd0+iIucbnP5qxxpbJ6UPC1eK89mB1MmOczA06RdgipKrxFNT3F66z4W
l3V3i6+sHznwjgpNv1xchmr0zVDP2Vf984TBo/4I7Rjl4tj4N4yoDLgyUZRpUeZv
uD/9cObv5W6I/+1ZdhSPPJCdTm5ajZOxTr/rg2D0umG9GkgijQ+VDCaNgNoeflFw
4/I+SeM4+NdMi3YLSWy1UWk3bN2k4+SaxtMf/PyGV+8Kl2tTkujrvOpnZ5WH19xA
LuMqKsq4t4dVGtLfcqfvhhSNeP8rGdXOxgciJvGu270pi633hM/PpEFXoftHoJwU
E1k89W3v+YgXvetK1l4Y/ZBHzR1nX+L/Ko6BT3qhUovFH8txkAgY31WydINGQOI7
oe+Kn5xF5HulUEuqm4bcFsnfbd/JuAm9TMSvE3rvj34XkZ25V3FYXhA7COm3DWXc
+cni3+3gFuEyfSKLjB7eOyVglOQqPggeEomCbGwxnzeQF3qhp6foondFRXXIsOBs
hRiUon1igDcKUAvKVtfX4CnHdCargNJgPcM7Rm6jGX8Ckn5lmOdZoug4hAqrMsUj
q8Nf2oJt6BiKOX6tQPv3WL5LYwRTJ2+LPGD2sEFo/WtvP5E8HjcmHVqSAYGCkYTi
jHHOAXuuKIf9i6fJ6EpM1CzZgqi3ar7NYqWtojikXYYAHE6Xzo0lihqgrThCBfiJ
7xNDHXnJ0/IXLvHYxF8tkrJyI4OXrLKZIdNE5eU84BQww2cuCbJEV6HTSr/+nWUV
aLeo1JuHJiOn039YkRAB7tj06QLKOujqZsahXsinD4iZmjBYyW+wgTNkM6ST8RNg
OmBV+oJIfvch8d/8+2EYFg+EHiNultM/eRHePAX2IrVngWWeHa+pYsM8G/OKQHqQ
+x/tOoskk+qSN3rRkQ5D+GtlCiO4hafbfoiY+47f65mxgRMquPUrtfgs10b+lIh8
8lRxRPI20Zarcb/dOoz//ZRMKcGUhrEN0sWi2E1r9Tulk8UT6DLe24JdSpopFx2k
dofRDtZGmciCfEtQv8dsGZA0uywklCwj0atz1e9bBwuZfwrS7JWZ6pcUwLLGdBHY
CBceNVpOQwWUEBtPUR7atmtCyxl/6tLXj3rFl+xlWSMNJlEAC9P1CCphnk+7SwAP
Vtx7TQfDt/hkhH7vUget22zYIgsS1bbhectgO9obfUTqB+A4ha+tBE7tkx3LRR+w
SjfXl5w3supULQ5DXAg1nRNgrCTTzU3Jl6cCDQZXTaaCUlZ0hSV7frHTNtIC60yC
AdGjd3VQZSXFfazz30IryxNHVoeWrtPDC1eBSHdPBJ7x7ulasxjgTRzVRqPLEkLt
t7TMHTclszjE0ThdkAGklgYiEe7f0t8TnO6/ik1rhMZlW7Yaaw075m/80QTmG9wU
Iybiox8DLOmeQxcXTURbzlUCsSaKKsKZC84r2ia32ynErGMKmW72szMZNHwhEAIH
xGo4qPBc0ZK6YTEWZuFTRYV0zJ0Sf2+GENMyje4XZZQfDh20W6U03cWBJtNyg/nJ
VMTapbXeYnthot6aB/evSuDz5FzkMrccRHTKNbfyYIvNs1WTbO/YdnS9Ftp93MOx
ULT2vrwFtRyXxxHWGdk3noKmWOQJ5SNetiA8L0spQ1Ar9eM/SeFwpQKbq55uA9Z2
0xcOB7+upQtiyn2ZWLK7NFe/B5yaLuCK8/dw48LxIHdByV/pLI0+XV3zqAQcfAdK
HDp+NhIdq2aDhfegBFwNObad4ywkMZVjc82s9yldoPqJ5RsiAzuqNoT98sT7QSZc
91gXpflBQlQHB0UOCN9vCr6yiv1dPU5u5+Z35vG/sixRXsMZjSVwF+OxCX7YHfA5
cjAIDMPHiE8v9P0BtSHe0yAjKX2w5oBcBUOX92yasflMb9ADgLEgi5N8TFVuuq3C
RSRJd/wv2I+qA3UIP4O4f8x/JgRm+KtiaONFzOktJC9lQLHzkuIJz3SJaqFiErpQ
1/tDZxHE345sNNbfdfn815WSRs/mHu35OaDzSqs6+zWtZ1CZEa0Ax2PBFYiCFUAT
ebXlnkiQtvVxqSKpqvt1Y7hnddn/NoNR7P1lVD4oOHlJ/vsmx/MVNtfADsDxvtTT
deC0RiX7rkngZzd/shm/xRKaf5NU77sMjifDqiR33q2Y6GsLZTdMVigDzhqCD/pY
XZmhEvr3lc9qyKGcQ+ZM6UGOnApdYmBTRBJLHu8Vs/ahwI7fduYX2As70ygBYKTK
eBx9opiUPXXr6CFY5gwK8zluZcbX968BOHOyLeOYeuiGRjpSVoKTSgAo796IzGyD
2TCLy7nF95hFVbXO1q7rYAyvTbyrUIn0Fv6HRTrsSPlwIb4+xiXybJjHgkdAP9rM
+y2E0P9ZF6p5xntmE9/TgpdlzjE9rbTLQwmejyvno/4fgAgXZKH66fpdvv6DWM9b
TDCYI2bj8/vrMzThOEaSTwnTY0UmK/koCX64HWU1iFphrZsISt1mMJaZ/va4Fd+S
0jrgfYsrVVEspDzEiq44QPODP3qkdkA8yn/Uk4KD5Uz913T52pFKVVBxkq2PVSYE
9RuXAEH266rM10PSNRGLyV9PpSr4e20yU0Al+TeS7Q7dxSLyf/nD0kkfmWuO5ycD
W+9piZ75xf8FE2LFzh+10lajdiG2hHpqweLL/2vSZC5883hgLDon1eFQzDT+C6Rr
sKvk6DqlePDS0+SAAHVjIUF+gEql1oLDjKiVk9jk1GN8bTDAQP6ON7mDKSJbvstT
775N3mc5ogVq9Hy9bokNDAchZUoBcrdY6uo1lr78Rq7gpXmFbdeFB4nUvsA8aZE9
dRlusZMwf3FOvvDJp34+WDFv6v/lbNIVscLGNVGU2xfq6l8O/k+5ZbRW1GEZbkPG
f0IihxcHahFtMadmApjlU0vvtstF5YsHw7nQ69IIeYO1i7lc5qBI4s5BxhOe+PUT
zn2sPQFzP78UOld2Iit6+12qVxo4wTWfIsjS44L72WHCzDg4a7sL3qnlkBpmecuj
SaHPf970L2OPXiYkoaqWEHK941wKTH54gQD7vJ4R9FuM5IF/Ktn32jSR2ffOqzH5
lVe4/XyeIddaVWOAxO7vHtSnpowbQNarvNzyixMLJYqW3jsBx3i5v+oKnsZiP+kH
EGFwBQbwquyeSghEhjY0LlKHn+zWTYHobHYaow1B1PvuM3pChN5pBlssxqzLooD2
JUXYeBHtzAO+wWiYICtEg90n3EL788d0Oflt5hUrXQjbPInU96mDuEvNKFSjnI+n
HlyUm4AgitgZQFXOA7ETcTwcUT/N2nblNiqF4ihYKUSHR4BMWAehEu8w1iJDOHKP
406IUrD+58PbkvT9MI6RdpN5+sPSTo3Mkkf78OhgmM9VmxOh64u7ZOQIHOeDeL7F
kORSMyIzdoBHKu2PXKYA7Du1yPL6ft28N1d1R6hW+MOfi7s28Heu5frRSDY8SbOk
ot1j58g7+8dyCaMfABHX8de3aM8zvZ7+Dznz6h/W0slc+Z2TAWAcJX7iUJdTl5Cv
QuXrSWOg6gfd0E5wDpi2jjT0XGq309+LAfEYADgE/V0lrQhjGNMPEj5DeJABLgfM
L8pAvWdRh1tSejhxtyzxlPP+gG81GS9Mi9YuwlCrYuRl3h5ah6CDA4dTxgD8IYT/
EWatbAuGZ7CllM6ZDi+C7RpgwmwW/eZ4z3sMekp987qt8/J+GmvNAKCB2uHZFSI7
Ua7IFnsE1HxSz9pmQBIhwYhY8mu02NBUIgeu119LHbHPc3nChHYgVpedWEQz683R
oTY5XGVocD6nwL27Mo0Yl0QlDfHGcZ4R6zZbRPR5PJZ98105T+4/jbsSInBH6jCy
OLV43pe3uIRtHmbtTU00Jpw1aitbnqD79zbDfE7Ql1o7z+A/Fmi5QPfo7o/eohak
7kwF4kx0pUPcsn/PmoPGv4VWK8oqIhLLBXizIqBpxcrgKcU1x0Gsn2E5iRwOQjJB
j+gFrAeN3CNt1GxeeWDcJprDotnLBgI2macv3Wu9VweekOuHy6gIfApIJ+VuqQNq
S7P7Bjv1PtTtQl1SaRH97tRzfoDGzjEvGBbW3wRUWOH8V4d3ENXTBXRcg9gbZnlu
3V8H1ZraWdXFU9QZggVjh3uJxttNwEpIpaB/Xv63nWz3f/qxR2RHUZ7SuBvW5KsK
HcuSXqcMjVhzM4aVozaC20+3wfa4dR/tOQYR5dGNjUCNWndXW38tLPlQX8r9FUOd
3m1WBs77FG497b3ecvYAcs/K4STDG0bwinm3UlXtr1TVDjT3UyMbFl5hkq4SCnGZ
6m5WMeRp8V8xiMbk08qbvpNpsxBIbnDrQvvqbTOpLoyQALMibdMbDKGGvWSi/tkH
UJFYjR+dpixtMU2mMovazcUS00Jsdkap/rNumEZsYKfDTJLcL5oJd1ObK9oCTiLM
XvcEIe6W8dcgAgaXxkkWxDHBl20pU26okSxwc0aGwzhprRVQAlKGKUz36jz4Tag8
/+9udjlG5xHudhzWBsHWoBeOQsCALGfgxTbXUi4hjuB/QQrrco3bmv/F4NubKKsD
LiPVVrTFkjHs45o4WAGXS55dF4Ra4CDH3FT3Lz4Jj1tLxbHteTfHuqHIFTimlbFo
vhp4ZHXajB/j2Ik3YaUXYATvYc11Bme+psyHBhwq5RQSmV1KfdulYbLr9awiAf2y
X+fYESb2KNKdxZOhgVc2PkwaSVpk4YQntBNec97FJEDtGIgZVpG0m6tjuoyaXJZq
0pON0ZJtUva0clAh6AicZN1YKILMrOsr7A541YzaAajrcg1ymjp8MVtQOabejAKV
18YcrACYAFtUf+9YAMuv8D/JB3yQ0AbwJ0Mr6ZwF2SU6/+zXyH0iLsGyTBge46ux
8S4t9us/WVrmQBZ+XEP0y+c1lXniUxBG/5dxo5R/yqSUWUHlbejByNiz0nGX6on1
zCUIr3aJcaVQgrdpE84XhVYo6JQLdZ4fZY14Zue3DxlPRlO6zaES4Xd89sWPlr+n
tpNJX68MEKe96E/344o5BXRnKtMJ56BfG44/SVSWqdzBszPY9NNEuio/v5FYX5wI
s2BVdyfKdBrA8W3n68k1ySPNLPmdxESa/LtpgLJ/OKa3vsdo7U4aDXalzdDRtc7V
I+ERMEcccQPxy8e1ylARfdKrlAqDFSQl4Ek52NQ8YlKGUGH8PoszYgt3QhwrDfLV
BFQqTjTFWWjHJSZ930VqbAMQVvhQu8kSUhapLQLp1lWwa8oZVbL1k2xA9LGIyXsR
L8E/WD1fKkn8jV7j4HJ8U6VBRw4rGWWOFBuII7ETNDtwVpbiYSIqnEtY0pNm2f61
yLLNT+8ir7LC8e/1Sdhd+X5JvsI2/tBbnrDuVtq5DYKfKii917iCM6d+kG0qTra8
3aLOHeXfSQDDn9z/jiIWEoD5xuHW1vdY8YUfBIDP83l3sJ6aMr1Bugqm0n7SN4vi
BPjqmcMYyjC8ctJJfe1CLnFQODIU15SY2M6XVjNxPe1HDR5b8fsy2CRIvWpg91j/
uKdG2NKRhPnPmes9lkDdcvmX/osW4bIXZFmOAtL0gR2dxNNlUJArxnfPaQypBSGN
ZhOqqEnZVwXV5SMFC7ZgAqXqxaieUqp+DxYFKHo1xF0cQVWK2mvLIqEue8rI7dUN
CyNvbPcavfWXcXEqpNLs4/img8l5f6Bkqa2O/cpsRhvCMKpGGQQl5eL6vC1NEVlF
uLxULoy4ZYQkvZ6MgcZTyqqExIXZUnPqKHSbel/M3KLjSd+ztIVvZYAu1YtU15DF
`protect end_protected