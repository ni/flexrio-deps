`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
hVdJHWSfELCmA4ds+csnOQAALbB3ps7EiTSHEDd//nts1r+JQrRE4d3bDPRJpiX2
Sl8d+xAK9BIi4i+3ruAzYvB6kuD7r+gs02Jsvd/1kn7JYK4xBxCjtdDFjVHOTEl1
sSh1oNiYUwLuwR1yKfP+xBhqxD2Dv6pCKhH1NdGilpJQ6cvivGkSunAu0tzP76T0
4x1pB179E7uIeRplfHWX03KzEBF+eVtfgXVp2W1BGjfAe43y1pCvNYZOh1+TY62g
EgAFgbo7pAujZxZy/YSiZjUr2mGp7o83qMXyusx8+rQ41D3X6rxfuP0RiId2pOpC
6oq5Dfkx04a1dk4s8w8cVg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="Sm9DkM+kBxuxXCFA+l3fFkxuSWV4xqRc4Nn7Ji3ukao="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
m2emGBqRy4AuduN4dffN8194qYvc9UXRqiQc56IrQYMiIVQPyh59I8SYabcDdspI
7AFHnvKD5YaF6tQfxWm+mlcmMEk2Y//aUjxeiGGs+RkKgbHitJF/K7nqg1dmKvDg
a/GaBCq4Bqh0EehlN4ntP5HxM4qcvSfh5m/Coe3drc4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uG91daMWA1mGkhgP3oZKMYye3UAomMWgG80HuuXg2E0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
c9NqBF2D1wSep1rW7utzHsk2j40aow1MnrccxUTvKej2Q1cyeDDbgAml4eTSXI8z
QYgCADtWi7S8BeChdv4B2VxKcS7CMq/DaQrOy1MKTfQzfAlK0iubmlTkljLy0Rwd
cTrJKn61EKbSa1l2NxJKw66NG5i9toezcB4XROs96zT1lupz8XpOQMtG3skiMyGE
dM2X2k2/dOzLIohCH7VOLoWiKFtUs2+IB2lDudOdL6UnzXOGUUJLB1Sap9SMZS8A
LmjNpq83TzkPLr9LSljn17zaWSpGRvYABoCCobDLz+aIUD7qOpU6aO6hLBxQ57Kd
6L7yMlxf2UFsVu+20ilkQW441LbmJg6ePCSQTTFk+PPHJvoUM+vYgTB3YAgfDFC2
aAlTa40eWvjcN4daC4BUSlqMrZzUvWNGyjk37YnXQJrcYPGkkryZkPlQtpfBDySC
Lki1wotb34iiAMsGBNqI+eyG4Wol5H6dN41VQPMriWz4LbKJLLCTON2YQTN76Icc
BbbM4SvmHf0xz97vNkH6Wc9BNG1sfOG2VAHl3HFLBFcXqjgEkW89gYqplp6eublJ
PdUB9T+kd0uwWUDDwZarm7/xBz/xb618iMrC22PJvErXBkw6jKG2MOdFujYmjMc3
pLk46V9kL63ZDEh1P/8GWu2TJq0BVjpyOOrIqwXWkvvT/9lk0K7ftTb4tPqH8NVI
4PzfUu2f00+ujMXbvH0kMX4eN8E5Qpc7h1wZ0AHjFjAiG0LYyL39kTOtU4totp5V
ouCT8/SvUTIqGm+y/maK8rIE8ctxIZrj7Dy2TP6PON2fbLR4D2AGZJj1umO8JcwK
pwJNHOYPR6HT3oULF2GmEXS9rcvUUQMJAYpJFbU1bS9gMBKpxjXZN1SYN46sL2lA
xm1lNV2//v4EJyrmejl3utinsaQuJIwvrGHEyxhi9DeRtxtMkO9MXhvR8+MjJQEy
/aPykguDd+8PJl+1IfG0AUNztVBRfn02LH24i/LlukPibM7NnT/eSZqB6ENm+CUY
w6nV7nHIv6HaBe6k4zily3JskQM9ypyNFlAMTFeqBNTr8YXPlhsEETldpX2uNkcE
THh+UX6yxE7sqkPal+EhYFFelY1XS8UZ6oPV6pXf2a7TX1piNz5iBcD0oAdWRqBJ
qFKYVGONoykRrVhlnpy3Y6dpz+tKGN5BC5FQRDID2OKla0sdw4XC/lSaQwNJz7PM
FnK6CJiiMZdqURsigBANIY69vd5UpnF5AU9pDdqD0FUtlQCgh3jRHcQbmstEF8fc
4aBaXajAmj6pm7D7gxlqidItzJ69OsfnfqfEfCSQ0NzeUwOLl6s574pJX4eXf9Ni
PYztVPwQLUATWo7XngUSTYOFcyd3Sy1U4NshXJBpV/GpQATPTQt38d6JF3K5JWR2
6R4HLPKTa/5LvQCtgYrJlYVL2Wt51woJAmEfTdQcsxoMbbNdaGcIpeiDuq2f5kXL
15PFSnIunGK9SpPmeORX6h/51m7QY9MjHpmniYDnQddIygS+f3H3pANYUOivVVDw
Xs7VWmZUNE/KXk36ltA3sGXLD+8GOzEsl+HB5fKKchisHDOLVRIMsiPPkbXS2vqj
+pfAwxAmMt0/M6pjSTbtLnx98Pp8oo7RhNN/B2gTJm8xgBFNQ38pqwgTHv6jAJb2
DaMO4GY8tLj5GznU1Dn7C5913rDf+0OSP6/l2gampm3fwmz9BwSTpOShYjR5rPIA
CRaoTMS6yyjKxHBxwK7P+fUf/TDKQerox+jwdyNjaNjwrvx58ZAr3HOyzctGyiIb
Xv7zBSI/gyXZVBrA27/Fw8wiyjcf9B7jSUBqU6GjMTJ1BpVhd3Wrt6r1YbUwgos0
GcqHcK/owzCNNHgGe+Aq/0yz6CiGm6dKSACUgYmif12imR4CffodFvxoZo17qlgK
YGyeYxloVmgNybv9evnHRJUIeHFLrCox32sWJQ7dmXYN5nGeOJFXuRvXdP1tL9Hq
RFi/aOv9F8tZ4baiFoT24ZSPeL+IdDr1qYrGNkTZ4p3/0ZDYKVDDji5RCFAxtz/X
KHdEuIOBttz+1rRJxTp7pjIRrHdIFpdJKUoqslCu9FgWNtjiehD3SChegSQJXoo2
7IQmnDz/DvxGm4HSluCYOefFWE1rebXRBT/JeMsoRAOAZjj1TJ99aGdEa96l4o0E
3QfKkbGu849ytyKKR/5UZAhCCzznB6E02mp8C6pUMWT3bceYkPVf39svMPNJ2wp3
3aQaYx+q1DoPHsyq4KKK146r4yTJc20Z20IBkOdlZ7Ys4Jf86hGqLW7p0OJCW9/F
igtWBYMJMAc3F7SX2ubBlh/ABrl1RcSD0dfZDtIDCSQlZK6X3tPKWP7XdU9oR6yD
BTSUQLWE3ffFuVdhtlDgdL1/CoVqPlaHzeK44RsyDrUUxh+N52QV3pyPITiUIs7T
tWvCIpDY1jol5IYfAMmtxwaV4ToN16C0cUX/FtZ6fRwIj3/+14pZjTiSEX0y4EeB
0meabifmtqh3rOvC6VdrsKkCIE6RjjVfrf1WSC1SVMG+M0HeeRih8viTz/8gpNUb
ekZL4IpC05EN/pHs++Rfzal4wO7DxNafpoPpKPT0X+HGiTF+FaXPJXcujt4raMen
2Sb7a0ZPiOWCSFTAslYL3mxX4by7Ov74veIIP2rPPnjhnnYqMLsVfh0HEby5MpOs
`protect end_protected