`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
CZ/1hjxIYH4XUI6J5JyuXbt9t1QeCxbwcXbZd4LgC66lEUdvX231wUQdOLhItmR9
/WGdBhBqs3DYXHSYjPhho3Iad0PJ9lpgfRG9+Trp1xNRv9zEIiRHAelIxOvBvRDb
Fb2Ed8QnQPFjnujps3b6a/eXe7WIfbcUNTAxbN7QEhV/dNjc2neexVke390MQlcl
xHGLKxFs26E1Xr80+zZYqwYuOo61hIP7BPo/DNJnl4nn5nUJ2xcHyFQQ541XaSvK
Kocec9GOiR2+4syotJDl372AKGGiMbeuX5fupm/OdgEL6PmgSclxI1bRZvBIzB2K
aJ4Ht9ppG+VK9PaidcPmQBL3qNXnzeaI2SZL0JxsxHHW36ZKqZZssv5jAXisdxVX
N3Qp9blramGy7/aDDDSt0Dx87VyQKDQxp64EsrPjnVs7iZowFyiNsAJp0hmyGTUS
Qfwv6b/xExXCf+mbk0afowHqOULooZCUo+ieK3YOPUd2RzFjQcWr7NezATxxEF6v
J9o0xYuE65ocmJ3+JX2DcS9tSL9eq91s/P+RUCR+5zbnTSv/sMJYOFalbmFzya/r
KyicEFuI32g8tUyJLan7rSoAqDm/Wlwjvg9fiu1I76KOvnP0NYAHVZ3FjD4WXVHF
gpigTaTPEI5jd3GnjEHRjCmbQ04YrLaJR5aao66wkyr/GQpeE6UuO+4710frRB2M
80uMCx3CpzOj1wFDoucuCqjLLtsptF8Wrg6Vjl1IqUCwIoNQQI+MTw3uoufx87s2
+BMG9/8tWoskJFx3xummXTxixYiAmAkU6RBg0COomyvNw51lW4WErt3mm6+pu9dY
1dl2+ZH12D+9TIz39tQOcTGsSAqjK1u8m3sRu0e8cVhB3uxn0a2w0y2gjtgD4fXA
qff50HkLYeHYDzQgTvbM5HErYFsE9L+LBuaSAEBcT+4G1hw9I5OvekxvjUC+Da1B
qH2VRcsMeqE9pxOAbLiXAffV+bMgHhsmlQgnVu0rQGqJE7AEtCyzHIuwdxw9wodu
li/nwRtESPodLgLC5jpo9lFHraKVE6OHd4pbWWwSbFEz3RYwG7kyTkeJxJDjJ1hL
PcFnSvJZDn9SqKA9M+Yhh4zeJq+lHeF3bPhugYWEyAqlWEw86TFw9sQQKXiQ511J
k7vQ/Kw1kVyhdubG/kX3mUNqe8Fna1hQjUtZa57PkCU0AfX9HJp+kYaPRl9W1SAx
xMRHP5EiIOFsTzINAjX6QDLHgjZVPXYLYmO+owSl24IXYi0lTdPYFlDa2BRkZjDR
4v1p9OcWNe35QtuFGfVqzl7dT4bmrQX8cns+rbqa9DrW0wWgLq3QPgzry+kFv3a2
KeAivluQi2fCGQ9xc8ZC3zQXb0euODVVBS2JEnwQBqnNMNbL6t0eeG20j7vioPei
3r45/+iizjcMrT1/cLNn1E8+kV+fb3ae5HeRdpHQEdvJKresf8NtI6UOkIv0Dp11
GaGiL2+M4CdTK1Hqw6ginMBMeNi8hYISpK2ZbC+2S5W4D2uFaYrLZ+SKFAqR76Ce
aQVibKWX+e3hlr7f9pfko4aWNq0mIo7ak6/G0lhZ8zMGXUxj7AfVRPx3Hcaws4US
20uJhPMW6bgMvHhpKhqWwskW10LIeJ1V9p8CGLEHv9HziRLZ+pLgxHdB6iFN77QF
bXres1t7Ki3V24xgdoxTejlXOI7CqXC3tL0IuoFYwn09TKTU0Gr3xn7tTTn0gqKR
v9HWJzLZYDxNdobotBZjoMpbEZIjf6DxLFTdw6cvAZ5zskrA5lAAvwkj7IK9gdDI
GebNZUCWvEBEfAeIpIeZd7ZnBN7GKfwN73+kpczu/Ez/WVSGWLTiAvg6h9MdlL9j
bUWEdXZQNVF5eO1o7uogEOsbefkaLmxJZegqHj2EvOggfDdbAUAPZtPsTBtbhk8Q
yRq42i60oaskCJ9QJhuH7XDYqxngl7kYHdgmzXAsTsSRkSH+GWo26BvalfQlMKFw
92jDKU3kLKmKPEDOtuyuKmElOTKyVD0pAdyaoTkrSYPVCKtQm5YfqnGEamy2ETpq
tG4XA4gqnDxtlA/hQac+tZU8tbwE1I6VuL5Og9Fhc0wRz+Dkvw7d7VCH6q8amr1i
ddzQY5jE1Ew60uujnpwIc55yqZYpWZNKUdCWzmyZeFvQZbUjzeXUBHmVQVZQOtqy
77qcb1S12IY7F2H9tNsbadAGd+9NY9Y2X8e2wedJmhcj7tWZJp2XFDL4fpb2DAMO
LhGO6XtGssvl76JwSbt5UwVVb3UNt75y7IWSN4T0HPa95MNQfnr9VJat0zSJ+aVx
oo9EeCY4ZRvBHqmeTzMMlU9vx5BEmEjrbiz86A9+kI+bCthOiZ1LqxmwFwWZfSbI
DgyxBG7dNeQCazMwkVfTYdIbExtuHN7Czni+3OcMP3w6ZqWT9/QmJqCvkvGBk93J
ereGqBHZxuctHPisiQPVdIQ23ruPTCOPqaortFZ0woHFkEKImv6pXlGFvNpCzorp
AO+5vOwKHsoa6ubjl+RpdEE44llW1FucdljMESotKg9GCA5FnVUt3Jc/iD0f6hzG
`protect end_protected