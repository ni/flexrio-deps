`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1456 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
dqtlaMM6dsCHKxM+hr1+dpxv+KxyiYWY9CkSbLOtYxXG+xV/t+VmJaCU+Sy3D0Y4
GB4brjWtzPr+nVtRifNpISIElPfhpe+dJxZ2KT0lc9DYxnbKzXObdATh4I4HPXX+
uAzyQNZACkIRzltkIge3QdhkHS2pzJqJsREZH2RsTFSWk2jWdYUpPopzizEARP0m
oJkLT4dsw5/+bapi0No7K29HxV60qz7c8ZqCja+0OSjm4jg2aN+fmQ1FN6J7zsex
EJr5g446Tc2R/DpwNJB/NDXBX8pptRgKbEYpLThpTItkGtNnG1pHh5LrWHfPy20N
ekiJEHedbVv5csOydq5tt85WwXlgBYjflyyiwXYPTweIIlXopGgOQEqRYpC1rFaE
GDTON2cBv51K+4n58hGDwsWMaBy/iOUWC7WX3yUvA0hYRvmIi9SDSpJ+AJ30qaPk
lxALp1aRDo+iufxyydc3lkXCvp0pY1zcEufh2jWwu4CwW7lhz5SAQEIjPUmqFEU1
LmnmSFzo7lX+oS0jx20+iZyXgHTocoEzrrlS67hjTdjRIg6ZVR3XYbhjDMc3p5Rj
Q7MbEzSHeroybe+VYYTlo38f04uffHC0JtZiNnz4o1+w/qhkRl2ourE0CKts+CxQ
QMQkoP4495lvYY5jTmcf0SHYIh/ULx+hhdgTSh37x73EZKVABPXhmQN4EPd9Duxs
wMM3NHvglhaU5T9jOZLSuYLKsK4WS8XmrSQtt1cbgaa2PUlPxOS7s4jmQd4GXBUM
2tentiuedxjJ5DElrEsHCKWdIFN3w42ZRV1flYCS4VQVl2BTCVUzR0Bnk1FccXrH
q9oC2hlwOsjjADgyvOLiV55r0sQq12Ntx5u0XFpidyieV5M9IxiYQm5J65qmu07J
QpuRDkgEYJrUEgHUuLb8kArl9mXd8RLsOyJOlDYPq8VKxC386/plIRoYOTENwS7b
nZimfGbPJLvOROEXh4uXMZ8XaWGgwJwojmIEtBTDESn0ICBWuWpN3Qa0CEyOmg7B
z10FXX6aAX+mnRbtWd8AU/wGoC0WYSOBKh37+pn0KOodS57/BTS/ACma4x6e3q1n
kBWBF+l87VMXvq1n9AlTdIoCR7DfUWfkAVE2upYHKxc+LSYTn+Lq63CbZ5cHg3BD
p+7ZXqD5dS6Veov8Nmn2KAaYyLGNfPp8/Jwp4pCtuxtIGZuiOaKA/CXluZ9T5EPp
TFqZlgTnwDv56bYBNaPHW+6U5I/2Uvhq83/4Ct7NIEEG3zQi7qsU92hPhGiQaLf9
t07ZB/4ipc+ktFrwJ1/4fldpGoz8x+Z4C37URNYRUeD9r6Lt9jFZVp93tDPhQDfy
lKTggUGwedi0jv2Rc9rgY6MpJ+/XypN8zOR9mO6FaFLkSIi/mi0RP8smCJvwmXIN
oR4eruWuShn1e8B+lhaP/OfYUwW/3h4INtMnP5YDe8cD+12aw8k9R56WIjGH/iDx
k2UODvFHIRt13+jQJyDwYYanBqb3fjRBBIKPSB3x91NwqxbdGRkyHri3yE/OcZNZ
+NQxybUQteLLZVAn+6I2E3Qf7hxUQUiZhF62JvTuOYI+HxgfzEspDNol06LMv6Nl
LyP1RZWxyMvlKOYTkSRvCbdApSXqpeeAxLk1J8w9Y7Kpm6xpjO8TSCkuEysd/Lq9
0k6+jYfFF/trT3AHf26CK7Xv+2FjgtWzj7Ft6hRro7uojhzz1BOKWbwlVwyq9uyk
0Ca94Wk3bPz4cfPS3GN6zVLjh/Js79xO25rmtxta0XEQWI95YxjwitPWly77/UWv
3nm5bpJ5p1vWl2VPsfD20A==
`protect end_protected