`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
gMcHP74wBZczB0bB0IzoP2xg5wC5NPjD/GsvSQ6VQgzYAsanETMwwsWi4yhFtJwv
5kY07u0WerSDf8woJ0stqW5xF501W3JLIS8KMiCOd55RHBOnavjYiaaLeu7oUCmB
TtTS1R4sO325rP2zOn9YwRbyyS5Ljn+PzFZZUmkt5xMca3p5NGqKtZW2dV6Babni
5HlLuF20Au601B75m2nv+ZRoGSrpkNElxoTibONmX8gBflpIVE7BehhHwaKSucEF
pp4QQ5zZAZjEC6aplZepouGVggAulz5AahlX5bf4opOVlB1J7IrgyjENtw6ysQ/q
DzybQ+ipztSXBGhmcCVU3A==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="jAI3OJE9Sh00Sic4PtM/KZ4WjwT98XM8AMZrZsQkxWQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hyw9IrFLPQsjvXplweG8O0lkaSLBN9Ijv4B5VdTRt6ipKJT9Kzsb5LxCKvkQyF9n
sGPOd5i74hRHnkHfYISGkfxGJCa55ieOyFShOsqTKRLxclm4oja9vTIey6yFm1BZ
54IDCG9h3PqfDiTD847UCSMRvFssyycwv+BRHQMQlFs=
`protect rights_digest_method = "sha256"
`protect end_toolblock="BnLuc3jxknmZOyxfJK70E5kp9u9O8IQ8cgkXv26kHA8="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
xABArkLxBOK6xG+7CdOOiGu0zbCbHMrEntFfAZEE/xRFxZaAZl1QLkuFI77OC2KL
XxG/mrHJzO3taVHgwRXNLDdc8ePbxbAiQfzV3NJLBO+gsBjmIymaCa480cPNpHLx
EiggSl0xPd/AJHEZui0eXuskMV2OnQSTC1K+4nH3vtca5RPtQDH15Q23FLCH6iJb
FaF/habi4FwxMXTxNv7Yr7pgE7lRLh1D/JudsCi6iz5+ah6bkSIEyjNQybIYbOaF
DZKH+9i4LhU1gVLQO/wW6fICdDZOV01dBs6JOK1QGwQBtdAAaY6uV6SXFCNsHiGH
31Op47akHWJCIf1/8KK5VYflQ1/n3WvfHYmiqfQ5oBGA5kkZTJXoD9L6cMdTRGIj
Arv7uPvFviezQ1E83pHKJ8W0AP3rs6RNFJHjNWY4yFIwLybPVo9vgXWB+EFWAlbS
8Eka243D47SR+BHFm2dimYgfKuBARRqaVtS3QrKcOMxtvTbV6w3jYZ51moWDmqDv
FwfDBD8R5+48MUtO7F2jz5rjI41xR6yrAfEv3hqMacqM0irbCkOYCvdxpoYXqgvp
ivy8NFUyw8Ev4UXMQ3g7nqS+/Giu0U1nrKHOrNuS4YSmzTXc58zmT5/EQMjuCO/0
VMC4afbvwBj6fYmlZQBSIim9iiR+LKqUFzOV0nrjOxXmPHxMwROqISzaa5w60sUj
A2Afo8RNcjnFsKobdAvcusEL9an0m+6ZscaNXEg1mMG3phU0iuoYOqeqyyz38ODu
Y653LAfqSFsA3en9zXFOdMLiBgaM4T9bvpLEr+7S6xTOYDLXV6cDebr+Pp4UuZT1
r1OUAKyTg3XRZ5hEj3tiQsodLpdIWwvEQwW8naYZQLmF7izTToNIX9KiUKt3IIl5
VY0aM5EkoyfB4ESHNuGBubCHXPZ77kGhC6qO4iCnofqqn48N+vyf1k5rubEzfjHT
fUNhz1wK2FTghwg6wrxYMPMVoftx/4BdZ4VyWFRhWNrAYiOrkPj82TdPrn2xeFgw
RUGzW5wF2uJoqvGfoP+BMZyEweqvkOxtoFZAuIgpfPYZh7VM8NfPoOlbQ7tpxk4S
tA16DmAf/+R34ja7S0RvRLIH1cHtObgAquK5PQbyK3q2jEqU6W86lK74fG8iPoRB
Owuq6BhW7ZM2G30FgQC9mrLruMQ38w72Hk/GlO2afYph2vR1doayF/oJ6Y/Q9QlC
jJAc//gu4H1AyGat6prAc6zqmhxhc0++1gMPOLdVtZFXs1PUEvYuZTk4Vnx7G73/
uZseEba76rtQv2EkezoB5u5+GkUyDlcjvuLfsPDYoK69Li5eT/39Okaf8HqydVA2
ybDvzb8WM/npdijES7Xk6m6nYAAO4KH4J8KLbfztPBz5MvMVSfJ0gMZhO/nGd/s2
XQ/FzvV9m+2kw5bsUXkEJ70UAz5rTlv158wRcQ84OvDW/kvqTYYCo4pfFeH/KUqr
Ff1yfiB1RjtWX22UEU6emXVZTRz4Vd9aToMC6rPT3Twlm7rqt/ydDO5NE1iEyWQS
i2kfQWboe+R6r7khgAHkrQE2X3HDjxAomxvb1w0hkw6lirFgUIHRE5Cnoxvvt+Wl
g7qo5hW85he/2u/Vr9q7W1xs6olGYYDQGbd7kd3HMzqqQ1i+jL86UEHsvLM3xB2+
CQiAdjHUr4fXTi033QVXLg8gQZvKNEVSEoTXMxdhVpg3vWM47gIGBlg+eeDnq39/
yqYpwcIRTsvlWXxToAkj6BjnPgtmlHEvDJmKLy8rpqTcMOnwHp1QjIZERDgFTswb
6Sa3qowN2qNX8m+iGtSJ63kkL2usmLd9JeLVZ3I2GJpQ6Kf9wC9ERLNOHforW8cf
GZceHqZ3qxMDnrsB3k1Iqp+kkw1tgDDPpsn92seS0ZXPWAAcAc61IZeC4uGN+oUG
ZsmtgTm4SSaoXiZI1qer37A6JQe/lVGWYZmsRfuEU828lkt+ASiYENGpzcwjzOUx
tXguM8Hsh8LI6uAqeuTC60jadVTue5Ieoil9Ffcd6WFUty9N/mOdktVTHFSISrWG
ksBjTEMFM5OR/oFGOmEFDejjTOmeroCHQI6LTAI0xxFFN0eeJlrzzlvUL/lEjzoo
NA1+lo3bKXoY0/gAE6ie9mjdOeW2jP6DFaLl9pVEpwIGzB4bvd+MCh9PccqG/jW1
WzvEH5sGqT/+nyDQwjk8QmUimL7L1ATDWdkteE49CdAzJHXzG/Q6TBTwxmb7Ydem
3HuMaNYPsfWzDeBKOjtBdgY5xGEZBa4vo7UeKQO2UZ9FR2rwMgBtTy4oLdbcw+Rx
GeQddS2WM+tkRS9tv535eMqZHxLyqsLPHMiap8sYg91pc3vfmZyQHqipnosKjln0
fEITsO8hkQoSVYt8HyB9HJCPXffSGZiC/m1nashiVCUS2F9CjxaCD8JbxDaZgwph
TWFcHo2aKoZJvcfhnhyvqqnAIlHaDLi9/HV8uA6W9UNSGKBbZKv1qMR4dYSkTLzm
PdTZGuuvxTWUtyv6GkWt8O11+ZsD6mWxO/VIqJ9d6pt8zFRw0yLWqEARj2AzkApQ
Sme1JFDxuUjM0/t49vbB5vBq+1WJGeSQd7W6uj17OPBnZ0rR5XGJx4VjW0oiEJwW
6Yx/O0ifWSkV4auWa+UGeuU0Ynj2JVNQ+zo5FzZwfrLpgN+4+VMdAMO7RjGu3xdG
`protect end_protected