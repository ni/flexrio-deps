`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4368 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzsNg3HQFZgJUVV1qQkjuV9ZgJ/4KU3IwJNRjIKpHCYuY
0Sk1H8yBguPIPjSr5+TKXrSh32zfVE2RfFCSYpuVl+pQSmL/i7+Yh34psRSsZOBM
ZDpfQdMUfYHEj1C4M31TLQRvRRfen0Lsh4qh+J0sGN0fkcf2nLbxgGOEy+vD7FU0
Qx9Lj69fns+B7IOHTjb0WcfHB39kFkZSrQpC7mLp0WBDMuRv+nWFRO/XyXhsNkZU
0odPu9qDxLaQXvHElE/mlZeAXn8t96nKzcFt9L0ZAilGqL/WLXqaGYtz+As8xzEe
FbC5uuJ897OOPqE4KA+8v+TolIiNZ2rITUGRh5cWENwTGs9XmgQuSef3vJ7VtsKC
1UTHnCUkO/db1O3VxUryWXuATulaY4DtIKRxIo5F19kqd3nrJs3hJVFvXKyLu01c
6ZmpE2n4bHFmYdA/HVmd4FOMyjoShT2m2aSP/l5YL8HZzZCyOIPSGwqcUE4tBzYd
KTmvCy8pAsAZPcKSDV/0SgN027rUiLy+5ABc4zx//QWIGod3eRvml5fOkhYlbSck
G/OjHt9DBHQYU76QnkdztVtjWejdVWZ2Wrxj22gXQIsfGsgsv6bf7Z9PumFL/QmD
F8CoILkeAU5dIJqjkErNO0bsbDxdlDVKWeEZO3kiZNL8t/Oufkxrykrt9CwM85Ao
7Nu1LJLV+T7xzmlQSsg5UPuunbHp9E6i+Lxv7AERwc8TSNLe49iS4Nb+vI1DEX+X
AsNJvrI/IPAqXed6vfpV88n39k8Tjrm7oFHky8DdgJZy67lCgDYqfUbWbB8yFSMG
1OK+ZNaGNC8cr45NXNgRQ5tJ9BU3G4KapoyNGycmDrwHWkGkgdPDRztCXdXQRjKh
xPx7Q7EL37oQXVTS2rvsqV3c8sftUFsH4AWty3qhXxGm3fY7rfydUBm20AcyZdFy
ym8yrZ9cQH7nMdSMq4vDQ4BfubLuYclRLiqS7t6iXLB0WsMBL5sxb7fmGILIC/Tk
igeg260NvkQVxOq3Iu5FLFRd/9Uuf41KGnBXPFues1AvTUkxqvovRheShA0zoywj
mBYBjY6LPbO561hECz8XFATbG8KjdcgXQnuTajtheh3T61Ou0ZRmfQeBJmyiHq1g
sn7sCzIK1aCXWiKe47nsxUvBeTdpxo/cEbbEH9o/yDkAT5VbbfMnon2p8mQ1AL3m
sk+4OGE3P2J8GMN/0rGoSTm4KFZRRtz7mil2IsY0ZUUnGQ1Wlzh1aq1/NRj4Fiwt
oYed4RGlglDuWDfqlMukEjpsoT8AtCz5WHpw7kp4oa2LmRcmt0bGu7p9Ix7NxHJI
xcPKRAF6Iu/GpLf7R5+xgGINIvdVhxYd74j9/wGs4afIx/CDAcQ0yJS6W1PC/C9D
n00/XwRWeTrEaOp/N4AYlCB6zKmRuVxkSni38iLXkGSJpeFNximur7+qS0zgbiTL
d5pL6vLDmBj37pUkFIoXORsHOBjxKpxClf0+G2mknpWkXozD+25JJbNGXMoTsfqk
mcgpEi63yoG1RazwhZ2KCEhLVwgmKL+QvDgZoRZ/J5QmHdX4f8DIblIcVkduLHRp
1NYWK8qPhvP7xJT+Hb6+XkBOBGaaff5JU61UczGot+wO/rcGoDNIdsSkolaKMldV
IPgLebq7o+4YlfXoNufJrOHxvow1x9AulqVg2X4cB1QwCJwoTdtaHqbeeng4eaYI
AEdfKyi91ZXSCCRNe9B48XzJxFL1I1szzqs3Qn8CzkoFEHFEf4lvJTizfJgM9AsU
n9FFhg55huOJGLCqO1yuACLUl334pipjwoidNI5/EbnsBdIyzvqIdPQkqq9L/G4r
FfpuMaoHMtjZ2jqHNo0pK4TvfTNIRBAgB3rwV8qnh7+UIbnE+x+c8US6HpOa89QX
nz4KTHk7UqiV3AnI3/vpx645VN1CuqAt+jhpWLVMa8hrvzCAtr5N4soQfz3Xpo0r
atk4G7SuHPJVbH2IfijJmEVR1vqlSzYAHLaYpdl6mkYnIsfkdNY+rffNW3Byev6j
82lmweFIK2Wil0oXQz9Pw3XvEU9O6bT/pBfgt2qQW0q7u9bhRdNh0+t+3OMYwqRs
j5Een8asvFyaREVV3/WI24ThlwPJXHaWH5jTtGOmqiuE1uZ47vrVklHLv7Lcz5x2
QqnGYJWb4UQreqhMRCz1VYDXWgsS8yEjs6yntEuelNk1aHMV1ZGYX5hUoTmcHTUT
ndKEhD1hPD+kilKPzdQTzApEzDYyABq6MCgg1K6awZT4+3w5SWt4ajv844kQqC5W
1UmsxPRPRjBeEcP53KewASRaCsfxE1tAdAxGqlCl09dJtNFdnj3cVDsAIDKtraWp
MX0kgqlOpeEAg8HWFV+8bfjAD1eENzg9ejfR4ENDhQ4MxaWOcyNS3Kz5Ie+MRjox
3wuzP2Gxr51XB9c3zxLIJ9mYH9FSeYOhYoPpdlfiK0SYeCXx2Spej0VD13E+umri
wVMuVylBiQfEA+tuZ7KyONs0o5dx6WiNJXo7RdGmyo3Hwgda6jUXFLczXQvjen3y
PB5OuAwfES1aQMl5Z5oggsnUJWU4a45vWgp0Xfty6pL/EuHUAbDKrHQTV2ZguuzH
tXhQ6OI9VvMoTBSR7R7N1x2WyDRPtevy/tHxmExDXIxyJ/LiHL1doWj/Pc/PRVPH
DSsr2l47XG28tl5KRnW6G5/EhNa0Qei8Ebu2j5qv+ohwfb5hH7xbprFGOQb/tLy0
fz7VJY6O/wsFZe6iF59Lj5taeynzsB6mbMedgbffkLDP4S+ZZ6lakAa97ckc5EhS
muzrrzyQKPi6Xn7UO9U6zJKGCsqBhRSVcPwFuyVjiFrb+rA441ZXCsmuRkkdT5fb
3I7lTTrfEjT/HQvsfrhviWtztEHXQtj8gK6PvxAw6BFaAd+JiDTkq/75Yzd4sRpA
742uLUypHUX7NVz30DTY8Jo7rRVUQEjeE5CNVgF1mbQeHaunZnoJgH9KNHlPnPaO
BGWnMRhJOidEdDpoHmunrG5HyjaKlGA1zRix9lszQTre6EZSvPMvbrNyvrWW8JGC
rR7TeZ5RngCq7CWB3GWkWkD6/NuzRnVLuTmFCyC77Kqk2KVMtcx02BqHyaLZHLNy
IEqKfZNBJenxYoBwh4AuAP8Zf1EicV47+e6B+ePjNpcv9EI3PFmlxnL7+x9pHOG2
frPky9IRoS6A3IYfK73sHEpyjic1lKpdHPR667h5pVHcR9G+NH/XxE05sFPC341e
1sPmDJdwMWqNBD17iZGeZfL2cfu1qu4ceAYWQBnaDsSj89QR0jwip+wo8f6/IFQi
XqQWGYRE/M+tTXSbR2M/dBv6rbkH9f9FeDb+DPv02TjC2FRS7sNeSXX6wTadPp3w
WhdEwzJKRyO8DS5nZ4fZtjSLlv1TQXqIZNhGuO2YYbs4WnSzTkKylg9AXNjVhR3O
66E/nOV3rWx1271XeJv+c4obQd+tztVsEV89plDKEz/bPusnnfUkJOFPBLlhkrVG
6SDkubJMwmYfqzQCBQALRwUeLwfXbZID3h5N/hPOLSd9dpTr/ejrTTAk0R90D98V
v+YtRSQicZTZ4sYWbtE9iL4HXYrSf0EkYEjvZeDVIlE0x0gkorvxnVFWvW7Hz2kL
jwmqsThcPVdZMUAImlzAZRnEj8NeQokLCG72gJBLn4ieeuJNHuJkem7/FLa1K32h
p0SnivUEKLP1tAY2YE1AU0Kd31ILd6QWFZe5f7pSP1HdL+U6kH7fiXojgyOm25HO
RC21fsD1YIN6fvNcNVYsLJoLTD045dpPMC4P+xz+roIkamNCIbHeH0EqsBALwfIf
Genl6gMZqEH5ylPLh7EEev+FvWz7ZAKS8W5eIwduwR+m1ReHVCNLlHtl6Y5EeoXY
oj903BS6UtqqHwpqPjSf/nzDvNUKGH6Kcv/QxJ0mteLDEZZhwmcuZpvALQx2pILS
wqDxDwYA65lS92JB8tUrFJbqzIYCRVMPik4PL14WhYmEYBNKkaC7NYDcuDUp2wCO
ud7mi/PsEq1DcThfGQH1VFrf3EFqsyNGeL6qlvWvKUpkFUojWLOsVdgxnXMGqCzR
VEIfUNHvMhROpsB3yimoNJAlazXPZ8y5d1f1QLrfqNraCyE0djTNOV0tmZQgF9VN
EVkpBQRKvFgCsnqXVwKPmRLe+5+gGawhQzQ5tGYp202mc50+pporA3Ozsv4U7nJA
2+O9MrrBpsYL+kNZkI9flqbGZ2wqltIbtvCjcIKzIv2hGLTv/HD0bq1J+Il+CgsS
HO3KC89MaNGypkYSorj9+FcpInqT5HsNUWXrzmVF8fX/3esdfw0SHUQys9IY4f7q
Sss8dZgMuBGOxstv1OO7LJi4AdWX6vB8zgU6YRaEXux+suc2Q7T1eqyqWKUOLKQY
pONPhl498r6yPMazsD0wfDK2ggMDMswMsVd2GCK+PDB/07pSoNAH/aSv+rPJf5tS
Cy92YhaaYXDXbTTD+EdeoBKambE07HuxvXC+8339NBPRgJ5Xo+GXUBnRYGqryZ0D
O7IsKj4O7JSUQbZTJSdBTgWqtPZB9UqFbADPHC8W602Kz7meN8AoNehfrefguGBf
6EzOw8Gw4hxHLgV7NLZOIv+6GWp3D0jaSz8SsELnpU1fFUvbhdzhUmTwroDTTpG5
380tETNMxX0ZeYza9wjN9lmcmhiimBbueQlr6im/NbdzNhecP1Wyh7gZrZMDg9Qz
zYmx4+6Qm8J1HHJwuzSojVNrgM5wXtdskM1K6QNGT+XA7Tfdfa641cMB/O6CmwrT
oasvZpCcPn3PdB2IdHUH+5FUG9fnFz7e6vkWQecfkpRc2cDzH7YkCknOnJ6TIzr0
+xUyavq+zW2jDkRipeQmcJnjbLxxEPHsqHJzpQ2kaMtV4JtkIafjerwpSgWQWNik
wP8GoQF2EpdHkMRwqg+YUPZGIH1jcJHlGjBO4zVB7qxuvnNT3fUxt+97tfsSUC+c
lsqngnRj7tls+kEYxwpDEhrnD3NwBGDfxfjmQRt9iFw2n+qs9if+MvRsGR20H9r4
n5kEDjpordHU3RvKkx8kJQycZyfm/f99oNLFqCoa16Cf54PlOkxfeJWfmiNfy5we
QQfhW8ElZp6aaxGmQH066qA78+2U9rMSXDqMGpg2fs3gGy+POQfvmGj1KafYLoYC
UFQEitmUKM+w8TJKxBjXy64LYpnslzjBXqSOPuPD97nM18PaRZK8Oq8SKVX1svhJ
kPeE9+DU0ho2buV++9706EKTEMg7GO2ldXwlPy425daAU5rBLYvJpcM6Of0cVfTT
AVCUDmoD+H+zV1Q3Zmimbjl0xj3l8cmPZpjhDfOR5dWuo0ezCt2qVu16VZkK0M6K
5ctIUhKpJCOFiVz2ALrJ5mMeKfoWhbOq20kfpPXeunPQBgwBv6KKbKr5jWsWExK0
8a0efkIu8Px2u0AoZ9Cx2xrgliJDL5gcaW2qoNA+Mma6MKYLXKJ0J5t1tX1tDIF2
z2rLu5iFYMsXjx3Bh5nkveTf8FeBAC5bkeBXkrpAerhMqrY03imhGDmffxUPu19W
a37ZmcJlBefESXoDVIc+cXFhZ7FRZ03+hx7UE+2WuD6rksQTwFzWv4vepYmKbigc
MMbgWgiAZpXpjUb70NLmqRiaMqv+QOz+wOfPOB+d2ld6Bm1kzf8IJYkExJoMqSp2
`protect end_protected