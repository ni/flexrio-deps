`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6272 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhEl66vkmqNIpUVBO9a3D9et2jagLaXHgpCw8XU+WudeV
UMm2lBGTBxc515BEC0lQCVpnkonfNFmyiTO6WTIU+l3CRuYQYiWu5eHFc9yOAEyf
oAZVUToxuPleCTG0sdCo8c8WANyNS7rwlG6cRVexcxCw2li3yEXFnm6XM2DwLWig
CIvGKsHo5JA8vsWXJN80KaLs6JbddY0a4StevHHuP8m9dxSwPDrA95FAlAkrJ2nR
AWnoIDI+/jcLz1oJRFMFSoAZLEb5lpPC9zLBLZwP3xH/c18Zf2QzskhFm9dFEoSt
v7gKtKXaAKkp+N2qmviKo6Wuc7ezZjXCCS8hLzyP+rug3toLlh3naM3awLENhBf+
JwifmceHM4p4CMj8tPEB+/CXmFsKXfTsr0nQt4MsNcNQU3+1y9k7XlO8072z7qcA
xwgifmuscMhWg5XCJKQy2H64b+4Pbjbi9GzSCLCNtIYAZ43ikqmb0jC/bU6XpaYg
W/TyYQaNs1aPWI2uz8juuAZglUyyy+/A+o+zboLxnXcYdGdJeTUmSIbuwQq5AxSK
7Ww7DivAdHe7Q/bS5Rwe8NhMMw4/uHWEuJr6gx55fxEtXmduPkDoTLEry3RV3Qn4
E4OnJsb9TmYlbD1DPmv2AWOlReKKEWGvZYUNn6l4WK3ipTndLI/sWdoE+iAyuZbl
6lI61QW3glsOMyoYXfRvJ+n/nS/N4NblmmUHY3GmEoMK8pcUtIA8IDrUHVzzoNjB
7B2TSm1csG6qyv+rdth+qgV2QMbzWtL5dWfkdxPOmOrzFgLuAcWSYAQKmjUbL6dt
fq1gouR6QhUb9jm9NCyofJvLoW4/3Bo2T0GMmMRs5f0AAWmub8GBEtwWv5wYPjn3
/VkUEQ0UkoV2IzdGsZEYFOiHkHys2lFtRFGSZtC41j+JW6IlkfRXM5lh067opuqF
HUloeGYD9NdWNgXAfa3f8H1JU+KRZQoz9GSgmV9VWL7g1Kv4dBgDIq8PzdLeXkPi
OMF9ttiE0onWYhDQP9UQx4S2VcFmjB3Z0lbQ5dALQ2XRx/nQ+Jv1aFIwqhLEsunL
ZPcxO0/2xtqm0k6rs6VhgzFnmSHIPGZVANuNsgULN6AQLtB9Gwz3TiXgLc/GGtGf
GXb+FL4vjLB4ASWT8PxwF0u2p7ldSYDy5b2bUtDb/XDMsd2xfJV7yvKSkePeYu8D
y+CGBlcENmpIOxz3Whoy62Sm/D8j2FMd9PNyET/MsvKeceO8vXsTaSGPw5M5IvlB
gFSzS5yq45GLff2gljFGdm1XNIjk4xaKAdeClHsq7EJ42+rHK/qgAGqMCmbaP7MH
rWZf3Eq8i4kG5wGvr3m+XfEiX8MuQ+WNh0LnxzWBLo/Xg0HE6EJp1+vPGXLdrZ30
427UhirT7hfYnsKMBG3FTkQ9G1rzxxXSSWy3NHL/cqySiURxnPk6qKudjY8OYKie
NN9CApuOTxndYNHe8uDvoEGHo41t8VMmGLBYn8Hs2aAuxPWrBW6+K9gVwaoLF5kb
clUKBdvrN9ejkjdI1fLnOg8KYjNEAMPkUCiXSR9qCzmRRbvRVP5l1XZWhsjOcb6b
UQHQldA4r/HVEQf1gZfTlb4YytAyO4LBh7djVnpwTYy8hgwBYDiHkeOlWd2n7lhE
DIjM7s/5g2n9kyBejYuEMPi9uncm6vespej8sk55aPgcdsxS9ooej0/dPzymc+J7
IV/LO4vTXisCM4PsVrbWCyXgfyH0GbSNcWJNGwjUM8iGo2vS6aagqSApWruqAZna
FxEky9uZhLH05ToLQVqOl3GVkF+9/nD0vKMh2itVmVvUJBGp4mrfSbSh+xatKxgm
JPpE1Qek06+mNnHgAECoqfxdQbMVCXGGOEhpSo5hs5BfW2CvBEZQZHj/mjXhO1UU
CEj4wNNMtDC2dAj+GS6p+4QWa8o9lyN654DcSMlqCDkuDK8M5lcZbCKxjqnsyFdh
O/Gvj2XJrZIWU4stHPLXasgC8C4pHkeuPA4AnP9PpmXPBgsMPpIF8kGH4AA2ybyg
eNS+LHMTfr5ddZSWlkiFcpNoynDUFdw4tWMZflNLSgXouB3sf74aZQXDnrpjD8Yr
bpPDcYY9NS404rCPhBnpgWNvp8aObKVJ700GWkXfMaTdMybzIdNqeI5eALhe/+sE
7lP+Welfxw4tomwU4ymcPc6UKiq1jPBsh8/bePBfhoIZzunKGBoAOJf5ZmMXCi21
2SJQYNEag9o06LQhfKC8B/LfAYr5pY4g5u9KEJoR9jqRkQmPp8KeBi+uQjp6QxKy
3Iwhd7LcS3RLsH5xX+KsPpKLcgC6O9JWx4a1PP9oIe6yi5C5vYkgRnmDB0BZdlxn
BgWjRA76umhfeN6Gj0GGOfqH1LPHCdQ4oPOvmgku7A41IEmADezoGbPr2v+Bz93z
aPCX2xQZ/jrohccR9qkz006Ffl0XPv7BOv00MmqUC7NfOpR+5s7CoQM8w3bNKekt
qQ172ksfb+GcEpjW16wdRIpvsQ1DHbMCGNLIYwakwL97mceYoXNPTxODn93VBC+w
+UbNmi5+LX05q5HdUARRBWin+zc9HTUkCU/G+QaqO6hUQXm+9Yhh1LoPGez7RgHt
Z5VdG1nljT9+dbLiYy2UcixkkHBxQyHSySbDU78c85Nb+dDa4s1z4IthLKZLfEnz
qd4hZs3p/zKT0rL6BQpqOL4NCHUbQ+MZLabIghpU2gtLz6KOxqR1/4XhRtezBwL+
Cdldu2Ld8TxZX3JpW+Xu4v+nhyn6v8t1aoW3LET15XhrCJ0imRIiJFCcpOuw2RUG
IWybsK0umW9NgYScIS9RJeHlGxe9xcoJUsikmESz4gJIMW6Uca05wQS16IBEmGpH
benVAh6zALIXh2M9BtjYohdGipv76bdvFRKFS9LvoKjMCnURpK+cBzovRM+vNQWf
RGcLjj/yEUqQSZz1tbE8B0WXtxmM0XBcNWSGFtjszBVCstpRw5qTzBIsX25j6mqK
h+8ZavEyKfBupPImQgIPs1bp1n0UCkZk4nkDxkzEI+RHH5aLxmT3JJdS2vw14/CO
b8th11lzKhpRZ4h925CW06kgTtxsJ30hfXZPGgmlG3g7balWyJp++Ht98XBMpAdg
xcthrbkEnqZfXGGUHbkTsVUMVKy+v9qXtPTdfd9ow4HXsi14D5jNi3+2XgYIR4FH
znBQxpRC6bD5c/9q4UAmB+Bjcm/u43/djDK9S85yqfWIRKogwCJk25lhHSe0ra3l
MJwTl8L+WUfu1OnvXSX+qPtg1hYKoeWCaueAMWxNRo1s9Ny9jKxCQH0o06Ft9x7l
dJWV/U69pfKBAPGD80sIELzmcaEPQMn2KFq6SjUT3s/DvPp/0a8TAX6gLwMuaefn
f8lmT4aKIYGRSOIcoscqtgrV8vQyPPF3a+slIJXzaeUb4teQ+XevF8ZfvFptiloU
5F9YgIy1+Xg0fzQ3jFekgIv+FrLfwP8IAvrELMxTBaRt5XlJGiZpjiQR7CEcMkdR
MGd6HUGwPvturkrjGANXOUsbJ1e0x0jyAxfhN3i/NkjUIvSrBQnIcxbF7qd1j28G
RJ8xsbZpVVeBmFKv5TI5QwY706HhK+41suv7gIdIkCfedECuq0xMu+U440NEGX57
dXAbmslv2EBUpbV37WWq61S83JPp6wJPvcbXTKCaOAcyyZ9TFc3KqLGqyT9NueK2
OFdtJb9Uw48lreFP7J21XhR24vT7Rva9zXItDxr2sHKXUtpqOQtGTxNC6y8VaPUx
m8qQ/uFgGKZ2bZOH9BQEasIzG7HLpjh/MNUcug722QkjAKQL5EbRUi1z4JAJPHok
xFgG5bNyl1uiSEa1Up3xGOe9yG6Zg8ZymyfFYK6CcvB2wtUDhyf/0JcGZ8pamXxK
5ZqbcRVoKCnctCRyXCe3AY4rnZSs2SRPDSk0jnMU5ldt4DV05P3aUWAWvG2RWUAT
RwpAKqA6NLe4ATlaRDA3NO4bIhW/VIbe6EGURdL1mpaHn78FiUSy2bgLzj3qMil6
AhP1y8K9PU61vWqwRgpILto1rAUqMVFw7gDBY+TiS2u7WFBAVoBDP7ursdiSFyen
53YJQQjP/bSzihO7FVXcSAY1Tyu+s2q7yBhySsbQRVY/Su4ovf0Eod4Y7Cn5yynT
ARVFY3B6DViZ0TSHJ0i3kunycHpM9tt7uT7ButvZsP6HhtgNvGiAG7U5gO843rry
SJBaNx2wCBRugaI/DgAa5E0HtfKNDR3jLEehH1E4/3T7wKi2E7gTByH/wR2QbiwZ
RKOvmF/a09ezT0HOM7ia0UWLfv47OSN6EG/lQHl4Y+0y0VrH4CrPvBdAlHN8wuhC
P5TlqtMQe4wYy4a4hoECSjgpOSQaIP/vBCOCA0WLU2Jkh4M+UVcSqbqI5LuxTeCW
G5zhh9OoZa04SuhgF0RBPQQ10XdU5lk9QhuQHEpxkfi2pxYy7pcPR60nkZegfEZc
El+GQfkF6rq1AdTe882xfx0KFeszYoWIrJVCgc/hWz1IdoN2sFz4QS+TssffcLzE
OYzQv7DC3vxE5FWMK6qUjbvi17oM7KclG8aPd4gYbAAy5d1GuPYHgz6qEKnia7k+
I2UjOjZBPB68CstStAGDWX/uwbLUuXmhPMC9CuQfnm3ejW3NJ6omIVyTO8Hhl7IL
lFoKt0ja7HlwxeOC2RyAMatuu1hdl5xwNYoiX5unvW9ae8SlSpGstLShrOLz60jV
EEPu+nwB7JTaxaHIusYhDLl94tn3B1W4aNhCUf9LHb1HIPldlnGgXAtwJLHIxVIJ
4mV/AcYWkUY41jOjdBKfmXXcbPHNV43I/krkhiAkHkbwqAg257u/0B92QTO/qtZ/
Y4FD2fez6U7TdwPC5ThupywhLvnTSLZ5X0YnVdu/9akXepuNObAL31oyucFj3SlK
P20MfyP/GiMJdhZzpotG22D9Imsd5qzUNxnnX1jUIwHiIVWBRzomU1E69irJlWNM
rZyrRXzvGYQoc89hztdk45Sob4XezDkADoE1IKX30l0F3PiI06YDr1OpltenAdIH
JEaJVxidGdyyfKfujhH6zD7jS8jlr92mIDRLYhWRUApKW/OEpygsUalEQe2H3mEV
GCISZ8upsVhnuVO1oe/hKCS7ESPEwvK5Wo/jML1I5Yt8b/cvvrnAvz0cRY17tttG
Zm+sk7wlnkTViiRsA267OrW1oGHbXKnl4rFFxqqIK5450kOGP1jenHZLpQV+bwms
k4xjBfuovcIOrC9v+/1bnDEBKgz9HbbTmHKqZtOG/vr10q3tedmuPH7OqlOTgjKT
n1kzy6xJwtCU/0IuAZhg6FF5CS53t0J5cjxNGf/EULk6DqVCAhKNcbCFLPOUNVnE
d8SqZ4BFZsLHQYYmtgxqpZqYc/WlGPRtsljwEZmal0dvH/Mdbw0WEtnWIuKdbjmJ
9Wes9rGFh1A/hWGJxe1YUiZI+Vi9IUFqW7qRWcV6L6BjkGJaNWchmRtk7tOIJCei
O+SM3tNYH9MxGVYe07LRka5Fs2QBMC9jTmwuJ2NQdsI/hu8w4WF/1qQmeFhmlWtb
W/0CyDGSVPSbB2a5j57lV5eQ3OabO33Bhxu7++yBqqRgUeV9Lq7qO+NTCpaqJUQq
K55Pze4l9l6bELmBc3KFf4TMjUo0zY2bTDfAAHiO/6qFhkOCARP9Q4cmclVUR26f
FbG0WkBHx38yJP2bJ2TsG2NT52y9OWEwhJ8qufn3gFNr7mrdr165tRMgZdliQbT7
PRs6LLGRJxeveHqHIq8cimYWEMaDIrMCEvLaQwpLsUDOtmRWwfz4QCeANo7r0f3S
+522aPEWqDwPbGjAFBBS/kppjqBZ6uI89EcueLPF/VBJ5ttR+yCcj05cc1p/NBfS
B4P3z4GYsHQi0xKGmZ02Fzrp1g/VBArhKsc5Ax/WOWaBAG7h79hvuvddQxcGO24e
AeGShO4PbwvvQ2v1LCtkilYx7YgGhw9+f4jlEfaj7trHBM6hC8ZYGtTJw6k8OQWF
CjfAQyMldzEXutHDUPFpw9cVa9GgvZVXI2sR/ovoTcTVeJgozRXe7qWm+xizzrVO
LVk1nU9ysPjM85wWya2WnbUqf4AxSUF8myIFX1qZw+Df2XHr1ge9zL00UbA9SKkB
xsTz6rRSvN+fuVvcFjpTDfIJS06rc9H16bsfkRsdUfTryUyF7vcmn5IYJOoIVuCm
Fq67s+LKs0QO0L4BJiY8WbKa1QgeAzvyr4NWskufS+h33dt/23uGYjxA1mL6/Ze+
JsRYGtLLASMVJjXaaNqDLmML6+pwja/dxVKsS9/MiZ+l0Ja+y785i/9iD+ZqTYAm
y/bCPady7+Ysfp7tWgAzE3t5YfKMXR+91g8J4vPMdCMYKRUNItIHKpj+MeqSoiPG
yimG42nea9Uge7eyS8pyOM5QIfSdohwTwmjjIanwHQ4Up5TlYj3Ktcg7c6uMPeSe
xSpadcstCDAZQq08jWQJ1mjTIspLQ7ilZJWIijmkfLEex49OLmszUHtdnWcQSXxe
sS+j7bsuzrk6JI3KuvdkWcGJb2hcIOmV8+O1x35hM188tRIo63Pn5SFf4fG/rRq4
0+nEPvxt4W4CcvSMdC1SxF6XH+n6lZRL4AKOfgZgQwxMVWrInZ5W0yCJZXUgA3zR
vhS2nhWYmBzAZBiUIQmS+5aPinrwi9uyiOgWoQxIbuLYLxCSV7hvJYHMNHitkKe3
QFZ+EMTTBCkFfLuHRHfrMP/RloTaSBVLBmG1AirD10oZFANlVdvisgliCozLqp25
yRwqK7LvR/etX89nLxFxsdnpdnRBEP9ZG9dqSgvJr6gC/+lwnxJOLWqmZ4XngfUY
uqpbQ8etZP1LcncZFkwpPPQ7a3W/wbEGsPr+cVJ0jfxi8IWwQ1PXwRYMy3pUJshe
L7IoKJDSTdRYbJg4aqJ0/4vPULPFVV1ReJwncs15j1h5bKXNVg/XkCwzO8CyQCs4
/tqI2HbTnM5TUM3UgI6w93c848h9WdqPBZkZpLo9Csp4O/pHobGk31c4/NOitA+P
zkurnhE6nFPFlGf83JSQSILWZN4myEzRAzGJ79/lF+Bg3kw1zHpJ8GTJlOnRVPv0
+3wa2Ez1t5uRC6SFBsFsoPGxgnq6WoIIWlHimpWANLj8x1rEv/8HtmaflTLdYJpo
O1PS90JCpw5zFOtVOAICk7y4lkEWzkXKoWAkvAXVVfr0yDnaiiWlKCuN6wpHOpxl
DIDXYkIF8rca6jKETJjXyNAx2K3ZN6IAoa5iniodiPBszmp29hqL+Ri3DfL0Lco/
vZopW1aL4BAPLvP2+CbJtgNYqCN/j+l6g4SeYPUkIszwkvR1fYIIf56LNo7NDWmK
+qqDCZT/6IEFe3t/DzEC4Um4KK7/Lqs+f4Ro3jbY/+62DzB+1jp2wlHRuZsXaG8A
ZW9FRqJvfbOqFXUPhgQEocXTsrlDXoPX9ToM5rp1WxWnYOZOnffzUvUs8KMQcTAs
umqWp+MhGOKy3z4W62t73fv0xWC4+bsM0+PXGIXmovxW1NgOQWD3LMsH8d2BTZxu
IkmUcTdXiObA8uTmk+IGnPY6Em1BFbTRImBWvuei7BtD5UEAjk7w5gGzMB+rjzLb
lsZnl7J0A3SQn7C9kKmw7wtkeouJ/3nPKixLu0oPcs+T4eq5nPVT/dpi6lGg9bQJ
0Y6SxQK0MbQsHyvx7h0Effj1j2BJitTkO4KdZEU/9lTly1p3fSI+DxMbKHpV7uGQ
FWMXJvsnGuIZ8FfY5cwEjeZbLBZHoz4yTziBamN4YdRfPCb9RmGfFJrV2CU629hr
IOYl/f/qXAFfSrKgZpcABNTwTX7hik9hIx2Im0mpziRsdc1kQUOOU33yOWxlOmTW
g9H6+riMSoZr9JYz0U7UxubIHr/mOQ15WyR6z2jIBuwnPE6EJCP+BsNc9AKzuyxK
uIEVc3X8Kcn3ay2U5quQRi0Bk8gCp+asHM+ApmCM68LqDHf34UWPQsJTdOS0qA7v
74kkdr7WrP1Hl8eWsTv8gOYDu7l6f8uZoT/QD0ifmjp4fYrKL2AXHMs3gQyPh9yV
9s4vDa3G5mZ0l8b8bpU6EumR0nXEArIZJ73SSH7L3wO4ongJIGlxsDVjwFpw7lqS
+zzGN4EyBh0vXjb60NQ9x5F5Jd+yi8PKD0u1tWtimoILhhpUETbJRvE62PdU50JU
aVd0nk1j6blDkJgWQFfv6P+y7cxZaAYd3rGgq0DXgb0=
`protect end_protected