`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36368 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
xl+hxsegM9+gPkvRB6CsqXeGfJRj3o9GKDYCOMwvml/xgoyOArlMiQ9jCwAvCkBG
eEgUwoJzv+wiBgvDm9GGQGLdSAl88Ds2iUIIaj7rxXg/7Y1NTYoPji79rhX7Dc6o
FHPDaLJhhfQdUXmXbYJ/QGWkUc8d3unxqDwkIO8pX1lGc38Ybn7lHz2Ocw3jvEFe
0Gd9Ns4w09VynkSTBnoxojh9SzkBVwFxZrq7nRbaZVuGHmKnZM90welM3pQdCpnk
MtNpe7m8pzUicXJUubBxwBTZZ6/diHAGGX31KmvCBm9PvoQJtriP58mAPIFDlX0N
ZE2+fLPd98GhlZmFsotYRlF7fCYvlyErFbdpFd+x0HZXlCkqVlXiGkGVBTW8EXef
rlui/46ZDAn2w2d/IfT2nt3DtkH7xondRE9ga9TBh/TydeNQ5jvwztT7nyER1Qo1
GJYpkTClfDQZj3o5o7laVAgAZOuGNisFWVk/RMibXCVqCEgDjw68axTVtAy3Ms5b
6ShSnfRZPQqyHfG13F/fRcTbPo8K9VMQZgIb0RS+TR4lsgtKMX82kx8dANdKCyZJ
XEMvhS2xQyNdgGutnVDXPqNd6ZsI83MCiao7QsvowETTv2Gt/jd5aX5ud1RBxaX8
FkxvNw8ACL7jgbewPyXsME3DabO3U3Jtaj1z/GSlucMqTLFjfaS6o5MXE3k8uL1W
PdEr+hgaL37ZOBgWFp6v+A3dbamh/aTNxvoGMIDrOeY3p7mWP+aEPOnfKNVW6n9F
sLznCJgNlhtib/p37oD144lPJYXVxDTr51Eo/iB2SykbCaMY18dCnexoSOqlHwjt
zHL4oels7ztiVCJeR5cQQoMRi8yGecV4kuyB956OupzwGQ5TJ4GY2WjbtjZj2AX2
UsI7c4ZaY7EVXkPE98AgpWDDLu8gN9YewV/D2E6VbN/LUQvFaPx4U7nut/t6fY4F
osupfI+WWhF+vsSHcasd4+K2vGXVQncqS/3b5ezNI37TxDZfoDkz1/VburZthDsu
PdZNONDKJ3oKbm8z+CYZAi4xgKvYfBnHMfk3lozEjcw9P0lrQlrYiQJwT53izh7P
yNC0l2qQFN9qwXqR/EqPPR+LHx/7wV4gYMZB2BT9k6h9lYDK5MZnAeDh9r/Qr/p9
DuC2dmDHm+sUUiA18JaPuO/4hjEtGdrvuwpun0w5qH8oqW97sL3u73oieOvbsKot
t3NqszMNBsrwp84Hq2Sit8M7Bt/L3QM99kr9wC2Rwm+J5WEYORxaym+7KeeS51Y/
y1/eZYcI7Gw22v/4lNuzHcz5YNy62d3kS1hwPX+FUnWLu00rtr54kScNSN7DLD3J
2gnLHrkoqkwRbZlpJHCsKWVudBxCc8pIooSAs9U7LiecTiG1LMfeJ40nEDwKBSbi
bLhJIYUcXnUhrlfbtYoeRsa3y1T0s5nqZuaEFY7/Z33uaPL+PS6pd4JyvN2FuXTo
/kpISDE5JNnwg4d1mN6oBhLqz5sryXpAAsMF9ewPKTRupaa2Dqw8A2J9PbVOJoCw
73ehvS46f90mgbJsZQIgX0q0ZBEd41RvDp4JZLCyptRG5EVtFlvPcK2U3taCEwm7
W+NovjCV027+s891qrmwWk14k8nW1/sxREkZ7rRt4UXFDcdh9T//ICYrY/sN1/bV
grDnw+p3XBiwl4qrH1iR43lFCwV+pCOjWOG/rz68UAOMxaDbf/Pl+uHX8fjNzp8Q
8G2841pqDopNFBJGjPXvWclQVqXmBd7GGFOmi9n5lORCJhlA4LcQ2iZeLLsnSy5L
b/1MB/02/0uToJ4iD0w1OY6PzmfHduERjfDrD0/adDkff100zfYYR2uaEvYSA6j4
424gk3734tEwJDRPGz2VoBgzYHNOKfMNu+5wRdW33P8cmF3+f93C+u1y8hWNFUNw
4UV9OT4xn/xwxJr528p7Ldn2iUm8SwKeWK5MyCSRFKZU1O0nVf1HI085VW4zSTx4
i28uAtUPhewILaXaSUHlFgRC5LGc8Z63emvKbSp2MVnMJPQ+gys4faBRRR0hCt9q
25PTijTACdxTS7Pu0voMZ6rpNq0jc4jJIn3YmgmoG/gj/n5JbY/XA3FBXHIGuEsr
kKHjespKmyULRnWloZefIbept4pjZHe/vIq7tWTzFtXSuPd7O+tPG8KppkdSg0rk
HLe1q7PIte9AqMWzsJ4ZrEPDuEktkPYS3oML7fCr5ijoSxuxXE6jnBlA5WKxvANu
3jWoqksuJaUEKK7j51f+FTg21TIH44J/KPkt8kDw4ZTtQPp0sKPsApINDzaISvwP
ZXPIIco0rNu6/ZaW+Z6L2K6cVq7hm2Dd9GDaSHzo8Ioss/v5dxZwe9Uea0aczFIw
627V1rVfq4b+3kvJLDBZ3sMJdnzuDNjTngLtusEGnKeCV+cGhCIZrMwsd2GmwDjK
ZL03vn3MLfsp+kImDtdPrMrU7tBVl46p1XXaRiSRM5xI3Iga0m1rE5+n+gwmaGgl
CziTQGBT1LBxoaAxZGVueK2tr35HXvvxCTvv8y1voVnsAtHtrNLUlWrxrQVhkeFf
dxQL1yab4oUma6M3XsWPshhx7eYqeGDE50E2s4OXhExX+ZV89lTmButhllcCKGyk
9TJghUNaKhh1JaJ8WUPqwdfth2r/28+pbAnVrNL1ucSlN3nvHRf2K5u0hc77bzKq
6naGYybHNUZNgtaJk5c7n52QVkyQeQhDVmef62PNM0s72mncnJD91Mr2rwS8lrJW
IaxsYj0OoSBDNWHXvRNLeAmPWKz6BU6KKqAhklPuTcXzGUroatmd22f6Lxk3Y1jz
IDXZoHWrSVzX1oue0XLQ+4b+nMb9eHJ5Ei2TFOmQu8YXxmbAHF5oq6qGFz05+dR1
0/Yh7QFbYiiHvf3LmKrXVZk+ZsKxSfVw+O5IkbbPh9zKC5olOe97FriVDzjlDzLq
OaYTAqJ9a0W5bV39vO877upG25Io+d6tmY4mPdqWHwKgI1xTwYZitvJBTuTedSUS
A3WA9Y7ZeNq4ZmimYZh2ZhK1ZpxrXIk8RW41FJrPxSmDlRrvsbBpWr/m4/K1uxsb
v3z+5q5CjI4XUNDpmTwOE1283Lg9yXOIMXwkSQi2/2kLWLkHcQqJPi4LP26+JaPq
srPz6+pyDfgTRRMohInmfFR0jzNzegbfIxtbrJNWeu8XAYwQAXztUHEUCEpc5jWM
NYw2AvoH+XWzPXilc/c199dJI/RgJ23FX29N6bmYAUOJdzP5dXLB5VaYj7W+umFc
I96lBWTcO1B/CPQGoNbKYMQSdZwPTpzy/8pVESeB67dHB0ViRl8m1QGAbTWpYQSA
RGIJxgrYqfyIvw9bRKy0gUy7JPP0wCyLdKK43/ft8CCLe7aqKULXxBkDNVexPJGc
iHlS0ZRPP4YfHwH9nnLAe2fpgzGnjrCJbb79dSnuFcikRtt/q/zN8ild2/UviFHd
ciWoZV5RHysREeKcM/vZEdVHHQOejqkJwtqgFs8tEX8drm8P6vWtuv37RcGSpJKY
sBYJSRKr84Goz38ieZj75PowT7Ng1/BbpsWB2bXUlZ5EaaZgnkYFEyFLaE/oOUjz
hgjbrrhEZt2M1b5LJAwhFnNVTfOOISJqvGLa3tX2HWYwcUdNuf3FSONy/kGpTlA/
QH3NgjxD4eI0NFnuORLLiG4imP46GyCqYJ3sOl6ZgJmo8Apzv0FR1aCjoGjhnIgG
LlZ9SvcGNPNbdApVlEjDEdKpEZk7pEWA2car/PANeffe0rIeSrX1zYaUhx4TWGq8
G/KXqFuhbOG3VyD8Mrex0u1GAU+gIgZVCfZCRFmYYhnIyhTnNpdVdZGUEsGZbh7B
TwPXC3bmNo4i2ELR1wNO+uDIxpfyykGaBq9lsIiNwbxVvhfaC2XFfbIOFGOlNkox
5KdRmOgQT1gUCURoJ35rNHF6+9dvEyaj1aiit4ttb7G8JAwSSLDRxyFSPNO/yw44
Tk0UrPwEuImS6h7ojDZf1fI+wE5zqurfxzyFheCtRWB66K0mtgCgAXTBYlPh4owz
qmlYYPLyeIFi9w6KG9/AjAhAYVxdLN+MR9aQ7aYpfBtxhzPeXP7AQWnmXFDwEyci
KooG5ybAhIgUDvJmzroPLKPTUS52kTKPKoUbn+4F9dzvcWEYmd9NjScxyN6IgGla
jKrxSXvzcfB3Xd2/glliCPQVUE2e1+MZFsOAPr0NRy1LQytUgiDsO9ZLIYF+qddl
MyWr/GBidqfc6wFJzhrMJn5lpe4VL7izYDDRGSFF7fNefbISlGMXs/xObQgrs/54
b1wz0isVByjkMYzYpH6kGmS7bmfsFLHXlCVLzJmV2t5jDjUKRxHa1Hmeav7CyPqo
5BgJHFbVKMsLbuHRkk2HKaXgdJ+JTDYICNEEUP47n45hRwEwZvO9DAYuCFlB6T/R
C9ylgPgesT2KBhhzZPoixl6k9FUdE0b0FwH8zAUXPT9BLN5LhOHYzfskLYcva4bb
WHBS2rU/IAdWlbbjxch1OU4eU594tAYiCX0EPzq5RIiqaOTFJ3+vKJf3nASNgH7e
AAHcNfw62wUed+is3r0eX77PSu1Iqc9V7i5z07kQW8buSNZ11g8x35/Dik0Pd9eo
hdhEN7MPT1e0GmDlqqT7AppKyo9g/TgQ9D2xhyrZdIbQ+6QIoASS6dOQ4EBoC2sX
VoOmm5xzEbMrtJHz85ncS3PeHoewmnIYGyIRlEF7338usMjiL60kmZCVayj0O8+D
pD7d8yBLaaVhILN1ErErbzHE1cDX2X0niASS/qm94/7h5QVJLuDiVWNdYx/cxpas
DZ9YqpTnT/pf848ujgcUWU7Eu33xxMV0Z46l+s8oa9lxQgymqecK6pqH27qQJbQQ
t7+nXk7TISdCUTNQA/MIz0yto0viKAKfxa6O00cMb9X7Ln/FWBFrFOeGnkB6CDNm
kCE3QE2CQX9sDo3gzucA3vw57odJ8VLAIqRWJDzOE50j2fW2RoQREva4KodcVRPO
iUZ5nRuFlDwUDQT08AB34qA404+rcA6WguxdFMyXWgsrQFv5ovcLb5UdYD3Fsvj+
yc9u9VMy7OUZShtRoxHIXEUIbN+DYpziEXfoo8GltAsMAzABZwjwKxF6eMv4/Qil
RAh1y6sFh6FIveTxC/G9OH6+UP603ovxEqVVDLTN2R7AjzgTebUW/4PZWA8SwsbI
8stdfMRYDDZjndvA2Hflr/EAWNxJPQYxGMHwpbQyUQxn6bADNOn80L4rptPGlmUy
uCzgqZ9juIcnclRrJzX71ERH+sh0oP7AyJdgLlN1wdhEEOnmkFmvYHMzYN+0Dm9d
eQb2IGYOAv60MLXMC7sMT9K6TWOAVvM6E+l2OjxWdshez/EF4k5imScfHmgh9JU8
7hRy1F1gGZJk6gvx6dY17BI9Uj2s4ZNx960vsZ+3tuMLgG6BUBHXX4+gMGGOUlGV
psM/aMAwYx+IIsPZYJV+fo46Xc60hI+kJB5wBKOdzhnaTjg6vPKst7wf3FWbPjXL
4L/CSPgg46LJi4b7eUjPAw6UlmJep1Q/NVmktbBOvhRYrbOEgvzg8QECjGId8La3
KDLjBYb/n+nw+DZclL0JdkSvaBTLAeEHGrvk+hfQYX3FZW8Nh93KYW3tYln8XVTj
3lQuFMWsPIwxsxGU6yHtxnon1Mms07QQGOivAgWmL1Z0sLeqJkLPSq07UbYM09NJ
D+B4KktDn5Bcpu2vMmzbiR5Oyr08aqKeyNkqP2Xck5KXcbUhXAWbSjT4btJbFVvA
T/5gAHumiAfNG2E4Zed2G7jxiAY7w14R86Td8TzaF6IvLQKfTq7tJkKb7k4ieRNy
oYg+ZgQE//GJtlbd6lZd0t/Io0iJjbCMNLVrceiqhj4VV5BQRlXWAw1XIRFNZaqT
jDfYvZ766HdFNwJZgiHmcTNJpvQNEQ3TXrSASXeJA0GufdsNoTrYFvqDII1yhoqP
/W30ajxyOSKjqliMX7TjhMumfcQZE9zZG0AtqKlwL+I64gr1WNWu6qgEbuq0Ec64
ZLxlz6yDghpoP6qaXpsYY7f65CVOW6KvpYGOor4vrH0Mnt1kuQA7ebZfXOmsQf1c
gHCX+u37xhYvChE7fj+CT9uqSA/q4iQZzl5POsWdkGtWY1H+f1O1kjwY1lqcWU2q
gRZLGVGGlfjI/ojtgjwayMSnaoDi11FYwWfBQa5nKimCV3GX09GJyy6GWN4F0sGl
V8btFOYEhiAz/+G+vdqpoM0Crv4TFXuH1j/xVOog9Xk/UwzwUJSmb3rJnfh/M02d
sMLnKGo24HA0SKhL/dehh4z44zmmT7AyBXc+L7EnB7l5RsShjVdcgJvx5JgCX3Qz
ppPOcF9A/XlAIqNU+9iebjpLHQn6n662LCh8bvr5Jqj/TAV60iM1YPEWiwEVrvht
NcABJXP75deJ5TI+yvsA56sNyNIISCsAl/nmA1/rjMUJSAmadEMU+aN2n/jt80uf
uH+uZjQ0mqmAbgULMNjBBf40BPEmYENVSMaU25mR7DdzNWGRAlzUKjrr2/nlR8p6
ek23azFz870W002VqTb+ukRpZ3u/e0hv5McTI8k5ZoR5OvRdxNxUAPzCLhnv6mjT
J88ejrAzLO6a4AykFUqoaX9pPXKWay67IDHmEzZpBqNjvQxw88k/LqqJ/+EdVOBS
yqnV3DPL2Qkhm7/tSxVRx08ReaU5qi9wmY8BO4nD+l7poazeJma8XI65w3AJ/FeX
2Xe3nc/TwedkGvioK31iHc47VDvV0z6GTo9OrrFo/AWtVQSssf1mkmT/T0q3BOGp
jrVv0GkbGYKoRfC3bNQcj9n5EIQc2u+uj875hgPV0y7KMJvqTgYMr5nOt96v6uCy
ddOIjJ0Og7Tiii/PsE5FDiqxx6wwlzktY+0olwO3AruZadHx6d7RTPU/zOvHYP60
c7g2n7Lx8212YBGgl8+7+0Ud+SsuvNwyYwXu+vcOAIa0gMddqVsiVwERw1bpaw6y
rqa/YhaptlFhyWODjCffemIE/9epNpon6G7j9U94cCphA9EjdnC8Ql2gJ/aH+p2j
teSDM8d2LOfQ7eGPm9rPLjoo32UVbK8/WGdhn/c7NfbQkbiA+zAcWVrv1Rw9tPWv
TPdc0m+CABq+aK8uWVlZo1faeb+slppH6jcI3LhafEEO6qaSFnoHzKpUBcWH9FK7
v4rkfQIvi0mnqFYn+9DWuR1U0xduvJikLskfbxZEgfsXq/AYxSM93tiFaZDDPIey
8slyV1zbQSp6KNhkDS6oJBiLQAPYx6o6pMQFyKpGmOHGbmu8XHM0cBTp1rtf9vR8
K3eoHlCA3KV7LzpqdTqrYwbfpByO/YWy3pX3UM1jJOjYXEEuZsT+LfOTHPSrRZ05
j+zvxtc2yYn0mEZg+FvmHIL7NZMG/QrnayAsnEVKlaCjt3cFElMJt+9KJ/lKf7hU
a0T3Pw34w1VtwmsyMCToRU+K+BWo0CAFhI59g2i9CYm3SbjzQ8Jg/MbqYD/y1mCd
d1U1W7cN7iohYAl46Bod3Isc8NQFZtCuxmaaOZaRmWKVMZbbg+oHdnDMGgehqAXD
mIPzJOBSyQm1P7Dim0RTJ4V2bozTkGZenesIrup7scJvp4IsCzyEOioBDAhNtf0K
uaSrVpKsEKQe+vwXg//dvnPfrUf/QAZHHr5iQhwc0oKOBmA/oQEbS2VM4bSCYmyt
UOUvsRhk1mm8XZ3sG4eA65spVtqskL+KFODbQB0X65XE3HThMCxgbqnGsg+EJUo7
51eeMsxTZXeHEzo7Ibt1qFBInk0uDA1j01QAsnnV927CkDPeOsxJEPvw5CdUsfGr
ztitv6Hv/TXK5SpBYcVCJSp8UtyktyAuSkXXxpxz6Jp4V5CDDFoy8qd56oodwyPL
/expe5JTtFe9ha/rBVi8THdh0dtxC8Ol/vn8T9O8XBXKMvH01go+5aAlilNHN+fW
i8P/PACIMTklAouBodQ6yHfIy5Rgg6ZVpwF1TZBso9O0xh2KCnmE/1zbcDuzWH9I
gRbvK79qrgdlW+/xBY6kaeYOo5Al5z+dUYy9dzXJ1J4dV+F8Buw9U4XSU3AXNLzl
uQIw7Q9EwTiRrtwBO/FMX57+C4gD2fY99OkSZ5spehrzCtIpf/UKhbHT+wJTnEwM
zVeiwKgorUpXToSlCEHcB8P5PDgTp/gr9nFaNBfBuwkw3q+lXDm4hpJ4oXc8c/dW
T7wroAzHxk+IsQdo8pH1IQgyX6N4o3Hh9xmIYoytVuMG73uCNn8y0VVTLc8TDL+9
pKx77sS4VbL2N5CS1J9XGxS7hpyzv2ceYkpkeIrT2l2X4QM99UtMcWFwH15UVHFA
DPtz5rsyDbvK09xZx8RDjbOGiySpNVS0c6W4YAa9TvaZDX/C2TgcxVXwSby/plc8
cNtQhRmF+zc7PBEpxgIOgBXvrGBVjCWTvwX5eVd2f/eaYK/CsW9GqKP3hnjs0aeA
98SAqIGHN75Pi8kiiuLsPtiAFxnFakz7kOzEp1eYvm/Vbm2quISzom/LX62Jsv1x
/sxNs6kVMTUE1b5vC3rEvCq6uBSqzv/6lQovkU21y5YRebgdew8uSHzD4q4jJUBK
2v0XfZSmAk/terY7zkq8yc+La04u14HQxiIFBWNuc+bcrzdUrZ6hqvKp3ovhfiZ9
V+gZ7jqXaAXQkGiNqugFYSF7OPno6Y1fwB7rpl4IXYKihDT3Zi/U+vu33dMjBL/9
JqdTeqszpxhewpwhyRmIVEk25NiZ1liOVFfGNqUPCdLrqKLiGyjXg0crvz+r72W0
j6sSTKWEDkqFphOsTSu7Xu2qnY+y4xHF0KnepUzWmdBlVDDk/VzJgqBIjSby6Spc
N2GumL/JcqfD15Vo7Bb4rGgoX0bpGzoN0x6ftMndsZ1cnFwohpgpuZyH1VCCUj/o
Nw7EVNmvx+NQISZcrBsTogWHXQggwpjcdHp8j+SlOBFkIZIYkqLk2tKbTudgiVvi
ZlEMaYZrCir5TbgqQl0cez2PHkJivsPDNSs3BF52VL7CtNDft9w9e0Pckf8l0gfe
r1xJJzoHzkRPiMIg+VsKjhLAi6N53gDlij0R8ynCdG+pNmHm2dHOD7Ir7AT1ZGwf
BHXvjj5Pq7SBzPp50Gl3QpmA+gV7bahu5DhBHtLcaOygrCynkKcq1XNww8zUIIOU
Ckl5H9hs5ENBbtGCKAVGWY5acG3K7UBZXvRR4HmwE+Mt/41c6qcNBj77sBGNqX/R
RCFOP31Vqghmzs7TgzCq+BkSOHlqrwwJi+iSltz5lLBJMdTY2pFPWUt5knMN1W8v
striJnIDbSMfMwVxCELH8ExhDEj0YpoKYJcyr2Iruln36J3GXNSPbwJk+kenP41K
3RkvQPt7B5CYdl7a5QhEIl58dX7lRCWrYqGAYPQ39UuHBx5Lgen8mngksTrso3/v
1kqewUbH2J5z+YQOU87+GylgOWaoESv0oOOhAWjmg5eya0b+SzUBvWvSIBtatvcb
TWQbZT1dlf9kqLrqpHOXbIT610S+MZc+JYfsv4Pk63dYiClbHNAH1u9BqShg485b
7GTUMrV6LjWie0aX0jCkNhYfTbuvc13ynE9gaR88MqrxB6EE4VEvb0uIeor92Gw4
6E4W+hPd5An0mdTqiEVlIDxLrgWwmGusqI2ozv6i0roz12Vk9khXVUrohMlHTVsc
nhLlTnSQaVDv9PCctrfNYn+2rGB7KaDr6wipskQYtIVsb8StgYy+5/LREam3IPcS
MBP7an4mEQx3/Sl460QvJh/op6UWRK+pNdolQydXFlJG1m9056xzuQaCvYKWhH/7
p9dCPJ021WvRM3O1ht/ZOEMykzOaWklXtcWi+4OaCqZ9YgXEdAhGlHDIkAn1vWG6
ttO6haYN5QfGxvhEHVLPadnCh4+4xqYtAnOEsrVdH5Gzx32xdcOzDW2jdxp2T/oA
lH1tw9KSkl4K/MjMmXNcVw7LTPjWPEiuKvZgzONsif53EmF4T7o/VKqFF4rQ08rw
wDtH6dQlNtZUZZS2Wz+/BjbGr9OOpQDeJa3G5b+Y7At1FvYkfaVqemIFqYMNe5UK
/mzznGYSOXj2RXHiOVmQHGxEL2TvLq40UGSSAyOkTM8DIT+YJ1GsNV8dbMVE/SxL
rEY4QxXV3nxennvA5hUDbTN33wq85Vc7hTtZC9cgSaTuAdk13Ap4Tq2yC13kubLR
WrGfmpLOddPo16WxusU/IN8Xn1oEBSnbST6WnsdZUDKlfWM1+GK0IuBNOOPKoXyi
eIywoCf8AgugEbHtZjFQSlKnx4wp4agAGmizEP5I80wiE8nidf8Pzi+VML1h9hR6
ngV4J0ZWa6e8tbK2Er2fhBX72mkRfpdxmCe+VX6ZfHnG8BlppCo5e7cOzrAulmp6
6agHtpRBZxAMWHrZc+ypBa9LsCRzKx30FOo8I9iN+Wf1euJzh0bfWiDOVWc0kKg/
8zP2eQSNvQwJET8v8HEv3QzYaAo3NGC0P+DgfN6oAu+xTcGZjtzdguXcVev2wJiG
9rvXu+4MWXV4ywIPolVTfRIn7u+PLTaODz8zuVMAxJE7W6fa+j4OKVNYzVTzsewj
DAqEOgVo5J9N9QVbYYlbMO1DX7F23N9PLydsgsKfZ46Z7QUEhjIgR+ntcixWTw3H
x1tb9tCar590jHj08RFtRj29EBIoUS1/Ke8uUBkRObFShw/ylCTpu8MQMAyrmobD
50eV/WgQQEol97qB6I95XEVf9vKoqTIj4sQSQ0k4oqd9jm7eRvv1LHugvroidFid
ohdIZssH9JkRRWd+poIaR/qmBmEvZsAXIeLFuR/Ov8VPjFiF/xz3VAxNT6sQsrWP
U3+iCeecKvggDP3jQ37X0iL2x6Yq9HJf6MlQv05qoptEcKppACCEVaHAhwgP60ZM
SeVjOOiR1MdfW35Kyq3ByfGTlfqk9MA3Wj/ZvHofC1SlrXupwcIU4ZnVBKpXWGyX
Sbdl6qr/P/C23FEGKAu76Fu5Q3FS6SdybMganPY3KP65GpCxcjxVBIdTE4bttwQ2
1yxG3QhqM3YLqbQJTirr1CghthWQBH5+EQPpDkXPGaoOnqyUKAGbmx1rCcNWDZvL
GuFqyTe5liuAvIyFYTKCPHcXDbUqaWm5rJ7Es3U2m4GIZ3ukg8qrbnF/ofCyf5Xn
hwygvN4YNZhfJ65XHRg/oXw8ow88qOHU0eC+5ST0EH4xVn/FNaQXUi1PU5oQ/Ffo
QayTVV0y7hrHHFXlQSsDIJFPIfVRdA2tnbWESLAEXDuES5cFrd+3/FYVIViJNYaP
O+EB4sYq3PiCYicWkvkus9mrlObrIvkhpN7rfWHFq3ZJxsiASA+/YVkZAnqGNLI4
il/MbNlN5un4fM0joPLlhFZmaWSdQCon8QPAlM7ZtXbN5xk2n9tYIcBQdO5s2rHh
Xn0l6ZwPkCGR3zqdI90MmeB3ghYM3rtqAL9dS59FsPGUg3hMV0YdDHNqnkA/qzkE
7qoxQxrZmg/XO0+xEQ3rfxYOLFP4XD7OB+gR/3j0oHgvgOv6X1Gqac+awyczI0Ig
zxrck2pbB1mHgE0bazL5qd3NU6dFdNDpl2Qm2IjD1N98SWnJdJIOUX1OAHCTPyxV
nn5mgDiScNKL3eTPs4vToefR5yOetFsgR/bveYc9cw/EHukXtGhuWDyl54r1NvwF
LdXvLH1MSwFeoKw+xm2riVDOPXe3U50qy0uBE0c6FSq7ohtxgkiNubbdslcETmBK
H0dtgaDOVZN136KNSNTi7lT7D4zFGt51UHN/2VEKvySh7fggi4A8sEVpef4H9U4t
jbWMUnrdYjmw+rL+BtcNtBZ0sMcUenZNyl9GWLWjJD8Z3DfNt6Roo/bl98RXFCJG
SgdyAS37j/4L+wl1vf6PS23X/IffJSkqrxggyc2hTrj7JP3IimaD3O5HL+j2ambk
OdO0jf2zdBFNE1ThBqOKtQkohlFGmyKAFaCcG8RsG/tZS4Z7pS5Q2Uvw5t3KXl0h
NPNMNq+BDlmlQPfoSEBJolvOm8iTb78w4h4q4OXhI9OFVQqULLRH/2o3UVfwVQX9
pHtTp1k/3vCl9NAHxugvmcKvpnK/qnyNyE8J2xPaFAdeQtq8MJm/fW5EBqTO3aUT
qLSCxgpnBp/ifZKXildJhwgJU9+pZr5Y4XHEIjAvUquzlbqn8cBKjQN4GyENqwJn
hoauLDjLPcU30QDW5/RGtTByZeUDw6B8hOmUiBgNQQTt4uHc0k7L+pzXLoa9EfCJ
wWpoIefh+y3kyXDjvTqW5fX9hiZpwNv7eNunUfk8eU1gIWiMroGzwBpd0p+UHaEU
dQBgXB89vdQpozZMhHdFgBRs6hteB/IDbZU7WJbG7x1skW5KWcaRWaEhpslztanJ
CWDTxssJfqkoQ5JV0O2fFIB1/abSjjX6DrOYXT/HYwDHXPCH+Ee5pX/ga5sTX3vv
v2tU/lullo6AnsiJnB2bl59Yx2wCtrQVm70syqE2yUG9yaseC+uhHYiY5SkQLnlv
5W5NFpekFZShdJX/2Gxz5rgivk+t5sM3gZ8hSXJlb6O3viTCR2/WoB+255seHYXy
uj57/8aj3Gw+rPdHIwCL1OvW1NVqoBvSeILRAdmIlAwKaTDJ0nJkSwdmxwrMaCKh
kVXVy/T5VuAtnwHIeqlyPe8Y/tk7sKWqUt7UmhzVFcoA7BxikI73Xqp3piMnpeC5
8V7L/hPYF9Fsaz3HiS7W/9MF1tIjF90YUz8TDvQMIVLJhlXbJBH1fqllvcF7eJE4
UqKiBpXSvl3L9D9uF/1RhphyvYV/Qv3Hx8SkfoBjJ4SJtOvfEYir8Ieap8J+Mv3N
yoCB5GJNptlywkfyGNDeP/j+OQRq1QveFy03L1s7wMG9hO+8jA38MrS0HaQ3taAh
1C092MxVhYlxdUk69tMscrNeFBOM3Xcqsch2sNWpXJXLJoLggKSXF0S3coGrF506
TIPBpEZHwfK7j0AA9JnckYC9IErLL53oKXA4HjBZTc8hUbf89ImuSX/scoqmrvxP
iGFTg3J8fMzcEpRPmFJED0/2nnowgvHVsdXvYK+OhWicvP2D1aCGb9zyEiLuy9Df
iXhWK94cPL/gGSRpK7KwsaoEpgFTmqCJ9nK9/5CeUkVT5i/MVimX/vNHUzzh6jTj
zezBfD7pfvZN00Q0X8NPYkR9kDu0t0YC/CcGr3e9li5/1CrJ3SYsSKmKlJheMbCp
xKqjQzbfvypVQs9huwdAXFBe84WHYEZ0IoXta5LJhrLixt1+A/Flg3TO6DK7EKik
D7WPUmQoMWcDVrH0cm5UEwzLQi6r5n/9uLPxkhLT4/AWvIaz0M3hOVRyRkzGUC1H
CR1gpECOkLb3C48gccVkiO8kbGCVjJOACtxshZzTM6YUNq4ZoDee81tH5Wub9ZiW
KFTwoebxhoeycH/n+kC0ey/A2PbJpXY0uX+j+NCrZzdnpdCItG/CSEZwm33LYJYx
unt4kLw8uAQ3+kzEg9WP6NeqY/7bSQf0dpjFAfPa7TAwSiggskHLwYx4vgsyLR7F
AGApBsLF2uK2t+j0BdfMbK2UpQpyLElssGvPc/lEo4qe5RD/VqqcIYiK3ybEjHa+
osuvlYQb0xJA2ilIzxv7sRxvEooT2doKM+fPyxadkPNraMia9XON6Vc3F1oRbACr
pijGgOEUFnGX7+e/YGcHYYQXQNJ23+CLYbf/Ib90dfEIqD2cH6h+qYYPyGTlibVQ
9kbwwrl9rRaP5cDo5rUepYew8nZugcrdD0s9IDMEn+zG1jY9kA3+AopH3KA18c6z
g+sKoyjrSwmyp/lZrGGF8Y4hPGdj15WfVqDNMx1FW2o9pqHeXv5hLiCAex7RDxVv
9fNm+MjosC3/vFbcfizrZgdR+ViXC01wzT6kaC9l0Gomii6uY16YSfIJsUnFbvhz
bc/N7N5qyxwvOaPg7hfbTwSlqwGnLm+VdqfAaCbBGfW2bAh8bj7giJ6S8cVG7IkV
xcXkn8Vk2juHr6/ZdNIGCjybu5LtRstF8ZUWSmsfaoODlOyAISvQMgNxaB7qRGRo
xlBKNUZ35D9fBB2cpO9jQhXKRRt04vsbw6bzJyZiOm5YHR/YKIV3vvCpKX+87iGI
aDa4u3RTdw0UZC8fCf+/jlShwvMfFEaH4PjooZykgJrDBWni981/IwnMLrMrWGi7
6euQURPhlzNaHo8ZmesKx97QKdaUOmbU0BDZ5hQWoh0GsaimrQ8MVStg4nGE4IrN
AYKOmAqALpcy4Lw1m0SrBPggpwKYSuPJYyWFY3eBrNRVbDfhdAH5W/tIEKMM5zQ3
rmQtpNacRwpqtckCSXDM2t/BSwD5izf+8waTlP6Oag9S9znqYgAgMsepHF6889cy
lkZ/nP4IWb0lNnZ+dKV6FqGwxprsOrfLq2Ksfpl5tC7anHBuU0C5aZtEfcwLtESS
DC3LToc7zjBl6MYWYylk7JMLqvPbXERKwPO5fIvUU17B9RfAGuABW6Y4fjsxqu1e
9D8ZMLOM2YZDcz/10ixeakCTrPwbrmRAel23SmXCRBW5DVMs40UHKYN/Oj3IrJxG
IR/gpo/L3FHVnMNIiS5KUO4+pTJtshpJWji+DudO3CO0Gpc/LspqR+s3sztGhzda
5/VUsP9KYd2y2uY5ywz8Y5UFPZvcR1YhQKOqwUgda7/LkKaGf/xyxMZQ1jyK0HG2
7DZ8hJGfTRlpskrJ75uHakEn3zaxRIbfhPzWV0mhb/9jHO0VzFnu/H4KWWMgAMmJ
F+AtgriAk4EVpEigta7a4tvLIFU+DoHbK8Qj/3vVpe8x9F7PF/xiR+RH4c37ZrR8
aSpSuxRhNydIlI6q5PxotGsR7raOQefcXDCKvVuK6BqQj2WJVjpx1OjuKlDNLmOo
JQm5r6FLfQl80LHXHeOYQgwg/DUHKttuyouffWZ+ZVxW37fmoA3Y+vGvBFaT4ym5
oFGzXBlrhuVclWV7zIVR3Bpx9SfFlN/z2OWuqXwcMUpdJFjXKkaX2MFmQXCmL/Hh
oZwRa7x4ne0n23oC9b0gH5aqFKhsutoOhpUN7WZXHBIno4Uxa9qxscSgHqCObX67
Hn2CNL1YxrKHmv4766bvvD527RPiyWCOJE1HQrHO/VX7yuuc5E0777wBVLD5CEFi
VhVmLNxl7X8ikOdas78mG8b3p4pA5DQov5ckAj3JpNWKox9LCyELLSmsN77NUDB4
R7H4mcpy1PtZhrwXU7he4LaLFs+C3GZjE3cYIaYE+rq5i2HiPtiLWx6cLI2Swi3J
+cI905XNXFtJsa/pjWrQNG2Ue1dUDFxMvRbYnPdecJMlOKJrLHYVBxEO9UxCPKG0
GwiDJuU7YHJ8ewaWwGr79+svpsiqITvUObaR0gkm4AwHfR+tCyFdE8nj3AfxwMFu
zdRAlhUjtVHag2XMZ8SE6TC5EKucv2yHR+Qn7h9FOZaw/n+PyH5bP6ZFYONOrzkI
RNp4rA5GBrBZqIT/g0lHi6MYdMjKJbBx81p2k+06CRy/h6Jhm6RyS+Ki4g6VPdZq
FesoTDrd/FGsfqqYM1YkC1Oh+Cpq/Fr3mWhghe5r83ac0cv8zR20696Xioq9N1Zm
IqBUjvTrFmYGsxgKeuTHwCOXfVQTqwnbdG1ZOpJ/2NHMAeAtbRzbl1L1F9YC/9X1
K9KaN8nIW42VFSNTMB00B0UbA/xZPmqsUmt0mPpptO8pHXds6F1X+9XJK3pxIj8u
JMeGF8L5pBqSP029RFMs1S45ti3QXCnJkNQ2AsQL14ZNxvrvSBoYzgFt/vxungRF
0BUOIULkXunYGy51xZsFG+e8JwYFkSa/X/Eai00OxEOazE0hf+nNKzvLZCxAREgj
nMnE/NyF1aubXbXyOSamTdxvpqgQ8QSke6cpJAwxojOfgpwUZFqJ1aqb3vr1gFmr
waIyMEKx5x6rcgkLPmcNVFuuTT9HO+RmF/zgBzhs+v1R9/920/K9bGooClUwrCmz
sCGXg1eXv8WxpZ4TMlV7QwbyjtnLgqw/p/HxN244PtSArWA/fxNORreLUudJdQPP
nlyqJzfsmUGfPsmZlUxLbdwM6YQdB7HhcByBhzvVvPFUxasPTM2mAqwvgIWaa7Kc
sKEATrsV0KslGUpB4SxMkh5xArlbqGMrWxNo/qtNY1BMtwgDsKuCpBBdks2jqquk
vme6ad8fkA0vzwjSFW/fdLwB/Dnxg+Xc6BRxq3SG5vHS2W/DVF5MVwIKLXIYUkOg
3GnSAOpnjICOgZWO1O/B6+6tjOXYXId7IHnVyqO035Z0i7+wqwoX3cKCHwLWTR/f
/uPDmKTKPemc3D2kp885J+9cn/gPo16rhK5yzgRFIsfs8YzkgsPJ7ivUUjJSCwZ6
dHca0kI0IF0wokNnKiuJ7MSkJQKzIyjShdjZYoW2vnc0mhSjOiNSsBBboXzgZxuK
lYbnjPeOsv/YAwJ5vs9BmezgzJ9DlxbSkg3E227RMcvUkgjHLWbs2G0QRzR+IGVI
IFt2uYfe/gmQQmmw8TxIPFl4GMnQlTTukMLHA6v14iMvQa1PkIWiOU9VrLWWBKft
4bj254Bd28gMScwxYUmWrNfsmGhacRwtyIspvyv5yO0TMz11B6pWa5AJP0P4fiP9
CXSEb3Rc04LxzMxXwPi0vzG5399UNmjjcIirc2/wz2I3MhRRLTEvuYu8E7IttZm1
MdGwPlCE0RGzoW8wTNJJcITukULfBUBC7CxRfI9sksSqmFZPWH3sPwnUbGAG/yvI
aeZHzni0D7OraLtuggmbFCJ10zDZjC99uULYOAzCc7khpjh/s+PNo5fH92I8YsFy
m0oP6026ytEciwL8OGpqxNjBxDvYzyNsKPC4VY+9uXpvPkmJkQ4gscEFJTzbNO96
mlbR/W4dugmPoqabdlZYWUKQQQy4kNpovRa3fZAyHiR7T5SORfrY6lPFn23UX9Dh
hMMYJIpn7mXrFRDmb77E9CE9/5urs9y9DBuGA3SQR9KzQ/lLYZZEAYs/RPC/aVPA
25XVhrWXFKgvJ7r4vMuLNNzYtgO3BzvE0nafNbO4ao5epeVCXhT8s9ksvpHyVl3m
zKtF+neKpU317SXiwCQhU/K/zic53PJ3E9Q3UdvY6zzs6RgV6EpjqzuBBHgsdcKW
Gnk9LHSJs6Ib7lasH+gZ9NnICOMQEhaVFuFqEkEpWBCICr71EFIontGm53yAXKvl
NJQpzW3Ig2B7Xs4lxzeLJUdDPIoQV6NJ8Y/3HcRFxmqd5fn8nLQMQ6QZi7gC7IAR
jryE1E7X0ZvEoeqEBza7FEHoWT88v8wIZrQ0yOsqdlyoQQnEI5DLZEhHSrzWVwms
HPMdADdvZCdH2lHMfD29F9CuIulqPXerUU4VIlf9fk79216NYoOayJ1lvxIfA8Hy
ckYplbNChmrO/04hcRLxJs5cNQr9OHZ87TE2k6pIB6PGkR5ISsM5bMQHaEyATNoe
Z0ZQWM/POU1QtKeviQ/okelApq5a/fSmC5RH655SHYGUo/Bu7yK8JW3O6RyPxesz
lYqJYfPflF4haHj6CFx6NYyvhl1YGBdUn6w2V4QGzvo9sd+X/2RsNegGUewfp9ii
WAMNTr6IVggEN5/yz94ZVctFyVWU6NUSO1FYqBORMECiIqXz5be4qEhRuiRZeYty
YEjkc+pf7YVhPmo/mx63590TaHCUOoskZk5uv0dBheMSctUJHqLjxPlPqCeAkg5J
pSU583NaNv3ki71arb73vNmLylWiwzD4Qknxp3rt6+zm+ShG/nPEhBfRJqxz072X
+/oX3r5sPIDurMMjKwnKm8Vqxp3RD00y6+vGeiBcwZytMvDt282Aevy3dyTZqOKG
qNpOZ2rP9+QUe6YvR/8FR8FtzHCPLHJ6peGgfB2KHqI/qtH1Bp2HroT0aQ2zIZaC
pGms+7loFRX+YvPhMDSKno3HCP11Rs/tl3xGujGzlqASZ5LLbCp9B1Sy7YdRzqn5
ys+b5Q1S0juCHRHiHk8RFZOc0iJUhpBqWbwGcuFG31PC677e6AybUHi05+Qu6VLd
ljlvWAtGATvqkcYKnTVCY/CmBmm2vIcWNd1y7k2/lHPaqXZ1JjHXboVM7+VUH7gj
XzF8IoJy7S/pfCMxZ+pzfweKyQOHS3Cy5/XEkdFRUaLbtPounbjZCNk/Y8lqefe4
8UkaW2u67SJrLXV5QoCRQDrUaL4K9O71+rrypkx8gnKFRKC8TmIyR0Jko/jlL0iv
PTKhjIHhSb4ddZ1Vm4oH/IM9UuhbcvtMdBIYXGqwYSg0ykg2RBMqXQCYryH/pRtN
rUG10eyRCc9/Yd6mofBFRrwKK1QznjrzOpgzW1+Xlq8ie8yFB4Z8qHMNu501U9ZB
szw/jLQHIVU/rCL5m2EEuFbmEuDJqstaoQowQ+zaidScNNtbiWug9glzMcG6zwbt
uuwsHWbJ0YhGPza1roXEYdiYypWz9LhbpGm4XDr7UCjV7JQBmULf65r5g0U7TJNr
LBWHubZpS38lcPjQ6YvPYkmpo2RIQ1Flxd4hKNzY/hqOp1uiCCs51pA2RYbUGZ2H
Fia0TQv5bQH7qHGnSZHfIkv4o+v0AIgVLeqbas8dXeZdwdttMyMTH0iTGKfQ8Wlq
97lPtWW5vNEcmiTZr/3xKCqzG43alH3wwpYDdQQMIV7w/AFZkBq3gPtneISUoRUF
3ig4Gtb3Rj7LFOrBiP9neCjozxy0jLXe/EZunGAxwPWM1InEjz/zAKpqWlsOWpLH
dTm3+tVgpOFxHKcx/sK0xAO7ENdNls5qZFiL5W0lcjRG7GZqSya/6vn8kykgEaCH
TTKJMJFGymRYd9vVx/itcgbO7NTscpWtOMUhOU1j9XfoVnbY4kUkhOqb74v7JFB1
amG6DAttNjoTdLCGZE7Fv5D7MFp8rv595NMjnHBE2VSPbuxhvx6PmWponEfHVQHp
k4q67LnVC/h7KpBAtnR7zjSMEBNHQ1vYaM7f6x6LR+tBqP7Q3fbMe/fbdIdih4wb
7uWtc77qo0zdR8+ZOJOycYfTXiTJgqx+xWjXMMM/5890Mh8bTcHBfsxYrZB64mLj
Jn+huBNGH1JMPiSEIoTcHy7US/aFdloC/56SGNd2yiQ2fcR4qkR8DzV+VLKWWDWm
APyazzejuX84CZHQDy+jWjnPK4Iycr1v6qYVQfIXBUfnbffm1HnhieaAS4WlNpAc
V4Fhw5gxKX2INrgRg/hZz9t5lRox4ZS6D1VljH8qCvXYt0h8NU3gCkj9yB448naF
mS3LtPuUazVdvRa/3W6aOq4P17AYWO2GuYhHH2SeGStrgtQ80laDLIJ3zYIDXkUt
lRR6eVsVANvWHWmrEogDClqVnd/lcXLLEaEmauAyczWHv+mLXAm8HjXEVSqMDVn5
7O0oAsaSm9DpHSfPwiwQNM7eW+uF39/IcKJXA20Kz+lqRxYSxsFNQVrmGmAkBb3F
6+BqHJzfbRyhnGLxFLlY5vvsgaSrZQRqH/MblFDxTKq2Q0KeE+XfYk9wOK6c/xJm
2sXA91BmswB8eDGxMQr9j+RVT2mhkYawISPB/jGTFD7sfo+jU0M4Ywn9KYn1s2KJ
568a7GhERqFDSJw4S36d7mmJnAZH1z4mpHQSFYUeCESckZVKgUWYjSSH/yhL+xo1
NtCReKg6X5yfZQTeZ7YqRWCHtTWCs2iqJtDNpuus06HbH1fsQPExUHomo4yLDma9
yc8SNSaRq2ONnpwCCNlnpL9EsM2aqBa+DiGCdjT39RGOEMwVs1xAQUfWDauHfZq/
5nQ0PLWAGu1TaNDa4V0XRSJ9gLsi9GT8yNpq6IJAgQ40WUaz/y42ubgJUOwNkjde
0jaxlH+s5CHgNCMF8pzhcJ0sDLbRpxq3RMGX6SLhB5SXPSBaGnyvAqYF97c7VIqF
iAbXTVobucdN6WtfUa1cJ9c20SI9JdooaRACdIJlU97xJ+10QOaXl2kT5uBTA1xS
2WeSwObN7hyt8w9nLNutD1/iBCnLjFmBP1zVOftCWi0nBWugU53epJUzQZPCCnoc
GXwztGDMdD70pxndymCuhPmGC0EypLoFgB+W+2vwtuUcvpWj/4eNzUWmh1s/iIQl
ZvGh0koQYuXe/UenMMMCwUeoyrsAiT22eIOwWQSwao23v8x95gwjIUdV64R7iPrm
Qfe4VRC/GFk/SpzfAtsfLwv4zB6pG4sLmdidwn04GIGcL/7Cq2KgiuOJawwTT3Hk
CkVi1T1wGZB69tj7G3+zY9avd46w0vD8KYq5yfowpzq/7tKZvPhnoVl5owjggHgC
CwAaCMTjwpPaZY4dyNy/Ebp4NTCB6lieldEhgu4OttwPRkGU831zJ4o3a8Nn/reJ
MaGIbtOUNUPUrRjnT1tJxntX8nwImPslh5JZvsr/M4xvXQXMz18HVCNyRM5WQmP7
XlaLKkCqFz9o4uknGq7wxWL8lSFpzv4/qUAEw7WRJeAirm6QbBB2ouF0uqEAd558
8lZO4oMVQW8DaCQCUkkUb84UysFPZuEuqmKi3OREG4EeuGv0+O28Hro8iScd740i
lJw9iriqvxoZmMfceKzUPPOJAq7m8zubreeHjsoO6AfAfY4b0jmsuQfu8e6EPwba
kOz3q5e46+rX2/JRBs13KAA8UaBoMW+mvZ87BNbTm78zPBIh5cCMpvCDMkz+6FzG
FU+V/23K+LzYyY0gVEULFotA/P1ChdH5JucHAuHLe0roNk7YWAKjw37veXFVpfyC
RrM2CW8NWlN0njWNyQ5EcB+lAo2sRPPd3X4SxEut8TXwGzhp8Kd/16PgaTNPcgtJ
2s9ThzSL66WriAhsytqdM+Vl7MchmkmNR6xZWLH1yrBK1/y4pgCxZgT6vLJHVnhu
J3ZYtlGO3lXzrJQYqvPOh7fyWS1LyVyM3vuQJNMNQyGg9Dn+YuIRbl/sXkbsLRyY
tWGGE1kyYu/cSDs1f2E7JM+Kz9Tos5SkpHJAup9ks19PwnTs1DbqC92UBPLU//61
1wV6nnYXrF4y6/FxNZeiDe2SYIiV2GL0ijyqUD8foY+dWEql895PjZyPYilFFzyI
VSVfrFiHKkhODxzUvcftwAn8AQE1PujgCZvC4D71eLEU6iV3/m2hryWPnpiGlvqP
OErIBmHRqWsZAS3Zwi2ErPDj0omCBgqEcAPYdva1DrxlO0kkJNX/78z4bdQeG9/3
qrxw0xQX+GQt/nWEmXC14IZQmLG4hyrcmti0XPPp1B99PXKwOApPcJZVeTN/k3zJ
yzlWplsjUwzP7OoaDfmWtNl3l+Qrj9T9su3dRNeUg7QBrZDHVgBtAni5F0fDYr0d
1sR6ZxSA7wgrPjRmOcqzLl9pXiJ3iKhfsUXp/8xXozpbWzPxNZwLc4rGooYxBmaX
izOSnIvaIEE2ECN/l05wJ66sC5hmmYJiLF/UfqRmDQFhvVMwE/QjL9ITIgt6RcUe
amscJrXBj2hZv0PwxOa79ERfXU4WWVDIeU+j5xmu3vU7OIR1ElCsY0UuLebkXYmj
LNwVpRTHJTEoMaQG+MXW7sjAIT7DBr/qlnEEJN9ibYCAF59FVKr530feAACMZZVq
y3pi2TZYYbRHkkGXcIqiIbslR7y5G+tTD5UCRAcCrHJ0AbT2FRQ0ZV9wGvU9ErLd
MLbcUkwNX/yZu4BBQmoBHICZSKzM3vWlDqKOszL4JmLb8wTjngqIkfN6xWKO3pH1
rSEIN1cCJ4OsgZCajf+Zqc7gG63fJQX2NJ6kfVZAUL3eQYIsWq0mtAH0iuKFRLMa
ItmrYZzb8Ta44UTQipsBqOPNdayhbkSnIo3YwME0OksyroILfqUHvk+rEBV+M4m2
s6Z5DJQYrVggtv/o2njxBPOcr9z6TRRoyrYRd7HIK6223ipxBTWZUSnxPvdoE+IF
Ruiz4sCFltqz8/kfIRg1XbL1bnNeDvy9Kf93u/cjUry7CNwJamj3Y+OsNwREVRFp
QHE9P+cNu9iDQcA7TXWYRnbaMw8i/MzST9V9K+Ktin9eyNqkvPbNC5CsbinpQt5u
k0qCMr3rmHwD9b+l3Co65cy51ymAl/gY9YO1z33NptR0hFzM4B3jIEPVOHgMfb3C
CTAceiq5dIOTmmIB2w8dO0ZD7H9DBuP3KkUiTsrEMrXyZs/UOwhRUgAEtODDI2L4
aybzd0uQvqnV9wvGHV/Tv9uayWxoZxEfharZPk3IzXJukPftF7xNOht4D6lwVw8j
ldFK9KYMTPrSLORHhLMJCxaf/zlMkNmTbsfAc/Z5DwOfxWl39rzC13FqU7t/Kz4w
oqDMjpcySAf85pQtUroRNZx1I2fxV9qEVJZlrvdpW28DRX38epQs9L4c+CefoseZ
5TUuyVwAuFHAsncTzJwQGf1khkrTmw4T8yrMupEQfnKJ3C5scAlR2zYy+OEdDMO6
bM4CzcVe4OgPxd+z1lSU4++Tg5J4klfS1LrtQQYBh1pDsZQGkshOvk32ZObRIVSU
pN43FiBRt8vm1lP/VYVcOyhlZBvRBix75L+eYB5Q/zy+otmA5X13aRzhnTXWhPjY
JFmMxjUQy5j4IdK8tQN6KbG7xmXnPocd+RorPqtMvE0b2ZnMnhzQ/BHT2UxDaMQq
hbFON81/j36AnTlxMXbzn1dRn0goA1Y0dvJxiSuBiJuKR9n2tBnOcILZhLGYqVFr
c5+oBvjn9VU0WmlImzr/LUquoRPdlvIh29wp4LPHOOGTdzVfHLHlmWeET6wMTcRw
EISSUMlqrbrbe7cVQbOyPzmkjjT6pTwKE5wQY+6DmDArKyGIKehgBiC0Tb+yw7/4
Btmn2IRMglpYzuBDxFVQSeu/ROuHs1kuc4Y9otsyjaGpn0TjF/ZgXX1Ah/DG27Aa
Aa7e5g2pMX0Ue00YEDtMZQ79TLw8GPocYpNv5GrPkfioZ08XTuV922Kz5UIegnrA
iJpdsoB5tBBxb5BLKe4HvkPNgJGM0Bu5Vsyb6kBXBiBWTKoefSmW1wynxdaiyxpR
e0NjO68dBsCopeIPrp1zf9Kq8oZloqqQ+fDCrQIKUxh9S5jzHUg+UL9yU9i5PrJU
+SwUmj7Vm+e6MtUG1wo8y4jlevFUMWbHxAw7zN1LKukXJyG0tjK0bMMml2uftQSb
x+ubqoerVAg8g7DDJP2VpCuX6pe27TkTl8IiYbunAu+kGp31UFkykoaGYPTj9P7g
YGBPtJ+fwRcdqZZhfAMgHtMXVNrL4e9Tb0zSNx2MgbBaSRgYPnVavjP7sybvZIxD
LJWDmBYFYKa1UgzbrfEvR5XcxD397UJwMu/VR5YVwLYr4t3JPMHdHvpFjr/7euY3
1fP92IjmP06wJbChjMQdlQknvaG7Vb1OCOtbcn696MBDuqEhUB4Jtlaqq/4K2r46
adpnLH1kv6sS+tPY6Ubt36TILq356+ySL7wCNihCcQ2bucm7akomi4r0aOSQWR2l
uZ3kZ7J2LekGqFxCboJ8wDCln1t6L4oq9p+UsK0+06fcEfTkATfym6/HnoX7IkRa
Ekf9ccJRBCQXoIDJD7JcXBK/qPubJGcNl0RzwOQc6mFEWYXdPLuEy7D5+QDKD32o
xCwGGe0bcC2u/lhQEXGYLPSFci9xjeG1O70QVo4475KPIMTexM8wQQjFnm569nI3
jisWvNo+N2gf1k4S9m8PuqU29BfiK7o9AnUComsaqarGvz0lj6IAxC9ergtcNq3m
qJVB8SOLYH4JxbiLbXuKzzJnXG/+tWwrlix1UJvkd8BPfUbiJsJmoo3MiAlbkl2s
P2nj8u+6NcAYwf+NLzsLVI5EbCfOmNbti6kz0mGlHUtCAFgcwf0LYmLEJQ4rTZpd
iVFPASVxxmHC3XwJ8sKQdjWIjVE9hC4nPTuOKIhAztXfNEM/W8QLkWaHPtDfPMXI
ofBaA0iEcMtoXdrqOk0lP+bRP9KPtXJJUxc5wHXK7HooHz0LYUhzqW4l5/ZtNiVS
SQk7eYWa+v6hWbpbm1+if5b9ZZA32HuQgvJoBv0flghGblNWYhBbNtQFdBvwnWcT
i0/nDknx6G5M5ERrnxptdorN+KCYjD0o44xco+WIyNQTcd8FqJ0AYZrIL89cMrLa
JlIy7zq786bs6tbq+zC3D7Ir9KnyZuj9yTkrG/0HaOZH858HAmr6ZbSXL15kzuR+
rg05X7EUVptshyXVT7DxpDOUoPmfZ4b5szyX9PFwIpRRf/b6RZlrPim0HrGZrqo1
aZur47PGV/2nX4CSuzzVIcnJ2j2HOKFuHxxrYK3BQwPaOguMQFZS6YcWLWGbJ7Yk
VVXyOWeb9wmup1btgtfX5NdkYYvr3PjsjrGLBQURAuQ1lS8pYTub1tjHlnpN44Fy
p4P5AHseyT91QkAAqJx41zkG6/Tcu5eTxX6NjSmFIr92vltUAoKOH6f5If0aBZjF
gTXm4xAoHAyVxmLbLS0Mj4mZmzRz/3/KnWfCKDNbFsdC3fCGz81x+6x3jacglCHn
qOKtpkOmfKEdSRAyvMBLXAlDG8R/CjYLbXZhpvc1N4uSgDJLSF5sJQcThc4fRU2u
TYPPhSHLLLL8QSHnbyY1hji6ELeC2jEy0UiFlIOTgMO5rPz0fABSNUdgprchplOu
j5OxCLkYf5lCdijhl75rxbjLpOLtMWgmLGU3J0EwaxUZfUIICEsYkg378Ckp4ueK
OMd2sOEZfiTAw7TJ5tp9LE8PcVSNiVHr/I7pSK/huzpkremwKLo5FtkaQxw4b5T3
6qPnv5hjowgpxQk8AwxUchX6h3OlNdi0GCd1NbJU/dGD1AOITlxJLTG1+RKQy22R
3uR7Jdt29K30NlT9FyRiJAtrRAKl8WUCrUeens4npnp6YdTKTvHITn5FKvZLr5O3
9Tzl3pFTbuwrNLpZJD/bLn52ugPZiQC2tcktlL/wXD4FYMEAimSTCYEn8pcgYBKT
M3NwQWofQECWUbrTQMunCW9S77GSC5diMSAtsew5qbcr7EN+BBa4H7C5+Yd4+fxO
JOyFIZYEMlVkMHdEEaSuMlx8+BVsX0Mo4l+bS5UD/SIXLEBjf/OWy7Qte/pcbdq5
/+D4hRPUGYRjpYrR3hrZaJuVtUC9tTxpFfo3DHFtb3HS08F/NT1XViNF3gJ8kIis
Aya9J3+NaThvLy0znW53UB7406CsvosGgR+7SngPxvKpMu4wklD5sGlCePTvz/b2
wniWct5/ro6YlGnsoJZUVjxZ0W1WoIETFwA8YaTa/0tPkS6QqvL/GXlAD61G/Y7p
96MN+2X2AG/6UoTPCHm7YdF1pDwddFi1kU2blFhtADsc7BldPihl/2wfowrk6K1h
UqSfwfZPAGR0YI7oO/ZoZGQNqQAfVLirINGOLvAG8DaY7OvbcMi8SL3k+64i1Bny
DbS3yTaTzJcJlp6cbX6z9ORaVuuclgOjeb/gZiYI91NzdfStG6ysvbRpjXSziLeL
IM/AaEvwB2YUxrBFLZiJWgYYdmDfuFPUZTdk1MnakS/Iexb8wMKVGgjGJgJJIQEZ
O/wTp1fDEk7mGbUfKvzQyh+aV3XW6iTA3Seyq4jtdwTBPWl6ahob4ucXLk2x5xme
JywcAXvSzeaY+nwFhGZyL2vPVwA0+dYtw1ap2J7ATgE8DQnjmRzpj++1T1YodiIG
nUYtx/rfFQQ5xGwz9Oggczjw97lL22Mg3RIAVUuUTtt0gKFt0vlhMVXerffEDBJU
OuxC01uoV/+/C69hTjFSUxPZGEkhZXBZpPipm5/yVzpRZNCWgxZiAkGuqlWYlSe6
ARm9E3/shU5/KQilpasugyU2KWHtw4FMLRzWk8JaPwO5DmCN+UWF6uPz9hIUhUmt
I0DKC0jJEGMKGZCtDsBrCUvhuvEu0TyYTEgil1t6WfMwM10nGtjRnokvK9fpg+il
yNpkDH2fCK4xzBEyN3Cx6FHnDTxzNKeNhZc1T/m9TUOf7ntPMdpYj8fRM1n2IoAB
QI7Xv1k3USyO+b6L25cVqSPpgxQwXfwhWVSeyDAf4tf23iwan1fLKbJ1gm3lmed2
GiScjKB5p4pdxtmM+xOYiWhZSmzyv6+QFO4vrpNJQrGUD/+FiQ8HANA27bFXeeaE
MkFft8Ykteiqe9gtIszpG3veLcA/Ow8m+W9RpclI8d1zPb+wnZpdm5bInMjFy3KZ
SyNnqmkvyNPKk4gPRL+weT3BboL0CDQNJtjrCjAcxodeJOhtyFScuxe98d9A9IBC
9OWgk8uK8i4YTRDFv62NRF2YVC+pSVQqj9hxa+F0QR8wdVah01sUxM2U3DGsQQBt
SxMxY/Wp/z0+tMSkQ+f3SNbdCCzn0NONB6bPlXyRa3w+d/wjPpBSFwdiSmH/fVJB
sw5Upmz8lg6M82sNiGYmI/12FZeGN/4aPoj9BzswSe2y+NRex7sDCNLya2WRkZzH
VXj/E4H4R6SlVOguHiI/urWvsPgaIjF0coYzOM/gjexfGGaJwDYV46zbJ8XtLHnM
Ypbp7KFQikPfEx6FwS9G7l2vkXot4wC5Orr/CbfbWjXLUbqo/LZqkeR0N30+mhMo
d1wS80Z24qWBoSJ1/qgc6OCinMNG/0HsU37h5/SCWu6utLgv9EHuBGCndTFOfeIb
nRi2Yb4ZIbXAX0QgKGCqVOzLJY3iM0ZF/v/4Sf7bv2Bhmf7cTeGHx4Lvq5klDFrx
z+QWaIlth7iY/pXb1b1pine2GJTKcmaLV037MdFJou+yHwaXHKzrJbm2DCJoDk/0
SaV+NrtixPPKkVuzeY0ASVe7v+KzFq1VwE9vdaMzjv2ts0du+/vtLFmTI/aoP2Sq
AV1/sE8aTutobFXDIk0EXXwYL/iF6NAiXMUgwOLh0LddVgo6iiin6d2WE1jq94E3
9FoctWfXY9UpCMwiMtCtGBjMiSe+1AwGqgAXhqfVlcg+5NFQJWAOlI38FlDruzzs
s7vbHSHmjUP5K8dAWQrKcpeNS7JZbBDQcvHPTBpTCkz2zq40qnkD3PewTd+9AFCI
Tpb6Y8afJRLaLLGqSJ9hT3Mx7JAJ5uLS2jRE8pUijMuM+I9VYU5eHQ+yBpuJwDZV
D5tQpiM8D54WhC7W7q/nyrSGOsCn6IMTHT22wLjxoYTZp1sIsuhLx863uGfHG27/
zuTTag5/4W/RbNjHOK/uyfHbv7sZ7RhYABmOHKCV4hBfGfH6KsHchlCDCws1e4In
ZeQCRKlKB69qKYdZLCoB8agYNUgMozPB9jI2I2Jbxi+Srky3x99R2JDElOvTbNWc
h+tQNhmxZAXcN0NT8cff/kw56LdRnH5xK60h09uxwKuFMStn7WO3jE9PvuH3zit+
+LEUyrBpc8RU+fzwPZyFbjSciz3Z092sgnXNYYZanfUNDgZ6AvhevQXL9Bnby53h
fcjagWuJBt6/6bGmUXLTrUg3SGEH9VbZD0Ra/4ZE8WuSJ0DkcqSDGpzjeBy4UWBG
gNOkpVaiBh2TzIsSULyGMQzoePRnsPd9h3WoOeNv6DUNrgFBKbGJ1iD5S+W3OFSq
VH+ro7KHXaMHVgE3yuT8rd18fJAeORr18H7d+wsY5ehsM5vWfiCXhdJg5pCWHGaD
oLgC2uoZEUqSI6IFTFHbHo4cO2oornaZxIQ9RJNuQmmuQWbPDW2tGwFUBz1q3ywO
I6Y2IalrHx0/iP0I6jOs/OKXDq+HVm6m1HoKSeOp21mEweNgHpicyZtj+Bi8pqNS
ed6pSZUeMt8pYEyHe2CrNkFkEF+vJJhY1YSFq/dQ10qwykfuzhFHgLPIPgs9DbsE
R6sjqxkFtXTySrGMMg0DgRAenT2UF0ZPc9YQUMQfvhOIJgf48aVcNkkzuj3wn/UH
W0HTS1RTJw/9K3z4xYkEhn2q3qVjmMUoZql14jUN5E2Satpj+fRsoky61jOnPWIv
+q8l7c90rza2nAa/kcFnb2qpYGHqaM85gVACyMmmgYIKd3lxigZZRkKtDpOBJiDl
5hSnStxnASI4cqrT1sGeNT94vHP6LBIbiFJ3bdKnCF90U/Rhgvd4Qaakg7I3dJIh
5bc0jqrSsKPMLZuPTGnHwZ1EoHT34+OK+CVnGrRR/J7KZuhEpcnAbQ9j127r4T6X
2wItJm0adD2vvi18wIxqqcTjaGFXhT5f+Yp1Or0n7dWjWAqerEX7XLryHqaSGAFG
T5177ColmvwKSPmR0N5qaF5E8l0tVFfpDwi+P+LH5AWFMEHG5WV3rl3vTX+n79+E
izaTp1+VGztWv2FsXe+cDat200XmrLzLJstyxdzThwpMpyFZPlEkRv/rVQYHhpFV
bjHS6kbFVLSNJtotWfFlXTVHnXmjpuBTBjrvOABGmJIXxvBd/b844dpI184oiCOA
hfJs2XQwVQVcviKbgm+7uXC2nZXohGNMKAXxxBs2hlThbIeUfkQCZu25bwZnzm2G
F34SjhIeXN+x0+oDe7ATD0GkcZkl+5rHfWFHMetjeUij58XahF5NFbrxni0rx6yy
M9ModUGSiL1W/Hk5I5k5rD6K7C58BMbEO3iQunJi785t0mEm30aOIUqr1jK7dLZs
7T8rv8eCXTy4Xh/CGSD0jAaQhwHhDf7QOFav05JBR8pN88Ab8ev23cKkJ7D7pkF8
jvehtyYB087kSIE6mkT6QrnIGDoccIj4yLKMuN80nd9+C3nbRmjQzLhagFGxp3fq
QXz6fSCrtHRgwR6wTsyO6s5m4TiVBelQf1SmCmrmw9w3OCJq5FPudrpFp1rW6Z94
3/RbBKzQypy4frRL4oXEnbIGRW76Uxet7b3T+W0nYeB6pW6RP3IX910yle8vp45K
g3w2SOnWBzGtVKkA+2m0TSrmo8gecOdOBv8IyDAWlw+iZaq+7ZkoSOT99HSB28Sy
8GYWqXxk2lUDPMwPK2irdN3dnUYNx2Vhs+hJZKz0xhh7hDlH/py+qOXjNTpDM6IR
hqR1COGs4IM9by4N1mSGwjxEjhdGUjOqQzvhwP2mS1OOayRC37u64VXA7EjAUU0S
CGknjwIyAqvGiS7NyeayjcHhPJrJwFql1lI9mKoDPgLkxuPIA164QLoHit2drmqm
R1Q6jdb0t8dmVB6WJTUXTPeBSVGc4rCZdFrkZgWQIpOX+Tp7tuMPTAPabwM9cT69
YcwxHXCmfFEkA5fekQWELBe/YBa+W+qB1nSIV+XyWZwiq/mn0zkszzfXm1Io54gP
cl3HA2E1Wi/oGUr02gTVh5AbYqSv7G9XV/V0niwTuoh+ptkgwIBcDO9i4grO5u4z
EELUkSxw/sDX+bSE7UXjwoQ/LlPFc7L8nEiFeEEccdWcSiKz45WNYw842tUPOySG
aTLFu8wXUC9rz97kma5f7ztJGoLIjwgb7wARdTw4wfk4jwZ6PKPGYmriuUhT7iZm
x5zn72vCXN6YpaO9qvMGaAuoHRyHsh0Z2eG9VWOUn0ndtuIzpAJdKoqsZKWx222U
RK/aNcPjWOfy27urmSVlQoP36zqziSke00k+QYfkqPOpc9EN6K7uk7hIhDfUu+Hq
6d9KWymgIwYQIZYucw1rw9VDLq51OWvb6NICOUtC4f8x8o2uiz6RPHrokmLTb8/z
fIJQJbb+MYZ+mp7ta/CfddhrpWpyDePVMRjjIx83rUo9uoptIDhPSkcSamlGo8Jg
nUQKGImqD0JAx/VEn40qenc5+gSc/X2oG/81iwwjekq241+P2oQUDBjHJcKl2x88
kBpIsuTRwAJPznPYzto+XjrmkvqGZdK/27GfkZqgtKyZx1Sg8zFX5hdV+GaWixJ4
je9aFh2xOlRS4HjFizoEfxIpO7tb5dxGi82wcffW6DVvoc9S5xqkAeHN2k8elIxi
6UKAbNAtcGMfCqJFxxsRv3Kbmm2lhJdDybefK8IxXYHXzxU52nRzJfMH0iBjWxnu
kr3kkaSgW0oTt3BZqSHC5P7P3Wc929CYTvCCdGfCTrkxj1fPMUhtChmCnIpAhWlK
Sj3hKcwbN+Vj0H2lWYHMr6fKblOnPfrk3Dnx6wMoOFNfLkTYexU2PX5ruDe9CGGY
zj/Bs0MwyKTYpTVTnJLSD/jVcPkmmY/NLmP3PRHZBiHGoqGM2OaCAZ4PNYYZKnYo
fGU35iiqauMRPJ2nn854UwN9Nbt2o0wKf0LPf7KcvF6N9BnJGpfsFRN/uoM5V0Xd
dopXrPyP+wP8Uxtlu8b8WKD+xcjs8o6XKi8P9Hdnng7LmRcUNsUejq+NL4KYlvV3
69G1zaSayMom4t2Q8E0vrRjNxT2pixoYDfix+utwhhK9tkCLjASg+cJr2TPec5Jf
xGoHn9O/fxnHyZCTJi2JpyuByJoISmHtNF46l5JpMenMzOi/WqGQjXHRTrC5OUQa
HKiPUntivjx/SEfwTznWrk7tQVD64lLLU53xXX546PpDkSIuHCO+/HOFL3zNRsLe
dwumMfJfaFG+b54Yj9Lsnzj2lRKn74an9AF3Hj396eEY0FY8Lx2gAqD+XEJGBOhO
gNWly0e5laZQLPWa2VZizQMUU/bj/34xL3rHhwqz2/93xDvvWf580m1p3jiblqXQ
ufEj6b9r5DNmscuIPsGGOYGU6pI3i+EPacygjb9AE9OmkCM6ef6zLHH+di1idPUL
aM7i48y16+XiTDAtKqPniAnZMGxtxfcPD/r6fvpmLKRQ4xSWI8nKYHkuA8i1ik2d
bq8Wt9RvaWEtt/twUOtpb5+YVp+R25pLdSYxpCJK5e1fexB05PxZTvULtJ2Ua6x6
siWP/JQMcedUrTZty3u4H5piVMfjpqcs5YTIvtP5B3fLdg4fRqMN4aC/7gelFcC3
Fuf6PFZ09/ygNfIg91Hm4cNKYDY1XJv4YzmrAFlUlt94P2O7+OCNtU+5jvK6MVBx
9mYIPc0vwRX69uDWTWQAqppG5P4zLBgXOZWMvSd79q+LyLqsSagQC0zajwTG+G6f
bsSmixBeJMLDZHqSwDaJDU2QYIDMfZVyVwQoG/HiwcrmPEYB60PAPPDHKeVOPeIc
hxaO7DJJg9d6OrR86z6ObL5a1b/6fLWUgIn/JrYOfS6EVjH1Ep3ZRK0zG4GWmw09
zaxIp/vwYknmHRgZ4UX9Td/Qe318+dMp2DVW8qylFj2xsm00Vo0x19LbM57iBFWd
+tC2hh36y4MhC/FmOvKdwOvcx+UB1sySU1++/Y6DLwDBaHMkuujuC/UP+R8NNHib
SOhBO4fM0qsR3veHY/7OZp827pHOKNnCu4lNGsq10DXNm3ZTYa7gSFodXPmgyCkC
iNu71w6gw5SC+vZ5w2Whv1dTUnVinQViecy62T5nWkrCZQUveXnRZ8l7YSOjf/Rv
qZrMG5ww3pObsc1XeXnIGzc3cQ9XlGtBLCRNU2ZW2DO7ojTi78Guo4Nz94CfMepH
WiE6/1X9mk320XBLoSfDHJRzwKWv7cxv9Ev+Q/qpg1TYfSPd7vMna7Me2Gte/J7S
PZfHkM6f6jgHXyXy/ui4hzj3FI+dxQwMeQ7lzVbRkzT1px13Qtd24bKnhclmMPij
wLCFmuEvpYdY3PiBXwTHiy8sR4wF1QiockbJA2EHXdQ36koSgj5o3eAoiN0u6po0
qvDRRASjml+TWn+qMb4kpez1xb8s7d/Hm0ld7STema/V9vwSPaaAN55D5giZR559
cnra/9umj6O4RtSjifmP4jzdp3/YJFJfddoeOvwn7fEety2Y9UjXCAIFFv3VleCf
sRkRNLdn9y5P2sX6yt8iO5xeHvAD1p9DFU7JlY1V1Dpd6f6F8VLbmF7h4l5h+d2i
LM0XaCe2B6JU+bWNAsVMUt16AZQBTxY6S/dp/DzC3xu4cxepyC+uxGfqBkv7ZrIQ
6y1FuewNeVTmSeWkxMLjwVJbEpB1TANt0LaLAzL1CTYFL7w3g9uulIU/r4l23XlK
zeyAd2XL/OSaFDqfK3mcIbqfzXjxATVMipn5CiqREbwc3n+SQCt/nm0km0DnDt57
YCPsDZRgbHkEGEnF9mq9eo3QjXvzQypfV5xGbELhK5ayIDZXiOK9+gKaXGSJwfi5
h4qGngJVTJo0Nf5+w7KJgC0JP0A4YFWiJOlfwfB/Qq6YgOCiUppF0PTAZLAiq9Pj
KjMM+bD1qO1aJbmH5PGT8KjE36j4Od2Od7eqk7rLpI5udCULaHoUdYSFo5SZZffq
rDUK4TmEp3KLNvrpIlFgyWcysFKVL2G3F4LAV9xmcU9X3Ja7Sh/SX/aWtDFFBmIF
fP7eyKLwiCQkcHvWqrNja8u/ietC65ARfAbHYsDc5HCEleWqK6EjZMB+fACYP357
xJ9LAl1PzmQuECG+QFEWuax0HpWghHOLJf5VSLsTMnZoZ7K4qxVR6L127ToTRLsQ
KAPJJrZyCDKZ+1wH1P1fyO/aDWmqrUF2T9fuOyhaWK8mG+boFaJPmVB5OGR/zWYw
8DhzMBVFr0ujLe6GoTGn1pFzP1EdWuCM0109fRjiYQjuiH46AFMWpgYqtgOFHBUC
MiQZcoSySoQyN+66I4LSkOH8iRF3zd3tjNx4OzZIxuNHvlPdtlxGx9M0sgiZJ0A6
WCiMOvUbF82WGnSQLLAte35IzUqJqDiJNsE4zdhcyKXyoLQTm0kH5EEjkjFAosPL
ri5ARmG4OBlAoTqEjeTOWko6eaK3xozXMJRfJ2r868m2LiWcJ7IbwGX4Mc2JT7sz
zQdRaDl6g6UzZc/tp5/taty2D/QfO+4OuotXnanurmxeKXOP8747epljWNaahFrO
b44Yv8YC4Sjar7OPxha3EBPhdmrw16JcOLwhT75pTZr+0RiHioMNXqXS2xnt+0xc
nHl8M1fszoWVC+TsI86QxoFdK9tGzBNHgods6MZv3VIHJjjt5Jcj2l2E3bn2GH/Q
tYxl6kpgngBtXqLzGPQC9Hf1vY8ORRTqrkSZpe3Fd3ixVim5bb8fP/tSpUkHzxte
XdKQ3LopT9pEkGaIRsClzv2zWpG5LhCppZfDPj4jHAoxOy8+jWu1oWvylT6E9Yfv
sG7UmcHBWND1blyrXmjDjR9jsF+I4lsNm0MNYPRpVhcGdS5HFZ4XBrkFS/j0eRUC
eQKWR8p5Y8Kq59VT5azcCcs6JOJs9A+L9UiIn/880QkJvS1/GNA+CZJADTh4mfat
c7PejwzEyUjMexf40nBp8V0HAQuzef9qwJzngCT+f10yMiEOqi+UwkjNpbE5F3CL
1ezHP45gXSPw+jmwv2ji4XcKQqeWwxUFcjUuG14zFB+/5yu8/ma0EiUOX2iT9zq/
g0NGCEZQX/OUgAE7/iBQr5FWZxxBTxYZEOA1+QC8AdCent1sHks8L4vAdAJaqaqw
K2+q03HpT+ocZbdBhmmjHfUPRXdA6quG93QwscufY/5RgUoReTwYzf9hOO/AIlkR
zJemaQtiEjnmG1ctHl1HkcXUCqrTkUCVxMxGQFwsEsSLm2t0KUlDLeOHt8YG5IRM
JzYJsNUfxKrFVFZEBej0EZDkV7+Dut79/SgYpbDO7KtiC84M7OpVlZJ8qymOzguK
QzhJN0j6aG9xcBRhAsrBxVGObhrXovCUrZAV7hkK73FvgpfkZe4YKy/8/Fo5cXU1
leE5Wy+kwxmnxQMm3TnyokGZOSFIikaYj1QT0B+tpZN1EErnA0DlMKDkoxpD2GSd
10BdUREiqLfs0t3hXi+9JKetzch1cRxQZN8WEYhKiS4ZIRiptgcCKwrukuwoG5U7
/e1oXH95kxqLVmNmm2E9TmUN2w1w6/5dOUExpnY9eArVsWNKw0QoX2SgSM2T5y1X
5JxQqU0G0V7v9bj//sKgysSHipnTiNerOzcgZ0d4n7punmDF6fi0J76yGWM39DmM
CHwuo1aJCppne3JzzWnThoDiT5vwiqj8P4FotVHW6fEMiwgUOgOkqTJJwcoGKqwz
zZX19yT/KwToENI4vvmGhf955JpH80+j5kk++h/yoqI595jkR0Vpxonkji6cAMuj
wg4yF+AC3FaT7+AySvVtHlvDW0xsw5b+O0/+MxLPBAgxfj7oAZX9Qj1WJcKjZUY+
V1+s5rTOS1JDesl0tC6NClmMCqG6Seq7kvqcGbnv5jBAn15dUR9NhSKcAdNX1IHG
6xjBCzLcMgEzlQUeiDyLhV/PFJhjplS9zuH77nZZ1N4BuLoAZPLfcP0gN4oUrWXO
2zBuluXk1YM8Ujx9saj1QVsnqgwWlq7Jf+ZHAlSGctbG7RYqUrvqqtrLWo4txCmJ
BzEHLX2eht4Ii7C9dtABeXjam2G/WqaRdfTe/XzyJD78pgS/6n71k+GK+vISvpEk
GCXL4GcvVwXa4SfHB/+UUYUfJabHEq9ZUKKm0RvOv7njpZC2mlDYGFmc3fJFnCRt
aunF2W7UL5tcLq230sXIINevkeWmKG8faaRYXTTN401gTv7KfChimhkA+lXFlswq
lLgGiRHv2tQCWuuVydGvsQzuidvtfibBmeFa9Wv35aBr+PXrUWM0iONlHwNwCDrM
SkqjErYxkYoBnlv+dwOzQlbVUWWKxbVcXGPzeXicU/Tm/gxBuZ8UNmYooJqG/TYF
wJ0aURkXNPMm/M/nUtoJMa+j0wLn9vxAtFnt0Fh8wZ40wV91xOuMwiM/L0fOSYrg
ws9q0H/csWrqCE7oPL3jGsIPoeFmfZEQyDzJDmFemCP7Zkhj22tMJ8x+bJ2wTklz
IsDFQkeA65WPN+uBAtxtDtATZlPLaCXwn+VKcN42upMqSLeea6rQ0M/Llb/6YGFX
mWp0SaGQF+nfQlOaV/f6ZzRZVelOtC6s7PBr1BNJQx3W/4f6dG9QiHIJad7fEWZr
x44FzoNJLAtydFd9QngmNZTV/yCsquqGI89nhYjqAwl3L5Xqk12FeMrBE5RKWTUq
ZIAqa8B/bafA9nY8waRYdwlKUVlCjUU5Lc44j/4Kmq6bjO9xlZeX82JyJANkG5hM
Hk3NoMKrGQY10O6v+pGGtGfkF70sWZZwoVj89ZuNmUeZBddXDu8lRjuC0aqL122g
t411SejS7rWI/Yry1P1lvg9QLTcSkXAiX5xS1B+NKL/FwsiCKySU5aoGFuhGmchL
WkFv/lGXbc/L0gNh1aasY1QNKlGc01WJsFDZx8tHmvKwF/BDYmsjzLWQs4fgNoeP
LX5tyot+wU7LZlbpSGUjD4e39M0o23Ps/f7Qz4mwFfLx05vh9kxfjoXDilosJjwO
eadQXz844AjFtd/SCZsy0yEUlUsOZiKHVw+Gd6UiVxSRUyp9uxQBMndE4bfTM8J5
TpkucWVzUtGJp3UOlJ67eGSIksnoqwnQM7zrPpTHldDfT7qsVkEN2m287PKYRftk
0Pc6Bdj9u5LUzFYkOSyl3bsdO7xZJFd/uK9262apXsaXd05Ts4oNXjYKz5knuNai
q7QED9rds8wuDzG4cm3MfM+v+mhpwfzWhW5GJzhNb65GR/g4eQrn9b2X7IVlThPs
7WZzyfBuQyvdzyPELjSUNoNvbQ4yAPo7DYUenwJMw842fJwojTlx6Xa3Gy+HldCa
MK+LcSlsy3/+AnuLE/fHQhFasaCmUwjIOz+g5sAvYNCLqQ3hwFXHg3xhoubjTPYg
ij2iAlGRgh/rr7KHFAzOfEJULsOTt+9FXCKOFfRK1PHM6mXg+T8obTwNu+seio+L
c2VPkDy2wq5D40eJ1JFqsizdx+lqK5kDDkaEtAudUEZ4MkXca7AVSLWvEb60Vhjt
cxDJ+0xfj2oEinUOvvDFApNyjCFqabHiIebIotL0nilSRH789E9EmfsVMM3riMoq
SsTPCo1l3lR12tugPa5OBO7ibewtaG4ArquFLQ3U7+MAe6Hdi+vXN+pTDQTye7PN
ZBy9E5WyYvxCyaj/RHvQfWAvxg66wN9nB1uv6qrgzOPkB/z9SdYPDMfbaEaxk1w/
zrz5YjF7OVdbhnh3MfoA/w/IibmpRlvp/4t7Lon1YxH1MHDoumrQa+hRZJVJUr+6
Yp2WCQ8OaES2hTwJKrauPd6wOLtZf7LR9sGKxKeDaRmbej+VL8KCdo45vGgE3SN4
IKKlycupme53oKd34T3HGpb9/qEoenC+SOsray+U/kkOFU2KPcwxxlNfdrWCYoWn
b+01PxJKa0+uaSXD5EsxuzcESb5PeuH8UyZdPLWyCvGXydBojixGd+PbOIprLJ5G
By2tiKcfzqQgDkOKmqYJJkgpWIOroRAZtM2UxXi6hIKzH+V17LNwV5dAFq1Aguw9
TldHl66et1IkkLBXDsMuXmN5SHnOjFi+QhRcLZ2nqDA4YVBAoqM2SSC0bymQmIlv
pGCCwJtpu/igXdAPa+u8eXdErEJO4tRL6MF7mP3c8qURD0FngRiqOnbGrDorYabX
S59AhvtIyBU2A1Pwwa215y4iClX/5mmVKjSY4dWQ0JAsZseksCm6jEWaxMcd6NfP
uUubsja07t0595fDEvC5opbj08qETVXxDyXMEh8RM2ExBj/UhxfVOzCEeZmW4P4P
CC9xsKajIcQr4hXQHwSzABP2UIcKi+aIhnkmYS9QJffLbJlqto4+v+cX23ybaDUH
0Gp9RQr5udP2Zrw+7Ya3eFb0KjXZW3SmlaBwEwrNoAZEtCeECJokecmUJYFJlj5D
mR5VJc+Y44rFBVTYF7RSgNnV2gU81liHluSuYsv+XUtjCL7tlwsEEmx5NXk7NYCK
YDLrbqKGr2CgZ360B4QWwqi6uKFiFpVJZKqagY9kz4cWjPPx2itqNA4MNpDEivpW
Mv0A8U4jr020kz3lfEjIc0BXZ3GOtpIbbWJzmpFQuZwBWX1JTs/8YKg1auaFCX5X
J54rx258GrGhz3jbPNQeNc6TQjRohONaWg9/3PakPkuFaGm7Td4J815FRVjZeHzz
zp4/RQqhSmRV2wNwn+eC+vxDXbTKKpBc7yieLWRLyQKvVUtpyytvJ9pPw8CvogeY
6giFd+J/1N7CrpA64Hb1RHp3AGTH739JyxRhbz1q0y8OLme5ov9R2ZnmZWkxSWy0
aWsoq5DcY82AMt6zKRfJAuBuInWLzGZHDmWdqLxxwPeJVfpTGzuflf85mosBCqPA
6bh2GaQX5iST3iEFKcvqJOnjXZz9S7oEZ94mR2OdaCikwYd2QFRgi0IEPGTdJ3fr
yC48Fj+9pf0X8W455t6cdaqw22isZX3ImF8zPlHuGNvXxstbWq7po/BRQNA3wqno
zfi/OBMtZYrS1vY9+2DQ7bkG0FQz4S8sfqUd3M9RgPYEEEij6fSyXBKyj4qtNEPC
SLvh58reJub2OY4R9UQZQ/HpeGCQ2b9WcFvIL/iNq4Y6MbIMuL7Fw+u3rK0z40Gx
KwoXMGogNV/kExRXfiZiKcif2zKwLpmH4rH7DAj1YZeyOnhD3t9f14Uq4dEPwOuw
WfXY67HafH6pRDdDABqYF4i2iktpez400qQ9lvqgnC5QV87hntHLBvRtFvNhpZVa
wJVSMtFWgCyVnqOWJ17fy77RqPW7eCBTifrVIM6PSJSWidf80PaTBMR7g6n9kmIR
+XPoBTo/nyj4pyxUsiJvFeZt7JmItuznNvNSiFGcmsKSD1GfSFEaqTNT4yUPCmaF
7tH92MmgtXoT7tWWYBI60Nva00kRKeQ9atNGMc/h9o0w0Xl6GZd1/DjWhP2neSoe
Q5ytzf4pb0ImuIalwtGP3y5YgBWmESvkGIIkdZTAwtNZChYXtDwOpaPo7RupKmdh
bu2pCdjVMvgU2ECn77enkiEreLN4CSRlCmbo5EFafCjLosrn7hpNksaEHRBYPVAE
esNdl63FZtYOjYtc47RMS+rfXpWmRngrqChoLOlzSMyUo6kYtBPICZzfzQdJmZhs
SPUA+9bGKSCunoNf/kNc2nEcG9Tq6ApOM9RZGqSwtJdkD6TL+tw9uRkvK1yMfmfm
Kp3yD6AYN23bjbO3Wjm37ybr1j/D7vme8IOVuK61i6ltziWXyq1d5+BdR1coRLxD
zQHrhGbpSTdxEmFS0Lg5xFPpyHc7XDq7gyI7hO/133Ux09T/7f0N37SSKwt4WYvc
exlM4BFWKVH4wuABSY2rTGR7XGG8/qvTmPApyuymQxkxW0hD9f2DSRqYDv7qVS/T
HwnPknzhaSMy/PEj0WUVztC6ZxUxG6UlOX2qWM/uFfVac8rVSluAU65r7TZPijPI
Mo6naK/wTsBhGuXgcTAC/WOCDT9d4tohsYsjzr4bkfH2bGPgdRLpLPAQ1+un+Lf5
MXxNTY6XH5J6HowlQJb3mMYwH3GAEIX3Qj0yg/AtzcHIQgQIwrgwIyV+eVi1+5UP
/sLcDNxWLVfS8TjpO3Mpc8qSDdoGZDKf9OBgpB0GfTuPWsYley9dXhwQ8FavUmrF
82FQrhxz48DMUiTa7+awlq/VKRGLGcppA2bN9o6SccBseUw+gqe7rClVNQ0w+6CY
Hk/TbhJfozBsbYaDhCJLx6ItTLdepDAGRw5OtWsL+9YFHyYd7MvRwhEA//6E9LqQ
RGv8TT3/2i9JXLrVEUjkKNNntMA1T8/3yrKviKEITfOT2KxC5uH3RUwLxqFWtKja
FXzzjZcjuFxcQLBKiEoXDcNAhfdiTlu/o0aLEu3zkSOaxo29z1DcGp5+IVHLuX7x
y1K5RGiafEmmx2pS0jN0a694xone2dHQfg0R78GNb+zudo6BRm52+FS0PS/jFbxj
CnZHGJFy7mYTflwtWulaTL9uoj/FnlAnnsNjVxv28/0v+nP5F1JANrlOLSmO/lBF
iKdkFgPXPvx8wtHHpLZ2tBN/yxBFeWmaqJPXLA6nUnyTe6grEkxNQ9gRF7bg3P/f
YBpMY7xOVcfcbvukOo3xyM5l37wAc2UULIUbGKlXTfXgOb8xaq/rxZdbdgu5tj6y
U70t5YnkQstl5Im2bAgTA/CKa9GJAonwVjG7ljpzJTBC1DzAzlWyD24fhI46dMuj
UN/+/XGM8BEwPW9gmd9gOkdoS5AulQSZdwXRcgrl7Hf2U0LEWgtcZQ0loao1gKsX
y+k2mFPdbR6hnqVhmHsCxAvVPqN9/shiiqJBOjC7Uwy49YUloc1bvAN97EUnLy4n
Dde1sy6wzKq9JoR99CSmCghzNKLesZSRcXT5H7unosziYfUsWtOjA1ndt2UScowL
E7YK6SFCLruPKt0aFp/P5CLZ7hklGYaHLAugbUZDGjL/dE/ehTb+31y8hevTWirb
oS0jGKYwVgwyfdstmPgdNkx7LnYsHWegJ9D8UdVhvBQbhwBkcHD/l/i1Hpli4r5V
GVKHmBUq/IC9QWe1WVDqh5pFOeXXA0hRzrpcvUeRkE+QOYmwj7f9Mbzm2iRFb6n6
tQxvY9cIUgVuqSsqBmF0au9/Tsr3xb0uhxOCLfX9rtUZyViKGvz28KtXFJhMFzaL
he9K0YErZKgZWKT0Rx0Bxs/IuuQYJ3SZRJX6uj6S9nfiVFQi0vEQYgOH+Tb/nIpC
ftd1oFkHWM5FvBsp8e5uKuyWle1PPiXbY0mf7HLZFq2mb20OU92TR0jg73QqC6Zh
O5CAyZQJ+63RX5kINiXZP5vVxEA6Pymo1bRN8ORQA9wWbETzrGFdkSEFrxdFGEZy
XU3gjWrijvqYZiH+8WPOlduGCjcw165FlV7+HfDaoGIxVmwtKKJvg89fuL6/EFvy
JYg6kvan0WVTCilcCPWzeiJclqqeqmtoyMBVv7HHLar2iWcC6jOhe0zbv/PjCLVp
xbLYxsFHSCpDGLjHIT6pc2hXzu7/gCi/GZVrrEK1ZHJQrfeBWTdOTlv3yWTraVe4
AL9dk3XW2xkoqDcdVKguHAHBgyxivLij1mP0vysmRPK2C9GvW3NpZyqmvn6PX289
1whROG59XP0x488EYprRxvUrzGKrR0pRlCENAGvAw3l+pBkw1zRrxLF9QdjTyxbc
GAUfS+Ke9DwLtLwCCRpujxOzPlX2pMe8QrBfijugRotfF/mgTQ5KiQjghYqw+7NI
Wl/KdKcwqS5EJ/IjBibgY37wOm9ngQ5yLJS2acJILwXsNP1UhG48dCtzi7wwG00C
7LpoOH5yJAv6QBzihY86l5utOcucCQ0JhbSIHWEj9jAycN0NKWeXF+j1NXB+a8BP
T6zniMCPeoukpPwuO9N2/DIObivLJ/rWCz5XsoICPmwOMGYX0wtI3fKz7dmIWRcM
B/1VUPgAO33n/kAOG7nR6yAf/4NkCo7jIjf7KW8RvxNLlh+JALQ1e6M3z08c1JjM
KQRlkz+GXqty+boq0sUQWNSI+jWS+lgACrorJI1RVKgXnEE7LFbyDszPB23uqHDj
5tMlyi8VxrBKCIa9+BccGjbDqq4ZUn9HIjkvzLZoZiHyXbnV3WIdwa4+DjTC6W8j
nADBt7u3ExVhN0kR7SpiMxup31WzPqqbJhTN/d3zNyD1Q7pl8rsh0w4mtBPlozTn
9kpxNWQ32Wu+d8ExfvnwXanIuugr3RUG+/6cyq5K7MZLVIhE27WCe5ePJ+Dv7Vpm
1fx5JNGCDuF0QjSIHjdHqqXxWC91VHygl1EmIZv1HbhCnRZsep3Mb1A5k3oVzZgP
kTew0I/Ump0/zsRdPObFP3uL7dOEF+uCANIgeZ9THfzLpSFDqbjZVJsLbXiegXNA
DGS+5SkY3lBCx8U+0/M1qtmgresXQkKVHqjX/AvTYFDK4u3nHrjRZTn+wv/LhEul
e9LT8TWDIbzre6qqsCTwc+DL32oT/D+bSKIpCkP3GbC/MzC5TG7yJR+YkpYa5Jgd
h7+aLxmG2/tXWWUK5oDwXrgUbI4J+MwsM1K3e+lYOs1d/j4Y9BoTHmhLzTF8pKsH
8TfskVk1gpvDQtFF4UrRYDQiQl9m841IjFcYcpCMe0FxrpsAFdk+riig94shl59F
ku1i9EkBlwy2ORJ9L6dS9LEOQ0OHZtg54acW4TbaiajxfFzjuo/JHBv4tLtYEP0D
eFuWxox6zELrPVnAI8P3vwyS8aiEHqyMOiZw7GDGDa8nGmeVgnEgWnldiWCZVtzs
lB13Yi2ekFlBPUpBIPc0MlUu1KjsB8hGIo/kNRuQhZS7HPcH+RN5t2QY2CZt7nQH
Vz7VntjqbpvOLhGUz6nHX1xAnWP8J8QUeREpIEpyN/KPXvy1MAC2++xEzmeRLKgO
9UPXBtrR3IJlBeva9V6AvD41c15jTd+LlGpu70pcI+LxQalKLERjKgeNXzz9HbC/
bswLwJfjFLTleho9BdSRbvieNeVzv/GiOoMd+oUVTwKnDxaKuFSiEtddIfDZTnlB
XdLR/R3qCglHpFoXJZPfzYGKHTJRRJNlZFDz9ULfKYLQYOZO/BA7gkRGGXlx489y
jSdRQ2AskOfcLOtcFVUrEINKycuYtJRF8+ygBGs+JLRqNccYMKt8DsCPYe7KzPmB
SHWdyVCygB7rVnZiHo25/J+eW/zjm+YSiAbBsuarTqExibUszFST49r6DcCO/lcf
Dv7jNOxb5aejf7K6UDHIqH3JHYeP9WiO2JtbeDjBvwjE3mibNfIE8POSzFI1Cma6
wJ0J3yOjoFEuKRv0ovd/75Nt9dK0StjQhSazNnB0riRPxRzxHdnY2bC7PPutspmS
QmKT0vLFfPwG7bL1cndwBasL8x4pFFxqIWcKwchUKnahA64jwRzu4NBPwRxWJn1p
MTftu7gTaDKSygQcCA1Zu/BCJnask/kcMx6pMldopA9SX2Z4qHegIcCN3XJAoeUQ
ZwZUFbHlk6ia5jXn3ZCxzS1mjxK8cdPpt+StLHpWyYIVY+UIj1sVy2LTFPzTx6m+
mZ+iU+IoD+cxWSdIsoUjHtqf+ay+9PXx0VZcXZPNBstpqe3bXk0QRwPBK/yZwJTO
ep6NR4r70M4CNPyR/EwGZSoj9aJV5RLGwYCMxokMXcmAfbKpGLHm40NJxWmPlyXp
Jx2bN3Bm5uJV8wNfk5qX/GZpnJV3VpuOQi19pipLWcnqh0xbFzQem3fyZWV09vLX
Cc2FJSZZ1kzKVYl3N+kRiV+AYLKSkwwpMY097BiOC0AiWL+R9j2tRR5oKRJrGJ9J
2oLdrvAOlbhx+xGAFR+4aqxnXjFf8fe5R9R8BnmFZigfo8NFOZ40Hm8VGwqyEqLK
csYjTZsh9sjGC4twX7d4eaMtr6OqbixHuN4kEKmgsNXntSyEzP0/p0s3vF4bk+Ew
qI+RoV9vCcA04Cgfs25XRdq9Qo6TubO5B6+K/4KhH0rf74yYDbgS5PltL/1/hddc
JM2oFARa4ivwy2pRaJe8NLNF8GgJz+vdFbZRud1No+aDY3rQKfsw8wNR89oL4SEo
YKOh+qh+T3dB3+b7J+tibiW+ZEEBd4t00aGEUFewSKkisbLU2GBiED0FRIQWlnn8
XnXSJ95U4J8SUSwBf871kDIiaIcXDg57qm4KXfVgZLd22LLtMpvuUTiVzmtoQZ6V
J1mDXdzd8U4ymyGm3i8M56rr2sGUbI7N4Va1AaMjYJoFlHwls+6W8eiPLRzfqYxc
L1foW5LY4ox39MwWHt3hoVpuzrnBEKMk7awk25E1K4Hqc+tvE/d7kgfDv9Z1kg+b
kg66T4/3yCXVzHj1ja2OlV9A/wrAscHG9DKMBs7wBshScNkuYyf3LdR3Cl1b+nGk
lOKOKA4TfQYMZMB0XxSQRHAexQ9+ndcPvOdvMr5ayEN4BLWOJgTd8umy8pSXJ9jO
MepyD0DwK+bqiQtOI+6d7T31JZEmMTUKGeTmk1jRmICjE/7y01+NKcVvOhsYqppD
3Qb4p5WEXUB9oBXDgc6SCpTJGNeLuJzNCxdW/ECnMWS/FeixEwsCUMHDFiq0qg5l
GhiVMl8lA04CClhvpHLBgRTNhxlah4Lv4p/AiPl2XZ7H0lBUC4NnQSCu/glVh7FC
5O7AR8XeLd+9+pJitBX6URe/J7s37YyepmUW8WEfe+F2ECAmSR9MZ8vlpKzpc9Q4
NsVL5Hd1JoNsCcOfzkokW5IalrFbRRFmpvx0zxwbG13unQ0Gfb8QHWzLi+qBJ3OC
BReHDB+q2ky+4MLXMPcejIiOpvdACNbMQXwRx6Z7f0FcZn3U+5jEaKuwCeVPaYLi
cBpCP1LazvMjDZrFgpaATGkhofl+j5QlGZLNh+0enxYtwcqGZDKZqIQ4mnoClq3I
kSpJmwul+VjxYn1rHSHtqwOYVUDOeJ2WvKY0s2sfGfGAkNapjq6ou/XZLXwgtdaB
kUMXqF0OHkGiTGh31hCYc9km2J54rsRqJeSrCXS/rAYkl24bSsO8hYlfDfdBl/sq
g0CEqmqNX3qktmxOLTWsnWrXvelKZMbyNWcBUeX3mK2sRkR0YfPj6a0a2z1weeLe
EMflIkPO9Y6JcI1FVnQtCOTjc/J+0yYh0WWXyfqqZag9lW1M+gKNxn0hmLAbaoM6
MmZqQbQooQlsONPAgiuafb1w21T0brmB7SUlJGCp4XULPvrHRnDacAMEw4r4hWce
UpNn6GHGRMQkptEpPvWoMUf36YSrc8pdBsyGRbW6OiwBCtyfuwWkdRHSaRIskaEI
adH2Q88Y6YN25wjGvp4HDGrIyN6AINw99F4cFlYKyo22HixpWYC9AXN2I6IAvLgJ
LpQi0nObzSlG1+9iZhyyVSX+v0gO2AIdiu37/7sYJT28Y4a6HNWXtcS9B11Xdaw8
Nlf9urL+uazZ8iyyOZYpLqJ3n37YF2NYKiooWI7Xd2svT3O//SkOfPRTOVoUhE9b
C6ROXkPBvj5zdyakWy3XG3WqujUISHSgWtQOKaep9I4Ak9igGwTSWYer7A9SPKtn
ucH34amC9GKvpvcPD9Jm+ESK0GV0NQNcQhPzLJDs4UNCqrqXoukjYNXmhlDVzQX2
C8ZZU9pD+JQEYtWPM8FiuKzmena1wU0x0PAUiAAraGg26LqIebkisCaLbG28Q1XO
Sz/auh9nIC6Y85ylF5F7Je8BPmcuOPSyLCrfY7HTsWWtvz+PLSL8jQDfi0t4GYXZ
TfqsN23gICbwCis+ybyfTLKPDMSWPIQmGWFmNUeNdKEc7sXLG/RZEI2qxkETfsol
TXkDjwSr94rGAZ/zM6eYb3ligc6CkdrxsgyCSXrqVBw2DYJiMK94qpk5hx4x3IBv
mvLOLpJrGe0pxlvJu0vGvVURUHMiwQY5POBgX5ZvIxl+R1IUAYgbbQ05fFPGlxvr
Yrdz5xGiD3kKoxtOIYEI+y9gdySJn2GU7Mi8MJWJmcJJQi6lCjVeUcIpG4qvydRS
/PKQFRAPuQEMi85tdp9LlqwWUmuZ9IgflJN+tj7SwnaD1pfxYQgV+8EIlOrdY6nk
54tDrh5s9UJWDnJoZtbD1qhI0nu0Zjjz+rEzJyJgDbg2uMR1S85k6/0y3j2llN/H
F99iNlAQuRsIsc1qTGuQmv+53q48iIzsl0AHs4ocTSk9jpuafgs1vxQ1IIvxPnZQ
xeof4UpZbQRfVSHZUR7qk1d0kzHYbK9GH1Cimr9zfQji1AXNZbPIszj3INdc8PHx
DBQ0cHlGTcAMK+P4wGETiolMrJJnCDqdxYLnwyUme9jx4Uw9scIyFz7IwvfbQofU
Ilz/Mv5ZEUML/BJH8lPIG319wBYGsq4bKTeFhxG99i2Hzqa5p4po1VdChJIrDY1K
XKqzgEDRWzuCBtKVGZ774M0K9L1RLw8vd05+Tz5p1ivBOwlfsuJxET/kw12lwgW8
Ret3b4TGOxVyolTWty81Msvgvr8HYJPURJadJHvDRkw2IJi3mNApozDXLKJJF8TP
XN5Bf51A/jFb4C41mzcvpEg/lVvORS0KugpIU918Wgzf2aEFCfVd/i9bxaBpU08R
hAf+XLzIvWrgSGIFbSYIGy2s5F8ELrYStwe3shFT5UE5dSLEowMZ0ACUwtW5Wafv
DPPop+PLxUxSCYpZFeOCB3Ef9eaDhU1bO3XTcHwZQTD5FXxC1BxyOAEVFOIDx3zW
4gbCQ0wem9i/zJ0P0SdQORT/QhwZYk7b3zJ8ecNzgogECxBbcz3AS7ibkPYmpA17
7uqBLQw/JDaMTLkQtr+41YGbKn0PKC37CIGZJ/L4Sp7cP5uN3aDuJkGqt2uFnTCz
7GMMtI1oH4td8HZgnbODrnvxmIiLx5SK/7NWL0Rzo7kqCrTRikZmL1/uPplqIJMK
pBhhzTK4+kXpprHRvWds21FOC5DeA0YXc805kqF2Bzkzwdl1HrZcxxzxIO7NYzW+
m8sN8Nvh1L1EXn+1K7apOZ7DxZ6wqf4F7Mo1Ol8E97814SA+EiIQeleKxjV4O2Zy
KxQJHmxjkOdF2bTnLFsP4j/gq5JakPIt0EDpTc1FHhWdC4rzr+nfjWIhhQ3nkmJn
FBFy/sbjYYu7iE9YZUD9CrYdfPAXnCFXPt3+vIOGF16mS3Msb6Z9XOyk7fCJ/ZVh
cGUtM7xF6YwthnYTEOM15c35wsioW7QUXwAvuQjqWNCrRSi/SjctNzf5qgqqQ7B+
kv3lb+Y7jSSeuI2kLmVSasHs37neCq7y8vFlXERvBzf1+vPZYphMtrg+ZQjygsBa
hDUooRuH0lS1ZKzEr2tkzKOQJ31ftv8Xj4l4H6u5DJNCCMCe5sm8JVQSbUUoI85u
2ixvgPSJ28f6ncUgEqcS2ZxSU29hsqY3/VntEQCBQS4PN2wBdU9uXhnUq9V0TGQe
SY8lQcO57+7EDU6+vtid7ivz4fenholyS5mWdohUbQcgJhEMqThC9HJdE4LYMgRs
xVeXjp4CV2wWHJFbiHHELKs0SqUNum4/zKFwlytJYP6Yd47DZK5bgeHCxmRX0VB1
P3NbIlsw704VvK8PZewLN+YwsXwECV1kGvjccXH/5mulZrZIUtzRi8GHu7noxtbz
FkZMCSCzwKKw4MU0A26rM+HEy87FM/NtrL11zIDPvMHkTj/7M433aGPeQ/FN7mpT
oRX16hrGd+WPvAADwC9ZC7wdM3Nli7YqcwsZBOr3U4ZA0q3fDA5nmSDvVN7T7/9a
bGlThRQaGH9gVTF6KYjJHVidwP2H0BVf/fsLOWgDo/UEu/S8Xmz2o+D9AwKaFtVo
yCb43WiOz1oI2qM2iszvEwDnc5wIkWbWLb05r5K4C2whIuUhjZ+hVd0vPMRqQlTj
xDIXWYrCphj9h5q2Klr249ol3+oI1XooFMKM9aKwbGBFmoc+U5aq24XH6Qxp+l3g
1hxAP9xHrdXyP2Y9l5XWUildO4wvaS82z/ma9qSYWQwAkEHHOB4jgvBg/27jbBUt
xySSOFv0hSGY+UzuitWcFVTyW50dePSeVl5IY80iWPxU0a5MFE4V2gZnAhH5EBm7
Z9/zmBqVpkcmIyFkjElicBAMl9JYpRJUxIYk5P5CBcl6WGc3fDrpsnADn6LQsgO+
zndRuDrC2FlwfKi7wZq967dGVsByDwvZG3C6miJ858tqqXvLPW4lF3EbUUKqQ2C1
JwWFevmgpnoIxE4iLKJvaYzEu26AmWD2xotvpEUbMGBOSqy+zNk9OR1y54DjkEmw
kiM3kKWMyYQzWMPIfHLtakiTNoKrbGqcmd8Oc+cWcf8M3tdUjxTxbhtinQEAm9su
gDJ4SWD5DMeuByfj3rYUzTFJ78rEQI923GiNNWjbArHVBR5zyeLG201syhZOEXK0
/8/BUvN7ZXCu9Cji9kRWfdoOeBGwifjuDxMrngXHDsd4ATcrYK+CdbJ8AUD2Waui
ua161Xlq5m8u2hOc/Za81Ays3aLF+peB9wVX77+/qzoqeAbEfh2Q90pJ4Iyb2Wbf
SOFTXt3B8ukzG/sFwa/JERIYqBEYh/e7odYtNRz4lfcTvDnf2phzd4KBvCBeCHmq
KNAswlKVPkQhkobGXaOb9j9QT7Ex8VKRPhFfc4zbrCcGmjdDDUDnGBMWHPeQKHfp
ap6HIFBZoheKpRSPJUmVcfl+bZ6JVH6q+3UwvdTNNpkulrkpWTf69Gu8ZTHyOy+4
zgk5OvCJsklgSiTxFiMwSQI0f3MI53QP4pHYkWx0C2AlfW21WCVB3cwq0FufanKA
fmWRnw3ZJXHkmfaHgPqWNnkkBECzv4elfRaTR384q4Om/56Tfw+u+FAMfCzGa3sG
p79Be/FqJrgRQq5q3O4Q32PLL80kBbuEjZJ5Fu4F/xBK5SbjBBDlsJDo8ubYFwjU
SK9rVCgn/CpWOd0YsvL0gOZCY7oQaPYY6uL+nZ2UQDUzXrBnRJzqU+FduPP7q/al
/4uNDLD/g5fRuFziwbk8p60iNKlhYgblYllR+c4yMnCcN+ewdJ+0k8sRzRpBuvUw
Dp9ymMyKB+aD5JX+MRBEVDlRQFKLpNUo5g5zRQI/6rI2mBIQeo1B5upNVpzY5iLJ
qemT3N7hgXrYdeGpm3oPV3xl30Dd3nRlgJQ60Ll0kjc/NeSWIud+mB5sUAR7jlK+
O9OBDNukUIoADLUT5DhHxsGAQMWgm0HZhyo/jPk3RcIjNG305gfw2WvmyDQZMr0i
bUBXKhpK8jzU6BembLod8R5StgwtaudU9oRyDD4yT5RQtfoHGQ3l1sHLitgBw2vK
B7Tu8PIzm4FXM/UaMvGW4Yr1LBJdzSnKYxA0Shlsb1OTWUjaH4h5AhXTW8WyWkEB
/eAEFyBVoya6UNylWiFC2dr2m/lqavqVipiDWYaewEhOiqYFW1DmD1mIKVgSkJz2
L/7yBbGE5I3Ho7iKnMcA9WQ09ypdO5Kuv1tcpFgi9DCoQyymeETh3jAEn2dyVFep
rvwNVRsYl/bl0AQsaJYMq2Wfc5J5qEob0HhePCaPWKESQj0gyAw03IC7hZnzNw4f
EP2RzALxgG7M0RTKPgCasP0tVvMxcZomcap3MG6Hu6Vr9ZOucOLcfL8Fe6dW6iFb
KEzKoOOfJyA0JHOvnplZaaDu4WX9HSV9YO5T2IGmkRlkWF36auX95gMOsPusj38l
//H9wo08oRiza2KywA9sjuOJaElxvbV1K7sbzG+oCqTcZrACk0a2gjjw9NOzWZ/q
TRnPuxw+JPvp/VcpHxSCUW9mSs9nN/ar8poa4yxzjWk/3hhuabAa9ZKLxMmiW9hS
gTrtLAhMZuxZsdqTxfPZYltEfNpSBmUiR4eWH8cGvn1h69cnBFyTsBJEFfegJI/D
XtckJXXppSkYbNPhIlLir9XYBL8KPNor4NVq7QthjUusSb1NsK6ltcXSPzGU8XCQ
TXqDaCm/huYlMtpEkSB0ODaNajbr2uFUDjGxpBneKRZD57Q8GPjUgXRjejhZ/XJF
UX0Q5ghleI8OC9qdnpx73vHSBCbQ6UcT2BikQ0yI3m11eDRwDeYDQFKBXNFHsOJH
dow/s2Bph92FessKGSBm9cHmss6sfPuPyFmUXUuphWVHM/HFfo5tf4738Ymi4A7f
NWij5LiLshTWJ2KSlPVNoEULq35/KAmTErzWl0xDTG3jEKcJYPKd+Qo5xmpLhyHl
8nV72u0IdyPFmY+bdmwill54/nLGqIS9vxp7lLnyYea7CMJiiKX4htnsSQzNFrzV
LcTcDDpahejlFdvtI0fOlDF2bKcKAAJL/HD7UGdF8BXE946EypxpV0fAEfTc7qW2
HqVTpYI7ucErt5eAsEHOt8z0ctcpui6DG5CNehzhoOR85O0hfavFVxKVsKUMfAnf
1QTu0PBE+m+yKvFC+mUMOu+5QH4SHMxW8ES6H1znZPc=
`protect end_protected