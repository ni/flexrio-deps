`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8432 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nn7oC/bbltaB6y9f4wbJdgh
0G6WvBg4Flfb54G2gjKn2xhmS1OPDhzh8Q6RnaYECbGantxN5mwnJvIc40zkl+Ht
a4RNsyeRwcGBOOf153etHtXkDAbyh+6XNlioxpQYhyeiTASoj9+DVWkMGLMomtBE
JZbNz/VVS+Vo9lXF9KdCA1lN48VTd9/kzQDhPAkDfI3+KVluhCJYewG+buYC5yNL
OSLvWCflgWn8rXrducvM+5tb9dTIpWb7ZqEFSRYUID8mhgh1DVOmZdZjkWPd/pjI
yEX3FGE6x2HIcwXEzqpAvntX5eLfFKlm5gsHEkpBWm1/9epARLlHqd/FyoHkbhlc
tr76uuFOKoqpetY6xC8Bjg7uxQw/xPZ99iyxCwFCX0HYzEuscfF4GgTfOn1q/RFN
/p20GsnVpRi0e1BwlW8dfc1mMh9SpXO0cFYx6Yfh1u/JSrmvTxP3xxHE6T1CtO7/
1OYO9qGrVXf125nJHKwDH4W8A7TkKcoxmG881jrQg9u207AemacnjFs2hWQKr1XE
4A7x68AWJNIHWXM7Pjo/npgSuF2OzEN6BzW0IHjAoYIt1QCV0K0kXkNw9F1PAZKl
BUqi2k6CKNKt1/lCrCvzAoLpPy37jF2Yt5kEvyTaRQ70EApT+PDejdIwc+Zv6ImM
fMBVD9K8EpEk6alnqw7HvSOwMtwn10wZrma/OmFnGX/zF8TKkppGtyweFavHJ48I
firMABv2v9QvMT2RVfYzTog3HNg0/DaernQJ3tl54u32t86Qp9as/Wygt8SY6+Te
+cdr1BOY6rXFtzqG1ME+Nf0wZ84cHJOlvSF3AwKt4hyE4JKdlfTfXzqyhdeRqqIf
sYv4w1o36QnwhrQnnmLcZR2XwOCWoGS+I59E6QoMz7d5i94iijD9Om/nBJdWeJ32
j58QNxWE7yjVztDDJHfvRw/qBTISoW6/4p4bXTLe4Hk1o4ZEpvGd0Z/AaBLUk8eY
UP31DaJjyz7VNli1y9Xe6ZWdpYe9jrrUdtS7aVXOO6yki+szII2j9J9HPzDBuZ1+
MVzOm+acq9HgIyLJUF1roYDhqVuc2sYu/Dug8Hq2akNCOCsftM5Z/lD8q1nwnEJs
MKt7gTMBp8q2ddNU28ir24AenlxA8Gn/RmcYsV63pX1BMJ7b5wyYRAH6jMaeaEjB
+E6HWHg+KpRTKTbgKc15BYYsZPWRcSiW+gspIBQeSdPUj6n84yrCcNweFs952W0v
ZpARTuPgOsxonNckaz/WWuYO+bV0n+lLdpAh+8EiwyeAq6p0fOS9kFweSgmeZczO
Dw81gM2eUaNJHZY4EIutplGpxtKn2vt+p6MMJApG6Jj5AD71Qcj2CHVsmKXl9Y/K
4JKz20Mjk/7zGaS1NVFcq5HE/1QIEZBBMwZaIP25LD6MmDoAGNsE0P8RRuqqq4vb
cJgPEeaw1s+TqB3IgPyXuzMivBxbXgjPTwaHi/jS/i9FiHiVSaKVaLyf07AR0xKe
qicEu/HuXGw5OzwSVU/u+4hMGpXN1edchFm047Qia88G7VtGSokLoj/t+HZfWKdX
uvSa3Qsn/kmfE6QyL5FVwONjo/rgLw1pzekMnw1Xd7pWy6Hag+4S+LlrkNXr3SuW
i5y6Y+XXj/Ceo8vSKzOYPBBmD6xbqXnf0CFqBV33avq4lU7JDCRRXTl9WRGDGiuT
qGXHjWoYtZLnhiDX6Isy3TYYAwfSWe+AtXR5o0Rke8HTp42G1KVdrpoD/9B71TCt
uWW2BHfMUfZNHdNUyc6HfmRKGyaWxxUSZjbFW4VGRwLuy7gyXIdS9pXgsPlI3SV3
tm5nFlZMFiZCrxIlprIS9na3EZW0mc2XRrghCtmU/d6lrDBKyQ8+FoJksVsFH3wq
wBf5SOZzzjvjAGsYeIhB/U2VegA15FitmZqQSfqYU3Y+u5GtWZE7rGe3FMtd+fST
uVD17+HE3aCEwC1Dslss+VueitrPZlgKdVc/t5tA70unZFcRT7IktER+CY6TejK9
BZhapzWKdxDEDMIlxq4FUWO7Vx4gyIyQA5uC/8UV+EgInP+I0qR/ZYneF5IRRgc5
WrzExAFA8hLLvjpHBVI0t/FUig+wo0xjuEO0pjE52pi8ruPJPnhUb7/BQeO7FG9e
DBU0CNY9R36rvgK1Z+qKiw0Fi+nn6CAxUFVh0vdhpOj1DPw05FUmA60j3IP4YxSp
yXBE3hswBvPlobKvQ+tLstgTG1tvmtvXEow3JMWhbNt5iA/yEeOytQqvrvH/DjGk
Po67a8z5C+QSWdJFISaaBSLkH3JBQYWVqKm6bVN/Fc/xw/YHcqDb/EkzBxqwz5DV
+OmQCDc1tWjRQl+9DjtcjuE0mcGdDY2iQSmHaY5ZY07uVBr3pDlT57iZ01vDt24F
ZuS2rvrTMzVSUR3HLHZuOghJSOV+7Of6FsvGgemRBdlw1As1kuvmBPj2X3VjF6wh
dUWvYe6+w+PZj2bErTkHkUhbbNqqLobzc82OGwJPis4/IrsE5fJEXzg6wOJwT+fJ
KNFg3551+6Ed4hk2adW+11Zl38rh+xcpgWEFYbTXNyKkN4xHL0A6Vw7W9O/ke6zD
fygh09xp1fdM4UKeclimLqZYBwIHjEfB6/tBlblsDsgmKmj1APrAlrpMFB35O4Lg
4kZopnLT08ttXT87mOW/TVZ3lwgvE24SUCXwpV28uP42qVVWHxLsFtnoINCWvsCm
8wei7XFG1XL0EGqPRRonZsleMx72eUG8mnaRdeNqtSd3vpY3+lB2M3XAUktGuvg7
2Acf8VJDT4/N7Lt2f+YiQa1qr9inJoLbDLIRJLC2EfHG/VdatcnoSJaCFw1fH8Tr
GkLz3ycTmYMM2H3x91IFV9GZrSpmvJeQJ2Ti5OdrWe+jJAWzBKnd4LxyRqddbsJI
eEVJjdckDnx+XK1E5X6J/xg6jvLl5AegasAG/cg0Wp0r9UjNRn9wZimAKMFE7sNy
vwzNxhVUEc3iFNfhGbMPkl+DelDqow5NVwtwjFA4WscCsB1/0YF6Lq01zt2oPAiy
xES3GcNcgfu0k4AeR6ATAE2V0k1Q1wDhe+kmuec/HNSqSXxD2Zmkao1QDW2NQ05Q
PyGi6zbhvopJIDM9dKOSYWNAY2StdB+SWiS/U69xA+LTXCZx3IOICqJjFLW0smOS
2BJIfNd4eyLQpCyxSOBDg6BiPlTz7Ba4inKPoH+7vD6Hs/q3JSmA2SVxvB0sZ034
JIzFrXqpcW9R6o/c8+UYQedQ9ewZPqPl9J0FY/Gu1oJ3Jseo/fZejmfRlORf7vJq
3Jy5l2XHsjNPLSvnFi9hYCWl7OETvgnhhJT7N42jiJ2Kuiw7wcUyoxRVnt3NYp46
zIjFX6QpAtFPtHvABPw8esHTiH01JWMcDl2B7MVP6NlMv6V3+gL8AIJH+3oxQBeg
0LjtFaO+ePGsG6XpScmOZ87BwLUGOrUOOevGbwFYtsmRN9Lv4VErA/61XyHJebNh
CUhSmjtplno+sBZ/Ey9H7ROv3fp4vSDQzDBUWh6LylTAyzkd7RuYZzAsDnWgZCIQ
lOjyxo2vtwvVVZpHuJk8KpgxkX8lJ87yIAkIhbvWgMJQ9Xn4Vqe57FyCjlpiLj48
gRoUhXroqoblwnQnygfMWTqyqzikifd7m1A2NwDKxyxtK/z1elZIlcskSh9fZ3Ot
t56YqT+nZtjs3rIF6mo1pPA4jrsxuLSsPJ7gEaJyekfbDIQn6CZ+3yo68nNWsVQ5
6Gs2GXle1cOit9lOTVOOvzcIsvUr76JWWGzddLht2Bar645+5xR4Bz7EZ8TP05t2
Rw9sMMLCMLd1iDjaflyNeOU1KH+blY2DgqnGafgPRedoiF25bFwJvh0sbCCn+S4s
SsVM8gRlzx3TbEw1K4lYmFkhvrEeF2x804uQKqKntRJAcAPlvWuRnojJxLpRwFq9
EnS6eN/C2BEaiCFpWFTvSM72NyPRQCElRytdkrLjKcj2lXT20XgrNmCDQ/GMJoAs
gbeQYxwa5r9DQHLthxNIJaJUftWXqBLdNeO23fdLPFrtLuVWN0uWXWWzpsUrYRA5
bvlYNyDeIXu/OXeZsnWyc4bJyNPsAsN6Mxr8IkvavXJ02bnO4sR7Gki/GRtIO59N
nT4LI+HKeDXw6Bhz81nzLlzWj87NrdreKSEaO8nPWWeyChLFvfjsQhj4b4dfq/iS
4YzBZbNot41l044omyCADPVk8UsgA3cuWFdp/Z72eamV7UqhhyoFfHexzzUEj/5d
AaVdpZoCKSLIaqAEHcNp1OomcVuvmLluVxm9djkbhYNRJ13S0LOlucAKprYVjdJy
QuNlZaXWwQbJyjioHtqELrYIwVS5J84ShXDhwWKC4w02K30515ErIxZDsCT0oFs7
MXBfPG4/WNn1eEhjCp595IzGlUjySnqZjTJbGG8r2SwzivtD150OLuMWNTVoFf1f
0e57+X6pWeBblG2OzddgTFs3j2R2CBvADYBEhAeEdFQLPDf/AGqe3kF6QgyZjlea
W4XkT13AuQEr1uVV0neN9auuZ4SbZnB7jZl3I2WoPWXVAHK/Fyp+QccyTvwWECtT
f5/j2Vg5VP96+u3/zGBtLIfV/gCOucBbqvUTGUfoD++XoZkJ4it0DKEXzOlOHZSU
4CPufDjY8zNz2tfwNuIXWscm9YZkCf8GyW/K+8M+4WHfkbP1j68vzJ2T9jk49+y2
/6z/jnHel/AkWdateZFivunuYBuH+mjm0orAWWqSW3ZpeVKhTdH0uDyClAFzF/m+
opjE1yQ4Bia6fYAvBwbhMZWph3aGjJfGGRTRmx3dARpZjMcqPhkCk+VP+fyRLtAB
WYePnu/JmM7wGLfLqIVfC9wCzzu/UtFt+o/hx8rM41hN1wo3dSoi411yDj1psI1t
pQ0E1Vkq1umnW4P8rIteh3wMqtWoeURg0JCErdcDF97IfhYqpD/+cyl/zL2vxgM2
yyoSV8Cf85NQWLSo0uDJiIkWFdcYy+AQZs0qHOXsWs7WLXs9an7luKD/z4ORUv6C
KikAyohvhtg4DyA7HpYhAV8GvqxiozNKCRnqefASx/mEireEOSuvn238TsmnN8QJ
D8pgBa7uqZ6O2SO93Yqr/X0TxOn9eEQnpjSqAzvCj8dqMgPlRefvJgBa3i0jTye7
nL6EGGrY8Frf9VKl+MWHhXLt7wCv6WMAKRh6g0b9zzMGwaI3/o+ibDkitR57INzU
4Dynqb+vehIN0JCTZQGnABCG1QkMMPiC2wTf28VGRiFV8Cwm0q4t2CuWljCcRIY6
s8cZTHUdejJLS4ZpriTMfeniobzieNLH0Gl+hFkViLOZGQb5DiYFHyiBDi0R2cr4
LKBGmn6GBzYQM6VBGsLuPPRXfAtGvzZcH/51Gwg2/zXBuUpwPSmofmVFJVg00HHM
J0ViJBmln0X/1Dya4jgsZoivJdJdDFChKjCOjsidxIM4Vb1P1OdFeTQ3/+slK28i
+MWjAYsuafN0x306tX1BKPlJMlTZdaGbXMTa6JUO7eoDEssBgLLIj+DRddPnMGlO
i9+IhDmZ74MVkfLCHeYNe5br8EOE0OAv/3VwsO+dLoGju9I/vOdXR5KJMpa+AIEl
vdzbX2F4cl7CLJPueQu1HlNHbLIiiVqfTk9QQQMBqxWnRvPXHD1CxCrxNZkpIw+F
fBE4BAkNk9C8g/qgRvQB859dJKenmNpLGtC0g4enJA0xGft/+v89xU3SPNkiZLUT
S3TzzbS/BqBUG6flaJ9kPl1VeXHUmj9j1FXdrLpOBjUAR0HdRkMv9q5qquO8kTOu
xb8Sqfhwhhs1HtbZOQYjx6/CeWRrA1nbHi7e3qawx/JQihZeIjbZpFejf7oG8lFB
6PEVtIL9x0V6tBsDe1cVqy5ry7UwmsFRzCvgYUDKszltupaC8OKcmf6I3gwVxRab
sZPCw3346iLsifbybvcBy+XXWtOfvOOx1GlIqzz+vzK275kglQsm8h7auCbzqFOc
FVGyabo15qyLaHjf5uI4SnokilluQ4GKfHdAeYqHUYEwpP0CkPXPDeNCI3cmwU/c
c0nEJsROVdi6VWFi78GqIEyZpHUNGgXDlSI/RWKUYn2KmxWouHClVkV1W1eR9onJ
8q2sArBNVGUFOh14mCl9/cUbv+utfQkLvpnLFpKojP2S8PzjXXovQDbEPIyLuIGh
VE1WzOBlhlmSyaResJogXvQ20Bz4+VO7GbvufoHke7wuGVwwmp2j31vr1QiF60Gp
SoxMXbeon2PZE+bkcyJ2obZVbmLtsfRq9ValBoL5mFfmxgjnBCjTrelKM/HZk+pT
uaqTLSRkRGBq8erxBUPZ5CutC8SsM/foQoob5VltYVIULS9kexlq8d4bILy7N510
C3Ajw0je+76C/iB6SDBAtcLOaiCbl9b0m6mFxlqOaa8bVcST39M3Di8V7JmK/4Yc
cpLdy8qoKQsrqaNFNbXwa+z7UZ8NaOSixOZu2BI9j3vsS/QhYXJcHCsXT4y9A4+8
IvnuNCiwzSSh/wpdLBIxjuxSZ/+37vExAMHpebIeJjM2A4dUB84/DM1QcN2+evFp
6mU6GyMXD1Ex0+HjyH++Lc0wiPRIGk2UlI3O1rI25fKtCettxjwdFE6LCyAyP1h8
6zNUpqaOOQPRASVv+ORiTriE4lLYUeTYQUHeTSfLZLT3XuabEFfmftk2L3sRWDrI
Vn3+/VbnQ6nTJvEGJwW+pj1H9KtczoLsuxmo4VQP8+uLv3Tc+EMfnKT3+RVukTaJ
UEI8Hegh6zunvgPB1CMLF4d3hXougxVt6oUdzKMuiJww53di4BnH2HVVNUe9PKu+
SHHl9KB7z30jagpoQ+TB7A+96uiGCNwZOJcUDKU6rtgeLJjU/M0xpZzTKKGqOep/
dn4UgmPx1zXKGJRbIVwd8CNtIPhIwBl8xEnl/qbAtJArSFCHtZNU3CsOWsryKzZG
PtY8+cU7dGpZ/+Qr73Y5ZLG390ao1ncAEzVPpP2GN6FaABjCSuFtEQ34AC1Tp+B2
uLpgpi9oclmbq4PGSthdmAmyzEZo98k1FgvJJ9z3s0T3ZWMiF2sc8ROjvZYphxDy
EW0Sv6d2b6ebW/bbxmWS5kz0Zl6zhmWeaWxeLAbI5p0rIP2Zqo6kFSY/OZzQBoVn
S5hDSzC7ZqWJk368p2JUL6lokjoiBm38ltWUaJBerGaJ2R/4oZiWe53jbAChLWhy
ZNLDhfMuug1kSx5fDx1xSBVGMcB/ZdxYKwG4EwyoM/l5do1ow6NZZq/JAPF1CZNC
dpkM3krLJM6fpFdR0iqGaHOPi/fX1/jBeofDB4l8GnPwW42BgcmeUZwNV7jToNsL
QPadC1I1DWBVzg+QXML1Yb6XJ9HhUiGzBXikjBiW7VeCrkxZZGm+JTtPwRiZwX5n
vuX2752aWqrHwGAA2IsKirpbNY5V7/vgQHl8mETPB/plNxHcIKqLRhq6iKsB6QgV
ZJdygpkHR8+cGL8nTsEghAdzaJ/qH6xOXjeSF/XrWhSphwUg9TcdeeEj4Ba1sOSg
jiJBvT/V8b9GQLSqOYzW3jm1oMHszz3xLQm7gRfSD41OZthAc8Q+EL7ZCH6Rnq5H
RpAoGzW8MrfLUa3kVXDUdOpcIQxNDsMIiyeAOKIxot7Yi0wizFVv8eF09mbSaGqL
L8zFuyGUeFeolaR5d/rNiBxotV7+iFbvGYM+XYEtOKByXAWoWsc/s0M/ueW3AC4Q
lYxwUthDGpzDqfgspBWrH44s1nt5WGhAN5ldQqh2yAng4bN6UFLoCegyxVwHdzAi
vprpP8GGQviBWU7Po3miX2Q3nY6Oaz514Dzy15e4j0NZFjg08WPkWs4cyo/qUO1r
MwXtRQqnjNrunkcV+4BIDaejJSRTuw1Oa6LH8w0y3pA1XId+bWuRzqYW5mNMbbaT
kIt8Sr9+xK63j3A2f2I10R3Xp2HlyrdkiUyQbDA8y237qRVtOZEPLVTUhXVZEyht
G8Ttkz6rDQY64TN98YOAPrmS6leRH1bapcPhCoWYGxy47m0rDlPl3vxDZDUl+Ytq
RWwbnzGDJqQ69o/T/CvmlJ894MmoOwRDY7GCBgmCGktml7uOBN+zQ85XraNpW9CU
cC1Zb7jbUWA/BvSDeIY387ZN72YZojogz1R4ccxUP6Cp76eeHy9HNBGnUkZtCFja
6qZwlo28MyUDifCthFTWfnEzT/sRTuL1aECtClnkhLI+SrT7MdzMwQ7TMi1m9wTQ
zqGvT6OXk174SNbl/90GH6o1Th28+bVKoROlgz40ZDuFqi5IeX6AmjoW51I8fkuK
ckxBZb+IqOC+1UdHHsJawzj47+6ioPCwNWmj8Wws8u3xZanBvmy8tWoPI7mie05q
oCX8MdP5/5Dr0DHl3yR/HctXlEs0iI/stWbI68WNICI0JDuBNUQFk+En8vGYRZTy
zjMv/K98/jjxGAc64V9P9n/zJA0DL+iimJ6x3J1C5kuF6r17fxMPMADVhYnKEvqE
Q7Ki/3DDhn4gmpQs3iT76l/5qt4g+AANALpmjdIvMqqwBBdSlBIAOSG3auO0+vMW
lVVRjMCn1lJDTdn08F6I3/rxu6VFSYaeWlcoD5PRM7TeJTH1W3leLsD8s9Zy0iaO
YXdUAvXBmO3ioeSDz3LyKy+SHBD5ZSfpe4SjT8S2bxexOjjSmkB4huGeTasVdx8B
7oFoJ9kWKN5dmSgXObxd+Gz3J/t2suNzIgV1+wRhFMjDtPHjQ/uYBGp40hmgDMhi
g/4TPBQ3BE58SMTrN+Mp9zNVoaLAHMN3pv5ucy38cSAUJRpvi3Om7BsOBFr5f+Nl
QQu3c1xfP/ocPM6hAcAm3v+OyEDDp23dwrEy0YY7VssYP4I+lxMJzOVVsDVXaqNs
c5H6bemh8TcaQWfaLaqQzVT+/zMyUib5edeGzgRd9dqIRRtNlAb1PLlhWnLCRChO
NZMR/TJPLe2M9wteUcHU+F31ETUymA7QtpqHu76goiiFQVKbcZJuvOujJIwVQQZ/
aftkoQx5N4632I7aoR3Jjd++d9xFVndnZIhhQSmBG0JWhyFYuxQf5QUGBto44LLJ
IV8T6wADiHSVHoI3BYwAvJxAwcnaB/dxEKv113NkLaPZTpoW51ZtkCPy5gixkCmF
HH6eKUOSF41wP6qquNoinz95ESbssId2iEVBOdIi4oVWuGQ0g6EUF2vcHQoFYJ8K
Nt8B+oNfrFsRDRKhswJUKpXUZylkkOyUTPgekCh2tWPhxtsErnxYz4Fn/qkR1xdt
Dpn0F2X+Z21+4lI0EjzWHxgS3tJfAw1IFhXNsWLSBUnEHCLK5x2Ck517SgyONFAQ
eQWgFWOhRcDeoU3x5vlhGQgyfiHKD3YwZK+2qPfXgtlUQpYH1xsPRjxRPkhJ9Dh4
7HAKkyjkow8JfF09HF241S0GtFJLQdYFgEA7oPH57w/Ik2QRp88+BO+7WefsEMND
+C19O1oY7PBJss6IfrcT36Ukwz8cIOMS9aMv1M5+E3HmEZ72s1ym2zL2wkwDqut/
54vVMgFK6izc9P6Clt1NfErn+Lxcx18bGSAahzAt/fDNs3ADSg9AB1dfFP5aKuTo
eDkrNdhnjGC9SfBWlN2ojITdpyTYSN8yP+uFi60cjb4NMwYFWxwQLbpft21SIpcA
MABDyHQoGRvPWqCSdsxv+ML6ds8dj9QYcSMWqlLwniSjXaQKwXnx4FyzK+hKghAX
iqh08p8xP1N2ZzfCPrcS1zz30RyBcGpEhaFjIvubJdJT+Eo/mhfqPBJ7+HK9qWQA
JtUzQeFKUhhsis0HoUfsAMxwbkEdoXokcTC4IfiszbSYDi52DVD8r8U9rrAJAvL9
LnZOmI+mFDFFSfWm3Mdag2MAeheZ8DjntE3wHVKdJieO88o35JYNWYEVDOoGUNDU
sIC+ENYKX/y1tSR0BupHi7D79YNiaDVTdQpabRmSqEIR1eEPu6t6abZr+HzVS/mc
ZTaw07LkWMCu5S5zC9s10mO+mwyi/XDL2X/H/DA8yDdHpNjuJqk96mw8Wfc5g27b
grxwusLspXf8WWvnQ1+1UXziCkIAbGmQCXp0PlrbFEAUgR5pib3Pl/VQ8p8l1VsO
Rjycu3A3XYuIW8w/MUwTxU2JjJcuemium9PtX2ckra2gH9iHJcxfsibcJ1NSQKEF
u6ZViE4zeWpJmiHQhF6yX/Y7yL6O674YsMflQQsP6+shJHmWrCt3MHozvyZhwZXY
0en4SoyFneZxq8PD4rwfMEWVZ6q2nK+EGmI7mYsaFmrMoCiFDDE0FBUsTZuH4ueM
2Ah1TGrctkp9otqTFPxyIqAbTWUCmfgRtXxV5K12JA5cepAFRgLxSpvGVfzpVn6r
MeC+u6a0w7QSKaODJYqiK7qq+fBFeSjJOPLZohvHUYko0djwUg0HE/h1uFF5e/hc
6YlrSiFsYdELocq080Ea2IdcsajUonqPWs8N/GdxIgolRXog81bCBzs+jEC1WWYz
qgdqRZ/Oybf1BOZNBgBotGxei/GeJhpOeKKKCJvCIUwQDG3r+DMsavTTkNGWnkyP
lHHE9BuawMJRugWbVDhkSBVaE6G29qAmPEkA24mAYJB1oJ9AFO4t3JZphO4Y43fk
1gPzrpq7RsBycDVhOpqdO4HznHvRjv7nlJFlVQaXxLpje44S23Mkpk0IyCkaYbYz
+8X5hKhCDwxNWdPGeUOC9DqmMU0ICwxXN8pLLMbWLOhupXsNKQPce25UIew3dis+
1nJ4CuKTJLNSwWFw45i0LvEENvNjlX/IRgPTlnSGI4+NdZq08FMxZh4fr4KTVl7X
aGYshQr7Qt95H8Ry03tALJoj9o2PSsIDM5BpvA7T62L1Ugrd3VY+E/wXgXRcbnne
CVX5XwSaQl45ABsRuo9wzGPrMYHlMeEhin2PRLgiKLuW32sAW8T+Uhsgg9mOePXD
C65GNyv1Zfl9l0+8UX00/p0nUTS0O6p8SR6XNflhVvegZxXd1xb0aIkvBOEHi3Sb
tpmazJqjmeqNkDiKYilAKQPflT5j2SuBGKWcNLfHtguaGoYRf9Xp5p0vMbfYp6v4
//bCcZZ86nua6EipXtiyEIEQl5pkL+d1b7+PYkEMSBJLJvqPgSsu3LbWSZ3WF4Mm
P3u37W0V+S2vkrk2rxqDA4/Ng6M36YefJxZ7X0PJe4Q=
`protect end_protected