`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5040 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
ht7yt7qgZZej0S2R+oiVFTDhGBfirsPc3d9Kv5NeE5eOX29fRaDn3KLZlvAJs5lX
XNacwUQgGlK7dtfg0UwvWgUJpbuFOnobPkd504cul0wvmerakNtwjDOdWXeECu6v
rKO/P6t0flvtcFEwyu5muPz5GrBuDlQCi/v0dkSypEFO6Xi6WpjVtgVSEO1Ub0bA
tSr2V+dQDXZgG5KHAxyo9nISGP3utXfv4V+HpYPQP1GlvUfxJMJp/lyQ6TaZ7213
jdaYMr6z7mKT9oLmhN9FoUItvhTeDMbXsGunn9KmKIx4GP82V02d58ix6qb2X4wo
MfEGG/YyW4ecKsQBA70p6LvkiGBnjpHHUJm29WxJ2nuocGrVeP3ONV4chrnALv4X
VMGysTc4N8fYcwJW7fAUL08cgpMzRKyuYf6AY02ovGj3GYxStpf5LP3WNcTtol7G
/4b5CZ6AQ9QYrcwgrEMD+Hk3Lr6z14472aEIICup+Z57rGbZ2Tn/1d0L0nliydFK
chlAmN3vf6cinuwBKeAPRk1MnoJ7ABQX+pW4QxUCE0luOMOxSbjNb+D1n+nFu2qj
hrr2y2oyvgWoHGbYXHryMM7iSbryzF+3vHfRIcMl2016zXRGKeVMn23WTPAQ7OJC
lulC1d2HoEPcB9C7mVoe49qngEMD92yDCsg0mnKCoTl0QejJe2TM9/Ph2WaV8hvy
58z5yGxU4Nf3og2+i0nVR4Agh1yVhWhYwa0uJ00TWr42bTzCwduyB3GaCdl+j8pu
J7zqnNpYc29uTN7a5wE9e5MkRJ/XmI1P9xXvbmxj2pDDZlCO6stFEMM8Rmx3Q/8C
1Pak4ydDG8lrKuGS27YTFQm534C5MxwD4tvZ9pPwyE4xdXR+pgUuzTVu0jMo+He0
tdeyeWy6hsu65iCNXb2hGVGydv/Fv7JDEpPK71WW8k0XjY5YFWW0+tOJGFU/WRtt
d0l6U8jwxOWfWsFPxFRZAYVpeqfBpgq0WUXPH75jOC86EAOGWhm9IDrXE9E/h6UU
f7qVu7wMLP/7u21CFOIcHKUAFH+pQu+ORI78NfTicGLr6qbhkb4STVWLsuRBaYH8
m+2/2iZL5LgYHmYkEHbM4NvLIZT83v+qOA/jgAPmCtwBxbCGrimXj9HNJCeFdjAJ
efxR0L7sGI9RhfSxQzI3oKNIfZ4Rd0HKExOh9JNGNyMt8PAY99yC/ZbkDlmdrzYZ
lg+0P8CGedppIdtZk8WJRCtrtRQZ2dG3PTPeEKJ97ourH3Nr3B/uQhNAGJKvIbsN
tmHDDPEzgGGPxHIpVC1ceG/x8yumJL3vP6doe3Q2of4yCF9osUbpdt8sMrXGfL6G
DhHufki+Y2FpNC1zVpi2j8ApVKt1PjL+A00CT1wnSuUhIA6S/8QfiiuuYyNp0yAM
T4Boon3yxHH9XMjWmsM//cx+HGVxtqOTsfh1MPAYpP8Op7vj269E+FB1mW0wG+9/
/fE4knGyBHlLdqmrfK7cLacRsJwCA05wO+tSpTF1q+flVk8StWHtP0EfYY3RTOgI
uScaG4NE800Tnhw9W08ihWghHGzFmyPJCeW9FIaCAe7k884cQAXYDixDgRfxkY6H
Jm4nzkw+oVCbIYSlgd46nCWmm7d7E8jE/gfgwgAbadIqI3JU36ZQwd2c2JjEBmkf
V+n2fylxcVKQ2GX7rR/XSe8ID9nbVniXIFIGHWbTcC71rrqVHYqCWq0LV7u//FFk
0Dkug1MFAq23oB26d156hqSjqczbNQ1voRFVsClf4SmTrq7bESzFB6scEu/k+dpI
+AzSxPeTgZ44ZVigodPzRIWwSLRm0C+UwEWAt9ANicdxUxPAIp7GIccVwJc+MnRH
TYESlZP9p7WBVvrzv9vmJXGKCMJTCI8exvsSwifPXzdObPHGKCqcyJDT342i5gVd
hluF2U9f71THKNTBgBBin2DxItd/h/a/dGS7V4TCaUBuuH480LN7MozEP1b36M8y
uC6QyB15kXFb9Zi6zAXacXROEWgwTPAImUcTDu5AXgy+x7jHmEtrMSx4yjFNuWJ7
0mFFe15AFVaFU/q7LJzWGvYeGEOMd2hDITU/l/V1QV0wBiCWKBS6W4IpZmpPDvxu
ixDYcg/vW5SsKMfpF+5BognxhyMb5B5dIY2YgtxplsfOx5EH/CJN0QCdQbAo/ewk
FZ+0gj7l6Y3/g7Qon2TGNubVid1sNxcd6Qzr3P4wsu36p+ZPz/QKX4FXXgDZtEQl
/z3CPwOkZypyNKvqbGp03IpBxjUTS8evyANHvAYFG+W7zzx/rcW49OcGl3a1tQl+
Yn5Ydhl5HhbAqqqfd7pNEVI89Ua2ZsLiKcqy/MOAFV78PCbs7PoA7vesx0D+tVlH
MkG/33ZX7XZh/N6Zl1k0kj4dyv7kBpBft6SjNdDKNgrD0QQkX+jVd+k0rs+3n2Zy
S6ewU85homAKuPmqrA4Kb6bnQBSoCLkJhWQT5riKvBZqIeAxcBPr0cG6Q2PK0eso
3DBFXPB/Pz3icZo3a+lx1tHTCSnGx+/MASAeU4Uz1JxLf8SNx+LQPkOcsXMSFr21
o/QPVsD2UAwgeAGIweUuPfCvoHXtpnPwRdQarxZMNKMlUrlNU/qrQwcc8juoDTmW
VA4+DsyHNWKQjKr9S4bZ9OEvoMxv4zwoFOEQ55maRJdfvdgIwRFsl2XFGIxks79F
Kyj1JX1kIeSb/L65VuMRrOJFvUVVP6CHrHcaXiT0GMvKxIsIwqjIG954RJIMecze
prCWRrh5U9pRuTm0Tvu7F20u+YCh666IA2pimGV5JoYWpUObCMSmmds0wmn1JPxh
pMSuKo+cTgKLwRkFvlzg35YJaSjcxd50z3GOOEz+4a8oVPN8evxR+tgHM0L/gavy
n2GuyyiE2waBZqidro9NFOwiTibmRzkqr2V2/uzxJUSEeYhPpzo2IJrTydZDsTws
Jj1IH6ho9Da+Ng3RpQX1VYW7cX+MrSMQujxQ0gHBoxGpGUrw8mxhVTpnpTZEBfpR
eYY+1Lw2Y0Dv3ibWWoEz5yzsmsf6j4+oIn+hBn5Fu8Lo/UvYhSZTPNzob9QxI/Y5
mPsryperwb3CA1RRww2FVXPjSUDOnxD7LMkEw2ZHCJuowywRHsOOVYzeqou5E3Xg
Tq94PmHKgjzjcrWUqDPbePOYgSwR2QcSMx0WnDwJ1mnuHBCnixuynRLm3S7/KQlF
2L27rEc7NcwO0WOTmcNFl4StAZRdzFTb8B0bW7XWdZLiD1QfcOnSeZp/Eodo+QuB
duK/Qp1HR86cArsA+jSueR+TtPq1ATcsEqrHvwrDSrIaWg9TlP83Fhl5SOptjjWX
JxFDiRB1sYrx/dxBxCMgLam1W5QoUdIkOiOiCKwKcqYGVGgbf9yNQBtkMvN9/KUH
138C/HNna3ekvsDghDsXr1yFe6bf7HVwrR/cpfEWr4QAyV42wUW/63zHRjRsImAP
HkY//lhxNb2uIeQygi1JmC8nbczyZ7TU4n0omQJd9QzWbRHfXmm86Ftg4bDFDrGy
UZDtWoGlURkV2x6PghY0+4fs1e6Zz9GwykNqfzqfDMAsPrQoglIxy7tYH3YJn79F
0kAHj23IuU4RtabWc9IN2l2XFyDd48MXlSRYVgacvP0KnWeLa65r4VCPQ9LYTWtO
RS334dl2rD2PXmB0qKuv6KngZgSBHE3C56nzDBRrVrbmLMTjZazDG2Pe7TkFqRHV
bJYX7pIbQS1DBV1MZrVArgEkhy4eXAtTD/rlODTZ4FuiD2ODvei47MNQDF2JhyYC
b4DehPzjUVzMsAwfigU68jHi5IS9vZjZrOZEWH4K2odeQdsP4JWqxCixtccCu1XN
wHUaNef60uxF+fKddG1AmmOENWEaPRqyu0oMOAuWgRAjznNcA0zpr27xyEZSRNfx
vlq/V1JWRRl7ZOlpslicE22l4Xta2iCs7WvdtJ2m09TArqyH3Sj8pKHaJJ09puub
QgMaJUWTkK9uJCxGhvOWuglZ+N2SN7fdrzr4bjyoRWUVTb3QdswXR88AmUxx5E3M
Z2hlEh1CUKndbJGIgWHndg/vuvt8S8sMrChZm6+dxljCdB5XrKP1Dwl1m5eGacJP
Osq//oOMjwcM0lBX6ZSoxL15hcGxgpqGwtf6BH+mdQUVXLo5DAmS8bTNVsbGYRkK
RXSeejZ24isFTsoEqOUEMkF+4+65i4KGA9nEaa34CerhTAxgbbI266frhxPS9bA5
cbf+mhsC42qvExjgeSBzAemhNFIW9BjFjQmSscuW8QW5eN0rqRUw3AlYo51tcYT/
BGRFE8HnJBg5SFN3h5BEBrmOTJmijIXOJ/WYCVBORgHte8Vj6UfLoREDlLzkisgM
LIzEWaFNWkW6D5mECy3osPArMfhnitXfjBWPg+PpOX2bzdUxpCOFNt6Rrc5bLXbO
VRjrJPBZKU0qUNOhugbXGbGDYQePlJ0iYizpzne6F4kjFQum77OxSBzdVAMtnp8g
5lzinAPkIhFl52d4shY7aT7lYpDvkPlXrAeOzImCeQL8wn7ZBDeZDq5RlJSspQly
9hwxwlKc4VNQ4g395X3l0LkKdV5wHs7rX9X2EBfIiKkHsylxWnWWi/o0rc7+HHdV
SAaGvqJGD3y9dngiIEiB8Psafl/ZGIoKNuT38LSIkBMKMuf4v3ZD7HjKA2WQIDN5
rxaX+XA85injdEVD51e/+lfzCcQAF6SZxOXUn/UhKH8Hsg9IgPD+ydQoPghcZWyd
nkdkti5oAHat6HTzTkvvhAxXrZSJf4buwfIIg4kBHwQpDOEA5JBQ+VJCq+x3rKG/
Jhx4BAY/C7Ybil3syOTFlatMKfbciCjX4MjTE0ce0b/qKGjBp/lVWdIiaCla30Xt
hKFqhcqbhVtZm5E8fX/x3lckrGypsyN4y71hU4d8wGuFj5HG9VEmVRVvyZ76Jh1q
pq73Oa9mdlp16xGWZjLyqucDr+iWvFxWvncB02+IZ1hG9Vz+T801HRBzeV8IBHil
1bMRr3VLZqXRntuHKJSbvvtpYaJoFRNe8brrQx/Ut+pzj/reWO/jvP/odb+BbBPj
BujEH1DI4BBNzq/gaYuC3TcvjuIpALNEFO5fgldEmvcNxzIZl3n4/6z+GytzwxqB
dY+lRp4SYQ9SnTbx2itUP7IzrWMiMWwFnQ9KBtRb9j0FSZtRyccN5au9lMxXTMt2
P3r/hOd8phhFo4qDc+mA847G+xHe/vgcIzNjs318xP9aR7BdaP/LhpoK0c/LxD7U
ueRjN1l4D7NF1qKaJ3CLTuZXWOEFh1KWbfWa0thZAf+8pF/MMiNvfpNh3nKCLUrI
lKhmT3cY4RCzTHx0AUVkFormLPUMUQcDMkhIqgkR4Zgi+YnLBx3avSAqydLHk0l2
lKtX7grP1SobjkDaGrodEYKQ/70NRKOIN+06cPl7eAlfQI025PO3ONH6tssSikWc
0KcKrq93HEnqoRuknt7TPACgOqpe0it596UjuARCB/jWqcoZMrQWSHmtiuIwuioR
byOrm3YRVxDJBe19I9UAIoKC1cJsmixrgYfjRlZGcCIbAaBTq5kd1k87wgY55fPe
IsAXKb2j2zY99nzFw1JQrAJy9OzJ49xkpfnbBm8MTHsAKL/QwDy5A71rHrjlpeU8
kav8sKh6ru8pIhvyDuRc+ghs9X9j87C8xehhhqdILh2ouYrqyU5F/dx6cqGUH2MB
uB1S/DknazMxYq/82oY4TxwfAsTEWV1Ld0L1nEBVlih+7sMQhgAP1aqWK4EU67G8
B95IfvHU+VPYKbji79nEakq5CJainHcA0uFCWl0kW70MgiCxkLQ7qHp3XJi3ZeiD
PDBNOuEU1+TCks3iX7ZPoWrF3FChaxXFH6xi/sofcsKFUSXiyS8P3XqdTAnvslPk
dqDet55F0jrWpxQIJKEyYbqpSGUxKPc2NGVfQAeVi0QMB67S9kxj2yjIfO1nqx7E
3YI4qTbvmi7iDpAAbZXHvax5kFoZnEaqv5sPVczrZ8SHZEWQwL8pqEDVJHiejiRk
4szvYKTZcxhNdDvN9eCI9nBklbI9bmaYLJ6ruawjh58zOsA48xRss2lH+NFOZkM6
x0qgPZGq0/JEMMHZeqoT3FppAzYbzEZa7F32kTT3mT+emJr9juSP++nAiL5dMZfF
9P7PiuKdNakR3BOMpRzh7+HRAYV4vVof93Pjn/4XB5x2FryQ3iSdHbAOlVdAnekj
1eH8zvLfAXLZpOt3l/OkNzIczHPNWipykXlOY17upQHH9/LeDCnvzu7WFGg99QKR
pQ1zF2gx3QLUJZS4hA5EtIfLfUIzdAWUoLZPasaqvKaECKdOqS2B4SGLUQrh28wV
J5VQMreUZE0GQfj9Sl0IDr2AvWxHx9vNC4lscRj/jnDByDgc+eldM4Pp+DxlyIdG
2Xdp/28euOs7Kz5LJydJW7qBItb3VBI3edBYKB0jJW0k4b/L7MhMYoAW6eKoDE+J
1CjMjkdo21qZ4yVrzP0wIR97gF1HHjgs2m+stCpdCF2ocmqkD9Cz7hoxTG9Tp3nZ
yJ+8Ey9snQMdszKywAiujlhJjUCWqjUwfgadyC6jnqm/s5f1iyoVjkEzCKNvQClG
`protect end_protected