`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 22016 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRpv2xRODiJMNLGiSdcH6P4QhuDRbVm+q8/H6fw52YOaN
Lm5QfnT4GNzUn0LF+8OS9XEiaZxa3ti/7GB0G0D6gwSMGaV00+FHbeznhqJR0n78
G1hZAh4aaiQ3WupFCMaCOJHDLUrxTZJqLQDjuau0019lGLK3FE6OZPF9VQG2u9fh
XDEi5Up6SJr287yKvJ2WHC0WBoDcqUmKcBoRmwxGRU8/JioGkZOgooIxD7zCo/TS
I+QtzBToFqEk7UdK5QaSeoIJyzuHDyTH5FcbwgZjIrfUPNAg2IWR8yVeXH5AEZU8
Nfaa4if4oSVR6K1OvyU/cKwklDMg8RRxKZAUud4589JXayF0GJyxKDl2rKOgiY+I
f/GVPH1Mn3VMRgUJCxutTI5gjVUiZhdPC/OS/WEmA0Qla87G7TAsvxYVzQbEKJvI
DoTMkYpjPfNe2cm+039Qkpu9mTb22CHKdappsV5EQ2BfytHoNIFOdDB7Oa1O4s7+
8Ck4jyJxwtjPNlABSkybiJ982+PYIGH2Zt+VCAT5bSK1Qh8uhixw4jYATwlC2Qpu
Ebi1yM2th6XuPOgrlIt9c9zWaGctOM9CW4JGZPMloi8ltUMrS0qcaFFCYv6ic/Bh
knY9TajuUQduoRpyh7r3TWEicDvAYvjPnOnwF0Mr6U1lw6VK4t2UU+XmeFabtavi
wZDnwglVLkFzDGlJrfPUZM8PsTP+QKKCzKWgBXwLuLfel+EA9ldo50lcUZljZwG/
JCyTaKcwNSwqhNP6jfAxB41JE44A97ZaGHS0P55ckIN5gZvS1ywcZO8Ev06Bz4qy
rz9DV+B0HnKTLKQ3pypNHtL1cBJ7fatbum0qi1xIt8Y3EOhT91CUtYNQF+d2RITi
t9x6eCPW79dWdr2qJ8PfUwLlNf0lMqqY0TnHFBCsekUdg2SAXghn/9CB+Ro5x7QA
+ynnfexDTvB5HXEzRamk96tei5Yxr6kJEUwrCjdXKBAnUuCIvuhFtxlIG9IW7zKU
LkVQsQ0ZHubZtxERx6WGgjKcZ6zytO0l7jFVDO5F6l4rGGFnuIr9Go649sQoUNLx
Ew5/8WYo0rR9+bmYLRJNYqtBNuypfTlmQwqzVaXvYukDKPaYBzTc2Ap2MZLYlW1g
/ecqxowRVSZvh6sRtyIlMEe/3/xD+nEQseTHICx2bc/M+skiCpaZRkMPiZqHEfeZ
GQZWwNqUlC0vjj6OApji0m0Yd0/lwAO8w0ukH4I4l6S/CMS8f7Id9VwrxivtHJRo
mxWVy2JABWplyUUeppzjVT6Te1KEBsA/HSdAXYLQgeqK++ZRRlgoC7bstNIU+0wT
GY+F0YvhsmNohy3jO5Yxa0gssOEFDoddiGKObThcd93lDYmdPXhRwtn0/zkZpoxJ
q4+jJ5lT/nm/ntAjsG9/IcyXMRPu+QEIAGuX/vEdoXygmK4fQXDzL/fB5YtRkCsF
8zEU8yo49etKjLe6Vovj9F+kfzPbvSc5MMgTHAKIq0TaRSb9Bn4zCHe2u8YBYU1y
prTV+1SN2fcy/q7ek1PrCO863FiCUfAnHPbhMBIe6ieaE6etKr8Q4506KcUk+F3V
l0hlbETZnq3FDySb934LsSnw7asaQCnOyWccCUk4z/Q7uhdQRPVbA9SRcs2EZb8Z
oFK9amFEiAJnkK0O8+8OeDbYE7e5ct+yHya+7JFMzXOrw4F6Va7LR9PYgbrTjUjK
wgOkJZCVNmnn+xzPw1YR1x9IiX2w4TCtxMU3hXNerqirvDrZY/3Mn+10amYkj7Ob
Tg5v132Ud7jK3lobSAZG1oxmfJTAuwE+fmaFIzRH0sYwM1dCkaZaVBa/XRAx0sGa
dtUoCtBWwp+qswwgqSCgXDpWFS9Cq+l5sR5fpXAzFuI4PGQ4nBrlRiCNHofnuG4U
zKlXkAEa42hH1ZHBWq4q+GRvI9RhBOVWHfjOXWU4+UkqdkzforFxlszCeWGAqbkg
Gd/FzbsMfm+mOxIrQelTQ7HDEd/gk4OQtLd1ODGCreYkyvzjEMb0WOfZI4LUUD+J
iof0PxwcGf1AoyMom6S1yGUUB58NVZ10oQVjRgXhMdlbCGhYuzSXr6CJowcGNyo5
GIaS+B7XzljiFFtWyIIrQNxUVI3Pu1Ok3C36uZuMhfsGftFuGgL5q2VEHFnZzHK1
R1nJWeaVfn+LH0j+33hX/xmMvnx5tSk5DJgkqT93sYlkRKSUgNC5zPVxsVY81SnO
q0tdmq7J5SXvyXPjAUmi8ig2/19Ec8Sr48ToBjgGU5U5Mq7HyqLPC2jxQmnuXNR9
GVSliZ3K+4C2cqHx1iJUAduwsjyCSKhXCkP+gzAdGkcqU6IHwCKV8Iu+RdV7OYgp
wokv6aeX+gCUDnEQj+Kno9L/Y/gxdbgu6PNQ23OdvL2IgnlrYVoZkReVbYzSPk2q
PoyisGRULRjQKzB06ZhAvl0aO8V5bfq3oi96G7/re/fJm4jdfG/Mkr3+89XOBD2D
uYnA6+XTD4mO6b9Zsx6ZdzkD3C2DTJmYkmciZ6cW09412YDQd4QOjlOEquAUsfKX
ZuEQ4NkF/xZHC1rsDsCibqEt/U7rq3JPz0L/rufTscPili8dDpqxcfD2ynniNPXJ
MaDdOVLHYK3jXOA3HY0evalaLTgGcItYfo6RkqfqhaxN/yVm/ROmkGDnrORJPcgM
JOzMk4X+0ONlUUh0Sd8uI7BoMnX9j/+EuUWBRr++scrsImhXwpv3FwYYMZnWS6t+
5S1Ywxylbdy8MIvWrzZX08Isqd4biv5EFcNLFbblc1xilWdtRf8lp74b06Wda8q1
ZTJq2Y/Acl2xSZICmYn/47m0NxKk/UPZgMQa5dbohXfKYj9rm/amY5YYjgYDbWU8
DqlC83Yx1l9fzxZku/v1MNoK01HNtuLwqp0wd0hGPYuykGFo7mHm+En1QBXYrdkk
zhOAKeNnaKqFtY1i9Ua2z6HBMol0+xyqYhCeVW6QcyjqeFRRBet3ZSK/Ma603u+U
fipfgAz2AFFp7LSfRX6PQRvVlhZO1rHDR+4MAeSpNZ2c5y/3XbqzEmGrNgC1yUrH
A9DbEl3XFTtbGs4vp9byucRe6clcmlUUf0iNSsob31apU8CPjO+i1FLHfWmyUQQD
tN0VpexA39pGlW8aUNe+EzL0OF6orAgVmxOboaKrRapKmFY+uvwolSI5awiWf/NU
NYJpAd2BPuqNV5egqC4Th+UOudMtxPvK2OgofhcMposmH/ArTFLovZQ5sDVTVBFs
OtLIFJv1reo7n78nb4Ojx3ZB33Pkj43c3eYUmB1+iAnnXipiLo4MLk4cshRjYc09
Yxz0Ex2jw89V/jlfPoD3MYyQ90C0fHKFaTAjegJ4pte0uGZmxtmUS5wXEUrWJ7ap
WY37oOGTXxgRH09eNFB8KCB4qPXtajyn4AhCwBbfA6Tlg2hnRej5dowMuFSRkqej
5jL8daSfFgSjDk0EuuKhzhsQiuA7/WBLXAzHThrubx4K2GrM0tmqT6rjoIEayyKC
Ln8Ek1IAnzT4+rVTDMLfJdZR695a3i9k7HtKOnaSx+gyDXyayeOc5y1ZexHPypXR
mCWvfLKw+Uixcw8l09uMTdaqx67sXiWcDvKcBu2lT0SHfNLWdie5nllmoLvVq2JS
dGloTd02WrL8plTwxhhCOp7zQOw3W0xJ1WbxBBkgbDi3KfwrgR+DNZphe/w2KqHY
pCR/iIF/yoNKrs/mP4dq7XVEFxwBBFuF12/3fle5KDXvIkvnhQGu1XRfIn0Y2W//
QPBwWOQw6AfwnZkX5PKpIcVWS+eTKFONNKse3XJpOth7Xz20TCNfFUF9MCQgIXvk
WVDbSbZTAHCuuVAU9Fy0HQ83mlkGJC5RlzAzVsdHv72vUZw/rD5MzGv1OBesJI4j
rRdXUkBboeB9Yl8aq4u7c+X8qD+FG96NiJt+CBKdqFOxt5v3CKwyFvrNC/8dlW8O
ymM/xUIry+PM/lEFPG8eEllADh+Izn24uvXwu4dTQEGUs9aIA4FU7KJLYGU6ZDD4
3OOpAV19A+St/kDl3qiHGiVR9X3PBjgrpD54s36hU9FxZUsC5eV17v2m5TYRrYtb
TYpYwd1LGVDX+ZsZ9T293fLGhY24m6WBToLZgwPWhD0tfdjG+DA1ZJUvOfrTeuTe
Qe9tqCkt5WDfs24VA7P3MNKSnMOCleyVmBYJ5HPbHCDqAvS1m/DTCzZwWyPgoENW
6seahkwDtUJE1iQhNfgdA0lVUHV8TRs3fYD/y3t6+N5Ip93K5ORnjUXoQcHaPzFZ
elO7aHmnnU/TUqTmuKoUNfq9o87wSWl/bTDhr+7B3sUwyX1IX5zvTYyXWbjP4YXr
tnkiM9VD9vOQu3TLKg5FVYh/h4M7kYGGFJto9MunQLgpgCEZWMk3jaIQfl/w1Xcu
t+nRR0+NnDS1qI4R+XGsHyZls/AHNYWouRWy2FpVBzBcDEJlyYBE/jq0xzofK/rK
ircTOFNnJU237WNakTHX3zssa0lvxgX9pUqzX9DJJuA/OXLg0R4h84L3JkuOY4y/
0vx4Re5nbkOjto9ZylSiJaKi32zEwVW875GXje7u12lui/71OGH6WEQfZvWsvgub
hT+LaDzz1Uvdkj50+s8XdI5tV6ILAo0BjTR7NBfiORkLkdvFmvlfKV9rU2kV65oH
dhupcAU6B2IY5yvqq8mgR6X98qvuEkkQ9L+6wrfI1qi5g/k7xFPjm1Hxt2un1GNb
VI9C8G7Wyv3V3xhgJDxH7k6rkzp0/cEgDhqOY3yagJZblYr1pKKe5XyBzFYEhmwp
FYaqSp4a2PodRX3sK+7+3u09WQTrmrOQUlFLshc/vAO+HTHxuGVzM3wShR3xS6op
JRraEdQRdhr+fs15wHOI7YuGexhPEcvbAnQNrqK1yOGEdyzK8ZUQ/uTBnJxbu1LG
6Q5dbvSRist3E0x+KCXCnKQJdOS7keLg6E8Mk1GewAjTuHrzsuFB9bYaqFTW8B10
HakXhYYb+w++5RIx5Gwaw47Ix06Jjh3tEe8Lrc34VLEnczVkLCADDMTjZyi/ycpC
H0rTOleBzq9TEfoY3InA9W8vUS74E//wf6x0uMCQPtHjcYdHvKhhRYRiAKyUIKGB
H35qt/eY9ieGjWG7ZkJFc+xcIyS3sInOF5D5W+K07bBS2AxYhL3vtFGZC4KL71PL
qwTjZYxTiNT6GqTVaV4CQO/Lq83eFbIYkZ5cgnN6TJgjtgRnudbNmCaPZbnh8Bdk
nlVJIDOZJsHXCnwrZuWcoukR48fd9wUOmN/T9jjLYQ62i3x1TSotac23M4OKKJBR
ybh8aZVleUBzwq7s40jwbuwpCwcLpuGXmL60CoiX+UYRxlD5GsXdNKJBdWrzfKnk
MTUETa/CJ+Uc54EtQ1S970n8dt6zDl8Amu5Nr7N361ZVEKgJLOmg9UF6ec39zMxh
uPQeOeLu2ALrrghIdXkqPK3Q7n9xRvjsfeJZMpEsSdsK4xcuiv6zwUEmMvip0UCW
BjxAL1dFeyH2Q7JAiWSmfUSffLBiKrT+qd6iId8bjIAqUYq4TG/YdCD3RjaJMvDt
p3deQMfr7Pqh7Zia8G8fRIxB5QCVkVOS1t3J35g/E055AQmvOwkTp7BAcpS8R8qt
RbEJX/QDCNAsdSnoyriVKMLcqqH4Z4kKa20ENEQbcuiWya5OdWE86Rxag+rK7B2C
RKb74QxizWPqoQGxyloOyiJ2jSarfJ+VlgAKRqTShwTpwIlOTieb2f7j9neSamiF
u2q3uax3VF73PG2lwpsAAeEEYh7AHs8g4sqPLfMRQBZTg/6ki53d92bo64oG/Qyt
CX2CUa/mnwenZGPqYqxqf58XDWmxsNdTjxbL0rwuThyckf1v/Xm30PnJDyD5cG3g
9RkbZoztIyOuFvGxYI61cnBwd41PvQUxFkYOR2sUzu7EI3ELN5JZGp+u/veQAYXN
ujMMUxQr6tkJacdUHE7vbS1Rg1pLw4I7Xd4AMk26fTaEJY32auxy58m7cOp0ZV3i
1+WsSmUAyTYouNdgzRyDTppPaaotgzoZbd3zeiILK6xTAuLFr+sBGZKv8J4KTq/X
NIr5PuWqzXulnE6VqUTjMEUZThrcSWLNSThkEurkXE2GAATFXNtAcUHyRyVuHS/8
5SPpODMGsVOOEGBgn19eRL3KYfhkM2gnpgPAW4+6uaXwyvwL0W7ThHU4i/UmRNIC
UOH2Q37KNdv3D7a07ogG2J+cO4YLZJCsz9HWO5WhjFXUDFUb7IPYHNcKliIc6vSY
AuyF4569g5gycn1Q3KFBTI0IwwGD+80gUKoGbtmBPAu5bAr2gLNGALsEv3HDLBEH
x6OSeAbMPa3GZmG4bbUhW16bGqO7KJ/jn5eGpOvDJvrBYeEe8V8n/a4Gq3gAluW+
eXQZp6iu+qEQbjTwkEtNZZIoKnDp0lMu3rXyHRBdJs3iBGebRlEACu9mQtOumhoY
1OuGsXwTWYbjkUcvVfG+HgIhFlTWiYlV/5/1fRwtTUT5/p0+kuWBI1MA/E5tUjsT
iBtxZBznmRb+B8y1L9nsBWO5tin1fzK/R0jBMTQxtqkbO6d/qa1PezQKdwTCxiq7
nOAK2MHrhgE+Cm6dgGqVeuf83tJqngUtaPSw7WtJgi7Zfx4/u73Kd0TmASg0VgEG
vKBlsvsCIFGy60ccKxBUk+8F9N0rrNmM6zk8RRIcDT8A3oGpauQCmEFIdZ2MdasL
35w/duLvP1PBle08sJIcOwqQDecQAsd8kN1qzXFY0oIFKmWUihtddYPeksU3hL1E
aVS4sTFeXWpl6C69ZO8WbxfmsGZ8exMw/IMiw/PazVrvxRiQdsSJqgSQ3OrRhvjo
mZkyvhK/8sss28KuXxvMN5ImQcF5pWexOmSz1oRXZuxvOQBLBRDP+hcrlFekbRVT
dK8cGXIF1e0BOPXt/2eLL67cO6O4/rvQ/uh5rHYGANZx2vUhtl1Dme5rmb87jxwh
fjrIJTDXlNI1zXKx8/uVK/jz6WX3TRDLMx4bzPniu4b6AzB01A/GFQtI48uOImOL
ZuWeSiskZLGGU/4dzMSnaaGep8rraDSZ4YLFnS9a+yHeYr+Fzq83U9diFq8zP6Aq
Ouj7Z5MK3PvFxdOsV53hh7YwDua5orJP94iddVumgGcq2efy3/HiXPQpE40sWzKj
VkrFZEg1O+iyklrRWudCS/GUAEWs7gcMf5T3Hnfbwl0dbLCkCHNJU4UyQvLQbVa8
qMAPHW3/rSSs+i8EWxMYnDjhwP98TX/e2BuDTs20oSVRcDucb0zbnLzr3F06kfq8
RNM8/G1R/Lg7CeycyKX7dPnpqsqwX9qEYa/pbhf0hrFzUT8oc0Ao1u/GU8IDcitE
PlqISfBGJXUYjF0L2SunRfCR+oRWx5Q+KdC6Bwb1sBSF5I4UCAGoMAB3Q4koQDxe
WBNx8dTGD0FfATWl7IHlVz4wsPcP9WX+6d6uuCTixT543xq35pTM7sMAZUtqeu2x
2qZSoYuyrh87KoOQfNP6hiEN1YajyrvblZjJFMr7oNm0pnySL5UTwxBNkqLSsalH
oIGFqievD9WUupOCPT9/WzixQ3uy0N1EyCWyWxt8Lhti2VhUrRabbvRUFsXkGOeK
1VbWXmwHohn8+kIjbkluTYVH4CUz/jvj7/NYBHwVRtfx+1pgJaXibNGJ2vWW2xar
A8dLE6ujlCTZHyc1dGH9xknI4xLchtaHs/gXJJSBgVZU7F5l+qmPPMrmLvyMsZox
6FK8X9ryfgGtyagsQfdQD8N/nwIF1mlw0ihPop9N942SBzE3xx1CbpdmpF79F3dc
gYnHfo7cOUEztD/KMdJVu8iIaIj/GqnMzGoIn3JmdugIMyoBB1kqeGi57Yrg/Vy3
3BrEIp/8UM+MUyhW3L2uJz3nsn/Neev08JSSpHQBfYNc7Dw7wtxReKGzZZePLIns
EG2vcw/SvBjNd/63ZCJM6TkqLRlB2De8la3IyHktGy1AOVmGy8MSYMpwgTsMX2OF
WBCavV71quuanjD9ovkeF4hg2hoaE7nVo1lwiAZrqvey1lhB77ohNwkHcz9CAQ1m
Ytrc9psIauhmUG1POSGv4/6b7t4jt2k0dyQ+mi34DZ6GlqdYcF+Zsn+Pg3IC52hW
ukC/5rZpK5L45ARCFs/e3q0UpMDFbhlaIftyvzj1w8tkUaRYJIC4PpLZYIHmh8Mf
5aTofBa7c0/TpMm2n7ZmksGNSPFJz2P7fO0SXg477gjWbZNymEOdpU8vhLqLOof2
vjoudGaOHUzO8tJS+giOxbpFUgDjWFgvU6iqNypIiI3PpwX1sq4gyJlKYfdxyTta
v9HhNO+uLLpbflEYjraB/Bnz9qB/tYFQSY2rsbPytwQL/5N4RdSCia/eBzObD0+p
VIGTgnE3JuBwmBnGxugBu9GaeO+vcrxx4r/BTKMZ39hO3wGDVnidLvFJN9O/Qa5g
iOqLi315mikSQku3GUhVfDMjzJO22OrcVxs+tp6AX+cP5LppjCNCCbGWnNv4plTH
xgu4qBl3pFr4MB8RQGdhNM/kP2wI0dpbrJrt85jGXmR1qocZtSYY1EHubfqPs1WJ
uwNhVtIHBMFgjW2mpJonPe4lYWCe/c06i2mB0PiPe8WL47AdblcIswIIFETFQRCv
cbvzbxJwJitUqVtG0DY0IpOIxRMBfbhpaEvRwyJFh2NQAyd+R8DiTxwDi/cAnK+4
4GYmBN303Y6nufV0wKfKw/rIijgZJAEkCRgiVefDG3c9wu+EmAR6v40WB8KjW7mb
iYH5Vwb5sxl7nrwJsxc19mdpNhDWrcEDhNatlTwzpp2WHCSKVXyEzTHLYFZtF4x4
OFVRCkb46cRHtw1O+mGWIUyLAlTWC2weW8r35Hikm+vHQmiKD8loD7dzyBHvCmfW
rsveEWwivybXIPekbM8mCXho/++nIvqKQnQQbodOtGb0P3pzGqlYw/pB7LGD44XB
A5RXikh/rp2JzAkjRWzAPWvTskVhKgmJtnZ98YwxZlg3CnQaG26JFMWbfAG3VFav
ez8tCvhZiqilWGJI6D8CxQOiVeJX53VlAx/gw0G7BALz6i4CrDiqIQcofWgahgDZ
OV2GOz4CwExvkb1lbu3L05WNI6nCHZxFlvHXjr97doldzihqxZCHOrmzvhfgg0Cc
9eKlKoJ1On/bqurI/lUJeG40JGOQtmCuh4Z6lZ9dw9SXzwHDfnw/+oDg7BQRmgx0
eHsQ3ydJWXv0SyMf+x+nBHa+PK56xZ6L7eysJe5nSNBN8+1GGAZPXsnnOBzlIdmK
8cnRzz7BsdJU6fpkqVjAmhxLVEJmm8GNQqg2oAfE4HxOqzlTQS3PmfXhxRdMPC6W
tjBupjVpqnZHsvk5l9yQUAZNKR3HMSsvlcskbVpPkG4+iCUXMSYjuOgeH7TiyA2W
ro0Vt0TA5ujYT8gRgjM9RIV6LhrfqNx9cHcTkB+pAm+HGafkE+Zn27vp1WmUoasN
MthGqoA8kf52cWcreqH9HRBRXKfKenxpHXqe2MDu4nxgzi+4do4vkwLB8SrcDlJs
0v9btpk4xPAGu/qo7O+6auSM0yKHlL1yvkpgFpG+/z9EL2WwzWMLjEcWnGYfwAat
iOijtC8YHnOeJNeZG49BTwnjvcu5aJkwl6mh68ap5vYs/oMPRNBIdSMStxa3KDDP
PsYkipwENPyuVMSFM3MxO4zHxLAUaQPMRCfohPJuu5nCr/UlfkTtUqEGR/Ghw0w0
bboRWI1sq1zOSncjJyclpAA+rSM88OefCAIyiOIfaqaQV7NpPiXhXZknSu/WgYOU
Aw5OaD3rcfSXF59uaxLv6HtIgYiYEqna1KsKNrwRnyFk+FzgFyINR0hxjWkx100a
3GXD7dyqqNd3OLeFXZm00fnWe9NT6Xo44eHNuwySDRy1RKAv6WSDSyc3+uUrYg7p
EUd2vBDK801lcxLuH/ix30ck5i9Q+iUzsZ6jWL9L7Dg2TJa75BuN6PWEGR8Y/Sgx
Ep4Rg+MI0MOf2sJ96F8RKFhTlUYE1uJe48A4LaMJwc9CGd50jam+frDimerQ1vfs
BSGs8xGpqSa2GwDsCazhkg6N5yfJAoPuaGFMecHWz28wxBNM5Cvlkj1O+ts2KNKV
cQ5bLsYLHjwIcgK0cgR9FyQmuW1hVqX9h5Ca8QzCTm/i/wx+32WiQa9C1zQcHSrM
wabSQWPGNMZv6FGYzymAOASYo9WtD/Uu0bgbN4GWwY+SjSL0MqeOsbiGpDDPlXMk
VSIuSP3WwU2T54H4JyHY/adHy71241KHTa8iE2Xjvb2BQsRBJf5jktG8FrGFhgGD
CXrbxNhYDM36vUFM9szNcEbo0a9Qaj4TKL0VuPDTXgNNFPKdGjlO/lkaB13yEjXC
c28/eJ96EgqYeVVnbfXKr5lBGIaqZnRGULkrXJThQSf7YPd/9TP6vfJVL+v3BpG0
JKk212E3km6T86as0LnDMsxnvZwCwCcXW68NoSLfylHWm9BYJjlkicQ6ghA4SKBa
l47iZUJB7TMY0paE4ev96KCWmZzMqdkU0yAbbhy80lfeP+4yAWOwyfBDW+fh3qjM
SZa6S6/yjuYtZtkLfeOd7eViuBJX2mkdaNhAih66ahZuWX5kII7EcX5Mm3fTUX5k
5gSioErUHUO7GGDCLKjzQmRsvrYjkzb0TdIF3nGuLDK3ho789I6NsSjTOI2HqnmK
o7ZFSPOPTR0MDiDOyW4OjN2JjT9XjcEVrrOit38O+nZYYp+FFT34iTFvYX7Mhx0a
YU78LdGtDXyBGpAjvbHRFfr+DPVGFaGRJomM9gcdpcZV4Ha/toMTN5uga4bR022z
UFH5kDhNs/wk/T8uQdvPri1rOoIHpMpn2f2VL3KioM1nZKQpna9P4JTscKI0VH8i
QdGUY4KuV+jRdzaf38B1ztdomb7LIC6s1QEc+Rn8Q7eyfpN3CUfCZyMO/AyCHurO
gYEBCLF6cGoyuCk0eftZZQ+xgE7fKhSSi0cSpUdu1Eh6P2MxW2IxuOcXeBCwhERK
MRWJQAA9shuXIDRG1xUxVlXh9Ayn3H/A2oHL7Wwn9EaO1Gk/WZEmuQoT6uT2c3+j
e/K9SaUzFhR1Wb1kEQEAczGrlyAY2uJm5Edhu+KBBgh4oll4MYq+jZd/aXjJB8BW
qkr/qhlr7ph7+uHTk/46v/JJO9U9CCvycvCyF0nVK20m3nPf6cxnHW/+fpo6l9m4
GnEzawI1QuioCY+QsQ0heSL6ZhQMXlIKn94yZ8pBWczRTxQSh+jaxBMTGs3YxqAz
+lYEimGIoU/H8SGgMXTZ1kHHb1JBiczCTxuqbm3Fbwy8Cxy8AI9Mf66avt5uer6D
AZusDL/ttNKadp8gVty6uKwnMsZPnHaU+wXH2+7qTrXKMyi9QD56kOX9dnaX0F7o
cAmGpuRWtfwLk/hN4zEh/aBXYHMii3nBxvmoaP9+Nui+WMC1RZ3GJkgLI7hQQnCQ
HGS2Nkin+GaJcz/rjBNG3Kaf+8p+CmbvnNgFc+69jgO68KQGgRAXsBZVxI58ZyHA
8+pck6iubclqA0/SYqL0AzShu+oxg+nhL18frCd6a62IyW+cW5Un0Ql79k4Wepv9
pZge0GO9NkfqSmdSkJ9TyvYIxRibgBrYMXe+MpUf+aSmezhsT+PxTBVBP7Vifi/t
KTVEZnXC2PCsWmgEvjX8E13ECHNu/weG7hY2bzRJ3p9JIDUE0PNNX72qH1dRkUAw
9LmDxJlrrMCbOYp8Jqs7OTOJvYb0birtZJkfhJetAmiuMRdf7BkbDtP8suBsQ0k0
gNiUBYlc27kEWDsWGFP0n+Faq8OSOrDm1dQRkbySRTU6wNR8IvRepNDIriR7pPYp
ogJglinhAKTiNPjgG6EaYf+sMz2CDCY4Gy5UhxonFpn7SRYO4JWIHpQd/8cCjOVt
WjSjKv90P1AlqfheyVvxHfi1RF4bL+N/zpqfsuC1rG51W5Y4TiCMA4vvum1dFY3u
G4IG4XORna0rhp3arlz4c/vXuFahAVUQ4uj25y08b56uzjNlcAYMDhVXNsFkPPnp
1WxT1s1196F7lMEcrzALGFqARTCfzBIZ24MtyrJgX/U/ZB4t1spVCt4c+B4Blq9u
IdSmPPza7efyL+djHL9NFZtVmTpCVhpiZHqWGaxOSpcHAVGchlkLnYM8B48dPfxD
Ox5QlJtvVjTBc5PuTdyQWel0WS5AYo2W4cu3hvPUyjol5xsHiPJx4TIzYOUg3oAW
Hpb6ePUJ9Nt9GEqKhY3iua5ABWFCdv56A5jcnGcAyKRS7vXGkOnhrtfMSy8es/BA
sYdlEZBbvhVKUcAi5PV3OZvpnF+49yvUC6P63fosD8/iR8DNPH8bpxwhOK2KxucW
sANYDgk2nHDIIjbDJ7Lyg1D39m0/RCeeVzGokv8KzzcSsBHPP8qd8U24tOYl6zuo
eQHj02sVulYZjr7C40rSyIm0WmKGiB2k9NsRYTi6/WAgKdmSca/YP4jtlTN1ALKj
Ad7YL3RB/VcPNq2DbvUJHUZ1ZO5OuCrebk3KlSgchT9hcAIVsji/ULff/8QAGVB7
g67mNEglqCsD1wv0NpQvOMJFQttU+kCwvPK3Ci+J7FPW+Gwdh7+wBo0TsYiQjwIM
eXE9xVhNOQqRPRMAeN8HEu7dWRAKWT1EtWy6jKRP3ndp7vME9AgTQ8NwLNyVeA3I
Gt62I+TFl8QD9hhmHmZFAOiARyeXNYwsEdz+HoeCq1GzjpO2Y3ckPFWDdg6h+5wS
kO2rhDUatylsI9dQkrQFJFFd/Hmy/Dk4KBrscqodgXSVdpSMgpoV7tRrTrukTvqP
6S8fVQ9Uvg6cWnvWyOFiqhFoGOeRHo/o2OPCTJ3T0HK5JQoen12PouWSpiJVLXMp
6QkGTUrFhObcx+fMvVFyUdSvT6UOzWnAWbyd6OnF5SKHKiivlmXJ4RVzMGblMSH7
FjxQeUn1jLmtOwkhBDWJPKoWce0RmrTXZy/K8YoAC0FezJEVvEAel6vWs/n0M3lC
2Z0kXUrttk8UhL0DMUHoLVOjcjz4FH5ftbv7iqQzsVDp7yix5QIIO7mJ5XbsDLPD
PRrkrS+tA3BIs3D/5rN4BjrGDuJuBSCHvzxFUEzjCpPidVWjOSrPnmCy6TmGqiNl
teErIhm6lFKQDTtx7AyvIMOmy7YtDVrVC3wXAproi6FMvKrzgpkqyNsel++c41a2
uVBnKI0lOhQemTdKDzFDfATlGYqkDRzM1eG/GpxU6ORdCrzjoiWXFxh5FP/D3OMU
HbJRWum3W4gEiZrD91QKwI0fPOuqGze22V77//8NQjJS6o9vKsxoz47oHUzbUkNb
fOWdRnuAXG6IlPeDUpaBRs854uXxfx4A6hhFCH1uUUsvK7FGgi0emXFaD8ICNEyQ
7EraXAnsVbUUETxiobmxnzVLmMc7XGGslXg/Rouz8tQ4zTvjsRXFQiPFCCSAsRTz
AK6HgtUyBBfiAQzYy2r8gzjkyyLZJShsAoCBwBRZCqhAnuNB8R34DWQgqRPmkW6T
XIHZKQj1iiXFPtyNfDoF1KzR8Qy5i53mD+7QwsAVD+MHTYma1DzEaKWZ3stOpb/t
P1J6JkzeqZUdoWW3RrUML2+8SGi6V232g3X5iiQnWc+FcOT71ateKPqyKFd9lMGd
8LUIrKyxse5ImS2ARsdE0MmEnMALmzRSxCmR7HvPTKOqrjXZLTgXthkhpGngdCV9
P0fy/pD13b31lF3T+/0OezuJuNG8w/jIkALL95ogGDPfWtHPES7NrP/5udu2GMR4
rvM3/kr6X3DMQKElmb+AI+eHapNPj6kg/yZcX49V8VQMkFPhK/z0bVJu66sdeaR+
Guhw37WKWvkilksq1VCdO35Au0UScsI8Om6DLg5oyJ9WVxTYPg1BJk1ULDZcNpe+
Hb8e0gLbHAeZXJh8BkitLdeGTv0QG7krvEb2nQaU7e8uSz/Clad5vVAo1bGeYpNO
ezrZAY1AUAIS6mj09Lj+RLoGYPcDEYVMzMoZjYfqcVrKNXOKvjEppKjBZ5B7951n
wbtyJNETOS16DIVDzXWhpjk75Rhcy/N/cLibm6JziEAAkMBelqwxcV+CHuxZVB45
pSvWWrmEr/qUsFkTCk65Hl4x9PLq6YohqE3hTyJY6VJ2qIcoax7TnfdIw08YpW1G
oAt/P44tyxKqdpEmV7nbkIrYXh6ymJPNG+7eKwhYpltKYkT17zb90x9EDmvcinaI
swFq7OdobnQ0bRbaHQCgkzI0R8YctL+r2A/LK7ipwMfHki7VkcAFec6TZlvt+COE
m3T44hPGUPO4zJ1ghy8q0HPX7ehLsYIAsJMReTrAa3uQEIamEmJM6boWbA2ioZCP
Rfn5InpWD4OFcnV9cgUBja2NLEzh0zzT0datL7F4tARVTgLK8jcAbfLPc87ISReQ
Cdj4sdarKYbTZYZxhGH141RnVXIjHuju6UeNYt3u3JZVlhtTL38o9XoWn81NMtd2
sa43nD3YGzuaio7rr8tf6KAdly78el/Ilxr8WDfoAFw/zJGjDJeQsoa35ozsQOSJ
da9NidXwVQmJELlRdSffVAhbnRRera1c/UKvMgA0ORIPVHYB6mH78pFqL7Sa2xpu
zHyp5UUHT0oH9B2pl8VdBPyNxc9/Fh7dNdqwxIgMVVg+e5GK76eYlBCvva/HOo4q
8M4QxetvUpsH/UoQn1qQ9MM+0hc0FxcmPWZNNgjabY8g6AgvP/QtCXMgik61MsvO
9OT/8ySWkOJO2aLKQZnEt5aE7DBa72xrcNKFEFGAxpSO9EZKSE5qeib9B48i8ZHk
hOqbiWuxGbvd9bgzVndzZo28i54VxWvtD0Py1ad3EoftPm+2AmVQ72EketB9IKmh
J7jqAe47lrttHVOB+w39U/PTj8E+IKCxEUPkKcrUReQofTb44clX5qRHZFrT4420
21lz0JS10hFjyZmBMc4wjwY2Q3sTwImSBp3gE2m0AFTGSy0nOdJtF3SMdOrkCbTc
h+7sWxeXhr25hARlXgIfdZ4sQFh4FlX2MuPLkj2vxq1UHhZY/LV4204N4E7iwCKh
vrqGNTsoYKL0mF6lCDnJUzx7GiOJfPY4pPiWEA+0TTaQ4UJB8mavs19jefv3ZYR7
FwEUD3DoxogDNgkkgR4AgcshVQXGQR0EvDxSMWpGtZTIOZiWovSW20+lIwchxdzn
0OVfoNF5F4/Z/xBLaQe0aMyzBx14NqwBdXfvzOfu72ffbkBolNKDePXxoXENxP2c
3W1DqQR1xTLjLlatrSw44gqua27+qa2B+o4yF0a6V8z0RxKYnygNDelekICNbphH
erJyIrAbTYo36ZfP4wF7OsuqT2ypERuFlCvdZHDqSImwDKzwQioyDeitbhz825J6
x8fBbXSgDRcX418k87F612Jk+z0w5rZMS1JAvf2d4veis9qZdCPR4HWNvxaq0Jef
ZBOROJs49Og4KlgNL7psS+sZDV3QTLsAW32Rjce0iugYpe0zZvo/gQoUU7qZBvn5
A3XtS8iuwZfbmz1/+5FOMM5qlWkGhus1kAnYqFA5LGjl55sHo4gBULu04TQ0499J
+5lvKAfl1hwcZedvrB5ZZHwda/WPZ5ZdUDxYvoNVNPJAyFoKmnztnZLYo0vWhcqa
6YpJG9nzKAJ3NOdM0x3bY11RYQ0243ftCjh6Z6A6hnmxxqdszMGA0pLu4qwKQ/6G
IAlMUqc4yFaIGzOG0PNngumUtvUJYJtIZ6QJbK88XelyTeS4sBR5CmC2M+VPXR+w
pJ0kuA4oR84+DX6ZI8T3MW44fdS0aGXKTJQ5NqfpnQsMbQOoDI1RMYGsttq3fJfZ
pu/cXjdqTUL/Qj5L8vhlKldnhf91PqEEAB9gLr/vLYjTYnn2MFhXZrjsiQmCRUqG
df3NFAn+ms6rC8J/ZQjtgLdGqDFVzD8V9KmJ2xLGe7259XwHCLC0xibEgQ4CZLkl
K1kCVRTB7yl1KR7uh7o4FweSd3+CWTB51bT5WTvKYjDQsb4PLAIaLyUWf/Jsfr5/
lnPYRy6azQlLiZ78EV6yEY+W5/9w04H2Nm998zyelNq2yEGwOllPja9fG06AktHh
YmY29L9zz+qIIBI+doBDZPG6keUt+2EtymAQeB9OwfPbvhw9HgySv+JE5+H+TTnn
NAdQmzVADBEAzhGG93u90euVD+k9jFaALjz+KJgZealIn6yqsrNq4HaImw0uWf8V
zXZNpyIaHRCycUramBE+elRYBvAQ9UtNz/00JsmTAnPug2iGz+CItRAMz4w6fL8W
zzWMbp+OWaBdWj3Kmt8zczFVaut7gTvSftCl55/l8N41RsEFDP1GgGIaxDWWFJXk
PpVox8wkSJwk7sXw2xwDxlWn1wuVhTccgaDQ0Kh9Fm4leupcJzXfybSksgVkmRKk
pIqMIG7e88hC+Yqvv61J0lVvo8Gb/6EUU8fvNH0cbknrauUOjYhQrHE0ALDn2LFu
l1pEY+d3W7c/x528qNw2ebjJ+oVtgET6KaeFFQQ29OE6vKnxfgdrErv0+Nyc+zaL
YPVpGYsjB+eQqrT6Ol6XH8jY/OHoOh0NG4bSAv80Vu/QrHIRsJCB3NysKoSeeCFO
ho6q6/lN7C778l9KWthHnuLdYNug4L89rEEa+kOpMNy8NSKeQg0TpTd8cwchBJHA
flVyrEJg9KlSrL7Me/iXFNCGj3N0mKFR0so6I8t3sMaz9C3DjO8DmxJ+wkNM64hz
elTK91YJ2iKEe1M8N6GiChi7IVVObgeEeH5oQot6lqChsAt7VTQbKCEJRpEjfCJ2
YhgCB6KJ3Zkc9TBsVovF5r5aAkYKOIhYUxsltKxo9OhvpOXPAX6xlrC3U6puvyx4
AbPSIgZzaXi0h5RR+gRWmu6aOEDwRC8HpPwAlKDagPyHD8e7cmWqMvmPl+oCr/j9
dU68OFaIOMy4UQOvm6nNHtU7RAc9MvZRcmjmr/yJIyOddas4Pt8OQWhaNRvnur31
z+oG25m3G10jxbtmY2imoh54dj3ujGMfgnHQomfQDwb56XSv6efUKqIw1p1gYuyA
Dvx04jzyW7jZHrsbH0lJEXy32z1VqwyAmrL95CyH5kma2uHIMIKNJCV3paIVSnIp
CrADunACs2w6HcncJYmKvbohpS6BQyLsy0q+AXVhfxpvvINdknXb8gnQOH65+dzP
7HzGGCX7xY1q6cf8PQ+NKnlg8n7O4QQRCLq2py03UXPHUB5oPWu1UE9Slu8jcILu
ZZKi9CZ6VDH2FiiD0nYDFsB9zfDaNRr68TcKS+AufGPv5fcJlkN2ndITZp3kq3kC
74ENBGIg8zvTD1sj3gjJlTLTx2ywzltD1TjMdk8hsSselguoi2s8B9IqGVt+61gc
ePs12ZPLM2a5xq3gOCk8qeo1Hss5/q7mpqdwFlHF4qFseVkFhY+oRJJMtxffBGC+
gIRFQQ9ScW4nTlN1SoKtKA9beULWcYrMaKdU2hqrcbBRjolthj37CXEkw6I9pv5f
5ECAwdAGB5L4oZFuYxKNCP3bvaUklVyR5fmFQ1VvixwoSjai7dhlBxteiX4thjZ/
Eisye1c0vmYwP/P7Q7oR3gUuEjBIXy5+ugQxkRWqmzIgVO+rH2IsYe36+QG9OENe
zJpIsXq6zltCII5waYOGFDRfTzGxcuMSAjGDSnFdcGcuYKJrkG+y1D9kNV5eAivQ
BbM545quvjhndVTXJ2WgNuUU9IouYpCDxq7oYIKzjFivW/INfScTRqaXdSPgVXIe
NwLLMDufvJFxioowbYgQHVNk9vakZPMxkOnKPxklXlM7d1pDECFFSRT6JLZjItXf
COJE22Yb1RrpIgLDdpYeouZTCJm3VuPqVNKQXyTR7IXDa/xPM3lemRQYXoaGEi8E
Va7holhruo6OFmQ06U8kgwf8tSnqvkE7TADcX58WGYfs+d94tXo3c7XqtH+JL1ey
4eiJJ7i4wxUJtD3JSUsCawWCmEjTW1pBHLoZTY4HWi9H6vuMuY2nFH8Y+9ZewMlG
afMw5zO0zxkYTojFhdFX13fdgInmLXuFKjsYBnGHlgrXR+lx9+TcobY65OaFU7/z
ysGhyyFjfyFK+sKOJNGXrqq/pQyCWU/9IbiGVXQgFv0eh/PYYJMD8bKVtwnGJ/Lc
4B9d06OKEC7M19CQ4/8qhs+bqgJMBDgNesmYO60iabApmp7fF7ZYD6LZQB2BcvAU
iMCPNpxbL3Yv2Q7Zh7vm3DW9vZn4JrpP/+viH7Y2/nAcEvN5gtz1tf4qKpFjcvrc
hw0Bv89yq0rwrPFSnH+/DqUX147ZC/AHf/y0fcOZ1Wz/Gw3NHwWccSUmrop1aDgS
dnodxrS68a0K8z2cMtcnrA2ppiHqq9nIvNl8xRD52OOaU5g2jm5hssde6cT7OxwG
kJiFC0hjZsdVyt4QYksfvGVJSSZEJTY+X3OlApt4dpJRrfdeaEoZGQr7ZjS6A2cp
NFMSQuhiwS6gdVmmw8PYP2sucrS0u0NoukOEKCi9M0dMCMXE07RwZoO5yAHzBScy
HvbvOm52Ydbs3DUkvMhYGcRgm+YgZ34UqmiihjRJXh8f95Vt3aQSSIg1bIdsB/AQ
G/zUkuCjk+ubkenZ450xKX1uuBnqS+Js92/PaUMAHV9l+HfUAFqEESWcvWSrnkZT
Wv0XDpAl6p76nUnOGoxw5sD535nZZgDVMN8QNnJGrQh1bSUtYld8TwyjbQYFIw0O
pBZKJDWqYvDlTx/6GAjyny7nPhYIyQul+3c9jAlVhdN2+6EoGcZgAUJtUylI85Bq
PX8agc6AGP2KwB2/L1xsGMXIaqERahiAk5A7im2vML+e0gBm8URNNeTDvl2xFyjU
kqDpW1r49huwzrigg5jtDslzYZwI1vIzqtknspdFf8vMIzhks9FJcx73pxIeSaa6
Mg+EHhnTCD/6D1YzBpyd4YobLaJBiX3ar+bHdw9e+e7+kwUUwD7svVVk8Ka2eHbD
niPca04l0M/ddDkRW1rdo1hD4UXtKJ7lR4btgf2EQgwuxu1bbsGVDu2wgCVHElPD
VBwjQCSZa1QizVHByAzrepKBS/rW/+zVxKGkU7OM+bmmi0vld7ZTe17eA8kbHzK1
Ubxgh2gZO7nLT26OL6rjqn0B7c9VnssLk5XtiSLs5MK7XFa7Zdc1CVcj+22u0nic
MPVtGEWtMlZGVVcQPWSujGDDl+nwN9dJRBgDesJ1TYRmHJia8dzd0W2sZMq0PnM4
A48D7d0Cj6WXAW3xHFYtJ9bOkosvA2ds+imFlFwAPspzUix7vPZbIjL5zstiKFOr
e6wCOobwSoeE/yvyOkh9wrMoZMsTsSU0oGD3seli6s3kxvWFq4q/VUBgkEJ1xKC+
qv+WJ3R5mkHlhxbAfo84RDIMshFxQuhwhLXFbjGwGkRyf56dxAYF43Y4ktb0VyoJ
UwYACzwjSNqSX2OvJLUcTIi1ynVWGcgphnZDRjXkK6lWhWT8K/jMVcxAfR09p8l1
8D8dKdUQMIRaDlVR1AAYQrWunW2iH3O6SPC9NSAZVsynzp4bH1Z0oxWPN+GJR7PG
pT5B1qO2E6qUgpq++um9YKUnXy/RSupjkcVFGbESRmiBpSppIk8TOS7JyVIG/HvE
jCP/v/iUi7RIeEtxdNTvuCZx3qGSaFPXPHSKOZN24wtk//8PrYr8RHpE3+AQQO4U
BY/dNp3gi1XGOyoN58z99paaE+I/AOi7UV+KEWFesQQWx6ltCPFfath694ROAQ0P
40NDmNaa8+RIlaHe/s3bkX9uLbDj4UzqbhC8SSErrJbx+95wjgv646TINot5a1tM
Xsx7qNfL5vg/MaTor8FHaJDwRy+kJ7K5EZZWj8wHcmkxoGMJf3l+V1sLT/1qW0ER
befvXfZKTW2noeGRrwdCB0w5g/FQTBawi78psNFDaiJ0iRt7GkJ+qNYo0ACb3CF9
zcY2+9Vyn3RW360GbsNgJRkKYlDL9An9r2svQndIsWaAEJruokEnXXQ52PilVT+1
NdHQJ6BsN98BujxxNvRLPlvjUZwCxaFOyX8xWquC9zZaGyarBQB2TtnwDHA3zV0k
AMvRTbkcT684NAWA5mbRQkZtsPnkzuP4qRzH+DAnrSjFckq+Vzx9CrUyOXAe4OAK
voEqxvLhWdH7wz52+ItzuQow8J5lAnGnjKGDboZAPpx1pbYtodKoon4bMSvqIVyR
2iKHnyTHgbwFxEZ+AZcN+PnIhgMfX0BSFQws0DKUxBQfyvG6ffBDqPiow+blCgPu
w4fn75JepqZ5JoBeyjkukUfy1wGukWZezDqlUy0aUicJl0jGlZWzrsdKJj23ZAj1
cp/MUjWg1yPg5pTdUH5ZpE2YsBVHMnM1T3GXOx30lxQfCjCk6IHFUaBMafA56FRh
husk1joY+8Lu+APVY57kzKXfTGjfxzCj7HoimAuKZoKcLTtu9innvu//khbTwWS4
ig59Q4rfyFWGYXABd7gKkWqBfR6Lrc/xyZe4FOB2U4sVFZG/D7LEylY5A3dkXYuk
oFGO0dOcBGiu+r63Wf2hB/twqdSCz287OfGNyNjgPWBIawu8fcVMU1GldMqSnO9Y
fvosOx6iz5jHzPhcLDIGx4MhII8sje1EkLR7QC6TYFam3dzoz7n3NMEvq+lNFZ/k
af4yzxoE/Nrlrjr5NzNl7vpgWgxTOKnB4UCFOB6aGe9HU9qxPP2YWEoTWzcw6+QX
9cuRRQq7oJtfN9R4nNnv1Kw6ILpBvk+jPNpBgepKLF2eqbwRhE+kdBCeD6COOAFe
4gBOlwn3gPfyNeVvgZVnOrvANAbudbn4SLBA4v1QoW4uoUnJBSffwxaiQe6aCj9a
79tTFqVpOPMpGi28CuGXlGAEbAa6UCW6qDR/lckK9MXVK4ea2gyLYKFCdspTZDhS
Y3VJ8RWkDrgAiLHUXEObrYOudCnVulaCKq+IlhZaFLB4sRgm3Xeq5Yy+m/hj9ZaF
wFJefRvzlLh7a9TiuQO+Ki37ubeuNe1nOBsYz3VzPR9s1ziWaA7jsKyvV9Zmu2e7
fglx5XnukXLdV+0EL1FgP+NDTOTeOEqBVPruNqfkIYTu2DIo9dcsxGLaPe1AUmJ3
EOKkfv3AGnbyF29MUIvWsW0m+3e6jErCkdvl/9OvLFJd9P3mt6inKo869vq3X5JY
f5BQitYL0koXwJG+Lp5FplqEDSitsdpYjYVESV9k+m27E5IFcbnFbU8rvSWNO1SB
5OtgkFZOtbc4Vn4XN8bI0tbJqb19iCUolskmVtCirH6EOJQEg2B2fkt2oR4+CWJa
X8H1GGii7jXx2M6JphqV04BsztzNc+kdUdLsRRkgS8dx+aeHcjXVmf7THjhODuLa
ADUXngmFfdn5g7NJ/K9SIMpgt9gPnUcYfGrqkl95MN9ldT0oBFHPUhStQjDW+Kd6
grAdtJiv+3Y0B76HEzcQtRgArc6ZiO94cpNs/RipjHablIn+ZMBDura+JigOxqjW
Xc2dHAQy1eTEyQF5vgnIO0DLE7h0xCeannDIoJst6fpiW3gMvSSg0cHrkCMZ+aPf
1lFCikrnFgMwwyLcjz0+kugRle+j+nWr466xuga8NPGRgnxrj1maYri9Ka83hBJQ
nkCdF3ZUSFuHO6oJsDg0p7Zx0a6l8u5xASQ3y/xY8Zua5qtdw6OWeEyjWNeJH/st
/jg0HjMeZ6Eyc32mvw96f4cygENF8Mx1clY/0MVBMjKFRUNoCTwZkqEA5Rl7r/ab
cAo8+TKBUZi+haQGPRcfIxu96Xwb/9scqQFEwQfa7k0peh/k1+bBmuL6gjrAwQuZ
9SANCrl+EegrnQATTrI3FpW4W1pY5Q5ZqBtcSjXGdRSgwH0oheoEyxw+WWqId8mS
3vPGMovPEmT6LczK8ZibS1Zj9470rU8auKbuih3TzdaCZ5a2Hwk+EMul0/Cqdst3
oBWp+10xf9j3/6AvG9XtgYI/QMr0XyhljnXdN3CXGu1lfd2cb/L/zU435su5T8bh
njkVpEbiQX5OZosqSmLUjA/8QKIHXKVQuy9Kx+H+uZOjuhnPG5hMacpS4WM1AU5+
NMyKywDu4+mZxQp1aeN0uL5w9rXdtWlZKUFKQexbEe+2Y2q1lIRiMRPe31/+Cywx
btUWOtn6igXHrw02fpxsUwb2QO3DOe5aX1dchYFoIaJTqowUleQDzZn0YWNLdtBT
v5UXr2nzYpo7l7wm6B27iL5mEyx8OfC3Nhx3RK/wcjSwxrAITMeNU2lhDVYW5CyZ
qO1STQ+ubJGd+j4SPfJf+fZHua2iIT+GlwfY/6TBksiHMOIODL8IgMY5+38qnkWN
Y7CMBCc9NhyZo2z4JZbhc1IUpQNxuFlvYmpQ1hANPR9rHousqrlMSf6F0DnHWfXw
AKlOs2tQN4aVrxfSI4t9I13t43LyrxnVSu4UwnS4KyLhdJmJqjIvD5Ajs39AiHik
jl/s0dAejeJDJKI1ze+zi9+eUlPdIrwBGhMiTHKV5mDsjSfkqtf/WWVSvEYvdUED
oxEarOEyjuUp1neYhGvOFS4kq44hh9LW6fB/yBLoZiDslstuXNhOUqmPcUGtJjUf
B6wRD0cHhx4iXEElAnZsPZ9OuaRII6XXmo6j/mQFQd5D9nbOfn9K8mlFiaUqKUZ8
96Cx9NDxwbEcG6bSP1c0sNXhuM7Ebojo0cy8ZQbLnjAEH+gEPOuKdVKYyIrDnRWm
FcPIkOsTtpAZm1+EBjZrWIYkTeCTum0e678/1VteoD+CpF3r7nH3jCr7XFh+2MBs
MCMKcZTLEMy7iwhtw4jmcRL/GJMTv9E2c5IlvGtJ4ViZV6YoMmhsz67t8nzIOUqR
eSyN1rGmUTn5xAtSsvhzOCob+JGNdeJSduTGYWa3lXnEZPrf1m+swI9Cf9QLcpgr
dOqfElxMbcDLTqy6oRUzPOdd15UlOBBIE3oX/x80pMLdXFyIEm3KNCyyq+6PsZ3n
PQ85V+N1udVlKF2rAxqa0NX7aB4yhnNabFKUXI5RkdfRuS+hZdM3p3QGMqFOf4v3
EbNi+o7w4TUpaR/dr7eZAfKT5oUp1tfWcV1uWl/YkNucq3hqcM+PhytwS/zDpc/9
whx/f5B0Z+Vphujl8rvW4ip5W1Sy5DZ8//SGA19wlRV1TAmiw9i+P9LcpO+oo2DJ
pUQ5uqlG5xY3WTzox5mDiEwJSzrVHACJm7WBgtv/cEHem6BBP6LY45FJhJ/9qZgW
rgNE95Efbz3GHYefhEqHvsQz0drxzBphnwI3Vj5/I+ha4gEVXyX5KqcA+qnRlY2k
+eB0TER4rFR0/+QnZkNV8uFOBpyykABUThJrcTTBRyWesyP+sqIQHEzeFa+IQFLh
ztfTRQHfhvQxSQaIlQNWfCLKDbfXTshaUhw58sGi3aMN1OMrkAXrcCW9pLhv0Ig/
5JOhyq8mW4VtBFD67NIAEEaJfYv1hAKQWdv89lO44KANmizm1KI1M9EeDDec6ZqV
r5eow/gQf6n4TwPgpemGf7ybyaQbpLLRxpQGiioOffOxC5oReJwBuBrW87LscZvW
bSGFmiQ7sHM8VPqQzdB+Wwtqoo2HYJiVqYbDFE57SNZ/jMOXPBDk8atAvGtwBi0B
hMBpnsiFJ7l+Ay4Q65kSGpBKf1DW5fUTxliLGFYZPF9F1+6ZZdUSEP3dOyrzKpnu
Wc/SqTr3LqEffchf7YCphW37cO25UfO6K5o7ZBOv60CNyfmco/OQVr9BBGVYOz0z
xGs+WiWpv8mP2x0C7uhlyEzLT8AHLSx3QZ6eJaFj2/bDL3tbvKAsk38YmkimhJ18
TsONMwjGN7qkyhNQ7xOT+PkhWCV3v9EUmlge9p0RUCUB5Cerm9+qCK6/q8RgmpCD
lcGjtzBXqhOpoZm/bqTY7ySRfuDGjpdWx9Qkk2Vcv4TPioADOVRKajfQhH5qfnhK
PZjULbC/cCzQ9DEqx7WBfIgxAiEWxzEbABc2fgAA0g4tEe1dyvP+9B1hMc0mZB2w
cyHL+zfgaZSRU7R7axNZM2L2AMdAbuav5Ve8RQsemUF50GFUmgT/rbAN55ngez9j
mCqHHo+C52UZJNM8C4LQjP0TF80odCI35BjaZjI6mN05PhvD1GjmVN85tL0QTaUl
s2qQ8nluKvvjc34iz6AEa8miAGTxSReUvjOzoO/tOzgCLlce4bN5b3sFI2v4caq4
PBXlCDxUWiLpEc9zTxg7GcZVfg0op4qGVb61KyIuUi4Ygpg5HHxVSnTKbD9mE/1O
GaOWevZDllLIjTnq52aHzFlDEmd0BTfymSMpuAe/li5M6Ut7LLKSir1cpxEP7lO4
utqcxI3wfCvAy8IbZqx9oGJU/dWivApZQ64+rKF/oA2CvXQfuOq55Qg9GEHbSmEa
jN6xBU1xOcXSOW7921lQSo0c9WFSbEaN11AYQxg99BsYew/I7cAo9E5Lh4KINVnR
srO+xXaYVoBr6Jw37qYsYaYTNGrC3gLLOuK/KQjGSZeagQmd3OEmSaC2cjzc62nt
ok3wIL0RxD/NJ/M6OzOTVp+HsXGR7lGx1+m74qalBwJTH6Xqgn5bOxixMM575SfK
dB4mvrMl1O5Ri94HQYnZmWY+xEQcEcRM5CYhWBG8uhAXKrYNq8B7DRLIeo6gAXqv
A0sO6uNKsIKs6/NgHKIxtjLyQ9N+959WI/MTOMVL66bC7CT59LEnB0O9lxHt4krt
X676CnVicSxI4VhaXTfsIHQ2ElN2/ePz2nhu1/Js4lXyMM/3dUlkcQ7VSjbKVJgR
rEc3yhyGzyBtreCoUGynEsyxTGx0ZfE7FtFSLNSOXvlYLBgS1cEsEofbaCwC3OUR
fEBpdW4bhObpRBpQXdsmnPt018+vUWtLYpyFcVBr9obK8EqGbdET/QINjJWNaNdC
KbEthuje1a4o/iU9RJAfnlWcsE/lrJyxX3S8gXNmH8cFncWnoa0MB5Z3YAPGhFK6
4QWoXtwbgb/+0My8paNqDom9KzQoLX9Uo1NYMUgTXYnRyG8u9ZRSAWJy3taLu60v
+roYRKKfZsHxoU+55L1yjoj5Us2deslnBedvZEMR2x6nxditBpZauOEeZ6Z8dZoT
H9gLgxbHHeTfuzzbRdP+m/HpEs1/FvtQCJaVRsbARXtrkDAlAm97C/STE7hUDHqi
La0IArOdKxoum5DOc+FuHi4Tj+RdP6P7VQKT+tbTNTbYyCR+086gOBqcU0csy9aC
1L6wqal7EylF1lRottPoTHWPQiuQBxNlR1p+A/TMK9sLGI4+7s7/V2wrCQ9KyoFU
PsXvl9a8w+uiu9rV52tPHySbVWX508l5UMFccpPJf4svyUXisGtu8qasukpSp3a1
38LBGde56wpFt/P3Qrp4hl/wn2ZsLCov/2IKCPrI6boKPSY0VZYs50lYDtkZhhS2
buTCjwQbXjsrRsznSveaagPj7CH7y5adDUobe4yne3GPsGny+bBs1TpXhvM9XuCs
hF3AlNh4kNiyTBoSu3jDZ+Lf6B0rgkAFH1Mvlp6R8YpMtAFksYRaPiDgi5Hy5INy
Vcqo6phCLk93yCSdEPmKrEhwEV8x8IEbq91G8I/o1UukNLVNW3O9S9odRPnQ6skV
wmHQHItICTp7MO+getB5K/pIgIwL4MHXKAoAHdMN4GBbeQy96WBXqfTrS9tZR/gA
Cdh25Iv0nP6fe2GiC/FQW005ExkjQHgkwgqAXw/VJX6uVAguPdt/pgdLniKWxwH1
KsMIU/nDBQZeh+nfXHJFsgKGNASe4rln0e6wlKUmeJBp05WjQ5oMOXdbdd8u06KT
aL35fjL7khAixmOd24JoUbbfmabsJveWAsPRX7eeT3NODuCWN6olX12RaHGUeFPI
YvypVonI8lg5YJBBsjiyRK4bND6lyiSl9XjR36exZIhYejvZVZ0qTfjsyvuiKKPE
9Mw3ZqZJvVudmMMM9HEZFDkU0O/DO+dYyiVW7a36HWfGrS0ok7GDqk8DdRDE8hBQ
AX0JYOr2hprPUpAkFq+MWDCvyA6TxRKSbz1/+CzlT1Fg7hehC77dVAa5tgu8A16y
nTXFxhiCyaQS2X/PWNqBAwQi9KqQAT2pHuFRpgoZCXJQpMKFkoTuStkr7pDeKohS
Gn2SZN6P3p1JB9sdEGEU9hJWzZKTqrI4FpltdcKWlKTG4HN5tA166pQKtkuO06mc
oNB9303nCsQnzG6bR6+eWSk8AzvSTd0utf203vJ0vU2pomYnuCUcSyx/YqCX0ctx
4O9CChANiMW554kQIa01wzrn7Nxjja6I+I6L8xbyajMsijm5opCT3Ft4RPSD/mph
40i70sRmCmH5YTwh2i2heS1EaYdJtH9Zt5IAYjnXaeGijV1Y/Cuuj41wR0Fklvih
4ggTCsd6Ju32YC27K44mohOvnWrhinPSBq91lzT0da1t/2twPrcyAhYs9j3yb5lw
1DhsHzOA9FFLpuaaIc2P8aSII58QJgCk1B3uQta5UasW3tmJatmXHb0JFHpIme/A
PG+p6nlu86v3VQ/Gz7avgjrH+Ef/cvB3MU7vR40w124g1zFqWeuxxu1erTpij8pm
Leeh5BaNQjyZDdVR5t9+Omp8h2VtGAYk+5ceblNE+fE7Oqy3p9zd96LNN1Ol+49P
8IBU0FdfTxq4xBfWelspEcVX348/aWlK64oDkDIr7BB0+7nH1pxN74LJwtQEdar3
zuVjKCwM4PSMWFOEU9dwXmewKuS5ucRQdWG3vcwMcPfQ45mIi9+X6x0cFk/BVNM+
VP+1r/CL1NXibwpr0XZeyVjwGT+fj4y+mZRAT0XVqTgIhlAv20XnuTf/YaZWRKF9
rY79fQlWPecx9Q0aiKxbwF8uiHfg5aZuRbHt91BVK9rJkECICadLxkWDDREAzu2a
M1/EvOwYCefaR+vJyKjbP8ILgNPiupyN0xx2WWsFfYPjQkBpY7SOrYuIpCTEBV6w
xDq/E2WWIzWg4DZdpGVIg04EAEm9BMmZLyn+IhVXnRGaBsBPtXP/+u8FS5dJQd4F
9MHnT41r6YePWRp27ikh2ogFzlCixwFBQMsQYQUIsAx+0AtUQHDBen6F37ux5SJU
NugKDlRlql5xH19axRFP0/x+I0BEdG61xU7Q2Ii1UF8DW37xJwbaQvMCchDsf1vm
PSBWp1VPdfoejQGCk1BIB+04w9ngl9bgvPsj8ocqD5Dns6Arb3uDwVTkBGbY9N10
jtU/MZKHpENYabom7XFuZeMTRA5u4VnJnWsRuQ9HYv4qjlV11H7RwF4lDZp+n2Zg
DJxuz9wQdZHNLrFnh7hOvNdLA0Tiob6dN5FLBPhxRJfdiH52whAH/9UIC0rdI9na
nk8B6Isj6vFztTjpokMPoEAhEMfg1FMWA9ci9RyVt7mcHt6kdknxMD4Hv5+D7cYZ
PYKd9lOuBQfm+hC1QPjLOvrNj/03sxQ2m/SEGWLX1x5LOwHOEOXksVpdKsf7YqUJ
ifL5JAyy13NdcA3tr3OR1VtTyO90PqxkYReODiIuL6HUY3VEOgW5AaSgG+175xNx
dFwLYPoSkiOvP7A2c2IRw6rGnI9e6S3m/Eba+l5W6xQxldVjV7NvwAykRy3GfPs/
nclI4v8G3eBM3nkYkzM6rrsF5ggVhoSG+xVQxOXYO+v+r+PL4jLpgtwSS1UE8jJI
3QQi7nWvbuAyP/1gGTpWmmUlHaq/i54hHjccYiss2VMpPcEJ+efiAz320MUomrQ4
RzMe6l4wm+kNPLmfXNgqQbIVjJB2g92h8CypzuMyD95FyuBEG9wdp24WKjP+4cSZ
4o1f5svtLGPjG8PU2tIndEZWbhyAMAic48nDSawvXxY5J3Ud04qCalBOClZOkbIj
DkVgGnvLvP8XsKUf+vEmz8PsBAHlYMj9r72htCG7rHXh2hT8QXkdrr7J6r9Lxhsd
ex2Uo2e9+Etq7GVlgWJHTcERQB2WDlXaYf+xp15uym1/VV5lww4SLqe86jHQURJn
e9v9+HGRQsveS54NWCJJdUGoXiNHE0o/aarUt+SdleYVBT3tjzD7YfgAKPAtLFsE
Mfo0cCEGn1hKiNGLT6+MpGx8HbDsjoXsMovk2avs00LPbVEyuXMIdNpJjiOB+tX4
YVPiy7Armf1Kj4T/dBcGXqPNrpEta//l8aew1AX9peLB8kHkJDBvrz+2xXBjb0qS
YOogsbPjM7mJvbxznQH06Ecb/DBw1WsSn9V3+F9tE1Z26c5wSSTejG3WlKQf4Vx9
cRLpVJwoAkOteLYZ2ja0Jdzf2+yGaTG7Nt2/gFBQxbjzZXh17ljO+vUY59TYyile
olw/WSLXRrB9Um9Kwtw8tmpJLSb/o5kuzzErHtiUPrzF0Dk1U0XaKHM0zs2BNHgZ
Z4qcHbuGTgpx3Eu+BUya0n8VQI8HsfJzH8OKt4S7vIJM9ga3dHgueFv4lKFNdR9J
nzaVIC38lrkDvMJGIRh7W1PvnAd9byOD+qiF/NmNhVQg+c1/7CMVw1RmW1WYGBcW
aG2cIkLmAXisWTtdaSiq/w3Nlc7dpT76eetucKb3t3wNKskBhu2N8HlB43wG6XSL
IA0Z6U6Bv+MKVDrR+D/CcjtcwMRltLOwF6XSjqonHnfJ/h0U1X4AftjNDsLKnQGN
5Xos7WZMjjyHXR88zgrlZnv+qKJuYreA7jcVhFJkt7T3U95uTJtGpOsoraDoMjxF
JBWiJUPqN/4L+FECaGGpkXQ2TBgkfzmSNhqxzVNWITzjnu+2Eojcv4h2FVXHgRrq
PCdo3y8VwNiQ0mt/AVdXDWo/DLxVv9KO6uAV7jVkAJDTwIVwUmSPLA/htu5amlsR
cyXaz/121UQ7hssh/0pJuBlDHOylXBGYjO7965wfL4Yl+46zrHnrrQUSonbrm5vK
VeGhzzW2yn4CuGK0K5BTWp+S5SXVjqjYmE9NJZ0zqPuRmCUTdi/zXPjF3BZZHKrr
Vr0O3l3vFRJSF4aGjenjpOenwzJ3nDaIB60dZ0uAuO6/CT+zd/tL1vxiupnd8cbj
g2i8PZwuykHdKfwNW+i8BE1ZKhCivvvI+Xp4cFYlQ8nsn/Ho6B+QvOF//ljAAk+2
rga5YaF+uBRcxA13Hf1/7v+pkYUM3ChG7xmwZmq5Ewxunt9Rq2RlVY7adtOYve70
n32e+xybVyJRWo1LjCsUE/iAGo/6Z3Dtk8NS565INSVuFRUrYXwqAunRZkWkXwhS
VNWLd8+6UvHDznyUoBNB82b2lWRReiENZY6+C1Is/QQEtkDyqpm8LD/02kuSLOiU
53Q6pZqH/X3RG6mfgypvJwUNHDJC8tFsBGVuEqrWkCA=
`protect end_protected