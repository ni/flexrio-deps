`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36768 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
YKazAXTwZvVeXonKKI9l+3QOkipZlw3tZCyICtnlQnFKHqHT9NBj/QJwb7FuQTRT
sm6oS2iP8BqNE1WzrHuhKA5mdqBCxhBD8p4wqNvMXfOb5YQJ8P6gIq3YxZjVVntL
g12B2izlHnA5as9/gUUFebmwNRdf82Nrg3aPKKFCODgCIQ+ycR85sUyPOvMoT7C6
HnlJPB+HZDM1sXbSd0/wmGJl68RuHUu275irjECTMILiFOJml0a2K7l2gzzotQu5
ZDtrWqd9k5vLy3l3159kL8EO67qENenI++jfZxPLvXoUBCSHT/INyvySx0RNz/05
EO0zp/z1EF/V0jRJrBhJcNKJOWHVeWGgModQbHnjeZ04y4/TLdMbLE+5zL8eadI4
E1DgPNZQr0N5xdErBboQJyeUm5/KA1cZE0VzhKIhA/Fj8xDHq3cNvkHdD2++WvoT
gAao0SBeDb0mKVfSQiW5NVxNYKe/22YVba0/aYi9TPym2t6niv/JTJuxtUF94brM
cjotkSprEBYmidWvKTWnhC0RxcsHhxDq69zNWkGYxF8QzApymXC7V7jqD+/f472T
u7Ur4U2MHr1Unzm1Gp+fQsVzlhj8nUGRTwmXvlB7J3bHwfcsOTbwiGA4yPbDX+B4
S3EsPMh206gSE0RxYDBJ+wqQy4kQQqkqiiepxs/HAlgIXjZygR8M4xaHPQ/9koau
J6PQ+fAuNw0nQYjirysTSqAWGI0ISCvRpPKc13TYX3+EEIp0DOYPmkVUA+7/pUk0
upS95GRGGf7sKl7X63On+MRTAYkbLDNixMTIo7eY+pkwDhUCV4qOm5TLqQ2umozU
bu+GU8OLKTN0FagZR3BUX/Vl2YPfoICFgXalNEroW33UKIJI5OoGg4bm8Wkd67l3
5CE6QaDotHbPoTNYH+RJHIcePDNipIHXY06VRoQG8W/s7rhAWL+wjMcmPWVHUJD6
y36l0gRqGE2ImNIQ26anp9mfUwY1kAAnt1uVUsigyhziqKFDxCEyoSexX89FeUhV
Cp3lL0+lVBVApy0Vhps0Z8XRvav7Ab+ZXowYlvkiUO82zWfO4wQODzChQwk1htCm
uaK+4hc4Es5sM4DemVu2SKrQ2uH3aKniooKZDeBxXl7FkKoov3EBJKGUFDlJFbMy
8UfD83mS+renv5E/+4nPRvDqnpDEU7rMnpG8cI6Zewse6GKEQfKcsj8CqeOqUsJX
0YXRiPQhStwKlXde26rAmi1RftqUQGTT9+auaphegUf3n0tvJYKXgtSsM2yl4LlP
QyX5bDeFsnrXM2h/7NHCWAXpnm22tTsyFQycoEEgVOhhSQ6bnxc8KY9vD7U2D5sS
l5hUO4zgM7ALalJhi3ZOoQ6sBVAzmCbAMEgHCIm/FAZ71KBs4v0UHd94BodhJrZz
38P8ureD8Qck/qfhoLdLKmZeUqFX/LEaPCZPOVj4q4San0Ob8Aa7xXMMmMbCJlrM
dXjnYGfEFK4hOSkVV4Ql/WJPofzl3NN06HwuouneVLBL4twwmPHAgr9fygeYo+y7
uqmYEP2NhZ0Z6JnGOll/LJlGOjxVsg3RvcAHUqSUfm/7xKXaGvAac4XlJ5bPulqt
zL/7ZqY9yDxSqnQ3PtBphTYT57jweeSv4Uteb3sxn8jgUrYb2odqkYJFXLRIuM9n
JOGpQcPp1SRyTVmerdPCndFzr68SVrle0/Puk+4DohFXcmiIhBdnkCu8sMFCni6d
cRrvavndjAQyl8UqZM5F6lltT2QJAx6LWOjZT5sJCuhEAXLstb6Dm0MMNPogbAbr
Sp3/0Y4FyESVQi2U8KszCHpqh56C9H+jrndqTBvk7WA2m/tLVHEt+/nYXT4STuAK
jKtX7z5hWnbs2lq/BEQ+ChIlW1LAhrM3xuAb///vUHdtYvo82JzNQbC8ZN44BIc3
YkennaLXzzB7XW+NLW+cWd/n3PeSGC1DfXfv82z9bcDmTIr4CnUagkrG9LeBQraT
d8KD//c3IPMrC8S+YSLaocxmb9+CEVcbycLgJx3QEglDSniEdmBVZhXWhEK8+S1I
PxfZgh9MLKCowMa+/chu47XzS5OJA90qS+olgdGzYlTjgZN+JlIubQBb+Zxu5Xa8
3LAKjURda17pcDO7kabNGo21q0e2uh1syzJZCTmXNMk/282O7TUgQIrVnRg+n93T
TpfIoIFhr14L+/ppfIw7Dv4ZLFH3pERSzx5P7NA0eBqxPmZ5UIDebHYWiVm8S2Id
JY1GNdNWTGl1HDMq+yq18otDwO7GRGxRsAQ6EB+dd5i2tVEYXJujPL321RY8bhKk
SLYj4RB4qiwMOLXlOvgNnXrZ2r5hbbvxoDQlxd80epMWqJyFsdLq5Wl++Wv5wxfc
ITKd+4KvwHF3VL3rXruHrT4ap2EhiTUBLuhZ58kkymnZGnUHMUVs0Uc9XTcj7grq
rXPTE2N+9VSXGtkLIq3BqVDVyYsoX49wXoMHojUSeBaGYyVGNDH0xAuPJENiL++O
Esa/xzqxCoz1XKApXue/SGCaPLJqrPK5hBcb7ZbGjyqxYM5pzGCZkvIBFJTnKqDF
q8p0SUIkya6AUQnKzvFo4c8LeqeY68QNteGDtgIR4hA5XPxTxW0Ei9BdVAwdpQVp
ooMplvLtn9sDEmqWjzkf9ucvQ4Ijtznx3aZhF5Uzm7bsv5EfXTTDhAK/man/B6tp
CZLVUIr5Mwk4IBoHGBBo+lCcsBAnWjrAJDtlh0u2cd8FtIdH8MsEW3KrnkeUx/xV
rP3rGhhM0bCLwg83gaGDTyZWym7YTA6kIlQv7cq8VtaomDSLrgtwPG+0ZCAfrVEO
8PE/NCMZGw923CoZuQlaJ4aI1g3CiIZ1xUIfkB5S3dtVZMWic3GIC5VF/rFaZsMQ
Ls2YwtevLgD8T1h8sMGX9fh8ucA3KKvPiNcTYCZ6U9KpRnoYZG6/ccXLUk/0JGhN
AG+WDEH3Nljowg0DVIExA2aPNrhHoE3/OXNZHaE86/1oOsnplh81bCPSpkRGc0eX
f0v9QwQ+OG3Xrd4aY+JeNdaTYQJJvOcdYN5I8kKj62KgnWQPI3pOOSrmUEAJZKnO
SO2dDNRxNuW62+vSmcULHoDIK8QnWT139aNubf02DgTXe3ITD+vwB9q3z/n/sPjS
ZaL0gP4nzej8Mitu+OxPzib5VfIorSaIuNpZdbF+EMSsulz0MKmvaMajeXkQ1tZB
LIBnchATYAHrbUZIOmumam9Pv+DG+uFcKJPF6ho139DcsmuRuoJpLK+tXPIydlIu
7r43DQxTcLoZ+W6IbO8z76K1guDh2EXoastc4qbVmivkQo1DUKkbkJUfcbevWdaG
fW9mG4ctxluhhV86We3FeoPozI4u0W6zXZOBlVPuG5NhQ6jD6IF7tmZjPb3iAuR/
k0iLXX9vHR2ljraGs0my+r3masUI7vHTY7qASW6udUN/oDIyHgq0bkABHtVegGlV
DJSJhUfnukc7UT6hgBG2lZmj7vdLtcdF7h5MyoSHhyU45uRtJG3qiFdDZ1NWly27
0OIPeBlvza8/lz+9IbUoMo/2B6j276alCzXWnGlS08G/0dAlvsiq2+z2H3BfxpjW
ZiMvMY6kjbesY6DUwtSenE5gtF8TxqB4Dmk4fWl17lj38dgcFmGWE6TRu1YZdU2b
XYs5FX1kBm5IGbKAWS7QKrkOyyOCCU+Sw/Eb6TGrHEoceGR7mhKyWDcZ5OtgRSGi
HmngiZqtr0l3sIwIVI7/HEltc4RvnZ7Q8kOp+scX8le2goZ1u2dkqs0FLy3QLnQF
HbgvQu/zCndaR8biEHNEPT2dk5LrhctaSz+XDeL7lk8o+leGdMWN9f64KS+oqWnU
plPmKjuLh6NW7PXNTp4t452bqoUvH8WTHqRyQMCcl8BMoXKW+ov6CEwl5MnYQPX2
XEmBFgzJc01FkyesG9AFoGBDQPaNY1/GJFtjKWBi08eSluCxnEVXaAZoptL4W0AU
RkJ95HjwrUf+snndhfFHIzPX7j1EZLiLpFNb6fQCywEw03z/pRAfafwElrsPMSKB
x5BD15S0lh5pKheAC9GVFmwPO+9xEXk4l0avOJhU/uZogNXGc5q6gQWstri7n0tj
ek3MwAlOx/AeELa9v1Xe09mX7fVXgIvnGPIZ374+1r0u9aQUfbpg8lYNf+wuuZAM
SHft0MTeJW9nAZpd/z4W/y+0X2FyWw2hpEyYwEHQPE7MMOudaPFcfW1O1xyXtgaV
MoSEr5X1WjkAeDDfGpLOVVFZ4230vEzN5wBDq053ICmtjKjyitHBCbR3rhxPTdMn
bF3RfYORWWixcP2En10g2hoIoj47t0yztp3XT6pepd752/eVmSsUVk8BhhYPTgYz
VW7423FoQe4DiFXSf2/9j4LJVnq4pyf8qLZtb7dOaPavOLLfqMlkvyrxDwU2y1Xj
LvvtNFlwd9/FZeN7MNE/WYRlg1foLt09BW8WobFtBv4zh6B5iXEvYlobbvHQxMQ7
KrBaB4SFjnXiY8Cqjg47FOQu3pJcRMMljtX608AVqBmF5OCKKoljOthRoqpq8JZu
Jx1kyyTBo6wl0zLlrLINvKf0mu+9SP9MiW+OzGeLqZusEEZHKAA5SI4akgQmEYiA
ZWKoqQ9+OeHuPHtt/knevwjwNnj9pi4llxymJoDKpvhR/hlYWdnY9fw3xw70t0ij
dV2lGn1R1poDIRuqoQY9Yuak7dCpLvViiD1WHA6+T9cwlkTgxvaxhq3XOPzr6cmS
DR1y3dy83XTv/VslMdSt0kpgDoiqbMk8UPBvwC0H6+WJ+4n3D3xWGi32qgyrEsT8
ML54P6sjIEdUvjIJCoceds/fzS/J4eShlydHOkO2zsOEMV5FqSchuzXcjpqR/hp+
Z4ADmG0VduC4yoEGMIfE0IjSpynhUk/KBmCi+sZdSUkyik+lZA8cGn+5+hm9BLib
Krf7YCsaZ5LMe6ULeIxX46mZceGxdnaOcErSZ+6hYW0n3wvzhiPfg98Ur2V8HNH+
3UgDXjJJ0/1cV5yY7+IeiE43GpkOd6Sc/FG9RATiuD7zSEDJHSoWw8j56MZeXFcJ
JQFchenMTTG83mGSQoe1hN2nXzKYvckDwTM6IpOl9FObMjdiace7CPE8r2z3d55h
juLongZAnpMeIuSenFWH3MBLArqCBJXSiUnGP150mN9x7gbf4jAWE9d5hYF32ZTK
L8B0Rf9xKZxpdvddihMABpgKltz1FaX2ZcfYPCM8AYvmwa9UOvFcR8Wv8vv1kUb6
+OKnafl74XsmrMneLXnmESAuRxxlkihmRvIlRrpfwamJQoSY21835aF+Xa+di64o
7zEbKS1yGdPzIaRO2CdDezn9oJazK2TccTtMX8JioilANzkXcTe//Z07ml8wl5nw
IxST7GT5OTbuYiJmv36AwKmB37GdcLC9RBVqJM1RU6c7347KBQHJ9nRp83NJdgam
vMlY2RYZ3uGngmjAVQmJsfYx9UM6EQIOoit0aWfNkJGqkjzzvZZfDUDb+Jzb9Nru
5ri2K/gg/AytVB77PCn+V+YKzrN2UsERzCTtw0QCg9a/V+XjR6wz0A/eH8hTuCzS
BPdQ/Z8z4RlRAbDvWX+WIgZtH9hsqpLQg0rB/4TgfZrgqH+RyKRXnHioI/pBY8Or
lXg4eC95Sazx/MTcniJsPjlbvZSfnbHq8TylbsV55TBHb3CBusaScllJWoV4oJWO
likgah+RkmsSbJ7DELgOYiAgEKRVSWiPsGiBrolfvYX4upAhSxYlcz8kQEl3o/Qn
0JD2XyM+ApXgBlY/JS4Pw9kuobXT0LtKwZLrcPn5lS/bfO93/Y1IpvcgDGIqJfN6
yOuMQESBbll/gVw00bWThKB5BvxP1OZ5Ij1hVZcxqBYkzfVCvw3h9VWi2mLLr2qY
oxMcNYFPcEOaYT8QqaQeeTdnER4OV5t63hGWdb0pztexU2ALXWnRzRQJDuyaMyPv
WesG6xckDDzCAsr0pF/TY/c1y7KoajAjWZBBQVFV1muClLJOUzWn3XC9Ct3TVas8
PW9cWmoig1EWY+zw8mIV0V7ICbw6EJDxtcWiSRjlOQhQZ8vuluw4pMB0dfHi7kHZ
DiAqZxyhPqXwPhzW0a899CNsjdiwAbv0+cuH4pFhUQD5cWtoIJNUSGFzPdLfMhrk
3VA148BVOclIJZ/iDQfe8dcJH2/lSUhLtFnaOhCVWr9t7YiSTDiCW2pEtoC8fKCD
U5jHHPG2iO4i8/YmZMF0XLxYsjKDk6UNNnFr7b/TmnDAWE286d21vk6/6k6/5rWn
8AJTEfUZmvQv4xV2VZ0WhEz8DkpWyJ9lgmVTUY5z4n02Nyflza4nc6k/e/drxTzr
UdQBfGZ5/uTpY2RNsCC76qgBpp6QXBSvYUan8YSPBb/d2tdJGYV/1QDMxhYXgAaK
Pxmos030nVUgMg0Ch3YwrIx41B8JugNqWk8AzmlATfXoWwBMD3+lAFFnNRMoHZ6a
eDOFdZkEvwLcjmNr2v7hTbVEMOcsBkairu+Bun8+Pa7KEX0HhVBDOK/YDUEBUWZm
54Gn8rPv/T2xeXBirmrxOShi40SLjVBVsd0KYGAvcy4raSaXNncz+L8vMnBYnA1U
uilQGwH8CpEiZQbfnSjY4wefGegqpbV7MwnyGokKJewxgi8OekExM8IMXqG6TCkf
Ovr3fskgFMyHBNPtkl0iT8r7MBApSvmw+RHXIZQf4DnhCdhBcQicz9BechK70QJJ
aSf/ZbYriiAFHK+T8rQWnPcSD0uUpCXU7Yy39fYQp+4qM0Pzbd9f0Hgj0bIJhf8u
DdeyWoL4FWr4Cdj0R9+NnvL1C8BXQQaPAOMVxOHsP+3ba8TOX1nuc5yVbH0ELbuS
0W6nwXtwNnzrP71gUHVifax/csgZCTQ4d8SuNTBM4vsGEqmM22W7W3r41/gfisAO
8yzFB+LrJTS8I51ZY96OxfzhPgs/HS3Momhh+YCjA167CgJpaExhtNgUTFy8tfuq
aWJV0NnfHSl+5Ck1C7GoROwyOKeORUpZVEo2DL8RZYcfsCKWaMMmPeLDHCG73BuW
YKpNtf3ifLFGNY8nEEKcxIbHs4wTDjWAM/9x+QXXYhqTzEznFYaOsqgO7tkHu781
PPDKzwSkkB9NxjfceSQF4NZyiUzZMtNq39l+SlngZBEqpwOP9iKSkXbJvGRqdD83
10cK/cI1/JOA85gzpBfFW9pagxnm7EEJCi4jpXCjIb+mgP1I9wvewT3NONdzFyao
4/qyiKNPhnozGHjcSIBBILz41feRT320IeaJFRs0L1Nqd1f0f5AljX15u/0ZIMsf
+guHkt60Vw2MiKqPsYwC56C89yGsj4rbBBDnTESdw0/JSbfGBjvmbBAaGc7JxTl6
cwsx0L+26jAtPEoLLggDlTabaFswbQK2ESEl5uuVBtk+2j5+16FK4X0HepNATMON
16/dzBHl7YvKkw2FfByJiIO9AK/TXVZ2u28RhwpOhM5p5STFt3sm+q4pgJ48XfYg
7aGzsp9rR9paP92SNoI+PPcBJ0uT6FxRqifXHCwqZfn1Bz7kcy2Fi8iauh9Lahlr
vxstSlupYKn22C244dnMS3EBfCiLgws4rHyIiuTMSE+5w+jEjT/93dW4CjYzms30
58sdKPqZFqemNRGMiCyxlFpGr2sWCCQlvxzWakywvOoY0JCwZtCHnYlhBzS9LENf
SHSg+5nibP9KkSPtqrrgb4rW4xPMxiBvCEBGPVSx8WfYYnZyWud2JsEnMKYqkcb1
SEVNAdf6Nc5TmtyFa2lX9ncP7F22TDL2vC7nc6dY6WUBNbD276LUL6u8STYFk8Mz
4r7WJgi4dbLh71Dqv3/mR+3hU9eeI9p9EYKhJtvtBgHpJ73ihcFduMjPk1YdNY8e
L8PHXo5VYendRq2wojOrnsqA1elHPvZEqB5LRXakW0MXRiEeYW1rGhCgXjYfwBBD
h2DzgTjSbL0mTnjnj1oYykbPkYvyiM9TlmOT9c5BBoLH4lfs0Ol+IwJb4zB5r7fP
C5JdhYhHlajZBgonlU6XNP1+dtyWesaI4sTUfqa4b0qGbYKrk6Ke8Wa3Ms6MMK/r
q8V0uNdMBQzyR2gTrZRRpn4xSKjIUFtvkT3tGfEBLt0Mm8NidHYdmPEO847JoZkt
Tzj5sj0kY4EIkG1KQFjrhUZRuIHqfqnf8PZWbKFRRCr4kQKq+4fBjB+MHfyJb4aD
CHWKxvf0z+/lXoTSNlfsUjKdJtYDaaF0Ii0BHf2EUfnAA/BEMYKLNevuoQg8K0LY
C9LBgdPL/8qRPXN2jl+xa+6t2Uyvmh1G3jgPEK4iKcOuofUpUwO1lk6Z9pxpfo/4
Z4yYq2sBcnZVI5L8mUhrsNl6WDR+piA58LU19Vf6kpOsDkWSEx+i9OlAJIKnM+3Q
mQHJFmtsubzx5fgGTNkxA+FAdqD391SjALW09BvwYBxiGuL+0YWs/HIAo4SEitUb
LYXyIZg7ccfrlIwH0zx2h+Fp0TJKdOZ5xgo6un+6trpZ7v79y9qIa96YjkSsIQNj
iZndzkkGDrN6tYCtAGdWCroIUlelRIP+PUgZsGDmm9unKamFKHH5vn5Wvh+ZAdwg
kKKfK1XkvKey1AI/qTqp0gNn8i7dHRL5vmp35pbdn+QDQt7UeLoeaE80jMBijO5P
6nUq7b6/tffNJms53Oh8p+dTsKtA8zMkr39tc3X9/6ssqCpQYK+sgiQWtB8bZFhk
3KIglpistP8ExMmOsENy9ZqvaFTGBd73ciklQsGEEQeDsuZXY8U+AHYDEcuo24vR
cN5vr8ebIvPSMTSuABKBFTKo69RBn61QTz0gYbK6O7TlQUzTpyIweegfDH2CbwjL
5mnHShcSjyForPVFqFXEsynTNyW5wMWAmv6xFdxGR1z9sdhQwVg1USE7l5i3gOTe
nVwKS72GYb4/dc0zAPGrayFIcVWFfH5l8XQVuuzUF6dleLjR9IWB2DA9Ci+esK9+
iTw0QF/R9MUTyPWoIfD1NKV7VY9mn25sqYvxyIjVvDG17oBHcNJbDou0YzfhwbzN
d0uRCQ+Hl3ZEeSZW/bZkx22vNLfIjkH5GpZRenvlkRewejGB9gsfSfzigc0tyAUX
st+N4fEdtvj2a09gwFY+b9953QNhZcWF+dPdND76ZtdXSQ89yW9UM+WxcO7yM5aY
DphlyqYBhFqAc9RiOLdVPDfn3oqNwgHfEcfW3NOzw494Ha6Y4Df/tzbFRXT8KBDs
hN9Kr29JbOvlVotxRONSu60Xnck0AIpBXmIQD375MUsdSrCFMDyxSqa/YEhl65RU
dJzPSJf/pIhwCat2NYHejbfxMfv9Q87iDyGwuAZVJOfxhTB957kFIJYAB4t8ysrf
rWUzQ5ubuvwgtXhyZVvB9G8rn+qVRqznU7LNB9n1OVSd2IezGQpp75tStbQ25hEP
xH4pezTp2JqgTSOEgyAcHAONEF+oHo4a+AP4upBPMiO9xTNiwx+zcRmX1S14Aovt
waWO98DwiY109M6qQiMIyWPX2QPH8jL4An0qAA+aFQC4YUJALn0TPuNKL/Ah2pFG
6r/d1ya5kTXtEyKObnaeCDssk9KkA/8JnL0blHccFL/1V7Qj747MO2+0oRIgixkb
1mGIIEhbZLWtKkSdO/tNQ/YdVCFb575tavrmwLz2s8NwHUn/ge5OzN50pBIpEgVS
EnwCRvy9h+cAk1/7vTrUsbwUfyi1lKUl82PAl/Xo3M2dxckzPM7SVVAh/hcmjaA1
oBg5WkGrYuc/uRgwM6yeXVq+T4mlV7yP3J7hBBmDsWa4Q192hlfBf3G9HJ0rawuJ
28400NHKJW+fmUfKwq9EdMSnB6c9WBzn5KBCtMsJvtVf70CO/h/XyX8o1wOx5dPb
pNYH0TIiS/o0VJztGacR01kGCnA++1TKMkfWCr4l/KHmUTEsRNTkIaZY1aq5YR43
sqTSQnKVX+3rRaVubXRnP4YaUYILMdJIKCOYGaOhrs9EX8i2tf5087jm27GtAo7c
CfDRAoR8GaZCTU5Pf8tf1MnmY8gnQrHhfQngxOvYBWpACJYG7nB57ZiaxUAKN98K
ez33TnGY5hafEPbXVsDhZEReYsqjehFbKXGS9Kj34LJwYT/qPrblrIj+dWAS4gp/
GDXgZcrq/2bdrQpxbSFTeD5Evkcsnm5abPPM0e4uiDp96aS1KPfRzWXVNt4H3tAm
2jhTQ5HLmUXX3ipdG5zQeGnezBDYLkph0wchFkZ9bEu824G1azISuffFSp8yE4rG
3osl0ldiURpx7lnJXcawiuIDFbbQx0Smg2UiK2VIA4oMPNFTy94nZFOJF/hyuEeh
lc6xjf8OZfuiVDM8ahAKtsu5otRKh+kyyi4yM8u6e+08rIue0QI2SxBJyGPKkiqk
rmrfZE4RjVY1SIsA3FZBnlP0IsQ+PXMzptat8ueL9K4D6QCOQo8Aabp4NnDcJSv0
oLMJE3h3GugAmKm/8o8FNNzaMeIfTv/c9QK96mzWvZpQRriVsS1tUzzKKAHnIkBR
lEeZcvaL5L1sBknfbPSwC75vSZ4BXylkDOuSJsepgq12kCUW4m70dGfUhQHeOw2r
cn2QFr65tiyqtDUnByyVsZxqEJeq8FwhgUysJDNLzaB4ASy281BaI5mr7fJJxJOg
WqqsuUsZFF1H6R42LTIXUxOqU3PHid3wYsUwcrMJKRiTZdFcpaalklEQBJ+SFPds
AmoL7A1wBirYXfjlxcT/icnRewouqTw0FqUCzRayFLJj7d+fe2BTJ3aszfiXdsXb
nzoyuBe2ND0SNQ2yXcQZJUjhDfXZ/HVWrmpfPwpxIGNt+kv1ozpfXJlI4SL2SvOk
vv3TXtS3odo9ZB8j8nONuEXs/JnqKPpGTKyCQflL8BAPfFqc0EqBhIEiBGIglyZV
J/7+rctFQAGjiUrqWm10aN3Y9ADxABJKH8/tlPrXIwVaM1qk4It0vM/N/5dAnhLv
DTZcIwjw3MKLpVRuQinAU0SxsjIj3735XrdkNLM9W78/Bst/D5JqN/mVZQAZyj9Q
KDrV4yx84cTRHxTnYA/G05u+tURlavsuAbRWuCC0bIhbI9rSLi7V8BofB1Fubehx
Hyz99WmNowsFbOfvEnlr0C0Nj1k0/UkxjmBawgjt6H7KlLvYBcYodVI/gufuBy77
GQVVmp/39rxhe5nOrpNvqQwEgVggwEbXnNiCDSPc4mWGgbA/rle04cjeHx/RDpqy
vQZDmaqiXj0z0tPZ05pwVw3+eYRgvsqzzpTUyCMbAGnY58XLxz8goSikKTAdJqRX
LPBazFVEWi7+2PM0Jllq+5sAJLiAx8jMEj/bhZ2e557tb2mhRenxYFXzPEHMrRlk
bdpFcEInZ1Is2QHWVBMlq9lOozctQG7IWcdHka9/7xx05Vd8MHUuX41P2o1nZvSl
S/Sri0AElwogjO4R2XqceFFBqNNSTz25Xj0ZMCDPL36dD34JE2tvAfYZf1tgS9ZA
vVgET+FBxvMnyD5EkRs7l+v7zqkOmI19jh3muX1yONB7etw6n7CSI2Z8XyVsHGlY
Lr16axNdCrKjBTkHjE6G8aTRwGd2g9C+86+4aERb8zoBjRNoaKeOWm+7KImcbtdg
a+Xp5fdOkQlY4n1dTwczFLaIt2YXN7wcLOjEUNNky5uDeNTxVAdfxJIgCwrVHCsi
3Q7qDudWMcI9ngNqyfzBUytlT9s0qT8RklBqYLN8+BhRduOvAfQ07KjpGfqQMLQ7
Q909JNnahHmhPYwUWR7q4IDPLXjnTU/cKfozooS3tHQtFnjRk+GBKepc6wzf9t16
z7WdFaX80FYxQb8YSTMTJGpRTuXjC6+1Gqzel5VLBu/DpuQRj27M6JQVEsVV8/ud
br0ZuLWZmKRdHrbvivnFMHx2sN/1En0x0BIhWgTnl83xnE7pT064uz3A0wgLsxme
AvD9FmAgUaRWekke7jeLAjUdCv07hvkbCaNCqk4m0WUFsWdYKqck2+xfgwzjCuIU
RbstsXURQnYa33ZjnzYPNvdHYSuRhhYo8EM3KD1QfBZuaMwpwP6jn0izLxc9x1og
7nftwVaoNn49QCiNBNcZxlTH5jQ9/bkuYlYPQ+BQHOXd4sX9hytZ3xxC6cH0JOGS
ChTEjQo7mzlPIpdF6F6lRMxmaVRVf+PzE8AyF45Grr4hCMxFM7CqjWeH7MKNFgV8
eEUerlpBLmmBIvwiAH+ja3Ax4fep7JTazxWSq4GBffqp9YfiwpMubJPNfTyxK2En
5lpFSkApf+yKF8DKDBr3ai9RSEgL/1w4IvTyYcOxwou1sGLOEfKCrhPqNOiSY204
HoynSdw0ezcyzwoi6IyuCtUwobRJ8kiXn9BbfTvjZy4nbbFXE0PPgM6dA055A6XG
cvlqInM85XHAKybwLewz4Mowqlh5psKKlLMAW2UaGGoNk+fF2mQLImQdafl34V0Q
13j9jK62KpD1QV+DfYNpgHOgtN+5F0F47aBxmP6iHA2WymI0yQu0rfu/6huDPoTt
bLfGObgwRlCCfcjZXuWM5u+gzVfNHhkLxZARfPTjxX8lFM8HqhlRnH2bYDUuBHlj
AkrxPYKBAiI3mOjwPz2NpP7XZC77+b0d47WT/DyECOzef5q8onq1ZUbQzFrhRmXQ
khmE6UtoyGVYFtlECYCXlbuP+4KdO7Nn6mOXHf75zuUbA00srXkIKeThlCO4x/cy
4B2ywUmXiV4t88I/Lg+E8mAhZU8hsH0350/M1XfUiTrTgpcpuJOeIULoiedCRyj2
+UcwCxKSVKOXvkM4mjnMgRxbA01AirPsj8ZnjJjQR+vMN2/P4ito7n3A2mjI+3ye
XhZwREjeWHdN3LL9jB6p+UH8zKrXkYySb2L6+c2Aar0Xq+dChZklHc/4N5zMSEGG
qgr16BaM51sgRfgGHnTNcRIc3hLmUGfoJ8F3oEWb3i6T1BBI9uQEzUDwLkK1RTsv
YEJ5O0mFQ7OkwBt8SI7Hg6idgHUq7G4EEz11ruNwKGLZcj/9mN5F9l/jmG9xOItr
EC3nvdXXlImTGjlWj0G2krN/Xb5XgE5gZIVommOihMOIkmcGEQd57hU+65uRn38L
4tqWQgGuwsJMnUVGqookLTu+JsmEPX40I9i01fjNUWj5TCJnxYWP/qsPlG+b2sX8
YNRlQyeZBDpuSvXRMVPYbXnX/C+AsfyUD2KQvCv42vSx/M3iyTb4INIP14u7S6Ss
hkKLjynoUVEGZyhyLjVdX/+9kKpfGdu9mXGVzcm04nMja5x3mEOOvbM6kOSlCP52
zDfFgzx2W9Z1FODHwHmQuwnR4L7qcAcgW3MWqlmrb1fnYZKWpYNB1lLmeyt72MKS
WG5kLW8yr19iM789y/L4QSpRf+U3Tvtba78fIoI8NVN8qEWG11zjJRZBbdjdNxPS
VbBHlANF5woNADAQUKcmCc1k3UaaPLvMbZxQNDmldB608uN2E26U7aeDvijNdsjW
ItNZrpwL9KBehZHWfoJ4uW5FosusgDqwcSD2imicQHv/AcHn+exL8i7A54FOGXHu
x7yj6wIbT/1fTDh2ivkunKSD88MRS83A+liysjd2BPmw6zjs8YiY6Pz4/5lMbCkX
SFeDlokIVfGXpnFXazspGT2t0oUfQRU1zUR2ZCPo6puJgHmg6bNOJk8+QwUId2sZ
Kh5ORuHxvXM4Xrxr0HDnHDVAqAucacvEgrDF6aW5Et2XGpzuWZykNTXhGIdZ9+tM
kBwoE6Ly43YWiX8K68GuARZ3/VbLKSsTdv/VbmYiwBMWvC44XF7iorCkDBW+4amJ
+jFZ0QUu8PyCuIEGWjALUQZVIhLrtZrN9cuUmtBmhYaR6p1RQdEmO0SVF8/MlaY7
PMDkg4EfwKa43CCt7zEvp7ZyJaRPZDEuEG/bZf7YvW+Yo655hBvRFa7DzDTe9uPV
2fOpAjNlJ4+ZcOZR6uAei6qNSFzYag7EHo7hMzjWtX77jjl74EFdgoniyiERp2Qb
gDiLlaxlRljYYmF/ycb9777wwNOU0w4nWt1Taa8epuntodNbRWO1n/HxzSNSKDze
2Rji2zKMOK93MQZzEzRr3G8mVBvccAMn2BnhTIjhKRq3FSuzO8d9h0e83pBN1suI
CFXtZWvO/HpGpX5IWRaGKkUdl+6m/Wo44jZ4HLSpo1SFk11OHaPSOhgxpraXZ1Sm
y9VzgMkLTMNcdhiZEwDcnYwrcNq4Frxw/8Rs8MmK2vkZEq5rBQ+P29VXQezZaEsX
IVmRBDrSlY+o5MMaQybN0/8Sa5PHF82bu6QYxZwZGNHMtk4p1qlUh+0UrBLxBTV0
mLtHY5WiqqE7TwYm1p41lGN5ctLPYVQuFqMNppEwvZK8rjhbxGRV/K7RfTl4f/LP
eyXwjpQ1gzylpu/mPDDoVi4Ysyeh36Tt0deAn4Dm2pZOh+iiXYsyxviELOD+7zL6
Y4Cm5eVopX02vM4Owy96vvbT5q4opEXkZ8wGEJi46OYKs1fKLK2ckkphkgc8DRCg
kNyRy85xA8EzCcDiNz5RiVk/vlFzZ8D4zdpg6/svjq5DPEOxD/XiIUxM6jqtruUm
POd7N3pQRQoM6kOJaB9VXvgh0PudjvbntH04KzfvHWTdgEiQHtsva0eJdbTWYxnh
QoaCvpG6TVDqys/mlOgTIrCOcxVU/VcwJd9P/syvVEcN/+q/ynpN/QSQKxaUBZLi
v+CMcUsyGsmt6h/E6LDoFTWCLyvsj/HDkGvssb6pmopYSAQGPr4lQ/amJoMDSLBA
Wjk5hz6tplBOxSJe1kk50tE6tVe3tXRDOtvkQ/v7/VdeAyC/Z0edeX17mvVXbOKM
QnPxflYVgxGRg95gPoOwV1ty2sgvHpz93hEXHGiPKE556l/BE6S220BjRRdWLZ7N
mY0ANwHbnOlw/aMdSX5ZDpuAAPmomEh2RfzPwQtjHML0De8vo1YoJaafgTOl6nIa
OJMhXDPqJKwpIoggyk0kSXn2BF7FC/BiYSkHk0Q1JbXjoiynuKIr9v8JFvwDJyOv
ZXYdShlAdmz6OINyIvyKU5F+GNFanqT5J42I9Jfp/TG/FbXRIaB8Px7g5jTVNW92
CPrS6GBf1KxjOm7Ss3ulu1ezXKkDqUtambt2pPrt5upj7/Vuo1e0+fbbJWpoh9n2
RhKNMp6ws7KEx+SFXgEJpnuTdmZksyDRxuVY2umvBqPVNzmosMRUt66Lz/vVsDM7
Cb8S6T1dNtjqSRlwf5ET/3wuXTKM6XlixP8meMT7FznRkm6uqStlEZIdoC9E+gV6
3LxaZpuqeBZtAqbGSbP+9SdtQOccyen7EjwXuFRMFiI1JMsH5yYQ9uGbaVsRgM5U
cEESdrVtJD5sZPiFh3dN9mZwV5W60DavEtnyh0w4U87tL4xl76o2MKlpT5NVroVQ
TAsj+cC10KTJRJ7yF01RDqGOZdVpUgibFW7Gh/w0GwV5jCjrpAOUFKVKzRcAmNo7
B/aEAk7tF5JEW8TYKRUK/N2goOZ8oSv4sXwPxX/9mt+eQgvuqaa5ZA+w3dMXZIKK
mqcXrklJEQOA1r7W62Rk70J4hqUqJUCfp7XzHcgJGhUPc1sTl3ZOHs7dbgn6R1gJ
dqV8gWqz26YCni2t7djSSBA1eMfrYFBtIGGrmcopNND6037pDcHtNhB5pRNYg2IO
gDbO/kcwcCQSPQJIwdFyG0PEoBwD1AfYswF9EyI2bDE6j9uZFhlKNLpYLlaYnew3
5HZAWoorDlwlFFU8XYd8GNhFqUd5jrEKvz4I1r2klK8YH6W2dbHsa85s0GK7dXc0
Ucjck1Hmp3e971C4yv63Sq/oF4xEFdEaG6T+JMgysepGRUYTzpZ2Vjk8VxiBEzIr
19W6C3Y0EfQ3U3cadx9NrsWhcBucSjl6NA6Ds6E+PbhghzulrXAhsUN6IqTjgV2s
z3HaS9gvAJvXvA0odVFqUs6NITYaAufjk8fETbVP530Awi8oa9hMWmRkRAvKzjHp
UTk4O/3lwNMKpMnnNHuDroCw31FYg/yprv23lUIUuFqkHgOCXNhEY7g6hc2ufz3q
eZO/taGpzchOjnx5X7ljpKhpjHgBfxMj6dBoc87Qzhkx5lViVJs5ivm0WSajR/w4
IEMjm1n1TBSlTHWhp7vyK6HtiOx5qxEl4mo4ae5rYOzOG7RFnoMClxRpexjDH9n4
6yy0gRjp5AxOXziQ2cWRD7+yo7i3hTZcvGj2BcTaeGgZjS7+VJ2sFBUW7p4AiKeh
82uUmEIlLydKX8TFcuxmte8p5j9RSskbd3bfcr+iDIyvn5FX8/5zHM3HVX8S8kpV
Tn5hB1DXmk+kJOh1p1nGcsL1QpJoqMNjqPtLIbHHWhOwppzWF5W34y6OpyijJ6rL
2MHUUZtPvJ+DCpjS8nnDZvlyjKxRVVDgXANWd9hW2z1M6ltNrnzIzm/6nWXK+a/R
m0ynk8UZ4rAeYWo1/AfiSExK7jCQqyI7aEc9dUAAg6gal6TQBQS6elFsrCAj1JzP
V3E5S8OWtMOJ6glWDzkYU/aHkmkrwcRj75FwFT2B35EYcuxDswOcCUGntL43fzsw
OfaPOnZECOEpAmUQJP42Y14Ofnrb7P/fH3SRPKQaUqqvjTzoQVibA3/M/wIw/nrn
GxJTY+6EvF+K3eadf8BJBC5mvJhKu/9OOu5S/VjnB5XtBxmiM5kDJIUQYTdmMnYm
GCEPJk5FFnuyF3fie90fMd/V3/Gmr2pzoCPye18BDnL1x1cmUIziL4Qz/ztG/Xdn
9lko6+4GMEYaM/EacryST5LfYpipJQuPgJufOIeu19/ap82A8GVzxIZy713oGXxX
HOe1RougFk1xHEUXhp7sbm0qGgEhqaAFpaDNky17RtVt54f4EpOyfWaYpsfXxlCb
JIGQ/2Ak6hmPY9Ug3PrkaSEVoyBKBIhB5mZGPwIoGgaRTHF72QdMhXnphBJlInEo
Z7MsooG9zPsRI7XVoUURcSC0dyYbAlMVxXI/iCyb9K/Ua1ns+I1aSZAJh/xrkxvR
/I0ad077emjF6TnV5g104/gTn5gCQdklRjoq+TRjDBh6WGrxvKRXENFxve1iRo4y
DIe13ZNcAThAU/nArQD5bVuOurZIdVr5y7SEHtBMh6udjH9XZZ8TsUjW8JjotHNH
gDl0WQ4EEwAnRvPiDC/rjp0zl7bUQAw+ePG5BrqecMZySAfe+5gz+sJrrlVE2ETV
SWymMWnEu2/OIviuh+yLWs5BMbubVbIE5Ib7Hv9v3fKjnM/Ho0uHuQnHoO3Rkxop
G9axk3sAOWySLn8Rt5Ip0FR9sufErQTIGWxpPR5vtu7OGm9xj618hGoBkCLED2oZ
orqHC+SCv82yRwx9pTj+gqltjyewF7rC5G/QjeAsqbzX7ZnLT8uZgtsgY1M5/JeU
D3btZfMXKzbZT+41Xw7kpy3m7STL+m/75JZ/RenBvhQhb4dLur5AjgF433Tnr2Im
kLjfaR5fDUi3gfNlYupvA2eXO6hRIr7yJD06W6bMQc0+WNEuLkF6oVnGQ5/ds3gM
rR27e583YRyaZ2XrLpmgQKKzMXQMoDP9uHwuB7M4EGZroK7lyHS31AsX4KcCzLw1
U9wRhuQQ2V2SXTZDl+ehOg+A4bFT63YaCHyayLG6XdU1FDRGpjEjYxJ9N7/MJI6/
IsibKeFb9rdI+aRPf0QDODJNwRgtiHfkF2/+2tXjJhPGh8U79LtTdP6uzzYk8hZZ
tfUHiRrlw6wMOu5bYvrxKua24xfCawyvYDWMQfLDPMWr+zhhDyRqwLnMK+Qfbex5
4aAu/STJs1Smf/9M2XqFXPI3SBrL2ZHn2X+uMQJYue56DyO44fxh1jdI45MEwukM
RtyA48BY4b2wSC/KWJ8V9ofKz3tDyOEoz8NoMqIweMj2LD8FO/hTWLbVxrcxT18b
xpss0Gqa1DaDoiRNqd/8xHe8mRgLO+MbMQZvmXSt2uXtL/M7XY22GInpaj8UoV0o
FpHPnN8/m8JpzurtqVGYpfBvYfAI29zuUg9N0KxBL1UrCAFfTTlpv0lzF5iSZux7
s+GDOb250JELj5gA+8mB7dM8BGTW9IxLUL96bAoF+mxIixgiF4FDTRbWe/hDg2Mv
o+Z3oZmcr7SASs0tkNb87Vw5X9imnutcL8urLl1yXxRNixSUe5C63GTRlTxhW9mD
YFnXqZ7JekO6dH7EpXpdXXDsSSRWICpox/oU/ghWESv9D9KKhT/Wio43cuhvmh9m
6/zxgj5ZRgBFNOhREKL/oSZ/ffEAvNmOJ3y9sekrXM/cnE70TYBEQ2+ZQS8VkOzu
F6bOiiuhMGt+c60yQHZ0LyqMEfpcOPJPhbd9kW8bACBBhemh0fpD013Cxs2C8UQJ
CDZDhRtj/6ctdO1iR0sQxNV242xB3CAUCZoA2egXADPKGIvt+f+xmRdysmqgKrQ7
+Mcgu9M2eJuuSqGY+kawLk9MkBMV0cNMPU1ILeplsPKOovqvIn0KK0BYcJQYYSgk
5b61ORZoZXvdkLO2lqlXPQY6oEun3nfCUPQn0ncOknEen7rDFiFP6Gff5hX3oD7E
6tJg0p50qeJJ7bTr6vSN7F+E5hgkD7z2aQCYrwSNHkS8jhVxNJOinJybtIz36nnI
AGg7pqN33fKV13NUlEocEdA9VXIVoYZMzkTcz3NfcSBVxSkiQiWeIZ7qkZxIKUAo
zwgeIXmpSh+2Mrzu6mggmZd3b7Bi3xJKl3t3pWKM8RzAn/Xev45BrX8GWMCKv/Eo
MmnDkq4mH5ofGQMO1LXnXddMz8/csI/ExHKUZW6v1Kfj4VYYGqkuEF0a6rIwtYXi
0o0qwgaMPBcls9vEfEuMcuqDMSiqNYtm3zh0k7i/JXW5rbzre3SE2m5t8b/cG7Yx
eEgHbTu4IHNNa9gthQHS23sxEmfrm/U5lLwZUGXC/+85YF6GuwOcNZtSBbI5pYW4
PYKOsmIhiZbbwRTEESrPRmc9Lc+0hrVqqQSauGfJqhpkZ5XEFwdEhDv4NYZ7gNd3
vPPKn8hz4ot3KvL+rdQXrrvNTrIW57oOOca2aWQf1VXrrXtKaeU1IFQCdlgEVn2U
k+6y3OsKmR/YhuHz9xObGcWFrBZuYAyYowojtTcTpAOulQ0cyzvoyA5QAn97wnSC
c1MHZw7k1GfJz278DUe50yfLR73sbZu+H4uiUV+k9IewQ0o19fyGLEAHS4V0qwSE
Du5BfsgTYQ5l5rnlrwC5vh88IrWxzxtJF0FDLpx1SfM3TJbDwRXKIx8Zja1Uul2l
lwu6lRpbjdISGwjhGo4ZyC0HWn4wQBxIdopFXdhEqMHhbjR1nwaZkXIZFKUSEsI7
Ef0OLM3axOGFuWqqgooEsjs3ykgnBwap8Skn0dF9y0ocJHrJ0X6BNdd17HfK+x7i
JH/v3P5siXzOP9rQclGI9CRIl2a3xlahi5QDN3Km9efuFzGP5JoqeHY5Jw9WsRYf
BRdpVx68KT0CLFyTXXNIa3Yvak3joyG6lR+7SIq38NJEh8a+mfITi2FvPxVIche+
NlrDhWJXXBYRlx89x9VPJOqksNF0OlWLgkPC+QQbs71APyLGJFDuGM5RM6R3JLhi
7QXZ0yEIG+JLCd5PHwN0oWPmW12QF5NsHVy9GdOq/L33CyE/7SKSstpec6A9nFqw
ucMNkWVc7wf9w065YzIfBtF/Zznj9ZU8vbDyuAnxz6tRbTgdGMTOyHEVvtJCqUBj
UJa16hmtrWxwp8woYzw5zUnItnylM2TCoCuXWhiyXfXMPgq1vgdjA5dXMrrNEZ48
qdMWA/r5HrO1nI64lf3QAP4n/76u90m1iYMBwmgHclthhFGhjll4zP+Xj2c7QDRw
p/agn8xBoI0ElTi4JKypri+ckdPWmDhevC5zbXNTRQkDs0Ptwd14J5NsazV+w+g5
9YkrDAwyF53FrzEvY0HYmnjKD/u7L6n7crw0f3eMSkOXVfUZrGZ7X9710si9JLzH
jjyP1HtNbyXC3iC5prp+dlesTPR0JD8ZLn+vqFg5hQXrivvgHYLqwqnMzPnMEBXp
pFJHm5Kr3FvCjJJg/ire/62AKstGEzt7uZIcsHtqUb30DOxp7BHj7E9hCRc3f5FJ
RPtKmuyLGj3XzYOW9TZBs881QBGUubLC2qWWvq3GjCgNV+84s02AoWHHxE597w3k
peLR0xngZ1WGGgJ2YdSxkguURyVxYBXFG0FEnu3zOvvx/bKmS+WwDRgZdGhfMBJd
BDSrHGH+5WVhleizptZbQ4lj0w3WJ6YKyi9raOx6AhRFVkxhLu8XTf+aHzv2FEgR
EKuBXRNd+qy0qc4R9nSKxxt9D0h+WW751swNTtMywTGqcag8egxH6Y+SKOng5YlB
V2wEBwnIFcwn3AHfK4VThgSLc/2vJKV0lqiTiCsvFEvGcZ4X0XWzQizATxGyZ+vW
OdbKIL1xhzRwyxLOTYBVVHi0Lk15F7asNW8sZSCgKQck/1Je3TOSRMr+B++YPbmQ
HE/g9dhjiC8D20pdV2F8OBTppx0FitTFoTchJv6mAwev1bpaPIEQ4BQ/2If369ox
DzAQ78XmfgpVOll+3qUJK6R/MklGLMiv3EOzLfNpmquWDXWTQsSd5ilPCQ1480oB
q8nSn7FeQqQipdy7s+eJHzo9/sLu89spghQUjVf8PvTBpG3OTB/oKzNDovoUAWAl
UAkvQYj+Ui+k517L5OAlNzad3IBSbnWuLRp0pY749fm7ksJz4JO678ZDSAzyUAB0
H/Ww2ZMtCst4i4B/PNp/MQX+6VBlJTpfVlmJAll5Wub3ldyjm+iX/1l0tR6JwPo7
wBsvplh4pT8IeKFHVJuHUpWkLkYuD7Ux6f/fNlHNkQEuss2AInLWNJWZwF+RIOKm
rfaj6TeJ8paIZwOQ9jNXxVRYpaldsBtxKDZVYWz497agucIk0KVRlJFqUd8Vde53
SD9/7yuBNC8KZjABSxTVl27+oKPtqk7wLDCWETKFcDjdpvL2ZCftsXhJqcu7nKKS
g9BiT/7ecnRbuKYkFWxj26m2yrNPvWJlFKyvwkOxU5S82sn0nXTZ68SvwqpS6UdD
6Ldr+R40nAL8gX7oDsxPZ3c+GsavuAaygilXTBTVDXARHW+0Qv4GfZoZ/mIuFjtI
qeUs0V8YWtHiuPStmGYiMvACN/qabRXQ4twDbxnBFhCI57EUn99T3AvrNCKXV61E
7TS5yPipHN0NzbO9IYOdATO7ldmxSZ0phWFwShJr4TwpYPxoNF/asEIFjdaIk0my
BAPtzIguNnIMoqk+B21po104aAx2NjuwJ5oXaYDJaEiebPvrEFMggz9WduXbrne+
0Nbl/mTnURLPPLLP0rgBc+GTGS42r12P0eXaTPkjDKmc7I4ZraDlk0v68SVzVCfE
LFy3PPnHhy73NiSOUP6iQjbfhQ1KwXDA/HRZTXZPU2QuGhzQpRE9Eb7IJKx4vn2I
vsYqQgLi/XBhtOT5wdSevo6laxXtO+rSEInNvanDgoqGwHxd+QMa6lzREFvjmAwC
lRbyK4BQjH9C85Ic+aXklP4YsH3NwOpjEi9Okz1Kv5KE0UngljmJ/Oj20nornDrP
ae+33vkGmRHRutLjhmSwqlXMVYccEqA7o1JkGEJQdk1aaXxxdFh4XJqUAFdBDMbJ
IWwkxOne32+SuzloF4c1M+RIpOxOBUmd2SUeX65CPAsxgOsF3zbyLBjEM1T7TYLl
I5w7Vhm1PeTTt7u61Giu3XgyNxSN3wTawXMoBP+zuC95IwW7ViQETBbdmHv6pqey
kEtDCCX4//t2DMEfEwAcDY+sMaL09eCXXYjaxW/rFFXL9Q7rRm36+MpI8xJU+g7j
NnXIWaXwLs70VqxgXzQCypWRkLsHozIibjxAtMGd8KVTg+TNj1NWXuil3olz8+Z7
WAzASfddmWTP2tiZQbbuYkbvEvugK23qKlZh28qUm/AZMwUzsDATLUYZio3yjcKR
bpHh8M6gHQhiUuJigiMt1SpRPrgzRJPzd9YBaGtk7CsI74OyRVTMmrjLBQH1LDeV
2Mm8SA1aWbTrVy6TCKhgIu0oUpZSTb0F9pS5OXW6YNhkmk+LUk9+8FMFGtsxWsj6
X3HKxVGLG20vK0Z0X7xmENg5yGNI9eh/Hf+F+kGgvg2hO/ONvdcRy3UEQHi1NdO/
I692t7EE9iy4AjI69P23eytPbZH6mgbKckDI8ZagfVau80oLhNmdYcJhgNHDj5VZ
4MTDcf8gSKMJ9o4OSucq+YEuNdJutT3xRpXDLO1aQMgcn+ZFMY1C00VzS2rqqdgQ
WcrfNZR02H6UF/n1VA9SSpdMS5FaF3NkQB/txuJuMzja3QZUqK6T+oF6NuVn81dq
S6z9QZmQErVhInB6Rd7+ox4+Gi3CfsvTZQtB23y42SYo1stWz9m1FRzHPfWgoWy6
OI+2M+Kf794JD74/OS0l4Ul3CJb2NieS4FSOVgqfI9KFKncCT9l7C4qDzhOEM/Ui
AUQMQsl2A6u981Q6VcVKbqBwtffDnC6XOZDdpQ1t8x2POan9fxkLwLofjGCVfh68
p1W32qZ4RMCIM4XlZ/BEE9e+8P8kgDRPF0/Ol2O8PeXTOnQjPQ7hEwgAjOU1TYKi
8xaOX8mhU6P9Da3yqAUGWKTBtyQvTiLDkCdtB8KCBUqgCzGftLUnQhUbtGMw2uPJ
t/zZJ6ajwYrgrsEY6iRNGkMWVM0p+wH2OU96rop+EOkNzr9Bw9VcdhAUui4IChKk
B6oVL4A3N7MyWd0wV33lXA88L2fhb14DMkSL+isnMVSHDZdK2362P3qRallAxJzW
tTSiZ7W8izqLqDZ44jtdN4ULVyLTK6XJnvJpq121kqMg3ZtMqebGx/lFjUrVjgvK
IAmhsZvxe62dMWBUE5CB2SCLNujrqr8QKwYNc2kBk6VaMEQT6IHOjbieMYjhCMPg
/pIBEryQGW+nLVAmT9gbbn3/FxyubE3dsKsmjaFLYbdskCnYc+NGxrNJXUCfVtZ0
UQuOH6IQCVEe9m7Hf1YhheRG7XuDpp68FuvDlvcZwWSvUXq3Y6l3WouvF0Yr3a0U
QuS7Dta50hJ40okEP+oXOY56wRBvQ951K7d1+WPdfMQBJxh3vcl8MwKwY2DKJ8vq
d5Sc2hCq40LZi5de7i3/yYekL1gYDbN72YbFeCxlDU5TwJfAWZSnUC24JU8o9iAL
O2ZsHXFweTCpQBrqhCzSVYqtJM+fOofiBN3pzoSVHoJsjQJKJAIoKyaEauP08Z4N
YKEqITiet5G+sxpgAaReDwvvZEhTiHrqzgfReyLEbFW8KIFgMfhSXLj3MiANdYGk
HJ4cXgrHOEfO4665dWGUP9cxn1ib404msSSr1i1cvcRJ8tEAQzslN7rwqGDTBNkB
s8g039oGatXajDaT5gIoU/NUVSFxpu6LIW8wSqaDah0rPfmUVjx5EMumPHZX/YCw
57PT69Y+28MWCpe+xiRij453WYD8sENhVP0qKhgEkZMoBkuEmf5bBHAyANL3DXez
frT60O8H3fBrPjvO/QAk0um97F9a+P1VWLEN6LLIfY7Ppg4hAmkfo16BBIJ62l8q
l2akd59M3WLueYOgUbXzg3CIV/bL3Wy0HRM3fsYG7eQgue9xPsw8cAlcpK85CBpS
wBKI8mf0L+tPtkWCx4wJSsROUl7k4lYEJydd/OmWQBltkcK3aqi+KZJA56YhbYhV
AVJvAfwzB/g6FmJ1+2R0YKljc3tNL5gJo99PMzx2ts5+9j0njNHzbQW561gWnO0q
ZiWQhmlQ6TPaszfWsbzdW3GXeFZbHfNjxz/0DLq+PFueYaea/up5myET5cx/s0FC
4QAoImlBhCYSAdUnC2fpbwO1QQFUmXywKENwwTFFC8yaD4bRZSsuxhJEvy7+TE90
5NOlf9Bvk0uh7tvutzfLAZ3c2M2/3h4FkTz04PmbCKyip0Ax2BLsKCav+Mivfndl
wKCjBTNeBnfXQp67ckPgtPhAPTjTvLQLGWTUWauFUGvOUO90QqzdG8h1WzGUOJzo
Lnhr34n+bb0FFyCIz0ECaeV2OIYQsDc8BUT8DKU5xHSg3eYe5scwmcPBQl9KZ/0r
A9jR73XRwNDXv1H4tNFUR5Yh+DxDmwV4xw9VowxrUHweV2G+n7PHEuH1yl7ppJ/k
Oy8DkBLrNzB/hHnsnmAOUqnLq9zW2Ot9AV2l+fdmdxUUf5jTgrsp0trBHp3mwSkz
dINHSofZXqfUYpNilBa/ppPQ3NcS87sh6p2OVz/NE/uYPPUXyEWRn971QhcwMuuA
tf+HcFcmEXCPNzg3Pd8+vfYNduKJFSl0jpinpNI1I7svunzTxiWn4OTTzXHuMX5h
zfMoJfNYoAGMsvj+JyIKAC8KgrdGoVXwg3yLzCZztYD5WwX2qxWQP3n1SP1W4ELy
KT7Jd3BnCNXMJuQORRH3UYrNlhRWog6hVJogPkBY8rTNYtXo7+3+K3jaLRAF3yS0
hj3a1XnUAUa7DwC7BN1b6u96sgiTL4qoy4T1jZYbWxMeQSwe035aMob01UtWgOX3
NrUrMwBp5pB4u+H3CrR4Ccm1fMowDQdNa1YhdavXj1xbqpB6slXXxS17W6/s0YR2
7WK70JBFNyyrahr1XPhjIYIkgOWIe6wFsGtuGVcEvDvLJknzc7etC38vCEXFTrFC
5G/Epa1IeV13YOQM5xN7NZCPYLUxe90vyRl7p09WFQHu1Agv3XQv6AhmQiI5chXi
q3a7dIJe9Nt5Dhtjk9w9q36ertoO7Umj906mei1RU2l84BbCooucoSFta/qA3Zeo
DOzNanPXTY5/CdnESmCR+CUlc/5mZ44oZmDMXSwMGhkImA4Gz3xS39DiwayFDRzN
HGKnG0dfXSoHr3Q5L70PP/Sw3oBq78qb4kHApma4sMy4rx/bP/X7ZdHWbmlBdQtr
JuI2yCOG50HMgYBzzHSPqu4fbCY2PoDP5lYeligwhTBjHgQryvWTpxgFgG2ZKpfK
nw0lnX42RMLROKe7SWWZ8m4qTlUuEMbIbp5U5I6fTZUHqvFmjR2ZohCTfswOAcmY
WAciK44Ve48l2zuSkUhOUBFeTjgnbQfxxuTTrkyfhnKpmgkOM7+rJqMgdP1V8pNu
602mKnuQ3Zb8Lb5dFft2Y3uPnmk8EnO6poBJHbKeIUXfFGnxYH4oT09LuqUprs/C
7q3Aj1bRmqtfsNVDNw2qdSQx0DUtyPreJoLhiNqtx+CCQFDNX0xFCoWo4fgSX8Pb
TvWc8dmdi0vOlViL9RvpFBSbc4kZrfFpLrOmLgS3jJJ9NEdDuMcolMzq1kFxhirZ
1W9Y5vliK7IxAlE8Wx8KhDNTtUprHx/CDj54q+00y6rzMVK/HdbVZqpszrGlycFD
unU6B8i/v0Vwb4X9lWkhHKI6sYRLlChyz/BkGcrPHadvdTNPDZSJwVhZ8Mj4A4iF
2XDfQhJh/2bvkmz1ePFxMLh3foklp95fpVUe9Kmwfbj9DQdez0WEje/gfBCiQA3B
y/LslVtI0a5k5loaFkW9RatyML4T+FFxsQ78jTa79DowOB04YKHxUXgq8SIffFvw
artHA1iOyqjROwDmp9h/TrOIC5fryhifWeCGktmSt8J1ERQHy25ipJuvEy0/1XHT
9jnh50S8W9j0NQm1cBv3a5hvIiYvrdF2E/3cPInB8exzqkN6/EU4dbg4EMb9gUW8
TGslqyXraQCSs9i3WWywZd6vQEpYmLzqfrbet+YSGa1gY3AKu1sYVcIf499hoBbT
nF8n1ABn6DEy2SuZEIBdavOdb/fmvi+huOvzSz1YQLRezfOPccG2MJN35tCDwOkH
r5usAA0BPJgvsw8+U6loekY0b1S2N0UyyhA4qItC2PprJyz3Vrma5b4189RgjD0n
gZUNoqSI5mqfYvTIMHL0OywmWJjt5wNqG0MnmudEDeYmPdW63uEjE10qLjMJk30K
t5EAO7FUlaCTVF1GugjImFp0FZ7eFxwEhwZvqyfi3ax/sXUw1f2QKl8/1R8hVSK8
kj0GNuVoh3GvF15R7/Z8R5QqM6ptWsyX1tiVCB8kEjb9FXcodmgiIXmLWMoaQCJr
a9oZNVxVG/mMQUgi2SkNqvTPkYt6NTAYHPof649sFqEd+3RvgO+FPEnQ0EKh4DWz
SYTv/h7NGBS6Wydv5ziuuDz2CtWxOOq81u/n5QnVoL5Hj8RUYfjuZHzN36Yap47J
p7Zh27sKz6/lO6nUEsDpZfvXCsksuQKcuuQH9DZq7gJ8ZeJqQKSyz/qjm+1akY9A
Xh+qrTrllmnSfzEJGpBhuyc3ur/CkrYvoxZV2l/sVm9uYBKEWQ1O0SKJfqGVu5K8
T5EE/ZXuUNPtw/jzPfuDtlZVc8h0ifLWxZzncJuT0nu7E8lO+9IkbUROKg7jWN+R
YPKqlHx51tdHTuLsLY0c46CecbWz3PjjPvTpk5sGZ3wIC1fiuP4UVquAeeR1iPNV
Q1zsmzQsu3GNkjkEt23G5P0W5K6POEj41QKb3J/KEDnWLV9WEuJIX5+2Yl5Wk9Zd
PeSRNAgYiR7AlC2s/tJEiP79nkf5cDWOOSm7Iwu2BxYzlYhTqrl7YquJofqqNusK
O2kDoOS8Ht/8j1eJODJv44LnIr13/UeDYkY7uTzpjGCO6HCW6E0goPNNlRWRefkq
VgvAuM2rjGZ7XrF/w06kgfi49fJI6QMgPO0Xv7L12ZqfliKX7NlS9DAbBB6uXikM
1i1XSm6IjzcWPY8QUkc6lzkSvfPtwoN2zrxPv3KnHfajvXdgNrSzR7UPSAVK4Qxh
l2LNjK0JmIxAP+QHujoODW5PoYUqTfjm7TDed+5z0mQ1fNAWWhH6WL3HMiPXqmq8
nIOSTlN5fpqfWJcVoE2V8pFJdtfwvGxWGY60K0jlKg+kpbdaD/0yFVpuestvFxpk
xU+h4r5mK17cVN26gyB8R1cOFsRJ67FO8oVOgzThLv0rGfgqktyQZcbUNTPVdQeg
fCUYJG5KIJQxiKSedrTXJqVLFrUqwH9kzo0ZX/4IM3BCO8fHYwZmfe/Po5rinlPK
wZTmCogSalWsiv7nyk5vGuY4eqvqRhQZsw7VcF+j26omPhNHYHWJIndMCgBS8Qon
FHxNre4YSvCjEk5f+vC5XYPDxygra5z2WmleZc8bd/GSbWjrWOAS9ySlMUrSHUbQ
u5JHddTa6UOnEt/qhavotiS57ZTcg0SO/p6G9p4feJ2W9Lk8mbpFer02KDconF8w
H4sxxZ15vJaOIjiC8d2shuAYqen/kkWW3qsqb3SAgvKmt37nhS+geXDoUbaEPJt/
VHCGZipFvYja7R0g5kOdMNMyW2IWvKSgM0OFVmWffjP4ue/vR00TLh0YKTR6HR0B
U2jRL9PZY+TEp8UUu2bowIsL4xgEIi2Yk6IucAJF7IZmfB7q6P7iVjpWrQNO5U5S
yCQaGETAHZSf94s1BSVcDZMci9mRZdBIBdiuleE7UaWGyeOcxojK6PIyI8z39ChN
LjwWeAslwr2v6Ds4P3bGS0HUUXRxYTKewe+ll7mA/VrNeT8m0bjfIbQqUVB+kpw6
us1ziARK8mAujDPK43ECke5HCCZuw5Lp1s9krGYmpiBUcypYWZFdiyyJK1wWpwcc
5I0L0gAPA6362+e+700N5NI67Iai2IayK2E6RpPylcjHwlLpKoaeWsu1wBF/FeGD
CsSa4tGsgrItr/7mK9K3CUwnh8hUDHtXKytjtZL8YEuFWdbUmhfr6zkCTfsCoyRW
Xsw35+zMobd+kuirMZQLViB5yL28936/fymJaCsUy62hZ/Mb6MwEI8q8mqE2O0v7
FYs6IRQFsp+ppEP/0BvQI9ulghUMNtPgPj2/K7hrrYsCQwafUK0HJXOo9P/apgpO
iNHcbtN+HXizJjfvK5esVYXckbl299u/PLIILtfqlJPyFNqjlxX8Z1QCflnotuXK
/1IYquPEVwMdgZTQkwYmsEYel838BKkmxUxc+DkoQZglMeuNApZlTJwF3DlA6pyq
Iq6Moa7fUcqXNgxkRoyw2vxX7v5k/0joeG8dGm7QV9kNu5OrOwgktqSTMqCi9Zg7
ODlWzEvbIlftTeoVA4PCSQDU61gg9Co4K4X/iUGBu0Ea5vAinHQ97QoSExIwizhI
9DjxHV1loQ/AERc2CWLMNpJxwdUzwK09vXircamUA4+5EF4nLJlNiEWf6NYpr4jB
WR23aq6ZC5LfmVo7WupIm8R8OiU+XyfDMdLAdjE4bjrC/sw81ERqCncVtW7TBFYG
jkv4DaXCU1Wnw8wz3ao3/m17nhUL/Y322oFoLQl24zu7woM3yILvx432LoyCJxBd
lXxrZtO4n0bqNXswZ+SFqH3jVgeZ1QLAOefgzA/ojr7Jlpulj24ANAYIYF6+Fs0U
+9Al6qv+RyI4wND+5kAgfA6z9/QgzJSkFWBdSr3cybdLDvXPn9pOnnwxC9IJ+3sY
nfduPJcIyFcU6pykIvMpbg7YjWN7JrPBBlf4e8fVwkK/c9XBTiY79GDf6fO7Xr5h
goGsa1hb+zShB2NPYDHeUEfVWgC67WDxE1bTPrSxMuJdqZFhLYYPMteBhCzZCgFT
n7n6PuGsggjaBl8/jl28btQzt1CJacDWJc2eRrsVmKfaUzeIRfndF3TFB4vUtocX
45a7d/Fie8p4rh1du3fWadadtkMUW+XpbvPLh/DyDrz/fNzjS/tKrNnMGhZ/8m6C
A2RMeWCNlrPsS9kB7pxd+r/PpaQR1GRY8db5N0UcUKtfU8PRxBl104RLTvTIiY4T
TkDItnl/eUEUUt6v2X7DynP15xIG+7QOs/YipjG+Vulcsk/LNwmJyeRtSIN3awFx
nbNqwzHUN8sg2yarRydBs++0bhFeYMRYRePeap50OJvvKkl+iLVli71kZNvQxxMY
3QKlQcn1kyUUZiIBwvU5cLyUKKcxXddtzQ+loAAR4yPCGEjhNeYMyg1DxH3+/mL5
ODKV4Bif8BwyZOMaw+kwWcjMENO+pLh0eHC2XAI2kZtd6Arsk7T9ptcuiaoa1xQ2
7IFUky0nlKmDkyV+hMIsCso6/gaMAIB2aLQCG3YQI/+CKbuzyXtNH6RakPWNhIcP
Gtw/Nx+DxBUmeeiK6AqRyWfqilpvKEUWAIrlL+wwWEYofdxNfR4hPo5dikr2Yh8U
yezV796jAQCZoxYFSzPws2NQYmlsEjoSMvsec34cU/xo+SWkSVrVllyJWqcnIVhR
PrWVLasAsRYklUHT/4YGaMgMvbATh1pZ27plkvWTyz2NzdYAD35p7AcWGLhZl2QV
jf1y3/XqvsuUhJsSwyGxoVXgL8PPAl7Pk8firCBJKQ2fiLREYazhhSR9Dt8/+a0u
GMnKdz//k21ADuu87sA6koEZboVdei0y//soIlfxxLd5hPJTFPAiNv48F+K2JUdy
PE0y89+Wv4KnLQZoHZ602+SHMh4VL9k5c4pC2B34FcwhfE1hQs09gVBScgs/Owk8
VC9m6Gs02pb/nK9ifdCeBpVGU79l2cpXQVXjKlcxF1Jp0zuj3v1YWP1GVU0bdk7J
4eQMPLJc3yVH0qFtAp7mRe+z4Mwmu+fZElRtAkrW7lB0h1zZ4+S8fM/pEKp4CNRA
4AmcN1Cj3Pf6XC7CJZmrx1WVEPLKmAdgu2Mn+GWI8zE6035Ydjv9QdO4mRcxdgR5
lFdR5nxCqi80aWtMLsZLzPkpxSqChy4qVY/nwPhLe05hmoQ3BFOmb4ZbpVzQhY8b
fw6OKWbBbLumGVNH9UnIIb5IEwYtuH6abfDwDJZ+Jimm07wpg+wZ80Xy7WWhRLMD
g8dqALtyTKhSOtsBcO9P0wLocTjcxuCLy/LqChe5/ZWLX+0/EKlzR8lAFlSz6nIH
47YU+xXusWW4jZavWyy3C0t1uAxi5ci+Jp3GKs/x6CphU97WTY1xz0e4tAQaBacB
8AKmkGV55tuiQAXKjot1WaZ96W/wX/h3wtEYrQNNzGiV7cQk3o2qOU58UZmbQjx9
dEV17qteK9q/9e4raJfIgeMvjwqQPLnd1IgwKmlynuzv1JZyg7vUrjFHc+6QPkSv
hiHMQLREOvK7/w7Nn8yrdTikkqd1O/A8ZiiJ9aVuCnLnPEH/Wnn1XrqIitYxFydv
S4mbZ3b64mjc1gG9A83JZURb+qD8mZcqNCOj4+tVaPp69gQRnThe7Yr0THcmKxLE
R0ZZ5nYMvTgYmAjkOEBjzoZOxhOctEkhjSubtzFphAmQ8QQ+msSXmnJ57/oz1Yy5
XLLgi18dSztLK4FElBUmXF94Nb4vEl12K8+JhtBNWpQp8/F8QS2AYOx8Mgsnx6ts
PG4enPZHjpCv41q3KuWn7WyOoOvp8M7PMYJTzKfbJrXw78jwSA+XpuUpzP/xSuhl
VZqbMDIfxKEiInq+yx4TA8BJkGjv4PnQzC66YegCKcXhe5v5wy3BpuxCFs+d2UU7
DYXVZZOpWvKFfquAmB3OmVRbH/MABmmc334QJ9R4EECr+rlotEqlyEg0/AmMDzGq
yzH/OLFgsftnO0IQ2IwXlWdvlHd8d138kOxSf1ejsRfbGn7CyACRUF/RRb6U4r31
JGZR0RYwsnkOWw6Aa9XlbnGSbO5kq4IRQ22IzWgjg17kbMgRlRCyUBRSgHdabHmP
I9zlRCIjT93UsDqhDeKQerEWhtTSmi/cwHGY9rssBPECQ7J5KkE8TG/3ZtmG7vLB
+13JtKQIzb9fmsJNTP8mh3bFKGyK7rP+ilj8k6pciXuO5jtH/SPRmkdbK9CTLdsA
JQFWgYkkZ2MSbOKsJiT6ymfw/14DA9nFI8TWfCpOgQPYGH7d0CWe9zTHslhFJVmL
QFrx1xr6Z7tjOQNFLBcaA0C0TXdoFOnd+ocOeVcLysAfRhgwPlAk4OfHHmV0WxS7
e2ad1eIUTaIjkhaddphrLkgOD/2kKjLfZRd6TynUaZbo2gYMwQ2/m7VK0LxNZuJU
RDOXgb855yRhWvBhoOtY87tdxO+yGM+ZShGX/y1McLHNkZNWTvTIRm7u3DHmH9QN
MrCRDNq7XmKanbZ/iT70cEV0yHj2VnSg7rgDJHxGDrVBPxewH5K+rqNfTWBFGVwN
QM7CIqHM7oAjH2WeBpY8TjYrD+6SZFADicdzmKVyUl8oEH2b03awOryqtvq8IF9g
LM580VmWdTN5/9OqmsN3JvxNYl6aeS3bIAdyv5q4m5+iWjDcmKLpg0WErcY18p59
cO5SCPUryuBMXBRBIQQJkgDCDLq8CkoQ4cvqipAPCTmF+UkF6U2cWUuerq9xphFR
6RVgT2LNpxsMfJpdsV0JRVVRMPok15dwsTTH3Qiq+lA12DiqeK6g/iXRhGEcvdbu
BdmHKg1RotXbDhCt6mOQl2mUP1hu0qDs7fOTF42gP8efRJzqaOmwQ+x2kGWhD4Be
IHOkU72KCnfUZ+pNAqgx6MLOgK6ApsXudTLyvywpoZQzIdxyEJX1n+hYxmM2vljm
t9sscQIDgAyyumN9T+l1xr6ZJzFK5DT9XknaMcKi/REsYGmCDgYZC5Mb2A18zRlr
amvdlnSrNhOTeJTbfWmopRmCTlKP4abm8pSmH8llgl/9ycYguQ1JrYsUG1Z3WaU2
41Xs+R3Tt5oNUaBdu2YF9MDBbYAI0lflWV3WGal78fYEJE5XnIOwNrjXqt/tmXcZ
aijK/KzHGSVxVdkSmFZmQoT+wUK+kmqUL/Q0mbtfG1SGjPlWJKtFiSLoU24kDPXD
pxuRTX/gM+uBYFVTjxf6SvBRqjiymmy52qg+QfkQegk/V0T2w9deYukjTQXeMQzo
8WbkkyOkbaD8nPNrA8qj2sxGFQOT0CcxL1NV0ffKYY8DPTixhLnoRzPaHJeEKp8y
JmqBgGfucc/4p/kUGeKFe+AI+jXJ+qzkPSajq7jH1CEu8ntE2JpnJL0wKHlXqxiP
IVzO6xnqCkxKbalMkl6od5rNmuyr4azfHqr9NVbEEOFDmfzD1cYWmnCsnudXJuIJ
SVFA4V0lqmGWuNsacS4eYs/1bY/CuX3LDBlg36v/rv4fjZRrXbI21xDr4G7MELtT
MFDkm5ki60SPGJc8GfVIrNzimGoM7J7GCvxY2VqBSM0TSrmzE+6QuNa+XT/7ZVpE
wfMSlx0aC5rfnMjumDcNa0/m1a9Kn5DOtei759qKEupWnVQDtDwrpiQRRyoswsOl
mrUiOPdK4a/+Gdv4ggzDMH6I3ZEeSMiU5fMnS/qWazBlxu7YLREuOD0wsUD4Kc9k
0WaN9zj8e5UToZHuvmz6OKAMUcTcTH+ELWaAca8UzmiP5x5Lnlpbpcx9PKhkcrQl
SAeXO6oZaKGf8kkm9ee8NL4LneTIyPrM72IMrGd6a+UZupOeX+dfEMfwQvFyZ1Xq
ck2DymeX/qUxNiK4WSP7zWRNyNZ7R7SvRWlnzygFVw8pwuymrFUjkizPOiVpGwZy
HshCIKoJjjcq4/yv7laC7TOzD4SKprtANWAAdHa8AXS3363fURJvOtaZFr/4PIzq
FZVzjGjQA0bDS/XDzfq/1M3LdWNHZdlf9IW1J32loeyOQipsQut6AMS1RJNfFM+J
trIQkEPX3jboAX9tPiyCMGldJwFTG+8tpmVq2haVe/AAy5OiGFs523srPgeccLel
uMwTSUaR71zFh98o9w5A5oRsf0qiK3GV8we1m5BRoVP8GtRa7OsCcnegeM3FtB12
pkQKJu5OyNoXfo1tMpbTBe9NGC1tZTSx3d9fzng/g0A/DXP8Tpzj0N/EXVJvOcek
I1jgfcF8uTN7xl8u09SXHCJ6N6otrz8W8ONAT++rYG3t4PWzQKHrcYPNJpM+qKzI
x5FWhPNBT/wZNNmtIdAiv9HfdK0NBDly6V6aKLFzptPeHqDAXu5WS1zfi/2F2hSM
P+2gxwUjO2OCywOwE/iNRN2NbkJm+I3mjmIK0pRdS8XtmAW+QtfHYLHHLcDY4AtH
glHmMbItQJJ3+ED/ablSELcvOLJEuzaD3xw2UTyS96S4DYSN5+YHFqSDrrm7y4VN
kCOdZX6C3Q91v5iFAl8bgejxt9JahVKAVDTFSbc053rCll2fQz+iWY7NsRJ96imm
thh6180MsrgM2gZTx9i99DsO9NzUYXO3nJslxlxXB1LsMZD/iozNjOsHaw31UG4g
wseaoo410slqVRAhFqRD9OrLeOmobhWsWREoCGFSq1p7JRLUWekksBbmh6Wl7Dju
PLGmpPmkD0BpGNqlo75dj5Al8QzBxQMuMULdKEBy35Jo03AJ0zf8VTITR530SnDJ
1m/ue0mzA3zHizw+fEZmUOJkbrXHEfIbFVouawOjbhfth7EuExz3cszJyETJPvHC
Koon0dAejRefnLySz5HmgCkR5TEHi3AyBlX41mk6MoboWWTxmbU0hGvyRcwx0OvH
zUxs9u6yXAMWddTigSmGqZqn2ynH3pZaV7l7jj8nq5tLcI3AmaEAl8pGsCTcciN0
MdSMVYqinTusrfG/Pt4OtHegM09ir/iRn7YY20UcSM+JdUfhMQErwxxzoDRvYncx
f+Y60eW5GBXcYDg0c/0o68sN2TRJSg4+DJ+2fC/tpOCuLjA9Ng603zYXDkWEWb9j
KVcad7eMBIg6gBY164akp15G2lZ4Nr2zF7kjZlfkRBPp30ymtznwjAfUiT6NmFn2
wKoF7+m9MTnOx5pntWb2BKE0KmVcu5TgK1GPTASDqONWsh1JhGQ6uij8U6EInQKE
ImffswmFcfWe0kfqnP1TvZ2UXg21ooEDCYLvUoThfYNyuif9sbvtVGuZk8bM529+
2x1BhDunuc8b4xyrRndb2lkvp+Z6sYADE7rPh+8nTLfWv2hAMJRyahI+Xb2/RodA
A8/4kR35N3e4iJNhawH3iR5kmtHE6OswyQ2F9t4ASw6CsM51tG1s6BQ8lsl1W7PX
DjiAm34xmef3xHNw1aWJomwSsESQW4zhB448fvdSceS7e3BJs+tzx6SVh5vCX/Ek
MgMVt+g/ig5Lvn9bTlomqEmwgoScuoSY1rLoA/etr9ABx6IbEXk4bc3siuPFzDh+
My4Wk86OL0XISD9I9EkUk7oEhd//xpEx3IyZuLnyNQ/RtVh10VFeB+Mo1vg9WK/W
Lh7U+5zfPvFdihRDirfFAxEBKXPWbxSDw92uLPxMl2XkoBMomi7MZ5NYJFDyld8g
LEzCZ29AiOtn/Oo1c8vGz+jp1BghQU4Q6pdMFe0jbjiaP4jcHEXEj9B+5MmPRKmK
kHN8vd9SrvxNmrInGke+WNHK7+p/5ARxkaP/0aa2Kp2i3W6+ipURQHUUQFlDXRS4
i0vlPuO8Gfwlues1+b2szTSwzOjr4YcMrmpDbDGCNBJSL1v0l3yeAYCRajc36YM6
trT2+CSacupwIv4iiN4cp0Os/K0vtN4kPAr0yhlN6DO93uUVzz4RrUg2JB+mNUGl
LNPcdr5xMLPizc38+RZWNJ+zs+MSFQO8KZWZ2T4MaxUXOEqrPY6B6JGaOQYxO1Mo
EzrZrJk1iS9P3Js1cRU8gI/8MMFZnKHgwN0m31NqD5Jp++HJZxaEpx0f2lEaHv+m
UIjhhJwoE3osUikZsX/OpAt9gdU6RRK9GT4OQ4CiK5N3phw1Bz43CiQtQqrJ62jm
hn1+BxjP5M4L2ZF+oatwfIEJ7VhxScBZ8nz1YBCcLQRaA0S7xgzKP17wsP3MM3uX
Ce1rDfBJf9dEqAhZqEIlNGmrzymMw1AbFqu9caneGu8dXDAmCkYedoe218zfghp2
2YJROg+OmqU1IWidn7IMv1mIu9jLuXX2aVMzzqXnG2820ApzNcrWjKMxRQkahIvn
E9HWAoWdAKMeG70SMFOMwRz5yEFSfZ8ucd3OALdDHN/kckmohGJSIbbLzbBii2CV
EL0GpZo4dLl8ECKg/aHXB+rW7IiB2XWae2rqR4AeQBRbPMl95HaYrumrM8F4jbyj
iJyJJZnNaWtaqNmIX9ZHrZcqToSJ9efOH8N55vc3Yh22AOxWO6vyqbJzcHefHW0W
APoxPeJ7e8yczu4wnPV+fLcF15NluvNGWdupSIr/mcDIHZQ5G52LaMZzpxRF7mub
TjoV1gyta6zEtdmFx6Ud/cUIIFTneTHDZfGFMo2yZgUmVxyonrHiTMEtKpikJlkT
EH30E3bzYm0Is0FzI/colkAaaGduqYkQTvgKOvMtAqw2YelEA1badEF22YEj2h1I
WxKwmKSWsAGFoWHQoGxC97j6/CPe/D/KyzJot3fzbqdgisaqePCTbLeuyzaK2JUj
sjiwPb2pdeTptGQ+DWCpKWbmVWAFrxqfW/VbxqiXnBiKcdcDUyyuxRW18yC7pPXP
UPmNCPxgtCXmvrv8NOiOvd3jg2ca1D2mILZ1mZarqK1T3+YJPzMq58MXYfJiMuD6
AatIrxYCWzJYacEhpmqy8gWLJy26xCWE/pIVUuCbqBJl+3No63EM5m+n5Q7o+72p
KF/WPzE4fcy/Tbejv5TH8dhguMrZRTIpkt9FLD0Onw2QrjHmszkqwMEEuB8OEVYs
5sp9JzroQABA9dL85Dmu48ycEfHBmBmBgKULrl4IlR06QW93Io3fFSGwB09z0Ps+
WSqTrbQ2VL85eQ9dWW59kYFe8qufTn88u5U98Cqm1/ej+dShTk8y42gljXaNdJwe
6n1Z8F6d8snDg2fZu69YwvADQoQNFpFX4nmohN3jCBo+E/iNZqxlRuXOH4eCE3JU
U+Ilp4JCnRn0S2zWtHWcYdCUagx88YBHlrP6X9vohzyWfK56uFeU4Cm4k20RkIfa
FwYPdZS17WoKcYFAoTMSUP25ReKdHAFUIUevTmlneTguHinNU8WpBuEY16ihvpZU
qJWupvRbY1SxtzxpsWUSCnqAZPrmroRQYwwEjeZpvEKjctlWIioUkAQyAr/yUn11
1b0bZMImzoIbGUq06XOE2kujq7inlcLiTj33r7pLb1Z10b4tnljy8M3s5j52TF0+
/9T+Zt7ZnEblpmqIQWoRVWJWyYE9m1OqsRrcZYsAQEgyeJdeKLImt9uH57oW4HVs
s7uAOZW4vwmaQTZPtFCXKl//uFEn6/tlSB6pNEZSf31SyxiTHJr8W0SpKxzOrrut
edi5ElE0O8i0Qd3U1xzXo364miCurVBfRPIkdkRIuvSDOOSycSP8MileY8sPo2BW
+a2TLIoTQJY4VkIS51eQX8CxdLvxbUF0Z3qeaQxdMqakbvh3jqq9q5ZnPwz+aG2N
VZ+fcDeKxzGXj1lWRkWzzEVwMA+yEjOfYoMKeQHE6ujWHWOVNTtPq2O3u1kDCBzt
GUPAcqYayaEJwTOdfi4625kWylUv4/q3CCrK1m3JXKGOUfGfUfP69OKOCXxH2yFg
J3W+Ke0ZzjhOXhV9e2iVaHfUFLU4ki6JMXFCVe94580ACeD3S87t0z0KphaW8T9/
esaei5weXrYVA22DW1xYV2hOUxN/8ZaX6DPBtjcmzJQrASvmCOTu9ELTJdwnN+gP
kiQgn9TTUYAnrj1aDxiPAfMHoHsFqW/dD9L1HR7o+tqLyjVHwdTBYm9fhLmxElz7
uBNDw7iXHYC8ECQL8UP/M0W6e+zp+UYPQPExutkdVRxE1ou6q9Snay+E/CvkZIKP
cBZd5hqacF9R0dVt80NlMafTBUM4zXIjeIJiNBR2KTsQiQQjgEz4R0nDvxTSoxYj
ydpeSRbBp1GpA4fc416F8p4ABHxi0UrF34lxfmI4YwwjsUlwaKt7IKxd+uDdBvgc
Qu2CD0NVGqCpIrEC8qlP/6cV3Vcn7Gjy2yzbMPB+TRH/KdmZe5jwNUPvRNDodKtt
Isz2a9xUyXZknXLkvXQIpGlw+I+3NyPEKyHRvIL5ZfsG3V6cSUBROR0W3mUxXOzh
6KjVUG3KrfrOFEczz7J4V38q/QstlmkAhq4utX2BGtm55h2sNYio7j5KIMHBb6OE
yHerCe4RuIXlSVt33iSNxqLxKaEJUOtIL05RpSIN8qOOtdoK2fPH825382sIx1QU
hoCaopXdVnNe1xZsz7WPLBdHoPBerDWcKCR0ZNTH3tvH9PdQ6U12jlEOi9SO0qj7
evbJQ1weXO12Wa0U5M/5DcZUuSmnsCqjifbv1GWqzbchlwmstAh1azhlJEW3Z6Ix
JxRujaz5Yi1/quWkPj6tkgTgjRLHsabSfZbGFndvvPddGlLVsZWT+U94ZPeNeCdx
DRmxBeMrW/ubmPjn2HQvW8UEKWld6vwcU3V6R+fnTukxlbon4Vol1ZtqjrzGmWJT
PGtbU91HQxEugU+xOTyOtJ/x5H/tjTOqwZczLhmrwuNgebBJh5+cry6vqouYJTkf
oqTYjjEcmSvyKT/cH6LvNsPdv+ArOEfOcX2BOoRfoWgDd2i/gDV2QszenvxP5wLv
3zdG5xu/1Eczc1gksUXsuAlZSkw3j3Xk0CXntPMAGZPI6JDppXcX7E7CVkU4kR2d
9gOZO1yryLyWwqFfpSJU9K8jSvfJBOgBrS8343fdyZTRHe4ZJQXbTqkatjkjzNSv
yzDrhXdto/6Ky4bin2L2q3Uf95RMww3p9bGmTC0I2xYmRKym+l8kG7cfmL6Bewr7
Q7F7lWROjDZJ1/1Ck4vll6vLvyuBLMCrOdTC7V8q6m5VKBRjevvIHcesU96c+RD7
0NtsIMOruIpn2YNX64YS8VPxcZURbMRQgq0xzWuSqaxhwllnHzj1Aur5SxIhz+GA
yb5qXy7+mUAMTxXIt0QReoA1FjD7u1C1C6xCSwf6GHfBV19N6o08LqqdC/1opCis
6EmldosedFyF3AWSkMZuxA9/5Fo3uKluyULLErhwLtWNFI4nF+SccwEjSpO9bdaa
o3GtncyyqRBRJpj4zIYdGkOLOndUOwRaQ22/y8reLKU8UfcFS7jFrnaLfIqX7Jan
HYUsfA46koF+LW+qBvViM/XhQAq71YnyEqvkGPcUvpVVFq+TSps578rvwHrttNzq
x6GiK93bo9AWMjfaHfodweCx5u9laQU7N5LJIFBa/Xd2Lcl9xRh0VGm1JQpaUVkh
f/Tl7OIqKkqy3EQJXzu+oojgY17DnhBLwBnWGr4NkZYZ3JZI1Ud2M9o7JtbqP2n9
Ih+8b7mW9s5SrAXqbc66qSZMMAMi4uZH6tA6khoCRmubtp+GdmVYgM+HSnTHrZf5
yBcTfETASgO5hHMjnlNu37VX/R0HtQGrhfy2A+RtadtBIphhTFu8viwV4v0EtBdp
H1FVsGuAhacKHEvqg9YUHBQDQnFnlm/e5IzHCHefn1oLhMUb/AS9oA900aOAlhVG
tbrbv+FdkIP37AM0gTkGz7dGugpD/YoeN2wbswojFAlsGVr0wDcKuvLUaqdqlIhb
twgF+xixA9lijykYrmofrKiu4uoboNCzcdcfxOvp0XDyjTkOk2GQTfPwyVrcO0D2
fTaNOP937teJNg1C6Abyruh1PEA9jw+9DEtOApR8RaSJr+MpdzKCIDLkzadCI4kk
G6ogPSfnYwtKidQKZx4ZGNGu8EKueoAaVKhp8E0+EE2jioiJL/Q3iqrfruyRhgae
wrRMIGxGUqT0MtRzojqCFzzjdIyRiQcdt9uNKGA90HxSiFzED5W0jr9xUXzAVOz+
pGYms14+k0/9WoQL3zmI3d0tIcuwdIfy3djBtGaGFRDlJ/rg6o3cDOm4vPLdDXYf
N1jCuJXDiRoJvxUjAFDT+PAQa0Sf6X70IGJpMNhx5OolSQgEObRcR1cvExi5venq
g2EOSElCwbFF42LFj5c/GhUf/CH85A+HiGQQypX7bcB4teKuXXaM5va8okPVHnbq
7Iq+NEqlqdGekbYKzyI5pbKahuCmZGmfZBXj74T4Lweu0XEJ0pjtRaW1GRW+Lm4B
xFn5xiDH/XEDR0PqNdB3qd25F+UW8qXIg6+L6DvCGsR7W8FRPMNa+am51r9HKNez
f5s5/F48G6EkmzGfRLVMOcON0pb0tgboqEC9ty1cjSp6F05M+tth/AhWTmUfOsBp
zOO1eNQJMlh1dli5OGj4mDFn+h1IEwZPMV/HqpyieukE6AfVsz7eWvyvNJoaMvBS
jczKWlF0pP8jzo3ngfaprLp8Wk/u9hosXfX1e/v8A5w8Qp9pvrzxPadpyHO82SkG
bJ4YVlKSGSOB+yLVLybZ7crJd+cUiu0HRUD7yh1/CCL/wS3iD1Cqkh0LdEcxAKDU
DcvqyV7Ryu9cIc2K2mjD5C6o0t5khcK0E9t0m76ykT1ng458MbRoReiNthc2X1D5
7ctsNZGpZ3i8kj88Yq2q3KDTx0nqK7KwxSWSGwQHeWnHnf9AYzzU3FwZtKY0mZ8l
JxfqrI2DZcspfpWnNc+jSXKSuMuvdIgwa9yvg0LZ1DHyw7T9FN9NxvPRqs/hy0tP
/ubKlU5YL6yrd7IBh5TXU5YqKKji7wnbfDqBSt3Az57R1dpKlPxOjNf6RAE9Oq3G
1pJhmwDQ18jOMWDLZGAuSeBy3Enp633YFbEvVVs4HzCoLQdol9q/aFI8jKZdf37d
c1HxdobC/+r6jPCwGKvWRG5uPIjXYTJtJXmw3GRVIv19iyiT2/kAiMPtr4E03Obz
M3eWjWm8EIDFLgt1Ev6CYP6yP0FvG6dAYfz4aED71Etok1xIyYAr+lqoU7scRrr6
zBpEbSGpD1Q7Oh+4QqHp6BDMqVZB9MwzjhmUPMYFg6c3VuuNYBjgAb7+iBXILhpR
r7DK19JTnKr2kzYfoQUAw6//Bxa7MeM20WtONwD9Y2KdLqSYpH8/Rw0TkC2jJcjY
7aIuOZhBRUsXdcGBFC+8BH3AloOOPa2Y39dWPpJMbsrfpMk50+5/wcl78gXYAloS
XZV5o8Wjzu+8Q0oNf2KUA4YH65MFuN+HWZQddZwLu6Huo7zKCQ3uJce5r4vkwVl8
xH2kJskwd60SeNk7G0h5CqpfA6T9kFHpMZEcJevEqkaJ6RVYDO5m+9K0e5RLJron
ksCtwwU3EFpvjjGjb4GP1SAwho7BUQEPQxlJSoy8rdY8NHR+Ti0lakdSHZnwDjjn
kW4DKVJUZArI1U/MuufNxpBxP9s6NFfMMhzJTTNSJLQHdxBOvjQZ7YH5F2oSHPe/
lGkUEJUrYQsDJsaUnmbkMfgzOC/JFGicO1T3F89KFwFUd5/LduuwaaXr6r8YRQOq
TbpqFgn8EJohuraxnzlMpTxuD4DvQYF11W9riW1cjqDUME+zz4F/NZNRnL+0wrmS
3DpDZBgWMcp5rj2/GIOq1nmbgXYIiUc1iOsrPL0a1BVDfuAc9Tyy68tAUMDvZAiH
dijXXIk63ck7qIA6tKjtqGFZCezTX1gbp30kWYfeUroU9rXe/R2kVy+FzEnuN6LL
o6ZSiZnLtqgjWd2u5AL+eC07VbX5vZ3ntPpZj9r7NrZGr8DIXfeL0eytd3R4AtDm
YcButi/ElwVCFKuTaeOpHtCg4jHezCKulh1bIQCWIlWcwQJW9c326u/R42bYhDE5
aVX5kIIpeEhK4tFfEgmQJkJKqFqz5lTRG7bS7eEuRbtE5bahpeN8YBOEgfyCXJat
5Gy0oMTStLzhVqfinim1NNtOnCRYd5v2B9sNnj1o4zpiBblEMy8l/3EN/ZgBPazT
aDGrm1ncEpW+icMk15YW+Vz3XfgKSVulnZviN5Uf9tOb0UcFUP0qUTi/K4lCsc43
GaC4t27UpENpKKDSa6S41kq5fHcVapejBS+vhsxjNxGR4U95GasEiEscwpDBb986
XzUerTDqOIM5iwo6IhfULDrJWM6zY4M0y+l5Wj2+4IF/68a4/lv6x+tcK5157B4j
qtlWj0MjoyAYKCo+QXLkdVIqYOn3dA5Z1X2c/mWO7fxm9FVX5Ac92yuipn+WS4JD
Eq6e/DOUVembb1uxW8OpUrnkBLr614R1/fj5wkEQ3KQ1talaaW04FJr0rl86ikph
KVambZuwwnqKd9wr5/rGAqkV9rtJ4ENynCQBYk981LlcYXWuA5WOTysUdJe1JlbR
kD5bt9si7PaMHrXGLf0aWL0X4/+LuqkqY3BB6O4nklF2C3mr7n1BqETblSEvlte2
rfASuvWZLZUgxfAwACMtPZFLqU8CF+RnNvRsKwyZ7CxdIGjkj4fbFx8naxznLhFF
/W3YnVSaRp5yZVtlZhOM+iYDThH1qvFOeG6IOLPCZSv+4BgAmYX+eELXPqj5h+2v
ovMXP5N8JVCag7woSWHIwzNucBAt7uOX3P0ZM15IpMLcPJYHB7bL88SNyzvwewFJ
Q24TSm7skcPOXJ53BAfx94A33eLbZMZFeWg3i1wfsfSp5kgKw4T/NXLVWqP0+wtV
gc50DGDbBs9rx0ZuStNbSxP3izqJ8NKYmdTG2qRfCvx4fhyUmNRyuhAt2VZKgTL6
zqjTDjzxpYzex8wr37WlDlKrrv16D/hQcCosakq3dHQsE/V65xH+3LuAF9Jto2nZ
q1rwdd4awie9X4ShTvxUbbhFtxTBSibryMMPEzPqxoFNzfG+7gWxlxbo74kefxkA
xdsMDLExxo2mV3mq8oeOKHJfAHpHF5KG07DwQ6kK3dBi/VvZr/WWZoG2UJb0A3pL
5Jt9SxMiyPtmVdRVgjc7RX1lzKkgbZWLB9grB9A1469/i0DR553nNxADLxAgErB1
RHXWC0kh74VnQu1H3BVlHeXlI4PlxTfMgMKu0OMOPZNw/BPy4yn6P6Q/7jHjHPsd
2Tbbv5oWjqut0EmCgKmrXOeoKSjOr1QoWVqVjCHPoU2tjSkaVVNLDz6wd25Km2A1
zG2imiHQUGaSsxVUfImDwxYeBiPU5NtUfSFQuME3K0OfUCQURPLAnf2fMAG37VE0
G6it8QFWeedgbLgIHDVpw2nK8vseg/6bU6Gf8zMu/FZ0el8RZSny4p8XZCH9fZkw
7EsvTJhO/SJf73leA65vb7qTBXn7pRwUZUCQw9rmogdQX4VTeh6gn8uH018m6z1P
eau3T7nihF+9anZwdQpZWSZg3GAEd3DXkwyaaMoUD1ZYQmFf7tnApo7T8W78P/T0
5xN8LiM+zi9VDQ3V+mcw2+9PD7Aqa42/maJknTBtCiyCSllhq88AMXbwB9ykavZf
2x2BE73xWG7K5Dp4WciproEDhP5pVrMPd7aKnhrBYSbOsHlsAOIVfUzACArW3iNN
P5YjHczhvJAS7iCNvdYRKmC2D8U8bqBSn9QfH3CPMS48xQBsZKiSy6K3UUz+kM/Q
82HW4OIXBs6yzLv9QsCbbupEVmj6BOwvfELNrVnTJIHIgCg0tj9ZwsAtGAOpR2S6
lMbHjI+RUZk+CGV5pXekM6bHdoEgf5HbccSznaW8bEZjyOHnTUhZjzx1kDQG8VjR
H0PnByLdtsKUBfvnGoqmI8W7fnnXOYqpYL8TV0QOTYp9jvyE7wl/erGK5KZVFazE
4eGUQmsbCMBAtcx666HTQfefYJeYd/3g3Q4Y6HIlWFtBKUV0oGhwIXaJaiwCDI5H
SQyavYEG25QJX3el6TbMr8i4X/lVQF/0YR5ao5Qd49HB5EHBwxfMqup8LKn/XiCR
a6bShYpRmfoxoEvzW8LNpBcgc7e0krfm1bztFk+PF9+ghKTgjxvQWi2f/ROJEHpS
M9S6dGU97Zesrg/+steeQTQuI2XZ5Q7Ta9SnnnpBzMyAJdlBNCfrdewHj2j56qhr
ZcdIBzRPZ6jNU5rArT5lwRjUG5OgXFwd5J17t06gFlpjupSKDm6SIzjdLLZfklKm
Bg6krWR0Bs2yQ4BL+xjSy1Ayl/5FML8abGhBtHtPGUhCQ0QFgs41m4ekWzdc7myC
q29stGVzca7vi2+gsrRRP+qCxTUvB2JBMepLru+vYam9bAPfNWJOGX+Eh0JThJcY
SUtmMBRKi0hbq+B+hbQbogpuweDIHGShOXkm5UEffP3uKpwC7fRunAkOkJ5pPw3R
muSNhzRRsZ0fSEfiGe9HBYLBNBecpY0QlHPp/ixczOroCdSO61/c1m1GNS1leaEZ
AUjZyF0Q1qhFFT3ZfqTWc8qtDJrkuTwP6GFI0a2eKqifcCWQnLQQNk03mhW9dlRN
KaqzPupgAMf9KAtwKV7+Smw1f92fOJjE3jiYGoEkciGeA/FA6B1490nWMQOaPx3w
7T2k/nUn4TM73QmHG5t8mIxb0kaKU9jcovk4r+J0YQib0yslCU2TdIRPmuTfgha9
yEutQUSs/cjmFQCB9bG6af7RTnYT5K2pyXLGrPlICHnWxnr+S6JNZiOHqie0ovtV
oTjRO24ko8L5VFixDHMmkt638PWBeSBUzony/2faU2SOtSqZdHLAowFPMg97YZoN
IXFWl4jBWeSd6IQoIKf70OGXBUSNbbTH1EnLsdH7RU5AMxF2RYTlruNgrM3QzzaK
JD6WwskNWSjjjarPB7hi9f+PrTxLZLc17YpNUp8uE2BDUpRqW8QPSPiiFx80hrYq
P97iVTDnfUaoXUvp/+Q5lMOYZKCfJ6WwtJKDlhXDLmoh0xHox8R+EBgSgwGEzZKa
DXKcskcAsw6fqZWAAXyfZQgcPX+O/qUXlL647Q8pHsjUPsIy7OHHk7QJg+S1U8Ss
6EX46g6pca5aD6AY9CECK7FggCaAOJ1gioViP1a2A78xM9j7dH6cLRjqQgLacbVq
VvHP0QGRwNCmknjuZI3v9qoDP4226lzqCBOI9q9b9TVzxlr2ms/DNoS7njyqUDbX
ibI6Y1IeTrya0QrwydvDKRWXBD3yuHY1ZJfWo5NI4dLKKvVOArqkqLVvuvy/FTnX
NNn3/cXJ9vsfwbGQtmAsW+4vkL7QlI2scdEi6d82Vti3Rsp6PsiayDL69soU8+do
pioUHhe+F6A1eYU7QTxC9WtqSW1S9RlM0AQ3QhHyl7kPkMvO/Pvcxf+ryBEolDAG
0lnaoE+LlUBlbs7nU/ahv56IaBHOQcZxZQKHebNiOM+5IdO/LsdgD3ZqqB8niJBB
eWed8bYKmYZwYoi3fee3cxXv1njInqFG11kih7y0ztuZg38kMTagkAZXMlgi2SMo
EH/bDqAZZNfofv75eo9qoIipDcQhOfIjWBhsaRo5UBZBIyemOpF9wVE7YUO7ehEd
iAFQiJsWnaSfAU5vKO5/GmSqcfXVEw/nYHzAYsUv8rr+wR3CxV6OTA7mYL1Hs0Hy
tD9SQi7L6Eatf9fomqWVe2D+f2ZpraL+UAsoHodReOTzQCFCngxboswVzolSBx0D
kIJNCUSfRVROoGd7HYs51E5/csYEPOMeNdqY6yumD+S0sr5poxQfihe8gAREoU7f
uSKdEH6EdwICicgtTJrEajeOLkBp0HhZ9nfLF3ZzyT2HCpm0+kifL5WBP3xCX+Yv
kIfaVFXbWLoczPGAX+HMbDLYd/JPQyOgo9jHxFgDiwIkIcv/Z9hx/QXBb1d3NQKk
n/ArWl6O1jzbHrYFqYQHnKzpST+57sOvhWuRaioBGnsj7rwwnSsaNZ7a+6NFBArk
C5EIxOzDac1Kqon11+DjV5fEmJhKjEAcdPUHdJ9vjavUbe+XyPvAZeji5sKReLGz
oaWDQMxSF4PxAopHxkMme22pr/lm8rgre4qVTAdmfmmsw8LinGvBFbiC3w8oegKA
EyCyPGFwf7Ra21Q1Qypc29iyPvXmfl41E/fBXCDd7JgSQeAtxVOjMaF407/TuapY
BkNrJ6Aq0fRzz2krM2yU8SzuJuzcls7XP+EinUzy/qqasUDk6wYZQ+HVV2NEOnS8
ptz6T6DNhQNFP5knfzvE0z57rZuoe8tfYk5A2DOsDS/Gy/Fbk7whPxAUJN6uUckV
O+84zk+BOqbk8BVuje6mMOYn5eCtxFhCS/ib4x6oVXSE2cg0wcTabqj7Q9Wg8atY
HkUzdNChIc4RgwH7C9k2qcnh6wGFADbWkTAxoY7fq7QFZb0+2EerfbpxbkWVPzQm
EsyUQwcGVSHuxq2vK0L3BPF+IOOUL6YtidjM3akqbV1jukJCizbJTje4NfSbBT/v
gpbgBnA1PRRkvQBps/Kbp8BbxTFhbNPEeTo42eTwpvQ8EQVy8BLjA9KUnRVbjkjo
JiVsdGFIwriJaACAEDc1pfThVeFgz36oF/pXPJxrlg235GVBwPoF9h+W/Ic17/i6
2OnrASj42LLUA2CU4i+YA7WOfCqbIEMuM2EEM9lJBIOHv89ku7oG1qvPtJSL1vsj
tHYTU1lff+6D6cCmyXJBObY2qK3PQR78JiTixS5WpvCiw2jlNwnmhLESicK9FFME
4mn7nkoiBV69t5n+tccjd1gHRgHOe5pT+0POmBKZkcBv5er61TsPW11xunqWrS/R
XeX9Ck71meR55Zhv7u0Y+94cZOLD0QrKrnJsmrZNfMV95mRStv6vt+myZk+gO3jQ
Hygbh8ky8697WGkghWW4sDKn+Nr2kVGosUJN5oufeYftdY1uLjBEczSly0znhCc8
bzPSduwK5oSi7MgYrmWnra/zgTHqlqdW3s1EcLX5ar4EeEtn+K7e1GAbXGj7fexv
4YzfWYMPHPWutwEcBD/A5lSKtfq0aAYOsDl1e7HPfk74wxxQ/o2c87e6Pu2Bkqdy
A/cSm0OCC44A2T+JZIprSKLlbUZPr1tJmbGSUED+a7WW8TFJb/rAxghWb7ZSHY04
UciLQaoFgnXydYo7W5P6PEHkeleaxkESilHG0xqGcCf4smue/D4YY169VWqYw5cF
A98ydT4hQ+1NNJTG2uY5ljbBiuMkudIiTGCwaDEnOzYU+aKYtpVL6FUMbfXhuhtT
AOdAQlnahnMqXm+k/Y1JLUQX3CB5DB9FqAsgc0vff4PDoQsXfIpx3lN2gvakl+pS
PPB67iwk6w6InmuqFEKDjovk/pLZq+E/e82CJ7Vv4gN9zr0hq3VWPJ/62SoToPzk
Cj8FqiUOMW8V6gOkBNPD6vIx8aHQmm8sICHihDHV4hH0ysWo5DfY1ifXUstUbkqO
gI0LWqTfGW9Yxh/niBiitjJNS4uRDmjzoXZUHgWSiAS3kAB8SiitmfhfFb9NTJFN
WhrdRYExikgukADnXx8AqQnnhLBfbW0XxfZpI8dhXFqNyleUotM4BK2/GYKeZ5wS
LlMQmqusQGY8jhWw96QASDZfPx6WiNGh4VCu9fs0xxI5pXAT8MF5Dk6b8hmJzT5R
E+Rq1nRe4F/KpoAc+oNiBxYuKTdTb7bIFwINrVgnB7/MAfDEJY2uq84fOeu1JagN
QBAjYx4v2GHL1SXBlvRQbE6mB8XRc3NfYs6Apc95rsjgyrBZ3k58AKl6COsIysSe
z+QYcYgjt3dU05eNPhedBqQbgOPf+zJyZ5otXPYd8TNjWxA7WFE1K5osz1Diu9XF
89bjg6k04uE1madhG+azMlyfIAD9P26MfZKJ9TLM2hL1LONZhqnFND03DFX1p49h
lnysZKQucgMIZn4IvFYInM4OV5xNtwoiqKckvD9XLhlHQpaH+0XZtAvtU5es81HX
mORCRolOgHdza+wTmgk801yjMus0tMZDqPHG4CYdwyykq5YHVeMw8xIslv6qJivQ
xF/WGqL4x49AvtM3ntRUWWrC+7/pmJDAWvzm9IkMBsIMaikAixlsnc9iQgrOAWLT
xkBNema1Yy647VvXLUZehjcF/YL6RWccBwdtrN0f302CictihuITHeBPTZZDqiOY
OuJdxC7SCG9oDv/H9/1rqbr3zbVRvsW1GEq9JNlh6qzavbz36Idx7i+6hobAOAie
aooYd2jmaFAxQOWd/kpXzYA71zVgTYfez8G8PogGJ8JQg+OC0a3bMZgTXS5lAHC7
xsYDAaK9OoeaD1TXLBobdDKhQXwOdvxHVhb8eGpSYY36vl7FnHqeP+r2GmroFnJ/
f3Miq2wGmtEH7gaskVL7JcIvLHEbukKhHK/lXaiHTjHx+QrQoFlmEF8MyoegNMHB
Okc9qyb+bm+WQ4HlL+hbVQFDt7PBgAO1YxiV1evr1nfXXXq16LPeYQLKLsrBYHo2
N/9CkZiWuE8SAWwIPCMV09J+jzdbEOu8iy/jds3YiDxpDOIh2n+auH0YKs+YX6Qc
lJ4GW6PnbVe2aWRd0x0c+JJVHEj10WWWp/oREMr4MQB2Nt1zlfqwBFZmih7gH6US
tfxApYLLbXHmKD4jT/DJ0Tpp3KPp+fzdGl9M5+H2htgjztPmW9+C5+pNoj/fGXZw
sAssO5xtSqwnO9MtuvjDbghsF4mwWSY+2iSCE8wnrBfIa3LvfZL+0wiJYDoYEXx5
VhLbQLRqUc62rqc1Fx3U2hSXdwMWAT/75XO2jsYW3NPIs2kzO+w2iSiZb2TUD9Ij
DUIqPHtY5ZfXoKypdTMU5qG1GuSTtEPjuncc+e7a6Smg7+ozcK+r+ZqhHV0XUqXH
Yl09g75j/Agg5GCQ5Hd99j6Rxgfq+IFy7dtjpqpHOo5ikp3WaMqikp9XKmvqHpfs
2icjTRghLAt3YXhrfjnA6oWRzTRaenND9kzZOYjQZro4zV0QYYjQQRdEbbfcR02g
4B0Yi1CxNxdIF7hV9z9uIaMujGHYM6hewt/U+0W/+lRJaANyhUaVRKVuk5taaBVc
454B9hOzfRdh6QkH4Kpbyi7xSNrKLxDQ95eTQcVHnsr6ldAwx4JAXq5NoOM3j0WF
R9Gx2Ooe0MG7xZsL9c0aREYeVqkpbVLmKWz0b+5fJ3A/Je+GTC7CtoGw31g48DVR
0JBIgE5wUAsUdtJWgWNV/L5mkRXQtqvWKlEHS/XcClpaxBanKy5kd1775MvMkoG3
6RlYrlj6gSD0CDWAMuLM399IS3GDjrPttYUJAdiDyORSrK+BKXPlZUp0QLEa7HvR
F88HOBpjB8Vni6vBMdcP0JO2zLfIR67sBIe7/A0MW27zB6PHVIxffLcooPHG4h78
AG0BSYqWhusfE1ipEHCvzS0yy7sJ/o5UgQDB1aD9DIMwhKGfMEoE+vCQ291rID5/
Gfhj2/KpdcOkDYKNdfTVxGAZphUn8QWuSenJvsAW7YriFVGy2zMFvbnXFXK8f2BI
eXUNJdoZHxQJRFNknjB4mnH4vUWx1b40t6zzHLXUPhhn+g7BigFPTAZHcpkVHGQC
canCXX0+GUrE0m5UFP0WUGM0xfZ9toQI00locVzh4Ar2Y4LklwBRqaWIYP6rRJA/
ysvxmu8OoDH7Z4CjSdJ8LlwzAz0OW5iEupHcYfX4L7JkGzIPOFGF9YqY9Ob+yrL0
/T4jBz1rLoGCG3T9BFUuZLDTfyzUp46Dw5ik/BusxTjgK+HGMPF/sqCcEZ9HZKDd
4D7OgPP7ecbYfHP/Ta79OWKoWp9TVZm030qMvcPL3QPLTKHLQQlTUoQyG2yiFlp9
BIrvmFxNjepFrroLeh4Ty603O1UFAzOCOJ8lMwtHCiNZmHTQ9CzWTwpJRe7fDkaU
gBYmgocAMNhmMLa6hXZjT5Lsn3Ffye1qIY7tHk/JuPctJTK+mB38s95r3IwchsOS
HC5rvuMR5ozWvCyw5ZHcR4CYzXWRObDqILnlXailu4J5sZHn1+RKCEIFYx3OFnDs
ALB2ZSdRj2e8ew6JhMeD0iw7bu4V0CKTPhQaE7i8C7Uxkcb8iEEbYeb4joWVF1vF
if/90yopNgfJCXdke0rFBqT6gulijZRQr0FvYrxWGSab7isHERWehlfaRyWIHLmL
dTMDSZvLaGeEh/AdlZgonDTC4+ey/bTVF20dmI5YZbvLa5lc54zVeHoxsOb/McDr
r5ujwDKT6ExEfh6MxlkejjGqnqm+PLQfFw0Ck+GcGifTcFK1AlE3dzzmKGFmH9p3
QKO7jxMOMxOG9RKdnDLNvpvYfKhwvvvOgrXzwwwgbZmGGn7hychMIpVQaTTt+zEY
Hy2R3u7cXMkFfOzI5dZj+2OEMK0w+rP7Q3Qvhw7xH9x08G1WNPEZJgVJxhNeqkOL
Rjsc+LJibIvn9MIjxjTyt18oI70RigDJW6OQv90ErSryQ2MNUpuwhrlLF99hK0G/
jPT0TQ8efRKSLEYx69543TYAofJ+Yp918lCTwX21GdkGi4A/cEfBAjI/vlUOviq7
hC58Xd0REe2azZ18uYUGcWBDk8zDseX5tFfIMbBzDRJMaAjvS++osOsKhFWrn/HA
`protect end_protected