`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10368 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
L2bRNdr1lLBT0eERw3vGlGkoZyuoLDUOvCJ2jqvihXqk6IY8v+AcUHT7wAASiZ2K
nWbc5cVruHgznFmT9e1wNrPMughMKbrFiHGdu8UbsOHH5oil65AjYlpd19xHoHJf
ThZxUrj4FfSyabqORh5+LZofqVQvInq0ZazNaeYjwI1OdiNaHRFAY4igP5pilfRW
1ooC8VX1YSMYht+lmcvfUe/WJko9r/iwMJWMypdRfO6bhdB7FMaBylbnsQ/CJ7RE
8akh6k60vIBmgSzvODCJ2jvTPhVZxLtoMKYHteA/K8lU3NpZwoxaSbBynzLC5+1Z
Wflh9H+MknX0F8j5MjiG/Ohpw/reYO8rEWlol1IY6KcJon40hAjXDoOs6u0sptAz
BRuzRg6ZpCBeKkG9uICX2n30QmfaANaa7FN4PPWlCzyqO6y4hJOEyTPy2anEl4e0
x92Yq7qFglggtfRSJI0nmZSRwj4tnS+LSRcBnfJd/mjhBE3IrG7Xaqs2AjCE+XOT
zoSeySrFMy0gefCV8oSee04Rt7nD6ptaoACTqTJr9uabI0U350rEeNy/di1jC0rK
tZt9cPPNhlbD1E8ARq+cA98yvZhL2i326/nGTMfcWzN20MRqj38XmWdzCg/aQnHB
rjPqW0jxC8y1ehJReyphbfQZUOhqM1r7QP2GqtFn5MEswyuaLZY469qefx6O5P8Z
xoMG4DedEh1bDmcqIlYuaOS4RP6EO0F/qDnrg9gAlBiVoOKBLmxPnZ+lLBpj49fc
srIhf+DNN/Perlq0Xcvi1WFPEfInRDfq+rMhXO88PMwv9em34UkmNeAb7682IF5B
Z2VM+7emaHWpURbOtnpIZdM6sWPzFTZT7wgUsqYDMn601iJjGc3iOw65LV+FOH1b
IxDe5rjI58c6KP2107pGwgVg/dJFqBOxAHQI/h6T0Zn7nD3hzT6rIVS2M/AleGpJ
GgeWofNpf5dZbhKzUeIo89MvC8eBIYshQF243wmFPk+Fntdcdgve4ljO1m7+ykH0
CDGS3OJrWnQ6P8GQUsfyUL4KaxOY6jNc3PcAYOm2JFWF5T3ZDmLykbJfPHh3L37I
6YyWRnfexWGScjj1dNPtujvft2hnla+8RlffQ1FRVYpmcaa6sk/mHc1gBy//4IEn
FWsLBuIWDEMZLUwTEFRVxhkdOsySgiCce/zHFdGmr6UEK6bBPyDvkInwIEL+Hq02
ke8T6m72zwOcnf7FOPcYtS1p1lhH4/wet8028VWPhKKKID5TOyDf9d+DEyu2C0W6
F8EwZTRDgN1r64dyABHjaO6B32OS+yHc6XCp1RQX1KUrkqxg8BmBbxQIqsrJQJIV
xr15J8oMj/zKnZpTOmfSzzofYsqhfana6DfGo8F7TXNC1qYB0cw0A0qJBisLSizi
Dj1rKcQDYzot6NWQrU82GgVO8+R+nnnTxFtagehkgK7/Q+zuPIeAC1N1sjj5UexR
yGffYJuS/mCuL5acW5OFxuiMPZMKK6ujA9IqEtI6tjJNOMyWYvb0s7MTE2y4Q6MU
G6HYfxfz42aGo1Lu54nnNjX7S7NWNAlql837ZJqyMexKRjSRcFG/b4SZZK4p9bFT
Ednl/vRC+BkmPIwXJiD2lx1qRkE26sV7UPZblIoA71LK3hzz+CBGRYo4/XCqYb43
LehY4D1Du7+W8wI9g4QAVmacrP+nCM17kqgpEXCAkudEBUW3a9D1Rk54HMYGLAXE
aO9IW5jlQP8hnAB8w2BCuOMbUaM+vIS/wPF2v3kjF/qPIoHbkPjCmvepNvrr2dHV
pgto0hYjRX9/uopDdbaIly0nFDp/6Q03wjDFy81mXYUnMVuYgXKpJepOtucLitN+
viCsj4QsbdjtxaBVyOCNZx+Nymf7QYfZlwSECYOJ5+NAS1ImxTSIZeGY5/ONdBzB
ZwiqOI5GZMbemsmY7m5d6p13X3DTEASQzFFMSvd4bPuKbf2CpIFO/hySHi7D+U83
4gNPLEDLQGEtU0uRjyfUQDyNUT1eNCggbKJIQRcfrbOpP79LFBO4TL2YH2QfS51S
+jk1ZFn6+uxA4GXO69o2KEIm+I1nInTFCjIKmbVI3b7vM6hs26qBwUYc5v7QgXHQ
w+HkMD9UY1pwCVlSY8Pvzn9hXJcE2TSF9CXK2X0gJI0BLxMu8qExScku0GhWRJxK
oEIGrx65c/A+36cKUU7OHqzWmXWA88rO2igfyBblaIAWDRPl+QibDoygBeR3zvJC
ozvG8gJVLwJmT/HVQm6MzRr32di/Ub9Li5eoT07RngkOgeo3fFw9AkfCvkJec0Hg
e6lRodLLPEQD62HQGvKemYuvSUsShkTo2f286agYSfNQI0jd8fvKTKFH2k3v08Vr
vq8JtYJOVClkVi+jU4nla/w8vHifsNWoFvUbg1xDIDnRwc/ZTQ6eeXQFclAur1h+
y51GTCbmSMd+kQAXw0A8skIPHu31UUki+iBLvFKUO9/MWgbqC3Bg+B9Rg7chQ2e9
9oFmqsKxlhNec8m1HIsT8wKg9riirS1Xxw9t2UqBs+wbXui0LrGkboQCfPIUQ0Yz
lcymDujv0mbcXskZilbXvqaWTymNpuKWV7G+wBW6IrxYbihfA4YldOMrrZd7qtsI
H4qJK7SjUdLjFxL4wsklHTL0zW0Az4KHnup8oP8x1mDwKKB250VIof4M/G9Br7c8
QkHXItY5Jb8lZGic5BOP3nXPXnWi7B+lGh/EAVXYujoP3pwh6GsbNme/PJPdr3LQ
RepbriGPuq0wlifAnEVhhOi+9NtnEn1kxN0OCO+sjqUbaQJC+i60ouCBFZels4vv
u7/cjlDWSl5e2m+trcdXhuPzzDAS4EUX7+lYtJikry/4htt21rwLswe4kgmEpMMI
No0OCcfGiRQFR+klcS4d5EWaWDy02XShebzAwcKixNc3ZbjdTL4j1ifv2W1S9QOO
VHTD2WSn+1FE8/SJFO5DF1ypGSx+wUljtBGHFhcEBM33u2z1HroQi2vKDBXxogl6
J28vZw7sWDWnZx/vMn985EyWkBWLAbqQ5LXpY/z3eKeTT0EQ5LZg/RXrXbhTNQU9
OIFEe4sOZ9quxpW0pd1etBa/ZIRGG7zwpQk8MY2p63EkHEaX4TaJ46x4seX4eSs2
HRLBhwUGCdq0yoDmg0wAN+MwcffdFiN/1lVrTYyeefcC1+NzI5MFBtZDxe81VqE1
HWk2Szr4yPv1ugEN0Q16O6eR0SOhoVAdvUEV0ElhwT/s6t+JLnDEL7ESF2zBFjES
4zMEoCyEs5JfG6RoJj2zRhgF1GfQ+6SHykB2kHZTy9BuRxnTDDCKt+QCZZeBD82M
I/Bm1fu9WDhZsxzumPrlHrOOKRPOunwGql4YtVTfQlY/EQLvPezeev6iOq2TVGbc
7/vokuFJfewUqyW7SE4Pn40qp6FwbRNFgVvDOCo9UZ1Yfv4xkgAEK5hhqDh9q7Ve
09KqQMs50beFIbUAVKHQoHomitTCVEwRm64DlB9uAddsxxtO0L9Pl9/TXwjzaSUY
EM7+dS5OcF2/ytZhNvqbB2/jMyvKoOLH+KES5dNZW/9lkcqw5NHYxEt4F56Y5zSL
ETjuha0sS3rSmij85Pz61Xfyr7q6fLy564Lyfr/sBrzac7A6yc6/srrZrMUXK/Zb
YowDott4QsE4T3HsbmhgliU/byJeXn6HxqIZGPPYYJvLldDYnxKdkWWxn7+jKtIQ
mLrZG9r+rC52PeMa4mHhEjezsEtrLJjYIncvcOa4UxcSeLd3YiDiZ1ab9onZm0wA
NSLvjATq6e44d67qduoswFzxYFm3lnOGtsl1V2Mldqdt/hXCvjbHKa/4+MoxAXyv
/pM34CKphOnaOFC+92LuMrulQb1/0rCIxOBf5ZHTh6zGPV+rng5/8ysuVasKpa6P
kwHjS2wK2gp5B8sQr3FqjemUtL1nPFmckNro3gFIAAL8gmhFgiuPxNGSLQIiHPot
KlpXOVcIJZAD51n8kRJe/Rl2jvngr465lz8nWam8F+uctfabTE+IlohyecGAOTMu
TFZjQ9joXgmi76iAxe/ZETVzM2x27OE11WDz3ptTqhUXxc+rqFvNdMsglQM4O/kW
Hd1ndMtKQ6z84DcUgmKZ5cucFCxt59u8kmNGc/3awfZZeGAY6Sb2oiPMO+JnpvDo
w4qiI5FBdO5Jt+69wP49MX6Q7EZlGtvF0Ya0+/1j9ZDtodO3b1B8Wesa/Ev5CbRN
zaZ3MV6HA4bmrKeb4Pp/UASXrhxqT43poPsfvxyr0zXGVM5JNVmgbTrfCDkzWUCc
ys7vuQzUinNgRrbX9pKPCeYKSmK5hba3CrqxSh+QNhRFWfyHmEdBj1aOcY24HrDG
3ZrSVGBpOR+noqzisu3Hd4kxFx4joa7nq3fMnOehj5umKkl6tRpjWKFyLlq2/Itx
cX+qzIqOWnvUiR06C3fDWeZP8tTU01HnmEsnA9AOViMVZ+ZiqhAYNxB0UhGWmmba
HyB3jA7loICz9HAfGpHSM+UtKB2k5MpBlWVWYRyljMef8wMC/fe5IsfmNHlHYWbf
43byfYtVqfCs0vpzsB+vulJP4VIL1Zqjew3zBCc5HFgENw+LozE0HoK0ENofOFql
qKHH7eexibNEZjkjW7kUnk6VYI/NVe10NuaHzclGHB7vMxSxMLPgowGiJZYMjPyT
/GXQODbnglRRvb9ofe4iB5AQYyj6wy60WpoN25xLzxWzRu6o6rMOayEmIDzrFjQH
a8NyKA5OEzgKaFyQWr3EDnOiesnAy3XFlz+23M+gj+RsXOWLG9T82RiBkJpBTr4M
kTX5Av3IS6Rn2NP2SU0NX1itfHFRDW7Mm+cOMkeWHIu+7f4CCWgs9MslSZekB94l
MxXBtjp3p52U22sx9SEqF3sjXJnFlt6+B6QCZwyjGyM7lwniM0T9/CSabmCKxR/P
3fHfTwy84Gr4AKU1di0a2+LTXH4BgbbzjqUkCJCq+GBpqFYose5hLXK4EV45xYqO
t79iNg8E29uGHVItit5guPTNuiq1mvHUBBed1myikgo8sWtUEMRl6ztRX5RqdZwS
DvKIdA202hh+8vbE01HJm9Yu33631NUBE7IhmdH94sjQpjBMq48P+o3svKpaSRzN
fKxNPFgcud+jZcvYBYFQKk1F6PLvAQL18co4b45JalfqSHtf78okXTnOOwxgADVY
x0he+POBbJFM9FKScx5xHoMHNPnE98afGuqvZXsvB+v1LjmjfoMmcBCxNvHOmvHz
g8zJ9QhUd0zxZojbsETkkaq1QXXZXUH80n81HTymJNferes2Vq2d9f6alz8WwnmV
4h8XXIEI+AqKSRl/0rttZBq1r3NO638aWXN0CJlPDfn9+V6hce0vMsiEfNxc8fqC
YgQVCNkE8h3AECpqJWvEkUBvIDbBsOcoFmndnI5C14bIXF3iEeW6/E7oWLhcfxgD
EmJYOMnru12dfZHwNIRLlgVQ8aK4OsYwVOzL+2L1PNIV/R26s5V2NLexb/4ajOFH
DtGTSkS1ZM2tYecJ8h0IRc4SvHhUHk3yMWOQC3FWxoIc34HuF+2wKlFLNVpEmTha
BuuuaH6IAy97treiTrEOojcVbb05kLfS+VdgSDVFHM/qj0dd9ZwlKFGJ+7Lys4N2
g/lbXaZahBlXJ7XhSaGZDiDHinzR1V2Y8a+gthMaYEyjVGoLgKK6rfR8/TZgPTZT
BDwtVwFlEjVgIqNGMSD6HiSyxueHyg51WmySdFbCJyXe3d927v+Qo8TlCO99iM6H
ht5VthhrQ3VPNvi7rIEmGOrODjSx33y1Jka9C0llzPoIVgtofwNbOZRIOcHgQDfj
137SeB9XCgxfvQ+W+gHsn6Vk9X3T15N0LV7Qq1wrcvnP8CG6rgerajopfAe7PHUl
U2Vo0PLV7xJfae7R3c7OYoW5c9LlJWBcaokU0LOubst9u59dXEkoFriAXPenhzRA
cRNetj5gTIc6N9EfX4g1gTn4692mJ96IcokuGwxG7NTr5EIuftyaGhdFvKgF7akm
0jI5/QKUNGFYvH2l4vrEemy3nwJZ9rxt5ci2KkvuXR33AwVt5NAsCocI6a81iLxO
BK5STzBef4xAtxXVSat4gpnY9DstgZQH/BiAjifExtsegfGKanpn8CQRc5f4ancG
m9fTbAlrbb5sI/jQaL8iGmcKOrYfjXofGr5bmrdJHYpkkU9e4fkTkpKcWj6i/M6O
5xWuGgcV/omyVuweulpSsHKJ++7mHVssBRj3QnmFLG4hCKrRbsUmkQUE/yrRdJ18
YZyGdMQWrPwhqRjdpq3h1euqmorwBSu3FkD4wg9vYx9ZObBmmpDsiUFML3JfSdwD
ZFQcnmv6dyFd8EK6hj5wQa8KAuy+fKefkoIhcVJf9qME9o6sQqWF3g7sgUsK+M8V
nqXGbwyCfk9yDzSw5Q4AK6hpwNnLwrLpwvb42wE/Nm+dAyDk6NRX0Uly/urziw9I
B/nE0ApwezX/pyq3rwMFukxBhIfof0imj6OuSsr7z3Sw7RXwBgPPaUPAKPHujZCR
ng+znge0VHHeCadgy8JFJwUj9LVNOi5zF3vzGOEoxqP3WrcnmV0b8x3OY35nWQxZ
NVkZxehyfr3kTfAeCo2EB6ioPy6gmVi8/uPknfK62czC+e9zhQA0cPEwGVrWRdLL
JuQM65gedq06ecj5CXd4M28CqpyVxLXKqsc7UPCOx0oXEZ/pK7muVhX83dBwcWmu
fdfJEu8TsfdCHHodKoBtnNz3EeK2mhW9+sW4u2711i/GRgCL7QEiTXBNSIZRjW+U
EI+E2Czt6fZYyD97bSGDfRRYot96Sb5k9OZpJjvWKo5jeplk0UDNMzWtFnQ+eoBd
LpLeQ+52Wz0yGq428JGg/Vh0Ia8+DKftCaGwD4XQl5GFpg1fFlCxDGH4LLvDZRi/
t5vb+05A3FzbGDtNg737kKpzFQ5HnQqerD0w2KATKR0faw36vGmMWg/qEM+4wPmB
3OAYYqvun0U4ZsyFU7aGejOmu9DnqxUYzaY4Rxpavc16Co7NL1yGusOYrk3Sk/QT
0wvLK5dMx2iClTAB0/RWhmeP8B39Yen6hKF5hISYIiWUSWxYljLo8eT9d2GkMGCS
ccLaIsTQW/zpR4EYz6jL1lLCguUFEzg9fAPwLbZlrZOrqmGKX1mVlhK9+iBMzjA7
eAYuDjYed8GAkPiO8CJC1WS98hJ+Dpmr1bN5/KfPjYIbyHgS+LmawkTADnnum7zY
xcj91dcg1dIPEGM0zXE/mhfz4s3COiJIkM2my70pBjSARM0oHL948kZJgUwLf7od
hz8U+ky7Bluh9bwbE9SpWorq42onl8G4m+LvmMZ/Y3UfmeD/XseJFC+gKxvYmpi6
zMehG/RzbhxoW85TR2ZtHWhiybvuL1BhVEto6Ir6s+FIPRWH1Cv4BPfIUILNMbOl
c4j717U/PAICl3a6tVffAhBjox/u1CpBvI/bCOs25nCsTkCNI5Mz3oPOfQvxChhq
K21XuheUlBttrNmq2jVQyXz/F7XrkR2HprkuE18NhRGvsruvvbSmMm4ZhW7j4heC
4QHTRPmP5amfbx9MEQlKMWwaYi7b1dDReK3QwgWxbAtizLggpr87uWmyo0MA+3uC
4GgrH2H4+6l85bLc6IdNbej0KCApkIRYLPxvh12O682Z82BCYEeXa4/T8y6tfabO
BpUBM3nsbwSYV0USLjjiby3Qgi41nfJm/1skfHr5EhtMDfI1NE27yeJRX3jwhuXb
BumMwzmSX528gmwGC1EZEFPf2SY4c2CjxMXnsHposrr6oLZYnQrmokWMOn1gmMNC
7po0+at7G0tnMBOyYpidkk9U2JPC8WjphPrUCh3eY4JhjJVW8gKUvnC4jYr4rbkn
8Uxj8nZDrPcejE+AN05nklcxP+01WbPgSPj727q2TXR+QDvgEVS+YUgh0L5mS5No
gicX/Kqj52/NVwXQVU84MczWURrn+GkwQtt9lbQ5oZ+jcIZ34tw7f0gQmXI6B2io
Q56cBOL8L0GMdFsEWnG1yh5ignnYpsspl2GKjq7RxoR8o6FKZFoe9POVPsjmhoWJ
g46KYpooat+qriJgAe+Ry/fwlStxuEv40fVVRc83e/62oG++e9zaHaEwRjCrI44M
OVD5aWfm19svcx/yXHzQb9YcmbCc8vD5vbfne4LI6ioZGB9hlMrjYGtp5We8VpSX
Rx+RloL6rksj2pYK0r3lSep49sRV8JwquShQ4DA2iHaM3Eya4BywbHqhB5O9rTcC
Aaj+rs32DOfnwB+CyNJqegWWk9GyKGrYtDoySqeYxt2JU2PxYV1xyeuqwgklXZB3
YTQZcLt2h7cBPYsMsBDpYzYuJ9Wt+lTs09+bhSNpdYJhJfgEDw3VVctHF6Krfcj8
Y+TLxaNCNoCSYk8MnUshDr/xyk6IsCsvvpL9gUf4lxRZwhLQXRHJNJxcz4mukXtT
69uCRziOJWSdWMYlNmx3h+ZHMdHqYR2UbM8f0OZBUSIIP46NFsOFaVdciX03CWsI
NA4iFhhAl+39R9Rm80H9KaIy+UXZc4l0wWneevg1yrQ1P/r3C4OKCf5MBNungRs/
BTDeGVqSFN53VqV4akfxo0PBqdrHemsVcdQsEtFy6wIzj6fR1JnQo5yyTJhW2Ux+
IxODJJVAjpAdrS14lBXA0NO7LhCF5EFVcFv8BIOVzV7XGBctzIl6aT5T3B0lNhh6
XXOUYWX93kv6GcKd3JEyqYogZ26dTBJOqPz4L4A/Pfv4VuZ0SXZXPuXuW/mIphRj
nCvRdMy4571qoEEzhPH73xHa03hciM+C//e8awH3T7JnemZ2TtNd7h9P3wD06Bbp
H9Fb2UYFRWtoyT/gnuFgeBJ19miWLF0yiqdLOXx0P+D/8t6YXJrs0hcRXdb7NcBW
2zB0vaHOxPWRVhYnptHp7vf496p2zy2rkWuft6LPSS/sluwP9RJHh0TB/ga9DuSB
/RWCN/1MJX3i90/xpBner0sP+bimSQzOXrgVmlYQCCyErJ01KNWEB7gBHfiOw0mE
AJidXQdx/+05HskTH6h5P7lrjLM0lK9oyKFCfxwenV+WJmmT7d5CHfeHLEyTrPb7
1Ie0LPSiV2dveLsEOJorEWBRKDsgcn6UA/yh58oqtQoce7Kw9UdfBAVWc48OEJzh
cE958BIAE1vH0SjR9nUv6aS0au1DS9MlDV2IiDGfHcIfl38ZOl9tUrbXM4APop53
1kmE0NAMiGN/vERWzSuKtXqY8c7nJRZ1RV+xsFvRLMxuAv4z5ntD387agpxInpo7
tX7dsI3Le5dAQsEcGyRoCXreRm80VuEW+4Jnq2yPyr9FYp0TqeET4dPV1w/rO5jv
hR2SQO1pUX3hzWKKewwb1BTdAaIRdO2fS5YE2IDWOTltUwiW9LggcBkowiTrsgsx
GacH1XEr664iRlICxCI8uVcu0LRLsaHQndBEAmH6io7Q7JJWHTnii0kAmaTnAwA7
+FGXT7e+qDHxqFoy7bmsNCEU8peOlBlQCDuo6V9+wjlo3Ltmhk7Y4+TTI15ti+8L
ot57rbQ+yNYg0fC5QoSG+ov4HXglR6QpH9C0llfwNxFYzbpYCT+P+VaYD7MIZpU0
S9EULHw8vGrVfh1gALWmaLPfSaVakj1HF/HH5AF6yM0h+wcARXeG59CY+2yKsEP7
unWmzp3oyPCMqE9qDWMt7ZDiGrD7sMoBc0kr6nOdXjzQgtGSVA+qWBzFaetOdzjw
TqGEbKqs52D2wtrP0GPakcLXY2t5k5juiHMDDLwerff+RL3hc4UgT//uVAfVhlNr
KB62Mdj4R83ABTSx7p4Neua3mxbNWiEijNrZL95Xye2GvAtGuBMOV+ur3HEeygUX
F+fSx/NX9sBRUJjvXqnfMgjjfn7gh0KIIwBcb+tvublU0dZPZ2hbixDRiYfFbsmk
TBlV4L3SFvhp5aZgdEMjJOm+kDRilZivOyUZwIQDEiQUi1ejVWSWBrpnsQCyb6M1
LtWMht5Rmq7iw/rB6JEgbDxPeN4DroTc4ZGy0XgWbvfNvJ/p86TBrweDAKDwzwnE
9B3tRiqQgYiv/hm92ofZrljHjV5/hbf430ukNBLQxUsSdngl0atrIhMMa+Wpd3WP
STlHUIFk3iYiuhNHn2mROaRLtA3jlga8YaOcPlzmmEFW6GyKa7HNDRkjwGTbsojW
ygWrzZOXWZuT1jTG1YQ6/GPuaHzyqoeTvFUjlcOxu60DbQLoiva9+KYvb3REIMPP
/ZOJACs/xtCT+qwzu21F0YBMWjf6uT9jUJz3Q/IEx+WViH0+bpysPLz2eRLCI//O
EUU/3CJ5/+5Nuq51Kh0XQRmBFg0QRhAxscXmgZN6n+xC9amuekSztKvL2MTtj+P0
3eNZC1KWSjgQN01t9CLToJLoMC1HhBDyTd100OrfqAmA8/m9cdj9FqAdVKPDEF/i
Hv4IwBD+HYD9XisWzerFwWWVmNcW0+3aoPNuSOJJIGCn18kERTYK+LE46zdJhdFn
zbjIapEP0d//aM+rZ5L1ZYNrYMAsv5lKmRpkWacaJp9uJ79f8D1+yPDgb8MU2l8u
IkONJUru1cFWfhrjQjveLWHgk0PJh5sdUhT+KEGkZT8Dy6DFy2VOsHM0I0nHK7iV
BNKU1A8uQ2BWQ759PjeaPkP4qjl+plla0ebHEFgZHxge+Bisyx120rk3Raxl+Y10
3SutXwvfCdeMA5rdGNPgwJTu/d6JfORbPxtfiQGhvJ0LDsS0Gxgjf+mXjh8rneT5
V/76/3qt0GbSZmLO8BKa3+0Norcn+TlzkWZ95HJme8HqAAFHTL9Ofaaqr0VVUoVI
icHd3QnwgZph0t6VvpmcPtupu2aJEvJ56OyGXlmdPn3GPAu/7UhRtXZu0kYMWeid
SUPLiNI6p711FqT7b7S0cRqC3YNeH4Td4jjeg/xttv1s05GbdZy057MdmRoYhsr0
9DJLE3IlgwPBWiktRnA+lsxHBXwR6uT6lTZe93oWil0s2X+dIKeATDzZIIwoDKaf
jA5ZXACEvcnMSqbWh91B2YiLHlwBua6EOJ8brDE365539A8AczKVmyYpTC2bWW/W
SwVH/KcG620I4xWCvw9+68uD2JYfT4BURnQm34nm3twiw+USbJtOKShshcYsvscR
/xQENAMEerFJEfRSTryifs0HgB8vexgz7cTedKSEwVog+VfAYGbhzpH+xfE1Muyt
gJXWQff1SaRJM7lEyNwKSSOEgd0hK6a6Jf6wtcBbf4yhYd3kObBpgPovzczR4ZWq
6RQbT9iVBCMVouBFCfN/bcIUMn4RTE4Rjf/YfIz8hMiEuSp0TkvSo4LOk5mS/Tnk
abeds1mSqFNhbeCF3r6fivnq5wG5uOvQKliEjOryoR44hFWkzRc/aTc5UjutW/vE
f8ERf2KMPDCts7IaxCBikhdzWASu10tmThWvXoG/uqedLt6iQC8xcGiVQVjOHimA
ZPVEju6sTneVqYJFsi61rPpikXssCpyjK2JqzbM6jwORbejjAIL8eCD87joDbejb
ZVHlagHDAvSMUPeLYji0u1dr8R8KJ7NfDY8B0Ke1fzpjQkBtXgeLFh0aGgXDUiL1
QsKOWCG2tFh9leIljzqx/nhIf5ptkcBPj4Ud8Trk4IwrAW/L//svN2lyH2pokGKO
o22oB+yeOJ4as8+rds3EBtuCmuXxs/ipQMerRkM3Pm/MRMbeDMslkfXO8XiZjlZQ
T9qQNxjI780QEe0aSJS2xk1wbRsslxfFpssRCFHs0Eu92qXgd2VQJYyZ149uGDwv
itHsfx+eCXXGcVJQH+2sXFmYRFblY7099f7IDU79sptG/JrV/0WuQUDDE2e+EzPV
/z9h/CQJf8YZklgupvwC4pJX9h4lofC0qgQhECYNQWEn4EdsBxIbr335F/c6nD7u
SQncsmxreeKWcX5hcl3hLiZoTHR2GpKRC0NcvjjDy9cny85z/tql4tc/ZbZ8tLS9
Q/lKylAoVVz63jjWwQxPzuRrNEXx+9KUlz5ESgyIXfx3u2LSu6T4jKE4+N2g2m+x
G189kB5nC+Iail1UUi7hg+NkD9W3kemjLt/E5jt6HhtU2gdYVhOYjCdC3WsVEGrB
5GeMuGwGsxI5N2nZUETAem1YIm2haF183AorGED68ExIX7tcxFI5FXJEGRLmILr6
NfNMZG2TWegLnYAD0gmW1K3BD1XOLA+EM5UuN+lFo9wcmFAkER0m8iCsUuh4bVdz
QVKuh+cT7XL426aRJf2kMq2jRvShpZR7gVcrQcxNoWpRTSp3Dwg/tWr+Imavb1jT
20b+YGAIr7CODVdDP80dXhmUqLcHufyNjds9/cy06MibgeiFHfUbQiCLojwi0Ips
Vy89et/RJsv2JR4QbD1cccIk63b702eKJ9gKUzX/CP41jZLIw/ud6yzh1UiD2sfY
W2Q96XV0GaeuLVL8X4+3d5u5JvnNz12KbRSgEk6Do3tJ8oI4zFnCI3zOofB/mQQG
347LJqPj+43oPYW5I0NTTsKMHlzpZXi4fjx4hBJvW/mOA/UDyN8DVL30lbQ2ColI
JwpFfuWL3fqkYAd/wzMaAexq6KOR0ljicmS9WIjHNhvvcyAO3kz7XrMeeGZlQDdP
ZQCkoSfZDROfX1HUHFFmd47MEaqgMvDL7vkwt6OB6UcJbofRWoxFzJJZVwFd/8EB
h3mWRsI65tD4Fi7rDOlTs0dNPJmVGLJmewfk5hGht9y4Nf4hkjBJpvO4Rxc8HBsV
W6kuxUBaUFQC/lXANe50SWjGde2wKkyfcxKlkL3J9fTw6xJSABo4bRiwSIpcQvpE
tPqCysqhd1sk/C6qinyZUMPN+M17ABEbgOwjaarus/PG5ksOSYSJReHKZxGiUMyb
EzKNzDoY63lVY2smUfV5Z8tGI2b784olhibOXWjpHzZ+VDAmefY2JstsFNpTOUaD
akFSAbcmyoqyH4iPQpmNmkchPqdJCDzujKF57PoP2GQpGF5qA06c9axPD9qH4Ukx
H5Xtb45XzTWBNlnx6IhFEJZTdoEBs4+NwiXEmLFdzLm3QTdK/+rltEwGw6upbAES
fRQbgSuyP2XWkeJRo6W8D0SvPlQeh8gSnMDYkQmN/lGHKXg1jK9emDCrQkY0fh+v
x1yVXXSVV+FQ7VE9x3Yxc6fOHnLAfot0B5HjoyltBxTremc0CaOaLTxCyTz01L8x
WV35zxYMK3YeOOv6sPzaLELB5q9k4hj6MPDPbzO0Au4bLc25DAbm6rQfnfPTd9kR
PEnSpFRZ1BJBfK6MVOaxG5oeeiCx1v2DsmeX+7S/RO6Z49fOfHQdAphf68/chBu1
klGhxnkXh/cEC4sHJcXSSW8N7TrJN9F2ht4ib+ONBBc8e9MaWUqdhiaMsqx/mzkf
9a6ya0nfvIvCBwESW2kfx08feUikhKLokZI3pqxsa8gEG4qWf2Cz9XC15+OwwKks
KgTTIqCIY3fBm4TiVmJigLAJ984XgkYQ86fLARDV9pzNgcb8uZSm7wC+iU8rAjIz
PYjlQhhPZPBfayTFmA2Rr3/R+xJfLNE7zdhDL4LJfUE1LXlaKsUJZVWsiy1QvRc1
tQ0NRP1bN6a2/KtZoCAmcslgRvn4ImtW/YNgHmuOqwcWzAECHrpJ/32Q4kXOaIJu
Z//svBcFBtI0lOxARhr0t8/Oqo7pyK1LMVb5kLGmuY2xwDluhs8IViEiueDFqmek
`protect end_protected