`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11232 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
ht7yt7qgZZej0S2R+oiVFU9Zfkm8FC86aMlFHVMxPeHiKluHnUpU9D7WO385UYRv
Uvk3wHUudwh5gMOvRQ/ifTuXk3cuEgvSWZ+YLJPXJ74rBIG69iYdLLzV4EtWBJs0
d6xnyfGA2MpQhITCa+Ei9jE2c47OQsmFnEAjnqvsS6dw8I8DZHSJYIpNzMHoJclI
DmGOk72to6ZR0khMcrql4vFdIrohplQ6Gjz17EG4X7skND5aHUj58WtXwjIhLXi5
f/djaq6Gc4rQiweh3x/2tBMLm4m17jfsgHnXW4vSYG2UVb46FTkvLid5AZm50g3x
ned/PZCjm4pzrV4fSYf7uw4hPRnuEw2y2/hXQw5RHbZtyHX0VHC4kvp214XVNXGf
xE8NsE40BhxqS23NMKkMirUtv3agJCe0JN9uBH8OuGXM3oYgsRU4ioSlEuVR07Tm
yB70Qx98S6bGD6iIiOTV2kZv+dDze7Kb2W5P1FHC0HqRokUnZg6wmGqmCV4R0fKm
5yQ6AbvAdi3WgbDTkrTdP/TtmCpKsKkVGKCv1mMWwYc0LlUe2A6TYDcLozTozjk1
roprlBdolyfZwbw5G2KB+YbEHdbiEsijtdTy7DUcagAQ1/lPpm1PYURhx6H8mAHw
OTFfmicdQC+ohtjOtMbm4H/cf7964II3h637gW/cuhw+SrOcC5OPH2VnAttt/T14
h3uJJOn/Rzh+glG4lR8gRtnboZDxNoytapPVt8rtkHFbwaEUDA8r9HjHnDz1sX4H
D6jEsZWYCjuHsx1Nkodl2N336r6tL/31dDqEnhYRikKwfOj9AOIh3l76aGnkcLxd
zIXBEaJ2K73e/Hl/xonGzP/3N6k0IG4VYh8gUhHycichXTO7MOV5i/4v06tc90GU
d+4A94nGSURpVSgz5jYItLBEq3HW8M/vJxbsoP8wO1K4LWrTpL76VNb8Q5sZLC/R
5jLPbas1PWC3Ru5rYD6SSPQkQSttfYJPji4O+5Hrbj+Q9FiSVsk6rnSi1SM8ttPx
5ysLwr/6+JzASVf8f+RDLzPQ/HRGwchp735brckjq/TCRh94tuHDS88mMCFas6Ii
rEPIVWDP2WQ+/gzRG+5ZrNtRzOmJmylVi7ndgpDDqFWc1PvVT5gJHb0q4EKa/boU
qSROPNRYG/UtrI6gWuYz0v+MJH6k6FJsY4EOYKs4+7AEko1HeZb5+jx7en45JjfV
lDfu/gLxk+/IbcJ5jwcAfTc0SvX9p7PjzAUnFguGWGQL4UQHabwQJqkHVjExKG3d
JC3jgnz2p8Y5VyrYdbe9a1nhA4/c/MQYOo6QG5UsU570HfN3YKbT2Uo3+6ra7zVF
Xelce9IziAMEbNff+28DN8EOwZCFrAQNiWfWqgo4vBynVCR48ImD1dfdFKz1P5Y5
P/QLdKxGi3CwgOdrYj6Jvkelb48TLCUjNpoI5x5ANszCoiBZJHDTs6H7GfZEp8td
4gMF009OPwkXK/0erzuS1RO+uc2OKfh+I0j/j86tT9xDbkc36ic1L349rCRuWSBr
DjaJHXXazKALTO/0YoIGb9QwbZugL1w+S11+pGvccmFfZM8UO/y81Ubvbu/5DCyW
mBtvXoMT6wznglcEdbejbwyxS/a0XJegmLDskcyeEpQ3OETeNfoeiann1Ri/3CLI
/UfkA2YbdnjBdqjwEo0SY3jboR+ZYqle8v0BAHDOTDxu9bow9NBOq6yDMeaZAD14
aPBnsgatmSvKnHl3LE7EdIFogc7C1X3eFSUD6rgHRU72qzMeROdEqND6OmjSx/g0
mePg8G3Il4rny79pUDnJ6i0WV8YebXfaQjXWgm6WG+GAlmw0+R8bK3ClaJY8ENhi
0a7/7mmsORz+5JOlSUnkCqT3yjWE20RzX4qEMA4QcPZmsAYNkEPWI/FLp9/7v1sw
tJxYk/tyXXTMr4x5WQqHy6APl0srZgc3pKc9dpuio6iF/8+eQpbM3WnquAxigWVp
42AJkw83rHxhdjhsogJtK31hicoPkQdFMY+i1wFa4Vw9QvCGfsmJWoVnFoA7yX6H
YZRu6fRgJIsqxAiwR/L5AkXs3OgLnYfKDsZECNI2ZFxuplYjn1t7yQk3tNJ9fwKu
M7rZ2Bp6RjLwc9zXIyWEzmo5RccRyyKJsmewnRZPRivB9VsYwbJ9q5xonAxRSnIz
AiLDCUIbzvwOM+hkKWunUisSMjqXHU0hF4qhOEzubqSomEuHtdBErbN4zOpcqTab
0Q7nU4z0mzvTiP27GpCGxDH1Kky/gSnrvWxSwGgbYnZVcfkBwnHehsfhqT/zll2F
ak34dbTxk0ZhtNPCb+ZMGuHNyilA0Df6zzBNtTN9TYJzQCKzTIvIqqF5TYcSczOp
ORtgrumH5goVserl1LiDOZC0iYY4k56bV5Ek4fo9XFnOD5BaUaXmOaiJrmDC1NxO
I3ssvbGU67lo7VqejQO28OSPLWctxTAueNXJ2sh3LcrDhLV5F8SI/3yd7zk3w5K8
AqlJORanD337N7pKhgtZk2ZTklYjeyW2kKCAIauDKvFDSUw/0XIm97oVh47CQCJr
se2EzXcOD5MF4ixP82YMR3c/spblUxasYxU302/TtQq3k+EQ5Pt6/2UNaAmtB3Lm
Np7wE+s6s2BiVfm5TtzSUstzbuccaiu5NgNB5lL3oNVMgH9ky+SWCZ3dFNiSiAS6
xklXaDwK9G8Htmm+LUr4Zh6TOWbVM4Xswko6dOOnm4DYcz34uv/5mZWukCIC6rZx
GL9LvkOBsHVPDrLLukb0cot5evPlrbjmN5naeOmQJy5ri/D7Kcaq4IRrNUzFGHjR
LoBGwdQ3Y88S3rCyxCpLDTN0JwSTMXepsncJ99etUhj6xDZ4985SdNO81Qh7u2aQ
8eOHNy92Bsdo8ErLasGyQ1of9bNNF+OmE7Trkmp2sDTIscW4aIgrC6SxpcehloDn
kYjVPJCvpzKfwslVnFiGC0i9oUM+jtdcDzEFCQS6CpA5PvY/c/IMq9O+CvJd+rRr
H86hNFrGUretuNsGa/vfai428M7dtV4vG3I8qRs0GvrbytfNm2ZGPQoqRmwx77zp
uVbGDgnAh1BlgeShTRA95b1LNxnQY3XiL0QwMNp9yImTS4Cqi4Rfjo39PnAs+c9x
zf750/dVUdmpRoJOcDPylGiuD5I+VXDdcwhrDyAJz4DD2FCzQq2H5x2vf+b+rAqq
TKWVrnhKxSjD3ZhpJi/41YW+nZuUIPlB/yq5FHD0/bgt8kFOPHdyE/LxM9+YzEZT
gzfCZfYdNEaXYpMDz5eQQILTUmtb7/hH9O0A8oY2l6NJzzAt6o0rmGw2zzNGadLX
6ySo7ZVrAGekaN0w/b9ePSyXM3XNsLyDiWgtsC2zKEepOfiWoJpVO0jRcsBvtnwp
FcHDJlGcUg78MCBnzTbD3+R5ivkAshSRdxmCJrdIMPQeHV4Fh5c7BZJD71Zx6R6S
LJF1Pqqf+oRpdHLHPJjjqvjDjFE3E+eIpXj6RSWShzZdOmL62rsI+w+Qkpaab4Y9
+pb+ifMR9wmh1Fj6LisQc0BI64Vrovyh2azksTcEhO0dR2oLcPUB86dt7CwghdQw
wa5sf0XsUFlTqy+B4WRZXbnMHNbByWNcJHhbGJ+qR6QUpP3Od5fWOdnCe08UMqB/
rtmcI9TnK5X7FcFDwRCcI998wuLLLcKDCW1ZuEJ44dLsqwPqP7h86A7XKvXVhvOS
qeB5TpFNdp0PgvaUXK9wT50IfMLn2PwQIcr7KXPpmtKdi4AN4HufCB44u77Vyc7o
P9Hmg/Df80Bn6cIv73DlERdZVqDy5Km92/c64IzRmLlvlrjKmQwzxA5N1aPHCxfl
TC5iPLj06l9Y2JCrEl+36FVhVwl9MR0lNVTKI9WWqUZCbEWDmbVtD4H2EuiLtN1p
6jfGycyyLPhSsjxIAvErCaWfRtC2i2fJtl/xH7G+ErC1dJiH7td1Yr5d2DVkuolw
CULZQHj4BVEALBr44z9mn6da0UTnqg368nQXxHtJZjgslGYb+rkqCS23fHbM1Opo
I2GLKdWB4MvbCxUneQz6jJ38aRWMvFurZsU/IZSTBCrNXAe11uNW0P56/+Pyj9dv
vStzeKdBAVzZBaFOTvLsL9Tf8ZiKnCn3tez94T/WxXPet3VXAWOnqH6EWDRQS1l3
12nxcO0Kiw8oVADoZjLCt5FnDLZwbifnLznkHPfQqpWB8sWyASs9WO9KBXDW+59c
sa6l4cb8uOv+NBbkxbSZYMC6MSl/ese7blj2mnoQEKFA/JbiMmJG+l/1C94mCxb3
gKlTwho7dFja/5gUcdOuwWIpgul/hNbSr8hO/mFluAAxLB8LeuyLYHbwgHSiKnLK
9ZPNKMGUBB38+8dC7XvL3cdN9N3LabApST6hfA0k+TOAoD5QkVBiZl7JbIr5I/EM
B+BJcXvV9T0d3OCOA0HlfFGuHlYFQZmKhHM6ru99Sqoi1Md6sBMRdNsPQ4ZF3Bzy
K2gphsr7ptDnWQ5du7e7vib0DLVGM6dXjVJncTj/lFqMUhO3zWIqa6d5Q0TH2ZoV
jYD59KhbEEmxGwSMMRBSqB5NiJFId4rrdHa3msD6zTctA5Rlyag3mebYUEFwQdzI
O2eT/r7X5F/dRhswrEWR/8MqGmgt45zVIx0hF7DLOhqmvOudNFwJbDtdpU647Ho3
XklJjfRoIqM0SVQFPAnzpytxd+gJkY4c0P8YcQ+JbZn5T7E4AiO059ZxPxfMe3sr
JRDA7D8dFD96AR1YhJTUtCJSnZQWRuM4DRltat5QvG029LSnGzVmH7Ejm2nx+cMR
49M4kD8zp9pa71oJjplI2Bw0Sv0532Vhd0DJEr0XmIbqiEfiTuEQM16sMVwLp60a
ZjlyyYrgx7et+PdOG3Hn5UKiGbuS8epQGUS/U5gx+Rfj6O/dFlV8BOnEVFLCevMP
j3CIAkl2DluWQ0IDNZEw36dzc1CO0Qt1JLf4xi6bAzIbJmf3jkKCZHH5n9XAkbmC
+o/uqGMn14e4352y93B4ftQU4fyC8YM5HcvaUIEJyxdNpQ5pe1ANdNSvnpIK9EnC
DDcu3MkuisxSR+1JDsKXw6yhKX1djKiVMCBoF68lhL3xDPVkdq8cPlawOvSpq07Y
U20sg6YJsGD7FyDUPbdibVkvVWyXE/ao49uP533kZ4nn/4rH+7/Q6yJGSUgjKYhm
0lSyirQyVYw0Fc1LAuSIi8LPBXzb16EfbdTv8GGrjbkevSuvX+0kyBtwTW8ggprQ
kmcetPJ9wNfl0Mwg1xAvfG/TS5afPmZtLBxG/6hbp4/8L0Fj3MIT2hExuPG2a0rF
lEJ8aTQQmaygHHztK5rgAGbLlg/sSqlSwBORN4Z0SLEZ2PWyVvUK8USEfkEv5lSh
o2Xw8KOSY2ho9pWPc2HYbREW5Wk96H8fNLTraRDkWfsYanQklaS8JyNcBtCEpkS9
6KTaSE4WZE4482LBB07rYs7oS+2wfk5zpUkN/Jx6XeKzP3ra0QcrL905c15+FUok
LOpk06QTTxW03XoS4tLmxDEmxuvvE+h0uL81vrhtRbhBQ+T8lhfpc7O30QWfsyAT
LGYQZKBPP8oJ/wR04M5ilyB5kVc9ifkNqP61aOE3mhs1uvneU26S+C2CG1sfDL0D
87a8JMXzWJkVADRxONX3lAAhHefHF5e8CgVSaebvT58c/aQPxSvkOVu2usn2MMrv
LRoqkRkxjKqqWDUgkn9nBsuR+bt1r6VqWlCEjq9a/MYaj11dj7LHUJVcqAPP1LFr
Km3wX+QwE/e0uKvib0ff/pu5BD7rTMbQYQ+JKk7h+ucZ2T/Sviocy/+kH64tzrvA
xOW3qupw2tLiXDDmFApwkl/j4ATNO6R8Aq2GAme5yjm79xN1mNA5uNuTIbeVKonI
zAg69O+2DWBOnvB1ykFmepaiI3wOUhsMaVaOAZiE2hNSDAIBOs8c1F+l2oyZOLa3
ZAB/cKJ3qbaX24rP1OIrv2kQeVNfvS4jlnPb/T2uNQXC2jb5nUC0YyCg459YQ7/G
3SHINVuOptEhiCxcX2RimDIvZWSIO/PquPaKikWt/mrGtSdVv0TOsyh6R0lXuvbU
fqF5dFaf8OJewM8bmGoph9LWuBNTdoZa6AbPr04ut5AuMmURBJ/Jp6u9WIQN3cuQ
eqaxdNdAdkB19qapicbxke03u6WzYHjYFnkNwHtNJ2zPK9bBioQ9WF2gHSkoMgp3
x1R/MR58Vb/48BYAYvdxqaIB4du7NnW9KzXB9/nIHYZlkRE+8krRNWAjIzDB0Xr9
RSmQYBKzrkuRH4H7iCJ3xzKQ782H19RjK17LkENRdSSHK9Amu/Iv7Sc06nGcR3ig
KznboPK2hKXkwqlvXX2VuV3A2h3HgOeiskfow6Vy3zuf1nVr47wIbA3zj6z2JOIp
GxmJ3miMa+nid+g6W3co9LpFVpuQVktvP0s9BGNRUlfDvdaI/IPmjQFtQnvmvtT1
tkhPXJapx3cKA86A67F8eWqfmQhkUUQFWuchH2vySOffDeHtKcJjEYXAP5JZQtpv
Iiv5ApCEgXz0NrBRDzgMeHyqos8Eu0/gHKwrIErrkahlnRHq8OZdn5V1ybUtxl9F
+6koitzyXDg0jOI4mPeuOeCfwSwpLWD4qoXTymnRzEVYsHYtC2hSlQ1PE+AbNeka
63yBre2Ct1rkQSobxt7nMn5Xtdhab9D5SxRRcj6+aTirq2L+F9Aun4eFa2lZ9rZu
0xBBJyMcVJKc8TrSCE6X4KG03u7szbhOfr7ivXhJofbhlHZEABBbSPIM36bYeOem
DdNZSWqutweNRwy3yLa8MNYOZUX8TDLuclEPP7YRQlTHCk3u4O553PqrQ/4bZASA
Bf8wxusS2SaUrNIb9i9isfLhUW4aoc3Vc6EW+Go8/o931ImzbV6yRIenotXK0X8i
CeQzPR3mqYx34RBS5V4LGxp0GSZwFX5Syp8G2r+G67vUqruCaJXgAqykySEY5D2R
e/9XDfLSsHeO57NZ7vZvf4asKW8j6NtJfzRQJfIbVp/R2sHS4LbsTC3+HpdTZDF+
1XUzloJKJ6D3RtLjNeV+I5rOGJglfCVaB+8R68FL3JzhYXiuAf4UgGbqa6Q8+3Ci
TEoz7mvXAikh65zQWM7u1Ojr9MVWcqAMVt+mmFrcDsVJJljxSaz1Me5kN+eMEIjd
7rEH7HBoBNHEs8S//Ob8cYb2sJpVubDMPoGTGssvbJ75hJNZaqdUyHDauGr9FydS
sBhY98zRrZBUJv4clxNPDNxF1muBwxEoOpd48Fj+hf4D4WhpRijPzIuZWx6fo5MC
aI6JYyjGD7rJLC7uLylRgdzlFP7Or6rlqM/n1JQNjzIZD09P06sYOZPlcMrPuWQK
lRl2BWpxCB8XohM0ijme+iabrCg8KplORK0gsd+ljKUHkPvk3mzAF4kJKIuwvVBX
0Ty0O6ZQhYd9OGM7Qaq8eZO/EuoxIFl6zRxPWD/vYkawYb6PUp4wu+B5hn88Im02
W/bc33ZSb3mGNdL/G6mBwfVvrBHatH1/ISBLuBmz4jURd1QS8tndEsRJCUkAscBM
eXIinZd1f1GMfnfMe6wOIiUbCAZLTTebI9/ZAh6GzwsNgGG/6MzPX5eqX9PSPcQx
jNAJOnuE4jXphbzmFsvQVh92YK38jF0F5qTE9QjuqvsndEuh4l0up01Wd4k8Dd1C
6F4i4z0QlSvilyPBZbTtFArAsYw8J+k6bRU8ewbAJgR5kbOJjf63zYgLIRLhdXse
R44rrhlOkq0+14IbOrSl57RD8Unc3zl7lp31H9YofFnfJX92CwDjwRNLF/G3nLES
u3zS9jPQtzXP4myn/IVXG/LXUY0qJPeiXrXjWP7R+pvIiX+ZSIeLOsA7TCn7YZjU
tDTM0r75PDFFSRwhoZ4aqwSG9in0F8itTMaEGa53Pf8w5B9RCARkyu8CwSVZgbq+
jhiTqclwT3gCTl2i/hneO4WdpPXTBu4o37Ge7915zibl3rFlsJhE6cwSJAjj3KdP
U6WdLKBOj1trcf8hD2rWWfiPqDtWWaro9ce4HqyS2gGgCGY/NGstdfJyqN07BWFe
tnwDY8vLhOxRKF2SG/tXCkcZxLBUDL5m8BqtHlZHfoy4MtkH+K6nlMNNbTNy0c8+
8XtARFvgDBgDYB68eRtAY+MxmsHi+2BdTJ6mCNkEjrLEEJOC2aSgMfW2lSJ8agWO
2r7D9ggDhikitu8r9oVpxI7XgE41kChl7M84uZXPQkNR4AXCRCC/jZGf7zbGfutc
IvNOEFVh2pv6sbnBS8uWRxYJky3yqhMHVLG6xvlBIWqPAlfT55HK5/qZA1bpZc5n
O5PNs929k7x27RQeqBU/qz4gjez10xXQquoIcbD9ASUkKjcMn+/HyFZRozGnhkC4
YL85l5fajFC89t4Em16SdjYUJGYYdpZR4EQc/sxzrgHeN3o3vwf1ku0/mIF4ORcA
NSzb3ZeePNu/sext2Nu0q2OCu5cjEwyfoqyh1n14gDx8I/UUoc9otWXa9W2NNZIl
BvJjlVNxh5JDNyF6r+e7LbgUPwoKDYPq7Zw1+abcfWn9XkgxqNpQ6Jy8o0aSAfsd
nN7+7N17MPrFYlqaV5SHKAteIXS7RH9STMLNoPPcVB2wup/GejhX+cRGP9g/hi3o
w1jv4HCa1o21hHfAfwLC+8iv2Nzo6lNQy5daWuwFX7qkaaYIR7cA9cLmTebkqvUd
/mEos1WlFgiKkPIvnOMpU7jjJlSMi0r9iT0O6zkJRNia6da6vWSwEcV7D1qKCX5S
BngG9p/+qDlGmHTRAKpbCFS3cMcMmYDqsRuhJ4UOGTzBcjVR9E5H06nS6D1sYOmv
svi634B6y4UprNiQUsWFC32li9xeFETax1LKRZvl2u6nbHw2SrQAJAv1y6IsqSre
rovtT1kBtDzLgmOq7h/vW1xPNPVk5Rp43f6VjJImTT7BqvTlwcuc+3S+YrfgsLf+
aZqw9hGoR9c1OzSMvZG1YxF/zPShSNL/MGRoIxE1NAcqgBmjMZd9Xa8praAOMdxf
VjomX5R8iga0oZRrxs7rYxBudhaaD8UjGeeHngUIpnd/a6cyJ91vunutCG6xtSdG
van4LHqKrWHfT5989u5Z0kTEBMBLSd59ekGFvNQPtbQxGdu1LGbN8WL11iM5emTj
F7Zau6BDdnfReT+sdYyPaOhRUQdoBXvyqqJQgUshFjru2w12MWbin5VjWH2LPgj8
8IxLkqD8Gd05Hlcge+gHMeCJWvbsRExPdfy3pgYzdg0GxUDL8qCNTdHu4VES5DLg
VuJS/mQooW82jFesdTObWw+vvqtSd41Mj4/SwzDDxudDtoOCW2pCdsy0V9B0hPzX
gLuWFFiv6rO7U1cqol7BIIQ7AO0SXKYCqdoiXgmnOsZKuvHmnx2qxsExu3iXIzYF
EpbIYrc7SoQBsgI58ibZD5MXbOXO2vQR4VsEMcf2pZTa8oPRqP0Axk/nGybG8ntm
V9xVLFNdpkjmBi4jZC+jb2mDuUn6xga+YK4IBOToIcTBrBYHwfrf8PcoThok/rTY
yo5e+ddWnPSXT6+D3SzRo50YrdFvG0qQbvFiZnlP0EI5gv3UFlZ87QcCjH+a1svz
54PUsfvbtWOm4XZylZOvkqO9nlbcyzfWVqtpCw0pFQIieLedWLzqYuIpaaOigigT
J6xY5FN28cmyHdk3j2MmS3awZTQPkhXBix+J877wYyT2xbnuT5BAwMvxaEvSjBZI
IyChyhKIG3h24DFHQlC33bdEiMSYYp+wkxZx/bagBmGtT2vmi+vgQ5EwTbFVw+KO
0LSGrxtGFVtcABjDno4l1jIZ1y/tnCaZUL/XcxGH7asLnrN8raQOCud4j821YmIi
fBje8zQmmULBKY0yCFwPrrSDnMqqGBKh8IK5dpDaS+Y/U1xrlJQgzO2KYYiE4FXz
0frklhosOjxM+wIX6ZwfAFDBLQHteI6yrqfmROvOWD2ePojdNKfKhkDh8Sv5YBJ/
hdi2iMuIVTHOR14Bfy5aFcF5GdKn21iX8VmlAriMgPX+TH3YiwutuooCdbl3we1P
qiKb/ciquAWJ/Zk0m3AxEtmCQI8GvWeaDYlgjVVcsZ5ZpW4CIVzvjVU7PKz/y9JU
GgTOQbenVH3D2FrGkWWmM4k1Wfo79Z5+HACuEkFrZ6EesWVTvA5OEa95M0RpxkY5
/Tyeg5W250i2nGBh9IM7sOpgNeg8ZX4izao155vjT60dDqSfLSvRGoi7NgJOx6aO
vTksTsRcHjyGL1Ef1VbXPqPLFmyAX+yhmTQMxmJ3PyBtivc2NnlKSoVRL6ClEI+Y
lTQfczFMKTBRyjOOPRGdNMh+6dp6B78yQM6FYfWQDaBXzE23Sxixcjo0EQIC/aBq
qD5TAE8vlaclttwHwCl7cn1P5ZyMDtH3WRb6/OmwRjj+gYYeioYjCFM8vUkACUe8
YIMOcNCu0mIS9cwqAme9VCJ7WnIbLB+o+OtaJL3lLQMCoDReFWzS9qcGHpdckC8e
uzwK82LSR/vSew8XVLigsxbtyoRyDj86jQV06qQUB8bqT+bxI7MkNjgq84lmFkf4
eWeX8Hd7OoVtHXb09fsGzh0Kmc59kK3mTH3sO+pTwKiOHiSpGNuQYZ5MMd01xm81
cYilBb4GmkryHcvDJKrb2gG2+0eTN9lGTKFaBOU6LmM3Ac7zMuKR8hgdjchfPXEi
2SMngoaj0iuNWH8iS84m2n7qkABN4JJ4Z1pSjC0cv049FIWKsqFfBMMLbmCGgczf
AVlim3ncY9LDwtJDVn/KI1TahoKrBa0nm2xhgUjT+GFz5Z++wbhA/MgN6stt4Vbx
85vyU87PhDNwKMoP6e2VT5kB5om//PncJuisJuwpV7d4Oyj+mFEQiSv9rkwgRwK1
g6uaU8xTgpj4T6D3gLtsT9phOABjd0ZAq2BsQX/54oNPS7gVnSdiPcheHm2HMy9Q
X/7evwOPP+JZY4FoBBnI+v8LpSJRdQZM+dMvcdCKhRfOJL5487ufP4cR+ktmhFpQ
VFabWnaUsu0HpD2MFVrTTxh9K53uKiWmRU7unK9eEqSp7nmhKcFPCx6pnEA9o3ye
9NFVBz6SYk0PrDdTOnSfxqYU6xYsxQHhszrUrU5dH5gTUjC2X3Qyyp9IiaISsEGK
RVrl09MTgmjyOee3DYhVPZOfWUQd8FkCDddyqrTe5Mou+2LG9chXfdAt6pqnEcOP
BiPdSiBwkR53IlRVUZ9yTBGi+Im30zwGh34kITDbOrJpJ/sG23oxlTyVCe5re8Zh
t/WelN3slHpeVx2iFSOo7FibH+Qm1sU6s5w6eUuKnTeWkw0Rqj1ymE1gnTdAzqQK
KolRxCq90nfaD8O+ekTr4gGd072/vhFrxvbVCYyy9ekwAkCB4Fra4hdLegB9j9z/
GixIp5CPL3UbGoruzawiyqi7s0ZWKrFSs3zQ4AEb7tqA8lhklcCOSzIP3Kt6ukWl
uIEwgcwy3cWgb1C5smlv15nCMVaAkW3glummLlF+vqFAsYp6A0Myssx3zmf8CKmT
WIf9+5+LQbCl2b4eaKaY6zP/u4uKaKMMZE5jRKSAqTYplDkJxRLjXCzTqKNyDSDJ
k1JYvYmBhAwxCTTIfXFQrcLzSGI0rIVaoGat4/wxe8JJGTEsGGqied0Z6ZlgODPc
+Tq7SoClVMhvXybDQyOx09FKjiP778wOR/DDWdJIqbPCXHI3sactCGnsmoN1wjwv
2rUjlV0Tn+K3a/1i5Pg5QkYtGdaZai+ZBrRRje0FgGq8ZICfFvtqAt5iySYgbNu2
CIGBukDvFsHNxUTaXIVVQZrXL5w2yDR+xiLSXCjWJ1EqPinKpwx4VwbryF8E/cme
NvnfFz2MWCBhqsjQwPCkhwC9wX2dsKMjaI4ldIlWpX2K0/7y/BVoNyrCImqT5Yu1
B2KR1RNvt/z+fp47s5yzoK8/k5dkGY+uG9odpM+0hMjXIWglvJxFqEqnvjsOkQQe
9apoUA31VS5f5JtmQiovW+yRyl0VdXw8WQqftQgngt5h4fJQuLzLDYw+he1yNihn
tgOdpCVUo9ew4O121zRcAP4uRnDKfzX0LiTuDT4fE6Mz1e7mAE5yx0Lyhb4WlfU6
Z1XWzvmUWxgxtZYKALSpkoMy1rcpeGf+p23vybgjfSOX0JA4NknioBf1++GOsXUU
sTeCe9Tf9/X1cWmzPi/88YxsnYJ8TwR87Ymzmva+aKWXiqcyunocGH3bfEj5WsQH
VBkaK+zx0wL7B25vV3iD82c8IJj0cZd6O0mXqrY43LO5gmuz0A0Qrd/KNL0/fRdz
ifEO1yDZLCxPwk8v+9P2DljMb95Q0WPd+HwfztVjG/WNSe1w6LvPPpFhMP0XW3pL
byFdrezUrygX87FNmiO54bfNo+xDRmvt0IN+gnPMpVlucQawwk5SoNb5K30OlSYH
vsC7uYA8Nt4H9bnJJTFsajPKS9hFIMbMKeAIdik/xU0fg0V4TTOCZk55/jU3Jyq7
eDcXHOkk6sfCC9UJtM+jxT06qIirj5ydyDLaagqnGK5cOilA+phKMVbiaupATbs0
mJyn8aAIe6+doKeVDGaqsLDDDR+4Pqu2uGvz2Mp+nv6J00yQIt1YmvMjBMzIMfEQ
vYYcHLVDsM5Ww04TAZtKl2PnySZKM5UgvQ6jycnpeHiVtr0CGQPiNxe9hOZQtTwl
Vcz4NvBWOKWwBB/WAocScU9bSdGkj+9ivUvRtTQNHdkOICSOqHQGI+0axhnOIg3g
zM9NO153DiQ6I3vBhRewV8afWdD695YN7nngEYLiU5ltNjUhRaK7uO1DHE5JXfmf
giY2MRRNy4NM4ZoRX5nvS6jCiqDdKESv/BCiTh/q/aPk6Qas5qsbnqEB8FBMzh+j
AC/xTj2shlRUlrQA57/zQyRmLPsU3Gy9F6S295WLY/OyttDNkjaCrlGUGj6Fdf4M
Uxa/G3C9R/12Z2XpmAkBMQu0j9sfk/bKJUp1G2JIw1z2O6Fgmf5nViklNup+zCvq
w/sNIKw+/zGCFCrV5k02x3EZCszfAuF6UxeHosNm90btMCstah8zhAlJR9U5pzuK
O8L7nhj7GAb5HcRn09xr8PEQHwoENAzwiQ+OILBM8mS81ZL51A3BT2h5jXfSdtip
0qTqBa0p9kA0ZcPefzuKUOOuMT6hUscxRLEf5LQPwjBNAuSQGVz2Dl+G0bODkf43
GbuYsFeTg/A4H1JVmYM7GjR1r7UWlQ9wMkbklfBmxhv/FLa3iHIU7g+dtKlPr3M0
JJNsHd4aoBZFPvFN+3ozalGEFj1PqKHL8HBg2GLVeA/C/EThxloFZ6kIolWfd5OT
O9nKRx6txct0NF2Ra3zp1LctsEE1BShN0affxiayQlbzwfyKUxliSQBOF1f0IfYw
8/m1OQDydJcyoej0ACp/p6Qdos3+teiP7/EEmCyElyygDdUs2WEnYisCl9x41yp9
dvzibOpr01X8S08qv5ymnRXZsgFED04Vz+Zr/FlOWMB+7a28VMZJsXOU2smguLRU
h6e/9MXngADRqRliVfiH2TzsbbG+YRFTF7/PQEfjTKDY509pFk7V5Lw3Tl3SCkXv
uS6KnCaqGB+RYfYY+5FkJsgv7oRZ/EsOj2g81w9+BxNp4glnnS2fIc7z6azSs4xJ
QCWm5jvGcxcogP59rBJDusXvrhHBVjAM/deb9E+0WDUEzOP4H2F2eHIeDZ8W5RVg
UnM+b7RJY92e3YwI5bcLr5xU7VBRUiidUoSzA1YQGNsYwyo4P9WPMaaP/syAW46Y
MJRGW8BWuJRUpghXKWNYNKoTZage3Uhpdg/wKQ6ZZZPAGPba+um9TBIoReslV3VJ
ntaadNL7nQlTQy8U+6hfOtmWHNJ0YDWUu4iIMsujOU3rUcrFbXYdwNUmv2dYn6lI
2vycgq12yzqZeIt7L3xrfLR6Aon8GAMr0RIT8z6CuOX8zACMfT57xOVIq9Z90r5m
BymIzPiE8l1485xF5GL0Ni5pRafnKKWrHwXAB7r+VnJFv1hMjKYRK0D2mA8hR5rj
Pmf759Fm2heJ3JxjTN6WO13x609vzjSyxpoLWPXlH74r2UlVT5G6Uj4pkeXtYeSF
MHeyyWaMyLNuThHvZu5RT2HVQkxpvTFkUHMYLWAH2QLQX1LtLhQ4B4575+G5j58n
q9ZUef7InCqGN47KdHX7Rq/XeNGnhx1jtIFOjEoNtVU5gve4Hgcmq+uPAaIgLq3k
bwJo0kKtm6X+8laaFc6LLe2U/4V5cw9XmF5FzWshu9YkOcyUe2pkGcfcwjvwaos+
p+334M02MxVgm+fW2D0JXM/HhlAu9QOLNB9TX2GRpFuNEOKVmzzwuc+BDXuJUXfy
QcSXZozxmzH/afASkUKk66FmzjbuK+1tl5cnsV0O1eO0RPGfNk6KpBmU9D22NFDR
w72Ie6mRiHupTek8X6Xmq8fVXlgWy/ZjH4ogrD2SFnFUrOoLMV+wn8SI7ZqqYpdz
FVT5VsRaJDWM56OZ+kD3p9FaCFq9FTeRu1NIJUXqBpFu3GNNOvDVWN4ZzOOpAUvR
/0eWqXa3xkcEVQvfUIxY7o/ikkkhPXHYItl5eDPDM4slzNtUc0GHkMdATHuqGbCo
NYsvVhbZyTxU0UqjdRcD7rImbjM1klUWHIH7tdT9BCM8LN92qVZoCmXxJS7Y18nO
cFvzp7nf5FOvONf3H+luA6+XGtn5xnEUdyKVq25uWlfbg4Mi4v3u9s+ygV8hgOKF
RMreNE1LwIhoo6yaKrIM3m80cHdcNVq83i22QkT44E8wTdWqCcSRdj1lairn42Vx
oeWBVq+uyGLmVieGmlL+0Dg55tx7PPjNy32E+VTSsnu+Y4aY08Ck9cGGfCSicWER
`protect end_protected