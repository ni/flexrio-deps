`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 19632 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRvSzIdqqwO5JLOHm2ufP7Er1fodAbHG0kpDIIj4Ba9VK
F4W01eowefxcxYxcjE1xNGJzw359TyO6XR2J2XH/Uq7Bur4R3JNQkNRc561sw494
rB19sKDcKwEWksqlMLi5A0rnpgt8hRjGFhtxwKDRDo8PZ6cJr9BNlMbK4GpRw94P
YqRYgTMs4x9fr3oe9xE1ejiUAm3lQ6AGcXQ5qlhaUT8Hyy29FG795wQSh2cKpD+K
A6pDVjz4rtDWdatnJqsB06FKQOmD4Kj0ush6MGPk/t/iWadjlGxAFsLsyVgnKUfU
PWLP4Or0tznOFUrbrMN0EMQKGUHMPyw3x6FoFrcw2GFuWlCT9hcQpi1Gr4Gl/Uqz
cuYZKQ7DQ0ZYdd2kpScWKaUfpoLrA0fTAeE6/FMKkNip/xun0Igc7qCFQqtyWOTj
W8EE67QWkQEPOtSH+uNzfJXB3WtnWsSI9WKHJ9TwNDGzL4J/GCIjDn0N38YMFLAz
RTLaUvHAKnwTvlYF88hH8a85vRwxU0+3OKQX/uvbXd2uZjMPg2nUU8BCgtYsYyJC
eFap6dXSRxBLXyTH5cHieKrQVyuOEakDnxFaFqZ+qS6FLSFFlFHhrto5z8KdpjuO
eUpQs2AJyzrcdffBYrwwDuw+t0juekF4bSp7PI1AwE2c73KL2/6YM9J5YWWoAhMm
O6G5wTXzkTNDHi7lRmNdG5xO/yYCNl/LkF8uN4/a4y8OyfIaBIp9ARclT2tiS1Si
jyaGy/IwX6hopdtf9gSM24+pc+0b8YV+yFG6JAEKbLj679oCs6r67CR606YKvMHg
fjY9Ze7SFFvkyOa/bed7xInnbL9WaEiNSOGWBtItiEYfDIz5SLYZFfkV8j84O+v3
kzSI950CyAU2a3t6gFxSIuMagYXqWEECEMIdOAlD7oicJMyRr6PojIrUwA8DoaDf
ciyXZ1GVbJvj4WMCaiHUpuZKTlwY+lcsYnaKnkPhdcr0pWIHMq+EaDSrJbBRoGLm
dZQRPuInY7ewjib0uUQkTG1tWD+jfy5X94uphC1n2FHVnzysLvV6pv/jpozPIlSR
8pQ5N5bvBQWgu7MSNL64usHMvNWFsJpA2Ck/+zPOST9D4EICXpQ4ChLueu6HYdeA
GZ/pwpvreEZSGkf/oT9RwLVP22yyOG67es/BOxBbk5IGlqmWdy0xS61nfKdWyM12
hjIv3StL5nim2ah57am/QRy694DMwCqz8rtfhsiHUPwLxvtr2XoNDFy0cNvWSlYv
9b4LuFcBb03q/hpzf++bMggfNEGQBX7Frpdi3HWN8Hs8i5rlg4kyH0P1Tvi+be4x
3aaXhV+Il6HAPI6anVqfXa+L+i3WYs47psTzYAdajKLtKe8AeXjI2HTG3GEMKPsi
tH5h6O87eLeCJFY7DtM3NrDAhSRlDbYuo8Y7noEftD4wUDtsUkkupbgN5QdOgscT
z5OT4V81/xRWgSNJC8sgIU5VsMmdwVE+OojpiISX9V7kZYDHBcf6AVGv5/dmP3XM
++e9gE0gVQNqtzR7jwwdybAaT8p3nsEjU0yLnSczX4VpY+MiASbuFbMhojpm+4DT
a6zWy4UtSXFOGCmQh5zZA2nZvJk7+IqyOCBayIhYw8stRJ8VrbowCK+QhcZ6PM2K
Hm6ImhPVg1SO1Om60IEu6/COLfVZDUVLPoOFjh+yzc37k5GZ41tMnX1wsLt25xWV
cLjfl2CYHd0fcAqpKoTB5VnF5dA4/D4ll6mLI9ufM7N9kiKOtbUk127UW/4p0vlx
pGYBb/Evr+qFujjB2yW7Xj8qbGAreI/mb04TgiVm7RqDRfoVRQD95kmddv1YJa2x
gyEQVx0W8UYhyWrPj+9NZ6HnRP/V2wpq7ep+Lv53qQlarJTV1g02piX0/NH9kmMT
lMEaPxhNLQnXxpRxhf3RX3uYfIQkH2cTRq8HSlttTdWEegiXV6xIkULJXBle2+f7
278uro1H3GQrtfxFUaHBk2LdLKGOJ0cMJvMsrpzzmzVoBF8oaw5NNvU+0Asi29wF
GDEtha4zNn3Lgj4DNWP9PzxIGAE7ZrNObd8tso2vv/oQnuakIMa8CiVa8ml9KaTB
C5zUug9uCTAVGQV+Seay94ZPX32peSw7XLvGszY4erRrMjya3+FRuRLr27sfDfC8
nydAVC2Lkkapt4mYvcQ7kGeBkJy5tJydTuyhQEXaus8WJ7pyM1DQOZ7t+d5M14v5
N6yVuh+T5UMNb4hoTurOmC+y78SZ0SBRTRoONfjQwPWwlvihsUi0RbWR1g0q6e9x
DUJ7e7s2G34IZzavd6JiA1C0iQ7J+gGriFfOLojuBZ+BF5zUyTgyRRUAGmIbggdg
WNN7PhLXtAr+7EzaDP46Lf5oI7AtJn4eshu9UHKo8lMn9GcJgR5I17Xn7uBYeEdX
Tc+IJxRHq4JhwL4D52BMNrYbT8Oie7cXW4Vr3PNyNIuM66EC+v3ojp91LmCFJEpR
BI2LFB/CAX3BVFOJq8dKEcMlogSBAU4D49yGCtREoPOO6z+ukHUGjwZm9cVydVNM
VdWRB+QPVPz4bRVVbP0JuvUhfUeo0wY+r8zkGzjK+FRJy+O+cwTC2GKgzhug4GR3
nmE3rNAR9rXkTS+qqcfKcElAn5lv67c4mK0+QAMAgv0sfbxkLuP3rbGCgOZN+qCz
Kf1eyhYNj2579ZNxM8IvC6Usg6eJ4mfPx6oia421qcHkqw/Ib2GBUdtcGBxmUXHX
fCbhm11hVCc2so+MUD4lr7bwxhI4tpD1fHW0ANZWoxUbgae3A8ENe714fbWWD3eb
T5HcYL+1wB0srNDHa/GVUxG7CO9ALWcEeGAwaMMoPo92sfdXMEFFnBW/Y4PxqKFi
4J4RA7Ocw5LVTHPMi59f5Shbbh1a5vPAg1AlH+PGWxzsHHnGnKBsMCId0f+LNbU4
qzdIm3EhiS7Vl8PK/EM46AwrZ5AiN3RpgwyQ0lQ9R0QlaPzkhHvj+Y31UXmLRQGp
onHZUBQhORuYoy2YsItYMRLaXiO5k1UV3GFR06br8rjOCxGCo7m4r0LwUtSIhEkZ
LIimCIWQQTyHUzHXKs4WlmBgUxw1rI/yZPCmBz+dkfeA9gM3nrVYE1rSwxB/55Z6
bFBDcGEGibpgBFemx2BMlvL+WzX1gcC0WBeO4wt1YE5r5Oe8qtzS9pnMYYtVXg5G
aZOOja5Qo63+mVqiA/h+sThegR9QHFdOzBJ1e/hQNPNLVf08ExCz4sT3zF6b+csE
QDCeq3Prctjqb8RfZYeFz3qGg/5ZCGsDdhWbkAUOFJ88CUM/CZEBCVz9WLXeoIQS
fWAHeH8scT/nkzDqva+jt/cjjO7J0dD26EjSoPkOPrb9jV0skOyeSXznWpnXf+Vy
O+XklHP0H1AeVFRFmE2X82RGK2sSgMC1VNXO7TMed6MnViEsFWJRS51DuIwKoC0b
slq5w4n1G9xqTmtNil6/Fj7WOfBqP32GfQGPkHTQRoj/1pBqFboyCqnfLGnBaAvH
YPuwnFI6+FQyUQ8WvzYBB3LP2BaW9vmCNUpyd5ge2mBHIarAij4gs+QQ7xLJvYr1
LNhdyS07IWWjPyCGlJjni7md10cUnSKxzblGBpI+Y8BG8N+nBSdiwJ9AuR+vXNww
9yn5qXKT6Nu7DFcLhlDDdeo3fpz2iaLdk0EVCKd9iDSDORXcjec0ZVD8uKWIscbY
gMRh2kSp0HzxFXFklvfh27SJowF0NQ4tRkwe4jRm0ro1nX9jRV6ifQrWbQDjV0G/
qsifIVyTWDkkIFomuH4+FrlcbgRtYSjm9klKDhqaDKCaKHIB5X0VPzBJKbSg/bIs
LibnnD2hXt4GLFTPvgdUVOajJGrXtIs27hhp4OpWxMlEeCrga39xnK8t+eImeN0c
aoID3geXc96Jwp+p2rnkF7+IQvuxNIBvWQnfbzItB8K91MkoNopn6bVNMboebFe9
A6uW5bEBhG+2ROW79Rj9dZlh9r+8Yd1lLQDItFGOc6Y/OZUopibBdoDpS+u6OwhF
7x8W3qKzg9sPD0sLwiBRF7r8tBphvO76P6nNkL4QkrWsVlRjg9uLscpkniOjpPH2
9uyGlgfWZ73Wy8wg28HNUf2N/ltKWLtS0TqrD5QE1xdKeFCJvhHV8qAsPpPsqvw6
u9M5NtodnbBH5dTp96QKS/Bd9/VBfxDT3+Nh5jBFmqXwKlVzHsm6TtQJSdf1XAN1
BoiOtd8Px2xpbkT0SIQV+VAq65pq924RPQmtFhkEfjsfCK4E/TBFwLAVHJusogrO
mCl8yfLw0Y4yIoeVTzZLjEtR22X/7Q9OW7rw0sqU0bYxUJWDeozs0ifWpEDmKELZ
uE/P88JMln4OwPiohgeiQZOEBdKbIbDyPPnh2TZqMb8WmoUOaTej/NmmuG5Szj4i
916oVPxXr4/HJBKmrEU1aZFbGulo4paPQi98BMlIs7Ihg9aX7SumFRRAL5ndpxlx
+itbD1IX+PD0Q1KQ8MpSItEI3pB4dme/DlvgNzVYtsw6p2GS0/I1fqBxNGNgDt8z
Av/EVnM59vhAFLUrfya0pi7AI3/RZDqyZmtkxfevqOnQq5uklThAzT5a+qvk5PBC
GfFUd1vPixg2Da8lvo6zjyfieh9b+3d/3ek3oS9FZB7BFsNSdh4HbxKizYUKKZlp
w7TYIXl9MiHfLXveh60W2H188KXK/jff65/9t6y9KxE/jbTas/HkDzDKfimTnVLU
gK7oV5cUF/eIx8hWjRVWDI6GadbeKUVAQFj/YHK4tAvK/VKmu+ssFL/tiGxu7Kyb
RuH5UUFRsQ5eEY+je9eTZFTjboY1z/YuXpV5VgP0TlcowVTsy3KDSH5M/XQ7juvH
JwD/JoFLbUBdQx0WxjQWyEcIbop3xC7s+TlUaeXvD62kAwZxEI8ht/hzbKy/N89I
5+Q9KqWntuvGBrkBw2a8FwFzD8zNdcP3YmLD5R+VEOmSNt6WSNjdsHaa6nKnmmSv
U0x9q/xE4eByiHuXnO5wALxNd2Aq+Om4lZ8Te0RpXveo4eiFmK2rRpiBb2308Zcj
CBTXZj4ysJ63624Y9B8O4wuZ9zoka7LJ+eoC6UNfme++4ddBfM/VlYE3G4ugpu/0
lMh/1rd033CfacS2/LKZGWXYPhCjwaUhGB9QZk8o7TXKIN2BqQB6elVpQuqbEQwr
GgIDcG5GzJQKx/DRENwUclTYiOO03dBVqxq4ByWUraZMk3prJCAH0dv8/rHgs8tT
LE5wRCHGDZNQ+t2o24ALlehbk6o7vBhJRDskB+iA/yzQf3QRb5NvAvBthJt6zwLo
EgP6ZfNqtWhXXr5dVhH7+maxJ8a5dKY7x+tlPPRcEShlOYYHKXxg5Ge3KzJn2ae9
hxgYXgWp77WvXMBLK7foBdJMcpCK4+hzdOMU0iNvLDnHs/oXKQEQnWhFRL35IQ5B
oCl9R8JHRKgH5hVHBtXIX3WhydWcrWAXqs/5OB854KvWVkc2bY/uBqDAr3ZlxySo
zOQK/06uNYWieEL43l6st52TZJkhPZvbo7YDwtiSTiOHMcv/F1RdYMjOO+6XEbpb
OwDchmUz9vsdnn23ijpO4Jap+9R/x9jbuPyPwKXvrsb6WxxgGa6xcRzkJLYtZr4e
EC8IIByxQSb12kkpINoZQSiv08dVEqAxqhqIi8bklcX4aT/vakGjSnK2KbrKyGvJ
ubbh1N6WlBHEeFhgYvdqj7o1yPkgW8r/bDA3n4dDfwjbINNYJGrJWfggpTC+TxfL
5BsxOeq65kw7+hL2CXptqYTpcH4acXsQsV77YEAql9DI1RcRzdcGBR8yai4cpR1Z
IQPFrwbCDDjQuTtFDZU7LmHbqtGYIBj3gtmRnne+T5sc4HbKlzTuFavBThBobv+S
q8w6mWBJSOpckdyKbjB162PQsrSAtYPwWqnSh83N/k8DrfcP2D9MIZzliC4P+2VH
hz/gM8TJRrJ+AzEtY3LXaMaCjemzh09du8/9QpHgrxaip1yy4v+9GxItMeBS5xcW
lGV2mgILi2yOeQh+Z+UeQXgRiSq+zyDBkcCDXwMwLX4YCswznCs5P2pU4qIHTkyT
J0sXbSrsZZUKB3i8yW1fILmhNq5WQila5Vv+lhtFHar5m2PRLSKcGnzwCWP6XFLc
2tMZzWEWB70xRNIi1Sx9KQj5gK6a3qatNQDV1nmg427ey7t5kws8PFQ2RtPKksWk
FjMvi9In9V7mcNtdASYlB3jIh26tpqV0Hqs76ZEv+NYskGr1BViqzTTuCRiLpKJx
8x/PslPr9f3zVYYtFZTaTYay4cD81sJWNtS1TgLb+BhUVNDT6UWw6AJvBz0dwl2Z
x0CitlJa+5+ysyt7UP8D9/YF2Xcb9584Lxt7CpI4KrFCjqDLbNk7IkVO2wo/ESSb
+2T7shjQ63NpnU6KV5iyrg02FIlpd5piC9H5uyf7an28pQz3kX6Cn02UOWUMdvqG
BOxI+Fq0B2fLjNv5jPaabBCd2X57P9/YRx0lKCfme02AJhirO+atAJ24Otaz+LOq
zaU3koXnVYmw9O4B285QugoyUPFR/ZZVgqn4PuAkbfcIojArdw8VMx31/8Cd5kSs
0IzMmjImN37b0MBiFSVt7QGVEBF/N4P+5T6mMWtcVqw38jQYDdrl7Jr8ELLMtJXh
uzL9KpGEc5UsykXwIzOQQZA1unsFgAEU97RX71DtVpTPbzm80Yhz5bz0JSH+eM6r
EccaHeyuJI8jfi3SqAZ642xJlRCz5Pf3cAIl5y1WyKXWIA6BF8/Ukhe/sDA8738e
n6ieYeFV/fpsF0uPYAlKZ11Eh0MHz2kTZI0iRtxKSWvwkXzJuRbSZcvjT1gC74A+
DVaQVK+6l7NUoAOM4M1mAU058pd/HaEycYwnpE/gai5Bbl07x12+x+YQr9DT8fMI
KOzZq+zy+Wlt4QMCnBS3xaUqYLPTLr0CXalpunQrPDZgA37G0uCCyn0MYEhjfTn3
qnzW4xAhPD5ezrvuwZrU5TZP26owHpDzOhmzYCfGY5/LPwMeqfgPG1Ni8zvIOgfO
0fLNSkwHGgfzwLpKnghE2ys9hM42Pxae2MjTyofFvys5qi8gvaNLUc67L/e6tLHW
mGOAXCaEEbo28v19laM2w3UvTZlJh4+HDrPWJVX3SgC1P26oPYVuTyRvYW2HfH/1
DXg55eOVkHjCMw9HKvxhWuEa0k/f9jOYkj2ZuUxDTQhSXKVJ1ONs9pwGbxYB+nTR
7rpRwoP3oURX7ozssF29zuOTuYDjhZGTxolfczQEL3D6lokobZDPKV3p54SI5McC
TmGbo/+MiZySTYYSAKmeRiSlUr3IKucgS/F6YM+/nvGnpEJim1ifls2TBfnrbVt5
IBXidHe/RHAWXb09DvD/X9qnHXmjGVmz3wnxtaYQoXQ5FG6gYjxUzLLtcU+iKOBl
9B1xLJudL/l37mw8f7zNgdu0B+CbORquSEONwtVU2kdeShLdEDq73hB883tVsyv1
fGOV/w5KHL8egjMp7niZPZR911aT6DufQYxbEXeZyQj/YesqrlTBVVXZZbo5CiBa
bHooUoTSofSf7/GIx8UX/iAtESt3t3lZJqqDxTfZs4GUimvjemH/KnfFcYAkKXLZ
WOg0I9VOw6vOt4aNE3lwG2ag+SHfTM9kYFI3UM2yvboKBpAjGD1bedCvvcsEXbB7
Fcv9dlwQeKJpMWKrlaWBYjGp6JEBLJx0Kmgl455oEhYUxgiigqL+Ri1ja7ku6IWF
5SIePV1eEa4X7gpXA9cNnfpnBvE8TwSLohZSLozDaAEo7pMQEvNWgLizMNwTRm4a
OUWCplVBLElAi3aPse7IFTWpetR84RKBZ1+t991XRy6Gb1wJaVMo6qnUxAFvqpkK
IsqUWk782pv8S4unvZOtSNg0NIpJV0UpbVfwUYQg37OfchmB9Z0Wnkk6FNq7jk1z
ZPmm2SGL0DFVKoOQEfGKlRj7X8nF+hj6tbwVKxE2dUIEvbTvFNoWPxczvBYN6GGo
3z6Mde1Z+wjRdx+BcBu+2ilVSKJouXFhUuV2vP8rGYX6KaBYamZH+fLxvrc/LmKX
RsbzdE32go/9FCVNMRCMZfR34hr/W3grYlTtxO7pDFjafljJBM3VImk39q/y5D5O
5DH+zDNmR+FVH8yHq1D6LbA2oWYlIDC0dtM/3y5HGOQVY3pFFy+KZQmIV8n0A1ng
OCp2/IG9LC4fzRzAnr8EgIDDBXw4+u6vrkPUXSmfqZznhOE84zHcD16IBYd1GaQe
dvajIr89qLPC7Zzbebd/IPzJ2iOC1QTVHGeyVlWjYCx6ijqN7UPHOqtp79l2kbSd
G4kP7t14VN67vo+Que5EQhd7Jv4st71R8TduhArLKEeiJFdHbbKHgL8UJQMr3h0f
f6GS8jsjwHmcgb7q/iTVTr/FUiFKUtMMT3iPRN707886Hg8SLJ5WwIPMP/wOYXYh
V2fCRgjdLSYH4008qC06GhL7rlWdvzuuKqIAnM2jrJ0UE1Ej65dSV2h1yfH9vCWY
tHo6mNe6iAKGIZNp7d+svpO1ylgoOp12B8ULyLLe7aECr37gZfz9rulEOXIgMAxR
e8UE8Hk378Wsu7wY/qkK/Cc9Lf7z9ZdpVkh7u/pazB/Ew3vjqq1/MhKOnUEX4XFw
T75QDY1UmD+S/2YLsqQZr91VLZb05haIjB0KfqCQwPG4TdlXlm56ZA2haL6Bpok1
vsv4tMtMnZIpCOreavN5i6E2g6fKYQCQuwRNReCJUlUq7qn8FYpw8NRS75ioKROp
98MSvRkwH5IjflbNi/BEIpoJSELv7pdoyJz/A5xjTibVIHOEnWkLIXiiM+jZzkoz
bTsSUSwXsfPHogT9X6GxJEHmaw2tN9ZeEWE7gYM9OP+WrWzkzMmZT5PXIR2VqIKt
8iBxphiunZUYL3UBCmmZTKwI4twI/8E5TW7F5WY1RSmzOhdRjRkWOFJi5STgAVet
h8s0v1I3SKSa9sJE3vYHtvYbPjY1jXVvlY0PohbB9NQAS7rcopbBhcs5vjaoAN82
j27j5ofIiBn0TQRukDmWf79YvCdJINXx4mLIYtHR8tqBBS1A8ixjMU21I91HBayz
54UvcBC0StBz3SdVwDd5Hp+DVYlfoWxg2ac4mR/Og150jEY1grYFoH5v38q4kgv1
WpdcQXWaG+bFDY3qOd5nejGxVe/Q4sDr86rtguaVkPRWEv0QYCtnnykR4qZE9xIX
zgnNMQiDRxINepe1xGwpC6LhnDqP1+HNbMt/20Tw6jx3d6ZYkcs54sWfObvfHlFj
odATjp4CPKT/Qupa1dhv4yYr38e2Q/CvAGDtSdzKzMuQrVgskdtuNuLF0F0DIXqJ
zqFLNxKtubcIHFkUB/Akr30BjGewDi6iV2UK2Yu/2wKVG+t5oEO77bqHrvLKQS73
IEPcuGloLaKBCQlX4OmHp7km3tN5tkDwBVvqlWyWyOPSj7CLdIiGkHz5iL5yTHFO
w2LD8g/xCvT/m8z/FTNv6cbQxN0QDYXAp/fuUkFZmiopQErs4ZsUD8UFA3wzvLzM
EJwut7gBa4KgFLOuYRKtvP/wsaja0qHg6XLcLeUvLDMxaOLxl9Kemkf5zRj1g5qg
fw0EYBeVVfYFkRbscruLlKT+5m1xYVpl5y58bczb78q++a3n1owZJxLlh3FmTw2N
Mb87awI/3jKvIrmszEijQ72k9EvqA7S9KSPogBeTjXB1USCE+EwJOX7CIeQtYWWT
5A9t/zs9Bzl/WP/llxN6tKo9WkqM066Z305jmAIRuhWdCPS22TLiW/2nTzUZysJS
CASnQ66nKx2liDdQCZ75JYSfJEdMYOomxq8/HzYYZyhlPExHAznUcc4A+O3z3MZ0
avw4uF1y9/sCc+l1OnsgKjDElUcQU4JByIvRr6L0mwlTdF1v/6vNIE+BFKd8K0Wu
t/gS6QksRpuHTMrNDECdJzQt8snHXfF2u0Wu+Mmm25pOFT8kzei3b7RY+eTsinUz
B+OebRbsSSW5G2/LtmdEr1k05+rJcbhjP6iZcGO/8FPko01K3XSwrD4Z/Flv7oxm
5lLN2sBlKPxEZ83+ewWgl9ztX8Ltm14SVRFuuK1Ycu99ZL6EWz/9CZqIQxsUk0ab
iz5PWz6F4Iyh05ttieTrtkcePDqxwXNRViCOV4HHI3PPzYcbJib53msMi/qOKvhz
72RVmTQCAmqJLLwW8UoClUPlp3uCTVX7MXN8O+Y6FUfBK73TQJwLDPk1KIaZQQXr
oUuR1+eOwi6Mm4EsPvyMvUk+Ng+OR3sCZPOfPSf5VtNj29AyPXy7qxaIbpc7AsrB
9fMc2OKTfd1AK14/OLt6EZuBT8mM8Zpqpg5aFqKvYgGEZ20FVN0Tgljj3D9I/KHw
IMOy/sfV7kalncUyvKLq4K/EHM21XGznEvTk0ZFE74Imfz551YkaZbm9K5W9xKBh
qZ95bRgNAXJ0Bw7oJGRWQmNK9yw5LvxcrDwOx/UP0UTI9F/HtFRfqSsasXU6YWoP
gI0RU0Jtmulqz5acHmrf1ZPPin9+oh2i6qpKR6km4tq+CZ1y/NP88rsCza3b+RWn
sI9Ue4zWm09mumklQ3qlk1l9YP0LqY0k7sZyEXwKzmgOeMr0hCtIHoMCCNArEsTk
TBTmyzfYSougOoc/6I4jVMEHmLKJYBktJpgj7/UC0MgB4wSgnPFM4gC7ouX5PAXO
OXpYFoKO6Pu0ZmQZpuRSRFgujkGxz6EBtd0cwS7uVZo/8P+P9Q/3U/ppPgPeNGmh
Cm4VnEDRRyPDbNbAXz4OVMtM/Zip+Dr5o+Nw74sJ4t4I5PHW4UpMyiFOU+g1gyy0
4qwj5iD0I0MpfIA3OfA3l8YbhXFwHEOzWmTShNG669SeeTeKD0laPpXr/TNshXLH
W5//OpNS3p+S/2o2S2LAmZa1buW+BWSEcn4Eva2BP6EcxdmYIpYuAAy53Y4zZEb/
HJuN6lO6atbEzwyxNkdMESwSdvZk3YmJIcogoTK3OLbqhG+ZEX3AzqfO9hW5LFGs
wGetXNuQH0fRWujU0/TfA8FdCXSwbb5ioO1ulsfSQCy9t48dJrVjd3UhrbfUhpq5
zSD39KyjIK4vD0a/ApSp6t34ZmkFGwEcn0NyWvg71U7hYGcwU3+zk1CdlgNgKjZX
sS0wV9wZ7zOQosDL2uAVbJ5xJfCnYHRulKBBFR3IS70+2lZtNSoh0PoJDzNjwsau
QZelKmuFsKLX1Z2X5hKnZ4Pz2BFBnoGZd/niHQJXEqt6FtAOB5pi4BKdD/Z9cDCY
+xCmpQL4iSVYHlLeXGOhkhsWfuVs2n+WBoX0nNv3qrfay4C0Une9cZR82WhQ0qRL
6WcQFSHGVQoRMEth2ZRYMBObDeyBMxii5lGDveaFjzEY2xim1Jix6yXM61BAgnbZ
zFI5b1UjZzmRHDUIfxvGhsCBndBGJZ9h3kCY4vclUxZpRtMnFxygQ48dYHeo2cB8
GYcWTSWQ16/KLHrvDxKGlbwVoK91t5qKocFanKXYMBrPyz6ooPUf+IMOX8vjb11u
mP7FzZxI9Hs7DIV7ZrdBNGy2TCkfndtY8Ah1Nn+av4E3IcoZpUYpphwVa+CfR7hs
g4xdnqgW9/DwbrfMaJHWPy18LpLDHqznZhzByN5QLHBTi/wJtjqPUqqBVEJba73Z
i7xm7Wktgd5MtvSlOcmIJIJmiVE6rI0SfSqxwILaXXCtjAW7MtnS6R3nUG1pp+PR
oetl1ZVaWr8F57ntUFQpy2PMnskwbpaxfjDf2eDTCqi5LHWBFMmjG73rK/UVlr3I
vUA+LN0UZN6DwenbHjgk90Yp/9ivf+YVSzqabaN0ZXlbt8L8AZKfUh240Qugeduo
J6jhbunvOJzdQ6aATt0+PGqh/b/2GJQbkdvz14lJKgLKLRbk4Lr8hj6viP5iWc57
UnXFn50O2tzd7c9OShl/T75pOJLMY11flYG7KgGzT6O9BB16hoD1a101yA+gitOZ
/isjWAmhleCCrhG9dNSFfrGCIROHB91khK627taPOE1/RPcU1m9eZ3WDNDnEvBDp
Mmja3xG4F4ET59BjOhwQDOgVh5smPlfShQSvT93J+mybm3dGVvRDgFrWfXyvell+
XGoVwB6fClGitjvdr/wFu5Y7CVH9+H4f4LQJ8yAxPzFr5Zo486Fbc0Ks1s6Bol7J
2tSJey4kq6IIo+siJLPYsIBuMPS4KkuvelNrUlRBw0Gsb7hWITU4J0EzEtLK7Hux
nxeG84yr95cEiZGfUd89FgMQmVBftvHCtdIeUZHH/3S86NsnheQjsdNYzK9r0V7i
RnPpg7I0AHri/yFQSlQFsySl1XuQUMUy3lqGv6fDgmoIPeZR3yJo7TfipY/j/wn2
ORngGWl8vpO8p268JKyxza1tSxtFh/Yv1syfx4hisuBPpLS2WMFrd8FCri7qn27F
ZiPIeWS/9WUEQsBpMSfbA6jo7YEmplRXUg/bNDIefN7Ku1CGkE9pF+svaFmGEBCe
yPtCq2MXASNnQRnDgszmG5qgzTxCpYbvN5XXYRjFuSB/cnNo8k9cm8wINnvGpwjf
73oq0IRjqd/3hXPJgOvHvjz3qMUaBFX1FC+FNggarYbT/TUYe/UqgwHc7kD5PSV6
IzmNps/ihLK7/PJiH1oWC0H4AgQgzfCWVrpdOqZlJQGVPAf6DxtgcfRIf1C5WGbQ
BrdAn60fwiR6r+5To1qTNburhbe2q+nvmLrkjmdCuyM16Y8fAWnUXa1feYjVtWfH
YquLYHA2d0hQRWTjV8fk0g08BicIGhW8n35jgAT+lZrTag2i6Qv2pscwsQv2IpiB
TeEbLesqqm/FEb8/Ho/qt8VzODozn4BFq8FQuKJzjnXJtZUa96KoPKeX1PC4Et0/
c2I3srZBF7Dk4qFTFbyY0p3wxP/8FfQALPikuaVoXBy6lLvwlFaRfyZMro08rT48
w3fGCV4C6d+fHOcQYGf2GHnIU3B5SM+D1EaTj6QGY1OGhOlulQQzgBfUi7wNQySi
VU+YlacI+aYvCH3Ia2RRLMnvgKasE2YpcFZv+ooPE/CzUhmRSp0ZL6ZGVQqgr8R7
1d+h1D/zA0a/0yvZuo58uB2bpb2g3pY4AcCqLIrErqEnlHTpa+Qwm8vIOMAnaULw
ev4iC18sSA7QGvz29SOY9y6cFqnx739mvoG+jTxbppFEaX8i+KvDeNas6pgONo1C
Dq3ndyv5T4HfAJRG2RkrIVzUokjcVPoDt4Dp8/H7jviVbqhwFHARC/d5llMELLNl
u9d1nVSyC1s8JCpExr2CbEIS1aF7jsZIpVGTBASQSFVrj9IwG2BTScbthV7j1Ru/
STF//44iuzOiLaf4Dk3c1lDnnPKdyVt3o7Sg7rEhLE42Qq/pV0S8VxHw27/9gDsk
G+ZOivL0zacNny3a3U6EsTaEl2VV5QS7LTE9wSbx/q3KJ34NBJ2DGqQA+sAO/NhF
J4UCk07z9Rh4Bk00zNNj36Cro8gj7hnqe2mmTE100jh6vZp8U7KDjI5doSx0Hwbs
5Ok7v+4GLDneGfV69q25iG2dt55AEYnX6ariy9XNtke/k3V0nOAQ7ywgqwaUQnff
6BNZcr7Dk1pOLBjcEfzzNiRf0HlJdIuOn7rxDfRSNa5ApidYQx96wSGccYNUCis1
eyQKGwK7M0lAzFO5YvKN6aGO5ll9+iow8IfuXGfOeCxZdBtOHJiRw6CShIb7rmNb
DSee1+iTRbr09dsydmmilV/awA2ggKGQJ5Urw0nhaB1VCtjOsCm5hGzoOg/zIax/
WeMKJth3s5apQaJ4AlXnE2E8Ig75cMdjLYYenYR/bEmR8T4V43TSJYrk45wdqL/c
NCVykL22u5zczvasUA4qJq5cVC6RhjcIhKM2jq6KMGFqaOKmltFt+oGLUiKv9aUo
6mKb0TLZYLaY5CxvBX+ab0XnX7gNlZzeEvCbY3EuEbSzSH7Li+E45k6xlk7drAaH
8eGr6PomkB0egU8s6a50eRrUPIENWYOT2RjQaTNy73AlOgPMNHT3k0xYSVDaPcTu
Sa6PW6YGKLn0oh8f4mjor9eVrZ/nN5byooUREw5ji00nkqMy05VIaYl5qiiY3Qph
7f5NvnOUHj1Uwr4RT6vae9JbL72OGXf0BdCIwuVrX4aNWTBLIe+TPVi+sEt9cSAz
gEtaLZ35IlN+XcdpUHie9LHiITeg/irwmUW/wy6UClgt9WkBNCNZIxfx5l0M1rcZ
8uqcv3id8Rt2pBnXFsVuyK5bc4liHyGknxKMKbrBXbLYkznhjmtt7CUuTHaJbYTF
UeU/ZCrgBvHmbosIw0YlNCuocnvwZdrQjV4QsUTV/zH2EJK76KHBU7jYu5j+aLJd
5ij788yeLGt8gu1Q5wQV1d5pJm5vAB6W2uWcGVKO2ETKhp8slkiyfdz+/mE/L68B
XXZNAMnDS1l8mEum2uvQ+DrUFWZx/2wfGnufS/BoJrPM+UARX7SsLmg+yEDpHB42
j2IZx2HMD6ArnO4xHm6yASIH6tv7VG60Bg88yluJGMl60PPc/bH5TC6mCozVYJjS
dd+zrKX77cyAVGrgHStOrouYPlGYlPW3PcEOEwAzIm+9Bafv+5ZL7kBnR2qLbW0s
cgaGfRgtBkjg6gcDpN0QPuUDyXZQcHGx3i5uwALI/P1eRWDcjJP/LU9+GJx64f+C
+3X8x4x4s+0PMISOu1SLuCsQnFpLGmPgYRmv3cWztj3Jd4jFUno3oH5qGXa1I0uU
6EKVVbvD9ZoXQxZqwxfOpwkusFEZuQ38KA2tM5Pu9hMfsjQkkCJ0AUHMugxfOQBJ
hoME4Tbe5csvFi5q84xVMGz6TzfWIdFe72ySS5Ws09T7B1bJXbJQz4aikL4i1fb/
ma/YYLZObzMHffccvb55SsbanLXpZy9LAtmq0g1bNAsPhdvvxS3FUOue0f/C0To/
gGrQRJqtSDIUVq/9TQNEI4OU5KDs4U63Ri2QjnJGRnt1OCh6UiYh9NRtp4nxd5zU
/v5jJZ/VoNnDTNZTTh6Hh+efi1NSWyNvDeq7qg2D66MPCkwG1mByZxgJIDbTuLCF
7MNQZROEdHbaBAzzsdOmr1RT+Q8ktLaBmVZ7nD9XuSpLxS6kCeZMATx2Pf5XSnIC
BWKCATUhdsXFF9MY62vXw0wAwfjRSExXB6LKExdo9801Xhy7lmj0zcWmcFjDooU2
7I5d9IKJHrV1qHGlqBYr1IEwPDSkr6FzuMgzH24q7rMnMv2tR5Vx89jxa+o6apR4
7ISJpkZUo44NnLAsMzUuUcs4+Z1edIAIgN9AhzOeW7mItL6SLSYY9MMq7me24LQ2
ZayvvyaHFJaorJZPKU26rcBrAOqWif+kU7EM7YF4xHU5IUMx1qQ9mzHFYjtDGRUZ
UIKNNOoGWspD3DPJZ26vEdDQUN1ckWh9m0QJ+l5Erm0oHYMIINcB0JcxTxVc9lJA
eYtTrUqtZwRlK9uv2eYr/w6PVe8/OUNGsntP960tAX5qEXakLGOkaqS5UHzXJ2g4
cVlJru9kHBGswcDSeo+PBHTOwvjOLtNFn/hSu53tyAuWpzdLvMJmPU1G+lUiUbnl
l2owjQOfj3k0dO4jrR8Z+w84qgx+cEtRxkNgzIcg/H5NyvOziur7bqhjIOIMyE9m
avp6xGS4/tIz86Zrt+ERB6IK+vGhzjqamO5DNXBnar6wpQe87CPIWiEN04uwv4GX
dU1XDuSq7igtN23HZ7R5CmRU6pyBThuI0qddYCJGExaj+yNFZdrFdAYczElmM1zW
afKgtpJo3w7Pu73AIdgoq+TOkSaymGkYJVs8+CsIKhUsYPMWcrKwiMUGKnmUUwrk
vbOxHfxlOGyMXZimM+CYgcY/cpR7Mw2cthZprATWY7p3dWfKH8yER8BPCNB7Jn44
0X2Xv5R+8j2knDC38xN6ntStCX3S4wB4ee29JAW+JimrNvH/QdNsQfzs2bOxIlOF
oB5SDGZs+K2y6nvpejUOXTkbBJ3F2aACvw8Nfq0P2I/XziGpJZNUYpef1Ux+cbX7
H4y6SF6ZJmI1e6+wnxZQW5DSCYkkWz9ZFKmPC+d34Ux/oZEu1poMlzVceSZLMhzE
upKC3ypYUva9xyGdDdK49w2LeseZpUsXsFbgUFpuw0FPUyzrXEGGojWi6r2x1zBv
R13qFJ7kLP3Lt4dnM0jM9m22k9x3h09b5tagHvkPEUnlxdf8+Q2Wt38dZQy8JEkN
ckLtNOOXASrlBGchyoEdXXsudDdlpH+vqkMBqyepkb98WfiiaYcvB1dhwahZzfca
EZA3bXG9DINg1z+PmU7f/xVGVEWNUKW41tSwJyety2PVb5lRETtc9Gy2U4mAx+E0
0+c9pvUqzQxNolhbncXJChqnCBWl7qtIAJskQB6NWRSGUczpajeYo8gABU/lPNMO
SGPdUEnTldQEYW2HTObaS63ktWReJT1acb7e9Q/5GDsCWsKs6R1mkDKWSw/YRpDF
TkEC3CAUHBm6lu2StW/D5bHAwntpCCcULTVslT+JLHeLnWXLL7QA0jde6O/p9+TT
xrdIMbk3QAJ2NQ06kxzUgWiibNq7JatOU+AD/yflVPiPzBeYDBOnuUMSAofWGqlI
MKoKlvb3IebqQJmBOEgpp4/owzfEZg7gjo7qhO4ikbzd6j+qr/C7JdJ1YbD0uay2
KTX1Mp+6jHpCMc2+E5Sv6d89jzLr3MPPShzUpuN8DMtFZHO/BURJVoIWVR3uquwl
IOyjus9d7Ud1APtWQVLVDXv9FXXhqsYonTcw5MfsETbs4wUwDi7P0zhSoJ4+04AL
MU5a12vw7ZdDq6/H54rXJc2axWB/MCzrKHpHIHuyvNtQHQ4nqcdAWtFSkwgedTDL
ADILE3ZVQR8Ztt/IeZ8Us961GSKLBW2iUtEWJGlsCpODbEEZATcqQWxOKJrcPr0H
dkPjO0ANMdXO+MX5bDe913PkdUYKAcvCI9vZcn3pUplmecWjmCEUF9TVsWyRoO9D
u0eFWnrco4hV8m9jOCveEc1VB+jmlqqOCfk81xKw4Y+3SgAZN+Vuig6xCkleWgtM
E3Kuk6IcPLZNhdsExLT6uCk4FgGVEwafzr2IP98lei1oKcq2s/5Hmqq6i8BCGyg1
AlEImDT393SqUOCZ8nUaw6aInU0o4q1euJBqQfgmMNe4RmRI44Dd2xbHsJTU9eEn
V4zmeGetJuR11W4DgRPjWvFaVi9wcbNxSUW2cqpCWJ2BlzLoizc0Q28VBGb0fABe
DXjy8PoDkse2Qc5AtNnGYe3rFhbnBZU3TKvsAaLyj7ceXnWrzuDwkrLQLLA0GN73
5Krs7ZvWlOJ7iXDX+k150TPdUrP/Io6wsceWIj+yLBXcLg0+XGUda/VXinaAP9Vb
Tyfs28VYLIVtk2sucAPtEfYWkbw+JibU8P8afxx/0iVEnF/ssOlM2QuN2E0feKCX
FUYqF9oIL6PlxHoSMkryZw9Yxbieqw1KQIEGRrdl+TkG6wFbWS4WVBNPIuQmn8Tf
JBs9uYduI//AhyqJlqi2yY5OcPVISbIXmmRchxqq4+TCEhsWdjiDkhFtik3dBy3v
B69u/X7WIHW0fm2pjNa2lqZvlwg/0Nv2WO24poivE1Re4vNm3DQzgepNDoGqrCUw
ZsOfj6dcRIthD7Sg314tfon7q4HSI9xErIYdkcEyhIiCd31t3sS+MQLHqpqOVG6q
Z1g/zBNxGE+iFYKr/mIE8jEAWqB9HFD/kIZmgeDKi41YlYF2aE0lMJMNsfvbDI4M
pJXhG4k9ibwMRAKioWbn3cLWce9w1PRvtiG8dw34sk4ztFYL0yiVN30h0v79OGrH
mU3pIzgrHw2YTcs/b5FdE4ht1YVupBTWlFQ8sEbyIcRx0lXZWQeeiEnApmVqwVVL
6c3t0u36BUQZdheTw3r6ubcERkj48hOd8t1iBlSowOudH8M7QhpomZXv7i+RcFLr
sKDW3osssHewBqDmnXYKpAs4Xp6LWN1V1qx6Fqq4Ip2maBZ8Fwkj5gAY7A4oQkRe
tlHoTXjqePvCX+n8+FrB6Pa9MyP1LsMgldopdWnpEs4IatIigHLgibm2ILXqN8GG
BEAuWEd62r9QCWBgdtSy4CX9UmYmm9jHsHI+b5J9bUo2d7VuV9Kb52vG05c4/7nV
DQsPE/1oTLSeeu/0nvOAKWv+gnf/TRibZXtjw/ueJWeRFwnLNdeMddMpXiKo9YnE
9w326GXxPRgM7n2xmsFHP8Pi1qjd2MhCSPeJYRjZFiU3CD4c32aDfp+hcKbvj+f+
pA2RvB0Qy5fKw1utzTQrajULBMqx3vfurEUOfnmNtFNnLbcs5LhFeJOcu6/NYcxG
x2F+cC5zCBx2hOdUrmWq8sEh1YQGHOkbA1AwhE4dYsHEVyurLRsEw8ERtz5WMPSg
W9lyGHnoY4ESjmsgb9OlOA9800C36JoLuSaLDZvs1+RJVesEeMP8FhG8X7PZNAuf
LxbxUxQox9znvx/jes68VVTU8YYi85cIs/GWsn7+El5ptJZR7SQs5pbSENM6nS2Z
od3ikZ2E4lPK5C7wyJ5ZLntiUAU6V1GbcxLeNsx/ZtiMxfMV9XvcNGdBgscsUXpy
tB8H1agnSnfvNwWFbI56G6SKHpCEZ+VtAElVlIgyeDxgDyW42Klrmmf076bVPdZz
S9EvDn6GPxTrSJMPWSyRBhR0aExqpiWmTDUIb6ie6mPWgBakOz0yExaHLRXiwL4Z
7TKqUzZHjblswDHeeQcOQFb4g+4xHsIx7utOeRYHwRvKyL4Acjm5kdQ45mhMT0l7
W3sAGYVNyMRJlPJtyblEGzFNAuV5Ow3Cagoh9VQ1GMvP69NB/cP8/MCHHYUgeLwU
TNtYxn9LUUWxAfmSxIN0r78YqMs/+tDGJFkMX9/xTwASULdIo3vnC3AbEqMWySyc
NoTsBfLhm9BEmOexOVyF6w66sMe3dR7D0u1y/Tx3XenBAJGV+W5JVKZwMgXBZxb7
8IiMSujHgLYgbNb04iwftUDjvong2Bmuoxs82scuKA8T/3oVV2Fg4ETU0M/UuRmO
tN1+EhH/jEslfaS/h190CrQomPuG1n0KuJ29y66Hwlmc0J5t8L+00xIeKAnv2UF2
FYO35E1NHkZ6peHYmBTsqiSIzXJvCpzQGHuiVNV4aFHpFrFCc/EIG5O7bGv/Yi4U
Ibt94kM/mJz33b/kSHK+cEEpiqYKrMl0HsiYC0L4CqDgnWGOHWmVGn7sKDfLJy4d
lo2u83quGdKZWA+MVbk9KnK43qYQSqeQjm/iWUUj1B0ryvU28j5FWri8lAgyKa4G
2G1wnDlK4vaYzXQRhsuXFByeFybXcYaaYYDnzuSzCjA/g9Mnzsx0iDO1rZA1xYN2
i7tr850WLyY2qPEk+VuEqM7zNEWJQd94HmoHIiLldljT5rQi2gES2glIsPYdFmhf
D8xV/MIr4iqe//ddQPU3phV3TvBZi3vIIdMjH7Zoh+8FJ36pMaZE/l93VjZk35wa
w7B0J4WhO0R8ySozMK8UqDpnQkE2G7MFLSUVmHwtbiEYSet5VC7foDwQE2UazWDz
snHvhunKPrPnPmc9KTJCWmilnPeUTCln2SZ0LKPuOY8f9p+58j0fj20Q6Ly6SrLe
B+x6qPy4AQt8RsC0HNhTuLTXws7RFl0Lv74znRsj5bh1bkkhWNtAElhVPy1AtMVv
urFhFnWvdVQxsJz+XR9b/lxsbS875Gta6EGgmXGFHWjEApnXHSeOVw2yq0ybQ5Cp
bc9e/3o+tTqwlLTbxTU++ASCGrLUn6vLfjcOl94NuwcTDjGW5IrviLA4VPhK5eLH
FedGERvbksmB128LFTotW1qW++v6mhtePXOeNb4HB24HhVJZ4BFUzcg9UK6IQvBt
ibA8eYsflRL9Tkt2issXEBV3VsuhW/ARXgPNdXJZXcZC4evaKhoijxtaEG5a7L6V
jV3uDPIyrLcZGHN0XFRSGsMndaubV6ot2fjdWDWFlKDqY8bkxbfIRjwPKY9uvErC
x2k7Z94QkjB8nXxwnRq+8Js271/7dzcSlrVIUoB4QWuvt5ZtcpI+C1lKbLRyEfEF
MhPUNLPsCqA+5uCjaQW80/TKHU9byHsX4ChB14F+98vriNkZv/XztZz7BfiFQ6as
bAWrXCPwuykGFWn/ekI361CQZL7zZhp8jr2buxHD1waGsSSFDNkY19DZ3q7CdUeW
agvou7+V0BpSwX6+4jYK5hbccwfHOsqsJLRhsEysQOJM+OkT7RGvSfz8ojGtBDF0
jzN3zhnEO33OHNpFi/A1qGVtUKrMMhpXVi2NCOg55cRMXsNu5BQUM71QTeLoxt3t
5pKCvQLJ/Le/UgwT6NhdHw+j6AVpzgyx6LKogDe7ol8TPfZs5Lva9LqUcajJ38rM
Mo9tmDqBQWRCLZl9lwOMagU+T1pIfdSInFJveL/mPM9iM79WJ9AL/+FaPaBGL7v9
r9AdOyaUobNniAOAG0qXvbesqKmfvFPKmZxEqGDzgbM09YTfUvYg7b5xMg7bF+3h
97uSOF1Dedv6fZDeE5315ZVOjS7Pn8LssqKKLtuS+bSaF4GoeIzLG4cYg1X17TYI
+5+3poH8RoVIC9rahOo5Ep+c3Ebwax7NSxhvUQIyJyb8pvR+0h/8Rs1a188NxMDC
brD4QeE5jDfLFU2QbpJHDzdHz/cR2skySIK1h1kkiCBiMyM1xgYEvsTKoWB4xgYX
XE0ND3+GCwEL0a5UsS7hHp/4UbgQ7cYXptoXelBEl5G+Ninun1Qqf3zX27rc0e3G
ZosOw3CKi21QOLxKTc3XJt262UEuUbgyX7+JY38Z6ukLzFAeZqAGksbcUbcWx9hi
2fyVu/pcxtKVwgjgNOSyEPJDR+nWsUJPmYdEV7m+Z8HHY7Yxcsdffuimo5YNxYjx
LpxrCYb9gWGXvF/n3RYOTdItmjulgcqa+qjyznLAXV+XCAOY3UiEju3EtzsXSpLo
E6sFQkphDH9w3uX5fWKM+vmC0c8u/5vrkBmjZc0bj8j841n6mfTuqvc/stPIgaoB
pb45MNtR0QK8HcCeXygi9I1y0ysOzMV5yVQI49rsAQ9IIfI9Mdr3vi53pBnVXWAC
e1dBKBibiC5pQvcIuUDBQ/IbTfpLbMqQcMmwtGyyyCRAQcpZIY9IdnY3MdHlMx9S
GTSrwnhXrvPS+tk++fRf4lsSCsZFgyfL2P+7QaxGRJLk0cKndKwWQYQ5PbCoeWSM
uOfBVJ1fKKg7/3n4nqg0ddB6AEsk0coWFGn5lYFpSXfDWqXUgPiw/sOhSxqxgLyc
BDVIu6koQuxxq/zcbZrhJLH9uVx/FinGsppWhpDzvhn3SsPMKxfNelxQDkcQUdmz
biep7FhEUBWH8X60Ol+Wn++IYyG99cCR4aTC+5zcuSFop2K7NewkGQn8fuwW7FRh
Z+2sUiRcydpRFbNzuiuBiW3nKc/AlcSmOaVGyXrbxcoCDWcBl46bV46Rqvowug8A
Fgqu3lWOoVifNQ0VFUEwTf0ql+EIxcUOM4oSGEZzM81GGilv176H2xpQP+9h99Nb
QpHKCfyrRPNf5bnnCcAwLl5ZbkXY8j1r3v92BXyF83Q24JRZdq2UfzYoBal+XmGe
ZTROEEllrGsckXUYqr8lVWVHrSalrZQ1iQ887lOMHrxXDGx8yrFtU5IZTzZhAll9
ITs1PbIp55Zmw9oacAKoyTTgqbp1Ggi7xnNe9yPY98XtC7a9ECXRQkV1rbsmhUDR
In9a/uJchF2MEOf4IqtFZqJ3wW9DaIMJMY0h8ePFwM09Ya31qpstXHlnEwKtuNTD
eOdXrzXZoPH8R0v229EQpulHre17SqS78xortAC4WFVdRuj+O+TDODigPC/MU4vc
X2oWLQjnf/w14p8SyfB1BnjwlkrxMuozMzmDAhjX2TUJ8D8jpQddksPf3nN51q5r
ORWDfPpqNSKG2fmqzr7MuWuAx1fNlUhTsIwmMS2UdCZ6S5phzPbVT9hj0we5WJN2
ZEF9PD/b7VZ5fhujXUkE5LkLt16+6/BtVGLxSVNqmcWA99BJ9zvA28oqKDXVnh0c
WuVGOoqWU6Gd8BvsqUDQF5Tq4JfQYtkAOWY6/pIOH1i460cVkiz4OsDGD390dOyD
x4CsyGNEG5zMWRWxh5CbsJZnwG6/Aegp3s57kL7t/7XXffZgkF1Z+PVeKtIAqCbl
P7FcVEODiolOycYWTynUvhkuKnKc88X5WfLdMzCzhiObIep/I347Kqnl95xdh8Gk
UmFgEbKh1zUczPZqbHDdcMqi90xSebyRKhQVHIbN27Kyjc5FVpzRk6mVq5LBLNcx
tHAo8GRJf/Xaai9DayANv48pg/3glWd+uB3zUXL1uc9awrtkbHJZy6G9yoXZcy/1
sdOgOwI2XpY0+DAuLCPN/+m6PFcHir6wOJ9/301wfHIOk8Qrix7mH7OxLTh0y8cm
SmjON8+y3rzli8Kls6zWqDkbp6o10/jeqKbQ8TJ9DykkN38z5qztmELYcdjkIHZS
Lkid4+NOT2VmbnuBN+m7iX4STNVnIuxt5MWivSj31X58wd3+4nD8Ssnrt7kyRwu5
Tr5wQIQJUMIXY1IQisIj7ny0in9lt0VqGPxXUADfoBIDqF3b1E/ZS24ZWaPJqd56
t6FYjEhrb/iX7D4CrDN/TUF8zmh96QJgLRqpkdC0vr1p5E29LR6g7O/R3XGSKQah
o/S1cNWUVMG70UuA6uI6P37m5hp9VmI4STT3pWR5ohIapmyH6Lzda6W1ACr2WOmz
DHNuDCpI/a8qFSfy/5X5rIOMsToEHMPoQkN0QrwipybHKCCmZlJ5cvcbeLTTydCK
wQ+TLMjLQP9RhSaF0xrlB70aBGwvUvQarKOGpai+n4jI63Z+HD5htDTfHZHACkVs
CSw14rlKG3X6dGOFhXpmpdJsTnWCdtwTQIWTd+l27WNjD4oiz8kM5nSTsUmtEvn8
Lqj11bH1JXM2FAv7ShA7asBUC7a5UhZC0SPlf4TOG2MgXfotC2raJqBpu5G9M/L9
zdiDnzbEAm92Pz8QyTEOZKG/xYLy5wdw0MWcXTo9A8jHrlrpvMlAtrT7nKVJyqZ9
FvrTkL7ktWWavOmH3xrdpS/4TJDOW9pR/QctKeztWjYkWqaSfbBcxs6gOHgHCp1a
wDf4K8qOLupCL+GbxSO/TA1WMsRGc9DBm7ReCYi21mGcLj9v7+vp5Z9G+qF4bBIf
CqhDI1XlCycPYXBASRG04GvmMtpgQ4H+BDDEfBD4eiiWdBMeTNnCK64Odg7xQYZW
TAUq/EPk0ScilgMGAUea4qH2QAMdlUkjDU1xQIzEqeG4FPu8rgSm1DN1MIgQa8f1
BG3u5L6zOjPTnCDb4doRk9QFkZ9Or3Nq3yNDX2LDU2YVkXwyEeuSScnc63PsA+dr
0buOBiBmf63nQ1ayAH5Az2C/QUHw+undijAh8j5mLuiwXUAEJZzkE/GVBRdIGf72
h5tS9A5gtgnKyRpkZr3X3vdDMSwY5mn0bhW+I5+aUT7Hi3BURJq2Il7S1V+13RUB
KHtJhyj3t5M2dJJzYDjhe+9UK1yzsKLU0gNadSntLjY9jTjP0XvwlpU1mImkXtN1
PDAQ7PBrNN5bHIEiPijeaQVMiNZLNuVhWfeGZWyd88pD1PSOKQ5jKy1m85RRWfKW
wc0ACcXfhtqucHuG/IDXRUq6Or7j7kX7Tni7rjcedWbG/ZBk1axFsoYEmzt8UMeA
3X3yfBtommZuM6GrSUnXSEu+m0ZiVAwMpsZTmytPCcGtb/SD+m5sR8sJiWmlqzIH
oIi0LoXklVK3VkYHCpMsJbBp2KtA/z7wu239nP/YkL9F/vMvKFYMtk586mUqyyrL
BCicY2mn6ccg7Gld4Ylmhl8BoVHBQy61urbjGvofNHubtxpbPTDvldVBqP27926k
YdYGsY9zlZNxFCwwWSoZ+eCk7He6JfIc0kslK3wP1WwzWBk5Yma3FRCVednyl8Zq
YdTgX8GyF4dZAcpZfsAIe2lq6CC7i8VG4T9ujAvRYGAhPEFevw+0O1xbD6SgR0PT
ZmfaNeE6WLjV84z3StLbXFFWpXnjk54PDO5MsXRsbWoi8MjmxJQA72032u+mxhVA
oJaEF6J6ll0SEk5PdciV82l0k35SUQzdPDm019MGVtVsqzqiJXehoN2QlzShUKtU
otl/DHGqdB16HsRflROWQlMASyP9oVX3XTs3p+ZE69gXp8Q1lhJQScDmIEx4Asj2
XyxatB+AKOnvy0GS47TzwhuErRDxGrdQ2sazyQZ5txtbN37aOgDQThpxnmfX3CMH
y2sur3AEkdnBvCMaR9QPixXA0Aa+WxyJFcmltFsyCokF9VzOAuFHXH7WTH38Y9FZ
fdzCxh/TcUGuOvtH/LDrwDOywjVoki0U9d5keUMUdYeSnueARswtqbL0gtvyGrzg
OVn32pv01OzuwuEVSNZ3XXYpMRaQW4BURQyI+thZa8MZBEqypFaWEyoLvLjv7RVa
M9XAJBtMXsMW7+ySrlQ00zYTQwkb1ZLQ2zSo4CKjWAbe5vvzULqkaXO+Qto0BHmV
5Dxb/G4QUVyVHMpVnwENBGT8ZRM6Z9wBVZwD0A7IA+8TEgRbCFBvFSPeh8BiWcsc
Rxz3koK5aAwnegybun3noKAB5A+O9OAAyQZ3hv2e1OMNFNQ5wpHNo3MfvmoGPjB8
z8Hyu5cEY+fp1vIef2Qk6kgMEJWi2Odum8KOrtEwyn3bmydz8fpKkUsDgSoODD2f
b7i2G5tqGyIaZIDL9X2JawyyODry/faWDENC+IlwNsiM5iNdmevkvZmxXLf14nQ0
eTUX4cFA/mJx8E+QakVZrl4HG7rrioJo2vEel3xm8zWJhPA5uIG95ZGrVfRiwQsA
Mdygxv/IUn3h07NSzsb89yuuGYVl/D2M/hIu+5BfsSb8k49nYsbo6ZoZBcf9K84O
PfNREWA9rSb16nM3poCRUyp2yQwPqRt7U1iiu4bYGgb+WSz9SeNA+PtAtUmxALjN
0kjlQnb6h/ehR+1PMc6HQyw58/I9ms9D06LaaxPO9v9MfFqmceRML2qAHnFPDFEL
JKAI7V/GaZcOOGVag7ZGgC8C9oxkCyvl3I/rFHMA6wugWAQXhL5v1Btyfq6c34pz
A6NSJ1dDd/TFLkdnB5w6j3DIGZx5/6HxEBluBST3FWGFW3fk5wJXTCwDrv3m2Ykk
Tdk78OGqNPp76qJygNLQuhHQ6bPhZxrHQAJJ3M/tl+9Ek3E3jlc81X7rrEWci8eP
IDiobQnsKA1zVpatt0r5oSeTd4V8ekMlZF6mI9NUe0o8rBUvXpUbwnvE7QvjPnOV
EMs7mLRq9GxjGiysJ1GAgZoghqJfhhRyfD4v9uSQ9SOgsUMpvgVHBWZTrkwIZTGe
vb6wJ1m1Hwabr/oby2w5P0HLuk4+5nzTB4wPnAI7got772uD0H3FRO3gP+wiQJTX
RbfAwUvebDyv/qxKLq16xmQE9hYwQ97IFq14Rx+UKu9eqNzeltbXdV2mXNk9OPmZ
ATN4gSYfHW2aDbNsOfJF05bg2sPF8yggLwiUWNGZHxyu/9QqSFH8Mx34KSPjTqkR
VgqGjhlP4shjvncDjqg3TOoEm34xQPbcVSKuYF/eR8eP6sEp8lZOh/BA3it+xrv1
t386I1OeYZrkqpcjd8y2sO4ULe/BZ9M5GJ3hPjB9H0bCrJtVyi9PYS5pMuNyvswO
uigxlDZop4ou7xpumjCNPLZ/4muAbAYZhDHFj7OUQKmGPT0USSm3thjMTrpCLfYu
sPo7WEw4D/D0MwM5vPiG00DUW45A96UZz9iCIm3itVAMDlEdu6Omk0R7nAoupw2i
PJ33D3FisGY9tMxXG6ZfPAw666Bcmmvp3KQN5heQOVJ4yJoRlYt3NoznOPmJi9Bj
A2jY3S7FQSd3NG+yxDr0hbmh9jAhNQQgouK4U8mjCINAOVSCV7gL30I8K+CO42nF
cUbcTjcIhDhWDjIMpwL9HbsXFA65Ub+Qs/IAG9E8JL2dfyAtZaLJ1G9yJvG7ahAS
hW3jA97uqs1s56dafQ+ES3bxRggJCtsj4FNb1DXVfgMW3iUIY7IzxKY+piE34i95
`protect end_protected