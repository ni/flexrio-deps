`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10368 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
LfLaKOw3utJqtz02pVdKfzJAd00IHyvKnC1DdN0hYf+I8NLfI96WrjxP9irNvTu7
jb0fMl7gbLU+Ti6QfSLnXgXRkHSn7ZZgmbDHjXSXHgs/wPPoG7tWvPoCmeVZ4t69
wpDUYLumPIRW+UizHbV4kmhVwbbOUV3XrFYNKpvJ2OVOqaxn0D7Bdkc8YQJSEhGQ
T/DAOjszHJ6bM+sgeMbaML53R/+8lX9y/anoZTX/14nl5kK6Ae/YYYsbbOT5MMbw
R7AEjzVX/MY1NcRez5IEbzDcqA4w12S4F/vyOMcvx6Mgo3pVcglyDUccQ0lYEhDW
wQGOQ9lztSNcGSRGJPSm1Np8VTogLNvHZPjBmyymI8/fHXzQdN4hpwszZCgS+uo1
oMj/JYI8dj0YUcXKW/umtNU0uDKvo57JPVdP1aG+XuWt+orl+1SpYeXWUtl3aEGN
XikC37Jn4dTv4vvuG75Fl1/tqgcLDF0O1dq3OD6F7uJsTEZfwMzQ6CzWHLQCpkBd
0nwTD/ZnZsQ4BAcKng8yiUhUUkn6AdunoMoAbTX2jEcZj+cPCz89j6Tvc1dNbBnM
dt9vYZ6xODgzdoLCpUO9yhPZNz1tMDgdS/0pVZPOiDzhShDCQ6dYF9l1BN2QEpca
AApLvHuiWqp8J+C3327HWtmd4V2c1HYxxo99R+/c7N2EEfgWnQnziL/zhFa81D9O
ZZBO6RnobSpnz4CDT+dSEmLv4KJ/mrMZGa6ocYMA+ftQp/ltHdYRreyHD099UPeD
XTBskKO7plEPCMPkMXlVOjidg3LeQWDr10sByttiXq+Py0fbQYu5u86GBLGslMzD
D8ClVRdL9wCV+zW0UoNE2LpIvzq5EykdwLS9CgKrKyTI3ZA4PlGJNG+VmWWZtPhn
BeK7baW2oGwb4NmIAH5T7kHP7dWSPGSQ1/YEOd/OP1mHWWR+FY2NIkn8NcRFur+I
PITU39he0MYtVC7a6q77k1CS3WeYmmfSXebeTIC4oKo62wfGYiyC+iSaZyB66UCl
K9mYUwlqYQrEu55Zr2ztBGJW8ceAZZGidRaOQAB4A4L25iYms8o8OMplaJTv66vV
wrTPKDWp/3Ow3J5gF+LkAetP6mNmE8Y8qtsuRpTHHTl4zjY93zlAqontmAcDoAUA
C6C9PDWmUusJVhx2L31+BD7G+5NXVf6v7JrVe78Pm1SPonIxXz07F9ipR+iv8Zwj
oiThuI0RXTelim7Y4b93bkxC0QF7Iam3n850WOaY9eJuULGS6dWn8R3zU4WYoJJc
tOlOzOUEfnCTy9y199MfZHB3C/H3yAv38VPtUVYStw3E+zxZDMoKjXCy61PLWMi0
cPwfxVqp6OfUKO77N4WE4XhukNE2YjSZJCBaB9mwRaTBBXrPBAorU9+VcuSjUYIG
aPI+u//wdEbE621qnVT7E5so9TH24zmVdcJMn4gUDNBNJ0ptbGPYxbL1J1if1Mnf
o/POFCOsBbinAvDmnpO7pmsk7W7ytnx7ArCh6bAhnu2jbKazQqvGo8fs6gYAFxAf
oa4hfgYyyp5Ga32TbUKBc9mAWVrTdz2rAr/gN8NUtlF8yaUorAYO6roF7d11ofSQ
n4uBvgsH2ULZ1G4wzBCq9AQj9BD9kaYv0/MAZG2IXUeePAEvDJJFh2dOSkIxTWhB
sohQuIitz2NZ0G4HnZEZH2snxLuwNyOntjO6KzTbMUk0dH6A0kExYSDEcyPn4Vgn
CMDqb76663ewkgVVzZxIAXpXLheauYCyxLp/HgheB4LvyqtAsDTb7RQIQ67p4HOz
tkJqQhVgS4//2s7mI1oPsDM4oYqEdXPS5AdzDAawJ7/R7fCF0Pohreue9St2u/dR
UnflGWDfeoZ9RR7MnqUOpmvtmeEEdzSnLg1928y43aFmLdl4P7yL5A/ghdXe+F6/
jJ43bz6q9AWznWv5xr+YjFd1IRJ04N6Yc2X6ZQKk+0FdLjxaV0KPUHY1HEJltEjv
U5ATkcTu7QPzwuZJpCC+JMZvli3eMI+1E/0zHw6D0nX+raLHrUJDG0TEsMoucVg6
git+Nrsvoia7cp76/wDlnZRVYCAydBtgp/YM1Z0tZtalzTVhdkSk7AwTO1oPK/nh
SFbPFjiJjUJANHMQWrFo4w44HGcRppjS3pIwHyzsMP7gxMm9v4jokNR1pLFqS74V
711iz3i00445GXiE4ADvjj7Pq8xFnBE4vmO1LH6Tp5gVDxaELNgGGQw4z80JeTTY
uGFgqd9zqFJ9O+u9sQL4xjEtstW7wgyEvFccjgDjzioVDLgGZP3WIfaWGLgauCLl
3I4MyPVynBEWrINCxcojDncDotJy+gtQtPCNofBQdPyRLEehNhuQuPElH578tDc7
RHgi1eIE9/Dv9fZh5UHQGIFfWXznyiyh2PwTqDwwGRqIWCPmkGAZPBNQJpmR534Z
Uyk0AlocGO9CfDwky90wr/oejAf/vYbFhpdaMQfWwT3QNhndopGZDVdkspSdkFuQ
ApuXItYULd4HLaKSEPZo0u2zHaLqSfuIosTBPhyMn/0nygQpfeDauzzi7V2mvKCm
qdv9oyo3AP4DhuTGM5H3W8LB15gK3XFnhhaYb369l/dyeLpIP9jjzUl0HquW8NMv
Bsji1UkL2umeQ7vM7WkWSkfvHXKizxHHsU1Stz4xG/tX7Pqm/Y88UCWq6atNscnO
FOXGKLXmWB+7zv9Qjii6zvOxVf7UUxeUyy0HvYz7T133rslK8Ko104F1hfeuuQML
gy+Ax+1761FaOo2iodLbbg108OSAo+Df18V0H5mky5slM9EA/PU6FGjwpzIQXhmu
DXZVfq03V7kPImIfBskWPZ2Em46fvdZc0cZkQCRL39MbBJAtaUqdIaLg/PhKCS5j
t2XPeexF+TJpx5bBYDhxc8RWVf1HjDx8H4VXV77PjPg5K56PYlVmWQmjlLW/wmzs
hgG5Xah6/FtwuyBm0r5T2/Q6uS+QIZn1sdJJZk4MgY44cnLHnN5ljavsYRGJEEQU
Usg0DE/zw9EK7ztM9iwdxPP9zO45aVOBVZT8ENkEyY53uCyk+Ntwt3kUFWC8Mk+Z
lKGIpgLgEUpqlzlkp4p/qP+XheBAAKfu/5abegHyglay08Ld6If3Eb9gETII+f++
+YhMxYDr/t4moCsTXMzOM10rEya5nomh6CPkXJwvsA8iEcpmmCCPfGwXUySM8xsB
6kos5nh+XZRFlTvU812vdUhbfLJY1WVaCa2Ebtq2kFQBqqrbFWGmmhIzgDSKk6d7
FlN2QzzeU6Sd4n06zWZs4qquQbBRF67ABeo72DycPd1+fEwuwE4EUywbOT6bRXtw
vv+9LQV+OrDHStnMuawd2lsaRXK0gBeIqIOQiJs+8GvzC5rBM57QE5GdFHmSUY6q
eXhjNmZwtenWBWqTVQcNSSm7O/b/smGdTTHWwBxjNRjkMm9C0om1wM+41GkUhZRJ
bVmRSmOgvdZT8Jug7PJhh6EZ9TmL5IAtScrHZNy06HzxPMiRpYaXEKfMB8uV0hZ1
iivZooFDxFPqhI4IpaIRPGOo/f54szYwLhUJ8jBTiAfx1kscLJnxth6+obEtdw6w
O6x/j1yYbqh39dbLTu1T7/sjVHVRqMpDgmcZ6U2aaEzxH60D8DsODn1jNL6fMOe+
ogj6tvBnGFdM+jwIbUUmR2ICLJmI/gEonzuTQzdW4mpjGbJ6lHajYsiO4H/kV7B9
/E/HngUwkSbMnZi5Hde/vqWrkN71QT3NjQDy1wzZWRnw0V6/L+7Mm//+e/Yqpyfs
swphQ4y4tQt8zkz3Oe1dJe7jVrFeu0/9D+aOME7+RujdunDu858ja4nugf/dhbxG
ThFySgDMYXnwy+Olu3qzLj9txT1ueY9/pTGIwiVDt8vIOyiPrAU7Cg7wrU10hms3
+hPH6ifL8Gx7Gh+mt1wtS51iwCpGfjba2rOi8bEtJbwoSa44wWNlJ6yDl+AXhm1U
3d/8iJavHJfKVVZ7zYymkeYO9heubNkFUDovg0V611s9svFVNNitNTILL+qaSq7c
2hbZyznMZBlwk8s2yUb6fYy4ZRPAxiAwcRCw3wg9ZGHSg83d45ytdhmsHJoW88/6
eKHt1GyXp7XuNE9vyNkjgJv7+Wx+u2zoEzWPpd8dFrwcQRqUw0as3RccGwmytUAE
bfaFLBWOa5z+zmdHVZlaebA1Jv0GveBjZ/LAvTUPNuEm8HOknnzt9aLxQI6c3GSb
Uq+hdsNc3K5+XUXvYLNS9fDyd6al6vEmpFQ33413Xf+2BvYUOG0rHGwp9g4XBk1B
nsITi4xMbS7gifnE0n/iAIqydd/9UZwJCB7Yj+8w7XflKcye5cSvVy6Agc6JCrFo
ihp8n4Vk0wVwBMs1gz08b89+REEAc5DPUMj1mfghZVoyV6ROXvabToLmUpOWJzEQ
uTrVvKPT+Fas34FDfCsKHlhuHJq3RLHh3995EREbDPziqeG0aQ1haa3F4hlEXtFU
/IOuXH7HY+E0eujiQXiXPO5VQvbvPHIr+J7Zu4PgDxMLcXDBCPgHN/k69f0ZRLXX
2mA7elxTEJXVMA/HSjsXnhHLwXip8ygEKYkqJLpYyMydpnihDz1W0SoaTfytappF
uOu0wwT0no+1Cn4yj6PYePTRJCWpYgF7WvW/2qPR3VXpsfaYgUEfQgc4qL0JETgc
oTv1ivqLt/CouiCmiC5bK3FMy/qIF49jzm6zK/A45CVIj5wHsAx3i/WFr+9//Ifd
sBEgGpfR2yp+rO/oeKDZgAmzWW9XQuBP/3eLj+JLggtZP5ePVC0Hanlxr9E8JssL
gaIeoVitROxFXzHbeBiztWkS7aoYi4kpUGS1d9+lOkwQ1Yg/ota2ujvgXKVb8UO8
ymufUwSrwcAqjkPnWz9Z9owtqS8p58W2D9jxGiMGOV92s5m/trtixVegJrZTtaEU
8ql//6poCTlwnMzsJPoCRMBNSVdAM3rpuDuWfhVoADtv3faY9bnzBdpjrbskyyQ4
QAbJ98UiVgzsQeKmGX5d0elyolBUh1XXr19bT9KOoB117gIhPX2JcY/Is6h0Cf31
R4fuwaQjdrqOKksEV/nfmlA+thc6lPcCU75g3Jzwp7LzbQ7D7LSgxsfF9XbL3a9m
rdBByQRZoluluYo6LeNDVNkpyjEwk3oBiZVOBj4Moccsy2n4h2RNuVfz/Qymwbxf
ZxsSA/B1LaflWKGORP3V/ZTnpoz6qKq+fh/aw1H+6zVwQL8WJeCIezbu8iIygYj5
Vh+RvxoEsKjSxinQIn8MKf4Bwljho8U6kyxlfIxh9LfHATNH6ConpgSVpP0lVpnL
ToZcJqoKAODNMjgPxTD0Z9IYTz44IAyq96m0fz5PVnqk/hu32qE/2QiO+XEXeBnd
IqA8FyxWN0dVsVu9JT/VjvYb1zJJsDjNZCQ8+rulv8nh4/rPLXay3JIBTOHJ0xRp
9i53W7kquHprupPH0QIBbwAP1YbNqLzxTIri27vUK+sgkE0U7CYPAJo9P22uycZ8
FvAfTKZsg+23siPD2DpB7YErylSYJaThvBWDK731SJLW2J5j2MiyeLHHVAfpvAn2
4TxC74yFZnPumf2C7qUuU549j/f0DyvEYt9yspyezMBpW6aIhskSDmEKif57mWaf
t5m+KzUJ4thzN5hBoQ4PWYSxkp5ePFTeyZhuN3pzU5sOJiT3qSeblh0s8zKOxRWk
EjCcHabPOcGeG/34jCmo6HWjM1uReed4kldpWiwUyiCy2+EihnBIVY9gb8VCeYpE
a/Sl7TUqJHELQAEQiWHrWNZn25/wPzi1b6d/LxNljls8D4eVfViU7H6k63VdI7EC
4WZ4pvuNARrYPd/8b8wUdED+65/k4HnvNjKJHl2GVXCWxgSFv9mYeMeDeaVOXZHI
p/l+sSnberwgxNY7P7vB694zrZ9MjQEutbfYpu18BeyDYpRjMO+LiaMFdkJUbax9
RQmguuUpArVa9A02TJX60tabc6fUvfodNhJmq2u+w+L1eT3OK4sRlwBJmPykdsEg
O8HwzGzNXWpXFj9yE+s9M6Fr6PlRmyvcqIA5jmUdH+ZqS4A8qbDUDqJ3y/ZQlH24
E/+QNtCLzjImUIE5WoiLsrm1L/4sA+cpMop9INjAfPWJBCo2TH7WBmzJg5w604jo
jkXFpVa35xRqX5JS3MlM8wriUxESMFtvWvh5k6pKGQe3ThXYG7NdGZrgOJ42Q/12
S5/C1NSogrqEBAFODjrMXma001kkDgeU+CX3GL33sUtelns/JEPeuiDQTNrVICNM
6WLKh8qmz7k/0dsuLOSdyF7xPWU3avyOmVw6ub289DJYqudIJY+XB1v3CrWBQJ1i
wnB1YKkK94/jyyiNfm2PduU6kDWpKyFrwbJFR2962P4iQcrvaLjT+4EnnxsrFaSk
SSzvREWvD/7xXHdqFZ5Cr4vK2oUdDNn4w1yIgjxdnbRpIkT+t5Nwdn4bhSRXblW6
+1u/oNsuPoT3dr4R1+ery/o5qZzhGDdeHHbWSHldRoT0wPxrPvqoC6e1WTYNsCXV
ukkGKtUwOa4JPt7ibYXQ9SMz8xzrRjDbDjWa7GORetXR+lhf8Jj8HTfu6QCt/8Og
2XoxVTcidzmBNE8Bh4oQ1mq6hMs4H0seu6wnh6Mq0SakKCWMRVq68ghBvdGpwUVG
HpZCI0b3bab5bvLrRPOK8ORza47kcITiP06b8lfyFCkjHijg8HtrymhrYE0hrwTD
l/A+e5cCY26xNnvvLvCFX6V6rpP/4hOD+7VuT0mSjttqh+3g/33t+eV9/SuXjT0L
rZfKX0BT0YzEcn1Ulqzp+8o7196cYf9SjIg0brag2PrBC5Bp844AYg6nlRZYr6q9
0QtCMNS0YyOXy6+jyAKL3LWf7avZiCaPFyxi3K22T7Bq/0wkDaF4XVE+rdn7nzfY
MkeblV/iuqvh0WZfAy79zLf+KQeZ1IuHV1h8ITXXLW4iAD3zAYXNLvg6k0K+ZXGE
hPqpKCL2tV+2hloiyKIP6DDXPy7dcHh2aBAr2RG3WqVBo8DkNXHSQ53owKx1LMTe
c59rEQJTJTHdB6FLNWEFUb/2kanWa9l9KIWWPzOBgaWW74n93v914brmUap8t5zw
RUpUDh5SLMx/b3a/wVArkF+LVjHAjZnjpeq4FPam5EYCb0c2CtQKoDSkpmvVw640
XRKjiZXbxAzFGUskHthBtHA9CzcAm5gUPb0MY9Vr51ZJXnT6qNoR3ZYH2cfJMOQT
9rp36GO1hCj0mqKIYRRvEll7Z0Y5ykkA7KTSB96Z04ZvbAiF/21SNquV9tYNETI7
u7nuXNov4cWn0YpsTulmzk8ZcORqd6VQf8Mp/0AeAVcm+rxLY390PoLpS+cqCahP
xEZ7ZfrIBtOx6hkfeSLb77Oahml88eU+mp0d13LSBtHElwthhU5+BlUY5/2XefA0
AjrB54IKRjmYE+dPqIRGb4OrqZKUFPAde2SdR6j1dyMGQ7uY6o++HfXJFVdzkgqL
QOFgg1JCeaeZh8y8U0xIx6e6baHAXuyIHER6nyeOuKZDNLEYu9mTQ8LnG1UIoOji
BVUMy8siAV1odqlXidTUgvHJC38Q1XHepvAvOWXMxQhLcQL+V9J7c3qNyC80ASkC
LD+9A7lwEboftFr/SsLyBRkGvm1OhcmSUfh5nWK6MKB/hWN+eewXFQLKWJUbsnCm
a6+ms95HogEHZ0ufIuzoNVWZG0Ahw3wKye8tkse6UxM2+26Iy0K730J2CgB58MNV
3pW+3WBR7zfl4qMhGjdz1RyVQdo4CJHDHutcndT7lSyM71oecPftwpfuU+S1tdYV
uOhc3CWGCw4YNlo5EUxS/V4hQKoASIT8u+FTGxqoOcSGKel/QqQbrLtzcKknK5aG
8mpKKT2n9oysD5omVg5n/9S1mj9gmdv548kI4E5GvkS0BJqzoqC6NCQaux8AHxjW
gLo0LC9pM/3WGioblN2Em2off/qMehauBWCotJ/mYFSY6z8LJMLz4r7YAPNcJ5NI
339+/2y0ZMMB33qnMz7jYEZgKFs+HdWwtiUR3/QdJDfW9IIh6JY/D5+Oe9P89dq2
hTYKEUOfGG+/0pWfzOQZBg7GQ0YFnpYCB5kET4K/jaGUprDOlPi3q0LViRKNlIsI
86EM0kkJWED3HGHL7xSq/KytBFgkD+gH+otwWM9EN+dU1MnQifEJELHW9HyBC5Pn
LSS29xWWA/XE8EEYuusRdNuhbH5kbP5fK1iztuG+eUpmcZSrNBQXb4n214yeb38a
7UNyELRzH0NU25J16BZP0fEigTmvfJxa2Ql7k6tGY0ifopfWXIdMArXBqjNjdsp7
yqYgptrZWqhosEmE7cvaxeB30o+x9Ozu1yC6QDv5lG2mzIoBmsNbtUPFJ3Ct2Dyt
bcADbs6py9IDx6Z7UjLKVaEDRuLbqNW9kCdAyAYJcLHTqyA224i6Rhnz/tVbFwSQ
0Lf5SECA0jFiLfRfx4KusiZEhoWWPj0Nht0uLoVEwDGKqsaxtxN8/Vlkn/De75Tr
rWahiCUUvabSt+DlPsR3rgReFKdDKt5K+fZCTeLB+w/jH1ddyvlM4eOqAOMAIpVX
C2SyT170KLQ4KDNsLihvOEv4Xf44qib0ztLos3tkbkPp86ntju+Xchg56S/mGKzN
nUZZKA8VI+1ZcqGlwyCxeQGdspgYIoCDxhQxjeiHxhwejQheHCJw5J3BMlVvihKU
d6yCgLF/7heRIN3vRAaTd/7RD/7enCT4EXl8GUvZnpHAxNhjOktV9dOUuxfhwQQd
q3jIk+Nc5mHUq1708wLxLyam266S9iO6c5KvzjhsYNOjPMlTFzqn/8+I5omjhjyW
EQr+/oRdknIEh6Ua0hdd9NOnEs4XkHsxB40PocBKHZO8HrgfXCCFnQMUIi2AP0b6
f96FwVzbeWy5oqy8wKAvBKTGOD+iHNCLPylqXbehHYPTpSEuQ9KytDLyFGijUhuG
+QDVcdjNrdiliSgTizXY+mq9ytaGW65bX+RzQlkRRA3nDd6Id2Xn5lHchwm25426
B98EC8+kzZNW76o2uISfxBeyQ1m4BnqQg31zqMdhZMkEqFmqFLtJhQUCdSFD+sHq
ubQzsGwRV5XGqZZBJQzxmjrescN9ihgiukAYXUiMRUm7UnhqoCGZpXImQmac5HUx
Hb6YUlOQJkwoJ1kB72/qDTazYQKFESSNqa4UlEQnEc5rU8Pa+paj2L3F+SZMF5/8
uubyRxI+tcFhdvsU9EiEyHVrBg53aUry7aKW1fTElaspN/Ux8u538VuwxdYibEjL
dElDv26nvuWbagrmOWrB4cgjoc2zWicR5YIVk5s4xe8Og/Nx+hPvDL2XRz0bLsuJ
YXr9PxDSX7ARdTMPKPTdzJpbs3LoYU6YmcUW1RH/ac4WKRMdNOn9g8ULTze6JgPS
WMP/BKt0PwByjjd9J+SbrevU+KQzRN0pyBU41PDv8WVGxdTK6xd42tzPQI/DDhGA
n2hp0OeXwB0a/xq1YxotUritoIsb7doNQ0LsZZckVnkw9KVYb/2TlERfq11Cu5+P
d0w1v/D6jtF+Afr+ClNY7MOH2yGd4JWL3MrRajVjIs3XqfdCPNgKrn9FCw9ZLrUH
mU0XIdbpCA27TzONQniR0z3m1g4sY8GjlPqrF5/5+NymC60wX3DGpuxpDVtSQHf8
YMlOvn9wkn6yoXgcE6Vn68c0ht9dPY4/crZKxvAnJq/2V1Ea3gH9GL/vMGZ8iWQ7
zuY5eJ18xP40kgtSJqx+KP1xVf+cgR10lkTi9b5SUCLxAeaK8Fhl6iiXT+RarAiH
7bHo05pkHh+QjdFJRCutO2NOz7MSXNzcALRIpw2EYtWeugclBoHbUXc5k9oYDIRd
zIhMUDUjGDsfnKxNoUmPebk1YjXyyP7i/aOVKw8MxQoO/0KauN0HCpAgfkXfi7A2
i03porn9X54X1AzjeLEMdQMiM55c9S1VofBPvoh7x7R55/2p1756uUUTALq42i6W
pAjgwZk3yNA76oI3yxv0Hh9aQp+4PjB51rGR/S3xFO+QaRiHJ9hqpE6ADFBHvUfm
d49+0U+X6rXeK486WpIsYKFp26y3HDzzDcrVulBOtZaG0JM9PIcMIqPBA4yMnsuY
HR//EwRlrzZu6J9IPf4WHb2izqJe2CfC/esg1sH6PYcCa/ZQnTwpNMvQpLLIZPoZ
O+e+u9Ye5gLrOtsbci14bey9G64Dscyo/EAr2EbkZXt/HHqqGEsPevSD5LCBbbcQ
JgEAUuBp0pEvo9BFu5BO/S8CGrNGldi6KTFh/Kr+KnV63Vi8J2tdPn3YkbnnbmuQ
8LaHT1mdRijJNArJDcVohRLVTP5BTfxxtz9Wb0m5E78uPMRsLw9EFvDVCN0tdqCu
D7xzCl8pFNhWotC8i3T5wNM6YabA24FzdDcJ4bTAwbv+zExUipWQvKQeV21gz4EF
xj8aGXaQrhvuXSgZ0gMXwW8VuQM7+MVS89GQQg28Re2Xnmh1CRapoJPxLlduXezK
ScKTyE2AZjWDAd0HLQo1WW7TvKSU19a9BO1P30lIE2fOF8pUhTadnVTNi/7BXQmc
q+mvRLbd5SKhJWpGYqGwOl4awkIVCj8QyCCjBHIVAHQf7jE0pthuLVtRcRCn5Tcw
/Jjc1WFrCX6oRcZ9qGUsxC48qPotfo88zrCgv9jIUsyMUe+ggr7Yy53iJoOHMyjF
D7/O0KRjIURAozeWHP5sRRLj2M3MR+VcP3ZW+Uxhzq4VR3AslEk0ylN1+27uWY3r
w9YANaFXqIWV0yr1LVkU1KbbM76z3H+S6iNbUj/Wy71gOvs20811meFN/+2SwjF+
4B3oMGdiC/PDmzLGV47JoRuBdIohCVMCsdtcoZ4xmahxwm6vbhFChBOfrr6SrP2j
cEZJ1dGc3PkpjyPXECGmEcg6LTqkL696vdtb7+6fQq0ar40v6l8QC2lm2LuSnj5p
L3tXAXIPfGdf5dVFhSQPX1N0pUYrp+b7G/GOCpaIIzVlhKD82X8nEF8hW6TGGJZU
6Pb1cAUQxzz7mvmQzTu8FTNg8JrlwZUuztv7PG1EQCKOKXgxevJMuSlaY5DTC/LE
//l12RE4WIek5gJpw/V1Z9MRw0aL+G1kf98sRuqUgAX14S228imljWOB5KqE0byM
JZZy1XBBXuFc5n5Pi6mNrhxU1b+z7KNR/Il8xfuFMCOhFOs2plfseAXg3xOAho54
fU9Zneswl1UGdCl7tvPuPwh8udtrFtHBGaUp/3UxvUNVJ/l5u5mex5Za2u+W/u0J
ncsOKgdDfXY8NlTVkCkwps/rjymIVD5qA5nx268Frge9eWd7w2XsNVAKBarxQ4yR
xA8M07DNlrGgvb+WTql4Cq1q3E2sN9qXdwDvsiV+47bidvtGqqrDXC9n7Qfcok52
p7Co/oC0Ib+M0W+KCF52RBh9C1eLMrbs6MiN3NTYCg9EU9vt6tDANNMMw8Yz/mE7
XVT19a5C/X3KapKt/EFVvxNr8n2Y4Dbi1y74XLeaxIWEW8I4zI3Bms+MI4dbfrcE
4mIaDBY67D4BVv7KigMhCn61kxPTJWWokX1Bu+5pgPLRPWGEa7oN5t0rSWOL84k7
PHGVLOOd66eEAJvnaxzpM3BYEM5NF3rKkd40loiO6+3K9twHOCczF6i4w46ktEet
Q5KP6QrQGJsAvBlgNMrF61zIpt/nINWBQ3QcH6E/KFCW+JW5Tlrs+oo5StyCDvoH
cZLemwICOX788l7G3wW9DEgd5xDKC/u8AQTfQq8PgmqlYy69FwfjdPjGHvJI82QY
blx1VflTaVx5wpPfMOK8ls2t3AxNfrzHIxUe067GLK0vMCkd5XirtHeTG1CbNk4J
zI+e/kf2mQmMkse2hZ4EsmY4qWPfb2ZHr6MhK3vPoHAFBp/fw8l4CipeJ81E5agh
Y+VpjYx+yI62WuAE0gaNGM07RlBk6skEn4CgojkSZIVJEwWDdiI/9VIWJh0hshFU
6tI+5jDfoCcKLuAq/3Q3jed0NZSpFnLdkqgceCrgVQxI441l5yZR6w4fgrNG52Cn
PpAr9s7DqKmI0fdus8xlvwAQvu963OXfGtQPw0WlPF1X/fISeaxe9gCwgL5U+R3P
HPgBR4rpfXCuJaVQvEQ3vfk2by3FkikUBq6HUKrbdLwb256HGXTOqWaluD6PdsVO
vYE2MtIO4omKfcheFS092/iBV8pbObSEXu9wGxbzcjaWI/64JsbNV7B6S5HiRsjO
MGgC5pDBsnqSii+cj/KJ/O86puR4QIzGx0DW4o1er82Y8sm6QkcWs1mT2TP+MTIg
VXD51gcxXyvEkAGR89pWab2qPKGS6ZZk1YjQ3+x7K6kX9mvvcSQejiIx//1ghHdA
gL90nwuLp7dkAZnVz8Yu+preSnYTr/jSr4VXJOcl0TmnaGQRKFk04wlmlzP7YWpY
hjeuK7RikPTfnu/MwGul/71Jxmbo0X2FqZDBROa57OsYLj/pK2fDhz39RTgOaVMC
YG88Cr/qtMbGZP8Vm7wwLtCYrhbkRti8khj3bZ/9jqo/o/Hy/Z35O28JJii/wkxa
vzMjFuIoEY7Whper/JNpuBndjLF2YuAFzsMQkpl3MW2UZ1ULrAJKWe05bZm/wkKa
sa4wUi/0zeDwedSQRJV9emfgUUmiXGQc6Lueox0TFK3SkU3Fljljs27FsOZrmx9j
FN8+Pr1iM/fU+ZjSPkS/OcoR56tmtCljmP7PfErPdrzNA0pPVJj4SIIBg3Vsihlj
3F27u6XAgKiYfjG3ICMu9bYa5Bfjfg9EU/Si3vdgo0jAtE/KGViKDvXy3DCouwNN
ly8utxBafcTY3KFHnqsamuBVor8RRP1I1oagVSvhx3VqLlSu+q48kX2sQoUUgFvs
QjPKTyQSfr9K+nl30vszRugk2jQ3d8HpDNRG6D6ChWryTQ3JqFZi80UolwZWciKk
oMu9Dts0xKiqqO6wRK0Bf6mQIQ+/ZLKtmNutyE7tCI543HR7QYl1mJptyoCBg4Yp
64rWVXwFcgwKc5ieyxloaKm/r279omeyWvJZjbMlhgCzJxYB9b0A7cNDtCmfTXgR
ZxRX9Wzio8nzvQ1WR0bRleOjrHC/Nj+jc7JGuux3JM9OwzmvsFq8RFy/qH4RFtol
7SDyvQKb1y09gJTdZ3hq7TuWF27na56s/8ECxSCewkZ/mmG7W7ccNqGKjCvxBIiM
kZxGclmyR4ZnVVIKI0C4aTbyx8uz2R+ndmnV2nSPc3y7KwRoj2pERG+4je9FQOSb
eUY6xjzkmrTk68OKjqWdGamu60XFPM1T5NSiU4pglRJ8md4ogjcvCgpoDv90HlSf
AYBwoRWXZ8RK7tgVlEZ+0g4b1DRvyRiF9DgIIYgTTbi9v4VB0bJRHKQdeToO76PS
aL+cIquYEcclMa0ki5heqY2UnIqIVNZWf2gZnUy/SDwvbeHlw8BRpot5lfqzeq/W
zPYAmAzkFqESOwrOULIFuEakE6FwPD2bL/MKP05sQiua62+52NZ6w1QoD2oUBvmc
FBxqa6xAsfHjvRml5f6B/zJbsRnx6NQxQy7Ds3M0eeGu2I6+MNjjCq4OCElciSEG
R4uIgwmWAan0uftsc8DVMRe1l54g+9Mdee6sq/PsVOmLTo2IjNq10zoF/oyFlz3E
SOh/eRQwK0FZyxdgOvB1fS/Q1LSzAq0gI4/3wPPT8x9pj3VZM/hW75gSiIQO0J+o
`protect end_protected