`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 55056 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aVlarhe+WUv8WRJlOJJnkAG53ou2yrz0BcDB15W/Sj+q
0SA+EygBYZmRAeXS5ded3MNiPSvSdZW9ELoDC8vWMWb0yKCQx8x/gXiWu9XhWO8b
VXQz3mfh2UblQjz6JpUa9I4efgvRQKrLVORhbi6rd+qoJ29gNdI+fEyUToRet18y
ouPHi+bAzQ6axjf9KyceSwhmNtb3z3DQaBu5QTQJd9QL9gUpbfH1Nq9hQgWGYcDj
WRCPLWs9itMPjc4iVumq9VMllP76HcNU8nB0qnYsowBx3ajWvT5awgUYbByH//h9
vnxqdfQ7JVv/tuF4MVi5+Ki80WaSIpg8akb5mNNPCYJx4XoHJXpLS5kWRRM+scsO
tPk2eEYhrsfMllyhRpA93xsOWdTkLhIDNr0Gl+K1hCLW+oDm5BeEFenk5nfcPnVQ
L4d24LGuekIWcdEZ48jT7EaLfPLDCsqSxzDHzuABOjrMSGi92DnA+Ridso8Xo7pw
0luvuvvG8gDYoCpeYSfcy0eucolSF82Y+Kk0pNrb5XV4Rs6LQ7IWTGasct07fej4
kZnw+IUwWp/HOT8uQro4mdoAYWWnCodBoTTA3dG6Gn/9/PyMH2sxiQ9B6izrqih5
DkzI8c3HNuYbaPMxjpRcLhFagfEt9lwnXoOwv/1tSbjHt1QdcCexxlEAWoqOWoVk
WSer1/7v6vQ8uiP4e+rFg4r3z2AfPdFk/pLMrAqQ8xvKoXzljiI4/PTOxpTKNCSF
0FC1ZCsy4Ww8XT0tn1QlDdkHW2YEmDgMna7htfWFyqHyRQt+WrF9/7TKxkgcfDNd
gdUFjztdbPMbPAQoA7EVhqpNT/dMMKy5RINQjTNO3iXORwL8hVsXk7CUpAZ+KJTQ
6iLNvdXfBdla6VF2jh/Q3lCHPWyX1+cTbbnswRrkw2pBnIJGtAZzNFFYcWN0ZLzF
ORuKFgFPOnwQRc67xTnSlSlAFNDGRIir08p2stCjLH7OYchlWblqe3laVm7cx18E
oURVWJM5H2Yjtz3v9NFQdQeDSaVyVfI1RdXcotd4jLyHqcT0HCe1EXDzSLPVs0L1
WN2bGk6cK5AhXeMNG01kxplCv2zpmJ9Tkl0y0DPrBIy03t1gbPszBA9q8fcrpZM5
tO8c8LEhilYGTuBXNmrtLkbFoNdB8tibVU7BUeMhMFapcp/YzyoYZpQjkQchSaxu
eZrqmBRGXcfrVyBcvm84+0hTQCCAbTcaCApHn/5Gj31DeGyVoSNeNjsUqHIwVfNS
I9x0Ean5RmzdHPTNo8uJ/SEPztL1a51udtRuBUGJhac4plaQ4PTNOob8sM+6haOY
1hsHHjMsWutJysBZ9dAUjDn2gNT6EGKwNSIwe43gZPkSMcl2yd730GH2ZIwkLLOs
nqAAhU4aJZQIu4VSuklzz+RYfOO0yLGolNihoxEsKyyrY+wiTxu9C19Ngb5bOTF3
RYBSKVprRZvJYX3iobbx4mfj/PFMSzgR0ryMnTDz2LYosYD3YMdRoUnIgncZ9e3e
LajArF3CJftRPxzgLfcaAAV5P3InhBBoHGuu8vV1binKLObUJJR2ulqWS5g4BmKH
aq6fAK3B69DcRdcjiPcm11GI5QMRTYobK6s+tKXA2f0WW2HsaRfkUCkPY96+7sd4
jMP7QQN+Wl1IUFxXKd5ll6VxgmFFCMD4h8RDRCI3/qoCBKgR1e6hg2r3S4aN7omD
kpSpahouvtVJIwA2toltpxr0EP/I7Rypklx3MAuv1rGCfQCIz7AogASUFeLodsz8
YzvMxvvc5IzynzencrlJgCAK8MHLHgrxy3iyE4hWjSsO9r4rKtQhb/Dz9GNQe1nz
XAVAuS6ND1wWcmU7TiNnvjusIExH6Cu29URjullROPUDSVgqV+hc+sOZag4eJa7Y
Z8csccLwJSre/M/FXnv+cJ1y6p1LDask+yewfTM61hzq1o8Bhv53JhZclPgXalQz
1fuXzTwQbC+6HkmnyLIlcxwcFkehjbPI/jeBSFQnxet+4S2R5T133HLLquRjJ8GP
B5dmUSmU5JmDtLXJFBBFCnOuqMPk0T5/QR6vCRtbAPTnDE8RR+JPV9JV1mFgIeoH
ZFR3h0eLbvQx04WarSAoP5OohFj/LWufOJLFTQxLG//tgvqXZ+ivsnM7TQKlBy0I
EutCnA4++XNAhGIild6aX5ksy+MrG/9hKDJlA9YKpVd/Od/7/Uj6rdfDcgwZ1k6K
gQRcCaBr1RLSCQ0EnzCEyfG1SkdSj4vkh+vsk09fLyKqCM9fYFJ0sUVY4Uo94w0s
KV2eOuLCPL+MBuYznL8xEQ51ai6+U/T87G1/8d25J756gTXSYsE+1YxFFsBDBTZQ
+k5BqP92oqaKiZo8YIw/7lkY5LWTU8HakwNWESoCzrsRqb3Ltf+bH6RZrhGBG0T9
728VpacY45aC5TwnJ4fFsR0ivfA6hUYAgy4LZAxUegMhYJyHp8oYr/mrRiKUzI00
FafM7UiZdBp7KvPaKz6kECs9RvoO0ojLDSrxM+F6gH/c1TtK3NB0tQoKhYCpBYM8
3Upwr94NsM8MYEmk3n/FaXtVQzqJlFebCxGfRvol82TyTDdjk011udBI3jT5LQak
UhhoVyDbNrp4FSsPZpQWqiEidUbwhk9ZwlAOL16HL6YX3deceIFbo5p2P1rDug1m
JHZe4KJ1xA1MKUd9Dj/+99HD66O/1cCqP6cBr/xeVh7dPRMX/9kE+izXWJGcMRfA
unTYta67f/0qEDGWw8xZZyL42HLvUmXV7WlILj4ys/PicBqnR4xVgShSD/Bwnnvq
0TF/tEYmc2QAf2U+cA5yD6BWKjUHc8NpSii0Cw+lmk+K7TqmRmx4JkeK7C/V0ify
Dh27VDbQ8hZ0qpUNHBpDpBZr7IRzqagvBLhHqVphS0FV9h3ucTbHE0nNEVZwKYNG
wXrtIq7P2beLdD7aqP1ESssgLjKlzaDVnE1wwyoEuvEXk5KHFQ4SF63R1D6dm3yU
NIy9alpAYmDgY+mwJECIs66ti0SfHTV4w2Tjb1GMVRsQbZliRQcPpyvrNCSyTsPE
xEIEyGFY2Z6HQahLrtCVZO4tGIs3W6ZjNc/SY8oPKRgAXZ/vk29lzJTC1ihOh9zu
CE3RmWBeZDiwjq3diyzgu8AGXyfyPWPJUs/l+3NI7l1nYgHk5bTde8Xe/bYQbBIT
YfCbHILmw6b83E/rESqk9KVTzTXTPrcRpitJWgXtXA9Lq3BExGXjxoTrXQv50ApZ
zuHjVG+uiQZG9XDzTC5TcAxQeYuDGsvLtKzEe44uPAr3+RVjvoDhD5iVqDzw5VDA
Spa8z+cLn+S/TISAHEvGfdKAPckYkI9otGt2LZCJ7JUlZnVlAVog314rb2BxgMxz
MljOFX8PwBxgEXu79HJbqjUYQkagZME56gknPNjljto3ZmVGq1x/Nlg52O3wjzvA
RTjlZK8lKF72E5ghOFcO8B7fksONoacuMmgHlWfusqCuYCA4HRiZ8Cwnalj3vjGY
8/8Vk8NbhqKg4ABW91JDdVR9LwrI2BxeL+uLUrUWTgvVUJO8VHxBX6+pVhO46Os4
hHJ7HcDDfqmPC0hlGUXjnNWFQXl9eQjUR3b8MZE6Ha1dv389nFGUXhE6xoT1Tqqi
yNCNnDs7eMUK/Dq9VgxCWfr9gTM3f+eLLJeYgXEdQTYkneD9ofTn1Q3w/92bIfD4
XrEj7d5zA2bKiDGhbpTMlmJ780NEhAFPllNsD7PjTZqQcfCZxe7rySEgM9ItemLw
ulFH70Ic/SgqirY46cKnXM6oc1DSqs4Nlj5vSjvRmyirBjrgxfL7y2BYddzJTZK7
1lhvxVXXiCHfOYK1+mZW5YkQgzAxEJvWd/SPE7V6QKQkU5hebOGbqNg8Td/XUjbs
thWDbSU0/eQ3fp0PVPluEOaiQ4BmpnTR26VpTi7Py97PNBbxE+N81viQCUlKHyl8
4quE4r+L8QlAwpRWIVlrsi21CdcZdRJ1Ti271UtDynEJPzVibwWhfFwAXw0cvqo8
o/nMYmVQeAuTs8n+mYmpFYTIChFLTlbZ8eTWqF99tLZuEubnqZlEdlXto/jnOE6j
BlAFJ1ldSpBed20cWxPungKgWb1kDX8IxcTLUVQBBvm+YYBjkPLSbBGwB6rhUaA5
yPbXSFVIPlHwMTApxORs9X6Bw/M2xAPnZm40c4P7qDSiozpzplYCqFOkxdQkjcCw
cPmAVPNewuONgxa7HXVKzcZelJ9BjnjIfkENmmcRoxuTDK/+HOZintpES4eF94ce
q6Qd4GSC8ptxR4/WxtBAZeAdUzUtgUARSl2wSjggqnfZFLjYnqyzuqLgnapV3yEV
sVDOctLxpTRFJ4SifNYaUMzFDoRy7ySHLBPXDaXcH7oWB9TDjFT8mJ4S80CORa36
IWYXx4Q0d9xH31EDYPHRNIszjffmX2r5CrCAaU0Qnr5V2awHyfF6NAcXlmabQqmD
ElIabvezOJ3Ver1xEkT+8mgHL1VSDjmS8S7XUmlCZ1ZRyFxQHx7c4SvFq3n6ek+l
RP4rk5UlmfIKC3XqSclq/LrPleSV2TWdkx7pT6aAJcZK6g5vCQMphnuoCcNFh6cR
227YQMMMZmRncz8Qq62JviHFR6iUoQq/RwPqH10zboApNbLPweugDmGbGY3MVw0C
bEckdp/Hn4HlUpWQ84vfMmAuI+JFP14Pu87yTkypABWWWd+5kirNFgkDS6z/LsjY
VSFQ4v/hqOxCQUhIl3AIHR1XjOqpdl5HtckMZMOt9OooMILDhQ9SqGcVPFcWDyb1
xTwu62zNmDlrUWlDZ5oQm1xUZ7t4sePXyC2voao0cDj72FGK9goQAxNZ45Z0VG3h
EThDtd1zsmbWzW9H6eROtsN6v7kH3Ql7432BxNiZR/OUv2A6tRyxOjyZJUHr1A48
f8PS9i5tk2XwhAhTDEZcew+o0mQu2gd279UDFNmjU8gi70vJ21Liz8J6g536P6e0
w/4SlpBJmS+nHWEDAXzVkQ0JKpCKNp6zsxbhe+xvzqMWbJejIhQa3alkUTEP/REA
SNPyV8JhddnFpzfBjU/IDt7iFIHQOfaiWAiyBJz+gOlvZWWlMEJLlCXVPBvuEj6g
LVntf1MO1uiiyxSHF6+iZ84OSCfWp6HPLp6vlCyn5zOFA8DIYXf9P+6TMOIya9jN
zCTtIYJwBnWeWJeDqV3KYz6+8oVNRH6YiXa1av7pYT7zkIchcmkNBUu/ny9GzLmV
1uEshgTauwemjctaEJ6uHdu30SbKJLOEm7b/pFjNDvNiwVag7ogRI29nn5nYYW72
uRqsdWvB2as5gZWCHHHIZEUagKZkhnzP3jSh8DAVsJgyMLhG+gy72IKQq/MTysMM
oDOZVKRVLWLdbq957dKxAnxgfLO4Up9HW+dEE2bNnX0zOllx+ixmvTBuUCYHdTHh
+V0rm5VNpc7mb6cSIfOlEnPNKEkNOhC0sfcC4Hb2SgO4ujTfLfX+qOZsNMhN+QQd
ioLcn/KKSPIvxrxZ48b7PXEuBtJDLDA/bsrIw4CnsQB8Ct+x2FN9PO94nm8P9ecT
dWgLtiJAUlM6eHT1uKHfQSGXysrozPM7sGseCtcfelBSEcJQTbi5DnkLX0TSQ+Us
y6mdDMmY63J+FdKRkYUkyCuxk2doBXQHAD+qpQeh2IEr5DSh8PDAHoc3O8Tg6mWI
YaQFEuUMCaTrc9JQBkAwcVOR0GJe5y0VspX4QgIOlTLcHeZjLhJGFLClAMk8+4vR
07DWhK3psLCaWDNw7BW7q7tCUBd5RsXsRp1PfJOuhYrdsOPVJqPBqiFryEqE0kNu
f24/0xeM7LtziZe6Zdj/L2Oohx3G3KoWgr2N3RYys/UAuR8ca8JeJBgaWTfyx6Dy
2/I0ZwywPtEjVtowH4aADpcQ64A9E6BxOTFMChbXfjfoQhqjXasnzv+akWXuk0/c
HjCZqVdZLEPB/oBCVSSkN5VpECb54ji4RHC/DSTXHzIS3AZxjxMHcujwi3jWFoIo
OjkgSMxijLkaAlBNfNWCmsyZUYIhT3/xP4Gzkv0vpjuk+maAbLzFvoQ1jwPtg9FH
f+YjnfDWO/JjugDZtQamGUs/SKvNYDrw9Ja8LuELZhYVotWrD1GHmkIDmR59+7X8
wuWt0rX5WZ98ERHJzGmznvPHtgFaSGt8QWMceRV5V07CfrZwXa21jXAH6WoED8WA
DWldebwB/H3skxS5vPJSe8D6pspla9J71p+qaOOhNFa569ANO/GK9ztFjk5Vphai
gVqifKmsQHSxVlcoO1CZpSd/0TwEJmaPenSAgIFeXS/bs+v1e0NFHi0C8gttUj8L
gAicYC+CYZdPGARyf0uiHUEOA8NDOfYn6AvaD2JDrnjHCgn/RSjJXdzuTukcid8R
n3HJgebhM92IJeuG1+q5qaMTo/jxNYSt9dCLxdX1z5Y44vtUsyoPpbQY/heTnR22
1VaUTmm0jQrf/qNT77IN4pCdwCgzee1Gb+2dhqPQC66JdueX/H0g9yAjOMn2JBit
/BXoCJgM7U+I2SoSIEjlVfm3AKVbkYv7n3Kl6Ctc5QL5AMCGqpfVvLamhk/UGBZF
RFrKs/H+FYOBQwNCyQQI0UutwC0YBxWFP0Voe/AhBYorvuPzryKZUYNsHPLHU7Bn
QSH569FmtgIKwB1eqBnRiKKiSboqkcG+rQ7D/t1agGRnDWc68K203B4RVej0nht+
cMvefe4yez46X6sEcH8bU/UGpYt8OubVGqnYY3NFQgDQd6ZJqPvx/eOsMjkVkr56
hoZsZLUcyW+TmHYFRtXrSgDRFUeckK3f4wNeHK+/J/+sq8fS7LcszKGveFvxXwXp
bPEembmg0/JjAfGfcA2jusJeT/Ps1Mu4C0oTysrCoVzAz50ECoCki2O2yX8hGExc
CXzKJqGusGWcAav+/luVeEXLeiQt1q1XR6Fja1kR0FOqvfimDMmellSYtFeGp2Eb
Zfo85MxuD6ipMwyUyzy7LZLsZnpiTDj7KHgR54l9XfUj4IpoplbfoIFmjbHoS11C
Kh8nZRyz3vipGR4kMWpB97u6XyYFtPK3ozxZxKq6leuV5zTE9DCPB6vV1vThWkp2
CWzG3lNEFZxO+rs3nx+SqHCbOgrb+YGfoTOOpECVDmYODZA29lMYfD+/ZdapPVI3
YpfwVUJUYywB0rdM0MHfiCb3NN5JmlGskHO9bGO3TOwfAG8JpRYjbzfMvTSNIzGU
hln2z53PcsZTbuyQu5LMoXbu8qDt1I3jZ53m2k/+pnS/IRYVBnzWgAEPg8i6Bskv
CJ0ZiaA202yKMj3fl/8RYYcW0FIhZ0vi3VGrq1Ml941MS02IcQ0h5YKayDtWaptC
upiaa8wydDic9r0E1CcawVEieRPSNDwMfw2GwKZFi/BIpyzeZzAXrHt4fcrnhiWF
4VH4XgxtOYnRS3gV6pRt01L9AFl233Tibm+WTzHf6G3N6CrXqKXQUBUgmdb404x3
P2N6nULKFgH8x+zvUnPjs6BADo0YbtiPNfNsMmC36zFEqiNM2K5rI3Te9TBD5Wxz
ogOPkmymDyjxIBxIckAoWpHElLRlkbVCj96HBWLSXmuoXomETfwLfjgV2JK0sgGz
5qVACrKoptxfu/c4N0mH7yCTZ7mloJrMUFI+9V3QKImmf/GlmSOAIXW9K9gueupW
x7DGNOGGxYD/c0bHtNrfShnQYJIYJ+AGMlbuJiTMMAVtc0mvi8BBXR9N6PbUE/G+
9YcnNhPm1Wamlc8eoMN1AOaIGsAEidTiYEY34M2Z3FSEhevFDYegCvvwLa5Nfncz
aN3hg3MOFYRk8ElD/m/ahkRmP8za65cd+XfDvQ9nI6RQQiZe7V/c1F5llH6meyZy
Jbc1vqGLBIXpt0HICCRRhShLWaYZqaQ+OR4ZVR1Kx0sAGP2FUCkHTR2HQ2IUF+QP
SRNBTZtGDW5tXWntwNAWf4miVhHg1wWMWD0Wv0VS3MsBC/eWydobCcAKoqt6b6sh
YlTngNLlf/ifUtaw04/j7/VMuD0jx3ieVlHm1l+O4cjPNmxehfSst8+h/qLly4W1
oI258cliidywlWj73yBDQt1EYU3kSUSStGiDE02AwJY3KORWRFMYFxNlMOTDD41e
+m0lVOe20KenSOuag/6IuEuOfnrXvfgtH7JsPyNKPlSkqiE5B3S2vAMuW8+GHKgS
vey7vT7ZwTAyKaP/k9kMfTRog/zPqAEqys7jw+Dx5yBgWYyRstStmtsVitVxRF7g
DIeN30GEVFQqmqkQI/PyBVZR6iqZ2BF/SZOWOs2nyMeve8+tFiPgqNBcvl7Tm8qh
aoEWSvOvP40hjCibphtB0+Ln5YkVTxIbXwXescaVp1iOiV9Xwxra2MOgLwvDdyPV
+C9m1FJKny++VnPPk2Bl+Q1PBZba2dKdbeCbGi9xO1H5Ucw8OKMedH0HVEB7/lJl
ehqZ6vvVIx4Dm8sZfGXD8xq/GHYlNLBYBOQiDb24v/1waQVncveF+qDMAOZl/yIM
nouljXs9d71nOB49M9jPlDjZ263LrwFhaKb8/00qewXzNRtzHt5g4ZkFCzHmCgBN
v0MUqhbmkXNOq4Ebw+ooYdrGvyO2AZsTJ+rlGQGcE25aIcR+TcaxbTmKvzNEJvhJ
A7grGBk7Bb0waLRFDesNJ3yjk1Rr0ZM0s956682WGMZSqlZFOKtoRiOw8YaeZsqZ
2ak3uZ0xz1k3VNB76rtuOrHO4+VGVt3/erMy08H9jJe52N9TErkyP1mukefOdm2v
WisR3CeRl7iLN7wbuNKHIf/Zq8HTOWIpBSgDQp75r0/jMf9HawmL+obfpq64tJT7
3LKCWCldIldEVQYMQXiqzfhe0SR65UDr0+dcm/GybZBxkJeKkHc4yexmaUUFBHJJ
h0KYrsG8iah4ANrEDCGnY4cQcuGCXuUcJzpv7UXW/pU4ZnVvVgVocTeFXmQSq6cU
YrjODT+KrSeRs5cbsd7JOzVGEp2ki7i3U2a5iWFD2U775WfVSlKp12yBENhoGvxa
yMWqSHjil1QEl5CA9z9AwFX23xdaL9qeTi2xxWbFcjrqZa0js63wS3wHbQtnPcqu
ZUpAFwg3CtnX3x33LneIF5YYrwTpTgoilNAxWfCVtSKYBiS7bAguWZPH9t8N+tW2
bn5Y+LbcXPA1ALX+vrQ5OX0VAJWSIjdiswMIvcCaBNzFnwWjKF4lK3vfl2nSzqmY
ebQr1cnhQzIJqc//2mexQ8qYacRoKsHaPpQiZuhI3su+ql2rk9paYjEzimZWvp6G
WFetvNNlt1yXCYRWzuc9nHSlibjR9M9Va3+p+waauU9EcuFmU19Ww5R1ssiOMYSI
Q819m9txUDjWI+S3cy2b2HQt2nEJ6UALesb5U0SYF2VXJqVu6QPNA9X2sGFrzUP4
gxTahoWoV4sds+IG7jAD1G0G2GPKsY7hDcLVpoXP5vNxJa1Vlbl4HpPbablKgNIz
Z4yoDhnYNg2ltTV+nwXhRjT6xJIENf7vrkubZ0Zob9JCc/h1cedpzxjkui5WoU8u
HiFv2a39hjpcHurgd+eXWe7+xVRe74onLaH/kv8ZBFCjPCME0zKeOIWvTksYXFLn
vjl3QupUg/BNHxalfQ0tv5A4l4nq1BHpTFvyvr2UHeiLWkbgk6uZF44E+PFChY7R
15HXB8aBHQJwxmEvGgwCPUODMLd9Gic/O0bp2irkV8fl5l0/ykuFzopCCw62SDS8
fCKgikSOp3yD96JuqCfDfPaFYI28NPFhvsoet55JXyFKoN0vtxuLCpsaklYd0CdL
FkqWmZpEq37HxOXtPQPh3iaBSPQ+VR/eFsFddVxdTdh++uUb3iCAooewGbx4OoYL
ftIxlgkmNmav8BMyqMumDDPZRNYZq9z+Kj+WIMZVHgUfbz4jrpmREqlWrQjDsoei
ZBjwCneMONb0bCwVgr01gOPzl7QcpUrAIy22dG4DFY8MiBkCP6YKYuekrZzcgDaO
utUtdyeZm7ZogrofL15F39hKdSqGAlCR6xk35Xy6mcfP/N9heU3/p8OTH+VOxOp0
ys3sOYw/SLqLjIsZF2e+HUiRCNGERIXK9cLhusLIh3E6mu+7QxtPBeHhpQln56u+
cFpx87nDk8TvbR0BuR2TG7CFAV1GYfrHslNHMmJs0crFVo+jLRqbsSJROTXDARop
0uv9qiZYSfWP4OiQEOTg7RBR/cS2Kvaxb/+22iUZEQRjc7cwjUcKX0jCw7Ck6wRx
DJxZWulXV14KkYoNNJUYZHDVvEFw+by2/dxfkoFrXEdw5X0EowpDvwz76pALEh9v
Fn2JH7AB54AUXo9vOquEVOkTAp8FEZGAE3N7PjSIXl9cMu9gPCjvHjhPOdvEeF4c
MngpdCjhhkTCxdebl2/1to0ukALYm4/SA9rHA6AZ/vATJp92uhWpDqoJD1AFFtIe
Vnftst58Xk3Br/V8ozzYSg6nCSXg0/D97DAAzn/FD4bD2QPe4OWss+2cMlM2oCut
5TP1wWaL3aXID/MAhecSLBxxaYEdktLu3mJ+PQ4vyHwBbo4OW/W/npg9ZFKyRhre
AKd/idYKlx12EZK4Bk3jqXMJfOEz5yZ2G66CffONV4yaNUukyzHcwwImtPGKVQCh
BSZZPZRdZFKzg10UlZealXDvKPLUSBfvealrS3OLYe4GI47nRjhzaMFL6p911rMj
YZnpei7x8nT4QJZRs+MFSyPLbBZEWe8zpqSDIyAmFNh2abPJTEru6GOPRSXtC/ZR
5cDOfmhFuavGklXJiJzWQKY7hliRVoL0GN00NI21fMOLOoA9L8ZbfYjmNXQqRA2M
t3GZ7xobCqXPMxi8oHE2RnbgmIbLYrw2cdHXouw0SW/CnPAtAb54hI8g310+rK4L
waIoTocujB78d1PPiJDwWXrJm61mzPRLP5pf5i9WpjblwFkU+CUxR+jI6BsLAr0X
jGhb50lWaSNxnFnUBlwILH7bGBC8h/XkFwkExr+HH9sSBOoFfgmVAfG9v+9IYMFx
06EZ5dfknVprbAbqrlLDTo+601XxKzS+uIv+9MRXlJ7ry3mlVMegcVGO82b/dyXZ
2s0Qd98PnEpJrcTsVJOtIAzqPEFw7m0zDT3L0Rqk9obK5ez0Pv/XhzAr4bwyI0UZ
oSrO0VkyheQ82J3IMSQL5HsKWWBWF7vkDJI1bIVBXNrwAdiVXAGTrFrIeQCqwbUF
NaCOvmi7gglh/Pw18jjouF5HvnQD9psNXOUOWTX1CCZnqqZeB4ofDMQ3jRR2zw+B
Cs7qv/GeZJwErfyboxdLRoWSsIZKL4HoypGrK897NR854aasD3jGfArzYHPZVX+S
z/e+qlpTPEmeBFdBKyZalkEGH+Rqg+4MqUIedaNONvnkbUGXIQNvhJNdd48vnner
zqUeGJeIE9GZXGUgPhI/zPhv0dJgKi3kh/WZgwRQ617zkfgtmrCB5xmhu5x/KQdq
UPkpWO3QcEiT0sRJc09AgdTxMmx4+jvUZglB5RfRjhIX5ZJxQxbL+BrZbeZhLQod
DqWevK+4ZHoqmT/fmIQ+QdH3KwhmB/OghPeDgLq5aHKS3M1UX3xNbja7UbGyI12O
ptuFzWBYsi5TrC7S0a1jDU2I//wStok3UoT/3TVV2bkvBh1qMvzuJ65DXm2M5OzH
pc3s9yIAbSzC4BfUbR/7wYrhvmkCZ94m0fUp8oBrePsF8aly/EBqaUoaP+u8829Y
V5j0gXNfxd20Kln8LyY29Gk7TeeYVErIIxCZiiATnHEjPLsLeXyCNrSZPrbfjJAE
M2bNdlzRUpW5AOZAu2/zfRFrMLDI4CHVLVeeqYLDM7zYBxEACMgjSFaaNGQVnG07
pBWsCfp1wqgFbXi6hoA4q89gg4rUTErTGTwvYqOqOUU0u7moYE4o8itqKl09Xk6t
Sw+vscnssun1YQVzIMjTY6av4H5FVtKdphKcj/LVa9s+48cKMNZ8xhi844SVaXc9
cxRbHPZR9VjYz/BJYL/U9ECtk3V1TL1ino5DNsSizoBVgfz6hWnfH/zYIXFGnPjs
W7Z4vZ9LRNctbHxpn2tq+N6leuIv38GE1ApCZ6NFkaoZ44ZmzuF/ADUp8dVpRyha
SsSSBpGveHl71RkF2Y+HqZw1IGfmhbRI8jtSBb6nCXOWsyxJsOQxsCBmt5wQGVEx
RsrHL5OE2qM1VOIBXArU/u0JDFGn/jqiejmZzkR58brEQ2bBagSqc7S0xY/meJoY
AUTKZGjgbvi4qZWON+P47nPNHnV6xCAPl/6NapbxET/n7ws8LrRhbOXiuOdu8ru5
XEez+rYZeavU86AMjGYnd3a44Z5miPoXJuM75gGINF7e3MtxJ3Rcc9hLrBVXS4rw
k11dASWTPcTO4ylQlA6805oUgEe097bOqIQGBmtb6xJzCEX5+WiERNlY5JDQ6kZ8
c4gLTjy6b6j6nQKsFEOYxN+m1NbxadKOQf5h+3B0m8WtBuGgQEjpK5UVlIQi/f68
StOKIa6WMlFWAW7Ma4U+Dpp7/ncYEdZ2GpizRdpvm+n8vdOsHEUevzulB0Fh2dUn
phk6N/NdnxnLIoLqgnDnGxPov1XWBHwXkR9C6Fr+6T92n9hwJJhdvEYXtaj+Id6Z
SIUjpcS8jnb/mLWYhsTkkITWWdyAYn7CQV7oGY5CTtblymIlugyGZnWzYe13AcHa
JAoSb+zy7zG/zfbpev60PtvtcCz8CnzCUhsPK8uq4mOS+5hwWYeCWqhPYYcUga/a
nEIsDeA/GJeBkPltHhGmLsjH/Xn121Ryoh4uxg2jbSJO3+XdC70/lrs2R8CjHwLn
S1KMRRUokqiGVz8b6M9cCX1NHxlUpLrU8bCqH+zxA744fG93SpPdQWUtvgDW1ZXB
dWeXpAEJ7x2p5mQEyRY6pj6oM9/Np3IkkcMzQBtTzGs+78MqGFJNlAfKrOXhyqWC
bwaenxgsIu4LRT9PVpeQ9A3H5psnM40Y8tWJLbnfDGczsVYFGrp3kS8K1dlFx6Ev
U5h3RtaccUtu21JahU8cU/Ad6Rs3MmFUUV1ZVdBVg+ZPup8NF5L7a6azxezRKACU
AJZD56TH75l1EatNnJUF9Fj9PLhLxjrGvv6Ypa9IvqV06XuUkPpkcD2xV3EMKjI2
9okmm4Z98NYJpbPnvyIDjTkQt5vOanEK5KdkPSlts5bXbM3YyRhm8BhDjr35tyQt
HnmaMJA1RLFUgUyH6JMfi84HFuh9QMOoCayWEhFjyGFBRKXdN8brjzC2Cl0wHJws
BAXmKAIRCSCHpClT9G+AJXAL8cj2TOo/cjYa8gizHOXFF2SedkQOd1bh3H7Lj35w
WQuCWW+7V1U0/nWKlhKpuKrYZeD7LM7uzeYfEJHAPMwEyTtY81wwE3e+h4QvLB0G
usHkFXojxFEwaKy0zowOLjENmyZmh/OK7NQlTrXNm2cPzbEIaP2Yu5UcFBtMXiVs
1wMu8dKrDsGsRfeTMhDwaPd9+bJBAlUM+gj979fJ5tpwxiahWCYDgW6gntyY5Gu+
bSCK8phF7MoeCFxIe4jKlJbwaScwIPk2R6B+5GC/j6hLQ/5y0SZ9/dw3wSH5N5Dq
NbFm3w3qYnWBwwU/uREl/4UrdDyNcnjclmEOyOTgmrK7S2ylCRBk7P6rMs6h8cFW
M96gQaU2+DqLtD+ScMNXBzfqZA9BgPOOqzoSV0ikQAf79W/h8yytXn+wy9nTIafs
biHpE9yeJqunAl3TGF2zi/PMdqfPcqq2oR8iZwU1G9E59j+JVSsieQiJXmLludwz
siIeAl4bfP0j0x02vNOdPoyTSIM9v3z76rrMnx0PX9TwU5WM99QFBstOMGSfTTWA
JLhDFB3qUwjwjVU8yy6KyV3oKVzCLS7BWEiLUMxJ8xLQmc+OIj46RabfffvdzySk
tEtBEmMEUYTVxkrWTufWJ1tnHlU2A67QoUY3fammWzjfuabPzVN6voggIw/qyNMq
3iGnkxpB44MFkwUt/3KEAw15cSxnA9St1Y4fs9vFaAyod34y5MfR2bmAvPD/namU
XwBEwa+xZbvewlX0qsS6DAf9Npv7VnqHIfYDmOmpY4VJLUQyJAIER5Tm5EIIj4bF
x4xUhgqSdhA9NFQL8aTuhVPCOXr8tUXtzXOHGdoRo5EkwFpEX3D18To3uS6M+eVP
/X1mpix4nQ7GvVD3+tK7nTrxdOdwtrRB5TeEQBNRVUW+AFdNJeUOLbakTCdZ1vrn
86ULM/WzcDrmXKUzxf2MWPVtwBOoOi2yCL9+WF0ADb8cEnmSQ+AceuN0vIiGhL75
zYs2ZjTCeSp66gKmqd8MrSbMi1qXUimthWBoFHsEwo6f9BAJG+Ws5su1Rxpjtpw+
3m34FQi/761ZqJlFVGPyv20cXBsDVUNyW1ABR+1GebPFvknBoHXQhn9Qbg+NdDaC
DCCYUoHZRqEuYR45rDzLOgTDZbU0RahkAMAQLnF4Z7cEIm6dSmSa/oXl53JWnXGn
0Uk50UisIZAXyKgutqJ4fvh0jAV9Wz6o6VUqPU3LAb9q7UBhU88egxc36XquSnUY
kRNaOKUNDxc9lVtX6hfLvbbLJbi3mTBRxp2tYuPDZV37G2ibXOHXeagJuvgeZMzK
4/b/n6xW7XhxiPGnUwGERXuCMFb+BE/wo8XOCwZ1+9CsBs/d/4MIFyNygZM/s8Rp
uakHXp5ho95qj1FshJKuYsJ0XtPkO8P1eIZeIerHzrk68NzyNzxEj/nW4QkvevRx
bQqWzMEPnE6UA4rWzGXkuhynT5afj9kn4EVTmnoEpabTDKEtpBwdjMaHMlk8RHlw
UOxZsPFYQ5jcL2Ou7/L+GyBvJPU9aw99pD/gNJXN/cLqST6gfXEQ91hNguZ/ustz
e9UWIUNG3YBPr+Z4YFgwyl9ijclSslZCKKYpYJtAMMeMYNvMwUr/eQwlzCd1F7uV
UuWQ7xuIxv4+x9W7xD4jy70HdhVwVS5PFunhHsBYbqmdLBPtwVrNwPxNiCBOf92I
E5Tuz2s0GfSshIUeEztBqatRr0BoJ+vnX1L+SyEvw/PLtxRqYj3GP5xtOzsB5Lbq
E9UEjVvOdVteDTWhL5SV5EaWnn7VA70gwpKqmHDoMjYT7Acr9dYXOIZYK9KnaYt5
KxF3i7NTFYyWkxdyTTejBAPVQ6yzIUCeRwZbOxptvjoS7D4UyBEmUh8QVpRq08Sj
Goe7RS8TZXCoC3nPBIEx1Z97JQFMK6TXNYmZmyZym1+Iq/hlRbuq0VrEtEFqbJik
TYb6y4aeW8lW6aR9yq5hBEeytd+hZENweeA6xOt2b8ENRA1Cg+o5R0gXWWLY402V
NQtYD/X274jRybaipyzx3XVI+ecqXToGElZ4wj2BCTLJsmffduqBWIZzKgmKlcLz
GPl6qUorhasqMZIthmqfKHd9SNjzV0oxSfjP0p/NK9s1ifVRbIOFl11V/JccY8yL
yyn6bgKM40V5zj6cthjiTeDdpEBbOb2u9yDYukviPM2IEVMs0IhFFudXgM6MhuuA
IvFRfcH1M4gs1fRStNPqtD8jQtZgFlTwZF8cZfl98WAO8vJDECv+vmtlk77heFLk
AYNJTza8iLxgDyzqRlzXn/8LWstHiinTcWIneamwLblqi4StVB61AOXU92GVsBSI
clScKOVNyUYEJS0nLWbhYUhnxmaQZuw73Wn7aZ9Ttg5XaSPtB+jbhNoSO9ZJkQGF
M0VV81q/CTiNldRR7BETGRP01nCrmu1oEv/IHQzv+1ipbfe8x8AhaScW8oiHJ/mk
fh+TTdzWwz4C0wWbQxbqKi73hD05GwqfeOblteKHcsvGUJsv/uhFHmPi6MhudSHX
TY/1jxEGjsDyh5kZCQjf2n2qLkVmVvUDUO1VxU3FKfrcK/vI7uLZ7kz20WDpJVnM
6UYv1dOBZS5xTUL5zmL1QlNYWU2rPXP7wxuG2gGE6z9wYGinK1v4wedRwU8EjKb3
cP9mWUH0tcYB7KeQUnOajGGOvAasy9ryhwINWjHSEWthLCn1J5rdWH4zd2F6Agh4
3crk9Br8LaTmOJPMXd28AVhSYEW7XXJFpHXF0bDVvacvgssUvH682rDiknI2ege3
suSM1NPoiK3AjTgIkPVXuWWbNLmzHhJOsm543UWN+iMFf4u+GcuPthl6n6V51WeQ
aDHXiO8vSek5Yg0WEeycl2HWLkpeuRd+jo0G4TEsGWPfrNOcPR24ULmCLk+ncicR
+io7wuQ9f4fP6pbsPGZAbwGFo+bTaX1R4L18fiGUXGPJuEYgKxuO73hnbELNFEWe
9JKcx++Fbi+S/abS10p7YARRZECjz2oOPZm+ln80BZPP145o8gSKcNDN4bqpwmYH
7t+Fvr66H/oqSbmEDKKzPlFQ/yM+v5/FsvPSbkvwKyEgir1EbhHRkvgG1J9ymWkb
Vkp9YXIuChVjm9A74KrivV5cmhW50qb8czoR6CsvYQz0GxQNYhT2bCR3t4qiXilL
7IozG2Svt67T+Mp361llYSULkqe8ElXHgQI+Gt5cqL4kga0uE/HJW+qYo9KcI4Sf
5RYO905NbioQQfy5hp1t6vcvWVc076wBM/THNfejee5d2TB+AMtgxd+qq77k6vjs
r7Slt/7sISz1p8fbqQkZpPPEN7p03loHe7ygSIIzqsbwlJvmlsjMq/rtpvfo54U6
rD95d4+6HpGK09MY7ZGpHNxL1TMzkovTaK65uzJWmzCglQMgj0bQPJYqE+300aoI
hXepQJz5MApLt5PUGyeLYqJ/Bs9b6Y6Xrcftk+XBwroN47dEstCXr5Cn3RU9XgRY
Yei/dUz5M6biHsAhs3ygIuUGlHFI2UJvxWPM5P4a1ZICBbaR/CdLeMC+FrAW8CN7
wQ/XYMX8Sobwx04RzJPh4SfTk2BSDe7yK/TTOkAlYbhVI+kNKxMxp29+kicWXpNP
8NyKLrvBubGutuFV633NaTVmh2tlYL4+f/QA41ZGSNlAz0l+eLE0aEKWbJOW9zwT
72rOfz/nEqxIMAp7vgkUZQ226X7oGvcwu3IKHBbTqPW0vW+b1eYBFfTyBbOdomTD
1i7DyjDNNBtCWSQdyZuoVyu1+1UahX08Sm9fB90zlEe8OhdTBE1jOaRpGHiGhK4J
jbmix4iXS3frGTMEUy2pHg0X3MrtSD9OB77rGh6Mp1ODtFrNcJjq3Rm/E6WMK8zK
ntxYSSSc2NXddyO2DuusssqBO97UrL+fN3WXLVK5+bu1ZCwoNaWhWZBqPqnQcJ4d
IQDVAkV0iubXw4tmEDEFVAav6jHt7CumYJnKoLLeUC9vVSUAvZ1DHRaEaxltoF7u
Abvo8Df8DIJ0OLldiFriyiSzEoiZCs60l2iugmdKMoAMvrU8bMTLXAXRDLm6ICSG
KfdBMdXDbe8g3li2vp2sksoeYQ82BXNDAOI+BgAQbXu2CbT7/PSgnPJDD6eV8wPL
oESuShOAbXrqT7O8D9niASG5DDXtF6igzeoz+klFcC53lqSspyiC8jqxeLH05+oq
2HLkWwm3GBW4IXOr9YkYXfyqVPqFGWBmH/sUjxn/WHVf4P89dU7eYXl1zmQ3XA0o
rXFhxHMBMtXKFQN8gtqTBH7r0cbfAQzchaznzEeoQ4ETdY6koaICmgGioBI7fWCs
12U7r7d0TCTGg9gT0beidmkAJP6qSut9PyJZVhgHMj+RzHajyH6kQJefbLDyWRt+
zE/ntBpSyBTITuE0O5YpgTKOtSRVUva8HOlgRsrhJkIPWmjEh2i9dZ9wcS1HGB41
wYYreEqLJ3EpStRKo7hniJMLH1G99lYaTGkiQhZhJsufojbS/IijoNVb98WjAQMs
KDqLPae9kD+m8L+55m2ZotJzMu46625nVRw8xaFHBSAP6HviyyerAhEWAU6xyxbc
mHGXXUcF6eh7ahXU+73sW2OR9HoC/FYNvbq6OD5fB5MiH2kEDV1YcHVJ4YB/nmCz
5LA98HN6GTx8vwDS/SjB2JYsSfiCq6Ts5OpTDAbOnAmRJiSabvEmithY4dAi3JPT
cnHyoxWEaJlQEo+IEh9Ry1MRLUL+hpoaJaSDuixYxefIBn+v2ozatVoTjlKgmIvF
45+uwrH7R/fD+hl6N3CucWX3wLZAx7VnsOIV/3pS/eihgfwvjAcZszVibdDd40Kv
Oxl9DO3HVPCIZm5mI2uY6kLWxqpmqWJAk7e+mtB9gc/VznoXYebdL1po8gCrFZnd
+90BSErfKJcOA/zHxMpoa4wIZvxEiWOqh5DLQ654Kh8OtODOlYAWDuKP3WPkzGxr
ShONXy63HvgxtocKRI1tWqSJmS/Miu/vD6isHoQtN7lsn+jyyldshtCWGBY0dwxM
dtrA9KmHQYwbe54LvvXosFnHJDqlCKOFF5ldyAohmU3th6Ixex17ay8LUwtdCGSE
cBMJIrPNE6BXfh2cjmhwhz9rGtnmbQsZwLp1yQDR85/z7C25CG3idtBg6lkQx26C
IdYHQzMqzQ1ULch5VyHQAd3vfH8kgiaznQelWap9D6yFdwDHe5OHfEQq+mZNZwZS
pe12E5ExPSAl7zjfVLbK9/JK06vltyIQmaL+kUDqaE8v2tt7AeA9URmlFBlM3ZjU
Tki/+u235c/aiGUCNEujrhUw9ky+86NN9XmaTUr8VXiT500z8FBrkq9YJ3K6Et+R
fB910P1G3Ck85mF+Rcc/LeDLHasS84uTjNdUr6TAxDtRu1tK0DyHQuFzGKP26lbk
235rTiPlpFDp+/qQCAS/oqexv4rWsO04TFEMSlvysAblCxUQBDxhI++wthk6h+du
revHuO1f4C2wfjT2SFsHagTprJmQESCYTxJYHlcFZETdCzH+cPOQvEftrULLNYnc
UuZvndlD8BFPKcCoZvEHWDlReIYeBKLPrYVZVHQcDVpv8GJi8pgtFdr6MjGyg0V/
nIrZMUhiSG65Qe3rytL56xstZfhQnCJPqzj+0KWxdhN7TyTGoo4SC2UeiHcu9z64
M95PAAHixQCq6b8lxWeUUgvhHkm/tBqusRBONSp7slZlmsUC8wnxfKeIDPNee8O/
xlGHnba/t9OdrC9tjukYh5D4vV50bQIFqN8SDa4oHlU8E6iXkJiaPlHCqvQVDMTV
R4FajG5XufUK+FLbIO0pxRlHiYnul3cM5X6PbluEr7C9PZl+0+3Oi0gOZFH7/YRE
IVdHbaHh4Tle+OmnwasPPPdh/ZuClbppMZINib3iiYaYstbBxMOOE764SCWFv4lX
QFtJIhivbjeGcf6VEZNvmuZXSTmNoWm3frfXi5nYtanSuB7AZxT8o3f3NmpwKBGP
irPyr6FfGRl6CAMuJLbYW+XYjs9E08K96nBLIr6WnaiZ4E+LpJv7zoCsuLWh8BVs
tziaiN2Zz2x2gCr53jPkGJwHRTAtNLYzMXgnCexi11JrJ0WGfY6aqLDAc6kk7OOK
H9fBn5jAfaCN/duEVCRg0hqDVA6ZSfHKiXkW+cWozeRJwRjYS7kUlbiqeqOlEf5U
CpnK1ypIbVpoyarvUihgjnaxcWKzOR+HRufMv6/FAZCF2kcGp5HBRJDAKWl4bWhn
i2E3hC3qOnWyH2CAEFIh12qMZJe4QW0ODW/Q6VA+hxklDKnCS4ySA4IS4u+NXgHx
Ti9kW4cQLn7WsphjR9tc0R2zv/ThCugAqo5+CoRIpIZU5GWhS2PrwOOgKqfZAJKG
35FCah607z8/dFyx9bT+mnqAQycbasawfDgxxeYsAE1DXf3lQ91FIr1khRfezcKP
DHjUVbmgRi+z33zJ8yBSKkWM5wXH4ONT5tNjEvonrnAAyW35kkL3n/zfFyhz4xEl
TSgdgjqB3+CyXQ1olJSy35V6cbWbYWCUCkbSt2Jsvx2aJ129J93gPBMHT5eZnLIA
3lRkhyCWBiBPRstJzueoxaxjImmDEBfbSwI17gHaYmSHKdC6ybKJyucWl5AH5/E7
EYZdZJy1fnN4eNMw75XOOUpnMVmH/k7FhrZINF5X1MeVIQpS7mXuOCJh3wmoCN9M
o2boa9tkmongSGBn+1yS2PxhzLdV/e36P8jn2Or0LSTcEmetqgeJPqfimt4FaXI2
9iqodqaiUiLg2L9ZVsu/rh6m8FZ/cba6Wfrg8TtAOxvVtHu+EKcVOKQLFum6aJMo
wJYEsE5lKJYerrtoNXnWw7pPXTPS7p/1CSUQZL18msgc7ygXDUbKyW8Sfj16AHo8
sqq9pYK5TawdibbE6HCjHdv24gx2tNUBUDBAJV+qBAyuQPenQTuYJutV3pEqiWnz
sh+7SQ6HJSMVULtdmV1a2SRc71doNEv9UBYZYRsTq0+92JaUQZXvSuzS5HvT7E9E
hIh04CcYefoezqxJVMcyyiTgzODhJ1pMOPGBaEuCSY57+fSUNCsRckGzluEDJ9wc
0zCvYK0WWglYbFkMZ+K+8xSuUJosV3fC+0kUk+PZYH3qsb6OuT3l0ba4jg0nbqnx
/U1gHSuUh9vMboAHW0zGne+F5ZJTlcvMfL05AzFjk1lS9lyoJ94fEEtn5IIyH/zU
213RWJ7zckoZTpOh1y/2Mh7RatJLuZcRr8nXjRbfWv4QqcGjAdZkP2MNkBljV/ec
Pf9ifaWfu7WPXlatT0WiSUdor33C2bdeqH5sTWP1QdrwgMu8BF8iK88BpB6zo66h
ggotiJQL6iwoYzUDGyz/XaCeqyX0pjpv3OSELTgEd5N4Cab/AWzXQ8FGBFRLXeam
uONOCew5t/FN4n4kEWtJm9D90wI48ap/RRqVb1b1/MdjVEhzH8VrYCYv/UI74Igu
Btf72XpnFXwqWWvkSEJXP9Jwo7rvgx3Ycu47/uOwqNhPeylj34NgL9EbdfJuQ0Lu
TvJ4cWxHQT/vaRbqU5HdJ6eniJAQg4kzHKOcTAEGaUiirtiZwq/w2q5z+NczDPx/
vrJ48L8FrifVo/tlNW4eaDDX3HWvjnifabxEY03pTyTBrvzRSrMCaGBYDIhaEb/2
RbzhJ3Mu1H7DJFIjCsouf9AlNFtE1TGyxh245cVV4cmMTOMMGuOPQUNbp3g3ttDh
qMF0kUJGYWg3Il2vdhQcfQUbZ8NLAlPXA3rcwZcurIT/HWD+Xe11sxhp7Opm4STX
Yji3ei5jqygnhNvZz0gpzgl8IIY5BtV9zJnADxvuuf/ZUba1LW0R18tg8g2Bl9re
zOjpISfLyJJMFl9lTnroYpx25mVEv4nEpLBe5xs7HHnr8wfNdnSoSDgSYv70Yf23
NRTkSxolV0eHGk1WhY6m1CcFaXWYu95jAdXQeFS2b0bGbm1W3umUaywl0cljdcGY
/mqqC1aL0psw9e+N10COh+VQzbaQ6D54jeI4UafdYqayDGVzIXqSU7z9lTgNUQz0
T4fbmWEcHss4H/S9AldsVdLuL7MOTBBLonYn0e2hLKV8lawHmUU9nKfLAOIqI242
S+gxumYeXHsMjIBDMb8KBeXUx0PdIPMnvyHGQ6loVawNmxfqLiYRL8onf0ZoeECc
N6l0zLIrINTJ7sVizi19i6zQb7hA6rpyHXsD3wg6thVbyGMjeCVDrUD3CAN4dKRx
sHNja2LmwDp+Bzm+uCv/xuDEO/0EJItOQjQeCMWETHjFYm1u/sUsU0bx2BV/qsQA
Ef/LU0b4KgSITvFwuIPphuq9nAX3sZlBJeBnIFV2c6R7xNrw6LTclv0KonR8geyw
Lbyg3CzbgYa1q3Un8qAj/pPPLZUEosI/S/uwnNbTuhhbJ4xH32vgc/JINw0jnRRk
88R4iLxi6RrwY1gVqBJtMJFmtlgCAkXbXbP5CNLqrJT7tS4dVb/7uRMHvV3EG8Kh
Lf8E/RGuvMbPk0l0q/Q3yqdINJSJrlnUsPiF/nMel4TThe66CfWNsD/b0MmkLDti
tuQcAwFx/rGd2lEkDpTh0jusiPMyK/P1n65ZECe8GeYiFUHGXBK8dWx6MoskfsXg
H0gd2uCMhBFyheqDzr9IxAJ3F3+D/eqPNAOJ0ObXXodSG+SPXcJpghf/tfyYOpzI
HY8ZOcrDkhSxpVZ0Z2xZ/KMzEpRQwK/8z+uDLkAnL2htOD6CApRnfKhIJ10ti339
n4a/i9A0OwC2UiFEoaPgdYrvxbAbCN99fvIy6MthflkgNTV7c6SEOmFUgMltlzgn
5zqdgrYASCI35UKLDZ3WkDVWVfIzlOXX+kzd5vffZGq2TIDxST+3ndxoXhRnspPN
RAykxuXy2xmP9Zo//rdZcO4gTUcS0QE9no0Q+UJMq16XX5OlJ6HLnBPW+/OBB+Pu
1qRvhLXiChu/FXAUk2DJSKS6mJDMNEax3qSIim/COwMQWki8OgcFMyjkgrQ4hSf8
UupDdZ3SHjWdVzcyaqi/MWY6jFXhToDKQXA7+Ld4Q/9fLpXtmxME13QDTyrNdM9U
+gYqAcDDRC4AaBNO14J70UxSvi4dpg7b4f/5l8GM43ftzH+hrSsUK8g0qOqvf4wp
mDBwu1id/aHof5s5GhYd1b66/UAutF7fKaF4jX6lFo5MLJ37OxGWQQ6Aw4W5MZRW
XdCTmsg/7KuzQvhroMH8wGMp7zFGBfdNXNxjpGigC5Wsatt3U2S2ApuwQ/C5Dfh4
N/g8kfKEO2ZWo0ChCPDDNG38+XBhWcJ34bEVdva3FZydNz7YEB/ApyYyYJL+LnAw
zx6LWig6HntoPdrOR0lYKVaT+Sz4oKuSyZNFh1+4chl3FsSZYa8sf2K6fryL6Ukz
DR7SE6AE3OC47QxlXSVgy5Q/B1K+Yi6JfjJORxLB5LwUQSqDo2aL2YMsaspjVJgK
6a3a3DBNItSrxUUHTfIocM505Y0Zbl8FNcWj2+p1GyWnn87Uh0s5U77eUqjDXuL3
prtifgUbkGASQVB6nUlF1EeD9s3sGr7q9GGc45CcTUH2282/3EqKXTugDE1r0eQW
tmgVkL4ZYULYJslor69Wu802dsamuWRxA85J6BJxsFofQ8pKxfwOXM4o4co9O2dZ
xy6hKSaBO86lbBAdqD0z09q+SYTivy4OZ+h7rzo+AwOPX1Vcz1ZAYrr+gX1RRCZW
1b4s7o4lI7hfePEi0omx3Qdzi1JOIZoQq1vapKwxTalS/40hBuwjRuTDaddZIrzQ
DhQe8l4AfqUheTgZY5bKEyCGUB81Dq4tez7so42TTIPximS4BuAxFxAm+qNwWunr
EMMMWwl7gn1zUGLI/4tkPqtZj3a1RD2ryMQiLwGrpe3szYaYpJE9DZp3e+m6Xm9Q
Qzacw1MzAbxYL9eAtwg5wEsP6oiMEoi8+40tuh8zaTRfriIYQ+WByxhEhLtM5RiH
Vg/JqlMujYkGxzWSNF5QfuE2Rv+VDm3VrKRp1e9lpZpEDU4Uyv0kDJoHn5IYNp9d
KwmUoXtZkqgzg3ATaOvWhdPlxwH/cb04ONh7SsbKmJkL+U6xkQExDHO0wWQh27ax
1xuyT4FuEkHRUp4K8BKrdLIBNLzyZ8IqOBAdOG9lUlKgpkGP2IJbmFgOcNnHBBQb
KzRznBb/+3z++8MrLipO38NdWh1w955C84JTSLRTMs0IJXmnpEPO0pjs99gWK5Eh
1odtmY5wP57JnnJ5Cg38UI00Ud/utAPOhsejSqe5PUIGK6b9gd0YIXzKKCSf8ka4
XwtbXAPbnvAJNSd1vCHWtj+muNisT34HWc1rIU7NtjpTAzHpwAAgrK/Wkh/Mx5YZ
hFT5Gin6/LptxhZczKiCRZwWfbcyP+EpfKsT4gA6eFfwUWRNGdWFM/J/b0dKfE15
Bmd4rKIeHXUu9eiGgRYSVZoThsr/UNKMBZ64+giNXXiHDTNoazWQb1vlkKNujoMk
brepo/8+0uyH/SsWPkfKti3Av+943B5ZEng+BKSUnCfaEsCW5COyJkGoktn3QCTu
a8xkmFmIJ2yIBJX8JPqhN+KAy3icwuOOsrfP3Qzf3zwe4y3908ekYyFC32AQ0Tkd
HaFmJXjhQQ9qh5kouocyz0Vc/m4uODzmgwcDwbY8xTuJ5jRk6od2JvEBXlBfCEjR
G3IQ9AqRgqYuqTqXOTQ5iy+4ecwfVrrGm52k5cZv9fw7xoT5+2e1B3UTIfLalkUC
otWvPsxAeQJHTV7aV1WuVBM/GxjR/HUrTiqQb9cyRz0PsNla7n9e1ZcK1f9eoak0
a6CU2Av9NzW/2F89FVecgVCrgevjzyZFEbTfATJG4OB6+AW+M5RQ8/3aAgLZKk8J
Yejf8tmJycyoyRXnkR/qmz+ayJ0SnaOgh1nlXBrcvycUOlaYVGSJsGeXk+rw/wT4
VMm+TBAyeOu5UOUz4tBUMS7PRvj8gRT3C73StydewGe21jPqNsBE4A2CfZHZ8NsR
jTV2VuAtCroGBdVvJsOQ6Wu9wWzm9y82hozxIemx40UVss2dqPj3CQHhg9O2qoro
LcLzMu3+5+ZbcjZx05Y/PeqjIEKVdQbn9EeCShoRpnkUxaOxqr8TNIYD/rnGLSMV
Txbc8NqlbnWrnWEer+zoOOVU4MgaJXuG9o7ZZYcCpLrXufRR62RbpQ8x5eyjYwrA
JBpYGWKn2CLX8/aoLPfytyKwC53ehUeBEmFALSIqtemTqZnOxu/YYgLH8k7Iw0fL
Eg8KLkSHiDn+sX3az03kd5JQZo8mfiDKAzi8gn/zpbMDYRZvz7dJ3Mi1IjK67NrC
4Isrz8dwWLZS0U/ulImyhG7286Bh+PLDezSyit25YkkYk+m5lCfn2y8cu4p/rOOz
yUG7iwZ8Q8PTApTmA0NT6QFpPbOqCHSZTHFliIchWE7c/mOlXmlibTPNoh+P45L6
/k8SNOdPFuNRan8MFeABDevJHZiZhSyP3DSdQN0qKAAyBWUncc/4SWVYMZ9SYs+1
fPCXixc8IXWtOJwaJuUNMuGSOjJhtlMSo5OfpJTtNjts+xGCxQCNKSQX3GnfAjm1
9IQwHcRIxQGmBpzSyMC0Y5E4E/Bw6ryzVtux84ILR2xN9fwU8Nb9M7xeUPwsmQWJ
o+vorU8O2Ifyz2/3f67lCF3HuFm2GHbYhMgM73KGlCtZ2fgjLZ6tyzCzM0hECf1U
V/0CXzOoNfOz1K4Sxq/NdEtzN5ImMjXicHIntCd2V9SwdkySOAmLCKzCIo7lUpCc
f7IvKIUDif6F5nVT+fITAPMGgJ/wO+5kmwtq9FM8A+QPpyjhuGdfjOwpR+/t/n3L
YUCnJEgXpjFHZbwyOw20tMZETs/Vb5rgY/mwdFzoOuXy6k440K9YYDgC6aln14SG
hylilSP/Q7RKojkG40tBd8g6TLDz9bsXTS8VBdaoSrnx6b2EX/VER5uRKihi9UWL
TW0/yOeA2tY3SHg1dQMZNymwtSJJqRa8n95mwGTmt5z7jftD3+sI2kV8DvS6l7VN
DYM37dQI3toohhVxkFWYVzTuivM9jp6laoetlnkXoawg/p+BtDt4euQ+NwVObtix
oneZZhxeIjuGFiDUpmVZQDIZkhH2pBX0tCTFkY34beoWqLfC3DkFZYlkNK5Z3wLH
Iu2N4u+OoAXFbnPcNusl41Mjqzx/JOk1vOFtbO9TZ0rZXs8wZFX+3st9BLJ22aGG
kpDyGHC1hzAsxkIrgdSp+rlbvsr8NrPWAB+o6putI6hTMPrF5xS+waSqLJduvz9z
7QabfPjA0BfAsL5fIC9w3iK8SC3Qb9wyCnckV8IhArZtWofr88oa7Ox2wiJAfBGj
9nqJawrstttv3nXdZ5kmgf9MDMDSqT2MUj+CLOZ5ikvv9/25e43VyRr/GO4jjtGq
6gHPw4iizSwT+yD0vdeG1j+r0uTHXp+0m/0ubmmKDcTK6OVefWul174qZcx4IzSm
fH/obj2BU0gO76N3631+w3spDICFv10VPQJf7Q/XaFfC24q1pjQkdHqyyeQIuNzs
t5Exg8VKpii9PDqh0DRkx20o/O6wDnwLVLLVlKuccM7o92ckJAhXAr5cM+xm/Dez
kbyeSiwKL6p0/hBUFROWHujy5ccrz6r/RgEedcoCC1GfF6gJ5rXeV3ZeGhb8I7AU
L3y8cFGMQkfJuaJ4lW5CHL8Qq7TB1zaALH8FqbkhtB/it/TVnC6U92HmoZ3FMY+U
hbSukwKbwJ4Qd6PNCHbuCjO5w0fy3uFMNgZr0X5jZuq1Y8ckSWuIujGcjGsEe9Vt
cVxNvF5gNE5Tf1fEG4ifO9LZxNx8EudKi5HZyydkmlXRFzJJfVoLbTPwrfixuCer
ohCFkI2QG0EvlPUhRfOXSnVvZKy1yzuq7vYArgIpjHUAl+EAj/neNs+8v4Xgc01y
hq6X6bQlghAW2cvNDftnrFmiZHWEW0cmXSR7g2Hw6Z/hUIdZbl8XGTxBzcgbE1pc
pJ+InTMrkZgnoA1azr1OSAbmAcZYBgjxQrd3nlFU/yDfHeCQ35dce4Y+nno3C6s8
CL2bTGdBSvT6PWByTK1pQU055f5uoXVPkVZdycnBRLCix0iLSOTGsP60/aoPkKnD
oUFgHEGc+Y7jqIinc9pGxqopLA8eXl3SX/2luo5hhCV+NgYS2/PtfRay5Ip8DpbS
JrsWWyxBxWcdKoWM+V7iWwx/hsUAXiPW2MDHVuTlMkgi3N1k+97CRukZg+adqyed
xwjExxliBGksrrQPafDWlI+v4irPYBLQ8xy3HTkId1gbo6V2x8E5kLrivVsmrlyU
SpwSztn49L/pDHPK1PwQQ7Mf9A140O5LOsh1KJcgbYE1SXLOZj/7OlIFh+QHkfYV
HYODhf/e3BMFGUW7cmJnycPxuPFHlU6LsU2s16baJj1EMEd0m4TSjhFsZh14ddpY
ZIy3Vjr0jK7pUo+TGpSAYKaAXAMpHyLQwAxB5fhHf0aARcQauZKFtsiicO80fYEW
aMENJVCeopjaBRN+bsVW5X8htuF43/+5Y0TEjJjTea1e6ZdZMHX7LuVRUAEcYVKS
KhLXa9uEvNSbSijZMsqiq9KaAZTsvpuPcaP7aZup6IdbAZyBdyxlfONGHqmpHwYT
malRujMFQbCf/PTivOCGG7d8issy2AOdvmEKymZoeTaWThANdP1HwIfX1hwJHbSE
JS0aUTxWY0wBnkwEEqsCsGPavprEXF9eAME2F6PaJWAFoEgv4SZ19az1wuWZhpaw
HRLm0tnJhucK5tqcBAEmhVpSjV/mtSaPkJBpdn4Zm+bRTNpWIR9Gei/J7BqWbHNG
sI1wHNev3jo2DUcOdBuFpcmkoG7JrhPBjtvl8bssPW7mPrJMnXuq8/7w6eEmIEYd
LzZYlXxq0lDPbOcsB5fUMoX0p1vBVSlDHTuCVyGnlorzHcmndzHD1Q8wLiXkgbaP
Rl/RptQnvLA9Otj4I8vLAMwVW89kLZctChZhfZLBtHNnFJYMDsQEfNAzMFi4V+O5
GzLm2O59lt6Y42FEEFh8/QTHTVbSb+sWacS3yjW8Q0C3fhkn5vwohp6+TnLVFI7s
W+E7+1ZLacsZX3OAIIOLBnDp1KuFgdeO2t4nHkF5dDolBIk2XCDEigSmeH07lkQR
7XLlj5BZ6BswNXzOHPpf9apA1imbkpik7XZklBek+/ZHzwfSB3AZESKtH+MT8Qos
WzZjVpSNX1NLTZZoTdAnSnAM7aaWesIReFT6H+peby/S/nwwt8Unv34iIrO7g5n0
tqkhqsfNMlyZD0YfwuTzBHQvcau+V79Ct/hShKCWLd+fe6XB0rkMU9Bl9gI8FUXn
SS/VgHvgvh/N7/Oq6GnsZG7ZfUz1t0i55woWBoz09u8o1IPuHK3fI489S2LSn6qT
o1KUxrZUTeinfkcwUWSdYUxktZcUQjY3xlWMmmzyVyVEwjoDV0nU0g8+72WU7cvG
rURWoTJLqUZsziQTRlZiVnXMtt+sU5SxtiZYJuw6urucwh0WRB4s8kjzaJlIV/RZ
gkVrk2mnjNG3qxpGvRK7XnV5c7uTB2MJX7rMgk3VYbdfKxI562PdbJcga5aiRI2Y
kL4nlstgZf7Ok/QHwulbU5lT26Sr17YurQSBdy0GnuaMNkRQ36ue/LV5SMgRYz6m
RXgQQlCm9tc86rdEzoYcxgBpiNep5zpZfsy97OJ7Wk64+joYMwnOedwG2ZwE2o5e
64Ylutfl+m+er8O5s14sONWM4KecqktGQzUXpghjKe1YfuPF+vsURE6zD8pOCuHL
q5oVGL+Hkj6g7G11IYtx850RPuI4zjvIay0d3GD3hb0iMApNfZcd4tQ0ZwI+VeBS
gR8Zm8lmsaX/8oo8EQg+bl2fNSIQvlhbMO0R6cNcmOEP9tgh2tKGMC6t9VY0mNlB
CxCq9I6xhvBFOIoDfSGiXiKMI6ZuoiJfDfKmm6J+BgSTszzFvRvTY45y0Fe7f/Qr
Q0rzPz0PIpe/H63Bdl3hg8fG6MLmJcUEO/+ZrHlTSTMy1CoQMB0IudGrIlyNqLl4
846nvdOdlbK3FpVlooQFOkObGX1Ujgjl9hYfgnJykUiSL4rbunj25lu3rNwIpozH
Xm7Cgb7dzH1CzZJbyZUiy3mab0kJumx5dzKtF2JdoSkv1wxj8YiSsU17hKWnSftE
jJqvFgzyQP3VmbULfHF3E3Df38hZ397BYq2Ir3SfpB5K03du2xK34+1SLLnj3JTq
N+isIziX1IYpgNQTCsHr9BHB7VDn6IgFBap8ubRpIlIsNTGZYJKETdl4XcyaU8H4
eUvS9S0oq8WEzY4sX9/eY0T7lXMSOGJiz9S4wWQt5o9xgrcI9tw9Gsj9sTvXWKvh
p8eUb3Xz9Pbq+CCvrKEJJzP/hnN0ijBB0t870VfRfu7A5EWQfQ95NPQRUhcu6NtH
aZCUuW9S2nT97ehfWnwYM/+yLFQApSBopZJ4t+KKCPkLMzivkjZ6obUwh7GTnmPm
qj1a1sL+YK4P3PhHEqNUd2wNjcASgQ96mKg0K2c1gY5nucWAgTFH8x6P2RvxYBqX
uY/J5O2nLB3pyFRMPsGdwMvi8PemKfXTugRbojkk38iXJ2PECCSvVis3/yphWaPn
orb/lISghfAd/nPYIKcHp/CK22LR3HxAJLczSl+c+mZBEjnzFxPqsgaFvRrOWRFe
kc3+Xrm2P2aWJJVSBwyVSdwd1HXjYmqh92uA+EqHurap06fkk9tN/YD2ojyNJdQu
mHkL5aieiIoImByJGn0viE+rgQtgGUdo6ppnowVsfYfXDqL4Ljo89qJWnbalsgQr
4yTVDrrYN3TBA2wtISAdIOUTyKYb7v+wp+QeDytLq/tvMBli6EDQFHDJVMqV3Azo
CO9VIgaWliC8NL+AgK1paE7fnsvnmxn/QfI3JDGhyQHn/1wQVxaAWE0KISu8NQ+q
RMeoa/mkn28sRJQuZwg1NiANMuLfD3W5SGA9T/A1fsaFPnBxegOcGW4omXZb77xB
YszXZ4DUbqC3kOT80QLIk7G1MeE137umOFwrwUaRMnuWSeMwByhc3NlghZulXqse
bslVXcFRWZ2QOLiWI6wgFogxXYxLYw7nfeNLyF7kHglvXPjzVdh6csWS7Qm9z/Th
zt6M8LZ+wJ4K7Wuvg+BY0yicbNnck8Pl4mFF8943i+gX1M+1fk/NgwEIo+I1khDn
wGkulmclfIJxVpNa6sW/uKdFfcivGw3QZtPq6JwAyelLKgankE5cmF84yKDCWWdx
admFfAqQ10GizVVlU4qLAvI6rAQxSX13JOEHTykzQ1pKrKKJ72J8VyHVMZHPffsa
ilSkZdUGrvcQjBcVy3kz7LfAyS+rF3aArKIHf1GWelMyfawVIYpWMvCLSIVhDSN2
Qf9xbEQyQ/0thOR16FnswlcwOtjpAWIT7cDoL6yLQXTil2ibd62hTHJ4/mBEWHgx
QYEa5Q7nD38ocGHmRQesD5guah36gkI07EZ7IwgMclPvgv/cpn7mJanEZGp/PJrQ
tIbiXFFvJV/Xb/rRZSrXc/Ku/q0nq3LYt2xGUAxXV7rdg0hQAEboSIpaR5YiyVFd
4/vd78hf1dd8ZNLnfJUavRQ0s2lM1aQchG2Opfub1zrlEeMGzSUW4kJpSm/4tjO1
YKo/2vYOXFVh79DkJDt3kwanL3Jz9S0oWGPGAGO9pgriYwdBc9sd55Yft4lH+wQA
XwyMWHZcuTWiIZJDa1UjH/mEhwLkAzP8oslPslpFlYlxGDdxV+CpfBpsOFnc237p
OW6Fp5rckvqp9sHs4lRakdXVllQ2aYbvfE2ld/jDHLc46UiPJfxHP/nrILms+rk/
OufUxh+mWpyuIGKWpilk0RYf/+TXtgRRZsQMEHDCMSrp52l6Wh9B7xndHts4aYuU
REAn1k3bHtRcJrEJk3EnNgTli/PYVdCKuXasgcIuCyBosYzwoxRhTuaxiD32qL64
Kdeh49/Mb93P6Q1xhSPBFSEqb3AEqKqPFPmlKnIw9sz4d1RDmWdr0ABmm1nRjNrs
vSz7NeHcS6QM1I+0ZYlicA5YAz8EbD/9XrXckEbngJaHRjPAg0sUsqOWMRe/G+vK
0icK04YxWvIC4n3+Zewjd7VI+kxe8KR8jeQsS33g0LVzXukEWTw5TfEwh33ve9qH
OQ09vYvEgHIjUGNLCj+o7ypXms2IGTbUVM3uEspbmTta/0BuSy5FkjrKt+hFgBY4
KJJwsY1cc0TN7MZpVcXPYRvEvntDgXQkRx5cDx4RVbIYJwxa8UZ+cPnj1M1ttBeW
h3oa8lxl2dPfDKimVSq2PUU18CEKbzqMh0+wlIPAMnMRz092T0Plm0PCWRfUN/w6
HsjvNl+r3Gk+GcsIWuiQ48/OB5u9XZgkaGd2df4eie3ah5a2WdP7CaX48g5/+BeF
+t2j0I88W2wE/8X2Vhxdv6vwsl/coDlfpYy5EjjBp/RpPe0hF+OY8Roob05LTYu8
GecuVbqNMdi/RA6rXVN2VYFtSt37h2TQQtWLDQnKTiR4miAz10ik2VFDGImcp379
K3uUOXHaxoPwcYO/nCh0v48ur89jEbNIsB+FIT13V68JCK/qfbc6Hl8Pmop138Fv
qk4hXr2BxggxVpSSHaJUwK1Eymyv3khD9qmfS1d4iVlcEtSPxnFxt1n8QVkVenNu
JZ9Hxwj54/lW/O4uKT28YsAfe2XpFpUrf7ivJUzmoAfow1tfpfDeSC+UAJr8T2x4
kO95JntJY09wv850ZUopafjKXEz+lQgSC0E7sY6SWgHtwckkqzgN/NLBVxu7cBYM
chZl1dEW8reU+P97zs29kbN600QNCqrBB4TqjXlet1epjLMXHokmU+QlPToCYpP5
W3iY1tT4ohztrZsEhZer2LrBFFGcwZAVw3ihmPD+ugvwtIJH+yua9zNCE3dbzVE1
9kz+Kd1dAHt3avMfpw33s6bShlwhC3LymJgXAtwj/W0blLg/OET9N45q1Y/euU4E
BSFPdMrUd3uadoMjb7XWlRbI/WdlvzWqde1keJOiAxOh/MJ6LycZOX9o9P8l0EqH
rbHcNQaekTIC8WJH6nMrKwT4jvpMKv9kGHkUw6r/7hMK1hlE4lNLh2QnvF+qCMhK
CthjGQAFXdKW/5y4iuPe3cFDQLxjipoHzLItupd/eWb4/P1JY1ZjRs3M317V2SM+
EMW52mkh/R3ujqZV6M/8gI27We4Pqm0J5rpZOv8jF1UqNtuIxTmlFk41f8myKeuP
8oqS3++5o1taaXbRdZavhTkPgECDbixm/vm8z1eR6667VkoDRG6YFX47EvrPPBgs
LkOkfENowvy4RjiKbKWx8Et6eCJDHOak642vfLzMTSUV9QuvgDF9+s/BQHeQO8xi
LxfkLPLLJzHT4PPAYTUqI3IyETAGy8VyRjRaaqP1N/FNQj1OrCIvh0+5NrSpZtxY
9IdwVn5HGwOC2rmj+KcTWyq2CjvyWqlFpLH1uJc90kxoQmZBm7ElxjB+kchlQnKz
I2fYgbZCCAdleNXcHbT++ekVZ6l0ModqQWtjsQh8fLQ+7evK0SsKyLT6vrxG50Vx
LLPMhF5nFtytWuiPTOsMjzlajR6al+9QOUtVEdmKOcM2yBfRmFikBL5EVJM5aDWi
RvJqON1qRsCjG1UXVPXwkcbPBN1ooMZ+zpQyMqFVFlJWjEmwzFwkICRZNzw913cw
s4RfXXOUkxvQMR0jVUPWLX2OYWeFkuEdLcZT+CDrAi2I0X4QRuqUUWnTFIiu53uv
oqCTAIfQpHetENg6hpKRNnYRmbnmpltqhy4teOlLOUWaGLDW9L3lD6pNCB1OVviu
+uDvTbdqzVzTMJxOfZ6XvyscZeNL0emayFhMvHnOBJaCJ0D2jG3PnUwq5LretRdb
7C+Iq8zDldl0DkEA/6/VuBR4TuWkJiRxtSUKOax/Y5PrianoIJCxoy+j9dtkwLAJ
u/xUf8p3n5H7hBoJ2OU6xBqGMRCUf2KAznwv8zkURkvC/TwLR5/FMfECrjige2YO
j1hMtupuRfe8xr1wATy7mHzExG0XIZhFMJMd7vxHrV67A6vIeVZ8bMvAhYnawInC
/GAhjs6zkARIkRi9bLejuFv+mEBZ+Cay1KZAOCK/d8fF251vLVMu2jo/5dP+HD/x
zW9suOIBjoC8wiG/47Jwy8CR/2ymFEIfjW+UZenmUOxiIX4UZ9YrEG+HGxEqKt+m
p+eK0n3/NbaivTovVvy1My7ojB+A8DdHPhkR9GHbwRFeKSLj0afHPpCsECC1DCF8
+04OMskR+h8+IPXG/ZUn6jw4jV23j2E157dUSti6af0KLbV/66iAGSiXeOxtlA+C
jvkgYV4S52qCZTwk8uMKRkZooAlohfxVwS29QTOXgO5QAS8IlPP1sJyFqXFwo5D+
CFTCeC5vMF5ntQog90uLhPod0516fSos56xRxGNDF5w7Oed21umbC2rsCsHkrnhr
ijJL9ykk5IFYc3TtcfNgAbYOnY9qDqBz7liltyXJI2BtnDKcRc2LTedRlyEHw7d5
mFzdUYig7z2vA+3//fkNujZK1DQVVwE1x1YKaHW7641tvPFT6ZbpCFggturjgsiH
jzYP2n7NTD18TVZ/VCoG7n6BItLu3ICmRBP1vsg3PauC4spRkXCRZ4KXMFZ6xgVk
oOl6hTieWHMISx8goALUFES/9d1zwUwwF6MQKpxuieZbN1FI7O0mBkzIDrgU+gC6
tzukJZf6a4pR0ZTmaPG0QeYFZ1cqTQrDUuJ3NiHBfSmaPWh79k7lWYU1Zc9XUWlB
KcPd7jAmwfmhx1Kgbh86U2bXWpRF4zRcITQt2P+VNrfDeB6P7wOyeF31iGnAiwDT
yYOVchQwYoJW0yEulEltTeJGEy3biTL+n1u8suqjw+IGDO7dFkiX76ApJnzgPET6
4yR/88dJvLVXSNd4uTtj9EmOplaIsaYK270rXYNeXLWF/gOwVNS/3KnXQRtq+Y8I
N/mmwJjoMib9B7Sj+DS0WoodhCw/qfZ+NBEMPV/z8ZbvEyMwopSFeipsT2BEi1hv
L9Qnudl0NR72v9nfXQM+fdWObeU06wMBf2wevtsH/EzToNi81epRjo40+nGoj3wl
QDVWC6KoIMGoPGGOPyQi8VykoKIvUcKvQrCP0MKYCxBZwru/BVdkayrnACTnYFCx
xXVxh3mITeXaaPP7HaicEgN+PPdDDSfI7u0K8i0UYhYf6g+4moLtpWUs0Evr21a3
P66Z6Yx06q69QdAhu8IZzQXZwYbgWudhrzs7i+8fT66yu6D1Hc0uyp9vGXHb468W
qfAFs6xlPQR/dA7GzN74WqJt7Er88EJM1gQ1s/dZrwQdOTNA1p2VhFh4Nh/SAgrk
O8ul6u1GYX0oHJppcwLrzu627RJq4Hv9DvwOlKVeflEXY8OAan7Ct3wPOghB157w
zkJTmcxaG6CWVknuXpkr+gC/CODTmEYcTMkNr39rrILMJuCg5LES9C8TKkNJOuMI
1n35cr/Z8Q5M572uD6OisMM63K+Fs+jmDDi/5z7DBY1MBunFJTC28ryFzkwLmq5h
3X00oQkoK/7Ls/9DERvJjjSZ5pHOu84phwHL9M0996PNq3XdHueUSJ27cOymtf2K
NTVTBrPyu5+m0xFpL1zbqH29YolJi7sfhkFso7qthM7/N531QkRDjSeONOOethcx
AMzHB7cd/acqyZ4QJFzGQZdD4+5vwTSTwaPp/wXHpwxELwCrNE8kBXGsTxeL/MHp
kEGzzVFebfPigoW2mkOt0+7szarudLccs1KnogvThLn82qDg3z2jR7cj8JosWYBH
rQbYJnKHtJXFse0/30BN1iXq/5iRN8jUFhYlQxMosG6WdwWLV24kA4aDD9l3gqXN
UH/CZd6V+YE5e+7SmFE4/P1ZNgfYaRDHY8NFpP6CZvdJN1K324FTLafyb88uK1LK
DJkkKcTc6sST9AK3qyBYwZoikTIP5RBig1XJZ1A0xFxkVgLtKpXshoY+L3vO83Bh
ZkQGsEEPz6xRJzqNO+4dmT6s9/qiUs1ygw5pBeuuoEQIVlbtJOP/72HEi9cxpiDV
e5H8DbqcDC+QA4VhXtRaVwJDZsEkZJQ+S0xOiYVGz8+k1Ri6Wh6NK9iGQIOzTl3I
boj/6kDYm5yzd5NgfbTb6n7Yf9vXZSlSRknyAH9qhNomVg38MxGSzr9P0R5xPfUF
Fts5UmuQORa2wLGk8g1tZgNsBm+yGJXvgsUmqPPHXHXqyor4WcEPNyGL3zi1OFpl
xyrQZC9q3xhRHHWtNRJD0lBjaR6CptTdFsJ4h3+1LXePZkXYMrRh3xJkJ20b5wnL
Sc+DZux5gS9ETi46oCDLjySkzzjcyzjZfDbLMuYzBWCP18Oli7sj9pg2jig9QCsy
IOHYpNUCdeb2gWcHWAHVxlo9XbR9KcOccw2nMglfK1oQWSbfPTTm5rggVKtNq6/4
HNCNf7djRNvGM8s/riMsLX45EZbDQAh5VTWoTec9HQwjx4W6uQyyllEcRDm9+xxF
XOc5cm910vHZYgEQz/YXKSZWyArFBEmzVO4ma7Z6hoch1kifIbLzX4UtLBm1jHIz
zETVTsiTMk4IM26B36Bnw14/fsFHtkQ7yDb1NHbqyeWxdRuQUt5L7ISFMAn66Kvh
KrZfZeGkxThzbB7PvJGDLS1/Y00uag3M1yTJolxHPT3411irOXKBPi6rNSx/XYZk
Y98ZIN2wEn6aA1mA327SVZ7yFbFGtHwIfR1lIgWKdiGQ7f7+V9v1wah3d7iWtiqN
6gxhV5pAcXMfXWe1BtwUI11D+St6/gALg+uBZW0Jvh/IqVYGB7pcQkivxFEhxAYl
OUOMgl6cfR+Pp3gFym6/cpdIOJV4Ilx/aMaVmy/0tMFJpCDrUoL56oy0SM5Zf9nx
3MMwIoxFUlTmGbx62bftDnz0nZ5YAygsmaKzAAAGiMLam61kvfFBXL0G+SBLMQQz
olPogCTP1xCGdzJMOoJ1nogoQBT98jbVBcp3f329ZYjrKPbO6PZ+l6cuxjLPMvEm
VKqW4I/ypHu9vzmK8uYTD2Fcbw/uc5P0gpgEn8VHNKT+dD4tdW2UKKCNDMJ1pEUY
RnhM1ilMwXoARbVP2gjsezsHC5HjHcHF3kB71sEr0MsY6azm7xdAOtUfeq6+AUDN
SDoNur7tD/eN7eVfuKhYWM7ID0sMXWTKe2VjjR0RaVlCDh3snbEzJYBwXFsAGNpW
JFX02WgekI9RiwDL46FxeZ3LVR/GE5PZAfN93Ppg7BXqqfAkK9PBjFyiFcyCfljb
Z2ZXNqyVRiMQOoh3GOylkaSWnCRd2muf3hs+p+Oge41cxw9bio2ZzytwMYiowETI
Ev0fewCGFPd9kIia6W15OOoSHUJ9GYqaMDNwX3KYibC/DJweMCwQoyQFRbBJt7at
fuSfoWJjkT+1gUXwGZtYuqpwGwqYO8ZN/2I46nfYO7H+T8gztM/mTNZ9A/zOcfZj
EqZBfN8UyxA6UbL2n2VpXUR+53nDq0JOsULI7h+hj6Aei0Z8hyd5zE/DUvAlGl71
kaCCBwVQt2NwkvMIINRy0MfgOY+EPye3aKoZ/P+iArp/EjnaKiAqRaajWSMYjG9b
G4TqdNGbunyMV4LwgBaDRlbCmYI7jYCJdiCNjgUOGUFU/42I2/dhCIB6qMFAtecR
jLFIl01KcRwbD0JjugSwGBdjDIhrLglhfgiUxZAbz3fKMeBZ4HnZ8juufuT5+laK
MRPkgjHJaa50krdWZtMjzftQig5SjoDKSqIrz3W9R4y0a9eAFk6HpjWS/W4ATFLp
fVNC0aQPtWM+ekvbeyfE7Koyz+IbdCq6txkf2hBL1My4+8Q8U7lopMzuIeUJFiHp
iGxpqAs7YJFbBRk15hvLziAVPSsxlmqDm4fQc8N2dtZhmQ78DbeZquY/7NPuIzVq
tSrFm5EYfocNMuOJp/gjwRwvCd/8EmCuDDUTKiE5GGwVvqujPjh+NXccxYN7Cn4I
g4ihMVZlqlKK3Pil3Ugk2lhqFORpVKhABbapE6DA818TKnedsK6NZAMTHMT9cxEd
CLoLfGsTa9madT2e7FmL47q6r7CCwc7T0G9CMj+IUIQwfp/YDmex6T5k+8FmVTXr
NQzsqB/v3Bpwa8zQdA8na8bitdHkQKFZQ+y+SSWSWFLUdJzaCs2LsS6Y/4o/ouG0
g5eHJSLVtoPq/C/Dtgf5j4HUIaNqmxfVOsbenxxRXR27Ev67dxz3MByfHvvapp9J
B2pz2WGPPUKGTz+aT24ihKekJYGszPvDU+9856A8yWc6PfCdKmdMQQQfQcpapVXl
g9dpDFNqIZdNssafmA4790+yGF2WMQ5UCzobAdm2+WPUdXaYiuB6iXk4P3xs4MHF
bVVN4CRjyhDMQryFkq0zZolhdidIlEMLsUL1Dkk4IkjSCG5DH0yVrl0yh5k7qJQo
Cm1v5Tql5fbWoZFCACfnWEy95noj2d26+L3K5bZ7TZdgiHutaVLuRtpVzhc83A9l
NpNER9yZWRTXNs7Cx+E01M7kCvmSFQa+L/Lk9DR+O1x0QihwUZ0ynldJKmXbr7Sv
9fOE0B4RNw51FiCzXtt9qvdZoBSRbCbhZC85abXda+hcrYoexsnIIPRKHOlcmnm7
LwjuDXj48CQtFbfxdzdmxdbbftcY2K5sQuw/cMqPt+Lt7B7usypY2dODODoodYhN
Tqaqs3RkeI+fIP2mPayR3hvJ/SiXJtZopxYrcgCvPygeb80j/fJxcrCMYaCg3Pwf
dFbQY7p1xWBUCLDQNFg067fZ0eFML5nvuYsBiyd31GOMf7gpRImVjSMithvl34ok
iZ1ulyEsYb4iCAJN0ZJIWLLTHgqK/kSZkJOC628R4UgBshi+dcScKHq3OHR7cFYk
pL5yer9Q/MrCDxgW7LSVHEEKhWFW+IC9cPzoKeP0kUg1qzkmEoUVVD+CeDPjBoRL
AFXJHiQBbCGAOPmGHKEv7vUV7YyBjCBWTyl28Y3b7yCUuvzSbaq6aJpS2VU75Vcv
jvKgcCPS4o/ftmX/jSY0m8IMnG4UBD1I/zqi0lNRW4rCLUptHxoHpA2GXUqnP/CB
xjUo/Nwj0hQcKNgInWaY4XXETw9Te+bfdWGCdq4crS71mmy64+g9cRIiKLPdzPsX
gYf6Cm98EM/2FbffGvSPhoQB7b/9TPCmNH+kHvqOY0iRC/nvJ7oazrrkfX7jSKok
3kN/jSmW1+suFYTOqJeHORFtCOzafL3iVyqlm4wiPH1HVfmBAnLjUTX8FhJKUbKs
VKoeeRKC5vGWACl7RgnoBlqWc33zwIG7fjIK1wu4f47WpSNlQct5jOgvTWUoyoew
rq7MQww56w18+jdRikt2XtLyGQ4+M7wJQypRSCIZEAIaZ2H6pYjVBZ0S45lZFcG2
vhto1UZRQI/uZu/v53CuWVJ3N8/TD9U0AArMTtKdiBchRcqvrhERFONhwxfT/6GJ
TU+TKkzXUE10e3b5xPm9Y2BIH824/FkifPpXQjI2EMtL3uwWkoSjkaucOMr3Itwc
LCGuXTdL7GMT9NnVS/OLP/mS4WrBBgG4opp0vmy5+R0RAVyxMVliCSTTKX3EsqDZ
azFzW/IOTOCxrI+/65KeSRFTpSbV2/CnC9K0gHRHRyvXe38wnL8BJRKdsEbNFZ0J
qszXLNqri1tMhh0Zc0t7mKN7VWrs7xwALE0FNenENHNftGb1LvPvYB9Ef2SLSUgo
YsftTyy/jOiBdZ9a5O20v2Ebs/AawciJ89wdD3q2R005dBbJ04+ZMyONodWoFcXo
ftvDhd+z6ZY0337bmfYMLlpVRgv4MayrN2Zs78NdmN5YNuOjSaleX2Cb6UTAtoPp
WPc+hkgVa4C1/F+R3jeQdJe6LfrZnvk4Uv3f630Y7FDYTeHjH+F/Dxk8Zxchg3rj
CzFH2kW14hM2AbykgUl4cATsxbIKdiKArz43C9+a/PBMlNhNC5PflG52W2f5Xo4I
6RYMVBV7om5dXPQbP5x0jOQmQ13D6xB2ueuF/jfcFH0KbnOwps6Al5u3QvnRQPdJ
bkdiurc8s7NQvIQsJNkRSKFrUhRrcpA1it3H0KVFGaCLYhg/zd0l/qXiS5ZcnYK2
38S1WycGphYOTg+aK5/XIdzwrf3w9Kp83az9hfFxIoit5AiWtRL4yjt3CrAPEstP
0OSsV2Pl5wmiYUSMO70ruc7kupREzVU6fFwpZYZShu61O8pmYYebCIE7Zx/yL3Bh
+HNVzugQQK/0xd23IFTDN2usvzyRKRqfMuQB90jgV9E9EVS2xlDr01xQi8/F+8jl
Dm5s9OcwZV6txYZqr1Lsun4mIARxAxSusNWatGhMXQkdZBMg3pcK99e9fDWvw9Dw
WyJx8UA+W8Jl16KMivd9qiiZ83PXNLWwR7y5xMCdEtaJr9Ybhor/WuAYsf7soZqQ
ivB3zfPYEH+Ycsnn3Li+TvFXeIVB7ZisBdPzFLk6jphwEQpcO/E7SdoVandBEJuF
hBsyYVip48xF12RqXNiEPY+1Qgimzc92zhr7MxzsVWwyHI8hP7k7ADZhOzJ+U/2r
6AQiKBOHAIS9ADqdbti8gRJ04T45/CtxLI8xuYOchp33+S6Io0O/vp3YgLQlLPom
Vp8fqwJcYL71D9HLBtayg9zazv5DoVKz4FNotOpACQW8sM9YaTXI0G/whl38JYit
eGniG8eXAzc6XNMqxyqSIUluuxwV3JJBF8V92U2l1Xm0LGI0IrYYtFW+nIbOAfuD
bXuDClRHzDfsBNisop9MVbNguOkpVazuxh8zcEq+5X6MYicdG/Zn3M/I5ay0ehuG
SMNbPHniu1dy2PDdzHcjK9YsjuQmOvncSocTLBixy10SBD6eGG1oGHhUccblpwpo
7nXIDNx1UNONAy90ZXdvBwxVWfVmyvfq7nsvy1LlhfiZmTxV4tTnWtPIlKIdIKV/
A9xhPvz7giv75lV9Zrt4KvwZlTsY/BLFBZAVelXVvuakZj+M8nrsIO3PusJOPQHi
Bo8kxR5gYIZFMj7s+39iLY3KL8ee9TnBik+rFPoFRkwadcAR+V2G/OSAX/ycYnz2
TOY/MUulHk1OIn8LsY2RgJkzf8mvfqejiAPGEwBQknEO/pMRLzJYngYVEHhu2gDc
PLlWDzCgjG4J8M0Tx1C5WNULUO4otb3oTY8/1Bi8Qsfmv0rkmASdVR+rPXkVsbze
SeYVTHp6ZkVJ6tBNyYlSP0N6hIFbmvomXkLfCuIysmeJ/DdaAqJNjwRtFr4quqCt
koMoa194AkoDJTodLVLgPLsSyp2L7D0V8seXg4iCZPLmrR2CRdz+aGUxNzQ2CMVm
d+K5Duvr10IoeUmzUgCkL1JVuZX623sXOfNL0UudgGiBxHW6VCL93d0N3ErMD1y/
BfDZypSXrgH1NnmsrIt+4SbzPVH+8dH+R9Yeui+Vbx8m0e90EQXhlQl2NqgR8PC0
/8VneTR4bemldvmnlzcsnFOYWqtqZFKX1Z965v/3raagcexJbaRHL+pQO5ZKExZM
1llvxq3Oh43N6WXiwEDQchekLCCnW8IhkqYoub+lTynLp7S4TCdfM8XKlvee50FP
AMNxP6/0J9NCPFcopsb+pXMHlFibRbLZriV/X2ypEvrWpTTUdsBq9GmHhF37ppZD
tjaJuVhfEl5XDNTOh3Cv204IAkBRbqs57m+b64v4sfL/wDKooKvbQxSAWSCmpk4r
2Axvh4mZwpmane5IYydSG7tlRCXDyTq6VBMtsuid8FlV83z6oFsl7EnfsgJSc3ni
ZiS7eDusUxmSa/DamlfbxWSgkvG4afNHM2GGi24C5fvVWnCrWN9nKIyzkSTpBcp5
hJo+wIjYxGioYoZsQnLTshWodNNrDAfbSnN+5j2sGQ37sDn5YeYkSfPlLW/SzMVs
5+q2M/QI17uwqYCYs2IV/DAEQeS5Lv8BqlW2qvIHzy+gvLxV3DMLi+opAfro12rk
pAxWpx6ZfZMfp/vtGOUHcQrFY26/KlURAsWQDqSgI96lncGdZ8L3OeF2aSTC3bT8
ifntRW6KQMTkjdcp0ywXUTZGRZy9Fva5XuXLycgfGIku3UAgDCxF25rZ0Olld/DO
OgW7pXJBDeWtYpDZ8cwSZX7NDoBHT1vOBaFa4Kr9yE4POdWIpc7SxegULH2zGEOb
H4NRJmS9DasyN02/YRtDqWLR49RcPFFRo/zS0862vE3PSxL4qQGrtpN5jua31Vk2
Kw082k44d+GiWENKeVg1oZHtUNBsvcDGj+S7qcS241zgRK/NHKcMKxlLAzFc3X67
v0F3AsRAViPlGntw5ylf8xR8+La9VKxP9Ck/Ni03bLQVBBJy4tvTVJ9s69OrwCnT
dReeFGpTy/BZOkWg+2Yn7U5nCz+imooHGsaOlnUv9jdO99NpIQZFulWZ32R4ifGg
4R+V8cFqozyKaMnFe/ZIHO1RiiCWxRAVfyLQfB97R4MSRc761Ro/xedMMK6tScPn
EwafjPSbhLKM0Zlv3KGEkPXla27wPnjyuqcPaKKej0/uK2WTuky+vQwshSFWar/g
/TSCQDEBa7y8dVqKRzBl9XLj7H2RSqeZys+g3rDt21xMw5nqEXbwUgADMjZOhb3r
oIQNEL0Y0w6wjT2UJuDI0pDRsJbTWqwuGlkxRKy6zvTIclK5fKrRB9gBeICecZqQ
2T4Sd9gCQs1sugeHciOrTI5D4dYKbdPmhOZbJW/o2h9N4kuQ055VnTB2wQ1UxGzi
MKrLqS8UwsowqCWthLFxrBA8mdymnZbWA23sS46YODOx4hegFveq3P3MheHvCl/C
w9fkfkCprp/VsDBhIqY/gFiGf2ULi5qxL0dxoMn4dbzwasw9li/pymBL1k6eSAMk
xv2N7QZcBXvqGxWK9/9swF53TwHOLUf5JipcVhRmGq4pqBIEtZZYxvEpxtCJln40
ygRj81ZuiOmeX99HWlGk/KusciXkBF8cdC2oYCUsKtFZKpQrZJyYD2Icp02pnHGC
O2ubJKmxKm1sF1vhktPWkYRzeviRnsiA8jk9oOD6XQKNUL1s2a3sq8fkSAMyGvwR
RQjqhAkc5ieXpnclPIdsWRNdbN9QAGsULw6HBXxYM7X9Ri67a9KeGUsK3urc6mFW
uLne1NtVN0fDco/fUxikP75k//cT5yMwPth8nYs89GIuoy+sH9XorzaNbInNl2Gq
aYI1Gd4idaQ0sOrr0BVGZJLithDg0qWdDg7k5gFbaLjr9D6ulSQKXUInjZTNhQeG
D5RpJSMW81A9MSNCfznjpNPXprtaNfiI1zCcpB85CyyiuokpdiVtv0+bgFk0t967
rMZ5GEpVOi6jUmzdiJQweNwim4Xqb0tOJR9P44NqB3jqVuPmXORRuhe7z4IuUDqp
O/J9miaWmhrl2y8yTNSmYHMJVmJ4WhZpabJOientg9BjQ6O/HWt9/UrZxQF8SowK
BS0e8tMNEx1BCES69Te+W6vJUvbyGrl0KXciMBvTxnVM9at4bGmF9JuVuiHlT69j
MJBE70bdbr01WXltk7RzrsA5dJDmCO8iVTzRcH1iBqTbd7yD01ThloJydH4fH7rS
2udxsy3xT8xkLGV7eVElV5CUi7U7ZMV0m/h112B+E5jSYP2mekXdf2HMv5nzB1G8
0sapYkKJXmRE/tCNgTs40OxNu569YUOC/1dfNqo45N6cmh8HmpVSIxN63/4/hjn6
yb/1lxqb9SwFoz7hOzBaOQXVSjM8T4jbQaU+cOIoQr+B3+y2XI7364o/hzeeCru4
as4EUKaFtABLeD0M1CBO44YPHgO5vVU48cgx+tAup5n6GXQKREfME3NMjqATxA1f
m3pPHRFeubmK4Zm4NO6gt7m2N93rIIySUB0w0giOrVUTJKk8mp2XhyHZKRWZZX5T
8aRyIwqJTgbtOQZHQrmMprbQEBk3eEkFJF+JlKTPM7xUC/+ocQOC9w2iEmoyCXLQ
Ca2nZRB3Hnj/afNffY2hGGz+ZAKZXrdcb6+WHD4iTPUReN4xYLGSPg3ZwXs5i8hQ
okyT76RCHquHEFd0vMip4kcBvWJZ0mmHDlL6X8AjHJWqQL5JGoIDFsVZFmzX7ZSz
iF0aqdoAse97AlLYqOJjf8S+39vSkrOJ6rwh+eWFcRSBgLvZwiWK1BBqwspPBrQT
J2iE6B6OOKf3tss8UU+Tj46BpC9qUlTDqadCauw8ZNkmMmEWw9RzKCn63U/RY9Lc
lwoFIR9HLj0TFaB8SnjGgq6n6GbkcqZn4eD/Wd8dffbhf21xckEI2uRLqd6iV1hY
EUo8XFVYNihm4eeCdFTayWUr/iZHxvfZymOLd4ecT/+OkTLs22Py/ckdxI4P0Rsv
slWI8KCHdSLaqRMpt2NNWPseXfuhNCscvRmDGoI7jeMspMfrNmZaPcf3Nx1PmaSf
5iRL0vtGiCF8Bm5/MAh0T6UvwsMjqPUh/tYP9YDv/Vei4YmXAGmP2OHKnyevpaYj
o34v4oT8g+NuTGYIeYU6iuiLmSbVlKTJXsXjOWxsF4giBLgcuJsRlSGtlE1Mlk0R
JV9URwofyONpjmJURdBj30vgzE3q8M0PtfUACTGVQemB8KiXrIBQ6KoEAsby8Szl
3TtWBLIigbuYMEG5yYaGg9uorQHaFljXEuB/I4f3oY4NefBMh+eBS96j60Qt8G0Y
Jh8vkYYFm/yG3SgwXlSF/irDWyiKtoZRB4nB7yxP2Qh/zukoIFHzEsOV8/nH9X4v
SI+dMwz1iwXsdsmwov1n+6qhJ6ULnB+cD3sCDFWxRJVHjTBrvkLgYwNztT4hZcGV
1amfmCkUAKNdoiG6xHs1uuZf6ZEvgGz0CAK2nXZZA9ybg68qoSc0fP6Wzf9C5wPI
g/1JWoPCb7qcUDGVXifnrTg4mAGVNaz4Galt/dhR33doOkZyMTch6dXl7BV9Hcda
P/S5s7Y1gyWQFJEYcaRz1tjEN/SGf9yMUxeBn8H4RJ0m+SHLNkyjipFW1F0IqmcW
TxBb8qrj4RC6SSmOioXTSQvTXdsPrQXCqzKOofeWKnBb6YDJE+/uxz1s5yuGEj0w
4ZdQEVauMT6rir5WHaHSTN196J7evL+l3/Mix8bOCEIz5oZlJaL3ulRE3pJm8ICq
njdUvMYaDeBltHJa5K5aZUcoKx2XYxllO+7FnbU69Y7cq+skfigNB2ykDSdJbNIQ
LY+S8xJOc9ka7vcCGmgDmywUvV86dnO07l6OttVM1r/0gP0WSd6GxgDHYuHOfyqd
6BjCxvhRyF5amCMYoLOrxvFaO2tAQ+zfPa+yKQ1dls3mw8muGhDp4/gK7aVR9be/
IeuKOP/+0mbH8gsZRt6XRjmY2VIXj1vemz4onegvbqsphnCe70hCr29PsHQNxZtC
G3BIYtASvmsn8WRsw/butM441I3v6GGsoMZTu1fhHhRiZ1odNAIwliYDiamcjkpI
Dm80F+QfxWByeBAOjKMsbZs/fjJhUyT4h3AU1Dh2yDqTbQAuh0MlwI71AmCfz3y/
xiPIDAgEC7YVozDdD30/+HWKWKeVQ3XWMHHQ7vViZyArTB2tV1Wj5SA0UN6C8Het
IY3E1aowzhzoxOdS+x2k73LAbT/SL7f8a7pqL8pfp2B9dn2vZMNNHWb0em6WDU8b
hagYR+SykF/WaRVqiiTMDxIPcND5cgwX1Lkt6Hf4SxWyiydF/SteCI9EB2cUFIh+
fqrI08bW78Zex7Lk3rtmpMjO/y2hfYA9oyExLvUDbUgFJpfBe1N1lS5qOxiCBJEr
K2aW5bpUg1hUKQgULn3MkHuESf9RFziXWllThQ5aYrBUhg+8uf4gJhp4Vb0VFjOq
z5gC0/DsScQbX/Etxq6RtLaPyc/sUkcYIp2eSTBTO/TSeo0Unnt2SAeQpcaNIput
wuphIo4uAWnRppuMGtnJK6VogonWZWAP3KzWN1a0htFhumqq+gPrBUW9xpcLFacI
7NDyxA5g0g3Y1n42WBGnr8UHU/5IvehmuRM9Lz4l8X8dV3yHIdrJ9Zn9gUOhGulN
qL3S09IbAhWWe+biuveCxAwQ3rRkRL4+/yjZrrQAIxyy/5S+6cT0k6uknvByCNJ1
PO1qWR80ZsLCF9XDyyaYuEiJNMaJ/8a1QvDFzyuVzUWIAM95D7bUGcYb+tkPeY75
xaEU7O+VAEzYu6OJf5WokzJA3H2j/nVodPL1RWtPT6GlWm4Xlw2fosxtxF1Ln7fP
TR34BF9pEiuCSPO+c4fXkJGTW/RcRsGzJDO3z6RR2/cqvlE3j6dn7DCL0TExk0L7
XkKpElipGauWCnnOM1FGa0T1KzbQcsOwTNK3oAq2oWzYOilVVk6zLK9XMEmlMF5J
enraJ1+AKMLevyDp1LF3Lk4cwZ08T2VGaoJNJm1CX7Rj3ALj/SeLDwKMg16+4PiY
bOMui5RmBOsxFNX/DKkysEmXnAxL08bK4R6yJ77bJA9i/JTuNU5dPrJprIUG/ZR1
Bx0rf+uiCpTH7pD4w//dsfcFeVtk6MepUE7pL1GhprgLwSf8RMv6cL3SKom6+JWT
J2zTDAMPqzgiqLKOZYpF7FPMk7P/rFfyS1ZjNbHuPCYkYkXJD4kfmhccUbQ9Aa4i
p3lSjBEQIZ9DICKvm6SyOY4bAIAz+zYeNmu4hRyNrhkTK9ilTwcYWWvJFDyOekqw
zVELrQatNZJmJDvR0KGlP/0p1cf+5R9qTcl7K0cqNknjpDwlv11S+HoYHgDiMMeG
v21xhKgPqi+Q/GDeKDAxrK2e8DneFpevVSfw6aWdCkHbVFPu1OxTRq0nq6Wqk+JY
zg6rEnyxasrqpyhsgYL1zpRhMFexsSk8IIygKMHwoHQ5KDu1l3/WwicKAAlsLGuf
4dg4ufVdVPCZkbsp7R53Z4C73GQfshtjiWvp6jnat3YfCSS2W1Uuq4sN7nkVYu8n
nUsJADlnqmHzqr9XvL9A8OUlFsbgGcI2+FmQ1qU/RPabDrLgtp7m6I4Ls6SUkd7c
y3tt8Ob5qnUmefTwnaxMXUx/oglt0mZQhx9dimE2Ji8Md2WcmBO+SVVBNxWWpoCX
sxKEkhkKGYDfPP6x/0uvnWQ6lSUwloiibOvi8MZdXNPJuFDhj2R43byzmZfEyB97
FFBwRjQ396cugZ9IjdP1GGGExRg4xIsrNjPKB7LggxwYj5KiYaomih/f3XaiQYNV
jfkDkIGZHM04uytQjxmGgRmwx4uaV456GSnUXePn4CH6PBajRadhk6Be5W/PhKZG
wAzsPHE45K6m47BMlcQSFTmn1gMNt2dAEh3F18cyiYp8QU+m9pMUUN4dFDoJ6HVo
9bZaVk2zLItb2+rqmBomjVghrIy0r2GgVy06PuPFScvEC7sao7gOO1kKlaoJRHHB
g0CFzsTErHavcyKu2LbmOtggQ4+/iVHuHul6zi2wwrgEI7fcOsiLlWp0Fb89Cbys
WZKgNdnSyGeAw9tQwz683WLaB1QFL+02nPfioxHOcZ/yW7ZEiwYeVzBRxuLR1TLh
20hAon9wqtzyRdKfL+RcJyEN55jDYcgauIWFKzKeoeBA9pdTNaHCBodM3BKZldgi
rgL96S/QOBvJJdCMkP3HS8atxaomnZvnjEhjp/tpB3B5HiygdFmsSAH5aPKzin1C
hgrahy2x/Y6KT9Kpf4Yi2swd8fz6K0hz9mNQ9bHefXuuXSDnpN6BCgFiHkzFz/TR
/VagXOIRCHzqe49LH/NY1m3d/3K6UJBNuYFT3L3Oh0Xqa+KUX5XHDKhf5TBxGQLI
WypPCFDnbjH+5Ftf+vPsm1izTzBXW5ffpNKL17v+F8n7bnfH5tYN/z3986IAJi89
zF3ZTGhPE/YAzFvinKDNYbfdEwoUFNoFqFx5pmj1Iipx6eakvcgcQRjKM6fhhdBh
7IBy/AtbG2nEvSzy6aLgXxiBqErWP15lJLfwAsC+oOyjxCd98Pk+pHgQxk3dHeRX
0D6tg7HNMQPooDIGBnPgv9j3x75vCwseBNbuqKmrST9syjn7GgUItmDxerfxtwtM
KCODaZMqA0Tg4eXlr5GoPv/3MeL7h7fDAi+jmRJLgw5i2DNChrb/tW/Jazo0Bqu1
o6p3eDlN5ECWJQxdPoEqAlqbQYr3jcwFluRU48eLc9M2XE+vQEIo2SxGmq6UXSai
8sD977JVB28BkM+FeFxKxxu34ASf0aOpRWSqaH2UwvZAWW8wTp3s1482jNZG60rT
whui9ULZSNLULvzBvm8RarmhhHm4oVJxRH9MNA2G5SNDLzWQ+j1Rn+wEWPGuA1V0
ylZ9dB6Z72QLnQmdlA1VaHDGmdqExStEJ9XG2PodnyXPze+ATitvzIpSMen92cqZ
sCvZ7vKhnaPRN/GFzxeeyCJTwxNWs+Hm3ckWrc6I2KIJCTKZaxHttIXtYWrNrQcf
CFfUOLOWDN5ooCj+CPQMl+axl8BPYSx89Mu8d64aRZyJgYZodi+gxaADTcyo4WOy
wN0mHmhqziEoLod3jgN1s8n7CWkbHs7Nj23nV5HGLPGTj01FDLurBchML3tY7WWM
WiJuieuL2985qBBbBrevhOT/KUhmadq886PGa5mIKoQyWR3qscaHs4qctGOVBxpz
cIWsm83y2sUqIR2JOxsyz87QaA+nPjq1PjH7BVZSXqktKjSfpwbmqTSC4sh0/HIw
TcIEOpX08OkdiQiGDrPMysn2dXjuAmuHeVY3R/rwSnUfFofjxYyFydpxvGC8Mvq9
ZlxAXbeCTkNxqOs/41XdsP7tkHvNrG298t+AlFu7+4zDj5+t7tJCHQ704npBqk30
3YRf8OpbnpnVbe8V9nHxpnKHb/BgmqdvdXi156YVnvF3fxUeXdEviVwxO02pIffO
y/Yzpc9/jxeNkDsxzOdtUGnC3jQszxKU75DvEXqnZa7TPTrikwLL2O6BAeJgewAI
Cr6Mu5mn39/FdpPP/nHNDomXFDROKzbgYhLw4VJaj6EbTohdYVSNNho+ORe4SqlF
g2C+JKEzxgq/SfNPxVMVCC7pbS0j3z1+FPkj1OttdazQZ2BkKnkTuPyIWEvAfGoo
fZTU9keh5kUC1b4lalm49Y/hCdndW3bYVRsQy2FSzgSZrMfpykhxMxLocEYmVE8b
BHaD2AK8j4zmNm3y0ugD2X9e+5RUKwI5slZ8Tc2AA3alISgvFOv72xNgjGlOERSU
Se7wbj4PkPfGjCXXLXW89wyWOxgboOQxtyQKZoaZBtZQq/bYqV18xHmqkAqn4mzz
keKhnuq2TBDhJwxE+xi1H09fp9+eymMBgdwpIOKeahUwxoqxoWSrQKVboyHEMfAK
yvUrCOJzZ9RiFsRGY2EY4QcoDiU28DWRhPy3joNQ9e8YkeO+L6l/EzAXTYdxk/mi
mFhMCjlLn4+9icoLkZswZ5bGnI1Qn35Z45XOQiMwy0tYRlWCSyvcfS7F9Xs8S70i
/umh1oyHzcbXwnx+wXQfLXKZjZmFCnQZnAoMdnyHgagoberQqu0Z6GfvQM8a6y8u
NtjdHr9Srx6QkPi/UhH3xcSPYxK1MtR6uCAXR9WkZ/zhoVqAa1h3AUsqsZ0SGQOV
i1y7WNcG/E2HMzOQYqpiGINZACk4UCVSfhuRso7JDtt3YiYbj7FaZcg0Nfoc88Ky
rFMK1H0CfIAr1S56NoOH/XxDCvatZSM1+mSaDZWSnshAkjT06jWA9yghEyTjCWSE
+KYOYmZizl5k3g06O34KP0YSc6WCOAEV7GXpEQHr5bMYYEh/gEusNgSQnITKHCRI
kONoByW1U13KB/VdRVGdws+wb67+aojVgEXtuL2zdxszJmkHE1e/4WObV6clDDcj
0taUvXdMJeEYxp/N2m0jBcQkNr7LNCCgJA3P+/rKvHo8pim3cFW234AXJ7YwqwFU
9ETbfBIsoEPb6tuADVTQMmZBIYuEcHl6wmDGQyI4NiEMZWPn67kO/OA5VKBZQ8Ed
HO5OAfF7BX9aHqH/+JMg2biMpMawOAQiP4UnLbDk1x6scBS77nwTYICQpMMhdLNs
DiwiR9qf0MGw7GeZNnnmeHRjUTv9suapGsue8P8d592o+NbGNWa+tih5eQopFw1E
LYZiRTpPfdlQ8gKszlQ2ltHC4hVyP6DY8ucMMin8B7MrgD7DX7MoJ44MHLNCJSYd
X2bFNO2IAHZUoUx6VDhdGvwI4L+ciLEeFv8b3DuYIDLMUeQqeHdt3e1+h8rMtdnc
WAQRq3ZNW5ejyqk4Bsz6q/yfSfkpsAvVSg1A07hfi3VmX1vZ0zh8cxFpkH/zjl4U
AWpC71WyDijUjXw4X9BOXH8NIYZpoqB46XbRdurTMY4X94mabwCzoZBGV6Z6Vi4Y
Ee1oi+42YGMlcQFjlEcgdjZ5yDNwgKQ2dRRZ5Wnxh5Q+AVhlcbCI8CO8NtxSH3bp
/IeE+4awvo2ta3wU6p5LVYZfjC5vCDBnOD+zAJKX1W5Uo+f8ShMnLzPRCtEI/yYE
S8GJoEWJWAzSWIP0NVJG7tiWfOJaF4s29fTJz5bZlh1GwWeoD99GfKKgHcawWLIu
JmXXjU/7f7vs72BADGTxA+++wxnSbmhFNd9UrSHMu0Wo6gB0YkEkBYeIAuRb9SXw
ZAemHiH4MVURWyluEuGQqluH/9ZvXwnkeZSFQIX7u4sZdVAiSmcaGEeiURGW8ugN
4R1jXKUHrub+eaz+lI7UYWWvHCotXpVn9u6b6Erj5UMgbIRtPWay4RKJHIyd0sl+
1uKzZAS6hHiV+5emBPcEmlyhj8nC7c1BzI2EQXNKpyxhrn1JvulO6elfJZPKfKgG
BaTrwZMGTF5wW2Nn5lVtJcJi7qPbRIcj7ZauQKmjijnz4f5HCMdTU/jlosNVlZzR
cKRsQSolCLjhIjVl9c8kQCZyTECjNgI1A3cJer3BvwvXnBa6ptP7yG8MOVjfgHtn
h3G9w5iQaLLs4MY00ccsMhyH9DqNo4HEYASP55IZNyet0zs2ivVPIz2hUE3pj7+L
wgm/3UI0WC1D1tdARqluWRMqO1AuvODZexTNCjruQEa/zypIco3Kk1l+pBc1lyUK
j3AHa5XFGuw3V4QeEMJRUuxZoNQFEzkAlIudsUsGjVF16dbvmBQGjd0B0H3CH46F
RuAF0uuxcdXG+f9BYbdZMe0ef6xwMzyZnokdurIBiUEioeO9JdaCItGgHBRjF0Ah
iKUoxHncSvtOI/9S6g0epcw/9jdeJVdx34P9t+GTi69jPmOZ/+4EJUax378TwM2r
Dz9KZrAEGmv+l7/1ToS4++GjB9OCp6buFo4xiaH1Dwg/ccbZNGCSQd+L7JWnSvWx
9BH6y1TUuJXe+gRafo9NAuygBpaVilvETzNhKcVtBPvdQyvzIwRrf5/ezznt3Wsp
eyJAbS73nHE9xdezdYwopEIcJy/7KtCDnV/EuWgXFc2/pQM1Kn6WmkoOwH5jivDe
0eTonRhCAR0wNYA4oNITKYHR5V04zLHglS0n96FG9xYM4jjdhsvpjnUP8/ygZBav
vT2xJXvciKF6R6EJc+JeOKX0d8w4Srt98rdiKyHkzPe2LoUu9YsN9Q30H6pdQagA
M1hM9/86vKV1rKpqW+K4LEAWv54KKrD/EfO/ibf+b6zZ/NCkHQt5Z7kviRd5phIc
v+L03vBI9CB6/Rs2Sji0QyznCXl4SIBhRDGU0LZqH2jr0YKddO1YftBkDHpkJk+H
emImfwt/RB1WId+4G7PSA9kwi+/9WPNuXazA9nGqXLwQP/XvTVVY8AFQlxtZq3iB
eVOi+t9tj/fgzKqCnYR+34gLvAHmlHcXS/Gd5nzlWC0cr63hh/B2PwZYVhGJn7Y7
Z3ZkZEixRphZ/f5d6X3fdjtXSTqBMfP8UPXUbZeo+X0tQsVHukAgqJgphd4iW7mG
1/1n6Sx2O76I6hetSgYcJn5kQBj89adoxZ9QB6tx8BMle4h/EqxSQDF6gDxO1n6L
qc73zU44+mu605NkWnzGBRGUKkS97Mx49FRO/tPZscXnLnP1ec4Sf1pars+26s0t
oVQu73egl21W6G/yewrZn4DDmm1WQXOykiMtIpyqhgF5H+fcdAsjWLBJD6SvRJXa
T4CZfA5ku2GEXPZ/LEAstAgsFQlJYhFfWaAUdHAB1OFnx6u7ofk9RzSB11Df5XfS
8UM1MVEebUY7AyxyWqy5oF093mc9hhH6OuUb1XcXeT7u3rAGgA9xAYv57gxEg6YH
/c+5eAxDrVEuhgxBFmFLW51RGkDk0Q0B4IBXffUGpaeXmydDeewf/jHB++dlnaNo
F7Xe2MT20BKGca+NMQVrnU/Z9F8Z5Pf3mPj8YO4c63rqA+8kedbcWZeKXJ7qqcpM
0HTaQVwjSWgMA7PHGGYXvJD8e1YPJYqIKWSCYo6p9ltN28q+zW0qssARBF0yhM0O
Mx9nscv8RTQactfTsRNG1xy5yaekhWOQYI+9hKIzQMuB49I2nseL9anNRsMswIEq
SROf3Sc8UjLHMTh9eQBG6HUiUCXPHZiStTwe9joj5+e9E3OeJKFJHKnbdKNYKLMx
AdhCRuY/ExaJQDVE2oM7PcX38LB7d61rZEfRuhzrlh2jw6N04tGIO1S4TLimcsYt
dfOR7JHN3qSbMJGAzHR9dSBDK3hKAhjgS5OqcZgZnYRqdwl2gfbMDBpiO0J1sA3M
bmODYJ2++BBj3BD/mXg/qHwnMEhLaHZBzMbb3tN068cwp0lCeWZsZibOPa2S7Eb8
fIjb1fbzl953lVtTGrTUIXibINhtfqaBlYbTe3yh1/DSkcSTEkwvml/Y2sxg4k+n
A7CbDj7T/B4F8WNLc7KZTEb++MAKAIgH3F1+rE/dtQ1HRiV4ic/YYT2cxDMsU3d5
Etn1UQ+HGQTm6+RQdwHGuRyPBqJcvnICOiZXNW2OG5EW5DrKm2hewCK7hQPMEOZz
+vcKlDPF7vqSTkXU4aNTr03e7HLiNN9P3FED2Wae18cA6NILvwJCmGmA5w/cPb8I
fRdvok/CXXkcQl+aJZruZYjj8lMQVhcqTtXGgJrxByT4o9QCfGZ5f5AXqVPaSo1A
pWrjYMVwE2fCpU1HnYIrHsh2XFBnTrlHkeQOXyPoBR1aymbCpBSTkIlbJ7HLMYCv
i9cbfZbddQ5GBcJuGUobOuHILLHjxw2WCvtX0KYrKMxUYcN+YHB0EwZN2fNZQfCI
I8gr7hwnTfqk+aP5Wn7G1siQQwdVp22EorkE7ys+TeMAuanyFBJwG37j4mTBt7OB
L5K6xJh5yLPcLUWuVimQfnuXaMdzPfYDoBL4S9QKrSuR2HJ4zp7pRdkkDDu+Yzvs
soCeKfWvYWXNiur3J80gTROkidkdJbIH6YH15ARJul3I6/e80DOV4TiHMdBTQyCO
ghZSAiAujGKFXzF5G9fuc20STbzxnsYLJ/+vAUYDrtr4U37xnORss/7sVm4vFiFp
yIaiMUZFFFB9n9AYME1xp4cHig9QDfy+8AF9IpmMQYLlUtKjVezCumY3S7tKB9PR
s28ZAE21iOvdLHIDsdwKiCGpHruQqYUOS8WCbqfbIBU/czuV3VjHfE4fBPxbvPql
QuK5its2k+L8mi9hrFEWxfhaSpgGC5GqCDnPV9uy/Hu0YLxP433bCEQOcf4WbhAb
n37z3pkcyabvDkMMiaVMdZj22JvDuGXeoNyuT86ww1HqJkih/LNowG3TIsPOY67C
QwCnox0+vEJIAwEW6Ei/YTFWehWn5RCXoGMrWN5gmgIu32xzqvbERXUiO7ODDy1b
v+34TSN9G3kr6lWW+Apj7fTkiu2XXbtrunba/1m3B4OrvLnjPKdMikc7yTvRIxEj
/x1kNiO1OpEmnXTi0ii2GRLBxMCEqBWQ7/M5fkIMve9pV5uXMF6noOkM7q8yDFQJ
68xalttF3H0RUH+vFOE3zvCZbfkturzIA8O2QHxTq1v2WuE76R5ikE7pFJV+vZ6p
WE631egFADKGCKxg9qFLDPgiFjQ4ALMnOTprFIlG1410QHXEvoOhfSuVREgLwwUv
SoT9rxfE4CZV5/SQjon80YK986kkPqirsa6tJpcxFG8EvDwbsB/8asJc0PF61cK+
Xf99+c5dV9+YxFj3tlTFVSr5WhGcR5g84PHztGKfjN34ytPs0KUid9BAKVzBhhX9
6gW5wpHcmqwuzkhuyB4R6nYjFlEppKkDq8TYzPjsSHv0q6mkXCh3NtRr7BQ4XTZY
rlhEWEBjkygBtKN0hwKfhepeOF6ULjr8jA2YX45t5C3gna8KWCuO2je7eQpTtQGU
4J7CXwdDhOOo/jIrpvThEiYwAl50wFCQbo0I1qHy6oDFrfKjyYX0mUG/HVEJmnBD
bxY/uUAzfR8QXTUzan6JGWwnyKK8QRwSfnKIoNAOmtK6IBx8IhcfhqNg0YzIeZmt
6jJZkCHH12Q6R4aNEOYkM76eOxahqjFMxZyUDXQv5fPymwyyeAdIy07Ex7sLCXQ/
fs/gbV57zXnY3jYgoZBVg0kqOPgYNMf5Ox3Jg3njwcfXUfpKvl/otaiHO5iqB4JW
f2gZwQ+3MuhQ/uczQNkwMYgxvG6eZJVb/pqiQNePvypoQv9cMPYPIVKoVLoW6h3I
MI1M8WWJ9Mf6u0mutSfyb5SWBuwOO7Rlnpr5/XYQiKphzeWgarxQLE4xpmQvxLve
LaHjG7y8+tUKdu16MhxRzqLlbh3FvlXAF1//s6kvnpwBnDDQdd6CcnRkyAuMKaqa
2VAaR8G+Mm7RIFuhZoDh3clyuA8NcWPS4TFzkca8o37BzZf1q3G/K2QyJj1WMqLP
BvqZtjCwxgYv3Bw2TbJO7xlvreTvbSmeJTcBUWE/SNHeqdhDNmkohSucQnQlmEi/
cOWGxA4LAqoQ0YbfmJotRBXM+kLAoKqy+pLP15YMv+rH62ilV4T/r3bOWbg9oEr+
Kn2NaERnVjgZ66udsRhiRSSFJKxSGhYJFrSlrvvOhikP7C7bIu/f6SPHpvbRCC+z
1/KQIiPiEBAUc9I/FI494YxoaWyzKLX+4cVvpf2dJAWvZUljxUQmOFQe0ujA+tFH
C2HwTqSmueON8rSfLKcpXYevDvtWLZTKOGWMtfnkSu9sSgF+Foj6uWVcbdCA7PFt
r9aH64fh+nX8uRTqH9unlV7hqlkik93mJO/l+L5DSNrvryZ8Cy5nzaXzlyb+f28m
ihN2tJdHisATMynhUbyLnmG3PW3KmKMUBYXPdI8VOoaoebe13Pt5El/osQ/UwKri
zH0Xz30XolXnNJJX4TJGTV5eqWhmXTeoHH0jJdW9oLEiekJw/SPdvMPKSXNMGwzP
Hmlqzg8DCAqliZZw39pE6MYwARu987oewUlZ0jtIZlKDbA2bTzBJzphCt3zVTzqy
BqUm9W6+XJEiVPk6UEeP7lFENwnDBEQLVBL4tijq+kMyA/VzYcEACK/j83VuTeRF
hJFanqNEUAeiZLrubXa6ZpJFdK9pNUcnMqAPRUo1dIC+PP7wbXYh7/gl7y2OoZ/W
33+1/hd3qVyOx5CLzF55CoIq9pAApI74YiUrF+gRK/P8KPdoilB2JMzHuxp5e6ig
8891RZ3kiGlyghV2MHZqd3R3UWufrNRmqNdkk71M9fPkkGcr6OgoVQ4z1QhVZZq8
Afsn55jwDLoSYj/uhLGe1QGa2lccIx2p+/ZP9COHB5oZ8VOSK9NJgpQnYg0ZqZc2
GDWl4prSbifyYs/TI7XKBBjmMEwNwyKbcS2XNdkFLu8KxHcvFjp8SqMPbPUHH3uQ
p2qDgcuRwKTskyAK17uSs6lEVrCUYLd7dEhjUpN2dW/dHdOBVns/J/SiOKqaLEJS
2Io7Lp010a5oYqDa7eIjLSq4b1lvz0IH1aq6hbmWUQY6YaRALHlHkpFgGFh+BneQ
oXYhWed58SNXVdgOjVl7b37U8KK6wcryXfzYrBj8IXnHzN3TzbkFzzfPwnryzdtL
eXWbFL21R5kdQCTkK7gmiFA40nnyiqcfQ+phM903KimZOSpQwi0pvdEotACU2RBr
Aza+irG8f+SOvmedsTaxarFFcfu3TbFkgQ+5qlgutFHBEXl5aO5Alf4I5Kx0N+WM
FkGrGXLWq5u8k3xnG9CazML8TFXSAwmorwO59/duLCWRjby1o2yPh9GHAhUZFBIo
EfMnt16JqdERHI9q+7hRjCzX1GMo31U6MFzpnXab4XWEhD5kGL2Nnyr7XfeL10nO
SPVd2MJa/lbWkvZD1m9qfCsWeM3V4Q4+2RPzjLFtn+gbr8t5oYCCDN2ispOJUnSa
9O76YnMMcSPcE/EtF8xEpic5WkEviChAqMeHfXVc8lk4ES8F6JnNXCRyquk5iEMs
HVeOE2HjBLtPhw5vsaFIksj/bYX53T5bUGG+cQ4hLbk1L2AMXSsqU/0qb7Y34tq9
K/Ie/hpBDGhn9oLzeF30FiT3YTmTSHi3nPMkYUr9NPsiKSXpyMRIzdUhV5qGyqf8
GfcbJVlZSo1Svh+xN7H3OOv5oJLrtdcYPb5DHBXhC/fh/8ZloWX4HIe13bxiLuHz
r/i8hQd+Afw8L/PJVL7k3ZY7eLjLiGinB9XUadSX06PGYUsovQd6O4xSJJSgLx85
QyAKNg2YFyV+Fbzv1zB1cv/k4Wgu9D2EHS+JG2+gaRiAYMMmyfkQ88FeN/vsWRMk
Tg6HokL0Xy2VgFLGkdqmUgsOeLSXFl8BbeKmQ2BfFSEB5qwt119aO762BjPzYZN5
4dEqglgPbYeL+9BYqt9PlsbKXc+HOOJX3ZgWTcJMeBJEvpmkYySV8ILFT6WY3xxu
a/Kjm4kMt/ARWKJgU781SrProE+wA/2rxY/EHLRFdCVGnt+8qxwtKT77ntnEuxR9
dz1tC0uK61uMi0E2NT+sTGp3TCIfTTX2IETbImpLK/40ofkwsCTuZsFUEmAhKDs4
f3UJ334VsqxDm116jDHMVK0WWebuaJXQzTVS6oxU4YTsWV9OQ2jD5mzhBJxEKQ4O
BRr6T8n7BMjj+PtFjE4XAuBBchzs86jyDnt+on4rb68vVm4TcWeLGirhsMQIW15W
G/jHQZ2d4dq4tGVaXJ3RRazY593A29bZccFEpOyzsIIYBoN2RGYBc2MuSQjdTdMo
UGQ1YQe01V0ALfvw6hPgVHsLlevNpbRcDCI8zaA6m0WBx5SSfR1Ll5tEho+Yfyww
jE9ISDngrXQbDjVX+3k+k/JurnTGDEOBfktgB8XaEeRp0MEcY2G4G2i1a2H6udlN
lThaXq8BsAhf6hbP4n92Bbbb2ugcSmZC7l0dGoisEu6DyY4nFHpQ38dZPXSzroek
Z3Kyy7IY0B7XzsPHDr7uq6+VqxfiVgBL3BbIU2UxbJfJdffO5iwq1VD36mp9IZZs
xQnNHl8hM6Z8yFi9JbF8Ma7XYwuHtlwpDn8CX/mG1nnNdpcfEhVk1OWRwgb4zhRD
xcn4a+FsrDtXwWdMtRb/xYVe2DhAsGoeK48+a/53CK3PYIthmKQTwH+/PQskOfM5
ZB5BtSGuO556PrlYWBK7UXDxm/ZtDrxvnTwe8kDKC+hmOh+5NVROqFLIY2z3e5h7
ZK7Cft/psiAlrqQXQSONX4VTPqsijfGMw5LV8W+3kbxbHOErVsHjrMkO4NwXQ6F+
ULXMkkbxy3jzGKef7nLCA9CF9jS7MsGVCuuxkCYlK9hc+fwArrevyJCHX7Qe+uOy
GdQGkRBT9Y22D2Ysq8+uLBPGhyOiJ2ofmrxyhaTzF7s9oFFuokQR4FPuRb/665gL
zp0Gwow5JeZVu1Nu7TpVxwDuR+OnH6+uY4+FTYNqP9f1iJJCbGWaRzXLswufpiCC
xq1t/xy8UkSl/O0w86Hh9TLSpSsvRd54LWcOHVTEnuCk9KFKTlQt4GnipKxFNZyr
u3c2/+iKw+DBVAFoOw4CxuHJtLnUPQ0x6oq4hAmT6Sozk+n57QIRJ+EHe4V2I0cn
rDrX/d1HEO9kT48cqS0nv79I6Pla1H4qUL3Q85I+CyCwDFVhtPjNYCfcvxcIZXTS
o049Nt0GicyQjgKhR1m4zHbLaQ6Uzbs5/69ZMxrkyrM+7ilI+7S62ya6WOF2oXE0
0NzOx/NlTSj38cJnkg6RswJk4zwbU7eo//lW0RHX9wKosRFjLxrtYEFyKIxPqXPD
cSahrI/vnt2S8pEORJGOr0R5oVFIm4ddYMThOoOXxgLjuIU2WRg8gibVBMfelmGu
iKAHbjxzjD+Q1jb70ovIrqMxrcekOfWclfNLPm0UjpJyRZMm4Mc1NT5Cq54OxHMv
qEtaG8ghBhFqFIa4lpA7lNFnXFgBItlPrkPfXihXGg93pZgQdj9qMvdSRM3AvwEN
+k9X9v1B0Q8ImH+gwM5CJtuYSLtrEVTgPgNTJmWmTFTuuQBt0XTXY8HX/XFZpRRU
jjo3ViIRv/1X4oYQbIvSsG6Xaut7vL4I3gLWmAUWeAfnyn6Yzqj3MspfxJ11QwS+
2sGSTd23olioOhkUoxfGAEa9s1kH8p86b1KNZ1umB/tFHtY+yAgBOSP0J0JAEQ8R
lV33TRY+dG2AlGuCqvGClqenBLrvn0w1y25jtApHAPbm2Dm3TiYNS4AKrVK5y37x
xYM8ctGOxvP1idqlihGBSO9W6GAdCIc0GMWPSax0MG/92iEKtfI/oNx+yK6PqJh8
tbgXQFSp7paw/DQ8PlE8o63S5kx6pD1zela0VKIU/NHI2Usi8aW8ae2y5a2WhtP/
3d/OW0BcJP2n4LXGKt6NIvUxUS2I5cbQD/OJYr8nngSHQm0ZCCcAvqYXPDXlh/s2
H3Sr5ipCG/cStZ/2g+ATAT+vPgoM9eRdjwcb7tuj7CCcOqzB+OOh8rtuOHdKm8p1
52De2Yh/WSx85bunwszTfPjEqOMeZsZZAdpCjKCp4pBIz1BAKLGj9zjxhy3S3RwO
cReT0TK01mChWwjvGD4wgyVyb8hP/0sSv6A3Xgr0/HYtFUhjBa6reu4/QSlpnR2T
wUT34QqYaZyJKEwsX8KYHkslaHOV3MvGUFbWJfxPC+FnvB6X5X2BphE33HI35+HE
vfdakzjeQfDJZ0eBXojWd7HnLMhqV0dExiXkuAypHbd+0LIXCc8/ZZUoHz8XlvOU
jEO5J9In/zdqbg4NVcD/C8o5Fd8UafxaEdJBrnZ1snZhLcQnCnyTE+7oK5FVrDpb
ENMcMH8VZXFnzgP29pRMNSwVv4dmznYok1RibWD+goonTXWX0aBeUZU3YRAZvKNM
kJ0rcRw5rLe9OBhaD8ZHmn2PfsMkTfYzyjOTmR1KTMQHBxxh2XHyYPdDT0ULniYV
WjHCAGTfqUl4CLDmadfWmGhzDvqyr/FEYPWcsXnYPOJzWBmED6/nYWHSH8YpDLAP
BCU5v/7y9JUMkXK7BlNJzJJ7XDcztGHJGtXNYV18bKVYePsprlQU6M8KjCP8i5mc
eIMe3uQcRolBVqkPFcATErhhnUnVu69648lrxCLABkqoKSB2Ob49EcULKlWwX47N
oi4BGNTDLBmpGT5susn9TMsMJjAto5zgygwQzOSV9SFk7N8j1CV76Te0hKUOb75w
392uL77jrjzZo3/KgLUIvMAhIUeeFF9UUd8FrgTNosiq46f8KQH7WLXfKqx6NJbC
xAVZDzUwzyPosVDfxyJCvH4kYvGSYp6+6GzgLEy6ew/LzikUT+tsj1OYp6ikR72w
gEY/auVcsH8x0/anhiR9WUH3tHzWZnkmCnFkn7FfWyjMHZOwmC1PKU2qzkFdAMRg
yDGACnSgQmRMFPtFGF5q/bt1JU91fwd8KDCPLixRW2KXU5tvX/rbUZsK8+GU9VMz
HduUm8RUADAFElTcZ3TtIgoGqfM6SptKndNw4Z92Qg50cAcd9c/nQsN9lit/2Lfl
tR2SeM7ezUclH8CJhMARttZu0Kh4wOVqQz0GPOTZe8ZvY0Vz4m6wUuZAeypnZXxu
/MgHMGwqmtDjREbwOYvuJx6gyiO/Q/bqtEwwwdjNEeCHT5U3sNYNJs1h2252fvYu
Wfwf3K2dY0YWp4gnnKiLGuVU/xYFDmnEiqBCWwtQEcCGjAVJlW4Tk1AXeiSmW2q8
wpTUFiRps9XCQIm3N1EscEnPqeecaukYWT8l4c23JddbsSP2MWCL80vgLdka0+kt
WRFhOIkj4hVBFpATQX2QZUbYBLH/U1m7ilf4e62TYT/DITQrBrmqjgWahlHKtPer
UhpwqlzgW0v0YRodhylZxsBOrNlaZdSuhP2OAob+jSsOfbfldZpS0+YK85iunvTf
+1TQUgIMjmc6jL6Mc9YTWf5uoXrLYKUHkL67GaFXS2kD/yghzKArWgtjcZEJAD5O
05+oV42mITOZqnYt2Vt/YOX3MN5oQMCtMa5xZ3MJk1ahDPBMSY8uXVvkm4wryk7M
6fOwX2ysRxHEb2/Ep87QZG4CHXNACRQTf15eOHTsw9F3DaOl+Vne77Jw8GgkngSQ
GM/iCr4nCttHhadO8eOe3ZuU5jN4OQXPJepurT+VGPnvPi6PmuY8R4G+UtYvGKn/
nuHj8mTHnW2V8l7j43h5A5lDZVXGSp2+TwIsEBRAgPXmzIxPyfVtMDtCQH/uUXt+
Ki1cN9ZDFsy4Ao+XWJfSVTOO/dD1vdwKUXalL4Ev64XQMev5H6uFqW03mdX35A9b
gAvfUzqfhEE6X2v8qUChNIt3kgftRgegYLYfQQVbAs9D6S48Jz5xgMM4obRgNx7T
q+5Lz0i5ZSIMUVwpVQ/aEABW0Y5bESZ63oTWBGZGfkNS33miyoVtvfks8pnWCJOJ
0ia2p31bj5qMHsbcvcXteRMHSiaO3iq0bymE/x6TYGzfjG8+Vz1NH+A0HmlCXMp4
eDelBFdmegUC7iCZZ38Iaz+XuIbStJ3eHeMSdCau65rdN/S1rwdiRdgiBJl9HNcD
MZm0P7G9Hc23PwU3YAHm53Z8WKSv+JR08+6rIPCjGjP1ubxUzf0YD6vjWY0zBGGn
Y7SpzigSFhD5GmiI5eX6WEVV1mKD6aWESXL7Wux3oW5rnGitWeT7l8GonkX1I0ty
Dc/BcPUBGxE+QjgmBFRjBF31DYjgeiqqDNyvC9lZcYa1rxyI0vDQQAMhHr/hbM14
ATHftW+WqA38cWp9poQppD71wm6AJEYiB1oEh7QzHdpVfHBdMrzBEytpz0s/MR6u
l7P6yb4EKXfwGQWtSUJU+xYHhDK7n0FH590XUPR6A2civerEUKaDbnRpKm08DjTr
pID+CQA75KHOuFR6GWGgGbDqX2GJeuXLZ4XLpvjeXoplO3iUFoqu+YaAZq0AvM5U
XWlp29bry1VDRBi/70gATrF+lVKQQkdj33SRXRGfwYBCoHLzevLa1S9g1+9lLi0N
OuM/60e/tlMHUhD89O1eL8c38QfjUPThBPHdX6eaza/fcRWZx3tTXHjzFDMJUqhr
KsrBNdHOvAykvDdXi2pURTnnxQ2SF6p1v0c50/nAxs2BGHHelshAIIA+6etnVuGe
6LqIttvBO2B1xZWPWb9nbJXnO7ViQOKE/9/5zHgf/XR+0AWFoOpWTcK8vPPsPH7L
dSxbhgQxnF6CqrDYY/2Bbv/3bFgTmpJS95w/1y2nWJhQ+XXwjJSTMpwOZA6DZpPl
0Fniz3dF7enO7kpv4KHA8YaJ1p3a7l6hz407JIFkGMwbwr3LZ6gU4BBbOtFHGQTs
JfjJUBtMtpxJmhg2oiRZxmL21NIOwIAIvPleY+8V1n5mC6pp1arJ9oyIGVmjDs5M
qzcFQvsR5xlzlVbIW9k9na9f3KiPiFDPd9Re1/CyJwkOdt5yojF3nG+JstBMswF5
AfTWZA44t3kldH0t9t9h9ZlA7DBDI9i5ullFiw2Nfi/nJASCRZ1+g/kUvrXVNBiH
SUCX9cYyCh5Yz7j90/Fdh8/s3jQRF0iIL5FbHq6pU7fzbohe0C0zF4FmrT3DB4pk
ZHMSxxyL9OGppAGwDYMBEtFjKy8w4zVoJH7Q922O71G/i66XJnse6BwnX30GTTLd
y8lMUfHlnGgToHOgHcn387YUGa3YBa4CiQ13z3mpNdy1991a2epE6oVjpKdZFkfd
yz8nZ2eFm9vATVROY51XhfacB0vst06zwaSB7B2/ugaIsYsMcAoAoP8X++oHdCgC
YySAkPS6Rt0YRD+5eBAJb14K3qOipOfiu9XkUdHKiqwDcibqDI5SwBFAzgGa42oD
yA5cIVUUMDoxhe6uBKuwe96jVV2PoKI1C1HtkxKz3iFyXhgJ7xGPMwI5DN5Um/IV
iuajazcwCYgSHtnrxkzax9Db7ihZt3MJjxMWEOL1SpnS0uSA/yxClNa7Rii5mAph
Zidrlz+8+oQZzXTZ6PJjqiA7+AnAMCoM5JkTQcbwLls25C5OR9Tz80+wHu25XuPw
EtjLuVdsG4D+1ibXgKddtAoNzgMOf4c8+SrXUljlm9YcqK3jTuvmuBRdt++p5bi4
LEk6VOz3NNQHIAf+wfTUU3YVz9pMwgm4ZmMZVE1Vb8arRxKs1147/qbqEfHW1VT6
qrdN3PXblVVoDdBRZsr1opY4W/8+3GKqY9sGJSKWpw9zAs4SFB3NdzSAW6maPww9
lhgyaSbJlQ8k0HiTv0WbuBuzH59Byl2UagRP3ok0eqbFiEcxiPKYvp4ByFuzWpig
9aJt610oWPoOEfBErkBG8fm4jIkg6MM/aOdHQcTkFIoVlI1a58DV5wVg2CTIhAge
hotKqOf5VwW5ikr+RerJ1lCzPBv+BmDxKo+pyy3k+Hb8+UVvCjVqSu/wMgrT/FSt
oCp24A1uZcNetteiUpwJnqLg40NlxpkKrjswaiLFQaN8fxv8IGhJpRfu0YhWMIFB
c1CW9WAM2PCFcb2qe55jRZEv4Wc+WO+mInKlVYVCDnfgKbUtTtaLP8IeBV1sEFTC
srspz47R3uzw4Bi2r9cJeE+0foavH9DlS6WR9Kb/OmLHtEtW6gnpSMPIgNL3EE/z
6jts3hgy4tIQ042ozKO/nXuUM7/G7fIWQRNKTd5ITfQ9qWcgQFrurzaCD07GkltK
RveV43DdTlH9hQ0f3NMuSrDycVjSISfPdur3Gk6ooZ5duM05wg9OdCI6LVmZ1aji
XwXs+kUDpXozT80U87BLJaeyUXJymqmmROL1lVhjqbyZl4hMMMFzeKizTxZxitfc
rUAt7UD0l6Q0SmqFoAgHFN5b+euZbwtds4LOZ14Ulbc7gF7N+aJS2ouiu7BVpDif
DRoYA1UdU9ReqXnQOTNLoW75aoXluDGCW4rn8m7H9jlbts+JqjcBeWzjZ8RknJrA
t3QQ7uhJg+WE87RvTqUJwI+m/ouXoeLANEDGzP9Y9J16gGFWESTBPbjnzTeMa+D3
jqibceys6dStT4MUWNDYKI1NzwI9veXnCjypcjL2L2rssXBcGPRYtHphEWQvUUet
H1yPZ0RyiuKQcdLLWxzzSPgE9PXJMUR23Ri/3sesKtchFk/c0JJu5Bv+VfnWZvbE
x7y8BKAAPTNwJaeAw7sO2fmeCA+/xfZkPoDcPhNAycgqTTG6ZqH528bnqdwHQDkC
xgvhLzYZ40vP24HhW2+JPFr+iksY3+aKUTQMSVmbDd+2FugqNDajTZTYWA8dQIpy
+g41PdpTGKmmfRiuRGt+S52otmtp3qghlOnLCNYFTfNA02V278ZeTxUDuoEiOMgj
cS5hGKhn5fwerel1GBkyjnC7Z1UBSsKBvZ/NgNWGJbXCsFQSRjGulInBtVZcTZBq
vBiM7KrF4Y9sel3cbKbLKYiDgUke/a7X1h3HNlytePZFJIsrMgyHikKSxSRds3sG
8P3h/cKrlz5VF+/PwEnVnDVKKSCrJTKCk7TGw9bWcSCf84J66yB+eT/beIEBxS63
q9VEzSOuK6fHUCVIe4Xyr8gVW99afCjZuJbCyR/2jX0enf0/NfT2Sah3sr55zfrh
Vu1shrrdLYZqgrW96yyJ5BPvkp5TtvyOR6IoFXvVI40EbRQjTTuIftvwf8ZjV48N
jyqRDyGhEb5j0EnYnc3xl1PqNiHZBr321CFyLOX9d/EB1uhDTnNb0B1yepOShHnc
+GSovose2S14nNe+j2RRwWstbi++y4Tnjm2KabRxbDU58vEur8OmqKb6/b/X6ona
uLWMIIFcV9OJFYnel17J7GQYGbV2f+V04eJH8TBiSb7TtTqqopgb3etP/pUU6S7C
wWYHRSxl9busd+ngGZI4qTsEKig3tuKkFDa9l9dGG5NZq170T3CkqGgwtqkxVirV
zcRsHZhDzDql1jaKW1Wyo5V5dMOqMBu4+PE1+hcX43L2itzdoxAw9g+8zitM1vot
cMRNDHMWdMC5uBuRckFA6uPYZqfzA0DFA9SuidyCM+2V5CbfLtVcexji56KHd1h4
YfkKhT3qiNfDTiWHNfEiFi5fx4e2qJmHGXlt+961tP7AtorrlgtP/oYyTA/uNQ6j
L3c5WRnOX6reJLZOhJhUhbvoWKAwyILIMsSEhD2adPexmuqSd4kkYjBrV985y/NO
YeA35M1Pwz1TYDref45TP4qTwl53SGTPwjA0ApCvNgU6ZOFjeF4ewfU8VQkmy0AA
fWkYzg4GxwjuQ+3FZe0M568/x3XhTsNeT+AOslSoZJLddkvX7/jqhezIZe6jtDGT
u5VZ5ynwRr9ZAldnmhB3dDv1F4JYkyP/IOfY3x9/yV8rGRGhgPtiZBrV7b2i6KqU
aB2Fn09jZzJOY3eEkixXGijlDy0+0DwL26eYWXj+xPixiOv2OXFRsViGFFJG5tZq
uZ49XyrZuLyHMHRzkHf4nWRdvn6jTaCJQFvzUA0GF9a+Z1JgyXqkzbD98cPd1kpn
ZmvT8T+zSaTdMzN8XACVfbZshAzUqI7/F/OkEswTiMY0sWWYLGcJCo7RsQSgYEDc
rdx8wpwQiMak04UzQJebdn+1CkZxY947kh1KEQrjyH3TQ9OgIqLxbULYLLzvODkx
PUi/6mN/RadWmAJU6HxEEhn8OY74RETUMY63SX+iD1h0YARfylvkmW6ZDhyj84xQ
1HGZU64LqHOJvLgSncCoc+w5FY/1QbKaciLkfFcq7cBqrJszPKct/tv/WAZHQNMO
3othyJWwNlT/+pv3Iw05NRmzGDZrzQ3+RTTT3WKCk1spkcU3WPQZ6/jZvGgWqUai
sonqvoHmsqo7pwyhxzirr+g8ufvJ8baloNCn0LywQzG+UC+puua9pQ100aAWBHgd
TCbk2aB88pdBQAuL110iR3vh7GZKizO2Xb8/OwSPoeMBKNRma4cE/TA3oTVSGkbi
a7Qt0/jCAqj62gpvDj3Cricn9inKPxO74uuzWYLHKBhf2AmQwNIy0z7/DIOv+khy
pWpxH+LR4xtQjj0YYb1KsOxQ1tUu3Pldm7W/D2NUoYy79fMK8ohouF8TdNsB/KTE
s6i9ntdKhCfIHexkdC5w09V+pd7+9f75nZwHDWTpWJMUgSCvBdv8wBymsnm2ywRt
FflfpMMCExsR058VtputL66R9nMogPbMCVCKQWq5BU5GRF9+G4vux5Hc2BrOqX1A
Pk9MGfudRezVmbt3unCJUUOoq84tW4/d2p825zaUUVN2oHVq77JUKBBDzoc0MKOd
S3+7Wh5kuB5BjgfCvxoQ8rt7H4zDxjsmtVShQ5jmCp/nZnyeGfwv2D+6vcFMW7iW
g+E0uuSRUUKRwMopZ22YniJaDGsAsMg0Gd9JC6a+nKP2MzznE0UvHz5GPh7pydkt
tYtFLl1rQqVDBaLkql0BFZzGK6aB7kHxLKCP/U2ZXlkcuv2XGGlyyDGwQW5uFQ/y
NdtB13WtzwO/L5ijq+7RoaRDAc6GHkklOqOGTVjQPn72sHObbgMA3reJMNf/VS9q
axhaGk4NiZ1C0OtkwriqbyaPSamHo6rhpeZCT478g/ZDmgzeI6VQszAqcZkyVadJ
sCQHj0eJA53BA6LTCbEsBuxjylDOb/agT/la4jYxkQQ2jtSWn0SqmLAaWDf5OzeE
lLIdzhlorRAgVYdGov2cPDJRXlZy+0ACMoFi/oU825hOEU6/KJzfTK6elH41F9Ek
+PRHCts859DyZmj9nqn7SoOSzipMQRl3wa2J72s1bMkniz4q0cHOicof/wLWG88p
znMUUUFDZ10qkAG+KQ3ZFWyjdKik7dHaPLsFwInAXOVVtZNBQmGk2kDLzwX9/CMb
/0yf0L5nkN4sEwHZr0+PFPTJL+hZ0liAxEkFRw11VQtlYmq3jmRoNnSJwdsYB6O5
eJDwPkcS4CvUXZ7Q1v8moK2297TWuhrJu3CoboWUIZfzdX1wG+Ri3mbLE0BBCK+3
i5lJGL9QRlOs1FMH39Ox5ODzJss7PUIM+mCoGnGNExPZl7br/JnC5BDvTHfxSQ1z
7Wvy8SCYXc/fZhIfm1SLPeHKO3ZFsjUe2FaiCuVcULHEhehd1oaHkjE/paT468B6
FU/z7aQO7E3BxHVxcp41JckW3iMyqddn6C5+4z0zAp0Fl1m9fRGvQbDEXlaTs+XG
2MR7VYFqZ7C6iUQ6rLZWpU6SO2HH2AisTIS7z+Ds8Y8FC5KYV7Uv0RcZla2xaizi
72i1qOP8VTxWJmaXP9KeVUVorlxfPmEirY3lRL+sIOC/iUymV8j3qW7S0EE1fGss
aRt10hwnSJ6M0X2TPPcvBU2U6ghbYbxv/sZkNakN1Q7B1c1LKM2i0s20xASLXpeb
ys7gSuC+KLiOXLNGhbpbWIlvJiDAqikEmUG1JLvi4woSQqWgMaykYrGzV6nSY1Ae
BWKatEX+2nyOaCa5WioSkqa5yygl65MwjYCoQAoZL0B/pnQj64TvH7Fm31vNPOek
QoSq2c2uCCREGFSWLd5h+OYsA7xKzxglriE+WqyS3dOYYhiwznNB7+r/Fek8Ve/r
/IT0Zxg82wMrRuB7j4AFTmhGIdRjlMczXtgbWCnVB/ZWlJP21g1sw2K8+M00zQ16
crXQBjKj0hVN2NB9WpXhLQA53Tiy7qRdztQl1euIRAN6qRGDfAqRVQxomsG0I5Bn
e1b3WhqAV5FEa7XpqeDQzJOlCpbhc9pum9kscTcKJh7kvvbS4DietL2jk2YYdzPQ
3nsZ0yMoD9LSHxJT/u9UbhZEYvYsDH+J09V2acbTHdys8CXBeqx9IjHAmrlCbFBK
00Afao5o3s6+FC2UU9WswYQZlR4cmniu45+94Ia6MeTu2q06Ono6Uf/tD7AJxEeQ
MxlouMjd5X3UAoNq5Gv3Qg9dduB8NJ5w4p/Xv85a6VOwB309qL288HVnytL77T1a
Ox8VbWlZfj1HW9Qx8WXL5yUxFHivtqykhhuvmdCF7lnhOTI35VIlXMro07KB8xfC
GKavqEY8XfiHneoDUVFejProh2qSy3VotJ+Vsit2T976QqtD9d2n2rKo10ubMd2E
6TMpSuFD1AxKtPPRU/rxudSHckWBuPIFh3zYdv7457YP+lWIIaBn6I9Uzuja6XHu
ODk2JlQoZyAxWW4Kq0tOiZGZG9UqUcO1zYLr71YyEhM4v7jXvvWiX1gvp1M0xa0Z
BGl/lq7aYP1lIcKO0wh3p28/Oti/C0+ofZTIzT7bc/9bd7eS2VSpoQiBp0YKNA1e
vSP1ZMVTZO26NqOBSx+yhrvTOCxAchXxXkfy138CVCC1W5tDe0uDWnYWCz68kcnh
2ZelHZpMGGPyJE71gDtn1Uq8fAUlx/7C0LecMwyC3cX8WSl6q9GLN6ft2/SWq+dR
SmfqMIjRT0kgosI3xlWMVIrlcKKyHvjs+PXb1KRzazhjznZlU0ict5YAwrHTVAkR
eba9DmhCd3QK6qD0x4vZRHQs0/Jho3ZMbbDIUzKGIt7BuPSVcP6G3DjDkqO5OME5
Abgi1A6WUZngQg0cbMc84JaCx8KgELwELW3Xkg186OlLcfD3mhWakJxX6ZaENObe
8zTWFcsagwjfyIgAn4gTtAH6hp2yxgg0S23eASb/dAKamiB8dMRNPxZhy5KRFRfl
k75G3XOpKa0f4L8CdOwWrgy7/HXkp4DjFZrjTHf78WiITa9jWXvpYyEyMQhpmCTH
DLaVsnmpBfPubBMJfmBbUKSVKQziz74rSzSVuF2iP/ekHYYyLZKZ0CM6Qt0DRCrp
VDSSH3kO4uqKgDG5hTwJ6t85gjMR3Cj9kZg4m5TQtRWJADMa/UH/UmgYrBspgMUF
Oj/wxjLQUehjGn3W1E/82azlpkIxxV8qgjHie0fUL461bwBs+q1sDFtnASolSK9i
kzqTrjVwOSQyonw5/MZtkzQGQgKNkhA2Xr9WzNfWjpe19dsn2zuSi2g4T6Zbco2j
WxlRe/LIaByj8D+hIHN4s8OGbo0xuXDrQ50srf8NUP9SC0168VuuyNvrUlew89i1
O4UFQgaA0bXAbELMGaW/RtNVNACsQoQHK3XHU4WarKk2GyBzfEczj78HJ+r6AJqG
zsTpP2EeXnAZKJlD8aRU/9GSJqOIUkcLxlKBWHgWsWqdk3ghO2ZsLudikdzTPLl6
brl8K8SzcODNTASP2x/SMoDcyA0vTI2uyPPfXHrqguo9c0iPJihzHmiP6zK1Fk7u
cHr094WL5tCwsG/oJSaShx666xB0NvFmF5ez90fIINKIKyUOSzERKFGx8Hf92JIU
FcSGzYvnN3AdcnGaxCnjWZ7t3tcRWpaj49hgDm1E4SH4Q8KpGz7gH9zHzWdTpX7w
CQ3wurrvDCCPDAdeXY0oIXEaNp7ZCSkSSXmJIjcuXpKDr8ojnyNvTsANkXID4xr5
8JJp7sT545+fseBWJOIeS5tN19jKQIsI/YAhoAqSh5E0uYxW9e9TMi32aVwOoQOX
AuIzskop2sDJs9SOehclY1rtNg/SpxiTPx22hRjzM3iyK2be7ucy4ZxJ6N+EOZyy
ySDQYgxcxab9ySboyGGjHtPchATHjmcjMCFmuMrfx214e2fotdqiPacP0jaN6RQ5
tS6xMtv3VhfBO+ROSVya1gx3JbcsJmW3pzhAWG52oI1z2mcEWS8PRXsi43wICZG0
0S20y+T3dpeK6U/UW/5vZX/ObO3vbhbtx7RL63UazhXsmO54Y+/7+Gwff8FnpJxV
pNeP+mghitVBcNpd8vdrP3EnPh+goVZr3re/JSGKvLdaLrOVm7uoQfHood4+FtyK
nqrj0SsitWxg2ncLY/+WYltaUJBPG6cPOTVSm7urbVhExstbvLPJs0OepWSLXi5K
Zw3bOlXJ4bYCqLkjd2QRzFuJGayPT4mLzSZZjLqXDk0H1TvWEskf5ZMU0z218hCK
p/BjFcWqP058olbrKW+KgqiZT5vdgqCbgYzdcyDcdsng3dnzqoO4VMg8dzRAlrJE
BzboulWDTt5coAXBY427dVU4xMEiIT3gkhcE6kBCsZ62KTXOwHMx8o5NRHm7S2t2
CaDBe3a5zypiqc+bYn65zOnVtbnm/XyixOG1ns/13bgry8qWrOVvVJAc/4HWp5QX
cSm0sr830/38QFMHL3v7/jgQjPgcxH6cXV+NKNmgxSa8lq5SGclx4vA7FaDpSBzD
mESC7tfNgk3iHO/r75JtH6qduBMbkxsGS1C+8PJEtyqNFdEF9Pg4J+3/kZmAphHO
Vgg5ahv1A2RVEAuLmjKIvOSmJlp02QlUol1D54JzI5WjuRJUne9WCxrc3n3kihsN
1F1ZUtkeHmgLJQlVgw9I6UObeU2E8hgJT+U3VVJwxbvEv6azoTjspL6QCUQQ2KeB
E2BDerE1zUUdkj1/xYcE9faHkgxAwnU1tWDf1lEBHEKSHwZSOxocI0Znm8CST1S1
TUglSf7wzMqyjIkm8S2q0+34L6bTQBClfBWeZ7/VYwcLX/7pgJaKfe9Bv5wR0Rn3
+NfrKNq6TWLM1PK3t5Oy+/5uxSxpWDX+MBf4w0UYpuItRiDFscok1a5YHMszfqJu
/eX/YCeaZxpmT9eVIrpd+kHhHdqTGtkTwmsFLe5BFOypsX5H4VNorWp5b/sKXv2T
ssJKn316pvak5m8pFfxenLM3S6i2bw5F0hJyy6GosNWX0g8JEpGE0MWQge/z7L74
mGA0irgTKcY9xbkMM4YrH66eJpNZQtRibsj/I4dQlntZWF9VUrI8cAv5QBMp+9DS
jOQQJ7fbd+A4cDsYmIUjnEscgmxpq/HgapprfyZstQOAej4hGgILXGAlrYje96eV
iwmYZlk1QFw8L71CkZB4ZgiXXvI7hUOb0zggpmDJOWeM3jaIBbpk1a+dcWmhKsaX
OhzOkpa/cyNjhmxCcFQYDsfduoY7G49WZ24W5GfZFij1gAZKKzV8CytWjVZ3k/Lu
COmiay16L0mcbmGKwuV200j24reoT6TsCgAQdG5yp3NTsCFARqdG2yqiO60u04FK
DxAfDzvdZJaENx0uuvmsj6nKQfChCGgSHK+UfyJhfcqy1EJIu6J9+DA6Nn3ZKi8J
W0EbdphNfCYrww8m0PvIYeLRAVfZMCPDW7VAgBi29UynJhNi1Mzginun31mOKL6S
DS+Mum5IHy4qaAW8yNhHW9So8KGw/7ufjHBUSLQLbv46AjMqxtR6DBUcYQYMx27D
YBtTLo34azfc5nMKBm481/7OpNgWOR9oKRL6iM5e9C/AZjDlgRgM1dlgdOec3QUr
CuiPXrE5qVxVjHsKwWdc1iY3T8Q9gOpA89RtlALUPF3F5bRiaXNmz9HKOKSHQqUn
20lf2RQDkbBxfXm243XbtAdUZckZGb2+RrFsNwll9mN61KZ8uE6eL2ldEZBy0s/j
ejLKpnhCNXNKSBLtQR2Mb5t4LdtEazPAD5/Mi+YelC1TEgy+qP//9SDyJRvkSx2y
B/IgyHh7FrA9AxKivQcBXR+3kuk95JWqASYaHEhj3MKor05JUQDoXnK3bL3EOWk9
QmgzyvUtv1UJ2soej4Vsj0QgZ+xLPNqbNAPinbQ4Wro+Va+wJ6tWtsiojDGPtfsm
GyBNvCQLrHpYi9A4294WVKe58Tz/gsv1F/d46R0PE3EP3+PHHuZjeCFu4dcZEmGt
xrs6h5YEmT9ArM0oRhYtsGgQafTRJ4dOS3iNBtlRU7iwr4OJ/NjfAPjOBaL4klcw
+G2ntHWE/pUvdFFDQiiu6jAJTGvD1cWIONwRE/rUb33Fn1UcMM2wXqH1IExKs2Gv
X3e4SrmvcvnfVHgceGwu1eLxFQ5noWdIePpiV/BEgX+3Op6T1YY/03MZpM/Wmyut
1cylwEuuwsgWrHkkR1yf34VLI2rvXNHtRKzGCQlIaBy+lTKQbhEc23TUHckKGT0Q
xH8jgf44tFoxHrTxLqjuXKagSv6CLz1IYLC3h4BanInuOABZwunfo8fLIUL8K4g+
j9fSJDLgbDafcb83A9vwcR8677TqRlbh7sc7+1KXY/nq26Jty2cd5oZLFrycsN+D
FZz6TE0hJy/8d0H4jPvGBJnbUDOQyi99RkTvM8Egg0mlxafSuXt5GydhKynUoi9V
9u6n24o3FcW3PaQ14AF9X/boEOq60PXCN3RMRtvUVytrU0zpkBzJ06/TIk27ASQK
zUGV5scx3NnUXSt1EmooppkLFetsIA61W+fDYaKaauUq7su6Hlu9r/c5ksSFkeJT
7dCwTH/jx8mNCUKX/W7EjdvOsaWhjvv/0eoKL/yTMji5SSFWbqGHslKOrIjmnUsf
onK/3Dq7/pTPBZYEVcHMlNkOoilJoOVgxQmtgh/v14AI7hkh7irwk47KwY8Ot5uN
BYTNmlGOTXydD7/gCeMgs7VVCptWhyjSxQeCbbGsjm+kD7wfNesdOBNiiu7CmtRE
NTm1U2LkbF0Bi6N2qSGC6s4VJ+1A2mjX4pDF3rAOvXEMJE/CaxOuA+XVhiISV5ap
5Bw+fFwuK3FidXJXHkVKM1gitjW8EDU3Vzght0pZL0lB5DesGNVvuJAb7wYDRXMu
i/+ZXOOIEvR5D3jDJpF24K4TTNFAs06wHKWp3VeNyOYpZ8Lt1+/y6e3roT4Jg7i3
pcS5RVZRttoxIS0rq9WI9zb9zENFto2JK1fbU4gX2+KaIU55ofiTrIR9ZKW4q31C
iHbb9K+1mWoQ0IACVliILS1fxSIvOYF+iHNohL30odlf7nev6YGrWQItwCt1UKET
Gjd65xBM5MXiLhz+gQ/ij1BUbdHT5gU26772icuz2LLIcd9aA3v+wH1wka4f9urI
BUdXY0TTXfipetKeaFrkdaF+IvmvYf0cZUjn5U2MScFoGtEyzp1o9sI2shekXWRl
AXa67l+DvrvwTRggZi86ugipR2lVwBztzvnzVR+TgiY4UKy0MhGt+8YlruY05PcX
g9CpBqQd4KIkynft957VMuY3MMpaaZ5h4Ww/+5HXFB2IoWjanYwxz1fF5Ps3SkbA
gM86SramtZ4bqjWG4xI2tSWdGcU5Yi46lI3io9d4s7FMpyXLIjHG4TGFCDfudv2T
rSgLW3734je6YknHIN1Z8RNSIDxxmmghhwqgdxEmpGctJO38Neo/9wiIjoqVUZs5
M6UD92K80C2JHBzC6bCpyDhAvr2oD/n+KF74JrnJaBNYvN9IllrhGdRfrBfQbBNt
Et71p8norI6NKE3GUXZPjja79Ca6DgBUo3FxXJjdMTQIUU9mKJ4A9M6CuAotRz9c
0Cow1Gy9obpe6JglccIvIoOkvQdidevr+ysMvsg4yAEOE9SIhAwEbbxVy5Zq9PDE
anE2Xf/i689/y2YDN1fpGZ0uAsKTDaOjd5UJzgA+zDJoqe1UgR+mElaqlW0J4qme
43mIa4HHTm5wSddt7azyM5iAw4005bXWNlSyqh/KlgHOPteMBc98QNcgRWB17PSs
jlNi+XQFMmQ5WpnB6Pb6Cslc78TKjRk25T/AiupEx5hdnGT9Qt6DgLa8BGAWB23T
G8uxUVS6Vg3RLjUoXGURM7OHAR+u1TuK36rjCI6gU5YOd90LsOZPxvQf2x6fUpct
fV7fHLWh+Nv37IEoknbV8DMWNnFok5QcfXJPx/yfxWmbMGjgDUXNnH00Bkvp6jb1
JAf1XUSGeeTeFk1Y8UYyCC/IRXNs7xF542TxFJnlsiIOwZdcqsTn04H08kBHIV1W
UXm9XHNudXIo22yTEcuB7Hx+MLUNucjnMKjtvIQcOTKUaj4ESuAb5Iz6FepnbCi4
+a2Xqb7uM9ZHEd+SzgR2QzTBVZP2YpZ5MDLB8VpQa2QqfZh4V9On5hL53XNB4JZn
Gar2CcH+tky/JpkpfdsHxP322qnhz8+7dzNT1yPuNT2+yli0sXdvk+ryTMDKDQQS
CM4Ou+lRST/8o4Cax5+jtaCqYFqfuKc3FSevXYPEBv9lk/b4SkOgvkx8ZMEU9ot8
yqMS1F89LecWotqJJaT3u2O2hyXYZpCDl8NFtThnkTMJtur4LTFJdxeQ+yV5l88J
oL1K1UcTOpdoHEa0saM4a4skPeP1awz8cRym3sg053WJk7yJY6VLdyYy3BfSiIQl
MQfPypVI/jNzdLyyQ2i2tLXBKvtTR1BYdiiKyK/A9AwNV93pcwAyA8WfmGFs188t
YLX0HfeDZevBMCc7E1121rEZBOwrh1oECPoSz/PUQV9kQcN1I7x8ocCdCj7Gc1Cr
ZgjyWOqunNYWMVRHLuKTnICSUFzrOgwCWNN7dr2xl6WBb6maL9j88DVat9b7ktKP
XqFRbrrM8xzETSizXdIeRnzx3pRqgnoBVfWzEnY5oLbbdfgAZpseElYT9OSaZ+3o
7ZCoCLNhpEk0AyBIRD7iMl8YbK6SnPl3EaNz5SoB1pb7+ghn/TMfN38zew3f8Qgq
7g4w+DEY0xQe1L/0BzvthcxXf2pJrCDdxfk/7RrgD2SlkaHCM0k1k1cyLtZ6eOgb
nN3t0fY9VYyfLNiCvgSkrwY40RIwQzDIQTAeDUtkbuJfbQ+Q5F/qOTpEckCI909w
wk2XWcgFCxFUtUXHdU+maXSThh1uWqsSKc4a/PX9MG7GCqI+RnnFmfT38B6/G/hl
Gi0lR7bz2uzi9hdVN42i8GCYbRSggWlqYMHqA1sjM9pignchlVDeI4BWw5GBdddR
FGMGw9101DHPcez8ua89cxQ5OARndut2DcSPw7D/e1qha07t7RtFvb6m49h5thnO
mnXrxj1cNBucLHCkzXg7SVNnTWXtxhqHZiL/zH77CfWiziDlMCgfB05mZeJ3oppX
hiSyjVUdHMs2gnde+KCQPuu+rhSZx4KY5tOgJdpGikeZ6WN7b/rzJWCWilxBA8hH
1WaCiJWI05o3DH0yojAP+4FAmGXY0th0vdQaGAxBCh/J7/ICW1a7/6OT9QGsPNTZ
mz5Ggr/BhA7sFLw1JIIHPoHMwMN5l0NyNxRMQR0fXc4HeR8m3X87LlUn+MyHFYls
ZAqYCFHzp4Mwu3RV54I4D6RUUiCHjFPAJF6t0Xfp9HlrNmGHIMS/AALW+xpM5Pud
igxRj7HDKOantQ3oYV/HC+HirEBs5uTCXPMEEIs0YCxRGgbBBcT5CP2Of+gXeRZm
4Sy030qOaqtspzq7VZpZKxLZxmEdVf7+hDLVmsfnQoCPQqUSdul92xMty8W6aPQi
v12gtZrRnafwtJ3F0GVeijY3m3HcaCK26sXoCspiXPBdy3n+EK3r0bEFD3/xSvMz
OM3ZJnxVH6MReCY70dUu9Upl0SUduYIRtvMzgdkkeSpuf6dwjhJYtOz+6cFR/M14
qbj5UiDVRdH2SybEnVONs8wDCLrAJgXjd+a+A5hLPleF6sxrj4/7UIbV4VoawqT5
7Ic6J9x32y4kL4bdhiO2BTn4TqaID4funoa4VmZAt8fVdRpdwRHhz3CP8hJIjWBq
HXYzK/w1cwIHnyxydzGn0M/VEdCZbYB/21kfnPpLuJakjX5IGVmMHUu9+ePNPaB0
py1xOd2y3CjKSaueAP3bgFFjFLp9wVPijWnRFxIuSgjxTrNE3jR+4yeRHHoxBYOT
8JtUW49l4j5VpK3MLgrXAQlYAOL6IgjYnZMB++LbIxL4r7gc1mqCyDt7N4jYpLQf
HzT5ZGtRjFHdyLdGYKSTJsR0JsUBGXtoQA7Rt6oNHbsAKd1UnUKVQH+H+h5szCrA
S8bqyvElzJ8mS0XplilyyFkR/nkG7wvNvVu5tDlezHnDxxYEHd2X9sh42xEs+UIM
wncCoOOH74Ck4uYmQ0B+o0TqV3S0hA30B4cAgDlKqomIfFyXehiDvaZ24sKfZXgh
BAMKlY1c/cv0h5VCukZNfK4w3dxXWIJ6S29ATTwv1ucQ/Bclrj/EePHWyy0jeo8S
`protect end_protected