`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3328 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
dnVBOIGMhMFpJZXzCENQ2I2z6L3Y7M6PBrtwF6NajXrsM+ncjGukHJa+TncOy5vc
lnmDNS5icGz9NiyxZRPbjIyirZ/IIk8FrnEJkqB4ISalWx3nFUZ7ke3w1mQvdlvC
fOfDiHV6/Sue18ol5KbsjQsXH8uN6ftCk6mAYYTVwa/msaatc76Sjl6ASuX/TuI7
9a4rjOlc6OyGVekbm5ffcyFRBjN8rlmyDJcIdlLJuarbOnZqD9Tze3UrMoUUffpd
W7OqFEAhMMX+I9D/aIbHa3GmvNxeiewWPwDqPgzp5ZwT2lSEL+yJzd/oGmIoglNS
Ww0EnbQ0KgtTxB2NWEnAozq3oaCxGQ+XA/GTuyfOXVId2Bhu7AzevEUEMm1o80Ia
smqkKhWtSmG+WFfduoexwe+/D+GRIqUsKKWSuAxF4MiFrsIEoI/GH8AMXGyf1UrU
MipVdXUvHbAvIL2np4a8MD5vwpPV89pny7N5onrj2uEPRPZt/+BpD0C/UodStRjG
LKlvxpGyvOHWq8QA0Ds4IAQ1gHRNXX8EkFWefqZh5RvNb3TNScfiqjBahnISLSV+
1mMWoiqDijQuZ6QFRgcEiv63WDAMbqGg6/ZhyJTn4Etf0ex/zk9ToPW+LqiIU3vm
NcrjlV4c1euBPnEOHPeFo9lKno1kTjn13pIwU/V+7BAd/4W+SQ1Kn+QA7/pL4CiT
l8858QQseZbGXGombehHxyDqAhWccSHwbsiZoGGBs26vLYCOUrLk6I8iM2kf9Wyw
0y3eH2NPeZkFvQVdESpLUq9ieEpGbpFdRgzx8ATVHagj5JLI3H8TZsO2zuAEUiMu
4NGe8xHjkP8vrKhfIaY5LbYmnVTJs31YBAltmhqET9WvXBKWkam2IArY3oYilPOT
RBU4L7XJBZXIkbwU2Je0JI6YZbh1Biuv6HlX75MTaXeKu2htw8SAzpSX73ImTy+m
P29X/gNLRR3e8rCUu5yN9LbnGkGxXS8o9pqn4rPsDVL9AQLlRl7A8zG6A43P5e26
wxTSDGCO7kq+xdz7Eu7wI+OOFb9XqvybPGlap6EvcamKPQVPGiKR1TrBzZme49g9
DjX0KuyRiibu6rHC09LviZ1fZEya+tHeDQ0dEZtoWCOwloaaCQvKbR9L/CXLm4A+
3KAXiJwNnAXLgBXpJD3BrILGjBd2jGYsdQAEb82DBCbaOgWaZX76UHxowLz18p12
sL0kfNrG9sxI9Be+1katOJ8MLSLGGBlxyhcXuf2F4N93SCIFhCr2WVnJnuDpCvFO
EBuedwzoMD030ujg9lI0BzuZP5aFk/AviO6T6NkBGhK34NnpphALmu11k74jZE5t
P6ohyIQEK7rmeEsIx28XshvR6SOGQauVD5v8AYJaTIIcNs6peSWgKiLknNbeOt9Z
g+nDa88GJhHHXibPlf7zqW6T5MeAeNQdkzr7v5DHzwXzzCiy1fmtwX1QKdyyjwg5
H5I8s3i3k83skL762qhtzgMlzj9saFDoXvPtTLLKuU8HBjP4rR2EaHOBAHZt6hOR
6BYNs6Owh4HTbk8MGnA6BRZEMNathGJEpEdWUcFyb66fjk9zdbI9UyE2PglYl6CR
4Npe2RTh1yio51AVQeIlDoOvgHST6B5uLQvacStSG1ILmYgqal/HO7Mzm318cZAr
EqbZ0PSPj8Q4c0MTTNcvs+JbQw9oG5BWR6FteuFojNRvCpavJpyP2qrI1j2WVxgL
OtSS9AboRGbUpydmz93dWKTOoFKXPb/PkaT+aGkcoEV98dosLR1AXyrsZlaSGRIh
Cnd6z8kWd1RsscKKaCH+LYnaR3ciZDYwHfRqeX5ccvB5DCrhRgGFux5yr/JRcixJ
7Mm8qxp4+AA3h1kO0hAwDvH48JXqB2hIEjRDCu1eOMlfDOpRTCzQBeYRPOVBTcnV
aQLFw/Y8AfgW4iX2lHk32x640E72KR+2L87shO/POB2/QFiIy9zCEeI+47XE043c
aJ9eNmxQpJpOw9riM9OHhSwOFQYdhGa9l6HMFCQ27FZEqexys9qNtAsxDWyKPxmx
ZS9HImEFRI1cXNh2xeDyOUplha8eMjHk61BcinTvA0Ryw3Av3QM5QWaQpf+N06uL
rw3Hh04xzAiajzbgClACHXY+nawrdAJ2vdfiNiYpTvCfV5oRph4kjQpJ51WySWY0
Rye+QTKheb1r9TghVH6O0naXUJ8G5SdtNoVDBXpzqQ4UBj5g2TBdMwBQXmwjOl2e
jJFI/ymleG++mGCJ0Duhs1Snghrw+O2uJMxuCQ4GVHLZBrx6goUmW4qJFbC1RlGB
1o5ThpjwzBMMtjyc88kT5O6TcWXp9/nnkmPR32xxmDEF14IaVmkbwBLqM8uf9QN3
GdSFM8G3aSRwSxt4aDNqKZGD9cXwAe8cAZkdFrdQBFhHPRGKAo+8a6az2orPMrHB
BVTp65r/xgAUE8hQKydY40BdQSFRVci32DC9oZdZJBPs3tWQtR7ID486NUxtxOIg
9KRF84WHXdBqadOPrT0cKxx8ooypXXYsUt4htJtPZZQIweTFXkth/y6iX5I0zWAj
ZSJA+pQsqiCdWLqACnWROJzy90JfStyPCl7Jr59c0aj7YTOSGkXRixIeEE4SwqcF
jMDA7VwXpU2izeGcNISSn9GwuEbRVNtUoJ3grNFWmQMannzMPosUsnXg5F68bjBL
kuxpuc7gxU2pV8EYBFrR+wYC+oCx0UhuuKwX1jGk2GwVf9bKIvqRYXDORpucrWcB
A5qJ53x9J2JebpfbNrZWaXkxRve9+oyADNRoVZcb6B+mRl62xZ8T2uj9FRtvbL5x
pyUw7IwfvwsUb62zoiH387ixhMRxswGD2c4FohZz9nMz7K/lFLAzMOirsDPP32tx
KtAhx9YiVFu5fPdlxgaZ7Nsy57CeZSy3CCWcn4ynTVVU+TGp0FMpGTRC/V4kggYN
pPTRlcq9wKguWa2BvD4DDpjMdtZYxWMI3gRUcwo2tHj+Sdc11m+CVO73/z8Oh2vv
oXdo3zHNCfbw8yKAOHvqXvVgScEvwQg/w1ShUzgqOq8rcgfyjLmCXbMfrlkxFSvr
HE5BKDZ4ciF07DTXZG/4mDpzSPfsM3UrCZixlC+C6z5oKVw35LVbJ1ZgCego84N+
MX05Z6AslawtgB4t3WFhNuCbbsVCy0p+GbFY9jNeBRVazoIYfC93NOBmGkHlzQXc
iU51eWMQGMnexdIvTc6E91KiXYHZZAouJNwjhvUhuqFExcmeA7xcYBeYWeHp84O4
zkXaxeFtb+h3Xje0q3p/eJGkvssuWU4PLB8YvYXIq0A4RXKubHvBmgCUv9NiaPWG
e5O1s6EzhgQRANGTeM8fl3fuB2Cud2OPtXlZXfP3ClqyiGUj9vzaCClbqkeYbIqK
Vilyn51W+5uHPKQquntQ4tH3pwX3S+9Wz5W9n4XpmLyKqcj5okP0fSM8S8CENYI6
OBF6yx7+OvA8ibM3oJ/uVOCqNcWIub2l306bgTjJVec6aFTgphG5geqCQ9BwcT0B
tP6ttKBhMOReXP79WuraKvaHB1lnc25A3Jjgy6az0uQLLwEVEgDpv+M3/Y/HFVd9
fyQBVsTIWb+A7RMthToBmIfdD27ZtAnDvh5uXYvLu6x7VwcaYO2+ZNQSDRK50Rfx
4sPBKEK1jATtm2Ck5KdD2CcBd/mpmqKOFYGzdXuFcKYsp2Z2BWWMTP5RnvG5aQHx
d1KxcCqwO2+sH3TPGQZMQA2Ph2Ut2qjI/wlGkdBjqHC4nipxpXOOtINYvdJl72Xj
MLNaTlgsIZUvpXNqN8lrekkVWHr21OrxCfsBIZ1A2mZM8wmwok2sdlr51wflSjyr
Cvt/p9Pz6YbPlM+1WQ+2Bl36BKCCFxG5E5n/sVoLk3IGNukjT8iXTXtwVUUgdmLb
LwraOf/feLgbFo1dXMtaD6Y45VBHS6OHTYw29Rw6pqpWbDVP8l8lpipmlp6k3JhI
PWWCAEIn709st9xYnHwr0NdD369EywYp6ZW6RPYPKYfuv7/Km3Ct0Jl0/El0iH50
Wqm+2VHYygRerynJUm6dSb8Bp7Dq6ucC0JdvFKW1Z+AxgPTJjqk90BjwyGxq634z
QkFFOikcx26k3+67PUUWAtZJTMI5/4XB18sO10egfbW9EBsGS15PYCyX1NDKeaJd
vSOvPVzBvP17gkOr5y7S0bq4/6n2kINvtFkK0mJgHw3gThOP48dn36BmbVQa42dC
fYVdieh5Jhkgty4utYr7Z/gkQNqLZe/5XQd69z0ozIpKkeI5o4jzy2G3RyyJhJp4
mCDy3IRQKj470ZOiWlgndA==
`protect end_protected