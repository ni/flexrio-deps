`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
hVdJHWSfELCmA4ds+csnOQAALbB3ps7EiTSHEDd//nts1r+JQrRE4d3bDPRJpiX2
Sl8d+xAK9BIi4i+3ruAzYvB6kuD7r+gs02Jsvd/1kn7JYK4xBxCjtdDFjVHOTEl1
sSh1oNiYUwLuwR1yKfP+xBhqxD2Dv6pCKhH1NdGilpJQ6cvivGkSunAu0tzP76T0
4x1pB179E7uIeRplfHWX03KzEBF+eVtfgXVp2W1BGjfAe43y1pCvNYZOh1+TY62g
EgAFgbo7pAujZxZy/YSiZjUr2mGp7o83qMXyusx8+rQ41D3X6rxfuP0RiId2pOpC
6oq5Dfkx04a1dk4s8w8cVg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="Sm9DkM+kBxuxXCFA+l3fFkxuSWV4xqRc4Nn7Ji3ukao="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
m2emGBqRy4AuduN4dffN8194qYvc9UXRqiQc56IrQYMiIVQPyh59I8SYabcDdspI
7AFHnvKD5YaF6tQfxWm+mlcmMEk2Y//aUjxeiGGs+RkKgbHitJF/K7nqg1dmKvDg
a/GaBCq4Bqh0EehlN4ntP5HxM4qcvSfh5m/Coe3drc4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uG91daMWA1mGkhgP3oZKMYye3UAomMWgG80HuuXg2E0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 57664 )
`protect data_block
c9NqBF2D1wSep1rW7utzHsk2j40aow1MnrccxUTvKej2Q1cyeDDbgAml4eTSXI8z
QYgCADtWi7S8BeChdv4B2VxKcS7CMq/DaQrOy1MKTfQzfAlK0iubmlTkljLy0Rwd
P94hdwjXt2a7F8/H2L+sTkyVpnYc3Qv+cSa+LUGzcOjkvvWQby9TvDPjpQeB+VK/
H72bN5ZBKyRfqSTKmENaSBMQF7d5IhOIbAqFKa6DLO/IUET9U2HeN4/tnPzMEvPF
i18+0CYV84PiIP0zZQvjw9EfPmTC4JCnIFF/b4MLwQQ2mnOagmiuLPGJhsAy4eos
VRdc20ocDQOalhAMvVpHiYeE2ZWxmL7E7MGTeFKFsgc8dV19foaSw4r62skzF/P8
mH1Mmb44cnIvtdU4pxsh9uYldSHnOPXq9MOZxBeS/UdKSPEi9UbxD8iq7+4+f19x
/QYIzYO/c1gCBgZ2isF++9lYBZ+VaP9ZDiwzS3d4oz2NJPB89cMnztPza1PUUeED
fvEIOzmkqLtcXyUWSK6trI62METvF56Q1fMuHlWcJoJW66iRAbACAtbo3tZkupim
tM+3q05jlU2uNRcdT1/kvdKsV+YRGqZyowp/zGHaUEl2nOSYMcjx3/LAPW2d943E
T3nRjKaScA+zNfk4RXWsocl1GkcHJ2i/6PEAlQDuw0Kdj8WXxXz+U1NCnQC32Waa
2ik1OJlfccBv/ldWdJ/hR9Gv0WQa1F3aplxpYZ0wYbaN7wF+Sed1lHnvxUwXyAZA
4Vw/n1e0gpxJQZYZ2kkS8qfmtZyT+zB6LpZ1tlNx9BODelnVm8ZrF9SMh99DB3ht
KEa8d3K+nhT0ZtGDUheGGKZ2BYM2nuF55RPryY2/ALGCcFwowBf72AhNPwWbP1q0
XiHJENPHp8rmuZ+BTZYK8nFjsZRwNH7ALr4+MoxL4PZRyE7emQarNp/V70MjYSRO
5utCMy4ImgBdWafXI1wrQD25IEd7hreyEwCAVETfuq1pb1NNahNzIyBQ+BxZqoY1
VyszZvMJE/gc2bl3mUt4tyB9qXuD61YIuJcYSN+nsrBCwGoXZnvF/oemBmbD+Xcz
DArvXXIo0txP3vWIzVC+LXDhjNP4St/VSUHXgZNf/RW4QM5DdV7r4eErmbskxUO9
6nm/F1By6Mun14Echvsf5Gs0HRDWSrFf+yqQnU/mu5l4cwpfJg8aLI29YsxKjnG2
j8obbWhAR4AzGOy/7UQgjqFPLjZEnqHa02ylltnRU/UTNGPDkNYei1+/ZSpnom7x
PzdLXaGXCYo451Iwh8w6m1l1aWcLPBDOxftRykDOWIqe+tRZZpdKdYmbicU6GFjx
5PrIrk7bcNgtFqo7hr2u0TOPGnHqwS1OH1Xa1DkUfxXI5UcuB8F6jEqGZBdGaMdg
s1i2Vg/AB7TL79eTcS3pAZ4cx9/uTux9xlFhlnhJKTVT+u5V3IEIqQaBIUNYUlzY
myt2wMKyRDdEm6t8imHN0y3RENaPS3hqV2bugL/9jxZY4Mjna0GSD/yMzChqdwlM
Qfe3ZI3s7Jfh7fy60TlL38Lqb4O4wmnzI9u5iBxpx+m5dzpeY3izLGUcl+3lhUjd
Fm33DTRVFUgBaq3kvnEn442H3DQl9HI4xpneFZbHlMoL0uBvZOXt5G2hEGZyXh1i
qJHBLVSqs4mtVfqGkdstbufrZ5iTVKEYIg8XpThXAu62hgJbKe+8UaqQVxVGtwfO
JeuSwPa7pjlKt+vKGyovADy4g0cPSEi55ev2wKSXw0xSt9iCeHgdSO80IrYrVEFQ
mnfFa4WPRS0gCndRvR0UwrFU8+KVx+SCtpI9yu76pbtiLdpY/X3IPGpeyKd4icR+
5HHePCi/e4VsI89jSqUG1MDT+zSoiyze6SS/Vtc0e6YVgK7mIyBj0LdkIgzm4qVm
4DNr4TiEHVPICw2XqYbCPNKMcZWXrw5TbwJkKoX1ynV8YBT0W1pEyHdOhkonzkrA
42zSzEDO2OJ7uKbk9k32mrgc9bkR1K363oHI+fk9SBSqepiRZ8FIe1zm1ci1WtKX
jW1XNu1kzqtipw8AAGj247FDwCRoRK7z/TPRvolozfLR0+NyX0Wykae+8YtK7gnX
b7PhOfpil0rwBjjYASJOK4hzPlzXR2kJhSg6s3eZwcaz2dKdhrKUUcsQ0qW7kXru
0Vsc7RFt070qA1E2fLN+tbi3UlC+BJy0+WueRz1pcgyh66AVgI6ZrgLDBpw71xod
syqvzCmwnu3HLBmv7g2ASkM5oUE1rbyOu1nFJ3AFiMQN03uUYhqtB5aBVuLZI8M6
a7vJhHuYv6T1bGEd/HB3t0yb8O8lCZVUa43tR6nrDqgV/jl8+vdbH2IzkcDEqu8J
kcUOke36gQigxF0hvlDhx5YwPGNKiXniclrM+uFjHnteJQOopEcix+TXVUY+CrVn
ig5z6haParJGrHjl+7yzFASZbEh35LsXBSFPfzh59W9Ujo3417sr/51hoqyCLHjz
xLu4rakmbQoPVUqAB+8IUdtuApYjmg7Dat6Gm+Y+sIX9x2uBjL6s6J3KV3icG/fk
n5jfLCpFvT+RSb3l1rZ6EXk2E3OTRCo1QCE9NIH7aqAzZddXJXuO1Nt88z/kSm5L
jpNuGM0xM7OIK9hwFl5YsrhFeBY6Ci9lw/AqTS04VGk3El/tTuwT6MXIHj9R0h+Q
4JNFIc95PnJN7oWqN94iYgklYGj7ZsrXOdBW2XHrdWWVvha5DoEXpfVotJp6gfyS
eYh//3hpAwlvSgDF2/9T3TQUsRDP6A9+RXcnKoj+BZfpspZCyGWlQOmWMGnyHuA9
qIPBPq+vmv4luXdgj7rDm5LPG3b5wozXh5LlzQvMTqYIQ2tKBjB6+UUkWzmQJ7n8
/OVDdiuwO3pZIqd+t2LwEQd0B1CqL/c2aPfGNtCp6M1Il3jti3ME1/g8BwZItb31
W0W0tdG8A7c1r9hlJfdzinYK+jRbaXnfX2kuc0xoPHafsCj9XyT0A2sLafc6TtQv
nwutEdSgcqOCFPjBrStzRC69nqO14VeDlJrPb96sitaCabftL/ovY1pU2EABzEBh
UU6CXCyIVbsv2ApKkpUKBcReo392Ey1rfn/C8m51oTic2I55ztKJKyX8IR5mTNzU
JjsJzLUa08SUUqMoolQ+ZHWDWfKC9UEEr1YpmhDeAQDlzZHtRa777Cf05d3qTJSQ
hkgsHc9k/yOhSkVkAMPcawgskbbxnFLx4VDkd9QozrK/aeDaAeEl6tEyThuimcpt
1WjniSesqVmYxxqE43LhLKt2Swnc7XPct9pM4IIRhpOxVsXSOvDGZu1qEN3lkxnN
hAfP87glNmCUUQA5l2xHgL905xdLTa+3PrH57B8dOiGWpUJIuNlLKOCEYb5zoJ6O
v6FSm8/mGomoTai01RiBMoJtiZnUfgFIBJgizCdR+5fATT6mwpGMSJT5eJYrFTHX
lgi6/27fgC/6bDlLktXjQwB7lUpFNTL4DHz0NkE76QO6hK/cPn+rgitPUxWVM04C
2wVVNeYo1zNLawNDF8mFgd2x8D8GRiF97iA9GuQ2MoAAyXiluHhvflnIg40IvlAn
AcI4Ohmu3WuxZmZEp/Vmq0eukxqgXCvgaWiEao3wnuu+csmFsXZCjzkGCQlQHFV6
XVeLUmBFwz1/8tUFenaP3/D57KqODhsYKeMBRz4jGacSYzu28hV9QNCPyHiBxrMO
UdHF1gqm7dQg6z7nRwGr9bzpLvoRr0Z2Tw8BLDvsMuTZ98vAdGSLBND1ezFfV0Ax
MHTtcDN7V8axJieSpHAlpFmDG7oeSkhXvHJ7jj3d4Ez2lva2iK6BDczLTGWwGxYg
rtYdY7mh4z2v6kYYdn/kARyI+Rn9i6QYmKXwMYuQ148VRnB/tvnwsQ5+Y9YRUSSz
rmsGCM4yStuAb4M4/dJx43HUPJOE/OfxOGlg3hSdj+AHCL/6T5aqa84iPNXKCJQY
OgIQv7kz+SuBh34wDpJBe7efiQ3IXIBOwkoyr6+2qtmnxMSDGH69LnEFLmn7kp5q
ZehEtkrJ4HYVUbMhcH5wldzOh71+4vGbex5Hd2xV/RTI4edoBKzAEzu8HKgyMZaV
dPq6LvFpabPmSznseApEPxW6cQYy1p1NzD6KIo86LH+HRDxt/6zltm0f5rbL3Kx0
16ssSQ/7AZ47Hvb5dPtb0H0+btSkcrBdORDqWjmNNbIpHEv8MGcS2BRAo75yD0wx
Z68d/8KhXoAfNmwDwUiUNrP1cIYJu02AMnhK0PmdRdGQzZeTW30ymzuIWTSBcJbD
m3VF9oFuC6FUd+slA+yQuV50Z7TmssNORA7U10EVRP4E8HLXD/DL+GBnInot079c
Vkv+irJVdNaioF6GQ1D/A4aP9RNrOC+rCIF2pdB5Dqr43T2PtOTczW1O0roUBUnp
pl5AC5jYccx4qMWizUKbWs2ucSRtMMgtTDShoO9D19+amcudX0vOItrHUABRXJmo
34EUbGxd7KcQlo0GSokr5NEcdkbEEg+B83PByB13PbJ89HWTzxJcHfKHZ9WYbF3q
nMUt2hU13V/jsbB4JdcrgmWmcVYZinyQK7C2cLEi3VAnEjnrrIchvxJJg0VyyYMH
qmzcJ0qxbwoqKGYmq/07OdrJEpEOj9jeoiFS5uPWuLRE7JHHjnDWHq9BUJfHrMVq
fi0nU0BaIxH+iMkEydW45GKo6oxi1MBy2N0f3R3Hb8CuYkmXLqY6KXKALldokk8W
Yb4pgzhdPQHZI4rvT54QAqI64jKLIuIFrRjViVCQSYN2xKSQxWqu3JAzdYtEloYp
ELWNOxZD9VyD/Mpn/veklnwVT7NSFlUHIVzvdA/QBvG6aPFkSsW2OK7qP0uevMar
dLFeOa2HZIfBu6y5tF9S2AOg4rzWkRUAh6hkhO6BEqXh2IdfH2NxanfQ+TXvSMkH
OSJbhwJtw9b0CBy1esTurtJiKsIPuw/WtPvlv1JBX1wXNgdg8lRlTVumaUfcLI7s
ba4T6kCt44keX44B6c7epuxFgvYW9BaC3Rs+TNQUX0j7mY5NswHlmuujI9jCxNra
WojdeoZJbia8VOuW5q0vBAcePIoZo5kjz4P28OdfyNS08WMBQXcErgRLfjXZDlls
/fv3akNe5scvzA6ENVuO7tLRTM3BhJCK+fyow8y2yGAceUv1S3P8pQHC5WkRU2Vm
rddZhuu54CN1IrXllf/avuIlzRig9FP2ZDa/IHRom7SPQjCycD9w+iHgR+YqZ/fL
cOzrLdsZ6vVIeUs/E35Ax2CqO/cQa4Rmf9gqvik0QVNPydtCb0tko4hZlUHrAQUZ
r02QkxXSg0XY9xiJwN1MOXTg1U86Z1U4iOzLpQK5Xzz2MqU7/wcdL+BLLAiDx676
CDY8ifFK6cOBrzXH/bcGgblkb93SHbYhQCf0GFLZkd48ggYVlwnYU95aKO485h7v
Nc4AnOToy6wj6PK6jdZzouNb327RfIFeko3L8+khUEr2YMxODdIiFlIwy+KIZ8cI
BplBpJzSNuoi9XJMyUvQJ/J7KYQNqp2aax9Nd4wdIgrRErW+RYgCw/U6AEcEYGBq
BRVGAcoIizjv8wQA2e4k8Ri51+QkiGCJ3bP5jj/rZ4pnyWvUR/roZ0B/es69mU8S
4eY5sggLbNJfMaOtOsArm2gXxnbH/uHTZMu+DO0s0YT8vXy95EfUCXwAIfk9o2WY
Hq7GkmGYBigsahRXr4DK2jzgoQVWgAIKyTmcd8215VhEeVQ39loEaALPyVRn+Ft7
U5ivOaTzXH1C2TNrVfUtKBxHlYGiat1Y/v2MCJEj1wOuDCQoNq0rEa0zlkegCUfg
8P4ge0JyQt94Uq7z3tc7JGrHhXJtgtJrWz+s0hrt+gJKpDsJP9ypgujDVTAkILd1
TSlY6UNMKRV8KIaCjVT3bp62ADlbhRS9UAxBoTA4DitoCLULTP+bjzhOr+m2VAx0
N6CPCxjz6r6Ulxw8AG0uR2r9omI5NqV8m66Z7Vv6QdzoihkVL9EX1TZ6lEc6xZ6F
DOQkoFSiX+FfgZ7CPUr4xi9OojaDltEo/ljbs5eBGJJw5gfWyepXKLKgaUAVKA5G
xYHUoCGubtEao8D4DCPLz3If4XctgW5hF+D2+utB7f0hmc7Grfnc+sjLjeXPFxQS
1h8ydIbkCVLRbZ6PVXPE/9p4sxPTgqZzsRorS23Up+B2df/8aKHgU0l42Mm7aqGq
CoWaG+WDtGVO9guSLpOlHKPbFk3+QGpUGlyWjx+8VaxriIq+gLjqBZi1RzHl/2yf
Q5I8C8//JkI45hLx+rehneUCYLVeso+4y4ynOj1goMLIxGU6micUirMpNtBl7SVr
9FflwYF0pdO0coEBfPgF11mG8gbCRVRWFOdpircMtPDaBeEipQDo3jGlCRumDukz
Rrsc49OXGLbmUSx0DHVnv8tCg6oTsNtQALTP5HaIG8W0OjJl8a5hFWtARX7zV2rj
tgj2/kvBzattVuA2ux78VCzfsuLZovv7Xw+4b21xfyhwx6uDs1HY2kt0BywbEjeQ
DmI6w3fBV5LgY+pAJWiQwwsfdyxO51kPe2R+J/VyrUh3nt3S/MZWdEIlxXfGZOwo
EYJFDB02ihaYzCgcOY0r47ZyIQsQzfSJlzftqs1HeMeSwgUn4fS4HpCCzZtrS7y+
5dFEnCefkPjdJJCCcqWxwFF6cVTlfdHYtLcurm7urMBIGKu3ZEg/FPmFaxLwLTex
/RT06nkvMKRdho1oU8AzTJijgatVoMaVxLzT0caH85649HQxx3zWxBuLliAtRVN2
g1pGbuj97ddmD3AYsiXAE3QOTareXXIbrfc+lkHyCcmchvY0KnnCR9wtVCi/Go31
7qMQdOwdJiIKSms2RCXhDXeP8fuY46hz/bXjZlU+3eyts/czui2hAd/UZ0vRUDxj
FxGz/IDhQh6rYZoTpGFe4tdu89AbaW/alYcHBkH9KtE6idFNRiTO6sLTE/wLAlvJ
GAK38MBSiacCeRXoMArFyAyURW8C5716lARc7Y5QJLOcip2lREg3ZpbfQEdEfCEO
24c+4y+o6ag4jvjFv7r17ePaU8mXoDvx5Ai6fkviQxNyLS5WApKyaADkZYBAecKM
SouwXrosX5VUcTrW3tui01kjm981W4Yyk7zPwLZimeDeZEhPxP1wiklclddjog/E
YYX1e+R96yi9waqBheTbwVq+dzK3WDHdCJpEAFju64mnGpSK+Sv4mkst6GkdyJfA
6mmbMcg4EqO6KliWaNRneqRLK6KrGtOZ1TNif6RW0Qi41hMS2w/qFMw+6vdIMrHO
aR4wU3YmTK54C7w4KTct6zJ+NahOdxxjlZRMCmwQc1zMPcT+euHP/Y5z6vVHNKl8
OhPNFwZF8dsW78jOYqmcFYApIzZ5gIf4PWtpJ8tqmtp0dhAzJBqoQSIlnnm0CdsF
LbFId131y9+oj6nk4R4M/l5Kj8Un1W0bYqNubf4gFp7tqmieuhL/OByN7neUDPcY
KTeo6LKjXe6bnEfuyvgPhAM49Q/RH+V/Mryp3SbbYynphSGnJG/uuKSqCcDDOzG0
FbNIlEX6f1BqIgOI2O1h5ceSSTxbG19BAlVXuiwTh2RxcROv04dcZZ7Kg0USN9E3
9Mr5NB3e+yCRjCiJ9wvA4fFT78/HfGJrU7FLZbU5uuu1/YSr/U7LxorYPG08YRc+
EAna++7Dp2GRpEmmrn2AD/ANmg2HZakShY3ZZkZMnLd8kiwCNhZ2czPMgsmjoKQ1
+EVNA36kbAnFKufsPKtikjsiGMDGnOvs0gNCIQJrtOH/kYTHFDgnWesXQ74XKo4v
A7qPEDjPGZkVe1cCzsSm0Kst5NWT+9KhbCHIoYswXSJO6aUUqGJJw1LC036T74jc
zpMEC79/DCH1KpW/lkDbEC2RYtc+pz+2Cx07ElwxNFalYeJqCZpusDUnm0QQSFiD
o3IyIO/xcWkOHH6xL0Dl7vz2KVGCfSOdROG6/UnWCtlwJJGGgPkBP/5glE49YVFn
/asMlubRnk/1ZFUyKQ5T28MR3qsHXrfSYp+sYcUEN99RUVx5Sz9UbSXAb/BimjPy
G2b7AyMmiJ6E2C0oKaVC8Lt25/eb+0n6RkyaKIaVVo/K+ljmdd+pcW2yn5BRDORv
ZWECCqd7zXB94ONgrats3e92DrcO/b16DqQgxyAooy5WNNc4hiQT9QU8fqe6gGlh
wBpRXch/3/Ac236LEOjqiFcY2ye4+iDBwngZVd6x0GDQzjHiNJMu5YgtnmQbbzVM
wk+9F8hktr0FrjNHPTHV5oKS/pLAAOvqiAJxeVrjrFyl340y2nX5iFoOcgluD8p4
RI8ySHRH0u7w05QoOqJ5ZnHsdxEGiEDBSQyJ89xu8fNTcHt8w223gxkbhuIFGxgG
AVM4lRT9PeahWT5dApjAMBBHrUiVuJdxM+rmImb4Dao5lm+D6b44vJvsZl9COHRM
rqPZiQKaI9cSbaJT2yVnovBxveLr8jwtgQZDCJA6CoOhnbtoAFtQVwTFU5YYDHPv
X5tFZdHPBu4guqfeHmN3QFa66Pbrg4DyX6xYmGu6sstTTddl6gj7ms6aAqy8Blql
WYqr9RbMYNN9xsoHbMqv1Lcppah7Y0oqpCCO1lZqYXDmnQx+FYf/gbYRHlvXPBwk
5rKUgbVQFoe3/mFGJowlAfRXpWichPuLIgOf4aHs9WcuZCy2SpijQ8EH2f048xaS
/pcy6XCJm+wEO7FubkazV9cBa7R4dKL92M3Zf1Vi0BqrCUDq1/YzZnXza7uo/a8J
l9esit/aIfxzufnPb++N4+kb2ZtLNSJ143w+pE2fzGiojAuq3A5EqjZGgKuzmE8y
Brr7s/EmWoquyGSth+xngR4UKX1yYhIJbeBPKfSSaBgPxUBaXltaSlRD/zYRQIHe
DaZOIzXWR+nTLnuKeKleCjBTzKjbTyoA0bu4gR6Z5epFcfx+pwG9Fcb6qkZjm9Z7
fZjkxgdUUFRBa6opQJyh4RlRr2ahUFXIhK9JVy8RSqrxr0e+ObFHe+tW/jtj0qvS
RQxex5bDSrXdFFudDjJFKbdIehNSEfJolkQjwPZHqRTW8XFBZUbhGBcDdtCXC14n
jmOlmG9PXZa+WZTd0RBc0czu9SXRorbQHer714xB8gYFQUzgQFHoG5IszQlQEgOa
TIu9lo9t3IGgENKpWTlM9YRvP0L1GJOXe9gB1ON57U6+SrDcl2i+azGOVdDfivgE
jpppI+HubnfJ56bAF8r1+8uYYL21h/ambWhnLf6qfjOSor5f2ol3clajCWdB6GQu
EnPetECK/eD1dzACid9KX8/s8VHkVQDDs6f49wqX9OOJSIWVyg3y4awfmsjFKebH
7v/Usayu8azY0iyY6iZHGDg6sqoct6y+5SZYPedB3SBMaaYtzYL1W2eiLW+SLz0l
eDRj71+o7nlbuw47+0IcS0vnvIuwsytZwr+TzzHXIxb9c9D7nymu5fPJKmc/yXio
15dYaO4cYJmWsvMaH1OBzP0smePBcapSxNNpjudlTrNLWayXSiPOzM4rgwnlDczr
zCLbTWuXj6sJnSXf3hXqZijXJknYpiGrpDI7BmkYGWtYd320Hf3Q6xcj87nPZKmg
2XLGiCPJgGWZ0iX67+v8KwWIlYqV/2aA4UJm36RI1CzMgYrj5cqHWcaHRQKEsDD4
IFMtCUVaX8es4IyHZtl9CfC7FCcF8EYR46XcpoxYzr8fvvdtFiXybXkQcw/X8ufI
Q8J/V///ApD/V/T0VJZuxGZQQidaLSzVsNz2ZO1nLviu3UxXtf2/x4jzr1ffW3kr
Cf9oqBuvhmyeNRRgmeYc6b0PPmFmpf//Mi7f+obmP7W+pUutkBDeN8veK713tG5a
jQmK8/NPfmyoKVLYoG5HnTKqgazSKfTvDdMAykJRtrM8OCx19Ghs7lMfq2fMok0V
oHgzGf/aE2zYNdjJFsgMB65unN58etnBzg8wIfl551ebpKbUIDdfKS5YZlIryl60
wcISR3oYHc7+mvnecTBhr8bKXXi7AJmr/XhuqQjxKD4NlI8BxcLcInhnZQKTaPoP
B0HEHAbnHC1Y4wo/QGpaFxRP8r0ojHgUSpgNi0mKSxqfzE2DdDihw8OTMudo+vqs
F2uG7ZlTvdKN0fLM3tvqBR0qy50Iz5v4fh/xNmXrb4YvVs7VvP+IVwV2FTcP8EM4
dHaidGjOVDKXUG1T2jTaw9nF4+xOHdeLrtoNcDnO3bpC9xN2oVGKs4k8tEREk7Cy
Sm3Hvlr3o66RPA4YjDFr2N4JJuWUwHHvc0zzzR6Gc6xm9EElzSmJEdIgO+cN6+H+
wpnKKBOq0puhK1wwRTjYdRmImCHg2qXYs0MZbmpwnN/hMCbl9eSGbRH0DTJ+eUBq
A7lGm5mUyWuWyb3lV/7USX06V/XLVsfdFGSPGzxqUOnjL/sd7XM7H8wgQ3IFP3hQ
Otm18ibHIvsMgBUUVCYKaqTkoLHzE8yETOR3W8fNRQ/+P38//qPx2mWREX9ilNOn
Zx6GWrQK5Uu3AJc0V/dGrHpliGchBFyxMOQWwEe5y5IV/PUNLC4IHMFhD4Lt74rI
uXt+OugNLux934zw4EvNGQj0o6gI1yM7qaR57MldQ+Yq6BFapzOgaqYH6kH/Y8Se
Ew4WOfCJ9+DQYrOEKgjlGBbXHKO4Z+O4di/XJeKPNe/g4ZSWHAOAZ4aHeDeeiuBf
URtsFGx6r9xv4Z/cg0OlvjD5J/7/u0RTt5DdrlBOsM/DdoyHTGeVhn3QI7qpPNfD
CJfD+RES0vA7/4F13UmYWes89viOSCQN6p0yOsHCuX8LNCBoLVGMov/IYHKM6JJK
jxBqBRTClWkPfbA53ExNVz7LHkwHma5AsfEB4je6JKrUYaySvA85ihR8KjS7CUBN
obcIAmHIw+zroarWPe55r0/FOHYoCzxk7afzSZZkv5SPnJdvY0yJAJ+Y0r3PMjSC
zugqzphmwwXGllhzhH3rveSM7Cn8bZGmKizhH2u747wo4B41OP4sYAe1VxuWk/zg
QA2ijTgupG1KHwzshYwkwYY7zNnF6/gbgdhvlVqRaTnc+lOVRLUyop4K4mXtdRJF
WBB83IyCqscQwdKk/pDr21b6Ix+ge5v5dbafv1Y9nC72fBIp/rThFvIEYwdpC+Vy
sPsDDHCfRquCRof7HbwIRUn3FQOivLPYTZJTezPyRhlYwk4g6SXTD3D2ECwadtOZ
wH6YwkdbyC+kSD1GRkjQSStsOb4A29ny3h9WOykjsFUtWqvt+EW9kamO7kmPT/4g
heCk8T1tTEYa2BX/PNkj9BK7U7EEZ9SrHV6s8MH731+TqjabHzDDGi4vjUnFk+nZ
jSxnbzV6h8bITtlZ5evvsroDKyUeZWHuOCUDReelSBpRDeYaa2r2eq06U4cqoyFs
35cVgU/wNA0rf/Uyq1JBXlaIP1WtoWXUHJ6t2nyPr1l2+5Z40K50X3X0zT5ClIL2
zLaML5WApKbREAmXGPvuWPGBJMdehF49WB1tFTb5BLULToRFs20XaNDRczekLeX7
w1XTRZC6CGWJD9kXoO+38WXoy/7TtYltW02hXXPDxlUOYAo4hLqmXLhYVzUdeWdv
hKVwZavwNNtpi9+ne3byLjIHGQLOabr2w5r3KMx+AMpgXtzzPCAvTBThQrsE1vpS
8mowjQf4ddrT3EKamB32UqMY+/41mJcpqfWD8NH5JJ/YYNJjkyVj/iHhoaLJkLjS
vQjVvXG3SVPtYMo5FMb/ciPYOptCA09AgIsZ9sowUnmVX/jvvTiMtabakqPtGO+z
+Q2m2mrXpl3Ebr0pJEFrtDhD4dTr2JgFvCU2WnbiiEzOy+CUVOsF+VTZGLWCdpSU
dlIDRMRTrdWcrEQckjErToHdMUHfphCAGCKEuhPINw7SPyBfKLSiGlRqKxwrHeKZ
0FN8NswEJQVWvhfbm5QZR/hh3su4Iv4vbkZ2J0IXGRnGM3X89ihctN7TYg0Kd9vx
GM02AhKLa9W6yNWKZN2sdEcSIUcjjR+hLYrYD15+cjAfYRab8qQazv2Z+UQt22Fy
609xpthh47q1sPRbTERYeomFP2rDrdxtuKdZNI5luUojpsc01BHIxNIMzDGXVj4A
FeXOmtBTcXKVB/0zi0yXqgv5F9f0xEeHcRO1HRcwJbud4NLy3EyKmy/HipNf+vwW
U2MY9qVBUMRSTpfFtfd8n7qEBy3CkJzLl7Xk9aSDIx3MtcTQwHCFKi7btxLkMXaP
ajx+C7MuZDnclbIPINeljrcnodTltLbQy0FnBipzNzagIliCXNUifG14xyuHUQpv
okMz9qqxBB54iguR0fZ0QWd2CVFQDsOSqrTQF5dGyjwOnocquoid5MzPRyEMp8NM
rcBULT9PXqDc30ssCZ1+cBHgzWd1X2wJbRlAUnWxO0TulaJjy7ek9p5heZ0oL4iQ
ssQd2EuLjQpZMIGNxhw4zUyXbbhnvi+wZfxM4D9zKP61wEftZGdlgIouYOz3JeMx
tErEH2yS5apiQ7ABLOlLXw1MlQilN9x2l3d3EsB7XJa1+x0EAtamjT7fgv+SwbsT
tjFJIi0L53FXXrJRGfvZMpl3hGr7Xgb7ZEGeEin6BQI4HPbJhqibTWOJnSD1Rik6
b40YK5pQ/TDVXVda2ongBzAMD8Ug6J7m7a3tiDsYVmol6/JyMGBR8wRAYWglbJDp
lvtVSyBx6ZdubCDu2ABQTz1XWSE28GaTFB6qZungal9QYpkVDKao1MV4uXO85E3T
4TvnRX695F46rWhMQlWpJ3WH4gEI4f+6opI2T7ahE7T9iiUg/R1hlRWUEv3xd/D5
KwWqaDrogL4jf7gHMiiYAY3P+er779XjP2e5ViCdG/m5UWbQyeW+7KuJIoHCQcAk
WEodnPsJ6mN5rfXz2Azu183AW8JMQzgextvGOkPaYvkF5I6hDQJ5Uu2Rag8ZArJ2
/EsbI1NBjYUniJ6495gfjyjxnRL8dq9rQ32ltx8atzVeAXC9wS7BVUprfZUfu2Bt
D2dYvdwpwk3knwFHS+QLUx6dlWSegqjGWyNF2aIpqrf5p7wPhLFIFdwYvQyLK2fO
+pL4/JJ6XhlOjQR6KdE01/9pEN+9Ic6VX8IZvpqcSlUjhpLbMGTEQkygmDJcKnZ+
/DvPxCtWGsIAL5N6LtdmP9nUJE2QNYbZhjDZXrDTn249aDL1C5uCix6FQf7rMA4A
UtlsQj4YenwbD9YRdB6PYOGIItCU0NCxiLAKy5x3GnCoIdh/868HqP2Sw/EZyvsW
oVqVEJUa+ZGkVFE57FipzEvA0C+KCl2Gc2w3ywo3kS1qbopBod5gohfXBoH+fTN3
liHCj0kXwrYsjwD2hkHK0o9c0EHLlTIXWGzvo0k3CtXWKueNaxB7bYT/dtxpXlOv
bvvOQzAsxBdoUY11TQHDZtTo9+wbVYNsZqlUhm0gKY5trj8txFbfev+15ChRKWLA
LDmyNPhuCu5/J9+qWJv+mDgAZ2T+MC0vzK8YBCsMuDxY/zB9WVCxQgdsyUGRkHLZ
6Qi+pYy360jOadGx7bRO6rCq78KnFuLrQCyjrVDHlzzHNCZPiJLpiH4Hb8Ou/cJY
CGWp8vI81UuD2P9ZPtzM9LkwCITNenA3UmBPSOVEFOXuyL5QNytiumhzK4MUN7UG
jpMDkKqOhRM4fNcNx/9DcrwnauVHrdUVQSITtG4+Rv4wR1tCE6xkG301G/UDN38T
MYtMYfq68vd4WX+Nft8Ghdo7Zk7WCTFS0wyIUOQhN8v/ayHaEnOInxm7H3dHFhN/
yabEONSBDKg4Wxgk8HMriNSgbSLNAR5rgAmROVtOxbM980TzB2gYhJzjQ3qMrfrU
iZuD+L5tmIYm3jfArac/HwhD5EFwOdyYrEykxqx+FS8HFXImUS+y16DV/CTUrfOt
aWiu7LaypqLB4SkzUMruI9BU5YLKWvkPqZrXn6ZAZd5ujfHVcWgcngYxAZGFhlRb
VTZ1+8XWZMpGe+zHwYkb4mqr0xyaCH85TVsd9ldnjxOiJ+yBrMIc0We/9QoqvFvU
tWzs2EtEt0R/ngZGc8NITeGbatVxmnfp6HsLa9g2r8Wsv71VfaGX6uVf7h2v3JFC
CofnrR/QvvzGZNsMCPr30b1iXoV1iBlCEsNLQnyYxfUkGWjNiRL73btQkPytmyMZ
ujd0QXEYse7h2gIt5VRUFtpZ9IASiw7nsCsP5RKKAQ1mc58XC2XKwrDk8FHtYA8b
o5Td/Eb3LfSpm2Q2cwmZY/hJYVgWABnJTmDxxqdk9SrppaomAbNNouxS/3PbmEH0
lRpRHPHop2H5QY1l261S+/tSfU+4bwmmqLJEH1cVTiB2NYWXHGScdKRkMXSAOKVW
8M4IBQJ8jzPRyETcjrBhON5B2NKa2A0XJodaU03pUVMa9BdBGbJ/F1AtBYbiQ5cq
lMtS5HYe0grnKlmTScwvVs+ow4flSITq8qpyHLEAg5MRxUzQF5VIT47ggcb5n11I
yEktQnfAYzjw3BaQ8n67+qUYwZ4vrJW9b5e+SWJW5YYnO4YFy9q165zLPenQzGlI
inQJ5VXbIJPdAdCSYn6436qd/1tYWvjfrOk8/gXe4troKav3JiJhb+c62iK/c3t7
opEXwdNZit4Z7n6mszKvTauOjreMZQbnh3R5bJ+KgS0qp/tDmpAtcN8+I/OdCB1H
LEqBDzuqWPWR8A39V0IAdg/R0HrDHhf/10pfccJCPd96WusUw25BUClLRdKiuN0k
NHEimsIvGrjfdXwx9bcHzIUvb1d6pwTNsbbusJIDUQiwe+i11Y2+6ECHgG+oTJzQ
zdlVLPOOBZxZVF6p2Kb74hbb388sx5uE1NiN92/GM+iYdodcO0W3K+w2sviLh4PN
9LQjRjqJ9sV+hI0XSRQiQAjBRMQxIWBXMuwtzYckacCYwTl8YC1vn4hkkohCWDjF
15PDF9aBejR8ucqSfCEG8v4N9SMc7B1r+UqDLxDmGvzhysEzCF7sHQRQH6Z7Cu4o
O9SinHqu3ubFdf4G4QeuRRutjRx4Zey1LL6WFyoRnlDWcE4Uf6g4M00Dp7IK0NUu
EWRp17Mpicpq27TH7gEZEHFH8r2pqIx2WTj7nRVisii0RdipKSHGKK7zI52DHjCf
+BDwooVtoGtFzDBD4kEw82sOJ7QVZLTSfcArzqnUgdD6Kk2b+3fizvitDdAoRx0C
f3AKKcUTlre58MScG9duC7dzKWdfU7XOjxt4bLkosEZbn1BvXprgeJxLY5ajMyU/
r5fFJEv5/TsQUqRD86re2gDBVwq858ZFTVXHeNtEUdY0t1nhq/WhGwKYi7mxrouQ
jY/O14H4tf2k0hBq8C2ig8cqguiUSLxFqDigygT8OZ8rKlLQcupUOWbWSkN5vrWQ
HH4aJATNwh9LExDylM6r2enW97NCweAhNykBcSQlfrOTGZQVH8bSPp9ntL92/qZ5
W6kNGfV0IoSh6Xp3gSBx/a7O2yIQASQiSufGjxT4KTDl28HR+fbus1WYnj6hUjXo
3u2n8xcb893ryKzIsErpfvEpKAp9GIXmyU4FDB0s+VGI8eLCNyOnVdN2HO56nFiy
cYpe8dp8M7gXCvGYc8nuH3VLxBqB0JIadrsOdXtB9b1p/C+YXNn6+W9On7pa9zyS
wqIzwWwKIMmUwRD5syidiq9LxYCR+w0fJtZSd3hQLxJhjqAUOZt7IgxLiSO3rgUf
ZxlX5Z3dPyjCa/4IYrQUemShoJRfbeAg99RU9I6vgJhcm0FvXktiW5oqZXLd5v0v
wu1R4aIXpLVzb69jITRAKQ3zSULgV/cAEX30ubjuIgcDYj5i1AMe2R+xISIVdV5L
E8gR1Ch4xui8lRotU/OfthraWZU/TSEpbkYdN9ChdTGx2hgohyM7Xf7VxjodtKmF
cvUmZc/SX8uclFKmiIGgPKxZSXJEykTmZq6ByGBHrNZLJ1zGUIGS+471Hsj6HlPq
pWjJoEvrh6vsGyBt1R881XTFNeq8BQ6Q37u2qL4SCksFUY8n/WsuluU3xOXJTPl0
BJwFXniYi/1BSxu502NqfKpj/VDSqNLuzPe89A1xe46UpjyR/+tk/owTperMftSZ
OYfZ/vrOXEce6bE3CcvonejoweFUycbkg1XoPtIw2i71nQUxxoy4fYbKoOsOgfNh
B0rH37GDZG1nUj1p896P881OPXmZIfw1vnbKrHMvHDhqPMpuMYPqKqspMuj3jFs2
SwjzrBtUw9SouLLWnINx1ABTwJsSp05rRAYPzEDdGJhFInccyVZLAQvMHDtc2C7h
O1uiUj9+7ZFMN2i1QvyNu53KNM3Z8LxVazSjflaN7ixWwykfcHuwq2NQvD2x+u9i
WqsqxI79f0sQYq8Gfkpjxymu7yhzcugT8WCOixofigrebnSBk3ZcG3WV7+1HdFtD
xepwCKeOOy/rR7Jw26LmbaVuPaAWDYFL0VkQynZRKE0laNk0QlfZ9ix8lkAx5UT4
o2cXUH96ywv51xbkv7szOKG/Z8yCPiORlkIv7DxaISno2h9Q4x16iS5tsR+NgMjZ
1G6UM0Ol/P7zK6ox7im7vFqiogyg9oeOW6f3/DmikrkhoyB6FgLwQMfgsioLpStl
trr1rWe96q3DRF4fg8WhLc4KWZiB/cMJqNafxV7gxCJizL2URtVTJlbZiczleK4I
thc+/hbsmu5yTqmot0xXsJp6FiV3Wvqy8mF8sQCeYelndQWmmWsxGlpxniRgUVa6
J0HC/4MHJ90dKHBH9eUPIQ4OJnBQ4t0LipKb9ucwEvvW2k7L6QXLJzBaEfd8g8ZY
88ASLLifZGHnjOWykgCWgGAKCaaS3fnDDC89qpPkroQWmUekFcgG3+woMzH3+RZF
VntAKrLPihbZRs262RBLTo9qyKMJxJIgBMkzceAlZj8PO13yEZ9G53ogQQ9kjHnb
OUAwlU05ZLD7c6fYpkf/3+C3ZjxqJhH+Ls4Ff61HQR7OeP8QGUsZM6nHZ41UVRQc
P+oR2VAV/ttXe8/MkKrKd9qfbDKHRu7v9h2rgvlOIx1eWdtD+36Eid0+9c9xxUco
xOKZkh7suiqfb+JJj7NANeuFLU/QMaqFgVfpIOHGRb3/+LKkB2d1zEg2FWo/3EAT
FDmZKIWG8aOdI9p4h7fDq+s3Y/NTCmTUgoNNBboR35pX7kBni4DrMAi7OjsGnFr7
k1YJ+uqH1+OabICOTz65GjnrCH5LsdFQrXFC4z71RvyOhhPPuv6MP6oe4GqvIOW4
RR83+p0HglUxu0G5Xx4164gmWIVFWNo7DB28/RSTzrHaIoTKnDyXreyABy2FKYYU
eVVrKxaWd7klzPxr/GMP6g048KmOpJmKZvn6SnIOnI+AaaA7owMdbSviFXNE/ou1
246E42e+zyaWzPfFUAAS/UCa2MS+84j5pZxy4ad7SNzFDL1LXouscMt05YW/dmg2
mNOGapj5jCR4MxYIe78YSY2MfnP1ydIu4RWJd9HTcyIDiVuKc92ng2APrqn+RoAp
PfhvbePvOYqDkGVnb5MYqeNQRXUywQkxIXle378RgTbrWsDz5AmZLDtGOgxRaDU4
+++zluAU8epcHp1xl+oPykhECLJ3j+xUqbHG3Mdih0lMEs6VoBwdOq2b8jM/Z17w
XB7/8i+EA0/Fd0LQhKfninzYvgA6v9TzL+6Yc05SpkZBvG1zBYw02fDmvkfBikXH
vw0eBDZePj68p3WytcVTZBBcvREYKcaoKxiM+Aht28xv5FdnU+4xdJqqHspops6k
NnejtY4ebh0aIW7xKhTKG40ZUaaAfONRiKFk1oQl/Ym9f5x/kKUKs8Qv1b+L60zL
5vDC7B9hTRBWbI9Cidgkzm2aXOt9lYBdGtSGSVBNfnFKUEukaJp1b5/OTW/nmqls
3uwnWKwHbB9uvtWJFKWl6OcapXaYjTtyWHUk8Ht13K8oUml43M2dQBJHMMv29VaG
Ji1epSrNbfRjzvQkyCNyN4hKpNTjGRfVZAy7r8DJONk7TIOEHH636nrwt9YGvu66
1vFixNprA9h9jyUO39YbkT3TEpuwmB3xUpXvoOBEWXrxWsxOo1+/fjCL5I3UG8vF
GvCtGtnwZIWSZtC5I7/Mp+gSvHEi0gUHgh48hg3eSkeVLc41fxNaVS7VKr+XL3hP
3Ikr+UqCunere8JLJI+rnviQllfuVBCZqOU0rh5JScXYT3Ptmx16q1DbPuhlLpAJ
dyEkRV5fMOti9t8gWwmnVynjhrKGzpaqCquzNGIhazuTUKjySdC6Kp0k3O1K3t/Z
K6eE0cgh0/+uSMMz0NEj5LKNHJ52Fm9gFU9PYbCZEB+wvrZ8QekxKjjlBVn3QSRC
bbJi5ILIPTXhRcK8oacAZqSAW6jHhmky+L4QlBdlXWMxw8PkkM06eJRAtMMObIv1
qErzrphzxrT2f16WwRQwZoVxQLzna59Iot1YJhklpKrCYhu3AbBwLabX+IyoVBaH
vXPHBCi8w+j9lhMcMdJi6uOI45tpMHW2xiNyC9pDWrNgx36MDJQBBwCOFNpfAd++
MEp/Vil+nt9YUeY7VTggJ2LcCBwv6sLxSprcs0hy2hSRI/apqB46QKAxeVIQiGZS
MB5I1Aagtqu4fREvO3BANM7p7vO/pxUkP7loxxydlyNtRxy2a27toBSaLUVuzkSW
KEPdxYGk3AnziNHfozNEtn4mYo+sYWK8EVFEkXAiBn9H5q2jpfr0kLxW/Gg4C20G
Fzzb3p3rHLImHl6L9wIyNmtqbZei05T2GTszuYmBbvBHJhZIXCenI049gS16RiCP
vo14WyJcOPqgbOxUd+M84Q6RP0ARks03S4MONqdWAhFhgnRR5EK4feIgTdhMywp3
8QNi+LEYe+cDjPtwe05B9IJgto+yFyBAgp1Ss3cYMHOsHfQ6Y2kGQ5o6k6m106FV
Qa6pE3uBJjOnW4SxpITIwiEuFtUI6RFK+M764KFd5m12gmLsTp8I4gsapgnFRfqU
SC3WG4mUnQ9W4w3y0rsEbZ6DBjy4PnuQoPPD7XNsUMd1AaQoNJGNIA3fJniG32FH
kYtXgtXFJhTfUdTEIoctk3RhyuumLmiQMvJDDKtpT4d7BRL/EfBjX+RtdhTleNPD
M2bmyuJMgVWtAEaGfGmd30szRCntzJRYmGZ2ai8wktHJowaGefxhymTY+IlXhZiF
gDiNNlBXnVoV7gmsZ6UAo3BTEkCNe+MK+KNS3A41bHhenzxJfVajGuEFClbnFEwN
WrJ29hDjBX0VYniSShsoPnqHxx6TWvB3Mqu1Z+m+M9ZkUpwuSJIUeD6dWdW8tF0M
TNZjV1eMaGewQSQDgA85ftRhqtiqREHSyJPN57A2PANBrB82B3X10+HrmrRp8wkf
9VIJ3Ufqj5BokadWgfNsY1MWLJDpJFHRbyyRY7jkB3FCJKKNEuZPLvU/e5MdsMho
PzwX76qob1GOVCcKOwiQSoPKk70D5dqB/Ok7y7ptlyjDuB4zyTo6fjUoOjzz4i8J
ZEMtHui0Ms2+ESiLqPkUYV8X7WCW/9DuOb79qSTtmY0P5zf9erwRObxo8uIHC8iT
dyXjn3R9GxnBnjhUY3nMAqFO30tshnmMXbWX2LaHXIM1/4J2MlLV/h0M4nKSvz3w
NsHuC12D6RgqT8twTZYWfLqPf0kIQteFF2ArHbb/ER0TtLncMbSzE2F6t5pJ9z5U
Wdo2ATUXVPSB5Zf40uug3va1Egtx769d6r2oA4x2l9/kDMZWNkmeVoCFMuUEbHwP
zriMabS1XNTt25xt0IX2x+3jTPX8aeydwo/sceECVytXlsyEuoU/GiDOCsqwix9l
6C0U0zT8DsVsFoc3+FIsPtkWA65HWnw29mJDaBW8duiatOxKr7VabZ7xRSLb/Tuv
WdRLHx7dGaA22mpAc6kPvYO8tU90nU6YkuaLN8m9hYpGRonDH7Zgj0cigekO4gup
cyEegVVbVpEs55RUz9sHnFa4qC/qnXo1gCQ6ZwYonkkdfVGdOFfW91tHiMsdWlGy
gUnB+3SnogjIDXjN3o0AVHkr6WW7uGp6Xcp8BywQKPSkNJHlqQQKSO4/ZtpLR6SR
/ty0SbuQauR3s2ZF/1dqgdCWkfcb+DM/lWIUno6ZgNYy9/5bGGtKxdSeEGF7+SIJ
hqu5/lHH2JF5WSKfcyu7EFvMgZxx+BmIV0/FiMpWQnQ0pr22qZW9QxCOTEs2xRPE
zRkWol+KMsM00X56L/CgnSuo4rSw/n2ifmRdoAUHPr4H9JBx32jfHxHKQ3KOTUiX
g3wrA/LuBh1oAefq7FBZuErFI+MaUh1aH4j8MWb/fU51Wob6JPCWAGO7lhOic5ms
tT8soQKhbn0IxnCcHykEUoRzC4gS6LbH48rk3kp8NIb501Px3A4mizLf4P86LKCt
SZPFINSrnUNohJ6fCBSgA2IQOG3sMZgCmGao4A4mR4KDW0/u3zlq3RTqmh8otNkt
/m15++Z5WMSu9DdTNaVNwc5yvKMNqHAHMLq7MWIp8CdUBiUV9yVJxjk+OYDdAOfL
94hjd3Q4/Xt0v6YZ7daq936RW0kJttmnTCQ2xdEyM0y4GkfGN+8rrSP5cE0JNPC1
EbFhCtHIdQ4+8rFNwfWI34hlXxz2aKXGlsukQMoGKsqu2VIS3jfGkCpxxYgWkTRx
xqdOCBq8ZTyk/7qKmQmsjq8U1xpjML/RC4wcACLqx9LTUWOMzTFw8eHWcvOHOCLd
DHSSxEBgDALftoi0JAEatwRqJzRDV1Qrg84gjXYOnEtejRAV66jRx2I/u2gfgxnZ
DwZU6AGZSjEqsRCSQONTk4zU3uGOJxlU0Jijr0vTzHShxPZ/ug75B/8QoHVc7I+3
iExIkpWDowW7WM5DU+/6b6FFny2TwlichvroX2IzwpC0xHzNV7Z9KKSdDCACrRES
a4D+f+IJa8FUOVoUAbhcJ0NmfFca0Vb0w2N4vDhzNZ4ALifnJ5de6Ob462qCnd+4
pTHn3YBVU+RtcPF5QC16gshIh5OK9YrsJKVjxfUJCaLCJXi35Bf5s9/tQ5nyDGuK
3xIgrbPUk27eP+HIvNXdqN0BUGNIYf8GaNOERnEwOf8zii/Vr0sOvn6lv/+vBs3L
liLiAz/N3kJO8CIfqggXRMk6fsfDb9TJWHWHTRcAxaVk6DYocd7Wqp+YcLzyUOUJ
YyplyjnwXafYQ5NFT0t0jBiyQtdGTQSJRIokTIr9v8S7d9CEQL9nODyI0Qj/K1Vv
BcSltj96wFvlcWafNHy+0kquzOr8+KUJ1E1y2oXh0kOywjYkpj1q1CrtjoUqVUFw
v6p5iFHO/PTOVLg0YDYykKxFvm66rw/6xgFpRO/MPHc684nwrmF1e9sZT5/FbLO9
ozc1kLbnQy6vwHQ2ajS0J3VoCQT/LgogJfczfP/QZ6JLjJnd4Ap30XQEAyRRbTo/
1TxV6ZBr8952VBghZtVdhwofM7AXTRhkinn7aGUJqpaQtiVgZxeArUL9InQIFn6N
FGa+f1d6/bS4XTSTmxwASoWpbBiqMkJ97TPtv/mgm3kWG/7u0Hc3nCJJPtxvPHNc
FQDVF7VaOFjlbJ0QD1W8ifQsu6LWke+g6Ky1s/xQ7GGigLNpaXOPP3lU3OwQFpvX
KQMFoMzWJ4rrtyvoF5NZnCgIkR3y2kd3WpcT2LP5Ec/7TpN2Ol74Srav+YuPBExK
0MMo1dm7KmgnYT3tqYBQhfhYWh8FcQ+8gtm//znQJRB3Ac6ZAMdkWsRpG0YgQBcV
GaAnjrY0ztRc8mpDnx2eImXDfz4B2BoXMspmXDRVXSf2ZQsrqgjVJptW+p9BLK4D
4zvItHTt3ENHhXdkxkAgSVV6zMX8MCE1ozqHLInpAgtwya3p+kpgmEJn+xCKiMbb
6VnmtsBL4B8ZrXB782kLeyUwVYRayffU+h22lzbUTfuGa99fEMP78IJ8zppi17Xs
32aStXifVWrcSBwiuUO2PyDYAyhYM/Jmj2+ZIhpFVqRe+y485rlB+Dqdf6dNzJKm
tvi9U2LWA5kwAsoE9QrWNFa7q+LM7frPA26viEoYWAu3P7kJcNJsnZUU9vNQq3vg
7Qp3fwXD3K01z0Gn1PRrnB76VLvdls+levtUEDt6oLszfNs6BOlb/9H54+GnF8FD
tmOxHdBs0hrtmDUdwt6/9e7uXlw3MKwtRjNzJrU96xHHpnJUUqjrpGEM5UYqbirT
wMiY+T2BDiYErVMcR59DBq0BXXxzCisoxUXyg6OXSLCvdgkBx7ytgdqfnFqEY/Fs
LGJEW+fVkFT198biFmVhv5WE1uK9lORCCf/TTg6tdMxRRKDmfHqyjLDZ0KjReJPE
5N84mhhu7Y8RF5MTmvMev563yiGQ4UyYRoeauIwtaAd9MBSNHlRW302hGcg4br8M
eA0nv67rtnb5WSLEZgGZ5zeeumYXr7WpWVEyx89kMp5saCK+w8Of9dim+lIYV0m6
cTaJi/HGPlhnUeKwFfvZyeM3j8aNH8UpBE588Vh3YACcm1un1amEzEUf/XvvQkRK
0H66v48eU2rn+WCqAMTOLy7Lc5JAZmT19RJ5Hvr62iDKyyKjQmdG3dmw5guI8cc6
b9Rg+AqIMHHbCD7xXxg81+4aJcZOwpnO2k4vbUzsz3wECTmWb3kvv5QvDQznS1/o
fp2ogfvGYnScUAdhSbh3B1lSyxUMVdtfqiBNUtf7v9yg6e+8c27Q9gZUKSqNd365
VTxRTiCVASrG3g+ebjtKmxBUN/dOZeQoXN/i+Z7xP3BDWrj66sBG+IGfDhGUHae7
j+GidoQEi+4ln8J08axlY53yjhd7NiQlFF9e5DvYpvMWQSPU8ty/C+JFntPvBK17
s+ky2nfj14cRyjMoqYpT9mqdx7GX5/2d92JIpWu7XLcJ+j19MfUr7/7vgABbHRF+
j1W2xISdN7UJco5nvc/neIiUGmcjEsT+oU2K7wPLCukKnngb5N0Z7rJxC52wKRRj
ESLmM9J8lWPYxzn7G9pIkWIQNzdFXwnQYIx/GTUZ+kCsUD0xTNZorDKX+pUE5dDI
MkD0M5iXykC1wn5yRApKB3eBpT3gPlmwFhUUFpdq/afc5WKvQMTuc2s83feOqnxF
XsD7AdfdmEl9Sa1U3eTAbPb6gl3eHPKDQ0TO/tWhczupskWImGmNI7TnTUPO6Guf
CcjGNDHsQOXJn7p41P34DZIwqv8q4C+3S8Ld88IQAGhc5vmgcDtKxVSskunV03o8
2bD3k9dcxlLXjRFtQBSeyvuR6OgBMuKg45jfydLR6Ewxm4wxmKzROm6VyxG0R1JC
hv1tJX7/isbkQtCMIo8AFGiHTKtZx5sUxU2CVkP9+FFy5W7Oc5mDSqP0K+yOFYiB
VD+MRV14dAJDnK93k8PdDwvSMhljHRliFC8NiTMCrAjO7dIEcuxAzXNoi4SlRjvp
wQi3WIR9h+ee0gBgvsc27eDtHffgh/W1XxNgdtdkgRrHJAuvbJxYCRnOp4t/QN33
BpWElihQlVmp1qvsg278AY0tVPjPzE1Bpf7yRHNgbtSYNUZ6MrR1oHVXFza26r23
orNDLi0zn+Cf8fSd8l7Ik+uAw8NBcOr8W401hvXS9qf5pMcrE+4ogag1PcebCibO
45QwMpbtHcTS12pCS4f6H0VNd6dTpHfVjVfrd0IKeIT41D1ec8g+Jq4m9fZWMW9W
P7GuEHdG+lIc8BBuSvLuYme9tw3GK6CwDFxn/YHO55mN16wvSFuLVGmgR70XVSUS
AUa93hegw6BAo1QsJUezn9u4gXbamQYRWpbvVSyyROx7SrKaiXIInXhkAEC+TJkS
jnacThDOZzNLfIKsa66p2d+29xrJuJbqtfnJgWIUWQfo+6NNqi/qgMvodJ56eueh
+70b0ZkbiGXVY0ypWd8HovNyyWlEvoxyazJMHCzmFvZiUQ2JU5GmWWLBoZAVVIBp
7g70NCaDrpGyfKQIQQI3yj7tzffk9mLzXy8lIb18yiX9ZAKoOhZSGaQUNRQZHcv1
ogsgya+QuAwT+eq1UZkM6BKrLqq6sMy6F0nqRYoiYbJNSPDnT7Mziya7uqHqaV1Q
tWSUyjBMZrcdcWMx0agO1yzqAqnzWT13nc71kR5vV4aOGoN5zYqw1XzXYXoVdnBv
t2exLiqRN+JR6UBfE5MeXCio0OMD06MS2AMJdPeMn7ECeg/mg9/FFIhFhJH/xU5c
MPblfSTI6XsFsgQn1Lpd+EV8w68wV3YfV0AOc+0fM0Iuv/aA4WtljKNlyTNNzcEe
pggS5J+982w/Kgg4KjMlikssoJzB0emLcw7u/6fIR4kbG59J9GF3+hwb6ArJxk5X
P/MpTKxyHvMXNjiSIe2q3uOBXfGvJStippLYDuewEqVC91sUQYgUXhdwLHJBKh5t
fsxbEgYvViAHmPjLlMS2w3a+PO3akEhW+wnu54AZkM7liZoiFwbfxAC08oBLcVaJ
7TJf7sMIrB8MEZLqaMImIitx1VCuVavBaoeOCBajX0vTv77QAqelCiSo0IBRxwc0
eYL8XYLVJ/G9JPmnbhPlT2KduJNbe6Cm02Tkzhh1IwXsrU6T0AErbCX98X/PDN17
7eZOzGDT8PLrDQsf8ctM7Dg4vD8q5jpms9B0LYTfWLv4Bm7V5ibH12lbY5CEEDT2
0WWjjV1xdAi/o/MmbfXwrAipG2RKhzK/LkYzNPmdAoky85VkwKBkbgX2MVDg51Jm
s69k/xxVxe7T61VdqRLj0DhPAV5unV1uylEh1dY7kmaiLVP9cQFMtPYbVrWFhuCk
wgy+NEJngVYUaBDdB/d/r097wKEP6+1yXIorajJ/Eke3RmSrx0H4BdZDNSGl27My
3ys26wDQaVLV3lxUvQdpBjP7w2TX//JkyXn/ACKtCdcZTwIVZ80hLipcrpGUjLcW
zoFuxNa5p5XHUbu6/QbuMS3fKoq3eX08f8I0waSYviIAqq4AT+5leYsjBziXo0EV
NGx5D4AX+4LgJfUB4thpp+GHyggSw3gb19OIqX0wCjRuTn13xumXzqoP9shV73yc
2shtUDtE/6JJiSTo70NhuOKUs3f9Tk5eLlZFmy5yd1DsJFJq6jwoBWgstEBvpHLy
wLBHhdbAkBCjrbDyYMHUyz4iKzhKv+UyotOF7bRkBfEjf2rXbkRp9jEM1MLbzSBJ
awjGL44UdWNZ5RRDDJTL385/ZsOWdbDx3aYs2y6KK4InVqro82PVXOh8zYrVxfUK
aJyzCk4DSkhLIMyPzHRYccWjsl3GAn3Y8PjaNGTQ3dRBtu2zWgRlKZaNjNJfo9Q8
5NV5M/v8UTeageutFA/NucbllS1mzUW8S5RRAo4bNNEXZCQ7vlZUQVzq/W3aFXaQ
rk9M7mwd1EbScuaRjmPIm/wqsBox9Gs+Rp3bUW3DrdNnnjdYAhh6O9xxsY1N8F6H
QQJqB3Qk++yCY5WiibZ9fvrYTO3JF12khdCVDLDgGyN8O07LCZAj0yZVaQEQ0RCq
MDSciMj9/zHRp6cKSob5s0+SA4hdIZAEHpWg747So/wdDSYDA220rAXKD6IUQ4jO
AvwrCjq4z5a8ealPxZZTx1+VVAd9+rxz8GZiyqqwLBU5HPCUArvWesccwOWVOkvI
U+8vf8OJ+IOHPX+QAJHJ6SJHa8KUMxVmVuwW+pQDdxjrp5QWyBLWLIbv6Pj77YDD
a0z4mDg+sbc+QAccruONyrHInGVH72M57cbbc2oAXr7Qr7PQBjSSTs8pYs9o4sjv
ZkFJCmpPpIx2SpjA3nWvmfMBORIIVdM7BvBEsENnxrMF04XZEKucxTZDbvHdaCJP
9NE3ECHfmOCs4wZ8thwgtlND1By6I6gGK0ughWLQVSP2gfsrKCNpgikzDvCE9zTy
PUS/Lqx1uxP5JxwcpmWiLU8YZUe0t06god5ycAsWgwbSBcYL7dWhQXToRqVdEfce
Fmn2ocpGyc8YktJwgRSOf756BzKENNw3cMpAWalT698hJ8SfxSFzMTb3pa08t5dX
ZI/Xr/k/FHHMVURkXdBok24FKKHJpu6ji611RZBYMFb7QGrmizbq2KUPfIgiseGP
F90L8ZXX3eTBYJMe0YzFx1C2Gv/7Z6ZNt5eikFvpfbJ635uK1mSwGgP3OzxjhcFX
5C4K96akAvVAE1wZw72e4B9o6YmnBSwsu+HmqphSTqnrHbtUFd8X3t3sacRNXJKM
8P1hQIFqh3zxa21KyYYmUQkVBQwlLqqNG3KePBsTWKtdPkOAWRLEqzOAjU1A3VZD
XXXdlHUscQmKm2ExcBypBnNpiEwEHthR1aQ8048qvA1GSStZ1lqnPEDF7C+tKbKb
2yJLd+mocO2oc2oQY97X9sZue/MPBISykBHDmT7r5QCECj3R09R36IuVIjLqpTxp
QQk5ct5E0+hciPhHS/pcILG15KtXVK5nkE2We/ZNe6ebmGLklrxMLYZp99FxJKVB
kQPOyAgZpIqFe8EA80fqk+cWmn9ys0AzuEMRsM3Yt9PDmltiq5lV5buwKJlobyce
45cuEmCzOmXjdwVeN+XRn1rRNZyAPw+lPcgv6H+2YM3liycEps6ObmVKBXd4o1Jb
mYnuq6lIYeJOUsWAX3pJ3BQDvB4QBZNg30iflqQ9n7s/imtqL6kXMCZHMmPFkCi3
yr3R9m//5cdBFUSfgJ1uKAYgi0UeFLeLIxF45MOcQiIKuJAYyXyIodVs5evQKLsC
kIxBdvKuinvr23PnlOoSdvXxE1hZdeImx0ayEXqsLWK7mP63k2ij0cfEypTEl388
/8WXyqDMPevoVkZW5UeaNOA/CdSPHF+vtERA46qmdrYn0+NcYl5gsIzETFGhQ+u7
AkYsqAQOHpStrAObMFu0jGaH8W/HzIVZWtI3Bm/Z/V4UxVPj5Py+zXr6utIIv8Jh
s0Ra/cpAva1oZ2AseCMKbbaK0jleKVJoUuzDCwu4E62dGbDb8xABIBC/r5pl7wbz
dL4J9N9bhNrGHk9Vs/5jNBYPDv58KUyyQ2+KiYLxHUrKO3eXH2TvRfq1N7BBetXb
/OrWdZZr39POE5IQGjoTmaAQxveF2LK+PvRQqTXJBAJu4mZOGEoRVut2lnZ9Tjc3
POGRSd08wUXZpEPGxnaB5yr+HuwEDGIyZub3VnB20pKgY8jtFdgXcNJaURlvAFoe
5amNZ0mPBEp/gCtjKg7Cgj4XSEZtK1o16vXSFeRldoRFEiX9UdWT/WtSIW7c7BWY
t8xToXz5OtT/OEI+1NOAwFq92Hy14VP2izzWwHtZixfwMB6naGP7aXuqRUImcde2
cYtoL1jDyJSphJubRZzQMHxWuPDRQoyvFsQgzJR0bHzzd2h1UWvsDqeKAVyA2TPx
zuS427D6qvJeXFuDoQttRMDr/QKwLGGwq+kQcEZYEqwYEIrFDY9iGaLOx1I+nhfa
o7uyDqipfp6VydQ5c2GqIgQhMY+JH7zEonu6eFUd61Grqf3eRPiV3FOsxsRUTKFo
P5nwCvHDKTLCGjwDvvoxfdINpZOCQ7UExLyEGK/6w8HkGZ0hAGEGuz3MPaHDMXCY
8nkQ8y4BAN6hrnW7YMGCJqqlmMLXGzXAKK4dqxpkIL52Opl/fkRse0uEks00ny5v
SY2BFCoaticqPmrn0wtNhrnfcucPl+q4+MP9Jc6Q8M6Fpq2AXH3963GUuaCnA4Xg
kuO2n26AekHk4Sb1iDbTr4dNeRnN4nMxMy+Ndp94DSkye/uyhQESka7LJUbz//3s
wo647GqTI8fjruEvUo5R5tOTIZXfEaGAlHEnMgTNMdIWBbiky2UIE6JrjQ5F532G
6CganjYoVEdlb9hiD2BwTD8cmAM7FP59hzW1LaoPrb52AFHviM8oPGmkGVRm0U9Z
OZadNPlhBC/3Lu5/6+C11gFXoHj6MqmSSYKqmPkE8srDNyuuE7yCZfG1Qey6BzeD
C/RKcDo+QD1qGKzDec36HvsmMbZq2wN03N0OMGa0iZ6RxbrLTriJS1iMJQsVGPiN
mQvjRAcxflIxTFP8/MUe3UmftHovXF2v68n/VltTcH0poA/ZYJMVwTeveJMT2YIi
pSzbldefVvZegbd0aBIa+IBYZdktOdKxiYE8ZMNeo9uCSn7IJ+EcGB1+gTP78cQ2
vJCrK4cjHcue/PS3zvUv9W6qu1d/YK0/qKLZAdj2ruprd8KPTnBA/05PbzWKDq3n
3rIM8hS4M4PLkifSnbH/swR6QlCnUw2RN37HsXkrmfKh+46DchzI2H5nG46Z/+bj
QFaRLPJ+GV/dgCWNiD57zFYbvBPBwrVMtPOEmizqsDk2tbQnm5f3vzOZx7W5MeLX
Xo37WKZ5L3Gq97qGlwptxZ4iIBasV6qutJb0BhXUfZA+3IxU4onxZrFY6m8pbE85
exZ0x5KAWzDVnPHpr48eJ6xgYZAl2CmdPUJjf5woOWRgdNlY+VEd/FBBP6ig56Ya
3bSxeaHGoywQxnMZR5Z7TCTVGYaW2NnKMnE44mB8tSDY+ZbchkOSFm75b+jm1djR
mCOsY8ewUnNyORYnXuZ8dleejlkWsWg3LlxZi7Nm4zZ29cVi2vx7SzjJ7pFvFaIF
BeLHY8lxWDUruNBVpd6cSzN/XAuoxLhpv2R0S/V4GciMQSQqm3YLoVNQ1u5+/jpV
gCbPbQRj4yC3wG03+Layw7MJPAbdQGGLQcZhIODuYm8P+L715QDoAn8XBc6w1t85
DCKHu/YIi8/rq3lLZ0sSfZAAZhENgSFlFo379Xsc1HfiGIH38NP+R0l+acv03k4M
Vagt5xTpZzScwFaqAA1etaWULGamsWP5DGruFYKGE56oPoLW/NbBZ76ox6+IuRXU
ZFefe+LWyQx1+mWZVREvJeE1CZ2U5ZRNS+fMFMLfyuCvkA4Nm6Zf2ppyTuHfsW6O
iIQZIcPrGjtnG8BQ8BJpIqMLfDmUuJmpMHoXPs2b0T06oXqnIN4sDtndj8eywHK0
1MZqQ/iefWXR4/7cKumxhaJLKh8x7+aGP5IFg/auu2ZG66EZ5UY1CeZPCZBARuvt
07/vW79fMcCnRpoLffUTaQauvmFuOFznIo0ubbhKF3ObhzMmQMuqt13BdRuQi5o8
nhK7pAPqKifYRvwoIy0WVct4vuKukezlT5tz5lIYPihwJDQrt1c7ia0aVGPVSqma
iA185o8IlSnd32ou/KERKP+oQ3l+hSUmQCozdA4IC1bVH95L6chpfaZiA0kcfecx
P5Ei9T46VmMvmoMI6A4DMAXs/kIPcfseeSrVllF/vySRX1LT/CJN1Hy5AecebiVk
ziYeSqYFNjt97Etj/X8Ek42ZGv/YH7iKE2zCKKPZWChCcBBaSfLaE8lIc75mtciL
g9pWv7odkRrlkZO/8y9aKdr/dAEpVeU2/v3KyivbkXN4Sdr+UrCLBnMDeLEbwnFT
mgeIT58WV1Ol4eICop0hrZPs1pIRGvCf90IpXzo6ogQXyUim7Z4J/ZRwe9gKvfkC
uToG4UkU8hL+m5xcUy9fCZoLbum4sFBrWgQKCirvlt3tXaBGOo16gGwzgcWRULWE
xB/8iAFEjcWl+bXRqWNuTxbb7OlTSTqjQSFVlHQ6Z5NEb5xnfmXCGJU71qFC4d2E
gzhRrOzfzmEH/VlJOzm58y2F7xfOe1pGrlItLhYPyijVfK2S2zfqvKHWJUBW29qO
6BPeIfTU/Go/YkG1gKpROg387pHDSYa3iDh1LoN98FXZRb2/RvYmen53rIvdYNYN
0WQRDwJrmKwUcqjZICyn+yD3vrsYSb/X1XJGg1gc2meB/G7cXkLx1/3RenXBnY7e
ROYTNGP3H7JwUBP2FsQiOzoA6psLq/UpHAJv1R1Aa2nifr87zfzJpva6b37CSlnV
E3h64In7EAeJQggvc0nHMM1lbEAgElNGcv/8GZOkv99q3rw1b4pAff6YrXy1H+Ha
/CdZ2/s1Zxvoq68+UYQiLIyCuecdpNcqa/jTrmA3SgCL2wQQraWtyMbuLNf5QfPq
5qWH6rgIb1NtMqv4zHfrtcRzagoC8lQxseNsaIjHAng4jqxw4wW/booZO0HhkLPc
L+14xVf0FursWfTpbH7VrfjVQK5rf41/7rlB+QOkPaTbB4Dy80aJeTX7uzkTvV5A
Ckacj8eNmAvULaVUxICFXrWuoUMTGdhVIytEpcDaZp1C0DOGNEwHKr5DVvMzD4vt
ZRLT8jg7fyaqKg1AjT7Rc5jU8d2SYyCc00/yp2uGYWCUGYy4bIwUMvIpdJ+qwmss
GVKR+zY884W0CbizrtlL9edKy3qFC4SQofC0ZdkcA7cwN3KSP2WG+t3huxIw+N/u
2rf7Ws9TdIpBMEjpbVG1HhiuThUeHFy4VIF/cq5Pccus8tOEht6dzIDSn2VC44KV
jSUrETQDjruOm0YefrqZJpJot5rsZ3LhhYgqInhifkxWV4sM+AgLbSeLZC0JdGYL
bWJB7YanaibfjuaMrIr0MgvCluZusCf0qT0DzHdgkLaqo7kLbDNCxFWfa+yjxFOn
aEUqzVSgD3nCt6Ux9nVldPxp4/xe2YznSSYC/NCdlKf3lo8rxej6sncEJW7Mhi3G
NJr7q+vqe/8jUBMaQD7zO+D+UaYIQVcs7Y6xNTN4o9LFMCgvUAu1uGO+BLEGrITT
L5P2xVg67hM0FV0yaL8URAdknU04FMCW/Tm66xzNmM09zitp+fJnto8e18FHqe42
U7atttzNbcQhhsT7dXLDXEEv0wMwpX6U6+ZprHGpt4HRqBVQa9HqNhm+Zg53NmIh
wliD9Y9/jqbG5hxACiNrLIZoWX7K38uUOyR959n+Cu8XZ7yaUk2+fMhshd2P8txk
p8Z71xtv1eSvubjzCmvsYlo9XDN4SklsKmO+p+Sq2LFn4VkGAjxiKP661p2pWTi6
Lc2kuee7321L2rtVHfxQdrXbl82zAocQKXDujcjvlfWXwnniQkIBhWd0p9jiTReR
ZjGfgv0QXZ0We64dkzNhs7+2rbiUtbMae/DrkeaLAcjrjSZ17lAftBZX7mWPBgeT
6aaqPDT5BF1sUqFv5B5r3TsnYFB3QMFQBt+eXaHjkCE5wh4mFaSUxTI0bRb0qIfR
tv9M4VdwWsTe2GSmifR3f5JIfy1aTnLw14A2hu3r/AXRaGRkROB4fkP2l13OgB4p
P+Pzu6kd5jzaxg0qsNg2hglx7J6irzeomKdNI1CZ2t7x2r7R9fkPamjYy6KqGg/z
LsKpBZaQ1irvV7TdYA39ODtxh5vgupQa1uHvoOCkkGLf4zpuIAkudYbY/Ouqi/de
wMTDbZKQ2DoTjwtQf7ZT1HP1Zo88cTlcgiK/qj90D1mnGe9nYEPHfhmMjfS+Ekok
lrXaWdb2XzXRz18OwzAHfKkjXXmXGsVOLWQ2Mm54t5oEglQyZngVqZ37F2pC5+vE
eB0QVgOk6boHCZ3s5OQ7MiZjGNBDuDF9z83PcixvI/2GKAOJQiZjbHUHabRncx6Z
8xDZCeb+Yr0kcreYoCUVm1pzQOsbp6EHylwAzHi9mBD2puFIqwPti2kgKtlXEP/u
jkmoG5ylV7ygT8XxdzD6ApoT+3AlvR2EPfQTtI5Pj7WH/uteg1+uoD9XCZV75elC
miT83oNK0qhho8+LbuNZM3X6wwjUgupYFIwhLabduoj14tS29+CmOJPeR50ouncH
BeNMnYATyy7PJWQs/WoJkIQoMsOSUbFp1YtdHU9Las8x+HJopsagPXyqjyqQ5NI7
DxnCtJLbRn6iS9fSvPlW+LrRJKhCls1/FK+Oj2PRd12oNKgnK3gzGXlycVcAIU+m
WB2wo2hiRSPcUyzGpVxNxjoAq6qxV6SefobIiaYkKk3MMnklgO+ojaq4CftgXTPK
7999B/Dicmw0h5KJAVHBGIRL09X4buBh95LGnuW9qYJilp5L4T7jjdyJWoeESeR2
AE9qKYn/BTWyhfz5U25LMa8TQCMQmm4elG5COLpR4nw0FdcnI5UAX2wuoCngf6M0
IV5fIgRQygZ+3wDilJL3WMcqFAoZEwh8O9r9a+Qyy7iuAOZjDfYw3ctRpkfuGpNa
Vz6XOsGXBCwS9eGLVI+iyljmB59+Rzsa5B/Y/4uywUD+xv04PRNuiO+4mtH+LUf0
FrwZCLR4+y14KaBFNPr/LH7QZS37d61Pu7x2JWIKdyGC3KGfKQU7sGOc5oupfgC2
A+N77b9FCqJqfEaj375YFkEuif4CW+1gqV0bjSKrFA8Tptia9faY7Xu3srp0f/Cf
ol/Lz6M+MLeO1amPoDNiCaNFjDaSp907FqDKukG7+sci1hOzO8SfEwiucSQJv9cl
UiQrTwwCTxRYPogh2BOzBMfVkiYtU2U4QVEKtpe1UnuP8vjeSse5pVl7y0EX7b5h
2e7UF2Gvo4C3dLik2y4FR0BNpxQ/6HjiYRxjpifEJGqqn85Vyf0tJO7NmKGMYijJ
aJzQRqeqttM6RFpB3VzMYOxVkBuAXVNbka2Zie8RPi9PXi3F4oCYUenH8W5J8OW6
ZrPhwjvieK1OK/vfCPuL8LVAv8QnnpF/VrzV2X5ufAdUJjNXPK+zWStegLSnO05X
KrErLJKVNjBn9Tw350yTI+ZwDmFcpuQIw5EtPFSmZXU3Hvv6zwGvBunaGt9Kzpb2
j/U+hdK2Rw0n8lEe6KbvJEh+e/9gzeHxNmloQ/Bh3YiW4LQM9FnZIEKy7L0yD0Pn
Pnf2mQ9ofFS+3KxA9bkf6N/fMTD4ejFlfnm+UVbuy2R0wMtwhe6TxH+6Pxa0SEy4
zg46ZubFx29Q0+5hQL0O89amExEn9PFLdnQ0bWPRiAL4FvCX14G6PdaKXS4XcC8a
SZ5hW9MJh4OLaHXDZSv1qzTAO9273im5JPyN2u5Rj1DC0w/G2NmivZ3a/Ycq2tbm
Xx/KD2T9zf7690GUghZ63p0tFRH2wNm0BzuqgburplcgnSWQEftgnpqLZyXiMWF+
/vy5k6LiBwFl+oQjIdQDTSDDi4lZ2Kiz8c8o/zSi4F/Rg1FOY3F8GcODiyr81/Gi
STAow7bxTK6FIZ1yafh2YZcpUYh7ZUZkMddEUw5+GmMox44sQrwyvbkgPVZSfeSh
+a3tmQdvoyyx6vqMVDWNQ02CnGMOEKtNgqAxJlbaZXZMlohr/Sn1CsKsuEUP8oBU
y6ZMtM/RjhaFzgyuj3YzVXOzbU2kTSIO0z+vbelCkhgK33obqOgXvZ7/YXRaHpJy
5W6FqLLvgB/U6C6Hakk68U9hUOa2vDE2lj4aMXLBKtjyIccQEYcbLw2LDNOXId4G
xbH4Wd4F/PbaHnuBcB1eILus+Bzmx6yoWVkIuQ9MweyNkluLHegSWbndai8SNrPP
ohqMsVOimy1UrSssyITxy+kd0aYPkI8397DNakY5pJNDARpJmqNkocRuuMZuAcjA
X227jpNIXbZyVLNj52y/bwSPT8eUGJci5KCsO0fDuyPktbVjsbRgrFJlqXt/pdc/
yhLBwkHdYXPI85E8eYhXiFxkG1fcEIGpjsT/qTn2XNJESI/RZIuzgwc0I8UJs2xD
97dzVa2ZDIQSZUHg8nL/fFp27gRcGhFLFDSSvuDqf1unrr+PBu+DKi0lzsmGh/az
vjdbVsK88aAF40uLNF+kdJEkVgW3b1JF5OW7sOZhcJtC9H6/pTDw4ZSTCvA5ii3S
hqprUd9zkfpNoM804XkP4EdQpLzsTIquh4cZ7vNfoN1/UFZxxCd+Jh9rw156zlqI
zSusXdXrAVUAjtVJKyMzDYq4hCkwRzzM99gipAqovkICs4GKsSR+Oz5Ff9QDCFaA
WS046CRjDSLVEgEsCfxtUoy42FNa+oLMdOPhEIa3YUX4TZHV+vOIFgKs8G32cfHi
6Az8jtVozAGonSIru/zJ8heZS3KspeCRG1GqrWMEzQIKgJoBWolM2FasDn2Q4waM
CUCMZHAQqUMedi3lSZxT2sHHcZ8Fhna+VlwTdKP4sCQhwAOvklGsUURv5HZXlX6d
8yWWt2wyD/6RWr0uCt8ZHgJDa5IHhIyM3fTTYSoyVDBDtIwOaqJ404tke1AA34m1
NrjsYZWKyptMlTovpXhuW+phNi5KjnJegLHKeNm+DQD40crbp6MoGbpznyDUJZoh
dzztvRHUAbAokhfUtS/ERBtM8hjtwwIGXNJZbosfCY8Ic3vX3Pc++h4FvCZAS/XL
wgBxaPVBJzniZQ8eN6TLNWnJ+ubSitdjgWSuVuNTxQtu58uNGy9/yInBPr71yN92
Df1et1hi9RzFYWf3dwPr3HNM196vsUxEHaoKUZ32akBuofMBYZsqohGxFTDUtyQD
3n8/S1D+HaHES50IsPeFQo+eOMW5ilz9fhrdp7j+1ua2HB8EUYApgC/wJiterUb7
rW79EX0FdggVmGxCZ+2PZcqDRg8bvxgP+pcY6UTg8umteCzs4P4BD9Si4LlfATtV
x/Skj/NHm604+GUNu/WuCfhVzXVxRX6xpzHMPBKEyGtc8c/G9zk3OlcFrYds8nxS
H1X/6IrikYPzVzktGz7dy0xjhLwkJFH6btIM9TpsVaJlifk2XgF/FDp3nLbzNBIx
yQw71OqzSBEHRrW39i314kdUjDwAVYXIiaMBET+yXARzATdytktux3ZRKKpBi2Nx
ARRYOe0a3xjVa/jFvaaeqtsb8tSKldlZNckGxAuwhsn+SNSugAfic9YY0bDLgE7A
qTkULRorSVS4nuGONDW2o78ifH/R0fjv+7H3oew8nf6gkOTd9UIHAR0QHKQ+Ug8A
fLWAONyGpE67y8TVSUrHvLAs+yRkx0GQvwi72/ODi1cmFBq8i4Xe2fw7CslTQsQP
1RaylI9WocfjidSMD3SJaXHegTepW+7gwYj3kEJI84ufoJS3CBDspN2CttTOXTVI
q/d5RqqnTzfcU/OI/2KRojk7HEPBu6p+PM1FbG2x/JfzixoTgH/6miNdoUFwMmF2
F0QRz0XR8q9+sHPdXlafInydVUaPZQ/FvAfHvyAu92X7uF/PMjZqNIgclhjNj1SM
gs8kFDU1su6S7tMEtPWEgFBTOk5NQ1mUWjwvNAxENZtpY2HNsdllC+aEgO/IxN1j
E+AX8ClnH6+d42b/AadWaWhWLaFjC5ApA8vSXbdjY7RqVGrbN3WHBRYsQe6UYraA
gcBRkadhoAL2a8bbsGnQHaQ0PsgZnEm+vqe+xv4ZPiJko8Wm7IXS9dnYThLjaAh7
vNUQbFprIx7hjne46ttTm21il8dZwmCYgrHZWPLNUTbv7dyvbQW29K1ZsKvgwhlC
/x+Jgizs3W/Gt2j99gjoHWuw+Yz7xAyaDu3yq8UxNnDiiRfBzpWbXPxmF1uy/kSJ
pUtFkwH6Sss/5aq4sRhNVxBxDXg586NygEq3WPrN6NWdZSCyiPXvkxCjTxYTbqKX
1lxo83ad8up4rUmwGr0SW4W3Wjg6x86atLI2i40Nuvjg3J3nYfKHHTwHO1BJYQaW
7013vpjHcDgCtVXRv2V+ZdfNcdirjOqkuYnzt+wXTChmYaRallDJTd4EFANMA8Hi
xsKZcRtCkoFp71S2sxEpuUKSlyF5k6FAFQ5WT2YvJn2ZpDqmiuNaXKn4nC8RqRKZ
jIhX2BYlz3D/c3LEmRZ4B/Yh/tuIYT08xiXxBMnsBtWRwQ3xfp66eRTxxaWvLCGX
0KcZkhpAk62kwCpkzwCrNFClnTym0ybBXK+JaM4YOw/m5QKiiNdHlZmj7PyryGZ1
j0uPRaxMkgZQ38qPg3Ye3VAk/9wMWEJbk2BCNVlmlTQ+TM92fn3IWc4cESIfoCXS
o0RlWYUXS78SgtB+zLSWL2Wyv16STT6SDsvdYW9G5a27vzuvRxVBlWBYE7BgpHeZ
bslincPxqBM4QQj4XMMxRAaVc5KkYB0kN01arWblxUpTKlZJPneTyB/8pOhZ4A96
RJX+OmwYdOr+Y8uRVNWJWpvqKplux2PRmCrpmoOARZ54a0M9FfStt0MfG9G1bdaU
oVlurxvuSDT+Wtq0Mv/K+7l19uKpAUjxjrf2l17ThZLPVx5EgMC1Fc5346zAAG+Q
gM9zBNVJd9QxoWzkXHqafeurclfT7DKjHrOHuThOfkFKJrIQPlnkFQv3UCPk2Z/q
Dqsci6d/P2AuOW4LlvDPyZ9Laagj+4DNgq5mkY3Zwilt/lSsZgT/gzE5c4LmUeY9
AEwwClxLmzAx5dkcWQwQDEIl1HJAqwZ9UWG7WkZcLZ44KQ+DSsfbNutn864YHx+y
HY8VDnvquH2qYE1xkwCuXlMZtHbgsDSo0Gar51KkfytYDwKDVt+nERq+jr9zKEiC
F5q4Fc45nivDViJ2bECtC8BS7hDSyub8mM/vJeELnsn2Z7A+OOpBqVHnt9Sd7euF
pwP8UDYY/owkUWtYDD+gyERt4DDRJZzBI2hopDo8gUzarz+7RnBm0wWrS+bvSB2R
Szq4bPI8NxpNTo1Y6ZNZW3mI4mbp9/tap/gsXXVPPkWV8WjgrT5kjwKomuFYCF0z
1lOMce+Aum7BJf1J0SSIvGpY1nfHDWOEpix6wNdpqe5SnHADj4qU8TvSVUk2g11N
CewiBtl0IAVRUnn6fZmIjxsb0ygERpkzOlH9jVMr4l0ThP7q5sZ769ivxXwan+S3
AFAuEJiYrKaYXyp9qbJJXxS3hyJ/y7FUaSCEAY4wIdy2CnXb0slrtjYp546VHYRi
ZbRhrwYLm67Lqj55KfRtfVS0PnrGwjwdshHXTNvmFLQgMH2n4m1jyH7sa/kdRO/r
c6op9d75J6Hr5nmjbAVZDf7Ca3BtBWgSJdtmzfq9kf/qXwhmSVtkQmk++Nyca8Kt
W/yg/tk545rJfxmwzhLZHx7XaMVjLp9qWpdfUHNFQoGSPuYCXCAWQeZBIxwOeB3S
4XBfUmr3YJGcEErK+Rr1Uh7QOiUFk7tDSjtrF87/7ZzNcgRUWl4ZQe8DLlTnWDFq
sL2eHTL9xE74HkxydgYK43Jkx+25pYPbRKBeYxcsduEgXDyXuoFwmP8CodvC983P
NxQ4c7otiXSxhDT7dwZW6kdEzHyhMtHSMTckom8gFL5IZ5WEaxDA+ckdEjJoceRJ
dyTcmuOtKe2UBvNmm0CqkT8PUrTpfwpIhh6OJsuqenKqTDj8/lZ0yBX3wlXntl3W
SGhPvK5Uim9FjZXuPrbvFt1LmzABV5++ydknqD7pfXOyPLpPGaNrwjD3PULNRfom
+tZ8cEoNf+SoBr4RVanDFNGP9h9dIySToMoRJwy38u/PmRjx6HB1L9JM0nkSE/vD
oNHcq+WUg+66KMVaP5U5HNtevJZIH/2LvlRDDbn5QbAnKa32f3V2o5H9O66h6urn
FyTx1HziBNsVqeq6WuOL+VMA0MHPQrHISVazYkFcOJ0LxFnMHM5zwqmLADsYVzSR
z5GIgToPFNkQLgEAcYMMX9JcQGokOo4uce75Rv0U0nXzpv20gcbE+1fJiEBcnLm8
T3A48KWG4gq6vB2o7cbTDY+0j+u14K5zWMhf2eCkk5LfTfhzQcYxXn7K5Vbk18nJ
ZTushxy7E7kWsuyURQdEz1AHmPEC+DDyU06rzivyoANJXqZFRYmxY+HwepCQD9az
XdpaacqxG5+QaO47hOocIiqujZi/j8+y8hNeMs04pwlgVekEDIoyXhUgAx3zMxPx
P+ZPFRgbszGwCe2yE+tAUU/vqZKeplGnD8prZ+7O2fUBHuj+V0Ej5OCmkllN6afO
S/0AL0GPc7hoV82qTelotoYel8PHVFOGeqtgepMs4QJlu3up4Ak2V4eGHPhDPzQd
mSI4JLTezwomSvTiZ3ClUNe7seNsxCEGfdL47PkUNlpJqcF+6pvZXWYejImWzBxK
q8NXE1OZFN/1CUXOi2JUnKtFRiXBoZJLpm/lRBAZP3ZpuzmIehTYEgNT1PHjq0mb
CviEOLCJGFKq61gv2pdU6E+e/Jr/4T2gX+h0uZvQrSXhsNHlEPQ02HheOCpojO6w
KrjLPfVJ1wLFIL5PznxdSkXSH/Apn6og4BmfZ5DnKyDGLJTBaVlqe4XmuyQbrARF
R3ywE65vNl2wpZhEg3OJC3QoK5LEBfL9LDlpj2aGUJ/UCOyRVYKM0UOzjEWjgNg+
fyxPejXOA/sB2CUJfhGnwZjCCSb2wp07oQ0ZpyhNRUDZ+xqPmNgMJNslMIJx3w9L
1s4eiuPFnYxkXgSNXXxHGmAPBAJPyEA7ESZmuXNIasQVulfxVUscZFY8bpD6qmhO
lCcIslD9X+B7QwlmldNuIBjSQvKIjLhS/qYYSC/4yHQoB6h8u32Fgt8QFUDbcCP7
FO1Nd/tzzaalXapJUpg1ixIrvbgo5sXqCtzXsy4F4c4tZ3vvpT+GrOr7k7Fsp9ne
8nu15dVfbrNuHwXAcD7CyVVRzZcnkHMc1I4U2B0nAUz14J/7bS9blxfBVqHAk0Ml
koOOHVpXQBBrT1dhdXHy/CnN/Wjcu7yS/FDmHBO5YLhU2V8oXxEtG/NNhU0kSXPf
W5ama1lcvyrwhVhpz7SlUBmaQ5PGChvbSO1n3MjURLLXmA1ESrajJsmyKqrvu5LG
kroAZp5KnYbZMFyuGClm5f5tH1oPgCxncmjgaL3fWtaOnNQ4mxVq+QLX9xCMCuBk
spd+RGQdzdSzrL64Ny+YHPHLq/mBKOd7InyZlG9g0aEpV8wl5VptCdXx89h1Xgm0
vbSBsYrL+O3ZMAoUeAZILLfHrkg5TzTKM5BYlNvaU4lP/5LKbd2axEbfXHRhSXp5
ELyQUGpFd36DL2IlzTi6l1NIH5xXjzbJOltmsnpfFQouhurUfcU2oMILvtqjuvf8
E20r8CyuTEeXGPauZk7JFm2mibhEn5yqQ62muLn+pgnqrXg/3iPoY9lYSF82Uc0o
/5yr+6D2ITTGxtIl9YP4KvB47qjXmv3kg2v1z0bU7UjnM94HRltBSejxjps53Npu
Y3+H+1U+uQ9TMCHBy00VAIBTZOAKzbmYUALLYGqDEBb5Z3BXW1CR0X93OLlCsj+n
cS7BnvP1nCl5b1SsczcRlsTomnJzx3DAK3d7P6FzEbqzwssrrfZ4H4NogtyV6ZZs
mBlKdffMF7mS3P4Av2z7VU+zukCD/26pXrU/BBEx3ao5NwJvy/bL0xYBLiODccoz
g3NK3N6lqDKF9URC8Ra4N+6jjf23ex4QCzIkloD7oxeg3y3OOFriTXdeYie2i0Rr
mOwcLfjzInq542MJ0JBPI7vOoRm+Sbn2n55mcHtvHws7qWOGFm920qjsTViHDmOX
hl+OK5dmWgoVIbyXVFLjlJMQi60Ud3Pj+Hg1aJIctodWtd3mbFYmO2pP+5OOPHWu
hNmpMCob0Y0TPHWs/ItM+VZjs6CPA+rzzdYfpQUhtP8PBHYb25GiL/VqQQEHwIJk
IoBe4jOyE5UcKqI39hjEnNNKhG5BpqaGu12HY6biuKlNpptYTnoaJUTrVGf/HDyg
h3zPPwnM/1SYHLCBr6++u8Jk1Si4Z+uxu4iQI1VY0x3l4neGAVxQZzRhFdIiPrH7
cFDUnbL+6f6ErxiA+TzIAAs7NLyq2AaVgbkEaE6ZBd8i2CaFo41UMU84OGwdiLuI
iyP9VpeVdVKzI7AbMvxKSqGEX2w5VQijZbxgKxqVsXOZc5GijTgyV38QPrpcOZXV
ivbcjQPzLG/uM6puwXozmteY1wN9rotODtEdo+ZmnPFM0/N/SQnDn8SjH6cHxfoJ
UijjskZ/RQzFMF7dk5QP4eXtKUaJ6fZrY3sVO365uwDFk3HNSCmMEyZKo9oILNqw
mxSQ0QuwkgzZCVIw8B/FLapWRjx49IDJuFclpjgnfHMbUC2Y7SrB5m5dfDwkVYYM
7zdBdyIVny5Q4kQnUX2dnuCJN/SUBApdUm5BEYDY+2+BcYSjP7S7V4b2SIfvPbId
r/VsCojNIz/9xxV8o1fUsE9K/y81qz/JO/oA8nJWKUqTYbqLLtrsrYfDWH+0z3AQ
fNSk2sqcCkDRAgGQMqQYyc9TQndXhLKqvo/yZYy/qhUC/EYq/0lms1+WKZuqYO4g
H36mutJlV+EgWlWsqYhdwR0BTi92N6F2Y+Pl7e01xBxQ8zEdyMYYMvFv8cmaOPvQ
pm3DMcJxD99Hr2okf/HP34n/k5axl1YhpBKI053LmqOxWg2y3t+6Fug2kXLaP6lK
egVjpstBHaHhy/qGvi4dtvzpVMzpr/CboWt1pzMWz8G95Qe7tiq4Wn7GFZJWEAJz
m/SCI+tj7K4EaJkQw4sruVfkKVeunRELlu8OK4ZD9Q/mkYLxinJuzJqquf6H0vyU
nXwEZCqO5TLWy9kKaJdtcfENJpsXb+/dqI4jqf7IQCLteTHfzTiCNVP1gHC/BhPY
USIxy6el+aj7N4rnQ8pyf+bY22wZB18K2TJlHLIbsTfQliwXfeyq/w2iVKhEo0NI
sFA6XmP+GvFuegSKPw/2fHRbMA8LSi5rw+dcACwQG0xPD5KtJ6DIisk5mamdGEW7
Z/e6SoHNQi2WeGv5e8k87fhihSDo0zTv0q/UA0BbRA2i8KHzrtd2A93XVMaP0aGj
uoQdZ5iZ5RMU2i93C+hX0sS1PbXkL6yNbUkphld923MtVXPUGvDqTZgC8m8TEgd9
y5kBgmQeGMKjV+UxqEd9JK9jEd6ys+fdCklUr2/002ZbVXdtKKeYKjaOqlAvge5m
qDTpmHb+9ShSPHgnKMz7DVzbnOp+MoLrrlPhj5Mrq5G9dK4Ewpm93BcVVL75iTTl
bsOyyDIK0pwCxWyhy0/V6RNaVpuYHe8iPGKiW4jS/gFq8r7FggT5uZS2S6HYkq0h
qRqqh0mJ6R0HoQObh6h00G+YIPPx/yGWXsJ0+m6OgOAhu/+57vcylkLCZI+J9riL
dA9KmIqTYix+xmxA+Hfi0h5g7M9WesxxuuJFQ/q1TWyFWe4RUEBKzDqYuRUzGgn7
CQFPXsI7/YHDCbn73mHAvUZ8d58zoHTjFeFfYhzX+fj4jz3QfJ3OpJjxODVNfEXD
O81jouL9yKk0rXkH31G+VbVJpxym0stRPKHM9+5vf2sU6RYD5ZW5cp3t3zL8eUxC
f4PGlq7X57mzLwKRWzGMs1U11/0BJ9Up6mErujFR+OjywFSps4a/uN6Sb6lMb/19
rbU09D0fMZuX53x5ywhoKebnTgyoTt82xfUx+l6fTaw0ZzE0WWm0BINO+Xy1chWv
+GC0vUjIfnv03wOXZ27dlaoZElAYceJ5/q2oocHC5aQG2E84xuYFNGC3V8vysA9U
6+3Sf8PBcndYXv9wZblpqSoG1rjHmx7//TRVyJhxKhOivQJ8uV0xUEOzDpu8CPN1
FSKiYBtT6e++x7DSzn+A4peaeK+C2YgfgdDQ0hKtK+MrhmAanT60zgC/vVIoKa4f
PBVxxIqZN5f9EHAV3Uf1pprYVioxdGnsdAgHFtp50HmHDpiby1JcOCNY0Hp6HkUr
xhhT17lGjPaqpKcsGC7APOVm22yEO34lLRaS2NkRYv22Gfly9uc89gRaT4qrQG16
Po0Fv0B8RsznJds4nyz3y4kDlERdKdv5sdI+/NKlgr8mnA4RCSgWq9upC6qxMjAX
uEdBuBDQz6D9QKA7I+9D0xV7I6Oq8bLMnMR35BlXVuqaAEW+1v7WaZo3l9GFSaHQ
2sSlBC9NhE0HsmBJddKzFpHgRYH8/jie9I4BTH28R0Wa5tQkzawJ9MT+YeB3w/cP
LndzzS9ENHhoi90ie9DRfQdj/ptyGeUUgnEJOFjZa3aqGXxGrsmA2m09qpjcPh4A
hF7BqTCKWFJfqwOGsRQowK4jaINRFZc4Nevghnn/vSP5PBn+74FK4RLb8PuOVpDO
xMKKbBHLjm+ch+Pkz6c1Vqv4BU1+gapq5vqQxZuNVS6+ywl2KBVnwiVXWcwJ+Gwm
oPWWwNHX83rHHp9KLuloJOeyk/3nVS+bKE4UFu4HLHsc/R2Y/uOSkuoq67vsLT+d
SYPfhWb9ZzBTWqEyUTh2FPBXj0haWJvrcGFTTKAmXCQrkjyMuLVsbv7VuZgOK7NB
AoHylrKZEeVyNJ53K5kVqYfQIYwX2BLs6mS0lCa/c0EI51v0baisVuEEya0PNl7T
ADLq9fPSijwZeViw/pDo+PQV38KLZkVUJCoqYEXoNlxGmMKG1fwogG9lBaAf5f0h
DYzTwQsOgNGgs/6gDz3lgQLL6HNukCSsmWVU+VVi6Pr8trarU3n5tqR2oOdWelLr
OeNp43Y9dRcNSe+RRPPdQl3fl+T/kqC4v/H4FCMmkG9hjLr8GHwSWDCUt2BF11r7
tgPcU96CiZCk4HzhW0P8l6iA6CSBjnPc/SCR3CJGGv8aAEjp/AK/wVU1hyH7pNQ5
K5XSD4wwicELoE56bHRwF58wvmXoXttw6h5e5CqAwxGnB4Ccn32XPKmS3Pq9Myjq
K/Jhg3XmOzEg1oHf1IJ6G93aE5GPvGpFcRje/rBYC9vvMdtF9uRBWm3HzRCAR7Uh
ruU9UGgkb2Lcj4fI2zm8Qi8RoRErLNzc0mwyl3UZfEe1qum6PiFhbxQTnRmYdqaJ
c0O1gBhs/TW4hO5TNUalVhqiwz+K5VJZEYK+0DbAbQrZA8Q/U6acX7AMW9KP7uGl
z8mTTXQhJBZHF9ysyLl21/msLCVlqJ+MQbaDBvZoDdQQMBafhA3B8/YETqCW+Ukp
wz3o8OKzr7ia9+TUugprhe06rZFy4+esPgr4yaez09wx+HES4h4AcSmop4sB1D+Q
wJ5CiTuRJ0/esnZg8pcKGIgDXlRLQsAFZiXmBH9lsQQkRDd31ey1lQQJpudvDOnA
V+YYvYFcuNcRejoX7o4w8eFk9F89MI2ScNmc1Z0p35ibxho0fvly0irSVPTBgmJQ
AfTcPyaHw6EZKJC/FdlG3rPNqoA8ribZg4x9dlBG9jaduuj3TTh+v93Sm1rRq3Ee
TWIQ6/Cis8w3feSWCArffOJEh9zuhzXormF3FvqiC64SH3EiVcPgoRMAJh1Fea++
lmapJ6eriN0rUj24WohiQd+rtZ3YtPoDME2bf68tAKy08iwQinkxvDkPk0lYqNVc
KVFP1IwJvzlnoIg9KDdr5squpmhlRNqw0NDWuXqTqy5coSpFWTZum896Y+zlIBQ7
PGXqVMeGbsczokMXqRVcjumxCiln9KOwMG4PGAy99/Efcv0kyF3l0FabpFca9kcY
jVxq6vX+W+NkUug4vH4FEZZmkPq1I/1PWbbyX5mCYNfuxRQXFMR7PnsiMgeB/Urr
OfzZVfow8byHlSNWmK0KHIPF/j/eVi6QJ0uIQLyLCoN8QSBVLIDHctqgm8OyGZ6R
a2b1tmNzhsd9WgOiPWP7rqHtACmIov4CzoenEFMXkncf92iVDk15DEJQZnnknHhj
dozGAd3BYJ/7/n1uQVAG3qOaF4J/VdxijNbHXp86i0h7oP9dFyKvzrCCdBFug/gy
BP0NFH25vS5gxi/8S854LNqDlwrdzxB2NSE8rNbX17R4GQvI7xfnnHH2sluCVfsL
DrMQkK5PuA6pFA+CJYvv0b4PAI5CSerQ2Xa+vfJvLjtkd++TALV3xnELk+8wK6in
HkyiPPJZYR++NAl8IeHtsrnLq4jOneS1OOVzUsm3ScgqiIg9rakfyu3UDx7tiqTS
9z3XtIm8e7RF214UeX4pCx6hWsA9HL193VGwzm4cjj2aW6hAEXf6OXybg5j2XdUk
sjrbDHhuaJdwLjgP6AGkhLukipWOBLWVDXBwN7USvwV1Mg7wDivAtznLNjyvbwbp
9Mwwwh58teF4wr+HCXqNe90K82BQ32SGo7kZ29BjVG0aghpLZ2fyFCkklxhxrPOC
Fbo7qFBUT4zABSH3rak5v9Ykl1OH/8apMPi/IfbivnOi4LPxp9xh/DQvbu3P5eJO
jgdjD5xlZzxKYm1KPuq5ejXNIFxcX5e+umlm8pn7tCVZqw+0N+KKliuao+1MaagE
3GuSMGkbasuWC/vj0F/JBDZexOXNCx7q7efB+ndnMWz83xMiatXKwbBFC4LAjxMe
F8aaHQI5xk6s5QTQqwh42ArkX3OWDpJGfc1Zh5S6KXEr49zk1oF6H6PDxqogh9YY
q6TEVZenUlpeG3qtlBq8Z/xX9t2am5qkiNtV6HqG9of8gENnZUhWvWvJ/ZSvEwZQ
S/BAvMcAwQk5Ihe3RCFy3Fp6NGfjR+TMuF8Vw9ltlbdtk8rYwS+58Jcq/go85M5P
csHP9ROaQaGnQjYmR0UkrVh8oUg1mTIN/4TOJYv8smCiAnbaLKvk7FgnOo1Aka1C
zif4hvS+NbVh/4aVBQLYx/0UHN5zfC8nxOn030UNREdWgxTwrY2jIR5h7hiqNd2L
JSuVveihnTZZFn+BNZ8rWA8lsQDEW0gdysLgyJrj8rsqLuwikwIVU0Rlrf3M6l5H
c+0HnPpNuHk11RAAZcyciKje5n37j3b/4ZnGqjoiR5fgAWtmAPyuR42IKeYqCmwp
W77P16jgl+a9v0n3EvC//db7wkyYodFp+ti0YOBH84aEl16HIWPWg4UbuYC+r2HY
c+pAxlKyGbMm3SLmR5uVM5xiVWF3xPKUr6tcuyBs340pbiBgzWxk/lu+rRoR6g6v
JWi5dvqZqjW6+cQ7D/azBUIsZ3qsCb8FUdMVGPhMkjBGqfDK/WJs1aUDl+iFSaW3
HPY6PAMO4ANRpJ2kuEZrtKrW/twL0Mj5Pke0klsH6+l3yo4IedkJCnEPXi1i8qdm
BVnnywgbtqxDxdwKr+keppd1Nw3Jv1CLBlvUwRIoMsFHLP/qT0f8Ai5TSg2LEgLz
ZQYYlconQnu68bGkTpU6Hug19uyBpJw1NujdF9KupViBVIb+kuGMd5hQTCOj3/+y
bpMltGEiRKMQOulFQ8e8IkCec9aQG4shHyKnLuU3H19R9akfqUcSggYKM3zmX8TI
aDf+lsu2L17dtjoOPEmdLpXsWQEnSFFCRyFX423Uu24WZMsFMGsxWsA804xdZV+c
zIZdBqPRVWz8BmznE1+xpIndhIwIFo/zbNGJlmzbLczY/+xi4dvazXU7p/fYGmte
P97iKQt6b3pzbIuAz5/cE0S7JeEgy1bUETZE5qNapRtxSCcWcQD5032eNMn+H0lR
snP90T4KiJxnPDow9qVkD6UrGyxJEBgEuyTazNoyKIn0ankzQHLvxpQXLurKBon4
WaEpzv5KgNqm3mAZVAxu03SXnW8/p+a5EjrM9kKQdNoKZ8kRmV6nR+qpOCmrGa1u
uWibu5mbvU0t4OUKfcEZ4V+126jV3IPL2pF+zwvUVcFTZUhnOCMcXArhUfZE0eku
p5o+a2JKPlf1luzVv04+N1qV7EPdMBHnGX6yyCFnG6zBa4kKcBp6D3OqYxZbwN/B
mMgFjA6ApMI57LOk7ZuuOfpwuYUQDxZZ+J6IbNHg89TdbSX1N8E2HU49ARpxBzpr
nCcVZ8FpEof7a5JbE4CQ8ywiHLOvD9Ec9qKpxNSfAOvWVsXZP4sSgfRwk3BdLY8/
hSqbcTOsqWFF6+1BSxFs3cHl4PUr1/eKo0Es1tNxTAaKjJqH2MyktnaHtCL2maUq
rZTYeCxE+nJbjHQmAq9GoQoSgBH4Lv6VbaLBsFUjJJunyDTX3HeYJwc+hpW6EjQN
W4Zftx1QK3uY/07UzoAgK8yCb2oj2HmVVeyO3RBqAHuDdxHZthE5+In3hOZyXKLh
3qZss7dBZGmZFJac8RAdC/qp8YPOwOA+c6weKxooGvawyQllXuJOxN06cQuAvz0a
hPx3BWVEyNe+7dRGudVNZTvw/KY8/89m27kK0JM3axNXnA3GwVuJseFJgNlD2CZj
kAR+R6d+SrP8MhAIXsMVTIs0qBq6vtqOpNgUE+h46FBzN8vF8UGIZZiNpad+cB4w
/w2CWXBdYlxG0vwoK0CPi1sW1WT8Elq56Rw3dabO+AgWKrsOZVnZcbZTlYl4Qnlt
4ZkCLbTaCVlO1DdDA7F71CfcyO7sAmc0a/MUW6k12IWpA4RJMsZqbZttB0cTpJq5
CPWytdiVLVyqBJbxaDbq3DV4c8b9UrYz7PHFhr+jNjCA6GjaZ9dUrPRllZIldvRc
qwygZ/Ue5xDGpCgJN8Vb4EaSxKMorJoXCMjJaXhRwkzFHf+iQQe/9LwW+rhbgSUF
4IxudBYcV+RxC+mUIJpxjrrIEkkQvBJ310SOLWCoQVUluvY7tqiwxFR3AZRvUdIW
zYDFtGxAotEmqnmtPf7daQI9q2NwfBbWlWOEYPcYRaU2EXl7+7kzoU/2j9ZgeXfM
8RXbqmLyD9+3w38EwAiJHzjs7ottRYGwsmciVxQ7TwsgKe1rRgqUuyhZzeg2J1Ny
wQuMPzbIX/OmBSEvN0pZQS50uZXdHWbkxFQKcn0x0ISsPtM+NJ7F8O/LP9h+hy4R
gk4GYNnk4BYTsoXzNHbBFJ+tuWDNsnncLrM1L8RU8ZZxwNOCQof4+sxK0I0FgzbH
MlgAnGPghO0fJkjXiEV8sl8DZX3T5UXqvE3WEO8Wc3NhWWo58tQwmK7wUzeKDJO2
fwBFkUJtcn4NfYLdJZPLpnCyplQKL08kk/pMQBDH2RmWjm/xPcripxI0BZ+lGY+G
5DWScLVvR2BBVfh6BihSfqfk7WO0dTu5U10EeP3w0LYP/ZKpDLI9lg1a/WIQG/Cz
ilDaT0pjhotDX3e6pBSY9+73ExlXx//ziqnicLuuSoJuvNd5JBs7VaoeYXrHNcVz
lthzMOIRYADCdZsPbye2mCFTIcxqHFngtJAZHfRZSPkPv76uHKhPPYjl+AvAIRjf
sf55mrWLRRvnYPUJf8uq+EVkyKdMMWpF3Wvve86fJKrZJGQeurhIOVUBUndzvuZL
WKmeUcgJ1gA0//H+Is9s7aMKfC+1+hj5YNW2K6zAmGx80Ob5aktV0uGDQn9eP+59
Muo6qmV2zusiBDCxdmnqD9HfV4JqkJTg4LFNMvv7xBRloIBF0Woo1AKfVonHcr2H
UmjVL7cr3Vd3uiMTCaihJB/3b/c1O01BxnL+Uh/oF8QvfbOBPxKtILetrDr/7aoF
I/6PYEMpNxA9vmQAUiatC8hWfmVHaqf5jMFV6/WZPegX8wHbXhp0xoTmzdaEqX7G
XLEljgmKJ6vSrp2dl+1TjalYLHwjakb4IBq6A4C+59srby04Fk/KMjV9/lOS3lhX
ZZZ2NG7gvHHNGZbSf42ljyn9k4dsQLu46DEUzaqfsvuAOJopWBQpRekw+I93AZE3
6iC7Y3DY9w4uVx2lbBHUhc72ii2eJjNB7Q/IoRPp29l9WrST2KDFaz+w8wo7yuLL
SjarjIBCipMUfJpXobaEIIJXPxfPvJE2HT4yoEat9sfk1MnCV8UAJ5CWOXKyo6CR
+rEelp2Uwi0XLiI4j2EZEmQwwETGF4lVnvmED/nnZ0iFP8rB04RiUUE+myuqcZ1X
br26MGy1zA35tBBk4BPj409GWF7702Cx9snM3N3stAogO5Y5bT6KX11sF1Rtoo2K
DW+85Rk6E6CfnUZccHnl3YXOCGi9hsX75yef1UtxZE5m5UDud1GRawyZu04m2PLg
xuwc69Rwn6yKZbI3WXxCvW22929eHcepRSjaHkRD/hwOFlaue/SdqYkMecpG+K/m
+m73d918naF89rgzIAfb+OaRhWjVA2L2t05IxAgqSzjfGgM4wlKdYHAeNbWGUSpb
kUjelMIICLFt3G8J5dO9U3PP6Cdz+lmI4gHBZQVGAiuMYv21LJmfb+kM0MTpsEOj
N2dypSJCqfpMcJcc3daBeklB7g3ORpoPir08WWJhxo+J4iu3p5CA+IaekbkYa7lh
ynMh2adjnqDFeM5FQKEMtEUlgoc6jJJb8wvRzhyQjLve797JGUKdGkinjcCTuyr+
eAKlSSe/QR0cLu4YDW5y4QXN9mdsjUSceN6wxDpNFuSMAbznNpYWX2gUz/ixD7nu
Jk3uCNlS/PtY1xmY5HuH7kZyWs89il52saPs01eOZPQ+1jC+ScU1YCHUK0seO6rY
gDJPY2vynR3UxrafpnRoYOjcUAMIplzZ1pY1i0uW/IQcPu+15ouFnIS2c/GLMbGl
5N9U8uFER+xGuNchcdnW6Ljhh7snBn7HYl/P5qI5hVCy3+Fh9ltQDmy2tgmnHoJs
aRCo0IYqwDyVvBgQjl3U7iqXu3DaTgomIrzSl+ZiJQY9D4TKWozLoPLcrGKaUWZW
fak0afgb15244t70h2k3AwtWc3karbqk2ClXXeoc9bB8EsvtxHZqQhorhjRGRk2n
C8GfRQ0MFE4h8KGItB+VtJj5VguDTf6bfIFrdFWkifpBlGwo5Edc27rBuQwOa1t0
YAqZ9N++iEG6pL4m+YhMbxoUIqSAdBC5e7WNlBmM4ZG07Z2WsAVAu7CItUCA9WOm
ds4VFTfEMxFAAdDV+W5WpNtr7v6qX8GX3QVOeix2N2bMbTK268y02eogEw8J9BYt
ygqr4AXFjvtAGPjnN6MpfhU4a9Wy9krwLWQ02hzml5g/2yf2NadF35sJ/tyr2tk2
rX4URNLmY5dE9ohwSCLtB6Xy9toNi+Yd0wVE9qGvUxpirgbuNYttcVb2ROzSvwF8
6ms40JBt8cjS8XGg+Ix5Xyj+DWRn9g0/44mHeFzKKv2U8QC8ogqKnhCI8LFi2S8C
y6BroKTe3gV9n6kgq88ZHdEdjMaUT9RBWFRzJ1E8cwE3cHy6BqVNruYsryWWy6Fs
6Ro5mkTh+4dYw4VKz8YPIRaC1Pajp/LGSTxEq1GlMFaAEiJH2yDCqFFQ/WoSsrjb
ypn/VsG1Biws/Mv58LGYqyI7R2oqwxBdEmVLPwIy11/+O44vpiyL0Q2RLTvVVBkY
VQ04kQ10ZxBuoPNKo3467+hx3M2c1NjFoWEYm4dgrFmJac15GtI+6LYgHACWnGnF
+zTZKJdKyjxek1/yY0BVdFw8r8rAQ0G9sxFR4Oha5zfRD4oRHLRXqFbolCTUbGjA
gNWHo/w1WHF4Tv5QUPba07/bbpTgS9mRq5jjj2Y/0L9BuUfbo9mU6BvlV9ETO8s0
TNZiZ9ligZX5d5vofzf8FVl9wTYg+gEizFarLILvISNE1Whs/ypTybdikWgUtjhH
lpf1pdOmSUYhaD4RE+bEczZYn5nGzL89wFMBeUBzU/CPqk8CX8cVa9WQSNUfcq8w
TrTbuxv1yEJE3QOx+qNcrCB5YzlBQL3zcOwzSGEuTRbsX1KFqB+V54TglxID296a
J1XzinVWEAnin4psSxMbw1KDhhF+GCxEFvpP1s2xqTekCDA6oPJaLEJ0hFeR2PSu
0dbQU8eFz0VHPFEVS5xa6LGArAXnVpKELCd/f4PpkOwmHZPt1DPkRLawlbpf20xS
5ZedYqwpGRShtU1u6LkKrlEpwYaOyFaY6U2voGkhy4H42bczTwrHIx+7BEujBZE8
dheq31sxpPDNlz4G8fm9q0uZaz5xIRZ8MI0ayT36LeaTOP6cbgCwujtYchSp8o6+
UimVgI/P3WjEwge2sdGWYtL91j1EpFDk88ttfyi/iMSLVcg4vx/0XmTjMs+psHgx
HLz//qdjv3bqlzGRwmT2EjPKyvjSinEzwVUeNeNB/9gt+EkKuBOAxtUMQKZoapIj
vbXUzAz1PxO2W18cOp2d8x/oZujQfmR9aArFlK0rtNGsZ97UJwlwD6aJGyL2rmt5
6BvepF3SZDbS7vrcCGEynzi+o9ADz9D6wvIkAdkIRvd08i2BxshXnOerjvSzpi50
FBt6lOgQKNRHsc3U2PEACJd/mB5mw8nX1fppkNUQs1fnCVr1zmu7sOAIbISbrYSM
55yaii+ryqATq+1lWScVcHUP/USyVxbyAJn9v2bG7yYVZ5QaBEg7zo/coST+gIMg
bIq7DinY09N3kjb8UcdHChpoNQvHeT5fXQVVIl0eUlb95V06IppMO+mYWKpl8jPI
mt8QSXuBWckaTt0uruwy2OxIdhWvP8niiM8VZpZEvAeZEzukCLgzxDJEJs0PMn/J
gUNlT8sV9GZgcFLoMODHxAWiYx5LsUlf0h6OBes6ZyOI3mI+LOhKYw2DMsDKMpS8
6fvAXOyY/Wrl4ZKHo2nnRifTle9NtLdfo7YLca1zWJK8etzbE4hpIHDMdAfLXRbv
PcaueVPfpdoHC8BFmbS0+T/g4Tff8JuMaopPKR9Y14ExKntpFF2sByg22FgeMYDs
oSKdUzaLVuId2hlVTAcHuo1xDSZlmfD/LWsEZpuxlmRk3dMOBWy+DpcFXJgqCQ8i
3cfobfBXUyJFpEvmOM/U1PFyk/ZDTLoxfnkXc44oWOQXjeNVW97tQwvnYntDjgYz
87Ogp546sX+M2h2qnoqx65dm1u8a5Wag0+2XwdjLcPvmYqhjNF7q+Z5djBwH5uRW
ULrLdgmX4hDBgNdViPbtuw4B8ilM4aH5NzPSfRZsYfnZjk6lAgM207HGF3fsH3fm
R10Ykk5DRtfeXOxGKBqYbtCoPKjqaigAYm5XX3SEROKV4kb9bLpH5JRSUK0uhlVp
TNNVFm2w9KCHNT9R+V74ine2fMwBfwNyT8yBqlikXs4U8psnWwuHRiuqrK5qeKo8
baZ+fn+PYM2KDIIk/9kLMuPBHIaXUVzo59d7rv3UFkZPPtTl8PtPrjcHyJF2hSjr
UxGvaYWV73KPjuex+fc26KqLtDT8wKmzmnn7Js9mAP39HmD9Qrjf6uQioHmtdDlx
7K6Yfk7+HCtD00rJekrpIbamct5X/g43ZFR2uYjZrEJ8/NTPduVjZf89bUDr3v6+
JZFO/80JoxugB9rYzBQAQpvqggngthFAWuuJXRxq46fUaQ/W3I3ok9S7U66dPtof
JjuITR+OBRqmm6dZo/plHEPp9tB7YXx2HYrqoEe0tQnnMnGF0mZXoQ8MwAZnpDuJ
Rfr14LF5kLqNQVPnZ09kj988wHCYwEnsKTS8ayhADbK4eTiIqbXfJMbqMEMQNUN6
MDkgyTIGdkTMX/5GA1Jeaj4NORJyZksZiJ5Xmu40K1VuDoJgBB/dDUaQ5P2tnFbX
SZJdm5e5jMm1vWsZHLSDq12gW3tCDOyPqL1bOvHBQciPP6SJOKoMUUeJaYEhHMnc
/DmPDv4/7TUe6cc3HeYXv4Er0jNxYEJuyMHYXxYCl5eoBdxf2Wi50ELkEJgLGlyo
49WfhKX0p9TWWm7N708w8HteH3HGy9JPOd/b5Mt/VfBSNd1I4oS+gc0dZsNwMGDr
R6VsSeS2ybFlouuK8myyhKORdCLw4NBleuBkuYdGG1HnIfjrXDbF66hbI/C6f7AB
/Ho0eoeaQ0wxLzm6U1hHMOto47Z/by6js/6AxTGfVq6CFWmZL5S/giRqN3qrPV0N
zdsm9O6uH91SK/xCGPBihPvd46Nws3kPQtGSWAGFdZeLjp+pr/MQvQoXF9awHRY9
GeMqDYomGC0jEXuGdrj+NpNBWH6vOR6tYtl34L87vPzov1CYJokKgK5pirGXD6d7
ZY9rCjOMn/1E/zh6PppYCSXFSfXoLB+nTtSLyKgZXt/PXGjRdfjbUFXaVRtzvNvc
78b0U57Z6nE4hMZjyWqLHb9hSzgNk4CxdUWE8+5ipZLqvJ0tZr0M518zOqv2jeEt
lqhy9gOfhwSy0nnH0y6OfBExIGlLyLAvHhhA+DNDIX9mR0HxvPOEsqpl5jfHUWlC
4kWnUvxtEG0DlcRnl2VrEVFv/yjg7iAjaDqKi3ddwTfAo6wgrZWUxZ1O/biLTi0/
Dq4rmfI6Ak2kpAYr+3uig0XgA0yb0uOMI29AoOofzQLC7+IRsmLufNTJqM0Mctya
kIkHgEZHrWaTlsgnnInPDPSXnLFGqmH3ecZwcwF/xEEz8OfInncPGWMJs0shcId9
ZaaarySsRVovDl2glnkDcO/735mHG8Jw0pfNZR0TIfPNDvGIRrq7EUIuxAK22/Yk
OEcjHa8ZgUvaU8FDILX80kNPF4nIcEM9TUYilh4gmrhGo90MyOXLqh3ANBdBwhR4
JLCpDFnfr2OB64kQlMe/Q0VjN/3qrAxJ94OZfsll2doGpv/eJ5EJ3UszmFAoE8Kx
5eOSgO36b2DL4rggAo0kLfp37x9Yp76RDFHhCDXLiiRK48eqFAI9LqCap1XPorEX
vMyYLJwaa2RwH4jV6FCgYZ32BYjPw8XmJiDzwGU25Eu1Llk8F2mtANlBkgOw85eK
Pafjg8+XE3nhgtSC4dlPrPdTMFgj+ogGH6JEG4NI/C4Xu8tobQp/YJ2Njd4doo4n
WvBhbDsVbM7RSqdljSzVgwcV7mrWTg1JBekSSb1w9GlvH2XEPNS/ODv5IxVRInGf
tjxaDZzwS405EKk6hkjPtt58xEsVbpoH8jcAP4tTPqF5yCDUEKUIRutqaU3GQ7Dp
7SAYHejj8BpnKP6l9byso+QD9kgxP2RbJ/Q6Au7SYHXnojOnE+Ibh5x0QHf0XOzp
kT7vfNsn7jTSg//QjXZ3ZwT/xOEJJ+qlK2wXJcR0n8XgdkIGS40mZ2KohdRkWnQ4
40A6jQReE10OI34L8Z+KVn9djO22ii+w/oSzoX/Bf2Uondi0EcjVwHX3V+0YeUuT
XrF9PXIMu2SZW+LXo8rAjG36U3d7SULk/y+7PqQBq0EX8F9ReKOQe0vu6OmeOtPF
lEuJrldr3ZHy0LW4yHqQtPI5Z/5xdL8ejsNiZ5Z8KoETCpjILgjns8UPfWrPxzKp
i7kcRhft0F/4Y8amSBeeAezTsfn4K6Xrx/xI2Jc198TE631lzGJ5VgQKjllHZmbn
/SdOOZyMvjROWyxgd6O5kRCNFs8Np3obQnPBGePtMu+hvtkTq2YBNteR5M+voQTf
TjOq5InuuFf7B2SB4Z9YDwLujaCqhU6S0ND1OFP6BNZ4jAgzqeilq31qpEgHrqDJ
bRdfu2ZgeIrHvxoXkEJlQUOKqgKEDGJTGkmXfIucscnvAePEn+hIpzb+9IHd5Zgz
BQ3gzB3sJRZW8AftjvThNMgq4QRgt+8Fyhhsg/DElQj29fLMoB2xTvpyMrVdfc16
nDYxHSZaVi4iRe3JWWxCVUQvHEbVI7GP7xx02ez2mrQO2A6+nSW05pUtlVgTCU34
MjKaiQfJE4xq0oO9R1LoI7vVlUZAZWgqpni3fhmsIv/BT0KqQ4UEX4MdXCCawSGf
VKegreY+qseijEoI37ADZAkK51qy2Vk9fvYNxF+H2gUatNBuJYgw3loas9QZ+S9w
VpWVGK19rLDkmx2AWPfeCzS3/oLn6ZH6I4h8c8tIqvkxkQqgSgTf/Zuy6H4cDPEO
l9kIYBzdZ2n/I6GZSe9+QlL+lzMA9iOmoS7PbUWPjbKK4SzO4aHt3G8dAx5xkEzH
u0VJOkmT50bO6CqwFE9Eag/VvjwrGdzlbNYIkBaFUWOCPPXR8pJJPIGYXWpcttM4
IijNBG7GbKjQak6+Nx3OZozNPyoTLvUyoIQZH27gzaZIEK1U1/48VAGBFA0fbIpn
wyZ/pk9Wivj6oXYo6+voTY3v+OHhwHIAjWXQWix/eZnneIfOqbbjBMeqR90aRqlS
FuYQwumOBVLB0eFe6iPGal43vrYRnq0SIFjU/r/T+gZoo/siYc05TPVXHkuCmi15
0JaiW4DNDM/BWYl4xqsjAc41YPbykz7Woh0+OYv+YIzr0T6CnPleHYRe+XeRHPCp
Id2YhNQebp9hVkbsRGndvtmUOEZIdQlSI83SnsmkeivJ2iTEEVvDRr6j2mcVgpVT
S8/wc/kZPN5yYVRVyf/X8h1UJvedZ/eatrNWxmMmf4joEeVmI7pUFbWkIrzcieNc
qjPEiQ82PpJoK3KopYDRCpVbVaVZ6ydqxSys70Uulu0w/iASWXeyy/1qlCp1+UvX
6sYC1MoEn4s0h7WAz2JxjebsCuBvLxzhv6oV4JX3+ekv6JmYVcwN2CKFZ0aI0MS6
5/LKHrG3uQeeqpuBj4d2OP8rT9R9wSrk+Oc7Vguvb4zFKMOLBiDpX3cjmU5VR0kh
96w0j44aEYnrOAe7xrmTg7fGmz3Yl6v8Erc0KHqfSiO1mfysrHE0lV+dmaQUJhuB
CcOdjDM7H20NlyDh1rsYAyvsNVI6YaCDZYZEcSHByx/SAGAlPErfYO2ub6fhmIKm
7UdATqEUEOCCaUoM4k21HEPAT0gj3H9n1MDfkmedp8IrBYi5fxe4Xw2ONsSWbyFa
5dRUn5qlh3Ogb4YxxuRu3yceIoWc1c6NWSEQeVZw8obwCc/gR+/BCSSUwJwiJooL
SZNYKYEiaeDqxAivwTo6XWLAWoxcmhTWhWZVGZvTaVkWGOxiWiv38dIb2Z5bf8jW
LW+Fgea0gXk/36UCrqnEbsUnZwk1Q6K/frphSyD0yBPsNs5aQdZUR9awqdk71yS6
HgwsCFp2BuFIaCesa7vuP2ExgAGOhTMLJQqZ9d61KB7smxCZouvPn7/GaYA1SUOf
DnQx5bW6RtCqMRP0HB8HvVP0mNutVYjq42jQQuFFNuMZPK+/It9TTDX8TdvJM1M2
EAhDnoCj8NRWw4TMCk0r/NIQCX2kUbRO/5xTz/CSS1MvzbGZp1rZY+wuv2SiGvYq
PKD3MJ761YmhwXVCUPbkQ8LTOya16UOk7jMG/hVlH0Poda///6cZgNfcSDrtgGPT
ezhyS1IN/mIo1emEds4mqROx4Dal7UGhP1MgR27vXfljxskGiMnA06yyyim1HrvK
AbzKid/EQcRma/pkRFsR2yxDrx5aXP2BZf14NVUUmGA2y9BXW4cCzKb2F4ORVQ+b
7g1R0OZkZjUyBvtogwyxG1W2SZJC8vv2oSHhGoIPbKsi9XPSfDb3y7DBlJir2FDY
5qel4Ko0AvUBDBx2F71iHE7GTOgkOvX4NuE6OM6VEW3KwKn8FJAvdsrp/fslmclx
esG5wRZHcPRsUc/bcCH40K8/9XvFaXGiIPmhGuVsHCNI5x7m6RDpLOxPP9HwMSi9
CHRc/4x/wG/+lU3ZyWnsv69W7fJyN2UrkTLqe4vmy7YDzQhi9DGudaOBT/BB1IXO
8WNxujW25RfgBxynSrETX9iZvMLdzlqElCvf5FpWXBhLYDSV3BOeCI8t11NVuwwu
G8vOT0CXT53k9Gc3HOr4jFQYodrvIvvUSYrdK8OkEEkjd3rCr4WG+FzezwAsxq0c
sRj9kb5OFBQZhnbiYTSenittSDX05fVV2wqTBKteM9glCF3basnhbCJuKTNknmpj
14U4YeIPpNTfAX2UoNMO5E7pOH6XSyNpczrjWFBG2zUGg/HNl7VKbdbcWn7FN+kH
gmvUKEm9ZIFk7flZCMDWERqy7YknIETAFvC2L7HcpKSewBKpDdISPaEU1WfWCqIm
+9c5r4iYsT0T0FQ05mhrslpv6E0elbpvDejyrgB8EmFnruaitdabe7PY3ipjsOrN
kqtHdIlqNznF2DJJ2QMiR32vPUDzR1e3dmroF7uTTjUQvPATjyBH4AW6igarzCU9
9vjMD7d6sVIHMZdOCrcq9Go45Y54w2HK1DEW0SPMYe1L0bDhdbJGbNP0yhoZdNWa
0/JNm25w8+EhUDmFlTAOG0J9GfGl0ANEpb5/vqSkjEuEA1Vt+HgIJ7b5NnluClwg
63YcpffavaVbxSSFVVu78neavcIDr2i3U71H0p2QG1+ct+/npGY9oZQGYaqX1gqA
xgmIHom4CeKIEJ8HXjycFsRRJMgHf8GX/fwl2hHs6RMbsNunTHULuz3712CQ/DdA
2UvNUBjtccx1REMZWzwxv9J2VZ5dv0exjsGK8+F/1/Fp0LGUPECOsJm63VpNBAaV
tq0Y0cLPK/DakSh/wRU7IxjEyovkiiFZhRz6S3+JYv9Y5R0GR4u3Abts0LcGsfVJ
p6aX36+TUQOsE5WKV1IelwAueER5ai1YNWp8YhRSAtRi9idKGo3GiMOl84vm67e6
rw3midMSTmognk0T9cUIkqrf1sp+tEf15za3yAARA3LKYhqiTh3lmzL9SucPL48D
sS1MLz904Ml8Dme4erNLhOOTTE1YH1Az2JwmVy2KXPlh92/cU29jxaXSQL4oUbU0
XRV6KXzJR5F/oxeu8qISc3f7PdGNYBfyqFFRTZhydUjhOXnSgWczJJVo1jh6UIBB
HO4K00dZ3MxE2h0iPmyC4Rq+MrVFXrhR7bwcY6wwlIWjAFGquKbhpYKMXqCe9Nof
LNO8u6UuVPcsdocEnKeWLNJDjGLz3vFtndZWAp8nwpVToCpZRdhR7oa3mmE2dbiZ
cBiwm1KNzzW3zRXaUgIuLBJ2Vs1I9fuvfe0AKfKcppYhJnn/f9+x/6ebBYzKh9WR
p3pAqvBMsV5ZyLq+8H3SOqEHiZ8k6eVbPPcOlk2RGd1z7ijjhnkbmYZlkQGgroMA
02jq6Z1lp2DsmvIKFVEZXI2ukKkXTdPiHHBJRhe45jLoQdGWc7JQrgFDUt5rH8jR
BaJfGIOHoxiZciuvGhYMVho/J20F9pf0hr3/CeBCNEKVKxjfhl5Dkav73k7g4Zzz
fw4t8JJbyCI/iiFFrGTM71+THdnAMPYeTFDpxSYMNc/56eaLzyLkvprbcnmr6Ce8
Z+UqhqaB7XZspOIQ3J8WVHVjcWIMqu5yKAEO2FscS40dnYH5ikOoI3l5eN2t1Bkg
w35vwvMeqt4HYlvrAQifJHE7h6JVHo8M3zkz8Vd57L9SG2Abbuyehp4pClJZ40sy
gqxhLYEd+O7e+i2M1Y2tNy2FOTFSBYzPSgs6RbiSbfG5EuxQJPOdRVysb0iYcCOs
P6qdB2JgAcSGvtbChgSOvWQ9pMAqtBPlq92ATtn+6IrICu76M9lVfoqTZGVaC1hK
G/uCgORNENuIH0dztiXGptFGIVypdfhX5GCV4lgRdU/m2/cEIZSKqVsx+P+MXsSv
Jy/4WcrLOsYi3+y9zA71nHYoPb+aRVDDFDwuwiq1UrWvCyiiZgCtlkT7qYDGxAXy
kj0sOc63kYz/Plzf0QxJepwsWZWGCU3ykeD+mcLlI10A6ijMSnScKoaHt0ArcFlq
8TE9W6mu4q2wLlx9SHEaKWGRt+D8sfvFRm1Pw4LMchmUXBvfgmP2J3EH/tV++hOr
+am9nyd0RAyHCDYcEdstilGdWa71asooezzxJtIfqLdZFr4Ysy6RkJIPCQaF55aa
50Q1Ah8XwzlVBRWn2b+7XFQC4DT2BhWYdAkFG6PyNLMvUYamP/alagp64jLDrr8g
eP61vrjyB/WmcxmXt0qWP9NWm9E4z6oVNi3rVzTZeLL0k45rclJUsuSYvIVB0hBM
+rcrZ56WKX1iuhXsZPVrXTlmt249BVLg3qRPe5jLvvJtXAHnULJQfwdZ664825kv
WKbCa9fIgR+sf60xLrHTj6dXIRhohWvhWgkx9Nx7xsL3N4JlyeLV6BzuUdXHD4tb
CHiLnuIy8oGe/R+NR22YOzGwuFJjDujJDCr0K/6OVtsNaWbHs/H0jigyG6uX1cIy
s/8nN7JHt7VuS8u5DRdiKhVSIwfUY1IrUReeFPn9/AraTOBTg+x38dh/DGnTRTvo
XAyRIQvUz+GGZu3ofzy4P5wNSM1JU/MuHx0tgbGmAGNtz0fho3jtxQ+6/RuBMZ/P
h8VVb66FRMYUUyBWe4ut+KFN7jEI/g3Qt1eQANshfFIKMOt8PrJXZzPe33ie0sHk
/rcZG4tCcl+y/IznTNlbFusJLwn/xMvTa2v56nXVoVpLFVD35POtMgR6t6y84g9K
79L6531YTcpm8raXxcpzu7O1erhim3xFlcl34NwJTb7stEt7xAe7OfcfuJTg/TeL
14LZbyiYzU2GejKYRIm20WUpgyIzQM67AQvoErW2pcOA/eeLPEbQk4BNkwHr0kdf
5zBGb18ynwyWBwffOkWzDVrSrapj9Y5QspnjQT73KUIhsjK8hu31d4Vgq07X2xev
lb6msPLWlUIMtFnRnukGdBXd5bVyg84Y0YQ/0eueSu/MXtBbgmkRpV0zE5NwQ3J5
PrOAR2SD189AKvs+b8WwjHXdybM0buvkLuHvZGLELICtoqSmrxQsyj0atDEp9e75
3P4nmwsPsnj+MQfxYGIHozJymkzhz6oNxjDd3gfW6e/vonx3ntjRfqK4JQ6xpY/K
FO290Ga8xf7L+1M6z9wDCFH9PuUjWNxwsQNocnknV6MR5q6G2QGWADDmGeAt/uQY
1wtjJJS7ygMMz0eIA4QfpBC3uV+nOtCMlINHE+ArhV4iyh2c1mU1n4jTfoYRlu3W
9+QwZYfvkBJx/zNgf6wsyAWA8f9A1lU+/wC6rkNGMyZFsB2lmRloht/ZBSQDo/8M
B4xdltHzhcjLQ/vgazRgcDCoZ827J/5GwKj1r8A4E3BqAScyYTtczWEWiyrYmHu0
bSXxFbPCq6tny/zBYbauWnCuVSD4D7DHXBd9SfNGV3wXXniRk9/yw52rOOA9grHy
sfQ4mr7B+gortw4RgsiQJo/yctAnV70tk48xR/asMtfWG27qee4wOUIos4xI1bHO
MAQ9bxj3LFofzwuYafMflvDCurYRsE0BMWZVR34H2honMH5ZUQbWAUj0IgrZubv/
ZLNnumZUgfq9SRIZfCWy4utLpzvKKabfTHmYwUHBhz9xROl/q6PRhoRrmgQmJ7vp
JNjsv2csTtYaQ3t3WFvHbCBQDYMWegaxkiys8ZjFjTDQJIBwNxn63fyjjbhdTooE
VYx5t6znr6VdnJhboGVnlWFQjaPhEcmSf7HBrbk1/1QoaiZ5p3KXC9mnqg4EdcAc
o+uujjhUvoh2VYaQcDBYUx6jIBUzy6pfJFpVBLlPNWKBp6WYnk3tRrDzvV0WN52G
gitfWXtjHPKfx7v29jw4f8GBDX3Ixm1pcmmPBdYXjxap/DEZntHgE/SEKAYtc/Ae
u+g/LH++aS75HZk0y+M/X547lamvtEx7sLhkD5b+oHfe4CglggiS9ycPDenbXqsM
BEanAX73ShkyKQT6z2ADsKLJodgqJjREJ+b6rN55wBQYqDOu4fdItX/YlvuF3vL0
VjNzKMmiUK9Ys2EpPfUfVDBMywAVXnA7oH3fLGxCwrnSnNsjLvhs2MawwHo2RYxb
DDIh3L9g9VB7gytNBscbr+n9+EUllylXWDsWO8w6zf5BBTIbyUY3B4HRYHTVrmci
jxST/FDH0KhnXvBSJD6w9UW/7tbJEXQn7VFZXRJryoFrsK6e51SicfZUbb39WRr/
QfsStimVBdUTQxM0BLCzhu/LDjCz6mivVnT0QaZ3Ij8JpeuizvhCwRJ9yv+Mz3Vt
SNyHvmGaN5Zm5VFhGlGDvwwbx2dl74lIDNU1YC3/f3Qy91V/iKH5DjBYtZvZ/H1Q
gps8hf0mpBnTkFw+XOY4WSMDjv//mJg6HsSUsEbUDxLL9QCinfoJed8zX2WRd6Wy
xL+wlW+ANP4uKw8nIVKM7z9pZuoU91EP1uhkk+LX3koXo3t1MhTvqgVw9y1LR+Z8
RFJNHkj2QzZyi0RHKawZpAwSSnUJjyLviDcN91TOPNxWJixLgiLJa0eKO0QuoFut
MiRiPGEtCMuO6L4PUfNaNi1NlZlq2xAYqvZkfepBACl+zyY2NjG2hWWR3PBG8Bsy
tkyZftbK0ulAeZ2SpDMC6iu8Jz3rbGIcgd8QXhXB4aFofCDqNSRTVEwgnFV1nFGr
c0Yuf3hHK9CsbKhBMnExBemKTRESNrAtBhstUG2iqKw417OUogMLH8cOMHmZ86vN
aBnt9NlRWxGrGIQRSnoSfTMKmbHOFLKRd22alM4ESpNmuTktX4SbNIMFzAP+mdE3
W8/CNwyxmTfAiJUVzt1Tsar2I8EsbxaIB5V/3STfhlgMLZf6XGufo0DNziJhP3UZ
NWjCKyPozZYR8FTf8qD23s3f1nmRMZ/IiAp1VXyWR9JClLuD10hE+9EiDOWjU6d/
+UHZKEZGG4yE2iKv+WJD6ShoBPBNcIBLqQ6FSyO8/APU0czzglSf3Ne8Bh9Gb0q0
qWgsGT/DBs0zyB1ZdVaHs+r4mpTneKe62gGt49/myhuFhCH9Vvvdtjq4WzuzxSfH
ZK+5ULb8VlhzkFgC5yMWJyO48U+FW5rlmUGbglyeRNnPQ6aEdCbNftmMaEBBKH18
W42y9VpgDpI+J5h6Go/vJy8+3ZmUcn+Uac7DxKKdRcBHz/SGTNvy6vpmTFA/2M1B
Rty9fxbHeORByoAERxE0TZwRFFHFuDnNIChQg9Llrkilg0pAPWj3jpoagggApyYs
GmDvtPaR/AtsTIIw3k/TnKX9n1otbHw6EtJDf3Ru6gm1eZWPPJF2u9ol1XUm5DbL
PCA76mPBq/awm7SBzMe5A6ilcAComOICLhJwrmjYP4eHEpcRTUa2VvGPhKUeKAxw
fQme2nBoGxSmhXgxsiqR8rDR0nsqkGDRv5tnI6QVW93olh42Q/5naMLy7b7RnAwm
uvyVUErh+hrsTjSWoQvSMYlNxTyE50s3pB1jVxXZUCvqwQZ2fenHTp3WOvSUxJc4
AACxrsBHodOao+dcCXuLSVbGmOsHcRPrPpcXq518Zb0OQ5Ec7sLp/eoVvng6/2zQ
tFgRBd3DIMPTgkwokT9/LojdcnzLBJGsWd7dBpuJWA02gWzLZl3f/bK8ceDfFA6O
AsvC1oOUarVIpSkrUDjpXFvGV5UQcmcuwNm7f2X+GXr7xdwEqxQEMDuzo8VGlSqh
jbiXnAL12JLZ0NQewQE3JM2SGPyzsY8wxGXSEeb00iH7dUXRXd56LBfXiqqML8/d
lEt47Hi3J5mo7z6QC4ztuBNk/xsvrH8p+4GywbSpxa4DrknLVmm5UcvzSenoNNCd
7INIyIce9WC1j1GVkAXE4u9wrZB+0pQfOZYNQxdjz3OLkJ31h/inRTkyAccm83hy
9mkFvINuH22LFRb8utPt/4WEAkwH7+EdyZaOJI3wJ3iDcrPtJt7aU+zEzAv5o5Os
ZwfsiBwgJtRT62QRzWbSdWtx8aAV1LMwCZXsA3JF3zJ5ILAtXtA3yyZPhHH+WcWc
5h3CnoOyk4W4RgwaW++1lxzbGFK0bPp5kpXs38jUEd+et0AGAeBKW7POalwGz3QA
pCz6bb5+vI6mPxs1E1uZ27V1mpHfc7rDJl5boJKiCvQL/ds4l4CFlePRrWD5OgjX
AHubVC5W+52qFtjUxUwGqY3jW+SJ5UlSUVJA/zDG25smh1GX56EUKP+xf8tjOfiq
9tAFmNLmapj4BfFGVHhK5Y+QgTEQA5iKEmOW14ruJhUftMwJEK45XCOTpkrnKcfR
hV8NSr2wTelosEYN/JYyHpjMLtyYdgHXHXts9bhV1ihUvHjUKxyQoQ/+JzC65LPE
QetBrJpoehSJLr7dvLuZOlbRF90rtax9NSe+vVdBY2ntwtc1h0bpyy6ZAk8/D3hi
SitLWJMJrsca6x2bz8lrPKLLH5ryojniDhHcA63E0RHcX8MHhX2CwVZnIYI2emPo
rsEQlEu3LajXreAS7SlpkcFwxDdhwUAtf8zVV5FAN1S4++BLhKoGLifK1mTn3rdk
HFl99PyXZmsyr3OF/bISYBZhJ9qxo5k6FH0wKkLX4DrpIt10t5WO9IcYJGiS2+1H
tTonqZRkP6GKuPCpaF3bNwD2veTOTcsbKKn6tuZIGVSGcu2gY/4mBqSzqRVnwFW3
g2Vo7IdNsZFYGrZeSIBOWX1QDJuNerz+CUeSpiaiS6vcsW82nNcvot3xkB0xXjHv
myuX1NnRAX0fI8/gWKyJTzW7eKqt4UGctPhe+ueBfKSw2zESHAkYJorJRSOq5L2a
WEJp/KthYM25T9qH51hDuo4kGrjBk68yccFzrtw1uF+vMghv3z58Hhdac8dGzZzO
FXMRzZZvndIP8ZKj4RyIkUMuauUB09TIYD7iRQNup19f31OCqBZAcZJzJZ+aqS0b
hOOfM3EiPhkAi9uO5pAwgJewalb4XYxt1hsykB2rtNSM7lfc72FGsTENRju+cbUV
RhmFzbwVhnwPjeto0c1YVPgCZdAYf94jJfOj9fSCAnGgbtCVOHX18vaC1Reem64t
5WXqUNcAWES3MVWnn9617XZvs5raRAoukY2NBO0PVN7ga/8gRCvxEymNPM0CjRth
JgFR2/iZWusuL6Fu4PwtHjnPFyBuQASenpFDzLMvP6RWIKz2AkaMTTaYUz/EsuW7
3eTnewEDwtlwmuL52ZgR8SE6JNLuzLxmAf10I0nc5BrVd9RthM6odV+UJBmmotq8
YLzXClSpAg2sQs33gf8bmVY4b/enHbIwiXpxiI215fhlXGEeTP3PycQL2g8XeMuX
+39LCVMIAPJQaMHmsS3Zow3UhscJruGgUII7IQ1BUXnme+oD/nhQ0dBAcTp/8f2r
DFF7v9vfCXJ5u8lM21lEsnE94m1e53zVM7tr+RVeUjS42a7aMNBIhA/sjHYLAjtq
Rz1dtCZfGyINYXoWZna9nmAY9lQiUY5Jp1/MEe5SuHN8U9vZ91Qq7nufbyyDCmu9
WSLd4cp5M0AvPALIQHER4c5+BfqFewPpn0O85R9h6+d9Su7i4kcM1BVD3Imem+i+
dWwVo5vnAx2S2BN9/knzStOvdhH5pamX+48oW2aeYwsTj1y9TQKyvzWKhssTce6E
UcpaeQ7Y3RveljqpuL3Wcb+1KeejK42h7r27ss4nwsKYO9p9+6aeOkEzXvptRpo7
EucJml2f0dvodLa7AMe2OVv1PmY1pCu7lngnLnfs6SNBkeD88aoP+DBl/9F8AIUn
KGbYao11ym7a3wRWK91bPdxcsLKQYT4etRYX3TBho/z15EJ/pWjN5Z42eenPEQAe
fASTuO8vCz28hqbHNZoQU3VJDU/iL/GdH89xwK33afPq7rYH6LRoVy+I2FoCk5EL
EVbmtchD5BFPRe+Lke8JsoLTSbYp78raDvThtONtMSFj/5bE9gNJIatdPp4oJU4D
yfu5P8UTMnUwEDpKr7oH7JMg1LdnetKEK+MrT8oXql717F/cq3DbHFPtchix0Aal
oJhciOxofeL4NLAKees0TLtTEf25Kp28eCPGnbivk+Kwv1qlz1oOJwJdRka2L6tg
XtNkiV5DFZVQMhMQ9zRIXUHec7rToMhV0RZQUk13+oj8OtpZqUWTb5KcuLqx8A4s
Vhpi5+Xudb+g7TPTp92cLDMplliUq5Ob0h3yCfJTsh9bH13625WpgGda/N8Z2GcV
Wm3u4aVloT4N/qePmCpU2pFGivKHi2RBzgYhwocICNeRIKTADBYurCab9c1e1CRO
3dZI9LVEEqM4BaFedQGX+u1pDc/3ftCBfCwGhAUL5n3U1QCG3PTnL+TpGOSIJ0wl
gcw4WndsWelwcFYA2Giyl2E7Ngm4C0bPvdnNHeclfuI4DdN0DCfqLENFeLsb+h+5
GzqcmlkPo5VgLPHq9vhjFKripliJr1bvwbdkpv3vSY1gOb8gbt102Y7k7w+3roZo
/FWevzJ6kn0JE7v8MsZHGdP2ifmeHMBQUjsMULWBPJFB7+Z3fjtMVA3NO83nI8XF
5MOQb1NDTCRSvOcKCVRR1YjjxS11GowOjCDKfKtJCScxBNEFWMCI2WR+zo974PsP
0AlAs7IzXu0Nu2HMpiJ673ZAeiLcgGLLrKSE5mQgfw2AQH6ezWUh5CGbMCCIHLo9
CHjEhJ5MbVkoo+RYjhaFi62BtdNXrNdONFN4ZbssjybHxE/ao7dutlpg3qrx/v5v
CdxXDsMEMm6ikr/Lg7Z2I3gQNbuJFvoAeNsij17RtpJ5fpp0VXzWfW9dws+ecJJf
CksWCxaWhPX7bGhblXcgH8j6zAGYhAMdytX4Jh03ZOal2dAY7+S3vhO/v/ePExZ8
Fk7tUMg+ArLyyGDemlbH03dHrCKx0nmmtYtgsoEIIaiVMbawi1dW9TGJxF1yT4ib
CnVWUJ3NCX0q+A4+e7FFQCQRZdXzKWNFY2wyU2H3h/nyh9k1AVfbaEFR3/NGGpVx
jZTw5XCv4n9AK9zrwOxym1ofzRXbX4P2Oce20OQJJr/biLqaywa/3VzMLi/zpuXk
i6W8vLejcC+wPgm2ws8TQCiUPGzhBNPP0L9DXN/LOTHxpstJeNJnW2sfSbVQrdIQ
F3VsrLE2GJaricThpWqEDtK8Rte2sBE5cOkI+GMrQ1dI/8/Muu5nvNmVxfaduPz1
WNjN/jOOflYf53VPi1W/PCIplQdN8lsQoNAreHJRQ8/05dSeFVxVbs3xWCZmlaFe
7BO97++irzHMfFzZZ/qpvDBSsOjhbVK+7UqTBJM+mb9FGek67xcR/BPbhrthWCrA
koR+MSwqiDcspakREGBZTa5nhKPT+ZY7pAqXNZWrThK9Rv8BFL8UdIuWqEW2piLl
oQ1a+ZT8wGQFI1rH1qcyXHe3YsDeOy70T04ITvx0fYDlyTha7iKUwXJtxlOUTT0A
wdejCLl47pO5zaAOzkMqC5VqI0dSDJcza8DJN4sj7lCSsR4KNQAJuqGNAjXvYI6Q
bO+y6E1bVyJ1lMWHMtnTXLVTjffJGcDTk5vslEz1Sq12Tyh2UiNfxWdPnKKAGRIC
xXigp4DO/Y1xaPOt7IaYj3RWsTAD8LpIzLgNDaBTV2tKYk1mWHfk6OlSGJmrHud2
AKEXz51P4k/lJfvCLVps+1vtyaXyN7VUWzT4VISXDAzqK0lMIRQ6RsmQvWPQmFvy
iajZYRSVZQKdE77kXuZxBRJtt5tYOATMIVbyiFiT7tzgqOhLSWjvT46d7/bqwAg2
2YFYhKtyoEh9qFXbzvNHnCpXBZSDcy+xc0YX5ROZxiPtnmCpLJyHGhHiv+GibKHs
JDa2SObMURSce7olRlboBGpZ2fOOmJtAmHDgF2lnQSnYLI/gduZfbZoAejJzSGza
+y4SuaO7pcRbqUVVmFnRq7JspUlst3GvvBvItmr/8Q+E98vnsLQjbHUQ6TgfVWTa
VF/7Psr1qqKxOTptmTpWOHCosdBjMEnsVgoor9d/sJrOnxQ02Ay+dr7Z6kt6v/SO
tYWLO3sz4z7DwvZTBfTp7sCFQaaaeZO9tPzxRMlSp+mEPH75rjfhxrxPnxjSX6uL
c8hMszL/FKuySnwv+rlmBwcHNmTzSXCVwRnB1bkbn4GcZ5LFGCBbPw3ILzQGmrkL
SMG5L+PrS0VS4rXoKlGh3T3AQQ+aeEN+v2mYgVAZdTKqkIQ024TGvv1pxhyHkf/W
0/LegvmJkDpW8pwXbac8g6BLHDWmI6zEYjeQFvFKnWq1O/LTykvNskd2QsHNglBW
gdQZ+DfvLZRktyipx407pQ9yAjDN3jJpJy3e9cBe9LGNhPUts337KvvhgmtdY+e8
w3DnEFjdUWmx9Ky/rYDWAVDFkoYtUTuJ55v5q+JsYT/Es0OjR9lYaF6HC6CwD8wX
zTWp5ztB9dk5mgHz28QidwSuQ2RAdf9V7xZ9RS0tUB7E+pFp9ioU+Tdji8jAhG9E
HDWpuB0IfkKFVIrVtfPwNDTkil99Bqt+cKs4pibAW6MezJ12E1UZuXkE6+hIL9OJ
0uVcS3zUJtXNryOFp0rsYPLocCUdJATpnaifoQQSlM463SSSL+PAiL1srYradtI7
lRD9X96jukTMH1NpgAjXjRK/d0koD6IQhdZp+kk9cV0b9JP5R5kAg6kLZLCQjoQX
bO5BwRzERwPcfBhlkiAT0s5EwPVAGluoNIEa72NY4T9z0BybEUj14PdGqZ8Tf7lr
F1bt1NkeT282vSAO+ksfgHK+Sz8wQAex0+wtMgDFGlSYgvoPNEci8sk96sukRp5Z
XlXwIJrMfLOpFBFsEWjfWgDSVkS15G9PwWXmM7P590xDcw/HqSo1dcHPjWbmmGI1
irIRzmBcUOkoSP3yiZQVHS6C1ueJBcTujD5yousvq7KM1yh95AJrooFYXP97s0xN
AyqlM8AwjCPTuMjs2oxsDdrM0lLeeiRTiPjdCWjfwId4FOUtrTNz8WLvsFSoaqMa
wt0SPYduem5rBohObCv/moOmah8gd8vuGBb3mmEaBFRb5xZ6gdC2ZxAA7pUrCAAL
RlmIfnhrAfgddU3ITRZI8rRI4CnjhGHphW1bNKr+SW0Id4eA6+enXtWlpKZOus8M
fisI5SqtBcICamMh1rDoBrA9ef3LPEdoWsJ5+JsPP+44ZBtUSIDkYGfp00mp7cLE
KQVHlrEtP9pYqKUdWNCkscGm0D+bR700M9Ytguvs1lKP4DYIIc1DatEfVBvQnoom
s1RQb/8sBvCCaSWlrV0D9PkDIwS1nQRdXdZ+aQDLwlH8neAE4qT8GTSVkxQbh5Mn
4LzxkfPiEOe9bOLIE0hSHrJKQvLtF/5NuNekuTQmiOlmoAFFgdvps1cY4u9PNGKw
jlHvpLxcMJJmRPEt92JgKHROnkN4B3hgplk9FWqfy6BEm+EC5vPQehUXXp22yn8k
zDpOgFZvX5TC4XhfVf2PDuiRjUkT7ldAZzoWv1W1XTYrZrpcZD2D1kN5cRE1L/U7
nTNbfIQkK/5TG4+ObtfICI0aZIR1C+j7yVi5GHHV4U9knS91IbuzVTJJoTI06Ir0
6TyNqe2GrZg2k3T0NvoiJuuseWS6ZUEQMNdoJTzkoUqIzs9UAKw5Z4TgU10fVIOg
rJevBSlZboDzCgx1Eo/Me+U1KB1DlVoynh2LfRqI+zVUiDXdMTk2LNe5tnhfccgP
tVOuGRwYTrGDHj1JwjsvFGvYD0U/Vp6WxGIux9O0cNEtm52rnbJ3LfL/7wKl8uV/
ErGmfkscu/2QbMlKp5JZMTiQyGChk+wFTAD50/7NFMFmhRzj6p2DJXwcE+GokCbo
EIUztvWsGunvKHsa31x0Y3c1nGBEaPpU1gaJ6W7o7Qy449LTx8js/NGJvCq0izLM
L3S+Yc7tczV9ZrMZo4VH7z9osOAy39gZWl/I0Hmzf+HvwzyJpcecFcZabM4NDaWk
YQ9KSPfezS9SGhIFqyhRfwywzte+LLMLGEyNh4qOvh18CYENuHSmVBnkrp7FB/Gp
juv88OWa3OaehkoWApNgJl7BnYAtTeI5IP7SgqUSW62AteZTG0ZKVFKcwMI0tOTU
t+vI+LKdcJzVFtcS4Lfm66Ar1/GFQx3aKNzWVvJk8li5zdrYEFoc78jJl9TijraJ
agB0jqlv32Askyv04yh17CYKUO8iyzcRkT3CUMPIY5wqv8JwwYnMecFnjU5gPGyB
Rq8J4jV5saZfCQaQK5P2Xh7F5LZmOw9X7EI9Olq5j7nFQ1TIp1gerk5TfTXv3nZT
P+1Bixg2HL1c7Hua/Wf9J22bQMQ2RQ7YAGIj5Xnh/cxQFK+xuYxeF0DGQ+X9K7fY
ajJ9QmA123oYqbxdh9+cGBuBmBA5yc8qy1S0zipHjmOHc6YS1wrnX64AO7j5cUTg
QRCsTza9imo675k9hBuHmhDEfzZ3i0ZangTjgM4OhHKv4Z5Ij+WDG/o2xgXfzxlE
SkJFmDfgMvGnP+zW7DUfeTA7KGy3RRHgmb6vVtV1LvdgliZfHJM85ZN9oCnlNrVV
KbWjbPiKYqzIPZHMWZ4F+N5JfzTe06mj49ODRDRNpC/gPOaeKogksFLqpqh7mMd2
f8qfyWrdLgmlM5QIEvoiU2Wduu4EfHKVARmyigAzSH2D6IrjYDYIm9JObW07+EDJ
UcjMG7sJldXVOIDLFV5yVb3YcVgsK7NUM/Ho/o/d5mMQaSFlMrhEnDof32jp92HG
xcptICezY7o1hBsqfUB2Lg4klmKdv2FxQ3dtxJ2UJu1hEcMJAkvtEO51xjbtmQsj
vHbeH79IMjcnxCUVHnjulzCzotKgnQOcWbLrolBGd12lX8U1DWXzHAkg76Wt32lh
XQP13x65l4Fi1RO80HXzTHHl2gLXAl82Vv/PAZNTUm+w+dHXbuPiiGLmW399unr6
5STFazAliVQwnXP/BRBheznO7RAUADq0sAG1gN4oaxAXqx/6fw1BTm2/TvRIAeVs
nHgttqFP1SbsQEMtMb1qBL9fRIDLoB6r8PTmTtXKWAiZLduShAv9PLDg22OrU9Uq
zuxxDjPxCzrkLeDQiGK+WIXynbiSI0Za0zX+KC3X1aGuz6ImrnyaMILoHSugfP8E
yGMa4lWA0lRDrYKlQ6bcElq1i/+yMugk+iQ10rc6n1xuu8ynPAjroD2X/4w2CYQl
wxRqshrcfxfeodz2J20rTSDy5DGA0HUsMGFpBtIIpSxRcT2pQbdarRLavKEYvAdE
uFna8wrpoEauruUC2RVV+lN6mrkjiwDxJ3wa76/vhU3HyCm0A3p7Asl/DBNUuHNf
3g+VVIAWS46UuI35Tfu8vwhDPisvvTn8XvPJApGPtQmswXrroq3JvlAG/1/c9siw
0T+intea5aZ9QVQiRC+okBHwsZkZiZXb+5haEVPYrjvsTdacuBDwbsNHbUZELnDc
0+8KK5wHRQYTuydy0YsrIx5YuIRQc9qPfTH4vOguRV2Qv6r2BqaHmLr/lWiPMGGv
n44Jzb6sQOO48m1s7bgAbPLOibsfsTSucrXHfDN6XLGGVpv8FKFyWNfVhE4NDk0c
yc1YS+xgjkiyLiST2XRFVTpTmV+LLG1ZMZBmwLbCK2eRZHm7enhUBtClRBVjYPnO
MB8RhPi+lYys1+Rj80JTrsuBQy8xHg/y+HKNH6fXdznBNsI9YaifSxQCR5JQWzm5
fL9Y1qIFKobbR7CPccAo2KInK21ZxIBuIeq8QiArfCYhK0FjfV03ZJzvKcV67h18
Sqq8Ae5Ltyt81yNLJd448fAMFtV7z79JXxJx8J+aSiIb5irZzI7dHWQQnV/nzqUY
/JDLGlUVKBLfDXkqM7xCt4qBuC4JLqRDBxjBgr9IVmCL7K9JtXFMwz4MMyAkuI8I
2+tH+3pDK4x2gNhIdFlQ1BhEG69EqfJ2DVNx08T4y9m9Sfkroa1VdSgfUyQQbzA5
CxI6d1nKqLpBk++OjDS95byqhrw2Zf9MaXzqAwqS9L2XrevxtZEr61dgLX3B6Oz2
10kyHlRo6HPIv+vyCZ5AREJi/TeyuBiHXcpianpxcjNY1cbTabLrvPauDstR3Qzh
jsfKiG2MwBy5x0CUl0Rac4Wg8LZRoRmUzjDUFKATDJajmb10+KyCNhA84urSTpj3
D73iEryMLwfIm+BYXHt9OsKU9LOED3q56qJBOXpNf3e4usgf0dJ4OC6mdpTt3fYF
L3oxPqU1A0KG9eifGVpjzUUXSqTlkQufDQ0Yweeabd05taHpM64QOmxvk5W6/FHm
K7sJgOXAIDC5SepfhnutVxIdCBmNQXkWSjepzGMPg3Zwgzm9OF6eHB+z7/xjLOv6
orEl4kDETmVo7gUfKnZUWULFxf7Mq/0cqY+P4Txut24VUIidOCv8hgcNhZonsDx8
PZ7NE4nNexJv012nWNVCnawXurWlmUMp38eIEzbkVVI46oEka57dxTE2Q+AmRRPQ
WQTsIUCXegnDa6p6OGQWAbAeJClTti8aBSH1OzVVp+F8oGzFqxvThdlgUUdxTGp4
usZeaExH3iFn7c7UximZ85KJCK7bglC2pgE8/E9sKHKlWAGO6IhZdFwDPfyoYKru
Hmcg1vVcx8DKJREohziHeuaW61L40RvW9+boWZ0NXYrftrV91+hbv+xGbPWqtw31
GCA2ESe0ETZI3kCm7DjhOwzdPO22oIqha9PLO8d+TRhQYEHt9iwjJH8q/iHvPNYr
VQI1jUcuczJSpzbvWn2ReTITEUc8r4Ru7Z/pkjeo0pwhCTaohgA860QSuFK+RsJR
zi7hs7/REHb7/HUITVq62fb+SRRtNZeOnRmj61PAT9OJDUpauFy8BillkHTLD429
pFIqAcy5xx7grOX0euoMQkIVxKuO+ddLXMMZqZShs7OORQR5kDXQHpDl16HPbtUc
tSMGXfZArDCnZzchm9gSxQXRoW1SGloMKiv/jsTIte0pSrhuUyT6z51aUW1lRScW
WJ6K0PV4NznjETppf3bozeU8CH128KQJorrQiu3//D+GpMzpj0lyJ4tjykFgnJ2Y
SPtT1tZHGxCOffkbwKFx5rY/yvJTkMATh7cCif3WhzDMK9Wbx7yvq/c94YDYY7iY
whrx6TK6MQNFe6lYx5MZ8pKG2sFFvjx5i7TT8yheVzbm+19LAMfXm5ExyKrWQ0QG
eSmP7klJWnLDy61D244YO3z+DWZSlA2cPCCuTLtbXKl9WfNzVLFse/xAYvTztOqX
u3m90u9f3qIs4NOEHFsoDaUlZI4RaKOq8v4K5O9cXfVTPeqak5C22/Fxh0RutLCf
WNe10KBQ08qVdg4IUHtRAxKoAhlVVKgGY6R+HhDUQUDDdv98C07NGFu83/vGTc95
z0OVpSfA4neTdLcIDVor131HXZe1QOhnVUcuLPsCAh15sTdW6SaUtE6MBDDydOgt
PR4Rn23iflfaMAs4l58gq+51gsrFu+24jcV7dnD+d6Sn8qgAoqRf2sgOO8cql0Os
QvoKQk5J9PcoRAtMxNafniSg8TULJ/J3/HiOh28eaPtiXTCbV1JneUC4VcOb9zjx
+kpQ9nziTsgSsxIPh9Fg1UWjeQatXtKQzm6YJB8QiFMNtt6jNg+LuZjABagccGuj
7Zhc2B5gx68qkz2DCRzgtEYwhRPINrXI7DZpUsJa3QZuPmR1+XjQjh/ANGlmgAH2
DU3gjm87ID7oUUh6RYebn8UY3g8s1V7dCHKXy4ZhPp15+Bieto3ZB1XtcnQXjbfH
pCy2mYrKwztnLbcKkry2cJMuNshEk/3q+lSLU+ULYP/Mjw7Cl0C/d/BYcXYhjljP
zH28VPD9KxHzp9GM9koY3+QuF5XrKwxXHd1RhbjyFZfFX6aYE1I7vz9mJdcKZMLU
+a8n+6VGFPSeYF5msMnTAsl23JdjeoGST2q3IIOHNoMFfxvW888N4v2qd6crMyoL
rlanpC5mnRealGcksitvT0yIuCuvVa8k/qWE6TpFgUhfgKw+PASMKHx8qEezN9Bo
PSKIgUQvHzCESZAbCq/5ZC6QbI/ArUDwJEJjyQAgBFaSxdbLLF5Hj19dYb5/rBBt
xIkIWzSGnKWQLV1xY9mzKis4tszRchsc+1j/pjALhVawnHkQ1eZGk7bHMjz3Fvb5
d3j6JbPmFLRhrgMSV5Z+K3Mu9vwHMmJUG5NxaqNmtM1m+CdOpHMKC1xqcuVFlj9U
HAfcdy06yEAiXG/z4nWKUa5otOlt2qqGKrdOlClo7oRyTn0hRDAmTTmhNcuf5sKG
2ohu47EVnCTBj46wV4AeL7WDKpAC+jhTd1RHZXODjJ7uoYfTZTqclStT8oyPDJJc
Oeeec6sIiLEN9zYbMl50ruru4Re3kc7xYCBeMmnFxHT3ET5yYynjDMLYGTaNSrv1
fORNWkPmC7cnfLafKxAAKMMkFoOiK9XdRNmGL+3TjYOUDV6Fsdy7BtdaIzjbomcg
PFKKtF+SS4r43JuiEtBpPlGkQiLaqbRoXgv0DHgfuMcqkFtkzT3RK7vcT0yT7abM
SQQIPovNvkewoiQs0dD3LJk1IrDF+5CoqKuj4odNAswViMa5hIi1/GuYs3Iq6xJU
q0wEC00fSetK6W8kT5UQL0IVsyiu+usa+seY/NDjsW0y9H8q+w9N7Glsn2Hr5Tqi
TKGK7K/3wWzQwaZDRQc8CT7OqXDoSH1b0YCxJ7cYAqwIWnGfZqxUaxGchwkiI/sU
oLlRnJ8RDwo3e1Ov3DsiE/dPanXh1D45dBZB5SpODvQXTM8Jsu7eZ/b8QYNQ3BcN
4xenjCfHcYOOQP8vQVDR+P6iY9OlD+dl8qTEgQQ17If/cgCjTLrWTOGCY4yNKlvN
wOHtEQou8aJv892tukGHWIe3Ypw1LuY+qvajHxWptvbmJ5n9x4FUH1GsHx8+TAfb
ggE8kqyYs3WKnJ/I5LXykghrk05NwkiofrnWW5hzBptSO8YG00QWyBqytlNN+glJ
2kui4jKFv7T5hFBKxjQIfsiE0DlWnervWHQDhG1HMjWFujJ8J+qyRfIrO2hATCu3
AWXIIug0RwiYN3BXWszeDT3/UwuYFnSbnN6aLarSVbfzvAaS1tqxJyNDJSKol8Nt
z1BuEWejx7rDfmMSys0zhoK4b6He8HfhIWgAQXl7drDzd2H8ZcjEaIXzsFmUMHVM
qzI7IPq58jRBqlun18D09TGssa+xlOWo11lweKYVvtGOmHFdufl7WNBRoJ1JjUbO
W15AB16fKyhGlZh+3dqTrcUHuyw5PSQ9wVrs6NAh9ZcLV2RkG86ulrXzKwv5iggt
2fybmh5pg5wITPbi2JVhtRric4rUaUl+ASFHG5252kzYlq8CgqOg5CAalCc1HAui
G9UJgZyUFDfF5kvFH4uM3oK4/yf/OLBOq9NgdMlVZhjO8mWGIX3mXZlzGC5gSb4z
hDNXYHFzEXu0dAEouQmEW5N1Hjo5Q0e61vr3xV1mHZIFgS1sYymV9kQXK6EM3cEp
A1v5eKBuxpOn+kC/31IrhYYxKKSD7qqOWChMfUg5uPMc1JahsBW/KZdZ9JrEQxpc
WJVJXJCKjjgA5HfPHjhzJgXmboIqUFB8WdMuKxLs0jczIihPpsR3thBvvQXlByYf
91bUDBK/UbStBlGJbXADadPBctQn+YhWp8A8myCT4ikqTbUOjG70qi5NQQ2D7OqB
TW4XJo7zclkJGDaXl6VYoyHWps5+vbdyz308VdYTvFNfEO45ZJVgTvZJcVpT9gbE
i5We4LRP83UPAZ96UYLda0HK+UpTsWf6Mbjxm+vMPbDj02tI61flYcPGg2uNylZm
GsZnDzFJMNs0+nvqb36zT+aO3BIeXJEmL+tXlYzwRnGZ0Kw6036qQsvVCMpe+4zt
fRT0QQaJQUrhj+fec0epypIK5L2cwUunjvlzZfRVrtn27K/GJpTYdxq3hyxuroFn
NjlIegT21IftxP8c6RTxW6lFBsuAotAyssO+0gFLK8HZ1Q++iGjX6RyiZwNQruqd
0v97Gz2ylVRRtV0ssW6sp70n2sni0d3SNVkBZ72mqUBHL7c+vwq4GrhzSrWQhnLt
IvrWl4USd0Hvx/85IzHwAMMxRQbCh7iE0UjnhQ2TzmfXmiCxsEgbioqPv5vj/lNn
9UFVPGc6eiI3j7UAyQidpdGI7on9gDQOBLfKcJXOSxdsHn77C/+mApFuySEDz14j
ekBFsINZ6VhNVXtJIEgfCSHAIezyOaY9RcvKNyf5v/As3V7Emc+PDZIdL85H30lw
23pEx2f6jaFRwp0x24g4Uc+IOunTOY+aIOVyysUOj25CxqYTNwTOH/Ks+fx8GKCP
p8VDvNPwdFzwvHQpdj/TrIRK/ovKAZKTPn8RJdOnZYZEDkBvrDA3DoN+DKAPCXS5
67SbEWjgWSYw8UoqkgpwX8j+DjRg9TyNDPbUHQkVEeHkK4PiU+llUEisDrm6Oc9b
k9iJ7hlmC/0N77p5+13egmSkOQVLZLUvE1FcEvBUOFmHDxguqFvnnIclZIWzNKgF
nF9TLRWBjkQYAFF/a4+nS41dJaj8uwMdx51Wo60f42GZSQfc+ffH5sEJbaAAScfH
mLxaXKmw7/bCkxAbgtRn8FMrLWQNMfmWDZpaBB7RNHlUWudihB4AJTLP4NjIo4Ha
ghtv+7mceVwnF9jZvSXUYKwQ8uimlyZCLVdyKHf5rEjCs+C2smg/awGQGCvHoxOi
tAnwQfNzd3grQQdZhrwTmhcwNruMdgOwQGrVb45zDq962bTMTyP4qdxJEv6hPgid
utez4WsehT/D1eg1e73lAp2eb5x4wNgtZQLJersxX5+EkYpdyZu3Qx1Lnzshb1Dv
qZLcyZPzxX5paxYcVHP29gfXMmlf/0Fmdf4wUd8peEW1/IgkK1HADvL7w47Juo48
U/Ps6SfLZkSo2JKYRkktOhbuW8Qo5H+BvPeCbvvf1CphT3WWhE1KvBPSj3/uz96I
WHj2DX+E8aRd6NzJFHa7zlWd4ROTRoJzsPWOsJq+vhMh6fSGfcocUJ23C5OMgwfE
u782I0Vase3vQwJ2icTbMDp81w3Gy0KgkvtyBE+vRvVawZDLhzqnunyhzgBLLeKR
MvE/5yz20x4tecFknVX52r3PDHLVHMVRMYawKS1aT+S+5cVPWKxigoe7bBvt7eTA
s5wfObxeQjXpDgCAvZZvMyfKAcB80CYTrN7zg2j6Y+p/yTqHcOlz8iNMxQnfhZ+9
IsYTl0KZ3X8UzgzJ7MX34esYzCK5DVKTKE8cPc3TMjuZUp7jSASpbPAeB0XqgSrL
MHRC/06HIFEa7H0R+jkn61yqxKEQZPg1nj0rRn7ogTpvUJhgbw+v5G9WhkOh2HTO
AKlpMpaxsTkrEUbjfBEhTPxXBg3TuUW+OtLkAMW2iC4RzYmX4P/Vd4QSb1E08f+c
AOt462sDAi2ffSRSSJAa/xKO0/+ILzE1MHA2TriyodjrmbpCsWsm/Ouu/TBSDt93
repZa1ARTHmLmnPk0QwyepBJh9Jm4g3XD1UONfUm2uuFsZf0+zILaGgz6NkPjha4
QmS5RFau5znJaHI/LXsR+7dR40XX+wbEtaN3WeyoMSJ3EvvUaJcc7wIlMEQf/mPB
x9sQt7nXUrkswy2zfnEus0B27gSuj9GIm/ED0lYQzMcXSDd8UjKz6loWoR8dbcnS
3aQCysWQ7TkoMGs4zFHw/EEcu/ZHe41VnEE+xmiY6nItAur8tXORB1G+rn/fFIUS
IfsFEzPGijSGHTQ5pzEm3P+ALlSFK0A54zZ05ASQplNc10zOOXL6sOg5lXbZXFTq
vHlyNvbL/5ZF5OwmMJn+jLGjKzBC2w12zTFkGmRP2whpuE6Dhm6JA+txKEsAeyLm
7g2HwdRmGEt3kqaaC5EyVAGKpf4ToJogFCYIcWdnf1FwMA+0lYduz0/qhDPudruv
EhlNqDNJtqnOnyIjbAOP901z6ZzrXvCLciMnj09XpJeA6flTjGcEGXjCAZgMwZDA
Y5DnXFpm6J5lA5WfkPV0wsEKgOnkBRaaZyEKIoioDd4FdOVqlTrP+5hOVlaeSlR0
5BNylVyMCCEFiyiE0QqXJjFdh38II90W7F2JDJy7QCbp7Qc9ZoUBwqbCQrBL0VLU
5Ga8BHP5lWOoIsc0UBOckQqkruakbG44uRb7Q1zb+vxHKn1/Z6SxjEeKJIBFX1D+
gZgo1Fz49sl367McwAOdh6A9qITJ9X4jR0lVrVgTbPQI3Glvsh2pJyEXWcfRuSxb
Jg1wBrKy3HS/uHOJkRs+X6XrD+C6os0sltoFH/n0XMQRkYAEQkM3R89amsH//sTJ
m0Vsdn97l0dT1CVcfl61Cag6P8PX7pZBWQs67RiQ0CtNY2OqYfbIC1Czdqi64RXp
6iqf36i2+FC4pSDJjLDJBdae8PlM8DbrXtP37ZfXOZ3Jot38wsPDO3NpIai0HsWo
4S98WCvrO/ngsmlIihvDjyL2TnCD3HOQmq4GUCzbBpJCW0r6zqs7KT7ACzqXUmjy
QrzglSXvqydU9tSvLxhz/01MHChh0GoxtoDfZvRGx7QFM8Z8QQava7w5GWX7fe1j
h0CvOcedJBPaD0ri3vZJ0bDlBiRJx7szvjhiV/kO6a1sjMsvyg1SfvGsVw91KBJS
FcIx0PovmgXh9grVhmezM9RzuXpAVP4YnbAWtsJoa43hXpeyuACjOuQ9PryZpHr9
3nguUW9tcLwSEZaLsaUaY1DIk1fnIFxiTHwvKcNNmW7/etc5Hn6sp2Fm+ito4xCA
hmYNnJwb2QFCIK5LVasvetk2VoShrz4x91yj3pv9BFkeLuQyEuOKlumFo+2gyKZP
gUip9anTbk8zml5FHdJ5yz/lEoNdkbSNGyK8rOqkHsasG0ixFRIck5PHZhCIJWex
cw4Zs5PHUyRAGH1xiWHDmUtNpTLnRq1FYwq3c5WvflDSi6B/k0jvpK2mXXwb6s76
TIILN83gzsYfknNHpThGZYQLLBOtHNZN9y9V859uiXT8tk3DCUdsI8jl7lNQQPuL
r7VS+jCrt5NP74xjSzpIGpHtI6RXm7aeiodaj6nEtIQEMv5RhRJyZI5CGVkV2WbZ
YccHcJatY/To3B0Ny1o/v4Dd/Ns9WNVpXipxL1FJIwI6Eha68SIFyOJaraAXmyGz
cC0cROsWC8Ic1H2bsJUIxeN31oIYxpSYVLgz1Y9ASQkOZI2vJBTdW09wthVV3D7u
lBaiTAXLm3fntIqwCZNhWK1lQw9Jc4PIN8sYt6k/t2T8pn5z4CxEk8FdRfsuzT2D
aFumsqQKMrCxq/F3X/XWSt/v1cCkYu9+4s4juBD9Giqac2F+MBXQFPcwDcLytaHI
1t5mCJa/1YlXtJGyOFTYrikco1Pf1Cy6jB5IYs3dWVO4VGfR2sH2YRLUFsmfx6gj
HqWbZdZpVB6jrlXclQCyrTYjuS81NC2nE0ZZtEqrFxnniYw62qqgAX7KJqxVPFPq
/DlTvO8A7Ylbl+U9N8kgfNbs8VTSympKnAgpw18HxDa9pNupiUQOPJChtraoWCmY
R6+Ao5oGVZq5ColMkmgqeptZ3J8PkToYzddR67vreJ+L3LKaxSM+641sEMX6dYgg
EXQNXcJovX0anZnj+5vOQCTFoi+9Nj1cRRtSbCddpMUnPtx0AsRMpQfRoutWC5zb
L4SgAck6ODhUXvI3TUbCACvd1AZ1+eh2ZnXx1C9b/Bdoa6PqNVPuu54NSaLv1/il
2tj+d1QMXg5/qyGUuFqD03s0anLOd+QZt6N5jDzYG3lb6q9PuPqwsvcRnWft097b
PTLqzaoZ/8zT8sgBH21pkjyln385wMiUw/HSXsoEXFSvdnllUEUM0QL2txUnyAuz
lb5Xv2OhFhyfhB/TmrjXigYjiX15J4p5rDWQCwRx9fvyjXXQd/POGbiR02F8GA1g
zVOlH74vBNHj12GrdoAuCQN4JSgSnu98GlZE3QvUK9tPx4rLU8adRrNSvbRoXaTU
WVuKxY6VKPWT8yClV/PEUgYxhM+3OrcPUkH5U6WKLp3jW7fvkNDXEV3XvBqAUptX
mxPggEsicLM629Qx0TvAbB5zvyyLlb5YZXwNLv4SX37dqZqWUOL7FKn6zFNnhwIx
Yvew9XAF/zI3xC6tq7u50Z7iqBXHg3MOzrVWsaTmxBe0wj+G8MJTw4PxEvzPwleN
VYeIfySZlStrJyA2ERuz0q6yJte45WGa+eVe6WU27Rlk5Z5kXAIzEbVK8F7L+yT6
mRskOquloH+gcgWP6l/Tfg==
`protect end_protected