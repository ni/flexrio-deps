`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61520 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRqFIMsr5emsPPVriiUzOHE6Mdmt4wM8IGdRVanZqj+XL
r0EgfexcE+aZ8r4Ir17I751pajoEHmULhHVJHIjRzavrAeMVnyM3r4dvpKfP3m1x
ENoxy12n+QUtcx58topsBXPt5RHtv0WUmSGlH14SEGD/TEib0dpH5IKqS2qEks0O
V9hK1PqqyWhmvRkEKWvvFGfHfWNRZueFJBg8HfFHnn3zY86TAiz+wy+ekboYk6la
Sb0vLFlDwR4cd5RdGY+GcLySVS+E7C8KTw8GNoRNKBacnVE2LSALZ1hDRp48Jy+X
LnOHqXg/tqF710TFD8kEQoZ5lElZUkD2zKUZkd6XBo9DTOxUaC9YhC3qfniwAxZ6
myOw2fsoWsKhlVk1TBAFkU8O9OU6bIQThkN6Xc5IBHjlGgIXpZ/WrFeK2RNb3plv
iOYKIB0bcdJCiooI7skBZ0vTjkOBQYispA7+FIPwyt9x14DgqjFqQMjuCgqZ/+ac
/ruIPO3/f0N8Cs01NwMEv4wT6BRKciQXt1eCZPMAZoH9KwjL1KVjT/KGaGBDZ1oU
SnPvSl6m5A0ZJ/MYkhXikNZc+uBXOWWH3mVXTJ14t5AqrvWgb0flLib8wX79r4Y6
BFjtYbzOoETqbuCLPBsmmJSjRhUvX95UqDK/8ailDESKIrEONuWWWTIgZWHPJRs4
7jz5imAva/R74hNpEFPdA1li8EhUoRDtBiudxyI656IuOevZuZgN6RmB5Sp6Gt2Z
qj/fKWgk9BJFDID/BBkl7CrOJD0GPofKKwxjt4kSeWHk2BB56iTE3T0eVtQHsrf0
nFI+5YLrK3+zqz0bJXSliPf5DWYF9O0mT8PxZWB7cyzQv1Plh4/eeBgPL4b6qbsk
eVLy5D0TyTuVV0/l1QGZHkyjmwCP+2M0rEsqaH3lhCxPtMh6FoFV3jHf7e14qVpH
hKePUOjZk7chn5CFYVLKMmG3uKoIJgY/Qk+0s0bIz3yUQACCvlwULjt0lSrpj4cg
z8ZOnOtAFsVUA6z8ik0TyRpc1zoDWHewooHJhIoyduUlP2sSEMe9ibQ2nEYiollK
iKTYNOUcIAr727BT8lPK8VNRg0kVFwhQFeYIROLqL4mbyIOHe3CpQhdFNaNya+nL
FPzijym3jQonFeZJIkfUkzz++QToZ8Lt0akxjwG5n5KR24BVvKhTsw+xkIo9jvwq
wgjeldw7S1ItOE1sHsqlBdxe1M+aSVgh+A6qC7vAY8c8TBh/mCdheFIx8stuo4Fh
RtDCfhPluVV158kAsV1RjEUCTHiGVKK8lLaeEsfqyxARGVaIK5OSi3bRYg4nOnjo
ImLRrh4CaLfrwPRzHfAdkvaydWKhuSKdcrAq9l8jCoswjlrwdKquoj67cMcFygfs
If+T2/hkeOm3LhF/qDKz5390SCGviBJe3QpbmjBKDzBrW6ENK4zxWDVDzx/3fiLY
UMFMphaZqx/0XAK/Ogm/R3T58tjoRZa+y9agb7Yxj90g1uZJ0mZvHxyDBpmz5YUO
xRriX9PLlO601t0W6THBq1VjwFAm2SBcVztwOYZuT8kun3SKuko2PWMcthBF7Q6T
jmz89vS3ZotMNFQ3gc16Xx+NCdzyHPww6q6gRPIxEnNY9fCqXTOkdzv/Nw+f955l
XSIoqMsUFR4vXmj+8IvAqkNtqfe+vOqNT5Zbo6ASs3da0k9OidC8lZ9qZmYYAj6r
PilTKz5tPIrSyYoxtrIpSBzmr42fm5DOhibMwjIXYX0QIAs7mr1q+VIVrkwe5kGL
s5v6nAyAHaB/XnppxfA5FJ31unnJbi9nNyFBPFdZL8o5T8pOAOuvf1dCB7ithr3M
ImyMeM5XbprNswRJFl8i7cyWVu3hGGSzJEhgp0iSvlxhaFxxgCnOm2ZVOcPVGQAE
RHP/Z2KuP/jKjReNIvKW1I132ukVMoiZr88Tq2vInkmSA6wN1JxdasVGUrvEVPUr
BfHD+ujOTOFLO4u7NTKuqG4HJFgXRfkFM6dhQ7wb1Qap5iphlYqpeExxn1znCSkn
l98irmWSgYY8LgCnJELm5ZNeAvJfPsajDFfPh702dUlLExjAMuc+SaYrZN8ZxKP7
LHqE087dUdB5DG4CtY9L+u2aXYRJEmVKEJt/juzwozn8wXU3yJv4e2ay4/xICJar
LdFpO0js6Id/e2dplalfOIAviSybiS1SyIe12qWLnc3R7zEeNkP0q0mkowQVCuFa
FW/qitQ78EC3ZO2CYCsbraKwWuXrla//HhD8eCm/JNpqI1xSDUW5O+/oVFB/ZTvG
+1UbtFCKbchrgepOBYoSy3dJ51f8n81SC3m4ZyqpDfH50UO5SP7bMTmLrcz5LazW
0PKS6okT54Ut7CBzLp9MW9ZjUzYsY4CQxnhaQcxO8QWRUuuvt4g/nYY0n0ZqVgae
yudAqc76vOs/3VgLIVb+0wmCXp6PY2OsgBGvyey+AvfPHlB980OlxqHUQ7n242k1
yWg9zJ2O7jloQSSJ/DHKWZgaDQAckZxG2QlmVr3ZbV3sgRtcqsgO1ndHTtkGdhYr
BBPdB9NnxUv3iXvyDctalGjWh/F1eo8MXmFzaBtPMpzfyvYeKliOF+JFBETT0D3B
4EbtjMFvRigSgtqBGTPvtoAWcqG8pF189FWAX7qQdMXNACmMFBHPQ95oMK/91mzG
VA/eln/Zel5wjZgsvRLXu5WsZHCf91ZTooQy/S1jg1lDdi1HwS7u3YM7J2hpxTJ1
4Ah6e5cvUgvJ3DuuxryKWMvUofdRFN8gzfC1cJDxWjgp5H4PyCEAcuaKaypS/cTK
gdH98MNh98ZM9tc1Ly045vrLdLwziumM5WzbO6N9n+HF5M80D/L5uqKu9Iw0bo++
yLQQ1xALc1wNMKQotzAGPud8zDChF7OTn6z6fzhWEWHi0X1HcVha2XeCMkEpl8uO
9t2UijRwNrz5YgJZjbtyD5F0v4ccTGChq70Uyk7HBMZOruWn6l27ZTPlM+Dzmmbd
1lRZk9CYwoIoPBmNcON3a0JAZisRV4FTw6Nu/7HDJ3hcsiakZf5x7nR/2KVovXxB
ETGU8IsAAznKjiV/3E/PqiIHfoDMZPgyLEqhfl6C4ZRvRC2XwF+cfi5rMiWtqBQW
mGLqgfODK6XPOQywSgqrNfrC3pp4KMraWC1fhdvxnDRswAoydn2n1Q/rukRxgf80
HkUzAM07/vZizkWsEEiYy49Y8Eo/2S9pX7WmuViHNX2I2Hksl9BMKF/eIGSp0PNE
/ekhYDaee0m/LHct8TtI3U0WRVgfAXhqZJGH0Ubk/U+tePruuRXrXGg3VOJ9qipz
ZUtYdhQVCGKJBKft2xI4dlxGg3aA413pGe8bC+xZHTqUASyl3EWVKsRnPuCVlixD
xex8Uh+buZih7Mh+wVnl5dP6GTRMyLL9p17uRBYm5B73SY26X/UTwWhprqgwB32C
hhM9aR//dGlbJBq+Hq+FxvnOrBDDof9PSZCcqJH3zPVVm9EFQDfVkdh/ane0Nh7C
YyphvFemLjfSEXRX4xMROcSB4lw4oc/uImovAEe7Gg5oMHh7l56+Cs3rWaS3lzLm
YZOZyUU6l7xz8qlK8kOONiXTp/LOxplZf9xCAerYA7iyZXhKjNI7W7AJ3vQXuKVq
OlpvZL4rThG5/bWtemLet0Rc5GpA2TIMzoX0huTWla7YcmCbQ83SxmlOHH5jIxdX
z8mYML4wKhoqf8DVLwISsWAkv3PVu/uv+O/3e6x+6Z/T17hzOpFfKI1As+gv7lIC
3DjhuGamE/up0IXdAGF/7FmaHkiusRAGWuFtdxbnpPF65cH0Itj0qg2g9sOZgi/6
pig+uv7vZoFNRi/IKEdkbg8sxLmVluEgt4qQDNH8ks7842U9affmkiDh5mDxCVnG
g9xikqG00O8d/NXjk+J/bc5nT31I4rX54GI+ssL0SjIl2MRwsO0ZfOkvLGzRevsS
stdYI3Vpz68/SFJNqa/kSGa/aUgF+JRLR3RW0BCGu3K6JBbqNKqjqcDfet2VD4dD
2h7tj1yCR8XqwZMN1+Tu+BExJ6Z7Jh1/dYqEk584MPavKvJX3PKvgTdNOUopuMB7
wjDCU6wA7heV1To4FRZO3pJe3/R2GA8JUvoRSJXSAGbK31i3oBBtWdZeu66RigkF
78p69rR3li2v6/tMBDFaqNnMdtswklEfb2tDK4sgZMrh+vpovrjMjaDwNaq+JPx4
c7OUxjrJ0pGgOtlQPJH3CnN2GNFvn1fo1OomrmY7wn5kASegkdUYS+rHkzd4b8y2
4dmNhWvb6AAVts/3fCq2rQJ0WSdU551K1Bfqjr9rKMxe7POm1yEckNfvd9RAVUHX
QirbPdpzp1reCu564mH/RfZHYzDGSVimekT20Qxk96LJERBedZEcN4JBEJ7RxGpN
IyMOCE4Fv+eUJ5n5v3KgidDrxh2I3tchXwz5+tDXt9imusuO/w3tuBALnWrvauu4
fuZqCGNLsFsDHYI5NvYronV9xmiw15zwOm84O5S+TyM0f5JWUdY8qy5yTgOPeQs7
k05kOm9mGBaEHeqcKJdoYYY7skIiXwA6j8jrCVv2HdSgK/VleTPJCPl0IWrNBdwX
xpFxVtPCbIvgUJIRsjukrobLhJwfoAEQ2cugfsBpbIcMdgmTQ2B4ugnMfxgQU9zT
+ITeVJ8C5Iq7dsI6hQh70SVEf65/jI4w7S0qQy7RV3VU+NjozTbbwGqS2P3Yk465
FpasqkuNnc25IsK/zqriC1C5h4uB6dF4EmMrHnGYHeSigvYGs4JTPH0szhhEgE3W
OAT46GySi6WUm2v5xn5Dz18cI2E8F0ZY2Xa8hrSrUQD8M8NN0ulQcJqK1LG5OBnv
uAb8sFrdEKuy+bhbabnJO9xKWoLtLBati2Bh7N7UBA0HLL/PTbskWSK1d51cEDaT
Ijz6RLQMEGR+y6gpYoOxTk96qdc7xd6/Oi8LgNHnlVdr2zSXjyE+dyfwGXmdKpMr
WBg9AedNIrP5qIjHHpV3sklq7fRk1T6tPLyxjHxsN+66qtMAJuNJmE7yqeVQukL3
oyKTLoF11F0bxJR9dGA05x13mFX4kQemQ1Rd6TBmsZNALrgmI10bdqorBkkMl+BM
VAkCzD3xPmJIvORiZD+7l9UmBFvu5Bs9YRpA14LiUo8/Ib9O6vKKvEDRTxQDNIcz
Gcwq3nhjfPYuwa5i2s7xjzR0QZUUPA8q2/VOnFowvNejFD1Yi0E2AlzdBl+JMgGw
sDaC7yGZa9RY30nIT0rBRM5UAiq1bHgLuAn+SswvsuMu/ciZlDHn0nRdeueb4BIM
uR9+8SdQjrOJMUSJZx+lm01whqzFHyPWto7Qw4+BJYVWVm5PoWJ5gGlODvLyHwwh
1r9a0v6Ze4YwyHRiP/THZk1pi141obPJ9C9jE7PLpapm1WliCDAj8gROiQVI44Ay
+kf5/7dW07+UiGsLRoeOs0SPnN5q1x85sOJyDVUzXhk2UhTzPxw7ev50O3FPSSE1
k7am9P0FDTIWM2Nfi2+hPXkvht5P9RRURZa317L8shPbVgmV8q4piEVHqacdO8mG
gMzVhwUX1DYtTI7Q8gqWZGn2k6pIUJFbReNCYzCjyvNki2T0jJgdbH/NmtTyDs9x
0bHAlYtmanyQfswgexxO8906ne4yc+dtiwu7DIqwuEjPXpEx8zIcnlalPT1QR58E
3lqZP1z6do3VAUydYXWYk2o/KqVABWXCYNASn7dc9vZcRQWbgxkGMaTX07AnOmEH
682uDibZ40e3JdGzp9U5s877D9r8VkpZpXBjirNvN/AFhHiVeFnNpwJdOJivzJgz
EX52JE6tNQlHxDW5gfoAao9j9gs5/srlJvEkwJaB0NykK3PXw4QwWfXcqEYjKc0X
EEn0JwgEWlQ47s5SD6On0EmsQsi0HUMfozlkvllSVacEDWt/fqB1XAyvEI8lU/gf
T1JwsssYtH7A40eoLGAeN9OqKXvASfXO5fRf6c4+pn8y39ZrplVnphItVPfTA+F3
5769WAPluxW/zLCmQUeTa+27ojTUxXzqS+HXotuin/QU1Nih644/ee2leKy7BoIY
rVfSayhZJTkMvQvTdGHDPmkiBhXKbLu92b8kYKbT/HiHPX4KjCBJZgYABp2Z0q1o
nKFpnjnDdD6dd/xy0VCybVGrR5i9AzPooTiEX0FIFry9KaUgF9ytO7dMA5/Ee9sx
mfLPpurGKyeKlOoxJ/91sNOfVWdt7wIPOUyLKnyUtap8f3weguH/rmyMvSCiPSq4
xsle71kAhtZi+k+vut+iCeoiDxRA97Qb8gF52+LT6+gIIVa7fM9Vuro7XIQFX632
8R0SktnagXPm0FoIX7+LtSiotVjZEqkbhf7Q025nNxEm5MIdUNLu8qktVBwc9TBP
0bcMIsKYzmf4HumoudbIPWzuQ+8YeLwBKPgQj7AalVdd8X0mtbY8cQp2K2biq9jf
bP4x8y8UH4S3TRXEsW1I0fjLFgiK4hcRLMSb00w5nkCVdwUxQQ0ewniGmMWgLlJx
NWXEs0PSZtUyr3OXLj1+WjENEEIRygVWF8gX2F+8S3JnDAr/GG1MwgUledK9In5l
tC7suDlXl1yp5gzYb7dQAqTzXpJqkNyFPtgz5EdfCtYnt5WAJ9MDktPQsGomlAMS
unYwhv5dWDmK7KO2G2pug4+ZeAzfe9Dzo2IAnSunDNzVq1OoHZiLKqOFZqUCN+R4
You0bQWm9QHE0JVuuBvQmgxVxD+bIUaFYv+te86GdGplRMnD0cXCqZKb5YJvWCRE
4sERSSNIaxHNc0oSDZUbWAhZ/m8voEMo5E9P1WDrVGYS+mErupRHTn0r8+DXe5PX
yvJKRlZ0Z7GMDp6wew1jZlauAFLQj5cp/uuAwSoLJlexdSnHSMdxMusecJCyROqY
0rcS0ehjq6sgx29bJr7Xsc3JLaxh9OuGxdi8Zu+5GjE5clVZVL25rmOyZuEaKPcM
NYJLXvvlYJq8uuger8VUe3zpmjg2mU02r1XhIiD6IT6WMWRz4S2wC8htZ5+UD1QH
RmNBs2WJTt5Dj1CzD+36HhBidprCtWHYWvTZsudSHewmUJ5OCSiQ8xCVxScJlBaU
kyaHEv76ZKaP/6V9+sj8R8QLQ9Q89JL+BzdwyXDbaxYV2YEMYCSKlybDg2Qdf/GI
DFLqzRU1pS7yzlBLWSTsowYFS1OxmbUaBwOHg7Plvtu75jQ+W3PMZegXC1a/TiOl
J8upQJL8WBreaoDuWcC5KnbSDuN6KmtOBADni1c/37nAc6mpw8GT0eSN3Z9ZRIYf
GzUlPvo8eOi4hcGS8wuGZyzhNXGOxJHRHzzteL/JNdjkExcc3B1BHohWyQH7wL4A
Nc1jh75KAZY/Ea+QbW8j3XsB1fniku8SN5wwCLq/Pc4CF3Meh6H7z7sCHYFiEVTK
WTsB3Dgt+9N99O7qj8t6Q0FshquEy0bglh0DC5oA8N14kmZ1bpdIUCISkwdGyDgJ
k7MGMBjsSjCSi4y7jI99eLhHmZdToxFcdxSzFGshe8gXCOh3xInfMw1zCkBPAk95
pymI/sD91pAqteWanByNVt7n9ww+txy7h8AJWhjepEr1xK3dccsJ/2t5M+//OQS5
gSjUYXQ4mQnyS9VO+Fky32J3BS7fFnzq/gd7PwiZ3JTuxFSiTGKMQSiO2bi+W7+D
RmTilBLCBkSGU01ZgZpbXRE0xqsZljz8X7Vfkm1R2Vm4/Jr6HoQs/etLGnU63a3t
O3WvBoeSQ+frJcmL535Co2wqXSK3e40ZaHfjpJzpKq/U32hnUAHVbSOEir6OVvEO
4f2FLf363EjGGre8AWMGk+o0XTh4Z8Sd4rLVyCNwca3A9LVkA8yTCwB3mYJCzt8X
O8BMtnD7b8ZAvL/cMIUWH1wBVIoRSDPqIn1UY91FIj8pgx085QI3z2+OxbSPAMd/
65R0Ev6cta1CywjtzkhGyVPC717n4oH6t9MHSe8cdw62aykyrTp86yKUUtvBMysF
no7UAdb2EAocXPJVsKxAUPuxqIL1gKA1mqnyyYLmD61r5zc6/mmwNT5w+XjNv2ZP
FefxKe23vsQTk40WqOAVfeT04qA1kRGokKxszgRs1GG+yIXkwzqdz85M1/PwNz4j
8b2s2X84jL2Q9yOdOX1y9DUH0P7r1ASqQIDO/ZBumGn2GzdJPvR0q4VnKAfsC3DD
k9BO62W4llf8lEpJZFyKPcIEcokJU1JNU8hVDwLu1tT9DsZ0yCRPqf9j1ficNR1O
F9IAgaSqCN9i7tPmg8UCS+/k8QkIdBiArcfsosAbLZXWJA6oRcFAH5CwtS3ThuRt
abyWE5Qx3OGBcY4Kzu9R2Fj4oRF19ZaBOrOF2YAmovF37b3G570uWLMJLhqo+2Vc
D/m74eP1BPEnp8dZmFvzHp5xEfWrEPshaGM/TthNa9ptg3Un8MphZWMTErj8QBUt
mDWWA5WxMbz2PmzWYVpBbWIb22C2bBBdCGQ/pCMBv1v38M2On08XwpKiD/AON1tg
sLbGhbCXb7Aclb7Pv1M1IveTasCld57As3gAGBfx/pd92F32aKEL/daE+LSJ/flT
3A5477/ZL9ugQ8X8r8EHSmg360lQ3aHvGX3Uv12caXWYiTopTm75xkuAaAFC+uHV
6Q9yjdctt6daWxPIpu7dzCO/PX/2gOh8J7SnbqzZpYu3dus9cvtEkAL+hzYcg4t8
2tTpcobg64jfC1OcymvMGVJV43ScTB3aEH+L9XIfO59DLIPhU1pdY8cegiw8MdRj
Vo9fa5WkhTJNCuXuNOMH0pbvpa0N7JKSNI773Px+tY9ojJiSMo9k5cePslzAwlp/
2lYM8VRybipI+71lbEjpjB8AnOPCs5lM6MkKdxGD1HmtwwKku0AVanEYFqCr8hbf
09wLnbEwWnJiYcVJznLkgaTIKS59WExKX5q4y1ulRBVYs/v7KvcKUV/U4YkUdqHS
4GV8wO2KJ2EJtVZqQXST2iBNJG2oCLipNu7Cr46+lRXziGsgRNXAkZU0QuSgB8Tg
NGS//MKB5OJCOoSGLQ2iKC4w5OaukLxk3hGN9Vn8a8X0NNhvHRsXTpKqnEhV35qW
Utrzg2QdVMThAwaetqSzkPo9B6DlilzDCJXDAMW9fO8LNvQGsWFRz5HXdllijjCQ
Ig2G99wqUczmhvCakXbRFYzvSM8ukcdoo2FKaM11yF8HR0jt5IXWhhLU1gKnlr/z
Z467t1hdvviOFgII0Rc2oZF0qk/c/0N/t3OfVa38VC0p6EvTC4sWj71lFBQcsGAC
ibP6BBb+JwNlef+VZeQfotkCYVwbz88DBbEi1Kid82ou9AdkwxJuFtZgFBodnpjz
Zw7ulcQebGkE3/2yr3XhT+2IYN0fst1YjIbDoLtxwYcC7qPx5m+XNhsOELgkvWKy
eUuQvh6pjnOtlxURpV3sZUVKTN5qYsMIO371a5TvMxWo5sby+MSoceHypz14WVVb
XzfhcnJV49UE+j+7H+JdzzB1F0+UTYV/4l1rbhOIQNGdp2I7XX4GdenIcjBD+byU
IfWGfsoMtwKNWg16q5h22VZcqXJyqEQ0B+fhXcWqWNRNd39AhciTWk820m+wEvzQ
4Y0vMTdHzyLGRR35JORcbLnEFgthdfPvexpeXOLi5ev+yxpWjf6WdcX9FFh+ixDk
tr52gYFZnytR+8g6MS4Q8RLtp9QEXXzKq4Q1Mmkr9PktgrYcge0aRI4TQkVY9zLF
QLDP7H6/CcSlcF8NPhWx7DocrVCweuDTCMDq5nCppW5Fo6fxa61plUctXBQAzaY8
+QyF5yaz2a+GqfQxleaOM04zwBsQme5Jgq9QIOnkgmbdCEF7NTemXZOtlmPtj2X1
jR7fRzzkXaRVuYHwC4L4kT/1XrnvpNPwmkWHY4Hm3TUyb7wl7cM8f2enxJ7AC1JB
ExXLiUkhOocwkJWufHV7ieMi2NXbCgnBZ23KJz7K/+dWf2+pAFDhk8YgwrZiz9Is
0dlnavFvRlhLeYnfZTF2lKCKfBYq7wbTYUBFJ3ct8tz8tlG9b0gP2zQR/sm5gazl
WU30uLYc80ZW532hGej/MqNBP0k870MiPGbvgGANocNtHZoWilcrghT5gOCczD4u
CjriB3NnseUPMAZq4eWw8wB0R0yXaCq1xujTiA9phXi27ajxl9y/S68IvmNXVlWV
Tl8cdctbYEQXguSZHCdrZkmkBAH6bNvaA+Si9Aq0LLfrgBMc7KjaRrjHlLBcoCv7
FAhwLvgiDZSeZGaMJaJvwUwOTxSyyCSiTUJoHexKvyn3Pp0RsBoPT1ovmLxjki7e
JTCaKDPmaaeVyPmPqRYG2Az7lrsbZE9Pb4mJ/q/VYxY5s/toSibJ/W4QVtkQKv11
sfexd1xOCc9gRgB0xUPOAP7845KxgaMF1cFxG/hxYh4vM8jXfg7NqfpLdxAS+38i
NslmLi2LvQwEM0CZtma+qb8FhCn6zR7WW0rdOxAGyXOxr5PQk9GAv4t/NCzRkWkh
E9xyJbZVnqpFcAjlcAoucQjRAtG2IYq86UhVZjL6LDHkYQvFtNhu8fCJNuSRuvyl
bCCEbxOX/mpCtf4bWVBdW9fqJPEDjgNbo0mS0xxZrRXj9fJxo70xAC1R6Vcpad5H
jYpt03+FNxQ7nqc1c50rnpHDr1kQRPvv1xcduVPyOxUkTDrR1BiwFpjt+x/ZpUIy
2OyfxWWXyfBxcOt88qIz9ea3Cr4WC+23Ye2lv65hW6Flskyt2Qx8CbLXXwcoqFW+
TcQD0z8WwVvBS+DHmnjHW4ao/visXFWwxgfwaoPjn28xEPa5cJ6nNp1vNPakjDSb
BdrIduCbkdQAwvqVdS+EGVZw9SdiU72P3066t4Pr9Do354qRAckNh3IkhM87a2JP
BUn/tq7JOyNp2H+e5bZKXSUkyO6L2TnFUhfLiQqDMDCyrs/LkOKUqYTD7leGtu2c
RptG5OF+771HjVyx6u2F5cIkdm5nOvvkSuMhHQrwE2P3WF4QdrrDenO6UKjUJgl4
7uFutbIXccXXt9OwMSRcmUh/fF5a/1c3cgRR3TWLiuwLkAeKWi/bJp3bEfZme0Cm
pCLJSgg8CM8/XartKeqVUz90pF6I/CxTMtzLwRZV+HHcTsUXkx65ooLt/Hyvp5BG
S2pf5lMjaMiuKTTC2VWefTQfFvxtZypjDcoNWfW9OvgedXZr90U9OcCtFh4x7o2W
Wbdr7gHL0cCJC/BoOQBpHwooByyo5QW+hvUw2J1NtisVvcwcmL40XcUcEpCmT18Z
vLN55MtxmzVekiNCQiHYXlNDpJwtCr2Be0CibG8YWCmz62bHUVE3Y6hncq9Oxxlc
ulN2NKGUtRPE3YUM/BslWiapSiKp70WPkfPKaLmRShYLFLUNG+kxwhUrTfdG7X3Q
4PXeCM/CUNIKNUAA4+ZZTZ2LzZcBtAOixNzsRAKzzZxvj5atkWAjphvR0TE7idKS
zJFphrmj3s1U/KmsA5YexqcvueiXo6i5YeYKMvhdfyI3J4cY6Z0afSuOvwDJ3zHT
R0cg0LbPtdM/YzT/x3EBRDtmekhtx6WNJtAdmdsjiwLaeJPC8QRiBVYo+9Jk6RPP
H1e1TvYjHN6478QUrhQBCrqoQtjoHBtKmUvL+6kvZ4RIsqsrvnBBl60Jq+m95y1k
wXlgY7vXcAJ4nsOPCWAScuyYTG4QfKX9kDxPFfrfjEoquPWE3+a6EBMdWbLVdBQJ
xR6SyL2Hog77PKZ2ou9J/cvOxFsF56n5JOyfAs+tTuns3qaKUShDT1hgvoa05I2l
h6HrODUPyg2mlZt8RCnXDAEnAAvlrKzeQ3x0OE+4HBCiUwVU2+hndePj3au7rgIX
UIdJvOPTsrrVPumxWbY5134buv7EtaXKP6AGP2YEM7B6Djozatj6URtqn8/3785e
uEvLPjJXaKTu1vSzp4Sz9RbP0yGCmAwhAP/YiHI8al3fzUaRRLahTQzfYb8eS4Mt
6oWLYHGfnXePTBasj0KuycZmXc1f09MHxc8eljs2slDnZ/KbvL/W74EbE8TAxq43
eeSHKmhNQTq3Uv5mJKFbC/WGWjvmeHphaOSLpHI5AVP6jLJEovonEb1F57zZCtNU
rVGWkNiBSA+3VZvUqWG/csswUrBa7ipQDSKdTeo/8X9tsIwJukcDNTPQbZi+O+ee
Qd2s9ODu5PDhHmsmLitWmAvlerA3kGaQnl+F3oBRTObY4yCFARvFxzqSFfPqfYiL
EUy0yAsXTo45wM3vsXvOmUhHgnWS07hcAYufdyobDOM+XgiFGntTwJOZ10ARCQ0b
ZUB/gVYorDkASq4VB09eNq67FGM9M0rwHuibjblvPR5Y5nAReRZs1VbomBURBT9i
LllTATi4F0PUKYU5ENY7eEBk9asWNg0IIfX1777bDfbO4vd2XIRZpxCgMLxa+Qpv
jNxWGpZvQXDcsSMxh5A3X4S3T47ITjnNzMzMp0p9nqfJUtcyg3Viz+7uTTVrBpIR
f6D8ecEnOg3VGKr7drGvMndTel9sAuQE0bQ89dSoh1Tz2R/36ldlfwwowXVkyHSd
4OKMOjMGAr1DYIt2y+EUP/0RHVU91xTJT2a3GKA5dypy4tyQyMrsUUzwYAnVG1w+
1vYevMUB83W7RTF4IzeirYdBA4jY2x9c71oA18rhHXtGp4CPK0I5b7zOq4T51nJk
lQipQ4MDXxJZNm0yaWsPWSJJwV42jTAePsAItPTbk+mpU6nbUuDCkESIcwwtOzue
VHqxJWz00KNJpkocIqITZhp8C2Li/XwEgqV6c8bOqRVWnH7s0rIhO3+NVxbY7ZDU
VOeQmz1X79dow6RcEqtBydzeqHGkkg01/8drrje15FlnRGdMegfZLLvpt48ooKE4
a4/okHr941V2/NF/vRH2vK2rdispJRbEVOlEKRFuTY7e4f1BZSrg6QLLMiXbDI4E
ZWwY9CRHuwZabt1dPGFcAjWBjuT/hoC7aW4qTUeo7r6+v5l0avRELOAB3sgvuTvt
RWMzS14GlHlTQgmqjLu4Mb/9IFWYbsciMr2779X4AwZSjkKnn9spCAh8H9A17z/7
3KS1w3WFMpjBcjxwE/QjnH1QIDZn6UOAEZZvMzIfA1OOLZGAI2AVVBIKNJjQMxSF
b3JZFBu6ozy1lae0/pxQ9AWivjVc7LBI4p+0LxXSNhi5z8oEK0Fi8U3RvhCROt89
HOXjMLVxB7i5zZczbhmyz/jn1BwOk6I45ELLedp2Oxx3NfEMDx1GcSQpKsohuYwK
a4KZe6yNAogEDQfY3vn2TGUYmvDIeJpM19p1k+KPITHhbL/4yMFOm6aL+invNKld
Wnmfo+CqaiAtDISpMyzb06QjbJq52mlKHZmkPA4D5ERQG7kSqP47QM/DOcIvd1/B
oZXfRjG6Tx5ZWnNAlbuzVQET/TUdopOMOq2wFGPlM7v1LYBc4UtfUYkjqy7p3cOx
Y9Lv+cdm9mqmevZMnN81xMRqvIM72aTUV+tcLmHWYsqNPFkCRhUAFbHk69r+4fKl
uDfnfbl9wfIAKub6CPayaLbjIlGvh0Q7w2H5QDjkKo9uoo+JWZfMBIhBHroau18Z
qxKyBvvVer/TAB5eL6cs65CPYD91TcQ4ZCyLiRjYlgBcJitFL3lhQaZ2koINwZWI
eJeV9AGaj6FLonCbPNi7FVlX54yL/JDTJ9DMIxHS4bkRDhz5SlMY1MsYp3/rUBsN
KiDGZoyx8cORkYtM20LsPXiAnBfRUqbKDCv/fT/l2e7TtHDAhw2NbaWh3RUKgdOC
Y6OqvgM82elZk0hNKTbQCQok8f2VWeKU9r/pm1uU1jBADqndSBQnC0ySqbpSzUsg
wDWGEq1ulv3J8ktmT5QxW4cILO1ZANgCCQq6xFfiEe6PPvUsS+CzILvyfijkd8jt
xj/WR4/bxji5Lneclk0gKzLSE1KY6Ua86QV30IXDzhe41c+z7ydcqWUjUqAxMDIf
7W+Ni7r25jpoBJewvPUcTFmOxs6RoZkLvil0//Ox6Al3mfqYuWT766oT3Np4fsSy
SS3g/6QOfTlarSgdie9HsnAjVNbaV3P82V/4IO7Q8hwFj2Sc6L+bWQh7NgBaXEKH
KdXqmOV3iqXJLGvdeZgL0YHMiVUnR0LirvcL1k6C2RmoggOauC0uSFsugwSrKESQ
l8UmTeGWleGgrYCEXlXHynpaUxQzNjAez0EbB05g5LldYO/+jQoF2bcCfTydFjE5
8/oMw8lVIMTPtB5DEQ4bPG3sTvxGlveMym3LlcjYpraYKRL2BD5kyNPW4ipA8Nyw
U0ZXH+DiwJn8SB8YZ3XbKXXL8ROloPDyQIvRDzETYAmHj9SKuI06l6Yas9CZJ49J
K6Fj6fw3k/O6wNEnIRA3fJDlnZT/2zNJk6Pr++j8gL++QQyNQWr413l7lECadGva
p6l9t//s0dk+yHfEw/3i4Sc7wLu9Oe8UtAUktLlEp33XWlf02CHCRnzOaS56+d/k
wAZk/Ed48ZD2OOwjqa3gsEcWusXMl038Disu3HXR5uupZ9av6hIZQRPCtkwUzLMz
bZYLnTV4fjWaE/ntboNmTvjRIlIK4rijBp+pkfjvyETL6+L2cHS/r3iemcklgiFF
v/4HCtu9/1A8Z1cg3JGeqoa9Rmvho7+6aFIJw6ld7RflbDsIbgJTSrgdHLPuuWRb
Y4qX9RMy6pr9Y+IOx6K4glNA2L7I5B4MK/Fyx8+bXir56rRfOVU+rnHobeX8myO4
yXox2XeaA9aKXVqdncTw58cQZK/kJo1y6s0igE+8Wd5j18w1SRwkEfBhqK1m3oFg
fAUpj0YaOIo1EUbYk4XR2wzmYujv8VLJLJp7zNa9Hld7YdFfKx8IyNXswyY9a5ht
ngskDNhABujaCecZpSoi0A5udmsrKuDRmChcJl2RbagZsWJ20rnl9wa2K2Z/Kib5
dXcKwRv7EqvzPDRUoOOSbOfD0ZhFGdL2ssaMl4K2xhsf1HndO8+YG74HAzz+E65j
oNSQPArHrDYQjanxF82SE2c7mQGI9o4Z2Un1xBZ3LJFyLW3+sP5USrjz6OXkNTqn
UHb8aKcvr4hwJDFwSHgL/8zbK1L7i/GcBKyjYAJenw7wcw2iY9kcXPlZJ/LRUWMB
1iUNwcbJOE2QDvlCFYo5jMbaSgbCS9xOf+pKzxVSgndevyKIzu/hqLVYCpX4za8x
pyd6IFsDVUevQ+afkw8LyXM/2cuQ2X9iRBembWT9CysawxCYWD9UMTMV1OasRqJJ
BHkWKDKxT4sFKyvzIg/4lT+yV3DvCMY010lTxwHjFqHNYHrKxGoxupv4c6sXj/Yv
37ZmvNfEKXU7NRHxKutoSX77VkBrZysz2BonD19wE9ydcF3KfAj6zQTF5pjdrgCm
Y0/VWDd0YY70SemDywos9sR4ZJ/q1yPIFp22bB4CYt+YFtFMWEe6lhPtzWgUlVR5
324RFdMlDrR8CeThasrxokcmrPUwu1KGmZ1LIJrQ4EQ6iFC/y/8Byip50om3QiG5
9+2n0inJhk+5TeNXH2DIgG8659kkXRYtIxuLyyphZmcVAgfmfykhHYXNCCZy2azv
WHajOKrW1FVc9RS7H32MGhc9ukgAQKRYgcRvwo8x37IXuNBGp0IM6dGCtKLLARDD
a7uVNghBl8T1PW+ga2AAJi6cI9U+P8wpKIePPSE5RZKgihQCXCP9vhRGlyJpQ7Oc
r9Fh7wvFjJXlvZjUHVnF9eiKWhaPW/SFItHcAdhQxLQxBBxHEuR/MR2482wI/dwM
RFz42KEeqxEhpNdYYWYgcAsIznk+ZOdFEJIbaC84WENQX/NdH4s0k5cWsLJxboC6
p0MdLGqAgVocFeCiRwlxdDFqyzS+twjjx2HxBdx6z+4nqYvUC+Mn+taJ33qsr6Hz
539M9gOrfJLEHaEm55UE38A7+cXSd4qtTmhWFI6s43q2xMtQVVbkT1AUawzKe/Hg
LEh0EexoDatDn8ExH27vZ3wFCirt6/tYXMYJKYT+ewutTuTVtweRMhUbbI+DvbuV
rtGDz4yyxQVBIj253ML/odNjLY2Scc5MPG7rQ5cv5rcTV+j8AOpf8LJEeTwB8kEl
v/AT08H7J+Fjg5FvPzF//3E8Y/umS6apyENYxt9BHx/ilo8zY6JiG0C43Kdnzfce
Qtr2+jtsvXA3VkX4AetFr3JDUzMIAHqKeSkr9DJZpLtzIJrqdPgLOXOKpx/KKpem
meySOolh+wydIQdJtRhd1DFy+4mkpuW8MpUOvnUZn56+ceOI9Rlb09WxsPc1ISkP
ZXWeqqCMbJjTaC2JK0B4Nx7Utq1zXmSTt9Mm/3YZ6cAOAx9OaebyBjM5TgkmRKS+
s4xBHlXrqK8OYARcwVZkMIRnUdt0I+DfALIl7G+aD1bK3oVG3ccF0jRtbI9tkUDl
svskhh4zLO6zS3pmTxDSKV7Zdo5ts1qbTBZNdHr+RH3J64xm/q2p8PhX2lmywAXo
MDcQAWLvWpueTfMRLNw2qEua5pi4hzqMCMKf1I6+ScLwrS0PFYoRtVUqBfEAD8yG
1tItV1FU0Jq45KK2MtyJO7sczPcTax0FIMuiMrewdYosWZwXWd11s1CBb4gAOkFA
TqE2Y7a2NXvraJj29HQMzQpMfYJbE5b1M8Fdhfez7O61vkgIi+XvKmaAe9Ym9vVl
SXCMmU/MP4GXEfNTkaNvCZ/8EEcbVr3LRsfAGd4yJCm3r4gmxtoBaBsVO2tc93Pb
vpI9wJ0NAkYPvk6kVJGdnvlYsdlIB8lapD16K+DVdBljTZF6hC/Vk2cwVmgxhBVJ
C/FU3syLLcO3JS9V+rMC5gV9p+CQSg7CkPEoXFWNkvTYxcYRO6EM6qog6fzI4qGW
FPvHuC+ZfmGJkhYzjJJORQoafFTucgp+xQnVfUkiovP/kKlX2q8Sdo/GbGUQTNxu
qR078qOgkhT3FeVYU4yKcQ0GWpzLzTGHbyctGDrPLEl4p2RF6VX0TGtnNuQCUj6e
r4VXpzTBO/s4wwbGCmO6FyfxiTuAImZZ08tOrDIxS3ATM7FC2vSgwp7XRzH4j1M6
eysIrfEAMB3XGzuniBGYqbksCMgxXPx1Q+y1j48mH6L0UFS4ko/0wXgDrRgTMWbz
VQ79D70MM+LIvf70aZZ7ufy3WWIgCFyJSLTsCLYH4ARwVEtYuo9bNjNZ1DA7Xfxa
2oCI00MT3j0Zqnj6gMOZjJqmWJ7/650i8o6B8J0+6IpDPdo2wffseWRH6I/quA3x
LLuMcmDWB4i8uInLLL8RTIiYKJurwXMnQ4NVeEH2yU8rGc2/sa8ZwM0MekJG7RQy
3W1GR4gcPU0+ot42PRxWcPIdayZekGl8l+nR/1VIc/kEsayl/mBqVBdS/lNIzYKa
SZNjQcnKpAdQpgz6EsXNF8R/vqxmNfs4HGsnV/tYvlvjzKJu7K8UhQq+MdhZScaw
Q3VZMsgiqRhcA9uisOveZ/1nUQCP/1eFtOrgEdK6P//E//6RxgXL/xjVPqJgZw+n
c5hZD7SHoVca/JGueZdUPArTFUqSqeCssEkoO/Yn0Qw0Kj/y0G2N66CCJMhQHnI7
+W9aVSjMhENZlOY2GY0wkHmfe+BNbxe0ueTnZoQ3YeRki4E0iFqOfAA29/ITva0G
8dqbpudAHaPN1OzxQb6ufbgS6T5zAc70fzT8InpmlHQMBHdqN7/LQHk4alhL6r1C
tJsyOej5DBS1+Q4WL1AhevwrDg/4Y3VGnNTA01X7FvCj2wqmYhv6YFAV7wVhMscw
Yv6HNSs/2gYLBTRDLTa1G3kJ1n/51cM9Htldh/lrnTd47wSZickNRS9XahC/94tR
H7Kw/pvdTJ9ZszlFCDywcU/adEtG07MreK/rGYD8LzruzRhIXHCWNB94z7N3KG6C
Gugxn2Fnbpx5PmqUlY3bU78PqmOjOyqM+u2N+XYZDs9Y1+y6FIWQKkZg1FeObkGs
F4SuYHPjWRqd0NQX2Lzljb2GMzf5XTJshWAWYMczyxSpTG9/3tFpBALKgHKUcsgf
at+xGt5/T0hJUSf/Ju0CuGsARCohRciQCAXsck8tT88V9zgTqXYhh1n1AKiKe/5/
5itGCnBnn3fWkKi+3c/7cWOfOwy/QSK7cgYntvDowawH4vlN2yrYo17imojryuXI
VCDXuwqEK5L0NvQJxrco2usrt7CFJzGMcn9GPkY9H/yIamySzsuCUeJaqPP7gWLv
czNrc4yjpAWi5myea0y/82dsP8KZyXZbn+nJcfCXa0l6JEb0PPKuTEmUD7iEQjlF
2CkZ2pnhEMAVyz9Dpx60gqB8bPaALa3RTc2na3rLPRZB6qvTgK2MbNnxWrWUG/T0
ZeEJH3jic2zlJxjo4cOkbmgWEkzpDEIaZOjDxXQBRtZ5U8vZjoTPzHPTLthSpizE
oL1qY5eWuur9OJz8K/qdSwMboZ7Zj5prFdxre+H8WSO8lvQZkcOmhmcy8pkPIbGx
QBSOMDTE+U7DhA8nAuChfl3pYo8YnFxHraPku5l0rKSr7V100tIAGw/+RzNXMrMk
4T4fFHMW5KlZId9/p/NmUq60rAc32m3hHTzU6sds44Y2YpEH1uxlITDUogrmwWV+
zw91LTMFCX13b+5LNVrM30Xi4r4kGB2Csi2mcg8O9sMMlVe/ifIaHlX5SmyD9SmH
bcEZfzx7VwrIFaxcmekYJgfwmbPgcs5dPCEyHXLx3+raH/85C3OT7FijUh9wCDIE
qOk/AyZInoHqXFlGsfn456za/4hcj5rEUbCtsyVQmx8EWIocYjzDsfFeACUHmMEH
rNK44MWobH0bgHk8h2L/hT6U4DH5zeAZ9DUruQO7tJv6FN9q8zB5soHH/oWCU05m
rwmk+kuX7VmjieXf7htH9gG1xg/C6Npr7rpZ0mPaMGndi+q7D2oK6Z41YUe8E5d1
c3ieWkSPXFLX0pWVIdgjBE7zaNoOAiYuQ0PEnlFwX7ECz3Vz3y9QZP3mG/U2KX8Z
PO6gBWjxTo7DcU8yInWkmmrQ7LWo1OmkaQv+tUTCKa29PPL5IE+nowkXkwYzHfbC
QouQqpHvnD+OWJhhKI5RJPGKfIkkwZg+QRdPUXHuuIgk1WvacsKOnyOYTgs5zlz0
+4CDbdd87lsQG0T+ckGDvbuPBW6JZabAWQlOecuRZiUpdD5fUbHaJzCFpZzb+5Zd
WdWvP4TiyU22l7f/3Si6bQFObJN/zlX8v2OVuwb43YyEUOqMQcyhwIbBgPzev8Tl
OyduTu6dJivwhA2dAqq2IYjxak53LD3R7b/iTZ+KmqkIEYxi/m8ZhQzvVrPDGy14
KR8irBMMH6/Dbit/X0zjSRI/+0q2SiEfTiDDHsVFBsyC5FdrOILY3JfxfTNYEJPd
eh3sYJXirUzA5fhw7Vox1xyfohRqc6TnuEyKznQqVBrGxJNgZUKN04SjOGrRRJzI
D4tLmLttjyukDhDA5H48tt+Q+aNDjQqryMythsb1a1sZdt8egbUwdmIuH+4fA+63
p2VvavqiCauXffZEjC0gt3mbcy40Xo30kuQzrG+kSvYKCTd9RVB42h5r1Hrw+wPb
BedNMFQp+51BSNHT4JXLpn1yxZZ0CO+x2LqnNTPR3LBxCe/08/a+NaD902X8d80b
LeVgBij4FyNiQeE/gF2ANx3CnXzBDyIJHcjgfY2nqmdZ0SSGOq2AgtJeOFq99KPK
BTEFAJw/LPLBw4MRBV2mRs53FJkXh45TU0hLsg7axDX5f7iiZKq0AkjJrn9R0Poj
t6GnN2ow3CBLb2lV0uf96PaRjHXZ7xJgAvQIEZJipFFwPDvWrwo8W+1NXOTvHr/Q
POHRM3gIwkVVtO+Se0+9diTSgxGat63Aa5ynmBdWtw35Zp8/00VY7nniW76rUt1v
LO0O4+HLZdBpsUpdgv1V10tLyBaVZtyOvowOvrBkjR3DS7+ktR9/eVC3N0CVxlJg
T3xr3pRy2bqVm//T0ouoQi5e1GlnQc9y4ZCcq218gEf1p8tEhUGgTYwjSeOaty+u
7Xfvj+CD89oTbAn1wfo6/ziZZZnWE8KZfRBXqIYmDKXacZ7lptstjoDM9+QCHonz
QKgSqDR8n6nJQLxCI4r0wKAylXTXULQQ0FV0bN013Zr9eAGbo5WbB1bD/p8/irra
iB+pEfaU9TXrrspWulFMcueIhIaGH4RVOkzXKiK6PyOG6sg2Oljxuast7m86XMaw
+U8RdZL8r46lQZQEf0UhgRA9zHn5k9TwZB6VAEeu3yDGziJcL7zUnngxaSyx8zpa
ttRNMr5Bn+Qq5H1sKHNgckXgC22BOJcx6Nsjy9UoaB9xc85YaE384xb+QG2Utj8D
KRy3e8lxsG3prmQqoisiEIyvdJXUjwRK9cdY1OA6aDpcZY5j18pl5De1sFcdmrEx
Ay61CWuSjaa0g7EWV+otp4hrhNpYbLwAu614eL+cff0e+br70jdsfaTm8sE5itgf
vASTU4TRzSRuprqtt+XJetu/BXxNHlxPFhhKkbhtD9D4f4tfQ9B778F4a7dGPnzh
SoMUYIZcwj6GQKsrb/g8Q+m0mD6L9Ri1h1S9ACTpdTn8jcI2Dj6tTpu0kzXTaKTg
Uvwd702JbOMPB6/CtMeR4pspk905KoRx2AQ6/0laTOoRR3flFbcHs4QUng8Q0RNj
InxwTX6qOOcwmiw25qAbzxyHDOk7g/HrgTGj/tUMNbrHOL8Gg3H5FCOI2/sbzzFu
34YCRFcuWd5Dc9z9gpC3taQy54h5tvn/olT9k7UnzLsoslCJ6WQhqD/JHf92EmNr
j5dGZ6ZYi4eQtbSQkIJVlLLMQzxfVeC/yvsxyBRy1t93k3TEbzJkJ6Ut7SDPIjHO
9WjGxIoVycrVL6xfTJhU25PozoifOyyPErVGNSbDY3nOBZal2bSltnhvGlqoA2CC
3QUm4urg5kRIOioZFevTaN+NOE1Lgk0CsiGxWkh+132DWeUinGGGgvGFiIhN/I1X
Tb0Zuv2/7sUe2D64mMdFEbL1JJy33beuYkBUnLsCgtf0g3vXFX4cczINx00GviuJ
PgcHkTBIouZyAtdpBVn/Z37gwzqYk9rDZiNMqnBEdmyLA6QHiqWcNukTp3KKwa4k
479Ccx4V+IRJZ69SxxzR/zOR3DeY0sO8ldiNhrRPzgc+c7Nk+qnR6Fts1mP4adyW
XZiGJDh3jsd9CgR5+7C9ykL0OIVR0h4t7+lkUnno1/5vEPyVYATqZ7exL+JgJgFK
ZIKDWhM6McaPlFRCFslXSAPANMBYsXgVHHX0Tu7LC/E5Smrtv0K+ZsIhsob3PtE/
Q29sNaeUUsRtC0q90eiJ1bjRatNcxUHq5zdIy+/XPKDlVnrt8EvnXvlIIPpHptiq
NJBDWiTF4cLBbjWht7bwFQnCJ9osppRk9H9sNWD7g97FbpexlOBFU69j1IOH8R5P
iCP3YDNM24nP/Omgjk5dH97WLhCjoBP5tqUfh7haErUyKb51/EIkI8uRttaLQOdD
NZD58kQ3b4yMg+dZmJ2NZ4XZr52M6Dqkr5auWu09Cqfv/1FR66aTDszq+6kl0h4+
68OUDIBZuNidtAjd5RGyAGsiDQTN9DOQWkYvIYlSecgq0a9Rm+76hzFhyZ3I6xhG
0hoc9aGeJB1nURgWHCRgadGa4QCgIbOaWtAyEiA6u5+4ZqUWhihFu1rrfN71FBb7
0hq1XUmzGs+OCSucrn23OlGwnvaQglUHfGIyzBhlare9+hpv34zDdGEpjAaJ0YrN
3xFZudS1S3Q5KFmkP9zBWwH7o1cJlO4ZYa76R1YOMerAaEkiCKexCuS2lkzK9wkc
zdL4KmhWi6K3c+aQGRSr77N/7uNPmYRRy61ugfVfOrBKnbN2R300QOgxheQG++Jb
W/6kwhl2IHi21PTCdx9813ugtit3On//OdkVFzzO+CKCtfM/f8FvET/wkQmTm0cA
3n02TPYEwum9UOfyiRRe30gRDUnrtaT1MLJPFHQqh4X7KjrMeHSemysBhpZS3vOn
Vacu5XmY5whzeClNxgJCAaGpNMcF0bkyBMPhfI61bHH8XIyFdnWzOHqYc+c9Quzh
5po4ZPbUHm3lG25vCqK/lmX4KTWWCmM4tQLPfMwN3L3MBj8+uM0dEwHIdtZu/pDv
2/3BVTOXK3XXLfvRGmGAvKTjV6RbVAprPCyQpl5rxwjDYp+B96ZEu8m1IjnmQi+w
p1GkzdTZmylCbwCV8bXiV9+yfVh5qW+qgobZA4TzSk9HW4vI7w7gqEt4nUX0LVqo
BtAtT6rnC/yL8rC3RumUDLqWmyuRof91EBaTwlORg72U77/HpV25kPSDEcwZ7Eqv
DX/Muyc8tLtg5lWkJF/QpMSbyWuVXT06A6Ud4bkOIHbOyLkysDlCqsMKIfu4+OpQ
nkeq36qIOPpxGlrDRSaRMjvIyjJVGl+eQv3iLKMX5p8ft41n9bKQzVSQ8p3UENmU
KmlJggdjL+Jve6PY3PUsk0Exqa+Ru2uEQFhZvpWnNIi2QgIAosZrNKON8Ao62b2J
dNFLcMh9rI7IyCCr9+my6ZVdMsG8VVOcC9ZpuvlSm9TdzDpREVChPYSalVx+3wWZ
y7pE2vpLAWPsXQvPtDzlx1lb5jLtzb/TW1WM1jTjrdRlVcFDRvEK7KimJi3C1rtv
Y1gE2dy+9gK3Hudsyb1/ZOm/W86UYbgyaXQ6nrbP/uFSzo/VpizGp7jEjpq0A+c2
dZi1eT8vWBfTZINReBl+EcHXJlLghPjI9gUeBxG7VdYpvtoYqvNzXrYw640uhOLR
Bl3IQMg42uMA6+I9zYLH16J3P0sCInwpRQtA0dB/7EWYYZrJ+Grw6AncpAEKHZy3
zBQoMWKkbgRE8OfxzhcKdEqCWEM8oa1bQNMXP7NJjQaD/33d4rVDFhHNS6FdUN1w
g6QVQVuhb5v9QlSCnqF8bTz2fMbgcV+SNtahc67hqEfRtYfl5RV4CpRsmyaufWk3
zvrHXHGT3MXt8QQJ1mxIrarXVkJyDDbdJV9nSferl4uQ9M37AjDlSPGDdwGTrVa2
6mdLCQEl6FO+XCcLH0zxlLRVRDO32lwpdI9v7+mb6YHB8gsTxr28dHE2efuWqn8G
CCC06JvumEJdeXvt0kjiF6CH8StA96V3U3z+kwKeQu2gmL2LxT8RxWxjnq6T1sjN
xSp8wEhiAnpNNhfDyseWdTxtWaQKz3T99K2l6Q7jMvJjQlBfORQ+dmjpw1LNxEbg
N0AZwmwJcU3h4Ln12gzn7pNcvP/CzheMEHhw/SyaEjVFX9euT5R9mw8leYppp7z6
9x0pOHrAk7HNuLnGFnAA7motz1MH7WrNc+PB3tpyLnOfNRP9pVXTOh3LVBvUo1tE
dohsdT4mr/lKc5UqLFHqjtUUxqk3nBjSAgTygqdyZYZU4CVO1u/NkVWwNPnuYHMO
6p6uGpNlDfWp28PQGze9sCit1tr6gLQUDun+FlJJ85iYQaMFwzy8HzBJ7ioqZxtf
t9P2melo43BDHgdnJDx+qC5qJId4nxNbXCipWZYankvsh2YLqw5PXkl4CwkTk9nl
qhrHRBiX7t/n73pyMa8Uq5QIKoLcseZuXqC2apd6tWbWpf3s0nBw1Ypo69P145gp
9x+LbYd2YjUDE+sS9iSTB2wbqTdR3NuT3cVNmZzHNMtuQcFIUdPyWHtVLKWWm7fS
gwphM5bmuwJwPIWvCEUuU6+7NIp9IgymqwwXqoDN9inlA4+3dbBpzW6aGogRngFg
AIy4vzwnqH+PXt6J1ic7IpiEyw3+Yc/O+MoCTaDO2BAyFfJWDfHY/jyn96SkgE0S
2H985R5uiHMFKsML7WqKuWqOcHsuuJPMLmzUGSf0zeevIhDx9nnbTPbRBig9sDy/
vRSjnPmMEK8IVyCRWf7FGsvkv0QH5AupNuNZ62WJK7P/KweMRvuWz4nzY+8cLsuM
Yjmbkq6X3JVp6EUrgxb+dEMc/6YhqbGiAiZcn/GKiH4q5dkrJhuAjiy2fZheVIk8
+3y6BV5L+dsoXh1Yp57rA+0R8hK12nwLFPKpoP3HlL4fiZOZsdFHpthcpu9dVL69
elKkzoeN/i9fgyyyOwMezP0zmUTkS96i2we2P7acp6dv8KDcUro6+ktIg750FWkP
2Q8j+GGsVqbqrTx/FYBnlmhml2dNtHqeor8cbRhXT43Ye/iU5F2aUNw8DpUzL2Vn
m8l40tkV2F5fb0dakKj2nEXEyhkQyi0ax2r9raQ+KXyIEPxLRvR/oV3Jn7HocHLM
1ufBiKei4YEhL86E9fshhOMHMS8kk5+4KAmmMtVDXdB5WXCuLIfi2ApI4v9florl
43cb98vXGCvWASqKo8ZhSLV9gx0t5NPkJyGdqaN2fvNXU1khH7lhVJYaEgDp8mm+
gICS98OkKA1TGLKsMmPUvIdWVJNAbeBhjMiyCmtFvl0qgx5SoDqfsoAtO4b+AEih
162w/xR7Eecz2YHU5lljePBxKBwKScpsRf3L8BNAdQU9TBra0PueXAbPrG8xPNN2
Gv6a8OORxEIHjQlsRityTfGYBSka5KWI7o2tIv2aVDCbwMHRUuUX5uLYpAUTNKDo
8W3IYEwfq9wjH4RnbeBoo8aMup2pbL+1CQl0rdIZ1U1aWYpM6RvjZIN/8/nJL12H
/AqobNDpPEY1jetqFrckUKlOgoBwhuoDccB1VvU/yjy/Owgt3YjXdSoJlsWOkOVt
ugP2p1EmVmpkEKfj12NKVa4HqvxXWxVq7hIP4SotvS48qW4HCLsSO/vd7emgSr5J
CfizzkMntm0kA3AF1Mh2SkajXk6hg83bH8IbE6YNJZtnpAIQzVcdYJL/QkzpGUxq
agObpcMlwVq0sNTg/1Mdu4z1ihi3Ruk5TDJC5mf6BwKzwX/mdhqzjsIt96uIu4gV
s1rC6nH5qL4Nl5rxLCi9JYpYfa8F0qvUx2KW5atiJymO0PZoHwv8QD2dmLWhORw8
aUUu3wDj/nU5iWXZIwOUXYY7udK7fpZYUqDJu22hZZWmNO4rMM00CGjgRJ5ASsa4
URh4sNoCfNIAkv4GUAFBuzB4Xhvy2DL7Xc1tZF2KHc2BtjjDy7/z4Q8rNAKU/vR2
QRB3Y9u4TL2IzYCYCyvAqG4GveqkP83+e+mQDi0JSCaqSGxl9azG7zYpf99oqcXC
BeXToEYorZPo6Nr1U2cjG7IexbeC4Ttyjph4S1F9HsPBUFq8f6jzhyutG3RFhFdZ
Gsug6U6IpqF339fUfI/OYqiX4S/f20q3zIj+0VggYhPgMgRvLyXZMpVOtfYrZs66
6vfwMXXW8k+dKUMT82GXQrtjnx1Uwqtr2880auoy+aO7dx4TILuQrnP45kyKk4Ty
Tpeqcl33Nn6Pf2vNQPK/xRA5KEyfOkLABJmr8cYsHfvntkIS0rCKbsiPeqq8t4E9
RUdTEWBO+Y7mhi+oUaz94bjwmxlUvtrqAtWv/ifM48b9hINOLazEGYZLpjbhkYsC
4z7Gd3cgZbwG7oRBb5lXc/+ABonGRyQ0vdqi8uDjFsYtGpPACf9RNhQ+Vhm2oCmX
IgbcWYz7YFvLaeCmCc1TCTQP6W11dgHHavA1EjNnFpBWdjkLuVB/hzyNY/UVpIbg
1ctUYXGFMFBfkYzmRcSCrzyf+Lx68ZwY91cC9G9RpHxD4BBl623oPJOmz4Cgx8Yr
85Qz6gdYOaYUXrgQxQ3+PzyIdLCxmJ3pC3NzPA3Fq8BMIbbyJ+Pb4Mw3ZtJ9Gk+t
U8R0Yu6DXq4XnDgDKHl9n4mMAnzM64S1i0g9TlbSssyVqpNAZOJ9ABPdPWj332Vh
xn4yimBsd0dn1CfFSn3lPo8mfId7uDPR+dM1Fh6i2Qov62opB9vKbwu2QND8bhhQ
LbhDyhvAq7hwnXXh/1BREvZDzsUfO7/RTqsGePVMAgfMkWsIb7/nIfJRQo4rhvCF
+4Jy33k5EOtr1HsFAI+gzsrJN/WOusYNdArpXBNZFClHnUJz4H4Dt5y0O+SlW8wN
G8g7P8NzSOiVs6Wj8DVNNKSwT8Qt3O2ZngrcB8V/Lz2FiotvBdyDEH3f5mESVRA3
CgXfp+6Fdy6E8mV4V0GIsGcLZJXYurTpGV6B9SxXA2iIFjXvfBxUim/VTXWhFDgx
XBkChuCEu7vls3CYsEBH5NMcKCYaLEKCq3OUAcgzdsmVKtVlGEYFp7xh4ZwoA0KF
zXR9O21ESi9qfPKBREJfAU9fFqDtoJ21toHWDxWsa4V8RPN+6uIepBD4hIkknUcm
PLX7Kqy0N2yi+oKb+9Ig9w/5hYzXT9gYHscqXzQiarwmvz5EAvB3HjEdEpaBTDDN
svL0vRT9k22hTpKC+0jWhKPY40CEwLHpr87TDuHze6hC49TYdWymuDE6CTCukgk6
M3gm9+qOZYMm4U/Q5HyaFDHvs9v8M6a+rpXfI5eKFXI91w7IBrTmUyrNz6/wXnVw
fPn5hExVDzXEW42Z3dILhfnXxiV8dk21z/o5YblKT3gxO3KN6udG96qc4p8Yd1GN
D7ZfTfM3+3jajlqhsFLr2Za5m71F8KFpOLbKvyvAS2fnGu1iY5y+LHrBLmwBXh7m
RTYBicuKnMdtPBSa4UV9KVQBQczj8eK1gTI5jT/atWDhHE0tVKZCT4VSBjZoT3Sb
uUOK2cHiinTpYk0xy5BdlpyFUBZlQBAPhGJ/s+xasCdV3pZ2xveM6p9ukrch6EBY
03pXswCR/VAlvZM3mMxcCBmbKD5b7kQGQqgxxr8muFHF7u+j0DjuMe5S+/Iq07bO
P2XfztcGO5tHpdzcHnZNFsnHtyiS6zilNxyLKhv6WB4by5INhSyCNfnjvjR6egR1
2ShQRHsE/rk1Uspq6bpSV+eug2wMuqdNGQY1f/iOcIBZOtLJf0vIdsbdb2SuRayo
DrlgMM/wYH+clq+tTMYc53wKJs2vKFXYfQLUWIlj7OnidPcz2jrhgFa5+E1Spjm3
h3nSK1fXnIuxQ2rSMKCNhy7nABjqm0CqmK1gUiXzh5PmUsATdH25Jl9StlpOMB4F
Nvc7VdnAF0CrkCh4zoO1VjlhVJa3GUVuyn3tHHJOB1BBM75eeOo/nXtEe1Ru03OO
8s3LNYDFVwVRTaNPfEZ8jRyEZQIRVkvHGb9J+oS/QHcpFuoXbtvLUPM+TM6KQ5G+
I8YpXavlfJO5OVH10i1ZZsbGdH+d0hS12Myt3tUt05JwipvxtPrx+Ac2MXqK96Q5
ef3G5ko1QyGL9SlP9oKyPJlpVWj+6c/pCjWEreS5WbQNr02VRK29moauD3Iib0RY
gAiIY0akfv+alXoxE9nybUw0lpCdxDAnnfpYPwvSm9+kGTeRDkHr+9ywo30bJgHA
wsgq9ZvALaKmPtT5NJXkuHJ1KGzU8V6j1gUiWIYkai0P/YtZN98lvwv8iXk7FO7s
jTDx66dj6CQl8YUYb9ta3WnOw4uHGdBNxvs+k+LMXy8x+oXUPszgXPI23puE2SrE
36FJ0hMV9uaRiZh3u9e9TA9ER+JFp1WKGHI9tuyX/IBIDbZwfw//JZYfIeLoTGX8
rlla3L/WP35FVBAdUGIhGCL2MX/LXJZP7fhzDZ+N+PG791J9guZpuQQE0POfAmK2
7zvE9LQFu2hkp4zW7PyXdV1QeAJYXs2+6tKT7dyROfJlqdZA65dT2zExn1a2xrWJ
baOxHKO+UPOsktj1wvmjp6jZc/RrYYT26F1OkpmBn1G7gTWVpi/d9RNQfeIVWdf0
f0ynlslDovP3b6xIo1t1xAv1KUzkTgUt6t90Lh80mUHPPKOCZyF6TiwJt+fXJ06B
KD4k3jmQ0eHLcL8Zh0ZXwXYYElM1Mr9BD1y3Pxx/T7JpxWIThtZj7dul37w8JNPE
Vv4Y/13m/5MCVOYkUIdLhluzLdwzgwu+wcl5hnY/Q4YH154mz3169fToXiIzGPzC
aH6gf5+7rO42fND26aVBrwyYNPrV6LEKGafxCQB2u8qSWhCvTT5VNFUKerKid1hm
kVlhAt3kiFngq4bnE8xKfV0vKgwMEcsA919t7vftg1+zFHP+SibBFO/DQKI9nSz7
xbCArdaVVYQgAU52OYD/JOPQqQBBf7D9asGKEYpKvyvhoQrrqPX8cnSku4j0klA3
ySYgyJBO3Pkm+QauFQ+wXEgVKFCXaHInwKRCI6Miu04JnIfKB8La4xcKbNXsjwoM
fASZ3Dg1a+266iGbSAAv2MY9+XLroYllm4j7n4wCNShGmey6UZ0b+BTdoEossRo+
cqZp9U6WbjStJd3JXhf6mkZBXZnWgHRoe4Qt/HKSFs9TRKwBJB6AS6EM+mdpnfei
oUfUll0UWMtaVSX0/WmVN+FmFQbeKJba+hbEl9vBgkLv7m6ieHj5Jt8uDEuNOnET
/JKGaJkvgKDqO7nHvODi1hNoUVoIe8CkeNsTIixtMEsU9CLtNhKtchxLArWowUoj
DyymniKAUlVxjZkZ8XSpPqxrVrZSSyZWhkdNhXBYXrkaFmrwTOYMPU6Zhtm3rR8B
8XrVprGbwj95fCTibR4asDaco0YPv3Mb+SrlfsLwjTdYpTepMNx2jysFpiMObMXf
sU/K5rcMLHuKbEpHBbnU2++Vy1dLh/acGf3YVTz6NI7KebjG5FuWgxkaiweSaAqn
W4MkX0zSXWG3Owiv9h3M6whTzjDrSxPQB2t3DFI/QGE+OqMVjKNaMbFQtI/QIAyG
POX+dbLh+ycIgPL6z5B1ujLmDedVw+qIsYGp0THZtwz+TXgq6ykdM7dXOrz3DEur
QhgofViZvMzH4rUuCxF6uBx+PeR4ujcQ3DCp6r0JXrshDd6r1CYJSQUyKJNJzdXh
BXcTBeo/BFNey0vtO/B9X10amw/geUJCE207E5Gh8+WlNZejivUBNmB1PTwYtBo1
MCPfjnRrZKIROwgRqmjoNJpeTtggbPG55scFZIctQEc59Ql8010rKwaTh8YG3PTn
3lzTjDqmsw1NzzGBXOY7i0yIa6+VTh3TzrC8uJXWAG6VMavyj6jRehKUOPyYqdQx
GvH2ibBjxHLITF7xzmvCgR9xG6Apj+u83ct1qW9E/UpMNsq5k7WbgpFhSfb5+XYh
07DF5+wOamzPJ4rj4UjH2cU4D0ZZh19mqUzYiKIWfzH0p5EU9BZ6WWD7YXPEVDAq
6Qgqhs79Zg0Aiyg4P427zXcgYeAUJjjL3zHGNxWU9IKUmsd+N/GjoiUjyN/pXOpw
CzRUVRxy5pvb9KjfLvqcmoUWRRrujEr5nxkJw4+SSNV/qUawuFMfpF5rcONrXBAT
Q3HDggg1aAAm6LXxwIptGrEyAo/CKZ5FiaK4ajOnrxSscJNIFDqIYq6DoyUZR3gi
QcDz1LIqZPQFZvZUI37fauXBc8PFizfjmRNeqaaDutkqXxEXJIjRuIHWQG02lIpz
xOBOpS3ZSFhqy3eHxUY2d1RfAay/vGLL10B9jI303QcZewYFeFFr4ecIGuuoTmJA
N5SouXy4F54FbRtYgDVqaTQHAYCUy1VjVcLeNh38z3fExHig9o+kMPsNFz3zqXCF
CRdy19fQyI28D/VMEYfA5q2DsntNTD/6uIwt8Yl4Pmo99c/0XdURrNP8IMlVNaRH
Re/nEY5IQIHAr+JDKBk37hBhulGDwmFA8ey8ClQp/cB7Gep0pDoyhPb42r3Bm3uk
c4iiCw/+zLPogjBpAQR4tUmoPdq1n65YN6+yMQGCcGPptuObWHw6HOcWVrTP6K+x
oqgY2mwWO08Spl5iDKAXuAkAmQNkko2rnftN/783di6Ob2ZcP4SbnrCALrLsD9Dp
FKdJGLWh7BW6uRFXsQg4El5yb8nWjfq4+sMOX5tJmC9VJsuWrLl9Ht44KVghScbw
2IpF3bxqvYma02rO+Wu1TDaoMJwU8v5o/ou1gNPnvel+5LzM4HD0Ja4MgObcMDcp
BxjJgWKtjLZjoKOQGNb84h7mIPUJXlJYhERjj6IJV7lQPr5Ox6fxS8Rh20CxEqTy
D7P68iMHXcztydBp+MUrMKyK8vz5Al9riIbFQQw3CKtIgJuOkK11GPc76dA57OS4
y1eHzvAd5Tms4NbKWam/ED5HuXx7JpNQzCCZQ8Km7jMC6rN3R/2+hXEjp5dP/0sl
ijebMg9za9AiurAF4awoBWQkprew9J/hopARa2k84b08GxkV/MWP0YuTk9r6R7rp
GhZ0gNhmcALpAAaLKpQScSA7D6WBuFeJMLOsDht3EuILYq+1IykuFf96nvzN/sG+
X2QKPTkjcJ+lOxWaQ3HuyxYL4X0quRwP1fRjKwU643fMmeFM3RsvwkB6KZrga2f0
rJFjBGe9CECtRA9MchdI8zUCLSObLJNRZrXqOqTfksSQtdtC9U3aeo3rz6MBFfME
5YZoYij0ZE67B5ITnwcUu7tsFdFfpmcJ6gVPVAWURPTgN4fu1qP7sUnsKk1Ceihf
8L1TQ6zo4KaxGynaGgeKOd/YEANojXK2m3/n7L0f0jsiz1LEKGMI6zubcxgZqGAf
fCCU53mwsxUxBj+TLG3O9n6pUAoR97WPbgLH3IqSiwuFBRBTCTejhGmtYGiL6UmZ
OSVYXpG5a51IP8L4tw0npd7DKdD87zcpTEWS/VnXlqwAexyif9+sfoFSMzlymOb+
/SpNOxfQUnpXBBDg1SxWt4cPx1x+f9k8j6qq/bBZxtZoH4TQeHvcLjhdRCqPpCl2
hf3xwMcX8IguOKfahrUwmSXPkkNmeJjJPxr2h+u41MVP5mhxAbTW8l0wRwSs0pAx
AVGvrH5doE+MJ/oooIRkQKYr76/Vt2KYars9vCZcgNBvVoTaLtOdR59Ytifn1z9J
ViSy5BSs/GDyaFPB6vU3WIWVkB0WlbgowTe2lK5Rn8wLCMYJdvMKyP1CKrB0ZOcE
XH8A0X2gbu8uAw8EsTVp1hzYF8pHd+M4Xtu5fgQWZ4uDQQz+JNXTmB2wzMVAW3/O
z6sPHV/d6aSOTGAnU3I85CCagAizplBVN8akWzXhk83bK+27mOQd+KVvO+wmiezt
y1Tq/VRRpFcGAXUhFTbbPjAakrTaA73NhCbC25YLyFLteyFDtrAHZg5MW0y5wQCH
VlqcL2z3F2GY8n9CbzzIUD1cTKlsI4xjN9U9KesnOiPDZRbBfKNdsDeVn91UQVz8
/R/3hPRwisjIkSUlHougrdrjXFIVDz834gmAt4aDtuS8UERgOqDSmdqEGTS2G/mH
hctleemz4NIbIpo6wATBYkIDVVhGevdkQ49czVgMaGpXmX5uYwBz7/f+0GlZT+Q4
fHwoGUFjEZdRbYxG9nTNiiPaIrXVGZ3IzRzwxDUeLxpAuJf30vLq0NSmm9F8i7Nt
ENSLnz0BOfWv18HlQEXWD3jUaOUk3yn9TtcS3KIXBnAx9jqEXcERmslUyCkO/0UQ
+GUKaTC2kCSRgVZ0NBOMShIVKA+JYeCzInkuwHOEQxJDwhcTDqJ5NhFhjL7T3vnk
Hg+JCIIoSgr5/LEoNmQehp7dHoS0JvBGmcyCzDNOKIu9JxgFijHOfBHzUpkSwbCZ
Hrr1uPDYtsFulOrP/8u7YuY7sTOn59tzGaH1Pb/p2hguy30hhSYzjOTLn1+pPKCh
kC+b9aXi81K7IRLdbmKkrlJSHcSz00K5ft/7+/CWNx3F5NIf3/XBdH1JFxnpWWBl
wQB2jkOYpGruDuaFwALPeRHcg/MNMnhxDEuCMQ8X5jtR+p8yeRuHHuOa/PBriLA+
FM46HsMlmOANg0Q+f4U7+d++CPOiYNTlpOmeX0tZv4AGgyHaIBhjYMEuU2KSIf/f
+oiw8/lDVnd+kG6OatL7zG5SjiJWlSIe+7ZbRM+CvRRM3sFh8dmP/kTnsQ51XaDt
LiTMqt2RU2pzkmn61YXVnthhk+pCLL9rgN0/N0evyzYy3PG5h9JP2HE47cPVgX+G
mppNfF/RnY2FQWmAJJJKgxLDngXl6xTzebO9RhfTGkx5ZPn/62E8Mnj42VUWMHOD
e9wo0q02IC0LFPfiqtjc4CvnYMMEBKm/vDdaHLQ5KqM9i+Ls4r+W+/Dldc6updIq
rFdu2HdxNMrs65ELAs74qIswdFCYM6a8Js2z0igzO05RKgSDT5KId7RUwGfnvsIn
5qaXRXXmf0iGOWI3/8iqyxe9Z8Sc/bWys0y+8JW7JmcVAMxmwt4CMGXiS/HlsoyF
Xhcte3tJyohF+QaRwX8/HbJpBvsaDaacueJUx0+9k8+D+70hbH3YUjCYoK9D7kce
MBivFCVRbZYWQ9/cOUk2om/NX3ImTQ8mAd3eWpmd3IU1Gk0e38Qb4BoYQHmW++kz
caxxXeW8/IaRSZmoeYFhD6tl7p5mh27cKa8Ec3X2GaDn7j7uIR49L4m5/jAbSHDl
xzq6nPdzsq5X/KWi8lziWBn2T1L7xtYtAx/goO0KmOVHHkPEKGrLaBjO2tocy6hI
pf7PFIumWW+ZURSlw928VA0cN2kb42LRuqpkhj0V3Y2P+GQxLywU6EZ7SN4hz9vF
MUoeD3ghzseA184kEmB6f1vKD83aqTfbSmlKefFKvVkAO/XGSgdgE6ZeESesztDo
wPyCJnIr9lsMOxfHiROqWw39LogxtnQhHoxnlEQbfllbQwIeIunVWW5stPtuGJKn
MFhl+Ve+9iHNJPPYwuoaW2Ju5RmCNSJ/wJoZvWwKoWMHOi3krqj5uO1lrVde5gaO
LLGsoioqiKErKPuwI3MNzyMOxsz/yu+hAFwoj9+hJAcxgRLszM7jWWrR1D53N9aI
mtOkxHXvAXYjiYO3UhSwOn1vJT8Px06vn13ngcr5q8Wz5XmbN0Mdmav9FJ5RJwW6
NyM0JLcVlJmPoX3nWSx2i09U20tbJZCs2bN1Fg2K+FPJI4jt4kYXLK9HcgYjbXN8
A0sE1fDgOxnGRjqQB8yYqp3G3a5UpBdv5eGGlWRjgZ/ykvfMC8fYTSA0T6PW3wOS
G+swf6kfumVqwY4TZtxhQOiJLqs+HAS/w92cYYEIVkQPbc9ZfOEXlZ+BjG8bNDjN
0/bfxLFCs7DHDUDFH4LDFvhv2XZHcmh7zmmCH9vwVu8mjCEQSH2tWzkwUXqV0H7k
n3l8xZnb/NceltWQAUjUAaMTb/eThfgt1k49he3f++87DF36Z6zOc9KRvdWxbh1X
saEphCtUbLFAa26Haohqz+OvHvtB5K62mZzmSrDUPnRbwmFMkm69ASaHydGbwQMG
Edf+Az9FNKG4yjbYM0ZXSMDtdTy0QIDgPNCBpYnOJmxuvpXWUrAvOkboEsF/caVR
/wiih9cqQmJ09WG+Irofi52x9ChCjPQ3ZrHztHQ05fvuQ1cpBJEiSJgk1LsUZhlb
0mbob6faob/BIP8xG/RgFtUpZsJIdK6qJ5oviPXl7hd9pSQMaN0/uD8xbadcAo0h
rMEZfVHfPFQIAQF34+LVB/+8YWJOP42a+6au2tnHtCR2wgPNA0H9jmgHLEf1fKVb
9dXlj/w7k3hFfvWy7/u5/Tqs67xwjDgPbnbwZddRiBUxXS/xExKyi4ivMXjzbFxj
aHNWIYMfl8bv+xG4kFiLUNd651cNewtxEfTz5GZb4Cm9kTdyaOXWZpGViKOs1wwD
a3wNitUB/uiqXAONaPee9+bT/Qb9xuX9Aj7fuP+f6LlRi2fH1PFBFCGunDa/zDCu
Zwd2HBPbRgaW4OB8NKModDYeMMheGHNwLB8xSLiyCk/gfKczOHjPfFVJD/w7zFEV
MYdhOveBzQ8t3e/06y+9DFjzA9/nmdbmXtvdU6eJ2dwYFauJ4eULbaCuk9kSx2c+
VhndZJQ9tlMoXRrVVpgJxsBmSAMERnNXbI2P4wZ83jLXIO2yRMgdsEkLlANVnMq5
ppLN1f38pM/20t0mIP7XUtqdDgG6wdiQc8uTcUHHQhy8Mv2YitnwV82w6x8DCAuT
6RwHufxfklcnp7/7XppWH6emivSD0EvtrCABG2QaOOOzuWa3TB2YbH+yoMtRKMUS
nAF7oOvFACOwlI/7Xf6vBRfqFEEzrEDize/82XpyFJNQxwP40g0GDbjlzsn2/Lrc
zBbaarUfRGUz4J3NswQd/gCbcDdcP2Itf8/Ti+TdI0MwRF4KlDpJoRM0+M3UZVze
WSafMGMl+PqYAD3bTU0xIbhtGTgStbCwpWad8sMsjaIvq1OkFCSZvmfiEY95Yjht
CK/CK6QgYLVDcMt0QbzRDaJYxgvVLmHZP+PuWONAM7D09f40obcS6XcJzWEMCxnq
O24nohWF3iIyQeo2eeBHQ3TGpmUxQTl8d//POPGK5uSp8bvwH3U/G+XXaanIRO7b
FfPwQJEjg4nBNZJ3zAcoYm86GSqL00MFoU3/aFJ7IS6eSFfIuhLchj+m+O84pBNe
J7mc2NEa5EcvaAstYI1VYR2aGCDMtbMmBIr/d4gd3/yLcNYxFYQmJjKtJ4rsQR4s
7ebCuG6t7YqEvWFDK0t6Ank2j57wMaQ5A3W/6DLwMzt0OM/gv6nTgTwhC5mVdgFe
VfJzmxeTAUmQmZm1e3mRwv2rr5JaGD4an7Q+LCv142Uz97HINpsthrsZWyzQeZHi
r/pOnMH9kzGDiGk9RfyqzLjVtg7Ra1FIMdoQojl8budlpEmoS5tbGEJv6dQ446q8
Nr3zb+jniGaCTiMem8WhoqbCSmwo9txZxwUdr4tIcq9Fsa+lzqPflgZJokoBdTL/
uIly8fOEb7NccwzO29PqLOmYHk27gQb5rSPm95Jir4vXiLMrratOQc9tEZZ6LqXu
iF/s/uly9GwROa/jKIz81lHxYRXe+HPTodlMrFJ3crvDXJdjqO5SbOWBoF76hn5r
aZ8RIRWgq9BA+sqZRD9tJBb30o4XVBBUN7Yyu4CMmC6BaQBg3VSRi7VmH2vdvWyu
ShTwEJLtzj8XhoDRlk5S7ZYUvdwLVDWemwrg8fTRJ+Do+sT6I4pDzHATpr/TCzRe
3u6bSDllQUN0+/zbJbMZjpalfDOIV8anR3n8CWpMXGwH+vX5oAMAN7p9fFpeofq/
akEFTRAlcSiBNMH23eJM9XKMMCTNq/gjq+78byXL0JgGaG2D9C8vpiK9xmcJgkwL
bICueeG14krvHx4OjZYGPKPMl668/forSgoRi0oAtBRXEN3WDhpD+kioF4CpS6e4
23nDNn1819qerflnlIpWVyBsgG7c5njPqWo/92ArUWmZoAoB/oakK9BKX0z0iQS7
mMNXtlXM7Qp4gouV+PhSk5YoFGbbPcBRQxjbIrNC1r791cQGxnELEJEQzrsqBSGY
mTmRJAofg0s3aaHUtTKBYUYnJJpKXphGKa06q623tTfaSdFUga7w4MGzoKBZuaYO
JfC0aNR5XLxYEZcz0bq198ogN26wNjgeMoXkIRQ7oEMxJxSWCd9knb+WaJ3U4iGQ
2NzhT8dEBh6roPLOmw0UMKZ4J2zSvAOFjNjY3yYjIiXgzhZLwieHH6oDNW3Dw9vZ
gXUzWSP+R95RQ0OSyF4QPAXVrTi4GaVM65id2CMJjKYE8dk0jcND+1jDmonKtw1E
CBvFecyp8eyZF0WmKjYDCrqlkTt4NpqkMn+IwzJMz+UC4GK15O0akDG7uYlNDeS1
diAolJGQrPvA8X3irIL1FWT7UIDQad2NqCYykvYBX8xawGs/3qr4Kw1t6ViWooR/
l+sL1zNU+xGsNO32VZm+sdpeMfb1MHy8q7nh6XfKAYebSPjb6n1Z3LWdk26wKb/O
KyFicatYR45zdQ9jRftkjKK+jJIEfDrRcZAPp4YP5y8cRyanj7eQisUUJpdulUaf
50tcWybQx/y00qwDLq5v1XPAN3QTMbNWDtsId46a8DEL/jfUEa79yhBSk2a7gnJF
I9/afH0DyhrOfmaGqboFaBhp2tHUHabWJQNT6xUxjVVmSuVey9+Uo5qR+RD8dooA
uEpH4H6fYfGCYLKeUtikwOtmcraVBHXANbH03cJF1by9QaMqYdZDEnTbabpbqJdI
bUQdDthacjIogjoL3uGzKU05CCYvUNJjsLqYwoq4XzZ0M9rmGnAJ7022FObJfZYY
RNPa0kNAxXkZ89KwXoBvVl1NlrkjxWo4CybjuHJJnp3VYS7BCTjn8LGSCLR1/1dm
XXuOg7Bgu1kpOJOHfsuLyC2uH0QQIJt/yIQeY1YGInj+2KEkFTr8Ykf2ztjg8EhW
KtaIw3ZLr2l4CNvtQr5dBPZkRyVexdrFgWZSxDMcLA06393uToS/sjbAIwTXnqDG
InwzDmR4JL6L1R0NW8tsUClksKrLIoumxKzK6buoBQ4jRSxRNMLhH1s56FRBzY0u
bs6gqvs5W4+UK/DYe8bwV5kJHjFQYUMtig3Cd+7RbwL6+9N2FLtHGsc8iozwsTpS
zJlgsgrQ3sTbbVvSLFSg2j82inH0dYozN47CxbSxlI5rujuikieGnfqmm/aJgtFv
RPzgbrV6OyaSa/FkTfgrALQMLLRKrwmZ0Avjyc9yrjSCopHJLANULimBQwGJhFuF
Q1tadgsATuhy2w5Q8LuhSY2AFmcnwZTwb1UVH0fzPX8/nqPi9agW/D9Rbs3PHMnk
1XfR6rdtxCEVNH5oAdQQAgeRgWXXBrcUIgAcOrqERnlJoEopvXer83lqTGTBAg19
8tKQqez0fKt7RhBA5wJ+WPHftN/w0Nfpz+OMjcmRPilpr+JK1xGr2tmu92ItpGCy
XZ5/bGphaqAwYVsvvD0Tdaw7SpKwjH6h2JlHNjyHZiRDS9LMALoXd8x4A+bBZBs9
LY09EX67Dfd9ih9rfJeho5TRUb6fxjtFYD/0ghOTXuOuZM9dSzN9UxEXD4YfBN1v
Ck7C29Ny53iG/VkaXLEbK5pij8xRpIDMRVkwU1j30A9xmVI//+kVDBmvLv5zmGmB
SfXy+8PKTNobrcrmesAHl25Dyg+4F2GoRRwxtiMPgSQElnxCFea2pLsl/LvnM1vn
+WJ3+Ba90LArnmz96FkVgsOEzMFJH2MfYzZHlcWCtuijcudIDHElhSt10OxcYkoS
ReyJ8twHIJwCVyD8MUqmNm4yALkRie1t0Bwl3N8CYQZMtxc/PekaKih+lq1J7Ks4
7SG4YdHVTC4Y2J+CSpa5i3+u4hBe8lO5joz+e1SVBkFNnGX9OLcmK0A6pezY5/Fz
pYuMiQDj6Pl5TVk1Nqn2wD8wiHPANIPlGvFh4jx0m898a0wyaoX5RlzMMmyG93IX
Y/6Eue7aj1QyBAMxPpqo4Bc2KtpHGpdVSa4YkhmVZVzpszMRMQ33KN0QoCPXUZ7W
VWVmusDcrxs4JawDvqxulZThGJeyDyTup7wqrVuNAGr1vhYUeFszzTU8t2Na3L2H
1M3P7VkjLxG1crGeDJEC+mGQhhEF0/uzzXPZlcort18+WYa8x97ZavaeeVJFotsZ
GM0Ld5aHHXVybro0gxjL47IBfVBSzlEz1J4NKRVohEEHk6PeXuquRKosaFctRlim
QK955eJOqistSobzO42ZezMiZzGUxPVCuVNC4aEg2uQo5GYKEcGjTsWutiZ2o/m8
8MOl2+gfybxiUmH5uifFjgF6DkrN5e0y73pKjEf+129EsnD+Bhi8xM7jVxRTPb3V
dGV+OwEi012QVGmxPrdPN/KOrHbhn31NWU/FL+b0IduMHj9NoDF5LdiQAsMH3dNQ
8EpGxG3qycsd4P+k2cdHvgRqdPQuSeF6SDaCcwtRxtTU+KaN4aBnNiLnXgoWX9p+
OJ0eU2ttDW1RqngfWictP9TRHDLQZKF6MKxrOkHf4mw4rFIFyp0jNNLq2eFC4vxy
ua46NiSw/Vd9Ur+l8ZQRmyBttpS+TWpm4LjIn8QcTA3iU9dFQ384qB4ZDHNuiceu
fX2S0TC4QHFkNBuFGAYEMRnOobuLLu5kRq/DiNVvx4ABrptmAZtz8AduKJRxosws
iz7PX08gpIt0AzlnCzW1CQUPy/AV1+pWUFWETCL+BbN8cp1RI7eiRDSPIHYpGmvC
DZhL15ZycP943pPvEB9sdXninY9vK+E/+hdw62lPNNpexjwgyQoNkjaVjVIMEqN8
0aiqtnHpSPW4VOD4+X0LLn/Xyvix4acyfeJL63jD0AILg1TV+XZ2BU8pv2ZXO5Mn
TAr6DV/jRKCyibJ4s0r0rMZa4rNBTaSKWCRiYP8kydQY812c0GqOwqRdikN43cEh
p0i5d3YbuucSL1/ofrVifv1tLTdweRoHvJOuCvF+94aZH+BohkOR43mQtBEq9iF0
cNy6hC6pmGK93ACfbg/siW3haGqCq08MNeAK+Y9Zhcb95ADfQFP4HX9nQtHIVq+e
DaxOs3WIt5+iScqwla+C7eK8GlPw2wyh5LUZs4yWQAdsEeND9RkRpvGa5vVPhpUW
ByoSmP2Au/WoWOXxcUTNQ3mVHx2psql5AVLqJVX1XHskC9V1tdLwz1JYMjtMfxXZ
ngmz5IjF6xvv/SXCujzOHOK238y9m35Ik4evIbQPLGEFl8EGDGgtIgzjHsQ8eKwI
bQcPrJvqDTyR/6Bc1xC/8dpS1x2MH7pdOL7+SFsTg5P+KKU+qoq7OAZ0uZSolx/F
aRZfKFD41eSkzCxnmUaJhUDN06X1mPaWLnFSqCdAj1qAOOZtiJaxNEE2vtI0fpUV
79o+o1tAXyAN2wg/yWLCahbXgUYsGtXGiNIOLPVIqlN0IeVRtpak2ws2jQQ+g9JU
b3pH+bQyP0+gy8nhrvEXBdemC6wIFOzNPvc1PsBZhHD8BoNohNrEGEjlt8Gp0lWJ
fWx2CbMS+j0MSUhylaHmEsUNPQtWtRNHwICNCDC0IPGikw+iyJD7EdISH0daH9kw
mI+jaEUGEehw7aLbQPauO4M3Trkwy2vlAXLQl7Hzni06iwk8FjADRgaElwoBxf3N
FEGyMhBfx/I9P2Ripapz4exZN0Ak5jjtHcdKFRaCUruXyk3fALeGX6kWtelhTJ4M
2oCRn4nvoG1RX8/cYM4yJXjmIE0rJUCGLx103CKRnP0ISxwTA4TowuM9Ht5RBl1Z
h0kI8BKcaCehg2vSoRLyzCqLkf4ZETgk+8K/Y3z3hZS0JUJ94JKdB5wnKqlLU57l
tLElHLvIDQeQa0FA/koJJAorJNs8veM31NHe6Lo43AyOgeytFTk3wSsyVMjSyMd1
GzTHQD059ZgfQk8vSZknxF8tkf4IFnB0gTgH87XV0ByzIswaDu9+MmYSVRvWozWt
ti55amdzvinvC+JmjME/AXbUWNkntFiMNZ73BNa28Wy0chuvWAThYhpidafQ9scN
n4R67Dzzdm8+ntvS0ohKkXNGcczPgMbNAdfxtCdrm+C7r0pTHuTEwPtGwmsNL+Hc
LxCo5+cmQvId9bmWqXsjsLYSnTH4png142uRfHo0/A779HZQT3QkKb4KLsbYGhTJ
W5T5/2UmXr1oiL1DUn5T8Dah7zomXlk4k5CxTlXw65l0j8LjMDtJLpzeYRFCE80s
x6zQiAthN62JPGmTDLyumTy3FcSsK2D+9+q1QthEqetL9X/THJMGGrNdKxVPblZu
iI1wT83VfaGEHFBTzExpS7VtRRcZObDfiDlfu9ZfHK4dx628Sn4kOjYF++0JfOOx
kHaNHXYcvuxnGjXueNPqdHl2oYIf9WQxf8QOu/u03swqdd4bKL/9vjwKMZRT4CYR
A3on914IScwaWMFZdhm5FzOiTROz22TR40qqZobveOqqGuawREuRarjgGZIEwfDe
7fJyARa0gK5U/bhy/61prHvtOrf/D2m6AmM/28d+q/IWYc/NYsJsxG77STA3XbqP
hoRChWI9OCxrry8ynr5zLhJieGJDVZRGCcscCMwBQgp3p+my0jFf+IpF/VN3QiWy
fCNrI69K6Vfm2RRncMeWMqBLyKZu0tUzqesI0zDmZjo/lvfmPMK6aPb16GZeNItG
YdBb3yFQZcLI9iAWJpWbl0UvpjCSbeHRXcsYjEqM+6SLJ2vnc5/F+SbvDZv8Gb4J
7svKwBzK3ndKKTeM6Vm5KgcCAnU14kJ1QBn9q4qjXu+xSsBTxfX+T7hRP1Vw8th+
TAcTKSrfsRc6NmW1GohcOdBqSEEoPrTG6XUCW0UybAqHoXxvylOaBIiPE+jXJD4b
JxC1DlsaXCo8tkFWAhCieHSjbYp5CzbLiRXR4lVj7tbEoUC3CyajwgpyZffRcIF0
TlfEIyYc7o55ggnE70Bxo9MhVjPWkeD0+iH5lgkwbJSuqc6TFMr0k5ggMLu/m7AT
f+y714B0DHf0eGuguVY6sY21mNjwtra7aHkuXKDeOf31keEr3k8PdnzMunkk0y6+
h6/NgFxRgd0kg9Ou9DCKPbrzfNbpqJQ0NBilwsUOMRhvp68CT03m3J9XBKFWoHUJ
Tt2AIjBKTkZ0UiXo0Uxs7+oalSo3Iv6kznj/K/NhA8wcrBAkh0g442NfsojME6qy
gBToHG4JHZLj5tB10eu7AHKn76kDV1Gqk7drrB+euoobI/EyYm7OyBdKwFNUjSLN
LTpgfYfV1buhDotrhPFg+HP0C13POaLIXsHnOmTAyDSPvvYfmw5N02RSHsXpisOa
0wKM34gRUTDcA8F75460RZxGxD61JyzNNakQrmtbO4bj7gcbT0NSpRWZncgLHgdI
Y/mwcCN9ZrvFGtV8zkfz/W5RUdu5vacKy1B2nPeeavAaaN8IYZT6PY2pO5WR68Ys
Z0a0cGsgOx4td5K+lQqIRyMC0387VNL2GrKRI/W/Uavrk5WXdk6qqKdCIrr+tt1s
fR2ysoJl1RjAuhj1ThH78w1gol3Yk2QuoNwt6QsgYCFoOHLWFIKAylF9neSFHDIX
CuKF3LwE12il0yV92lf6YC5kyUpCOtqmKACSSP+cReVF7Ss+0XFi6GNNONZf7SLj
bSQe6IEBHvpSx8BdQH5eAlr2Iq3Vto281HLhz9m/V3KfdMyxWMvYbiBAgy10Tmqa
+PNTSQXK/S3pWC6LfeRIrWu2eXQrIe5op60bfM/+b7+1iBeJ7pOzd5fabyVibw1N
jFqJjsV9lDfmHSn8jF2ZgIS+Dq3+kBWw6HCYnfQHrNBfNgphptgWtjzEZy6+5jss
zpaFf6YgjOUiaVHzjzZRlBZFVA1RGKEf2ZCw9RXQ+jqGVdVHGWcRM8I+WCwdZGP5
SGNmD5g1RBM4laDIP41+c09rwBDniKLtTeuZFnLlAZ00utGdN3N6ZEz8+DueKfDa
jOP5RWlMlsbcTGRAU7Mp+tiHsn8w6z08d7f6c4mdUlpjnwW+UzFrJNM+tzMTt4BU
zMJxYroBi6H3FwaStIY+HQP2oBc+heU//ocfTnM1G5bY/gRBbLCFYBX5qfSygfkd
n7tdRaNQIMnBCZuD7cfiP7jKeuX43zdwsddL2aSSsstF0Gcx1L6X+stb21u6PR7d
0EMjUPcoPqZiA8+IR0dKMVtlyJya3N7VQjPL9CPNAtZW+JdwHBAIknocXBgK5g3T
Tr33GP9SenqLuZTEB2q44WFOmZtE1c/yFCsj9oyGYweDnVpPTrj+vCarwTseaaIa
L2tOZmLYfuANMBJSuLqJl4gVrobipaICoyll5T9l9usqdARYHl7beiqIEK8ISvrj
1vKyMUJwZGfxAqp2Rou/bZ8gb1RpMHtq/vvFE/+l+lfy/qUWPN5AYTcj2Jb13cjn
rybK+cxTLLEDXk36Ialb2DdjISVi4WE1XMwOv96yKRnLSKYE5XiyXQqMHvS9krhJ
YT0zXa7fwD4D5FMpZZSKTFc5FHE4fvFT50uKRV8ib1K47xGI2YrP8k+rosXiZTid
h+auQ/Y/0QdKUs2lDM+PTAPKBX3G9bBHJX/eeZl/Hb9f4kWiz6Equ8ohBYDE2Rc3
+phaG/T1mtBNWbbKt0Aa6Qt7/LQnxNCAXexeRZw8+x5iE5NSHyfcF0QTPBGEJQ7r
9fzE0uoz4VRgv2eY9Y/y5L7a3XbspInVMUQ/MfLlhOIb682VcXVeliqXqu4i/gzC
ebD178bFC7PsoSQCSJmvPJ8DqqVK3Fsp9eLNaWmo2eXoKTRrzqL3QUpeg/rhEhqm
d+5gPngw7GtCRT4pYV9JkAOneXlEDbvKrLbRzE6FHCFFdOMoU5jnLl+bwoHNifpi
vFwB8rmMhF7DqSc6ZwCvS+PIiBhwVa3CpeYM77P2kHxhfyu7CXOP5IyLOOLaTZCu
jIVy3A6r/KtLE52M/5L6XgUsPZLyrqJyDBbsiA/9nd1KJA5jGxuIk0ibixU/KQNY
+0AAyDKE4XuZgCzeZd2kboiTcCuI8AT+8Rg74dieWDVtXkonuuOZzcxDqceYSsNg
ZZtFVJeIc/6n7WtMXHVGCfhYGL1396SuDpHScsj2bMV4PNrsvvUALHYRZ6uRT54Q
/ev4rhoTlFw9bITHVMcAu9zvv2bqW5qHHNiIrnWb+TT+8ZP/YUwAKnCssp5VMYhH
k/Ekjgy4MppfZZXWqdwT/Zissx5IqTm7RFIKvzNsS79jkLXfHxRbbl6lIduwayb3
DbgPjf2Qh0S+m6HV7ytJjgRFjFc6i1qDXfejtxxLDrAoVfJYyb6FQ3ky3rO3Cdbh
8sqY2wNnkvsrI1z/Lqjypp3WbhKOEy4TkuJd6ZsEUAasfDiT5v1EUgyraEJO9A9G
drnxs1X8H1mv9wSwFiXTZ5MeCXorxRpnZTH8p/8f7lrM24/7AJzumcZsGE7FAVhn
FusDOktYyhelWWDuwdBAXhzSL2DdD4KQuVGSwyVPQ2U5NlS28j79yJNOCoERgsoz
1FdTfCarXDhHDZAAqZoa4xLFSvl8X/ipq/a+HQ1obeHC6/tXjawRjX2mlTKlR/Ej
3VYGI/a4rT4YBbGPtT0es8cvfAQfHiktbl/DjapXajNKb/apA8422TUcQTjN2fSy
Z7BuANebk9Dzl/oVB1hK5AtSoOM+xGe14b67J3WJg+A+VwSIuZ3UZr0fWs2U16Ag
F94Wdg86693orlXytnjO956nO5gb5yqVF7ZHz6Moxh45U+B6gnTds4lXdXRek3GM
ttfLowL8iSihRjUpXRsZ1ysUYptPUiq0C7h6vlwQyIpMVJAuv0rI6uMkh/NYNByW
qEMbR/1iFbolDAVSbR3NnVJulV7UhW8io7jkiAsG2NS9ozvgnNF5opTMOHmQNLfH
4D7hxQRMass9tIfcdxlXft6fFBCC73T50giySaBVgKkVKdbBIDQHjvLIMeDzTmSD
HMyf4lCFHqOllIXrDj/v7U2PueSNI66ckq4xLBRH1qa4KiICSUibf0YJdJPWY4g0
fRAkZLuI2PxgsAJKNnb17FWCDxdBkT4mPFIhYMJOW98AMc6kULCCL80X532NHxBy
fR8ftenhXe5tEA3kDuqo1qaU+byNbSrmnJklS/whIhmeEukgWywdZoci6VzkY1AB
aFt4zHjb9dlHvhX2TozuCgRmX6kLGH5JqaW9IDyYY8cCTiTKHObMA3kouK/eSbde
++Dx0Oh7tt5JcYLqEx9+X0FrD486MoSChP2xofrv51+yNiI914zfiI7rMzheuVuc
XMzSqzN2D0Ek3YzZZefHungbmFFfF7o+8az3Mh2uwNHuOOgprm8An1qxpqUNWg1d
nrOITIB4vz8tQk29COe8ymEDCMtUuMxPzShcs64p5YEJcjCqhmAviHtfuJqgCZNW
8H+vo09v3RN3j1Gnz544vv82V/NEn7TTgXgdaQCnmWdgNjuJKvtLb9h+gBRgkMDw
AS85cd3aK9ritJFimK5KTSZeMTsR5wAGH8GV5ixglmK1hRyZDit3bD1bGOliytUe
a/PMNsesABkkCKhnedzd6vLrdHPt41veW1NcRXLOeQVRdCu3rF9JYXfODH/ONRS0
+dCNki62d6NFY9/OUBfvunztNxxLadDUaUI74gOlvSVAQvXpgldxur4oW0ceGVL6
0Igortc5rgGo7ALtWaubdKmS/Ajg5a30Nzc/XL4EGRDJCa/b2JpAG4T4JU2myQkF
j9nAL4qylZLDf05x67frZSd3EtLjjufov2wwb608u43dS8x82hAGpSUPV1JtPKXz
lJbjxxfWZiyrRzLPUMUKmzhu7hNYxb+2Cdj+KTPsufp8+Ed4RVh4a3wsfPSuK4Jy
FfJ0DTnrKX4j2WEosCtyZTLfxOm4WpzZpw4AktNhc9JQzwNVck6utxkDgkf2Z+2c
XrPusOXYDbr5Zafbc/PtLukInBWiW/DbI4i1TbdxED3mK1LPG2EQthvqljkIK+m2
8GRgiUCZLN/xDfI1xoxPgLdrjiix7s8fUFVrV84UmTC/Y/LiK3YF1mwxpmwzLynq
3TM0WXDmx/MELH9etiKRSIabqbZcHI4Y8J3TEI6hqc4p4TTKoMWsIRXoj/IlUfCT
xZMgHwfQZ5oR1Q3jy999zwIaEziRMlVEdaOcd5OZRrd/SxLbOSYpkNqIjhdshGOE
4FzgKShbmBpcmz3qTlNjSw/Yt9SRkBL9JuFlpHmhFK80IZ0EOXvDAIKMt6EpS1NQ
+Sa3Hbfspu2XKI2O5tTNw2LJslOp/dR0IdgsNKI0LbW3mFcbODKycaW+zUw4gBkx
P6ANBQr390SglHRowNU4ShcGmYERNA+b0Cwg2SYOe5VT5ftFWLP0tKRQwGAKKLoH
LshjI4OmHGPbOBmFou3JbqK8w4XMta//o2hjVGKxrSVXEqVlQSnTWxM1dp5y+JIH
9E/IYdyD5pRcgMNzcQpLim7dvKMUAtSWQx5oCB7cyHrPam8CxTH05atTpS10nwp0
U1fCZviujURtqkd/KYxgB63quBk4T5a6axNSGsmWyb2QWlSykjdLGsNjdxJ4J5l+
P2JNaw3v071t5lJ2wmGJeRYY6NjG4wZDDRllAvOlePhFQF7RPhhfpg2hCdBTR4Pl
Ri28xxq8nYrc2JBHTO5wYAXLhsx9t5ODp2pYLijCnVdkqZ1WJHjGV2nEwDHu8roO
UCHPljEXen0e6bkDSTmPhVKd+063hEVJa903jIbG7dDVscYa12/mLf0PIkiYrVsP
idi2fVr8kiRkr498C2lUbFyHmWYYrN5Y8xEZxq03FbVJuwXpdiA6XaRyz9CsBnEL
0J93OZjtph4YNxgwfCSCwWkibvuPDV2M0GPsdreBsbEU27JxWNK6kl1kxOuVxhUr
TA3jOe+9I8UW+ZXYKk7Fynj5iHORex5saMNJs+cjMcGeRlbYKbFm69Y8ldcMVWCh
vv8u4SWAhaQu3NHkU8G0PnfHseCbre2BfmRHHi4jWRxNM2r7oJmesI2X04es3eD6
r97ZfSug4edrRESmo3pReCVe/qrBDQV8Kv41J+/5SCES5FuIJWoKkMkzV0EapCVE
Z9WztsoN9e+nbSLi7NEFD3T7uhWJtAFftyenvlrEV5Jhh6IL4IL8ZJ4r/mdeo6uR
O6cfHfTMi5D+oxlHjN3DF0sDnTUVjLmw9cTbVyICOPwmGGeBa+AInDiM74yQLe06
UtaKnYQZLUGvFhoS20k2k+JrypU2v3H+g0wF89oy7sD7TtQYftOGBk0gNE+XKKin
UtJrIDIAbd8Q39MLQ2Ns7KBQiP4BKKxTBF1HvZt47QituqtfzjXxtaAMBIv95m95
b4JToacSDOrLvNtZJWPsWcf54Ezj/SCGPLt6DmptPSy+GOlr2jbI7nV86wQdJY53
to5NfH/S1wEdrSAQugI9AzXveC97G9cfIMYwEnvBVl856Fqeg+QOEFwzpuxONfW8
5QNiWin2XQGEJtDei0DTFLtF9R8VM31jf/Mr7CKw4bUMRaaQ6mFBgc9fDATyGKv0
6pfoU41BvkYA+09B+IcijuqzWxxn40K0hCY80qBcOq+ysXvsfHQG88dC77makOR/
VWvxrfyK0aiXrlW4+71Dd46uuB9i2IBJyGlwSZWjeFOPFr/IFDQcRny8JPYQIcY1
JS/FgEVPR9zzM2hB3UQOTXz655444O5eci1zn4MHg/IRZ/dpd5Fy8ewrsiMCCqhd
VUMf3J1xHuKFbh8QyXdMsN7IIc2lBXMxLF6l45wZZsAkj7r1160gNltIDaDkUEj5
J1YCrhnOosXLssMw17l3uEluDwycBob6CdOAeN9RDHIa9y8VvNdVReoTJLUurWLQ
a31QH4KyuMytPWtp+yPyvaEi0fG/cZE0IVtXsy3cYeUVNR3xGR5DtN5lZVy9A3X0
AfZmaaElUFfiCm6+jngdsppwC/P9v85+6naEAl8Afg02z7Qmaa5afVEN7HfIozCb
w8QJ+mMId1nbvSxKlRLanILg57bUzR6qqQJd0LCG3q/RwQSWIrSbS44e2/gDHmof
ILtPz5QvkNuRmjG9h1AG+gjtn339VqwyCqtC+5OfLhNpzRNrIGXGKDQ17kjy0l+G
V5nQVEnO4IcDBNZGtN0Sz7XM3NMYk9R1ef4F0d6XSdtL/i9ZV6JbBxrS/7TCbm4j
FajjPg4upRMObbuuVGoEEyZhfkafMoQzGRZwwe0NIbhy9pxQBgfaQbg7RaCwDFht
FhUPfECn9+D3Z+7x5hsEotr08JqiFZIPoSuDBwdNrlHDV72TS8ZqJpvL9Kx6mT2G
0bfWu9Zzqcse5itJyGgK8oNNRoBCs7+eOO9uJsSTefWprHQJA31t8Z8rVi8eNUjy
epVj4PvCqkTYV2ie+1MwkX5cBV7PgwHFaav7XCuB+XdPLwgG4wKa4GCS3PKS0dWj
1rUTLO0YdNh2D+8sWjzhSepQvY36GCkio4uE64tjZifV6Bm03SmDxxsX9r8EPBE2
fpl4s7ARR4KNGn1kdA7O5Uu5notYgQJTSEgyKM1dAThXC1QIQD57i02neLlgQYq/
0MpZNGo9aUuI/HNKBmbMFeEsdJ6ZQEfZ00fyzch+uE+8fblrCRsTmX06ml0iST8C
Euzn/GToNiG1rHARcNdELfcIRtS22ShI0clB5SiqASLkBIP2HOc4g74owxsXkXUg
6jeryDngH+F6wCsfGAlK3ryTle0HaYEKE+Vb1/DRNJzLjeuk6X+Sc5RdhBmdwPPr
LscDLsTjpjCqIGYIbKF4NtfKOYPxWb1VwrvOgPLGb8IYaJz43K1Wtcm/rp/vwhSi
y1K7THXKS74JAyWx/8nl9m8p3ti2r6smQaDD3LiKVILMhRqVMgX3GSy9kOatQ83s
IXSw/rBEUcMlVn24HJmXd42uZ1LssNAjlteCyyFp4II5LkQ6KSeJwDNEIzPHllY5
i99X4cQh1sWT01jTt6vEJr+GcTEtWWUuuF9BJWse6MsIqoUFIyVIdDa/apQUYKtI
EZiH29SWmWK4nADxHq4wqa2PapAIcbfp2RGmvW5NaQy5AKaKMYJvqtaWtxrTC64I
Nar1b0xWrXR6McPrrv7qU4H6T2Oiuc586PfKOHRfX4JvAc+xkr8VAjUej6/0NED4
kHJqnZvg37KYSXLeR1eRsH3kRrvI9yqFVRex5nZoJ23cV7zdnuhJwl2uEBGAUDNA
lA6PyuBDdJJDwDaiEl5oNJDCJNA58jzaNi/Grp4lRGYRmHzLILY8ZgJ4y/R3ylU4
BRRIbm1+jV9IzQDJROUeG5lkbCeSatT6hysi3S/XN3fwweW6cBTlWYovMdFV0IVL
jVwhQaRVExwunRLffWJKNZ9VcElLlpwUgV79hgIxK19PLuDNdVuCaiQAhEtJtP3r
5clFxk7CCstg1p7P5oIx00DM30LB3sJLm0Jnc8Er8jCSD7Te1MmcrHSkkqZUHqir
CNaplxjifTwXqn88Mt3//v4JrWPUwZb1Q9SPnr5gp8Pb8aP9vqvEsTvxms/shHYM
wCFQvuptHyjc1TNr/2VDvTC24YPPsUmxQ5DkuLzVOgENIRB0Xyd18+UYqZyuseN/
ZmDOxyxdBg+OK52lp7r88NkMaVy+MLhUIW3/y/GHrh2bD9aos77eIi+dMZfDHW4X
aDH20AAqenGV0Dw3NVZM9TALGlQW9IpVjHY40bRTaZticNjoO9aNNp+Vi88T0zgs
Jb+eRj08CLTenlwvXJ4ZpdmmybwRiGqUkWAOWXf3aJc6a1FaWp7LpyZrTHb6P5rv
T7elU3ryTw9f9EH/NTS5YyVfRzSFgiyZi2tjAcArzC+le+4bIXtoEHLNUkkwAUHo
F1/Ma28DMEbwBqtZLiHL4CY6ybAjUBG6/H7rke+6A7kGps6dXnJL6uZOcnQzcWRb
oQV/QCegUOUeuWlJXkQ0y/io4RWokBYSV1sVVkQeYIGMIctMX6neI9Tuctqgjejz
5kX+IN0qj1vozfpWhFqxeQ7Z9ph87wrj2aIC5OB267KJttuWnnSOqyawLsEQ+XyB
9Ly0ezr+TqT1/mnoGN/H5/0XHoMLuKvftm7/4Eset66JNY/R3blMse1ePlcHIV6Z
/hdN44TfVI+IxAqXyr59cRvsgzT0NcJ8kM1yopCCeqZcTNhYVzO/XQhV7V9wywj7
lxA5jF8Nrtma1fg/S4Z/4PGNW01xZwapWmqeb0JxyjoKYFAXJ/59vM2fGzcpiHlF
+Caowy634WYzS0vh4LgUWsMwD+8eolxotvf6ShlJhdrPtwmFClR7b/duVYitCEXZ
BO6l6Ka8uLnU6drAmvR7Pi3jMItgoFHUu2V6DkQMzYAovnSU9SrRZKygPDLNBiyg
p4x/I7cayOaqEBS25X9VjjL/kzFFtP5xArruOEUQtvo4nwre/lTn6wTc3Fux77t0
wcHtY2TiuS9AjcjTg1v7bM3UvsqZxO2u9N4ZmPQjM4muW3R9K4ZdBOO8jqA3HG+9
xBVmW2t+DkLQU9iGdnk8CS9aRMikXIya1z0ujx9mKsudDw2zDATog7PYtdR/cF2S
T50IrGWkkmkL+MnOApSr1738J4Jcyn/jVWjx6t5Y4JJKTiBfejY/ZDpUg28lKfAu
fNgtAqRRkU1hOogPiT1tyg+pAv7xxXaxkeGZWqcPnIGyD1KofMPAaOE4rYZ3/zAz
6DYz/5Ye9EdeNCfu2vDZZ48xnhUGD3hzgIc07cMFr8yiQEnfJ+/so6N5cfsYzLF2
3oky5brO9ygcdC72zmv5ZFtr2A3OyxD830WSNe4VZn01a/EmEUrpawTfodZlTi2X
fbj5deRZu+pLHw22ICpLtIgiSyZAwffZqWuRCq0xbbz7mJ4TCvGXbeoNVmeGHqJG
s9uqVaI6+Elx+4QFHhHLu6lEaB7PiZipyzswgCaaNS+PdaXTeX77w9fMO37Vi3dY
ALkOfpVUaipGPMExR7iSEoF2Su1+7RiofEAc/mcvcDVFCYU07M+IQTpahBvLSxAh
0EMd4E7NFIf5bJ6yMbam73lz7XTbFhrRatm1sIHVgQ67QD5DTfFE/sTp26JCmPaZ
ruQE6zD8gNT12mJuZlQgNUggogqLFkgDeeHa4EV67KyNvVqYGAwrW31sbrKcDkss
G7MawWMhadaLJO2sZG90eXii2gU609hyHYOycAfVdxHMJQnjz0jq7BfpPYi/xib1
GoSJlBy0PQPowVo5p8crZ4SaTCTeiQedRj+ehVTo5S1+yeevN23QL0yFYJxdsGgk
CJ70d4g5k8XU4+BAG/S/DF050eTN8XknTsTTUWTGr1gh+mc7jQLQUUgoyrZtjrBU
/U8g27M6BeX2AbKJbC0AzVtIslGHpOE5tBx4uVxAvdTa5Yh7M1E4iAUlLW9HdPUt
C5wfVsqTqilUGlZPfAlAzagMV92FnVOmF+NFgMWGTf5R4fRNLBm3JSusckx8nD84
UyKvdaEQhEA1qx2QgA48PxKmK+uq1e9QeF2Ha7O5urFH2LMvJ19fmJfH1Pwfsoju
4vOpEu+hs9BKdHvIM8dHeBFJVCGVRlx0OVP7Al/g6onkhXY4pPpf7e6psIcFbYAz
d6D0GSHdsfEG4EMkbDOU6y+Unnz8yOkf5tgr2pd2QLgOeWr14bDVnK6cY7jGUpiR
u+PXjanFyx/1O6gMXtxQ5gH24pBNnm4RvybNxOgOA/GcnZNrMDXpOZ4krj8l6mvc
DPVuaT82M2ZcGT5C3mKgcv+0f7OUBdHvnF24MY6nX9QklVcxWvLKgO1CJo41Nou8
bdSsZKnrnIIzlaVnbkdlOr84r31sEWpJVBFNH8hJ7zRBBEGgFpVIS6AS7l91QkGO
3O9/9i3D5sO/epRNH9gTrr2ulOvhkcQdq/sFAIe2cTad52cABmPZxK1G4UiuklZ4
LZSsbkB6nw4TJ5tIr/awxzvXTMwvpRSCpEq3am0LF0ssRQqNHt9lEU6bBdjgTa+u
n/1yTb9WBHHk70dWsAxMetknMmYpjkzIkQTdDouLt8tHK0+cEyTd1t/P7EP7YywL
hu2kYGADV5MI1C96ofHVsZk1ItVEo0dDHW3gEGeaOVfGQe3Dilkb7tHAmeolIWbQ
Km0Utx8Ckp+Y/VHRBh+Ww6Xzz84w5K3R+/pkUkdCJ3rnbbMc51kAj2Zb5D80QA8p
bDt9wxVx4DIwIn07fczzj1ptn18t7C2ILRySvQ3u+YOcJc3VoKGgUApTaQW0GCv7
SBm6DmWsdcm4V7Y8QkTZOjZZVso+frXFJOi7SZbhSMEpBh5fZj7Hm6IvEO35g/Lp
gc5OH13Z2Hcf3LW88T9NuE4lwvksW/i7GzOt2kj3kwHaMUVwFZtf3APDzjfS7wt8
+hUp4CtbLExdTHBahiU/0RVMpXJF2bNzIZ9JUr/CqWFxW6NVvU7QqX25NV4Pxd5z
xISk/DlvI1BVIu+9Q5lgj0akPxMiirxAlZjs3ZjrNuL/qVEd/+sT5CpbfArxy4XB
MTjhg4EwXg3FDjpB/pyDE+Oga7LBqryIWTLnHM9WRPzi4zW4fLo/mkwpsIMuLYA2
+r9+PzjhqCm9jEMNnU8D7MUQeRZ9L08d+hfHSiWHq9PQVqQxGpNT1rUVh9EgcvbM
Tk7JZz3u5FbkvP3Tzn/TdPPGD4BjvCn41THuHxuKtE5KBYOjrRNF1qc1ydjBkb80
Mrjsu9rvQyepxqkIl09QhQoIVpHZxOD701mXClIJg7LVgWOStQ6zp4M14DvMJlmi
g+OHmYsuybeWGKaDr6s/hiMm9WI1zWVWzq7OewTuo1G6KtCcN8dE2QqtbNejpqBt
Xas8EgCvNHOTZrS11WlKvO9ntQ6zQpMDT4NSlrIvsDvUBOf3jRpbS//BEthiYqc6
iSJEnb14idXHiGFvxxsHoCQn+M7OM6cMlQ2cDfeCqVHE0ov5z01ca7va1qW8rvHL
tGYGaA9V74V+z4pBBqMC+84Ka8PM7jaszwZyy9pkFXjFIsosVK5bzwJhDACnn3Kj
y0foayGwDaTZba4gGtdLcZnZhSLIm4EE8T7YjbHp2jlRJTK1d3eoUTEZ5e2YN3X9
RqX7NwyC0KOV7erJwLNi4mymD7PyyvGJxQUoGU6fVhyuqq0KRax4iqFrFpQXK7Zn
h0grgwd51AL9SCpoOz/UEdDiW0h6eEztiHkEAmIJaLXX/9X3xs2lYBnjqhQdf97s
8YtJ81Brt4a98AyF/dJHHTHOJWOy9kYDgw7Cn8MT0nv6nxE6o+E/bNS20ZX0evKw
YrQTUhDvfCgSwHwzAhhrSjeXo7vH6bu9Dyo4QrdHXORbQ7/kes8g+8vqPE5GEvSB
wRLkZg3hdSd/VOx/XktOxQbVXTKErto+kbKR6vdZi56zm3h7Yw2pxVxconY0SzVU
cjYnGoQ5yEsICX3mfw02CfUOgsbbRx8Nl0P8pkNqO3Sy4wvz8fDRsGOb2twSALFG
c9XmQkGSPOlaCUwknB+HQsdV4F4t1uSl7OK4zGhaSc+8zkPkTwlV9TY1Zwewgqoc
rk9tf16uK3wX5GqLDBUTXykxgfDLFU13T78HTpb4UccjfdlEsOwevwz4qjc8JMgf
xaZ8qaOo32EELsDQkNZKEDJbrM+2XNllCAjRGgqlhik6B4ue5FbXZWaXqaiCCljs
EcUAaAc/+iigQ1ASKw+czzHsUp0BxQpwsqTzV9UVeZj/UV3kcDWWVcVLUdYPm1VW
+8c34Tfxa6Dl5LzAIrXIOXyXUtPTGYtRParqoQ4ef6c6dah34addIUVNuIB4X15u
cXqCSGDSALyxyKc+U5VhmT+uafPVqrsKX0SxZiT0g5MRmdq0vUcrq4mSCvCfTleu
UjpKExZmTfU9s150FuvMavwCDbgqcpMY4Ry4NBpzE0GowfZAJaMSw3YREMX/JKfC
7oz8DeLq7KWCqkW7ZRzeEMnH++uELPXts3Nt7bykcPw5VomdwUa9N0fMGrCZIvX4
kV+uxiuRkE6oTFXuTp2SN03cpiCvOagpu4XQ+DJJRLs8ZriJv8wXaD8lo7PiRZ+/
DUif/r3jJ+WgeVgeTJ08ZGualikYXV1UqDgDaeAZoZc9gTnE/vOTS1YLhp0NfTq4
g0RzuUrRXLRo5124NRP3uEUvNglPmrKkd0LIGKxMaFc6A05jhGfTSgKxfR0F/AUr
PVpoMqJ+TM4qHfBRzEQEel/QwlBnfvM9Q13UyuQpyl4QPnuVITuV4tvZmzSqI3+F
bMLPZoWz1vH71+ry2pM6RwfzuoiYg3+DM+CY0S2cKrC83UWJ2al5a0dY5mkObIOI
zxd1ilxkZzYSut5U/ffyp4Sdi4mdVZcQGfTNmwqmEBUC1f+kOXbu3oMknTECDpGL
gYou35xFnEE7PNOQsvhvTtE8sdUdc7HUjW/A+1aH/i+9VH0YMnWd4TbVwSU5b207
MPotImHDvlv/NLJTSr3cSuLzpTIhqo1v3EhHQkZZYWD2WEMskNAIHHTNAsj4tTRS
moxNITROv85lpo6S0HAQPTDtnh2c6BO5IDyRcW1DzkbrcrpTeOGofI8xsXF2GZTc
J7EvAyj2Nzc738CAiHyEA3v01yHKSSw8yCXx0ZmzdDS4MUzvJWeW6G24gaW8zP5p
Goo8y8fXqjgAJnC4osi8HBaPE2A+xl5BSma4k8LgTOQzE+3Vv/VJWOli6n0uzRZG
pwGTBU1++ZJjbc4b0Nx3pP+r5jXutR8zJsXGsgE1vTD4deQqXcwvlwKOQlOlMjax
BUBdDb8MXU2ZNH3wcO8RIVyikic4VhhshXby+lwS3CsOq4ytcrcgQFg6drYzHImW
B/L92worEHMkYh06zXYf6XVTvmzM0xhREBaIlkay051NM7DzXNWnNp8SVmrz0uwu
gxWKja+pm4Q6BR4KMkLapSje9LfHYvqqFGPKrEDihEqQY5oqJorKKcvbC9WWsa05
Mz/CynKq2mic2JzEevoUlGoDM0u4pPMHQEAvxd9G5qeZIyCWUgjCZXSAF+GXfQZn
zzS2efiydfJp3p3gsVh05N/6mzN6m1hmmFI1NdpAckzx4YsduoFUY1JQaPkTb1DE
T4IyD6+hfUk1Cnx+4pGnSPcvhQrOh2xTXP6tWTvZy6GPmUZheXCu5j5N8vfH8u69
uxzFYZ5qwynJjzv1OWstWFNh911Ksf+uvmU9vhAJv59CFPjcpBTqOA1k/DKiDPug
ho+iDPLuakCW3xDHoy/SpodHE9ahWrE7EW5viIapIChKYlJn/x2/oqDAVqT78tA5
AwRidU5Kq3xiYdj5B+NDn/T2iv8EKDXOCDxt1uQVDowSlzZnDETd2Ecq1KWv1M0Q
292WN86zYNH/7pT/asNYAQy/sUZihhRBq9tLSppw9t3Mup+RcqWlu3fifv0M1iGw
1WfG/NplFqwkpcD4mM98vyBL0Yam7e+cmc8FrRagVWqVkPqLflL4P2lxpOcEmq36
1dGaG9P2fiw9YSMRjwKgS+IbsGuk03DcnOwIrlM3Qp8pgx6mPkrcKaP6hEG2mfaC
oOibiPwOYBg/B6VvPRqWgxXTIRfU1Y+OT211HkReUUjRZagsl4XewzYDcOHpCZ7l
aHnU8VOEzYpp7hj4dwdsagJETW/T2PPJk8OeWfBDuUDznaMwFx1p/t4VfotWq3zc
Uzv1qUbUiDZf6JMHU42UVc2yf/gjQ+shX3T8Vp6Ebk2JjP0VnHIG4MQrr8gYqwIx
hjqBiTD6uVYVYwQ7KuxHRuNAiKIW7DOQWsj5TW70KuWrJtwJsbeIjY4DwQ5usihG
qmPuBE7VbU4j2C6HhhPNAIFvT0YFQdwwcTxNqhz6V8uvl2lCHUgHwUMfjE1HWTgH
Zht1NT5A1M9kqYreQyr0qsXoFWpibb/Pt9RGkV0rGrqyb0DeWs7brWAXwfB9dMOl
b8LbrcGXN7C9I35xIzCSwrN257Rgtovkvhryg0lxRMWM1VldT2t0Qb/X1ljinEfT
1dlMn8HKGffE2OwJ/XxRoyAbBF1urz89Cy54U+DchoNQmsmXl/aURD/o53xc3kq0
aMkIcmiDsb98HWB+UURHRDjioQNuEzUVsWEbVRBq9N+OCC71/ofPUrk/6Py1h7hO
VlBDUj87JMZjfqhItZXlubnSjBl7ppgw45whxJptNMOjHGdQ/wv/506W/jiEOVZx
Vyog2WpVt4A3ESRsEnOhYAPG4ropZylDSsx1aysU06rJMHkTsQ4z1P51eNV0ae3Z
wKFnVmDNvD6gv79PfytQRcoOuFAhosD0bsOYTjChF3oZL/6IlpNzkjhlAXe9FfO3
kwx0ZSh8ic8Z2/N9f+qfvFgi5gwtv9nWiFdQu3eBxes/QkXDmgJoQDwbAL5Sqm5n
eqToK6DC0NmVs3QdnKfvg+7QPJ9hGyhbgJRrER2dxvUX76lga4/wx9xQ4A0drRGr
Al7BezWWJv+zzGMz4qsylawJ7LXlAO6OL/Omk3JmuvAw12TZlhs9v6S7qXZ31/gt
qoYVdyAjz3RL8AyCS9ExIABvwyODqumjN1U0ghvRSndL+AlAzEf2l1DSekyANC7T
LkWM5jD8iMHnXeNBwcVt7pnla6mBolxtMR1cMRuI2Lai/FOqMvCzIHw3/TOozyW3
lXDr5rqWPU+I/uMrOsFiDmW3OvckK69RLzwtBSxs1wKaaLGtLlc6WV/U7DSz2OQm
t/WuKxeHjwzSPTxg2/xNDDlR0OpzM3+mvc9kAwnumVB9waECLmgKFlFhoJaZyO9K
+eMyR53rQXVJZBJxrMZrmr7ILNrwWOFD95rdEjd1i1tqMDbs9SOmfzGKd6v+N4TF
KdZM6xcaFSmFkXajIqkb0e59yS99lYmSu7T2z+EeBjLOWsIbyLtxvAv91FLpfo3B
txJwoVSDGw2XryNJ6sX8Fw167qDuFN8/e+FY8p/Ib+xZTq98J4MShTdhPSQ366nk
tjsqwAy5f+IBitoCB7ylrr7HANk3yxUMY4FJCauG/oLqbPyzrld/QfRm37keVwvB
sATT5dCdwwfjYIr5LuJPKqKcZa9B5i6Y9kDKeZZr3xuv0+lpSp0X2zOL6fvSLkc+
wifACUF7i2CjCukmerbgvNywSQ2qBSegEdKvZ5qPifQ/yaDfzfaUoxTsziYFvLOx
Zkr1s3xBwlqOKBA2fZJrn05RnJL+88bPJ4AZsFDUI1IIGBZAguK3k0gxRTrh5COY
o4a1qw5k7OUT5hyCsv7px8b0evYpYMSXQIT3MAXp8daJtOQYyLElJYuANRkxvACt
X5HMzWkLsXZ5somMRS+JXxTWkgSTJ2HVtslrnEA2lDqWPBKlICwgw/eR0AtCqULE
xBQ0u0SLtc8XNZWDtI9nGKQb1V14bgRDpogpGdyhv1qdaEjrnET+VaDItCpPa8bX
O3iCNjnHVTDF2au7vUi29fBln2GnIFWfpVa4p5dwZ/3r/gh9m4Gqh02KEAzeC0lO
j/1PGk49fzHVhL10ra2ml0SfJZfJ43El6mibNs5SZXYsU+yw3jAk8vCjwH2TSwrZ
YwBdwFbNTK6v7rXEodk0l4ODaDO+UZgAczS3iyhQSUpXN5ZRabGqslyaZEI83A2j
Jhq6quPnU2G1pj2WZHDZ0EUWjOFnX5SvkGZXFV1+55GEOOSUjYV2dcg+doB4sN3T
mAfemJfP1/y3cHcXB4G4GNCinteqquBhXQ2DK2Qmbvi9x1xRDOQuuhPXMPOcr+GY
o+GGzmF4w/KUKhsVTjKqJUbRPCgEmTPforAXZk1wttulsM+mf7GDbbwblFPh04BO
058CnfmqcT583fFjbbalLNx6pgAsY4IO3RW8YZctDjDVBb7TeTVrK4gSf+CI7gXN
+3hovrySQzbWaHhNxw6MMJFbuukzMNU4eZkjphZRgo2mMlsB/a/zbd9nBiliXNG7
XlI+4gfrpXyBBlkVKJwKohC/RPyHY0cg/i8inGnz+u3e1vHlwx2tLUJZrbzM0vVj
LdYaIjoHyMmjI21fMEjiXlwsKJc44huPFkcKSnxpLInGletrW2D6r0Que5NmUS8y
iHrvaNUqh2/cO0NPq4QJfN+74FMtcTWC2gefA1qgUGqmDVbGrY3l0l5Rtki2fjV/
PHxlT5H1LqhFsfMvCccY3BCFqRpLV7K1Tw7acyPHd0om69GzF/KaYsgg5GYhpEvW
GJeZqfdv6n+daQZyqoEGo6Vol/E97g6FcI+ObV8YjBMX28AqI2qNVZIKl9xMalvW
s7N8erauUGE0sQNp8vtbMKHfMT8gkr9eKPiu886Ubr1MrfnR4sW+ex1XQ0Xklaol
KdcAUqCdY7TmjNQdQiyabfpY9PsIqyBZ09hLCfotetNgHhG0MDXNKuiuiYnpIi2t
S5VgjgIpVwqfSDAPubfXJGV0mYS4v9kRlyPit9/tqxkJkCmXGM1bjt4rLBWzDevD
RqUIjfS9BYhsS7PjqrrEWAGO+XTjhHkDtpjt3b5mILbmyI3fgUZQUKvYP3Nej3Ol
EXBsBc4E4aw4nrQqhMRleRPOsrHg+nK4Pmp767952MEGJeSyi2PQXyA069reWEG9
YkfK+aiYf4whkPl8GbQTp7zFAUz9KTsOFXWA/8tLn3TNNS6gx+FxWTeufbQVeWjj
mjWTERhXayGVjLd8M6zjrzaHPZhXG01V0F5sMndOOeqTRGozZJss2ahtZLm0czLZ
bKvQ5aNFllir8BqV1z+yGSGKxVYXpbzeI/Slg0/+jboQHODFkQsfyh8HRjiNX1vO
dKjRSRm7IJXKnahQwu13jSbtoS9OMZTi7Ca+zTg9WVGrn5UNqiLFb55/5PmYWSb8
zCuBBWg0crIv2bwRnoFOFsd2Sn9GtS5bRsm4DpEVQaEkH9k6v18E6Sl6S5GFWksy
Clz7EbBqeQTe3Kl5X4y8QPxCnkd2hC8eO9njDZ6OQEUmn7OblwhZESzsLC4KhbJJ
8WPGlKuPqDOFGtuktQXOKX7+ip0Ge8oCJ0kinenFJnng9fzZi4GffttE7HuZY508
J29LJQoMaVZ/+/s7r8UNFFPrdKoxUZZ243pXrcxuVlqTzpkFB6nM22bfFcVYm6NM
SHlIxuHmTd3jyBjHDBOcQSuF0TE8apvj1fODOiy7KxSx2bQ+62ZX8V++Pf7/B9VR
BnVfQum/lvUfwI9IATF7DlUptiESmun5Uuw4lP4SW9ONCQeOnBAx+JJpuwBAoTL2
teYqqLchE9WEsAdZP7dA4ZkFPZhdLW4gjKHP2Mnxs7Vfoa03Skkku4xtnddPboh0
KWFNYy+bpeejP9TOVB4YBzmQEc9X8mOC9cmj4SKQBax/D2a9Po5TL2i942JwpauN
lZvvD5rF6ekkPtuRmHuHkO7oX863wEReMcgj4ERJbJ/lVxKo8w2ue2d/mJ//fiyk
DTGCkpqRxFShAMXgPXj97D91silDQO0Z0gfTKekejmFVYq+nJMTrMBWDlnhB6o53
ODiVIwXKsylgAOrocurL0PYz1yCS2FzAgnE2DUn+R5lCOo+ertRIlS2PsfUHTpBK
cTb8ALckbiv+AEzdxfKKHwyxZ1CL5KtwfGQ5h8fgVZpmd6m6uB9oCq2WLam8HjiJ
VXtK+ml0WEHRKVArWjT3XWRDtjOg3DdkXg4wqq8nYS6PQEcrX1A9Bup8kKrkSUMj
Qb9KwnEAxvLbV+3iNuFrPT6PPU7Ds7hdBsUXvjUhJo42hWvffsXgSwgOEe7rJ5EK
AE1iVrcTMOx74LZK7MwEk0IGL4sejf9c8ZziPo8FjUb3fhe+FX7hvVNxs70dRl7u
AhsWpZUDKfNk5I81HH2O4ioJFrXsxXP2unIeuF0uU2ktJZNk4IpPT/uXC9zFTWmW
aFOilXnHy4RUQCcSrxkaMwUzq2eCj6ixQd+qid2opHfQR0fnsbpoLt/bU1cIb4xV
FEqk856xsPKKmYtOgUMjwYDzfxWrjFSin8M3ye0PA+CwhRdgZJEim8uHdxgju7lB
DYtj3fbchcSniEE9UFULMdJS4RiINrxai0fMEcm2QOhK2SzAob9IQEhY7wsizMgL
741iuV6tijgpquUjjLTgcJsDTz6pylMLjJxVoB4PSkJSGKyDxB6naUIBBzPXoTBp
XhR/ncL7MN5HsuGCZIOviosQxZWraSOBGNqRDaMbw4s+fvSaEYwBLk+Lh8xXD1fy
21pkw3JF2uk7kYr6u9xnKRBES1ytexALPpcyvAkmdiJoharmp4hL2n0G1ks5RO3I
GPMhB0arkUlrkjDlRFFm5W66QNJnFF13nbmN785gECvFg3uiDB0qIt0CV2LG40ah
XnIcUc5m2Hxh+wi8XVGJSfyrvUfJ2Lqr0lf51zyvUTzcxUNowwOzkZhXPyGzWlAA
EWoVJEZbq6kpjQxMRbgxaBgS/Qs0hUKSOGRKupmBN/T0Y8HvzAGHlzs1P5J9EVi9
DCFUHRmjdzykx3XLZyI5JpvirVWTRAnLvpudT/3NMLVtnAehz2jqDDAgGGeegQuQ
PXQXGgCPxEeNXSg0/vMJJj7eS+/EJyoHLcm4wVLG7WUwFyUfwLdaAREDR0IPbgAI
kHQRtfrwBwITQRKYS7Aybc9bsSvbUrDIOkfOvPWrhBniHit9uYhkxpTMEFJgqNlK
pouYnFCR9UTs+rlHAGpfWPc4Dn/i0rn1XKXJ91PybVwaeSlEpG0+f5U1U2aTuS57
p/X/EuHZCxVhDAtsAma26W6rfZDwXZ0yGJ5myPJceAgQY7Q4IcEvss/oy7egmvND
utfRsp2dMiqyOGIlL/psO0tE6r5k5AWQuFvEnlgLhYFQGWdK+Ackgi3u1zryR7O8
lodxUlzBnXb0uamvysaRxwTDWd7uhmWLLYUdZ8n2fvk6gfS7PEEZmeNx/UUI3GAc
cdwbgKsAsOXe7u+LM8MInZJMr5mr9Dm8G0PsrlVCpDE5PThDFKWlCHFKCgTa4eV3
3dB1+Fg/evYjZDIQfsxrL8HqULkniqsqmwPRwDcciJ/1kJ9bxPelJYJmSNtwXo2g
yx+I5R6lbw6QtTFswpC7pdwzmlxPaNX91v7r5Su8tlijUGK7urUKb6BiL4+QKpq/
74K3d/G6spks5qDYS8dacX7fDy6/9/Sns95nHeGY8BAOToMRjFkOfog1RLBS/s0R
YBs4n8jFmQu8owC9MicE4y8+fm4ZUb3mpvH8blbW9JaxpkfFnMeHT4QgAV5Rby8K
O3v/infC41F45Hm75TGmJfbXCj5VtJYAtPUx/wb8C4Z6bMOx+uTXtYjzJAHF7Xre
33QT7x7B2bKu7fNGRiadf3fxJytFcxOjK1w+daEgO+2GX1xOqITW5WDo1MV++OBu
2NNymO18awtUyndhpjjyY2z5EiDwvSbMZPAtSnEm1BiUJCpcus2o7LphV+JYfm97
IvyEGu7PjscbboUbsluPB82kUQ3Ee5JN0I1Rv7brewrsYLY6qRqutFB9kKUNYq+C
/ZfbTKXioIbyERUQizM1yZ+XuuG3Tn8T+iZSMnUhnX42xdM0fcxTQHFJtID4Eq8q
FSWxW8ne2EkRnmGg15zocR9ZeIqUzQMtUofREdXECpqPHeyui5aMezKuusPj2NT6
t4IQEbd8FMASFHTpUinQhFhrX+1jrTJRWpQnugGPMOUImQ9hafw2QIhEENKoEQJH
OS6M0Iczuui5pSIbscRP/f//Z14RVL+GPVuzsdnw7+XH8ASfIPGgfGSgpTnt04U2
ricz8FgYwnaD1imU1C5JyvO5DdAC2stScT2cwnZ1dUl+QxBQLcJD/apx/NR1u111
69HJmzRqm7UrTqez3KffYCTZDADOIHPiP/DbC6W/QOXyuX5kPlFtJT/9lavA25Ft
IOJGZRhSYycAAgb1/fgE6MWFLLdvXzsow/Tumled9ABDvE3kmoQhGs4docPsT+yS
osCSufmpBjnF5Lq/vUJo64plyXbrxFNdhRFxw4D/w2wg3uH9MrOe5TLYJunUyT+A
1OsTwbYd2i1+ebKyP/fnc/3PfubiKYEwUe5A2yxmCCNY4WJ87baLYekSAvN3c5LW
QdRKCfWmyZZoQ1iUuepodFzTEL9gf4/Rs1Z5e6C2jUzVIQe0mKPfGnlVp0sTiSEm
+oAND1PmLRMWrAEAVJsgSXX3mRM9SPgDdiU6uxmMVlr48nhN3VFuvZhk7DHFmf/h
2q56esAJE/XuRYHD7cHZKHQYU2eLA1w7IlOLXjoLr2sgbUxGsTNOJM7a6XzBhRNp
0wgPeN59t0jwUpTgdAaAw5NVAMWxHBGqD3wwhJM9NEpDEm36Q3idgM8zDRBz2m3G
OwPfhPJNF9aYwcJKraTKqzCS5lRCcuK1KB+bnxLp2COQvaFxUe2Lba62Mn9qgFhL
PlWgrdY0Md3gjQyenESHwhS6BMWNpuRuFRUFqS4zwg2o+VkLkrw9/7W60bJ15pJB
nQCOH/ShBvC5ts54FStjWbdorObN/Eb8rQ1LzMO32BO/sb4v0PN5nXhusr4tRPq4
n9oKz2l5Sr4j1Jhoou4I8ZElkiy1AlhTGMl2kp4lPEADjILyhy0f8cLUssKygceN
uVmH64tFK+HyJpa1t8/S3vilr5NMx7OseIAS01fvP86qwQ7rL+SimZdG8xaZC4ui
+JOt+p+1T/Do00lBWzKtCL8KagTudhXgZXSujk69KqOOPrZ3JlrPWErSsb/OvltO
Ata7ZyfXFatD+iXCwt561OD5EDbSc6rNoi3onwxj5XONiQVKUxsDwVMQN4TA+DbB
ae1Mcvubr46rFkEYcdBg3ZUnj/ewuj7aUeyy8UmmbgtBQG7MSQJ5UHWkD6G3XMW3
8tufnxINLixvkTloEaJk5ekH3Rh8p5qnJErdjVBP2gX5ZDJhWT1kdGUQ7m/70B69
BDE/Z1nj/jRXzvXJhQBFnj36tsWXGdLzGOYd1XLmiVItR1G+ynlfrphVYp8uB6su
7wD6SDZ1ZXzdoOOrbLRrrblSj5Wgh+Xt1+gKKeKBqSHGNYkuVangGwzg9JEamy7o
OkBuVRn709rd5ioiVgUBV/++OJtGldK/BEB7/H3ERjlpFJMx5tfTm46CCJ4K1QXX
Z89Nc1eHqkOdWzi8/ONGiHeWcIFb2lyCkUDJVX4QD4Zb8enLQf2jfGX7amN3m0N+
o+lxJsM+Q/A/U4RjytEgBv60pYVqbmcyD/a4MQMZ7ynFAp+NjV3ngi9r1dLIt4Aw
XTlhWlihbbiIDy8y/HkO7t3UbFqz0+zGSxCzq3pK7aVVfpkyB1tZKXC3AW+tiwdz
hNyfLOjSLGOEI0X8fqk+x1SveSC2UlOxIrj8lubAKokCUfndCLfS+m3T1mjvUThG
CpZ/sfZd2DofV5iCJDpZ5Y65lWDoXZdu21MChb6AaLUkmXxEksgPCZNy6IldFI6a
gnUw+3lKhGaRp/iv6XIkL2SfWsWUa0jk0vIyWNV3UMcNcuiQB5T3N/FcKcM5iaVK
VEnHYOkfKJdTZl2O2CYnlQcLsB8+WSFgPOkiepM2bsPz5FztpJevxX/oyvEwCk1P
aR+Ijwg8P3G/OQ9BFQGRB4njE8r6Et7QGJqIGBmz+0PnDP3Ixn7RRiXM6I0Llqo0
/DlS392wOWMoJr82V+KDKcGOdPeUSLLcwx/jlg5tQGunTADkWwDwt7wPiqabSfQ/
pk8hpC39E+W3wM6iQP6uOj3dTnSMN9kRZyLmghxghhbexbX5Vv8TNFRJEML18vJJ
OYdwAg5xL2R8woRt4jyhnSaxP5EBTOuajs65q7m+BtwyxQXU2LsqtYC9AHTlr/8V
GXZu6ziarBNpG4327Z0wCxLCpFWwjAwIE3PAvaul2q7zmxdzp9ZeVqY9GGtnmXA1
9GiOgpszPKzlfj/+GUpYwq2YSiDIuy1IZmpjGVAMQSeTnDXJ6UmrygHilX7WkTBy
MhMvx+OUmyQ81mY2OnUEc4Td4AtIpHQ2RfvSea0bZ9nzkL6Wti9X1YAe2aUWXKin
fCzO1sGJDIYAD0dTJ/7JL1gOoSstj0qp/af2yAbS5JAPerucdE4+sDiEzeAcJGSK
dqKEGapTsuu7mhTV+zsjz2asH3TPhg1OOswdih+OT8zB/zitVJMhOoT9NSXKRO2S
dIn6jh5JeKsPPDGowA4cyV4qSZwtPfl/zn/5mTur+m8fcEzwrqEsJn9bha4ssGa1
8EPW/fBxYAadVq64Pxu4sqsoGAmu74jfzWujS7XWXH8vTtB1bLiO2g4/iCUWA1O1
aA/JE12nHMN5BT/MZlJ6hkn828LoiNgJkzBT4fy2aXzORaFxTmv/MDwHCytLao2Z
Cg6DgFo59nE4+Kkef2HGo6QQmEe9BdvOdgQt0+1vrr+Clu//E299CiURavok7nEX
CVvQ3WEtHJtjh/6AynWfs+Cxoi5m57VTCRQ1BEJeLYG5K3xzZMmjbijXJqoj8je7
np541OzvTNDLzRy/xIz+45w55ml5Zg66GXnrR+x/qmWre93ZyXEXby5GB2nC2JAH
9+LaBi5ckSp8HzdZqfaOKj/3T0V6R48HovQQsW/Hg37SyWV8xUXmvF++NwzdABfV
LY/U6z/8m44bkVnBWRcocOSME/eQ7V1y9DQVSAasfvAWCr0iRs2WyWlunB3razxS
Qsm8/OYre+ZwavG8QVfUw9ltpjtDtNJ8PXlYssngsllZNrIuIe+JYqmwKFX2uDLo
zcvKT4GaVy4+bST+Z4z1Jux9kiLVBmtizL7J4MI4au75fs+x4qV2E/OaB3OOtUlJ
uVxA6zAO2SjCr8vMvMNXKXDzio3MnKBqFm4gBiPUvOtL9oSRdN1/CsQXqxHVHsTt
Mayrs9Xth2NSd0I88mPNihgZbsYTjfYABHung9QdPOmZZ2aYVCkEjaWRInyE0DDx
Fi8bGP3rr42at14zG99iCUtI8VpkwWW2FcnatE53TwOKVLj+X7UmaAgZqSLh5QbV
x2CEsfteH1fHcNPd/2te7hNC42tfpmLdvHDF341uRRYLXLWvedi309jrPWvz5UUe
FFNclroL31lsyHycuOgRkdaBT4XGy1tLbNzhIZyjzn7zUTdFp6dRazWzdcYm1IRZ
Y4shyR2RSut73kfF4L/AnjOXTsCeSzvv2t6053n/xsuIFOac6SP2Jv0U50vZ3S/J
brsya3YTpt/lwxbbClkF5++YDhuU79ak2hGgQFuDP/xeENHCRqj+UVvObz1vnPFy
H7QSVMRNBjRJ2G31ZPS4r83GauOgGqO7hFQxeY9Oeq+WYgdN9y+JYvpXSm9e6BMm
giwRn7Znl8IBd3oKIEq8DSgmO3sX0UdrhS0v/275O93a6IzXDFcYRF2b7vYVC2rm
nuFBFDy5R4yvzE2e8ZN3Zz6Hq2COFQc6oA5BiNarc9dIQCq8YbS3Yb49peWxOVyy
UyBahZq5GBz372HrGPFP+bgbj4/6lpYkmIyslha5yboIBEF3Nhbmh3jlBvQNoyJX
GKUSmOSQsLr233rK4wlqAL8VxAbEwpRbr7oxLMxsYbMxdKym3oqwvESIxhS/BpQ2
gE6oJqK02naV0E3gLHegbzXjMTdMc+43/+crLN8H7+57cKDq6rQuQ5TL4CORqQ1L
kZpEGRdQCGX99GPU5P6cgMKZRKdilLVCZOEL9Kx/djYkBfz7+/pdaOB2sVieUles
0NCDCfOYGZX2qVXtAFYKA0OyKiHGFYgg/05UBurr6qmS9zwkQeCkSDtYS6RWVDu5
xd0qPvk3KkSDhGbBOL6m0VstA5NzG0AP5EVwAy0VzqNA1w30iCeEGaM8/G8RFmnY
bGw7M99H/hcaaplqNlKH56plyfmWWTU6EYDDu2X9BkinoX9HjMwR9uLoPqE7pzQM
PWD6aPeT80i8eJwhOzf214iheBswy6UVMrgBWftPws8aFQKJUidrPVuOTbF+NaZH
EJQNdgitOL6wfqZOqnSglmVd1kmIz5ehV60ilg51vH+FcZGVPd1Dd2erETPrkb6W
tOcH1k5aFai6LUdsshm5PK2D026DcjILWV/2TFCIt7AQH0HoBhtEnzHC9giynyiT
GtyyQ3S0ECyHDrlgJY/v8sdFFJORyZqFLgR39e15usbPSXN9eBxdvYtF1v3nflwC
nc8sOK166faI/wCJZSnmg//2jDZPfnD+xWp3BywlbGOcrK2lVw2w7rkq2b0UMz3v
8XIR363BO0k8/JcPHMdCJIAVp9lXIe4oE57IO4R/0fHb141dg9jiqJkLsWVptFcV
YmHvE9E2/vEUTWyHf0X03X/qVOgJuQUht+ZB2vRGdVWdTuCNqkFmY2YU8/KtaaoI
QHUrHcCsIGafjJrpQQBjP9Aga6/sfjOruxWRtlBiLAzPs4w8lFW/rwW7AwqMf0OJ
DZUsCKyl+G5lVQ2v11xAiAGUzB0rXhnsD7x+KiCNblmdqD40NboTqMsDSRSPMwBn
xXDCqSvq7SZ9m+zSAufbSIwREAxS5ZhlQCO8f+cQtyPuAymKJyFNZ7Z8wjnvybb/
4ySRg7aJDlapBYqYdUgMxORXgLYuzlHw6Iv/7tB5WXR3QG0td6B7WYJqOfXFHdBZ
OYScF/FLIaDQrTzlt1CZ8GrZSKOcaIkcw1HlSuRvFG6abCj13/pk3++5YHEquv9K
r4qp1XaIA351juOnERLGAFSuLsB7TyfgvhJTZQ8ZAFtnkQ25fA+SPtBSzggxQcHJ
tl5epqAl5MXBZZyS5DPhXqzsA7QvdykRyeiD8fKsp+rvERYKz0/Fpx92ECgWiDh/
jSSF7QPuYJ1Wlx632dTjeeedjf6tOYmiompoMfY46I7fkEgOf+dMLM36LQQm3pVh
Fp3LvGS1jDcHfUP/qptrL6VxR/nPa6XTWZugPtl4PIy8g+Lv7XAB/AAO5pcMVx4Q
t3kBB8050I4WGAazwZLWHYCnLFUkI9FKcibzBvP+UcWLNVwkhoP7phu4ITtB2i6p
7sLzRCJ5RicbfjYZ5MrKhc1X+q9NoGbIc6wLY7Jk/p8RMFERlhjpDdWCq6y3Cogw
9WTjJGxlpU2bz4fFdJ6f+cttxQSQnbgjkD6oXnQvAVEUOXdQpn0bDlATploJx9qx
087NsA4t+BZGrzN8PddjTfIgBvoVK5N32zHHZjD0weKvVCDjv9vWe7FAVKoQvEdO
hFHnt9/qY6nYZcF6oR0VyP17T5bxLYFaO4ddmhEK/6ZbrVfZEVowc2xIaaKSYiuK
Sm64wxhl3LnC8++HucXGux9br6Gp7esNiSTnH4LYzQ+ezq6On/tTG6wiPW05e09a
4LYIIV+RyMstd9t/pgqBKeU1GQE2lEIyIlWXr0XAShFxWLnSBpf7utaOYlxlGXJ6
OSJyfyVc9BfjxmzF4h62+WoP3RujHA2Kqa6U/TOzGOrIDEDUrDLXoucwUEL8elQS
b4n9yskkXKNbLuKDtGmSO4PJXz8oFbu5sFv9in0ZisOacohyyF5agya0o5xiEX8I
Cv0NpP2dPoPWd/LT7dCU2yVUFyp2lIF2ezjvzQImvbWL3yXlKfA/JbLzjZHXhIJk
IEL+iYV8+NOplY+yzoU042/dOnFbi1+c/N+jpeewUsbhHclM+7JHpFS+6aidWfuM
JrIFY0oc0m9vOaQG79P5hAqnSjivgODM4qLAhLS0NhQMonqilTbYsNgKke+AN4S8
wp5FGKxqPMRitMO2TFhPiBy1s1mQdheBTK9NgybL8ciGYzeNUbYJilDbvDcPwoHq
Wz36T4UQeXHVY3i0bVT1Rq1lizK9f2oAgcuyslxW+fHYYYcD1qUBvAvahwcjHjW2
8IDniHEniim74ye0nQbx+1l4K2+jdpYPZ+99bPdAkILzBGm+V1BNve/VwGzROqBa
V89f9tvk+dSI890ErOCPsNZKTCRdvwerne7/RKubAncW8TWoMJYB6ZZPYgOY+2Ig
uMkdklANPGkBn0mUpYtgT89hTQOTbLrJkjDYCYgmyG+T6NrLZFQnJtiAcwL4m0HR
JORnws17Y2LACyakINLivO+ait88C7p1sPUl77yXzlPKeCC3BZlq9Ef/yy4QwLd3
bgsVRcoR05HQJN4mgMhIg9N1GMovufuQaiHnlKYL3Hk89xITGvLnq1H8DzOySum0
dyT/obbegcET84YZ4Tsc3h1vMzHG/aobkwy3+zVgaYCG7lsT6EnuQtMFEXFmaT05
qS10WsfQT2bsz6MVqHOwuCNgy3diEIAXqAsaWRjdmNY7cfVAz4uCiqb9d9KfmO9h
GytXMpvc1HQfNJV6PUzK2bErVOqiLfjpj+tvTeQOzMk3H1altcGDl1hnc6e6ZVjk
0b/ACIJuSn1hHFm7Hv58qt2a7SiNZh9ftrHGfukrcanhk/btUCW/Ux+ptpXRnxwB
Nwsgd7W/VkcTn6S+0fv3YC6AnhADBW1eMHiFkZwXMDPr/k3q1lr4J0SFFYWFIox0
b1M/91TQxkOtfI4SyVQ5r+yoImi8Qe7kkALKsnFNtcEu5/GPEbF29uShtKj0UASn
VH8Wq1X1z0sRFH1QqTsqikiLBfknvWEkTgpLyaFwSIV3As3jpEWZhsZkJJr4aa8m
6GEu48r0iroNpNO0vuE1dTfzRy+QevVOEOf/sUGLKpSo5XOYhQcL3H/KtTlV0wN3
g9nnBX/uWl1RdN/7/Ba4ZhqK1ZT400v4DcSTaDO/MOIt+0lWnLpjMvEPPOIJWVqn
+Hjc7GkJKZkgF6iRhWGMrpgzsRxAjEryd2cdEGWEQqcSQyk/Bj9PxWP5xVMZZI3H
tdOkfEtGhxaDZe+e1aWgD5Sef29OtIJ3GIeEwIKXxgK9nBezpZf/9ECsx2e944Y/
J22+V69MaNXXqEcO4DcFpGFYJB5rm78GXztvw7+qVbisFsZi2v9QLIFQwAhp+Sv4
x0l/u+hwin/b95nb+fVOxRqTUkW69ZKBHI+1DMhO5emECBA2HBDtlWp5uPr6lH+l
7ue6bdS3bi5Pi0NC74NduTFcApMnpi0F1DHq3fmUpanHexWEJHz8CICahv/Lp26u
XsYnzMg0QiDS++mXowdyZ/eF7xyjw834WAAyZRUODmprmj29XbdoeRDwhOcWy69n
b063y+aws+iA84AUOF7AZy5HHdMJmJi/G1MCFTYwYNC0atE6j9/JiBgMwovIoiMM
Sxp/zV+b3qu4ltF0d6s3P5rZMfz1IPZLjo7IfGzsBprrQT/xSKB9XTURITOo+q6A
Shwm2NsQozLft5ujvB2Dr/wtSWC3evHTi8XZqOpVlKqM0oRau1nUPpWWCUyVzSpW
PIXX2Jx/B+UI5oPmYoLR0mNGKDttZ4KetR2PJfdenY935IdsLxZcPr17ua5KJLtA
IBrEQ8a01VP3oD6mm1477YD0d0tC9isEPsUwwxupy1L+T2mqLZX4UBYeck/+kEqm
YKuKa05VhtdtKY2q06vrjO0GQCBgikA7Z96XHcWnvNxR2obFXs2ccEFfKuzN43A5
fA1Jt4TfELmQoyEjv5SLLOLc+9qnZ+kmlGJUt090TzSjcQrUZG5b4x1+p/Z0KES7
W9QSyHOP/APB243QTCgp7/6wmiE2AJR7P9o3c0EhfaWuVESVUvt6XXxRvKj6yKUv
0Fj2esDamYQCPzu37gc0miXjMHUF85N3/oEf1FLvvlKwQZIMApZYc5kT/wZegYLd
Vj+8Fagwpr3Pd+0LG1J1piYVP0LnlVzyxNosTwXXVH+/KTKCa8P5IgIfwStkVC61
U2VTrlCcibq/lCi8cOhyKF1jeGwyj0uCR+ia4W7suUIPLvAxjc2ehJh9VYLY5qJO
iUuaoPZkHgUw9tqrdIgIbpLTUdnt6klGi8OC80x9AHZ49ySTSPD/6fd6o6s7b2i3
1PFR2BXHyJvl/EYdaOSjbbPck+auE6ovOeUxaI7zTGGbA21a2Tyc6IRVQDmd0+0j
yxv4wJUFqQwWAOeUEj7CjuHJRFobouW2wbwBShmjpohqKOwIFPcpeEzKicq6EFdy
NV+fxSHPwFSucBeUutXsT2WbBoOhoOl0TQHwN3s9bfZM2etbRRAMm3hz7siVYWHG
AKE8mbHwMcEIbo/dt2SArgJvFjCRdGdWRBaeP7IZC0IZ6Wjum7ZKDRT/K7YpsTdH
UCPXhcCf6yluyf12yowqcyrtxmW/oJhehAf1HPv/L4CBXUXgGYfaFX9tPxYB0Tia
UTn3wfLzobkxthZgOfs9hQwFYGmR98kHp+oRRe3rQcXPL8Gnja7YM8btB8uJhCHW
XZBtPt4XpRD/bXw6M7HGps4lTKL8taC48P5FD006zb5LjRuYk4aT3xKg1bZLkrA/
gD9jDSOcZ8/ZZxNw0/cM1cPEmv0ik/SGGSHkihXteh+gdeHi2F0O81D5UHZuAz1f
Lh0UpAzXviTgXFo6geH5SWf1a/+3JpktHpwnjmhYEb0ov/odTliehtiPLTJqel+L
igR8M2Ud2sEC6994ZvfIQ31ylTdLkxbD9s7hvOgSN5RHJOJ6REFarnrBZZ5BHZHZ
ZfbA3YS5G0ADmu30IvU3+Tr3BM2HtWUwRsD8b22U6j7yiuVPpnWEPhbUaIOClay0
wFmEkpQvOwo8kZToroioH0wJ4Y2MgUUokZTWHYl8bG6Bj2b5oTNMlkMZaElAOEGo
yyKLEn4Ajq6ld80YltjXmdpk1IUUjRPmnftsS87JGqgHBj1DBfhIm0gFp9LrYbYX
8SQz6WE7IE7Vgm3lXGjbLvIsM4CfkayeN/Vjhu0ZEBsmGJhpNYL3j1IHhZPeZhWu
/z+wPSIxCgvksyDllyiDTCSbyOqz6g+0tkq9TSoL3WLkD7toxO5Z5b65w6NGaLBQ
Ly3P+nEbT4K7yprtDUyQv461c1QjruzFTVYh8cTyBsC9ijmFRcVhxfC/Y5GS3Itf
qEV25GIqDcz+iEYVluxDmqswdiy1MTY7qtFood7fxOAYLNrb6Rez/Tmesqf8Hd9B
thpq+xmJKeuSP5SyJwwh2kBcILhdwc9F3cyVZhXdgo0lSSmpWLMw+SzYe82+Fz3T
iKoXl9Y4vQvI2vkh0ccVR38WHWUXzNpvei79z2ck0/WFOSAk+RyjhP12npJGicCB
XDYCIrSoHNA/Rgp+IMcn9OYb6NmUGIJjkurTpsZe9AVN8L6Dq4LN655xL62HSic8
m72WrLBKRmfPWBtlEuAMkoawcKquGUMh3vOa9TLnDW6eXWKAiUDEtxG+BCdrtHcm
tCT8iVjJwj/+rMbx/wODR9CNsuwqPm6FZjMRWtbkz8MHxKzBKMRUDIiuhosCVLDB
8VuHD87nZcBgDNHB3VbCjwDon15uAvT2dT+lwv69G/2BiASEMmnTm2ZCJeziAr0s
DSYuMUQ6+GK0QlJ3NIG2VtgnV7pwRT9zSIrR52wfQykWq+3m2jnjDzNIemMg3Vnx
bjAJuNJKnb388v9KOKGGATvMo4TLf1bvj1FGHhmWPZg1FaGRdFc8S+JEcw6XIdUS
4RLk38DP6DazxWLH+wD2FNEMc165R1g7GnoGgU/5Xs92YUCdbX24U2aSeJGIOFAA
JCGX8VEtkFCko9cSEiKGoi3MWJZ18qYp+ZNoutNWlu3jX4ucSNw4/C1bxN7smsYY
ptJsNWFWOXs/2Q/HDw7NOuqiuQKanBeQVFeUoh4vxTugWMOa3GrcGed+y6ZVTDUw
s9v1RvA5TCT9J8TLr3DHsoyHRDWLzDGhJA3QJZAYXxubCJScpjqj1XsMzGyUxPDz
eRFJHUqn1+SwbmOweMfXJKQB0egicHXeCN6eXG00IcnoxFTRS64Qzbo4HXyI7Exf
mq6eHEuECn8bfZeYX+4D/M/rWsHrDjQOlEFSyWi5vxlkXzu1mP9kmVjL3cEbvw2G
ZV1jvBa8ptR8PcQdG9pxujC3DVXxpV+JLeUO8K2aGn+nh93cfQe2Phaj42N25pW8
XKwZY5pYXYuVHXw/ygfD05b4Oe5XsWQmbsn4hQpojQKqpruBDw6H9M0ScumDf++0
a6FXnYnEyu3juyesrGD0CC00hag24cqi5lUK4kicHHeagfvXaUasfG2D4Ae3PvZW
BvE+nbgWYHKx18pNrqLiaIFLcNd9AJSTAu6orOMVfuZ+SAK0QrEt6GquO/orWbFz
gKnqsXU7SVQJfVx3zS16HopIJ2Aaotqw4sdXsFzmO8ev7wq0zaKmHW61FxEtStCi
HzNkX6/B0qhD5R1q9shRcP27Hhaksw9cYk+EO4R6FbjDXIHxMYQetT+4IemAJQrR
NDqSO9gyGh1uiP7oFynd6RidZBpH8aCU9um1A51BQkz4qmnbpLoS5apiiFRHFdNn
VGUCW6fLkSfK8Ta0mmleRQSsmM8LsLgH2kEFojDv65HVjK22ctir2RWwG5NNKiho
jMlovbXUlf1HZQM4sE6m59mRD9OPLGDa+awLAYaclf68Zdd5Uz78gXZDYGuxtQ7g
xLbQu98Gy1UEeK7Bfd3TIzMSunRBt/h1VMsYt7s6keahgF7455nU/v2oVJK+VJyf
P0htadXLUvina8FY6p2ILq6DIDV/N0voJVp4F0XAd1+PYfyPX65Zqu4WGl9+pGtA
HlR2xJo33mfco2ghkR20x963hsjrB/dZAKUWi+iOs5VPQ5UoTHn5B+arewX9PLO0
Dm59ztw+HvXziAn5VgzWEntwPfQRnyEQXfmF7tKmGRfdBKzKUC469HH1uXC04fdN
qBtFWlwc81qeRzb02+qNXfaj3Hg9FoAo4akRt9NARLy5Hqf8iQeeH56RHqOtjl4J
MPPQ7lnL6Pwd/UXBDzN5OU6eURAWuypkJMczDZI+STbWAdBUk2vHy50B59V3wx2w
eP0rEISiUuzKcypjUHwPg9UGNTCkHF4WaHVdh0Fq/mGIMEoac+e965oYd4kG56Ph
qpCyBnuBqh4GfmoBhDBvzOAWgrHwpXudY1rdPAyVaGxhj4tbYuQd3gl8WfORQIb4
r7yQG1bp9610sJzFKkztFUntGIrQVOGgw1rR+i/Hzx2brFTMRxRfsfWsSIqcFtxc
OdeXxVUZV6ttnkPE9CZDrpgj4O2dEac6wnjX1zdw5DGdRKKsKvReejrCKGBGNzEx
JTKQIiVng/5NC6aTCzrpUgnIliNPfjSt25JCeCA7vXRh0A2KLNdHu0fjs7WXkyv+
1LccCXGkJuKDOHvMImwWHfVLx7yykYv2ncEvhqfKo5j1toVecnJi/7leOVlYraTp
dMvqqdj3/67SmjQh2IkOPt3zcrAEgnKbMjxiuQkGmUnotzJh/6x2FjQS2iR3pNiw
5JgoGQrqNhjnms34hYd/Ana5Z91+daoSTiTQAd5J4yADE4AhXLwTwZKnQ/ZIqxeG
Lu9UYBlquEVX81YHYux85lDn6sxcWkUnB3HBh7oNN4RuZ5WHDR5qfSxZy7iGchrW
MOmG6xzYwlq0Tyg/WJ/T1RmgsYmxfNSFKlog2cxSXIb0KD6F5v1ZBU/5Yw9f3JTM
4FWmNXelnwRrchOM8zFjAqmGuqOEz84eqMjB2ped7IRX22tmYeZi8vxlG7o3Rr3Q
NCAnDmrf1wEY9oIgUY47caNokpvtht893xaLtOeZSaGYkFird4ovMMpST/jBmSym
tA9LiDeepwayvcbiJkBUFtBKrp9nM8NcDMjL6vM9weuTI4Buq6RlkZnT8t0Wut45
biCus6i3DCM1eOb5PdDCrjZbZdaTJSqLBzT/yTEofi+fOv/GteAbePDDoazdsbIf
Z1OkyR+e2svMPyZpHN363Dan38mZphminROURAkyROOpr673OIq6wMi5A7r9XIYn
AdU2la3DwxFhG6pYF8sFRyMRECTZf4EV1NMing/8R/qLO7c59dEcBsl3gnrijFyd
nHiciMIJ/j0o3D9KU1dL5EmmciIrHZ5aB55vu/ibEik2pY/i/+xSRE4oir8+RSim
TsVCJpv/HCgo5yNVHqLxAOo5cVcroN4p1v0H7VXaif67pemdyOsgksGipYgHEVTq
tUFoYyxPef76t+22BM6pM0b5XOGBT7zN+7JtjRmaun71eKxaeOfHC0oJjAdGAlU5
61HI3c5gltf7docpgzL7yueDZ9/+M6ej5CAKwfAd1WpYY9vtmwxNRlOTBujv++nk
FP3eTL40sHPNKI78jldNi5YveA8lcidWSvCGNqbM52T1N8EhVoTuJ55F429CTWX5
MyHOo79viBTK3e2+mxhMVZsovEzqM6KQyUoJTNvtSjxEadKvJmXiiMcmY/YKRR6I
iPyxug/2XOyci+YldQNs0CNl9rNYXEnvJIVYNgkoe/oGLTqOCzUvtF8lsopzPXpE
eb3vutOClI+mp4Jb+LW4LFwS8J2iHbBqP97P3Fdez42UhKudQiGHL9joymL3oQeu
Qdtcrg05gc9znr/Dh2xhO3O5Kxu8OfTJxLzUVnKI1A9G1Ccmwb+WM6MeG4LdEgAK
gbevhdokICsEHY2Wt3cUVQP9YNguEc1tvk7mpt1XCfnoejyv89HnH6t1CAMD2OoT
If7WDccp8mEdytkvmKSDKRVftIxHaB/yudf0GVUZFcHL+2tXsNO0ricNfjvNSCaT
2IFYXiEs3UoBMNL6oGqzwLtDz2YgXQUEXDunCCeT4QN4m5VSCFdtbEbzFPO3xVUD
fLi1BrwaiReEWOeroGU54+S9IEB81LRyV32xMuUdvPWV0tLY6fCjzREqF90BZhVp
BHCYQSjOAP3YEHEBdBkQbRkAS/Mqt5lJvAaq0EBEas2E1+3zR4KfwEwXByv9T9zb
QtcxhzoU2sotVgNbehziaGLvFDQ9d1YAKOYxpwiW/4guf0qFIR/kw6DM+/uioblj
b6g68CFBMsQF/iNTxqLtVVRepu1AHmpcfPY22SSJxiMI7lI0Q76o+rJ5HLYEPkko
4Sw5HwmJr/nEt2eFWDC1fDrEoWZ7RmVHWjwLrwJ9GXJjqAEDpqwmCWDisxb3YV3P
uD+Q/4fzgI1IeyG2DlR7Paa+57bQTNBNNUhrzyXiArQI5zQAYDN8Grud6knXtQ3J
6h6AKeyCZ9iJgzGSIszmt+kRxQdHIsJAnsX/wFmRvTvWKDGHvsc01Wyt823q8pf2
L3Ym/98juxdH5rxRge+p4Uynsra7oQvevMFDVvBhu0362KL2ZLfpoZ/C1izr06h5
GJC9M4RpLjT25bhs6SSqfMCp1IXt/hSGzxtBx3Ghtv8Y/lMRml5RfUsdX1c7IYz9
TUuzdNHjDRqnF09ZGOQtaxC2ND50zIFXTGqxsWNYRpaM7LrREIxzNcIDNd/tGEJQ
H57mglSbgMAKRjgYmBFTwyJG4RiXTqwtOyj7kpQj2Up69XWxYe1CxRtwAOgaLpQv
qYr9ubgOIsE8XaHGu3IrkHLuE5Q+oJwZgPoGGNoxZyc21WnVRoq4/tQdDgiTNUhQ
6W5KFurnvL9GcZzAQpj16VYMl2eJiwLnOqQrU7qLiqCcIPp7iMDwtE2sOWLfF4y+
00ocizp5A4byBL/41R5LHgch0x6OXwDbL2ChXNXjPggG5Z5Myzc0dnP5bCDD21lS
mqUNNRk9g6djLf4GEgKhUo8rboIqnksg4J3nJPMsegGMEHJzd9FIGAiDOZ76MeqM
zRd3K9L54V2SgcMTMyHQauiiUZfAsfRMXmkX6bcDkVINoFSFb5OdNE45O6z/x2vZ
u1v2U/SSZThGajKNUIRuXLjxAYtOq1J1mXZUOY6JcRNTVwekloCMtruRoCOXGZ7E
qo7GW9nHCBurHZP30tewvCySx2eomLM0hnMEPlOXwTmTmck/cHjFCUYc0WbyNF7z
Xj8RuyP3z1fZZ75RSg8AtQDa9VPHS0bcW4tS86s5N+2wGlLLHjEcz9CdO8NWwvg1
SNSDnCVvYKFbUnbgCbF3pSEIpKdMxN2ltUJvorrs2qB2AIN7KgssQUpyFGxVhI1N
ydsPVURiEswhfLsIcTeZagz8JkQE13TgFY7WF+LVN/nYv7nbyHMcIsEJxzNBbxCS
TWxrDqxv7X7L/2NnIJuDNMyleB+8iO+4XbgHbQydsCrg4abC4/QN05LqtjSJMmEz
0Pg/kQJ0FO0dIvSX7uhSI5MBENPNgi9WQnh/ph3JkaybEl3YWgQ5yE3L2aI1XCRu
9Fx/ZAUXlSqlrWCzq9c5MQAzzJ6/28JnFG9Z81KhqDJixXSvt/H/hp1Zc+1SavkZ
GAE/+0eGS955bXO2a92ReOUj4SH39cn63i9WN4L4P9adsSPafVpAwZYaZiRJ5LDc
An34CW9E4WmwpFTZkg09cNZX92faaBqNrLgu2ELBKzcwIUkoC1Y4jepkVqN3N0Pp
FjerBjXXFsXFmtdvj/W9hN7NNGVO1IMeX0L2T6G7yatCEpXLCkCXc9iRofCvD601
jXbgVNlD6VKwYjuHXTOFe4Jw244mqHpFg6RDA8zhFbuJUs5oAqfq4nQ7PPLXuXDm
Hn1C2rSl+QoSuRstS1wvsjNsjIMo1VB9X2VmOVAyRU09iesHEWu2Tz9HqEsUIgCM
zl1NHRAowdA0Y3L0lzivo+nnxB2SC0O1hSFOcL0gqa/8HSv/CNeH3i9iMwxl+28f
eGH3em/5DEylcRfPcxA/q3re+i+PgJNzddo/9rsF1cyDWZr5Eo70Mg4PfzcEQTCB
5IfTjM7YCy1HXhCBvMVlFTav5MQpQzU/+L6FetznR/Wxjht65XsKAwV+7uz777Ud
rG6+9g9ehcQ2wJ6up1MxA7Q6voyzvCJKYzrq9F4qY7amZnlxKYYRvBY63st3j1Xf
h0OhylRC1lIepU5ruXkEKcuSR20OPxAKq1MeTkilqF1OTeIbw2lZHA2Lw8vipZUf
qBUDNZ39tDKeVrVtj1ykCHY+A6lZJn1A9wDbVXy15K4tmg4exo1oM1pblZQOfjgj
KMlYngwhgZYCVMcmpsaMTZTvB5PzTgSewDoK24oJR6tADjgAYNrlK5TOfE5/Dwxl
/lnjshK16V3AVC4IX0jHUt2ZfADGKPjS3aMY5GRknZ+SvK6ssK1pPg/wF46cD83e
pZgm4uETsHZRwdmmupljFnZFW9QH6dB4WgYubOBsAbjTWTHvCNIDxLMqxCGxgfZI
v0F1xK0pTRsspqhjnKuhB6fDuuCMzlHaIfWMSHeNLfLmE6Q3G0nhy3eAVRjlwyFH
Bokd5R/dzo7AqucsctVOeJJh1pEZGdETTzOm9x7fL90UIt7BQrcsCdxFB6PrhI31
ocCfFJg0lIjX2Qg21nqUz4dLqi+OhqoxVGxD8jbsfSut+IYVTY3NLxo2mVEof9G2
Qd8Lx1SckeDu5KezF6ZFVNSMp7ZQVZDfxMUztl1a+30tTb+7av2fODZM4iTF98GZ
LzZmGM8Ct4FoLwCkbQNtAmkUkctZ3qUq7zGq/p8849gBhd7NCqGCb30WWNqDKEue
9p+k3XduVFGyMJCrbQ2v7/lY76f8zPT8WDWfp9kQalp81iobIzEP5yMoFnoTaIbj
lOLp8oQC+CLa8H6MyE/7UakXg8rthwjb3WCNeC8wikRSyXF5x4MggQdYMxhEwefb
k3Cz1VGRFzVUZOnQAt51TIb6o+aEWGRFU/v/V98gZwcfIXdY61Z2+9wBLJaceSZN
Rwh25nG4YIV1AXrdf1bMh/9fp91IAZEGCMrZRia9nhhed+0ESxVoVswgppduuGhB
3evvHaKloyYyUBeHVIN5rf9kM1NZrnV9n9582CLr+wXgZTpUH60BLQnb9eY6SYMR
7nhCKTe7KM6jtkN+KM8Z4dG2/VBdcvQhVLXwYl5N8EnwkmuTDY3FSb2AQNMKeY0x
CWKyAOVZHUeIxRVKVtvbf5ZY0kuKubhezEfV5cjsA8WqdRL9kwlEcdthAxySk4Ep
S32Kktdtuyh61ih91/QTA1gi8owQf9Brfr/PcuK0qbVANBtG+BwDwRIBIvCMpLkW
dKFwlcCUYKx322iEZOCvOBwVENFalJqHuiEeqkezxVaFUmaJpXqP7k341k5aUO6/
Zllj3UYQmhWs3M0xqYC3OaaTXCe+3w8J15xf4ucGGDjHTcYsSQ5qNYpz7asLhAzg
J1AIUARacqD5kciCeXKnwOi4gK0UVJAzNxbn93HCl1eXTv+j8SdW/fFCrsqAGvVV
E7+y83cdna9mDc9frb0ljJisNOEQDVLpINFH3owxFEV5nmjb0U4Ca+m5pQJ7EuMI
JIl3Trbf9bdNCh9TRq7r8/i5Dr8r7elt5CoesIAPERw3JqKeJ7ea6kyd6isfsofb
frviTNkaATmPRcFXDcL8HxyJWCu4wEJSE2x4/Z6PpyC9j8aYI7IdpUiWjc5BoUEb
6m6BNqY3Wv0CuypsAR8zL62NoIWD2f8S3pC+TvTNzUO4urLUc1eeNpEtsOQ0nWpI
CYYTUrhYEjnFDLsjFfq3cXhNXbyQ+Aq/fooDB0y00Lu56achZy1pxoHCoBVt9QX/
oGxEN+JPpbdhMCxqtHGLMiByunY2aVRsJdOw/lx1142MgyEtSEJaw90Ya3Gv8oQ1
JadT/6No0VqqIpUSi66OkD6unf3Vrgwn4cl+yZZ5xXRKGFjYb1HkZn5+cXebFCmm
gD7lcCcFjti9Mw0Qarc8PAG4a9k1WAygpXDZRINb2lFvLiRBMZ9H0SbfBDiMisZk
39ht9VQaIuQDF/yTAi1xy6BaAmONI2nLQFkziGRCUrwclMQ4rZtW/Mx6XZzWhche
CWn8dJj7iAa0Fh/hbM5xxG0bPg92Dg/DUGpdc5L9DuCpfXFmETEZ81J0zlOZGY0Y
qBAwTCuDCmbrf5+GosNCSfu5dty+U2mB7RNHBMwht5zceNAVr/VysSxjXuuTAfgx
FStrjwG/0RgBa1Bc8AFC93qvMxTlRyEcB0Q5ss8vyAKCDJHhWpfxaWXwmiW8OwHG
WdtVgLVtkANl+4oDUzFfUVjg0NIixxtkCp0oj7/zgu+o8HeuNHrSKH/bYahU2g9R
UnTJQz9UEpYGpt7FLWfB7ef3K25oQu7J2KUWA7pmSx0CLOZtt4VUd7zlEUhVc5gr
gHYbLkZlG9PNjXFI+dKm8WW3MIMLgEFTS8/zRbX6ainZ4LRr+y4HOl28/VlAkEkl
XUhi3JOi9OiHdDGRnNcl8mX2jAydSfZi3zXCAmxRC9z2vXNDHOePuWKu1s2ucutk
hU+WhLdnOIrAVDo8GCalSXBxCIxh+/d18qGm90Y5+9WyzvsBBtCNaz50tcEi89xx
OrMqw35hLCVxcTyhndYNEQV+h0pbv5b8HPePXH5mtZiaxQ29uP3Lg8UZL1lC0xLz
LdjV+Xf92b/c4IyKeRdp4hhQifBedIkuNwcMBZgWGtEj9t8rrUPuPopQUDKR9Ysy
R23BbC54b29wb1Ctkie255WRtv+hysu9mjWHovZvL0AFoFdbhGuW8rqm7+/YmGZ8
ERLwlaObwXX6NECqiB1NaKVy0A2Y+EuHG5Q89RisClTa3acCHMl4V2WNIEw+eZX3
TmIms0Cmtj/4SNwzZwDuSjY65Xqpc4CMzAo6/qG8i0vfhk2P/RobOob933u7ozwV
av1Hu+epEs5ixXd7BvVpzptAwrupEV0bFrtN5IHBwS98IeaQkk2vtn5/fRUXJ+In
wLJ62MBVYtuDc+hmE3TKv/D2vcg5ewnrcVsj2KO5MiQa/6auiAOPU3ekcI47LU4l
QlLrb0Ch8eqGHCYcEvieJfzgVVdKSw1QzNbOJAIiLakofg+hx3/r2E2CFqUt1kIF
CGFxW2lGqM6q3A81EkbZ9c2coYVNrhIwreyCBZFP7JkxSDXKWRwS87PZt9Ubr25n
ecl+qVAK9AUOUC98gDtZ2OfVjoGN6sMo5PmE3Yvfq9/e6ILHzWElEaCw3Kk/bV/U
CwqYiHINU7+HYo26pufRaI74+y/ae/ud/sG7v1wv7QtquKc6cE2WXX3ax/NKERpk
aqp6JOZUKqawxM5ALz/jj9SXUILGv+6fjroBiyJdQ6QuxEkpmrAUYX1TC9HwnI3D
L+jLt2HSIqm/bV8v/FpmqPNV2wfzHqIEpHyQVqSJmo0xYsbw2wC2DhlaEyZkwbJh
OvBlOEWvISvJ2TUyHMvKFe1gFAo3c4N6VXFVVGCCgtmCFRC7WQoiu3CSas1K0t1j
9Md3r/TgHuLiId7aK3Fdnu4zsF3z5XJ93LVxQQw4KncfeCPM89prl9JtwFywnMXZ
kqUscYTpUIxYrr9rRczmIHGtsjgpFEqJ04Ji93xI4pkvf+CxovkMKwkLU/ayFc9o
tpsW1k2+g/uDm0CTv/diJgbRertWphaiwjHbiyEc0sINLCWDdyDFSiJeY9BN0x4x
xDOiX/rgqR0OFUKqLGrkXznH4jGYxQhO/73QLRfrkVzR3E5aosATmAgS0JhQX45Q
ORtgqYzz7EoHsPL+U6wZtR2UWTFi0EkmTD2wpngLHD5XdBMv7OJ4ewVsbHZ2tank
bxF19KwH6ZLBbwcGaHWdMf1DAI5kuXSJ5FQQgEgHkUhvzTHlRThlFgCVsPB2Ogjs
ZagpYEkYb0/0DIEi5Pn7n0rlXr1Npgkn/E45nAXmrOJdFS50R+VAZJ1KYtCxWvAI
YbDozRZjoPpNlBT+MDK528vxf53Ue9wFE2HfbUpqzzkv0aw+/+nStSB7wukB/RXT
2YGNCyCP1pDEFWXXAngyg9iqxig7ox99RwqYSIvysoctM11YVLNWOUsaFBJbIADU
+Xb73vDEC2MYNOUKsEGOtlSmoFBinx8ppIZYCYer64HZWks2W8gRIaCsqBvqIRRc
QBp086nHQBRgRJzPbjCn/s6F2uAIywUqlqUgu8sXz1+fi5ealtgxtOGHpmjLMSEY
agYUprxKWSSvrl6xcoQEeSy8fTeJm2lNAiFbiPI38nuQ4R/WeMHWMVMNwKWCIK5s
LT3TrRKCueTMXbKP+EOVxrbBiUadkuj7ykqeIk5B+SxXq/uk2Ksc2dKi+mF2J7jP
qPN4L15ejpCQI71ET/yjKPERKMBOD7RO/BOdOzddFu+DcBHcVkFZnJDQuNF6IGzw
KUprnZkakJoBvwfDbP5thOD51oUS2TKdDfTYVqw+FKG10OhUmU1AbdoSr+1cw7Vg
8lRfXrGuTOtUYpiFtXLAyy90Y01TI1s0styuVtHnSB8ye8hZrPIsFG6DeYoAfwWb
YlTZYxfhMk5D2Sop9mNOPceCGdMO+Rp+Yu1FSzmf4B/MJ3QIjRx9wlMtxcexJ3cu
KuVbdor3aw/+eQWt+L1uNt91kfft/A+Q2V0a1+Qs9MkGNTPsPGhQ0yFT5jYJrzZk
hQyz478q+78kMi0Yccd3Dctp+spKnkXLXDvJHa6/iPDO0AWq8EBxZAscJzyLf5Z5
AfNTDfBsbhg41rtYI7aNkTjgyvN0wrtVpfTULTgttTekFAppHaWsnCZKmcpvhDgs
gPyE9T4wqmkwkdFn4lkXlM7rrIahcTxuILgKsqJzVWYMmKtow8xy/D7WNu4f1fzV
7+3ZWY1DuGMspGeJOLfjM8xcyXrxehSpq+LQcgCOtPGpoci5Y7HsZ/JXxmdZhnXR
yQWnldwLau0ghEEEKiQ7SIaeLz2LUF/W34j3yNehjW2+UpWf1vceLMm5hHQtYz/2
TK0ijDjfk6pYlTAI+i5nUEbHHQE4uq/z5voHYk2uDhDYSMWM0bsv5tkwIyDi5zO8
nEqcE5kyGoHpJGiatywGthff3g+a7sHFWGGVIsNx5JKVFbE2HPlRIH48FYGCDgSh
FZHDI7YzT2t4bYjaUPHG0kdgb7hctQJ9vGMg4JYo7M9ltQN9E6Qa0fmWa7yUeuEh
WTYHmVyxDAV0sJzkzjCvxdx09dm4zKQ+PR4D2/AJ5lm9Q1jC+F1gWLJgZx2PrRZB
janng6IVL8QMjHKMo8Z3ukJcsrT98gFu8d+eUiv+AsvbEZpoPOkNrgNwY2hkpWs4
Vgoo1+QFbUdJ4dxmxXcRPQCwvod1nbKoV+/eItFZGPAUZCB6TLlCdQD1b92i9p+0
LoZVhE57sV7J3w49Ket4r7P2mM9h9hEY0k9LYCA2vDfQzNgNTkbvqwvTo8IiU6Zm
5d7p+J87EMLKfGA6cf8vAec6hWL5NyPKF9uBSkaBIbVY5SGYpYDR/adIYdzqYY1a
lJCm0mqRwSXORv+MIM/OoDoDkqBZWeK1ZkvYB5BcTbwdjNd7PHLXbj5j8AfB86BV
P/uVcZGoptr5G/23Zjxhd5S/rjFT8nztkRRE1hihbUsb2unX7VUBmfsl3PNrxY2c
I2rr78y1TIQkgN8KChDaa3S2FkWJQAIlH09qv3cCXIG9DbScqGRezg7cyejTBg2X
Iy4QR1WNWUDrjVoMMv3RWbm9JvUdkfGDlzZqD4NXmW5KqTI7JAyW4ly4i0KFZt9W
1IPkmYpROkZ2N+ewFJI1E4BvuQgl5MgAafgs5rEZBA6EPGeoisQl2wdTwZ9QKY05
gy0LnXANj5UZGT1ShS5i8VELY1q4wOksWWOGOcr44CgutsDLdoaYRJB5XpHA9kQR
YUIN8PJM7FS49uCRG23WvQk9Igzg2j//0FmKFbw18p+NcwhsrgjKVDdZSAbg/ZjU
gshpmQQwVYwg7JJ9AobPiQDXufmzEJz2kcynpkbBgYrutE+lC2JQzK2ZzIEZ1zSU
o/wwSOCZBn51vq+A6WhWsCbdsf/QNTLIvhCjemLz09H14tzCXzFmCUW7UGU8Boqb
dyg2ksnsJro0CeRFATfmku6Pu4CseCOL5t4sslTCV+e4fIo/A/xwqJssFkRhGIrg
fF/JDAb9GAsIa9jt4/rAmrWA+yS7k2TqXA4rT/70D80WRNplN3fG1oVYu49GL65J
D7s+ovCWYRaON3q9ew3Q8ZVHU4g9iIQvCaIAh6pv2RxgMYI7mpDmZchA67N1vECy
yo5aRuptBjWLTo4Mzu3BUrC/P/tXpw58SvF0ARJx2Y7DqwvZjeC6sHrN3lo/SdZx
PCN6OCNqEG09SmY1cfMu0naCGBws0o2A4pLlfpmoF5flinOSnQ8rI2t5E1Jg2VQ+
n/GZQqJ4aRP6gVd5HJbIwDcooH3tMK7Ynhm10G6NCINIR+47LcnoRbJ6LBC40Dp1
NoyhGOn3jHAslaPt89Z8Nb8BR8wXG5qNc94oIVVwZA7GerWRbvLZ9462G42Dg+No
EokzJuwHPNZ8MtV9VFDgVQTHC1FqyEWgWXJnMr+cntM5VervO1EEscfeLZ+u751L
foy3B4O+7hkh3mOGxXwttqGTYtc4L0RqdaB84xagXeirVKtFqPG3G7oeQlLqu4cc
HNH8on1aRHMZZqNXI47LFgTqjl8S06rrkLFm/lvPH+2Y2bk2ldHz+L3+kqQT1CcY
uLGaIcpt7UAVhegcfrPcyVEYQaGWGMvwwru6Fw9Ll5xY/Uhh9DlqplJGlVW2WjFu
niS1wSuFvuwMhgWa2Xdry2+SZs5xCyLWSiRRnDaaYoDNjrePhlFbS0EDrM6QFvOQ
2pWfY1LsnyDOxyQn68GTeNSb0DCAyGKzAHoIAIsYbXfiJKpH7dG4MOkBk7lI054V
Ba6aJRHUYgXqPsjWmUoTFGSn2BSAalweqJyE4T8MjFRDj5JHP77nqMYK6VB1I4Va
lHmyyMYGMO94P16HWSwJq+x4QJFqlip5Gl8scmvKUVOLD8IHQipRxOLrhdriMUEC
RlsUYd9HUfKJgH6PmFY2frqX4vf1XFSq6Ac7Ts8AzqoneE5BMHd4N4CS0Ro+xl8C
HmsqJIb+NmbllkMr+wt57R7luKqild3wW7eqeBbhS+xZi2DlmuvQZAb9tm+tbXKh
whdspXoZvkuDYB+5r8TIsff52ueFfNaDWwlp8f+yKeqIHJWH0WFa2oYjJAl/hwZo
pF5vdZNJOfbfz0Omx3JeqP9ZaeH2+NkOIpVqjQ+lQKvIUFqNcR5Ib+8FGZygSgZ5
Kc+VFvDgb19bUyx7IrkGMu2g6WUJZu/E0Yk0wRsCvZZSG1DqzWZZG35zye85fFP9
gNjEGTGy6VfJFh+V1aQ/YcSDc+cHKjMh1wrZi9xF6xf2hHF8FZ6DR/JJpQKe/5iY
V2Es2blIZX5sXM8sxt4GB4UXn76bax/t1NMt+H40KwgcYIrMr236JcD1NhwSZ/X+
U4wserIvPdiTH4jNyAuILzTtYaqYM1FBoKITiCe0usg=
`protect end_protected