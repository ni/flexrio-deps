`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6048 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
cIEcm3T3CtIEatkHUC/ntiwbDTx51UmRZLG1WpClOKD4OePIndij5cJVZ+8uR1X2
fGV7r8UtiI9h5qQTMM07+0WuY/gdslhCEyKADjjS6Tgjl5JojToDZdOdlfMJVD0m
tQ6W9cDtDCYpXtgcxTUQdbR0sxbnLPfiwd+zfzhv/UCLn7s7DBP2V03MfyuAqPcB
L7LYSgvcjUWjkR8r9Jcd9Ss6mJcw6C2xTKiFmJkJV8rVwI1fyRYP0P1w0IwI09gG
z1xouSCOzHyu9V8AX1bR5wbb6xXLB00YyMuC2neD6cS5ttv5l//JQmSJndJ4/keI
m+fElI1+0CigXzuMqYup+OxoYQvAtEJ8ZCwSLmViN0F6MmwKIfcNSHbby0uwEWZ7
rxm5aYJeEXbtCUkzEE8ZnRKEhuBjCVa3aap+BLrPuxmlow/uvesw1LmueGC+z1Qy
n55Awmo2aD3zf88CUNL1kl46wI4N6fy1haMb8USaVE3egMlW6tVL62PDc/zN+L+8
3Fx4IG2o6tWlNV0EWBKD8NGbsX89krKQ4tinK9wofBhFDePPEbwCgqt2Iw9mAEBc
IPwbgjL47lz332aaTNIipa/fw4CK3aCmXjpWOiYZTNdiG1AK8EGzwU1okpOtWiPp
0ZEPqXbHXz7GOAw8u+loB21acszNsDakdpfm8Z8nsZ3pccmqbHhfB4biJmEC4X2D
s2rqLZqgSlHpll74+iANUr5NS1k3FDG0dg2yzR/DZq93mcQ1sfUauSK2mHcgJqnF
Kk/LX3K6zvJu/p6XklD1CSQpJaKCKmWPCcvx0qkakCAF4Kq+mBbqkfxquaxkOAGw
WkkQYZxBfms16hvskhc6WFOInCl1JtaF6fjlME8owpzn4aRYizBnjEG9L4N0YGI3
iI2xbc/Bvd0xue4/ZHM+aS1ZAPgSsPXbtnV2ilUyBuoCV4c1gyEk0qnYe42R+CkA
Pict2vFkWTHrkG9l8uei8el0ShMXu0avPqNjS1s+xqY9xLkK1BGTKBXTc32WH+pl
pIGWWUwhD+474pDhAO3Yg+CHIW5UFP3x/Z88LoZRPb5+ri0nJPV0EDgK0JujQFtI
A556CCdjz/T0vA+MYE3JgcOtqJvSWsDXXNuTyzGdj1A+CH0Sk2O0qi7dPB3ocRdG
qv5FW/HMRpilM/bDBen1lU5mni0xklh1Y4k7ZbggMlhzllb+i2RCDbcz+f+XLgx7
bm900WryBA8/OAq4g8w1U/zOd0mUCktGT0w91dUh9WzWm5lF/TFk1Y9sOJHDZQG5
LrhIXkaPIu3/Pl67YFhG9jKxfCEVbzyw692UJGf5xVdkZImKyjVPdzh+QR91DRel
mxgs1Xv/+dvxzMNZzPpTy5Em61F47WpSWXlW27WSlqQlKzShpRU6f5zEK+zZS4wv
xxFrTyTFAZYAzsRxUrJ7rzl4RxbXccb5447fvYaPwmIOzFJqt5hgBWeOt3ZvjMts
tE96LGPsA/FH29+OqC9PoplcnHE4NLxZv5YeV0S4ZRy7/1Z4GQWlCZS6lw4lYL3p
3I6OC5SXLVjkBm75jy/QG0T1RLSppknRG6GjDPqxUu8hDqmUmI+X8sv5UWuEU9zd
JDPq9+MhbOzezONCOyZxMJElTwYUOm4DLx1Da1mgETMl1+tHdaNDOXw0swehYRWY
Sz6BDrFPx7t1Z80k1SN9vAAgq8WkuQcBBTIpzJWhNy3/NgfJj2Omd0ZgFIynuSXi
Bc3MLs7DTkDiLvLrHFwETIUzT2C1C2xKYHIAtudEQIr7s9uQXekinwqYkMnMMBU9
lBhcK7TuyHdMg4wj3bOhKaZCaWQo9hCQmJAy/wI6JRh9PYDArQPjrwQ7qTj85d6I
Xuauv98mwJsQBmiRIiD/dY6BdG69pH8Pq6SpEAI8ffoX6PX4jDHHwMDGn7R+jVGu
sTXG7DLxd2vlSln/gdUzTFCVCUMd1kfYLhTdByM8D7iUMICr5WHPYFu502rBI/ER
NMsgZZFYFMwx67XQrT8dzB5gmIlKGUnPyEdHMGbAgYbOBtYQYrVzQBa7LtFGm90S
qLPQrWby5+e4jWQkYOXt2aNaivOCC+7gREMOPipfDaI6o8/2fV6i1FOnCmMgsBMX
u/3OKyK2kAdHmcBxixZeQ8A6uKcgB4dw9or3eNlA/Pi/n6XEau05agfyPgrsdovf
HwtyHs+C2YbGpYr0L+bg5ZtooJOuI1svN8saRkdJIo+dZn3ZS8Bl9F8VocYLrzP3
aBsT5w0FRVXIjHMTdESyNr18PWdEu2H363HA1Ad3pMZEGoxgWt38Ej8X8q6hC5Z1
811bWGY6UQcGWlZ8NNMHm6vO5jUET0Qf5mwc+6P3eE5s3UU97BdUJ+vmEVHvpEGk
xsFAPNZYN7WhM03GeoNCoLSM0FG3mLPEwO0xjiHkIHWq0OD1DC3/FzZ0sNVrHqwY
GiK/QETFmxWr+/juLyQRPixSPCIEgfr+7uKdUPTq55AspmcDmrxA3D4giWsP1hqN
BZzZfbaNhvq7/yXIlh0Ynr+A0ncDR7n/An4ZlVoWMylJeGkT5ye6J7nhoXMF6Hif
+qZUFuh0q8V2F5wsVDmvGxp/YOGdfPB2rxJiYkRI0FoAK4mhiuYqKvhHqkHzuKEj
Jg1pI6uCF6Ryhk4iBtyBoiKu7cxvqFH92luPzVRCk4rpktp6wOFACF/QYmyXas6V
Boqxcsgx1BaUft9wsrflD1n4mndPJTCJrziY6k5NKeBTPGYUOjVrnvxc3e3uyT/2
KGc7yRYCadlWD5nkzJRiEoCFDlDrDC4O483Uwa8m6dPIh2JTO3Zs9Jd4UhiPJeAQ
PvihM1yoyhfMlZPp1cS6p5+ns/5v0Ep6rGeVbU+/D2erDmjXRwOaH++QWhaHh3A8
ZtMR+tKU2dWTfpum0RSRTHor5SUOHWryr3xKbtAeAggxgxcIMnoBGEbZgZQ7WVbP
KKYIaLhSBJW8BOI3vaUOX7ReEf0EdLyxzTNMCVO5X+Tj6WqvdfPqL/TLsQkw9+fu
MoxJA+cIWtWq5MSluUH7fc3r9BJFFgcqkwWbZS3r0zaxzbOVdxDsL1ziCnj/oVeI
QT6YIDJlh9flGslY2J94MBSyiMZulA7hTKuHz2VzVqLVfw9fvs7R6BOFqzEOI+N6
vRSB52hktFXgEfknUlpuFFdCJ7IZZcDduW0xcDB4PDQuNszfL9UkMRFuhkvBxVB7
pHJTDiEtynhDqE5RtAYCM9cI6mkXgT4qCINsJ1jZZN+P1TVwd9e7yIXBc9vqyz4s
vThm61Glkl6fBrAgRg+Rm8n7V72elDri6uDTRZlSHv6+m+U5N5EuumZ2qUYVvYH4
slSOUnZNAzJYMxWrPauOR526U/fRTg81uOaCpduJWZZruMAjtfaE8awrDfWO2OEY
z8idht5x4JxsQCSV7M47UA7D2LZgnZ5UBWLFMvC8ReRkr7GnsIEYKPnTc448VxPP
7X6/7zjS3JTItXhE90bSBhsufDORD+vEdkb9Q90aD4DrZjasTrFQzx5YmcCQ7skm
iuUoNTWxVvBc8uwn5LBwxxnJuJ1kxFa00jbERvLEghPFuz4+m0K35G+hVcGIoWBr
vSavq/kkzjVYQx9UCdX+mbmu0qj/1rTlGWP6L94+sD+MgO/XEoS8YBewo0uaA2Q8
Rkrv64vCBknNa13pbz5W++2aIJ8QGyRFO9g8Q3FnTK6/2v78ljTGZMxUxStfVhc6
Qx8pgeZ+S6146TZlTPozXwCbdnBVz1RfuZxzCXwHdIre/GbUkjlR8gUYg+0bpgzS
8s9QOwglYYrZ8V0I01s/ADCrDYyHcuEDSrClEXKHF4ybw4jEFJk1x7yk/EZIxYAT
207mxm2oF9yFohsT7FduRcXwwQFjp7iK/jc5doFyExL7lsmYm5XBaY096THDPKnJ
+lWpL4uzlIiVtDb4DXkMJkD+dgShBFtR1/1JL2rAE4kqdrNvdyp6YksPZiOHMISx
7NRMuZun+fTkwax955rEg9oksfR7pScsqHjvYpiu8L37p5JRI91OMT8vYfPJyd3+
4rn5QqQlfwzGivQuM9oNARVYAKESKqWOUePcpxCwhcQsubbjZ5Jx8tqeoZo4YFx0
xl0uLj5HnSBiM7m/KKoDaPaMdcdRhTym4ncQYN+8Zmk79miF6NGiSO07LomgMZ4e
q/wQkwGKEeVJ1YjdnjAyxAPzR2YoF4XHxxTiLgokrhr4/RfNI5SMu+8GoKNnQPGP
8By+ZvgfZpIoxaRm7Y5/BiUKaksaHbN7ZXMk6vDdzvx9XWD5Li8Ux8pKAi4ojnry
/9Kl9YOwMucvBC7arFEgH9fVVx2CYVLlgargIK5Jvm2cBswiDmFPJ82D5kgJ/Z3s
1WgSo3ntP3iu274wiBh/djUhpdLLII8AgLVOX/cBlX3kPdQVJwE06xsG3FXiDpk4
XCVdGFAGudqihrxXVUIS2s0nsNn4Gh7xgAI3vH/V0o2Xn10XHZ4lAMYmAcjoJv5e
c+nO97PdtpGb0Poh9LaO3U/goTnCvyS5aREp1D4M58Eqr52uLwWyYP8u4bMwvpWv
DOAn4tgBx2NuJJ6s8yKZ+pWYdg2X5TFxKr2gs+Waxj573Hyu+Ifj/trzi3TIXzqc
B2FXrMWKH3DZGUBw49W5nT5rW3tUDqZB2XUKsVdLG69iUQHUe7ln5u9LdhUKcC+v
SP+aoztO9CG+Mb2WamRcTkuNxGFjRpfdVIm87YBkIz+l/pQQOyXTL734Rp4XTEqZ
srazvRAxUtVtJna/W17CRNh3958hj1PySfSTYbY31duwGKulrkjeQ9ExTver0TuN
/ff4Y5DiyWfCzMeFPD89lQKDT2FyFaOCIhD6ZHl7i0dZBAfCI6uz5qB1RM0mXn8G
HHx9x5aLDRCn2ph9FNW5gnZ/oaO1HTvXAhp2FKNxEVrEw+o/dI/ubwQRNW9ZOJC/
KZEs3T8yOLpJZfgY1O4ADiLxYtgYttDgsohDl1jsBfGEwoSeC2ysAUfx56YKQddm
B19E+N69AMwdgpwzNkE8sgea4w9oy1En4XmJrS9rjHkq290DroFGK8EKN885E/bs
iqlk6PKWcutr6vnNSam68hWGPPjsymAUG1wL+a0OOyhVrexCZAyYSFBafiVhCzVD
zuIshUdQSvljFF8qO8QnEAwvl8p3qObc5HO7NnnYlipeIWWC6yrpQVmLOoaIx0Oy
aikTU07umIwhjPzLWS5XclFhnR+Ucj5L7oO8yNTEtE/245P7TvLySFWiJg1mQ/Z1
P50c4+lbOPCzTwQOCqxlRk7Sc+gFMs9FqU91xCWCTZaDzt8UZ3yF1eKA2KYuBcgd
JTGUuxgaO0oXSQ4ogpywTmIYPTA1BR/Ma0KPPeAHjv606PcPB7ClqqapPriwZYPw
EEN36pY2lNCfCPcmg6OSR6ojSAHN3hoJPTFPZFbDCGRqxekm+Zpt4r7BjyAF6pvs
3NrV2JDV70tFbMhRf0DH5UXow7rnwRbdPtscpDIkOCBuOqtfIGsUpqDpj+Q9cG9D
in3tH0dC0kuzd5rT7S4QK6okOrdixcH4+IjQD068tMXV5mMNeEo4gWcKUQBqzJ92
BDcf/FhJ/2ajlboipU24hWdty2rHtAyFHymNGhOE4USFYpUIIDEYBHeOMqgjOM1L
mKnwNqtl8tPGQQIWusEmRvd4XvvV2HaTDpEMHtLZ81ZQlXmZJORYYyfPIK1nnuQ5
+AieCRgFb3ZFGvOBVR/v+bbmFpFtZ8ob26qhT5oGPjXNawmgNZbMER9Fw3EYBhFA
45FX3ptRlshoijP1tKQpjvxKZMJaNRfydL3O3+lmtALE6N29LUkaDOIY11t7AlzX
b0iGZm3io8jUPYw4v1fonMPgXD08sR1CmpK5AYlYWHcX04HMyjdFnTX9R4JGYp3r
ZySx7yqJ8/kqr+SITh00dymhtunBYtHopReMfsRJaNv5NhXftBu+lUMezGHbBcGf
wJllBaYkRY2jYWqFwy/TO8x+UCV4vVzmdhI9RzG2//QBvNMiTA4aWPObP8XhSQBK
wbdmeXMmF9znowcfouwEu/L/O2h8NC4yEyp9p2U1AZuAsudlewcuivDzuG6CteJ4
dzj+S1eOUNKDgS1y0Vfh8c/2F/4ApETbUFz7LuepKe4Dympsbtq0VA6B4rtF2aBc
+EtSPzrBACzhFYB1oh1pw+h+CFmdY3b0Vs5CMPH+txIdlK+SxwpBxLaT9ZmNf//9
XCfg0fwsy7b18b5x0idZbsuf8rdO7cK6UDjuut8V0z5kWng88JTRnfzqHgjdPpVT
VTXwG3UU7BT1ESLci2p7ZWHC6m4EGJVB07mQXqlbQ0NeN4FEKorp/9MUxA+mJPTj
vlKGhXlEYMjb5gEmir9AfxUhXnO15fT4vgzyFR2c1zb8yuhVsnJ7bzSvoja54KMP
+rO+G7EnR+wAzk0jloGKjmjuUgpLZlboKNFUJDh697bLR6HcSanvPoCW1XFvmxvU
oUxONm73CJmsXevLgDPbiEVjwT9pCa8wbsycfCSNRaHheqpzCesJimSnTKIovFF6
2GVcl/Y3THUWT4yZ8gf1MqEDksRXjWoNSDl/jkJ+zBcryjXTjPpfBaAjlFw9z+x2
afAliKXgfdquT/A9vpMyMtOQfnqhM8e0mLHm/RD6Nt9Js8DiRvjU7OHJgJljztwd
RSjNp/dUZx88Bpl5ZNxAf6VtKbzSXAsELU0LkyfbqroFDakfsxWJSgCXWRGA4OSi
O89OnCM3FeJ2Haindgvh2cOM2ST949KkOHDXW6AyvhOnuy+e8ZpZAs6no1hq7A0B
/G+pMJE5dIL+CpQ+qTxnLQx8RXrK92usYFgNTZ5DoKFJRzcXW9xzOdBqVJjJfWKa
f4bPD3rN1ko3gxRTm/VCnBZYRoVFHa+qFBuS8B87EfSeB6tP01wbmqZ6hryhZdC6
/TaQSJHvQUK58PfoVWSOGLh4YQRyOP67DeYq81R7bqModnK18UzdRUpF9SvGzDiQ
0dgdLBUxlbj5EZhQpKDtIosMsraPUJWOgDdQtHYMCzamIUXVRlzW5nvC7Xeqc40w
FF5OCpMj343PgVW/ll6Mvkfs/HDxJmBaka8ZMIFt3pGCtS1H+HR0rXg3Sm66Wy3A
/fmU4llGZ5dPKnObvGPg0wY/TDm6HhMZ1lkputACZBVSrkFHZMafn1cO6wY4d/ya
S3jHQDk8VZuvS5Nt4PAXaN0GyzUgZ2XffN5qfsts+/fgjQ1dJuuUciudTuw4EdwX
FZDZDit9LjhDPBpRqFvsaVBOqFgVkHj9FYaHxOhNIiP13ZjJ4myCROmD6pJKQqlM
2juCq2mudKqywpBXZdAjuvz32H15KVDcRCLvvBciq2ugtYqyX+WvbPk8LkAxYcNl
58P9YATyh9dQUgfl2HRpf+LRiYdwEwYH5WYIpbPMWvoEByqK0TDEnpup+XnlJQL1
BbXYEvVp2zb60odypfrx6tIZMJWdKq1p2ocKYNDal8S+ktnX5Z2RcZjeeYeY+XRM
uzwUfawE/6ezgBAd1+UvZm4vQVgf2ErkrXaMT41ilhAO7Iu70xCe+QlEYrzIBD2o
Xnfo1oOAxnF1aQAQpz5iPrrWqjRi7bJlbFPQJ/34rlh+/VO7Ng6AxqDbp4uMmukG
Zdv+9jnmeoL4MRZUxgMkm/RexWoe8wLdcerFLwjpPReY45umytI7ko3dnAsnSQUq
KBtPUHKKQ+0seKiiWNdivFRdbf2g2WX0WV5adKIE9iENhT7d3wPxkF+SJQrxx6Hj
Wu8IVmFKNwzxWa3VF71kJ4xdqgHFmTujt6jEwGRStj7JSkvJocgeqU/j2eZQ5d8D
+19UrTxz6WBD9tPJ4pXAfsIOwhUlOfFbnhHAvqTEyRTZnLAPQVef1NpNoZCjh9fL
PjQi/datTGvi9UwWLiGoT+qnbJ6TFLnuIPJhQQHpTqsXRjpZdk3kqa8fjhHsU3GG
`protect end_protected