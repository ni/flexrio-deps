`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 33072 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
HDP29p0vLOrNPcWDOvry+eDDmy9r/VB01AA/OuRIVl74oUI9yLRb1tRgr+z/gwfZ
9eDTdEka6zD44Mm/0j1/YW+pHRfYCU0gv0gzva7hfH00UtwrLXteVadlfUrlA4le
pEcnBlAQD8depzwqB2CaDmE9rCUR/owRI4OKj2VvJsdv76qurFFG3Bz7DsamrTQY
XsmzVh9vu4CZKyNHWc35LvikO0brqbNBFbuzCIAhLeAAlG7hlcU35DU8WqHO5Wz1
io9uoyudNAOoDUJnd5YpgSnKwQYRt/d1UTVPh5M4dOgMxo7n6OyL56K8W0NqqcUg
LxU6euq4n0mlq8oL9aanT1BH52LXsvU65fZt9CCOKfmxahP/vqrhjlxYRisuXtjk
pF3ECQ7MTShVLGqCsobjAYw3pvtLjbQcjAj6voADoDkHNdbmJwsxsImgLeK8IRic
nxu7bfdWZ0VUK0xVh11nSwGiL13U1j087Oreadm0isO7FwWa8n1KTYZ9iSSMgMwD
iy0oqNn50WkBWa4kO6ry/9+uwoAhD9ETX7bkw+WP0rOzK3MOfBU2LsylpUUMoDwR
oRDWupMlKNdUR3GWGGbxkTKtX0wEqwUTaNvZRx7yCk4Q9gM2grdOVN0zFQRFy5OS
x+8D78tLD2PgV1ngbzx/vlMbTcpu7vUwaD5fAWM6ieJKPq2DyqdRiEvcGTtnhBlN
zYfIQRD1/CsF2rPNfOGSbMIx/SXY/QLVRIHxfuZ1vpLcuQG3s9xeW/4vsjffwnYo
ebL01l0zbMu8rfae3lS5a7tLaj3KyEgVxjKTTXpffa88mPeQrEoSynRHfyF/tbGd
sEJ5bxkvfDviAg4FWZb8DaP2qbGK7x1dqeQBJM/gMMPWd2zfvHETxDE6odPliwu2
fr9FMRgVq/rvbiNO7neX6c8mfy3ndexvsBRmMbPojuQJ1+as+XegSmg8HPqnqhHU
DMkvEtBJjhG+HHMgVhr8bFDZZ6VqxcG1lcrKYneG+iDAZz5uDIMxs9Lo+uCVuSXI
q6w5TL4+bxo+4u0EAQk23GjR3cMCHkFvpGnxzG7Rq++jIPMVIULqcONfjbqI2I3L
2w60sf93BEJdnjVUVYsUZnIHDexLgcdH08PT7xnbVjK7n/VTCMpgahZHZ9lh1xeB
zwb2Cd4MtC59ZbYsK7HcU0zrqSOpNL0FJABAqdY4VjbVp/q4Txc1CmO+H45Ktk8Q
dQx72+jPOXTW7pMukNC5YWuxKN5DZQw0whizlxR/BTqtdxZ2HHZLGRAqSvhdKqTD
67A6KdRYRAGiIZBngozAYyRp4QBr/ehvae6g3f+JxifeW2dWvutVP/aIeqUU4eQg
cGLK7REUkBqaHVE57597txOiYKCYOuh6k0EKnW+O68jqHKdcwAxaZlsg4bvCFLxu
wkfg7nn6ksVEp1815IZaBozr72PLaQkHdJFjdh9tBudVSjp7c1nzokLRDvuKRj+Y
SjUbc/yevJdKXdpPa9na9MOieceaz+OyrfYDqaqKiYI5rlp6UuU4GuCzNX+pRghn
Xou/b26DgA5VVOLLFXslrOoJQ+raAoUG/PdjhSwhbDr8bJQdFYlcnfrh0d3H3URb
AJ25WEBjturrKnpUWm2XYvwi4Y6eJPMbb31xDx000yQbFYtWDqBKr7uhDKmW/H/h
VwHUCeGVf/YadSB4s5L6kIsYmxAgTJ/jJwNlMSl50EjSqWVmtdYuDt/qFBWuXzHF
8u78M2f/OifIVDKXfIg4PO6B7X2FHG7xlviaidNULRP8roXY/Cqp/7aLdPjRL48q
P0PWzFUUsE3V3seUwwmtqPq3/RDCOIvmQ8+rmHnLkFXPcX3tlVyPh/Xro8vk6d8w
u9Pr+1kXTqQKYMo/+Rn7WWL5IUkV8IGgGCfn4OVz0Bm/TNYdxGisop73mtvrqg03
2+UQ4pPccCrWNxs7mR9LxoFTE69MMdV5IvfvNX9yuhcjq7OJrDcEG0hNZhDsUa72
atXEwheo+B2Ism+d/io88IRJQxyiKSSezn+fD9YPt2PdvLbFY6+3WcYA/HN27huj
gcyu6XCLLAegDYYl1uJD2dbjiHeFb5BvUs9UknkWth63uF8fN/JnIW0h5/iW8uYi
3laU8rYYkxqAEDpxG5GiaDhG8LVLMiKqDhx4jUAECKCMXIn1E2gU/AXnWqlfjzWy
yNNcNp0y5irmycvu9t6oD4HnPaOqMTvplwwbQzEFRmiPsBdaChcVsvQ8WXMuurZ/
IXpeaEYBDREBhTS0aC5Foxzp0LSXVZM34zJM1v1ZpIpPIElbAgH3S5BmtyoLt3CG
QzjtN5RC9KH35/MNhLKqs5lsiH0xZ+4p+pu07Uit7X171juZPWUEHKbwQfe5Ps2Q
hMJMmYtWNcqU9AsoK7uX6aekxsP0InBOET4VbrJS4YhTf75utEEzsHyLFOSvnqgq
kCOAeMiQEVrWARmvKVKV0lHuFBkTvLoGRj4S7WulVAKWhXrGsNNp+6y2P2A64/iu
tm6yVo2QLrKlXSiLInT6Hlyu8TUOfMKFp/zaRZD0nzr37pZhJFje7b7u/5+pW/+F
nbPUrhc0l1gtEL7+1drJkJ53XgaRlq/saWAxTaA5YzFZ6XJFyqTF5tP4YEZNo3Zg
ZJqwy6A1ypNFwRPaVMHe/NGfIQnyj4zsypEFr/r1E/e9S1uiFMsGqcM3gXjKSKwG
PfNlyAPP8Gq139iUPaLLHEe7a6OhFOAf9rUwDeR7AEHtb7OSDNmzsdKRThJdIAoi
nXsu1rPOCQAbLyiMpljEEwtM82IvNuw+HfcjAcd6QD9iYJhsEe8VznSqt33i9bFz
u+NboZpFXF09vCv+lVLDR/pU7tNypBI2R5Z6h0VZjqehliGEtLI+pWSRQRRPYbJI
VIrhuphtx5+74PITVArxfcbDlHtM0MvznK3B3WL/xyoEc3Q/IgdJcfQre1qT/wFu
7NunbBZ9/GzYHpwDtGl64DnSR3uoxkUNDqmaW1XfbtYenl/E9BAHhzEOSb+2tM2d
RwCg9DwmjBiwhNeaHVxEvXdsSns7ZCsgy4vU6KZkQO5DKPRGuKk94Q3635L4zF2V
j+WspIGR7rVfCQ0YPDeBSKkigQTgLiJOH6fQ8mCo3TqpG35L1KUu+uPqHV8gks0a
Zfd/sIVVPIRchpEOnh/qzp2f8PO1VDBbx4CZzLVpZsn8M+bIeyUqArBPUchGdjrI
GRdyY8+5HtFx3pIiLDjAOVuxrxs7S8Ns6a1EC9R0ZOK/tSBNrqxreMpo7GvFzmt5
mS4jXIR5Tul/AwQ20kAm3e3tYHz1UEwR0DSdkuLBnBwrAlI1XfAEoAinGmUbZ/Ic
FO3YIDBA/b9Egr6c3umyIcpWoZdm6UM0I7qp/KkoBDa21oAxtwnKNg+2YBL6lnyZ
kd6yd1/2N7us7YGSEUAojDlDxwrpptEJeKSbGdN0zit3uaaeTh/HcrVgL6Rwqd6X
hmsP3Wf3bDNwLjS+nAXT+gJk/MVa6FU7agl/3ds1Bq75FIYB4s4Dvlv8QWuryluw
jorrZV10KwA/IUfykTn9PoIj1kIMbgSjAPI9t9aw8KSijsN3YS2giSjY/7lYqnD7
t3ed3WhI3Jm3Y+W9IyE8KOCkx5rEqad+75yRItoCVu++lxsrqMXxdkyRjrcTzrmL
NnGm/2tI7v4/XGuYRp/PmuLMDvePJqeZik1tguYMNtKNYvwNTqgiVInswkrXRIAc
MNIqEuFmI7BbD8arosPstueg/wSrOK81/hLzh5oRiGkp+HU3oElb6JrG2dkMuiCP
gy3F+YPaMbim4soLu+VQHPPLB6y2Vb8MvdhyK9UuySOwhMpt7tXiKGJ20363uHkD
wfwpt+CJWFu4YN0tkoNEOyUr7lAaKOMed/JvZ0nEYloOL8KNG5yy9sgq/rR/wp05
va+IY9EaYr3ts28SqBX6cWdr1FYia6/0yHiSktEkETdhOvTztj+f+/ikGQCaxTmT
Hox/hSlCzF0kH8g9Kn3KmNGAy6e732/3f6Kh1UVEvkKn9gM9nZSeIaKqZzsO8Vpj
GsrbGZpuAM39xk0lDYAgYvo1DN2HRbdv3cQLCq7l2ZGfFrmu8NJ1jBP8GemRrFWb
rtz2FMyDQAsGIiduh//kuJmvrBxlDQ4h/mQAVzAZJbsuAHapA5WMTUDjGnmhpzux
Nlw3qDOL95jkat7JfNPLBIEBFlE1QyXC8hfxNeJ+dSRCkkMkSYeXLAh7Pjcf2aky
O5GpnPOVEn9xCHTe7g1a2KG16eBUDi4WuIEHbl/YUNceGqPUW5Qn/Rxe/8OIDvER
uuSGs2p+WIlKbTsmjMHjtrIb2JABOVUYQIjopZY7j42xVG9RmqsmuSYm/GaIlSpb
KvaQ5PbRAuXy3Ucfp00/IS/UPbbbBWQvnrcbKSkF4tgOOEJCrXElzoYXwPu/wtHc
HEVb1HCLDb0JHYWImm6ztkwqd/ceXZE7424P8Z9nFa9C87jq74hZVNSIB9q+t3h2
MS7k59tKGxMxiPO2bvneSSuBoR92PndtEJE0b+2ROnj1/m4nM0AE6aAB95SSgt9H
5UKIz+nxYa1keOd6uRiIRwWPfrrZA84zedEXSFJQ7NajbFDDtuDGhsDg8Dk2J95b
fm3/qTXwYZjC9aqwhAfbCJiUUZm1Sr83JWDARN8/mTeNxtFvtoszPHFghaEOPrSN
5r7kH5NbylcUD5hLERFhZmKqzFYrUfq/6nnwVM7Ww0Oy7OofmTDIoSoC5WLoelUb
E695t2bh/15tSqhZGzri8NWUC+FpOjZ0/GrDYKidlpk+NYh9SZPbw6ywHYNE703P
LPvut8sYlie2AZ2adPXY2TR67xFIx6TeUwkh8THdzu3le1+Kb/4fcSkijOqaYA4S
h/wZGEePZp7nouGX2qQQwYOy9zLCuD0SvtYY4k1bCUXxMTVU1ef45sP5awfszZTI
8rtl/nJAyA3iwG888lO3zIIdp0Os82YlVXvWbLMXzunHc1nmeS5nyvrpZXiJceQr
4mJJAdKTfowYwkMOM7olYqz8EiE4YfeTIUOrWNxi83FoYRNRbsJxHsB13z6LRXU+
H8y9lX+OaTpbcBuThzHhb3K3aA9vCurfOZYiX3Dyf+dhiNex77+uNl237xlas37r
JpnXVx7ZFFRNhIA0qIlCuI7z4EH4PuahiooK6k1Ak8jYt3MvRve1JlJfqga3ugMo
riKQfAlMd9zxYgbBkTbgytkt2SRvyi64338P0TMqP1UIR6mdj+6BstDv/S+/cjv8
ghpxUIHFynazhvocMXsBM2HmExsMy1SrCbjs6g/FCEsupyFT7uPfBBi9eSVeTXAT
P733ixVdgPABUZofP+9Ssh/zVaCCjhDiC7q7TkVUtGEOtqtF/pb8EQeCAxr7Ghl5
X2kZ+r45t0M3Kfp+lfPBJJY+h24le0cL9TaAcCF27qfE3WqHEdHcKXc4G+fPPQwg
dBs4sz8JKGWSYjSuTChrfzR+HpUG+J3ezH8nt3wS4RLD+LPHJCL2s1seUigL01y3
5Npykdt2+ejgd0sDaLMy02Yx459fGZsW+d/Egk02Bld3Natarxs5xLLJv28xu2OT
ZV5vM9lwbOw4mNslm+YlrkqP+6Zeuy0N+VeX+20kLW1ASbF79WoZ05m27EwiND5t
3n/SGEyLFn76CgmsuXKvNYvV6T4fyle95RvCYQeBwvjxJSDPvOhS7/cLtxOclpqP
7rSEFZnEGcTMeD49s8greSKuhHQCRMrM2iJNc1nxoUr1bwFLORCaqip9I/SVH3Mk
XrWRFR68jL3eXA5JaeCXTGp3nWzFxpBIMuIJUiTxWURLM5VDPw+vEu33czzGHFkZ
UrxZ6PoeX78nartkCITkckQxNDJ5igLmETJsn3j6c/wkRHlewB387QwbovNyxVNz
b7sNdH5O3U2OxLOCOqssyHcDoKDg2p4GnL5mr9xAHDRt3eL0OrG2THXNQ8U8cU4o
qq6M8asmSIexB+gFIoBb6TRACmWmIp/WmAs9VqtIYEpkHCjnDo1RbVkBANom4jAd
2WKlWvLD2mmwXla7/sfKNLxbuQy1T87oECk6OcfaASNCDahxB1VmOJnctUmw2n9Y
CZFJ3rOupFNTmB6lPd5ukucIAX/JkUxlnmNk4Sezv5fbTkJjlH+0Y3V5RR8aIZiS
ylPePH/Moe2sZg4HBhm+DE3t0JXJhXXJfcPzO52wdVvtB57BCm4sw2ftoHCM+e1Q
jt6dpoo543Onwnw2oHg+NYnzVFd/b9UK71VUjPPiLZzW2SHVNpPscV4npDHINoPc
fXLQnhPT09yDhGHEZOWdgAg43grWRqNqLs2TBd2ZJ0dFNjEAXPVz0lpfEzYP6e+P
GBlBwz4VrO8Ait3+ntHeDPp9Is8NFHtfTkP1ICSnqJQM3qyvJHDZVGV+WT4/3UCo
0kJ7lln0lltU0ypgZRQlbbqmy6OQGdLE4Pz2FCaZkcpVMFAcqDvSCLyTWTXLOssS
NXpPu5NL55lkTKU4JftHNPPvESNWa3VEfx97/3NMWo82dJGLlxKbQKETsMCg4suD
KCeAdHkJoE5k43GXCxEcoNSlIKjbMJt6yLq5bJf8TBFg2vZHuHIfFUOW/tYv9mix
5SgWfyfuHQY1GyuZNe9gHFrNYP8bQhhFLrplsMVOWwZnZYII5qGvTnLn2ROx/5B4
M1L892m8Jo8jPl5+IK/AAjFTADryG8X66zv+kgLnx5lAM3V3S93wMIHrjByJ9uot
SqZMEmhQLznv9hp65c98RZUqtrAxewlrfQdJz/Ec14/rLs9VKaQANnGAHHsiqseA
VlVI9M64wyb9+aG9YF/xr1AFhJ7QO7S9CFTFQkAtnCZagZpHmI6/DkPyvvPL5Mhd
glm4iMv/zu2cPSSa37eqlvxjlqC/EWGlyggmLtOgYpiguf9BUrg3vFfjeU9f4yJv
RCDgTS3EnJkwlVosVUtukFekHq3FNqQKTymRYPeQhTahaQM86f2op+5D5J4X3ppZ
UckvRlFls9c0X4VPwzrEL+LfJGHP59kG1LLjjDk+jVhnMXPReXEDYACh9FaYuGZY
7P1dFXchMGw+HSYPO8Uk3sHawd3of/5530jidGqVx7XmnppKSx7nUxCKijrsuunj
0bOoY8khsKuzhBBsIKi3yvOSSBpMTFrglDYRkI0HskbM7gLLACqaKWNjr7f59gcB
mmd9kdOx3xrEUgYM6bXiNV+1u6/ljipQscOkNC2OI2xBZjxO+RpoSzPca4u3e+iV
dyen2vFAoj+IkkXR33UvGE0FbAjd7rUEGgj/7QENJ3bdTBOS+dL4Fhp2CfmpDkW3
cZKlD6PzDhomeVdtAHsODBsiIrM7R/gkZYUR/ykjKedbibVLRRTZa0O6L7jtoRgM
nIEnjZX4kHL06FRaK7GtHyP7hj0lf6jCcBLj5gnr9h5rEfo5S4Dp3rMT4Xs7h8Zw
YGZ7rhyXSygOSvZRG0jR9T74vOf21FBrVMKKvkFa9gz//cV1ApjPLhuB0wGGuWDY
MlxGCaY6uG9lipYZ5BhA2BNPCaGSag8GbiCvyqQGqfR+BGj+/qTFirwg+3OHarSF
m6V0w2xP2OuHWC5APrxdQ9qPTKoLHeGoh2ah+Th0aUzUwxNXRoBPzzuphfcB/I1M
iaZV6+C2QEG6LhKdcJCmeRZn1nOc2IpcZ1lIbokasqRq3CupmdX0TP/nAHJ/J76N
zG8Ota/e1jtF2AL8byRnr8HmdV2J/ituy3YvI0GPRLGS07/c5dnhILJoqzEcryE+
M1ZzP5Y0sF+IcTC6BJc7czoXS3c4/jhlHkw5Wa5N2qZ3jO/81fHmPeQDIXAWsAEC
OEOGyXHCX04eNEinYdYxcS8/l1VCYyUYN+AGo99X6uuCMAHjJN6H5t+63+XWK61K
68cOCdTKjXHACeEnb9JyU5eFi62eg0wg0jyGt81brawDnWbaa1WvWf2Cc5hiDKO2
YxIwGvnEO4fns2LAuRrPH3K14V3ghkb7uTQkwwNzKm912FuOYzKm8Jl86OFkD3qP
pTt/R/hLpg3NP4rff1w3t8CjUR3HNj/g9Y9hl24K0ZjMmOE//b/05G7j5pv4yUFb
/gpbKqC2ebJgkFzRgRjO4Wm8202MrnJYbBeDPw0VKVn5OK1VJY55GGyjuVPPCg4z
BjSjPXaJQS0YTA+CAiF2S1D6LV94Lv1BRs8tLZGdPJPN0qlEcDPKoUO6pkz6SUNZ
qfd73MoF09LG+Qo32RxwDUEpNeDWA6Lh3ji8RTArO3t+uz3h5we3/jbCQNdKisXu
z57O/3ilpvBrN+Vijq6al9pwMjw2oh6qE8e2yrNY4EwjzPy9gDiS34mRzCT9z+cR
H3uZ/BUgZj1VuR3RLS5405jZHpiAF7eddW2xcWdcXubIGJ9yJ9URhQkhImq+g6Rm
nsKq3RAxj2htjPp2M4LMGzeKKPNkEmw0mqcjbketNMIjrWzLBUOVGQCYHUtr8Nxf
1GFPPgO4E9TXQPNfaPth4RQxrrpANt7O6FhzWgsSWqvFtWpGJrg/9df06e7wkMfJ
z900WwsOX9KcYb+gjbkY+M1GxqozMhx/jtD2aED8oHlSr7q7hUD1lJKuARNb9WCc
KdyoNhUctN9qCXwLER/KvBiwQoCAdgZ6ZBLOUYKRJUTdewLXvWuSdu0NAS8+nX2J
MsSdSx6IiZu4sywJDjxaLvMVW8xJm10uQTlkEx6yXZx8tdt6ano05tLeIY/GcjO3
NCyX3G4dhckTKEvBTIX98UGnwbs2Zz0/0ca+ZpOSj9pSXz3PQFUEU8VyHm/4lKGB
kapR4yGo6QkgKSCPIa7zVKiPuiVkdw2359MI2fIFUPESbr5potMn1s3/qt60So2v
/HCeYJItSeBmwpGoealxLgedMZxE/aGCoTIMwXtFuFvpJHSJzTyItHsa1NPGy9Bl
Nw9Kft/EwtpTiq4ofTa/BAat1YGUlSkz/iQsALCFmJb6nnpEo/lqAqEITdT8sAuM
y0Rx2tm2rom+TKR0d7RF0M/yInBVxIv7rVfZ4FBqV9Rkn+cljqifuSnmPCaVdOzy
iHwo+0DW5netPzFopKcRIDj1QCAcPFSnDKUDWcbvX7LEwOny3dPBb9mhbRTR5eLn
p4yc8ttevj+t9vPRxGbPP5fklt9rfDQ+6vsv+c8AWnfPWC3GmPQAtOb0+cWbH6FN
sl1N2DyMidTkEc4uZyw37DkDSYraCXKOAtosC+ukGMt5Kte1c2G7+jsii/+Rap70
61s6DkvFqEz7NsUA6ojoP1u26K+k1tq37y2j81gOFrMX+S9hjFR4VQsQYE/l9eRL
bVj5Qu0tnYxFdsKov0zah6L1GbPZhJ8uAbH891TuqRLldtVjAEPvzz7ZDwcCL6mQ
koLvoxmPyM7gdvWeNO9T3mfvSthwbPupWqOvftjh/J+Hn0sWBv79Sbh4sIKq18By
FN+H/YO198vbc3L9GgGv/eLPsPh9t54NWTRSNDKfJHphpMbKCTwTzTHckImD99L8
RIv+UDb7gcpXV+aWjMOJ0RoGfMk73CZqOZSeTEjzVDQhE48Wqt9/q8jBm2+TjuNm
io3tfwPDpaDT4Xg3q3Yj2xG/U+2t+QdyRDVduKl+Hp5SDZyp2L4otpXdUaw4QbSg
OXC38UqJ7aEx7qcsPRJf0HBjfH7UZgXERG+8DTGtLLGudoJFqd1W5+6yQB2WyxB2
HLeavd5E4RfH4mwPW07c2Kf6Clc+JSXQjFL6/rTiulp5U0aWVyP+yXwqbDWmWhct
FtsiVfEDdE/eLretZK92CMovvrRQetlsSC1Q2ifpVLcU9/mH7Z4Zm5CnUUvl6qOh
qWRVugvUR95o4+BQidbokQt1z8Vs7QfG3dXJBXPKMwdcYaljciuqJExVPV8J15ou
F3FZ5nt1vjNYrQHbX9HB1C7wA89HnrQmXSu8LDayt+46EggDsuopqPaWUWERVRFu
425/Xfkb3HS3zlUpt+b2jTA0PG2YDP/5EQSBIGvpn5ScS9UVFwRi5tnbzkU13aJe
8N6MJD5g5aJqQ9s6SkMWHxxQrfvAcUoKFboeyUNtYgsdzp4j4qIGaCveK6e/ieKy
xMmZe1KECP6vEOjtFNnlutzNfPirq0WacNVRR3dalCaE2rtBqvmQDg0Pg0V5FWjb
EE/RnXmRrGzMtmsSCLXfiUyUb8aOSVNq+6tq5E+QMwG9//yJeN1Hokt1Rs3HIcEp
IFApwFXQCYA5DGw/GVZpJImc6bgt4yVLjHlQuPEfQOykl9g8lBwHv9xkpt5iR5C2
wlyzg2cAPSqctb+G7qe4uj0JYqwt5zUM8czM5oo7CfDolwxNctCv3bHgfZx8QZuE
cOODhb4jZrvoB1aa9SuqcijVd36sH3Gcg2HJ18R+zieA5VlauzK5+b85yCF7dWz8
IXqknf8rFnZxJE/EY8iTXJALtZvbcRBoZRp6h/L+8D8fJT2sk8goZV3gdMjes79e
cuK8egqVBabCD9BdMmDJZV788ZKk8Or+tafB/O7C9PzTs+2xV8lJKNCqu+o0hZs7
CTZ8JguWox4hVA0QWMU6Owz31tAC+bsdV2ERKH02Js6aPWBpJ229m24Fa3fkQChx
bJbqXs5JClslN84Fo0OsSrVU3ttmNj4ecdUazL4JO3LXYc1mRFUtnjD8pdaA3rNf
I/kuFbF/vlLzwrlDIUqE9YxKF9iiOVYncl7/unuIA2HjXZLL+GTK1rJmLxC5Bm6Y
XrDHF3uMgUYEqTIoL5LblHTftnxzmNeTFkvdNWN7ZZa7b/iellMk7moOgsDEtP4i
YyowlopIn9zwhiL5lF18y/IsAHMLJ1bcGzY7EbDal6esU4XWjzs4yO3pZg8TjaB1
zZm8uStZKao/VK8qF4wYUzLfFC+wgoHqp8IgXmif6lj1ne03qlHwiDrsFZ6LUOKb
OCVesKyIJHPufq1waVPOZrZl23kjQpXNuEs+FwSJBLlXgyoZMBl7axyIP7oRLHcT
2hsl/3pZgvSK0E/R+lNn8obMXGxUfJZqzrsvxDxlZFV/DFL1amM+0Ea72ljT81im
Egd8qCGCZKURH9dQuB+UJbrqtSV13QZoYxiSeTiixEOiZkKcSAFXOgNLRALUKsVC
nlZP7CRLpPx6yG//WUy8tPLAVZ9LEdf5h07hR7RdY7SRIPn5BcYtDJaTGyjdW4hK
ySofMuJ19R0KO37KakmiJ7wEKtV2jRaNjyzyQvMxRwn1IFz2h/oxD/OjzQm/Tj+/
Q9S4pvpAEAHxc4MPzMv1oLy74IUA5lWnP6cBhMaMbPnQVefnTktltx+lRIwqRnoZ
C+5NKxu1XxTtYKDjOkxpTRzzHCw0i6ADrhe8+SAXgm0udZi0S7hb1M5BClVB7NEN
WORVUKujlZA/4R6hrGXnj9rFhZMxCVA/3AmeFHGaavDs8UHvAbRKHTYAHc09ol1C
3k2MmLfHiO7rq/sF0NZpeyI43q2OO+v7iueRqE2b+xjPFzJ51u9lUrohhkKKa7Ff
ve1/56ZNdNH7+5sXrNDCMlWeTiwCOZjjeCG+6d4NEriL188zIl/PekfAbK8RkDly
5fsfa3rn0OZXWnKW+/PCvl5w3sbAz7ZFF9N0vNSbxr7GpT1WrwJjWxbwHh64DtFp
CrwjBLQGOUAX8JVq1z3KAUN+iOsIWPIE2kJq9yM3e9eu56oS2X2BL9Y2GptGr9kI
4HP+0iNvGAVk627efUhQAJMQSeCKE3rYvYJqqqfwia1h3kwqlARDkTatabep05hx
nNWTi6BoSgxBGRxEhjre1ChpHUS+2qj9E14ixXoavxiepANdfmBMPsd/BeiI1lCs
lfI7i/KXqfnfw6+0Lyn6CWX+JoS+JtkXYqGhxTid0vs6AbJe8A4w5t9/LaLs83N1
RHyzl6ihURcecP/jXWpscd4bfiLjCbALX1T8N5y1/O5+zhA8UZEyRgYxO9fBnWdr
7wwaCtJF5wDI/2ormYPdXgb3BwIPBenOHH3K7tsy7VL9qrMoDZeiF7jF2p50d0Ax
GKo6UUbz6l95eTfztNHk6f12vrzNIcI7/gBB2y6GSU2PyPgbs+81KYFMD/ljLSFl
3xUnVxJTZtiGVxMiq08sIERTeSEDSI/on4Ohb8nKiy3JKgtKMGiyDZ+rQyxdnBXb
juAxmP8+SyDD876AuQde+ospTRn/eavgFxuFvVSailovM/VBNSMLEEL9gEsgKFvc
qdObRCiXltknJS8zE9TRzVQPIhnyjXSFR1euaR+IX6e+RGL64CynniZtoyaLmzqA
4x9FO5PGxveFuW4aUjk/U1Af1aj4IcqOc+XkhcsEbcR7vGb6xWNhTRITfodSaGdm
UjMvWS2WQ8w0dYGn84GCyI9byTqkGFpy06bgnzFjkndSkSs+ChFHMbSTZITlcYvF
MepH2goy3IEve1BI+sQMt6x6qqDP/mY4rx1Zx5iEg4rPGvwWqjwIIESNjzFvt/pJ
gVog6A95s0qc7jR3cFHzzcSLbgWmul5kg3AqZ2XNlVGua+uEDB9f7L/+Gbk7HREp
nIR6bicwgjb3UnXKNGK9GAS3TqDFmFw6z9YR2Aws5uBdSmnNjVG4IKYfyyGHZS4a
HwlFSKWItYujU++upRFZ/BSgyBJQhJe97gxoJIsWfLEhPBR9JpR1476EUilDO+6Z
NeKqZoQEgIZstGpI26QmbeAGqVRr1m6xSu1kWVD6rV9koArUkqUk2801jBI6wT2a
pZu1kwFonMTgThp7U1cJb3vp9NI+lZ11ratc0b6sVP+4uv2Fb051Wo3QTuPkoAnc
B29pnQslsm+hSf3JtoafKizaus62AsmtblVdUcgXX5XgxgxIy4rJy4euzuVvsix3
h70gOh7ygGLwAJKBhN4IMT2NxG/FGL6klrG1LKro67Eah/HxQKKltCpFQzm7dmd/
GP0WTppzMrciVJXtl/nPuXu1Mx4NiEgIuxoA4zF4Y5JKEcPgTJsn158ZMQEdEZbs
yNfS7jec/tdhiheyzw69JIma1U7160f4nn5IjHIGsajeplA/0+CpXFIHjcG48cIk
wcRYsACtUNWhpJzJy8ZOyLJiJDJfIM1/U9fpVT3DrlX2GtpSpqBv2aTowlhzbMjS
ocpGUNkFFVE2ACry3Lc+6tATlA75LyCqmmIfF25pBExAVLnnAWA2I1IFinHenJeJ
sdhWmIjUTVY7Oi5BIDm+fchA3JL+HhfqbTSIOUmio0RVEHCij/swTMuXHFqeUQP7
d1L6Pkz8IHdZ4ZzGxGsTuA3NSHJkKuRWXtZ1nHIi4Z2r9pCnD9EYgrawOGqONWIy
Qkt1MmSOTN30sR+M4uBDt7VBORDp50grvghVX0+iawN7pr6NZiaWdAVHzyA3ubzu
tCA6YpuA3dlNhfOpfC2gJWfJ1+oD1RnG6y2TAfBFItGR4/HjBn+Fy1n/MKJ/rwEv
aPvnfeWrbj1zSKlhSMHWy16xiU0XlYfulDHaWfGLiYTlBE5prRgDpjmGBtA6sVTO
zZz2HYbXvfE5GzPoRSFh3E73Tv9zkk16Bmmsv4IVYyRQ9za2OZDyc16lmIB/MMxg
vheyt1g00Mh5ZCanoNAyuDOOSQKikVzN96j3g+cXoUJaC1h/l1wuTbwfF4v3aJXk
1AfsHIRVHDNYF/+6bakMPVbUiwiTS68CP5jWMi82YK4KhYvhgKNNArdRzPA8K8Ss
BYTl5QaeJ/X/Ps7dtyxuvBmYoYM7VphE/Gyw6cdouAWKgS8tMR6xQ2SiDDTh1kY6
DEvspKPSvwHdegXijFahZLr+LL0+MfPR2bdXt8tScsVCV+6Y0N3+T84/ur/3b2fa
xHdPmUKdVDfQwlWmXNRcmeWQEa35gXyBTzt8MaNxnwWA7eMjlJXsUccJSfwX5kCL
9Wmp48HLMqjX9WwQr8csROTQ+u0IpgTfK4Mmxpi7fUqn9/OU5Cq6zBO6SGrq7AsG
bU15gXUAc8Rf5HTn7eIDJiL2/vej144Qh78KPDgysnyVIOz13fEDFAtWVsNt7+Fw
wXlQlBMTKiY0sEYdg+Cf+2YGqFMiDVym5YHx1YmYlSpwOSSHVwk24LH8Ebd41gaR
C/Xa52+/YQelDbFrDANcd/q6lgc/OvncKT7sFFzZEbDmw1sx5jfZPYWHXtRnWIPN
WLFOJ+de/Cjhd9Y/VjxAmzN1yvXcOEE4UleEIYZotHyoXE2xC+x2HY0N020vjJA5
tqqLtHZ+UtQxBFOyCHh6UJPLNHHt88g98a9AoK1WV5EgQmM+AWkrzsYlVpIMB8Un
72VejvdcPVqxipud3Rnoiw3RNy5I3x1vuyACGlv/bT5WyC6O9eWim6ju49eDEwpw
H+FBTwBteL9nxJZ8dSlrFrugi8fm98DsTKFg1ZHPRjDR9gGta83N2ILjMs63a0ak
eHpvpZE9XxIcg7ffI9WJIQQfJZOzpwHuuFxOyLmfVz8DxggA9pdUq2F+Ee1Hn3Dq
JXF+Fh75cr10NuwtzHn12Yuv3YPPO0Pc+e+YXjJpEWwaDrzgbzJ24ZZa0yG/f0Mw
2vWRAbABaRkdM81f2Fw+aQhNf38o9lYBJPFgZtfeYLZ/YdVZebxXjONZz1id1T/M
m4TDDOVIFZpoJkHdSV8EdWdUl+VVd9jnZ+Xb44qd7sOJW4vHqleMkxB6C58ph0Fu
F3praXqF/vRHI5ms/UWIoRPeyzwuBuJk2/k08xxws3RlFNDpcczhiX4iwXvExul8
ZSnWI3xrSAOwbIbsqJ4QkAqE/Nc9Ik2XZ/ahMrU2jSEo/5RjDTPxVBCt1RwxCIt7
qfDUZtWt2PwRYcEgfpPDBC6XII/qk6CgJW6jTKX++q061INYXtG4liwUdXW3Lkt2
KoOXsjYr5V2WYmLdTNq3oSpIZvmtOAyOBxlFWaBDzk/f+EkqAhLFQmcxb/Xg4eJ3
3nyRpSVsyKq2MbN8NmzauefcvX8skW+XhYPOCj2sc84gep6URa3+PlalDbkcOQyo
iobr9FL/zv0Op8Fctz2IzcVFaMfq7tyo1EV5tDn5gmzFiD62LGPC9Jtf6tPE5B9f
M+QMiJ02QkPjiiIr9Pyrxs1nTzx93HU4zmeFg9EVwwr8k7cv93I0Dc+4NiNzf+kT
4ytAm6cYsXhDj6ZfTjaqIHk8p0x7vvhVXJbhUmccXsL6EgaHbcxuq4ij7VmFDQSr
S6eVS5p29ZB4vhP2lHqCmTDlPj010+QUWUSHYGA8pXbYNVtS5sR8LYFilVdakv4w
mglsVGBiuxZ1By1ul5pwA3VG7zSPHY6HbAKBlatTlZ9v0ZE7fREwlIEmrWrBN35q
RqyNUSU3M1ve7BvBwiV0OAQBGr0fNsEkGF5rDK2kOisYatbcGzWTDjUdHV+LhOBK
ju6efuWTQMkVXRz59Xbc1XbRgagiq2J4zW8MbMGGzLps8v2gvXYcjtRS3MWnDQ0B
2bjOo0CXe5OGTQGZHp/3WIUxiSUOSaZ502xhjBzP9Kh4SqWS4hP5SrZORd7ku4/O
+9fsJM0e1b598aAJ063NEC9AbzmcuMWqX4vs/5IyahnadOs3q9bjAizZbQWxYO86
0hD2Xtlpurt1mczjvhYkKQraYzaN5g8DDaM6+LQTdjsXEK6Nq0OXYgESS4BL5RD5
KA6fVI+7lanCVhlcHZomXYsc6UAWpoBGKwUMAuKVYm3YIYn/wTwSUkagkFqcikjs
H8rk9bg9Puh5/mNSlYbUFaYyCX7zq7uddU2uA2Q6ZO7RaMA4SfNAi89rCGNXDZIP
VEiR/XaNEeGcywCemNCu4Zzb7aWyTjIDyHxopmTPWFdHul5y7woaON+Ip0h7UDWT
B2OnE4gohCrYa4zG8YnRqeGhtPn0pWd4N3QGBLNhPgdurjKxKcmACW3f5KZclPN1
f7VQ5NzxCsY9jytvCe1OCCSNTSQXwbRQedNMtPSLYDPRRBz/uImr9WymIy+bP8nN
0KuDnlNGV6NBKnoJSEZnSoJfOHnbEXeHBSg8R7+P6YCNuoAFePv4p2or9ubHxBIg
OtY9Pphwz9UQPWZuZOV3fGCqZ1DVfdQE+HbRV6ShaiSSH3hQcBHQEEp/FIo/Fj69
XGtV/JMMhegx1qc81R5PDBQBFmy8oTl1+5+VEDKGVI8Wm7u8TQ7neSeSttijltxr
MP+gkqqtjze+BhrR7kiOA0fDyc2C6wbUgZJtyxYxzBZ+IdJ1vhVVuyx36R2Y6mzJ
w+9OuUQ+VMqDuQdmJt3DMt3aOEy9sIpEE2t8Fg83ZNEbYPKqhxuSlI2+Vv1R0J8D
b9yWCf/85oDd7e8CLq3UbPnDz5f9DZIlOoo8Up9Yz50VnLYsAlzVPqo/uKqrDjp0
qniBqWC2bXj6G/27lsXGT9sv7YJtlfApXxo1OWtyFnmkJX6/42HMrWAXDUSwThBw
UinotORTNWiPjP7iAj5ZjM/3ULDUHz11LIZ03JyuSdlTBULAcXfzUwXsYXtsFdjg
ckSsmPbYW+NotBZ2F5Ccaq3KJZda2wvrUm35sSJLT72HaR63Z1W6n1gV+maDRPBh
qi/QWbwov5ZLG6N0KpHegzjjoKCSHCnB4DH1NwUxJLhtL2b1DWKOOMAyfDx8tpbj
ms9VHN7ye/LySs0UV46y8oXrCl+VXuWNgUBIAP8KmbWKErCNZSn8BfuJShq0v9KV
rRh89V3hSdu6mitUmIVaBGKxuqnmSykdrGh5Ey/jGdqb6GKg8m4pR/omUYssPnQV
Ng705GN2eBE6o0WdkjcRHIdlIKHQr2Cfw4USVk241UL2eBBF1HZaQIMIScPxHvyo
WIOM3kmsnV9saFD3uerxdLA63RGgfNGqJAbQutOS+8p84TPyWKkBjj8mSRcKa5pA
ub+fmpfZgnAHhlreaO+v+FdPMYJBAcBxe9inY4GU4uvqM+kJkT2XkRay1YYB9Lx9
ae75JoHh0jGiO4w1GG8/NE/SS+12b6j/6+i3pyrpC5rPUu7aI5w+tVCkfEALOTeK
eg2PQK6ed5ypTJsFvbObY/+xrG+lrWtK/VcbA9ZOmPXu9TsT52SvPh7rGskNQTDj
+jSbjEArA57Lbmvb1Sipum9tJUyUdcxv+ltpAbGrDLPhRk7q0Ez1qeveJipo96+I
/ZCByZ4sKQr03azvooHHrTPVmC3a50/anqlfgWWO9Lr7cVLlGO1WsQxoWHbvMcOE
COK8Hor0aYyQBOuM5W8aEew9uOYGO25Q3GzGRvfk/A4Tzx+8B+47/x7IOXwVzUyr
CIlvGM9+e6m1nm9lgqFE3rJDtBkVQdbm7g6Q7hAY6HvZMSwT8nQLNQ6PST4tR9XK
eusGb8ce3xY6zAgB3YQU15ihgNub16sz+rUBaf5231TLLRmQwn8UTr6TKAthXGRK
9kWcYSdXZ6J41qsr9erHnfNP+xjT+YpeCHH64n9yN/wi7/WBzU8dBRnA9vKYDtIW
cRjAZmY2PzBM3mfdaEoPEfcgaoQYUiVW/LGcDzjgYTQhGkJ0bn4VteIUhcDdN4lS
RggxeBerfLXtzJ7I3s9noMXqD3Z5X5Grghv8m4KA4kNtNiy8zkubyILihFeGSi0G
hQ3XGuG9I8A1FGZL1zR/IpMiWcZwL8uh2G7PPCa7tX6CGt0SwnIE57Aui56Ve4pa
PO7MQ70t8BM2rBB2E7dXi05b5MNKF4CSKSv7d7E2nzVfIEKW74WStG5xC7Z1Zl7X
TOyrp5qHlXmExOPbdjgaRpAavqK7exoD8vIG8xJHmoNXWqfymtooRypQ3Lyf2xC1
7Yc8s9fiy3Hprqst1Vs0g+ynGK03/W/S8Mz1HNl7bXhiQMdY4z/Nku6PyAa7KxFd
QqgAOCBnHwuMf98Rs9tivMhTZFc4mqGjKiqbkFUUkjcyV4qKo7ENM6F5qyLKLVQc
XyBiSOTXSBz25sPfCTgDLZTV8rDiZ8aJ/Z9gwWzOYdj/KhOd7yMvTAAy7zF8BqeY
NFVuEYMzVZUqPIQH3k156A4f9+OSMBtZJ/nJceoGbbUIhywN3f0DtTqDaBHHdOe8
aqRXiiDhbDx/ym3YlYs77QiooUGH9vd3mi/ub0LlisaFOLmO58KTAHE/gp86xgyQ
m0cju4XPu92rP9ztit3C0/xc5WJjerTETPDdB4Dxwj6L2ezqP50+E7ZEgkBMJrd/
V08ZVBaZZMm/7FC9CV+jEnL3MKn42sPzFzyXqzVZyWDdoEpeYvZ5H5FpYmteE6xm
HsiSumOK1mT20Ah0oihC6AHCZFTa/JHDxsOTYV5lMmNL0QW2t6lB5+5vwesxGN2T
n3kERdsD3b/AGX5nnYaT3S3j5NWJgwUCn6FYqFFZwNwVCNYzEGTlUkMNLEgOtfrx
Ngi6te8eEi2Bp0SY/Wxcj74WiriHl5p+QIDxT4epySzgiS4L9FZLdyjhG3NlX8OI
HfJ9anGSJ/m6stJifpJnIspXG3sDDQ28nm1KbROnJO2MApm6MGOFq2ZcJ2NURgAb
qnTrzMQkoHqKItxg0WjgOE15rFFrGUrgAziBs9PjOg5eYomipRY5npK4ZAcW/pkq
Nus7BrueQJvfsvxjoBvK8hHik8qXr8JZg6JvJXJR5YFm8jK8QMnXHf+EG/perfxs
da4qe/9Xql7UM2nSkYAXQyokPrTPPgtMF8CncXwNn8blTF2Zzb0+F1dRxRlsFCVZ
5K1ZUA3TeDTXmaHgYRzbPD9bPhvmlnK57R4QmVBTX2QIrPDYeh3SlVTebNMaodu3
yDCq6ooJins53NtjttR5wkIt5xKB9mSeSfuDeGEcgkxb9n/Til97wWeN1UlilrGn
WDK8iAO9BBCIHhctQK88fp/Kg6VZwOZlAgNyT4dSRD54AgaZNlmc47IQT7LQnIIC
Vr7KDFs7Y7lqg83WG7LaVBnC6wiukvlm0cwXZmuvrKEPCj5iMv4O7ts0pyQEmLO6
VDZN5ar/miQdr4gCMbO8z28ZQYo+vZr99Qg/DoXSpE3z2VRR7HJh8oeIIlRcjnUP
bY9Ky0UzHNjhKzPCFUSLQPXoWYlnoweyLYMTcVHh5M/NZiPVO1KqLt1v8VxFQJoK
wFHuGGcHxaveO468ajzvOF7Tu5WNX32iCNqClC6tApsHjbAd5yU0K2EX8yWmDcIu
WT3S8/HINwkYOA5azgD0QdJ1YabzwSBozgfI7RtJrJVgtoX8RAqUGzkDeUBgPNrA
y4WDBfvhEz/GsLG6tcNgs/9XMzbtYcSds85wAX4DCrdnjFh8u8gIMuzeHtblF1wV
G5CtjjeuruxsTiyhiK8HOwmw5IZJyzOz3RSoJnTRh34GN5YuYHx0DLkAwc2D/59X
fX2uv1nCJoJUOWA/RE3xwPcj6J3086TKMOvnnv2YZh2sn29RpkHD3pUhpMALF27n
U2OsPUfHi5XWjDvQ7le8wcRTBPx84SS/bT6TAJCeAhUm/iRrt3uEOmJkI7bfgdvm
pB2ccHx1U3cJxUsP4saMoXVKO/9JvmgggF2YbvKqJP/SDC/8PR8uWZ1LU1kE4Qsh
C1AUGMROqklzqTB5YEAjHgf4SzsH1CWf53I1v/fOOCVqbmMF0O26UxRMswuVK8ZI
IZ7lofXC6MiEACYAd5LYj7MWzADgNxmw2dQmlWq39Iae0Ay6rYpE1tb4DFKsBH1T
SjJSPFq5MnxX90CmaWDCH0cMHgxPuGC9CwEofb1N0gGIT97Rh7yDHGl+sn+HH+E+
W9tBxkg9S2VXV2e6dXl6s3bK2GZqOrjhqccf/bD66Nqn6c/iYTAqgpoynfayLM88
D+8F6KJd0Hna7V06Q+2Hll9eFjlF6dOyw91R3ZNxJD547B7e1X5vEDWzOzgHCdM+
fgnnKdYv70wWZjMDGcEwNmqYjH5quFGrXAi9StmDxAVUlnENIz6Kuqi1pvWVUVe4
tu6ZH75YQ6g7sIYtFdkLx6AokSX7aHezo7wK8Jzs4CqEloC+zTm1T2y42MLYD4Eb
efiATXDhMnk2uj2WC2fkZ6bTZgxIBiH/WDVMgRVQlaay8jG/p4j2srbed/MP1Js3
zVm9q5qZQ1h3wr8493dLTZUprRucefP4RMlCbz2dsRZmf4MgGi5x6Xtxh81EDUNg
jHSZOgE/OcEMdocvi5bn08he2tH197m9mnbCf56ZKxOIO4gUYfart+61uiF88/3H
1NX71wpkUqyoE5YQn/cZ5eJRiZOn1ui5+eZBS7YugnHI3cVre5XWey84fYe5dIUu
NbVUtC18EXrnfchN2/0fCMwOPd/FdEDk+ssBacgraeSnalr/FVN6Ellpf8rLcUXr
mdfIUUgEyjL4U5kvX4yXcO5FOcHSZI+bG0YhTHXE8X7+9oktb4i5kIRcfILsF1Dj
x6V06Y3/tYSWiLqeUfNA0YZLG3GYSd9YCupfPCXx+b430xvL2XsBVCyPU8Wk6Vef
2RRlpTj5rVQ1yYRZlnFrIlFqGtLaPqA74WRzCUjUIUjZS14WCVkvY5p4yyEmHAcu
+/eSHK5HdhOxZmwFGUdSrEH1wbAljHWrPKwCkSeZWrkooBDwPm5bfZfHSKCDVGql
3UWF3PcrRE3WbPkvcfi6kOUUwDHLTbNk448UI6r7E5I9m5WwlHuOaluDG42pCtJj
oUhp77llEabSe2BEAacqNwbhaglaGsfYdAYpmX3VGghxvUMAb/mNztXgic69drFc
W9PlXztCMDudoJ9XTcamrvV+XKepcjFYqtGlzCivLLRq3NKC8PBBmzaXz5mQdM9o
QpsR8AIdrtFVUOFyn13Y+efWrzDUsRtNWMOWdLo1q4h3Z2f+KITqUnMfj3QJq51I
AGibw8u7tF+3BMYVpmU1iZjYJHxlI9AHIQrSiSZ8HuFuGhqnh/hGBL0lw0DA5ItF
juX8BIQ7sOjAuxrILZunFY3XYDfo5KSESyoGu/AskjPXg74ckl5HEDaHu+d7Y6Kw
mkyucO/UdazpZpjEFQWpnWyT9IyA+Sw2ZqzDrki/H7TM+a07cjPxZKnJPJXLjlQZ
kWYM4ja+PuXJeyn/YWmUAnY+oDrXVyKzvTB4xymfkbu+W1oNZgqbHCgKMJ7q8iiN
FQ4ucsuAkOTe+hqmmmSFHQ85no5SeDHte6PL/1E/5kWqNvYzbPKeVy6rC4L8AvoJ
oVlFbI4luCavyMg/rNRQvE60NVPHVvDOaRVkpN6at5xm0lqgzRtXi1Dtxouh47nj
hHOdwbBiF07UkPQoJvxTLinuGlzakkzEogcHqiixSSW/OKvT3/KK3EJ13NduxzT/
k0W9WE6WyBVJtLjY3rmCAoARBlzNLDxSCOePnEWrZrUSE7JIqPdYQ4/mp8thxF/H
615A3u6sSQXzW6JUZs4PTOwBt56j1t6CsENV1w3U5QyrMP2kxyNtAJU+UKBnq67R
belTM8dArEbo+sMHBeMfQO5viKTAJ4Wkbx357DkxBs3AbbqkPgjT4mhj7yxZrsng
4tpyruuAd4U4nbXj2F05sKZz5mD/QbFlgx54LEcfh4kt751xND+sQ8QtF1SZuq4Q
3y+sF3E2IBq4nw4sUlGbbzo0qYSmCpLKAcNlHd1jmvTKvv9nseIdOq+kbOccrNd5
iYBrr21SxqTQT/vHuBxUjHcpgZMlLy+Rb0EecD0/ztcnDNX9UDNQyL5FoTjsxMjm
lT98EBrIeE0Ij++yidy1nPzgLBSLB6RTzTkE74B/jr1l/ryNnSFKqh2rGPlI33qf
6yLNSR5lzPBFgzTcT7EaE71SYi8EqOjuhQ+KGuziRW62dgmdBsLofhaue95z3KuI
Cx+q3uX8VdEg5lYf6r5djNccdN+0pHwoGmM7e4A89Hnhh1xAbicKC9CkLln4RZCx
N8+OpNc8kCq/6878HFf4hUam0XbuGQZwk1q7hJTnjkuEXlGYT5GH5IWVXk/MQxou
i6pW+C7554aPixRSNvab/CoRtW7UBS0HBoR3468vd4LcMT+TCNKCPt2QIhM/So7g
XogldVg0g/1T9Dty7bemawqLuWjvOIKiNGkA1DuVSHR5BcbKnh4GuCK1Z1yp3n1E
A6INPGkzuMW/qUULcl7C5JV5M0LgThXUdMg2u8ZqUWArTwnSGAiEbKTtYV082klT
vTK9OHTWu4bqRC/oL5S7QeE/BYOt3qiCqzhqS+5t5nnECPX+tOF4cNw6mWe9MbRC
p4maSytiWjK3DYT6yhM0VbTivtkn8d9MwyNdHVpP2JwOWYaEAlu4An5qQRbuDFHW
f8hYEMLY/XiPNIypNLAOc64mQegxIa7c+yFqB0HD0e+sG/N4A4vokuONcLWynYlp
/okOBjWWW4XK2ztseAFrK6Hp7YtT/ioqB1LbFI/UgsSAxgB6szVyZ2Sj30z5ksB3
836v5jg21Jgz5bL0cRvdcWqwIbsiyM0SsjIcsziqIoabw4X5zZla59VE1XEG/vXX
rZU45KFojFNaHAkUXXyVMNY1J9VOyESZ7snaLBc3K33/Q1kUKB6/J73OQhYyzwy8
+jzrvYP2Ba78kFZQ7LdKLmyTj9CFuERrjFiJnI+OROnxVxS55pFOMCd3nY1TdXy9
XZ4k2dcpVMhNVplMkoNdHPuVkqsbPqRKwNWacHBIasOUk6d2AzGj0U5ufALOqkW4
qUBNknvDCGfKM3v6mqAMKpHnixvTd4n1i01t/uYGKehFoD2kTaO/gJqDmk+pGQ1O
BxmIb1tnUbhlOMYrLUhLmXlH9B/60qQeVfWWZTxkIgVtLMnsFk+B3AH4hP5UxyQK
GmjRrcJ7F9/8D7Zr6YKJUwwiyFqJ1zRK3BXJd3HMhimMuvglhbOsO1KICOetut+M
9Iu05lIuFARx3MPedmDJuLs05vNKnW2bRUuunjkk6I+iFp4c55xzKSWt3U/PpLnL
bcBe00XH9m8tYSsrt2N5RPRfVWYeuZiYqQ/+CnVma+MFq+PzcROntZfb0mIyZIrH
QMy+PgCwGY95jKq1Mn4Cc6bZpca8+gCvZuo8ODAGti8Y6TMHjRN7lKGvRuTKEX5V
ffwiMYcxTrIPWxtP5q3gWY0tJd/DLQy6ZWz+MnhgfQnM/M+IPFqdJrwPEF9fHF+0
yet7GlHm/WtctBi78YTOICh0N1DrtiROitOPeO+9QV4lumIO8XHF76qJrIHx8VXg
vIK1nAitdFSvZieMNyL86xZFlBWtgeMvNE9Vrdfh0vZLzc+yrZQzAkwAX+cPjZ5m
yCTCtm3FAKUUA4S/RRT0ac4og6CqCNUo7j+8rgVPLsjlbDUwrwEXa+XRyTF1yX1s
gyOdd8sr0EvMtvi+Y55YL6MvRkOTZZ5N9yv6XxNdNNO9zd9oyDj88rFjgjdvomz4
lYIw7pWoEerp9J+D8D6VBNg7sK67DI3i9ukGzLmXJtNtbuFVrlOOStxyEN2G+u/8
xzQscsej7W/r6zt/IvSjYaVRK4nDN909eCrv4R/elcMssE7UmD94icsnFGH+cWN4
VFk+IHq6+/BKto2o1s9NVoYuXeYBD74urbyC2bjAEZ0pp2roE6Cv9hhHjdIFl0wy
L4H98lNzrMlBBdIlM+MMemhq2XJBxG47zZ7nUzAK2Oldjelnwo9vtu8md2Wp8HHb
0ECs8Wg2mQit8VKYDOHOLz8licXVHvWgi64afTq/dIzy3pnlZzfH+Zldv/p08cc1
50IIbdp/uTYL0CaTPcxlKdMfkuOvPdmc6CG5cQ1QgZFVk0TUo/XszMLuKQRoZu0m
tKuUTaqVQW19oHErItFCgPyPDtaRjk6G9Bpuh/cgVAGHjX2t117N5cJpJv7mj3tP
dT46xIwOFh6RvcQeXdguW80n/V556o6Q9u8Oy8zuKKsbv55zAIRXQHbuBHiyM87X
LlhOsdbMRxwKBVl9rAZwwe8wnC/Lo+8+GDVgngOxkZIjyyaSL61K0edY1J4mIc0K
sCMI4xQMwffmB8YhtCckPgVHqEpC9turNYrsQ5m4PWNmjJ33kPrL4uCemIxLncX/
EVXmWuY7B2wl30FuKNjBVNofla1baVXVJONiJwCmSLaFPMoeLbXvlgJlpKRU5wuh
iOUWi1dh0hhCHPnCI+VIelzLsfT5fbqAtCMwmOxWJk0T94LWvQw1F28oL/qMK5m+
BkQ0ilO0Q+RNLpOffo21i1EBltmFO/bmQ0LP3jRc+H8OJTJgxFowzq/7s+1vhqVC
EQJZQn0SHPJAgZvBxk6p6UX6wfD2HeE17YGzXRjeLxZwUGx/uo754hjf3WE6/fl0
YW8J2qPZplZoY6cwMmv1qUPj66qFvL5MREbcmYW6h11xX/cEnncJggx1RLVMInO9
QZ6FDmgVjeE7cHHG1jtCNKQsJcwnyd0rWtEBQ3m3OLrF7F+ITwh6kdNIDul+Vcfm
gEtj5I7fQKmJnUYV4S1TvW495hPTatPMp5VSqlxl6pg6K9Apso2oedxDChol/8GR
XC+P8EWsP6DptGvB1SsrYqZYfY+iccwrr/P1uK4lFHeyxK9hYzeHoJrY99kNBfMu
BLlO5DUh0dJwsy2fqpYw2WqXiBPhqpf0//vy6tB2hr1b+i7TJBiUZXgr12knXIbz
MkZfzlMW6/zEY0CQhdftKq9/ds4ZczNld2F4RV0CpWFVLteAu7sENs+rC26ZcDfi
WBWlDXnWb7OTaS4huZzJCrZEH3GOX9AAL8kPY9Vd+qyxNLGICAlUPnY75s4hLa2C
sfmqmL+Aa77AKtLtK9i3DUbvXqWgDyTXvD4ulidJZArfwQwbf1hf8cr47vW6sOev
nSl1xm23+gJA5V68XIXi1TkwK1B0fO1cu+JnRup4fFEdJR7VAQT8jA3Y5n9B7r6w
G+VJbDpin9rrQCwl2h6aLWQy63LDAWK0ylKA7gviIhK+KLTh2aoRJrvu6xcAoZok
qGCoJy12meuh2jIh84rx14oFZJnWguO3gnlhJD90QHWo6zScsy1qeEe32nuoSMJB
eyDIBbllXR08jVLciIYMY2E3ZNv5+vEb7TNHRcTc5FQWq5PCz3u3dgFsYgWzMEA9
rH2tlOBLdVEY61KdDm6WC/a4Q9ugpeDUbPYeIB9AeNf1spnPhc7IuLR9aUt0Mx2n
oXngMZxa0n0sXuyQO+6quGoGu2RzxjZKybSADofiR1mDXz/PCrJ4JRZSojBip1yP
bosK0s4VWwGSEDqY+r646mZhDnQRo7kzz6JjkuNxnn6R4zUvFie/k4wWqWxeXOX1
UEahLrYB4u47ivTyzNayWLR9Z5n6Ws6zYhrGZK14Gegoa1EvNBLVaakBNZa6fKdX
EiE8dDFBb4YHKnVm0nyYJzQRKTDosWAONJFOdVP3+zUn8nBuzVgsSfQOCaTnfek0
G5mwYCyWid3x/T+CY591axFNrg5mWUCwlhM7PDx1HCgwm1i1Rjg3aDDpmlaI0YdG
7jjFxOJtP+kD1OPIXOYND0LsfckYiu9QRcgCxgrFPbVBszbhqUBOOtrsQXnr50UP
2QEqKn0GzAR3GxoTvpRUaNnz0s8g5lEOElJT2bM/ProK+v8GjyJxHQZWsFjnOZeg
SWLBBsGppHIMN0ixaUxSJG92n7xnCIO2TZUhN6AfP7Vqo3m5y3Ib124hKcmgGFQu
EQkW5K7M6MFnr6dwgYqc+pciRR/Z3hMQaLU/8HNQD+E66im2/k0gpWitz4sBom3Q
DD5DxbkN5lWjySYY3QFqJ9ZffntwnKPuG3LhHFW+OdoI/X4FZ2+3+tPfv9rj3s3+
+0wWhVE2VWxtJnFT/WBghnq9YaAqnZ+iiri8ajlpZtJjDU6rLFahUAq/thRcd3OR
Al/cGRbrNrxxiGf3Zx/h+yznqqlQ4ow05232uEN8Hq/ixzDu2N3JIuSr4rdF0HGe
t8KlDdOTV7ASTu2DQvj6U/y+xdOT2ECJgWAGLWkx4p74+ZwKoohWdtTl0a+tIEmY
LFvhSofekSWSB3GlF4iGPpi1cuOwIZm13jU9Cuad2UaTfsUGhD9Z1oaY5h8NJm40
lT879olKvQibadmfHHirqWDFGJI4JsgdfIjrsXbTUpXUIV7MMDaKsDVoRjY6iN8p
+dT/q9kD5bN3MxEIRsbVK1J7+/bI2okSM6BzvWLuBivfqSN9ZpDbuFD9fVf2goKU
7842hIvP3O7SAhG1YG+4vFD7DsrcHsf3eWMDOIjZFSfjxkeSvy19nJgA1C0sDEOi
7bFWbBjFCcddO5WfIKfs24lc4JUXutDl+cJEz/QrIZp8LV0fz873P+MnxA+LtLBl
eXGoiIyZNmXYuVeEt9xolDX8YUXuRYuNP9J5E5vuSsEU2/3j3+xD+7nbI0ob/UEg
z0kpFtNnDNT1L9vY5BFpnQSQVBi6yoMkoXWrWxr/bycylFNEBKuZDiRok2ti3smI
ezCA62JBTOf5b8sg/CJcwobnsAR+R2sB0P+Zrf5qLrC+u5v9EsDMHepylxIOxGwh
yGKfFD44joqLLaujH/z/LpaogdRVGqhjdnGnyg3zcUZCqtSm5h9kl10767Yex+am
0q56+oImLmKQL0Xm8j8ZFR0UV605qSuZA0JyMMh4tDbFv1vHA3rqp163maF2jHHE
6h6SFAjOiXYC9PVtKwTRhPIHr07ExuGRRyE+LxAXl9Ad0ewz8gxfVPWh/WzMgMan
ymWJViCZPGwuEue7pYJakmqWwAFPnJnZfA1ZdRANxVrgbuYIHlw6vko7GgsbFraU
ooriMO3CUuNz8YpaapP/qMk2Z+4dS9/1H7kCjCi5XV7u5oamDyx5jULMtFA1i2xE
F5c9a54salzFMv34wonBmEgu1Z40Y11AkQ4Gg39qXlsF7OQSoWL338vzyyjaRVJ2
hsmPD0Rp+ZzIPp/GvVqq2miMabu42FbzJPyQjONQ6FLc0IEY+/rX6+REGG56GGNi
PPgoAT+mL1keppLDmK5uadXT2c+Wa4X48K5HfgfosoyOJ+oteEfozQGbOGj66LXf
MozH0sUfehdHbOvA8XmZR6vsHm1PN3u3F6Uv4CTCs9WdulsTg5MLDDAefKExRMBT
bnTeCQbSvvotnY3s38ONN2xnigugavge/afjws0Fx0J6kiGvd9NUTHnOQRsrn2so
c5kxs+NjWtlVfiUNL++fQGpzkWP9Gs+NbEiA72eQshZkkupLt7PNSxcvE5EOMkrA
jafPrvngYb/bACoErm/6gknWE1w7btdRu0GVTFy0+RT1gNj7UOdvWmrJPr6VJm/h
6xzoBvMbgPnvWNhelIeB7maAgdlrckFQnCKo8RlzkwTSkxkez7coMdQlWDcaZTfC
LSWgaY1T0q0HMpCco8lInBcG6KVSyjuDYC//WahYB315Wzzf0a5FskWhXRv0N/Z+
5SIKOmYEy6bltyBsXIFkYmOOcI2CcHbNtvawUD/SyVvTwnGSU+4/bzY/qXgIokY+
j3pRSMhN9RrJYGstp7PO+7ifJt+fd1naIgn9vnu6hZCRT/svDgdDArMVYO9aqqnL
rckX3SzDRg42eM0pEDoLE0Tkg5VSWlh1koBipjhADgjfxF4ZMQI78BGA747//APT
jI30RZqhTDHnWv0c32MGqT/q2FqrrhJYxiIRMofLJH6nQbroMLiAUd9iAMlhRAs5
D3Z29oZ6/CMGQ1pMvOLPNNe4q0fgLNdYd3M/PEDGLCiq1rkeZxAvRg4o3pPv6++a
iZ6Btfpp8z/UD+HAQlgro/+VolFaE5CHEY4sgAl4SzGq7GFf+BpNr4WC1kazft9A
oj3N/fL/Y7UR5sfCGYQWYLWSrumJtkMiTTdJNaq8UTJDRBqrG/Jx0oQY5f7GFE/f
hl2i/l187BN57wUZMuj0RT59bFaGfEH4peV/ENRrchQpICV585glhqEqulyY2fYy
e6GMvDUMsyYdMl4XG3ra8eNnbtxa3rAA4XA3EQDEiRpWA5Vzn60Z4E0pj/3qXmX7
lKeCyGlklGCvLtHeCcrYCzbGJ1BLv04FQN/sUEmZaQu5Rwi6/OFDfvdH0VwWEe/7
38SQVYVNsyDstauhUDTEirt7oI1r/IKNabeazFRMurzcp/ioZsUm67SqOn0XdBJL
kA3bwaMQLDZ9V9ubn1vBco9FgDpKaWL4g4fLR7FrC13EkOHpJIsuXIMPw3jyQxYp
7DAptQ3SOD9+XDf5m1WmNovvIGPlKSzeuzJTZ8yJup/gSPooJj10501iFWrIsMeb
+atBDO+4YgRczu2ftNOZLs91/gn9pS8ewrw0zyHVVQLMV1JkKM+tTF8xSIa13Ikr
RB5o1u1+Acd8dUmnfHSFL5gqfp6aAzWWBszu1RgEbrUqMEntci1idoOOXMPzyiAL
FiPkT9q+psiQne5itKkcON7Fh79HSReLa27uvLTm2zi0vBsDMFqe9BVbc7PvAfMN
KVD+KUGhodu2HczEFBerr4Jf5xAvght/0QawA0/3Rn0Z+m/eQxrYYr9vRP8q9xOq
DnBGuNHSRTKI3o4Bq8rZnral+O6VIf4s6OZoIqOnVlS2/dySBHKDdAgREyDKm0dq
7LaUbwOyvghf1Xkvdo7CuI3cODx7gySPotiBBzu0QpBOAR3lkkG1bJjscxVe2YpY
J6mVX8qYrm+o+uF6KiEQGWyjQYwLUoWyIu1/uWvWIZPa4vpu2Kr6iCI+lVTPV6N/
or/0KgWSDqqShfrwHtyOsF+/ruzXC8TLwn1PMpCstjVEXCqtNQ0GoL+HBnZ7D7IX
clVDqjgWK89GoiHikVENtFY6RLwvuBD337nHjZ1wUMfahmXClo7OpXr7/44J5dBz
1q7UX8RWpL47D5cai8m987Yv3RcYIbmxy1CVXs51x/A1oL5THlINg58cmojYVGLh
dKqaptLvlRYaAJxWM+ORKAikP6K98wnuORd4fQX1LYo+igJmCBHT7qQ58MxTyB5b
TbJ9WJZQhyHAxVIMEoC6Tqk5TrXDPSOFb2C77Ysi0EChQgplEeJ6CWpdgdsVShAY
Hik3LSftxXTDGKTtTtkR7eKoahlBdgnQw8L2Hxd1A/8WtamnFXsrOND7WZZ+2lMf
rc6ptjQ6WHRtAgIR3lad27UoaP69uzhZU1FPzIfBPJCN7h+0Q3kgDek76E2fb63G
BKenZXEeU4CV97CYF+N8lD6slP+zaPABxpfRv9CUxNyu2MdAEhqLvfXzfMoQgCVm
cX4ebYLj4vXB+49LEI/wkYkiZY+IO4AA2QrcN6s5Kmii0XaRDS7e621DyvT2GZsI
Y7gjknunnqzbOnDM5glyuw6Bq9GtyrLHpi7sl49F8omRBVfh366cyNNrw/21kEb5
In3TCdBxIWRujZL274CztW2tVSt5Pe0EBzFs47acEFarddXK3cLQS67TfNW9yaVU
FO/sgAmKszksIB9A/zF1KuW1rLHVvmN7qjYRXr65OhITAdT0NLfGbOWZvEuYPWcU
hF5F4Yck3LBL4Lwnmwr3bO9LouXVXx/o1Myla4krHPM4N026Hto+eXyats3Qqclf
iVDm2soUlLaiOQhxQGUjz8JsqlT87s8NStLeyXShexJ04g0EkYZpSJNFHIfUB5YN
o5K9kPLo6utj3ev0ApPs49VGacDIQ9pna7iy+dQsylgjK9QAwWku53gKwE4N7HaC
M1F3FhPlGmCUMEZBtjqX2+Jpe4SDVJAI2ELKixMCJd3ZkWuii9xuVw4wHt5hEl4/
nR5TC5RHNKmXkDt3+ny63x1hufP8vbkITxZLXDJmJgtM/NCUv3CYSXnpStX6Y9/I
AqB69HVG9dRSKsMQVnQwa6UBBCFzLUf7M73KtwOTaRC+FPofILd/RvJDnp4/uX1B
CKHWhBnBZ4xoALJ9AkMv0qQ4wJu1GTjRhLuvZlmeOj4xO+eoQB3kETAHSx5CHYRw
R9AqTkSjJV8sTEaHwyywMNSzoUi1OdEnFRbnoicLnqN70JjXYYiVVb1NCsKV6YUS
4j//1A0s3LqJoJhTTkf0Z6fvvNeMuhncSsUTHQNcscLJkVgKdpT00HEgXy3LAf/f
cKRqUegCB7i6/VojwJhNijHsZB5JsImQ8IWSakiIpSVCk6/+6s9f1Ep5O4+L7IXC
h7hX85S1GuIKBqZsvrv2QVo7Cu66QIspnx8TWckagc67FIeM6QQ6YdBG2Ns9iI8c
HII6zM6V4pClEpgGabnpCi6RU0IJYzU5fDhjl2fQbuPCAL2LRSBeb+hFaoiJo2LE
W82WqL/kgY6WTGj634kcUZ2fdKvZ0lvdpaObbkej2akERv9WXJfWMw/49ZF5CF22
We954YCGy4N7LfZ4tYfcCN6TinbK4goJ8pxSmfbaNlnpXA6lab8pTA+DHiDZHnz3
Cgyhzx8bOoryZCgyJ+feWfAquU6ygYSchIIFr7CTkLSVkOcvCJY8Akw9BUQz+elO
lmnWurCSOiZdtGvuykHUHA4kGRKwtzYhwxQtvxuGXyCVSNCY0jsz4CoAIFa6wHNG
TdBzOmUxxo2eYtZ/QHd7XdMX59MWWJFb3eFh0m3OmGd+M84s9STmUpYbutt7IJJl
FO9OBBU8xq2YZOg0esdiwBW7Ha1pNQbxsqG3nY49vUp4AExfWDHXLfVl0d9DQXfR
rNC5vqTPfpvrqv3M6t6ftczZjSeMLaAowcG3d4CJyPUIiBg4DM4Xx/sjVEYR/c7Y
tE5EEVyg5DnBVeFHGUDsk3B1ikIro9j9ni3uTzzRoeeSJWbcGyF9GMZp0et7Knj/
RQn/ZXsEFYfDnT0FBRxD7SSiG7Rf/ftbNJBSkwQhwD70SSazKmAHYiBwYxqWrBks
XzFnjhT5w9n18ObRWXGCUeh10Hawsa/Wsy02xefKDY5YdH8HTPxmAdafv77vPKkW
Z/5amX+vNzgMfzVSLFj/nilyj2gjCcbK+57q7IYpS0qN4DdDgzUiGHpjgi7NN24B
Bo8nxBjmlMDSA4+9zT9wViPRgOVgwV+RWM3+9ExH3jXlR6d2JDsAng3fiSjOyxOy
wWyo8Q1IKoAHOQ5ac9mKRNwFhybLF1Ffgk3z2Wjzo0KeteSs89aK1m+WjkMmwkxF
ZjTmNBgmMfi4ItntlixEbl+C8+Dq+eiqL8nzG2pBb7svuCPcEta6cgjog6LGZM56
nXGRNZf4heFd94x/rQUfwpTXUmJx2Lt/oSvqTFXPeDOaL++44prDZElTSp3pa2Qr
xIdYVZ34zf/GlUFFbUxbRjqL5aVWZeKnZiaC5Go9+60hQRO6tT0DqAXIJiVOBRCV
AgSu5SVMyp1J/NEj5+3GJdJCHWF9BYitXsRpnmU6ER7LZogFj+1qIQWNzPErHtd2
e6+LTDnwnoa9Hc1EZfgcrB9vK5TG98SlUYrtqxghtgKSag2lWbhkl+EPG4xa5tO5
KVar2iW+35DWaIMxvRrh3shwwAKef8EwhY6q2wE4+9FMSip2IED1s9v/bQ1oig/s
MLiY1JLoAh/S5JDahopC1qaorLwyHPVoc2h95g7K/74xY0gZgLW3KguM1MYJ26CC
OeQYs/7xkudT8fv088YIZ2OWLeUG1CWYe1hMy8poWPQ3I9i+mcDU8asDUIsliDCY
+mysN24JUhoQkj1jxF0k36gg3xinVrK5UEgqPtlQVJ2Y07MIINTYD3gP96qbx75P
OHQAbnZ6Ta5ChBm7MZ6TFhCWh1Ad2pKEI5HYD6seplDhi4ZQcGOvkDu0GrABe2No
nqnG66g7ynr/kwpOKzZp44HoH1jWQikzWA99gcE6LgLwgF13s+qVTjIioLe8H+kF
gcViQ4JbJRHJE5xiN1Ql1JjdLq9mszPpTMPvTeH4mkUNiU6mJUuaIUgwHD3AUilJ
OS9RR0XS6DoCVtYZnE+6NjvoZYTuhbV1wpP1wdA41vevf+l9Dj9PFNyobrfJfTzS
GSGDF5ErbZ339dlyV51LGiRYnOhuyZ+umdWWpxiLQidWseJZ4gP/5yyZasy8QbX8
zfy7jZX+hXfRrNwHlzYHPXY9j63nT3TwnyNbeYYiOAdixWm3lbqwDFKBoJdOKfOc
tkJRpTU2zTcwXl3u3rfqTAYpCXgtfESvx6vQfyjvAbp5FO0UwZnY+duGecJmx6VC
3c0hxsKNfuy8ct+SUP9EIKPZCVVs6QEANeUaOO8lfwNA6+qlqXmCH5P6r8tuw5wq
5IFXjb/P4CBKD03I44DNeOqczyrRMJYbFIG6eIg31FP9nA2RHwUVWm2Vqm2L3lZt
SHsk8fv43EX00ZNlofk+BN5qK7UxETv37LDwbC+L0i7wCGZV8rxf3p8RsB4EIb7W
s1Dxj0vuxTzzTRUf7Hp2/SyoTpRyeHlWCJMO0Wm7Ft3SrIvZvAWV7p+wjafQGjM1
r0R/wniG1rS6KA0kjtiiKBXPgZIJkdQo+c+oe8BFi2K2qoJ306k3X/gPkJnMAIsC
VarKgz2tRokoEiLXtItedMvFPjSsLzQBbLUayU8buxUEzQHhU/7k5KF+rWBLQUXU
wA1ds3eqPdb/dOKvAekqiHK4FHfl5cKq3M5KWdGCcnx5e/3iYPDA8kpH8GnW/5b5
+TuBdL1QaMR1JNZxtv6VlZljKEYEeXYdD+gfFfD6hhCZlg2n5FVbv+WHlo4Efu6f
PdTzqnWueJNqMKOkDFGPrTw9f3WvbIG23z3mbJVKGx/+nHdnHgE0zXDkP5EOsHby
Z+Kr+cEL3qSYgUfJ7162xtigTGg7/4NdTbnjyODYPRnudbSKtHpLgWR6XQ27HE16
YugT3rgaOXXZYjZrl3bklCotOciwseJ/753EA3AfHfl87NtBPn+gtA+/+m1XOhLt
D3idsNmONwd2jR4Twd4sZM1htkTHcCr68iHfOviEHpaBwSl7GiA0eNjLis+Lv/a6
VDaXRFZDaD11+QVGO3mXq4vUA2UTznHwkhGe6MuQxtqxDTMxJUv7T3ixZNV+D0bM
DQz2RSuv0RKrnTM3OuA1F4b/rR4UOfsFh0NcwnymztlW2Oys+vzThgNnYp2tx1+l
e0dQjzqPZ1gOSbjEaJxnXP+R4bLTGSqTYTmKgk0hQ0J+gon5j8B4ZNXEyCtrLd60
zOs4Rc3ibg39VrZEKicT+7fgQ0dPO3PhJdCHvjBdxzpolon3fvBJ1BKczRsRtrba
34og94VV+6FONlUupMTITNQzm9A5U3/MqOyOTjXqwGW+DE923a1qX38QaBNifsNu
VMyisf2cVg3Ne4k8ZuRg2/gtlf+TsuukPfRCJcAwFnHV9ZfCVmpiJW9CGmZqrYWE
FA63Z9M289GXmRPGpo5hrheEva8Y1Pwb/zS4Xdrt1w8szWLjzzcuGsS8s2BfRfHd
LZlvgY1Z36zOHJLlM51UOZOyaEahchjD7JuCq3aZX6+vzILgTtOIgefYr9KgM8SU
XExIxvMNxX2dh6UziC2IC7Te4KcU1A/yGscNHoc+DOcKWV1e/d+Q8l2Z29ifnpa6
MSz6W7o4Ho8wAA+WMHQ9V0OS2Z7HXH3zz6oSCZbBsjHK/+MTC6maOMAhcKia2qEt
3PU4HA2yDb/PbM19CmWkjxMUUV8n+lf1Adwzgo+EPe01AIaXcEmleRO1c+PLHdVF
sCql3J4lE752eKu4dVvWobMhYt0YD/acNizDfiEcmrY0CS+Tu+qCnOg9i8wmcCR6
J0FtdS6AcEKxHlwyN6obdnjZzBkTkWbrXzF4cnAXRJN16OHOvEdPISfyo6ZZ97FE
9LPHc7ZW0qcyCI44AIlJ1eYaWD0kJRcEde0vXGK7xVSVYh0VAzQeHXOSP1BJByWZ
XafXnSVH+8xTlWnDx8xaQ2nG429/MPe+dtm8TGHcAcqwPHfwupiUWXkW4hK4DHed
Ftd5XQOirv/8FTiRvngZ+2y69PDrBYcsGGedaybvz4cNi8EfPkdWd4evCHeD1HGd
qLbfxnJQhU6+UTcLW1LKorOltBWHJCqy5iio132u27Cotwfw00Yln7FTokALpRTP
BWwpUZyeG74ygYEu0ftrLG+JiaizPfpbrVzLL0P1TpitiUqSlThcGBVTTURCf3Xa
NZVCue5kJuv68IQx9D1w/aDdBG3dUNf2W5zdXErzSMtsMxqbMEAGtqe+oOv9n23x
lopE5q1yJ9vABPdk9B8nUvAbWMkH0fbg1MTxWk/ZjYb4M51PEY5zc7YuC7YvQz6Z
G7+kRBWIVBP5LjrLVi0/yYNAg1Tc+oHD8tgJMmnbTvhxkFkq0p8sj/ztnf6Du64b
n/jZXZJITLCqng2wV1/pdGYEvE4Rb90bx5lHBOTEvYeFtbT+kdnUIPJKgXMCAXzn
UI5QSiWvwDJHkaJsOjyFKHZb9YdKoJE+Kv10HYFLOZn/qSspR/jtQyH98HEVMlpD
YG1EK8JVrOtbjmGq85BBSh7ifHEgaAUCjvwx54GEQfY4x67JEVg7/43YNIFIx2ry
qt0jD39DBDTI3OtWy5UjM5IHxfDywIiUWnLiX1wBrsPFPS4fNrwZuHibFqDubOdI
k69kB7z0svtzreGmKjoBY61DsVJqS1kGsBtBL2My8L6txc9ezikv9wGmEFtf4ckF
H23Jbkr2Y2izwb20H+fB0WRftsuPgQIPgptHJv/SXEspzsV0WzauXds0f85eh7tk
KvBiY7JC7MsAsPZyQR2wsaFTj200ikHHRMLlbfiprEP3792ehEMNa1oJD/CMDV8q
bBhWouIm916tnIPnSdLd4dTX9PqiEG73YoQMgPTnvBe/vaGyQlFbMX+k3/5gjakz
ycj9VaydulldHwbNhfqRkui+g53ToUGGj0jwfZGqN1G9mut9Swemp44XINhpPXGw
l4SW4M7bJvnH7SjxLf4o1s9zW7sqIno2GNkhBH6QVQRzC0EUpmCN8DTYXBrf4AD7
B2rlWkWmXrxO5sha/vB770ed+ZOcmj+wlF3D2hQeKpy8BKY//Ow1Vn2JvD1xcWxW
vE8md/aFpyCe0gIkV8FjCPNBc1PYlDZPoUBQD0TK4fSSUnnLYIDs2t5JrMkWxLTl
ftt9czCr8XzMk3BMVSJruvc8THmg9n6SvqdrKOGCsFEqRIrjmSLn/Vyy3y14OamP
+d4csPEmkCc4GDUfGdQ5qnW9ZAELjetcDqGLcng9zgFp7M8B1D5SQnK3lDmLdZwg
YtV3mjwQmRlEAsNPJH46E0l/Jcvad1nsiv1It+1xnVFpwtGkFurgFeRvIwQp8nYH
3WYyBle/VONe5NcECH+I8mitV+6zH7MIE2GUZikG4LAyuB8ds3A99CrvHfzx1c4S
ePSv0MGizKWcmgHQdGowH99PcfK+CgDwPob/pcMPkQxRsGqMCWwzd0J+WvGeBL/F
BkKneAQEre68aRgCF3Ue2lYMM+e/fI73uo4bYkr5bZ2AnWl+VrONlQe2/OixEFhW
iJkQhD/TLdCvw010nbKjk6q+TLXwkyK00TLc9F79asDmmLphO6ixnH20I8iynw7T
QoOoDXC/6K9g1gL4QWOl+/MmrlWGTGBG8e1eZWKIYbU120wWEetQNMTFrgQyGVga
tzv+LcQwHGyQ6LpuvWFj+3oPnGvAdTce6zhWIMIPsHpu5MVe1vVkDG/msDNrhF0e
qzAmmGivfrKA6RCfi9562CykmzyaaJvIsq0PDrxf9BSVTv+w7cF/J0fkBXwOLykE
EqzbF0qHXg5TlNyxlA+fkSsgfUhVe+FLAC4ncJGZUIZcotxg2W/6XBVPqev+j8xU
2AfL2mwHEifXHPYg8sekNGPsvIAl6rv9XjiiEnRfs9vmoEb45JIcH8TmWlbRHSUy
SzIqXjyqKFBXs3QEklCHc5AfeIYgyyU/HE3QJdXMpnTZ5Jg2Y9NevUpZqVIHa76e
SRrnGZpkVgXGqI+kYuO06EGGn1W1P5CHMM8wrEiwmJTKpwloQjxXeIrhz1ajvO7n
0kfA0nDZ+HcrrkcxXU6CrNb2Eznh1mjJQxzB8Ih+3MkempAaIwdmdpxvn+QaNekv
ksNsTBnO84X5ebGfFmqxkfO/xh+YSjycdtg4f/l+yrA5wtIMJciUK19LjmymDL8U
O1YksQp8ELT9Oe4XPhiuEQStkRtbgd1+F+kz3J+rgWCikVP69ZOKH00iW353YSaj
YlOQSI8cXX6K24hB2gTWmiEyLBrtiIyUkh29xxrNqlFzozVYejNAF3jmuwvuf5tn
bCBuxME9OD2yeWA0R87uo/toq+ysl7RU8PGaIRAFZQ1BN/4td565JNqQuZ9pznR/
oZpU1dl6JVx2sTDC4WFkHJKCy/7dnP5z+nXaf44Wy6QuOpKDd0LkEH3rxI3NCAXh
HLn8xfyFUokyO5UGQbkzl31TFfdG8BsNXu7DgyIdv658vD+h571wLY3bqlroeyuL
6b3mS9Q4stbVzm9ko8ZkhkMh6IWT615r0O6vHumNGK8CW5HONQ/8FKQp6+fSBvcB
HhOWooGjr+gb5zVaYQw3KGDzGmCDulw0TqFhQFfmQ6WmmHaGLZuDG/n3kkdIYLUV
+0UU30x0HxDQ/nSs+SBEJoLUyPxYjjHUReJWI4+izzICjgY+chM5VlKG9KqM0Z6y
f22gVV0Ia064dtfAJd+BYFFTvKQkVE6CRuN754va3GDWbMhNYW0SOA/WnwtAtUjn
ZZBKxt7AIgJwR2zeoOw0aUjIbl9LaRuhnUzFAuhIVxai5vopnVQbfcL0EVXCGh9I
FDUgm9E2gJcbSexngLIMm6Ty+DvlBwLRJqornXyaOf23E0luqNneC/TsQQo/Lfst
YXSmrJqzfuj/JY4hNfPg8Ji9/8MSm0USFmvaEQT7OzHfYi9YyHzLEnT8d5lNfrf8
kGSsOsovwIBr21bs6lSNZ3Mhf24oLex3qEFzFnZ4sGtgRpVO1dBPFGttwlWRUw05
whgT9TkTcMlOZ6W2xpvXiPmlfQrItd7jTQP3mL8ByvQU8nSVYNV3XLuDGvYTsGfs
4IVKSAUk6vmYDn7cK9a47dhGIJIjvuewrCojQ4+QvCNQushs2louy9UWQ2v1MaOR
01fE996A5FxCvCQx4OEAIH9scmby4miJ76R90NTLVKNmx7dTlfYAzYX1I18NdGQQ
rVXwXKQGVgTKIJFYNgt5Fv1I0jbz27ldGSn5dTIlTMfNRgnGiTRp707rcaHZ8BEr
ToKuRC3Iy+UIGzh1OwY4fDlPy8SZIqvdIWpZ7miRAdqHUcW9WuDcxMpuTsSv2z0k
ZfOAnuxWNtc0KEL1g0BALhxyVH+Z4EuG90Z/EKSGERddNJTceJSImTInrMkRI1TE
/j5+hNU0LQkIJsR4E4w/0M0SxO8K2hcf//bT97tU3eq24uc1wY8xifrivsojGayB
/h8TuS/pBaYg01rvD/Fyhk5vnNKsNsCnDuVeSrcePX+boXXpOP4yoDwI223pN+nr
4SLBN5Rh3ikTXvu52o/n1+JaPyJy2/WE5/m5i7NPQghGtHWrg2BEjv7BN7boROHr
mVL/keJ2XpRcvWZc1gxJX9FQu2dHYh6uxxXt50MJcRcy87pdwZGmQc+zLvZXDbcB
+lAxlQamJxdTNqhQSFlmQzIzS4vo04UsWLQ1DAr+Q5YAZZWGj88ryCwmOyPhDtuJ
p3P9UhmO7joOla1G13NJ66FUx102E6sAksqP5lvcCe4QffoOojyizADnTRxsJ/Uq
6usB8IE3wDfbiMGZC4qBa5VOwn5VE7DO3Cv8MA612DRRM/fpreE9xk/ZZKrnzWQg
tGUMK61H4LLQ8TJFc6ybc63rnNjZRBgp5ArnbY1oEex9ZqUCnSLCf1TbEzgsQpGO
Tg33sHy8woJFXuQ951cE4YOzm8Y3oef8Od3SHdaYUadL+XohS8LZM/r6uP1DlI2U
BmfFjffERFThWx/B4Pi6zoc19hCnK5ms9t0rn3LV6DugNYdqTy17DFqWNH8/Bndw
NdBqhSGOOMi9pfLt4V41iczG2/Ro9/KAWs46v+1UtlT1Rc59rAUjKDGlgV6ZQWTV
wtD7R1JX1PeJU4+RHaHe0h2gTN6KxJgCN7inoNbRd/HnKu9S2HdklJDkQlG5wG43
JqmiUnq8BceUymj1zR4evxhVef75p0SQf/gs2e3xP6GqZ54L/g20z1hA69eTwRXa
Mb3IniNYyQh88Fq1+VLNhugSrLJ4kP/nLl2PxhXN7ep49SeFhiTn+ZyG7YR9PU6z
3T7QULkTRebILUSCpQ4uraoPctB2OsxcSXgkIUQCpCYyNGjfdbchtmPGvf7YmxO1
2B7lXuvWPiqEh7AmPerwiiu3gWc8qcO6Y77Q9GN8JKoZqsM+azPkFASBDYNLi+6E
7vldfgSAWDB/Thr2n3uBEoowjLNNcVgFmUUqESdv19jhfWxQgOp41LY6QzE1QkDp
QDeBsDrY3I4jjDG+5JX7PKdDwlGQtJH6e+CKPskaIaMC3TMu5pA/g2c8JMnJH5J2
5ykRPP3z2eIzeiDWpoi7fw7DmKtRRUsVKwl9h9muIftt49sXD1LBgqYs/q2Zynba
FzESKJjk+a2BzetivsU9xacu2JgoFf1ZXnvzqMIrGcQRzXBoaQTswhB/sX5zlCuC
bJu+LHyBIMZxqCl5iImfpPDmPb2QbWvqqlFhMz86DQ2kJeJ5uC18eEmMb/1/CvLd
teFdjRwxleHQnS/vXJiw6wJfOeF5XFCUG/JWRUiS2kSyXhPX0vPWfJavv6tjZo1B
W43ic7Bpuf+ACQVSb0q8iTrHrat7cC6ccYNjbj/10j9KW8gugIKfTdS6Y3bntSxB
52y701bfG+IVU6AxIZPE0TX+roFXoL1jkeIfRwCUWcJzIBPJxhdsgtVhKjMsd/af
iuAII+yjJmwwmeES+QvcYshBq8xdcpB81JD64RKvW4CQNiYwnE9SRe7wQf18YEmz
cn617o6j5/QSNFyAwwa8mLW+BOztcofaRiRGr1uVBd7dz5Sz1BeSHRr2VmAjH4Q6
wAdZ7gfgTb7HHo+SZxk4NWJk1MS0jx5MVbUVBW0spwxwnZxsoOYca31VAqeugjqj
yfGTOV2FbsI0RqYkk7D4aTQHMK/XMzdhR5RNaKQ5ZW1gnFqSCrB0pMIOawFHYnRN
2Ml/myafzDqcX4wY/jiBTwx6nD6l/Oeo1Jl7e78VUXcnT35S/hKj0/l3mbz6V94E
3dmfrhXClJG9HJI4Lwa9rxtOpOpBwAYxF4kWlkf7G/X8g2NPTP7VcYNFckuylRiz
ar6iG17b1FMoVI0vjYPqf+yhwii7PQDmjet0nzkSlH1zRGgQkrrKwqiHw0zeusv5
elH8A8dLuCHn+mLZrQWPokrurvMLoRVY06SuiNmJuLhJn5kEJMbzWMcL0VoL7z1U
uRWlRBzsHmAFEKX29l929PoAeloQIWaMXDhzIbho3ZTk4ihlqISlueCFJ8U4Kx+j
1XW6BHJ/eLzsWJSHGdH+CuLeNeraPGZl3ogsT62p193xDOT165YOXo4tsLRFb8IV
OCTyB8GX/yd1Ief0s4yGCfQ2w4rYbxgliTMX67ajgxhoxErjYqHSPfPVGmH4rqyU
UMnufbmoJtCxdgdZ/1h0u9IzXV3p/zKQcoUs5kndLa2PxGXOSSL2vafOqDS9/Mor
TuA4MxrvHWfZod41Fbq37+Q8Gjt8kRyK0WaOJ2oE3eEIkls013unjrObSc43Xsz5
KkHonJgaF0jf1vyEeWVs7N90bInDZOTreAY2ot/mQoyF+Z+fORV9mu+e7GAkWfVl
USPi7n8KA7zugnL0dJ3Gg6SQMmGN2z1q2mlBdzTyS448c8U2rSngffIsYiGbQH7V
OJBswmntH1FI4b1gV4kzJg1q1Dl2KOej+SEmyWrLM7vq8NU12OTJ+FR+ArFFi92G
vhhe1ewpoMyF3OStTMxKjuKnHKYCayOxYvKHa4V84vL4t+N5QCGHjCCjOMD2eltB
MMgSaHGJu6THpt2tuNgKpOmq2D7L+FiZXDFz80AVAiijgSNNRyc8GNAqVkHO6Z7N
mIB0ecAW2u+U79tTwd2tdhH1lbFbQDYhblwF+/EQpFWeOAoU7D6fSts/pBVkNgzr
8FDRrC7nWZy+FK/AaZRz1EdchhomhqQWoYgZymr2GJjdiw8lQWEcdOBgPc2JFNHM
2ikNfuI/TKwgICm2xoogFolAsTNCmxzDKBrSE8UzXibHmgiyIdrtQ1lWL5korYxu
oYnSE5vZ2S6k+d9zdx62FmQnhiwUDTTYwG+LqKX9zWKqhvwhkO9np0xZs9DPwyHX
kezvjnipLKK44kM6wlAHHyNY7uHh0SvAEmzKORGxCNSbnq3XyusZNqqTBFMxPuyF
x1lflh9ZKEmqtPf0/XohAzJsEe1IsdrQ+SNo0j3zDqzK0Nd2xqvv9XwDK5rvH+eQ
WaKS2J8yl2bhV5nCAQkUXN/x8RmFbciNpzLACCp8jXltnB1MsCwdO5RceRbcCEa9
SWdav4bfnSaRMwq4KvirINo8gQ+m4gvKCHhjp7e0cBCgx1G2ntdhIHr0sH/LdMsa
1H+ki6Z23lbamxU2JfSRxiusTbeTa9cbybUNKvgNSuzQ28Wq2/6QAllpqFWoRkQD
ji8t0Rd2kId7ZTI52uGt0Llgco6H1RVtRVlMR016/yvom0YikU4FsDZrKCNYKCsC
rtDW3oAOnOjxkPM/viP7BjCcH10stibmyDrvVxQDRs0sWDk11Giai74GzUzArqFd
lrMph2WkC9XkF6pe0ryBB1PvrAgqDUQy8OHHXYgVWBoX3uOhk2mJhV2UphvO9Waj
dEjJKPPUQKnyCr60nsga87Dub6VCVWuiQv0bOgFuaKpFWj6Fz7wmzRzPxd4xj4eM
qFltZgcuBqsKnULk3oPZ+aMZ/nxPyCuCCW2+blu1E37pC2yX/kOb2yhK9cM9EeCg
nWbjwHvzZGx6wN9dTfshMxUrKYU86hTg1wDm+GIWeIesEf4T87jBUNoMBGJnWqHp
VLfFczi1NO8Xq2NASC6HtnKIGESPNfWrWjawFEcM4ih3YNCYqtCnqbr6Q4ukgNKO
itdKxMnXAepC9qAWSBABUO+Un1J6m5CwhHjK6Z6KrSKKHv0+QKhZm5Z6KIXya3ku
xBsZ1pEvBxDpi3npaXute0ivRT72squEGasSS2sWAPKznOXF0AsuM+PwoHqU0oyE
dV8OOqHqKDwWBp/TggM8gbQAET6A1lGIfAP28WRipi8O9JXJ72znnrC6BbPAQKkW
wgpGHf7CV6btng4iPzOrTQVYKV1HXwfUk9Ag57kj8r4FbRQ/5Se3I2Dr45EqP8SX
Djo63hipUvJfCwRVV3j1eD0tV6QIQTgcaySsDmFNUsVOVstqx5iD7b8Brn3NQQ0J
XwA0Ni3+tgsGcTUgGozmiP98n05YXQwBvM5Zhl/aibwl8ZCqHLeX06nIWWT2zc8d
BsX9SOUtZArqJs7bclcKrNKwCu9nOxXO/4IQ2ycd75q/gc4C+onCoymc+1z95Nlp
mABomivq47diQFnHEZCs8jMzKQLymbYwd2YZJ+j4OoduHeolbKs47RRsOwrtc07M
5JMHIQ8/JlfRzYqse0ARFpxmvLVfXRUPdThDP0qeMHvu6BnOdbwXgAOMrnDLjn9c
S74+qy2Q2wJq3L9ZtKTDCHCOys2ORzzG8oP2Q7xtLM2QC5CA5M1SqMP2C9DaVetz
wl/NqrA6Urns/wKQA15cAPr39LsN5GlXCAx9u/7wDSeuka8xSbf2rFk3FeDT0j+T
fVyK5PBMXqyUHG5gkUpdBSvSDBPnQRfryTnORLd7WBH5FQ7yWQgqc8RWc/o0Ggq6
1frV5wtdMh7Al+HYemNehl3RZ+Qrbpu8MJTnDlSIYR5GBzihAMGUROYBNLoXpiw7
bsepiICk9CW0DMo26v7U0HQdcoDkpiL+AifB3EvgEMEDtYWjS66rOmT450Wfq7/w
rvhvD8Lhhk3atSVBjvCb7FhGlMOiKzX0NRvYS3VRk9moAY1n3nT+pBSm6R/RN68P
xaoqrdpzj5abKiG+XMNZ/PytmDD/RTzT/dwX3Zv5QEfKoMCwn5G9tUcabG0mAd4Z
s/4pfP+UF7a0DeUHPmk/RwCFMFcr1VC5Yxutm95NRhEs7m1LuhoRDeNg/NHweInN
og9M/c7lXnmw9vVG5EJpdGz6CSBsjKOJbwECE5x73HxZDug/kBzCDWZ16x5+FKQL
lh8BDeLPkyRVGlMXzh4Au6hn56ZddZcVs2e7otwRo2Nthurx4E8ANBlL20lLVs+Z
E8LUGwLMF0GtnuYajs0WWE1oKfYuimBCX/puT5LdJJXhOMYL4xbUzL5nNkjm6Bfd
0eeHGS+08l+4mwCZdccJI/Ln7//4l2TmOu5Ap8OdD9mWs1MXgwNN0wfUp/l0QDIu
yPHVhD/9eWSloLu+BqlJasMh66zJmPW5syFz6qsiXzmXL0t/30Sb1+TFrj5kEZQp
1FROH0MqlTsf9sD4CQOwnGJtPIeFoXyhvnb5R8MAX9widfL+otfyJwZvrapFL1N7
aoefeHdmTsRs8IWTnTrCgSmNHK0nfB8ueiS9VVKSJ32c7Ai5QhFv3kZM+y+2M8Hj
YIBy3mk/IVwwc0od9AhjQFhd4RdcdJNOK8BpB/saKC049BZ63WKMKesJ8BGXadm6
ERHi7yazDjwclVk9Yms4V/Vm6OqjlotDFualfGQRIOgjhBAuA6eaOddOY6AS0qmz
0nl7Wy4ZExpLPWzbmTTyFzaRDCVtncKazoTfgV/NB+z/opX+DtVuDXVSdd75BXB+
Ac4C7lmIH5nSwOOoq8VDiBqjA2POyBmyPDj9RKpHB2foaO0WO22I7pe9QzEniZdS
swJsq9bJ23mv6rB6HYVTvLgamcVPF/1muQ4OAqr7u1RAyYwsGUrNpEqJFa+VwMWC
UV54DhlVt4vSr+YPPlxiWf7B88z/0mjw+L3xxMr3CxRE/Z96pwfkNMMmPSA0W7Uy
ybjJt5uX+tANVt/WV4FshO7B6tCkD6ll0hOlea52BQDsTQExRsPuFpNfQxpfx/L7
CR+Ig1cGC5EQlZgx3JJU9fWiZ6UsUDukNOATP8ww0r/5AKrl5SxGtHIwem/acPkg
JN7g5fGc2IpoVnbFdRvNRW7r2uI0dMPGSQyyZeqcv3MjHnn91CU6CQky0c/eo+p+
go3KQ9YtDIIe7RPbKc9j1bL+0U7bCjuUBkWz1zrUVN9jjMjkZpLmI1Wn6I3oeKr1
DnLwsEk6A0blF53kW631whdZeq1f2XWatYoO0WbJ64wPR4XR4g5Hv5jbDPUh0H+4
gBeNolbtTaOwKWc+9HHFjaRRQCvRW69y791rf2nwAnaYGmcwQog5NvFaM4UNOqZi
OWteTDuacAkNMkSUJv/6ha2R/jD9WTxxbUghcT13yXgUGba/Dj6BsKcfPCCSUlzr
I5j+4tw4Pcs3LIfbywsMi3WMkFFJylW/ph2gO3YufeBxyXlmbns5DoZsvL0BhLFI
wzjvJJassQ5iTNJbDQj0AyZWeb9+dHIqNsUc8FO1gyk5ihUWxyIAnuwCKIYYsFjh
uHwDFb26KoZofMw84eWmyHafUezQdeEwlmgAP+93NgJ/4dkMJozVEnI2M8pRCfGI
Bzd2qFqsAwc+bfN4CE7SdyDwOgir4cpzLN4E4iF1KR+nkGLUYxX74yfnK8DTSEJL
aEzjV1Xflu0xiDUALHydAhTAkGLMHWPmJHfALRKdCwa2FNvaPFyL5JLC5yc32sax
GWRr2KyHtp6avV1J2gVRz6HMY33a01Lsb4xKamn/9d2HeQKk2O986C5uNqS6R711
aAr6BBuNHzlk2NdtuMKiSigWDA1773bMks/tlcfaqD8/ax66xAGcovG/5YztZ71L
YQ1QDUNAzd3Z5F7KUi3IawKwKNKhEc4MffF5rRitS7PeEcLVGMVqRcgzj3VHTFjJ
dsuOQyizcmLdtWfMWuQtJSQlkUPuqi6hJUEj7Ii+3tu/BdigUVbJ5eHoPQREaSEt
hN8ePUotCFLszrfQzoE8k+3GZtvuTGYOgXaIW+6i2WPwdXLJ2YH409MV//aSQwEX
N5Cg0eJ5IkRcNwVx6SpiFUJMxa5K0LGRtBnf4f713iCy0Sx9HfUWmNBsWeNPyIgU
0+0BAU6AFxdCvHkfyfh0j5z520QGlZqETq5qvur1QE9b3N6utONfh4u3YuNkKwnX
1mFmwulsPSDZKVIA/zeSHi5HpRKcvR9XF83OoxguA2F3ac+mF/SNgUYB0rEvfC5D
5dwKvCNOZdaDMvBIahPdCvon02x5n2TV5tAi39c2/0Xd8jo4YLMmQAdYYgMn5N/N
ltvhi9Y3I/mSBixS8ANyEC7XrfWvocQSWkw5IgcL3SSwfQHpkQJq6kNRvxCCYZsA
`protect end_protected