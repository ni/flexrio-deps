`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
Uy4DmKguuKHGYwV9sMd7gnnNEVLW9+X0c8RF3AeSDPX2LQlDvSp3Roqej+xsziIf
elteFIK6HRZJjkGs2TPpXtzASg/EQISNrnGr0N8gL65gVPvfzbPqPxgleuL6KafI
0r5T7/epK5OzG8Is9ssd4iHpE/ppcNUMD3caxjqlTFzbb186Y2g6AV1tl08AFtCq
h8ocsNYzLMQpxdtoINgFqsWOuwZT9SFV0BPmZiH6DDbKVN/KtqVdI75s5A9y1e8m
orlh1k7OVgDaLAfi9izIiEZI1BFzS+AgxQVPN3E4hdn4kiHFc9ihO4qEleSK1f+9
Hm+fx9H19jgCjr8WUDCFKBqZl+bqvAsJpWG1/0pS2ccaw0LawQGR4PoksgER6kfg
uFWbgHdnxOfsoCKhj4Qoo52hDm4FBQzZB6CKBTS10evUECEFMuKXhGhV8RT9Yc/B
+K31CPN4YDqoWR1e8nQJ8Z9txN3ZITvq/8jiT9+dgR8mMer9BU4NOGBdrHWw9hGt
t1QXCmN6THChfCL6oZzPRn6jZ9Ny2bT/Kor8saoAnfOiOBIc3QGFmfBidMwDTdAv
o8P3T7OHOLVkyJIq9oJi7A9jCGjDTvBW3m+RlAVQYVT8NmrTvTnxs2SFA/hgLlHK
My0Oom1NvFySw+SBcLZrFaYOYqn1Z9mid886FOBCU94au8KmkZuTev3yEsILxn9p
Ql3WP9SPdqUBJf/2fUWEccYePmC2HMY7R+IU+MkRbLwStVqNIQF253oyLBuaB+MT
YGWhhShWkpiq1S55VcQ00+tngjDfAWLZiNi2DUPhoilpd+S+67zUffQryx9Dnxjy
+3VecydgDVt7/1R0VZz1eTPDLgEE9pnyzjF24+Xft2V9z2foYMdAh5cS1LDbN7q8
4TR2nRlazvyf4M3tz+S3A+azkFqHrHSfN/Iy1rMwCxeyIff7adtQzyUoFojsoGL6
zCtZ3Z/5hpdqBq+UI8BxocCscZEC/E1/dCennHCz3+4KMTF6icC/4BJsp3wfvggx
3G8MzC64L5LKIVtuLlQCtdwGIwjRr6flrLN4YVIW27Ws+0eXWur3TM16WeWYICcQ
YC60vbySMiWZ/uqZjpgRhzwP9EYG1/pI4PBOgY/B55WPyQb27x8olSp5QtZzSeRC
rTeZRfU5aj91w6hUgh4IKPn2wKpuhI4/S411qzQ5kVivxtcP5NTLkcqYgk1Q80KO
+78JP4VKBMuOx0+nF4G3AViZxMRgBc2tNWIyUvD7Y/xtv9QzlciJDMLCjCGSCX0f
drgD+e0OxQ8+7MYemhbK9NNdM8Vni1ZrBX27QNiqWW69y92QQx6Ijaiwu8tpZSnQ
DV/fy1vzGiWdkD3QL5V5IQayPjGp8vF6p2oRRKs6NULRaMId4uRuRQlYqOQfXiar
WKyQ2UUKw0L1oRvRTnr4r7PKVKhNKcx+j71FMe80yka28D/2TXDoGCRUNmQdc7f3
43jM2iTuOgMPMhuFDkqMT33OGtL2AvyhhXqGmSQ8+vx5VtJDHiTC1WGy8wyMLdDk
DZxLBhbhkjnAyj7ZICJNtQU+XFPa3BGl9+hepk14i/R1O1T70f87vbK03iFjqJg+
yUhoqGb7TBM/PLeE02Bwakz8IRer/F7cHtfy/fv9rFyqDyAmgd2QGKyKqaKqJ4be
EvGHs8ucWuC3KwxM0Zh0NuCrFLJuxFeoufx8RF34AwzhxnlyDh85AccOswxJdWb2
7EJ6h3m8Fegix3fH15tiVQ9PfC5Q+LtCzlvG56im7oLTwQzfgPVWYfEkUc8L/Cfi
UnDqg/4UKNO7D+QLS1sdpokxtaADI4ePto2v1zp5/7tiZwhL0VB9lduubwO8CCoa
6qMtl4m17p/wdNQ2L9zBgfy/a54huXXbM36c2LTlhxMhw6eRuuNPHttyVXJNuEPB
AQ7/MD5+lpv2tnuIKzPnY0cl0fkM8CNp/LLUBCnoWRaq0sWnbYs/qr6MFkEHU/P4
kodMpd4rtQDPwKZNz8zXspGxoa1Fmw1Yfd09orwI7/I8N+GZheFgUtQkjQXOv8xm
OfE2KifFFCOvb9BVz+aC7c8NoVSRw557Mpi6DKB81b5vaVzlMzaDVEaO4Um6KrR7
yyPGmndlC2wdn/kDcYL/nshPWQ6HgTnkNTUak0ourXGBxc8IlNv7PkpOt/8tZKJ+
ks0oZoTKFf7QAEk66XqT01D0oqw98b2RbMYqpwiHyFxKEF2gDPwNOohUYGmtRg5c
9aBsZU0lVk3q19RM6nYMCYwcWCDdD6mPoNzSzPR8GsflRhTHm+0F8fYxzUgJEvO2
fbqGTtcbV36+Pb1+AG1F20EhAL1pseJrsLvIAxlYr+zhITMUz2cYBWnCzP6gJ+8W
yuc4+ortVbieISqygva9GK5T1hyH3PIH0f9GzRk1pg/RVTChcLxu0hJuaBX/cfIt
SEs4DSmMLtcRrI6bRpjiKg+6jK+Sr/0JX/6vX6l21mlz8qRU8KFt4WUEbOYLxlx5
3bwft15pYYsu1uERoLHAWDg5LGH8pHZzZJzGpgwShgE9e7PWFasY0dVwMeqiaDDi
`protect end_protected