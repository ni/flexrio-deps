`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11232 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
cjljSPzTIRTXBX/bLgom+fTL6s16uTa2x/Nz9CgPb1B1WfnIFbz0zHFqzhjIM8KN
edbHSi4IFzIVF+D6+2LYD4Rjm3Ix8W5EMJJ/7t3tIgCKhbyG0OyuIASnGaAsHwaU
if3jNdo2vSCAH89agR5ohtEk/tWoJU4SyJxfJI0VHRh1tZVUqnCUfsOiaBVaBFd0
g/0z7P6llIzcGyDGPk4IHvGLyaBAwjUzKLHPa0QJgR+/0HpbUpecqzLwwQv2r++a
oOyQjOck3WScVNPEWHMtwvjuKwyl9fn3+mnfRO+8Y1+3iFaQax5Q8ucegvbNZxgS
8+bGD/Q8PjTDamA7GjUPgxBJIPBmYGVz03IxALjY+VzWuDJE8qCuSc7oP2oE9lC8
UD2TtuoRd87RErKCJZwwcc4WsTdkjs790pGervDEKTIJoGJcKhXKqDN0uDf6lVvD
agxlgl+/uE0XxQLFYUYQYpFc3a9kd9kebDQflG+a1OYkFBBuIcnUK3NeMu/NsK4P
d4MP9SltFSxOoea9U7U5guf/G9wRZrgB5Cp13fL5jQYEBuaPSoDkoh3A8giu/6dO
3BuV+zUkgeWHu3D+t5fm8JwBp9Hbxv+y3QdXVtnIWh1kTCpkjU/XwYvFYzdZ5hGC
PHb7qof3cKGXkZ8QCHBqss3hujq8ecOnyOdECd7iFMiR/k/oy3mTzdp66pE4pt39
VvPeFrLbdD4pKfRo8wa5LOI3oGz63/HktLmCiL/ZEvgIT9RVxZ/NU0sSl8Dq0W+r
EQY4hgk1C9Fbk3NKFPbu+QIAORBlvpyldK3yvEygQlJbjMffhzJ37j9NnBdN7tzu
zVWz8bnra7cvLOg4CCLwuOgoiDi5KSKpNkl7/il9DEwBxfde2dRtxH6eyJjAZ6x0
mKHYs75Y9mVO+VDZIxLy/ZXLc55E6ARmuWwi5uolrMgQGjYkc2MqGACIHncHGmmY
Bpwz6Yq+qevjlxwwSjeirFia9sooWiRdTSPphG/FHs12NEBcNYp2+YdggjG4MKtC
5ZQQwvD6BtsfPr+S2fypbiTKXROvSvG4uWVbajCyVm5srLyT7QwCZJdvVy2wbEnu
Uirxz3fwL1OkaLPHiyNdKNEQb4EOPARpTDzzBDFuIstflsXaSEMHE8t8mxUa1zkV
NxwKW/oc6SFgDbbhOGzs5HZnq1EmeQnmWzu84oTsoyM7mr561Zte8NG1NdIU/X84
8Uflpjnoc4pqrFQ1QZvEe2CLZ+X9BghjOWpZ2eP4lNplBX7TCsiTiNSrSkiJ7aB1
MFUEeeaHaeoVRoqbq+na/POx4JSswzO7t8FU64y6C+Jvav9MSLKHU3HSLvBXoyYj
xOo5maMDG71mOOAYgFrEqlFY9ZhqnL9Irerwa8Tu2N8JnCUNDEIZauEmKHaHu5LE
KOfydF0nf+rwAPrXDCXJ2ErOGQfTyVnPWnmYVTiPuHHowwB/tvbDjEzkb/QFo2sO
YmN7l1gskJOu9+G8KMzUCpt/B9pYbQlWh8X1ZjNxp2uSsC5BhNWIhyzHDjTSViyu
dWkCYj6l+q9DnJie/mpe3HEMtTkrNWFe0SDa2zJ8lpalLl/RsuV8vtJv4fDyjm/R
3/39PPeSk3nxMFMGKeVhCu23cE/zBvv3ZI5sH1eqvHCSOTDYgo393CpFfjC7BPmV
5mIVPR6OfEmx//slPwo1ZNv9zl7UYPIAJVIhUmMNUSzoZz0fCGyn53hwGaps+gno
MGlUxhBpUfIOSJDxqYYC2TfUE41W7ldyfUIU7+wR/xRvxH1FUJHtX338JsTcUG9u
tPZf9Vu2MvhTHgr8s5os9Sej45ObDW1nVLlblBzIPVbJJ3hja6smg+KjkjXq5Z3V
iThXF+QQNnRk+EGXhSvHL73o+1WeGS1N8y2TsUd6S2XynMC6G50TAo62RmbStyqT
yHezRQa4R8atHRxPlUJ+prl4oRJhWd8S1/oOy+RMMgmkDtaZtipNxQ7Tvc4WOSf+
k16jfWcjASeQfX57si20m5hA43jx2SyXeXPkNDKbgQDcbWZFINUmcS4KX9DHmpEj
fSPM9hZX606q7yEd8eLEWOGk1j9QV1QKTU+n9urqFOMKJNM5FS5gblhiXE22nf2/
clrJsLtv/z1bodW0lnwTFJjKKz1Tb52OT1ijbQkJ3Kg8wwhk6duRfIKKtc4riCI7
S6K8CypcAnvv/u9CNe1ns1tRCuPouEWJNgaS4XOCJ+439yZM5APCCh/guCfByrj9
JuqmKuoj8GZePzVbmM953Jz1gU+b6E53JmeBtbh7tzz5zNhZ94yjjvLA1N+cpcn/
c/MU7jUp98JL7VzyQ0ljohMI4EY1c9QRageWrhwN+lobBtNFAukDp8yPrnpkaqCZ
IkERzwJwbNvOB9eyv9U8LRR6UB5jXJ7dX1lnuy8sTamTkZVQ9Ig5ihGvSAMr8yfr
6cxGmzDV61zYYccF0bR/6kbUXa7sD07nVs+2u7O7VxIbNHvtcSCNXJ/tGk1JHJnQ
82+daCUwtSZEus+zx84L2D6Cr6ijypbWeT46JxI2l26sn1oqinFIurN2EE6NJLHa
8i8I/R8mRowwdWw6Hw7K7QdIyx/lHM9nELUypFEl7Elh5nWsZjcjYXkz8adUIUj2
fmEK/1sYyaM9rEyMYlw1lEdJjeZvk+B0iT5U+Zedg8CRF8OcqNvlJ3OKWxEmWTVs
nZWfYnF58m1+zZ94LiRbJa0bdXN68bSpwp4sVafTgBqep6XiKWkvUUDMoXsLD31b
7/50jc7uubpNkhAz8nCt4aEjpgv8QhuoZbuU7MiWpt2lEs9NJFehR9WCalOh6HC4
vUULE1ebiQ5F9j7NI1LQ07VHY1dfQME207t/rOAvsnF39ptMZC7XVHt65hKQMBBI
49pye1jUIvmXIPBnTDtgSfEIC1KBQefkDRJUGHEHsiBPJQqu+kvRAuDw7HjkZ2zM
epoEf1W1Hb61mM4D3q2zQGiml1qMhQ/K8I2g17iFdAk5Ec4khilQMAQPr9URyc7Y
ZFAy09DQbINKH3RjzC4LxDSgn9LTwHpt7Mq5+7fnPshdOdsnANKYt3K6pNPDnmiE
lGQM1NfFk1yKUw1u0MA/0imO+zvsQtaCmiW3WmdC1cdKvt96Fidp7kuPLcvM4dLo
3iG7meaJvf2xwelZzyJqS2AzVXL3/qkcnPE0THbSGXw3BcexEduEJ1TLrth4VG1u
CANcGB6MFSbiKqZWDRJ7KV7JpeVqRglGcdrY/UONEbmCoTAdEIOyMxddlVZcGi7C
XWdSg33ByovsXEipJ9rlehhooV+FuamI1EMD3bDOxZKPbisY+Xp64N1kQ0v3wydB
6Hm+8G+JIYaRaX9ChQE2w4LkJbZYiXLrbggclGm5xNyYc1cGri/FKQmwbDluW4gQ
O6UDnOsekRZwfeQSJG5C8cEIqQPBTRiIUrAps/VcEfQE7xcVlepYxvFWvRPpW59g
RbuuUaR3RKwjoE3D6k4/h6RLIkBQeYKPnwiRDZdPGvb+aRpqK1bhdCEvsAj4cGpA
GoMswc08Ddj8tru6l/3SYEH58ywXyDD3qGZ0EX0dKDVmckh+nVyKZ2tufK8qKcKj
f042egM1GxJQw0lFf7h8HyJI7D/0nS+DyRiHPxrNTsAT5eIrBi7btme+JMDuxJLY
eRbF9seckQAnZ4J1+A0/h5TC7bNUxy9alNzS/NCfyNuaF8fPo/i0KKof3n9NGj/V
r38zHhAOz47X8v4Vo98CN0ph5HLEE/LLAJMyyN/ebEzjCGe+CVSwvGRdFAmLIKJy
u7+ldniMcL6+y9+ttq/XAdnPrpCEwFNlYq37gpVYW16sWCxgfdfz8f1iHyV2JEof
FORgj0ZnqJe1wzyisHH+nXBh1sNpHwDIl5aEpKRPspTFUYK8Ck8NuU9RiFpZdanK
i8vWLrpE+aRA59p0Mb9YHPEm40LJvb2QH1utSU8gWJwVvhAJcA3E1yNwudOemzbm
hDqRHP+D4Geo+JU0QWiY6I9bFkJr49kIflP22gUwtFAIQeH3+oA1Dmk1R69o8eke
K5DIqJ1yLg9NqgO1pE+ouJMF79aV5QfmIhQAR0BYrY7/VVgGlRLjKEm5V0BDtgPW
RsfVgFkbsa+LlQhH05uu+ipxUxRkUMSWsJfl0jqkycWyVTQWLtMqX8ZMH70lpXgy
TFEXQ20LkCuBth12FYnrSAaXnS8Fjfgr9M+ecIUZ8ZI0gRrqUS60iEkKJtsoQHPA
HJ2P3sQXlyWKIZhvSCAG8NCCroVy4EycyGNwOxAGuC90Sz0Sbc8IlCJGK4m72wzn
MMNWtjKdS6VTU5PZgj8kKE9V3aZdDYWdzuaw0pnAmoVhARZKiEuh5xOW1Utca4Qq
xFI3mGE3/d+4YiAtXymk9/dI12fOk151544j+GhYMCgxp/3UFCCOwr2laLnjnaDS
k0ap2FoahqI4c8LcErJZwi3VbJrsM9ManqV5qsi4E+jq4PXLnnw+6S5sT6vlwFcm
iBMRFjqcCMpMf4eCGdSY3KisS0bH53WTtlI1SJelxzlitp+HFMPvpbvPGAKakzZz
iz9qFHyvSuFiNDMRsbH2tL14V+aO87tQ++NN7O7mqvSqsLwMYI+wbw42+BMvZVmV
o8l3r7XgtQ5jqIHiRMmIqolFwfRSzHQdkeJb9ASWsx3Y8KxFKzOGYvmF4Ahko+rC
SY7qE9CexHD1r2OldmR1bV1i42hmIyWGa1xNoYcT9Pzpt3nuKenyG3LoCm42DMZT
Yro9TBwFm+cxwIzq6fWV0zZayoiDMKqQSdicfdSUuFgF2HNR98dir46g6tXcOozD
nPN0FRdd4TjtKLvzAQYFbnJ1exKm0J3qy5F43LRk8MxAzYuANjrQe77dE7GksBfm
GAdtDiJghfybOMjLACfeUxnf8wjMmh/NI/FZQbCb0eZA40S0Z2OH/sSH8Lvp98rO
FbmQmpEc8o45twbC968BJnqbTw7pLLDATZehNwJCc6W7DguqtZh93qpLJ21JRw+/
ZeuU1Q1o0JzLQXQJp8i+9A8iLuaHnJztVAYQo0XwWrKFGKeSWPXvgJlilvl54RaI
XTmGWnPfz2vkoYq/G4OLXUX3+oi4dX9sPMBFMMHKEZresCz5QeQ7w0vFNBUrGUFB
babbcKUescOZIFfTPZF01JCuN3ifBPH2EiRxz3he1ylkj9g7ANYzLVzJMopKxjGz
9j/Qvk7xY2vRjfEbP2a3GixEYj4poER1qA2yb0mpHk/9Vgiztmqsv3UGsxzj+kG1
WFLJxGuk209UL8lYgY8F3q940D/Z4oiZeF1b3EzioYyPBQvuFUGlTZciOH3ZBmYy
7wVe7IfQZoa7WC83eQafgsl6g3KSgf0qyiRaqvoGkHXnQX1EHDyff9+rd/EM1qVs
vek4BucMdeCCe0CaN2FNc1xe+0CdAO5oisVgxxZFLB9X8gvagawe7uBM/r0xrwyW
jY0gPMPwNYKeDSm4emXjXF5DpAsJdTG6lAMj6XWhSjz1zCwXRgwzsm1RpJ7m9Vv9
xvsRfV4Rv2tmoZe9hHq5zx1HAalaz5NySfxBGEGY76RE26aLE1sXLbRsKoeFgsDU
/o1B33rOrBa1amYWWMpYvYYEN69ENx5FLIy5EpcrWNHmCB5xZD2C9+Ol0hK8B/DT
vpodlY8fbc54eBO7gvV0QLryzzUrJjcheJO6c8CQp9G2hKg6x0RYzKR9KjIhPGqf
M7tMGA+oBqyp6Sv/J2A5eK9q2uI/vt3XO/yKiH1/fxANdNRlLZ0sASZFOsntj3Tk
r+qP9bphJvP/PLl0yfd91hhwAHKEMhN2ntuQkBUIEwlbvQPmvLZ9pEx1NgpyUDfs
uhAz0pZnQD73fokTApCAPA2aL+Nr5GPbrTS81iu1vuTtw+Y3XWlpf/HXN2sLGSi0
+9qj0Yo/n8dXV1jQkMxwJfXSsgbxoLmk0I3rPL/n/TDVjmFS4ZFfqJ3M7TK8mio5
O9u+bJsqmm/wOjdJSh/oBqOER1oopD0xQr+wjg6+RF+21KuBQLjgOTh4qquPcCog
JXeUplbBvLseFtzN1XCLqPEwXbbj/uXTOUO2tNhc7biRwgq9YzRaDqOqAU+49Zb3
xKhSC7Evp/kewKjKoh3IiXjkBlfHadaZySj1Uv+Y6bTKuvKTRmS0nSuC4mEwzbf4
YpDsWNtLcsod/EDLFnRcJhLeqMPl5FI6PukkJ6/GWfpZiVDxA7P+O3pgvkDrABc4
O1PPMpo4Rrk+AXJJKGsTBl4nBCNYx7y3Cdop8WFKo+fokdjzlMteHEsSJmgHhFJl
6gYk8fGs/Xmz/GjmsOzneZyHiiW9IyujMVZjjNzOPNHluJSBZyEig1tNmVDZ6yOH
Ee1bzT7+nQijW9gke8pmtv6sObPNC5pkslfZIUkIxG/Jv6nDlqYfkrUsmxVbRFhx
SBSx5lxv7nhCzuvPBqt2HL5K5wgkVHS6KNvjrwUbQTH6uM/F1zHcsl6tHZFjrg2E
HFsFKu8My0hyD4cqpfyDiIo6ZpDjxW5xDUcYZjYQ4fk7jqbap5TyhaR0Ydbbixz+
T/Rk6v4UU8IL4D35yRdGqoHhuKffDeUwOsqc+Ev+YggQUYqcB7shsmnP8mApbXLC
f1nAWAacMIkple3qCNctXDxi465IFI2k7rQ1hutrm7tiwGBBhnQns/HCEGG+Umkl
ICiZ1E7OJt1u6F/+klEWDtOPUIE0Yb5aHbA7FH/ap9lB9pBbWBEkVglMDtS1A2Lh
I8Ae8iZiq8YDcejRAifrqg3ISxECOGkKLLDpuVIO43dpYl6SAz+yPHuFu50D6uJf
gFOaQ/vVgRUNTB1DoUEQZd8gap9QIs+TMD9fOW5mAXblnDhocwj5rDCyudU9YgUn
7qMCNG0wKVdEDY0icgmNSnz3WICagW/M3lXHaDyiEbEXB+QFjE5T9Tg0E1UD+rjj
P22Gcmb6YmYFe12cR8/y8eWNYaaU3cqHAr3PppBftachaMAk/JXFzIvDMpwWKkxy
HG5x6gpaapVGG5kZcczvJCkD4vfAglHKHBRkd6MPbrCdNlYuKSc1XZii8WW+xhO3
gPjrtUt3e5ATVkLi92a8OslGgj1BrrLTbjF0MUL2bm/ce97AQHIj07JcJW+zasbK
gA3EVHBzj/sObn/qLtc6WRu2ygdA3fqa0nweTy0do8A7+qVG8/h86AWCNRmYFKsb
x7sH60GlpaV5X0VyVx6vvkAwq5NflmkXTkykx0HjvydTF51Ou87sMLcM64f+Fvwb
5cPv3u59f5QXv1fVfnt6btDGATxgxARysptacMi1ntMFhrc11Qv2OXAkrqPt/pY2
3eT5dAzG6zAdXYRSk2gc9ZgnwRZWX/lSLbnj/3bH2TLv4GjpqPVutS/ZKvdw3F+h
YImXsCz3qFElCEH5hWznYYMfGF0p14RY6tPfV/OvVwvGqh65dVQzRGzayuLoCexw
I+sRYqEmGG6Dw6+8LIt6Us49M13y5j8YxUdrL1RKC9eI7ObWBsGqvfI+kjPNXCUX
4F0C82rSqqozXxd7gW2gU29VN6zGdUVecmEl2P2B0a04LAz48QkvQvzzLa9NnYjw
BBfM2x8nL7whjLjWJ9NAkY0nsGaQHB0XwpUG7BiSaDc1Of6UurhEkXMfL6cWgYOO
rTXPK3po5KhSA4sEgCdwWbVp4aG/VDBUGjoDnaiUzTrNCFdrDx80tHvMtJXVaQcU
S2Ee15igvKAxNqSxzi0xoP882itW8/SUqp93dp+NC8QzFfoWTpq3S/ynE/f6hBWY
CRg9+YJm5+L5vyS143qUuCebakA2deEBsM+UwKBPFo5T0YllkzvfuR7B6VVWkbsD
YfjPWjHMkE2F6j0o0uqhVGc6UnGkZ4tojUuB++m3bfkRiLPcNTUe8fU/4FwIuua3
vvDuuOvyg0hU56EdGvWEZOFRhHdACo4NdmM7mB6OlCsrzco4xloG95TQ1v0qICW7
5RliEZaqnJIzF3OUkKILbGDSvaglpyIwDifd16A2KaMj709h6Q/pzXhrJfLF+IkW
Ie2WC9eUGWZWnCe25xanGchc49xvptrh2KSbYyEy/LzAslcRnkjx8vE6HvVl1sH9
/y83XLcjSASvUCYG5folGMxYJeN54wDaPzuOh0snmc4u3+B0gkZ6BOMoQjOXi4ti
rYFhMq+FIYq0klgdd/Kz48DAP2gt+ySuZmxvLnUAut+mCcWaMQPcr20GqUqk30Rr
qtB3V4Sa1LooAsPlNkvCYrvHQy1DxJU7nyKeFswTOgZwt6AC9HImMoA1G0W6flNv
DjuihH64KVzUu05LLq/cdFRVQJSFfqnU7LJo9TktFdUK16sj1jueoVdybJWHcYSv
jEC3rk5OVw9Pm6ViiJPN3vjnbZejQpHlrXP4I8Fmp91jiFc5aGE6ZGGHh9uRTEAK
bqDokxQiT4fUD0IKHTYf3MdHN+RIYavp5cYfH5A23EG/e81KkljaVjAH2obK+7EF
aJA6mrxCeRkNO7PLUtxOsq4m0H0Hky/2Vkkef83+dRs2zlshJ+Lkvw62RLzh5/IH
IgLF4LB+26PP0+jM5KDZoD7qPXVG+X0XTW9/cHySHs5IJ94iEaiP01WJs1cLLYAg
apMBMY+PAO2Ba7tPx5T6RKjZqhRc7Gem2+1V5BwNQQ0HEikNdqEwu7BPF9/MfWVf
tfpCD/kWQmgmsynrWL2zOcDGcMNFSpAdJoGIzUDvl8mRtdf8wxh7Vc2m2835oKTk
AWe38o8xxkgD0l8PjbGq3XABte+Cq/xZDCilZJZgD0FgQ7kRVRCpskIwrobNdz8T
Hh1rzHgngOM7g7DzSutnGeggGtqqAe0UCuDOnznRB9WHJhCb9j4VkKRrtB2IYKZb
g+20LFDUaqf7xjjxpcwMhtB4xjl1GGPZPuhiI1utOasR5kRSOapQWKVCtNgKPcXz
Cv8o+2LPOeU8KiGD5NSFVLIl/tQCGnw/HVMkoNBmZNPjg1e8m6MWR1wRSaJeYfdv
WSd9H83adsFo6uCd5D24pk92HM/qnF59TKu8hDquFe35IRVQtNoiPsexLScbKI2Q
g/+DNa8MNb/Fv7VwxuXtHzRb+kdr5rckKGzRKcL+BTpWNSRgRniwMBp8CIMAnInu
AZAefZ9hG37e9CmPeXEJ4Hasi2H9jokiWoriV28vKqAbwoI+zfzB9uEb5dOJk1o0
VPRXWtEdvP8KUOfSSqLcLLy75Mxrp1cLNVaQZrxvrwWvL1k4Dh95Nh3EiC8DxynY
5hQju+LAzCb6tulU0VtbAWdAuDEUSRd1U4Zihy2uxsWgE01o/x9iOdhWJ8mGHCC5
Di7LesJnlKCUNncgxj7fVbZXb4YLNlHq0/wJFi4uafOaSqHE8zSDJgIwwyNT/qnT
VcCIay5Qs9r1KozJu32ouHcinP0jYjx4Qp9WGHqkGIA1Nj34h3+VS+8/0DF6AgwB
BtjgX/9O2xrFaEdMdvAtEXI6WMkOwxtlxEGtp80idmIKU9OXoSHIhd8ILlcfb0dW
KjUA9RIRjZhKiF6yAg3MkNWz8cRP5kZQpLqGShc1OdH4Mj7PXC8AfV63YCy9Fzly
rVFI7z6Ui4hlutqElAUXZ5zgkz9TQJyuQ8OgUlZ6x2eUGXjJbOeeIrtPlLR1/Uox
qES/ctN697UDrQ6i023Z7Lh+UFZ3c0/8WdUZFCCrPTX6i8PsUrMcYyNTS2voLj9S
qcWN/FWHs9UUc+3vL8WXRKlvxkbTpjEikO9bUiVTLtbvYzt2AAEWfTfb4GBnxGvw
Ky6t7KqYY7u7EisQ2vnO4XrBpTrXHeP14Z1f7oIO259xDgi9sAnOpXuAIc8Wtb/1
T1SYjIatJJsHdClQBFjnpLI44NDr/zhoft+UQmzhwRlLCv1hjrtl27GRySX0oJUL
rrS//vDOuvXgfqEAUSMx3wkPMF56qf6Ig/9vhmQUNHMfK/AClWSPg4SrN+DwpGlg
aL/riVr3GGNn9cSx+1FDd9YUq8FBKRSmNP/jP3y5Kq7a4mYBQuHkUh4fIUIGAAHD
KE3Dkt5YICLZdJolsPOnMfumknebga3ZbLNtllrfNCnlqvl9ot4XprHVK2+tsevG
I6sbGU//qQNRrG9E9ucKPljdtM3BZPQdLfNXdvFo6Xku8sJC0lF3VvV9pUOuQUep
j0ZCxyxu4pVsIy23XyeaYBxdy3+5zy1eJoBke7slDlR1XS3bWd4QeTRXjKfcixRG
LqQZdvg3W9LnA1gn5LQWdfhxLnsWFMtpghQLeSCLw7fPlJ8As3TJ53RDPBdnGZr+
V377inUao50Hq3be6AosdtEJmIOjdDuKtHSOtcsf9PyZItS00UXA37jQwBnjV9Lt
osVnSdFgtX8Ase+nIqVJwRQ+n6TYQ8qXyJQDwnwVuoAdwmbAxgfOodacMaYsOZZK
w3THY5FOcOMzmU9soJoL89z8t/R35wQOBpJ8j4rTX5/3CsKhEVbr0p1ULtQWCEb3
zV6la4Ln3R072GRz9/ALH06CTYOcjYfiE0j3VjgHILkHxk5LTSCrMOUVTpkQOJP7
RIuwPUhVvivTvS55gholmpZJckPKg9ZRsBXEejjdpupF/ye7n3IsZMnM4tl/h8Rq
2FZYiy1aC06vYl3S8Qs6PtmixCO2ir0Dp1b3N0Gm1D5z87wKUXENCiTMJVfbjohw
M8tf/fUJrh99kTfqH4XyLvrqPLjDSdejjJuO5sfNnHk7m1cuorbgy5BI7DQVCa0F
1ElSLPCQsf36Ozhx7+FefeKyEqWMxpp/xObGQCjMhLQ0ZdV4SMw0BrD/LAKh2Wcv
psRrtkh/fRVnyYIzTs3/YAbt8cOolcFTv6nDTgfNTINJPuqEZqoI/e5bqMtpTw4s
oghdykkEbUJda3H6x/fMkDJeK+z6oTDnInkZzoP01Uhea1MFFWD4ESAYi4h8+wUh
DgSVDaB1uyFyY5TJ3uU+6eNffyJE2IwV8SWjtCRb1DyrAa5TVYEszpAaBQHi4Dii
bEPPObgGZRX9MLvrrCQ/Ax8PUjsxz9YQ1Z7jCRkbrKDmDuQdhVafYd4Kjv9EdkPm
00QRLbPZh2nfz5dXqoaUj3lH2dA28yHf2enhHdAEGb9LLs4I5XAzZCcY4A8ZxgHw
pbfnxKkdKaUP7gB7vcrW4DnS3RPOTuv3keevjIbZShSgDw09zvx7K4a0HnBbpv6g
2P865O6QeebfXUhI0W5x3ekbUrcogPLMhBbE+fXlPiQg8WegovTlZpRlJEDo16yj
/e0tWMRwInJBm/WRGCIfYfmfPbFsXf0Ct+jPqZGD5iuzpNFv0haiq+FUC3AWT5UF
BIrSjFpArz16T1WSigcID6vV4Zn2tQ0azkeEnJZMaezLEtc5ojx0G3uh6bASlFFV
mGUJ/ZBGP5jEX/q4rV2Le8WWnWTpHWClfHCPvQm0y+jd3aiM70HZD9kLVe4xUXzw
Pl26O3N8Uk/u3MKVr5NrLVniJn2OpyiZI9Ch/UAvXf0M95beEpQ3kcU0x0f1lJc4
iQ4PZ/TYFA6yAFoNI+iockdnbilaWfl+sucommmKSvGmbyE1nnEFeA6gnSyqbXMN
B/0pT3lb4deggsH3Ry3As9R5yZ++R9rfun+ZuLCCpL35hyKNgLbsIcdUnKwImZHo
bhNK3wgGIxoaUoEQjsMDQPCEyrGKxf0ZEIIhQEqlQE/dTTVSGSPUUVwwZUfszKm1
FbSOrKNEYDWXJ+p3mq1j3SATO2G72s5KgdAdhzs/N5jdIlHcTTCb9vzvwF4jZ0cA
Y0dRu4uN1BO+jl/ikGL3Bd7uFcaXeEEPpwywDNsT0v6XrGMRRHxeyFg+ub7Cfm/o
OInS/7jx0zCCLbTCwJeedjOqPeTWFX5luBlISf8xWvtGFnkx0Wj3hP91g3+tOYWZ
yyGsyRzChlx+/uaUqeZOJ+V7HGAUiO5aixOVJT6f/taW1YMrqboNw2WeRLoUd4FP
bbEQZt1jXMol+5krWOhxJBMjZmt1cX5JwNMWrjxCXOoVejOXsjjVjiGhrdDW/AuC
k8TlCkf5oEEfXPsL2SWykJ5kQMav5GfnDt1jaMVdPv6yvK+2HwbmT0EC5wIwtikE
yYnc5ePmzobECSvh3DqniV1LBFsBYmNG3YUk6LefI6tRukKbaABx2nayzp0aDZ9u
/sL4QxYoIXsx9ETVXyd2Cfpdma6jpBtUOON1xL1nBHTDoOZDJUAnkyGluL4Gv/Y0
vJ6YKjtW7GYKFYOLXg05VRZGr8E6BYk6WBWeYw5qb3fYDc0UsdXFDNAiWeb658gm
+2SH5hQHcKhL3qrEEMiAtRg6bAf6dfZcHXL6K+JeWkDyN4qNZ4SikHkWECDxED0T
u/gYa5LlmEaooyBDD5IT4WdHu8vO14e1bi7OpVeEU7HE0Un9I42FqxDzvzeb9DHR
INuAwUGA/nwj3xDxhYwg0ctYB5KPeREVil+m7lQ6k64DgPQVP5+bZwAv1ZzimJ4s
WNPxdyrEz/cTDVs9fhEtyhC1KtiGqkLeECGtn6cXbCssgaEgpnKufd+X5PwFmic7
bzewEUE2lUtpf1WzCq/qMhvHSA+dNUXICLX4Xj1VD9rE9X3QwUOoqi8QAM3rfj1i
BN6Wg2KQFGuCluIH/rzH5YxSgSZIkoa4azVv1lmxslaTI+8caXprsAPfWtl6xBwY
2sF0DciyCBRe8La9LdYgYvcihrncj+KJcfHe/dDzN1Q2qpzNPZnH6FqC2dXe3ZAa
82gtXuBjSxDHawidIV6CFK61arCzcmrrBga7LtuXEknipKlybh4HoGWxqD9dIkxF
gEA0VrhV9HLxVwQ/vIvK7fWh6Y4HF1DAWhcR5P8xUbyklGiRA01a6hmwtcKTHY7h
VkMGZYnzP6xhrij/h/gczAXM152/YV0TU4UXWPmGeGGYvGfpG8WjiTJc3VXOKncz
ZAtxBl7NMHYUEz8T0gSut4xE7o/vEf2AKbgcm/YE4uPUrvzNOajHjX/n7KSaCURH
NCwYZppTFNhWRbfAqSkn4M55V6UA0XOEVIoZrptveM9yEHX9LbQEqbQCEcwFAf4O
Md1gYUaQ+cQbw1ZBvJff0z3rRo3CSqEu/3HJgd5yUembZTwVFgAnBnVcK6DbBa1E
9j/zTthG3gpMhxsCExQaeBl+v4umSY75FjXYcFiom012kukC5fsAjzfKjYDTQgCl
JB0dQMjGsbK/X3Y8l9D1QB4alRWAgEaCPtbmrO1YEwjGigds3nHVwzpfDLY83mQq
ook42bARUsef10pO/OCkuXTF5s+AAGkLhIWok4sRqN1eVZjcbya2i+0P0VBuEGdT
44v6rGn+z0lRRRkCfFFFSe2+xz4gkdbBY56GZpWrH6paB3jGdynHBNMKZZC4xI49
dStqZtv1+FMkNxdsahIjObsMN1A1CyCzIDOfTVwyzGAOXEX2BsC9t6j9LlVqiWk1
A79E72BGVcdGXcv7dcvj3X/PHtjJkk6oLOlY4OFSfKAlpY7eigeBFt7wt5HCiH7S
qBZYr3b6Zwh5kwCqbEVMmebGvuPuLKxeSFD+/KMQjq+HA8LkLLEi7T/j5vG0GZoV
8EZyYSDPmVMO/tZ7PoMchiwCiRE5GOQ8dByZSeLte8Jbg2Ois6lNn3lzzOMh7aL2
sKHnaHyyLPuTfhAYNrExHPFMFi+9c0LQ6fJQFYYFuEm+GVO68PI0AlRs6WBo8BYA
9VzS4B3VmRcPjH72bFOowJrhOzZjAQAIJgoVK7gexzTu4cQ8sFExOvW2i+J+1dc2
+j1QkrQR/9r4vWHRQPOABLRu0zlkfzG8wdNW5/NHGxVMDCC3Cn0VmXJUxtZtSMK4
Kg2Osx80m+T6xEOl2hQa6mnDNT3r6Gz82Q/P1qA3ye9ceL927KxJ4T0noxNmvSCE
bIn+H6S2rWEL7cGG3r0/dY0ljyW1L6F2qd6u0k7TU+stCW1j7Cgw+MfrPrCLzjjr
c93IyXHwuhhafiwS9LTnb7KLJ2jgJJpus0YAyn7E3CM3FMFRNj/Dof0onqOYYWl+
roIyFfxwKqC6JgVQd7sPgfvUxNSwRNhxHr25X5eCkCUe6fX5WBXFGWkeAs7OGi/i
rg65AAVcrnemAMbZweR0p6CVwLtPq+d1MwQBP6aRZvd45RjINsV8tYzkqwlvpRaD
By0yeZI8aGZ0wfivGNRbEwalHzbgBKNnCkirCoM+9CKPz6bUYjnKjyHwhOn2g/E9
C45kEyNBZopmrtwMuWJsn7nwHdSjDxGx43/F5JazeTof5Kqfuza9eR9kh/uZ5iz2
RjZg3B1TFDlEX/yCb7C1DqWHyP9WSnimzgVHX4AbRDwTUeNkwzrdOjJIosGEgnoe
ux2fdx5LnP7ROcTvVoCOInuz+dvsF0jmbXFUwth6zkXL6pXOCguXdRkTcYnlM84b
K7s9/zabrar3GZQns/r5Ywq6ECkkGesGkLpWLr5gFzcjetNHrVLRnVL0SY0A1tTp
5+X/9svXHPVfOetO6SouQBCbclgyTMN5ZfO9s8sUY+KrDmL9YwvPbHSMdzSflfe2
mdWo7jtpp35pvnHcsFx3I02x1hD6NuL/co2ads35hW1nU2c4fTwozTp4k9hebTnI
9vjqQ3XT0351u/qmpJEztlxPirHgyVBRsixO0zPdwWygHqQX9HHmqycFHi5Ft/dz
yqmbusTczg8NKasu5VfwJvJiuDQMqRER00rlK9/yQ/Nw6c2aBp2ebrNiuZ+RiVst
K2m9/tkPHEcb4ceQBhHSs39BmtIHUbR/zZwCL88JNOqa2XWNJJKJwsXQKZkT9lca
Yjqm4jVcQkTP1ifQJWwxVYt30SOtwN6f3y88qrkElDs219aiWVp986fRA6yF2k08
O5npaDfTn80Yo8J+AGLE//tgqoZnySL6KXW9P1b3dFbSpoFu6isVZkDwAoFRXUE/
`protect end_protected