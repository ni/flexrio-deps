`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
rSYIM4JmoURNDQ6iqvASxECMvoifzx+aFGlaKMLJ8f1ItXFa/9ZhwTWkdBxGFov6
srcZLrgr/a8FqSW1DwBGGkJSc1B7FbdqXaA/yQmlCxNDSF/KHwmC4M6szqDhyHnT
ip9WvnFG6+r3sx7yh4dbkmzqkYabfGWQj77BY0efq62cvtevQXNg1nMnSScQwzP7
Dq+DSI8mJAdaa2nx0nkJ9m+trlggxNBbawZhoo0hQ8Yt5/dMMl0dfuebsVc2A7jY
3JkL7NPal6uRHl172pfwPd5J9VCWIM9i5fjIyidhmOV4yje0+qL5cHKGkqabIJji
OSj5Tl+V843LKkigH7x2YmsU6wXvkzdAC2tUCyD1YDhlRciP+zSiK01RU37OLK2a
P9cEFvJ3Uns44UkglQ4HqBa5BVUXlUTS8kpC6Pp7QWL9xr2KtTnwhr73ifQgWdSF
tdBAN5yPuUt0ENIpTrqgeSphvhX+/j4utd/w63Uh7dRmQNLTm5fb4YajuexyE2Jm
iZOGcSKcAeUZWdDymNdbf+0+44ND5mukeRkUNBGh14RvSnVAFe3PNvBPI3HAnbLh
F4zjXsGSuPyRzWCQ/IT8AMZpOMPjf6SAxo5mUtsMa7bJgVJQxf3p9XtCxHXUpJWo
URUCucB6B9dnDWyvawrWAf0lOaYILTwpyyx+WOt9XMMsccNXUxd0sWm8nv6lPCBX
sQAI1QaSDa0Y2v/GEa833NM7qrOcYgJExQKM+lBkUmQzYdCHQcQGnNB0P+S0lQh6
KlQnf7ToDbmx7xs4KDphq489KP4waXNrbwcPj1rOfHSK33hRnl1P6i85wf0mHTq/
hZPCXdp6VvyZX+RMg9hztFnypKxFdYzh1mHQaCvSatxMMx29sXMh/H43bhuxPBNM
l0o/sB5Nl0V8UJV4f3hydoP41M3uSDfNFMs0Y3IvxUgVFbhHoQw1xolzeXI0c4RN
Xg6AZP8USrKRhTSpCyBIuVgqizUfhBd3KvuiwYdeqqeSftVP5HPfryMPwLhqQhO2
4ncYvH3O2K1cWmmENhDHo2Zpox+hC/5XvYw4YjSD+3Vc5k488ToP7eR53aEpLkyp
J6+QSeUBcSc9LFt751uSmafs6+9lk+AUzAS7Qr1jH2RwmzfPb5Ifnw4o7pszNHQA
DjEfjHGSVlffuIMj8tlORyUy0/FXOSibX3h8188ylsPnlavr6P/L8RnKzNRvpsM5
Zu849TikpTAZH0OjPNmGsiPk2FoESEaS4ywdq5bKgTYKf8qbEZknWiX71odpAHYf
ErYnsP5VYzx8QdCAjKgwnlu6L1hq+11K1YJ3p4EFne3uqiZleIJHX47mLPxWJdmU
SWxUieuhMtHM9PfGa9s/23XStuuvX9mSU0DQ+ABWU/59nKYeLUU0wtG4S16Gf5Ay
/kmqKtt3BvfzLbXpJ+P4NtauTImNXEMEeJR3rLJpqdkaS4yl7vxN0qSYwqopCSKA
Dy8rfhINmHnHy2r0tKE3pEcVJlqzEkIyahvZe4hBZazY2mPPKh9aa1x/CNwj0wXA
PHuhkg4h84Ek8NxvrzigesFM8nyu/M1LJbv/U4iQ7BxQV76VppKLSP9whOjIsa+f
xzH2EyZQse0XpAN0sCZriqrBaszbzVKcMG0ltM3BciZWiMH9kjO7EsFYxml+xYJ5
On4cC+AGAHK84JsjK6o05VgJ93SRLsRRD+WIFAIoQSu4skNLq0SDhV/V7zRFbTtu
SoNE+iXZ5WTzqZ/XJjR27sk/v1eIii6QaPBmkJ/eDFPUJzZowxCTE90MaEKvRnat
RHlKoYHuwWTQ4GK4Hn+yA2AvCE/OfWYgf+8LWBfYvkiMh8AAp645aNI0Kw+7lrub
FDI1NVKpQdfHk9ieHoSHib+nVC1Xbknfo5CLSd/ZmR3ro6frFifTKUiLQD5zWpgc
gIJHBgLkO/k64BNhO9QvCpCFe97XN3qcxC/weRfSYojN6oTWLeS8XVJUkAWlHVUe
pMlw3paQ4cjkBV1xEXukZ7MwIPyCOK2huviifbQC6GYDpDmQCPg9g03L49NOjdCb
z0Pm5R8i+nCrs6EYLLgEnvg7lQ4zUz3b1WEVNmhnDjSfBFAS83Jsw4cEBABxY0x8
yGB1POsikX8XenR/P3rkd83TnB4N6Lz/00bSKYaQbVD0kw/tbXhnOxgTPfzlC4cJ
8g8zKbVT23Vgzqm5wImI0Vdc/x7u7z6df9naWSKgmgTghZNBA0aTT6SEXiqwbwfA
mAI9c5qRRVFcM1lrUfOUTJu1PKqYJ1QVamkyaZCC9ZsJb0KcXSDZ7rhlJy3zeC5B
vzjKewUDakz3jy8vInrglhTsORsHS8rctprXx4xEPfQSnbC+lVeoPh39lVRm8bDc
27+vWtYhZMWzGo+90Wt31zrKhaICQCsBbSuY1792T/P9UOspUcvEx0N+OL1nKvQ+
XGcUpXygnetYjLBzPkGgeSEuhtQIFHaDX2V6n4X1T6VwLGQeidDJW4WoPD98jYqQ
CLA/jHq0Hy8gfD3YH4VypFreajIQojL6pVg+a1OiEfVU8xlol5HoybxtBJuDn2tl
g3b7UNKdAPxWJnmMnKOPwz78z1IHjQcyRNzpvKdRjgL0HeZkXAiiQdj9p9nux8+z
BI8NKhNpONBxEjv7dY/IAapZKMhQJa5i4u5/nJ+C/zRAuJuE7B0mR6zvIiWKXBAp
paNjEwOxEy8actaRv15NlhoS4Yp37bEjqO59FtvJf5QcW6k1za97oRfm1UPWaHZ8
e5IblqBX+pNXbtRHyswPLk0Y3HlhUllBsw5X/exPAxYMKwGBU1hWwPh2fF0+/Ic3
BLC2M7z0qTIGcQm8IqC+eDp4GWeoKxz+JpYMoR60F9JdIhd7TxbREccU2g9OGdyJ
D3vtfsjTR3rcUzJSu5jA9ZnS88fH8Jg7ozvCJ4ZFQl5zDGzwGahTAP4VjYvlhSti
ZcGNNb5M3MNvRcLsrcW4nxRPcCaqM1WEAgMc4x62h2fKDg7yL07uuvOYhsHcISIc
5zcB/GhMnZcz8mgfsl9kKGvz+3PIkILQPl90SlhCn75t9PD4gFc+38gncj19VoYN
AF4MI9O0K3Rtv9EXujydoTWLPJEaYtXh1UMLKoS90Ohoq4a0UcLZ192iSE/IVtYm
EdraG59jYvEWoiPdUgvNixTHvSzRVBEDBAq8hO9gsKChWzPQ8WEVJQxPDy6ydzn5
Teokucnqo/fpp8lSh/ZfnnkOU+a0h3z6glXqNZC5ljGkf+khQd6HMXzhqgkC0DWh
vsveEX6BfekKj206/PnHfvoyfAiY/QSk14UapKmOWPMTve/icv5Vb4GKmJx24cTk
KhaVXamFl76L3wdnWwp7L+XRHLk8XUApp9c41P3DoBLgxBoQofwVm8ZU+w7GeoqX
VCEgHYEKjH73y233nGz63HA/wLDLbStWOza8zxWfb3Ko3EwwiySImSc4ch3Ax51Q
dG2z4CZxPPKhihpNCQWgYnmj9W+jAgwv3+yTQaSp27UrDK5jo7BjkwNMXyzUFcSs
IQGXN0mWAFrLwDkBum9eEXQFGOwJbFBK+eVBszHdGTkCj86ML4ZqHLikdJobftq8
JXYACOUu8JB9rup1tcnYnBTDI/8biEM+Md9x1qJcZO1MU7JXWOUs5BvDX5s6FjAO
7Fck5PN/ncQw+2hoDdK/CoXf6IvucA13JtpkGZY4dj0dFrl2EmFVHJQ4rDa7InSS
Nuvp20eOA6yKrALemgQcrMFTDjNILoqLbAeyQILyz/5oVn8UMJvMZXRNkSc/JcHK
V7XZdY4Drbae88g03WMGrfDarxiq56w+FT/xanorlTG3mGiDH7+nueHfnxkfB68u
Xu1pTHnhIz+c2H/0XI6/+uNQe8FnWMnOED9Omn/l9JlFHpDuHv2ev45O8sezv868
FyPW/wQISXr6BdM90mnWRR6AHXZsOzedJKu80SmtmP5B96ErjPkeij44HiYoviRZ
ENsKMM62xktQQ3SjfTL0lm3vQa+7lHr6yOwBMEFNMxAmXOUX3RnB7fZSsr0Mhchn
LJl2EsmrMCiQqORm0+4Lw0ANhfbTC/6EB6lOsMPS/BW1mlH9LYvzQMZ0OZWrrNOz
zItl8+N/AHAsOUyoYN/gPuz32AQ9qKTzOU0G6+Puc4benTkcKAtSyAJ6pgIMlaCV
WpheLfYVbW8jHyMa/axdmu/ZJys7vLNHppXtfyEUO/V0KsHHcDXCJEmbZA1BqWVz
x66yKNchzbbn+Xcon+wsV8adErEA1SVn8oHE7fJTMM1jwzJJWy+xfnxj8BEXQpiE
NR5R0yAR/dwYRk+r/3jS6e8RzY0IIp+Ra9IiOP8W/EoUpXwJFsHpogWsV4cwpjq+
clvrhNoe1zJL+5YfPHMh1JKmjJ1FirgwRQkZ9kyFFq+enisOz3jWnRunZYSPV60C
UGZBlKbC+VeEvEIjg6mW5h9nloqAcuvPWMVNNwBEape9WRqo82Gwb+yCcuMcEq8C
5Un7wjhGhrmFhH00W3zcub5+g6XTN1lv1TXhDehLqqq/Hk6YFu268ghT6q9rq34U
Pp7vs9l1mFegUDTAypgiQyS7ZYB6wkAG+mD+k0xRXSg0vK0O6UZk37EVAbv3PgFZ
otiYsgDZGUDQZK2VHvq80ct9gMnWJF8nzYejLd7+QpqepBlAafhUwo2hkZInE0uJ
EJpMHfN/WqQ1TenyZb+7+h2lx4ezoLAcs7kfWP1tN70icJqhqbm0MeNkRkzrBwgp
rdD/A2ZoOXIzLVmzdE56dcdD3whV49VTapr9k2H2MqAEUhVsLCEJSfWLhc1xjd1f
odswbWrs7+/wI7X6Z/p2YrN9SWmse0Lx5BCSkydUGSHbnHh7jBzN+Ir5hc0TiNIr
mlUFxUkBlDhjYxzhYbwtVonLT4c95WHctmpW/AGBVu3Om7tHBiOO6rilZJge17v8
mFG5SjHLdpKqncV2O8DaPYaSo7Ago5v7lslIAdwMNkPBtHQOicII8Pm45yCQBz/N
sZuy55Yi3xfomMw9C64zcnNQ6SR2B2qE9T5cgI6mdCN/COlvUfmxk4SwkAwadPRZ
m0umM2JpoJQSE+D9lWKaDyEpGftU3rlVTTgEYno4LH5m9VQHhH4o1jMq+IAImLqW
jxUMybMYPy0JehMXTu1a4KzN6rgmEnqxulVhgINQRMTrrqwtO1xzM1zeMAF94fNp
vsXudMjekdzGVpFJ4iaR9E1Rn7lOc64FYsuQyshOjrcYehCE4Sz8SLvg7fVJc16c
igJGWMYfvoI8xJ7VjH9DkgSirodAmivr+KHvYM7PDqfovQF9t4fbA9KvaWCRwFzI
LLm9x/WPw3BLp0qAqLWIW92jOZjm1ZFs5p1PgTAUB2vmjFtWe2e+k//9aqzxJfxB
yCJeM/NXTSBqVN5NMS/TDbmr79oOjSuG0p6XR3DswS9X/XXff2ne4f9bP8X+58TH
fJHiKEH+9wT0pdl7ouHvs+WJn7wArpnE2KM6LRBwaHBORvwnqsO2d+nUsSbOQoWh
hd3QzcJOf+IShlW+6Mp3vSZlQWyekCN+8SWkIDVWIzt7oflCHcTmJXRSfVMxlxkP
7LIkTRjNclO1GOcCH/PKit0XUNwj2KnrfQmk5b0Xpc+0UKrLC0rJSpuHLQiVUZzc
i+lyYeromsLhbOY24JEURc2jzZYE65WQRjjUgrm9MvaUXJgw3s1nmCeiYVH+IlGS
7ox8OPUJ1gOmZsffo1EFkmfRMZv/tP1EZzThUxKpq+Wn50dOsMFGiabag28FAs9s
dMqFkARNTyjsxsgW6T6h4m/smGzX3u8ZtGrhxFhrqabqtev+ydbwNb+Im6ukr4ko
F1ewLKOOlG9OQ2HMl7XJEIvG+cZZEM9PL3hYeqcTiK9C08Wa/0EH2IVpA78UUKln
1BF2aSZ8pLkXwU+fhIxSkqdcrC9Qkq0Zk5TxvvPoxp6yKoJYJgacvCkQJDFd2I69
3BeiPRtB320+3rBIuW0iFjYFq+YN0GeDk9esF7v15MYOjaiC/25Ce7ajompsa5pY
IWi/xIAMusU/yAzjCmd7pWfix9tR0/DZeF26mWnAhbH44VyPjziWz4Kgl2UJlw9Y
87Qw5hqAaY7Rlq0oFpwbwHkHwrODPX+zRlDyrdVlcI+LWx8K3LnKCU4AdyL8pC/V
3f7XbfKZEyfF/Yhj+SXTFZ6RaZOEKL1v2VwvJN7JtRqolpBbaHrFUCHIIRHtg7j0
Spk0c2ydCX0FrucEtMDBk++0WsOcofv5+yfxHZw57XHIU77O+2/jOmn1cQdpi3oL
xf2okXgs6SjE659i9RuGMFfn4TsuJl0tz/iHM/DNoQZ2cd1fseeu6WzC/l5dXzbR
MzedOYcJLzKvqUNzgU5l0jpGhUqQwwq3i23ohW02prMyEEutLsN0K7903xwYJix5
KSe2QWKYFoZw7TwunY5NOtLuelDoU3G7YZ5Z+alelk64Wy2UHr02iY06GqZq7JvB
lyQtawuL23Y8V15HOAku0YNsAnAkrnTKtY4t+Q4D5rj+mzj+x9RyYBnud8XpUqVa
i10ZyMUArZTFyYUmj1GIhv0vGO8x5XCUkIyKffPAZEigfyJs+ZrkToqk2UpBbWGK
jnK+ogifFSFnQkdtq4MApjv1WjPcPmvcoQv5+8N+yu20/rwlr0eDI82qPKLvAZNe
aZZ9Td7/Brn9FnzyIki7hIMc4NItkuI7bXpPbIgdOsKgjqQkj3xDvkfxVbvh+4zk
+ed5R36MYNEzOfBbq9xuFlVHpjys5qwDOWTUG9zGIhYIbghQ0CyKnWinQEnPVJ7x
yJLw0r1CmxoEcdF5oPqtVRIndJ2Vw56Gse/ie7YNbZKPE4GUgA52Q483x6LBb83V
/D9voY7YYBNB7DvtIkRnDPRP0pJHIcHrdu+FmzNV0LOd2DT4lhs6t6unjjjJA8/x
GZICAjVxI93WDpytyxlqq/O2STBkDRqMxMwlHuEiCqq6hLdH8/x4BWe9qY9LTrjK
zKfqjIfWY3xcj1mRFuY0TwWbeD8cHdlbWQQw6xwKweMMGzNwLgVfxKMfM3EodV/b
9/xzQYXLMPBU1pESEYcSUTzWC2DkW2J94YSG2ZO5nFBjzfdqeWbXW19k6xBJibRd
NH9RpALOC5+EVUGa6fdBajqNkQ3XAppNwFDn5HTz5ia9w9kuwR7VGSNTsqPtdIqM
HPVHyk5IqwmogTb575swYEg3srviH0c28V1LIu7Gdq694JADUkT2KeHd3vdKQyYF
U43QoNqa4KnySid81M0sPINexkjoseNHyQB722FHBRuonKpws4AIYmWP51crg99j
4a4wVzGhJ+WYXJN87N1Qj2kKRV4u4h9W+tx0tBWJOWlJ5iql+v5P5sE/t47Ny46l
gheyjczLjuz0zfJ/5MbGat95JFVJwp2JR2sqBTof5j+cdb12PXypyaT27gUVWmR2
iQcYwSuKEijjBWhrTfQBNXCC+Kvhj79k3eDJQLo0wrdnsMpOmp9GxuhJLEJjtd/0
XT11segphyGVtMlF+59JprkLjEQFQfMHQPQoWHAq5EfxPKcmM+er4vk/HfRZ6Y5J
IG0v0qU69l5WTnd/BlT44a8ITzDTlK1rjIFxclZtib7f4QNQ3GF0ASCSFAhkLS2F
HiLMy5i7DQ2g1DMI8AGcDe3aAJppydWc8ytFVBWMM1T4BCsiApJ679nIhJKgEBfy
nQh8nSAq7AcXO8dQ3BWk5JxoUjXgp4i5t75DFexr6ztB7UsEmRrXDlCauOrDAAAf
2b9jhzIA1pRl4eaVHJbbZlEbUlDdEjo3ls4V4FyehWCdRSpGKZXlkYOoB7Te/OFI
KHT9QwdFrHu+B/+DzNJy/lnV9X4pKtASmBOwmaPPXWHbAa87vQzPCIvL/rNm2Epa
X81k3ryVCKl3oMPbqdnaekglLkqdnxedWId6nNDj+01lmmt+Nl0Pogaphr9Lc0ic
1SmsG35VTt57KHedR+IbMUas6yBSoi4mhsdB6BW8Bd1Yo7Ofksa6Q5BWOgz2B136
PmaOhV7EUIbylByZX6ooE2fZJ6CW/Ns4xYvkGMeCUirJ7auOeUkf5JwfDiZK1Dlm
mmUTzcqJOW9AJW/xrVygZ0gpyygIvGwpauaZmL4nL67s40lRNyK08Asv+Uu+q8v9
g32ulutKlthh9IypNYDcetkquEZ4BBhp6nyxj+P40jzBXae2bASX70OJ8Td9jd/l
TLX6wJ7yKfSlQ/RbWhp72Z5ItnGj1+xf83fJVPvqEgxiA60Jk3nb2OL9yAJl5IWs
aWbU8NFbRs/CKXPDuoPfKSG15RLZ5G+3RnO+A5Ach+Rgpi0Mt/A+UaWPl4ce2t7K
iieL4PVd5e5QJ/faGe1BNk9tK9NQu9+Q+JG38I5B+GTtcRjJrfuf5DojoGNcGKf6
wDyEwdVe/lWMZjvJMTgoUtb5AypDLMcFw2uK9v+WiUtalgASM9lTVWnyRO/+JQ2L
wh/i95VbXQ56/bqvpZv8e1RoZxD+7P1J32s7+a3zW6Sv1bRhBqkPVqzazGaWsPX5
Dc2hU5jXF1oEAHQjCd1tiIRuHSNbcseK0/rtBZU/xTBXXVC47tMwNMVSs0zHP8Gz
2l5fKWs3R9VENpFrxdxq68zwJKNUU1yGD6mwl/yP1DUd5MrFWlOheL/mQBR3JzdT
rBc+6T5or2q2x3Rg8ROVAMqPVCA82eEUvHHlQuiA/EZD7TIgJ43VZc02MfI+x4st
37EP9TS0bRIM6a92vYOSdgNy2HxfoKZ3KO6gq7lJN+cJ2wM0r5SoxAVgtq3FBJqE
c9DrK5dpeHBnQ3jisgiFIHOLpmbQtoRNM3TWdDUcL5joxEVmmpCr1GHPlQNEDHY0
/gLyL5uZu6xbNCAfRww7Zgfp40GIODt8OupAUwHtF3IjGKsH9rToKawrjxjzYC6c
l5gp7UaRjD9xtVfWdtdkzIOe1l5D0zpAHVfcJKcpBl4Z+G5gcCRR0cxxRW19UMiP
eyvIALPSo60JoL6gNV1YlBuBhPoIvG8SnoRz0X23kTqb9dD6k33HgRMi10Un90P8
0HwzzFpKVE2/WoMc5Yr4f1vEsbEo6lomPr7VD7DCNqq9klPO1LP2/+b8cpmrn4RG
ZMed/bbzHNgobusxLSTfG3C1VHRKVDHKDusq/zw+IGL+2P3AFX46DqOBpx2lsw4M
a7No9+dtlRK1YrmowqjYJQYsQ3qxW8QGUOsDlhvnCe3+6p/eZQ3RsYM+5zptDLMZ
HDVSPR1/ZZb2OskCmAXRtPVd+v/B+YrIKSlIYfSHF4c3aTvvWy8N5Hsvb6uU8zu2
VAgkCF9VnqjVx8yMsh83uEcLHSMx+Pw3ksaOaEXy3SJyCXss/EDlExG+qFWcJqtk
/HMmXdpU+FbnAcJ4eA6MFu6vEVYj7nEQZbUlF2u4mSWHCD6PtYGngIoSgOxkz2Dw
HYcwBZ99kznyNC7gBVnCiujvPrkeHwoG7lxfunMNNjPCYsQh9ezKbcvBEelxRrgR
5sZCeatHQ+ALSwwxXFL19go08diA/F2FdI1KejQm5vLhJ5ksr1lc8LAkDHiD+7BC
+sArTgqLnpzQiF9Iggfjq4gl3VduBupjpcesbx5QtSDLQiXLg4NGg0ngZUDAdnVb
QgnIugyjaXUq6Qov2pvm/VVCOsfDt5pxP9ql4doeSHhzX/JHMctOoYZbBN4f3u7N
CpyuKUQF37zKJTjg/USQdlLT899RK44bnXN0vT/sSs3gDY6YiYsM8F/T9EgRmoRh
m15mPbZh8U9gItFfpGCUoOB/rLdbVfPvoIocky1Zyok3BbpzeL9iW5z2gX8Dm4km
llKRPnAgNDUmRqOUcMMIECfjZOVOeqGEOIP3mUe3F+Zd82PQJm/T/y29b4AZRHRN
o924rpACcOvJVRivW7iPVKcX1yyMdRDIEm38LTyOD6taNYp5lEhaeoxKDJbpW66b
jrVkJJVqZshg0+bI2A1YjcuZQJoHF/lvRiO9i6UyuWuFqztxh4Nlu0xykQZpB3mo
9DrJ6Unha7Q21wclV+hEy5jI0Q0QIIR8FFAkunLMo3hOHfJTxth+5dw2n2HxsGa8
BNRPKYDieuoWYBr90Ei5ANwtBryAQug5OL2CJ9d1b912tu9PuWWWtrW2xRf3EtJu
d36tfjgCRlAwJTqJBn8a6IPbelUppC6H671u28KiWnUkNEanxge5wqDRk6D5J3/q
+/9jHRvFGKuq6e1khzFzVfjehLb3rGPDCi17Wvc9TGrO3K0H+Tp5mnc9HXepkSkM
hpTKna4RUkzo51yCzypgD6yG6VSkHUGyl8Aa/jAukZvc8VvLCmoUtnjEEDBAzVFX
1waoXhUVgVOTjRxZaFas1MuSlociJdQZmMxKNiDQHy6K1/EuBl5RwCFLdU0/TXTU
sQ3ePOxBmJalluJQPoSDou9AFXjtRSuyyNkjXIxMNIy+THln5jRPKECVU115+nHJ
M4FvEaDBoMnenleuKCadIHhma8ycqCMArXq8g6tKgtBVqVSgZpgPsPsY/27NCKrg
n8u7K5gvEqUsjHXpJcVsARVWnB+imQ6/o0zWPCSN/8xVC4Fl3a7Tl3Dtw9Pt4Gm0
lJzwhtc9xfbCn0dyKYxh0BV9baelfNZTwjgT6GyKs11BwJWJThpgxYPsZAmbb8yx
ThWNXSsr1dJMExthHCZOyNy46MdfcYq2qdfqmIebE6rmvMaBxq7nZqhn6uz315oN
Byzr1hDD4pgmPWS7uqRI/6fYT/BNBhJB8pD/Npb6T0CBwVU+LjbcnVhsTPeEt7Hx
7qTIp7aTwHQ0UwdL4yEUAZ0X3gGAOntUoEOhzf7uXW6a7KQiH+eOGi15WjtZGPJg
0dAA8xUVkc8tOEzgv5gVgzD5GUJoxWFW7gGMKcVa8nRsp6q1Z8rQY6ReEEov/zGC
oiFhNKlB5FSi8I9Zs4kiWjSZfW9jioCRpzVh+w90P4Ddd8c7L+pRtzJIGjEgffmA
7dUUsWtI3hPlDdwXTQh3eCe0+EzVAMTZpmDdC8BR8AiFUQ3kNsYJj/+bKYdDYEgh
j8sByXqxrR9IS2VMxQyPeD9wBCVjTTaiKudkCSeimtt/IKYkhGOLhuBMTqHOlH4s
tFB/7caMBLgUN+A6z3KXRakOHvSk2AsPQPEL8pDd+W7T1Rs0wikVXIYsVYd6zFzj
AGNQ17z/pu8E9Xx1gXJ8536t4vZJtvY/voR2zRr2DvWFU7Xy7u8+sf/IqWbgeQWP
QEs06TO9SpSzRrHUa1rxYYya4ncfGfNN3U89QnBu5LFnNaVbvpavJCE7KjUcfbcZ
V3jnkMlezolFOy6nBRIPt8Kslb5p3nphq0C7pm0EgSUfxUBJh7v/9c84nqGUoDMp
X+MBKiMPv4ieJVt0L25fG2Yxsjudogk+5DERNHx7aVUMWz3+0sGKYobZeb8j+92s
UeJ9Sl8JKkn20R2QKCMRHc+1X6m4tm1FPIcpitok9h8vKu+XGeB9hgIs/kv5laSr
7m1Cjjxd9ksDkvefB05GLqFLPYr2F+chhtWQ58i5pH/CH6NZObitJdDDm8qMUwfL
sCvpbrHaXXqg7Ik88JOpAny+WIEL1qXjFy39s4nHlh2y8lWc1eU+wTQKhTcF9+WV
Ps6mmDAK3q4XjuvXv05/m1SbiLXj6LFDCTtyntm6pVXD6T2l3ZLeOt3JALfL+bn3
f1duQ4QrC+sWjTe0egIn1OMEWnM1zpixM09ItcTgL6YjiUt06qkDCaZ8stuy1vbQ
ZT5OASxzrowl2DrqhvlXnnNGT3GDExaxygaeqPhlwuewlG+436Z2IvoMEbIolcyL
Dkvxq33VmC4XVIYw8gJ8DNGakkVB1n19iC3pVTRDovU0fNK0uMCf8QKugHyQ+3BL
zSmnkXkwiOi2XW0pWzn9EV6IAjEvrCquVO/ZKrgpb0KbmpB9AfOc6Dycz3NGgszj
Zv8jWLx5p55TrXb+Oyq2X0RcEJbboISKUrRwRGC2YfbSVBis3Htt6h/Pi2HdFZtV
6DqAe9lGwvy54D1JmSZrwLJALSOawK1eL0p+V8qUOJXuD8H7WEpD3B5J+gISfkm/
NoxgnWG7Xk1Y/EcItBDwNL0BK4PTFyLP3v8OiIDlvW/KnGa9iiwNfc5WBK09vlYW
MRfcnB7iCYMQIhf1SolRHosEYTmXujrSFulLK2TGfalQ84cMnz20naTOqa5r/8oB
jpXTAuf0+IJ+FiMs2xdnM2LxDyUdAkEbJ28MfTZnlXZozuXevM4R6wSHwbfH2LSB
AJ5eQYisgYG3yWOvHK5/51CWnY5VMxRoRY8yaUTY74xm0gR04hThxn+lBM03DmdL
ZMUAWtoQf1XX1dYbiqzdjtdbL24knrYX1MNBOXitqg901d9Wrn5DmneXUFbekBCZ
v+zrB9WDarmfZHC+w8ioHhmSVE1+MvOTKb/inmHu+04UPw6R7UYvxew94D43ijpx
7wvjrA4oKk4ABYWMcptANN0jcWRPiAIbRxghdgl9epYIY2rtnylcZEyKkaG2Wq0w
Odanfq0wn5Hhq3YCbiv9UPQ6Ep/v/AAO4sjf7+9yfC/u4gB6WpqU0XB17qxrizSk
yO6kycixz5imaZFU9ORAc38XAR+tq6Al8B8DQN5dhQvpSUYkS4LGUMqU5xkx2JPz
/rJnKEmzf6mXlrN3RQ113fRrL4mCFTq/NOM+SXtyHPCB0YcdE0sUTPox7Nfo0pgo
Ge7N74+KO3fEvJg2/u9em6hxjcearpFouMJn444CIopgGzkKaMbVRjjCOkj9k02P
zso3PNpVkhoJv2BwOji9xSN7gG0w+r845x6Anqi/8iSC6w0MD0k2lCndUxoj9aLM
NEJtXTJXFtrLDNCixHE79SRW74iDH7Jv63jBcIGYURZZ0y+RGzG+cHVI6M3tseB1
/X/W9ZVyOffsrIQqNhd2i8/4T5AKTk4MIbZGVh5OeZo+UMKrwQDK//BThj3xzfKO
P7FmslrtDDT4yaCqW8WWtVMgNM5GsgsOswYlfesExasBb6ppYLODddPFlMOLnTzO
6aMLMoI3hk/Q0SrEPBJL0rDxS+prmmXyq3obPxs1rTYtpKeDCFXioiYg+REwWmTv
pJk02rj0oPQJsFazFC8wBbT22xxiboAerQjCGey9fyIJHjNPwKy1P9EFrjXfCAvG
tPHFq4Nri/Hlbwljx5hOqqRcOVjGLE2YIdOZzq6Di/3zxkeYZW/BAI7Dz37V/BFE
GjHNXjoY5/HniNyrEvCKx67Tq05+hj4dZ01M0EkyO866w5ZZK6wv+4P/DhgV3BPU
8fOUFrTTyYv2QnhrmUtQwrxmEvvnR4dpyPeaakIPUdOkTYIKJJ/n9jsNKQbiw73O
WBP6O9ebVcXwL1/9JiNfaj11ksIXQktQz0idqikau9AjoUQobP2qyh1KFzg5wLhx
8x22PMgxUcJuNLbd2WF0KQUlJCqKmlTKsdROZ3Av5XMThd3Rn7ewqdtRR8uvO5dI
qzZDRBL9Wk2YcSZ7wQdpVBo3CiXt51v5MN1ulmxRi+SDwqQpr+BvId0sYL6/qQ0o
gJ8eN8A6aMH18eQm6W1PuP/g9F+ymywvklQLrJKX2LijkKU6js7BaG7Cd2hQVwjm
srkBQYDh3yOXb9SwQcAIwC4dGxiHSx+0yCO0TkcEtRin1qyIgpLrjuxkfslUjrgy
2l6HwwldXEGiJJkosmBq1B0TK6FBbBbQBvxOMh8lkmF3AiyNwpU6ylsDKCL+s0bC
MGo4lLfBR0w7Eh6QJBx/gPq57BUzRkxfsrFQKPYlBq2IEdSYHYQkLhN6PjDtHHGT
1smHoa45lc34Rp99jiA0V6PJijSKGpgl+j51gcHlT3/rB9Waox8yWgueo3gAMhwm
u+n0Q19CuWBTwUJlFtep3zcD/dNvtL1Fm2OHd+tMw4qtWeukSezgYXpEaiv1eKsC
8LeuA7dadHZCIC7aluOPWX+wPjCjaun67JMAs3vgHx0Q/wbs2a/fmnGiaibH0m+K
+ulkqcyU+rbHaX7vBrWx4f19kdjWuXni+FWq4xmO5N/qcoAZXnADdOWmicoI/sus
tyYHlWJx7COqTmTpxUh9yr1AT4iwqCiV+N7EAm/s7Up5I9A9HjJCb0xKGwMV67i3
CSWv0rKfqV7FFQXj1axuLj5KA1GNsI2uOKzNiotGoXWcp7eqTVe/GFFt0Y+dywDS
S07tozxM5uXik/mmb1YLMKaHqdSovIPe8lsDgeGdmPmcTZ3rttX7WFh6A+DICXaI
vG/VjQatAE/nI5NGo0vaJhAUbpGu7nxUoI1NffI6zV55ONsc47VmsRSNc3lax+0k
Gax+G0ipSZzy61QXtWbmqFRGgM/xc/21fVdyXM64ybA9UUIkypBezEEXG2K0Wlzc
QdFGocAQE72JLxdbZPKPzmCYPC43HH6gqIF3gNLGwpunBYWifg5a4AzAz/R3AbXn
Qi1HeSJoHqDjK9qUKuaCmFINyg2eH64ts496vy5aFEfa83lrvYIr2gBrWudHSVq8
OuR0TG7lNumWv5vCxdHZ8SnF/ZG6Rrhlraujfr+vVwiL9VsoNVDDaEPg6TXxfI27
357r8LtqzSwR13Yq3dAhVpeOus+tQ+3gaSCXHFwMnSXfObjr+GajmQJvwtvEyxKl
BFqWO4iWRVPWiR+JYuxgIqiQlZBOdkCLA4kSaQ4vJykSBwZqFnZ2swp0wCTjV6CJ
81U8tEVjT+8s2rPFCtsMkZZRDFC5XCW4yDELzaQSMCk2Fm4cO7MljgTK0+ns56C5
+AVugy5Wrctphr9pyV7gSblP3/xPHMIz9iEbqHHzb3g2M7p/O7S6Hm0jbs8tTg0r
eXldKJRDlE0AThNTd7wsD5/ZYaRvvFAg8TaCp6zMProajuKO32XXiEOEVzl2GxMf
ydwF4KI4xW/c5LHBoIQdbeIDXKpimY12K8YOiJiXA3uRmt4ygdQZIIHE9fJODJ50
9LTvUb0wXJdvOyr2WhZxwvOd6DavvzE/iEyc7Zs158PUr4hE1Dq3ZTKQ5p1KCDql
hRxdfBYJhUbXk070u4WRq9X6oJyJqUHmYWpEBIgTCr1qorzPxnM7dljGbUZg89il
/+DfBDMCjkVPzAfENAV6gZPnpmyZP3cLpFgsfTjrBtth0NQr3GrfpNX72fC0St9d
tAWpyMScAXh60KZ4nsO4vz1lISUW+L/0iewv6YwYUY7aP34Bmv8tw0MqX3o4ODn5
GL8LapgGZo6MUGJsHQoLlPQNjQFp/e7vvZzbGQthywHRw+Vn1zy1ENiw2g2XfKcg
tdiLPonGlsr3iFnV6/sQfVewxjZtgiB/20Ac8bGZWfEI8cyW/Gt4ds2p+DanPwEP
LfyhbwoF2+724i04cPp7Q+kMHYu8SYc8HOSiHdZ7XfmhaNm07Zg9J3obIJ2xDi/9
wil+Epy2Rwspfe1u8QaTunelb7SfBF7u3dTFW51vqweT2/+Ko60isD8G740WyVAt
o4HptMd1Y2lmBwQlDOA++yzfsnZTemiKwETbEbYNJvG0eNxS55FAEhJY0hJHLWN4
RxPHnGf57GlYRljtwY/Y2e/vz7eZrJRaDeaot4xKFt4uZ+y+6xConkgaenGzianq
Q5JfeQjEODdXnCuzcXO1KXyjCn/6NHqcZbxh5Yfs5pLq0Pqq9b1k8eBfHgamvJ2d
GCY9k588YGmHjfP7S5iXcZunbbegdezTsSMPcu+XhgKzFEsIMuuTVVugF5ieNGTc
hCm4BdHaHt3n2JwDFWQvB3wZsi0J3xZkFvd6v7scLWBClrlQf/QSJhb36jmDCu5b
5aaJBXFdqE9kR1z0BP4Wolu/2KAIobCPN/BZiiOGt84GqNFQQuRAxA1mSD8B7roG
debxg3KGQ2+Yj3z8iH8/gEKZxe3M+8LUoGr+ALRjcVY6yaimHu1SfCnVShJANmUe
eW29aMnGGkhm5JqW/B/L5MRa28pEarIcobqOiZE+2zqvmREEn+jeM/rq0JMdDP10
dwVrsKtbx1Dypdh6Tmq+Qok/4vJ6nPnQ3V2u3x9TgPUZVvZVPgy4dOzVhk3cfSur
HNq4iWsSafP/uJv6bPhvTZqEbl8f3asYa7AohJWv59dXcEI+lyrephYmkWtg16f6
Y1a4hgmXMZB6gGJmq0FL3xRW+bD8Ic+GvU3Qa9OYR7E1lPlSNBMML8UdsufpevFc
wlT9RlST1nDJoH+3PWKX3NzXF6s8Mq5/bU34x4r+z+zAueXbGc7qTdmV5DWuNBTm
+siE+J6G265XnqldsGXp2izK4R+dcf5rw81DoU8JWhdNTN46osVgBoRAw5VSbGJv
WcHlD2IV+zZ7XAIpmznJ/SAoryNu2qZYO1R6dwYSIOgy/1mha2JXlvr9XpOHUZid
Ss5kVHgK34QGBVkq8h11BsvBAXtyk6YZuanO8yhi85x4UbKk97q+0s/6aKvbw8MP
lNmWF/UQGBv8yTcYBDqvCsW8ZOwjcBQ8lbwG2l5AIKp+0FlyMxkvHxjxvUznsDaV
0LCCTNP0maz5GyMe7l/0GVaXrbxJQr81FZWd94gC9f1L6kL8ePQxomo79eoFmgaw
O5wj1iqR1hR+h5lKFNqGmHCjluqCJXEnYXePSIr8O6gY4s+FHecncJ+p54Ls2kjN
EtKz4NZ8LKq0ygpE91tSg3mtS8IzYLS7BJ5w2/ZBaABdM6c+kxC26PK6y/pGkTWa
fZmQtCVIq+U2yrvzkWvo04+eh7sWgavRS8DPZsurUAoB5uhsLPpWnxIGyoAlEDoK
Vt8KIOyKgsVj5giQN7fiL2QIT8sTiNRhL7GAmSZ2v4Fvox1BVexvx6zHMhktC4TW
/R2+OKdMrYMHtgIJsINUJzUsb3PIlsyW4XT03DDHxQhtzsIe9m4/edEksGTNb2LX
eT9GP27skxMlAntlUk4buR49HC7ox0f+hT1qVC+OoSVxi4Tb7H9bhzya1wy3Hd5G
CUHBy1UsIG08fgOWRUCypVKXmfhAkrRYnqtafaqsz1Ju8vCAzS2rV+eARdM4C+4j
7cavWzkfB1ZH9dBisQyNwgnvxyEI5GXLjxRS0zOOmmgyz6oCmvBFMJfoSJo61Xov
4F4yjIB6H7GEvhkKzGzzgvhHEejksFjVdFhgOPG5iDviHNF1OVkQmV4ybaxl60wz
KfihsgvRSu4ww8fmjQNQFSLP2P0pZamP8UGTqmuLNKC6viT7gUItEHSfFV9Ft8wM
lHVESHSMzXgdTY33Eh+K5M0pK4hvP1eL7S+j7O/rp8bkhwiiiQkubEDPsSpWf4+k
BBlFbPVa5j8hfD/SRo1YKOyxY2o6S0RPqS2kL5p2qt/UNA6vTUofB3Aun1o8TNct
hf3r85odDBAvP/Ki2EflXPwsn6agyygbvR9OxAUwG6kNa2nwanu/bKApsaaxNEu7
1wKL8Jk6lZsxfJZm1WtWk+lw2NIj6+INctD08LkfrjOdnFtWz13WqMAvAU+3+fyv
lM9QXcalmkR9p0HqizWT5R6AhwZdUjNGoZkv0CTAdq7srQTEJwCJ1DpwcGyEHxlz
AcUmDkLL91cYXffxLxNVQysu97lhIJVSB+i8K21qU2qomExF0UILGoqnjC9APWaT
Kfm5ngYtwTaHDLrSSdx1qDyZolD259+JfG9mNWFvwGmoH/u4mF5Ie+7Y2tFPsDz0
4d5KSBCtNPj86yujRSxSrIg8QNAdyicGuF3JRxB9jk2Z3t/SaZv663qK96C+2BLh
EoJRdK/Tb5BYNwitUTIvkP0P5yUbX/89YRIDhSY+GMm4VtkYq2HeJRC9lN+hcAf8
15G8vd1BJ21tCOjcjLChj57rPhCb1IyWLz9W4yXRox0mBDQ71c+k9gJEuV+3wwfn
qnnYlwNB86ruobdQfcN9sd6xkotyn1AKPL4AGjZrzlo6335G8gpV+Wp8+rSg3sDQ
TOYMgAJVcgox7bNok7/xAyJaMRfGgYHKalFWc7EJfwYmoTyUp4HO9ufP/neZhcBD
Agwf16vtskRrVbWlABLjKBrXYJa0onTYyqt6wnbdamdLP8EvYOBRENKEiK2DjYQK
yEPT0bZcHT88wLJxA7JzDsqA0GmlalXtb9zRidM0Jx9N/btUda1zzIXsKaw7wA1J
bIQxlrrsm6Iiw422PZ+Ag9mraegk2hdIric8SNtHmCtrBJpkPrp0uMKr5h2Cksya
TVXGeLyTaYETplql1jMRfLKTzNHUCJ5aVeI36IWAc0U3icIqDdf4+GtpOL2xpZ/0
cQUIzKonsQJuooqqdon3+shQrIsC7PA4a+2e96CYqejX/P/6YANTvBiSTRSJiHXZ
yyuFxKtyIQQa/Seu9Ir0jpO6grhyoOEvYZgYqM9B6MecjnzACmNcu6E/5yKKK7t/
vpouEKJTfStGup24ulOKco8IQa3rZrr+nMWHekadTi9qOKbgjxHxG39e5Qr9/BG5
Qrpp7Mirt7hgOcutOkf31vLv6PC2O5OnDjqqW5CmXjYD3ouI43fUk0jgguaKhVKJ
PWu8RHqkhFuumPkAtVYoA7gnP/qL+22RDF6ZzAF8cnidjrv+AWJLJ9QC9573kXc2
yvjt0e2pA/VYKB/aRjrx9LBL/VYKje7nPhopaRXKhq2lI52Yh45ZktB77B+A0Yuo
Ipd67MTUtiUucZekuC/B5v2bON454iV8SbOIXgNMTJbtbFljCGgL5pJpc39eD1hg
jPjAZoeCV2jkIEmzUMk23VrqpxsLRRPy6u4OIn8hC3QaU+gq+aegsY6qsw4plhT4
IO4J39f6ZunynC9iRKOU9+S2APWagLzE8ZqGH2ncQNln3axJDCGondky5zdvrAyw
62qVGNdwUMMPZ+/78AdwHkG/EioIV3KT5plj0z+hm/0vHEzFTlxcqB8IVvNCBHNL
AkWBskOfDbrncK2Hh23k3GZYWpwW+X4PafoQOTqoIbCoKGFd24XuP2eQrCDFqLv7
/tEU7XJHWa+u51NyWL4DsE8vRLrqhf73QpA1C4tnceuzKBaq3OgJaLz2XC5ibwV7
JpgR+52GA64YRGFrV4pM+2Uua9ilai4eOVHQSFekl0PzmZaFe0ocD4VsnvaxhcXV
OYg5Cgro/iBkqjSB6T9uomqdEunVNYWW3/bW/XWS0cPSkclxfRl6cNHaSl45b1YR
9On+UoR8u2B/hqiP7XphAAJqs9Z1TyCQxo4aN6xqK8p6zMYt6EttpDmT9vhzfd8h
tEaUE/aSs0kSK6e1LenFxE7KSC4HTWH+C33JA2qlzFP6WINZMNxicnpbXcrsHA5y
BMkXCA7TqiiSMm1xDbBF4UpmgLD1iQEHJg9Nf5Ycw3G4d2Jdl3kXQY5S47dwaUTZ
HoACWyYJorYf++/hY4ytKiEYtoe7uASA3mLs0GjtXJuIi9M4IcUP47JIu9F03KMP
rRZ8s7D2oT8E+9SMcpiv/6c3xKhwifwHBDtj66HTXLzRNlXyiFrpX7/0+qETDiVY
Fp+YZ3DbU+rz6G3H8omRh5/2BiqjZ3W3HzG7cb2USiuuumySSNqCFn3jvDql3aOF
gcUOg0UzNvu+MaTwcqLOyEbr01hiXUHGiCgyVfmKJtLalutp9APZrxOBqIdax4dN
09foD5t0kHVrRqcF5YgAp97++8IuHgGsqf0MQ8P2lGJl0HuR6NpReQTtPhILmRUk
F7XnM0vwroJwCQdxy9m9RNUGt2WSjlGNPyo1Z33ZZ+6RAzh0zDdNlCjmq/MQv2vf
y9uSr6YvqBBtN03qj+7eZsV7ELMOfjv2zUpP3PTgXUl8kOrPOzFUYR6tZmSgT9De
spfrn8E+iJEzlRBJR2FFYnT5SJDBEv45YLvq1BO9INaHvZbg/n4xLKx+6CJCoIgc
qe3HMujPZE3iRijVnjBaT6uc7nIHH6k6mEixHxqF7ae7Yh6YYQPHLmPcZ6ZlJnG9
1xbHvyCSAeXXKtTyTqMrV0Zd4+a+aS3I9lifC6DGwUggG18Pdz6wj2G8t5sGAf/i
E3maYXR9GtSSVEfe2GBK8X+QlKxWMgfVc8JOt0deU+pLNyELPYarRZvAyC9wwVfr
9LpS1bR8+BqsTprM/PHvyg4tXsA+ivkscjHJ59AMYYF7mBRBg9aSIhrdF8EIBqqW
TL9gPKYbV5NmnFh44CMfPt+bfUXknK2gnOhlwiQtDJOrAF89tcXt9RAwuyNRt0/N
SKFjZoNz4SxUvHMujBJIhVBB2GSF1EpkSsnTEFQO/CTenaQ5vTsmF8X60RIccPWw
5qtml75ZANJNIv8JCNMnU92SkF9SQ9aIK3Zid2rqpcVNZmiw9gYZzZy9xvtURl4u
6x3DtYrI1BM4QhEAHrvcjq+3UKWfHh8bJxiS18uhVviHDV+tvpL+qLmRBOaRtCCx
x/jlkOn/yXLOPPasMyf1Bhs+8g1W882elWGUzUPDyieXkre09u/hFukTSlsbp3aR
VOaw/SlpJX1jmlZnXanH87B8w+LjHuGVxXQ+BRx6pxG6TSzp5cEMgt/s5U8BIsxU
A17U630T9lk8ewHi+y/zIh7ooV20tNdgTupJlZjDvw4mOVHwXkwRRYmdtbiYyM+g
8G6Lm3m/CfHvB/3lRZkijdnlwrP++YGmkv6N4GWORtuy1mp7HkP/FWqTbD9/dalP
bKoQ+36AZ1TwIR0fCMgc67jhp992J3A2NY2QNdiJ5KNZQRriE5a4cK8tWX7TRrWW
pjsCtHtKLP7xAAx7ILDl7QiXdct4i0rVvdPwjV8SudMMISjpKVl/RTPaSm/QHwZC
AvPTqXV5+2831YWbMkEspO5vZD1n6t1cnaGdF1Xb8AQkfEnMBV0uDd1UCbqSvzkv
3QWtgrZi6eS4iIMsTFlW0T3afIVKbTONsrET/oznn34ZE6w1cWcyqmh5jMHUFMVt
hBdeweOn+IltY98IHTm5iFRHU7fFvWjRM14nU/ZrlaLEAPQWfzky2oYPzVN1UMcm
8OSoMZRvWt7Z++vFVUQyxxsaCajsUSBSNfLS4R/7YtV1nu4vP318gB+vZI9gcgk0
R5PubkTxgbB9dC+sqG69iFo5GYMExA/HZaRNTArnxMEeuAazTP0bdVUQthFWgpXx
vQsBll7adL+HZOnDnZUOib5XngZPL1d3xWQKLIl4V+1t4MXUtJQc1y9wsGVc5LtN
9HZw6oGNEzcFOhWaYaThHz92NlG/VO4n+CD7QDYKDSiwMX9+cBykyaYpaK3s+rgM
Opoh4PY1sAnWofO05A3KH+LhhIPMzvH4LVkZL9UTIlSBMtKswBccEsY+GfHza6h0
RHr2N9cPCmH/gUB2gNu0ZSdA0C3nhY8CJX8IhpY4QxEAJl6me1tb7/MxMNjhYjta
jjv3HN2kJU6B1CDY+LYg92zIoH+TV3PXBoWfaVWKm69wH0BiVxeGOQnIu9ZH80UU
BvjwMUU6nZQ9C/mhw6mg3HudCfo5dinXoxzgAGTMIA34OwTLmAdCVsbwSpIIJbzf
wV1uyJ2TZsVaUrYmIqYJ178t+gohvF/gnkea/Czr3GKEriEeazNX1s8zqekfW9rW
Dr8htSliMU03hDaaT3WVpdzIe+rsHpjpnbO5nr+RYR44bkKAQlLjbDiHHlk4oRKR
ti1vWlhj63ORBBuetruluKTkm9UXfltxOHTvNQi2il+vWcGYeufjf7K77bAOnzVK
6Po7lzCEY12JOalmEF4LRMFN1VcP3x6vj/uNxheau0YyTEtLc4SWeQ4R+HI+JLn9
/FsmQu/mkqmuSy1+CXUw0Q+yBTJi18GnBy8JNDZf4+yqfdZqxF+yvYiLDM11raU/
k2EMDXK5hVhFWmso3AASEgFcHGXVShqMIjPANLVhRuk28MINTLYrlB/+gNXs3XtQ
GivXREAmomPvePz7kuMONW38cfbW50f0iGtm3UKg3iAVcFVEF6Avk9167qccxJRl
WT69sYl/2fx/lL+2CuXHsj0lUBRw3E0FK5z+Gh28u3jjimR+KMpZQO4/Wrx+SJhG
2kQQ+VgDxznUZPHdxuH2Sl6pnnKZ46qwLIUDXLBcM9g1jiilnv35ARTvDBtOQrFN
2Bvo7TCjRH96bePOW8rH1GYEmw8P6s2y+jijLWBC6K+wX9zXLQJhfnplsfOjPVi/
4jGg2zO+ptywD2rstrOwv4bAlgPX33fn1kOejYufSuY7n4UM/shFt/LEFQ15YL27
V7l+vDmPzoid0ibE/9S86MWBW+RFGagzIV2rf++diWUu55BflZn3PcUcRzY9Bnx1
47uwJRuJeWtl7IgEA+VUTAih+i7HwEDkuueEZoyMiw5MfsJSKL9GtN485SmZIHSF
p0FEgJTTZEM7cqC1qDPoKboMARZ0smol4Rh1nbGQFMRUfMXtL4Nh5m/+/hR1xLnO
FxVXnaQBVO1WsFgzSnuBZM8iCtdOFxdZYuezeR9hRmEemJXk3uJBtE2IPfIxO9DR
60ncL1zProKV44Wz/e86NWSc7KFQAh41bTDT3rgi+21PxLuVi1D7Nq/B9F73ZRAb
nJmXaxCpVbJdHrnac2hKfz2LD3cDnaxzd9S8/NfZ8Zz586koOMZhmRiw8eFxML0o
lGJ9ggEPX+d1Ktm6ksr4kkIP69c+bU9tdEBaTCC3ll0pvFFv3tYnpA3s4Udu1DU+
JKpVfex3/ZVFwG0CtNaBOpToliKuHYOdCWyfIrP+NnaZRrY7Y0dNRyqrfA//3ZTj
PNYYVOY3FHXFWdBx3RqkLBbHHBjKwu6jLYKh4F7Cu03LUDTQi5ZyAV3E8h49Hf0C
0LnzOKRJ9u88O7JkKDNpv9J1x3/EwAS9peWBuQ8yt9t3VPoMZB3EMls04JG6WEnK
EwdtRBHf5kAHBCR9W83BaQZn8laDWImEW7QWFqDIIzE+VouRd+Jub5XA2jpdlkVV
8zfS2GHmxWeY0222KQh87n1R7GQr5zh19Z3ZCk9PsXgm4r53fMAHopI7booRYQU7
smS8oaARDjKkxC2/ubJqMOmXX9cHdo3WEPODbuCA8DXvx6jdLny6KQLsTBuNwih5
sIGI4Vs2N7qkKPTRzIZ9uIoCf/l6O+NUJtr7SpFZdeA76VJ2gtwiUyrwJbLneMDY
XR36aimDfI8djfnwo41d1G1CIpp8N8s1CHAPpYNX3zufIRDw+iigfMlUUSp6Y1iD
rkLI+D3MNQdh78Ib4FMBjMblUykP/pKJXeMdOuU5rLBDmTimWPoXffshHQnJMru0
cM6zo6VZEvJi2kLPv0RlSqe06SrzU0vIdxJsDuelZXudbDCnL+2ZZTUvpKbStAyQ
r3fl5QqYDB6dMXNlsUjyxYUKW0XqOvPMn/88vuRD0wowA5zkhTbZ44RGa+PgUnNI
nZ5MwCmghef/Ix48Mf9NEoHiAEqbh+l6wq9O00bwUgq4GL15EQKu3bwlnsWWZo7n
387kmCNLgkvXsFBIDMIUayUbeamUigFmqu2UKyCQrZHrySKhCO45m5JpQrOiSFDq
DhWXXU9CsYmNwgZiWtFQ655zFiqVwFm/OoHmCVWhkDNS8CeAavs8d+fjc4YeGfGH
eeguzpD4o+QArI/8CC+TUiD33BCfoNRA903tN8hWwJBj/UXs++opL/bqgHz/7DW0
+AqBjNA6yGo2ODbXO4LWo0Z38Awi3vsnTtoBGdQuhQuI6qNSJ07i6zKmmGiPLFmk
1KsixMcQdu+o9UfD09wOIeBL4E9A9uwS2z6TDMTfMf5cJ9tPmeuYf+37U79vLmWt
Gcwpg0evmPiF17CsFFu9TJ26GWVgegcecqrtKi0t4oJkYrAooa/eIcjEjUfo/x87
M9a7ijMhwCU5VwIMwHSaWY3Wo0bbqzE4vMNs/D4YaTws7ywC8U15lHw4beatVYNi
4o3RZ3UWldafhoVSCzCXd4x70cYfY435KqUxOHicZ1sTR+DHm2Ykj3hQs+ENEF93
2v5PqlxexNR84oi6KrpCC9VfPM1qPoPlNNfe1NJ2BF+osf6chtYMLctADbMSPBtQ
P012aojsq9A+VpzpYatijdi6W5QLPLBrdjRp5q/pdcYCfXy/JQyq7BX+yz7olwhT
D7T4eR0Z+nYABxuY4oS6Nwxuh3bUTiXzADVyDiTtyIJe+qpiqWDQLdEdZg7H7Gai
RilKIhzrG8uUrKp52Q/e3Y+wZMjee3DPjh1a016Y77e/2UQuadQMMQAujBFQzT0S
Q/xSZVoxkM1TyjeNUfqjVlVXEC6QZjAnLGhpg+t6268seobZbyt90oQOYr9GVhKe
7Q5SajXDapPlp8mbZv3dMG13Q8NGT/Sj/AnxcJNyYxDhhXky7JYGtXFMoftr5gFn
/ksDI7jV67OrXOKhs6oU9t0q3W4stNyaDb2FXMrueoBUOyIQx74AZLnqrBDXQHK5
iGBjnxL/A2bxu4z30A26DKEa2ENr+oAO6QD8CgGstWChH/9k67jT57OvDtpTwW2J
AALCJE8ozRRDaO8c2OpIWwZTB62e2yMX3ft69jsq2WzLHNk2Z2Zd4ptgs30E8OHV
IoW58+sS8ExeGq+Z3COSqml6lL4WxiIsFpxYJPlPw684h6HgSqCZ85iY71Z+FjJn
8Jyt1F+nd6pfiCSo3w5A1uA6QEVXDom7JpTnHNVUyE4qiSWBFfaJC9zd1egyHFme
A4EA7WoN2OcsYSnHFNyF/pugwf8M3O6vGsBNFuafGes8KoToD3chUjAsc/RhEyP5
NjyXfc/PfSjQ5DtrX1delcARA2W+ND72R+rtuS0ZE3G/8IogogfWALN81LVOK71A
0NW9742hJSyPCaItzqxcB/uyHxvbd4UwvPCv/gQ/TiOAXSBms90zbhP6ga8YEInd
H/FzLZiuaWelvZVrL5r9s2WJwGFMIuG2DbtnzGxTZyU0saw5KWenU3PjLXHgmOtY
nme+oO7t6EMGYfRLoUKr3wKaGWsA48tFBCuoUnwXxAHZ7ajdgAu7c3w+P5Uyg3Xv
seQ8QphVwHXJR9jFB/FQaGKAw8WWE3lJyZRkmybdHZ9Vmo/OXB0uCpfbEVkj46et
+Aj0pJE3ASH+znYxy0cIlf7FkruyhlVTbRFohE+zDCe/Jqzimp1BEAsPz6mTh8C+
Zl1xPPLaYQkq0U6nJP8Pw+LzoR1JCa0eOewjfT7Jrcrmm88Ly1BoOIpjeh39dPGD
3jHdePTWszxK2b36SWA4qN7dEvK4r7FZot4Y/ZvR1aO7zGWRi8aZ1/2ofxJWeXL5
0RDUR4kZzH32kLih0JqnB8tWhew+WRpI5YnM91mS14t4XNySon345dGS36+7oo2R
2SH0MwJEQM9NOJjrnGqTjaGxmIVXW0pSsusnI9dVqlx22FM9KfBcVR9F25wDWDhQ
CiYpSFgMZQUO5+MaOdwDW6IgXn75en5n0y6oTs1LBfQMW5hzz+qpB/MDr5Jb9jSl
NSBYgBy2OiyWCbYGB/GMHVNJMyT/ixQH0OousVgJwLvp9BCkXexhBzBokMaRaZ9B
003Yu9MuAxKeFUMWL2IekK/DTwmlokHez36wJpR2NWEluVTkYOchdObZNKNE9rs+
J5V9Rribzz7nzIPEbGSqQuywOmDlFTyK+jZgre1SY1dJwlHbciKxO7Ra5TDdzsnF
/xh3dud3B0mybpMuYJhwCxaXWjpu6TI4QYgYQKYWmjHEWuJPUDQ3/IR4V4mjpLr5
DREIOHYC2x8KuZV/ma6E7bD8L+NpeNoVz2XPt2oc4p3DkQij6ELepe8MPhcbcPCn
Z4SHhLLUORg8GkG5gLudAi8vYGRlpS6RQdMMvpmtZ5es4vjunq3GuiLSPJ3pRpys
bfWbnnTheNZJTQGx1z0qDymYvXmw77XBH+puGj04dl7L+HpKkLAjrLcSO0FqHcyf
Fyf5ym2medLTBIzKtddoEAUCKCB5WyhamIt/3XJ5C2OBvcbj828bMS3Ctb1H5Dgk
DD9HDolSHI2Q7XvqqLKN/S+Gu31zrptlrS8n7oJkoFZLRVGV6NVt7qDTBLNkp3W/
UBWQp/SPDG1/EudT01QATaRUQdOyRAjNcAIC56dCJq9oBQjZKKV1u4DO0KA8o/HX
b4PQlrGf0QsZlYFGayk5LUZI0ljeJ87VGz4qKGSvF6JFRj7/KYRK0vjZ3M3Vyegg
zPt2Lez3+CIJ+NhinuIUs1PtTGI3Y/xCQ/oiuDfaY3rdBffp67vEzOyqKzbn/l+e
qAxhk8ZbMXlrrHkE1zvtsD09yfZBVbmUh5UjYDbtzOXZQ9URL6oeSsJ+lMsfG/v5
Fzmn3Mtf+ZtLevsLX7HtPBoH+iLWDrhxsW5wTgcLLUk1/PRdE3VIBjfM60NlUhBe
CeTCBHUgJpfUn6GdRGSDeE1CZTBh1lt3HGLc9ieSjqQ/iWos13apm3s4QzK1pPbh
y+vmQmEiaxSqTZuoSeBLRqv8rhTthOwjmE9bFRYQba4/tPuDotcgQ8e/deChkcy0
QFklL6Wd41i5TqF1jppG/EJ4sFcXroY2vIcWt2y+naq/cJ7hdjyDOwqTdmW4Dt8P
FXqTM1zpzraMXZQh5U7ruxKZWB9VUi5X9ofjz7Wf5XYRKAlvc7BsacoCE6XRjkJb
HtTeXd+E4LESEyQKDUiRGuOe89d6VCieJD67hV58QD2KUNlhgVG3i2vnoQXXaXFO
L6rPeY0hRIK9M5j1v1BP1rrsW+2NecbU/4um4YjPLhq5ojXRp84yd0CZnA/lHppS
vIIkb2q7OofVAjbDym3/zIZujJ/CEzXXDa+DyX8fXtiMZGy5ZJbFyshkoZqMd6yd
s5wCbUirL0K8y96md4Zkq4aYPMBcjAyqWM2QnYzMGDOAezhihWu3Wj+9+UOa0cqI
T0JNsNS382l1bdzqeBdx4aenwyqSU8Qtt6n7yaQWF4x7pprcMdct2FzPQm/ROphg
zb9KtyAozlzqwgzwa4flAay2vyCM1lgIi5yhm0z2qh+Ue1CYJb5RvbmLWBvq6wWO
1TUDEK2p40JPNxrVr37Fm4l5UsPmnb2OxQXlBy1l9KI9MJrNe3Y8UPj6AReKPAMv
ai2MgJM09e6HbiiW6T/dgUtdzLphE5j1FykCmn8GSo7r3bpeYVqOeyx40sj9k27e
nJkFt+sUGEA6Z9T4z0SZn3GLJHwL+3j0+WajbFufvQs/1GSoKrNi9rcs1K7jppTM
LGFOjVBXBYErDPBRFDkHcSJl1Qf2yccC/YnBs/r3YpJdToCi43KGDX0rIxD1szSR
BadNPR0x/xmzveCu+uVDRZcdW6LSOyLX3bTWiqVjN1scsiP1l6gCrtpj6A6j6DPy
pvG/9ENYiPT/eA1FBJ9qpT9zmbpLTXmcsAtBZfvR8d3x2O7a8zdiEuF0/UvoeCNH
tqsQJVjfeedgLDxTtVdIGCFQXkSFFuCcDKPnlO6E2jYs1dxOF/o2DSHOgNTWJgmS
d0JkZqvmc8x1Im+BNY37Q1EiNZPzg0lyubaev5u4Rak7+F16qelYV/FFPBGhtLdl
4yU10dgBZb50djIvCLxiNf5cu9bzegFD3ItlhgrFrQnxTjNnYRCGEsF2YMgndHdP
F+IoMm5pkgxW9gIKieP5365j0c+F0cxuKofRZUodj5WXSu4EjRTG5uZLgvJYpArj
diGr4hHejRxSxjwz5UaFp61VWI8g78fAL6zG8lQosBcUiwzcqovgMJME7YWE0V32
Aqpw8lcwPsUuk26IDWcE52ABSehYQ4yUNf62FwFIxb9RA5HNZM4idjHSs5fwoKTj
HrkAeUNQnbtVZtA/yk6y8g4dP4xlppxSh/Pk6HK5OX0uM1SPVK8dqWs2dRyFgtbE
VoiFiYLp6fFLlNBfXMe6TxPWhthR8p2elqKe11K/9v2Ckc6LbdVGd7NcUvLn9Srj
APSYwz6EnlXbiD8QngUNtvJSm/iPJUbfsvYSXTQeepwlDGGQvMM4Np5mM9XM//B7
JATv0lXGavQ/mxLMZ7K8L2WQT+7gJwOTg1AnDmZwf7+iLucy0N4YL7g8V19owPuw
8aPAspn/OZhKIVbJkzrF3VvAT7mUxKLnO6MvnqNY5eeYVMl/ibBwq8LOjmskRPtm
wcvorQh1CD9FzQpTjdBZNSAD3TUMt8zWajvPluRxjn/BHweARd3f2gRrlp5FG1xQ
LYkdQF5UI8DYvZhFkPYq2ldxSzJwQWsCxIw0sK0feSs/xYY/+sX9xaJsRjg0V3z6
ySfAhPRSgIgf0m4L6hyI2Inu9v6Sh7VViOzPdlb8EBfK2+n27PBYYOPcSkdAxxGO
9z+wk2LXvqsILWrMME0szBjCXtbGC74yy1L+d0JO2r8CYaS/n/iEyJVfBvQT6IlQ
RZ1HxhgC3KfQsXtfiQHSehVyoqF6qayc0jJsaQq7ELAk3lVTMYXV6SDZgwVeTw1C
E05Iz9bDbIv23HdS9J8Ot1Abe002CugGa+KPYJLradWppkBCm0+BiaVSyyQNCBMx
H5YeRm+JY9QlxDk06WFIgYKnVYkxqeM6NhcziQcLszK2khBiR2JKii4Df8yLIAph
aVgmdxkYH7WDVaXE5KWN/NHlXwdMf/kt7eSLipEksVZ7ZnUk3Lg3hq0RMVjr2KwJ
OZNJvRFTKpQ4L5HPmsRZ0Czbd/6NsNoY0i8OPH3iE7bshVTbFd4g6Vt9S6oowvNv
qUe40dbccFN3qrLMvI83ApZakMPTl2J6V2Kt1bLKTQhL86S+l2M8hsOpgVZsstjm
Dj+mmJpdmZwYQRclyHo0O65HaJZpcy7JUY9+k2cB4/g+ZBT7mNAntD2bTGiJB+9+
etHUNXaKr8vL4V+KK3nDogjNYmWdpIQQxGV4r2HzSPTWQ6AoNxec/w5aOHqO/kV5
3leSM95g1oS6mKCA2xVzoupEBX7+z/OgpmXA4kzEfYvvs1ATohrXctfS6KpR5q2k
LcvDY6WQvYu1hZAt6phq65inF+9h/JDRnZr02o2Aig30NUtwS/xyX1Nc9xqMhsxx
5eLMfQR/5pTMtWyA4bAE3eJKnVRhY15VMxXc1EUjiGoT+2Z179LwZalDy4ZOwa7u
ZACLMrNEgz+HjWdp62E0r6NNBwaGQxU/+wQSVKJqUhUIeC+KT3QKJNKw4z1hvGAf
Cv1EOn1yqtaLD/yCw56+9hTOW1hVv7R+/WOueLHdKLd9077/N3eggefaEJb48qCF
N9KaaA+/aZd0BnNutzG6LI42NslAWd3CsU+Ad+tnOQch5f9Ae1rrGUCov6EcYpJm
HoOZozZe690WROxvP1GxiNlr+XkV2Butf2xFT6OCJ1tJxzgyOdlaB3SqdO5gANbs
6avM4NPSF3bDV1CndQYBCyGRPDUpxPEUz8JquCWVJHi2OF9p+LkafWmbd4kXReQz
soevR3qDBNYbO4CccVB7+xrrLsakwzRia7ZWhpt9gPk6ZCtlXqUfW1xgWty57dwz
spS+Zk+1kvJoEZfuI6hS/vgXgA2nKZAxSuTLWUgc0GMsdXCPUlQ44J2HQwLo/CR+
TYyKP3+FQ6Z0JEIJfIYc0c6PeTf+7Zh6IW3rE2JeZewHG19EGm9vXyW+jPsw9QLg
AV2BZFbP1opmKrrnCvAhsNweNtDJsA0QQ22cx02vIjdqlG9DpE6n2JpFHcJxI4Yx
qjKMC49JSVgDaTq7fmk+5FhuZMUiZYHKVne6yMikCNWOkxInQn/4WKGcvBU92vC8
aRn01GrjXgQQ3Mw1wXfQOhVY8eCL2Y3Y75l94oJtO2PNKr0TEoiX6JAgVFplyH8p
cxRGiuAiDgn6q0HsvLom8fj5up6X/X3m9+nrRi6apVjAYGFt0WRbyaIF2lap/djW
T0jsuZEFeeHue4GrkmM2p79jaOq/5ZC3CT5uAdSWZw5k22fWPW11J34lnFt8PDBP
WCgteQZ9UB+5smeBPou+nMU8a+vLk54qBZDzGuNSYRb6urVgaUj3AR2bE+MySPII
7/Uw/43VLByxwP06KNZ5RRgU7ki+Sq1oYbcHHelw79HN8HPyTe+5dcYz0GJbN0TS
mQ6JhkDxiPtMa2RGGEfHst/j/I86fiSqHVD8cCsAcZjjr+OEoL3npHWrrspb0hhA
YOwmQm/y4LPhgikQJh4G3Pj1arZesKi7rHfclk9DgnGcnvCUKu+3rEn9NkMDRYmp
2/PbO0EfqknH87puTsGxmziaFRRl7VFok3rhMh8Fz1z6OHGFYo+iZX/Q4u9P0hLS
UI/MzXYrIh3G/Lq/DDqF/04rKpehWMKsZaJrGJfFkx13Wh61ba3e46uCgMaannkc
OUev0EKnzoQji0KdMFqquXyYxHyZXTBmSfj33FwZTN8dV/7JTiwDIZGHnEXComHY
Ce5bcHQNpgVKe9OoqfGcLsUJN/LzgZi6t85N+2kGla4QFnpE0mu2DXjRHEpcNcYC
sgXCHvW4sv6UGUy/a0hyfca9zNB7ewLeZ1YtB+ONTmXKX72hue3C/ldFVFdlv6Ku
zrYzNF4nF86EP4g/sX4/qA2eBxo+hgpdhGO7ZaiaIc9o58fhoiFMV7ijqJp1UQ4Y
R/YbnRkTVgXWBVQSWXEn7AKjI+mTaIfZPmtjVRqdHum+P69aIZ3Lz/1r1GAW8r27
9QugoIFZb0fzSJJl1aHsiQCPAFi9DNPVH1MQZOaVeIkEszsL8cOmWrTHb66xzSfN
z0r+duKVWVl+CukI9GPC2ND9R67764vjJ+W1tRKQddmR8euoNNsxqYmQOJOauLDl
SZ/StFoVq0Z5KwIN2bxZzKI2fnIG579w7OuM99RDmaWnqtjzZkinEiNlxlDK4o2A
Qmiec9MKTeMNZVqZcWoBzakFTM1z86MmxSiNfU02wnCn6C4btLQY7rq0tex68RVw
nGFh5p/lQvlfd+UM3phHATxZVl6AC0xwOnZGe2UDaQXqG4Bvk4IX5dn1Z54RgBS1
VUpDyxRqBnYqCG4ebGJFDkWoJ4GqyVHPTEVzHncf6cru0LhmZBGquWiXEr75wQGh
SHM3V+4UpsQl6WB3LbuBcuI/361m/edHJbDFRZfiSWj2snwaewuSgR//IEtvdN1L
mE6v+U6Lh714sNvsa6h2tNrW7qBn6SDgjOE2VHxOmlYg94uHvU59LMDjRX4moX5q
tyyzFAiLkIbS+SV/XbDpXWOZY9yaR8+GEtSI2V6ijw06irkyxpQGIaP1q2lG6UhB
PXIuh4CfQXEiRtLrRZ+0/E6WX+Va3lL02T9sGEkQFzh9ehC24Pq9rKgENoktkp/z
GNbGwX7HIlC9tqFu1hRSmEBx0d7b4OE4JXfJOPmtXzBiCBiyCmTE+1q8M76oPu81
uHteA0QudGJbGqsF1iUQ87Vlmvy9MdvITP+BkTQZ4ABOysoTfVekM9VlkxHe1BmM
NFYiLH7sXyEHh5B5l0RepU0AUOgfQQa+LXGj7K3TCm5fROK2bgL0NxZ+O3yRR3az
z70qg7sFswMkkBZWFuqaKa92i846S8atzBhQ43ZQpm415AWfNOazpqM5+I9zM13d
rshGp7jII1fel4ROXI93FQO1vMXDNs4ndiZaa0euGrpn0iU8NVNDjY4ULreNQ5tG
`protect end_protected