`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 26864 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRvSzIdqqwO5JLOHm2ufP7EpPiMK+Qq1h7p6l90CUpAjN
g0iC6fuMZ5J8rgquZavA9P+HxYrPQ1PvXp00D2el5eG8+xbP9hxsyY8LH+tVrnCt
XVMZSfm/5bOvsaapYhQuit9qRZ59O0DdFAm3LB8bVG7tFe2frg5oe4fuy7NCMtsV
nO58f6vQN8oX5oavuypVFrZhhlVYWPql4sVmryeDQayK9sHJpRx0ixfNobiMteTi
nIeaQYcCAnWV/xCU9sdB8xzBkFAKmamH3sriujIJTRNjt1hnJSTZpJZtLgkdO/+g
l78q7EV0QJjVO+lyhLM+yvzHIkiXIW+Qw1xHaql53gBy6rdIb03CHVpyMRuyL8s/
Ys1H2AGG18dmk2x6k9VhN3IJ7iXG5ZtSMsbP4/9qxi/Yf0QqGNooEv/a8LBhVwbL
5n29NY9Y7SXAlZFV7pqfTV5n5ObR6J/dKMp9ecgnZpJKftKl8V46GTjSQfpOE4/q
1LdYUg1EyoOW5EVZB2a+3inpTJl/3+WCAfclLZexIlJ/bSaqxmnOppmxC6UCBwIy
h0Rin3chC8sUQ9yw3sCj3OWUeWTKwfnv0O4KSepitbxrrwPIOZHw5ozNylHDGoHK
puhwZ43V7hq66GuSKi5serfh5d0iKr9Wv9esB8JMduWe52IhRCnalZJwk5XF1ZG/
b5mX4++zbARsZOUULvy86uC3EgKMlI1PXvcBSfknex4vu0ufzfuaq5RoCOF4jij3
SKHfYrNuf9/vTASKCKmIXQksYl4yNd8/4VLgNT4wKSdJUVCXnji+7HMZHefgHlCP
lepP+MkwkqymwmhuFpzzOzdb+zpmUzM1jvAhqxY6iKMn2WaKWKz7AnkYtfXHQCU2
EVbHlby0t9FMBMVV3620M7PslOrfC2bjEm79BYTy1O95s5GkFgqfIMIEfu88YlFw
I7mOZQyW3MutsfEBDgrguuf3rUJ+oJZaEwaXlyRDOVbjKXoO6IBpJWSr2Mjgj1bX
sJdfNAMQ0B3QILzGB8IHJNXK9r/5pY94ZnD6sj3345mfB/O4CS+Y7woEzpbPkaDz
noZ8MulHWZWF7qRfOVoz+Y5cxrzYY/KxLba94h1CtTag2JHOHmq/NucCHOLc7zS9
J1LGGC8lXf5cbMJtlUQXxoutamMedJFSGbIIVc39gHUqG0su836of2mIIv2Ysg+r
ZQ5qylnBj8wofa/ebq+yhsRhZm/FUggq4rxZ4yYqHiqVQ0k5wN6cVFhiWCOdkilE
PGmpOayHrYET2CuAx6taKWrnYY7HdgkqjHEsuXvS2pLDgOV178kidbeyrwZlP2eN
FVvA26sVKe2AFe2aWQ9imybVPDVoGxVGEaiBVjzjgARqvspXNQ7wnh1MVhXaFGmo
o4k+Z3Em2O7Rl89vHbrPWvVXvoOyz/8baPwifN21sFEMGqybUJpxlUfPRdjr9IAQ
+b2s8qsr94fpHufMIdVRCpKILcwOWm9BMikVP6sAjkRn+wPIfO/Y16I4qhEC2SQ2
vEdyA53b7HWA/F1qgmzMI/zQeF6pJ+wKzLiZOLclRkMBZ6TZwBwIrIDFoUzW9R3D
SCztO3OMyJOoT/oR/JWuobhKfKEmND0F74RtAni2fnWg+Wafc8rPCVQ9dgzJfD98
TmC3NeGUCAbARC5ha/EC40QYxLYWYPVIEI5bPJ15bCoVNloMGvkqT9xX81MMVJLk
OJM1rWwr4vRLDWGheKMX55BL9J0zme5W+BpbD88uPjqK6ItDdOC5qn5NCtABrwUc
shUZYXcak/t0RxCgJ5iCgdWRowl7XTja5HYoVawYZsUD9k9QZ4hZiOUaq6KJ73Nf
2uDy4KyGzWr3Ck86k24OYraS0oFpXpS8NopGthcjvUB9/ZR6UBx35S/Bp7Ommzgy
W1vLi3DcFVTAkOcj3XISVosvrO414M/umwf+BM8iiVHn7rglD/DJd774wVM5GaFY
rV6qD33oxt3SjTkZTpeJcG5VwwihIjmI59OjGeyCSV76GbZz2Cn58gid0+cjL1nV
jzZksnz9qgJsa1V7SSFLR7QkYyGMCi2wbG4qxoOk81QMQNpt6toz9iT/hkVgUKuD
X49wT3SgevTy2F8PWBtUGAyZfa8jHHJ2qy5vrnnI+SIX/X8EnOBhh728Aaqrwlgt
Hh8ml+52ql3zmfvkUyhfLXLFhkmtfvuDx5I9bcFL9UxIgAOQcVuXGWYKOFJbAk0G
v1mls0a/Nr7WMn2YvCSfsipcKWN4t/pedz9z25IsIDkg3r1x+8ks8gevFjOPg88U
dUpgOJZNKlRPZOennngX+3d61odNG/zDQgzVWKaBXsZ2/TsHQY9Dk1I3AxCNShY8
zd8Oh4XWkxPlp9jPEqYfwA4zDPWQKEwuGxFnSCcIJIDRNrUGb8DRAtMUGc27wROE
sqr6IMMnq9BUYxmoHw/KL4Xat/JPIJRm+qq1ZALDxkaQH+yQDLZLtBiRvCnirB9c
A+BhjyHv+k9B7cI/qNb3fibVdyurRZDaai2Thn9fbfOobmLl3zNSb7ywdIBalhXI
T0NsfNbo+15Zj7KJOXRUM4BcjRMPZISPI23vea79aif5FBPQyda6DpZm8QkXpnn+
OugM9B2LmYCo5lCVe6ejJhbQl/FEIjT4DvSybcQnAPmdlfUd10n5179VDIALr5fw
FXP87txbe0vslWxCY57r0WbKpMDhnVeEf+vAZOh4yuCJQqJnQ3SywTcMrQnOlvuT
wlW4mkL9BsHQTflLmNBs3DGERsUTdUJfPdHGzSJh9vTSyKhgN0t+hKBVXK//yehN
K1EfG7A+05rdHIjBy/2hfCxBBmUslh+KayLJxFFFzo086K+FkbJ28zr4+C3+iTAg
uJ/5J2Ha25hkjEtkMv41WdbuVljt7EJKUeXEMmIh0+p57bErD395OVIgfWp0T4qJ
Tre3nYRVdlfODdSYVPhgbJ/lWMADn3f9Vce/5nUZML/egohiOKP9GM2gGtP34jaR
XefM2wwngnXYJdtSGy4Pyb+VGJ7hcP/4nuXbKqxa9ZnzMFq9kJ6IGRmukqTp+HRF
iXxHKHIfhMFZyRtAgrJVJha/NoWTwCqe7ve+hexrYD2elFMqAGRx2RjmVU5SeN6Z
qj6b4Wy7adlo7sFsm0l8ndEWW/R7JIi7LNt3TFUAuPM7OBdutjnd1HKw4hQOZ081
vj5JO2fj9unLqhwK9/FqpqUwl25LD7i7Meqdx0EsBvLBfTb59PbwdJFFuJdzs639
4WNzpk/ed9/BgPWrStPQTCh9azQ+fAHqEiJjAip7y+YbsFiGBPwUL55xxTWaI8dI
t0rNGG2IPUJt0OW3vS4eikI1swMpYZ/xKs1t8U7Hy8jD2qx/VtOYT4qf4sGUb4Ke
1V9M1Y4btc1omEuJxweavLBZ6D3PNkzX0IHZVgNX2q3QdXGi8IU61zKMSH7zYxvM
XXl60+A3WIS5dCSKFMY3fbO2qlrJKR/WKc2yGK0nRqSHm6KjBGU+3vja3Mr9kTor
ck4CZph0iq+0dzrJayVp+dCgpShsau8tAT3usQhZ1MiAwuIIzKCiqeUl3sQXv9zo
CfIQC2NLYkVrrcsfhdvb2X9PWYjZ5NQG/3l6eIfOawqIMClGw8EpjnPJUsei0wYC
xfpL7hiOxd0le19MwSVI7IQ77Lw05Y0Id/BYhPxNvnmW3gEoRkzZgMLKVgZPWihI
hV1MacKERGzz2qY5YIi5gV36JHDUsHW2wWqEv1r7YVuAvKwddclm+AUaxgW0BKNN
ZSTmd6+JqwOEf4F6evHlD8j8qgtDl+O7VQlQ4PguiGWYLQ4IPgHOixCaLiTX7wls
wI1sUz0c8po8fnLlk4+GwEgzxpz7eHcRxdP3otDgK1cXgVol+M7asOr7oKqQTbY1
LrneNTroudHFrQC/fr1bpm/+//uG6ZgFuKKmUMs6rYZ9sdbXQ8jdVyHsPySvrc5Q
hZdRT5FHQF76D811C4zcxgu8qH7LF09HyeEBue5B7+/IV7l2jwKvAhyMrIH90mPO
qSOSffd/B48BkfTNIzoDOIOuaNYSqDCpCgwjjtaapNoR1TbcZWjsDwsl4dAwQ29/
H6T/lMMmKJF6VG/SOqrbo9BbVSWMyAcTBsXV6X1a0V4xDK3BqyrdpwKeZNYULwnf
a5mzOYZIJ+mpr99nUdTNLYC1KDoUuo+v3ZFUz/ykiFEhQYLV4FOE3PuR5j+IgkgB
+DZ5QigfzVIUpLMkVBLt5y1x1HRc0qU53YZHEewIP2uG7hRB9Sst0IH160qmekis
XaF6vSOgvhPUeq4v1Ik/i0aYssuu3A+j8W3LTuVo9hr7yxYAiYlnMJHV4VN3gRNt
efh2m2tlTyT9xTDv4xO/8ZH8cPlADbBhiVOh05eCfR0lUspunleLLjDcDqIvXWho
JLW4DrX0OoWpKbesseumbqkMVGdC3TY0T4WJfzi407ddU4TZHgsOlwvhOrjU9RIb
tGrtVivZbm7aOwrD9l6R+fnxAws2HoJE03XE/UtKrtuCzaDeZfq4vKS1lE8IaVqO
4W3SU5UhgO894fKth+RnLkF5NSy3zDB1W9QNpxrUkMBLztxPOtxSmHqIQQBFvb2V
cHcBuxtPprg5EN5FmCcq0soKDQEJCBqeftPTdNVOpM+Pjasq2NsEIBcjlA3WW8a8
C7i5ieteXrs3IYjL2sfgwFaqqNSruTzueZoe+kQHxcHpQFpFQFgpBWL9YzoS8ECy
eUwUBoeCYXVV4DTJ2h1IexmR2Hbi18o+hbeFsRYZlOCZJKxG9ypWw69IrY1BQIC3
PYyr6xvjHeTHPAVq4B+agHSoZ5IcbQajX9Xa5IXbyKWkTsS2hYH2Nuhwq97Rv/nb
yJTr8SyHvHTaynA4KElJZU/d+OoAAbtHQFVJVYLGCs5zuhBsLhmEo1BfWcbBIOwo
rOe98pTqxbIk+Z2O1pFpUguY6LzyRitxqKqMHlJvjsJoIIQ+rPRChou00DaDfVHF
C2Yj6j8sJEAYQ8o4nH22X1tLDwOig8CYKNodfGIZPqP0IIsF5IjOzPRJTUF/XrE4
2cAKidP6HNSNXrwGbR0RXXOvZ8HGHizLEVB+34oZ/FZTSJ4IFSP/ooKmtCFp7RVm
asWGj46RG4bki7bRoSRuhs4POi/4i3loi94glEWPyLCqogJPiK05nXQadGuce5iv
VqQzuGEbQtiFeRmtSL9ZSwentx0eD82tEV1xelehOZDxgH0F6UAtehEnL0s0MJBn
zFUK6JvYFEd978z0fJgrrNlv/KOKzfl8uM0A9eeNNoitlfxPJ447WMB2IrPToMpW
FN06R51kK8rKRRACEqlHYaaKLQdKCkttR5GLoutjXaCALOJIl433qlOR0/oKF88t
RGD6f4Xd0oeChNe5wA5Fo516wsNJnw9UlasnTeEMdYk/kUsXcG3hrdWW4IqHzWfh
b9ks1hfXaV4h/5f/dxEqf00OK+QRlTJRkLU6NnnyWSqAbST7gP6gWyRSOpzm1V0T
h+EvZ1FUMFyLHCsYdchU55N0er0fkyEAb+gLIbIBsvKpggFk6FkM+bSOJcC0cCrH
G0JdcjiVhWkGTdWMNUcouW5n2iOfZAnMOE68FdcMmMwYnzaZ2P+A5Hrf6MdAWyE7
diio3UUqSAo2XTBS99c9Ky6M3rkrlD+AGljTxjGe246CiDBQ85c4lgzXRK94RIKI
pPJaW7W2N/0ih9M5UYy9O0FZUSy2E3f9/2LA0HkyY6tuXTG8V6wKW5A6Qz2daFH8
IQz1Pbytt85vpnesIIDm8zjCRaU+hV9yBc0tMBMRr4TZ536Q10+P7C6XtCNIKgEO
32I2mIWelCR7j5mNedbeW4BqpTstjYxmwnMIzt6+wcxGLTZHPp/ma5ltGJGqIvGt
dJjBcy1sYO/9OyvbyrTaSPvINa96Kis6JExl4TZ6xnXCSoA8PuhK4gLdFf/kq8lo
xSTE0r+qyqRsMqEiUYFvF/ln+S9daT+1Tq61v7UkDMHaOIm8y1iE/khVvNWrIpKb
lVpivI9B/Zd+Agn5ID3jpb6lxHit+TpZNbsns0m6wzk6KKDHXUeq7079g/IJCqyn
vX3b47g8qvBhg4tnjXjd6IzItHgZpshUFNIQq11y+FVIuMHmcueFflwwicgooG5h
2/p8fNcKeFFZIkptYImin3O8+5UtYgLwSJJ8k/zEMbH6IoQX9rHM7NkX/IEimCcG
w8I7/QaZa9YEdaEqVxYutwqZAF6FWl9m9g8j8RE9l+rBwu4N1ULfPX2QS/eB2gUl
2WlunZwFLTWixGrLecen1fRSvNqtIl8n45Fh/s4dEhsSQhmRtzuSv7W/Zv0dy+Q6
vAjZieMXFLZ+HBDdL743uXGIQuu+MTfSnZxbZ74btzUwjRUWi9SxlVGTszMmau2f
4AjmsWLgZgbnpUsNPgPe4a4HqdL5bKiMEgOGpAFjMaQw5SyRQ92IxZHwTWCLfu3V
WriuQhWtZ6x5/GDXmIQdz2XMbdIODIYmYZYBrqC1LK2tz49ZzpEvVMsySSAiIq/2
HMV7OTqusN9k+NWhbqe/JbkaKt2LXu5sGhdDnYd8tySLRVByGWrZucimJldijlGT
TN506bPEJMWgu3xIjrUWLUw8PVsq2jvbXabSxqAHQ8k9WUVJfKAu0TaqiZeycyt1
DYERZ2D9nVCDeW2ZnGmcpPLfv+eRd2b2BhDWTUg8eIB98yVmumP0hdmoYx6+R8xn
PDyAVGdwkiYjVTyoBihX1h6TS+GSPFWuUcu2RWAVFt756GgvkYlAF2ut/3imLn1G
gWXBGfkqvlsbuuNwqkoIbj2hOLWCrBLkSPnQRou3K5Z0vhWK2sqSpopo/a/2ouy7
1U0lITzIRpZlVSjjCsF5xGSgTTL5go82I9gTnWn2z11VaLH6/bNz+N01g773H6hq
GjTJlmM5hGIFynPrXCa90w6V/8q0CS5Bekdkj+nJVdxr6cxVh/bwSXBT+QQf6v8R
yCnnEI4zJbHNbPPf6TrSQ1Mj0g/SdlTV0U9ubghu0qPcBthQm4TDSCI+cdqHccEw
vrhUQtydf+ujTOANroxsLR+hcyGgcu6mdhhPFMEGq6Y5fn02Zo8ifEmolJorSfZH
Idda20OXiDvhu/P0Y0mRF8Fi7FYyV1SoJ9l4T5MZDgV72jaGwmvPJjFYgdH6fArS
PYr+myYSyZD3uE1jtVucfhIJx/DIQRSOZzripIQ1czJ5hwvIoW+AoR1Vy+Lw5aVF
59fecfh+i4nolyCzSZhhAVdxAh76aDEaAWggqG4uf+1jhmrwSqE0CMQ9SJZnT3jx
RWIogznkhqEm9obWvjuGjC7vwvSOgiPzDozAkNv3Fvbpr1YMB3x1yw5PgssJSKxv
pcEV6i0DFsiRHKaGMBv3OIVJ7lwgq3vfxmdku0m1DY7Sb0tbhzMMOkBA0lwIaQRa
0zzlfyuO6PP3wNaBgKkAnQCBBvTMW8rncH8pul28sEo0h3aHFEjeBNBE3i8LBuLZ
R+f+SfPgGZro89ZeRt+ztorZWj6Mct7QkzrzbSysiKRhMHWNzIut/4uQvGldtNLj
YfCfT0LhDGwh1lEb4NlqEaeHt2qw2IGfA/7g0C19Ps+lARGnLawEwieOtNT8CZAD
mjWpZHO5VUDybDyYUn/gnjaDgGInYqtAxO2lwMfzCfSIBt0gFWgjRVEvjW0vURte
iZnZL3EiUScKh3IFXlbOCSq2EFSH6nJxgx/zbYhMiAbioG9ye0JTNk8nt/Dp7AoN
ntMmFrAIumT6PwwZXfEqA7gwWhdGIvp6PjcQiabAeICQoHBZl0OD2L99CVUV3PFW
yp0z7cxKcIIOcNeobaqx28e0ZcZXiTUXh/bJsJ/qbX7kZbu8FWQVyBdRR+25PXOM
+eJWqk+Jf5Mq04MyBsy2Zi1Gn9bf/0X6HotMGHJkq3gDLCDUFF22HKtr7hoy6tpr
8uU27ZV/KXN3LQpusyHJpg52iDVARWRgclRExSkGt0JaH7Ne2IYVJXB9ct+oXFDe
SPlZJRfLwQicr37f18W4nKrqwjNkqnmpEdDNIEu/qwSxuKpWolgXRPBsvdLJhDSa
j87HhJEjOFSlzcxlz20362qP69iY99NjKrRuhKkLU0c6chM+5r2lpL3HBtJscqxi
6gowHuebF5IA/59eYsFsAgwTD13biSVkdkrWiwrrnmB2V8bSSRcS9OUymPJlB7/S
Iu6acxysFo0bo9IhCX1I9+LTqNRcNYzgusdEmOdM6H2W1tPHi6dT7CJvhYeGI03c
Vswk01YVUxWwpeWgrg2kLBvmZjd9TK1G26TB1uZYF0D6L46Uh2u+d1liubQuGItI
mx0IoLbMtnCYaeECAGizo2A543c9jI/9IAhpfQwtfZfBJ+QuR6vFfZvgko8QyzHz
FYxtfNUzx5AtW/9KrQ4BqKNEolMyCcVCEzhcBoSC0XQV8GnCotoEB7lyvxfoKMza
nclz2m8zkZKiJ1L8gw5Id2A1Z1J18oZeb/qfKn/yfhetI2X56Rkl/5SsG521Z+OQ
p58LqJlO4hgrNMNk9NongKfBkFCWGjelhd1dtXTmCAwGGY2Dx5nhZf8yaT7kP+FI
I5wmo2vSrNjwgzsZ+A6/IqxobeesFp26I0c1b/WQC0r7KpvSAo+2z3qKP+iBY7Oc
Y/cWY/vQVv0z8lAbWNVgD6IMuvLRtal1BjjwetbapiENbFkk+SUEatRDCNNaXe1h
tIZJkHeYukcGcKX3IxKtwmLH73iQuL75ncLjtiFNLcEwcdcnGKvFRoHB7dQ7Oz78
YzFPDa3QQRn5QpE9OILoBlRn3LyfwhowcqPkhyqgLzgI+wE6grdB/MneM9+E9ZgT
i6Zsz9kLWCyhkkrbGMxfzw16N2TSyp+4m5dLoPnUj5RYqdE9Eb6UF1r3u03Lc11C
LNik7m0re4YoYvgLzY5yevTCDdGHkVOSU3qv77EW3vsb3Ph7i3Omk9pdDl3n7OTr
ruaJs8LqkxixXGfqJhRPwlv6uHzGKRKijPpnANbRDTz9mfnEM+h7wut90zvtx2HT
S9p9entiOddfEVhD0Obm3oEEkdQdPtp4F4+HObxkq7Xlqy+pTtr/tkjZ6N/VV0Q/
ZAGczt0hVJ/z5VymH0ZcaN/omcILzVCOcW7ALebpn17KwW19819BRf2ChOd7a5d3
myFwkG0rnJn5TMcKxCu0hMoIl44GksUAsxx0lB5m8mq5XNoL65mOV+sbVEk9SEFa
SNk3yAi+kU61fQMEOjcnWdVviIaLgTI9eO50s42HYlrbF3RRCeY5/h4hemcGVx4l
Zq//hQiEi5ExEEiSv9WiFqELK8RHvgXHbJ2Cob2hj8DFas13+8vtxMbYWpcUJIJI
FcQ2HQYE/ASH4TeRvy25ZrLADCEIlq9U+3G7O0nkpiI1obrjInBcfVHJLLkjDkms
m9AEsE0UPTLF+sfZg5bkt2vES6ofAWytYCK0GlUXXCE/MOTOznQluy74CtA7Lvt3
UnHMvV1t13ePo0XmpfJh5K8nfOamr1E05eyIR7eOpNLXWwGRado3G6/mFWzhRs+E
+eqAYed2RCUt2ydwRjatJMETzJTVUpRLEYxlOLrtevUaEcrLuMMjxpX9dT2Y/nl0
ZkeFiCMVDO+ANRIWKlXxNr5YtBJX+U6uxF5uNwb3iXUBIFJredlVc4MEFoptZDnX
Tpmtiu4lszL5ooisLIw9gC2UwdJNMO0LL009kY6v8rQ8l12gx9fklfWR9Hc+yMXg
2TTGlezukdjgUr2rTZdlz99odDNsDfdQAZPk9dGVLaTU0p5Mk7RlZqSdfQ1K9hOr
g11cxKXf21jCFVmhcByr6QhKhB2ilkqKC7aqgoV56w3YnYdQ64DQOAgGR5+0BF4w
Lmfpi8wTDqDnBpqtjKqlNXxYyVaXqUseKWWDOG8DJx+0dr9XZstFtBEqXGDGokVA
0rhfjVcgpB41NYCRviKOpb1qrqXg+A89pXwcw+ZdoicpYjV2IfPAEaeLSodr3lQd
22QC2sSbZzbPAYQPJ+EOX4AHRU9GqVSRnACGSWMFNZXvEBvjDc5C5aIFgEUZevYj
KyvoCu2MjfJgMEMuBNSH/YVvJsdn5T3YMC9qdl7Q4HHc2Mw4z+F5OGPmbQ8qslXu
omGNEVVpb8ZiE2Kt1gp3R1KiVDhIIzo7cOYwO5vZ04OlTxK03Ap9Zhga5LNLjFPy
IV1pBuyfyIPK+Wi3bihgHeuHbBwh335ci8VIYWSaKhND/yrfYnNVMN840kAcd48S
0bovywUU2HIBCuui7Y/uB/uF0dZBWrK8LAR3asnVjS+0rPldkAkL2923sPgRwuYv
VhR23he4CVX7FH0ICVMUbjKfKxpDUxgJ776lhDPtb2C0vUnqJdyCY84i4hADvYiE
bDwYfZ2qfSEj/jql2ltM8NX/uFNNws1GgVw95kOlidXmhXT6xWrVVrFvVmlPLGKB
sPjetUUY+ugEuiHMojA27+WcVbEIClCEbL1ug0B1KqY8IkBlNQLfaBGXV7aqa9kU
3HXWfuVCwgVdveLu2lHPuJrv/q0wM4wUyHOWrcKlM2ykiKP552M22k4GglBW+IRT
txprnp4FJaPjP3q8cFxTiwBCz/ASvzae8i64lttwdB8cRcCU3YwKoFL+f6J+wz+c
HL51dymJeqp6k2bPrfVdvRPcvJD1meSNJcQDLiqPpbR/9uvkvxPswqorVwLCGeeK
GHYqCAVL8jnmrSf2KVaOTcnBKY4+Fljb+4nprh8d7Jm68yvpBYWsJP1mXz2v7qqk
YxRFKMCri/uo4cofm5SKFdGn864Xf22kFXVrRHIAk+R/PmeGlL5Y/wp/1lFhby8i
ugzm5wweUDKuzwhfIwusqNq5n9ZwdQJeqYaAtXX9n8VExDgVbS/yPJLo0g4L+8CT
j8wrJZLGNpFTk2ABXSZAZeMwoPD1YpXUvvVxrTuHchKH3KadwhkrVtCHlA09/XDP
IzGf4JkL6OKis09KqiqaDlO8yazx9zdYZP5LI1nMEg9NMzt2ypngEkkG/MYrcNJC
sdCdfCH5+HEnuKYIv4275pfnfXlPM0dai03S5LBywEVukhnsplorEnfTLYhoqA3k
pYwLJepXsKz/u/ZpKzq3aNbJTIFICUatjtZiLgG/azwsUFsAHvSEHsYLM8cu6OlF
/nFCn7oFJKd4n61dMNO2mYh1r40HWlKurEb+fCpwvpKUvYnWJxcUkfYGxVXzk3Nf
tUQVzD9QLquNN13FwmdWDingjW1Wi1GZoTV8kxq7Xb66faHEGVDUCuZS8nqzCeHY
IChXqor6GgSp0KohZmxmOIOapktrjwnRPezdxbWpSsUjqn20Eq5H8TcRDBBg9e05
r+0n1kKMVydl6YeXlaAi+bgKe8sI2fzENHJwEO6LibyWADUkhfGYxB0iKQnriOJQ
/iIbk9qLYM+5B/47r58seppYFcJkVogGHly+BHzxF1fIPOWkdC7JhDzpy9KGPVuP
gxMw7H3YmYhunolibX9LWmcTvLV/kINBiDPHXOcgK/1ou+C/MTZbdXpWKqN0Pko4
sNBPDurjrSjPGM1Sa8zSnRjHce4bg9ESNJ0INAd1vtHBrGxvNKmD7uieGrqBocKb
wZ6eeDx9Xc82s+bnop+Qs+HfU7dLVqG4Oa3fD51VPYIESw1t45YrvZvsO49Eo2Sc
ESeKqmZmNYG9RC6wzvWdhe7JT18znk6WhgsZ3SG4kEiWi2NoEhJL40xYnZbSL37u
7X5dI35r1maJBCH7oxmzfWIDmrdylCMJT/AyDYx698ovWn1iSbvpDzeO+UK7zGal
v8wK/39L6vb82P8LwtFHCh/l/nXMBDPz/22kCa5JfQiC2Q+vQ9WAmkP9iuvEfq20
sBDQNHu+CiQaIIy4NGz7OXUVn/eisWLsqWi3W4veejP9GD1ieCPOAnC03dCffMBF
VTKdsj9KHS+PdaOv2r2xN33qQ5XKnZJu5k/XVPpSjEqRUCiK0KtsPac2kWLdUrCB
6qbUdPOtoad1XLPaWoBEkshHXGA560dL+0gyhkawMJRGG9BEXCrr8eqFUi+KiLHJ
VTdLdY9+lbRJA+uaKRhzNBbEfOQVPxE33LkJwL23teJa03tx8WbZYTOPAP3Bn+Nu
VFVzp2VcycjWfHNE/61N/pIbhbGhi/Kb29BKOWSJQhE7p8iLhXk1UgEk+NzOgeom
ZtjA01h3V61/dQkzNXikv6CNW0j3wcjLaU36XhXFP3b1uD8z3DxfNJm71ND9f7fl
0c243hyZcy8B5V2AXJm8cTa+lWI+G426Syj7dK9s46yjbFgEEAubeM4TUmn9xE6I
iX4znsJ83TGAhJylkA5EC+tmCQtCQpAOgPutSFCF5WQ6kAn+aQW7VIs9AvO8I/tW
mmFZq9qZW8DK/2bjA4uHt6wZJxc3UBppN5E8wTHN4WrKAkIBNIlhwssMDzY/QY0R
w1erfIb3sX3C9t01FjrEZofSK8PizcRATC/GveyGzN4tSecsnFZqBTmNeUBj4Jr3
3cPNHoNSsGKfnjjlenncPADCCUfwyFFvZYnUNnTP/CrvLzOk6Ssjwp3GeGew1SEj
BzhgtctdmXlxNqhWJNqDSHeQuekShcVAgwq01Q18w/+f/wApEgopAhe+JAPPLbHc
O7a9j8iJnhBP5FX6SxR/AB19IyjiLExQeiBaj+kcKx3jzuTizgEJ6VM7pcs/HTtI
F99oGosvIurzyBOHUJeVrYpOno0clxWEbfimzY36izN/9KZvd5MjE6oxlqC+sklh
TofHMoWH8Tjq1a71pLBYj2pHtCIByujkYAzaiTM/a+5TI+VT0HudydlnCq9h28N5
Xg9sSRXagX6m8uc4k8+N1sa0aC+p/n+xV46xc7Hfv+t5IqT0atRRz3GR81QlHpbg
e915NtnK4o27ruh5H/vRGtmtRTnHYnZVm/dJvcPfBg3XNfkiLRCJuD5W8tPm5ASf
QBGg+9vcQp0F7KAH84QFiwgwTS47YNwiiZgthSo2Q6L6nXPe3YY8fnqyvjhAVmhr
ZT46wA+eIeJFUtKvueqX6/WiDo3rblFFArna7xik7l87XJC1Lycb7zvKvoJZ97o4
E4+sjmc9BPmn6dzRh47Gzr+nMvgsr0Z/xMZWg8Cr0G4YPydILVBJDiRbIvenrtqW
BDvwIZrIearmlrqL2UJ8zyuD7ropgRuwl5/CLnH2DQs3kdahwPeuMvn1LrE2Hxqi
9H5njHpX1BZ95owd7X8f0u7Y+yGIeTiu17XjYpWZDCxUzkbLw8wLq4woQE78brWt
5ZhHlbdv/+OCi5EHqIzGEKj0R+F6EOJdvhHWX3/Pi9oJjQuQhGZWP/EKvCIQSuPy
Ud+Q9Ov4INm1VM1wGvgZORxr3Pite5I2tR3lNFBzhrrkizMxzH06QwUn3MjbFY71
LzSaw3IQZsjUr14YMqg/6M1DlOFwaE5GwecV3G7X6IYPKZn3wO3C0IIs9syw6qE0
6Wi4nZz1z3GP6uDuKmTq2283Tc1o7guycRY5qtLCISY3n6EGm3DsMmjaJE6x6KB4
qnCTWxP4HZ+g6Fl7EwYPMo6y3yuBnAsg3F/JpT+HGbi/2V03o4uWxNmbJEGN1Uyq
iEm0L2Sdtir9qXR4Azgm9MOuKR/UQW+0PLHdvZhA0Xtshr5m751zJDaAa+BCoHRE
hCgoFjigmOeOAjaKpqQfsE6XbaNRiL27AFLb02YRedd4+IfCNY0ock8qGwaPj85c
S9ldnzk/uNoQLTN8UCK5bN9Y/mswONu67CmyqMhjBFjjVpYcPEYrU7hA30O7blAf
yozCykTo1mk3pKHeYriMSv5CiqmLGOe8U3gUCUgREiwHm5ZvISkay100yQJt1xJ2
43ei73BQk8DJbqCJ4KXcZdlfqo+hd1vOcCGPv/QO6wqQ7vS+lnoO0g8zOhO0TGuV
rllv1vhDPbh3yPlh+Wb8Dxp8XgVvDWuR7bWGXoFzJwd2GEff2sw0uUcaLHAfNPN4
nZFmx+iCK//8QAF3a0ZQkFDjTPo5H4UW+a16BgKKNiJaydyqo0tTppC8f38jCTG9
Qg7edKy8USuUhlBr2K47LuiDO46CzNdL3eV+86xbCOogCDyyyjNKTb7iLRO13gKK
Ex4iUSwUHYw3xeY4zl0Yh0qG2I4IagktDrsBIs33ZleRydwxrhgEESAXxjc28xrX
S26IfZJLeQfDg6CRzb3rOaMfvcIsmXh5LeTwjEOgPVGyqzXS4ddmcOik+0MGltfZ
DuzW82zRA8FN/aopG6LpiMTTp1MSIjbEmLZVQHsI3A5N4XT2//kWTCfExaA5uxQN
1BVhHSNFSayvx0IEc9tA20USapX6csefjIIcMVfWR3J5JXhR8OqFpGAMlJtj97yb
nqQXSwfx+e/vwOj95axyxohH+a1UySxONLyI7heggqrwxxA+oC/fDVTbjiFhSvxy
GRMwoOd8PaXciy/Sp6lk1OKxOFD00ntMioXrD22r011K52bJ+4BEiaEI/jCvB1Or
LvAQEO6QtmnPsWlvF/0eTXqSIIBXPYqRhaY2dR9Bt+zGGhF561J6rjYogOAo07C1
lMgmSL5KZFkyejVWDqe+FaOA802lt+KPA1+VYjzNlgPOus/UZO8a1oQqaLHqWC4M
qxKI3+DdXnO7FBQf0RaeHsbIOQtX9iTWU4RskRPQ0TSlSCDK5e8ekDLIIcI3e4kq
f7KLyMn9Vm4Wdx3sDlhWolc3dBXkykeEwjOEn4WiZP91pCv8z3XA1TwvveRiCrG+
ELWMf8AKYYmFoXhGXKSONSWJrUTFKeMot5wiu3/qE8JTs2BjJwfISZ33SXHyoqol
TUh2ZGPNoZxMxla3+XtFlJ+qtSbxajtKjE+XCXgSKuus72UmriB02lOi/JpTdFmv
SfIfnP17lruuDGcJjONQfOfIbZeJbJxKQHaxIS97QANFY//yXDmWe7luLkDVM7qT
3OCdrnifTUbW8eiW7NHnbwZuKEs6xp86wA/l/n4x7z2b1/EGNMNcWdF2iq6Sn9QZ
w9rH8+VZLZ7reryDfIrATTwTdQUBNNViASXD4dYMMHR6bf7aIi8E3igKezwar5hx
mzeuxizo0DeY3QIshA1tLzOeGH9E20An10nFlhZH717DrMO6aJsqjfKcWJDlk9Kj
ZSE/ZgTuaC/4YQvbGG/SH1PFhzQv+8fMw0LaOaez7k2VgXccK47xfi/mO/jQImqv
WLETeOQzVgqqnrKWJ8+ahaWLZKXKp8x32BaSAcNB2KCMGC9RCLJ0w90XlnzBllJV
30OFrNqzKxs3oFkO0l5JfvjwkWCS1TOFSMnK0qeQvKhoXBde6BzybcRuyBwwecSy
BdRKQsxPkhQT5By5F/1ZQHTNeirnnHFLc3qfypWHhrnN0svGcvIvY0+KFeDntYS6
WxkF9ru5V30mfLJ7FctFcqPIrnZCsu2I5BfgT7hUyvtUA1kRbgPJJhyYvZP1TobH
bpSCj32+pyJrIrh+MLaew0Mm9hZfZJmPj+z3bp3FivPZ9OTGsGFDirpvizskpYyy
IcU2fjP1t7CpW8fXA820GWidNjcb7CzN6dyaTKqGhUbMnzYYoxEgk8xrfaS8gQDU
aegvuX3cNjnQ/bnJ5w0WvehipA12bJ7IpV+qiA7we6CNSi9vayeu9G9IN40EDsmn
K7hW3uljQRBkyxECJlhIip/Ta6o3FrL6RQgCrIK2MIXDDVXUYaxIhxemD6N2LdUS
vjsDNIzwO7LHFDaCX9bzVRJU1kuKHcsFy2CcmagUcOljQZSxauzS7CbBRO0RmUYc
1wLCUl618LHFAhi0Cq1WPcOUikhuf+7as8WFaePbFzJVz9li5U8gHNJzD5LdtIFG
5UsTOX522JGxOi50UH7ay8+JOlYYoXZzNJkFoVOREdydNZ8AZRLb44d4o7//1vUY
E6m1EEUqtEx/1u/FXyb5RFml5mwW+Ip9eaCsfnDkibhJzpqh/NKoGaX59yVSdWk+
z2E2/X+cdZ4ywZ3bPJxMvy6aAGjACpZMQAlPzRdTp8L6hJt8QwGpbwV14yK5TgEG
9vSsmz3JZ9RN7UD8Xhpigjd3GVAwQxn/LnbBE7LyF+Y9yKGO3+/DiE+9Yxk5bLJ1
DaFizj32lR1eDqS9OvZyotGHrAr8UOCKFfd8lCzCWBlInmSq56N+aSSIGJaNayx9
XLg0WdBb1sTG5Vn1S7Xq4b5+VfmlR+YPvPJc6V7ObkUVvUMp4401/4Nr4phB7q90
Q4SIIW5N4R5gwFiNJW3b5n3FVuhQY9pQLySccgDEs0oTbVMS62D5wke2PUz3pvn4
BhFERoj/0URhgmRScDd3claduDKPdouBU1t31n7l+v/rI/dNEtVUIQbNEnPgEUr0
LG1XcKqjCUIhhEDjCGabtwpgMjbY57X8KFlqpwB3br+7x67LZZqjoprfl80LKSCH
JgxKvY5wrJzvmHoe4byqng7K7FZzeV2cAkHWFhyIxbRJnKGxSqBlpE4x6XKKGkWT
EWtHkCEy/OYpYA4x472fG0HBi9e8iRlu6D2jtf3/9+1st0QXg0Hn7oTDh4Nn0Q+H
PhP+9ZUjo2cBnyIhyvYYylrKpsLGGIN6TuuHJezo7agciuZZpmdSKONspXyyk6Oc
irKuklt5z+2b082N7Q8oTRE70r1OllvI6iELgTmjpVw4EyA4M8fWpM/UCwomjmCP
pInTNYr/ycc4rSde/deLhTNmWboriBJ+fo5pvSRh6wKUXUlChn/7qYKFIGINfqyJ
5Ia8dihjfM9Zmu3SBqz79AhS4NubGrTuK+yaPfbiTwqvlqwaUUmqj6bP8jDsDNSz
aJJfcnwRBjzikqG22JyuUFxnoYFCkw0hhhziz70qU3Jq2lHYmtFLcphksZfDOEPj
NwxiUIU/wAcUtaMgMAN+Gz5cD74qFku4j17p+68TMKReTY8jA73p1ZzE2ybSVQQM
8kzYC+spsPp2dTxVZSbHC3BC+KNAgu4jASPRo565HcAiIDARwdlEJmNWxYWMv//Z
Pwk0IGYHZqu0MfLW7GKojNgbCUBYOjcEQHniJFFJd7lJUqJow81nT8h7amX1GzGU
Cq0M+uFCqmNblpd287Qltgeqo2hgfTTp1G+nCkCnIk1UdAPd7Z32BeF5RwCb5yG0
o/Kd2fBiNb10JKGlNXl6NT7Vg3amprddD+8vLQwwaUZ7pZOrNezEVdlSN6Ic45pa
c1ZWl9MatoKvuLWLqa68GKcjIA4CaJtbh9gowNtxwlwF82/809nyqklBIZLKuFY0
gFZYafCPykJWT8HihAlK3gVlppXp6/K/oo988FG8SQDm/kFBKL7hDv1TZHedasdn
Al+UJBLsPQXWpnmR5OKk/iIjlAi05QDIpnXLk1Xszej2At+eEa5PdtyhtV2LXcg+
w861EnHNBEU8rCHHBvxH4wvIvA2F5JzR+1ks37tn8WH66z9Rm9WO3EAupVILO2vi
0btLTwzBZJGBM8fFXRWUOooLPCxJIm6pg1v9p40wXgFjeHR/qt4I1qCCUi+vKPV4
6zjttCo4XT6YA5gKgDguGplFNwmrdjtJv8zCGqSZSZ2gw2ujgZsdzcR6HL3fid5A
Xk5JXBg3AApMqGbsSYLEcxo77BG2zR3t3hW6KnwFuh4NvLYb4PJd7LyJRJTo1P2Y
eUm02jKCQdooYJJ55Q5a+Ri0l/33aBwTByDat+qVz0U4jWRu1henKZrDOcclWfEM
nh12wjPozJVPn7fwTvif2GHx/Tujh9OFzTuWii16AsbV83qQcY6YpgL1LTxETTbo
Qes9YxEjOrfSqG3KK46nH3ERiU4Ka970wlJERW2BepYON8T3EvjEJgMcI/j9UnDD
w6xkdtX0cI1tTaKxeuamUbCGuVEY60JAkkpIQKcnqXUFixM0HenrEOKzdZDpQI6y
1KdhjsKf3q1Y/CF0LIo8TXPYER2zKnEoVi5AtUmxHUyxTzpryHW2j25Peds48lQw
CLR1nf6xAXZrUtPDieu7jgmjnSMqZK8KnalpHtrMKKAf0Il7vedy26toBdrxhVz6
ICMgOaybmGBNued+z3US+xWU/jl3ydVhZ5G+DOVefUgu70d7pkHiU5T2H/tyfJE1
5ykayp4QDDcNbWi0s5Up3k3fsi5/N+hqe51Ud+XVdSZ5jG7AocqTTdjnzE+x6DlK
W3+SSLJIwV9k7xokggi90vAL1Q1bJJ75SPPlPxQjN9m+pAN+b1UkQ2594p9aKWmu
xGcS9RHfdDrw+SVhOIPaHZxUm1tqV4djD2Y+Yj148DLoyaT9Qgj0XkM2yU6mCE5Q
NF071NNyLBxf8WQF4bqw3Ymqd2TMs7YpvL5Rt7Q9guK2NfLx46akTe3jfV7lceNk
05ga7FBvBf1/Akr9CD5U858kMpySgFRV+jSBCf1K01vbmPUieF99G2fiWChSlJ77
oyi6Bn02Z38qx+6sBVR6QPsPR0uoyNnhtZ/19VvKa8ihd7Z8v0KMBXHJTM8j4n8H
m/OQQaLAdgXicvPHs+44KebJkkOVY3x5p4oibusQZuyk8SPl7DlbWdU7nB5GJZRL
qZRxIK5j31YxRqAK2ifY9SHbqtuZhldX9FMB3/RkeQPzxY+v1D+/o27yVXyCM71r
UXSfKmmuil4+1COZCM2J+/n2XZV1f48MFolez2cYBW+Cnqqxtl4WFrrMwDgOsGCs
1gqTujJBIn2eECoItqBI7+S8wtaZxFeYDCv4bRTEVymjsLNS6cnaYWVdLBZid1Kl
Be749+xOHBvLIpuolgmjUxUc9lrYz5Jwa/qi2G7qyjb7gP2n5Vme9rHKAxBnLDVr
EYP2JZc7mjp8FDl5XuGCgHWG3fC8hZM9nFFCycUaKAaRWqZP9bxweNCakfWaXc1Z
5qB/jbjrrpHPlkNkkOB/H88MnBgdLuxEAmDNqx1sPb2cpJmIdQUakhWfIt0Ti2I5
DrhJgW1HAC0tLvHLlUUomDCwzD3GFQnPilLMflmyuBQFUl/MIYrr9idSoEXGgLnT
eWUOXp/vnrA9D78fpYZ0VrEcW8RJoViY7cr8jNz5hYxxYcfLeDo+lgju3+bpnLBf
VKtNSKUG5lmq2HejjDDapmsG1ytiFruMqpypzb1d9WlyNKtWB+RzwxZr9Sr47tU/
Nb6ug5UqSq7JoNMXRkKIbNFrA7B4+Qqpcpq5Y6O1nl7lPjZq5loP81YzswfdtEVX
XO1uSd7/CioQlNbSYBGIEYHWvxdNgWje+TVcIh1WPY1ILQVJ2bSdesfZPWw201tS
PceGhQy3cb4DlxH+RiHuV1c9TU6bb0CQYgWAxBm/H+RkZx/7HUv0/yesmsxRucKC
8grUpG2WY5/JxhByNrRSZM/OppGyULEayScomi+SVVIMuspddy+vgZv9B7bOsYYf
F3ORamAlREWDCNsAV3w2Iuw1w0EWGnpwC+etrXvRmb9FFzixCCU7WW3FtM2qm3m2
SdM88Yh8uacgssEIFv/p6/zsCbwooqq6GGXskVDhzcvSVRPoUjUZ/Vx+rtzVitmB
Kb2Jzf7CnWRoANsfbUWjcpr5F99Xn1XAjkeIXpSx1slOI+45e67XpG/P7bPL/bgi
wahkWser7VV0JD+VqBogHFdrzHEnSEgYr601gwgRaJseCJmOL35qGTzMEulPlzS/
WiB/rlGxaucGqDm1wN4iNs7+khNHaO6MSuLowEr6ssYsF456wdjYPO7v/NtVhST0
7ozIB8K7G6VPWzuNinyCspwc77w111tmudG0XDNepUNhhxEALPhigZXo+uBGI+rn
/0ivcjpN8g8E0jbrMswzvUdp9QKqp7O+ClFAEv/Cxu39yRzn/llIwbaEUHrUCONK
p2ZYRZMTWrD04kb08SNQRgz6OSAuCGEZRrauYjh6NX8QwnYwxezfycXrwFaADy6B
xRvVzDTA8/oxwIjk6GqGVFBcJAnN0AM2GEWS5mcIJyl4C/LPsBYQzOu+L7DZeErS
2nT6lv3BKEz6JeezEqqK4BkMJx9K5wT3f+urpngS6RHjug2NAJAXCpwS3hqF1y5U
i3q2nJRrO3R4L1CLj7f+eJV0xORBfFCstNdPl5W7jWInhjTa77Sr3C0bc1vv+ZMR
mjif1mEoU2ZtL0+ZsbTu5+YeyYUlHZANs6qxXpmVSKJFXswqztxnDSmVKuTmc+BV
LjfArjE3UhTBXjBgw48RkZGvZOQhJODqr7qUfDXFve9CiMGRqyJO5pgHuSlzs/u8
JqRCyYlVqbyGzPSEJdMPBxwbLxcoN7Jm/xMxnJrK+Kc43PIl6VleUbTviS2U18lt
POjQiJ9NutXd7s4N04w9JAsJx/PJTyjoUnwk5Du/fsrEBXgd5UBzdpcA2P5AxQC9
5N6YSLPqj8XIFBrYcC6eIGeaJaVnB5BSVmLlkNfWbv2LK/W2IMz7Qzk2HRqUL2UG
WjLv8EcOS9iW2OU9BIf2yJaV8DtQJc3mlC4y8bHyg7Li0rx3IeQWE/bZ8kADtgTX
7P01fohI9P4o6+W5CF2bsdB0YUkM6PUQ82ysc8TzBCbLJIpQ/tO+1Dr34h1DTH8z
YMGCVnTDmoF4miyYkZ+kyZfNqXO+cpAd1YUreiTHnjpToew6qmPKu/ILjpfBm2GU
bK7hpvwWQdZCNb0j4dCazddBjf9ui1h1jdmkhxLNplK2bjOJfVaE2cX5gdfjiZYr
n/OZiGKEoCOq0tWJFc0NtaUJX29f9UmDQs3g0USvcrnipsDEQ5iuA/WS7xbhXaZU
gcl/CJUCi6UDq7tNahlzIIphWqDCAa8Yn9kT1S7GJ89jdRLrwhuTRSDhGO5FbpO7
t8oerlyjAhBXobo13wxw3/D1hO8HREJevNH2nfjxASW7AbtjT4Sk/sdISjtboJ2D
bHJeKoSE0sD192XYTo8VAio/eelSAAW3ga73R0Ou2Xn4BnxGqTJ622+genSbR9zs
BONtydhjsIPI782nXnu8fmmkgACXUszSP/HPPqTWXyj34Zhm65DpMIrN8WnVN9hZ
mSDpNUV0i5YTYPq0Y6AlmADH3OtLuCKUr3uW24GTbJYMOCLsdAL9kJx41Sk3Dq/A
phFtoFx/lBaYzXQf9BK43z+dc6nWcXztMAK/L/lJDkdU4EKDILPnmch7sp+2A3l0
buE2DyrN6wUHXOEPqanyfv6CFaDY8M9x65JP6k+GcKIHzUCTIfqV5co479QtrLZR
wVs34v1x9yXZ00WxDq3+msY4pI8mcvZcDMyzmMTP/5mKwrzQc4+c43ViwTtWTSFV
A78ZGWDD5bOMM2jkMfYwGnSGnYHZaK25MRP4Gnh9WpzStyr3cBMjQowaWroCXHuS
8TLVn86uYEbyRkzU/apvTZDNOK2DlaYnx5gSh3gmLyQ/pJh4mfq/ntGFnclD56Hd
a3D3HEwBghtTSJagqKFvOrF0SyS7r4TK5eaHqItWA3pFWZnDTpw/FoRaf22InTrx
ZECjI204OggngLMAS/iqx8hOYD3kh3tLS6CPcq/Ui0kzQCQaD4EKtCzZYRYeny0r
qWCCcxC2l7QaYvAZJPzBC9TtmvjbrNaXJIgsQG4ZsBAqUTZUUGAxHUBRABicDX6l
9Rgw+WqbGLqczBx6qwmjCAm+evZrGbwBJQFQ9ncsDfkv7iEyj7kFRJYHXqUA/QiC
u13XX1nTFjvL5eKTQYDIx8vuQaVgA6/xeK+37jpjL+zs/MKyBAOeIyP36BFd23el
QNokOMhOHGMcLaJh5OPb6dNOzEGKXqxUklxywk7cyKOspHC2tHry7Nxa+nQtgJR7
icnlIC8D2NHKdtb53GqJkncrBwYMRtUrim3E0Gbx4d/rAEsfIekunjLC9gStPyQ7
OmKbMgky6SafHpoRo34wyIlSYwQpRjIlmjXbhi2h0lsjpmvT2FFzkrga92hTGOCc
CdtvoxG53J+pW3K7BAaeXH0Ezm2hB62MnAxA25oUlxND2c8/NjS0JkaL8ZRLCP+F
opuo9VPnJ3M1nxB3W1UrRPx7yLYP/MnBpnyKkssSwnRhEH4+g1yNLPcVYUkkmuBv
qUZ9RiaMZM4yWQ2e8B6/oCHA7u2CPqD+VuGkAqAFupJsJTZUk1QyRi0TWaHbfSqD
Us1Wuc0ZNvnEGGRjrLuEGD79zBr6zQm0b3fM+GKIP3T8daOZuju8+ID4YsoHj/JW
YLnvw91yIXjwFOwjiXiQ5PPtZ4GTa/za5qzVfLs9/tR3sR+j1b+KPHC3P6Kino9y
xdl4KbSmod6EP/7uE0KZQDg3jkPef6J75tlaikn9QqXAcXimUBuFAmBR0FQkRmR/
wjvLXJEEdo/lToMCNiygl9KGjo51c19tuQ2Ek4i428hFxPNJrl0tHJGreHF9rTbK
t4NHY0ymTMRzLdYC4vRSnjlXLK+qoTdeGpKVdGQQn6KJjFTs7b1KSq6F2Oh+U3dl
7EdBUN9hTVOzMYOlv6sWx+SNYR6Qus16WJK5kqboMbI9V747Y6r1ZJ8hXSzOoFjo
pEVL558Y+dvxpMHnwVhBS8kL/6Qqe43zZuKPWdBkOgYA37I/yx7o3NBoYaO7JY36
vTChWvidT7RyuYyZv/LIJtMn+LlP4S9ulDIu03WQVJUFJ9aSPJmExS9yIy1dj0ZF
MDeWd/De8daiHiZn5LP/4YF0/Ah5xB1Pe7Oh+zcgV+8vxE5um6LNthAhgvuBHqai
zn6qB+8d4+qk3CdtFmeJznANrCBl94pZBI0fWMW0OHPOOdr8hDl4CfsmbsszVHXB
uw4MpaMi1KnFoBRjGRyL1dNIbaI9zWpZMpL6aHmHdsRGgjYXaZ2QVLHbCPOL9x6k
AvQUQ38tfcTlmW/WFyZ/wPlWujSpgYcMCkPsdbzd9/9NnnGbvNMzAcMvdnO+BvPD
HfjmYTsGeVnWZ4RKLF7kTS01WB8ioVZmcIQFxsvZzPBg8noGysId81mdtzdilyod
XN3HAIqflQ/5abIEgb4LTBI6Aq2sor3aDIlKN2Rs4di02LxQZpaXPdaLeB7m8yMF
qg2uAXqtUcEAlyNtu/bBI3Yzr84kUI+s4PxUZgTGoiaFFKlfbBEcO+v1VANKwdJ9
hWVjVcFyRxsfzRdSbCIvnb03q/N4TJ+ryQqOttfhANC1IczZQqGghhD50OyDURVe
wJFKqldnKa514lrO4kjqWzPK5FuSHUL2KmDKPXz/tQkehmFfXqG04YG87nfjyf5n
U6nWVJzKcRhEFhCQY7+2ilrPLZRlkFhNzTEfUscn76GUOh37zspvkNdbnsLH4M/x
4PvTCaV2a/6uxe37eedBQFSa3ELADv2Ln5a/WTEbPAkYpx1CI5WnspNp6EPYdzet
jShzGfAPNccGww1fviWuiuLsMBRA3AN89knK+ymRADMZR3s0Vqs5nJLudP1ZbPjG
8ruDC48sjHK1YtHKeT3yXVCGAAVN8oZqP5rWg5fYQsZ/m40EKnbvEBCnzz2IlLyy
sm7xd/H8ckj5WOH8dixJT0DZFRGVmEb/we+mciWBolteTbUTfJub9tvgHXxU9Si5
UUjty4gxDKAG4cl/RwCCtzd0h0eEr/y1eUHPkL0UiunbkiKQYFwq7W5Qqj0Wbh9K
CPOwWb7C+sTmkmhFYMfLRnd0w/kf9pUOQvtQTDUbqlI1HJbJPmz9j4MGDvTlgcrd
KeWVC38/EN1WvHROFCD2encdmEfJtXLqCKOITsuGFDVEFgiJgbu31z0W3Ue9ZbAb
X5blEK06KJ4VFhEYlgjlmaqlzgZju1deaCjRQM5ZxX0jLWmNzH/pKcpDjT/ZurqB
6M0/rdAFPe7erdfgR6fJC2TrElWTywA60TazvLBoTPJYHwLVoUgP5EnHQo/TdZ7t
fCq/kM9In2ShZ/wXn0h6Xrb7zGkxX9LqmrGIeiwS+IF7kobWoqba294z6eNpcC5t
UWWSpJZftEN15JgTdsugqcG8NwQgT3FetNrKvC7aLhNya9DbHO+lcD+d1+cYRcIB
wfEMIO3L9KGQh8nTATe2J9mNuFzJKqwa11c2RBG+Fool9eK0nFM5+dR6mO+9LZF8
0BZQjSVvDi/oVTWa1pmgfhI9ON30eI7ivQVEXd/6nzNexXaTHCpCWOnXW+lZCRxl
8fq+oKYDyr50v/CGFBtXCBTw1xnhhVxK74PwSo4bWlaLGaNKUzAmGhBb5lCExbXl
q52WC1Wtla1ml+xDDs7FHRC41AeJflkRKutbHM0+Ye1n7QnsnZZGKUuUAzfGJcDp
4YjVOVGDtzzgDW6WY9ozCl3bS3hTqU7ySi/5ZjgRHbvK7Bjfhieu3j1rwGAZjC6D
ui2E5dao6p3V5TTpb2nxRogdeZIkZIt9DKttU/2qDKw3jGG1UrscmRAI8AO3tq4W
YlS8yJy61cBFgSV5FurpOxZSw191TrH6y/6CLdAeoVpeiz9WyoVXMzOVD6ZTYkad
a7p7uz1VH3y7xi+T2Pg1yugWu0y0a31ZHYUcwgTrbXnOS88dUBAYrzqTdS6550wp
WWxHiUWIYoCIsToK6lJ5gi5kI4i1JxiT6poOdfIpOW7VEijY3qpNe0F4jrRWlCvf
7dLSKLUcHkyuYcF6Ilv6kzomiUnBM/7e1v/1+7p0nj1yInlNxHJTZb36WDc/urNh
atowNgogfJWiYhkgZEyvJ/milK7ra2kT+jHSTky+c7cooodGkWpanjMIeT/HYw5s
p2pURrbF82B8y8Q53YxpO4aSbddOHiUYp9J4YlTEynF1Y2ZnDLhrzpSX33EHNhZP
CgWZ+3PjF3Ag/dVwJkmkBRlF4J/va7mYFU0a0ZoHbcSrIYF1WgCetq7og1/SeXf7
BfWrx+i8491RryXWcvaQpqB8NwrZd6IqZ4LKLn4n7LOlBosd4U+jfvjlkR2ns+FA
zsZvzelPxurdPCBioo2M9YHiHgZXzsnDOBNVDzg81xvrUcLIzAb+JmMzSElaQFjj
8wHQ+apJpyTNCG/VVBOs2LZhlmbfWj6kuF3y+QXsb2rii3qp7L/m48qnCLcqOorx
EfIf5A4frO4AgNdCYq667AZhqc/wyY6KZQ1TiJ3bK1ZfvbLgvOTCn4dKxhlI1jSy
0WDRoXRLsEtjaTh/GBMmXhrsRMkuPVCzuJjLuL0RXyHJvD649Z1vROg7uqNl7E18
XAlYe1A9AUBgTDRJ+8fX7IBr09372jGCA2MSIe4FmXsbVwAGs6saQDwvgWOB1X9N
w4W+hN6lj9JyClAw2VRhqqWAtvyjRUh4uC6Rbis+M7c722KSe2gFRMlMM92bZoXO
aLoMFPPc1u0aCAuwGpyreb2pUZfaK5/1QbaZiAH8pOGAC6qhmbqAX3KNY6GrgRkK
RU064h242Gz85N+TeOFI5syLPk+/gAoaIMZ6lIpepR6zwzgaGcT7zC2/Eep4hrml
MFvaj/06SZgZBmaZAzYDZac9kNKoKd4rklndOKCkz3Z2AOgJPWRX9ByB7C5TZICl
l9kxGph5np8P3AlOXhcuCo+pQynlrST18bkAu5YxfnDBLhH36g1sPnB61lgAaSvb
zR5Enh3+xjbHGQQaHl8iHRMmmt9NPxJrMcDcmMFBWlY8JL7Gtf5hFSZikYAsrVrC
rBXzsMR7W0UiR9p/kGfRmQtUJSRCyXGY4Dmd1U5hD1P7QiYik4h0VEwtFFC1Tg+G
PUk/pqGj5Gs+iQZcwpB4FW2iwJOyuQxyw8PzcD2mWgfb2Znz/+D7me8leazjkVl6
P9PKmQG+wNIvlj1PJOvGc68PTrU09SDppWFp0IPrnwVcVNBykMyF6ubZvXt66Iun
hzAXt386Wkp1cOWZdQrcm4X6et4c4ZKhgLvbWqDD5WK+eqA1Pb8UWXMlC5zd9MNZ
NwPnjI7BGBCa6kJyKHJW9/5U2nkWosyhgnPx3CFlGfe9U0X/dxRzzJu3+OOIZGg0
3qXxPzm0KaxuMv6ycCaG1TgLgx3xQCSk+c78vxVBNM1DbeD5otT5E7M5DilL+iUG
kosLqAFkxK4qx7ioYS3Njh7E0jNzDzjKNseELJxG2NxpG6xhaFilCTXZ7hUkBxyh
aU2hG9aXabtN5SqwjxM+Yc8IijSSB5oHEUaR27TGExt1eP4hVTxoN1ICMQK+MQwj
Bgp+Yd1eU+B3pitpZFCUn/kvVKsw81RabLSTMJeqYaKJpuDSJ9UW1bxyIMOr3FAA
Yy1LX7ifgX0aFlGorW8fKEQ1kaPtpXOIBGHYxq/b6kQdK9P8i+/q0sOcfIwVamvE
LfwySSLlyNM32/B3CdgaUNuhIRTkXru0H+RTHNdYwefS/MPNWkjEKSj2kh6YWFSX
C5iRIZvjsqCJe+m3RMvUDX4dGbVQCSSTjaFVMV0GIk2GEOaJ26DW9fHSQ4PK4iJT
kgMnCdn2lY0C50ogX/VYm2y7jK9dkzF4IJDzZ3OuB3ofx8Ka1IFNjGmF8SJTSL1/
bhoAut3P4UgVIB/xBggpLGqlWjDjCoGnyuskpxDLDsep785uVpnVMmQ1OyrGyBYo
XG53Q9X8RIzdWF6P5fEQEQfIn0ZFeVJkvrbxem/TdA4N8rstsg7kpuyISD4OQf7V
piWz388A8gF9Bwz+mnkVT4fLkFGifh2uGzyU+9HI7sDdt01jDdgYAoswME8OHX0z
pQg0e/NONki3WTVmbK5WPUSTx38bQfnZNShpZ2C5vq1+gwfExMKNqNw455A6jUVW
rh0xkfMJSj1Jm3JUfYCKO3IpA9Cb/CPTvBXIPe2Vd4g0YNWiuiZSrz3pKImFLo97
u5GtF7C385hZnyVB1Uo14+qUtO576uUhNJ2BNfX+k29F3XqajY0Tt38flapagqYk
C4rkICxN7xUKu+EU83knlCJJNwwE5n3KKDsgP7ZHCyxGO9HW4ForYvQer4vfZPCe
PgPkepXC4GOKzDX9hg48HxhqAm6Di5HPaOWNWDiC8rZL1HtYkgjCJSK61VMDLFQQ
uV3PG5tSZRj/AXCfr1waNGOKus5vS9SXkYN/OVBg5t022ZRkJ8TImDLSo+dC1dNj
byOjveizJNcCiO/T2IzPXbRKfadWQA5bv6ANCUdHGSLN+7lFO2JEI46rgcslmxuB
OhLBCjMH2h9483VXUwZHw4Z9vPO19Nexm4gfXLPEjsQrssq6mvBarrnJ1uBdJ+E/
uz8aegSL92n/AvW19xAJzOyUdNqhxPi2qXT5z+T7a7vvyKqbyA5EBH5XnTsJoWbo
6gEQo4z/8eE/RzhX2tKNnXoE6rDrwKl9tliz4hEJUtE4lmCXbfPxbF3HGE/gEibf
aWZ4mv/2EPbS1eyrSypipPcXEUXp69003zXut4XSrawpgK3ZlisScMS+iyktFTGp
t87Wu+Ktl/GWGCvZlZ0Fp5IbfDiu5lefkJPYg6OZmxyEMetRvfxeUrGD+lA2aU4e
XnQvo3cC5PUBD9vVSTqnzVj5eblSC6E5keSnT94POzjJFE9h1oVUVDbC3JVq4q1/
/fuqY2lWSbHkKVg/pUgQ8+P88QLebPzPMYXwOIIiJtS6BC3ZCS2rGzYaUI1BL/Ev
6fdP5ZjWRqThqzuPW7q1lXRHCX423u2ekS+tpFCwB0OtZMLpOKt61M6FtenhQ81k
9MxPIq57qPcqBBb/IMFz75dyK6CLa3b3RiTfgHt5CUVdLYik1cLO5UYpnGocel1U
g37d/cO6o2b5ksNCYp3EG9BfEiDZx3SHCYbw4WiujZyZtZUXbRfH/9zcZERdC2VC
JMsBVC7lP3pXfOLwqNzhcuKo91K2tCLHN1A9sFz7RwDzG2nq5TrxmQhiCEJ6OMjd
47VFUnvKD86cRKoL4evUSPS3j6X/nO2wzFIV/WySTg9+UEoB91jQ6qlPPHDURrUk
ER26PZN2IRRsJC1DyIfc3tsoRjN5IM3By8kwCdYuVLL8YlBnSdA+SOy8YsPV54ka
OsGPqepWSC7ydyZRAkv4v+l5niBlPGw/ia4NB6xTpiMhmzmRRKwFjWvYERbpK62I
6+ambxIO8Xyq4hUi7xhE6c65rxQpCQrqt/prYU9fuadTyEw+L3YsrLl4Fo7XiT0s
iW4H4W9noU+dD5Fq8bwhY1b7gTnQXcZrj43DSKAgI+MR2ZkS7bUYY9vV6hwqFDpq
QLLIEbTwEVmfHYQV7W8RjP66aKKeijKXYRty+JDmXrVG0dZIm0heWqQ3Rtm2xPgY
3F21qyxk+QD5Af6c5svaQyoadudXMLRDfpVlspYbJ5W7YTF1Y1ro4shRjOJf7tet
Tx9pNytIRbjjGV0HXh+OO+IhksFRZdigXvqfXmnaQ25N39irsb+PlDA/XJY88s/8
CdgDxowK/VJZFLmvXkzOtQvbdiuC8ysYKRi1SX3lsZNZjYQBixi+1cxRyJiAJimd
cJKVYfR/spejfXWA9c/8lnE5Ia6Aen3BXmteTJTGb4lCkOUWplfMs3K4eYuxQVBI
pRyIfzwVEHP2E2Oh/A2Gfe6MBtJxdmySOTyr2ZFUck65DcnEtpBvR2qmxnCUBRWm
hts2ROik3yKvurRzDNTOTvStmD3DBu9z/5HVuLIlYrXezGPdP+gJnZ8vLRpIIofy
x1kLp1Gkm5Jg5ex3JYI5znBWMQehSfEcO/WuWA17bWty8Z5ZGl4bvrmDlbCEARiz
aaYUGtYy1jZVGxppLftnl5lVTC5uOtOo5L8fY1t+qn14e5GwWiCpQakmPTby0veG
Z0dHToC9w6hkFvLLTZ+4DDd/1Bco0X+06xdpgTWTIW98cGszC6Vu/TA3ntooYA0t
mVKCK+m4WX/M3GgRDGaAT62ksl7Md5AssKklj24ZYPNAOzCoa+2HdIrJTuy7fXOK
b1sPB7cn3bI+VzISSwmAm0eSW0c3FCe8uXJjho0BMfMC+gSjViLBXRwrX5Jjj0TS
KihiYpfYRSvg5jQUA7kH8WwLKZwaovL0rrpC18DN8M0lf/XCaMeD1RQmmU4f4oJH
7eKKDsvL0/gx3XN9qT52pysZAUkTjNGtZYVlVU5qcpRKp1XbUXH+uJtfboUoh+CY
9lrEzveMqLjzTzxPDtcx49jNF5LgVminKVsz05jrw9R0SvfBRKmFK6V6z9xMdeGI
uh+/pQSpLbp3ZKDsvcpxL37ozftz22PkeOVpXxPjErmoBQ7+i8xTQ9k1hTsYO9RL
3J5/pvcgisk5V74hYuyKCioM1LbWNXgqNla/Gojz3ZGUM8WLUqxAlSD4J1zuzLpw
DuRCrM6nW4uO8h3u++3cGnKhhHgVoHJGxo5A79K2Gjc2MHkTUmxrEZf6MNduXioY
8u0degSXd9Ozm7FTxaL0NRaUo5prgy3va5QOOp0EEghZERNG60txNOSmNpB25TdJ
1CvLh68pL0I2ZNa+h6lqR6GpFCHl0+c8yErmpok4y+J5Y+sD0HUDiEsPxNA8Qe96
8+kgXp418nCiC9sRVVcegWvPJWkhOuVRAu3KUIaDhAQ6gGyToCCKfH+hG5KFpq5Y
DEGPGNdFxieraG7Um/NvE0giIAwLVem9JsuZx3uqnbOK+70loT2RnlWone8519OY
Jz8nSKuXwsBRaKUjC7/lZaTNFFLG2fXUghfAQRrXBjYoOiD9RLiWUrfz7Jq13VY/
k6eFy10Lhwy29GNwTuKFYKF8phCMmRS3Kew5pV+f3i64J7KVwva9i/XPVT5jdlwh
MaL6DTKed6slS1ehrQAJS3YSEFwIMu4MAeBlLs8R+1ANE9CWsxSFoakpTS9lMCuo
VEBWZQZzn0xx8d2OYsW/Hi9B5nIgltrPTBgSQ6/KaCiuqZgBS4n2YVFqyuXzhgCE
tDm4r0n7fJc9zEcwcWYBQWrg4FblvVIR94WZ5+cNfDhnPKRHkYy5NFGbrEDkTerM
2mzpUXoksJ05/1cJMI8gADgbcQQIRHViB7N02Y5oufN1az7Jio5SgzMPvKTQ9teD
Vh9Vhc2WcPP47fEzp8x2xcR0CsF99Q0smSrQIp6+EBS4K1dCcrmnJlH6hhqUa8AG
0gNAzviKr97ezCNe5KNF0hBN/9DZlGgwE7zDX/WvuolK3fx+TN65Gw/oVl6eNS95
JnIOJHS25OFj/iTQvORUhHJws9lDGCNYYVTbGLAmZWwqO8wFRJZR5nZPfmMEcuVh
fkhvrjJCbDRemrjb1yJnVnV5ZEHsqXKR/IN9lW843GEiOELyLwA3CwEqSyfMJOBP
qDyEC9eJI7ad90vm0MZS3xCA1OOG8HgTTw29/j69zMSeM7xt25WYu348yrOcU/AC
N9MONSuIKsqAZJjK4bCx4hvxQe78dIzOwALNkxS1xM8EkJrJJRP4oY3f0tnE4anO
yYse2sK+ytJCMOKaXgJfV0uNlvILRgUhUK3lV8FwLPqF6XqRyt6ZlnAzr3Nsuu5r
GAx5m0TU/DUJHlijwdANCNImw00dnSabonb5fOXes7NDwOOFkd+2qR7DvlN1RFhN
7C/ENneP8EbkEWOPhIxiqVB6rMmTk5T7yh3hnGKQaLLFOKzo4TTAmp5uBLCbFJju
2uFcckz8TC2gWKz6BsB5AZervLy+i/TZTlRWcbbOoUmJGfF+nGTDLpZAjMiZ+7+Q
OFXcb37Sxw3Ra1BnQaApLjyW/NFi4yXkkuIW0XBdLoj8wYTgD61eL2jQ3z/mnDLa
MdpqrfT62gSKZ97ORT5Yox4+7qB6IzeTDnXPc9FbXhXzKn03u3mI35R78Wsqaw1o
wz0VUyzcy7OGkM7YsnbpNirl8JX+Ct3tEleTabesz5AY8uNTwZ6x1vtoJ9or008b
X+ePRIaQbYmdykjhQAAfhwwYC4s2QVI8DZDwvcmJmcOHj1vJZaZgQZfNuNy2F4Iu
qDjaNbkWFZY9ziVBACu+d3Aby5EA6C01MG1cLrZcam2GTAF1LbEUI5mRV6ELrxBx
90N/GlGuSmEhSKgqHHwx8dgRHVQRpgv1w1ePyYLtU5jYKNxcs/OIMqEhaHnr9w2Y
da/xdyYRPA+uPRwUdsiGMmqluEd9DCrnf+bQ97qD7bLdW4qd+X8ccbcOKsCDZ/l8
mszEbjGXUN5EbdTmkuNHuBPh/Az5sF5veGRIDyolhtIeEaW2rHmF5dvXcc6zqCQk
UcS0N/MFOXS+a4DYWezUtXqQZ9RNr+Su/OtmJITvIHqVZJDOvGCA69pkvJED8vQo
9LNN2yTiJ7TBWtSDc9q3jAu7uuuf60odYlkv6HFQ8H8PdvHun6LIzWqSZgsvpuZR
UtpE3O7fXNlJSa67hxMp/XFrgG7uOfpOKEgCOzMdhpdWnpEkAZ41e9vUbpV9TDin
u+aqJUuzpgKzrC57FVcrxlAB/vDyyLLg+drAW2mzkV/5AP03Q8zqBBQ3Dtfcjf7d
0o5bBS4FHdyOdiPeb+gdnTyNjRXcIGuh8sDl36BXS2JqCmpkcy9XG64ko38sFv/b
TpDbpcJ0N9OUDhScaDsTrMKL3QPSMzW2487AWEt2OsbW7NsPpV4O5U2SgDAVIO3r
O6Km6bdftrkKn9/CWxQiEtA53WR6SEQRYAwij8mmhOra4iyFxy2mayb7oZaRPMTM
c6Oorc9/zvLD+tUjx1JddNCp17zQsiVGw6lji/T0wIzg57ZnctPAmtopdPws30Le
U8GX3ViGIt0MuEUUWq6LSj9l0IF7Ci4UOuRb/O928bcCH5QHMXAuzWoLU8RE+inD
fuXOvARI+HMP5YGb+GJtHsFCJFEzB9h2bhRS9VVdXmVr5ig52aEZwzB+rQjH1dpj
mkiFLvYGh20SsMw21YcDtyVfv9oKJdehVZOnc+XiLLfQMsooSAWIYb9NMCkxFRBQ
yX6Y4fmZfRZcLz5hUTsPWxoexYEQSuc3LU5bIrkz1ZW+ihZqSWhPPigVwmrpfT4T
uvvKGahi/5SW/mNl4lKuJIJPoS0xCD4kQm1pPiSO23cEDOWWByrBGfvYLhVOCyYI
I7qffM6w51SiKc3Vkvtfe+9GgyqtkrXmHy5pYFezW05sCVLB2C8aPi6OoM6Sq3Vh
AC/VgmADgv0CTeCzBkZrReRndGB9ZtGbnWur0BkBhQV5iH5tEpiafFwRvHju8uZd
dSoZeH8MBsG8/kMmoffrSf2cyXOyQKUpWrjNznrshMMIKexl5VXXE6AMheFIyN6d
6+Pq8wze7QVPgPJP9wpxspifyPeEgdHO/SIaiod59jqxzbEoeNQPEb+IPhj/I0/m
KbZ2GtCfRAvBCkSzqi3VpgiD27COZCYwsMPxzYinRQT617fuq0kNkvhKIW6unz4q
fzmV8sgQLOBkA3Swl20n1VzoAlpm51K3jjUAMcg+c2I/a4/Wq4kRM6EVP33Z3xh9
oMn3qR891ciUcajPCLTdc8m6nH+az3hEAKmQTL5Awws/uehdm28h0jSb0mmFxtxR
bSdKfdSeTwnikz9642d+TgP42PMfkQKmt83r/euLZndBhwHWM65wQo3bZupxVmFT
+FoTVTC4cl9RvdkJstDM/Pa1HkLdCwOwWTFAdHMtISJPFu+7K+8T8l0f3+jlho9w
CRI06EZ+XKkS2JrZrKHVBn/z8DMeEi6A99Y0ecua+s+yvY2q0drVCyY+O033Fofb
z7VvYJRV7bJoHLr8FXoT+6dB7JKclRswpPUls/xkzxYm0F1TRNVvnuVxTT+pBSaI
RjWcZ/Q85NH+miCGCwhGrgqaLYVbVXYdjp270GrF0GbPDwaMQsnRfZU1s8X8Jfbo
hZaOFVINftX/O9y+5TiL/8efoEzQ9VVFQAaBXKrsNskCUjSEmE75FvEkS+8+07Fk
hRIadnntURnOIsXsZtpr8sJQlzEmCwDoAKttsoieDahECdDhZr/tJWJlH1S1tups
MZUqVv5jYF+pRieL0DhQNEypKDPm2I0Hb/YX7Rao5q+y2cIgLug16F6dhkMBEmXj
9zWqObFexC8Ok1BOwqYAkAGi9NzIOQ2ZsaYNwpbmNrBCtXUb2+J9VK+8uBtRuimB
7aF1kPE+vJ4dncIUn4r15KGw4Bt4cbGCRJHnZpASvlSF7KaSSCrFDmj/lIRF5rJl
fHbqp2BGgnnVVE3q+3o3lxBtJEPbRoi9vqD+gpXYds54+w///VbN/xw+6m7CIHzt
IyUCJNAbZzAwCTJntFZxWbV2fjsTjQBrc7YUofdUMlVPa3miYMxVZgUKaXoazPo3
mHWCamRBjSEcCJW4qnBKVWGGoTi0h2Z+6GQdJ78f/c0EjbgJhYC2Pb/nQS5do8Mu
FrHtcFkyT3zaveArZKsjL2GAngsmTW2bG1joSwHG6R4fgq/USh1l5u9+WmI6V0Lo
oUd1vu+YqjzAZPfqPAWbtNKGvnrnc0AOdjcCrFuYcO/Ut2cE841sbkB6dZwjiL5S
vTfNoLTXdkY+faBQnlm12NqvO+wFr+ENSzNNn+rvSI5rUNSdCvDDZoqIixWrDInZ
RjNmpyn7cSk7LGEc955LIKeYPb3mb2BQFA/WDs+YXpbDdw/ZtMVUz/ezPS+zciSa
3jx9LeUKrGeb2wyrpjm+iFh6AHkTnWMMsGqIKz8bUOk7VsgJjUV/XpzO/Pg7Dr4c
RhqsVsW2uxdiOAnBhrAgbc2Lphc+XP1KxaBZw+pWZNRU6I023Vqsw6hTeg9g9VEs
zRaAyHZ5xk2aR4asx5N42pRbttC16LOG5bK88OTdNKTroDStV8w9BISZmT5nQb8D
Y2gjDOy78ZpCA52PZj31tw60y7Vd+RL7YDL8kNj3EtQ8JQ48+9Ha8EMM4Nw211S+
r21AV+KH+LrzgAL1CQtR6QOetYvD9SvQzXqg0KhRsR6h6qCFLsZ5SsUGMG4M73M3
rD4G6rsXYnThV9iizzbySnzj2BP4uKDKeW1WvN9wXZER73ww8s/XZMuH3kOOyc5o
WZCuFTazfXVT3DGeZ3a7A+7MqX/883X/g3ef6eWsTtCZIvAGYsn9tSjZB0qdeWZ1
o5Jaz2YS5DvSUzvcG7ghCKdOnc2DO3xBG2F7chxPKE334BsXnyH4SkWSTpxRC+2e
YVG2hVcOlGyIFxCbnRnz+ewLgk+gC/gX+ISzgIBo648FrSHlVrbEgCfqE5Lmxnjs
0GbNzfKQXuAAYttEPXCca+jvl7ySyWFkvHUKvQFK1XB69JqKlhUko9O1H+BZRj0E
o275tmsnMdOgk+9taA+ZjUUJS48cDk/04V2A6xJiRBdWVGmnpewfrFkEhW8e0qVx
bRoY+LGgFh7s2dvgQfU6kT4hMMiTr0Tf1HJM7vpqS4sO++xPYkvaklxZRpKAwIkC
mjwo6R/sr5/xROGiNviG1gK+dY89Waz2qOhGZkuIMdY0Yl8N+2wueg7ZAyevmHC7
h5+JLyaRx0a4eC8lzOExq+rRDhHq0tmrbbFwiq6IRpdAPxyi6B4vWzxHe/gZY8vx
SRjCoTMnxse9JOSXwhBo5NkJZqX71Sv74JREZMMuX4tXvGlCyKdchTxbzMZRmhHE
DsJUJCDLljUOFxA7YH9BZZkx8gl/TWvqjGI5Ctp0/s/vV7/p8EbTsG3cYK4pLtu1
whQnOS2wYUnCd4AOWj4wtiv9ZU07a8esofQP3SIGT6zaPN05N+GXe0UH1SHASduw
5pm+yZjI1Nxes8KngThqDzG+kd51QsowQkminOUgGByTM9RyIRD6YJhzVkPgx4BD
t15ciKMiGctbqhfUK/Pua6jPu/NDL2pu4BTS045J49+znHfnbKuctdR6KbbeofZQ
D8/GvNyOYgAW7cdP/KVGSdsXvxnLobyDTEJtsxotCOsjCYJi72QFQRjjh1mDRq6B
1usdnhSM4yqewDClBvuM6TlgZOBaUyjy4K1Mz6uyDYtLQySUclFdrdYKgjcPTE/d
OtmhKu7Pvn7kxailadeeXeDwh9GLOzrrUFD0nIxc8mH3v2o55n9yKKIvuLpdwSDz
y1//VERHYmh5i7GF91rEKTA9cGwBQvjXOeeHxCMwgYpiHy31fxe8qjS7fqIy+dV1
Sj3loNFRRbsoeSNnLO3/Z7IuP3janLcGPT0ld6v/RP1H88N8vpwd/KJiWO094J7o
d7nPPjIQTwEpk9cT3BSSaIZnkFXZor3lRkWIM/2n/KNM7fZwE13exUtjuCdGoSJs
JCFDcgBJXpvv0vw50Y+2gfhIxuYfYM8Q3DUesmEzDpo85bI0dmI+v7i6TBrJ6U9g
rdUA8JS9c+8WZJIC5NT7IhbJ/1xzfsDn+2e/t0XAd7CBoL6jgMh9iWFUUSPm4tsR
Nlh2+fVAw/JR+JCZh8PauNpcq5bGEQIUAnoZLvFUVoB5aVFcG5jo3UsvOW4tqTWU
oclBfyk7TqJ/zDVmVmfGe2XHwf0/qBEidSJMCRXeTjks/n9370f8gfQXJvxk07WB
E56skoYSDh96oS8VLSEyrADsw8/uJMtOiPwWJtqzJzXhiQI6+015BowfXsnji76h
ubOlaBTYb3+Fr4rY5q3L1LxZwIGhqIGqBHwSzi3HDv2t3sHtz/OaiJ8em7pDPY38
X4g+kmC4wAP3g3CTdiEq9bQ0gR4NqiQ+zmYhdeP6SomAINkAtd9eCfbXeBh79VGm
xAS0jUN63MDDwP/diTyQpFGWCfL01thkuM8pfbwfyDyJuNr0aqbzw2IA0xrI4sDQ
6EIOXYNSYkTUmpcjBJJHnUq8DXhBt5S1fYW/evCXvgUa1RVP7QtzhsDJjwAbyPld
my80APHr7gaUobKESNF7CFy765qLTLqrDp6jPVoZXrlYihWktXhLv/e67wQI05hL
5IlJAV22jdTQLc/eXIu9JuYgo8WEunNzweK8t4BgvlPfOu/3YpYtr3XE+zMkHaAQ
8m3TjaIa8W9dlCWa8WSlR3Sn9xiRA0nKZI+fUtX7YGvr23FeLqa6dPiWNew2oH7u
nHPfdUdHJxWZaRiCyLBkF1N/hOsZqHkYwTWPTGiL6M8=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 26864 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aXtofNDQzja9NaCJV9U+TSZPT+mQJgRhpeTKbPOaCnky
F0sgbNeWLgrEOwp/YcnBCZ1QgHVpDx691gKem1NsWxCfTkmFLcmJKG0gIqtXWfLX
POUQCg0Zxbn6u+SsKXyCbapYSgbeZ817oBLxwBSIZpwxiW4kQ3KLn8xaeSwl9eor
kVXB8lKoV9u3hBAp70SK+IBTBiV8wL5aqLCXFvDPePt0Es1XzeT2g4AxyQRzdycl
jmmE1t3dWnrrsEOHKNSWAqZoegmpfoLkoml58/oU5ki8qvoln7re3ntoV27DFuW3
tPcoYKUfUIYDOUc0Heo7JdUPNfUYXJIYE1evbPc7oD1qbDpwF62BgEdjaitFjMuD
31DVMA9mv4G2AX3JZ1pnVfB8/LzgXPeDzMLJqGP0gHqeX1kB4fYCctSV7gILTsRm
fXbFFlFIgLeiCXctfeesZPCSr/29yKT2DnhtHoqIimSvNThuxpPu4jrgjVZAW6oi
Ebz4sMsBT1A574LkqL+qgDrjt0YY/n7XZt0B9SfTLgmEAzVKlIAGnyTCfzxoJ4u2
xYL71iUnMDnFJHzjGrxJrPJXT+p4zF1ZGCcWPVtE0NNUhJiFlgwUIsR+c3lCURnx
PotMTigTglUuQZKym1lSSD858qhkC6r2tPUyHKuScrc9roXq8UXPgZk9XaNdDhUC
opLoPk83gUTrXvLMm3J78fT9msgmsi6u1IZqgSUr49hxpDIenUlFo0wbhVerM2ij
odBkIW4D7uteoTP4EwTSdCmfLPSWZkQNggNjhQhj6KAG9Xl4x9Gq2Qw9aJ4X3SYY
tQjLve5tNNkYg3pgaCE7SzNBPVngeLD9qhHugSyv9PoLJaal4hxuKT9Sb7u7L86i
TRQ+4/i+W/8VFyM1uJFPZdusMLT4Apfvj9jOJ79a8XBMQ6fDnXO3qqFu7EEOBpp5
wENEqkgYQE8nMIZVbwss6QH2XYMWbFVXH+V/heqWYrk0cNPsWrQWQl6y6B37G//x
ygn1KiygP1hC8eTggOnEFFVe/1FCp6I6TVrLlu/URPGeehm9sKWpiSzQeficOGlK
ZmCGxeiz/iHu0NBLyCrD1KNls9SdhN+F0CdSvSEtXzlMt2OtlddUtkUf53ZsEuo6
WjIeDgjs/c/bbWf8E1PwFvuH8PUMsQwAH3JcJ+s0VXat2ceT4uYlxdHyk4qtiJpG
w/l9aBN/YePHXq92jTJ3JuPgA/9VlFwQ72bTgz29vixN9Kq6ukhYEGaaYgN0DAh5
/TrVOBYnHHPP1sTiuy92eVksS1QTJiSdLGjPEKrqkoRyzWhpqlQuklJn6Cy1Y6T/
8mLPgdH7pEvxVdoeF/SuScNdKNOfgVF/9CQkycNemwvliz6gJ+v2MWZF0BHLCo1Z
7PWTJ73cs6wIPbIe9KIyrMfe7ZAE4th4RNQaXLF8vwH7q7IX2HBSLzOKcyc7Z6B3
7Fqko7q7iyF3+BFQSHct3POXQdyJf10VI5ZWUOVECVY77i3EMu16n5SX/smIDN6z
rJeaYoBtysimErp8FNAYrZV+HTlwx9oeP/CZxWesKdancHqg2ankjJ/dYFyaI8hs
H/+swBuX4p8rtv1pM6Ic4nmPvsYJqTSz2U7SG6yWq0AbOoJ6Q30HHRQej00cJFM5
opjADdz0CCoZQ5rwBtowcrYdtxgjQKn6kPqnGTqMQxKv6kqI0Tc7I0XUuMBYG7rf
6OCb6W0Bxido4Svh/dEBbAnA2Cpne1Q6aeBGYj+tK4LafxaEdZ458XNIsBLK6dC1
js/6EUk168Ir4uh/R34K1sqCFaCKskMU5PNMuzKWq2x5rBO5UuhaSXFOfppYORz+
nYd4kwxx3wge0dXZnwYPTPXSVjFmU8owE+gmAyV1yPpqGySaxbRZMCzvDyf77Xu9
9nKNQ0W68sN9umGYgv1auDU2iVwE2CoD94NvTP6b/sV+azAmKS2n4a4HsFqnLyTM
e3AVUr2gEXipuNr40TKizB1W1Gi3/LePN44ajEOhKJh/Wyem/OKVaY9bYhzh9aie
15G1XvkHX44h+3hyoazJBnY2kRvg6C5Zg3w+iagLAzSp4sTD42aq9raySbRyCH97
RFJZBiZsizjZque8DFxLH2X3pYXFXjs57Pm6jSRrTzhapZP0J+MfgPrF6CR8ZlR/
wpZ9cLXDv/Jqh/SmgqCVFjYNSITlHXRTr2LXT0uKYrxDx+w6x7QJQsgn3ggTERzX
J78KuAUkADaPTr19LSy1SUtuByC7mlJpAaJMyuZ8UeLjtox3Vk4g4eTL4mYcWzaX
h0hyB+Dokw4keBpUcFRANET04CXDIFcz/52VtnxG4MIuJR6Dp1goB273yUzL1qIs
VbSyiHpLa3njKBDAOBXNZTA114B5ikmFpiDPbpNx9qb1kseaoqfnCkwSD3/vWU2p
j6gP8QhVlCiKlQcsjZZMfSyEzhMYhSpDOMv9T9aoiO/7WGFz4YENmdiWW1eKfdO7
MOO37CKscDcn5aYowuOXRuZaifEYCr2qwiswtBip+dq0SF2gtRveaYpIYhBdWL2/
zVrlsUmkhO4kY/7Bj4Rg97E+NUPQ9JdyYl8A014fAREzlLkN7UucRJ5FyWvOyj/N
x4wWC/MLhZ+yG/myBlnmFRZSId04Esa2J1C8gs7+GGt5kOVH+KF6j6P8RRR0xz1Y
DlV4oYxvd5pvcGbeP2QUHjVoybfOM1U6uCu6U+LfmRdPfnTlN6MHYfeISfOUV5j6
n1h240YZzjQwi9w+1V+Yh+M1XUXnQ3BH5hnaoqz683f1EH6goN2dyJNHFIdfxDG6
rGAsgKIMj6zPoLiASwqxbQDO2voO/7FcghsGwgkD01j6LKzhU0tWhLIYyRmthjXr
B/V80ccQlFOPQHt6ZB0DH9K9C2VFBNS/4o95xqTE8C6niNnHY46wnVAWPDzD0BpH
0BvI6evDYvKiL82RCbEay8wRoyiwM3AVEEdIMEZ1hawI/mEY3tiSP3FgI24kbc8r
KzevB1LBOH6qSCBeYWg5o10vJGTMPslZtRqMIWcYMlCd7iDm8LodZU9QR0qLI0z1
imVPfGGesv/j+yjbBjGVJBs9CCH5mhES1BrgTj9QvyQOb/yCDfzVcjEuWvz7nV8c
qPLzUrUD1RdWenGrpjchHgT+7FZ5tLODMMt5ilupykHHmDhQVGtMcgd8gmx5ZqO2
fOT4nWyBpbJqK+1F9xtuRf4WSimsaM3CpEJVAW1dcgKFvqR8D/heNqdczRyP7NTG
IEtcDGW7bhu1Kd1oY2DHRyoKxkNQ8ur3QlrdWUUryi89GJSa3htHeYIl4KqUkijf
98QCMMPX0Ffk6IHCbKL4BDdH7BmRK2tTNPIAZ5P/TOhRjpVEHaFMLWLxAKhJOi+s
h9738YiqdeZ7eHbJKsycmErQYsQYowWJ8UqXfTUh1VZlAjNVr6BDsbKNP6eruFl3
o+696oo/kg8G3ZS32YeCDYi61bDx28GRmDppQiZ+fQ3mav/DgeIE/5oHsiD6HZHv
1FaFMwTGhdiRRLDDR/v16aKDqA6FMbPVwEOWGRPNKGVzg3/NK/txrElH0WoJLhss
7+nTtyrJ+m+IoKWdCxuSTPxoJLW44Ou0SPKHyiFHwAdJWvPsElNM9E4+rZ83Bb43
rRUEj8hiHIQ6La+OYpflETXL0AgQdEsJucwaJX9XfsakMUiUYFCr5OSkBGnvWWR8
HLuK+/OeTsUOAOEmA9El1sxFqKF1hQc4H6oZaDUW8SDBVoADoIm5yXKkYogxTDIT
dQ/DPorCrk/WLjedIbDsYGStxn7bpiy01j7hmabZ2jhNsVVblOjllRpwiNy1XCSr
VVeQl09Ss5wuphMnre6N9zsbpAxXbxISnGdiO319cDC/5FXA/wLN96ozk0XCv5bz
i5RPo6+4Mev60NVTvonhHvH7JLc8xZbeoj4Vn77J7gqxHadMvUnAzl0/yj84guC1
k1MBC0cmawqBW4Aa4SsTzk8eXaXcDyz8PRkZY5F32rrlbmhDx6FpCWlpfmEPD9hX
BS1gojpKMThvcI+kCL4pDaRMo10fEmTIgPxmVcG5WaMcMKGL2nvbh5d/w/NM6aux
reLKjE/3rzm1gEN7BJ7rG0iqQiuL+UgYpmawssYC4nDiPjvxhFlBMUDvt1SQVsb9
NSuFqO3RntC3xgimJzMAig2oFwSlyYjUu0X5Apv0KsV0KijNDNehqC/wAOWDecLH
n+oFBrvPc+EHDT5NiUc1u5KtKZRLrNREYJ/N23Udcs62duRJgsr1AduA4He1khG2
EK0eeck/tg7diKlopNpaY7YcTA8MScY410ZTrfQnVM5qcuKqAhWzW8pE93C6F1gd
sLdHTYwqeGExaMHfugQjXKnTmjCIXV2d8+qNUujyUq7INrcU/88pUGjdz39BLoPZ
G7ysnZXjyDhyhyLVCtudLqKW+dTRdKT2c9vec1yACslHp84A8G5ppGWCtECbQPl+
IxmwlzAvN1g1SDKMIeuEPImr/3YZOTi+354MhuT36EBbifvlAjNCzAhhcWx+Kn40
PwWQfTr+IgasJZI4sEYXa9JEnbLoCAo7AwCMix+bhlxWt6j5UeEW/GV8pGCJ+fnq
584a1GRUQGypiqiLmSt7owWTOMImiXbbmGEfZ/SWHnCEScRYhN0+pBAUNc1KsI/k
PZDPzpBrdVFE4FV228kgaIiP1I9Ii+1GsplSp5NOFBonnzg9J3Jc8BRWP/2bqjej
W5hUiueggw+NOOmtWhJPTm4tZVhPaJ7GBTnucsGJBi7007K3Qmn+C6NQUsYtG6F8
M9HA8QW8t29MwIfRVG98Mpd0S0pwN2To+sQdL6H8XCjHvtaYkZgu5DnjUC1E7/oT
jiTx/boBRsiIAicjjCcujwGhUH8Rmhiki2+w1PIGyFBIeH+ayrrcdLZEuHDJh+LA
xEKS7cUivJfDAf9bMYJl1IdksK0OewexQGRD7WOd7iSxG4rpijNWgFX8PAb+z7LV
GJmsYpwKsWQTWTedQJfa3iDWtQ3U7tDIHTvFgM4I0rCzBiGVX86N37tdMnDL9oV3
OgXrqByTOUJJ1Y/YdV9/duXKmoAQcLNxbzD+nuj/B3GgZgZGppRmKdQT+kae1vD4
/1jNhia8ezROdSoF9Z49j4hBP3b++q0j2lGqu7Jg4gMU9hdkm0oxxCox3f8vQZIy
OmngmpCla5ifPthMsWSacEKElEwYPhZQzN4s1ubaE7+Fje91vOahi3AJxelWnzHw
9XnEBquJbWyznOXBLVSjRtPib6MiZpPBz7zFxxgaoqTnq2xen5hXEw8RIWl9+htk
RWHD96ejT6g4G9i5ZfdgrVgaN/0tLkDmHvaH4Dt3WY8dqKSTIIrLKBfRCCNUPnA0
T2jgE8UjvR7UhxwVzU595QlIE0Xo8N6Uu+WR1tbSsGhYL7n06Edbdm1det1SPwCD
U7m/BTwRE6FXqkvfTKvjJRGWgmNy9kpcHCs7ANmKVf/ASoU/5NCDAobHzzWiCfGq
T8kOFUF+PMQ7JrP6G1KjBcADBQaKSm7EkjNV0WSrlWc98m7qIqOSVvzolv5BL64H
3gEN+8/0jX9XFlqzLeaqYt+j3Ose6EdHx655mOF+7jfJZ+CL9szdaHkEqKNGWbkw
/NSJRG134+lWOEEc/txO7cxBBbdnFzbxuWgNEu5/S/zEQfO+6Mh2fTdAKZHlzKc8
WQfqoH2TbqXNpxQ47LuYCviqY/EF0G4KKGBTR3T4J+ug0c4uSg3kNX9MWg3rbjm6
NYlNhV74cyzs3YKJ/mH5/IcdCUkZWr79Tjcxv7EK2XTsPtI+3f932hpmYWeA/D1u
xJldWp0bDJvYqrjmlZD9OCVQg83JwZ/HF07Q74tyHrJLc3Ujw3mars/3VHWDasq3
m5t/Q0A64pbc1djdWPtbAXIASYPL6zc01DLJKRsswfJdcvHD0rKlLVrL0kSIubhp
B9S/FSpkTJyCwcIgUX5URvhaMCZ4HfhWHM6lXmWayXIv4IMqeKosZpPl9z7ZuiYw
OryD0VsvCZC4oVk/HufWyghQ7Qgmhs2M1Lgo5MjYJ+J7We4hXQbpZF7fY05XXU4k
+69bUvslNL+qBGsoWKaTQXfWiIluzIkDAVEB8EbkBqQednT2j1P3feEWYcriq8PH
m+ybXo27T0H9DViKFZP4611fWCemztn8yUA/aNy4kgQ+M2l6t8u2H3bfxAhCuQeG
CgvwFR3DkQmmwf4wjoQhikbLQzkQPx6k5mvX0RTGcwCOeIy7XOR1UpO76pvSdzBN
6bffEep9Ky0rJQ5SOzzT72/iHRClU7pR6HPcwul8Cmh3VgkCoFup3eAIzD+C82vC
kiU8ZrM8Rr5dB6UonVkNyN59Q5pbOR4EWZ04WJxK3NCkvzqh65a+sh4KbRcNOyjQ
Va0HwGxCSgIwcJK+nMx7XkDEmVgY9DL6KHcGuoj7c4iLS2vBZlhnTMnOVE5tnmIz
rLLmqE64neZzYxxZMA2w9zxFcELFyKMlnZ4l0qUqn9LDxdXXaQ8AxzHX93sgCm0a
fXwbC6QffPVGi9dgi/34D3erYcY0McH8XNkNQKS+0kMHQonZXs2oWZ21cj+UV1UT
C4Tjy6RrDjz1JXvJVaFis5tbVH7qyUnvoClYDDxOFwgagq6U5WYIbxF1N3FqbusJ
k1TjPnEO/mvqHJvuKdCoLJLypIbV/XL8s2S/TVmRdI2OzprFO3GMhMjRlUDUDTFw
hZTR/dmkKvnoPxMtG7dz0plbaxw3LFuHjG0ubcih0X0nx18L+9XQr5jL0sUfIwTi
d/rLAUQUfpjmEx3qnMZMSvQt3mGXf4VY5kGlQtDHCxbj+TKJSa6XF7z/5NWY8xFW
c2GkFEkFzxhc8E5aWajs18cqwnVUjR+YYUMO7YqcdCEg4zeBBoKcOlUKVEtow1ti
kNXUr1TMVVepa6xnYrKtkDDQj6UCVffIfAxCPyfOHmqqbtxyGkG9XbBQOqXmzABy
vHps+4Z1qlEpDibZrf9lYL3XTWpqQ9+Tb7mpX7fhDW6JdqBQdy1Lv/NFswNxvalJ
hXKgk0FQPax8968/eEa1vJF2dqNql1tfl8PN/7zIuaBXR3ExpviiRAMbWe0E5rRL
Sals0HV1biq7du/fpbDPzcxzIQj/v8oWqFPhKJK2fAT/fgl2Ad6hi7p5Bh5fAgjf
thouNEz50GGAt40R6VHcKFvAh0Ju1Ztawja9GdpQhuPCYz7D7XJkxhC4oRRBBK5R
6poLx4pOsBfI+PK7InuSTjmseFegBRt6xfGE8cSU9+u1PkPBs3ZuU/0dFLpSRTBd
TCqXrnD4useQrYmoU2Ynt1egWs0H5XJ2ZRXDLJ5splknAVO7bWz3tD2zDZDKLLsj
kId65Wgxcb5dI0rWTfS5ViL9eAxHhvNC5StQoxT7smwsy+o31iUatT7/WwagzSsv
LD791BtUO3VJa4SqaW6ZvIdAXIXeO/3QPQTKNuDokJjifM8tNYUK36nm5CBush3i
SC6iLw8/75FCHyZKAs0VukKVKi+faQRHSrIMMgQUwAwM4dpg5+E8d6fnhMyDP65s
qgZKrIvvSSic9r5dD0ja3psTAXyzzuNlIvFla2zBPS+yzyjbi2tSJRCEfjcRkA24
Ok+OpdOJw9vCiY+V3v3OcYwwLWvrbVV4z3AfKbqI6FUKtibzEPGezA/q6T6o5dbM
Xmockm43YjSXdpeUtHrRdcRDAVFteTnn79lQUl/C6jxqYSTRwmAp+UraPAKO/LlA
wXESzKRlm4FNgjMYjc8aBo6Y/cHRMLOSFQfcIOh6bYoNASQI7sKTSh1F1nOikBe+
s8uO7pd+rLzRZ4+wwhxt3Ronw9BeNeVkbiz1Pu2nxhqXPEiQx/7x/NsiUo0+W0v/
xcNO7BbIAOA8xOE5VdnuS8FAuDY54v5W5bnGxmPrEKPtQN2MdNy3Z0/chVSfAZ/7
G8FfdMJBUvrxvgoNwpHhb+sHpQ0mfhcM+QxMK+NkDsIoQwDNmYhrj/bZ99m0DvC3
Kc1bcUmsGUvvqAbYXfInzXY7SHwWvuiVwJq4McAkFjZdADAePZFR+4yQYY0vmPpd
1PSWmRBZUvQgDLloOn3rAHpYMzw7TApyuHSQMrADFVhxgTAnwZJDOyJQq39pA0xS
NuCDZ88u+C2Z1d/jLzGuNolaDw3+uUvfdoGW7yiVbNFcdnvLb9g3cyffqt5HQbsh
mjlU0IdjTKl3k6I2vJkY088dJMGt3sGc7cKKUV7zpEtw2yn17FCwSvntkTTatLRx
bV7tcRBPTq1vcIrbmo7b1Gwk4Lx5KCO/dBMRAXxS0aDARfUcZ3G+VJ8/ZrUpBuk8
EaFyfq4WKKuyQbnqCSnD/19J3SlFGtwJt6W2wQ/pXMoB0bSe3spFjUquUnh+NQve
2DItM7HIle7dgxpuaIgt1LtulMoU8pa7jTpqRzKytnLr41lMErYLRs2Y5flv7f/A
4SRLpYeIFI08nFMKXE+g4KJ86PEz2Aq2Z9c153KyVDBVl4yFyMqGfg5VOZOmEqxk
Vz0xgWDogkZ9b7EqBB4pJqMvNrYLihU9SACaa16DnU77B5HKoUqT5ae3CsY6vAn3
sxOkHfqG0S95U8UaqTPmhgul2oQ16mo1p4Sge37OCt7hQIwXPQGdYTO0O9q2BwDq
TcNxsmares2L0akYmfJsOfFyiLwpGQWG3Kcmn4jgT98pCPQyz2mWWIvjRaJRYCbu
3wYqvlNHMbg2tsdv5S7JQX72WZ1GhiyngAi4g0IRDkKKG+aPH1UG9jOuv0ahNSo5
yRdyDEAszgjskKFZMmy/a74/tLLtUUVHDT//J6PaXq6stXAyyZNipSj8bqVSzGjC
Pv18Q/9BjNlrk5c1Ni7NTK4y9/3h2d9ND6yAzAy5kXWinbE6UKfCqK1ZA5jNPiP4
56Itn3xKpWp97mysehB8H885zYDZsd+ni8n0XWk7rzt9TZRUB7zMQzsucbo0LpNM
4fgd7khi10HCVXskmb+AUSTnb16igU6Wl4tisVpBpMxoflExqd2SPUV1I5SUq83g
LFH/kYm9oH3LEAtzm1A4B75vkffdSlbMoyGFVcDxpJmkO8UBvCAW+IiIyfa4QBmB
G485Zil8XlLohwyFY8Sm+GiyNs5ZA8C/OAM+feiffbSypFW17TFATZPcNhFMyzML
woq6gU/y43rVsps7kLCPdDzpSw4ozD8S+4agDrSmpwvDg35ffyyVpMXBXA8EEI2G
ftfbhwkKpSpyzv0uz9t7iIcma9j1ubV/NEj+VGYUM3jXxtm/o/ILjGsqYE3UUP+x
2ogvi8fFgY6nIxG4Y8Z9Flr5KUA3HVNiCjndTAj5Qp+SOzMzfp9Ds6aYQZoaqcdj
ST4bXwGFWhQ8J2CITSb+nCIhfIpKDrbnS/RVz4/1xpstgqQjQygyvEyMmQ+xJB98
jjUKBLq5kQ4VMr9fN6QBNa90rFCMS7nYSBXt/cNz4qlWymYQzlktioiPCNMVIW71
0LXno5fSGlhdspAeKOS93Mx+N1xaZh/H8gvutrg63sk6QisiX8s9PzfsJJe1BM88
LWPiionxC3C+bHMCPgEz9xaf0w3d73pGBZK4ZAZn0eFpAnsQ8fhPxA9iXZNigtqY
arJC3pWZb5zTXk2w2ukdL+NpJ3yYIlL8ioZGmhcbj1+6EoHBi5MErAaqw1P/mrPq
xsolLgOR5fqdnKsBYVK+1TZHQagX6/hMUG0LECxKxcS1rOE63hVaGjPfaUQjxHAF
e+7d/V0n/R1sQvDCeoYofymRWwZ8l/ar9t9c5FM7tQvuG49qiunuNy9LHL40eJHl
KVyLvAhCcnuIAjUb5Ppyl6A2dtXExsszJ8DSG2JUdDl/+1URrK+XPUJmlVrpGruG
8kDr5ifDAMmmfXu+bCXJrImW14V2ZLOJUrbmttpeNVuDRkCHlZUqvq6OOjzMeaxV
a4Pbumh6HzxwFFjdGF+VL0BastKqEpozRE4YpOVAnRx7z+w4EL/uqldoUyfRXRFv
Z5bWFUOxmBGDAJ2w7L/xNqWVxvPDY6zpYo5qpCgUBTy6q3yYDuFF/7spX5K47iic
AEzCUPynkPn39zVkAxVxj/wwKpqLkON9L1QDnH5P5LZe1suO3LHiy1VZqaRHH3aD
WuuBMEMsR+HPWGVD7Zx5z/+/U0v/nkP1/6VvF9tb0cxr9tNxWUmx/pm2NPjF5yTy
JyyKIBcbHrmKOt+usHF01oxBjSUiEpvFjLspvkdhNn+TyD4G7U02JM2LihNL/LCa
xETXeJDP7OHNMB4ch6DlvCC5P5WX+Ku0Qeiq4O5RvXRITeM4ogJ3NW5dt23gJoId
h/SQa2nhM4MFhgSJCqkR2ELnibj4FcnpVCdedE3bgFNx9EnIwp+oMcDFX8ad0Wzs
T8GaFEdgcWk33SxaRnQYkSQVla8+UB/a0D0eXGALa30xMPXZkz9c+/KtQQnYdVs+
99id4LnCpxqS0R6nvBye2pC5Zg+O/7Y9oDcBw3VE9s1a+2/bfEWO75Fe+gehKZ88
DR481Qqn84XrplKl/B0aZqK2cOI2HMFaIrxLeBHQglLbo2dGYor0RyftKc710tBO
m6HFGkc9pqbIkAqHo/NJ16z4Fogv5nxtgWEX3n95yGxrNpQQmHjxGQ/fDr8N+jWt
IRT/gSsIQLYT7iEoxI4B7FgNbVgZL4g29KWYGLO8qlazvnsZjWtZub3i5TT3VJH5
z1h1Hefh/5C9yhMYpzpBT77zH8JM10GqUe5zb+NxO2536Q7JtoffaamXlc8GzgSn
JNKoPMEKvME6Z06ZqHU9Z96ZWzWg6ziQBxyBC8cWDsooA5o8+hQASUaZXbQrfbGU
Toefd5WauvgVrewIDqCctAAPSaIt5P8udTYUqqpVSnXl8jfNyOP/reVej8YthcH9
Qif1YKHLA2hqHLCj+5LEow2+2SlaEcWzu60XJcIm2qEbmhjolugafAlpDIKumnED
iXQ+Ov67trprelFFIh6AbxPa9r6znzFrwdXMbcriC2ERZwYIsXRgPgtZJuHEY498
pJiCLTlatADNWnscT3vT3ka8jp58BpgwbctXuUXvPSfMhctZ6R7wi4A7t/aHZahO
OeoEI9rKZTL1MB479HowbHsZLuVoNHMwafDOu4bmlbzCI9HDXAcUW0DUiOgXOd/F
OU6RNDunrd22h/PX31OFt6o3jmnDgkudBT5IzA6cfYOsx96h+ngAkEMaO6LdDbSr
lXkLfwMRgZkGT55gtPlbziytZkGFRpuKlon9UlpEGua9kYvQuMLutgRqBKfJ9WKW
ILKXIHoIdVDNwDMlQIrgZmBOYYlL/dvUL5uBKlpHz1aQ1MKF1q8VAlrOptXYREW5
ZzPGVO6al+FLP70S4flI8rDIf/5JFtTBd7IHDHCoqCDNIvspHNTEZ2MxuEq5hCOq
3b+PAUST+NSxfCYrOOml9CfFrzGcy8FyImrzcq8AotqKtMJJER0xH6DJq2eZ0Pap
n0fFHPBWpR/37zAFkuwZoZds54Ss+XBxcHHDQxjCjpPSNO/0yf7tvQoh+nthNfdX
nZ0QFQhq02qRZ1lUhK9jZkaZfgZwZXd2E8oEr560Bbaihlx9GiJQKsDT0Bhofiod
H2WKW9/ouaVR9pNxPOWYH95LiwKCrxZU+2ja8O0wdUBQJf+0Y/gU3TaeGrcrS6/Z
I1HmPtYdXKKn4zc/TxBA7OFd6qHmHO7e98nXYCLkQzJT7ZII4KIc9hHq58PYgzqm
upAjmd0qOGD+mD4+HFVjmx1YXXuB/3p0UUDgbJD3sVqN9f8acaYJ07fN0c4ugPNw
KIdxMlwTDocxtD4KiBhZAmTv9bS1+5PcMH5bQ/k2DjAkCp7l1XNwJ0V5W5OeXEfM
gxuc0q6iImQF1qGTFYATvbR+rt0U3LeM/tZXsrATRbKj9n95mG3tD7ALKeGQeARV
VZJPxaJOnq4eE1N4/D105sNhil32c8VNxKPULbU8lp79deD7gDNHZTHqWF/jnXFF
L5UEiGoD9a6v03vxrr5KjPC8sHU+pVF5xDlBezgsknBITAyUmi6iv1L4xUKV/PuO
BjxAC+dvaNCpSRhN6TSr6eDBEdF7qxBiY7EKBe9DN5cvZzwTby+iWxTC1vK3qCQy
BWgvboBY+q9bQ+3ckc9zOZmZ3D6ZVn913edEi7NUlbv+N/et3F7Nn1TaaFBiNZWu
jk3tMmT2VtXSZbV39JSjfmiG28Ig9LejMqNRqFOpu9ckJSdla/sFduyaM3rIUecj
kL4pd1C+8TXcpMupfjj7P92UT/1pr9Nu4L0xE/EJLk0c3uh0Zf9/j+ou822aork0
sp8lSs1D2S5G/X+5RKUAmhZsZff/4MU4zwpBBGRPsV0xCFghqtf6gNmTQQVDnOv7
wmerpkyqI6DNOaMgbCfZHNYjm8RTPuyB3fUVB08HFm8BzpS6cEBeeI7OKYw3t2eR
5fbDece8AzP1PRRi/o+ZH0uNLu7QlOvBhZEWnS2JIxuf4respuAnOpxhbk1aViJB
ucMiIvgk8UjVExyUSqK23vKG+Uujt4XGSrv5ZWhkHWX7DjZRE0AHPohu9Ywvgvxk
njplfs1nkJCEeMDV+aB+AnLhhjugVvx4rVMx+Cv3ZpjVTYAdCk7wH00R1ufFQR6C
PF+/jt9GrXy8nwlOzFac1pgzZSuX+Rqun+DDW6tE5rTGgbz9pKtgmeP0HMeoBb4h
lGMgFpVL8gxrliwx9TyNu5gPxxQg2WrmXvvuGYLqWuqtPUfdvjuCbSlCRIuPDdyr
vH8tyiJGgR21xG6VmBHJ9Jx5Ub7yyeR/rzL8YfbVhGrWsdRfU3Tw06PrDtK/qPML
+0FBDURXi7A1b7sbKkWFHpyL632F2PbAPUw0IKY+RaLPs+CqjBzjM+b9IZCCgVjc
LuzpA0mL9w+vBCyVUq7hrH9fCO8l0/wTrH4SYjljmhGJkRjqH84YnaJ/j8NySrYK
j6BbH8WEtsGPOpx4AqFOcGKbhLzqQcCHEHIONHfYNIrgy2Zjzlzb1PsREoD5HCm+
Br6LAlcWGMXErdSDp0GH37ia/c+jovz+wzJj+Vu1U8f6x91f6hngsiFQHsfIPpZu
rhTKFCPZ3GFwF8189F+wPQ77dWhzeDGgei5Mc0bvLOztqNPcYnFFwnhGDiuQwb4D
mgIFDNWPXGCGLx1p30VuLfBTvG9AnYzzqEmIBwgbz73y8C6NeZQ3fU6RCPLaDsc6
0Divj8Od8z92HZuVBiNfY1kiQSNShj0kKxpzdcHyApLtFEKXdGFBzO2Pqk1yttmO
ltLITRrgv6IqlvwLEVJK5kkOL69Qx9W3wsCovpQ3OcR4wg3Y55lFGzp5KuxNqJmi
tC9M7u8q8MHvZjZprc88nuB7dBVjEcRYzsS2U/PCUPfVvBxUEU1JcnhmHHqMPpVn
zUnDRnxuIE0RONtNV5Csjnvjdy9cD2F9YvXTjzbE/5dceZFpMbsmb3/0fTn3ll1s
2jbJ23+SJPl7ws085y8tKMTcXD3Bm2gBS/r1ZOKnTgY8XNLl1CMzUv8u+IFKrRPa
l21AEN4X7BIthQEHw8KRtRrJvU9OAEgV7Qa5sV2N6Hf02Dhus9QmkqWgl6xe5i+V
8cSZAj4qpoNBryHvj282TbYdaaMLb0/CyHdUkTzw0QP6j5t3YdBWjTmdP5Vw73b8
73OewZelbamHcvf4j5vAim1HXVBLpdv69KGaKibYSmvGqCEkc6QZrKfEu9J0J2NJ
EFBeN+EZ721wfW1yCh15zmN/vDs8H59fI0vvu72NOv0YeidaTssUKoPbPoTPS/UM
LHPPwk1q0MKxmP8PZe4Np1XFgYGtba+JP4tGeaIHlcbQ3ku69q97RBnSZ2SExfgJ
oXFqxkvtNITSwS6Uc8Z8PLdMcxUcIfEi86k8EKXyeA4WQ3aeKeCF5KrFku54Y1oM
tH24cQarcj5pB1AS80nQMriuxHUNem8fH1FSrvkEaVbA3l/LUXoz+vkFRoR61WRK
rEyUxmpBUYyQfp6H0GV9jeXjfMZRVANJiHrMFxRVgLerYyCXX7Xr+ArR1nYRwp83
h3fz9SYfwR4S/2KfVxWGTGmNa0n2iH7DPUQpAP6sjXtv/ibfIOEGP8klLI3pNRDQ
Dp8790tqkQwQdnqtwYnODty/XQg0U1KUUzZg3NYNkGQ7WmR4HQCsxAuniIGxOETg
UaT24nLaWj/5xnf4kiSPZD6LKvXiOexrj7CrRqH3tkVeiYBfllq2DV3MJc11gILs
FG5yD1na2Va/MXUw4isqbctHQwfEJNMoKscuhpDmWhd7BfBEFuj8vaUmJ2I2N+3g
Eb5OYaI8iApMUAEPzAAxJAMxWxQDVQhwQC/3nvscv/BeZ46n4+2M7DmCiG8PxEhN
bQM8jZ7STv/d0Y/6LIxZ6SYsPggpzHzyRm1BiUietpvxbSFiKBroobBYfzKDfwIO
8mU2Q2ZMc+LOs6EBpGlReN5C2MPwQTnXSAWW55Uoph/5EhDM/v5viZsPZuNpQeco
GD7EVx06lhqYcgQNGB97WfsSmBNSUWRf30aAGRxPXOvjzb+Qymt49oF53MXq2VuX
yM/RGplbCkcK3XvRxfC4U1732asuEBtJV+td/0sKTilZ6GsOL/+711d+XDE0eAvR
8Q+hhVQDQHXbxsn4jiHNpw4weX9Qb9xp7yJyE+k6lf49OxC6Ro6PYA9Y90tgBeZH
wgrLeCqdpj/UwEc9U0Gl12shd3eZ5FiiA925feBHLxxFeGKLqsUq1m5ybnZ9b2H5
87ZGeNKpbnmVZ/1Or16nWt7Hj28a4bxJwBoSQGAR5EgEAVsppAZbiI/U3AEr8ZkI
GLVPVPQrDDS0X17KiqCUaNbClalfwsMoSfU1cG6zO1IZkm29C0mcGJwR+FQkDa54
bF8mv9L4PQ6ZgC6XzQaUTrTttSNN06Q2Q13y7S7erTVERi0aM3G92lJNht0RpgNw
RrnCrPjM8MybCmxPMdfhe15g6k0ncUTSN8MUfU9olScXXWdG1GHTa/GUojaw9Guw
gmOAYfMe5RTqaK8HiuCSrXA53Oy3qYomQ6iyHrgAvVwy5nHXTbEx+nXd7jcZCjqj
aWge1SKReGbbkmriE6+L4Rl07Q9lnjB3YMJl4WLyS35xpshJjkIqmROzOK/vx07q
xHjLPiU6N1FVEmEv40+MMS19MjzkaYNZr4N6kw1YOZDJ0pba4B+1uQoACMwfCQwF
UR0e50BZOSTjvcF2hUrGGbDPQUO7z3HJliyKqenJ8METamSZbCakI4E55r7jsHFt
hdg8LLmHx3UuZD1uPhWy7KGA7BVBzafdP0WOYBeK5GDtPAZGfjJtajYWu+P3WYyI
pyyVYEW6B4+hEbSEhV1ubNw4+YQGU8h/3b8BZxAhu7rBJEMWJWc9u0f3ermVbfY0
95Pzs3OZbFJHpm+QlHIt4sfdma/rEH9uBaZG4504VQlefPQAINbJD3NgFUYy875B
Fl5W5qW12mu3aqTo/Y1IdFk2NuEf1rvcPQ9DI8N9WntsSiCHfpOjEp2YXHZEa4PA
5UeNMG5dgPxih3Dbp4M0C0x2FumnjezOmkchf8KUcN1IAI7Bdi8790u11KqDtayP
IEH5stfDNmt0MMfLxMCMXo4aKOP8xYcPb5K3/qUEfkUp40CsKHrz4PaCOZ/1eyvt
13q+i6OYNsJI7E7HaZbAv8c2UxmMwyBC7ESGTNx3CYvNsEP5lVv20VmlGe7DUsn1
n8wpyteajI32Nj49BSn1qUNIg1LNmX1hkhGN+W+KdTICtRSEvfvJdQ4rbBKsG5xG
aiGmChglNskX78dliWYyj1DTQ7xW8mBURKK7vwIp78aOamrCSmXsxAR9bg/5LfTd
+B9BbsJHuv7ZiOEx3UBelecP7QYXI6xhVBjRyX/gBx2MsIkXX7jcQcHbwNxT9pZ3
qGIC9dMzwdZ2u51npx8yPKJaAFCkzQaJh37D5B491Te1Qdxl7mTrlBb7DC9lrB+O
qz9bIVRuRQDOHAhDMU3ZiczV3QALUDmMP4QcyVvLxtbSG3RoK8uMhT3Q26mAMIYv
fg21DHPTcew7b8Bq19qZD1KFZyEREMKb5jkCyQko6RFRR+EmhM44BAtJ28O+r/ZQ
72su2qCylldecwJcibIvPavwGYWjmkW7/sp6l1A6ghtLmfiI/VhVBHTZW7xVssci
zYnW3tNJYS6c56TaKcJSy5jfxeKpld9BL2zDSA/MnctfIKKKU65ZjMjXcJsAJvKC
jqeHtfXhyMROjz4iNv6u5wUIXXzsodagBu43+0hw/pifZnh9mZn+CEggn6deCmgq
E7SBM+x1zx4flqYVBPVZw7b1hzPzMDVemfn0KZWe2KuSNwh+qf3OsrvSLj6sPFkC
Rl/G44KMAAS5HCY7euM3tkyL2yN1or2+N9Gq2rUKeJhp/CebXsZDzUmuEpxktfg4
YRNtSRGA3O35N4HlkoSyNiZjbJQULOsd9Qu8M4eSphygfvSpVjaj0H6nduQlN62y
XmrQ046zVBu5PU+nmUb+yOOTgcZxnVNs3EqYODSOpm4jALXJKQ2bMedCsghScM7J
qSAR2o/cT9pPex7ffQ0n4VBQHvRhWXbByWkMof1iCZul0G+/Ucu1KNVI65FTe9z4
b7TBml4OGkXV8WdG6l4RjlXf7C1aZqzZmo18YrtiC/YTd9CI4Zmw7Ne7D6uTdLXJ
dCYaAmEnSyLHqk8JNsq010+SxSlUE7Ku1JdlEmjuDTE4M7WTNWfxGAejj/AR/cXM
7CwJg9zL+tAIqrUruRgABo46vQ/f/RJ8hZLPQWcV6s4AAs5BvxXeMFXwYHXHmWus
OtqIZNemK3KQW0+mfhTJywwuLSjWO9QR2HeM2kg/dTqGZdUZ9J78daFHaiMhsQUD
Q6MXFAY1g9uNg3KahwGY5t/7ZOxq+nlYxrjcAT9h913ebY+XFAVNdQrrhjU5zVcg
OTXItnnNin+6BBezHhVC2HRfl/zzx7nxsIJGtvYODrw7ZXa4LEHyeUY2+B5zPdqB
1oFuN3aZJBvd0aKK1KIz3F0Q9S2RdsKf1CUo69Lvb1oiu1i4jJIxBbT3nd2ASeWX
5twtybrc8wBmWKIkuMefFE40N3x9U7ANZyqsbEI8/23wNHhUuZ7RdkpUrqoqr560
ijEJh4Zc4VaHBKUse2EA/G8YeY+Z2g1wq6mdpbECx5oY3eSF+xt31hCrCtbj+4Os
a//BURg9ycBAe/wLbUbIBPVyfWR14sJeDprFqYrJNEdWgk61OCbGxY5VOdftBWoi
/j6v2cEWIlbsHMywqLT0gmiwVg1rmozo9oabMN8S2DGeECR6Y3g20SCkhgT3ZWW5
K7EwbPV7Lls0aBKX5nIufVvxXxnTlFlC2F4Yq8WI5ZgrtAWnWp71sOWYwqoBjoZE
S5jsKPwM9YWNiwi+wz0KV4z+6rB03SgAi1RaHsBDNMvNlGdT/7gPwlqEOBklQAhU
TTF10T2/ibwerZufanXkQsifvxwiRSiJM2hVVeiLJiv65eqgPYERTmX3QHoj5lQx
wUziaPM5x+8P244wLzFYL9LVDXNBbx2ISEg70wsGRm5+y+eZSIMLM7i6iJRDqT2i
nkjKiTtNy8755GaWNXqSiRtw2PUFtFntIR0H8Tc1ZgBDy+UodMGuuXmIw0Ut9cQq
88Q8e/aFy8grWqJqVkxiW5f4YXc+9syEXC/n0DIIzqR1OBiSng7ko11BS7oSrCfi
X6Y4k49vKWKFEKUz+LoiAUdeCcXTyhXLxEtpJ6ddT5R2BAUjUT++gz6BhbBcwOcE
hFO7fg7vTS8v5E57yP/17xtU3pe0R7wHs6MNENuQkEpW9ZXLqIEdrjrwpvVFHj0B
n06GXQxO0tl7FmOd3Y3vPRiOd65oo0ytN6IYG5jkCOZwTXo6dYpy5y+RzDzP1nJ5
JaN5EBC2XV71RNuJgJ/V2vvYsMQvJmQ6Sk5EMyTg/XPqYeuxVHGPETxMEj5TZ79w
4ZPvFj6qpLDM4vnScqQK32NEsYgbAumdEVJqwRBQUFmX7a54p8xpAdDDHbOOszkO
Z0AE6ldzVw7eI6v5GbekWdPfNM8W9DxK612Sb3j7n4HsrniJml/Y9qTgmTgozMoB
mXsRveeTXJX4dXbxj0qXtaj7A5oIju0i5mD43tqPps9QmqcqkyS2stsmqRLqe4U3
o1pXhAp/E1DyNf25Pp4WzBRbqbwvMgx0ZhiUnrLoMhDYs877iPuaDiU4aEgNHcGx
cTiHIh5a3P/JOwjG6dG+LH3468NCF3MbF+QBean/HMnZy+CCGtqAOtau5lzr/vqq
oY/VTu22MGwTFLLRVXPi1UzvkoE9iXRkrrAsTrNngECHJnBcTUt9eXm3cxdNFrBM
qrPyXG9fAyxKbqaDMbn6RZE/q4T8WhU/YZxBUw4gzUWD04H0CRpk1twIPcWwkSv3
lbcvv2FPvgoTE4a9ZgAfe5DAR6vv6Px26+sGbXIGRRcqyGob8dKAGBeXR0+/yVNp
Wz7Z2sn2umECTGkL6pO5dMukM6KJ4yNa7yLgM3z5TbYbFaHn3pR6jkXYnRqxH22E
V0isixRVOkYINV++OynJA16eLEqMt/4Ygt3GFTNhuR8Pu1ce/NuXkzvU0ZXb7cGV
xu+dmozxtf/8Uwf8nlf8vRbM+tNQ7Hy0aZXF/UEBgncBEXe5uX88ktJXYGmbpq3U
qopEy8O97l/KKIbUwQAbX+lr6pIYGAkrSUvN0Atar3rvVKK/3B3yaiExlAaAdeyP
XW6NQsqFfKStP9HI0VMssNKRRON2zsHe7sd/FjsyR2dlTkOdJpAHKLhqssze6Wla
86AFYTG8oopthFQK6gHydIbGthgK0KrEQ+1JGZiMtge8ECS9c3LBoJE5wh6g+KFi
iNkb4s38/L8mZen3WqOs+enry4TD5lxe3u4A9MUPYa1j5PZTCf0MfGpmcW5d5VLH
Kz/zLoDHii6z+wXXXA4QxcONFf2XXqO2w1AQHhbTzykPFihHZEcO9nXqewJ27qxj
s4+jRfgyZcMNWJ/Eqv7BOskUptQtS0eq9clgb12b2pwY1FsecKQpSM/dOzo0IH/3
MI/0QriZnqp/KDWdWUmZsIN7UX56wNNvtq5RCECjHa5cTCxcVitoN6oaiXs78K75
3fNMqyMAKh6O6hrc3lB4Tb1w7Q3hv1KjU5sZfx0OmgiZwsVfyoOpTTBNqospiGgN
QbKWLyLKWfmf1cv675RwpdmvOK6YrU4wkF8pUA4Ax6/VRcbJUE+5xpn8VxxQc8UG
oNf+5xasDWSoaQ/wy4Z6RrCAFeWTzh90qY5tso4FVjsuGDelZndtBc1QqzDsC9z1
hW+uZpHRAKoTCZ6+z6T2+iwrnKLDsVTxfdpi9EWAnfcA4tuo99MBYz1uwwc2tLc2
GsT7waUvf/VF4Xw6hPiEJ6v8FBUaPlydKUNZJB0BeANw5kKEXS1DGpHsRCQqewAP
sJe+Jf5Lug9lT+5MPWOpirNNzxet72TajWjkeEU6TbKhU6znf6FVd/8iV893BVJt
trnGbXKAE+izD7eenysgkPgyyn1AYKvBsHKhQBK+Uz90OzAKvbm6IC3gchnapKul
+22Wg4JwtStT2sBgf6VAIlpzswYl9s3hOqsAul2jWV8/cpib5NRQBACisCOCAHz4
rgFTFpaeHRSyTFMM6eA76MvfvWGDRrsUDKquEtsYdWJWnFpo5NLHcbdorghHE7W8
7PvHIrZDYNCSMdotcDNO55W76qiVbYhvzMYwyWx7r5hZEtF21sfHJd9/nOFcIA5k
un6RzTJG4Lf3TIR3YHAeX9EyMkU+/govJTshXqTgxpv4OBEqNVYyzuW8DmsbxPGh
TmKrtyn1IsongBoXtQ0RIkfkf79v6iZjAzJp6HtobKHegQ0tN6eF3kl8cQJeLfFd
+ORk5VRqRzoWFrSlNxns05L7by2MbDIueRgggkd5fqmRR00pk3LbDdqP6buzHVuP
2NJfp5JxtZGT4DtCe6YatL+IrHS0rwXyTJzMbSnEyDzSDOLAJAYFr9oAfT/PfU4O
rlQJNTt7koKFf83rYQLvWt7xpQ2Cpl69zzXyu9G7kWyKgrP4cPxhIGwC68mddLB0
YgjRz5z9vuq/HVFBBbo1GVFMqTD2MAL1gaz6Xza9BVE8iZpy9BoyqpGDCl/dH4Kn
i/oAyUy+MiRN9mRwzAqDsAiJKIvwwGGjLP6njCgoN0JsYHB/EabOP3Vywp1mFGXQ
c/zEzE2ZscJp/nwXNWwnSGITfxYDy0izruf/h6bVngiv/gfKwWQGlo+BhYjddltg
JAo0vVmDZ+Z4DxXklCF39YAIRYFYjdsl9ZEzYm70sSJAhKWxhE2Z01B8yUZIDwGe
77+SjB/f39o3tZdc0TIqkE4DUVRqKwe8TP8WJj5r7DeOqNtXIfb6azKPNdX8avFq
8XI3+slQ7R01ZJnHuCbMnC3Dm+ZaFRIfV8LkM0JpruLjoIRUfbSjH0GT/H4ZBD3A
FVY3BS0ReDJ4pdss52Hyz6AZhWcXFYPH2mmtsBYF0YN+8DFNVaz9aWUyZlwxW4Da
UwbDVEjxw2XxIIABR25elVHKxbLd8dk/UoXrOow3LACI9q3mjrkln6u7xLEvKU14
eq2AFJNvKEWFefY/71ipYKj5HOucNv8W95Pnq/u4Cn1a0QNWiynlnFeB/bR0ICiw
SeemxsiU97GGXL+PC7+TrElyEJtjB8cFyz/DC+VtvHIAqzwo/6UC/axwO5fRnU01
7egVzEn/GwISt0zbZLhJCqHfzPYT/76KpU/Gs7qYeCllcu97/2ltTXviOagytBlK
tvQLEj7Z5YNa7NpU42E6jMiVGkrxH4Lch/vAybE8yjNGwuCO01x7udRbmoWa6oQi
YHesylFz7DUE8ppO8Z5MPxrRJlpy35GF3OhU93Owy7S/gix0AeYOhePOOMetzfGQ
doTSmitiBezFGkEg+imSr9/cjz1jCrg4bC4dFXh4GzeY7L5urp0IrxcEkBxGetS+
zziYsapP13gvPA9SwrLAtfMSizd6ZQXHxy7WFC46ILyPdS4rMZhRZ17XXdtSE+25
lAeMmb91iIUhV5Q8bA6r6ICATM2E/057+9s4qJ6vJjzU/GYlENypaFiUGN4llzPM
Iw+PZgXuaEu4vMRjDzF2KoCE3fB+Dbh9qfBCki2ExcmIwoL8p/9lkMZ0xVd31OAg
97K8KCaIkLB0vpYVhLK7wFEE7QTIYgTD5xbQUUM7BRRObo4CKVAtEQqC/TRqtW3X
YPprPMT97Vb8QhdYrJN4h8wxhTC65gMxis9CeIxZ9AHwDmB9Dwgdw2R5FByt/T1m
qHOQ4vicMmS7LyQvUmRKMHBUzGg3k5T30bP+mQhczjmwmQ7bDv1uU/UcxV7ztDNB
o60EKmT0U2DPrbMJjMvUttylJ7dSJxL+KIezE5TI1+6wmbuYPb/cuQ0U4g//DFPU
xvUN2bti+kB2ALWeUpRKUbNqhxTpUc7RGHUwI7uYsP55Pme0htxLgIuhPXTIHHaC
pVMqT9Sll/ltSg/W5daCL8LBNPPlLWJslQSOcYcLSMHpilL/CUd5oYduJH8FYIBK
HmM2v/NP0BcnIKPd3d+dPjD4vDBXE+G6x7L+nfavTbcBjRNeGp/e+2gtq/iDOu/6
tzYLOL4CeXj+aSknwUoFR7XPMoKGRcI43AuPWfdjwDdNz+ncRSs9d1m/jEjCyZQQ
qrsJwDNAkEHObWA9+dEz0sZ5daVRoLoKKuew04gW2sE1WpJ756O9SSSrOWsWxXi+
CaS0FyW0eJgMzWWYbVnWPxkvfIXfV63KBPwkOGemR6D/DLU9u45AAJEtz1Efxpjm
ehIN/Tn1xz1YFNjZWuLd8cLsMuFk6mUz7EvBm1+WexmFw637RjEODYcoV5y3Br2r
EZbPmS99AkOz//0rPF1OnkX1OwFTyW5UPRvG7Z2FM2Yzru0adeobe6PHkp8enDcu
kCak7nz+8pESvJ11k/9Yrdz+QMcD1a/J77DO/GAXtvgUtRtP865UDBOOlewyczAe
gZJgZ5CVeKR41jZZ3tubdGzcspV4TjX50/Ic2Iv8I4LH3OSl2dBghfGTwyR0gKvO
jJVhVngocPcMTNWWd1ji4pYa417KMcJSGyoG/btQ5Vhcc4sjw+QfQ7cDAIoFiumr
PHQ6YHRXAf6kXTlZMzJkuxeehWfIwvsi6bYHk32K3xHUq3X2p/PCexJMkHZIhOby
9X6jtX8hNCDwjWQvV+/MFWMwbGAcl6oiW1Cl9KT9uV7ApPT3XXggdDNdl4IHfnCt
3esoyDPdDZL2GZgWtYTTKa5telcAAuwWmxRQ2uPE1SbMrl8UDfFMG8ETnaJ16cn3
Cn7lA2i70nrD1BMwk9EJT7iO3tn8w/2SOig7yQ4lrcZ0kmxk1TQ77vN/CeB0YFCh
T8Bh7MPr2Z1RODrOFKZEWYKZFdjq0HiZGjQVJFtPghwpZ9HGYbzKxAZI31NXJim6
jXyjwOQ8UgPXTUzGs8kcu7jyKN/2lfKhJ9/kppGRbUXRyJHJV4Q5FwGVPPFQ2tsJ
m7Tihgss0scRwy42WAQQX5LKlcIrL7NShbOvq7ERAxk7xPngnfN4pQTmB6o6jebi
nRWBiyfARJTXZWmRPyvMzAS46FWjaKlf63zvOLMJD/nzRuczJWmZMXB+SZdzqfeB
AQE/ELaNRO7uM3tjupXw2pJ+MB2V8aRXTxns8lOoOvoW5K7AWMGaHbvtyyNPr51L
3g7PPJVxoBcQmaL/qC4i2t0asBuVt3lNr/odOzYcl1xBzr7eC/u9nMqf/t/GeYul
We9gSxrWYzt0bHGvXgB8US8fvQJvXn4qxlsQYQFzVlo2r1Y83f3zCBXo3u//5r+N
UsjBmjiv5ic3T2G2lVl9BUQ7tMczSwZAG+R6y+2B7nkCcQ2g6i+qnr23nP6LXEAI
3xNhL7XIiWAubHCcNJgSLUZxxJnMMkrJzfbulJakbd4uxigKDf9yjt7vce8nM6Wh
cXrP95I7V1M9Dmu32oGbMEWdMfW9XLPBIxBRQyU4WLKJVQwpaLtckB3M+F+7FStc
coYfqU27z/dfXkkIQyaOIsaCi2dZIe/zRTkTcIF1+yLYeJJa3DCdlD46M23AwBO0
6IQTCEQk16T3Vc88cEbm+/cihHD2lydyWi8fQ8u/piUL39bLwPaOSXtRnFpr1ea1
l5fdtLLHjutrM9APTrkx7cSvTiuwLK26XtMU++0T5ruYBzQ10a4Ob7nCqzfcesDz
QfpXWbpvfeHFG6KMM4FywpTSdp8xHMNex/JII2DSCciU4WM9Uzpa5qbWTee4weWA
sswcc3MHIydF05wXpMIxXw90LboxPwyAm3vABpW9Kb70mfC62t87thOIzDpwYVDV
SqUWPo8nRTiMQPxN3UsOw2awN79jN+CIZzK5fxKKHEqF2JLT0rcBFQz85P3qUJEg
3KfcNqpO1m5y5CsZoYxciOJS3qoWNWmXUTp4SuAxRnSJtq7tO3k4dEcPKHSpMn9B
HouGAoI7c9jTMzex0B87xtYr0xWp8CF2QFsAsU3hYUeVh+JyE4liQMVRJS64vTx1
QpZ3rkyYhrQDw8NCsmm4gDMA8Tnp9U4wVY07S7GlHrVNfahKKLZ362WD5KpBVjq+
ufZHgidH2UzPTHBZQmOraMYRQz2C4l4TH+7srrDvrhXpozpkRpXStLUvF+GuMuKA
ZREO8J+BdHtscNQ1ZVvv8y1tNzNgnbJ+A/gNoocdU7srf4XzgVVgly9XTQobYsnD
wVFAs/IK4twEgqr4+63hc9lJ3Q7REfCpBdlIVqAUYwvpz0ahG+YLxrfNZnTnJ6ZH
rKT9unf0yKaVyPi2c4eZbh2FshWEe+/HlYJVcWESPBEWx0iqXGOkbgP7GeYvYGjj
LDeDRAiUkGVGsElwMVeAO7r/5oZ2CLqdlSd5kUAUYW2aVgmOZF/tyyclJ4Ki3PNR
SMNwDXt5SVbVPexmFvP6bFVTJcb5b9h8lk7q7+3VhIrTPnWeWxuCKfVW9GUxYqBS
A+CI98/R+vjCPfezukiJdI85KHrHtTUAe5X+YxaRsR9f36zY14RFGZ4VIwm77PlW
a3bie8MUA5pcWXcm4xvh7UwT90votSlCzA6VCBq5bXXDdQysuwo4sUqGQ3xd+Noj
yENnuPNH30hj1hkerVmEpM5rF+HE+k2qqG+h215/ygDDNrKfvYjY9Twi46XUnTvG
znuHqE55akJyYKMBf3GYGr7MLFaokgxWZnE4hQkNsGTbj9Yu5LXDbVI7K+5qJEfE
Bzet95Exbzs5LH99TxOLiG8OzL8F4ToinilvhpLjVSORWTmYHW73NXgKBhwn7Y4w
DaUWJG4ewbJGs2jUvj6oBXh13FkAErY4hSvgrJyjjC1OOxMID0PYfE7ovy4hsGp2
c1U4P1g1WIGlnCOW4ugMND9pCvGYM4OnboraFRPycUx5UdYu6TQZWVw5LLWkLfS7
U3zM95jW1gm04G2RTOEVBPlvqaCKvBUKIcQRs0zYcLNrfHs46hwKd+DjEG26H4ix
lbDVx5qX0/bvE3EzWWR5uu7kr2GnIa6ZQ9NUB5/yMHj8ic7bLCcZoPJ0uTnKNpDM
6vr0/foPcOAqb1TfzjLAI7qhc6sTwyv7ibMud1Zf1AupIxoZwBls7rhmgaiix31y
NQ8pGDZT3LIDFbBIDN5M6R5dzITdsmD+Ib81EwTWUPWUiYkIDu72auXdLifE6aAu
M49NwgsiDWT3Ca/Ppt+hWenw1wF5qJ/D2WASDQ7DMxRxCNjIDuYIDvwujwKxNeuI
WKvFO7sRtW26+pcvOld0LX/+JFZtCyRiLA12nMdknTMd4uLUTCpHaImdzwQUpzwb
kqba4oxrO6wIxEOQaqLg2rJxY1rI+Wm7DZZ+wC/27mEPBhOe0mxVARKcn3MUYjeT
TNb8N95cyyCnlcNN9Uo2zA7GGU5KnyDQPrHX1/3seQbz97SSs6z15R3f/LYUFkaN
x5DcORLSch7P0nxbHYtfUDvfAgB4Tq0YwxfXVtkVVuu/jDKSUYhIv4HyuQyxlAuz
KVyuCCgEKqPcfrg+gWDjig/mYeJIb7zkeJ8sYwD5sJB0tGOb6v+jxjREYip7yH+H
SrNaQKVBi8Y60vEHxTj5dS2noxDM9mlJ1ni0MyX5zXTOLjsT7WTPa4ABVnJ0wPwD
1u00xt5afbJ5HcEKwKa/G+sFe5FcoHzy0qJIZ5RjDFl65O+5AiDPIDSW9cSIylMa
/EQpi8idzs/t3QiykuV81g2Y9CRM+7VaNoIpvnxmoWtvaap7jG3aENxi4veMSrOF
6SX7maznEC2+VAIt9QUKw5IQQNSx9Z7paSVkQtMV8MUWYLbsZOSraFwGUtr/pXsq
9VkOPqL/VVA+naZgIcB6d1X2HmGAVa6xIro9F4hb9tdd/hy1iFlTT3/oGldMceIp
6WpjZpQ5+urpHsHkMNPDeeDuSD2sglSBM94NZQKnU5nGmv/oDFcC/eCNhDoiNFgT
Xui+mcwpGWNaVr+l772/P4kQSSOxplI1Cq4lqg7elMY+vDWaJXsEUZuQVp1jlfeC
iKFen9UD9lO5RmUJGCUyedXMoEalWb/RvXt3m1YiOv8kzf8+y9XQBYjeHD+9d37z
hQxSXh4ODiG+3qiCEW5DhEwIUXvpMPc2tP/pTbreIFnWiIN7sfspKGtptewlo4nk
bjT5kaxNEq1RGVPZ2BqURKLIpTCsXkbZ+t27n/1YLL8j1lpEDaPGWUgbkh8Wgntm
XCGNCnAc4EDjshgxNy5YWn1xzsL9g3k9f6f7KOSephu53t9M0vkveILd40A9AM7b
5+OHG7FAhe+ibJ5GLEAGotlVSETdP+GH4gkm4n3iet/57V6VQkE0gsuYqYRWT/C+
gK8VgTWLW1qmVFsC/6lmHodGGL61ApyhA/DpTqUuaBQSfw3j8uwrFKeNjbi/EBu1
YMBATECU+Uk8YiMIAg9hEnpXcySGCRNQqGuGEk3drH+TVB07rmPpsTv09cP1KkV3
X2so05VLbb2uya7kKOAcuhWey1ESy0FkTAbP9/1WK0QyyijAietqtVi3YIzezKsw
TbssdtKT+o0NC801oQRX3q0R0HDXigI1WjWjHjBqEk870hedIo1kJhtekJP3TcJ8
IqxEbg7dMJzfqts3p0cqscc20gpu1gIEeSUtrTl+oGtkVs7K1IVUBGh3BexiM0uJ
8KPPeuT4tKhQiZCGjOSoTj45I3ALKLL4fp41PH94PjW7tWet4EMTLia5X7CoLsXd
KA9rgC/oU+qEOn7eps+TcL1CGbIvRUx/wx1741dpVWdoaO6fwCZb23UAhrkiPaCt
MbwoXdD2OnqlHzC5FpmoRKvBI+a9k9MGF0P0Oc1vG88QUFa9WlD4AHg+xUbWwogW
EkN6swZyNQAXF9t7w0K2aEc9M3hDIHHSktCDPvCbI7E22IiwJ17DDljViAUFhj3N
oXrufCqy2dmEXK1zzKCzeBzCxm4RKhSuvR22Z24johAgAUNX6gbt4gTa7z8MhN5U
6ihoRQPjFidTV2EA0R1FZPdv8PVx2/Swu5OJ56Nh7OqQlEPDaFH0NL89Kc+HMsDD
r/dpFfMT64h/r3ZsM4iCXyFUKOQ4bbvfbbdkxJXWFF624sbcgqfN+irlcExgJBKu
NKMQchpC48JJBg/hjlFC9fwp+bJc3ao225fVZcVenWzFmhhcqMdl8fePv8bxzlol
y9OezehHEyzV+GQJMfOU1aa0XUQ1sCQlEW7dqDNAM1FeEPCWGYuDZ+Wj1t87QYeV
mGfo/bnYTlnarefPIS6F0wH3AHBidpC3hGtEbdEWi4CJPM3kAnnId13cmRlaVO75
huoS4Pd81FRYjH2J6WLkRkQiB1uJg85e6WDqLSygmYyBNaAJJL0TlZa6g+FMCSsQ
PAvp+Zro6FqWaRhDP3xTXLy3R9S7sBsO4YD85ZiONFdG5PmIkYcXvBWvSjBuJXpp
3F9c8wSMobQMKx8w+f3Mjyhu9Lj/HMLGGYzLWh+mf6vb4FI3BEqXhxLbHIvC7uAJ
djC3QA/3tLbEWSbYo5xWwuAO2ZvCf1PBe229ipq/E+RSP8K5GZA3uCqbOCicBJWl
ok3M+50i21PDQ2fEOcH0aC0gRoaE33KhTJsNcdQpEJxxsxJ7hozELxpHgvbcu/zT
tPMEiKpqzyw70+vdKD8bySDOjtvBV0wMNQkQDmFA7ddoB16BU1OJkX8f5EvJCo7o
SFLZicPPLSAhe+O7zz2wVBsf4yH6bHjHbBZ32KpvGcr7XAjW7xLmACzwsa0T2g5w
AlCQfLU+toJoqQ+00MOSG9SEGmVaXveEiyPovWZ5ddqp7UyVZS+UUIi5vLIJS3hm
RrhRcOh/iRO+7FcMWU4baaTLoBWYGrJb2E2RCG0YKtNCYiM2k9EO7QwXL0lqgJxe
bxLkINSg6vGbNoscQfnVo9nf0MhbRZsr1+SgnACQm7aWaQhS/oKUF9gp7uKB4nA8
a946yyjU8pTxT1ouDK97pmWcH3ZE9yXKri0hlN8ScKW/msr4GC9OZGqyDintjWWL
ZUQNXspUBzS0cyBcymC9ud/zbyUqz383fwGXyR+8HNqdVebaojeavWBiOh2LT3RU
NJrnDmhWDkPPS8z4ZftzliHaTSSKmmMcjGkn2XuQTiMKx4R7/ux/I/rVz29CGd3G
7FquSnyKlUDYx3pLelMgd1u532bwIgNmzOMNn6/KCP06ifNEV9HmRESaiUGvXPDg
0u0DIR4SOsGAFFOEnJpod73X1avRcOhvIIYNonxeArkRFDToHPETpZs2r+/YvLLT
APstGb5XechDYNq4OjKFE+rgLe1lppzJhr1FL7oG4HEF6nIDj0b22GwNKXTf7ZQM
fEOg3SF7PvJ/WkJSZ0wMZTohUL7x6jZBfhyeA1x0OMUiV0X28qv9TyTpt1pnmySR
GlgxEN/GgaepJkGfpkXt+3Hw2K2LYG1byTjCaR2n9twHZ4L7FOHnc8DgXK692L60
AhUrL32UDWtRHDDk/2ES+Nerlh8Gi4JEF1/CM63zP90G7Qps/w4dlaEy35QH45Ia
GzixWWtzrLGT8Fqjx9QosO4tYYlnTd/z4oFF0/NTrpSzgcqVxjChTACWXolBZJEG
7vRMHIDTKQbPX85b3+mJ0L/No1zuYyBJQXoHjzj8NlbBuK0AH26yItGONB9c+iER
VCr7zVnP4KpseJ9BknSr66xaczd0wpd1hQ0z12g77F2BT79FJ4AywAMY7kmox02a
wHU7HRl3ACJcvdHuMyCgRu6HFpNges+9D3mI9WS2cOqOxDxWffM/ZihK6YdkNJRu
mHj1RvXBqVRXWY8YeVkxxdFoxzBotOAxh3unVJQg4uYHeI7nlnGm+w3d1gyfMkBp
6V4UabTU8bLh7rEUO4tkDg//aUZMEamvFV3gYSypM+yonTIJZXloLB8kI34Kot/5
FEOUyn4HxakjxnGsYrM+s6V/ozETFFRCQ24e2GiWCSUYt6/WQMCplbfYcNqYVCiK
iAve/rKKmb8SGslXuFz6webuo5V34Nc5X2vmEUudIqCC5IH/txc+GgJMe8MszpD8
I0Old3KM0g+dqzpiHkaEI6VOUh6xbN8uYLbi/UNi2Gd5J33ZoEmzrLbMnKtSFi1F
bxLrvLhkT3flCjI0vY0Gtds+kD2uJ2To9G3GfKnFG0Ru3KRTjzcTuEQnG3BDdTiz
dobdPqsata61VEgJDabyOLmTF1ppoE0xH+M1+bXh242tFw7DAgv6tQ4qZskkOo/A
n78WM1QyNv4NXzSWNS1NtDIfubMOLYhjBoGuZ2MLPkFeR7wAYk3okH0xuVCp0qtC
c2shpcKkylfLtrreJXMfLLNsy6pkojLFqEaAEgfKbKv3Ow0DzbxMuEFdwOiYnVdi
WE/2pT65EG1my9bh0Un76/W0QThTQ5uer2SC7zcdIzWrtLRudxQzKlEZFm+wfOnb
REF5BdPjit8i5mSExOF2OWBViaJUDOVxt91fn4JU8qqtT7FNo+ALYalmBoyQhceY
/zF37Fs8mNneZOMCQzHS91unsb+9FEejoPCjaddkc3YY56V2Q1c/ZIw1cS8I4vmv
/y8y2sWdUy0Wf0u/X/SuN6QG8VCTKVLU70cE70Ip+T5HpexYxHLzEYvSzl/VyOc8
eb1zj1zqyEhG4gdilKeNhyIIO8QktQlZJfJJYh50LSdkR8Zhsci3H+yHbPUqs+wc
fcI3O8EiNMbDmJfB5zdz6F8g8TIVTa7R+zqd+DMfveTu2oPXRu0dfX31roIwc0EA
pElZ7MnOLlD2KVGGFPLiPQyeCf7PpBU1ecq8/qkR4TAOV4nXNjxm4XjIFx3lj1Mf
AKb5Eck+9HiKsjXDe2JZIIxj8Aj7qkURxDeKra8PZCO9au3NvMIRBWz0IE042dZz
pl4TqF8H7LtXTS7lLBVLiRrUuv44fpuQFzq1Bc85/voWbvUMTLBYtnJxPudZvwY1
G05jPkxSkiquhZRAaIr87PVjeH4LJ12h6Ew+N28/IWGO/NhMOmu/SCdTEkUFUNR0
f3Sd0esjFx928iVX93tdSqomIbA4wNYqsNfbA930D9QMKJ5UQiKBAzAFxWbmCTHE
KqvFROyjchpTkWbgXfY9Z7hNqbI6kAd2m11z8Dny4pSeQsZdiufqKHOIvyLXxIGJ
vtZaOgw4M5rhPIut0QyHnIAbSBKDSZ4Jzkss+0ZU44BSW8qvIyhmdul6uQtc/FWW
oydxtKjEOz3U3GW73A2sZQdcMAaRE5B2QT/czOFoUbFY5SOOXE9ORwfE39/8Tpec
sLGFlz9P3oitoxGs8tnj8Ox1RKcc3xV28WcrrRnjl40pJlxVBdPobFivvV+PYghI
tZX7tUWEL5/ip+5LNv6hk6/U3Xi25sl9DfA3605R6hOAn5H+aBlCLo05Mpp7f+D7
Cgoq6HKC48qLMeKFLY843qm3yvStBtK268eHY4Nwq/Wa3N/NLBle2r8SrAyZ2RAl
bWg2WGc3C74xQdPsWhU5yd98LfOQy2xA+kl7q61A1cmgt7xKtTzbUfFzUsP1yS8n
UWRWWxYj6Kr6goZLFKsGrmSmYoxAd6bnjQd+pMU8SIKifQcI86cXesHXyKNrqxW8
WUSxBwEswKhGH6PbM72vbFzss8I81eYv+d5L0kOe5s8X8yKlJVVQFObV1JyHI8hp
pBhYVRW+OJ8wURERyQSGfdXy1plFawZXngXZcAtquSFlPLKjMIrlL8Yvyom6Huus
vZcEdJfR1mR1+G069rjyFRQ0pRApYf76/8iKrf0mGBpHMY6hDUZoYGoanVKhzYVq
vRYjDDGP2edP9PVcR/ss3RyORRuIs0g22ozk7MM81MOzMWgz18Lm05xszTUA3Bqt
SOcYGbJmLK3dEILQszN5XZaAzZm0x1Im5SsA9mUxymoYQfHsOTZHo0P2wecjgfI/
bXlXri3T7opPCal5eJMRfnyD+2iL5xmRVz1ZYStaa4TqnVJAHtct91DFPBknGSYT
EGT7yCufugfOYH1F6hQQYJIXK8w5DG2pFahi/iQCXHA+LdBnDFWym5/Qa1wrdUq6
RV76KgzhnfoHITV7n/3GAuXS+dYsv1qipN4jnad4VRTeP/dfS7B3M0e+TnMQEbAg
MMFRYXMIhfG1/6ZSg1LwLhTi/frEksTJGU5v+Y29KOL87sFFFP4alQ+SJydoAKOr
PwOn63+KJna5PbHOLIATKfaw6W5dDQMWz13pQDlvGGBSXyzV4+b17gDdE/HCA4sP
xlCth5mogmeREDP99CNogSAUOM/hT81Iphwip+kExwXRetWoGzDNlhteoh8qTnJE
rdrvbHGbjq0fEBUedbIsdjrgl2s7KIg/520FNU0uOa0GwvE9C2D+pyrgF+At0b1f
4nNZzsZlRNmttTpmHc/QWdXOJd1WI34CrHeYiOqbrca3xs2HCzfYL/oexEGQd9Fr
WXW08zSJ4b++XzImYS+dhzitOGp4ALqJB/AkUdj/Meky0HUF0e0FIKQlSmFPWIit
Nnu7AvMo3aYvpa+tg9WQjnFV7+znWQlRWOGMxMLaG0G+qZ9a8cg7Ip3vEWTC5UDv
UDDhyGySkhb5H73dVvGbGX12Qx2atYPOQTV19LUCDLClZ4shUTZj/chrTeIWKxdd
BkocHo6COWdS5TJ+yQFR8N8U4G82Bt1zfHFUv33zi6VkJJLjNO8QJzOLBVAxcnBt
VVEBruE5NmAfPQODg6MubmHsp4qW0GkiZvxPuN4NQNKyvQLzwzgReIjLJmfXxHPS
q0w4uTlWW3uhMvpo5OgiHEWCHce6pLZZYv51rmJt8ss8JdsJrxHGaMGrH1BoVZtc
4sRd4IY4C/6DWRiVmBMPsrQz00RpXDL1MiqRIlTE7bH/lrGfYHhq2ImfuwMV7Y5U
aJG21gWpQ9w5b47jkOCVYPeCtz8N4nwkDXqin6GouWpPzqR9bh+pRO3HciD8ut/w
BlYjq3vrPxP4GOl5jHBvv5oKqAjJkvF+Gmejn0ieUNTeVYD1qpVbKG7vPKVKk99k
E0rJ4QiyOhUb2ZlYPjRpxTrIs71xRXMJUBZM0ZNV1HD9DSOyf/9B0BpB7M5OO3AB
SKmaixcVS0hSL3fIz6exYT/bTr/ZEHZ1qN4V5oW3z2M8YugeSR+KC8K2A+oTL/h8
waSX82pdRkkRAhhaWMJ8Ok0XvoPj7dZ7YwSPpbTFH5iPP6m2QBHNFQpLasTI/lnI
L+lphmDpwknTYN787YaWMtjWLshyDTAZWCQ2JE+ngTKKq26Jt36BYNYQJNsQWZDY
At0Xzh5+wHPEG2sU+bsnG+bw3/NcetS58fIicpvdF/YcgAnZtDlH8/ZfktMDsi0O
Ir0daQKTojN6q4aMQd6vbuUU+G78pUA5AKCTkpUWt9gwmJhA3tVu7XwCW91t2Ttb
wiLG6mrjPXZfGtUhdK14Q2yPx/vNyO9GB7nVDfK3dPDXdEhNZL7CQLrjWM6flA3d
JzjzWmR4r3+7V5kiSp12ZA6nsH8pQg8Z4TY6C0MEk1Iyev4LP9l3jQMduyhW/Uq2
PtbIVUZOAUYeyLfbFqPodag3ofYRZ9dD1JBgaFBaJD4WVtA7e60romKsFgT4d/Y6
6WGuuK4ruV5hjXODSZUMHLRsG1LrSe7QXJYBb+QAixaB33vhl1ahnW1evvvEquon
BuLXD/N8oE+qAVigEkuzC8uIGVrzKmioMJhhQhKap3+N1e0j3rjPwATQkAFp+OQ0
jGw197ImToTYgdwyM7MS6I0rsuwy3wjfK8W0jYeRh6gfl1/UAwccSv6mr3+1JuYT
4QSrlOZEQNsIRKr98HNbFtbJYcBNQWMZ+YhrWGaYgf7nMlzm6sXRoeRaJg+wmdga
pn+02g44o8EpnzJrlTOPvX40M3z7g9ebkhKPlJkDXGcRiVFx5GlCw9NCiI870Wad
nx0xTFL82X9ZWQB74R1q6gAruILAQBi8uT6L7zZHNPfQT8LjmbNPPfsy6LV+nCaV
FSgXBcdzdLXrW1s6Ck4R81azolzvj7O0xD+qr1yjVH8qTxYjI6ewTzb4R+lLKy0T
WyaDK/wR+6Y8plGJw5VkMEQ6KBzKRosU70JHr4JSfhHoEvdCivAC36mCWHNxIlwX
vy9qPnN/MLlFZzPnK4RJdU/Nh+ELMCWvbhNihh9EB8HlFo/oGWeYZFdkIkJJavcO
xd/Jcnxknogi+Ierv5g5/sEXlQuMeslge0lzr8rAiSk+G8UenfuUwGC46epFxSxy
YvS85l2ykvm7j2TmKGOETKvPwT1yiKCSHeEttxZeO6RKSYKSuALtwN0QtaY2pu4i
fSnOlp6FiHh8mKAuO8wpPd0/g20Mg+NC4wQ3onB6GbR9yXq1olgRIyrZSGYwD4gY
DNCuT53zxxtxjXTPOXuH3jt7J7FmDGu0tS8/a/051yW0OQuKNwtFTRO9KiuVB1gE
Mn4ovuzuIGgLGjleY7w7gc3Dbv0gk4nqwmTnrSwUiFTAet2X0pjzxOyjZp5DQGfL
ZLlKFxdrg9zla5W/TkYY2Ii86YD2FlrBdLVHAoDtR3nq5krQCK1+P6w3DoTWMKji
bvZHKX1vH3Px+3yDOxN5cH55/gzSJaSuycOJBc+aCKcm2Zi3X2951s1tmQJEKXdA
1pUFp7lxuXSr8w2rRcsQfWMUYpUjlTCWI9GP0rFQBnxcgIO/RSX01yJK4caBxE4K
6qvs9/8+LkxpFpTKh1pVWiCob4z6dfE+AkERt5AG8E97Z/ZDovQ1sTCPlobf+gks
Z6Zd+NSY0T28znQfNffUIW9f5zRdMYqkdH/AlS8l63k2vA9C9yfSf2DmHtI8wCde
qdAQaIWnqtneeMWnnC1aDrww7r4EUrluIe7NEkGB7SHVip8oGRaIq59vZA4Zoig9
kJcTYV8GEvH5xBJeGggvj5uzBxJMAqtUcqCeWOgLpJgWVeHsdEvqcTSiGebM3InD
+vz0c6jlLybrUHS2GpnkUHJCXn/mi4HrjKg+ucu//pQhjfof+G+iSpkBkooxwg5j
rh5rRciu2CXflLHiN/7Sa88AI613YJbxuuO04odp7hrUAt3t4T1gy1k9DZ0EwK8l
JDMEbtHwR3Q8LxowC4NrdKa/Mua7iUhr8DBAWeUSInJZsttRd1t1vxbyRA4tBYbc
vyIDhFbUpM/A2vYFRkGukV6LAvxkSce98lhAySsgWfvuLZyMWwNACTXnh5/w4NoP
Zms722o+gY2P7JSo31LXhDaj0mvniGmR9XhAcEoZSkDlLczjKEVjpzK1IIMyQNnV
AZbYiRZLUyFdPWv13jZBvSH6FZnXiZojB07a8ox6kTmwwH0fpnXptZOHM9oYELfd
OD2rib00I5X/n0hSWtKbAqucG3MeuXBuQ1cDeoypX6h6LJnM09JtxCWlvTCINM5+
EXhaWeLpsU5+/TxCGEYd8GocUdb1k0fozMBdPUQSklfovE0eaRGRbvhQFzM8ft5f
91l4+zQDDFjfIW9UELia8hfpH3l8aOnsdQO5tsnqlA2wA+JM0qdIYcnTYh0eMndG
Y+/Zb1ubGcUgSsoPzyswy+BeEleyvcEHPDDEUVPI68j5hgXE6yG0fogDgh4pIse5
fnTrs8zKJRoS3ieq/YbqETLVbdFF/03tiWjJVmois1slh9vpfaBvo/HgMsj5+zFW
xDx6Gg35/Lcar+2Nd4TwNMR3ZYq7wWW6I1aZ8G2ry56mn+dXqkTU/2L6U923rLMd
JfDADTu2BJIjgfIHgF8jhCcfjYv0TwQhHG/zc0Svt1oBhzEjT+GmuhhUFqHGdO2s
eg/cPvnVEkgXfnSox3jWe0ah+8pNQa0ajvNFEjlGEtsQ8UW3VX71IIi/+FA8iMQA
r1NKEftGHA6fbtFY3kaIb0O2NGkPYne3xS8Xn5t2Q7COsnesqKd62jJYzM/GsBQf
LY4G3X55XmxR7Aa/X6tBKiEmT9FxSgoTDQigwgoq2qYsfopbh8YvfHzSjnx5rR/W
0byLBsrWiEmgMasRVZG9Rb2famWWVS7sinYX8nl+XI99xJokBsMNb+aLQcGNpTlD
PZL0Mx1QPAgEZKZ0Q0Tf6ezYq+qMVTKQk/RXUhk1p4mH8AQLG8A9PPdfdHtPFVjp
UH5FwQKu1Rlrv1F3nByaFJq7i5Nm59NWmMaGrgZEtLqpB52IgfWR2n4t/u/4aN5d
ry6rGdVV0wCi5LYZOJPn7ayj1T/XZJj7OcYeuDbcwxqwbG1UcDf0bB0+O1EphXcq
v2c8RRXTPnLW62D500RZHebfRQ+8VqGJ1XGoUCdFKBAT6dDmFcyQJgLIov/kDBON
1EkvxrC9LZzjk/B0yzZYFCMMdM5gWzIHZ2D8aElYmyWoQDAkAe0AtPtWgDkAN7JW
2XQylSDEcimOj8Z5iMCe+VcOlaGZl9cQPlKrZaxKj1ud2TXSyd9fzSIbEqvqzMj/
AUP9B9kNH9+vpfblW6KuT7MrbnIpD1Mt1wbw4+knDpB9agQHuvn6uop+qMUuFsrQ
HMch9VtP+1jO+V72+iUqlsSNWE42OqFmNYf6nsOAg5RJ6jJ2wm5eBXBoW3fYV1wD
i7vVtuEvaWHRQBhkDTez+8bUQX/Q6tu41/9LPO550mbIzmStfBX8wu44l4deJ1oq
50TdLM6ayEU7y8OFJj7ITAdTc+ycKAc5qVa/CZ23iFzqrjytgortWZvzfw7W4ykM
o42Rwg1FpMPxwi5PVVzHt99fMPKtrARYHiORuHcIF3HjwzNYUcNfxoAQ8Js5RtDv
kj9EHpqRLhXtkZZrTcwRvC2IueybcUe0yxWwrTA1tCs2HxXK9eOADZOxSjDSU04Z
+F2m+mqwLqE0Z98cKYaG7iy4CmDw3kt/stI/QWHkL2GejDjfYj96VWALBjgpKEBK
ecJKrlTQYept1CXTPmCtNm4o3MpGrwjxskGjF3wcCmLzJsqMEIMpQIUzf9+NW2zu
zO0Ad2k5vcO0jHgv/hOV9HhSFv8KIKY7cSTqeu+C8zIi1qXNv0GYSDkYUA6WHl1b
kSHJ81GtQQREb5fAzoBnkPycoVakW6iBYte37pl9nRX0tqHfUq5pQeuNjI4xyt1j
WPBskJV6AHt6huNAqZ7K5RhpUAFXlF1tBsMuDIL3w9n5X97FwcMpbp1w6cG7/R0n
f8w+PLW+GCMTyooLvrEEuura4L8Isn4AYCWPCZaSfV1bV1IpTSuOzH4olp2bqjTs
KMidRBhZBdtKOvquklasAs/poucKc8KJYszjh1e/N4CrLAcDUW8sh2xQNISaF1k0
sIeKakOxkjh7mU6eksDVy5fy6BHZ6kisNG5bMYV7Nqk=
>>>>>>> main
`protect end_protected