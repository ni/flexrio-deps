`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36368 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
xI6xg28eTBkT3MzzlHKeZNELVK2GGNaMEpodwayc4vU/1QO50Jt8f8ACjaFzhjto
EyWsCYOAMxc7hOVgoC8oNbSI+3lTOyykj96NN7ltvXXLw6KNtz+kdzejYn8oAW4H
bW3NqdqVGeiWKBQcixS9cvcUj6nUVFoAhoAmI7ELzk7EumJSId697BQR+77AAbYY
gmo8+dbqLWxEsGUjTPKqyyhYKkBLZROQOtaS7Eu3pHWaBaFTgz0ioq/4GcjjILke
3SUl1FJWT2f6bZEgXCgtzD/6yf8e9xrZqGNYkJ60NGzOnhfoNc6NkpPzBc9D2ttM
cif3IdwPbQWn3RaH061TpzWVh+F3CxRNznMWsYHL9MaT0S7U5rzt5G26CqsWJpum
AQzCp/p8BiXBiHB9xyCUntPbvAz7efEspi0LrGtyByGNNlVrRUpCPaIt2hKwavP+
SZnz7Q3hnJbFdgfkZhiRLC5Ofx5gSlQtOLQ634mHZOqoOwFv+mwHjgSSk+kRzBqY
L+H7Q7EZe3nZ8h6SmR7g0QTpci2KQQ+3nfVbSNLb2/g2SSiUAlKfU6yimo2zn4RA
uMKBcSwsVN21bBS/lEx6GPSw9uCCvpE+/jsk2JSF/f/Vtz/oWjf3DshWSf45+jfA
NbYcm5JG+8yYabeEt2l+hhlWeJaF6FYWif1B9r0Lz4fBCv7xceGWM3WJjwnA1Ciz
pN95uCjpFlv+/qWkvTDer7wh9poxbubMwUCreq7nn0OOq2fKMCNA+XwqVVzae9A4
g+NKMZiUn4KlTMXKKA/BG41EKfcqz6KhPShzX1Ol5SE0JqzN97U9Z/y8i49Ef+WA
L7wKoPNU0zFRyqAeNRKb23W1jvvNJhxWLmPPVQLTnW6T6+B02RKemSXDf8vQY/xj
fBDxOPgSufJ1gq9lwQE4/KkZVrjH+LPSMFvZml/04wfaatIVC95mktfhZI8HEBdi
GV0jL909/423pY1c2R1Sq166C3Ij1LuwVIro3WKZFPKItDqPhrBvsZkWrEvrp16X
nONFSL7LNZI+zgRR9AA91cOM3M0xlvls+yj19rGpKlls55U6hJL6dZfTxjF/mY3k
kpx+QgkSHP/QrOCEqMsgxBPTYvpB4pY+wLUmwyTO6Oq+SdvRviFXlgfPy9DZgULP
w8Cb2RuSiiDRFjAFCdVUQFymfMth6iELMeNvpkDDhrzu7mPnFR0Q+Fi3C1NRWa07
idQr4Te/i9HRdSQoARuONXPagsizuS84+sbenq06wjTR8H7djTwHW+K5y+cpU5cg
Z6cEPVvmo3Vm4wx+CtR5CRG9+G7GYK9bH823WWREubT1V/JaKzVamAATn3FDxE+o
LRCOJCQOQKIRY1Nm2NUVyfUBvfDw7u8QqxD2VA8Lo2POq+GExAjmXRVwFVGU6UmZ
SKtO/z+kxjqe/CJEpQX4TdQa00HObg/oU1Zm/ysdAfC5xtN4JsyI/YfQ/GGW4BNG
Ilk/yWjXB5o0uZFS43DNXJ4F7uaF7vh2kxEtw9dRDuTnRwJzat01+SoNHXrZVcbz
CodMhgJPYoj2hit4Va+zSes5XD/f/bgbtGW9VJn5hovz99e5o6fQXT0cVm5ceYMg
koNktf3NYzYWxTmTE2EwTCP2piR3oBm/61NsoGtwvpvLTAp1PNvb1JXSKQvQG4GA
Y86utvJrczTUkgVgtKQHP0SS4zWY/YOxwHPI9MUHsQMTlk0WaFTJExMzQwvg0ekl
BkRyYz0g+6U6mOoznixLTK76ofzTsL/InQTR3xaJTQQljXilkLdncy5Onw+4Fl4e
pkK2D3BgFYhOnVlSBlDaMFDVC71balG+ny7uPxFQkDmdfTDbX289iWE9lqJcBDP7
/a+aV0KGhl09HNjpG469CjOPW8OCrSWUcC+amNkW5GoP4AczPLwUrYQTR2Hpqqd2
sZ9qHql2iFzM9YIZwoTVyKe7v+d4VutO9YeM6Q2UL9VZtynl76WksiLxHXxWLQg8
+DA98L3dNp4YJvfyGscFxODJpFABQq0jU6HTwVyOvdmdvlbjIsj8gZ87MpJLGHOW
Onka1r0s99/lIXwSESCuCw01iUIe5/jkRiRdL7bSZlyZY64digy0jBxeIdcm0C8N
1s/wiDpEhKG3VLvlbzhEs1MX/Zr1yDE7V2GutIZv/ziZ3RQS/JrNvpfp7O+9WHI5
jL3y9MBY2DeN+OeMKI3NxpMOXel+k83A4bPwJQxdGXgH5X4vhDVBrdYnmnpLHDCf
uR4bn7s+2Hle1y568ondEkdw7/AWe+pgKfx/9whL8yrynWbnQFzYcKPxPbixrCAF
t9urn1pnMluzL3cSQdwEapl8GRARcgcRTAIum3X1UWJsEtolGdUzVSNaf1msVPWU
Yl7NXSD2HFq4wtTTOG99E/iAH53GkzKi9kcJaiYyj8VLRbmZY9BaEPO2M0YnjdAo
9i9JOhTC+heggWDrM/nERnz/8hWyd31K3fhgaXI7LIqi+7330/ELeWAo8ye/Blnl
CwJ/3B1GenYBK/9TY3eFBeOVapPNpXtiLHC2NAUcGH6OkBgon14VdPsG2vabX9bK
m+9uIHjv8ngfxEtSlBf/NLjM1qY4wadnd95YNIiU4eQjLxg8GnDWdYqee2ZkHSQH
7IkOyjlLmJrcjcdlC/OpWWtKMXjoHE5G/ORKXDiPzNOAlXBMQVSYGjZs96Ag6KLg
ea7aB411d9gE75/5A3S8wMllXyaZvXp36hb+DagblZd+IqqwqIg01l5PiYlVcA1C
WjbcZbUBLssURoxXDbOZU1o3aOiTkQ7rqTqco0cEUU/21g1LX96iTCzO+I3sJz6m
Vaov6Nq0tY8avrl1zvu2u2Km7OUQGldmG8ZYBWHfUp1Fbo+gDW1HcVh+WRafUyM8
Dph6LI8Ru+F/kVJNuWZmWMIvqRC3Vx+g6Gg8auPTFe6yL5blwk5sel8nfpVgWcUF
inHa6jMJ060jqzAdKPp+8CjIPwvTbT8aFtYG9a/jCLs5W0gzFqRzNmbcYIl32Sa8
uxcDT/zQknWfchNiSBGdikcq27TEBA3DQBPiX9Zm+hfz0bu7lWLes6ekKHKspSml
VWyKTR5sL05v07PTfL4EQhzYCb8gloYQthe+dLnpytPRTPyurcuHcoK9LQSSD/1v
T5Be2cNi3XoYibZwowwvdTKzoXGanm1wm879JVcT2A1fokODr8tx5QYtWeYLx3LG
N7tCBKb92Hbn0wFbhNFHLRgAvCEDufhwWgcfHhCGAq1/D6mwvFYLyGTZGFXLH0Dh
IBcqUJXeAUYJuPe/vF0U7Z6ZwL+A4c//ubxqBOu94VxAVdsDNEUaPZ6a6Y4GBVWF
y+kKtBghPZK1yzSH5iqsdWs4wmrnj/plKFfqPrbKzO2bJykIwqLHncQh+0pzYguL
JQKBvKDn7xdfslB3pyHD4jx3hfi6eGzEZKMCDcodvJtOZtpPNkjGUBcYE7OEm2fV
8AaAIMTdPfXBW9eNq3giwGxQYBihStMAy9tfgHS9YB87Kf5CdYsViOqvNXsvTkMT
PjrDw5MXMdjghxfLpqYQftmKWfaFU0xqY5HOnlS9iJkUveMKL9apoTJuHdNO2rNt
ZBgL//o1Vsotmf5nq23qLNHdtnH7ZQGHkhrdhSQv7pYnIArjikxoC2elnfy5Z8HK
UuXPdSh6MGagR+CnED+ZupXsfeAfV4BUki+GG+zAGe8ZAta+9bT3poMb2sliUSZf
srkVA+pwZV/V8hFXVLap2lkPGngGMMSgfGxRQ0NudHfhEUYYg5I/7mU8UUsFlrck
SOxcjZFmFJcZyPzhAes07EfZ3/T0tCZlE7z7BGwLg7mdK4czDlQTL2SyU1T2PYuK
gO51kCOhWlP6xrwjpb0Km1MlmJ8ZnWmWPZmM69c2eoER6GewxzHOPPyIwq2GuRmc
7+6/DcDcH1kGhar9TgoLXt+LpIJp6q3jL/j8wPz6gMy4IY+qIt1Dl1OVHH1zxA/d
wgBoJCcPh8UiEx4weWjEuLeZunTEB5euqbHTnzYzbLeGza0wEidmQ8+vyo7MW+PL
RKH8opRda4/CussZFkIMp9Ra6umZxer0XQni1fbd0CLr20KeFArETaMTM3taOM5f
YLLNfhKRvNDV/PGvOByHGFVOfXW6VNbzUVOWjMF0eb2f4y7gBbcITngWR1/HYsV+
v761esg9jg1lq5PhSG80h5OZIfZwBkYn32uJE90+TllJ9CmNYm02Wdq4DNlV8jmx
3cRuFC1jRxaSNX5MDw6xYED+s1IcRlUwGBZ7eRHyrM4xbIzYCkFs16TxvktHb/Sf
8TJc+ySYdNPDzhJDC5dokXFD19hxaIjXFte81hKs4UuD2uCSqEFfhTukJR7GjXsh
0NZ481Tx/19FLQukBqGDaoZtd6uwSuGRZsGLeuJBXQtl5dibVsUopUHfj0Z9wCXP
LPi2RkMlp4z69HyXxhpX7qD3IgjQcHWoXlSnUYgw4HWBxBYmBMUP0mrvzlkWlpOp
UjxNhsWKW3l/NEX74D1hV7aaZ6Qo3OJaFjdwTCMs9xQXDKyYYF6WsUIyEPHAhWBu
xA2t2IUC4v+PKZAu96LR7UzWjRTaZaquwd3oVQRpPETrcGEzVW/1bOrXeu23PaSt
7A15jXF5YIICgnpb16j37ovJR/GVekCkg+NVJmaAnd3xP+rLWcCDFFMBuVpuZAW9
knWT0dkaKFId11OHgUi7YOyYkwotOJfVziDlT737SCGTHEy8wXnmL9/8tUsll1+W
TXr8fCO6IYVWcD8ANWyNgaIM4UmT6BAJIXQ7n+JqPyR9eKI4DDO8k+J5LIpj7XFr
l0YbXSUjXyAQ/5oS9gJpZUXcdVm8RmffD/darCqsXRx9x4HNaCpYl+MMpLyo0k7i
Eo5XGtl3d08d6IJ+WaSCcT1ZuCwwcsSCONIn20267B6LDBUTMUJLTIPvfltt6f+6
L9taJ1A8FPJwuJ93vjAKhcd07v4mGqljDqkXsbaBsnwvrZb5HDLte4KRjI8UeUBd
6/iDPYPM8drVxuIuGfbzhpYm9Yi9VKWbD6EvdEFIlr/3oDsnWzUyZLob2hWIosUY
d/q3fDhgub85S8U5gZ5HCYW+XZxBI0t7Pn6yaMyRKs/kVAZfeapPjwAb7Y7/osxQ
MUqECSuZBQ6q5ZlcDLjWZ6//k9TiZXt2+mq+WQS3VaFzDQXf1s2EGnhozEG10kaS
T42b2aigaqGRnPbzPW3suM+DVYNF5OSyqKTTonj+rMbgNDkseRyJ0GBc5UOV2oI1
4GHy3sEF7APNGhOnbNMKuor8KjyTJM3CJHkYUNKOSf1dkPhaEBZRVY38gCfMqVhC
AcNcVEiUr5CTYWKsnwsyrCw/0IAHD/HydymHvovI6s9YpnO+jgARCYpKYFJQpIzq
6WY8+x7FgYU4pDMDPgADFhbKEPh7siFjewo1WA15f/fDW21hY3Se7UwBOUvz8WCx
KRfacEKnl3ptbZsSQrlUf+K4FdC1j3fFw4NpziwGv8uQhW6JAtTjAjeZOXib+s2R
CBWHcMCHcYex+GXPRvK+8bEg0x10nzH4I1e2GhvoI2dlztiQJSGq0qDkwTU6ozFi
+jW5LYg7TsFSMyFatCGPUtvzTUy+YAsV0ySz5VWzBy27JoGvHG3AHPIUoQooVhc3
J0p02Ou1WSrTqqwOrhK8B+6EAU2nOAYiYlnHbz8QaEGPgNhfOvQaVKeOqtf76jhH
QGcQxiAp+WVsLbW/ZCeh3ZxfP+WvIVnInyqz99MoBVjYuRKofp5Ndq3PKFJ85QBU
ZaHxzGrK+NLpTnS733tL6O6k8EtMC+R85pRT7XEf1dOnuVayFwPvuBkzYoSxetAk
+bD+/bPGy6bx0JJR/gA1YRByuGRvCeks654FLEYk1ksLPShYQrOKnhgCADkaLRju
vjAhEXk6MM3rbEp/cv333vs0/c90cDHgkbfjhTIRe6zQMIqjKtAqYUnydY51Ad84
iC5EMuKybsx17dQogRbKnCHDIGnFKfbbrANcDZQ0jjSbe3U8SXccTFA5R1Ds+BGF
lX6/rEYvqZifOusEvBmvyHLBMYiOFuHvzDZuIem6KfSjlkMKU0xqjYZJzarmlYpb
er8oWbJSKVRwl++wArN9MFmeqwciek4QJK8cxqVDc0szKZvCia/UZpoquPLAS7Nv
/RL+jueymiwaNgjctw4XQ0y2xdhAuGh6a+HLFm6/K9iNEH8XUYvpQTmpIs9Pn5fn
isHX9WVBayQ6rNejopakV1xNWogATVLZl0HXWXYR6S7c/bKgJg+mNMl0b1T/Yaei
jhOXMpKoJlfh/Kb2UwU7RlnViuQbq60QTy7cHvbvLiRZ9wqXYc0NDFYT7fykZfQA
cNGjeqI/zNgn36uYJ9aKDK+I8y5wCglWDezYzPub2V1kmQDpYcWGI1mANQnwDX5a
bCq8eyTGM2yq86jTbB1SRAnAyJVbgIM/pzYF0YIQ0h3CIBE96aJvF8oy6VNjGaUp
f8yVBKd71HC6cCytbONcJUe4yZYCWM1TxjvZlTP1Ux3JQ0xyopteZOiJUWgGHm8s
VKRsEkl59JrKTddIKcZoWLO9shaghFsTHSh9q3kOD26EZiXc9qu1yzPaoYsQt2R7
sYc2fTaXrUaCnlg0HinMWMCkhtcmRfCuiB5Prr6ZaMOK6DiiGinpXV4XQ+5YXUem
JAbdnI4FTWle9lyWl/qRttCcGjE2BlR83HAQgazXg868OvfbATlztkxjjKVboqg1
j3PxaIViwbwzPkaWmhARaXHdlRmoeWrk94Ulz9CCC4TDwgLurWs7l+iTcL1HYbcj
6ZRC+gnaK3Z22vsjAq2ncMUryJm9rspUqOeU4kTmiufY9uxvcKoqYTHHaD/dZAiv
NCYf/SNjmcgfvPzilBzo3B04Lfum9+VMwDcAi3LfkkyMdic0dZeQEkMj24wa0YqL
2ALVAGvHnZINTe4h2OHQQ3NZ1VzRCAqetnf4tprKF/TVy6WTK6MZmUoapjWscELy
56QjhmrXB1K5B7dLpPzGnuIODjALngcc43iK0uVXls+9S51oDmouIPKeEDveC9sH
WtyX0c1qeGOaGzH5er3JkMvVP+AoTvQFJew2eCtOkHyzYmJxC6pTBYvf6zx6JHXL
bL/hzybFhutPG2S0UtDKOkiD4QDXvfHvpRvxkxf6BMzquEqIgQS6EXVBI6LLZizk
OFZLziO9vDq+OtlCIknntDcQH7wgH3GTEv0eEfL5e3kjDzFawmKS/yGKvMqex8av
jPhm5f9QGlACZE+5SFylMa9yYV5CN89xZrvoJFROgvzwdIvsin+VR/ZtRcMUC9Z7
GljSLPxO0PJrHrji11lwKqJkLCj1hMGZNRvplqR1cH/81ZrjGdwPT8CVA7+IW0+Q
d6b3APpHYcNXsS/r8SGu9i1MUma2U3EQYluHGSA1lbAEVKSOwKKJs04joG8brRyF
uR97N9MIDWVWij3/MhNhrSve6Xl2j75GzyzTuL3gBnb6oJAkYduVv1M5mZUOLbAg
baFqLp17cIUWEs4mzwn7+8+GLJmgRU9eX8QoN7isKMg0DkDHLY78pkpLZI6jyLT+
jRrMwylomgvKvxTMUn9oavePEtm6QR19L7Dbo76pWhqlRJTx0tVogZlYMY6SCA0t
/KZDIAs+vhTZDWUN3i9WX1d3qt43qfGU3UY3NU6/f55LzFrH87LNVTOQtqDM9TVc
d8+0Ypkyz8QbKXUZgb1gQneZUzKjseUxYgTuxQUHmltOi15CcuHmbrjcY3uI4ysb
tOJ6/BhNzh3gLNerAjpPW4JZaQ/GZHscqTkfrNoZQaE/Tgt8iVln6MVddDEpuudE
tp4kksfmz0kwbzW64P7U6HH2VXuG2Q77QsN48BqWgvdHWtAovlc95kICwDJlUNYo
IlN6FhSbnAMEarq0FyW2EwtD/ukooIWLd3hTJ+/z+P3Rwn591imsXhpViH3/7V0H
gdzyXkGpDd+iAOQk7GVCRx9v0V90Fg7c9hbALYmHS74tdZixSh85WKA2qThYK4/2
0+aCl33spKYm9HTuRxx6fdQ20wNzeNjpa3AoaSuGfgU2wRhmM07MhM+ddbJXoUTS
mSrdiB+2uyLEBnJ7tB59+FVRG3e9tB6tVb7OojzEQlBXr9yEaimoTe9+j+zD+sRM
rR04Al6dWuIf0c5EpZNBG3eMwYOCLDyekRx4HxYootJGxYP532ZFko6SXCL9LIut
+19v1tWhofPBbRP1lCsyNWRyM5bbd7MKZoCbxWyMRGPjNRupNenftoGOV4WW2sAn
K/bMdeNl1dUe87Rj9PeynPYTWs8fvzfQArYmWBB24aByymv5etVkUoHenguBdOQe
FhGGfynTqSvL928ueEfKFZ/A1mTs7X37m3iiAPLL5L17ikDNA//K5seIadXm5/zs
NfUmDSckadw15PBac4dLnJS4FdCTeViZDFjd0WNoKYyTxJsCxZ3zzK3Tbg7XvnLQ
VyCN9q3XtKW3W07HL0wXz0OWCRmgcfU6menP5lw01iYP9mFyQLoMy8bdbFYbT0wX
MxxS37ZSCvNUv5dc/Yn1BsAl0LB4frNTlZV6ijnEAmvVgnb7I4O59dZCBxUmGHwG
gyOeRZ5DJq7+Cy7qyq7NMPkrjpEf6PiEmrOc49F0zFSu/Ma6ZykndlbtV51lREOo
e2Uw8ZoE/ed98ftAyd+z2pWf0egSNvBU3iXVcS3bi+eNOtupk4xP+s/tNWBZQB4r
7sI8E1ApL/HEI31cmdcXB20urodvJ3QGcwyn/+phASY7REr/2uXHjHkpzkXKjH+d
Kmqnf5HbF3y9oC7sysqjcR0wdQZbeJOsxL925NysyGZ3LymXeqXOuhiVPlEFY3Hy
WhVmEIn0uM/RUakabO4IiE7LSigf6n5zIRyzuky5xNLHp0N4l7aT9EguZAfpY6rH
2YHUgGdQIvdm0gYVocyAG71WRVEMXFAhED1WYt6nB27odsByzJdJYglyAc/tbIe9
eoyCEZGrMTLJjMClF11uoPm7uvZd5lELh88kAQMmaUjhydb9mdn1Pawvg4dShBe3
NIyhn/sa77dOFTF+mnZm4Jqo7ShySSCRob2m/RCVR/lpVslnKH2YYr/CI9DmvhaM
IU/a7PN/UTJ3emfsdo2l8+ov2RJ1YaxjnhOs1arZwI92WRtv8dPr9R8kfMpDiXou
JdMcG+DsWfxfw1WrPLw4PiZkd7CLi/sZumEAKlclcP4nWAtWYKrg/2X4hWXD0Xmy
KgF+beZen7i+l5DSB2Y9wrv9gk9ail3qonKXv8xVQTY3SkRcr/q2FbbNm3ZzgdSH
qzhU/qTi7F9oVOlTKXscCaVXiKzSHKKcuxBZyXw8YTQM9g/UgngXgKHbvQA5FC7g
28JSnfmILXV6NThb/OLOgnHpuomyDRBGVdjLEghFqBFJbnqZvXqRWZ8/8FvW+tIy
dxLftXhSmC5oGUbOnrPupgj0DlPoAS7OO1WCn43N0La+2/dCUhzLRZu6H/mxDxaP
afzhSaeiJOsGqgvZEAh3DaE8WeHGLwRqXiHjPfkv1zsvKVwXAX9MC46kRZ/UO+8H
j36/n1GIYeVnX5kCc/sxyu4A7xFbeE9NK6mrvCE2miYoHy2TZUZpFU1+9oSTFtAz
baa0iQdVg9MAkJwRh9F7sj03WqtCvX3Jsbn7q3hto1LNtts+bIRgdmD0qMjGzsf6
ZgnzgvSjxYLQuNLWm2H6elJsFNBXMffVQBJfHhRnJWLFr/FGYD27MyFJryA53eJe
Uq02e0ynQXqK14DeQlkcNOoe54pbKbW3O0EAYmuJezfkMW9pm5aTpG/udF7bk4kG
q3DybVgitcbao3km32GvSfDvspOkWg0/DIXymbbMH6rInVGGWe+E9V9UdGe/WuJj
wKhkUASgU+m/qh54cfaPC0OXecmXmMBleIvn6PFSGIsJcmyYgOJF8Pk8R0Faf3tp
fNpIMBF/dZycxM/IIjAX5Wasps+rPgCukpQQr2byn9iNSGt0CEJDdSpCFee8sX3e
mlbNh2vB5Mr9bsjCutfLgTm+mbwIIVS20K3UiOqffBAUIp1SFmYue8KGB50LUkhT
HgV0e07pezRuwprgMNmbuYyVWH+Xp1cdM38gX6oqh8f+mZSQhZUcKd9dxm2Xx73P
bgDKeaRu74fthZQcxBy9onrKFDpSPhUOLnaCYPEoSzOa7TTo4C7FwruIceUDbm11
rEWpurzhvXoiR+oUbMhJJVKxcjGRmjOAok+r8FVkjDelWMjCY4ijMBzZiNO/o8E+
JPs/Tgsn71vp/LVwwWloXZ2OBcO/KpGiigH1HxHU7ZGT1RnFPq3jTuq2meBItlf8
rVM8u2T0nk3vOK18RHast6SH+T+TGu9gMh3yVGenPCCfhxa82HmOGcwQzKvHE1cC
cz4i5VgyRNDOVCJ6w6TkOgvfkx1NuAjKnXdgVnFUm7ZO1/86HRSQBGf8gloIcT74
69U3Ei1bkicP5FaeN6fJx+7ehudp5z96332dabVQ1f4p5/yQiJYLltHfk2/SklpR
hm9+0Ai7qKCdZ+YcCVvylGg1DXTSukI279LYPO6DQtA+wu+g9rMq10vFzlHcUdDI
qF7fgZEB3Q7DhrIm7XjzmkzsqdMOF1W3x7plcUxpK6918UjNjPJSiMBfeCIxJY8F
yE6ykpFVI9A0Hd59n4yfvjYLuGvrqosXOateepy+skXx0RBhpfOLkBOm/TzsJr9R
unX6P1Mns+i2kw5CkbmO3z57fDhYMs7gj0gaKcGkccuL/AuhYU+KI/ggu+X+egV9
GhjrQJztmrhsMJTNl15uiJSJs1FfjnwWgDPprkSKb4wQcAUwiIY0zHEOKXF7DFsP
ZqmpQj7y7VGM3xQrdaHcObIAb1KkcYKTFjj0bwVLb1zvZW1HCw+Q83oBiRIAQJsN
s8oTLasITojS2GQ/Bo/QcP5ljkp0rxqMG07cDpBr510jlEDABYak2ByeD3Qf0HLN
FlPhUmxbbCHyv5xSlSTUbcDTIz+eqP2AoGR5YagQzotF7jLTxYD4JsogROm9wEQt
ShpB9FPi9JrvwFiOqcLSN8GgnxuX7JBnyUhKIiNF3IPrDy68kIMLSOnyWfHqR9dj
rtvXtIqesd7ZRvLSuNLZCcXAaRFImdKOSQBKpfRRbe0r8sp+su7/Oqw8kOBRPNJL
eoOCRGoIZbaiC9HK3cxkqa/cGWFdNOLcP9ynnIe9OH55DJqINuc1vuJAKbXc9hHp
4qGsrGh02C36DeN/8JY0LhoxXS91b6hI2zcVVFp01UdoVo1+HqHQfW6TJFmI6LXF
12wnXFMq+ZUyDbQ2+XxQea+4sMdfxKURHKCucpwLgP3SNXwmVBRdfh+0m8J0Jhlx
fAz2kmWlGFkvRdPlGLTuxItcGX04mJ6T9KZTuZli1DZkYCT2ZiF6/f+Ox96/3yGR
7TqzaXA3BGfw0HB+Lrc08i5QyCcrD7YnPNJiu65Ks+70OGTKX0gtIczlViGWoEeb
cVtuwO/gOnWOLEGAJqcGIA/q1rWAk4ybivlwI+5YIbYgsIb8ebg65Vu5upPcdthf
4oIIAOUDyjjIJPsJdHlsD++MhYq2iVlmqe7OFQOMmWl92iddJsbwr8cABBMunPdw
v3uLntBLn3S49PZ30VG8BG7IP0innmT22oRvzCBLNqjtcMZeGx9fgrRgwUGrGNfL
0JJEeaIwWyJFDNq45OsyD3epdQMUaU5swel0kGEAUf2GIJelgjVskwOobqknIaZy
iazirE+OvdRmljlJoazuJOmAW1QamtrsCF7Vb+Fg0NKcZsyIOboxvE958r5RyOri
9pOMvtrKgKSGlxcWODIdhAT7WF1lUtrNiOC1Aaf/MFSr3AL57T9oA89OF70oZKxt
jPeiZWlE2YoqYHO2+y0bH4mXW4gl6W3FnTLCab6K44pzrPmSy/oE5q9/hRaCOza1
JlupFxMFHYln0LpW/YLY3EYSa0cpqttTxn8Pq6Q9NfO1N2LSQaWwXVtFS16/bG7o
dwLlS6fNLjLaSPyd+p4C5zvqqAoyUthO0wK7IMQkE+/nEvjMrA0Xr08N44nJ6Ijv
BbVH6YMkdrYRdIFl5DAbS6hHkf93k8V4qOlsk58mH/ePra7E8VhBVbSimBFxB7/K
ZMQ5mn+cjoBleHMGojYxd6JEDbzYb4p7+FyURuhG/xw6qGHLvsrPEwmNo4uJMb16
QT43HG5nxRxgwpC6qtAvFQUDM6urWVWg4MM6ryaQsOEtzL6+IHX9yERpTVNADhBf
/vQLkBmsmK6alq6EA++AULI6ORfYBrNUj6/faxJWssK1UUL27/4un/UeLpsQhXpP
EeJoU+8cuYskeh9Pdk2EpkGmfiLzYt+kfONctyF+MXBQ05xL3YDHqKcE27h5XX7l
P/5E7rJS9XyfBuZoLLRW/K2A5fFvrpNc0QMgoiatOtDU0xyX9S5/WrmZKb5uoxS4
oiH4724g/2lDwYpiu1kh/S1ANIkbRsFe+cCQINylLw72prHpmvMQNgGup8Gv8h0X
+vniKT9+nB7WnVyuOiR//ggHXrd55O8wWNyezkCoscapLEzw8X9RbniEzFjiLhXD
JSIa+NaDax0bScORoLqXy0D8LrkyrXV/NXc5qdiRYab80nUv3iTQNrIxyQYmgsJo
CVDl+PXGQcazo3J4qYF1BJJLJIA+M6nLNuDJAh9aGNbTBMozMUZNA066/zL7PGp0
XVqQS9noND2Un/1SDKz0QRKBGwhAiDN0cQHcYTgcyiBb/LHfoPHAlotLXowrjGN4
vAScY185yNyAgUVOF/kD2jd+o8dutIEMCOsfE1nMIJEbqdwDPJVSnXv0BiDNAVdx
DxY2QJcd2I7nOuQvmdRPtlCB8rYGhW/x7Ta0ebdO2o0EghEjpAHx3mdgXKX0RVdB
lw0CiD8sjv/M9riVhr4tZHp8fvWQ8XjSC8npO9UAwd3lHxQ9j1WJK8AKLPnWk3Gw
W/Rmcc5u7FCtEL3B18RLZPF/UYWonHf9euOu4+g/xRvhtGsMAXlL/53D1tzxncUW
tAJhNcY/0XdiTPJgHvJGnM5tCuvRo/k40uK+5BbFUjNWvDhm/crJP+7bZuTBN2Tr
Gi1JzNmVeFoLqB+L5wJkoCarqacSbit3jShiMt7xO1ngJVFtwKsKdAwY9vxj+u7H
xxjcpjaOefTPpTOR7zmzl5iKnnntb8/ZC33rufb2BizK2aE3xPvDl4Oo25jdrwcx
0ib9hbcivw1q2rXLD4Njne5mLdJXqppVqt9gAwOIkLRxKzRbb+XBP9YvaPRf2IbB
tLDSAwalTvJUtaFb/2+hWpoZ9oR+Bx7/wA1rvJXjK8SMBIGtNSPHQ6mmf5n/wKHW
iZ9Kiil+yBj4wrpn7u0YagFoN3M8PDl00z8HI2qM3ekIM1RRa/Xp0FhfhKLT1aTh
C5Sq09kCPMpBAn7uDEIU3cMq7XZeZaEKXBi6P6N6ZWDzzKDN3qNqr7Gi/ZtCOdRR
z+dDR4M5TKtmAZSpIEYRY3nORD2U+yj4su0BDDd5PCCqexJBTsUHuVlzfaqmr9j0
WyhrChez8w/M4FvcIPIX5QNdkWFjLEw4L/RAUNEN67+Ck0+Y6kIa/5Tomb4IoGfj
lx36+5tbdOIGWklj6x002XGhGK9dPW0BrPzGrMVY/lAOVnNLgaYqdey3w5np2u3d
FgwWXiyQPBxq4HFbFOwA8FRu7l01q6f0bzmPtOjP/cRchWXPqSqOlj6e9ey2sFkI
yf+enNdlFAo/pd5rr010SQw7Z27zadgKUDRXIvYFc7ZbfPylTZ0aT76I3TroTduq
u5obQ9omQ8rsxbbQmOzv10ZW/Peg5WSd9klJpYNxwaFvN2PY9MT+o8H65oyiM6rC
YPPDqZtGPIH2/j65aTO+ItyQrR/aqp0v/FQgfHrQFI4lZ0bM4UGtud3m5k4a2DWO
jjAKxpkWEyPFDdqrhCzImM9k9aOXHE/1bc0iefJx2osbKGpmNgBG9nTOx+pO9yst
CqKn+x6xwcoTHamCbZeKymj0SzZxqJErKo01t+JgTRB2UWRPOd1p5qEHTDvYtolL
A5h1t3Trl8gkdce33iHWDj/z9ZoXa4QJmp5gF2A8krIllJBKGRownaFJIHVt+GBv
EuWfIYZVtnW8rj991Ohdeqnho2Z4LKOWbpkB7Dh7YUIuHJyYlHlCMtLWHas/z9zb
xMu9wCk/JDBP3haSsfzU/VfHqGdweAsK3oL/UjmbhyRRBu81lpfH3/bqGA7eSmK+
ReQq/m7tgv4EpWlgWK1AiUBmexIt82s7Y//mnJFheQN2sWJQLJlyZnnMKUhNerc/
1SJpUw57tfk21hQh8CKh8nPF9KlIZL0ZsYQTuMgQdtgNyRwXuUFh1pcElxDV8230
x71RSw16ZQPf73k47mzMbfDc+iVrmWwszLdPJ1J5lrXflHH7ko4nXc+VX5Asp/Uk
sGAVkIWJu8ZPRWRZGq2pvZGgvzLIYlVf19yf29Au29ZtWU0iIaNwJbfWBkCYmOOG
CGlX5HKKbI3nq4WEzU3FPuv94ob4JuxcSOkG6v4OlTBv/Nru4m/6ALdC9dX1o4Ps
Q+oiGdd+26re73R7h2VSUie97hqvsQdI/X5V0jdOq/4Tt50cHemEYX5RJF1ZxphX
ovNa8EzqvzIlUKxsb+aeRxARq0nV9RW5Z77NTf0Na0mz4afSPS12G10qw6NUC3Op
rr8FxC0jcWJT5D8qAG+0bhRHSuZ0NYCF5r1BZ0KoVivgzFCxP0KNV1CPbKvUB+L5
I8rivFxq7+QezRxpxjcBLTD7HWcVp9bvBFMIp8FPn6b7vtFbGR5F2TgB+jP1gEcL
Ksnrw0qF8/r1ck17HDsv4eqVWixdVrEEj/VIfJUTST6jIkDKYBGo7Rs+PYaLOeJI
6INnLXv/zeAfsP7WMg8x/HqtpP4J/O8hBf/q9iZAD88THRm07vGbPisD7Bi5fuqH
P27XtXeZbDeYXYwiDQipPke85AbHx4JMlFHS6domR8XJZom9UzaHpkjgPrRSOiCN
Pa6n5Uk5m0SbX9cplD2FNfUCPTO2QpLPhZ2jdaIMmnC6VJYuKOCCnGY6Ez0a2mDI
FXbC5nUHswmByY2E+1eNiPNpBXqiQ4R/xs5mMWbgbmYJDuxo4JqyhvAYHX2C9Lul
G8tgAUpNxiHfmHu2tcfAEfU9C2tgnxeXswxuzwnItMXxCrIom37n9eYEOh8CLDww
uoQ2q11Blt28vo1dSAT8J1C2LPAXlsNiwJFLF8be0OvG1AWDN9Kjnp/iksFQ3nUz
aKB+SoTny33yi0zk3T7UX/SNW/K3yR3rq6ktD2iiat72DIvMku40X8YDDYM5C20/
GPxUf+uW2coZbf61k2syRcdKOrFxu3vmcpYllmu4G0f2PCT0OKhgbEqr4DzIGRHo
eIouwk5QlIXmMUffBL65vvJD214UiD//bErcnyXBPedbVkH0x1rf+a23KJuvwo72
u1SPMWd39eLO5bZERvds3mKSOPPuhjzIkPT73eC6hGFsOQLGmMfz7i5weODjk8Ev
5tHjb1PZj6uHcqCzLpfMj2iQSEFFoJDbg1FQp7SH3NnvPpiA5F3CifIcpPSJhytB
4fiehRtktHDWsoQs3eRWFoVsCeSOzBt3xzUIx1hcu/wUKypDHIrlEpMdhowlleK/
p6PufgHKLxaemO0jFsj0Pm4iAoH2o6Uz/tyQvXKF4Ob3FP4vKJhMEjcnHsXJYQ7w
W201ec+jNJTxi9m/ae4TS+380XHb9BfB13Tf+Cb3yo768rhpcxJNKzLI9EXN7KpD
6QQtyAWLbQ4DM1atIe0M660cCmoftlcUg+Qzf92dJGXBihDo4a/9nRb2ueZMw/IL
N4uJ31VAo/ALvD8XKnZz6ZkV1Y5Q8We15EAw+o8WlMAU0OBBYkcwkFOpHKUsCNQN
IOT5XSz1/O2SZHhpW4gXXybtm6LDbiLogYqtoL4bFBlsrcrWe0Dx3oU/dF9GceWo
C6Nyugom/VtzDMDPMwxUSZMrofTbmQxEVP7tv77fSGJ0nlsW3cz0bTS1Ljahsq2H
dEH/oygKRR1SSniQvVFEKqCtKkIJzOjw1lh6VF7c7XPz4z6t8hsZebc4op0ph5x4
OS9A4PGcWosGEiJk+To+xN44p+mh6VNSfQTFqUdLg532gEGA9vXB07rW6RsHp1po
Kb1ikSp0RB+m53ubkY6KmZCbrV0CEFcPbAoV2ONTGu2TBy9P69EOWL3cGOC1uT3a
38Ng69+yz38WwYo7/IqYXoGjFrGwbW45sdd63RRaXfbVO2tMiMI5GHbxs5vu+RY9
PbZodeVd4F6LenVzy4IXN5h4g9LEH86R4WITKmoSLAaOQu8SVw2Jsd8D4gAibItp
WAVl7EosWNFiC164L69aU3BwO/pUHSPeDSxUWTGVr8ESNw7FVASVJ/aZiohuNooI
7D9dIUu/ON06T3L+q46ExCntFFUnUZnPchNwXqApdPeMiiK4+POFK7nLEvIgxuyH
GCc/SNjK9MCReYt5i3rb9Qq6dtsfnlnSmapgasuEVbYLOxkS/hx8ZlONEY0/nwL/
/rjrB3IeFld+iUNKqKax2ka72OnAbP6RF5QaZcWjIQbTAUUPivuzH+u7MQgeiSnR
DwqY8EAuYUQD4dqCw2GvnimxEjc9iidQPc+r/izJp/S2g3etmJc5ypMgWGEf33vP
mvwTsBLrhwZLNy94xh5rF+esyfSuW61mUn2UinosHZa5ncOp5h1i5eNwg0VReMcw
B5ug4BxgfDKHK2FhEkSQWQTzaGzcrObBDtUw6E3ljs2NhTLomgoE6VrOJ/r3xzJK
oNf6pvbo5vQ7oJ0Lxx+fuJdS4KfXLNCbaFR2sBmezVzyW9AxoB2Nnr8Oiw3yvxCy
Y0x7il2Y61dDUiaVWR62Bc5xFTgtYDthNkdLrvljxAUuxLOqLbT0Vkt532YzJcD/
bZthKtHZxFBZP4D4E02gx/HkpbzO+GpZxuJAXkKN8uZmPoQAuv1c7wWdxoDxAy0m
KDq0rGyqfCuRe7lOrU2cHWj24iXdAGEHO+NAkcDJ9KJVJiaLoIzL71dWbqPSA6n2
MFlnGzb30UWMETjkA7pW8kj8k9+ujTC5lcj19sTuGx6hvKeutWCEcEw+1MekhJUk
RVuDiIiGmqGgSpO7AQVvCDutsHX+gMHHMv8p6EpydxgFTjCRH/AcE8dINjwsdZqz
1Plevb3o3aSSSJCcq17AcxqsPfmrRb8i9OkvhparscX16DK8PJ40pXFUhjDvD/GU
vY7Ft/fODJamxIkAznDtHMHhxwiW8NiTRvwjTLiert1BUDLqHCaCxATzEStzLTTh
2Dt1VxRo32ShZdxf7qMBPKTYMariGXiORPLyWdY8uoyAhej03oZFIeme9gIzoQlb
pqojDUd1ZybHhIhvPLiGt2aLCOEmgdZWaOMw9TXIEg0CDc+RZJGhsQw2E7pGfLkc
3uf1MD1G77Fov8nANG7j2K39BrAlc7GnC18LO7vHSqgQNSd+v55pLFxVLqInYhd8
WUszkKH6jiTFx0Cruz25YzksPf48l+WfHDUIih0H/R+ZVBcp4WXDJxBLdmgcT1do
qfp8rErRg8MU7tOH+Znfa3W7yRZc7MEezkc9T10ir5scN3b6aspLsW8zRasIWCPu
JNNicyJ9BwX52N82TfoWVlCZaKfGygpc1pGxD9R+Isd21JMOcfAgX/tWBhA+hA1s
xSysksRKwR11UDNCrSTMRsTZQWStRPiC3WEF5OtSpEhWdSyBrjjmoTY8bSOWwd5+
TCLSxOJH/EieF9kNzKPGeQIIJ8/oVUBe2KU/5Kqwkozf7kvKLFLMpBU04NmjQckK
pKZTxPzoFL49FzNzvMiHlGj7s6639UgI2KvBwXGMRsGYrBuwVXrj5r11LMxGXAMZ
eMC95abNsqiXGjXz4k7re5UWgUfmVV63K9KDNQQzP5kD5ndFjj9D++336rcxnOku
3xD88fCuaetelLMEj7HxIbB7N58uQ2XPwAWOfY0vvNYmnzIgy5sp3R/f0JQjiX98
hi0WPPBU2HHF2TZIhfALXfLgMM0X7/HUNIkeXc7RhLIEOW7XyQbUkpFLAGs0Iuai
lIWehqdq1UlvpWFW42+kCvPIP1IWEg0jCmzFXmXBgfnppksy8aTqiBxZJGjNwg+t
7ydSorsZpD6q329/Rk/GlopGjeHv64iupDYxrqG2y1xy8+qP65EkV62edEODpbNz
Vlbsql8qwZ/hy9XjsHU/Q5YqhMsNR3F/PtRGHNvafkB526w5d2dO8Gi9pftnqWQH
8MqjjNqnLRj6mEc9M0EUvqwBD3/qiAYM06/UWlGzP6/fuFaqJEiw0x0Kww0r/C7K
dDOdiVPp2ukuy3h3HOVzrjGn7Qs/c7INetxxEwNcES4y6vu9tuiSinlV2e9uXOU3
apN2g9mGPFDpcDGqyZFRhqxfqU8ujkxWI116NnzC3KVNoW1guAURrkOSMqx4WxA+
Iya6DaaKRLYPovvshLAFxXrFx9Z4EjLQbWmc0x42xMhQuOmcL7dRoOZ6oldCww7V
Yi2vj9ggO9SZ7LMqQFL1hv4SpJ0WItnoXz/2FcCTaDbGt68lVDRVSiXsYHOCjVtV
5ONuoUTBhCRZxzcZd+9DedGdJ4MA9e0Ks8FNM0b0X6TFln8g9fh3MQvuzxnWd5EJ
c8UKGcLDlPirdTIs9orHGQd5kH13OA3dSoQNged0b4xDxmXGt5UnlGUGeiimTYKR
xGw7vwVHu5veehZ7ccaR4vLCUWshNx+y8YuELomNacQr1KCkhuJWaIlfiq3M66gW
GmaiSDB053vy5fjyMjfpvolkDovuecm+nIp2BVEqEcqZMetfdpvWsfm2dxGo/yCZ
TFg2f6SML3LYK8wrCZrkZcFy0olrQEN4nF2ttgUwYN8C1ykK4jkoRZlsxBjfFkm+
lmRITMo8jkA6uwZuol+TcoUAXcsgDEUi7HIJsakF0ihOd0Tf5VjM70r1MvDfWi2x
gxWPdwTmY+Fxf6Xh3HfspaHiNnardagc3VP8WhlqpQoIcBdJJjUvqXY8OkzmIpCH
0R7rQ40ph3qdC4gq4Pt4KiOB+Hfbt5R6kb/0bXXKg8SlZ8d3TBf+VU58AqlQLX3F
KrX8adFhgq4m2GNXreOTlEeIfwrGOgGzFAp0T8OaMFNZwMkwp6Rs9ghf/fxFrdzR
nseD2mgcPX40x/oFzZI1PuiCJiFteCroSYW6MCjbVrZ8vp3d82407aa7AScG8Jwq
vrBDPbTpClRgOyT10pjshDl6BcBtyj0yzmc8JsKXmgpur55BijQoDPveWoILcW2a
xMVRv0u8lOb9NAEJ76ahjOfe/sKhzxa2T+jGu7bWBEo6yxHmeNsbPSZI+Y9b1fCS
di6et1Bew4E8AJmZ01QOwdPAg/4nMjwCnhOJzQJJsu6tEbFQ9NJcPEz3tAN+34W4
8YfDTwxMj66rlyH7l+tCk8kXh95n4MsKfGj4YCYNwtvpX6T+/aVVTkDYrCA21Esl
aecL0iMXkHwvIa6GMnegEu+BMhGg530pUCqery0x84i18HwwqByXgh16AZDwBjlg
IL3C/zwIcr5pdwOSGyqNulBIaod4d1UlwDIJt7e/mOpiwA/eIqK/B6NJ7vcVh2qc
LtXRFPOxEyx1uHhrljErboX6Ds2u+UOq0O+I/9CgSKUvIzXVuj9BwWJRnPab1v8C
C07HdlGQAf2RPI9tVCK4n7xSy85+0hF/lgI85qKyq690cOHLXWbWX0vXapo9eXgd
c5JBYjlgNSREmbsMPXilsgA2lw2vOGdIK3CL7Ma4I3S2lsVH/rHzXlZqWh8T9vqZ
9eHyyNxc9AeF5nJv/88vBzYdBLMvHgU+zqS1cQ/z0mkD1sQPCk8m6N70UawARcJK
UhyGj5YmculJSCimjIY7L545SZrt8u3/T4Vd029Beom7o2c+Aky1ZyypM+912jHm
c5PKDEKvGB7URIZrIVrbAn2izrajGq/O2xaDFuQtzme6QUcojQJD8k9A+b5ob5Dx
QSMp3QuD6GN/Ea56gHIPPHJchERL1j2BXmNB47cR7uG/9BSqeRYUyK7AjJ/rtwOI
tkj/MXdiyZsqHho4++jQd6CJaN3h2ihNZUIXrDtC9FZOwyAc9TNpFaNogSL7z+u4
pJ7kJtH8AevrXZTCePeQA8+2TBdjAi7/wyRZYPAn2G/aAi5K/u2+Pe152lt8M8Mh
TWYC7/bVZs8aL3ydcXesYIBOZNDge2qtkrimgqrp4TaVZerV26ygDwOHPkzkt7K5
QAIr/Paom1tg2X3PaAlTExa8/IrcJokkVheudAiyY9eEIVYTlR4W2WXj3OgK2LTS
sd+JWpFhupCJxdjt1RNVu/MrFgFi9vc0uGr8uwvcy1jnDEPxWtuN1foZDDk/7Gdq
dD8i9d/AZ2j/dWRIGVYJXiV/i64ZSjwG+DuBm7WuiDB7Xh6ogXADPjpDcncEJxsK
Ury142RwE/OaCOKujN5HmzCUQNw3Yfan9hl605C5aaaTwNeiJtmZ/X4hTQN2i5cm
eqLpSjETtsyXmtCMrGa2axi0EYQjMH1nRUpgSx+IZj6Ij31XTTgFXVokSI07yft4
1RqejkHjW31wNy5lEE3oBouZom+KHJcZRCQxAMXp03lPHvsT5stTeuRGaTwrL2P7
3tse8q+WRHho0DoFldg20Q4417md9vPJjRJWQAC4Xhv0JfX1VIvnSmIelpBc6TQj
D824IRf914mAUy9GZqPbkeWfmFaRwEZsdr+sE4kwdB4GRQX49w9w67Ucq97nkLva
vKQxosH/LPIhbbjDA71p9LNKBdUHKzcmhFDDgwL6zWIRSRwuQ11j/ibfOUNFZQN2
S52ReX4flc7rZIYNwMtGwXjS+DKnmxW91J2Jqvm5kzLTym6f/C4bbPRO8GuR3FZz
d2t59YapA2kEhGDuMayhSqcnxcmKfa3SQyC9jC0x+ojJXxNNCuodDioQ2NuY8iSR
QZZZBwkURLdeUknRHBcC6C1G4GOVHrPOW54b3vHkgm3B15Go7kJRju1kdE/EYvrI
1zk8O9wIZR4XjbfOmZr0PX2bBDvFQLBuNhbQ4sJZMmTGdDyJjFfqFW+KEd7FnCSA
QvZu8KztbUW07o4N5xttSMOBH6wwX9cnxF9fTok8rjUzb1hB/lbk0Y5HWWPlEHEb
KGDGuvQertL+4gjvZ4Qa5gL6XEasImKeG88yLkGEsaFdQNv24c1w52fReKZR2Em/
ZJrSa4fEMlt6korFV2xKhiSIH0tfEEhQKbFlKM3HPnz4tFZq2y1H49g8WW/7QpJZ
/3R+mcfXPYA7YbD3Ed7V7wsUUVk4+HBr7oNXYnEpiNuDz1epYKEJ+u1HcuAy+5sH
9e1fYmO/ikuQy6Bd2vrQlD+pwiiApkBdF1cCLW1OS36/lknCtKtL+HWvW6sMOe2i
3XY4Qk+m2bHeYwQWyGt4r9h0fLoTCI90y1VLxzhFJAB38B7C+VlvCZP95khp3Q7v
Cc5429qYfpVr2bwG0a//KED4FIdnAOSJFvnkQvqUjgsLn9QcEl+w0tcpHtEMFeqg
w0wceS1wI73QEIrjMHHVSiWsuz2KHJPXkuf3VI/hJbg2E9u6Bx/4dRMD24JvE91Y
V1nZJ+F9ZBscGuu7V7deLsm8W9jASNtdcqaYAof33yuR3zjPcwKHOkdG5xKRz/zc
2SS41gWSxZNv+L4aAQ3D7Lc9q/ay90gQvYyRxTY1KzyrPjtEUMYMbhCaOdixnOX3
HwVy1fHJGXcvG2wGXLtDfGJRCRAfAZaeBA6HAmr2OOKJD6bB5N0LMwSzYTz4zhp4
7Yx1WOeh6rNhfzjXqLm1VJMFILb5OzHjLVaXnJwwMDBTACdRspAXd37QgQ/FNOrU
dxcyqj4XeCKc6LNu4WJSTQahnFu2fesnf/bK3Cd4t37ZTGurOE3eABshLEVzZldp
c7Q3xbspaTW7vFMVmmKq6rekjtov1kzE73VzbXWmxQebqKJLQaLvP11LRZ0k6Q4W
8FHVasUCIAhuTOWKPQ6Ck2kVjxZdqRohtcIY48IEh5MoFGjbAcqQHg7ilpSfAkeb
Lp2bBXDaXHjYZjZZqw+Noj7HZOwCMHaXgsRHrP6ZTSFa0/cPhbNrwAT9iXUNt9Qp
nDiOx2qjEqr6laI7kn288YbrndVtFZFVeKvLpJUnyN67fNjWTWs7uu2kFBLnhtij
9umIRMV4rABiKBP5qzlPheG/Rk9IgHxd3q1MU/MN5iD1Fnz8GnvQ0FvHS07PnzCD
g+F7OE0JIQ9QU8Wh8rMZ/Wit/3tS0pjMSQF5a2fmDAEoDY5ZMiNvL7NlDq3V6UY7
n3MHBb/6YIPZB1YUTgVl4tJ/BumtiVDkgW+IY0OBNDG1nPw5GMlyLEI4upKcM10j
vQUEcX+3JBr+mfNh1WAQ6DJaTF6ujZcpHPZA3OQHWVXSjZ/5oVsH2HkOgfY7kGyZ
zYRWEXxWwGcnh4unscWdk91hBJmgs81PxQXy8GtzPYIxjjRV8P2CXWBKlq1RmP5d
4M+L0b0d06a6SnIIFEIjtaP1P81pfEc29zmReNJSe0x9sRH+tXR0gvXQir/wy/Vs
2D7Zvb+6bAloyuDdLkzxhhDOc3ZeA1dvAXVZzYaXQlA2wn5p2t1Cn+oxBUy9vWOp
guYo8hUWHqz2tDPR6jaz0q+XucwRh/JQ26zTgXHo3ceeVI+/YyecmbzXCjDecYRn
QTC6GeYDSoa12cBSX6sxxqqa/azcMAc7V1LOe53d0FTDFp1MDtoZDhiGLlxUsy4e
n0LsXoM9FDZEQUedxORfWVJEwezx7dvk3tQ2kfypMgiHNAF+o28jz+BoRQl0T69h
L/hQUeWkMalenk5oC2NKTmm7N4BN9umzXUUFWLmirKfPxctJdfgezHJV+j/zLPl+
wQV0QpZ3ShKomqZ5GtVeNKhTt+oUYPAGOiSNHDvqbLEaXtQegn46/8jt0X6EdLdF
QOVZq8KIyGa5ThV9tL6msve/uU3loqwcMjVeA1c1LHTu/UtuwWZgMwSHGObsUWzA
yQS3JoEhby85i0LV8+JUXKcGKP7RzcPSsy0YXnZZby4ZhgIG4u7B7riQjjB6XPuQ
LL15yQM9qG/+IK1JQXAvQGCqu+CZow69Hn7EGT/0+u7jzepXhw9S0KPbDgB/by+t
NgiU2exgz9s5ZB+1hPZOETNEFrCWx9UMfsPogv8TPuA3wn54gocRlkBShjxUWre+
Ah7yNf21l0oA3Q4nZUowIi9dIOeXH99SaBvcGCQfXL+V388q9msA/XQFrEs8EbjY
ELVG1k3v/YDO707xNGX2u4PxxREbuugrCwVBl8NYWZbkSW+o8nzpiT991j3od0rv
i63t/xMQyh/JLyJz28z2xAXUOSdRJCAJtMct2dvMnHbBSE7dMn0QbW1NLIu69oYC
fGSXB2pRVs9Rq+Cl4xepqG3nimO9WnC1EZfNtnZ0fgT4l6ZouhgZX0aK7jHuKeAD
vk5volYg/wC1I/wqqIINgAFf11VKFPX4VpdQLJqt/ugKNKzt3Z1ULwqZ3XSYbeN5
K1b6GOc4/Oe79MpXjAEdY93X0mLwP1f6S/8oZ7jQGI3QxgGSEi8vt7oYH0sXJzqX
cvVU/F34uyUfrLeMY/+uFRwpqedZY00hQvSawvBtQaD7Kl/6jNOf4NZ/TYb7DeLT
whzjBev1Kld2fMRhfotsLmJE936GicBpzP6vRONqh3A4WLaTdb0ma+d2H9CtR7jZ
GYVj3DipyLelB0ZfHuuoE0JixLVU/PFEFvwVor+PZwCmJ/RPgpV0NvpIENS4nOd/
XD/rEBVxnbR1Dx/9WIsR+UG8Z2CXp+kSR6YCktq7a6cZ1Ua0P6WuX03/pBwCRu0O
nUqf08IqJdLwA/XUcyet19bVtoES9KnA32Dv36+KNVlIcRMHzAZNdUR7iW11VhFg
E/6wuKm4JvH4M3/I8U28yWgsBPtfL0CP8dZRV76Jj87Oh/mx3ZzCrHra/6882vk5
1t+d1im3fBcF42eXA2LcDmf0Jc7OL+V6Aa/5dhlrxJlEDKqJnlEM09vPMfUtiUXU
SYdDwKcp83jlO8Mw9E6Imu2ouzQVmQ+GaUBQInOXPfKxOJw+OWbP2oPz/F1cw3yw
hJzlo0CwwDGDYkNDMgsynIrDeKgvpVy/JfC/z1vsfCD4zWdp70aqy2/Us6vjNUqz
bk5GAKt2wEh56GY0AWed0yG64yuq99srvsp26dbzrC0uf/IftWnJT0E2YX415uLb
SctJ8I3SwAyBvjkqVBZ1A5BBtDtpOy3+JmxkK4ZZdn3K0TJLhMySFmBY9N1RcGKT
dKruzB4iQ7/7rVfw2g7ouWuqxnqVmZdjqF6GKvWejWyOKN8jKg28LD2ShShC3LR2
9E0pKgERv1IKNP3Ta1k/60Onei4xbxNWsenLKlnLj3M/0Zf2PHxww9GpbdDORWXg
66qGyYcWg6a4DPEckX1zFR+3mw9SCiCvMZ7HAbV4cKBr6wb9Oakzi8JCWB0zVFMM
BQmMMCG6GciM/DXNz1tIv7+EODkJ9Ar4hywnKeg1YAJjsC3Jb0q1QvNtFYM1EEFn
laGMlM1m2jUTqAUJkOhbDTy8YhkIFISfnl1ECA9ebml4skqubCMlS7A9WJ+dDikD
xThuUcepuT6VF6LZ2Gn6SfXmIpuK+nCX61vjeI/TBLXionf1NutCJ7mPTgKwL53/
mwnZWWff769XgLGjH5KRKTeutS282p0yyKp20h6gMMQjYg3naBEVZkAOvFHopgWO
egEGNqpU/KEfU9yR3rsUst4gsAi4f5ba0jtjNSxFuje/q3uGtFN8JIbfGJ1sEyTU
OET0uN8AAP/DyVxlENsA9EtLoC1lXQp+nygu/x/2mEmXkQihyRzO2N4I8h3RwrNU
qre3yRDy7NwKGgMXXCO2Nu/NiI8p3j2kCTHWXV0iZwrwAlJ7kYbHGRdSisC3ro1y
zelupY7GUxbG2Q0Ij7fj6ypijzcYwUT7b2cMiwq8odnS+fN1qShqMuhO4Ism/+HV
U61jtUgBDkwGskagJ+XjWhFfz7ToIAIvxUEzyngLOtUAvJnHdzTBo4UhFE1Bssf/
jlcmTsld0PZ+9lyX6eh/iUBHKQ2X7E3CpX7t3EDNbrCgIWA9wqJJuW4GH6Zn3fKY
H2/qE4AerjpWBorjRF2nLUZk2osFjuTE+VMbfnXplRJWpxJ1ttVahVXLO/iTZpvV
xqlg9kRcGUMNx0UUMRjHgsc4kgqjcYgKdkRQ0yU4wpPbUTHxTcW+A8gZp0bDEOMg
mV/GBqemN5VVj+xYxfjzKwy7Eb4QuoMwCw3TgS9OOhIgpHUL5cqrga5Ap+A63i9i
2XoEd66wxnwQmxESqLNsCt4I5SNXV9QU6UlD4Nkm7axfJyM5gChbwJ9BRRrVlKmd
ERlUQNjjzizOhyxr9qxJf8p5VWiiac6ncIf6+CyBrPBEAkF+IPlqrJ0Yh3l0WaYA
SOhg4DCj8ASgxe5gGgDLo1x1PuCm/KMl8DSz0csyjbGliPHLAgbXIaVdAkCipd+v
jYsgz9yJPIJy8Ms9f1zqM4O3753qDqUcU7x5q+HKAQMzRb/1W1mZ4jOikUYmV2PL
ikNwuskXPIcvmb+Z+9jnxNmNjIrHwSaxjB8Q0l2q02DeofPc1hqYqiXFIJRgVxDx
tbhtiDDwfdZynq37PUOcEzW8gwtRsc5Lxux2hYLzTZL0avIM2afouzT89R/zoLkS
kgDexF3XuXG7ecvtVRFfgzjmKSIap5pyLSHhA3PG0z6V8Cr2V3wzzTfo470HcBqi
FqhE7XphwHP/wBLoyUgOZTm2zFj4JrzH9DYGemo5zcQ6WRPT36vLO0YbQkxOuEbp
7nRx/ba1KzhzcJnXcNIERnUI2a6F9OckeE4gP96GIvGgNdx9MnunqhFE4TYwTgZY
j1CBBTq0Gu4tckbsFvG6c6YK9RigvDuj+jIKrrRch7JdtitwuNZLfEuAmwi3y439
nxY2C865cs3Uz6LJn5LLW1KqMw75QaQzMN+9I5lim+j7HTYEKJHS10DrVsqR/EAG
pX33LTT6YVZCtrsEDiadkZIxfzGoTrtk5Y1CdIz6LuC1C6DICQcCEpyRd8o6c9kq
6kY0gKn6/F9cBMhNUqwQyvt2/UlTXpGgDrKAEKgEOFH9HJ5Ox3uvUcZC0Hx5sM64
/WzPNo17Hpu1NhGHVcjl73rLoMXIKvqv7NLvsedWCnpJ0hGRhivMgQQXaXUCPHic
WDxIVJP3ajoLF9/5vg2trNGEDeWZ3laN9BtAzvMRhUsVV0jUE4MvnFgcJj5OKwVc
7Nm2PAKVCP2v78Ovk/Agi5YuUyTACb+9/PZeBxnK0OuAaH1BtGOhicNraaisfogI
oJktnasWyZ6w46DbTc9IGEUXySZ+WAd+6EYVaq1KsNvvSHQ4TLbedKXHEVJqzZ8x
uaQ9SWW9LSsXpH643mQHYmv+EbiSHQa2Bj+2dt7aklWCemz7nHRxNHS3bRHxmTmQ
yDV/848CBQAPoBGWjFSyG01WuktXA94apkMUXZizAVyjotywgjSlwnBhctOUCowi
LR/DEd3vsLBQJ3pYWcAac7pDd2MnkKCPflgIVW8QMAC6rah9sjAMzEmZ5rA4X2zV
7jQrx4vagc7YiIKxxtzYGarEqcxvjZkDHtWN897UObGJ/VFs91S8aDtaFHgD4vrJ
OGHg03Pu6VrrJS1yr9F9huwd5ybWCwllQ4LAV0vN7FFky2aHN3ihQfdsrgMuDShU
pm70r5efaOlTMgIoNfEGFyzp/BzYAZoUm7ID7y1b5T8EMC2JF7R0eev6KKAWnBXJ
ZfC/qTL46CGZXRrsaHEL+To+r7Pc2cPnkgA5ZKYXbygze/Oq7IZqGmllPinPJYCy
Q6CMIns8nmRtjby4Lk28TB4OqSN+R6DFGgK/e9ifGJKEKxLwKBXO8yodVKdaO+OE
0w3fnaB47GHzh4WDzFTE3VKx/64Zd0yhv+sm6bPJQGzE36N3Ms/vASkUdUDz3LH3
OhlJNTKNJrptg43T7iAg4wxzvYIry/JFlELhIEDYVQCckkqAFrfOvyG4efqiQ3MV
9qxyg/1/Wg0HNsKbK7sbAzbj5SOBV/G3U2S7VHjYoUbOJAEO33DN0iWW4qC5hShs
DJ0G3Ly92gsw3cLY7k7+HCQqzZpSzAv7f5tQY6F7risXhBsezYcnnHLYf2CerowG
0omm1RocGeKPMM5hsQaaU+7T1mYwvtduZ1QaFjB4tIHbcUkEYidzL1JqEy5vbC51
DuJCcgvtE6lVZvb3fAPePds+dvUz/NPdq6beC0IQaPshWiOyAg9wXRtmPIe6JOWy
76/dHe03MlAg8xsYLjlKGwbjczoGmL/bhQQNMksY5K69CB1cOpXZhLV70gSkCQ8i
PpRTo7LzE31UJ8POH3Nq+0JGpRMAZbOd0XSVAxwyZ2EsyWpVuol7Lr/SLUcSr7Yo
qXXQqU4MKmqjumYxcTYNu1uBiC1Vvf4queDa8VvVj3zG4C5i9QRRVwrb4vm8vTIB
eI0vAT7TCyku9gjyRgoT/4GfgYCSrQMWHI69L3hBdXrgYE+5UAhpjhkbEgCAF01m
kMc1aa5nPQhoJJNnbz2QqVMBQmHrSMMh/NAUOWZ4DvLpfrO79TwpvfigmUVh6IFP
05TfVj5Hu3/VUfOA8qBJ2MBM+Zk1Gp7vCvk/HpmjYuereZnbIV4XXoEMLPxNG53N
DcdDMJH+M6TQeH/DeR0IgDVVNq6lKO69r4E35VAgWS7jRNNeP196rPZGR3Ut6eZI
qCS3y+juTsANP2pa0e6HO73vqPKVYdtVcZlHXAvE/LeYYZsXi8bE85wOriSjRkFj
FhybBNInOxigSdn3y6v51VxGo0t7Kn2LyX41gf+hJabJXXTIx54vogJsPLWC6P8l
3MS8dgZc9VoxZH1JO2bx981ZmPKqBhu0mXrpaWJHaEbCxc6zD6ZviQKUJ7lX7NWX
VqbIAj/gxWh9LMOjr9rtoJIghdklRd8kXdZwGPM+0tjjaJ6FmZ1XP1wnAAULi5fR
D3av534p4MuXEuis3rIyFTlb0w00QAS9UcjwdytnkFho0TqOcEBdacaxBpltTtCG
4ZU2nzF0SlPZ1NfzI+ozpDyI7BhoWkRdD744NHZHccqz1WxdF9b/Z8PVwDPMmmcZ
PqLXrHSqhAc6JiJlLqlzvkJJp/va6bFTiS19arddE00n8gGooRPtpwwY6FiyaRo5
qlTWVysCg4Yc9LD9QJwKJnbXv6KeTsKBBAca79rh+Yq4Ah06h5mzrMyMTQT0Fd/x
htLcsf6TdrS1cX0KJDPmkIO8knap2J4XO18uhDdjd+jmIdlp98epAu0+osRyDOR+
k7FBAbTv6vnjLo6pJnStEAuxRGd6LqXA5gJk4NFUXEctIMqufhmn3ybsjHSwRONx
9Of7hwajssD4INykrAKjrwiBR+Rpdqbp+8QWsjX4eC669NF7GWHuOGM2oQDyX0Rj
zqIAs71DYhx+26eSSt5JS5BZvTl1GUybi/gORMiffdMMcPvImGLyoS3+wfrkxqL4
kA2ecHsraXPw8tzMjOyKDXS53isYipxccA7MMV+8p8b5BgLUVR08n2ahBW7zCjn5
TmT9dTZOKr+mk4ldW8Md6qP5neIUW7gGSt2SpOXgCu/WAlTrmE9KfvIoIiZX0KMZ
Jwcrl/nDtPWB6YiMC9E0ceskN4t6eMM2lOlic8zSO1SxjK8qH4+tshAbbCE4aP3r
GwBQR4f4StJgzVFAmDOkYwHUHr4g+JUd3xSN4mkoRBLWaO4P/OnacZbe3zK3RxTz
M0/uX4N3O/+JLInSnOY3q9i2aLW5g2/EiRxJBBQVUT89uJqKyX2p6GTjACPGg0Wz
tncbrGxlSofzI9u8uPTE4ZOQIhglDpiCa+U4hjYaKH+7FMRPM3qC4HHuLKtDr9lY
YituAWw2iH24eESfQjzF540SfS2flek0z/r/bSwXlMTsPQ8xVBkzD/cytEaJpUj2
UHLlbcC5p0gNy4/xalS/hQQOnZihk++uv0XU+yMqFQj5lVzLAEN2bG+fcFUT20hp
jP9Ca8jriLIEeF/Yp6xUtCopMvRPKOCC4sTZGF+Z67i0+c6Um8B/qunH+pIHyM1p
Ptai36cBiiFnubHiWoEPthiqOmkpGVW2xSNLyfBmaLiU9fUSOOPXELuLZB/dVVAS
zuwaSdKHx8N00+2tdDhyfng/NlhPOdNZJlAfOkJQ0CpLHKdvNZpancFyt2yl4Wu+
y+0oRdkZZ4f+DB5/7SeZffXdmW+WGDhuq6ywX3ojQjv4gflWi7c/idb7Srqb9/fG
bjoEhweaIa6Jln9++rfufzkvIs6csgrcaCW2vruZFeaJL72zBtUUlWdUVoHJ7hDt
ZgmQos/N/qam1QQ1RG3a8+Ix669Vls9qlLSsBeD8gxVeIpjKVmn3b4X2h0pRhhvx
TQN94QCfCKATXooEQ955yQnCQpId/ks4ZPUH+LPsD3xSHOBnHb/Wu4avO08klHeK
WqQDBbPO8vZgyU4Nv+VX8T0a7lrPlBgtNfSjUEJO09EJVFPygse+Agsnq5IFA+gt
lvWxVlZh9zIAqb9yRKDHLaWWrn0jEpH7tG6r+e2+sennj87gON+ciMgixrPQqGSc
wqv4v7z+yM/hbfCsrOQ1RlAPeosMJJN7NVCl4ODG2gxH9FgYVR8dQ74jhz4+8dfY
TyZLwb6eMZLN18jmFuHNXUXzJ1GiyYYzCCFCqdfVH0O1pJ8X5oFGwpSGTQu5pNry
rdxhHm1zERLe65KEcjKYU2XLChSMxnMmtDLZBKdO3WsOEF/XXRzWGOSm4DNENDK7
F8sX+agh4IKfZe3n+YY8JVF/PO/SWXz+wQCkTvQXBwFNbXx86G//Y4vJWupICADg
EUmKYGisQ7wxVHdxvGImQVUviqtHpGf0OIWX+hCpZOKQ2KHa1nmHMilad6ATsvpb
PQVymJeAXRMgMVOEVtFKR7gEsc68EvGKTGd1ndKGTLP1pZ0t1j6nDCr8Zio3DZmU
YdpLVJFhsJ3VczIQk2QID2Ezxlaa3j43Pov3hS+dO8yfE9pUFVS5rkh9nPPEfKA9
YXIRbkb8SDsnMBmTfarZ8MHxQ19DNQufLN7gfFAw8bqqcaUlOzTNXglMoGkIca5y
O5zsmGIyDIfCmJiCXu6tA4bryaj7hAZl8UZUnCQn6RyORerhczvaDQ2JBPWGV5ev
ym9NVTW73pf2UluJmfL+t3BaywFrMC1lRd9UU4zRIe9E9HswAOPI+YMjeuydHXzg
7/RxmsbjyKtDtVDahZhLt7S7oJ7Z5fm489wM8Ovanl637zc2AQ2HjeTDlgkwmIzP
nnYc5DB/Yix3eVJxLuD8B3L498Ttcqei8eLt5URbHjeNX3mG3QW4agMRg4JNtAXI
OZbsZy/VaoYAwn0DajTRoKVfCa2Ahdi32FGdHUjyTfyrSGU4RHwy3vSYlNPMGOPq
JF4DHrqfuR4mnW0MPrxQZh++o4MgoQ/xHy2OjL8nEH/MO9N4ZNgYf+5OOe15d2qt
uwMrIaFKtACYK2Sx1DxDjOgxkFLDtVg99Ni6FxS/59Rs5F70CDIntc902ijTjjct
XdGy0O/ZWER3FRuH/NUmzSBRxgp0xH0kiw6NSIZRf+TpPku7ugvE9RGm3HOUwYAU
di2q/KOLC7N97roKV87K3g0yDGPogrjefOi8lnRDAEBHetvNLPjpAlgIHxpFsh9K
uKr//9ytwEjiG84GtR0tVS9AUNvC30u/HUiVSHlnHdc/BhXYmTn1T0xz2LF8L/CB
99uAZ7kkt9lp32O77jSONEN7kc3+ijGdCY3U6RALVio5ctC9CVTJ4i4gQ7rBEPOZ
pr1xvyp9v5PducmuGPrJqAdI/11oH9SHBv8UwZJUBkZmZAtsjZUgKSBcY3AqvZvm
sjqIyW1J+rlDH5k2BymmMlE7A6nsUngSOIk1c0njCDbEZoWxkV2kWzHrE3DQMuQm
Hb0PzGh8JZ1IwXpER1z6KuPxAmi5xsKot7/MmY847EUaNSn57V9XorposyiWHrnr
mHp928rF6JLgbh03p4ReUlzepNRgZutms29hIb6Y6xECfPYIfVLDsQgUD8e1rXp0
5NTHgwoK7QgNnaJMlInGecMlIKYzaJHDfiP+oUstV/rbr/n+pMb3mKMs+yQCkmI6
jjTpCQ4OkZFlA165g9n019GmdPY1qIHlkt21bmFBBuiCioKZv7edbEPCJls6V2tt
jAfRyliQSxhyydU69+3UuiYY69nthdsrCRbuwUCuTqrI7GBYVzjBo56gb9UL1yHT
xx5bCkWdk76Ppsm/etWIWHEIhTMjJozo7ihkgJNnM8sk8FQb709+vikH+/FmRwFT
QeK7xakqkjeNQlxWEVjozKBaFTBVSA0VfvSy1tNeqBeKbEN0TEhT4UqfHmDdREwx
a8x3tdx0bOLIdx6u4mETE9oMGob9l3acL9+9gd9O2MCrmEh5eXAU04s8oCrvSfDP
J92iLJrJNpdLH1YGTPdk67v69p2BVVuEfba4ElFXZoaW4DgYb07+fVSNJ5eOWSx6
O/cH0TAO9ZOG5tqIB7MzAQDsz+JeIfI0JbJ46Yiofd0YTDQzXr4xb9eJRqvDWfDM
ViYqVEXGkAbcx25sBj7jSY+wbMTj7cUcRlCsrusoeD9Sb5lYV5bXmVb027fhsIU3
sA140I5mh6hlvFKpZwimZhGiQktmQiMFKZkEjkc7ryPsEzCAMDRixe94b1VM9kAz
odcJFQsg7dKbKBCXSvasNRpbDM42eQ/inObnxIlOdCGbs+zFpLQkM4/jpvT1+iHE
ktfCpAK+tXfR6WXZD6wC0UypiE52ETsVltPh0PqAwFF79dnsBmjyQWWbj362//QB
lzmOObbT2CHYkcruyuC+vLQJgl0memDWXBuIYoDS2gDPEOzkBYikhmKQ7A8aWpk7
V1Ez5vwhfYFisqtLrlZ0PM9kGj6AL9hBKduzs2PAoY7DrK1t7qR2qOcRmPDFeXBk
/kxumCExizSRTKLz+RTpEXMRO1J5Bp6irm41bbvGf3VXBGsANAWAITmytnEGOg75
4rRUkNImQO3BqQCQqYvQQmFiJhZgVS+gmpxK5aP7GUi7Eoue9GXF1HrMieko19X4
kJ1Y24SrRWtTJ6Pqy8zS579HhRj7zZfYoYwy2iRho4QzfcJyU4HXu80RXdQrjU0Z
gQJ64LCD0NdwB2hc9o0YSoBNd5nfFMovCJnw7WPDfcolrBBnmuIdW/gZ4KgqJbgC
UpsekqnIjwGEm6xpQVDSGA++0K8bm1miCWrOmr2T9qEeAXr/JzJf4BlWMa+BSIHs
R9ol92Jo08n78WcBzWYhaZEm9j02exxYeGsJwQOTIJ9KPu4QEtbML1AVOgWElxv1
l60/kA00PKLLewvi7n33duia1qIJOtbqK84M2esFny1Sl8/jLFx1E1LUn35IpbWW
qUgo/7cqNeQN7uQ9TGc1aC6MP5GR6/M3cYVm82kAQITOnhtshj4Gx680BftLT+TJ
0hMW9BCDvCdR1bIMdkwntcwYb+qcC3IdV+qdd4pcBDjriJeL92VjDdvaOZXkqEQx
fzt9xvgbBEfvVC1HOjkYmvP8Q75w3T6APFUDoi1kB2QCngULIJBzqRUcEKG2/YVa
SLdAZngeKz+sGwkjccSH6gYk6FH5UI/oV9C1yRSELQZqdaaIB+LQ4yrAXx5xi35M
H+R+K4KIQGVOvrXAGec+iCvRgZJpTL9oF0XEyp2XAQMlTMz5RlgOCN+2Hoj/CmJd
yJmnomPcrXt8n6VEh1up47KJVrQq6F/uGHDNYo0AzX7ubnHedMZ3OLukDKgJrWcT
K8Aqs3/0gtAsAhYI1lnXyBXxuwB6AGTa2GttOh8RQkzMa1ezklPHX0el1eDf3LJn
ieff3XY+l/V0zaNK4vt5q/G7dNJRCV1ruDuPyLIWmuL7G/BguU2H7xubsJk12ika
kJUJEBwsqsm3G/Q12UWIf8AqdbK7Q7FFxbS4qSwvzruobon3xJZPXw1QoefRDVfl
iqMl7e75Xl3vLtp3u5MW1vH9LAqYNlqQ+/jkZCfi0QSTon0Ggs80GLXZq0evb0tE
xlTp5pGpkbDxfZMSBfO7O6TiXJCmdQYcOMeYSDks6AS4lfMwbQGLVPXIAxf55/rP
P2wMPhScaeUaQSxyCkXasaqXXfbbMas8iqFeEOLG/KZ9FLcE6hoSavTJDnsgqEnn
0h1r6am5iixF8TGV/rqXJ3kdhaDf9IaADdB8Cy5Nr/VS9/uONJsPuAWUHzUCvPKo
jId1WS/6xsxZ3HDqv6r2uV1bXCdZyZ88wZtbYBEr3ij2iHR7A1cF6GRCHmnQy4pv
DCmrNcpd+1xv98wyCpUgK43EOKvt+J05daOjYktbfihtq21YbxWm1nfBH7InAIZM
hnmTXkHntJ38JPGbptbfQpxzfgt3Z0OaIxHQyRaItrXNeJPOtgtFwO2Bq5a4an+6
zkJV/eaqO09Ub5cwnZQxyJs8KAWhwfr/rHByBlAoXHKMJQ2ukbgYpKwl95ou8TU3
vw/s5tNzm860LYo2JEeYZmedjpBbIGKv5weeKRUJ4K6N+X4Nx/lqhcK47WT/F5Lr
wMfAm28yLZqECP8uzH5jKbFD1V9N/F34VseqHpZi2W0oPC/vuQXwK+WAXxsRAs32
Oq5/t+PlUnVm2iLz1ciIgokS53fPk99hFaV1ZzXLni3WuD7By+IN99TQhQrZHYAv
pWqwusjmDlk05+ul6G2SFRWE1PvtJCWa8eHbk7qXxUO0GnPibQQ+zQWhgX9uV9Va
1shCjwee+TuHRuOmUJ8x8J3TqFPFk6886TpG3Ll2BPRLdNPpnVEeflXjd0vkgJ0N
zRZ3NZMLN4sswNc6frs4RokNw+WkFmspDY3sVaavXA3F/BfwCUMu3NGk7JCJmQSh
nhDWF/0reJ5RKhwqy73nYpED8e0yE0h0l3OMkvq2T+YXH+IgMUXerfks4fxL56j0
o91BOPN36izrujjcHmMHGjw8j4vG3vRAaj7rOmCGcpPZMHFnwHCNuesS3CiYABj4
dCvgoB0Ko1CpxO+bZf6YWlDqSgn9WzHEZsVhLJOW61HZrA1Degy3Pju/imGFvcwh
ulVWK2w9Xt+fCo4Q80LMbvkFrvCNASehlNoTna/NULeqeVNhrSpy4SMcru2yv7j0
CP9tZsNS+3QbanPQRP/GG1Zeoq47/SQU6WbUqLebwHnzAtu1CnH/htmGia3dnANK
SppqH6D3Pm0yryt2WkVlvE2aNyyG3+TBMXkD649v21BRMIh7BkP+daLhv4lE529y
mQzFJEMWPg8Iq3jIt5Vbsx3zPZVHTnYI7Fp+uifI8NYziiLrHMUBTj9Glf8f6wAF
b3B3Arn4i3gQ4CYwS0gz1vzmsAPKf70lmgdIgJgHIgAxlsSn7/thcn1zmoBBfjs2
oZmZfyGYWOHP1tAEBp1uRbPajQ/eBZcev4dxW8iTETZimzQS/94rqJMn2ZnEc3D3
jRJwoXjjPeB/wwb/bA3xXNNDmJtWMPpCEatCeyzH9jrZ78uLf7J9JNCNpDXnwr1b
j3qobH7p20wXJKLLvWsV6Rygl0V2iywtv1VSn2ra126CU7dJWocxNHKbZvlxfCXb
AbngWZdGKKSGql6Eg/KdKGA9woA42qOUSFvmXFzuDW4uT3QsOSWO6nZQtETpO644
H1lRK0aiy1rv1NqAQnWde7htlstD/PWks8EdpSlrB5iShasxEGhWkwZky2O77B1O
53BOh9PRmxO7IIFllX+sIdga7mnnN4quYvOSm//wjRNTW5ARmPw6Xg7xjfUaYWG2
DW8VvbOcHMNfyudBYWEPqy6uJfcPiprWftGh797Cl7i02KS0J0jUwaK3K3313Ft+
gaSf+IZ5fdFIeHkrUf7H7y4ca/0c+x2cQM/m3yB6qN9xYdZYWNbnYNoNZ84faSaM
RXaxoeXLevPpDZ/8lAZgARaQj7T80j3CcED5ZyN1Qlyo2bb1mRkevISsYBTSGT28
MzVFUAn0bB4VK7KkAEdweI0noEKnhcuTeNSyHUCnYzM1/PXsBNGnnvv8oD+hkLNy
l+T98G0DWNTRtSYmIosHGi79YK0bcPK0dLmH4kr95NeGd62zOaQyzZmzjEJ75rio
54WnkJ9xiyK5Q/j1vwG0oWqCxwqemhRsTRzm1P0AspLOEz6sSz4FPtsosfkKiRFR
s0E+WT4LsilWosll39KXlDuRk/a9LyWrL+Zh1uc+4KSvgDdfFokSLxPRDeHqCzKX
2LnuYA/kZo4xF6pOV0cAZYK9tDCyE5hZbt+yIgdvYRgjgZO/vOzzXDFb+ZS/2Sa8
jESUlDtL75fRu6+KO4GKaxRThjbPhi+cE4XDQUFfL6yuJrXB1FPK9s9+cB5RqDwd
cRQfOymxLGX0ubS3QR++B1i4LPqBWJhrwjLSyxL4fl0ipTeOZ+eU5ZntstZmMe0H
rN4SDGzPf7G/57cpyinWlotl4vthEviaBDwuNjx5BwrU2g999o8CIgtePENXarG6
XVVwHpSITggqYYlsYIw99KFMPZAVVVPW1vMpLKEJM4x584DD8sG0pkegHBi4+JIj
kgBXl/ee1kKK8F+24hF1bDEiMK0lxOWMaANrpGR3niEe7/Bdnw2pA02+5wREbta2
mUp9Dfw6MDa2UfIQ/Scd9GUdvNVqkRIWOsllkN2vXfLi7Uu1ZjnSdBEzGlEbzLrC
2lwgI+ci8F4/0q0j+fNPWpgGDMY99qHlM/mNIUIOAak+FrFJWH7jbWWPS3CsMS4w
ItSCK4hIlTpYD9oRzcc8G05eZPSoGc0MytGsLxCK00PodSUH42QcAgYzL6eVRgmA
Ce9gSuLrwHbN9X9e5AAqrGAQQo04fUgKAIy95o/4inbYPZJaUuFzLO/k16CpZ8nZ
Hc7jjfhKsbrpJS/F6UI6EsVzYFnZrTEf45mBatrcaR0DDG2bMVkckXic+juwGeKi
GFVY1JGjqYuCZVz6fqYbzuZ0+TnUjhBWTpMbTGMfniV+Mfq26UKNhT/eK8xSZRhW
LTE7RlYWeY8Jg7w6oFEcRBcdcG7ZTZRNpYfu8Uu7l5SRlwnlcCLenpCd6u+BhOy6
p9dkX429XwjRLB8fh62qQWcNJZTT1uBAmEv+uIEf2niDrQDTnxRiIloABFC0oDws
vmYvli92oVNME6L5K9llK7ZsObZXdD2MN+2T++CfcKe/E6NWsF/myHq7ZabnrFpW
JBvG9AZ2ez20hbzTol+8Qz7kXR6v1RCTG/v57j82zn3fBcMxmO+QQzCpEu6ayfc9
KuitXuVNPgLM0NNBpv6uFWuTSqZ3EqlakoGm0WFtYeYL27XzHIeLR6UUOLtPk1kY
+NqeAcfKHWRjLuMfrMJkEJ+wc+n9hOyY+vWJ+x1TstZ4MyiiY7d3tJl3cWIA/gZW
KKwQytiIlmdK/QyA2LgHSw6mdh9/EilC4P6uVdx6ilI+5qhBND9v13WGSZo4/z9s
S8ihxwRuNCbvRRwCvrdDnsRpFxFF2a4nfU4rjA4TAY03uB4Q9kyUmSdYygIPhFqF
nUlD4tm/87n9hk+CLeoK7c5WpnbyX0J6/29k4hcq9pMV/gP8TDlC94niSev9Unce
lHUkxbpee/uKRRGzwzmmx96ZnhHA/szsZytLLbOBmH2U6R4WGA7P3hPebJyEYgpM
K837QX7560RPChzMe7L+wAAgImjGv8/B86ZKAmf/KiQAKb77uIyPnjuoIkSNc3ti
C3BKFpMa7yegiyUR6OrbUlbwjv78FGg73pQVanG3wrVvMfvWIqVzTUzNH8krO1xv
caDOoJSGWcDRjqSStZcyAZvtGXHZJ/dRkChXVSy+42HArbWO5OqQkenv4FpZldUU
0kSmaORAHRXid2dMbcfgaTf5/UeMd/Z5yIQGTX3ibJZ/ndYoSTihsSis/aCz3K+C
k7Udb1KXWWqSRZKDJRwiQzVsPY7OxkDR+aoX/TqkcTYGpEodczwySu/r8to2jR8f
q29woOFAL6HSUR9udPvzaTHXgz/O8MWNLmCTisfAq1hp+yNAZpBc6os+FPsLi6tX
Du6casWvlI+v3egIAzR92J/FSTtB2pBxT+7Eg5pessWmXyTyUojGo2dGgPKDp/NW
dsa7bRn218EpWyRLD0fd22daXKhVC651fa2auw+O+eva2+8tXjR+roNulrI8fbW+
wsv+v0c4ML5kYXBB65GgPE5jgn9QUaq2DnqI5ADGEUF6elqZbk9owiy60SZd4dP9
40OLwYOoJpCr6+y9MVMXFCtesywm4smyWC6S7aBjwuWKkHbM/kcyXMSslcp8/sTs
ehuddKkAQUkGG/bBYotTmr0iwMKB2yz4G5lj0LaNqfY9zOGwuxlGurk2rqh5/MrF
Blc2G5BiNUmhLr4C2+XqcaCsV0wr5ycfGjyHSUP5+9AAZV+o2o1fc+zsABBfrqPx
YWOYpI4W6F3szgYxgA3R+eJtU+VaVZF7xLDA2moPZXXZpqpeVyGkBBOPlrVzA8QZ
tB3hj9Y6iUSl0j3AgVjcDoJHsddSMbS+NOmf8kO9W3Vme8x0VHC/FIW56OxXLN4B
H7NfEDD5Ca2FHmNYXYA/qlXFF+a+dpWI5z9prq63KoG45snKBk+YuIStQ8KHQxJ6
S20mEfqPZNTesCnOUgUpP6zRnONnpa/DJDQV1XVTX5nwFlVYqH8aA6M172n49PQD
FyMtNl1vv1R6a6iVSQjizMLk3LvcaxTx8R/8i+6OeFRdL9Az5SzWwZ0XeQcWhEzj
TxS4e5OoqtxLbbtBokUAgt+eAky3H/W+7gT+s/vt745lh+AtTVyr4feeXXG6L/An
rRoemLs6MVfGFlCIt/whdB9jsznstp4hFjI0B1fQ/FEwSNiKCaG6/ZfSKpO7ipJ/
/Euei101xBC1Z7iKptD7uergjzgiCDpIV7BQkFvnNN/EqIYqMYso0elFOjPOjoz8
QOrGQYmQYVuoVygSZi8TusOi8ER7/4QvwXEkvy831P7OQKMEghGr7UBlGZEVHBvg
CkArMFmtWJprXkhKrxHNYCkivy2FHJnge/u6oF+I8bJWcoUCHbfW1kowti4BXXGn
Jje6b9z67T6YkEsM2tE8hpC15Quk/iH9LujBZA5dUd8CSqWiZoxQCoRvnaFgIPgy
QkQkykTehjt9tgsMNXWHK6E/Y+iTcegdvIVkGlwEeYMRz9lYJI3ZjaB1uKzgVfMy
MeAzVt24fjqhtV/gzhDmXPLJvFqx34RI1F2VK03pxA2PsL2mNd17Syp7FXfT0jhN
cWRta/XBXTDt4qhrPFv3GAhyskuZfArFrd6DBFJf8L+NQtgRVsIkNRl0kdIdt88w
VIBogomVyBSFHn6SBYdmiYazLZKdyZtXZve78f4ns10g0owqytzYYOEvCgd+25j2
1TFxQirkm+UDDJS+8L4wOwKIijR6G5u2Fa9ZkP1Z0+efgovOHMJwHPFQsOtGvR8u
vDQ21L5oCJKOK+C0u9+IbXxmpk31x5E92blL6Bpt48FB/FwjOW//T/XTirWVbM8H
uD7Lo4umnWZ7z79E6sy9nfpwBAFaDQxAlMfE/luHcj1CW305wRzZDy5n21IuNWnt
dzT70U2Qgnn60o7PNkfA9Z6ovL+tWsh3HBHzY4R43f9UJj2oEWWR9KWAPFjbPJb/
K39/S32Ms6zHHddWFv34NnNDqNIZS0zynbIx9gJVvAWdUZP9VdPYTfntoOkp0MGN
maG3GvKTdyMjhDkoinr0KTbU6hgnVruz+DhA/3LBbM5ogElmwbzLdxHfMMug+ILl
uQBOt+Pbh6YhVpVOnt6qVHD6hP6j63UMw9Pvw/eTlTZ9dXuMASN+oCcPbiJ7KW8g
cHs5IcmiETdXXsUb19+v44qRZC555mfxcBkTCta4a19DcWbtkgQVsya+a0UPklHE
ESshO8HBHvqYwWdgVAR4LkVrvd5Y/zAJ+u8F5csvotpXcDqU0gZHfLGoWVCYkG7S
Ugqj1YmAvhadWLySh/niEN39Ze25fXtqdety1qsYUsM30SCkRKZtl7ntaaQzA4n5
7r0vBZZPZ0wD5eiGJgBbf3m7WidsAP075Y429gWwt6/XWpSQ5VIlVES/OgYJxaBR
Ra9yfb2quJKYSp110PM3H1gsK4BA1RgNFfFD6CQNRCSlkvG25Xh/qnGJRt417a2G
gMW1cuoKs6F9LZmCNxeoXiWoBmq3xCPhw3vgDUA+q+KiRiWLEf3/697DsJICzugQ
RIFbZK4EwPtXez4WNxXzPpaRrhonLdj34p+CghK2Lod4uOo1xghmmUbIiFuNteX3
wPhr5TSMA5VhSICWcLcc6NKH2jBeGYc0oCCxBb7FtTrmwZX3l+2fVmkrX9U0278n
hJmIUh44unmKC7OSYQ5ZrcB+N7axi/TFCYC1Dgz21jrkqNlt7G7F6/SpARzX5Gel
WeuyOshR8WsvKs8Gk8FKQwK6vAmbUAWJG7O00T2+eWs3hfbpScAX2iV1mBNMDyhP
1J9GYt1Aaaofxmzf6zdYyCtJ09VdQt+tMoYkv+eo6kwiddq1StRszFVa/PlO1lVt
F2TRjHLPtutW5RxQ4L81yhGln5G4Rf7d2a0Y0f/DCumB9SiTRAHnMVW8viVmLyEd
SAc6t8H79k4xJVxh7ZsxU1OR8n0s9BhD0ZYRjpBP5r8+Fxu1siB3XMgHcmbki/Ly
sNQcbpXblhWlVlAdCCME2zuEecqWyy/tFcPfIaI771HDhwNwXYZ4ZD0ofDdcaAk8
AkLeChl7U9ZtyWafBxeBrPwf+JBmE0Wxd4j5Fc2ciPQ4eMrGh3/oTojXh0LweB6R
34QtJzr+awAWlKd0sibGnoRP+K8kvrOnD/OGQ9bTHIE4GYgPYI9U4wHqCGwz0Ate
f9aS7KpCJ3HvYrWM2ZCo/WZsP1s7m8hdjx2TxUL+MJNqGHyi+bDLOTOHQy5TAd1j
z+g5HLMR94ili+7zMhkv5Tmdktmzxj/KeJv4KG1aMEjG9Rc+S7U9UYw/y/G9igQq
0VlwCjKe/K8IY/FK2hInX4hmnqtUzCsJcwwpt9lEVWtCyIjtIFGDP4cAAL04ZXgC
Z2NvYFRnGwRX2NaqBaYy64arwGWF7hTXkf+WlexGYr1EY5+SfIWHWBjjIM1Olmew
POFsCXRNe3am27gGFm8TW4o4VIAjrZ6W5TzYD4NsAnpEsnCspX9YWuBjhTYSe8gt
i4vaVcMEzVu/15HWJ83jwN/fGxl6Az/RPfuKwuCipHUg3UzOFHdX8IzoVJs+U0IS
YYZ82tkXvkJIvZItOLI6DGKi+8hSA7ek2MIAcoYrdvO7t1AT8bxe28T+tQ1rC58P
EBg8nEv678nkooAxleahZVp4Slgh7fs0FW98OEN3ERShQlO0L979cQYyuY13LT5N
c0PhiI+37ZZjhfX/zIO6bd3tdL1TWJtWW2DVT59OGJ44aPkHUEWAuFRaZ2wqvOsD
wV69yrHc3AV+0YmOSjHt/9RvtDy5xPijXR2YYn7gOb923nvmSJ+wnhFpDn2AFtDr
elcEIzdXDtXxH9WJJG6Jb6SY+dFPxw2gl0ip9Ff6GsRI330EhLpTr9eLK7gU/yia
VyKmzlHNp3BsWGrGqhpkcWVF8lSDYuD4pGMylcw2n1sJGCLERhWueg4nFJIgLsfg
0ABtAiI9r3SKJmjmI2ZAhwHBmjQzh2uy00ITxYQwFX20cWF6Rh0iQGB6Y95B1hJf
YvihR+dPqijdsqwNjy6ic8kEK6hPCOgM4F3QriMLdjjxIbMvQFycGwk+2TnsAlje
GjOmOjdAHHMqkwlsog3f4aMPHlLkNoTfrzCC+eKcOLhD9sS9QMgcvaRmXyiBf0lf
Q+ZbeB4hy0un6HwgLC7ybefrEZMrx15bAptrwsOJfrkLgzziQHOf30o+p1RCVPbO
4ia3Bi3wSlnaU5RztcwfgAnKJjAd40FZ+P8GFKNXOqbgQXJR5s0K3Ej64JBwpKfd
Rw+7Yrng0FzWRFnvdhvrdFqcycCuDXcAJVHjbUTSW1Hok8h1TAWlsMATvLCZ40Ik
9qCuRTD2r9CZ7JouDET1xZSyUjsc8tgMDFRLrizyqXf2wd+xfZqm4v2U9nnm8p4u
Adeb2Pz5PrJ3rLwO0UeGeLItk7XV1rt2nZaUBIlsnJZmMKFvRjU6cTs9O306RxAY
q7CDxmbJCSETJ6pNyE428v38DIU3CzrPnHcgP+FiJiXNiOs2lplqQf+GeBWhVAZa
UypbYDHPRu0P9kU6pCEuEKoaFpUOp0g+0gb7MumyVF4fYHENjUwfqC9jlkUVVSde
M/J4tG4DjrGMJw538CYZiJXkXLvYJVtc2RVqzcku43ETrwCYOpRDYFdJfRiIXNYj
HoztVWma8YXI48lD5/o1a5SpdKUUeNC9JCax6U68AoZPgyKudomEHGgNhH3VcELa
qwCXiM4Yso3HBomMOS1VMHXZpN7uoCELiBCCNZijvyZjuAm/6NzM1M0aQcLfNlls
uPRWEOPBpn2aRgssPcVSOq7fu8D2pAcLB+dIUu8Fcyn0+37jRXkI5SQFpfe8+1pJ
KeCJI8PXYGhl0ELNEgLNrQz0cRAm0IM+al9Ubitrh7OYxwym+Y2sflnkH0AJF032
U3iZ1wa3gtAVmKZiEnVEY2ESTsMF168WMYL4u3pBbESwKwCnjd6aSXB1Zjf7L1L7
fak3uOxKrKqxNlE1/l9EwWUJWMzhw+aENKJaPLkO7m4cEBRthmhRDGkkQDzYuhgI
J5lHVtMsTFADgybE4yGQczRj43+KixQvOpHRaLloJNTihtEeN7n2LGZFYV2OCdEJ
esldxEc6Wv5Cy/RlsVWzSPH4CHzfZvhtejsvDyeQMSufoLY0pL8aqnaugxaVgB7J
cwjT8x+Vc1Buz3mNSonQPTgkQ6EcVOrZF0x2rFhmC5yJqic2W14qsmodUit3qWX2
j/zhi3+ugwAO1hQlXhUJcl9ZDXzsEFeAEam0UoJMQuMJLuY8v8xJQ7xizSsda1TW
75PuN/Ad0LPGdvr2yTZvQC5OZyEx0VnIrxd7Cy1P2JPFoFzSQO4e8xZyw8NWU+bt
DCgMc+f9sRx8Upntk6iGZKcHTG1f1A9aeNf+hnmsCT/xWhB0RI+RE7KSr+h5zIiX
jlZEe+7nYXSx2yfiukONRzbTrKYu0coJIPzoouQ0XtFOYeERGphVVunqpmLTYp1d
WZyLP2/Q9TOx8ZbGbGT37wCsoOW7KK7c00S1UR6Cm+EtgmG6W3rzX33rwL6cFnJ2
bzeJCnYx8MN/LRXeq9wzXXud3lrQFS/WWjYOP6HfSC+7BMhmi2osfbv8YpwL/Vcg
vRBvJrzfncQCwWKdFZOUT+9S6tCIU7mS/lf8Qufj8a/1f7qxW8K/3393Co5ap/7q
/ZJDl6lsOxnYpTkkcSxHr/wggAqAfNNGk5Bq80lqytoDqLCOPIkQCePwenLP5eAw
iy+S7OD0wg7CQrtcpgLUD3X6cOkeFP5o1Ogde/pohoaO3JV2fqJfClbzNeADojpa
71MCG6zQLgHVyuSZ2gGSPpQn0PXEHetrX/cUCABOkz6yi5qJQEbOR2VyEzzufm5f
DamZzfk8xIf/W2EoUbE60WjX6SZmkW41fb5+6FURETEgxqTR7q+xUWqPq7vU3Bjx
2mcc0AlCK1LIMJv+qaUHs2eURiDlHKQAQjrJnTv9k/8pfb9yKWMn4KUI9wQRoIIq
GrYc1pvLHT+E1yEOS8We+z0qeZA9VDybqpuCKkRrMtD/3NCBEJksZ7y1aEe5Owvt
Iev5NCcomFwk8MoVWhKvXkRmKgbS1M6M80W8JFgK3Mmg4XGhD4kUFPYJcCYgWNND
EQLENFzjeqi2BEO22ejKtVfBCsh5UAp7SOED1+z1004AyacMeSO+We+ws2i407+n
UxX+sOhn8XYkQPnhOCKsw2cR8DAjqNtSUHU5qtRg8oQNCJirYvHsdOg8WqkPNfnU
YIK2trRKvX5nyJVWFCx59Tey2d7UW9jY/G7eJuQ+15viC3I02/Xo+Z/xeE8qG37F
VzwcfyO1wuzjjgThvBnjtaI4P5Gas2fHqzEwLlEMnRruBWxD3DDBihTXL+vbSCdC
W6/iUXcINjHbYsW7GABaOk3WJXdBWAcMfM4ncEQUbto+uAsLcnsPCPFtroWilqN8
XlDsH/xrgTaw25sWPJRu1q6gdVcFbBq7eSGqkQDBgsByjPawRvXFUj5xnhRLc3BZ
O1JPD3PyRZEu6rd8hDBZvV6CCX4yaLVYc5xtRjWQ7crYUBFPtZfwFh/XrJ2KWc+X
P85ByIF9uXH6Es/+z4X/55/PqCq47U6Muwv+apd8NfnhtEyuve4XUM5JLLtFI9qG
e10GpeJX6gvdyozlGfMSXtTNDRdNeTU1Mv1wkWymRZsh9TpB8a09IM5s5/ufkn3L
RaE8WH2v4Xy1mki2JDFwQBtoOQ32tchuUDg8ed+O5LNfHs17hivX2po1Mwt3MF//
4qPnMT211VqSEl9AffOKZtRM86N54ZHLdLzS9IQidImkRO89ujdE9YRF40xmAIE+
1mjRlFB1LjPk2kWpHYD7NDv5Ph6mQyx6R+uF1gYIFpGCahSSzJmHsLNCGpgPAooV
HfM3Ok7nFzhGN/dvFjuJSb5GJYBBAad8NevS4Fc1l2rUsCJCPI6INk+1Rq7489bL
8WB6DcIhQq+jRj9wrhs75BGX7rpg4/uvFpjyyPlIoBIGcC74Cz7BowM/yHrsTHCe
FMFMJ/3r6vaz4w41DuHpAKESN3uN5Ps0FAn5P+ISCc0dz8N8rYREugIeTVAoZl++
1KolskXfZx/3XsLtCkXFy1/ueZDrZAHyrPWjfhbkLLmekCUDkA714CI/6zPa2ZCR
kmORzJ8Isdrw3SKBeEBmwSZGq8kBR3Dv8e9ZVtGpn/JvqDZB3KcSdBkTIoztDTjV
1yWlvIxKeAKzFfW8l21tKOEX/ObtrOuqbRWNIetT9X7jvLR/HqwYXvGLBNeG8SBI
fc9ABrb885hyIpgo2NrqDtmsTMRAd4u5wqXYQcEJ++rAdr+xsXSDkAPLY7xSZGh+
WTweYvyaTqVt10DPxJJAbLIC/QvQ7bxm257APwzaG9LIw6IAA76PFMZ8Mdo7DTtt
7FoxuoYLoBa648MGhLtST2wgDaTJJwOxg104bU7T++cGIDNEPaf60THUjn6jVkXC
9mmpY+ikyuKOROWw6WUuwLk446o3IV/sZLGUq0KZ7lAegnAfGm/fV80mrpCnplJb
6qWn6gwVPbf++jKwnIYu51dtVfv3MtIgKDe5Pk15DUkjporXDM2oCVp8SKQMR0/4
AOcZjT27fNsuA32KoMREQH8lXxQRZ0RvW7UdfJhshcrqszlnRHiwzuOCMfl3EwM6
JKwbNFsERPmTWG5GHF0PT07EEDJtntFi3pVguqgGG+zL/bFHIpbrMHLvjJHVTivS
DwjMsKgYV7aBg/wK/ian1rwi/YaNnAEafayYMCYqe07wKKmSH2k08oqK1Og+hxyw
EzleTPKwBllJ78Q4t0Dnh6Pw3jG+m3jYbnbMNUZ9oHQplrhAh3f0uG26EyzX9b1C
RatmoGK9dB2RxcFfhwwREETKtD7zQSknXMDgJGe/+AJVCzr2JwmW4wr0Wzp5vc5g
bO+d1xpVE7rfskCvmtsho6IkITCioGMI25dV2oiN845Zd+1M1rRenBhOFFaXgEcl
foQ544zcUAxgdvXxhLex3iO8uLrv/oq8h8wf3++JQbr5ZEHArVyC5A/2KcuBKJMK
G4j1jt1hvS1ALUKX6ptD8suvQpbMARJ55yxdaBaBb4zhgPTrADboLmC9j0NdWFDy
95kAgrOIxXaBvxfC2H0XVhARn3DlE8jEZI9fIQyygLCrNPIOy9HnxLmPjurGxdWF
vk3TtaKns+kd0Q88xaTk0gnU9u3FUMynYMLTqBdQ+7RxvMr7vIT8eJT3FRTG5l1J
p4zlyc2EjKTee7d9HR5T7QuGoVB77pdbUOnee2RbhEa4ueoNMB9UCHkAuOIVe/KF
YjMQy90o5KURyzPnV3KPPIQIV8GlnLmxnHmeEwPyFyAl/PS+CAXW4d+Lr2Ag/+ST
pPz/WSs2H7TLzQWCHHVbW+3uSW4Nm/JjXnIiwOO/zLnfpCoGCpnmeZ0Sx5Oc0pv+
QXZ0Y413LhWRudqXfCqZR4ohfDjxpFsrdR4h6ZxOUr0TyPVZ2grKrf54f5I+Zt23
A6T6XnhvpVQckJ5qY/z9FnWsSsxq3+wcjmWPNFsnjUKhsb3DAmojf0etunv9NpMN
FZh6TWncwC81fLLULSVtS0Zrn0Odv1iibRCNhniqsI2vTn00/QVPdi6iG9xqrGZy
JCDaalL1cm8Q90IVgTivjPmjHboWjKBvw3uJMij8Hbl6p7pIucHWXPzCAn/SAVjx
vWeeHyY6go4KGD8t62JzwDQrF0CcaM1Nl6KU9DkdhINBgJwHzpCnKgzTWEtJM/6V
Z256wg03dsgCX57uEuq4IlWbpyQD8dBh8AU/NNiFG5lYrJc86vZLYjUDrYy76kfh
P3I1cyq1REfLGGAOq1QJSXUPxDASLoEAvCOKsiQmhUqA5ZCt2M07nRRGQVBQmCpT
teGnC2JlRxJXsEH7HBod7OFR5Q5Aeof77cvndmBGMePf8D4lEAa/pI4M5eNPmZLI
p/4HNl+x0ZWoE1ezIfbBAQE1oQuMyvgelyAWFfMtWaeZ8k0Y9ffiz4fSJJELaoH7
IvQzemI52N3FzdEatH4vca0gBReMETOHupb7GE2Uib7p6UsWPxs3tNw5HpB7CqgE
VPwdKGKMG4hqBtgRAw9aNPnwWt4MSRkmMVDxZlTYsC4zGkD+jOsTSVLj3y1+llvt
Hilsmo/q8JonzSwuyS1LylvyzHdcpMOgT60PK2gtB+hclIPKUIkYOB4PFCn4Ly9V
rG8RPzxj/EfVrJDfQECMbYbuY8LVecHXlOQ/mi9yJYqee62PCvybJj/+Kl5FySAs
X83Xacmz8f0qPqrEI4+bqiPftiK7t5OjvZpMXd60NHnouhyrm16r4cOKCY1xBcMU
mb8Ss+M6fYz6F5iVZb9BZg5owqCCIcemQ2vgz0400VnO4eRxps8bZMiS7ISoam+L
2I0qqVMfgPW8zRevHQI4eZve7MGmvPX315BD1ABnDzRMaghAYuPd2XyfT1HUvgnW
ilOLi1h8+4KZkyLXFy0sskkQ6CHR5uXugoMyd60wV43oOZ023IWKehNZu9xR1ZZ5
n2MVAfpW3x4nh3hOMELJnteJl8QJ7F3IrhhyHDlTHRemmVDu3eYQt+jnfePEC2N9
0dTh85suhjXdFpsv9yUb8+8aB2g1GmbRYIt+4/YHkjmi0a1fbtvgMCz6dttr4SYF
Ckkc4UEU3f7f+ZQwWjgkOANFfjD3XU4JVvWhx87lqDYXd0dRFw70tHXq7Q1oQxvO
Dirs+S5JB0VMkVt1gxvuPHf3lGMsb11W3EWFBIvYGCG80NfrZWb1w23O0LwSCMGU
z4YKjqYv8bBC1aBpjIkqed59hpw/4GmTBMl8pgQvNtljrwvIPjokclmZDaQGu8QN
NYC8DcBjsHbNVAJeMyfU/rWAGr0hmJu0f6T12+NB/dVcNfvMpuySbSO4/ADbLXQ3
FyYlfWQiyzdVRZJCdZtFNuSSFZtkkuD+esgLXpInOBZtojp1S01i5lOE7yL0dwoR
wLV8BEdS/w68bn9ZhcI/cJQoSJ3Fw7QGNJ1Wh9ty+prUnjuma8EC7GtL/B9tMo5M
EiesmBhw9eNu7SVJztInY8gqiddtnMhjk+r/Eoi0mbsz5t5zx3ZqREp9dwu8gvyC
Uh3t6vNaKxaI9Ywa4WSAD5alN2PdpYbEZYbn0xZWWgSrYat3NLi7G68ychYCtamw
/oDZjMGY+kxRtXHLyphY1Ooo4iHndYVJorGEBfIjSnz3IIWqn/RfaNUVbz53dWr4
2JKAzPgGdAI+MCciO188PZvBdP/cJaCWj5xsDWh/PL3WP6NKWEra53Y2QTCBP/BK
r45wb7lp3PDg9jwye3C0VX/a0ipMMYvRRBp+l77R2WS0qLmJXxJQH0rFgIOa3loA
IOTU4TcVZrHRJPBtSrncs35eH+ee7tUB/98vZh0GeMgVtDbmwRQVTkDBHh7qVQ9c
xduqTi81L+LpEJlgtQN9L61mKy3Dgy4jfBjZjwWhWRekL7wnC7mIWvtO2gFMHzPC
jlln9/ZMyWL3C3couMxdf1XTIA1lAMaH1em1pbI1kAmb75egChUbLhIKQ/HLXOlI
1OxjcisMT+chE+49oNP4WubxW/5P6kYuqJfdFsjDNHzxkrz64sZgipvU/daFgb21
KwmA9pe5F9o+Nm9KrNZMb9c2DfXTqHF1cGKU9+YhGIk0J3E+GHpbYjk8qIUrosXI
JAfhfZ3ljas4IzDE0LDspC7TXhWAAHvccpfuuB7BebZHe6cg9NuPGhmKYN4mp7fv
05tJ1d9LHs0rVi0s+46cv55Mt+QgOh6nQOnHSaUMXb4X9Fjk+Pxei/k2b0dYTkK9
vcUTHgAZDnKQ6fzNtWXGlwMGXqWxcvDv9ytwskGyGTGUoKzK+g5ripcx2cu8zQ6U
1xXwhYo/nec4lC8ekSYZdho0Ax6jXipTQ75eQ+Cl/FDBwR1PsanGsr0xy5qOIXB2
4kKNR8SeiCe0xk46sIBX9JmOJLEzebOHkp1JYxwb+d1ZaKlHUWwGvdA9j1oeedhN
dNOswroCvLZhXTSLl4JfWu6EaRTPDupoyzjtzGr4n3ycEFyacYQurljhfAciq5yc
O6Sq5vxQ2QYQgoC7t1fkVkBztpy4IJENwhrEPzPl4MaDvx0BgaDQpwnhO7Uizqeg
pyMy5LiFRlc4E8uED1kQ09D5nNbdp+XcWFjANsuk2PQ6AhV34AYL9Ek3UzlJg0k3
PE8XJvu9K7o5jdwLw22Z5KsdTEZyzu13iEk3cWUF1iNtnHJvKms7RDF5KvnRuv3v
JBDEsbAxImXMPvw+hQ5bc0JADB2FrZltluhqQid2iSMeHWYVYgAbCECh6WC49UUl
G/ijgl078JoePTESA5B9RQvmD21I1Vc+ONoK3ApbIyUu2TbNFaWMxm0XO6xtSXkI
V5JxSNN4QYBxL8eZ4ugGkUb1xrIHINO+1SzGEg6xr3EUsCV/i6sh9fBCZ62b3jdX
dMHqLL9wnXGsWesmwLJwyyFn++NwJfivH4pqtZERwcABl5la50rDxXYZPOsLwQlL
gWop0xGaFrXKzfnFGej7bKLOG9I91BkMvALRhTmHyX8O9+fXk4XP8E+PXFVcKpU8
4Gh5N4WnPT1MymhapW5Kmvx6tBwoOiB98KR4sD3JxWrX3aJGg1eCARgQRtk3jmma
jU9eRJmGniyMI/4OzBjivG4xxHqa2w7s2UxphKxrCFzcrxtE6Ny39Wio/Ka21x49
yTW8NpR6NZbdXl9xJZaQ3IJHAw5fbNbxBdGjdgbqkxY=
`protect end_protected