`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5744 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
LfLaKOw3utJqtz02pVdKf2SIZXmC7ZNdD17pU3lAS6gCwhGXvHb3rmlv7+YM0SAx
O9CUWp93iNUj7pz/pVlIIOkT/S8F8p+dMPSmVWDjZy65IpETrRPP/WcojYXMYlqz
XLiAySrt+F7hKB/64HPcxIHa2n+FiB1WZ9Z3b66JrScdaCQad93a3nSFCrZVhqLe
igKF1p8dBAPBz/gcdD+8BhEXHADpqIk5yyTY2khdrTpn0nsgmP8+6y8V9Zdw633g
MbPQNoQQ2ysMjfgBdCC1OSJ+waUZ7qijJ5FVY4kAIwZQa8cm6dvh9iTg03xzpT6K
GKNCjTGs5lE3cP+8bGADeyg5nfbspUGnUDaZZxBqA4qF8EOcLk8AWc1ckGaXlhC8
10qIE0qElL4TV4kaYCeNiEVT2FqzTbqVG2WARpnLqXJwK8psvLNO0y1Q+iY3E9lt
bMgDsgKwtVKk7aFyzw3t8IQnP1Orvzkm7dQox32Qkaqsp0UoyN5xudNaDTAfJL2W
kPnueTuCJCbscUrccR0G0pRTmckLj9Fu65orPWd6Z4VAlLzVPWZTFAmRa2XVBC6o
0A0fZzFH8Y1GBUTDzUmSjCZfd8J/9bPgTlU5H31uHyUg890Di06AcfZG8RioTW7L
3KghjVFBg25EZP3Mp/AjyeMX0/Q+uUrsCelhrEES7Z0LPrfvtgkwKL7kh9mtS9+p
dxC6CRn5PRN3uPN0rA3M9VDZwJTztpTPWHC95GBeFPrjhNXIP8XMMHU+nyXD7cnx
m/j26cN0oI7yeGTQBC1v3ES49bWq6NQwZrYkManNB5gOCIPtS8NFE11mlwWghyU2
Io5pYS5vZjUXndoTe0PF0rv43Yo54CkDwXJQrK9tbi7sPRnWXSRf8pUMEZ9n4Bij
8KAh1lxBpImWCUTpEl0LLiVV7gamhnqFuGGAN48HXR0WUtlX24NczowVBEIJrJQI
O6qExP+HBZewB1HVhYE2SqcN9dM9ruPopclOe7HQy7KkdDvTs8LFSp/YTKjBBFOK
660hVtkMVci2TLBer+EAYtZnyVWgy+VrR5w3tXWmVVE2QnnCifYeJQpkorb9Nc05
TXbUIL+9RILvdhoHJfHmBRHi+KtBXU4ZFGfsaCSaZYnz1477f10Z0FW2AZLVh5U6
dmfRLUa1qbZg806wSytpWD5Q5Er6aN0gQpLpQh6bVg8uQUVhRCRj44C2rpdmzUZK
BxcKawifivnglcr8DkDaRUACz0pth3J1bbll0fTT25EWfWOr8wWTmnPQg7SHlmhZ
3tbthu8WiDWOXnftelm3KbS5kUiL5fDUZczSPeMIJNB2EcImqfGtA0YIvgclZqUT
3KI5ERY2ZkoFsTjmo3BizsTvcYZKT3RHMNDCO+KZShNawDSegCLH5YjXVnu3V+vs
5ASWrhS5HjCZNW793xi0Rhx5+8vys95hw8ILwyP66CbM5ldRP24OtvlRudK0+PsA
UIuaTzhUTif1dhL6TJm8R5RkoyYzfyOdjXUeIkYUEbHUJKMln85EG9Y4MbtWRbX/
LIcJQrHOazhR/XajUF6EkmQAXAlD/gM3Uvq5owF6IFDfphCTSk6/4mebIhDlr60/
nitWnXCHMLrfCrlmadMOq35LZbTUvARShxmeVuC0tBZdrUzr9MXesylNKUVKMIW3
D9d1lNsA/UFt4w9+2/XKsyo9/wban/DzJp8gI3yrIJTj/xKKQf/Su/xyyTFxdBx7
n9LA7fz++m/FUyzn0wGtpHvOOmbSoDVvCJTugY9r0UpuhIRLRzb6IB4YrWkfCukY
olwXXpBlFz0wdwYMiCRqfBoqX151J1XVb0CL+dlMndUwhLBvZpGbUGWRb+OO4tlC
mwhBLQtaIM+oglYaXlJKZfMvlpDF88+0hwzyf6whAEbE0faqo4nUmNdCtXwqlOc6
ADmHR7thIvJWlzAGHIKW+TvRIkvalBHlN0XdDZzrIKmG5AbNAzVa7z8hEKPyp99v
FL1AN165qOPx5EbUPpy5JrS18RgZHLatZPXjL54TqKTMS7djbOFfLOCxj3HId+wj
Mdpm+2JpT0J2yEqy91urEtqzM4lZKsE+wsjxSWWZB7+/wez50rsGFCvqz8itXTS0
wdo0XK8MasPV8y0iA2azLvFvx6N3IyVFKEf0CAMjgCPzLBxdRGtnSEkGizmrOaEl
nD6NUQKOzJ5uBt+4xwQKXBxAwpvxbjZCoP6NQvAMTOV0X2hkklZn/FL4cgHUwX6t
Q3n/AHiguWJzBRgBNg8wCpE+5Gyy5w48vqWy3N9C4qV1WIjEYwL6IaduOOn3grnr
UF/8V2RhM+Ug7iMp64jTSYc2KHqiyD/g4+tOhPqEDVnFUclodSpo14qWSnHmE8yU
PfudqMht/BAezbcgi2KdQqugRy5kd+nNgsnfjtJPEpDvY61ZwMswaUotwjMdE6rQ
Z19PidAsSvPC9FXo3LPBfymVMTWBT51XybQ0fnlnM8dt0AdL8YpkiV98y5fCP7P1
2tegwhaIuPT+joqd8fB2a1gOBPLDmS+TPHtPnghJJNz1LUurcGYUUw19lI9do2dW
LtFbfUcK4ioygE5HKfoK+ELQ+4NaTuIQfwxYtXi2r+uo9N1KqWqDXw4D7NdxR68f
7Dlu/2WcqUAyocnC5Td9Jt9TlMwlHsdI+xxMAFRdI/Ge6HmWhszFRSj1FbRV/cQE
lhI8NDjk+djKHgncYWK9wPIS+2UlXSd3n3OMvOfW3jJXjHVAQRDU6/xcW5Nym64t
W511/PWre3ByOrSlA/0DIXYtEf2NjUTGLFR0TuGXqkV1TkugUOsnQlrARhcBWA+X
vweXRu+G/gyg2bYB6/008t0braF09v0Uhf9C1r29zg1BfFuQMSXpj8/VHjiwNx/E
PGultDWzF1Oq6eITiqEmJyKWGpoglnrSWaREYTGGJMeaMHVGrBYkNHZEpi1z1vZE
bcaIQYB9qn+EC61+mGrAvsFGsc1Rt8ZdQdAXKYoVjM2PxQ6KqibOugGYvxlWJ/M9
5jrR45GBWpIieS47XliT7CtCKq5yieqDEP9efBVAAWjdqVzMnKDf7/FX85nsIqws
0/6ycTdCGAmMoN+XhRnS2M2lTQTUBPpTE+X03J7a5ClT9OL2Q1Av/UUivUgM49lx
67Tu6xSRFWl5s4CTL80D4y4uheNuYe5BJk0+aV2f9jGV+JRSlTZQ54kCX3WKFMS1
EbyNn/FV+ggP0kcskJteguGcIpIfjlFWfdcmkCf85m+pH9sT0ddAkbUUmuB6ISfK
L+OdBfJOISnUvLAen5SmaM+FGiTeTXD4Fi0e8saPSaV3IatSGFRbPRBSccea7gGS
kW8NARwNflRh7u2l6YNcdRbdMH0yTB00hZIV/BMZQ/ory8+7aYJtrg5oj0SQroM4
JJn//yBdBBFxDELy36F3CxVaZQ0gTBxU6az+oEiLb+3W2uvMZH4KsejkkcoGIqC0
h12hQ24TCo7hXLfLllG/DPSwJy3sXFX+P27LkPp1/5zfu8U+NZmTzLbdwbcikBvb
OsdmPuvmnQTxh0FZvAwRuuXIsfyDOan55BGWs1O+aq3T3t3SHUWtHjydBprwG4i/
BBxMlT3pkMj/RTyX2xbIfONL6ldAz4HeLuAmXIth59736KgTv9lX/PgSggaGeK+S
63WgH2itJlcTPSBS8pMOcSEvP6eOHOpa225t0W9mc8cqyR6NIKy3B4eo5E/MK/r6
bGyuf6uTGb7NpeDn15z6ZmdhHdxikxVMOpoOfGltzh/DkPvfvZs0Cvip4Z18pOoN
5sToJxbzSnmtH855u1s2yqqQi9ZwvxiXcyjVi1Ms1NWSKhdK3eNjl/HvXT7BgiPG
z+y8IOOp3cCg0aUnfquMaqZt4w7Ifl95pIPUMY2DZ3QOpySD5q/Q560pzUj+o+Hk
01agteNMsnzznSQYi9HbzEwBtElzuOm8IuNCa4nLxGMVbiH3CKk156OMmDfash03
7zF0XiX069Ud3wsdEGLjOr7Rs3TL/u9tkyH2Z7/uiNdqkgbw8shQxdmSEhw+lGup
ZCpVG05AkLmkuhMLT6YZ3XrqoeIuyflMyuz5bV7gN5uIyN7YEbaU7dwiFVS3nYBj
jgVfm0vH2o8CpBye7CcbkySZtAb8Iw5IM8dxZ9KXMZUAdMMbScQA2D0HgdvW/EwB
BpG3ftYfMlb4Iq9Ibx0RNRGwxABMW2mJ44FY1Lyhljs/ZXAKVGi4SfbnOOvgCrjY
52C3MX+rebBX2JidIPRvInhpyzOA7ETo+/aQTmiHdKwKNGa+QS5UO7cr4A66rtFu
mgPxLNLXkbQlal1MTSMERfoNSe+aqkvrkc1D+JhVtsJwC47cg2/T/fz8/3SWGVz+
LexUdobxpYkQGSPLTH+X7ykemMB6UpRYeIGe5AsOYPGvlz5jZJJ+fhTqusapeo2N
HOIts6Ju96eWepOQxZXRukTek6CKvZq9Nz4gamtiquSkcGfVShdu9NbPj/Eu2AY6
TYUQVXnxGQPALLFAqu0/QA1SYHQUwfnyZlOhNfB9AbSm7Bv1u1Zn8TB3fAnXBoUv
33EeB/cethA1g8T5edcyB/694n/2NhMsOqLk2xiDxlD/8IOMUUMlUykrq/0wpQhD
dX7sWh6t4w3p3fqFDNmPJ1PH40mKgY9qqEEVSnlybbPuJWYWhwY2jPNIB3Ceedk7
gXJYsAyE0ikdfJwpqbMkhI44ZtUZraNm/ORpXoeeJKob3cGafCHM64e9I+VtpmF9
vezha0AIlwFkA6GA5+xZKYAfwtZr4x2uuvHUpKH4o0ca47+5bjT2uo0UrBq80uWW
IxCPIrNfwSvXx8WFa075qeHbNFbfunYtR/nlh4h15dDJJk+oWt2Rji/E/RKpa0/D
A4P50I2ef9JHyGSLQATcNU24EpnPm/izaE53CWevzlrruewK6k+QQn8htRsHypef
wxqDWbu/MmKHFhIklBAYYIJXZIz+EWnlfomvAHdjw6KV4ptjZV4i3FeX8XmFbUpb
feP3m5cTaoYUBSk3QToCJscXdgrf+GuaLFVG1v4Fu+Gr9jLnlBXMRmsas4AqHI3O
PDgNl53ZrolNGweix0e3YX6q6BimhX92//ZKg19X32F8IkWnAPB2n8tRRXjWEK2V
KPaJoNbpJUPWp+Exd2y+XHVaMVwB3eqDCup0d8E6A7BmoiRfEnTgwh7E1TKqyT6D
/0FLyRfjLJTAoDrCLSlf6zSHqEozd72GdTOHnc9Z+rfwhr0a7LDQZ00pu4r7S1GB
6r4S88anZBOsqX7y7w2v6SX4dSStNROkXqVhpzMn+Owqgd/iIavhX5EEZrQrqNwY
TyURM0Liv90h0blF60hdi37l/WObAzG3Z/7gBKfNxe/gD3PBgrmY4LlRcF+nQods
En9/pNOkNnkI+yV8RsfNFw5kmkCwjmhsiWwOfj9VJ4CJ+0huF0qy37sv6/RhIyJo
UtvBJxTIhW9k13jomnamQVDP3R9KXXmGGIF9O9ICG6uLotYqMMGiLKi2qBVWVRST
I0hveMVDsnuC7XJp2jsPRnyUgSLdZ7lMNFauEI+Q7J4ZJj4tAjOay0z6s2Zc8oYe
VTj+jkX9ERc1buIa43DZr88LqBkp5LBFUVj6tweHeFjbt6Qo4AR9MISq7Lop6pdy
8V5vrt3adeYo8wa9jmtLiezpbWHcXQGMWdhoFnfrgA6eAGZIXg0kHjN9kj/9eQz1
67KHnwQGKXCzv0DJRBzXnGsvvFHt2Uu2cKA8u8JfBEf6lDDV1DRMbqoAfELarno+
jUZ4pa9wyAmixeQrmbWzhkSiFgkJn1zoP3KrQtI+9Cn0xLCtz0RDGYR7m1NirO0f
7Qrz3J6kZBGfsWsOJyljbbxI470VOD0Xx95qiyjz7qtkCMRxm1SWHKe8MmGxlOOl
1tsEKaRspleUUsj3AXz53JgVdUhQUVgtcv/WwUo9CTLDb/+HMmfZXB4A11HgAQz1
1ilQf5fPBDrZ5d6M5eKdzK61UU6mHE4T6P/GSRcBkFxjCIkwWVHooF7CMCa3Sv4V
KY3gj7J+//kcKh7s+zKhkwBgH6xrwW8aViDvIJF7s1rOcw+EU5ePbSKo4WkTA9u8
m19rqD01e3Kn84DFf+9nTiRmJU0BTmQ+uUuxDEv9XA7sbVfdIW0aiosyyqjD5zUE
DbLEsczzPSPb/8gifcHRUvjSkCB6go2tIs1Jkgv6e2gZJ6h5XQDOw/Ac0DTBgQqL
Rjqd7CY20ecflwYUti1uc+9f4MpdOhXNoQNxRkmRBxbhaxaUsLceNHVwCWzCVfd9
IGyix8RYJzGg16UYz81LafHeRZ9a52nyl/iB6CWhm7UrJUNrmLPyZH/DCD4k/SzO
J7r1vdnKQS+x3ggTbpKD3CfB/KpjxBZ/V5ogow8wMUAYhlqtWyWzFnLk2AfbCvBb
/jWihxq30ftAYK96MVgnwyIhWldIqvsC0jlNB0zIj7CWKnuC6zuPhY1/9ECgl87k
Vwg8TUw8vid0jAFSSSAHl4Iz8PNLnkBrIUOCn0mgsoQPktZPLG1H3VIEdx0+UfgO
AfZTKp0C4DN9vl7/6Hr9HTnYNDIJ5bC+LcOISQevQ/TcOCfg/HNaqepZA4R7L/L/
v7KGdvzVMmwJ1E4H7GBZ7wxWKb1FCe7xx/rDQdeILl2A+rWZtE9d856JtjZICUYV
bU0D8ofCg4lu5wtuFl4D+zTbbEOies3mRLdWVk5WwmmsGjznegASiVsA4I1RrUIY
kK4/1BGsdXf3Qhw/3gV7J29Ktvnfc0QeHGYw/Q9vsOUHrrcQ0koZJUnRDWgor2SF
+uEah3ERuOvUk+NJGcMlDnr7eGlPHNHL5e6QaRlF2/ju3T6uChQckUa+PVs9KJ+I
1agFqYEf46tqsxpogIX4i6jaZ2bAAmV5QPIUa4eLg/YT+uN49qFuQFF68DH/S9uW
boek6FU4uS3s7yH2gL6OPHwnS+6EhalT3HFsohYRGjBJi+NQZnp382AYkyowHYo6
Faj4QwEteFLy7T9ULFeIFMAZYciiuwgqmqHKHrfN3n8M7vNXHIHoELnaB36gXq2L
N4ex5t4I8aTVHE1C56zhuhq/Ra4lnbzqaSccYFeVlkna3NmEYh7qVawRqc0CDpRP
w1d/ARmdwwW8qBUOaHlyGgl2lSltvr39OwwJqsW1UZtzVgS+0QWheVpY8jayd+dX
yVFbXSJrAHqVSlX7SPfqfVdTuDlxO5UWAEzQLhw1YAD1MxXfBTjdOS/hpqeh4wCs
Xzk65PY8M0Ose0hz/wWrg267zjxWIjmmLxLomCk8Ana95MVDfKfDbk+VewMMya5B
lV6Tm7yC97Rfclfd6Dq+bfkR9r0guCWHkbj8nfHxtlR9ynAOelnbPFG32rSP5fVk
5HL/Vq0fzl5u/hMrfoBtp0GQfYABAXuuLYiQHKurn5mmYhk47iEnlTg49ZCn4lMC
c85eJCcciYlw9VXa9OBCrlrN0/jMDw7uo9x9TKbOlvDA5sthMY8JigJ7J95swhMR
9aUQMydXjDZMMlkjz/wHxMXESAo/aPWtYyJNMUTRjlg=
`protect end_protected