`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
hVdJHWSfELCmA4ds+csnOQAALbB3ps7EiTSHEDd//nts1r+JQrRE4d3bDPRJpiX2
Sl8d+xAK9BIi4i+3ruAzYvB6kuD7r+gs02Jsvd/1kn7JYK4xBxCjtdDFjVHOTEl1
sSh1oNiYUwLuwR1yKfP+xBhqxD2Dv6pCKhH1NdGilpJQ6cvivGkSunAu0tzP76T0
4x1pB179E7uIeRplfHWX03KzEBF+eVtfgXVp2W1BGjfAe43y1pCvNYZOh1+TY62g
EgAFgbo7pAujZxZy/YSiZjUr2mGp7o83qMXyusx8+rQ41D3X6rxfuP0RiId2pOpC
6oq5Dfkx04a1dk4s8w8cVg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="Sm9DkM+kBxuxXCFA+l3fFkxuSWV4xqRc4Nn7Ji3ukao="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
m2emGBqRy4AuduN4dffN8194qYvc9UXRqiQc56IrQYMiIVQPyh59I8SYabcDdspI
7AFHnvKD5YaF6tQfxWm+mlcmMEk2Y//aUjxeiGGs+RkKgbHitJF/K7nqg1dmKvDg
a/GaBCq4Bqh0EehlN4ntP5HxM4qcvSfh5m/Coe3drc4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uG91daMWA1mGkhgP3oZKMYye3UAomMWgG80HuuXg2E0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1456 )
`protect data_block
c9NqBF2D1wSep1rW7utzHsk2j40aow1MnrccxUTvKej2Q1cyeDDbgAml4eTSXI8z
QYgCADtWi7S8BeChdv4B2VxKcS7CMq/DaQrOy1MKTfQzfAlK0iubmlTkljLy0Rwd
cTrJKn61EKbSa1l2NxJKw6z/Ec4s9iHLNPgu+vjrcFRKqe/NVBFYFOTgsLBpgnR/
zrE/MZIaYUnMWG7fDZgLJO+PzunP1BIYQ2iT8VWwfMatMDcfia70vX++xEe/V5TU
V/gNEan+FY/5P/BY344THdtkwHijQxWe/Gz+fwW1J6ms0lVBypCJDgAabUAXYQeG
g1J8m/57LPtfegm+6vP//P05Rg1pAsBIAwieYz9rLuuygjKejY0sxIXY5DTMNCAx
7drcXZJhuBfRpXLVdKbCCxpTha9xs2dugiC3nuCyl6E4exIGogA0SIyFjf7u2p6o
9Ks+RLtD87R+0D41tkfJ113K7Lw9x+AdW2aXJV7NRDjijB+lURJqwSOIzTTPopGm
utfK5lcWapERc2ROFt8xq47jrdlVVTzzHiyiQ4cIKl6zNPi2h1Zoo+ypVg2VeCYM
TscQsKJafE7hbtOrR3Rz08TWpWI6VZwKwWmWzeg3jXT5byzLYu5ayl9wwC81kN3b
rQb6OUMjMBP88dZ4DMX1A7T6KBe0o3t3byzqiFNjjuFykq3gsYxIRp2YZknFznzN
XwMfRqpXLiIQS57Md5dKwFCGN52ciH1vS3P5dUhQkNN+aoN/yPCgt/Mv5aHvVstd
uwjbWdoAWsClek+UrD6ZcnZ4jQyUUjVrSUOJrAhNk3rMKWahFoGwnqgQB2Sx+wF4
VJ7mVrD/7nDWM21QR4jUAHKmmt9h2dV9r6G2muztIioB/jwj7Y5Vq5AUYfP4LkpB
xb/45fpVIqFv8ZlgHyEJuKNljq7vZxHk3T726G6EMxbs8W6GyPNZxa31nVbNACC0
0vF01LpXGoPJ1xrczExURVrUBc6jVYN8SsZRDSnhU3QTXZsHPUfYKVjLaHt11u2x
+tAc2SbHctEh6e8WAQYK6PMOeEmD4OhC5T1HeQepD4AJ0ZH4G7+DhElQM7EysTgW
VydT2r2TtZMdxFn+A4S5rpcXMBQ+jrMv72FiroPcduKm7ZUpnI/M8MMr3zI/7ayI
MlhVE/szteKA9KwVZWawegVnqzC4bZ7Yo+txFsluqxOMRMoRfZS0v/9dQMDd9i5h
AQufvWuHujbcVN0XaLC0FPpWagmhC2tBgr84enA1R83VSFEfBXhoIdIux207aDB1
GEHJacqsooQrf/kU38J5QyQ9L7H50PMSpiz7v+6mEd9U15/VRX+Lb6uBhcTX4MET
gwopqSfLKD4bg4WiOetk8cl9yW01Ugi1cgKc3j3BOTLaEEWnnW4JLDaCayW6sRAZ
YuJDSUa4LGOWwQ7v+3p2FPQfY/fTn69/EqQxLimbbeOygZC0Tb3n4rWypA/CcPhv
jf9VvxYkHwQcfvbcC/jkuC7bfoAx5Sj6Kns09IXODqJu9qpYcV3JFYeeWH+lZgMh
Ar9F2wnL7KeztxfFf6V2WfmRb9pbeWTemEh82Bwv0basiA9DqYZ7Rb75O1urBZLy
rCgWKXXBmm+ND4PNWJyvzAQKJQBjtjP2Grsz3Zon5FiT/ZgMxDvlkowZgJR40JyU
A6pc7/jUSoftz/iqeLbhsvoe8uKjU+uO5pX46pmjRpey2qODIwt+1GdCvBKHp9j+
iRRA33oPRPOEhAZSrQ17XTi19V+b6dsGKh/1DT0DIpEya/UNaAzo+ScDssGt88Kn
JbvnrMFhwxTsgUwlUaZ7Vmwkbz6Fc6Lh6Yvb1aOZpXDwGVWAKwY5L/Y2TNg1gIzx
wpZokAbUzRUV/+juLbw2V5s6YBsYtpa7m/ZTLw49JjLyGav7O1uigyyE3Y4c/rMX
wbaT00nwhhmXFZ/oP56MhA==
`protect end_protected