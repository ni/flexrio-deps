`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11328 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1wB2ShNYedzmkmBWjqK4Mg3
8iDfXbv5M0vDNkp8sRs0MKOWyhBwqeRD/Axt+WhJVoaNd7LJr5CVJUW5C1bR9Sfr
Mya3hZnbv99vXgj4RblPNpXDbYEJ+AhLawMA/9UT3meTp4jaIAHAZatMSStIMnLq
cpGc000PEHrz1gIMIHW6y/C66gups4jJrra/aEDQ9nb2+aQfU7xhEcX4/KQd9FDq
VTy4ndfRL6BxqRac6Tc4uzhDiVuADe4TRFlUJtKlVSemCVEkNN0P71yNtkfztEnx
CXrC1NS3BnigT46pQaFKSrxqaMfy7k4wNYNlqyCGRXS3Yvc9sqem0UgqNwPtwcWI
jN2XAaox/ejJgxaPYpAdPvpAnqke+2AQIIFkPi8dwGnkqrZEaOfQtp+j8KMPs7vC
X+sKpEPAwtjCD8rsSD2aEKJgcmFYAvA+hlPZBhUZjJLlLABbxmkWJz6zyYAP4KgK
7+DNwWKl5AUvC0mfrdf4tDWzAb60lWaJtoW0UUongaH1s/E57zvb8ffdPlAxu+rb
RCYQD3H2jnWX70/cL+YN+zydD7m6Gll3ZMpuS8a6ay7Qh3b8z8uAHF3FPlqZ6uLj
buJAI2u+0s4+nf//iW+bRgo+Jf9f3MCS6FBZcpevZSvhs8lHSIvA+xYlk02/JIV+
i7opL7BRQDRalhWrr1MjTQOcuYaSMNPcTZscg1foOuXo2VlkTqxMxYSKlQlmfxd0
RZj6hh41pcGsVHo9kXUxlRHu/vMPDEmzhUHYs9t+ZEYsktDoK8FwihYtbHOKGobh
2EB0gD3+k+am2qGsMq2x5mJP7q1Fc7kEaAoicxd26x3Qwu26upd+79Mx2Nf0UNdw
PYAKbLwPvTvL/YfQLoWisXtPLashHeDPsen60wJ9hkBLCejRYiR/8heip3n+rw+4
eTksA6FLf18fez3M0h8ljt28Y3B7uXfeSoDfUoR7qUM+l2YsBwZERMyuzxeO8exi
pVgSPBKrIpZXhl2JTGZ0n6i0UtvFnCfKZbfDSudrtrFA/NKP78QWV64ECgvDnFvC
X/HKmib43VE3rmfcGLfEtlfTC+5kEo1AwadezYuqujvIxIlsM0SsM4dNNkqxGnn+
o8MVmTuqLiwbLPpKHVLeLnwhCDtPl5eDYHAeVNzboFahh8sY9wYHkrpIVRPOyxB/
zQ+Ikw9xVaOoMyY97Wbhye9F2nWhushMR5/ZoRhhmbWXxkOMwlWG7G+3Pg1q+r0j
gmkjYSVN3DfMiaXbPRmsG62Xz31BMOzlilgiO5XdRmSqZdnubKhXp3Wr0Q1+s6sm
QdHFB2u/6Bx5wpAljsxIs6+dmVdoaYGQuTf0raNfiATD1eYwyht+/NTcFJ98Vdeh
hY9DlYS75CIvj1aWKmPwGOD/TPM6fdHGoQ09Vh2SXMq8kyVRzO3qckucRzLMZcye
VdoSRQ+nVuCCcIh3fvmMRCW6bEFZSpaxF9DvW52oq1GrPZZ+SAcihgOvo5EoRY3p
YGj/OyPLGTiup2D9IUQEQFhHhHyHtJFjU43E4OHObmeZPDTHhw3ECLeAFXnSwBKk
Txoz+EOKZ857IcbyOxtw2tUf9jVevrRNMB5/RHhqTSZnZaGN34Tb8JUjGJLnDJDL
q05OJlJQnuSYm/EQLjfcpV6nCBjlm6O3KsvU4xkT/nAbya6wsiGPrdR+NwxDs8S+
yH5rJvmG6gbHUDN9QRzpmqRt2D6kc+gkYi7mEzp3z4IVxXCHC9wIxQevEI3PKQ+V
TwOQ/9O6nl8Jpo4a6cWVvHIFv9UxDWAB99DPXm7d5bEswyRE4pdousT3tYuqo3CV
o2QYXhQ8ABEXrQnJpEaxDl0SB49sERga5Xeyxh3lBnXCnTtCAjQ520m/gInRoq9d
fKu5YM0V73DUvUC+FUVgbXxGgTXicsOzgbjSrVz9roGT2IhWUpWy13NSywqBv8PT
PaVbW8JDZqyVQydZZjRAReOwUeryoRucTAUCTuMMl05tMH3W/Bjdxec48P+rDKMy
yzYvHqtrzChCGFWcFtQ/ZNi1WGLdWL1NsvoMPjJ/gHNuGWGWSDlgWYnlVSMF/9ol
w2q/ZJn0SngHvx+gEMxd3vQ7dxPkX3b9XjfXc+R43L4TU0JlI41yodBBvY1oIiyi
vSf0MANVEMPm7zY0f9iDnPwtOrS+q0E0rQDCw8BneWmKF318wRdcfwqilrHpBkDC
OhqT3DyxAHRUwRL+gqi/Was2z4JlX/Ar15/ejYU9d9ZIYT3VhO7MWrbv9kWwGCfW
MrLkhnx3+Wb7FWlIETI1HMAYWB6VTA5y3c7gnOmXFkMsIA0EAH2dEJeGEMb+DKfo
H8ot+4fEF9f2UZDWuq+sEZ1PE9jbggIcFxpea8AdwZaRajxAF5Qwo1va/5Y7cnOY
z1dVT9KopmbsSRLf1+0/8XSMxtLeXo/KaTzxLbYZu6daTmPlN23gIHY1FQKB6/mJ
Yoz6DzVQzybZI8EcPvImzabd5ISVeNbe7dgs6t68fv6iW16jOyUF7Avn8759Mzd6
EjZFWxIDMTNXUMtRNNgF4Y4ml6v+piqly4o7+/tj/7XqxlgoDjmNZKX2Dy55NteK
2AgU14TY3yx5UCI5LXuREXtss87+WBU1vfkmE1f/uuRM4MpXQbZ/5BwdtuqKOWca
/ne+1Z5BDn+tJV26Ax1dYrvcwR1NBHf9ms9TIG1bok7a+xlN/27B/5k32rIn5VMH
Kz+mUeCv0dA31dvscvbQ132mwplUNG5fYFolYxIcOagvCrH37x8irVS3RgJSJrBD
LGQEmbBURxuvWV6Ki+RHHsX73J53bXFQ79LQDxv6t9IiQRlPLFVyoE3CNvJXovzL
y+v4b172nBDMmxIfL0YzUsVS88jf97lWYucQ2yY6RK44hjn1pDJEvv1pRwf4ykii
IrQQn6TMBZJvADr8LxHMH/1M4JzelJyZc8uTDAf3gzWBM7xEMXzRIe5qnnmmYtNA
GajQmLjvoC+klse0fTe0HsHzRoZBFVaqTaG78hIybWZZfpkZZmJELwdBcJdBsB08
em/VJ/SKTbXK0Ep+CTM46oQOb9KPv35oIRVRI2FkOIwbBH5zC3hdC0y/eHTBV57D
pEVGun86zL3dsT+WBmbp8+cFsb7np7BZ2kOY3jsMpq2s+XwOYzn+LdOhzCR5TgDx
xcVgtv9ox90OIYHg5ocLanDiqyqnhqI4RsW9lEDFS38Is70d2aWZZLRShM7eYl5Q
oKnlf3g8+LmI3+pWNpHBsUds6s3cj6M0tzcQtmLRH/w3llgT38ugMZ6qs5N9t0rB
gQ5G0y0Z0PRfdsbvcrZeVRbrJwgV5JewjtgotCG9gsSvdtt4EF1gdjwdHqREYm99
IJKL/qSD1Xcvzho9OGGe7pSWXeZUJolpARl85VU/j4vd5n6+ap9j1fowHQqKDXZ/
gFC3TU+6yxdDDakEraIMHcGA/ktaXD/iD8U39MNi/+ZRGJiSwrFO9e6trL5pOi+i
bhn2xHj5/NK/HhRCMQDLxM+RDlpqjcrar/bS9trBHA6NM84kPHhueidfz9QXfqsv
S1bEWT2My8OHdNOb0vDNvDYfxEY35EbFcbENRQjiA5GWhM775OWtJ+rEOA9nFMZj
5iUtTLPaZAhYmomtYqLlhAWeGwrvxrrKPIKzciBqCn9y4JizVOqB3LC+zClhkRku
dqmJSr/BFC9pt7AjPK/IPrig2sozSTHcrFs3cDl0G7miHJq1NZ0NxY8q98wrakCs
NXQVgHmNc3J0NLPMSBkw7+cz8E3OR44rBHjIQrwpGOSUzfcRQQu1z1HJFkM6cYl9
2pB+IS8abQ8mcqvWyHFvEzGcYMf/lArrCVPZPze0iL9hEQZc9oxx8O549oE0nR1J
eecTCEqxi1J8fi+MBJm/eaY2ySvQWNa2qMmH4qXAfde7HyQeRi8g/KPh6TpO8yCU
JSRJeR8qT7e+v2SwuucRGAewbT74KSbelS+bQae9ubblWuvG9UwybXz5MrmsHkOi
VyYJAt7pR/QqTmqMa3V0MZlB9UylLoiESE16NXu6pS0ADLk1RMTKqQwXK7ftbenk
lvihU32ezc4iXWIzPvjUQyqG2is9HE1COiKsCx9iaQQQRg0yxcsffO3rsqt0VLxz
XNx4lLbcQerFtV9L6g2QYuR2IEQPtbrhvl3O2uTsImvbqlGMvlSejRCzka1ahQSB
qlYx+T/f/pXp9Wwjo1prPPgrFC8PZbP8p9MmlXTu4r9xYfaZKmNOx+DVtld+WrCH
wPHRuV1LcEr6rTJqlgj4k3S0ERvF/mr1OZX8G+0IXUl6hEtLdOLke6R0Za6l3ny2
umL8IrOA6TJpbXVvRW+EPv4H8juU1YsAHMYAJDTvcBUONZmo3assEnypOn9QHOuU
vMEg3e53e5kezGFr44l5Cim4bFEgV5c1IFkU4pHxIXD4T+piP4nrLyiQjrebEG7V
pyDl3Le0sa2xbb30j15vzeAvK6QvWfzFJnoWbeMPcOOyQypWV7aKpXjSEWOXnLo0
ogQXqJa4gjTdLPS0rUkKnuS9UTuMicsw+JQRwBpwia/8YsXumyhzYrx/CFPdbAYU
ZhY7o42KTfauvgBU3++tfLcHthZRBq/zbGfPPv3HQ3m6gWs9oZlHvb4YzE5h1FdB
dDJuzBkKEwad+YrDLF7u54aHcB2aOKpCbMpThULzi3ZEHlq45+hNRwTUqIUwdAtX
+Kmawl36QfJEOdVCc5VG5AR2WG0+39z6E1CB4HwvDMW793Vfp8DHO47KYQM4bxx6
u+T2oi1ar3kpOO39c/NM1c9mKS/wzvh24dopeHJqK6mKVApHeeEipyQ7H8ITICLf
h7UIbryr4CjYR3UX9iyGykC7PnEfiXMP2PuDMxOJpvJBr+dbNHKt5x/xcWlX0/Og
tLmRIh0em0UGhHnD1fOqfAgRnBGiBZq4Va3pNG3F0J67DZjz+vpJOF1wnYcKrKgL
PF6D/OsGvJ8aL41vlnsL15tkCzpbLqhCYMdV3S630pOnUYE6Td2G3y+1+oYM1+Es
DK01eB/CIcqP5huOc4cO+zhLUMKG4Yxar4X2xd6WfUxK9ohOhilG2gHbuAXWYEHd
3b6ThIxMMI8VT7Pcw6i4u9Oct36Qv0X8qtJ14uWMSEf7M2ppG2X78Eh10419krJC
gEJFrp0AC+aT0mjE8emsse7ZUae0Ssi+HMyL2OvIHg1EBmuwIHBMZf63l4pUL8FW
yQR1qyv5U//y5bL7oEcYEU16tY7smMth2nZcQO7jHwx+gCknJ/oZ5nDi0SNEiEr0
O33EH383YCMaHrmkaAxrJSstnI/a/VILSxQy5cnC2FF3pnXkYGuFfgmdvCBtyJTJ
hi+H7TW8vazmXC6OQ++QR/g30cuMYRi5w5pyxfs+nvzgbgSYfQuKnV24jYwFOwPA
r+vWFEcjQwgTy7BR+aShrrJXdfZ7OokfICptJeq46FYX7vLtNIq8gOV0xGM9tiKC
1MCDKgxkmU1XK/hvPO/Q5pW+A53Bm3aQdpjON24fq7i+xM3cFFJds8tm47yPNwDR
wZ7KAxpZuZ2yTAOQbwdx0qQ3tTtd5G7+aZAkTjhXTGvgb46WpDvWCV5a/5cuw1/7
gBe539j5qjK+9mtnBdnNZX51Sr5aJU5E8eMK4e6aeDX1XLr5GdgC+SfcFNiJsKoW
GUCV8Pgi53iEVjeN8a10xmRJAZDkc3tRebluJ4H729o/TUA7p69J2RLYsndfoC8Y
kdrUfEcOIs3ijltpFa+zce0pW7RMR1XafDmjmIIzfQiaflrpaVEQg2QAgR0W4mSQ
4N7zSvRPFVbymLMjxoT+6q3AOLzbS3OYB0hSyX4jbsmHb74NdvdA92Y/r3RmGgnf
GlIC81dVeReoO8cBDU56MlaJH2Zz/A0NBPa1vL7YkpgahzGUtmIEZf/mmZIz7zBU
VlDacVVQnnBozqX/02yyJwXE48dC0yCc6EENWikb54Jln13P34BOuYQb74CRUftv
Wl+vi6o2Lt1Gp9tXXrm+20tr1AQN/SnpIzPYzc9MDRiRsvl5YB6+NglSDnudXGF6
ETw6vy6C0UvGbDgDX2x57HcU8KfqgCcSfktEdb7OIxXg4gpggsCStaZj+YjDFG5z
oKRRu7+wXDhGFvG2cbWDTv/0RNCrqrB4cEfN5lIEI9vf8MMZWQQv4+x+lt+v6t9W
fIs1bH5MwLL+zufLVW3y8a5rmjnd5/ivazFi7tjTSYG70drXpW5nuQ4MfcysL3Ro
vdFv8Y88ENZgnzmXhJdGre4xw7oC6yIeg5QzfYRjsoQ/kwb8JjRUq7TluDNpnilT
CPJH2yUjfMeKvtHV8VNn8c6QU4vr5rFKYuJ0bi0pt8lcjo6H8u6Vq9agur7wtEeX
OOKz+aFY/c7ln6w5tdxqcrMZK84ylYRob2UEMug3XmTg8ln1JX9/ISX5a6PkbrAN
Uk4Oyebc4j9Q0iMcroeWgz099XUmttgT8eLGkvgMcuCAh+QVu4EHKX2/DSTQb78q
s8Ct8AA8neJtaREhpmUsOLCq0PuVajDd5Ah2MKVqBBjAbtYQTxWjqdzxql3x4pOu
zBVN718S8tpElt9nLuiHsZ6n2HSS1m3A4W7ILOFAfN+Zqsab97ACePvU4bnc2EqO
vpUWdx0dZHXCnbLzx5wTlDCkpa7RxAuQz8VGcSZ7VOCcEaqamfHr/YY28n41ryNv
vN9Pa9UcGIpE0y4WDv0hsz0/oPLhD3ewBWInIR9ru9w0nL/3w7cWhuLGhlI08kuQ
pNUBGAwnpo0W5ALjH+UCswDHYjRG4IPCx6SHoc4wOI03/T9QQa4DLcoYizVTokq/
OeMnUtsgZDDLHUT8fmM1fpxfZcPmz8fTKkSgBlp+WgkgYgzpoeKfk7Il6aoCyp4H
XHV6lUc+ZG2b6SFlnpqCjpOqKvQLkxbqQBbZHZIKR7sLICmAEXSxifGjIMFvM9LE
/mEHkP4vBLR9bV/f+fEPQJjZtwo4Og22s5UPZ4CtJQvJE4EBjxv/9Y/jF+DyQLuQ
hmXZWOVfGS2wcqoCWMP9sNUeXFdLSLCCKnm5APQ2LeVB5IAzn6Ba2qHLLGedkqSQ
5ACH6W1rmdxigdu7FGrm+V9aEvv1bgtg9jRFxZACg7DJtssb3Ubp5GxzbyL1d/l8
+byBeTQzxrXaJKqkrFLUEsfcxx7ZsnbDCARM28UL5UfWkhhFKXLKXngDApiCUCts
rdnGqRZTrr6wYgmpcBsh9K0W+pYN9YylW8ZmnOGnmDe/WTdSx2xAuiHRT3iNtl1p
EuKkE7bf5PMEdTDIiGHDFVeeyQQB5BIUU9lXm519Zawpt2tkDNIJQYhR9Jm5rrEb
YdQiDRbaQopWidTQOt/D0dth5zthHef8cS8bfxKjzB5y9T1VMZI1l8Wk/ExSJeDF
F/MTJVbBurnQL6s6hXJex6niJBOnTgTzuKU/y4nH1y7T1FXYTVI2z2nPmV0uYmaV
r47MQuRDWVg6MuYSJT/8YWReggSRP1nBs2ytKb3UNsP/3339ghJF6cMjRxYxcNgW
2HGGdUAu5p0fxCk52gfIwUYiyFv+IKt+XQsdtNlj/7O5TNFxD1fqdlrvIyHWu+mo
0IfEftYQU4RtsiGw1d3i3tkAbkLVCq+QMb3siIYymiq34A9MkGiKU6LFKuo3vkOS
3iPij2+gdG6aIuHaXdx/+VTyfX11mtUzV7S65P0/qQH3c9Afs2/m2mX4TSWb5SIZ
fEI9CBPzho4Cm5LJoI9nxsFmmwrfBfhsx7vJIjd0qLI/aPGrb/MAcDnZODNoHysS
UCS1LuQj7Y0fQDUtishZ20UyMhD8El9CiGCstXz9orfMUd8eyXBr8fMWXRhbqlEz
KmOWwIuKFsVuzDflmNVVUhxnCDU+OGaxaY5YkujuZ/LnKnalIRNjXiYNP3qCbniC
9OLZBD8YkbSbumc8yP8501RBiV2U2Kx5HRetfPdfjk7DVT4/FvqUhtFXnAdiZ+iC
dSKvIp6FMUJE0DN0G52IsPLvriZmrni2VfwHHnBoMCpAc4L7Q12z+Yqsn6tdz3BH
sopwopZn20/IrntoJBwck/RGGKA7mfIX7tH/zAV+08UYhghYJbMsjdW+VXg7YUOa
vGQkPo+iKblJx0B81wggyC55GPyzp/UPI1vhS8ZwbGCoNU7Na8VodcITq0p+hqod
VFRwWlcHthOBdEy38sL79f/kKxV2zk5JRfwcJcKOAqvltuqOiyrW53Cgm+OsgUuO
wsOpsH40uaF1miB2z1EZEWXCU9Nr9zOW83CTlOIOamIgGm0J1+3q6B5h5ZjhAo24
5tnCUn5jRMe7sQI8Mnw6BBv2XrpEUNlqC0BoASGzUYW81X6XTnU7M+9M6b/DuRn7
uiPivk0DsKmEpkwZk6aMT2jno6P12uCcjA+y2k4jLqz1ST5cmzpg+XxC/sPco/Yv
M2z/C6f87QFThSNSY/zM/v5L0OTkyau5ZFTN7a0I/OxQqbtehmW9+pn1ISTgbVre
qJSPOkZd+GvDQaIkr9xhHT42uXilF9ya3OoaR5JVY3mz8XycWggXiG9eijmnFNM9
lt7hx69TcGSK6y54ofvFMZ7fRHdDOmgbpIGO2c0vI+6TCirh03hac3aFtRNqYYju
aQZWFBKp3H2cEN7POvZrL4058e0Tpxu0qdR2fWJCTFvFDa9W7SHQFswI3J068uvv
Ni2rSgJTW4zwc0oTdjd10qYTB1mzn9is4jc3fsBfTWYfDG9/TEPCtF4Z2TnEUHIw
dKZH8L3M6CPUNXmRqRKHp4B8kwInsyGbL6CRSJ4NLNywlUFLIfNn2V+jvbGbeLaC
QLV7rEnljtW83RNh7VWEpAjKxJs12mdRiG66sr8qVRB8ePkAFRdRFWhRMCyUl0v7
hXmfpHSupeqSEcTrDUS/z7BelHSXQxj0EnPqwV4snNguiz3e3JIEhHcWwIs6VeBw
qnrRv0R7gVA7oT6ujFAboi70ZmtjohEMsiu1aRzG1sDPlVV1OFNKur7puiZDHz/x
2YXgq8jV7B+0f0WSqlOFWLC+ocUylguqJrIpIkD/z9U3XGto5c4WNLevhZXPDqYT
xLAoQf6KVKZ8teKGyKEyOIJu3IJ241psOj6gPYviUtFWJDMNioVEgG+T1qL4leCk
Xo/d4GEVRrVsHTB/9dSmpkGg+FZNR85L1onSP3kKeaxPLau+9piz6XVKo2gDa1Gq
VVu3XUx6rep7ora4Il5kzLdq0PWbzOxCT/3QyNCbglIIkPXcBJBTXYhv7PZ7zlPy
NdPxqcHRULuK08VoNabAx4PBJ2RA+1xLQh/Hz5znKc7KlNIPxXRVTzArsBkY1/Bz
8B3MG5JuQscGukufBihcq212IvsvQbfrYKhQM0dYPnRHq64hbScsKeDIHtM83cq/
X66zNUrpBB/P8gdeo4dBxCYJY0sjy5/NHzRNOkIsbygXjCnNUa9b78MC0cHwzf6a
qZr2QPVgpuS9A0eLeG4DhjWIu16R1TFDOwEvArk9uacpxoIbmfE61+1q4pDlwn5I
Z7Da37ISwFgf6rqBmPZ6b0L4ArmJKZjPsXCKLNfUEmzqOVws1GPM3ee4E6m8Acvt
gHhHLVfFyGtnsasf4L0CmjRNG5CE4cLbirTpnC+jzqqHDWo9JnSgLQywP2fBvjwD
18s7YtNstX2jxAZKqCRJ2CSjlBpLj3GoapudD7g1yMFY+TTd9boMmg06l6ba64al
iHfZvNwcgS9yGpnMp/tN3mkV2E9El5wMZsu3B7F9WaeJVwxZZE1SIbl0gHCgRrCn
KuBnOhUYHPxWD+adXcss6Nr4ocsuBDS3PEJbw/7wpsWzjq1qb5FVOCrTiMGGQQZD
GkTRvdfjKOvSq8UysSiAsGnbLEFm1nI5C8jBtp0TC+EoSvnOhLbaQ3hmiMox0LKn
RUb0CISuarwTQLqVVUeW0XlnEmUWyxKX483gyrSytUnqro8rrnY763AwtPkNhZgN
5KX+UgzlwFQNNUo6R9tgvLBbPLNRBBTrOG5WSG9t/xqBnSGIo8a8RpaUmkdU1qLV
cRBa4rGWC8fuNFPftG4TdpUJXePDkdQq7lH68Uz5Fc0miEcr5JvT7kwGGD0AAXXb
w/yu0sF2DuwN0aHTIxjgbDHW4x9xYHlRYlm+dylXZ+FPsxPy0uJp8ryuaNu67L0z
onjxQwapLpqmfUDRJ9tkmeFyO6+Qi3Dk3nI08nnZAbABlHmxD7KO0T67D8OE0OLU
uD9Rki23d2YJ+3JUXnbb3Uw35n6cQ5rNUvk5nw5LekEn2+eOpA8GprP4POK+LAhm
ZZWqJEUR/6cqlcj9UTfw+ABO55+wPutyxW1BUYAUZags8a6VameKIkSQWzvwYHTi
ZiG9IYCH4UGufWjB0irNOuyXcWOKV3NFhtz/WrxdGuULsltDTNHh/FBLfsQgod9v
6hTmPka4yUE1Xa2JOtle4uR3wkDVUbiHcFqFMgulm3zmHuwumryP+5WHs8UAKyNx
OGPYPeeVZo1eOn8HbW0SRBKUWjKZaglz753MOhJREtyR1zzN3+oLegDXmY7FI1Vi
1zpQRZIw2HyytkQ5RExlJGWtvchZuQRx45b8qLkZ1vSMfT8Q1dnvABwRoBKR5hsT
nIW228NIP95M+QBcZbEZ1kBI4y+d3K4ZZYb05OTsIUzclf7ICbIrnvBm76KX083c
Qig3LJl7GALWdUUAmS1RnMsbx8XkVa9X3j9EqgfFqISD57TfvXVFqLvQIssOVa0k
lJ7jJEBRh4mWUsFE5X8WsYV4lVtS0o65biu1053hJFhXubYKhg2chKWTNUl91MfT
OlSmF/P3emGcc4xnGTF2qCaIns8SYOoX/oHU3bBcUuy6kOF92En8ZhlVq/GCcBei
aOcSUhXIMGyEdFFlWXJZaxyFDFFMMnHOmjjjA0ZRA3+D0Ys4HYsvg5EbWt+9BrKr
XZmOVOkJu158MHxygJ/Prb5gKMCC2y7ekYmbBobvSiKahgEIBxmbcPKYETConfO2
sOZ0V+cIoqjQjt/XWblO1FQpFgXoyyMxObYZjaSyySilfc3NtmHZntRnoIlM89SL
Guct0Hdmfy9Rl+aJ1gtT8romILPGsPjbF4YNDzaLVMJIi+3FJfejl29rqV+Ne7o3
v1/vcy4Q30gWUuNDVDWahHVKRY4meolNp/KUh8yGjF2Vg9uAk10qSj/L6WUmiC+T
JnZUN+cfdmTZcX3zgmMSpPyV1xZlyhx1aAPAukOFKwjEeeWfesSOr5OSJ+C5rpw7
RJtYGtho3IzZLuT7v3z9aUXXgd8D2rwTQe6Msj45VNjNbX1R4veMGJkCVUjCk9tY
jGSgKF1/K9C52ZdMZTWpuojPxrMjCFM4+xE5NfF13I04iB6fDZQ504A/b7R0onAi
I9U8DOKRDclHq0D5Of7YcuaIqV716H3uEezntsiyKrbLdM+/aXHsdGKJDRED7NvN
VycqutGr+PB29s6g2mRzaZ90RRUd2F+5Yx6z+BwTyOTlthaPUNYVkZGhYI5kdXPu
sfcPzgiIOIiret9DqmPzWQrfOt9UiLxZh2j/5vvhhtEctt3N6cQxH/fT8mMsjJub
5kDZUV+axerp+4hMR+LXIrL4ZG+Ek8r+5nH9TEjKTjKHYnzb5dL7WDMtOdh0VKnh
R2NWQwcomkkcNBUoP4n4Fkdq2opu+snWtHeDMSjF/Uvm6oEHcgodm08SqMZbemWw
zEX4PVPVFrT4tpegv0m0GZUePWq8QUsbT6o60vNFXsMjxaR3I1mvNYomcgQqnFIu
UdWIFvDbf7/OmmpeY6JG/tr8VsGzUisBMMjmJh7/9wB5f3Ok6I6FlzmJ01g5gAbf
mXIobgPNHKp92lohxjlIaR2nnCBSe4t2n7loaeQLwTvmG9R/z+p68DK9I3EFL82r
IOWQ7mNlBe3yLZ3b//e5S2td0iwLHy2nCOhsaSnD1HNT3Q7Ltv3+/iCAsWvsORx0
mb6gyLvlqleVzyx5tmw/J1Uk99Q05UPdYeqdQJxIaJHFBl3zBW8M/S1C1a6KucLI
wr4lagnpxwPOAypw2dPG5Cb5Ufg1CnRa1iLHZornXX2FxkscvYxFMGHjIijkgMl/
4sT6plUFYWNrITySR8JK43E7Ajz0qNAF+1vd6TXEsrRI8af0px7jqC9ivOMuK1r8
tbKJWvvUZg/9LIs292a097J8F4P9j1BdPtNU42VTpMhUoQxFAf5gLi/bbsU+XUI4
LgvSA1Ckh4wi3gBbyy79FnOBcEPAq0MVY9a0JTnCx8PzaJNm1wwHkYiEqzmMyk5G
L3ARml4Yh8HuVokYFyKnY3ceMdmTVomZwe5st8+w5ac1Aprips8xQgBzx5Yp7WmD
NdQG0Ljv4Syf5H6Mj96/SHuBgNFU0PIPk2r6dGAsBaHakL0SWs/4EO30P5DUTya2
uilvveqrQQOx+cNUlSCC51/LQWO+EYzpBjNKk4YJLYPFhlom9gfXod8csN6/KIA3
/8fzsUvmmiJy96M4N+vQEnW2NZUS8XT8GvFVe2V4BENw8Ze5+p3wF7P8yAJYVBwX
6n6zWHw5W42RYOxBMtuWl2vGoChuB8gVvXUgaohMbLNa4k2xDhY7GogqBAHalQh3
qWjrijv9TWw6QDbONvBZo6y8RQZRCE9mXHem4dI3TTyxKCk7bIer9nBy3xH4IDZx
Rzq6vXWZF9lo77rdchnv4y4GKPDy6cZczG36RTtmjSv+M4vZFnVC4TfPsCFutFlT
64kj17ZzyrV9cj/w9T8OoATRdR09xAwPkL6UWiPZzI/LNTwu5znwvMJAHquKtDex
dZN28pC0E7OxH0bD837R5dzXPUY4MudpW5eBzK7o/vjhPoBQptm3N7VIY/YK5rD2
hMc9l+TrWbs/XQQ7vn3jsWvDbQ6aH4bB9IjnSlEhqeDJelUwWSVexkFXRp8+6KwA
suT9MvvaB05dlaE+Eoy16mLozkeRYfVOz6IpMuVWlmBhopw3pEnL9Ufx1+Dy9MaN
qT0PxL4QCS4UyQpx/BRjFtydFbBrmR7zcnFHuGuzXzZ9XcI9T4owaJqIF7gXkqtn
W/WPprne0B6q+1cKOLi+CI0/Q7EaDOnWllCbk3/K1jxsNsi7WaTSmKmZ8UXesmaZ
ROp1er5eK/8gAGrkcbn3fzS5fSDWAOB+aJ4zbafOE9YhOAiWR+4X0I68/q98DDjd
ISirrcPab9APVxBVUWXDQXM+h53yfLp5Wys0lZbOrP9sq7Gbq6XDSwdEJJdJk3Xd
AJsex3LYcHHHIuEDrIJVGXZw7BaBXi/353Hu7h38TPli9Kws5qDPTwcKvhC9wPoi
+l+HyF8iJxcTQxfwLRj6sujrahCnZ+Y7Vsa+Qlmd7TZGZeAVG56psO1jeXLducLs
oEQYcpvnZ+qQ78iiHyz77ck0AFDbxe85LCICMoN4VLHDsdsgDbQ5K22fZRGuI2KM
odxaXqPvSZ4qppw7/YTaG4edaEe/w55qZSeyFwnUqo8IUihUKocRUagJic5bY6RM
o4sue6mqaXG5pZj0MUHC3HOI3oBW76eeRqwaQ13GkHhqyFnVW9Dsb3vjafEsg4fa
op2nbMb/ah0a7eqnXf6gYUEJZFgmK9IZNZreas+Z+cC5mNld1C0XKbqLpJXcvAld
W+Dc4ed5o5BogLPvO/nI2MhFnahJvnEJpF/7B2ZclFhLxtDEZkuhJg7t2Y/YPf8E
mk9YLqjodFYobsWvR8nSwh3DrnZeED2bLD7S3nJsySr8f/bzvoLcUiJANuWsh2r+
sDyWRznlLBjmUAGC9CBad0s4gy7Oda+G8/m0B8bKsis65la3dGR3crnmZkxFrV5h
yvaubIyci39lZNzFGbcbG07ToSk5yRoFqLAvbSLCUc6HaoXJSoaaLSDAvaDcmAtk
qxn0daxvHHz8As6D8g465YzEQhd23tH8sfLKSEUWihsyPTSgM52BaMzQ04us5ptE
zWspAc5SpMwVxX3cUF13/a4HT2KHso2Xb8quP+QT5LPqEMX+00Wn7Iulb+ItyFXp
04ObLcY3825p6ZVr8dO9KaMkqzf8jtO5wEgV8HRDeBJSWREqxG2nYBGZ4UtXsn3P
Q5mjbUs/o5moOlJgP37dFt/mnjW6nUnNBdYsFNYat1T4wJgOWH2fIaBcHoM509wn
yKykGzi2KOm1YqDOrqRLBbG0DHtc6XhJH39uwQq2BO/9FGy+LZojpqVLdFGez2iz
kz/tZy4ExsA2kAB5//wNCcLbjVg9HO+APpXEuuTYaXydFJHniapCUtdiDM+1oFnJ
XagPKEWg4OtlWHChSfCTXBlAYOLh5tTiBZ2QKnahUdxLBv7ZCAM6ukf5u3vYTrpK
WgD8/RGsQPYJTtKw1dwqNV8BUWZfhiFVX4u8lfu8VQ0lB3O3mbyWF+VjIkyUMRLK
1SHO0C7B3QqWuuWCacgDrQonNtZITistTfSNinxPY/k45t67BwDvcZM7xpzIwo2/
lCPher9qh6CRApZIYIlHXxgLPku0UFtnu4qqswsEcbEmf2vaOntIaSGxK3GzZ/8v
orfvYuPJHeZbj/IukxrRKfvxaCOHjFIzqgYP089tW2a9+9//34tTAqDq7jyc6E8u
bW9SZ8W3QyqqsiraUwnQoRlSV7ss6+3sJN3URp02GEmVidkp340JUGNEy0ZXYoRQ
RIXrQinA4EyhjjoJPv9Mv3V+Ec5PlVfOvLrogYBAmDg1+FRw1th3ktzh4+2DBeAM
54iYOD2Gz0Tc2VQkA3kRFj7+D5yXE7aPLvEHs5B/ai1X261zbl8GT9m+wb0OiDjX
RAl+S44BvvWeHEwDAAklSw+CwYYKO7iQE8xxxzA/hgir1BkhcsTR5rhdA18eN1QF
AQAKZuKqVvEeE25agyFkODlk+hcHqQE89pXxttE26Gm3OMGc3ywp1OpvrEj0Z3Vw
KYBaWv6yGaqt4xejXdWnZkXFD6nOnUJ064uwI/t9ZFFmWS6osUKQyA3Golp5E+bi
4Phso02djRyDh6x/CwDrwkuRpWB4n14GUZnuhB/lVjBckwvPYWg2jUcoZXKz9lI2
`protect end_protected