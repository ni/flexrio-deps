`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2128 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
00DMXaSvPYDqrb17AiDXX2mD2h4oHK43wZL3OfRSmBp6RIIMXXHKssOIp3lycCRW
qdGRBwVRZqmSzrEMmAr/CZ1u+b8L610X6JnoznYAAMl/8fMaQAmsPqcBmSZadU2O
Zc+CNlaXKCi1lY372BXnLjFIGB4r64HGw7z4ZPPYB3LLguIwzuT1g54Foo+NnS1c
8vFIXLanF5/KUKK39m1itDgGc8rIuEiysKQL58T/Mc3omTN4Dwh+gfOQig4R1LxM
vUPok/YXrlD0a2GfybFZT5Cy16zEfn54h28X31vn0EOrvaZFkj1d6dr+oHfCw0mi
YuN/UHW1tVb+7iSkTCe+HJX1sCZlG6wDHsY3xs1bN3CaMp5yCIf9xXdPcJHW9LGR
UFU7epeK0/xg8GU93S53lKcJexoos4r35uT+IrVEjkhpAlLNR+4WYl/idk5eYegM
/fEGw9iJJimxKayNmqWow4vC0HVz6NuGkUZDAHGToWvul2lbIbF53wcnrr3kIVaS
1fw5ypHJOOYe9y29FLTLNIWP9CdKIyudHQ3NKhJSfVOvdK7B76AD76C6ICmblYsk
zI//dSntAS/kbj9sRc5MTzWZRYz+RV+R+ZVpYDp82A3UkO1NZbKKiu6jLpcJbEcZ
kSFDoSppQyXFXBJx7mi0eu8OUpCEwOegvOCl7vK1xI/g+WGnrfhEQK8yX2kz2ZYk
ErqImJ/4akcl40hgniHaePs0rP4Z16or8k3J81nnRAVXDNQCATr0Bdqp9QxPnsG2
jIsCiZMccXUx3AA3fNvWo6Ilm071qY8z/SIMvrZffZ5R8laoO7dVqeyCSaUuOOfl
SgjV3ME3LrRrQwOxKA1LmVDob21yZzJ+PxELr+hqEmaMxtS778dtgixXC71/H0IO
nakafFirdDw9harqcTpP/1XW/bXb9tCIAwTNmA31XWQigs9sT02tJuzicK4j+xr6
icMtU+m6iDewMN1tZ/HSqZ+vgyBkO4U/a6VuYlGRJ/cmHjBg2rHKZxbJEuP97SDW
NiTeAmtHu3jSjppJ2xIyADdw6B5dUWIpbsEA8QDVhp44XnFZXYpFcQAG046Vj94b
AzqQsvFU6vKPmavK2PI5MSlSPqq6HNrAczoFwqo4qu0PeCS12ip6u2lkqtgHLxMA
PCABJbkZ9hNguwAc7WY2Gforl0b3gZpVaMMyox6NsewRPAb5b8iv9cKKl9kZCggX
fdXTNjx4/raybekjaQy2v0XkXzbEToB5u2xROgsBVn0CJAJH+ygUAmLnuo4IfwsR
cOdOLvvBqDGqxwypZ04iMzYjA4FgWA5U3ABBhzPFxmsw64JBbIdLrFm+iu/wERB9
S/qB/QqbsdSOSdoH6XWem45HHn3hAx3O1cka5CgPDnj46QEVlihQG7CDPjtsOrDs
J42zlKurh8jjaJDu5wgsEG6cAie4uAexUTKCDBVPuNRrAx7gKqUkAmy6aKAUC/u+
kzZYZOBnXik5X4daOW8j0uGCJoQZUVPEz8AslkWc5DurV5F8BfKmgsmr6gc6q3PT
iIHdOM3RCQwBR9Jg+j1rqK098QZhaqCwFByc9IVCBDaXHBwaIsTPExCQ12zs+Tm/
3Xkv1Yu3/UH6h5D8VIreOVT2A241jt62D2RgPyW3QrAsyLimaqBVHQPMbvKH3/15
QdeY221U5irSI+6TB0Vx/GmdMiPWls7fYbFNUEAJcvTY/pF0LOAy2lhosOZQec4o
JggEmzxNgqzpUqBTxY8Q78oidajl0qg/R745PRB12WR6+Vrq4Y5VDxXR2dmuM7Mp
NxLHLmP9IRLhoQ4wnnxw+r/Chn/5mAxckd9HMHDNFA1s6vP1w/x10mD0tAOnQfQa
BZQZdlmQ5BhZquXacL6ku/Gv6rhObhNJrbwkZD+tcg+ZWWc/SjaqAKrwsmIYFY+t
Zer++JW914pQoiTeBDfoX9NMhZmAlRl1aYadEKz/7k7EgKyLcZ9gmtbtjvMnGy3q
vZZfUAtQrhHbJFoj11y/XLd0kMRB6cv9diVLwOznnuhOW6LJS6O4H30eIF1p941m
Avh5lwfZsT9jbAXSsuDk51uiTTVouWW3kdqexw5j04OHn00QrCE01E+apmGn5nhK
97F1Aa32s7m9iHFQRAEpWCl0+w9TANU7+Q22Bp1MjnNGHq+X6QNLUAUsbQiv+qXj
jTRWZJQ2EkQNtXwOIOA6NyjGkjekUbFuIcT0S9mtOt1cISVus3D622mCFWLLXD83
9uWohavRI14ABwFHmJoJz0l7g4uNzXGaAHzY+vMgp2fjTd9MpyXXzcLB+ZtN1Cry
42I5NUBDSQjB32S0yjM+wzpMIy1ahv0vbNF/hHHVaP9Gfg8jgpeDI5lEWiA48da6
fKbfScOSEytVd0zwnXS4mDtWfXoKbcd7YVpNvqMU20CR2mxtNri8kQdOPZ+eLMb+
nq9ZuKvrQmGclUDtdJXmNnciJ09029/kGvBlX6cpb9Xj1RQyCUcZQ/kXBjfuBS1u
LJgIOtV7aH/ko4nqoepd6Cf4YZrsRVuB6c4hHmOBDCBhdyS4tZjIhydrVn9n7kWL
4aVMrIqG7TcV0KPoMZNdAmjDCbuVp9t8YlgBMO4xvuHqUp8yu4MrtRMKn5ZHXvSN
2wksSGi6ca1j/RGCK6+3re1uHcMGkF1avbVCRiMjnytja9AMEanp4rWCHIPI1ASr
q3EvVTGFefJmkSJXWnAWzQ==
`protect end_protected