`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20320 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTLkTmGIPhou9gzYhuquNWHaQglcJPF2HHF8re6T0msPw
MLd+HKnk/7Xr5auvEzc/g0LZylnVdAJldUhqGEOUWN9/KTPq+OtPqgkLGKUOmG7S
Z7t9j0sv2PEXSTyHpUXoQenBOjhxPr0dcAASNwVYShNQdeefFBDP4K9+/VEbwhs2
lk76mUyf0ZydvgoGwVhCkOuu+jHOx9e1O+DV9GMOjsOOnuHo4+3VjfZNKUZFRBuK
dlbMh+w8+od5v1CFf/pANJa/PivcvvChf9fnTt6z66MhbtAaxx1pM4652wii4hPR
+aHtTORU9B+5oqTkLprl0R7pEDELOlxmRzXz4+63QS11ttvu286RTSQc+MYkX2HE
V1cuI3chXSpDQJIXtX5C3GfHB6gPZgDxi4pLeiTME3nPWMkxA4SiaDAJjDfAOV6K
iZo2wP3dr1gPED67xmDSYnRgDDG6Z2q6LJyVfppl1jqJ1M0SQcyqfCW7iXmhj7aW
tlOOUkhx6wp4sUpaNMy9sxO0CirpG1Xt/jkOSAcnd+FK4TUnaNKt+UMXrVNIBj1A
1ERW/LpzgDQypSYLO56tsBKPYyQ0Jvl8Ht8Xik5xF7oYWIJcbMmTiq0ncQmRUSCh
hJNaVqIySZmuNQG4evPlKpm+OfnROjCIwDlMId+hxKBxg4/ihpVR9o+xk6IJzYAW
7C8Nb70nlAziTEKB1utcDV/iWp8IRqQomwJWO1wWH8pE0d2yC/DhvYX0l0d0JEg/
07tGvJam/wzhmA45lPUzyPFCnblfwizqiqtQh/nSGHySGn/2wpb3N+qn7843Janj
dIpZEPdmsw2dwZN7AutPLnpDq41EJ696J893NrqNu0rXIiTwhNfvJmz4DY0V+MIh
WlttVd8JSvQ9BAFZzHHwMGX+1o+UMJMvvPuM549Y+/OtTjFN3r/8BHx8Zon80pBw
nRqKdABDyE+tefP6MTHdx/xTkougDj0t+gvxE20usJevu4iqqlrNl+ev3fVS/MNv
8giYK+FEjZp9B6wgXOZ26gDVgooVQDSU5irHLEmoT39ESHsjTprWTsEBK+OYE5Ws
4tNycC4wPfbCHpUdHumGfFVpzXVhxYkrBtUMpzsbTGibAVLwSXoYzND2rJ8XoSjW
oZGYNVfvWDLSTAA0nNkLy+iHbb9YVbwYzFasHbnU9fVWhRQkieAq3ArhOIFM/Rpa
StzX/1OvZ3NlHgEmn8C6PZPc3Zoj1YHsOdf77zSnlbjBdX1SRaRQqn/FAXO2JyYN
zziQM0FBEUvCj4yTo0NvZeffz3BTpFC70hhYlRiYS/hfqe2LRcyyXhQwTTFRd1j8
jCmxss2k7foMPg63OrZdfVQAJs47hQhNqaEkmNspZiBT5H9CgaTEf34KvQV7x5Bq
/rnN7UwXTIRDH7yYGu8EovDvEuiYfNKkfAVomcmXxP83kka8FAKLe4Zo+8XNlrG0
O0XHvs9LstXUHGLAQYtpe9zmmGcRHWK+mY4mzO4WwAijUrQpZmCRT99yVOjAEV2i
0z084H7LicQUtz0jj3w1r633sNLReSKb9/20EyCiBl56VlpVmlmsyAWFd4trzjwq
fC+n8czqRixMuVUSyp/OG/EZpu0JmsPWP47wSTxMEXgUbmCBeRRM0C5qqZO+A3Zi
yPZNhhbh0/Vha9hP8NJyz9eqHYZSO13jB8RAck8XbH24Ox+mafRXHg2TTbHw1s7F
tss8wYn0Xbqnu3BESXXDGxvJxDuKxLDECr0Z2v2OoknBhFu7j630F6eDIe4I8rPW
l3PbyDf6yga0GBnrKi7o9WQr/mFZcDCJfO150C8xomo8UPTvNdytmQyRdlpuuT0k
L5oyFuCBP+W2tJvncw+0kO1txG8c2EBOKDaImRNZo/+SLgsmkQ9BWE319S9c1jTm
MaouRRtVkUzgz/ZTx/1Y4rgpie91lQuJhBU5iPH+I9ASq8MHLciIjthycLDeseON
/Mnfmm59TRIn93NuJzRQ+FPrJEEO0ywxIc2wcO3pOjT4wZX238KPNqIdgjUV2ygD
Mb4Db47mWNKK8k7lC7VWZDLZQJqXQY4AblKCLW0mdX/7XGXz6L7deXOZVtvAmeqA
4iTGRn0IyYhodJnmk2PLgUdls65cyCrJMTc6Lh2zucrlHmoIWeBZwP0s2bPSTsZq
2COa79Rr27CHpLrQAiTO6CtceYABGtmK+gBtlxNRzMo0HTPOw8lLbprW7k3jC3uC
rNBayLRSmzjasIW7rBmgJSy5og+M0IzuxZ4K0HSXND+cj9of15LdSEpXic7OxSJ1
5/nydFOrd/sU7ackDEtJ+fvPZIJFLhSSnuOcT/Tu1dTJaJ6H2/9sQnBvv7siV068
0jdHYMTLLNEZRq2Q3D3zXoth7Wg11fc+QEg0sJBxTAi7c3e8T6qYRolbcWnmLbLS
hVJEY+KIviQVFFFp9FJPtwOqw5pgV4Jz89ndXle1NtBk5yAp+hw18pcIz3+IZiv5
dwGo02PLcX1BG5IGyjm227iYZsr5PoXavYiA0bbbMU8Fv5Ys/rOjDl/PLiE8agzP
1qeFC8+s4lBu2/LjWie9wl4Ny93QxLxbw/KdOC5/q4QDtI/d0ITU9HQG+z+2eujx
wn5rnwGfTB2BZoU36kuIqncNNGH20AfePnaDpgtBNFEr1gqjRi98mdFRzOHYjILy
aWWMs6IIXCpJt1wz/bFdZSbeflvagCBqO2QGhToU+ZJtrEQffQHwCSAg5stTagFq
0TL7qnbCVlk1CLFyNsA3y2rcKcmVnPC8+qzeAXpXI5LhtKO+4WH7EI8eztVPlWHs
mMnKUyCTBF2tl0/wBuC2iceedpfA8KVNsuWRX7SPyoD9mp3U7RMjC9+LYszrwGFR
95o8ZpxeSfIum17lAczEDDVI3MVkeos/frKqVIqOrvDcMgHAG8ObzhPDIElHBbT9
QXj4Ww7J/sgSKeyTz9pfIBOfLOdKFpZXu4IThbw69HdPLBrhxjPhCo5Gu0OL8Ahx
iF9F8wDSuPwYt6IOuMEbsObjmAHwtHLIgkXgNN+voy8agaykn9auRjnqsd1Z5qT4
U7k/gNkWyvhURChS5Ddbym5tF9mHOtThRpmj5nxoPcbm6W5/fLnTlt1TISQWs5EJ
0ublR356pKjJpCI4pg3WCJAX7Nf9Ki0maKgf+mt72GRJ4ry4xvC/d9AUFhOQ9A0y
Y0TPvw6Up/Xik/yS34BZVEkOJBTB/JpEdXpSEguEQPOGDUeo23NGGvPCRZTLz2xo
W85sCVrrmgf4lIwvqztg+e3vFMAJD1+3eTggVnx7hPJDOpX26gPxnKxuGNGDqGcH
9GAY117qOtj69uVO88u9wn6AItx5M4f1+A5xPBrBCTkSGrKnpnz41YbmjtmxZ0Kk
My9s8Z+5q+C8RadJRZS9og+4TYry9efrpS2NWosLq/DYdt6zPI9k7lBND+IzuYD+
iTuVXQeDtEm8LZgahaaK7TPeIFQGRzmRaSgWY5PtVAXfurc1APXFwoFqA7AwRE7/
84roF7We9F7jwtrYGD7VqR2GqG+Jh3CiwHNNvk+isMeXXs79y3syX2mFl+yt0vKa
xH2HC97OShSZUfs2iYqfC+jbYP4rpI7UueOj0FZQ3e21nC8cR1VhnvHQy1XLywgN
gHvd+zPL/5EP0RsPt4RNj9fXQ/sU9WDVYa1Zvzypw5QE0qLmgx9chadmuhAXUz+s
HTlH/iHLcTLqfw+ztUte0YII04BcuEWbV3D9SQg83yPmnLNjsNPnG9mjRySOJmg5
1aEWU1tEVCS6ADMlfh7OumGtYYMUmCUsHQIVrYfefiv5hULl+bdAORtMh7Cizotc
fYWlgJ4bJwMQj7kyGqmfrsWBCmRfH1OTibCz5F3oN0MvBTWHOH0Ipvi0KWQaqtVa
KSo3HlqjqLjUrH3Dem7AoJYyJw8gCGqr/H8Xt5fqLAoKp/+6XoWHX/QAbE3gPfNv
MBKzFGGHe8by1+LeQQumF3jk4LenLv4hQOkyNf9XC5eSKjN9PTYlDzGuFN0s7WUt
T0y99HBCrUKn3ICxW3m7NWAusTNlMbtHjor5rUUU6KZXVyERcTol5SPRDfY5EjF9
uNr2luExeEWJ6Qx838qM3CIR8D+j08xlEldgmWzDdq2H7soTBttRlwAYkNOBIadW
gA2/yKX9FRxmqbInj3ByPl9eM46GUhEmY5EaJod0TtBHckf6Ka+ZsM2NGi+2jrhp
ya1PZ1w3PlPaDKjff8F+ZRj5CE1d6HVssVAPY27+BdcH/OPFlSZCFqAxUbR4MFN/
pb69sCx3V8nRjXNPmkgC8vX3YCya5tkZrEOU7qvmaNvtDdi0KB5TytTvjVrt8Lgz
KU5j+2+KcaLv4gDB1rO+ZZGZ6J+LyLy7IHpQ0nq4QKTIqTZh2xHzaPZ0EaRUk8iN
WxZ1tbFnFQ0FkdvwlePFhtBFMic5NzhACcLNgchkbNbBvgl5xni6IjCtgEbr78Ii
6Xt/FZDLbkp/byvpU2sQZnuLvg+wcnwLbOCAdxAfKhA3hxX30snkZRtMoJXYrQwo
5IBTHfKW+Kk3VVi61WicGVRbxTYg7XxP7SPyDgcKNenP+eFA3/GdxCz1BQFnpfKD
jKiv/M5tdnpke73YGrR+WlOv8AMDzDxCcw6BUP8abcGxT0qywlhtu4JXEB43PQBh
dMf2AGL+C0bpZxN8CMl83PdYTXFc1No8ueCbvOjXn4vI6IJaHtER3OmNquM+EgdP
oeFMEBMInvJcm/aL27U5DsYmLbc0QHYjVTpZtauKhJGrgg0ZJb+qJKzIEfFvXca3
WDi8gYttNAkfdRn7Ki3mbXpGtQ4+NZWgkzvXbfMgd7yNKiOgZtgzLN2b+y1tDvLM
8QgXYumg1ItdsXQfrXRRsbxaYKhs1gU5CXsMyqdwVqgLaP12Viuk2lJr94Qlmq7n
sP9XaOkzXDg+erl79rsT7WjogDY6+LeF74pjeiD408KwFcbUUIgFKfow2jgoWqoq
+PtOSvGKBJFtujXDOSAQbO+4/+AJ1dWQM5tQBhr1aUx5nk+lSyNIGwdQ/3sL+a09
24LKAASHXExage7MZXhoYaObTr/3Ypu4T8hiRVViRkEayutWtKd4MdMxUhPP9wGG
yG4sp25P6ghWAGH9RNhCWELB2RwNkXWgaJg4Dt4Hcs5Q2sqLviN93qgPH5v/jk02
EfaHjBYnv6lxQSBP/K0upf6xjORs1QtDRP01vYUQJ81NEovzrrPhVAOvX2UXczmM
QlMeGslFLp/04kNs1S+m++s1tpfrkLSbsjt+9byu81QRajidTzqu828u1Pljihvi
58q4j1SJHm9zVGc9rmX+/85yWa0QEtI/iW11JmZLSoISYV22JyqA9pAEEafTqub0
Rr7JcW4cnPRMQaAvl8AdwGJIzKagiWOGUbdWlDz4I3TuFY7/M5u6CODoqip6qNmn
UN3usv2icuvEiiUE7urbGa7QbHm49NsSUota4X/Qfuiz2QKUu9Va2idFe1kUnlOD
O02iGMAjyPGk0tS31CD8r6DEdZCF2BHRJA99BE20qH6qp2qaSvBqC11wzCEG+dvA
QJcvwCXF9936N5sVYJ3ACY50iXKu4lS5TNvNt8y2gJcvWoDytNg/hVMiJecH7fQG
FkW++Lzz7Da3bHoTt1890FQ0zm+ytMhgB4WeJ7tWivAVoKUWsKemdp0BxMYELgOO
mvPwzU2UmfCyWSp7qHoZZG6BuRyKt2tn/VBkwfcehp0sXShoBChc/mJqczhpDZkz
kk8b8owAvchhfaPtOd/5XrKe0Bs69TqdKcUCWtA3QxKgyucyENwAlaD+cG/Cyvfa
is2DNTE7Fs/otgw/TkK5aXLNQQDEpp91BC9/mkOrEnPfy9i/49LNHvpQWaErKml8
kZBmLbcLxBTAPCpv0Zcez4X2f1zFPgsSS51qiSNmkVJPCt5hh12vHVaHQkSH9+Ra
ryj8pMALx0tuORfHqZuSyR0vtHC0dO7b9GjhNxuCcaMs5UIXPANKtqdcQgXLpLB1
o6YrLsV5MjInmbDVm590SXRWDSWi8EgGyyrQpigZ95DsPMOuqgsULKFQDscZOsGq
LgPS1sqHXdykTbYbuv+ZIZyHPMMsmqQwD3XXVmlYIWcZOEY497OKk5Qz+mxZ3PP7
ssgqSSqTyU60h3otT8RuiqEjwLLbpv2KYAoKup2i9mWY8eAQU3K9J7wumW05EvKb
S/gpFB5q3BuZgRVJ94hDaIVxgRAGcSophCtrLIaxXG/dIkUJ27ow6otx8yk5zg35
ub9tAWfrsWMi2qQG9znuu/pFP7vr17q8WfxMyILWqOISSB0qmdzKnTb4YfsFcE5A
C18vLgbMY6xphU3W1iyH8u6qj5UYyDPt0CmaLng+4f9CeWe4znrNzsDvoGm8isz+
aX4qOu9LfGPjhm6lkj6BL9oV9Bk4aZohVG+zuWzB253u26o7Kp0y3cGhRu2DbaI5
9sTa2lvM2/u67wT9qZ/baARB9u+Q/jceQOETecRy819Fref0+mQu5YUq5uf6km5l
Nj2b/FEZyQ3QU61u2DClpBg/BzRGUU1NReOgTdpDixwSfFzEICfxDQSkQ/tLoCDn
V4Tstd2Tg2fg2395J7FOkrOKWhC/BMWtCiDNpf5S8DHxjrth3jQrzrW/P0ShssUd
Hg5QHDXEwx4rRzoQjp4bSGmmNuYOvb1U5i9UPdRLBUenlKcOeuIBmYJkX79uyCP8
sXAdaD8SdKfWhe8qtHSpOlDcOB14V7nuT7XAyavIy78f6NvYUEVbjDq7Jr6PUVTM
UP2wslxCbUVC8ycOgmZWypou1+xQa9s6gRep3p4uawVPTV+2lnECHKxv6K9V86jI
XGYzJ1LimlXBsCuTsy2YVuspb40eMznaj8E19jI97ciMCXowFHmk3XlbpIEoRJfj
Uw50MdV3MpCGZoWuDdGwdeWCCrL2mmwMdghE9PboR2Rq4zCj4AqJMTn//OkTc9D0
8UimWs+kPMlXgKUJg3ZBoLwmDb+2oGEcxtVlKno+TN5IJbZwY457qujA1dRbNSnP
IBZ7VlVqaZZhCvLA4KIqUb3/Q+4xcTjXmIUrR3sRV6bdWEW3w/D98uL943t/RtvU
A+qeEtD7xxtX2w+NtmCXjlz1Y/oObjeP/pScEo2uYZFDAxEPq1QOiZ3rsM+yBZ7v
vXF6PS0qQafCI4gHgXSJmHG3IHuocYfFX+FrT2UH2rNWX1pH2U8EV8EyZ8S5jAE0
cRhOv8cs4HfH7OUUTiqrMLuF3E8FKcdrwtxLNPDiQZWM12DXKm8w1C1/ACMUoJpK
Vox1nos42mfWKV/jHMYWwvr5vC4Xy2eaiXc5sTd9/G7U3wxElAFRMxGVlyKifOBI
cG60z8sM6egtFouXtg56JfnzyZ1n51N3AXpgKKGwIsPoRh/cDjT6L555iGvDJSnA
r7dL2/tHAAAT16/SBrpU6/OpArWD/xyLiSPdKQJ6oKXWT1xPjf2lPYU4ULhnL7vS
fbCej9k8deCOGTalIc4YPWUCvv1BJOLgE8o370VdbA9VMRhlJI9QwUIJFb/n52tF
fFvGRyAkRYWdxAO3snjmxdIj7qTBsMpugMzTfgJhv2QluIsy2gocmoIvbKzc3ECf
NqNOUZauQyoFmyZVFbJ0fZ3KS9M7N4cF5bNuiM6H7UR4vqvOhN+9W00Ti0JpeOQe
CuqXjbTMMPR48VNQv29+Yj8d/BpR/7c4gbqOqF/yuKHkfVI+AAo7qs8f/FDuTR7Q
xbXgadK6d4UPicGQ3IuxRMdr74LIj3vHIeJWCARqyKuDjqKYta2eAPFVAoNZi/bb
cHlekx6rObEq5sGQHqlYafJr1ZLGn+IsT3OZMn0suEqrZsNlATqjhY0B0GcCyR6h
rGjK/gmur2PeUJKzBXK3dsn0GATRXJC02kmxnmx7XFYVd0QvqdOHHEwN/8F70ZYl
q17Lm5haUJBXsPhdvVAQRx0OW9pmbDhrMs8UwCb2Hj1emgZ8+F9OjAmuCk1DbQBC
vbfvlE5nKkBCPN56aX+qOq7C4ZQ3Vs540VCqVDnX6xPNzrIIM86r5X2SCfAePgPQ
hjYRHCZVwPQGyO2Tnlar0XPoZ15TNupivZ7cY4cOHxAEn+Wg2bx76bnS/tdK667W
hQSB+KS6ICDjGPdAWsFr/sUtA5omroYQrG40/A/l+A7pta8dGBK5AVXYW7UDJSH+
VoFvfwA/GghNV0BTXKHiL82Q0/I64NkoBkzEUdKChtoaW65tKHsrr2xTo1fqT+Ph
c/sMG9Bp7JmM5jLgTjsok6UO61X6Uz4KnCQv5cUbnl9/JJbNmAQEzQD46QYgu4du
T3aotRuFT72X9bx9nHbypBpE3JIwabIYNTAcroCpf7bwHT8Sdfc3nye7fXOmyra/
YcD8AbjsWWP6E8U4NQBbcs32m/qmiAiMrz9Ncfd10uMdP+ZCr2rBQRuFqubegxBU
O1BKNVAjMFuPBHKScp2DUy26cQaJFOV8luHX/4xUqJhqSdKcSdkowR5IMcJZ/P8M
nohS11YPe7H546cTZgA5O2S0xPMNNs4VohpSgprstwUP+M0/V6lvXEDo5rx9a8Za
dE9EpePvsi041Tc12YKsZGcdJYDuAB0ii99myxZjIP9NVfbQyL+s3ncWNsygeBAA
oBmExwmA0qHuSRtyByKboUL42LrO7tVernU+P9D0UfDOvJCyJt60PKhMHiFIPUNj
uBQ0ZsR4QOiWoH+pLOUuY/J1iIZNvC1z+ZevYg6d1hyoJDzAVJ2+xUX6/US8qDB4
Xd3j1DP7eRh3daaMgEOnU/OY9WHMUOnn9cngigrDgYUVxgx3vgB8R+E19h0rrV5H
dqJuULyIxf5gIzrX23A7hDOWitmNzuXF5r9CldWUQx1+Oiu+a9iqZuiuttbh87kC
gPdowkN/FhccMopVfK4cq77+XfUKCnesO3eCMyJzQ6LKAV1YIUBD0cWFQUDOnL28
7bjcPYhKzwxAzqIx+76+UWcBQDJ6fQFFYu3/gvjDIKdCdpcAnoQPjMTdtLWSmezd
3ksRfYxn0MoqQzfOrrS9eAqQZC9wvDWEN3ig1qTj6nYlJH90l3mwVza9d483D3Ol
XgVAlSnUQTmJzTn41fvjt/jTWOqHWZ2o4zeH2RkQ16tjq7dxkDk6iBSAeY2eReP6
ABd0XmXKxy683VVcbsqLnroOts5V8iM5Sz7PqPWzbE5eiJF1VRJfu+QzKQBpfHBH
OD4vz7oRcSqUUhansSMajxxRqkB3ZP0eU4V0GfU31dRuXbGmNCRFMNEt4ZRomDcs
mRIBJL7CqPoRtjrQWHOex1nfEUXD6/AJonxi3z/eMnxS3uhU2Uj2nKtb9DIQ/NBr
sgESlX93nxF0XRkLPlrty3pDutHOOyNoQtSmviXBwQOmnbwmmhc73IN83jYcusHQ
JsJdSGqlC9+4AX/HA+04Qup1I7oH4ocgH8nvZ0+HdLcJG/11uW+Iz/ZVy+w3/HKB
444r4ZNd/iXyg3GU2rnhbuA0moLQaIUizJYxjRPu+zXwLo25k67348Mq2rORrPeH
iEoGwIvUdPk4N7NN9W2ntAqDAkmNuSNx/OtG28mC2ufvQXAAOGy4kS3mWQj8BAtE
kcbPeVrOi8ZVeyPLidnTccW3QASoP3Wg+5D8cbb19FkJM1br5WQV2ydf0v89RZnJ
fZkC6mJxJoH3WlfC1ERNfOHD0QkxOvQ95nzVlIjemYjwArfJ/v9EZ5FMLf90C7vK
1/EWyfAlahpXf7Ir5rpNi1Fi0bHfpwQCXB6kMbXjHi2BAO6Om4Ot7qUEuoNAzoEn
uwswagchuL3/6FBFa18hTVlxHGKWECA6PzXkPHrwES2xoWKnZ7Wv9MqPWZB5zR6J
9b4rTIlNHEK9jQLyBCeGvAHvILt7U7vXR4S7sbF/vnuR4zW+5FQuWXX5sb4gdzLk
rNt+xnfv4xqqff+aoF2B6ufQ1pH6UNhqpQRlhHpfd5MkP312eF1dpmPNzBW0nPu8
i19rZ/qxSMCufWpecTo9k4nOGmPhHnFp5TJeV8T/n7Evk6W5g4tShE1RUj4rMR3S
Bb5XGN6AqBiCBdSVTMqf+PNGXqMTkkgOK0WK1EQA4+ZzZyTfMY/pv8ZQT53579KU
jAhCFvHrVuM+BqrTOGdpWf6RC7a3gKauscbBxET+PBHPHSSYYUIa0+W6SLY6ABDq
WJtV/kIazlKb8+NXqVow98uoxfxdzexuinamp5d9XLBC91iXdXAWS0jZSO8FCbVF
1kyPVNpXnmMbzsz5cEDS5/uFxaDRyqITSZRfl35tTHt+Z6P2339+3uKNupZtRpyK
v4zeWpvWC0hWPpmuNG500ekesCsa741spMptZDCMeQChutwvn0mRICojpfipwi+v
Np4q4rsyjRjdFl0aJJky1SQSRineJ1kyK6o2qQfSHUCJn+0wJ6GcQDGjJtY8ajMU
wh6r7I5VFjUnf0juwoMDFqj1yahZuSGm5zR9IdPvtsgFdRIwnG1W0VdbUDaSzEPj
R+J8DOpPCQDLBJxlwyd7yaDow6MYtQZ4rS7iIAhcDGLJtLnfVksPnYqOfCuJ0SUK
LfSH0V2dglZWKkprCHZ3bx6rQJ83XC2cz3fTx268ZJuxoHjSgQchN6z/8bW0+Gh3
TwQx2r+zHaU/kD8PFWEhB0vmZ649pOgwUlgG4TVn++S5xDbtGYgFBYsweB9iN2vn
/BXrogFMrufwIsrU50bGjiH02JFFRQGY5K7xeynu9hoin75TAgLbvu1zG1dRB275
11S3Pn0CkuNksStbOnftXCI/xPg2GeWWVymgOAx/+OVb6XVh4FBLwOwoAfmJH0vp
j7KLpjk9Ezw7xrAIwZITUoOe5cMqctWqdBqlH0H0AfzbZbSiIL+qwjHtHYOB2jvd
wLZ0a5+4qOijLELUfC3an3qSj770+lXveR3R5f/YFigYk0/ajba6ph8MBYkCH869
zvx6R4E5ulDVNVcE7J0fxZcGFVFpr+LSSVXhczVGLZdOjPnlqQYddcSBStKWGm6u
RG49+qRByl3gcM7143aLwNwWo9E8OCF59Fpx1It3j40eUOsOjHGbl8y0ocG3Owky
+jW/0w/2RhFTrrFrsPmp3b1k02UvAHAx4O8lhqNSUjqNXxY2vESmsYvUn/UvDbxs
npjaMfzRqt4PsmjKKPhpPqKasT56CtDxV2/78xbtJAR2uCnxNWI4ucqZel4JdZiI
CHbF8/u9wHjLTLewjmhbSCnsxlbi3jDHs/OiYd/EMB/9zOHiIeH6/U2wSpEOH8pQ
ResoKKuL0QTuE2PmOxXZ4PsZxS/0HHL9j7zcwMwiy6GR0f0i42RbTNCcAcIvsz83
lfEct0ejquUx+6UnXmbnWaGes1tGLJabYFcmNLo486okLv4Gyr6BWVDKo7IAA2RG
Vi14DchR94dd+di+bDAmOCVFCyD78wIKj+yOM8Ul0k0j+jy/84Qzq/u7hlDDLbFZ
LLw2V3lHvODIpDM1uh2LMWT0s+6Z9lc8Kr2FQ+24YbwOB/QqDyYvzcbXbBTWlgVU
RpXvy8bw0T4cX05n+Dw5F/a37QqL4l9duJvYTQzp/+OMfMphmeeYbuvCmGla0Gyk
rUEKHKR5nWuZQLHHkitV7XsTErfkmoERd90epQ7bFWyBXKLZ2wKe8tsUnkMVGYAG
8lZoDyDGitwudoh9d0Fm0v/128B5Eq7Gkicq/14WlqgEupG/DRT0hiU8UpEcEul9
sur/kuvc9I09+JEGTCacdUdng+b+xzGct6gy9biuL9gtPosovybSpHxvB6pY0J8w
w3dpKL3M1FK5ejAccI8+7l0U006839VMrP72REroZG2XhPVGbjI0HQvvFXqphbP2
s7wPXS0LfMMMa4P9LRQpY4dih+/Nkejo64gu0U95cL0e55xSxLxopwW1Go2Xb/1k
N4M2XVr04q3La9h47j+O3xMBfJu9vwzcMvcrhdTrbX41p/H9ik0vuPngXs1uAJoT
gnhBBrZgYFaA4pDy3ans6YjDBiK4Zf7IlfEfPZOtEONLrNs+wcfDdhXbIfAUKMK1
VmxOBNiX1B78ijh27QKXA/RJj4r3310FhtTH80kOX7aaI+nZNy0QApT7z8oh2Yey
OPqi3ByphEIoi6YjdvzPJ0i2eBGbg4S9UihKsvSwzPB37g7JJu1mT735LD06gUm/
qddq/8X/RjouxSVWAL4vzRLXCkP1U6xmaIodOTEAFqAY+sVr6U7qpvcOHPCkQhbU
FBIPg+d8yTOsEvwSD3N9Wxip6u34iyvEmJwGT0QIogGLVysg1Ft1xHML3qZC6QOh
jFjuYhUgj57+UtVFLoOTgnlFzy/ZwwqMgGHPsHlY5MeDBMc6flwgbHhQx2mZf6cw
F4x03aUvNyKn9XL65bQrH8HIFYyEcmkv7Ukb7KOTytjvm05S2kFFrYHoZtDYU/L5
u4/FngrJVy7EpbYvmZmkNLAeMqqdYAY0nkhBdkHPw5QJxSDGM2cLSDt3NyN0wn5e
fDegiOyLSzzQzAgoNa9s+s0QCipEM0CzSNaJNvL0H0OO79cL03RuSZFbiV+x1hW1
Q/M7hd7apD2Afxoo+t+ysxd/tu60O9+/rAvvoVO7/iKCe2l4Iq+CA4J2we76lOXO
2UrtszyW5cDEJ72eqqZrFf9bhMxUQg3MkQNCMuGGzf3D+sNrbqshKh71Z9XWOv5s
9/OnbUtBEt+zb20S7deJlzMeIMPcQILEZZX9v5edkCj3Dw7Qn4d05vBeUIvI2uTr
NGyPBzecyCE+HGzXSMbC5sWYeZJ/lC/eMNXMKVgBvJ1NQpYdxK5GMEm30nEeYb1V
M6RatOG8j6zts78S/x9QkFbaFNGPX/+gg2CFhcGKXjC4DioPPMyELCv25xOznCaw
hCYbvLqmzHIi9MSaFJKlFANmOYuF4WGR1KTsZsQc9xIcxIrxY2wEq2B2Y+Qs7jGr
JkoYra8OHcAtolE7w7alz8ltEFAPU4ElMytBEge94VGmiQOZsiTjFpnDi8692n21
+T5RH9HjAZI1siRkIp0aDPkeeGTcStAXHgAByinpLX9rKqvLJXK+y2IUcVSUWwt8
/lTqwOe/SaDHVFVzw8ypVMPbnTvScstXcnHyfxMcG8PYwRVQuso0rL0Bkxq61QVK
YX90Stu3Hcio0AwUvP6/YF8+GaL+ArM3CqmkzjvhZxzpyYEdaVDFHl/PfYu3jnKv
hb5HWthmNoBvLUXadTCDrBPt1yPav8a2FAn3CN1WzH18C1o0IqI92ESfQ/fOvMvu
MLF82Fns7087IAgL9yCTpEYo3KAvZFKwaQToYFp4qe+ZAtYyje2odvJpfSXMRnkK
Lgk2WTpmgQsacy0hZtI1gfgS/pULci7ZaHGsaw/Z2OdGpTC3aDHinGpU7xr3m/Jd
2kJiem/si49+q79zkFHpPHe5NJaRUm+nesp+I5WjNAN36/uhjTQkMEqO5f9u/Lgx
AdtMgrJCRtbC4bGVwfLwFCBG8o3WnE2lzQfllnIS7hUqQNJQ7Kwkty98OoIvfcJ6
nhWJU2WmmnDRE/8hd8ayWx63BjhDHn6rW56n3RCHqeit+X8iUaa6yF6pxs/Gq14g
hYJvtdw5WvlltWswqsaBuxlNayGo/WZ4V+q3046By38qeB4f3VjHGDFUMtwtIj2S
V/VSrA/3s0k9S81aN20bd8LA4HEa4K0M3d+LNHEUmB/leLThyGj/6Kv6WsTSm22Q
HzjMG+i1ZXqLP+X/JxE1prf84suyMM9Zf3GqG2XfrZg/bmJqTcaIMp+1CTLxX0xG
BGkdqtTPn3WhMvN5FHAh3sMDuAWNLoHdZTvxXd3zEofiVlz6i2d6hoSuJe73+mpE
byRl+PRFl1F8WjFXXzw3+nHnoTInmE7/RbCOA6g9SsKugbSOPTSuXgGhzpeRNEuM
NM8Txoww90VuSS31y3khvT2NmxGkMn+ApH3vVapSta+yWUOreJbMGmYxAthi6y8i
Cpq/6G/w+Oze5ZIc2ce+IuM+PE13a+LN3gMajI6IV3LoJZgcfjlhDjmSYwZSQotw
yY3KXlAYiqvswJCRF3vhYooJmk6rrv2d2QMXO5fEdTXofCbPVZ1FqXH8NmSGGt79
K7D++mPQvyJGQBp0fTIfUF58D3/79MGFX41UF2Yx+Vn8YJPPGwFNw/jqhBHZLhAP
NGy9qydeQ07gZ9+WtgDkIHTCr3JI7t67OBZmnJQj9wtpfREb6pknwLtd/TIy6jcY
0Tz+QdB4VZw6+xuJ6cflAwDndT3JTeFLrpunDAFqjTBNooEZLZq7fcxy2Swhz346
Rlpo4OrwBg1SWY8TEOwhimWbvYj2EXzJbJGHVpVfoYVaaOratBdD9sp0IPkKlN4f
UbdZwuRRzsDgkIBszm0iPWVSmNTxxNJLTqISKetguDvM90uJ6k/wVoPsg1S5YwNv
fQkgEo4Z+0WdyyjKBBB0qB61mBoKFCa/WovrjmRld/1ysYNHfmSBXiWg4//Hu1d2
XeA1POXIxtJpg0OfGGVc1EZvqTtJ05wz+baDDk0B0GOnwdf55LA1OOmXvG7gFEAv
e8F+bYztldq6z5YuqkVDaLaGe+z35i9EjbmpsIim+27YNWn4xGmqK+FFM22692K6
xKYys4fYNV8uDH6bKrJdLOI5bYTWrtN/Ii3CzVreEeg9LCFWL/C5Nkl68JcgjK9y
W9Tb4GkXnlo6CIthFXkJenosALZbQgSQMYCSf9385jJaIKUJnRas5ldzis2R6Fyg
93MRT87dM0GkE/NAmETof3EQ2yoj59Zepp36zY7XKNOdozQSiKDgsV3LwPM5VG/3
CKSbraqNWZ+PBSYE0bjy4ygdI/6VH+MDKWKH3ME64DAb7yYHO2Dxl54ZxT1x5Vmw
5PiNmAvYH1kwp3rVFYv0Tf/i4nBxvL/Yv71eqGV/WTIi76JFhf7djsLrYoNZRlXw
FVr2g8+zo5Kl7AGLWz0fK+a8ANcrtevuKH12yrLzEZely1fH9u59GIizXKSopyY5
HPqxbzJvjXJd2kYlrWFXCyUmnwlBqotc3ivwEyEDNt7+/ASt3+eMyfuo4PqHApeI
/MBJPPIBhmwic27/SAeOczGkcZ4HILPKlv4JdiTfNWMJYtk6gaQ9ga4kP/ceOFKU
TFv5GnFFBaocOcVZ/QMZF5B+19lCUB0qdgKDqBEmTj0/zpbv3OoU8WZtbJPToJm8
nWAZIzWRvAuQ6a1MSuA6uaqelAruPtf2ZLd/UyOdMtlIZd1I/wxcJq5eoenSsp9B
jquxKdamz32riiqEi8MK3zrNhfItSV9ELBu7zyQ+D4egCGxO2LYL+GOZELdMCsX5
zqpC7RDHbMLj9EsqKxVSsJob6VnDdc5tcwuehThbc/bodbG9NtFsZHDADBrq019H
Nyv/1sTMIPQ8TM1DANka5NxZPhOWlze263alBIFaDtb8lEHoiewk44LXlpjzPz4s
5FDMHFiFtpTGvO1A54W4mLKHyk76futdQ+8jUajQR2KLq2nQjzI9CXXgcOeATVne
dCj1SWUgxGSBYBOM5VotPENR+W15yFvlslJdGH+uKIw4CRNyREVil33gGZoT1nq/
D4GFPgb81C9xe4L6HU+1beq//ohx9L42tEJrk5rzbksvmha6JnBIRgA5L0sO94d5
R9qkUVKUGGUpDC2+SbWQMxf9sDCKzjQ5+Xe+W63M0ccE2nBrGbHRyePKv0m+qLx0
QxJUYKL5/8/0c9kxnuhgDtg/YNNffHjXhNdeVYak5G8wg0/zGT1ng0AiPQUNR0Hj
P4VRmxqhP+CEKqu899uXPMrdnMBJAOySH4+fgAJfm/HxM3r4zXavjQT+deprgZU/
NUslU0N88qkkIILPRx3L08K3dSiwdLpe83ZiG2WV6eGsS5XwsTWRvP2HOYb4z+Q6
iZX32RhfDFqJGZnaQZSGnA38P7AGQ7u0qg9cseF8yApsAcpqNUEu5mpFolD7/IPg
6/kFUEQ5+ImQC0+iod9gPmExNchCrO3q/yhQlBEJZee9GMVYkVdihEeEBmOqOh9o
vV1N/Ky2eWVbiTOu8QIfaFQBzSKsSbEFEVXiCqh1iLrBq+6RMzpVyVo/Ghkpt3Fb
viTf4jAy+HnMf9XUD+6eckFYJ1R9jDMIijkKjZS98UyhGfFQoQBl0YPuAebN7G/R
U0V8GeALImCcY9S7ErZB0aJi5mMKqHc/hYCLmIwrFEZ890jriWy9juckjiL5jbF8
TDPA6P+BGVF7d6trhT/s7+UFnLOyaZwfcyCxwo63mf0bnFW84jyA/dtlkTdKVSZi
bxbNiIgcSc6Io0bfQnijtge5+Co46hTuld3XsPI7Kd5Ontop46y1ou3xVOpt0x6C
s6eUe+Igv058Fowoo3A0Tclra0Vogi+paUeonvPWtdkR9bQMnV21ej9lu+x4MMcr
/g9nZ0K2GXxPAskk1ry61KYzt3ztAodfW4fdDuCZ5eKMiYpmgETB9xtwaD/eYDCS
h1IYaLdzeaSmiqgMfJv/j+0YyiUp088BPJ931R7gRjFxoOEw6EOfAmJ4ZQvpc3wC
a8M9d+nZHsDRI6UCnkljz6HwEdM+Y56DtjNK0/wIe0TZYgzZjrGW5zSBvxaJz/WB
/8s3q7ah7i9Cgqt4hWDjFS8mT0Lq9pLM5Q4fGkI0y508WYKMCyLWHbS3S77h7YLW
q8NS+/1idkMVneOvym2roqVtr5BNamJgGGLrlyI9j6St0b0DvWJYCbWv4XXcZyxR
7HsCUmotMQywCF0FnIJe/tsafdjD9HVN31shoET+PuKbarCw6JvPOgFV/qYdo9f6
/VyLEW2S361erctCJj/jbDFultJndHWG6Ipj80ju3soA3YprDm3dtmRIZF59r1n8
WvqlUGTYnSFm0hz2lGOkxMziql5VH6k5T0JSnMKA87Apwu+YW9jvIKeQ4/3oz1YP
w17N+ewHqpMvHBas9gR1ai2ajkCxrIgwX9YA7X1gfIIoq8OJA45zYfbv+QTAhmko
rfmw+HsP3Y+zPM+ObEcYSRZWbHd+l4PaCNGmCI/XaNxq6asHUwS7DBSaZMpfSt0O
Y1Ks2sjonGrdQAOJJyc1mb8YUtfV+KovLl1gCOX48ff67BOWiWjje2fxYOGXAbKU
wpn5ek32gLJYrKMklkBRyqtR3sVNA8ccSnQLrukCOIoqiqx32NlOcuh/GdJxyk/K
sOlsZpsS24NIBvKbMKIF4hiYV6pGRlfv/sJYsRWMO/bRZmD9c8/Pnh53XUuDsom5
HXSO0hyPUInYzHGVNQ4hTZilycx5+/0o2JO973O3HU4J2PdefLRZOoxFgkmDuJNa
TF/AlG7iPj8CzRMdQ498B2/GPpna+wi34VOLg8YhJxXDRZAQQwGgxcMzmW+hfzL4
HhseAhJZI+/mkjbEBCvVd9ZuIm/b6zZkgB/VVmYS5jLeHMih7Ke/6uKhygOJnCCU
sSPPCn9DFmQm3fdSHtuGXEwFUIDcjDAz3+2KGYwve9ZgcSaJljw/BcXONCEatbwF
b1L9sj428HQJVIo9D+C5+ZxKXmYbCqhl28Pb3nPVatgZcHFQE+LUKSuZSenzxDRv
CBzo9EGeUrsXxtWht/xVx9XnZWsZeqpasDRHjY8TP6iltYCqABfGkYG0HqFvQVdZ
Aiipi05cpiHPnNfsRKPP3C6BMVqlXndfAPAGIO9nzur53shNrHLEs3hKXb9XWZ0c
ac73/tfK0TO58+lTI8ujW7l6VYNj1YuIwEYEtHHq3n4sfH0UL2CGA3AZ1gRSfoyZ
60iwhCSGSr5D6YY7VXh/iKOXrisQTnUzGIm66G9lqZ3ZyhCgVqHnj487XjLxwn+O
shunU8WSI5IRT2ykXsQT5gu1fcjNpNgd06AwLqhfRdbV8B/dlbMaecSiOLW3kNGK
o4jC/8i57tbmBbFdZ3xzMeU/B3S6SGWhpChEDB/l0ti/4POExhlPrABP3uNbG4mb
iyk6r0hTJPGRFNVcSRgPgJjzABKmwdGNnyvNOMEJ87D6ADgmMnehajnf6BRQeCLn
7I6QOm5agp4nLPM9LWKtT9tigwjav36xzleE0RomNn5z0sYoBQi50a3MnR6kJPQI
TNXtYDAD494+Pu9gXggMBbEnSQM3HA6Et0sS8xSrgh0CNiWXjaubgwqEBED7y6qy
5Y8f9uYs3JVwmJZnuimTgaUsBS1VIg9yGLeMMMsxrpElBJZchGUg0hcupV0y9pqx
9IwZOBEtQ+OecZMl2HVe8xMIE7PKSR7tpeIvPEdgEwJ/gXGu/RLK6KXaFmj99VQE
3GZ60qI9h4U/8F17KPTnfQ5fRDkyLWKSx3RvdhdMvw9UlA7Bi0qR0yXI3iNoiMc1
NgQomEotrk+rtHYmG7PAu3whoTzAosB/colpI0/OeUgLFsw9yU75722JRRfbLW3j
Brfm1qqWvsfVZRu3lmpW7FTnvcauiuZR0PE6MmBFs+htcUskWDEfCcEcPOPXYwVA
b5vJiWNQMguCXGurLqTKaWpxyHq/1uUN6wlTwmqFMDnyj7N7ry+bQnOM6G19cl15
FGKIDxEW6kWd2eHzpa5Gq7I5ydM6Jd+0tUwf6O00hsIZVMiL+0+ouHe7BsLx0d3x
fKYwoJDRDVC2PmhVqkZoJi2ivvLHZ2yIU7USDhJPWRADYOfQ1JP+fZBqT8/6E5wW
ICeJELTQot7ofS79VtibiPXXEv3mb8tGpHD7+ZTNhIAIiX7dQKRO69Kpule4rnAh
InwOcTPo2dQ4T7sSbNQ6HDDR0tAMBJmCI1FiG5JXBhi/XaxT532/TD7f2jGPj4b8
u/EvGUqRg13mlgAQKK0Jgz0qrd6lNmyG/L4+6GKzYkVQwPRkIK4ShL0XwKHITVGR
kISOlyEcShLn7QaXznZrQvRnKz2l/9sdkVYJUHZpwIXgcDIfdmfaeODHXb9TlGfB
C240qdIV2C2N4TtXcas+94UCVOieBUFtxxOp9fJs585APs2dQuMc/HTXYnjAsafz
e6TcGcKq8QkAZpc2NSDdo52magRUHaYwh669kkSTShlG/pVLVi03cYG3rEZNqg/i
fP6I4CgYdTzA5JjJQ4eK/Aq671UsZE3QcMFMIiLxEoALR1F3B2GoOqalNuGkw5zo
NZj7UJ8soyOabp95ICKB2CTDB0QDE/YCfQPOAVVW+opapLU7kRzrXm3991vntKk0
dWDaAr+LY4sU0rCY10t3eDOVcUzG0UVyTUKDfwKmCmeuPO3p8b/sY8d/ygU4Yzlu
1fsrR5bqsSBYTsW68PzkIarND6F0JIp1uZCMU/Q9gtQZmXFRY5CodS2PhRiMJCXh
fjsCQAcwQDVWiHmqqBkdOtjG8kXDKk75jMeeRBnbROXgaj9kh8CIkl8yUwvxWDh0
qPrbh4OibQf2r05T3E6t3Ti44ZpmyIu0HvR+N9SyHeYp+kNyipHcQ2EfFm1GF634
fvI/d9F5IK4bN/qRpmvmfT3gJXC9+W/SVrUxCf4KAKi1+OqJFP2nvuRoczxlvQA1
BODPtt6xkodKMQcAh69zI2Qon1GFcEF+cjU8VQiAKnFNmb7CziwyLYtRk56US5b4
kurfRbpVau/ge89IYd/Rz7v6AezOBBul/iqZZdCtx9A0LkDxPYq3qSwwByNls5gc
p4NsOsYCyi/B+i1P/n0B3BbvB3QtlmZX6ZRcCfGUUG7wk+6RNIb0g/CFQYcCd4eJ
naraMG2oCMfZq6hfc/XQTUxtdDdflhQUJ5BMJVzKRijrXCbDeI16zDAVtw1+wdNT
6W++CDqIjnGVpDzPt09DsmmKwTQryYfC8uuflU4cpx55XKNZlgzDaQeKUoXmQ2V7
4Ke3gw6Hxi/WclYQecQOFhyyftHBlA2MN+zVcIisCMiC4ValoG/91ggohdCXWrDJ
f50La8pYydyJ7dSTS1G4SJEEWWbgMrQURJpLrjo9TP6U3D4Y1nKhFOIZUTZ3Z4BF
8PBCKz4BbycRpwSMsnEsmcKDFGPnqcbQhAdsQoOJljSwxzhGsQZxP7HIRClMjCQv
mOwdhlRF0aNVWilOXEtjJPZ/kJRCt1B3RkjVpUP1Mkd1FKkAah22hvvlZCFtcm80
y1CRKW11eszOjQfoIwOGn6/IatKJRckHPLQfbwAHZQYPr/bhx4x4s1DoSBLwmqi6
Jrwn4oM+EzXwrRLAr5xb+wQ8MaspCJI8qMrhILh6PEpbXrPFkXP85jziJQZr3NGH
weFKpJIQ0McmkkWZbpkM9qzwa7v1b9WHbCUN+KOVRbhGS35JKOclmf/7rUwbaygN
RZ4Uk6De6OlqJYUvbcKwtikkeaGQXbwcs1Ahj8tfZCAiwmjvTWb0FhDbYuls7LcY
7g204HEnZsJnIMrL9Qa1J3LmVvcCSJtFwgeKVsViGd3DhMDq2kZPUHraXns4vhmD
J4kzS517hgNrUt+sPxrmMyLGy+pa/SDSdMyUn19UTtMSJcwJv5WYPB7IGqlVvnLr
oOVIKVLmu61RPn9//wcnASJiVV14EZIOsmcYCgTCbL7c2+CIi54B1SP2qOmHNHLx
PDSJTw+WGldIWM0T9KCWivmlzwmdEDx6ultWN6PlaadcPA/IaRHHGKH4+1jn1PfA
cWR4daExtA6RmUqD7IK+a7U1Y49/SGuM86qxyHZKwpEvF5zAHq8by1bCdykQ+AAw
Vg3oHYK6LlFQlChiElDO8nMeq2ePVZH3ny3Bq7szxvv+wIONM4sK4VzC6h50T3WM
rLLodN2m8axdQUdf9gn9+Om+e73ikXqbkuPCxh1PnZAt9shYs/vbvbI1v7u+oHka
mpTfViEGQ3ysutpCoicpNKCxbiwa5eL9Bgj4627i12Ow59tNXKf0HS/6LRCKiEhm
O3ibVAb3xDagfwXQAxOT+ZrtPPDeJB8f5MaL2jFHscEfZKJbVOYgXjv4L18d0b8d
gDzouRw6sSCtjhsuSJfxBGqPSN4OwCz/vWUn9hp5RC7pAEiluH2H9X6WKuvW6fOc
0bskPRkAfKRwfVkUjMoCE+M0ggOrLVl3HVNnYoGRS+UZkMo/DMiOvpUmjG139Jt/
nK7DwNdRjq/iq2uetkT+eFRjcLKuUwkJs2TZhjhzTTaL7wgv3plCucipqrYu3G8v
syKI7Sgc1C66gKrb8Xit+rv6VFcjbySKfR3tD8+1VXV/ipoNjwN0LsVncoSO8Ktb
b0LKK+f8PFUDFVWku7rwQwJhHdwnCgJJ/aMH6ClgSo7zSr3x0bb+L3DWl7k/j0/2
qXPa3yen0Simvec5BE4NWX7rt0e8yMZjAx3FbnfQcew8VRKAXAiw2Q1lZV0yWcG3
PJvi5jgDLSVlFkoqcJFm9cr1uwpBCjXVYTpY1sqXll3cWOkz5PFocQCgbnJ5gjq6
Mmazwjlu2mMDEDhG3JtHvulO1UUsEN86goYn3znsBMP5DIVFc9F3Z9h4Nry4wSLZ
hWuwwY5BvTVTt8waRwowm1xTv9ApV6Z7MbwTHfsxIrJsfGm3xB4Z8Cro9NW+VvL/
xzlhEtnEXYJsyfVoIMBljrrAuaHnRtb0tJiVDgcdEvTWj4QoyC508ewd544zDbI5
5bkzwu5e0MOsH32dREDA2PTvswP8kU/4HsfvD7vbZBK4Vc/9XPVvSeLMydVuvhgr
fIlb830CUHFCCzhNWhjsP6TNDwkLLejaVsRAcMqlLsfCqTOGdTbXSqzv0lmbwHG/
d29gYMborPJecKl6nyJVgOm+qI1djBnmCMV32yb2K9TFv6LV9Ipb1b+hzu3ELQPN
GpzgVU1m8Y5leyiXyZRuAKKnN3OdU4TvosYHZ6meC1glpad1p+t43FA1elmy4vK6
DHYV0DRazB7RZV+3xRmk98KPiP15evy6MMBGiLjM9GGL88iOQbTdsG2a6KDMHUzt
4wasBwOLBmRjd21W9utuvt/rfluq7Mip1app7wBu3PShji0CmX75zfCT42JQ2MBi
ft/s6j41ERQtuRC3Wg3nlelA+iNF/UdoZRoYM2SyIh36iJZKQq0tSHkWlwJV9P2D
extQfjRsousuh8ERxsUk0kSRr9RFNCkFDrQ4o7h6/psYHnuqbh8DdYvvzXUalg6u
/f4xIuHIxhBhyLea2ZavP8EPfrGKiICAq5QkIIoQunFJHDTk4KXZmVxnLDYDK6K3
gsKxRNKpalT1IaNe6EH591yiO1QKFaV35nY0h92ADcVaC0pyTTw2jagJNk1tuc54
IguHhX+q+Gasy73ljBny5uOgi/ECdrheLn5AkYWULHme8PZtASewA6qiNq2l8JE5
nyHydj8xOAw04m+AbAINeGTJcjzWZhi0bSZYC/IsPAs9e1bsIOZXBxA0Cno9hdyq
oUiVgCu+YTeQDrq28/dKjfPASbcejZgweDDDOjdPBFAVF6XgJZ44PVbHAtEau46u
4VIF5wbEF4ubq8ruhHrRkWTfmDW/RGwuVPOhSnaaj+bXGLONpriNqjfw1mNbwmK+
AyeG4a8+5Z5hNjHgZLMbicIZx8GuZvhFOUuzB6UxIVbc0j0NLiZTP+/lNsmB2Lnd
QUhU2qIBFjgJYML45orkRYlWAs9BHEbNX1euIH5hxY05OpPOL20lRxWrGUH8PJG1
ouo9pzGjgF7j+2QKvSz/iz549cjXoZB8p21fRAT0oPlZKqqXHqfaoIUvEzmT/Se7
4pK91qRqjicKjjM88zqp5kx+oA/SqGz2U+BCQMKIbWPyxXDjoZe89ZR/H2IQv2Zg
hdqLFKuMPk6hWdYx22qGWL+ze+xjaaPy1fzCRIfFp8XqZ+MEBnfJuaA2DM9CsdWO
cV+C9sa7rZ4VP9M69UeJanGPgfJ2/xDeSq527hKOFPZjFGrJf4b95cv0HJ0fP0Wy
Qn6lxTWxRSu9vl2RpQDTn4fcVo5K4+fEUo/zfMrI+nni0PWOwM1MvFtUn8FNEOq3
1bSMEdVvK+wAK40uETLHfi8h7vI8SU497tkOp6vFog72lVh14moLYfP6OzutA7G2
prSxUmJCbbN5iw4qTg1ai6x2EOKBWOBAjFb/dxMm9MHiT0AT268nBmu/KBWD5Aaf
Ntzdf1cOK4cEhDBM7N8LGy+XYITwvhlyTON/Gsew7RfhPa7eDFAK+7dvUzwGtsV6
kSFOAv+MWsrthgRJCIhMuC74Y+Iwo3+n0fsdAHvXbBdVlG7JNafrCTtbGd14mcEs
ex0hGGFd9ZzQ7seLdWz9c278e+sgX+n/akZ1nDv5/EdHnRSJ7/keR2lCSENKkJA6
gh8bzLvK7dIpwTu3+4IoC0cLCT+LDH2892OI7QBOM+YjjCJdhUu2zLW6nFGRGASN
/jyXIs8/qram4bsZ5Fs2W6E/a2bljLLo0IHatmt536TlynAahFBr4AmIJDmpvRfz
m719c2Epc74ls3ccdhgRcB27jHF3X3A0fM8wr7SgTl4MFDL+KGlQfcLIJaB+dHoI
Ny2v153zBzWCQRKroy0tFqlFZT3ROpymHeQNTSqfPOYKW5O/mSwU059AwTTyxhSq
VCS2v7E6fMkbLGTLcVOV03Vdl3kMoOCbdXEZaT9dZ9rQGkf17ExET+n7owlguWbJ
Mz09VATyhEKo72le/B45Lq/QewNykEiDUoHfR4bzEyrZupG2k54VqhGHlafRc+Pl
nhO3t2FvYXOM0sxDMHaDZmusxb/bJSuz2xQ9iJKirwXcPufBM4i4Qvy51J3wDRC8
G5HVoGb/YvW2TMR6ou/B2Y/l9un59v7FdDin1IhCfe30/gMca3KJc+/uIJaa932C
uTjefY0IQtscm+t9vqx2s1Wi8bRaXwjGBXsjdfeBl78YBWfhDmswFgwdXfn/8hIx
0fRhjQLmJbrmpXG6BCUqRfWIUwfFG0/Mw4NeAkjXf29mnVyk0rfaezcwgNVAbCFC
WV4pQ5JaTGps+QRX6YU3CIptrP1k2YMNXsWCaosTjMaQ9IUMfQBQFCHeW2+Q71nV
FW0BSPKIPUsZHu0L4FCJ8+YaaZfmg15otHOWinwVuBelHbHvb4j3xGFxgheec1/i
utL6/CZIgJ86vMcPuOnJcTE62eAei4sDfXHSnpmFlMAJ7ksy72WGb8DV1opIJhfU
9l7dNf7nSIxoRn1pIXcup3rydYBPAdut5lkhQYei49NGeH//QjLaBjVMASL4d5lO
er9tVdbFMVYKpiFLnXU4CG1zg2pQs4nXWFa9DugLvZcLpw9rHw7SCltKw+OaRTQh
Ek54RnRhPsLPnmxrYgUAkshilNBIEqYSaA1ZTMXqmIzTLBWtkRAcuBmcyQXp6tZT
jA+hpRxD3/U8pVjwznF9rBiLJ3Yz7OrKWiWys/BBNwybKNPRTdHQdBRqVIeg7+vl
H1upA/IBYjy3rmEGcg0D/YJg0sEfW9x7ELaKZs/62pqZ9VERvm5rfubNv+NwlBuV
Or+yJKSX9HKtBZoNPMzt90uTWNqghtOCxlq/9OUwlDOuyjpF6Lnp0DDBVuixAVls
yI1qW9XWZGkT8e3/XLRcHxvSIg94VwcayJZGXrBmAu68jHUxxJ7CZhVO5avO7sHx
d2vAEck8gcdcsPzHry6XS21U04jiUO1KX4pA4EaSaCExCfBGT1XVywi1u13Wbl67
2AlYaiWZwDMc7ouWUZY7LtR+pFzePYr/s1U/zTJgcoCDQ1ghXoEWNCaTeiELnUpS
KzEHn6SRYkg8Qese0gytJKMKg4JtUimW9zD0jp2EDXbtKosvRV/z6jJfqQf882CW
AS7cDhiDJ7nwuHvxzd+b3Vtk+OoWgu71P+O7SP9nBivtWBQrq9Q9YtzAfgdu9S36
6L7U7H2LlI7uLsYVIAA3BAf+X36JRf2MyYaKEM1TEiVDkw3v5lWLbfdgQ2cBPkPR
HJO0+eqLFvPJn6o+XopsA2MoogwdUCWuOMmfhuCUfSSIuXJF2CLOVUTzYxhCWVgE
L9npQZAqbzSVmg52+CQatFMNE26p9aKUhGu5hdvrMO6P8BBTWWczJwh86Yb145oP
dEX6kzt2t10hv8685S9yxli+FHBsChR23Lw0pq9+1hVthITtbacp6yqPW66rwG3P
TXJJlNLRo+q9uYcRy74F3a5JnVZDMGt1sZVdI9h+265vuQLSq8yhCBQ6H9iTrBmv
FtVq7yzpiaH+XgfE5lGc5nfyyoClNw0xJb5J24oPtwNQ+9UM5iIIvjOxHiomBKEr
WuHM9JVOYQOHHvZlxqbu+o2pmxk0ScZU2pKBOZ+Qh+ifLLnRmrCMwEAA2U4RtNvf
duac20OfcbqP54OojvKpSAeQL9c9y63u0UgarbIAJz1rAoAixvjDIhujJ1aE98bY
AyKKxq95V9Yi3Hz8gqgUZZfleRcSHqJObfWOCzXUwHtg49GaQSlsYkE3y5b9oSbm
fmJqGPOaJxajvQiC+BEUvP5gNhLEg6GK7dImbyItD0KECJcgvjRVtYPFFXcLfjZH
97CX23f9KffBelgtlTsRgZDUW4UG8IIYEp/vMmTVlIn1Vpg1HCRLFmGDXen0RRVg
0llzuQjHN+m4kIuZUm86iITmgEfVCZUSBOgdQ+i1FDxrJ0XwHrgyThlT9q8W/p8+
6E1iYPB5dIPRe2Q7jVkbyPA+P2w+G7wzoJKfI1wnnpX7ZpDR5ZDR23WeHsaVNzzu
AuW5LOBUcv1T0icAni9GJ2tmfslg2LeJcljZdJEh4z3RT1LFZH2DKxAZEg1xU8tw
bi2HrB/BeWVXcSDFdsf3vw8y5KJXH9y2w5IAzYgCwYFVMKgYq9ZcK+TRHrb25XnM
+bHdMHrVvVz6tZUcP4JeUSIRmQC99YuPz4UiM5FG0UhX7WVTa9RsFw++YTY7BDnI
YvqYrxh14FU/pNbbv3Wqw/FXPLiHe55pEP1JixeL2PSdqimDCQNksRPzvjCzFcn4
XQfu1MZiC+SGCLCWM+4eMO/TH/I2O2sUuGLiafO5Jc0DI+SotelJlJXnJ80Akfbn
+m/k5C68WUccpirTgKxGIRdg6ysxn/PEdWUzCOiqMjy7Xhr1VuEBMleZdM/gwZEP
/AFPcexYAmOpo///JUupdIZmGpfuQzkg7Og0ImBq+dmjKoMCYPthH75ugt2ZRCw1
GsGo/B0V06SIfOuhgWieIUGNLse0yoXU4Ua7ieFdy6NKv32L7NX85GbzubKVxXT9
QDIsAD2UqmnKvbSG0l8hVx+BmpcB/IssJl/EHpopgI3dtIHGXvPB4sygF1kD2lLD
bgfNKIPTReJl4LKLxVFHV+DOs+XNBOdfD9jC4POIdtb3ax+RvrfL1M9pbYAIPHHH
MdoSQ1F1bjAwPPY3xQtO4ksBKD/w6NaeLnRmzr3pmD1oJphxRxDjywfWIuQjVyWB
tkdeWqpY5sFpPdJZ6/jz2qDyzwsEP0GYSxPqbD6hPYMJJeo8VDyZ8lGL3gdL4Udn
XsvOTLgRolFTGMAoHIP77KJ8ggV/WgEALPDijREM82FtL54SKkrlIjJs7tQ+GCNV
G37EXUNBshOQm76FAjF1AeHUGN48qojXy1sPpwLfQHJ4DbBqqKrJRatyMaRU75FR
tRfH114TP1odO0aAGp3jGscG3FFQEneTN3ISkSERQhL8gwCwijCwZ1gQEQk/Gr/r
NH4ib1bm/fxRLp+BiK1Z2TApOfNF6paI0adoOjTdBhTocW7V5xos8buV0/ymalMU
jsRXQudACGKcwjeHQNFjHG6lptGMHP/r280RtoZt1wM1Z7kkEhtBQCrbaia8nH4o
9rj5wdMfbQU24FxC0SYz9YJ6gLxZRJcU4L0dscuwhCWR6duPHK2pGWirVgE+hJ19
B2yn40oNsj/F+BDndQ/1L5mxHewtOHn8vTalsJz1xsynWB3UQLWsubk0mwSaaVjK
Ox/sSuWSDi6X08vfHsftg8yADNN8eh+sdw/WXSgH8dBViG1Ge43ISX8WkeGRHzfg
wuk+LsGbQi0POKlHY0U3fTKph9MRCJBM5nOyuwY8d4IUBrFEmvh+75/TbITA0tCm
Ymr8hxEeNUziTLEROblOLow3EcYehWTD91brpmxrh4Abdwc5W9CdnaNf+Q7kAt6p
P62H2XTnZd8nEMZ0P8/RvQ==
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20320 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
lmOQgIOM5jiJrGbWpsW/8hKFM6woPzsG2Er+pN8s9dH/idUYN2l2Nopk0NcXiKvL
nZO4YFl0nLsyJtCjo5D5bjqtKkrGYC3lUC6/NFCSA55Q1qQG1NbXKvd+FTCJjt3m
Kq/QuzBhax0ikzSnXYmPMTfYy0/kyhJDNEZ4/iah0PvPc9mYMFTvTZH9DdiV/qVG
3xBKUtBHjMDCiU5s1kWcgQxLiKX27ZkuWEmeH8lYGYla8LYlEawXWo3q7hGFPZt6
pceJ8oe1H61VpzBoFhivH+UAYyZy15GAz2wC4UXTo58CvcNk44wW1NXoSXn69z6r
XfAIrWvelKpEIhPC2a0qdBN+uOxOZ4ZMHS3oFjf9XAjtj6bu4XAkCrrPJC1zLOfG
YHpyzmrv48oRwM8Spo5tzCwNImlmPDF+b2QK01WtISA2/515KUL+I/LCt5XIa6dM
D0ZnBocH63KHSZvKHieZ5DOZsRg7m15obCSs2xx/Zu7fDKTnvGmoelBJ3no/Zx7i
Q0ILiRAn1zzxUhdTIToVnQ19RzKYOdI9nO/7oG/J53Vlu2F86tDOS0t2QW0cMup9
rlwbKPl03nqlQZfeGLerf3AJDs94TIHWR/5drUfTeX/RtfzL9X9rWQ/Hca2yUN7x
ztMFlFKYBspKhhoj9nOEDOXfWsSMr4h/GzGacF9Tx3b2LaZqUlkqbUDGHUaBgNS7
awSRMRIc28m0LUMPUucklULYwprS0S57UtyPJ3XhQShW9+2eY3wPZFULKQkUi/mD
h1zoIcV/soQan97Tom7RlyGOfWDPWM2A6FdWdDnYek8L+HcyCb/m9spekWVy3t58
itWy0XDOTGqeofqNwJ5nOwMMY7rLN0mKle/rno7PBK5aoCoK+nt1IKab4QHzAO4E
jzecKYuGmxo07SL/+rmBdYdho+h1UoOl/ytAiywIRKHu3HBlAmO2Zq0ZpnuXYrMH
tPBlGSrX/XUeisaxwK0MjZ7SuKUawIuDTaO3aOb1eNZKIIs1xrVkt1TLStOBN4nE
FDsW3FTqSHe8NV89nXXzx2p0A/14sroiHktUKcVaIztjnYWhgeSHFayNWjDaMUfK
yLISRbfYzfExCprsYF7dQZGe0euSKNjr0UodtJOUe76vGRgb6ZjEqutXB662lvHG
IixEPkZIsS6YIY8mpCsvrsS5sGbmrbswLDPk6EehKM8GHGE+NPYy8uv6m0rArwDf
g0P0DzWb+EqQiNZtqNqqjWeIyT6+TjuYGyumH+bwmEXPZaWwbc7Z6USdCkFh25ZM
FFKxpzPudA2Y8zz0RWICzjWZ2kgyxkw0uovlciOJbOTExf5jgid37mQCiWWVm8fh
sGiXvovxFlVztqcXBXRyDgEwNtA+Zv/l3VWnQPT13MkChMlIsAlGYnU7vVKbk6uH
rIe9oFJM5RugtuD7EzDVEY0W7MWW2YT2JovaIVwq+iaxTUy3UDwEQmi6e5M3gRcw
jyOYQCg4t+NDr/nDmV4falFzFxCRchpb9vIIWXb4VtqFdSXMiNSdg3vLAHx+MpEh
86aRGQkLiuVZh3WUOePPUEbZot4HECLQ9vLI4R8GFxBDjyeCjoQ54J4ZBPhOLYMO
JuiAu/TuHp586XFByClvM+ExjEJelQutg2uqFWugri2I00pf8Dyon/sTTiX9EpQl
7yKQ/mlEjjf+BxTa5YhICANmz4LT1l0DN1IWmSSg3V/z+EgEXGun2DEuMzlYwlCE
zV5N2pXtbbTvFMm50fe4BmRsGSjDwzInuKN3tA0JvH0EDA4W/VbhbMxwzpqUN9dN
RkDSGc079Uq8k8UINA2fcoPc1MBa8n16rnn4NAwgfZ/fjxieCf6Ua8OX9IIKsSu7
P0QM1ppRmn9J44us9W4UG4GAQjVvQ8uiCqhOvR2Am9/1AJXiwcNKrd0p/D8PUjdc
cCc5ESr6yaEh2O05EOnLWilEnst9nkU3keAtoU+Fb7oiQ8kOlDj0cJGPgDHTZNNS
/kD5mVRvGhV7qce076ETNdVz2NQTipjvrQ4HyuFWfRzg7ZKFkVexBhQyHUXEaEK6
xhKIZ3E/O4fpOyVYU9CUYe29lqh6aazBD7AeT/F3vUeyrMqoSpQYl+WHfHep3zLr
Uvymw0+QjpgU8ksbq+9G/sZiT1Q+3RdfNgYSxRG0QkBny/tkV8MdNeIuS3cyDHBv
XqyAz6ymdYYOsZ0vfqAkkoY5qHVDM/pFqVMgzj4kqqmQ+TlCJMTEBnBbKZFHrmrx
3HD4r8ZO/3vVs3Ar6X1irRkdPQ/8jTUD+bsZYzMFda+sJI0SrwN9HPa2qzr6FHgK
pTYTBf1T4lLpimM4fooQWGrL7dKluR/fiVRaSZHr6A4KcLIvaJyA36avdn2pCXaW
xhjwDQDA2j40JrJG49nQXZZYPHzwJolR3KDGYWmP1aiK1N4zRpu08/3tJ8IUb+Gf
74/5CMV0j8u1e1zuyQ0VNz7b8pkNsHT7FcEuddi3vCV14P1WuE5s8D4fOZI4rSuB
LyhJjdEWITosDDsohrtYiZIvtJaGPwEO1BUyVcLbRe1Fh8nT4L+GhGL/pG86ko1w
X7duVLJukkYVl9QAdIi5XZKgu7wODgHvWmksszlW15ukdBZ1OVHu+9EIZ7ETNEWR
Mm83lAFqED9Hve/+wwrGGJNR2ENDZAIzGpeQBECE2HRf4GE5AQWtgOAarqaOgnMq
I4sFRDcmzHRIy+tg/wzyuNWpsDEvEJCmOrN/gqLF4S18egBB/Xu4nxuweSwV/kC7
Ra57mguPx3pNt/MrrqcrH0+7UQLK40zBLWpG1lEn5LXsz1nhMmv87HHEOJWJstFd
ICSnJrrxWxr6Tom2FgxbmWJQ+1uNOOgzRQ1G1qtENFw3bt1Tp/k0+BVapLA9iqj4
WcOjPrcCvU+xfh4LEtwt4L8BgD5GiXDceC9CjxMYyBH3v2p+vCugTQS+RfN6pmlJ
nTTf497osJFMPhz354f/4sQ9jXWoTbKDHBSLltIxsu2CETPkad73uH34u+BrLOY1
8JIdhqr+j8GnfO+ijmwO5rfRLSMKOWkW5EfZc3/hPETSq7qH69Aj/14iq/Cetn2Y
vX22eyIy03F12gyXmKkkDVSyl3VCJW+T1M9+J6kScqd1HObilrpUFYwp7Zj+ac0h
RxF6kYru8YW28d1WvpKtSdR5TFLYn7hWAWnaUmfzjVVU3+fAhnvhGUE6gGS49rCA
AIS2iuNrkRgJJvycaIfnntqlNEuK13kdLKzots2tqD3kQVFld79E3yph5nQijkHT
Zj2mr8JZD0/i2kW34nv1RDKO3FEs+HmqWbiFeLHpILLD+TOPqEBjWo91vW/GX46Q
8SP3HBph+78sOlFypVAc1DYKmOenJLnX7HXAnHdsSmk2rFKpSLh8L11X1m1mMZzb
TbBBNuOiVhmAuPw95b6XyTWCPMXBt+jwWq3OPJYZ7rA4Ofks/zjeD5gLmsd34xTK
ivtkbeGdIB9vqREf/Xgxd5jXD7vBhm3nE9geyrmtIZzJzB62I3bgzwdqgbx74hu1
vZ/hjHqQj0W/BhkWzVjR/5HGEvBb4RgTak+0WJWxkIMcJwAIYPOPiDUr7JkKoMWb
X61ikJItpd7Po6UwLJ8lW5z6HjiMFAOOze4Klhr0q5JWAnIP9+/vcyXXDGAJK3mP
Q53T+41qfonl8jYybPUDQHKqC5vez93Ov6bWF9o3pXh5y0xVdwO6LIcfzXH0JXTQ
EARxsuut01ikVR1CAPfwyKXHmX0TaspqYuhnaDQSfkIQSXGDGQLsk8KkMm9BFW5Q
Eqb4fOoQEzqPAM1rz9QWQ0rnMerx6FnqbcATumK7Sw6DZrAnuGG/lpEGk0D7e2bK
rxTyHxCzqs99p9GODNqTI1lqgDoLqIVeCV+AllMymYSH1dLMEcHPC/sKEYGgnHGa
PV17h5gaLSYCEW3Egdioqhb5AjQmahr2ZGaPaNk26Sf+mk3fVJ3uQKDZfe1QMkr6
KjeQujM2cWuNl5JRvXQJwnswu37Q6PAjMYhm006L77eu4vQUgkei5z79mb9lf5om
r0b1UXZ2HsylRnvaZUv2QawnBpIOcw7emkSxDjbWZrfi8Hg8vFq1lXmkn96q4ZB1
rl/NDzBTHX1P6+jm0BrlBthVEgOPtlBIJOHFzioO5Y6C64c/tzcmxWx07Nayh99Y
7r21OL0iC2nQqzg0PzQubkEW4Y9XW3gDA4YJHlZ085pA/PEUifuXh7Q0+4ogmEl2
6ICPC/FkNZCVKFiJumW2btXst9OhMa2jItMxaTZt3VyoK9Q8oFb641E+fz/nsuf7
kOk8F1iWFs/b5xUMbx0OKCiMPJhOHaqnVOtZ4gi3nq4btK97pClSWWTCBzDXjwwb
c2f6SacAV1ypJTmVErdowcNmSYQkPYy9df1oWoF2TcacJWh/gr1OoaTh+PbNGsBy
ZfoPvUR4+qQ9ThJ62CXB9PB3tnUQongjJzYV4/0wtrCRX5w1mAGmjHWFm8vp39RA
B/+dm5CebiEi8mLFDjFTNfQzjr40TV8SwOlRtGOvvuRMfOjRdPbQeI5txEy37pD2
Od1BWn0V2PE0S+FkBOOYOHjgKNqMF1utZ6Vi6N4KzYfiJIKupkkX4P4U1KegWBFk
QRnmn4OXi7kBb8wIxYyvkwICllYQSW9/xnYLAe+yrrv1mrKfi5WFKmhzPEozVkfW
2OLZAI0enQCUXJPducLrQOqHaUDEePhXZI4YrYr5ynGeHASiOGaJHL78YtoLRBGm
VAy13CCZz3ALszlFSz+Tzkj49oG/Sv1tUAb0jVASj4h0GKJ8c1z71lxSbKMpK6mC
jJtWUz9KTv6eNxtM/zAJcJ+lZAWK08bZZfR6/9Kyilq2x1M1gUGElqOi4YZ608/v
PelchoG31bUGNjv1dKtVoWLnx0MlC35OOCUgPh7i6OUlMSe8KQLM82IRq0LXWvW7
PjM8Ko1IGC3cvy4oob5ytRZfkMq6Said7us16/9JJgC7OD+a7Qe09lFXQqiyLr+X
FMo836uLrxRmZdlf9OM9vp4uMgxn2I0dO5lOGqUtCd6UmJR5ddg5QA90mRLobZv1
QULDAD6rJKZkVhu7De7neMdHu2teH4wjLNCVRs68Bs/wIUYPThGJISgMr12yYjzw
YtOefng1NvFO/w+qINNKIKHd/KfrUGwuWNPsWloM7+JAKxkEL8vfZRxOLdZlNa5y
x+MwZg+4MHsyRZ5iJPYq0kZCkGr+ARLkTYRLp8jVg68x2CoOmwyjVFMq+vLLTQGB
AoIjlHt/kEKciSoQJRb29cSw+TFD00X89h39zzv6ul29X+Va2F7Bu/+p2Joxolzr
+WO3ut+tPl10XLbmMJhcpxdTq5kRm/bRUYXgIMWCZKN5FUMOEQIU9XHT3Ind5QSL
XKQ5hZD5GoYEnvv4uNIlvRhiNQ1/1tX+7Udw6q1FsvpVAhkXAoBOGQpTX2VHUV8y
o6m+wyuBSdiT722pvOQojYidQN2H4xt9XNkRvqyes1KZ5JunWcNw1zY4FYmhV+gu
poPDUA+FYZ54+QhEZdEJCaFPmiJlBOZsAs2BvEOMy1PsQRvNk4Lrv3O4tyFvtq6q
FU30/2SuaV+YJ/58Jk0em8cJhpp/LGpmhpHyCaWjxQb9xXdfnqKokFutedBvdYy2
EDkVJr4kPmXOYXw7OL7DWiWgcZuv++hZaYYt7O+bfVWZgz7N3oBDzRb0DMH1QhiK
GBxj0tNdeTZn1tzbDmwDlpUcfTT38yNN731AEfpUvGyuJFaKUeoK3iCIk4fEfdbT
64Zb/r/v5vyPBC3lVfHsSM0j2/hCKKz7OKY31pCwLMh0sEFIb5CucOgmWhITxG/d
LtMy/VU0eVulYQWZcNunjW1WXnWJgY9zkHezhvZRKy1oyy9RQoDygRJuYyVO/lTI
bIItaHQMuLBPsHcHno6sjEtpoJfnPCoYrngw7aedLy+P9X6HLgYzLjgHYAZKIrbo
fvPDMDhAD2LoZpWFEAS8+92H3bcEhfkqcTrUGrUXcWyzOzco9C5gHw0bCThAZ95e
hkTcv+9zu5oT9XuWTXp+/9CFQm9f8pE+5BQ3GC60WVv5+YLGq1IJry82fKbRSDv1
xrQASaLbKdWLRGJPPsxvEy5ZVEikfSSxLFYG3OtpYNq6NLzhPvc2HJze6OKp9NZ6
8Q08cgsf2smr9awgtcJ05QY/G5t1rdzobladQ5ZNU2+x6EkW0xuTbjKJi0QIofSg
LvDlHM2PHn/IHVc4Ir+DMZiYXKig7slpwEEjOuM0VktDhE+LSyn/xojC0SC2PKK+
fR5twWogQ6xfDNOm+bX26PMvdrG0uXEk3dUvbbxSShapizR4qgKJhi4KUps0/qat
CQ0XnNrTPD2CBNrJHYdfI4i8i82FjEURcPx5puBhfJdTyZyjj1bb13E/YGQGCGot
sGRQ12jV5RGycxNxp3lF4LfS6KfYMDIbo/yKk4MHC00bCHrTO1hUPXwB0eCE2bsF
DZOHWcVnxnercugny4InSg4kqlwGPKK8dDiy0HqS39EQAAmXr8UCTb5H2D5NW8NN
HS0juYE/53hUJQ1hdtqlihKaWpvS39GHykEkflgyTQlpn3M+Q71wRgtTDSma91cK
jkfz7ZnrODVr/G/sE1lzJ22U/WpOezg1CjgCkLB607dm2cyofTD7x9mVA9+IOXMd
yn9plvLR2r8euGVuWgtk5NZ1YrL0xLE1sr1f7CMBl3ERW3vj87i0Xkz2A+raSgCY
/Haze+NFO4oHf6ya06HKPNfxuR6SyoFxbSkaS5FtguScnj5JKD5q/wccrbup2hCh
SUGRiax4y8OOiy6FctADmaZKyKnulPA2TRMhuV/A+tuM612uK65Y5gGny2P4Q4uy
FHNZJNWlSZOSFGGRrX0eGnewPNsunxDoFRa5eHI9bLYp8mhf+rWccr/0Xyx0Kb4J
TrKKWyAHruD/KiCiItNDO74DaxFcc9tlRFWjeE4SjjqeVbwA76160MZ2Ot/cQKVk
TMRv7SmRccJ1NXGMBKoqu+EmizFFtBirb6ZhOh6Bj10/s9OxqkhMBTll76U5iMbD
/Nsv5VIYzOL5gbwRQh9gA10119uJJxmQ7vq5il4tZVXDvwEXNynyrdJfEaL+G5Yj
jMPlQn1HN3l3kM5Ub7QMMZyPpI44jDRzY2BzP6PrrCMGpnj63NCxvzlSJZVFu57i
vzwOdYlY09fC0dxv6xWITwiH0fCGWpK8n54MkNgb4t+cFz5wI4djUvRlvfBNcBzx
PIA1tGId+yru924+JImcv3OR64CZjcIfFdW/S3vBk3+VsesqfcG/T6MZqphEh48s
6AG1s88XPlLZC+G6XhUitVhrihZw6jbpG7Fu/xRgmm4hw/IMmdJIZVzTKuHG647I
q6sF5VUhowJDMGDaGslTl67OiHX6oNqRHuKmrJS+urxXHazYIrf8blAjwQ8r4iKK
RfHdKt/loasZHimS11FZM7zooKTvH/S2OSFckftg/BHy+lRpsPyQhy/JuYL09czd
0SwiI7YPsRTUgU73UxXj21emntZgfcBIQ+98YlaJChEcra1wW/2+7dYq7Y+elwM3
gQcwOcHtox3tQa0Nrlin0LD77JeZGKQRj7rkM6u1uClgxxpYwkoRr8Zdr4S1j3EM
z+lWt1NV747uWicnZsDhzOQvwIVIM7uvNvmtqs7c5rToT7OULRJpve43jD+sOvXN
kIiGfDUGOXmkcXtpqLZsvhpO5gt5IA781mxY5Y+yiYvbfYWyYY0LEvgSWIxBw9YI
Z1LwYzxPIWbdB3e/1HMjwI3CafyKk25SUWxX+wUs6vwDkAlmKqgoCuFWESke9qY3
zAIwS0zUuj+Bt1tFTmUx5GcE1EvJyiCRtLbtfkHnLQhba9GIw0Fvd48bNBJQhybY
K4exHJPKLs1sUPtTY4b7+j9uewcWMUf3zvaXctRbtFJFvONhHfdjst5mHwFS6BdC
wVFvwpEnR8U63wLExbUbRHp42fn9fYWB2tbffKy4qAslSAY2fUXlRD9Vp9JcF63b
IGCt16ib4Sd2BcG03SrK6FQrRvQ0oVc+5DXbKnSxsMerP/Orp8v1hGQ0M/aaQIex
A9MNtfhJQ2b7pT9Ibe2hLpbYAy40ZWSgoMOv0Kw0a65PivjBdB0WofdmMvMwGoJe
ioRH0b/vBKL/YNob7LhULaOalQhqfMngGnfzeItr1rNM7DnDHG9Drbhkg2gezC9C
CelhmUiapqilx+59v7gNbMQQYCkdxQ/ghX9qlmmg4uUfmOZ1KaR/bUh2qAsR1nne
TY4TlMQ1i/4bSsE8lFqOLCxzMbmiweF0XXtmzM+vsw/k8iIKOE42Hp/9FtP2bAG8
0mUaUQ4utIn0f/LzQtp8s6h8ZLwrSMQ2frBNr8cYOTWzLS1aR1g+H4V2+JAstOwW
joIJ35yPKIALBEtR9vMX2dOB4EXByLJRoKbsrO7grBKtV/m+YDcdCGHBYr3d1wMH
pgKOUGNbHLrHsCJPuyuFbgWCGSFAQxTaK4gWTwRfwG7FHULxWXAFLb6IGU4moyzV
DyugvuvJQPmlO0mJQP/50aNS8FOgjVx4n/0wa1v/l5HkI9SyT7gHqw7o+MgINF39
2m3VdFOhrnsvpY4Bab29fo1Y4IBW7pSITsP7VPKAHUSh2W8cIhHV62tRfuYZY+b7
Rwd/eI2sEX5lOlbf8KsAYlinwTO6v3wHF8HMP7IUBF34xb7AVJm3txy6Q9cF+IDu
sV7SotBG9+pzrBLs+Ozmh73bsE4GK2E9sjdZQCPsxpnHX321OvHSF976ZYHJY6UX
JGJS1UZgyUjWp9SvCGxyndkeEHWfi9w7aIHPie94hmLgJiBQ6/d4omYEbJzZD93n
WpnsiSxm3SplBdXDJH3V0DNvvrohKTRQ2vEMDxPPn6dG6nj7W+fylcFifgyWaK38
nHpGQg4OJFWoTPIaPwogt9i6nBNLsui96aElgnC4B9GWwxJBBx2HH9Cv7WQ1TaEy
SXtlF7ZVyTHIeQemHQk8IBDZF5FAwKq/tASs7PXsVpItzACqylu3d4TY2IIepykv
8nBs6UpBrnQN2MLWcjm3ca2XNPTtojrpTZZXulM2X0KF0IusE3UXYQX4dFjwkqJQ
IY5EQzQciXaLJ1uNt6+ixObJojSP9CLRUImIM/TrbevmgtqZzmzCfuKQc/XeJaCX
+cgSD6OhI2pHeyFS03QKEy7WzA1MZhxu2PMgXGqBep0IJ8TfQocSZAq4youzDIY0
MC0auQhS43r5dr/EWUJ+H/FL448WNhMj+D7MjTAjqCT9os1OSkoZC+EBnT+HLlNL
z4w4FPr23Ly77KAKDJqIAbpsz5/GsnWkDKwwvf1nlMvDFLH9R2g93kZMrcMNYo7S
ulrp4IYc8K4Jazoa2ddF7qP2LMHW64yTxWI/LCUMvStA+dDS18Ni9trpQJ3cRPRa
3Gga5mWn2rKE5k8KcYFjb9vw81LTsRjeMyaCCIDmQp5xBJb8CuAHvRHufqNLJjLh
e8iY5Z92UgZrvfeOTJOfULbaHQgxU1wrYjvCHRjsuK8mrcoJ8S9MoolqzzWHX7MN
PXCllVMb4WVziDtvtvI9qynY1QcypFep4pa1GGr3THrHALpwGXm9SIDl7I1hyvx1
RZ69KuNjTM4NLeSGg+pl/7nYYdQuaxI997XaRB9UZe757S2tZy4JhpDMmhBeWG11
xA8jkjPDOkc/fDgr2sX7V9SHYQiYDyxyX5irtCXCYm/TRwjhFIvG7JDigU/28OR+
F+WcIva2uRwlW+FxuKrtriwD1bfCS7pqUm5x5nOnPcAlPAcR3Q7euB05PmSz094S
cUoDc/ach46R7/X4VAEI2gq5GDbE/d7DqREsj6Vf/JVVucFOTnY8374w5kao1RFC
YTlyQEtZGD90F7dLxu7GJe5T5S/W1TcXbc26ClyR4KRpB4lAkv8JQQBvSeVT7zW1
YZHzoQgmvfDMc8APXn5xYu3weYPumncQ1Krb2Y6sSPGNykVOtoMqABB9O845M6RU
NfCT04G8/8KMzRzq0NxbnFmxtzXKuaDpg1+gutt6kKP+rSOSh9TvcgUEYILo3mBq
rrM48DBB2zgly7sWgWF+UAJ1a+VHoOv8r2dsPlmhh4j2SH5MDWIx/3o0GhEBs+zP
zFo47x7f7vFrwDi9BMQkXSFKRB9bON2vboDbXiBAeQZx7eQ5hlw/sBhcMxZyBWmY
HaEo7SxyxfjfFThgX/CX1he4vPFOUlzK8TJbf6buOfg+HwzEfD150rId6oOi0zEA
io7HxAkv7nzyf/fWM6tFZqZuWJi3jfCnJ8DA5Bh5TArpri4WPe0yhXP7Td65R8hn
dlUEMNObhRcUlwU5p7ZJe4CMCt66sG9udZYjw5neIYMn5QG1C/WOOPK0l5uP0u8P
wCNAg4NeMb8UNh/bsolKrLnL1CQKq1Toig6/UI0JtEpVJZh7l+9Dc7H5xitI/hIe
TkopiSBEq9ux8ao+49dJdEQvLw7Q9R5ZuS5sR/CGWxyaWmXadGYk2Mt3Qt71ph27
/qrUhCHVukJ1ZsiOU8q1+b+mqZl7lqOUHgMlwPy4izeVCOhMN6BNhBQNGPUgW9ON
R5EyO5l6TNh+CQz3XCCKJt6W7k2pbzAvN2z3fNTiWzFLJZSbi4GKyS1UsT6F3tEp
L4tuQk31KJHy/zl3QyTUOV6OesmnzelMEMhSb4Tb+iE7ZOdZd61Uw0gyDqaKbqiI
y6dApwCT0tfHyGhJnNfAp3c9ivGBD3HWhcqIVMxh+hRQs0lfubn8X7WwRgoXh7tV
A4zRcrx6FD6w4ohLNlF/QAhroBL3O7XVUDVsTjSqe76kOe3oQg8LFGW6Ej5Gltqp
sTtoKwxLpp1lASnVceyMqzABClLZtI4x8rlR3IR64FhUt1jfrHYV5nhhZdWEnjLF
Q++AgqoITo13WNPndeKPywklhyHlaA/QgGYiQ/OU5yBXVIKM0rGIpwiM88/1CMza
cAoCDF8k+vLr3x1YL94jPAXAUW39PG5EmPUtmoCXx+v7LIWnK1aLOliCdFf2OPAR
P/7/nD/tF4wlA2zvz8u+xUxhLlO0fIcFzgnA1IHfXNVg1bRM6+Ad58wPc/Vbv+Jy
TxhgRKJyh03yRcj6dty1Na/IT20ZL5CmnW9ZVNPV600lcPSLsJpzX+7ppNB0xAtN
KvX04jPa8BttU/hnAvvXvgzgUsQHtzLCzXA+ApzMJpKjaj2ThD0w52scqe+D9OqD
bmU1NzwjBN0bX1cDpwkQJEpFE+NpSPirF7FZCnyhEWgWo1J695W3kIUkNl0O9b6b
tSJhW47hW4bKc61cfvbp2gflON769aT5TX1f/5ODXWnsMADN+ibYbV6TylzXwVr3
j9efmJNOtu/Lw0lq3HRG0qO2oFyZdB7q+QgDMk9waqS4dtOUAYEoELTRSsMOgkMp
RoUCFCDKJ6hCukM8STYS9zO1siFA0XT7dXElPNWKbjpCgdSnr702L8tFkQXHfbEn
rBmDS3h9ZjKdRkXfEJ+AVotz2VUdUzQOL8VN+wWF6pKDjvetmF5XpoojDvSRbd2Y
9xjWXEhhiAWq0ycykoqo1abl6ixcTbR5L2xSoGtspVNAQBmAgDnWVWKVGu7PoN9k
9eeCvlH3bpnddkTmdIifw+66XNQ3dZksVeyGrUAfE07ZPkfAYFl3AVmfwA3P5YIX
i0pq90vh7KzJr9d6sw2zVrwKZpQQ08jN2GFsF0ZysIAaJez4XvY7fQk6/NT4Tktt
s88XiE5Pd+kckmGLL5vdyjf3WW7rJcbXPZfjn3U/EQ5YA7ybjlrxCMRtldhhn97Q
SUz8LMtweNnHkuRq94akeJQdAQYDD246Gl4c1ChT0qIbrjHAst2DIvdeiYjD8OSt
JfX1ubhcaKt8ss1Hg7aMEdWLFbW7EnN915OMORv4HCJvdPhaQoEaU3HKgHHrwbzn
kg4RErQMxZCIOKCrMxo/EkA5DAEIFpKs55Z/xyJX9CNHhiPecV5Xmicagx0lpK/O
vKAor+BgUUaKbmpueZ09mIJzD7sIssDO+oLyXS7Y1oWp/0cDC//RitgYH0vQzXvo
TUJuiGqsX880Meori9PNu6n46MB3mcHF73cvdPjeYsZ68xxBdCLTiGZkCXAMZoWC
L/zUVrt2ENmsdWNXnoxn+e9Go/hoIw1nIwOhKWyEQ5WUHphcCO7Pry4icu9DNxfB
9/UucFYcHv2+J7LlcDrT3D+UzOB5e6WLOgp/9VTfToAfsI7cfSk7KnN0YV1/tCGN
vIuvO8K9qCRc80ncgvPr6Uy0TKjn5BlWTHepUYqS22lMAWaR7wJ4fpdAq4cGFf/J
IkzYiHzUKd0q+zCxDLlrYIv8nA4BZ5h9oF0i3umVl+V/wn2a3MlJenHgHgJHKYkD
vWbn0tZgUeA1zklqWl9n8IWEiDZMnMakBG0Lo4LAKBxtYfV5kFX7Opvjh2G8cHhi
4vzefnM7agLegeMfqvmxW3EgcAVZioMsmkwh2322Tqp/1cFpK9idhy6hdpeso5NP
lcClAXxe1p0O1m/JS0fEBbv/VxrYfAuV0PI+gKDTFSUz1H+FCXLLGu3QJS+SKbMs
mxtmO8JJoQAq22+RPVSM01US8MIJmm9eQz37wnCWqOl0lR2FwePB5HYYZEHKFzLd
4voFlcnXQSkaVrzZhnj7QvIe4cbF1QI4jw3pBj0ZJzWzFeETJGKwN8fZrC2RDZgb
crBS7OIc1yBoPtbBUKCN4u8K/x/mOzaosCDuJXUQNLKufEs0PlTYYjjVVGmrEtp7
/qezlw2xVE83/u0JZkD0vQpfyNutvpX0hZZ47flRABjMsWehx0WN9cR8aTCAOfaG
/jW/fAXKM1qxHgKBnMm0D9hhtazd5jLyP2xj8M+9k/t4cWfoItmcit8pf7Wguh5K
9GQZXeu0pvrmlG83mty8YnHohZ3crwjVD5kjt7fjKdvfJHrW8XIM5HfmDKLEHBp1
b3QpjemPCXqjZQXkHTPAwC3YNRgQsJzYuecyZktA/NolLvwi0d6bfpqPD22lGhps
xQ4G34vRCFQMM0r4dWUwSQCKfl1+qE3Y8vz4lx5r2e//gktchGPUht4/ZmPuEj/Y
4hoCU/TMsmP6mBUp0YlYBFxfrvifVaXiSL7UUMdH+dOldB1ttYkb7e11o6YuyM+L
8G2KgKcUtlsiT/UaTAzOqnpdIGnB2k0lCgTAdM89vy7WhYbwNsOsnWacVk2hNlDp
2qUNMDi8uhdSoEevkR5+eJfpckIghmjEXpMnnsPgzx+xbMQv/sXTkR5Fz44kCIGd
E8B+iS4hozaL6/5U7NGGf7GbwEFNDqIdUx7MyEyZYLsd5CLp1Z6L6qoWy1wYOR3x
DkuP1E2/+h1kuwmEx8ERD9nY1OnKmphPVHWAPjbJMupY21nqIr6LpyZQVVNd5clJ
VM45TEkQNlvZggIYFueQHU/M2xKtDSntW/sojMeb5lgcX+znBRMdDJFOqi+UulB5
J1bBrdSQOdYRBjR4QuqSY6PdwUvKX3p7LjFQSyRPHoKvyXy6is8HUs/aGPBKhuVj
AlN033hNrod3UKO6w60qGREqUPSkzFfhxWcJxGv3Si+dpb2OeryeT/ktb6xhmqOJ
3encKkN1sNdkzfbb5SCFYbX7c/ZmcLoNai7J6DH4J7Wq9A5NkZsVU56mvhk8KIt6
NBxOzXeZuVhe+Tac8wqs6xNi3VfRfVLOEQP8nfrLRBguM7FCVsxCjtJn6Vokc/jy
sQ+jHRpfy4z1MAINx4k7s+hfXkhRDZ8CCGKg0NcvGpl38fF08wEUs8GTRpwPY/Qy
EClkd3p/FSa9f2HjUh3pzcE/droMCxeclccgXWagz6JEcJWJ+plmgqe4T9PdxTRu
tiV4iFp43YGDbM24Jm2i7ifv3x2qjSsQnbikD4QNFeQagMBvNJgk0bVLdnk7gx0x
tS6yWBr0zIzu+GKzN+P2Ck0D1EguDZcDfQiRoGtdEj2lp/OKBfoJKKnHT8T4p4EO
WoWc/1bG20vdPWUpdqg5eq8VkmLO4Cgf7SX2WYVRssZyb2CZdrZfK/H1RA+xC0dX
CYev7/JS9CKrp+nwxF5bNcse53gWq1bw8jjbrFjgADzoZo66PDAn5ynPX74d3Pz2
KIVeGV/4zCUrFhlgOAYtFsLQmY+3s7BC3WmLPMYlzvpj4OH32L1neCjQnFR4/E0f
f+SeHNWH75JBvec0KNjdXXK+vl4cZiUAHvsxgPDK2DWbWL02m6jvCDf9cCgWSr/V
0PJpkTwExc7mqlGE0jAM+m/k68NNBe2tQjd7IznkY5A401+2sr434TcQ3a7yBGhW
d9lYaZ+sUsXnm/W5zICU12EcFIPV5MIGLxZuZCSviqS4zUrmIX+btSxmhTtY0Zzu
qbKzkn0X4082uEJ25kiOHJ2LobjNcprEqZ3ZGj9a4PQfWRWL7DoEr+ivxHkleT9T
1LPOtPTqzP1JQpU5IMXUqryoC2/u/gcIdPrYfKcJezwVXGHSWaQ3zeASFIAA+Vz2
O/UygFyCIrwfNhOxYPBAVLsHcdMHyvkEAi0HtB1bxYeeOYN+EW6qcTjqXE/kdtVU
kf8bYgt4dqTqBRPp4cTId4RlwyMcbE2NvnDMmUzJzY0eFBMA24UN3WgsVEMrwvaP
Ko2sCFU37l16ezjhJgUG8/KsDvEPQbMfxz+AFuCVuYVfWBXKGFsFdKcHVaodrSDb
e1JbYhQTN2LxCdi3rU4MbrNBYW6mO02U7QMb8Byd7akWtcKuSRo3BeVp9amKLU6U
4E/J9ycK4RpFXTFnm5pBN5Xp0IJy2um3QDF8nTDdxgawBNEUim+m9+ndUSXWpJcS
Y/m1TE+oSwJysOen5pmVu8fk3nRBppNwaJ8+Li31HUljuCEkReOhsfihhBrl/8LP
75z/4OaMCkxJjO+uJxtLZac7TUSinPWc0bUw/y1bM9atVaWufgBHZbbsu4CTtrmL
jx5Ml3cUs9Xkmh3CjUPWO1jh4nv0dT6sc75rx0zJP+Ea/aiov/CaGDYQCHxHfOGk
jr873nuuhjEMT1Dpmn9WtqP0ykt20SU/uFeG1rt3D9qk/F9jDG54R9Apk1vMLnF2
46HoEUqTFLar/KW64cYPBpNMvvfm9kcGtiJ+GGYIoWEg0rGfSUirORvgtgBys8c6
NQIfEcnN2aGNNC/scsq7iHXl1yglS8ohM9IF++LjnXAREiUKuwFX19wZG+PJJ+3m
HqRqoTHWgqaWssWI13S972DInxTHFVcVPmISeDWYlYNS1l1JsKPAbDhmh00VOq1l
QeHKVrclDyzrcv0MfZoFoXN4Cu2A7OeJjYOvG3mGcvGWWJDfWEkwaj5ZOhi8Lup6
iI+HmQQbm36zcEntxpurc+xR17LvIQgnI3DqSZ8b+amz2QXao/SpeYInjvDvG+Nv
OjqU5Y1YIgYymsKQ1YADr9Qf3kBJC8UU3wwq3WP4M5cweVywW15SJSH7HwvfARqD
U8PJhbj+/zs941lLdP2118cHC+mouRut2m0wQn4ee4aD9rfx8Omjas7ojvagMPI/
/Ru1mb/i/wT66reUFaOqSelgoJuzU0zrjtK+cL69DpFaMxTPvfFL/TmNi3xAEaaG
muNlfUmdyvVfFUGWBWEZKWUw3IQOfR4Odj4mjVwnNcco6I2wVxeJeup6lVbG9WGU
EmSJR7YKx0TRfIpFDztpC4IkJ9W81pXj7/msQAtCoALTs+2imKIoeNmThmL4e+oM
dY31ajIZjRGmfCsGzRwX74q/Wu+WHnffDZiwZB81YHr++yJIADTJdADHex+y9GF9
H0b58xar0nE4n4V+bv6b7usMrcK7oWpr7ybamMLRRLUChqsplWiN6VHkEH6DZ7TU
i5JluBHZbIIAGUa9nY7IbTsMUtbqLNWp5Rt+L4ODemFRHjYQewZmd19JfAfXocos
0a4XwWih5HtQ4nNbzEhubdBMQCN1Afply3XODrwx9rYxGCn/vFD0UZN9ICN7g1IO
l1lYl55K7nOUdxWRILb7TkFsnvj7QaP94n6qs/sPaExKS68Z574nf9lsfG72iQpF
cUPRGHC1qPPjmwVkvHhHABj1si1UpFueM9pMgAx9vhm7BIsvdDsU5UYJ0VYcCRT3
Xi+U2RunYzPhNxppIq+OCiuPH7r89/f7/WxoRxhGOQoZnbNNMftp6Iv5ubtoIDOK
ZtsHkTr/QfaS0dZKNtmNjM32luhgmKatAsVtjtmvaN1kprtJmouRzEGPRA/cocjD
A/w+JTYQh5WXRzz9HJawYAnDOOLZfylmiY3w21/LXCCkjxN3qcxptkja9+p+hGHC
JcxNy/q6sONK6xI77mXZj5Fw3juPh41/TcSbJ5wfvhKUDWrxo3gAj7x7BDp/5RUV
ZLA/d9YMmZBnOQ2l0CX106eZcJGr9HnwVTPAOET3tLLJlKMgqokvIpZUYqkXQY1F
pfakk2bNwvbk+OP2sxLxaDxWQ08qFIjP5c6GtYBt+Z7r52T+NeGD0jSTs+ybYqg0
bU1DRdbBt1uWwW4pYicAZ+d3LdudLn2nVyJmFGEXV8LtoVUuAys38WIlf+LocVA5
jrQmKUxLlQ0ViJERZIOT5B+/Wp6BGNeQoxvnW1UDQ4JuA2IlsPAwr9Fc6D6zIRMk
2KPpUFgEjjBrK+4UPzTcR6Oo77IUDFODRV6N/BF5nojxKASZ4ZbYAesWywEch0KJ
GR3owq+FlDb0pE4aCpZnO/UojzmqCs7isGvknmf+lh1KhRXFRANw5Z5BoSncuwlf
TXY3YibwYHKKqIHSiPXSt9JKJJ7S1PPUAz8hUJKLpPmRIvhacRHLdD4rsnJwerfZ
OQWY0KBQg+hjp/lhbZLLOxObrfIngBIYxkWKqRq1XlNLazk3c/V2MizepYTG0jYl
5HfgJGd3yFpUqx9WDuCz3DUKha4SoUqzoJJX3p4nSIl8ovCKlwReEfeAfHA0H17k
tYwQGExhllRPOo3AWQVN/IQkSY17eekFslEn+YNtO5+v+GUB73opPMDxZyOw8GtX
QogZ5PXX6smbLuo7vL6d/trKaUWd1a+EQmOIWUG/0093Fd6qAr0TjT6Qt8VzsWdc
kYclAsUXmWMhsVzdZhu2sasSfP0NqWM1S29A16i7HS6Q/2o9Y6hvALIMZcf0Ua8G
lGs7NwFCKWQac5KyXiZ9PbdiJdVRMChDTz4VtCFrg/s9bnk3QdvAiFtOhF7szMf2
Y62xxnNSHI/rP2hfSqmoOr2HDad4uf2OSLc/KjGmah1SVnqRBm7b0sW7JNDo3+wm
dUAHmpNhn8ZPvtARd4J2ZvBKRlln+lwjfU4oc1N/ni+0TbaCCJl4uP11C6QcuTEw
m26Om5bK9X9UdtGD9MguGaWo1pLn9TeGL6fzP1+nUhTp14kKBEuIQhrfLVjE5pYo
euY+0Q4Yo6BdFGDolfhIT60RLQxqvo3/mE/bBFQn6/jhk4hdgDseOVlONoHgMfVp
UBgZf1pdblgfI1VVu/WVl5BMcj8xA9+H678uSv56v6DHFyphGsaZiadEgsf/8YFU
D3XF38u5uNvTFu1Gi5LRRY5vOn/hrplU0lJePp2X4wp5kueG2rBbeK19eZ7hOU3u
AWXooszHsBNSzhn3I0yf5FjHLJNi6cZnbPtXsEIak0PebYDJjvO0HYY+OKFvo4AR
tuOoOUOI2dCypk0RKQOzNYRLwk71GYltteqcv0WJra1Z5CYrirPT82UPFJoGkU5b
qqNmpr3UUbYvSnasEyHHMcHvqMDG/d8p5/0VyCYodfGUFBxlWhgNuLpHYv3NQIOr
DcvEVFX3GdcAschZTZz8AZkOUvaY+NJ6MTF2Q7EoxrpT2Q5b/gGsubFvrclGi+ru
xCVeVSApTQtPbna5A4EE7IA09tAKo1rvWYeNQvqTG4mRUT7p6jKPM7ovyVIrnoM3
3V8Nfmr3OqY9OREzsQM8ln3uKeMMT8f8/5y36qN2Mqawtxth3OilQuLuWHNMc/6J
fuju0rI0YNYAb5pCb97Bn7od/UZHTuxgVz56+TxsxaiAgeN1JU4q6o7QaOw49wYG
eeqNHJycUDhQ+ZoXHQi86jIeXqIIM6OmrWGOPvNCHGZo7cZdAXT8ge/e88OUm7/e
hEBUK5ZV3GmOfxHEGIyHRK2OJuTQB6GZOB1yPAd6nP2KBtBdJgwzCXr7rBcxgX/4
hTK1nVQPmBjQXzPuWCWR+JBYPWQrBAMxqhoJQ9W/c5nzFVwIfSv9j6uJq8GB7q11
OTmdCsinSYILFv4O35qGE6W4Kr7I3bU1S2re8O8FokfT3n+6Dpbh/n3DADyGtOAj
+BNkQHlRstTZeyBcKAWspHPTmRBq3kNOZPoKpxKLAmUeECS9SnS9k6oJv6qXPZbE
PbNtXacZoU7lq9Qxv+W2ZimKakkxggEQFnb9KM2x11Cpgc+Nj15Rb6oxtIXG5fwM
B8XqkIYEI/odtaykfp6mmilvWs68+30W/2gR+xdAmDThztACtddef2p+Tgtwa5AE
RGOR8hhMukgNneTKt6xk+bBTdy4UY/Z57gAHl2X2d+SC28AMiLxDYQPuZq4dUgNX
wWhJyBstCq17JUvHUBbJ2Suru5kTptqLO80JdLAl47bpdpq8UdCkCZiBKstRTJEK
ROeaGCSX3xC5ywFDkBKrYyEgHtxj93x0wiSDHTaSzj4NFsSzhGSDSRmexzRTpxJe
dEgGqxvzJKwd6ortlkEqyU9bfTITXpMVVp/BBXVjUkyXUVZxp0nwqtjL7B87ogIW
wlfZiPOYi0k1krVBEqtRNs4ur8wRscMwPBgVitgKwb82dsLmQW4/xmBKDwEKN9Re
D77lnDyltakRTNb0WqyeL4JhTsP3tb/gjAXl4G58mRwDd5GPDluMWFs0goHrMrsb
uaQ+aCSVrsqyU/wY6Dh3uuFiGXxZfjydXEAmpS+S+cUzLG+1zgZMA/cil5cuNVhZ
Q/bUewGILzDYuUZv6dleyfqay7Jquki6WDCRqYzpZ0AKIJ96kIRMpjfNy8PY+upQ
BrNqnDJXII8TmixP9LR8wZUfW7Zrr+qbQQaQmYVCGe+2vm134q14U6pZUA0ehMlj
BBkAFdR/BVUGculfNDVqjECy8Nu4sMx5do6PQrYxhWQwpOLJ5juxVzQBj649IipS
bFhHo5ziVxOait7EofiI3Riziqb+h3z3f83+Zq1YHb0jk9T02rQL+AGOIBheGkOR
yIMmh4VWej/truyRo3NVZCMCEhtcy1/uaQtlbrJ97l+TrfYK93p2XUAQoeLmAH/z
PBfiGGhrDvzQRzEe8VgawK8VuakHRhJtdR9ZlEF5aMbx6b3y6xbfRIdeQAGa2DTs
gZHpHACLKDZC9+/nmDtvaFbeQVEomaoSWmFlaa/Ht6YWmHSIb+lkApPKuUtaSSgZ
E4hTd6Hl4a1xvBURaAAST7AdTZwdWl+zvp7lroOTHD53Gecj1b2clEUjeYX8F/Yy
YbUXuAfp57XsvWZ8aUVtcuTyjA5Gotr5ep8m1JCNfRLO5lQLoeEkVsWHtcn/mxWQ
XX1QseFK4TT8COLD1gccIDX6Cw1mC/xLURR/i23UYICYvJWUmw9G88B5gsUAF6Wa
BYUszubeYw+KgU2xN3zYgs+7OJdzG23HmUat6XqYUNgAG5OI7+ino1EstnanjbYe
OXQT8pw57O9maj3el+vACS06h8DNTxza/m2NGrmB75KS30ySbCf10rjP7xa8tv4n
xIquYMdHPzZ+jH3AY1EOT4JLw4RqnOtGnyr66e0gwJPyFYbqZorVIJkaCBVvphz8
Fic1j9tC07/TdHLB+FcnC9raoqu3W+6N7Zv4rFrryKX9TCnjE/PKBJZSqPCCY5lM
4yc3sydbfHtk+KhAt6xyqh4qbtcXGMMYqIjzm0e0in85JWbXX46rgrv8EQxy1+nN
z09WQhEyIaaGpfKzMxEx10Im6ev5TOau6Tr9GVRnm/joJsBpartdr8yCKt87a8Ya
jQPotpsj594ygoZAqIqC1aZXV+GLlIzu04ryDOMmCDVTC/dCmuHfYUeiw1OBBIa5
S8m8aGMxrNIcGUDhfc07UYz5ta5yqFX/7hXbNmh0vXTC0tqyXGqd0NGfQJPeWa/U
aNbLsgitRdeQDUWEr4jD8F3nZCMtPGpkKXVtQz6MeBydLXFJb1/ApfMMD3MdKejh
GyZHgs+NXh1jErEdlZ41biY4LjZtETNx76Kj9w1aW/AdTrsyLdIWK2bEwyxQfipW
NEOfRDAoAMFFIVYignC59ER/mRBHWQxtZzA4LlF7MsM38q2nu5bf4KyXypdL0B+Y
KE8GOC3JsmdbRtuwBIoDZBcjSrcbnKgvs0mOXyts8tgjQzQ07NK/tOntzWPRuo66
98ZYy59uSWTZPnWJ9QuxQ9rRsohSQmfL5R0GUmIXA/e3Tr644eu6byEXfZqdhFPO
+opByCnqKVm61Vn7Yc1EatECK3nuSYU38WjVx8GZsM0jZZV4N35Zj2nbF0LjWlmf
81YGH7X9t7yvAre8rIH6gX21HGm+jja4fURzoYeO9Fjs8cBCn6XZ8UKuz86+x3Vg
WxyzdfUsGqOrU3rxozp1vdvJaPshUHjZ3qLCp7Hhw3cEwPKXTnd8TksGBhmBz0Zj
b/m3aid85en064fn7gJVJpiyfy7wmW4a58Mz9FBr2Dd9wc5XJVX41DfTIJX/X2SZ
8PKFq18/F7j5Uen5ec5mPoF5dYKURbovx/8onhkdkq+ReiUGEQQ3TmyzRCt4ryZG
T4kHIssPYRJxQQuY0+vO9fKC190v3CEKgosNwDzBI7q0cVBDc/1pkL0qqNeNrQWU
oenEtpxptmHBjPTiHK9w/MXKe5pmnNryEcggi6aokk5X/if63vi9rbz3vv4cKcyx
6wJgn8TlW32jlM3M4NzsHvNqOBop/Ivxc7P+WgnEw4y/d8PuF/XVaJic0AElIOTa
yzcackMsfAl99MLmcNmnQRfZeDBn7qmjW6LXj0xVknu/hNPVj2cC0DzALb+nqpv9
oL7Wx8lPn3Z41hlmN6pvmSMKV9HmPtu2DckndNUVNM/wGf4NLczXXm13EGZ+vmTp
BVr+BvStFeaaV3DhG/zpwwqTbkz/Cd3LVmuUmfSSEaHQMKpL2xRWBRfJrkvUtSf3
UcQLM1SRTC9jRn5gt2LMSKehgX3/WQYk/FQJGQGUjalBl92XiqMBY0pS9p56mzmp
d58Q9CPwMwAcWbzDSUbLUawL8hXGhBFjSDwY/QBGs7aWBE4dH8Z23/lseA6MeLy2
3LEelOupEywYDZ6zK6sPmR8LPTG75NV4MG9xN7XzjgZkbs4xhl3eFl8exgcDaMpL
gHpSlozFAfCsTLSzMPZGIyk4+cslP2NmSg99zXQXcp0Csx9Gha+WveIPZCEo8yFw
gZeKuWY6g+uLc0WPTtfgLEXsNEz1PgYigwKEN3WgxPT5QBiwiw00s+GhQUpthvwj
Eo2r5UxQurYqvaWA0i4a9z2O1AGsR5/L2pysNnZoRnYJrAZZcwPb3Ayn1wPLlMCF
Lmi528gJVIB3BxCChDwWGO+6yh8ku+62VRF0Ps1LlCtlX+mkGBXbM3az+mzmxQZr
rAgszOQUeEdCLhTGJnovzG93YtajX0BLx/v27HuMM7LNHTokLnl4071pEHKpxkPo
OLmue6oqr+wOvKe5ATg1HYy/8ORYakjnEp7ytvyhQjjZBK4hUZ5+gjprsrKCctdX
ATQTp9aI8rc89fh6Rfjdkk9Nl99IrhGea2FhjFCscxi3lQe8JcJY3GuZL718ENDW
tFZ+FMoYspCOFH6VwncKbZcN3hv4YWVnjVaE389sP1PYVPCXGn2oWz+XYgOfCjCy
EbO1+kT0WTAlgLVIAvjIOH0mc6Dz6bpqh0ruJqqqutjdXgvaYPrtJ20sz0txHD/z
Ky7TnPFA8ZuevfUz4iZVqtoEJrYoelgFjREyvbfQjjvHErd9sWdi9zZ3uSfdOGz7
Vg5EiDMpyBOe2eOEAaghBaRsJr0LuFf7tCuwkSK3UF9weiBbPRTSSxTfVDhHKm6p
vmN0oGuY3abhEo7hmJs9xPHwJ0HL1EriZWsHaj+ffyclje+RnAUj8Tqy/9K/iZ/K
yz3gX18gA4T2UyHMnZ4HEcEWEqWt0NUJsUurhTvFFKnu56l1oD9+tyGGZ8dwujMa
YZ6/BTLouvQHHnHGuJbuZLArXR2afspZMqxadz2Q4Rmf+6VV1GDq8PNsDt9TwEjP
Fxu31jq6hm8h2oQRQ7OKl1UnWa7eyg37DY6BVD0WVhvu25WWcb9JYHI/N0+olkG8
2oi11M/sKv7UHCkh9rqZ6VQVNqDfn8PbKMz1P/6jm9hRSMQVFmZ2pgMaz8kMJHHE
Iz6IQC2oDwtt8MCuLcsBvXg5YecSLA4I+dlRjiynuPn+Xn8aDfdjqWSwoVPy2G2V
f/Yokx5URb5KFKSSOtGRi4JWSo8MIv2mr0RxLDUhQbT6kAfAsXVrNdEJaIfc0nQF
QTi3fCY6CNfMz+/9HU7q5u3nRuLg2CxV8yfmKN/sS4c5wPJyL9MgK1bgm1mH/cga
+tuuznYTF4vqbVDnihh2E8QMvzBlAmZuFXgulkFaDp/6+hjSMW9P9h2KOodY11XI
WmhBoJ+3gFIYqQSksN6hSXK8RccVxAZ6eVrvJEFyAc7K16K9HYrLP5EEmW2npibS
ZVLH6mg7Wb+peCqTUe8Hj54OReiHRHgUKdlrU7+X2i4rGsyIHKkse+UGJ88E/LQO
bDErMV7HH10DoO9wJ85768QCyVbHPRDeliClRJIEnsI23DL7BGCgiH9z8NAeCzQB
MQxisyizxBYfAxVwuPE7QFGdOk1EaeCA4vRy4ARxEQT4BRBwwHi27mImeRqR+iwi
MT2jqmbhO4zFkBeN8A2btPlleuOA0Mti5VSvgFZYlcorgpH0cuKyhNoDpElvPlWl
k2Rf7tyWNBo77VDBh82rtK+LOhjWrrAX8gXHw7iEAJxYuqgGhUNeeRRrDYe/KfT/
/dLiAtiIlCyKNXlu6TcaoCsvD/pUU3RXXp+GgTmegwZaDcihxysCH7c/ZZyZMrKL
NbSTWgtehwgszhZ+Vsv7OQFGPfWMIOhoEfyj6juZmow4WwDtye36/77jM79Vu93E
cYXIZLTb7IxVJJMnZJMYCdjwcWR/7EDFmlhIUjGv8silN8iz3jLPd740T10WUYgc
pQ4yT1Jfshmux4FNdGkLr06dXhbaKEXICvUl8dr64AnVUK/b5o+TDJ4xV7Iy2bwG
UZb0KYcntEai4r0woPJX0iXPM5eb1S5L4FdVe4Bor1H3zs7YcwJRBoT4sbxeqYZa
1dRjdnXhfHvMpsGShVk/Ya1LwKYtVRrQMO7i2DiEQnBMYcc2Pdig2ozIL++ru2g8
3Fn6dC50WBgq51d9M3Px7qm1gaQbhe1fNCwsW9k4xgVR15CDKFP23wpHT920wyJ+
ahj3YhhgBTXwfYNW3x9WyS4C8IFnF0iBSki5ayHuTyAKSRzi1zvkJZP90GIJsvrM
b1izCrv1GtCn3b7cmarN4t/i7oJksHCEqhYv3pgJXVX8CqzgcT7RsLaHXcZFDnEv
0xgzVR+JsQcLzBejWY0hp8J8l64v42I6TW7/Moe2ghOL/VyvxxM9OGUKoYKJbSWj
NKRnysyuse+W8LjxQ0vEtqNDufdmlwP6evaCcTsfZBUzrKCNF1tims2PptY89dgA
ZXgFmnEowgPSsdGvW+5hAKM2Yn1Ume0evx8Vkn7qsfi5cIaVt4070aEF4ng6u8Vt
MzlMRu6dEWcrOleXN3qckAZrEKU0MP01uXJou/F3tn98m0phGcchQAOip8pw8odk
IPHLEnU35qLemSe55a2iNjuTmIU+UJXODpRMLQ9AtVpOAmlVJOJUZOfkZPj4yfJX
9QpxEZUo5ZZ7s3CJgJMC6Yo70bW1/F2KVwlVuAtc1u+y1SiVxKtd9T9sG69EOqfn
emOxakbW5kKuWa/YvP+6vPX1LO/g7CJtVX+N2HinjbPZusIxLL8siEN+DWdzWGfd
z5ZMslpfJ3iLU6wgKAo9t8+H2ZHg++zUMP3T3ATt40RGhZHD320aAVgDEyu2O0wS
sMtppyRDlfgdZFEuJllWPvBaHb5ef6A63oTaw/3st+OtRfkR9l/dEaZOniS5LKvi
ScPmM6JjmnwaLhHKR2IFyMSYoXlU2MIPGLBegBOa2uybGfT12iC+Wk7sUIs347rW
T0BehCguTpnFoUh2KAY539a/kPhC5Q29MUxBkOnMWFTWtnWX0pqJ9q4OZXyILzT3
1rqMpM/Xso1NezZhSNZ3qrq+k66b6ALbaiKQMQv1iJ5TxNE1WXYxC4DR4l3+Bqz9
5fo5E7mPgMIzx40OY67TN8yfwookXXPDFEY/VpaWO5G1TRjcSC3pIOo3fyZM+qY3
y0FFFPjpgwKuMj/M14CDmCeG7bqQlLuOp6D0PJdZTSkBvwyPLbnsgJBMFk9OdOo2
4BIcCzGeFLG/06Et4hlxufZdokAtTuUs+/8s5uJV6aXx+ARqZjIbW7/Ls7QO9ZNP
BC4a3apsZbfIiYp+aps2o61f0U6WhLNASUKloxz4Tkjtp0IC3YCmnxKdHDqv3vkN
M2+9G/JB3X/ucIlb5A1NTxGg+ACn4H2CElDw5cm3MATQQ8lf9CyNpBtYTWKqeltn
sxoyVRHFzZSHmADMvUuDv090cnMkq8Ihh08NkwPWqR8pHLekkSRr623YbCCvMhCK
GfXxNHBYlb1uzdXR4SLDtlW5p2P7FxRu3yYRLkMmHg/fafV5LhSL1FtrFKtzwSZU
oMT5Vx9y+yhSuUUOAoPQwRTFDPl7E/LW/9eAiMVTunvB1IfVJF8wKo7WiJptuEQs
s/aRaR97ArlfcnEDfHCxc0an6WdScPEQTJvXOTNEyAP+QrefX23Ed5n8kI5YjZ70
/C5cM/UgxMVpCgweAH0td2pXTcuVCi597J5aNYHjKzi3lHGvtNfWPVS4ONnq66D0
2tfifV5zRgi2gk0NdSkc35BWyUW9HIo1YKBrxpbsmqhAGw3JyBMN2nhrSBvFUE9A
LKiNkS5ZNygLGwnxV8VQI86vfGEaSBc/JbnQl7WV6sMCDxp6KAm7FYz4z7q1yZYG
p2dKLuZr+1UAsPJrh+oY/s0LtaTOgwTOPnDUoEd9n9vRRe16dgVTZv1iqRnDoypH
zIjc1dFD6NxJ4w+Kt7jW7i1DbqnQE19n2/tPHIWyXEu0/u/GS5yIPHAboU7zShbc
IvMjk+IzPjU+R2++QS9E+44YBSCtGevrqnw3T4rEkXnPottQUYL+sJl5IjwS04Ec
Ct6Vbsz3ae6iUpJ1OTTfED0b2D8L1jO7dWDx+hP2L4NfMn9o8Hx/lAyWlZ0LcXTG
1GYk+OjCg0GRT5qZ+uKxdSWFKMD43+7Jgrk4TkoE4VL2aRzJJk5OuzQWLI8WwHcX
nwbcoeAyKM2WX0LdVWzLRhnA+/z2z+V4Hd0UzX29qx+C1IITX4UByLfCXIj6uJMw
MQxpp4O4NNSCi4q9JQeuZE77Xxxq0ZkJ3hoigNvp1lFj3FM0PCUr0OtEW7PX5QmR
Ehw9mq65lWO0pTlLu6eRNAms5tZCHx4HeY8WgRBaA3kCdaJDtRCze6kJAbLrS39z
DZHx6NAwTZD85PmwX8nagrhwm1g8M77kObkcLFIBLSmzoo+mV0GvhyhMoFth68qY
EPI9vdJEoiKwBeOV4vyOQYMdSZR3oik5WYr90C8m0nX7gjX/2I+FOE7zzWcqYJby
yES8JkSHdXjx9Z/G0MH4GKDuVgm/54RYrhc9JSUzCrO5a0UW0+8TVst2v9mo49Xj
RjJpZyfM/vsSBIXsiFlDg4DGtEz+8md8izSCmoRCAdIyCdv9SRxZNq8oEpBFLLJQ
RJ7nlfjmcqPaDXg+Y0XONFrusMKpdgv9YbXDCNgTfOr7a4ba6I6gJrHQL91IcFcW
prsU/GvtISSNPVjANtBeYXQ6XTIDq/zCLcT5Ww4vLDNdoV6vvw6rLpKStap9un8b
vIZE2eeOmNirTshXKyqY9Yhro6TLN0Lxm8tMOV5Esk6gklKQOFQfgjo/nEfskCl1
XB8t0Me39qC2mk8We3UNW/g3TxUcd43IDEdOssR9WUEK0VBHZQTZiYSInMrWUsR1
/0cHlUlJdME22FGse4un9PKAevgVLhc2lidfY8bcV8cEZrR4ZjXWQtAhDxPCneHU
IxTpgebWsMnTse4vwe9Ryr4CSoTbGbuQTifN163NS+rEZK50Lfkt2WtczaZ5FKBa
wK9QeVjG9+6FkOtCskpyaIabqrR8mhLyH6sEh81T2ZuoFNk+9qoUPcmtXuD9+MAv
KqNz8iIWxIUfVvLuLPaVcTqeuH8EPxk1H1PSRbV9to/XkLjbzvk7hh34hvRcQmxN
dW8vtT5fhPlO89Pmd3dSNl1PzVeZ1UCYEdAJbGx1IQA8yjM1wlDlGkMti1dS5LeS
tzvFbkf3poj8g2GZPBqSCkWWkwDHw4GdxjLSqDQD5rT/k9Q6D+GKCNjFS/9BPTVB
d86T/N+1UK8bf7LgJIarSx5jNS3qa2mjzcZbgFDPWW+FMGi0VqjqCsR78Wf0/zmo
zuJjFyc3CPoLKBf6LxazcIJit/U0y5DijltrQsbJD+Z68JsqsxaK+B/q/oPjAIqT
l6BuvyMLtz2GSQshp+MSBHlRndkgdXT3VwofI2qMtZNfsdSvCYitI7xoq+M8XvmT
PpYj3D3DblrU7fXPCesz1L7a4/8HKleLbYggrVEP5q8ACkPTvfSAu7mk26VLniwR
/TU9JieOqqz/BPsd6EtWIWUdIqXx5PuqjMVb5t0OjGcShDLK9E0srXKu3SOUOdKd
oWPyq8aQjGnAzLJTU7TKqpm0Bh42NPpp0MgpymqSdBkQ2hwr5USsdHMUtRXkCulj
i3GpPy8w0WKYr+WEB/8t/Mjny5ktl9KgYszwA0SkJjGUT3AZA3yraDUdZJwgomOg
XjIysuKL2ppf0zPkKxxqa4OhQJlbgAHYMShP5tGfz6MXWQgGsTDIM7NquaJsFQO6
M2EJ+wlH+EHPsce9q+QC9A==
>>>>>>> main
`protect end_protected