`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3792 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
wcmpwSk7Xh2DEFViwcIwodbbDLmZ7V8Ty/vbMb+w9eH4srpA+IXKl2anIFkEV710
RxmiAy+V7M4e12UY2XF2CEVO9hpct/RAr/q1T3Yb26Say27qMG8Ro/oFD2zC4pXs
ADWesRj2ZUE/rdXo9CRb3Z/qKVvKYZf45oaHpO0WegaegP6an16Q2m0TTVeatoJs
0+Sk9Otv6qaOe08hEmxszEYzQajP0SnL2XQx3Am3wpZc/34CKCgutEEqdyS3wXby
FLQ6RGjsSRTp79YxgB1a7vqbpZ/knOAhDisNr2oNgu1+EQtp2rH2skl7BW5Tpj8J
0Nes8N26ECjyn/hja9d7O+RTkAweIDF89/MGV5xeaf8ksVrShivDlSE6zTVJ1upN
6KgQyrGcTPStPGGJCEDYU07M4+wH4h5NlUAjZ/fTRX3cVMt/g9fuCXKFhYEQ6rPC
NaaKLLqQRghGhLHHqtouPkYCoWc5M1HpvKWvOLo5MT+Wgx6vQRT94qo45JRYFLFK
U35FlwUB8EF0PmN54Z/4FHTrFjbSoBf4AGWY6gZsR4ulps4GSjp9cin9EhHQe7Lu
uVY5lMqyIvCmGp9Oalo7HN3PQjm/GdaOc1Q4Ie+fA2rvWvoaHKD+tcfJ+KBDEnZz
b3KYQVHiIpt5Kefh6/sgKG2xuxgYQ1EL2HPmBKF9G6c+1uznHbonpVi6+sZP4PaO
G6wANZFnQXn5LeS33naY3HAHR8r0GsXdOHW61pCgFsAm/+QivX7YMjBXg0lmN/RR
1eXQpuE9jqxGPKXhlAQmTgckH0BMoWeXkVhlJcd7EanHND7mGNbBcNvyZvGSpsJR
sH5MlmLyNWPBdtk4kmm6Zxam7J5yIaOQF4Zf3X150JhLrGVSVOX+nF4VekuYGJ07
1Xv/J6mqiemUWILlwdM9WRA+nXdzPmbTD57CekL6RwdXkz+gIP5D6Jj2IFyatBD7
6vJopS4FHQh78xQkk5ERPVLUP/O2kMmu60/5heJGJ9IuC6CvR0durUifpO5HnTcg
FJjgY0rQ4CUdwgpbf2AseWzpwW6Vwlruf6lueyz/i+57ng5gQSa8C47ifMySedM2
Kp+Satx6Uk98jRDfvnyOos9+R++JCPCEbPaUZWURv8+d4z7YCXJqL9ELa2jY9ztm
GMEYcyIq5d9/jQbvA9icUv3K454zaRURhHt6uZUCA7vL0TF6hrT2nJN7qFhAaUPc
wryvIMfUXOAp92hx4GlYdy1uIcvspwnP2daY8IydfrXORa8zXF9QLN0bD0H5/aAy
onW+G8PTxKkqC7g69mcAa+f3T9h7MSb0zGUz9G14h71MGb6l2GK8HTIMPeV2UGFN
+bGefMWOEo8UioyDMwdYl8HQ0yl5u3pldmUPHyCjaLqTicE5llX+/MEHiSJBc/1N
q9LGuGnaOe5UmZW3GSjh6kXEMLM+6nr94l6uQ9lnHla8vfwbGK3Gvm6sBhQHBkjF
RvMF8G45Bj/I2xdOkQ2FoG1JIC37YQ3BN4+KKpby4Fe/zkDBIGH24OkktV+KTNT7
ppsmGwSnOadU0Aq1UyGE6BAWBcaMsTYpv9eWS8HCmEoy4Y3jbRuxvKb23IwcCPlL
X0EugwE9u/arv7lfw2JOSbnTn10NpM4YY8+Aet23G6CwenwNI/pq/whGJfA3xEFn
Z6WtH3F67nMEM/jxPfSodrOy+6D4RuWK2y2VVO45CBHkn68ZsbQSOPTM7bnUhrRx
SywQaQZkHK9g3gJeJHDdjbbFlMu5SgN99E4UIwwWh5GmxTl3RcoukwEs/lOghm34
J6EfcQV/WNSGqdhklWyfy01PK1ZeOMuo+BeSYud4+zwODYYG4TpCi4ERr4IxExGy
4orbSR8U3UcwYxSXyn2ig1LNjcRpiciYEKgkNwZe5nKLQ7DKo+ELENH8p4MnI4vg
4l690brd6phg1dnspcDN5mdPF+EgqrAYFDemvT/BakltT9czeBi1saBZFKwd+iPL
PpNAd2TGow09ElfWmJHLcui06bKf3c/fL5dA3/1avU9jpH2OthJG3MTzS/v380TE
5PSLLBQZb1LNAk+KZjOw9jS7Uw73HQ+IL2FQKQ2RV4+BOg2m5w2BUU4n3JmWUR8f
84eblI0E2LLAOAEwKvq4db72FgPdCWoTkp+OzXxMWvv1YniHo1/LfBUOS7z4UWMq
YrofU8ANEf00xJiQaKaz47ancQ3/5neEvWwBx1eiH6Y8qCppIEKMgg0GwdnTGDGd
q2JvHAHGpBrw5WpHFPv9E7hJwkuBBlqxfiNKmO6AlpyrlrEZ4rD9vqhi0w3Bt7XM
BWSfL9tnTPm7sisoB0Qrt+nIb/VHfPrfoC17kxrZb+ksfdK1BJd27o+8entbdwpO
yvwv5J3der4/4q9p7DA2frzf0np6FfOVJAPeQHZXyvgv3Qspw5ls58rHLug7Ae+4
FTWmHQnqxK0J1YyRLXprgRf6WDN8uR6RMap+5fWy1iDU6iYqnsVj4W/mkU7GVcfR
lBiOL7bDWOro43g2nDa/dWsGOWfXv2NgiQJ85mvam0TZyAkJom/ztlqEw7JeBLoM
qyyv6Ae9yFdvLtPOQSmmfOnnF80imDznT/tS71QVivayziNNjSiFvOUoPIm1a4GG
aEFjQq2c0Rsdj+INonMCsqoDSWH+/zhD0QfOpPM9B9vuQuB9lAmtmrQfRsWSokTJ
O27AW6CI5jntK3zuH2VKhSw0x8o/aIf3UjGnJyc8SIddgRi/pfFYFzFKwSHUKq7T
5V8k5sfC2Q6fEhHVE8Sv8OzqowGDSEEyDjqfE330ZjPdmTEU86oNV0x/8n5gj3Ch
TdpiPLZJcGl5N/SANoDHLoPaW8Bl4kGoh7MazOW22kAowNJofKfHjesT9hGf6EP1
8tKnFdJgo72gQFvYryRcqXN8MBNschuYETwKEjU4K2Oxgq4I9LiVPS69A9bj5If4
qxjH6xidV0djTOijwuqZilpF/UgwK08H2iC09Se9cGXyQePo91NLdRXxxKM5XzNF
lQP/Q8IrO8Xdvk21C8Non5nSAAcqM5r46N4eludx62bexA9lucSpHy2q3VvOHBB3
ju3/aDb923SBM+FsybhU1UQih7WE5wJYcmeBrGBMxZcci+kTvQEuOslOwsl5rcVh
vai6y5wvs8HC32w7WzfuantqG6AfswSW9SSeUF+zMLrYcsONI/E79zBThAAiJanP
YfzuC9odA8HWZNvGmrfqPCPu/V2cTp/p2R6oc5+aolOrMqBAaAsEkeIM7oKmyJJd
q2GVMV9ixXyVgQJdsUGSqEYM8UfYjCwPAqAHO9LOIHN6vCAmvO6npVRB2Kbe+7fA
Dhcxpa9XC2VhXqCKJ9mTCz9ec7oCvdzBV31NrC0Yz7YDQXuD6h81vefS7ZhhMnxK
JN1bPnWQxhkn/X3sUH5qTRhduzsfVSL3z1AZfFC9zkVldJO/ilTzB/yeXmhGvcBt
IV3u7kTrc1Ijk80Q6cS51ziz0lUbRYi+kUiUvD8vroa8QKzf+K46o+PxwBD2FQRu
XEDGE1iJRilv1SRrY9cjfr1SBXoTYgqO3/SK+vggonNIeGn8o81PvNmlQf8YHpFb
I+jOf9heQbxapiw1Q5op7mf20LPo/YMWVz1XH4DkWcwDj+qKXGmjuZjcukC7ZXrp
B/KnLc7p27zGI3zD6u8H7RdI8X1yld2OF/pwRp2M4bp2g07l7ltsvvnexR3dTnBL
Xk0dszLRa8JbZGQlBTWVvA458l93G+4ac8KkRF1d1O6RJUuo9OvLwlh3Pxhwla7E
jLCxA2wWB5GGvgtMG8OC5JFreLuNogwOwH0JEj6nntHhfIN1+C6VGdjXQME3bCpM
QEc4BPaeDopOcHyHB3XomEcZV/zy6pJAMnOcdcaDoLl3lbI4cZUmjBrWC4hRgnwD
jK9KAwM3uQ8qI3A7oU9KW0duN8xr+I3lIoIcp9U4lAZ3WnqaSoYCDkKKVpdM4VZR
PVjM14knzjKbNN+/bwWunrpEiOIwbSqmkn3DkqvllhgQbmqb6VCi/RTKAebkkqE9
S3WetQnDDWPlyfWkiXlJAmH7T02BG9gTWDyS+NcsuhCjyfgrZxWGJYhsGjcUsuAW
81eIh1WGG095JLOYJBBKDboSqqY0qZd6AaYngIX/+4SKYmbz73VfH7EvEvBiVVP+
D0YWZTEBMYE7z+bRPFigAtfVZd8SCTfoZdlfnf1HbRnKsah6f0QyP4IyMPqOmue7
JTQJjMlQEhPAbTN4DfxdBOjkVfRcDJBmnJcL3F1jCnpiWWrybVUy0MEs0oecFYzF
9Oc8WgijxiBru3sfITNEKgGotdLpD9MMxBFkCJV8bHOJvq7BF7OOrNhcye38xdFR
EKQTSNNbs3069xwALH/fbd9kEdvzvQEK1wI7GP6Nmi3BwP+pxOVeB6AEewbK/Lvz
3fl3I+GKqAP1JAeAi2tC8mugPyHl12PbtvuUsxxgeSpr71hd7xKHRRzoUVJejfdZ
tGYq1iSqKzWuCsNsntAzQFiYJCMOJ9VpIJuzeP8uM/id9LCcpVUT8XFpUq7t+R9J
I2ysYA6FjGbDFbYtaONyJ+6YN5ceB9SrIYHnjkDMN6JnUEFeb+WW/SMhDN+JyoQW
r4Y1ayJg72q4e1XG6UQjtHAmawR/KQZgUsZMsZM5+9ZZ1vcY+NhlBF0FHgUAuLXf
CusKbVH0NPKtNotUfh4p0IM6+cZf64Mx2i7W3rkVnF4LphuDHBuTGAxd3P3fOgQ+
QfqJf+Jn/GgSdQCGndA6+ZHKsvAW3VayamIj1MkM5oiM2VHUTu9ryHJXRc4hE9fq
zlaM8XaNxTsK8//7QvT/yIyQbUCpbSnUiFCVwJJhG9B7DoR9+HUceEgWRdrkgS/j
TbqoCzAPR617WYiVIqN2UR84mA/w0LpfmhSYePFjWQ5vbslPRhktRtuLVyBW1HNh
`protect end_protected