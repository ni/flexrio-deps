`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1744 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
xsYj4ZwXcxl9cxOXlpzXHdTeGkd+v4WO0XoKt5XYAYAMUWumAXEAVHyIMySiNXRg
V4eiEUoaxg/rwXdRmvOZBDuiE5PmjmJsdLKasDUVJdKjBPpI/eTWk2WgRXC/syyE
zpTK29BSezSLml1nk3EM6KenNj6G9H7onrPOUZ2u8IRIW2lA85t3WdE/9OWEkQ22
U8iawpYinq17L6cD8M15eRzUmXRT6qKCvinZ/zIjOXaw/eZnooR2JpfSh5fj/gi/
cYmX6yNWghkrJSlHRPE5/6iTJHI6fZy97B4lTEEyUMoImSkXFs05hTdOCT6zEudF
UIpY2XSwSS4Xc7+pfdnwsKGfcaoelHrt/hVRx92g5pg7Bq6QBHOzyvgJ/JcG3aFS
P8yiNs0OyUDUTcD6neZ/l4rznkSHzEsMDJNapEuPCkM8Syz/lb3rtqmQZKMCjQJJ
iS5CRL16xYcc483bioaOgwhEztQJ0y/D5uSZIdRsDElyIILQiPNTb1ahzAvF1I7E
yKcozAuN9wsqpQWOgwEtgXhMyBvicR1WAMLGuYcZG3iymwig9TlYcMmj4chpuNqb
aGeAifHdxfNhWDZjbGFSNKrLDNzSDXheDiCiLLzZlyZf0lAKD5wTYUZd664BLTjb
zUZyDsraoVRmGUg6VNA8iKOX/3wF7I++4Ym9hh6E42jDTQpJpKYN9tMoZBBwqQQ5
sfslOTobzdUlB4/aYE1lPJ5TH6qPRO6cFsF14tO3eflLIwOEEWUwM7OHvSjhr+E2
d1d4+iZX7AsznDCXp8OO+BjH45gwxnnihNNAgAKvARO9A9iuMhdC7FlIXbwkP7aQ
3J3coeP9fZHHJKst/wzkwQMBp7HpQrbh6MfZuVk3RIQWk1/JzZJcjOI78i7+K2vZ
9/75YyBxua0RderRcpFHeN3/4aUEl5XSLGifTPgUGHtRukUZBXDEGnlHHBq3LSac
ehUuXNr8z5+ApL8Lnj3erIK4UmK32jKQ1Qv4J9H3Rn1TP+txTZ3CcS2qtdz2esPB
pGwflMwv/wp1kd2x4yrr4q7BxLSGmoKp/e7AHDO+W442+lHtAuY3nKmEZP61FJY9
EstJE7MQ7wO7HG9kgLPuw7gy1nvGE1U7q8PUnWWGHEAP/RZNvKx/u5i0Dj6yriow
zCUS98XdNIryXG+l0JD9bN6pHhemDEgO7+IBc7tctUz68OtuwOaRQp+86YLhR/sK
YNiJv+XAO4CPELA9aIROOf5BaCP7z3qaME98JXpehWb0+feYyzEeJR+tJbqIHXpz
JfG6qSWrqnELxzxrkv95BlNGtNvnG/o3uwH5q5DP/BUEFWyNnsQGepUafjADDTdJ
d2/2q83bcsTh0VICG7FiEuBmJ0CXBzqpmVqxCngdtEbXlMIYyXzGvjGIc8ecdyg4
cdVW+VLOCjobZTsot3Zqo0/F1EA/bg1dpFHxu7DHvhCrDN2b1MNQqL6q6YzuLFlb
V64Eq9fXSdxOhrx4SnQjjIiOLOHVuVJ384+cfAB1LUDU2UW4yHz1niYPtgyf8aWw
Cpuif0rRJIPY5MqhQObL6M3oiWp2NSgeU3Gz7CqcKJpNRztRZAhTcDSMskaJAhzk
pJrh0IH2myfC/NLyn8yTfyb5l41zem+zaJQ52H6Uu3wh66IsSXtGLiBZI64ICFVv
ImXf5dabqGH2XSD2B0vctm51leP52rW7/UWB4bTx9WFvG8DmSbzmGkcgGAlGIssB
btXMbyct2mWd/4V6vDehVptf0rV3txG/mkUKrqZPI5yagQaF9x62WQvbBdMBRhok
rANy2J5mJiohwjvDTSinYCRuCnD+kIv1dD9pIsqViqdByOPb+oEluYoQ66Xyi30b
wCM66D4HQTGdev9jGcKBOJD3R+tX7mFlkdSkMXd8pxrvsQkxiaZx7UT7ZsUOSXMJ
+iP4IbzkkVsQYQiOgfuiP/2wMBTRqulEn5kY5CLEw4EskQGPJklUTwlRBD3YBSXw
azIGI7eU8Wd2INBmpMU7PxpxKnad4aiLe7mqFZF/7UZLTYTOken3grYMgD1zg46A
UPhS5vQoKWKpLoa2ir1FE2iP5YJTJQFsA93IgXGtk84bF13HbGqM0V3t1iZS80cK
HAWrA4PGogh3F5+/gPd8zbv0LbLVm75viG7wpe08z7rdCfo3shX2wU8BWlXNWv2J
OqY9blh+m4o4ZNrqoyBqgQ==
`protect end_protected