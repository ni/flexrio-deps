`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10368 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
FTGcP7VlpSOhasofAJvqcB1qG1wsgtH1+m0gFKduqxaefRtnMhIaUPS/2X9ELH4M
z2mOF4k7UxJxfQ7nIIQ9adh4GXcwE7rVEFqW/8taOAycmitPsGEnzXk1FZbySjXi
vhJEiFl2JkADmFe3I8LbP7OHD5oyM1chRHGpWM188NO8mWRzYmUE94M9l5vdK33q
teqcdkBTcI2z/zJFaDxYyV9L63lk23LuFMZeH4S+xUaKtWMbLvkN/GYk85qJEQpX
CCB5Wbau8k0ZfsYGFT8o0eLMU8OF1nTj7NMT2ri5+2AYkJGUQzkIeBX74KSwZnDr
VdWqQ3xb5K+Guh6dhXQQskMVkmhSnPMyHP0loRYHrXkDNxbez/kxWVUZ+GZHhkO6
aNin3oc6nHixbz3+SFmJ4eL/VWXGdx1C3OJZmXHLM1LfaPSqDX4YblykZO/Sc5ri
Zxrn+3SkE3h4j//bvklD+fwivXkZUauT7kNpGmaXH8C3SCMQe3/CIvg9pQvUL+eD
ZC/gbayu+Zt+HhW53eyad8ihJzhWTXWDAJMFdnv3dgb5eXM7MRMFcULwGLDSLVQt
kerchM410MTLow0eT++iLSk16udZkf/PzqyvwpyockFtM+ydpemTZigmuUWM7KTz
cJDuMZYZLvHcE+B/aEo4cZziO8PiuwdvqNUyodU2m794/Wk4bELis81vIWfFHguJ
3ZgB7upC40jIX/fB0L3z3eNV4JFV/xO+803pVsB0d96iJMV7TbLmVjWddTGmZgDl
iihDM5phr8WP5M3cNIb9jodm3cL8ydZMFIp1PUQg0edGEeTnxICL90WnVw+AcMjJ
/VU+VjRI5/X21SLk4n2BUHuMIq21dkQ5Tca99FNpwAvDm69Y8kQLyLrpdSmyYIcn
7QmT2eRYOjkqZEZEQaZwIY5DhwUtTha1R1hbqG1nA+SSIPeZgkSHpgJcwEHUPX9R
DFdBBDJ+KudrOEo6MFd5WdCv8acyA8S1T00/e3IcbLks0xZaYX1H+f46029xiW+E
auXl/PRaMSH5VKyIxRqStsGT9EWWT3PbIo6qWdoxU7tB/Ynrsc1MhGqVrMkv0hUI
emtHTOkiOAGvAle/1QVV7wIIGeIWeb5ETNBEnDuUZ/kkQ4fn26i+aF4Amm2FzSgi
Is8W1JxSKizKM7BZvO6RBejBrPaSEOxk0GpSzN8LCPmG6ykaitHzQrJFMNYm47/O
cGPSHe+vmF9xuhsRhIqvvXr/AnHS5f0PucunBMDUMte465iHbkrGkIO0lRaH1mpz
BhIph1bU6zpzTcFDs6EFDkk2XFTPuSa6hNwomAewWYOuH8wsFlEYn7Cal854M6/R
2saomtcQywR/X7bXLb2+E5YE7pFxo073jHUx5f6y+WVnvfqX7o+jlPEByrwfE1OB
Xby+wxQaf9NBccF1TIPmkodP1mhpbn0pHfkx4laZNLYi8Ou2QfqQ0l6LpligwFuH
gCVfWEym4QQrikiKrr46K375q0Lrsyhp3BHkriV7xZH5l7FrFdbepozpD2CjMkYe
pW0LT3WgCDZdo0UKuZugkjtFovV1BXooulZ7t+ixcUQwI4KeIO5ihVdQUFyrJXSy
wgpk+jMbe/AnqinJe97bqrQtUax5O7fcHyRepHQ2YxYMCw/51s+z3WcnAmg/Co10
/zK17UFVMTiMcdgVKvI05anbtGLIibz4Cv8Hd4//mbD+94yN5X5UCfApyj5G2BDs
bYfjGyjOWstEC1o9c6aLBFKUa9ScFZRRNIw07UI2LNPwy3065h42umnCIuF834Pd
uF6ASQ9vjtqo+MI/Y6c/EBhQtUKqegaTEsT2yGjEScMY6mpV4qkFem33uq2MqRWS
iG8w20b6dYUFg33LO6eyGOYjVlUpMT8rK3ia3Uup4ArqOOooTryblYybvIYeegPL
ZkT/6PHN8wpiaJBynikHE0KZ83QsXbdinjgkHEl/16Xhs0F1ZOvGbL2T2hoKdVrZ
AF8qZOPP0ooJi/3bOeVCQ3X6GWO6t25jygAbB2DYwQjD5WW3n8uuUpnh9l9LYxPP
SlnIBJaEoY6Z/h4ldeVPRExBl9O+VzvMZOMPlT+efenYQV/AT/+0wjPIBNYgfoM1
KGPcNbB3R4JlzeTE6rhZCHDcvw8TZ9582C7QB49I0SmDUItS6S7QWQ2Nqmd/A1Xx
2lLRtYO9LSc5K4q55haC56wUMfa3KQHnkUsbt6hnWMGc6xEmuRlcuDb0A4ZVQFLW
bvSZtFD3BoHIN5gCHI56L6kJYNj+jLipe/hzjpQFAyAO4wHBdXhQwDSg0o/ffrff
2ZnwazWIiV20M2rHjuijzY6BtUM3cB471+YWMNJESGVI+qig9LFq0llvKgNbufVc
n1OlPwXdDbiCibKttWft04ZLF/WFSCHapG6jS1vOvbF4UL/31dYBkvUo+omRohPc
jxpzB0ql2GUhaONLCcGx3eseMgK3VBUznab17ViArF5rrLxoSdICu32w/WGPS6N0
96/on50CgYzKBdmii4XxEaKPi77Y12ObRA3FxdULs3Yc33ihfiEfS2lTFpBQOrDv
XV8c2oMtolnFkQbWF1v7b6zQk032NxFNuSoVqMKRiM+yqNMAKSxKuYFIOGTc6CHJ
ky+nJKB4Xp7fXlOIa/S+arQizjrFzwBh73koOZtl5hkEwBSKm5l9x6Ze+9r+lt9m
exybiiNF3m1JUgXqLW26DoXPVFWuUl3oNLGJU9KxF0exDtp4DUcQtHD8DVYJD6Us
uLU4O1PzRAhaVBbS2EpOwOjblQugvtnabhZlVD/RXXIIaEmA14935pQOX+KWAT15
ppRnaftg6Vie4tuZWJEhMOprqxvMxU45vPAyGUJU4hDfTzeOd1kXVx7QcllTJ+Ge
7SokLcP77ZwvuRsDiguNZ5Xrfsh4ZeuhfJZuCnNW9gGyea8mlT/ozqRhjQkIuItQ
B0bL/r1e/p7eEPkhrW/9nKuZjf6E8TYtRsn1mGIjbsxTyQEyrzVtEy8H+PX06XZZ
Z7gpnq1Q0C0Rd5zxvc8SBdCq7f8SvQA8ROqK5VWaWVHTLWiOn1Q9ANu68noehsug
CRnptr46e5oQesDtLeiTaMEyeFJRvflpL02GS8eBbr6dt5ceCLZ+IkzolQYy+wyt
hXiFrvzUAZq8Kim4RsFtIVEd4Uq1jLPx0TABfjHt6w7UTUrIiqW6vctBIixjfRFO
Wv6ZVwLKfVJMcRbUp7tQhoFZ9qWEhU765WVG0zXCWddpoL1y/68CV7PBvuzmKLSa
DiLdsFzUavOTzH6TqkrRh+juk+3d+CarO2PHs6N3fbC/I6GFIP2nLElcM6GUVixf
dJfzlDOdfDGUiyp5ZequJX0m55ylBhwQK2TLWCMqQuaoqitqtBeWWz+0GUk5frE/
pTS8o7ZBzOXwP+MiEPrULZP0UEOzIp+bpaCQYv6BiS9cDyLis3AxG6ar/V0OhuEp
wS4X9FUWD7gBwEDypE+0RFtm8KGHjRulI6YThwcx9HLyGieHfxgsSo9zV+GUDkVy
WbLGASisgWZ6/oQOks4D9AuLdAFXI1UxvyBAuNmlbmrARKRlGV/BSz+OIJNoeQtj
wslwDNn5Dm9vFyi7nlV4XBHJeaNYjy1Vg/IfBjiTY03Eg/8fYrmkZws9DGlihvkj
7s1JjhcN8OGHMQTJdPPQusKk+cunNLlg/UaLEiilx84sxmKqakhCEvbqxnjDdjGX
kdAV6ADCR0SBv0zUsUfDHzSy6AauCj3XMQcLBDk1EHCQNHf9engizgH0CR4BYgXG
tGceDKKNfsLn9hv/VOZaLcFc7M1Q/ElfcMqHd5jWhj+Ao4Moby0P3wLnmGtt7ITT
elhVocpPhNYWsbA9Hx81El+DWY8+189x1LFc0gVLT6X7tUY1vVkpCeW+5rYj5dYb
T/sDLMI6v046D4Mff2alV6KFjwPw+yiC0Qq2AZQAMdcblcp4Z/7rlegaJvSU+bCv
zroOnYiTJp/LhRtrKPdPzaJ1O/KgBXERW2lk8ZwVVX09AJf5AQuRoZLNVakonzKa
3VUBbH+QloI1gSG9PNIvnVJbP5//8xa+ERDYv2ba4VbNIg3GcwtXPW7fwIfIcAqJ
LINFOQ5mmEbX2pPEgunqlh9LkUafnFI6i6IbinwrPnJibzY+74SRfgImKQOV6/Ss
9kCxOo/3TSaEIKWwjdkka75uKVSc5XVmKOk9Oky8+No6JFlB9Ogz0d+m473R8lJv
EXwGjPJl2RpPd8iTpznFTcF+ckTtYibgvH2oWogvIeLIBbhLt0vFoXgXfLXlESGv
lwaQVKUM96xPSRPonWiRkQ5NOS9CsdgZb7rzTo2YubO5CfU4NnYyxPUI5ee8EeAY
GjWBGL/gUxdBkJAM28Tzb4wwdvsq7MM5ONzA1JpwloYBYTYkAApaiFh4CmvhIU+v
Y+gi4YP7R507f/nxEQYY+JYpbSnlPuIst033JF77Z6ULd997y3/nQxTTf9ge1jkN
yhCMipvQcXgO9t2jTEsLrZgyuHvWCyS8A7PoxTpdAzA30m4aQdfP+XMx1g1joFHy
+S6S30pzMTMgD8X9okCDwYRktfy73jOfoGc0EWr+trRhB9pFCL5VKSHNsOn9h5mX
lo7xWUyw0gkrNM+vXGdZTYbVfOuXGqMlQr+kkRrr8jR3RlfJUUnN9Mo+RKf9GoF/
ZMrdlsMY5Kf0KkhZ6pnNG5wz8W09slhZrWnI4cV+sg76zRsWcDqNofSK/tjOu9BE
D+x1j6UGQ+B7LJ+GplzMXFjIYVruHYWePGObJrs5cyRRFILbWuZVLoKced2ZAoox
Qw8s/1Bho3rwReVVNqU13liAbtU8UDzbHx4IKea+dSXvxbtehBf1A+ZkV+JSCoSn
umNLuks9OQd/P6O50Fwj+27ACvGgGmQlC2keNXia4ucrrvUVWuXZUxFpeXG6vFlt
3zRGxxCNVNHZ1SsDSNrDWHsvVoExjRaYMEvh7ZLkx4obY5pxH3wn2eHU4hRtnqsw
uf1ap2d2+EEUQZ1ViHO+j7XOLHGKaPZYW2QSQOTSXL5KVxeOrOPO1dgguLGChH8g
n+Y8tyWtctOHTHUWmPePSTWqqRKP/kWrGG+GznJ9GpoNqGqIGd7bpyof6OPdAu/L
DW7vcKwE3YpG2CUg4t6zI2YifTK8aVlMvdyVN0Pnk7wBxMuUJhs2hAWwedQ6M9WJ
MF3jkFkqugINOWW7ryungvSPJzAQpX5x0lLpApHDQTESA+MZWspU8orgv1Izeb2a
l/VgTZBZivb+wdE6hkOj37nZfCmGjz4tHLVBBIQaO4GfsPje5QZolR8nupEfQQGB
Q6rzKAbhAO27bupdVcVrzeKtPQlflUajOvrevRBGFqryrluG34cClOI8GkI1PvQ+
nHqNcbCbgR6bwLOcdhstRX8Ixkbojpd5RIRHPflXa5w38T6okrYaoXV/GZi9y14Y
ipAcnB6ns429TCKlIu6kAiAwYN0MDNuMa2j2efUXm1gLKJpQh36tMKyudRpDo/FQ
Dpb7uh8w6Wa0fL+DYJJ2NP+zoLj1wRMbjtrS5Uj3p3Y9hekHzb91dRVzB+8gqo46
qfqt+xFI7JWyCgdVYkxQeTU4Vip9oKHym3vjZv3b5eGfnUEcoHsWKH3Qny3kQ6Pt
wh8wESlAwJMeN9Lnk8p7YA+hARDEIYHPAwzZogzuKd/Mkf3mQwVRrnwoAb3XKiy/
MKn4apf6/6ictuwQK6wATBsn9YoY4FBcXILXnzI4TYMFN6QH+KS5mE+aZKPSDRq6
IXCnbvQ42l7wA6rYrTj2dQlCGBGArXwEFRg9Begjw0gAXtAnz1ph19HUCprj/Kbw
1bz589FPeYVk+7+3hbGO+mrTKOhJi4P8v3tnTcckOvyB+f4zCR0+DhyFb7G/yIJk
GugfoeiAPAiuA0vtxK6ieBhQBSm7w6ELuIOUYYlVrhi3OGUje8kCf2BIniNdNB7m
ie1GEIGPne3QBDJkWZYMc/ofd+p3t8ngiGtZxNB/2l1hz2ALxQNJrxl0YrCCy3Rc
Y2maBW1cp/MoOLI0FlYTJ92LOaNvkJ1Gez9FcMgiP5ogk232GxfUlG8Fk46JE53B
1rELGDKDqVFLFg7lDTcIw0A939ySk24hmdZBuleJW57OywaIKFqf53PazQIOuJeF
iVca3Irl6cAesvdHciDf8sCe0zeMMTGupJb+cMCiScLAh+Bo0+cWB9u0Y38I6fjf
uLzVQwOpCFVcxUoSbjO/oCbzYO5Mh5yxRbDuy5UOY8WYeR2Nu0XObOzgLzuErlIk
4E2RvhX2YNXNzkT7DfSlvtfdgdtroq62dT7yVsqee24zOmQW9ZEDo2DRlx5idUK3
izj3Wy8GAGdyPpnkwucZmamD799ZDqkkgpoPfEe6LqZtYF+8t9mXQ1wRGYq7byy3
RJjhrPX0kBRN9VJDr+PTdR3Kd/jaodDv2WCVn47NNDPdZ63f+GY57pjbU7h3hfq/
RNp/L2i1E1R+3F3Ti0g4LFAWwbNT45bx08CYbZBZNOTX73Kr0FsKpWoeIVv6jIis
pWvd3HMjy17WfCJQODS3g5AXLqUt1owjjFEtO1EV96cyaoVVkjFCYxlvxjUmMPQ9
/nLSNHOcCy4lkgNqOqPTuFVpNV+Oc/AsyFDh7siaMggMXJbbZ208vNejpH/Bt+Uj
/7VFt9t1BgcjaIJbQlLox/x/AAuJryJJIKbBR1upm78Xd7zepD2NgI/KgpeEkla8
E+trrX1KPjlhOLv3CCXqJJkxopEQhtGR//SDljjLNgUkmBkHWhK3FF1inKb+PkMD
7nxngNf4QzJ8vGDjsGvxVY281bZjMruyT9QHvy9kzMZXmpN0TADuSSaoScN8AQWX
vNpmciUr571fFfTgMzd2sQGKFu5EL/5tu6QIogSPXx/vdjkjxHj1M2fGVvRSifLF
RbLC4QsPdzWkjMGh8dYg7zug5PbJF7D3M1/3YxT42DXJ1X2iEoV2Vhbzga16x7Y0
SZu52yb8Bv6uZ3NOMWdBAjbAXy4XCxN8E6qT/2j3XAkujCkUV52515q1k8S8jYjc
6vm6pspAYYustJJ4hzbT5+bgMQpM4MVSVYAgPBV2vfNXaoxxgdZrCEeERNnYQ2DL
DPLZb6Oqm3zRt8Asqpkj4POVVJMtT/AwrEmk2qw1XX5eRXgkTF6RHTh5CV1ZEft5
rSoFZNzSIxJWJaxk93O6AIJ7jzmrcfIX1uoAWFNp1nf/i4J9qPl5P1o7nl2crJWQ
rQMGs8gFywu2UP2keBEUg/IGWMrJKMLoU1DwQ1XjjT+suKkEANAWm7bO0bDqJpSi
637Vj9/KlmqekMzss3e2r47LuthdtBOJg19wFxzrydfiAd3xokwbF3Agq333pF96
ygI/kjSo5yPb1hJTdsfPh7Zaam3Uv5NYWGqrnt0YC6ojzytKA0Xnh5NDNyGzE0yf
2gexLM/p5ty2PmlyQv658ynoiDuAjHaQIeiayFbSBAJ1Iuq9MP7tZtmQrz4BLeN4
R4BxhJ52pRtsh0JLYGf6XzCE1EStNbda5IxpunoBf3tsGE2tD8yexQsvDbNvMVrl
xdUifpAzs410uEnG4FpNrmiVcstmyn7fTysXaGfdGT7ZFBdU8EcgFaqVTBJPLDlJ
w4YC/7WIKV1TA0QBOpIWdiLLtYEByflRUhXSva1D/Dcf6skIRaqb6lMKEIESy6j2
Bh4G5S33iL6FrLOEYM5GRhenuXa8PsJ9ilBIHkuBiEaEN0Bc6uwHm9XDraYY8y1n
bcYG7qzbF2JQrSJttfVc9hURsDZ5V/ZqnU6YQdSIYB10vZpWMU0ZFRzb9Q39IQbR
jtCaIQEBqaS7npjr3LEPZsXlLQWfASGJdI4/HrFesauURCfzl47kxAr+diHnc79m
ZDyvtyz+vM26y4yNcABineGtzFV6HKfmZel+uLHzxdNfn6XFOZvH+pd852YAKhkL
SwDwzrXeadGj4Wyib70dov+387alEg0emK5n8gGqyNFIgeFBH+4c9pXj7MMcxQ0f
MlJZjYRRPa+A6thbvQZfnF0Xh4+2nHdCPBoB2NvLfP/HIIpjRZJesQDL6OKZgIW9
LlHcIfQefevBJsGS0otl4QkLdXXGoj4C1AQhyNHTExTCE5gqTuw64GDR7Ikq40Sl
+09I1QBX64j5/j7EiUdc4LX043e9DbIho9tqcY61mBR3g1XJm+eiqN9KHRfve3eL
hO6maPEzRF/zg1IAMNygsDKtRA0uovsF+gQx87ON0hmZw40Bfa89XLyP5o/QScx7
DajxolaYDN/rKOdx/RD5D5eJFmypLjBI3duqK1laBn2lWsyAY2SPswUsAv4WJWMc
Q29WxXVFkEcYWCJW9xupzw5YMtqQ8XsZeHypMKooeO0l/3Tp3JWaYBa504MV5fuP
yqT88wqnOw5WlkQHTI5Pu70Qx7F31aaQlvRcQqY5NHWlVw7NPAcXT9MUCvvsBc+T
EIPX+hmO8eDaft7hzBuX7bXiLV2TX1vgGRJth+HVBFVtxLi6tN+Eg3XP8l/CmZim
DaXw/zQ94umK0SB467djubwsoMO8cJx8PD4Gdj3fopzFutLLvgrRetMyhnePdQrY
3quH5ZCB07cnsf3fOd8AZdWWhunPqqp/Jh7UW8EdfqsWERh9ZqVG6DRMEUKd/9t3
WO4p2h/1oukIJPgbjXettSh3Uu+xw42AzBeG2l94eo/1qckTgFZbxtceq3RA5R9b
4GZOyEwdXYMrqiEZR5MgJRLy1hSa4NWY26nZVLVm7F0XsN5MdXW5xrd8NzWXLJ+w
6ob+pm8kpgFCHbFF/P5rNo1gW4ebssdqmfpLLDY7ga5lj8M7wQxV2chsF+ILzBbp
iyh26sQHi5pa3xu5C86qLya7Dalh2OPtVTWlziDAD1LhBfVV9JpQ5HiA0/eobTvL
Dx+VzD0tTCaBzP5hm3bqhpUN5LHCNO7Qvsp7dwVIxnalFDHnRb26c+SbFj145jZJ
4sYzC/kgX8qEMHiD4Rt70X4N7YrGiDjh4Cyhj6gn+LwOCGLKFeZLvJxMfS0IEpND
7v0W+uPIkRQ4DTGMR4gnVqEF91KXG1/ijchRxsSRNH717czg8AgnhGDNQy53FD79
x0T6P8g7LjviuA+CdmjztZjBuJjxXG36SOddGTcTWKWlANDRJMTbvpIZiC9F8F8G
/5KuDP9zRIFGgwimYvjC43yERmwdt/hwEbGKZ/LevwGSKSKnc3jGe5R+polPzBOs
xWBBX1FgPrT0A66Uzg8rR25OdjkHxW8OfsQSRQz845R56I/tCcBNYUfTNtEHt4+s
AY1j2uip0vDHAuxuhLKz0jBv/IgPOSdWFmTBtUBcoiw0BT2PqHbhriVEjajf6VVs
BJAYhLKM2bvbqSU60nQzaZmqAB/Xed+wYvtcy6O6/ovyW1kiy7n9ir7G/TpUKYdW
9/eor8NrFFDRZYrUb7PKye8UMgm7L8NwSWvIEFHd/TD5hTHffowuhR14v3vCP33Q
6An4B+XDKiaAo5irE/3gzMPadrqJlgFap2z55Ff/djGyf0ZpX+ap50C9QiDIcX13
fqcZ42JYAtMhuBNFroBpA0RVnJRW5MOE+qNBGW7u3UOMNYL4iYVsI0zyC3w+PJO2
4JfJ+3JuCaFVIGXb+DSOldZPE8rKenAGj2+QRUs/v2bGiKcoI8JA5+d272H5BP89
Q2SZHC/Q0b+IAlegJ4r+XRsCl3dfCDH0usw7maIEbLesgn5TBaHgcWTOQQ+89ej2
sb2ARDO3kwg2q+4Z+CBwt6cmsGxZgjQWecbHyN6bBzfPPzp26ltFblv2WxHYTJ/p
U7WWkL3nBgGH7OhFBKJqyHa0zTvA5nA43fStpziI5VWToOVhvGHbY3e+RdrsCVrJ
Q+0TErpTW7FsNs4yTrG+Xq8ktA5ztzOpVYrM6Mgz/K+b2rqxVUq+oA2cMFnSbF1O
vbLl2bjlB77hUvEK7AJyxU2xAOCT7LHrlJgkMPm+xBLc5DvpPjZA/gnl0dcF5cBw
Sw3+0nqXYc9ekr8Ti9xPBJHesytgJ93mBNnR4+3Zw1MjpinMU3fz6y4HCN6U6lKr
3kvrAgbZWD2VroyGI9BKXlTzZRc6B8o1IskPNSg9pF578EVl3eODSkGUbIVE/UvC
dyyJl923XNDbJ8xqXNZu/E4j3ptBBvzS0INwRj4dSkq5NXKxzO6EzM5bgNo3Q4ei
Haxk6jU2qD1ruvXNrN81r/yjLUyhfwQqYF45hcy9zf5nlvo5svufRPmTYn9VqYvh
MjV9cSPWvYrVsfmfhVaz/suE6NgdkX/pjxQ+3MmDQvYwlDOtUUsuwYvWnJe7ZHIU
YQW0hO4P3LZaLG341qfyr7Xxn+aMith3owbn/Yw1X1rwY+TuznEWHGhITjoz7yXx
+bOjTNl68bWAErVxG0tb+FSjcCkkPF/0I1ACKVEgCmWOdZBeeQShs2rc/L0ybMEf
uM1aCW/+tYXUttGVVCbMLfsY8emP0vpr/NABhSlJNJb6s4lF9v8nyMJyE2YmcFJl
qgMjO2w38m61Jg5L4GaaTc0EVv8o1iz5VExiXajgbYwZJzgOXq++Tl8tbA0tuynA
lpMBXX9VsS/0eFqqn8a8EmUnOAyI+mm29A503hmHvqSjySC6tt7V5q8U9SZTLdKe
cB7BmbQ3wkmMMZvdImDhdZQJZeaWlCj6xLTxitiBZ635l/jcYQ50J9fz79Rw8Mfl
XlR1lqjMuD+xMx4KIDRD+tsdnpaWNJDwxxY8wE1Di+76oXgIyrcCxlO5Djhs72wz
yPImPbxeM++2St+kmjjqZ2vnV/bv/kFIKoRZpgnmQLSr7PLiOWYb3bnPjB0fGjuU
CYUnKS2+LSPYx9CQjIPmArhW6X8IruExPK1QQe9rrS6Os/gysgdgJCDMYcQJ0jN+
1St9PRdrlkDaV+l9UWWm56ByUQgkq9zXkpHr4xVNEDMoPbcbultDH0PC+cFRNtlw
a4vp3QA+12AeSEqbVyrHUvjxcSRoBBPrbDEq/d7IvO3C+mQPDQ0B0vdQa6632lkF
kUojyq4AbnAw9/0qcrzU1XjSBzqiunOuxQESrfR84YfQQbK6JZwlB0MaS5Q38etQ
j7IMvexBWGuqIjxzeqfwT/bqk7cUG7hVyAjzjUV7eSFK5w6dbN07dteeL/p7RyVC
A/cuI8DnpV+yO7YXvGMKIyw8BCSKtnWACyCNY+joTwssByhQAof2CyqeQS6KSC9v
G5vLXJup2+WB5SMNooR+zdIz7hsAmrSuRUJMjX7ebAM9RTasZRrsZLR04fFivCcS
3GlvGsrA5a7lW8z4Rg3Zw7jUaFwoKV9hXZnJocWmpRFUcRoozL59OkJaG9ESzUlv
4CzBGmqNQPZIq2vWCEdg4ufTM88Z3E8MxW5/VnmRrlhnYYcLgoJjndVnxwrhAxyr
qrRGcZJDB7sV8IWczIIDCK4W4Xl3semqaEKNR3BBLafebBEd5RyAwc5DyIKfhMVB
YCFsiLFbcDJpT85Uy2kfRHFkQFk3XuOF1hADBY/To+AJMaOGkyG/QqLqdm2AMHDY
HVrF2yYTvbDf6M/YtRB6T6y2HMiFtuATpdKSqAB5I7Tl93F/+ZtBncrejLkYP0CG
z2wf5nSKwRj+cwXAszwWAXzoQY4IYGTqA1+wQLffFLyK5qICrUbWOPxSOHfpFkjF
d3AhjLzjc0iCgok35lnq9pOYLpE44hV86FDnQVy2u1lykCGns1niZmouumyediQo
Tjzinin+E9DD6/ZFDvKsAZRwMkpBfk4H+ExSYWDmylHqTqxZy9aXn2PF8O8Gh6Au
lXnZQChQ3BtALNuj+mfy5mKReigKAWn1LrXtYiuXu4Ob5g0lCHzJkiOHwbHgVcRH
jAITgEWWrx1QMEIEUE6+XoAA6mYpz5qlpEzL9PnlRHE0aY9EvXvTvB1zbl7sIcrw
rbek7tGfAD5XhpIUZx3icoIPfkje1SfOrWnJIcWzjm424q6dh6ELlUHPmhG74jRG
l9uoqVGboeW0zFNxJJh8qwGk5xlXItmjh4l5kq4g7+quORHLu3feutSkHNCTwI5x
v1IuqKARFrW6YUnCV0RLd8+pr8KXdqOxHZTJu7EIDXB2aINL5R8c/sJ2QgnQBM52
OlExOowtPeu9Zslf8zjUW8nSgBOQsQxbWkapwFo0/c7J7xmWjgGkVEqjIZzOe3Qb
SuZqQvOuhINqiwy2VEKX5eFdikRTqY3KTOORlY+Y9COX6BSC0NBQ95bz6/EljOxK
9u7i4fg4+3VtngCTstw1LDTwuNniiTNnVL310EPAeA4rmjSRWy5sUYZkUdY5mUoa
sxboeR+5Ajw/JAZUz7pfVy9xt7dTx0zexpdHWOJsxLYaszcQ4xY8GAcY7vQF8uqe
aPC2Tkveb3Oe4B4NK82H/dJuIFT02tCeriMZ7a6nNO1/WVUl7UhUcvTG5IMSID5+
0EGUkmFc+GzWi3pFHBGEQrsU4sEMd3Aza89IzyrqF4USqI1q9RUXR3AnKC6pi93d
6/sMIO6MnWSpa/wFazNKysisencxk1z5ZeytMqOHesPk06BHcXzaNCFJwdvtG4dQ
fqIE3WOT/IVoOENh6TyMGML3vZTK6Lz+MkiCkFNi2w7nqQ3mpFt6zzg1jgJfO9gP
yuGstaO+SjvwM6xyzThHvXLx9BDldhdYI5LiqPIh+/UtV5tM25m+SSuWtj0CFBZS
QFUcQtqZcNQFPVgqEW2gQ+3j8nr7VDHmhP7uHCVVvG7RuYWqKS8FxI8y+IwTO5kU
9hzW+yd4neZCvJPRan3Uo+flWCtP+VFN3w9/eH1XKX/JNhnZNOXE9q2DlIU4olS1
5gfF3YGT+Jpb6VzoNlZxbI7x39196ZDMOO0KhtFWbgCMxqZtghZ1dUO/BbFE+G39
HN5H8NOWywC+TmiPDPk7Rbw0JSG1jRgoToVb/6wEfSqmlhBbUfhBm3pFCkfcj6vv
/orhxiTQRsMQIznrNBTJa0TpG+iEk55H5aUwt0b9ITwWVWc6eBDQUxOci/Xhzz9V
PEKaTXZPZu/FPkaCa/h3zO4pC4cijVcfvlVNKhcQFo2q4A+4Wx0Oit3DfCzUPaKC
H+eKI5hjQsyC058SNcbk3ZnSZZicvsedwai2mfsvMT9aJSDgzoDCuFwv7lCULeNE
mt46BQ5kOKQiRF4I+ZmFWj0YZ8i/7XxXoUUGt9nWDVbnO9BNEHe91zZQQoGoDJRG
AVl3RyYhYk8MEOoEVLGXPkmEyD33zkqBKR3/Xy8HKNocKPxvQ7CFFqXNBd7h+4LM
5JyiLtCZhH255lgSwWK6KUfMZ3H5KnfBhp8t5RN8JYdFvpWhLOW77ZZJ9HKZaiy4
FLFgEvyU09uqX5uOr33RPG2blCkqdc5UBwoZJSCBsSS1QmxwFjwHtgLsGe5SukMV
2kli7gve500DLDWqJVH02lvPMKgM0gEm1BhQu9bIJ7TjZNt/Uyp+NuQo4gPq8XCX
eobRYSIeZejis9umOc3AgwieTm7jofffk5OUWVSxST2vOoG2lp39d8dF8YiIrsIo
/iet7MNsl5OEuCEwzMjXUsK2Y/UhpDE/LJSTNxYjBVJ1LLVph3x4to/RG2GORFhu
x4iBU59qhfyEHZvf77GBaGw89DFcK3jtagEukUykUEimIyWo2hSd8ULsC1sBmzah
C6vtQbOYDjMMjvqoZiTn2PfPPLade7EKOwuP2k97hQ0bKzQ0APKmqz3vnbmLOmRZ
`protect end_protected