`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
xl+hxsegM9+gPkvRB6CsqaNG93a57NZqZTKN1Rlh5q2g8sqFTyT1K5p+EXZZrbGf
dbSLPs7nYLXbdyf++LWl3Q1uRJ2smdwH2D24PdDwvv+G/2bBB5aPwIRzteLGkOPn
uy22x4ICM8CtgdR2x6fg14W9e132vKqiUmYiVlWBc6Jpj4E+mR9JFlrUo3mbsr8S
k6aXBaSs/wMgs8w83o5rp9w6WQbVLTLHaIrRwPlsPbY7gwUab/CdvKI5tW7Fi29W
FFE5vQ96pc99tyz6u3IxLrgWAvOJbOAnYAJI1++tYNHjDjx3x5rk2qCwVg84GLgv
degBhQJsVU2RYSVAFgDN0+I2Exde95pkiauYhFI8EsOsnSHey5kbS4Sdn6F/h+az
7bygMpnaMcRg3ZRrIkIm+ZKD5YopNd7ptl66jZah5OU0dlZXPDIl3qm3DcHAiRXt
taqRaLkA3Z4TXIjcRTh/dUSTTiqh+8/2uEVxwiRH1i8lgyXjo8p0cN9BRzM3sGdA
bGakU9BIdO1kkst0xOOOZ3QNOsXM6rHXU/dVo6+/wcDxCNxKq6W8xzhgzJiEi/Mf
0o+XeL04yNNkvAW2Zf4Oq2thg5Sd2nqM7I4O2HeswIGBQHNGE++8Aacj5z14vEXM
qUixnKrfigbIpN75HQ690bNsbf+7iIotsE5g7N99y+b3Vz2l+NsTO57KOq0sAcCw
7Xu2gkczjYvj6J4KDRiVoBHoPPi1EllQAJ4Vq6dcRC8vkecSDqO5mChG88/FDURH
6yBNBQtzdIpaP9O1uoZA2VSXZGSxrpye70lS/OUP5ATJfZ1tB73mKtEkOrB3Twi0
nloBhTRoh2OXZdcHaGX9bqr9CAnZ4U6q5Y9fu1tyx4VraiG5HGKneXMupmTWmLBp
8C8C2/qJlxneoLBGJ2N08r2iisXeHZz5bSWN8N99Nuu35Z+Mbhu2smpjVFJ6G9Hg
Ed394w1mU5nHWifP9qfO6toBYGY3sETUmf8lVumNlqxO5QDTfEMBZkeCt4IBTX4h
ztoii6OJlcmOc0zqNCEG7mTiW6SsivpE+DzZYu3d9olWjHY6b4doVk6liAZSSfbd
ll03NVBAFOm5Dq455wMIhRqRh+pGH9IN8RiTV0heOcPmbWiz9L6lCyrt5A0HvwPq
XMAmsVbdcnh4ZUfJg1zTuE74RixjObSBA0oXA+cjQzx+ER0ZPR7hOjGIqFEHXslh
HlpwMM6Z6Pns0UgrCYWhXn0O+i8vxsfhJiE0vgVii3a4sJYFOFCTdJD9qUhboQF5
cjNufwdbvlXvjRyvCOspc1dJSKTIsCKD+NM5pxSmev2mD8tbOlY691ceC0ntvF+f
6MWVq2//VczyyqFmdNPioJVtZD4S7Xkz+NcV9Wx+Sg87P0cH+pnbKOegOT5ulL/e
7Lee3Cg2fvcczBw7LpjlsIju43tHGMya3ZEsnzct5B+tJlVMAj7J5hWiR2gDW+Oo
p5CyOf91+tuK7+UVR+l6ZvKBwsxoI4G5KlpSxwFr8DYNBZoZs01wqqEHDX3jy5U2
y3Eusxs2fQB46r2Fz2RmvBSJj+NRVZkfz/wKyIuiNEgvYr8V8AxjjTlUWpJkAvjb
1K9eRzPRXeo7pPVYE5GF+WA9qTRzlDHv9K0UbvRs1VFLzciLZDss1/bKuXrgFsyL
MZc28m35zWJu4WMofEvhnKrX1C0eTyGP/OmjS9R6QSaaLkv4REbL5FJJm8nkFxcD
sji739AE133KcfPDt/sKIZGqmaDfOSPXAHxk1BtoaavXtUAGXB2jfm4Q+kQssq4M
V/LfZw2VVZa1OGSmgZcn7kj6A9EAll9b872pK9p3+pE6CSMA9NokyQ+XIv+I9rc0
vVqn1Nmvs566CJs918LZFaPOnaXOmGaJmANU9EDiAdHeHpKa4N3gz/QNj9tohjLN
J7tm3x9VEnE6xdrrFXUvGH8e8+kB9f+rYCMmkr/odeGSY4x07Pq1jrGvBepUMEV8
sGA0821hWWiWzG/cU3cGYoMr5hKIoNrGWH8y7XsQVR34bCXHvTCnFgnonzR5ohcn
XTBtXjl76cekLhcKDVn86zSUKZXskBRqVaxEDv4YgR0Bsf/tL6vK/KtV15awKR0G
/PAQaGfxYTICvgmFtVIOju1l0HRRIpUPJYLSTOyLysAV7uD6WiJ6HeSx4aIYQWqr
57kBi8qAvFmjhenldsH9Q827/79tTwj2nNGAlaIeNmNXzBLQWKtKP3Bl90e/ZhRj
yFkMdNOkiz1yfPPGHjYrwSHc4YVqz83xGLw9I9Vv+C0TXWMNUbpuyAExnNvnmcFu
ymGd8h3aPAQcWvzt2d1LsV3m1LnHV0y2UxrijEEkxGxzz3D6t/5UbZCWtMHLRUh8
gOhv17aRKQPnhnOZpxhlsja06Y8KTroq6ICkVRXErbKWd+GdAc7MEjPi0MlSclkk
tQnDizYk+/Am6BJCiXQ0kccGZbEjTwuHhqPLgBSbcAS/rnh2L9f5jmDTBf6qJreH
xqn+LMCCpCkGKCQFelzlgmnoANzwYXJ7bWHrFKnsZEvtp/iHMWpLgz3LYiIuzFPc
`protect end_protected