`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9056 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
YKazAXTwZvVeXonKKI9l+8U9Shdem0a/bKmHlnYg5N40aHEtRSzFUg51UDmTufd0
m8dPFVBHDvWWeReM4T/h9bplONEI5W9V1UwTbshKTl/ky+WuSrPnxmfEw4mVbit8
cUThP4ZP+wJskfWvSsZun0Ttw/ItKy8p11Qf9UpllxaH15N3SBVuCG23KJ0C6IoG
pUqaW77r2VnsTJBKOUl9YpI6aU7dnD1MZbLE3015JTY1oKhaUTllmj3KIg3ZkWif
BNnquD/WCGoCaBPcLBnrOsdk1pb3YiYM3qL9U+s4CQIiKXTbarcJVRVpsj8oGdFx
9bV1+3qchrg5XVZHc3sr42pnapbi9JF6aYFFmK97mwkhB9ZsS2/PxDDyDzZNbHIg
fMCQe14E48NB2NqKHNsQb5ZANbkdh13T7NZm3VYsb7T1r2pR9BXubdrH/rmxogyl
N6BccpMpGMk1dJH6cKN1Q5N7PZ8M4uTRVOUBT8CiPsHQKW0majESlNOqprHOP6Mo
NSOdHK9mmaHqUmL7/8iGdeV1V63ZM99o2Nuqr83NXCUQjLggoFeeNErMBhD9fUDD
6r/6rkREZ0GYx5GhtsfHyxahnhBEdk48dBYXE8dnj8rY/rk1lQ6SDpZf9bPnZX5f
/XWGCICrIG2oGywvjjc9MI5VktjH8K8Cu77dbpBHHJKilQV49V8ugxVm4M4CEhEB
/ORNUyxDoWqOO7kxyWHWodzF4WoK8IvUxwxxJihbD+t2mqxppm6lh5zsWSXXTOCk
YnAUXNhsNvbalMI4nzrMaeQAdqkmgDhleJEX4wQ24BGErbnvfv+Px1s2dbFC1dmx
UB0bU3eVLLJ6gE9AxyS7HXLOWjAMkrbcaiTl/FpQjblANfoSy/ciVNR6ZbZDW2By
7YZOVTZhnt9fjYtJpNQ8pbeUKTvFxtlFEP9lG3mc07nxCytjvpVdr+uws2jaXrum
EqhpsHZ6bzorAfjXNCpYgkhLMk3XxRCdJZRA/EvIQqWfNAyPRTq2OXaOewl/9d+B
SGmBcw8W4MRzA16B8KsgbL19XdXM1Cf5r1BBf4xoB92xk6JD0FTjo8kWdHYg9oGW
HQFv7QIlnUYAXFNr3tRN4M/11JFngU0ZZ2aGKllfVmD7JDPROJHrLowktHicccLY
kOQhJ9+IIcWjMxoHcWPiwkdbYzhi8v5Da7+kWQifaeZm3CtYK00ZEDlEFV0VzsLT
cNs0Vbrktf4SwpkJDPWK6ESmK4STTkXR9PmlzM4k0dCyUj9vnDlEwF6TT9rdLncF
RAoDf/JqHh4/W5Bipw77CxVq2Skxo3/V8Y5ubWsPVIbkpsfcGwKUbnVpBRUGGwx/
TrQXUK8qWy1dO+YILxJ66cyuVkPyohmpP4hFHmhZ2Q6w9/UR8UDp9S1w5o4gDD/W
2QxPGWsfKwjqIt2IG/e5PI8gTt/hyodb6gIZKKvmnV4IDK+iR8UviEGBI7GxAwP8
D7ISz0ByNYo8XqaVY4UP8QVw9YL1FqJBtTJrwN9DNrK3GBeIqFdL9lQRbkbqnDCl
6IXLfgEQqNMluh11t0+oKDyw2uci2Y7boojIJFbxEsyfXyo53FkqleBFwvNwssKT
nKeoaJXXJYTJyvJf5eAZrJQoyTcM0VNMtUhxoO0bLzS9JnRmTV5XQ6PtDbTnEs/c
yZ0o6nYRe/Lca2c3JIoK9Jfu4YYekI+X3VYQlBal0VuyB/qwffV0ZlygVROJhYMo
mbiUWExEClvO62RXQuBr22YvK707PND5DeRrHTFmTZL85hmncJGrwu/I4npfYBbB
wjOazcN5PN2Iarm7gS12vmb+MJQ/73iwbOotR9Y8c7MJGucnmBMV4lhj4jmYkW0j
y423VJL+I9vKbDZmyJeM2Do5oy0hevG+vjx7TozIpkxaT4yYYptlD5p9VPVs9dY1
NQM28Zen5Ykhub9370ciBbpQ8E7nInmAyCnw561lyFYTRPbGUZnI46NN/dEQCWcC
Rtc7+nclzrY4atYWXapianXiC2QqLOYXJSa9kUyjq1ex+Eg2kKjdmue5eGa7aum6
DFo8wMfCbHAGc1g67wK2B+2QNIW9xYPGUuQgmdhOGKv+CJ4rArdL90I/pT05CrRG
VkhzjOhxRKFGQx3Lfpri4fl6dRjxZ6Gsgl0Xce6PpIMPFHxUgNJOu6zkP3J0B05B
t7ZzpaVyAZwereXKwXsuTflJojr8BRr0VzXUGZHIUJLoswfMCde9hWA1CcvApxBI
LdFN6GQKnV1RxcdDqLldgf5gEhlZTxGwnCJN3K68AuEKr5CEHY3miYmV4NoKjH90
FclPnsB9vLZq0yUF0bV2iZrY5aSSNfZKC/Ea3NKtgs5I4Wefp8ddf79UcOV6Qrn8
qULXk4jmSVfXcRHHcmPfnUEpyfYjN83JSrNZ4Xr0uyocRFr9d2Zk7Q2Z4PIlrYZf
IhhOQPCGXHNCerN+nzBTMGurhD6sVAoQ0UuAlQ9XER70NROgpomaDMRKPkU6wUqS
htWLFe1gDXMMKD3n0bIYDExMxRrSMgOFr8u4VK49oQvThxw0WaYHgPh2rzXbTxFf
dYdlhb8jRqyPjt7Gqs1gVcg+RWM3S8xGhG04d6POSzKymKyWcxg8asXpVO4ptxgw
uTO3/57PMtQ9DgDi5L7EKCMV8SZ+mURR4y1Mc02ybNZ5ZV8ZzoOIO9QX0ZfrGgxe
wSrDOyySwa4iJbDJfthcc4tIMYRR3O3AYI2wJDWfZTgv6XtwZzIOjRicw1qFe1yC
Js2ir8xoj9lqualUg05B9Wa6JfxCnBZoK0Aokj2xQ5J89+CQx3BIcuqXKWHx7X9g
yziF76hmAhA6n9AVytHP9eQRItk8WEbXv4D0tQ/ZpAShYlifiFqL6lWB+R/UlUsL
N+oZN12Ek5jkbn1dNHfLH9HyYVPN31hFSV2PEvUvCRvjqXR+nDiIIsjY4zjYLzF/
ie4FQ5I5/2nPu0gwKAgJRs9cVkZeUsk9pmse0w/ika5GaBVB4UFA9dyHzwPzzDp3
2nIdsZMTOv8q1uaaM/Lll1qmDeN9+CJAw/+E/ikKUacm9tFqPzTnLsRuJv1s3OQm
GgW97uC9VGHpAhhSfUKR5UOrGEEvl43elq2TGiylDkVB5n4PtkX/D1ucM1bZiAKN
4KUsKe6h1VjClj+2Qt2r3HkxH9kOUoXZ/07shFmZcVCtDaF2yCANqIT3qEpAzxEL
brLTrnVz4myku3Fj4tc/c1SzpM08sjHITXUW6+e1pa2O1FRncT1i2jyxwBVo0ChP
2dyS/689kzzcdPqoZaZKWUWWBQ8I6CyqSEruW+NfaAvnejjk1BSd+USf/fJJivk2
jhdvZMdrCL82kSKfkLeGcJzRDqruH/mjVFwM4Siz/XbqhAo0oPTE/rF2mcftrfOL
yMLjDW3LXoApWh7hHp9dZinSVefLf1V7/1kz2GsqJhoHzF1VFw1014jjpJigEazD
VAdG79cYQVsDh+VXJUsOEe+4YXQ0ugkgouXaN9YS/fXLNqVCD0yynABAuYcKsVD0
qHD67ZrJZ/3o3MluRIg0F3vvdsRkcQtF/3W/4Tc6yNPdKoWe/R23gfp1vCMLo4WH
NN0iccOec2b0Z0+im6ATrNNSbhB8qjuj6Uld1WWJL9lhbhDavQvly9/gKmjhSrRn
TSsY9tOuxJW/a0n3CsMrwJnS+2QYCPxhZKuYytoP9ZkeIGKrcPwtNJm418RUPfrl
woKGtIG20iFPYle15LPFirG1TSu5RyMjaiLyq7LwK3VtG2fbTyzbHBkvhvh0m3SJ
LnIYddfh/OTie1MXjgcIowGCicWeMNB13WH5m3hqqeNreWml6DbReRd/7CmAklYc
jNpxOmdho7kI/n1j4XVu+6diUWt6h7GyHxKmLizoPUBNCPkQ3AzzUsYRUu8lvbNa
GDmqDJXjZ3EOlA5dwKqnqJxKIpl3Ho3G04EVeogDGv8rpWIWUnFJRk3tbdrp8Ft7
PuwhIAx+aO3Bfn54Bdgsuayt8uFW9Ks8RtKK1wk/4EE083lSy31HExvwJYYYjIvE
tEVIIfIRYagr99YRNoA7pSlgFox/yB0ROLCvMrn7j4676n6dt8gc+GXpPd/Yd+pE
qWjWCBEjvOw3Umottt1B6vxhmc0MmWwF2jVwGuPX1zwePYDfBqAbExlCIytNhY38
4x6eLg03LLyYY5r9WM/9uyKfHuAFYQ0VapJOJ+/vxRZBEuDJeOP7IGpCTBo4gml+
K6CRaxvDWLHtcn7kP5v/Aeh6fbJ0xLfPTfemWOcNGxfduocAzvJ90hzuz1VOTHtK
THNH7fSj6NG26c84TQeBuNVm1symcoeLRO7J5VqKS3FEvSWM3qQe1K0n+Kzfxutf
z38GjmfUcekSoOO2zR5BbGUx4NKeDcqLAP5QBXwctxdR0r3XYkhRhoOE11FVnwxb
kUfFeCNS3i5QhNsLJ+rm/Ay0RRO77L8Fljln11rVoGFNGW+aGNVoySVkQ9YEWik0
GvufQGKUGyFZzg/Dh8nTvX59XVXsXJ3UHz26WSBSieBB3Yrzh8ZFHll2gt3Rm2J7
UtA78tPHmga+d4C2iMWr63SJC3jWtaY3zvlpHDUxKcZNeohJfCcQ18fPulu2/+mj
ySiZJAxWn/aBKCI2HnKY7BLvjZMO1U3ISSy16mYXysMvklW6Cwl8IelB/YxuXB4c
VGrXwZPTRr3dkfimXc3IM2fhq+sAHIrHFEi8hjG7BCEFoetiqdtwwFJdNeTo/Gvb
KqxjeunvHnj90zkWCcEPV7i3QChJxD/11cDfrAurYtnj5TRsK7fk6hE42r2L0Cnr
yFDhDGS1AzaT7Yc97x1u6plVLtbPkkdPJTHytlO2lnntt87/6OtCINYz9OU+9rj4
57nu2yDJarz9RpWPNED1CAtHanaKfZ46Y6u9iwmbULRtfZCMujZWYBuuqqzwn3gR
H7wje4exbwO2Mf/NJHnJlM5JRtNAFqtE03YaLdvB8mNGWjnF1YO/F2d8r3eyXbE1
xWQQLPE1sJL3Af6/7i4szkDhDsCDao0atz/+J2gihJlpbwr78xug6PGuO6E2Twyw
6YhQa4CZUCSaMd4dLxRAwTJjkQsNBsitheLjldg2V6w3Z0wlvDq5J5qMjypPdEVx
CFz9Tu8IHrvlUauXpdvKRJAH4XM1i6PCjXxZIMJeHVOV1G66zI1/SifoLM86Tiae
n/JAzx1Ab/Zb8iBnIUHixG+s5SVinyNUb6SSumRtYzRP7RnH//ZGDHH2ATu3j9//
gfc0W3BvcxaBuYJNd8657PD+chhz1tZ8+tWCaMg7+IfsXhSUBv4Vb9HDqkNnKH6T
7R0/mdk7oKZR3kTnZaSh83bAcFk0/FZeGjpdWoRnXPFHT78vIuI9ARRjve+9Jvok
/WHjGss2QF+jT1c2pSLNA/kEah760Fjgn7rJwD5rueFUSSXpp7aqWAN3xVkX87v4
s9YTKxOn3OfEfnAB7OrqD7qyEclVXOJb76ycjVDULuLLk8rN2EmH0xjpavYpi77y
ZB11L1uAufCXuZhoSQ9HwfAjXFGsOl+ko8lwSUN4o+XwOJ2CoPtRNcO0L5Qkrgek
VPgZ+d46DJug0T3EamepNoozVgyhdj+3h6HBJ9ZnTp9gvoPBO3RPkfw8TBPQJSyL
P7ebtMcBet/pP0RQ+VF3RLLuaeDSnoUyBjb2Qu54dUYB8dVzKmJR4ySfrgOX/5X2
O/9Xc+uOQjnBIXqowsosrJ/8YqRjpYdeqSnLu7RNq+aRWGlmenau2z3FVmr7VjeL
AWELSRQAodIRcWnGGe/c4Ebf81oAiwIJxPDD56NhH5a2gTEEskY4tq4lcezIqv1a
Nw2PZhaoYTNLfNOA1elHx8hhts1+htCXFTPXCdrPG0+CCMaEnM+MHWhpLx711LHg
NS0vana3l2QKHg5bepks4tQa0nL1hvLYHxI1ecsO8QgoD0WQA6zcLcyCQ7SDoaQa
mkZG0vrF/Upq9/SMlIjIdcL9ZB9KArOTlww9mBWVvBWbTVqiF2OnjGyxnKQSu9Kr
Xcxhpctf9W4XFRTGaLZ0uAjtfF+e2LZefFKLN9hSCyTtTZ8w2Mo3/ZzuRRC1z0nZ
o78mz3X8mjU3PlZKUN4HDkOsXfVML3dgHdX8TTIp1Y3MwGFsSZVO5ighh6tRM5Yx
ApnlOJtXUGAWMM86jB+QncZKQJxs/EJN2SyJ9m9108/kdKSw9PkvHzEbTDFvrGQ2
8z/0rMnoDTNiztntqdCQr2QM7MTFOGDQl9WiiEtWI8u98lJcwQs+WRiGSrrpxyoo
rcyEodaKNYZPDm6jR7+2yGOtWn9Pi3UvxX9a7hytoecAW7vChzqbkMB562ayFi6I
IJNUST9IPiuuXI7f7WpXQ/yFknb965BJrOTbqKbCknstPqqXyXQaKt5Vvj7icPW/
yjO+7i1K7UiWWsVxBXWt9jetW1jeBjWo8R/HhYaSlMCY/1vPFt6IKQQOu52lLH8T
lJavUowOvfs4Fa8Hb77xERRmiLxj0uUYYFHjKKyweAm/rD6yTS9n/tlwDVtJmgx4
tylAb/u0u1QiMCPp/VcOifE6LHaf77rftejY/AJyK1MkExE55YtKbduJ5y9xGVY7
rJKE6loGgkkvDJjMjFkfcNFTLXQnxDuibzAVgrH1B33wdWmKFTR9fsDNhmHrdO2Q
UDx2YkK/ybWgiPkY1SssGdsrjSmzGKzVdHPDuToSIiI+v/fciP9aK4UG7tC3c6y8
l1vUO8O6/UDlYmOLRu7wwGIGaxPC7Njjww74NwqXX/vsMsBUNUr7i5xlDQ5dHNwx
IWWgn/VP03x3MRHGFoWDHT/Ko2QXMbIR7xpk+fkGOqe322FHM/5M1o8LPeQ8b/FU
FlNIPSGrjmgrKqUoqgMGfsiBNa2+zFNN1z1mBBQdLeSFmJKiBxxhUZ5wsoXbRaK9
l1QaSacBgUFDaUNly64mmkSX+7loOYKCVHkwn1FXJ6eVmQnu/wpXtBNTj2IbLSw8
bCCufaaULbVppus1K7pIT6G0kMteq+FbZ6EmwA7Ed4zO5UjYrNDHOLho8ClE3y/7
lsy7rRruOt7HG92AB/kAj8iTQQ9Mhq61ivh1f42Ai+KG7e1W3v6RU41ettXGZMOC
KPf+rU8kXL+Ja+OTS+/AUJAm5uiVWpFTDJ4T8vmk3SUjuwavbUiT3MfriUdZeues
yic2bpPXEM8qGiq3aPD3ez8J93VYiU/UcW0JTppkG633bwy7s+ZjCF/CBb0vACOz
Znj/AiO5iEobdNG3KrIgLojJIO/53QbvKCoUSRVHXpR6FjymwI/tp65qr421FC1W
Pm+P6BPegqZncEohshfeYxjKube+Rb8paIlms5Fbn2UE5VcS6mL4Fd7nzrmGaQpS
F+XjATsiLICUZbT6JOrWzUGV/gVJU+jlwT6eR5WmQY9OaJwRh+Jf74VeqYisvfxG
8550LYMzu3upMFrj++MXG7kD8V/cCeQ4PCzkbST2OGWhxhihmkU9CzvHW3yzsdDr
ZKLpXKKlAmBK+zDw8/mvv+mkFh9ElgeBe9FLoC5OHjeLJSonZNZxxS8/FEkV5T94
/kEcwET4asOxAqeX5lbAqjITB+S81Mb7QM55sMjrn2dbhfKCLMzadqufsbJEKILy
fputtg56oCijeUI3eLqBLaj35YlBCWgvqfJ0MgOcKercY/Ks1k2Fm9L11bNueZgt
5pFt0RNMFQFOsABDQwj/IJ00jB+TMVgVE2bDbYJdPfqZB3u9maLSHXM3JkKDxNEj
ea4afVgBjX/Wq16m1sIAFci6S88EMhwI01AW4DO41GJD8j7hF+F8hOvBsPOZaoU1
KVlG7RIqxLOso9R16A1W+zXhUfTur6VlbHceDr2E7yWjIvZ6eAZ33e+0QNKjI5C1
hLsYfr1QGV9ld7XZISV97jUxqZRqvi3aBmq+W6ySIg8Y2S9snLL4f1n7QmZJU3lO
8oLASG8GWJQGbibEQZXr8d5tE7LULKktaQXWuiZ+gl8N0NrTxgCqs608ZvamLLcE
O6Yyl9G6+BhuUkvK9+E68fDd+V/gAaSCBYVZ0GVgqqZ9vu+o9xdNMVV1N6Ph510b
4ltaCe08ZwXc16pww/lE9MH5MCFp8HnNOQ1uekXPVQdqGOv6g+yBJs1dWJdllk/+
AhuusYz2Y/RGr4TH4/bG5US+Itv8fhSlH5drhetuV3kj8PG89vcbnCdFFuX+wvtT
PzGmNlpLDbUo0gIUy16ISKvPrVgZEI4zeIfRKZIYQAjajnw32YKY29SDZhoDaeWA
NfcyR9x+7kWVm3CBRY77/mKIVyfHfR4zPCC1x7SXN9/p7g3Z00bZpWe7oKBFwhUm
SmhqCXbNoS7EbRfCguwltDCn3uGQfyiRM3p65dEPGATXY9ZY1p047DzQ/1iGyQhG
qCBRjGOzPzmlB2GiUo83T5He8HClfNTrW7c0qPvLpaPMoJ3UzkuOe5Nduq+Rbd0u
xNnAKFdlTiVv+zeF490CX2ejT1Cxe+hqXWh0e0Iup48WMPn68F2YY31nmHjWJeCx
PsYX9zVicndfyt9m1nrNnjBAqBkapeT4FwXxzCo2jXM3DRq30bVGt3Stu9k0J5XM
Uh1qAmquaE7Kl0WhX0qoz45rCJg3Y7uFooJVN+tFTItcjwNjFnXgxONqCJiAXoC1
GHLC8Pn+mv2CSm/PdE4noTtOzEtS+pJFsynukU/7vzTDiCM15LRNCBnon5nnlCgS
j8YOSmQqOKaV0cY2sc3vka/25tpNiX2ZXlqEcCtGcJ1vBJW7qhpk2WPi8a51NKzh
nxQcR9q4p3DJB6qHhiJk+YBfW3OmvlN7zlFog/Z6qbv+AA7VxuyZw1TC/Q0s8Ltl
U/UyXpx2GVdTbPoxDUqDx2CH2wWMqPb6MjuD7UJveyUze2p7CtqRf/WSYE/in8bF
GZM0lM+4T1MekAfsnPvLbvZYIn0ss0dhg7Z7Udk8rtDmaNNct6XdPiUB7N8pfhGr
t+I0jUZV0xo4p8eSB8lju2mDR0XWIXbcG/Chxr4z7N6qGlEEhTMBK2pNW+jpnfMU
VhuRLadw24SxZ2lV/xk788xQewDEwTY3u65s/bXwdvAeLpoww5DV0KXPCAyuG7Ob
4NNe4Vq0wYaJqNKf72yV90kkoOI1OT/f4QeyQImGlc7Awny61R+Bn+zbKYYKyd4P
Gol9E2Bz5w4RGBvfcd45OE2UU1POzy+WAF635sOpvPuFV0bZafLvODJy1N5Jlvjj
fan047URMr9x+t9SM2BViINYy01sZL5PLB/3G0GF4/8JrVMobcZFqgoOgoIQvdtA
BJ5ySncCihAeNIFtaTKb9OrAvNe7rIMDrCf5C+AzESRY7xT7pdaBN7mm2c/SGL+f
teQppbCn1DXm1wVzjWsJI0iobub9EKTvP7r4xfQoS2yRU4I7d8GjRzC5m0zq5l0E
SPxQD3LFA+fhu0H2IbhMyQb/OGlFeQW7+ijHBqI78frE2RZug/p4naU2pSeZ2TuS
LxnyeVGTXze9L7qyeQ+NPpr1NwgEjzeqECvI59By/3osDjVU+abT6ywZFc4bUPHY
q1FWJ6/sKZPfzN/RioX+gFJtDeUu7+pa5UkGqjGW6EbNwTmFP78I5+xjZzpV9yJR
6AgLVP1oZxI01a3CXdFpcp9h3O70hktcGd+QqfnqHa09h6MG2cUTsVVFW7ecxMBt
RFB12pImnFEfjpWXsEuiYZCHp/GQZFCWv8ylwnEV/MSzfaQg1wZzNUE1upQpX4/R
ZuvI4BJhoJHv35p+vc8eiOqKcQPn8sbVI3nJ7KB2BlugUWijYxqUrYQGL64bCHWz
mEn29r8v/CRHRNLm4Ee4tfcZ8N1PkDVkn5ueDjQRBx3e2WupBffNN6tU+NnLYkuW
kq3+efWXBKOfRZ+l4XLQ5uOClrCpnanzRTZB3BP96TnfUa9IiDAyNfQSMq+pmGpD
BTK6GTF8LfjYeV5LmMiehd0utQC+RKNSv6vtMadX9F2+iC4lTR9l+H7CRJLFsW8m
KBHn1uj3MAQF4fA6v4u85Vyj6cKgItpX1MkVZGDHW93rFGToBj/xB4ZR+xfIxRYW
HF3FCkivTgz9bh+/uqIdhyLzG264c6+x8g7b85TMW4NXh1worKujLxgCA2Ww/PmS
UNMGGRePLDYgbaL8DSkVyVMVX1Tc4Xdoe1NbxxTw9eGAC/1U95dN0OO3bC8gMNqs
lvdFigRhnuI/fVBtw020MN8Y2laG7LtZZQdXhy8r2i/oJiis6Fg1zWqrz/i7tFyZ
c2KZkSb5RSxRuSCj4EtNqfBvW7oa10hiN8xj7WUR/nrVI5VFCoA6hjD+P9n1qzPP
mAWSP53Cpjf0RGNT5c0vI+bTcbpa1EBMG+k/9gORHPfTo+AyhKcFT8e17LxSoc/n
8a+TYiGWBOPl6FAFJcOBp7an2x2ED6ME8ghluln7mnMY6EuNcizv9FeWRg5LLFnc
gHXGfQax3m1W2qiZ94n06covA7HV/+1g1OHtbWBn1+BqzRmmghrv1PjzwUzCRnUP
5fYnPgW7W+5GXQj3tfAbuxL1tDBPPToQXiAWWMsVHvJGX4VuEuRTvuAkv4QPC56U
FV8hTTPm7K+GN2nHkk+rnnlzmoevqZDVdNBSDWhurbiXREypuu58AePvaaW4okl9
jkQ2fsk9hA0SML3YaxpH3E+KFMO3foJ6g1R3QgYzYMfVzz26wkH8aJWB+wph4G/E
sJH6TFK70H2mBSCweZsI3UiekvVIW03q+ilAQk5EF4ZMLKYmOu/Qp1LjdkDPCE8U
CBD8ck/H+W8DhVZTgVnB8f+x517oY4cvMcWZfjrL9O5WnE3AH6QQpWmBGLOfSAHp
BxHcIhDd3Dk4IU2Alqg6cCYbIr+/8Xv78AhdaMXIwXJWsk/d8bF628MXvJT+LV0F
U8zwysHExiUsTRelCBpqQwbRyKn+nhYlLsEzfEMNYvAxzlwANAupgqZfMEhtMLUF
xG1nGQ4z71snodtZSKVyyWvq96NjjnUdAcOCvyck9FvMFxQAyj9FmJDCgC952vR2
5d95n7Gul2YQCb7VelG7NW83YO5npTxIS/oK1tnVj7PqrDhi3rwow8QECztHGzZZ
5hoQNfLTWTdn8rkVZToC6RHTLlunQQXXK1XoG6CkB+jvnfBmgW+BnPSGK5d0MBHq
mTTc8gHIwKY6HZG7pL37GEbrWmd30MqICfkeYWdoS3rj2DvXj8FClePrmAZJvbj1
tqXwVNp+EWLlWcLugo+CL3LStFzYaQaOKrGndqxDG9/22JorT/1q7e5e7C3fHcHQ
71QADqQ2aeHU8gBNsFyMa1p0QqajSTfjgysmOafFRY553Dttgauywc0jp/CQToV8
8vATL6KBRSr7zOtzYObx5JMnCgZqMWiHKEHr8aDOQmycaRYcd5EiAI49DirYbFmS
58IEpqSgjGdx5j2fEIqYzakmeCmrRv+KyCgAl51ZMpiN44vJKHl9tIRfxPDbwrQT
haFFTWEmWqZqIjCtMhiw9fXwfEDQujkJjZ9twAZaV3tXfx9ytiK5CV07hS9c61UE
4l2ujKqLq93nUENjFXsuzgfKa0hwxGe0eBu7Iru2EmDBYOpnnIxb82RDByfLhdts
i4NN9jXa9WKYeesttYFt3yFGnBSLLgsvX9ufZXxkyS3rYwjRMI84BhrBGA1w2Cmc
xcS91ol2P+c29yVvMvseqCsl9MNdmU4DmsWS4kiFbLAVlIKwfWzxBJisVy8C7srT
h7zpVUiraMONKcElEQB+btwumqdvsr1Nm08+EuEhVzilFs+CayEXJrnXKGU0xw84
1S+NLM+/P7SU0rO12f8W8g/NROGjus+GChaTpeWTUgSNWD/BwkvGTAvTAiccoalc
BQt+2JbNKFWtHxZN3u8be2sZtoWLPpqziCoU4z8tlw4nbPF7qlH04PWx3pplrHKX
rq0dowvYTqKEf6d+kjYLPo3fBu00DXFo8nAjNwtHFa8=
`protect end_protected