`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11488 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
0ivLeOT4zMq5S+D+IkEISBcC9ZT9DZV2X5f9kmsw82KDyrddO6aGJop+nTExFE6k
dAMHbVJkaiFiogP7FJpN42Pr4U0YaJR/UaFEry/PCc4iE9IUVMUMgyKlITfOjQAh
kATl7rsvHeM8kKHohpwwbNrhH5VXfueyMNuupk+rAevwEu5/Tg9rVU/0y8U7SDpN
wP2wfh1pxWCByn4B7kiHjYZ6qFThiVueC/fujgwwoej1ck5EzOWc3JI5qQ+sQIbV
rRJpIIj8nBrIHvULeBRnkjmilQyOjbLO5ZEaGwBdiMBuie8cW5PXPZvAkZQVcoV0
+FC+YqyFypX8hzIFarXvbsJ7mWM9zHR6093cFnbmm9oMBEFA0kKy7pWi2TLu9S/C
RcurJ7Cw745kCOtNSJT6GLEDcneLxkt7+74ge6JH1p8SClo/Oj7x17UBjCMXzlTV
S+ASl9URw1wkfQlYw1Er3ZKvLE04MKB1dKSg+NuyBQ8s9tQw4XjY1r8Z5t5OymkX
+NgH7+jSR5nxg5PK5TZGtELY8rr1k5JKpo63a23xKWC3XqK3ziV6y1OWcxFrzx1w
SYT87nR1QJDp4hzNicaNsiMBbR2R00tL/x8mBqiHcmd+am6+vCBEgbrHslGU3aBs
n82/nBCv8/0fCEJ8YBecQRN1d13PEyUX7yyO490Zr4UEZ+uBS5RgT6O/eFtz4M0p
G1tYXA1nNl7eT7Uwpl+HKhLr9ZFqXcZLHm41P6jtJAWs8Y50oLRbLexyzgVJDzPk
L1MBRN6uoq2ifCE+m6sqEq35CWq9JCy/jTmrInRthmR47ygpW+3cSL8AA+gmwCAZ
VL5TR3JeNjv+xYmMij6aE3CK6hnZIn5BPkkARB11tciCLhxLzIaw1r08pmfpo545
dCoNAqtTD0AjWPTrN6x/j0chPndEc9lQgC4C/cZamSIJUNuvZCT0H4i02lIij7Y9
knH/VUUswGTPdsCJJqRwK7vB6Ms7vCm0+cL5nc8aA4lVgAwz/gQc9Jlf2azBcB1o
X1B5m5NVCcq1Rp0pgQLkoJtw6gg5Ui9X4yOYcUGDnePWaQ+r3OSI0Ig966FxCkj6
dCGN/VTW55easxIhP/ye4byvQLiUy27Sm7VB/5ZZyFi8dXJ8RntTeEXjVOh/XUIV
mlGP3hj9NrwLkka96Fwo2P2claWhXT0BzaMuScXEc5rT8P9x94ncUYPm+X5SCIBD
LBPyEqDBMpaFQOVWeHxWLW1yhWS6EHUFOwzBrZWK2voqmyF6UvePu4MwaCdwfGM0
Ay9cfrHEwfl3ZTPiKOES34Z2sFuJ3NsKPIR18FhMxcVQJJwX38wmMWJ20OqFS4FJ
4ks+4x26yxi3y8NuKFzEcushHn2Cn+UmVchS2sRIhKKRBHwpRc2nmyH7fGOEqWFX
/HrmTv1VD35NywVXZexIIKtB0wzPsMuGvJ+/kd6IY58X0tEGnRHLTZXZnVdi8KgJ
5qLr4LteZl78TVKDon6L6mCbRPglV7vWko1XahhURJWMisDI9I7LClW5L0Jf1L2Y
d6VXB5yRKhMSHGhhtOt1OY0Mqj/AUrK8Y3I3db59fqjF6nDvVOVWQRdGO+MIRQoW
9ykAo/yDNAK0n4Cb3mBK2ULShrEPBiaIkOP31v+RwgLGY8OVIYntQrD3Hemg3kFn
XBUSExoRKZCMQos/781jUdkgIvrC2O+WnYWH4cu4MXj9B8aZmS9RlOwIiylMONkl
comwWf8Dcg0VfXybpjQuyqVU6iqf0uwAzd0Kr82O0fzomS/607p4T7mDbQDh6PeS
tu+3mmVRKPPtnbpu+BXsmkODFDg/FS6/Gu7vYtUe7A/ox94wLZz8h6DIsOXEJXQj
5b/NtcxdfuV3DwI6fY5zww0FLN40253mRNRXTo0AhfOG0Syboq50U779zvSLftQ0
SfSTA9KpZy6nI6ki+5cD5LF/8+4PBrP0roga5cvBNWSJEBfsdqtcgT5lClooSPQ5
XakSE/qyBiPVGxLSvLAY1iHZ2cFMz0m74WHDejqJ0a2CospmgLwu/s+qNBwQo7cl
K0RRxe4K8RlVfPYOMUO31e+RR9TZoSMvoaXNmb6eru2O9AAV0n5jFAwWCqIe/hc8
EOwUOugyz9YrQlUEr2cDiA6cFQChZ2IL3l8ieI9XVIhTPGesv7IhlLmJ6n+JSFKu
jN9tV+6fim0cajI5RQz897EVQuHguLHjXksv5hgi5zfbTOtye9hH0f5dpmTYu2Eg
SkzACOJxLYhH4yk4LzK6t7GtxESH1Iaav/YYYQ97qjBGpuvkv+mM3355PcHmuCEP
X5vs5zKM4dsVfaAHiRbW3mW4KvQq7LHDNOLYn1obYXlKy9o6V+VTGrahmNpU19Ic
I1+5qa80pRkGUzXDk/ePs+RfN0pnOnypFcmq1awrDVU7xgQqzBGzFkJQW2IHn1a8
E7DKRjiL8Gcz5mHKPPsWBhxe0HLqpzF+qDdoSLQqqPostMxnOVwh8W0EE2gWhcek
TE4AZWputYFbr5pxKEeZ10otADxt6h6JfnCioy+7dayG8Lzq8fYVkf7LYaS6BTzn
JmGVwkK+jy7alQKozOO4w3PYQEBi9u6sudg2f+eVu/T+SPyJnW+P50ycbWHPX0gh
INEUQV3S9FMQFO/D7uAHOX1tYc0e2mLI0HCdYQpUhLFKSrbBg9W3Yad6LblTkoh3
thKsKDZXWgXj7F9VyOb6Yh0TtT9QGmIQCTOtLVIbPrWvDQMPpAGn5UpYs0eMzYw5
tyKu3m2QVoslV/FKhAatmeT/qN7MatFjznQhJftrKHJ8UG+ExtzFtwLL0u2XF9it
SINsdZBNyQ2xy3v3ePXrA1OJwwH5tS5iiDgkAzIqR1EgYZV8FPpAu7GDlnfIQRlx
nWAY6rgHwBsq5hH9y+02H2Hp2nK5sO1mLbAo/3W7n9c+rpYjzEDFMZy7Mz4uW5q+
Ars3Xhn7PV5H6hMyls/dPDBZ8Nm7SSImIBSmvVZVEcojTAEgpNtQFNbEyk4rg8zW
l9LpFncMs/Kv4kknat6GeB/pjNFPDHLn05lalNyvR0L4Ej6mJYWKQE4m+OxsYe05
tfU+ii7PWXhL527i2XDLqk/P99QFGth7UseR2H7zvtExFEzuvs4FANPL/uL8IUTR
uQ4Utfur909vdbBHKBA8Vib4l7VEOhQtwU02NamEWi1Fw9mPZaDw0sck4Rs7oNw8
IBk9a4SDN5BVVbfYTW3H/cmvHnxdBrOHpZg2mqQAbb3jD76Roh0xMn77iZchU/Ow
EYrx+kDMVEuWXHw9mf/JMdJogWGWA+TfX+xIgzbRujJp5mCB2xhkkm4RaWD6RLIP
5jaescXRKm2eILPZbc2CBNGCWSw9e6stK/3AAP6AHkpo5zvEGacInIceV9OoCnGN
81botL7WQJTzRWg83wqKKS6bLz4cE7TkHZm4ty+HcSSI87a53FvcPn6XYjoKRfNd
JNFuwZR2/vCVyOubN/e5k03t8CUAXqzAREwlggZrM5sI//hVQT2eed8YSdFa3z+X
zNxaFB6oOOStUrHozyv3Xll37+gNUvxSKyi0lHg2PH9ZkRcYaQ0Bf9pNXG7A3/Kd
CPRKEP0OP4CVt6LGcFPQahaApUEIAy55bvjEVoPnduIbwldkdfmfzeAuuiH8gf43
iyfPtknUb3iH/uXFsV75VoMpEq3pZZElV9sBCu6wiFUNT7eLmUuufZe0DIDgWMs9
ERww08TP5tX5xC+M7Nk/GTc5tq0+mRnKJMEB1cbtYsi91HN0NFMht82kTwaO8iQn
HbareKsa6SjcjiWVraTmhye+qlg32PE2rUGgfqSigWz3L9gCY0rh/rCWAN+TQG4U
nx8gPMGz2o9GTPprzA0JV3ggLP1qNQOxyivYPzSY9YPEN/jfTr65GJPLS8EWShxY
vwOtc8Cv2i3AAUbA9cygKwix2TpuGI8QHyDeHlOaizamAX9NHd6VsAnkjidT1Gkq
l7GGp+D9scowCgvo95H2yzjxfkobZjwBXyKxqt2TAf9VxiDExbqFLYBWVTFoeoDU
ZWMZ+el7R2WBr6BvdtqwiYoy79fw4d0ytNWtIIic2f08yp2BdNvh2xH+4Jwfiwia
fz9wnXo3Ho31SbS38TiAO4viOmnf2RLxlferxsMWsbnnxRqdKW6AwVJJYiHYGqE8
kd66Mx0mAe1J/KkulwbGP+sLGXzCnDNMvUmI2yZO8xRfwBzvloMX9JSKRPZ9Xk0d
uPoERxR+h3G4zItg96dtOHP9zLBZRj5aJSdHcKElWQxK0v0Ro0B8k+vv7Yapv3Bt
Y9rfasX17ZoJGISvF+JyVVWTVPWzhyJcYr86o3WWlsFrFno4t3wBW8s9flF1mX3p
HRCCMUjz0/5vALhnKQkep7GRiCQGr5EMZL11SJjwym6Dw90pdhx6mpJJA9UltRbZ
8nnvk57dq92UXMBxZmRQD5HeHopMG4Sh9HvBXgOGzkY+fEFGnvChjRcl3IjU35D+
uub9yDKjvR++XRxEzLz8TJISsZRqZ9R/WPqSzzrxa1JU6F44GA6MV6okE0sh4hOd
HQVLFHjFEq/66rKHjJACwRd3LQYQ4sQQU3KACa8L54hq12IiNKSFGw01Sf0kDjPV
gL/W8LRM2GX+z5oQMrWLL31JQKqis+7ZBy+jox04scguKxH/59qbXeE+OzmfFosH
M2qLELuJFoFYsr5SHpmUmtN4nAaWTfmmkfT49He6MXE5mZsPrFJhwlgnjWTQ/pHx
/Yk1hZTRnqKa94898GCKHXOG8eNg+Z6srhlHVKd3vc0Jf6JSL2ebe8bIBe8CjjAS
gh3TSA0wCv7yOkca7QvIGtl3UZgnuvzn4Cug5N2xDuTTzP5eIcUUvfRyXJ/HQHcn
d0klDk+z07nCTkKAJxEteg3g2tbQqVgGuxkvxx7dZWWAZLLmAh+GZzNtIFwW3zTM
3TDSR8UxFQEASgl8s6hN3nP9rP0HftoJ2m4KD61nMyhhNJ5YbO1nFC1ZL3dJXfy6
tOjjNujatUgbVM+6/HIWcapPThYc8MIKezfpV/xk3c60zCINJAZ2xLO9jhSlJmD4
rjlQS1v/+8dceuho0KPxPVFVke/FZTCyWHlALLcx7NmVx2knmtQtTCYsehQti9y8
r3fVDycjn9tPBj/zO+/i2IoZA5+iYgz0OLLcPp+NvsUIHc5MqumuZitJp5s1ik8h
qmLosq87aKjiZuDpQW6Q54uSfP+eFML7iZleeIUznR9ajueRUsBCsRHsTrYk6d2m
eXbZE4LPV6yuYrcbRRyjEjtwlgDAF5YtmhoO9tSuDst3RO6Swj9gFr95yPWjWiL/
LHCEf/8koCHvuOECKytezr0U67box/dII4DPNJU6M0IcF5IBynJF6FlkbygwZrr+
AURfEwSHX9BTVO6NDy+V9VkjYRwu4mweLi9gHNKCr89X9rHa9YkugT1kinslvcQC
vj0U+N+dZ8RnAwQ7gMqkSprx3NMfMiiN9mIkAwVKSEVmt9L7v8yK+c7eZBW0rt8x
GFW+kY+Dg1YpIa6CsoIVpclrsa1T1fQOcvyeTu+l5EdrPE33KHSrtANTDx/2kfWt
UxY1IUznIZLagx+scKy2Dx+AFANAmivCMRvbEvQDOhX1Iz8qmXplR5Qg5cURRtLt
VDC02lXqPjCVYTTLmCMLPfqkWAzF138RnmgVpPFnPfxN+TFzVNmXqjDnnT9bVF8e
0uF0PAeunwEGvOqmlgy7+ENy9/aDEOhEW5strcN2zVzcihloXhqfz+PbtLEexUfY
RPVCnFLN86A+DosCbcBigjjEeLoqz6YhNYIOTlp8fxUYmxTiyIbP5pqJNxiGK+Hj
4Df2baEQUNN8nFzbJAb8Wh7Jli6lDww2Psc2VoRKQsugOj4jjo2U8O5l/t5LxRN2
/soOkoqZ/sFeYkhiwtuTMDSJyuWL/c3KSTNeJjhKnTT5W/X4/kKFM/znorPT0sK2
Fu3g+9wtxVb0mCAVuDFOWPXdUnU7861tHwtU5ov0lPMUJW4UTh596XXQHD70bhjX
C7ckHPQC4hbdMczWEa//7DfXAU3qnVAagshfu2fDuGXPQ+iQ4tPjEm42/dmDqr1P
LXmOKH58eWXc27EJjWCfDA1JI8b3CZd/SwsmpfybGUYEMvo4S0JfxGWyRtWWW9gD
v0o9gy3Yxx9/4cHxa+mqa6WiGHkdVmMDKlSoRJhXNQUK0d6d5TdADNAaJa5B5Y8c
WUmXbcM325Pc9EIU550zAd2OrXZJlrdTV8G4cEpECqKgFgw4sLK6ovjdnJOs90pC
u2nhFh+7oMI4QH9YdljnG8YYmZOW+3x6qDInVqt/vKqiMK0HLaMeO+9jMYuvRRWJ
UOvzvG6J8Pb50sNSXVIzpejg8yny2QGn0IiIgiDlnDkfZYPIBUU+TCsmIQiYwMeT
kKktGCVK3MK9iGQnHT+Bh+lmWym7BJdM0pOnFWnI1KlsRdXa/X6O4nYsmLeGrQsF
kmSqvE5G06ly+lfMYG86z/IxqDtsYqvqSTSxscCFtcAS79Ecr0e4Csl6v+mWJNNU
ljJUedNHnVxSMiNAScWjShpw8FtuUw1otMyvKR98ooDjU9vc3GY2J3lK1SpcKikU
IOtV5r7XE62UEXj0voLzwGw99ue0chlI7V741KTlcm/KFDUmayoq6JUWvXbUnVLG
GCSMhuShDwQ4FHVa8Hq/Uk3trN8z2CiMmk4xijHgsSGvVqNRsoZGKpjsdaccRwlu
hRX3t1NS2YJY2yOcW8VHOcEIwIQ02xlHwrn9mQn7/dATJipS6TafR0EN83QS0C6r
a3RcQTJkSbbOxorLPQdnXoKTdgvJRXW7/IwiqIeqb1QuueA53Ycixq/W1xPs9Lij
R+TSQj++FuZPyjugek0JYnCVEkg+Q9ZhMhmZH2MxZwpNmA4vmIVgMbibBEi2rDFU
VPGQOr6guBUPm3qHVv8+wW0xJeNUTnP0P9JlVnKuGZKJWAUdzGmzl3bP6rw9KgZO
NFMJrx2d1fHl/PZDgg0qCYRMQK4kx+Y7uwCSDnuHrRdwzKoDxWGE5anDayxdLiIa
6UxPOuVfHSK+uYGd2S77l3+JUDZCHpG2X7e6J8weM7JJypGLIz0CoGf6WZT29z61
YFjw13sm5UwUFcLAsUgsDaPqG1o/BFasdqIs/mgvjDrZJrB5oUziysNR4mJUfnfz
kCImvS8BZ06gAx7emmi22K6AURLvnLK1kJWEMsVt6/I01hdwXwBe8hEBZcaotDZe
tVkZcx6d/kuhk559nRraOgesCLQHxIowoFG5uZokPBRsGmXjvE4cWRihyuSXQBra
U+P8yPThO31FX0f9Y1xv3XnVVJM00JTikMGUhAljudp6jXtsYUm4mtmeB0k3kDVP
OzbsXWqBJ02zeXqWS0wZcooH06KE9YzjPN+AAuX1RNJfzWaq5Frplj6Y6fU5yff6
KUgQ0KZhUy0j4j2oXq5JH+qd+C2ur0HyCc63F3cJePmsEQJFaNIqmqapc57d3AUs
BtvJX1HZdqdlb5YdiLx0+MUwZb5hWBDWtTEL7a+I14pXJAzpqKtxKWKU8CAN8/+j
mvdcKqlNdNDbwe585Zwa4vfB4WQQf7yzOKOF5G77jWDSFeqz9Y+8lGhYr2+EGWyq
4kPpufOcd9a2leUYVe9d4ELvGdpDQQTltzvU37Xun6a7gVpekSg8XEd/Uymns8AN
aRBL0QKLVWxy12sD8lJHF0VUXPjWThw8Vpob/PsvV/ODNwkvFR54AFQWzIN3QFe1
Ohndu/tFptdZeGsfgQ0zl8juaJR9/v4634fjmkAV6A+aehI0fLVHGO1wuXSnX6XV
1dD26LmwF2s2cSMfbxrge8JM78QS9w3rAwnZK9BHyzq6PIT8mSTWECxQFhMKRuZ6
nOpWhMvoS1fCXpqbaODWBC7MUkzROXNXfYuXZSC4BhGZXrG/LQoQL6rorKdPFMen
xdk7RXXDIw2qtqUeJ5KC7Hjlt9/Y51v6cafYX5kBcZCbqh3eyW16lmoeNwZs1JEr
tOhLrQKCbH2JifkmxPXw6lVU77IykvHk0JT+hgx7AiJL3QdisC56RjRa11PPEMfo
3p0hbMDIbLJ5eBa9eARv5K7DhFV0KD34XnYsDblsHBmn8mkh27gHZFoKMxGYXF53
wvN2nKNc2/jxw/lYshxgkXBDTfOWUcPERT9bdewjhhOAlN4/hO+J5bcXgmy4IHd8
JOPPOJ8gKR0jqABpjgbNtj0n5HrepZ94ckpewmo2XJEFiRLfLLpsCZNB19jhmiHg
58wzYq42XAH8+4VAGSJhgNU0+bOqCGPz874mBvg/D4/TprLU6Vs6xZNDGQD5WAkQ
ct1j8HamduHH7/oLC9PNeLg07wMeLmQE/pkP5Wb0PBkwq9odY+Wm87oiP1YbQkvv
Qa0rftF0pfmAi27hIQheTOcz4HkjXFuYpOpbm2a38HvT568vUAR7Oe0YdnYhYt/k
cnk440FCrEdbsQD0nDRXstbGGE8JpFNiWzrAvT8vkFyKe8dCFm0fpNT1/iH0VJJ6
gAz4nFzlWRv070KqP9gsCn7p747UIy/8fRIUDl43be6AgDG1SiMrr8eby+WxExj/
FrJDuPsEvt2shkMvMWIXemYmitDckBdPGOm33Yrd+Oy0c4uO8rs0BHZGIhzri5nJ
pplfEr21sZmSLlBRDYMB8d5FcW1HceR4L5ffb26HlpuDiKJIi5uIaMTMCM65yfv0
CGiCNJARNQl4sNdKrY2Aiuu+YG5jmvSbES5ZfZGURG3np2qgiYSqUIm1azSbOvDS
aDa/rDo1xs3rxOrSYl1NYCT5OjuuNzDB7gz/sVchKluM/lKh753nHQyfBZumxngQ
OY/KGRIBdNIDkJEYn9lkj+RUkxRPZj8cIS2wm1zmh88pxQWWLE9pvXuv9Lm0o1+z
y10XtvKGIXj8pyIgAJyqpi07rqV9aq0eEHO58mlUZTjeFRRaVon8aq0EvrOPXmeR
Uhbz7XE9zPpZ2zWFOQHOPuBp6Ik32OlbwmyhGbA4OVweSo6scyCgjRhydkx41pg7
Af+7vRGVXdxY9z4JSXL25oB9tjNe4iNB6ZvPycop5dHlX8yJn2UqgJUiy7+LMbMz
w3M7hg0cOHjc/Y/JcYYEdR+ee1NT7/Rrg7DqKkNCF31hl4JwM/HQz5tRSg9sbzBS
o1ajMCOreNUfPsHMkzZMjQPbAr1suFGatcRyHjh30b2x9ucE1K49cLNQsMyPzlNX
ztz+MpS+bblOl6bkwiE9A2aB+z2PaiuuYGZq46votHNnr43xkkdxRW8DdN+77AUT
05sgS2o1ybFHouW/P/eN+waovHCeka+i3MAIlihF6jMy8H+GJe7RaZaNu3yXAB25
273me+p4bzH3pfiJNYBGXAKv9siQk0TEKoxH6cRXtTml2r9P54mSX4CB500jFJyH
ilNAZg4cKXYMdP1vK87d51BTGw8rnkLetlCW8fQQCWCTMSey18OGbbLHNIfk4sRz
gmJ6wXSBuiiu5nmUrgrCjfCds6PkeSha9j/qJm13pXOXL9h3BOJlkxXjSQTKPrWa
0milvVMFwaJrvWuVjdlGle+l7I0cvfiSCGsVMxkmfCAqQisneu3XY310A8u24J54
9ddf/r08Cv3cu1K/im3QWF0CA8jb/J11CZ1OWBsSQKexNH0vOO94BLXui9QwjqVc
wk7yh4i85msgaBrMBGIQ1oW9ISREcN4gwK2atkosftN6aceC5Dwy/PYn061Y3QN+
lvSJT0fVV2vc4Ra3sVTuoUHacRC4JHoxeTXfeszPDSwDT7Y9p7Tv17aft+2JpART
L2hPzgWUBE1KZryELvP9azrsG2MsYyx+G2vpxT3kuCYTIITPgxylPQrEk9qKtIjv
e9zmbUAv/42c61XZjyJDBNXQFAJsaTQonllo36ie7PeXE+9wu2CO1ULn8p8C/dSC
ZQKlOkNX3owI/w7ephuTjqDeUPs4hzaJFgPHE9cgermJxzK5c2R2M7G5Xs6HZ65k
O3/+iVm3d4tdn4pM7kA5J1xpQNogUkJ7oKCRsAnFpRcZBW4wTp5/ssqhiZtu5sJc
OsrNLiyaHqe8K1WsOnBZd6pM+P8abrfvJW1Xhyu3MEFa3hL01pSOeyBJ9QqNhk8J
3HRSnp/bcCVXeLyfryfaszCrvSqYmBX0Ji0OUlv8KK/T+mo6J5z8bQvshZEzXRiD
Ru6+4GZUAk5w+MLkEfTlcMdiKgGYHqUUbGfnk3L834tiAAA0teF0UuMqk2YKl0k3
8wwSq62OYYVHbQgPHNbaoPppa9G3VsV/HeCzrwp+1mKFfHD2UHpdD4TbY4G1Clki
KC7kTstNKS10Wk/3Yut/T6yjLD2pUMKTd/ZEKVVvcN+o9feYnjsgPkHxbbvVvxtE
/RgsrSXv0Gn1t396krOzNbi4WbXYhvgHhyrgbzjw9LXBRrRdVhbHSdY04W52if7i
nqGrVvBKAeICJcnjxpikP8oCn8eaEI6YCSzjSgatsCe6bV/q18o/8AvJ7WKudYku
eq4HXrFvL7fwufhTwKRaWmBQAKnfwZUGbFwJpnZoRg3+xLYNcfD86g00xNVu1xBB
HuswJs3VgHS0rqtib1aNwlQd+HOvIl+BgrH+CRlZ1qBKS3Eoljt1VOv5m7KqyB2O
11LorU61xcY3uryZyMttItEvD41hS3TZIHFAroOSEfRCud9PJoqxe+X+Yx/WQbIb
vL3pcn2StzMr8Ci5WwvW9z6iQW4gRy6MjY/xCPtH+nUTOcf71Hg8Ps14yOjpT8fA
isEDQbs/oulo69LRmxMpLiufx//8yRh2lbXkYqhLZBhUcKyoJEqRlvKxEhpVhT4q
RYl9yFmKqcRodu0DM7LoZIcTuXK1EABr7aDGlnIhwlUK2KDu7WJACtm1ePYxGvQl
apStNwjU6FJdpaFt95nEqxeWGzYQj3uJ2fNrDfLsJCMkvltoJ8Ui24GLeLkxD1qS
wb2D2g2MfpoW7zZ4WRua9aCLnp76JAIAvfTS+K5/ifDxTJcTNr5Ekr08giI7TuSv
CwosJzPVEnH9Mf+BNDDFbS5G2tnkHOD0/2I2/BI1xJgATPoeQtND4Y1faYGRigwF
sCWEAxALDe25Aq0k8aIeWbSwP29YdBx/IMTGz+L0N7Px/KmI2YHn/Zx2rs67N1TH
Qq0Bbo31aj3kasf1v2I8sYM/UO1E27PRyxje7QyCDwMoFQw0Rs1FxDloS0IxiVuU
iZTOip9ma+0JJPpP67NwjwHsSF0JjlxK1yTETndfYq1SkEcquvoFv+Nx/nxdG47l
AZC0so6rz/4eCCwcMbo2wEDN7WlhH1bZ5W6ht0U/psZ9qOaBfFMggfkWwc1YsCAH
cQ6cpojvQMYyIjNSYAJGXD3ylpz9R+ISz4qyp2uHoMvvjoXbolWTSpZ3C+WQ/n/V
6lDT+qv9DjIyHOmMhiThTIlPcBgGNfOdD5ChXR9C8eHuMd4tovlF4K0dDWy8o8+U
G/MLDy5ff8ANGK467wq+/TbnQS0LLesU7Ss0FrpDSa4TKsyFq9/e7V+M3FbB4jRa
kYX7MH4DsbVQdumJOxo4u2CribqCGZIvd4OH2jUWcyI/N86xeUWCKRB5X1LsNOZL
qxrSVAVIVzBIR6wpQqentY7rvhCOH1+Uc10JDIFrl7b5a2FLvgxuWQzViAjjLNqD
rRylu8iDGY3ka6B/iH9elQHpzApgJGEevqPv8cD/kk2OM3mKvoFGMtfgK4081U+B
jQo2NWh4jzU5BZHqwNBQZNy8jvVPE/KVzRvABb/29CRye/AYdAm1fY+NurWQkgyV
Rjo3XP8lhRtC7BdRWXZE9AlhsDl5xUTVhqGgO3XobQL3EhOM+LjOg4MpK82Bn34D
rbVfnAsHeFiRHewEoyDQtR0tGdk5LCuGcy4U2O06bJMIO91HzpjMhJKCVi05Ea2d
gxRprM+fDT8NRA3EeM6kXNfLuLqR6QtsU7khhBZAwi/eIFCHKf7WWtzpO10EYOFj
jjxxGFVaELUGgelvju8lpnPglHTQZO6YFJuAJ8wOXvsKmtMjMv+xbgknk7n+WLwN
M3Rnka6IB9lNwKCvyvLTJWGpRmwY5FRBSfYbyjacojVA0xLzxartRxMiTFBQxwbp
DuQETjNGbOd1ySXL2n5JPrmIUMI+wH+ZyZ16590Mma12LFvlntPgKvEkt9tKrS9Y
U5h8tTSAA5N3ZN3Yh4RvQ15obI9TvwGB6ZJdi2EtGol63i1AautO4Aj/Se5mL5Pg
nKiicO8F19F2bEpW2e0zw/JarYaHZgdNoya0IKXH6lOV9m7akQONHNzoXfqI9oju
KrIIRDTAmQHEfg+QVePHtp5aSpqzoZL76tv77ZEpOhuvygq9wd3y/EfV66Q0gT5v
CpI1myLmhtDuPXHp57Nv4Xn+PCCRibyK4+USl5gU+D5zbWhQhiYUeBGB8YHaFoOO
1T6qmZ6wMBf3XdBx2IlKGHKmMxearC/CodMqVNcffV5UQ9UFuVe6ySKe4LzmqAES
nVtqkqXTN1aeNb43UbWPwmHyaaEsdOGQCGkzeTsAi/4EKyweQU4sRQ22oG74ztU3
/WVbXzGVzZle7Q9ZDxI6R0Vsi9HpxAjiyS6PX5OZEaXi4uYe1+lNPG8we/PYtcAe
IRruJVHcOWhv5iNLuFvgBG15tLyFzKewPRfZL4uDuFCgmc16v8sSHf+ogdTGNF7F
68kyM7O82h+MZpi4aesgIGBUT13afnHbJkfHP4Q7mCEoPhKUc15qZ25U/j7Tq5lp
csXLahP/TpiTtUkbA9rrOGOIK0Juc47tw+2FZF3CcvHQFeAMW0hysPrdqeN+mucZ
RhhFB4A+rUnuodz78Cc9J16VsIbismRU1GdlWH/kxz4zQLiAuR0Bl2ktRjHESTSa
nHAhHM82HjD2/PlDS+5L73y0HBJWxdVi2yObhdGQWkztElqp+UljvfXtDDMA5lTt
7MN633rjwo5aH74PQ6rnwZZrlh3+IrG+ogKA2yiYfYjWBDXTvPljpHsOB1SftDDJ
PwR1dNFDi3w4wQW5aetGrjQ4OD4sAF1yx5hHshmkcfQy8OOCLyaXq86DuKPGy3bX
H+grO22zizX5A8e1ejEVzEiftWV8rG/AEp1e5sd1xjUpHhvxqzYRdlaBv2slWIoh
ZyHoza4XDOLxbb2pjNOlYXuO01fgtBbjQ48xMuIbwgzNya5Y6TyZYfBiIW9E/VyD
PK44yafcdQvlBTI7dChdhig0ThseR7QFTDGOhhQIdfNSNS2axWfmVeCaJCLIiK6h
nycbbO4ljq3o/leP1jXYwZF1deRo/OXWPehuUZz3/HRY2KX1yLStdXPNsezB+ntz
aWQem+Y9J3Zj28yzkrV0oy7+igl68Ymu8xTMSbyw7b5pF4CtfWdOgcVi3a/bHw1R
gTDJMVu37UiSR7bU/2PybHoTC+VUrMUvpWJw7Bi/D+A7efUh3Ve/0LU+jNUbQtQz
mmhcoNal4UoJ3FnzznGU/L1HVFdL6d+a5JdpLIbFwWchgfgPnp9t0WRiRxvZ08UL
pCNL8qc78EUVrueHPV4lYRWQ6dgRusaKqdCF1DrcwXMDsqq8LUQHGw5WWUdp2cuI
Fg53s8g7OjmLyZwuTAR2xaNGtJP09l2mAAzwc0MvWxaoMhjjwZ8CQE23K8TtbZa4
UjV16VGk9Um2WXduz95p9yN4S0WTka8PCnTP8hneBHals69BVdfqH+SrBSd5Fo7F
KBK7V8o1FqRVDXr7EDiCjU7PrTSTqlH/ENSw7ihFt+eFKZxTIcXDaz+DGlGBb9kw
8yGT2T7GuiR1RbxUEpG9AfDKe+3ZwQKAGzjjFDy2TGp7hd+JTfHdglhk7WiBcYye
HeQVPQLsdmyZx2a7glXMTszIVu5LdQP55JDUOYSIpcsYKronZoP2c05VSuJlCiqi
BJuv6gXwJ8Clsbair97y11yPCGTm/CMdtTW7X6HRbHORNdq6RSvVvD15usI/uPyu
Wm3QZxkQCXk2fFwm37Jvw5JYpqVYdU6Hori+eN6n7+PIWkjLEUMQeSMDzBN1r5xx
xDPzM3X05g48aRDxJ4OGF0R5MUuUm7Dfsei9lQBZLEh0cil/iq2diOlLNquQZ3W4
47nQhSvHGDYj+Cfmkvwmwnn/TLkJMf6lQrqEVy8GMo80YQkK0xc1DVRaaszO/wMF
AfWRiWpf6Sna6scIvfqi0R6sHWMEP18ymSqbWlEvKZ3taG5neId5HFK9xZ2imMQl
hKKvFJAgmaJ/+gO2s/fe28Icw4LEGv2q5SZe9ZlOrgcS4evJKj4yn6DmaVa6LiIY
dVGOqzfuPFH8GQ3n/OJy0t/DKBmqO3ylYlXeSEBZKYdIlmoAcXbkj7fkhdUj6NJq
OcNdl6vY6JUkkKxeUBxiyZdZIQ9zCZgNvDrVRIh1SqYn3bMR2556sThYBw3+BvFL
Ej+uSmwyxc9JeWPTbnnlRROkt66hU0K1tUscQUPe2VzYYRjf3RCLLKfLVbo4bIb6
9F/VXzuLGhrCHLiXK/PBLCZGoQXTYvS1vkukKbTYNMnYp369nCT5HCJfp1YarNpg
WrAnCj9MnWNJXxqeLMP4GK3JyBJf4k4Kaj7yjLOPY5b9FpP0TwKjEqVvVBxyW/I7
P//cntyH++DWYbbK6hucJLNHPhBT1+Ml1C1kfpjTcyQAjYHJGrev7JF34LIKjAiR
MfCbcOsDlT75sI3Wv10E1QMV4a2pI3rytJ6PcbR0lgfuayOCXWNCKnttY5C4Wohp
XLcZTVG+30o1GKUX1P1MtCU696TBu8iqxIk2fn7kZh5eaFEk1fNf+69lUMwfKjtw
ZFgzGUkmYUhcZbHwd9nRDnaINWx0MkeX7igfVd7X5BU4LjVFetIb5NeumlaPghGf
lVW7jZjb9w2ZZQdta68hec7pH3yfAbb8RZneT7+kqW1c9TCT49gkOBUqAYVmK7xs
/pooRkr/xASiWeqcLO+ed8tIisSgE9KBuG8OTBBsg8GPX+gGr2dMSIpNFyuhb/ZP
2eAOt+ovn+HJcKMNHE6MN5sl0FYr+J2m4wNNK422v/njfhftPy5kQ9LyUIRa8d+w
by0b7yIB6zoUt9+cLDgyKyUJTXQ8wdGQ4577F3QjuPBA09+tVLTLTDAP3mERZ2Ph
7aE5Y4Pg7ygh1zZ7CT12TH6KtQ8bKmeU6H0bH6uxejMvQTnbWhzK1whMBwzgx3Js
v6qLBPx8X1TdA87C+y3yhA==
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11488 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
4NAZGBPmQSC1EoH0Jm8NyLK/7KbYLLTPz93jnnJuxsRmBsewLkwdtDz1Mdp4q3Dx
bvnkUEb//uzywt+/Y88qMVL6Z10uczieyHkPIgbI583r8DqcPYe/S1p2s+W0lm7m
ZrQSVrdE3X7WqB3t+1xXg273+Eah3IZmLQU1oSpTAMuv2aYdxL+Qvvg3tkuDsrgG
1ha4zvjNGXQVERxX8JLrPx3ZNnvpQq5UqVpsFaikOFqUPFPm4NBigKUsUR0Ktkd2
VAxCL1lldJPh6jPZxNezRPO40Vq69pCIqiZux5AZAvQQR9cOhj9ZeZQaseS7Ja6W
nyQVhASR39o+mw29rrDJDOo4FwYJN7O/YGfBUNFCTixW5TJDbPrTAAUIUqjOWVi4
3RnYk1mDnO1ANaUQWfySjku7N7VChC2xmG1uHNtFTF3gpy7GxfFXhB/5ot4TxSn7
xCTGnYtSYZ5v7aOf0+s5miOe5IqjrfCNjk0JUcjbfqWgc1nMn8Ga94QyUsVrI3vY
v7q9SnNkfWGPuY8Z2h/XHxNl3fAZ+W9/CVgN9GqTgix8Onz6vXW32gCgDh63xs/J
LMak4+e5e5KC/KMGeqztQ63Sr5JDq2aQbz6K4limeVpIl7CpACQSiZHNHBF7+ovS
j4zI9SvmkeQvu65mIJaOJVkRddLBFP7ikSymaNRCOiCN4lGxcDDfskdggipTQ7kE
gR9cOgeKnIc+I8A48HfCDEi4F32QoRTR6UGUSEeLY1hMN2HJxXcRHXZ+KfXYq3Z8
OJwGpllIeAYFlT8B00ocY3q18iYfjUMC5gNpSf+GU2b5OU8lJyYakPSUH1x0taSR
yjNK82l8/K3DBLe3DB/vSoyWdlm6FulU+km5M73G83m0NQs8CUb6WMulCBUIk+gm
gLJsZI/dlsJWuRn4kJ6HE6dNSwQ6ZYc7xdZ6ItOQEMBAeQsSBtCjwesMJBuduZZZ
Dc5/D9SOx2awZk+rpMXghtCmf4qUXM7tdSXnqK7dUrEHnlwEYqRJNwF48K6pkdv8
BJ8nV2aMGG4vP0JnxIc6ubinpvTzJN7ovDnzikulVJA5mBKZP2lO6cs3y1PF9wbj
Ad3zPcQ5zRqivERfwYi0GqxC3CB9bh07H/wZsLRcvFGxfuGr6jGJkFlSDiXURe+Q
Jz10T5CxKFh8e2Evhq6IwWerybcTQ91Jxpj+bfG4qzxRLw71NVzZPFJZ/CBYw27V
bwtTA21Vsm5srYkwYt2fN0Cip/c67UoCJ+mPZS686HXX7HtutGjdFmsFLzBnItQd
U9P0Ef8Qx7fg1hR4X1ZewJu2IjaBsvyW5u9kUt27usqq95tYIfqvfRIPeRiuIes4
7dFfcBCR8bEmJ89V1lIQVtJpe+IzxbBfMsbt4Wly9obHOHmxnCu66Cn5dMLyiDbp
0vRUD2+QgnrLNtKgh0HWTqvJX2ErV4+xDpZs11ioc8V9bLYnFFeRfpm8o40w9H6d
GVto+eBWf/9cf2X328PobAo84ZSv8XGT5Dz+BNRjZIU+mrJadzEGz1WSoeFXGPnm
8Hyh+J+tTY3X+0r3xdw9gIHsxjAmuI+naDL4g3RkYu6fbxLIySmRT26G1i3oxOKY
w9x4ySoqZhl0pFEN0XhuvIaFh85EHB3e3UQbq9Iedrr4JeA3QzNocnsYl0yVFeyQ
xOiKWD50kEsfs6aKgVDekCI1ZI5ENpSlq8qmgKhW0UcVDJmKw5qiZeanfiOnv196
/5TQO3v2ZdQehb7Tw05NuVW1voN9dLFRFIm4ubVOeOeXPlJftOhTaR60A3G/CLUk
SgnaS+5QAeeAZOyU+5Il6NBvCHr2mio7mp9LfIHRFIMg35GW/1hlPO1F3hDnSnAb
zyoZPmLWGzbsPyGg3+fVSXlrbyx8FepUJCbGjzGLJqEL2GJSgNnGWvsnBuR01vf3
WLQDvA4IgHy/4zhJnQlbyjX/qf6nCOvhglNBdr5RkEdxLy32mNl0IBHlrW8OiSFE
i5Evywq1sS4YsDSwjU/kObxGX8NJKxZLEkAphCpb//5Q5shHmpfj51O80xjLApin
3EiAU+AehrOCOu9RkKhnjsNGPhXIwZ+s2lqh4yXy2vA78WKeYRanely7a9jxPjeX
qKe+9p7YiXRDWw+sqxBB8p5OuQJHCxR8P0W28l5jzGb25QJDfSqkAZDxJBmC+w2c
QvcXMg1Eeoo5FJhf2o7npe0BrUnUbENO5ymhq2cvoNeiJLJCtyYBVIqt35LkwRKo
CpkSD0Z+xCR50JTyCLFmB0ffQGGEGXWrlhcBk7adpR+tgUNYIKX4C37T+EIMmQ1E
0k1qm5zL8DlFESYPgLYmx4f0gDDCcDS0Dj1nWFvtqzpbpZZUlKoD1zsar19ZbBME
Frb7wI+/TAmDueOP/+meQtD5LMLllzSxeI/HIJN7CR5fcdS0UCXH78+/VFuSGZ8X
oDAx4YguySJnYbnBy9m2dGWNB9WnNxZ+u/aCq9ootaEv46iptkufUfHiJkoMsJD3
JPLJPC4RpPZ8gv/eE0yNLaTn3Vtfw1Mj3BLnxvr+z5XWpVhZQw/6P+pbF1S+Kk2V
qWjuuUdkuhUooJXMcVfcrdmZzNM2PbxRkZljKZN0TMKtoprAQRJWvjEVgUDYjIFm
6hi7sOEfDSY5nPmIMHSOIPvIZTzUYQeq/3l82MJPX6iw9riasD43DfpAZec8d252
4++SVIfkUcYmJ5UMRfgRsdEc9QIempMRFCUwNQ9eIXJmSQbXK43EPjRvj1Su+8kC
BnhcSZVzlgy9ZY7mrfxRAwmFneX3n6ALhsU7drG/n5F2ZekjnYTzeoM0DgZMLppx
7zD/ispvabNaLQVZrG/4fFkrGrk7aPmHrY7zqqjVA7qOcX75LMbWBpzqKcoiGL+5
Nbm2udYkGW5Xo6koZ0QR9buRC5Cg9ZsnlFSKvz12ZKzKU6X91OYVyA9mJ1OhK0vc
LWjoLy4wA2v+OWJSrILjpiV3g4wGr4oaZdwKkqNoNbkCBZuF1BRQkSpokFAXgQTm
lOijA22GP+spt7oOwbwcANnpUYkkadfn1jrm59nnWWMutxnG4a++278S6ScNF85L
S0Md8JMR/eD3QQ0l5ACgE6b/9Kr9AIJvx7ox0XrqCOxPOECf1fihAvLrS00Kx/il
3HQyoswZbUPlnSSKhQFnppps+ZK1tGp47vUjc6kBvyMZk0G4ovSuW7di0nDhMeME
er7hGYVvRbAItcpVVyOEJEe1L43jSXMxvUGxkCF3BATsFqDbDDoPbsArs2DaEt3Q
UcJ2xpBjgV4eYWKrpDgqR6xx5lf55tHmEtdcQegBDIWMLLHVER1SI/1+Mqg59bwb
mfO736M6gLwpu0dxUsPc9la87c1R/N9386poOP0A//IWD4DUK4xlM0dfSKYaOXJf
hjOU4L8B72W+0aB0jR4Zpm6y4/w3pWAYua2S7EN7DqPCYDyP1I7QJI/i7VG87FkZ
/KUXI3K45hCjvWr9wxO8CVtXP1iyMqIRdzNM27nN7DNv5bA99xghR6iTu3cfZdwu
bXiHYEAGh/ZGcrCSVhTsOvHr9yT/Ny4GRziCPQxRlAOkPDDQMYNIKFGWnoODfOWQ
0zyK0p5iT+OSC9MeqO+Z8fdZgzP2ARQKAzmmzADiiUZ5mPHtDsEPl0ZQ6ToogVUL
RHU1HvCK4ojaojg1wa3PIg46rI/kT4+jq8HvKjR+8JpK7nq+pYndXT+g63f4oNRI
r0ortY9NMqy4+WhRj4ugoP36yPIFFuIBgbTrzpMKQtYOPmsl8c2P3qJs0Z1V4MqP
8HTlFVhyo6DwHUiOLX8uVGdunjaQRcJRyCrMPpegk15rCOTn+y6CryXYBHmwVVI3
+6A989h5I0DAmnfoXnaqawWsgZx9I/sJ81+JeK8GPQtFTbNpgWGywJEde75YeIsG
Edu4aW+PtXIHfiNXWIn0fhHwLhX/h8w6Gg3smVecODmh+HLS9BdDRzWxAUNbUjoa
JMtOrXeJhhj58qeUJswhaqeOuFzkeDgD94eAcFPobQdl8isdkjcXTcCotufxYt72
+z/5+GENR9vwRtIN9ylPewrfV9QBCSOVB55eEc9pTydfsfmmAjpUa3xsaJrizPtF
4mZR2yOW4ia8i4AuWTYZLyvBk0gVFh7usfLwtA5eqVomlxj26SJcXW5utk+g4JP9
SNqTYcogbUbJb97rI1lPDlQXGaladRv114lIVP6wkxrhyM2/3SikR1ErH3FQz2oq
j77MyrcViQzw725uUAgH7iYHlMF4VLQPvs2LeeP0w07FAeIl2pAuZpBen9Uc/+XG
M+dji0YPH0tLogXv0R7IzP+ShnjnRPCSuptjNGPKaNzRvg/VY3sM+VedQ0Xgz9pI
L1Y47Ac0TwWTdMrLj3eUM8xNeO1clFunbK12p+P8xFc4M19RZrHz8bdy1/xcOkJ3
kGpGi+4+M5nSls/GtsRpTgQnIMXtm+kzhAS23mQvrg06WZyrVJ/Es5VFvksh9tPy
DUifGVfT6kOy2iWquaCUN3kdb8sfNdrQO4uNmVucRxxFI/75YbWNlyFR92cPFb1T
tFDLJw1x2BZrZsm2YpStWPUjOGjOtptY+pv0vPx0/jjmFSYAPAWB9iXUcIMxNo/g
h+m4hfddHCc0lUoY6yymvmpOgbHMHBNNcTL1Iom45PEOj41rUJonslvawjcXxPPy
sACe9x3QwBMChTaOx/RfukSVkHITDCXofUznzn6noXzZ0/7JR8x8Qc5+R4z13gfA
PRGCgJP6FIR8f9eJ/VsNXikiNbdRn53EP7mXT0tywXu8VbtPsSCgO7zUJz5uehqP
xzLLgBDJtM+OSwjz9urRsIIwBCeSpiDyU2kVimAAa/GmFok0yprGlBSuvkis0aJ+
OwX80382738V1Ys31y86U2FJ/ykgAVkrHTwpjKdWjMWpu0+rY5cYoSRpIz99/Jl2
x27rOsA8fcRJ4zmrKVSrZqfw0mH9q5QtbUKAkGKkazOoTx1HwtnjBbRPtRMd0Ln3
LXC+l/xT2hMduasdM/Ogeng+TCVPMNHzSoJMj1j5oimD8DrXCUzSBZXUfiI1rrCs
6Iqt7skrl2VpopTBGfYq94R4L5l1FG0H4MdW9kUHPvtWTND2/rwSjznNgga55UOy
HUqJ9UJZML4+yERVLOj+YXsoIvYh6gkwIL/HtkrrsxeAejBwo9H2uwTl6uv4W5s0
5MCVeut4i9zwPRCuN0zatVGLJBPKGSsdwihfxu8ri3AmxGAZWOAhp1Vg0A4I0J3F
eYy136sgcUa8xs4/OasncyVA3CVJysoSr0foymu/kzLaNArB2debk54b+jrv8aak
Zl0DxQt1SUAx2HjJgo7GZf/yK919mMvsPrAJ8fEw10OnsTKVNrOxQx2CNWX0+GJv
bOZWHfIxTF/WIOZ9CmEHoIosY34db1N/YpeVJEU3OzCKBmN8ABlIRAjB2a1xEuQU
EuIuVsqBJCDfdqAlrarmIMrbOZJWlgeduaGM24kc0LeIrmMbr566+sdWJ/eQpeB6
RqQIC3EI3kGvVLA0FfPhiG7MXQ83BhWmgRcP3Mn9ki9dgfvmf6Qpva9JCv/o1GXH
htYeOS//+CRj+VTn7mXz9WI5w29oq33iaujagWu5yUXR5TQY18pLoMeYI558tKqN
KTO24TQfSXwehug6PDTGfIyROfxF1LNY9eUKfpFv8E4dcBgM0eG34v7HYD6+SQtY
781EOBnotr2IFHAc08u61dR1mv7cdRV6DCEERMXESZBeH+0xKUI6/x+CX0mWaH5Y
YR+XYX+zIYZj339+FONMytccneU4ihyu/C0i217E/X5qvKDhZp1jXxDcXFJqOsPZ
JJezyjGDNOMVB/ZHx8xwTHdh8Bs57xNrk35dtucmsmCRWKoVaCRQ4OuR8G97tuFR
knAQ0ZJrEBoGURBZb57ZdV/zZuV5dncziCA7K3Car9jxW+x6vOdoKHNMO9GZiPGX
gtQ9HmS5ABNtkz2PgfxnEOqgLvi56Z2YTEHXCzslhyvWpDzkm9kiT7E48jmf5K5g
qjm6kKo6VbFnl70DBZrk3pLGVzqkwLO2/xyJp0vnxK/b7xz+rTNQ4WkrECnWU4Hs
jtEhABczmUsFZxcsmfwln5fU7Cz1k+UguCkydS3PqPjwYSJ2l32DXfnviWQMTCYT
7cX37ivr7Cb/eKNPsT46+qyDL5RfkUvJZhYU//OCDYMkhHvfLjQvJLMlJGMWcaXv
q3hUOa3NSh2DGtXJ+MVM4CcjIeNEDc2oSdY1KxBy0ofAopcpPUV/tz7zxuSQBEqe
UhGm8otLhpzd6w7coYElMfeysjJel76oMZRs0l2+ybQ3xm7yDQvDtwkSDpjJ8/dw
AX1hZcu3yUmqAgsO3W/OYJBxmPyuQUxkfYjIyACK4zxMLqisADzdHWHcFKvn0H4S
XbD2/mGAl6J0WXAyOuA7Q6dJ7Ee5x5binrm5DSXT82wVtsfESaYlkxIHXfyOnUNV
8y1Z3DpiIX+V+4Y1Z00RrcbuVV+TfoX6P7nTuoAb/kR8vHDAHOrL0Y87B/1E1Qsw
Bzhc7b6+8toGd8pTL26VXubh/eQNg82uXiI8MQAcK/h3LLXW43YJ9WcLDjtQuOgO
KhKp8cy4GfgFvEBMAPkMDLY90U4UI9z2qdgymx9c7mLuLdPxgE64L1DD4tWzItt4
ujiH/J7sr1sPlf+gsBBrXPbP5UA2b06zzm4E91UTQFB/Up+E+WT+Nsebde45YYWN
zq3PpcwC8yezLM52NODN6XxPJTXugZeyzQnc4QJRAXD6dEeFMPpZs7/pora6muOI
Y0YIio/+3zUhlQ3KJOSoYHpBnYnmyW8GrNbl38MJ0+wxDnYTglmzjuF3qqP2WAza
vFmNA8kChZ/4It2bFQgXyQB/K9hEYz+QUoMsRZ2iid4MysjBa4GDA8bORmVX9TDm
U33afCYHMWPPRF+nxNK4YppGIPBYXD0G4n4XkJj7AmwYl3pscOCZ6ZE7opLS8ZBr
NU9sCa56mYJHymyR8aoc8w3kW+3s+tiAKnuizpMt0ITT9hiz2EMoKwcUqi3FHOjw
TGtaXXDOA3VLA7ULYdHFaGEq9qYfif6TORjgOlS0PUMEvDSQQc35/+gA6LzLfgVz
rp3sjyRG9p9Pc21/DKITm66MKJj84V4sz068ycm2qjtoWwMrLHunJs4VwQfAa3mY
NeCs2VBZva7ul6AFOYbFjTEF8w4+IPnZW8rT/gSv7e8lEsFPK53DDFsohQII60Wg
tTnZZZAnpnU8We8gSg/EOoqzQZr5eY33R1Nxf+ywBdKJYSqGjjBar62VZTtbQjvF
bRYRw6mVaoisllNBa2PjDHxeDzT76Tld8v56rkCqzBRU5JIQnUamQGqUIKw1iQr5
94S01t0oDt3PUr6QS/GV39jWWQ2MJW1+3ZPv7aKaFm9clXrG+I+QeT0zY6H22Ebz
Xu7iy/wnDsxtJ0GHywrt0227GUgkv59GRU6LQFPSRS8ISB/IZ5CYRoZr6E9gtuP1
3E10Igu5gKZoY47nLruMz7nR1r/egz6teFQKrHbxo/VuYJ9R5VxxQIAEZcMxlfTy
EwU3oOQi+XEBWCbCHAvoACSkkuf/jbF/zKHaLrLyT9e1QdxHJU+/wr61RBg6P6Oe
SkqMNBMb6hUxRNVXAooGmdCmOqSJ5kmhfK6AtBa0ReQGku4JFDQmCyQNF3vnSbPi
NgPzc0pSJSrT1oIK7jMCoc6BTfSchBubjBdG+QmP4j3wFEPXd3HXCa6hily9sXbF
suplh2TYAxi9/atrp9o9eV4VjUkrtXK1BZ88fttRzj0/mAoKyfXAbVbvl0GEqNPH
cluK6medYfB5oPb9zJZLiK6kH3zks0wl39Vn8V6knpCKJe8Jb4ZQ2jL7NSNnKQb2
L6EkrvE0ICgi6Ek82OwGtlAV/oluqJkK785ffUbnZlgwW1kinTs/ZVMr3CRKA/7y
I5dFn9hJD/oJtnhpW60qBonZ9FqiHMJ/wrbu43KM4ZY8paxl2mmHVS7FnBiWYX88
F6hpFG6WYekzPz7XaRhx5TvdWGUId5LKhUzydBv7ZCNq1M3+aH8RX+S1sxWJCtl3
cNQGJVNXnEXcISy5Fh2H+D/aSXg9Wg9pZfnZnsEz6WMRtt4XFNqr6dZ+H6oz1I9F
6addIWICqNm3wSHmUOX05nYPBuo1a1wEusASExjdhByY1kQfkZFHxVpXpRq7/h2X
MlvKoepArpK4jZMeqdkwmt1qQNUe+BlVC9Y1ImiRo88GZurmKLLWFCeI4CSJJ6lG
WunqI+bZNbnwIAQ2Jb2NShBhdRpQED9WHzLYnCLBoY1pc1Kdf8AbcEdDXC2PMh8z
V1KHm2uN2IfhZ55Cr+O4SaeS6AvVpAne59L+I6T4S8c3T/ha4PTDpfhFCn5+FJWV
T56wUO8ZbY+YwDDo8m9gZODlC7C0V0Ghnatyp4W1B8j8WvjorFyNSin0wmM4xYjP
2yoCXAqnezBQWcZOkQjmATSGxvjazaRm/Ne3xk6Gzj4hjQxVJTmyWhmTvRshmPTS
gAJ89IarDPzWZR4U54atY552wd4Is7YVLDWSRQVgQo2O88z71zgE4cctJPH93gWD
wbsFxCtzUm9VDjJPE2TH2PwNU1xnwzL7WknLpos11qvlFFnySSLQtUS7l1KDJg2S
EA8XLW1lJSYoWn2YbcSq4VFIGkfMs7oSNeJJz8eVAzW1BvDIl0dOROoYkhU56SQD
662JyQ3F2LW6KdwzSQ0j07SVwNG5wAaoIrlDiNYBQsohVakBXjIx720sQav1IIr3
YosOSTWx1Wmg4MLtGgdvodQJfxJfGFIKPXxk1DSEoY8wtaBeyVgW7YZEoW8hNNYJ
WGJTzTg5k/wldRojgOQA/tdtKqoxmd/sEzh4dRtkNiUayGFnjZXU0/+aNssnvK0d
WQBAADJZ197s7n2n+a2zG7BEXonT83n4cHOXm8+cTHnK0Y607erIHhlXMGnQy4Kh
PG6rSJuthzwe2PcEvJKI50YP6qJEwgy+yLX5LpDWFvxVVdjO61i5OYmpDToQbpd5
gHfVTMKdMs7B0j21q5u9y0o74XAKf0go59lUym5nadf7WJ0pjQsV7RXT52qBOkcq
i4pa/HurklI/GyDw0ES5MsxyQSlXBHf7PqNqoWr5sE3jyuyMfMuGdnbQFA8O7vi4
1cNA2/t1f4YscY+RWKc6rKPFMt1yWmDDq5BLYOFzB588B7yC5wVmklEPUyZoetWO
km/G7VOB8bQDJ0DH7blm+ixCfvZJE/cBhO19bSlzV9j4C3TxuizlQ83hxmAiTr4V
RAsLOZNCmPsPmcI1UwbuufALaYob2LDAWfAqs0FiXcd5XSetXRT0vGfFbJ7gNC0O
E/PLKbjpvbNflCVJVySU61IMA8heUpc8QdlM+c83hvXzH3Qo4Xc/L+21yP9NzVpY
p4nWaVmz4m4LHj2yHzGW3bmG50tE63oYpjGS1JEIdya8mHWUAd6wgulCeqo8FQLb
53wMBZBPdPBLG6tB9Xi9ZlbUAycdiSW8aUOgyhdDSEHQ2FhwNImup0+VbO+4LnZ8
9r1KeP/gc14Go6hRudM+eLA0djSmVsoi8hACftFd4YoSe5rAkUX68yiu7vjfRJ2O
dBbrC77694gOiYD9m3oB7b1h/Ig5k90IG2k3zJDgFHEBILskL2NhC3euP8uYZGza
AeKGz45iZdrL+l9sycSl0dE+vdgzUnnoVv8P7pg9IZ5cuQcXwpLTAVy3vcKvMMws
VLzcBX0uvizk3sY/x9/Q4GKj6w14deguxk1Pw5uv4KWVBnd7BSon7FJhEC20JGNl
P/mNOLLZqv5GeCW8G1SbSU3o6bf6qIFvY7FlLh9JHIxR7ES3lKZRNR5sMATqLAN5
Ejzb38X2Nt/Gof/dGFjz+MrhSEbc1fC4tOSTe1sQRicm4qlRTZuhznjidSKrN6Qv
46lVhGeRRcZeUsmQut0q24aspBPO9IT/+FDtG+muBlnivIUQ8q9/CBZIsRHMxli+
/LApeUrxEQ5oasRckUf9qrQikMXspUkmKuc9Gyn+m2FtRDmfRGfIWoyh5Y9Lo5IV
+VVXUhtvrJfRpIdI+C888JUS5quV8+R0oR3+5UOq2i0QU65IW1xor8GyGenU1j11
Ia8k77sIDB5OUxZZHc7VPU7fo9EzBRl1nXY46egPZqGE3O7aH84r1yTE4dZc84pu
2cE/IHYClQunYwp22YDeUAhsP+e6pWQgFLY83xfElDzjtq7kBd9B0tq9jT2GSNos
2Kja4cTp3kSJ4RzDTPaiNJQIy0IUg+74MQRIiR9+0uGz6wPQ0CklbBd/LLq48iqM
J/1A4YWhKXhkoBaOtyKzUd4K8yGnTlHnP6dCo5RaaYP5nPn7W34e6G1o7Ok0phrr
YrKSaKpF7WCyYD4PryPSro60jByftn4D+9HMBWvd7r8TZw6k3M6fGx6dHWqd8FD8
e4rOnGTrtTYUBA79+Auznikt1n/BjZVOvAqMkaGJu9t+bNNxXIxk/foRhmcwb1F9
Fia12K0bGuLBA+icuhONvbHQk0zCWNS2WXwFlQHYAXvqxLMm+Lca0r7phRdD4LYy
kfdID8uMz6qVrRrelon/MFKXJEIhu0XKMP6g7YiiwU00xfmBuEQsko8vHEawAybc
20LfRQLEV7Rbo7+igV9lEvnVYZBSClpvrJFuPla4lQbCRbQWKW44ujOKg5SvRtGg
lMnsub14O1LG9XFd0L0z7ARRyHJookPRPLx5pmryQs/t+I45NlqB4wyJvLU9XJhV
sNAfbLIg2Zxj+dZV9y6UES1+3kHrCxjw3f/uINNls1Fzc02Hq1K6OhFcO33wsEmv
tPSEl6i8TpE2CZFNXrGUwiEVOx6rgYF7JzOnHzT8MC0FuGbZTvQsOCxWI/3EPKL1
0j7jOdcqeB1gJjuWQKyL2AGqtJbG3rLghdfmQjJ12pNNjYRCjQBgGzEve/2qGzyz
hzJlAnMd2/eVzJwiWADwF8Bfzn0blNWQzsB7ZJ/HLMwoFSSWU3mcX60nJqyVAApD
AhPOQk9OdQLJO/c/Yh641HzwwcU6+RoCbw5gRxVSO8Z1LVmNd8jva5ZeWZamBHHd
xD/CcYpmNasfeSxWVXVXdTRApJAXjQoEiNed5ZoUnF8W5W4SXJlzKjzZrmLD3w1u
70mQhkQiK96KSEX9kGJrCJ/+88dkYjXmOIrRAE3bjAPQnVvZfVVwLEzfIaPjjTf/
mpegA88f5/IhYR7pjuag203QGiatjN71FxRROb9jhjDYf1Ebw1YqnJhE2s1i5xLP
g3KtSufDdU8ewASwYrjh4KhV44USBdNajE40s5stv4Z6G66zkCC9IgU986RascsA
pStuzXIFOR84NO7uEsdvJKAyfhkZUvi3tzrkhwFI9OH+unmPGFBjyNGKCmqdPpmW
f0DKPBwxZub4+7m1Tr8wjIT1KRIfxJ3RWT7P/7OYijFgPBHDXLOgz37dmedWJAuK
5vrnUqqbH2S3yFUNWLrBYjMArAEvBZOsTtIFmrgXrKtg/sSzpxrKDUsjOyOjtcSt
dNu9bBk2PH9E4TdkbpiFSdsCJdSmluhjUOxoiaaleuulxxx50DfaMKazH72wArLr
/ehSN8fWnqYdjPJo8L6qa1skeLF3ZMow6yPlqxukyfaetBFIeKkzEfYSXWf2VQou
Sme5t6Jm/rdpJQac+3ZdUBdh0jtekPOsaKDmpraJBvkLqNoC/6PdMZwMZnQe2BtL
1lgEXGO0qQbXXIVf4dp2Hif8DxIH7oFJyMjZxdLFygf9oYUeLoXxumZY9nEX61nZ
PU/M/L340AsKbgmIZtXfdgLhyXPPuhgmiuzilylhS20ekjmV0jSgLwIcwESaIe3t
aAw7dztbcZpJFpsWInXBT0ag+7NilLqQpFpf1figH3fukw5dHIqy4kUEvjmDTAsB
Ci3QcSrdyZjSaLWLi/c4G7212oVhvSVXjiyszO/tLnkaVEYZPjLC6Jv2YPs4IN5B
um5pzmHor0l3EZXaNWZbNxQNVFiXG+2TNdVdshjLy0XXhr3mMC5aaPWCOX/jSN5W
v8rNIud6JPDf8Ctkch6DV7foVHB2Sm69yv0J789yAV2Q40uKV0gHuVgfeOI2hFxW
WWmC49m9L8/YuPrz7lJbmBq7Wl25Sx9MN/4b8UWBM7ixP0ivgmszwFy4dm0Jnp1v
2Wf8cdEjnMnQAqVPnoZTnw8510uwbYX4QVFing71jGdtMz7X3jZSyhsu5wSSgxUm
HNJqEavyO2Br7VNJP558sg3pPpgHnPRidU53pWxneuCkGscmjIxGGXbvlchaOJ5X
VboR7pY2E0yczVidi+9Hj4m64nqIVZmEh310T7daL4lqxcf4oXkUdhInRrwSR234
iX0rDfnyE4C9p4c6TM/9HxbudbNQlrynM50QOh3YxaDZh6tjGEspHUe7OdqZyMJh
2WdPpkZHEGUIqoDNpejKluFaPFg+PQBABQcTL5ExsjJ85z85Yew6baoODiDCRs2a
vU62Jyw/o+h5gd8T8/M9DyxyFxctU11syOr1CrFnWnEaXBkB5BZhSjMnZl/K4vM2
+9Vq2/XASCvHnerci/ahAluP1uk9ljSzjhIeNG0mprQJKymIUFtXnMcDOXOSNM5Q
OfSLgRvT/Z1buDS2NeyfCxHbJLCG0l+DA4tSe+XmU5b1jW5wyuffBn+owib3StDx
1AvrwDUhBLYU7FFxLV8r3C4k+si3o+fT1eKPfPE7QqA/nMMc2f3cDXJOTq0dS1oJ
rHCwlDthe6L28l8IErK8aScSJqhdjLWT1XEfxHKpanKUTkjEXxeQWIu8bSkATLxk
Gd8O7Uepsu9Gz1zfomhY2o+CVvhfu/s/goMLESU8mcklUltMunAXGpAhJfOVvUR7
RvPWxgc+WK6G+3w9NLzUaeIoi9YdqjuNc2eiLGqgF8GFlKddRMp+KqvH00FUM/bu
ih4dcB5BbAsZdB9u8kr8EI1NlPRMSXvCtQcs7JA/8b/q0ptISipI2VtoNStswzAc
IMYL0HZpBbB8+2iTZlxvTY5ALYRUQp2fxai8rz6UXYVZJF/Ism7dCfLezKJJ+ksC
F0c3HFHZDiQkTvRatGoSAeI5urdDbQw0g8yxsa20c/aZEkGTSPLQ77ZhJzeWgxH4
QTCz1KNgo8ijebhC/phD+mlUU7XOsRgpjDH21eNmuhzOn2q4y96HZ5uKhBcX76oW
Kq3pso7H78WzXr/YytssGnR8F+R4OR7Tes9SZRRtAe24rkiOcSd2U/AI/2Yfr6zJ
mM9DsSwo2YKg7WHJyWLCNRpCOlg86USnDddSmf1/dMZoGXOEyd2opBhIjCLBqzs8
OfZyaT/pMiGRxv55TAR0wJuti7KsEY4Xqvx+/Gbl3DwXkrPvNDCGfjdNfOQE4UDl
ObCVKJPFUxn9xT20r7Bjmdcui72SaNjQhY8p0h3mrlPws0fDK4I2BQw1yW5/V4nE
kQI8Cic/z/Ok199CMAEwQOTXWIeyKurEwf+8eKEH7v9EK5PZpt6AqXUb35RzE835
PUWhaGrlgrnSnYW/0vRhPO1+iOpkvTxUf+84PScz5WkO+xmjcC/ZpOP+W3mo/RZm
1eyJrgyOqyBeBMZICpkAdngH2eWbkyhodKyP6sS+Ci2G/AYrmdp1D9l8CWmEhhMS
5Ba7rV1XaxArdcvSMj+U56ejJ44HGzZ6MxoxX+RaLiZ6A80X1fn1ax5ErpEqUTUI
Yjj3jI2wgz4Rtxp0ER/fyG4yhj+GxQhf8Y07CXOjcF36gBtZ14ncicc2kgtR3KPU
ZBiWzQ1jW2lwcamEtjQrmOMOksmeBW7cLJTkRON5DuLFrXLzYODse3IYJSEUiAiG
DsKFzsNCBgKGzFRL2zlZa1l7I+fCn/tOVNi5UyR2QViivSV4uXu9k24QUM3Yr5cs
IKBkk6YH/wFVGwId6eXjKAbYp4WJh9AkmLBZafDpECgMGTdE9dOQIZjn0Z9iLPp8
2e8H2AB6wuRBPS2h4cvP3QX2B/1c7kN6Gq6lpAYmv3G7rb4tm6i9XS1GB4niZQlF
E4d3oExUnv6Lz3GOyRJ1IcV+XkX409S8A3qkKxnX+VaRwx6dSIpWgMV3bzW2XO3U
Wg3izF0dClg1wU53bpjMuq5nOdETp/1j6ItyZkdJfnFUrq/9mGsu7chUdn1ptAoO
4PgEaMvu1cu7P+lgkfBUCYf4RDWP0vbE7cMWl4+MUYxenZfGVWqGglskirSy6uLT
/yeBJcL3wW2AwlcUuN2wSXjboxDVCBhxYMqEIPOl/iLjgi9p5klOMer8Ku/sHo8+
cBsk7y33CFVrV+/UD25HlZiG1y5ovteJMWIoouMGR2WH3HbLEg6tcWt6UF4luA1i
WZoct89qOOTDNE0MwBrySBykxZKVQ/jsAee2oAKBKNPATfC9YXeQeax7eaPc2ZQ6
jrys/NBwN+LtMuP/uZFXSVJfOTy0oBp6F6iD5lr6+krMSgg/AL/RRT7F5Y3x+0Da
rVCGiu/Srjz0RLZ6uq1pDb/6AMEW6H3evXHLos467SOnwOIelfpmLvq896fgw5E7
o3P/CNCf6D8l9dthGTse170XbF/zbRgDWS/wmNm4OnDzTMBqkSzNJd+IDXBocRqu
bYAMLAUXmqz6njiVzI+KVv1muKyizOslEa+aHQIk0wVNz3tuxLgP2/3lwtzMw+/H
UPZiCPs8jG7v2JJZa0CulxVF4XDKAgIXY4qprQ/4W5NNbi3a6O3MsxyafMgdegsa
6IeoYSMJjmaiwDk75VxSB3kgQy4Kf76VUqoTbdrIsx40l46hmFQFm/+FxxnDU/mW
HQXDGEewbuCnmZ/1rw4Ce5bUUueCsQUbYcFiDw/r6rDyN9yFu5KsHLwOvLI0qfvQ
e/EyfbA8VnpYZVjsk1MOc5uwTPmX3T/+bJCGXhtafcGxmijBWlLIaiKl1zRIbXms
o2/HBJKSRn2SrHXoI8qF5PTT+V5hYVqerOuLxpmWuBu1UjJ3pEBJG7B3VvlzXFJl
u201T90NJybBZ+W0yPqC9R6xsJh/GU+Tou/pQKadBKpA8UZaxQB4HSzNSnYbCU94
j/qJCv6fN7/lv/ax2PY2bU9LBfy8IA/CDBCVad8USeh+jLD0D8zaJQFibObTKaGy
QQ8DyTyexyJpL5/8hRyvYCAO3E1FOLMKE3yjCtKx397e9sdgudDH9Pkq8FR/Dodl
ZbRFAkdYg3Sy6B6gAJnNlQ==
>>>>>>> main
`protect end_protected