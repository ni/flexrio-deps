`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 33072 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
0ivLeOT4zMq5S+D+IkEISAGbXovjuQHwtL3OpGyyXYbkYNGwFO7M7kAbU6iEo9XN
/U02e92woUWLyhTwXcv1mLOQxt6waD7nuXRtJr69HjubsW4NCbfGvXWv6VPN7266
RZximzOMcRvgeNy6Lqket7j3ShPfhdENIi1U1KxASmBqbUNYKxuTV0V64S1C+Sgx
jMSRkyLBB0HXjsiLQvKM7p5g9ooVOR8gwLz2OLnz5xMAFprjuPb2YXWO+zbWyHmh
HythInBI56ofzgL5dOXhB8MiNyHbPlHI92vvVTskNzb6OiIgUmwiDeQ6ZU17I8lv
JVMNMg5zz1MwTG6LaLiMrMR5TmKBAcNQ5m/CvHlMCy18TxLIjPT3YVOdUVZbdMES
d13sngHDMSPLrQYSrZcu0pK9PBR+aKXx3eTzpPxDqvrdgDXaFERh8gEjUbVtGAH8
CQWk2nsZ3h0j8Lc4S96mSSTFwWoq9WHeaKdSsOIVrDzFlsuEY86d5tC6tBEBsyKS
8B3UwIFrY9rIzqWiGCmxF6+PNUAdEA9CqI7bxzwc5TqSC0p9COY4N1C0IIULDWKV
19VEau4nH5wn8Hkq3pzzxJy33xQaA59SYuJrTHvCTmFhMbzZ6RsdUf7Dvd3HhhqM
0BoHBNzHSyr4fJ/fW+L3eoOvLYxqs8U9jVz/wHiwFroEiuVY8LP8DpOAW1tEurY0
1CMo2QL7/yyvngBQuxu9uhoc4bVf4ipts2GNOtNuFYNNQX78iK3+PRAN5GGUd4If
MVrwpzgGHg6fLvWwA2shZAvxz/QbOLajNNldBOVytkxxtIY9COnazirZx9SSAeAC
1dUcekE8vpuEhVtZvzfjhNcNpkMaPfE5rYIRzjsyEkMZPl5J3E1fJQSY/5cVp9Uy
AhVKuOl4cHaUVUZ46UPMqyExzpaAFIOZixvj+ULjuS2gF0hvK9IBxapr5oJN9U4G
b1r318oZaSHztlamm+9loK5qqWggxDEXlK2QcjAuHyxQaZw94ZdYUsZCC06ONMZ/
YmBdqLpQ0xqb8LK0vDsfOC9VSlAbI4vQ+2FWjyJzIgMrXrv5gTVMt/PVBJsQnj/E
v+OQTC6wABvbhCJtGuu4ZBCTz2yXssYa7rP9iCg0rZKhGfnxwtrTqbKxo5LidG4H
gDuWj/d62/EYsnIGfpN2xwu1ba3E0tQMgI4v0cftaLInwUzrs4woxgJ7wxAvUhFv
Kvsnxx+w8RLzT3h+H+cxT4RbUdeU50uCwF9PskBAlIWW09egJq+V8kr5/GTjp7tz
nGk2OtOGe5EQrLfyfc6aU3AKZncmJklEEIo9qEAY5CNElfjN20TrnZFTLPfUA9pr
0ttQiROj4KtmR2XftEfmbK8iwMequp5BNB13+tIaR30MydhGLmkzNpJRf6jh/1zy
n1cKMM9hTPaixmlF6eOC8vvYQBvs2X/uwnfgcHyVo7YvtyjCJzkITfaGaKqcqGeB
alOZQR3Tad5aQ/O08b28Eu8RBqpo0cPWp4MHKRmmEbELWvuFqo9UZowS5+1/AHDW
JeRki8JOk1PLTQiMfaxs/WA7FI3Hjp4CD/9jt3TZtJQRcXjTgWRSEKQybKrtuWMf
2FrMTeu1ZfmnibOURpkQonLS5Cgoy3btf3pYMaOEzO1cV+hCmWdqOodB+RVeOxz1
3yLz116btfrQscKbIFObDzN41S8V09FHgy+CLTx/uz9WNu3AunpkUXudJpE+nNHd
Qg02wNOC77+Z+1Qoxe1vDTe2K1q2442jbdx5uJ9yuaaShldUP0kRz/udc6ewLI70
2m4z2BMsaBNiBGMCzaTBnNhdyKHbTkYvpiyEgtGRJZBiZZlawsBmfcX5v3i7Hm96
gP5XRk+GKlaS0u4pxC2gV0+yf3khnnJ0JP5vr+/CCxngOnYhOCs0UfsGyDZ9pH6g
8qc2k/VaNX38OA6cZNrRq25/YseVXr+nE0PlyVXaFsHwnZqEN7MwWKnWKRQodxKz
uVCDC/xphSu5PsB9mP46I4AQTpUxxXrWCoYU8GMdLRzl8sUMilXRE+YCyNoIylkU
IVFvg9xFV1bWQYE+3WAMWkDnzKsfAy82yq0i0iH+5esBMjRIY1LByN0ALyZ/Id3I
shkxpKbn57Vr+jTG/r2fI5RUuKebRC2mD5rM7GhelVHv9B5v7kgWyaA8XpBq7ZiY
0EWfzcTSH21w57TfrrRSkaayYi/nHaBXh8uHlCMk2GvtEYof1eEemv0DGtQKhpLI
cIAXv3JHIpZlXOByemvuDMm2hR+RafBv5h5JI8oG9m1vuGFf+IL845j4mrqOEt5+
Qu77ALjpYkTH+LzF0OKcI5Bq9ImwWTGTUqBk9bD/gvu9nl57S5+ib7YaY7iWfPhw
SIdExghozGK1s5EabHpbQI+RI7B+8xVPMuB2YSP3bAYmQELmjzHKKiA1ldhvTm8S
H3dzO33/feCXorTZ+VoY6WLYv0juP/0o5+nrc6Jp+u/ZPYm/whh98AULqdcReoex
hydXaqGmd3kFJQqhfICvT8yl/UBVP6a1+qrvPwzrGUA0IHk9KVhQDdj6wvN8wGUJ
uJJwWP+Dzk1d0tHcvkrfD+Y74bTeW8jC/0BQS72e3I8R553OLY0ltZE/h4CCbEOY
R6pVJip0bes/00MWnAS7xsGsqwhel9NBGXEEHXOJkkQHGbnEIe1cLUIzE1HOt4I4
5oaPVr4DMYaFzmMqjBziTnyibu6SdL2vC9Y1MNEbef1DLVENwM0X32i/JFsI3Hnw
bnc5RhfxKxvBf8PxLdJPFcPgtoB2HS4FVW6s6MgF+4yDyueAaq5Q04tF5HDXYiE7
il6VnelcAPPWEKX7nvTLeW6xcSAqxDm7WrQ7R7PEsjxKT5MlS9Tz6H30Az1AA32G
H9bVSdyArhiNVG5R6V7Mga62KOplrhf6eg+JBJyhhMme8J+yY0z6OABNwzOoCbko
a+/RNC8PTuLA/xmxIM2PlBeK8GPMmNM9p7N8Oa6De8ootQg/BTj+iXkXmDJmKp49
+g+p53RfWFnRb52CWu1wMTna2dcOdYVF8hWBX0OWBoDBf/a7xNlREIVklgKOIdVh
QLMZiIA/9DBsw1QUR+AACLDxZR9lWpblqQ1AI/4o4xLwNUCYtlSvF8DrAgMj1tLi
bVJm+/VsPrAlrgM+5Shj4nRHwRYcKZokGWOJBWQo1b/wkPBEWqOHcT/R8ZQ/RzEo
iQZC9rCXsNPelYQs/ZlhIGvUNyi8tETWWqO5/o3lMMud5jMIBvO8k5OzpMOHEjFq
FHyFrU4WZLhvv2EDLTx0QOgBxsvMPNAKVdhTz6m3LpgZzreFUimqM6ecGdghuP0k
fkhS3jNmLN9Blrrznbht8mg/B6LffvMNycR2Evitw/JtCZKvke7CeNrg6DU4SMfn
f1Bd6e53ET9QICnmapJKqUxT1w0B4BpkzoIhrT5CjNPZ5WlSvj7Ep3Tyq7eVR0WW
HbetmymUJ2tuz4HNbRJZDzVoKsP2XacCQZVZ4xJO0sJfavCXmxi7+SLpsUIF2nDk
Oo1Z1ymOKq5wX5FFmNv7DwWbeIFl/2U/rhnEwfLCOcSXpY8IwQcuXRjNbWa/7Ljd
5GpkMga77W38fZUsBIo058ZsxKD28k3pwGXE+1XWb3MMzEGpUxQz0XNAl0OBmDYg
y0A53zFMDxW0gnij0POPo04cOWe0bic07K2GXANO/wrw0Z3uS4q/A36wr8tN9itg
2dqAsJpysMq8otwo8Z3Dh13gGCe8dffQ0ubTGXSSdt7PzCGCZFj05OGLQtNb3uIx
BMOmafOwYIAD6AuO+VFtle+EiTomGQeXgl/0Zk5q6031wlMfXISbJwP8h3HWCIZu
QWYF+oKoqAOd1xKinTSoWd/dzepp/a8xFuDyoRnfsjuW5hXUTnPJyDeQQJ38giOQ
xUV32SvBeB1fekVkq2VG4N41gButXxyrMYNo7HwcmiAny6xUVDalQf/NvjBB+yQb
7syLKNxzkmQi33umDED9M5FELGMcvCzH/HPxsF2PrbIzlhu6dtSvz6lh9XbhYruI
XZS6SFSqwc7jDXaezqtToEkZloi54nIVTTTUWworFNQa/UWRNwbXvLfuF0Bf4gea
f+lua/ffXQbpUx6gcRSEbc2Sfaijrt2QG0lEOxkxz97+Dy9tLMisL3buHDmaL2or
i5wbs6Kz52ndySo5IIhblbcM2tC6gR4GDW8d1CJi1lpBB/OWzzxe41rhl0MC2NSs
Fe9IXo0gSQJyNcEusaLoPZv2boKixP8hCMXVP/nSV0G1lh+0PHRnxyd3WCkoqg10
SZCEtqZwFKWc78JV/IM34AtnRSPjTFNN9o0ColHqzETzOTuZI42meUqUSLvCIESV
CZvW2LRgZt/YyLXZl6xRu80GA/zKbV5AshzKqwI97b8pjwXgDa5cSsafv24KSSqx
X/srPrafGydffWetI9nz04I5yAnaIIxGkj+cl2QC6tOhsaz/WiZG0VqSMgluEm9m
Md9nBoZF6YJAWMtutjApUTuSmA3SCtA61syxk+649SjGx/gB4bUJDIf7bLhRvp3t
lkRc2TPb4p2MkRzgYn5FjoYrtKARX8jjGZjza4hUwGW3+DjXx4ORzFzwrtImPPvg
eDhDd0b6D4zrcfjm6rfBudISAFxigNMukXW+wIGKd/QPRCewqYyDED7BZccE5SHf
31YUi6+2GeAi6aa3cBYBL2s5OXXTvOUXleKFr9W8abb4jLTzfAEW8UXZc2e1yY8q
2w3fvCiGBiuycFI+AgZ6qFqEOpXM5dHmSIE9erqwShRqFGAweFJawdVs/q5OcL2b
H/mrANqzSDsClsnD3akIcAGU+ZTnDXbHogEGd2AzG07bvFycFFUoaAIl3HWO4Pe1
oj0f8+ZYNA0c7p0T/8byHZEx6nvAoQHa6+UNXYwWEqG/Tmgdq12teikCFKc8cNmg
fyNLEzVoFsx8tMIHjy+D2qJWrxLafSyvKY9d9w2v9s3bxGGW0VzeR07kniM26wus
HPg04AOHNN+Nekm2j6O29CkM9lwmD4aiJGjgnrxQ1PalPXyKZ/M3iybP7hZbsFQc
PNDfk9P2bO9YsMPEcDOVrSw6Ox+gMQqlXuZ/FBG+UfV/7ytwR12xmJ2Ji9PittIZ
XT9aqB3js8+DR7kA5vtzDIMedqvKr7nKB8hWCblcrSkKTY6rcasY4znmHuw+8yFx
YwA/v/2ioW95XYXC/zEBF7AsPcU06XLfVj5s//xsrIqu7BOfWjRpJgkOWDNx3w9s
urZfAFlkn66A3xC9CHsN4+oyAiAZHL8iaSbHcpu2Nn5ByOPMxBod9iATEbRAKwYz
TM7clbmeAhZT9zXg7JLLRGv+gR6ZRFYQyPk/YAtOORLWhwy7PCMhnu03M1r+J9yI
MI0m3yWdcMHLx9PQn8/APCg6VIMCGoas/w29FPpG79JO51Qrf3jxqQ2ae43QKpM2
QHZwGe1vIjLQbaAHdqsahqwecv9oI5FIFN9WV3rrKEKi+qG766nvR/DzoCR8pAXq
vrZ0KdqqlZZuOtUl6FM03TekWvCp5d/nxkGBswPw3bWtfYd2jkAn57RRepA2/QUU
4pZN/m+wYo2KVHjWd1fP4QPFnvBnAegq7S6C0vc2JpjZi0IDI3MpksSCzbI7CrcN
21IlITQdbNOcot3BSJK/X6XIll4OkzVtiLGWReui2c2Xuq+JiDaT+vEKYOcDshCB
YeslWpk2hdDhCh1jbL6iRk87IGOW1Hy2mK8SjpLAa8N5r/HneaM5cfYxQBbDfw1G
sDRMls9mLuhYx8uYtDzmkFUpBLyq16Wcy1Y6el9nzRIs/SihH6e6tmQiT2gOcMWB
Kh+g+EdVcv/TmB3VoBdkAVVC/S4Tpk9wiNQlAl7KZ/EqUSp7vBuQum5iKpH29+kg
EWpiAvD4orvPA07L9Fyocug7zwZLh2gEcIshZo72e+QwEzaWGp7/AtJrqLAwKfej
eH1IRiG7knDp0qA4DA+q5w/G0xT0W3utQFRXtj1JR11sFr8+n34u/0QJd4Cgz9ry
htWU+0hHZyzMqGcnQEs789ELpJvjlfkTyyKB0wUpDSW+yniTTrq16m3PqUoQwdTY
3vUBoM6Od5ojoqaaa5bSr/I+XkHOcm8DSfpSP8VKpaau8Bsb4vu32+iBIP1KPJta
17fyWUyc6XXhUeJ3SIaKhzXfjplVrkyGOLjBigB6hfGw5tTELTjSqfCrBvRy5Io6
q/ifDNyJ+pJcrPgO1WTcT2EDStFyORB0t3XZsp5WlOSqQrdUdM3a5MChfIUYtOc9
3cx0pcG5CrwWTMRQW3MhrG+L0BxagA5F0BN/W/oAGgJi5ngVqI7mkMAc8AtYmR/f
WlMywaG/48oGFOxgawQLQqkzqEQGxe8mOnDAtiJIzKivmsvXaX3+bq+nM5hS+pmw
43Q9Wa+9dhbGO72WDg0Ga/zpnyWfsVQABqy55D7bywlZ6pry3cYUPpKKjXdW04NG
ZCR3HdeE337K5QfdnhPFs9hElKp5xLyTKp4WyirpvwSFFkjT4Lm1VWRweY3yUWhg
Inz5PtHAM/9XdgXI7a25OUrbM1WlJPKUbyftq6wSw3PQsgWuq7U1+7Ua2RsIZ/QI
xI6on10dASICdudQn6cQQoDfOLTdnKlSdqC9tjcuae1oEWDQFuKBsioTE3dZweRK
XMTMI4AIRAQfZWbBzddotuIxhzz25CmZrUDCLxogccJAl3CB9c9Rm5nUjKmxklBB
gSMUT89A/Mc/lPtqfauAaA15I78PLYliFtxOcwhxDeZwRsIwG7i16/mU4GzFjycM
SPEL1ejrNVZr3l2O0EX+wzdb0Vo22N3cq5feb2Kqu39KPl8v5+dmjmO4u3cQSnC1
D2wD6w3La0HvQnjwJkd8kYpcgy/Vv05kwTv8IOFp25U3QxSThGOfxttdLOJMaClF
gj99eUf0rgRU98MxBNwH3/xYAmDsIRUeX1b0FekhbZFB/xkuHUf2TPNNRAnn0K2N
THC5VAPTH39s6woPFNalL884vNvrQgZGX6d/ApL0TEuN/eCZvfx7mEHaFo59cqYC
+18B3PdoA3W1a4JTBWSnmOUfH57Js885NzQ5LCojvlnDc6QkNOrCSCicP9jR7NAx
JxBx7MdJEnTraukkxhsJtBpHZyQ43V6j9FTqYQPcsNaU5LQg2QET4Ytvh6AeJg1B
caiYH83XaxdqwMYmnDFuRNguajjj37Tg5EY21jOp3PzE625joTfegZtuy3eLYojs
gV/4AJZikTLKPeXQh8yrs+2usadzkGfMEDbu0XGEJ/2bdAMs5igbW67To0SCaQA3
TZ4x7X991KP9ExizHCzygRKyvXBG5otiqOAAPc2vOii0tKU1kpKlUreXIgMknB3L
Di7wzmwfC2BhWcH/AdEBpFKbT4f8DvFZNpzRbhScag0/NIXG0wsEwPeLSanQrBCM
h9NGVgvPyuY70vm00rbg5Ba/stEc8371FK2oPUgfdhnQuJt+dFIllcGn/G7EUVnf
vA7VZJ8ExtKp9n9zWUISg6Bq7EFPMLuERhi2G44+1vbwjXUEfMw02Ny2QeM5OS1/
nfOcDJD5Nr9Fhi4GsaHfYZfSZYHazXX0uHyvwxJWv1z01WwMz5dHoplk/5XaB3r3
bc5Am7zVRMhojGhu6woHQ84GFp2m+EFBytU6+YdZJp5N2OdaOzGkbIRVUDUrOPQt
FJJjrrtvKfqm4e3I0BzY/HvC6R1pC2hPaswxUDete+sNF796/LAR/yP8OL/n0BPo
PMp14OLY4WfxYscM0vUiCgzo9jkh3qHl97GbG5dvc3FJnTHM0PKBBHap5Uiu+EiM
5VdVPi4+IhxkFLLs3FKR6p4ZMIjBjnbooyDbS14GvJ7uupojxtSJxccxbT9tOica
MMwRQxIARF5CEBChK751yEjDGY3G86Oell4HIt/3OfS173BM7xnyRwQZa5AIs1aX
BFl9uy1eyYcdXKjBKKqDwE/huheMYoIVT/4qcWkWQol+qR8/Vx0KqtihZzsTJ/bw
D+/xD1qahU8QW8bh42mCgtfOH7nwsfzR36Z7WWVwRugAZOHES6pbTPkYqknlvV+S
jUrMUcjHqli6yJGpnjeEqxyoHA8R4gRCj4yqkF7He8N32ExLJX3o7PIOntD5H3ka
QhIF8oyO+4v+4XuUS9N3okzKyDU87D4BxBqnBries2EyM/hDDB4aqwTU9s56Kscj
jLFPzaiE2me5qPdV5njT4F+pse3vzyOpn34Ed3RNtAQ4n9GO5VU1Jd/a+mU9K3yy
mV7vvB4vHI84Lch8ShtdWU2/p55a7JwmlTl3MHMIbQ6cAuWK/MAj/LaZTl9cvneZ
7Olpjt4PhOzyl7lTg9vjILfiblgBYa2DSBQSU2NF6UoTEQWAqwrqTt4MXQJ+l2Gg
WCaeTB2TwUnHLY32CGppO3AHEe4txWzI3uKTBysvv3awCn8oTPWRPUihk15QyGsM
aBiT1oIeIN/o6yn5MJp33U/ZLzV+FnGQDhHjj8JXlGpqhSHnLi5z4y6PhQl5o59u
MqyH2in0vUIwJ5sExwLTAhF6CUIgFjdHh6gHy2ZkNU3qssTMuWqTErAKpspc+a4R
Xthy1BucXWToCUlp0Rt3SdwIuAKJsVp02RBYMZOtSmcCk8HYvjEeqCY/09EA+8Id
bA7mQGzIoMMTYRfVVrcZu0u6Yi/+jzCCYSRH71iM3mqi6+qRgG1uA4WKtsQrsZcq
+NXqqjyyUWZ1Lh/6Nw9bDJoG/RN3OFmJqKygeZJmKlpmVLWtOCNfeNCJdODVNs1n
waN5droRy0/PFdScwAyVZ2iQuvQB6ttKwSAJQ3QXxcNUIDK8LwT0xCSpc1RYHHf+
JKWy9/2ZOGwypgQ5cJprJ9tR6pdcxomy5narj5IaI9gCzlEM0w33Tmg6ds7l1mus
i50ayRNXWCJkRuyn1VO46bwdIIEm/wzBMx1sd3ztqdNoaOezDZNsef79YP+uGw74
iu4/KqDVx+8LHRTMHuOTKV1WJG4fbCphi5DxeyHOChT/GNiGPqPeLGlEkm7JBxoi
uMPOaAqkjSbkAw2VJPk+wc+4QG28QaIzDHzE8Bqa9wcovrSgcGDYmzbl6rM6bdXm
1z7KQZWhTUSXSyyzFsOGBJ0iJv5feeUeY00nSFwpweS/eSFAwLesxPrmzgjuHh4k
h2/NJIG2Qs6THlG7ceUtCwNwlepepVPZVtt9JhK8e5T6HmIa6Lyi2iS3gLVXO5Ne
3jKs+J1e/LCWRjmMEFQVEa1iFSL+y3NQ6Q+TFoBCAuSVGuEEWiDIS2sEceBCiETW
znH3gpdYKhwuiGCAALFImtIQqUigb2goWScvcDfvun1CrXVVk+Af8yZcf8rcunyz
wkrQ1AOrhxGYdj/D0jw7/LJ5adwrWga/8exzfKcjfSxB6g/GAG6Lhz+N/HlAzWqX
vF+EeTRUnGDyc46Rjpy2SC109r/GsPLzIthWoRiYvo2Sg7ROnaZJ0gE00g8K0lMZ
61ggKD/s+tn+z2nZN3+TKlEBpX6glDAj0CTnVisVNLTewmvoMTxiSjbPmBrh3e5W
m/UdCDSKlJoOy1cQ4xfnSqn91dbT9Mk2/zZGZG74O0Di+G626/7++Le46wJpVmwJ
wdV1+n8JLUkugwS/RE7Np2wdm9qg+yvcbeexgvqwP1NayYpf6jVgcsAyd2J0jcIj
qTY3Oa+DAfS99edjjsi1aYubyopi+DB/ta+OBHWeb4CHOtbzr++nyGn4QZH32U2a
CD5oS5UdEIDsMuG0ks8OWj/MdJoa1MqS+TaK7Rxk2cyAFCUzosv5AbrlyVVUy33M
adLsKDTsMn7l0Nc9vFzR3GJkATMd9FFsO3VCoSiRYDUt9+MVObM/JuUmXsn2UTZe
QVVAoCp687DsWrzIdBKo9IdEyTxXxxOvRU8f5nV5yxhevee6hDh/sUaW7aH8TyWW
TxRuSktz0nOFntUgB/es8313ZFrUg+gjHGLy5dGZ/Hmv4gB8gvU5ONRJ/72Qb7J6
UgupTny4h4GZFXeOvvVBn62lhM/WYgxC61zuGqn91xf7yfBOi5Ah72yoA2HaxvmG
iszc97JfnU+jRCl6S5odrjxCpvIzLUaP+Jzl+0yvhHYUHXaCRxnwmO1EePR8Taue
wVvM9iPXWyaPPH48dFXUb7VOlQbFDvLLExLGJqwolqOuNsY1P98BS7oHCeL0H7L0
DynXywWPhRy+K4I9EWadlIi05L6qKRq4ZfmQSFrPq7c0jnDTXvQl72fv5G51iTRN
krXY3+13PYKcD0sqcQI0V8emohAyMzDpifE6rCOQfDck41NmXlbt+2uqrvC0G1rO
CKdmbrTmnamr1Q5wwmiYl4OrmTNKkeqyI+inRdNTp6zq6YR66YokE+h/nI01fhmY
YqPvl0+0Yz0AsMSJcyq2Qa+euXPLS+sV0mrQK3nnuVHo0S5UlI9X3OejCPx9sRBu
098qVksbE/QbpVVIz7+QzHg+bSYhTxeUzZLpF38vUhkbjfUt/sl+pUDjY6xFClXl
/6NjObxYdbcdO2dxotcsTkRJ5UUncGpijr6Rw5pxMeNqMbMh7VNPCPVjKHnS601Q
zW2AwDiBPGyK6JvMZUrswip0AoVibHXXqG+7Yd8d3OqOXhko+5oFOFnwfrd4sQHl
LM1izG6IRp5BdH8emuq3Fs/6OuXK6YTSUiP4IF0HYV7cvCt7zsTvKOtaJ03LvgLZ
eRZeXXFSM8DbKnglLK8ITBLnOxlbqTSXvNwKJSlctTk87SgvkVIMFk9RVsTO9H5h
XAW95vdhS+d/WU4IlSZg7bhTPfVf8wvnDz3nheE++0XMJYf9pDT/6SjNiDW+2XXU
C7IDhY3VbrJ2uLVMC/UI1O9LWClO+cWRE3zZI5ApM34QLjK8w09+zcGcHJulp3iy
mc3LBNbh7m9nTuNWHlelsu51Av6Nr2WF6XVuhKbjcOdq68Q9lcaI0Hr1TIgXjNhh
tU/NxTAWYCSvXDxPwxuzi+f/G9/JDFpWNcyZ0S/cjWuhgOrnaZ2feTCPfP3Bd2Ot
47S6Dtj9rCpQpBOiNZUPEnfVeZZHtbuCV40KyRd8w0k8XwO/KdpGMvRQhRopdgEs
ydUQK6Q4eIvykHzArqmdxEC3RBUfiVRb7EFMQzWCqQ7esxQqCwD4k0O5CIl2NnG3
DlZXsnoG9zcmxZp5emY0xpqi8icWHs6ytMxOjn4XEeE4uAZjC347+khHnziHw71a
Ilq7g4/vMLFTICGn27FTv+8ImAszY5OGJ7YcESnJm2OxB7CphV5Z7TcaOzYz3Wcp
U0NUaGnjJq+sxJXCe9FEkAWA1v075Do2UsiEwOuVCfF9bq7e3pO7waKWjsnZxUzc
kRWIncTEy7fqi2whUn3zV0q6h7Tbjm6HdpQ51FAMSpj4gg+ghuvu99v0QyRaxNc9
mMEE8jDz22osM+Xm0e9QssCg0D5NUBiXMLxrFznvqqHTnSXLlMzLqa8avmQp4XCN
8qJrx3HSsxDdcVfuap76p0K6QJjBhSc9yljjKwN8P2jqA3z4Yw6TPOPte/OR+Q4f
C+7MHk1piHRcJ01Vho3Ocw0A8jku3oBW59qeQKQOx+8byMwpfGKzhR79haY6bBvo
7sKfvNVscf0jstK4LMmrDaMn830/RA1tAFC3+NZWo5axKhMSx26K1FrAnGRbzbt/
qUkeYBLsMhKj40OAlTKuL/K1jSApKZIcij5Vz7egrVGcY/zzBhvVExbdUs8PZlBd
uyNeLFkjLSrsYMeaPZXjepWOrSeSERWAk5ewgJzGOp4m9vtYRhrqxlp85d9IT/bH
v8rXwjc+Xv73hHoRomM3j9VxQ/zgBt31WbiaiIb+Z0u0wXjwhdfxrX7Wr7FW65Bf
1XN68eT5uCXDFPTGZYWwKwqMFcvMWYk9TOxiW2+GdVW6DpeCgcr3Lmu+VjLeUZUE
FBZSUTZsu8UQ9+mnNz9u6qIK4Vc7NVGPNqGz1H5HZV82FkmnP6sXy08c8uX+vV/i
9vhMtKzJkroqEfythF9W3UVuhqQo2Ot1BBEO7sX/Ptt3xWQfSq5kGbCHjbngjG0q
zoKLqcMd3KCRG6sLibJ4g84fN9hetooNfQwoQBTh92mNCgY5VmBxixb/q4veplD6
Rrl49N9x/BmFrPK9grY59FlSzM6H4W7TIYfPLzeAq8qScDrMTI3Rqm7hAMladYD6
R0Ct4wAXai1egQiSe0Py/v5DenOaTBRkZIKCrHbIoZevTs77KTL2bqDdG5mHQwz9
f2KIy2QrzACVSKT0mHwTqsF1fB4w9xlJg0P3aT5gG6w+ec+P670kK9ixarQcrMIe
aSprApj/b7qZSFBSH2IyFuPocaAlyUb30apk513UOoOfe8wka17Uj66WNa7QbjlF
uLYe74FGdXOyBCzzP0oqWiTHNVH/uxuEsK/GbDcqnZ7djQJ7hWvKg/LaMn/OXrpA
4QZFSpIP4u0hpShBvU9Y5HZ6qW5LrB0exIp3AQRq/0gwN3zTPYZqvqSNiCnbMxIr
3FdBqMQhOI2Sjnhlu5L1ewsqVTNsiQbuQAOnuigqZvLw+Seu6uwfjw39jAz4SIMk
ap4A467+C//ESwHKdIC8CXxZsTNqEr/GkT4p0oC/85usJ49DsjE9UzjXUtq+hESW
s7sumtJyxlpUmNirpCKC7px++UK3VwpXV/JIQxq6iiu+JCUJHGChqyn8MKrlxThi
u6SMSk6nwwgidrgCcYbIKFnZUo7+fqphFphbXVdbBvRmgJNL5QKbgBuoaAVXWSz0
25ZMnzO4NjcfGbkGZpNg397q7lR12YyuLaFhHMni8fGIneLL2oHmhMJgW4xrqgj1
HPIPVK/aP/enFYjbxfu+Pxvx67hKe38ggzVebyV0Yy9zS+x7o64wIwWZf4l2FUgS
xVGjRcp3tVJAVvYDX8v67uAhjd1RHdSc73rj0xOL1Rm/Hy9gxsDKhGNfmsts2eAn
idGItYHtFFKnIeMpmBZt+7H/mYeFDl0E2sK1s3thSBgFEG1AUSiXnP87tvp1oXHJ
o7Tu0ekDqh+4Nv6AidzRy49oBCFVGD/rBnxbL+Q3ug1eo49YfRtj8TSwmbSSJ5DZ
FHzAu9Qnm+2En/fGvYkLMUV31VX8VP1fbrHU1i4kFcqUNQyGlgCvM9Xq0r68EAvu
H1TFuP5tWGrWwk0dl6f5pAJQWiR1SFapY0z7jE4wAIRZyYsCZFzNSh7BLusLiS8N
YUD5SjuXhCCaTPIeDMC57d1BR4BSrMxZnCmHFDUm2GVH+5C7oRVqEzjterItqCGj
UEsrSIFFct6QofC/Tsl1gZ2gVqZ7+PO8LgHPCStMb+HEszS3gwGX+4BPuNRc+kuQ
iLIhe75fT0Crd7sqlkXpZ5ISKu0+d3KP65aRria9NRUT/MRC8UkgbmcfEtDWmD+S
ThEjC8aILdsqyCR/gV5BhyhpMgZ+Ddl2aWIP1mDYhB1M92sKCfRJX2sUEdeGfXOq
DSDxhvp11UhusISjP9lHG7nXiCkhP6GNDoGXDslWYLgLCJwxPUUnW3RqORynbc8p
bwc8gCmCac/MawoK8eXC7ijxHP60nR64dKIGHn9ZIS3lsV90SyETwwj9yvJV74pW
PAcsTySm0anUYRXGXSdKn+PRfXZRakx3kioWEejiYGcsSGge9ZnYtggB6t1LWZJv
M9LWbDhI85h5nyJGiQMSETi0eZw0Z2BcgaLmqAQswhuW7supdu+VHnUcZ1ubccGo
YIe1MPOCJCGaWnZLBgNa3ITMxojF8rXqoyOgZYZ1njtzVZPabaePyxLWGxZfasxF
2CBB5X5T8v2z8Z4Q9JBpDCLG6JjLGgtOd9iTvJj+f7JcfJ8U7Jb2g5lyu+AJc7H5
bsleIcfY1E+CijFv9SCbDFJ+KdVZBf0n6eqr1315xzYANHBCOSb1HQ1HlmT6/lDX
rUqbwgWD9XxUeiAuQqU0HkSI176ZcJteq1vycflmwJm3/Ob0f6q9PzZgm+Qdz9wm
XNo75o2KTXAuS3RqtShJNVWGTy+U4tNz8yds5V1bIHz+G6kUVZ9Fc/+7FGMnWxyi
iaOSYagHqw4EYegjfMGvrVtovO+zPFFFyOGZAh4P+NPf57MxMMiyrqtmqxFxvQ8J
puqwDdvbKNZ6+MHyDXuGF6LfgH6HPnCzaKCQSm9vTHRkZNN2UN/QaZFQiVOe3Z5U
Nc0jD1itBXfiNcfm8rhSHFziMKvxa9lO9OLlEDKsjOmziwORfxwx3AbYxn1P2+V9
NoQ3qn9MWcdXKIBXxOBu9issQoK2fQv56VGGDmC8TdY4BSpEeW8T9B6/xBB/nDSa
m4yOTTo9L/oLD+5yrHXbDjrkH9IC2Ed5cPndj5R329gBx5uWvkSZg6C5zBuWs7VX
3L+7gULLTsOXuWObUEZB1cja86G0ra1jga3OxBqpkUHdarqlF8RkRPhoMd+i2Yq/
kZLQxPv0Qe+ya26nOwxzFA9t8gQAXWiJH5owZykSTtxWQGGLU5rfBqJuVfHu/s9U
9+4cxPzB+DyqtaYTuvXpofwnlN3qgvsVu5c58HaTKqelmFHPxcZF6RGN5tvrg+ky
khh3fo3tSUVzs1jKesNcEvgr/40Y1zYPdqLxs3OrphDfK9XLUUjUVuaLvUcUBRRy
lousWJaML1ctGjm/6kpMIV6TtnpjajuFdXGl6d7CK4Fug8CNr1Pk8NlAM7qBnALN
wXBlLla+UWFn0CvbMqFw7Mb7f9q09t/NqZ16qHM2aaSfHe0407IsImGp1MJlYGnb
t6jqyo2kvBlwVRZyse6ZGPusFwDjTLxRc9/rSsdMYdAFBtTqaaaOgtz9xqZyAjCU
Ce/jhuU7xOWkJhEcTa6ZSgunKfDV8oU4nnzkDeZDiGmkdXwWXece4FbkitjJ7C1E
CTXXuErS0sl0ULR7GmsL0MfTwf3c2Y/bPCfweVoNuhQBiWTCQrDL/HmxSB/tzgq+
oVl50VUnPv5IS1YqTTbeC6bKhrBynSvelOT/w7hR9hfjWRSwT3KSPg0tAmX+XDt5
7kGnB0NWAIriyqIlrHxNciD2F6e7cpYGuK1Q5QywM7QGYi7PdUVk68eE/BRGbCVI
N8S8dOWBSnij25vmbWfISad9nN1jm5u74GZ5z69cX96PuP9q/pD5uW2C/yVNrf0J
jstoGTd8XYi01xookbU9EHjKlhHry58skLTrs466B8qykdXxwcr9BTmhzR/fzDiC
sxLBiJdK1JJfuWRQ/K/LlojTU7uJSKAbrQU5s7OGds7JKsoevpADyXRy+SR+Fwyv
BdDUCcSgGE3iKVzp1VGINIR112kDqmIb61UchQTnP0GWRdPoACFO3Low/hrKtNQR
R6mRwR1NYSUpfgQT2kA8WE3MxquE/YD85OeqjXLRjs8GtDOWpxbQuVDkNsCEMM/f
+BQCTNGUkHgkUKOeaStUCBlp3MLjmSw72OcH8FdqKk/lrr1bi7cn5/FF7RV9Wv1E
pLn6gQZO3IjZlMFVzTx8nMLnK8gQtNRC5bIWl8TUzu3NMaRvUA3KvHmVIaFT1zZe
URRRDqJSX9Juk5+a+x+F6RHvTwr0tDxybWO7r1x+9sXtXpAVwP2i5FNqIAQf9GXd
W7o6uaTSqc/L1jIME+ok7C+ziH2y9Iu/2dWsSaGR7Ikm6VXvtD123JHorDEHJrN2
BDsPJfaQkpCPPrc6/F7S0tb97jmuqjG9J04RQGHDyH/AcWoy7yL+z7ct9faT3pXU
qcH0rwTloqGPx/G19n19HJXFBJ1b59XXNna3pOAkuCj8M9x6qMTtGPYbh9poI3h0
Yfs+j8bTRspCGSUjolUICZvCWC9PvhtJsebwQm8dJY4ZUrcM9yoJgo90PrrkGLKB
5LN5fEE6+g7FW91gbtMTG4Dte0jMCGJWVJjq+FPlfnevnpAjwT6V8TXw0M6T+WAS
/x3JfG/D/PXG/nha5rLjOmvnu/Ms7v951yXacliJY1TlTQ0+YU1b9Jo3AKwfDU+8
a6B6HJQwXr4neKgxhvLzP5N3EVEH25rY3SuE+ihW3r+qiEbs6uCLqEWsAlVqeQ5E
/CqdPC2L5RPmryVcWdMSJrnSShkNMYlTUHm6fAgz/XEguGR8dtIKE30sN/l0scB6
Chbrgpj6kmZhw7P5if5t1Yv/fowDeNE8hnm5JmwQRIpomLKCFRjGN+rIlkxpM+qQ
afPyTtGOBpWQUjKbCUsYg/u+5mMRWSH8GbweVAPrgLnt0S8xXEaw1Q4tus/2Be8w
XgfxJUk6LsQORzqgYNCZ1xj5n/Bb1QFbTBAD/+zIDJbmUxRF+w6BE8/ZpKof+AMm
23Kq/bs8CWLCjLkEvT1KDgnJ7zpQN4LEmdNptI1m1HsxUHVsPd5BqSzF4iHX+jnp
DeSEZLqfOr9a1oE59wnJ1E+8YPxxQdFkZA+98VkNGkHsQLheYZs86CsJxX0VAqwb
kymRZ53Yyx2Gt+pET+hozS8yu+JelSjaMEo/hSH/pm/6ImRIWnJuEE0qrANaK/xB
GLpJzXB3QjzvJVhpKGL3KEhXy+Zyuuu4quPq/+MoeHJQPyMmXoj1/uM+qJoxl5SY
/Hzk+aYRGIzWo94bGJCKRH4qhyaAJv7AkG4bEr1KjtqpYrhsWluCjI/rdRfm1BUn
9EF9FJGA6PYHQLSwnXTA0En+r1p6+JfQiQCwlCsfOJca8hwIqoQZbxaVVUvKIyH8
m5piZ6ZpvRPN3PY4mz0S3fA7slsrVgu/R+bGYI+Lg4TKa4YdkZXjztG5oa/wg9V8
zUAjtnT3ao7n+Zci/VVSQJ3cZip3aivuVx4iZy88b5wQiyBXBNQOhSu930sQfKq3
e/blIQfoPHmW4LxW53ThY/Tfudk9mXjCcI6aUVGO4VAhsSSsHXqx1VuUfGKh+wOu
oDJjUE00PPxhDWmSPt71xtGL+VDd9RHqBHjz2GIyQjVm5TiPRho5i0v8L0knOVQU
ipV5FIXhe79X+xpQN8S0etaizKQNSOfX+/3re86zIGDNcdPm3DgiOkqJSaU664kK
mM7Fi9rUlZh+7Qi2e0p8f+xa22vy/aD9UH/12jYqeTXomirjjts5XXK7TDrf/R1c
DeoSKCXQbINs71WeC2Nsm2q+p/y8eX6X/qUqPgy7jBpmz8zMYhnC2kTR/FXjAyyy
sfro9YASw2Ayka5swK/Dc0+1ilD+/duo1rezA+Vr8yRnYA1tUCX/5rQsKb7mbXfx
MWv7wytKUvCoYlWF4SSPIcZzwTnLTHKVtZSP5XXurD5rmEhLAb+KuRfDLhNoEZPB
58wbtrq3cUbdrmkBVn8QrIGOKiQTzQtsI5rcVHnMdGfZKSx9873/9TU1wtgCJdUD
n01p/alXpqPAWRNNX3u5d5vazrnWQB+PiBAenCAiElttXN2bgkxPdmimwV7v9K8s
cQ896xwnJYWAK+inhlznHTaiQwjXVIWNQy6tJBBG50So0qHV2jl60FV3fYkBg/AH
GaSfPorUfmE//KyR2BFLQwSPEFoT6a9bPGWcPMiX46LnnsBJDDJsYsNWOmVkoOTU
zRi2vXIJ2CzP6cL5vRGgpASSwAlEeblPNVhB6VO2ZGk6ty1QKpmzPsEEcbVUQZ7b
zBL1I69SIswd10QhpWf3xnDH7/oMwYUB+dbfWy3LtcbhUJ/Myd73r1vDx3N9efbc
O5l0PhCzHZPXGcp7XwVRbX3ZxaqvZgyggYw+p0RxDtMBnj3wFvwGt01kdlGiXhiH
INUIfKlclDyJLe/G2EX3Og7hPIdcxtPyLmyKhjRJat2KYnxsCS02ENLd1m+Uaw13
cCVD3idIJaqLSZVwaS9SbKS/fs1wEyBIcaAqS6aFSu2qU/HxLwh8LDvyhv05j5BF
07Lvb9Kskaa4AAaU/FKDyoNVEQ3Kvks5CIXoEWS58sDlXI2tqyAgOD51ZF6yaCw7
pJangQt8MUU9PYjbIlbh/rD622d2usMGZKRg8b9wq24ErdrPGe0ijbistI4yFQu6
z4lxfn0RslA0tgfDHOQHK3e7BlxolKPVqUtLD8E1sCC4W4cbNuyGdwmLCm0ew4XN
OsVnB0HkRfYx80F4kJvFsYPAWsn7v5WS1hw8d7T8kdqm/Qp5c3LgcUWNZeaHiKGO
TeZms0ymBIffEz9ymscU7/LEESU4h5Y+ReNCguQxFMlIP771j8/xR+pVa8NmJJfD
2fDHslpyLKs+texymQxW4eCM4R122UDyOG08o3iIqwMSlt6GVkGb2kXLyId7B9rD
gjKftc88QCQVs9gNWZelVStqa80vurx00Bn6o5ldx3J+qAKG7OrMpsVvQknB8a1S
hEQvulfUUDgXQbp6NrpCzWGlDZiIAe1Ga/e8NTmCeIQ+82Kq6Gf9G5k8Z7z2Xcay
rTInd0BR8gnw1gWRBXAH9qxi5kUqQct6jY6tbFlNYS+OpjisjONfiAQWcjaaoREn
ia9iB774+xjhvM9K5l/ZMuFd9hMM3HeqQeKUeR8bXGsWbKeQt2PnsIFlZgR8Jo7l
0/Aan8LEuPlfhb7X1/T7H8q9Ec3VhVBQbbYudGHeRLlncL3b/4BLQd5vaCKpr4UR
VyEFT5Kl+Ci420mSLOCnICz43nAygl5LMSkcVLvWoBORbchUThLRYGRGkoD8BtIQ
LuhEn6RH7yv+Gh4Ru4di0pHEemjuaZyyNA0msV++YDAuulgK1pcHxvLicOkbE5Wk
0JnP9Sv4sxXHTJk5+k4gptNULyfK4Th4188XED+YYHj3zlG1L13nanYLH+M+vCWu
SJ+OoD3zUAUmGDnjagMzvwpRao2oIqzrWZloaP0NGWnctt0Od7m2lRVbQiHb4sLd
wdk0zVaKFborszFxpEiqiw6TG1jenTyHxLGpenc9uAg2WH7kX33U/L5UyRJsEx4z
+nOyYApm/i0JD8KPEHTR6D8li2etq4Fs/irOd2qL3Jjyk5o7Ws6Rw7M6vLlsZEIL
+I8SBg3hNlbom8jr65yR4Q9u44O3/jtNSMSTzR0yOjtqqjqCIX4khRaaThE/S62R
EWVr+qL4UXeTAgiBg3s5L+AY5qCjxnJiuZ8dmvefk8O8iDU8Oh0bwe7LyKo2xWSw
H0A3WjD+tY8nA6VaYTRl/fYKwOUsvSCDfYoQtmJVnM5vhojxvfa+50hBDjEiA6hX
vGD+oMjxBEePgBGv3qQvACbBN4vDeOgolLeH4M+a9sHCE7qGV1CcQLoOKL/fWMU5
wtMWbiez38SbHxjhuhj3tRhl7vue6T4xWXd1eidXhntqvRbWxxVQ7k9USALM+Vie
uw4bOVLWR3w4gb68tNFkLRoxUpgZqtb9Ihg5MXERj2O1OoMTkBnsVVgcTOsxF+8X
g1nSN6NxNK2Jp4n1FUqgdgPVzE5Yw7ZPbSMft2ATlBpj0r18LVI0PmUCW0hSN2Rp
LMP9mllqsgeTkirP9M9koBbl5jeCCnuDx4vSW2VSkdH+kK6k17kkxXAcpP3s9vTo
cjWSc0ft9m6r2lAfIRWwgi2qLQyvyvrDRp6TsMW+Eqg8HE6exaTQzym3BOQzpytt
E4m1/2+6qs/HrO+8uk5T6/2GJAhv3cqC+08gq9bv12FNss8IKuPR/DdqaGZLJld6
mqv3j1DBrPUU3Jen2mMBFvtLvBqmiQ7rjiDSg9u2j4xJgsDyuK0EfyOUorW6SY/R
91/VY4slzkrzGGlJRCctlpGBWahCszadNu/nfnGrJJAvtZyazwyf7ueL/Co4Htw8
gZb2c4RriTjtgkESX2VFTcc3b9OuWwDzNkhJ/CZpsc+r+BlFSdkvKi54dTXFnoIa
KGfg+SCD75yPMFzaa7rg1UCifqvKSIEwhHh40VGKTQsb2xHgEsEwiEb9os33i1OG
TV8qahX/JF/hqkyAzi+PwP0gNJnJ2rX37mxl+BapapBNllmVfFmHbMEMJzaYCIYj
BXOPUdeinV6WvzR8FmivDvGSn/Lb0hEabM3hJ1pPjY6ZrlBiNwEf8tESu+z8YR39
gaq3nvztIrGmaOGdycxMXKI8LHYFgYoQPvhTpjnsyoXDAQBslxfBH/HyDCQMqce+
KC/EhOsBh+vmchmyU6iWNOJb6rsoz44Uxk5u7cFXKP8TBV1jBMX/3e6kEGM8Yq0A
HdkAPiDeWNJAVw74zmAd5al+I+UGQskmNObcgVwUS4Ogz7n9LQz4aVLtPqZTZUht
yKt8cpBUyUj07ph3a3+taW2jGQBSGLax1FRu35G2rS8EuF+Mtu1pWmyt3VVjg2Nm
7nmt65pWZfs92bGw9LVfUsPOgTuf+CpjQkAAT+Rhe8oneklR8racPuh8txpmzzeB
kUmyo+HXeKEDqVcG/lnsfaqHy64PTa0gQb13j/kE4U0o1tJT5g6tlGftGkqj+IGC
Z5HjdNnmsWEVSP99gKmbdawJNm6dkQlWq6rkvzljEyYV+s4XEFSZcpvFJntXwnQx
PrwusnplIfujU2TxbRA7q6vgMGp9NCoOEMUyi0GaQ2NAm4CXkX9HTXIsiiryH+6d
z9GbL54jm/mTIj34pYGA9rPkNUqnxz9IHwpAnMrizipglnm72/FkFQ7v0yqRtrZy
tza83GD+7CzzsWn8cn3+rrfd4A7PvpzqyJkoU153x4bG0SjcUqnXrCnu4/G0JDrd
yzcVp2qZlmXajYBGQri4wR2uPRqxX361xBvkwjf3D/kK85f+wfRBaViYv32rePFp
Y5d2CuHv5cNqvtSN2F7uA6eqdZxAuQolUPpBhn2ZM8KgxEs4jBNsr7/UbCqHzyh3
SFs8N5PWcUTEStPE9dJULyXJ42+QkPJe4mw6F2JEuU4l/k5MicLWbbRMHhnds96G
P8KEUZwDDpXXl+jsNFiz+TqXOaCfaIogfQVq0PEwtK9oTOT7wiaEtdWRvs/EOi4E
M87Njl16wIoKjAJpArTKZyFxxI2C/EmCf7B0XUHhyxYGJctac6TqDGGF27QnAtOv
ZNxQbdBqf5hXowMkc0l3ozGk5ZTwEfKUkvGn9+VJ8WdyDJLzI659ZgrHTnEMUTAh
V/P80OeMSnmIIAvq93TI/IQs5QJGL+dsbG0zRm+07vG+PpY+/fvIrAQaOGgMrcnp
SywQHjre+7kBdNJwriyshfnWqDVPY8aVyXf/dRq+3PrpnvwiJDd3isMrnO1k6/sZ
ufosgvqJYntK2h5tYO1G3efPZHy6p6ifE7aFnXcK7MEid+XOje9eTx8uEsq79cG7
HQpZFx93e2TNjBzODUPggtHyTRWAzaEAHdjKRqvlheDkPGWv7w0yq/d/eEt/uRP6
fKvUKu+H56W2Z9gcd12Kfj8XQbvecOtuf+8yFvRZDRKygjJKsUBFA2GCKojPXl2z
46lf8IJ0T6fEJ8+JULcDXgRN524M8+M0SNy9nSW8LiyfVmH1TDNB9VaN4N2lGQbc
OweseI+V1nQHUUnnw79ceR/E7XihEGGLZtVm9sA742UbOVrc+okdBWRHUA4707MQ
Km6MwUdC+EX9yawxm/wMKDO2DC9Xn2zd/nkgIRWxfoiBdwPiQOe0tM6PdKeqThnA
fYSkjq6BD1+U3oDQ2SsZ8LHlVOclQvh4FTPE3pauyqvST4H2XenlbgfgKBxCWp5G
ZMk3NG6PbCBAHPyjyUW7Nwa4HD8hzM0XSrlOvmHB4nyTwASqGwMFDUBOHDe4YqkS
Trr20Db/j//FYn3b0OF0Dr4ETkpbyLG4cZQ8Tom4BBe0YZkPNyM+M8lCpwSG8PLq
sDMKwZE6vR05/1wnHNxGsdmoeHOUXbLxedvmhv/EOqY02hK+IPhyI4NPxyFdKIEk
iTjMET3s/PFXKe3jFpXNO8ZMuhPQBsbrx48/I+2tucJrJZx/4yVkAk0Du6Mh24kU
nkGHpnQoaSWYLgcNMAqyUJvrtUi0cOBP6Mx3mMBkAEyIvBwtZVmp1eTBJc2Jp+aX
w3ozgQIaX/vMf8AH9NWhnX3eD+27wazBy7HL6TiTNhoV83H/Qt+scMV+AHzLHkXg
VSLlh3wzKPJgnBc4dwb7HQVbLZ+noQF0wnitvsGOiGzBQtX97EgF2QTJMxzcRR+E
+hohPdD4APo8KcTZ2oGLlMWeEdNQPtEbEUsM8tA587LqwjrJmltayrfXcLMRaenW
VZ3dkH4Nju5LNxZ7OPmiWle/2U9Ehgx20/1slEjZ3llg9DlHK5ShZCw0NRWMhfl+
H7Yr1WOs+o38K5llDVTgg37GxOcNB9OLvigiUawtnR3OfAu6k1Nvdu5+mMLg6Rbs
v/TLz6LM/by4Kn+RGKRPnp/9WbALXxLGpNpiMKzdIFD08miLlHp7LzYoLMOtQ/QH
udtY+RbPRI6Yc+8ohJuIK3g7GFfAXIcBpbWi/O9tWt1iDj1wG/Hpwc3+9cCMajTI
sIwEuINWKb3gy8yHi8lWAnwfWOE6WHGJ/lfNtcFmh7rnnbZLDAoYUE+vOqm1bhki
veX4UiQvskbebrTZrrq3s2P8DIF83TkqsDTtniwrJh9uJdH+/9ti6bPorFb4IM1w
2NeNxCwdEmuaRYrZFznmHaQvb7L9ZcfYzi/t0kIxJ/eofOwUsG9g+MxPTwpdWLzL
XPfno8CGG6kcxivzJ0SePT6hnXDNixlR9OOC+MI1f5XTNPfOy92xc9/Rs6JiDy18
RQX+9oIc8ze1lr0NI30Uje55Mv8cdgl2JKJopHCQCQzPWs1octIMeHtFp2bgQLDA
nSUMNUcyuNfcn7gcSet163StPNQmY7z6hJCuAvm7jhOAtUs7H7F76AAHh9jj4Gw5
sN5O96ibAFr2IJtnSocVg5aWAHISiR0G5d4bV3eggAN8XebVyBGNAHfmk50Dqv8y
jmTeXEly6B0eFHsd6DiyuqrTuen/0Idb7GIgbrIYxrjZIhyyjNjw2UVgufdNqNKa
O+zQG9YwiQrpEXoSEXkF88YuOOsh/OmFXKWBLblriVlEyjzVk76Q4WY4226kaAOB
Vi3QlPwhkYv0Lv18lio2wf8OcqZL75O/1F2y2bbhVN3Zpl54h5hfU/cbqEqU58/C
298NFlFrN8dosnXRso0oMxu6/KOL3mb5MXSP00fBmLTQuKSiYfmZc6Qgp9GTszNi
IqqJYWd073pSM6NzMmvGJfysLE7c59ZFzSkpNnLvTzCbXXdl9a+42xTF8Hfo1lI2
KrYdmDA0GVfh846HAOT78r4lF8qgn2daSaBR0VFxvWA5VtjT0NWcQSFmoekmwDdQ
vymXYHs34Z/fQTSAFRRQBruNvbHgWsr/bajEu6aK9GjF4dECgnePva48mo0Fl5xA
XJQi1zWRgVG9iNOeC/j+lfRUO7VMDQIeP1RMAH2RChcSfK6fs32sUoGwjJGlGNYr
idwqY4wgDjBSdhKWpH0oQ1DTwNyPjaAeuoeL2G36Pl795CMCMZNjOEWHwUhTk6pC
RSRquh+3quL6OJkRH+7N0lNudWcWRjqLVhdjIBBH3i0ataySL6RUC36GJg/UJOt8
Oz4k0+TDcWTGLNkGlfxsYiLj1vUpRNGJ7kfzNoenYRY4FdRoHBovSJUWBDVHTs3E
m5wROSZZUrtha1M8AZjW1CnkxAfeVy4/uAlw96t5h+IzXLo0yFyKQuQidT15DA2H
CiK1z046wM00b7EahrOvBEgrK+PLg6Hk1HW800PCgkL/wPIK4AWquFZsgA4l1k/l
4wyJgundMNU8e72+dQsor0FR4AbW55b/meIuMr+5O0y8mwuUTyBz2OGwohz9WmPl
89ejQm37z0IYHdaoTiaOb82Mf23KeO5DYcDiyb7qF/lMdRzoC8QTF65DGX79hM1C
/niPT4O2U8eESVeXI3w1FokLGpRR4CvHjGiAUbIxAPbuYAnVCztjNglydyNZhHlL
fJOPSFviQegBU2ZdUNwSNr5GeF5NjvqVBB0CEV7YGCB7QIwJ+KUkkTg1R8DDS0Rh
g+0fLBjQblgmhqgSYXlpZ1Ni+7yBmFBH/b6RBo/km9hIYlTUURkbt92E3KNjBUU7
JamDTShNT4XB0hYDb6inP+wqf7xbAwLZeo6d5fWeHs6N/wkPwr1Yi3a543sEthyW
e235yIvD8ZKVaI2ZJyXr+tA6oCuJeWd532tEmttoQgLxoROFgOmgbPY/2MdXZ1Fg
TM0wNf7qRQAfDGWIXQ37oWpMss43yUXCo+yHrUmHb2X5+RxCWnrL5y84n7MPpbTC
K+rRcrwtQb4U3RLzrjfX0UQ+SZj71kXjlyIs/crOYSbe5Saay+7BgtEzNBv+ofQG
PBKd79ogki3Tyz+K5QhH9xH27yGtgaPaq6fTXfLS5lDRH6uLH0eJ5DOyADUHn4ra
C94vBV08FiTeZRszgmYMLtGv82lYYR8bUUXCJpOSghBHQw3uBA6by01WUFqOdak7
j3Zh0V/bkxZ1LDnsbf1RgUPUg3P+AjQkTFWLjeOZ/KhBqq5D0lz4BxAvn/6/u5wz
t/UwUxEQ3RMFyM35F8APa5kkGsmYgOE54F1Yzo99XvDIsBV49OxcFmG7CiqHcijq
ycc0NqDBEsBlLEbk0Mv2FhIZ5g5IJz/SspPIUH601Em+iLcfJBi5nRSFAa8MIto4
kkfrxxcPxNaCZoQJFiA62eSbDvgeFwM81MmC8TBA1tUEl7nD0gU7hIqI9RLguHPf
vNtNYSmacMEi0RDYpDE0ke9jtZkYA+n3e62mIWPFORDQ7rRuNYvnPaI2nVbHhY84
gPj70YhfhuBa3hk0sQiYLncvwmcyV16m1o2CveuKeQPyU2suEN/dQ4KQQH1R0u1J
NhZYqVnkvFZnXke5W3osyRWqAOqvvuAdgaWsz8iQX/xUavVW3lawZ8aWB/hWnenC
6YGo3YVZsAKHAdnWrc+wpNe5wTDsquuAWD/Ms06X0fQMYAQwm+LvagTpoe8YFtVx
DW+PjyA3pcjJwwRJ0/YLm9J+QgCDeI47nwBmS8n4dHD/J8o32+xvEAU2usBa/vR8
1D6M9ITY6SSPkHQwu9A7rI+FvMs8fzL6ywX/brNG2EueFM8HG6Kr+p8Q1v0voTGl
qe0B2bPsQDtyJKzZKOgvqs+E4I0OTm76Goy1FySSNc6FLkPYxURFmYWXY6rzhUaL
qE+acCB9EUCnbLyJZF0Ci7bn24OPMOUU1xsa17iLMT0kIYcbiQ2SSkBO/r6nc3iu
W4i3ktXPBR+cWRmTLsJZPnbJh57ncd9IV4v3c7q6nI+WmRq3mQb/shUkNT+67Ir3
GQ00OzZfu4mfJ4KcHgkNRC6zgPTcEAx+YZWQfb2S3n0+iVLKlLzhe83Ux1/8LeVU
dAI9IV33aBv7dozvy/uY/O0ueqvQAf8FzNBsMuK0rrClFpI8isBIacR0h9ngBPsO
t3Xwq5TSnLXYe8UP7dLHxVZS3fEMkg2z8pBo8NUt5WkEIKVe9ImHVqyejNB1yk1e
4koJ+pRAv7bJfR/FA8EF3fOuTtrWtFWwjzg0VkAC53G/KRmaFv5smHw0jreA073W
gfSV3ZCuU2ZlvP8aljfdx3ngemzCDmp3DNvsnxHZIaaVM9/Nw4u9WWppkbSCExp/
zXa/Kx/JjVgeIjmjG9h9OqSnMKM2KdAChx7Z8KH5V8Sq/WxhtUc5bJRkmCkxO6w7
dT7mGrgWZveLJXj7rrX5z2hESU/z6Bf+Lgta9uj9IMoSybzlvGC0KJxaRIxUYoeE
m6RZl1TK/pI02mub89/CbLjoXV5wHYgfYuVoEq+qFD0EDpuxjOnaIIPJa5ZsBAmh
zm3bOAX/ePbKAXvv0wMvCLWSLsqa20xk3CrNxkzuzyYi/fGNePT/ZG0xzh9eICg0
qqbpAFqT6L/zwpQ2UNAyJ8KkYhQIVkoyJ2+iQgReC0a8WCM890bJH+RQBYOt2XeQ
UsyO/2tSOYu782TtEpOw+hWVVSIY7yU4JZBEsbB13MXt5E0jqF8gJutIBXmwK6OE
4FetRsece38GxhiJMODy3FVRqMr1Jafwzu0wibV4poj6jn0qxc6WRXO3Zc4fmiCy
FuQN0vTqmcOfOsxkRzCawLnuO3KJh/bSamTpYExk2GVnL3f++NHVXqCQ029z1pjs
VcWQkc0fRc88KMLU42FcZgWiL59H7De6gydq76xplDoYrZXLQXmCpMlxqDT313EZ
ULs3pRJ9rm16j1xH/55bw/+1bNaSxYBnEaaGqSOyMICYD/6hVUCs6exyNPxIVNa/
7X3HoJcLdAP5rKl/hMpMdjFTL8nUM4Lxr2f0Sw3tjrIf+5xwPx7pA+3j5gxbSG1z
diHeL2l//2vPPpNPAOZFCLwU6uuE5YyS1ky3gJ5v39yJNIaCnHe9rzkr9Ncqcntm
bnEQjD1QVee3v52TlukFkaQoWvKqmTQ8HXP5nEgXL9YezCGvsq0f8y9Ynsiu39bU
4e6IfjryP++RZ+kw8kJH5WLnsYDGh4kdek77EdQQLLp9zB9xsJt6zb/Lvf7fOsOT
B4uYeMdu7cfcuAF77Z+3U4yOBhoSjk8OhXAPi+1CsYQYVGTVnoVeE73pf026lLq3
lB0vtF+ESx+SEpEYAD75zhlXn4zdDUVyRiGumYj3Y13Lg9er9gu8XG0z1s2/HmGm
g2pMGqWoxkhTzzZhP7yQeleNWEJ2O8VDMw94L23xs95zdWoetpgJRGD8Jw2ng2rz
45xiOlIxANgmeV7JzPxD63OFO1dMOFUn2HeDLDRCzI/N1Gisf5W/+8g53o/ZS56b
P4swYAl5hKMe7RHBmOOC4xSEQuNqWoMxrYOeB27CGcNba9uma3earUQ8HKwFXvcc
c8H2jj5m8rxRKmK5aoQYZUM0qDjjU+KBR8fNDCXBBFmUP7uRwIHlwmex25XXpmfu
PuMuQqRWjLxOEuUchtrLBMI6s4tyefMfCuqnsAOepOtr1Ftbz2z5YwtxPC/4GxzX
XDAK6r8FCS7+OoHHezDxYuiZh1avMzUJjyWhCcxaJ+NK9KCynj0GzkMGx6SdkeeE
h88MJlLNY0WFxN56I/u+464tzb+agENBYJwdFIMt4/QOTAwednDN64OUcIApQ2/c
sYi4N80sK0cx0SUnSYSDsVjqW9KmQLL18iVZkpXkzn3vjLIj9CWcDtrbJcdWa0OZ
YcXL0B25ZpibXdnUG7mQg4XmNwYBN/SMK92xPqNMbX5h6+nE+/IYcq01pinEOu4Q
b3vTLiY3udAUP/uLRCum6aHP7MUTDOvdlcW3n+XnUYU6YBsKWjFMkI/Pd7oo+tqz
6Vx+KgfJDipAiG2pa+qak8ugJrY8OLnsb4mJZdRZMoXkJjbpxZ8S92D/X2lYR2rN
nMVBiVZcVfhEKY/sWvSHC7X4swYkLvFANdhzWaEl81IAFGDeUzfy304eV0i7F3TK
YfXpJDobd5W6vkTWqcVu0tjcBhPeVQ4xyEbhZ0rSfZBsK8HYBEq/M2bax/cbRG0Q
ySNTg2OOnHTh3TFbcOxb+rTWPY4rFFzW2vtmiwb0xIAZeVtUVl4Otl68Z8t92pFY
Q2Rv/p3C8d3fwD7fwqxX+LZ+hfSV5YpbPsJPxCm/thlbJJG38gkoiBp7ZLghUO48
LTQqrdL+5B/qaDlLn3Gqt3m1Au/YbziYiA6gFix5090j8r5xKCMYlvfXF59bNyU/
pkkfaOJC9az9S7jJl8KWZCyZCeOYs3Lk/f+OAvGCQ8WAdt0FH2v2miNRcgCQBRXN
ydPxrJfpLO8jBoDGCOQGaWPoQpj2XZvRLQ4gmIgAUDmmAXFs+d4kp1Vkk850Ches
Na5zIVeOO0ufTJ7PThltxTPIFO5zI/ujz5zhVSzyqJLEYzmrebfsLDYLFUtR9taT
zKUn7E9gNgbWkDXR4ZFqBYygcYNOKniqezUorT+T/YwRHG4Zw3xf3A98En0XJdlI
gbA11ajBgGgO9N4AeVNH8+L68sBvyBy505akjtqiW5brJE8FzHDNw+j3qmhD3NN+
AkjsS3kxct7nHBVPboBmNvuBzrj4gDkqKh85POVmVKpG3Qaa3cEQwoFtAdpoDnRJ
nzVjqR2cBipcDc6qYu7mL5zhbp2eOdiGmb3db2JX2r1jmuv6RpIHiVBI1i3Th0+x
JNj8neB4snKp6lVoYIsS9CcGFN4BAwrBopbZ2sySqG0fO34FOc2YTK3oa+OHyMzh
1ukVt/0OHkePKc2iSD7p/qAHFKYl7zyEFH72KifHYloBpXvPD8ukGBlWbVU24/8e
5rRY4sz4hxAxbqFLA11ynhy/GoJn3/9Vh6ZeoXFlihL1t0NvPv+hwF5kYdmcrdHi
S/xxUMmYGqONzihf4L5jdnQ68+71nDAj/sVcgH9BBsjrELv1DJFcMWG+qkE00ayo
zF8DyCt7BPC5NsiEXTRxHQhofZKrcRKvSX76Ll6nmWrq9aHpQ6nQY9UwzhD0zJep
bVBVNz2iNi+6X+MH+PGLb5oP+VpPyi4THVGzr/qHblhWVVrNKlaiUCfn5FwqnLGI
gmAm0k4GN6j7+28pc8k0P8dT99s2mwaE9upu11uMd610a/QvSAANLn+kVlihCphh
Y0xVK/E59vuc43XwTzUwJMCVShfr6Fl2/EX3kuzXg8vZaJM6JqHChrDN7gKhaR7H
cInNAmZ+yQs+lDUkDg9ZAZNRbHrn9DnJEtEAZX2oaeB51kZ6BfrFMGo/yaeKo6L6
gsAg3mgi7UWPX+uVjg+yMIcWfF2/suf6BmVYCaj/qWdWqwKFY6RgNCVnknbH0NS7
+PpYk6ARLrRjwQrxRUU8jYAknyj/Wt+Z4sl++Q72Jzf/FiopGoz7lXOQw1VPCAaq
vPqjvDg7hrg5eXeMX+Lm4+gvIJlmqHh7YG5Xbl9jcN0Kmo5mazu53clEsMdO0Q7/
Pv/c/1CjF/7wDT7DrWXaxBW64Bh002sWtBOWeQ4jMq7fqrB+kWnQ7w6Zm8PkwXXJ
En9VzOj/95QKZkPhCifd6OEq6ORC6uSMru6QMO+3u26dbj/AwbLnGOaq72fT+ksM
eLQLdS1lFUTO/n7OeDUwY6xo7WokZWJKU1SGksWJl95EGuqafF6V0dmnvdNFw6Q+
QPXb4UyRTTAKAFMVV5ZaXcKVad8olfAxTZt/6boQyfOvHifUwizoWQOfmfX8Uw0K
mbIs2ok9+yK5XKhJ1eHLU3sV5yy7Ks8l/Gnkp6TvEs1mUwZVJjPGQxEzHpOqgF5n
f6rytk02ykGTVJzO1YOjOB/afQRAlZqAT4KvTqspBU0GleWd37QWr1geRgpVq21/
6GT6j6kDDlsbvU4yp3+JQZgs4ns5r+xBM162h3exbSQAF8iLvlI6XJLzSsdpiRps
AjrhmYDe9JTYbSZyLGoyRja6QpitT2rRzXkDePxrNkjWQQFnJ0Fj0r0AxSX/Nzhq
onYPByMN3Ri9tfIPUrPbF/0lRU03bRfybOWf5LMQkIPxD1XbmKUYbo/EMCTSzmnF
UbqR5lgLZ6c1jZXRatO5gB6b1bMYSGfy7EoRRtjpuuhdVrL/qPx1VwEXdstRUPSe
CPUJ70lIjkHKUxhw67pCrgcHGgJfjM5yokbCj8qCSaYh62YgkPkJWZ33zglXQo5u
Zay7uaaXep4VsD8Yb+0kCo6p1fT1h3arNvhleBg2KaCjQNgBCD+eAS+F0+PmjSHi
BRbHwWxiW6eHySaPmY/+Jv5uIQRTzLDUdKVR00q79TsBvAtQFGsQ7O/HPcGT9qZ4
tJQzzsehNCuv3Qg7BUhDeYUIUKy/9eRUX2HqQ9gvHnha80JZjl052PL7thCXw9db
jyXXgNEWmsGER6mNF7EwwzwUDZ2eLf6+zrCXu3I9/+GOlt+/wGWcz2JV4zEqq8Si
NSAnjhR7Ac33Svlq4qsd5/8QRt4ITNamYbDGoYyU3keIEN5azpQEicY3o/cMbbeF
4fbcuezDm8s2rFBP153aykksiMtTkeig25Vsm4Xy/na93wWnUL9GzjeSzdCYKVl7
bBlHSOKRcPLPdvZ1GP08d9IPEI2DIF5m9za8rPlIMQOjz39xEhafPbalGEwpyOe7
IXINAGjEnpGBsjHpJQPfiAEsvyPz16S/uni+Mm/NXd0B002+UFYaMufqHV4knqRl
2xf7L+xCrMk+dlOfooiauVNrWYAhhCcGJUnmczxXl++L6M0hOP7QTcCKjaaAnGSI
vFK+Xrl90+S2uWz0BT0lLttVLYzEIIBliH4eMogt0g2lMKljhlh/5axAwIwOh9Cf
IyxEpOGvqbH57j46tFwT51qfrjbmqq3YMV6RlnEvt6Imb5Luhw4FkHu5+4YcfUHv
1IyHRHj1PXjUPP+7VbtLBZLhHZ+2oivvms1kGf2hOjxDDnjAj2bx8E9qJvBnYq5O
hlAKck3Ddsi6qitK2GRxr2C/mLHXfBDeaMya1cIEMOKQdA43oG6rA6oXg4T4/X9W
9Q6f93GIS5PXbi7FtY6jdeaNRsr6l3WND0LI6LqxtQt1eSEe+UR/jyMSlZ6AB/LR
pAjMkmK/UuZlOp8JSXLFcG4XvqnZxZErQiQPyIOEGBwi/A7TCcns8VJD1FZpXnEu
CE/bnGE8izoyCC1I3UaRs7ddI2cDTSAofCch+tQJMVUZW9kQOE06z0QNH6BoRgCN
cIlfaw9vzFQak/OYpdopI4VSvZKZ1nAAqXu87LqO4MM2VfteKLJuIzCV4BTBFAHH
fDzJuwO+TDDnaa8w96ZcMhqFkJ8O+FWN/lXyfRuTLv0xS6DEK36dgE/IZDVgvLOl
ibuFEPLsKjbbJJrN3RgFrZ08g1tNxo4XTiwEIIzfJGFLtySRpbF8wGLX5Nefk7gN
3MoZhwVK/KFBgbFdSu+Uccy9JW5ErcFhext/NticIklFwLX0iTx2tX4vfKWHxHov
vJCZCuVI2AxSeg07Jbj8P8S58vJKIERLAFUOCWayJcORnOHnE1ctcA2QucgI1wGk
+iUkInjy6f8PisRKzxOZsQnsHIxOkiux+CAE5ic+ylMRLEZ2IlNsHlIE8UkwoDua
NNGIttEvgPcZxe/NCHB1vzagD7EzTDnRiA/f3Ys0fqDu0xh14W96vc81zrUcx5Vq
gbCEQQ10eOTCCrFQwQNkw5Ntlre3PVUkOSiM0vmwSIZb9dL4NwNZJTyBjJyH411r
ztAosj+v3pMTzICvUSWCHfyAtvEDt7ua0HehIa5759di9frEBowS92BeNe1R4F/W
5H/Ate1aFsZvidJrDKXu0KpO30FyahRsYx/H+WKHAzvzmZVbC3kRSOdQTcnze4vE
XzqhpqL0/EvWTu7edWq4MUuYJlr68SAvpL51MCxtV/Zo0sgcF0v6d3tN+a6VCMbY
5TQ4p4Rgc2ZAHIZLYUX/zHq3iyG7PwzxSEhLuj2GLe1bjEanD6RrM1mujAzboMP/
hrVTqjGRV28PzqmyqmiJAxE65eFo6iTxSiUGAqypNoNNkcf9ZRXgY502YaFZ0JfJ
NAR4r9dbMSVT7F6dkXAAJuoVaXYsEKSVROM/umy10fY5tJLC4hfLxnuumqHav0CI
U8K2BWLlrQQTqROJQbQYcWgeSFnqbHLktOC2V9gE9GQ12G2VoyU+uUgkQF5Xj3oF
Hu8fuTI5byV0yM8noLUjzyYPBTHVH9EHxu60xvBcs4flHk1l62dk3xMKe27vjXzd
fIRewOEuD/mixs5RATz2EfwexK9JuDx4qGC65PWEa9mCaJB8WPoN7E7Nosl7C0lY
YX6rHmI4RFmPCAoG2+lTzxBhK2P6rZt5nLDx3svaXIGICG7y+FUqyiFwBcD91auE
T/nXe+iV900ng7yPnYfTbmgwS+MBe/q7+aJzkkHZwgf43t4tqaWw2HbQNpf3w2lj
Bdv8VhJA3K1YMX5eDspjWsdfUybIhxcWc5xnyF3uR35Az5vhEaXjKPM5pbbAyDmW
dJUmMABavvsivNMAQtZbQfsSLGAWp6e/0CcxUynVBJAXgDRcxTEC84h2Sb2W/eWn
SGb5kb1P8g22aGKM1fcSuViU27obvNJ7BLG8Z/+viCo2/k3HKXQo+cbcKf/L8hZp
Tfujh4oUmeunrb2MdjACLruD2r8IzFt2m3L3lRIibZ/7tb1+YcU7WYCbRzgpZQcB
Sb95H+NfcnCL14doT2AAUNXiqkZG5ER1IoptStVAS7BbBvMxskYzzj+42FoOrJYd
CjIaHJuh5pr2GoCtsK4HZJjrhd4rg6mjcFbCDAYNZremDzTBnL6FXU8c+zaVLWZO
r3sb4klo7LDzgPfzjBKdT6hR4aKd7z+oYc2WmXomHcsPzM0en6teFf0/vXSqB3yW
8s5zzeoL2Ne78v1VW2A7Zi7ZkPCV82/M7vaeW9UFm4AtszjLs4N2CUVv4+ZgK7u9
BwFvM2o3FQsN/pG0Cmzs9ML0lhDruIqyijsLdxtpGA/bt+DN2dHK1BJLlsFW5Fk/
DeeLH3z3N4EwGXittWSigqwBMNe/nINvx3ko51hgHgNqoPFrr1yDiJVx8y9BIivj
xNENP9oBvf0aozLXYKp/DrnRUQ+GFYeSwx2PtHKwbpc93rtrgIjylYJ6A+6MRaBO
ICbTymc+t2f6QINeCmvUFrayRCMAEvFyLWnDdAWprqPbD33Cx3eGylC1lWBH8giT
6iAKXLGWv/ZfLUWQT1Fwyd46EcUx7YPbhYtHT9qTsVQf60XYuBzZnE5v4KNeR4hd
pfqzbhVUEGEVYRgVc/sa6t050b30l2cD1RngmADqd60ej/k7bgMYuPo8hW7inqtE
oNJrefpPzWFCKAvArG3XlGl8KLNTR0O3lXJQ2gexRkIOYIBIlqlC7BKr004vh1XL
P4gVvmx5mLb3eNKaZO6FvfNn/WQBRBMxUc9TrG6j2NNDj/npX0wlr73qmGpsE0RB
6VecL2Rvlcmn7KxNYQhVEGGpuMpEAEsHtuCIiigXaQuApPxwtAvLxws/fQX+sQ+l
18FoQK+HoNpH+bjGMvUA/Qx/4fj9arRbB1R6qWW9lSo9sFukk4U5Yzc+YdBRJdI8
V4hAbSlKOtpQHA/eSC3avtOVoPVAHJU9zVrkRns1xekU6YrQMhvj6w+6pX3PS7zH
njOFCNrmd/MG6vGgJbhi0v3Bmt6f8lX991okyYEzjbKXYg24/fodEzeliPDNXj6U
7vFTLcWfVDdcVjE5olA4/Np+ero/RoSnpgfWhdsAiUcq8akAQQ+dD3QbT8MUT0cH
B9twREqkjSz8myPcS7kJ8z8P9T0v7nGQEKhjCP3rn4cgpSzT1MYecctxTG8i2fsG
ztbHcFTCXWkITUsGT2ADY+K4C3s1iNY0eEvWbjYJ1J6pTb2qt+5QGndss/Et49rc
Zz0JtKybNXkg3nqiMxU/hZVUX2asHnJFwJo33hw7eyn3Ro4RvGIivpQpweuATcz1
R1BRGO+FbaCCWh4mY/SG+6GMVeGSg9YvK9qfi7xvGQqu/54sUOFaTc42XpsdR6n+
iCk074AoFCTVJ98daF1Pycy+xB/OFHE3wACYrAmjhewwfdHL+PGWaftnFd0UWrEF
OHNCiJHntLII/yeDMdheuTGKx6Ms71qC+M5rYqWHGs29kyJ0ZD53V6+LVAOW0XUa
0EI36PED7yw3QHuCQCbRbZALtPEcfrNjEg+w2uJ07sMEeNfwyA1uFjxa4MEcIG7r
leWBT+RbfwCelkAGgQsVtnTr2VxZsrLYykj3W51c1Ypb8mdB8NW1WclPhRlDSzWd
OqSbtBpRK3XoZhUwYzYk9airte4CPPXQRXtjZd9t3B6m5mw7QnuM2k4zfaERfVtX
SawM8iyigl9vrRaGAz1S/lTrwOx7YL/lpffwGtU2H4TNbB5+Agi1iXbmc3lKgImS
hRhzz0uAQqx3wI1j0o1pk0R8KUVU3RJ5tGI7OBc9/0X8b94bZqcvJ1hZ08aX8/Qe
PBu8iYHbBuktmM3bXZn6tNTdHSJmRqYF3On13XvCathfIoKimwk21h5t4G/DTYT1
lsP8jkd9ke3i7SrtK5XVjDV8WVpAqkTNYW//exOU7kgJ6GEok7F8jy8GZpGejz0L
O8+5nsKb0HSiV9gf75VcRevDxkQZ1z/uD1njwvyuYpIQI+E6+HUb4OGMQOw3g+bN
KaJCG39tlVFFiLQBKwoklIQPX6fDVEZeAPjP6DL9kJZWf+fbE1z9eC/1TyZh/6qq
lIAJ4ddUdRVvQaltOsStDPReUdZn9C3TVPCn2smlFuHCsQ8rKKHsGzYmtaRv5uKx
YWo84r4EaH4Td+yhHVA9OqniRjGfc+sfFXTqb2ETDMoEr8mFOUIb7IcDOS7qwCSZ
+cb/ccNXR03xn/oMpEAE7XdRL3GXI1GfnKywrjowcULx7FxxKIttlEHSdACuwYZP
BvAsGsiI88I5C+UojHHTZvAgwVhf6DL2sugWfR5r09vXGDktHiZI5dAw2KG+OjUF
aSakqSNVemHLpH371tu9ZnNtOQWjXRa0KI897shptBW7zKX1Rga8depSeAltBXTj
SrQPJ++ll9rVTHSFb0vSUjUMn1PBcWJocojnUm3G5xlwu/D+t369nzJ+FdVf+jMd
q0OkcdNrZ1QBIUzp4vV9OYduTxB0ydhcyk7IsaGqtLbL2+afk2pCzfyQpJ53rFwC
2rWpqJVwf24EIyaVSA3E2e82ein0lO44sfNszSL6XQhjHjMPLsgDF5dpa3LUHqUk
Ks13cOi4lggmBh3jm+KtZIpxQmwReT8jVcDimQ+kqiv/HNl25aksXXaSQgJvwT5k
XXaiyl4OY9kahveML6ZLTPgkpfsWW7C49JQ6DQQNOk26SjOknRPmolvmpBavCjMP
DPBczLlByMnf9yKcUfHZV3aKL8jyJXY4zGRy1OZvbWazlA7k/1zvUUK3lPv69+HV
cCKM5C0MDq0J2AAxh8uR84s480Bq66/736/vA7S0N30E7ZG6wknoYln4twbipKY7
KsFZbzeR19eE8E86186BEf46vfXQ0QRjA47/dTN0QYetdejq+/Y5mvCwg8VcxDTZ
VbqgkYODC7WZ1hc5hfrteNOH7kxuFVekdnYGxkV+ordvrWzctCdUG2YhsxryfoOn
PwDfuxkLRFPqSw7swCGVhv9RrZOWUNfiskaJFF1QUn1nN+8TIUwNqapYD8kjQHIF
f7zLPkj37eQhGRlhvxOW74cTHeAFZCFTrt1zfLCHMn53nola07+jZxgwB2OL1ePE
7C5R4eStaIjHd6lDRb8IY4soDKFFTZrTrQ0Ur4z6xL4T8OEARNsZT4gtqmU/ps8k
ztKQgIsIPOJUt3E2X0804GkLd1laXWPo+pyFPkc8qIdIURi+xzi52rrj6xEbB7Uq
W50qZfSaGhncstOJTkgJmCXqjGvIMFjEKmezYNQ6hQQ5JLFoTT8ePAq+evqZXKG3
VrTDHyQfDh7E4dJZZ6qhy0guWFJfus5ibhUtUCzlwQYirHA58uQ7h5R8GEA6Hmcn
N4SoyKz2y4g9H/oeTh5H0dfNTISnlBGCsN0ZkL86kkm976QNWkBQdF9unkbW75UZ
tePMZ4+36qjtt2JR7Xvz3wiVlTnYuSyRTeb/+MQtVUai8xlou6sRjt6q7Y8/mbk7
+DvQESDSjCt7TJA7/qn6D/IY7QgbhRKKWDViMNFDFMtuan+e6Fk+7VoJlt2V7eNd
U/bGtDPP7+E7Ax/F5ZeY0WJxia7JP65Aw9EIsaY4SKNk4oJBnplVWejpbM3Ve1Ne
MKQ7uUD2cg1wp4g8YjJH7N+C75oW+vXBz7Lr+VTwXH3BeVuAeiEaE1mwtvjgJN4y
Wk4Er30t1BCnUZ/knU/VH4L4R0WaTkbhih0p8ZK/gzSnxtkVCOvP0ZvS635Jqz1+
OObBXjt+zkIXPx6A8dmLXJY3c2rEurzK7oPdpTRfOB5djzY98zY+chThilT4UeVT
9kZTBs5luEKXHtO/UnhDM4hizj7ZForYRrTLzgajjIC6QA49+SCsvg161kk80K6U
83lhZNM9UJqkk6pfRBqetnCsQvyVV9t0BWr3hPv7RTa90APetVVohG0Zg4kW8GNd
hk5mOW+iCoPNTPDsQcYFhiI+ZZfrLfRrQcvq2O8OgreGXdPGRgJniCPrsYvr+v2E
SI38yHHRNzkhKQbP2WRamm8UWLPzvpv/xEsf2aOoHatH27rRnNQDGsGvPhVaWHA2
T0S5TcR4BQ+W+tXOk+lns1ao7fQFP8n8PcXmaglCr1xCUAOmo2e9aB2zlQy5ZbvB
yHaJlP2QECyhRnjOlUg40vAC9rugU1mmIw/v8ZGGLBvMllhBLIbQXsLOlxA/lJ2k
MOGxHITc4T0Q09+LXFdBo+k7d3fI1Wmji/S41QloYMKB4SOP6t/t4oYwCyQviwjg
HEXCzVaDed5iz1vw/eMgnR98Yg7+Jk14M9R52MpQo5T+eSfI4n76Eo7gHn1JWfJG
z99MovQ5fEGaSxjvDfYMIyHft5PvYzb2z1QDk8cxjuMgBtzFsxJqswwwACjpW708
YUqx9bTbmSPLrb1UhQOpvejY78DsiP4XT4NmpNVusFTxYnmCK5jsCIwZ08X0ifgr
DuEvNEJmw5kTZ57j3t0vRNrE2dkdv1Uis4Wxi3zg027iLhQVKB4kFBHGhDPBhPYb
xjQVEwRoj0vNUPnbpJ/IefUyF0SxJGSEmuNFskYNBEVirVkZqe6wPSQU97w9V5w1
MDuOH9GlkxOYqcLceNSMnEe+SLwvTU3ZbU+2UmvNpKw8sJdiQPjGXXeHP9IubFI3
bf1UWQV0j0hu7LRWZH12oUOCDwT/bIxqou3HWrvQU6RCus8+YYM/UoU4ZEFDIsFm
sqfBPa419Pa3GiZolByI+ElpUT/Jcawt8xZhbkq4Iy+UV9ScWPGmDJyY7ZdcsaJX
3KiN9i3CyelB/PI3xqFHekZAHPrUhKTvn06LgegtduGa5pBIbBLFtMwgcTDoD9Of
QL7si50EVEDNSMOVfaNFwCxl0VwtuA9fJkR/XXvBV3bPsiVlU4k+hOmoGl8XjXxg
z16FLQ3hVcop5nxpsY7EVRXULWrwm9ug4BIzz0k4Yjj0mpfcuWsouiNb8mHliVpl
Iqylzo9KsKqtWJAyxvTXOiBtm7S9IxH7XQYqiSRdStMa54tmXdGC57p+rwM2ITGC
a/FJGWvloJ5ccmrEjTU1KSdGKPlzggCgIbrztED1o+Jb0yIVcHVimVlZE4fVAT9U
zKUJoN7FDEJMXdB1WZGr1d8lIoa3os7TadtTMcfYfWGjfAgs5k3DyejzZ8MBQMkp
bNRKYdNViCTpLkLlY1o2XLgspyAhkwDfFk+svuZX0wSp5UmaWe80FFoA3/uTWQpI
hNjq/cNmsesv9K2SMCdzxXJpIMqL6PPzqPRCCrvM9UEpRlzDajZgOk5l2eMnrhuq
gz0Vq+aFIyOeRkDoxohpmKrzUX1fTDgPF5WL2yE0VQJ27moiX9m5hjj6YXNjxBiT
InbF/ryBqZ1JCOedR6EiupIfEZgKvuL8/p8JZHUuqFC2KoMCTyjRwsYktww4bBNU
M6lO+ArKM1dZ/iq6LxG0uL0Akni5i1fPt6cZ7ag33Plryt1RfBdEghRzGw+UT/pl
2R5LXHdfZDThgyAmj4/YwhxeL/fuxK8TJeOLCq54rZFR8qlyvwiiXgNZeSSR2vDA
iQufCyz0tI1YK6HUgymq7YzUYT1BBa9c0QqCp+P0yjzRf+3jqpYlG+zIuNid8GQq
PYNMsj9IOH+ovRC0fzr/9u3bsUkaXhXSUMlIM+X2VrfsFbArNSdFmyxKRtYKGXd8
7jCJQqcPj08OhwrwoE5viumZszO6naYkGeNEpsA7VsmyEjSnfnVZvZflgsswHFoQ
4poVISrOXpDxn549QQhsy0F6fw0LZQZYcQCcpqgaJWmd6iBT9CY7Yp0BWesmSDTj
sM3n+9jQXT7r+ujPZi8RpIIzEPo5Zio/Nn4RuUkCDDunko+xaw3H2O8nxhmcHQGr
1/O/KmIHoKWzvrM7wcWgNzTo7DCiebqLjoYpgNpKvzq2IlstlUbDfuUwm7juj85S
dimXxIHvci4rCKjvDbh9MA+r/C/XRRG+7kd8Gj4Ep1B7vo8bZy0W4aUdsIaZIjnE
7/D0ESTE5YXbej8VUjujLA+YXS0mwVTKq2t9YOx99rtups7Z5PcH4yKazIFIIZZR
+2hnO6z/j0ykx2fJ2QGeW0bo1OvXTEjDUpcTaXBKjSiwXSfTchs+8T9f3pCdCO4h
+Ol8YXkkXrhRhK/B5BbgNlnnxOl9fL463UqUPz2bVGpycLWsRRRHvS5mLErYWalg
Tcl3f+vSxqGgRD1vw6Wli3wOMy3ObpzeVrB7BbjEDKbuoVB+2+JtJsMlAdrZjVSJ
BeO6U8v0yqpy+E81jNznNqrAfLy9jwbcIoYQCEJ0T5Pt2C95J//ihLoTiF0C8SK2
cP7P5vvrTFPaWEFd7mLn9J3RFqp3gC8e+Pz6UTI4XFOLyWJuVe0O9YAbLfWuWhes
kZo92j2oAbwea0TpuNDGtz/R0v7u5XPJlq2k+J5ZnjLzLI1oBXWxE7Rp/zzNHtHU
klMZ102BSbc8acJyhZw+mmRIR+rbC73o08l/00RfztNLCRoEGBsGKPxsmsS4rfnD
S50z7c+uSRENLZCG7jO6g+uQLGmmXe9rEFVMMMogLcFaFvmB/YJb8epHuZa5SVBj
vnHskf8bH941Wil02ihiDrDZz+JngWZScDOv61Et78fxrXVX513Z7bqmgI/6oBqc
dv6gOjPWdPy45rANTciM/5w6juJ6BsiwsZnwbPpJWvBnePPM/Ebs2KCOjfzeRl3Z
93Txhsur30ffQpvapKlKLP6z84TNWg/cgTHdnSJ/v0+v8JfcZN9RD04MGzP5XmcE
Uw3LeGzDPOzo/HsMGRvu2Ut3CijntLX8mE9QbKIR8PeQl1BgO9QsD6jsakA7d0Pw
jxJI7+l0zMP7bUM1BeFl1apd67WaTr9aeiODeZ45NDlCr2knkBoq83c4J+4XryaB
FpZQVA1xzCLPtNqDv1QWL5DwXH9rDp6nD31kkEMlkDgtAg3Q4HVHbZ8Tq6YSmNDN
1v3TnJ+SlvHFXb6N3k8cW5QBl/ebVEfi9oj/l+Q7XNrGODc+wCjC/mKh8KHkrkgg
pNmRBXlp7o0aKvzumGhhXDtf1m1OuQLvLM6HCjhTJmX9JwijMdtnLsS3moYtKSvm
fS3MOGV3OFtRe4sC2fcdSz7BP2qqvxqQx9cC3W7JnfPezFtqP9uGG1nBJMFrHD1k
rtocLuZFDx8cPQqt0wLd8hCGzrLiQ39bKLH/1JspG5O6hoNXfGImAqRQVCuUtIrd
Fo9TFFoYZAeNOsW3eoihmx5mHMTTI7xkNGxZIOofz3gJKYuMhrEU1Wh3h3c+YWC7
Hv2wFUX0KxNGdlpoje6V6vGr7rOoivf0WPdBBLAZqKmBKmaPjzGrli4DAKSleJXa
2lNxHUyVcjYDXGfVec4z9503FgNFc9+RTtb8FxxJ53bL8LYhLxK90fm3XvpgEeEB
vKLksFd8QEzZZ8wHz/22orH9g/nyJus8vjjMqrBKTlj6qBnFzXGxcvNMMgnPZnev
U0yxkxh7wa5jOwT/Dai+nb2ph7/xqcCP9OqeAbDSyJ0hnrQJ2+AMUPl2MIgGkkdw
Iro870IwETbEA6uJGfFHLhzkV1PtxErmIBCCdEGFv49zcgBKxZtERHveFVaWzUZ6
gYZiGnYaBwuBi8B1MmYN+rrTQ/YD1MULjMh4ssUJhbAc9Au0eZvN2ZXi8rPXXCp/
E4g/5jWsL1M0n2kfi/bmGRpkSUQiE6eF0LG3x4cCooG+NPDXi4wYUvfNUB+NF3Ys
PZRssEjS1hftYEbfNfR+/oYkC8Ut25M8VsRkRtLGlC+cQwL+dCc4ULXpSRKSBmX9
ucM7O05+byzzLax7l/GWzDpyk1GYYQ4/yzGc4JgpW05PdmSFfpK0PrjNhz75ESwW
1JovpTKiqitdD7ZY/++y0MtUeN6rrVGUI9rJJvM9asCBfVH3/B/zV97z511pyHd0
qs4Ygg8Nia5JUfpgmXmCjX+a5AwrBghOisWxUAWIvP2cW0ptSEBjRhiqseQYRgdP
EeiFUg3s7A+/S7BVkMOU393A3DGccx1FR0naxEnZNP6/abeiW/7ZWn/GLF2gBhAJ
pzB8Er25SSnacKTvVrgsJSFKPwsOjM5dbiwY/lnYR9uARKNRGc+pWp8Hdhkh8WBK
SW/bkUn7GFgzQgzzyJEYhBv9gI0pIEg7+H32htdB597ON+Tf972QXE+AMZ3F63NC
73ESwrR3m7LLQCAqvXrgd5nxmJwZT19En930vwedqnmJ3utuIEcqVkUo10u/fKpS
F4MvdGkR4Tk0qrr2nWflL2pDPwGy5r6mFCaGinKFQe8m/6wBBxHlpvFvlzQkb/hN
ojYOEtymQFw7B9HYb9jBIwO2dJtAanBHbE2VPYEMypvbGfz9uvdRErR+48pZilnA
kH9Mx6vx2jP8jDf9rErnXG6Km0oTd8bJ8L5RFZjpJzqIkGO80gEfnb0YhVN6F/xf
JO40pTyz8bR5EMaRh4craIccp90esSlBe1zwG2wthoyQH5OEf0En61Xgim+5ldPS
zhbPGx30yJD0G03Dx0qmIq5EIgzzwZB5x95e0Irryk/afX4EtELdahGR6gHGW7dx
NW43GCaIcEWPVQ39zAYfG6tnN7xOvJm6gF2VeGXoTKY92x6s1vdD0WgYf71d1gdW
TIxZPQEiRytmnunEffCn6lnbjW0r1LZoYN4oiA/yamSED+3XLSxU8I8SXNXP3snP
LnWkyJuJO6arv/a20lzK0q2jENp1d21nKBj9eKESax8Wl17cbYJuPKnQ9aC2x1xB
tIB1MoJ4PV2Cp6GnTyS1k77bzSTHgrDi/qD7UzMaYnChSb0NO8kHOnKOJ1oie587
TombZhD0fdN/Ac+mzcWz2kdwCrV0ox7FyZazyCu2A8J4fBqQJw7QIvvLgsX7AkqX
Mt7GuAxSMBNiPmXVoZDjAADFTCLsnhnyoepHwtuuxlfpSB9+prGu3yfw6BipJV3b
SAxcpQiBnxvXijYml4rY1p7HXniM1bYa8CFFtke5frBcr07aAhQs3qMMpwoBhGZ9
u2tBPqjakE7P/GbIgxB/UX+uRrL7p9n+z1hcifbZnhGY/u0/bKhM9L5HzBK1o3Ee
DSaeRsIgimwi1Klhojb8GR8/aMUvm9ijfxsdBkIUj5wsDdMbwK5J1DkbdcKmjjKz
2Wv7Lr9I5JNbidhL/TENKU8s83MgBiFcoZ3952kqO0cdSmGkirgounNpXHNts0Qx
l0KSoq3KLs3xtBb2TmvfpuR2kV9Ri7owhUY+Ivtai/jAubTIyWyyvSdaVXZns8Zq
cAT3AxRMGcKtLpF5/JJlFOBEsvvD729TltebHiI7hzkPtfAR7uydr4ZrXw4fSlgN
RZkxF87gn27ENhrpavHIG5b7VEjHsrnusRtvxPTUsb45i0UL/ZSZcY+GtMgDBzOE
rRL4Ru81UeqGx+BrUiXCnfrzdaubU5zjllCrQ110Js1JH//qOY252vANtPBlH0RY
+PmthiWZ1iN7MPTv1BsVGWRXwedlTG2mV85aBozJjQfRsDtk8/qXXXcmzSgzjzG7
HWXkZr55iWpbig/hQimOzVF7m21fIyMPbZuJLnDafeG3gtdRFtEQ2bLPiH5VomiQ
U8YetXhxe5E1/X1S8w0XvL5q7W58fssXPxJHY53AhwD9eGHLhCiM02kgtliKxVCb
/Moz0dLTnhbAGkhXQ/71vSSG3EMxAAy7NnQaRn5lcz9cvbtWeC3vYJFq4D5/ITrs
bBneIrfE18yx0ft0UnRtGqnTUPGHAm5uH1uwign0syxgAkPpcXya4iJzR3mF2JxB
9vhDn6l2YeKxF7/BipzAK0AzrIt4eFHoIvMIxSRjw8hy4zPnccA6Ga1MjLsiICKI
PjT9MvTV6eMM/6N4aGEG95z0vsEwh7jTHDY19VwHxv9qiXzEgMdOcAS27l2l4yRF
K6HMAGvh83Y2/VUtYG+ZLftMR6n54EvqsAmj4jR9BLb9J1Li0LGaJBtkoJJ4B/3J
uNK3qmbYNvVo7ZWiOHvYjDjrbqzyfqCqzuMZ1vKUQcY6/ctteMTHeHMwhcQFH0KI
B+CKK5qLmZTNtCvIBeJNf8LNiYiz7pNFYvv4FS00SlBrPVh+NJjYpmT5xzK2YQci
DrIVBp4d5VAYCf0TdKxcGsuXl9B1YUYaKBYPLCFxr+QcsBZhKd5m+IIMm+P2vQAN
ZPKU/4xhrpc+Hi2lvvkF9VXbVuRJKlGvvmJ1NcQmo4l4QFCCiAof9jVi160LYPvH
moXMhrS8L80NzzmfkEeNpjubVb94TPDaiWOEtN9bIDX4Vorou50EmHS0Qt/Tg4+s
JnulHSL3NqcSG0dEWl8kKyLorWMMCSbk5YUEqFmFyel4qmVBFklQLqu8YEUcHorv
Oelo4bzYJeojoBY8pqXhysQnybruJ7RxNfdxZ6SIMUOHrnK6WoAmrLIyGAyZ2Gbc
z1K3YShYRySzT5HMS0CXtqi/g3ung+qFU0jfBkuOaXBwcGfrfZtXRoUdAtX+WX8J
46bPvHpOpneggO+vdR1xuEmkcPc1Auee3z/AcWkrMI7GDpRo5JarHW63Tmbh+g/X
o03RgKP4zeaqi65n/neZoGhr5o+VreQW9r5gg2EtoM//4j8izygFam0lJO5itZr4
imJJx3HhhXhzYTKaQSS/GsBCR7DlMIKb7JijgXmxZ6rLSYFf5YYI2HW2oQBUpavQ
z2E4+G87TE652SNlVp3BZKfqTAgIL3UeuGCKxLtYEQAjzWJit8eHU6zdI4nFEg56
YjeKP+bbSp5qSm5hzJptLhwEEtR0zi7jNQ98vdR3fvRqz/pGfNWWvRMBc/mnAfHp
wMVA+ok3Wi5xHzAsGYxnIZjBW3QchNUTkN+yc/ifsTdPdGkzOZZ0QXqyVCgSdro/
nphBAmqefWdphCzy7yVy9GeXHOuz1BwAB/SN7N6x9Qga5gmHf6tYkyW2TdkoYLV5
J7omdQL5pjP3g7IyvBjpk8qFWiCE0zsuTCJfo3W3MkSBqNXwot5kRlQNlBKvuIE3
3UP+WuQDmioFP+s6XfTH5LTG4eiuGgInJSn8g5NWGJNil4R5lVnddt9MYrJuPhN5
6rERARAROy+4aFU1GVadD4Ee44YtIFbY+WRYQNUuLx7kJ9bNhf+d6BS5alTLsx53
V5Vp9XzCe8Bm5MFA54JP6Eswk0gUGHpusD7VUwW/JDQDP/w0696XkW0A2CGtJu4a
XOMl2iD9nH7mvLk9fVaAzM/BINycfJwzp2TQP0neo6vFksALjzpgJWvMhinV11Jo
xxerwxa0W3czXYjNGTiMvR9OM37DJQ+UGNRXu794onWrevs42f7d4/Aco7Tm+kb8
Shx+6RBicQmCf8g08ZtqxnJwvnqY7yvS6/AseCI3ptsuCfhq6DnUjoKbJaL1Mqck
fgars4lDCTKa0Qmrn5bIipUMHsdj/oBTsOYN8UmJpNvqt6+Knq4xFJuPtgBfgcJy
VfCYRVsiu3WWH+WB+zdiYOro1ECKPaCdQhueD/9E3Am1RPGnNncPySq0VbUAPHo2
Mzn1EeF0mpH+LtDTlz+h9eeemZCwPZ9MfzJB5aRyRACPnTKJDiToXadP87OknEg9
AztZ4w9V5qEPrRLlHV6mtfo7XWHGc5FPpFWYi8/fxfoJxhXIdosxa2BFlkv0Kyh/
gfmDNViDi4/Xj0Vfow5J0Px4gJlnEaZGHWf0lpzuXE98QbW0tB6qIXMVlJe+5vt5
/J2MwNqHCCg17Pn1CaGZjCtV3oJG+DXFom9h52+mDuyenf6l1QjPEJo4GTyPNuyp
t/1jfyEqfMNFGj73H+dEj5viFTygvsBWTqFKnTcWw4IxoTqhVi161tZPsMIOf4Fj
K5rV/TKzFoFv//DrzLfdDIywK3e5kFYtGKAubAEpVXO7+Zc9bnrqi2EcOBAVIoBJ
3J8/QbAgbHxGEuKYyzUgfJsOgyNEnxdYzt4eTHA5UEBmC0cjMGLVmQaerizcgVWi
G3BS/HMM6FdBggq0PAxLBxk1sbkkj5HOu7kXeBGhCEQSp2mTvvyS97pePCnrsyT8
B/DsxARYKAgpp0iuE9WS0NhJdwDuvH9kDp5KfZW48IZb3NgAW2N3f2W8/TelBpz9
AhvIEGgUtNn/5/iHWvtoID+Tu9GcGGveWPp1pVN3dczmkvcY/MYwHSmyIk4Eqr2y
`protect end_protected