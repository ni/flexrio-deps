`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23952 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aYEGshOCBNLOAFPz/YVL0JBlYK501538q4n5LbYg8NYY
flB1IfPO2fNtbKgT+SOHHRb97TYj+4U9y+XOtPTgSn9pj6+7OCCldju3wYwxVxe5
+VKUj9ToOZTnRv8AMGOpd1suz9kw2NLHpLgaPIMbC4O7ZEQj08XCf+Fs6JlXIQ5y
x2wF3CrKYEGTsGe5QrJgS98X6b2H5WtMDpnL+D/WasJ5hM7c5isSGeP7LmPqIl7a
Qcqn3AEa+BgW7EtYUOKP+GJzNvAuxVnqKjCoIrqXgj2Yil1oS5SbYBwG3DsGsUyU
NhgVRFe8xmVGYOBwo7+BW2TBtlkVPdbyUCGi2seMxUWgtNZWnmc3vyvwqU87g7vC
t06jH36pOr2emxQ5VJuiyPV+gL5FB+E3RidOppmr0s3Owozm9ThD2Baxx2fokhvS
hr01XrQE/QtcmEY1LvWe4RWCTOwd0EcOx3aQ552ryiHthdAZmcvzEAu5AWV4QLnj
5pZONCVB6r9hhOQgvbbcbzkZlSDw2eqWivrWTEYlpLevYBTL5YyFfafblDroUkhA
BsWA+7cWlUlYpsAiNn65FCnffdo4JMWf64YGChpDUY0/rx15NcMUSbQ27+PKK6oh
+GdKnnEH9JqqT6bTNRNKKBWdI3E4awth39nYLKA3TGkUlQaGxCgzjK2MeepBG2sP
/UOCSxIu7qQPjf+IPBJV8WcU2Kpc04SNacZ9vx+cZpzh6vVOwdFt9tIhXQWC9zxO
wg1eUoFkLsyycV2OsNOdZ0a26svWvqhROQFb3AMPaE6Vy/YyhXiEGWZrgY0uQ//n
xHZKavqsXYXQICwyPl1/TQlMtOouShNvoRQG9YGDinALVxYVBrefBeKEYLCPyMGf
RY97476YPd2RwSNx9t/AhrZtdQlXpLyLGThEU9GMKt5RawkrIer7aO1Oq3t5Zue9
Gnq6ruM4SnClgjAtIONj44Yr2NuqzEP5dvNFrGbWAwi18Fae4JWR/ZS1+pszjMJF
HKn7HektXhiICKU18Q8uw3RfFxRKqyFaxAM5W//nCRuNcvezgN2ympQUS1NVDegu
lhm6kgQlUh5m17PMO3B5WXBp3hmhUiWPs0HG8w4kYJ2g7SLyLVkF+4DIS+DBcFyD
TIBYMXwFVsKcUGxU0HWndy8asiUWbm17jqqyXYrJ3WDsO9CkQBHAtzJGS8QIyCAz
tLRjxkp8KqHaV7GUEKDO97VPy8oMvChJ9TG4qeIuGhp9DA7p7VUXJgfrVCVNEiiO
DxGZoioq2gzePvFRVn8eM0A5/gO0iHQfECd1eRF7Z02YYJjmchAlPlOYOPQcncew
LIIkhcR0EAW5Ti00NENeWDaORYQfUcfooDorngTqpm20XfrWRNrYL9l1ZwqTopyO
o866tywWnZDAVQDNaBl8rhHgsDXIHBnGYz7Ot0vPT26RIn6SRhG9Xc8iX07YfizS
YO34sAS/M7dJ8aGP1SWmeYpl+yM9G8NWOVivg5C+dPYFYZXjGx7xlb+ilDkCa6SP
5Rjj3WWLDGF10jIbmL0a1VEpgB88VK946PxscSiSfyVZnssrn57WAIou02ViFl6S
ru/D6ij2Yth/QRZ0j+U4XW2dixBI7TDYf2R4PwdOjIIqBMINdt0XEUBzwU/kkA0Q
8QTYY/SHqehTrU4NKPe7n94uv7mAKbshiiJEe8XkkSlgsgpnGM4YZSkgilAU0muy
C6zG1n4d3+HdjYviDdghlnCalmxahtROuCtmpFaOUB+xC0k2n8RMKs6nGc/0ALpo
klyLkA46hrrKSe7TL/vBghE+UUtQu5sib9rxmyhTe86BpxSlUjeAUCj3SLHnncdt
fps6W6aZ+m7SmcuDrxDrvczSdEFQbhxiLUvVm0DxC/pVKPtrGjBKRL7Wyulz8q/y
Mh/v4rxD469q58mTrmzoRrsM+D7vfhGkgRCgE2hc1Dv3wF5wz5MKlq52y3mLmCYf
yF/a3OVyK426Zecfou4mSz52r3zDJ2H50RFClLkiovXqjGzA5xLt9cNTOZVBiLm9
Z42SLpxDCvvoo3MJppQniBlXzCQBFPrPxtlC9bllkXLz58zHK4sIcLDbwJI5W2Dk
S+ryIkbS0PooC89RnDIPqiZMTVZ/syn+1foPES+C+ZXvX2GW6YwibIy3dPzErXvC
Sfs90k9yhROKnLmM0g+w2RKuZ+i6lm2GAQHrdaHJ7l/Y17gXgZr4aajw6AHbF8Yn
z1gGAlHgPD3fA+3l8YmxPROf8LEgo16ZJlzfX3wCzsJBTdPkW1+GFhzar0/NbPlN
HCQ4MHUtsJ/eJgYdD/vqIyh7AocbKYlItZNKhnnrHaWYv47l6gSuo5UXEHvwOzih
D5/aIybIacEr8MQa2ZSG+RW5PlRYYQa/EkpM5KGU0PeImGIxBfxZhRwXQ9OFIX1K
N0SK2c7a5VNwuB8ezDYl6ZO6jzIR9rDwpoaGniEvsC0cNtbBDf8DQCd+4IxYOoNc
q+95c9Xhi6eTezb/v0ulRfax0zKaJK0fp3ADI6TTx8wY+m8pH5iVWmDUGmNTwRyk
RgDISzWAkV404IW8LWLlw+4NLmfODSHcak9mVe51NI7cwLTai533DzlPR9eKZhMi
MaMtEOfB/k5FEQleuvAAiNNjjsdNg63KQXf/87lnLguxYLZWQ3zwldTucX1IQx2B
dK+WqLu+4Rq+TLt/MA+LVIOtN3JxyT5YM2uGWykAIICRi5nivj9X0Arxdfxqp3Ld
Hh5QnI99C8hQMCpFQyY3C+4nPuyxcaD/98zx2rOJVIMZLYfwId5WcsztoEJ15h7p
+LCTvZxXf+bTkThIRzLW0GFowWwGE91g5xXn+4zh3HuUyfeC7rcBmx8ejApsXrfZ
fMXftD4+UP1wVyyC3xjFDZFxhi9RVe5bFNZEqcjyGk4hT2lDHiX0Qx0oPZvfN6vY
Ixbg9mGq1I2KEFLJiQ9KGllUGBi4CAe9sawqaLW7ml4QPbG3oxng2FHKuMv0/T4Q
lItwc4seVKOWONqBsvDIwqhrVLTbHtoFgXkz0zVRVryIZPeOmAFElmmiy4bok92L
vitKUdFd0WWv8Qo0m8SPxd+IOfpXZaeffGW9UgUn6Y7uWLIRr5OPLRKHeVTrCkzZ
m83rCvNkcgqc0ZuQM3AaG0qB+E2lM8JbRxXNPCw1l1GG46qEfyFRopr8fFv/nEE6
qYyRTay7HunF9QWgM2q9V/3dIK/OTWti7Vp+AdVMwipT8Xk85IXu2YQeRkSVoWIr
PEyTALU7ClqKGLEP2h1LVMF5aL0jw6Gz9oYGeT8kzv/vQxfvc1YqVs4iskdJe4WC
0RPhm1WtPfV7yCDF0wxJ2lMNGcnCe+hwwq1t8fuJWXvpv5IXtSBnUtC0GHB6TtIL
5AP+iRJyfOcI3AemfjTfVFdd8okqyuR1Gr5nhprHfJEh2jLzW9kftJyQCRL3LeMO
tZxpbSvCthb1sHU1kUXy/xwh0C/XTscVNPUjvXACeUyDKFG2hvwkM+LXB0Ffz2f+
Yo+7KE/6gSaqmyCCK0ZQuj0zEDKw1htD892qPdmuOswHFoOcZVWWXe3NgXooZOx4
BXJNkIYGF01asL4NwsWOalJ3oZLj55JYBqP5kZZxSNUDSKZcJLbTJvHCHfe7lp4q
O65xhZW5jNEYXJ5onVDznHGnTCXIuktZhhIYK0YS74orjKoXPWTAIW7SB30/uktd
y6cHQAlRG4MbqUHCkawhR17j3kOPx82P0OdXeXqj8eGf68lqBCNh3xQZHp2tv0X9
iL+OtxU40xvvRRIgRz0xW95l82zGApxThV+x5VBjSo+6ylkX+AgzICWTHUztAM8t
Bv/ygaF2FwSIWpwCki2rJGZSvTQJhvOV4p7amEQrZOTRtio+f7Upzk40TxxZPyrY
Z77oHFbs2o7tMgyia9v408ZKuabZFKAlnTSc5+yCoJYCmMGgvJ4nuen+GVovsPgr
aHEZkiFAIHcyNOSl5XQniGFa9xOIIuEs8ZxDGfrv516lAwwy2F15g1OV1vVdB//+
EKwAE67YW84TeOf9L01Jm2JbiKkaDeTKgbXp1zPgMgWYOt0k0qNtPM836ynIDNJs
dPcPSWXVtLo6c1jCOlRkT0epNCiT4cvu/JH9QOK46romKqODPrgwiuyarq5NwM7t
oTlFNcZANvopXmJg+zh0UjQ0OaYg/o8YunhdpJOKQstZDtfrRXZTg+I88CWnzuhg
/ZQunB3b8B+/uEd3tXw5qc/0+3/yF6mc46yTMdfQSW9ksJeF26cyGFkN3aA8Q+WY
st1T4bl1nFFF8oF7qeqJJkz/vy2YYbD3qT8s18MRy5qA22PcGMQQgityLlh8QQve
hPNApdLAeY5/nffF0ZNPkMJ2f1siipny3g1pkBMgPTzv+JhbRE3ZjjBde26AEkzK
g600hrOHiupxSxRNWLQV2o2Zj9jp5H0P3uoCTPuMJQrJri6QvzZc2YV0bOkesYJJ
mNeoe4hpcfF6FL2VnJc/6c82VUrQ0Ex2uEK6Hz3+XRMOZyhGI1Er6NmAq/tnlyvk
vqzW5YvG+SiMHLZcQS40r9nmKEyeOm1NpNWUSGrKBdQU2/T3lShBC4Fx8Xsx42gs
HYeKZjHqI5DL3bgSOhHv6S/rnsddYlUrm+gHZMg29JL0F+NGYwNfew1eIy2psdol
+IHf0zP/vu5nWvCk4jNNHH8w05mQl0S2PF8RKpE4wAKINXCuey+qDLpcCtSLK70O
3U2QTyBVaiRkWFEfNdJKMXVpQRjr3PK+qCGx/h7Yr8zycVPzjwhh88+roLU7omkb
Q4ek33K+c+i75jzN0f4B1QN+WJFHkpHpuOxawk6P8zmzNIbMJaSxCaVjoyMm/BXb
Pfu1Oy+/yz7/OVEf3boNrpxmDcukGGkoao9RS1KjVeQVMyufMDdmkiXJh7lVWHWI
ddMCzyiQZeHTr+LELISGLMTzoH1ei83EEtqPd52RW8jdoLjaZAfwN+cIrQHp6fki
Xdf+3Nl4I7NvOLwwHiXvIQn0Xw9Hy6dy44/ueZ+qdYpYUIXBLpU9GZmHnpZawxMp
OgMg9KPyRoD6fOJF1jKNbhks+hPYQZ04rmmKtcw/88iuMvPoT5qN5TyZBhsN+fRB
HS9hj3HNRFpjVng0JkDlZTz3q/DbmGeizPYmdimUwJe0vzcEw1S005okDSxXPxvS
pV+M1OsZ2byKAljKKyna9uGWToWYD0CHAx4JYt59h3Uu5/dKKSWLD5tAMmFWYso2
Fe9ohLPlzPc5QrZWfn3yfBoLcZsBr7RpbwBTuY6kDpHCwNCiHp9LUsIETgc8Gzbb
TNMb5LdMHQU4wbZwL3KeQQq+KLcYhOja6QLtESNpEhKyUmm7UGfTn8zPGnT1PL0P
8tccmZYdkFT9V6wMR9BGAV14zWqWJkrpwxlltQP8gdFCJTeZAJH6EgcwE5AcWXsh
w7mowJ7/xw+SJXtAm4FuJqMBjEHMFm+rKhXvFvK6CxzctNZhe3gjLJASWlioxvCF
/ueB6j+t8YUeMqRDpdCzH3CxYUCcrpGzBJWCBcsSOsl3iyniOU3yu19H2UrznU2k
4Y34H0lOB9OMKSurQ+itK65LZ9Wwbs0gfzySo1m+IAoK91VWMS5zVLnMxiardcgY
C1aGqlK2re3W9zOJXkSrr4i+Pqu7FG6RNBQ8te9Y+jR25cMUW7lfvmNXRZ8eZYS+
D3AYIiRNfrF0NKSjqXAWrF7nvl8PbEaUUgzUDyG1KuYu2c4YlY26WwsOKVevoH2H
kANFgRm6BS0XlQEM5pON72NF6IeaX+Zd+2OJRszszkYHdla4vNmeLEk4J0XzD/X5
ErZwXgjjCKdSqlyic/VUIckTN344fEzo9AiuSgxsA69LZFHsTpgxsrcnLxFLe/hC
mxJirjFpuVPc6O0vCjih+xVS8dQo33sg9rDg0V2TRGYVJq4CFCVEVz4iWbZw2MlE
NhWWQk6grdEWmuWJJr+647Mnd97cdnqckca15hixXAsS3c6tQLVGqa3Mio8uaaEQ
+j2aPDm5uvtiKg5cm414JBbqz79yC+WVuKuO5kf21SZgTS/Fd0Vo0IyfCuO2QeJ3
J8BIR6tOekWvFAWqARR/l6+LgxK5BJti2/n8LMzYs2SrF7S+3lZj0wAPuMwYIQUs
TMie2/cCipwgLwP9EPPQ2Yokc/6mHu5ThGXPQfb0VKMLp9CkBNzhYdOEiMh21xhY
90snzaZbw97zPirKcMttgHkFQJ6xXnUC59iG0RaQWpMCOD+pYYuaW/IbAs4Fx/6g
hiSFGkGV+1/a59JYlcaEwz5UVBOTYeG0YJOiI82db0aCMANTdf6hAjyGBuQwQv92
X+bs0Vr2syQyCqmPND/2aTyB2nrj5hHCT0Skuwqm06IFm8nED8ZdbvsU1PI169li
tH69bec+5OpEWzKfwNXbTV9zPsruVTiYgGc4lYzaQXRvikifqANBd9vWwfiWLqM2
CDf9TofMT6KMt2QoHBZ6KeU9c7RQlcUDAyg9IEqpHyq2OYSy/Bz8MeKut4hlvHys
8v6uFTqTJu1+NFV68N9sQ8e/7S6zk8ncWakvx7F3zWIN3mwnppW7sC7EWmux3mZg
O8X5PGfiac5YrFjA+bcP+DXyGAyK+f3SuL3ffQxKEljxxKbPcU7tEMbklxt83r9J
Uli0DaUFY4hZi92QEzD/D/24PNxVvb4Ow+TAYZnfMraAaovCtlULUkdX7eVfu2GT
fuBAaC0bKddjDSYYdfndyHlwWzR5vXex/7S2gMuEkIbkZXOBKyscCQC35vv1lPvZ
CBe6xhcNpnk6b3YwL0gnlOOPaJCcGIoiVCw/JZU1O7DJJyXSVkkw59RyNuUIwk4W
MKbD+9FOcaD79vuJ4MlCA6V7KSA6nXd45iIuFPE+5sXmj3/53vKj6euZPUxuh8rJ
OiFOByvIgyUjAeoPHlnKuL+W8eehwkbEzgHvWbFRb6SQmK8VcJyf01v6RojpM9H4
J6C2qAzoi6b8gG8iHRT81BMa1xh2sxskvfUAxPk9t8V+ztvxpH2RxVQZZhV0pOJQ
2XvT8iRqALoqfHgA4hgulUobJZh0F8Hf8H//HbCLn/Q/evTzRxiFEsTGs/1Rf9YK
NA9bh2kM+MOATmiXUVyzL0aWCOCoudXpkxU1OE2t6aAaFNitzJuzjE77U6TXK12r
UPHXGJ7MIvs5kWplh4jdtH32YlmIL2XMEfOiT9m3FDIYs4OrbXQrMnHnmwZfzJ30
kDaAt4JD6CK2FDlAtCkKvK2bdOgEArs6VKwGudZ8qhDQ1MuqP2GkGVp3szi3kjfG
G0sm0EC6g8mGsgcS9C24KpyvystDIq+x9RqcXAhOtKTyfqcxgZuCArlCmzQ7Auc3
ZPQJhAMxvzVGW8O1l8SvHU0cD4C6Hb4wHnzLKtwOQVFMZ/Camtt0DGP1jWE6kTb0
gmHPA8hraAlh6X8QZNzQWaYD/ntDFUkCgSXBE0bfacYCXeYoRqyiAgHmHpnqs9Kl
GW8QDPudcmmZ/085Eu+p/gCLF8PygPufBJVLGwaVRvJg870cgzUsRJhXuk17eNxX
bT2Q6kP5OKHVqEd/+h+9KDxS5MF/mWtqvO6zDg2hHtdMTR2S293ISMBp/D0WPxXC
eQ6uVzN2N06wif9RIU274I9voAHXaEPee9dL6uEVfmZlrw403LG7HU1xfCDuDx91
eK7SDE7Ipy2wV2brzhHjj6ZrinMQdNHlzdJGzymI0CR2uvVFw+ltVG4/ONrmr14h
ancqkqx6aQ8Fdy02ClANgIVH0FejvJ0RjqmpSHWDPHmJH7aCdXcLdaXQq6ff0xgl
PtxDxvLV6LbFxMQOJeXOiA/VbTasrjGjZHAlCRnG/Cvwr7ei7X9wSmQp3FXWrz/8
Bfu3H9A1GBBzDw7LM3dZ3+PoQuj2Hriaw/Xn9DNewm/jdnta6ACvESJphcCUrXhq
1xgO0J5ycmbvSkhK9H5CYLpOKehHIaAOm+j7MsXs5wMKs5TEy9BCaE4OVwrB3OuF
HX/0eTYh2KGANpjaqjfVAKSCRfyKXpxDhJuAx7t5c8VYRmvh0e6RJyYShLQQPX9a
AHYB3mHOymXb1uX4DUwgo3q9MB3FyVgf/6KdtE0HbmCNJS4lNsE65a9dwRZws6Zs
mIRgVq59ramilKQyqIJlLHD4oeZeGzaftXYzzk29NMJLiJFPTPRTRN0qJj2QcPHk
q9KOhafoVytFlSctvF07dWFUaii6Y0br+vt+Qb5iaw2+13ogwRwJw+i4z1WQ6ruV
OdBzqP67fLWeB3TuLsdon/kjSf/nVL/aKGOS1AnC37i/z/gj+he7kO9Ap34RIDqu
1p1FBmkPylivA+f6SNqR7SMHWIk0wCtqeQvio7si4k0yaLRXt3QJOKiuGsbhj+I9
/rSdQlbNN0VVPBg0/6S3JtNhsgZVsOFNR0YuxL49qgIZhxayZNMPllwsNILH19uw
5B1sNqYT3shdOF73MM/svdtXuew2FydfNWZ/WPmkvv5mzKvdLI+gAI9/+hMdRXwx
XDqNZq6DiDlzzhkiXUgi05ak21S+7qKJOVCdge9m4D4FZctspTRrevgxR28KRzuc
YderN6kTJnpKsM1mFrLEOn7o1cnIpNz/FNOBgpONsT20zfGr33SeXp4RlTloxIgX
lm44rExRumxOfffXlk2U1v/H2CaIb7iB9VgYvNsYJ54A0Vg6E180GfcgPHoUVzqc
6zQhR+zD8dpBy9frfDj9jlHLTWsasgn1+ICeNtMqNE/FybhEeow2iuqCsFBXMQU8
w2epbZjKYkZd8cAgnrxXQzNo7n6nXZcQ0jUXDQv2N+S78mo11zE4kw0xWkHHc3Ze
nne0fEvVZzedVbNKfIHYiCbt9dAgkZLD4RHGWZatFOGfDuz8kYBZxa27HDUwDeB1
aNbll058lJr3bKZ7n3/AmYz8CLExBcObhY6nXScvKk9OUZ2wpJ7ZwrnfArvUjD5B
zYdJigWalD0TbBOhbhfOl6qaLPupwnq9TGJvwwD7g5HVD8T7ywqHbtZLrpbYkYqu
HYvwzPgeRWcdkAZURwWLqinOP/78FQtQe1gOla/4V+m5tsiD2vxBfQkocgNG1Geu
LP5XAsJcFupRfa5d+Vk8Lqb8UTOHNz3J10ymS7/koStKXd1E9niHiLE8xWs5j1Dr
8jY/NWlxcRohOMqY2WVe3gJf6Ci/t3VjiaAqIYt2/jrvRe06UppXdjRxs36pfWAh
/MfkFA3ufDDtXBLW6+5hOJ99rW3PBLqSQ8Yl+Wctm9TZ7l6oG8JEUK+Iax8fwauP
1iknGTwmWv0RsFGtWITGjFzR7aY3RsUS+FOok9PnaxTpog2uV6DAEIVUoCn8lkku
Dprk+kLZQBZPUGaIVEnUD7PegS+X8SGfKmDjjREFCcJm5RP5aQC2Q0hrTtCPlAi/
Ba/CkM9ARx9eKFKDYysHSC1x3HtOOKxjYWYHVAvYYmPu/Uri1wrbbRRz2aVcFmYY
LbKz4H8zJ6W5U3FcBALCzuCaBSYCgNSWUeF94xQQj2aP9cVbX7aPhoys/TkxJUrN
Cw1yBVr/kLY9bSQ0NiVfg/UHcfWsjBpOzoV+604QjqSMoURZO6xNawubkATByX4G
A1srIQLFv2hiKSYInjy+skA5fErLE4bmGffTOKVdEaMoAUBx5iW3Md8BKdh01GmN
/aZwbHS7jDPoqEdSElfqhapQzEiJlEsc/mz8VElXlvBdAEep6PUU8utuWdLNk9Ok
SFQnNYjvWmmKfgpzr6pkAUw95Uj6t/0G7syTs4nLW3/6su3+w3bDSvD0dLIPjB0F
MU8Ivk4H31tJ72uzd4yyWJm7DEYXGKhDttaWaOHWW11Q0bK7eIt2gnnCwrdXJ4Of
m0vBq/mJ1KFiu6IyP4BWYJ/ihDR7oxzMz/0F3WX5xi4lm29vTozJOJIrswvfYPaJ
Viq4LuJFu04A3mYJBwz6PCgREXKpR1oy6tqrcJ6oAZqARTiQQz1MLwrJUgKtezFv
QKfxgNEuIZ1FvW73lBlmEaisOlGPSdmxm0luwxdlxNRk4EhPhOmuyjrXm/s2+1/x
EVabHwNV+FbNRqWoyaYiZpTM5zspbBXHmelGWX7RatWQVFNDs3hIq4o6c33TlRyh
4VkPNIo4cgi7rkNIe/9jBqIjFEhtngBsVcqx/aYUpbvYME5TuTW9csZE6aDbV5a/
X+yBCl425DFfWoGMvSVeAbCnPKf0CoViZRe41LTwKxtRrTBpjngqQ7helg3CF4dq
T5RM2+iOFaSQFXWCHaUoLxX0RfxUe995J8bk3b+WWc6nOb2nwWjEkH0JfTP8AcpS
qZChjyIJGjGt9z7ZTDZjxMAAredB+0Uv2lU6frWHAn7WIVAKu7ZF/0n75bLmGGS+
zyiSqYTcXTI7XwuPz8TaALpRA5TRNIu37BJ9LiJxld8+AbE7bm4eZAVZZsq/lZMV
zX2Q9yFvufpETTQS9r3n2Po0u4XYdKLxkLLJPhSmaU6CZQ7/gInisOlZdQ/wMHOE
ZBaejIbx2EjOxc9EAC9Zw7bv6q39u3Cp854KvW4htig1bgpjfF8o6BDJGkwv6wD0
Dp8PtNWrmMrCLC5HFz4zSPo9OKNa1oW6AaUqNIb2qyNJgXlvUpSPgx/3IIwXwNPd
elUvreYQcMKHB2D1xgQQkal6vcv745T81VUgpnQFXgei8WaBioJsjMgs6CbrB+mb
XS7gsx+j2VKHhYQJBFtY9aClow4ViYnD0JLp1mGfW8DblsQeBiwPpuTItIeRpxoK
SKd1DxCoW5aWccN+dvVqNnbRFfEeZxgSrEqGaRTpZvn1/AhJuOVJ728m9/NDDBSV
npDmko4maIa+wrWaIqUlUYAY7ARq7QPMWdR9Uq0obf8lXzx8xvT73BuRqyO0rldK
i7xtCugfMH4K2EM0g1fpK0UqwEGf6zT3rmqF7D844JONm6p6BGv8YlV4bCW4ah6u
hMOX44D2ZMuXXoA3wxVJBX93sZF1d5KnVf84NJugq/imL9B1HXtDp8iC+DBVWo78
v5Qez1wjTXppohTyQzkLbUjEvUnDe+sQ/0LIlc7T6ex9wpV3Jjn1is2Ec69pdonw
f1YqpsHgLRhUvNriMyUmkJFNLomX/i74mB2/328XovPnQ5ron/ugUAO8y1QKgl4F
wUxPvBrBedNNLANQ/CPHO0GnQylMlehmtMvkGeXpFws3j3bbFToXaiGre8rhUEpw
fd4VzrLG7KsMCmZHSmXOzdfb/eTOCwb3BOFOd1IBOfMoNIKRq1xaiNuVHaiKtj3Q
zPkmN63iD5CLdtBVMeYMKgTlRhHEdBq2/vO0D1zqTji/hSyhILuh4Ryn5ehwZVnq
jAJ/qFvb1UznkNuokHPdawO+ECQef7bAIDJLVMxYR5u33m5Bv/H3aE60jcxOUqWd
C0rtstsS/mHXNHe5eREg53Ftrs2S+nzVZSnMsCBe6uoBVa0vc7wwZNxE/Zw0kjNz
NeMPF8oF3jCrpIZ8p41D0q32PnSra5gE42bUGMnih89bnYeY8gmdDokPEKyy5VBi
dRV7JJbtyryM32g6KvC+IRWmB/uYTR0IeXCZkAWR0lrVq1VXZ9Epwd/AtEYbJyb4
AIcd5bwYMtOmMqUr9VeDuN36+mqIvxaFvQmh5iierFi5lxWQgrZYbTXqqYm4s9za
vJmfPmwB6bzCEavHUgBRa9WE/qhPBLXUObMSQNirhHbTjs7ZRjRdPZCqIpjwGDLV
/n7OQskwoQJNUUUPXmV3aAOpK5OGHwVUQB/CoQ49pW7NW550u5oogIz2CsKtHEdg
r4R/+7df0OBJgD/p+MZ1a+2YpF7SJHLJPcnoxcQo9qlFQiLbZKHNLZSUC+rySPPb
F8VaHzbtiOYJmoU7JqWmdjHyVvIguXS1OmPmPjERwyu5cDfA4yJtrqdJ96/YSkzA
FG9naQFhg2JtpUmIw1vkOGx1GNnjuZy9hN36Lpi6wwWMC5GTZ/xwUQl3QGfWzMf5
wV2nbAI/MC/u84I817Om2Q7kj1RuEulHLkBmwrJJpCR9cgj2aDeMiqLPWDVFPCgb
lnWmvIOf4OFxO582MfWK4BYL2GBzeY95JxsEey1QWR2LN0b7HFS9h9u7at4YdnjM
75ZVbtVoh2DmRynLYZZ5O4ZI/GzTHNmgfio1oij8BntFU3jd4d4jAV5e/pPpjtyE
n2Imf8B78EbQsqlMWEQnt4lm8RufLK6SkaS0uXKPvfsyJjfDXcu2xosIgVEW+LgW
/vjNRpKJF/8Y2uyYTRdbvHJzSQPcG0runb484jwtXNOgd3Hdtf94+KPUPUnHOc8W
Ide9kxLsoNbT77HqXCem5fyRdgdJLnBnVACON0o5T1skcNLRQdnWwJbHSSuCVIgp
zKjj1RvCg2ExY7EbktdeQKO+m5korT6llO8oSyZlo7cAwvkKErtRGnxOvFKb51Q2
snrIb5nw5e4tC11XdLiNiUdk0FOhnx7PbSUj+EyjoYDIDkxzkL3gLC0U29qXn1vr
GiPKGY51y9Yd29B4WAkV5p7yJpH+F4Z9N26v+CVvPZW0Xsf3WpNRr7y7dHI2uF55
bDPx8o1Yk4QKp/pG8m8ppxrn1zBaO+Gve62/xqkI4SNZCnkY+MZLyFI3oJ1D/7wA
bJg6XwAiu1Ruhq0ahHYBYu4A1iZkghdaKforp72orQ4eXpc0NUGUzhmji/8nEh96
WH7q2WOOtRofU1+TJfGuaLsRSEQ3J6OYkAJqFY27GUPr7m7GTv3u9Sxnz4y0yvjT
bKRLPm6MCUjtgNzTq5DMeY/Ca6m0ZGeL3OXzHQgtlu+vL+sPDeGI7P2Kb26ZU0qO
Kw4Dj601xObWLn0bjEoO9+22JxcLirOEmowsvP7ThVmqHaZrfBO0io8W2IL1qLc8
thOLqwQdiZfIsZ6pq7FDUGoX5W/OjS8Uqugs0OfZJH7t1J5WA5uP/M3x407la34i
h4MaKCwpTl7OzZhXT8u92V3Jw/b+yhkz3fmJ3GvspQw5RqOIZiW5aK/PWjHfA66t
JjkEUqvftB1Ou3s4gXY8/Ly3VCy1DYmFLU9Xb5RoA/BgmhAGzONINgfub5Pce0ex
XOKbq5gcCT3IigzOWQjvyQ04+cZRz088Q0/XcUk3cbEFrTxhD9e76cR24W7B/8rQ
c7WWItaWWXG3DpCHDwojDda0wyFKtsSusb1f21f49GI51wR1VJcp1pUEcvnHDNLC
xskg5k7Kv3nnWCSvliPRwaKExsJW4Rc21UxHucz2kzrl5mRA4FKZ1PvaqoD9K90e
xcILvf2toxi3AAQVu5iT+pcPcAcO3w1lZsE66pVPf9Yv8NiGoX1dqCDOFZTkP0rZ
xWusSdXW4C6t+ifVcskeDYy+uiZC8H70LoMPgMyQtMXdrOoTh8QE1fw0ZxX58Eyi
O6Cb/vqEP+yajqTwYEZfdppIBlrhnz75ZDEw5rYDC11/R+GCZSDQhUjzGN47nRFA
bP04fGXKhNSS5JOtCKhhDbGYdN928OLv2CpXWw2iL66YviT33T1NMAHgk6eHxooy
U6vYv2BcYy1aV1ZvFlsHdFBTVFe2mXg64HhLSD/ZAGPaZIrVxW7XIp1XkjXtX3fD
5sUG+9WCQoS2V1MBjg1NdQzFDaFuVwnjfxp7qJcrv5QtARpqg+BUnUpTm3ratBVZ
RBUXZsakLwPrQAadX8+KLPDaYtJAZfzw0gyeCJ0/tIcCqvbhF75eAKCaCmQ8ZwVm
e2UcOkoJCZdtiO+W1vrc77ILCbHco1HLOx5cKZ03MRWUL1fngBRpFGDmTAiJQ3kQ
e53pwco7r9FKr/P7jZFFoV6UAf8yMv+E7vUsoKrGcLT+/NvW7wpsCDpOsQIsNLBD
as/Hf0Rd+kU78APthj5hA0o9jPuoL4IDXgsIzyGpyKC0reH/2hlVkpSrq3h6E1NG
7QZjGXZWv0pfL+XHRL7rXogBYiGjAnO/NYzY2V0exP6Km9Eo42lJWiLWlUAii6P8
S95QUul/P2Ac5js/g+6soL2Vif03UXYiDOKmapC8NGME66Jp7b5QSaGwOOdxMs5H
OBAoSsdGsVJLSbIVwHI/wH04dKJdNZm2PvLqtvYLZp9vyeXvzVb4CaXcmVMcbrSZ
zJdSZURAUMoPomMQ7Vj4jS0ByLmUUhclp0sZ3UGUFfbRzDsmtSbpYqvZSEHjrxUi
HGnNJGk5iW5AzoVNiOuwsh9SlQA7sKK1UQJw5+7F1KUdD41U8CMBSMyJ/k6a9S41
1TvEIxUrr85jTxlW2Iajo7+6D5u8oofq0++VV8Pu+p9btVYiAwxC5ebe/2/A23rw
tjNlY838hYzNDRUW/HZB2zeSi6mNUGYQCQgUu6ImKQDul20bvEYbnPtzCLq14CTn
x9U82CaF3IDu/QyzOSWQowlS+a0uX4FQxCe9EU82S8KyBtwXnwvqENqWvg+CHgZn
Qm5JGJ7Sf2gEcK1LZRTZ9AlDZafH0G92hc3XYcpJanGdjd0hPxw66c7Rl0sIdNn7
ZHseHj/42yHXZbh92V08eMuIBfrPb0NqrfCwuP9evV4CeNMWwdkbS0POSBNZzvp4
EbYcFrA6F/jPm/aDJViEEJ7dgtx2fJGGW9PzTM+OT1QKrXLaeOj7858DBGYMQgmU
0zm1ir4E88P3uNGj7CQv7jP6Cvz0lD/d0XdBtpOuG4DCcNdPrO2xVtE6GSb54aIJ
z4TYLfWvahEm5YvAAnFreKg6LecFu0qnsX7T3lY3umpf32qaujKeeq1kq6x2Lk8F
Tu4BtuAOCf55/Ykt5Z0Bx6tEQOvA/Xg7JeW5EabIT+79KVQ9nNqRR5PQHtLlJOqw
HHxY/23O4RwKxmYr/o2HuYwGQqIL0rCt1Tdu4FxztNnUJD/Gn/3/dDPIZ0ZiOSMu
L4QK6pRBVoenzvOHwSWdkXYGkpb5r3jtrx+fEFJMRkyYim3KgxPDvBk85QwAGILa
Q9UqlqOgjqWriTtyKvhYCedJNuNTZPEtiPT3iuL4r/JVk6VbTFTawbBGiFgDA8sn
XnQLXxex/SKY9rWP6tL6+aiD1CJcXxv78IR//93UhP/gmrpArUKnwEDqXwin2ktV
CABczQcheEYs3z3ITo6vlLOIdB3yezeLrWAA1tUOJ6yYROEtcDw1L5bbwictjO7Q
3dFy2VEwgwTnxX5K4ry0ZtRObgoOodFZKj7nG12D6eJ+9cROXmzBowzyohI46bG+
jX/IG9Ts5pdG3GJ56UYszpJcpMEOpBwahY6lYmRowSYqpZZVz9KqIbVrA7s3EafO
BhJHx2SiYAWJUDs6xLLUAW5p47ri7UQFHEWxFrqjaw5AerxhbaPG8FA8cxZr9dxZ
20T45gNLJW8grzhKMudRPXPz4FFDXhIfVbgNH8x0bN6zAm34cVgU+Cp4dqFWtJH4
BjsodqBgq69rGU5V8GoKrEGnFgz0Dp8SmoPQaltGJnP9lKVeDF5fdYNNHNkWMWZp
5KWcJaJ9PAXfRRsF927xWBxj7WFxft7eyELnFN1zbE1Uv4txdwN7V8Lt/zeXNSQS
DwA9WDzfw+EkV6gu1fRpMHleI9BIWgxr3CSQlw9RXOxB7Vi+QyECgBb4BsemLGIG
9HOKd6362jL5Y4662pNTDABQ6sCxUtOzZ8GPtri5sMWJLCPLvmOuMxskDWGYYcRI
+uSGU2Odkxi7tuy4nHKpNaHDWMDEdN54OBFYD25ME+PzgkWaus5rQ0JMOQZl20v4
eYx5D9ICbnHrB/dtbV5GS8opYRmjBOlg4K2pCh/Bvvyo+2enwgFp3o0sWvgBSnfd
2hzT46/OmVjPo8Gr2wQsMQjZICXmf5VvkyJcNcaIsj/V67gCUG4A6S+GUeXUGqaz
9fqHmJNsXH/NN8yhKyoUsGCizqztLMGOPQq5o1HS7jhNXVLfKfmh0JrjVrLc96go
DXVfTKCgtPhIATYcvNcmXn2IMUGogCWUhSoi0Ueg3kcI/j3cyEYi1iY3xFpexD8O
wadE+pYalW85Dh/McCMgC/RSf53P6+O4dszFgDXu5VUX9NvmgrOIUL3IsxiTZsFe
dSpZQo7d3/xdsQhv3Q35ggdWz/pI3kZtt3bZJX+PpMDAoYuhxQvfcbp194S1Al8G
S5Z6uBDy1E2v8gItGR6vKI2oe7h+PW5dsJURmf0zEvCeRETu7QLx96oYIkgoj8if
6LxgLgrCQTADI/X585AlIv2/SpeDoy+CAGupOz0Zf/89pYugZA5FM+TVX4zPCZ8/
Xr7cm5uk+4ncAjLBULxBRsbv9CJt4xSZomG+GrEBiPpZDfV7KDwAt1IU3ohb0i25
qMN1ihi5oJOcm/u0Uo540tU6hUEGqJtl0KKMPpatkTg9In8jSluh5HiFTDLk17uA
scTt5xc7XMnlHVjjNcg1NL274Jam2/doZrCYo31em4zyF+9AitDegLbIp4tD/WCf
wNWzS4soYSbHp4MpOx8tkkBW2baqWGtGZNP9ewcX2G6VQq/x0Uk9agpmPRgswAEa
54o9UHu+NBtqjMOmZ3CIu/EyCffznknvORRjXd2iCb/CvMrTXIRVzGL0s1/EiT8S
RqKjBNOm0MTFCY985HGgPlc8D29mOZLRgi7N83IvGVSBCaxYnNFLxZvpK1mK3cjl
YH6hLCeAd2fnNyTkH3Cm/dRFMbxAXH1Q4eSpAqy0hueJr7RwjVHpTu6U6kOR6hr1
Sf8eL60EMqunjk4lArcVLLybB3TfsbTHNHS81RvFhyDm+2v+OZqLZmlivTWCw+sJ
Kr/Fy2pFp+StAs0Zgpgr+QxurggMayXvS2KfMPkXcn7/tI7ERw5txc3tMxyr7E6C
ChjSFw+rmI6Qa+zZvVRUpBT82HfHhp4POLiPXTFHOcLVOeS3r3rPVccY3LoUhDja
dDCml43UBSNwbQWkV8ADSjQVeQiQ4s8pE7eJCS/q+h7h6/EOSFsp27DCdWBWJn5Y
bWcPr/J0vCb39kw2904PwjuoLyFGnDP9e8BaAaQE5KHryMneDzDTYbFiU7McKWiW
sjzm4sEQeeZs+ii5c1pnqUPTAvCFHfOkbnRgCArEaxq2B0T82YMV6V+ydJlxNSxv
4aF+MZyLTW/oMYef3q0/G3nN8UbZBVc7PszvxnB/95VlF2jvLw9l8Y9YHVRt/Imm
Xq9WbPyVL2TuGRsqS9wDjm6x9pLJZneIvs5lRsR2BS7yFdcRGadMKgwzkui5N1R5
53A5C39dbagIyjQcruRDdsaDVhrDTueBq/OtqvBkpH6YuorW7/OOqqwPiUenvyv1
qufUSOESy4jON5mXiZIgZFFek9Yb9TtTbYgwWnQjxCzH7Z+y3fYSm04MKak+4yuV
df8UJK+QEYpSlHpJQFGO+4hpCzqbd/BeYl1NZwQJNArQQyRQ5KIkVAJv3KwKwnZC
yCnLaC4R2NeH2MsiSxF8Ij3hQD8yaADuWhS7nCMNkqRh7OdeKvHQ8YhwcfDtSKtp
tm5uqdazXAc/874W9KA5x1Ue+LTQZV9FA9sTbka7/l9s/8lIsisTKhMSncYdC8zx
zGDsqUskxLaAJQiPQvRzlWFdBmMOfcKr5byakNQ/gJOe9yMy4FgtmOL3xchq2i9B
j6Oq13roA5ZFPnnqqQyNevcLiV9iOHC9crWyYGe2gP8ChTiHWJX5hoqgD5VgPxAD
38SvIu2NBJbhx3BiIEx/NeQLkIz+CHVOss6ry1RlyRdHQ3Fm0NoKPIImOI8sRaS8
ivIvf0M/nqZwOcWNKDdDAdsS0d5Olyy5lyzW9G8l6fRld9TEjID5oF5MwT8it64G
3XIOlexwxpX5s+75guYjv6MhrHQYAKmj+Kd7wcHy3s6VeYpbc5l8rQcszoo7t7ag
XMadjWymzneLweJFPuN6oW36hJc2bYixnd02Ty8tKr1vbDFG11LGce9BvkyAvTzN
+lvVc9j3O6zaBTCkzHJ1X/SFkdmWZaJ1niRzgA9a3LAsw4bjgth3dNhrhDvSdZ86
UPgCOYI+XBINz5CIrHiGQ+Vmn9FODEgvko/GpaUZvH0cD7mhcMdZvL2jGZ3t63uq
l81dG05phfbyAJ91BKr9XbxzxyNdaxGP5cT3L/FihlZoMyrZrovRWUf/LJZnnZyi
jbvEitk+RxjxiK3ebnhYbKjIRUqMDVLh7dF+dC/dHZUI03sZAimOdqXQ9g/fsH1t
H8xn1L+1Mcfy0YmkJjkoYf98mj7vgj01Ko4MuAftJFi0xEvOPxJIdQNoA0YLS3jz
cWpCiN2byEzBTellEauGWtVMVUvC1Bbp3Mpl0Y5hMf1w1YjOMLmBaWEiAYnnjM8B
80WnKE0Js07y8RM37ZRbslay6ri/PyfZlWpQd96yFRbdqh57vRdCunYaDxqdut2E
w21HqzHIDmgDc5QTg99fTa/t7CZgd8Er8JMtrcnUmvZDyriuFiusbBRjTgiW6G1A
xYkD6Eznzg2M2DE97xr05OyM5gSMK3TtwvHwwu/2XGxnsOrpB6sNjBT2+alhVl22
x82wtnrPFODV2Tu1vDaEkpqhI1cP9jHIf3hTRRzSqg1IyJwqdvuTgricnxon4yzE
cuJsuodOTZlUQhzvmzeClwfEUtW82wwzgPr93jBGJVQdDixpBGqqIbjgQQLow4Wg
r370615EmhtOUrskDeraLtfAglXawQHP54JqkimoqsdvYbukS2K4kNTwrBgA15Ap
XLgFEweXbJHZrk0c/F8FTOZPaOOda+R9QSG3tITPSR2SJ+YsB4+sVu/exKixw75n
3Ie+R7D0tb7pHBYCtJbThNUDtWgftlUQC6K1Do0LV7kY20pU/hcb87NkcsQmYzR7
lRC5iviSbT1MipZcUTFTBboy4gBXyrXx6iKVJJ58dLLAA1yiTk9B4FfUFDYRMCEb
iAChmVBfjZLTt6SjeUM3x7zGiHiykdJ82ehRr1GgAuXtmMnthoGUldFkpdPZjphP
A83OpirMMYHzyoFqFEV4ShmvRvTicCRA9qplpSbHE5SXVl54Qz0PoWUBziCcCA1o
eK6XFh8PUN4znDzZJxI8u6TEV9+7BvPFtyNJrM7jNe8vka7s5NmlrNSxar3vO3Lh
2nldnFpVGHl9qTA6Dnl7SVEv+vNb9/UZTqvuEtpKI/rU+bUdq7jS5Smku0uMovFT
tV7Pc6x3rqIohyo+53wiOTvTsos92HOMZaX5VMchf2cefEzTYk8KStszg7Nii68f
s3l1xkkWpyB/k5IFDHUwauKZEERfjZqCDFtUod8qEFK8rbXLbezcxLpAzIUxfI1W
wk/ExyrBciCvGNxPwbLPxO1JnUZ0yqBy70HiX2CxHyC2nOLeZ83QpP5UWUCK1gCX
f659btXmelm2qDceeX8RlDPG6GXctTLEID8Z4n+be/+JUgMg6VjPxo2EOZqbRfPy
63QnxvyKd9ZjF+3VbIo8DUahIlfTVfs4Mm6Dpuu3giIX9HsdL6qlO/aaxPGw2BeM
XDzTao8o7K6zu5GZeMmVKJkwxuATbYSZJqrzAVfF8aS1gOEwL4WH1odV84wug3So
JpfNbs5qy4GuSvAytgv9j4paExl6TJ1lY6Yx5uMlinhUFYvPxVFmMUuAVhPDJK8d
aM/ZHbi/rA3rPCo2iD/as7bn3krLulbY28lxBliQJEiWwYyOcUshMyJVVy+t83/K
DNs/FAx8W3hkJBVcMX1VGU7Pq/mmaN53ODpN5QropDXwUR9dXF7rvMSDkkPFzbht
ivSDELatRLuqkShtg4JZ+aVtu/xdHEsWm8u3wY564ELwOES0henuFW1r4HUcvLpG
YlTVHWhn8VljPLz5t4UpO0QHTdN/f/OaChMLI+l4WT8BBAPYPJMaEOCUF4ogx33K
K0g61eQKr/VIoedsf0Hr/jRVknXxrD4D93wApZvP88vayLE0Iv77sEo783pK9YmW
kfV0Yr+04cC16hBNT9RcCdOC34oEIU97IiOA+jXGXBwe4z1xv6mq9rngfkKV2g4B
46vOHG33TspK35KbhZtkmRX2qmdIN9cg8HuKRBW3StDJVAfxiRRl5v0smMUkVBTn
jS+rpSzKh0D4WAh3FOQzZrT9ZZ+dl+T9HLQvd02HWo2WQLZHhr5rhZkhUD9be7yK
zpO7WfVW+F6cv3Zv6ZqXBgjdW6/PdZy3Y4VywupxLHGuPXGFEaieHvB98AOPX/06
YQbD+BtvVJ5TYnRiLqJp1Jyz0XKDocBj2ea+7AHV1LGKfrfgz5VgwtXmcGcBnyai
cSrEq4Yf4Rqa9U1CG0u7MxIJ2QwzSl9NesgI+/ewgpoxuIKkpXd7RqYi3HE7hxQz
mJdr2eX5iGRYYUoJRy+0LSyEabjB4Meoi+iaU9ciWajkdemc88KstWtRa8jc+6GN
We0NbvS0gnlJ40TzCBFSoK4xEJX6USxPHyVSMiTFw/kCOxobfeYU7uWT9Y7aY9yf
XnPIanwZyxoWdM6+wNhP8O9F1O9zyW3fHBwSLjCXh05eriFJ8Wvsa3LAlGe/eYs4
MJzZrYbEvB0WEKs4siwx7jbldrKkVJZwqpgHxMxRQ9j9FD4cG39ctVoHX+mZcMGf
Sbwme99BOAyYmzSu+BMjDYi/7hwgbiMltdUMYu5W/1jIT1jZSOaAtM6sp+y2ZhAU
mGXsBfQR6p9Gg0MRZMutmQxOgkVROP18aM+F3sbmtPEM/1IrS05RDrFxV2xzSBQp
sfRjpuAZUfwst2WZHFshou3SWvyosQDcZr+OqH8M+Xr6IVKdVHh1xZ1A1pYYEz73
BPL2e2XjIFpDODzMksZjIR4+cxSvLOkxBH5jF3uPpsNxZrGuDcZYcjjreZrHdmzt
gn2jNZlBCF52a6M5fUAPqNBpQrrcbkBE124XJfASxU5Cs7TEacDyGndGNizYraY7
wpwpKynrAIKRfj6bxnsp9DgGWtO47dl2htuLxsH/4zmbLQw2PXl62iRu2TmhthRR
nOQBCUG2ThiMM6RZIBRwi5n1ltqS+FWSWWaOSYheTtF84cMms+zwpyMfWiwffOY2
q1XRtfyGio9M8Nd2U/Z10J9i84nO4BtjZVLk0BTz2D4zp7fuzwZMCZiGOoPNP0T3
25V37oqxqbeBcezbvhlT1FNtHzHVei3pmIs/l8+Ajc6BkNlaL8dAKN7dA9hzQntk
Q97cpOTy9YhcnRXl3l+vLx3gzK9ULKqE7b2XLmH8c62aFL98Wj76Nh4GdfcJaqlC
M6gkbQYvX+r+RSrW0CGb8bjSSWSmPTQCVk4s1MXdVZzYs09cUPP1zKjBKOYKFgNS
uxMV8RS8QGw6kNDUCxUOqa/AFzIBWIrmztVpo+1/MKSGzjIsJOMk/F5vrYscMdwv
ytSs8ixyrjTVcB3ZMh7KR3dF5GaFnRM2kq3PCx1Vr+enrPAJa1R3u1IYGYRWL5IY
X1UzcTQsAceY4uCIVxeW6jtSQJJwEaBoezf/nyrLLKxZOgJ9NWNVtYzZuBNBo1z9
RwygrzuZ9hd9Bt80v73+ho9UpWd99zTPWKCW+HVG+C3INDvOk4J7kAcVQtVdkH3/
88I/1FxBWS7m4xwQQbrbb0F17dSsGD5tshtG2eA8QfSAoX7A99vka+BJBURwFl4/
fDw+Qi2iKF6Qt7Tsz60XVyffjIvRjTwcsvAKuUcoHtZzL62mFqFW+IuNt9sY5kNG
sR+zrfxokKmO3dVIqkn8MSs6+f760X7aX3UZr8mxtssao4F3TvSy0LDqOtQ4TGaG
FNCwmTz07fikozH7TO6H2f+QqZxhuPWWZGj5WjcaefiAaCqwzcoenyPSCPBMzS/b
F8ghQbuIbulgtEglvqUjmeXyuUHP9yIAmWZ2NXF3wlzkVpzSAR2J9+gzx4peHjU/
ub/z4cTmRn0vSdQM+tZqIUQXrOtNQkEBpuJTuyxd4I5J6ZsjRIjdOCryME6jJNb/
p89EjJtjKso/llTsVj66J6zQKDQGHy6c83b5tVdCua9GsD9LgCopwCRVGzDXX8iL
X72z1VIQWjA7QYmxHeXL24tClDpYqDmXEoTZpYPIDxIORMRnIdwD0oKRtdkwxMG4
hm3VQ+fZRZZHeRY7FDFttMw1RRILOIVJMWBmvUhERRfvlNsq3VLS8Riz4EygKndn
8CnUGl+RTs9ZgyMFBRv9aYsbnuSos++RCJnZI0IIK0f6UtU9eiYuC2NkrvPa9rO/
vSmIYzNhF3ErAuBucBcV3uovvKxVaDIYTF9DhSdJys0OQDMo7lCqcH+FvcF/t/LI
6N/JE4OXdKw46lf9Wf3thye7GQpGM1xYNyWP+izKeSx1MYC7yflV2vIcFqDdYFSP
zv1ybapUssUHlEEOi4QlQUD8LqLo7JYHDUWkyjvlqW/4yK8QZwu79Ngs2CAnZrXa
+tueatEF5Yd9m0fz4svQyvHUce+7V1jjusZwy/EUWew/BEvumyaZr/Zj012wQtKD
0NahCf6h30AhhSnJNWS2sFGOlovXf3NxpygKQkyD0Y3F6ZrsDbpL3qhZDj9mWbj2
w6o8v+ll/Z0iAJk6231qbqI407aZI7q9PIsM1/KF1ZdAwXYskWW5rLYWB6DqCsw0
M2lHs4yHuhb1BKc2nLzodVNnHZGjGnb7sb2PW0OxpsPQKuk8lDV38QLHOgHc2WKT
JAb9AJ6hKcY7NARif2EjkDvwx4t0397WBDQqf2/Iq7BObr8ffxuHqcDJcAxyJcAU
jz3pLL27pHRHBODHUCsvwhWFy3Ynt28zmYKfKs9mipuh82tmTOA2RrozsrLZhG8K
U0UX2pxgox9KNjD8n8Rj8MNs15zuUKw+PdGlbFuSbAdeDIX3L6+GoUKF9Za6EMv+
DvzkT4E8cL5meHMN86Us6uMFzG1E9Lq0RMrbtrfB+j99lsSSgoOr5avXu0yZpgpJ
m1nSZjS53E1rppu95N8tSxx6gVMV5noHz+eQPRyCFiZUwNwwMSdnGgNq8DJjJFkX
nKKFu0MDFvcAwQv4Rng3rhsWananbEJBLU51TCnnKpl8tzPySr1clNXMGrgZvNza
i6FfEDc6kYp0VTTCZaqgJoy04smXXiWjDqANFsX+mjJE7VgSg8ssYcF3nnbwxb/e
gvRU7BGQbgPm9H+R2QI4Cl7aQFurocm617OA3G88DTo7iQ+LNjWEAI6snlOgX8J9
2YcUgJxNATuLfn2fJ9zF3WvMprTDyYpvCvsSYrpx8gmfDIy72smCrTyJjROdeWgs
aFKHJdmiMSHejxYju2gYNqAOWdxT4Wd6hSkX+sAiPREHcxOuIxm7jDM+leUPilvm
fOHXL8hJhYWAthZO0dvon2pSog6GIME3182GlpSznaRapPEmDai1Res7ThkbXXMy
DXOhB2IRntRJ293bWUr9ieiZcA/JoQfzi6z+Fnfyip51JvTjQjes5tQxWZvbUuew
EJ4ZTlrk8cq5JuArkvDbqIGxxyDf8dm6dmKPofXDqlnsOUUMm8FEnt5xD7XiKY2t
9kE1Rb31J2IYrfxiz04cbKu4++UNLe89E2D+T6QqF79+0Jp5daFPEXufwx3Kdwyq
be/ZAoFPjaxwaUsfflPuof3dVG7EJpNEgA/6XvMxNoFcRwLX8ygHrziM7SvknZNi
k621f8VBsULtKGOUrlI0ooJHkYa155yZWyRysKmHl/lkmTJIktOaTBrmCK87jjo5
nk+GdkYPEp9kIP+Lk5zbnaga/IEsZ+2n+M7pJsOLLUuDEjkuUGGilzCobVRWK8qP
LHRy0EHdVWpzRVtW7od+Wasx8OPvwevzlrGhp5fqTxkw1QDAwI7zxcEn2GsaR2XA
UqYcjs9Q+CHDzg19nb7lNMY7wCUZEeCHyFOlZ+eO/1CGerOGMnVk4XeMS/wKnodh
9KGNIqLRsTLQvEKAIaYlmnnij8aCqdIA1jjOwuFlz8j+7lmtoosye8tgJpnBY6/0
Xc36H1YH22K8MtwewRGoWMkgF49HKM7EpRg3RbBGMu0KOY6X0547+aRqPfufzjbR
6EE43tFovdxkoRnN042a1m/yW541InPaGgNnwP7o8lWgaCsJIavuDF57Lx2mug67
Mjt7FyLs5DyI8FYz6pbZ08DSA2hcOzkjCpt66qDOenh3NsvKljY5AIFRm7moHydB
RiCvecsaSHyzRp/O3/7SpD+BRED+pN5+3fdH9AQhujKUcXq+ocVJ51D3/M97D9zj
wiWIBDdITpj7M/EsGDZu8z7jSWmLGc6NAE9RNRV5jtB8sWB9jMySAKsayKJI5EPA
mn+n318aJUrbQAGgcwd9YW/WBVENaMbSEYxiNmw1TrqL2KQT837a2wCLIygnEebp
86yjeL8r5wTlbx8NiIa++fOBVH6GmGmApJsjzWRWCGWseXgiw/PxBrtpW/xwLJN+
+/mrxor1duN8xa0Cj/ZdUiUle4SwQHKc5m5CAgXDQAcOssxGYQf581qOSPbyHwc9
RGTGesa7dT0QkckN4sL7R1RAkv5WuQpM3mvnkY9zBOnI2GYI9gKae36gtjV8shxG
GW0zMGeEMhOOO5ZrEr9EqEKNZ7yO993sS+oHeOp1bT19C1ufTMNehMXQk9ePQcvX
ZOi2N/2zuvf7ajnGWIunXLMZnSCdL/hriBllonmohvzL8S4Z9HllV7Fv3i9jkVO8
VGqwG4+U2nG1Kx1vZt34hSGL4aT6tdsLf0LKdRyoYrVnqRNfD+pGH8Dzp+BqB/An
V9StMM5aV4GOQi+ht53lhWy45zB6rgofQq5l94hEpkv8ER3MLnEmjzVpjKQRPxqi
sFRy7fvo+oVPOVBPJo1Taga1qGf3WVdpufhvZYaHR1MoL5MUSS4RI8U0u5noMrSQ
xMRu/FX3d64vFvMBS94S5H0bUrwEJ9UK//xtSENEQ4prvluvbziMmlXF4X8zXn3L
we9X11aFvZCsKyTbrXlBji2/Uozv/wM0C71sElyQYGyUi7pZZ7u8xyBkhVlNEX0j
BSV2JIzZwHkqaG6V8GF/PmD2pL6kd9/aNa85jj0zJis+RxYSATos+oZdjq5A69yZ
fqqmCNgBH6sLp507PW5+efM+iA5IpcosExeFrrhpF8ziClem+h3vU0eayb/gf0YB
RiTdBN2ZyaBE8D7jMkUsq90w5/bHb3pe8bftcKqhYm4TJSrDgMV+cziZ65IdBEkl
C2FGMfDcxvPaxStiHJL52KPN5ddTkiptzwK64Q9iBBJJsRJaVSYbFayKRGZJkD54
TXGu0kHyAuYW65i1yX/UJkDhDxbuu9rTS9iVskJLqxfp3+blVkz3k8pvsvEAU9LB
5gom/iCB+Z9nZgv+nb1kDcQCq9C2HDJe2DRC2pF60UkXynDMsUqOd+JpaDd7PtFn
pwqKtP0qYpBP3L8W/aKt6iSCox2WARdI5vYyDIL8XKT3c6QHe7XQ7+DhExh+Z8Rr
6nYas3s2kodEQ0D4XY8Os5aIg5y3yRJuzhwGcw/oDZa5qCpxyxeS1wXfMEnTTIZ/
KrygVID2kJDebv02Ac5SoGP3TkFNJny+6wKQDXbMI8IaNXF86FB4d8bqJCxFbKib
1znW9QG/99REEkkbFnWVXnguVWvJg5MXMTXsjVS7VtazbZ1Bq3rNImU7ZJ0duete
O1xlnuv2ZTsqmY1+Dmr9oEYcJ6jj2ZY29ELKPv9bKhSo+rN2ykH5sT5L7jtkcD7f
uEPUqCMFIxoC1MqDMU60Hf0yDpgHBHMQV+wHFWvxzCOebddVuffLuamABlm4kEJX
Q/TxFzyWqEuAaxGLURNeJGatRUNWumABYhVdh2pfRsuhf8z+DxkalBDr5OT8rfZ9
vtKryAKLo0L4P27szfYDJjMEVv1cNJhMDMg5Aj6X7t5PBWjwAN0HSNXKaUO+B8Pk
la2srIMRk/hxBGtQlS8rnB6cjfHV5YcGSkLQMBl9uwnbQGElsQmZdm9vI3e0AhQN
rX/+YtrpahQ2CpqVgY8JHveaJqwaqiIYFcZeGUoyhLO3yKGE9mjsD4e5pPJtOK8d
puuJwnA76k+6+1Z0Za5vp7NHzIVtbikTjBYLg910LOE8BsYIsUWopUGn3EWiY/oM
0S12n1sdCmMddIz9ogVEK4G/c3hWw4SbS+run3u4Rit6dUj6hOnIWM2NSS2Z+XKw
3YId5U1fk7z5GGVYbIFgAGGw9HXYLcbdr1FVMMvipq2reNa7YMdDWskSOLqZH/C4
n51oEgylFyhhjDak9aNOS67VF+i2qQmSICEd3HYR3y6a2YbZKjgayaHqh1yJy7mH
flJfUeNSrsVEYiAHRg37RvqaRhHGYLfuKRhX7H2JLC/jf0NOB2PtVgDRWYbh825K
rNIHxG2Yh/Bj0vmR2pCymQ+a7cRmHoFfxFh6QL7sOcKlzQc266r2Xo42Df8YV9WG
0nFktoXMMUqk12DsZdH7a3muwsR5vTsbyI2qkWLkjPC0fF+68iA1mtjY7/6SxQ3H
QdFKMjiEMe8aC1trKZs4gMrpw8OrT6PrBvK8Ux6cEqcoFzUVM8li92ZiPsw/UMXu
8rd7wUAjKfNEikFIXFlYvrDNJVfWpV7jCOep9HxtdehM3/RhKWd3sMQoFphVANC7
M6gD0zKEp4RkvlzNYoiztRw7v5rQdzKGc6QdTXV4CRRIxrm+sEkV217/1FNNzZ9a
liW10IGba8FvlPe5USQOGo+Rzx06Za+ww/XpyJM31Hqjw5JbV5Gjj5cmZV0u+6ke
P6zatRHHeLnqeLHp7J7XNQyXwPiI0vX8F7aQgi7xZhABv5LlwQrplXaLS6Jtrmvk
bTX9rR2mFrKZmC6lwZMB6gY/HFEs7ixCVveAhMnN7b/mTHYPGP+WzUfAG4V1eJFD
/yNvAeW6kMu8bpUQ2ljecHZjfE1UnKlYueCwXbSW3W8j1q/yiqbyd6fR/VtpM0Ke
t/+ovtq19eUw4NKWoKBExdoS9J9QY9ZQPrkx82xKDtZTyC3H4TCGtHwDHpihdVTS
vFSGTr2b0z1KctJPSJBZ34qm4K14n6+BJ1aPhvrpcwBunsKJo00ETDkzhLLtSiqu
eJF3laOentdUPVUyli+x+fAj+2bv0ZnJT7OeH+43Sk5s4bd5uH2hScRXH++q0S5U
HzIkkCr2pCmaQQ883iOtjktAE7bHX5/6P7oUF/fv4NgvzQtb6RrgKShOzIM5PSaA
Qcfaf/pE/s6kn0JrC0K2likkLNSLLCUdZV/eptucSBDpCd6ElBgDOTOEC2sKYvdN
4K2qQJqWFt6czL8FyzOi24xR/yRUy4n+YH3pwz9PzRTP9A2jSBZCv6FQ2Xbi3s5x
jx7f3t5lGkyu7icI7ofis1w4Ju7BMNxm60deGFWudXcPu/hdqm9ApKXK6fKRqVjM
Wm3V13SL5nR7R37iPyvonxVKsl7FjwuSyQ8YTiacUWuyj0UnAxeG0rdZO21IOuw8
jGpCz3JLlVOxq8Ay7Ils3yalb0GC0/JqTIz24vzFUJYeVWi9OAErztQYF1Jg1lM9
DdQbhNiu0OOUh5QOMLc5D90jCEHfdqgE+GVUdGq6v59Dm5wQLbwXL9NT8uRHnzVv
huVaxwnlQ+sPqL9p+UgR6MfUkG+8jdQrtSd7HcZCQCNVnwpzY8CYa/PfRjLh2dD7
zwqAC9OV4COS/Eb3dZdlbobHSEUU29+8ipVtCq1s66JQmK+h6n8O4YkDOLAqSXhg
lMzhdseQX/TsA8VxhhGysbtwY+4tKFF1xO5s0+gyHyX6p2mhbjZSYT9EPh1ssHmt
L94y4HYM2zsMcvGOvEfZHLCMZTsE+qtVoehSSxP5OfOBpulzwjdwi7cAZu3js6tp
7f+OTM0UQTJuQjqsI1UXx10XCx9uSMKowv5OZrXbKH3g3rL4ou/a0W5YOVJe4JV1
V13zLP3vB22WxRUik4PoaZ3PNk9v2GOF0qKIhvgpQEJvS5pR6jB38I/TPg2jmPGM
48l93s5hsN2vq4Wfno5vP1hCpzkirW7K6qoVAOLIpK3H9CsX9A5gkJtH9p30jBK2
g5LAvqsNu5CKaODBfpq5JoIlo7e2xdSHMaNeKpESKtNXBBja0DpVAXOGLt1e8x4Q
sE1Xu6e0H6UZF7TrQ4R7TtGBtdH8WktooXCXOiU9wDqXYDL6DphSk2K2PxcSFY2+
ZGNLUjXhCVRDPmI3DZnDG0z0Q32bG//lUw8C43ieMcIEoqYVg+We6b1elHbnVg3I
cjYL/WH3fWzdTzP12j9oCZqRrNP/ht9cQU+GO0a705aQfSUBkE2fqDSMYCYVfyD2
UN8V4wRyCXzGx4h70C2Zn6pfux2fwE4XBSey3xkeUhSjB+7L1+BlIGY5OYwOmJW9
iIb5YS4THMVLrFwYnEariThEjvQfVnc/caU0sKSNO35JFbJ9tXNcTx6ci6KHXKu2
9ihfjlwfJXbSY7WooId7zEZE9iMVvK3A4LLuS5eNi6xoxyFsd6TQ7SXVMeGMjo10
EP6M+v7h3GFHX94Q4XK2mb/xh5LbRWoKoTIL0RVOGEPAE37r9GgvEdtnPgohk9Zn
wgGzpupyMuXNVuc2jMlTcwOvZeZiGUYcpNq2gBg5e48lZM7qr/LNaKldmgQB/0cz
WXXfF6OOIJYEMbTNLje2lZJ02Qu2IP7Kex8gukurF2OkdH2qKrGGu6VkduPMGAvc
ZrWdoVfjWh2eRzgplxwAR4Ugx/CheVm6V6itugA4HlSosttvCbF/pM5nIf0htjFB
R2hBPprwYe4uz/hgSPYbmoS0lF1NLlGv5vOoCTHkYnPvWx0JKCclRTm58kNKlyn/
sEhNQmVBoiDeIXBgxdOoJ/HZoxFMgCOr63tjFrLAkJNjeSuvWof/Xs3ake9tidBE
rrpudEh6Os3kPsYJhIlWY+EHz9NOur49nnVOneP5Vm348hlJztqtcyFFu4MKRS/l
xNzxFFGpZKMtQUAB88dfMeNAut8HGXDVi9bS3facvbh5hOjJqrLWUxDQWhBLOZLL
yY/tAncFputHTKdRozTzkxkq9wX0WWawWIKUuuy5jzC297ntsje/39+oqYC//rw0
DER37SIitErJQbyNGj0438MEy/5JQWRBS4OwuZTep6pweAadMCUfys3Pej+VXLaI
vYY+LSHcPbK4t/dij4zfVHAxFE+jyPyHWVbLJ7+GuTu84GyH7V2DZLcIjuX7k0OI
KfI4zfTkK1sVvOHqczV8BRbKXvZQvv2BzltgCSH1vV4lrbey4OnOaAazmvbIGRDJ
X5hhpbkNmKUsQYN8TvOJi7IbpAWBiW7UEhsQ87xq4T/wD6tHeup42uk29Y2NbsuB
KbJKP+GhnkI1Qm5YVGIRLiQUJHtDs/B5tDOwt1DZB+ZS66OamlPgO4oIwTq+nsOc
QvsvMCLCyj6AvqSBB3y3qA2SPj7zjfOD+X6zQU/P01HRkEQrb6zldHp+sLaPAGol
q69/QZTti4atf2bChzGi6TO+vtbiTJn60uomAeIcXU4oQzX1EwVAK64spE3IKlsf
+SOmv5M/Ve4dggIED525BkmCUfzjmqj1D9wm+jDZgkw/gfRxuxYHZS1k5WSTXe2y
onNgcUoLQVYfhKTilhPTo3D24+ZiSEf7uFiRDBZxqHPnu/9EstoHnxv7yHGSSAB2
p3yEC8EQdmKPJnQ5rtVvOvtv8yOh8yOah8M0FTYs9JtdJDgO51WMz5xcNOBu5uzY
bMSTp7fPYUWUIiqsc9ouRG3rA4l0rO5yW88vNRfxkDClJNhWf+RtFp7fXpKH1hlz
G8TPWpU2pLxDPUrZYn6N3nSu9N616mAYKf1oqWz1k9jClDO0lPVnnPb/apW+BXqB
uTrfTN/inGkbJOnIa1OovMm6hZzuxQo1ekg4snr8iq5XT9ClUQEkIzuy6YnjB0aR
PEe4AYHpbiU+sA/zJ6UqOmI0rgPJrfEAJsWioTw4HMRJET8kwPn5XYOdoCZuoWgC
6PCgwvE/M1qbjxLvCLrJBD5GmbI95OV9GtTIyRzRpiURPfE4D1pUa36sA5R9OOmG
Mh13dWQf5U+QGRXNLOVgLojGWEC7CBCyHlG8YtxyR7Ee9V6gwjC452vXsL4pPk0n
rCZivhYJBEaj/aqeOAkBuK8gYNj0pdpdrl6KHuXUyW2J6rNT3OdP1ukDIisZWJfW
RVPTyKFnWgYwGzujvzimB8IF0nSh6arPl0LHTmchU8k/lvQgDSnXjKM6Zk9qN8bC
0k9MgHize3ISjZ2HYDRt+Fayz+JGIkIo4oDLvBpwrHD2RoMUTDLgXvFrs+AaOOxC
WqwPEQAGS/vmpF/0oMMR02GE5eQLgBVQuk04ZYzxPmuGQetnRMTvfxMGNxSgrlfF
QxCgMCLscPokWLSTQv6CdKBpB8b74m9r6bH+g1sIdJQe7yrXDz5OaakuySpFM5xY
XE1vzdauF5Zk4aFO0DlBuV/Yy5vKaroyo1eI0atAAHJYb925Rq3FRoiMSrPUY5eB
uyp3apXvcFZA26AISyXnWo2CWW4QBEvaKGW1GW3pvfWRrAnAl2YL8IZIuw6tKdd6
HPkH4I8vf1aa2B6rkqovTn6zgILh47wsxgJXaUmkATpxxsxibpXOprfz76uHhpJc
zJHb1Nj1LfHQwgDrLljGi3eRxJ79dEdYeeEJkB2ArZw/oZ2FMPkh2Aiox0Fhur8T
DSlolO35fcZW0FYcwmVu4YBQ8BgTS+eCLvZFa1XwrXukoGFByKR1ZFWBOemwus1n
IAXj3xtXgJvHqqxa93K1kIwEYFTLzYxJ2U4cVC77HYi7n2UDuYibnv8/McKwm3xa
dGacoTm39zNwDaypesA/LEAdFfNaeYU1UrEYVIaaLjdOerEvs25ImJwEk3qzb8Mq
OTNwrqX0JOVvYyUEpRDwB/rGHwPsziANXTdD6eObwMd0C2LcywPyX+R7Vgf/z2Ll
Y3lI9/B2/x0OmiH4g3RBRmgnqti5xErt3fQSqgBYtNV+xRMzoqE4xJVPGWz6LHPZ
/uwfoPHiA0CBl6jROkQ+F1pWGU5b2ELRcqhPbE6CQlzF2jEy1PIhICj/WTji6EUS
03xN+yzEcB0wem0YxCYMJqOxdsyfKWrFG1tOr59bvppzgOzl/RfKb4x5DU8BXOWV
m0rocVh1qN5ES5br1dwi6b0qEJZdHC8ixHs+L0EsKawiOjY9+gmKuDlaQlU/1Mqf
p6RAwvVZF3bNh6Wshm0/eh6rYDTEGqZWiZHSC3kuSIzsGljqLK88kV4yzGxyAecE
/qb+9dgH2RMkwN48jMOjxX6mA722NkvI7Dsr4a4bRaOO7eq7fM881fah/p1mW2zl
477f9ZxYZH0eiTHKf/POcj0TnlcQuoLsvIDSjvyEamikciuwi0Yn1axTG7k6cAfi
zZvyrkhyLzBPxOH6laxMLs0Omsa1Aub3gMOuI6vRe4u3Qayn48PyolesYaW0UUSJ
vEPNwT8TAyi0i77qS5H0E8XfgawNrTlwE9Nj3QYTj1BbJUNO/CYrHxXWCf73tBcY
pA9ye3giu+QIJb0/Q95mdabsq/9iOSlloQBG28PuH9K1H8/vRCHMZjJET9ojK+xB
LKBOLBYKNuTnyjwzPjYcLZtatNIZLGsxpvW0tu0a/JOSb5kDXdIknnwr7+vOoNXZ
Txa4tB8iNjeZplwh6eVECZi/k5LupF83Ma+SDsePyRSU5I4TKbO3Q2I1K6cJhFJj
sDN6kWA09yKR0BGiMnTZs7VsVCslDaD3bVq1h4NbFkz3PfBWxlODG9C0EsZU6Q2i
aKTGsoTutjGwAS0l8aQXO/wD4lent3l15XYzScjlPr/3xJ3inLUOruYx8t+6MJ1k
R3Cn5+zbPCLUqluVLaA8mi0lUWOjEQsPAqwsxjIcfrxgp36eHHgkEpj4qd3BhWod
OWU4v6d3zuoYG2XJv+2va/MzSF2e84jwysjFwf/VzbaYGIkOfHtmQTgFeEUW8STD
nPAZQ53NkcvmETpGR9S6TmDL54Uo9avGgZpt5caYj6yp2sJGFa1XXiKcP62yVnpj
`protect end_protected