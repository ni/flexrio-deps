`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 38064 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/clt2ISG0lyjZMFR0pnYo0pZDC9GSCYCxcgBJz06EzD0
3gJfsz3BXYXkqvFvd0lCXGes8rcu8Oy+SheaO+HhM/BzOMS/1uiewLXrfq6SNuFY
CPU76663c+NgxoIcvEQlKLHFXIMnNdFL+p0xvOpTVrUrXXWAMtmd5LVANpvEs353
KG9bC9gkpAOGhS5SgYOULgyGMRbni8GKFocCCLuNm0YwLiIvUP2595I/eo1j5sH8
EPFOBoGX9ktdjlzhqpTr9VvnAl2Xt/A5PyiHhPQghphg3dj71xx4zggkR08Zzcen
70Le1zxXuxBPub66DJtRi7vhs9dECfKP3VYhQ33LyLY1NVPD+F5xFIGfFMu388DY
DRpSuQrtwIAm71VDBHu58hpUeWWKBFAd/1m63ZLW9FvrpcZmCSCu6Lj+Q6mR/6wz
0o/CMHGkHRNo6AiNKFbZKj6R+AJTOzlEQjc9PHoejDZWASdt2rkgdA+JfjtFHCDC
ikokaRAA4lIVFaH4OpaNAoIWcr1eCp09ZzpyBRCgCBGgjboF4U+j6nVEr+7doO8/
oks7ObbrM8GsvSm85FgLjIXoCPp3U3oBodLD47iQ2jAtD0LB6yBAzcaXJKjfTxvc
+eia7Z8VzXYPrglNYKA8ym+jJ1uk0C3eXVF5Eqc2oDUpVDY715KmiyNEgBW5lwRu
6lZn9b4le57mdFkSyNJXzkdCFdHTeyNL3m1wmoZbF9Pcf3rgSzAcHghXB3+DCgzR
6kxcd9InijIGbOr4JeVvRzHJfcYuAulCWazD7VqSGbgtBXSX3nFjZ/Zr1QGktbE1
P3SN3OYDuIXo+iVV1j9pQNqFdIA1pZvsz6LYcVTwfLTEluM8GBnn8jLtbPNibunI
Bg0ysjYWddycplIQByy3F9QKPE66xSx3yUVpU4idAdQkMP1tLU/vssZvjOXVNnAp
UBYfYz4HUVmH+CiXoW6OHbhfD3XJxweVPdtJSt9whMPDlaxaMDdC2cmLf72zAluM
Alp4yqGB0F3KTe9Z4a3NxeR+rpuYyc/QT/shXMV7Fj2S0JAR4x3RuQKrkobvz59f
auFwRBRdhY+2IregHIdicOeInEpfX4VMOFmAIkidD240uObVV89+F2WczFmGiYh5
+QQQUsA0BWHeCB6SJ/zegs0gdvvweUzchHEIJ6zE9vR1UgMMtbzdIA0DikPXyLxx
W5O6allNoG17PGZ7gm+Z6yGCh1yWO9ZGzjn/KzrHpD1PtPgS/E10Ofllu6BLgm3r
kmziBOI+8CINWQcJHhIRusdfxYaEhF4wgTcS/wMqLzQ/gEQft6DfJGjHa0Y7J6ON
hjcQkF+d9Z4yBIThKVG5QUH7fEdIuJYFJE6yM77QVkpowpMGWF+jL2BqxGooa42B
b1impa4pxM3GRi97ketFDeUZuaL/4NaUosc6qjJUWzLu5UwZGj2SXIUbTxVtsFUV
kkPHHYampOc5T9jak3y3aKPf5osgGwGKOB675xtNtpyMj4+SXlN6fAONKtqqAyne
y7tSpAHFRplHB3tWCBIX6bhI+lnsfyym4/l12CK8DrHhiXClmkWKrqrFN4UjcOy4
hAeF8VFhVreCMGQSjg+A7iVNlzWM74uFeEBIu/1dDStuxM8XmmyPur9WBfr46KpX
HiZq7my95vwT3hSBWwuIXa3CkFGBDrJMJ2Ge38nehUjd2bPd4atM2RMSx4+Lwu/3
eqpEoOJWdSZu5rWzUjrtzuGFKD8nCzL/EMGDtnOT4ZE6Vaj2y1cszmBI3H2zTUkS
rnAEJAXbKHyPOs93huFK4msaYUe6ZYotB3/6dSNRJJI9K9BIm1VvEGaG5LVV50Wh
KRCibgbjxd+QShJ/IjX+io4ipUmCSq9w3L6VKf35T82QPmUVMI2iu0SdPsDSYtzF
EkxbT1lUe1WBVmnWrdwdfGClm+nidJF4qd1mzLS7WOjj7Jt+s15izwRnSUhZAy2K
OhM8fM+OgZqyiXEVKCHQa2NmdBTuTocn61uiYb0TicpWFWhE+DTtIZt7ro3kjigM
8nCP5ualKc5gEQ7C69NtRFdSCvaPoE5KnPc3sx/m6of2C0LlQ/CUFoPH3E0IpOpI
u3kTFI3m8ILMn6GbXfXlDSm9d3iG/hAlvvMI1ec8+fF/FpBiJ2ISJyIx9b2JPDNh
t84PrziypVSY+7sXh+wWuszx02YkTbLCcL/3G8o3z6jnx0r2amLB1Ywo0agWhUAK
bUTZysB0ULewfr2n+X3hytEVEznjn2s3wo1hLNDGyLwjXU3F4I6odIFEqgVQustc
BbCho+so34fmKlBB0rzR0o58P+hjKRAaPAt5htIFWbj5qwIedOIhjRlbe8n0NezW
QYwPhlSXC9jPKuL22TeVgk1jGNebQwianVSYnNORKcVHYFrvc5qG2lrydCt6t/bg
QPHgoNdLx0vF2tH5AkNqcoarUNZ+KyUNltadEoVVRZ0hBNlgwhCUpy/rPBvUFz6Q
FP/OnOomnYjwKbNVcWlOGvbEk/8So0k//MCzCIcl/0W5hGxruTx1IyvsT8odCqHH
YsnavS5CYIw+zPERCGUj19e/K9Xg/6Q9zCYheSd5hSoevgKtEKcyyykqJgVW0fVB
fE7zDXwpK1eXEQI83ol5nmXyvfqD3oBT/YQJgdWPB5kYNb1Zq5KQ/NRIM2zV0IBT
/TKGD/uv/IXVRSRsUvN+1W3lMvHs8azrfUDLMr4VmP4F9fZceHonK+IJmqy8Jz0K
as5947CRxeCKwgJg08bIvAo6VxzyS1YIw+vr0fW2Kgwe+B9IZnUjKSq/+KJn4Hsd
xqZipmXuSTWd+HTn+Jk7qzBgSW99Vno0PDoh6IdKh6BTEY9/+3w4CslEg+aKStHW
I8MYG8H0mPGynAz3Khv9U99hlRSCtZ+VyXqcw2EunRIgbHkMXwz2GYGSXslW1M9c
lP+1kPyAYHW8Y3pC8mrbV50In8YtHSqTE1zH3afC+kqloYcrMc7Ug919hIPhiaGW
64gQaQTR0B+1Ph+6mdUP8dm7u234IkmNwxJr2BH02zN5Pk/BUi9ysXxQDlxL+2K6
gbVwnVRAbHjebAGaLwy1NTp9KNdDF+jDMVKl+l45LqpnIQABG3EWyzv7RLsQ0rEW
EbJ4TtWOUQtuOmSBfs8WH6y371LJpHO8lYz8dwomax2DVzxo2xrfP4xSbuWDvKf/
aBEF1iCr+NfeV8KNtoJhTjSNPbLbNc+K1j6JFYZclPYkVpsmBWc+JTBUxr8DfbVY
npbGymoR5RIt4FMR6R4YpRDMS9mi+QumXAB9WiH5L+9sLKR723m5EJG9OAYk6NAk
NVXLgXunfphkvbXd9ZMUfuD8R0M26xudObCzRCTiiM4/KdzuMcAK+hVeliQuwCzu
M1cjfexpYpesVcoZPQAG0gTS735erhXLsK/2JeBRNTjeBNVT87YjeIlOf79A56bm
k0aQF1QSUWsYXk/wk6+mng4B69P2yV0zv100ZCRM2iF5CSOsY5vAfU4oOzVCSoKj
XlZXWHeExGgafEXI7LPU4vCsKyNPlqC6L92SebOCPVfA1wR0/8DRhmTfMSGNWlQZ
NwN5/T4mn1kZvaB0rD65VjNK2AUM8l65w6WCZl55C05FV7xUPaixMNOapyGCifeo
sZd1wg5kgg+jFYWVanYSiARHJqMNwjdRi78yA7hv9ASRTDLUd4WlUxEE+hG9lmEy
qhA1iDcb9615LGcGAKbekIqj3YqLdaQyDqzWvSkquzQp40qvtfGKBrTweicRMSNz
aPGVL9Qy1XBE5Di7vRXd8V8shCEl1TTW4S8xJQFGP2CCCJ590SuVE2BcMUTPFLLW
f4nOeLAKN0afntGZXhRZ0RceKXtZ/LRUiiX7Z8B85aHTYsihlZjBC/3Q953Bj5Sx
0+haGxgGfhn7IFtsjJABDcBvqw4b1SHxUDKv2VY3B9JNFfIttwbC4SwDVcrbaHMe
iZRhavSpuzgyXWXf/hGfyg8RF3/jYsybmEnsWoZT5WnRGtYU/3wz5MpHVTF/TFIP
Ou2+fnmL6YSQTuz7WB33Ts5dW+PcFORnDHxA5o8KzbJhYL8EdDa2RDnRpn2+A+HS
Xh2KvAAbW+GKMwNaauW8kTOyD4/GSTnkCBcNggGR/LmY3SmJt7ukKPySafGtzrSe
ta/kGCFZcZKMpZRxUTSx5+6eUesPBwSPL34Z0F7CgXhlIB32Bmyd8bAjdg/f/hua
R7C/VhJuivGAoFKBxtjj1H/EpE2bSe4vsqCA/ZjzkzidQOzglek7hnhSFkRi61Bz
WnxXjUOMwF1MgErCHD9UDwu11jxvXUZZWgbQNKn8EzZccW+/KruAo13oZHFMLPc+
CETVnz4pb5Z9kdi97KCKl8zYvGr85gMudRZU3HTMdiWXNz/gM4SHqGcvNiomRUpp
zIRbaY1D7IHzBfJKn0DQC08NrsTEs88Bi1wJLazDGrlPV4h01hM/fXOPWa3mmdNH
Rzd7lTJ+vbNol11qeQkxbMrS5i2MbJF3tcAwXxrKvQ7c//N0O4rA//qkPnyCkARq
b66UxjH1FY5L7BHK/NQIguG2aMWHSI0MZy8wkNcPUbjB7+M4BCFjbbkPi4cWe0to
6slm84SNUgYhJqkiHGW2rUa1k1/vgoXWU+p6iYv/QoRMyIGxgtiDmu4+BouH4oGv
EnuLHA7dHwoleWu4bEPuqOFp5RWRNMu9b44VymK5gpHTesxEDdxJF6BM5NjsmTUz
RWZhyW46HfOzFG0FPkeAHrBJXS9GjIcSopaS7yO/EbPst8bSiJZJCU5Nbh3IZoDo
KAHdga4oAPV3en+Iugf7gNA1+uaIz2N/oYh2r0gm2+RYE0uZLhk8MrBQ9YPcj3o7
hQIzUyfqtX+vZiOC9SoVXk3D7BVqpgev6N7cVUoomCYswLkZ5JJkHx8ya7gsCU0W
TRuH2rkS436B4oqQZj5nHbCL/i44Qrxj4Y5OtIowa8RxLIj3+08m9eu6Zuglf3DD
7XsBNOMt7awLCGCwIa/wd0tZjN9a0upwfAKMan8PmcFhsr8ns/ZLlPylLSARrLN1
LG7umR6ytjhJ5/L4FeanWfbaws+a2bC7MD30MbUxjicMSCFJXt6/cV8ljweFVgDy
wjz54IkxYCOOmcsJRgYI7zo62szH1M+GLj5vuc27rmI1L2/nHr1oK04yHzbBlesF
pKTS1dW57+GroIxhDZ6W5mQHXqzgD8CuJsIxcajK6z5fVMZ/zEScj/t3gnwZpUbd
qjD3QBD8dUU4jUY6d83nwUO8VWaez+Lpf1hperfHokwgBCVrNsRqli24LxEa/Odt
iKIAk1dBOP9TahrBUF/Vx4ua6Kzunvizc8s+/amyaneydSepIVV090Lhmf01TmjK
ZqsoO3PDUYLitrgOB0OAup5/y4pz1f0g47DdUN9z9fkLvYhJygSHVmLsBEWSWr6Z
vCMtyHpLNZJb2rLpyyi/Ne7oD0k3inR9t/cJVOTjCBYrirNomeF/1j+ziG8zwP7r
XZ4AF5Qy4/cHS30lJ3O1NWdAMOHZsqEe0/RuHdZtPtoWr3BJmkrd4msVcKB6QwRc
Y+LH5ZykKg3Jwe5CSsAs+Wd4W9SbqrwiYsduOo/kNGsKpUV2FCgEjlqoL01A+rBp
ujCj4K+5AT1NsNN4tfgqKkfx3axSQ9GRhh9cC/1SBjAVvu9j2pXQ5N2ocbQWvhVn
ANMxSq/rSRmAjYjbBoNJ1MvcyaaCRUMQE4gaon4u0AJqGZuJUuLkconWqRDQi0Di
46K/rmnF8AszpE/mGYiy5PrEMewurx3Vos1tc8BpiUmp40YrOr759q74MBCGkVxm
3q3QqXsh3NcfGZVZ3vDadmgfkl25GRWX7AiVUocnLuTNEukmCk/3OK72wzK3896q
1mAhgJ6Ubhu6F/Ka0OFCu1ZDJs1H4Rh+OwcVqecfwKdsD9x96PTQieiObMxgtBVB
qFrw8yemZ8KymgZQIjPY/4MmGiktZjoXLcsUYu0eGVnL3ZNrw0Cu43/uVGhXTMOo
htaFBGtbi8jEXGN159ftYCJT8AeiQ82ENVeosHdfl7HvOeFWm2vSXALjOqVJZPtn
6hD9bQEHEmIw7XhrQSqDTFehaqnsLdIM2TgSuIvDH/oACX3z+mflh3fkQZrv5w7t
KhJ4JlMpeHVfApe9vmrb45j6QkJktzJJ44VdAj+YQUwV6vLbOo9gUb961/QEfoQK
PiKPJv3QtjGFgry4+Dlv+9O2zVOlGMI5KEQsA8kPoS1ZFnbL+9OSEgZIrKh5YBZM
igY+oKtbc+cU5m8iKrrk2gNdLu0YyjHh3abnmZxoCvCF3aLGujBFCHyHhUlAuP9B
6DGaQsy9GS2HgSGFkgCZHcDnMshVKranNAytpuvdVab9zISlQfOyEwud1ym92Q2D
s1BDHtdvRnOp4ZzSdGhlEUrWMFY2Ia6eLHpuE8ChIfPfr37eP/ElHbT4O1+wi8Fs
Fyncy82V90ChckzX2XnBsDO9rsFoqHSArQOLTe6YB39D30CM9VLG+Do7RAvVftTX
B1zufQIruwdGr592O/KiZevpSFUoFcVQq9bIVATOpYUcF5H5QhDQcP5JyRyTaX4L
pKW02S+zlP8XuXCDeTedlMNaux+F3u/wQtnOVcb5dG5l+2pyYILhlcl62P1/LjuM
/5lx9/8rc0mmKYbZwjTTMTZpcGkBtXvMSCRlvZJl9FqUyCpvzDv1XKMu3wi1FI1f
IQ6XQDbxDDTOuj0SwW5SFn1vHnk2oyQQIivE+w/zVb1nNfdOBx8xGffBmkyHtKQ2
niTgcjSEV8kA+xzyNi3NL5HzFCar+VIRroXNGSnTBi9DgWymwtUmIxGRYNFxaXUD
r6F4G4ktlCCTWJJZMAr9pPd5sa501i9UlriHCkwoSh0LfiixYylvvcAMyDNk/Y/D
jLMpgiC5UeUX41xjlUiMfabrJoAv+kC9d61+T9aeYKolqWfTKNFMIbIZ90PaXXOn
uL81MkarALbOF5CiGWkEif6FOTl52OwS67ZkJY3OFLmJeHo1OEcwjUHwn8eYQZmP
odsEVlaznKkWGc5vlDLvuwV6JGABFY0P101h+mJkuWty+NOYJh9Hn4jZqWN+z2+9
9KUfhamG427RFk0+grEleWqvG+ES40ScsgkegRThPIh3QHMnQ37Mjji0voKsMu0Z
WE2dy0+q9nL3d8LQho7heMrzbQfV8915KTVUdObRrnL+yhVMczKbYQUkfu3VRSXy
nd9c2yccLdmW8x4EIq3nQVJqWMER4xZaJ4rXS92wOEnVpGLJe8YuT8Ua2Jl1uwRI
LptEqfK5SMOuAIyvRhINMFOs5QYLvGqllgO8SoZit5IVH0kQnodYO/AZWE7QpXzK
5+vPUAYeopQMmGc9EHj4Uy2Z0oIOutwpPh1P4TGhb9c5FhqOpDnlcUZAhGI0pV4h
RH/6z2StJrsksVRt2dcrNClFZuDPakteO0y2nR3m5N6smsxD2O9FCC5hsdCmnGw1
j0GKWDHsC25kyor7+zueaNInSFvOB3ukC2pUdix93xRdRnjPr5il0YZzxcZ6GR2J
D3pVBPGWO6IIsDpg8I0zG3HxN+7UZh7k07o5F5UrvqBIjR8CnS2xVznmp80WUpOd
Rk1QUQOqWsFfAix8eQnUT6bobwTWqgvOxOxQXzrYeFxkyeR1HLQ1a433+RT6ASGX
4my2JppT065UjqVzCfqQTc4aJje8zma2anRMCUSffPQna4sSYsMimAQrIxOJm/LP
4zg2OheEstvz6Sc5Y4ZVht+E2g8yi54O0NWbioHM8bwfIhSccXqv9QHGpOXN5Y3B
HP5pU2t/Z4ls4Fd5HN+IkBJTU1r9reg77XwVO0NQLiQP7FhNMOGYKg9zk3oTEHvI
+GnKhO9Sy6CnUDIKS+MCAi0kXTp9sevprbuFDCGOfBSDQggnLvVNyoftMR4VWY0T
sWfxI5Iwgzr4Qnwh0pVbMPmX8my8p5R87lnVRlAmX6/9tNxrTMZ250bHxLYyHtI6
DQsw0GWuMmMpXAniq+So0QRNA2tQun8bhUKdWOTC1BQF6AwOFb8pvRs8izFA3zd5
HW4X7AJ0W9+dBJ5wF69VeFeKZm0K21eIG6e7jX8oyde5X/RDDBT3m++qISwEXMG1
YMfGaNGFDC07lKFu+CLS6AfySGuxICfZTgAMK/Ew6pHidC4SlH10KaJmpAG8MyF2
OBvd0cOjSR3R/9Zm3OYNwDbyWME+qt4MU0NYfLjgeIJ9LhUqphS9XxW9HehtlxOI
a6t9MosHBvroW7lcF72jRJNbkKGa+tKUBXZVX80Y7dOtjV2F20JtG0P69AhnTyg7
MKfuvlKgklhRYiUZCsdtcrxpncPLuiBtr5gdYugdcwqN7udZncK0fs/EzkLhqF+4
FVqi628hqqnbs72YEbhT0Tq0yoZJb2sROqQHs25HSow45NfdyMuixMIg0sfS6ak/
N+9+uJ71t5tTM/EtBEaH1lZUkyK6NAmNiw70Ck0ArnTOdhZK6I5Up9Ei6yDZ5Atu
quQD4xdThP5Pu6THxnpSu0/VnMiDGhb6RhOihZnl9ErIRNHlXQNwl7BOnRps6i2X
ykay7lrhPIGANDWXR+Mm7kXjdMPci2dvnYQ/YgBqpXX2ZP1S1K3dwwNbTZMJUwNW
pqA7ljUCg/OdKxGAE9htsFjz2HWewlfhV+R7XwsQ0/LN+E+PMp8W9lXk5zXWRn5E
gxt9jW4+ciDSdHuBXtxYLThBE4+sYhkLmpfk0tMQNcnhDwnhd30tjrQE/bN5KjGl
sbLr0yWCATIHIDfCdaoAkku39mjCSkvqHcSSHrfu9tDyoQm7+gIj5O9SZa3Q8c0j
lE54o7kRcVvVfCb7YtPFu4qHDgvMF9FsnTo+/qt2nXTlA79KJ/fVFq0NxjeaG9hh
M0mf4+UhX87I1T4SsYltSZct7KLH0X1Sp6vE8nYu5bCNqgGB0wxBns/DKZOz59sd
Raq+6dutGZq8OWp+zwcfdFYrXK81101MTatlbsLnvjkFp0o/MGzbRjGQ4Q5KpS7s
2Xxu2UFl+bEmXjabR8Q0epBWvy8JmRoFVq3CXiu8oTFaQwVkmWQRNBmkkKru/MWG
B2nzbay8dQWQR4e0H7gIGt9U+ytgzi3nwGiAX0tVaSQkftGurxxGg4E73pDliC6n
Bh/QDms/jdrVjGos5F5ZZz7UWiMQOPh/b12mcUGXsMDaK0i1K9VUuEUlbswV4ASq
JhbdzCvNKxAKXne0zcHE3NX3AzGDsQZ5JO2isvRF129BrESWAAKl9bpsgtf0KZ1N
AAFQ/wYL8RMt2kZ803KVoHu9yohK5vUH4V5YshVTpzgvYduPVgpIse5cm1YATuKd
knCzOZWekoZkCOrwmPVny75FYwFkrC9GuEMqai+jUyfugOwkNLLyusMhsg7POegS
WrooacatnYYfMoH/qqiqsv17QwlxcTER8tN0QioHpNQd/AKP9Lh4EZp/+1+W3LOJ
wS9/Inyq3MhcVL5fSmZ88hWsYb/4KP1KnsRDAP/ycjhykNa4Slo5vynCAhV+ciPZ
z8nDkGWadJPx4Czcb09O3l5vM9JHpRkHecOCOz/P8cIPB8AFBT0SBxUsyfNoWcvZ
E/xcqXV0d/8l+qGiVFwyioQBonTub2VfmnQ0Cg5SY0rj+AR5Isgv5yFM8a5Q8rWN
fPsfaCpe1itFpqn3ef1OTbzQyJ9f3Ha+IxTZ8q5kWa6Fz+0v2zDSV1p1IUbCd/tD
Fptx3IAgzIMt6qJ3gPJUtZLyBQr/8vXoK2R6jWdbcEoIax+w3obrMg9oA0c94rUO
FC78/0mfWyVGk3uwHlDnvvWHfQDyrxaMiJs3tXyHsRAIt5DeG0jaidokDlqVRSXR
lsi5Bf0mJjF5WPRig5z7DSYAc3sT3ldQUXWpb+ruanhyiDD5PdIf0nW7qFoXZo02
ycBzXE0nI03BisNxM8QGsAyH5IpZHuSGP9ILjbznAHdGfI56Cbbsl/I2t0ELtWWT
O0Qqe7yChjH9IcOEXyLWAWZrblKwNVv85vCbhy7NHUMGzWsEbj7SYokE/gBk14eR
2Fnd+lqDXUkNbXMYcc/BB4CqC7mtxAY66kEihki3jDgQCOuvPS8kW5SuDSpwCWfR
keOcK86Qu3/NxsCSYh7enQ92rPggo1YtdF8HrtRhyRwzFb7yaAquxA0KU6UdWuV1
7D5ngIxWfSuuq8XDeaCGmwa9Vahi9KiSgvT35h/cPtWNK174gP5WJZKYVegUxJUc
aa9ugnBHIbvZSPgJeFkwIaEI5qA7yb7KuEBV1AeUy2mARrbPwJ8S6EI82t4gpf7S
nPSrXVDCPL3gs1JmLXgFdxLAga9JpqTlqfDkX7ux4PDMUuBsMIYIGpG23exPhBHU
9GtPnIApo/RNbc3bVTxt1+u0cwCy+cEW2gZegdp1fXitoTj5/jav2ym+yvSqdiqs
L/MuSGWUVGkpZuWEamlQv7ryDT4zFdWt2I6uRQOp0sSsENyBYiCoZtGooWCmcFqV
Z0ZT3QKt/eOY0pBnG5V+LnBQZ93I0+rLSFdkQDlKyQU0gKBBw67uYwWix6VrTfce
O67sj/2TI3jn6F1aj14VxOVR6KBG+EU7sDfEXZN0ocoSWtApS7sRjs4XUWdHYl3E
R7v2rWN/y5IN1kxHIz5PvkDSVyAhAl8Xq+UO4+c8QSd/yI/wuZZfSU++MbUClWqe
VRG7Fdtts7KdQ86c9VZdVz4IEQAOXWBLNw4rOBimPCFIoeLWQNMKglXEMUJzJ7M6
63xYhULBxjeuCCjDY4TtLKk4vlUa9dQYe4aXiMjuTH6YIRb08EZbBmSz+SU+ld2j
nnpRyGW8A6Xv1akpZXuXGyQ5RtFXQYvtimu4CjbpgAt3fq4mZGiC9Yh0rPqBans4
9XmHq+iJ64BG30qGo8hvi3todIduVWswpAozt41XYNcohyiU5vFXOTqp69zTdgHC
xrTz0gLOM3oZXQ92RIoiivPhbZhcpXWEiyADrl3uuTa92SeXfTIhDU13VVrB29Zn
z/hu343jDwIW2F2GdIb2NUyJgNPeFyufh80ee8h0bH/P5bOUIZ/Bmq5qK/b1Xs72
ojJ9LOPITXK4kdCImvUh+CPRVBdGGO9oQICJ7FfR4CloBuHUOEjq5IEgOAoJ1R15
HpzZo76eqUFNlS5F0qA1T7MqTT6UmsemIi/pnH+weydK9K3Ln9Ol7RCO+miPxT5u
DlENalH1Ac3FXPCOzqrqF3VLFxtOn8BHA+S9zv9DJIRs+HK8lYu9w24Jbc6viMpV
Jm5KUEsGPL+uEGl5iuTbjZOEgro/uuy4tJ+Tl2+VaCNM9/OHc7v0DeX/K73wsIDA
2IWOupcqMPz4T6Szu/0BqjCDySeAhC3EmHt7jgS2TfalSzW2D8mT0jK9AhbEyg6A
sTn8Vq9e7IdRrtfmL284bz4yDlWUVEZib8tpeTJ+fWpPRtk978gyHQ0D2xklvvgo
Ns6ob+Aodh41JzTJngSVPc3Bi20+G1UTxz1gte3g2G8ExaZdIbWT2ph3kRzLls7C
uiOJt+AaZc43Y8kTJxwzam3PULBJ63Sx+A1SkfzPeDfjriwBOLHBAfjg2ly+yI3W
fzN0Ly/eTZXL6lY6nNynWwylrgdOWii03Ss3bzhqo2qba9/6hnJy1+A618UMdDVJ
EiEe6bGjLzW7jC5Jav2dQAAN8W010w29tKThNZKBXTkRGJvdOAY4vpMIf8QzvJr/
uuGAzEN0ZNApRDd3/bRJW7X1WZ9TM6+mUHD4mjAeZhtVJUT0YZQTilFGwNBbGlZ7
z2kRUxEADYaSzyE0m0yLFvOVQS59JMJRoNwjqVytHGHthxUQXXKdHTcmlQ3Iora2
qHeXn2Ks3+IAFQAiFGYYAaKkegjAJhYr8expOiOZg42zO8wxbH5ukQhUye0RFde7
IyjON6OFNTdl7nYYTMJHtu2zDaABtOc7b1ECy0L6hM6ZpPWQo6AGj3zRBpZQTU11
ztTRq1r1YaMGeSqH+BsOYo2cBNLAQpGyLlnZHgawRVZGdKTkn7BpiXtet+pPSBSu
AmuQ44gu8rfsSjqk3pKXR5dNjoNe65TYeuf6WUrsWrguxvdj/yFz2Ku8LKUYUepZ
QFTksYN6YfuyHbfL9KH2ajk0hkKLZ5slicOtUgcOk7IR+Idmbb6PTJfFCMWiqukT
cIpWy0zx1ZuQL2At5dlNepkGkIMrEIQ1978SAgjS3o+g75dgp6IpR27y8Jqj+q/e
bk7V6pZ2WHqxXvlOMEKihZ9IpSwXy0LUOxlU9HEEgXVNwfgu57E9P8aFh6S8fGRd
Nj2xcvULtIeSEca0whmXqdSDyMeQa55BqYdxaewsUoAE8cvpitxawpIDIYKcO5JQ
qIaU7BZZdpyW3IYHTuzCKFcuzKxj0FNz8PZXOKU/y70SJxI6Me4HTPzDNyhsVwmy
GzaMa+Lz4CzSqhha26fUpgrdikJylYlpD7uacMPgMrM467GDe9kniLqrh8iGa1mK
aRBx4siqP0UavLsZcz9aYJwoeTLzckS5tY2HXyVZ3K1adu7MGglhblUu0A4pxMoB
bzbdn4c4gVHQQS1rqTuSp6gZ0HjXz0n/QnRJHqBg+9RxnLbChg/y/43zPJe0GyyK
tIo4zVZBwdxVXjwsyz3+U0n8CnYj7K3hFFRuV1aeW9+upVzS24q3BBt9k1laP5cf
+/0wdqH+KdqshhCvqY8BuTuU9HpUcYMMhIlDFsxT6+oSl/WROyRt2q01U35tyfdk
iCTBwWR/m1FQNl3tFK6x3n9SjkWSViOpXNmiUfi8Q3CPbw6qM9/oN5qGqV5rQK7Y
OcjjzRCRgAQMzLM0/sj1xD4CQ5FDl971D8hbYqq+E1oYAFJVHcB7PkMNm7JQCpRe
Wxezbz9vI9Q6Arbd/dTaCD3xSc5tnwmPy3LCqoTOxC2xO5nv8GWxDHYu15vEChKy
kvVmmKdPGXfhR0tRzCpYFmdKZn3GjzLe0Ckqw3Pj6ZmRjyZCv+LFlAH+vxJzZcUx
dxgQoSsQ6DWyP4udi6/cA1Dsvkx2bME6QUBJnMv1WkWChI+fysHSzdcp9hcoImVU
Gt8438sCZMdTJzY9KqYfL83qC/lWVU2GxstPgrc7gLSJ8eTlIbDb8iFcVHSXPARn
neVh89O+z0/8L5Fe/+NJbbksld6V4PhloN2lX1m9t43PgUADsn/tYqlNn77Yxb0O
EsjERgum4RTr3+tjw1sEtYHoinePrtkndwor+kYc8Fg9O0mPr/WHOqI0w2J2OLRZ
nZ5yj/7UhwK5eDF7qBZfEfyWMCiBWxZzjgAeoGHQXAmt8OgjaKZnlYfaj6UYMtqo
YxQM7RHpBCV/KIvsq/GDkotD2TkmqkRG9hyne87GUTXOxYEwb6vvrQyKmhuz1zD/
3FTGVj1ypZv83fYiVLCLBQ+Xza2lNcz+xmBGZfZ/lxf5kZFpT6vNkt2M9QkpMpF0
4D5O/ChfYBPRN0J5w0p8ApeE46+xi1BinLnuTi8ObBwxfq9DkB5A/M9bPkWFvYU/
gT1hD15ZfAiZv1c/piXV63/tDadq+BSsnKQn0q7Hyephv6bd5z9QhvW3gxolKzAV
+aaybiNJCzWa9Z58RY6tD/r+OlqnzWAzwZvDfaThy95M7cOeBLRerow4fC1s9GMz
25lO68dB7OTX+0ll3fLEwdGFJk8B4Db7bWMqynqevcQp+AEoqibYzGB0n0hbDvZv
H7wtkkVpv0kmOyTd2YdNAMpO8aa0djRLeJWqZ+mCqi5Hyjz5gTjhEe92pvWB0J6L
6sKt++67U8mSnpzAKqR7vOZ0GMQ5wCOuOacUSpbmZSY/BvyT2ARPHNiPMbuxjhaZ
leq7RHYXdkRdFmzWh0RRxiGtopmIbrvYlP5IDi/s+5pBz3C2LuFZ8PEGgprXFYz5
Obq/8dgamPoONiw3kgh+0KJ0MM8ryBQsnIXk8KWx0Fgb23QMjoqHrTMiYVBpc/gm
U8FdGwdZDhFZaWVMqxaxlrMXw/uYC7+RyqyEdsjeWB8xwVm1dasU/QrO/5bG9fDB
o46uovI8pOnDB3+s+LMWiN22WHlwSrNNDtns6thZpALsB+ybIItYWFjtBX9ilG2q
Qi89xM2Pxe8ysfifR2ANwe8dkyD2ZFpu+4pEbJDUnpKI7mFzjNK5SQupMlxUMG2i
lD/r2jYfYNXeLN+zLcweWA+aqac1iSZElxs6cWk3W+Y64hnZogxCJ+sidxGSUEJs
kbUt2FoeNyiY+lPYsM9LrQeaP7I/mi75q5Qeal2s7j7yOiR0pNH3Ivgq491bT6+x
coNlSIyWqViSUmbIYA0myvZheMTNX5p2FadB7L3OHGprcgQblZwl8FCvn5p49o5Y
GgQq+y+qKM4w/GIYgAEMCV3WM3PhjhD+vAQ3Oejgkn6xkhNepeGnFeMDM7TXrx4y
e/as7Y+9TGKfWk0EIBfby0JEdEnGcZSIG6D5jFm0t8s18m42j93vXY+oCMaYHaBg
p3cd8VxQChrBaD0WYW1gLl5PaCS7LBFTguFryhgpXn320IZIbu1qU4kSiZecP6Bx
CbahPK/+7nZdIRykNw5TfnfLzcJZHxCoJfsNnz8v4tpeSZ6pBOl4Jj4CvVv291Mk
L9wtixGkBvdjJpW+HNboeHa5phWMGSz7toe9+6l7VQ5BA0sG29VM/AFRJ5lp8sCm
aR4Zg4/Kug1FcMw1Bk9WY3lOAyS3lVLiAq1c/OKfDwompcy9JnbJy6CjaBR9T0xK
/c3wWvDXLp3B9yCVYE2Qm0MDjXJpM7GnQ3ZgEPOk/C+Nlv1XUMHTB0nLPD04G4UF
GsTOiIZRosNj0uvk1eNMESeAreLwgRbzVfnOC1rJIsTHwvjC8Qwtp5DPnxa6dRl+
v5fpBrEyl4oTbqcXwnp/pMILfOkdSUC3EbprsFMXaH3GhZUYgZJb2uP17+OmLRvV
aiE3/yDJglKBhrDbQASj1u1CEAadvVXIPDM5BuOGlZYkM87UY4MoJhQAqLbDTzWr
uL3AgKxngGhyKK0LVbJhrrA8SO+Kg+2klRg+xPokYjmwjYAHt/bCgBLGA6Kd5lCI
8XmXckr7VMAkozezRPilJvYKhIVo3WcZ7I26PJiKI9NBsq/+SKcO3cZuMqYHfqE6
ZboEcdr4dCG00GRxYwurPNlWazjLbwqxHgOZ1cea2DXae+1hRwL1IA07DuCmystV
8q+wJvvqY9WSBACuBTCXqvgJxxDCpZ47ECtnL9QrrX9oMtHU4Ktzcwx1B8QD6FPF
X9GQAj3LajcnEbu7UYQL38VGkxulEGE2WeCWxaAwtEvMSAbPrp8ixL7b4/R4O8IG
Xfy+jBEOa4U9S0kSURmKkl82Py5rnsN72umQhgZBe1hw/9B61kp5Vxpw+daQ39i7
27vtbTnr2TDQ2CUOE5uq4Lqus3FtfVE4ANqVeWC+a8f4yaFlI+1Hmc7Y01A9kc1T
wL7i8Hk+Lc56cqLBVXiHrqgHbCsE07DLt1/GCC50ZHF33mDbn9tBSACvf9u0Qm4Q
EsqWPARfqKN+1hDJyDmWkmleXKIgnp+KYSroeFqyfYWPrXBwRAsUV74QdFcrUjNm
9IYzutqWfbEtnOEzTR0L/1VQapw6fYGTPdp+ALP+vubLP4GrnU6WQm1orTxiVbDi
y+6saGr37sJdBhQhUG8p6flhrLkHW+6BBQO58GxKZ+v6ddPh6/v/s2EAdZHyEjEp
uq+EufCtXDUKq4927Cn4e6gjOkTsNth33Jo+1Mp9ZP9hBXvXSOAnhu6Qgjqeonlq
qDxrgUgoBTge7lIrZj8XXMvsBtherLZhgpeNUb8mfDy/C4eZaHx0r90VGH5nIHvQ
xwB9wj+osFl9IMlfdJNMPjcvvgDKzGcZm6GkEaE6VASNyPiAPdNaMtHtfwQXUjHq
8I1V9s/OaNQFVZX7LeKu2i7Qx1+GiFST5+Rjs/utHTy9+C152nR3Pt+L1lq9tPwW
zSajHHMs/svTrr8gkLgFTbUK0rxJaNKGysQi4az+YCU994UZo64G7p1VMNczWvRb
LeD8/VUQWuWjSdZON5GWWA7/2FbJcxecjuqXa57wiaGqpOSWD/sYRpFkhbkFFiia
66ToLJVSosFBdTwlTA0g+s+0C6cuGuPTWEhafTU4iXyKrNi+VJxlZFuEWwkZmt9h
sFviLDTGuwZsJC1BR7ws/tHMA5So3pI2vL8LdDn2d8N9H7BxLZFpulTQ7W/l3IdE
9KXRNpdlnlwkXcoo6MlRNV+7x642B4pLiM7R84xAXJnCudI8pxaTnJu4ThFr3qQF
sBiADareiEw7U5uHbzkx+wi/fONGRDQUZTmOmDjaUIW6r6ObIcIhGFsqS0wLXKYR
9Y3k1wjcTYI6mO8c5rg+cPqOOKTbh31avuiIEzFwgQ30CBvzycgDjKdlxTEQLpHI
nfC5sVIE1pKpqrV6c5PIm5Uqf27o8/KQtcplZ7PUOtKppzMH/nsr6Ei+IEu7U3sb
05Ps6ZiRDkZdc9VeKm8lbcMT4B8mGHHDCw2C6xtRjnwVq1orC0HM+k8BGp2yLLwH
5tO2gQUe5eIl4C5CZH6g8ZZBiHKl+NoR1Yfrce4uJgO3M3reQm/z/QdC904UW/Pp
+hktjgLjNgpaKNdTG1adaNAKztEBQ9GhOTGNb1YPkv8jXYgVRlPeqc2dQ3qTX5FC
OhAjMokku3lxjg/xuXp8dzfIqWW/pG574Uf4SPaKu+o0WjjWqgzFzpc2NUaKOC2k
48sD4RYUhRM97pEDD6EOvweUQT2/qjbfuBMHDUByZ4Y87j5OTBHIRC9lgE+sK7IK
UNlwP/uQtz7qN1FOLAhW7Ar8z/iRSCVtM0+6EvGULFMzjv7HLzYONuX8N4GPB8k/
0nEqfhp6xWEupygfjKr3H318dwENSiBWp+0kaJuDQSw1mHnh31DXn3f10N4cfWPh
jN+MOK1AclpqMKVFIfouMXXcvimJBC3nKZLWQOGkdrDYvA8EORwClEM/NR8xJtxV
xfoKS3YnOTk00Hvt0gC9zS7WH9j41VxNqjYFD0oYqZtTqFhCoG9iJvehK9IKlOq7
/KXFKMmCFaUOhcga1o9T21wyoxqe1V7Q3W4VkWPzK8Lf4SEB2SM1hqlJVHgOQL51
q+dfWzbOS/7EpY1GIB1mJ1+txr1dYi+CV9JBPYc6MBmOkp7kFWuCZiDRKdRXsJJd
NSopPmMWH+VxwKVogeTk3ms81dHeGpSwTxdIXhlLOOaSyQXJtb62EZrYK1tys0Xf
GpLotu5AKFO+GgbpXMPWMl2yDTD1P6ordoTC+PNTfpnSmLAzsMxjK6gT6cwrFVOi
w1BMlmEekQsYYNz9BPiyZmDODJRuZH8HJGx8t7g4RTdoDJOLTTIG0QOX1eDcgxXQ
089ENmdN2MJeHgBAJQMlWnSCv7wIO415jkq2gN2DJZxIG7FzmDpcGX2khx/5GtQH
tkNhfywsi7jLwRO+KfLSa1FutFVoHD0p8E/UaD3f4d40B3WlVZl5rkTKCuFEItHT
KvzBvYacEknjV91mEfTigOkdKTL8SrXEPq2qJorFxSFO5mr5sZfmdqjOpIF8ZE0H
GXDciTo10g8ZtcodkkKs69w4IxfbN4LjQIytBqx1Q4CkytEOSysTYTOjpHzB5DgG
iTL+A4xvjuyW3FzruUubpeoTKFOfLro76FABHsiwL9iUDqW29LcbhRv70i3uRS3r
Rl3pkYDXasF2ixFqwbHh5oyPdIyx3i1J9Pfhp94QBYN66Laoro9FCvFEFTRm3lsq
HTtBk5WSWdtLMSQ+odvzyyq7D41XYvFGg8f/hFmjt/T59Dl6f2SlC5MOjTc0oDI2
ThpHwL6F9d2K60w3G78lv+fd4+11+lUjnhv/tGvowh+PLHl0YxQZt4L6oH2gcO5m
3sI5XHtgSDdTY0kDSsWqBBEMrM8Y//+bETuOpDKCd3Cf/VhwSLBT+LIijt+MMLxy
1Iy5a7zBoQm36EN5MTvgeYJbMG3Z4w9z2XF0v7LvSCh1OdOYYxOAIfAbvazdfHC3
URAE+LwlbL2hXNZMwG0BL5H3u49qGPPpGnyftTSI8DTOBVJ6LM5cOAwuwsvIVbv8
M0x94H1/7uFXBK6RPSIqBrlG88zJWGV6Ysd+qvF/oFTzbf2zkL6YKLcnV0A8tjgj
OlQIB2SpGpU6MU0S8tmgi0kyPIV4ul+bcamq+pwEGl7gxQd/1hzoJYk7Gi/QvS4/
9rESEnVgzQFICdib82PwaX/abKjSAQFNL++qSXN34j7nZ/PKe32AR4g0r6MpC04n
xwyVA0bkbLYf5AJDm9A0vwABEfEuLLLn+Q3tLcHSLnB64XVDwHEUdsrveOY3wxfx
aCrmuZTIOh8Gscw9EseYNfzTsehNjYOFgJG7qZsmrLLxeUWfZrMNW9uOHNnsfyyn
dUFhfmF81cR9apMmXXzHYznIg6lFkaNtn174E4nI+AIpT4n4Y24iQdBNh8n6Fh73
E8zMC/uXOWaM7DGOv4xqERNj3j1wzWguNnfE+7H32BnWNY93ol6Plcmr6qC1Rf6S
2+IDVtWfGa2Sz3j3/wco67cLMbV8TOwW2pk8USj4ULyGkNljhxBJJ/JeK+qUWX8m
HQudZKW9/QdIBJFrbSE3Rtso8AN9MYPeId4GE51TmHOc3y9ZswI/CWqkHyIWOjWO
wmLys6pJGNyI+3hC7wFAX6hpOaMJwAW5GJSO/tn0AxVG/K88Ulzt+gmcmOL5PqRk
TvMN6QSgLzjMmjfDf+pud+vxHP7g8b9E8RHoYvbJWdZle+QRzS0ZmrJY8PFOS7TI
JSytoFlbH2vhv6jQyE5IQr2+7LZr2CYeCl5YTyfSZpmINmJXPLGEvX6HogeNwfUw
Td6xnOx7OtXtNOa/apzi7iyNUOF3sQEd2QeFA6WPxMdXyXFCmr2e7d2jfakuCgwZ
r9BAQTMYPo65SdaV0dOd5edNniu+ZmGb9mdCZ4bKy1BW8d3GeDXALSDXU+WfIaE9
4+oQnZZiwvMFzF8twWvWnA8ntUsqmMToxY+HYl1t30GEGNbR8QFu8SBOeoY7wfSl
w0FkWF5qFdi89aKgf78F0ZFTjCyiT6zOqeWTJGw2edl2+KeWV7n8+DphjncPY8pO
J18Uh0x+Jj6M29LD1Yj1BQbww1PF8B+6CcLXnguuHKwj2mltYeHZg9mB+ZfjAnaR
Z9WuLxzjhXu+x1NaXvH7TJSlP7SRLK34a/OjWzBgh8au1XEviS9sZJi6javvZYgW
EfsMQlS5O1UIVpTpZdLWtR1EIDAWUH4AhmIPsrQL4r5eYfrZQ3p5MLUqHn7ND39b
m+k67D1P1VP26JJKTtgpFp7+nD6qtlCsRLCRJQN2SUuAkoxLW1iX0u6S+uTkjqfK
3Jp1AZYhujq0N3l006eCw7Z9PSFd/luFTHk4mLF1rEr6Nlt5Q9qvnWHqTDsoP3E3
pu0uTZ/n+oFjG3W++ZEh9LGvmA/iefnjLo2Xv0UA0V10OABeqq7J5kO/2d1PAtrV
umju6NZUxUJwRwQ32wMzozx9iBtcV/mUhyI0I+OJpqSl+B3LWde92CnexMjy9Ira
VRxWz8PFXTreUfg86ZyoLSu+AWuprZTPkclwnxQ/6WH6R2F5O7Y9mWLoAhCaYjsA
Q4z8GxxBq0r8AeSHWI0X8dJ4c9MvksskAeWXe6rFO7RcDtOYd8tM5hosIPyVB2MM
GCbfjl2jiUbxkhcM6CfQgAqDb8/SAO8ipzwlYUTSUFKxGwSn/Jlpt0ZRboUbvYd5
SrWrs4uTM9O83kIqnNMsW5+LsDlix7opzk2mTvsxNqyBaK8XH5qiaxtoglBMJAO4
QYTvqGPynkib6TMJrkCNodfrNu/gWcj6FQNFfKALU+ppW1QJJlO9djyEcYrYC7q6
1kwFm+sL4cVDrpg1AYjsy7j7+3pxvXQ9ZguyJRTha3j2EWiM3vSXB232iy3PFocy
uLxCrS9fMj9QLWxhHtv9ApcniHZotT7dRQ3l/I6eSiiIsgCl0oe6jZqbTJ0cRnAc
8zUUu1YwtNX77RMR6I3rjRtGlvVUU1NgGxy7oBN3qssBip+d5FDZ+VxWEFe1lzI3
0cOVbR29vsX68xkFN5pp2Q9E3DFicySMSW8x4YzlLvFuS7c+NvU0gY5PsSiPjLZb
CEppgLnlhZK1WuKHb2HQHftupmil1STCo+C2gaO0wumqWGaUMUhgnulgn1KYHWE9
/r1aET5fnZP5c9/4GTGVMzHWnvGwggcoQS2Y1k3pg8S34heb9m8nAU+mqtMsjIN8
KMcri4Jj5uqk5Ou2Jogaz3zDothDS5Y3ILpKY+qTZwbpbp7zx6iaZKCq/xijZz1U
2r5CfUgfsuni4lHVYW3rH75+XqntTKYjTvcxGzqwUPsDkkovdtnwMP54T0+mhW9y
duktTjFdx6A0DhH9z3UzObX7t0YVWtkGzf908qNerMsASuWa/yFvJbryaTmZ0jZf
U4ycd2ab9uqcdGQXfZgdwk7mnBXY7YXt7MiVI55D+4HaQ5Fm47KQ3VNDKlhUmgNH
QcvQgEIEgiqZeK4jlQOPnFjowaTRkfydkIdfWJnB2TW/XgiJMVLbSNV1+dLk7lps
oHXE4+viDF1qOIfeWwgl2Zs8ssBcI2YmVd4tthrCFgN5P4EVv8Rl8IJcKKp//90T
YLPuh8ELF7Vs5/8/jWt2pjWZP8sys2n440fX3BcvhzSad6wnybaRGNnVa9g5GXEE
+fc7p0Pk45zrF0Mq3tpdzktals+5g3Kvvfi9ameufBVhuF1HBciQU0Je2YnyhMey
SWwM5fIHnC76kZmElq8WpC0D3vIsMBE8XCf/xp0f/84UYNSB1a7ZzwuDDT/KFcnX
mnHexCvFTowwdmLuEMfJVr+trB9V4xzrjAj1zlvIDUEeV3v80HY2M00xjAypzHhp
FUKWjZdaKT0hOM/d6sd2svzpJn4+V/RdUYx9Q4lrLF8ZF0oNpsK5YhgAzBV7WKrf
d9bxbpsVKsIjmeGFDGr+keyU3ijnU//Fph25zb4cBxz9RSzO99Yj5h/Mh+yOBo4U
J41SLdhGn8+j8s4tiUutmpuDtwH9lrDF1lQlJRueZRBfbh3fOy4RirwcB7XMJ/de
33tc5KZ0Lwef0QVIEnFGYHnLOE/opb4oOQykX7aF+nWK564Bx9cpmhdAclvu1ows
ZOBYfMAxgu3m91vSipDUHtWmxfmY5e6GUo3ERG1Gwy1qsQMjh+UI51Wu3OlbpMJi
6kXmo28UI7TBq9W8oD2dtgUipiqfCThcUgdFr9Aj5jAxpgfBzCt6ikKRTaWJnT51
jkplk/PwClEpXqPbO6mw/sD00UyR/d18v49ACHDkfl2eTgWRzMWRM8BfVcy82gsu
dI/x3ZgP0Ggj24YuPXIe2yDJ0wNtLE8O2BV+T+Npn2DSklFPeDNsXQaPk/19sv2y
iTuTbjLL36KcipwYa9dV+bHHJhav3a4tkwIeoSqr0imZzNliuiwtoP7hF4p5jNl0
VZWDE+hg1yraVn9o1QbtzK2Z048Dnw8Ed2XYcbdW8mYvTgDEpfhT2+CyudLS6CcB
AFc0Oa7NLhmcZcKWOw4Y0gsG3s08+wWod4jtDVnQm/YF41o0FTJDJ/+c7UZobYM9
eDkKbPBydzhsVwo4KE+40bMOO/GRq9tlkmOKTnTb7vn0YLy0lFHkVr0mhPrTM+xf
xjSam6yR7eklLxJYLAtqsxddL8Kg0FW0Jdbp7I7CN4r7pzx4irKEHIthgiYRWRsz
7C5JFAe/ux/a0/2S9toxzuRGRmDOkjOhHoRQ3s3lmlPQKmh3otc+Aluvfc/VBoZA
Bk2egCRAmLI/h5OKbTu/7vgrOszq48Z5LjeWD/2YKGQjsbwT86kz1tF0BVi+tJYO
RFjjRwFNbfQqJgI8ZSkyHo4hyIAxsKM3X+GDaitqWlkrJ2/iU+dGLUWot3X8mR1U
h9WNNn/n7uCKa0qch13KX7noJHyUomc/3cO+xx9bD1BvCTtNmuzSeyJzTL7h3HY4
tvlJWNi/JO2nI0J228e5WxoqzJgUtHt9R+yynUJ2MDtVBc2NG9/hFE3vMY076PKF
kAJsq5dDmo8VvNWhSYtWRg0sRd31TfUfRM8TwFOyHf55C35D7qLPYhi7VRgXNlTP
GegJkB4YMop7QwWpljs7ZGnlyAbQuwre1k9NYJCRUSCEQTqejVGCZ63LEpmudAeD
hgIS02WfbOM7VKpwkgOf0n/67IPL/lrtKEkXXTasdOqZyBr0LXxZ66puFEaWqPvl
xvol+ghe81ei6+l7o+BeN91hy1mzFfuZvCcttdFLGrkjTTObn10A4BYO7M5z6b0/
8/ty93T7iTYyg/kRFYqLLh0wLvYCXvpoKiJPrxD6rdxY4xZB6dq5ah3IBFMSM8eg
5faFt9hxOJ6jtOy/dfE75ENRy3TIRYxrAvMveNcALxOgQM7vLZ+pSgp3p791QV1a
JPFMrXO+b6o+5GkFE4k5syCKfG1VL4a0SiAgaLu8HP3tgmwkihFlt8PW5pr707BA
EsjTCkOVlOd8le6ZQPAOeIPqQu8PgoniLJXuT/m7+0xHRSoLrwNSDTiQDCxeMFKe
Z2mmtp/zlGhYhH4oC4bkdUm2HNlo4WDD/9Uo/pUhoYTwROMWq2tzhTq0DyVltvB+
L8Ew1/UgrFMI3Sq9eaWopy+qZX9vSLPgMGngawyXvzeb4BpH8xYub/TU8bjNMCZH
hdX++yvkFilPOcnpw3Dgj8L7R8zET3QiPLTTnhQbbZselhNlnmCzTMHxnFCNWRqK
K391ApDKZEcTU4MhGDw0HJWv/rUlFZbJmHEz9m5VRJAS+Eezi39Pk5XkI6aYDG20
leHcfhqhWCVX8RHg6A130FMTNVSKDkR0JUZXq6+MoeQpVl/+ux3u0LZji7kZqNaT
TPtqxsfIC7U6+Bi+qIpRzx1Hvd7eV4mZCoROw2sM5jVMFBtE036MbYN1vgwhpU/G
EXzcJJ4prC6dBqwu+3DJ8QWZUJBgvV++fX8E1z9ehZ6HR35APQBycKteF8vCwm/K
HyvFlLWWgKzaKaGSdmnvll69/dZtNOlFF4+ytQkNCN44FrsxGli6g7YNGmrsseYq
UanTacnIfpwpjk1kN5RoWAu/jtVgTuZ5l6te4bnlMu4NmE/gmqWLbQiLrI5J3zwp
pr487GL0gIyot/26qxSztN2Kz6HtfQ9Uh9rUqfP0/IJrZeBPj8xaSsZxV7Yq8NEX
3pfe42uKw3rwuU8oLnp+JHhLrMjaHxOo6w+v3pBxOQp6Yzqmaa07oIfV+JCw0z3Y
nKY5ZNS/vCdO05SnnDZGu3wbnHRzJy76DJdjFAecBXrd3BAfQOIXyTtMLAEeLCx8
J/LB3a//GjdSGxUcg9TtNiIVwFsY5wmH75FcaHtGp1MyVmlPXKazJGCNoRwJq/p/
l0SyO8tD2dNgMBe1b6RvEss4A4mYxvUJsFUWf6WuFnnlDPv5r9cKeuF2NVQxTsEc
bFnWbdn0L/R/d6xra6ZuB6IVYI6+CNwM9EN3aYJnpIRX4iSBtLX8eJA2eLCnUTJi
RjXXojaLEMVR4m1fJeI95MVhqtMCSx2RlsJPS/uEjOcXqsy0P4iGagXKNDZSvMbJ
41pPRlULRuYrBk9UORQ/XjKLeI8q7L2L9JCLJy2GaeLP+Fg2j32yHFeGh/Z6a0ow
KmMxjx8MVKTP2VhhtBt4N78vcSfGkqQL1IEWjXESY7jorJczSXN71d0nQGu6UwCt
SWMnyz9Twp7Mi2TTkQ6TYCUBJQ8zxwPebtC7wlAKN38ZpWatX8zhNaq/kSgwTGuo
qvVWyeXH9P5asZKof9FGN5vB6jkdpHo0iX/rNROlwtjUjpD2TamhJNecDjltL+c8
UbR3fRbaOb4kaDRdY0rFSH7Fvm/O6GLaAJDTWP+vFATMj3MHQyCsjk1sGBkbLoqg
I5UAP4JN/Koc6Bvz/ra5SaNNOiQcJS4M09k6ftSw6HXYaAATXffpuyw/WnFmbMr/
0JdTAyqPmR8Yjub3w24U6mmk3vz3V1esBgztKgBWogggEX0gNIwiuQ/cU3Bi/SRi
E7sqg4HidpXv2s9Z1peFzX2rjthfWmZtqieIgdFNgDtePK6Ne7uJa0T8nXJIFma0
MkJEGYMX7zPfkeA1YOiFAzTqvr6+IPYW//VeZhTWY3aTIFlG5Glp3pMb6YThh2x6
Xm/Eg7Z86ed8wOUK8c872UUEJ3WDWi1QcwZ4qmWWq9tUCBCy6tMFYvAdT1sQyQTA
G0DzZln81W/R7VS7sHQ+qdN3gVnv6W0cejtcx6algDb4h7Id78KqdXxO7LSikbcn
9VnC+yeVt5EqSBXkeKTJEHnL3oIOen1kq2+3R+l3kKY+HEdR3uqe+TcHs2oEkZpS
bPpKEFBrFhS+HhttX1abCV18M7Y9AG9tInkgosj5K4sqvpcqkdiObvVo3bR/GWkI
zCXt/fZL5eBmqf3nvx6KJW1hGJIs3TdbZhNprgSeSPhE9eeBanbWPq2kimZprnO0
Ily8j5qPZuUdH2I2i//p79/i5wg5a9IybLIBL1P4JV9qvzyEh+1JLxxhXO1LxyFu
FHK7RHec5rC3fGY8ElzyaSoCzRhtupYZK5m7qCZ6ZlhDHNzeRe2ZD6SjCCXcvS5v
s3UmwlFtG014sIvSHrqrK/B3nfyNNGUuwrARFS9VVzfmeK+HFenVFiPlVSA0yKXY
YoDs3YuHp2qIiovMhSZc8ri5fhS7kqoTJgLoDf2Cvh4HX5hJC19KrYzgFwfErY1T
70F2T487ZXnvRJiQ/T3HrEI4I5vB2/CmJGJh1SEycl787xj9rOrykjH+Uoo+MRDd
8XIUMYe/CKCgY+hdvESqSjMsLCqkM+cDTaT5XKhnVP4gaKBIEd96G92XMGuBdsCI
nEJY6yKaMaExbyVcf0Lb4cxGSHEw8tyauCpyZjIV9M5urpzEyWhtqH83LQancpkO
k2JJVatssB31TEviM6i95/KqhxGfz679kd/b9Je1KQ/iMcTIn6gwbNEnOsjqR9Md
i+cwTZDfwAFgDb7rObaX9Y89Ua3bQ6vuOGwZThbxsMDY7xAEClGNQVsB69j5Q0z6
FyvWZoIOzaMAMF8odcspv7p4Z/OLGxeVy+MVm2q1wkLEW3J4uxjKtOCOXMy6H8e3
z4pyFxr+iNJ0pS/MIGIze/4AMZ7J3oFf16kxgpcjQvJB45VFnZtyfuqccfmNVkUy
twhMuMSks67rZRJ+q3/T2I9uBYnL6r5MB03zgTwVVXM9fLYXkjhI9LR7+ksXveKG
zlYkX/4bAk3BiaVgOFrnnfcZFUDyHkE6M3bORB4DP+AZ9hwEVm3shKSJ8r9ZofF+
9WhL+KpF4O0htbsNmMpruLNF98dbjQJnxI3re5zIAI/pRe3aeIUbYZYqK61qG9Vx
Fj00zxkI8YvkL65bl4mEJSMeDRFr9o+lNpMhe79JHEF+T5qCLVi6/xZS75FAT3qG
J6gwLzpvKY485bq8cRJRFufV1x/Q32YaDar2+7haudA5NtZKx8XBigaHK/g0d9B2
/03oBRaNFwj+EYKSUQ89VBUDG84QE8w0woXWPXDVK7vjD8QdeQlwZ8g+0OAVADZ3
r1G4c2Is5goti8yykKRQXp0a3JVCx46OHucG2WBMore1DxYanTVfWlYRaXYEGQWJ
MVSaO4O/SbszmswXv8h01ZsIn0uDH2zMkwsSw8SVsxzDizW+MR9nZwGCnNPvdG4o
RnORpS3M0q09Z5oJR6/WUsLgsYbbSdBqhjKvvfe/Jt9rrm7TDDDDwUDCwDzMkLxy
FjnQlvTmcAMKVhd7sw13LrK9kW+eZRK36dyzZFwqjdhKHgKHwcTwH8Jq8BAtusTU
2bgxaUSJeaHf2ICxLMxMoTBrnn3+UcRDtTwPLmdAnWxzNSYix/6NDCMLa3vzlmca
B6guq5rxiy+VRzuRXB/7vheD+F15LhUyT/6pK37kLR8AX/5xKxovk7RWia9D0pSX
naYTqCzI6ivlEvE0/BJCBieAk1KtxqM0AfZCrd8kFzTyjl2BmSiPrn5uNVECT6jC
RhTcX0CmhQC0yUPrGMIZV/FwmfGUHd3p3wv82La2XPk75qXDoAjnCKoL1W6CbE4G
md93LtmjCYc5hVVtIKJmLYrXDa4KBUtKMctplMR3C9IDY9VLgMaUeHNuaZQm6g99
4QUEhlyNxrPnLiA7t1W4f+s3CnLIPrYMjk7FujP1t15aRUsR2Em+oas5iUmRO0Bk
ZcEu2JZt67hQEr9vofk0QP2jd+mzf9UatDx+NMiPVZ9Urp+gZYal0J+VdbEVZT2y
SIT0n7I7K/V/0lpPSg8ocyYo8iQLbbY9FwHHBT28rk+knZHCBsrUkdNedpraTsXS
iH3CkcdURFl3D3jz7aZU+1Zu17DPXAwKtEW2o7rlQh7J61iugIWRgIcW1OXnZV6R
PTnJYFSbhOCvq4FE0Acla/q+Im6choHl/XAq0uzllokg2sZeRmzmIBEDNEdY3q2/
QSBXWsdQZltGQbl3u34Y4QTDz1L1eN+PzC47wMZ/9VaDjL4nV8ftr11XLo4iPage
KIES+OsPmROGonwvZCcx2fz57etGbTrDsVko82nArnKJwy8f8XMB1BkrGNhQOfnB
wWkp/17eXrgWv7x7Ng/W+RkxzL00ACJlcdvGP/rBk4xADZbg8IZpOlt9dExT+jnb
JUX1NEOI8C4Zun0sn4NQmPqlzfDbr+Jql/FYGdG+cBkTwwizErpJXpZHa92e9KXe
NEq2lAN0B63ZWEHS1Fj9Jg8nFoXmUwy+HljhzxwcZRlb1aiYci7+Ixo4TWX1uj7X
9ur8NzvyCS0e1cXZ4LaWm00SF4KsDE/udpQg/YskiCslPerBYWZ/idYAs8KC8OL/
T5tGia7d0spaGcQCiU1NKYGmt986eo/y3+d6Rm2CIvstAD+x5oHrufTGDbQqSErZ
Uuli/DOmZU+wbZCK7ELlf0WZOomMUd/mNPBuBzRehH7XEVbWvg96V4n4oWilus5N
r+HI/7EMp7JDtPbBU9qAST5wYi6ZN29l3GBUxZm2zp4zllS5A5hOo2v1bXqP/a3x
5tO5pgcQFiluhAjee9mFUMgodx1Iggznvjlak3Q+3yYv7CD6Jjz/H/lb05ijah3e
vE9URw7HsiFdwbL/HcjMCsNVfKs7IM908r2GN8DzyZY4qnyeoKoS6O/tAsR0ai/l
TV97ezJCRE7uS+Z/y6B6ncXxdi4HukKstMXtI2hRGYZI1IN2m3uSgKEXtcpsrnc+
GvkcIS+DQr7wvR7LoFCZPXbjmjpTO3LCVI/fBBIwmRRerrRSW8eplUHi6sk9iGnL
FQ6lkgTuULi8I5E/89XCKt2tm8FT86lhThI6PhHhnVzf62pgASLntu1w/JSmuj2B
hse2rXrdgjXWLhy0eHHoRtFP96NqTtNN2uQRZgCItzRoWMX0ncpEEmQjndW9NUob
GBDseG5HTzoCY5d9clLhLYIGQ1Y1iV6ED/6DFH/JVq4zcGxR9NI2b+ZE+zGvkATF
BU0gjbzIW5v4xrCmHb+4F3IfDHmymsCjaJAtLhldcrYe8l+xziII1Yzr071bw3L0
ICLbSOM8Q3CQdVqwsIoXt+YsFj+q+o4M0GQBP8j1B0WgKMxD7L9UThA6M38Mft8+
1Qdn7EAG19vEQF06HZttM8R/5vppwXYBgW/GsAA0cZmEonSAZYR0S+UMJ69r4blV
StL+eMeNKD/FJ7Fl7Yt80kjmbrfunMGHypcy5pH7eIvz4jW8Th+RQLSPsHw29Mdd
Rzgzr6lVu03tAkapRWLtbaceF1CvY6+K2PhTiVeSAQJDnN+JM38Iog+tHoONsuyF
4qK9m6eCHRMFfvMACb8kI78TmAJixpW+NTBEX95olkBC+5GfR5jQELVWS2bLd6px
RzMjyDvYhI+o9lcqPK97WinRsOx1awvf0PO5nbodUY7eKt1vt3paCmdGO7I+lmCt
0D+W8xMs0yUnkN3stdn8kgFk6u6fUGw/0hGiAGrtN5pLj1n829qk4+BuMWViFhz3
RHc5gCvo+e4DKkOyFesRvQgm2oP3EXJiuxMjHE04fAvgEK7/s1b2Pbt0mcLdqAyC
YnEJ3V2tbPjCFIaTua0EeHCfIb7iGFeZxl5CzYS/OJ3VoYx7+wsBk3sV6LoyX+od
y9B4sEYrlcirdc2vlrWnOpL+x/5imEiq2ANxnVlE+RMIMBPlcBcYfBSIqm6/9hku
eeV7oJPeE+R0DFETLyG9YApGP8CibvfLKd2q2L5ep9xd2/pqaRC6/N9OVq/Yr7Uy
6eKWjc45tcQH5JiKlh1cltr78JP/Yd10gKwPKg1kPAN6jS6fy/bYfnzSrUYjfkRi
WNtlssWRQUuqT2XCp8AVA7J9ugUQ+Y0j/YN9OTIiLO+sLhvkmJcr2ODZTcy/sYbz
HxJ5Y0vLFEc/03eXNxdu9u8fhhCzzaObtspHiSL9PKBh7+d4cd2h2ew+pmUW7lkm
pTKwfwW1tV2g9R0WYQLRR18Ub/siqjf2mmAvN34EIOee+I28yST6yhB9bbUMRY7c
7nVJ8gTg4cZKi87VG2/3IJ29IoRUVkCNC48ATBdP2JAXYGq1eCZRyDbUO60Z9gwB
5Tv4Qoaeu5tuwp5HSUk485mGOHElAaYHfx92ZQhhZkCoptRzwPtmhKLUZ7OXBdN/
mrX1lNGeguymaLWk4kJN6eD6yxpgp1LdfIcpEw2ToZCyOOunOZJD4TVVEaJZgf09
fixeOeUUFbyD6akm4fB6e5hHPlwEklqbAhwNDXTVpdTacBQCntoRynRXZDDkapX7
sp1ujhcTwbUm3HwlqhVCiqXLW14jTAGx77g2qOE+m+Xv8WHONkqUcQYk656jZbBq
5a07U8jK4JJxM3uXObKPCgh93sCsyJjM5KvsNK18j+xLd16+e8z7CMfBYOAniMCL
7WgI3+/qSephUFyv40l21mkEIHUixuuGiq/l7tjsUqSPl5dHxqAvKkvVS60pXslQ
X4S/qc5WJqzedl3N1KqPgRBZg1KsDez7G8VefojlOKcF7Qhw0/9qd6m3G+r+awoQ
vARLFcUUKQyQ4aIfj4MfaGoL2cL8z+GvJVL717PfEjfKE4yeKLB4xMIuNMm4C/nb
jI44kA+K4G/iasOjZc4+8KerLVLyjkVpjkxSPCNoZpqGU2PVHLAVc38IxZl10ARS
vQ3KGuin73lPwyRDL39all7oT+mfWzghYr0BRYlhCbSffV+CjKOoUn37rjAdRRBx
i6a91T2kR8maPb0cOzl5mKlLRRAAkvd1OjfRQvFFn17rIjnDJ+sVMuyWSnbxaEn2
DSmwO2TyJqkuAjNjx8pjf0ScfLl8XbnCfFTNxs9uIursjFLIzWa/SW/M7t/HMEvI
Hin9cGbuS9HkzUp0uHVtBqXssKK8p4jbryYdobm6nS+OIhzVPI5bolsEYxi0i2Uw
9V44cy2YQ++eTYGz0bPqK8RZYRdI8uqNSQ29pNdl57aqEN1AsX9p0kBxQCYbcIAm
ZcfiOjshcehZm53pAmeQuypuIvCKLWgvw5nC5Bw2cwEFUHFk36z8P9aJGIsa3ctD
2+/l0Sp1WtWhQ9HVwnTgMTu/rCLSxJqa/IttqrKCsBUKB+XADDd6lcVm53qqyBr7
TJhw0TpbDViksIvNRMFhSgC7606zC9KtK31R0uHEO9dS62e13h953VlLjDpbo4f4
YHhnz7MCWaG6LK84vf+YctSuTo0IYPQMeumfj9J46Cw4w01lC+OeVbwOUQRraQ9B
yAUWHWgtE87dSfZospmAXGwyxYluzac2kCDCkUa21fb4K5EkfEh8NkQXi+jCa5zv
hADmA9XDKxZK6+jRNhlPwFyFTuXBOTV0s0Gg7+nqnpQA5DMb0MfOgt+KKOoyT6Kl
JMzuIOFFlZDrvf+y3Tqrep5ylQrQQjlX3U0G+0+nXS5yQFQZUbrFUXXuNbpW7w5r
rLym1IGbSAwgZ4Rbcg68qzyYXkJqjEWWiSTYL6vdWDouJiIaY+SwCxiWhht9B/zW
WhyG/WsScXZBaMCU7dBK5jgFIDi2uruwki8thsP3WTCj1bHkqsk46Q/z7GUa6LUa
2KGbdrmj/XyhUoPmutea+Cw7wE9sjND7fVRealXc4hbNPOBB5tX1E7WwffoCAl0C
xd2UwWcD6YgbzQt+WrjD8NpGH00uJ0EUrYhcsilRTNAZGcE5cpEo3aK4yYUfJL5e
QBqAQ6liDKigUj3wVTvOBOcqnnViiaCmTsZpnCLSDdCcSyb+10ObTkebY2m5Innk
/xvsw78wUocLOj8V62f48mPOTEnW+0mH15uVdW+ohnfAGfeNCRY7osIFUTmuwYT7
bVM19N4TuMNiL3XuwSkpd6NHAWQ4Ph3lBBgXsKTiulAwVh7k+i4tWaesya9WXE3u
FeTn8MoxLuhabSaElTmcwrkur9i4rzhbozsfI6QXglH6bfi2YU3bSVbYE1iI2w0z
IMg5nm6jrjsjY4KPAGTN/0kGoE7MSd759+WIJvuazFD/vrBKmoWcurKrZxhldbSE
kEqrgUwvJYET+T/NRn0dEK+A1DqQxkFA8iE79Simg2y6QPN7wvfm3qkgiTgFlRH+
tH6A77Z+EIFaxwsCirii+23/lmvvFj4HhxdgNil/9iXi99//cBmSU9kfGHVqpgNm
Sw5xmURCDLzz5q/iAeBwAXDFPRs6ya3h1Suvq3JVdCIqskh2PF+X44BP/eMWbopf
WwakYE7rkkNZ8r/J8/rvHqb+gvIyb3m5tpBmwb3UUt4DiVFB1w1mZUKp4dyEGDZn
Qt2MgJy0qq7SIr2LyCvgGTW8ar8kzq762ExMjB+nQZjGQ48anPt9/DZHNnZ+OXeW
9XKoAzMqItdrCvWIDns5NQpLYy/MkMSnXKjwjDuxgrJJGPyaHUua+sK0BdCSxyfJ
NZ94OkUxwCVtvwptvDMRF20GFqkWsEq9Assv5Tf+N+UiEQygjywKMU+a88RZco2z
lklBJzhD0n67/sxHCNQ768b5xghJTiXkI2kzN17auuUtgMoucA4I+TFK9s8h/erh
Hnc5RlNro0ZmtsAh1KSQ3sgfM36XE89Z15mT8Vs+57yF14rawuQ5D6lnRUKvri00
6MiqI46hnszgFE1gx2XIhVdWlTsEkmd3WqH5YaVodgolcy69yp1+g9pKGtVYAaOt
iZj3p678ER4vo0inQ+Yw9p4J3XcRay5iJAckd9Bp4AhQMu6MfxA/Vx0xH9lig2A+
Un2FBEfc0xUKMgKr+2rhkiF3KHgOtF+fqEzI/sbrtHAbyuu/xs+CNIhxiUeKYOPG
xuneE3TPWyUT0yGiqYa3G4gLlVuhMm4olUklaX2VimXhsb1PnC1ezEeOuJhmXR2a
vHWf0t5gXgQeHk4qBfolRNA53KXym55sAA+/UjoLnFqnmQ5GbqugTaxP1bGO6vRY
g1vdzr+6r4ez/DMmuQjv2lfOrphO1BKDbJW55LcdaTjDFfxi0dGaZv1LYEdY7byp
OtTvI/rFgz0oRZCQLYyyas/9+ro59WKuRmgPyk1ziAxMQ+542iOo1NRT3knx5HmM
lRl71ul/7y+1mqmmV1uvRzFigIkJ8WKBZXcZ81RaUqIng9lKL5/GGXzLUEB3pngL
PQ2AOJMGVecZI26ipot+ezUHknGf+2MHb48sPeYaGl0K7gIt1AqwaiXy1quGjH53
7hKRe5UZGl5bA/V02I2eG67lTIhnMt3/HDEKOy3AslcAiakw1geTAl40ZK6EOula
Zdxa9LLpTvm+I8GQdLAzp5sbMocYcz9xLe8eAc5U7ML2H+dEttIdzJqWB4mo0u0P
t9EDC8sTz2igDCd0pR4MgOzb9iMvK5wuhqH+qf3wp/Naqe1mYNrlt2hjPUjOOuxB
KVIxHUCcy00Oguvx8nsP4KWzcrnSEWwpXi83+fFSp3bh6CKpd1v+/iDRJ6lVA6ZP
bHLoCfahlTzP+WpXO6IXZ/uvhKtUNZzQm4wltSYAaKOl91i5iYnjFUgEGZNBi3/D
/seWPkza7bGH5NABE7D824oKQg+ZEUCzY5pitcVe2TW++dvq8B4atbf830K0Xszo
QwSleNtSPav8DL7+itNcMmNd2PzLKWw/JiiG+DlcN19kJrPIg1DEkGy4uZtMdRpU
1Gu9Nz5cWq6HQgSK9BZMt+gUWr37N2beXvZejR9NOuLcjBnxk4Rbmns3aLTXGsO+
VRZAa4QewJE/XAhX6bWpG+rTA+fzN+M8m5cxxZn+KZIsudGkT/fvJJ6NCDJppxmL
61hFQCPPKEcjszESsQC55hVWTGRBggqA9qVuEyQLH7Ud0YpYJeiDH3bYqiKgpdS9
P0yg9QsrzhQxGN1mdsD2+4KPni/Y/O5NpkGrXcPHpuA10qsDJascoLIxQOvY7OIC
TfvEUUiAAW/Z3FUgqtHoma6b7LWDd3AwR2n9P9Pk+gbMZ308953E/dW84da61/CP
EHI03YMVz5W3sbi6SPhwTImX9ziW8EiHVvSHJEUZl6KwU/8LbuEkapo8m0G/1dNS
l0146mDxeNvy8dswMmPI7LvHZTYuyQHLqf2yVFvy9AMM8UwVpOqBsm6wpP1tYHmM
KGH2bP7x+wlLq5agNpUsjWTNWf4FUhLw/qKQq1smpWoD5XY5VV3hAzgRLi5z26JS
QD+GwROMsIRXfejPSk6Tzmy65IWtO/aD3YUe3tzto1rY5K1TYD3FePilJdLW+D/R
fjkojqqDHdY9Howe6t0mxAck7FJ6abmf1A6lik07lYIIeOvTAiF7Ysddv80BeXky
OCx6vSquNYG0dnUZtRlJ8s0W0PjiTe8kz26t9Chh/TxgFmnx4lZzh+TuXtJTdX5s
W7oa8PAP9/9/0GvJEm5h1TFDoMcMT11KrR2VcCiXf1DkQocmzfjJkErPOupWq9Be
X0DeJ/yA8h55P5Pg6AtKbf79p1KP+gmDXjoRQpZ2JF78H5SLLR8c/NjuSQmq5hCo
B2ciOPx2l5sSMaX0tZmxZHh9XjCJ0EF8X9ltmjopjQURVPHPzAdbdRhtsSkfFtSx
G9+vrcmNtYVxtoKkwET12y9OjamK0HURAnZxLWB/znMnUzfbU44+EYc3P/TfqXCP
zWLsTqAHmbmLiPHj6DTYOtng/lIt3C1t0d18KXZL+o2cVkXMKXBmViIyj7fOo7QC
mFHz9ERnaUGyt00tHzHWiPX4f6wl4QCfGzm1kkg5bQjkuKJUtYNtircnJ3hS8HGs
+GVShGT9lpCEb1XoNQwUGuuL4stcmikgyX/+l1Nl69BkDIxNzb3MadgTU5nnmlsu
VlxYUDlZp5Pa41A36mTU+fJQ0PFi6qzg9nG4xUaM6LBF6/ABL0KgH9A1zlck0t9p
T2Y0GDb/MgxMoMCQYrijcPrTw/EJPTJRTOpnSxoRu+rO4WQNBl33SBnj+VepXN74
Q9mlBG08MNLDzfF6a72MbUAmcgDX768s6AI5nbkm0uARDB2g7SqiJ7inTuLmn3Ob
1fUhcc7UliORxdkUmkwtdhV+uLqiHK27EV9iBOT7EIozYYTV2nfzesrv6QgXGHpq
CST+s7uOVXgME5QbK1d5imGnVvdeTwMW9ipTZSxAEpfacMXFYNLoyj6CEzYRu4OQ
FmG3HBq6+Bp46Llumg3Ei5xzLvJFjfGwbW7AI+gwjcp0xGsH+M5g+zraBG5jWup8
37PzNMdD7qAKmoiCBMVk46yeceTQ58W379BnitRdEf0xeCjwa3rWEVkonE/XlSIp
vrYyqIqZr4yeqVL3Y0HAJi3crXP34xspR7z/rAmXWdPZqT0xn1wPqo2+tWI4NWq2
NGuHYJDQN8tqLmJtnhmgG4ceAUQeXdZUsT9dhIjqF9DXE597p+apwRXcbCgZlnKM
iZTh58KW2ymnwPTdtowSWa30tZBq1dZ54+nIzLL5sAcuHsZyXCfUdjybRA1VzHGG
aMXgBEnXkiw2zCG/K7y/5m8ux60twuWCriY0V1/IYB+Wlcf7qNRQGGhiFPhdmVid
qmi3vU1RqpPW3DYlByzeEN9MdUtYCajMBU/GhbLRQLXIB21m/40H7xAdNCMBGqoq
uSOajPacKhYdQxf3XGO9T7lXhxRobOsGY/DsN2Kd/Iq03f+s2r+VwYWG+HGX5gdf
iLlxBwVqD3Gscf+JG7qMap/+ZoIZrDryos4T2uBEFNKiEPBOO1u/uJgGcS9JHpHC
bBUkUWQzn95wbihuOn+JoL/ofkYa0EPzmLk+7QEVuUnw1j8AhyjMP2envoPWd8lu
EQba48PEonO3JirVC2PGDi5eeSOynGoCtnD+hu4MP12q9NdBG24g+ehWswnVHOH7
qYXY9sRPQke8b3f8hVugB+Ax/c4iq56X2Fvm8nm8cjyTGh3EpPI2PhHXd/ZKzrma
+HqxpA+s++h5+zsY6dXQuf67PwZW/Vx7Y3ZxYVCYnRCtEhwKGFzCyvNzhXeI7tVO
oNaeEFR6w2dZi78Y0Sc+90/q4M/GEMcb3pLbolXPRSPcucX9I7O/lkcjCxHKnGgO
lVepS9TRq/UKbbSD5/FNYShNYQt246BfZSu83LqX/BgBvUigLghCx/WBI5zTKbzc
JCzndD5gobxLwnurvJlg2OqOlAgZSljlHT5goMKCmxpGFuLcCTThT2wFPmwcbK9/
PLk6PRWpYPFJXhJlTEfHHFRU/Zr7Ttz3DfEk2RrEGtvuF+fmLfeqrsmqbXvuWR1k
vEJvg7V/tOE8fimCIwg6Ug7evbmtGxZ1OBNWjNOwIu3sEqTqOAYMVCAay7kGo7Fc
4DW7b0iZ9XtCeybPrxXxoMSxUhcoWz+2MYpdBZAoG28BbePYr3LkKVtGSwUrrsx+
UIHzqwQYmw5mZodhaq0xX+SYC0MJgBLG2QSniFSUymSAjHlpkEhZCogKH7+s+txO
Mm9iYhKvTpHVKCi58x62IRY0cN6G4iAkMBl1dNEpQU700NTtQb2CM+L/7Ke1rFZc
6Pg4PsdJ5ebtfinzQCMQZLSLNDABWThPw4/UN/lhPgsRC36VChrcE5p5vQxwDeeZ
R0Y4HJ67Eb0nKKHi0clG6SZIG4lmHXFBK9d3pAg/wLW53/UFuCfRkXVOLFv7KACu
VgrebiW08Li7SdSpkvlxvrL+k9roP1CMVk1+4rxb8juwZmIfDZVJzbBE48NWS6Sh
9azw7U0aMHJx7zykyn4Cz+f1Z35QophekEhanHD6U99QN6vo+eS3XIY6HYohzcac
DjbV4QtxnyYmISD4hhsk47LEmM5oUxpwJ3pdTI15kdO/y2wDiYJSAwCKonD7l+LN
acrGxA3TfKgVBYfX/tea07Pd9Ow4wBCIN0ak01sO60DGare7pQqL8vH1JM6EH/S+
k4i+4Qd535hWd6/cTDb2dR/383WC/+1Z4XuhMMgWFo0VbStHpWBoX5Yn26lXw8Wg
Tox2MdLTIcTpmZJkT0EFr7Alx2UwEyjn03Gl7aRBzZ4WKwAaakmWxZQB0C4u9MjL
BJq43pDlPeXvyJMFgUXCPqi48yF/UXF+gnxmIOzNdKSoDaUNRzVRnGFRDnJTgUkA
Zb/JGD8+/DrmGKA919N2mURWD9L7RyVFA8wyn0L2ZQ/VIMUittD2uEkDctH8XsQ2
ffHEphNeYEoieMjhEFdiFgE3y3ii6nHrnjWca6OiAkbogBPdfWoMul8uXGtsKjc6
fQbxMZRr7t+//UlkFpLkDuRICkAYo4sj3lM7rCZNEcWy1UZ+WdauXIuvwqK0ui12
YRdrM+N80iLAxmEOaa9XP0HKrgJt6bZNLUmA/YYDf5JoX8r1cHVhe0ybWhmh50D/
l+ovufuzHligVqPugFSc0aeUTX44MMCTir3ftIHzctwscBbNtb9W0SnceK17DGe6
tZBG/N4+oi2eNL6ulOhBb6vP2UDM1SyAST8Oi70omZGzcWYLJIXAnCEF/WI+EZIk
Wu7Hvb/EFMYBd8OWfApddQfYSfNWGKD3N9fjwfJ896CmxtB31nBhnUeirJI3OU/I
I7Ld2N4EZzMRFRnqHQYeV96vRZtLwAiOhV9ZulYksNiRPt8vOvfg8qVeNEKeLiXI
5Zf3uxR6l/HAQP9HrHJLyTfrY6CCtfn1Dg++JgE3sdqzAe1LnbE6wghDsNN019OK
CnM1lk/9JBS7JlpKkRDnYjVlk1EqWNbvbk5ZKT6dj8JL79PdlnjBwI39caK4pDJw
EedkgLG/4pKflAD0IAHxBfkIqadKZrzNRBn9WxMkEJJZHA8tYgUPt/qUqFPJGArm
ILK3m5i0J05RLC9SRzywTZoK26m6ftvWIoQJesjWeLkskO1nDjS8aLvT8q1KSONH
JXEcBXExDafk/EQphn8UzN2LMBR8RZpjTM/z+QjglsLzSA1YrjvgUkwu6O3qd4Ak
hWJIbJlypxlIUPdRs7HddICjcm2teJDUZZnUjbapxFpTPtjuOqeLDtfKkGuLKGkc
YuX3YlYU7tqaJSyTfMZOP/h492cLlP5VKJjYa2rkdb4X7eMC7Gmex6g/HtTtEiRd
0M1jouksFXdxAYd+aNlPKItH7unrvKZbC9c+ARMZku92/1GWNsULbZex5iQeFOgL
tf4DrNN1ohdGJNTU4IyBcoF3GGe4BHABb3Ski9zk1tRsFRno9st/qL3Ua+Dovbtn
ow8Y0bVm4qe9nkSbnpgF3LVVmADcVlEhriNqbbUxgYVe0nXypeXK2HOqn8TBKtpx
8q8pDBHeh9sdPdE9mNTRHjR+SJIK58jOLjlJlF6e3HdikMyF9Q1iOFxGiMgm7L6E
hbqqeY6frlAwMoCWIFI63NurjJwtdQ70lOlntnhxt9sot71j1GGB0VJeb6p6OBaT
GeNJR/Ek4xfvJnGpS56agQKcmksr8wWpOXK75AYjDOHjW/RsvJIxTzmATR+kxeR5
uKQO6xckiC/RRy6NhtvTklK91dUzv9Nw51iXYlnSW0Hu/AZxLNpU2ivogJKqYwbV
ByCK31YSHPxIi8/Bc1E4I/CxvmEzy5eLjpdZNUf6xGNFvVdzMw99b77Nz5oOQL75
xr3dRQZNrWu4yN2SH6Kx0M132PAarAOHFGX7aCvJDRMm6UcQ8bZotRh9AeCBD776
mgxdRhOUJvKQg0DTph2Bdpu9oqduTwlGZEsZoOyQctVGWoe2EnUNEVe0zOT0rCx9
BaiR3Ye2gdQgC4DPvT+qb9kCshI2TfLpr7NtrCNXaF9WXDKnHKCph6ZwYPE+hbd5
Hmm0bsiFRLS7mrYlNFkgnV7htfe//gO6gwJcynWYXLtXj8eD/AVBPF5VjqR1AxJV
I9wG+5SWD6kVR8694Y3uksCXm+Xh9AoBKBxDWI4W54+CrH1rNDttxgGIvKEUQSz2
tHTJ9wW4cShevkKEQGRml15DfXGF5QMc6TzOKy21E8xtmJUDiXeMEAHqeepegfIX
KR7p/B25oiisUyA6hrPSgofxS3U7LyG5Lo/0FfYeiGxiLcKgHxZZz9w2estEy8FA
xpMLoo4kcKo2SUejqulNoEh8Qfx8dpCjzWzENZPsDLEeNSsLA5suKrRj/8H934Uf
V0PTxC+WsHO2okRQAp1OeYHy6V5IEk5ZriNu6BoC4PVULk48vWQgvSyBvyZYdRdZ
VmOiykVNOtUta2gD7lYV9jECgcUYKc/GZ8SPb82Cq/PTm6zmnDP/xypFsadxqbeV
j4Z+aaCbdSQnz+4cNc89eKFKIF42QixViVPIwgri57tjK5nBanpXBihI3l1YydXS
3v2ZMo7Z4lvoMoCf7als4d6qS6ADDoPcKFpM1fCrYe6tUPvEZh9lzgJCvlmZ2TP7
UyPJeA4HVcc0tQgnRiRDAiqJfZyek4a/dumXhSpqtGRhxMl7fK2TelW6YjOpgonX
qZK1alRD3XoW6FK4A6Flo3rgHauXv3Ig7TTmym6VSQD6wk5pa+iXsfiFC/dpGiAV
rpGF/ANKz8/UNaVYwnl9/pjk+LRKTg31DNQ8EL0No495licGu+IkbARCWyzxEXlg
/n3j1ycRZiBP8AA1Q5NhD4Khze/Fv6R5JwBhapqbcdC7iC4DQeFO5KT3EZOad60J
1iXAUuwLcpdE96QO2e1dQvTi4He9TtvZ/KXj40gn2OkWmwDdor5cFFusGvjogagL
a3H86jCjL5dE4JGUzEsTiZCYiVTNE3zhWtagccJ3jVyTIk3GzBKY/V1kLOxBrMMn
5mcIhMigY+fLYuslw+fxU149fTSoW0NfIKPdjN6S4qg00uXT2dBekU998NbR0Gv6
vVO7cw4chF2DfjB/pe1eU7VZkbPkH6BjpcdBc0ThZndkHxZ08kfd80N8UpWtCKMD
JzqwHbaARcZ8lhtkSzDV8e8/QPmTQ5YwiUvUKHo9v5aOU+Ir7N/URqdT0NdXIMnQ
K+HFZ6CFXYR9I7qH6vYlylxldbNVSpOpU6VDiqdLpHQsJ91YmSy3gacAJ7yGEEzh
cMgMvUCF8AE7aPwSrO62Mcz7cescynjpu0cnQmYeq5khwSRKeXd+JVTHIAKTVhAk
CUHjER8QcGvHGMllFCVHCaLNg59du7jMGi+uU/mocfZOVQsaFoaVwbwKC/bzb10J
6zp93hIQDsoMkGAMwX8L5ZqpDiOU9Lx9yuNuwKl98yi0Jf40yyVliURJQwLSy0ah
qRYUaoADixoagcm/ub/UYK8+Ih3d3Ayb1t35KejCvc3ukNX7iA41pRMnlhAEdGbj
YE5Voh9xI1TQXAPkEksAv2XyGfzuWdUJNwsxyVEFvZ651BppeDUJixAPvT/k9KyR
ciW9VZD5+knbdFAbQi/Ry5UtvtM2oxcZ6NEDCP8jXavA1Ab8SolZBEr/k163E3on
GqoHOvfnzCjZCg2qyPh6qcuP/t6tHO+Ib/EJ+tSFFoLMiqV43Omgs2QCzdfgeD6S
dfxtbh4ELZ/fc0Jfklip1Qyr1gMEhRoH0ze0H/tmd2vqnj1Qr/8Ri9Le3qRrTf1a
GDBi7uGIwlyacerhado+FYK9e8Ot+1ZAK4qkSKTrxsuv85ce+LogbocBnh8NItDB
pwOwrGQ21kPhFWAHpM6RIHNwjRiFddlJ8adS8vW5QLx52+dEn2IzaebrkKinxInZ
2V5cjoG0qAQnVIslBLrQf/atLX21cGGsiRpekTsQ6vBhKOEs3bBHTRVRmgMS89Lp
3LMf72BvHN/ypMCughgXH3rrXWiE5XuRAUsmtzNQ7gcPP7IO9HxpfLZrQU6a0lIp
GvV7oc4Ppv5hWCcFozLIS+gKbE57ncQ0KeUDTgxH2ts/XEzzoLSwaAEHtyJ+NOmU
PoovpxliV2V5ZH5FLBq3Cl3ZjvG7Ao18767wzjEHA3t9JCG5OmsrH0lMis68RBNx
1UJHlfB1+Trkk3VqLOmqu8gcOoIvSxRSs3av6UQkWMOlRYuZ62gG2PnkKs1AuxO4
DPt2WhV2Q+NT13xELvCs5QAtuud28vFmyrNvN81wpLg4R1GdUnGDCxpqZ+inQfsV
GviPJ5x7PUuwSZoqLT0kXTGefLhPDM6DTKocnLyitq2s7TorUYd5IcCNILI9218e
AjsuA8706rLaf8mcQtMJ944eqlBwk5etK/toveq6eGzc54xmSeQDJobu4p1ZD/7v
zbyVtAephAlKBApFh5sfDqEEOU1xn7Q2ET7f2SiDzgaPNaJ5TSGoATADRh+fONZA
JLooATQh+mpm8y3wsTJDEgELcF3hwT0BsS6WPcCipsZxlqZZ1l8i1KczqZmZhFO6
1PqdH5n7AVZKrnM6Kx2iFvE6S99LmSGnfzp1FRrM0o5Yk0P/h8FnQw1ApONQEoNh
cEBpLLyUrdjc838cTZSDmQayW+EGKD6Cu/S0upQbiQWZXDjHBdwkHNYqTOgiY6BO
JkSqGtG7g+7u/yuM7QeVLcIjtVMjKA0pLCAwdoQ7tDViPpJ3INOtgkwL+PyxqwrK
SuH+2Gw920MmavnTyF9U3OF1AoMFnmBnmeJyUhDDy/KgFSkXjSCShork5jrq59wl
8UQw/JYaO2hxkV1c53IAVzjnWaRY8VS410U/5gjwmiHrRDuR6lKDk+nuufO57K4S
FWDNiCodAeCTidpLKsp0uV1NMTcYsDduK+QXSM873EE7kdLuq+xHSNDjznO2wYew
k1Fiwjiqw0O99SzHCMCTzVGjD8svOeORXUyHdmsq0pYbXIoR316cV+ePxfQ1VQdg
Huw29JN6KBjAhE4i/I51oJABbvyn0pWsqYJ4eC4NFerBUWQuNKkoMLS5bmPzHapH
egoLn8OJs5TXNONUbW2yz9eOj7xqmWWyeSjbElJNjOAg5hG079iLe/1+dc6xeYfA
RVicH9XxJswOdJWtvFxkqIDaqiApavnsLMtLt4EEpBAwUHx1ufsxV56O69q+hhBF
nDwgm2ByNZ7s+Um8PJqb7hrRwswwk7jR2dOnorx46BvwWqmqsb+xcZe4pTc0Jljx
5LHWqyqShwWcnPE/RbMGc8rg7A+dSX4PBI8lH5QmgTl+wqwhIlS3HJQuA5aMbugx
XXZFIE4zfN6at5xv2LUXEkJBVFKha/McpxoGvwVSE3wX9DIKu2jU/VbgUxvG/o0y
vcktKp0z99NSBsRX1wir0vOVIduMy6NW7sw7DoaqHgl0VJwatp0DDssevn2I6n2o
gIscHG0Es9dtXh3tEZ8IJ/pjRRoaRYq9nZq8nBH8n7QeygsNzLCGWYVCp85zfO+G
aQJVj5zlXwe6lkKUs9QctyZcxJcDwvHVoe8tN7zM5DFCSB0J43WJxhaDnt55egEg
klRusKesWL5KCjK6ctB6mmeisDclp8iHHazSwC8lR1X38zNwWnvvmRra9wS8WOrP
rLjkq46ebxB+H8FtVEGzrM9UrBilH4ixLi9iKinZGaMmkCGfYEIDqMMErHvqdOLI
A+SGUtW/8jBTqPCEIZn32KYxM+ZwWYO2EDFNBWHtNCBAouk43Og0uULTVxMkihBr
nSHzgX2VR6bJ/mG5CO4Fk1TwufdnVqRJ6m8PQpla+yDHu4ai7r9fDcjjWBy6/DUU
CPsZAavCu/IsCfLT5grKNBpVVQc5mky8MGbSk8vrCN3XVI8exU4a5POlDLAp6K4p
CvHptZb4K3vpyb3oFg+EaUUJIqo0/gHCy7P2pyjexjjXESo3TlZ7IkENraObSuyL
1zr0ltC7/IIQ6DrvXqOV05nGxjOQyVQBL7fnLhHA4Bj0MxyFATjDdH8rph996y0H
tpOJeM+zAAD81Mih+Ij31sVudYevjmxlH6cKX7e8z45HhKxoGS6hL4A+YqFGYxJV
0Tx6d1WZtL0qFj+1W6Qzr3FsStYhmV6flUIveWkOPFzW08Snd1ww2TaShs0h4Xno
pyxeWqzFMiI1fYylIukDdhAd/oHm5zrdppVh5NfGg79w7TldEfuNvBXcS2fD3m8v
d9xPGbcp90XOwHM2qwz6ZF9J6H+jPu6JKes730n1XSKTgYR1k7D7An/8opbrOyge
rFKJfAbPidlYIFTXIqlNXN1xs7slXqt+hCceI7LmIcZEEaApNq5v2dMNw0xQLbev
h2/5PaW94l90n4mAqcoXOhKoFUwYdUJADWflMbJZ4JUU3ErBGwn8D7EurwgDI6Rp
/qLeM/GbBpWDVYMPMJkM9LkWKHSTMUUsRNucMQpyM6fSPrwGx2+TGWbWfS3YxWOA
YWKXLUQ+xUBtqHU1+Da+7Q6C9VNX8Cs2KM+AkFSEzTvzdijhTk1N+agB3XVXrP7d
+x2laThhuPPqADE+KhGE88zfft40G0SqfXEkiI6ljbxsLbrmHjYFTPRiWn605eXh
aDNEGcYPxWUtJfs85aIjcBfoiRMp04MWwkt+NOIudvZ6zzQNuVi/6uqJScR+AIcE
AfLFvd5cTN7R5U4RsGU2J7EWZRhyIAcvav3pRXjyN4RdODmWx9o4KVaBL0KRaXiJ
qB4/TvafVnmNy3Zcr5NiCiyat+LSL0WIkixh74Koq8OEjlphY+Vpn9ujwGN2iHyI
i9/F9u0NDIibPIao8bvfSPmG3OpadGxuvh6j/hVLstFTVGK4+tvDUKarNnPUyKA6
WEqHsYFntztySR/fbsc8Azaa4iAGIkaNAwH36FLLsgxlc3NNc/PyzmpW/h//YtK1
rPFzF2Iow69mm4LyJHeDl8rn6DbWkqJAzpMXJ5dA0UQpgxTPcha0turXMEvMDCzd
6edma8mtWcTBQn2RM2j9PdL+muGo0JeMmWhkmy1tIr228OSawvVTlmS5tfFFE/dZ
/i3+ARfR35TNz8Rn9Ii6hGDbsYysiXybl+CSArliu7BinvzmWrXyh1aVALAI8LfL
lfP/PSsfRmImAAKA41Pqisy/jbxfgvBn2cwgnUee34BFw7iKCq9NjxC8PEMD+sEs
odw2bylWIfl9/FN66bRsvFlm9ke4rNRRvSOp0+R04/uCzLIOSffdCZ0cIe6ayPY5
72Co3g+KbQ4kTAqCxJAxZi/Ulr5CgDsOZfiahVI/61DRo18BZx9FlRyOgicsWo5n
54MFJb2eOqCTrOfWpLZaozKObviJ17df0kFA8lBL1F5Po1XISWIKWki39podsvTd
mRBNI3sUQk88e3qnv8jAIWGLRQHBqrAKHULYyIMve9DoO84FP56ZxvSgnIuc/PYw
UPd75Qx3FQ2P/zmvN8veKvSztdjSSpl0jHvQRCDK4Bdwj7T1wBtk4RgTCD+Z2vn+
U3W3HXuN120s7aaAb3bssXGmtELuYnxbzF0lVvJaeamnGyChcqsor0LDXXHab6kw
1H/jK8lSi6o7WtPNgQA0ZRHVkmRW7GYSeWgRQHKpKM5/NIQ33KvdH/mwAfpKXOvt
Sku9rxrgAkarwcvPKcnYuf7k5lWj1tjMkw3oFZpwo7McTwy2sWT6++TrOBnGzgM6
MiALf28ip0w4NvWocF7b1wYQ2Jm/Cj7HYiJEhE1gV4yRy9+wHPDueA5w6N1OU58k
rE1PHBXaVLJStP4Rg0OyImIVNdhw7u3JF8xggKntdFFnHRmIeptctipVmVp2hh67
YxX8hCgY0zbYO6G0bw71yxcy8jsZT28abXc7r1Ms3emg3YUpB0JtvFDf4Zl5ruJ+
KO1dbR7Id/+jg6Z7+mFchjG2uRObGBX233l6ub3JzFsX88meg0AwHKsCdZdAgc96
hawpmDq90hplHB+50VlMuqzVeDvJre5RRf2SqWu7oQMZ6y++toxa/XqSP4Oi3pBX
m1uS2STy5TuaEpbUUEE8wX8xS3WAUqLrcOazUZ+CYqvrF80G/ppHOm33qvygnNv7
8JkrkgySCkciOf7KM/rcVnBu2/c2c9cOunnmp+FZkFNJUvMaaEqjazC8JaLjnMkN
Xvjwee67geNAitjS+ve/d3TUU2v2LlYzXq/E6JHvB6g8q2ObRO1+Qb6YkHmY1Lpc
+W3rSCvl5Wccem/W/5gz6FmRPo8psI3mNbK60P4DgPbbXrpJQha5/j9yFV1G841h
oMjaDzz2tNQM2X0tQTmHyCE2y+QU/AaA2iLqGY+RAFKuAR2DusN+Sc40ZJaKOq4X
7G1nMjG9Uq65DSiPAMDLAlS49x5ILyNUX2i0NXmGCHVHDczTLD+NHA/32r1FYfE1
cE5l46NY49xZsMNVTGD0kFwL/GCDR8BFGjhEKu32Riye9LlS2FQ/WmIPHuakzS+h
Nv26cvOLjZ19o6bD07hi2rAF8OZi5tlTpFC/+nnof1BRkafsLMsMRxEPxUmi29mT
doQdtTx47bqZaZGrMH1sLSgmxdwoGoCVdBLuMregMM/+KDudYWDZqaODmfP5ibiK
AEiyNxiCHuN1uteT3UyLK4FE2cmY4XX+kBi4iRuydzh8c8h76Hc8Bw4w//v4eLFL
LygefHT3mg4xLTpzvJ328ubaOZXR1Ir7jqiY7qQw48I18fWfBj3j0+UoekskaRXZ
8RK72RsRLIHRv+ejo0b3NcFd4ohvCA/s9WHWtoGXbBC+0ooo98SHteT2SRjkbPB9
dOyaSLjNyxRFcAXU63Sft2DLvcuk9JbjpRbMhEaZGCSlB/TOHi0lHZ/d0RIdr8Ik
UQJDuRsI0DmQffkJ84JT98SFaPQcW/qt14z1mbzlx+PzqqcDpdSNnSRnzjg7QQ1N
rrJkNaST+GfLh36OexJVsWhtcsKs2r844iB1+sdCvSmhlgKMcw7GC3YUzAC3IiLj
cK4IZda2IR46GyH7ZaopzB4OrIiqwV99e8glRgJ4qU54HKaumoSSwCtUjKlvTAco
5gMXQfLOxgGMDjFHmAdlvOlEO+ZxbYp0EuiK719xj7PV8AtLHlXegGN+3k942VL6
It2eKGcVr+B89lwWphEV1zSVImpXOO/5iCpItVoyAkjzJifvDWESkS84dRPGotiT
mTgq365QsB8DH826lhwpUIYjWEOQ9C4A3RPUbkuSBXNNVHI2S/Z+nVo8+LUEKZQ/
QjF6Bd3MPr8/h6q3g4pKIax8DyRqrfxAjql6I/+oZDRZXV1zO828QxgcGaMcUq4G
pin3RANBcd6msOYcR9jX0s0Q+AMtpdfLVVY55p72mNKLzPIux8VOH3kE9MydaJdj
daFr/jVEFcdkzDSHjM7FC3PjPMsvf9VNkLrae5O+CX8AjrFUfi/K32wriueguhDF
kpCh93aDUsECod0lQLd7NxxxSvnWQ6NSnUOacxNNp/YA3xoXp+K0VdQ9fBPdxhvt
K2fU1oO+ewPkVTYIaIH1Dxg+GY3TxK1T/UglK8aBH0xmsX3gLjkHJwpf301vjMuK
WloCyCO0kYEXCvS8XLYs+Hf0mXC2YcyXb2ufOr1Y1DlZzEYpwJ7Z6rB+MA7j3jq2
UUu0UhbP61ixGuDHtoIovXbcCG/Znqo1ewsvgVdsWiUlsKZ1Pbs9ew6VHHenrN3J
y0YNsyph+pLCd2wUk2u8FJvEkmby0VqddE8g+PMuSx6YYLiZGJ1iqvirICd2xlXV
WfU7iQZzSUAVbEf5UIeNt4lpxhQldB0zY/Ekgi/31N09RAZgrbMW/42x7wLB/JbL
7za/hAZ+h2ymi6ve6bcP4s5F89uM5/oSU8Jo5Z1hN6uWqi5Y+sOJW80l3WCmbo2I
q+sdyPxHJK6POFzcENNjT3SckugTKFyGfXo0nwARz4Xi4J5S1HJWZCAGDgK2Pni4
Qls/g7kTRBzLIXgNLNFjhLV0Vyqua3IXq7rQj8L6UymxBuwuKpYG0RgHixgJqZ5L
EqdfhUe07wJV/M5B54nPVERBeTDTvVbw6FEjw418hz4ZZno0qPPio/TXcIBaSX29
pf7/9abyJVDvvn07KPcTzcnUmrVPeWagKEZO1eeHd9x6VojbBBLwZqrWruJLpI85
qCgPE5LDc26q+Z0tR32lwVtZpy5Lvn5enuFN2quMgPrZig/qkLh1iaADzRZiFcFE
oUciqLhkY1SR+Fd3Xdd0huBQdeD2cjwIkn+LGL93QcyQMVH2eSw1fFYGLYphNniK
QVIq5meh95wSyPfwmVjXukCN4zJ2CQPq7FKmOWsS8CzDy4AUBW7qvW/emK7bWg7W
84h4AVXpLNrukLv8QRz9UecOWRCwdd3/OTpESGiRxRPzd3md2UVx1lqDq1OscWOw
8WdcUCguQtsQKpn6oJVOpMxe5JVq0dyjFUqD+IodwyoRGBLbi3Z+9jgfop01nNYa
PPV85OzP9H0/brF+KzcHVWmcclDXlJJ1KIQwNHug/J+b1xfVxeVmu/oy3SXEcXom
x/9t9W0073us7zLeq9/tsdYUI/CzkLL42Ja69fQbM8Kjz7Cxi7gqAzMbB+/AeiIE
/6EdNlQ1nyXotKgiDF+8gzRy01ov9Os5flLafZVeeQxn7NDH0GIJ0X2IXsxW6Lrr
tz7JBCrABQti5irtiAClzQYfnOTC8o5nTqfK8/keMpstaWobPRxlIdHb8eHDheiE
vWLXXIQJyPa5zcMnMsoG5zDhPCsQQL1z4Vm1rkdaPInG1Mp+FPwHAAedliJ9b+hZ
hWZkGx6F8xnSxWNSyV6RWnu4JLnCE45ATsi6h6DVDQaqlCiSvPzom+78lNw/NnEx
moDNCj2HeAtd+IfrgmKDZkfxj1KvosNPdZtW5ZD5KVyOlAB5u5Yepfz6tFeI8Fkr
yNfTfhFFWEnGtvVqSW4YT5ckfF0MckInhDo+j30O83e3/iudk1YTR9VrMiB+u3v0
OvHxvRMYfcMR6hfiFdo5/07A2h4jVjVYYTYl+AXFH/+jE88H/RbIN0WDm3YrSiG9
+Sh0s18CnmiOpH2d6aSa4xurTha9nMwGi3fsyGHGcwU6zJw/cWik6S8GYHOd+rYT
cSTjtDXpv9Aex/t8HrqpCLV7eFRcAexLvkE1SMTVEUUXz3UoYgzJr00C53fW+N9p
MaSY3uDSRIMoL55IKyBz12bAlxFCkkPe89YQJlCenFkb2IX0TBaV1E7TilNmaNe1
cEYzq4Ofv5BcZMASjF+nc0JTxRgYaZvVQ2kbSH44qMpVoFTyigcqskxrf8t1Cpm0
mkxMilIypKwzf/7XqHddK2ONfr8yWk4gb6h+pdyMrtrXHNj8qlxq8Jm8wOxbp+sB
VwVORHie1jXFWvjGhKqB8rJ9Jg3gTMpIL4SJlvMtDlU6u68fS9aXXE0UuNB1g9+Z
pB7yXcuB2b/G1y6LuS6kOMhxsp/dLgI5mJEN/N6gtLD+j0pXDcARHpL6aLJdvkb/
hhfA4kqCbXQpq++Qw7YIqPIG/bnOgGvic8LTZnmbOGyyok6IVAhJVw2HMB+C/jq5
UpQtqIyJ+Guu9iIk9EG67f2xdcxB8QEe2ICt4biYzo1XWlN79ICHFG4TWcjS/iVO
t0MpDZU0K8QqVwVgwuf4Gvd0G76jD3ggmd+i9eGd11co38viw4Zv4qSMmW54musZ
U8ChRVuhQsc6TmQJghmiOJuCWsZytYoUbwZ9hxVwBuFDYj10kYhMCoziktwm7Emw
HcRoR5lL5b1s6qaD7QGJZNKjj/JKeLCUwpWJgKRc0Gr2t1DxrY9OrF07muvHrjAq
McQfnT0aLB88ZLOWcGHdrlzPtAnAlMKB9b3akcN1zF0vchpVArKxRwkOYXbVtfi3
M5FsJDzKDxdLiO+6B/Et914cZaDeWkwGnr/6gXQjOGoYHHQtuu9YM23t8NVOPZgT
p5xbrh8O/9KarIF5y5Pu5XBS9VmS9NhD7LT3EVVUjwPbHpB+Za1+uRYggQbkzaAd
hQGhaBSOmuhTd6Dr1GwQy1KWRhjGnl8dP76fE12bORK+Pt2E5+dchdnxPScCnRo1
OOhNBWaFvjbEO0a6ODfzSAmVz9BTW8nrXXqrd1PPLU2ygbJl9nio+O61b864OuzM
neHtKrg/Y8v3X5xNake2QnuuWKog+iNTl9mbVNIGnSSFLeEbw+CM5aSz7Abz/XU2
fMNZLbp7y0p/VyybpuZPIKLTXpPLfVST/0fhtZaRh6vtuB9w+zJVSb+i8j2fL0de
nh+yqZAyUp6rm5rRfzJ4P5tfm1OLS7r0ZWNmvW75i5ZIKrUsi66PPBheADxJfMWx
V2bB+0JcVN6EItjtTF6+4uOz0tUusqOEnY7+AS3QsP7Jr3pUhmTNaQE6pAoGxBiG
Bt9nVWRjQkZP5ConEeUv4N2Uk3J5gbH1YYGyHVd1yiZ2tG6yT2mK1lB0JAtfmwtP
kJ5p1ad92Q2a7tDf9wHLhAnr4QP7/bZGs3PhdYRqkT2qEON59XhFtekQZVZ6lwWR
NRvB8Gmm9qGqq83T1FHZAw2LY4cha8TeuTJEWOoXCRN049IZ9J66twTN9GISTPSP
If0pcQHlhTaQkHE2ueyrgDE/OZvxPI425rnAZ5g6hapbY3Dh/hwHIN0AA5u0Ubbc
/ulDC1UCXdrgucvnHTKZS10GiVmQ/Mg0aQbfLsTqf9edAoeLuTvSvFiykWcnP689
NS3iyMbar+pOwnc9ndCTy9x11LRH8GnOVvRUdS6mTc1Pkt8Y9lSKsmOWeWwNOKqc
eW8FvjifutD9rsemHDqxFlXXOyKxyuAvwykIJSnFApFPuK8Jw/6adUF6af58xFUt
BNoWk9cS6Fp+w+Z8iW1VLdNf53WlrANtFeOg09VttCggBTJdtx7POlh/84LTJx1S
u/llGbCk/cf1av7Mzi+mmEyliaKpmYtlDgoSQ1wcTAlnyNpxQK5lybfc/l67j/qR
UJ+aG67M+azjR8cFSjwKmcYpu0X4oFrg4crkGDDXOOYwvl+Tm99pscDa6qSk0uqd
5ShmHW5d1Cp2ya3GzxcqFD1YjSZfEcROVsOVjnRdLpOAFK+UJvmbYgJb4VZsKHEl
hklaFzYQ3Zdd6geMiZvvgjCGw1M1vYMyQ2kp1KiFu0s/ZVloQEFr0wQGAC6nNbTR
hGe2lNeTVyhCxUjlnYxzQCVERSW76gH79EBB8cBtgcEeVPoM5gQKOBVR06emsqlh
OnKTZ4XfqK9ZPgsbc5Qc7131tYDmmKKE8+xVzVWfkvXvk0svqCwCMjZkYd9NSSZY
H8zoePvpVAae8nIQ5CahJOt/C8PoFITkN5Po/DMFqdVMoMzk4nFdzdguiYkZHptz
VLiGKT4sGVDSyWgLQFlDnzJllBIobqLxZdbQ0dD9twHHvZ4BzfRdR+quXVRiF3xE
Wk9jzVLTc5HLx/eVIQnc2pTYIU3uvwCdIZX1dKKaGiSbG33e2waa/sFnuPlFj9Ak
dp3rhQFYX8s1JzseNni7XhH3iFFysyarg/qvT20IpulVu2ZemXuhfXmw6RYSOwEI
mmwp49Vl3O46WIbHiGgLuasbNg+cq7Jv0NN8Kzlt5IqYoOaRygHfjQRR13q6AiUS
tzcUtanSKzgGaNKSTfQvVzaBwUzScQNjzwOr600y6ZJrKYBigmf9oCeCDsjNvQC4
vBw/ovZ5xvt//6lstEDowVQ67buoUcYw2nk2JXn7sMSN5MK+VX7NQpJNnCv/nqf2
cblkoFcyR9v0nxWRJ4doAwt76b7zy4l1yCgGFYjECZ5qf1NE/cR8K+56UjWUkGaF
sGQFdgzgpw+T0KxKzva/q1s23GaDBcrAUaz1eUOpk/+vFYmo9QJecuUcy0uImtQ9
b+pDEM6EQEQuWmfbc22RFDRNZ9qoIxm6TkI19jxpyKxBcbK60VScVGxthxkNuLbw
BjB0W+pV+qLkJutyVsFBUTZFF57MpWonIt0E5VBedoOmD+dbjaM/jKxUmJAxNPLF
qAq+zTxQnjv+cyrfK2aPQGmc3f9BvB0VkoK7d7M78HnqSXsC2mwnZFbVK9hiTadz
TF/hINOStms2HSdyxkLziDNPGGedlNM1uulNXV9i0T0GZOrf6eheiXxINiCDAo9s
HlLwvr+V1aOserlOSVjRkytdRnS94iBcPCdb1OX0D3Yjje3qDB8Sg7dKUO9+Ncp+
0b2SDwPxtT6u21IUEDP+Wc+8RwEOPT84wQ4SuGBhsgSISzLCbBqgUb+7azN3qR5G
lyI50xi0y5Xw+rYfYgNJkCv3XdDMOWwiBa5NHuTVbN+8Ie8cXk8JN6Ob/EHH5m+3
YygKsasTWmwEceVtvDEBv8RAyLtXkjbESnVDqj9joK/qV2uenCvIULk3yyks8ZvD
vlIvBK4nhZNVIdTxnYfneu4oYahuKGZSoC1rn6D0byzqRKwXp5tI7CGSOCd0YEcW
Yn4S0my/Cy3RxtjrRaEyoNmFtG0FQbQWYoXMfENaHH7Qxk/fA04kEZmYwFzAsuxv
bUT+WCGqi3UYue8B/WLuIyytifkG9MpTFhiLBpUYsXL6EXJD656+aXDqsyQYH0Fa
tianEQpsVJ5NgKeJviimHwWR7Ws970EpHoKlsuEnQ34a1D6MtPvGnW9kEaQpz47v
dg6HDhvzKJATpkvbhMQyLAwKy3v0FK9CjNYwrxPqOHRqOA+U81y5HPv6MCFDvJxb
+tfR6JYcPyGRMLEK8HlyeZADZ8ylFxuPjUzBDI++rfAe902YEiADqfLvh/QlZQH4
5OecYmdDrOHlxvBO1QlKTzVnp2U6keMczv/mG/bMU5t3OKbdhKUdFIHySbNPzEVY
K353dZM1doNZDkE0iq2FoRLg4Twe4a6MvuQsloZR0rGmsY/sw55ZYX6RcIE8ZD5Z
ffkxuTZ29L5vS1X9csWLzMBKAV2bogTVClCs5uV9O3tet5iig1QNgGxZq0yhrQP5
1zZkArsnj+wPvntynZZO/jVsZEPnb5HX9XuqlY2S56eari2vrRKj+fKuJLORonm8
lIEhh3ztNfFBsWHfQ7JnWafwxqIHDJVCHC3Exli6Afw3VZKMgGP9PvpU9rd3hFMk
7TKVEccdMfCO1PQmgny9WlKFIkRwYy0U4x4RUN0YW23uzJ/+vY5yQrb3Y/O1u918
pxlVGGqkks3SNx4bEw7D8ERto6l/Hw4UQkhVJ4bNt32kOF19cqkcR0WePALlx+lC
qSLFjQ651DOowtXuG80UvFDbGUWkcEubz4GAKmv2XuvMstdzhxQjZXjqf292R56R
N0kXHOdshZd+qSoJJ9hHt9xXjCyzHfkimiENPPeh6xXEsWLBVcaZ4mm8irZKH4cg
WkHqL6MPyPP8SznsibiCzIIn0Wi1nqJ2coA2QdMHlGO/JKEn9K9FyQypxTr4TZ22
+GxZwU05DLINRatWT4L83+YjE/itFLpxJLZ2lVDjywbaBfuoZGpJXKU2f7GNOKnO
ViNiT3yrT0j+MSQVH73FeLTtcylUDHq52Zdxd/hkzXk01Cfzlr+/QEj4GoKXF8cF
ZwVedJ7AWDuj03Qj5vTZFDtCsq+VGAwgqE2vDqjcg/srN2b/xyqj3Dpg2YWJcKej
`protect end_protected