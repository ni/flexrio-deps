`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 45040 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
rC6KPz1bEhpOMfeLdNDaqEPQ1+wFTqU24/ZMLJMHvNoEuCBgpn/JaYYStWuWAeuN
CLoMQVy2OUhW7cT8eurvBtsSBECi0hP3y69X3KT9pNcKjD3+xjQpL9OW3b7zjK+M
9lPMofMeQu1DjxEzdNA5mhSCHWZMhHzA+k1qaynElrid1h5o5k9g79+D45KpgGgi
Mjcv9md1zkIcO61lCIr3Tqe1Q2IHjs+q51jzHqpGNeD+Olji4zv4CjhDY5X3UpSP
/+oHfE27gt16KjZGyfJyRQ9XhNpH1nK+RFmrn596tO8SkIKWK/5UGjoV5MugV3Sp
5ePSyjdb43E8IRTNeImtDMQedELaAGmLkxT7v7U6oOA29aIzFW6droO9s9Yg4BGL
fvjh7QqpZh31yqUQqub3OSWVeuT7aCIFLEQ4u4cnIrzJ7L89PSJrKq1ve8GrDo0/
PC3v/BGU4NUcVAwM5+vCZkWGQN7CMPUMv7omkVqyzp/Thl4MJlE8WXhFNyC32h9p
tiWyafXzHlf3oEEVVTcMpUO6swgEITFs8rwCNcqkWLLDi+gXEUnMHWpvxzmHnPie
k5zlwsGeqM2xHPX1Rawz6J7ixAjLUL25cFGJFtUDHELmwzdUL49SjNBGSV+qM8a5
qsGB38CcEC/AzV0lduYmvpitvOrILy7avukSm2yXhPAx1rN01+B2XOXKQJbw+zAu
0vI3XwPPMx+a0tnU71sU24uuTCOe8DDtUn94QRPDOThx9ibe8i5g5V0M/SLnGgc5
jSq1IkkyaZX8KUnIcPDxuit5jgMD+hH9Ey3FrQRne/1q/RzbtovuHk5xjv0F7r9y
4zy4NdQAt1+uqGRlBzi0Ia2eh3vhodzna94t4WaNFI10ZeinvS7uWKts6sQjv8o4
GQum9Y61eImev1J5N3OaMhneHQ0bepOgw3WuvNTeTsY7bGTR0XATcevlYlN6k3os
U9zbtJz2r5a5UkYFJGA/S2BQpF54J9D3d7XkgljcFoI+5HYa+NVR7k5FKlZicX8U
yTEOrJwEujIqFRNuGmOlFrLE5663NsqB+6wbQwZXItq8CZw3MNa0kIAjS4SaMTdf
byGFqm72VNVaXx4XjuA6FSvYyetVRnTQlHI0IG8rflVoRePhhgk7s356o2BlNods
MTGSf7baqnGviG8EgoZEBEpO4tlxX9vMD35u+V+A0J77GLc6Cl3aYyqnHNDBnp22
W582mWBTAw3zEjVxlyCfrGyJzbjuYLE59yyaQgo7VzrqgZMAgZnxFyX26wDPAxtR
mqnZ5O+yGgRnzKftva0w5MNaxKQFU5DKJiWPGPU+tRHJ6dyw3m/3qo1hAFTSrRDa
zPU2j4jXXzBROpB6cha2hMJFhT8nnJ+sv3dX1iB40rr0eq9Im5dkcPfYLafSVT+8
Kx6Vi6oYK4FBL6Tns9G/EFZrHhsNliHF1yaMMpsU6O3agsrCFxx7I+WP7QbHfKsI
1xKW5ceBmfxSYT+y1sHdaqwp/rXukTsMp5PBe8begxcRf4YIjKbQvMZ+P8tbxcc7
Y0bx9kuqGGQA6aTMbUdLgSy7EX3ul2FcpAJ/sbxwEUwE+wRCy3mbqCl1aLkg9/WV
ERx2svazK2m49bSA440h1hLHR05IuMjSEkY2yOURn8hhu2cv3oIdLU7ns9CcFz1H
+vuLhPEZa4uLq8Vd6FrHsPxuLZ0CXO8Z7PQkMb7ufTZPuti3QgS2pb+pjmvAfmeb
mNwvCHeiLplBNI/sD17oc35Pxm5+FbJ470l1Ft5agpujzJvVwewSVSwDMPmKLi9X
nhp7OTj/oMsiAjssazFUBRne748PuizD4d4EUfme9AJKnCsllhU4/hbLwwONe7ve
4qOpMpdS6JQeArMlAHYxd9JGBHDebkY6y/w9YLdajuybRk56lEmeBj9347e1f3Jh
QeFRNdG3YQ7FIwskSrP5yME1Ar3WHK1XK/SqjmXQPferPlAd4BEKeJKmQA+jEYKQ
vG3bri07zOA11+B5lZnrQ4EPTr4K2ApMLSsHK4zyu1bcMYCK3GG0TAeepml4rn4k
Pgbf1bUa2iJUbHS6+QjN/BC0yBB31ic48v0muYVsSloteLKnfdxqEQM7icj1LnPu
JBh+JHLisDe5QlsI1UIU9GyxO+HG5RedYwASyUCe9axqoavIyvhlF9LjH8IeMOmx
NVRxLfREs7A1fx1k+HnrdLeH/DE38SE2UJ0mUaKVWqztBwPGdy82WMYOvxEq2cdO
g7PUjczQcm6+czI0Ms4hIlcWEfNbT9JbAToEJpliao+zIgSD2cyt3AlTwQScj4lg
CAuiwWzO500rYFM72vYTSALcmCHA+gJMTLsNt2B6SAPGvcSRgQWgHnvL2o3m225b
KXOMh9dyAaZsSrFCtfNNxT2Ch+ulka4ow46/V3myeO/L+uzgxEm0YksWyZpyaYsF
qRVzJBU9qF4EalfwS0KeOmIEkSvKe6vnuC0vVaiUKI8LU0McWxkSsRCNibdooRlj
pme6qb8dp3cIaRHP5fNQAdzOgVKexn30ZWgN+qL1V0Xy6ieTMafWw9qPtAu4UfmD
L6L4UM6OC61bPAoGt3HrdVQAxopob5z8hgp87VgIQRre+VdVaak/TdHbPztUK/lN
5U1ac+xSrblM0RTDXHbykJAmkfskvm/mrJ+VN9FtwTY/NE/50ykKbMSkU1la4dSM
dhp9nhYrAwGLadd9ryW9zB5XvCevFqnzslUMq37EUe+TylRs2QuxXuuEYmh+x3VZ
rLjkhrBTkvWykYrH6WBQ9aqvDiPe97nAu6OwD8F0YWm6CRYgQsdcXd2IyJ0/BMbh
FUtq83InxO1qJWWGcXWqQnhsSwzRas9gQ8mQsf+QfQMIJzWIZf9ZwQrJzlW+UIHh
QqeQPYSBm++S958utW3K2Z7p82QLcCTIaC5ju9nhJrVZ3SEIheRuEK0U3iCtPr27
xctXoQ1PCfuek7ktBGPhcGCkZsUIhm06dd9/anoK9rkTgY4/nk7Pr8HuwEp5+6sh
M2GasA1D/ym7pYPD2Q140484RezA5gEMZpvmIljKZbpPjAVftl1sGnKotoHGIlYL
S86jJok9/rkSOsKRlG8xY0xY6TYOQr5AUCJp33zZrmK5jGXHZ7IVSQqwUs4crJlN
ZnuWpGwxEbPyqxOhuy2fhzTJGGnyC6irMuCc9DykjkITC60lJ5IXbNpbWC8sLMEm
mUn58Mhjuzg4F5fLSEMb7eKacqFF5e2kh2QaRVd4EE4Y+c6Z2SNngTgx0cET+Dsf
UKaPjWKGINbkeLoQi0DVE/WZfRjf5TGDb/mzkSReqbs2xZbq1LJjFrc6Hf0ziuyL
Atouh1NKaqudebfoiDol4GNsH9tUKJsRNUTBiHWzBEKA6C1i+Beh6LerYtQCHyuc
9rvxX03Xx6HiMBWySPR7U8jKm1UnR3lKJ7JZi6NMC7IP7aLRxILUdNPEHyBbkFGG
V3NCX08LeZpERWzmxAa4m16Demwd1feDXffqEZEtAztYra9mjRkGB7J6Wd3LWI8c
fizyphMqqgA8MTJ8RTUTKk/ymgYNMGUujbuvHmpGrIyTAaDEwZLA7OS65Hs3gvlU
L+HIHScCbu6Sf/itJRgRp/lcNF1KgW4O76K3lQ7Fn97EhB68mBwbD7pEtFl9Zlj7
K8Aea7Uo+iwYYd3iB2vHaqhelWVZTNiiyxlilDqrSLihJYWrqdES9pGMyI6BKnv5
69Bqdsl9HnZZZ91aSpWoMyU8uE2fyszH70108EfheeNNuCYlnnZoJ5swU7IJUcIR
uDpqLMH+omMold2rRfdQMtBG5neGbvrL2zcABgpLfhEN37SdvubVojoMTxxPMfJ/
oq3YF+UIV24eMvDq/d4T+ia1flpzE2nXaM0KU+Bo6wPYpgCb83tBucW7/RewKXlV
CbbTiSpTe1P8KcHoU5G6WMLTrr7pVdRRw0x1/vSXN8Gy9k5NXlX6Tndfh+BXIA7e
988lHHr1DpeisUx3lPbBJxJe2oZ2DmNWGBviinvsl7guqTZp0qp4Q7eX3BHCdQFK
0IOitl9nP4npBV2mBqiZy0X7LSkifXdho0jfshcdKlW4GC0ZYgGIicWI7V5kLnEB
vto2+6/64UnN02t3+4I0opXyoI/+unSTLaVwqamdhLGQKPt0CTZq+Qb1iGF7M08Q
bZkYkoXmb64TN54nZhEzoCMa9tfUVWCUXvQjkloYrNzdwCeJXSepMa2sK9XWjSSf
n2bGCEDqCPCZ4wGU9IWdMa/CfRUf4+rH5qVd9b1/eYjwX8eUnty9QbsGPUUeEO87
YU/eCUAW/ORic3vPA8E2COfCsr33+07iyDJtucEzx0FxOMpBSJs8lsEHz0+G4hXj
mkMpUn6RSzqE87YVTc4hoBPm38vw9E1qdhMsqj9Zsol9zU0jn5WEkundsc+e4lXQ
67SVb59+gbHgtYtS/P8AFINXlBK11Qg+kmKRxBlfcE7Yk6kNXwnwK/PNz/oxj+VR
UMpw2V++RjV0aIsA1GliuA3w/ayzC0YFxU2+RmdiHtlMCcto4aMZtbljCWJ4uDhH
jiLuhBIAxs+V3KAylgpHXY1Y0x8xEJXkbV55Ao+LYIBqF3kPu8x1tIUguDlzabKV
HJS33evwnuXGszxjgQK2bY3jdF4FXbVVmIm92cf5Fc5Rm6i3uatN/gwwahiPEo5E
pwaNPLtxffbYMGqjuOAi7pPuYSvCXZHIwPvIxMl+3WgS1v2bzznbUbiL1NPLg27F
6A/ATX7r58+PlBFyZF7Fn9ahQKDhacPKu95wl/qHMlgEq0rs+a0oA/zCAe10VLHB
WyegySz6wTXmPrXBA6cHGJFSsFJBBkBn3Oeo9aTRrTzAFPhhwj/xsg2j3bc6WdAs
r4QzF/HZpHqbixSONFFKalofsJm39ZSgGCK0V3IhOcQmtzSikj7MIhEGujkizVAf
eDz/iS8qW42ansAtF+Tpzui6PKuez1NvovxRvmXqmPl+fgIJow+ULoMtykY7ODUx
tpZHfmvwZvLHXtjg/KhiZEkLhY0hW1zfj8cBELkPxyBUF5/SerUBn95QPOdwmvs+
Pq8Y5gun/OKMlQTPHhEsuy2pcsgPBxq47NRFy0TJ7OqHm8xMSaWD4zQhj8yqS+oq
3pDBO2xkPYD+XNDNEdOoatt+4nuUh4slCGjEDmxe/L6NajczuCnLElMapD/rW6gF
rIn2O1w/GZM8iivxWxp61yr2JzZO4nc8w4IC5eeYyNpxmyerXSjoGLsP8X4bERTu
he7qY8/Kuk0Bl1uTNNLQgDq4N3nny93j4KBDoTQQ2l2oo8AsX8BOrkO0icXDnEZE
98JMYHM8Td7fuOqrJadD9AZD8te4EVI8jO4BfqZbxxWyA2h0QGqqvf1A/NnnTg0h
UaeIVtp0EGhHNNa/U+hWbj6r1C57ZivAmagVKjOIDsE1vZZXPvwlQzM5ZEyVHu0F
UapHeVPoiMzaS0vUdb+vLW9KuE4ke7yMyQQlnsw3dW2Nyy16acAb1tvmYtD9gYs4
/7Rn6SUd3Ucpslra6iaODq32dQ1ogliTgdncZoBLUnywo0BnrwXd32LSAdHdVPQD
L/1eT9rNR7LEE3OxnDeF9M2WYoI3tAM6Pr79CGR0SyiUe4ufMSB2C1r0ZoyEF+z3
NASWLsxOtqf+yUkKZ39gV8lDrD/6rUPet7b8hAXfEx5zEoA6hI5xZXejCz4ByJTv
PooeLunizRqeq6I8Z14kWklWeh6+tLQrJEN4dJjPtEFy9XbTL0us3r3WyxRD/E2C
gezpCM2Q9M+iFXhgtD5VmtyyEcTcPJvRVdpD8xqt9aGWZYFghjJyWku18fGMDwFP
lwStZlfvLr3byEz4icf++L9cAEuDDdONo+p5vJ1CC+qoKHpHYaA4u4MKobtuxVA4
c31yOWhhpJ1pPbVsriCSEmnIPXn0fl25C+TAcYDly5UgWVgzzipVn+qrH2OSmxLL
4Q92Fe4xktsWFNMZohgZwj3YIvvucPrmf1GCdEa2fduMPnD8vo4vwg9z3r7zqGQ6
z2O8wPmbvfiBigVv1CQSQuhp3zw28hOVeuimtn5IHP3rx8qHjGUnRfwb9mUCnEtX
k1+iGjB9JniI8O6DKQ3oRg3gALY4FeDvaO8XOc19ehUROVZA1QisYsKfwK+8GTHF
XItKnxpbDaEQ49UpY39QQAObErRes1NRKVbxja3VTx9bjbUqUwBTwqglsgDdUKuD
CCIDeiQYK5+AQOzgiawnsnnRI22rm4Pewd+uuzYUkd2+ylMlvbEtmAptoZl0RBNF
lhdnStcLKLH5j2QknbdU1/PjE8U/5GFKDhaJ5lIKLBl9Nv2yS7I1ypLzg4kab3NJ
48N8lMlfKnuocPo5sBOv7ok/Jm+lnMR8eHE2CeyBziAj1J865TMpyYpXPf8aS5Dn
TCGB2jBXCPDEtHax2yb+qenczZ3ZYbnnTu+LGqHSbbmhFBIHY6ciTBmQV0XGkIZU
icdRIxGHFJtdHpqxXaRZ4v4AlCwr9xBY40KBGEqT/4eAijYRqbhQ9kqtj7vg3MoW
2Vb2qUECiWmnhSkI3lZX9P5mGn0m4r5kcgtebpggqiPM/J7gCIMiJsd/w5hHQhM0
6ssj3LBWuX1VMyMiX3a6aX/mQI6Z0mFt/sF7Jf/JO0GkUR2TKbBKTqxFwPs+hkk2
Zrm28Fl1EamJuo6h9znFgC226KUFNQ1FdR1BoSmLFseepXnn+ktMIgD1NFnuiOOC
f1dcwxyhHm+ZXkDLhvWg2KUkCysIItO7548W+O7tdMVHrMv3YLph7qjNl/C5BUQI
NJU28JW+ZdmXeQfEFmXLhAKlyNM4JEJtFH7uupbnRjlQK6zjmAayhZhPJ14CVq5X
7tFzxIPTCmS9vAKzyvF/e+/CYzilyWLypsQodlOT9ABwFzZTBaFi23yTXEIMIgsW
tDeQsmcufb8taRQ8CpJlV14yMFnsMOmzkk8vmIHPdogWTU7iKQR+mWnaJb9jBuPR
4l4sHaVp2hMYAJFqokyHbLtPPqOnNV/pHTNW5vChxRxTR/x/3b+vaNCBOLhx7w+m
FSz3N1G/mOozRK4SqOwFGENLHNSVwLhgXUA7E/K8y8b1w+HCu2Q/4xqyXprG3uFj
d/R5llifw6m39FX+8LaODMLqX8F5xw3rOHoFQJE+eAI16uzjE8DIbrOLfm4V4J/q
a9MDYWV5MPrGc8rqchWVULZ2h83Xt78wZ4BfdPTlVkHhVWsiNM1svN843kvYI4mE
R1pCEB98OMvUloI0znjxyAYIz4u0HpFtz0Iqz0FD9VVQtQ11Ja/4OEKLLO97ydri
gzzPH9vUR+OQ9QaSotbN7iFgaHsHIePq+0nlb01t2fYGFbCm8JojAGC6yPIk6gMM
Jy0JGMQ8cxrZb+FAEi40GiuEiNO8duO3U6nBoODZR/0CHDR5m3gd2tjkHeCUfREu
UM5zHV7M02yFPSOeEg+npIBzriFjLT0/6nX3gyjHsoKhIkk16QFWGNaxvATym5mQ
KlfDYxI7i8HX4oUFLkRzWbjUGGbamDqAKp8mbeT563kiQSJM3AcQUMEumwEUn38/
ug/9sXj04i7ftG4+zAkXYTP4sDpNw8LY2C4Guoq/sMIO6rqZlmP8D83hNs/KO6yy
3N2K8VQebJnmn/5sHdY9aTa+QvEg4vygDR2ous7wxyu7qKtzybITf9/Ak1L7k8db
278NDUK35ePcVw0jmy8cD9813VNtGm5V3LxUk2s/dRSl03dSlvOgFDg0oLE/1SMv
Tt7IzanCTAAsBCDdyDt9EGUptGmmbUJYQ+1YfoXG39PJQEL79Qxz4/kMrPPt/PzZ
z2R6VQC67iaB4n2RjBZcA9LUyQzVMiT9C90RkNj37LObQC+cjmnbQm227+PjkNlH
oN9+PnGivwTAo3sNHLbR3br1S2K/0s3lFzxMXgTN0NaQ4XD9AdGXnw9dTNVFIhRa
UphHJZOYv1yAJwIfKkMHIfN+mJUzUMI5x1uiAKnvNBSCVpCDYneZuLhEkQh3XN75
YyiuKe3S8kFCULWFHPkp5JzbKOfk91IYp6QKRIPYtbNu35Qkk+q6SIpF7rXHnYJ+
df5QJDPn+NoQsj+rMWNf6/ScxzF+B/Oz9SzowvGh1u/vQlyXBD5SW6y3vfdDsysp
3Tl3i+OAUJsoDEY9+ThsJG9RQ1cGPiXkujh4DTbqhOYZT3Xj9qIAUZKms2HKMN1i
V8VE9h/FLnWcypEobbc8t0+mLSKHyA11YGrkA/PLrihMWqyzIWT/tqaJ32De/fY7
0nIDxA6GeePr6N61jJueOz3UjtyTyBJq80Drl2SMefCmpN5aLg0mu2Vt+qPL1o6X
F8Ueb2MLV6pbjwC6USVi0mtAotIkgrcG++A8bzifoVUYI6SwI6FXef1GQ2ClcDJ2
k8yqnkd12A1wr3RFkbPG/OanYjD7kWsjjWwTw/0Uw8pVL+xhH8dSrycj+vksl4iH
O+PksrvXzZZc+/AL5KFI+p7l4vflkIgapHWjzXCdUH6dK+rWWE9ebIlo/b9Kd2yE
xaSvNLQ/A3skaukncSGOS+F68NbRZzmDmmxlNkuKeUKEu6mORP25v4yb1i8RJoWh
CA+Hgn3zyFyTljJaZjEnfUZoh1coBHxqrq5cOgDfwzIa9M6nyY37gSzaobvJTnYh
zyw2UzRvDpf0ZazPt3Keix3rfPLRwqv4TqVwEwMxfuPJRrve9BVNgkEJTz3tJOev
eoxQuyPgibn1xbAFAJIV2CkPLRE9AuEP1GJvSSpXqVp2y3jJJmi+IEGasSLF4t4H
fckATNNYQaQIsLuFsYnRzyIjzSg6aNDtQq/9wJiOcxScPHG1XRGBU2y+lolBj+Cn
WxqApWlZZQidxxlW3O7b5CI+iGyuyiZDBx9wZiypOWFQFzVJiiE0v3ChyeisO36p
nDo4wqLxoC/vV+TXsV1IIN4ufWqUf3dbMJ9inlM5r1ylh8f2qvSP5Ylhr+bNFvVr
SiFybcQ641RzkdZph20MZ61zjdXigJCXpBJ/T5n2Ck+3VHltPBIrGhne2zSrf67e
w+TzqZhIqjHTZ4zIFMAvZzMV/ou9/b4T10Ksdn6H97utrTDQIyJOKnjTjh9g0s4m
v5UesBKLYNFpjoIOt45Q5kpLaXhditYLpmq4hEKGwc+2F0BbNIc+Gkd5rlFasyCQ
kid82yJlqMoNCRrEz3zKEnbORlGa7rgYtrwORDj9phxH3eHrtuBGvTcSI/ocmOac
1G85bpH858OiotCODvo7CFRx1uOSpcPF5enejU1ezWPTF3QXRJMQsaTesATQjcR5
n4ia3cp56ALCnkG5Hj88vOGix+4AkT3+9LylsgL8WQGVAEH+Pz1sbh7kwUwu46BY
nsDNpl0MZe76D8ehta57MrvFtZ9KWsFseYz5xnHQMIDwD2AsgTCsQNLIztWrGy1R
mklTDGpWLq8a5Azreoa956+Sz48XgvZVl3eqCH8nu485qFZD+/AhkC5YdK7N6EAK
HEQuq/c7btj5CYXvqBq6fAyg5hJvoekEUXOs50oscjHlsVv7WZf9Sqg7cNEUkvYb
hE77qpKY+0jkTFym1fvB2PxeO8O30BJClAKDozRv+RRhH81GW7eJcXIT57e4z24N
e0YiFSiL9Pce2pb2TP2b75nRqwe2nWV7kTO1AS/Fyy/GAuxITHhQfQYYquIilbSe
zVZqJTsWPt0KEh6PqS15Pv4X/BDlv9PSksVGqIxvt2uZDw7gTrMoHCQeVVHM96fu
Rb1w9steiIGJic6V46EEa+TFG7C/t1oGwfshJl9z/00Z89UrDRTQ+VJHpcDTLyRG
v1ghiRCpHeU3syWPiutfiKMBJ4wYqomfgUuuanBeR9ltG3iu+d68c2miuOEYgIVQ
UfNcUraz3Oc34SknH3uyWGC2WPZ/QJvYYyloGo89m5R2ZJpb2czIZRyYucTuX6hL
sWjgMgKgpaqHMfR7qp9FuIqUOQVDZcaN1o21RfTyo0YtymH1QQIXSlAHUO/tRE54
8y3/zEQwBtFticLMGUbTlDBZ5m6y36HzFShkuYAqpsDMaPJNC2mhU44BGfABkxAw
VT9WrUYpBFFOk7q7tj0MIPfHpIqJohOhQdnXKeLXlWOocT/oRtlDFUZ5Pb6BOSmA
8g0HvJ2i+d/7XkJNoIDV7mzCfpM4/6fdvGl9C8miEh0mdIncpIBxVHN0QZbYlKOn
1Dsi/Wo6e/qJfyEGAm/4wyADW/6RzXrIdUKk+tzRULAHzrv/6LQQ0mhmAcQFHEXb
tdtaMgEAvqcrsQlO/4S2UfB39wcSooC15e7JI/M83glgPlRPGY7B4ra+p5UAKi/C
8kQ3DKyaa8KS7fXGq768dK+ehEqT2TKRSA2fxR3iRrRJHfAwMKnQgl+ASHhbXFVI
1cuQtYQHmHfUKHQ1Zq/T0FEtTH42oJ2jGWk+DX/BCLCwqmx/e7qbAuMZ7+F+x4wv
emKhHYyH6ccJr67C2xOmVwN+hViYzFuChZpYvkuiVPFmn5ZjxSFtxE8ZeIc1Kuae
Zk0m0xo3LFNHbGv3kIcaRCMEyJtPF6+FzGvACS4vkE5sBxk4YScUtwIR1NcABz0C
mn3JMTE+x7I4yZF7Xa3z3oi1OVUtll63xK347lPjbRwzY5VOtCbDJ88cxhiXxPON
5IKs/VUtsVeCuNBymaYqqsFIjndY0hnMnmFTERo4a7uT/9IMA3awZQvVJXKoF4Gh
wl8YPM2fgUHzIIKaNeQFE1XpEooPJAMLf92YvUQvhTpF9qMWiBIxcIqgcktqBpP3
CKjZHNyMQOQ0LVL7MfnUszsKbhxQVrieOJe0ee8B1iCkoVT4XdCbxVY9E3RzkIv8
UA7mhjhyyZ7hRdXtVKOJtj/3HE+OhPvLA7SvXmK9THpm119YkKLWg/6euzIfU8OF
VYT1Wl7RzIZiiG9NdTTJsX8d1vb/ZWfNDcT3SZUnBnb2mXEEXvtriWsoqZffy8wo
QJKgmVCS1CDX0nu5DTq7j2+DvwtSYwugun6XjODmo6uLsfCAefnUNKbM84cqonR0
qWv6lp2RJFMWXgp++yCa1T+MMYxY0Evj6YUwmQYOE/ipH0o2y9yKhgYVC/7s10mX
fMlS3/pscXzjOkuhd64jN5bMqoaYBWLKrnN9ma4AZd3Q0cJ6xGCZcr69Ux+uDxCZ
nlLbNFWmhENSjb9RcJqZcDjjouxCwgM9EQ3ltoP7l7BUoWXvEd3Pxvqkmls1j7hB
WRk+wOhyFqunGvntpVdqXAcTeCm9oTpSgghy9MWbreFjOtABtraGjK7+kuRjRRfZ
rorrs3TZW1XCFQy8KpBbaeqq6RbxyvGNHn7ikQY556n7h1THkJ/ejdgFaX/9CcOi
Y3R0dvLyypBxioRfhXq0WjOiQxDByAhzi/aviqLx+n+iH4nfM2t8lDhSrubn9Wv7
LZreanaU63HzkEApB5AjfGwFgDYYkM5a/0yx35p5ZPE7CCzNB4pIE7upmv5niVoH
OkJ11lYXOIqOJB01nFL0fMfKxdE6GNCkRnw51DLDNFxkFdW47UNJ09ZkQt2y1pyx
+YcIJdqUOqjcl041oID/MU/1tWi7glN6z7HnYdzWMcs+bqWAp2cBKYCcm6dDQ3gk
nZYoiTDxjKIItjiR4FN9ZqycscEOz4IHvdPrgjYJkfng1CtEBchHZtW1MPhoepg6
GFiEvVUnkJjLS7gunpJK6Zz77dU7lPOlWruarrW/PKo5CpNCl8T2WNruV81uxU1i
h9UqzKgSxkruIKjcVvUA14rJlu9fYjkJuJPeNB7AgVYw7HkalV5pYgMS9bOm8jXA
gRdbL7Ly76WyW2rgGZU4u9gow8nlkrgrLntIao32lslt3O3q0zMqvmB6y/gBW6TM
9sOelbGEUQ2vD7SyzrgMsdqJ9n8HsV1PmduA3UygKqwVeeO/D8TaczmK0SYz6MNW
utEuoMIks3hAF+Hr6bGeR8DfW2dxGBuV9NW/c8ira0iY45wVNS3mWSaOVaZg4tV7
m/CNaNrlRZAZJlG6Mq7cTi5BpI0XCTqIL6RpLiuZGaQoHiPo1WtuA4c8WJcSWut+
rk0kx9QQHdyVlY0QYHHQBK3KQPXcypjVLXxL6HuV7WQEwsHFuYKe+ZdvVmu2Rvrj
+em+tS4nz6IVyv8G8weJmL7VqzjopLGgb12xYbLLWMoxQqljZqrQ6HcrJxXiszkw
7AUBrxnCQGZD/nNtHs9lyoB52Ll2uwiHBZ5HQWkUIPnBCR5hT9yyLmnpDWgeT9Ba
uPN+LbIV+ZfjQd2Mx+KLU/2V21nLzKH7q5lDM/ooQNv6Gp4T8r81IhyiMYWG+EpH
IL3HLMpx2fXyN+y41k7cQY12TBqLJAJj59hxHwb/rFZv801OFI8HqDN1qjWNlB3E
SDr/RZVt1vmuGs3bqkMm2AijoQym/bwQQD7uCtEY72+L/hl4TV00PHowHPOP2/QL
UgWrTR4oKfnkr+7/ru+pyVB3Xxac+z84kMOOROIhWL3fqX5vK9hQV4L2upjKYpLZ
YgG1JceWSPsYGJXZIg+g9v8uE9gTxbrbTU0TQzFN3+j0RtJCKBSI6AHUWoD8i1c3
SePGbGMtNO5PKzJdl4ozkY81etMrze9CmgDbukFbWS2HKqbo1PReLQJqk4qxariA
hpIrX6h67eH8kcNAOGwZyEYxJmkB0QMDHSi55TpTyc0QESSC7deI+BsZ9ilu/e6J
/wgpGEF0a2sUAw75y9dkvLESOUHILxE5RnuYOrji/9uje/dFBt+zGFsq5JM/ALys
ACRfRaZ7KmzS/OkMz4GqsaOiA1DRDV/lIKgXzxPThV91vuOUDv2lu/pNYUrfbicC
I8wGnj/Rer9SSDp3pdIr/1eZGJgitqrzTL7aakmISOkcKWv7pxaviHEbZpufxtJ7
l0guPaxD69EQpfiF/Ab790FI0APMjve0ahkVrfLcrpOtpQV6pWAhooy5zv9vVYfP
JAl0RG8P+WHhr8dNBkgzx9dqmMOdX8YxsEcoX9ytpT5acSGNLUU9HiCUU0eztsyK
XliXU3Vn8xe+l2W731/5z+s7Hhg3JGJ17T8/AVFJvObYAkgfvlyd7Z2N+QY7O8If
69S6d6VIi2pOnHHT7XKve15a2VF4gy6NJN87I6oWrZkLF79zpySTi1hdY/FJaKt8
/r3euUrixTXx98vWYfnJuvYBXTjjBI+0mSHZtJ+COUOL3VmUlgRHFMMMjsvJsR34
bYjY70j0b3J8qZXHBNUYsBj3N0EwKsN0Bd/28BDyGFZR5sjkcf88+daL6/85iwE+
BFILqeDtRjH+NjYkfXwy3ElROU8FTbOI/BO9n20cO6OnF9igFIwP9CgjXObqySbO
Vaowp9zjEWaYEDYxCe9TqEzEiFhvKEjssT+elsxcx/IAVelgpn1hS36yJHNDLiiA
sqqforVXDsFIAE/cFYwx4Aood0Oj+1ePI+61eqQmLvd7vrdKGwRbcj6CR1t/qhTT
Ss4Ceh2mDXZgXlvvQM/i4QokEOqwzbSBLrj9BS4/F5oIp1oEcKg2OUi1P4nmarBE
K+KTWeXNLBwhv56xSSq7wGe9Q5lDCITjmajLZPUsYmM+589xiVzmTNXkhe+pPTNC
yL2FPXYViGk8bouCNe3pTx5ShwkYAo43QRSGamR0Ih1vET/ozQqriKG6vNXZXUMR
6cIe9Yn026/Dhw91N45tgnhtSVX3NWbWjMzm2U1+4GUbCPiBIxu1b/HSyoja8X64
WizXa8cb3rWhw66T6GTPycQCRS35hJxDQGcT6aCuzjWDlASj1Xmmd74xeTd1kDPl
HR2Tj6jDX0DXwkBEMnXe6X+9jT286yeqUHP0977BWRnI38hw/bOS8opXPwcKIE4w
UEp1xRGjuc8lXn/0GfMHcutD14eAatbhtaRpkYIQ+6b6hVk4Il6Uewq5Rrl1NbWe
FQzffBUeh8rmwg5s9uUhJKYIviGhYwcjojKlPZVcG7A5aBo3+XPqqpiaXqN/y99z
OZ699rlA0W4FiSK9s4ExH6Wxj+P0mhB4j/xbPfQkZpt9CwYmxqigX+GMUjB/p34W
RWWTheLVPL+MBnJuR6V8Mvv/5nhMby6k9YkgvXxCKNW/g9WNnwPkLQM9tlXc/hEq
3WW8RN0HjLyf13wrVRijBauK9qpS3fsYizEdqsnzK5DvoS3hHIkHCiBzvq5WXGRS
autM2V9HCjkKrGt4LzOK6Ig546pCoWAtGooOgJP6r28LtDTJhwdHDCv1TTVaIAkE
UVOxoLRaknHCZZ127U4sfy1IxQWZfNPsScEzxFPuOGb3rCTHphsPT5+1STgGQ+yI
iS6k8nCOtwgT+aZQtk2aodA5htKBrf7G3uSrSg9f/Mi9foxCYnD/8xRHANcCH4zU
LSw+BfeWEzxI06YqsjOlX82mZQ/nv11+xoyn4UlmN2U4+JaMhNgUAj3UkJ5m5INA
l4jviNQtmJGEikDmMddbYpDrF8JVrmiCQ2Rk35+AlZTQDrFlt/E3FCRWpPkbcND2
Tw7yNieDipyBbtoSs8TbIB/DadXT8Hq2B0C55vgEjOIO9zIGqLhEgKvxEglH3u3v
5KQN7EVr5zNCHgSWJvjTRj7pK9NlZQOmc2oorMr49jrqIMchll6INGhxGy5usRcz
5OVJ/Ws5uNnLPrewrcrcIMIqdcGdnk5OQ4FUJh9qOCsnVpRlBYvtfOIOCPTSPtGN
/P+eqtcL4uxA3y5Edu9IUCaV6LvsVKnz9l8zFbSKZ6yfSxbZzQ32GwCCGzq00mRg
gqjV0nMgfvq5VGtjlUzKv2Zw+QqIuIU5OXGVS8ESxcJg8ahzTvgc3bHGWgAJZ2MO
AZVrE3XTKzQPwfxMm7ZeMpICyVv01iYFOf7+ANUPwgrQXtss9FqZe/dx3mfQ2cO5
LPhAlWOjCvREXby4SsGsxvP47d5Pl0sO5imQMiJR19/5esMg9gAeuViOx7sb+dw4
p8V/0H4fdaS5lKCszHCiqQ8jilrWHxIc0dbaZqJOB1J4GsHyUZH+XgMeN65R5BE8
hLpY8z27GssiasnqSzHu2oLDMVsuOo8yPgwFJR6s6sFv4Cz3LyR61DTqrBiMo3td
lWdKDFV6TaA1FqNArf00VZTqw+GhuOQX5T7uQyZkX2pf2pVU3Id+M5x4UdJR81Ew
ypeIhq91Cz8A/QX0euPmn8/Xl00oxnAfyrV4i3drAh4sghm6+tYvRYU0tsgy5/hm
BSX8z0jvFDo8gnWT+nQSGwZX830RUP2jFKDoujEfKc7hGX1FRraH/OKel1zHbCK5
kmiCKue9111MnMOf0D38zViK10XIBq9/QcZmHkrfOuqSgG7aERjEs7HJAINAZbmh
PpA4FLxHlDItpXnJ98vXjq4VgbnfPvm3d0RYNxc3Cf2ST1ZGICtVl2fSebkED4lR
tLyVtRviHmMOPmt6hRkKhepSPumz6yHtgU4VZdR8nymOkTGX8bVvyT2H92zOzktH
0I8q5Gdksw3rtzpm2QtQVFX5N3eQRkgsWGTg1QOgJBgl8agk6I+udMhgVyHaWmCf
qbSMtlEoy+yc1k39h7DNKVozAYwGvvsFyOq7enpsV2yfDBuvy5DMCMypcVXYN/iS
KoohnAPFV+Oc6i7f1KGVrOibEz5NWJ3Ju44iNhYtHOsnh4grJ+bts+t2r6AAPang
hx2QEShIW6Qjlc5kk/wzvFRFcIl38hKatq3gT5dc+bFUNjj6yuWO5uWVM8/M7DzA
HP80cFph+lvubp36RNpm3w3tHK9aqsxUo9Tpq5n8i5UjDVyHMW5dEQHubG7Pno8i
qD/E10FuWkNqYL3iGNqcQJ8Ni5iIl4c+PFydC7QWKhAjvDWyyA++odV5Edl8khDE
aDFckVdvsZMryJc11VsX2LLCycM5YR5I25CjDUxzbbbczV0/CEHr8blLBNFYjfPi
MylhjmgT36VHbiCI8A1+cpeZd4dMuFczsAIt9bF8TYxYQ0Iz+CrqI6IDk1rYrhm/
i/prIfsnR5hxQT8UR5m1HTllRgPp9e8SclU5Ny4kiil7b1avsqlkEU8Xyo6DYCU8
k6IWJnjTe701ETPAjq2vAodAZfQlzV7Fml5SHP1gKmjRcxTXSR4iCMe6lleRAMH7
aYWSyzCRg8hLIQxk/fugzH3XlOPCjAE2wFOQGolweeMMEMUNIhWdu4V6lPtE84Cf
O+hot+HRcnns/8Yr3qJIyl1WHA8ZaNGstgy/jGdDB/tfxcBITBnu/vzn5Z28kF4G
ZNb2emeCpkHeUpaaIvbjOzcKpxQ59GULg6ZqjaOMuG3A3pceQHg8iOfKlO5hfG+g
fIaMqdtiMn/P8gSbkixj+YS7YICO2lyW8Jl3M52sF3NQfQe2Zh7j9brIX9oAwLTO
V/cqGj+9Fb6C2NXfI3qi2X4dHDABFl9WEEB1Scf4aMhoAqmQh1mGiwvSfzJFIoHb
h2vV9uLiisK+OxHuFV5KwBIPNrUjvaLT0XNERqnd9OGlv8SFmIHf6k8q95HLerYE
0jCxVsp4NhZ2SdQizcyP681OtVw/REBqPIihETDAe5K0EDZ826Gpw34XhvFF5HRp
xF9Hzj7HGUIKSHFFQ8QSevWFyxRk7FgTAG5YpJ9jgrVL06bQa00mwru9PrxpM751
N8H+1fUPoDHc1xoj6eODAtCHKpIqvIWZSTLIaIZBhlDQX4AP+NAJAU/P2QidqU/5
0wPyQblliLAAxrJBOG6S0VWrXnN/mrtHP9y9hwySzwtQLPYu8jhWgfMo/g4AwSJK
YId1j20HdrMNEY3MYmYr6wB+zZVKM12f7L9KpCIyqjTQNAXmtuTdawg6s3c1gXUT
gkF2U7SwxT0ozycPHCUIgcIH2PXsolMZl/VeCNO9S5zjyK8OHusFVSZNtP25Zmk5
lWr3b8CjY2gTB/9x+mGH7kt3qnZ9sHdqTxxObKxmxOQ+TjC+pvdpCpbGZ2jYTamj
pAM6sF4pWbJYlTgfLfYYd6ZtH74ShRgjaWCw2zWKq6AOZrIjnGmwsyVsUqlrDbdZ
U+Sl84vc6bFQrCcpTpxK/G2+Cs+ZEeO4bRANA9FckaR05pHsv7aKUuvT5jAbqQoJ
zBryDRynVRbUIHsBnVkL4mU+6hcUQbkecQlT9VLTjC17WuHAtCO944xzUgumNryp
whYSFJA5M9Z9CvnyXLZago+kEEYuehdCrrLbj/qNkW91f7j18ILc67YBwHm5qElg
hTVO3HB9/SPkXsDtDUVOAtt3SJzsZfzZm2qgyowBsS8Y4o0qlCfWL6jNdT27yO15
uieKdozg+D6zA3fHwGzZjxoPI6A4UUoIGkUeb4wocYZitydcRMTZ4Sxz9YIlWHiP
YGDET1yOo6d4FMPe3Mp/G2AuJIZfDGwmmMUctEtrtg71LRotXXW/R0svoV0oDNc/
TV37jZQ8vHTqSxf7xWIG9mPn2HCCHt5fa7suCEDzEnHdwh8gRX5iV+ImhrHTsUW+
EsWVv2r2gcOu42Du+fyGAusFeJYPlcoCnLHfs3l5v/UPz6Bi4L17uWuTjLkDFV3Q
i9y7zHW1RSbvj37QXp1ST21R2sig9tCRAwKe/a6kx0J67UfAxFySonU8iJ0CUIiv
IfbN7lfCq2GZnzQuG6jvTHL6etogpYDIjxzEy63IXRYOJX1onSpTVkXBiqYP2jRI
Gm8Jr9sVhmK1lnUEHLiTAtijSfxU4EcpoxB2ARYwuI59tH/UazwOtAp5EOjk0leJ
icIB3vmMGn6DJwocsR1n/JE8RgAfM5aSipQTVA/T99g294gUY8uEumjHegwbutzW
QyLtSQVNVv0HDw2bUbK1BwehXVy/SOI29C++jcuRHT3KKXnWcFEJvhy8p/ee4nFd
t+49NVfSEJC1zg6f5kFtrGvSn+F2H9JgmJrZUzQNr6Q7yFKSkxcFviIRbiuSxKeL
LHKukuRL7C3GRrlEY3VN2LCoHOAymSJEzI04VQG/NllwQE5pkF2EpqgjVk2yBshq
ob7D6aBwOYmpNF3r5gzUP/uezpbExzT3yrmw8XF/njqrnWLq9kKdmOI71Gqay/pd
wg4ZUjcipr2Fdm8B6+ogLIgYCDRhl0w4hKC2IPMGwgIFkvZ+DdCN9F2p97+9ugQK
zc26aL4YWuXSxw7tJsaBPP604GFhEVmdMEcW27SXY/QPiJaGSdydKhxCd93HlsMR
IR3fg+rURQ7msO0zTcaOQ0tEXZ21RdY46685rdz+QMCyDLDj9TRAbiIviJoE55XX
CNq3PMDd7u+hCdXTQ+YcHMLqYEecA9g2Fcy/BuXajjcs0X61XPwE76ANC7nInd6H
AcwX1sjKy6hCj6Yh1Jj6O7bJzpK3KPp+hMiDS42DsBS+5E3jMoT7ARSoThTkjxe3
ZdRJbiP4sVVYrCJ9uSFhIYxN34w3tHOsna+Ic980vXYHWEZSrE6wu4XUsbPXDrHo
7zFVe6IqBDhnLjnu/nvH0EJMqOik4brgdxBY7rK8tR4wV0vFQT1Tjas3CuuxOClZ
FK1NZvr0dZ6phPyO+z4xJ34gX9cA42u0AmXwVsRxKSVlGkWS5HIa+QLsV7U7KLFk
exMflZGXuxIjJZhbH/3YfGhGGIe6+IUSWvvk41fpUsIrHQ59cTqiIZO1huGfwfhs
nJwxeMwoKvrfZimjKgU0Xlj2RbiHyGwOHB/hQ8dTx2/kq3SK2aALSwDekTEuH3eX
FPsIyMiw0+RDOQH24Zd+nlwU+fqgMjPgpV9uFZdDaileex8zv6k65CZQRRnuzrO/
d9c3RxRg/W4SZwzQ7g0+n1ywgVzwRUhfprKjn+N6Dx+eN5CvC4yiByhO3d0t441q
08NyLkaCz1JdHUl554FUQLCwuVeOhKw6lTpEbBYKjjym+NXBfFaNsybm3sPhMIwM
Ens9OyTws6ChiFr4fTU0UugfdPr7sV+apbiDJwNqPzIuksxJiU/udiUe23Ada0HA
Dwx1/DIANwyPbyvnMD/Qgo0I8CG5pDxwA6tWS/P6RBhy3Q1Zm/t06iNJ6fGMhkPC
fKa2QH6u/ICygSATc1ED8X+6nud+2vmiaCWm4rIVGNJP3lhQgPMj6xlK2/1h99tA
TrTfmJ87LUrBk791uLrxhzBoEudriBOeWwZtW4Qs78qw0gM2iwZY0XPyt6f40pai
EQtTQfHPA6zbrcTLErI9dkrBsCP9CdtuDVBajz1kxLU687BzkpaO0SgPTWZ1y8qd
wYHdBQ5BrvL22WwCs/uuohggZRJ0eKIvm8pYvZLR0PLRSOEPUyl5obmCAjHMjK8R
fY/h/8j/q6fYTmW9zw5gxiSdIqv4nySKROo593+gqic8c0d317YlnCjn9k9JOksm
UBho99KTZJPUFxqAY9N2mVMrftSsJY9RQ8LcvLWAZwlRKTk6JeydSoM3nNhIR+a/
Umhn1NXw7+ZJStSXEvWoMXQUzqwWUYYlNjN+ymzAx+A9+ilmNi51APD5v2ZPy0ia
QS2BYIINn8t/syQYPqomDFLSP+X7j2OQuqAAMfwCiaSUhFLTj4keUWPvCzotVVnO
k4Y0gcpEafNYFhusM4T//IAJ6oOfLjXnMXStB/Lsc+aYmiW1L0LJyVa+19izT9Pk
f7m2AtCvKUMkHhhON/oBKK4kA15L0AXKfpISfXQkLCn1rZzxhbJgEqud3rZDkjCJ
811tqRkJH5oGf0cR2qwj3pUj71/LTuGV8783mHYHWobq6ChVqYOJBz0Opk6cmr38
MGxN1iYBrvNfpn2asKFgHEHbxePA4wTPXMooLFFK/4pT90kq1gUi00TCM06bvOZl
IYt5zYuyc2Thfm5Y2rjAEtOaG7kvZW9tSsWyOs0faIAZ8TKuWsEytylMPbwcgx0Y
PIKpbrtbbSs0uAq1Puqw6+5ZaYdZaKBA13e3gMne9otVZKP9l5D00RED4TZW1AOl
fK3wu/f+MUjOWip3HM2PvbbzF4Mc7JCkzpgR2/ZzOW79pneUmcgALhTrdFRKAtwS
c1IbwzW81cLzUimb6dvaW7u3nbzZrDitjMPBjybVhrl/DubMd7hkWOyfISzvDq3T
t1KTfQexTt1vMq1H7DSSYPIiqnViLagzLuLo6HUqREVp1zRFomo3Y6ku0+Jh4PDm
3xUIPsC8XobEBSAvR1ukbdFor/DvRjHhu6IydcfLrzxdlsxTO+5xm7E45KuABedV
9/7EJ546Wul0+U2FFuv0Wl2VciVTL+n2PfnTjOU9eTD81g9BMAXGwR+5sAQetSwe
GVPISqnANh3qq+z/xP0hxf1TEFJj4drqeRCnkRU/te3Oz5Uezy8as737h0lBy8D5
JW1Bw0Ufm7BufyONOvU+hdUdOMQ5UnGqjI3qVqa89fw+MQX2J1xoTna+SMC11dm6
i29DIWnNwsYAUGCCIG8D4mb3CjZsUWsUOwDXxG4a5wd2090eT6fsHEpLYqF03hPs
76CMZV+Snf96BGEkcQNIRhtGo2XwtcQak626qnvpK85thNSK6O3zYduORZnNgJkn
42J9mI96vVon12ZteCHglSeFtE46+AKiw6o6qT/C9sU7MwsF+eLLAyf/yODj+mTx
l/fLF5+u4TB2tNv4tmpnsVB8ABxdJF9q0OIacTTMVqKHNw4an8/ExgwXITK9gC8I
2kSf66PVMHFeh0FqXorA01ZsG/9SyQY56B7HqSXsMZJHsD9itCFND/HB7JZgRHV0
cbSQP0ec1PZCyib6dEc+drVTXFX2B5LwgrBx6bQhERnt8n1aLG1gTygUgTlBLr5x
jxvnhfQFPnpHp9eFSQ9wvy0vrsmAsemaujA3eTm04I3Kgo1ymGbqkjnLlrKn7Wjn
ToGtRxSfrcbH/+lR3x5ZDm5Fpjv+OOp1gvTsO1k7H/7xIQoIhULGLjNE7cRR/pia
LZi6abk/ha6I7Ez7b3trl+QmQwNF1N5miwjAM9paP5VTlNiUYfP3BDdZmk8njAAr
K4E7UYW4m31NI+STxJX35lQYNdioKLKy4+Y5/alVX0pF4ObNV77MZR2vL8tGoP9Z
zMpuY6qE41UHgj9T0yUjtbhuwWfdsdtI3V9GYTeRAobZRW+J4ZKngm0u03k9ZAK/
26V8RJ4EBVd8lq8aG/WZNcPaOfMtuE0BXiYbcvKGSI8h1w00JhjtvruHrbDNXg/0
QF3apEovOoZV3MX0MKk/DZtcBCf9Eag2Y6iOKuDYLDQd+tbHAVXfbqY7G4iSut2r
dNPAttS69Api+aRYPlV/EkVN0FnVp3ZhMk1lzdmlEbFxbY1EDlK8Ty+1Fv65ckw+
6d/JcNWr9J1LCh8+8zOWKMI8Zm8TYJhATzsInfC55HUEQmUwnL72KDuVQ7N3KmCG
74itIrNxuzc83dEOVYMMl5StS0BQxS137EeKNP5Jf7LJtwboVcfR3iocJAms9A0p
uJGVXL+YspvxedgRxdTbeawH9vDUm57VF4ZnYd+h58MFHEJOWfQ/DL39uNHvioa3
TGMzcSIB6siFwroqizxTrh4hmaVJ6vxp/sI/1M4/F8x+/pK8QEj9FekzxwBUiSlV
LBrxhlRBEkV6aBhVPX2v8DItaYqSuhXzxLPElisH7KB/dXEDvC4/atcFuxekaU7N
0GytysK8Lo5dkSL0j6CWLkFzgQFeYWj3F7bKYGk9VtyPDujh7KcnQCeMvjJUieLb
PwV9ITMr5+GWPayAQkEPd7MMkRI3EpF+fiGpeMn+mn3v3WGqTYePuNcjVCHdpNIs
At1SX2poK0q15DtjEsWPe7efHS8ARVAQE2kAUEGAvBxU7O3fYg19UeyNf7ByvvF2
o0ePawKCKJmhX9itk3qMsAmskAXiSWJdv5E/nF4bR5Hg1L6akV+IhOG/SrRiSiLV
Fujb2zgYDBL2IGELeODXKeAROi/3DBijvtAlbDLz8b9Ckk2eX4PxrTIQaA6lJ2iv
uqdlAVjTHPBdBdWGiHD65pYlGw9n6cWxOe/uHNGNJRexL6y9SJnmdjXv8h+KPJp9
aQQ/Y7YiNc2WoWt4ooXlN9kgK2Ait+Pu/OXDYwb+g+8Q7q6f+Bl5gDahN/2F7TOp
nUD3i3RVU3hgnHDypzl4v0RYektAiH6t3voq277in3LgdZhxG0kxkP9T5SWUYsik
QhhvGkzcVwMfaOZZAFqCr8Ey6cSdgqe9eitAp8dC77ui+LPl3UgULLUZGWZdqXm/
8zfPLNFvXozPVfvVIZEnnKwnehUgoayxgv4RasTupMALRoUN2xj4fgk4H9sVgMPI
LD3fWMP2znuLib/gbERu8SsPB3iWDdsGItChdx7KDGkKZplWbLtKcmpEFTg4WhLn
v4HGmL8yyPtxm5hXxoTvasIMUxkYEDUemOvHud1baH9D/koVnnOa4rNUGFG/N+GM
T+bgsXhSFPUmexJiZYJnu5U2Cb/Wx9ALjzHr+Vx3Nc6aZT2tmmXdf3OhhMMl9j11
/RgwW+HVy++LGcBNx6qCMPwg4CxbjPp/EaFaMJJynTw7nAVBsCKvxaZZLIOEGFBU
uqJw5KYm+yvxiPjIX9C3MkC29TYl2x78V7ocN87ItdO1Pfz7wr0Q/MOsBZK6mkuP
Kdtq18sG2atfzkqTKwv4rAyXd/gaOMphMfv6k+o3cvhzO57J4FL4RzebTD1SJLIg
EIsxYfHoiG0TNqUgasb6v6qBlQvZDPXqPSxYe5/KrgoZhM8tP9xy0AyKa9x3IKvQ
TjfHg58JDBwhoe1ejLB/SjIbkMMXGn1/d5xw4Z1AD5FhwQcj6OJPhCVxbsOdf92+
3eOntkpk1KD3Rydd5kVTBs+oRBJ9yOQtvXez1jVoIXbzoq4v90kcbxGdIT0dOPjo
YsaIpn2M09QKAKbtjC9VT3o5eA8kkUTqkLjuJGL6gwyw1LYqkcvvy7WlzdHdYgaN
vfLpMRUWtArGY+FKpBTqgwDTIQ6mm9sL3wvlFa7n+ivxziigZnICOSt4unTMPDTB
7SMaOywx8FH0wP4Vur798E0mX+8rwqoeAz42gwtDMV3jzEoilQpil2juwGmwwWrf
4TbtDbfdWQQTeqdM27XOWCqtczTL+gxUk2WyM0tBNqs5dMTqHyaa81vgQ6Lx43c1
TNUpEFFAYhMsXoqRp+UZqDMDhaUAG5qMfy5bZWgBX4aDN5bXZCNOXfXC6yjxnVoR
qnBIcZRXRXBA6X6pOclmUUmCLd1ySvld76tC/SuNLARX3Cxum8A/S1bv4whfy7wG
PACtK3aoKZcOaUyrM7FnaRZkzcsr1XvJk0RBGfWgtYCYpHVqZsK8E/5qNXScYXwC
+Hb1Ee6x3ul4kixO28nuZJGcNfghx06dVn6ESH0QSFvOEZvuNS7HWDQ4JjVENB5f
bZeD625NkrCPSmokFJAxdFiB4IE5+jc5gfACAHQkMCFsRPmiA27aJy6nFQmvcpaJ
6bs54ADQ13ZRsk5zzFCmBmmB3HuST08BC4OimSBQO4Sa4rZ395bkHrB4SH1jjTCF
Kah4fpd8GFnGHytMAdJSDd1aR8tT2XI+koPzHUqq5eK8wG1XpitnQX+f98+/zhP9
o+VfyNJ4hai81Q4BSVtQJbLPMngf9WrIEkh6Oil/k3ASiGNTIagbjH4lw3/FRyz2
WoMYOvBHX2UEePVunoD3OkBIal4UJJhpAlxq4k6u8/H8/u0LlpJlQPWN3SVH1doj
9Y1Kq6LWTOUBXZPrKkNq+ZhWoOQ1fAJTN1mv5PeZsqHU8gu6ZW3xjOFUv/yvzIUI
RRgqbYCg3cNHXYb9K1Fdp9BK0qp/Ex5Gos2C3zC4WbZ4zQyY+SKQlR2GvsCbJLMT
gVp2/rqaUB3kkS6aUPXQQCBabgMvDPTUYQgLs73dfrVXLuXLPLkMex1keR4ZcKTe
PSUxYAgcKiM8qAdvZ9AePQr74+tgLd1LzXu1xlIuvfE+yahuOvhKo+pYOzw2JWtu
1T4lKG97280Ai3hqHSLHIpmZk1iROuvXxfcOtprViX2pq+9Smk6xPI7axeXOawFI
6Y3UkvaIm2K7nZCulsk9Ukh8Raw06qM01ND88pJv7NF1nk2yZn7GZ528sQ3uKfiU
UPFv8gdlL20VwQGCPQuN6A0Jpc6ucHt9INwSW/vkonKzbEfBivavO1F44NvxKRnn
nUBDe07GNZr01Dl9trd3cBiKa6tEzxhMWhrVvHG9ku8GgfJlIkWelHotgML0IoOW
BmqeySjIiIAFsemfJRmoBibFAAt+vyUMaEuSOYyOECOstoCG3zuyUpIe0TWqX1oP
rKBxUjUwvVM1n1vCiq9RDdx5KD2fAazKxWygNYlwUWwh6mscsSMwI+xlbTNjFmru
eYxZ3+D33Hn6g7PCmRQR8jhqyr6J10ojDuDo6oXQPxpn+Hj2mzfMzA1ihGfthkEo
/Z5aNPyLQhJt77ee1p9mY8f488X+yvWodCVP4QgytZujkBrJsOqil2RSlrVV+9lU
bDhNm2rQX6j8KYjdXC343kUY80gI9ljkDtHdcbbOfUrGvP7hin7gey93ki2Gkopw
rh2EIMoJ2BZCL8y5kyPvqA8ofMZBQ7NhWdPjv4SegIQPwD7Y/+aE3uEE3YXacRFy
Tluhje9vNZKhtChy8WFNHbGg6VHlnENjBsWqhaOyaaaDGmY8Ekk5ooqH1VEGrDwu
4OixZa3+ZrejZM3nttTP3LWjRp5Cj2qHbZ5xIaHtHCfOrI81E5YyfPOEaUIvwbXC
3uxrKZEXvw42CVxdUVUQvnZ9v36u8YpaGpUEg/N7oZ1QUwWqjv0gOrPc2IGV7dsd
IsEjWIK8clb+AaDRo9FaNxz1fux0OQMg2XJIRh1v8bp9SiYWK+nPbCrFS2Tx8efz
+TBpI5D8RL3UZCfXDlTWHiXiaeyEQSFTNqW5wM63mbp5RHhuHA66HC8NvJOYC/JB
DyJzS+c2SRCM6fosiEQ4T0hBNZmC4DGifYc9EEQFhqhg++reGWq8ZyHxovMpyDqC
yjW4a6eKBXNNRGqdjWrlpX3cakwNAscz77toqBJpaE0h8qKtE6ApMEHH3cZefrkr
QWI1dMTiJu+7+1f/FSaxiPcsX9PspAXLPsFp/X/GaOUL8azbvun8Rulg9oCoUdVZ
9rqm31q0c8/bqRuUPt/UHtDTCebfKn+i4PhhY9yhKaLoHYXbeoOxwENgErdAuGX9
GnXeVz/+vL2HrIqP/4LSPi/I/RPM4+xgJTR7zHoDgw6igdeOJB6b7Pi6ienNhDip
uMff3oOK/AETkkolyP1Hkm9XeHbE7ZSyjjUwqN+MWueQWIChl0bcGd8gX0vAkQm2
MF5wpuzVm+RT2x9/DinTmXDWmWYxsRJux9cvc9Rku0Cqk2mUAN3VgdcXcNh8YCrR
x1rVXCQF+PWiWKQZFKrtZ3Ktb4PbPKcXTc2TdeDtSeMX7yBXbaSjI8oqV8rOWT/7
7MItxO1jm5QwnQQ0PNbFuBN7HoyH2LTv2+BvL2+AOf8JbT4tR++5skBhwhHiDItG
0gU/oeEma14wDkqqJagQ9sBt37mimbJ3eX0MDBhWpx7q/40sL6bCAU6xGfLgV5en
mkIxjpaYt04TjeMjGkCJcdK7/ifAM//C3j98N8Wf0ke9KCugbENKpHSJMR78lHcb
giyXNATx/jB2UP7tp2nZj1pmvbZGj5sR9ba+WuySKnRCj3VXISYOSYQQzlXReqgn
oBS9b7KbtMM4YHvgNoBMEb1rFQQUYPiVp0Ut2COf+gEMDnU8UlWueJ1Uq3mwWvX7
466Yv/zZgIesOzhLgskeUyAqU4AnRD/IttJaOrVVj/TZEuziEu5/bq0rVL55WnVf
TdpLwThYkaXchdFHavbdutix5SnGQfyaNu77mB86LUk2PyrdiJyuVAbYGqCN51WH
IkDqbsRSWGLrOJY6I/+TkXAiJ95DU7NyoouWCmt5TTRYFDLj6+ehWNrn+9rlKsuk
1T+ht/tscVkYGsiKnh+J4Kfye4G2nRknZK8VaG+m1FGI1BlEj38Yqs52Wf7VF6+Y
3kL3WAU4D9nt8uIbDlqye+K8MJqkAQghl5aq5gOKjREffYQT4KMfmf3/qJ/y7qvZ
9sTiATFw1jFR/FgS8DrvRdHymOU5RYOU26Oc3a+F/vczYifnW81YJDTSLZ1NzVgB
3zvU2/EtQPVGjaAdCm8PdPedLJAFKPp3HZ/V7aOyGaHoYkh3ojDaep0Zu6rA+Yg+
GVS5jDreGzIb93TqY77tFPPXnbMH91DJ+uoeqFjfUEkPzXMyXxw91sd5MVHF9f5n
NyI4Sb/LfU04IGnyeJ6csuThwZOhPbAITFJmRbcmydZTojVqkwtUZDMJ++odXcWZ
iva93BCx4QfZdtSVMqTkCKRLwjKvL7FupOrWxU2lbdwSN4FBEGrqKeEsWtGl2Yqy
ywXmbdKebFPrQnjZsDoH6NzWknOPAqClHq+aaeIRPX8Ij7kSMimEp3ug8Ksl1QiB
9MVDTNdi9Iny+Xgx3/ybs/TqVmAzLZD7Ers9oVyDyaG6IvSSOYYetU9tj1KuVwK1
Q5tnUj1FxM17Avnz9Vtt964DTvYDxgRqJYrVy4gowcCsl9qxGhGgmhljGG0IOtUH
C7Afc/eapMIH040mlAUwW6sqWbHplfQoRdh/sEyP3ZjxNuu4Jpa6grJGR1hDlKcC
puA+QODnvLFUs+4/EzXGnQ+W7yjyGZvHgYJmPxCl+iSG/U7x6LFIAwYSDrqcQyqR
q77A0Kyrb8b8ZdpisFXk4uIIBntucw8IMZ7bKu7HqBGbmzIrScpeE0Li16IsHNDm
2V6DM0O95+MVFz8SFcSVrq0CzV3Ie7BXFSXf0hWPc528KboO9viLjU8usGlzxAbb
7zBqVtlJSVvXnjxJW1+NfEsyezffL7fO+x1SuoP3j42hI13MGD/xWcwpWQEv4EI9
wLM1NTCWL6QjN+U2aZdp3FNiPA6ECDFFcid/HNMSZwr77H5Qw1hEM9pm7WF7Mwbn
U/Dm5sNQ3xb4xHfgWDPpmeqaP448YNvo6vOj5gXLdRZ5/J8sAn9msu/YSNfQtkF8
pjMtTEzRgy+N8jdU4H02Ja5A5bEzKAxG/th7W/qrCJ3L+iNtYQmfI7C7UNa+HUNx
khTQSyD9oeuQx9U9cKEKKyz8PckNce5c2ivM0gZrNXmm2mAod5ZJLNo8K4e40ePA
NsIBQzVulFeq7DmOj94wmTILLeQpv4QCZLifszMO+9+Do2RLWBIczDqNA5zR8h0W
k7cq4A9nUsA5TgTpz6mzIVrc0Hwcn/hC73JDBEv0VamYPr+czBux1VoHBYEwrd60
CQ1hmZUhQciT6PrOKFpJKzyYFwoIwoVYMjKWQU8o56/zoxPLlYpUD/nQs9urK5mM
qttJYRVXAnWgBuVpAyxG6uwWcvyT/BN+hoc8lWSwcsk9B5egcJPdBivwoiVXwQdb
BjrDcA1rwXYXZBKZLnDRPqgJXofUQnLxk2G5UWrI/TBGn8fklUS4HLAgCG6vXGzl
u5tyJhWnB6wsNCwqDlSogJUFckPfEBbHSrzHzRYdT3krO/+auDjfVRPVrE658sIA
anDg/cxCdwXpTMQmdw2w2hA6LAfam2BkSdkhFLIUE/pKkEc0eZ1NOMcHPnMK0WMF
AsS/601C107e2fREhDJPDVWE7qvgbiTIbqn7JFXkWipfzlRbqtGBQ/cIPYulg+DE
ICcCRWhWbFB/9gF31OhYYkVf0Fn93fW03SzXPrH1WxrwAHxeghgXSP/hBAIROhg0
4S8cUKbcllScG1fY8H+EimWLf/8+uZ1zYw82m7JwpIdzxhlWQt3RZlYbzKo/gZXn
AJxPW8OjEk+mtX5s++Ok/Tap26P8SdCym+/mwDj8iIenGC4JNzvjj+vCVAt1tNDS
EBa0seK0/bhQGOoiWoA7GaY6Hoyl3o3wPk3jm03qktGDaXvxudG4ZqjcifTZ5XWD
l0DMggjcEmmmqi3EGEonPg9JmbBD+tEVJGTWUoFwU07m5dBbacsihsqsYmosXeh6
sH9AiJf9fqRatGL3IzVWqVhdr7nB0hAWurN46rvEpjH1Oy1e0MiX1xKj+Ro0EC18
XCh9fhXUjrhD90YeMnAHCkUQSL6E+Ppq8SiNNbSOIxAWrzFYMGSVycYTQZhhjIMr
QifVN72Y6fj2HNMgNakAM4zR/xiRLMAQ+BqJGgYHw+galSlnVUOUoP/qiKly5GNg
P+mZwwA2z1vwifQ8kduxhvGwnim7ET9ZNSEdMTBnx802sDZSW9m/cHFKjT5b7uNb
Q2Q6kKu0GeNQJ9vQGPCwczoxZEeP/AJAicw9/VwS7NOn8+DC4OaOzQuZaUy63QYx
HdzEgPlm8RexJsk4dcN+EjyfmmNKUyMkWkQ50m7RVUEg5xmtf6REPALb1AEMJuK7
nB8r+PUJ9p7xnW+M13Oilr0V4E8ZHeHj67kKVw7RoW9lqeZZLfx5mOFFvgheXKQZ
OoLNPCtuR/x5RnNchyZhdJ8jRBPZd1UokS3Vsgxxf5lMVZmco/t1vaK4l54ZVc6W
vloyGw3l+hT5SPctxbBKp5Sy39VO2IqFjZMCI7e1o1OZBvHQsSy/yGimNtwXjrFP
ee6a84PFNAwsfaAQpiCkDc4iHGhOSIGhGHTCZ79vx3Rc4Is4fZ0+GPWcBLE/BN9Q
YVvI4GaBXOQ/br3UsoUYThLBqo1KMYKsqTg4z+qbWOxQKWXj20ISylZCiZ6GVf8R
5nUQgKu64kqJZCkMmbONXy0SmCi2dWZ4hse2NMmaQAWqYINs/eIiyKD24L8evsOr
DdpucOPuqshCa6E8E0rN3tI6yUxFIXlJVY15O7erR64gdwFNjcxHpQcj3S4Y4d3a
j6wAChl3CR5XQzUD5Q4DrXxHa/0jxP/fsHdqUMIkdB6+eFsEGW+pR84QUnNUimVR
1uKEoGE9JEXrxv5j1QyxbIienevG79+6wEMhozyJltPj7E/upM7uOZbptExLD3RF
CN3FC7kCeCZdLtYVSCgRGpyOUZDu/0jH5gkKegQS7dis5bXdZL2AzXQByuQyde6i
OA15VnV2Ksxp5QvPeeKJ3ZUanb2RkrAq1+B9Wq35eVhZcf1lFHrPANS7ps9ZMJfg
glXVvYNq1PdNdmk2shZMfD1J4hldHmhVl/5i9gn/q1zSjvon7gWOyND5ZJKDbnOd
Mn/dV+mcPKMVrap4qWEvbRjRoujmx9i2WNznl4U4IuTydatJgEDG4WcM7z4TUpv0
vPamsIOtVno1TN7gnWWYrfqJahlMPNWiwbAi6C9cX04B+R/Q5r9vV1afmTeIeFYm
39/3bHCM9tjfeUcymgWaI6I1H+XReRAQi2uL+suan123ZjA5qbvgLGTgZlz3KI4d
mC87zABBDAEcgiKGit8tOJqwgaTRRCbpi17UqjlrTUxCPHQAUq4MctNociDv4Yrc
l7jQLZd9/w6bfCDskplipfLZzvX8ZjVeIz2yHr0LUXZEmpbymxqdILEmFPF9cKE0
mYX0XgyjwqTQaIKxotOGeFAkp/w36l78tG6E1/Q45Jytb0tDsnSCdHjU568uN+cV
wGTs/2A69Xva2GBA3gKgihC63yhXzPkPCKfs1Nj7CkHwPl779iP0J7lV5m/29cVD
Kz1MWBn4jIGn2IynazrI5VE4wagRJbFnNuE4o3q7ussd67y9g9666LoBmLwqQdDw
Cr2luQo0Dx2S38P+it3lmPfA+UbxMLN5K/jETskBCEm8nzX5EgawKpmmHEkc5xIP
detNKW/PAOFdgBNRM7inl669NZ/iPDyngcC3ZGQWVtfUfgSmIUGvZS9MdNbOJ5tF
Uo7mT0Fp+QaUxgEI2qNpBkV526Xmzn9+Oolmxcv5YFhsZZSgL+f0mGJLSn3pgsns
4wo+s5XBVcV4BjciqF202ySeoiCS67dpCcmQnXViXOi1kNaUo+J17nfsc1Snx1b3
Ynh4e3LGaUMRlmQVhb00Fd9rVYSKPQ2ArInlgowKxvJ41IQx9qmFd8K+3szeuoyM
7a/aEdzANHqdNMXaNt6plSnzhpfdiQybhMaznXLx+Q4QGrJcG0Bpw/fWUWothinF
k/17n9KxwhRlAVMreUiOTUJ1TZTe1pKlbiMfZA5ngweG76cTZTr4akKkvUqPzBxp
ZvoTbo1j9tvfWNGVuDFnlKPE3PePFuoQS0ox8iJw7VKwpeBWEwo7UIS98R4RUcEc
YX61Amov/y9SuhPQX7/FrRsWuP46tTVTLnGnankqbDGH2Of4IRBkNBR4aRsRgOkN
UyuxqHC+eUgSWyln6V2MULBwxrJZkRcODR0HaU0Rj9SkiX5OxR9XxtCYFjXJyHQf
619QsNzONtLh5SqJvW9oIpd158AEdamVZTGOl7z9ofq1xw8EPlGzgfUtA+uRNFCU
fMni+DKR/6FFN43alE1CccJJytIQddQ1i30SsONQu+vg9rzRxlKZQ8VA5ynPpLfk
cgh0eIuLc78xWmxDBxqW/a6WvmmZ+x+bemgUhCRSA1GU3nQODyg+rJfBWJdLEaWE
MQrv4wjhZqFZngNODE3Lu+SS/onQmv+oNeB28kPz8Miq6y38cOnDToaZ6amXHMNK
Y/YaCUQdvxvU0f1zHVU6BnELEXmoFdN3d/8flMz/qMu1feMtjjEGNF0tfcPnYka5
shBSOd8CIVejAuxSDThRllMMpa2r+Cn3aLYSjMaxkYWcXN5Jaj8nGR/tCZ9GNhbk
Pl05qeCUyazPci3y7MKEOsEIm8lw1Z2k+2gk6JVsu2oilmo9A+X4xbRXxfIwvRJv
gxGoy9yol8mzSHqj+JQtow7iRYlFINqwN05ckyaPtqIXPM9wnVVo5xf7ugIJ07HC
qUjArF8xVL3YJrc+Ts/BezhTp0ia6ocpUPmJ6ZLDhtdU2MPFcxEETOOBCpgkxOS4
0UhhLsPCGL/VCW80XfD6QDAn+NdaJ5P4UPbronos4fWs/v8Pcp4XfEl+mxkzORaX
pHDq1PljaGOqoCKu5anMHK+zqy6VHQTispZ4Yw/lwC7+Fk+DjoS8HbyOeD1/J7xy
O2xcdbmw3pS5950G+2TbK5n0QgHdkyoO8ZQMiB9OJvrapaK/HdHvdjEOrvGsMPnb
n82aaQocUzgOBwT4JRJ1NWhmcj4emERJRFZMJyziOhGmbLF6SpoPU0qLWrt/JIUT
D3L1RdYqCuFYwujjQBGP5Wya+PSii2XeJczkD9MSjLWHf7gzWMTtb7aWSWFBK5Qc
seoT6c+y6QhbhxC52h9kJnIoP/7GCNm4drimTy/ZA1ZbX4VxJudN4AN+XEa9suwz
CfJPOaRnbEHYIRlB4w/dl6Me78/IfT3AgWFENcPUGGR6XKxs8REVkoxsQ1ulgj0D
J09QzYUco8cHo9U4Xi+QZwMQrh8RpF9xmddNH5Pz5sIOuXbDl/F1jy1xQiK62FrU
lfjEO1MQMvFzfiir5ogyI7NaQRrSYpRGVmOu5TCuuoRhmQpaC5ckeNKaESvYBlkQ
S0212ydfSshguC9Ta4xXACpdzqFja7btuaHl3cnMW3fkVwxY+R1TTghPIXKlNSJI
qqK2VNCcY/sTPctyPRywwFCWc1qt1IwLUh8szlKZuDqKp2StXthjcGQtD/BfXmu9
NUSb+e3lJvuT/H+ycq2ltXXWoNk+oNVCexFvSknGoYbnC0k2mGJMF5iOT8L+Ny5u
EEQM5Bnsac9uyiMN9xPLTzmFKciy8vJ1LR0htlV4+NZ1mOQUrPNX7ohjFVlgCf+6
CPuO751WFvOYpAjw94CU1I93vC7aVUxUGvyExeYOSZi40YID4/9LyHC3OtAQHtxP
5KpcG4dWyx73/CW/3OVKx/KVTQr5Q2cSF2NtPkFmhvYryLLu8LKHr2MrBXPcgDKq
UYjIvxDn1B1e86gjnF1YcNRStwLtI01g6suKS3N49RdZ7FkkQag25JXVOYg5NNCP
XvcIytSDIufmqPBKOfx6ngE1XR7dVqSuHmLe6N5QZ6etSVtYwjAEEXYdcewW1wDe
jowEzZrudWFII6hiamenMZvGqOFNpSbLleBeJ69jTdDGhVKJ5Fc6dCuHsNM1kzLO
J73T+zVFg+I/vVugazMQPzYDXj14C2fqJh8xP4QcxwyH/RxSZwGbd7MntAlKr5Xm
3B/FuiDuQXI93/0A+xI4l8uPhkXuUgRkWAOj/X55D3tiH066S6JSC6y6+BgKd6Ro
jE2vFIIA88RrUnEBEvzoa5nnxp6tkcXArufAxtMdw7LosQNG1UVW+13jXfbLWn/I
tD1m78RdbKCZZ+9u8gN1pl1o4lPeqcRihwwvLVlrfjRsmm590euRjaGU0AXeIEJ0
NwdmmPCbhQgfEcWPqdeIH7trFtmB8bvUsi+7giODDLmHU8xzAC4rpei9L+3kV2Fg
+QR/bmZ/T4wpG2RiT8o1e9jcE42Z0rCszt7Of47ucYeWszUDaFl727VVyEBNrI6T
jvmlj4GIz1v/Ac4TrW0+nPEwhJgvXATT8x0iQBo/PozSQE43JBcRLaUfMnhXQZX5
ElThbmlG3n32/NpsGTB+bJIJWM+yeMP+G6yd3Sg+GZ74wXf9viUzQbCqQSRwa/dB
FY7VYY8NWpnoMtyPC1E/byn8cdeNm1mEsSWdBcKcMBChI+TBvVk/s8DHz999Syui
ZQtGTaGCJQGHcWZc03VTc04FBDMB3h/Vm4pWnBni7OejXLpUosOSl6tgr4WQkx4C
D2tyl/BCSLsZ1Lr8tqsnZcLRhTwE2yr41L0+7WuKBmJAQFnY0C+ZJLw2Zwm2D8hb
lgU/BoZRklevMtlKvf3Bq8ZDaD4qfVx1T8vFQKCrVxlK+Gn3tzC6/bFBEJfONOBO
tU/rG4iVeYIFz7T8kKj7rsoyVw43To1NaqzYRXmtZkJk2jhEvucwBI+izCcUifGg
S/PLfMqEauSBvne2xUactev2ese85Lf8WU72iqotgR2OaIncJPA/zc9vC9wjG+ZN
iyuWL/3+gMLGWmavSCy5qCH8fnTcqyKUXuPPje39ZfxNb6DSSCM+tXdO2Lr4+cfp
lc393XkASY0dp5Xai+v1MklpN0cGf/Qs+J/1qTc1r5AiAgF0KcImDxTYHEOxnzNS
Y0HZZHRbr+l0Z4qeBwpZ6BZopFgfviINg34XYl2+CsAM5ukBdEQIbwD/KSULrkEO
uU/9Rsj4aFBi+vedfzLe9d7xjsLvvxMpmEowDVlYEVx0vmm+/MV83AuUz8X7o/LZ
Cnej9hJYglFdMfShhLu9est3RjIFzFz43mq2ZftxpgYqfCDnsOA8cT/spLBUxFRK
2ztZDg+VcboEim4ayk/3690vB3sFVSVnxe7FklGAuTuHb9x+rVgAcYVKlwaD1dqF
Cd16alo0e5WUUBUUQuI5m0COas5lUBlqWIEarw8voycvmlFHurRGGNYuqX9s7kG1
gu+P8sRD0y7IsL3jhDhQQ7BnpAU8M1UiHEpgRCjCC4SjGdKMvUfHeSfVNMP8AjV/
Ds3bMMJmP3ypPG/3LjmYn08QaNjoeHrfiBrf13IJizYvg88o9zjvYlzzL81I4Tfa
iQzuW3qzDTiCoJJKiBw8VGjkR/qzjg4V+rhRRxIsiYAwEdbGqjuYB0mQzGHrugXH
ZHjK0/pGB4R2rrZsNlosRTLkPKKzRloq+m/IEDCAhSgIdEVb+lQhzHtNZmLi4Gpx
mxI22++jMqZJ8n/g/SX/6gKQP7ekkBe2L+HwkTqvneMiaQeMHG+xvOe4+TLVHR2V
XLvroBn/MuascAMqr0nke/OYJ1WMfI3CWybAvlzTWPsIhXnK6EvCHg9MiLGGiEqt
BfTU2KgQ5G+x7H6UL/H0G5XkyzRC4pY8kGWcpNgaYsPKt7/PnZJzpiazYh7P9Z72
b6wnjBxbeC7mdpzt5zN59m7b8Tl18pU9I70cRhtvuYj9izVKXw/ScBvvq0usbl4l
JAodRkczWO3Vr47K9mi1DtGXPFRyJDVwKP+95tl3dPfXPM5f+VQzhpDxfq/i68zH
y/yAnNl/PoSTTisIjt4cAKkF2fAaeRvPGCC72Uj+WFVQvPkmMqAk04Re0JaH6Di2
VLk6xThO2FLU+Jm14DjNRhza90XlWS9Vc3iwvhHqpefDdisARbe8LeyNAvDm0Mv4
MlVTVGrWprD0R4kv+L0kc/7bAfFbTqLmFBrZDXGmOifsPkM6YB/82tgwQasVtQHv
dWs5ORcdkZYYaANcWIgFjllhqFwxHxcX9WRApfYNO+uUlI1/TszftNAEhUKgQxjT
RgHnKGfRStTHh/SxYqtlRFUCJa1LEZ5jNxPQpRqyBoKzeNWtGIkdCYUwH6h2iYpk
9ian1HFcI81cOZ7ko5mOBfXFV1HpruBQRaDkGwiyQ56+S9cDTkb9LvLHAFJVgUIv
0L85HfOOtzzOrnmYOgEgQwPMI43frEYfl+em4CUwbpYlI3fcITyJrNjLH+h9H4BN
PT6Pil2Hl/k3OxKnBieTUfVJoFQ89oEaUaBhT0J0WHOZp0mbYvnKbrorOFunlF0y
qT2aSBouEmkULzPv1bDYXxp+yguTyhiQ9zauzsaYk/Vzuo+26ZOHDQuszprlCs0E
6I7VcG9v565GJ6PT8l92QIfu16Axk+ZU8Dl4q1NNihZNcQ4K6ZIXKQKFNeW7lu4q
nY4KSrMlOOaKKd00noo9ymxn41ciQsAD3QoT7pklzs/sERD0bmx7avV5EhH4gDbe
OKB/ViKDaM/vAd/Euu2nwxEtPG/bb2jXfoRRf6Br2kqeNQTPeMzBMMQ++zJoRPts
gukC+zFarm8E6QyeQnjUg8SRuK4vGSjTkg3Fx3F351v9aByYezCAy9dbcO0mRN/V
GZTWq8X3Wtx4UqeAlCoGf9GzAiPQXRZ/IYfON33bb//oq6FNJ/zjGs78WVH9uXk/
61Ndxo5DNnrq0uCfAdqjooAumM7G0WKiSwQVlHlFVXf0q091QdVCNmOoGSlgxkLR
vdc/jtRugroizrh3wAeFIgBUZ8ezFhzB3VJH4v0B1q2rzdqPCih0k6mWVWwT6Lh2
PF0uNARXJkGCNJfg1fQq8KOTEeQ+XNkwQA1BGzJ4sLQNRhDHeGLPxv9raPRTVpNz
+IG2anFy3OBQOJ7yVEkSeCsVRjJ9ovUKNAsOSgT+0ZfO2bhoInlto0q8gBkKjvfo
IyB90lJAzZBwUcxiAIwJiztQ+0kQ0CLI5iWjKI39WkelQ+QdEA6YDg5db93cNfqR
o3Iqtpy35iqZ+atG7xogxwtLHFrwye3YpwUh3k3eA9WuVrznH7i89npYaEcjC9X3
Ss9h5S4Gmt7TiOKu1nF4F+nDhePca63hWUrm/niZnq2Wa4ivoh9aYU352kCIXsAR
1wlBtCwwJ6NaVkb7dEnlrLsUZzY7s3NMZVJ8ap1eT9R+d6bUAI9LE3Yw/Jtiq42m
F/ExaDZYjtJOGngaLb6IDuI1veirDumOx1kHZpS5p2jA8RWl/culRqwMlqo69Pim
2kxmE40nhFMG/5EuGbAAoDh2NneOYhH+ycFT0XjnSsAPztEQpoaeeBSn1adSZKgC
WByR9McXU+bn3M4B+q3r9dObMtCBsAGyj/7RNkYwfZ6bG9o1RUtn1cBHmWe5mQjI
XMcFjsTpS/6vKVwhxNxS8YFsuv0jrpSYwBaTGnLieXgDk5IKZ7/HFq67Y3M81nyo
0/rnaCo7qXoPL/j9Xh++bNXzEFq40AGcPwhDv8BGCxtwvjx7LVRZrZLO0ZoFcQeK
xqEsRyIqsBT6HATNVfQUdYjPPI2FTku9DnsEbVzfWUUs9AHrJW4YfDANVwZ4nxaC
Ah5d2JPgi4o7xsCfjG0YqNQ0iyz1hax3IR1HohxABZsXF88XRsJCBwweapC3fooE
8wbxNkj4yLUbID0UBXgkTDIrE67GbIn+0LCaLc8qeSir/cGda5o4jtJ5VoGm4VrW
Rz6y5A34BDoXR9Zli4vx3VuncsibTQU+ezvROYK0AgppKGRn+hHJ7u9QTDUM9xRx
woMDp2HfGTwTozBWfNGeqXmuEVBOOJqKQv+k/coyEMDSl9kyBKYfVWJFdVOU78MS
K9r6ZEpw7+AWDiHLz5kFmvLK0Du3hkZGQt8GkY08yHFNeGwwIO02ZaN0hyai8btW
WTmUcGDuUF783a8cQDVnMZ3sWIVquPCmW3YBxWSXUXIpFYC8uKm62VY+/mp/wvF5
ftjHjL9gJielKgtRrtPUu+yLOAu9ZF7frrOOKUXQSS10rjxRYXTDToFQdB497wP4
V/MKyIUZoJ2Dz/2h7uhO52EMQKn8+bG+3gnnIKTBLoS2O6KQHe6ThjrNvm2TJi68
bEbRUWxEHVqNNiow4RnQA+/rdL25RMgYOVdvBJyR7wmVwCs46tcAisJKybUk6d4C
kPomgh3cphOiqCA1m3au5WaUaS4+YcBLBHPz+F2E/UBFEFZ6+5c1mVgmhvE0GiIQ
WO805sAsI6j3fKsMiR3htHT8eDvRkSMNXcNubXpiPnuek0O4hv7AHhtc7PHIHo/a
AknUHSBLUUBLyef0enqQmdvGblmfJayefRqcBNeu63g4kTq4JYzyajZFZivl12/b
w1cajXsSP1zKwLRQJx6pQSHKZQNmfatsrbOHbBSt5F05n6XqpWJUpa0WtUMDJ7WQ
OIkM+Tlv3mYcVb0aST/JxvpZ8NP8NZdjyJeUZ0oestGGicYNdJGQa1F2MZANfgcv
7X7vfNVju16R/bO9KSqG/evG0PmdyIFUPvrqVmnbQSL5eQiwXD+gEjjt4Eikfb03
IdiUutkc0E295dNG8BxVI9UOxjbJwmPE9RYMVV22OYUpuU0HZ7XgJW69RUYwi5Ck
KwqAMuX9vqlZ47WhpLClF9RZ6PW1wbJvNxoP0l976SZrwV7ywiUu03QdzmhyKDb2
bljUdMujv5isMrZCopj1Ev44kW4JN3pMSQubfdKGIwi3mUMoQVXKHmra6Jc4fCQ0
lQIIru537Tvs9GuHCcxNN9aovyDNy5hnhSwam3D5XUQUlSkgU8pqG8OCDMWTantl
79+JxVDYYYaDVXa68OJ98a3T8eiK6Yb/+6poIm60RAa0LGDM6PLiWqVcUTXavTjS
h8VHp1EbHGccUfzIn/Ju2fezS3QLFVsMjZz60GguCSEevGYAvOIiJd8Kf5MYgmjt
jDx8g5PxE9orNP3V3GgAuoUYwZOgVyUDHZ8sIobLEe2oG8EisqALMglpm3+oRGYR
Tr09cZBJ0Fp425qb98QBT6Mz48hQ6uNZ3fxIVBibI/XMUii3jeLxW9ESaUHNZ50I
242lwJghCQEuVvvA413SqcaOO5sbz58bVw0umwMY6AvNxKx7sRnF7gmZCKaubIBX
PXynzD8IiRKl9qhfnCqlXEALfH75H4tiWFdD9X5dVTG9BMnSbmwvtCsn4b7AWwbm
8tzhN+zujM0AuAby1ZY2S88c/JJO3h8bJ/ZvVPMUZwILaRtNDwq5LQxQ2nU0aYG8
Nk6ZQft11OA/PHan+hj/3p6mL87MdN9pZDKwWu8K6hqS537TM1UZW0w+siyH31zu
p6m8lBU8bLkNUYJifBOH/uSTUU0EB2ejzIWfr+wIxghZYD4E1lF6RbNvTJ5FId8X
VUaCfEh865QPF/YRBtzljO/YTqQpIl82BhJEj67q4y7+9K2LET/lEK5ftqhWEuhS
9xWezcRTARUXkOQbGOYAfyh/sXPtt3hTY+gmaSdz1XKZfEdAenmTL+jjRBsv9FGE
5/LaN/EYFb+ZLfySA0hNl9faWhdzKwIBgBe5f0UXRXhyrhexKUcjvKzwH+rRQgsp
OHduXnN5z7nSfJv96saX0dLYWElJ4Rop3K/NgTEPG0MvBZQT5PQzRQxNTCrHVkVc
BeNhyA3WiUl0Fzb+v0g8P0CmAWwE59J843mf8dfvpx2Y6KuzXlR20XoeuT6weZe9
aDe9QJN1UBkVaave9MRQhGE8Zbdie/LUlTmk1zL6AXRtSA1vM4A5eNKDZHNtaRC0
8vA9z+EVYTNOzPDTrNoIyMfPIeuuLYheQCwB11V7bTesJvInoETLF5+S5+oJ4EuS
5KtsMzgwORkdeKoJjaVc/J+EQGI2HoaAzFrvxnDLue8eDryzmoGye1JF0gCyjaxu
UDxSO6wvzYlp7TUELtnia8lR+dNqWDAHDUZYM8UZuP7WBIc+5PEFSvuEIPjv+8VY
IqMbBcJ5jPA5LQ4MlrjCH4Nq3gKe7Mj2fRKjVFebQCsQrqcvdRNiN1WMwV4qEa0S
VGPVwPa4lYJSMDIst21s+UuiNjchGUVb64lffmaA/YukiU6BrVh0owpWdLmFUYrF
J54aLVMzI6TUzsg1yAUR6EOveBUvNMprWiz9PBDbwnl5cdQ0fe4JlxvtgV1lelWt
JmcN9RvDMqFFqfFu4MiBgZ6IZJ1spXUlgfmO7aDcII3Ly1L+PqsSZKFdskZ3+r26
ZbAsbIEzZT3CTPaLQgqxLTKMIGdxdC+rG3nW/ng9KvF/h0H67VK6Fa+x4fp15qNt
MYDjX974lpv6ZTp8xSyhWeqTk0fegeymQ8ZUtPjGk7qrsX8pqv7PRAMObm6kA0xd
z9vpgGtHu/dTgApfYFCEkjomIdnjVWLqGBTfJSmLWExPvi0Zdgx33gIIOQHjYu3M
EcZdD/hHQgWIltVwIV6z0jsbmh5tQ5+9/r7o2n4g2FLoZbaxAZ/35ggozdEox4Xh
78cO9OLYZofak2/0dPYLmwYB9aI7ZeV8/Bf7Im13aSUm2hLHrNqxATYXdXN42bqR
vhh6dEjixnD8/vjZ/padclaHq6m6jrEQCMfE5+aRxNS6gspKenV1FJ1ziwMX73Dw
Mo9w41UBe5fIz2xOZ7X8UJfja4r/qiKTRwmq+D+y6Cq2f1hZvJ1cpVXFHOoIVsSr
2NLKJT+sI0UOACS9El+2yga8yxNLRzyX3+38FK9BDjPt1PX+kVNRf/0/ObWRjc71
7ajM/hBRSHnWRKtn7IaaVmOBat+mDcb0/MXrMN25SnrR1kXzTVk8eETQ98OJ7keM
KujDP//sQ2phUUV9KJwfDQso7dxueQ+cj+lCY73puyDThXPsfySN7CAGgXKqZjER
UBs+u53AudXbC7u7YZ9NIj36s7JWNLEsbhdfLWyjrL7lEvTHCA8Etr3vIEfL+ir9
7Ek+Zc2i/exCMkC7Zcwivdp9UqYfQqLT9RtZ13ek529j+FqCfHDf+URgWXL+dMm8
UyXumEBkmdQiapMYI++1mDpkhtXjfB+rI2zFyfBmDqPakTka0gUS+BYQnPr2gJzS
SpjkjWfmZ7eDj+8r4aDRFIVlLtYbWMl3WlRtpdrd0U5vEghcGv//8TKXEnsZrrMU
GQX1ek4oaRFTGTO5UxXoJwbSUVrCWpxVJZ7CkJrAQ15oW9fFTlCER4vWnl1INygK
W2s9Dtcn2jwALibbRKK++KbX6f1P4PN/Q4qLWGBzdJVS8nHx+VOd+Ly5JX/9u3dl
iXupuQWMLsvF6rlPBZRtBbitp8JtPuzCMpGoIso2qfOQldI/cU6nTkt1prhNIL/N
kEVG8th/KFtw4Vlo02PqxByvNgLFQnHIegQSZmcJKtm385u4h9Yf9sv1XwBuh2Ym
cnp9A6zPd5HvKeXaKj+6D/gmzaAVqLOsyzu5OcACDxEYNPm+TURW6tbS8iqyYWqj
yZxX8RDwv4e4drFN9cMY6TM5nY+UIdPXdfAPBR2qgHr0OJctrLbhx6fuWh8SKu9i
7bbI+ipPWwpkuB6KuQzcRHp0jlKgaHL3MY1U5k0z+sz7Q38J6iqGa8CIS9vfJ1NR
ej3HRHZvlAdmm0f5tiNTmPVV86VbyhQw1i0ZyzUMYw96Lj36B+QfZSjwnOds+qcP
oyOzXOlaRh6YPCfDxx1jBC00ZUepr8PNq3RI1WDnimZZ2GqkqrBIwCHmXQcMZ2Y4
U80b5VOO1Oa7CexyxNPu1an4ok+U3u05/TcfltShznOKEvHBa5dQ7RxnHcxm4Bo3
kim0xzMKBrgum/Oe1LTAtYOux6/EPcce+IdQd9vXP2TN8nMd/1jvcveDVkmXe8fP
Q1WlrfoTHgRgbhWYuCG5Zq3qdvtgaeClBa4ylXp7ULytkT9o7PXJNO8FX800CycS
p20QXIcdDI0yh/1o76NG0UEwUk3qAtBeyJUmHu6D4u3HwH1wNoTaOuHhGBc1ywHh
7tpjbKIaM4rSnXXNAi49YIZrzntuPCilBD/oeVxC3E14mU8mOBJsLiDhUty9GcwT
WX5tN1UbOeBQTCOZqhUiDcu+Mu5sVbDcWS+WGmsnJEBlFQ1HjsDlXG2z7tye4lvd
7pGIwrP+WnTkIl84yCp1gzlSAuHks1ci3C/B1vyZ/UjWJNG4VMYIxzUubbBPUw/F
0XqqxkA+MD5tol0xBmNAQNSfnkmJQIJQlU8I/sy56kEDEta4R/CQ+iZhqIn+1eSH
qpuvRpvkvbMZbwvhrSdMkM8gtFwFBD53Ix/gqAtM9lcI4e0TPJxbqKSffGBzx1EK
b9B32kQrgwEvz3xk6Y2uU35Qd4EgOssT1rCU/UdLqP0h1k0S0Gj35TqFy+KhwDS+
jL1QCvjlmMe8/CXZdInyK5+ZUuuxHybOAQ1bKOrWoZuTCxIM8Z6b6n5RuIPAuaMS
8uLn4xF27wlJbCRyQ/93LIppdFW0lXT3S5apKV2SfX0XOSKnPLfdGjc7he3s1fMw
C0ou5ki3b/chYJd0KhGOa6zuWjXrJ5V877OX/484E+gT6WParpr5/g0vO0E8y1NG
090naE7gjNid5ijZaBaL+O9PiuVNQ9X7a8X8tHQslsuFFBON97VhgyPKZFkScecy
HsrCqvfP7MU+Fjwr5z58cWg7X4h47K1LKnKs6sXSgCV5EMKA8MZCFYB3xhrnZLU0
EzNg4E0b6piC2d38Mewf736c6ixkj1X9pOI5JgHVg3VGj3flUysLBt5zJ0cOZfOk
mkQT2Qve1DdYJkf+YXqlixbdnH5i9dAMJhLuySM4grpXwCz0Svbq/bLrDDJkPNup
eNbiof37GwdhrNvUB9eMhEX3pWcyVARNcAXLDZZ7mT2kUD0e0SNf+oL5XgCBqvBM
kR1sN3I6qiJNPyRiH3KeAPNtgmJnbYnBi9QvpermeMcWBkw93pXM6Uzfq55cCRko
Q0uJ+Wq7axCZqvx2dw87AK1jzxFC0aydQt24vn6nutCbgC02uD6Ns0RFGX3Ufmt5
+GGZ8ERk0AAK7XsbiKHhZHIp2amrgoZMxZoFE44DpDlM1ryw92nGN5+Ic1Kj2i11
zVe6I0g3qwX7qhcvljMmdefPPH1ssmsXB9uPXYOfJBji947p0H5/gtQvW0KMLxdF
8eoLyH6HLHb0EIyU6mM+fH5ZupcxitNFQ+Z5RHmv8w62+WHu4vgZkpRMJnUNFKys
l50gVfLLcwQ+NzGW7vZQphgKgg42jOUYhU7oY4V0AdwDpLt/t2BjzlNv0z+jcelp
9fZztFLOV9Fo8o4diQWUohVWfzfGypvaPA435KhyKAmAtuZn0ImTu74JGH6CqhhU
eTYF9g2QmyvIT04yc+TCd9YlgVkFKuH7jBdfOUyxSYHg0nA9hhuGFvpl0/3A/0Bh
j98HmJc0eTM+1Qg9xs+NRggUwTcWRDmYFgVwtUS7A9G5lmZ6NCuXyA1BMUEufxH6
8ZKKAHNa4NIfy+z5PpmHygxEcxEajStcv9O5iU72VjL5Z5QjM9XidkusEl9mudmv
E3uVbBGgHb+9ai4Qu+NYGSoyf1GSeiSzbTWD9+X5lx89gQu7AqZCAO3g886IdgDS
vBgXWRbITrvAcOfKI/1H/eqzKZHq2JXHnn8jNS2htwkzusHzL3DHunBc+bTe8OQy
kPl+h0lv6/Kh/a1GxHaGl7ha6otns30gdDvcD7xEQuPRkL3WeG2mSaBxV95L4nqa
XDQ6SbC32vyDhc/qe5GOmt3s0PXrGz+GFsCAkEnbgCHWx36WFknHdpzAKwLrrJ0K
u+EsPthdhFtXwdnalkMVhET1pvFVVFTviJZ9JTMrwIHO8l+dwDyR3akZb4BEomFp
YFcoO6pdv0km0vjScywEqpGVuLmoTwlYzROIs+RGV+EDOUWGkJkuGX7/IU+eiI5b
HZj+ilWEtCZS+/LfUTzU8r48G+6ZER3DjNV0JvULYPh0z/XfFMQ0XO06L7koskeq
7wgYX1BNkQbWIPMzu0IzSeC/wPN0+n4I+cfPl6ifmwYItgo4TMVfnELFkHzOpc4+
G+QypeYkGg5m3UxEjQHB52bQTiO5fc1l4v8YvrbKRB+vpioLtbHsEZUYqzmc8tkO
6211ZVeKjSk/vs8FaGAtu//E02XCZ8oQMg7y+S+jX0vA2kJsbvTIG/QgDQwQsnN0
DIt60JYxwNjuVAwvyriJ1v7dJOe9Nk3l/VZEI2dRZCs4rWiw5waTxx6krIysjKt/
cjh/uC0o1gjDUvtnhRj8v1bC9NCK1XQmlk6Qc9COqehSXogVLvqpxPca9hLeFV1i
+qkwNbPBQbcT9wAA4pXaRF+YkQZ0heuZFD7kXhZY52g4Lgy+43GqHFHIYOVTBVs8
Uf2x2VIUpNpx0hNIP91fwDqzpebPkCxZ3JARQBeLfMKR05gMYPRZw1DOfEn7MIhs
1zbVvpIqLPNwaB5cm97feVOtLWz0HluhAZM+FNw4ymSDmn1wPPinlxwsMdi2jbhm
Qr0NopmczKrgLo4a6jMUkxCGLM7++NFBElllWEO6fX72pbMLSvlTNheo0a2hpQWR
0psFA7QDLxd0yYimSDY0GGPNj5nlb0zEQN4/IVTo1x3R3fBRhlPrx1vLrYoADllQ
E8gHDJCtJzdieNNO7BA0rKIP6615QhtrXZU33xt9vM2cbggYajFPbSvcMwjPjOTa
9ldPo0cKs2HKaWuOv5526/5IkXijNVja7LWNJlN2r6Iqn0avq1ShXlmQCyoqtaaj
3DwbMCioHnCRObezrS4lrQSSobf9h8tnfLRsyDUkIbzngdXpCTF6OCAIJWtW3bSC
ubjhiVBo6ix+0ExNIxotquFloAOKh6xhsqai6d1yOnxru1C9zk2zONg424iKAEbz
um9OUwm8DIcAZSABYP7wl74HY3JC+jPktkXuZXtU7czSsIQvUAx89C9JCt/Z3uyR
RIdXNKuqqjdZLtcHXHFpqxBcprzy6h/rdZvNm5EoL4Nox7e5vPrpYGNsnu39y5AQ
+/QDyPWSEYC/09uu6DcoFGvZ0Taqz8tt9wOqs5tVfKU/Kk92cwIAes6xGb/2f/J9
r7v1ZYDAwxjAMI1H9+HBPLHhYZayOinA3PwJdJcWH5cjz/ELw+JJYIIKq6n3Uwjv
K3LDJhfg/NDsPGltDNpaFQWcqD1XrlYfJxuXXaM/ZCbAD1LUWmQcs3ZxlNA9vYzw
q0EUWThKIMIdAiqX2ySRRDEU0mLThxiMQJvUBXIXAOh58xKqxIAeR/+NKNATVzPX
kzFmq1gBbYq/OT7ANLvxi6xpQqoLFez85EwHyRMINYi3F8JEpD5F5joRPfn6fgMi
LtQPUiXre65ytLsDJLczLh6ZrJR7NlHVpTdCeGHC3CD3+iA7Bk5yM6H2icGNUkjt
yh3n1d+kOVNpGYdCURX1Lw5chzcBV6wCdTHplyij/ln+81mHsP4zAmasZWYTXerb
+Z0XzS3wcEn7DibohA+xXghDpCR70SIud/MhAK/E1PFKl9s4k9dht22vzN2mctR/
S9jaeaIRoG+4tbmq+PCXHM+1CzeMLD4TOmpG8dsd4etAWa1bs/8E3lXE8jkt1+8y
uUMQMVU8wABwjcAoLfCEn52hYooixNwJgiP5xfjtayTy5VsEESJ+KLIN3cTw2Ua8
00fYGgehm0Gq0ceLTLWIo24R94ntSx5sTMmcJaKKb0411QH4qEBO7+SpdNVd7An/
nRfO4HNrDIE9hqHlQaqAEmw1pgZzqcatdCqAyx2LCJsVb1qAE5icqFB+UGoizHaJ
einm/dO7cRMUhpqppHGc0gR2z4LxkNRujiXo2qgDw0HhRo00eudZ14nPtS++SsrT
sZsBfBodsS9L/NKGBi/DEG0V/0QemtR/fcBqjxhT8ADrdsYqqk/VQ1MW+DeP2RBD
L0Zvp6WPxuKWzxwsoksyvot881g0dnhdcJ3HYVQ7yOp1VvBg8Lgx2vLGTQojdfak
6my99OyQXwkbGDLzzvxUE5SlX2JLo2uiuBuntVT0/fnCht6Ia/Jn1CE56nygtGUq
MMbWrB551nqFb9FmVKmua29iqr/ciRbKqOlXmhPOJkwPa5XEtLM9N1Wfk9funPyS
KdGmpKO5V42rcz4ygBYT09MxapMOFT+TKVlP225qzy3bqyFS3ndar05ZZwpuDMWG
nH9bCd/PZdRTHIshkEBu8OwR4RPVMWaXqQdztCMQ7iNVXUjrfgdXogXH2oeXOJQb
r9I7+0RYFIP7OygAKpbmrU1p/lH+JOdoxv7vzjOSOtg+t5dXnlcOGOqbXS4VsNux
AufNGHTU/JOoSCsr6nZGjwpNUmMwIN7nSsGqMGMFW5wPkak/zZdh31xhsynbZ4+2
UMoeGrmjnC2hpZrHOGzo52DnMEXXD0IYuYpGm3wX5/64LWXYahuJM/ibmCkfZjbW
27mCBo1QU12fQsqDl/6IyRqImCYu9e3cCF2sjSm6NnlK3FA/tZdF91Zaw5PLNYjw
4PWDfu9kxduvn2hgAkn4t7Rf6V8p6ytMdGPT0AUr2k9+tD3uxRMD4/7UQOab+t9W
QVqxS0fMM+1hLVqwO1e6QLpr2DTaGp1NKH6jMo9Tbtl74QzyAf4KPBiGkPhMj9X6
z+Sk5kJiE98LaUmNbrF5Y4KZuaZP8avBzAPUQZo7qCVEASrqZMasS2+xakFl8Squ
sevcSep0+78EsqwGtqyoVq4oFJtWDwugEq3OeTXllx2lMjut5T+81ruuPfAw+DMv
wokqlJVfAKsXqXglUmpa+EUKsz/MKZAkoxcSCTV6pTqRQk0WvBIp79SktGEoPoFv
kRT1YHz4zsCdQVWk0HWEZvzhNZVBT7W0JKqHj3rmSIH66TPGXyO4jqzwUrypBNi0
RarqOeqX+zdnoTOBDdtkhnxsj9ywxt95+Ok6lFDVPqDerrKvq5uM74riL6WfhkYI
xYa6oDEo7oRFeRs8P62yv3XU+xFO9C2OWzZCj33fw1k/9fSOmzeCX0W2IjeLhXYd
CP1Ea+uymY2Y11h9GnG29K4ioYNSFRQjK5I04A9gv9lThY5vGjz9ay/K1/YtievT
udNIrqFVQvLBmxF/YKtymwi4ra1MK8dKk0vNQ5j0vOHc+/wpYCPO4d2+lqAIMCge
oGAeBk6DE+CKK4RoyJ1KZ3F1wIkDjm7ZammDaXzwzkRyQ5QWy9xKCmu2mykN9Khx
xX5nte6o/5qQaR7Gsx6pMrdwx+9iunmWYoK8wkdaywmJF2dlQvWhi3hdnaFBCXHl
EUCf1pDf+GNC1eOJTegD1Hln3W3FWWXTK+lYqFfnNgLpaXodxnb02S+QqzT2+ca1
aTbm9Rwrv2NceLABCYzu2ME9SaOh0P3xxg/9imkFjg+FZ+LEX8ZzRhqFv57Ay4yK
NR82B1RST+to0MGcKSGyHKSGun/99z0Qw913Z3Gvi8N+ijuDeo+LkB9nRE2z1Wxt
xTZSvJ3G5jAZndA8UIqkeCdwzdEhB4/a/sykatkLizTna6qirq13TKmASu4PLG38
bfEyRGjNd2Z2jA8kJFWlMEZOpGg9InVhcFsYnt5dCDsoINWlcGJpTVkOYHF60VCK
Q19hVUKv9z+X78wsKKDmvVEqCJq0OyYRFdg/5fXisRHg5FzUjL9fMLsqYTJSaFrR
ckTIQLbk+VOh/5WWHcmi05NlFYvl4YSn6syYPDLx/bChMbnd3mswwr9f+gSdIgPL
v2nXkRtKDYecLYZFBiJbkq1H8V+gUKjAIeJRXHbw8e2kc+oImgvvmhFCvUiHie4J
g/5OqGM9yuK8fU3uKYY3upqaskS9dL/qd5F1v4XQrIazKhU1LeFtVgOZda/JNvrI
MuBscs0xGSXM6CA+UaLKK+sUNOeGmmVVIRyLPwaqrjG6MDqIwK1OtqY+ojc5wCJe
F9ziSbxk7SIT8jSkpF9qtTjt1RS7lZUaHjhQ5EKrxkoG5ycAmukTXIMLQmyWNgEE
5YjlafFuhshsRMIBfSp+Fp5TrdMuWsJFQ1lvwWI3I7zEkGWlGpboShfmlJNQonw6
xTj2XOYhbUX5is24JycmXOUgbid3H2HP4xu0m87bW6SB6ohT7qTSW0c2p89sgxD4
65uUdYE1+ONKsOJqm5EkRNCjiZcrTxZU/QgVRoMMl5tL7jhdb7Fav1Xg5VcftaPv
sTg26Wuyzzl1W9aSGHP5hwINHQRPSqs644DTRa37gOIwLoL7haVJTHvNupkqYqs9
i0dg4XAahnMNrdEOLZHVDQYPYEKSrpNQtA9iaKqraTrUYXmtO9WxBEjN4MJj/5li
JGHFyJdhNoYXtt238yh8VsyVnsQUdomhMK0idJhsL1x0q+kzS5lnFuTDeCLfDh/F
GhvxxoZ2rb/U3SrEgHVAB5/08yDUyAxvwuBRY+bG+LAspqrb0eNh4pdYiID4KU9U
iDe+KgLiId4Ny85I5XtGQlizG1LNgXkwCtpkECNkrHd3LtTNDPSQsLi5/DoWAxlW
UkzPm24whfcMGJH8L6v2Q0EOvyQwpEj5FBcXM03ZUUkIz/A9J+NIvI59RS6SelO8
/6jXgqWka9K4s97ZZYvIU3XDbXNXVeiSZ0Y1Q4johQhdvIsCiRsevrzpoPIa5OIw
wvTIJDVhjdezWKBYquYNd+AwTlW1ZCGlxoFgSIrGD3TAf4Oyv+m6DbV2GSpYokbe
Ba3a9VjXSIoAU/RUpZaEwo8cPZkM0RtBJ8XJDU9V2AWVWJOqp48fKIKl3zMXDS1+
dw8V1BblMrg7fPMgmLUvI7r52l4kw1BKx6E2Fy3ac1Nj3I/bQ2EZUIWpDLLtsvhw
ts5k7IiunXoV1pGxwoIBTT+5JH9RQN8lMU8az3pgpsBYJHRL+gQkLEiR2CQOsZ0l
Yw26tOCcW9pwfiXXRfQtiXdh0cTDFlvOiFJshKD3gAWKPeU9U5PX5T1xIZKplDsO
MNoYTUgqPJEcZfDG3+AVnz2zXC+wu0v7IzO7hmyw0Hdnivgw/60fFsaXCvFivo3c
hUPhL9Yt6ZzGEq0Niv0+PfXFailI0MN4VnV/FHl738eiuBQgTBwY1Zk97xLl/F6w
I8EpqvDQM62YgQmYB+yxr3qEZIqdYR2/UQPrtB+KcHt0vr4s8Fh+cFOp4lSgM1jP
uQ1+YtRYPPhwyqP95khhpm3ZPrd7ZwBJSqkyZbJqwpvrMgsI36qzsZ1z8CobVz6G
AlwKezWiUfWvCsgSoxmKe8P3tzQKudDc75eRund1bkG7NnO47Ll4EDUjjhJr8wmQ
c4Ht2S6bbBpbi51AIS47ehB1SF08C8y7GvAtSpOjQjV5WfEgGFeG1VPYhw3DiYhk
+pRr8uH2mVvHo1oAsJpiScJ/OdXbmC5KGyq5wNWBG5rWL9vbLP7VCe7As7jn6Q+Q
GsqciU3CWO11ZhWqIwRc7aqRfajYmj6Y2Z7XV7EXsA0lYXI7Pwe4LEfSM45T7YHS
bGfDIpgvoumFsa9mqA1fGtxX03IFp9UxkEQk0PTV6HLjAJZVMONu91Ca/SzX4s/R
krAI+LC02Nn8uSlvL+2evjE0t/+PgoYu1YsW+XdFSkur+65zQ6W67yaairyYSusT
Y54U37K4BCOLHVGWf1Oub6V7MfnuJ++stDnYn7PRJsTrYzJgJPg31T3KIWsMSKX4
Iut2Q18BJZzO9cAEQCzX0MGIOHmnBczXgK0tm2VVrpmeAGv7zk3M4WaBXokPvhA5
kqdofVqhoXuPl4Nq2xM6j2LWY5uHJP9igSL+QvtPV1pgiMjPzSjtrGR1VEQyE6Uk
Np2b8M90lznxyjAujL2gLbl1KUsC6qpH3Dvo0wyGmJZ3rrYF1BvuckWQYkttRvgH
mOaVy+ZKsElXaS+LBUqzxQ8WNflGsbxRUa014I3qfRSFo999luEhQtGwRIGSochl
sZ+2rPZVtXS1Wx1QhSPxWyPD6b0NpB44gCe+syvxKGk5Thu0gNMT3TdDWl7sXHRG
mdC6IyW5UrbWqbO+O3/NOBXB/47d08OxeSZ9cnq4uEtaTSSeSuC5Ec/2af+l8pYB
PT2NvPsIR1eSKx9yEOKJDzz9gEVK9Tl/A9eqbtsoKrge6752Kbl7BQin581l7kNs
qxZykzXM+XcEnxG4MC13hieZYCm+MIt551RXFUKKc9eoHQDmruPZvN+GHruyz99j
2jVN+9Z6Edr+uTJmu1Y3tLtZNb8klFUDQ3/EBr1/VWYF4wJf4UGl2dxDJjlQFWj4
qWSiEJlxyzPnifMLnrH34dG5VM0lA6YRUbQWJejuouketSZYFB6cYzbCqbukA26E
uHrWNAaBV09fw7Y9D+i4XvmtNdA09K8Px1z74g92FoikszMxkyKq+7XwDGmiLinX
mdK9KLKdQGa8UoHdtWZk2nYz8RJmxYqO0GP8X+7pr4rrW4jxfhqDp3321UGfOEKg
GEcbjIlE+GRuyIboMSA1wEMbK+v1ckO+GSjXkfbXfETUmXNCXCY3EOYRJBaPtJtJ
QeVXcvVKdBeUVGdSyumYvYNgOghEfKUEt3KPBlpL0U5eDmP7XqEr6J5Lje0qGzJs
7DHHVUBQNUZK0h1H31FwOSmME4frtU5eCrLG05jRIHCEOguAq2ejkGpoAD9yAKb8
wBVjFbNFABoB8miV6ApHUMeqm/E1WylyZH3eEoLpSyDqTt8AGI59kQGnA3JQk2Yj
ylJpyrF31bWMcz4yPLVClHQs4qQmYRZEDgpdqcXH8o4u/GINAByHgHldaey+9zn9
5hKt4bD7qv6QrvjSOXCdCX7c3C9V3+XaVICp6pZesPpi5OpJ3hHXX9S8+6XtADvr
+fjb+pYfqXo7Pu5V9u+Mofs7hOSexkzQN89DsYazUt2jLkb9Qv9dUiFyp9cTgCr9
ns/SIXoH59YYlGC60NvQAO37sXCNTQoRxOZ5KE2lpX7RqH19bNZNor8VMfPnLI/N
GBwV/CIkKIVHPjv09WlFMLdtDgWds76Ouh4rSHu3Ork+npuDi58FqpBMiHigzlor
9I7j+S/8LItBH1ZZa+f0iVAH88qzV3JrR43GXlUlfv1ABwoiXyJrsT7oCmh7rlPu
Wa4zYjhQSYo5/lAvIjtu+dTAbQ5bydFDYhrhVeY9cD1v7RUlbAS6jODJtYkxDN2M
ueNAGbLZmlrq45l78l/BvDdTUbqkXLgY0cit7cFkTcQWlSX4Gih73xg1oKxZWlIS
eppazifsCFXm1Bk+ak3Hd0S0ul2yUoXOcz3CcyfR4JlRHTxSjuYYVn1eHmQwOCSZ
l756xYpfL90mMQMMnGF1mSHjNUtDl/DfJt/Qcw7NMt6IwSAeIb7sZxuutwQ4ZqnG
4FLc/T+I+U/zJ/uNoJr2Mt0ZAGbMAm3G6aPy4TQxpbfK6QGiN6TgeltVB7gUzKHy
LovE0F7m94kAt/o8RX2igUl+IQaf5BU+UZ22f87J0neBE5gh1jzbrwkoxg3QjZ3u
5DtNYLZ7h6IrOfAV6o5wKVzJwx5DVsCfuL2k8HN6qCJYZdTZAvbSkCKnFRnhhLy8
MstVSEZAd91rmDTsYsL4Q6e5+0bJ+IRnns7yeYyogyPz0pM9krSnSzW8eMrguaOa
6a0m4M0Dvi49C+Msbs0wI2Y0T+taaNjtZoN5Nltn/rU3uBPUFJKirAnNKLAtWGGe
pJw0Mh35ZuOFrcUEr6M+pxKwFhnnU1yQXhbMyzLLD9uzSIRNASONHO2T6DNOKq85
AhqVCwRRjoCakW2zWoMKd0GXkjGisqBt90u97u6Mvh181NdwhV7Pu1ZxA/kELigq
l8iNpKer18SW0x2rZnvBf3xFH06tPkRhl0/Fb71UjuvPq/7/+4VqRsMJbNa6a4vn
7voRTQISfSOysgzPPCaNoR2ZQ9UIF/tp3zLz8gugn74ERhERnGN8G9kvZwOz8l0r
HbzTx/71tzZKlUatj9eQ8rmhiKwyARrVwGqTBdjUkI5EWycvBWxEgzwtcoxRHUPc
pwKYlToB9N+ywjNBznDm+e0+x1FPsEzvb5hlkYd6vt9bBFUi16s1rxibdN8lRY/W
ck8jzE+d1t920mL1odSl0SJV5fsm9ly8vDdllsRK3s8SF0Qft/Hi/rTHQqjdCrE3
2CKuWTfdggkJaVoe/tGtkWCcfRjVCDAm3iWqAh094vgbh3WGvtknTGvplqKZY0PC
K808APU/MQ1GEh33l2QajJbIEJ4yR36JSUudIaYQfBepIIup00+bgxpg8Tp5ahjL
xKbmy80YAo+M6K1ZizXDSk9lpBe6roMBXWAXyHhRC0TeBMSPFKt+c3YMRo0A/Ssu
apQs3bNPREgyelyZisB9TX3teZEbhLMTXR0krfjIKtsxhSJAAjjllo5HcY/q36la
o2EWFCriDJ2mKIdJC4+voLj6UV4lGk9SP+jjcTHu2ktiXyfWuGcTWys2djHk58yX
cejQUKLax0yGx+XApew4ARxveRKiyf7DMSZ/naab7PzCb1262cTA2uKxARe4nkgE
LNxvpmg/6LNNN7l5h2KGZRRUI4lKOBNn/wQ7Ef8IAVTPV0i6TNB4xZZq5sf/bbk8
Jzb+2ldHR1VH/0A30Qvcoe0+JevxeU4DETcoOQQlJ/7rP2oUXWsnXs47wH1kcogy
2uxvc/Qo1tWu1BSinr+KzLZxxulHIN+xXekZdVFJM9/7KcoAee+vZjVVKIcnJEJC
uG9JfpeC5pQ605BLlU9UIs2A/+vuxzCnA9POXyau+y+fopuqSG9lDTYqUJpYJwFU
qm/1V3ibbp1yTEAba/C6Swhk0EQjRJiaXTD9rIykuZuVawv6sCZcI+zkcyHuWoiM
kzI3jD80lbYdAd6wgkRNQ9knZtZnPTIKuOQxsRuq3tveqmtrFJ6K7OlRtfWWXUa9
xBt+2qh9omJu7KcamRDYMqM8roW7BB3m+5YOQCjQdDRnYfPKTbRi7aquwz3zok3O
FvA7smhYH6kjlR4D7fnErbKzfBmG2h+3b9g6JVG6wtOIMSHwHWlpYVuJZxx0xBVI
jf6v1tqD+Pku6tgRQZjkJQ+oFEBoWyGORSoGXKFelUS8uYTN3RhbrAmrHXH1XxvN
zdHGTjxqAMgiJ9QxtVITDv0ZCjumHwq567eq9QZwlg1iZgaam/Tf7rUxyrpIK130
+TXCtytO3GEs0GOF1CcmfGAk15D/7VkMPKNCa9ir1SC4aGcR2YlD+HpNtIZ0XaYk
T7Rq9tBkdqGuToR2UjXh/1IhkrNRLcrDe9oe44/Zqx4mPaiH37X3ietComoS9dm6
vZ1h6TaVraQvJ/EDipxIEpXTugjc3E2+dpFfUD1QyrrXqZfSeOcNI6/bfIN188T4
Hh0/74iIA949iPBhH/vG3plz7Wn0wbhTf+ivUgJh/TqEfhpIQC9pBgZL6d7MOCsc
WGmsL6SX0Hae/5BYf/NtDHiz5UBLbpn/bnGwe8b37QufLiM7nmF7bRaYUeXSrCQY
SdZTnx3oWqaQ7mh9/pLdhggLCDb/qRZw6Vx3aIt241GATbmdg/YQHvCkAp/ynH8f
dbm4NM5TDEeNVrOHo53ZjHMDFnVgXmdHzai+Kyh6Cq8Xtxev1fuLEZPwEus4kUwC
hag8Tl56IeQHn6tbykoq6n0Ih6ET/VcGBxvI5tc5Z8TcnNn6hXJhQ3X8eLGVYP/q
djKpvSe25ioDZPzpkhf5kB7D/RdrX+f8gnu0c+NBHc+8inie8y2X2H3u6MykIbOD
wcc4eCMw97rdtb8MhUrV+e9/yP2wiAKlb+VVvz4XRtZl4M2/xJo3oKM03DL+S3Dj
meMG8IVxrgjtqkqUz9p8Ktn7D+kCwPb7KoF3oUcyob+z3eO00i3JUPK3RWN6FMSW
hkmu4wtC/JlJHZj/WHsTjtGjJsU33AkFqgxZIlWmz5pWFcGEYIfLOKtuvnccri2X
oya0yonOWXdD+zUt5wXddEK+xeuJKwmUxgKnNNUKNloW1aNYHsTbPcqfZqDjuCMm
4iAFVaojT6r1UG/LX48U+aX2m3tvxlXOKgoTBZI20DSUkJIRizEvw8h5Kv4AF6Cp
x/oyCU34p8eCQQGMXx1SThWmJC5d3hLcD9lS7zoNLUbPKhCusV+wBh+xZ1OkM0mG
SahLRVZuGGzhHBKHsWacB747iejrGv4g/CMoHZAjS75e0yVE7kx9G5Yi7wQGMBZU
ezA7/z9du8I727pKSE1yxZFCEzw9bsKmxhrefymXWBIjvhW4lEbj2KEAST/rfaew
5jcqiyOAlsuLQo0DUzl30dLclvn9YsFtqhngW0lOIUQQtFZ0Mv026XfSzx1UEcDD
jYPICAOotlRtW9ztY6TOdoxAoUhmwyOXlo6ms5Z1TfYbz1GOP0KftdK4MSqcApn8
ilcMij5iKkzcf+ZYoopj4MIB3vfTiIA0M/P/SPS+z0jplwTj/qbjKmEh5z35cIiS
KKmTOgT68XY4Phn3TdQvbpbgTy8a4q9mdiSFoKVHqwo45TF1OvBJwBxfKt5IcwfC
MHhatKZYsBCGtsEFR/xO+WR925wK53hpvlGdMoAu7bdNeTWj/HM7eAHuj82ZrLYG
lJQDIn7bdgqFlArJQYxRZ3bB05sv0pXIjSdZRxsOPTzpmkOPT/cNonCOOWqCJzp9
yIdiv3uWmg9qidvsjcSX0L0rPCiTKHQkpVh7wC4oVNCgorunoejYAFs8ZAHdqBsm
MdQrLDBeV8qlvR0mBsux6coi8Pqjy+QfFmz9zPHeIn5u/Q3NswO8uI3ADZsGjx0Z
x+WmYQWxLAfbwZw57/Tn3l6pThbeL7WIuoks/bEAc3j7qw843PWF7q4XMosxu1nx
wY29KWj2wc9nms9mUoFJIvh/rtLwS+RLD+yFV6ScWi7rVPORl7KhS11AsyjoyWRe
CM2LkfIQNwPZQNcQxCjxIMGL8kkoKtkBbn24HG/IobASiER7f1HU0RzwXBx+cEqD
L28Mcxm2BaN4XovEWVma5onKNdzkXxnJbrbjyWSYUUMmzAeQb+OcGnFMdsqplijk
zYfFwrxaAw6rK5pjGzWJ5Z1q06SDgvaFzLjc5aBP2H/fWVKEzTfa6bz4QunWrQBb
HuLpED1W9P+nrSHQWAsHlaEI9ATkFLNjQv9zuIx4r/WR5ADbs8LNG+FfnuaKdS4t
xaMso7ODKKAHwpkAB9LB6HkhPH9EFxVMPnS8yXGxbCkRi7ImlslKQpp9v6Zu5Wz7
RJ2UQYTfxHm7+lpDnazk8FBU6e2GPOkW+J4Ws34MXUN4QDm36unU0wMYrB8f3Yv7
11VbWaSogco4kIqXTiSZbJeQsYqUUDirpvNAxtxXOSjaPYA/RpQbz/3E3DVrH578
87C7gGfNMSHuIjxsL8KDHIw36XlTJmZe5lOvqi7ET5TPcBs4GcfRzqEYmIULsis6
l5yMCxZR83a4c5tkZ8S3Am98RaPnUwr30cH46bt9AYn/6BFJZpq97w9lRJ6s974j
M0dUGDbjJIhTyiyYVlYW+uk7oAz5F+rSPBwqqk8x0ig3TyIKpTknD9A364QOhR+d
1mlDDYE9TqHIAxjWPNB0jo9jb0NWq7fYprrhna+xY/i9FRQ1F8Bt1nCeakfsnZyS
1JKyjn/iFdtDucqw0hjfzEUsSnCo0hD38+K6NCSvDLBjlTrISLbnDQBR5s+cJNuD
E2mHOEVKtb7lrYsbyu7PbD5p/gBfA8D5JtjKw+CMJOwn7laUYu3Zfhh/b0CbxjEc
xw9EUcNSlahHXkWIatNtnZTCgMDIM5Wwo2+0rMuSBLYHT/lRE1EcK+6/nhk4uR2I
51O97QuhUKzuyIpnpX0IsvNY7tezXIB0nHpIn/0s3vVSx+1oFLoxpnRdAeDW5vFt
+ZMNG/fmTCMgZ+XqnPpj+ho5/z8rwl7ZJGAj3eYedZIUGeBoByUZAJrVa46jlXv+
UOmu8WsazW+ZIdIAnZPy0i4RyQGofv107lw5+v03GcgWaE6HlhZma7A9qG4CwTZM
NKtFWcHkfGDfVup3xmm7LhEbiIdl65mhZk8WiTOoUGXKcS2Gx+yEZOKjogPMvgR2
Pg1FYZkq8PFX1l+oPnSLLcPtmDRsyPlhtbzDJCb/CA2A55bSPet7+rlQvX/RPREP
FcLkMH/LtmCP2a0MNathh1Ov3S73rvoTVpEADUrZD6PD0g2v5fiT4lLQz1rrMOqX
tS/WOQ/L4SLD8zKpJ1wQLPCfnW2LMGCF8tpKRDVn5UF5yGAPuEjS/0ZjtB401FA8
SJgw5a/d2TUYNghFubZHu90I6OFZeOai+rnfrbLagD8ToWxRegALxp4Ey5IVKKkJ
TuoYA9MyImnqEarVKsF5fOdwDEPXvHUEVQ4vKCIIjgTKt638TzKdfAAdUWPTD+oB
X1ZIhJlBPdHA/RPLDSKF0TjlyPBC101Ce9gpwHW858EWfOm6ZiH+Q8qOy42MmaLk
gMKy8a+6bk64tOHLRXb51/qCnXX/peQJ/v5xPfQiicx0W+Oi7cDgmRluDfCWupR/
UZwfiZ7ZL/haes15UEmrlLRSBaTpZdZMn9rQsp1gNZSMWnfwCUyCrEwVMmGGjImM
OlYXR7p3G2p1bYIdni76uESwk+mgNJfLGsA+UXOOfnrhEr0Go6UJs4ocxnPq9a6u
UJM1NLqd1wHVFY/6Z4E35ze22bot3oGfGaf/19rzZNHE/5Tg09VG+A+1gVasH3iD
6gjfOAZVvDAIvZhiyXmtmk9jkBSzHI4fWUp7N8h3ZMtpxMFSCaVxYTP8aTVKwL8k
c2eulLZACr+evu7go7pPx/YuUip3CZ9vtv5xcveUx0QZXixTodQ5D/HUKwCwvugV
RvKVQnupVqj2L4SNqtCOOXcitMN8CvS0OJIjI+KNy//Yd/GYGq30uISwM/5jP6PC
weWa7Std5vLm9MjCeNFYkr6c6AhpsFZ85KSQxkO/3/DWZeRZl9WOafn7AqUMuVi/
b8m+3rzJroDoTGRvDqnmdmeJLbU7Rj+DMS+y+Pg3XY4PaVNeo8QbwxQpDGNqDiZa
aoV62G7KuWQGwLAAOIALJ1t+3v3NjB2TU1cn4q0wMw7w0xlPNp6RoLbExViPQoK4
ULXcN9MbIt39Wi/6mgUutV9qbpBCop2zOPoNF0/0xEm1Td/q6zK4AeOFEmqqgU6f
gVk0r+TGH7xYG9gEFQ3c++eJ7ADPypg+/2gfoguoJaL9Ola9gMfXE27ym5EpWaMV
+qBDc2mvCjUJLnqgUl6V4APgscxAYBsUiPHrF8y4J23ju/axxKG4kLBWNTXszQ2x
nd2mZv9Ordjsqj346K+LmttCeO268hiTZ9MNqP2NZBaNeCtbD1TC80X0X4z+lG2p
sUCgy+gHGHekv2J+jpHXwab9UY41up18jJXHR6E37A00s8DHJgcVvjMUD4jbY+7D
DPRa4aZ1BtJR6IjeTnRxLZVZMHsp3iyMf4/7o4Vr2lU8m4YYqUaaLviPCxg/Llrj
RtnKUCeK0eUClvlwZYNy2tKcrBxilQEzAJLCHyO1DO/nL7BpYqTLOTFtATd1MkS9
ABep/iwwNkQQK7X+UtabhM49N1D8pEyGUNzLN4mD45SuqUCg8Y2/xeU9xxrfKlBB
URxoWpn2A3K4cD8bb9TchYh9cK+YwzB4/22ZNK37Vxx0QcLHZCKa6jhs+foCPjqX
XqNAvNBSIPsHlpWavNe8jwBt79WH8ek+HGgv4dvw3e6afHsrtZMo2iKVFk6yZPyz
SfSH79350noOpC3Wo/pcTYcM3ivcsvOKVXOM+nai+1aBdyj7c8BmntI0K5ofqFan
W46Xr40icPCcwXOhJ4HrjMC4MBx9SlSMAiWZllnjOEkbOPsgMOjXdkzk0LpktZ2S
7T7PQ/8RMRTNm4zoLdINBFI1KF4Ezvzp0mgtrw5IuL3Iak9Crt8wl97y0Nc3cAVF
AV2QKeA3RouuCH8GwgwHCp6mRS59JA4H0YL8ZFghZgko3fc3wbScct7r4GBfker0
n4TNEXXifvZ3nzYj3e4OSmXYJkXgpsRpYeRMfI3g6xKsVsStps/p48BgMCbk0wPn
vO7xE6evNpI6c4ZVVyrRj0BspXfNxHvlaSemibGxknwxc18p6mDFW89wZ1/pbjLv
IZs32qkS5WLBnXsBbXHNdoR6+BJj1iL7QPRTNYSObRzTT5qTYmOsRZbqHOU9OhXB
gnJtN42F9WK2KzcMhBwdKRDrN5KIBZAvBgySxPhKwRVpVpMQ4WtNY/QkPqWqzbIt
BwLIjf6g35OB1boMMutT47+i0ze6kSKotiuoQxF1KhwYxm+nZ22EDUtrplXEEX9C
LXpbd8/z3Pm07QCKwDz6oyyGaeN+x99/80uv3fbjpGQGOMMg+ML2h1NV4P5HqDUR
yg7OEc4+/EJstI97iO2hBuKmMSWs8nb4ZtXfYvCTfoZJj1CmOygi8CcZ92teYxcv
aZ2+qM58CbLlBqc7VBZHkRBeFDz2R1p3iy4TigNwMAVuZOU+586gytQN0T/AdKIO
4PQWH7Oj0e+zosgAgrQZ088E41J0eCcxujXAcT3PP6HjZFU/1KYSgOPOjgADnf99
/+gr1vWmN7MmSGdeIvEogxsW2g4rlzmfRi2p/IVA8TprdHQOzibtCYB8DkH8aaKJ
VH1WsNTwxSbS13M/AB1M1ROB9ybwSB9eXyG6iNY+NmeUOSFawQg4aCQhexzG6Jqr
XRddOpMqJrSV2J4ktJFsFF3JISScIhTZVvH/244KEA+Xyu5VB9RiWiX4cjej286Q
qtmAkcYFHW1hO4F4pMkaCOwfy8ljrdZIB8m7ns52h2JG97rN9N2KXt0cIOvvSBFY
v6WC3cXiBqcPtcVXQ67TfC4OyihJDdFsZQ6d997ySu/66y7+8tdb/2QNTR94zjHn
1ZaZue1K0wlCctOXZ5wUW2qhsXh79hyx3KIrLM+c7i3gw+oT+5nmOYnTRV755leR
zGVFfsVY96QOnQgpUU65DX2fOlXnHqT+kT2o3iPIwrTir6sQ5as0sQbd8xlDTXNx
ek/wJSXAagZWei67FyMhBoW1t6cLjGcVO5Poxrd48fXk8soIwLsxCUxKjdVt4NmB
3Rxg8gebAFgQ+sGl+y/gVakjr7CeI/3xiIjUsS3xQq00q1YKDBl89tDktektpXDb
s3ZqkuIlJr/Y0sOOd95ZR64K1+Ts4LjtohWgFaF/UNA00AAX/gCq7DIPKmuGUwH4
R4QlmQ/w6uvvB6KuU/KyqjpsKyNMbnZc/AXmvLcnpaTHbxnYF77ZBlUf6l+2opyN
KP3pIoM2khTDF7dhfQiuEmpOM+h2J0HjwANVTpChUUoGtKasFVR9rI+5ir1rx7rq
QcddSEk2yg2KzD72kwoMk2csrQg0TOrAanhdH2hGL0KjJ8Fu+jzMzQErMUEJy648
bidTDgQHL2LqIB4QPd++fDS9LHmgukwOLtM4mGovhj/X+O9KktCi+07X3J+p/1Sw
Bc37nQnF6GBAuPO4gMhny30QdX/G+AliaDGixgpAD9FmyBA/U++JDEsON+1hrog2
Fho1twloDyfgI3jkDzkq0X3yu3xwZ13OkcoK11MWkD48FnYL7NEjeyuHSLC8ZK0z
Yom49MKuPk//wBotg6qxyJlSUYZdP4YbY7E2uPVZLPeysJR+afTz+/u6XuwoZc0m
0kKIV+KOmC74I3XruvKgPG7ckLWyrI4cHclZzoiH15pXWfFMdVd1xsAvDLePUq6r
+WhCmeCAyMIYPaQ/PjKK3FIpaYZwlxYlciLbxRgkqxILfdXuiXD1/jWnSHiIhflB
0rulfMWHRqN0Go882rtS6KTFs+RcWQhjv8/QqdNaZYy2EO82Jf22p+zKxFam7L5m
v7JtEEvjArf33Lq92/mB25G0C3UvNyE5nMkOeJ79swFeK8IW0dl/YxT3XTiuVU4P
P9R3DLMQJ8kKzcQp172laYtGuYUrXZejaKqv3uwrrHNEmxVUwUmGyru42xp4VNwt
IWBVE/QiVmb+PC1OqY51j9M0NXKZGb7QUxRHLf2b7maME9nKK/iUO+C0GzlrW83P
13BG3gMYgCDPuoIg8k/NZa/RSlYyjTkuDjXDBaaq7MwgnS8xc3aUSBplPymGSgtp
v0FyFRKpCWAO2dE+k7cT0ad9I4x2wB4V+CJ1FLxrfrz99KUvWXQ/xoE2zVh1kpi7
0YHzuipCfwjGl9QfktZdWU+FhX8UCY8R2FD/bALGp6+//vTuBhKqoGeBWPkJXPBN
IQzpbqcAG4ozh7u7Gg0uRbd5sQyJWscBbkkSxNRqdBhUixD0V8BMDhieMtjccPg8
0QnA5L/5wAJslfyoFJhA0WEenpMQbDge57OSrxtUzRRsF1EapRh0GTs0pTCq91i3
WhQcvp513Q6wyxsFz9U28ZnVPyxFu4X+dHamZ/xNhGQtWqRqp+ZKlkZR3nskswFc
X5wpoVdj+Q6KjxaFUSMdS2gTJQhqzVGu4LOgdbpx0AUv5Rzb5v8PUiZkkPaYUeun
DviQjcQkh6PCd9pdbSNhb9PmYvVqVSupK+qe5ZHcr8J1QkLqHgIH4GULXiCHFbwr
hmllDpd1auv8iqhqyx39XfqkG7cd95CjCctY00o26hwPTPmUiNqyKX99Q2GPcgkO
pqTcqiFLLlwGr3jCze41/2wts2LP2wjmf2z+zLypC+arkW+hgSThgkiwrMkj/y8j
RPh2wjsfu7JLY20O4pKJNaZV03bMIWHwNy26tiJsnKOJXKRtj8kVdIRxAfNLgFDk
Bm4OfsaBTDxDBYB2WymEMmWItwykMkG6fSCEEdcujBzzq5KVwrznL7Pev1G4e6Rr
60qYP8EbzMQszG8m6rLdQEvJCXOjT7Tx7byLE+hFHMd3M2+ZtwTtstQDRhRHUyUL
UxyFc/A01gvTpHjtnCS7KTaKL/nxu7jvlBQ5GssIm9Hk4FVkspoA/Tjljh2EITRv
nZA8DOj7wBBJSQC5wh91xUtK0bBNYgdTlRCPB5/TMWd2nUjzY6vmfZkREaKech/a
tqx4Rkm2pgNLFCkO/zMLKqS9qtdG7G9h6K4JPPXEikGNlxDqO5spebq7BWnLL7uI
F3MwRU7hKF0cSHj+z38y0xQ26Pp7pp6DkuYKbxy8+F5eVSFbiwrbbsw9d6nx/B3d
ae2R0/5MavLnN0xvcN5KQSe3ZQWYmICGFwq2zrb1lSQ9t4bOKtBNMiOgILV6A/oO
niwSfGTeFXncWXB8mJa41l76z4LDyn2bhfsVNN6icH6l6BybN2hAnuird3aWNisu
sxSHjPJn7qxNVjiIyx1w45wdY4zTXgFxZyQUbZDbB48NlZ+lP6ZlqJSFRDdGIkqt
ILrdP7Lu7kZuuub0wR2xcKk0h/Dct2xWG/wyqkiXDd24aMx74wAi5fHb1Td37Ojn
zdbFCOGo0zZbvUbWlTxv8ZHxmdR/KMp6fcyFFowjNt8PJSyK2CU+H57mosc/DMes
x9yZ8doj/5oUd9kWjWkmIwIVbKvk9GkWRXhUdT4ex6qN+XK01m3anha7yvX0Q8hT
Hfg9VQq7SKOCAAYX6q014Q6qoBQEMU9tDdTKphSN+FwJRT033Wfp2rElkeacZGgl
lIfnVgUFTbKnUnHbnsMEEzFkj2Vmgp3GrE7M4uaqqYujfoyJe2ZdxezrA9+XWieG
NtPSv2F8UZqTyAZROj9CTA/XKxN9z+8RGl/mSjV7nmdICehvsaHDuPjK3zUAbzS7
RKPvBri6QxbuAa1bJoAIs2sshwLnq0V1/1pgZ7nQxT03iRggdW5WX5ljDRA2QP1g
Kh+3KCGkKKAh0aQjHm15Tt8tqpVUNnDVxkiTeum3xSESiAUOZ0Zz1nwmgH1DzsmL
SQHCOfe01MCV6nsnEq0x+k2tG14hTA3AimRwcznsKGi/PeU59+1eJCoQmJh8i3dH
Q2OIm5g2p4aMlFmQAaGj4Zcp63+cvIqyQlhgpppTLfgW/ZKpQtDCdnveDdwXYjEU
DuucvY+Gi2WcrQXgNhzWqq242eXPoUTdydtAPPvzuRecKrYtzQ4tUjCWSjoSgDya
A32VKSTHijQ9UzGrKssTwdVuNAbZ83KRiK4hb69Jg91QdJidkUQv4Z5utkLCd8Pc
EefzAKT/WY3vst521ZT5aw==
`protect end_protected