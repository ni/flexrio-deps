`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
gMcHP74wBZczB0bB0IzoP2xg5wC5NPjD/GsvSQ6VQgzYAsanETMwwsWi4yhFtJwv
5kY07u0WerSDf8woJ0stqW5xF501W3JLIS8KMiCOd55RHBOnavjYiaaLeu7oUCmB
TtTS1R4sO325rP2zOn9YwRbyyS5Ljn+PzFZZUmkt5xMca3p5NGqKtZW2dV6Babni
5HlLuF20Au601B75m2nv+ZRoGSrpkNElxoTibONmX8gBflpIVE7BehhHwaKSucEF
pp4QQ5zZAZjEC6aplZepouGVggAulz5AahlX5bf4opOVlB1J7IrgyjENtw6ysQ/q
DzybQ+ipztSXBGhmcCVU3A==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="jAI3OJE9Sh00Sic4PtM/KZ4WjwT98XM8AMZrZsQkxWQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hyw9IrFLPQsjvXplweG8O0lkaSLBN9Ijv4B5VdTRt6ipKJT9Kzsb5LxCKvkQyF9n
sGPOd5i74hRHnkHfYISGkfxGJCa55ieOyFShOsqTKRLxclm4oja9vTIey6yFm1BZ
54IDCG9h3PqfDiTD847UCSMRvFssyycwv+BRHQMQlFs=
`protect rights_digest_method = "sha256"
`protect end_toolblock="BnLuc3jxknmZOyxfJK70E5kp9u9O8IQ8cgkXv26kHA8="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
xABArkLxBOK6xG+7CdOOiGu0zbCbHMrEntFfAZEE/xRFxZaAZl1QLkuFI77OC2KL
XxG/mrHJzO3taVHgwRXNLDdc8ePbxbAiQfzV3NJLBO+gsBjmIymaCa480cPNpHLx
0+LIRl85m3WFWTFxk3QeDa7DWiPaB9wwuZf+FAdmyJQLYnBm48Qe4WRUw0fQQClK
vq+H/SP+AwQMFhJdbg6anrloPn5750TH7szip54/znWs6BYy3Qlu9/CTrrHlfH9i
HbStHgiPBaur6hvxUPiD25yyuqZfTUVyMmmAnGZTlz2qmZmRLVNMOwi1+bBGqXqx
OunAgRYi2phjWk2nytfGsv7AKWPwWPE7bvhO0qzeMfg5HQ0CBT4MoLQDJhaxix4a
ZeEm77L9wjWY79PwCdWyorc6cKsf0+nEnm8YxxbCMo/RGobgJHT20HK1guRYlqmA
u9ztjWDWjE+ZKK/D6cXfsHEZWz43UYFcVE5xlGWrJdGipjgQWlCynfHdXqhEJbh7
sppsyODcHm5rIGCzo1QFohLkTAOWYKFRa1ktO0vCPdVsRwbYRylrEUncU/ZYE89M
eoN9+jtCxsmqowipUdRqzZcvFDJH79QsqbyKjHU93oaVeSVyRj5nIDm4nndJPiLx
3tTXlbla5TAmhf8IvuKqsz5Q3RwqyvUmWpWvTt2SwXq6oJpPxhyzjkKjgrJtrO0G
elb+gSzCkoJiiq1iSdmPujkYlwryBRf42JC0MHYq6CLhXTv9XpVADJOhgPsZo1+m
qayJZU6ZB23c/hF41DY1me65Jjg0TA1EdfDqkbK/rssE5hkpS+wDbkJJs232cMkc
0T6FGbu4gIi9DIH1ypjyBcPawRBbOjnAA7t0dR9N+b9gZaZti5Y4sCrIppWwxki4
5RilWJfEyj7k9gIdv7DKLZpe4mkenJgZbQYUMfPPTGctpiLqMMLMTzvq1Im7fsdx
ji5NpGs/1NXLZADIJ0RofG0797lyUW7Vi4M2Ug5rOVQRAq2HlQX7vEmIu1tUAZ4d
6XrhNKx3mq1qSwDEI0zfcPJRP8gqIJYxVfPh7QqvttkG+neazpKLIjyiTsAN/o6U
AoTCBlM5bWed3HzC7xdGSPj9p1c98DFK0X/yptYNER03vQO2pulzPm/HMomyx4Rr
IilKbsLmDote3pWULsD815ruyq7jRzFHAUzOxfds06wXxhdvIsu4QBt8goudhwrt
mVgOc2QEN47jdpVgB/MpJr2ue2xA3DtJl1mKD9CpY30JTJVQqxxTavbvlGrzdzhk
ngIdRdOS/f8PizQ1a68tE9kiZ3rUOJDSDGeIxJCzy8LyZOgC9I9TdVuOP1VXs2TW
BJ+1FvIGtvcRpx00k2MrZI9gwIQoxuyT/QtP2TKGdGeyaSWZnKasJNeTqbWYGozi
AjNWf9IPVT/O2tMMMrlSwzLHc1RIi1O+vgNMh5ooaMSoYPe+8rjKipdf9MSLefqf
hHr9VbnF1LzZ1F5FkM/7DGkJqZhnPOmVEIOGZ05kmS24Ilpm1ruOtnJYA0IY8aPh
WaFT5iPcnRILUPSk7C4sAwyNGpnc5GI6fm09GeJVmhmjLWO4f4IP+lmkMgaQsFla
wRQfL2HOgbQ2Hqv+9NpkgtHmoMf9euG8aM7D0U27VetOXY99qnUzSu0nCVK03LQ5
pnN5ahdA9vg0OEhMhtl46EidFWHpCNvE+u8mTqJqdO73EujSSixRJPnYbeZft5I5
vYVCfsvJQH/Tg2n5l985KoZ93RAD2QST/7fC8SmF2W8aS5m0iCfCbrMFupredhvl
aVYTVbrlk6Rnjhlg7ZlAcupyX1Q0KFRGGObSsu0uaiZqiSpMVM5BO04LwmWoXqdK
wrC1yqgojm3IieKapgyVzKiaNugSidZVcbtRZyjaeUD9txfjrdTNuiZi092lds0B
5+v9awfTGW4anwgoy6Ri/wfX0Q/Hy94fkigj4Li/9NQViWCvBsCodJzWMZobVk84
6eJb5GB/q+3S5+t8qOyLW9tYoXSuRkrg1jtsdIEg0nQSaNClX1XQN70XJInNmjG6
CLevFW19sYrn6JDYJpqKcfj5+/le3Nh5htyHLo+TSQbKPpyj+4WC2bqtuJsQ5xZz
u68aeB+VYkGqI3DlMFUx2etYVNWXSj7N8ryP25H4zK5KVHGisDddl2h+KzvH0mHX
KxQOCJtKnSYLjcKqTLgrKPO+z9M//Pov+0AZjbe1PqjYXufzd0K4zohjuQO9dbOO
yLY65p4L2UteK9ATe2m7ZtKwgaEwZO6AEkOo2L0477i5hNoa8Xskm/HzRos+mP9W
PydF8ouOBt5sienqQql/BETbk1krhsvD4GWn2NZYB5OnwDUSWUIWZdKeOVRsfqdU
z/x0p2aWzNyUEk+PnZEb7e4RNe6Rj5cVg1WauSNaZet7WcIhCjiQS5NtO/gA70pR
hPTA6RyWgDlwoYkuVgmXQES1iChvKsYAXwUguPlvj0XiN/Thbj0w9dwXF2q7UJa3
ik4UMtZdduLmBZK9yDfGieR9pVl0zgZInpu6Ai/yggWt+vjp3wp73EprELLn7CAP
PV4nLZSmZ2OWIswAhoo+nK5LdzvuNW5kG3oEZeMJG8s4JVl5US7UB/4Noc4t5KAs
51ZI48MABWkOskl1yC+sq5eU+5IVwhTuFT/+MdLye5lruue87rs0kTxkqJk91Gak
MUeWoiaeRVqVS/6d30uKIY57boYcrMpO8epC9hGF9uUPLPtw063Obi/W7Go0LD1W
QHYGsiGJVEBtBLFG9rrpwYFJRmgNvJ+s9HSRO0JvnChxyYU8KS57Vl7W7pRvxwzS
Jsv0es/r7YdtFPGT7e75n0PuW4gmYv7n3tntcIzGKCQ1hmY/HEHP8wstXTkiX6xj
wxd6MjZsl4LwmUuURHwGZWxIQRR55wMWpM4NcJbIgPp7Zglz6unnh5Dz7v3Z9Cx4
yi1gblqwr2Bq+a2QGTZLi7OHJD/Ysi05FmIWbJp35lS8DiIkTenCR66ys0pSuly7
600eN9Bxm3GdmCTos6qZaYJVFWNfZddjg9NrtGoqKav0XXqnv2ae942K7TIxO8L3
hWH5y8hB08qfb8qZp8e59jPrGPNF6gqAHQRVhtXXM+RLj9d3yELPBsHQTcRvpl5X
eUzDNPj2F5p5/0Pdt3oL7+7Nld/5EFxtspmvAb22UIhvzgsXLBgS7tS6S5UgjJOR
IQvZ0gwusMnQlb80TmQ18QDCcQJqcMDQWbpIj0/tDmIHAg6TtGo1w0kOPtNvUAZd
29z3lyWeuKhvctuQPCEHOgCSQNIPDmd63VEkHGSE4sCqynjGy6N1Kdb+aE59obBx
BCIVKrKy/AVAIgM5y0wXLuo9b2bDhArIaEtKTFGdqd0aMbZMKI1Hkmt07vcaanlW
moO/gRBNDAFKRRnTbjJ+7RwBR4MMwdCTEJPRawQIPhg+1CNSoJBQrpqTPHZe8agz
6zUVOKXB2TI2zblUeUwsUETs25C7zQg8swsf87gSKVmhPjIVXt3EA3WkeHRcOs+u
2IMPDGNkn1hKoT9I1LJEB6BxrHX551W36u1ArW4Ou3TaMuPIUbAPRPeEZweswQ3L
s9fx/zys6aQrCSC9gte8p9I645BOBxeqmfdEu7eeOGfx+eWJ8jJoz1t3KJy/Ib6W
gAi100v7Ljw+ermnmJiB6d6ywqcC2MzGt3N6AW7oljpGDoJXk4OefodWxhqIyDw3
OVCe3z7KVvkTNLLL3fZ1JwpYDEbr9uZEj6SoVywTNzwq/HiWoZUNfKwatIAOhsey
vSx3qjyUzsuq17Rbi1OqYeFzq2NIcqPPvEIOzUA8k5DlE8SX4FIOymiYNQmOEepr
RMG0FYzKq6JtP02TTEbn4JFQP0Xi96L3UcVD9G13G6OGs85RbiB5BZUaIgSL+DlI
8E26dpMUC0/x5h4bKs2RpSARfy6/Yiv8PLtqRjnpzaMZWj8VMzu5oVzFdpgcO09M
6A9F/n1kKifWf19phjDbqg1UDP4Zd2hufrkW66duGOJVntzo8KO3lyibkW/l0tov
8y+qHGsu0gZpb5SsriSk2butH5ndPxx+uuQEllCXcM1YR0KIwzAGUEhILYUT/pJQ
VyWQF+e1gtJfFKE1TLvyxOpUJVeRGdsGY5EEmEqpxDmZ/kLT9mb+xQcJOAwg0UsI
mtWiasMzMLqeWTqM8aeaYJf5YSOyT2i/L4acEQ4ELxIygXXddqo9xQI8J/e9JICT
nlbuYsq3u5PCakvDHMIroSNNfiDQMdcsVjKzMamzGVtaFoaTuHDptBTDGzH7jAVg
vUfX4BeqCfF3oWPKVMe3QAn/2qixHZirdms+wH7DFHCEj1xivIlEwGlZLk5GAvC4
/5g8nRfs0FXYA2Gr8cvmztrwLwO6rvs/bqTVAcm1DkVgM2vmrljxQ/F92wu6mFtV
P6Lnjhy18kk5Rn6qxvM+V2l1G+1V3PH7HA/f4+ZQM2mY798ue0iEHwkvfnGGSc6Y
ph6FUHziNhhAolj8Uq8LlZTN8LqhSF1V+EeeBJU+Xgoww2agZi68PhR5APNANHCT
79LzSVWQWKsOzkNad0eKtc3NvBFbqeNVKeYDp+UVFLl8/rf7TeE6AQ0t/tBy7eyr
IoKQpmG5n1RsKYCkOmAWnO+5DMPndeoOwRYey4LQL1vLeNMJkNlECpb4tcQe0gV4
D7VDCixDq95tB68p4JVt4FhsAo+n4PEOBmjS/hCW+8M5/xa0FOI1pYtcnIrqmWVb
RJimQyvSxtXNXoOFBgreHtYu3DuPkW8bivtDtvALVmycEFCPdxOpWyBE6pPex/Gx
vl7++H2mm3s2FwsLKZ0Y9oIYa8/L7WirYjA+LRDEkBZfpaA3J6qFGgOyWPxdnvBs
WPRj+bk5TO+gEKQCQRZAeEAGY/CtIRgibjnw/exJoM82ilXmaCwvf3KEjuqf6jLP
2U0z6UZrog1/5MOnONxuZqG9kyl6GqYJFw5gJeifWSgZFjf+Rk+mKoKVCiCXszsz
dIhL6VV6i738it6jJrmqF9WnunmtZ/snnQoIYzw3xi4Keus4c8ph3CyGjec4rJ34
bGmCSGEWQYCFo6oowRHkRIUnPDYPXRPv92Q3kAtpRboRUDvEZAPcBZf4O9Teavvp
66/rXuv8W+/Qo4cieTV4kiGKs0dLJ4ofb4nQ/H9JkO9OBDcITLB8frsah/WYpwh/
BIJAM037IcDz4SJ3OpkoW2TVdIXmza6xwKGCtJ7xrP9wQME6FAeeE8gFm8RV3uFQ
r3ap6HkUTXdnw64+/o75yISVmsn0WWQMC1DUnO7fL9vTf5T6sWzT3+FFfln00vRc
prlu+do1R5vOVm3LJDHED9cgr84P94w96/uSV2a4BnjXp0sZL541Ks5lMsg1aqMV
/ybhxRrkdYCPOcdFLnJJ1+cDtBXWmanYHdbcFW3sp1oHfEaec9+940fi4JkuCEZX
3yHCi2DzdOBdIr0Aq9d6v85EEmlIFYiPmtdDa7TR6qQYx1t9I284nns3kw1H75dM
5/xFlRpz0G0H4gM8MOSgQYyJxJ6mgx+cIpJUMiXt7XsDC3Zu/aI7HFBpafieRzp7
ViwEURYprvv9cgHpdJIqdyt18VXuy7hGoOpggG8pIxyt1SUN716cfvgffp/mHjtK
pPm5jsfVJa1ERumzSjF2bvSyYVo/M+FS9YaYSNfYThJ2Mbr3jvUqxV4e/xdYIBYS
jo076WMcRQaERG3X9YUbbk5akwyN/QJAsbzWXw6wiVbiun9n8hZCDajZyVPMCZd4
iVcjMJvM5RabNuJDQueMnT6ueUTLgl9MS/5P8uCn8Selbvn613gpMRx6ogzWhWp0
Zq3yFdBGUPlpKxfq2GogGr9C4i/A+VVgf3uY5wk74KSK6jbDfRtu5nTCfJccN06u
akHDr91DQia8JAuPp/WSq+fqyhe0U7jredZVK768e8HqgBp5L1qZz0DIov9UsDfv
hz+MEjuvpgiLlGo6pZMswwPLsgneOCPc0nOZNI99VnPhgVzCaxZK4CGi8TYVXbBu
hjYPyFq+bpeI5bK9mRpWejVmqd49SugQgXpQJC7LmcgW38yYgO12vd0ky1qhkzsE
RCXs3kvI3nk61jWq2y0lfC8IrNFbQfYTv2RFcznh313BZVRvpw0TDsrFSwbQCbjh
6E8t5tzYpqVAT1WqCSQ5ZVzxS7oPeIfWgQp9TmAeYVoq1yTz0XvI4ievIcEnP1aG
QsyIX/7A3scFG6SHHryvaBj6ehcl+iKg472Ov8+A4R97v7Qj95QzEzGPgxfXzW7Q
0sZeyAIsBJW6i7DU1S284GnTPsnn9b3AlbBwAFUDxR0Fi/0/kghpiCr/zrSGVcyP
8uGIwLkkyRblWj/eiexsh75D5yruLTRhq9R1caMQt1XDNGlz5fif/ECk3cEgORZ4
jaumU2mxFRGAo2X7ijK9tXOtcn2lwVEgILeUvGyVg/IVjHf8Jse+Trt6iegPPSuo
Rh+5W8wPAbabW3srRDfI+NEXq0LKaq+/kafCKUl6NVy6XfZXdXaC/ueoPOVcJ2B4
I7eHkXXPGYg3Pb6zNG4Yi7Z/odg1CIrKByBECI7nda0cGUfpRbAtXHrSjyjJWvnD
AhkMT4nX+tsyO862beOcGT+t9NeB0BF2sFA0us3zDnk8xx6fUjPcGUeic2Eh5RQA
8eiFPa29eFxuTsrfLGijQd7vdANqVkSRHhnyjiRCQQuUohCe/55hXLjS/0aVncm/
r+8NrEGgOp6zG/smmzHHFR8qKL7VDnM1z8KW7g6RLuBKFE0njXbuggQ/Q7n8FijL
fpAmS1hd1kUgVJr05rNmeySSSAjTkELNpkhuQ6rFXkzdVZr0zoyAR5b6WnbSAJ3Y
7CtkpZKBQAxnwLcLQNR8s5Zim2lwGR4KRxZ3uy713HkjFZKM7ThecJFintTYCOQR
Dw/VEqeyBWoNbZwRwaqEXXe022CZOavZzRq9zznKjJL/MRAsJ/9CO5MWlbwPqRQb
CGSwuWzPbELWpKs7ZvnXsFjxTqIBqyDzJaGAfyYFHJoz2aZQisSwmHWc6fiX8024
NZssWno9vdZsc/fvafQ55APUoIYSA7kA7tFRmtrfv2toTbwCzGoUS1QcBH2VPxLP
DZBesGHTj6ji6Nc0jWRozLIDdGxtEPekQJ7+N+q/6vuExyYFL4mR23zfoBv7t7zT
OYVacZMzv5jH0uKbB9tuMTPoW35UXDsI9IN78XldvnX1eq/KEICSPzeUPBhwBJuC
A0qGoPFr0sKXvJinpKPruZgh9SmJe8rDe961lvBxE4/pwCD+PAXN30JBZ90JpTB5
RpCJ9mBeyeOoNuvpQ905rUobxHgsVy4PbDDFfoQ8cZ+9tP1d13jl7gd4UlAeAKka
5nsclNDuuHLqcnC98dueV9GfwsXudyowDVlyoeAJURbd8QG8LrQj1UBh/BrCcl40
sFeRUjv9LHdGtetdCOLsyb2qrzOYyfruE79FNCaVV6SYxLwZLMav2I8ml5aLpiZM
YZV8415+oKw7k5b5apcVw/sCwU9pXHwOt6XWUwphwrxVkv+jwukEsaye6TmUTXwg
p2BHg6wBZ0BFDhocHYsdehZS1biNOUUleUunjFT5FG65seV7+nEMRQ0HbndlRGdo
nF9gqaMLoztPjCClrQGSFg7Y0JQlZ8ozss5e/8VHXhoW0nTm1I9R6vzwtvzQMkhs
fRC7EzK4aZgo38IwICI80zTo6zgRVGUI3DpI63ZRhXK9FePOmRwX0/Fi/Vyf86BF
4QD56ueZcHnYJRgwwOXQ/DJ/KSBJgpYK5INJIoxSBgNBxXblwS1hMxS7M7B49SOj
FgZL3bLhXxZw+quSWEOE2lknLhEPo/Iea0VbI25WVoBh23aJ0Lw2nqu5opmjamt/
7fMdjw5c1UwHixpoHdSqnOMcAesCGx78GFLXXYZ4aCgWzs6D54LyF+mNQEiiLsVc
ZTVqohWr6mX/JwgsG0zn5kYB/ckkLyRjWDLhlrR0Lc2R0hkc7ipgl//XU0fpbQbx
AG+SNC4aenV5U6rHwPpr9s0INhxzCW9oeUwRyDNJ+gAWJj4PJRNMbpQYpPpKzl03
Efck9NF8yeUyjHjhWaJCUMAT2EPvy0V92pY7rhmBknDV1ssRHGE8VozG/s73fhrO
jRpPIzMCTAXiccPXEM4wwOdhIxa/frWdu7jTwkTgVjSm255G0GoDZgIruxt60yAD
biNtmI7JCG+zPDJGzi8yExvar9EgOIROBbAOONaV8AcH98JwFw1v5WJi85G4WEFw
tm1Fa6jydw172JidbxH23X0IYZ6jASHV3Q8aC9yw6BdFL1inIdF/qTq9yI9Mk2Gf
FNvfq23UQVHbYqWH0bQT4AK0FQEhE68QCdirkDhoTDBDX1Rs7IazTGqNIzKeA4cC
3qbelIa9fY72kVu8opV6JEArcIZIZjPY0Xu2Mv9Mbv103gP7v4FTc1Zwj8WN6jDM
GLI007fQZfqVJri8lVwkDe9azmY7GBUeSEoTq0XHkXDDYoEorkpoPccwUUhsV06U
PUdYO2uyQThw8qURZ8khKOfoE/gwgoKfa+EQS3f+2+HFj+Zx8wulGz8OTYBfjfX/
ZOo+jqrV09LP5iKtiKdKJIHkUEPQ4yo7VDdHc7kAEPNE4kTAPT0H53GHsekjF9oz
pw6N6BFkVBc08eSLiMB7YvPlkngIKoOj2Mbvum8x5w+5OMCH1O5Nct6GoVMbSGQA
eDAlHV/i7Wscg0pvIVLySBeI7Uh97mTqrhFZn5qYSE2nh8q/rGVhFHZbneqDS3VU
ZxTfrpM2LG2P7cPAmJw8BwGMYHc1f7wZkIkSJTb61Z3/IvnNjJ1yWckvgKPFD6zq
iq5DFGN04DYlEFz+Soxchc2g/dycmpki7xWWpWcrEnSXySBUa5J3/YG0Z/L8GzY2
CiMxHNq0HenLCjXvqrnpnG5DCp+myjK8/FedsW8FsGm1Zupqt5dNtRLU3uIDCNJ5
glfo5SDFfNaBhoYed7ApVcmB/Uy0FPLFw4rSBm2kBc79o7MbAS2Bopdu9GUJ4J3n
ZOXUfsM12ViRDd4hRzdrsRMctHVHVs6nA61OjNIT/hjBHVIot0Mmg7o6GwGzHnyj
jO0CHaNaA4v/9IToPd4P2PMfs+wPK12EhzKc5rXg/Dm6seg+J/6kkHfKNeKtpeco
UW2SdZKcvx4AQcgIYZjcPWyKFS+nkPjfeggLragnDK2PPUwir8YVLd0qiK7zBZ1+
xMkYLDq8PdeRonm4MdY9kv2J/nR9Jz4ISDkXyq1tY8mduAkM8OBV8mxbilc2qwHP
ccpd1c5zNq0S+0AVqGSbzX2oonr8DxWv3sts456g23vNlv+l4e2lCP8RXmfym3MF
M9oodLSC07Mfr1NLP3KbzlM5sdcYOXPxoAhTlFIqfqKuzr+IcPWdoR4YVEWGVm1+
z7fKKOc5cXub3OLOrYtwBRHQYS6f1aFKhBZ52qhDs5AB18cZRcjrXhkXbq3nGeMP
Phy4wXeaJiy18WM3pEpIPvmw61c8HRISSUqe5iBFX4LD4CxoxB/2fXzep1SWzJjE
GnhPEJp+MEVOwx6YC9KuqPLlOup0Eoj4ygmxEzBqK7Vhpb34KjVaiEKNDzfLEUTc
ltY8iel2sKHogzddw25OxqKa+d0HvQz8dfS49D0Bl/gYT/V5xvpiJ77KwMN93Sc3
aXv/6H9FORP4Uc+OYNHWVTfqdHlHpIvyvK2DQFDRmmUNRoXDeK6QkPaW5PX/nPJk
v/570dNMZ2Zu8NxsUw70W2wQ3FdhP5eENUH27DG2n+8cnBo3xVCH6BWyxMxS4Zzi
+lQDmn2Uvyn6nejXO7PBky4QD1U30UurBwmxZgpr/0aKZxG6ea0OpR+SJtY2A4AQ
IJ/BEsYUyxV3Wt7Qv6fJ/G4zxVFGaS8c8HjLcpCnHXOv/ORyQJPi+VgbAEcng/ZT
o1z6770n4SLac+e7eYoXfRZOIE5vHvovNjk5yRORbyKh90P2NzqWL+n9TlpITY3q
acwmin6mB64L60Qm0NIBm6BqOGxzdx/HZKmuLaFM5y+eMUhv2mNXGMcUMIZo2ny3
0eoteJazSNhykH0uH3mjiwn3NE2FzwWGEuHBVQ9OIX5b06WpRxbYpGK/0qL0y5dQ
B+CL7RLf+CKzAJSQxaC2RxXJMioodd7PNBvyCQX0DlNBXEmg8/eBEOfbpBlRgdNg
Ar0GbEH1OujOql27CpkWnPF5jhLrOQALm8gwATAotSiMAkltUqiJSe+46oidY0LT
TKopaGGm9bMUYDnFfEVNVmzt2ZXSJjE2ep8/4bonNoU52bZnRj96dnM3WfzS6GRU
+48+rnL4TYpzxoNRTe8aZGmqMq9BdgwEJysnK7bCTi2Fq+HvDzYSX0pFwYkR/RxE
msLX9PzqT2SCRuwrqBXdq7DosZZIgLsk+JyY8AuIdBw2/iusJBY0eGbw9mQIvgdD
qzYAbjt+tdOJjZuKxBmYwQrf3ISLdGoTEOOmIYqSEmMOS1iFSVdi3AsN/+gFgG96
HiH2+qNMp1PRRDFZwH1veryy1BVVRpBI69fmOy07el+YZTUN5g7O9j3UKUfWnhoo
KHxAPudDv/kCI6hc94teBoTV37PKS3lJgS7Q0QVaR9a3ix/GSaHKzXu0itCPZLoQ
/GVUw8c0u+kr0l6fUDTOBHgG17Ys0szOY4CjwBsVeDKMw0EDEfXB4b1maMID4XGA
4DEEAwR+f8mS8qmG/YuHpjxGA/N6q1gQFLc/qnWWpl0SLmSPM5hV9/ihwuvKW98Y
UuT14RkKatTdANOHVf+KYxyaSRbJyqCZI95a2HeHcKPSvG7qkVjOlPsfseOcZM3V
NPKZi6ROYVcYO8yEqIWuTPzBuI/S7kiinzxAMLEVokKVt/reXJPwEX1JzXiVTXtn
wZ4DPZcpYBG6iSNzZuNFe1VajWGu5UhZkQzJBsKl/YgUnFY79Wl9OG9npwigcmB/
d2tBb9/9ddkBwn6ZJioIXa09z5QoVCYHTs7Sxxuaa0swR4516nEGYhfQ7dGz2Wa2
upB5AXofaR/jvRNqgZofI7KE5Qs6k0PkmZ7sbm5jUDzwQ268ur0MyHbjnUhOORez
sJtNRVkJy6ezWnAp2rsvcLZGmcVRO10P1/pJ8t0J8tC97rXQ3OcN66QZ+LVumNdK
noSqcua+gvDqi/eVWBe58Bht4ogM9/VSCjqklZuLR2SytBnPQuqZKB/dgUjexOC/
JhHxMoIwypx2SoeAnrf8azCpXM9pQ2H6F4uqVk+qEvatODZpg/EH0XUgHjizEoPv
Tvs2lXzIvuSikgwnRvAft6vIGjm37ydG0PSSK6BTDL8n4AWkRHD0xEP/gsXBMomo
Px6NXZuXDamRZiJJcG+0eu/cpvtBb6Qko3IqUkOZbPgd0FUVSMARAVT4vJqUmH31
IDrzresft/Ty3CLrrzX+yzGnrlysRQGrj40nsE5ZKlZPl/qmh7LHoJulltFeFJfG
xy3G525LeEXX2aUyEcw3184zPgO8DRXSKylD/u5oTI/ZWRelAC2d/qReIhy9YZ1Z
pyr0IyZqpZoqNdYBJq6ZlfoBs3ObQ08/Uxczxoj1Hc1XNKg8xVw8XfGVpSA7HtJF
YKGpXoR2SAYY4DRYdehxpqFqA5/vB5xLzQ5eZpzCxiAZd1kh/6F2YoP7TKO303HY
i9OJBQrDgw3SqnyCo1aq2fi5hHau1hIB4jjpq+hBJDsxthLC6576rToDJ518VemP
sc16uT2NXHiNp3xV79Kmm2Wsrs3S+ywugtJlkA0xXN3LfeYsSpdHklneCRgKhdR4
tK1QSjZD2EgS7DNDq7kohmHEQc6IhG2S8gwmrypRhzRPTgEsY11Dh4nAbu4nhgWf
kjNGgzNVWAVHmWHJAG6J7TeN1Xst0A3I4W84qh1uLf13cCtd/i6y+AR3x5d4Kmd8
W6vem+WpbWFDD+/KJex8+lGMNfU3gprVb1iWMplXbBlURuN+931Ujq1HUHmyKLDf
vIbYo7KZqAuBW0XVq8rotIUssgcQmLs3mca5JqEdRXFGm4tn61IupK6duikD//Ho
Xcz4f9gsemhGKoobcEp9gCTidlpjzG4L19r+AiPGgb9WSIZDAB3Fgb+ADP1CmV8s
HS3ItkHeKpfw6KkFFqb7zJKXkg7fElYqNvuoWd7YJkwpBbAEzHf2i/K7j0kXPHub
MGcq0ww9jSH+B8l+r5XRy3v4UdbWViGDUfR8JZt01CRe4JcJUtnSRnwyiBdY1LoG
2o0593oXBLu0B89msGhSi+jhajYf6kCxB8fM17pAxyGgViy55ni1No9bNq60GJbB
VxHxX4h7qHAr409ZavyQXsalv/AcEGVDbl7D77ERKcAHWWpK6IqcXuM62FAlzUxF
WNDHl11uZyr9bJ3jtJEap8YLP+0ppt+5DhedN+GIymLaKTYmR1jpb8vHaR6/Bg9e
+gijyn+7aXKFbiuIZB2wOB9oG8oG9T2T8BVJ4SYiTzrmpYrEITO/trWiP0tH+a+V
KqyxO9m692GpUxvacYL8km4p/AAayygbPszvE4i4WkD/DYxrrOjPi/lBz68YptKP
tUGbN0fLrN2Yeqay8lYKnjqa8Rqn8oAcaa0L6+/S2/VBXGimLAVgrtYsESeUIHzT
EMLSHWCZAaBsRLxZlqT66DPFoIgwf7OQUZlz9iocCMRy5FtZ56rvNVRx8j6bgrr6
9kyxYqG8ddpo8/8k4uQUHZIsdhZEIEtuAOukNR37o8XO69tczQUcXpZyrn8zrQ77
yfvrWouxTdjhkgOOgpsnoLJDhakpAB2if0UZwdB+0Xbg4TZry/AFAAx82/F0yUK9
R8OAnV3Wq8/x7zV5+Jg/+78+LxE/4Pmp5c8SiW5JTmyGy56sm4/7zBYXCORTv8E1
6aS4LLkUz+0zFrvYzUzZHcOvpnsLutzUwd+PT/dx7pSX9f0Cmc3JANYJNOSkUNn3
orl+ufF2Bp4+ALfXxltEemoFKSQolPf+d+sBpDAaIJIeOypPvN7aeuAfx5VzTHEW
CDTMMUvcgS6MuKf4ZxY3A7mJGOPuPENpf+YgQATMZ73gStleVBQCyXtua+rVr3iV
YKLXNGTIKWZL3KSY1jRANGIIulE2X1OBj5AB+NzelrhfIZBIN/eZGFxPALBUWbXo
xP/WLu8/gRMiMrCuYbnGLDF43XR/rnvX0jfj8aDqT8n3rAKSeoUAZw4APRJkXj8k
mDauBvz4R5KDqkYU2WDQj1ZZ9CdGlcYjieCpBOjWVbIruuMe4814cDPxmlR2hQ//
zhNad+HszTGI5bHhTpo2taazb+koOIlW0rDmvyKqBsoeUChXcEGXo77I4cDcyXuB
1Kw9eO8IesNWHXZGsluTWo41lJKr7tIBiby1nkTk3jz4dhw205akkrkfBBLT+z7r
iw4w7gKlI4bAr1BIN63/IX+o2YfYXQ+ZgRqg2m7X+N/uN8qGRATpuqYYQGPgKGZ4
lnVW1dL9hHVpUGoW/QYSeLBAV8qZ1UQ6qZhk/bvVvxp5hoM6wICO95y8rWI1dXR6
KxH2HsrD2ERZTuzqp5JL37Zrf3nln8S50z3TO/M0P8gvj4zz/LQDpIWQow77uMRR
iIBxc/b7n+P5m41W5szzBcX5nOXVtFEAVSXuMeYtj2ZaX88KUEKZdcx3yLmTCIlC
7QymX69ofLBFPIDYAfP7F48njd+o7KweCVD2lQFjcrM2/0ovKrxBSEJ2AELr7Dam
k+lkbYO4LuGHFtCdcr5l4JamxjKd7pW1++T8IObqqkzepCuuDIMc110Byx8JAZQL
RhsMwPC/CYCYBlgCbDz+c9X9nU+xWou+m+dgVvzdpnDce7GV0XRrTafsqs37CHxo
sYGkbA1USNT9kxyGNpgy9Qn332/mPXf+U1ZmTiAg/FHFvN86TvejKyddieX6wwy8
XinTdIlVbTkr1Vb9bwUTFyV9X9uggD5NlcI0r5nMkIR7s5XxThzB23XszxYERC/w
lVbx40Ueyb8jbzJYQh0P7HXuQ9HLxBRr9wBWVZz1d3P8BxcH8K0B8XMbnvhSKVuN
6HzjTT6EuR7s0+A5Ah78ojnBKZ1OAQkIB0ohD9vAPZJlolpF2O6sMEJiF0zYrgBQ
KiwHfbQuAWLorwCmgWL/fHgctR/6KYYXqFIUTonvUB3FHihPcWAFoq5Srr4gZaEj
qJB9SyT0fI7vjCSJqIBPa77GIGbN33DAZQ9WNxdPQwc/sFvliGXrwMPw6Rmi+Dg2
+Ub4tyVXCxVQUyR6GaR9BQq5gbMUOdlkFtMIl/6suYI7R2LbnlOc/t1U8neb6hKU
FYzKgTHQ/xP939k2bKvdV8q6vnsetyPZH+fn007odGMdDeNeNdwVPEFsUxDh3T0X
g1zMS4iMdgpN3QSE++8KwbgfLCISD10da5YjSPI/2miYWTsrIWFNnm7D8mSW4gph
+snykHix24UqW9AokpOkfIFJvEpDKpdpiOQURYVo80tLv+LO5xBAohkpkcwcLs10
gEhOA8tIuQsr9vYQ4zv2WQiKHEH1rBo9RP76GWjCR8tsDA+QKm52jCZS9VQZMf7E
EsvJxkjk69nDOw7nnQi8tFpixRs+KpC6ejMTg9e93XA9oBxzWLibPNPd4BUNHncc
qBuUZFHHh7ZBGqnx2GhU+bVEkkM2X3wzrJ3g0YMzXI5LfzppH589U0zbTjPV0UH7
xXKZzGLWvmlxWmfniP/S6xwipruQs60+vjGKg8Qbvm/DjlL3EPXqXbo+meYCgFyx
ADBzfG8QzUE7PWO+WuWfpsZleEd2mAIUxpemiqp5rgJnJ9i3KpYjoaFDMIPoPMl7
bk4tB3bKLjhS6y1JY2L3dCkR7cVQWjP2IOCFz2S+yEVXWqstYEKyGc3LXEi3PQIQ
/ggEPeEw05TRGOev/wBDJQCLVzdAxEruAfxIZ+Q7gLm5FNtKgPOdcAphvBCSZtwN
fGfxqn/vmX/mFHxGvHGtEvGRSYb5rLEc9nZYAM5v+oiFBbz1mf8VuCS2KVyqfilp
qPBR1ztfcs0HiHHkm2HUx11e3hU9SYEbfm0j2lKxE0V/aNvMM8cDbX5EM5Ow/lwY
om5VyeOiEBlZA+xTQw2+kK8d+W+N87V7ZaqZLQg7v/Aypyg8Y0bPjxqnJcJgTxGL
7KUGIj71kUOGHM7j7g2kAxZH3RwtCkOED/aG1a042+fsTwHhBtoLXAlWfSH90zsj
FtO+/2EZsZ7x46xdYJidaA+PO/lLV54BgsHGYA6lrj5BDu9T8irASnDIpVb+uYrt
Xr89uXIxmoYJW7HfjnJ+1+L0BEqk/D27A65kq5Im+Od9K0B/w9x5qCOOU0+GyWU8
PSz6fvRv/TOpgFcPyEoq4oGGg/kNwuQUvJK96Q/GO4jnTbw6O0Il4NWmQi5+QTP3
PMHItmRIJORPoHrU4nrEigMfxbs2hFdgd1ED7tISXHMFLilcOKGcbZDVm9dNWdLo
afzNZN1oyoXvz/Wg+XOk/n1qb8ndGw5cE3YYvR6pnHrfwe/Ktx9dOohJA5abFzGh
dZ6C7JHKyjLTF18bMt/jmG/6AK/5WiNJv6+r/Apcr6fICUIwlPBfsCj2hTjRZrM6
yPAPk+9Vt7Gq7toUzF6tDuUmuM3EdpYShZYAPBi7lipi6zVlsW6mAiosMihZRtLf
2gBM8UGqW9FCoc1xJAC8xW9GLAwoMTStnDZDtGI8EJjMb/+ov/pPiKlZKdDYHdOb
U/DHLxJioXplVKBi7scT0S9sQiYd4evYmZiHm6pLYfVkYFmPtM7sAk/61SN0G5bo
HjWlqhMLuO9Sri1FNfMsC/T6jCD2VjA41NM/uQP5fCehXoxreWRg3pWZbyxoYRfl
bNxokblVpcsVCQ1/w1A0G1OkQ0ZGTO46LFz0NHMWnNakNz3sWNdszDEQxsGNyCw0
SHPvALL+YCgUhWKXLiWqXEEHZyM2Fxa96XBzknzm6G26yz/LqisBzLn4Wfs+n8QT
TBADa2ezUebNvSxyUG63hRq1GGfUyGxcLFB+d99PK3DFkJRj67J/TL/bk8LiryWK
JASqDxMq2GY0J31q/UpV3NyY3YSjrUp/Zn/LyRcNgsDW7D7v9c9pmf7ygzwErN3J
VmeAOI7/ADeIQTC2bSdk0yGcyLTEtcz66bRKcnvaCLyilv+T/mnas5mDgoksWZsG
KXnKTE6QX4n5Dl+dF8lVok9thSqLyfjz6hyL4PjPs4f6S3XS4juHq7Bm1AfkdeXy
IwYOTQqXNrhSdGj1jPqIy5VDyoX6sR0rrBHq0D8f8GapE9B0+ppAXduV+ZREbeaK
kFuI+v7mLAdRmD76rfGPU19WV6Q/nPILQtaHRUieXl0r0nYjqYviBrJTrotyl2Hb
2IbiHlkBLG8nvXZUt2xviKVYZk1bMMvbEPBqP5gx4jfCk1uxnCdOTOGN2KLXMneI
yNH6IDi5fqptaqqLzbjdiczp/R4slFs37rdPqbff5JYZZnswiVTumSTY3U+3gc69
cq+UFtcgdLqPGZt4Utz67IeSs5xxY4wqogeYNTD3u/KlLEdjpmotLzeEQVy9rFs7
YlRpqi8F/hTiHNRpQDbJ6GpJYwVnM86IGLCh4tQrv/LigFOgykWR0VibHW/WhnzJ
lF1JoJw0XN1h0tKXcmwCpOjDaEuc82G/woGfETdn6KGmrjvzprQC8AYzjGawu3O3
9r5XRFxo3VqmRJLYRakTg1Djo8IcMvVqT38IDB4bTZfGSvfhX/OB79V8Acf/8IM8
ERpkifQdDe2zNv8ZXSFiX99XgGxkMwI7/iJ/CvtfpNCsPyOHs0GZzRaUQlef+VA9
/nQwd/YqDmGZRCsND9uSdYFdo87toqV2tt07R2fqJtP7FR4u6QLoslsWvokppmCM
GrnOHUsLcSt7OPdsdUp5a2geUZXRi8NjkyDtV/h1oHG061KEPNQ0Cu1eHAiDg7GU
IaoqaaR2DmUXmNZB8gUIEIm7gfscXDwpC+d+B+FUkX4gbKc+TclFDy4sD/hm70gg
/h2wP2ZCkX0Pf4/AsfHv95t18+U4WMRXFnFNI+aYZJk+ORsK5Ad/lqD8il/IHJVf
as7wcvouV7HV52kDDjIGpKETRUfxkADmaxkSltldMYyP1LQPLMoWTCOBrbz3qBjO
REYzJgrFN3SoE/VyPcE23tMe37JhL9e243yscNbRrFmm82A31lRx3UsaR+ydWrNy
ZmRzIBFUAqTLOUod4qKrUfndmNB+KacHsXhG3mG6sjnPFtB08GdA04Fv9kWYp8Ut
+hdszXKOK/PYeEwhuoYB7VnmdOMRmZ41MkVO3g5IUBptiSeUC7JzL6LGkakpKcxo
HMXSz3svr2A1OZrdzF5ObKJ5d5AJggGxUDShrXiB6dqKRoq1/C0kENBvNOawfXNM
kZ+D1OxAt4PrABOM61nCUtiQWhSNQXXP8gt5Wkv+qlNJY3HNcsq2/xz8kFmycG5j
j+TZapLApuGt1ZJn0vNE+Z4jLMumqxgD805xquUknR9+8nxiUOHYQroSI0ze6ie7
t2GfxZXsuGLEUYA0wGXHmoNTIWLEnBMWWi38ublT5ITJomv3abhVhaCAlbOnuG0B
xNs0lMyaVPvj+ysy9nr2fi1JZi2INaSmAbIRvqgCj0gIJaeVSNz1SrlMPOC0TKrw
6mUDlC/murnh0kZWhEkC2XZLdpbbL83WzkS/JWauM0xZqMjpe3WZn2eApdZU7BaE
OmNR5FOd3tsqmnz9MD9Eg6133Zmes9S+lEukP49u/q1sB3sYTBHTmAWD4DiyhkVu
kny+rtvOew9aAmAqM6vhSb5d/hFiSIQpaNFnV1H+T57LdfGByHb/6gBjf0iaof6e
3pS7agKu5TQHQxhKJCLw/9gxfkSjkAnR+xJUhNlyXybNKxudIbgrkYxlFM0+OJfI
1j526bfpxkEGLDCh/8wmK/g7mU1y0d0y4QATl/8ncoXnTXUUf8Rb4Ry8be1B5bE/
wM3OmqUPpR05Nxa/LVVPh3EYAEwGuuoPFaJWw3JaAgDLsBaWjJQS3lJDxLT9TeXa
vuRJgzfE6kD3jtI9pPe2CnI0+hYHCWU4svd8d0xp4GiWw9i+5nPE/je53nX24Tnp
/IYfmk60A+5/MSniUB2qBIKomsztUAo/lXv0TqMakTv2PMZBRKyfKVDeJttg1xoY
JBjRGAT+SBcuy96eRy9XncoTZ0Z1zkzRfj6fbQwx0IWrtkZewhvUokgPA3O0i7k3
wHF+H8BLhomRzBwGuBJV70GqtnQugqE94mj1hDNjXaQcOisRQt+siQ/BFSIK2GIE
+NsclLjURQZicJ5J7QRFrWNGNMb8xuPlqqzSnzSGVm8YJjioz9xo598KUc8LvFhT
GewsbpT2y/c9PIbp6p1TnM0eVzeiloBeWhJtlMY1O+Onwgz0KVTAHaV/1nBTMa3E
jsuOchlk8WAH/EfbVIaFKxpyWdMgXo+tQe1+oQTzNs/4mxjjx63obSOnNZHBtk1H
euuYVhf19oW+Rh9K/aFW/6ctSw1PV4K1lP+/N7kiuJIOpRcVyawWIawii++Wsx3p
Weyu0pkBHm0JE4xxLm+Te4VipjOKzu0Sjh0rOD0f3/vHrV6PGbwMBUjLlAgEY2EK
nbJjSqauvkEWXA7tPpQBVuRrs3WpPAoNjfChxA/ODjfEuef5hpiUITv4h9hFwL1H
5vThN0+bOqQk0SGaCi5jmXIo9aIuJ/Cv+wuFzYbiSEqpdXhWadECjyAJu1wPpFQI
IKepyX2F2kxK0K6isIhw+FENSfHbQcKDIlNBVmw7yGDx0fYM9e5f8UHp1pv+aKbu
wjQQYAodtKHgziYCrnjTK4nUrdDb/tcX2O9urnD4hBYRKRlELni3YzczYmL3CL/T
9vMxUNp8ee9GITmpaSNpNYT1OTo5vo7Sf4YEwOhWF8aY3SIW89P6T5n0CeSdL4hp
FDhdjmTcFLb6MecJxTHwUKGk5wQLsXkVWD2I78uiVjWnPcc0xlfsZjj7Se5dkYUk
nV+clnqir30NPTwxhsELm0bIcnRaZ/Svw6sA1gm6Gda6Oaez0jrsZ2VsgiB0u8j0
g9GFsp4sL/SJ1pBq7GR0E43IN3Aw2oR4AvS25TWed7hfh7CKljenSEz6tVIGYCDk
R1sI4ThgaAgynZbMzGOi9uRGWgVSiBxQIA8NB1OJnQvPCyqFLiRQR0P/nPe0rmKB
xfYXUb2PkWAKplx4qKKFUzYtuSV71z50O8ZcS3yuz3fhcNvx3F+32EGPkqUcrX18
gkHEjP2bnTb3s6BrRvCRiLIbYc9phOEtoAFnTQG8FzVDJKhYccRHo9OP6OMFQzq/
j7tVu964rFAtNwVCR3cTkaIBUmOxDyjAlb3NTgsy7nwnvpRJJkmGau4fQ+NmoDuh
z25PbTQbpgiQRCllK7WwKrHdpQC+4oC772s+OlkPegZYfLPR3j2FwRgfTljgzfaZ
o8WTrr13S4ua/XY1IAFUUZImvZwnsIsNgcwHGh3eSd4efbVsbTC7DN6phGfx850p
hSgD/wGBKfpuBQ/g/RowiepvRpkjGELeVGVm/PLGr7FY26dZq9R2VEWTo9ldzLE4
MUPou0WhtCV2W4ZsWvexQcy3qiBMbdrePsyZZ+5u+RNHxh+KK/LJvVG0Ka6ajAfb
XEuJO3IqSrFC/V5EVDSSHBtqU2rlQVyCmSCk7GwkeUwzEny55RCGgBCc4d33zGUr
9RWWi7V/0zDRPyyAYt29Z2ndJmO3W3stqhqXosFMe9Zc+V/c/owUpQrKxG+Q5ooS
fr/waV7t3Bes+bAk0DtvUWTLkUKkvp5507k1fE0cHQZajGB2oO8nj+z1qyk0MQ94
cDdzoTjNfnXJ3mW+EF53d3SIxrKLZdyVgBxUFbAqP1hUpFpQD6nINKuDGkDu0wTb
1xiz/8OQx6BZv+1bKmVtj1UB+vOv23M5dUWW6f9ajRjAHNYyMpAOJdvdzlJ0+3Re
cqGEZPeS0+7qWVY5IgtdPv0hyfDCpruYLKURw0Rll4C/+Y646I6RIQuv5/Mc+OTe
E/IOuvpxMc+7srIr6EK2O5jUjRWlRKUFCtPvkdwukCIEXQO1q/C4xBRs1MbXJ3/y
lWWGy6frAZ9ZN8XFKqRRiXKfvGYwScIxNM9ut8cHYM1IB8+lgScKow6h6IXXlc1o
7fJBEBxn5jGX1mvhOOQn2ED5vvxw6sV4JhWSiejmzTEYNQ1VRtTRCfZzNJ42EyU0
Wj9pxev6471D9Rra+HDPX70XJagWimKHLgdapiiGUcolMLfkREjBBjJn7jtJf8yW
TlF3xCX/Cq3fiMkHogvUGvhtJiHB2z3vOCo6Xfxa5NNDinL4uEMGnPWG6KXJ0scb
PNiP3XgRAHxDOJjGRAdmw3sBjh0JjCful7pvHwFSyDUyQeIZdQDgqZbEiWxSogaB
aJjd5mzmzhXMG6InUcu/hclBYytoYWGbeZvaG+OmrdDOZDAGOXkIitNr9hVXYXpv
ARlIo+0jYJEvPO9CjOuFOAxdbOBNrK596yYPzshzHLTJs9bXV7uLr0/2egJ+DDrl
MUaJ99KlZghQc/3KxxywZmr19S9fHliTrcTgW7bMftEgaixDm+oWhOcpX08BiQl+
YcMJGTLJ0OCbMIWbTa7IZVYpaXf2jOJ07UzHkAV613/v6NfREzGUEarJvcLTfCJk
pl7lzELs5PYuzlD5OJJ7ey+5bCJxPgI4OwgDTAeYgHvKdN3jLO/I7ipE5Z5GcB85
LPOWAX5SNkTRYR3zQDqqc94NKSwKscjg7KpRhQFp9dBnGCypNEPKSiH3sgH8mL/Y
HgK6Hxyl+k9/vdDB5wBBFpHF9UtakZiZ2GVieXZ53vfNJMXtMntlpc7fmWggXV8h
FzhOoI97/xdsYEcXcbFWuxZYv25G8izkInhuufMvb8iZrrBkLSqL3A4KE0Ny0l8S
qQvYqFtlMI5CHiKsr83M41kXTC8n51JveWpCW9uEhJ6NrhQf5WrPYI9Kl1AjKOzJ
42YTZWpRml24YF7R47fgaQ1RzftgSfpgaj8JJCcxsNxnpBQOqM/6X3Spyg+rJkgs
PyyNnbme4mckbSHPKYjxYKOGCW/mn8NMD8yC5ogdhxvZ/XCjhzJRbUivASQDymMa
JKPd/QR/E1g4qtqM2GkK4wwI0AYaajU8zU+/omRnVRw0CQ++fHfO0zA6dKFr6O25
unZ6SPg2R+90A/hhbW18KPrLDByUEfy/iLx4ZcfZFLt6mfdieoZ8IahaBSFwLvh/
gBszDROMDqNJR4QCJ7uKRfGieIVvb93vmyh6Xn3BAjvmE5su1opcAECGFoxwDxpa
5ahNbpXYXKkIBRvtTpPKyT4S3I/bker09Z5YD8PUNFDgvNBsxWorF9YmiwWQXrHE
QONr7go6qk5WxT/HGgdD/1ayMK5GlxWEdQMKwyTDQGCkfBjL1Pa3qvKHfHPzXZES
hEK8LkXn0o3XBH1Rd172X6GcaNuxjnwtESSbklzoaooj9dBUqWFKqFlyuZpu0oeS
1zbGAr1J/Jnz53OmtiFGw1/r2hliAYoZomYR2ocVpU8fAw71B+GCBqdg8kf84rcd
eu1y+2VhuwE5qLrFBnXUl/KhETjh0Jq2/p6hyXZIMB4Uk0mckrdCIeCEIR7Zwxqn
JoW9vkhHpW2IPGvy2ZUAEtBupn8YKgGA/pvZu93/3J0M8n10lQPxJUeHvOp2a474
sLv4NruB9O+RiNNvMAvtEp9TYI1KMwwuCn9APiMG97VBGDOsBnLW8yt/RP0WEgQZ
v7zsunit9Vbyq9aZG9/SAlDLaQFlir2p+B7CmwBauZ9I6TsqrkOMmAK3cZsMfYOM
wTUanmLO0vb1y4G99gWVA1FjzHhT2RzwUriTNIxrX8cMaBFJhOJH9mEWtIqdh1Z/
+WJ9sTZbUsFRoO7kABTONiefQwGlJGslwvWZprJhFbIlFOkgx7s1Ebf5ChaMtey/
VxrXQBjB4+sTDmJIFJLIpu4fMCFcipLG/nKDQc7koKVsYG8QFupeTSrIhH9yfg6Q
LuMR3+4GWzVMUatVsmiCrWaPVN4EI12eo54Sxjv1B4om2CwD/ThNzL4+4pF6HLRd
IinpI2YtLmd7MpUQQuiWUUcN8fUEUL4rCuoR7H0rUNkTLJBGNCtdGbazUDXCXAxC
K32l923uLERy9u/7kwEgYIMPLhjhdroRj24OloYqqNN00xwLXKIcIkXJnXazZLgT
sWokh2zb3sg0tlC2JfNVBKUf9gCvAWW9XLivgO01ZAhgOmMRjmEGUA8FUL9bHTrb
3lw5Jbl/WwuNqkI28XpMy1/XUDws+/ldkGIsRPxeZgNog85yzAoD8Ltrq3KUU6yQ
a1iGXgTktAXe8hbYiCkLvHRu6TWJs/LFAjyfi296oooJZLe47hy5Cr/O9th48nvZ
fs83w6kjFXTinB6QyXfi9+ICkef28OhMwpmTIPjyNXbFmXD/K/fhQEO7mOwz6w+3
6Ahs92AAHnaumiEkPef7zgUsd4eMLDs2s+idNrWU3rj+nUBux9x5kW1YQswAV4lK
6k1qSrPjAQ8ZRBoabolw3eboP9h8a5UKDdQIMsobkRFPHaQ+7RC2FyQCl+zt7Yyp
ieBh0uKzygRNYuuMOeo2DjVcuS10hzm7Ng/pqeJXxcPZ33sv3cABjnCD35VYSOAf
2cqlehcUMonnpI/QfwKgrcMRchWVw/QA4WkM0TKU23MczfxHxbDql/r+i4x4G6oE
qBZV+DuWA/R6AES4YoImDhkTZVOrLPHGFxPoV4ytRHlwhr9uLJc+LaHHhJhJ4Tsd
sDLBaIkakfxaYN1TaveeoEUcTHP8gq+MFo5OeW+v8x0zq2tLtXT3FOMA4Tg7kGct
B/Nl82DgR8wwwFHErgCTwFwCFFs6sm07JyzXP787vPus/lRi/0Y44zFclbTi7SDo
jFEqbsXyQ4WA5IgLgSol3Fpvlg+IIbCEA/deoBfa7bn31PUvngtcjEYBuIX7bxZo
m/a0mutBxcIP1L2pnEXH3eX/ei1CpWpt32T/0kJkhEM0KyBwi45xM9dErWzp3nK4
YnBEKQNwwWoQMNG8GRD6TMxWDWd8Qa+kkfW6g2HYA9oEFlR9mFe44g+FA12him9z
Z+0WtGxDjyJVEoYosYIHnH8xbLwj7JlL7TGCKbFJVNp/vMvx+obfd6XuWw+baI0r
k1vGl+1eIm6AFlUM/awYvwub6YOjC44us7S6mjKbfgspbXCkrj/lQLYOXyfoAeAc
uMoGlVFqAHEQDVidaav2yuLXE20bos0eZjoH8Mcg2PQqzEBnZYBjQh6uYwO9jdUy
i2t9K/WH0jzhM7W6D6KNvMSt3Hn1oDuF40Mx5rOYpkf2IGdXjBrGYjnHepnjj3H9
2q7rcBNWeNyOF0CVUoieI0N/TqHXW1yrARFhardOkWlB9wg2BRa+vBu3EeYf+5J9
uFoB4j3Cj1B3NRDyT/fkIE5zfXIAFyc0SmbymHKizw2lyUBsnQiatW5n3EUIu38K
HrrDBw8mlLEdJibAizlhe44ZVQ5WYPBO+IhXlT5qkoIlfIUG1o6WOkSzERuS+uxR
gcbhqmF6o9CWbFtbrol7bGwF3pq9xL7epsijbjkHkQdFSnZLstY2SsXxYzIS/URF
OFrtCKkqBshR2fVmVzMLqwvs8DRfGh0H/qt0Jma5wV4GmAz8RPqdUokupBdys+aP
9i/MNYHMWU6vN/osf8BCxeMG1CVTkXI8PMftse2Hs7qysmMspMbTQ8OjbO+WST2l
Gaf9a0lB71l36beq0DkaDphe7wHpD3jlMMY1t8e+seaHVGLYGmEJouWzlhm8Qi5F
dcOsUHjbosqE0ICIC0PpgnRGhD1dnSObVAmfEKJGdYJa63kW1zXnmIS29eEeR/qi
bK8eFkNR6B8Xz6l9p23od/RQGBKcKDhLsN9P7BMfyKqVrrcT0Dez95gJtKizbjNX
wZMCzEkHxJ1RU8wGjNMAI0Tum2YzrgIa7/2v3YinQCh4bPhuZgARJPdKz+AzsNY2
oVBDck+LtuGUnTRcotYW6NxTmHT8BtXBvay69sv3vPyTVom4HsmPOrAJmLtO84PE
bEzi7Wo8Y7aNBP3gKIC7n7eBt8WB+2K9XAGyZHMIcd50v0GPQvryAtVFKS1FYqHM
zKYOETsacwI06Ei35rHR7f8d8qE7QIs7fvHEp2L/QE9Xa/mOdBpjuQbVr+71Fo9Z
atrnB4O87p2gMx79vNSW6fwTQ7Nf0vbGwCZfe/+xgbsEQrQdCSMmMJCtAkEJ9yV4
xe0YWnJvkwgO4GPKIl0NSrK+MhG5g6OTKRuLAmAOZhyViLoU1p4D2lKvXfmtXOOw
eD6WDYUGbdAeqdDJIrLy3m0QseYkUOzoGg20ndCtJUTGjAyG4b79lRnZ4k5cVt/Y
uywWuZHFaJ/Zd2woYdO3kRyltBtxSuTIZOneArtgzUtfViRS8eGIK9ZeH7xDdgR2
3/S1+N6kiPVYlB3X6TsT9njKGfdhb0XqELVf2WFJNwIVW8rAHQCkxk3MjH0XflBf
i6mk0dcHh+UykUlVn19I6CNiNSbQN8qg6qHnKAk6XysILCAjKzp3ueAnxzElxG3r
IW6xJVwcz0gXVj2S9PqL2IhaTOeBt2O72+WddiYLuFdSat31ehTtdbuPnyKbh9+J
/dsm6vw+C/JmmZKfmtQiVenWOlED8zyqpvFx32a3xhhiNinnKK2pYuK5LSCFRohm
Cj6UiJZUbLYNHhylpO8bUSc8yHxSvftj47h+MwtpBQl9hTdpQOEOdvr8+chk8Y9k
R4rmj2iPxt2CxBfgc3GFh320qQT1ihWGDhuXWKOBZaXEDBnrHYtaniojv+anlekn
JjG18PzKqaWr8VJrBuvKrsTckvHskL7kpApmJuzN50M9Wfq5tUAymHTkPf83FC9x
j1XKiLN4FYqkIO2TZ5bHHCl7HVHPeL8aRJ/zAKmTkZY0AYxqize60KUWvD91TD4G
AWQdaZGuoYY6LFxtukpn0+qvBN5ozmMH5vUx96rGpeip9s7wCISd6/MRhs+sBaVJ
Pz0/1Se6PoFIn5eX81A4rGNJBSIDKLL9B1GswwL9TrBdId1juyFllvwpaR7dev6E
lvLfBo83K3ITN9CT/CKE6h46IcKCZxIXl/6loTNUBtsklD5XenefMFKSytgHf41j
MUWDCX2UGTZyMXVPTCclZEFAWdqcEbAap/jidbNOjW1mgU0K+gNtG0u8b5x72gjc
GubMkr8JkK25CAiLvOwPyKP+3aZgF/ADrB2t8XbM5fYxYwZ2t6QWu0PnS985ETGz
WClSg4igjOiD9PHp620+EdmdszYGeGvXCcRwJkhK7nMKFBuZBwkMBVTtg/tLSSV+
AYNhRdlflQ1Vp+11v4qc4qftEJYYUSEjPl6LPGREwfLSftCRbGHPGEox532NgW37
P2w0VP8l6F+RYHWJsOiQ9cpXokeTGKn5raCoAvWOL7cB5mB1JXqgehlzWXEOxt7A
pvRT8xKv6Ya+nXTBsbg3WxZPDWKgZ3yT2g2AThXwap7MwOSOHkjhS5RPUqAn0/+y
gGnsd8/jfaBKUNjABP0RLXri4B06ZXypSOE1mBmEj30inUgsJrJGncugWHOQ6qoW
kQv4MFfGSOprdCCGN4s1mNcA/Q4jGrcVVvapUPFASi8E3cQZkGpvXCsWGcBeaaZ1
GnAKPCdIqaTQGp5hW6R/ndtPZ4Zjq6dInjQIuocC1EBqIQPF83xK+DGJwQnEH4Ok
YrltWxJiPAzLvf/8Xd/RqWqIYJor0kPUUgmmNFmIsON92ZmY1KYwfQ0Pp2foV0ri
VOvI6cknV4higNe4gPOIez1NNqsVfb8pXtxZXSH8fswrudtbzX4W/2BPldOJGAzZ
gd1EjYbLWfj5Ku7yl2uVjqf9DIPzPkqqPocIUyBFRKXX9cxNbXnBRTsE1a+2H8OQ
Teu/IZLcolI4pgdpcC28AnLoSfZE5zFQ/jTjeBC9jBtKM6wZs1AXq5rc/HipZmY8
8uZls7TammlYqS6s3ndRCkkDG0QV19HNlFFBRn3N80ntZTYrcmTSTz/ehacYRQr7
De8SaVCbWIT8apVhdPd+0LAojqcKujfu74VnIBP0YHLAv6urWWVUKvF+Ff+OJ0dR
LSlh46x3qHoWO1htqauQySVoqQIzfKltFsl7uXgt79AGlQi7DCwXW7e82Xx6IN+F
DSAW6nx5Kum7B690xiX3TlK6vmUlpU8HUud1ScZ9zJ6ovoQwMzl3lS+iGsGmv/S7
YJkp79PSm0bmar4XTsVROO6GYcwlFPI5v3SEVUtDU7x0Gl4vofAHbg/q3R2HF+nr
LFaHXTYe9nKwEcV9Mw24IG5OIiRRxmad0Zm4wT3O7/KfjKq3yPLLEiNh2EED5LQG
n+TCMN4DY0zDZcv8FnevwlrZxl7EfjAR4eUL3k+4GuQ3kgaaRq56HaSJszycFWqV
hiVQrIyS29d4LwWbExhplcBORMvsA43Sm9mEjHy1igMDVpqycjYAAMa5JUlgOqIG
Ntl0aEsnOShWihBwdLdd4+Fi/pWiKp6NwSIrCzBnXjofmmfdJv5HeIeelCuXzFnG
9WXCGaisW+IpCskOyt7fZfB1VH/3CVbgs3XTHWRacOmMVyUoy9PtCLFAtQlrcpkU
WOoZvNbpWG7R9l5+rnnj8TC61crXiBhrYdznF//Kbl0BNeI9Q+NHR264lm9raIhg
E1MpN7JtGfws+1+j/dlEwd+MCXx3SOLSCNYbWcxuKMftgVhislL4HSVfFWBh5eU1
vLbvNlczA8rL5H6Czd7ySNcUFc+ghdTRv7m79Rne9HGaTs56vT8sg6EkV2tJ8h7Y
ooikB8JTnyCR8anRyWNo3yyopWxmBS+V4smwmthVpnqzqtjNtYq902q4xfiSFBxA
39/v4xvFhHyFYgE0RXvVzL/fTICSmgk4SsduWQoQL4CPayj5nKgnIxN25M/Ax0sG
n8H+7iu0swWvU2Ggxv02L1s7U1bLPOFEqmRp/GYKOnjcKW6EGUHrXnFLJlsQq81i
BaetjILZyoedftHrRnv4W/ONBSvEFfk9QkISyjwY7hUmczgKKLjsLc6xKgA8n8ja
dcCjR3mB+qHJCXrQFGGQJVTlvyh3IXjiMtSDUAY8mru8hfplLj+029hHr5n4YFa7
o87b293kezrOP1xNExXRsQTP7UCETG14bmK6fWkkwx8eYOpxubxFlJMJmq73JJBE
9CBSmIPMBbvIKxyA+29yYYtnjZptf5hHZAPhwk/ofRVKf7dKrEpREMtKHyBT6NI9
TpoS9fbvLth3lQNvDq9JM0o9LzGJdqt5b75QW2s78yAlw5g64fUvkqXggNguKOo2
AKgnlb4JviVwForwDnRwwVLNun/RKxnY0Irq/h+5/K6MoOygoLQozeOtwT4ucLLX
OfRkcQ0B2sL1oc1zTgNJnGvU/pzgHTWNdJMulzj3lqlWaOtMZ9bSXUFjt+o53WZ/
3asf+t5++JtiLd1zzKDj94RU38pGq+jsmUUc0ecCEHi2qTHAyRDaGpAn/HHNiGEo
HgWyHUV2r+x2zVQ/4DDHNVeTHPD+aWhgwzlHRRLQaR8UjHekfm6bXID16WypJThX
kAKxytGM+oEMirisl7ljyhfcehovIxZJSzYEnCfmdrUCzBNhol7MljFVBRpwvq3s
QGvmZY4aUp48irCrmIuXiSBfGHZMryU2PM9DUoLkw8UZG06uDZiTohqUdsPs8yXy
yWpdmPe6u0lWkwkXZ9SEL4t63Blw/XF1X4w/wFfEEEJrB/O2HdBzSAZNriJOpGF9
FtFqivyfSB91Og+5tWLuxG8FDucF0rVpqW0QjhuRXoVK0zPyw8oG+MSdGjiuW7oF
UgcP2e8qhctxpxflGulgSk1fLCjDGQcUhH/yEDvGVr4WC9Irsd+il7ZN395flZNL
C4QX49Cu+tQ9DEeVkIWqa6F3Fu26AgHcCC1URU2h/C8v8cRrZWtU3eY5rYsIifeh
rmYiCaa6idHnqFG1i7NfMO7K7qC7tc9LpIp1i8xW/llzRbUcbMl+0nNQkwM5rtlu
wq2d2ED43dw6MpezP5Beq6OlQRKo7B2c76o04agI7sIXi7+ZS5ErrNtxgSQDtmjY
DHmA8U7pW9HAuiskUpPSVc+beon/aJYsDeOCVMFxayEzcTRmIMGV6YhtScbfShWL
JosWehBfgyP/joz0rk0lAaEv0bMODZ5cqNMnsOp4uFBEDDg+4Qu3PLMPNPA9mKbe
J/vYMeCfFWIiGtil5oSsw6oMUaHKdGDI/6UikLS3Cg5kBn85TsdPoQABtAC8OVlE
2sWc+gtahwqVL2NYq7uV5eigHlcrpifC9s2XUG3nCyWt+tUFM0vypEXwYObVF2YF
cEWEKVyt4A3tWIMqZ4jF8RoxP5wtO4+Ip/sHjqkJ4qB4YArdbyNsaCjl9fCiTUAS
BN5c5tNPkbr4e6Bqe+gzUJliQO+hANUGfq4Hw31WGhV5KeVdFs5Gqi0YwW2CKtPp
FQP9B3teOQc4GR6QzIkLxogMkfy+PT10ojVCFuywjCyUSy1jsi15TmsTwPB6IrcR
abj0MWnWlQeA8D2UpkTQfX23/R1TZx+h/sSbzupWBfUXLMWdk5+5FFSGx4I7w+fa
iS2ExwnAfzg4BwgsJ21vwR8eFSBZ/iTx504ErCWJg6TBNesOAGYTOdhQbmBzQJHh
24Wm6obKJcgRV6qWNpain1sn1Fw8llf5vrRTCl1gqbhqbCUm7GAE+MuJur6l8ycx
P0WJYBzv69QM/8N6IYziOukRvvZqMhT40KV1lq7A2gviXRgVoukz2LQcehc6xp1d
FDBifTq/Xv4Cj7jWci3U03M8JZ/AHDhLtsIPIjWPLimuzj0zSWbKqExgC0FWlye1
1cq4RsIjJuij5JSBvflXTpM38+OSpI2lqTPKlQtpSyOlgDSgwk+HZvye2d7j+KTz
7LI9RLC+OZS0VrWZCjUqEPubn7DHAzOQ8cLE1hZi7HQD9rajIghBHEe3ZJiiFasZ
YM/wXqCIrVXG25XASV4LsLM7CRtWS2a0F31cqhrtDMMvg2x5vhl3sl11AaoSgyI1
UMzpnYz1XSbNvPOrD8z54CyIqPFfqhsRltJGdlEp2NrG027bCbU6i1VGaGw/79Os
Zom9KHMV5MLNsKDXej6yRsroxATSuZdpgJD3fTQfgGskwHrbOzshS0tDv27J2436
+mKT1wTeS7bxFp+AoQgqo7epNsoqyRswRs5y0nZXmCKqVgSDMSFcXI6rmVt8Tvt3
NA2VDGy7Xrhws2DR/lOnozYr6he6LYcumU3ZBt9r/RFcHC1wY5bwq8YihT+m4CTW
OX0clLII2suUZICy3K+WTOxGVY58bYyS/Tt9vcBQWF3FAWtiKfcUojyd+TFlY4aV
+AK1jxfEJOrOobwCnyhnp9rjGf83YCsZwRAzAW8PX4RaPNDPKKufHEaAMEqR5SMp
6tnvH0D86jmEV4uIMLk/4ViPMkixAWuDLgl2K989xT/e9zKSuDuP417Qo7HYO4Ev
60fBc8eLvyggkalm1lyKmnXCRm6MDa0Pq64jbjE5CvBA+NGoJdnMfNiWMOCAehH0
wwUynroZz5gE0EyNOPfnkPBzLbss32ZhOusVhgVjbeHnwam+45cAT6IzpghryJqS
jnvpdkQR8xn/UNP6b22en8zdrc6BtidoETGjrb8LLseiTVyfndP4J2ooLyi2KTE1
uDi/0fATPRfcS/t7n+clFM9mdZa/8PoiqCaXezMqiYPET60uctcYu06zjWCGdvai
DaO9SLWGtPavzfXi/Fo6cjOu4GHMnZau4KhFNsRvPbQiE0nK6JwjLJMdUh/LwvqM
gj2JpQqw814F1GE0bMSi5OttZeMlyX6CQiNdRUMxKEZSU5j36EZxEH2/P1CHHgcx
utwjUyFD0w/1ergxqein/Z5K/IlwXCI1JHYfXkGDaBhZpwGYCRBuJk07b5HpQpqP
OmAEoayzsvBbcXYA0hCTObHoHqzOPtb+UjzVsX0liM1iQUNMX4zVP8vx+IXvwVX5
+BtMGkzMxUQQQTW+8b3KpbWHIZ7EJ2DqL0Uxw2/CDdfVx97lBfIFY5+xrytOGQc1
euxvN/aA7u3J9NgNUjl/fWMTBL7Fxvty9cT51KOOAGcpo7kpu0AfdTqdf4+2P+st
9oK4Q2ZG0bsKR9UIvvvTiRQP2FdSgfE/aLTDLoQwC3hPjdJyWQ7CCjJwuarcHkRp
dVh/+IrYZNKH/LLrAvaH1KhyEf4/tc8+/UDHVKQr9Fo2/1BzDFh0+Q8vuYiQc2n7
zE4xtoHcVC89oPBYOnBM9efW9XGuTs1zf6wVW0104Fl2y3cr6/FyYHeOdd82SFCS
/c+oSjJe1/ybl7C5j7HbT1gkELYTBNuo2T9ws4lh/7goQnuh8+R95Gn0uYPRbqlc
8MehD572mR+8dCSj/coRtRAOX47dMCsVq+fjYIym6th5MjDSrpbUdcQvUAo0y9q7
cXx4LDqMDKZmvM1aMfUtAvr9A6pcJSWPoOppmiONUcBiWS54fW/VFP/UoHQn0tKH
d3vJjfI1jajoNgYh72Hj8wGSCT+Wc6O/lPgHfDX9g+cuoS6JA2X8lVoqBnd892jN
9IwXuaIIQ7RRDe/fLw+ZE0AZvIhEvVS6N/qq5FJgzWr5ZYN4SDphBVeMwx6qkhL6
tS5wuV0pzng+JBv+rs1ho45cgQyDL/ZqrtN8PeYaEmDJNWkMsPDhJuqHN28H+NuJ
39p1HW/1lWmc5pdwm7r7Mz3NGYvKdXfkKqGRKjzr5AUhbS4fHZODhrsiTk73vdYr
K/8GWN8tGshgOT4U/Yrg4NUH5Eyv68iCYy3hJmWVykZyoftNWpToLscH1oJZUTk/
pYnSvgsxGtDIaLN0o7QBYsPwzhvJXjblxqC4NooM50zLKlnow8+hFBZJNr+p3JH/
uygfk3En5krjC9MZ54P7SouTREdksrNtqHmwTL6QG5T6l33dfO7vrPmQIDTUgPmG
5OH7QY0F5RSRvZYK89ZOr/yMZYha/JKEZbZx5pJ4hyXPoqWxN1Q2KUQrgRMY4CBi
z8gBfqjGJNlRBwem+D4bacRr8ocsCl1gcFI196onNPYfOQDry4hxTtpHzkaCvFCd
+IZ5LTsK5TIAZhBMDaLMgEA7sNPkaQgTqKsJiaH/1OI7UwYyfHdAX0S9vGW0nmsG
al0FGsrI61K/zyyJeebDuGZnjUxwU5ij9LJTfOASlX7w/kHQgi940AMe5lZgMdTL
V8qZQpX/fvvKEF+iwhrDSIAnW2z1jLarAOqril03h5VHPkuO2i3BAR5pK7k+P4Do
cPIIkct72ygzhIhdSRo9pyLSoEAtL43sd/pgKbZFLuqz6zWEWXXF0d5oZANoLf4R
QT4wYTzaED4i4+fkRishnRMogxXEAGarEBmQw+IfxEiYOcnKH9ERjozywucjqK3j
b8p7wmwNBM754jALACdsCyYphmdcuOAU5KXLf5rqSuel3ViSz924LQ9L8kUDQGbU
fMftBchTQNDEjT9mkwga1DSOUAiPxzToXKef2TVI5g8RmXc/JxCYXEU+lxRtW1+0
1a4WBGZeACYI3c7sWByts/T6dCsmi/h8KLsEzdjg18QEgGrmYdvSGQWCYRharDUL
fnMksyKKKKAZJ4Lgp39yTO09KElcY0WYnFlZ+UTH+mqJtGMbqOe5JiJDtVPDtWZK
OHmbjUuewWi7WDtSOVt7ChOxKQAfy2uM9tUiQDijZlasmyVXDlvW9wTBYpaDU6vf
NYjatLuCUK78Dr5mIY4wY+iOgaVcIiNx9tbjZ9cUFHMBeA+dKohzwrduYwZUHlC5
sm06SyXb+A47QZg12+H91yXx81UQZyQAC+LJTRTqv3MFqMc3Y+B3v1o5iEN6BM4m
mWFP9Lv2RgFxy7XalCjGZGEUsulRtI5dKK+6jomLwvhed1WnASHJ4AGBc1iYDxO0
+6fEil4ytTQYfNxrgYnfcrz/BvZmJRFqKSbp2z+SJGi4D6ZD3rp/5lXl8pTQy2qT
G6pn+5ORyiSw5rkFkeueHYVDm0wHfAc5N9St5LAXclDuOWvbxckLoZ0+krQUxGUp
je2LZv5t7WTPB3dv9VBQyXYHnJ2TYAXsES+BDzaLrl6KV3IyE8lpqrdnMCVsuaiE
7MRzNdPXIxq4n3xixvRRaVVX1p3TZBwhfaHQ1DuwCbX6Zcp1Pp2PqdRs6p6TbDc4
Ws1+MVrQQ8KTbE470WSbj4K5wIsUC1S/Ty7VgJGUnAr9FqKVCLTtdIZxqEILy1sa
9Vzl81BGkajN2JrDCipBi+2xLkWBJl4H/NfEWIXsGImQGF/ysE1CdmV3XausM0xf
AOK/yo42F+bGTkUgL9L+N0/qG2VHeWJLxrTTZJz/U1cAFGn7ODVW8/wPItuKjHYE
PW/nJuRK+nO5nbHtJsWys33Bj6TiWO8H8ZyxDcAgfAv6zHyCSnaoX1k7S4okDngf
IH4dk+LdBpPpiRvs/3ShDXiKxWIZDWYvUv89ezDE31FeKJw8FJ2FY/OMmJBxBy+l
OKA1xpj1GiVjTuXFrE8ugFTiX/ycA6SF89V/LdPigDxonlfkQxysGzeeZoNgIwHv
BqJDmc0dM76Rwod2T23Rk4zOZSXoC97BYifDFVt5D17XR4Qg5LlZUyBCilKgxyq1
Y73BZcThnkJdQJb0lVfGFg3GAksgGwJo4d5OfIJ2P1a7XsiyJlPJSoacELyfsvN2
hXu5arTXpZ5kM+0+xKwqUzKXEfeObM8pYx7ehudz26+p46vAslmdsWFxkEnr/WM9
9Ti+BuSpQ0iXbeWWasnEiI/q7JEMN96Baa8KaxzglEawLIOFpM7s5td9BJyVGAbh
VuX1Df/zLlUx3vnd5kLAg7D1+4J9B+h4ZZGaJM+qu+8KJLLVMvEC/ZQrv1I8Tu/z
vbkK0E/zukXrcysaRw6/atbmXECj7XlEjxjCdsYimLkOcjUhvAlQphy0xhcsdnDm
H80oJpsCnRu/uGz76eSDqSLnf/3qsvoN9mKWQkq2uAG5k781u+C2/4/c0uHPqomu
SO0nHNLJOmE3Pri+vTCz+U9mKM3pxindlEAtHiSdDOxCy5dIo/BzsRfSIU6cu4jy
NbBXIvN5zS8oLPtaSyGXvt763HMoIfmm3X8410vI8Dup3UE2Fq6GyZ6w/fJA559w
2bxjKeQ4PgHixhLM1zJacCPPLXRRnTPTCz0+OZzmUxW23MJBJpSqnkyQaV5PPM/T
/5wc+6Es8/e2vP9kX3icdccucTIfMh9Agwdjz6tLcBqBRV+o9DHxg125DZXmalwo
q5oXQLUBrHsDLSE5mU+CTPDmAdv8JcSoYI24Qk8m66wOw+r3N0jyEWMK2d6gClHR
vWUz/I46hSwM1dZZV4+w+cYbvazNj8Mj4SGlERil10SU86jJW5JuId/tOP0Bw7Lh
Vb1mIloRyZ61riC6ghN+Em/fkPFvoxXMT9eqjRCardlaVAiBtVfOwYO93NRDVNNH
F2kYR2BprGrEKye/kLgDWgr5OuhU3DYAWgw5kLGY/1QZpmhBACyAREJZpTCPVh6N
UsE66vxwWuSffhqTvbt+1NK1T+IuhsPFdbuuYZaRjjBWexbbiuatk8iMpEFaFVLC
gCajw9iqD5gHg0aWlCD/NRiUm4ObiAXmEZnDVGHTxFwNDARmABG1n8alYHyzZwiN
UFMiGHMFMXQmWEM+2lNwxKgM89I7ajsNbAgjviqY++R9joN+GfMoC9KrybXjiat6
akaIw/1tjlPZnJFe/2QX3BIqP8O1irB7/2CFCMZTrDtuBbuFx7NV0cxCWObFAImw
oeT+9cxQzC8cqX07PAaSgVwCHyLKzjBbFVzHQ1RkZZkW8qYG2vtJEtGt0Q468e0R
ji8Km7MenoZSuTMeJdMNiKzPQehTpVS/NciABZUravAAxbjOhNfoR7Qq9Z5iZugs
ET5vapuSJ/qKEQh0xqFgIw/LbrGcqgZZpcgha7YVlw4vyUVT0r5OmTZbjAJs6lBG
PahjUvBj0Y6vel+JskUR/HNI6eXZ0M4xj1UIQzygrIUfBQv6Z0GBr8KsdsXdkKy5
h0IeZzFfSr+axlWwauYHDApOK/SCr1uPOD5N2PjiBB3d/AjG3wh/tzv1yxfeAFsQ
M/wiMHMPxUo8zy41hYgPrMw/l1eR8eBnh2TmIu+10D7VHKBprAK7thoZVv9nsA1N
/K+8ukXKUpsqDvGvxqguL00PSnLG0wCyCT4daj6CNQs2+hgpB0YsF04DdJ3zfMfi
3JXUVk57hXkYpELawtvnT5ClPbbyzBUZeIxE85xrqLJKrQWgLe41p7KGTb6CamXj
XUJmUvMa2Wr94snJLtgCrhHaSzaHcbzfNaWshjt0zZpoiBf/uZ7DWQ3axcgy0uWF
ks1+4PihxWjCDFlS2FDR5mahUPlN+OXyrEzKyeAlwP/PhfKQ53JE0qL5gEGX1dTL
DaFfp31o6kPhdcABxq7goKhlvc2bn+6m1JECLT2Q3t0nCPkxBcxn7KNXvHlw4vnE
pZJauhm0fq4bu6rq7VClUds+on1ROM7a2Z3z2GMmWUwqxIaU9pTRGvNespIq8wuu
A6EORmlrPoCKFUM21BOSlzbcuvUN4PYPYHHCbMtMKsHg8pAIZZydSeXHzOYyLZsd
C3VdEZuS+JN7cywOVhcWWQ3Ad30yshrlyjQy18DkRUzY4ANfKxBk9xfOnKyRSLDO
TpQmqRoiiYT1W/9UJgzOQD2cEHCNrGdCGGO23eKhRG36d0tTLJY5+WfsUroskbpY
WD7x5pyp2QCxh42eiRTvL4GkEaNhS+++kGKi3DkrfcIgi0ELzd+4w0rPZk0/vTK2
qaHBO/j07Z8G0HkhId2/bUfW1XaI4x+B/VRAwkf5hUvNvmQaGmbLh89ghDzT/Dj3
AwfLirXQpmIrX6U95BIek7bn7neKettHDkK2OJ9pxHUWBw/yqUhJlw3mVZ9R+uZK
6a9q6KxnYL+BUTw0HviA+r/haRr+slCYpp7Wt0Hu6IzqLIO5+61kp8FS1FAeXGSi
lJs7B5CJwCPLhLr/IbaZ6H7VgDsVtCzzagtVNRrPifgS2C0s4z+JOKEv4ONJwH84
QBhIFTDp6fqHCR4g4IlLoSBleRtp/Yck6eXbJVzG1D3PkiqOogA2CyuMZ4k7ZEr7
V5LKYbDtIr81DJrEE+o9vivHW7KPyImNHm5X9aFfYtbVuTDa83X3BNLDpFmSDX1f
PgDdsgFvmFc5QKihAoyfymSSGV1qQfXnWVKI9BG4ldajgVC04HRmpEHJPGhye1ef
jxKEmOcmCBtdEldpMG73Ly3VY9ApDzsOAMrcMnfy78WRgL9wJmsCKM6nYLKKIdU6
Cg78r6uSx1KiSIsU3Q3JFGrvsRBYC5Emnu4DALk8Ta5mINGWLWg+ecnrGoAxkglg
aqJ0K14EX03e0y4GZYthsC4um2i5yNJFX5ne1aWBFxtH4oryyYhPEZQCckWKL5Ru
OIPubD7gF4ujyX3xJCf77iPDalCRfrvubPpi9fmHyUQLhdSqY5uvO0oUXJGrWeqB
613M4F7rQa13kI9gkLcoEfzGJyuiegGo966D6w8pzOJ7XMgy2t/hHXc+MaUzyLBN
WO2inHhHXmTB3ZToI066WZCiqZJ7JmtHE7PeMcGx3CKZBWxKIODqD2LXnh+K0HJV
3QCzSh26r9kVgAtPwSdr6zAVoz2+uYwsa5yg3OF9qApJ9htYKkCCLLcwUcU6PhU4
BUA+C87FoXziAsD8Riu8+4seY/VijzYQf45NXnZIPuwdVTInBwiaoZRfk6IewUYA
4HdjPJmjnGVhyJiv+V3Kq2rE3Vc5fi5MhysAre8hbpLMvMUPcWPfz5nkyooBxo2d
E+uSfJN/xz5Zr8+d5OkA+TUgpaLPzGnXx9XPWxCiLnrD+ofy0FaoHFRFTNs4G33E
k5QdsPDq9l9MzLa2bE9+rcTY+c2MPCGdfc2kEJHOrxKt0RjAi9U0t3v6QZSSLJcY
cEBlRqHHZYzxNaQ8CiO92TzYqDnEnz80H/A8cxpv3v8NaDMOWgOSZoQmxnwSVYsV
Z0rhqFFfLXJLjNhvGdaWrhAzezwOEh2XElyM+gIPiUpWNlp3ICUxxrMegoPJUIb8
RCwILdQKRxy+5ZvbAcRXtOCU5YGmmTlGp1zhxeUsvPUz2Bw3IQOGHWRJ3utkRRfJ
+PJhrAiHWZOVhihaGudMmPJGjbjhCvUcnMz9S8O6QZuigQbPBTG+1hkhlfoRZsvC
BkH/IdZxSlZgb0ov/wV03q/iMlRHb1HHbpz/6FwgPlL9+CgkmICZQWUPT9pVk/sD
0iqQc2AC8gr0lfZJM2ZNqrGQuOmfAdQU+5xGlwH9B9ymRc/2VsP6QFvCj0TEypFQ
2AUtv+7KEbVKp9+3EBh6nQ2ogdnFglDpKa+zR1Je1fl4XCCoLrKa8bZcx95Lnsjx
K1Fyw3+2P8MmTzGNiNYqhC+FTGqQoONpWScC6awZM+Ceq6CF49tL/61ykxOU3QBQ
+dxNgSSGecnRoRWLvfQeSuibU874fmgh45QW63tp1/dKAmAQ7dKw0lSh5qEbsXah
xe9ZuJ+CJzVbmq+EQbZDBqAbBJOLHQ51y+rUjP4MD8qxQrnl6Rn2C/z0q3qI68WS
IGEbQCkyPPB+oALkB5vwsm5u3i1sOPgkQ6EymLiuKBJmwkuiVvkT1LYYupudpZCL
mBO41aLuyxfO4EmUYvs39bRfe66iV6eKUseHFAhegSrvcwga3Rh9UHRXxG6pGWmM
5jM4WEgk7+nwPeEIQ7VU65rdPWXBhU/6QiUzTOErYmkf/5J6GYEuqhSibtWcHfH5
gTtWCDW2B1vR3uEJszd0Z0+Zby86XmUTeyJ34H15x7urxyUM9YUfLT9rKv5x+dyI
ryZqsyHk/MBAV56OQXVGJ+j3VNGxV7T3DtMPbPNxrY8dkAQysUoetoyHxcdldHUH
8529F9CihJX5iCXkyx3dzs4qx2xOwPsHXgNzN63immKK1naLc0HRpuihji5IKx8V
DdiNsjutG6OTxD/DO/tSAtbPARt2ARXnryIHbGhC1q8NH9x7nzALpXP/90CnibUs
BfPVD2IZSVs3ET9TFprezjXfdiT/9o3RTFX9kYvhd4yJuZnQJ3FCxmY3fiUkzjt2
Y7X0mLrtR9QmTCmXrPiwM1IaR0KR78jvCwfQc1wnNleQofQHliSywPwq0jQPVMyG
vYCylr1breLM2oEMtmqPTXu3OWvkY8GNZdv+Rq6x5d/0Bhrrt1ndsccRjrz2vRep
0p/3zrdDeQpywZpYbiildKphKBTtfWO6Pa+vJzmOHjyZp/qesixh32UkHyU1vdTb
DNm7TC4MI1NDTb0v8rWc8rgWPyPCffPeRM510TPS05fgy9D3gxxpIfrfX+TtuaFj
wewwu+Rhwm97ihXEOaTJX57yL5gYU61F62G0bPtW74Tragaohbow35PYlK9NFrsF
LOzOIYKf0sTWbIDM5nWR6cVvSZUTHsyBTr8AkhvGFnUsq6kDJFivM29r8mcMlThE
GOIvD1zR47s8UQq0SSEUsFFtRbZZfMuAyujDGRbTM4CAqYt2EWPGnEjBYbffNvwr
n+cCf3ZU+NWOtEmLNjct+2VYCfPA704MQQurMCbI6BaqNnUhW8dgO1CVv0PDxRrz
prqq+62/aotK73JxAgfQSYTImIPO1wXhpB2B36uNoLX2vrtJ2lzylyYFMQxnDUIW
SYodLOm3eNDE8fayQMwDl3ZjBX0yh8UqTFbCwiLtH8oMkEdl7uN3+EenA/Dkgrwh
snNP0ExdNoI2I557lqXiSav8WZSpAw2GzbXiGOWUqGO0vEF9BjWAnVeyeMQPG8z7
ooMnhY30q7g+bwEjRbeBszoENScjDSjKu3ONU9jNwWsLioTMaqavpajYmQxemneC
s8Pybo/c0k3+V0X3PzLlb7Len2P4w8pObt+VwvwgewY8Sv29YKcNcqjc4rkVQuk6
VBoedUY7JWnHjN2qSoaWWlPWWSWjOX5Q7jfBENU5SpA3jIOkuv/j1m//jXrPzRhz
1fdBqV+0Baafps1UOOsDjwVys9ds/FpJ8CscbWbt0aAUcdpaiYqCIHkP3yEmolIg
hvDqBDGlG9CKAOzp5bx5VyXpP6p/aScoFsOLkO84i07HSqCXuLOiLsIL5JHqhPcW
xQs8pk5oT3gbb1i/SQ8l3NdCKAGDLz8VN3Q7WNlS2SmiD/a+H8unNtg/JvuZ6qZX
FE4+RjHIoLEITKtZY0Z13qsNHHqYK8PqIq2l9SKnRogAUOBu572NuWPW0Ls0faS4
PjCWz1oJQRX11KCoBaqrK/JJbzwg/jvclaTkyk988bEpFWg5NGRoFbqbA5Oc+wqp
KKblBfAJWjawUHM7nlCy+PWUD5F+H0m0FId81IWj4KR4edjRak04iWn18mEGtmcZ
r+gCRv4ZtLCPipzIFUjDmZ0WFJb6HxcP8hh2eNHZE3DVblP9RsaDb8b1BTmzwb0H
Gmy9lAYH/1uC5rRGXinTJj6lhXVgNmESvoC1Qpp/uvJV7frF1C+A368Lj+kCUBRb
zTj7CHv0sfdYwJABqwm/u3kpZdmbKpcOg16drMvl9N0ar4mnZ6AcnpBhs9Y7Ip9p
xy6I0zRU6AZJvGcwRq8JJ5d1XlNvinJnTfZPXerPQwb+VVndY1BtJXBs63ZqYLws
7H0UlL5yGomlHvFGg+0gTh0bm+pmEHeJZOgjzIjomfgUIiOkZ2E1AdODHn1Ohz6D
2qO+JpMMCOzR/wtWFhy5y4d5YBY95iV3D5xKI+GM9qdxzKrdgHCWpQGgm+429Qs/
94aOLiRkm0DDhNd4UZ1nAgHvCKnpBg6ZI5/qI0/cMGHszKm1bMqjMxUVlBO9f7Hf
4AuBYrpOiMrvwnhD4RNp48YzZziAISgebRvzGiAOHWWFsqCMOBoVKHcF3Oxjq47F
k34OSuUsO60oVP4aF1vxLFgEzDaUsXClf79VojTjP+bOlpufqEuxRmhSchc0jwrN
40ZPqFWtTS5RhxHFYqHlOwKwohvET1F4VkMWlzWz8lgEiBUCxt44aR8lr0jq3o/i
oXeQeZsGsq278FObMuP5To1AcQA3MLxbzUrE95YuuC8Yy24phcaDcCK+bU9traF7
L8Ju0L0xTUz8RCQrGu1V1E2NsK91B/3L1JbsvUnjhuTwTAddEKfCDgeJTxPmEWNn
rhUzsuL2AdMEj5QhPhQgTBVWztDFZ37rTCRq3OcLx78vzLeLqQlHAyX2zBuqmK1m
NmeftGXS0/pbjFyaY7evQPmhweJApauCDYKGMIv1XcThrs1bJkvCgGAZOuuReTqa
jVfZT+CwWZmf3GRLnT0srhm6OXLauGvrYM9QiAyEO49i8rCfJM0or4VCHcOLYWrC
lRPD2KDVGzsGbLv6bA56jc8LzSw6NCi3UVxZqyoGTnlzUPVtlvyBc3q9apfJTR/4
zQ/TvdOJVpWXHiyHIzb/DeOVTg1rUVjEtq9nOPS0nolEq4D9n/Fv4lV4sZTbB+Re
Ba5LYSKpb0Vu5GfjctmePshr2tHXlMGytPmT9M5HwBL2tW6FJ6DWeKUpOtl80hdu
rcnB7y6fuCqPZ2+Hry/yNo10+DqERXyH2iXEbutafUqTDPnuC1wFyqaJO8smOTFX
F0C7EQk3BIqV7WTN7utw+spbAtsh70O8KZC79DpwqdBBZV8f15Un/spANseYsv3X
gdO1BZU3DuFNHhUBEBSLc3vCYCxZU7gHOA3LXIUfAoj+m8VkldeGcIDKk/cMXtVU
50BE4AsInd3RYCiDrL4lz6riqtC3oLKK4U4D2tc64BKVy62HLceKrLaS4JM8dbAE
cH3iW/lvnK1vvdxyWvHmvy+nucFDjHiDzL9dc+MNVbqh3S6YDhaLRBTlQcg90Pxh
3jJAlcq3t6eYYxa/BUC/XPoctYsHVnJj0qh8sGQE44lopts152if1aoaAts6snLB
8o5kmcPnHkHdR0+EAWuRuc9Fuxq/sqfSinA59vz8FDlS2ggVC5RGHsJEl9OEUvmB
PyaMpFAex8w7rR1TG76YKIIoYQR/aA91YDqA7gMmIZ7otzkLXcrzu9lOknbzYWE2
n+Nk4tB+GhxLYM1q3bEbOBoaddXQ2/oAC7CpktSickY3PMIK7hEWbNz/2bcmoIr7
E6YU7SYqTVSTeyIdfPdEn4ZU3Bkvgo+rY8WysFMCtjDQASPvmDRyKbiPh0pyTBk2
G+Aa4U9EQmBPhi50jiwEpH1TQVSB1ljYI6D/3ssqjtPpe8kBGo8PKEbWTAcJSkxM
RJ2cR4jtsT2cwt6MuuG3L60d6a2SsRocfl6qA7sck0qgJIgSvUGX0e3qAINZSK5y
Uo7fMYSex8D8sxHLaqbGMwf2s1kNZDLob+BfaMh6toTLMjOSEfOGXEV7keys+/Ue
v+j74qa2fT1ALe+YClawscMUyYTFPYg35rDQPqqZuq6MSO1PZRmrH7WNAHNz8toR
l0zShRBxkgy+xPdEqlfkWBcDtw9Uiut+xXhM5tN85Pl7qhz4tlrgHWyvYbWRo+9T
d11RTh037XQVzMtpe1v6WD2zbTJ1K1wIkUjABND7Y2qmfQ8/gIKnOD69VnnJvvBt
KL73pJXvRifQ+Wf+koPpa5mQa8zOASty1F7lBxmPFMcLlZCylcKKVkAw2v7XexL8
g2h9O42RhftZd7zl1FXnPLCOXrRNd5oubhMbs4cmWecJNJzdpdvOVpCx5JMw6484
07XDvsMyGHRfRmQtMh0r9uTwWulnEJrp50F6/Td/pqpQgoVba2fN8XYoHSCJQv6X
Xl4ohAeJ5Brn/FZhwlTCcgWRvcrCbo0X3JNdPUhWndae3H1cM06Hzx//74CuLL2p
cG7UEbBVUzHPf5TWlmaXJ1bZGIKEuM/qRXn/p81Ainq0uA8hBZ/TTpdk3VlFLZnB
L44/viTBUAWzANQ8KBS+2dXt7gzw3HUp8TKCBDHei1iBhAO/Ud82ofqABXfxTNX1
WhohKPkFubQT+HRTA25yrrd/oWAF7L2h/1xbgwhYebV+HHudwFx4RiWEXyQR6GmH
QTzvb7xQB4/bxwNHetx2MCFnasf5TPiDcQZ4aegnHtc7NK23I6rQvDtKndj6DJfq
g4hIzueFFNe77zxs3GPwXlW0pcZCt+BnUVmsflglq/ddq4xN60fsiQDsxEQo3mTW
3XKDQV8+jtoMN9/dqPp5aNC3y2U7sB/atrFJUaJYwwcLLbjAYqIIIW4U/MGZyCGF
CELQR7u71HofKXqJigjIFgDdYexpWubLDHMq/cjnzSH26YkP7Z6YG5NC2P9j+VYK
FMCDjMWVzCc+whK2+3XXXZk+4UvdROIoPges45kai0UhxvIn5GC/LAO9Schb3h5n
39WpM/0ukCRh7gkRka4qYjcQGXwDDNf6dfDPFFhOq4OkGtiU0oa0gpjrR9QVZpNC
yx4N520MyohZO6WX9U1t5CWlh4pH22HnDFUvb99CLu0P01kJDvNIyyvM54GJcDd/
jgKTL7WCCyDjakfk/niti+m/zbRTPOcdOrAUf5VUbLvdAvsnPK34zhpAFGBwMYwt
21Ew5pdCgqV/YwvyQ5jlVVKawQ+diS9nv4pGepllFV9IDb093gnBRtBBG2tF6azS
WnqGXyFMJiyS2MNV+zJU9o+DiUjVXKbUIBjE/KAH2En4qShvZ9rFsExAQ9cWlR/2
Io4OQ7rFCOISAxXKphwnC7pRSV9Dr14sCMRXJK3uF+q5Qtwnn+l74oDoXccQfZSJ
iMXy5mBt0GBw6oSdsgzsuSLF8UGzxXsUy9UDKHYM9qKKnHjLK/o1kCcll31tsFts
Vjp1zOlV5Ttd7A4IbwZ1p5wjuG3GnlshmZ8p7ta4YHXA1nhZfzsvs4dxcosJFoWb
2mHCYgu5dxoSMCftAYY7GFldtKGhgN/mGfmt8593neD1oDlajhfY4nmdzHTa63T/
uS5tp9ZoV8OCXKbI5p/tRHovCzbV//FkzdROUMah3JmkygfUvFLcO2WkN4jPZ+5U
HFLMjDFiwYm9UpybkvpkwnX1EvUqWuv1CBsNneNMQe4b1+mb1uO56DrzBP/VEF7c
/oGoOISmPlBFU09k5Rt/wiHMozm2nIYlFTyg5rg0LId93UUgpA5RWbuoKwginI7Z
rZ7ddGR6iwjkl7XcwprCSNigmHb8n4BkxwxmAuZBvvGRIWtgqbNfRLuVtUFPKA0d
bBtdq+i02sNg1R0ylADwePk9TsczWiky/ro5ioTXJrbwK59DJ0feWskMkJyrUzZU
ytIP9UQgZIJTD9dqk/QOLYXCxfznH99R8WtKGcm/fzIHUvW7bK6RrZkMEDdTFrvU
YA7kITBF+ERZzoB+TQLUsLFPnUP+7LHw6ftyx6j4Ha6cF7ad1b9T/Jcat3KNdRX/
TvacVk9yPiFgjsQiy2tmKB1HPuVhTYF362w8Yxev8wE+uO8L9MMGjtGhPBeaAmcj
zl2M+L4GtQmd5hHjniW7KW/MnzrF9OrIlnkjPUKVoL6upYmKesRSalMK2rmqdkVh
aY+ePo9UXQK0SHxhnfQTcNuLZk7ZjF1/ZAhWFHQzG8uwlThTJgnEb4XHLjKypaV0
g2Nu02PQfqmQd5jghVeiRnGwNnd8ST1U/PtpDa9u/5bjzSKj8RvvOSHgoP6bAH+6
kDaNafEtUe2CkEAhe0YcWJw8bVKY86C5uXdq5bJoWLlFZYIkNf8UcMcmxx/Dpyxz
KupyTalSMDmAYK7FO4Ml6QrkxvYTvIveGVMn+kdYxEBNcaHWUCby9Nxgi4xW86D9
l3tmnABNFKbmA4qOSxeTVve65mMJk3llgHFv0aGr90JrXQ6Qd/QSCTIfWhj4vSHD
dh0y7IRGHc0Xu2AZyMvq+776sVbLdGs2G6R60QAdbSg0yHX9lm04nXIXarYXNSaJ
O62qs3WSlKQ/cD36QyUI2/qIGobK5akQjQ933OqdPp9dDTfg4ogJy/0/XN3KCc8w
3fCNEnc3D3NUko//kRajjqtD+oDI6hWOswNmQzYH2AOO0vqCGn1zZxkFuIYjg6qd
qpaKaksjlA53n6gZwKw1ZAuNEwxBkDkXSBYwRVxYLqwqelHnvThsLlFEmnZ8K891
Zn+Fdp5I8GLJfBBu/YSQBfIbhScoe6lfq4qtQTAQswJnUK/KFnjhKD8qqNCJVuRG
O0lZlPpaffOgFQgVYb+3+FkMoZX1jkbK96kSQOcdA4YDLkbIyzssaDht4hlHXtRd
OuUSs9ERL2MoYE1HJqiTqT3RDPo+eMcH464fs4GHdGlv+p0DxMOPSqOntApEhz40
cdvDV+Cq+MAOwZXSzTsqHMTpxs6/+Qg3RhhIsdpB8kPPktZuCSu//TcLsZzZ47pw
F/OymKorh+bNAwwV9xwDtInOkoBNfwCH1D1RiYS2e1E5GaCSzqDdxAyp3XnElYXv
tYXUDlkPKaYYDvlUds+mdkE2U2z33xThMjcx+uy/1iaOsD0iqIGw4jOb0vHiUu2W
P7tVwEJVFb8wYI3VZoc/s53bsjYlFwqXQTDg5z7wIYqz6RYvT4LKN+7/No2cX33Y
CeWxDjmMoG7RdvsluQe1E6Wadh6oA6LRktQx0l7BUeXMCPbWPvaEEMWbJ1XVr+lP
44+RnCWkxgG27bO0xsgyhIcmn5MFLZBrJNaTDMMT7I91hdLmne/ycEhGqitvsmvp
TPa+EKMdECXPoSVY7XXQ0bQtAQPyqY3DEwjho7zHs5WjT2seH+cZaZIEUp5N4gWG
BvQ05clz9z7JyrrAp6ZWLMqLXs+wrqvl58yg16gI+eLuEbl+3d4iNBQKwCfpr/YG
dJ3Xpe1FXupG9vXZOyMDvXCHmbP4RhrJVL0VHAb2rD9aXVViDFEg4gK1X/gb36Cd
S+JEBWUAR4sVEvedar057tWJ2XVBzL647suBbSU1hb5ufQTOh73fkefzTvija1vH
e9brI6CHhshHMWK+67eCKn0KXt8rx6XdI2MvU/yrRYv4/Cg1aru/SgXoS1XPeVgk
nWqNOjgn3PP9JEYqljvGA02JwvRzNtVbPItfXD35i4vUsm3IwlNr4C+LWnoX+7X7
QtsBNW0NTHrgU3IaXmqL3+R2C7s8I8LJ5I+/jXDjMOjpsb+XyKqz3E/p0pK5Hz1i
aCUyhAs8lQcGZsSZikLDr6chCsP16fYL/wkZRrHFnQWm090LCfmbR1HQ24Ac240S
GmI430ARNLTB8fUGIwIAvqROLeciS6HhAxut8XlGH6EN66CAeYCIVhy0JrPf8KXK
5waVcEE7k2nbQ8/ekn5QRGCo9+vO5jql+9Khfyid/52Rj82IxyEUvH3T40LKEzxO
zoh5X8WvsYZeVTXrv9gaPNRPgzO/GTnLwaYGclWuHNcI5tbZcaGXfEEOKJLqTOrU
0KkisvgG2OVNAW63sZm3d7ZEzcfCmAZ6tWHMqgTliKOa38sFX4GFy62JSfp3VWnP
JJ2mrsGipLDbwG97jHyT0knvq4XTgevlRZOQmOoBSuCT5xSkptl2h/BvYoXIUFn9
F6g3ZA8gL+OqA3d5I7pISWDQbQHUTw43RAhrKR6CA/T94onjRr00Be+/Lw8LJCFS
IglvPg6+NCBoho1Y8kSPnIrxEYWf5IbhQbFfM8rCk6MhheKFpIwlsyEIH7u4Yps/
e4qA8gdagZxvYi+tJ7pP3y6jxX3IcdKW2hQaj502NhGkZRmkgI9ywvcFd84iSUwe
PxqmsUogn9z7d1OFu/53Ra9+cAx/oeESQrtF0Lm5zao2edBqTnuii5ZReNZDwYF4
W92UqGuzUeTyP4lazq9/ku190X1MTnmQwvl5J9pOAqdcIE5eJ9QCYUGlKTYtEe4O
Hr+ltfHo+kvvibKov8qx2KoEUkimmaLqJbDp2hRGfQG142EGJo94gbuZK+GfFo5+
SMs8nT17O0f0hQxJqgG/pUrUdhoSjQqXRo04igzBaEGCjp95jP4esFAWCQ7b39s1
/ct7IPl9SrCqVpOsATOfgvpPiHWv/bqhdw8QZ9WUjLtBBpEelV8zMwOiNZJojUJz
aO3Yd4aMf/QP9FdunIVhYbXMn4O+alxtuRb17fItin4xoy7qP/jbq1J3i4tKCkXw
ppDAut5uCJSL91AwuwDHD8U3aYPrCGZFE5zmsAPLkIZkgD4f6/Dw+cWeXkOsN0x3
dGsY84BzL3vDnWD+J5bKJ7voNPu9UuHRsMuykvquphwX8Ywq4scwYaV4cTfSIBqF
HMi1VryXTu3wpWSESBvI5SXbL9dDhdOO7Xn0BKql/NNCHN2rl2kJtdBwgQqEG8NG
g4IRDyEPFtRQAJFgFNzpn2loWxytVMzdZ3WQpU40Eyms3pTgrbQxGknxtSJhDpcR
M8ZuS03jTAVF929oXNRu/OMNFtJloXtp8fww10oUhvqz7zu37H/y5PWGHO+0T+bp
af54y5XpbP6bqXl64woHfuVctlR1qtprHFC7/HyZqeHiuxmNRiOg5yX6ENhBmCw7
fCy666fL3W6U0hBAtulV0/HcsLr9fQDH/TuZf8wj8LD0lJbaKC8wzaTlAbg59MKb
43FVtvT0WzmXMb99vYd5S/nKwnHkM3StUe+X5PHm3gHDGtKr5V98JVEo+P8sjDzC
XQtTnBPIF+qzPNwgOqg2o6flk92pYeicDNkTydEnVB/DUv+oFp84U64OYHhdV9hd
0EB8wDOrG/Apb3axtYOtSrPKIPbXEhpCtAOh7MTWgHW/cT8HjGz0IB2OLgaTMJYQ
enwCSFOcdmt/saxGBNvYh38lhkcdZQcfGY36msyFthdeoZQaNDqeZM+oVrLGW3s3
RenL2Mkaf4dssC/lF2tgVwzLvic3SLq5ikqFYxftTc4LgQSFlccagmEQvHc+7WgM
slgPchMZVjqnp2FHAoPXPqaw5WoPSH8POXOGTR/qKb3ZQniIIqwUDyOx5lehnkRW
pVWUZOZkUANGwnWBZmjInGVpZxNNtisB0DEQDnODlaGfPte23O7NPWDoIR1Vlq82
hnZ7jKI3sOpTKZxXyf69UfyqRZ4kG1KEFvfICosW6n7Ki4VG0w9zps6WRMA0mx15
io9kcvb67egPAtRD4FI+FPeUxMkviVrinD63GnBm65OHTwSyiitvWPr7AVeYhKZg
DIjChpj3I2Za4TTkD0VNpAcI19T4zbMeTP8UvDo+vbp9q8kzplKt5h+mLN5zbfcm
po6zVODtAX1fsqzsEd3MliTNwrLOXiVuT+GoL7hQrCRCdY4jaqRZHaDRK+iVaJAK
j8xwwkdJZtvmKn5LO93bF6UpmsCyYu6WWQ/JFrba1OrGwg39ijhMDy6fKVDBY9NR
g4v870YAmwvxWsuKmqN+V/C/dmmHvLTI5P0MOPp+wNEKhm/jY+4GlMKi+1RWKLyJ
uH+jPC7ym7v+2ks+idPDScZmBK9/YmLlfLHj7aaSozZuqBogW952UGreFKL6Mq3U
7ca3XcUwpfgZwMSOO+eqpNqcoA2wR2hPmr6Zw3nKSLGmyIVmxsMegVtdBrvbRGhT
C1vsSpTCAXi87SEnd/kSsOj5zEA4pZI5M7m7vGK6iClXtRKv8PI94EehDVOF4HE3
Qk/mDCzBmT0AZIdO93cYqQTJEmgATHG8VpfMWR4e0szrCLVilXhzRCd9HsZ3i1ad
8V8S/JCXDlq/WoGZpfsNWTSuxCuqrNzI/aTrgtGa6gGqTy3tK8mERyY8TopuY1eq
AVvtm+vUzSyeSESWSNEv3q/33H59V/FeGU91TajMaT+TviOMDGw8DR8Lpa2tKHGy
SU5p12vLW3u278XvIIzPa5SOXu/INf1+v4tHoGNkP8IKX27S5d8XRlIEu8AsyRqq
MBzdmPsZ4i9V6gE3vGzz2tEWmEGDSzPgYi7UAI0oYnnGGU7L0cHM/+f1P05KQvos
EWLM6IkG5/lkSGzbtu+iTcaJcoBbV/bbEEUb3jRnRLzVytXqa2DGqsxoDI11bw5E
nGz6el3ozOLrQ+cvn54NIuwkznxs5U8o9DMVmSW1NZt4YHsthTSAj6wR7AsZcNHI
y2zmDk/yz4oDkQ1+rRuEEYGh/021yBQ2N2Il0F7OC5auEZUv7KdbeR2S+CB18slU
BEaK4y8n1yrgHfPq0Ki5cNohRdnzAMl0fPgW7bxe++vEuSeyWjMaoy1gUJtwpYB4
n8loNIGEuruAdJISu4YFv4Uk+XFmCNzDB3u/+lIbwmv2Gva/J5hCkiQAx8Z+jDua
XYyg0XJJxddiLRxNwB2hgKKl4Dlqd5TtZc8fsUqh11WbVkGXOtdmZuR91YXftUF2
Axpd7x0RjRQQyOQzmw7ljo0rwWhq6QXCA8ERky4Egtz+DYQtTmyYQBqol5yiht0w
+SgwXZEY5LJn6V7y/0D03UvdhL7cN5oi9S8A0VmcOq672E9vCPCvc7mlXuE8iuOP
x4lcV9TEMRqNcVLVHgCskjKjgXSi9hdZ/NCRV80dt1ZUMLAzr9X9rt7ZNVL6zX8B
38bQz2kEVYAhCt7TizhS6CV+Lk5enMrg0/u8Wvd8b5gJTuLywWlu6h7eN93eLOjc
hyXoEoPlRQDoMQKVBOl4Chg5f67vm+CP4lMZDp7+eP0zjVUuKg8hwwRJWcmNTVk5
xZtnFnyLUFoq9wtCQkOqFyyeeI2S0mvUMUW5NBE4FsUeIHGwPT8kcOvPRiePYixb
5buKn53rtkyLU3pe9e0ixZdH06rntVa+UTxG6Rn1Vghv8AslUmJ2IEj39+yDMP6m
rNkZNYSN5CFNhmUXvJuCrzJcoA5TIIaL94yWiSJBuuoRXU7o7l4H17ni3nV9NILq
3jU3IBRjKBeNOGfP3EYGBUjL7/xhp3ZefGnzrvK5mvaXXZkJvQjSYeef/aMziC/9
FnXQApVoILHhFv6cFWQP9MyuWQG6h3EoYYCnJCgQnGit+DMWDtXHdZ+daKwQGX+4
FhBkMcSRQNZmE5DSffuF0ZAfDnIld7KbYruspKLtp1pKX/hksltieovKk7IeYo+R
DhOMB3wReP+x8WDTMF1tN3uxATU3FdVT86EBqRP9+oLjFhxzleB/SdqJo7rBMbFe
uiomkHKQeQFyZl0USxXvLsYGrANsCQU5SenL7M1mcdKmkL3OwFLyCsGG8qNGTpvm
nvS+T5d9gfaUlFgx3n9oGOxv0ah6rbHUuoFEBXkfGfg4zefK2WhesFLMA3x3GtxT
7hj1+bYorALwlYzIEdQOhhTpTIBd5u2rwN6fOmq0n+zM83Ce6ACY4j/9bMD+UL8M
dONa7IiPKG8ZQet3PZGC+C5ImGF2xeQ/p8bj/adq9nWqZl56Ifdb97g0PY9eu3lI
tH2wtvo/LF4nUsBkonzRLw47UOv5J+MwmLySZH6FAmCRsuN/cxfh1FLMsVFTxTFe
RPfiXjsbgtiAK6HOIqZyIy3ved/yTB1j6dTbAfMBW+xx6JlOUj2Xcn61T06CEgZO
xBD/OjBD4+rizn3xHXQZ8hbF/2LHXXO6g3YAUS5bHc8ns8d3cu8vYYBGMpq38CNs
ACOQRyVk00+t4JTfxabBpMShY7lsFqubXL36fAQ/DvFK+w9/nJHVj1Rluq5XPgnG
d01Z0sfJ/IkdhFmza4qlf+NCu3mtSoPVV5fJegukhM2fT5R29l/QgIxzoNxDgsOF
6AbTL5RpJAjx83TCdqR6/mZFjqsJEa4vv8bFHk1IJJlMFW1fq5NKHufghRlf9Ip3
L/Fy9YiQ+BmNRkloDU2tUgp7N48lvb95nGP0zTuRa0qOF3XT5veUIRSsUlwJYPF1
qmaKi0K82dIrIaDDW+54V5JC/Elxw9y+xkfXgxVurgziHa/NgrjeXwSB1ZouWXVM
nMDfSYYaQkZVDd2DygtFeV0XcY5NLcrUjbraydbOo5BpAIp19eMk9x7lDDfPIs+H
RdWAD1/Im1nV9Ad8erLzPfQq66OkJSrxOjmIkBgzP9WdZlL9F5G58CSCMv6pb5h2
xAGZYQhqPd0JLeG3C6T05J29UGmF4tL3qL1UUs3O/pju05cg6NSTR9ZK2toMvXIm
OV7eUDM3WAMM1DHgwloRuGiwFSJ/9rXcyxQF+EuP6hKmk9pU4Gv2kQV2ImAHhdvl
kBliYgCe+Y0qe+C7rVlbgvFjQhyiT/X6ft99WbDEKuoZazbkR5ZY0rDSrjTt0vTf
9KzSBlJolV+roCbMZBplij2Rw0UPEE62aW3KeOhYBXIB3RyM52Idq5ADjdAmivw0
dMIr8TYw1vzbCxzxGTsruRvpIL/Fa5xImosRRktoM9ncdrPwJjuW3dZPJQlSDI4+
7nvivFMAysbnRQmD2g55i5vDaBb30laxwWl1ygAWGkqWo/k3FOQW0LMpnWGqo3rE
r53wmBggtfASdbWlJEZcsW00KDqoIJNiNXWCLNcy+Zrn5z2r+aW3h4OK/z4omblv
D51fvHQNC6zi6htJJx0cAkv6MXABNIMwKwrviCofXG9IoR3fOBugYl8UfNJ0Q09i
mtpK1JBBikEvsHwQ2MTm2+Yk1RZoKda1rQDfS87HXjddv3w8j5yKZv1MtvPXBsoc
TJIYDssxOTPNm7qpZYAFVPSXkeZenRfne6gCPCXSnKuBs/K0uzzixQzQUf0AH2IV
ddsoUaokErsSpjxXFT2xLuONDE3cQm7HUMvzLqA6pk/1GA2JEW4PPw7S8ilcB5ll
YIs3y8eonelj+hjd8cuVXLfu3AVf1betImyp5G0yMPd4uM3nLxqBiw9vDe/cqfSO
hjkhRuWnUzIkOHopU2y5npwpnMrDXDhJLwftNjCdttbVaY+zKdLlM5h0IxfXn1WP
axMN+CQfyxxl87xAbgm8l1iLi9+0zfdh0nlcj72iQuFpuyevgqxFMbTwkCbMCJPO
xyaylVUfEFA4DYh8BwzxdNVu9P3DDNc4A9MKyagYf2VOzMhMf6+zGhffdZbfOhDE
ed/TxZx6E8CXZWxIVXmUMRmncCwwsN3TRgrqrq32PjXfa3kD3NLBb7yzGJYJx7mB
S3ast1BLm/BrST3Xj6AXBBcmgw3Q3QlQXlbGS0DrhdmwJpEc6w4ZpxJbwPgv2+Zj
rvF1ddinULdHFyHcTyZ2VjHjpuAHsJACnSWU5uEiY7O3Sj7+wEx+H+PxExK7P9c5
Nh9cd4QM/8zMUFz0OikiE5J3z9bumBQp+sXnOjhtfDPOkWYxLZqRqEKERa8BWcGA
L4u4pmlIICTO020aFa954ZJBn6qiLQkx0WnT6TAo+k1hJtBlp3ffK4INAlyOghsv
M9ctZybliT8rNlPIw54K4dxt5y3RAywCMR/KTQ7vlxjSjjiRuFSgFfLOdWvNjS/d
NmF4DwtGdbSVZjJ1q90YDRKkolGIq3HJCl8TZzPinniyKMIcmHBD3p80NfbKp+1R
scc2E91+wGHqqGDIwQEdLOObV58hByUyYsdyUbRGrXVImg/6QOHp0MDDEJkvkRB+
sI/+4nMZ9SypesmqXWdVSSBHpUyHkvTsHsR4BCFZ5re9jXh2V3h/0XUqqODN8qWA
NM4mcdOj1q5nnbjuANqTKoT9DefcNzDb5X5D/Qqy0Eqvyi5Bxdz2ARjGMktGxXUd
pfLigLte6uL3jkRC3iDqo+MOAsC7pj3XXFK8nVzlDzjwWQ7zosj2DvrbGm7enT2k
dDBFqkTFwmmitt5yNYqW7bReAnIWkkY8YyOehwWvzfvDRTxc36UYsOP91xpadQhh
psC8IGT/GK4Gaz+IORPt7yOLF0tVUffFAoHjeVy7ff213jEdJMeWtzLz/oC6w58w
kp/eZMM4xF3aHPnmIKInfkodRE5NlXSKjs4ML8q8eqcqDnPEyOIz+toYJqLJY/u0
Q0AHuwBh4skutksAXJr/tTxacXx0DF7XduzyBR5kgq/31gX79tO3xDcQ+KT2sGcS
Mh4YXVfj7GngdDLl4K30QZUyRjjX+FZErHNerlW7zMBCNFEQBtIVPagUurT3G/Fa
CitMxRoYnQX0O2jH9rcxx+uHLSNrWnOy3DPlIClqhsa5nfx19oDUw8v5H2patyYy
s+1WwzEnU8E2tA7jIHVrT+Vee7TXmRBDyucgTQ2/0DIGjKhzI3hu5d1P6hRJXETk
Xj4ZXFCusVrPwtTFajK0QgExYG+O70oKDYUVEvkmuCO0whQ4TlvnGqzkniKKJS21
uw373imxZu4ki4yRRmUqUAIlQtAbDbJSfBbKs/imTwg7cFthZtfRMOhBsjdU4J+7
ncxIhtWyQrr6d6L+CGKoqklg6GdyZxdwUc9UD03ZKUO4B+iwxC5tqChfobajUBH6
IG6r+hv501Oybi68ShyV1JXrA10Woxzzt1zzDZRZodlLXnXRwxyObGmEzMezBRmG
hxTMzmX1tx2nxA2LLiHxUapFwHtOMYT44yMA/zA8UYH/d2Kb6fdmOdz17RBhhzXd
ZScRWiJ1uNSUTae+2e/fBnx3axoj1JoGQQzT6hFLi8/YrUtZvprPCD2nSuY2ppmn
5F6+/SE/zI/3vkDuVBm/cMRUgIpG/JFFtDmVC88hb2GNDE1GGtdLt4EsHhVN8BQI
+q/8Um07hyqCPrvgt7uD1hpfiZfcuGLF9scAg24XaUPTUrnwwTvsoR0aD9Rpt2Hp
RlNSqrOCo06FkYZxMBg0lDjyDSGXjmO+Kn5zlvNDlKshUWlLIDXjLElHbkD4Aeji
fp6pAmRyN0p1ZpzyrQJ9ykpmYklS8uE7VXwzvVhIrAEbAwYpHpodA7HzSCmMQf65
yaTqwdKF6xllMr8WLBSJrx5TLDfRQ76hMmuCqfAPwYkiAj6GuH8eq5jFwznao0cx
BAu9xjMhtQDPLt0aaSSshbhckfFBKF6O2tDq98oHvZn7h8UG177Zjpl1PLAcy/2A
GvlPRFNrIiz5Q+7NGWzhtK54/KkfinSt3RALxqnZ+gUU3m+YMAskiloC4xDs5ETK
QMEF9IqWg7doqKNf4phDrJtyYNX9irKzSWEfcKDKKEDjfHuZ4LIWig6gZs0MUWp7
Y2FWIalm6jziptF0Rn2dRltK6TUJBbUzcdIjsk25jxGta70i+vLoRcwbmuoqgKuk
JSKEUElAq0ZgK7HJHIH8O8zRujrZcmbl3iWzyS1maIZ0VN9vm1eVjYOkSyHJTRVU
rvhR3N+fpZV7oWkouXgL+cYvf6FUivwVDsDEfGny9u7P4YKScpnSycqP/Su6pq/+
brtsjUu8U7EMj+pltAktlU0OlusjwyO/xYPHmhHWILmlXZewUdVCtYhvkO9appVv
dqhd6XAblvBdMApfXZRzyZnBo0o/6j8OLNdjYC1zcEOfD9kvVV6+cDZMt2e460xZ
gLppDahKN4kHNDNiz7uRB/ljqBNXs8OnDhCPGOobehlLMkSq0p3Nlx3DnHBLjzt2
044vlQkBEpUCftnKekiIqQEA0wRZDFAUUU4F+zGli2ahCJIyqk9JLAfbOH2kyTcF
zr2vNx1QVkWwJFQqUyuKJl3O9XHLKZhA+tuvBZLXmbymVOWbT5dOYzDZYzgONxCU
WcxsqIcJzFm8TMu+1U28huiSV7r/Q6xyR0PfLSifbp3DMN/F9LKS5xp/gW5l2s1s
h0ffIHkxZugrkK7GwXa3F4bmFyZEpSJjpXfjSQgabS7tmcd7gQpkiPWZ0ZSdnPnx
UqqADCkKDBfP9EZ8c5irYyGH0T08I3Nii7RHrUo+Mr1dAslGM81oA7E04zu31feB
JkACV5ho6O35FvBDflbg2pkt39ogaZkCavubbIN2VVdcahJbt6jqWFfiZVXrNJXC
LMIk/jZLapr/se6Osy4D2zQLHsdnleuNUm43NnMjm/TuAqrdtw/vu21lcPrcdQiZ
YUBqE2W3OV9eWKFqMS/21u6G3UvQnut+BdEQWYmmuuJeXDaXtOXIwiARqb2RBT8A
Mgrv9EIDIlGx9Uuwf/OHzYxqCqicny57ceNGv1qjvO58WJ3ptAucWbUwlinod0Kx
rwfGpJTjBO2a6vehVulmKAqm+Ih1IZEOIEtbpt5PysV95LOnxhy0G7xTg1XZDtcY
bRPcyMZIHswk2RK91QTwdwVpYs54tb1jMerh2eZw7BEu2DcNSyUQvikFBaa95kjy
h1OxVHc+j1ptkq6I0sJQcsJP4rMh3cL84qzw/6e14EcsvPcN+IOOatWODPU0TlAe
h8sWRZsmy8jlQAnbgeza8X3GnSks2TZrvIDxHysHjX9Amrs4xdb5BypHnRRPxq3G
ayY4xB3fKK30GJKwnY/KyJEocF2WKCPxk9damlRZjB+DM7T6mNlayMmIow1dHu1Q
T2rZFZJuLohURbUWXT4O4iP39TKqcuvp6IbB00m31izhcN1f3zCb7VboKliU8Xso
/WM6h/DmdpY6AXU+dolN56BOWxSu74MIdGRA9Gk02AfWzugrDqbZWzGLBvKR07be
7vsB8YHQkAObDZmqTuzQYeEStf46hjdAHiXsgRhwgI90pWwNmqfCDqqaekbGvzy9
pTg1q+8jrwCtpura+HjqcomBnf9J9LAmWIAL4EW344n166GYgomEpwwvkW6tOP68
sBVorWXfLHdW0/NWHLjTDkEs9r9wveRH/eBe7mHcY2p0fB5flA+SnUUsz9HhvBz7
yLaqmXmLgosdj47VhfwmucIU9msejn/JyN9lUb6aBqu9l59Rtu6HLPM0BN+lTx66
qDZR4hScIsjMNpVChXNEa2dxQtuMO4d6cO5SAcz+Y+MvdH/5etKG0exk5dzkCGiF
9GDuG2KjA5/n3gGhcpLHlmEuf7gyfG22pxVqUJMZnvTtaB/VNCg57sOKhiRQboDq
0DOUY4kgnU8ZtkA9Z6TAzfTF3NKyy3c8TRqxi34SldwqZRkn23Jx/gDmMT2wWRmO
JwTVv9lULtMgUmwhqq3ryj/eGLO/vRfgXe4queSfT3aHLUbs/nZo2haqw+1mqxrk
FNTt2bFMz0WbSkKHqJko3nVh6N/wIfILGJXSszlf8mO8aD0cPGlnn31VdWwF6oYk
oaJWsBX5WarL+/+ZGJ8OBp3PZ+a9moj4WXVjN+VVUm9UvmFpeG3ziP/ZmZ+j6fUl
D66mqVwVCUUJj0BCCh7IFEuEhKfOpEB3g0rRP0UjH1F7ajHandI2+BBL49iEJqov
N1dD/vcDJ3hL8ulgIK1zWhI9sp+EQE9UDaTKfAdC8DxRAYLJXYIkHaUtU8pmRdjY
QLelcSn9MZj09iThYvymcrUCMMDlkBm0TVE3lF+rEco73B5w5VRKqFFBRfPm2y5+
gO8dBQtb0NzwgTGKh+NSFMXrhRSXcvlgZfqdnCA/oygnzM0gM5E2iSDVvak9gpny
2q1+RPpJkD+9fdPYI9Fo3dXSMkcRVrnRrmlCBEoxwck1U1QkT1rrwMv+bAvWTWvX
R+S356WU96Pe5/SbJwGrXxu+z9/eEdZd4wLLWEBRjAlobJFYJzSVgHaXHGYLRfoW
58bWT6mHk8rb03uPdGVquK7RQ314dRRxp4etV7aJulzHI8P5hpEkkBwBUARR2ggX
vC1hA+e8JaSuVsx/5p8f2u3YXBVuvZVWl/Iow9TkEyqg3acM8UD4+pu3ykp+XVIk
e7YBlRwQHbuRbikSDRkq8Wm3ltJlE4qVge7X2Tx9CYbhZzc6nGw/gQDBhYQpr7Jl
CjLRd8001pp8KAym1aAPjIcKvrNoj7FdEUggAH+GSVMZHwBD4CMb6UfxSFRbZMQA
I4yiEIghgUI6+RzTiq20Jit6/LmuVTDn5QQrF5jX1lIpscEP29hvcAvKw+wHsemA
s+y3dGejNT8sSX5ovhE3KemkzjZq7lm79HumGHXBHgg1/FWko+W3og3KJgX2EyE7
FbqZMd5BdwGzodcN2fF+4HW9RXZxig1be/Oilm57XmV8hsyc/eT7ljSB2z/2ekz4
gOHdF3WJlzOpatHeNrTcYKi40GpqUKWUXEnsHX8W5dFWE0T8vfwIVt4X8Tlb5gfj
PDJwyeJojjH1lMMvxTdwR+A8mn3oydBY4R7LBu/nY503y2HdMfQRpjaACgrRlCF/
+NxgOZ9gWTXFCOGSdk8ExsB5Sp02Q0/hQtuarFeXKwgictfeLW/jvpb9LAnZuUTA
xAIbeE9oRdFXQNn7C4vkuxiL1eyP3HZoRsORyTTkqmxg1kMCS4Y5r//2nUgI4zmI
uyiRoxXwDnXB8XAo+/qcd20eiWU2TaFBpzvd3sPkN4xYTX3Rk1gg6KoKi3u/y2rq
oIaCnmHamN2LYyslWBswRPQkRhHEqiRdFwa+fWea6N5L5OhAY2ZpZhE4496Vcn/Q
ytxXElylbYAIyLKb8Os7Fep1F0QTPW3CTnfxdOIUMCZQ7mPBbVIMw2qkrlwLMA1o
/f5VYHrELk1EboFBqc2MsS6RS2vSMMsjAIJ+tWSusyV5ed9DOQnfzG7ibBR9aGrn
rASOM3x88ML3OgJZggni/NoFM5IPpXpbP5GpOaCvEwomsSLvSrh1ErL9RUpOL6CQ
Cd+SMsTduy7PNEo5qmNeCRnPxtFTIFV5IU6RmeBubAuH1Jfrn61LV0RiPSF3v8wF
tAS3+P0pPG81GaLwnnnC87nxzrbTtKRjq7Ln2fsk8Ea0M/8oHZLT2bmstbHIuK6e
hXXkwqHmYOHtEMLh5ZshKSKb0fmSAFZFVFoC6Z3T2JP+0V2lELTP6LpXKLy3aRX2
rC5edi9hYC4nRQm2fPflu+OlKsjiDTEmq9P5iohGRYOwaXMCei4nKNYTf/fIQw2n
gprkwoWSD09cr2xtv9QvOF8qfYCB6jAYIeBSVB7xxr7NlFZQNivDfo3b4OTLUDzg
OYqHCkQ3d/qkKqTh9bW1+6nYLxvIpdSlkOP2uwYvkluB9xge3UuIodQy2o1VdTcu
v4j7mXnfhA1smDr37gKvgfXABT8Be0ZuT13Hq5nIjTaST5qj88aAScXifXcOdFa/
pX5oqbK4OQd6PA4Gt7FU2hItINzfrIsu861eLSKJJLd2/s316xlGpSoq1AlC6LGG
1U/5oSKRSF7NEzj6sx/TySaPWEa6qVVBolhrXegTUm5zWeNaBXnT+Nw/XfBifxzF
FWudgVRtUUKTnsT8v1j6oilvwjrI8zj7GIu6NDSUZzhaMSTmb+K6rTzSL0ic56cz
fXfU3L6nWcdvTtBI0j3LktTg/tjClU38wRKJcnuernMqpa6kVIVc9UX37tAlVxNN
q+Gp+m7vPiawwznSrF674RSWxrm13NXYRUVXxlYkPWwNn6FSQMcjJoJmltOYkF/k
jdkvYMK65DiGZ1MUM1gRzodAzGNWAPerfvicXv4Wotanm7LP4cAEHC90Z84xVQuL
elv958AmtQG0HTiAAPBGOSmaywZsf9c0wDmXTP8U3+yFT5MNm10E6NmQcyhGAM6A
aDbslG6XaUqheGAYAiYpsG5X7qYXF7GqM95nAbH5JKdArEdWR1UxAmdaCoNRtM9m
RfsfVtI0ErJah5PkXLyAovtXixUrsPjXNqYX4wiAnnfG1ir1szgplpGredxl3ECz
MEZoi5lGVFoVqg9m8IDzu0daYE2WnpGxrs7y4LmcPZ9lJYExFkIUxGso8zmlo6u/
s2wZ8eHs2PaMGBeLspItxARGZOzhSIKlKoZ5jauyH733aGInbdGTkBW01BCVJJOU
WMgBDMaR2/HAtXKjrcAA7xSZlmw65KetGrNl8le/v2qmg3EuLKX6kvPPSEk5lVaR
DJ/lCJkHoGS00MYPl7DjENf1wHjiDQbwcl7XNyBcXKob9np2V55iAx6JroW5JcKb
3kilpnrd2U9o2MvcCqL0YG0xxjXiVxmN45qkfF//VyxZI0rNDeWLyqMoWBzzlUu9
mggGkU7Lo6G/kqwTHl2kpVntH23pTppFLCGuniPgRaQmx21axJ6hOOt02VGFipCe
AoddpCnsRwNuB+jTgDSWMPg6VmzR9HgKdlpEwA+uEOAnsmxpepuYXNMshuXV4Sha
lIPDmAe1Ridsnklh2qgyOP6LZ9UULM1R8xg3rjfHUsTRjqYOJi84Lg2R4HTiEZwi
qMEuV6dppl1S/Yseix54N9RHfDcKnQae7QrizEITQ2UiQReYgD7FtH1Xe0F1eduB
TVE/q9Mk7wvvrd0uoAwFfHj9VkN2aRH6+Fx242+8ImGVRLRB/hvZoWgw0CGnCQJg
Of95wjmoQq0PMXb+aZvGIMXPUsjRHz6wk64pwbqWqpvY73TWyhanfzUsQ1j+xxac
d645Lk5FJn1efXzP4kVXyBdmG0NgI3B1X2ogq9eijaI6F01iMwXet05NUqj37bEp
zjgjOoRSWpLQEMzcSuBTVcVq0t/NFOtXq3NKJQhbyX2IWBU6o8fe319Dq3J9h9l5
qNBXg6ARlQe6+Geg4xG+NFyP2Rujrtt+awjt5F7w+AAtiJgWnMgeP2sGY+ERON1x
sITEto1Mc52q915zE9YrTqmaZAM4+lSkFdHxBeIvxfe7Qh1UGko2iGqsmorLxBGU
zLSGqHzorW0fN6qpYZY57/y1s5C1wZ6CvBDA38flnE5NJ4YmWbUoPIKGlSo3d5TQ
46iU8zrgUU/ppRb2Wd+w4hO6wMTIii5nUyITtIbC79BTCFzL5I54/N5WUVHIN9Cq
vR3YlA48ZMv8DOzDqSuMIAW4mL9ZQb973eS8iwc8ilCjiwfZag5eN/hztwVBKXQK
07NZiUajUqS9mRCdcO6JVqllB2ubECctnQOR03+2IBZ/leLuSsBs8U7ZZAUP+kRr
G5ooMmr/7c0xRxtCvNEiMxLIU3vEnApZHXtZmOxqf2jh18IL3zcy/mYeRqNXVZw+
PFy/IiWG3gkIYUj1f0as0GSnD2wcBpu880hBIb45/TEI1pAbws99jGwSSWrgizyk
sjcSfRRKU+zg6MAMWy+UVEjqSuqvHnjfd1qWUCh2VPS9Zdyw99oNG5YHYkNybKb/
VwiCdxvvPmiWYbT0Kl/Z4K7ztJDoj7X7SZ9LewqRTOOwYpArth41Pqmka9giJ8/D
KutHK0+KCQ0bOlJeWJZQkLNQSAVSmn8dizeWXydMNczvAe9BKh4zpkoUsiONYf8O
+Qz60cfWeJZ/hiUu6nVuj4t0KFcypWjnEnO/F8Yr9y+nWO/TDnNMT9feSNuM55UQ
x9dTVx/2OWMazwvnvII8DT/aXgFO2lVBELueXcGHOwGvzYmOLdYpjIJXiAJW2qeH
vjyEQAXWXU5u2lUxJaHrrnSBkcw8RYmmVfzs9R1brJbCTW7U+tBre1nmJ96gGJ2l
2XZggKc8Bm+lr2uHfUT8Rp48qONs3s4qj0tw0Ww4BMpnWkEsXCyspECWZDopDhkL
hKabHEkxZhm8T0ctbvehuobjq3ZzV/gx8+ra985zB6LZBO6SZXXIjjZEadL2rUeU
IrYmUy0ICRAhp9Qeo27J0Aezvlsxv8TsSTun2KcDnXPrxYuMHC5Uu5KjLaw4TUui
XyTgKkFv2sfLTXf4anutnCL12dV/ZbvjuzMolcT0+/3ZB1/BHusnnQlq2M5+gkCk
Q96Nvz14NLYcAHgiu2r+CRHyYeZW2B4sssMWyzmdvRapUydtRdnAhO+2OpCeAjg/
igbfPawxmHXWJJsr7+pY90PBsMP+li2tHSw/29hp2oV9g9qRZ0wJROaiaBdic/vr
9cVoAL1MhicqafMOO/wqQLsAzFYsthvkJs3ZugA0LGDXemJNQNDeguKBH2D24d9T
rlxQCApZceoStFe+rFWYioNjKsXcR1Npcyhmw8FFG3DkkNKeU1vaBqssd/Nt4Ha+
n88BKJp68JeIYu06tTYpXNsxxGv73INxYuYsogsSgxvjefJzUqtTeOerK/8fm7tI
VVpU44Hkrcs46bjJ6n6qBoSbd7WRjUezLC/xFPFzxm7ODL/oZyfFeh0HBMuJ2Rrw
01iTpIae0i9WJJBDa3DamEalaE9iNzfWsGumylgcaxa21T9ATRgnA2OcOmhXzntS
SIpcnY6r60MlPOy1RNvvPc09eHxxzEuBPgTB21k36k7FShHc8fZVVDT7KBc/alR2
q0UURlhSNVsDzFhlnm+89XPNy9pVfjZmeH+zZngzmtLh/jEAqcNzaQtijPYqlL63
fbE7afA309SAlZzj+8Pz/k3Ln15pd27ER7JzmRS0eP0MZHYo/FiL+jn567iWkVuo
YZ/OaW3eRcTLdMBWGePsERp801dGPnif+dyoH8BNBDDk58cqBwKik/tIvuifJP/b
UvWvWfiPIin6M3uh1MetYV+3lUrNHK/wVAGgrPnC8Rl5HRmbUYL7Hv09xT9Qwz37
TdtADo7omvrPqI4mX0KV5ZfsAmoWFiY8ChZoYIgPFtQpm7fo4mlfo2IDJpvAI0Vv
cQDKZqgwERE6GWeByt90l5BUv+voYfOWkNTgfqmj/Yh3gD7dSg/Dev7tgmf1UUqK
vSDn9NfqScK9phxFu0d39wJSdECMmauhSFlxJcRKxNZaMkdWM324V/z+1Sq1JEZ5
YjtGpj+W8uu2zQQWx2/AZ/PF5A6ypCGKwgBx6esfmK2kXmx9U+mWb2VTLIKL0APm
KB0rode9Ir7du/H5Up21B/usp0pbyvWum2s8dGDDGQReSi/8Wrl3Ke2litr1VUTt
dd/0yGCPZwKXLeYuLJPiJLfgEuoPtk5vuDUTLiP8PkqbfV/NUHPPeXHg87m6RbVU
tCMWgzuQfTqRxJ2Q1JJ3Pk0XVy5iNoIgopXf6mZEt0ikQkrAgBzp3S1Mq6vP83Aw
TB943YByj73owZoE2wRFz9HmlpPQa3zmeYgMSabF1ZVCWn6fQTsuwyAnHLHTmNkF
tUBpp1ZG8abQk0tfkJCsLas06RMJ9sCb77a4fimteH0LkBAw4hQ2iNsGS6thrvLI
VHpwyEiKCUyeNhEWj5/8N8uqNB/ncU5EbWVYsg51UHplmSlNq2enH2zjQgsHn07C
fpUCMAcC2nLjx0alzfE11y1Z638zAreAmLI/qSdvV0rW9x737z8CIH6edbzKHwmH
gRbDDcZ9vnU3riPTIjKYwGRrB6C0uQMNVA5F86v63FOT1sn+/gjjcO1dgjmiw2hB
BsBrimI0bWaS7pok1hl/4kapf4c2a2nNIGNY3HmllhtlQAwfEBZBnlXuNHcVFekf
1Wz0POKFOoIIVpKIc5L0NxO/SWPbpX21pn/sndF2sberkoWFdFlexvAkYwdsKIq2
YkFzSL5VEnZyaGeE2VeYqJQFO7dvvu3eR19C6rYvR7nmB1Mr5zSfmhMebYld3uDR
0bxT3QgBDSVnO7Idw/p3YEUdUxfawWzCmQudc6JwxD4Uw9nMM1sbhe7utif5VYym
Xhm2hKFMoGgScZLfxA3r8J4KcQttdDDzMNc1Jw2x7FycIosWfqe2yoxUT2TSg98L
A1bYrG0ZSVtEP1o0lLXgGbBRnkYzcCszl1FKnLMZOv6u//7qG6DinR+bMnKxltjb
MmMTgHVJ+Gj1MEGpbsqFM1Sw9dMPOqOv+HRWhfbTVdsO2GDzkQiMXTcuqOPE3WDs
reO75Phc1tnpsP1DTWlp/JrIuAUFQwnUqRjUZ4DmxuTgO5PXN01DFfsnWdREfLOt
WUiSv3KokywbGEvxJvFsFqQAn1tKT6gFU6TqgT8jaDg2rufatBaFqZ/0sdZL1lSe
gjC3kwomKSUnI1twvE6rpp2stkfJ9giZuj3uGkS7TEIAxs5VVCH9N+mfOT/LNrqX
Bha4pJAcOG1YuBw5HlwQSyRllylKVhUWG9zgjD9lZkiydHWqbzklEmlwfvzvGXH4
hlvsw05/g6tmuU7IsAC/iighwwQVV6rJERGxXXG7auhC5CmNC3gRAqTg3TMpacTy
rXBjReqEfQ3jAMrTPVcCyuob9K8Ctj1eMeaB2Et7V2BZ8D7gEDCABbOxuPxZcACs
w2o60NRYwgTJaNMT+tfF0xCrBQzGx68SrmzzC0kL/nI7G4a0Kn/mHnKNatmpOmJf
1W9maumK111ufGr0ekbgFs/WOcaazuhkkvgw1M/aNcP8oHkEDLK9nNhB/CFfJMB0
cWQ+jBS9ljkWfm8uCaNq7SqEFpwhtlqsxRNJ4Gx9lAw9BdCuPTMZwZbGGai4UcC2
cltYeSkx6tXvlfThELiC5HSae3XIv6LIhXv6ZcvSM7ekYQduiYd4Cfy6Q+XNRCq5
q+9UVUyMHmAZK6Bn+4HjGF+fZdzS13jp1YWzR837DUpu8gGcYuOK2/QebN6YH5Br
nbOyuN1W2fta8OO9i/zd/X3z4sKQDpIdUiMR21+pvdsDJBUiA58fIUUIgn50D5BP
lPdecDpejcpexTVbHJ/9TQwFBoNsEu5oLIC9swcYJjkivb9J37T23rtCxW6Cu6l/
2sXz8I8wm1VJZH7nzRsht3hCDwOdpqrBTrqTNuaViDl2bFDfSNRAoNelqqP9X5R/
IcxvIZ2rCC75E6zXDsqqmqqLTRHqsObktWXmKDrWHWrL+ZzYw+SH3N8sRbIAzPry
+8z/efyu18HjUjsIfRgwqkafVQQ4A2P3U+r07/ephTf64sUodmHiDWBr5U7U6f+E
KmGn8ysHrMZG3ZgCqhzy1ooNGsnew62QnEhYtnfcuSkeWLvTzEY6dVngRqYwb5jT
KO6QSWYpWxzrTtNgYXecfyU/t3BtCR3zt11jKpwRzFl8lCVzf+QRMbiCGRtmOt6n
+lgwDNhiH93EhrGtiNxCD56g0WlWuAaB0pDW0dYgMnY7CUlOuwTjdKL2B4sU2qmy
5/HGkP/Y7Vn95Ux31N1s9Swi6/zg6b2BHtw2jN5EcZpW2JSiotR5yhZt3lRCRmwt
CZE3kfm2+h3VLmKM6l76WR/r5szeBm6yAfz0gjYqb/NCeY42J7Z4RYl8vP7BaHvu
MR/Mk13r27YV6fBGrvcEW4WlkdAd8CCbJWKqbNTcptrQDl86jtWHAxDMJGaEBMvI
ysxeJsu0BMoV50CsaEuB02tw+cQ858S8dV5f3EUJ6/VdUigg9vDvQkqSJU5PgAyq
hLGVfhB1Ld9nG3NhvoTaxUlZv4vLJBt0DmMA3gfvu9c41meAAC52ki8viOO3FNyc
LxMhFMulC/hq9GpOsXdI4ELQYfKgdVLjx9TFiltgruemxo4UUNUtBzj68bnkzQmS
cIWlaO7eKUB6esDODDiCZzI3lkhPhI8dBFzzlNv5uSq1Cz4v+aFjSepkgwB9ZTNe
CAjAiRqrC52jMMevtAGDyzFtSYt7reyi9WUaHEM5WQbfmv4X+o3EraNMB8QCGrDH
Ias7jcHodX/IJDO7a97hcZe3l9QDGsbggwjs0z2viJIErrJGctFVslni5fKxZ5Ic
b5kuCxphRkNUp8P0+WZYxJMtzl+R1lLhd+QgqKTAoR3iux0MDUx81EjZ3frU7d8f
WENu6Z7ZfxwKRdd8GIztze0Lj9ge+L/fd2rT0c7SdJCrpWsPvvm4uCakZugNVpdr
5FmN7EdxEj73Iu40VHJWpaHxQcI1cqag/NzOK/dNeL9q7GriT+9o+iBp7eLPBc5t
HG5Wm4hw7whMJaSkw1wPZSUFLZAPavMTy4PapJAOQ3HvwvqzNmJVt0mOHTc1Zmoj
AKzDWyL5bbaiIfZdcIkfnUftLSSBY0TMBh/vBldC5MybtP3tncR/8bcm/nE6S/ow
OQjMX5JEP3Ip5R2hua26GKUL9EDvm0uAb0A18fPS2oUkD7pppgF+zOozd9/RNpxS
eet43MtBgRibrJ4TJMLAYCVtSdngM9uS88fSeflKY7gT9fxX5f/2SwlMjUKMQiHk
V0gQra2MMFUCIx7k6MdccgX/gpB3a5wHePnG0VPwzgMDPWaN1jWGVGYT433Rjhvz
L5wrrsSaGujpNEI//gOSf1aCQPm49BuFxUicJ6jHJswsQVGZapL4dyel/0BJd5D5
rj/hhCMHXBi33J7NhV7FG5klRpiOuV9/PesKkdxw1z4EHP3pAaUd6h5erot1xFll
3cQ1NN6IJ/rrVJiCsQAqI55mzNWU+9lu8//EBp6D/RVGo852sWLIgb3TmyRwrNyv
il9CqqInjAMcuBDKQfGku0I70xQBaV/UmpqDocmL97zkD2bj8pKTQ8qyBSFMzMlu
NR7NugwobBbFjSGB21JKa7/beawrPh//EbDaWJBWDx1CwEbqm+iEhcknyvXN0TnJ
UTAkLiPYUxy+iQiYsP1+K32G3m6tQm+ibittUSYWigfdKfpRtau6kT/8jNS5TKMY
k8lwKbln8uOUbkNI0aqM2GsRIXeFAl3lPnO52APdoB3j96fS6q98elCsGDOXRFMb
EoG1JK7RMTHOgri6HPm8r4OT1EsMsEoA0Sx4lCmU88CzNtCypOIKg4OdyaQSxYmC
7/RRBBFrNqlQBNVB63AQ5AcMPHjaTDuXtScNWVmNDWjDFQbWe3qWAqHf+TjAjmK/
w3pIah1sM9xCCbCa4BHMwYg5QVgmj7XS4c5bhgMr5RiT4hZlNeMCHUUCWNqd4wvi
fWcT0AR8zCa8VFsoBwRPQvqyz+YJsLIf4C/DTfGZoIrqXSsiYP0ihsZpU+Sgw7n0
M6EbKyNucSvQpTnJaNl8E8MuO8dmgG5F/T2sIDdpugL6uq+L6sJu1OFr1L3aFl9P
iLUufdLtvUTF/GS1T8T2FNl7ZaRttIuVdJitUa5qlpMLFkza8pmKjNGAA51T72oU
ytHFd+LRc/ny+sLoWvW1FsZxN5vlqAEu1/mSltAvjw2mE40WVnwQ45/Z8vYixOjN
zBQdYvMTzhLvIMyQBfjrQ3yXHtFWfmnFiqwFw9sG9EXqmBCwGPZ/HM6l0AC9/PUY
Ut/4AOnh2xSWh/neeFwW9gjpFZYVslu5OutjBnr8z+W0UV9Mit/BtuyL3vsTaDO8
gFNQE5+1ssXmOQCBwJ6fg0IpyzxOXF3E+091jTW/ncLQ921/vpMDPB3jVb38kWv7
mwsxM6Qdx6VBUVDIIVVsSntp4QbAumlOvTXbWOFGXhYD/vNaI89vUzwHrnHi8NRe
KUuFO9+YLwUM+/XDFcGxVURwSzwnGj5eHqazTL3tUTsxoihbi0JWlJMTsLd5oMgA
Qzk10SfKBqZA7yL785WTR2PLdwX+CCgbuBuQr2BScKZRa337DtcrNJvk68WYYg3l
hgGyd6malAehJyac12cZtu+cSCguUHEQebpg8aIRT6RDWnKfBvIVvwRudgFv+uqw
E2E038QWMU0YPMo5BTY0rFYKwEH1w7HWeRAcanlJ7RaP3Xm2GLM1Czl3W8nIrfED
iQuDozsEffTzpHjdQj29izaLV5M6OEcElo26cCU6J7h8Yf2VsYkm+EvvArLkJtiI
aVakoUm2StnA67quwRpi2hHnX1jA2ahh8osTGKbkV//uqSAzAszSc6VhScjckpEB
/lRdm0c1AKyOr8GiLis6uG3ZPocQW9yZD+exSpwG4nvPcL7Enx8IwXvrEzft0PIq
YiGYrC9WieYs3WJUz3SUzviI3SpTTeCGJZcwpwMoF32XmjSfQtgWYH1P/EPisWtA
NTRLxFyYWv7/REn/4c0glQlVct/RR2s0XTTdYxHQQQfPJnLEspu/BkbTt1fnlB0y
GjbZCPZt+aLoN8b9E3e+xlhKNEgBj4AC/1srnRqN+h+VqLAZ9ohHJklZn8Fdt4nE
Nxtg3uYw8MQMjJgF/fzDXH+GIwZIzYWZ5AhI5J9yhnj3PHnPwzQ8kIuV0imZUuiX
HSpsBaG1NhLHHltlTcozwLNmxHa/MwqCtVii58rv5r3BkaYUWzytd92Uf55MlVxs
iSuNi3i4vrlWTp/L4pJbcErtoWX/lR8h1kUnBDjqp/vuHlnxSLt932nSWqINc5Rz
MNUu8pdHyYXatO4ZTUUSuz1qDyQlbVpgGaTGkzjldD9aGD2zfUzO9SK2gWHc1/9U
IpA18dv7sx9KIBurbmTtSZlHZA1eSO/1Azdy7ylpkOmiZElfJts9ahcOVUfijLhB
tjfOqixbx7jnPpMpbTm9Yc4LY8wOhH5ggF8mS0Njgt7D6z51zRAOAn10fxP650tT
t5NSV4AYQx3JAwMPU9+pmipmZQpss7I4RaVjyPYxVtDZLqXmjoaw0PC+uYRXcqL2
z3aoaysNjhQd4KnWPcEjmY4byXHUIc+Mlr/XmmTY/kl+0qikMGbTRwiIl+0ImwTx
syh1PS2wDNJ70gOfqDFkx3ihPv+mmBmigbsclao7BUx4zmHP58KZSbf2NZ3P3m92
lxT6SRHYRocCItpE4YVmYXGmvx7nk9spWhG+KReSTKkjUGz/WImoJoiREAMbGr1P
fbpL9JrlN/2wWn/KMM/pbh4Ngvj6RzLjZURPvI329AlRiNOYARnY0Wruehg7gCSk
7LJ1PsJPSI55iDvToSVtLvbX0grqxIZd4pfkXd76708aYEYMuFIIGQyDjHIfRSpz
3DkInm1G+sQMXNHKSU9TWxHR7AIXpnJ+yaDkbjjbJOHJ7TmJutpd2KKdWcIWBbHc
dECDkLgfishnc39R6PwBXALNQ9xLmDH8tSTKnsunk017gee0t/2HUmDHQrzIqurU
9TVXfc8MNsxOi3dvSkapsSA1JKRqypkVZrZQPGeuRuO0399LmQoHE0Lmd1GxR5Jt
98UgtelxnQ6LU6a804HotCzdCtLC0FM7lChgLHKzzO0U9f4lN43pJ+hAARshpFex
1+PVGHuBa9wILZzSYMHG8oBfe/GpLxJG26F+vNqq0wtqah3i9wR32a5woKoQ4lMY
vLw8C3Mr+Yz/6wnPthX/KpqYIRsEbV1j5U1295J5qO5gJgDx61I4i4VZ076aUsQp
UOzt6sfD9+f63E8ETIUrXLcum+D4GzEcU4+W+sP+S7bL4kd13sk4qb1kJSVa9T4/
OWaSYnHPKrACdijJp6yIc3TRrMeOuOpinXYYEhnjSeUgqJGw1ISwLM2OQvPUsrOM
FbfJu2XkFNaJW5AaNrmcNTs6n9tLM/QUdFipdEjVtZ+GCOhJtXBVK87qpQybsCcu
fnCzJCifOHdZ2rxi/feTWIhZvlyYAAPibObuCPryLKafu0lJGiMos9lVEwGGSuAO
u5YcEv7INhWnH422+qRmYfZp94+6ouNwhGC7mwXCt6dvpBKzKnJa77KHBPZemxX/
B4UBpknl5uCKv+z33KC20nz4P0ZrexoR6Kp9YGZsguVLgRxyI9hCtIWRsKyx0s5R
kPUUwO3lTjx0BfkYpL7Wx1Hm18laRX8Ds35ioOPY9Ekuhwtv7h/4rQRTJ7HZQGuy
y8qHxs0cpFkq9rplUBJmJzkwpFNIbrWpOGu6DRUtUBFHF8MLLonCIQfGcx5vleGV
QVnjMIyeQx+8zeMr0Mb2ZnhcAz9Q9AJhIHlQ6OmbdQVIUcXAMY+RXGQSR6Gv3W1h
auEvYPFV1JGGQNrOXynlsaITGY5jtgfjHjhyJ1mfUGzH6XTT3fNZdIfr2vkfHjzz
ONcLm74NsEnTxcBvFJR/90wPyG1/dRwUhSJ5J7HuGDXTTt88b/k/Cx4RQJ2tX+Ri
Ott+rNLKapAOsiCZyf70FPIAFfRBU9OvY40YX7Ru7DqpjeFYI0OKTnoSBR6kPQnG
SiAcqJX6bqd0ZOcD2CzhtivCF8n13+vP8vIXSIYUYK9IHn/1TBR71wiLF7ZgAyUb
DGcHfjrjTr/24bVMI5X4CFbEMtkR8BeaELKwdnbzDBufPkby8KqB/1AfEAbXMPFP
5kkImUCDKe53BuTGJdXCDlaeF82BGhpDCzVFq62S5s8xJLYaAeiWTC+kj5sCZ9Xs
s5LK+dVyf4KIpo1PPQuiGfXUmB6Utj6oIVsLdirV1qzBXOmPsChOdZbSM0hCVIZF
OGpnMD8jb3eolAJBAJCqPtSSrWk++tLYvoyWJlZaP+Y9am5PmIqKasZW2UIUSXqV
m7WAT7nfrIgK6LcZN8VzKYVnFQ6B+8DdJIP/1BoUU42HJ5TpkPRZqmEoY2JNrNpe
J1hY8zWNS+AQBRsnJU1lidN4ozzxV2YruxS7BUMKggInaI/ciUw7vnuepadjYKCh
YPDkUQpMJP5rZOeODKa9DKrTzTFLQJQVcnsDm40lkyHRolk46ECcQIO7Kaf1M8vC
npur9BTpUxk7dwrsTbSVSQaFipQ0z4vtJZH8c6KSt8gTToTQeqbym7IhROX0eE/F
e9fIGN0wfcVixsHxPVubKjWlaka5n34nEkVKtzpevjd1gaGQ5v1INhTdDUGOHedw
naz3F2CWBKjYfSAAuzpQcz4bl+HXD+igQp8UsntQHTJtfnB+7XVor8C7Q/f2/V1+
T85F9IAM/I9STbQYjTfq+F5R22pY2ipuDwuPMOra5dhsZ8TIZIkMDIT3x+LFUfmL
3kLFvSWQJKJGZqaE7vHT0D40LsBu5XwvnamK2ZoINktHVMHMJwCU3SSaZ6a+/aTW
NEiVpA8PGLhnhk8zvtgB6uwgR0gqn0kEI2rvJQSlTezxvHzl8oGAazwc/0+HryZM
IN26AxLZdViaOLlLtqCOKTiXpnrvj2ZUSzSjRZi5bItlNGoPt3DxHtYbLU7QKc3U
tzmI2DTnQUY2RMO/VQFje/Amn9ZHpqG5tfKTaPaGtFxViU7QjWWqJdjZ6yXfKUcE
PiOisrsQ0/nyDS6dBFQdWe7P1NgMNoo1hcUmMCR/lS+8FkgyZXnLyTK3iyhgpR/i
O1Vqv2N9xJxnAVKrotfdxA==
`protect end_protected