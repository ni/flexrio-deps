`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 41760 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aUNorLKGzTZ27kyxtY/WKeVjx0eGuUvSSqqZKaYfxgZM
nbjRpjlgCxYgqhQw/Q/zfrpIsqd5qqGiMdxAQPutCIOUn0UB+fkjaTmKMLCIcTKj
1naUQou33gXhXQmizbNBxSigY3ctPuyH5yvopzz/hmev6WdQCtfzMtalgEPNZOJA
K8vvTh3CndRNK8XpNqYbAlCoBDIF357iMbp/MRim/MwWX1LHg4fZ38o/nd93VH6e
6WhUuaT2SX6LLBo542LT3U0GvMB5+TntV37zsuOko1QG88CNynxnCy1iRzGFRDSj
zMlfvcBxwtzzHwU9+iekCwH9tvuI45rIKXi5Wq7mpGq1kGVmxCfeYu/9aXaMI3ot
js2aJzb49gXtR09IAMo6NlK/GsaaK4xcwDTgmdguFSByh6c5RJGsR0gIZbWKK+Ak
SCH7LmZ8ONuWt8HUqogpGGduPMV7tb8YsQRth1+4d/WEFhHnris9wrqJyC52rCjf
11PhEuIHOgWJxGL4cSqy0RIyqN0ACnujvN4+CgqjduVQQQ9K/sXfQubokAIe8/uS
Htf/hrafMk0hYpPgGWsGtarpUHZztKljxqbJh36MecUbFhaY9UBgNKjy+dfRF0n9
qP/+SJyxBIt40T4tNNK0q0XCQoq9Iw3RKqlFgcT/Pz5je8RyyAkaPhJY9gks878Z
LJqpy0LL75xkoQCSlh0Pt8evkEDNsJTxtnDAtOMyLRN2pZQbswANUr+QOVZxzIok
ipPfv7+EdfhwdFJUJQpYRTgMspyWjJxLgJYWAoiv68oQ70rCC46gBQjqaLGSrDMJ
4l/DdMS3iPZseXIb6zyTo10hdvsEfMioQZ3P3zKEzMcup+Tla34iEPtjUaKG0Gpx
iBCcautbnU7qlP3kTpEqYabkM2qwR8uuJoE7sUOx4LJQVEXorpX3afS91M+Dmyvb
zo4lNG4m6eWAb6bY9UczBL0vYcUsH9ukQSHZvWGJiIMHtmHz1zcYR2ihi4YI/oRb
0POj/O96B5dDjGPXy6s45gNDJi+oLpOth6FNAOVsHhJwZV34VNii4Z32pQ7xb7+A
O6lWm6eBb1/5c+85z251pneiX4dO6Oa4EhNMZ/k4GoVgN2h2ogUvCHbNX7LNgT+p
eMvx3fVwHaJbg3Wb9IlRW6fGk0ZLVDI2RvLzCQ4L4nIhmMxqLn4uiXqIInmXWdrY
i/5pynGXHiUAJsx5Ox6wXHCpZOAz7NtFvYI3jcUzG/Kf41VEpBJw1MMz/jfJ2fVV
4pb6LOrnP+nPDY8FQZcc1A7z3fplaD3XXwr4c9Ot43a7BAHhPyDAW9yJt51QFlHN
VxbtYz18PD5TA7TJMQrWLsImyAECs3EzpathiH9D113gyD2CsoarwyE5vSVe6boH
7GRmvUydjovEWDzHnrinLSmodTjjPsW8lyWmtKQcXUNNfsjqmUi7U6Ex8zMM5Gip
mxAqWx1n+vFYRWporbhGlNByZ+4TB3cCByP+IgIGun0uG0ReUkBBIFSENkY5+2ta
RXJSPPhY79YgbRc8zSCIX2bLr4n5mIE9F9CSbbf1pWhru9QCd/7zUIPxIQ3n5bjD
Exyo0Q/GLVRKrTiJHHzxePO3yrs7r11WYOWqJHdSYFhr1LQWkkk6XBsazY0ZDO6/
vDgxwUAmKfn+AYQEyEYCW0wJuyiU4Vfs8pfllbfsvIB6e0NSEJ3HTLZaM6ylD0gr
7TNG2z9mfSu7nYq6UlpzldwqiuDTLiyOfwFu1RDtm6pXh9n2Y+9lwEedR82/00rO
QyC6d0Hd2tYZzLseipdyiDJNLx6CidIHqSbdVIizN9n5yDu2lbJcepdkQM91JMDk
npXMVuqSRgY61/M+G4Vo4PqycGP3cBJoAJvWYiBMpkC1CFfaH+PfWKhWvHi09Z8u
tjrLaudxXPigBANb2EKQhBsW70/jlS7w/2Q9UDkxhMNV307rYv+9g8ilumKFQQmJ
vFHfmlZkmo7q+PKXy6cx1aMWgMnsJGwF0UJXUbGLVjroD72wAQolziZH6HGsY9zK
Isa0JxMrlb74MLJh+nYv9DO/tUkb0yAcB5HShKrmwaR2q/6JP8OehyUoOj6PdAZ+
7RJwF2laWOU9rvME+GFppZc0G80k0FzPffvgHFcF1f2iCx801p/61O+Fm8CGGL/A
qvA9ZvAtkSQ3vJPU5Jzh5c4GCSsqRmfS+lJi8i7MdTNn7jyjJfwHm1vsOPwVKTF/
sj/+n77URYImGUl6UiuH+xEF0vT4tvcytFvF4i5mdLHVWQ8qNVt41zAZP7Ly8KJj
/rATIlRutTPPlgMqhhyeoXoP/bo5uDkdTFmNgza7tC718yexHTVIxNv4Mhuwf09M
uRyLVcvunnxlRW4zNXRq8f9v8Zwi3yIcg5iM0pbZlRmc50U2llT6gWuLH3owGN7T
Pm4jWTrIMuD0QAt8j2YfBvuG90YcBppRX4Fq4EaEuaQPzThVvWcOqE7ecp/Fsbgq
4Ar+7DtNYlW8zakpnFIuNp9SRNzwlujG28v9p8oVW1gpjIOVwmdxwJspmjD003iJ
QWNclDIiphYpuHQYBPUmn515jje/O9mm66/c429HltDenLc/tsECv3FvoMhe1TG1
JrecmTpJF55r9HSI6C+TROgVsfRlRs/y09/l9GVoNbG5cK/hjD8Am6DP4YXB6PKb
FtWs9u7wDbJpWSIVgk3x+9HGsY6rzW5JODC8WBVl/3keGjoVnJxCHnvOimELfrGV
knV0gkKQgBfdDYDeutjpBPZCAUAi4c8djqKLdFP7adEM7dUoGchEjUQ/5rnEt/va
/PGALP4w6HdYQzo8aATQhdjTbu2r+4x2afsXCpt1SpmLEIG5mMHs8ZZ4Pcvb3d4x
291ge0cRu5foCOFvnlz0rUBNKbFvGXW2zeL7MbDFKJvvG0buIktMufhP8Ri+ZrOs
QHCPldY0J73/1PYT2DdkoZUzVa3NLjtBhnrdfMvswo0dxKA3hlTeA+h/w3nlQo5a
a6xcRXtkAqhuEVf76VHaYx6olAqkC7GnzNURnWMgKrdAKbTfBTj7v6nRf0CsOP3O
xVB2cNUoetbZEYkjpQrjtWTY4bIFXM9MhkwNf3JWsLLuH+syyrDGhqBwVi0i9zp9
wbOYBtZ40TVUUtTjV7Fyk8Ccd6OUNiXbDvDEXLEELwR/88pxpOEimEtxmXQyTaT0
dGmA1b6+K4R+lP5aiy0XAzQiFORkJTyMtMCSNy7ZRB/3nPT0WrDadDSPFePP7CbJ
V9CgphS+jzdWRKLLGJ/UzgJ5j9qTho65UdA4B0ml3r7XBXcMBTD9cR0IbB8zpia5
Bd1uzeucLnwyhxjAgjRSeKDZm8G4wMEVSEGMTYsMVSCA/XGsrGl3bQ64Aypm5k8L
ZmEKOb7UK5QjmMhAmnDC82AlNAzfY2N1PQwR7RteG2XvDNNENLxzXC/wfDF6TA7i
YqJvZUWrxm/UGV5RbIT/Dj4kzzr2fYCmexPOmuvY427IOdaJVvIxYEikstNhiWSE
Rr6oKgOnYF38qo4lyGIRkiELSuyQL2lBgSxW8YwM3DYr+PMmmo4wvSDUVydC0SNU
7hZAVrdPb2M+fMXALc1TAKHP7nB2S52zcdbOaoLxVo/6wZ0tpkQoactlltmZb0pp
jCFbDZsDaC5VW/8yvSWrkaKhyemEaby9TZ+jFwUjBYhwNFVySN3yDf4c1afvzWW3
fcSnn2KdCYAKRMrf7BeM/7NsNeASQa1JHHyyYtwlv0Enzrl653SPgXO52xEL3edd
woaRgquVC/A3KrOn08iNuP0MCCI8cAh5k7LxpLp4vrt+H424rPX4zJGi05i4SR4c
4GPaewFOigD+79EUmtV5KK1uFtOMoNwh10bSQOWg5TRYKcP4CQkjEjPDbOOvNnFE
/l5/0Y+qkPuqZBz7rmUs7zp45HBQCKbmpmc+UWm/XW1IjGeXVHMBgRm17PGZdb/n
WuCXQd8BfocsQZeefCccjtrELdPX9jLR9e4Nbt4H4JOf+7fHYwsLJcH4f1tTkGsc
XDNMWLZZfaM0FcbpKp4JHHaW2zyMdFzjH7xzaXHIrmpvrdFDBU4SuDnGGJ+JFP2c
6t9TX5gPd5KSky54nxkOeu2dQjLu/qzIFPFdoRWqBG41vYLh6xxiW7W4l5Zz50LU
xQxrojcXWJ9bf0d1ja7pkNwcsp9uaSV9FmCigNErRtT6W/zi1Ch44O1HXAqoR6Od
7Db2CRbCjFf+APhRnmZlO1lvwOv5RWhqqju20Q1Ii64SIYWWHN9HJP0EsG6OOXqG
3hDgyLcvKiUYysjswbhrgrKa0TrlGEr6YIpsLCJaVPofI47WvIc1uhTXmgdy7G6w
zQ4L1IIWhqcskPEz27bs86xf9iWzF14jrjqx4IN/UVaOW9MaLkUkK3Gm9GR+LQN7
3rttECgWOmbP0T6efOi001b2vPcrcSjpGSxmD6M5PO03W3hP0tq+KGcPun5hICK1
CoWeG7vpcFAI8eDZ+w1QXXnSdKoxINGJcoMQwgi/KShttEuNbdHuywG3p/R+Ubt5
ZOzTZf01TOAVr9UO7CJ4OHvFC3q8f02dMrfEC5UI7jS+JaQNRm7BFpopRMDeDCW0
e0CzLDzzi093hBA1/t/G8NvzDcZ+kUwXeVTK9Uz41s3XvbSVVB7lbQPcoahvrC8+
nmMtN0tATXB1IuBbSK9pi3uO8C8H5N9p0FjZfWvnsS1J5HGJVOiMwgFKQtTvKgaN
tz6hGvrypKhfjuepjPMyL2JDHLODSvWRa6rFLRdJJuD1rYmZUAt5kqzh5dX48BHX
OPmNW48ihbcBL4acNHRvYjKhaIXn++OCjxiZkP7W24J6qqx9UIybvexz+eqnzOYH
41KQEuVMFFmX0ArhWvnw4Bn5q7kjHUZIi/cllAOi9du8ow3lKLXt+rOqyAPzvNqU
7pNeawfJBazYep40both6agfF+Au1c3GZpOc74IfHBScGPRX7SPTy+cllKmcLE1A
vTxi/NaB8UI2G/ktswz3QNTNwv61tzNt7gM/NTpZvJJNBMSNQRJuOUzJwxnkR6t/
iy2mgRuvjHpyoQPfIrQPypn9PbvUC+4K0KuHnJQPaDipy/gH2yL7Li2rcN2mTtcJ
QRC7+RYYb45oSGRppeVooM9z76w7wRa0+R6aBTVr6F5TQ6FwIgJXoShQIZcl1IXY
H6ofXsioIyDnWgwjRxlFm1AwCdEZqAcdncY1wPUAcXilnhLT1CwQIkxHh/9zDoq8
8jLxuaRL4i6/7BtdCatdBZQ/rYkJBKr0JfvVchBPgQclj2dJ16KSyFS4FnkCKUoS
RxPpbIXYwBLDoea/lNiCA9ahMBs3/J4rfKyC9FpMaXyFbrS3kLv/pwQq5V+sZ7OR
XELHu6pHBEWg588DXXZ2X4z5QAFtMHAaI7nSX7CGD2pxMd1px3Pslewurp1pYP6m
sVEe/hKblQdobelMmk+qQ+RZT+0HRYUnPmU+paTXC9heifOa25j17AEure8MOi2K
TANd/YA1n4Okd5m7KOkvuPIylZb3fECncVlwo/AT1Ur0JSzx644cWqo5EYbw5Ilh
VP48mw+6xC6bKfxRZZ+sLpSdkFu+6C58UGv1k23cqJE1jZstnEYfFQEXjkHn7NOh
85jwKm7o6zADTg/ps5xcaoXmMNXJ+3Pg13rLFeWS7uUf17nqxv+cOssuB8h9RUMM
9D4t/T91zmJ5z2Vt65ZLRi20aToPpxyh2UzMXEj8kJMOW/+BhQosdydyRdW3Tm4L
F0QKNpHxofaXthBk3DZWIL+PIxWgLPQJhEy7zWkp3XGDgMv/Od72VgbdJr6QPB9w
tCaNLpmGP4iI7P9XPtvzxCS3pIBGJPUqUFwH/+oz0We6YJiXrJzTi1F4f8MnqVfP
hM8HCdXNRYVPH9MZ7rZ5djFL/DdhiJp3V/vCGE8lFb21KUBKSP/dikNTHCynr5Pf
lNPkjd2Wp97HWE5E1BYU//D1CdDSmheO8NsFVMpJaC0GHz1FOxvK7gHa/j1lOFET
PP1X4aq7+FU7myF5CEU+crKA93lEtpfKGBTpQfTGIXCqpK/EkCoUtNDnELn3DN9h
2bz/m9kqLskQIBq61SSSEB9hDmXnkvlyB4VwPDjRL4cufZCWbYgGLs3atbIWw9iV
Jd2Ewkj8W52UVOEF3n+kUsXYzAekIfJ6FUMgScFPnMfZQ/BVx5jTa/B+nJ7Bh6h4
9UBWRtgSlIt5jOvy105uI8lngpl36QbbHiA4QAIuAcRA6zBcjF6NIolVpHaTFxJA
4IDIFNEykPAakgam8DoO+AWCpr/zoF+g1sNiXnkmHXOco77PtU3KBHI0ZcwrY+9X
U+ZlZvhIDXB3DssUbAo2OyUxarDrpiTvLRoM4XbzB7HiiG5vXRQqjEqaBWYImdRa
+qlR2ZOU6HEFSvrDYhGDHQWr+vqEim3dPLmmrR+4a/iFxub0NJlCDCQNsMdAN+Y7
fwmu07fqF6ZinG4Q0aMmsTTc0Y73ftzNUr1BFc/2t/Pl7b2OX9Gv/YDhvvAeYGLG
5TWJaae3ZDHaow0e6PsGN/cxTGZUG8QRbtShB7CZ3qBhXzi2ONCnS3rJUAtFPbrb
FIZ4/MV70UhNCqFLYpjBn1U8bdCzoauxT+XOKkAK47brWUr3oMPkGwrtbfQ7Yx8w
0hlnvBUYYYIRbgz1zyx188iaXabaFKqfVbSDymfwL3jkKDVtYH4Tv7pikfmDFuUy
S9HTgmA1IUWWaVr6toebI9j0cbCwYLkiTzbYueKuoSvgS5gYhotK1PmRjaUzTXFi
68/nYtj8DMMgo5OABZr+dqcibdKOF4a03DMV9Bpe+hBErceEeWsW8VkAzIxfpsg2
50P+FixSHYArdNNIxU2I44ogW14LRZqkvKJzVTWUqlYshZaSP2mvUV402RXeYeiP
2He5Yeg0B2wI5tGK/uzvkQ3DAM2+RcGRWTXq+FDFJ08/E2oDq3Xpr/S+AROFjMqQ
0VTNRpMWybJCtWnoaJZ6++90UIHKrejuzGJ4KzgdpHjJtu8mMR6CTPr3Q8claEfC
R+Fqa80Cbgc61hxe2T9GmQtDzuL5gptaXgXSIs9UjlLekVRZ226eMsWwAuE2Vqxs
jAmBwiV+mJHeYNBE5Zqm6eF9IfAgh7nCFMpT+g/tjG4Pobo645aYTTDYoMgCd8R7
caf+fdaJH1shzA1YRZrPz+GjwidtL+K6MZBHGQIuaPObReHj4qVTRHivNi6PTydx
YG5XElVWxCKrekZw7qJByrgzPX9IgXrSIn335ygImZBKHE+kBlRrA7TJPHJH0m2S
pc96RqUz3bs19k5Xtm9WFVuM1C0IujJloIgeBe7JEbCPzCb2XFsKKfGhkzc3tzMQ
F7mFfFusZEo6264RK0k3W3xP10qJMu+oUGcPcxmSqPtmMrzPaswtw+cp2LoPOgWG
39hN+Hf8eicGo4MQii5bBbE6RG4p0nGVkdj11JeqRZDLPdddjhxtQeDvK0A+NDyk
RIsthv+xrrJyVXuLl/3XsvEOPDFMMRqeKyf/nS2lTYTf+TB6/3aEnFI5juWmTfmG
rv/lU/TtMXY3yI7LjCfJFEtTJi+Q9cOIIgjyUn+EFk4R1q67J7SM2apLVljGT5N1
a8DfLt9XGTqcsU0r4VjnZ777FcK7DNce5tuiyLBLDkeI9O2v/qWUeMs0wzjS0JzX
eoFdpSU25rIMt9YKWLrh6PxqBX/JAWr7HhVQKIn4YhtE79cFbvGtosigZCP2MeKp
mmrh/rVYQCtC2dR7jXaZEWvAFZP0sqrx5ZL/dOudas/Jz6ErP5+0vIHmhzswBJ8O
0StX4Tnl+PXb33oYPTpb7Gn+eGFmDCmUWYN25ZhYStoS6ZwX4JWWHqE7deolYufn
O5XWKSzn+aRuL3+heM61UV7RZQQCbEHJW2UWuQroGkHwU9+EI36WA0zdkhJNtKcs
65i6rmltU7ROiENT+MHRsrynH6d+SMoMYDb47x1s1Pzcnfn+Ie26SjhNRfXJF+fL
tbe8+xZMtBVakadqpGHIH9WBWb8t8HipqTj5nRKem1SmlDDQCzoj99YDGzEH0Yna
ByFaVYTfGGnqmXnhfutHSh0824Kt5cTylw3U4yS2ag5SnPRMKhI61Bok+RN6qGpU
ic9ZZA1oetg/Bh5DyfsqU+BxyY+upm6bTTK35uYj9kk9Zb4R05g71MZ4i5+N4p1B
vEHnWp4fXPKg/5uZV7MOcG9HozbIunKgaOFexYAKq5CvelbMqkG9AGqQOqGa3UoZ
FTx9mBB9AYDzgG9mmwH3qRXKshPge3zpMlhlHBzD4bKt7Zk5XrHZ7BVAsKJWxAxo
WkwkyvZ5TZ5vG367U56/V271tRZhElSUTneoYdDsf34OCJ0NM0nlR41HHCGP0h8t
McbaEFaHqSj7snEfPxXZfHc5MhZE2VIor2tKhl7T6a6JeJJoyQ7LTNah0PYcBiLY
mF2Xsb+VfLUvIIVHnCkF7VbOShTLfvAFl7X6gADLpCgE3Dh16CSSToP41g4ct+b0
RLwcO1/Hnvban3JXyVARIz1NGhnnxpsx/6h5xwIfq2PFVzfa4/v1i8VfZrLvIdR7
8B+4fHABxKSlNvkistWOuItIXQDgAG82DQhLCcy84yG9fVH82Kaeu7D/GmVpJ0ZO
5zIaFZvOFpASVbX+FKi1eqiTcxiJDZfDDLymvQAhihks/VHbQD8yIS++4bNaSRmL
LHrl1uNh9NSkI4vG21YPG5icWempyZ+9N0yTwRNzDOtBvYfmRw4VBpaLNFvGyuvJ
++DEwqEmg18JmInRzJNjgb7CI2Cc2ZdU7QmwR5hNz7kmDH5+69kERqDCfRWdEc3G
VNQCakHs3cQbgjnQXLpn9Kn0OtCJcBP8iRPPjf+uhZysUvVIPPZBDWRH0Mb1W8NW
/fZ585J5bncumySRimOCR142Yd52TjsUTDvcJXURei/OEKOjn+AASkZTDTNVoJa2
bEbC/I9FUc8qC5+c0KrYKQltGrV6K6SjrpEcQVGOvo0hZYTlWB1mO2Ar7J6aX4K2
V73tAAptWLN7jL5NBIFHpxl5NI6rChGOs1/P/FF6uuhSqknLGN7kU0BpFHp8e4gz
T7KRwbbwMteWoxyjdNgeZ5/wU5R23ef093ksH1VL7ZdHl/udMCqgXkJiAM6yTVuI
JINmxS2p+AkxFMaGakWnXbrKpQlVnGmMDAGP45WcMLH8Eglu5X9Qbv9UN6CvCTmp
hJqSpIb9iRKoGl26P7LjWmbaZ0V3Zno8RUCofwO4RrDvtiLyAM49CX159CNnWTbU
+I1S6+cfIeM3h7j1JQ7Xi4sOKdUCHATsPSPkJ+7HcIKrwaWCB5sX8lkQVPHkIXRd
ikdoeTdrhH1ZNByMf+pC4uJJ0uleW9WW8uaDtNhuEHUH0vhb+3sysB1jG//Ri3G5
S3ylkPs6eZfyG+yOFWHWUUUF0Xg1H98DTClas746DQZijkVRYLQrBaygt6wBn2Hg
AzlYvvv5IvP5HEUWhhQaklkDAJKiZyutswxpkJhG82g7lDVNkVp7JA0AlViAJAQc
zj4Yuy9UwSYYfYkyRV6BWvquV/U6xna76CAGOSr5eTSV2LBiqSG9SljMZY33Fc/F
kbfFwweLWmRdfgrCvTgOXlREkYswmWT6r7jgSHgtLnnsiV+yvttD72dWMhA7gkrW
GTrl9n7/uIrNZiZVsq+/ncDKoGu5RRgyxcCwRsuUmqT+JofR2mjiMwVJYkZ9P8r7
ihTK4X8tYeM0+fh6Mdq1h9KIW0nq5yHqRZqa9gY0zfT9xV9/93+JbK6irCQ8WYVn
CvCmOloZzaXWI9djk3UgGJv/F1TnZuXgTER/GxjUtaT7v1bEmEBB6zpfDBorpsB2
rU1OEw2vFSo9CvEtu67A07N185UfYDExvwS6B4yfXe5ZUKugX5tZ+tt+IOS1GJ1H
sHCaZTX6QZiG8M8qWHFAOXMlFt9h0sgT4q+OqpACysjxZlULmxlwInS4U+o/XDQo
bDV+O/LPqHVM6x+uopZYcvO7jQ1WGFcViTYmDflUQSbZ1voD/mqNcGnOG/ZW1kR7
ajOQuTMn7J8AIPouO6kmYl3bg1oXW7N0o+e/M547YCJCvo8n/DWTdpMnjBUtVMsy
cmCpYO9kp0zzzqjMz2NGzIXEqNbNM4rqicHB2LC+zKV0Js+78Lp51EwJug9PMjR7
uYPX/2GAR6KXrNRcXdS+rbOEgEXldhh8L5C3x0cTaSkIU4Kx+NMTq4zLPM2FVesg
T/ak/VnQXCi34kLVILR8m1lz/ayQ97kuCg3tFgWKsjSNseG1gEFNPY0rBzxXHi9u
9unPVZWY20vnwCZw1bMJa/CkpumSWNYTvXG5R4g3rWlPkS5jaqSkCljixu4clslV
gfDmGXQ4neLPxVRsMws9hzzScBuxgytj8mhi9BeSsjEGUslww9cqjeY5pc14c9jh
LD4wTPqOqqkrM8SYSFnBl33ucBAqiWYPe8ZNm+pdmxBlD9G+K/mJ4rgCPC5ndiBC
XWycXc0Ubr9FbnZu0iop9TyZRfI+HloFlKn920CIJPICZCFA2yBYtPcUUw//jn0z
KkKS0neBSXJ4djIiF7QIOFAsCfni0I+aXN6+y2WVvhNGyXzmL/WLmdsTQ16Zy4rX
W4W58BCV9udyeupKkLVpSXE6R+14ZsyAjNvxWxGmzkGCLFVy7/s1Nr+lGEbBSTzF
Nr7S/0G8G/h0MBDPf72pku9OKm+B8lEnbvXSifZcb4D1KOCws63XSCYiMI3jGqqV
rVWAnkKJvqd+qqY8/HRL5m6zbvq5IkyZaxqNchO3uhQLxYpj8YBFLSf5W6+7jcKV
wDlOj3bUM0zh3JLstZDgx9fH6qFTpgcJIw3a3/t8g+1cKlI72Bd0KeQ+ds6NkdhC
jBT9CepnUYfmA3aNWEg6hJUdOExPtY+rGC6XbRZ01jb4ko2ZHFDtFDA8rf0pVjej
fq84iIr/sApO/8QctI3O4WQTEqw177JiWdT1r6Yq1OlFLSuMkJj1GPvGmWOFVk+n
z2YKCLsmAfvpLqheOMizm9P7UMlOXl7nZcCXU2W5uSQdRE7Obd4kBKsa8fAVTKh9
z7UOMGWszpCsl7iUkSiNgFcBx7Opjpian8Ii3SjbiFiS+X0ZRO++zIRxTHEpENXp
n3cKxwXeEv/UIQKHs/lUfbufMwV1bJpvLuStPOsAj6zBXH1PElfKd0n7cP448sC9
yYCdDYFn1oVioRyKHq0ZyZd2Tzyc1plXRHo5EfljVXU0/mi+8RTXIgYkB0luspmC
Mcxu8kionHfI8AUfH1T90YgQ7lIfsMJWBGjnQqTJo36p2MR1lRhjCMR9xG6EPzUJ
qCyVWBphLVlvyINWwt72QvvyLVRmgRFVrm+z8uqomTO9rgmEvDHYVQ+qpS5AnNnW
gp8xQO7kN61txmGqDfeN+O54EYgwUolTUtx4iyU4boqa8JrWb7XgyEbCOz+4R+Dg
hCL0pp3dHm7t4fmoWFk/XAFSmHENMG5HOBol56tKkg8EosQTsxTp5eh2RhX0qy/k
buE5NWpq659JAe80L6Fw++ZvbffrLkDqeEDQE3yO75WssZuCCgn/oVALNszZ30D7
iKkTKNAk6qPeOYSceQHQTsh85EkPZM8NJ45SWJrG95U0waPX2waGNGLgrKu/gY4T
+C3SDGlepCoEJFT+T7ckutd343IAJwZHUDyArP1bHyJWViU2kGPsonhYWd4lqwOL
Asea8sUrQ16tOsjRMvW33pqb+R5ZzEdw8czf2bq56U5RNoT7/O/yLk6x8h1PGP7V
xeRnmm7GaGSLB+IFEC4AyphHpXabm5rDXkWfngkgHeYt1l9hO0txxMcoeUF67ATe
llqbvCRQ/tnx7DehFq9sKtStCt3Yfz3Gh7RkHbWm2Qyyk0lSWBgZu0LiQF12D24w
6CAgkrW3BSQWkk43JS9ynwRDkR5PaPtxc99WqSKCyrXlNAApK5txOWbb3biHM1qU
Dv36aEHVPqXhmdwr/kowMXA74xRDpcJ8xZbgC1vE2kM5H6EQv33tPrjcco59zHMW
NWB55eBQmzz3tYJQX2RFUzAnJVLp1gZcf3iKVr8wVnvpsbhnrG3FD8hkBUGGBq1j
0t077xSBW57u8Uw30wgPFPWIn28wGB7mc1AydxIDtyzc/UsaB+kVdCg0OBa49YCY
0ZBmvPQ0mk53jVpDurHpu4vjln8hoN/54F8y0VaCJurVtmp8Vl3jp9kSitMpc5KQ
02qAxDa2fXui6wlerz+Kcbm5T0vnUZw1b75TuOyd/BFHfnJL6HvWoj6XzqKUG2s9
uLL0/Xl4H4EZA39oam0y3dTc3yqwaSpmOK20hRlEnInWm51HyOKppQUe4HzcBqqF
ZI3RYDSw72wPbQncg5B8IRztYHseGH7Qpm9RpxFBMPJSN2Edg7XjnylgtHxOzQAY
hzBmylsUrbSfbwoxPkDNJvwDfM6T+JJUfT+04KQ43WCOzn1E7GE50iN5b7oJejvh
N3/9R6EHtXe2xqITCTVPr7jDK0CCvWvBhtovXxHDvd3wF7wkGTVYO8BsHL8hedop
Nmsxm2kH8CvPhxc9/Ldg9tXxuTfrWje56TEyy598DLIh5YAXnGvc4vO+nH2Kg/Fp
dGVlV+Ntocfx0uOftqst0Pwj8gyB1tgLB/jFYDIYBJ8zs73guvQQINyw3JD4tGuO
XihTdKfuzW2KcQ9bf8TYSt7fHT6VOE2TOmS6r6m99zpmEgV9Egufjzn6w8S65Izr
A9imjGAf1yFFgmpcWJGO8vL4ezU/UTxL4QCzhfTAJ0+TWHLanNcYYu0d5QfyMJyJ
IZh5GdUelhvv7yjPZLsk73UP0gx1YhTxowtbHgfgxWWnLDYV8ODKKIZnxLwrVWPE
JlHuUfTlbnLRAznNYwYA230MfYKP3lH6BM/wJ3kKNCg3ETVNX5bveJX7XUZPJjfk
C/qmGH4BInpROAkmhD55T1feHSTlVBQROiZt6VLV3ZtEy5uT01orVtj/DULv7S+W
YpR8DhAo+nk/tCtGnVFI8hJfo8ARkfR0e7Hh3FlsZFeFGUkA+eaq8nWtxufw/iyG
q4k51wfcAtgBInJCWH/afOSfghF1baaGLpP/yrYrYNp70iZtXbyY4SVknBqQYzlG
BiqJWuZPUk31e2dfvMQlSrg3tKsoVCGJuB1cafrTdrWv4NHklObPbLkCQpC2joCA
t5hwLR5HgHT27zJlHssBAeie3NDTTz37EX2S70IZGvF9j+Qo97Nk1/b52a20zIUz
nXR421iBfa1KGOE42w3UjznX+96INpFYoyTXafT07qU03vj/wn/M3EL+ypscYZI2
NOkOgYVCVuPtVHbGzqNM/hl1i6aO7mpDYFVESpU1jz9fLOsELunTG/xf1qgc5Um0
A8MFuL8CG8JGV2TwnBgmeQRKZ+0DWdzPda5O2YZdnhmRgkAdCXmmqdvZYLRoEHj8
sx7wrGwm+Z+oCDcoxdqNISK8kvfYpr/DbBGZJgWEQikH4sLRlvfmvko9FGd3SJbZ
zaYPr9obQfYsTsTfTvIBUzWsPgypFoBcSNefUe5c7e2ZXQyhJuwjIQIlq3SsmnND
ggrMzhloqAEaJGEWA2UFKB2c7ZD3EKHeHzWyU2Dn/8cYNlLxGZ9uNtV6MecolbM+
MCjGugghsJ6kPR9JVna/t7FlHdeegCbtFTtBPsXJuB32AzzI43aYntwPwBa9sFza
Rv2NdT9p2GTTou+F3dpR+lr6C4qXgWBuJcC8e4cztEu5qKr4XU/rJdbpjtyu9w1T
H0WJoMWU+ZR+lUSZbkt2hM7x6kfBrRsFhT8Ma7DF6Mo1IXjCIvcQQdBuXTURc4Mo
BXegAX2xym+4hIL7tyG4LudzoYlnL0t6A/lO1g1WkHxPUzFokvZWy9S6FDg+KQrl
ZkJ+BWZ8b79ndPW3ituG8IyCle6kugxj9ERk5EgjIf+GUvOE1roUb/TJC/Zgyhno
xSkeR5zQwWvtooAY8hMX47PBA5/IAzA8Q/gT4pbaDqfl4QOtzVBAxfXg1gzUJ9vH
Q9PuRoGHsA0OuRuscQoK+OqVQC1kxLqwKeichTeuQGzxHWWI8KMXAkSv9MCguPip
cqv0fgrGwwfSDrIpqpsovtuSObGUTHeJLA3x/kOjyCus1mQSnpT6xF66gfEahn00
792bHcV0cssR7LfVUJ7P3ErMqtHP2/4ck5DegE7iX4OiuPuMcmfdWLK1J3ovTnYw
JQaMSp02WflKSb6W2pRO/cP9fYbYaGMLMoUbgtN4S1pxtFTxJxjgMsQjcCzHTIG7
UW952dOS8wvjELK5N5Rj9Ls0+mjuCSMZY//EDvlreY1CfwWLByVutwYYwk8hQdgF
2X7NONn/pqG0KFfhZoWfVfw3tOMpvRVc1sPUMcgwHFly1cUrUbgaYCcCGknWKa0x
ugv+y6TiYmFpmQhbp1zJsGGat0F6PP+ZN7v8WWP8eOhKM3P45y6wMIs1bJDn7bzB
m4DP6zNvdNQt5MoQ2WeGAZTJhfPx1AEa4hcWm9cyT5z2IFGzOo6SHFuMWdTG9mMb
TajbXwKoajCerlxACpHH07dKvMVZSULCY8WX8ZjA46QpfaDNsX5ury8ouNjx29qf
X57tBJYZQ0w3xyjOrrrQ+xWWc14PjbIUw4oT1pzLh8wmUvLNQnN+4yFZFmN9ceBT
RCVQSqH6ycDBaBvcQHd9j9iRVcvnCwxaGWwFXHp0RN1L1QA/06B2sgk+yVrxQiIC
Am+8WJ0V+IT4x/zr/7n601PXJHpu+DYb7aivNLCsmv1a8yrEwJ+puFS5sJNQ3PpH
VmvXuC9kQqMJg1uURhN1szCcRKJ+5IrnLt7jO/EfQM9QdCBNMUe6VuWQr6rFUDED
fvpUUpow19JpsMv4PzWX+binE4j2gCV2aDCjMHrSiibr4gjwp/SNtuKqnRY4/Rpc
XR69NcFKJJOehJzGSfxpxXlQLYpFElgOsJku/HZPNkmEe159NgS4A9XVLlgOlF/d
OQnnkWFlK0PysQPAevw39/1AqZwzBnSIDAPDtXPVKCt0jTkuYanZrv7T8KWUt5oN
B9WKTKGgOKfbPMKTlm1wIWhtHlObjBh1IjG/yWJ8nbjCUXwBncfip08Ooh3PgKSK
Cfr9VdjGyARP6RMromsfwLaoQu+hbkqLCqGXRv2y4q6y3jxxv1EG1RvC8PSw7yge
P7R/lGggiRUlG7sgli29xJOdnX1AuLNiMfgUXDGkce+2IR08co+l1lmkJAbwOOGO
fcNk5G9coxcnEZ6u99O8F6orWMdJFIUDHFl1BgRrflnpBdKk+EQ5OBlKqXLTn6id
YMzmCpZ6skIAqbBQihie26ZqfKBuXoTyJEQMQw3EDLJCdVLomLCOPv0cnqaDzG18
iVF8QD/KGDnpayD42loZpdDUsnllERL7xXwAm2trq55rb0w/XY3v34nyQg1JUE6u
cFHdKxkfPW0Wv3waxsGxYkM2Y2LnNX6ExWIYmB+5swF4PH29lXQw/3UtvhT4qHdo
xROsJdoJWuoPTh0E0DE1DBzPFc8L86eorsOGN2ftHOF1fPkKkl73co/sZdr2Jjqz
4ZjotOIgftgpSHwWvoo477UcippE37aSD3ppbf9qyGi1gylzmcrXOOhPHwwVe3s9
VavP8VAPj+cdZss6gUr44UGNiGbV/6ihnZAvLh0OJs60nOlM6pYKej3wNIAe9+1b
hPKMhN1Hnlhie+dtBnejB1+3zjVtOxKns0ZxtuMPoVNqt/BqP+kFJE8fnf5fJhNW
oq+xOdtf4LmndMe7X8GWDzhQPMT539CC6NKujHotp3aGnNd3nFI3r7xlNGejYvzo
XWGf94eB6m97az4byF3jOT0scZpJGvf9JT0MY5CaV9cvDjfhrLxeqKhsGd9HaXoY
OOYuA6Dw7DsqzRIirPbKkQMs4b/FqSpxd/ppcAoKkrtxe85ZNqw0evg3uc56+QUH
lABkFquInDX0uV5lb37shsOf2D+p0Q9v3Jm6hm6tw4Xh6Sq7MrgR6yceoa2EOb1B
wDUJt1C1Q2w2OqgpbqTAp15MNLPFpepulMJlMd7N9QascQx4gGJVGNbi5LN2w/7J
hKkdTv2oB6K8X5CWB7IvE+8XBHDCJZ7/MkjFf2dNgV6ncOucqLq+NyyB5nJ1+ovx
/GhmKXy8wbNXtEPczf4LZEtR2LuzYpbSpqicJj+s4yqtfEAfOZTpsqpDWFIIz1qu
PLG+nutEGhDuX41CZaDPx/U+/ZJcPMbaYJyi3bepLCoHWBlArpFsYSx7yK3s9vL2
vIaBiGTTgU8wwycVV1ANqBcbXzcbe2ZX0RuPsOX0hwWW7loN+IJ+QBjrWmRY4qoD
PGsi1V89X5MvKao1cXUQ3+qKq1ISqS95qq6S3p0ZpezDBuSzqjmVz4j628AS9Fsw
q7c+lfrbdcTI127bJlJ6oI1D4xNiI6uUChHpQeKvlBZA5Wb6EcQsrdE6xWnQdHpS
aF+S4hFWGTvKg6dlNfVoMPs+PkcffEWKmyqn+aLEPiscrVRod9V2mhIQr4JynaB3
gUrtR1+Vn0Zr238il9eNE95J9ci+QbCZRWWznMiLJGNZFvJwA5/+8PwfHRcLH9ae
ZKqa7rf4gjqYYBNy7TxOUSUvJsFIOrA+WupC/PP4kB0imYowTn4/dTxX9PaYcqqV
+e3uG/Kj3JIaqkzOEk8EdIjQBde2Dc145zzixJex1mq/OQEsvTdY2sy7ft+H6W/J
hME7pqVKPStjBtOFIipwCusX2rbZLGrmj5xGc+gV1h0gEmkzzpnHX0ael+nZKCNw
Pv9FglC12Zlsvc7+gCTPiwj8hu7h6e8WqxaimPSzmq69N812ICr8TEh2+KAnVOSM
qI0xR6YfX74CCjdi1FEA7doXW7ZZKlkRNqO7Bz33YZaLLcydfdFVQp6EK/sMed4y
8rJtUa8DcmF6uC0dCbo/Ifd5rc0x2APcI/kmLG/ASzJP0z0njaBGsz5wE/Lugu33
iy3rm8+XKlg3e178kJ7DMZX4Dt2RaXoFJa6P++m4Sr6CwRrzS9S6JhrYVb/OHD6u
4F19va4pGam/H+GtfoSABkeZLwvwdpyaxCVBkl2AUZCtU3++oNjxYiIIpxWJ05Vw
JExZDHhMUKkRT8z6v6yOvEh5AZbU+l08Dx0fHF9E/LW/QQj8YNoQKNWH7LqWnn37
gNy2n5xl/njm/58a+AXMwLYCNsREV+CmvfYBImd4vluxVfbOi89Gd8JyK+xPTwaA
TeNNzrouY02Izh14/Ibo3tVXwVcRygCADOOxkaxqZF1iqMk5nq447OyPGwbSy9u8
QmIEjNJ++oXQ9OHK0EsQIGUkFHpx7oQpUfy/DhAqpi3D7vTX/eF/iHdtCkPtfKnV
6zd5xIhdR/Fx06AXOHLWRloHMirt1WlIubMATQbJcC+ilmnBFOrvG/4w63yPEt0g
Zle0qtrYUADWD+zAjbJn4sqImJ1ERShQqyKkYNQ+jhW3YB++tP5NO0C43TlZYdKh
sfmnr2Nn/AihV/KuvfR9fmuuu0BoFfQxEhOUa4PoqN9jD3NYvGEDeZFI7ahYtM9x
/DGcaRJY3+U8WrTJ5ZIz2cu/HOq9S44Zpi9xJNlIiF5Pg9KTwqDCiHpA506XsZKf
LuXzgYw0OKtJXNToDulM3mphurLPVRT9mx2HWS7YReAxB1mcDqUrxIa95wjHJg2x
Q8RDxx6OofkLfl2CEU96ZgMvpo4Vm5PQ7zmYHTtUOI+gFqDr4NRfYy9a5u2QwPFC
eYfiEKRvdi72dFO97pa+CCmMST5mdLzbpGZKU/Hjylo6I7owAwiOOKp4HhAPnAZL
9XkL4PfWjCBVHWmaZueJ9faoDN2qR8i+hYsdGf9H5qPireH5UaB4CmBl/ItTaQB2
zYtGsgr7LJvtu1sCfgUjniyWuZZOKX9sbY7fjy7zBOg3zXLSe6XN8lM4Lp0P45I0
f28F0v9+84sNZFGF11s3Dvxc7T+JVeHIq1+e/iRVWUy4QX6wKY+ERFg29I5Dzhz4
aPs2D9BYCGDbm6gpUpvqAmRLiqQpY0/yIBTqPsGJz/nY8ppZ+qVSaMLYtN3VuNN2
ETt9MhSmvcChle7BjD4gYrZ3WjytDEFVECqlFdUT/VJr9C7Hm0TwD1kdxzvZikx9
3murUJIw6gDlSN6fZZRO6kl7ZvZdYLX+Pj9qOBvVpvTQr+AOsT1BoCRF6ek2686H
ujYxFlJndokDUgjFAhsyeML+XF1NuPkO0pBeW8q3ffUtEUfdQV3sXpgU6qsq99eA
URxeeWfoor8u707mMyLervhQmYQKYRFWjpD1oRUdWW9tmmzU8v0XbbNIJsZ4cSI0
/iTX+e8eDJ5xr+CyLuWQ3Ml4Y5DD4jN8ifKPQEPgeabEAy0VBIqsH7mAspDsenK4
kN17fBkFCp8tjZ5T4Di+lrmyfK0qGDtNB3w5HtsbnlZwxjKzS3/tzNRtcFkZgE40
oug5DJVur4g81B6oJMJ6qc2YoSB2PYs3m8VZfO1MO0YcGaPpjXPQ0eHylruT0zdL
mg6kCrshIy8r0XdGYGbDznEw6aeemxBXktged5NUiLZToby9zAawXXJukV3XMqcl
Ig2alnWcWK/N8KRtTyhY9jfBJ7o3yWgKrWqOHnnsueBrd/9NypOa0mdk3gXhzjOn
ZHeA5/cgo9RuqWeI0CpF7UBeDTeABX43PVCOXimyBoELYpAa9N5gMdockAfQB4uj
+wiTUl3gOkT/IhepXIZ7Eki7tIcq82SXp892MKd7YeX0zYNBV3ZHJL8SdBDW8AEa
bS0iP/jCiJXEJOWhm0SypACzz5y+eEHMtsqUhmA4bcbk+3VBCSmskHQECxbeaXwf
4olEi094c8jC/q+N3BxJWvCHQDNK68X80YFRQCgRg/NOJuIEE+rD4NO0EdfXyeJt
Rg3fumZXY81/vZ42GavEJeELhwoqnTzfPz8buv0/y9QYEGVkmgbhNayAaEawwyrR
1p456K+it/FKBIntlxKrY9RWJKVpNExFzagV9EuaJNCos/P2D0970pULM0gsM5MC
jYFqb2aUqp70L4L7RiWFXWOoAb7lKAU0IbnyDjFY2FDulRrPomkpgV2RG6iT+mcc
gzH0SzZr/P0s0BCO0Relw1p8J1Vs3Wa/KFDuZfPcJmg8L8IIWGW9Cnc0vVgqnsCq
nyY8HUe1j4XAJr4zrcdcLa6AjjbUEe9GJIU/VQHTPRIqWJ0qKR+K3cxGnxRJyP6X
K5g3hCIXqN/rMlgoDuD5CoVXA+mtGuVBj+qcPZaz28RYYxHMjgCu57hUTkqiCsn1
R4v/xGNxvXbZqRqa4SPVlzOcIDwvFU2zFn5uUBoO1uYGO0lhWxpM/Ub5NMWvPHW2
frNObCm9+MQiDgKHEZCn7FtbSsj6mFlF9XYIexS+7plncb8bnyZeQk13e961zwD/
s5RIdpkUXTa7zRfqfKTeY6JlWS+N1drhSa6FeqjQEVz3q0fBs6wctfZ7yOFgihoE
1x+n4nVO98Bl6xisL4G74nhGOtjG2M3lyWM7IHZZU228MKnQPyacVcIrJ+/42ALi
RywLhiJ2B0mtRQoHQs4rv0xHstDKNlEbIpegx5HKrmypYoImVmpaQJaEL8X7jwRc
JTPoZn4QZZwJSqw/rBwVy+VQKNTz79ywgrauBwg4AtzymXrcvFBSrbAtP6I9aBV8
9Nn+uTNvxguLgpKpOkSBST0xKDeWN+JVh8kWdAasTxiYC5070LTJLFOBQ6QiQIz0
E2lDMIrcnYKjbK3TS9SzCEIG9ychRJb5fQWQrVMgQvlFJHoDL/0QSxPTxhHn6vwG
aMMCZ1lf3HlZpFNbu/E2cGtDnJm3habd5SrdHQ/13HZLNLJBc0xjoLjf4W52MJKm
+5LO2HW7rwmw2hXl3M5l9fyYlgfTmzEwyAvsWSgy0SEI/bDlduCglODgEEXfrrIv
0uJNstDxoKJq/ysaSRQolXbcOGsZitE+ESRd+B5dvxeBm4parOBHfIySPyeznf0t
Bw4OGG6uwGn1Ks/SgQpyI2t6uqPzEUKLEvO2745Zlx12oWO6xtNhXkFuJZfls6nP
btfSM38ycqwX1BarIdWYbNEfckQU6RabeuZRY5Lbnc64r+wrzyDnobpowbxEzJaA
EeAnMWLOs7zzNB5CK9ER6EqVqgyiKDjGXKAtojzg1EYBHqpZWtrlxBPE0NphPHWM
+lIEkpQxeMTwr7LIr29PNbHK+/iXElGyvrC3bYctXNHX+bGlO12nS1RR9GpeobZL
lPb8EGSqgJWSyVuenCVYbOm/paTxk/2pTYN/wVvreQjo5/I/+584IjaCt5yjF/DO
jRDb20jT/J58fFm3sJ38VhTE+IsCqWSAFqIhquT9A2LzntiZMOXh29hKxvQIbg6X
WO4mgBD4KgQG+ZfXYM2fi66ro6L9DwZDzijE8uCTbjbwuzKbgNokTWojuCcv5AI7
cuHC+Hsb7wmi5o9KAVUXze4Aq7ZHtopwxOhgudrCegyvTtpK1Rllx0Biy7xMPnje
GwerM8TSZodz4Fluc+wKYsaSj59/AlWRxgkcnTE6h82tJbOzuIz8Nbc73UmfEX22
c028a8hbvtKGI8bhIyivGmEB52v0ECEDipijvMdR57Xl9p3GCt0FTvfmT50Gk9Hi
+WaMnykMt/GPGTQ9/HjvuWudvjYfTnmKdtgJVBbfAsQj7QM/EtQvdymUK3BTBT+Q
/CDTmvtPr/XHVW0Qhjahbi1NzilS2ZlQxk+6kkSGhAqz1QTvVd3Hx3Cf8T21VscC
XfouXNNhkavbTB9NJQ23rnS904ixapwIodHS2Q0AH2kTUwxv1V2Pd1aQEQz+8xg1
cuEs9ccCMGQNDKxkDdQQlo6LbRL2ZFbD5jpCuHSQEOHhgqlivij6edHJtN6HvXKq
c96UirfCbGikjgLx/Gd72GBSId6TYojQt3ncgguFAkMcalPVGZVqBbKN/RcT53Gv
Jt/yICD2oDmRlwmJFzOnCXRnYF6LMS1sa1eD8O4YspmDFictdZ6srMKHxBc9MlTq
EfyuHTNEjLUgHBZQ5uIbVIhzPWInez3/TIXV13Gp3Blq+sByjjOkWrY/nZ4aNGYO
rloxkG71XwVPG3ATIPdVu4KfeTSEELfXBhkF7bNSJaQq1tPbR2BVoqAYRcmU8Ai2
6JCT8JYLkxy6JGyGm9bvp5UNS5tp+nxBsRYyFEannY235Fr0ZisM6iAvjl6k5vC0
nMom5IZj1qJlrqcP7ZFUvd756xZA2cdq9s0A1WiGIQXR8L4mPgrhW9zKG17r68GO
l9dy42flltDRg89DDSpiZWGlRIYS96TKiC8bnFWsuOwVMgq2lA+bKKRwZ+TPyA6l
l523d9FhRZEaDSALgdxsIhCPOcUQ1/1NO5ARg+RSsezQy4gfpl4TJLmqvO+OQDg+
rTVirrELqDBGloN+CfsyO3kFVSbS0JkZWaDSGjgZ5TVGZSQ7t1nRj/FJDGUFd6+7
pKdymUnjrXsuc5lrb4QX65cQaFXECGJWBepKL5MYJfPYs252clJuqfCow/xkobUi
Ia1J1s+cDIU6zgGTfmoQf2Yv/iG0LBmQW+pxPQy1hwriO0OsLLRFGV5Lwrbx9SOC
1ViYdlaKiZykUpVBI5xdRzmlY2NQqD34RhE0ZKQai5TZqz6myEvbCoc2sV8MlgFc
tEpJY0OY/A3br7024jsE66mg6d7nspTgZ1ldNS6uROSzX/CTIJ1L2h7K3N6AChlk
e+nu2RGI4ZahCwroLe8Do8Txr0X7HtGKSsUEXrqMTQqKe4N0DB9EYK4DtLWXbC2U
W15kYcDA2pIMDC/SkE3qcgLxWzHey0F8HpJUsfhAKDjm73jgjB5zWUktLUkYr/3J
65Sbowcp2u7Jb9zpeFEBd/W1e4fRzHFzK5qxgi0TJu2hPZ9etLwGc3N9b6Dn1spG
Zb5pNMHQ40IRsszhIs5dkpMPwcnBpCUAXVXim9lmFg9JYiP/T3ImB+c4SGan5QxC
7vOFUGOLdzp0cNtYrq3Rp2qsyJIqMHvs1+dhKowj8Nu5g1jo5/+1bFUlNiSnGy87
Rq4GHYT4HUz5SqQgqqRl0+Sx3uVt33y0OtkC2rEgQG0mZVqmGGisKr3omwJo3gpt
Do6JezIGFTfmzBcnKgvtJsZV5VAaXNzRd+zufNtWwWWCV5kmS1TXqvzZNP+U8g+/
tvKGiqLpOwajbeseXJtLerTrOfQhOjc1YcBWaeuHkHWDdRSeJYaPy5GCC+iboCEx
GEFCh3+5ANqjvjkQC6P46TmhSqKy45WCw73xo89V0O7L5EhWKIBl3qc4RkLpz3o/
U0THXvSJyoDVT5Kf347lXjdkfARbow6bdLATknqS2+LTL5HIz2/R8St/9s7tKjY+
CLjGPZtw/OqIbp6cMBJBnPS33JuNKfSEE5EpYOJg/8TxO8W1Gv/J27gx8vI2JBSJ
xstTY4SjZyhH1QA+G+LncoqkJQrGpFrblfXgoJdYPKOlAB4J7fkJ/UE9e4frvANc
TUCloCnM5vt7G5rDOwRcoZLTOBvaN5K9VApl30kd0lIHodtOwx13ipJXmCz3eJ1B
7lQVvfEuEIyYMWcO7Pp+a8zTGldFhcWAVzBJvD0bvM5i00WR8aq8GlZwQC94+fP2
z3eOodmgCOFR+e2dIdp3MLvVNhQsDtEjGZVX7oBVz+RLhOC0cBHbQvzg+wrU3GPL
gpVvbBIo4rGVCxuCIZIYOMuCJ3Ns9d/3604v1qXsdPEFLezCLOuUpJwJuL4vxl7t
COuzGDT4XDgugLD0kkSyMQ85ezCLWHOV75Z2KSp1YhmKc6n6PFMe93GFg6oFiWfm
cCCNiZ8tklGesB9jGC48dJnzaNtufv+4qbC7pxIxz3uHyKakZ8QncRIemnXCoCbA
ufe0+fKcMrldyWP/cXtlgqlV1ErfEVJXaImKXKjfq7hSoZeDggb8ikEiIye/d0CN
QKxixzCbmIN49lmFhCsSW8oYLWUTuboYtJPzEeSWjQ2o35s/gn7SrEgp7HpYIjgC
TtT2Ot/IotsNjg5/jLVJkTwReEEzCic6VVGeJQicloLzgzHujXE8nxB6Yz+hgkiT
ChVN3HUsO0qAryjtNweffJDsjg9Thp+6H75fprRPwyYHNDKTQYDTFrLjKMREAKyo
25UlBViYbJqAKLBihY+y5OQWvn1mGVgre2mU7Zj6knfMJpqD1RxeSSI9Inrps8Id
mPV86PGml8wv/PlO6HEOKc9scFNtlwu2pV5TmQprpyR+N0roz9yhi5wt+q+cbDcK
9EscsDeOIiDVuqkuGd5cU5L+2hnPzrXErC9DAbRi+2RU2zbiOECCIHvHn4ebugBP
/F0CfjJijaJCmlpz6K8lHkLAHUpk1j07Z1wpHdqEDLA4vRhX6M3pY8tsHIF0w11P
wKBvI28WaCuoWZsaiKUKxdQG/D2FwwguLW1DpQCkptr+dnSj5cx0GkfKLgLP78rR
RtWi+4oVNJTXtpe0kgniUCvHgpEELnTimhRZVVncDkS3s3+YaD4PN/j3KiF+J+KU
gUZY8EWixnp+7YBa4nuD946fASWT0M0/5jTrGe3n5zU7qIIBTS7inzKg2LPNenrd
R5GXeN1T8toPARPGSBaq/dmKkjNeZ44Y7APvnRqlXA8r0wKuNcKQoBxmRzZdnBap
DEf3DNZ7A5GlAyG0SHUVOLd98n17PB9wBh4WGEHRXIjDDnHTrmENhLZsVvxqV6YA
IU/fqnw7yctbg6NgrIlFqn2JIeok0Zud0BwvUnCn/jfKkLgOVklrn9+42Pp30fan
KzVW9zpwAfRHA7eFwWZrIfpNAkyGjoyVXBx+Av9OXHdRZomOOnorJ6aHZmJTPcjY
yG5vT7kgCrFlly9VKhApDIauqbrExIbwDldV0Jmhw8DV8/fwdry364gEBIosUiJU
1X1Sa753wfW6x45o4u9cjDn6Cjh0qVCsaKo0SgXj2AGnjIDitdzkiEIpBVj7eVm9
GwL9KX21cuDBcjGdPkWjbHzOmuWR63AocC63K2WhJ3ym7bMIPkqnzaGguKgJVuoS
5hE7g0qKRBwrm9hPJ54HlXfsRtfc93pChA9LLu+cTY+InZ+42wCJ08E9RdHCktS+
OUVdProG2OK0I6N6zh74sX4gQTT6E/51RM8C/TvHdMu6T4d9NNNxYu3L+ZdYZAsy
5PTzbFpz/7ZH88p4QanxhrRxyqeUYbOrhVl3MD6VsHRaqIWafcMqjKw4jG8/IsX9
C91HwHZ35iXX5o4qixv5gC3nLd2JF/l1apszph/OYA6n9MwUzZrND04PyK1tGVNB
1QrzHUUm6/07hJ4oYV3lLp9XGldgxtY3z9c0MapHnDYNrSzsHfjBA1sY9c/eBsAA
+oj02MGd1xyzY13coecIfaRZEZw2HcwK5iXtdGxVl07GY2Jmk7MrLJsL4h87AIyI
/vDPeidyr14azJftNek1SYPEbR22Qutgsj6MVlSdhAuq5aVie9UPBwSiapCEuGoV
n2JVY7/T51kzHUFR4OSLDh88n+mhmy/NCrnAyAhy327hZoOAzHWzKEjKHkv2+bVu
BjHHgzTugD9OcNr0Rp5LA10DlV2ynen9W181rkibP7gf/csP9M8sm3z4AMdTsSog
Mjej3H3N4h/PCnAbF/Zy5c+2reVaI5HwLKwUWVjFkot9BjVQuoaw3ztybA5yPjwc
HfBJIAevgV5soG8WlUlJC13+mqEJhErG13b9IzrbLbNLrC1NJBLSAS6jjPLeaJ6S
YRXaXQhipEiWnwyE2zP6TgC5pv4K2HwqghBt3PnjlSkHnv114oAdgSaejt+zgGpr
o2Wp5fNLsiHeaVpKfH/UXYa6+KzL9xu0VJjj5X7VNkiKcBSHlrAIUlXyrSScOVrB
UI4S9x0Qe/xUGx7oImWAlqRq9nr1Q/hKZ9ZaEBXKonIXWVWUz9P9V62oYrrKSpgp
87v1ucdbbFZoczMWUYdfheX+R+5BN/myuXA4wWBte3lEBqL2oYfS6pgCU2ICcO5t
Emsd2muhZO06qeeky5ivq0/AD9sS0POvYBziMR0ELBOuO8kyzljIl4h71zywOiaZ
hTejZGUiPawfA9Gal2Uu01/gY80VUgjHfp8xz1IUXiebu4ZDQJX2C4upEgzjYxbI
vP9ad7CcDSzsOFB0lI5fhjmEuKpC+id7jTXe5tZOsI33tJZea09zUyxkkMsCzuX5
bpM7K0MLHKKFpDyGiE5piFtdQ8JsrMiqYEzuVJzkxvhlUp84rmnQXWmGVqAh0sTs
iY+FO5AZkjoZOUE0pTMSi7hvu/9JAMiOm35939sSLbhRrJN8i/HLwOz1Ga6o0lEo
GtUT0Sr0VWXxo4O/D80nH1HUVeetJLd3h8WG+lFhH7F2wtSbaUa9P36LIXtRYibk
uiPPDwyzPqnHoA2rHCKwTtrc7phcwxs5sUYw0Aqa9DqP7TkLhs3T5XViDzR4ubeT
406GkVXHvocnC3LBJncAgzCUjAhkr6EENM4tdUMzJpgzf+EfoFRgwqyF3uT3uwJq
END9p5tdXLHOiGjnIgUZZwR7ZiKrK9ed285EftroeUw5GmMYslC2IkoZX2245x4G
Ou4WT/i+nzn+sL1kqsFm47kOXhbPZnK9XPGHOJts9OK6CkhWS22e4D7kVLslZsjk
gDvDhUAtV4CY5NW3tOUYuhcKzorIlIAO2MDUuDUOyE1NhGH3GCJ9w0CMtF1p08tg
jWNZpU9DPdQUA9CVq/WLs4zgiRodAyQDcOsfj5YoxW0Jqcmo9D8MmYcOlozMRGBH
ZIcgTc/+GxyhwEda5MhqKYMoq01X3ojxNPXrIjToIfEckrm0KcF2mxV6SALjc5I8
DXxxqI/FUTzS8VQML/g1Xr0cp1cQ6ueJ4+9jYDG4oXnCthttuaan9orho8IP2Wgj
gJTwcFQqSa3NX0zKr4nButJaP1BO23C1AFMTBvbTpoo5TcXob9/z26IVq4npYV+T
+1M5iY/23K2fSG+73eB5b2J3NswOxh3S3fIuSUEFhRWzA11hYEqRHWHDxgr8HO7G
B2TznPk5yY7Ryxc9CgEopOpvqYyPiJ6FvVIvYa0/R6BsgwoK9lXl0ASDoAKi+OMT
EUSqlit9J0XHeDmF7n4y6l/tYWIQchKrJqNxLoc8eJwoPlz86FnkU4/8PV2lX9x4
K2T49wCW/zSWAhgSSiXkXppvvvTPQBIwF25I7ripWLxkjZ7ULEsfIpgrJh156SKb
I1lrkXVhjRuXpCZoic+yWzTaCfy/GtmGNn17bUi6pxW783hYiAfRkGzw9M+AttIK
UaV2lFOd6AtrYIssyJYXNIXKOlmAb1xsveeYg0ya7AhI7X6BKgouL/k+fquijRPI
2AvJTPiibmgPMzTKalwIiylgwiV81OWt5s85Ibv49wHBnnrjvkhHNmR0pMrZvtKs
SLWT6JrDIevwUZyjhSQPvVYiNbl7f8gaVs0s2R23Awa7Isk0+dDV+ge6amOEhxBX
EVSQzFZc1PuungSLe+LVvWETUl3azW5AZ5tzV6si2N1gpqKfepopM4y2d+NzQ+4u
Z7NcnzPfMDb33lhyL4ZuYYtF01Hl5nRRxNA4lodz2YN4Pn5SNsbXOuXrV3u/ouoo
xnHvBIwLzdM0ErDFR79sBAsdPgmFw8IT6Lf9ogsF/QEpS8ItrcLpLYcfizR2xad2
uEh8mmf7duCoI5c+TGk/scycugKHmdAi5xdSWpWyHJx4b8RAk0M45vYgR250zybV
5e65a+7rauqSPFRrvOP0ECpiLHWd91lxt/gDuu7GbxsR/N/lWmPnmCHAQGVBp9yB
1QJm7IM84z0QQ0cBQSxVOkDCE3uShisVgnSTujlI0FQ7NE9d2nOav36CpTCnhhg+
6j/Ap0o16vIAaKGtwZfLGKzfStZs0GN0dhaRN4IAbWWE9npiTYyo6cc4HM7fxAY4
zZHb2aLGOihEl4vrFjZk2oGA8vbxYgtc5pIW36/vMuL0zZCZohXLK6IYqPncuHgL
hZFP3u5vYkup3hFKlLSOAvzWhsfl75iU0jzmsbJDWFVHP94CVq54Ac0xFJHr75Zs
L1TU44tU17XKnAysiD6oRpu3HXI5Hr96H+VSAt5TBm9sE7O8RZsNG4A6wFszWr7i
/pYdoWw0BKt4DDkOv1VvKeiQG376it8K+miDW7cK/tIhdOxH2Gdydrye04Lx7Nqw
VCgwuQKg6MTXxT9Nk0y3S5fEWjm8i671vAFopPI07AByVbzUy2kGl9G30r7TbUGA
c2QQMduad5HYG+MxdP0yJ+Ip1bzgIXii0fBRlkXDCFGaUMs/sNYQ2RruXh4hOke2
V85LHqSKi0hbFW0ip3d36rI1nNVwG9Cwj1ASRz3Q1F1Rw9gw2Toy1LCgwP09Rph5
lhupNmfWEDwPpYM0G3tQjDX6f1PCmA3yoE1hhp1eAsoQJK3Uz+ndI0m7tiwqU0Ud
e/YlPgWtB7XWOxEBAEKk8ezImtjZ0hLgHpKTSrX1OD/wUh3ArEa1Qi8I1De17+GD
H7Jvjp+fNTkPmAz9OP2lrXe6OUf9NsNc/qx06j+j2rThFzkLSQQvf2yNzFZepKrd
xZWwEiMIy787S+fOM/8D/f/RTKfhcx0PIaVRdq48GcNDVBonz+j0oVyrkG/+o2zM
ApaxcY3y5cqiQEEjqm3NIVTLtVeXRgH4STddcEtAYtcR8/SLQBy18vyA/Ae8P6Qd
XUE0qGv7na3T12t3xik/HiMoThttiVjBmuxu/DeVOwOYQyQH0boTIMDkDgjxCllJ
0YvFeHmKA+WddGHFOJT2zLZKge+CRCAL+X3JVqsYBOicO4eupznbV5O11N5bi9gu
Nyfzc7MM8cmYI2FnVzOVbroPC5J90WWap500aN+UZ4RaPUzkdZ+wTeWgTrd9sMRK
oUrY5/GcUpB23HvMy4NwzU4+s5OXktSLexBq/3O3zIVYsJddj/+YHY0mFMULAppi
yuHwB8mUx1tnrZSsRPzLKbtYfEz7bDCszigSN+/Te9yLJvsZy3w3z+mgY5tjGA1b
7rqI0E+XEYCLjFkkev3RNAdIxvXZYeAzkW53rI/y44xWDJ1o7hPsdMW/qM/kkf7J
swet/hurIqgQEDO6m+tJvBvpt13SiNOaJbp+FStlHsY6einFzsg4kX7hGecBD46w
KmDp4YTw620ykG73RL0NdHP4pI8PlNzSCH25+J6+M0XhtxSIeg5pOVVbN/elL20M
qSbRp28AgBjCmN22j86W8qExrBBypjiLh5pRvQj8vAIfcV6gPPYQ2A8zj6RKf3Di
qZtheCvjziSJboWpJG4GVKQaOsM/VpjstJwgVPmFcdRaoJnyG+E6YPivKBqJAln9
0UT7R/C6GoiUr1D3WsnR31Jjs8kIDO/SveO50NAFSx/w86KQFeru84qZrvmIuUcW
e+obYvyJWbEwlvszdT7EZibVytZ2FFUr9jbOlEP9H8CPpXF5n5Mp/tbz8luOhykZ
+LdAXNc0Zn9RlqECjQ4SGrhj7iQz9DuBLwQBLP7ncPkQEiRk/brOXKxOrt4s60Dp
jArRsElHL6Ak9JABX7+3NjM2q2b2oXwm1vtPmdYlrLjq1ix+GclSKXSgWpbiL5Vq
Stu2ZRsyLTnOgjsO6QYNBKLoZj9olq46Bsw6AdCgMQ/6CMHbdw1EvBXoEXd2ogop
8+1UlcVIgvKNEhu+KuBGXK1MEf1FL1SCKXFbBmV133iaxo2INZihAqbYFR4547UK
MZprt6yZjTKwmaC4TwVmLIRvvCPCLadhbUGEVQpkvko7ScUll3M2EKwZB1D92mUG
4KzHM1TPDucDST6BKdrTeszU0+QLFfnWTCTNezk0zhLU5OA9hz8Ph0ym+jNE6l/p
NfRu+fwQkOZHndB5YFd4LvQt3ZBHx/RIAyzoMln5P7jw3VEc39YsjgUnyVevh3ro
8HismgvoxAWVP+sXlVa1j+jysxEYtQ9piEep1ICp6IS4mZohvtI6q2iE967xgMDM
gj+sQrvbLfT2u13gWhGrkiwfCvwQ2uo2cjP8h9r1ygFy9i8QZJ9LHxb4JRW5Fhtf
a6LdUVQczOJbriyW/Uh7kPZbcKxedsNfnxyNjV9iC1E30kf9ZyLkZ632WyIc7p8s
N/pdiGCQV8eyvMYX7CT5OecjaqWaX07NEIYGE2qbelmdKOb+i0bWB0y5dwfbb5lb
zY6GJBC+iphjMwkWu1WUXua0wlTnOVgJgu3ots4FC8ztE/DNLUO+9NkvJLVwNa6F
RalHRKKJbtgaKCi/5b7K2bHL4aIMXCfj61sqpf3mCLLdqZeb5a1xOk1ENiVpIS1N
fh1yFBeXfBKT7mNxy2yZRrUEK5Cqtz8T1yiHj00uR1N4+fVQyiZLjtgATHTrqgi9
5ZDJoSEC1FZxqbVikDtWPhnEpB39+bARUqFWtojf4WiuU3SZS+JX+wVB0tP1ABH8
QdNfVPK/dGGwDPycEmCdHlx2KBB2XPZj56YEINHHmGwck+6C8oX7JviW4/H70d+F
dHrwMkChpXPEbJkX/ht/i5f/7ScEDgflZh6E0iJVBOXJGYz+rXGYdoUYNWbXFGmP
kVfwmULCD2NqEbeTgPZbubiJi0zDEgJpj+QvgxN7r2B2v1OGbAwmy9ZWqDC9HCnj
2Q8zwuqIFAgJtMmxgDEIElVvzMnl7jj+GPABc1uc7DOcVcTsyTjb0jpleLzIjc8R
oMXJmGg+WgEe7IOT7gPmA/qVN2QU0hsBfvhlt/zZPjWzwmaxEd5xPFjYW+vjv1lE
GKKkkEt85MoU3uyXYa2KZMEyZzV2riS324NmPKCiXA/iBuWkmaJ8itK+3IhF/kv6
IONsoZP3IIDZY+sV5/juE94s00XWIM/d5wEG3yRDncPa/36n/1UXO0DwUooEefJK
vWsMMVFW5EwiAvmFG5Llx1Th4ZpPUj9rZSIjNKfz5cdlRJ/qXyYFKnc+TvfxjVH9
69oEJSo9a9khyid7XH3k4BpZyprkzaVYRy8LMIAf2thwJuwfJOuqJmSG7udwRRZu
bOQTdQjJelkxL6qKhEMHKWEXPocVBFR63nhqUUscfGR4Vc44UunKZGOtMp/yYyzk
4izIrvNzT1VVM0tc0gU1tEFF0sv5qEq7RiKUXU0a8FOtCMCNciNp/CsKp2V7+F6h
WCqwIJw6f9xu/yzHsVmDezNCZmLOu/rMmIvf+0f7GpCXUvsaFgUOW6stNEQAkj75
FAcoCEhPgTwgBy8tYGwKLNg6kF+IUuGEhv+CJLUnpEtkLWQ0zFIieOYrhm2L4xXc
5HPLa1433NxcFBgSfUQvJBW92VUW7rPbY1cCJfeKlJC0HxQI2mQFt/BFdQK8ykz8
IFQYFCDmwqtPWWJCZ6lr0HTOOHLRSvIVpPOiu2eGESX8EPBBmAE9I91fz0Y2LyKa
oNZiyhp9x6jyc66FfP0rkJNhrCVwyBOCgkpopsKlzzTMhOdIl5UdXFiLpBD2DxFp
3Nb/B+AgBtOd75t+il3GYHfvdkLuqBvTK90E11WxZU1BY4e4La+0DbuPbhlZbcMT
1E/yveeo+LrJA/l/Bs9b1LRamQGnI+b1KXjRm5eTHfCayDeOMUo1oniualANJExG
67TmB9rtXin6Uaw3WbilmGZ3/s0qXM5Nzuf5KsxbEyu1a4DzyJg0oSeRsOeb2FPb
ud2dJ/jRVdXERZ2KMu5cUEHLdi2s1x94W5Z6cwSDur1FG2CcpImBOvSmm5vT8U2B
D4zF8dbE9rH2YYXVJm23r++P4aFT/z1Ury6xDlmuMnoSFbdWcootwiY24CymjUS3
gN5RpGX9mJ0GyCkO6GbA0aVzAodrSJjxniF+87LmArvEVkfWgeSAtW8VzBU1Dwzz
jNC8jEpu9Xt4Mg0TKYZBnWxqvPreHgFeShLLoB3HMqfmHhFlMTfCB2cQ2CEf8aY0
tPbPxZIbu574fzC+SRyHvP1NxkwjyebKdMVSYvhDvTOcODjoQsEpm3mJ87ZrBShC
lUgnpJT7NrjkcDojorkx5F9YAGW6KsA6Fu9waWDHiSnlGcWgS7vD/XJ/Pj4lHmIr
Icm+atM7j6/nldqOx2AikR+HZAMRkTFrq4ciPrMINoVTf1jQBDcjZ7/AYDtXgS+Q
Y+PSB4ZlEZNPQLnQbMAbHjleSsdKGItw5odDv6VCtqLf/oqN7FhcyYYSJn+mLsbt
N+CB/ZV/xzw4Sgj891T6httgPjiQhmbY/gJgHX7hEwtRG9gm1JEkK/y434E69vL8
e28mPK0D8l/AhfkubjWuqv0iz3P/UBeV8MMBE8mrXgPjQa2PcE+gxKVuwNdCseYl
UdVKeTWxzXKklxa+IMDMdkFIuqy3r+wuIP83OYBwwUMQP6BzcRcaCR/omFAcK56u
B5qF8BodaDi9uszGl5Pu3NVhxy+iqdYXMT+8vtra90M5M5yhqTvSuIdwnAqk+LZw
GMGDtcL/Akv7RCtCttcWsXoribU4i7mRpNxppkN6Rt0qIZNTLl+o2V6+BmiEzxxr
eOAkiZnwRM7ilS8qIOPMExFBiGy+oOxWZnxe+bC9s8VaZfBYpF1rzYB0x5IQWHF7
h8AqTW3Wisw+OUHkwFLrHagQeGS+fttDy0nG62ARRvHt04AnzA5RxbxDrfb++Wny
T1t81tnzuDHAva9ZTMCdsRr1dv7oEe4RVETj6jGHrvwJp3parn05mLLBgccVJTmE
giRhbMahdVuXvnpIkhnUM9nqzHzsDRk0G0gKGz7Hmyq1CnFeZHIDXRVIcoRtlcV3
8FdBoBEeKbloODNtRdEGi0M0stC2yGuWIrVjuPJ5f6l4XuChzvKvpeBsDtpY60Kx
kCe0ueXC5AESHoxwdP+itSpw3s1jf6TWd8qlIG0w4IavodjUtoTSHGf0279Xjk9d
1E4WuB5lNEH8FcKBpa7vQ8U1OK6b9yS/3oSP0VFWRcTmTviUwMVJet5eyi7XPiNQ
AvH8nln9jOKI49iU/16vw7JZgvZt31javGhqKwikCpBlSvH02UGjby4isSKTELha
7T33p9bbUCSUn7tPluVTH+9/0/DqwmxikZrKdAG/uRAxo+BzexBab+EWivHxe7Ai
qO5Xp5a8MinDelkvqQ1w5yIyNf3E8z/+pL//x4mvhy54lB4b+T5nMKhwAUGOJ/xI
XvYN7j2s+Y9AxJMIVEvANOYr3EdDq3gdydhsgM/E5GRs/x68InNV/G33fATEtkn0
EDSxGsdu1gsFg07M0W2pXkjJKbZ8FNjMFRauD6iqSmXVNyoKXXsjLx48vsNDGQrx
dpE5/pHX4vcQHWEfSPPlVRSR6mtgyfTvpprbXAZP4y+kR/m8mkeAD3ssm8Jx5D+/
Wn2nHBcBlbhPrD7BDAby8f+glE7iqUnCrv65U5rUnhZBjNfnP1re8s9DIVN/Bah1
bQC1AGR8sKxxGA+93xJ3Kcg6u/qicbM34VnrSx3iVuM0aeeztsc7oy0kNCcsnwsX
VzpGFNUdwSE4/wtjS8jisV9X6P+yMvJasLhFk4BpKrRWU0AbgJ/SAP3KXrILQmDW
jYOG/ahhCtYKl2xgeK0JWEMwtyltb0QPVI24+HCF2iXwnH7ybmc5AayISx2I1I2X
cg/hO3oOle2CJ1qQtQMbnQHV+tXuq0gouA0072qPNQntQStfvO2Le2TUkOFpHvZM
gtcxUe3q51thd6gG4LhiMcrBAHK4bDjCCWSzNT2BbTib5DToWlBAiBSLTixK70vl
9rgY/iMNU1MDmChfPcGG+Cu9VMaMMI1TXS2alHJ2chL+ZDrK6FfHC/1epPr7P6+v
7XELd6uzFoz7S1LUe6CxH8jD795sE0GLjnFJ8imodDTLA8eiiRr4e3Dw+KzJzA2J
xNXotc5NBYqwc1n//2zodZ1llNTha6N0cyleZRNkULgyhRMl/MA33WZ7krKkJp2D
WBLy2NvoqCs27oldSK+RngVHaQQrM6FiOWRtnPMB9PZp7zcC8+jYpGrqDn040JKW
XB4jMQS/8vA8axpoBfzPHqdjOqS4gqxHRABSeV2o85YfnJVlPyYrTlpXbX6P7Pfa
WF8PCdb+e/aVgk37hmpKCCVL89laFWTtpriLaujmm96MH756BlIpPN7DMZ6gHdsa
w14OywsfSA7+CLc6Ebzzkz5KGITfjrv8Np/IMQxon68/tu76JiYvw8MI3rsdmTLo
n1vAIgRfm3SO4lTkIoejwC1Y0uhaSHyuU3E+07BtVSwmpnbF6IXwYkfjLKd/YBTA
AbTh+Tms+2FmYC0UdE85lEd20nNZwPWmTBAEIs8OZMbxAmo4FxgjgMr2gYOpa8WO
6S+drl2+koY6m37f9EVKy6sMVnJXSWqhCQ2+oqI7G1EFa8TwWc1huxQLPBZhgoRT
FXUezQEtWxHivXfXcAgMLdN16y4M7UwXlXOLsFt+Xgq05GeSL2GoR7cjZS3kYL7h
XAloMXkyfQzJWu0qhuUIvuS7UC4BFHwnwnMjWHnkhlM6oYMO+G5nhTRCdLQpXlHx
g6P4x1bPQnb8gSXPFku00muDshXWZSAT0vQplQTkM+9pyCT6ZCrTjrUar3X6Jm7r
RsOvaz1nKAHio2ibWNb1VLRbovRuOUmyOkVY7kExNjizzVoQHL3/nXIRt+IkrjWM
DPlXMg8GD3qd7ZgBXzAKaIXzixalmQTipI6F22aih52dZ7mtsZ+v9h4Fl/XU3loF
4agLodImyC+6n3uBU46+LSpFn1cqou5UATQadKoY1O5SIpHbeKwqW1bMK+2H2kMM
v7aVuXxICRCM+XBmJaAJeb0rb1de316+oz4YnC9Z/7y9aA1/KerA3BJYrTDGU5Mh
Npi3vlhNXeJXegXmYiHZf6xtwo4EdvPtr31odkWa5LIEs65nvJga4FKhpsJHJjZ5
SINIE0EZbnGwCuj33hr23u/OOHY8gBGNtfVlPv3qYjM3uqySu0Tu9hsTMpcB7CPB
if2aNDm/olz6kRKNgtSW7WvEOlyHvQKMVgW2XVadwmjuFjnn6gQHbAXNMqkMmV/a
r7vRmD+6KtHbQU3SgBnwOSPpnj5TAVZUQZBL7o99apDPc+EmEflc887jEihlWnNp
G4j1MgC6u2LoTKaFwpNT/ZAbRA5+CEGiOKvRAYbFnZKGDUm4LN55AmB+h/u4Aoky
+Z8XRHY+EiAtUCXEWISwSvbI3Lz6iVvEbndvxGkW0LCVESbYxK+7YOxq+6qCf6Sd
3xQaPDVSbdyXUe5kiPX7DBC07rwAeyX8rft7OG9q3Hw9aGgfzzAidCMoOCDezyfv
dRXcNEYaCQ5POJndTqo3SgqvU6U4SUGkCyKC2Fqn0y2jlGEB72CTKUjuAtaJ0x1m
ou63ndSJnIUpLpINY6GCCahq7oHFN9rFtn+7Zca+9RHpmwQTqq4sP/OJNkAywTAC
ugjL60ETsVWM+U5l+1OqZHtUt44MpLrwu+/udQkXtCs5YS2TzB01L4yLkrQE4ucB
Qcew7iFrib4rrGBvBJgHvFBSAGkV36tb9UVgR6EAdB6xJTtbOdVdD2WsMEhn0sQ9
ZKRKjE8Bs7DbI9BqLDb5rSAzglJeUH667ma7WJAudbaPmNQojaesoDftSGdbkLkl
Qw9SVozo0bftdhEpZklwRNbVI0VMWr1nOl3zEJcoNGQBIqge5d8IMevu2BhQnkoZ
eyGWwZP10wzoajsIMuzLEdo0hx08IQiLuj9EvWoDYG6WTRpMCvCs4lhpQdgB+eUP
nBCoo8JSw7SWm+rsI63tTSxTrA49Jw2d0lg4rwSJMi9pfgIdrVos21Nu7HkeQfCH
7rhZj7Z6YMmLHxZnmvfMVDWvWvuWZYREn/1zY2yNTmNP+peTcIgH4B6DXPg3zImz
YFw1a1ITK82ZkU8UBx6SVrepd2+l3oxf3WL1zs4GwWuU/RfHSgbxYcmSceOrqLN2
2O3Qd/SaG3lzgRQw8E13l1Z3F/ohp7cfmKqYkQ/LzTEdDS69lnjP6IBUcTcNFDNS
+2ZKlViwaz2r+vjMtA8WsOh2OMtfpWrDkbyr6i++dDdme0MATgpdo5+eeOpEhT07
asR7a3Ti7/t5+hy7Y+ThlBtm2K+Hjzhu4lhSx32Zu62HXZCT0ZVbtACZJMoV/yLq
6WvoUoh0JgxEFtP1oT1LFYCbZJ4/5f3IuVaImKfeedcG+H0Q+fFXoT3/GRSiM9xF
btwuVXpzmMN2zJiLDAKuPN6nhEs6AzDVTTCIc/ZSpeH7AYwtHFG9PDp63EHrYzeH
1JbqENa5olBwizv1OonkpLtke+WLB6EEe7OIdJRVqWdLrA8ckW6h0BzL7WAAwl+e
JRLxcmzNclzr3vgGO1mBMjOyg9I24IjCBGkstzKz/+xZWO7Rj+Myc0EDv4sTvZsP
ZZrSZecsD4vZx16OXoa2p9SePx0Ufz3cuvZ9JhusuYsZX7ct80FguzPpTHZCTXMj
/ARXnsqqr/15l0POnV+6f6HjNJS3+xEJbM42p9Ul6MBHdIRxXKV2P6vmTKByUJQH
TEcE3oguCSWTcGoHSWzmhRVlSfVBoyNLaC3BFqhIsJqQmS5OqH/AyfzN5agSboOu
uCRx311VTABkLQDt7a8vq8rABnm91ff+sLlRvGNMxpU3Ri8LbVMPWVxLWKUUwKEE
RJb1j1WyGZz/voN74EYpMcvtRKSlrMGd/qFc5nPQVgHRMEtlYtlQnSGwxmZbJiN6
hPbdKVluWCtLaZSfK2CYXtul6tfA4HYT09vod3f5ByChCS/C3BZtgQjK4EMRopax
Lpr9jIweb/4QcegIjwBdJZ0h2uVAs2s2yANTSTPh1g5XUvJ1Zb7lA6ZCZyIQ/Cms
+fwVPd6N5P+ItVlILlBF16yCTNzNnTN5qgtt9n5CVZQTROm6Obl7Vh37ksgOY9tw
N55xm7lWc66fHElTcxVoxpbjpZTRwK5AErg6jyAADBauTQO7WHg0Tb+9aEPXoFay
vzeuf6xoAkdmgvxX1oK4e7RCFHaQu9WqCZQ7MPPya42xRJZtd/FkXzS7Mab+6AQv
ScYlra0q5dVUpBzi91kw2pIhquw0USfRdb87PkBI/ubRp0lxTez69EsjgRzmtmRi
7Ud2HFq/Hu4nI5gKSRgJW/YHfgRJcUGB1WC7cqdMWOdXDpMPQN0C2UFBCVL+d9kK
HYWyWbyrlXFKF3T1/CA2/qZx7h4gkJSewjHKuCp0oikjnGKTtviOx+aVjVZi1wrp
tyDZVGFey+2PwtW2L/jYrBJduJfZj9wTYQ8c+f5VGcIa/8vuqLDbboaj/r4dmNBs
jL/LJQwi+Hp8eaXU1VfLitwuxr4f8s0dIPhdc3oosVfcfDo4W+a97PukzxAF7QMl
rxraCYF434uDTARugPaiXu03UUd1kBB+kXxvd/npg1bjjbpTB97i14giUj03uY1y
pgFrLE7X21jvq4cXcQ2/MtElQQ2irYuMMYPHsnud7SvmHGTp5m97FudU0Rj1LwYJ
1oi7qsiGpsop/6BxSg6+ZvyOp/oY0+fHv5djS1Y7mN7MC+HmWMcLMKEStPae18Jm
be8lYpctdAr0cxttaLjefoZceEXSwRxr/vlBXP9P/0D9hGWKW790y2F6Kx37wT/j
6Z5AzXlYweOdUNjowdqhEXPl6ykuxHumGfcxX2MHAaT5lt0uGgcVSI/mXRpIDsCZ
rkh6J/8hS3Yj8r+hX+GyXxZ7gBek/0KGzcVDhkR5a3bHsm0TkcCLgZCKVgE5zGxO
47IRhw4qk/rBdPBYCI+oFxwG7Nt0o5wBrKIV4pF1EsZQyK+4orUXy1TTymWv5gVs
IATYcTjWJJ+zlY4yuBqepgPL3Vabrn7LOg4Zy4oGsvGdpy39BIrX4w6FNjfxdVOJ
Nyq9IavcJxR1PsxNwGFkRwSEKQ/hYqib5p1i7KlDwDynbrKgt6gcx/CtMuvoqFrj
axZWUqajn+m9cwiuWY6F5q30JHLnIAqOH8TQhMHoDbCcC0XcDCVdVz7ZkSNnMDAS
vT+0Ay+DOHAyLGJbjNJB9qhIFQnMJD60QXo5IFuyjLvOw6PvmA+95UQf1SmpNpPp
1F+qPtuVuQK6GTkOhaQj/NdVQ7DViYIdczOGqMxmTanejrLQmytYbwZUr93tg/6S
SVY3Ze9InKytUuIK2YvH73DYt/cfT40bDssYyH7k67397bxOC5dNRs0uJnuN6WO7
oa6il3aVTygR8Sj4o/+KTYc6g4G0tP883eL0dAFjBB9HkBk70EIhORFl6PWBaY02
WvcK/ObwZMt0f4a5Ez3ddvyV0GFc4gPK+/ge6h0RiRtQZE+hzK4UVJ+VccfY+BQ5
Jh7iTXAw9oXPgS1DeR3G0RN3E8poJO85aJI9bmlphueep4VJkCSPKI3dVsrHQKCR
xvXeBC792knFQAUZmpFOMnvZ31tcmgPvmiqxRoXN9PS9/T3arVrbDoxq0zQHTc4Y
fEO0C2BY2sjHQfHoJl5zfLZunkqYuSix/5q/grzlB1rddC9NBjQZt7DnZFib/RV6
fM6EK0mpeVZv/hAx7OKSJcmwdnw3kSXH57ClRlyK3jx8GTZzv9dDTnMVvh4G1FmU
sTzqonp/YhtWzGGc1ICZ2lek1QGbFSuQoEjA7RRRZT8GJoK11n4q6+1nOxZAhX7G
MKRFpVDxt8zvHW+tGBdoLwEXwAwH/2BAY1XzMxJTdq83t5QnE2qTiFdhx2y/8fIr
IA1jjwAMX96ZtxgorbuOouEWJQzu/k52ntlnEG5yuGASzc9FERmhQUkFCTfWkeXB
eSsokd9yE4n46hqda/fdmX7hyyWScqn83XLsA/Jsp7e1uwWOxPeo5FtsRN36R7Tg
Fc+Gkubiumud7bZYXnHZb/ReAc3y9ltO0yzcXYSNqHsQ9iTFN28rfem/HoJ0/40l
7LUKwz1cUT3ejwH1VyHY/QoYY7Biue3LjXls4iBkh0NhGdTP0gYfG3n7haJmiw4S
T2BLiF7tWcoZzwiToo/UjVunlNbRPTX/EWqApzgZ7ZGagYmQJ5XYfAZ6qoc4PWfs
vZDWZcqRoym7fbdZ0V9Lndok7SAa3q2zGhIWic2EpaY/eUFIIKEp7OeUioJXooU6
Fo8efUVplOwqfv9DwltqJMhpYryJJEMcQhWPF7AeEddRznA3/dPaH4j8F8Ub76Wm
nAia2yeW7g2ltNl4ItkNJfNT1RGDjsj+Xsrhim2A28+TzL/++grg5Je+1XopdIO1
kFbnyq306TX0mcbFvHFSZqLZwkYXCCE3Z34kTk+bLNpwuLRKijXrqvX7Fl1T8xc4
/kIyHO0d/TzkjplBzmFUAdccsUWwmRtkLU5VndWhrLhRYC6Ui+GEgRUNv75bd2nN
fgao53ErgfUekwaXHhx+07wRFbTS0+yb+12erH9bQd7LEqMEgt/iWGZJSROVlAvP
m2lVEirG7QldbgZvGX0FnQ43O/fy1uSd8XbZ2mpJegxDC5Nr5BKLSCNVBP2jRUx1
wUMGhKILWDxEVxWCSbuEhc4hVMH01L2wVyjurwGq4xqDdYVZkfq9BK/hVvPpscDo
4iyiqqQPlzTBfEBiorUcolimIi9q2Ga0E854bv9qGaCxwogSN2h6rK9XQbDxEA8R
Ozt9P2m2oxmhPAYea7NuAPlyj2nZHvXQU2eVwLJKIDSZR39k+C6G4TBnTWCxSJJs
GhCxSon9PNFGdpokBBo+6aF8Qz2uyi4qB9ezqyXte3TnFwxgEIsr5HgTa1feiTHw
4wb3KyhSvx+kVMugI0WTbmjhEFmExjZKqsuwwhUefY2d5m3oslDOEKnKSB+kwSpx
ax0cM5ctVYb8FYJcHXccaUeYz+7/QqRvpbFpuhqtZIUOGiWf6gcOmZv98kDUOx8/
ynjpQJkNY2ZnYJbWFzOaTXiIN0pWqGVQ6zASCD846aukmnWnpkSqWpXJiqbkR2yt
sGwxfjJnrCdkJADgiJflhhXydWalDT1x6emoZ6je/amI2L24aSA9NLSmcs937uqm
TKzCrX8HNXpqO6wyJ+JQc8sEfJdR4jZ/dqXq2tlXTP0EGXjnO/upb1K6W8haMgjW
gs3qg5+tGOBfSe+5SuUihAw0QglF6D6eu0u+2T/rBN8vJhSp/FOXRg1mzBcWsDjQ
yXIEXZNjY9klqsDB1cVv1sXdQ7n6KNVqTMp8CJs7O1CpdeiBH583KY1DgoLjAHB7
Ks/qUFaYyJdwcMG2PZUjIfg17+O6iO0MDqyJ+Xao0VUwb7DbIOkk4/DBwYQMyeNZ
bdAhgTuorbisa03bQN34l6orTwc6+mI31cgHHZDrgmBpOFbI3xojTqT/9JjFlh1x
jAGmxhqnQTn9lNECgtAWkvVf2mTniJoweVLnjzvdEYPr5rF50oEWoZdfYAYa+7Yf
WjEfKSyhtD6DSfvkuWz4Myr7pdbwyXhn3TQMC/K4zIYKulTModaudjDP2aqI8mQU
Gily6VqiZ8IMol7AXl2eiF6Xod/bE4oeglvDFDIiH1Nh7bg7nty3F7nkLtmUeMRN
35/IsFJIvYj5FiMB6BgJt4PuVNc1i/9NTAi4aJGpZnoFfzMP7Rqwt95frpRmfGCS
VRQMdqa2EFRKAzohnVNrd/KqaX/0vLzxVRsJMaQlGb+FRA1E+jYeLHFla8BUIbBu
l9sGJSyJhD7Jk00Ybi6YyyCJ6TyMohYwO/1qRkvj+ueusVPB/3lxGaXoB/aw0JAP
bqQ+Q/I8dYicNhyXWhpkxCP0ZB/7Pq5hXv8tP6JfOdmQ9I7AT73Dmtc9RHG+sCCu
XHbr6HvThJg6vmfGtl/t5GejCRCEe9KUYSWVmOADVE65VbP2HcXICsG+Aw90eYQk
dTfB24Kg9YU/+4d9QevG3VoMqdCDytY4ZIZPIsN0EcfZjym5NjUnxuulZgGjwjgc
ukuGzMcx6XwxOzJFAUdoP63bTZdcdKPuZgOUupqFRf4WBeIMHmkmCqRH9KkDa85e
Jcof9QLhs0kjC1nCr+9GIvGQaGzmou9HWbhZNlb0bTEGKB78fF5b8AU+MzSsI/Mz
mvm1ZHyq0PDEoDjn5obE2azAMUpaWn3jkgiYKCS+Xgy5Q3bcX4HkHxjVZr7O4Pn4
FiG2gXpeSjZ45jMZNrWVwrODEyEd6/ud2hB5+K0itC/8xpZ1/2kKjc7g0eW854gJ
nlL21o0QRbpCZJiifXRra/SemSX+M3VT3O0SGYpqsOiWxVoP3lM+Z7TmSsoQ5E0c
FZ13TSpszpDCEZebddYcsm5FXdi+D0M3n4rU0QYRJj6Td9Fu2VGwPyMG/VFbi7yE
ssV1WVzsvJ8LbRXirzmMF1yzEmSru9zUzhj4Pb7gue1wX1alkkLvCVW/vRsjqBSq
PjsB8w2MrObeN0yZsy447p6dO5TqQGiHLN8gJ9/f6NzmqOs8tIRwdyzcZDF5uFhJ
ObuZ3sahWPiR0nzN6Y9GasS9CDlzxcXUcts5+8q6D563BCK2ZtowDfa2CkYRFMEq
Nj4A78WXnr5/3Evwfqyr9g7mZRaU9BqEclOMBAgp43eySic2PHoRK11E9iCuHE2x
viRkiwu5pe4LXuQV4jlsIeosvR8LmdJUQI8+krSgNxroJmOVCSQNYeiueRPF6GAO
fq0UHO5bC2c0u4dPCKzR2E3/Lo7EWrthRQ1EomzdrLZBjBvnik0ZUrn8dpex7lem
5tG8/4avAOf8qiZC2okczlZwX7c9ms+sNqCMfxhrZyenf8KVw+65oS7mhlUnE+2d
IwaDGqO5e6NnLLnCpKcMbxTrYe9irfFEzpI9llJ1ZXCNz6FfjziIer9SmblZfq1w
zfgzewdut75KCTwr8alViNNfZo4zVwOHSuHYo/rOFuUoyy9ackE3/JmXPEZB2SSV
/LtqRa2B/ZXBOVJ4K0Ew+9y27vaNW/qhgLiFlVwSVfv8P8EbN2/ss4IhJcXUvkXR
59j2YeraBYWuy9iOEiROY2GKISCvNgwhTCwO8UZQX+YZLcJI0PUm/r6ZBF64BwhV
WOaV3q2zEmqzQuyJbsIoZdcqzJ0Hvgl4IxSPFkJG01NAfBuTMji0qHzL/BozlolX
342iunV2sKHgue/ZhmznAEuNyd7TCJFTs3CFg22f59qqWfaEuCFtQrhaeO5DbPnt
V4l/w4k0H507qt4pR+bDXPPn4ycTVEiDGjbS0UAI4BoF5CwHLLXeak1aA9ViDxq3
daqaRI+a6JOCD4D3K4wE5AdHGY8V1q87kwZfCBO31jhAyb3mD/Utuc52vdD8AigB
hECnvGTtITpniE8xeH+yEHNWej1Wk66RTCsHKB/90GaSNIzXNfhA+xDlqJuxIfmW
l7Dr7bhp1m/bbL39ZyhSGb0GI7rF7iCfTT/nYNE97Ia8GFNjBcbYn2dEn6Toxgbc
4Hz2tvEjbMrhSP6uaBzWxL7jLq4+NVJgGboXhoLpAZgnBYnmQc0Q52YbI9+zBczp
3GEyVvjy3IbOPLWxa+vAw6tsTnk5p0Ov+KQ4AzfSsVF4s5GeNk5mfoHsn4S9DfDZ
6MoNBVVRy1l2M/gIfQxU+IEq0Yy+uYnvmQhx8KL2l9eUnPS6K/vIehYOuOQh+ftv
6DEB8kqgV+E/hGRaCb6UnPlpLwuw2SZS+5pwkfmg9N/MWLMs6hnMV7wKBWHD9Wqb
OHH9s6G/CYNx8NwOEbCpjiSVYh+zLAsaCqconFiX6QMeIa1SB/3bwlDEq9wq8DgI
TWPq3QUtpiCnwYPYtnAT291IidDqahUfvVtXTMNTeEXD5ziwi60gWylgsn5Frtwm
G8mecy6ZJh8kCRar75+YUIwbuAW+Lsul1kC3vbMsK0GyGLnrOPEjW+i0LZuyjfaC
12Vekg0SI4HcBfKwaCEfZQ0NDK/FHzAoIPaiVSs7NwNvLIwE5SnePET+ppWae/8Q
ftKEzBoMxp8fl4w8PXmRR9egZeL51EhNEYARgaAvE6Uqmo+5jMOjPk3wCb9nawtq
uAU2tnLx/VaRZtVLb7Ed08CPbZc3L9KYvqEoesavOhQ9shqE/qri4XX00C6ftRzH
NwIz285VDHYRx6MFwhKWfbWjeIH4zBMBFvleSNwhf5uIBmCaYgjYyweKfRji+jNs
X7OGqFPN3aFIWC98coeErniQG2eNmPdo0Kz21BKxPkepdoQH6wV3voDnhRCDK+U6
B4abCR+i51gjIqTwemCs/7YR79izYn+j3LBZvG4KbNu4G6Mj90qqqcD2Hc/wmQ1p
cubFo97A/Dr/E4Rq5hCAZ+117B8oYlWK3Qck4bDx30BuBIHX0+nCQwxpcCqT9YJh
YXfVe8ZFy3Nd1P47IF7iEcN8XzD8drlG6GzFDpA8vwDJOOwzg0b4vtkO058v5DxB
bflz71dFcu8BwaJvw+h3ITtVNce2NLFU00cGuX4AmKe9YO8GrdVpyC55VlaobDSX
DERMXYrbvL9vDdBcwoH/PnFq0akylEyfm9s9mVDpLX+ELNJImKjLRqO4eBm+NNNw
OtjXKgucDTyRxDQg/YfxK2yA7zK32P6Iz4lcRNrtDbRN6DwjcPYwdQThFvE08Ew4
608GKx8PqE9KWT0oWglyZu1VnPLzORdG54bpJO9jFymSrmcYd7sLBAwd2vGy7IME
fcCGmeFE3Qm+SvPQV2w2FXdd4ji9sYYvcuTOlE4RrrXw+oN8cLyfY4p4HmzAT/Y3
fPl1Spe0MCp/LwV8BDuRLTJA++B7o8lDvtk5ote2Zm6zwsCGDKUYhXfPJBcxW6Nr
5R0IdkpkuEbht0ehN522aiZljquThCHs93+pVIyf18aqwUenmsaPmvDhdTPULJUR
9c5cB6BP2xx3F701jeRySDoztP6NkyqR07d963ZrTJ42Le+dZj6VAEG4e++Fdg1r
NRqAchFwzAqs7IVW8FmjxaOqE9g1OY7meLNkATgFDLXeJM/xc30besBrI80GH9Vp
sF4eV3oSNlfyfC6Az0NnslQc7Ms9Gw12IQKFhTUve4jAF90MPbktsh4mVFtYqfv7
8Guu2yCOrzUfvsXQWXKa1s8rwVjmrC60x2yi1xWZ3Bi8PRcZtBKh4PoVGWTmZ0/S
lx5q6ep5ML3y38GbfRpzcy4xYa435nuLbWWM+AZESxR2Hkf576CRhYG4YxNpouhF
2RS0DL2qoJ8FHZEU37ykkz3pMriGqwQwHPi2JlOpIqhJORUNrZw/nXSni91OomcU
6zhTrLVhqE4Ew33GbN+0Ksme+VeL/6Fxvcg4LUNN9HgM3KlWfwDN05DegKkyNPzJ
j55VS1ULycKj5dDl2BxleQqF9xFf1ZsxPnSYSm7TUJipYakmpuaa64BLyMw2lFyO
W139876p+C6oyWSO+MiNGrrrYnlkc3zibfdqHq6R0CUK+i21KlcETv6T8m1urrvt
VjYsZQ3YH/blmmOYDMActgNDtEA5qENxMCB3QAzuDPYXKSqfE2pX1RK9fPvlMlHf
U520Sl057BAaeIGvAN2dp6O0g8y/OUFkix0NHb7zntj2YbMbq0Jape+eLq5IE9Xv
PVsF0jtWl49xrwdhmFKXFXc+gPDZ0X67Lx14cw7qtFQmZLXV/Vq/6GdWCNbZyuxT
6uha6ENVtDCOdiDwX1Ezd06Q5v5LoTVsBCgBvrhH+2lkF9N4ZnAZJGB7IGZgUk3n
CgGxyLNRxJJV6z/L0rL12CLkAHMGnOjBb95njc1k1hRqCh5xZY4YJK5zu3Llb/U2
eEB8TeRFx3OVsryvvxiXMMGgKAchRCb9HMkxlraEAjLA24wLUBBFP0F8e+gQb/52
6w10Ljqk0iOn5r7Kw+6ZPI/NC/zoyogGklF+b5YbPqPVi0DILYEbgBAX/9OwCwPa
+3PnhAlkY+leddP+Sappym4cIPhP7LzsEQZe3tbki4M3a06Blkid7zSNL2ha9Ugx
8RfCQYQztgN4KPLnq3cvhzbA0fsrJisV5r3S+d6dt2s1w/0blXA6UrK+7oueeZGF
sSmUbKXLsATNCA/Ev5EM/tQ2PNb99CdkkcPTlCcg+ANd9b+u4KyQjs28+Nrkju6A
a1b/92qHPVwGZU8WzqD2Qqd1NcpfcW2OvaSIwW1YpnnOoUBUXJwVyJVVFemmJD1W
vcbCZdFP6FGfpsYqBIf9m7eeZXPgnPmV7e6Oc8GNfTTX6a7wkfjjHRjl4vBiOFyK
w/VfA3SVW2FZHRfj76jCj7kpavJP8Z6Ct7Q5lubPsOI/7K4L4I/GXW8I3QDxepPZ
cHFS914QFEj3+oliFm6y1DJW3QwgpvaCKcZP1rVKFqOVeIZR6aafWDmG00q0Ahkg
dl8ZJ7+tgau/gVAfDK31pKCGTFuuHZpsx0ZGX/txVIqy8Ws3d9CCWBxZvaTO9sPF
ztOf7K7DSotHQ/w6N+KkIPDKNAw+nYSkEFppRu5NFZF7P1Y00/Hl6Gk5gWqiSOHs
1/jxm2BywoNTWqf/TdmsUD95s3/geORmXzsv3gsiY7dv240ZYyB/F3ZYS81sn5Yo
092NrcPtsDXbpiq5XKBrmdqHu29ClY7NuvXHjAL+ku+5K/UrkV+0JqvjyIsqnrjE
xg2PLkm+vqxiOVWqxgf2YQpJXO0lnbdx/OkcBydDCbQpg1y1jJTVNMEwpN8ssm05
QsRgI7evF5AvlrVT4Dvgf88c4DGbMU40QtoM6IKwcZ+xV/rUwqOwCuktmLP0XL9o
nyxS8HIa8cLKm5W2omD1jdTm4Wozgh4wSzOUpdNeN+Vx8l5F/+/cts+qf2QS3eRL
49qVt9IJJzwoIVdWGJnSo/rrWMFttx757YhxUVX+MF+7wsh7n3IZ2A0z53PzvPtK
EfDMnpXTOkzR+4tKxVJhCD6A78tVW0XOQJT6Uw3rRGVpdus/0F3BeB79b1O0FHSx
pvjS6jePTHzjP+JfSEO6oek5u9nwyyWY13kouIcw5zRbgY1J9Go4SoVJJnyqeKWh
52z4TdlCe1bRto4hXWTF99NWOIBjuJn4uDCHw4Ix+rBn0Sfc/qE+Y5jXE+dnHnDc
7OcdkZcvzZSK/ZWhTYTSqa6fe97c/Q027vE0pEFY7HYEg67NnEuxhZ6Gv13eSZbo
XBQXek+g8SBH9Lzqc+i1Pwz4rpaaxk7hiXwGDe1V9sWVBu/NThLlmgIv3p6DH4Ut
6mHwGIa2Z7gmUeOXzkUPxq33QrcZFYvlHmeHkspHHIlg0oZ3LXlcAufWveqnbGLV
0ViJ0MIZpI4baXfI8X7i6NF+F5KMzUoacF1voVdNXNO/HbD8+811gzQqbGCZ4Hx0
ANVy4gYBQZHlffI0jqyFz08LB0wVTDxa/77LkY1fMZE8cHE7gbFSDcEfZ1nsMzME
PCTYSfBD997cnLzpg3LFamNglwGIRqv3RoxwxYUAn7HVa8L2mCjKJ09kCKDnZadY
vEcn69W3Y3DWO9yGDaOHdz4kpFMlhhKS0EokTLcDKWC+BuZifNnkvZ9Rov8Nfelo
SvcRFcvDcPkvvcDzrZwQLyR89sG8v9v1USvZddIFGvF/8RCNMHnq7w8FZxe8oBRs
mwXjaV2nTM1isdUS0ARzhSiqMY8Yvoc09p6msHDhocGQ0ryjljZzaaDQ++HLo6kc
+tJVzY1NLxTsLmdZJzbn9wbGUeMObqcRMLHESt+ruAGPPb6E6ucWau/OVXzQvSU7
mhCeoFtKt5uttE3LiataDfRLXvonb9qSdr+r5IoZllU20IBqyCko8i5vXhHi4pOP
LydCbdrTQv5DwUIfi+EjfNWRg4kZXMD2z4soKNpFeONHvNXtu0Rzpk3WSrE6QIM5
jCm7KhpfEoofJ5ryFsmkKzbwuBXI2cOGa2CzYuluHkDgrmNsE5tLpbgYe7ALJ7NU
36LtqHaKHjdj6taTtakcEOQRzGlykkPkmnQSSLUTBTIeux3OF2XnXOHcAgTMd9g8
3zMTifaBKn7PCC0e5jsj4CMTzQtSirNooMTzweophFQ642m8aE885oi6QnO/BrKD
7yULy8l3L5nuwfVkicuDwWu1ZrYOGSNVJiphCg8+B6bVmV0ElbeQhYCLnHvvfV01
2Q6yptUZvBSnlzwetsoMYNByCdQC9jgTRIYoFLwXSIA/1OGMnjhztjtf6FPUmpqT
gxQzdaSOrCrb4g7GXfqebYBkrjr1QoQPcNmdLMrY2EYuEZxMTy1QT8B7PQZ85TMD
xBBY6kZ+UvF0hXdnFkIUthk/KcqUM57Tbi2G0YenPNboKBYaxQGl9dxZkfqI1g9y
mGMyD5e4+xbF4f7oF3jGNi/NVKPCN1eA7m33A8FvPbDlutpgfAS67/sbLFvGu1IE
kaBa2AhxI5aFhkrqyhcBuHjVpPFOc0ZZLX41YOKYlSMAteAPGJehzb+gxccinRXe
QHVluBOpv2AySquB9adMKhWcq5XHlVaHFQ+bt38H/2vyHNDyuVj0pxUITrESbq53
R0trSualsPitSsR2cY2wb12uVUq7BrmcNiTVLN/aEo0lQWgUW66hr7ErDhWji+5r
5+gvowr8KUR3fk7VzY15HL6kR+caKVHLJWR228xQ15UYbCrMQQK92p5Qz2rTm975
g9/BOwVXfsd5wK1g6mQw3dRlXOp+EwuZQe8xdGi+/d83hOHvhtW312yh0+zhqgwH
0X91uu0yiKbQdcxsCIMlXJ+B1oAvc+2mrH3FI+B5gXfcKvR2CDzOBYjHByA+YS/d
CzTx6h87+JGvkmxN79aeUBLjJC6ladqR51rGt5/cQqZ19J/iM+YT2XKXEPKxbxoC
EQBqrlsmJImhzK5TeIanC5fd7PQbQpHVPe0a84/oa0Xxhnf3qyBGWsYmTIEG/5DV
8zKJ7dxo9pRFEHZ6w9TYi4ypqgc1iPiXblZoQWAm8s9Oe0e7p2ojkBAVFqIUBLJd
w1b99GrFzhXmcpPSlZS/omWn4NS1T8ZG7LgV4Gmsu2QMHzQB+G1IxFZLKZF6kKrJ
17Pg4V6fn3U5TN1lUryBl5hKWKHCYVVgPv0bLnuDgJw87y6CdtzjgL4DOjwzyqXp
rMkYPjv27Y/CN6j+C08pw2MmJW7GLrXai1g5PlHrjuE2/zkTYwA0WHVyQD55d9uo
8vsmWVV1Ze3dLoJhJWLDSK8pNXP9CQ3D4Ol9L8hH9iBUBo92Ke3ZJhU6dhF//vVY
GAwKS4XgFktmVBXZrUCVE3bdYqbqNmmdVNvzxSZFD2T8fI+fauI/As+C2pdlx7Hb
UR8y0yQttuq7B5fgxgXOFJz7VU2HgJ8iqpLoimv3AHgVbh4YuNJPGmFHRoV5rXUI
lbDx3QvjLaBSZrj2vIedPqBWZs3crYoQaL8YYnZKOU2im7UivxSRf2q0Igo1/cpZ
DH/xNCOfOIQ1PDGDuRC0fpr5X2OsT8Mw/a3xcCds7/wO2LByHjF1sody/3Rg5vnI
EfvBhowc1Om4EkZGv7XYyK+nTJlI587szWFx6+jRkgrGyRal6Ql80fj9AaESEwx0
8XgVqej3P5ahfz57pWEOLsI7R6uQh7dIA8XBHqnUfxnC/ImZ0fg6PFOB55lLeZwV
cacjqnaj3xiS5lk5jF9TbcLdnlgbgEiUbYgU3WHf2wOexXuT7UPx3adOzSotwXda
hTazshvoV0YJepDU6oBoG+ZaM7S8UfJCICldfVd5OFKGg5MqMiFmiaglw7tWzTmY
3KAelKgTKmc77c936fuzdIiq/gd6n5luC74Q7v0K/mF0s88C8kZQCXBQfHAqwjdI
c1wMHV++ix+7LbuNT2A+3ye+xdPAt1ueGQvmZSybya4D5JCfa8XEgxscSAmOyY2P
dbDhVf9otoyQxfwvdXptX2iT6MTcBxnn6COwKYdpuOsNCDXKJ35x7OZcR0oWy/Ic
Nco05okVAp4bo/WfMdCLzzd1PL3rCRPiSCyd/ffrYIZGz9R/5RALWBwg3gmQWhIk
fhfUsJF2fTIoiXcq73amwiXGAL3erLsyzTHeCJlGfsQHFRIW9GbvJnQj069huMJm
9WlgaBjsEFkEm8HJJBLPfNbTsH2bR2RbR2QFf7RDJOsuSoxSxa8JbnrimYIoYqlc
EqloCB8K9S+ohlhBdjOVPK4ilMD5FFeQyWRqTdpwSrsD9ASrZozReBz2FAuW6l6Y
0T88+0xRcBpsySHJhraQVjygt8ASUIE3jiXym31pbvnf7e2lbVO3w+gAgavU1W4k
XyG2UWFiJ63j6cmGwZPi1ZA7vORWYQlZo5poeghKNykX7P7HGV++0QhGFqbNFp0B
voNjnhY6gbI/IOLqV16O4jQu/cmiMG8kVuvTSjRuhyP4WnzotqL1zZZeRGGnXyqj
9E9gFGepMCm367W/X3ERKxwkV/g4/EJ/76lSCQ35UJhh2eQpxMQbR723WPoD7Hd0
8XitTC50TakXKmet9UcF0LQq6WVM40yQyXjrvVmM5tQVVwKb7PV7OSg/5OUxNd8V
AMlgeMrunwpV+G5H47CjYVABwKGUYRdC1uJX5ntHw0OF8n+SAiyRgXKhoIUgfWVG
Khr54Tfnk4tFg2nBDipoEJrpxySml/oPHEo3UTyzDzpWsWvlMzfbAeqKRKRlDkbD
K/K4KrK3xY8ijVAJZycTYZ0Pnl0Vph4cM+kOToAUIcrY2sYShEESbsUY9lAg/Sl8
78NiYto6RcvVyXs8lwB+uEhnncpJYg36ibQK/9TIwskNyndDZvsYCl/Llx1n2cJo
6eCpUl0F149dxiDtcfGdef0De7ef8QBE/b4k852xuAdVInMVsp8IsAxcJM/HCDJ0
K1kKgBIxCZrv3wcVO+4qMqUUFeeTh9is37fgGQVqHo6wtlEzLz3RGyNS/hg42ckW
MJkjnFyisLXhTu0XjdEf8RcKyMfWGecn4+08pZSua1Q2mBjfCoDY+0MGeUJjrVIS
niuaPAjJL+RLtnpWW7x9sO5A56aTrMrpxGpOlFz9F8QIdTdI11C0Ywz5FMiR7Plm
kFzGkm5gsS6MYGwMmc0Pw4Xo14rYMuGf+O2ZkrLfxohyY3wpgMsDFnfPyNZnTMCI
N9550TFdSb7u66qIiJ3Pmq/lWhyZ7sWS6tCmvErJfhvm/hmUki8IB9kZzwvfFdT8
1GEJd7hDAglY3qCcDfCdCQZaKsUVFmtJbWRrBDRSQaa9NZIsRb2oZsS8P4t2K5wm
bI3ioWhuvmp25UUQefsO09f8U4d5w1l9rwiov1GqJKYScBIUb4QLUWdSTOkyRfzT
ESpi8juh78Uc4Zssbb0T48botE3fQw+6JbNrt2wMjjcKj/1YaHIQwylClajMJ+WO
tT3NlNsgdPaggGUpdKGTOqpBY86vAHgHLIKQ9TCNC1jvS2la029hzGZvs5t7Nkgd
fhllaPsj8BxrSVp5AJRK9+25gg2zRO3SXl8MJpdii237vpHSJGN/uCxvrTrZdNZ6
FOcrY1KEMOx5D5G9AUGlUXWR4iQEURuWNanROaudI/K7VSTIq6F9nP2Y7GvY0e+M
XETQuGyYLoIZbmgKaVx0j/7ad9dSatX7SfwOCApEd/RhdZPGuKppFyKrPbI9dshE
9VmgE1tEhtiMrOp5lWNea7+tI0TX3Hxjz3KEj5On/lDMkCSAkSn1j3vmgI36t7nW
BkAGkv4kF7p+xGd8S1NiwQCd2eouS9mWQGidNc5qATgKqeXzzkTsRF/RZhZ6eo+V
QgAmmOBOL8XcMfBI3B2bATuYEnoN262VsTXyZDANzeV0d7xOXL/uC3zdOW8WwCVP
b7QyfftJeMFQT/phJ6C7xiVvgU4KYGhRSRLkMHfJ0dRTGMwR24N4xowGMNSKUQL4
X9VaecRGcl+0vqp7iPWCA59n7deXH2BH5NXJw0zUtxr6zVNdme6VhanmvzOhMzeV
tDdLz3VvT9P/eNwk5NYFL7tzn90xBIqlb6BBIR32AqaW2fBI2+AN1iF2hg4yWQrO
k9TqWXZxzyjZpykFII4ErRO7EWqFc1/LcF/1L6P7SxksKMk8y4+8lHsBeUOy9lIJ
gKo31WGT5ieh52H0ga4lYE7ZAWZdtGqLNPOaDBqsfrarqbdyCu69BE+o+Fdi8He3
IdJlYuWGvbaaGL882Y0lZ2SPk9Rd8g88sFXzDGZq69uNWl17n8y1G9t3w/9Il/0x
W+k+OtjConzR47XxnXQhJFUHx79MLeeHJ+N9t56TkswFUC0Zej0ejCWZ5AsJEqkE
XiChtoMBz3L26wyuz6JuQYHCSOChPNUkbjbyNN0TfXPzC3JzvUFy45NG0MfkHJ2P
diQZ00zGWxUtPgMq3tUo++3VCCebPEB3b10eGhyGtjlBPYezp9J3shuLwy0/zE+4
3LYCST+2ANyCjmcdCVvuYIxBXj/sPj0DUXzPU6uV0EGLL5aPr4m90cNctfi6ZBVK
0N/mjn90ZSLRub42mImzZ7Ci3FiuFPkmXG28719B8fEYH8QC/SLp9RRSgF5tey+t
9+8afzG2qD5EqX0Br2prT1uw3Oh3ReepSx8af/wPV5BXIVe8IvhTOwZ+bpvdAIyh
rwUZT4M7qj1VFDzki7I9spdhTPwrqMYNu3wTkt5q5/EqCJU4kd9lnY9aHfPFpJAk
9voFwWJR/y3xFjXRX/gHmJiB6D4cJQ5r0Jkb/kPYjtx/2th2ACbqD7dYHV3HHm2d
9K8J9MsGLp0b4brhjdr3QoTOTKMvwu4BsY17adknytfag+yIt1DD88vq9eDhIl7A
8DOU48V4PdPZ0otSdXueoqhVqiBfpoZAo3ZrQU/jgaVdrIwtfNb6tdACWD5gMS/F
rOGxInLEPO0S9WYb19G58c20ARr/16j2Kf6+DGkkjLOdvW4z7WM7605j+0+ITYay
zRutvF+R3MVGkLdqpgb5BNaLIGLVFzVE8spXQbAG5+jQYn4W7qCWRq5FU6M1HUtN
H5cCxLmwAbZV7ZT+FAp//vaYscr714Z9J2dLqfQM+ufcD4aXq3W1C3uv9uQkgtDf
wLjSRWWvCQEpGseb9uVNWFDtE8TwMzRRrD/j+Q2HJQNo8pE9DtvwvYE/0f7mCxai
af8ibyGsAfZuwTtFsBa84kZQu3rsuCQdK1xQy2c6VFVTNPwfpzrorEACJmySzRQT
+kS53g/Eod6Wd2vv973rdtFEaBdMCG2JRKvVSSVA66YZt5KBgEDXkbU0USo+solX
aVF8tUaF3CSqo4628uvnQhihPOyyRp9Z0XphWwBwUISMwI8AcHtYnljo3V4h4Tpe
fmMz0bWBF2dUWdDM3JdknCrrZscbm9dQEXvVi8Y+6YHfLUd8V/OpIWLKM4lKIo64
1SMuOGjmyWwgTnUbgQL2bY6yQpUj5jIMvZRuCb73RPQSOCe0w6Re2EQp9D5O4cAH
rQpykt7zLNi6utMvAVO0i/amg7BEQeTvmSv4Qp2RB8OnYcgAoC38XhdVSicUwwEr
nRe6/md3ezx3uL6tmp3s2nzJIyF49fFFJo1PpgQK0PqsDCPtpazGBvAML9ClXLWU
9lVMM9XYbootE+U5sj5A78dP4KT9yqsDhIm+i4w6c4a4nJYteefSlAeLuWpc0t8y
DChRmXCPxbJLA2c4IBInXGVlbNqqZoW2e++qX9SdZKJ2F2G3bIrYHPcNphA/yna9
ecxejWRBybihJZ12ZE3535yEVq9oghlJU8hfEIhyuOnqzhumSe/oL5HyUULoLn2l
2tya2VwTgbQYdIi1DUDGgF5yyf0ZIxmuc2rhaGzPdUIt/rL5vD7METICMifa+l/k
3dW6xMZptHNW13uGcmJhdrDlJa21sqKNmwfactH/lTrNLqoRvcj70Z7pzuY4r4AW
jNa/QVdUf70cn/49giHUMMI05KMOYx+LKe89New+jTCb+HuVvQch6bfQAa81pUZ9
DUOT5SzWQjvx290GH0waGyCQBZ9svqH0lcAbsdhw+4XyZL3uqxMm7mOQn27DWsXW
YYb3l08u3fTbDm17/H+8LtbO+DO9J8ccYYRFbvWq44t/yaoUmiBRPuBrN6V9S2pP
X63iuUwTby+l72IQLaUYmYZLzfuUK1UgwfpsOdJmrFH3OITUJpxtoxMXxTU+OpJM
CaDLfNnFO424CRhoFihVlwV3BpM/ORq8/y9XAqbcBECO/id0GaQz9tg/VfEwcNzc
csq0v8DMBvkYU+INoDJ5KWtNEqM8yOvdZTYzcYMURiS515JBl3Al/8dz2+Afjo/s
nV+uMTmTnQz7IL7De1NCIQW0fAFFMoT9+/olVDvv5MQOifsPa2rywh9HPA2l7fCG
EGUd3WlwJNXxl6QSncymeW4EGGwH6UFVd8o5b1frV+va2eSvBvn9lsp3EGzyTQC9
X/McxXD43DWQIc+aSKtMT/XpvWT+QSmVBU2ypcd9t4PhVXoLxF3VM4CDgwRGPyB5
S39ZRsM1jMwnbkqndigio+NmH0nlZCEvffNbGfk7oi3wU0YCynirgJnKvkVkioqa
laZJniiE4rhKbKCaMit4Vg0GqnC7FoNWrk6fPo1P4FdmMxncnjnH1yJW2sNCFhz6
Rz7mA9Mv5juPBdtmLUeaYOHp40qnsiH3B+sGTNBBW7ftpUD5ZfrRYRnH3vMroiQR
yxB+Vg1r+A/GXAu3rD7+LM23g4frHNltfWyIfIh22HPPy1aeCxdNfAMaCEzCeP5h
9k9+51dCrITw0Hi6DDVrxWoMYcVeS/x6CfFHqtC+5I7T8vvYP6FEWhH5VCioMdF4
KFOcSLja3RrNAaO70KMdzCrxmkSExGSt1GEiMJ+xloXP2WVCQIE76nAT4/GhLe3E
sk5YH8iD63JvaVn4384Vo2NttUu8ttobAvHcJOMo6t58GypWADDTGbBb0gzRJRB/
D1pydELJ9ykJpiDVsEj/4+JlQzaCtiylEPZF3n+pTJDRCB+X10RWfHSPwaRzZR+V
YM5xOPaJ+Ggg5Jpg3VOqRZpozCb5I0mKX9nEwj26BleSBx+AQz3tWlHVudwpoIB8
aXTMwzgvWf7Q3BQknog4j6VM0C4J/5Ino9N4DbHaQsILerUhVgMVJZksUotMdAB8
SaZH4G3QAcHSGmJyIrlx4QI9kSdYQ9Jid9h+A3EUj/1QQcBLT3oE9jNpRiokK68s
Fd9CGT1w6CXHdplEFDaOsOOuSbXMxqbFLuwQAyQCTIH8iyOgh5tIAUnCGoh4/KRR
3YmUBRze2A0fnoFCJghfrD51QUbJYcY3vVBqSJEE+rri5zfaFw2Kqq1cMfHdtNp8
H4FQ1w9U5l3dlq48UQw63fMH9/TOc4m8Vv/MJ0ZgSa4Ax5uCSb7kX60NqG1hr65+
hZts5ncR+3XBxY7adnttc6mMDv0V8agGJCZ4Iik9niTlBntXaO5dQBSsuYEuT5nU
UG9CasqwYB9Cxq40TW+GbC9xmVqlmYbKQZfsCUbBBoEJ9CnMzwlb9hSnauGoKwLT
gTJH5pmElYYRuqDWuD2SMrRU0fGwc2z3/XzfADO5AKdR1FJNGF39Sm995qh1CQpx
0sII3zE15QVFhQ+4MCYNN/2GrGDjQY8ptH4zfTknsFRWtxMf71XEFJJkgo7WHkYP
JBy8ESl2nnmLM85828YtG5YHHVg3mZCQPMnSK+/S8suWMAlb09d4ItvoJJ4bY3zX
vHfDnQBznq4OhfDWc+PNhQUf4WC2Wk1Qp5uJFY2UqystM8NKDfCNymXX+XmFAz/+
194O9UT9YZwHwcnuWgy2j04wBRRwMQ0dwegeHIFoqDtBT5Cv7n3X2IftpFR+KBV2
xosKIV3f0AloHc3MUoulBeDGkpLd64aUA3Z5Kux+xzxQtoW7iVViGlv+BSctKg6G
qy9OCQXp66NqlN2Vb37KKbxvFzzGwGABpQQc+GwiPwrzZhLxprXzBa6r1WZ/5v5T
eJtNWrh7cyszz6am7la52dd6O5cuASew7zHuewwrj+d5fv1c9r66Luy/YLKwcPyQ
CIKVvTYrb6R/7wXJYae6S+TuPiVTCAdx3BDN1JGXOtAcmtoJT7JeJNEGwNueherg
GXarnLLPI9iVC6WNVjOEF6LxTT3XaAlkqshhSoA9nw1BC79U35vN67me6VedyRWw
/r+vpl932KsqbDp1KsVBVDV8C7QeBUalfRsgwj2OLiftFNWCj0Qvpj1XNZp/Mjvf
ik+8OGeBnEEpQGE9EMG7B4d9E1C8apWlYvAXEeiuyj1YOPoK1pn+hkyWUDuo8kPk
/+iaJ27OUl5oBScnip5lsfnzFg+dorzatVeAWHQlOgFpWNLZIeucPg4jLt69RTST
DnRtiwmePWqV8PSJ0bN7kggqAmoR8Uiu1IyJHap6KebRyqzs0sm67Law7Hhst+Jm
ZTowhJnl6oklH6aHPeL46F8c3VCnEcAaHqPkh8Bd/XDkFlw8//GOR6OcysmrR7pD
JZdYzxdWygWpIws9Fc1lRzlKgklN0P6a+OZduFA0/yIphVlZr/GHIwZZets752Z+
MrFyd9xZovLOHi2E9FLIhV4ZuBkJyAaz3S57k1qsEMcDseQBJeQDxHQq1GfnU9GB
OYuQIJHNWFgljJ1nZSRb5NETz36iZ4RbEsR/Dz/xSAQWVMMCcpMzdsHUOeKhXsTb
B+QVuoeI/RjfR2h8/A5m5/n/agUgBwB0fvaIwkd6HYytGSOiKdaDD1nk1z31Atr6
neFkyOfxv5oey+187ot9/RnvWLjz+rpaC3YPbHTR8YG/SInR0+3sdefXPYQFVxJv
GpvbSHqUuzXXlG+Q1uVudCC8Jvyyu/grOrht+XG3/21K7IvfvjRhe1uBdGc7PVeh
X5mLVHXgZHMKgaxZl98RQrXPHrlGTJYsy9BOS4sgp5LyxDWtFoWdLjMFobFJ0kEd
EfSvOl0gT3nMw2m6jKQHhAl8fy0fYUUjMssJVjR4zJAI9H75VKee38BAKycDtVt0
dd3hcnk0x0lR3pw665t3i+a9cBI+x7Xujqw3j8U/yXVZqGe8gxxByMVlrxU2eQNJ
MPzceM21gtEI7ZqFmDZlUyco6M9yChvgYExONKZEmpjR+qPByeoRSAKVeSdV0Gt+
cQLPxYN/kTQ/ldVHNGVEqBQsFWJGNngoUVldLD5wknvLUMpZf23eBsQjN573Jzip
tsU7rpub0Z2A/X+kbzuBzx66cVFNQtJ6eyno1vQ9WqO0Gwqjypo5o1r0z1ZAxVrc
yx4raIDvYWgh4ffJGsTwGVwyIyDk1+7GLMScQkzDc++9SxpEtyjf+i30K5lJj5r0
gXA14UA8sF+/BVZEVVOFBt/1OIEW2cKTtBvTAuXmU51I/GIc/gL9v2yS7aVnpjZz
Iy9owtgo7/LPCazeNULOSiIyJW1XGhf2jJqb9OE7kVG2T6i5Nn2L/GrAIhGb2qiX
QGw8GXEbWkHn3iXmNQtN5nvrVha81GelqC3DJeJSHLm2A+v0rOI39yfwF5gFssNV
+iERk7pLusBTisYE27ycrIeF8Px9mvJh+e/tw3ZsHec9H/VPiNoeCbPe1Gkiu3m3
pUfMy1+GRGEE+ooHrQ9SulV4TrrYCVWTVyCb10AtZTmWAE8D3YM/FsN6KP9mYiNq
UhBJriVyUDV1ph4Bc7cq7rSHeo+yolmGD08Ng7kBv1X2gE5dqodnpAiTr6BPvbjx
RPsiL5btb8NUsROqdJ/SgEEfikbu1P1VfCTAaQz7/XjPOv3EJ3DGMWM0RLVwe/Rd
4B0/REp7GY9fVDrB4qGuwDfh6f28sKiR7aAqatKijq1eSlObGvYuhmeXdS2M9DlW
8FrRSEVp0S3fbweu4R2zfKwlEVDZaNWWOtuTTcxX5pH7ThaIfG54ymPsyDkrZKfu
uZVIsH9oPdTgPkNbBOvNLuaw8DQVAW8qmceX+b6lswzetwfuCa2PgHcRYi9HfOcW
`protect end_protected