`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 38064 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhKhfkQ1RWny5iJ5zpOL+J6n22O/UCwa3pitUyyRK2+2O
+nk3oq7qNLyVXq5jOjGxRMFyhObnOO0yxDYfjVnz87mQica17ynm/Eo8Vzxkya4P
pm5lIyt+yveaFj645+qHCjXi8KQggXJySK/qOT5+FVm6MLMA6jGyi3dHhs9857cb
8BilGYT6pWZFohWPutpbhJfFBg6xuDiA0pDGrMtcugOj4y+5zAA51o1jpGhYnk3E
U1GJqqL4d2HZWc4yVmvFEC4ve2HFyqAczqzXM4xCp4v6b/As1cl51kjJDpZiFY0I
OTnJL4MjcDW43OzkLImSV7m0hLOka1gufI3O1ZIVlX9EyE/yZWiR2SFgHVIFohfQ
nBxFrkA+crRsg92A7UXFuxb7EAJqD+OIZ0RZZ5gpAC8gMXakn3NoO93gs2rVqLxY
hg3Fnd8NxHEVtRS2IuQqGMPzztuGuuqrVKkV1sC1LKk+UlmPzoI43TIY+jxMTJAw
uSiKn9Qmxq2MokGsR6J+J5ve3LoNlfSlLg9Kvpu2JpxHFALBkHWbyWjIWsN7JwNJ
bc39zdYHpEqfgZtCvQcL5jKHPlZVTvirXA/wZEx7Y7w05zkqsN1ZG7wbPDZqzGxc
zf8IRct88ShLEvYGtPX9EV0XGF0T3Ei5I6gVV7JM4H6dZcFfF76hrSognYXSzhTf
QPWN1nROcR/+Z684MNtPkSySWfymlXrZAoCG7UIgfv5XenmztGgYfnj5VZ4tTqNF
FppDWuqZMWdtCNNUFXK1nU6ZpywGdS//5QYL0gLUiInvI9kNquZIyq8Xw34r4VEx
6U2Ck0ev5Vj4J2zopwQ0fGhRON5pH/B48qWXO+tmLVHIQ9pwQSmqN0JKi8NDyr01
GpVNe0jnLAhQ80dAE6PDj/1irKedn1PmZc5Xw2v6c9aNysV+WqXLDYKAF9V8Bq4N
csOip6Dz8UzNTO2shqvB0mz/6RGnr/ETM1xsW7eZ7Q81a/gvVpAeEE6s4NWY3nA8
OlCiMYs8gl088Su1WUrKnGXdDAZ7SRxpOKw4vkjxJvjfWaj5cTHqj+pBDUb7MrLK
HuvRz6Rtby66I7S+bn5UZEiMEbSC3eEcBFlzjQBIjkCaIT3Pa1Xpjy3juncv5oz+
Y2EHNrjgb3ikOzG0on1XrJ+9nOW24XDi8ar4wTIWRiouhUK+rX8pier/BeGJvKxL
yl5pa2s6KDywZ3pL5MCfzPirCShin+YC/T69qkWuXRjnhWhUsWc/cw7okgSsivaZ
yPD1MCjEBDUIO21U8nI2YIcZryndBQgXQKBZOMLdeVUzxi0BU+cO/cqMtA/NC0N9
vUn47OJ1fAoDpplxSUuhrzw2gfcGGBqRNim/IV3GbcOIFPnBUSK4MUJyXzyVZmfx
ZmGfz35ALbeAE20ZtbAI9o+yQ8r/2ZHjE4oEBtWBKs4B1nwpGyAlMvB9DY766r2s
+REJlfFVBGCbI0Q7GQpzFIRrOVBQv/EDkgy2NKQRwPQCYwWOfq2lOwg4xEvbyZ3m
t598ReNYO6yKgwNrccc7qhuB/vJ6Aw2TekWI24JF/339RloRwX+EioFm+bz7TBt6
LYcgVqfkvbYE3M3KDSq/zddABIUVdHMFpBoOo4qDWiNG+cu5F3vVclke+B+MTXhv
LhUFUTXabSGp61EC8RjSDeivRNEfAiVF9InYVzZAKrFtZ7w+kRrpEIDI27aMOt4O
yYeNYMFABMSv3iKtWjJmAyp9eMOqBVtVd7Zc78Iyb5aCqe/XuzpkBEcJJM7xYsJV
J7d51LpTeqguhkEzlPQHrDAi6mToJgoGpTiUNWPPTIO1/jMr6oV7ox/Y0MkH6Cjv
9x7NTaG4zpNvkdlhuL0p/UVsPgdiXm9YPJ2ha2i5dyYbM6eJ/hL9xayWac12GRoN
oW6+Kpw1aUFWccjmpGYzRqhiUT5vN4ypqWCiRfEFnYZqMXUhTP2qbhHIeWB6RIZ4
h/sSSKDM9ozicRjRN3++2NDb97GiZVqpxZOOtDO66Vr98p1oKGtrAimKkwvvtuLo
fObe9zwDF7xe+91aGV6lIfenqjxMbXwLA+B1JyEc5cN75NiHDcnCA+BUX1CGwwNQ
staPP9Rg3T8LmVChq9hCp4qvTOFPzENPTjp4cATnC2SeKUkYdnzI/TOicPxiNCdD
cMWl0ncGrOpIvb1PFNEpn0qujidyFBwLWYIfpD3kk5ddi4Ty4/sRKMoiEjTvAD0e
ay4GMtaP2h8GVhzmAky7gqPxQ6tyGWWpFPIj3sIlKxU1nxyfcrSr7StVgCpesuw1
GKrWasljcivRgvR0ivJNy+UE3SV8R7Afc90aN90TYkNH0jZjV38w0wXekJexjnPf
UYgHntFQxef4QXqzzjFAP/5ZlI1s2E8Fj7RacFzVJaYBR6FoYzMJ/qF0zZp1Non2
gnVZkP+/F9sI+h/yI0bo0tROsvePhzpBkwCA4VbcR3rfCYIKeVgv8ne9SDwqIwO/
EJsTBIuX+r4kQ30MslhZ4E0kb4DGRG+ugFBDe71aTZYWESWkCQnWfomhx1Msod0V
Ik18H58iWQv/8vw7StlwL+TaNds5OW5LES3lS7PehEKbV8xE6gCV+V3i+Fc8oWuE
x9nwqyOcbvBvtWURIpJv2e5tHyxUjJYI6HDdZEHq60oBSiIgg9z4WsA4IPnpwkfz
5LdsOgKambmHtqAy7YVe89L5ewtEc9epZMdu//iusjYSor2tpHwxZ6miLBxNEby0
X6xsnP9733A7C61qjyvi0vmYQF+bJJpM2SAY61RzcKLjtU6wjhH/crAUaNmFszZg
d74D8gi4/HPXiGZM/AM6/e6GZO9cSyAQAUv4rGtdii77iB5k6uX3WWcYemPE1/Po
hcUAzaNPV7godZus6cqcehAlouSBa6+0UrcxVmay9sVn7ASW1bvWeA6z6ovdV8tn
Tp8GaMT3uZvv9SZ19sXtzNebzLX19wXxc7Tvon7cbWLRKHECKJtfkdqeVBlZs0IA
lKmFbY3CYccSM3/E2gHJtyohDoJcBwyZx+f2T7uDUszg7vrYDBqPj6qLikdyn5I2
vNU/Q7/dygQbdBptxqmy89R8mCBiomXsBiBJoUOi1E4mlNrFDjzeb+vcYSwYkkEB
EAxYP7B1tFYXLw5IzzekLBONPfV62ha7JpgEsaZ6BIuWJ1PVEBYegETIdT5FqC4V
CytPkpbZnovE1qnlN6t9cXrh4XgQR5LWxDM5uMMvxVb0QwyX7IRq5mcL6RuM9Trb
qGTSHL/AF6bvWlt5kvsiXQUdWlqw++Axpa6K7zFrqPlajmc3U3isuQ8G86+AbaUW
lFBp8WBdxcnpFUp6njxssZfByDfdEirxXobZBDjEBjpKfqmkWt4YWKFsMYAP6qID
i/IvalqDg5WVxWUIKGx4A2wOiXqXb1QgPYcam+bTtwdDrPPd8oM7YiRsjj5D40Ro
Hv20SfKLNixXolv9PI4yR7euWiTaAOpQgj8RvJqiKXwWamwhKfAPfzJENLYXkzFf
F9X/9VozjuRP3cojryWS3Gi7znXgf5IVzDjuR4IKpVVIljhIWi1msV1tj9DgCX1a
AjuMe5RyAKQ0phK8Y9eH5Wf+bxicSUrZQtgpQk/vvEFIpiNK2nWLAAAmEX1Bxaf/
hvwWh5bCdcovHHzpE/zoqqxnM/gnHs93UC3ssrEqgW14x3czi6J3lYdknAMUuCRZ
Q1xUty9OG5GYQ3KnPnU37Jo7GcnYlzctwbVXiehhJ907mFnwImAMcAM3n9l7zDf5
PSdM6w0z4M4FsxOSuIJrbv5G5YwLIjEXy9f+7Rn+xT/omdu2TgUja4MQC0xxTmBs
X2maS7HPhA9LZp7hsehbFvLnDTclHqzJOynbIwK+qswpKQX+O2iQtvb2Ok17OCS9
dorhyeKP4pgG6n8I3QR49SNSTAMUSYpa8Qae+DdxAJH6NX9MX8D9Kr0yjrxf4P+s
3fp0XzGuXdtzYQ4bpP26Ve10y0ih7wDDrx2ExKV732/VMQ45L7y9eCMLg+ch5vpe
Cskv7OF+R/+NRZCzQyYcw8Pi7gVdDXJOEwCoQ3JfpDHLXgmw5VXqlZ1XWQGffwh7
H8g9y0XKEDQJHIDO0uq0+qdb7YuHmLD4FPV768Y0fNNKA2uQG6TbBM2XDi3ShrNz
iDTdyFGHQWMNcm4k/6QwNUGbWv6i7Qp5lcecP7L36VRY/0rK2fB30YdyXWFfPCVn
qBCBVT00dYeHtfHXgQXRotRGzQCd536WfZ2+6SmfGA/IiEW1XThOg+ZT7DFZLWZu
dCcdEU6VrAX49Y78xAx71neO1AGBmIustuRZSVSUnD8voeNPKHEFxPYERpumleou
mNslwzeTwVyq3Jlz4eWPyUU0Ajw3GsGpUQsAWaW+6rqrYkhVcfZYPiwMaGxzHLsC
J39tpOGWYzfCIaNZyrmrIDhUrhuYbTzwVuVLctf9R6jRQwrjV+i+InwkBm0Nh0K1
PbzG5vt+y1T8PqaScLanqAW5nq5HQvR9v2vzyFVEMXU5Mmg0H0xDcSBklkODwhm/
SE11XUvltH+lHK3La3iYBrnaEnZKua9EVGVc4NnKpuw2ao87pq+TTLDumzNm6L9/
CpZb3Z+7O3HC/r6+im6dpz6ZgwAjdHq61M3d10VHDw+VcdLDyzbRDlJ/c7vg0196
LXBcYK1TYd1QBaqioUT+LQnZ1bou3akc5SwGAKrHGuA1DcQTBf1e1ILq2nOGPs9T
k49U8EYuZn4SZiAWG4drK54Py8q/nFV6nRj5BdyN81kSu9zSnAUC8eB2Ku514GFe
mAdJmCgiSqBrcIW3Fwj0BFqwXwgepnVH26Yy20qBEHXMF/tcBiA0AmJ2x2RO9r7C
NurfaSJajBAWweDkWnLby7hnwZNg84y0VowELgUdYF2JrRtWeLgjuKYhD/3RYVyK
zm0Emc+0AO2yZeWRE6AM4BVpflZiU0jaY4Zg5mbA6rerZxfnWlHMdUb0xfQipSCu
IsoR84iF5u/4GwB/g8qjTAcbxmdlDNIyUuQZ3+NUUfEqqwI+AbyqlRp7QU9bSBqx
dfp28p3dgvJDfy65DXLG22V535k0PKayhftlm8A3GCNs8ekGRfDR8TuqFKptk2Qt
0cdyKRr7xCIJ2l3v9oLvLbudYkYbp6HH47ZcGIlaEtjIuhueZ9dSq5+11rVtyaaf
I4dBI4idAUpBjMk0L4pFQKFedRRuqwcO+JDFUnZGxSSQsMR+oi6DUHFOI55TuJ36
l6bDZ+xWQHMmMe4TwbbjJ8RYUERjtCXmtJgIol16yFoXdQvTDGxChhS9j0OHZnP8
RIn+RJDQQ4fw2AtwWIG73WkBR7uqi+Pu37h4U/Q2nmpvh9/rlzJ2ujb+aVZ0IFFc
DJBfkU8joR4/IMyt6YWRHQXHAGFNxR6MFL/2WyYxq51uDe15zQ8fanQl6+UJyi34
TmQ60quM3fi1Uq44LN8hDMsnx68w+nN1ArbGSujzQCLpRjGwuEwpJyblQcIKtRfo
pzt/v4BhlGK6FQaqS13kprdg9idhfntodetM/AWHSb0tnDjWT3+7thR3Cg0N6JRU
ztdMPYDw73br578J98XtCqlSH+mdhVe8sUkNS5uhtKeAjQzNhARTFQEwIdAi+Npb
VXEtEff84Qgtl7o61azmdHkxZM9pZno2vROnGVRLrhysz7qIs3BFaNuAn73CdCrq
2iGFSkXciCwHelLm8vGCX7f96jDyfjZpThDKMJNe477ZYMKql8l3ycyjkk/OD5AS
1mAVtF/r2zKXEMW+AyPnvSYjEVdnS0M0WtK2nzWJtmI/cMEzlJcbdLzITFvasjVR
9FqyRHARww/J+PUSRrOJJK5RcqQmVoG2JleOVFZLVuqVI+LC2SD1gaHj6y2uUovV
ydJctZiwmjjjGoFqcPLvbbODja8Gf/U2eb9E5ufpk+sl9HCjExXiJxkT1Uf3HQrT
h6Mbr53KwHo5JzAEY/TSZJy7Piht1stj2ow6OlyNBVNrLOjhMfbz23pvEIADC3Iq
+XqPF1x4oTxv3JBimSAjYA/vCipuudseIzNh/M7OWZGS+OqRI79P5FPnA8tILvQw
l0DrzpmGsZpmqY3Uoky3JEayEJt18BC4J7hE8ftIcpiXMWXanqreSDSWDZjki3x4
n14WTQ3GNO3QneoKwrTjXpDFYuYVQ0TxCFHNkuxZbIaFTRIDy3TCjgTOzyKDuSJR
F+M9LY66ao4fvnLAZiM772qQhcDnk/Bq8Rsr2aoTfrqnkH68mJs+fOFq4CwvF5ll
DnviupkBcYTWnAMfbnqWov5EmGSKvd7671z4y/XxR5b53+K6Xm8qYRhjhM27B3JT
LlwsUtLfErLf4KQExFd4+Z7xtA1tPaz2NH5XEoHk3kJBZU49nLjrNrX4luAl9nTS
v70yzFz6WQ7l0QPREYQMR9es37REBle7uMlWrfOv7DnvygX0aHDLmnYsboNww03u
0ebj3oCtbLcGsthjWdWgrNFbB0xlBsNLSXLh+kfJsz2E7zPu+yRl8sYN/dUqNEAb
2rPRomF6lv/+CVfSlqgDI+Gdxb7TuAJ0cmtgD3qB4rJTKcy2PP42YtrAY6Ti1pzz
JE7SWJS8Njer64sUyJVkX0j2dU94p+gJsF1T9DA9x8vukJASqPlbrQxJwDoJsYk+
qaUwxHvPYNx2kheVtAXVOTEyU3dN9bIkwW/MOCDG6e11zQhVNDf9o0aMF+fYgPS1
atEQI+rdQDrYYq3U3rzufbtfsm4owuLAlj3uERVhNxvmgjYCrj0595525tlkIMZG
nnyvoP3AWmWDylQikZkxFYYMNaLMWoAFmu7lQwySu9jjzlKMrWOvlA4oEbLPcZbS
6FcRiU2N/6V9JblZ2JUHXPn+zQ84rT3hqZUAi+tZ8Xts83ldpDffjr0MRCZ9hVPd
hdGImBjxztlDItIQo9k5n2GO5oTq0vQS8tNyqfp1LnBX42Pf6rmh/Sg8PHNYFsrX
R4MgtrbN81Bz4EaeMN9PIuAxFyIN3rls1X42jiKWi+VGh9LBvHWOOCkU3Oaj+MEu
IpCg1Wb/r3ELX+b4VDtEsPOxj1Em14tHX128mW8Lvvh2qiBha/XT64fDuRNqeVch
1PsRJzpgmIpsNG3uAm9J+pQNdgQWqPnzRvWROaPczkcjLF1/XaqlkVwWYuZLAUrR
gdn0ZLChINuxkCVC4ILg3dPirgvXhiN3S2GkNT1X/tHnPyaMrfbec7jAvsPTUzGx
12HH8Th/X1WV5yAwXFVO15r00oGA0i9OFqP0eIm5gY65DIhbVdyCsgCy8qZzJjD2
npvBBVPsNye64MuOGu1KPpdFG5g9pTtIlMF1e+qZLsm5zUHE1sNEM2PQLG+nQ9Pm
T5ULirz68C3Kp5bHSqgCG84f5OJtmUVsmAYvu4sB4/eWmtUuySDvrH7qLiC6281V
QEOcR1isDeQmYDh10gwFi46PREKVuXtAoEUGtw/1wKxYEl6iVqKs3AgsNDpwHpAc
9ioWLfZirs8em1qXaXsG/yW0tve0G9j4Ib039tvCca39bGX8XhgEkqsZiYTHL1x4
I+NKMThKjrVb5OqYcZ93Yg7qJdmkwYGo+Cty6k6Znh9FePc6p5MmSgiQPN4YY7Ak
GWLqLZSBQci+fhldWPtnY+bvxTKhrkXNK5e05j4hPciHYxIjpuQR739yu08Wmot2
yZkZxQgp8HmgRYq+bcUwRxewUFP9IYSYC2NDt021T9TKUcfIRTswh6uQoEcrvnc2
unsL4LTgw7vKnrIx28MRq8iV6eVV+okG1BIyyQYZTYISUZ4/VGGVwZjXo929IML0
35sriq0wglyop405ktKtnq3aCXvanqTngfSRXAV92kweIk79RlKAJ3zlEJUEcfnI
mLGlrZuJ8iKvjbzycyh7rk7pa6hVpOBdTgYGgsxBmZtfPd06xQdrzZQoYtIFnycn
KSzM8ikm5r4AlvK1O/Gvd2EmIgP9/uiwxeA/hDmdlr0pdMHz6Dij8Ps9kVEvQiKt
Kj28/pO760MsUOWwJ1urL9J7Jj9cJCGw60TuJRMlv26NOUAVKGBLSOVSNkoNWutY
nukTbt6YDbhmQ0tIr97J0EWxiosMdw/R90G6VfOsEr1tSmNtr3dlkIzWjkbm+OJA
oISvcx9OxBvl/xc5gndJ1xgRccJYuF0Mo9D3GfA+qysyCfbPWF/P7WbmU3LV7vHi
8YJU93CwwdIGpjIZBlTSZDUB3eqfy7xnOE2uULGJvy7Ra9ScVS++FkqnmkZQvdtX
/8u+ffycZIfj3LPEViC9vAfz+nGBPtspwKC2P4/LDycTDdLByGX+dIh/GvYLIuLG
epb1ujqJfL/pcY+BHetUhv4vYKQuGABavMWnoVnuB7345Vhzgc5QTO3/OTH9W9+R
gsdJeVjNfzzTg4Y+IvRzQpR421KTStgQdML3BDYwgMz7+Ce7lx6aD7NAjD4R7X/A
DGzEWfeoKbosQP+OZ7TFtoF8ubSuzTtp60dx5pnFxWuAM8L7Bj+6Hw+WsMjLgBh3
i1uAXh0DjW+tq9uZCcR+qwcL9U0eBFsV43MNLwxVa/HHicNZEXCMKeNHLLy//iO3
fjL+nxZWKLXYYxAf7MLVpyjuGh5ck3tqTm3Lm5h4xqHLov5K8TbF76TrFq7rO6oS
5LILOcObwaOQi646Anouq03OmLqpdxdPH81wRqIlYEjdBc9ku+q4qlZVszsBoe8Z
Eit5b6UC0Zq68H0kPczHuTfU1F9V0sbvBppPlMuhVqZksktYbtCIceD4SkbjXF2K
iaY+JWjHw7lJ25havN5cW+RCUnjslSAZublRHX+04JW3Nj5Z/uORzo7NK/3T46YU
NEt/XQ+ldbeJrgH5mJotaRcsFgdAt4PmaF0WIfXKI9p6OKWyVX8g4deKNDBvXzaL
4NeooJnx3il+BfT3us6MC/QjlYrsJLXi4c1Qr9zj7zbObkgSAiQbtTvIzevwIXPF
SQWfL353mQEDUPDVRdSEJg7kQHu+N92zyy+SWm5ntdoffEpQD6eiV+BD7C/4Cboo
RGgqBP7v5WokNKDLEz9ZF4ZkG2d7j8DUKJMrHcJcpn75ahTKeev+SNMQTi+1lwL4
HoOP2YEe+Y3Y2OyIeMKfQ4Ixos16zKSoRYCVM1x31Kk9XAazBXkQ+vHi32WcS1Oy
XdWtcpVTLVwXQo0BcH/dBio6UDsPnCjrwyGMSw0YHfwR/gzW67K4qShm2KkXxnB4
58M235eTvNnd/ikepYoAFFP0mu+hCHI0BBnwoSIMRvVrkdojJTB+aJQ9FTTLvUBh
j5AQ+4osXQbsQNSxSQIUHeFgoBjI83xeEQvBRu7XPL/qJCVYBnne7KT4CNeKjZ1F
txEWkK4zlvSiazDNYYZcsi8rHY4RQo7nZ22v1Uo0Q+Y8PbdU+kFHE9l5lEx0VgUW
PpfC9kjt0BcPC4Vo+hH8xiq/eQz9EP0FBJDcu57x998keUE9qqpTd78dOarEtlTV
SLnKxC7CpiQMs5joEiRZZDRc6mHRRayDuXUp9JriB3BhU4U3CTAJgoFOP0vNziuS
agQx6a9Z+TJMgdScIxOZpUeBwg7HIiEuGBVGwLe2X+QSkYSfiYUFCXhJWBHZZRph
MJFAI3Z9RoonQYLQVap308Sz+wOld+1iZNgD8GD5+wYO+dOhOeKruQQzR8OFYOu6
rsejmVElzTZjKsItBzgEdzWXM4ILeekWjPyi0uUJ3JaPRsIq7pYkxZ2gYsXDhMLp
SCTO5GPUiy+VfVaOLWJ0p3zU1HVFf0ZvBlaKTAI83AaVw5t6SgKit15AebtHaSK2
9ZTjV5+IEWbfb4x8kSA630XPbOQkJcpbdsdpz4Q+pjT+uY/6MctbpMTqhmGiS7Uu
KFpSkSWpgwTkP0UbGyPZVZRVfOK6pbj+MXFMny1nn3mDSElqyW3/y7ZDxey0dg3+
kd/QBcQjp5WCCHGQ2K2Y1s7yXyDAlQdneMOwKDP78pQAkszGraK0/CuPG0rhcP+N
FVmWtX5ctxQIEVlNv2m0oIsc9wxJLqylria1qnG21WOlweq9P7BM0z1bNDMTMhnJ
qYeVNQxyl88sn+NkIeCCJd0ZhZQ50e8DSkz9W5LMf6pDziPAVHPjdXZYVEiquTlC
+/DSKszC66sZN2wWGFowc/jqG11xRp39fnK516PhRog1Z3M/XRo+U39fxIZMp4+S
vWAWTVLy4rDGqPXGJpoKjRMzI1uOEzmWef7XCH8Xry19BMulY7xTSp7sY8tJM5lz
X2XarWgS2b13+KOxTM7fRHgchLanHBpTil3R0kOkC6Wadq0rLySXXzNw3E3F8zPS
7cPKlw2XMhT/Ak8Q+Ys5uofFz5A2D4xhQNn0Q63BlRUSn8IfKmczAeR8mx6J9hKt
GeE6mVTYoUs3BRtFSG7x+No2zz/sXivPY3AoACHiKWH32Two+fVTKZPGdjGzoBKT
AwCykX8Syf1Ig7SmqUXwAoDYVqMhFVXyboqh4io9MMo4XI7FZP6ur4kjoULfTuY3
1+rQnhDQYpD17F+D5kNSkm73LfzO4V+daQ/ICWjtymblzCNuqoyjOCfq2oUqVTuv
RTbBEjdBsb0RDonc4o3SisbC7Bs/ijgpmes6XGFHQ8F2uec373iOgm89dfTkmrsH
SnEJc+/kfoEV6wkSUJ5AiI5j6xD0K6c0PefykqR9eKrmSYNZnFSuHGRqLbk4zME5
4ofiqx0xv1InkxFX86LYCTzalmYjzUAe9FqFcla2dQSRWUHkYP0VE2ZM3hqATSMA
mkNIULiesbFHoUAG0FJgST5jh5pvLSkJtIfawhp2aqD+1RneLbWgOqyevquVeKPx
AT/9+XtB+b4H2obTTMKboFjsR/sNVPZf+WAqDVWbkRks/hrrZmqJZ9Dse3yl81bh
Ed68MnkM510FkUkV2G5PfjRivyKLTMUO7RtqUvy+FmgUZmZBs77k4j/EPBO/XZBs
FnLx1VY4iYcVjSqRLLx+jJvD9QDee+D6N7JozYPBSvSjltlrPN7a8Y9vWcLRdNjM
foBPqW8kpO+cIwOaQ/JsztowZnfSK2+zEouctFveetka4e9pq1qYS06waXd8pdxf
SlT0giPslXkD2aEI4hK6RANFD9xaW7I2PvZxFHZV0XdAQUucWvTtaRhg6eSZkEzq
0JPUKEozZxMArSe+SpPyWMjhpHSGB4NufNDd7fm/dp31wJxkNUIuI+RVOxUcl2T4
t6cpPN3FmCvDbWB5uOk1t2bkrFGW5RWbeCtr3QHnnekYCRpL3I3Y9a+WS9fsPdJ0
Ib+Ha5L/dxkL/vIIDI57L4hvXaZSOmTAh4AUDcvzQa/taKd2icj1I6j/LxqNQ+cK
MYVZ1csq6wP2X/tdgs/eOXC86UNHz3rzZm6pDCwhQnVBfc+lL1SdyJu9Hrbz8+3l
eqTZZ/i/nuDGAeKKDZO8fbrqJBhEbIc6Av9bS+5NB71jvARTNN3H84Wm1wHJW2s8
9b8bj89cd1YJj3WzZGsYwH2tgO3uo1/58MqYNPPfJmMmRwZutrJJjziW2hGz/qfI
8vXeb9mH4qW1VxIkYtx/suGbq3mnoXCo4J9QW6fQ+6DfEvlHUcWBpa9LRTe+0REG
QCDXFPT0ZI/Y/J96zJCzpNLTqGOzwvAPnlrI3c03T5B4778DYZ3FGFJ+mxWHS0T6
hWGbb+Ik3KPHzDh4GuNWFxpvQVFrfzYoPWz2bFS1DSWpoQHjDgz0CaqYLxr4FjZ+
PntaCjrzABi1YmsPfqTCHb+wsj2sEUyDSjKYpwwTXqjX/vTMpkUo/2OH4EocZpJe
aecou39fUGPbrqTGuUYKqSsYZQs2jNj1y1O8r4pULWowQpNqAyHUAmQ95/OZYZ+9
R2l7k0zsfdAm/ncBkVje957F0FyQsYlij4mMHARsYIUPEkx3T0jvptNPSMKW4Z4n
fid6SB+55NTneinpdO8kA3Bk4h9OPEE9UgwQHkVLnphy0fGFj2axoe6d4102iJvK
Hme+cfdtUl4+yVC6ec7vC0RWnpT8/ePt3fN0YX27dDpZLqe1J0XmtTzfgIbXWtTC
9mOGPSIjZNStO9xQLR6k3uA/R63BEx+FPCudj7Il+kbVgWzsgfLoa1l0jZwD+2B+
p9CI6efHMClfrcstC6rLkfxB/sgviyQT5NmR0UNLtfQeabE8EPhsOp1YfDZi1WcC
1sP4GMS9a0qBwp6BbCvya7bapZruJ0tMIimk+ZxO2zLTZWGZhO1TCupl+sCFoxU6
3SvbxVoArzNh6pBvx/CptSwDBKumdwDErVdis30Tzt4C1LacTTCNwfbvUdj8kvc3
NFoKmSqgH18HrCxaGLR+/c2s8HOS48wthfn6Levlvn2YZEG5omdamQMPqgWvdKxq
wNS/AsnJvwQrrqXE/saIt05npOZo80e05MdX3OFvSITStJP4UK5KhHLqss1sgMef
MJDM8FZyVi3ejsI1yeoYwLWqhEV6jA1iquv2gzj6Svj8h3fVyOALZ+suzR0Gx/tk
tIUlgSBHFR8xtjuVIrtgJiRv5T0Po/K5xuC5MEBwb7CJAlqynlZPjFvQIbD+Pvql
Jr4BBxysF8Cj/Z5HX9oUC7rhc7VB5i8uR7KHhWo7/QIbfmFHfc0/KzFpK5rbO+r0
NcQlfV7p6QxtHcBHCJqrWd1RfaILojIbRWYCX4Kx0oYhnBAwD1Av62amMuXheDd+
5yqVtAUynABRHoov11aq4WF005oAKfUYa3vLd4Q+1XmKJhNN4gRHX8BcpzqoZbzA
KcCPyz6roelzv/Ok0CZTu9IQYPDEmOwn/p8FPpFwEfVEz8v5UFMbwJlswfL9UnAZ
M6hZnYp3wrqWNEw8ybmvkvQO+mpe0AyWashGfDdOG37Jac7sR/ERFKAscfHimPxd
KhyT3JhQ7HWLiHH0b1iq0hOkIRG7chCRgVuNTGqZh3W5toa0/QDry0NlpKXfzcHj
CUui9b0tn5muh5oZkOWlsioqAWT/Ar37PVaLRoQbm+3Mio3cY4BDewJvECROxlma
jOqD0xDp1EiGq9PSFiTy0uzQqwDTq91j66ebHxngjTN/Q6eXnaL1r+6l2aS7wqse
73v3IpzhYL3i6e26QV9PRL0mOvvfnRRRi/Pj5b5kHsD91B/cSANqjdSJd2p3Hw8/
wH3RYJFDT6XYlsIKXVHUQsWEINzdDwyIaHpVtggyqY9rRUFQKgYr5ex4oqt7JSmf
0d4Ins5ZOPcPU2LuINgLbi+kdmhV9Of2T50UMUzu4cOjEnBzeUEjYjYS558gwZkT
FtDYUKyjZYjnlxxmM+m0ZklXkkZvTxmi6HT9evVzYWjV1XKrEzBDRS+tpaHbyK/p
09ib00rm526PDQAd/QGQoGETpu8gmAckjtL/vzOFAeD15jQ5S/ZgOssVVCcDmnxg
FgklVqMW/mePhyWYyuhKLXBdgTf9uPl78Dp1H942BEI5BXxY/5IFQ2E5IKRR7/ID
V3al2tCOwgef6/th/9yl8Oetdn96kK+UoSbFfOfGUfHrqTWYvKFlsnG8UMK0csmW
O55mdSthYEoEGoB2h7YkhyWjn1kkVZHevRciU4BIv8D0TOCmWT1/Tq0gFBF95dFo
kLfq1HPAbbimEed0lCXnzSr5/T56QtJxXKf+Ua/4t2ZaMJ32pHY+WZRjhZDLCCK5
pFJAC34B5RxlKTeYAE/rM05DmeNAUIv5TXhUyoJz0dn2wtmONOX1oeG74VE1HeE8
sKt7or+eZcTrV9WUQ+wQb07apzZf7RDsUYtPHfSFsspecmOvD/Rg0n5RDBjlhRPk
QyyEiM7vnBekqdXD9P7Xo4iNPyoYsOUzahJjgqbL6jgb3gCA0pOt79yVRl9gHA0Y
hMn3MapSf1SldkTOraVfTpQ40dvQtAuNXJUTCmbTNekcnAGKKfUmNAmxIor07PxD
qRsVCXKbgplm1DWgsQjFPEhpxBw6WwNRgAyH6M1ex4TX2A/Xrkd4arQNIWkDhalw
UM+kQGRjILO4ogpb1s8v4M1y4tXJ39x0Gg6C3Ra7IQ7o8W2ZjJVFweKmMLnNjqcz
T2m5IJ7AIF2Iy9VYOtfXKFTUoYx3dKd0N59QkUrz+4TqO2dmFRGJMn1FObMPBcSq
e5h483jvHU7GDIuJUg46uqY42YomUv8VbP9J6oCTxkQoryxoybSReqLjRIZBY8lU
WdkuwcMkic83M1ifK4uL6fFj7dRi0LY70KBAlKUsFAkFkU5b0qO18HYBUnviUWg+
BHR7z1OyHRcyQyA2Ol+FpvGIp0aW1JWqNaX2AszhNmbfAwTyrGNmpdqhHDcSOFbG
K3E8+76p38zcH78m7QmZSSVx1g2Oj4VpAHRxvDTp44/KBVTzsk8XRQsJL9t/5PFd
LzXCU00Md4K2+fB2Ud7TrFABpOq/1OyLDmKo2ulpqLR5y8MEZ+BgUZQqWqzUqtcS
ds7y0hqoXacG9bfnuV8J13k2K3Er0jC24oe4lnHJtMMS6Yb8qNb//+2HCnvyM7yO
v1yWIqne8cGUTNBEvabVZMImtGylJPlzONAR3c63y2xpmzSPjJk2ujrHAzK0VnL3
C0ztNIN0ll16ltkouhZUp+PT16P9CYXmLOFh8ziViPaG3uo8vcESoEd7n9UNQccy
O7xg6EYAM0wGOZ8zrMIh7fBmMkxUd013dfFFlGNoH5+loTm3rCjuwAp0yNYi3IoI
cyGIwAFFJC4faP1dL59yvgRFgaen+tswrdGa7Jksq1XAL+htEn/iVGK43KHOs1oe
oQ3GTl4waNy1sik6qaY3lTSqUJZRx2G/ZHPk0s7O4V7wvriIy2QSt9jp8q3VEkqM
m4md+jr8pdL59qHHvnz3vEc55sgxbVegyrNZBjRr1nbQQglS0b2irUa5HzgDQ5KO
J5ZngBOF8kIw1SJNMCeIolcrP1T0Z+gNiOcY/G5OlclvEEskBj2uycN2M14eKhWl
LD6ZxAH+9n2QCGL82FQfYtrHmXHtmQI/Us9fbliZ2P0GHPr6OCExcHMcnLYaD0ZN
eF3hiSYNFOJqfBfA+RgEnUwXagL0ktU/jK6zmaar1R43j3OHD+nrM4xGc0GTVYr2
D3c6flGLy0puy78ddYm8nQl9YB2617Q8cZQ6wfWxPz9dinpb6Ib+yfOkF1gY2rBA
1yXBwqF19wr45bXFVWneu9nCqQsB7cYVJthLP0sblcedB/GYq7QTuwsQv+0u+f5Z
tQZwoA2WKURK28AH8fzwcGkqmQTRBr3ix0CM/Fdxxrw7Y6Tw84hg0wdQtxKPB0Wm
KNRvNn0ZmlyjNikzIb30/rQsBXnJX/NzAvItU+2tgE2fkdE8HLnEMfxWTJjbXQlc
RFD8jgFbieafK9AZ6Wuyg72n/POulf84DgDAhk2Py4oOF38ByAWsf7R3lQbjdg2S
TQuhrPqwxEsGr6DLiYU7q4vR1DrqY69n2/eIULs50qgy7APBLax+t9ZfKoe+Cr3D
61Jpe7YvJYQVmpWozhRKCmigrhH1DEUlK+swLqHpff5tBEyEnLwf88Fnx1myhXVg
qElQYzf1d/+9BSiOyh5xn7+YB9qMgILDv9HLrtOq7EQ5UHSliuzVKfC+wu28Zg4e
2UTxfnvr4yYANEejTpiBoLEJ7h/Kmtsh+kecCIId4eW1TPxHKZkm9PxMacW4wFiq
TG7C0asJv1xD0dfF5qbh0tgYHYgOc8MSedbMRx2QMzIt4rO/GT2mmLYtncxvUV8B
imxwwxVZM9EeqkyvdcDbOPXiuekpbztTcL95ZlYIYdRegm1uF25zmoowBqBM+FSh
Oic+yo5UwIvmE6MZeNwRJJ3Pfw0z0UDtljDVlZUoD31JxbyroTQ6fCrmY/K0h3Om
VOA6lE9q1Z3pjAO+XV2NACVWeMSNPlWxG67ogRRlZ+dk9ePnPrzJJ/Ruo+ueWUKO
FMF4iB4EuAwe1lCSFvy95YR68EshDNDGtigcjJafT/vZzQ/XpcSh0ze5klFUiIPH
sOSVA+NmG48J9Kh1umWjQmNfex/+05ym80NHO8zGsvy12/FsViku3jgATCrFC1W0
IbP3wz9UTgvMc/Z/HvGaYzjabtOHwIlKlM5hSRItZI+IP+LZnReYqHl5+LKzLgPR
9ZU+fXbf+RY/JS7f7GMYVVh1RVCQMDDRAbCh+9ZSN+Y+EcwNZ8Ma1q8zqNYDIEHg
A6yzux48T5C9JDUmmMGPXJaXuToyrFkVEDZ7FgAJB5pt6jW05AICHey1OacwDKwp
pGe3puZVwT8M64sh4Ug12P2rP/wL2Ax1b5oRvLKjsWrQuLgqJcw94UTgaCVQ79Cl
TaJ2t9Sx6u57UOiujv1mxuAOSxA0bC9MgBE8AYmtzPo5fpXRNSAm7lr9PQfhtpoo
eI7dB8eSMpyokNiFiAaEbVk1GW8H95M9hmdNdUy/xIt0YbTFtyFMtCnoQPpbCzTj
3kgQGIXI8OeHsA5aXWxBoDvHqx3jju6H8CAxr1tDRFYgtvuTQ5428S7M0EZmXEwM
MznB5yUDXwBN/VCBz9cnAt5huFIYhKbhCDDoSUPmglIVT+peXMcHwi2GU6eRLZOa
xePLzurMQuxdXcopgDRx6lgNtGfMcMyK74Qn3/Ql6cXNFkjD59Y8CAHvmGOVaUfJ
dXIlNK0QktILiOkM99LdTyfRrfyNZ6IARYPfdb7OgWgvHmN432k7q477W9OpQSqi
tDSTnwlAKU7GJmT2uscl/j0u3GsugWHb8lkqaqk8egOX04Us1PVXtGfZXZNE47Vf
YTD9HBLREO3fVDRSVP+TnWmpvlUOksDpwyb3LjiovUKPKE3OnaeDT0U9NrhXcS9i
91jp8ZBJO9QBGy2n7+bZzJqCPK3Dk8cSW4cDilEZHG6rK1tHWqKoITK2aDvYMiEa
+rDo4Tv8ITgx0s8b7/DNrov+WaYhrmO4mWLiAHPY7KLgcKoKmLQxMakhs9DftB5K
0u/rRu1RvPRETxfKHOgcdBXnsRZKUa4sPR25MEv7ZgOObcFBPqCk/ZvTvX/gtxyx
MX8jafo3ttz1wmnOGGIHViRHu5OYRyP2/zznWh4MjoImqkail5oZjsswjrAI9bLw
BtG+AhhP6BKBNgyrv1nStBn8/WuKXt4HUiLqO+SNdSJxu3GCdMlwihgFNFlqTBpk
KPIddzqudKu+PzDvJEKXmt2sSx1o/QtJxOd+ZBqo2R6VKVPC39UCqN3P6f2oIDqu
p/iWnDFztKMAOLuHFdAlJg8ppwbPv8pwlQGYYaaB5+36gY3JWdS4pel0+F8lKkY0
WcvjuMf36SOLSqCLW5nnY3gOtgJ6o4lqcxk088mUSsEHajF7CP0Wy3fpBQWav/M7
7RLU0yzkZ9rDXGrUbwZXkQSJxghpjkWF00e7RXRSoXV1A2NWJ5TcE8q55obwRXnK
LQYdTyKY89qJx3fx2uIk2kb2NMsIGzMckTAaTseNBEUC6wXKIaXL86hMKxlZk7DF
YrTurfDXsqzdPGiBW48+BnuEsBByGJsnZprgyRE4aqlproDJIESPXu9f91w0zJ64
j72PPM1vJwbIzz1ldBXfHqg9YJp1mdjCh7Hd15vvmvqtwzdcKqZQNADF75YUbaOB
kyZ7eOqtryTPzknkFWeuSTwzTCHzzsJ1rsVgIqIdwY77RewtiDWDfYS3gtUZ2rhK
tIqgyOX5ejwwpC2jkUDensNKJ1C2h2KUKAevxydprR7oBz3KqYHMA9FtI1dXpRdE
0thiVscijhh9TfQ2GLognWnDdKSEnO/Tv0hpr+hwRWGCIvi6XZ8oGOiOCtL4uxVG
bGJSb0R06ZPuvIezmf/dnwOn895Q7AaPPgZTuGFif9EL4yax/EGFi81+mYxTW+zZ
iNQLGY08MG+Vgj123odfCvNusBVw9WBWlj5uS+qetU0w4DiM31qO43Je7QmsWlHo
nb/Ij+7javkkvcN1QxLdtFYvnUTgGuMMf1stAmKHCHt4OySSBHdRaoXybzhJpPoq
T0sdR5sZ2mdsz23BBUF3RaNreDUdDZT2aO+QpASuT9YUJCt8WaVb7LHvH3HyRXE0
CYHbWJ1FypXPdW8NoNjqSmPL42Giq+VlTXgHJ67CrEd9sfoN+qBAUHxrjkmC1ZKm
eXKC1SNPNWeTyvvCEhqxY9QPkYMDkQSXr6Es2waPQMCxXfBhKTgjHoQIErDDptIJ
zrojN+3WmbwtkfIp9dKLHZVVSJ3eFKEbnc8f8kfWPFc9sh82GHmtarxINoKyZT9d
eG+yzG05lWeAU90JLhVSX0cV/l01EkkC6izvAMTHb45lbAwmqWGIR7+5SkngIBjo
UeXzgL/K4iI9dk3WYvFjRweHW22Vj02WVx9Eln/T1Ys81zr2BSoukgbUX1VswdIt
TC7AAcn9qVx0r+UyReY5QeGuNfdrBWzAqvOEqBmOvNhqpKGtZSWicHDlHDHIlmVA
8dC8KFwPUgk3NHE3RK+3RiAHfYqHs/1t/tJfyxJQYxplk+wtfe5n5dcJDeNa29MH
8UJEsdAsN7mss3sO5SedMLy+rSOkxChLlQq5JxVcUWOWInZA6CpnPQBYvwNrJvWT
zC6t+uAyKHvcrpjV4YwmAoDQTI+qboPlRzj4BerxekBbHlMg9bpp9K/NCjez6wLq
h5TfUtXDHM4iyUvc4MYHXWeoXd9iEJ5YgoM4WV12RhGj6+UPXLO1k2e5VSFRl8Xn
Qk32lhmQffqdm0NKvYY6ek3BFj/sxiYRONyONrJkmbnZXjzvdBEBN6zXumHXAhKZ
JBct39bQCxiGuCWzSi2WJfHKlg1oTuhTBfYHNzXSFfi0n7S5QyrzAqOt62DENDVL
MuLJk764GKJfR8ZkBWtCzR0eT95tj1Z8PqKPvypIfurupW6hzqpAFr/iADe95JqB
xMagVkOoBmghNMjjRn5m9MsohSNOgfnCuvspKv4KROnkXf241ji6/lqpoAOaPdrq
353QbYf81y2eD/JvVhlwD00zapGpBT7RSxDQZLpt2M0GeLrq46LRg8QXYq44RzdK
8SJQT+8ahQF4sK7lo+UG9Nkrv1FbzH/k0lz0y9skeG95Akzl3cnvQAkY96NTDPkv
ZrgeL3RqiAtxowXj9jNJ0gO3SMMBP6b/ZjpPjGex1tZ4JtrlrFHpQZGUo7ygh5si
pFim2SKHL2I3CR4YvcJlU82ZfhzEJ7rcYbjocQT2w3cmcr82rxR83zepu+44CvzF
tFtbQS1ALAJyazQnmFsmUwpFzyyxBchEIwDHsA+7HRCXvR5MFehotPZtABEnCD6M
pZlq107Bd69KyrTbsmj1dPdcQNJrxwwAgJnDCcAgHJP+FSMGbACkRehhqH6donCa
EMSUml0EawFRVr8Xna/jxZFw7F92xR8h09+Yi/EjckzI4qHcMBjtpHTKjH4fQEnh
RMxDEFwwiakGctel/t6WrBiTjqTVHf4Z2AX8eQH+3GJmT8NzJixvEDiKL5v//65U
JznzJPvXIeN+UIVqRX8mjkuELT2Dp9vZhWdB6ACr0pSYK0a60accOCuXWx84Hy9f
VWCYU/fwMQ6Ox7WifjXkIEi+M1dZxJVRYO4IaDjORBQYxYtHbvsSzqNBuSk4vaSo
3UCb3wzpV4w96QX737zfu1G0GLD9ur/B+IgglWwsENSljlMMv8zWcSxY05Se7btk
aI5khFrtN5DDe48+Be+qgWmF4yoePmOj7nsKyytD6m4Xw5+5NYDIAtnNtccUBSpE
IdTdL+aLWzTLSUenO9Z0kdus3ZghuUVy+clbU4DJQ8apMY1U3If1640366cfFj5q
9z+rKxRdEs/maY8xbMIbc5FaB6Y/fTxQ1D/LkRTdQpJUmmrgagOdxqot4sA9QZSz
kX4wKYdtgSVHnSuLWDgbZPT8mQXL5tFmbqCHcK7v6AokB7SgZjkV99As1wuiTUhJ
JGHD0sMBuMWxhCSoXsaOmeOb8wFzvdFHU9N9kDQc9PLf1tB7+S3Bwn+U0zG2V7lA
ucezuv4iwSwuOhcnKStOYox3YdcqgXgoU9ze6PRrzphAyb3Y8YUWdX/K4Y5xCqfd
CJZz2sbgxcRCCrqa3fBcWVXBcaVW9SP11SLUPUeNPyTWUFv4thv7NmTlV5y4PteI
zJXHrQzfkfYazK8CS59LvgY7bcRAr4zMV2m80fhmeamkQCb1wemI6qyEGD6C0c3f
PJtxzq+4l7kRSIx495eyrRDAzGeNVTZRSc6F5F6cJEFqsTW0OOEa4LuNUn2sd7Kn
fsNCfpJqXSX57ewO5dUFDC4LHpH1QKyIv2GQqeaLpGDQ2KnZGGuXi3hPhoSGb9lh
bsV5CYlOStFgIws03EAN6zSvr0JMsDcsS/tmYfFH10QJFh3YNwPaH9IYFlJPqp6c
TBeJo7wWCd4PLzQKij4w1AmvNHLiWH8PjcSBvzh+meR8vevH1gwEfOTDovd9GQJ+
ETUDxb7pupZcGZCnXba8croyAhlsx5Vj07fNhYD8MkVnnRYUs0PoFt9jrQh1aYNn
hSd/aACbGam4Qj4Rp4TOb1ntqEMLrjjo/d3bjwWjpwk1/4WgOqNIxcFFLnHaf3ID
JrVO8mQn5B42mHOVnHrqR2zcSwGLSF6VySQi4fdz+6HS+kYwU2+CyidjutIDTS5F
0CnB7Lj31qMufv9cZqXfjge4ESX46DtFVmjnilPoSI5sKQjJTZOkTE6Z6pCXtFO0
46D5+2wo146CURRjhHtqLTQnMo1AJ0heacwAlO2bQO6eL+EiOhosU0iu+A/3NIDB
Idh73yaJbispgd158915QX2ntG9Gyarseynq6sJznnel64gWngQfNWv6kaG6e3Mp
oiSTi1/FZA3tGzOImm9nF9zh7qsY58f/dnj/tOQENA2q2mV4OaQYjDQ++8LOSHeM
FsPGwOO8mGFjMCxwRIELNFuVLImY8ZpQdOZVvehSXXTubV+dDXIa2I3SGKEEkeRF
+WquRx2kGqS1FZlwKMNsQ+i/AogpSP5iOGMyPhaW7sf0JKhnu/b3cZIW4+ehLiE6
fnRLheb37hTnSJugv85aq2Caxrqa6Qk+n2B6NVyD+HFRMf23CABR9gNHcNnoEaSQ
v+BvdW327Sw9v87NUjiPXmDFIVhDKYOKdminJRKaePZmGDd0zUpj55SWCUkUhD+V
xhwlpBhDLwwXvzbXwTGpVydDW5/cExFzmZaGfsonxtjpimFHNadR/+sQxlfib4XD
bVODfBA12/3zS/pfeyrANZI3MZ1reX6+kGZj0CdPZJYYZCC2WhAVergdh+BqoUmq
2JUJGsDhRZAhTkZ+4ihDPO/vMSIgPomed4gB/j2eFKatRTi/ylprzRIo5RPY7s+Z
ykIg2DhX2C0u/wOLO3eX1siiF/U/n339Jm2E9Tb4IxqkmPCMSkbVRfT42dyARNrl
I9KH9WV8hBONnoWndhsqCb0tWv2AMDSZO2Y6SSqLn7wFEKPHCNljKv+SPQSWJE2q
576JYzL8LRPnk+FzEq6xPJ0kQ9wSBCbteur8kx/b2zc8ZH/9xrjO5v5wy/f8eJcE
ErGQX6SPIewYyg5FxRJh9rxqAWZD2uPL9UgPzrPfIboa0N5o7QVQt0OhnS0clk3T
X5iabBEt0peHNPvvkjs68WXtr3bxq9k46gkUmb0c6q17Ll4sJQ8A2q3f7MXmek2p
tMtkJXJWqcvMSOhToNRr35TW+jssdSHtCc5bcTgCrE2dBHEjqaLnqe1BkgNq/8FZ
RXnG20mrILjWELKhuxeBsQBjQM2v0aIfmhWP1bdb2mA7vzZGh3hAsR+mTM1Kmncr
Kws9BDjltPuKM/sp+NWKxhvc4gySHU+DAtmgtBmgRE75N6Ume3XkNbgbxRJszQIv
hpEpl4u1gOZfIBTrWe58MdbYs6tHls6MB9BLn6X5CKd5wl0pRFbuCD/f+fAzltfM
URwLiJPoGiPhn4F8wlgwfUBPbkabw2QdejKtLH4oXsF6EQBInB8OsQJdmcj04BFT
m5t8FxCug3/UOCqnruEXhuhvfSf2HVh+1Jt85b4VrEWDiPPKIcSqw+otkC7IR4iE
Lx64l20nPdC3ZjU6hWlgd5n4v8jtG7la2gO9a4tEPWMojgO71nzz1gd4pQYTWHh2
3Nr7DZVmieXWPCITjkfhdP06DR9UPSx8CQRTZzYzoKps/YIkf9c9EOqTq7AGgzkQ
2EBlK6sJU7kwLsMQfXwP/MjzivG9cqee2e/ha8T2rEJGcG0AE10vuc8188iEiCMq
BZ9EXvkw/fO8JjHUvwKCSahvx7vwocJ2m9VBDGak5A+ykO2Bsa5f0hXyLjSzvcrb
dN/VTtm1VxiEwc+BpNWSda6MOCKAWtLvKCEhwfRS/ee77blqNfICPkF8PJ7DJADw
uiWHWl6NrD+6wc+sgc/osHklvb0uv/ENJeJajQyipAgD7z/T1Z4jhWrtaSXnDZGZ
XYMHif4Q6M/UBqBepfBtyA6TSWiiT6k3sGU3so0AL9Vso3Z9BAPETIwe4umyBIj0
v1BN47p1Y4T7rMhQNSGPxhVNEDz2L2g+5R9BWcMDsR0fKTu9KomrBNKlkGgwf784
AN4Yj08dEUaTk0LmGJmNcjATz/jwfwSKodRu8uy2L59sf4B9HVgHGe7arjUZFOqs
3scl5pcx4vBnEV4V+N5dqxaOFuGWdS4YwcbtWsut+i+nhmA6xR83rvZZrfIVD5DN
v8an+S9c7mwexbxbeNuWSePRqEAoeR/WFn4o071RYEbcosKLZ+6VWZ3XoiIyKm0z
slRWQuaxs4oHYX7WlDk99tHEUkR+b//1F+RYL3ES2FQBZUgKYN0bOGEHdiliDbpW
d/lpKGNiJnfaaZ5QDma799GQDnJwawGJNl4avyhOE/OFyYrV6gQAQ5xFdvxXIqTb
DEDqheai46tZ9LD7T3heL24q1ohqUchbRepBS/tmHGa0Nzc4CRfxVdfMCPJhzF9A
j+MdGhBEIXnXYk9dYAXZFlPvpuurPHo+FMjbLnIhbxEgQ4cBO+b59Hb/DkRuVi99
r8m8ycypVza4MYbF1okgF8sHqkAYa6u6Vu6XCq5TgmRntaltX+BLwgmSW8B1cwNN
Pde0+uJmDPQ9zrplYjbAaftGuwFyaJUBSIS77l0QjYCtIetTL62y4T9X7VZHYce/
wsRfCGknCBLoU4eSe2KrPZK3k49JYPml2IYl9/SBhytQXX/E6LVjBaKnWUVj6lJ+
VmoNPOayyn2HpgLAEtmPhCR5fHwxTexVcdtnObVTqOvr26OIe3C+zjNv4nwnKqQW
9dzkIem0zEWDdmarbh0puT8X07Ok9tnbDsFy4agIuX6Xmh/Ziy8NZXPucvl2Cpqa
kpDRZxHZxT6EX69P5JmDrCIvW9miIAhVKqqO3ac+UW4tpwU6IXJahuYlqB59drW2
SCyEePiQWXMOf2pdMK4UQF37LCBQY7PMJx5bSVRHhO6J4ePwYfMcfIWyUvM2mlj8
21s3w8q6brx2syVY0pQiL05fab3L3+vNS0GGTKmHtYpyk0pnjbWmuQpC+rdLwXEU
R/JfWfXuG/NPku+Jmka6t4bwi1ut6+5tx+6a5tdDo8wuwRGnCFDkD79GPJCNPZoo
dDjQ92wpNhklpFZVUqHhX7sdQf5dvw7TuLnVJVhlzPKIHbDeXwnmcytiszsNxUZ8
GPslN4VW3jcCeWQKciFAO1nklnL0WbD62ivil54Q2st4cqEEhv0rf0wqsutlnXMf
hnoEaLCNwBx83O2BuS5bOcN1AqETNk+cCo4QS9qvcNy8KyDMhoXfBOfRy+L0o25b
3gYAK/0gwxNBUxUOfO+TN8RNaPl3WJ/9Ak0w5ecmju9+XQ+h5e8ea4xMWNK7C8Rr
tBpx8yIcOpO6WSVx/klbkXWaZ5sDqdzFH0VDKJXdnurW2GC5lydjBUbv26Wezfg0
0wBXEN41E56rhh04iOMa1hYFFhHroiUoW7mFskdSBoZNNOnVuSVemJH1+4NknEM+
MiNtFhAsuDO20FyjfrLqeNKkcAtzFpUeyuhSRWFRVDKSUb4TwwEptgkjF7GCN+1i
CpljoDkKKgqjmoaHeUxuu2CtMHYcY4f5ecBTtBbEkVsadpaapHcQFbn9yLIztq6U
IZZzVAXRKXIbN6mYieIljTrN+jPAAwFHl7A9x+YO2XI9ftBg2OFCSIUp85QVk8a+
dKaK7UWYhxl/gdjyZn9aLBOQ2VTLinvLdrOIlh9jvP/klzfbsOj6OX7RS2cqhozz
4AyDCCHVciCoTdGJj59242tPs6oCZsVo2mFmlSrxG6gIfNqt+U0u/QdGEU2dS8H0
UvdL4kp3dowMdRknTlCNAq9BSIjJRyTfFAl4aoktxoPQYpittGGeM9FkCjdkIA9F
D3vNti6hdn7kQLa3IJMexhKHLH5XCWZLJFZfaGY6F36yHY6DcYqHtEs4ECKwNyJw
nBaN1z7jlBqfH3cQl7noTw1uF/9451FYalFermUwRXhUtQnLgRKaih3zfDDyn9Pa
KKQoYDn6U8j1yqlPXcRm0Oa3bpKBzjUo/0kPEd3DmxJlIyoJRVaQbxQHLVFhFMTj
FBLhFlK8a2msXIz2KedG4mXVFlXSqkUQyPvDa4jiWEN3zavLVUvZ/QzxB75PRUX+
KUENoVtipSuOHT20HIHcJV2tvSXmmARFNjpaDabQEAdBUfC+U3vWUeaQzYWH2k2K
cDDvPV4r6JWoLSoszOxz5xzIH4JdHgWNaSIoSNptDtbFW1heOVWdfQSwNgAapGco
KAi46IrIMciedco2I0X2oyvTvpNCTjclnD8puKu/EEFD2F/MhpeOXxn/6SGFVnvk
p1m5PvvbR6Ll52ss9h9k9qCel9HL11DSJnPv5Csjzenq1IvsJplSSrIcjAzO3U/L
FuIIXSvR6328x6XbWSHRalkKiTDF09GzCtZVxMM1mBAwwPrXrOOzy0bszRL2MttO
/Sw6tOgR2d3ZB8/LSdlC+W9RRzkQua4hQzmufTGaESjAqvDKt+kS0kSAwQ3aZfdN
tavn+2ihaAQ9X+VGPV2XmsHlK4myHnqUAva3leRLsNyE62TL5W9o+wWhLtVtYAlT
GvG4g40yvJhHz0aUPsb2IYc16SfFeTMWkTiQ8rqeqceDuqBp3ImYFyLEhvLv0LAZ
erNf8BYfABBsVr2tlzPEDF8QneXmb85Be4dHyZAv75/SPOe2bhb60MqFIUxIrGHQ
F6isGjEDXsGXhNhOwNcFvbpawZTs4HGkIGl6GXMif0bgOIFrRD5rLLlp2pRlbmci
RHlhnBxoK2W8GjBDK/14tVIyaz8uz/tSVNM1NASnS473z8WxqwGB1mvntiIq7cQ4
CdV5Jq+omzvxyZJgE/jTfXoI2LQwLmiviDTGaDgbydYmrtG9ycdT9ElMfnqwWBbL
WJ7hggdyMpCSQ83x1aEEfBzs8CZ6OFLyMBUd6NqkltR9wQLryLo9jUyZekwkfGLC
tuC9IKOs/DToTB4ves5kj2uYpAaGX5Bu4Ljn/E3RCwmip7jT8lD0ozpWvO4QvgaU
zQc3adr4pfqNxcURVeu8AsVdys9xNSsFUc9Lb09oHlKYjRoNsSfrBhFcPRtSGjUK
rV8Ul4GK698aiP/OgFJhwqyDVElRZdPaa+jkwx0Fo26KiwJ3P0MQU0QeKlc/MlL0
a1BKR8TVpYRUWP4FTBVkwW+HyS1euoyW34RtZ/9sB6nRGbTKgzdayyywNpnMs5JK
/cetJsyUW45N9p9f841R/LC29J9Q2Rn897P+jQ4sOJlGSSrZnNkfxDjV/EPhEBZ8
2hxux2zHsmGnrv7Pajkq3BFnv+qN3Vjnlb332/hzDRD/7xUqd+uaJ7ufKziLg+8h
yxuVRkO0XBjEwYv0sRQexx7uFhL2xTuRRgXv/zuK/qO3RZ1QM6r3z8+fjbu09Vni
RS1ywEo7nRh21tAr7+gdWKxzAjERNpvTioTSC4NtbQLQor7XzzBuTiwoLrn9tLIz
qg9ZWbyUYm+z1xz/yxgJw6MpSLApEPGRDEJ7Z8KIYBOPuEg7Cppq1TvsGv52R4yi
LtSE1uSV/16TJGfQqWRNCuQEOwNFXZq5/V+2JSpkRSPgm9EQJfAEbyL5hPVzpO2M
jWi6VYZo1RYKdSMEOpNLHO2kNkoLopjKgMNfUbxutUAs17DZmRZm34x9HTcIrais
yJ9tffrOaZfnfWMtYvLuX1uxFwzHuOF5eGiuo8sAu465WhD2sHc7lQIDWRDWJZS6
iUWxojOIDDXjVLVNrIo+rjEGl8ZplE9cqTQ8u9qV2C3ukx6AqqDL1/Nh+7nErAU+
F3md5l5STu9PWj5vSYg984jh+6LhAbqkAtHE/DBtkpTR5VwBZwwJmI61DjBLV+3t
/diVPdcEY5F+jxEP2frkxik/Oqj6IJsrJjOX+nPjAXAQlpW1uDgFOBNqBz21fzf6
AtjFidQ+HbyKEaV7Xex5AH0hSnfnTFPm+vOrufd5cr8c1BBXaXnMEeAD5MU/288K
T1nZ5UpuzdOslJZzWhvqFLR663mklZTOx0Of85dEExmvV76qipoLUxTSLc9zfPMb
SgT7w4Vi6laaiDzQ0F/kC6lp+yoW3w9F61HjGUeDDLmcM0uPEP7Qn+g3PeO5wJLG
M0/yqz8nydDotH5n3qm25nPi0NZw/vUODP1IN1FJKHrCVxSYGALgbjvrVF/2oV6V
Iwl90Jr40ko0qfaBapf/JxV0pDhg9lh/j7zgj5XUSTM6kJMrdpYYXxP3xP6ZicX6
XWbJwQha1QgBsa+89MHm7cwbGHGx/D3A2xL2j73rbzLMXUdo+HTJ8gc77FkscTC5
puB8in944hDFn/3AZ8mQCgABSvbXmLOUVv/YyAK9LLK+BLJYT77as447n+XAdCgJ
UnBM6bOe6yGlxNA+p//X910sdh7RGBOWYHsSnmyJYbfshDFKLtYPyaCBwvfHOG5x
Xj27sSIfH1oFF1BMW8vXDbLpZJeLCyvv8R+eeYGh0chzTFHCfp4OSWdNzgqmrUQ5
bI1jbqlfxCX7DmlwW+YPvar1qzMfJhUAG1Yzn60wAcpPQpEobgsGEGl/QgPz8kdh
B6LQ6RwLAFKcWRM5DrdHNJV7/kwLRgvfPsIbfnQPfty+1iHdZbua9eKLD1SWsC1F
TL0J6g46RNQVblXkZACiujkLqK0i/D8r8ZjLdQhRatVb+E8GeePd8lE+7/KrvxV1
WYSpZrQlVhNXL8aFkNFAD9jAsl7HWIjZ5vgx6WDMzgaIr5mdSdsvOaDf3a+CAyy/
E66zYeYfDhWzTLD3hH9YeAcsoJxggoH7payRwukSYNyl5opTq+jrXJNvif3/U+Ou
GKin79VkEVxGAeFHx4lMwLnsoD/UudeElazlFh211sbikWuUetS5erEsA34iMOFf
pHVYW7PKtAZnJmz8hkRiTT9xzmDtPE9bcl5NCkxqjtfoHdhlCQ6jHPJjX1ihgNiN
trRBU545wsQTQXQb4QwgxZqGS3kqMdkdj6thRpINYZqz5KU/Nw9CVdwKgdLx9/98
BYY8yE+PoZQiDYL6R5mALrF9SAqcv0ezskMfYYBexdO9Ztqmh3v7T9yv50U3kKG9
pUNAvp0wlX+h/kpCGx/Lggg0/OWYRxPar6jYPvcnRuqHVp6zCQyiQjFiZLsyfqBb
OWMKgYpD5BdUmZ+1Xhw5WcWOpFKr6s00TCBOxZUTSfB+69zzLyF9laOWrLG8fI5u
rGKr9lUTWLZ5wcksJezW8qPwVmHud3KcvqhzCm4AkATOQYMTzZjI+sJv1mIhNWmO
vrGtLC35cpwnd4gN62WN9fYOju19rjrrH33LQ0yPFptV5OznyN+EnxcVeB+C1d6k
TAaOP6XoBxOBqj76AS9glD0m4abojB5VNJjgWcS7oJ/gLqhrQRkU0V/HQ9V3wSfO
N0Yt+yImgF1SpEGZF3YmpO8/NxSbAd8hVJJep74psjzD1hw9u9PaxzMVYWPjdBmx
OHWcstFVCUkeusQtra3l9HvLZwoOSwz66kwkIofkJ3Z8vuHmgivzqB0etT7ebFtC
DG+/9dSEwxEMwUPCNRVMC+IpmiXvfqFm9OyGGtk1cJKjFpwdHHS7Dv6afl/1sov9
U4XA0Tjzgx3fT43GjGekAN39d9Zx/KJbAP9Jsk+NuIP2H/83Kfwnkms3fXMKdMjZ
KIggFz7qsSrky04+A9UgkWEQFS8JkuT/tn34Oz+ks+s33ab/Uk41ekGHmxpotGGz
VMQl0zWkQss9nvMK65R/BMbWyzl0uOKOpoeDj+BTbQ0lDg8ry6xxiKqOXCFJRrfP
HFbaF5/kk5QSgw24fNTo8leQe/AS3NpbEPTLO0B6yx+NtWKW2VoYEu2TDzpm5ra3
s2uLQ4irQlpQqnrW1SP1bu7x4fVlH7uAIjUgGL5h5+N5n7mhGjB44O6eZo4/FGH7
tIpdkPzenSKGJ+99N2MRgbkjo8SAbI2u4JPRIWiLWM4bCY0sd1zmCBQ0IqidqrEm
CLnMUFum+WJ4FvJxv2S1FE/a/YtgqwYQd3o3Ok3ysEupp5RnNluwJgZoyhQV+odq
faJRPlaMPEcfsYj+8x0jhp62YjzrQuvo6tKoaCvEUItKLForRMhUVcB2CVdSrr8t
cmKWfvRLRckGwsuJf8HyNVo99c3TYibE5cOeT6MzrmpifYqNpXUj7ajDptYjCb3/
XOYyFgRrXXf6GWE29qp3Q5MKfRhRwYmi/OUv8Id2onMZ10cCNYyipdSfwkPwPgrf
PIWs2jpbRcpl8Q9kPScpQ1IYwyiuAGBJqlN4uzzvt+1XA5AyfxAmp/VxwIdYrXE6
nwucLGkwETG/BgROgjgG+PMGHSs01VqgIoAJUhrWIAwjKCMckKiVHywvFHAy+q+j
Nfojp+/hdcjg1poW58p8GbIAeGyWXAzsSWrokW9009022MWVPFk3OQ2lAl/Pn14K
2FPcSOOEp2ZeLgX2mg1NE6zrAFIySwLCJyjA3pY2henAYEX2XQ01GfboRoKq45U/
PGu8EZBY8svo6QyS+tkhbBtUbAoroRSD2fmXoyefpvXr9Q50S+tbydNv16dm+LJK
bNqLnluh+TkJVlaqH7CoBDjI/e6i0UGoJAw/ez4EulNcDN649NwM/Qw4Ix5he3vA
nXQMa2YlJV9ikUJ7y195tqBYwA9XVXBOEjjhfuN2sIv+B0YCGbccomLBy4Il84Ho
OYn92HAALM3DWhAArBAsYvdK8aWJiE4ma+fI7xhIb1pOqs2f5PaFTPJjcTYakV90
eGePhjl6mY7e84qOyTUc/pdon4bOfrUi453+YLIyvsDrYgFYbx9dXED2jTpBxr98
wV5en6JcrDycC8ThnwETNt0d3Gmi3ym8HnfRBaIZ7d/Q/bsEzEBbM55n+1jDsN49
CrhZA+7+0Uuj3NmvU+i4rgypECt2PzFp+HaCfRUFqBG2NZFqNFi+j83jIpFhf+dp
k6IywH8cFSvMG8mEftILMGciGsGkq+7mJY41SGhJZnfqYfgDdGSl+ud2bWNI4Wvr
WCZ5+FPsyr0viBjRz4R4CH9rntj8yf9LHo3oWIfB9aI60uIlpgaz0ugRmRTp1hDE
X7cM1k8sg+xAkxs1PZhOzJuPG+uwmqHfvPgTv44Xu+tu2GhdLzHVfQz4oiNBZMh7
mDmOgx3kFOzmhHxJc1/QA9NzECdvhG5R4Vuy8ixrbqnh4L9zE94JkhIvefWW1dOE
AARFwBe9yv3+Dpg9V4f4hnQgNPbe+j81TmnBpkHRpTJx8xV6DwTdtSMLOWoOnCuB
1/cBVoMbPeKeom/YmyG9wWWVlvvFN3SOZJolmJYkaYzvpaBb7z5neLSfwEBzsuWo
Z184yHIg1eoOYKNvPo01kuTLn+GPutE4rFZS5tst+eTC54r3ph1djPVMMV11AuQJ
P+Kv7U38hSDeQykwKOQ5rTDt4vL0NbJoIPIXPQYPpj7E3glCQhvbpSkplGOfiKPs
9coazBpK66aPCeJX4HV6CjTsxXgiGUZVXvhnqIyzE5T2k+UFctKRe/TlVxq5q8g5
RQdVRY6xiSH5FNyrdc63fbTfYp15EAYz2wRGSBUYwgPNvJ4cXvpN3xIW4mC5dh0W
1Yxy77IwnqJAJKTn/7Phs9s4hoVLmkpYJjoA/RnmMxHXvlyYRamLPkWxKIVFvBg1
COp75GEPXJvCF+hB2VSGfCjgWh66yfNEVF35Om6sP9CgS6X3VOYhhyZdslJJEutW
NBvKRtcNtRRcPNzaFkuakbTHQmXCQ+6klGnSJF8jDWCXdVVVFYVQ9XumuzxmK115
Zgck5KK2DlH2nzhAIC+ZI8fNMiA42XR641r7+1IU9iTKF4W26HmYqzQw6vs2kSkB
UGtB08G7Nkm6d92AjE79Ogq0gY4jEDJkztHDTj46MF7BsWj9sB9BGKN3bKYOiujE
Z7x6eGzYOGIagPxzH6mJHvp/AgOHT0YsJIYvBCCIRbmpxevss4ltC/mJBGv5d9BZ
Fa79lH9Q58DyjLpT/Q+Hw8/687z5wqVzJuFfHnLisi8W2BT25qseoA7A+fez+Gms
GwAu5ytTwObsz7IjFK9G5b9X/RK5SCkHHMUpDWDo/qgkx/3c34k+8V4ybY/ZguAz
xb7hIjt0+i9gqbrH0U4zHkrtkX5e1Y2xAMfFp6HiwaMOX2TZObk+Cyg1+htwDDSN
bMkJ02eX+sPDq1Q7C35fFz9EAwkA9ts01iIZYtdOeq9yRsboEo4ixCLv3Tr1GDYV
6XkZfZo5O4mOqbvvSn52X9BidT6C8yT/oIcX2rPsFXCfBSed5fc1BzAsOYpJiMIZ
vN+i/U6h5cTOXo+HNaglq8iYL/BrHDwzYY+JJh8mcnIoKU6ZV+HvGA830jw6C4fI
5btR6uR+Mz6RfWj5uBxCe07ejqmewHrl3zngU05nPGOCjqIdk+2YYFp00wYAMP5g
4ehuXRcBgQFHgilW70BgvtD2q6V/HkovFwWAPOIgdR4+wzW3fTOxePOmkAM0/+en
sywEkOHdIBHRKH7Vmc05F71EBwI+jtDo8tAnT4JRy/VYbtxpaCCEB6OCnbFhQw1S
sDn18vbS4ng+94AmFQHh4N4dxCby+xcSoMKAOGFL/jnd3uyd0b7POX61wNEg4hU2
L/dWmIoAlc4cPhmiKL83kOilFxSXsGlXijG5BKL8V8CdFuM2vUcrCKOEqV5USATn
ES8y3ot9DV7kwRYHrX3OetYwG4NSsS/1joq0hHt1/5dheYI28WrW03w8wkIMSK8g
TO+N6uq0c9Rss92124tRoiyLjoc798J8QzhBCDAvixA9T8m6j4pgThJ5XWJOJqpA
ZNLvaECk9JOHG2UQpyOn7Grc0QEP5/m+h30nj+wIu2LQ5FskWski6E5p0Y3FPeWS
D0p/aLP8cRTnZrbF8T0pGmGUOqyODYQihg3OiccDkdGHk58cJ7/akUbe34gLln5N
4mqObqBPcl8IR7zXI+A0zCiT/swWiincK95Qns7T/+1EasaeHJtP4XP58kYDrB6Q
jlWILksXJ/y3x5omkVQLMzApPzdUG8eUzPA66PxtwZbABUVkbAv9XT2bt2F21H5J
6AVUSfc9RozlLG82nsdco3gPMuxhoBwPNZei2NTP4glz5CWmB0k26XdVKKB0yLKN
uQZhFyWAk+NwxWt6cThztwznlUDS15X8fh2iW/xQcN0JZzczCRl91xBX+dd1Sh9F
m/Gc2wdoBEPZzNuG4/4lmeFS7SnnYbPBGeSPJC8cpyZns+4npCNT6XZaR+6o5By3
Yp5b4buf2xlWC95kKCyXPStT0UwiofbuA+8mnxlodbF8EVKnIn8CvSldxmNxT8zx
Ao6NWa/dNqw1Out+HMQuwNKjHZSM/sQGJdhrPOgT55Hj5c2yp521xNKfhjLfxpVL
f8DH9CC2qN+mCQ/ShHzm9oHkLOBHFrusEGv6/VBLB2gu0TvQVEgqMcDxvp5TbUlA
CF/QB+AmPv8PDfYNEUFIKhv9lsMIPo5JsKe3+oNDplaR2slJLVRD3eeADPi4orxA
3oyphhzkqqMxX22Uej3HRL4qKzZInJjD3IRsK1kR/VcpGWNEZu8CI9frCOoz/i+j
8/3QonFaDDtAYpdCzXNu4zCnCUJc9iJa/brdQq63bMWuVj9ONaH8x3+11uNBT09U
AUkIOPMsLmKifhntF2g3dl1FOr8kCNHuhwfBc66PJqWwLb1yo7OhulvTJdEXM0iM
nmYKxMhoclU4ievHH8m/2AUjxDMTlN9TO6gu3olnMKzlUlGaBmM34qngz5eMvW9u
uK262rL/gNIFsRmmOlnECe+a9XqP96lG7cAH7P6ewwQ+Qc3k/+TC6IQV+iVHmues
kflEqrOjGL60wZpaEQb9vZ2zhqDMfITOVdgKhaTMWWMZnv8AQ7DFlItEoiEPIbs+
uqr5Rfi7L/gEes4Gq8VIyd8IIcPu8XH687tnY9pb4HclllgYGAaLPBBkUC7ZwkTW
4sR5jzK6L37qcd3QhzHneZHom2iA8GjhwxxNjNuTFR9iPgCF2ZQDn4QleGYQEO5i
YHNDEbo6GqIFoG58HU6z/j2EMnW4UtETUEVj82AMrD2aQCIAxnCQ/pAdQacAAk2X
XSuWDdrkz7jPFYITaaLAqzw92KejtCJXwPKKlh2V1EDYrV9JtCeGq/TIFDAmJfIr
Itro7p6gT3xSQ8xgZ0NJbGAMofdq5JkKqUY752tCvexE07vBnkswwdlgBR2FrB4o
gV9AtYzE8lTRwR0H/FC7oNq3O02boRmipE8mj3vFpUhKz7V1oaCYTDXHLEiUFR6P
iuMDzDg34b0AogJLnLK+9LTN0sLkNU7tt9V+MHWSP0rSLCTWnkQ28m5m1uwRI3d9
8lCiVfnUNnXSyXnokFj6fmah0MckaqwludHZcZ3uSl4Fp7a546Onut9nKOBdO9Fb
+pvjghXwOCuMZvdJFpQxzcRSAVRNHi3a0ktRPeFUrauicaUni12xyjQ/gtM0TAB/
yddUgMfRJhAHSYeaiJJnqaoQpUrmFmbHtLX6CWr6+hW5dj9DxGaKzOH9n/OGHiiY
uWbxeEd6lCh04+XnASw7zSfXztJvoFbDFPVa/b0Wpkqu4TF5OG/1HFyNNWfl1hDU
u5/dSyhXjaD0r3D8y19XU3dJoga5aJQ+QHqI4zHO9a+fl6siJtjHx6sfplXAj2pg
YAr6VuHMsNM2S8zhsKVTKuXnQghyRvzadwpC+jfAECdLt6ghRp8WxN3sr4mhdQ5Q
FT43J8eJ2ZbcguekV2b0IQG9zDkhWkIAlkpTum04yUumSS41LgaHPP/YJFp8uYB2
p/J16KqqJdUQQWoYpBHTAsXzwxV2o9l6jZktsbF5boygY+ERwdBJ5PaZDNOunbch
/Dd/reWTLP2cSIdtEC5ootsItKKKi1sMb8/v1kvYJeLDQG9NHenew1gmMbtmzsXj
Mi8S9zYtgnBBIWME21BfjyLkQBnzwn+iW0gwZyNuZfCC1VaRfqWxAp5scyRXAcDq
WqYByLoI7NepYZtF8RbO8U1dfwzZ3pHgB9qH7Rb9U5keysvSblKzRw9OrMCuy89t
2t74fqIxb0BbUh1Ee6UwLAjpUDo130MmH4jcpWeTfsL7TwjpgaqFgBbHPx3jW5EV
zIce4D+QFW4LZ0N5B2PnD6pWw5EYW62tOmhfPDjm380ozpQhE+3MhZ7sMjNpdruJ
O8N3lr5zFEvLPN6/N6o8ci2o1E7NZdfd5SpSsEKkH5T6l4DACQKFl8qmSaChwW1/
CbNEB6dUE+fI+FIz5CA+9/1nkUetp9S34+DWF32XVfVO3oE88/UfwInPsDs6FSFQ
VJ0xUfmlk7F/0lTTxrwrKHW3TjTtsMN0nBVvgWIZZdCfi3wXoDvKzGsI+fkZSxei
1fR7VYJx0INREXfl1ikgDJv+Fk8EUpLAqZxmMX6Hhx03BTPfFXZCkTxgCKxoyzNC
knHuu69kkohSLEWMlOieSTPr/B1kaa1+PoWeHHkOHAjt4t4m8CXm84QWAnyFl31i
oUemrIJVw1C/C1Dgrvx7k9yZTHLDBxif+cwsM9rLL6x1bKPjyXDs6aW5dCdLxEb/
yyyG2/ZrhO94/hEATD3UHmkqmTtq9V9+/+jllDr9mL1Tnu6ADiaB0kZs50JgX5Yd
uFSFtItxD3OjnQgsT1YyPUzPoYL5HoDxcw72goon5tDUqfMJ0RGtU78J2GuSUBWh
4MWzz4o6SWlUtEVFIru3WP8rTROjFIsKCtuEk+8RaaxgJ1LI0yA5LEcKNDBw261T
OZeHNDvfalDzIHFrPr/x8Rr5PxVvlu3DsoSj7+gDfrUypDG6xHbW+8GSwzgFinbI
1Mp68qM6BrRXSCTbymXvWKhs89m3XUNkvrg5zFNNeBIhH/mb8GP7EltN8kGsDQkC
uwhIDJeDbf1y+DXKYiX5/pDJOw+doGkpENTWiND3jnYozVmLL60a0eyDq9QoTqEx
FBqIBGyI0xMPKGZzF+KXRqPjl+wn8t6397XWolQ+uihce8mGTazDepqcxyQOhRec
dCIY1yd4kElV5q0bheKUNhW6ShZafWGdqk8KDNTniERkTS56PFCzBAMZ9qznGA7L
Xrw0sixaIQh/e+cqus2YCReyS+wHoqnlMAaenJqD6HxOLJ/0hwTKhzrxckdFtePE
J3zQXYS8tK2qTGLSoQ5BJnENOSCfDBNXv06soxGnRFTVGm2lTCtjx8bW1tedqaUv
ZryRM8c297jJIido8VEPzttGSxNsdpREpuyinGYeCFNowxSEttlYUBvnYrY4xzAg
9aeCG88wE1nuKlx7jQvdrCokLAB3Q6OTPlHjSQPW6/mXgHeLB4GYfgwfa1QzeNBp
HmnOOFCVaC4tagYQpsHcccluyM+YaaZJjncLX/PmsHbFIoUaZg3tTRI5aI6pkm/6
CEIRGQ4bZOzlk6C3j/qJgurhCBZRDosBWRcSYNStj48dcMKqYVivVcAeVRBVjwfn
6e9TjrwYTTDhY5jA9mLVEZCRrlOHHvQtqiIdxIZosVPE60/0esAPO+wRXF/w6JWH
kl5qGbaXAGZdy3sKi+hm+i+gO2Eshw1zf9UPapmOboeNwpB25LOIwqABCmUPI7TN
oD/XyEBgkLF/8qmbMMsgxStgp+WkG+dTsRMsjhjLupAWWSjSlZJDG7UpJTjXgw4s
ASTIh2b9zbIrV+RuE2VCG0ibqsxyPU3HmpBeEa670guPyZIYgAxQw8JrvBgEuQGj
teHyHhMBL99KoOt7amt0cmcujWrdpYX+ZMzr2bx5hdry3kwuF4P0UHGL2e77zqGO
ctI2yRujVkHQzeyHAst7XAR+t8vPwMPL9QFXDBG47yPcDMOKhu5B/2k6clklXaxA
R3l4qF2erU8VQlKgBDMJH9Cof1qSVZT9mGvQwB0wBghjWb+kJLNuHLHgEWEUtMls
m/G37zOG0MdTm77hjqrImhi0Ps02jS0FRZdkO3GS2GzCPn6zIWcDgM/MnUQudiNW
m96XyI7NF/U3wXfNd7Nw6BAVBFPU0pFrQAZV3KRZo6Z7m/cjF1DbPQ7Qa2jc2HT3
H3iYgj8PY1DacAG5wd2YQtUpaVNbhNN4CecVhwXi31Pwspffk00w0D0pdAMvav6o
nN4sFjEYWVxR155UffM77x5FE0DFtlNEFSg3iPvYfBkOR/akyofVClmTJ0Q/NiEv
PDMAI+ZpLJ/cVtz5V65vfDrHLYp28YOkXM+VOOyQWZju1JG3r5mf4aLpxppsTAl8
vIA3V0cOWM2kupd+qA+udTso8+O4HaLgSBOCDRYYWmvy7GO97CWXbVMtpiWE1QVi
mx1pefZdZpg1X+e46sAw1Qf30Cqc4xxeN6rXz+Oq6KsLDWS+ft/txSojMLIU9Thp
pWYcrKVtIT0rthIW0zy4jQUrRZB+LGTaAubGt87dqykGEvMdt0Z5xGH0yvURuXLg
HWR7lmjgjzT0s6N/5ETafTgOhfsubpz8M+G9WypLMoXC7RqDlLXlrSRd6qx9qB7n
Y4Lq6MXRV2EqU1FE5N8LnHki1PVnfFDKUMBCRC2ayy3orU5fD+FYzP/jf7xNgtH0
n+8SGT5TpNN9jVso+IKZcdZB7AAH74LNOGMYCNvcOxymw6INqvo1CLxFKB8A/Ga3
QtvHNOioa10nN0z882gxuprw1g4ED/wyTtLL55QAsOnh8Y+T7ri2XLXGzOPs/qVq
cClN5ectT98jt4YUesyR5bLAyxCyDrhheS2fo1uBT1TkrkjciqLzX/YmghXXfJT2
U0jBTUwIoX7lIjleBZoMmk7AO6wcMUZEbZzEgnk9zjLaaTRvARpb+ylf+9iXA4LN
D7JJv1C/Ak5bJDEu/Pkvjr3FVawutpmKIzqUqxKdMKcVOWjC3IaPjQIynqDQSjUX
n1Q9nZPGm8Tdjv3OWHIHr4Is/wFgkNAX8WeuN8lEfRtfhBdIyUeUpK10IENqfFF5
IsHZ8Jm182qgsRZVi43n7QkuP8jsF5PcfKnt4UrHBSQuwRCwtsI9C0bO+IY1DjpS
VKJ2aLGmDa9A4lU5OLaaxCWGg1v194IaAZ3Of/YHEBIj1z55eNR93Yq0W7PHBBz/
bHpN0DDi8vJoDE+acaVMNmyjybhFqsYMzvsqZ7O+G1U2qFNP2RXC06GKb2vRIaLT
sas45iiZxkEeRgFmvaWEgOE90W/v1lkHrZ0SbM8eoN4WG7Qy2Rbqg8q2EkTBKCb5
TalcMQx6M/hNRSQ3Z2Yw3kyU6GraiXeuBY4hqvkoNjdzL7pGsUI7C0GWB/KsbCmM
yFVjzPO5SMPCxaecGHWKH4jsCvCCBUwXdTKcJKdkpu8xZBk7yVxx7p6bS1vzBbO7
R0enSLByNWCkPX+Zv9tqRkEga9a6iBvK1X3KLKo7/ILoKdXvmeDpHCIpgToji0t0
eep5zQ6VdJFCW1Bo30pQf6SL/WVclDCM7SJcQcnNv0Fe9/8NzgM3jLcDpZMtUvfW
/NgUjfWtBrQiBqc5oKBfi9FSoJQjMHr9hi5ggU2OHQ6t3YbjN+lj0zUS9pvEC291
AmKzD3+uQ4k1bdJUK5nr1Kk2XSjYYzVtkXtMtEXz8Jqun1O5t/jFf+5JQ1oKe0Rs
Fi5LcSJmwWy8I1wlDZfazSKTpsR8w8wK29PnhNJyuugk//KBIOff8QCMxql97YIb
GXksJrMGowRcXSOFKOGLP/CjDfNUXf2NJKnsYtoVxWvFuHSmNQJkm6IbL1rH2ri4
zBMO90ufzIaj5hu7ySeK8z2ClHQ4r05trX4Wl8iu7AwGVD59YxzFIvSKMCDxGE7u
xcPa94H3hbbrJ1dHY9OaCWiSQXEgAsFL1honkvhbw7dmik7cLmAkrSLTVIWpWCAk
/jyGt0wzIgAb8Gq8/Y7rdrz2RQYPcgC012BxOPBAVblNdZU7DL4F2m00Ij8nFpKT
Yc2XSEFBXkPYfiy9pq3Sv5nZ6r/1cjECbF1pjzs5hMu4cAE4KVAVPsqaHd/ho0iI
x4ay5ANa1gIX5UoPLTHmuHXtJPcYJmBh8bZEPemonJ6TvAIHRyOG6oEOPCE9/foP
1ezv6iTzP/9/PE9LWSZd++Xzs/8jvgcEcEDWhBxMV5WyZu3s1WGJbBU+mPxOD2Qa
Ja2Lf26alNgaYvINxVGlAfF2QJc5byxd0nbHsf3YZ7McWJq0jpd8hFz04qEib6d4
w6r/5S07QTjJ7NWX652LPvOeHJ5JmGgYKOiNsvW2To4w2olDa39WHBDWeUp3h5uf
DNG0juIePTvzftcHtLsEHeBJhb5sJpMnY2SRKVLSAeBGLb4Ey961JqFJRwuAYs7H
BJ7r/IOiJEJptLOJrNNWmPRKQbL13C190aY1fz5MLjSffBM7a3CCuFAwNb0YnY4m
szKygfE4au++HQ1N5nYBe2B8euh4u8iYiesgKCHQyzFlaJ1vrfnNE0EGTBzLEbp5
k0zhHQTNdYzMNAsVAWQ02oJsgzYkJWgu2rn+Q0FYFZMTXvmv+56HZMa6QSZARY+J
dMyDMqVPzUvqtZrQsBQDLaO/wsWm6utjg5mkYuPstheJwuhHSTZMUr3c35/us1Ti
u9KS79JidW0qHdhpYxHciWQVXCAclxLnt71vm0OYx5PIVtHbQkqiZoNO14gFleKg
FySwgHr8m+l9H0YRpHcEN6SwMTBEEfeQ2+v9FnQV/MMQCyvjdbBBKnYgmo0WgD5M
dk50ThpNz3FfrVuUiRGg2Cej5bKlyOXmXtJ71tWRTJAwlE/vLtt75G4M5WKV1lfk
Qrs3mteMeuGXmoeE1g/MxTzy3xiMeeMkJZ7/3Kt7RBqVU1Bc1LA9/mwNr1KIIcVv
Ee60WHTBfaoYQza8cgxwrZ3642xEjgRSXazV66Jq3llzrD2OGr2Jv0nHgZBqZkRT
B5NCdIetkVVWIv0B8wsYUQPuqNCrgcThwYuqYyHauWHhvmkllEzrkuSbZYmWPYrG
O1/xrooxWcHnJ4cHLzvCpwW5ZKwGjoyrv5T+vWWowF3miCNu4O0TlyDuPtoIkSwI
nKTeLDE/JmpezNNv+LwqBo2LxKNkiPpUnKOxftQSnOx3bwoVcclOBdAy9GSjywzZ
Seo49gA4dM2srQQCtJfDqT2sWvfXj9W+t1Or6OP3L+O3LDZLf0Hl2tLNRw4Ncba4
dqWkkuXF4HhvptW3oR/2es2SlpxP99Gmg5MDX8J1TUIqhIL254NSu5ERanqrg4F+
B+Kg7sn/GehP8xucpYR5gSaacOyOvhnNlDlnXx+FAS0//xexcBrwW0eX3AJ8SykC
nWYZ93MFAgNbEnlYvKt8ZtnLGd8gGF8MoFS2sDf9Cl76YNEUzOeiBQNOOLsbagp8
r3wz8xJbCV3n7cyObTtjM5WxxpLozKhW1huuczcJJBUUB7Qn/m8ajl4tkzXMll+N
0CKE9UCZyURAA8i155Pwb4AQxbYfk/czjef4DwS9xJinrYLHkZq76+ReqZHMd/Ls
yTv4dhMJKVj2Y7x27dxWFdLNbvh3/nu1C+o7HYhZsOrThwRkOiz3l+J8Z54duuoO
4GTDxqzCHNntGEO3jasv7L1O4qq1VqV1hKLM4A+erbMXVtIo1tbOIUWm5N8N9dee
quVpbRYBUlL7thuXPE8GqVSIiJ27gHkj4o+X1LqQ6Q3rnl5PQpUT7wK2G2KZ7FxZ
MDaMeSdXIb4V7sQ8XpszInWWunz6kO2A/VPLQ4jj1yI8fPO3BkP1ElatzdC0QlIU
pGo3MBgg3ZqDOtmkZ0xbJi1XmEL225DzPtodsXOqku0bd7lbvocqzmK1+AMwx2Yh
w4UOMzt8P5YrT+Oag3KHo0xpa9cBF0KmAJ0Uh9fS+EqK0pzV5I50B2iiv6IvUP4/
9ndqceCkvURFIGM4YZLtaA2BJKLzkgWuSkmtP4LedMadWKqH0FeVvviyIUagaTQJ
Z70MUrUNd8AucJFkrzRM7NNV5i0/8yFS52A5mH7WdtT9H6TwTyu17M4dlLAZj/hN
MvdxaSYTWmL6XG/puh7B3zl4IMnzxZxwCJpHF6rqSLu/hYJ70neuVESLjrfVSuOR
C99N4txe2i6qNCN5VtaL8QTAjIDDDq4Mt7kdg1Jp4zsQNjAurEtoQSR5oG50IpmX
jdmpKAMdUeQJ7pAIp4/VrYT5cBkkUBm65pTr23Wm9MS4XXdAVW1nXW86R/8skQOH
nKBa1pEYihYglUT2WV7uMgBtFJFZlIyaYaoSnSiQANOOy8ckAiTf8zJb0YoOpR3v
wwgG+EWFWatTrACI09JCt4A5wOlN4TWBuojrqt7gUIWu86xkaZPy5fzlcDIdq61z
GedAEbGUfj1vxEAesJ8XooLIl/eZfBblb6auLXbmDf/M81NmOGTtzK7EWbRtARJO
D6j60UZmVd5lzQcTqX9KlS+yx8doWCHFgOZzmOZQS8qc2skSaojSLGutqwNT3hPq
HaQTZO/eW5H6tGrOfEhhkl8OmrJc5uThJWzy9m2lcOFOcJU3v6FcOH1vj4F5Zqcc
w1BaNeRauyGK/H+IjAyfVmY8r0WHkWCl5fZUdFWfGPzs7OAYn8TqrigEj+ybtOw6
PrANE2F6Ann8gPoLIsPg8zVAHA+TZylzQq1qRKuNLxByMLgTGRT4TbpePQ/GyhLO
WZKkKLwSL9iS9488RV7zD4KLVXBickYLlStYlflSwER62o6fej54HgmmjkZw3c28
Vawx+cmcFhLZ5rUiDdXc3AFYO53gaGsZoMEGx0zXko7eQN0xV3iXvHHE8NkgV2lY
xMYlchiD8AvURY0fsR9SuCe7N/9gHePwi4ftld0H/DElEJSCA+21a+hm5Ojt03Tl
I+eiajQ740Q2ftuQIaHVwN6ZzqkLUAJgT0S8cXKw9cqRYCa2pr42LS8RTbhOPsTE
Vkb9jBIceuG6TlCRTHDOKk/oEyPBxEaYE8UPF3MXqrZFyZutxWmmmDxWagLwKyHP
gMkaCMLphHam2tG6adW9fxl8eD/7b9NTNXuOQ/rWNACRkWkgW0Y4bYj8PbUY3gRj
WMo7fES7oQn80WwzI0DZKweC1ryVJ7CMA3u8V2Nh+HFVxr4BpJDgv5n8eNThxHR3
lizojITftDAOR5BrtS0xITiqZsUxuVrIbL5PXJSljTLrNrAzjQRxuW9kmVWEtvm4
YLwcsLNxe21FVEkoRL+Lsbm25VpmFGxbtl068gP9mvc0CljXQnlIJOh0vFtFNNk2
OY75UKmFEHEl1iN7m3yp+u1wrsJiWKw8rMY8MvdHsKabvBW3NwomzyZH3dz/I5Jx
RlHz7XcQyJSwH2Sw08IjWyQIo9l5DSe05n0lCztEf3B74WVrC4qY0NSXBMrNCyGp
dUAX3RMc7yM0Wo/NMc1fqxcc4Ys3bw0Dew6rHWiQYJoXAKtGmUC4tAH8FPv1ORP6
kwiwdBxyr7ApOZVtiXaa/nrLQet9orLwxnfEgL1nq7sqVcpxJ7FUkqy7TNmW83sX
2htMGNTUcGl0I7GaTCxYZw2IVO9M2z9XgfyH59hmY3FtJw9qrbiKmUed9AQ4QWWE
WbGktXKeazslBEzvMBLTZ4TGgTVnnlHRW77iNBBRIv3mArTAKEFt54QJLhkpSl3W
RxLU7+gZR8QIXWdXBi0forMYdSaC8CQaSCuwNFtLey3Ch0teHSBBxkue0Zaek5oO
CIKJeYlcnbYlaRQ00CrWbp0B2PqLvSjL1K6n+HXGwMsda8YWz6ex57WhDkM6tEHp
Vur2LQybLjoUIu42GkbpK+npj3/YFZvg/nJsGyzLXk651TGyyKmpK/aKxCLTqZlx
M4l11CgbpuITaYk35HTCXrMQRNF//aVwSdYPd5T9AeuUKbYxkWCwHrD9n//xIAGM
MDtp3o0o3bk3WELmpcxfqL83JBKiMVZY+jRfIBGaMGqNkqtXVu80VQFZu8beg6c3
gmuTn6EZWeTauewWQnzUqaKm2crlmxCSZP6yoFKhDuewmcH0fseGKd1v4NtNzuPt
oD2bWYa3nHPQMTqWVEkXs7eOETBsD2zHEbnNzsk9GtCrv0NhQhJsqMu92zBD9Hsl
o6GshEx10RwzY1c2kFDwODm11tagOMgBoJkZJvxTIKG7KZdOCJmDQJuxEjyNa54K
++Dbg+aIxnx/IwflqJwCv7XsgL97t0qicvYuSm2Vn1YAzBu/dehQdRmSeMRrzvaP
Kxvkj/Umujh5ctHfJ/XwoeQP0IhR8B2N7TQ6dFWSUqMcEEm4TbUb4o+37n5Empsi
B+JjPPstuP+n0k44mOELU65l9qZJ7nVFtlQaIhE6hokqOQ7ZGy1665/8YlWIiysP
MBf1eka5MWXPj1A4zb+YLwXPVpU43Nz5f0QxwL+7frwWet5bH/+kLSR8vCdx8FwC
g2Vr6ZwghAuPj5iSba9zenm5xqRY/PnP66t/K827wm7kmLpG401o3mE7iIe7dbG0
6AooeyXCpyo72+56H+qNMD/Ed53rDfiXW54GETWgCxQug/PyNoGNlz5gKdEwg0rG
UnSXwrDVnfkluRbJL52f8T023saRfrCVtOfCcM2KOvaIcxHovfyFHPgxyfhOKA+D
GGQjhhf4f6elnqbO6laXzcSCZ4/SkG2VeYr8LVj+iiHT3LwbfQoxvQ4eJ+ieIbAj
zJYYp3aWti16eWgymfsB3aSuBbkL/+s80M1lHBmvzt10p8godNlm8ScFLm2XS06B
RAbjXkSRgUnbRFdln+S3Qyxa3olYUWPOP5gryCYTQwIoDYsfMiMTgovLKEpEyKDH
PVLwq8geEg1ybJvxpcqWg4yk+6f9Rbn2/5Lekunq6m7Zd9qHVzGnhN0E+BfRYZ7t
n2opSmhQEoA4wm/o/JBx1HccZDnNP+aCmLpXB7Fpbj5SB30+BkEptA6LouaDBgbH
j5MchLprqFk9tUtF5dTpVipKbK/NFMhIJnly2Ah+Wsxd+MmP3miEDxd+Ppi/DLMp
Yx7xsCPI0sqS3OBk/EBfs2fae/odwFcpzWsgiRM7z9JdLFh1Zdn9+rcYJekgs8au
abv7iq5kL1Ou6BSE8UGAR8lAbkPlB/x2hlxQ+8NXrLTxEGvSfGiKkPe1hW9QQxNh
l6vYB9mF/r+Y31Z2gRjEzIutrr2Sb4VVMG10SdXPlMG4BnOsFHcmghYOQxja7CNK
VMNz8s9vKtE+ASipTzpK/tP+Mb2TdAWJSL6ferQ/vlz8+fMsjk6kh6RlVA3ZTYL6
EBnYdQeICmqvFGTD8rBzKt13mUa1C62hse1HR+sU6XfRZbNgZWvxn+sBgid4eEUS
GGFtD96pXrTrMWIf/1URmBXzozOGNkDEsQjg2jQU1jt0Wpz67pCXnc4xdmyDaZNi
FP7ycb+9mcK8lFL1IZMwC8k0+T2wAxcb1hW7vUyZxLhN9NwKH2goiykT06lFF6P0
8kpvobV11pcYO9L2eNqSd8vIeBiG7DSMGFjJEaSZDzxPrbQ+BpW1Ubmdcp3oRqF3
nnrOOniJMsBGji4iyLWGOoLAyX2aRJ0R0cOJkUwsvOBuyPBtW6/O+Ly851lczuMb
3+AB1h+iDqGtqb2YbxwF8OdKV6eL7OBXB9fZg3sv5LvzxokTxLS/gBlSgucp7CO3
ST0l5OGPDLy5zXvLSfyNs+cMzWUhhnLI19++ks0TOhN1K0mPYQfxTCL5C9aGMR5Z
D9b+HPxg8QUK6sR+6+EEGDkqlThtY1Tyh29iDJx665CIGzyJaxcV69rsoMQiw47U
gIsE8bOis0dg8wysXMnYCdQPNblrxK9MpxAD/3/iAI/d228c5UtjpBAjXIp0pt+e
80av4C8C2iOjgchLMK6FnQV2oHb4zhtOOD1dcqEbXOnD5sxczKIUfCMwzMX85S8y
kQJUZyOcCxeeGbkgSj0u3JHlQoE4g9mOLHeOL/fxgZdsvjW68SXDu3clNjd0w0Xw
uhtERyiiKxtP7ApUgj/0hNb5CPuZ4Uv56KKN54+TBkNFbBCoZGupbc9gosGIOJ5b
X6WihirWW8DfrOGku5l00fA54xIPvEmebscsuSBZPH91B5PExCQ8NKAxseRQhnlu
x4SucH8K0kvnf8GrEVGwv6RUSlg1XZKS0UY021ynXYorZffSpJFyYABjRCT50D6I
3gbORpu1EigD3uM/ZlbsAYAVreW5qgdI7WmRRSeQviAIXcdA89CYEt8UzTAwkT6x
3H/aHupkJRWZVwgGMRn3/KIiw0N3CVts22SwiRzm+4n23tY3p0CWPzkY2/3jWeaz
RGp3A7m/rbLrXOt0r3k2uRJqIfL++ze5v4gkJjlQfIUT2dhPe6To6wBbKDK5/oGx
V2JBvvqZZ8A5jVtEtxRtvetOJ0C79daGwJdwgpPVHNNEad/2k0VEL2KG0ei6cxDF
4dD7Lx9quJvzngPoYBOe8sS07jtSPxX/NvxHwWRJkxSQ6i3vYZmsme3K+iJq41do
yqieDu7gOJD48RltaGEWH9nTreoa7xiqHKX6Zdy7rz19McsO2ToqyEztkSfVs1Qu
URpLc/Vq6IxAep+InxtE3iOOXpn7AnIm6ywNw64dujk6l52Bb/MsyuZ76qqU6KO1
Y02l7qnl4vsoj/+X2bppdjkrIq2P9MfmdPqWyO1WhowQJj5YkelLTzxtiq3LaRsp
OvSu6bgB/E/aEgewE03qlKyz4/iqBuXQ+dfCbpp48MeOoed1lHIcjuWSRO4hfPLk
wbyF2TS3OS4qvAJb/7BlSOm0Z8m5hbOXqlfDSIOeFo6wEwEbtpAv75SarvVnYnAi
oXCiilex93Ez2jLeGNWS7ViBxoO8HKT+Hmnfs4HupX1pD15QPnurMQU3JMoa+rLF
/SYU0NcBRL35HxnPMEHFWaqlMnm7tgqqgrtnldgfv/Vvw5X9Tny9AVPSARCNSbSi
aRPZXmzt4uCRADORx/8d7zxxejdPSAp2A3KA8CRpbvd/b/LvCHF5ht9pbTctbUkL
8T39bZcwAQkI0HhlzT2ry1X7Ja3CXMb4ZgD3th2S1vgWyTAxC06VVUoD6nsuHZoW
z/6+anaQtBGCtJ4hZErxRgnf3NGxn5CEbZNbLwDpC0ubVPmE0DxoDE2xCLEDOePf
D3NXMrqJIOdGQbd1rQdQ5LMgtoc1iaVxlQb2aIROhZSnIdAG2is4ipfrnIT8lA0d
Je3loeNVrgGxTc00tCiQK4e8LpEOOfrUxS2RgS/WF+QnpPiUtsO81q3ri+ORMA08
iqq6D5sFs+2vFbzcEnHqVDa5CfEARw7B6FSx7Jo1KMC01tTTO/4NUN6+hD9SVyPh
CsefwuBbaSXWpeyit7UxcS3kxp3rD+fwR1AzLGF8hnMliuKNnKpljJM8Jf80rbZf
4xeJzGduLzKjUe05/LXptKf41JnXYMSKSGq7Nd1Hm769TeKchfjsOOfXQQv722Lk
HKN2MosPh0ooW02XafxdkkArtSb09mTKfToAD2bDDRAHNm3x39oQVXfujbqLoBFB
uaZHueAJanHdGY4TIFVeXc90j4rZkpCECxgmee3jsfDMniPVNgNTiIzQHKnYV6AD
OBCx8rmsjzx+WGdNP6UBxiVEeu+/0XgtVwBgKWkofdL8+DIkvHvhfOwWhiNaMpg3
lPB2VF9cVyb0B9eb3E54KrpFNH+sgq11vNeaWL90JR+KhEng9fydZL0/XUh0ZQYX
qWZybWFS5Bd3uIkLH2aDd3NgEJgmGAUEfWaCWj7/Dr2UwjJd7vo9dEmLnefOgT3S
CoTUPzvwLOj1LaSrMBUaAVTjk5it30m/2Sv21c5apIoQU7Vw4qEOJoxZebZozCU4
HTsqobqfDIAVcfLzqpkB+T3fo2UgiWdUM6WJkTpWaoXwxO5VTNWtBEwmCiruGKpk
Bx6/JIIgvQNiDZYwTWK0dI0WO2EyJUjM6FEpiAvCP3P+B4GQoBeEYnjY443CPm3e
2MdQyLSr9bdgSQvD71sKoF2gydRYnpUNgmSimITd5ZdQytqhDmmA6kmffb3EErVY
NESuBEgPvFdY6ezUtEUMAFmwiWVGAXqfILruhq/LYhYCKicmuzP+zVFATthxoy+X
fkRq/5e4cSrKMkN9tDDwNxIp9PoTY81qDPNrx6FWerKgVMeLb+F7bKy/5zQ99z9v
ikeSEfoXeS63hvoHPuzqtLuczLHLMA6GP8toKJk/J7+4tXmAqxLmySxb6u47jJNc
bREe2OTInxnqkTW+EA4302lIMVG3N7FLcFyWfM3dnDYC4DnahSftzzUc3BEvFaiy
h34cm/NX7xBQNGiaME6H4dTLu/L66rqm0HH1bl9OgQr6Qkh4MTNhkVztkI3Zx69N
5lujRKWMtJknIRxh6qnWt6kzh7QHS5xEmj70OiMHdeuw7xM0Iir/dL720bMuQGh0
4RN5QPBclrPmY/hQ1zeNDrssJqR44IZ9z72sV0u4+hAI0AFyQB8SouAtq/Yfh5ub
VMDYw+EsCWbpWleM04mD3wWdLZs1rLCC3sLgFDOOmW/I92GaTGQ7rRz5KDhFnqdh
+ezL7vJzJOwW+1RWMI98xTrNdUPHqMxAJx4M5asNsHEVzmM6rF7Z0ndFeee46LJB
OCDHcrUNkcn281eo9fokxBicCny6giE7ErFii0y0WKvIADLSOtOD3VmpTr6Kvn0y
DOpqQB4ovY97gsFoVp5yGJS/9LHV4wZZX5XDUGU1xrJGXfh2X51fWKE/9xnSDO4Z
djuyDJEZffEEwOfpIceiRoiPhtnPwEEFfskzA3fh/jCbj9JR/LrN+iost3cW3ofQ
XLPs/z5BetZ0gohkTnThEu6kLZgMzEsdvJhrhdSY1eSmJNIdFhfZ+GqNoAwRcVkp
SLibbBQSvVwsTmH0qHfJPFAJjyAJFXVkYIlOe0ZhNu/KzlLb+mQgykbPAYxgUOBP
Bj+RovXgHM43Pljb8o0TifQVrM5bX3aV03c2puICbVJRnn1Q7ID9avPYNlxI1ns1
vzw3v59mwIiRfhBO0Pt6MqVnER35RVx0de3OF9RmIeqZySzyR9h3cOlj0rujt8ng
7O/rb2Yq1bSl2PaqpLIjDa4vXMz00jQjD2r1mRiCNIncFGlWaUFl4oyEjn+pd5Pa
hxBX0O8xKC7e3gp9DZE3Hl75B6kjVNJ2fHgbzg+DybC7H1ds9uRTJYiapu1KXxSs
q3gwgJRSgXrC4paDeJ/5ZEo16ix3Hr7i38Vmnruai4T/L9zw6Hl4Z81vJ7KLKUYA
7NB0+CZNMs/pXtsXRWV5rKfy8ildp8xSlENngFkxxz6VGk05l3WnD1xtP7crAmmO
egFTgQlUKGxP9ZbB9DBukebr7jgKaFG4oMjbr2ygaEsXU0c+YUe4X7chjjUPmO7G
DTAv83HTXybSDu1QWS4N26SlaVfELMD1C3ZcGRJzvg5022GM4y8QlDnwGqHnqEd6
l/JT+tQ6SieBGj/qZKIbbkApY3jjkNlZVexyczyOGH/48/2p86JntpgFXcpKDIyQ
uD5pfNvdELiufr0VcUaU5LNWqTe6GdxSpMKgvts0HO8QSTJwA6jVQOWd9wmqEhS6
lDhOu3VFgNItCYPM4OrtvA2v1r9obetsZceJBzha2CKXXxI6joJKPTx/Pou5xigd
zU+iyHQTW1Nvqw9FZcRptpuVakcHumke7bJxqfvcEBtzs+J21yj78Y59hUqX9DHI
dwKzk1GXfrhVjr8VLv2kJkGyAaq/LSC4iDdlAAdyNNQ1q8NDCJMUhOzML3PbxYmX
Jqj6WYrd0okNuDceHxVeMOmriBVEA36HxKh98V5RuJlrt0AHu5otF1XkeKlmLPSG
X+k+eZnsLrnPr0WFce3cC6RDkhNZqRYhPTHZ22ofIflL44EQu7v6PwZsLt9EujhV
iSGbD1LtACxUdmxuOLWmkdNzpBufHzOJ59q15fLXXILz+Yigo0BVq7n3BxOw344Q
14JybXe7ggWeMGNOTeThtOW5XxRfw+59nvID9QoNvscOEWIY/v1brAPeRzg5pp4y
f/nZ29uKQ3QkdWQH8lfztbp32HBLAPddgl80tVuW9XWUB82HNsK6ebFTOKzQn0EE
15ZAj48qp4ads3ekC0bnKej57D2Wx4R0Cmyk1czfeGTs9EuPgGyqB0KuXQ1Ne4Af
p6H4BcdRJTc2OziBqIqvKeoDdgCY+3xYI5xIT+sohxinMXG8xh/aCES00Gs6ISgm
/wquJjor0o095R9xTbq5CU7OeF5WiP5gz70B1hjEH7sXpqaLR6BcbrULMnYIvUGk
2wzt4dmevgX/f77zwKScfaXQAYQ1uHNRCFV4y/uXpkjmUlH+x6p6ICKJO0frpoUy
SBr3u8eIR4x1u3AET8cED/DqLjMZjfncSZsPWZ5lklYVGmgrFznIwUNxwcOhLDHF
UCFDnbxa7lBoRqfQYGzMK9jO/5R1eSVAqJNTfPSRfrsEMLJJjwF3JcMXLfp4B5PV
LJyH2rYs3C3WSneyh/RuaFDqZzLyLqLR1daErMOMFRtl7YVMv5NIuUXMGrdvsIol
FdRtkOjZj+oCHftBKPm9rZ08i1wpvlqMSBBpTvWioK8x6bPQc96L7zfVfADL9EfI
/AYcbM9F2Gzho8oeMqa4Y8SdToigQoIhG1/W1oFRRgYfoI1K+oI7pKK6Vx0wYdBH
XBxBGmb+8Zc7/3wwJM9HgNioUS+BcpTVtS4G6d9Fr6jAGq70L4lRXMKbPJpVPRq1
XmOD2lxiRw1QHrJJxqqacKJeu3Xm6ECMNe0DHNET7O52LvqYICuiZyXo7Ib4GBtv
82SXAbC7Sozxm25g6bI1ryHnWE4npVqygVEZOEuSo8KMHIUCUNMV5DsMn5RYDFmW
DuG4QRnM2CXsSCRx8CRhbvQgqIX+qHPW2MQvwOblW5SfOrkBNSKXOEQcQ4BZs3pD
6mCBFCKwOVLNClayWNrqaMkL4tkUohytjbSCn/Xl3Pmg6gwmoluhF5KE7ILsERF9
sthWSY/TfkNIdbpEyNzoHybz2J509PJix2Dac8vUApkHyOtaa9JZs9UO/pVMP1TX
/thw7JOj7fQLcwPCZyCmpEsV75yE23qAb1lzrtiR2HDdoaucGIYCyY4KyvjqV6iE
tOz0flQ01qwdOdx3XHzpuOL0FfT6+h9TbwxKekWfL1LCrlfmaCB5G1vHv9XpGN05
HZl+6wNOUP8Ia5ZuRqGmgf/DxuCWuVJmTDQDnDV7x8aHcwJA65OiEw69ndNq71OH
+iSuqfqafEb8Wjpc2XIrdx3gGF1rLStuk4fxZ8RmyRMNiyY5/Kk1Mc2QohO0u7ud
rvamVF8mbgTY2chs0c81BOIqlA4tj6xmR/EnZnQifP+Ba0lWID8F1Z4eG1q+6CHt
q/ADYX2yIn9jz3lL53x6kk90frIdYfLhzaYHp61BQHHkq2IdJN6TfGQ1IY5YWYMu
CQcdz/fX58pB22aiduTP+JmJjyu9dM3XpX9iZuGr1tsxyLv1YisYtJK4LWKfkPeY
NaNj7vxd+Sqn900Jk4yyXSSrdrkI7wA+Rx8B7UEspCTmNQ5H86WZYIWCVWTy62Um
NV/0TlptFf+29UDFxoYQE9Qby199nxCkozAXpA8w+U8F6bnWecjNagqdeHLvlQ0K
TsB07vgjW2eorqu2jADV220CSKXMx3IRC50Mru/idXBkvkZeBA+I+wvQedBARBNF
COBPjYeLO+kWB4OhuQB+LdSpOtu3WstZekKtGh/NTx+nzXTGosKE1aHc8lEE0gvu
5lGG4bSakeWmumaJ43CiuSa5WnmC80OnfvzJIoGiqezC4rhVnzK+zJ6oOl8FZgtI
mUkejS2sfq1wleTn8r3RfdWycYHU/2hRBP4eg5MuPMJLHKDM4GUDNWMw9tTIlncv
qESU3qm5VZjvbCFflTekRerTY7ampmrTR+Knx162rz2+ho9q9u9Z1nqKK5QdfGzb
cWjqf1mezQHyxb8fRANqTYoNlIE+9l4Ubta0rwC5ESSvayCpg96ODeaCnJwYLgwD
tFo1seP8XA+pmbGGIWt/0C1t/qHj9UmStH7znIFIh0KCqi0batvo03xnRIWP4vVk
I0LpMpVE8txhUAv7Rw7mfGw1fFlRBaTIW0Ac/Qdd53O/fB66DUvzSz7FwB0BUP+W
ZrVI7TB1mO5Yh0lSkSNapLDuQIZBVnCZGV7z6JhzPjCBqORWlLcaJxv7+F4y0Qyy
A9L4ntefGtxfe8ArV274WQb8cjNFGQeII1eDLX77+WyqkTMkpV7XH1PzOdN5ftjj
b7BJv8aEp/afJGeiUwysxG2f5Zt5TINvTmpNBQyizqTqlf/gAI1l5fEjc6JxCkZS
xPHB/lWBKGllUnguh3DoqgLW9jJSRO/hjRFYgaDOcxR9l97l7jFoawgoNKjkExSe
cbrCBgCfWexS2RnIjPL0ej27iHZiXi+rvqqMEUxr8J8i6rPbmyGnPVu7fL45vHrg
9JBw02lUemhQIXgbXx0bMiCHOITFDY0vbub1iOkHKQ/qXejhzwLJPJdM40AFatoG
OYbIvW4/6oj2NemcPkCV46Psf3w1WsbLQNNclgXKPZ7WjQ8g+MJFK4y4njjp0v9z
WajuNUVz4gmJOb2EHXS7y5Y5/9cnKhT7zj5Tj+fqLLQNms7X6P+tjM8jl92vKKsn
1va4/Vk7fQFNNVU2+NYzHdmKfCNKwKtmFj528AbAsbhkKiCmqnhAeK95xPqF9o0U
XujyF5zzqATYZBlYhM6KCOMguB8gIAneD/HErX/qlk7WQ1q2YEzBCqIqiBVucbg6
2DN7mNuCJLyHmaAD4pjGzB9eCCRsgy/bVuf8ApFIFQVAj/dFaBq33gUrAffJdiaV
xQVVqkILe84icJDlo9h/WnLd2suDqzmMJrynLi2YfeXgMD31Mo+4QXqHE/GA0xhy
z8/pU/yISiO26Gc2zSAxPC7xwuDPKjwHLXhQTp8F9qm3TpODz690/BqvSYvuYZOU
oKtJ1vP92dLqJJpdNGx98SFKjg7BYqR6Ka+F200gFXmZhMFiJK9l/+1lITcUi4me
tHDA2LroOXYSPvbdeJmaAS4MQaxu1nBmwdsTP8L4EWP7uGnn1ZbWOuAYIgkRb2EM
lELW7Th1pvQgtH/tKvV5Kqx8yVPwxL6gWD200NVxNuVA4/8pG0A0dhs+puRomHfC
OT/eM/qTlNpT8RS3D8DhEOjNMnaFuFwVFFLR1Cx1uwVnDeCDM+OINb1ci3ulkm85
QYwlSi5LDdCmh6gjvG2r1v51/DMImcra13jrMrpgNBxdA+Johmp8pTAE7dgkhi3y
gZQ3gXzzYyqxZUDXTKp5V8wTf+HVmGYGs7ON+nhLrH32Yc31s6jqaRmdBaZOuHC9
Cr74S8NnY4TYdNzmkQ3ioHz8x5tmcR8MzG1DJW8RuybiL+0QttHETJMv6Ipk14MW
`protect end_protected