`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16560 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzkZGdUrjzQR9gfRaWjj8jjKPQ5zYSxUQ6qNMK6eBQEmY
8aarPPWMufzi2OM10fFeRo+2ocuUnaWsAq1tIAW1m2ZvkBSj5CRp8nRC5CRLxczD
/O7vO7YqEcGnoJkN54R4lhlLvvuPtsTdo1sr1pHmlhbMczP8w/A9bemnY/PcOB/i
T7elRLV0FVFlocwaM1gM8PXPfGuk31WsIeo23mdK/X0Zab9dD6qkWHVUMf1QggYJ
GH0eT9zeC1V/JG7P4EJCiwbmVHqQGkI6Gu8IMEr0TjDioWpvpD7r3NJedvs9+Rgs
TZc6SPs2Az7VLBn/U+B+k1BohZ6DR3v7rK1fgBDXN9gMEw7cQEphC3+/H0hdhkLv
sjKeBqCU47ZcUsTRZPBkmuCj19zwbrzFOfSkt/9SiXa+q+2igJ4IrtNsgtcBiXxD
wvNp1Ynt58rEtt0iQw2NiHIo3c6iikFez054Eesa9TmiaM/cd4oc0W20LU6Z85QC
xwLVhhXLvi5tCOs4sV8j6/JSUhERDe68KoS9oX+IqZCHNYlXoaVZZqiQ8giBipdf
XpLQ7iTjpU+V+GndXYMDnC0TotsfD0cU84y7OWBig3hhOrDMDKxrPHoCfOwJ8mB8
ZETjiQmOIRoyJ1F3H09ZbDYxQqPKl95bUx9PjnXzZKj9fS5N8Xx3B5OMqjHGQug9
wtY9IwqemjpDJvIj9zuSxrmkOOXsqfCojEYssgE2HuwiSGCvL6P48ytlmYQh60jA
OsR+cyTKCqfdE+tAGmcUUJUG/Ff7h+QUG2647SAcGVn8ejKZ3i2p5wwcS/dbZvw8
mOJqG81T9xSP/z1exYRyzTbI/OcKOYCYH9lv1dTdKglURM/SK9B0lR5Vl/d/Sing
c/vj1F0okzgwqRXWDpG3WUHL6MCFuu3GFRFM8ase96Nm/gEKQL4dOp9Yxwc+qLMy
ApqV9nfUL9mQuovielTHWNzWJO1RP/pl04Ycx1Gu4UY8u5l1dfkK7zoHYRQYK788
kTATf5S3myGxqIaAlGUqJN00jAk82UogNRJMi37tKgcFl5F0IlNoTwSGELwqp2oY
CgnyQasfTR5oLbV+ClGd5GXwYZi6lo2YrVYHEgudA5KnQqMUwLpL5JvCQC3X0K13
b5j+Mr2qeRrKtQdX63+1bF20b0pAlaoHp/xK0oIlFCl1vLgm0CEwHUZEj6+R1iS7
VXVybURizVg72uxYSb76JtZYkr4I8/airVKu8bxu6wJfDE4qY9OJKNzsqtY0KpCY
HDleq9dN6sZzTMKpSsq//zoNmSiJIbgBgIMqqpHX01rm8kiBef5mslbraV5UYct+
aTAza4hEHbh+wdrzEraCj/MrkegnDFy3FWwMNCiDnUheschh54XTea6D3NERCRAq
aTZEqdwvjYLWMeXhXmaax435T9eTp0Zvsabcju38muXyFLHqFSM4gTbJnjV232+g
1h21yFbJDaZel+TgeqLGImGDNah9suUnc7PVdJJFdhFB1cK7sqxdVr8X39/VXBAR
8UnvFo65spVHWnYm/DmZLqoNyCa7gY8i98w6BELpyrEbX6z+6b3FikIHlq5SINmf
pLR97zqZlhiRnhL7TW9pkQbv5DXafCrwlTHDww6P6SdZS5vUV3PPjjWHF3Sk6nk1
k0DRjkgjWcSp/Kp9UTJvFjKk3k5slkkk7Q0mGqsLn0brXHCOqrVIoZEGFfSZRQdN
1ZkTGxb185/ki0EfpW1iSXbk9HoxmRg037xQr042glEgC8Iz786pSkXufRDv/txC
VqYpUxGPI++Sx4zXMY6O8TKLsiG1h1Tg7A50sLXO+l8Lb2Jduks2OeXtSFuz+ojG
dWkZdpr6acut0GVQoax7hVQbWOxui+QcjVVHFsg5Mg1o6rKtoa74OARwliF0kxsH
IrA6hZU/Bl0dDcNS0tZw5eNK+ZCTNtyNohXje/CGOXbdE4Db/H36iDoq5NC2cyX6
Ig9d+RWy0BGAV5UcE9Y8SfUuoGqGdpf1PdR3k9NJmQjUa/5vvUxER8LhUreu/pFY
y/bLl/Ajmyyj+1BKvqTzaKEIpuFF1EcQjogj9S9RonOES1TBGcw68Cx0u2+uBfL/
KbkbNSYT/3iCqyD91KN8UpGEtEqxwpMncEsD4gE2mThkicLk341br0Kg7zvffEcT
/kZkrOlLysoTnULL+KIsNLY3pUQ4Yci5jsQz16OhIRXxh+/jA3VgsEeXRQJyVFUR
P486DPN/FXLQfCYpRKjUbnGt9L7o9cAxUh7S36VbFs+XpKHqYq8BUEnNp2CV4T0D
9rGF40bZfONZEsv3/qyA0hBdopC2/7vww+Upn+ZaAFRHpMK2Ku4EkHJBRIiS9NyL
37EGqToLKNQ+gOLT5B6DIHI9au75bM3Pi2bX2cIdKe8yLO/Z+wPZnFtplrHsVkgI
c95Zr2cy2ZE2dfUkKg/gfi4WTDWq6VeS1R6llXb1MnS/vY3WAisyTSrWs1ek4P5F
Nk7XNz0PJO4Em8b7UC0joR1W46G+MfVuujF7fbVDxmkTDkUFiKaoHrsf1iEJh1bP
hKJy7ua6BBYKIORe1h1z1KijcrlwDuwOA9KXd3js+dK10MedHusiGVlfdNyvfUHy
MyqmJTVVftFJtRyljZByiLNFbEbeGk7ns8ZVl62TMhoqrWacqtLpozQdEKlc51O5
DJ+6IWovGYSkF0xsHV4mBBviOQtya19DO8sOCmYgfyXt1jLJyEuvjlFN3dEnQNIC
YcmkbxvewBpKOaosj9/pZUD8vCh4/dA8OXG7smjHSl0IsUUYVRTpNIxlHbiAv6pK
JfuTphTURpDdDnRMVXtZ3SpCGAazgLE4/jvdCiv9Aq1ltGNJF6GTdJRVDyhj5FB+
t8DJ7eiyLysNjON4r7JArdNTjNG4dKCbmp550zv+5rX3WpYuBZHT3rPOpbxNOj+5
FsUgcWpofga1f5zQBNVYxNZm8aO5w0u2q2wZC9dMDWkPHmV8ohb+uWegGgQtl2uM
C4WEl9vxnFnrQF5aolYlv4sSwkBTdLsDxYs69pESDx56J22a1hJwD422TI3YkKhb
mOgKfDywUDdKucGGIaqIKBzlyx1V5p7IOooE+TUiBMLJRUzx31bTmyNM94+5+fEL
cngc/0gw4BJjvxXJ5MxR7jh0wM4wpBQxZ17oQJ42gm+MQ/X2It0h7kmcS/a/T7eF
x2zcl67bwVw5zW+xhpVio7Zy8W8su5lbw09ggeaBQ+S3M1WwyL00QqmfwfE1cQvP
mR2DGoz8zaeSZ8qq1SlodX1tHfZ2IJqib3Tsc1CDoH1faN+oezEO8IDCqNXPC3Ab
Z8TBc+wt2GNr8B3Zvaz8oEA5i7ctUx4YKzUWL7LXf2XCkqQxJO9q7mzF37Iho9OQ
Xag2ridIBuR4q1kgt83Sdrn7ilCbVoa7WMi7EM1UVoHsfwqoCsnWelNDo0IPKc1s
0ZzhnSXYtmdL76Yx3ashzyoR3WIHU9j92x6M1ixj+E4+ueeLHM0qfoT7WFklS4qT
vokXYVhz92MOyrhTI9Z0qXPVO5u7n/naQ9udLg7hqBMuiQDbCXmomeMwMYtmnO8v
kat911QaCD0J7GBiUkBapNOL3SIy714ingtRGwEHMjhhVPFQBV4NdjzVu3O/e4Pm
FjVjm+JSF2JMs4vrClZxH9lbcIJ51RuE8D0Ax4CzXAqwnqXSBKcEX+izsEs5n1l0
9SPifY/xVuKWe4hQsM5O5AYLdO5xA3LT3LqnMT3YgNTfvPYC2sYOR3fIGYUyIZPp
OIaWLpHuuFX8P3bUMLq1kAdhJTFnoKEmQ52fnvxjpFfEclbLy6ycH3ctXjyv0YPS
r5pK+9KWIlpK96XXj5bL7xm0o9IeoHCqret9qcQbaDnh0A9mRaMgu6hb5538B0f7
M/0MoQlJGij+juGtajkPNFGNGU2E1kKm5MFvlUDF+4pzt2SZ4qusVZA4U82SKRTh
AIzpZtEZsFB+11i9YDU71wHWVy3up8YEagie8WYtUjPFb7WlExUhkpgD+Rq7D4Wy
zAd7GfgFA8vYZjx2dirQ2F0rfDl4YBiWIyeD/t1fmGtvawbzGK1JDHMj1155KgIw
g8/4LZpeoshzaUjwIjll/9LNR+Iqb17MW5QPs1y982JJNG/BwI3p1dyLYCYtXcgc
Agyp1PbcrRwoqBs3Dtb9oi/DZbHUyS2bCfbUxMGPZVYhA7WpqeY20VU/QRfpftkU
5ijBN/jqvqtK6EALxP5icJ03/TaBHl25oSZ3UJ2Ww/A2jzIaaCldhoQhdXlzMwr8
ucmBQRFfQR8GEvKiiKDC5ZQt3gpVS0/dvCLjUkOWrRmhC3vuTB46v/J8PSSm/3h3
B316ExM/WaqgjvuUHw7SbvXFyKTEmOeN259V6IRVEY11x1NahApDGiQMz5UDnUlw
3gzQnijyrmU8PMhHrmly8DYAexOMf2zKJefCBGeQI6Nc3OWripuon9fAjHoTBEkA
SByoAHMhm9GrSl8KfmNGI/Mfq+QShZYjryEXFL8PvY+QvH48uaR0y9lU9rUH8fGX
4b1iOmzTt+zkR2jsTig0I1fmmBkcMnxabG91TmoqepS1HmU7bJG/bSYjiEkpEWxF
xzLXSJRmwfisnolV4XAHUKCpAKspEFvnKm2ybhl80OcJ3Mq4dTa3dVXhVB6pzSLT
xABP0mpTJoqWPp14VBHfgOPVzVoppoZUb7VdAqYc8dntopFHqokTHucbh5t6NmQz
cQe777v+9/hJJkWQQnf1IxgGntYiRzwMcvnBe1K7ghpWSQE0XWIy4D9m9w0ZcrTZ
yWtpYHB6sNgKwwOejg8m1IwRMqTScsTnABUkVWcWNKV8S9OM1UzPz6yMc1mZQAVm
P2Qom+SfBe+CaWwFcZKgBcMSrBwgEIH06FsaFymne1a/maoYR+jbW4ZfqGQXrhSZ
q6iYwwL7AVDG/Ad9aNpQYv7zpxweljg8I+3Ph4N8aqNzp+y4hnKzIltBpXYRkrWb
rPrElg06hbXzu43SR4+5Iz5bOP3kaWMH3pEU2Tu3xWOZ4dL7y+NzzHaSQ4kgEJPw
ZfRNAz0mytZFGes+DVR1rXhtyZWkt196DZ00W385pJmaXepM/1HuGtZlUCq0iSM1
vZljIgc2m9ZqzOUtzGAOUXpzcc5iUU/zWZ+9d4ZMdf7sSVcY+dP4OTAob4OdhRrG
bwXdxUBD9cX7Lkd/dTiw8B+GUa59DrRoT2qXlspfgK6aX3v2kt0FJA5dm5SQjbec
fyNjEc21fwRcuieEiQFo9GglPNPpl4HHemfHVMQYS032t2RfVN9gAf1lwA57ymU+
sOoCn8jlyYAjfIohuP568xFh6QKDQQnicbK98boOHyqI4tPgfeUtfaJL9FsMxtlk
t5qPKhwPQLz6WFjg663VpTfy5ujNMboYtbhDaDG7cKb9V2AsowQsxZvqHbzstomK
iSjC/iMxMfa1j4F1J1QfXoUkECXj/vwniuQpGHXXB3+49T4ShA53ZkaVj17F21v4
cJF3lKu+hN4Rx+nfyYjapmQz953bi0R3ciVSQ4BZ2z6iWb1J/IWaG5DFR1u1F+Lb
+USDQgX/RBrVcfrJ012qLM/0amBPmJn2Nf2lPPOWZgnPRFjC42ae9QbCnjTExss+
rr+Ut9N7wKqa2Td/P9J0wk06v5aj+xy6VYmZpYNRiV5Ze5uyOXhWWVlU2x0RK1eE
06pIzOaC5L3XTSGeo3bCF+Ov2fw7w226KDW6D28QP90eo+vr9qjxqz00TRgfJ3ME
Fgl2DgYGSor5S8LcR2atOs6ThdwXfYHZMnlGVSOlF4Zgt2N4s1Rpwvy+HvAJyPk0
qL2DwXruAndQHCiotHrC1bs8000b7g7mB5sY3lOmUOCvngPXRqqk+xsrOdYBwyjR
7VNBWfov/4PHpgYri6TqDyyjscHgUM5gTpuoFNpyKI5OjMjVXMTi6SvE6PNnbUeH
6447bFqKSETRqgWN4yhMVpRwlRjfuX0/9OofkOyoJK02bnDmmPkKY1CDvz246BVV
k/VjJdTvt6nR6BXPgxJlIgIRJ6+dT0/7wszS+a3tV1501Atl/kmYTznU9/gtwbXu
kvzGI/jLpgCNXm/+c+QHEDzUz9UHdybzIR3YkUjc9qfKHOCUUCuKcPMHyLKhOwFw
VrDQYJ0DYgsPuj9DK7SXfgbFH4Mm7PYadgigAxR4ALSBpNGlkonvwoZjWIKcCZgy
LOmG0Nsi0ML4rC29MWP62lXw0s0OrSUzrfo6Ur1xzIo38G2WT4oc/QYdZDG2T8KM
b+OIzS/ayJhcucObQfu3W04/3lF7xDn7dUeyz8blHLrInZLc1qa+9Dky4N1Lbrl/
vCrNmYwJdeVC0YYh6AMj2hf7UKrDk4ODmBO895jErClG6+DkDEXB1LFbApQ/pVST
wKdxmrh7qiPh3SlWDW0Xj/1SSWr8oi6mXhO2KHo/BZ026PH0PksVGjAbjOLudSSA
IYbvqO/OtoSTMr3qNr4UGiycPskMsemZrYmPeRO7q2Z7gkYnFU4KXEWsXYrmYXuI
gqwdqttDRJeELIx3MQlavf0zRGwJsNTmLfMUQDP01CoTzhAnWBLKbuO9C7AeTD0w
PZctlCQITQuRm8u9l/dnOoLQM9GkYRyGav/U1J8Hww7sqla3LbIjQ5hEJpiqZNNd
OOzTgc8kl+NXPzbyYJzTEaBluFLufYS2RAZF18eb2nBPkMgrXDj0/jNBenXRznUf
cyx4IpU3jsbB3ei55zdKfWeAVkMSi6NQ/kPI4/6/EpbhhSclqVW2DqjrFZlBKcAP
XhrJe0NJLSMBAs9a8wLsCiknCQJ1SAY+Bs1/9OEtatOZQsguxp//XiJfI0ETzm8z
KUU0ja6/vajZOwvQLzpFCdUXtdvBvDf9QH2fShe5EcFfGPS227sJ1AnrFevlem2h
g8rhT1KB2bvTG6aFWv5wr9AIZkrCtq4e8Xxx7DcgiL7h/L1T1kmKQecYUIvLInPD
HBFN8wpVq+6BFvnGldtDcdiKi27SyhtO+B0aGCM5BsUvjWjqNvBHxtmVCuxxEQ+p
ZjySnhiaabkCt/Yarxw1S16rZKqrd8yJ8GMwch7yoTeGMKNfwbjglEaDd1CqaK4Q
d73blOGfc4FJoXAUIb+NLok3ONJeqMLO/gfvBcJuiL58D/UjM5OYbD6FPqECuFus
dRAIvccjgLgqxL6AjWZKCG2qIbXmc/ERS9vbWoqRKxeEKCGvZtPcLvsLJG1jcOJC
s/yOeSUHrCGPckfvxO1kRi+iBhcZetQe5T8p1T8hm6pU9ALHdQ9U53sNi/re2DVL
CD0Q17WrLlDSgyXPIM8Q2AvLLN10mUjYKqeKDGM8ZT1ejm8kMZgSc1/Buc2eYr6E
ej38WhsRvqDNw+TOPXZuJ67pTE6YhBaQZcFQpi81wmHCbTgBqOGmd08bYcslopLO
tAjDHKEmaycJjxrl2cInTKBsIQNLJfr5keG1DyyJz4izzfTw8HoA6M9tlQosQTbr
5uajvv2PybnksEfTw4cfqDzsGOzjKQn5kgCBX7G1YxXzI8ikHYtWX6p8uTgaB4Fm
vpCekLVwFRz/i3qEgN/wWZWA9MrVi/NN3ikhQVw5oPuPvoZLhgWLK/t0Hc9b9z2+
EqgJ/vPJEiyPFZyGViw7+ubTSl9SgTR/bHvkVpWQoU37skPqwLJp6OhC/vIsjJu3
+eh8Ut6m8GZFHLCm2xtIx0K07+VxV8RADz2vhCmjJSOepzm6uTZz6X7Nz8QGpSUR
fxYsSaeePs84BEaqFziBGFt5TxE/lHW7q9YwMJ3JGXbUt0uyabScYEw6Kouhb6o8
ohznueMhuA5a8+qUKEfRf0hQRO6vuUSddi2IfyRgTWDwg9669FKgnfmwqBLdtsA3
1QeAuUxVLksfOVkF6vZ8WuXefTelAQGH7EdVOlS2IhMleXPL2NtqFejUnr+ThwJo
qp369KQojkZ5X4XynIGQ5Pg5SQvPPNj/hwksCEdd8QXW1lqwl51B31pUd0MIeOBd
/7AN+psoKf3IA8iOPzP87NDYgn5G40DUY2wyrL3fhh3uFSPXewjJD3OINMgbzZqd
lSaO60HEI4Q2BWfZTN/m2E/PoGwzCTA0lagTIol2ePVUFlKumNIsm+exSA5owTG4
He0goRlpNU6plXyhayKpEloFsv243esliJ3+hrh1IA+vszlNJySVadylsUCBlmKy
PKKt+MVToXiMF3JdflekWIJqEdnfjK5t+uEyuBdaAjUdImn8VIUY26AkBO76Awzc
rm9D/vde/fPRGGlN9Oan/TpavdU7y8F2Cz2jMU8LALrczokYVACqvm+vKdhnctfU
/TTe5HncF5f0gbiShldUqsjbZBbcvTP45JtIR7fUVUo7NScU6wFhsQ21krXyKhGF
WUAHvkN/kdWPSJs24rK35I49Qow2JOyG5gcpNkEuuYAnbApNk0ZH52DVuoEj46wx
n5acARExdwnWvciYEpIGjxkjzaajTApL+WUIMSUXoQLCXFxp17UPX3zNhEkT7yoR
9/iRqligVVZloEKk9sWU1iDduZMvTINm2D6XdlgJqiO+c9ZBgToFSNu3CN/fb5GC
1WJ41cssPAUb3kRNOhyok+wvBnhIOHSlVRbKbWT5RyGqA1BQCLTbp2Isr2+IviSu
XtytKoAIn/WKezM9cxRB3p0Hba2mDd+rzJniCnFlqjW2rV2uJ2t7WPfbatk3zjuH
ke7/F1gzP6aaudIZMFg8OH3/38m1dYbihJ5mcaPcvOjaYG8zT6kYpRvBYOfq9pfA
dDXRODUJBsJa7dhm51+ZwPE+raWxrIZWqaMKkfmqa9Qg7Db9HsGVb4OJSVBkxi8K
PFdBVnEeqvreJiehPkOJWzNO695DiltcwEtYQYw8/mfvPJ1v58vjECGeD225AWKX
tTed/C08jV6vY3EsaaBTh4PXolXC5n3Q6cgbLO4PVD6dt2vPQcdnviieRmkTYJ0d
wBRn06zYRlzEdT4s5B60Cjn5RWzV8kJTCshHXCYqGDHS3WFR58Cd3R+8c4qihZ2/
PAuw1PnB0tZjNegaWtiR4uQ7xiWkxCzDrmmjuazciF+0ai5xiDXvzwhFpf0cmrgw
3jmnsg841Drvlx01dUENh9FderKJ/RPg91tykdJ/FeATbSTf/rIOGtBhwfHQpAlT
HM/nOJIALDEMfxRAuK+EUBCpx+/BbiWsNIINIwVh6KKfBo6l+a9qNTn2o0Pox7Ry
ZLtvYGBH1fsJmMH4N9rk4piNQ03hYJBC+SwymBKFyeJyQHVNdHhj7gBHTZHe8Fm7
O0omqdhMigvh5K2Nebj2cFH1lsSfsEAuAmhopsny5z8yV4CwSaUcU+uba+dQKgLq
r+JUo/RZ6OMTpJU5uIdZyFBRWjJBf81KScB2y53nvSBEQ3e5JHvmn5Ub5D6Ry12I
oebgovvzTxn3W+wDR9TSU3P9VcTUu5lEg/Q/JglDj5MGEj4wuXzfXGAdF0cuRMJc
T5dKLeN7DAKMCQS9iEX1+Yhm6sVh0JKwvlyB5Ae9mARRCCWAZgKDzJBorL6doE2F
ciGETsg5MdvVwbK35SNy5lJWCdq7d85viDv/jtZTMgb3oGUFINtyONul03bgcJVR
fahHANVT0eJyd4Vp4UrkOLqrIHkZ8RpF8qPwUWGYSn8Y0uhcUIS4j8n55SyhryHN
m+8odTYeM3OX5KPG8apaFGJDdtVgmSusQ3j4MjOESSgxzTeDZDc4PzEPwrmBAGMl
5oMvWTwD5yCetcACBmUbvulEIKiEOe++i8rSUFWDHG8+cUXKeQ30IF+jvcKA0Gg/
WdM8aFMet9SscHaPqi9HxW3cTIaEF1YF8Vovo02xyD3md/Rax740CDnxD0Ss79Z1
qYB8bpw7+/627Oa1xQKROo5wrIwEYmKVC4Wc+ggh+RtSQE6zAdJaqInRHwDnSbTP
Swui6Z480UoiijPMnBPL7PD8IkEDED+QR9XhF/5gIKsVpItZxyV3dgwRJVrDXz5m
26CCROZLwXEMmO5Hd5whUiEr62VTId0hRz5bo3diYvggRUfoF0/aBPoZqEONrhU5
ej6XJAiL/IDtlkrxDC7ePesR9fJslLaf8YHpFNUkle1W+eBaK/djNt3PlP6U1oA8
p79VxB+6U6o4PRrwwjQlz3A2xWBdvZvE5diZTD81F5XPpY+KdVURcf7USRD29kKg
ImJ8mWroWFuml3CINZ4X2HjnfCN1/8F+Dpdc73EfDgC5PzWJBm1kFfOZ6SwZoWeR
X4LkHgV9pqk6YwvNbJq4kdp0ZC4OHiVDtBgoA4FbcbM9MmO1NjMg8SfI+ewylWlA
gTGmhaCIONxlVnWhhW8HfDtEkhs+olInbnQek2cEIHlz4QXYxVNu/s4JEHXPyJ/J
Hddq8efXmLB4hixfJr0uz784s2A7uv1br9piGVPpqYZB/tn9L3zK1X3GI790DKA1
EPEyh99Khxz8zRkmjlxsbOOE7dnbs/yIv1kcEkFXZXrbjOzncb8BdoAecK+To6QH
lgWjMoWkmmCh6uvP5QtjDa7afSsKTwikbSpIanzSfzAMRnf6aM/xH+rfzO+elu9L
laEpb0QgnOPcLOScYVH8lt8rW/Y7vd1Xo7eL2a89eLvlFCcJUaJdw+BQJfujDujW
x9fnl5XAQGOInlK2uc7ua52xWT9HDK3ntYS3H+8RSJsnPirMRpYAgBMydazeL3HE
npmBxRkOxXctlWxDsbvi/Rm3u5S8FcFIcpUGwndS4sD7vGAHDk1Lae+uLBm2SqUr
BlafBBNKI+FCGvl0frieMG13AEVoJKBMQ27c204qrmqE4TqF2n2bFpTos6vSNN6u
mTz52YRxkhN4+xugL9/NgBi5TYXPq5D540dGpWbTx290h/W2HWGTvnP7/EisNew9
bDNzlpgKamwtk6tSY10GowDF40T4gnlqtkGMno3XsX7CTlrkfQjDkvS2hkrTp31z
R5XD9Qjex2h9ReiMuIvGHePBCXuq2chrjnNe0fuaLV6qU1ICYAlhvCbUVRSgj5/A
W9BEqMPIzgynvPiAgwCJCZGaW1s4WAorlTVAcdBkXKA3zDwOIcW+mlafNqPK/yMd
jswx2PAWbTybFWyP2SqBceOdTwZwy2KTtJP+diiwA2uTZ6UW0gKS9h2peLDFufHV
8Wnzmo2GBJoquzUmu7XBU+l8on+zbdjB14u3ng0QJ4Mfy79f2TYo7knoGw4yVmrj
F5hiBiApjcAXXjXZ+A+6kKFi0FBYLXsQaa89RSAraALTSiddA5Wro1/BaipVXJsZ
S+ehQzAIjSIjmnhi6dmdBJbS9NUSQwrftVcgs6uISewm1Zyiyhau8Vu+anZFKNk3
Fovzrk09TbU8aNBfUBDMCAGxYb+UoHBVV4nbNtJrx3dRcwLOkG5YNFI57+xRn3hu
Fwf1PlcSKCzmctK+3vwpICyDZ4rKc/C+J7n7MYElmfK1YuURHS5LI12NK89eRAv/
iUDf3F8H81/XNqECgGdOqWZgOLloMd1TP2k7M1KCiRTYVBYMgCBtaDp+goIOTCbu
wgWJeKD22H2V8rtQqWsNOkj4jG0eLQ8bdGBsoHoEbrDXl4QRaCRrw7IiBZyKjM5I
ToRM7DLaVTc9qQ5k7WrIvOmNVu7piGOvewrLiGWsNyra8z5/uI7xhU+eRLLUmiBO
hXCWEH4IHv9HkZA/bAJk1mheLsmp8zCd8jMKMX5f1J0l6CsRNCR5uIMyd4/lU7Fl
Cl9kMU/WS3zuiJB+R/QCtBlIVdjffhEhJn9OdWt65giVK45IZ+y0oMs4dn0S/ZM7
C+oy2+6bvjond9oul4mWJ47Qm6ZLkLVFNPxm6K3GTr2ftdqBXOmQDaoxkgWKWUzb
DfUxnkZRDaM2ndxUGZdTx2Tn1DL9sUSa7pExxYAUDtvDMSyUdXaswsIs+ffjnjtF
XqoLyC06Te4Z6rDVXvGsEclrjPtcf+t4NfJQZGryfT7vH0mEsBH7zdd9OluPxwRI
yVcm3Rv7PJ2L7GkWk8/IhJ9qpQ/xFeAZ96kV0OqAKBOoxXpT8rB3qehk5wpCzNwR
X+iLfncyRJt0kYC0Yur7TB1i8BVcF/3c0s2wqSW9nx8HiaZDbqnQrz43waQOweWE
uIoanBS07svbcaPjzAUbvvMnCSzLRrXNLScR6P6WkW6hj+YvxAYpcrwdEYprMpJ8
oSBDQrAZKfTDvbiNze6AtRBRGVCgF+o+PjjTqz6noO5xwvyb62qf5bcp1hE1VWIG
ugEVSCjdsOcFUnPw+oxCXQIsdxHnu8Y3ZPQlu+R44ubaBMll6E7aBi0f01hTU9aA
jz/XY0ZRCuD7S9vMaONLgKBjJ1/6In5TcQ78Ry99Xu9Rl7cOCggB7cRxUn1P77sI
EAsZRP9HpogktepDfTMTMCUwDmA8e4HzZJLAZCSD55Y9ZEcbK8JqFKXgr+PLrhy7
PBfWW3jcGnNBzFbuCNK2V5giYieoBgY3htuLziIXCtaJqtRcKIQBUYH81lYHPg1T
DSOIBm9ygZTKrgbAycriZHFaN2aXuqqPBZBPrdIRQ/lv6RrkSPrJ/ziure5gOKOh
PZ8lVpOQc7S5jWaiZO/oDaQ21X7LgrRt7IZYvPNnjoFuidJfptoLwuG75Kd1OaaD
fY7dwbSCEDbaG6Nd+XnkSFoXoy22FqdoPqqNmWgVLcQD7M/l+nIj+z1rhnbWR2vZ
HjapZ1uMIvQN7QQLDvrsVnWrYWX9Y+Qt36rfK5G5pJiehZbee/NQlb+ynkAueWaq
j0pSpoTYCXin3wATS5E3y0HuAVPyNKysFlJo9UOd/3lFqPVI4ee55f4tocsE3Lnf
eD+DdE9pYXkjiq4l/VZ6bEVXVTtYCIO+XivfbQw3ay/RLVdClDD1I6uPTq36dUtS
PBOoe7ds4eLJIdehLanrgft8rYmv6SUhbs0Hn+9v0cQNbOmEzi1TjxA4Yb8nMi6H
VctaUJqyE+X1nDLV06GmCpmJoRrsOeQ08cmf0lKRRCb9isgP7rHuIt7GhkeJHy0o
SE3L2TvVKQVW4YP5CCqFmH1/CN3x39iXTQg+x61YqguacYFUwxUgbJItBkUXJbyZ
OC1ClWOXUbT+sO0TlRyON91XkNrsRrUcvo/Q1V5zhGb03HkbdgW0KRhCsbAHs8TD
61AZM3h99qT4Gf07bLHKwSVEbw0Vh4Sf4A965FyNlRvvLXNjLliBeQB5n9g4MCGn
KHPTJDNwh/BxgDEUqS29FhARVeJvtsgXXMl/Le6H0xaVhIeyEfrOGZomQE3E134C
KLWZITVxKl9SZZ69QYYpbH4x3c4XYYlRJ4OJUkTTuVZtDfoE1T51GI09QjrdERKi
Ho9snnHTHnSGmi4fM5ToWB9jDRv4zrKCBTDeXmKXbh5Dx5/yp/AvnTl96yjs/fGf
igGh6N5H5V12tnx5MMyN6IkoLX6B6H/nmhlOfDE0JKzZeuPxF462ppBi7TUCjXc6
kDWT99PSCAo0jj4l7glSgBBviuzuLgcV54REjWnuiJ1oFZQYqayAaow5PJgZZ4nD
n5lmRqawd61gMmKiylWgcVFktIwLSHftCmWGsFuXK8laeuLvRKx6oJFroDd+G6Vg
HcQKnVNEWTT+hTtQpFBGZLl5ZLbnzpeyIZtEJbdwHbgDC/MiEg7so91ifXKwgOpj
OOXRauU4kjE+sYvGslb8cpUi9vgjY/bLtBHbsomTWl4rSEPZMc0h/faEVbDRig6m
Zt3bujKHm/MO6DAiyQ884WnHt39TL8ROR901EXvM1vmJd8XoZtHrDe6iA/pxKh8e
UqgA6CzDSHoz2FPXqofYNGcGP6YL7n64aVASOocXarepWEXCzN59viiPU2JRH2sx
iseMMpDg/7sfXgCMCdSlEYvXdfSJNjb/zkAVUmQEKNqWHLY4F9ZUPzE8EpACYvh6
uvLR7EgyPuGzHhh1Ilrj3zzsauz1MhlD6ElKDRkoezbCXvzGJFg121f2b9Ozbvyn
4dC3ZJdsKnPg3AbSesLhNqLOTpwMgCrX57WRDe49fhzDfWzeX9WGZ2XjvVt89rjE
rsrUpgiWGv5HjsB3Xqf5zBLPZ6rhJJXeHVM8DUmgQxBl7KTPHBGLmb4F7512sBpx
h/QnhTO/NRR8NKrjUD4phlA8fF7ASHF8wv83E8wsLnsie9187/g9uMp59kAk/KIb
f+0bHqxUP/nG1rhQgfcMNcvyWMVKdC1tTEZR6q7dri7oDVsMX5Z7HG4HadH8Zqmg
rLnN8vqM0MaahHypfuidwYPKOOXl30gjv/ZfoYxlS9zpS6XGAhhxDyJ0BycsMde7
F68r51vJad5kUFm9fUIxajbHRH+JxRbgvruPcUu/kVynPnObPx32AF0CdVTNYiDX
pi7Bh1lCaOHNq/g4YKT1niQ+xIgRiw83Vcos1bGKD832q2eZx4dtGPLuFCx+yYnd
/DfJTd3nfr7xTl9N/l7eBDQvRCVkkRMjpvhrTzfVF3IWjmIIMMssjZGU449NQKvT
v4Zt82Zk4pImj9pjBrmUJkFKwZtYPxlRwT6OGab6FY83JPGpuTCYe4dmSmZ4W2VO
SNy6BW/vb0dELYrQKaPTlfxRuh9zmUct7u1MOLph3M5KC7ZOMbg0Wvezo6wKdS9C
b8FkFwWv8/vnEP7QSvhPqfgtRV/0CxAuxKS0sNevafvu/rwItfpH9nM4v2g5KWKi
IY6XNOrzx4cbIcCcJRpSZ24/iGsdYrdtZQhzLl9FevgKulWqf3cKXtzvGw990dDy
dJF3y+KYs0B/Pd0ybAPXVML0TZPBNMJBbb3fOOo8sdoR8pbUYbqNXbZeWVqyPoto
sUvym0KXFS/8oK2vh1bbb2Lr+hUotXJrBmL0MC2+0jOkASAzxt+DedQx/6Pp4hOn
INiy48aCauVSuQtMUba4kaich4MSJhaMbEdhmrEWyluCWkiwbTug9ipZTTTMF9mn
UwTS9r2MJH9oA7JWh7n9zNx8HoRCY+/g+VMsutAWKu65e+1VSOY+Ty9KOjmHML5V
ToTs1V51RdTapUIXhHuP8AP4tq02cpPrQqs5Q1yL9e6iMBOC/MnPzeo/6xCqF4CN
thLOoWieeo2mfQ4GQekT05EwAgJgAjS0xXCzlOWK2KqErBUA8g176apiC9jKXfmO
EMb6MDsZ1fFMoa8QbHICc8OloNiTLET6TYriE2YC9qYbiyAEAvcl5yQWjEzFKC0l
pT439PRJZihktSprUv2nrufxaWwBP7W7WwvB/ZQE9eouPePQp/KITu7S+6Bztkw9
pPKiF53iVGQEXwGcLXJXKaFKfCAcXxHcg9robs/09l2L2DF+uatEL2XqxSDpDLVG
cUrzE+y39aDe6XLxeN220Rxz7JFDHyV00RDvkAPntvZcBZM5vV1brS0n8AEenog5
vkTkVTApa4YpidJ+g7hRwObssKV/j3Qlbe0ul1uCQpuc2P2n4+ZdC0eZRafXF7SO
JiMJRMxdvEd9K6o8kqt3FzralkQDWfwhxRVNgp0Dasu2JALIwFIX871GZw6z7wES
TVU7d7sEHWNbtNmby+FvDBgNnl/a1w4sCf98LDfHKYcEpo7e2zfh8ucaYuDCBKYE
gJw5HQpy8SXf8dRqbp/BmM1DVElixB62lCyFZlqbOlhmzUni5NzYaKt00HrUU1ay
KWVs7OJsubEsdmAAHDpxmJ+GJwgxsjROvo/Zv9gGV0oZM9R/l4p6A8S3M3dthSX1
P4X2Xhfm6LZShTW1NSkGA97Gy1QhVPpjUs1o5KJDtMlKQ41e28XT9lWC1i9OjpTQ
YEF6FWKiCsPUgcfx6xdI1qE7I8NX3nek9wnauj8wMOqknrIN1q7DtizNNzoveBpW
xZbhqetp59dfLU4bWdVTn3RIofzlmTgzIZAWNJT/0oC9ka/lf+K+hlGqyp8ced+Y
jFBfwNelMQcDEZqF20GM/lxpk4hxssvb3aLj6whFczwbuFxkXI9eaG6cUjCseS4R
SjE3HyB1yHjH6VvoA3lmQdqqMxUZjSzDlNaxQDETDZEIddUD2XTd5JCGQZzbBnu+
Q6q1kxy/eG4AKFxnxat7b4f3456608luKigJatDV9qJtEVhk0amYTNDSna/Lz/YD
SO8AhwPBvTQhPlubIpoGLkqlRLAlMPiagwdP+FIq+F2qa4993SmAxaEeGePlpWty
GjaPVcNcLxHLRr8IRhq9/VhwxO3R/4XG/161XDXakPKqWdVkVk2h+km94o9uCvcf
nF4rHnnTQpX2uqeY/K/CJnOrQSbVhAg4d5N7tLRd37IoF+nnZI1j/TcjxkQq5DR+
KTBKvaN9LrkF9rU9BFAxE4hzh7a9S5NZBqx2qL+3e9PH4mA/gLi++TWDb48P5Rtv
shXmJglS7S7tNH/7Sy4h/Sb/ipYJL92sbWmDDxBpGYuJl6tISaZ4yF1eHkJTVgxE
6/7Z6v2JL2SGQAS4jUebHZJ8wm6KyGkzgmK5wJZxQMfk3A0MsLttc66Fq8AV12jV
fVAlLxcZWc/USzfbeTrg+ohVMS3pVbgn9MF8IPHEYu41MVvNkFnv0VDZMhX/Rnwm
72gYcbXezYUYgMmDm2QH5/s6q8cwPk/82YJFich9oYJsX69XvR6cOgyFA9zlXIBD
9gukFXgK3FrBWasp8W9UARIO2u2ct1HC6cJbz0bzxEITORmqD+z33yjHyZJR8Qwu
PbejTlEEXiCm9V+u0JyuOXAOpzuUuRKPibmUaivSwyvbOLEADNTEg3yvnxg1nGeG
bgoOALedEP+BrzSnVqM9P47zVUIqyOVpxbOA1QA9Lv4ndfhTGSybSeV+0HPDcRAz
ySD9QlNkNGOKmGw3CdhAAtZYabCv2KE+eJGhKqYrOKjligRafqqQ8VyyKYDIIdE1
GuCSBE6dD30hDQFkMF1JqBlf2SQTkdzGY9WWdH2JFHgcDSL0Pb2y4T6VFuGI/ktz
jFHmsLiprFRZRj+fqZJVsWIBt6BZphVvcOxMGFhEMqI+cpsJrL+gZ37P3vKqNLug
Bz9mCdz8JkNQgmM3/NuKxfsLU/FAijhzu0iJkCXi8mmYOW+Ppq77d8VQ3udk9r3i
ChqJWFgB2TVZJmq+ACmNry9MnOE9gry+/n+wPk2+nYNKmamDP/+PSxjtdAcup4T5
gCkq+GkRf5JeJ/sw2AqpDFESv4DBtyIAmHehfuoD7gnBNSJmqY+CCveJKtQ6/HLn
VZM6uD+zobjbHFHquP6q2Ss22zKvbllhMvKV57gYmXvLHP0V0E0O+DD08aPGUmms
BkmdoyH1R3kYXz9ZKIYfoR7W6JG4IQtylOs+4Ci0KWtlG+r6wgfwJxyQkI4YqKC9
yd3i3syj+ds07X4MULwdSOWiQgLtFms0Az0fzBm0IIGCan/H3GhCkSgQrYLMa77i
ye2vbuSukqYyn+ZdnE3ZRH4a5ozGX0y4w708OjVF3yFLPuFYMf5VluvHz9xPyRlN
k7p5aeJ/ts6O4HCVa9any98QAkE3gwOem8QzipBAW7bJnqvpdK4ro++Q1ofI12uU
pUd+YrKcyNlTwaNN0isZ5DKbHM29UKnlVZthm/n/KNp0OsTOxEFS8eC4gbkG7rTq
VBRx9GC7aX91mt/1FLEFE1FvS3P9fm2BoMKpf4GfXy3/FJ5lQe/QCnNNx0F6JBEr
u0Bhl0y5feNO8iynps/Wsu0hj0INno7a+iIojzkAkZp8Qq0O8vy/78Mel4e0MLTv
yredeLRVDqcKlkyKV9DyTgDoZDeI6II7p9+S/+XopQ6tR38VND2IBqWSyA9EJTNS
qcRo8icrtN1kdpNkyxSO0cGX2oFXiL7kFhB1xRt2TRgJr4CI8UAUh/KNeUZipe4R
gnuzoh7eMWZvpKZ6+rH/ZMdmE21gKBbkONbfBOxsbwcoPIfY1M9rVG61upqTIx4h
cmFO4Xud7PMrkehORsQjXTrGFWVHfFNlYAFH1W9tIDEdlkf2V+PoXXM5zHVXXAn7
H5LyrpBgcdX7JsbMGhprGbsPVqPNOaSLc99q+NCtMObUyl/tmwoJBf3aeckbSTTN
xhOzCLfLu7iwR9ahAAWQqhKNn/wLC55NYptGqz7OjZ6ozpRcidLVyIIWPI5gL+Wb
xxw4n6joPxOiv8L3ZlJWwwz3/DQ/2xhdVVm0P1MCsKUzjLRkygSY1Rh+cyTVAJhZ
IDs3Pfjyr7qvbzEe7IcekRNRBpJTnDazKnEoFa+yDWbWh2zaXLIl9riOKi62nSr3
kTes7iRDZJWIpibxHE1KAsWiavMBCFvLEmv11Go5GveiaDM3pKsFKbYgus1rFau7
B3xnc8u9oKihSxRjQ/b9IRpfCV0IaX1Sih/31GDHAvewxXOj3yNTVNcq8uBN8B0D
I+Z4uLPCVgr6hclKKrS76VuqL4iq9dlo0LDS3rGoH6BOgQLz0GUaXEqKiUbLp2SD
yoY2SXH/BlstOkvn/SDR4o/2kwwUcxU7k2qzqdnIsece8VqerMBQxElgg5MMRC+R
eRz3r5T6NXlNj+oJNw26h26J8s0/Yl09s4JEXmAti6MkqtRtUdD1ZJQyR8FnJue3
wdJOKzU6jpnJD8Ps7BIWTmmRCqv0AnzsXQ6c8fuDTwbw2DfEzqwmi81zsa5Rfoh6
DxHUyksNs+MSkhZihyK2tQquN622ESsF3jRwI1HKo6wjkTafL4sFLmQ+NBW91UY/
BrBRAbk3EEsL5+zWoscYi3y0aW0HHPpGUru5TGkyVNVOrxowV840chCNERIDpPVc
w5H5O3PZW/U4rBAr4UfgVJffEkpqlyNSnIz9998Jka8iHLQAtR3uuDoxExY64vej
CyWVMIeRd30oEb8T1PRDG6fTevYJc2ijY+brTMsn5+dd1GdKZX1tMEpbK2ZoUvSB
DDW9E2ksfED9q1BlwDN6NRBwh22qeIxuu+K/BOUDt1Gp/yTtnGAFIqApemhZjtxW
chu41MqYExlV7ndPTwz4VBOWcpvuCoKttJC8VVvKLZdGmNLpshz4JFS7WVA264pf
VXOpvt2w3FuVz0J2wfFlQlLqVPsWzM220Zb6yc39Iq10FF5k95ZEJjFb4MLXiEUR
kYFdG+fzs8xP9RluDV4vNEriIvF5qaWxtWb4kbTJmJ86ck8BgiMqUAUZDtIrj9lV
sQzZVyQOOM6F8wVLUNFmXdkVmnSV0z0boCxSzkhqvLoGXOsU1f98+xAJETbBQjTW
s+Hq2JTYz2lw+lLz+bsLiMcqNOlFRpYkpcqIJXpI5HVW21oa5vayiWcOLuNJPQqj
Oa5es0qMqCNttEpUGqYWKR8scnh/RPq8acVOR+kCwfSNOOuEh9ldmJVyChp+ip9/
WTDOHj4eStkfzCgNW2z6TOjywlY4mIx1fYrc9ecyZpamKVNEJrqT3sVqw98bZJnE
W5/qu3PVzHSqcVds45cmwLmaOGhTQ7d7gqdQJc4BGqwUq6+8wRVsHo7aol7CAmrF
e4tcdllqvUOzG1sYSKvWXOmS+7A6u4G5krxb94pw+Cr3vQ7nausBqEwkEVhy3EKa
LWw/g1EgdKeFP+8LfU2gWoBHH3QBSsvPyDM5+SvTqsEnOWpLvkw63YjXEZXSnjOS
BID1gwS5hZU19C9oZT0N0aU887XTFhNxmTSuCUMoA9hrsaH0vB7AZ9ynxIuxNFDY
/eUamRmEZGtMAmZeEMdO7YOmKdDH/79zsJnMOwMQhZBNpoan59fXHJH8keyOe2l4
7PjlgDBEC8BxBVvd3qxebQxF8gjDQCT+0E4F7A6ALYSOWbAzAHwrw7yKaCSQ23tG
C0Gjp2Vf4DYVJfKOj1jVLe+fVMjITznPa1yJjbwGyyBymB7phUCGonKBtqLpmp20
UGnwlJnGvwbIrsdDa6csjX0xYKsVxD/0AGI/J72PwdxejBcK0Gq70JnFnWtNid59
VCx1zc40ALsNB3j07yARkCYitKWnkcdkdsmpU6e/id8fuBibb8wCw1eLhZ39U8sM
IsLxvJ+KK6apQEZsU6yKuaj80NydrvvQeeKq6jS0pegnrRrFu7Z/02rJnxcLJt0F
mHEh1M6/N7zhmbATrm33Ob7N7EzYzJwKkro9ghSVjUv/Tl97kJ58p47EyQ8eHeX7
Ff6/POyaWh8XkCdyqB7bP2ZHYC9n3HObVcnnRBI4mcRbrq+Y6ynM0uII67AI8h3Z
m/NDKwkpI3kwl6afCmhcEMXMsqBpDc4b7Ci+HFfxYcU5qKpftan9M6wJMhl6Kk5E
7UV6U98mmRoDNSoVmQDQsXpy+o/zEOJHF0uIx0DBhnPXD377HdDX9Wmu9Hgn6UU5
oiYWxU+Ul751xQkaP3glun1VpE2WC+NNP0/teDcFrcunmaEx99xXjlaOJ+JicWYz
3AGyro26pPervxCVYElAqIGm9XkRaXF1e7FoNgFzXLrovXLgp+/zMh5oXPiMQ/B/
jeg7kfb9pS8vNUttNfr2eqhBdZAOceSkV7oZ+PpAbR8m0tpAaKWaa6tDlQOb8ObW
ocH3ApAPMUTFn0Ga7Uahzt+YExVG1Roh69Ip6mJoZl50AzQywYBsqh0pZXCEWGG4
Fsc2TY0HEyshlEDCrCT9J1rOSm2xaFnvoLDej2IHHtgzgGreNXP+wGVYIkfNYyPc
JXQKUhOQqqj4PDIHWwin9MNcRtVrWab8njG3sgZAP8XcSp97acA6dSdKI82KJZL3
gAJAP/CBFJZ13kQaeLqV48z1G5sOVlpK9vbHLXmQgdPebRPSuX/oxuBZWtYgYyyb
9rALeVzM2oHqC+en5OzTKRVCCnoJxtL87IiclmxHyhVg1rdHKmPMQMs9TTKVUwrB
qjN5eJEk8ypDyOHYjKmMmIGcKsQ2BKbBfUla2PGSebkd6N6FPCrbyM4cunyEPIvG
ojet1B57SxAlJ4L+jI3H+zcdrefb8hZyXoqYHzTWij6lXphfS6iJOBV70p01U15q
I62TwJ8hNAJ8wWIlLCbTeG6Ow5LITB/G6wEmnhJAIwLFwAdCOwGOPGfM8qj5e84x
Wacd+FE+uJhBkVLQfXJ753QKxqqOoJxJwxiyT3e6BeuePHmJ5y5XA47gin3/g/yC
WwsstlgcEDtFs0xJrYe04DgecPkqyG4ltcz1SgBhKs3LYkjr3sVjc7qjMWWxP+vN
d8QJQLrsI5QXuV4CrW5hu7m7O5vHy3DYIW+SQ8fIu/mYMJRGv6gHFDyVqBWsVA54
ekGAA6WMjP3w2mIoCoUgPD446gR1EkfhhZbIgKkcTQV9o9ktRYmxkz2TnD3Rbkec
+1YFi2mRmPy38CQG4b3yTIgfhJ8fJuw+cAFN3aTJrOHz7wJ1Ray7gaNNkPAvWlmW
sbvMbiHioWjMKqQHJ4fw5Rv9To2TMOKcbXBIYzin2W7BUJ5rJpuQL8/sB5vcH9tq
uQaa35w+LWaXijCNCWzWlcCfO4goDJRFuDBSw5QI8IuVhtaJ2PXcmjiuDazgJYLj
4H1O76KGO72O3k/ym+qsr8RLmrOWgjF427xGKYxQqkwwDZyDPHxUB9gx5Kyqq4fp
rwqU8peXjM1zhfWwr1t4XQnpCjoU/BuVRmfiukoEI/astYmQZXbaBvyI/WHsXfsi
NvqmqrKhmkDtRCerG9FEbd8TJu1gIV67JjGdyOIfmnLyb1aZLshR2EcPTzmUpIEy
J4tTuXUlVpfEbl+LaJy+/jGt904g4pqEFBGi0LWQb7D6lRrjVhT91oUAQkdVa6Sb
ESIitxHhanPq403zhsxsov94oWA3XpxQHcq/z1X02eQSnIgTpWlHMtBJ9hBQMBir
01Et9syM9QJKZoDv3N9QxpmEX/Wr5vO3SEDXMHWYuxnERGS8bLPDFGE5vj/9qFjK
otiisvtlR0KXUmIrsy5T9VCWyw1ExqwWiSozyt5pRG4XMkkqxpi9tS2fDiaVMaXj
xl9mvUHYS+wCcPGjwKS4hAl0qAAUTmmP8uu1htTvyuO2tsp9hqDtokPUKWhKMmgF
V6iPC7mjqZ9zQZZ+seKEdxUpKRmNoRw1saPxB1E8npsIuHGBD/JfIO9JlOQHwnl8
`protect end_protected