`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
gMcHP74wBZczB0bB0IzoP2xg5wC5NPjD/GsvSQ6VQgzYAsanETMwwsWi4yhFtJwv
5kY07u0WerSDf8woJ0stqW5xF501W3JLIS8KMiCOd55RHBOnavjYiaaLeu7oUCmB
TtTS1R4sO325rP2zOn9YwRbyyS5Ljn+PzFZZUmkt5xMca3p5NGqKtZW2dV6Babni
5HlLuF20Au601B75m2nv+ZRoGSrpkNElxoTibONmX8gBflpIVE7BehhHwaKSucEF
pp4QQ5zZAZjEC6aplZepouGVggAulz5AahlX5bf4opOVlB1J7IrgyjENtw6ysQ/q
DzybQ+ipztSXBGhmcCVU3A==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="jAI3OJE9Sh00Sic4PtM/KZ4WjwT98XM8AMZrZsQkxWQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hyw9IrFLPQsjvXplweG8O0lkaSLBN9Ijv4B5VdTRt6ipKJT9Kzsb5LxCKvkQyF9n
sGPOd5i74hRHnkHfYISGkfxGJCa55ieOyFShOsqTKRLxclm4oja9vTIey6yFm1BZ
54IDCG9h3PqfDiTD847UCSMRvFssyycwv+BRHQMQlFs=
`protect rights_digest_method = "sha256"
`protect end_toolblock="BnLuc3jxknmZOyxfJK70E5kp9u9O8IQ8cgkXv26kHA8="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 43504 )
`protect data_block
xABArkLxBOK6xG+7CdOOiGu0zbCbHMrEntFfAZEE/xRFxZaAZl1QLkuFI77OC2KL
XxG/mrHJzO3taVHgwRXNLDdc8ePbxbAiQfzV3NJLBO+gsBjmIymaCa480cPNpHLx
I+PQ7Uk5spYgOrbeCMwyHMeNH49DbhbU8Hr6xtjBwfOfQg+c5FxPup+0gpoWm8y4
ujvcvYDsv2JvupSMIIPSDmK6XxUPWLPYev7QbOfEYA58EznKVCZWASQsXtl2lcFz
VwhN99NMoR67q6G7qEWiX5KEj02bcsyezGZWfKC3fXtjiwA8rHSa3Cws2OWS/OEi
SETK9aijKeY7x1ho19HTRo1mfIPf/lLag9Xbwo+0zg3D4hxDcnUZ6mYg50zSbmQG
QuPUlLKncGkJlqr1H1VuL57icUibSVGMwz9StjVfpdE1tMfZNv0GZWqpke9vfazH
u/rQJ5XBEij/PB2r75qpZeDA3POMwUD8H5VvP77P0SreBsZAVPXvrUEI/wYSB+3b
aH27K8m522mPFHrQEbG3KfYieMtrOEL4PuDoUr5NsczNkjCvmtniN3b7ThQw5CDS
3zs/NZdKSwDLS0ktwS2MY/ymfvULcF5oxYaXq8LekH4CJ+HdQF7bmdX26XiFmYk3
KoH2sjncIdZto3lmmTkYcNpCt3JMGoR3PwcJbUmd9HXd8n80ok0fiDKw4LLSCw/q
5OwCcix/5gRtn9cgVuMSj8G672pZt0ZXHZhZScOr5BduW6pM293sRpf4gDkDQTeX
5Qiz57/1dsJDfHJS6HOvHqY7FZAFFv07BK9OM8LmVR+UMq/nzlU2FMp7PRfIos5G
ijmsa3sxHid6+zFrb/7fKEtM5b7OB8NycoOhWY7kOqa+ybSYznlAobBHq0uLf1Xo
JbJ/t+vJeeRk5jWzzX5dqGEi//9epk6UXS3ZsHVU1n4s2RA3paCAwhHXcdHKIkcV
OEvennrSuhw80BvA0JBFaB5xuxYcqD/M1A02EPOA55PJizB4CAcPMjvpqcVPaioy
HXivvn3knoXwaz2qGg2eFBu3zYGi1oyNYvLzgzzbjlPS+mkXEem9IFASwBWdrPLA
GSEDaZubAerBn+7pvsXNdmi6KIAifcHIJYtYzkR+6tHC8sRe5L9PkOR9tZL2aW8U
KySTbrsFdiIaszp3D01M/sbEE1qyVE+SbXayYJX3BkLZOieePaUl6KQQ8nFfE526
1n5nMlvBTeS6xjk1esBnPf6G84WopP+OJhOVmkvG6QhkHEPJ+/DFiUO2a7GSNVpE
cfy7oo7oauCKdf1/cddYqXJVSrMvmYubKV7VGSX5E358B+igxA3Mliyi9zWLXcoz
OhpLQ31k9VcFrwDoB094ZXcSqUYZShhhzM1OiWUYZgmqus6JJFjofdI3gPaDD/9s
jGEmoTjQJ0sRKVrh+abs3y0w0z0HBseBGSE6Ed9JFMQaTsi8cimTfSH3cGSroX9F
b+T9Nc0WhLZM9oC1MFaY4X5L2pkmpJ5RVwdTA/yDJIBnp1orU1KTLxSRs8O3Sha0
JOVliPsmNjWay8KFrth0rzoOzNYtNy2gaKunWqXnuvjnyqn7hbjrSZ2NCa0ndoAt
gy8Hgxtvpk8dVkcJPPrGPnIUIbiIHI9L7ygFFGnbM3REh3FoMiIQtWZbT+smDneX
1jyYpDNC77kh2Gndc/QIq+jct5+Q0jmU5aV7yBdnBfyEPELa180a0Dlg6P8R6/IQ
V/Zuu1Apf2T/bv7qKHc5FmYkSwp2lfXXmhXjb0jY5FHmsjTa1giaIytSH3tuSpbp
ZLlnFDRLqEOYupOUXHDqAwF+gemuOxp3N7RMv0wMc0jOpM2yckolPYAE57VmD7eQ
YmAh9QEtkfC2cK6Ca04xpQVRytQkED+l6zKBV4fJk6renYIn+xnfLUr1NomRVtKP
pg4JdzDcuBzXw9PeT8UKIkK2Ohox0DUCDrAzVFuu2+ed2kfmyHqo07PxA7ygiCSD
h94fx3GDf2G480jdOlJiqX8q/tFYXpCssxutGJ0smW1f+hviPvIxPSgaBZW4czqc
AVueypFvgbWiJBqZiE2bthSfGspKfdt7C62vOg9IBjvHM+R4GyfGFgM72B3lk3RK
HOFmdPriFcSJRFaKlSz6Qj4giYYlU46bGiYuv3qD77EXRTlY56R2J/SOL+YtWYJT
Mqc3WyC20UKviBsqfn6hVwu/T+SbRALrL6dZEwfSdPtty9vV2tQBjrThGPsT/UrL
XNOheISGqdhn5i/WnZWMe37X13Uw18I7LcjL0jviuCZPXFssKWsghtZxeggRSNP3
IoF4jflb/+fj22C7qTt+3/ZQ26o7zg/wXqCfEsbPBpBoIj1DFrrFzTOWKQ4rWFse
kem5RCMmvs1GpTdA0fR9CWHmbzUsw9BT9LP6BVJcYNH25sQ4ovDBAXBrCkse29Lt
iEna5v6/rVbgUqv6w+usvorAksZqnUz5hLuDj8OLXrAacrwawnjJAEmZN252LmlX
+3iMNxs1hsoUAzazT5Wze4fBcvghmOM4i37HvvTyHJ5lrOmuRGHrJZMDqqOuMTCL
A/eQiFBOdtoq2ixHN9wo3+pIbC9Lq/1IXEEEOUr2MrgqHjs6ATWDLBzEa9r/Y3c7
ManGsK8pBv/RYHKJH8XY9rky/4777znqVmTnkdRstGWmZVc6mEpMIkHkoy9ERBiy
TO5ziW5GrZZO7MzKSQXRjk9MixBSt1mAgu4AjIguLCnqQvlPc3JU3ySNOaoY2wJI
813KGgK4JBo/AbeM8nJ7gdo4Vr9CK87KsRZ5GsDT+53FFETylyFZjO0o5Gx70Iwb
GBmaCfuIYWpm/23lJaR+QckeF0bTVfAKRT8vtVFJZhUhcgyE0EmcftOEsLwP1RIA
i5BGfCU7Ugg0oQVrdWYdzee8kxLz3izMRvdL+DYfYmZpRwqp5TnFBoo3j5M3noT2
3zL6i1U3OIhdMx188wzLdKYdeMu3H8UDjHo9zHy4YBdMarOIF+DlYMQbDtpO+e2P
fJBXoJ13RDcSinZgC2KlQNMIhbDs1WfBmtRQYQZIfKLGK0Vhb12B93y81ROeV4c1
VXpTvVBYZliLSt8euzJUTYSeDZvaud7RkoBvHaF2okcm6jetfPjlJXT5WA0NeWRF
e6F6TaVr1JV+qJjzWLacV8eYDp/mUbNDBNUdVgUMszjxzUWuEt960Nt6csBHvOnK
em9SOmsZX/NV/qcKHx3yK/wAtGSXPKIlUndrUerNkM+Umi8qntJNuPaxKP4NHP1F
vrjwFVbBPZeAORyN5qBA8bDf3zQtDVec4Jgmj+JoWMvybCxZts6aoN26avvN3Yh7
IMcxKdecbiYeNTKfa+qKYZtbN2HbipHQjD26QWrWUnPPKBURj+JioQz5WJ6o6erd
SWso5a+pKNn2x6QhwyC5xSX8ceO5NfsbgK78p9wg+egORIe/JftSCXFypJ5d92nZ
xTKwHxLrF4RARXP3PoZSk5pL9twOLUr/5y80zEnlWvC6n8pYgR5SVkNECWcSsoLo
g/HDzeSYMP0aUDlqKuz41xEnSTABx+tJ5cuiJTwSqo4xbfcRN2UqaGqK0EqCJ1Ss
kkbSry8TBmN6wpLginBQvTpAz/CciOEC5aexpVLf7U4nidlhoDmjmCCNP2QHTf1b
T4Bm4jdEyPYlHoon72qzDNxGvN0Kbxgu7OCVu+S7O744DMAL8Yj0p4jVHBGwbcqE
tv8WsZrnCMkNSzgz6BT5KPLfpEmPcyKEMJz+cs6eg6IywciVbJHW0CM0bZqcBgGM
BFsWoMvp6FuX0EpRWjoUopeFlRuM4x/0SOx9Rt7Q+/jAYptbr7/ZBarT09Dl+/z1
JmgJgzcpdr1h21P4XiVcN7t9i+tOWjF66heJA/igMXK5IUq3Z6AsgSDPImULfy1+
GCvmhKy8YanndzCXEcn8KhEzA5ma0N6Z0CsDFqaWqe2jkUUYEzhzHx98txI/Z93u
ZAa6Zu4JBii43ndUlInN/HXJYIrb6/89mVESEnTg15aJ+q06KJfS/LLlc7ruwozk
3WhCs8zn/q1t63r5rWRNqek8W/uReybo6Q6LL7sUDKZO3X0Jrn20GL//YvYTvc86
Ds0JClpsO6372tOMdgTtVqvDdps22G+gWETqFS8k5XQlZkuB9oEqVExryNs0jHqa
odJWmQlZfczMwOcx3k8HGQBy8pQP0UZuuuYIQGiatgvNqigrd/ihptQuo6+CxlJ/
fStGboHGNQVFqly5iY9A0ThS/tothVGWiZiGP/Ul31CiWxrRGjG6eMeFc8agXaOW
92zrUVbL5QvSOT6ZMHHcWZlPVPdeWr2XDOPh12eTTS9W/x8f0k/ZtURhOwGsmG/1
dJCpM7XCtNH2HUzX0N/9ita78GgSybw+ZJmgx/QYkJ850dyHkXRjMKFtnUe3QJX1
x8CdVu3k6DuUKZ+zMb7peXsBYYg4WDAVkoXwigaR2R5VjpGX2MLkkGpaursdhfqM
zZFv032N35T56RpMQM75qnUC/0AHuo1TvBqJgl1xhfwb05X+aO4plue6hGFsoeG8
cDlQMdT/G6ylYyRfQ4rZdd9qzgHoQIP5OZpcLC7AP/NNTlOybswrcxgpi9N49LWR
xYql4uEz8aRaXc4M50JoMvYap01ggLgy2+Px/f1olAgQ8qWQEGr39txrmTBKa8fq
w/0yG9CrRsuoy+pEtLa/OZIFOEA7UXaaK8rPhThOpFpQVfcGm6Txaf76zXCIPNXj
1PTLTT1qoiXXQPr4szoxpl8i7KQ0KB9Oc+OarN08WEgNnXwt+L4yyUVO2sgQNqMw
hW62RftkwX4/mdBN6HU2kDlrjhmU0zO5BdN3ed3aFkOBXbiwJ/KaRe4YAFrhTCPr
83A+/y1PGLf2HamSfDGdTqokmvdS3AxiBvpFCJ/Wm16qCbSugqxSOlpnjbFytspp
kRZQW+ayyoV2oRehEtOgi6cffX3oQZsNbK7uJKPHcfFnoj7kiYVQXvUS/IP65Bhq
n3fK57BQ0GAm03kmEs/Ti1+apeO5Z8jnD541CRyr115HOdv5jBeUw2bnWj4VokXu
Q+o2TohmVgS0ioYHybjKSK0klixnuauoVVK4IF1lt1Qe2lu0eDFotFytjm/wTlHt
tgK8r7Y9USllHibz+RzER2jlUflwomYYqxqVi38H1p8Lsn6bSzy1iHmDdcShCFSr
+CO3zVMXl5dzDGD7tqYYfQyAE242LzP8ry4CWt8BrDimnZ2sp/wOF45+Drf8ITSf
e7AJrbFSpA9NmcA6Dgk2a2tnvyDK/d2Tw+x22SCSyywORxuLkSZe+Czw+EKqzVHr
XNV7vy2v0APu1DUu5nL5XPCxis5w+OoL8XHVTdwm/oXolc1SXshRP0xcW+l+UN/d
XcO1iUFIIV0DzeIkDonLQH4nINRqFWbNvAheZGZCvES65RkDAaa163uy2zHe35PN
az7kL198rul+fMgJjtuJXqKqRBUwQVw9ZP2VuBIwaBg6Ubd+GrepsaUbI9vXoc2N
Hhr2iDYO47ELxxPNw2iW/H6epI4ZJ29qcQIkeIW0MBXucDRyjpWf0B2rY4plvU+R
39vqntUjKVqq1SV0gRyybQudTpQhLXk+G5mUw3nRgKIac4hihZiV3RBcqnk85Sse
vGlaLuI6CpjmXZGiTzaqCPNwZoIi2ZqD2YY8sJa+4P3p+U7BGi6gZ0dkTaR8HYCY
KRMssYFTVgCBwXIMW7iBPotbVhCye8GdMVkc19OHNHKpr+DYv7jB3GGplkmUa1pq
EWZqFWjkGJC+96O+Gh+i+MVYOcnI6uFaQlHDdIRv7Mc6TPYXRZNJ8NcR6aHKOIai
cZH0Obo7VvW3pc+bLJbAsJxwqR3Tikbpvk9VbKEDbhPA3NY9vKMj++k7FjDMAdw+
/uh1m7Di5XUVlKd9ltsWA5nhZxLpk+FzGFRc+wAtv89NEA997OzgMP9c4W8ueMBZ
JEW5SxNCgeVI0fky7KrfCRPFTm4ZxdFWptW+obGK6o0ov0XwaKU24vd1nqhvLR5w
GcDaGA5O/bGPJmuxCArxB3NrltzZRZwVlgMIXAVyTmNk2KOmTs/F9kvxdwGDIP6r
m1SmqBzzr6+T0alvfW/T7OK1p+SVQp11RM1Lx07cEhzAm30Z+NorgwqxFK4tgVxP
MLdQE83u3Z84E4yt9++NVoUw6RoWKbvFXRpMibjEifsSZkQQ6hAsDKZ6tRnimA5+
lX/kc2NJ8W9cDjpfwSS/6TBsQv9CH3NPOzi6iRif/L/SgBY9DwU1WK+6lBNF2d82
eAxb67P8k+GftqPVdBYvOnNUFMFhBLv4bW5Ibv0rIMcrabCf0YrMA5mgZhuWS87U
v+BYhqKzVnUOoAkS6osQoSpOgB2U330tL9Lusn+dYTdJR8GOgNV8Zn5R4lywsbh8
gDdtFImPWo+tOY/rartOiLbOQD3xs+vxKIbjMJAvOSTHc6tkCsdRttE2NnZgE144
OvmEv+e2lkquCID321GGflnO7VOfb7NWJbd9u8HVn8vSvR1hEgyJkd3ZsLRtPEUR
83KivSmnH/OyjoN2rbHC85ONGNTl3s+fvGkYmEDW+MthhqvDoJ6sBAGDm6DdBB8W
ia5vcQVu0yYJ3qfVfrZeiO9WAWd0ZPZGM3ePlnO0hmWAl1bj6ZtlrzA7nfbC/hpj
/dUa55zYUAxECTyeyIZproeuY2pXgpjXQO81/XlB1xz7KzZtKoNU34qS3jT0EXkI
/XiWDiv+lpcVoI414OHeP4zunkGAAtR+b2IxHnX5WjKC5RV3s1APZvbh8oFUMK4v
CJBHT++J84OnVgI8a//VQX4fPyzOKX9rpF5f6aTBx7a9fzqmM2iAwHRC9n5gvVz0
gLtN9+nIhosR3xC4jCwFHl0GDZqzooaMRzmua+2I0bDvtCxDmLJOtKmLx/ZsiOEi
CbnR0yBh/u603qrukgUGyvq0K9kPYdZj0FZBe+5WRKE9slezafNWZbtM4Xgdwwa5
5o5jKuHY/SKhNUh/PiNWF/tygaJ4Lve9F8xFxirlp7VIfKsOFgwbM5iEOwlWrPxF
+q4q/DpxWONxTmuqJAFMV+w6QLukOrMgqgcGNlml2SLfDSPW3GOt76I5BQvIFnJg
OOmprtdaPfFqq0jK4DSy0ukbHJS9gNfAgKS1Z2vVCFPtrsjWdEQ0V0AjPG6O6umW
34RB6yr5zEJITi80rrDamDX4EA5MQw+L754+afYg9ZvMTaWtPH0EjW6mb8hOYP/8
flItEdxzthQ2IzSMzJTSXnEl0CBpanwtKuGI1cr6Uz7Z63jUNz1NX/cEYNy+/QOv
HBTJJQIXi4tDaTK/aew/SaGUKEo2nNSkxor3rF2IuRpqQJdNn1Kx8BKgSKCnROT6
g7j+q6YUswc9BYqDaBkWPS8/XY2JOtck0wixdAHfpO7Ifzw6OZVhoaZCClmSIzg2
bn+BqbGSbxrtzv6hVFU6w+zQstMzERahnRWfqbMZLxOuR4wURYy/n+Lq66arogmu
V3Og4zDKq0ANj9pqAsmEnGTSkUxwXmIis6c4aMMIuVNkPwaLj3uI9LMjcdGFipWh
3wE02JOhOIW2K+VR9nbac5U2vaxR6pn/JtwjSu1BBWtHT6gDD7EXOrnvfR8Fi0ho
kVY5DZY2l5RgNGA+pwE4i4kSg4TMf8CPL665XRH8aKfqU092WcuS4tn6hSPB2vZZ
EbKXrlzMOWKpR390tx0MsJGh/uNDSLwmKa/Z3RNSHcHon+whYUF49Ca2CaC5pv+B
VCORtkUGY0MaDpTKJCfWA3BkPD9eeukTMnnZe/HGN5RO3qLpRm1yMlTnqJUnszfJ
ptRLvwW7LhquPMVaVrrzj9ckTDDrAuTTsms4AguKs5zymAg+UrG5eQpbOJaGl/y1
6F11c/0Pq1tpzeysqZHop3Ro6RtGfoAeUb7fcrQIRbN9unIX895+C14QPVfYP6dx
2w/JWhgtKvKEFWZJBuI+qC/icqwnxpaoPg3SWvDNx8dBfGvwK1RCQIuP+2a3ivpj
2KE3uxhuFO3900QBq9ICaMkCnfPglwduJkNgnm+aA/7CCyuFgrvk5jXPDqQpNkxb
uZOuhTfzhyawrlRmBAmPhGhcft0w2o6g2eCaTUl+UGvUmzY8ibu1JEgA4KRrwfkm
FKanLCrz6EVk+smdcukc2FtDGuyPIiDgAxBOfBaNbjF7N3ZMx1mVOFnF0GTJHweR
OrdXQt95WDDIuA/Y5qvnlfj5/dZQnykPjcmToUVD7bp+D2BCapI66GwdCwZFLYuJ
E8AmzsfqLSr0LNDW+3QAPvQSQqo5nRi9OtvVWujDBgmx8x+nXEHE9N90J0SCjIL4
4lYVfknop6mPIZTi1uttCFwTy7aSP8fU8Iu7tM1UJUNudHUGXM3XQu9o8foJVwBk
oyXiglnjzmqOyAXzHNmzeGYwDi1iWYOD9+/9STyYJKtYoWhdws1t5dFmgeagPX0S
qVlEotMyHWC3IVh05VTe/MWutpkScWVxMjbmGDVy9cmkVoLyN+bU3JTq/pWj/kPX
uJICGgy5bhBeAEsB/jdxrIhL4d7LpMY3Eu5TNaroyoPU2RgArKdagBlBW5SQv9Qq
wlm/CPgiCdh0yrmAe97nYM/YSpReZSEwWq0Xs4UPfxL+F2bO7LpKQwbDGWbmdqMO
aWOxeHj+F8RkglqOTlk4mOTChwFk7KumIgDe6mWGSlFGfYfUBcHQ/Z/V6kZtn6GC
2fIr13l76ow0mLylqyWKzaThhXzi0gFAr4oEMF4T3apw3DIdqsmPrcCKw5h4Z6Gq
Se+yDJ3GJs5hydC1/56M256tC7PfNL1DfrbO0HCN0SF2F6OBO3wZA63/xoKwMQlQ
xePGtbfnoLEz39OzhdAXVDrVgtFk5NdxDBUNvjEHRdXU4+6/RmiRNqkNiygiYYlB
foYH3lBX5hAR0x+T4DSzVVW82waTUlA8qzdHTpBRcrqsl5BG9V5CK1jpKMlCCpQ8
nY2oFwZ6tzRAd3f8kVmZ0HoHOjcsz5Oyv0eSy93eMF8jfZknepPw9V5AG6y5iPsY
Of26lVnbJuyQ5IJqEuN5yEK3lguxcXaxA++54vrCXQhzoRkdi2nLnkJ1PuNx0ZIt
216C1c8J5fvrD/4vW8Dbk60dHpkL6pmbG0B2crzlTAEtbUrIBJfBNOuM9FtP3bIw
BjfvVcdw0ap3cnc1PyJhIMM5we+t8lR9D+lR9ARPOa5JQb0TexQbq05Od23s5eCZ
xiL00+93ZwklNjYuT+ye8rBJNxJnDwfXCwbsHIzNHXp0YuFrXtYFMY6MW3Y/Ca0j
z8Mh9g0c+PUBJfMBxdrXIqkOKOavFIYmgoCawcA1H/kYCju+QlS62mMgk7lGjFYq
pH0HWxVRgjMCREOJCytTtVzEMZRqejB6tXwv4CNQynTvlZGSWl2izL2i6RoLPZbG
b6by04xhrPAeaJrciEdPUhEaIu6tcxDDqSl/KuS7+Y4i2uuY7xYgNM9gCfSP8jge
Pn7t6cg5kmRmF+4iPjXN0sbufzgJ6o8CYVb4ybeoXP5wDdJb087Oxfxso0K4s3Vj
p9q7EDsufGEPaiTN5OpN+AZCQi7xnu8nXrEhtNuLmYRoO72qimMleWzg9+GhCNkv
9PVJngs/fzPNXRQ9kEvCsjsxBboIGQlJFjNKnhrlbT0l3uICKcN0hSL9D2N2sxlk
1vKhEw89ibFryH8+HfVGRxYFqhQizSe97sPwKngkLUSZqeavCz6M8YUgssTcAuwO
GDeNItHHqz7y9uRyUrEvuJc5jed/HPRmsp3PtaHVRnJPOHDc+Mx5+dY92EcUUb4W
8cFZkW+sqndrLB81LAoILqTHCQoZMfUbBBuiFX/oIxnhvkIjdAO1loKQBJFlAN4T
fwJmGAGpXR9v7B1fkVlQxcAXQDodV5z4/gDzwNRGhkzhVD6nylPmNLx9jDK/6Y8S
/b8Hybnz3mAB9cYJEWvWAlZC5fCD8uBovUF4MByRQiDnXqJWpe2P6uIGQc3BdXUq
Eb0TukmkpqhPX4droJMlCRhZu0qo/bvi2nhTAAKqcZzfHLCKyCX2MD9XkbFukIeh
TVYpQ2diVyXN/2zymZWfDq5ui56Qjv5wIMKb5JBoDN2rUeEEIJe5POeh3gu7GEJ7
4k1pi+pRmvHzoeXPkLQcSThzBXrb+IXGhQUAC1/5knbrwVo/QPvKCalfQznoIybh
AKvFBMHSG5DRvUXTu2PKAYGA72nW1ym6iqOaziitAvrI+bpjPM502dE67N9Xrnu3
bcs8cgTbkLi/zJaIKYgkiZjQZnSDXp05Jl12TSPceGib1sny1xMZSk1pYC06inIL
Dm0W7p1sgG1CmRhshCRJhBkWlBQpKxNTZi/moDL/gZbAmP5p2qsleR0VNMDV2U6O
AiZt3ohgFOJL9Gj4Wb01kbQ8ypkf941HBvvZhTW2AhqRl1fAadhKXOJZPnUi7kuU
dBEZxOPLy8pZVx0wiKxm6jl6/py6PIRzMJh/V5DmA5x810qgQeIIQwk7xUtYKwNC
Vm2FoXrSBDdeaOeK8TY7fa9RkyBCwqrAQmqiG2U+X3Q5nNjB/X0Gey0XOfuyiV64
IzNd5ePGmSR4AjGl9o7RY9vbm+jWljPEV9HJXXvJ6tfbFTMXCOJgFDGwafTMqCoF
0T6hSQnCyYFZn3p+NF1Dj37aITBJbhclgBhfgR5ahH0jllwyhTjYuioxmYo8HwUC
AxE73bfGgo5mQzP+tZ/CYJrMBh2Bnvha7dEXzYuNanF2wLs+7zuRsKTb5iys94pI
cLOWZfrfOsyy5XRGeb2G4JvMHP371sIzu2XgPP9am4dzlhu+HQWcUK9nIFqbM5Fc
eVC+y8HtDYQA5QEh8wIERz7HvwspkP9xG863W3xjXRGO1ODgd14CX+vwdJFL10dt
YXxrZ197jQBRI29iCPJyTxcACSbLNgaHslayFdYv9L91hB2DQXC1FKvLDxEk+sld
1WpmH4/HkViLPEVwQlAUPhYGQf0MRQivNiPWfvDuZACG1FtmISnKauc5NNsvXOsN
8dlzijfKXzgAqLDW/99Oeoc7OLTOtGc00AYPvEZao6gK2uME+zGFa4AecpcBiA07
IUhc6r0p8E1uT7KnLM141hFSAhFwLX42SoM+piE1/PQzB5ZBvEgJ+cno1nD+oYVF
x+Sp++bHsrqShK4Fd7OzXm++rRRTYu7pSNlGQJ87SYiOLHuNJe/NFmCLgN8jAP2B
M3ouhYD+7nlhQPWjGHB3XFU8HdnBBxxXAUnHyfJEY5T18Hj6UFx+jlX2E2gOhIjS
jTtRP9qNrUR1KXCBXVRTE/mesc6AKCRqR/4aE0ABAM+DBeJxwluQOLYCJcpJ+8/u
iRb1qx0dT11881m7bgE0gc7VHeGXFvM2lDh9r8z72K0+eu6E79jLIZYgFk1P70zu
rC4Rl+1hA6GxtYQXLXj8EL48KIFCYqLCbxHT3EXJlZk0NeapCe5I9blypnY8ztPM
BISVtYQePHjqlBDlWELP9qe0/Zwq50+cgRMHQH4hdSLZLMmlk2TwCY65VCPktLa8
OpvIv82raj/epjRZHvqrhU+5nqIFCvtnv9eHeg2wzTpEAjO6K1uGKNnsB/jbDzGl
Z8b9eLHmRMFnxGPTJ2W/CjhrPNh/qVx203/ETo5kbk02bYSuaJ9SgGQQUatzmAzH
bzyLFEj8LFqTo12D1U0u43oXfnCYM70xz4JJCAbRlqr/oxifeCAgvQ3sg81exK3w
mlB3YAIy1f1wSLRvOElB81618zUsN82w4MPBCVdMXpWmKfuy6H+rxWBHsqP2+nYS
gxr2rBhaLjLY4zoydPNC/ofxuS54kEDhpHgLHmXs9HvcnHPEqRduL9ry7NoQe5IP
Mo2nRfbWGRRwF1erbYMyvsr2oP9JyUIfFYxDgSDJ2zI/0IjP+fdH/6oICo9uGVEw
xzc1qCzIvtbdW4PRG2LGH8nBLQYcNXZ64ENcyMUjv8LC44GUCIrA63qB+GFx/ApA
DD/yUgBJ6uiHIrFYqLzlv8Wd3S+SysyL7RXupY/x+jgKJICfyBB0uxLIVm90f21J
v6mkBt4KxUucAygFsoTFuuDq0ttmdUdh88DQPkL1JISjKW1iRZrGofru0+ncmyRC
xnH3llTZHJ/lGYoXoRkmNUNAvzYQfG8uZkBY5MwoCh4nro2mf1jYKAONm18xBRrV
kgcWHB4v4ZWqM2uNz62cKmMUeEKY0si8IXNEhMJNJMHW6eAM0sJEyQqw78OFHdSY
QCoAKzdRYKIpsDMtjI9+5XJWhWZUdpbm7ju/dWP0lT9Z3fdvKtfNYp9O4I9XUo7J
2ZSYrzcyKOHc19vTyx4wK9ooOzaX0DcDiQEbSd205WMx1WE4e1NTdaituOOZe8Po
nZSBeKcZ2lFEL64nN0H6E8PKRaHQ/S+ko4eMst2CUYSMyuLQaVZivV8EyaXVam60
2mSo1mcQhUYn4q0b3pfkxLMSsG1Dl2+wMFLEBjCyxKUXlgmNNS+1rVbA4M03kkLB
0DtfAQAk3bsueXGBopTqxtAjTZ6aNt1f7vSsZrqWZW3Ne4ueMOmrM7p0tuXr8qoQ
NqSUijqbwwRAqykEfyBMB4MV1yVhbD5cStgGcrD0HbvdaMuDvsW3qPZUkQ+V+R1w
GXNIK5+LFjJaUBU3vEAzOXFG4+Q0aEPVoIydV8pkJYXd2Df/Hp7OyzuXi8zz3e+5
i4PExXXSyKiDBycVzz0+aDmA+6Q34GJksEwkapWcG4fwayYpMC/qsX/9utjieX/4
JYF9M7db0plYC7z0bi8j0WtYcaqyJo3wR1Xh5CIDeaYsYYa7qTb886orjPJL1JL3
9SyFiJFI2NsTuajsLObstIU1cJOkKiu3uK4Vdxmq9xr46E17EwXSg/ICZMenlwwa
IQl62s50ikhvCGnOgBNePCa2Twi0Dy5gLZBpeiEo9ZYSNrMKik9+fKuZVvQ9vJJZ
dxEd1rO9uGB8Y9Zt5mstHo4V1XX+FDVk4m3OsKMUYRWsWUonuGoTj+1ShsOyjGLr
sFZ0+avgmGJHqDE7fwtM9i5yu7jvdA3gS1BxegcBD9YJVSFmjiSEFPoLne/wNfoM
AhZ4Flm0WDd57jPXOAXIAV+0HoHDJqizUhODX7tA9yceXLfcemR2U9GxZl0isAS5
gME4x5Jj00KE7ojdYIPGZcoRACuvhTUSc+s+ZbR0Bh2/ECBXdHa01MgihdlA0GTb
U2vmkjkJwDhX2tTnRixM1CqfFykBXVp/SlbDrCLlM2Xf+JWjfgwl2nRRhFG4Xnsc
tojWsrSBF0brY6uDjImVh8JsrvPIDpnQV7xYEYsZ4eAWqtoUMI8C2Se81nbhx54X
w6oD4RMiNKEqse6qz1/xdWzPtR5QEbih0GU2bL/Rpjl7Ka2GsLU/oZlnAFoebdTj
4fqM3y6WwYCcuJ7jYK+3V4oV/yUuhTWNfieSkCes14ELRyBPWppHdAAIWm/awvRp
7MNFOENUQAr/PU6e8YxZnwzldZjbg7An/KUpOfkXExeN8Da5yDnYggK4asuGWEp1
BGTc+yS1Ls3dc9aaeIHdDwwFrpFXdmKQgLCvoidGtaCvygzMMd8qrAEZHz8zcM23
9U8gIFifazfNIphs9f+N12QdtdP9XmIqKyr/2D/RYuTfKzpSlWzIoRKrf8CxB/AK
0qUDQD3GErLXqcZLGrLFcQboRdTg/5CG/AbT9Si+fumBpq9xT1dxfmyJnKONnVh5
k7WWo7TzDZk0UawpOr5NfjwCl/cm5PNYrYDrVggucZUz7WQGCDtCxXq6PzZk9KLd
ZTBLER2kuxpYeCtAmLn7cREjCnweSnn245j1jEGpd/HmLGUCtlFcoHdeGLRDemot
pC1AnvYjm1q4hxXO3a2no+gTK1VamDhSIMyA1WHKPOia0r/I5kSQCzu22F5vhiBC
GZdaGJXpdRJ99O6AWmRsPL+c1UAyO1vY7ni3iDnpJz6RzYJ2+j02FyFnHN/QjOmJ
MyVTL4Bgnrp0oYoOxbGHbSmMpeFzmpDU/K9tbDi9QjPwey7dTyv5tGnhSN9ZJpH6
v0XMuek/XWuNQl1lyqcBZXjlCXDWgQ7O4ybgONFTC6A+bPZw4bzhmi565XmezisL
quqmYRmv7tqix84c35azB3kfHgkygBKzVk5INY4aorQS88Lv65nV+FsE9TvdtH17
NvVv9+40J+zAVmuJQOrt9nYP+vIASrOVZkg3wTNn6WOXUIxaVOISa58ur841Th3A
RPjJCfEXdHTMESa5IJLGIILKorn0+7TQDBhRyMonVGI1o9pTPJ3y56aZF6IEhGju
EhPM91U/62EZFUIB0dhGHShxBrJ2Z6wSYaMR+MROnK5ilgp50sY3H/cx5PkNziQq
Vcr8OwEmgY7aw50gsAcBdH+BT6e094LC2MCSohjQKYLMg9CqgnCfuqLgSmGEmjOE
OM3HR5JBei+rcWdBHe4Crdok8CCuuunG8vRSKsNAQ2kMTOjqSukI+ZqgugG/2q5n
H5Qzr4cXnLxQOS8/0cc6a6AQ7x3pdspYA+CbIRE8RRiJUw+TSDDEmTsNVc95V1OU
bgmGTy0/6vOgoddZ/brpvxb7eO/nSYE9bza8+CzNwVCgkGrFYo3xk7Z5il2TiCWl
ZkX/q7FD1CXQRJsaIYSMIITBzELmaci+36Vo3npp6d2KL/3YJ9LhUXBqXZKq5YLz
R1jzWt/8CbirlhuIVYrB8uXpwj71bbpPsoAybOykL4ySRh5zM09bEA44gF0h4cC6
ME2FmZtc1saazZ1cllWy9fR4egGjdEX1LaN431pojwEdkTxf1PLFW3Icv8UV0FxB
pzTOORC49asA28f7QNcjBlujrFssvIx8/eNzTOBv4h4I4ji+4Y/yt6DWfBKO8mex
dEzKnMEjfdoRD/KNDPM8RXyLtXyFwYbgJyhgw9fYD/73e4fiC58y3eeSKH6PHr5E
wIrIbBI13p8/vWi+5vsC5oB8+MgLIPUuKwyivLqqv96pHtY1znT4gEHoUOOtlB5N
VswAalwz7hY98cvohrjCLXrH8dxPdBtNoU5D3OVxoHdZOtnD9VzyF1DyXtG+zCSa
v4UiZTxLgKuyW78QdBwpyco71NOuOOlSpVg+UMZ2Hq2IsUl7nez5dsSh+zrjHUnv
4cTj9uwvQ90QSTyEkfEBDTPeBLlculDaIlDk+HLKlWjn79Hvkuq5pynQrN5scEY7
qFHG9hqvBx6uSZibGgewBBXXGnHpcpLDluHLqiSPyUGWTTnyUmuLt84c6kMEWQq9
9+vUf+0knMJpf44ji/qHRHrPUeF3/t8hCN9T1s141gJ6+/SUmtp+dghzbtHTenyG
QN1amxlWNJlzcYlgmdqlpLlPDeqLfl4rQsM1SksK3qEkhiZwGn423oHHQF97VLKQ
rVXFUOcorDu9Q50NzLQUcrOKP9I1LtAP+TNMmqqhOd1cx+J9K76/ak4f2PXoglce
zt1G1Uq59fSaqqvaAcwoWGT+Av3+L3iPCUJ2Pz9OvbLPuf19EMxqu83CreYltLvw
olN9ha4fivkaTsc4oOjssIgr/YzumsnSMYKO8gnx4Zhle55uYZzrOzauZq6dHr4c
WH/CNzLIZy6AXx+6KRlfkCzyUie0Opg0+k2hon4FQQ1V544x2HhG5L1BEMvAUd7B
sTYm/CLlVX7MObMzJUzL4wO1yx4zpd4F4qlAO4xEWufo3fQwFLm/ZnciyjhtPNYX
FenIG5Q9/i1OKiZOtCqe1euQM7Qpay/39OBRNE82rEQcXp8dWJIBJFGEIBwHb7Ip
EV8o3oDXg3Eh/Z/rM4RssjCCTy4ROICyhNbCklUnY4zhwhzYA4b+owc06Rot+wev
jlqbUB9FS6dw9ftg/KpRADq4qLeMwdZJk9yvMkmVlYWEkBvE+x6WPSC+k6iJcWDA
XavKCoJEJZGiIGuOavcFNQLT1oem/GLtJWcr+TG+BkiHOj/03rJrKD9odn21FxxI
lewZsyqbxQ5hK9fVtysHhAqFDrjxgSE00RVb2zpPfk9yH3nf/UNACVQV8R9RHvQw
qh81AeHPuWVxSNGMWOF0pa2na1F43jg/ujp18O1UuEXKOHEW84JSePH/J8awUiTz
f7z91ruIyJQwVU2AtYYRN5wS6nNWeoCdFeBLuscu7zPFivXZkFL4cuikg0S9hHGr
xDGfGvrqUUc54NjpJWwkhHh0ph25iX1/s/HhyF2LumRF22OSuROOvjMm1rgZSmjZ
bO5eiSeDhmCzSAWun5FoA4miWZ3SS7PfRLaSOUrpQ7Xb+02S/t80shCwQ0AG2ivM
luAPqPHV9MMl3YMVYhStgFSgEuRoWhD5V15GdHPz0hI4yBnGEazMoJ6FjgBHcrut
Ed3zlZTcflM1oHq89KkkJxLTNOnlntv0asc+nMQvRVBS5P/9ICl83oIDO3x8+nXZ
cpUIt+Rmx1WbMKTjYiZ9BEswZRLw3/eWy77Sztx3I14Fnjwk6wENj6m3a5SQcm5q
fy9NDvMhVroNjPs/RwGBKMjrpM78nEdbM+uAv0z1ig0AE9YBp+YLFPNxiNWpniCU
cyiTA0r+BHOmnvpeLqYfMJYWNTyd4QT7JvhZs5JuMlIH0TcMsSq6KU1O/t+jm/K0
cSu4eigwq2Ro8YnRl0IUVzp1hmNgWQ9RcGxatsn9I0Cl78F66hyBVokylmmbpOIF
CJ3Di1jNhQNWEZ53P+mvdDb2yScOXmu+FOT5LeeXHjkfRArSylaEjzf9B7TPltf5
ZMcxy5rbvTccWTJt7vXE8CFUAENbJ1MKGDguyD8fqRLqNZLR74BUZQYFz3GtCsLQ
GPjf+bYxlCEL1jEJuFZ95OzNQlWmMnnL6sWEIGogFWGHpC5ZnhjqFUXNAyuSSOV2
D98ffYpRRT6FnXLr0ktV3eLaZwR7UovZfc4LQ8KB0dOUJFKeTYp2/Gm/yY9Duq00
zHSI4lMZohxua7IcrwxXdac6KspkUU3qATZUduWxsDjrOZ4DSNGD9NqSJZhjMJkd
F5Fej2Kl+ZnuhrSLuPT7jzJtuMszJGBYsvuuwcxMvmB1mQIrem+4fr2lbGKFvZd4
PpFzA7rZvxfbdHi79UlX8cFwOn5enQdnywiNcOLDGDepraQZxlMlvpdFjWT6666j
/OZcPhfsZzVgICsRxSmJhX8BVVYhaEeyg2F12UcKPUOmEB10V8mpgsGMcvy5onIh
iT9auoZ9jnVW3cp4vhCZbI27YANd9P1wztmRFN9DLyNfRkyyOlpDGoUvMYbQ7186
bX35TQUMWpINNJm20H4LmSYAp0Sab6nRuGqfcsETIEYGo9DYYwIAnOuFGcofzhZP
PAxsdNoioGWno5t1hTL5L8OEYWTM455VMWh/0XKsbgY5E34HPOalvygtZeROc64m
gzoxMd5/T7rcZa4E8jjeIuNl8zeWGbc4mCBoxfhOmKgcmoAOMfFiWBYqQEmAop/1
OLc9xjOYpuNNWZU/wGOEUptk8F4notQRDnZ5qwwo916K4p8wbQ4uPT68zw5xcFDP
dvG3BU9B7aXB31MeMmJJQQCymXWIc9/w7/r5gIrGk/KThg7ne0CErksP0TIJpX/L
IgDQ3TmNAhp3RSAqOEW+tvPBjXJ3mZe4FmdKFN8RWfMWr/2tUUj8Uut36uMjGxgH
nv/xRGKwAqf85CSVnZEQTDD4+0K8OlVUbd7Gr/eVsdLxf/s974YixR89V2Sze5L5
4wit8RV5rWAY34LeW44abQ98Y+Nd7EEFp/8DkH5BTpEhdKUhOEioGScx/JPaZqfD
bQF2RxNlR+uNB6dRDJgqJ1hUmxYg3Mu/OfmaMXReDv1FX0rVcL1n/C3OX0oyTxFb
k8BA0TFMTNP0kY5e2xsMg+7S3HG8gZc3yYJWr16XoER6oQu1T80vzzNKNAFBTEvq
mv2krNtwQlUfJ4p8Ctqz3J9241RFrQh7R/vlAygwX6bOG8Lco6y4mkSCM0hGbl+m
VtR+JFww9O6Sg+lhvUwwpKz1+EyoQ/OLHl2s23J0ioAzWkB3CJqT2/mqSgAn7VK9
sTydbGjz6ZWKfBrbbjARrYkJ9JSxlUMZD/xN43Zfmj3jFJ50zm8yaKfGZvHvwQVq
zpKKsSl8ybkYrQbnAuoL0VrxgzatrssmCFlM9AC0+4gRVT4zytyNA19YLH+YGEtR
dkLisVGgvI14neyT27C7/OeR2atM90oXtJzdHpwluwAkilhFHhqOQBJ18+U6Zxbu
I9ncKO7SoHCPeL0Y95OoTYAggpebOhnaC62+t9L54DTlCbE13NX5XEzczQU6YRJA
SH2mYdIiskTw6PJekLrkBHopMyPFaxj6doXVUqsVM0OYLjMp0ghttbWrwazgymKA
NUJ0GQaQH/6vx4EQ21FB/Q0YziWEzajvVb3zz7aOCyCabMam75vTqEj9z1OwnYFx
Tx7f9/MKe4PeRkMHLwe7OSL7QNBkuDBgXik4su2TL43URnGVnTSRSHbBxiXM0Tvv
QJ/bXFFjRkIBUqGFaIYHrMAqsXB62wXud8FPp3ilAOU9x6mF0mWFRH+EhYWYB8ed
q5SRRwK+1ksVnstWnhgmObsPMMCEIbK2XAitsnDIG2H7AVwi8QIxw1rH/L9+bKJR
Rmb4XZFk07VJ50qF7ZExJXimwT0r+OxUvmq8cHr5SEV/w9yNKyVJqafvmP0V7gdP
ZdNtf/PLJc/h69Mayxy+T3+UgKNMSHnfjvserppTm03ZEU5Tyjx2sxmRtPndXHWo
Ch5V7c5ClQkMmgjdiW87ICVAgo+Nrl4IgbWFTYT0oX0JU6PQiXgoaUkuoWZEfBmV
4plkqU5t9bADf3I3N5p/DSQXOuB0tLWA37FAJx+EKCdf6tv6kSqEdVftSUwBugBO
OZurzVJMv6Y0ja/LcLfQ5CCApJHh8vDBQcIYh3Mm63fHtLlAsO16pf8DedTAKy6F
qXyHsrCO7GurAn3meEr5/T2Wxs9//oVbmineEF8SX4CriOnRzephPl6Q2b5/XNgW
DtjMnC5vybwxOWG5yLhGAI+S3qe55UMIu0NsEO696vydnnp0/BNgeW5k7rvyGO3x
XK4rnYGLpg/V0BDv6X7WzpE7OushG/guBNGxh0cnXwLtbZVPh31dwp1SD6l5kmIb
XIgdLArzZXT4rUQb4DtfFzm+RoqOzjYmjTdM9gWDUYKHS2q4BZUjbF7ZXHRVJOfM
ZJh2xlcergTucsk8yP1OIz3VG1phqbttQiFtQhFGHJSsF++3rQUu53GYLb3w9jew
n5eZeKnyyiAVzP2tABpt6s7/yHkgjZ62zsiYxe5mmd0+FAdnVO/qxfwVfE/lOJo6
4g8xxaIclrcKDVIcygS1VMpMfrghUVRo6GrDqHgRff/O2cu+yATUvPzbjGwTJ7sx
IFSZp5Y2zhs56oWFhTQPfvd+E7Ltf0EaYs4+Cc+7mibZboWQqj3DlplBdCvfAjQ7
W07C+ezURRZnXP9auFP4AlZ45+GZ+qsc4RA4XgM9nLCfLiJ7ho6lXbnjq3j89Ozx
ikzx/bQyjwWtyv6xuSpCPo+jGgV+2QE8l/v3TZdCh/JOunWSMEam6xBye0oUDr8R
qCrjGqpH4gjynmvtNNmQ5YnMzNPNCTA8PS0/o7jmzxjjo/oPeUQ9sfunw79l62Bb
uGrJ8Ox14Me52t2oj+0LEaQBHpuVpd2nmg/tUAciip+VuhVMQEVadrugryjPpvWg
pYuiSr1ujfnT7+p1lBFFjs+UlHmYBuGE664akhMCjmZJHMab2dZgBMuqezff7NYM
BYfiRoXFyYpb/IMv1euMqnw3yGdLZMlKUkgvez/NEGuRM9LkFP0ZPT6p3T92l+5x
u5dASAy+jONTwfWhd242shIJTOgepKSUg7CzGZC+MDfXnUPR3O5LAJJevFaRy/xh
XTMMBTsjdelDkXekVJkMlAQGtbSkLw/gcsBcclYfFihnRY95OgxCBuJVeIY1R5mw
mNcBMt4/RQr5hIuthC5g6lLk+khdzLQd5NfvDnM2D7LsnRAf+xQ4p8U+0vTl3TB6
TnNeiGucBaj9tAYl48ShMFngivs0/0XBLIAi/xKP9IOJQUCIO3FqLV4JmJGqqF87
vfkzp07t/79fDf8BSXQysZjB6bbuORNkpEw0+R6hrj4M31I64YpVJvLL1QWOWFAd
vGW9TLmoZP2QPKWq4IHD6e1K4iG9/3Zae/SIh25mgvHu7p5asmHt44qGfud1K4tS
37d3WmG17Mz0RzrJjiPv1l8vS9+4Gur4QbjTJtRfTHDvFVZgLi9GbF1+E6aI1sVn
cEHLiFca+Em4kVl3JqPZC6TPtFJTISFnAmMO4jqDeRILm6d5rYgob6r8sU2HPGhO
GRfTONiKyUnx4UIc7rBvnWnXjioDzReCtpfbChlna/4h1RWZhuEMcIzL7nCj7TY/
UXZt7dwW5zliwENnVSc5u5+mUW1W/+gArxlDbnj6rXIX3+2u8jw/G6ZRbOzTc1z8
PISBVxaegWngAtxXPwB9Xjz+U+5NXawurhzzlSf1UGU7hMuqa4lEWdmxOOZRmwkD
qSNEXd1gkEd/5hSUuKnX4LRDfYQ8FAuIXUSEzXeOwUmX2V8mxHpLUs0JXb2HPVP1
LFL2qCUF20AvMxd74qYLTwMgZ+IqeaFGgaluteTGi95GeGJzrhgnkVYoblXF2eAw
1iVBeRcZBcwqv46xIj2Pn6UsDpCj0yDsQuVObquVVYuC5dQH5od/iOocOrn4herq
QRDw4DbRMXifNkzSmRy4MMalqNGQJPX/FF+aQ/+vVdbmYJUf0hBkX4hrigbYu/wZ
+4p9ukh9IVndTlzH2SsQS9KqtNGMd7PKkgojrJYufn6jPxr6HUyr8jLOYuVwylWQ
5XpeYNGlgDClqeU8kvIRAlJ5S541VeJfAmwViSql0cyWyu+Sh+rATPhkfS2a/tZN
x1aJj6/ayE/WotzWVeFHEST5nL9Zmlql8PxzrrJOZEZW7nA+eRTWBMji78thCKYD
a4XNiFzR7+C0p0ohS9FJrTSQaX+v2VycBWtaXLVdZovSmn/2XjtI47UPjPFPCsxe
AWAKk7FWD73FVSclStiLnBMlUemPn2NISPnQ3YuqqfhzhiomjbH64pFCvF23ei6I
aFl8Z8J3ODgF1hMlG60zaPAYrhijSXK44wRbVRsLoMJuyV5t4Rh4qxOlInzc3AOl
TpqlboWEFtay3UIueQShkIEAs0TE4UIERyjh2DehnS1hFFbSoObC1jv/VftJ3p7k
xj1/nTP6WBG41oku1jiFya9LeLy5QY0jwVThuQr9x5KaTrosnd3xdg+m5b51Toms
yZEphEGFgO9toKysjF3u0JcPMZsvjBVA9HUsZAemvV2NeVZLN7+oRHmgU9gQe5b2
A2/oeHdK4gHu5htdXVWGV6jqjXQCewgtE+uBlYdL5fJXRUADZryXXQdTYizNsa3t
2tGZLrWJ8BN86lPSVpwkyup35Y/bBkZsISYMJovfZpXAo5RVAz58XUW3aUQVm6vd
YS8iZl3otPnh9ysmWrDAuKA/Ot4ka+Qlgm9U51CDqmPiQJBEJS51iEf8SR7ozosP
wUfF297Zlh9UWyYRbjh4U5Kikyguk5+J5Z4GxGDvEgFTgyS0HADCobgAtp+zXigb
cHmeTWDvQbiIUZdAiPZya/+O/vmttCmZrD2eRl73gkwZKAStZONTxgGMIputN2M0
t1d+VIIlXUuZJFJtXr/TmM0aQUy9Fk0YyLAABFUwyy/sQsY6vF7LrMXwB87hiR4Q
WcBsUe+G24pzieH6fDFNuiKthEqkYyvmMthy7PNL+WqVoc1BL9XTfzl5ySQ1lTnu
+YUo9sLfyCugo2o0w09vzeVz2k59aIxPVMdCJxSECIdsXXY56TlSAwqp1HanWh89
6peLGJNGzFPln5mED2T0GCTA0Qw2xTDLt7XJUK9bM3ks/xVGQo9C2Dd+HbJ3DQ3S
NDKIJsxd/mAdJp23LCaiX2jH9VT4dBNvpdCVzGhGtMN/G0UlBuRJ1KGPRVle2FmL
kY/K1z9k21cdqd9qnFoSXLrk8DCTUl2Uo7Fhhb0+HDFWfCQ2PVDwge5nED2ZUlvL
WmuMKOVEY+fB17FsAnSxFs9hpn+pha8oernstn34eGY9FtxYKMGPTgpF3ExeWjtd
Zqg1eOJUB4YfSCHFM/IrsE7IPOwAO6uaUul2VrKwEET0/1pJ/bSakWS/OR67L0bY
ebXlY9/ltcJBqN7G7s338JalJ/MybRamIz7BNF0ZrTj1k5BnYEpObnJ/382N39RC
VxEtsnep6/L//k99lMkj2dGNwZ7eu4yxSFdrnx5ShYw/EG0zCXYGsX24wwlt+tFO
o9h84uz4DoeV/RbWR4UdACtx0lvFV1nq8PpStgp5YAXkYAzhC+C+VeNbFFPoT1gp
oCFy3NuzjVU/8xF/ySqhtZKMVfZXux/CR+0NI9q+WSxldeHzaAkJoMF7a4GZot2t
/1OGFnkasx/xfUUQ9HIeq0tFMP91NuWDGqP2l30sGRgVUYzdfhIP8VXfWzKstbTU
vWi62mTh8tR90bAzfHjbCKmdsXIxTA9zUCPi/H7tSFcANN6teGObt3txDd1jK8Nd
wccH7kkZ6sMIFADhGElcU7pmpGGKMU+4bLUGxCDmCpDwtteUOO7dXSTSAFsYLv7y
WBwv8G4R2MK+lorTBAnOoadPsPcc3mU8rUuDLg8JCO+YsTRNWZMtpxocvcu0GBqo
9Zq04qgMKrB65LH9tTxhpfKl84gE8BPT7Va1dC5rnxHYSNjZ+HOOIi02j7Bd17as
r++9UNfoLLImqMv/jU9yIwcJa3hv4KoeoxMk4/Na40/Auyrkvmp7jgmjGrTMiWU0
jpGm0B+rlNVR/RksIvI37Jpn11+gntN0/cut7W8t9n2ID9J/lXm6kZGkhXQlWzXW
4CGQikRjMWWq8KWX4vWDkY7KWudkNqJcXirdoQCbchd+8LZXsWPQ/O/bgjXappXI
A6y1PEoo2KFOB2IMKWtEam480KcaA6g/6ZWwDH9eNHzhphHTb6paOckIiCyx+cM3
VVaJpKralliFKXTAvuBzI5tNTbdkSFEi+YDxUK7CoD5ftgLZiNClmxClUL/jzjj0
eDwiSSKa/JTpZ81Pgv83mSRIBzdvpr1zxV6wzwoqh3bOykM5SrRUTxcpO0XXRpYU
7mS1wUkLN0/98Izg/euEs93ZLHVxdzcXYjQYPBkdjSH/z/tfJxAUXHbseoHxgitu
QDCADm2RW72g+QXdnjav1ZyQvIsgzuth/QFWk+4dbw10zY6+9kf2XSNeacH81yeH
QKpZIdO0J/eiSBdj0KINzZC0V+KOCeZIKiQVJLWtlREIY7DnRelMu8owrExpHrXw
va+AQyfmuXcrtPuiq7CLEmqt853bl0jQTCgKenoWlzkv3OZWsCSRNQyDamRJcYMT
nswABNg5kQ0IQpzy9tOg5ZjYChdMDUfEuZcOTbq7vNqaDVY5nMcoy8h/CjWi088G
Xs/zIwEqLmmoLCgkmz5SFq1iWW743S5YHy806WPCNc5QOE/DUstVccwO9ECDryQm
vEBdw2QTOm1X8gXDltNqIczIVew0+ya7Igt5dcNVt3KdV5yijM4HnunyJl6veAb+
T1L5Gm5hawiOYLo4iogAwEbX5mUa0Wp/nFIDVgBT55AazOuP+wEIfZPCR6ZI3lQ4
WGJl6rK4OpBlkWIRtDri5bUul0fb4dDYq6XB12gYKlpT50pS4ztIVGQZrbZ8HAsY
AnVYXLE35YNZV1K65N190D/deVxZoHhrYWsex2Bs5j/+dBsQ4SpzXUQpJf+BBVQp
aFe4H0KAA3ns4tVR8VGVSw1XdsjqWrDIUaM3ZWJwshiTZSRfmngoe9I0U+OM2FVu
Z3/7LaKeN+eop58/TulykOSsnuRtnxUhiCVxsxNJydJOyVxhQx1FEquE/5c2hXdA
2Jmv0tLbX6UE7a0btav84neRUUnQ7tAkXmHWNKL4XtNF/2gX/UDzhhH/Qi7pM5/6
cIgzRQKyKF/laPH+Z1+2so/2C0/PdQKq9L52AeOatN67XJ1zlebhesO6XEeovzcz
nz6/38D1pHFRJDFzdnnce+wxO5NMYiNEPVhAbaC5psBlfCLNihNlZIZ4p+tcO8qZ
De46t3iwq/2Lirv6YR84yj4oxHgVZJrRpcl92CZZC/slxBEn3+Ds8+xyrqrSTiz1
ywV+LPMbtCfan3UN44v3MYY6ItT0YtJ1Cn1o892IcGNZ4laMwyZxqAgTU0nEBo5J
oTpWX5vbAV6yuK4IvnbhzA2L9t4VpX/PzTeR06kWkSPGZ56MVpzdHhCwChMvAxgS
jI3ulCd96zN17TeohJE4UyVQCYaqrExfMnftoWbvvJvHYkfXBGBrW0Zy0oWGap7E
hn5znIJPbLxfOHN2onlrbzD6mftwp/Qh9f6VFigyWIrI89iX2+cUuc6UnCUAV7Hs
9+Dpd0veZ4jV2H8Pk5UxfYRoJhiK1HJvMj7CG0z3yXMkIVG19m80JHo6k1aW6LH+
Xnw7RZQq4+LoGfNmji+ijJaczcAgiO/p+kbSAP4TW4yzUam1Rwa4rWX4ZridIIvB
Q1vmcM0AE3j2+o1MPjpDoiXwSDWXp9Z8DbQNgTZrXkkavp3NxNoJB0ByIL2dqwkO
nxlvDimYoUmC1amzrykW41LxCTXkodZEECvVDRAGbFAS2iycL73wGyoAYQMSq9Y+
jdyJ3F/KuzLOxbu+L3jSLTdEmMUwrEGTEIEfH/msIe+gXNZdjN772H9SVG1Cy7/4
Ya/vdnY2ST8pZgyBnfHaEfz5T4Ws1LvgRC1HROrcvJ7I7x/d6EUaOjjxsB8woE7l
wOM5FWKhUta/YhwsULuAEDW5FhYvIsGsfzX5rnouNt77B+7a4RY3hDt5OHiPVqBw
Bn5ZGPjVmFADIpUgDREyLoC7/BM4y8uOYQRWhjCWp2iMEWd18rY/QHoQy615bY/p
1IDI8OfWZAsfvpFdagJdXs2kmrBdxvBQJagA0No+nP6byXv2x4rbJ3knDRP+Pio8
zwD0jszorOqQo3ObXO7Ot9FPrp6DnGJdywju9Xu7X+yQbGXyzJFCtvexVyaHTTxe
p6TiQKS9dj1iHpHXYFlxiyVo5jiEy8isowJnIgW9wGe3K2SWWWZMop4pxElJBv6/
Zvh7+dqOvTo1bT1W8tRzxV9GkCP6o6XNfey072l9aiC4rnwKSyR3R0zVap9s/g33
HXonG7DzdgCVmED0/+V/w/pmN9fPBL2KzAoCgNg9+1aIGkA4qfcDanWf3wrTHviM
Bd2WRNIgJAy9jBp8t18V+LpARIPKI/s65dtjyibHeyPFpm+vkMAEvqjS7wp9P5Fw
Kw7tbrFPoQe0dSDUZmyMNWKLuLTlcijXCzTTnP+TRuIFSy73kfiNXL1QKVu4lP3I
w/qkOXspj+igxPu9qgaMcJy86AylcfwveFoAQuZA6UY/32RwziYJ9o+0VmVrFbWi
E5P01eXdXPbVXSuFCfaO7dqxrv9abbA4u+FdFb3Nc/JOPtcg0nhfLn3IkpsWVkP8
vTvNqzoVX+U42OVigJJHvu9O1smCYoHUn+dRGj1k3MV51UmIxiM1J5fe2b8murcI
kx2ik4umT0ZIoh2tPu0vsJPmWPvWlOwOOQt3kSEVUOhwkneXI5iRs/gcMp97fFR7
4zdrJuaieX/r3i+QerNv/A6qKkx6nraJJ7xirAgWSKpjyNtaX2YFUOxLFUJaTgmm
08W3fHTqPyBX3zuMFT6W4fGaBT7Ib3oax2EkVM1xkbNr4VHX1spIQhDlwSf4qpHT
lqwgNDvThMTnsg6Gw+U4JnQEno3/S4tbdB73sMTHXrt3DUCcp1v+6PspujMVRx0K
9Wdr95Hb0QuPV9scbvsm604Yf4QJRG7Q1P09QIwq8ku5quEppOAIlRH8UJWMHXQc
C86i40HmvHyambZ2C25mWfBbWCFwCyAwQVBXzvw8CjraCmWTw2aPYBjkMTv+DlUn
qwUxnXGnr2sZ2gvAqozOGjDR4XlmItlgyCHAjo2BzvLrwdIyARuLVItr/GKMYGdo
Ny/8BHQPx4kmfHM9bD9LdC0KlVXmWx6AgF48gkmG9lETDm5XxkvxCK+JV6dCjoZf
pgizzjGGw7EBICpDjg2c9e1jGlRPjLeflooACs+V1hhR/kK4a0odzTQUG0titORA
yiwv2JEHFd3zcfLAgVx+kKRFjafd+ZcwuaR79W07jAqbfthtd/gIFy6tSwCKphHO
bi04JFEJ096QvxkErZgIlynskbYUaG/lNVTjcMV6biZax2nzwX5EzGtUmBZs6nZ1
3YhI0wUjX5H3CgqutZH9e9AoDvnH5PiKjFwT/nKZ7bjTPPf0VgNwyPdLKieS3mV5
pZTkVA1FlZJQ2Suh7DGPnJu15RFXEJrY/m5Xuy+0Enz421k0YP1ou4n55a8PDJPT
0IpuB+GyVLyrIYY44sf4RJeCD+LULbiC4pXMz6n11pVxFmAQIvvcwvFN980fvWoc
z//WPZWqFdOuC+8ScroO0JUWWq3ibj0YGwfChVZZZjw49omSqOraRAKgt7YBI+rN
P/ZKvjmFhoVcQFDjBpaMqW29d0ebLnpLbiLnFXS1jlCLU+KlWzxSgXpVfjfXooUm
MPyNco5GGIUg6MRPYwjitijtIvys2lWSYmxFWLsto5JXEC2wvd6Queww4tSfnGDm
xo0HX/CtWFUIlLVIv/ZJNtVCwth/1lTu2iQD7q25s4OS2jzK90N6fYoLEh+2+id4
VJnzz6Z3XQOzanL7v1dcOcjunmWN6Irhq8Hnyxsnc4avrdBhVPsGPb/8bjdaK8YH
DqWRLBh41p/whEz1F8WKhAF9AQ/XaQ2G5y6AjrhMHGqy57mF7P1VQxPOe3JPVsRs
fqyhYjJUMAxemP1HNOXLy54yhsu//O7rdOElZUla2RWdB0sAqCUrYJ1nkjTgsG9q
DnRthusVPoGO1VU/KXLUIhHxCrLk/0khelYD//w9JCTd7h2lyh80Cb8seKhxbZBQ
Wb/Qd+KGr4Ihjw27huvrk/0iSqJQa/V2UJ86UsEBmP05MIyWahS4PLlWlgCtXPHE
HqPh3LlJvbg/rQ0CWdxJnZPzN7r7ZlnzVdiGsZ44FWLRl3sgBBawam/CN5Oswfvm
DnS1jBbWK7DPwZ6JM+lVez0Q2bybl4PF2VnITX2P5f283WpRB6E9CT4bRGi1zekV
ciyQaloX6fXe8vSUorLehq8LCna/EpO6LKqt/jQrnVwuNrCkhN/ddqK79M2zmaza
ZcKU0CFYLrEa2EyvB7gD7jMKkN1s/vANJD51kXGFTNIft33NfLXVwXMSiSZJk+gf
+jVfpYamxyuLJ+7X3DoS90kuSpF0S57KsWDv4EnlmoAnzfLPpzF5PPJV6EcPl8QI
80IxKMie/pU+aSGekutATZfiJ9Gy1imkVhO45qaPxKi31dxWhbLBazUkIhfonwbB
vScgiloPX6UtB9mqthfBi+ah5fiQ84cmgNSUcBJmyr9cN7bm/sWLj6GeSOrALKWv
WDb2ORD9KQTN9LV4lXA7WbOVzmrPgA2Sv7KK7ONTgJwgQvBPTR8YU7E+V0tJi2dW
BKEySYubGmmq/jP4nHd1cSMBoeHBPb1Vpq6nOAPgTpd+28Um6xhki2ZUj9tmHlHA
DSZFKEL/i6xkPCYN5geTh3mA379MQjnuHaEP1bwnFRFwlfXzHHJPFcCuwJioXox8
NpPUFFa3yA5idOoLldDjk4/lZWLjq0/Q1oEz/L/pmIzN+3y5VHxFitrz3kdJkbaG
13Os1ZpW2GAqSyFYnh6Iooh5Kb53y8NysRuPjStLtG9BhRIUK8u8dCMsCaDHGNDm
caYlKHqC4SNay04lI9QvpVEmzh3hi6P/1v+8eFdx7i0ZwQmyXdnCR4fl9hih3oMS
cBF6ai3v4C50P8xUR4ecdkV+OMu2h2YQ0s1EGjZWYMnji5EkyThC+Unew7QQZbPU
JdtougR2rsBbK49oTwggNUJAJ0xGaGiMVKneEorNIOt9GebKPY95jwdiJZDTKc3R
bkgTUMNEyXaHqyNymCUKG7o01LTzOk5f3iQ4m3kUAoDY2tyBeuMk5VrX0A34QSz2
AorHZtHLD2zDkrfxR63aHda9z1x6v1jrdDLzkHKz4gX6ZkOXUqeJngvXeNi93tHS
GrNOPN9bhn8bGUKkVUQPGKlCMXtYAXK906Zg0uk9+9YMrBa/3D2OnS887te2tfih
lXFmF5bLnUbyDxoXxQJkNYeOCUwPhYCOqUWCiMN/moLW9ozY1ijP1eH1+RmhFTc0
VyruD82DoWdh0fvnAFQ5BOtcgkNkshFrYmcpobCpyDyB28VTs3sIO67wWkihT7NN
YREojxNguXdVo9pJ7VkVx+8mIyULv+8CYviyhx2C7OxRH+Nazg+22+Vz3X2H8GPM
H4V2B84GD734TbK/wWzLxzUEeAKQR0bZESC6gf217ffJ0dTbhvQVlZ1vNE/GMMDZ
j1UeFwZhvvykLIFBgrLuKSlelyOeZvEsB9gcfsK8aZpODYLXbX65jWDfoXtpBsIx
qa+G6R+XX/MWNQ3RkliV4BO+9LiOPr2MOHMA2WYV+cDea6ImoCVMoXbnpXhCxah0
D50E7apYPsLSBBazISywprtVLIEY7iYCjzWKDp/8D21SNdBFFDkpyyBqIaqGWpmR
SFbgW97aDUTH0Xo0EiP1c7O/zzDmQ4Vo5Ilv5HprCK2AVZTeiU9EXGwDyn4F1zoG
+B8E6R50hLZb/i9oWQHHbZ0LVxuaQMBxEbgispEAymcWEB6wYoAohhJoloPmmifq
i9GButsxt8MTp5IRJ21A1R3HIUItekc88By9vLpWHufUKiAjfPhaj2nsirKnJFBm
sB7gzq7b+aBNL29NEJkfLpk7RDkqghNT0fm3lSQ9vqIzQwFn6/Am5hO/jnTCvB4E
kMeTJHJ9i7+I8AoV//cx3WUb2g3DLYxCeljjKdnwStOuBscc3acgBpx0PEOWiGD+
BGrVsxaXFt1WX7dgAiq0gFnNjDfZRimufjMKNQeayN/OA1mPJcjO5PKlj0fXL26d
Cm4jynnJTSwrJsSeDmo3H90UJ91LyAJQ3l03jcywkFHqszLIcBljai+QE4S1Ubto
TkrPGyWqCjnE2yrZOE4shiSL5VbDzDYYwwDRz0Ppfq73XcS+A4jMW0kerrUf7J7n
EU6nij3jS/VoLRJoaOJQ3Gow6YirXtnDS8Ahtea6+0LEJ4RN2uPOkyUIAaweKKyh
LCgwQrJLqNXoZdaUbjvOO4HdJQwFCGRbC0cfsW73VdXtacTGV40eaneGlhk5Y5sT
6ueStK1SgADbYM2NxNAEWuXUVH+OceJwIaEFhuFOr8746X80e7g+1PHdmNTVTeUm
Pyg7afMO24Mmgarzq0CZgT0dd1/JU6ofHi8/k/6mWVdX5ov3IlVOgKjhWGNI/TQW
SgU3b4cqZg6+e6BvYGwsard07FxRim7HoVsEN1i9ELyq5mAKg+qj/J0H8Ie7q2a8
2NiO2RuQSwMyFJS7C91hxI5LJoDVmAepm1HXomkmhtE1w1zFTvR31v1rCl+hDL4I
YVYjhAgQr2Q7biA/kVBdIj4JN1+PmLPisON3WAejF9hapq88IpjBnpCimcekaSe8
jz0podWRt+sKVYDojCRCCHfLuFD4qdLLi+GkKdDsc8ZsN/f5McbY5+9Pa0E7Z1Dw
Z93tpANS3UV8GqLqPrFggBnvhA0iiSv4cdqGi7iCB5yeTNRMt5xfPJytjvko2/3B
AzJ1G14sq0N9BuyUY+Tq7KPuv2dSaTHu4Zv1MkOuECcn3UNP8xa0uLrUv3sXNLgc
PPOWErThaBxucJMHwtEIXzcuExKjCYWBZCRO9x8bhpm7/Rtin4WMHigudVqRKN0G
4/w+CA5yV52WdlQYJsWTE2KcMjliQBdbPGAiK/LoqJZsk2FssWmajfDZ3nFSEYS+
Q9wfD9mn1ziNUbwPIYmZbYMRfg7D6+gyGoPDB7QQi5zuV24Sb7/dP6t68UFX6I0B
wCBfmHA+MYjAE/MTSZdpUKN0OlqSFf8gs4BJOtHvuAFxie2uRkbSlOh6kFT067Ll
DSZyzNLkPx43WJGhYBZGYonJQsPJLwOZz8hFH3nINKeCt6YJCrvYdSl8X6b5KzzC
aL1hflSEWv2GIleK2Yvz4aW71Sl9iwibqfQe+G7r12iGEtwDYsl4iWfmxlX6hOW3
22nrhJIXCa62DCK4AfTTDXgeADnQuuj/yqaTlT0CkJm2y/FID9Bnu3Uw9CdzdXZY
9zWDVLZoL6u0ozNKZ0Y9EU6XpejOoebylZIcaDhzS2XN2+xeJlrxIdv03Ie4sSW+
z1TiVdonLil1XIFcTZWzuDtx3A4BgVeVqnxIXiAPJjaEAr/mbjgsQrsAApti0CKR
YzWMPc5lpp3IEqmZdqDpMWSe9EWPbdP6qxB23Ofa5B3UTymFcigjpU3G6FGl993Y
WtN1SwuWnG5at/n0NTx/7mP7H7C3Csns12nQbRw+EpK0CB5RsnMRf7N6UVKDrzDn
2o5oFO4TM+34zv1XX7tlpn1TEiPd9SxaOpTNG8pEUQwHkRx7cfoa6/au7lx51sr3
TdeGDczWpvlJYtc7czY2YXT5Cx141g38dT7v9efNlCPcibIkdoRgCZLiZftO8b7c
JSXPBvuPTPwW2LRhLG3sFPJ5/TVM6mCqUXu21v5gFWpyEz5V2NIw0/iKB3PI4xXR
FRMhChxzhbMPAjS+uLH6Vfzn8Ijx7XrCbpSr2rQYw+ElV8/lM7nL8v3szGy+wv9u
KtPdxUj++nszhoX3B9EDn/V6MLac6rhlncPXFuQa3nTNGDn1AGPi8yTd66zCh1db
7HQ3SzuULnqhHP9Vwerdi6tvrtuyr8XqEegDV6YoQl8EXKtlQwWUMN8qR19b10rY
pXugoWiMu1FzSaiJVl1P8JLkASCxmkj7tS0oZ+r5T4caN2JVkvQD8bJ5KXNOsXOa
b6VEuxWJh4B5PIyXnaYDvYIrJ/m5brtjGNQEPVUUj8RtGswQ5yNm7ZulfjRvvQH3
H/7Yf/49bxa/O6YHO9r+bfRxhH2d9+xLIV8s0aXuVqN0bZyNyTA11iGlw6HGcEmg
iED+mDJG4B+ogY0Aib7FaqnBpeGaJmIh3MHpQfyl02YnFHAa5po+e3Vg6AjqC1Hi
LgxxdlxSK/m1GXKQVtgOvJjTnlVT63sz9u52D04BlzBk7+pL6QNKafAupj0hO2BZ
xwfu5NXYk2aMhQhRpZVyphRwN6HZQrjvvBG4YVnZGUqC4MjeTahEiRBUADaZ5Xp+
8ijCODmKq/GY+i5uF8Tcl+EtcJUJV/xFQ27VV2wJkk0uVHtj6DOaq22Xlo9HaEX4
ZBiDJ8y1wgci99Qy7AHaeQEadbSzzTuaq6t1sIO1Yx2HmOjeTDie9HFKCQPnTaqF
Zor7zr+cnnxMrkjD3NZRqAYnopqPBrcYnbj8Vf+hYeKMLkp4tKjeuS2zP5/61CrY
ThpfpgntQtdK78fX5jk+yL4avbmBggwq6o86/HRAnsreRaXGSkzOPYGhxOC4uD0g
0kRJuVBbJBhSBCGjO2ZYpxPbGXpmH+Ljze5dKWYF1T0Ta8tE/2uyurFSfOPczeIl
bsTmaHp50aO73dw0iRDpPIcmPpGxC+9a8+wCRc3i9zhcrgNPnvAoU/TkB1+wJUs4
FY2dPU2X7BMDT7SqDjNEulvlPGPtLqAyH80N1UYhd0Ehg5Cc13/1LMIL0nZ1lrTD
gO75a5GJ+fFBKo+B+n5B1Q+XhUpE3RllSwsofkGN1rKnGtC6WEuv6lfPR6bT8hGu
2MFeGIxouiwX2m2wvHpPyO8KWhJ8XZUQiu6hYTr+I/NrzNvfeKStdtQvvGwXeOzF
b12n7NK3xajm8olfzRCPd8h3LKPs2RIjpLccTNUOvYBp7BCjQfpJauP2a/r2cFik
lKX3FBYWjBMCXXFqiHDVtoyTHUmeU6oLwwuB8/sbly4Tg42YVmS5XE97xjfirX54
ZtCTz+CiNLWMZzr10kJibX6yNHHCLrYKdIkGi/usIkOC9Q6SiZ0+/7yeqdcoHsGJ
pVNIx0+mw8GmkjOh0/2aS0UUaAZLMs1aBx9H7onF6Jf5VxuNNRw/ZQWHqzMsQE1q
5qU2y6ruimpZNV0puFbsgkYo+siA9NIjCh02Hqrg2AGQXMYJcccLMVrFaL/uHUFq
dB/1eJMFR8f96Swvdr//R4ThP8Y55JlF1xl+ozeL2S5aYobKjxw8Of2KUGhRmKl+
WHv2D0FHlP96jR2UMs1uBfr7Tw/r6IYQEnRUkBROcn+pcAMm+i6/KMAZFDvHHZ01
tfpZWnKeWUouu62OPd53uVYC0vmAZXG4vTNtoOhk3HD8He1+VegEfnEgbDya82Fo
Z/KPcmSRZqsDc3x6tv+wcUQu94N2d0zZ1d3cempfmQ87lQNaEx1BexL0DncDk5xq
vqXOvwJB1bEv8uJ8mr73JMXZPSURifDtAU4pMOmISV+4Tn3hotpALgoiZCYsDZ1a
jv4jbq1jV3JI2Xi8/tupLE3yZz8zxNAYlGpQ0KlBxllT/ONdxwF2NeujgwuXtkfo
AZ6hYRasLxDfuZa5YKWck/ZprBjIuQB2nDFzw/uBpbbQlhgESaLFS3yi76o+bZ7Q
bfYwFgMnGeq23ZQ5o0hUEywj+6RKrTRZGedj4AEF/i82LMqKwhjBSKR9I40qiZsf
G/0bREJc0y/oZDkFeDxnrPbOAhXlBoYpe5Wmo9WVZCnVTik0RGyYXVq9F/zkxSN5
0URFRXrsDGDE5d7e1CX/WTLbjtnLYMnmva8h6heRyjolzAr/3VYHuLddY/b4BaVC
hxyQzpLMN1LyAr8sPXZPuF8nE4F4JCyzDhtziwUbNGZ7GJxK56bbKxQixUdb3XrI
+9XU/pISFmcpDyvSGSmq2JZKKyAZ21YoiDjjgJUVleJYINC2FTq3Rqr37Nu0oACB
yzNF86WJJiWYolBRfExDWQrd4FwN8NtTOtU5bhGt2C0E1Xyu+GcG1f9ySNMCCnBd
GkHxlBTdL4B6YuXFwRH8cMhuY/uk0xL3VI52BvTVIWnvwLPtJuDZuk79KyI2Wxvd
2wlI75vy5qxXgWPCw3ExofFFKlZFEWGJJ3zlNToi8IzPQfGkOxriUzYhsDP6CW3+
O1PY+qZDv17/G1BVsGiCLCFaTOmsqN2mR3NHGTn8NNRKXWuvFBbqdl620twFCoHJ
6zFRfkrt2Xua80ZhTylQ2SA4H1Zku6kKX561UQtrxoMvl1BjJ83LWX/A0dHN3zsq
D9zmxb17gLS9hZ3HyHCPH0hCZFMbaifeS+pbfNMS1z4g6iyH5SxoyAw0hPU2wwgo
bmv3fHHYMTkO08Qmq1Fqew0hog6ZgG7kVgtyqzH4aIPBwwEhkYid4J95myTVJyJ0
M3/9QN9w4flELtV6NUvUGHjOHDdNopcJkxaUGWttbn0x0CsowCJTckV3qSGzy5KN
Kl4gSCXk39iHD2pYVmDoK6rV4sFG1LSouSoNXw1txcyLo+Rkn3AmeT88PgKU/F9n
iuRzJRUhojzeb0PjkrIYDzxTyh36lzxLOTnkoPkosDjrB4ty5VL+O3Bdhph7gtmZ
hltxugOf800M5fSPdUX3fJZ8sJmZTCxX0gKIvvgvecXX1J0tQj1xMTvE1uHk+PST
LotnflL0Kq4Ijxrz6QEuzdweofpvlS6U5bUHuiwNNlnVD0qYJYJpmu8m/56dITqV
95DMDzrMbZsZFyMjB8iBBy/nSHo1f1PCaxcj+B+VSa1bBAMI/PwmiJAKGgp6FdsS
+LMwsDik/0OLj8+eAIxy9pSiW3jG6mgzOiBZnXpIjlmNyTp84ia8xNshf8KMeql/
h7PkrG1xil+2FRY1ez0EBiaGT4yUfotqmNQXeowftd5iQLvu/zNj2gnpxFYwPvAQ
SDWxXTIFpIBLUl+NpJtydrkX4AzS8WCEFFu3V+ejo5rKQuMkl+T2ofAM/9HdmCUk
sE6fz6/N9SnwgRn0+gRWQERESO6LeXIbzFvzg/WqfAohbpeRoJy2hI0Nq/TFqcZY
h8R4s/hCz7F04K5eYRZaK59VWW13OlECDCALRu/g4W8f3PYr39g9QtY9hIzbkDql
w+Mi60KTM4xqPL5zZ2mzCW53PV+31QeBH+kAomnOVlxWd7kUS9jfLpebyUeu+lhA
9cJzgm1uOgbXrjsGt/L+HsVxdqJOfEwpgru3EsTHDGuRLHWd/4H6cwPwWea0GAlH
VoY7jTElsqQ2QM5dkx5R/LwK6M8tILJ+7jm7sM7q+oRJrOMvmDNAx3bjNLTGZW5k
o+rnzzxQojR7vni4gK284JGQdstnlM2F44TlM64vYMoy4RFcFPWRMr7K9D65QoLj
pRUbc4aW0opbsI0IKjVuyyQT5f05HaltpqVHumn9VETpjZ5XEAlC5XL4m8IcZiMr
q9QG7do6TkPJ56Fu6AXbUT0jAoJuAu2dMiaOoXiVfGmG9e4DEIXr2V67ZbiC1Wn+
LTz2bEr7RrTrvfQGoXXfZEx6VMLGxrLMN21EYSfCcoS0aLd1xHCs7kKQYiUaHOqw
JXOxlYQaOTVTVNj7mwwQHKl1v3mbL5GptYPMaQ69faQts1g9skhJ9W+hd2NH0iG3
8babWl+sqW1YEhBsRHxx3graM3gWEBksTA5f3WfiCoLjkNppMTk5w6fc8AbnDpXw
2vXsY3hCUPWZQDkKa5mQmdd8NoghqDAD/VKZqH3bCvOZqSH682pnN0qVYqKqzX9C
e4GeUhm1z3mQenOGjByG/CRINtoR+a3MWaUkJrc1g+wuhOMTYYp/6hKdVCLtGySw
+6/VR8NpL5yrb+OdZMplD2hSkjU+4eFkJH8qPUNFMPRPVarCzZUAOyBmGb4q2jsz
mFQXRP3Rnx8EU0d1RrpTBX4W54BrLEual2B50ygO9JCZ24Otwd3RwCNcV8IR0y94
WYylz9QQLuVevw+Xsy3hUr3FD9K6wDmaZsl2KNH73uQECIirxvqkRrtdJT3H6ehj
BEOmMJtawfVlRr6HtxOfmIbs+sZaWhMfjkRJmO9tS9vY/SCI8cLcsztX0ipx7lAe
yxvIEo3Xldw6oxdejrn0lG0Qw3BzDWgwyGbJf0ZJNJKvw84c8U1Wzmfg/AY7YhDD
Uyi6lVdjn/OBRmFy9wAKVRF6Lh90nLUozJrRbUZXH9Kz/HT0cnTv6EB5M4uWRQfy
Mxp95GLu9mJotc/moG6EDwei3JjgmyVqnkv7INXXORr5OVk5E3QWEjZWsp2jr4/t
oVWO61hTxamzfheU+vxxTcTiht8rkFzNpxZ2dbJW5uQmYZgqMyYaEAMBcCuC+8Ep
VoDYEI5CyaJJStZAuCi30I6BvmyYjLG6FDc4+e1mXxNJKYmc99HEeTlgfBHwqdoD
U9TqA/5w6UXdPMu5MBdc2I94f0WABlq020er+fOSnZUcDF3BGIg6lwPt32OlJxKg
ynlEdZgXtCaqES2yRkiq1X0zT9Ey//KpfYqi9rCGR2BwGX9zOsjlGlhfifI2M0rx
b6hon8rsOPzu4tQ0GlCcEM8o2uVhV+qUGthIm38nNg4y/AfrlKDuwhYhJ2oYk/Dt
0TNe8o6M2qjj7N+zY0Tl0vB66wIqfvrqEeLApLfUvbgV2BfGW9Ggdn5HbdWOdHb5
Tw3TIj7QOycgPCfwWdkNH14qEs9x92gWwRnv3BF3/abG8p3foQi/YXsl7GE6NZ5H
UdgkhVfrYCB4TqNc4iZeqKpj/J+aDFvronN4Cg0kOnzvMlLaGH/2oX/ntHGOxDn4
92yWj1IAdnUFD+5Pl8NbNqyf2XXCuP/ZYRX81QiL/zn0YRV5wa0GW66WN5vRFKcZ
9sKDPATix0hWeCMZHYJVygzK7n/V5353y2bfmgO54FqY3rxTng3c1rw2S0nFsius
AbAxZDVUZYkHfrexPiWmBK11lzvkWLwLtj8Vvohz+nkydXEiveSaoteKwNLUYHSP
XEKOZH2ei9So3mPQYqyue8eFZp7IIaz1/+6ZDsMDE/ZExWkcdjbpYuAMhVOOMMlR
lAHHh/sqNS97Pmv/XbuELVSD0TLJe2z/PuYpMiiXjMMvy0pgJx6P+Wvt1eIyTVwk
AL08UVK+L1ENRIt4ERI3fS2UvbwebbrMglbQFhZ+Qp+0sPPe0VY1wq3ykOFUZ+jc
UktwMAhMZgYB96IKlUfDxnVjc5kEHMeAie0Tfm+swuq2I3FkOVPeDWtlAEwS/SM5
mxMT008yDr+OijHBED0duEHYUQOHsgKZaFgrkorKJvY83TmMOWo9VJts79XbXdqf
CoHd/YuFQ/S9SxU5srMnUBBC08jai3ojZ5LASOpfixhaiWK+HH7e8M7fJHYj2NgO
+rFVNdLxflrJAKLXAANxqZICVpKAVu+6FtsVHFeUiDLydW+x8YMIeLwxRuVC6XEE
AIgBSbnrUDBVn43lq9IOGU0iW4qErRg/Edxs8VopkwQLvsjLuWsfOaYeY5OCw8zJ
ldk1G85LEyv119cmC6+YyxiovaMgOz7uMzNQoXEKspLGPxG2AeQBRuAeS0i2keDu
0OzzhpB+drgb1tYxLSkQOPbv+PKuj1pLDUCpRwiNFYSfd2zfPob3HwdA/0s3eMrM
yEfav5lfruHBq1vRLi/xucOF+xEv5KaVTjexU4VJrRM34bJUNhmwvO1z0ff4oh8A
FxPWcqW3URfhqqAz0tqWmc+s7sn9vBwIsK9vlkjcD2ua79t6bdQejyTCNdMZJGYJ
yVQ2ZguuETETbahc7mPrdgwpEv126IhJdClJeTYPsJ7wDU05f2v6wtK3lfYLlc+z
o64++2xcBtvVJt92UGtDfMSi5mrWrX9+tITbQRapg6ET/VwZNBK/epeq2x+OJogt
vEW62QP6Ah56LEO7LvjWMQpFn4a3/5qQ6tnEjf9y7+px+iNz15c2/VAUMqu8HDbZ
juYTPaQF4HR6Cx1eSnKrLRk09U22GOMs83sss6a+h0ahVa1wf68Ia8Vx0fyYyFid
GEFtnoux5rd1P72tSQZRN7gqQc0pOOJuB2M08K4DrVV7j/MH0k2Ahoz/n04MeyX0
S0zEN15dcI0o6hqCCxufalV5cYK68ddftFUGE8oczXhOtFkCFk+6HE8KXmwYkgic
Uppa1xR4oc998IR+quUOtOaQkBHFaA5RMCENwH+sUtqHHH/CTaKDtwY3Dai1vYX6
zLr05r6RK+D3n4fwLsrnjIDf9BoPGITRPXqYr5D5r914nLTIm0Mrg+NY2xf9cyDl
MwlIO9R3uLwJajCX8YAK3+Mbz69eyZVOQ3kErB77VihTsBUkkUdeqJmcV+3yDEIJ
Vm2NdPbJmJeOe0UlICXNKpMjlzdNqDTmO2v/J26Uk9OarB7xovS6AlwO4qdo0uK7
//dBis4XpAm8C+fzfIa4IfEl2JimYnT2ogubJmh+f8rXwELSIb5uCei+FZyncY7H
VxHMECxXOf8mgjhEG5ilRRI/hEpKw90YEqUjGqpp1f0FwwFMBXhuJjpyACDx+hUd
xVLUu/cf/nNrdFkok5NO1iReLWjPognhYQSWbbLR5+gmBxasWVfBAscRowRm3tJy
vPkkOGDTZqnCEzOuPGrIZ49a3Gu3RA24vTlsEdNinarapace0nXQIsEYtU6n/fB7
ZlR++pBbR3FU9D8VFG6Y5SPHHMFRaZFgElfHhCT2+AigAV73eMUiCPQ0JIJMhmBA
BREyXK9mTwz9jn7j0VzLW0OTX/ld7ZDLiTuJmeeBtueUGM/J3+yoIKvOl/Sd1U8s
BGx3Yl8Pojv5FGJNTL7vikr2V0+S8m1pnlEhBHn5qt/nHGLfITro8CWAUzLTpAHK
ofj85Jn2qCeYQfiGHsbeKWQ9NPpsZXXUrzYw1CZarPvZxeEjmvFGchhNpYBScr+R
zTfgUYvsoMg2sWD+Bz+DMhbcf8o4bdRacKWH++IdrqeRf4niDKn5bkxUBu+VddEV
soijjZfHMS5/uA4DBoVpiM4HaVdjE9uEGQxRC3x+QNY74164k/Xe6vITdiItoSgd
98htxNXnx9CcO9VW5ZoLd3yPhPTUqMC87Wg09qXdaIE3/2iBh+OnXRuRrYFnSS9F
mE0y6+vgkuSKnQSvOC7WWjAwitCXYPKvqjdRXTcZr1B922qmS4FBW6cZlkx9955H
PxejZHq1ainLtte0Dtug8i6McXLjth6y2DdiGT1VyAN0FW49m9fYC0uqGjQFw55K
RctvqX9U8il5dhdt2y7/e5ISukBBBDr7QBoh+KUHWYWeHtGQBkGqsIn/1g4Rdq6l
tjiKbZ+dtVEn6ykX+dyT/0uR6rRPgfTdO1UIHgeGs6vfsvYnmCDktk5OgbsqtBsJ
3jbb9OsBoxy2YDBbgRldqT+KKD86NoY5tgSEJnKMV4Ht4EGvyFIZeuK+p1yCEOca
srYU06Mt3p2DpORegIaKVsKywKF9S6sUdtqKaC0SKs53tPwxCTR1ZE0k7aZaYZEF
nTGc2I1rmt6J6qyBTpD0l0IOkEbzMbkjrnF8yJJyvmy7tgaSqzoeFViFRZHgGuhN
mrojgY1L+QAvurZRwIJFXSS4rNsHrR9Y/urTxdUHt7xx+Q13bI3wmlssBLTpRadZ
o3cP8uBW5fTZRwPQpDkE6zLh9qg2YGASnscAe8Jka9UylByz9mKVjwDAZaVwhK2A
wbk/bs4OfwHFRi8njbtGmtxzzI235MISdoYv6vISyuZtYZ1Z4uw/Ch7pH3lXVXx4
vcyI2DuyPhlJgPX/bXRJ9KeSYSs+sP3RnrsNhxmGrN3+9R1Xy9ruNBu3Ms8dUyBs
5Lwwmf0+bNYA6GDeF6Ri8mI09V1JXVmH5lhSmJWlet1+NScUOKRlUFD54dpq9DZQ
+QBas5M4K5PPDXfdLSmWPrXts+0DvOuFnwfUL/2hzPlvF7TACU7FrPHAbKpuFUFY
7HA8QBMr9vpw5E1g8frI2ntJvNGZZ3v0mzIsmRK4AoEAXrMvVNnpQHwqN0UpFrh2
n6q8xKIJnkJ69rR7agHQ66QIbCBRHcRPmCvl2sbRW8dIlHs+jztPKogZId1cqRh2
87x4GLjAdV2U5FUUFcBfmfZscNJL0hHkBH4Rp4DYDhLUAFoSU3DMl/lZz4vbGEc2
Pe0e8V4u37ZE5wcuidkfR7TRV1H4FnV93JMW2hc/JNpTfvBPk8vCVnU2aZ3XO/0H
ZcY0OynC2ns0NyoV/O7cmQKRrBcwxqEKUz+A4J4HnEBq3LFY3z7zcCI72tdDwoi5
G1rZ1et04khaadqfnF+Qj/8eEaenFr3JJY+OxsXAlq0Tc4X7m5kk8FvWathyASfi
zR4wQxCyglQAUnNKXa3Glcv8wLrrL6e/+xeg27cZ4XvRbUthWx0VKBZIo6r4xTYJ
lpNOrERP/R3EQMMay9V7jT3La/X5VDMTRRiVWuHmr9o0TuUf/SS8ADX7i4NHu9Fx
McU7zfRLfQ48A11Hiz1YIahOSmo3+lcxzncJrxzZq9F7up24kcUrJglcMIfn+Wc4
okL22lXDf7vv7V6uKYssxIEwNVUQML/lf5J7rnyf7Kyf8T9uur3xuroefRAP6Ld0
P/w53lYLy58IBpTNkZGeZUAfS4vg5MQ0Ikc/Suq+R/gKBEF8Sd1nM8bELHdsqYAP
mXe+24XAG0TZoKHBoGKFgqdkjTPaZ/dAyapliactmKm/p9jqH7gewqZqZ/vSKkBE
gen2bnQy9xO5f+SiAXMtU6jRmLyLFM5Dcb/N7RDURMcQ/NF2kh3IIbcWxFRPRVX/
oPcSN8esMfXoUlUHzdSxDGUwL2Tg0VJ78iPADvDHPRhGFJSThgfUm0NbskgSRhUN
A3IsMz9rX9qZifDf3XJ0/ScTJ+MegDRhL+ETzD8R5It1bbM304qJrTBLLp0xNrTM
lw04FOM5YBsI++5WPrSeSrAub56fLeP1PMbuT6+DxmuOE/6KR1jDZYIT4oPkgNH1
c8NSBrPucmc0FwRrJGgRYRj+pqPsQfSHduP+qohkq4T/PjDb6A9RQnCqfR/XWQbX
h72L+h7kGzK1i8Tajtyz0DfLX/pFMs5xlHi6LhfUJwS5uFm5kcYZypOpTlCAUAlj
ri5zDeDMjP7jlsj3MSFVpu65dTLG7jzQ9tKYAK7vzb2mkv4vGlY2ZFo+HpoE4myF
9qz+/WCmZTzJllpu9NT8AAoZ0duo52uFiGv+S+U2VnWXIGuK2Cx8hGuhYWAcWXjp
CIGCZ7WI9oxWKzhwJRrXRwUyi1zIPgZvJO+Eiw+vvnhatXpN7aPmQJG0VOSsdsuQ
2rvhFW8on4ukDD2hz1JvwNxxxeyG6xe+5Kv2shgAZFp5I7ZhpC2mS7EfT0fCR7oX
qbta18xvgueBbIpzlPubyWtDuR4enIGR8qdp0Q6KxV258dFMqVYnv4p2FzRbmpos
6CrzdksMR/fnL3XyAkw+igJbJTnPFIKZJb+7Cyfqh4WyYe57794eZ3sl/WUrIoRh
vhalCp6whLVFgqh42HzqinQwg5wG8kHG/zaS4nh3xjdAAwu0I/8r3I7G62vmp9uP
yrdCnu1LmkO2g7qX8Cc2/fLdj1x8HwTrnOdyALRKJOGOvVjC+zA5Dbt5S8ZVB8n3
FCHeH11ji2MlD2HcvsA/uAHWYbIn6DvsrFuRaGAm7uSXS4nOf9tN3y8yKooyb/gf
FBrEIFbTtrWzcIBIWh48IVCkZ2DIjzhQkGcc3KuwLX0bwoj2qgKpM7xpz0cOTS18
sn1O9oMyKmkPzFW8a7rIVsjpFcc6E/Sec/NjJsn35OAMVb1MZjRuBfrPnhsrywB9
ZW+8wyB7hxApNQzv+kv5jNsWi9V9BBrCHNOBE9h1Xe+m6eCScJMGCyh0RzbB9eLZ
eVQc4sw1RAtjSFzkIOsSpEwvgOuFaSBUp87Xi+8osqVovzIJfwj0C1uFbRKGhy08
U8H/y0bVONaaenMi67eig4AW/6xRbOYOhdsKAODTCKItAz9okdXuWevXh1ugbBMC
xPH8HRF1wW/ahE7XYaOQylwyHLxuzNiUzlMlmJ+HKI46/C9Qud9zbN0mXxHLwXxG
Smfll2169wFTizLpIYmgABKZMW/clgRW/9IHHU3nPKLberjd329/j2bzP0QvGxB4
nEi/ECJtIRwlJgNS0x7B02bojFjuvbv8TwTN2apwQ8gGQYkYg6rxhxO1Sy7f5NLC
Y6TNQgx21S4GNhJrzbDtDPQUiJ1riYMosYjmxPHKfgi40oi2WsKRUtlJfl85/Lgw
FWs7va3XQZ/am4998QnCEL5UwoE+9rm4if2ou7hk7II6WYO23eBjI3WPgxFJZ7Co
aAn3Iuvjq9KXQVDL6ANQQhOmoPu+OBByn9Xx+T2V6Gd92AYR+jhEpi075sSgK0UK
1hlA+v0mmuuE0rW3mjpfZpkGjRL1ncdLvviiQSaiORlKXasjpggnarc82ctiqxQf
Q3PD/N9JOZuSvePWk0heoY8Pemz/WeiFZXDZl3UDKZ7FIvT9a+Dto0Gr19nsxKjj
pSC6RmGNrTk9Z2k2VUYNw6vbkZoBR1soT2IW+giaHNmlxdziaHWtmbJiZg9t5MyX
FM8JaQCzS/gI9zCmhHSB/k4Ua5rd3cNiI4YilUANTh+AGRsMxS7zh3WgAvwlmRYS
oTocoebGW3XlkrOdCou/c0uHGk4FNmFpGmsB4ck3k14h3ouIRfPB6nDWdWbJcV43
3FWLui1g66x7Sc5y5jrFUPAhpJixHxc+w3Xy2siknHq7dzc3fwApPwftUhA7LncB
B0Yf7gQdPw3piZQU733NL8fE4NjjGtCnKdF78J3Y2eor03cPvkEUVT1tWc8UxoTu
GhwUCt0kBU/hrME+hgWEWI9acbRZVkrQVA4daSqbK3zp0aY09eOlic2+v6e6sG5h
bY1G/rYDDc9ojjlU7a9++yMkkxyM/C75d8Ly0WXinS7STXxAZU7AdnH7N0UeP67q
AWegNTr7IJYQoTXtCxFJCt+55zKnzi+vXW3uTjo//LPN4bRbFtg5P6BhU0et1MF5
Hiiw0vYZ8etWkTij3Zgljf5Ppd3M6djimLOY8dV3QQGI/7sq99zcjAMmySfs63ED
sYJq3FtK/LdwyuMlYSbQ0/+vu3alX5MleUhBjjtik6BTIDsJ2hmVQq85aaEaCwK3
r7wd8gCko21xwr25Un6Pa9G2whPjrrAFWI9lIYB9LDkPLTwLk5Nx57QPuRh+Pv9z
slAtxZnTluZcUNixEzTbuiafC7u6QtSifzZLSWgbUqIFou+Fp0uKJNsF1hJGigMC
wEAuyq6ydzFT8wH88mJm9qIUuAriA2Htor25Slvp4F9kZtz4v7dTaLRY9SDCcsoj
gZ3NE9jg7Xd/X+aFfCASaeta6H2orF/aNugnZZfasekDpFpJMBQE2/lsNHZ4sk8u
f4/aoEt7gAJyqG20WzkMceJ3VBULIKFRwEPpEd2RkIZ1/HUDvBGusVh6cJRShs3t
vYXWW0SbTjx7uPN+LjA/WC7jHpoQ46RGvk+5sxbtB1f0l8wDKsHJn46rMEsCIGB8
xYigSqAZvzqQPGPZJbYJUK53SVLE7CrhNRDHYE/PlI6xsEObFi7pwxIsfz6hcFt9
l/YapdDI9JVWJOfFLlDAuQGOpHeT39UV9r5B0tgjmmv77gCirj01aOXkU1RqXxyj
qRIr/WtwZMv/jp+if8/Z9CsFsuHpU8++aGsACFGWU1SqJmlkd5aLUgktbLnqF4Fq
mPoEJS0QL6NW4wDGUvroBI2YVcKOXeofdAU69SauPjsAUwbEKhgKm/OYzrf+5TRC
r98j2yN1I4TOG8gjhDK2ciBhEUzbonFgg384AEiP3/LT7ys1QEXRgGkFBa9i0AGy
t0Rq0EMsFvxX17k8g73lvYYF/qRyEuzoukQ7FajUnMB037hcH39pkcSON04AiuA6
tv7bXN157BzK9Uvyd+jCDpsFoh/ZYjzkWr2lu3jNVe3b8YSI0ALrWCv4NNJbRpCT
ChZWB0GpUsrGg6JbWdXdKZ9eFtwYu+0JiFc4r3gM72OOIW0KKx3vMGC/9vo2CRy9
83mTIxjB1JGE0TMYmXVMOKlzHxvyU9n8HTL4kV6C+dvjBAolkfqcL6tkDw7dwAOt
krX3TAym34OqcmFYQjSAvy9LIPGO0/Y0yd1P4emdBN0U3uDTEtjBzkfIQ4wW6sr2
P9x1HHc1rUr4D1GRDqcwVAi1LRJngUzEJuwHuvZPWJMrgrHddPY5fCTEsutcPu2X
15R9RChRreRGgKJUlBVf0/SCJ5lCYPbod+81J2ELYN5WXi1NBncLFQiZ8wKaThqB
FAkLpTLsbibw+v3sqkfHo/+j1VFV5fvY7fdLtG1zPQFtIOdFysKtEL/b1uAUV0Nd
HGo8exfhfQKWO8Xcv5jt8fZ+QeZ0N0l/xw8ftk1jkEvYRKhvQYpvNDYaRz+p+gtl
RoEF4MkE28/z2qvz2kA8FwFXsyMKLjo23U8ZdrMRY/uMFMNEPGL7MdbpvJFbUQhc
cYoQZZmo3uq8Urwc3KUFVId503z9a2A1Bf7AGflAJyNWd8UAwE8GYnscB69PNBAx
TaPeebYje77SKHgD5X8ZFe+rqYHcNj11v174oiYgK0VRs9eZaJT1+dAdedW6io/m
LpZ7RId8XbyUgUVLK74bBJF+6L5Lj+ZY6ndkxv1bX0jtuKgDqQTLzpiCDyb7EDx/
yjfw+vjsBvaMH+nhCWmphsvKizNv5Ft4PpCZ/Z2/4jaRvgnzRwtHju+RULC4iB72
4ozxVNizsItcuXIRWJCwh9vEb9J3xmPocgPncopSs8IK5ivh/sMILCkbYurdZO+g
xmPlR+IAWClApTMi+nPKfT9ecfb/FYb+eJp2aZYq3zLT2fDDejm0NY3FFRWdysEo
8WXpgTmSduZHQhTpl471mcYhKHFLGXIdjoxRIuR6aa/p/1EuEvbnDvxZS4zYeq/R
dd9h9RpAhlAn13FSSW/48ut7/dZblyQAj/aqp5uSUJT94JIzNr5YDx2+naFZ6cXf
qCyYgA9f4JT6F7UMFTlhD7ik9t1MWGjvDOil4ZdCqDNKd9lDJ14zKiCfnun05qXe
jJepS1cG/WPZJwAA+iOI0/KsqU7TdhswIPOb/FEafYYlBG6OT290bpR6mZrKXTVH
yDrD4it6EI90Ivcq4sXay66UxziQKrCXUY0DjqNbNWMGzAcwp6tz7cu0CY4fdZKs
Zx1i85r97C0of2pBKH8fDPzwgr27+A7f7ibHK/fy4PihqIlDbSkPZNrbDym7m6OE
eudzYETB+nkpD64LWxGnhqRWp3aF0bDdAgqoU5nE9g4XVs3E5Ib4BZ3wXigfGAWY
Qhwm0lZL+1EtxC2fB0Mvqtq/EFZOD+i0IZsT18PsljcVQPtWq9TtfICqfQy4exKH
4j+H5fT7NrGWKgjj4E/YGeRa+dvo2YRR7qppkRrRoFpOcERA2ZK525762+1cCSI5
fsKoXhrvE1ejcewkXMOtxNfVCFUT12rDd5NGlJX81byzIKNgzspo5wSt2yjZk/k1
OtZltU1lugfqwubqANHXXgps99Xncl6y/W9dDrGhDejQpiI28o1K8q/e5HyAEn38
XVmsq05ogV/KCDlzfhSZ3WtPJmSce748mk0C5XGVXXugoksEM19px6XbB1WEed+Y
qN61w2I8lS3AifiM3rUSesy7TNP9CAvM0jeSpOI73uKQwH95iTCtm2Degw6gWsNJ
DpZV0/STCbHZv+WIU3/BG+3DVcvwK+7xe4S5jBVN3T+/oc5dBNh9o6Ul3xCz5iUx
vmsN9MPqKjvuSWU1UYWIulAVe3fS1jd5gNYr/Xvd7CLs8dQuLXYi32gEMx8kAjOX
2ykyrQ6U/p3m5xcWtNKbpqnqt70s0hxsy2lTOxdl4VRoXZbcCpSObGrb+09ZywDk
S8+L8WEjC0HgKA+P1MBQ0HALM6Gbj1S7PI/seasyoUHQVdZ6NSLGzmwy08kewYGw
T+slXpfAWnwbZ5RhmaSlfE/ihgkUMKTTiG/hP9/ENhlZYWcuL84AWrUNYWzapWJO
mkn0iAEUC4iM0aN5MHKZ9QIFDtTw/MaexydHbXq6teSwLPVpp9wo6zzjoW63qPr6
OboQ+bghpKb9gobtgxBK/J+g+KWsaVjCqfII+AN5HhGJiLFO6RxnyI4tSOMtHns4
Iioy7+zK04CpXt7BPwM43CtbL2eDaYZn3IKtymkf8G9JzN68Q3OmOCnWn9sfR8/I
IVQNW01l2S0XA3qskjUVG+lGi5C0KbP4DDz8cxF8n8Gvb+RO1J3N9mx8oyt7vvNt
3opYI7R8LUfGHioWFBv/tV1PEOTvSVBlZbHCqJ4SH0yZGfAgmN8q2ijeJi0wXA/q
1Bo1TB3rq1Sv2P2C6SSgx8KuWL/ZaLDlFry2BMIr/a81SMu5LdjRbeByYZ74v4l5
kgJBRjb3vx+4nM5c31znXGXG5BOStM+Zo5PhVqHyPav1w7LkSaJT6FD+Xk3N214M
ywIjo3KclYgZRRMy3d1f4jennZN4WbkVqApiXLixskRITZkfZVWrqCNhzEaj3QZV
lyOol43Al+2yoNQen0g1dSIQX7VrnXDoNJRx8sa8mefoGW7/QOhL4mGbn5wbsQxc
LZublnsUZZ91uN+erQxR83huG2qalIc0hH+68T5nJgQ1xvmuiU/Vz9pqIGW9OQSB
CfgnA/jvgY/3xPdulVoTmg0NHbZhYlXcKSh5ycirSqnJ4RL20HjN128fxUYDXByC
TGCeK4IJmECuD2re3jzOgYPrL9ccLk3MGaSwLh4gzsMr9WReGeoLx0c9vA3IHsqX
3zJsDguccgIlQjbOr85pLH7Lk3VBCed2lzcVh102MJ0xHOPz3YMqI88scspZ8ogE
4CEMC0m7TH8xYLYJ2gNssR/ZSGQSg9v7ajqjXdXGFquw6b1ZZJFzuX/XEL7gUY6d
Lwp3qW52XKViakhpR57bUwsPWAMniIB/V0GLnKzGAjStndi0V6FPR7TKy3bpuPd1
IyFaMKyYhzRS9gIHWIHOVEl0HbFCeyiX2BM2j0kr/qk4v41MBzb0h5OLhoR6OM8d
MJzkx3t1z3x9py1Cum+E6QmYtXJUnvMtK6jfw15GN1NjZDpo4ug6MVeYvGSlM5JV
F4C/cDFP9BScroIaWP/osATBRfe051/EAjNNqYZGKPvPXU5fmxf7O/ItONLD2/nj
LaV9Tk7arnqg6BppylloWuCL0AW+jlZ83LogV8mCx3hoF9ySa2EbUhN0ib6L/yCi
IGYHg1YrzsOwHbdPA7+q4Y3yB7CndziUIN1YF8fTppKBl3wXfPQ9MY0xrFBboZCA
xWjlX8c0oGFz/qg+UyFzKI2VmPVjVlnLCe9mCA+i3FbTV9mEAUVTWz5K4LMuE+hj
LiRLCsVPzHOOB01ObitMAe1EJxtM/BQdLI2kdJIadL5l0WmsDGWh4TdGCB003duC
QZRLzMhjJvLql3r7SJ7k+YW8IoZLuV4NBohEz3bKd51xTc/k0cz1TAfhuwvwOTrl
IrnoxbfrhthR5kKVRQsjms+gZ2Gmygxb4Arv/Cr+Hir8a/5J1jFmk8RyP1QHvVgt
XlmiDDp5KOu8bEscpOobONZQdjis9JuSKx7Rqryqq2pRaxKN2So9NtLvuL61fqro
LRu0BlOYkvtMyiG15dWTrz1hoUOwXzmZ5cbzlvV0mHRQyoxM5Fk5AKvdvZH3ODE3
wWnSZoKzrJ5HZPKadDic3mpUXWNzCnri8ULBcOssQrRbEWuV6H6t73H+R9YQ+Rn/
FWyzezMQy2lZOuFziMIbN82com52JZd/kiOKDRCILIX37bVKNQ1/Uw5190LA6nKg
PPb8Xx1nWnufM96QG3hdQ1w2w9842TqIVRPKW/zfJ+8NFfLKkDVVD0puyC4COPJg
CvZLQcePvIt0QkSHS79Vs+rxkCfNnxLaT8JwQ8ajYZsekt5446ETwacGQq8Uy8J5
jZeByOy9SQZ/4EMGwAEaTvDN3qFFmB77+XyIemwKn6vAJ5r1VL9Z1oU8XyicJrko
0elrlFqyLpAW0rPLmY0wlrruzKt9sNhHmYnSFKys18BhwtxM7i3MLXpARSzscA1R
ThSCtTXYalgbiF3CY7zgtYLUHsedPw7GbIW6+HXmF718Cv2T3ZI3r8YmDDs/Wgxl
dt8iQY5rQZBZJ92PGbA7e0SXOYfg55GQegrYNLbMNB0zZyA7PwE2CxhrJilIFV0H
pDn3u+mSO4PiTKB840yj7+tBNaldL9QS+JSogEFvzjAxanek0Ph61cl8W0WRqEqP
z8tT1pkwQ5xx4oZsYGV5Gnb7xtoEpBS0dPFdIE5k1RR/ir6Qo+dJoMTaaQ3otbQk
bjkbN4geWF4rU0nkhgIaPaXy21MFkGQrL2WYFNhymaBdMAR3c5W4m9W73b/AqjE4
N0wjEu+Qfh/ylFJDerSNvYamRmu6L+NHdSbKbDV4F/Q8rziZpPfP/pDgJr7TqgpN
pNq0oIpAD6TNi4QsAMlksfDqatngbf0OCITrEmhohcaGxAEqQoLiCYVM/nZ0W74h
lTtmzmtb1IOr8Pgiit/QB6WSFrA/GH1e/k3OTW4l5uXvQEDzlVEWmGP4adlNBlj4
LQYzyN1nn30drGMJxlghPyApKnikc8sKM5sEj4AyfkVMbJqIvjj/IS0MNx3EOsq3
6WPTGpQERHQju4nRyXh3sRq3RdnSADwCA6vBg+D5jfEm0NM0K/FMt/8tNOucKUdf
vrd9r6klxgiGBApoIlDJCSXxXuToroiQSRWfMnrs7rermzc9qyW7CY7Y7RorNvfp
AVwMI2NJ0Bg0QcB9+e4bg32kmUmCH94ImCOdqqJKZAuWIFk8tXQb1VuHRnBhmUa6
0VFxFo2O5rKvY7nPf8DfdKvknXnLUQ1pWqLH6NGV3yLxxAu7Q+gMuq3EeFpdddjh
NYTFAvjtwyihBj47z8CsY8Aym9mSauoFNfTvsVEbFALq2i36vQaditWaft4MnnCq
Yodk0i92A9rv8rCtwFTeLh+2h8P3wk1FfO6X6r6WRYfwr34ypzOFugTF8BJVOzb0
xOXST8iPwXBMO9lN8qWe7fOAMneYge9J9dhNrUFDGPAkg7GnklU7h/K74IhFvheg
bC2qXouGfXU/KwcPuy0/ZXR3AESfxZHH3GSKwGFG+IeyhKIdpc/ZfZwsVyG6IrIr
ZblCwTkRBm0qF82cQKsu3V029sVPqUsED6wj2t9JfB5yzLTVtZsbIKaO3wm+Ju3+
2RrhbZmmr/up/l1WUZdeyNi+UFvcvq6xz9WsQ1AYrRMhIfofAQz0RVM7Z0rNWXYF
7XJBTlJeJsdKjQ9+epgyoqhvHeLK3ssVT3UotTjJEwKfPG07V0RKZ/1UsA0jRWfH
cFrVrQ2HT6+smQNsGiKfCqwPs7k2iunUnCEYhElIcUfjJXRjKfRLV4ZV8XXtr0p9
5LLdnVytvKID0CCdumRQx1GXQhC5IAK7Y3AzU9LuZhZvN462DUDB8xhTJKG6TwPJ
nXfYiiC7sr3gxPtSNrOODD0A15OTP6zPMLoclhkkf9YyT28kz5wb/NgsCAKPEmF6
IgRKQeWHhoH0cEt1aUdjCBxGSXouSkrKjQXYd3hzAN3THBv9I5nFSYNYklSqrTZk
nMKaDb8R+mxhqrQL//7Nbmcmn78QnS1qp2AjOzJZo9x3+lUaExG/XK4+6DiSB3jG
AS5gw3lj5QIGnLa0BWUoNoQs2kWkD2LYoTc8vb3xz6tW6rvOr2N7HNWmbmi3hDkA
JecaQns3Ku/Jy/7F1rTvZgV/DkHlgYIu8r0rmYGbn5ZV15VNjCeoO+o6mPBhCUoM
IFKsYl29RCQpyCxrFwZT1cA3n6qowduyT4u/mun/7f8tC19c1gAQ+xnbbMk2283v
pKroeunEVcX5GkZgSnXLxn9AXRuUITU6N9Kb5ZVLjmJEK34AN/6/Ka0w6NCxz/BC
IICo190sZ8pLa1V8gMyKIfP1mBuwErPVa8VNIiGztdA0D/yUqbwcVum+dxwmoiKT
cPXY/QGdnChP9e3EIqNuWsWZxDVa3CM93cSvsqv2CzRxoRIdEoXtbImT7He713dh
/VQNcUjpU1Wm1Knb8zne/daJpmGJ96NeD9MkJUdRlzC9DLBYzylooHMIKufOU2eV
jNoQ3mjsjrut7+1QfE0vtDtEtSZKH01X2w+u0cV90WTwLPfJCNrbbIA8EaQgQB1u
E/1XZ0PR8I0sHDcb0PRIpFSuV/Dyb0CkTmmK37Tacb0so1WJJUGvFcmaLqnJI/VT
t77IWYAoVYsRMmMZ95znylSpNyh/qZtCSnberQWbqKOrN9W5x++nTvW3zF+3uYg1
jIpZ6B8RuAf4yVbCDaxiJHVazBWg0bxv9VUsT3cKCya2dWl5b9inScOjNqVOAbnA
M6n+NN2+uSBM/0epKOIKGCO8G3tJZwF4Fc0DHdIjL4z4jB7/zZuhgIcdH7Fp2wz4
wyLUe9b4vVU34dv6irayeHxBdewzMkHi/rLTuRTrDC8LK/NruGzoVmznap2P2B3J
C4oj1zk5Z30mYY3gnvKWrBtdB9r35+8/pbQ2BIEw3629F22pzX5wsYQIlzKnT1Cs
bpMq+pvJqbqAkgD4xUmSvA7GrJgbZNwnJyW3Wz9DCM1y8dGoErjpNAJqY8G0DvQB
Mk89jmDbbNUo0N2LdXv0oCKxqHTrUsVH/njxmNBVBMTUP41Y4YTJ5NsR1E7KFCSh
XIvVV0vMd/OZXzZ1GL1p0nMauFZTUTgpIONvmlpmbNmkqfvW6SJssqEQOIwKDLfF
KtKkJ1uR0vnXUvlGuMjXh+He+LgmoXwDyIfrS13X23/cm4nLq7Bd+ylVSMDZULEf
yqrV/kJszByNtQQZO8T1ziWW77bS4IR1kWHnBI8U4IAjXU8ZlrT0VqTO9J2dt6Cs
ad34DVNrutlv8UCxdxMuKG0dkMio1/zP0GiEzS9faXEIAOIHfCjP/98wAsU4/134
PFe1IsNthJm/nQdzDwXFUyoVNapRyPRN+dRhaToQQFRd9Y7bkmhwURBHJUGbknXy
0htUK70kiUxjOIA8aCFtcJdSe8shjrAjvf5VNL7jHIYldetx4P0AipSxoGVg/NRO
CuCY5p/WyinQIwPtosx5oCy47qqFqSp4SoAI+F4fS80chA0jfkeepqd0X2lMYKQ5
xuasj6e6ii6qDyRAuV+Yd0JLm28d/uGnvh+R5OBOB6oEjFZurqc7vCsA5JcZi+fG
YLHWb9rh8KlwRItFcKgXnATMPCBnn9gAcl1z+d5xeXimpcGyw5P2nfXIxbc0jYtE
qbMhVJjm1ZOp4oSgMyJTO6MH3DQorTNswah+83L/PMs+2Ay19QJRl2i1/oG0WXhR
Prt1uou3hMUtPPzcT1qEeH1CFAKkrcyXSuv5d0NWArM0J4Gp5gyOtiZd/admK8SF
BwSOJxpAVO7aOvCBMAbAiYfE9HUVNnvP0jLN6YHcsdcC/Q9Fk8FxicmrW8Sqv6Jn
UMl+az78TyYNWvMJ+xSLBseg/97DTHKHEEU500MvaHgu4fZqC2uDkQIvbdZm7vA6
Fjuw7NamDARFzu+nSqn4wnzHPr0CoXQZFvP49w05H78ImNEOxoaXi2aq8VIAjEtr
TxPvc3xtN+lCZK6Fz8+aLTkSy29BJiMCJ+pK3KToKNCAcWIUj+wCTA/jy/zLi+4w
KjcxsihD7gHfQ+jiXUilQ5KdeBLVX+kEv5OJ+MdoHH0uooOXy49fnLMk68iwAcSE
ZHljrgeFwDFSwxCTeY20YHEjt/o90AQUF1LUQwXckPF3ZGUQEL3XRLDIukjj5O/y
oeI7q2KPSKaphz2J9JjDr2mqFZqLpVcNJbejQnJ4rK9YJ5ceXdqGgPAE3aQM17R6
0CENPv585pZoooLj3nvGUkXU8MaQP31x8Zs4ahG8JYemHQjuzg/DVqd+FbKZuX/l
+fTsXRtQsxVuLW+/HEssCpAJfaN6IVUOQaBQstjLJzVTwQV/nj1/9FI/N8WdIaoq
FxKVfx6bkstYXPmEDtyVd7bWcwlrE+Zng4vaFTo9r53zt5VsT7rYr8cX4kYfDWwT
acTOaPZqjXLIl//xG5gidsSFxsm2kTQ8alSvaCTq2IR/XM2mMfwRPQsLmk0m4ATr
mjMJ9E2olIScNJQtLF/h1BIRCVNGGb2Xs/AwPRatdgO4bHVPdoCa6Elch8hEHArH
7QFqD6rh0At2dcyjCMfj3MnENEKZaDoQDvFAOPjm/Xiw7G6BwnCyfMZsgpt74Qom
LzaXuWXWG6Sz3So5PT/QKn6ivyBvzDhU55pUOZZIs5CtAs5LaoE9DGLnuxnPRrWQ
8uz6UHGanOVJcYbluDn9QIADGYg0wD3Ife7NSA+aIhCAzIVy2cLhk7EYh2N6U0HO
ChRjKDL3ksuCWN4V8XrnSEHTr1avquD9hQbnt7SfSU923ETvo9wEsS46PP1LMZGd
YLFXJPUV3T8asJpW97oJoCVlbS+zFY/H01GFvsgpgFEgG9JxLar/4Btg7wbFcDQ6
+RHRg017orKsTlWgUoLbpAe5LcKonSCFmNiKlpQJbeTukcw0UvWmMLwfcp6o6dXp
iTSe2CT5xHeazjvxQmxSv+kDQwxrb78ooMBCUmoMwRPqUIwgC+n58JPbAO01r9p3
J+3yvuXb0LngEIX7sD3LuNNPQIVUFh76VkDmR5nFnjKs/TarfKvkUzWFkcJxU9Cm
gBP957rnS0uAo90IK7S45ze3TyoIsTG2XORdjwbwl4YRvPF7qhrW1ROO5jXP3h4s
l9ocAiW5bmE16SWGQg1C0ULNA+5TKNncMH4OljWo9C0UF9Jsa5/f4t56fVWDQ/a3
i5a2JA3CBAj4ZDrdvwmIBhkMCtxqNJwz4dU5RsorBwkxNQHCWLzUjkQHcQEXBVmp
wJu8g5SCo4lMaUVLayZH9Ag5cOJhlEJ/ZWlRZ/UrYVIjFMudmG/5bsXjCGNTVVVF
rnUv6XPfK57Os0N8BiMmoTgNQZpIueTwjIw/a73fOwvjB/jiqmpe2g/+403mVZSK
uiONtWFnV/uBMoFAfURWUmPvyUyBCfLW9NqD0y+Po4iqqXmjPIq+CwYIs/BIWj1z
Heypdmy70tZ/jNoH1QTJn0mrV0WF+lQdmMmxsFuTtcYHURgie1VXHaWE8aWk6nQN
ItbDhbPRImkXuP54P35jiZFPFNDQH3CuoU9HnfOxJeiVIDtByamBeIFOnNWNxnvv
akdvMjMVciNjyJuWSDLhlrtBPa4VcvdgtFNIaMCmKp32YFLkqnwms9jT87IBoXoL
8A6X1UUs6CLzyZ07mB3ul4j7ROTSF3QlXucIHKCEdr4vy7JgeoPLtU+Jti9dMi8G
mblVIMJ8JhglKj6e+xSY08r2HilCd25N2ZABetd1dmuSYeRWiqAheqj1KoqDU6/1
idr7XB/LiJ40Mv1NYxGcqUGNPSxMV0HkehnAUJKt92XkyqiNDIaQSDDugcqV6iJv
DPBJyIGn/T2d7CGR6QPIlGu3Deh2t1N+KveFA2AviEfQ8WhAQGwFu5F8Aljo97hU
jO1uFIgWYLgzIJlM5Wf0+YHhsmigiR2jcQKqBjAVetyfkB9QkN4I9S87JHiSdxAu
QxsrBp673c1f1PlzoH82/o7cR0bHPn9SeuQYep+RGJpXulswXvcj9aYyns1eEDjz
15hUt7Mv+NS9c1yCNtbqm64Gzdx9ERR8UXjLgz/bDsIKpR4KG1/oMjJY6r9yib3q
lC5rGfWhFL375SHFa4oT0KbaCX+mOUqnzBpWbNZoM5isjBfa5tayo72FClMh4xcZ
skt6tf2wscBWQkPJiQMBbYvp3LgzzNQG8HA5vu+HByp6FFbW1mCS5PLtj1YcJ9M3
+g72ugCCea39LYZNs+sB81nann2NKK3+GxVuIkWnHtZm9clXA3Stflad94VCKg0h
WYAl2MoDU+DYREjIe22TQYRR4X7Wn8o7nEofoZAyp0LikRBD4ggFrHpnJSy64fo9
QgFjJHnCgOwfrqSe4gTIvRVoJT9khN7+aMF36I+ynMcC0g2bzhLZ35Xq6jO7rezr
1TaUB0wO5rO6pNHyveAzgLtO/VR78oGT1b84F8YiY+Y4RP7KqoEGM3vJez0XPs7p
6yKxZGz0g37+z8Ur5ImfBSIImNWTGa8lFn2xMf5q6wwaIsYhGyN13LmOspYyzoBq
4NyYae1SYXkQHf7QLuSMD7tdMbbxz9+z7nkssku5o2lxJnfdqlQu2M09O9H/45X+
7FNtKtIeBJUTFr4dvhGgCOzdyOREoVer2zpm25C2w8toa5w4N4aaO0HVgOw2Rt25
7BLchfeJK6pekjq2loHlaCW5SqeNJC2uQijQoFv5bRyHQk7EA07j7dxcAEi/lJYA
Pdl/BJ1YeO7/5lwyjDf3UgcFXUxb+q045um/bINWNv15I7S4+65JWjiDKauK6puT
qSuR3FdC4uaff9cGZs2SdOOAt/f/VdhUwtZogkNB4FZ9H9KFgJcWS3TdgFM/Dtb4
Uq7ktGvN78NQp9QdOK6SSyqKV+G0b2ySLUbsomhL+Ajbw4NpsFdchGhltVfVjVh/
LsfMoxIPoBtSZ46513d8zJzXUBJVGUQ0YY2OGE149dwD9jOw0CLpAzU7+2bGkYoP
gh2pIQCqy52rJyx7sDrDmKWkykv3nEAb1wsfJY4bShPp00s/EzhUmn95pBOkh/Uf
7Je5RMj3G32723RtAirArFj5bBJKHgQr9jclJ0h/K2asjG3B+q4M/O2TEGYUnBfY
NKTyg2BdWugjcP6LfjTq8z2Eix+XxFMG7j0/SqMcNESR3D4nPn2T47H5KfmICWPs
utRsExjSAdzfKIE4ibklp8UKq5RlG9I3YTCTddec8JVWjagxKXcbVlsmpec2MZ1m
jgAjpRQA5gfBnF4D+6S27gO3k+5Lh0QyEOJIupCnwEqQ5TGTEheZnxZ/Xn7VPo4J
jovZcinv3BZryIdrxIGHMOo2klZY/H+kH2u6vVJ9PBM5DUmXLyDBmUTFhvcwRKY/
G064CYjE+R/LNNPL6uV3xb/iNR2MKOqvL2SeHIzVLe6CcoS5iQyZ7anszFNLkdJO
VFIxwSDPwQWeuA0E4Izm2ViHkdYZbf6j0zOJxH6bGWrXF2txdM1iJ/S/lZZMARAb
6k6iK9YfJimusGzt4y20QNg4Bl86ns5heKrzoh2KeLH8ZFKyJGTmgLPdx3bNJDLM
q4fExOupyn+mjwYm50B4UgZDyzFB0vz/CoZqKPjM0WDLSBdPQWcZ01w4EwuVYZp0
5q/x9ico/RqcOE8pJLfaj5788L8lGTDlJIITnVMxFPQKsck5o3YvHFjn8Q+R5WpO
NN8GEjKghFJG2mlkI2npYs1w8HgQ7T6kld0lcUTQxOnLwQe95Pt2k+eDe7fU9KSl
17Ue3DRsoIQ8g4nNVbKtMENBQJcPd7MLnrX2dM/yNySwwIebgMbUsrEfnQlCcYED
zj6KWuDwcX3F2sR4blRjZe90pGeVgOWKibZPU2BQEGVbZnJ3K3YynmlVPi/6xjAd
BGwlUKhQ+Mpeg9HgSubCZKlzDIbyQ2DdL//69tmTZ5JiAIcm3R3U1SJR3nMfjT3M
XBKHjuCamNTOtwiPCyJe5HPq8EZRX7VkPRYwjWvPyAC934J28+Fu4hXftmTJ3feT
syMb9/fkng3n8BguOPviNbakzBkokbE31+CQMZALj15bw+B469JwuA+aHwH1NTZ4
CR3gBMp3JmroBs84kKBcME8ZAhxsReiKl5hAJoDNzxJLL82qsLVFLqT7ochOaBoP
gqHno1bKUdjSbVtNCoQrbNElO82U2QYjcmKi8v3nd/Dpr32R4oeEo/tcDaZOoc98
wfMFHTYy4S0p9N+mxcOuw/tvTUAyGwfFYC5vux1LWf7Lx9ZASUq6PUCHOmtN8PRD
pKAYHKo3A+/ZkiuiSz4XMHyDUBSLoJ/w674OKr4Tkn9ihTQupHLqH9FCPqqjbFjE
EhILY1feZwsuar1BbI47R318GYOoL7lYaBoD/wQVxHFkJmsDtRgLJFC2M47PgMD+
sDDeUGcsBmqd6MGbII9Jc20+OvuCZT4t6biPd100/qkASOToA1tq6vgyEzmuWzMW
HplEQVbXf2tOErES/YrT/n277UlF4E2Re4iDaJ4SWQQoLD5b4QzImTgtRjXSIwoU
lTMIsyK7wzx/RIzMiEXwm2HTDzHeakpIPacR648+Qq6XeB0oMuUchMwCVJe04b55
dppI5RsIhE+OxoTTd8yAoxYmWYDwm8jSHMWhribP9bJXV/v/oIiXc28HTb+Cec1d
HQRsP/2I0xUXa/RZgM0QLud8ij3I+23W9wTIV47p99X5gbuY3bGEk0NxxkVvc7jy
L9ZI1ovA8wHHHNmxhTAXqtsCqu6nFSWBafS/EmTu0HhZvl/IhVQloKc5TfojnueZ
CEYeXxw0f/QgyfVqD7277+NJH+tmThIguxaUyyrAv4GmlJeO7/vkXsS8jWMyRPll
wpYsadI+54o+EIQ8H/2tpxSPIyNrHuGs+G9aYXkAvwU7s6JI1+F9fOaDSEduvJ8W
1ofjQoY+kFr7vSti+hWLvefy6nPilg3/hZmlH5vUGrLr7w+UGVvc0dct+8g6R/M8
C/sK4jQ7ZYHt1pUw6OavPJ8QskT+ICBlpywwsQe4uvxU4dPWDE7Ch6c5u8sFAQ9s
nEBRYVWmlaA5onWUb02T1g7EsfkZSh5HJUxacrE7xeXHSdtanVw3ASSme8dhgeiB
tfUXy/0vQAMGfmoUcMDxvpBeRPdQGzpLkoPB2+X1pvmAku8lK9l/nyr5nhXp26LY
xTShry2hofZC6HmOtRUvlJ57QQMOTxvqK1edkqbBONqn2R8uFfvplTq6WAOAyWgC
5OPxVPAy9Evc/S4zATKBEiTEb6ZKJehlqiv6IZ9MI+KVu+lqdjsymVp+GZ+qAA6R
v9a7ZRgYCJ56R/0HJ0+gNBdh9XfBs2YQgKZ8SiWT+j0sSH/CJAFsqRL/50/PFO0M
0DXQnAN1haW2Am9MJbfDV8pgvpXF5A9Cg8rBnIRSfDd//vxg5Chm8gsSEIPWbXb4
Vb8KoR7VHd81hhh3HIxjYTOLhPaMvmG5wYTLnDsmDs34XJDTRuKi/IowFOgwG7gw
8IsUmAHdrgBkTB5oN2he+5j4Q5ZY9savlLv6yyHNKXnE0KHY7M1ickxZKbmQ2ft1
JNJOFSiB7bA0/o1YLmzgsJ3gjiWG7x9ndH2P4z8GBu2zU1fRpY9CVsXmyRzVDdH+
BuJfz3LtKsW1MNlNbE4g1K/5qeapuNokSKCwKTCj6o7rrOUS1xLZDakKAJEjFSmq
glCp6QrJHNwlfapxyS8w+KJdequqkjsXCN5dPtLVaax/GEQeytBDneizhdkwc65r
XLWf0D/s9sDcK5+CU4GnYKuzBuIGOYT2422Rs25T9ODrbeHbNGuxzhOKmhbz5tu7
oLzqHQsZx+MYpwRedFmcX8aPOCVnafU6ufAjBk5UHYtdkKSJvnCfefhqlwNNDJ2i
1xTKAtxaXM7sDXYvvXA3TJTv9q+CuhkZIGXzjtkXpnEc3iOBlElgWVhbnds+coSu
pEfsuYK12Tqnkc49ArtmlS36iKS9ZlPJ9C58juip1qKpivVgGDaDxSpxpx3bm7yp
JfZgqCmmvCvNl5tuJthkc09urmIHiPS9OuDSdhNZrAZZ4PQ+rKOLu9aVCsRYja67
qA5AKwZofNq2HMxflZm+guar4NbqdkKGHd6DL798NImAcDH/rTk5b1IvC66VrvHV
xOrJDpco/e5b590wc7PQqAQ5j32IQ7Ki8khbzsFK7ais4BpMv9+PIaRj5fUt2i8Z
bUxf4jTA1pmWpNSqSa/zXlLXa73wTiJZh+csYPwpQvwlFGm3ogywaM3yMevnKD7J
9R7He1hhgQzbk1B1Ocg6z6hbB5xLX0x/QogB1mVZ9yBG6Ky1XKy3l0+qzbHZBU3H
HONkYr/YlnvwudGzAbBatHsYZm6timE2XniqljwZ4GERTR6T0b5eDxbhGUaxQojC
Z8JTVzevsr9Y5izTyXBHmlLlXWCyvZZYJoVmo6TyXz3/sjdMx644PKEGkI+xMoNh
5yVLfBappOcP2qi96JKbuC3Frw3VsCFnImrQZT7RgrdaW7xITKQctKQmQzNfiLn6
QgjWMeXyv+0aBB/WFta/y+9Hk204a9AAtON7j5K11ajRJTBiOdQrWQOymtl2k1SG
Cy5votaDfAsxH7F6fvC0Mm4dl0jEh9NQsqJP4lZ+NaoGAIIycjFc/19PKS6kYabE
Wsx+NkSDNemjOFDljUD0JG84Q4n5cUP2AcEu6S9i3BZ5n1pFKNoX14NgOEIInyiX
v9z1Fo9adSSwk+7qe3veOPJifZbY77SuaTfSK1KK4xmdoraHapmVIEgskqkGvz6t
mgNY5/kwCyIy8flRZKdIaxXSQH3+CkVD0PgS3YoAlqplusjTa+fYkB3GiUsiyUil
17+SCGE+L/ld1Sgnk4uvn+EReJlgtGNwISieYLBWq/Os+jFMqjBUfW6As1XfOVnK
X1ViIavrbEw1uY6WXRPp5U5eEXqoud4kakxruWJnPGM+DMJa4yFANIMthZIFM8I1
EsTrPKa4cTcmoaX+GWBdEFrwK+ByL/GGyGXze+1QOsxJ1mkHpFgmiIpWs7XPlmnx
13a6oHNjwaq8zrWnKKpthwIVOwO1medye4XEb7UaAIzVn5MWAaslP08fwNVidZEg
67+oXkMTqD7KihSFwP9gM4wc7xQL+hqIg8i4EjLg2MCOMeZJb+g+TbiMUHH2RQD2
B4FdWCKxxt2+jwAuubbRZCpI0XOX6y5XejeV7Wy4lgGGxTqdnhj0ohagd+Mq/STb
3gdl9sQXiAKfGU6Xq69Sb86WCHfb7AF9OfmA+mXd+e08GOuFz44inwZDRIPedbpa
7K51+1efS3+fzSrZLa9zOgzQC6bQCkAFJF2IE0A3I5Cv2ozXWj8zBs1r2uUuX1KX
2LTZnGtltYqnWS63VAO+G+7rTX3oorhmq4lRJF4p8DSiYtQ8O1u3PI6hQNEyDykU
bNxpaQRkjmkqCQ/85PBQ10N0ONpDFopL78hwpUPnFIVSZB8etnOrS/DD2IwMy/HZ
NMXpq7wLpoX8EN9OOU7wdQ==
`protect end_protected