`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9776 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
FTGcP7VlpSOhasofAJvqcMnvgHTKGwA2k8ltk9O2uvOhLR68vJn7chtYaENswd5P
tpa7wENf7DezwL72FQKo06lM0HBltAVJhcWwprm2yYEcPTb5SFqqxv/Ea6Thp1Hr
aXn7mVLdsDu7VKvl7ExwJDSzWAaU0anGnAAgHnZvHenG+EhMI0qHAqp32BkU0tQa
JMbPnU9agS1I6Okelg6qsFJl1Qr7GBCcLfXLqXeqWiWN0gkhk3l3QPqxklMiy3GA
ce2P0R6EIH1kiFDrt2qif9X2M6S8FFY3U1zuSz3PH8QUSLzDFUW9/WhUW2fSylqZ
o48HmrUTKcmYvhc6D7glphVeF/It6iq6cGuxJ2CVW/kwrg4p4PP0y4Wz5LGtIgJt
BZcXBMXfN++1gk2Cp/3RXK+xIn8VNM1gWsC0xuFuCACdvtCGlQAFqYvIR2kG6wiO
Z83ZUP0VmczRh7LlTbyMS6GNM2LM1AbIcShEE4NxmK9afPbhlNESm13fZhPNpLui
W/qrGs+HG4weKm4vEhiBlrpuAYgJLuXaD7nVvy8ToQM1oJaS0NuTCopbQum6xIHv
SJyHmYmkwNFPVJs9NyF9kMmrJw+ywvZsmYRCM4rLRUFutfqu2/ZOnG+5LT28mljv
ksQgg33aIDPxWtxi2fLwRRyRQIMgk5H73jOnrD8Morp+T0kl1j2zgbqbJ7fWG1Cu
ZKiBO5ymfyaSGiIPABR58UYHpvUOtAHCzbg1u2OfWlaXvNcHIF8HfgOCU1OWNGKC
0h53FvW2VXnHiUjzGCuvq/C7wm3ztE8N+ol3Th8sVkXhtllwaGdLeeRDekUGXOAO
M+2GpYNTHIS2jVu7afBPF1CB1gfaYt//3b0SOKTXVTFzHo5wvu0KKh0eJRZv6hmc
SePl5on/pT5xnI7hZEA+xe8iTCpMKIaK+3+fgtSm9LTR3E89rzux6fE3PU8csnVJ
lgS+YUyZmiyx01kavbazuxFiWDUgAPQLrJObMCPKbWcLYJBDei36oI2Xel2bteI6
trJ1zG6TfzXFYT3QHFf79QJEw+WurwbxtYAmwRjSWO9nUTvP4pekLV3vqvf9R/20
9EeOfuEK/ykKIXgTBInsJf+ZwGd23xZ+p/LyXCS+FhmZvs3JlVGJ1PAALrvkmGg9
Ijot3p/OQYzmvjvQBEuFCILdDmfdBapzIXDvaR9FQhOlS6kV1l3guO1Xihhu9aaM
V/1rwvMQ8dqmajYgHOYNm1wf9KMN2F5WRcmFLK4nbV+X23HtF/ORMRk25hNT+0yZ
r9gsCa7lTHGTRmIW0XUsygUbixS9tryvBAdA6rpfgG6/Z1eIhOMPADUDQIkQWgvn
I+hGfRfPhgbwFrEOnKvpqhyBCj0V+icKYgPtKLYDClHI8ljffI4BaRF2GxOY29ns
wGeMWHBoQyDIgc0fNUSW8eVCHYsWBjTCuIJ2wcPW4CwDntZlgzgxgFkXZFMBv+lB
J2K9XXC4l4Aik2XHfisBRJ/foR58AO5KB9x8dNm1+Qi8aAG5ONruFH5/pogujT4k
TSOgaNuY6gSu6lAlQiLGZcsXuTV3mgK474O0fJr6uyxSyuAdsDIoH9ksiv+qVKFm
Foogf21sGOJNu40EcU0MZdd5E6jqvI+8ALMnezJpqg2UMwTgkMgJLkFCKVwsZdEF
5ocKnms59Yq8fsbJBEXetgpph2M+YyhSat1ckXaAlU6VeNmEi8VkI6lhkhidsg9I
iunEZrj/16paVM2lr2nYSXoiQcaEILQNzb81Q7iBUaEEkVaaWGZQwepRDPUW5Vb3
Figsg4qSKcGWH4KqXh7m1r2Ew+UOJeUzaMIf/AJWEACQhqSE5Mlra5M+mz94ex9e
C3LEo5vTotuECisbKExtDaJSR4wObYdwpEogUZnchGIxcj1JFoPZhkjLo+jSWqhO
StDL2/KTOuBcUM7G96PD8n0VnaTfFuEvZLv39X6mUG3EnbpEGV81j6NPNsE/3LoS
/MAnB4JheeDga183jS5cSbhdFqhHSedilJiW7EtyM/PWsobwMtsCK9o1TMFR3Rys
lxMI4O1MzYQbEl8s4fNPDZoqAh6OMplDIPBWmoHPXZEMaXX41laRaMElw6/93OFs
dYo73c4KpRIH2PGlIJ1Pjm4MLRdUZfc8wBb344AsWUOBNckR9JS4ltx4YjOVaUwQ
gY1pxZeJqIkHuPF/lUWyHr3LANxz2brwOLWny25BBVReWS0y1wH9wcDcSuOMOMIA
v5ZLFBBBdEENG1jxz5iO6bUnwhrd6Ljm46vjJqfKtsKoNcJEB5Gc1HqZFJ6PiVtG
K23SO6USm7Z2pEiHN8FhSXktVJQXdTjNkHrlBk78gv26HZzgoDgVo/i/8vYxMbYm
6J70ieaV0HiVVPFYB1HNKlISCiMzcJyobwuSdXO6x3PStTlUpbAK+28qvD9ntVx6
KyrF1tjeqGk+dcOjNPLq+ef5SRneFRGhRYA7jOtXHLEe0yB0RFT0c2yS+1tubWth
QpWAXjGN0dJpb4ZscqTQOvEmYb4HvWzmgInchsaK67V+uMit2D3hQj3iZ5gHAqNA
jjm020TRzcVplI+dDDkMKlZfGBcV0On7y1yamG7S2t0F4dyR2S8lNUE+dLuRRXzR
QRMuB+RTpyiKrnggoT5ypBsSHQDtAdXhLBDO5dkAE4Rbe79eoGo4pTr8H7rtC0jJ
iI/7/4//QQJm59BVbJk1+xudqJESRF1kH8i9en1pK5KdLlChgd2k+ABSN4NaYxj/
IMECOnj+bSEtFJ0IkKmgmdNbQ7EU9uU4ShZvA3D+5Rp4nRa3nHHY4EluorfleFHU
KU8M/XQC2Ql0BiYRJKtnjoPS+4Ac7ladpoj7D8GCfsnndwmZOw8UpOPVgZh/dtBc
o6e9H9NWK+WLP+uNFql/RjLQ3Cx4wILmQ9zURpUEnuz8bAtLYwcMY2j+mIxrGNxN
942ltLCo8Nr3g0UgNhTBXuBMduqfHLA1+uqxhVTDh99yF5xj0YHu32xGLYaURgRB
jrQC/OrxwrHFM2ZGr87pnrGBHHoCSMb5yYYyo7m1ISnHkuxAhD2iYd7H5rRZGMjw
AE96BkQ7XB028lQ0yz/jGK1ZPi4wCaXTTiqHORH3exlhIFmpaBTUHNPN05JMEyce
FyQL2AxV6kPcazI/WN6XAKbK6jVKSk1+PqPWbLfIm9TG3jWBd/+hNL0RbZrunzTd
lCb73RxXGxZXV4+LQMKuZJjJRNa0Ufo1Y6o/Lff0QXG6kC/Jfk++JRCjQHl63DrG
iekvIV7YmF/875NtQfw+ZMshjMapamrkaNARjltncPKI8oWpm6zoyZ4jPNL2iYH0
tK+p7XChOhuTEQ5UIZ2ca8Y1oWHaEhpEw19dSzuWHXDMswPXlkDHuqx/+22o6uRN
QACpoq48hWsCEIqHgaZZWTBUVHHoqn8xqJx2MGHB+NjCuG3m85DKD8cGd1LkJwr0
NGfz2O/oEhaP8UWHxqD6TE6f2VHnyfIQz60wWeBSt+h9E4VrstQhVhSMBuQ9gO7X
oKKoZmajXaxq99NSFLI/l6KMCELczPx6vlGZT4lWkrEAyNGN8wXmGUqVdnunfR1Q
5IowDiwKTEns4njdIk9ACxIjjSTrah5dHpJwGvhhhnsOwYG9Uk/1KORA1CINfxZu
jLQZvDvrZilPyJ5Hn+/d9KGHZEMKcwWyECrrxG/nsBPaC+G2Gid8PJncx6eUspFd
nEhSnRY2t33pdmhSThzjJ+I6KYoavJKsgIB5m2q1nZcGMyWNicsL3ObOYKN1vjC8
1qn8Ut2lv3efS9T0p7XyrEDyEIyLdod/9dcOBRF1N15Lbigvc/aFvsaczc2sUeZb
V8k78BQOwi3PLYtaDyi+/4DhAyJTb+AP+jwZHRxZXZOcIdmc+ZzaHEYxqjy4yTD4
VO9MtFIBiJNknXhqapsdmLzFVxmAC6EuX4sO+V521yFKK+o2yaJnG4KBlU5CY0Fh
j9h31GFg+zuzGZIZ4Fz7TpOsMdcRcYTLNwLoMWWOlWBkt3bFApCIi5kyVoew2OPU
4IsSLZtra153W8sENq5zxOfpdOKFhCn3b2FYuQkKOlyF+JYitJhUftNdxHxjrKf3
Qcy9OD83zCD5by31fjwB5kxmiQqPEPxpUx0INfodQNbR5AGOYzGeul+53b5N9meB
5XB2uCFkLEMRAxHk2aEL042ZV6jVq+2qui+O62hzzhZicDo6bwJQSyN37dhe/VIG
zQSSoUofFOzmMwbUZzG3UufrfkpJ8E1ZUx95EQC1PrMmxz8nrwkAkXVaszWpddeM
O5xRMbq1apPMpua4g+gvQJMXrcZrHT38eaEWnFumL2oadCgNhY7kW7XQplUtVSz9
BlX6uHc29L4bA+bAvGe2TXXHNCqwJMjQauhPkF5EirKntj064OXkUUDnooUVgi6F
eCQ7PK1t/HKtkDnWwciKpIDBASEpTHmbramw+B8Sxh5ckRJsS3yjHBpkHTga1pxz
Nc1czE8XO1PN2NJ2SnnHmziMAsVv23l7kuwyqZdzLLDA1FoQCdXZHj9epLjJEsFg
lXxsOcvbqcVBJf0K0rxtFwjTs0mX8VUu/xcbrsnx8GqpfNngabTUEtmUX4LP7wmt
gFjUr1lGUHnRc5TfleQJ9e9+QpdTNqrffmMNXfGjBHD8TPbqZEP8LZNcrCyPapwJ
VT6w4vbiNsM7D5syhYkt3A1HJuZLukFpCD/TBbB2VE+t+zZTm+jWu6BsfUnGUKz/
7yNxEeB831i70XRlxKHkB4Sk8cK2WflRpM28bnj6ic+cDi51FGy+zzETTvZbQbC+
s26DgZdSfob5jXIli4pxSCJ82sPoj6LSC4PCHIImLzkNGgKktIKp4gjTOXb/BIrF
chVAFBso4h/inZhxIwpDaBQj7R6dLC3Ur1gfUUhqhUwl74Qlj8MUop+ai6VQHVuZ
PNmArs2R3f7wUdRPMMGXCux7VqB+NGj6KBIewmTWeaHcuSrbnjau3B6U1f+92tRx
9g53JmhOmX755IStbMu/9cctT4MlkgZWRQXbDH7/PCsU/7I5hyPqqepufPc+CSDs
zhwhZIpLze7K2OfrX2Xi2zGg/ZUP3DYM8GzPLmUvFdx/UUWpr3VsJEan3+RwujBF
RUXvM11a3GKcfumb11lpVf65QSuRyg7ZU5QOeL/0zyFvWjG77efZufLUUXCajmV0
4Xn7490PsavmwQo6pLwT3slZwQDVZEvDWx9SH93azAjsAXWAxqzU9P/d1eFGj4ns
6t05O+QQLumP4FWR8odM6mFwv46yBrAly8D/hwBq5YxVGbbo9EbDa43Rr3LFtjmM
hzhNAWaL5eoNngmADhdP5Gm8i6vxU/eS2a6y1LWNeGUlSgpQQQ4vZhDhfWR6KbVS
yJFmMiF6tDF6PmtwWFt+VBFhUyoJv8OIQlFzjq8yf3F7XAosbfwCq4qKTIat0gsM
CT6T96+t2k4jYnD6UhcQrA/lGI4AmzY/ywh8BOZkpOKxDmqileCWX8XoRmfbJ3e8
pYQ3IbyjjYjg8yfIzPF2dGvAmaPc3fhiTGucgaiOy1F7b95p6MoTLnYq4JeDgbRQ
RwLxKeZSo7aYPM+OxPfM4n/IMr2gpG3fxihl1393c+VTzqdclIbJKjPM/9tB89ej
ikYiyZtExH15hbyahCMKHP54zZCAeyXQMhgPropT0JdMRCuG2BZD7Y92gIzQoxBc
IIhwMj3bDW81UHsod1NporzXS+Vkfql+lDBWBKwKqo20JyhMblHUqqkE9yPbjCVw
K5TlDXy74LLKTMTLwnTpvwGB3zBQKwJ+8IEpwlJn/sBhgAt1vjkPwlT0vmLPgAqE
XVMMadCnfx+wi78gOKp4tZpt4S8ZhpGhqiEc7nMMQFFkRsGkZfvalDjbeXfMwVOX
P3qvufcOiz5VfZIaSxLNEkFNyLr+Uo3N9UzFR3ZMPFSH8ObfSj31L6atbkgANvCi
I26I9X0+5GAWqL4TDAdHD1dmeb5pUKx7xOYagJrnvFqty70O90vLumSaiN+RWOW8
vagvrZUvjz3pO00tpxLZdktDTyt7+o7fnKsomsglV7HBee9hN74W31Gj9dL76xRx
KdTKEtPVqJsnNskkqQ4SlLDUeqYi5xhKsvhjcFzpuIhHE5a3TchaLqqMjrgQuYF/
//6DhlwvIRL+io64oQQT02A+jUgI1r3KPuhCxx0AaJnSal4HlvjfnX8wj2/fjE0T
uo/UtUBCpqosTkiolETeAAMUqyvIrcYxDhYV4iB4pGunxtj8WClTACvUnc4xsk2Q
9BhqkwPd7ZfdbLVrh96Nc6201PM0U63rP3WE5/WPofwKah2sx4vrSVkh3yt/WPnP
f3wdHU999HiINR8AC9yyi/Ri2nx4a3OwgAtXdV+2IWKxGxP9baaBzWgFqfAg21bk
/GI2cx4IPw7YvUA0SQmtZCh22vojZKDsSJDdkc9uqFDtWXZe4P+jLe/B1Rzpq6q7
6hVoO2y+VzoqtmbH8k0TePDUi940Qecgo+uep4eRC2lG2TJrM9OpNW+68o6yRohq
2P9HSPDsTbDXzJu9tsALH7hkLXq5RqfdH+7EEVHKIxo0fDWw/pbZho6kHVAVDaef
Iym4Y4ViuQTo1wx93M29OPbB33Ix3lwP7Va6BDUmrYeoudBUybab8Taicpi2zHA5
vG4nwQM1tUzSvr9CI/KBfBAGN1aS+S1G7mQrYJ8l3msh2Hn95WIJpUNe/UhwlZAo
wV6X+9C6NaVllPACqlH8KXE9w2H8oDbz6MmHk8dh/4Zg7LvDmGTg8KX1TtEyuryM
Fcx+ASMyd2ZB5MvUI+my51HEP/V+AhwXhhNKzc3ZVhQx9Xzz0flD/sutGbW2tAi8
pGgFr/Pz1kJODPfr6uPd2JC+PuRJsOFR0OZYuERCD+4t+RKA19haTIMUVG8VtJbA
6wQGnQFv+uJpKP/BNgZ/ruBT25Xvr7eGxEPwJzg1sHcM08i4ik/hxBtu96RIlUOL
BbqiDunyUiqj45bGELLvlyLYffM+U0J8QLxI+uPCLYWgxWUyo9GTu9If7QTYrWGo
8JkuIk47U2sYNnEs0Ag7QwWyGun4yoSByI1khc6DzxUwXmS3gId6el8m5xbP0pZh
Udbi9FFZE85Pc57/PHW6A6e5VhCRUV5k3OOmXl/POVf7DNfLek6zmWGydteoy8LK
r8Mwu8kcuUPCINvoGVAjgB29q96Dk41SplZ7Gil3XoTj5oCrr0Rnbp/R70VPPryG
Y0KThfBRtLiW4i+Ty7SVBoEYMN50MXKLypQmPIblWizkUizIkV1cyNkNYAyM+SXJ
bfsf3gCJkeUhnQqillC/uOuL4usdbhVfnoJpJQnlOtU9thKAv2VWBoJmXxOt49pf
8a517pMOGQWLVsCPsw3n5bLxZ2UXMMHT5WATSHMi6WX/rMDczur7AJ8vuNPisrqk
oAcelaw7xii9wbJudFw4sCKUTJUpUI8A3+Y1Fam/PHmv8nVYvPX2DoHmMstE6hJJ
CHjbiXVFI5A+0kpOH83LOZJ5cdCG1FJ0mvHp33X82Y4gGU7anlXz3P0At/jdbYYE
aB6PRMzLP9sedwhI25vY18k1eOw2TFtI9qIUX4fIOGFAAZNnumTVzTg0QGjmnloQ
mA4QQE3jku+u4OuSWW/4vjqpHgi94fyQBKyW4f62pa3GMq7vSQ3LsDgegjZS30Q3
sqrldPnvl97gUiDliQF8B1fMJJN7FTn4yNU95kFr1Rshs6RmHhNOMty/K1hcpikO
SnV+maaRpvpRqYFyoGGn57iFWzweUua1Zf+Ylk7pr9WV5q4LV922TDn1sJi9VkQD
fNZNzpIlaX8hBnQ2IOphP+nGRjW68aniY4QJPmewW3AQxaGCENV7WSy359XfxYjA
bg6m2ffS0JWVT/WCvWXMPQLloD+IS/Aw8PQe45wXI6L4R02aKQl/yRlWmEzbfEXg
FkM/tjyqpnUc/tB2daX+StwKNOCDhr3uptNpfi9AolNbngEiXqhYsMOFO7cSthIo
fnjsuUc5qIQUVFgdtuQ1f1jv516nkpKeVUiEwidVdx0V+5fNdNOY4M6wOfmUPEpn
ZSAt6XBI1u0APwcQWYafQtb6ZQgO5aek2BlTtln0qAu/yO741a/hgZmNbd8dlPys
g07z1PHq5iiGk3Yj87d9kKXjwd2I/V0Vphh2zJjwbOJTLY/zUcCqb7yVuEpRnPOJ
MzuXj+Dpw2Aq1dzrhQIXdVbuNsSlwubUsCRmGXAskDQerBaBXNvT6Yl1sdxxemNQ
z/A6TwVsjPVnMbfMMs08jLq4GsUqZON6ANnOqDwIzN40N2/31kyYyHoXCQPJkYdG
Raf57J30W/rzuXRC3SKziDOqgWgVZujzo1CiheOWTDiArFtH6H93U9l3MhmoaG3g
YDvuBbmvEDs+Dslv9NphcToc1UGqKdTpT9Mu0Ecw09VkbtbKSbnjZCzef4BSiHmr
BPOS5kJ6sFZFWC+qJyRUub0O3k+NRiVJOTihltK/f/+VnBgL+4GmhP5gbqB+gx5s
cPbeVQjYX/ooSiuExuNFVnUFIv6C8/LZpLEOZd1bLHyKlZlTELCl8GgUHGU3sxyp
c3dkttkhHYXyEw/D29AZBmvz9DBgwqSgpVbABKBFfuLyIPh4TwQ4sqbDghRyFRRH
2wBmzFADcyL7wlYDL13r+QX/UX4IvqqcyiyByE6R92ZlVTMdUCfEyCy12OGiB9cU
nlFzr0aqvorEqBN97zr1/uDWFgJzbPwap3bprlHoz6ErDqwzMjerm4OG5ndlV6Hb
bBhNji8zlAywC5B0VLuhF3zeIev9XgCc+A77nzL+Cy98416ObPqcsKtolQbtaTAf
YdVEBBgKu92qPZcQCQXS1yT60U8DgbefVgVOCvXJMt6wXXa6wg/jfJ1UcUCrfwA1
MQkMESIcuC1VNN2PK3AAKIpMgai+L3VhQMM/Z3HBvavzRSwwoNVJ373h+SyofKUb
YHYzGwIkAhN2KaGzze5uV25jEu8w4hxBVEnOGvQVtl7+mqS1lKrEzpS0C9nYOYSF
neT5p4Har7BfBrImp1huDvJq+bb8FIdLA/TcGzPrVm2v6v42bqcrz+YSL1ZqiQR4
vXOpgoHIxFk6FlWbxL/Kb1YcOJKs69fETrJ5ggNgx4vguFQVnAegUDMtP1ddAWgB
0F09GJkqfAabMaOAEAMg1y3dViSc5+dlseGrWulYtmrHtI0UAdSSRsmca509k9Xo
Rz7y9K6y9lssAlB/2ELB4h8Lv+3vwwFRgO9jlMFaHasP9URuzyZJqMSTOIg2b8MS
27MftTMSw8GTqbqo8BH3KuGBGHMz4lY6cYtR10Ik7hLxyqDSzcOcSd4aqew6DH9N
yIYJv5FPEJUZFabTnBiJBe9UHqGtjQuMtGqjz31B0+zWC/W7ZjeaGWHxybwyaiK4
sgMmqy9M6/T3NiEg3Zz5ipdDknnqyF/yIXgb+n+7sehpAaU4IV17AHRA27mbY/E1
7bciIMlU2BNi8vzLDcP24FVm1Jh7yRzUT24OSFLKetMVn8UOVLdCwCZqt5ZR9p/y
dTyf3UtM2nu2TdsTWIR9NvipKZlniMKAvd/G6IUkDGhzvowbFzo9rqhhTv2/3a3h
tIVqSzk+qcPgrfXeoiPnNEL4bMrGHLXnUK0fEwY/kFfPu0eakx1d53MGNQy+ht6B
VtFSSt0AMqFLTanIfrGPmgnSVyp7cQCEenQFDdxJ3cRy9n3LQ77xmFQktJs+nGor
0mLBZujKFR3jxP4AlgecGkt7uv3JVgJBUx3yNC/hX9lI26aqWu5S5qMlpn/H0OUa
YFruCOELYVomfJ1kVvtTtyz0+r9DF8IALSyewWexODk164edJ0iVHzWMT9pUqANf
CEVUrGZABKxXKPyU25seZVv+RhaHecV1urXExqWhkMMqzV+yhNulRX23DccW57Qf
UjSChu2z6wYRsC7AVsEtMTbRWt6b+xF/qMRF0OpQYZ03rcfANd7CuNAZ4WaSvfit
GfWpwaYP0sWgnk9Co1MFWyR3pQsHOBEAEICPDEvtZIswgLJC6/KsGvKUw1qnnTvK
5311pf1yfVK9eY57hMqgju7DNjpdHDFeAoynWCcEj7c7rDSEDKdPsvyQ2BHx5SnN
Xjb6AqdNJ4rHzVobMUEf1u10g62p6rhxfr/17hgDvaRt9v4J9Q1R0BIt+taJjzx0
w2ZRtfhR9JXkLXG8ZQzNnj6hHm0lQogSTlO3WbowfoLIZID4+eqwcjfpS79ApbCV
1ag6RjQQZtMGNbGt1CAgFbN5twHL4oNEbHSEPErfRFWWWZ408SnskMyyJoQr2ZAP
mHpD6NmEuo9JgjOl/Sh6earEomFd8AJZOdHy5KmEAx4SdxnjjTz7smlz7UbA6mDT
wwBsTQ9hP6Z/rdjAYU5+Im/NC1cWpujXKSEU5ier/Yo+Rpdge9hBrNDpmQwqEZJr
nX+893OPRmP+CgrhMXFx/G5RT+sUUN3Q/sjeT4ph+OQIKE0IHfD/ljHK0aqE9kB9
oFQPku7u3BvhXMNMfqHfdGo3Qpz8dcIAtRglPbXiJ5nZZQA+wzDAtNwoDmPGzeEX
JsRM6gOg353BK2RWaUzZ4RpPmq4G9IL+GdB7KsFRplf8TS0kU9H3vf+PB2D8v4t0
QU/n6OdMepKuF1ilF5vEnFE/IUkpn9GUNhqw16FN6r8i7BKDXFoisiWgXYXQ1lI/
8X/kvwV4jmiz/eA0/AS/sPttus0si02Nf+xFabpgCzT2kyPXgNFtpcR8Al8nZq1/
ch77uwkO4hqp+0v3wM2lL4RnIS2ueeGU4R0fY8yOjJoSOCzrKiZUse2jL1t0FH0O
3oLSuYDKbsUwDsmnDhhOhlBJt5o1LMOm+ZSg+DtngboBhuNUv+OcE/1OwgrPPtHy
yt3MI4FyExXJnn/h9jLwVH32cod5ksR0C8f7f7Z8ol97kjPuQDhol9oae4edOAXX
DUXM65uOUddPUjv2eygnPpex7KP7e1qs2j+WG6zYuLDLBA+Y18YxuT3EEXlmkbBu
wHBKwr6LvMqSZ4cP3kElQy42Y+SmAgwgc/6TPST2ij3dysv9nMCjeQN/8O3gbiZp
++RIMsl0QPztSVfhoJL537QferOIt7OGrK01/UBXRz8FNqyb4pExgMavV9PuJIFD
UqBoUM7kne4HeJxey6RlLotDOIucft4Kq0DP2Z5DXqU3pxFPlVgu06+x0DinpXPb
fiYthGHzZE1GU2hlE3rezrJIiP9tOsmAC5MHL0hcZ6NzPdNzHsCAclKPY/ImjzVt
p2AT++9AZ5xnwWMYn+yNx4xY5YYuP1XXE9ntvyCvJ2gpaDkx6+700NkKxSc0QTh3
/oev0/b0C61xL7Z7Jw+uSCVS97F9F/64QqD+cZFv0WYVfiQEe+NVZQRck5OLneDh
m4IN0a1ESPioVDGxUqBEEvERbUvQ6sDBR71+QmSST4rT61cxstNrv6VSEDiiAssX
7wJvfaaXj6geRXec4g8N9UIRdiRXC4OUi2yOQsSHy7gNc6sRnVJ/jqmOAx1hwhuX
8aJ/K55do4CZRksFmzHNrTLv6JXgklySuB4IdLQzhX0lsdyPA5t4+/C7FRNPx3qU
zMYKDxc5aPEZ61t0SJ71jZw8be+UgmWgXJ46EaxgnVRZB6IUC17Jr6Do7rl1fsGQ
gUKHuarS5zc+AWW3feIu4YCR1RcHlDdQ0IK1q9+KCSNaURiR1XwBf/fbn9TxJ2ZA
yN5Lrzydhv7wyV4iH4rMkZXDVXcA7MGj7cGSvBuwtekzJCfZxqjqVCCFPLWwkOpq
Dy0WwyEfblqViaTjRxyhrVtWGL3prI1/gAaiikSwx6Fn0vV9PVdRk5LfOIKBJa44
OF2dnqwZnj0HB459x1t8p5IIgA2gamlOp1yJZk73XJ44rs7/NAjeGyheQAvIEvOF
LYs0iKk7Red3GlGHRJeVhKNPP6Hv2YymQwgRUvrbhozv4vS1Ms6s5jvfmwTy2k20
UesoDCFGSF1uwPZmdlN9TT7xIfBeb4p1rgbJVrhwRmCpHBTXMN/0qE6lvo9h6nGA
75vs04QSmoL1FjNiASiAuaD8UxYMxeGVt3elbZITWmkGwipSC9HC8/Ry6wuA+HML
iB/Id8kqLd8afp43AwzSAvegbDe1Hj//YsuNwIcl5Ws3s92i0kzCeKaQ89zq5pEE
CJjuGM0XVye4VG1w6ccNIHh/JxzA+K7L1KrJtpd5+hjVmPmC/O8lwn1j3hEX2AUZ
CTJoLPpDEdp0xtApQvP7Xem+7+TFspoi/7j4qzQO832mY5MMdqw/frRNjo8j6QvK
iBhHE//llyy47fh2o2yZeUvIqg2uZFvFnZoAor8oiAIdTackWIqHTnKWKWswmCWA
t7+lKGKiRNlVD9QmeAUqaTenQz5BXmuOoq4AJBthoIo8FHzSsqHoTWigeBoPuZro
ig+AcgKwFqFKVhzXsGdLaqIGE9SViCjQR9PBSO+gs89GxFtD6CAC9YUvHgM3iLeJ
ydfBUEquoJSwhzJU8vpAOBIGL4eSh6A7pMTq4BplxOwv+Lq7d6BpSAMN9cX2PKCG
CvrOMZOuozWmLPxnAJ5/h43CsNdaLTMWyfdaKb9y35T96o5BupPgBFyUcYow+u+/
6SOdkH0gY1hgqfvhtrXNp0LQMxGCxnnD7MkeGIrWnpRU1tsvWAiKbWeJ7aJQNgA8
n2jWb3eQSkNOWLOcyCni265BuXfrACSsDYfGFmwP5hdrXyO7I/YteJjLR7i66OfV
HruL44COk8POHCm0JTHkgBQ98RDhu1At00cpLl1LIP1I2bas+7hfydbfl8hS4weI
DLXc050zlO33r8mLs21KzBnbehU/Bi1QKzjfQe1h7FaxIOKA901I2H/7L/bDMQtY
pvq9v/SrevnRLerVD7sdk0koWhP9wA5ksOo+3eQ8D3E=
`protect end_protected