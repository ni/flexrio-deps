`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6848 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpugOI2aylgiaIfwy/uT9JvFMZlI8EUQ5zOxQYIgzaCBiV
0Y+SZwGS7YypsgLmWR5N20YD/NkyneAhxq8JTa0Wb9aqqReU8JzMK2FvrECpT3+b
BB5Ae1s9lOcut5fLX2TOyhXN95rbWaaXGeyf52/STBVbWEJW0DA2R/RkTdaAiR6J
cWg5WNWUcQrlerMMxvRSHSLeZlGKt11Ysxucv4fmTM8ejFyNtG89jFG3gjC6xEUc
nKhFkiXzLg7No6oHPv44NmERncxqsyYlGQh4BNFGwbMrzSyybFkHO6E6t9Uwzvgd
WGwFcWAtpWs8b46j7XqOBuw+AB6Rr1xverSOIaxEGbGWkrKB+hvgTdacjBValtXE
zqHQGxcl9vTn6RhYN/QqLMrlLdqQkUebo8x3xqunTiLyF7BM1oQTGGQIGEk6fhF5
nLS9GdE/HZEJy92JH8pcGwzzSYmq7B5GHfn4NbCQl5oT5UhiEREfH3Bjjm7FpdCV
foFOIZh2YzT7egpLKkiGZMkXWekwe4gTxe/Hy94qAdhfYkWtD6Ty4CXLJkc6qMOV
S9aICRY/2num/B+4rqrCpq9FGUiIB4YJjpFYR+W4vmK2h4d5lmgaUmFW/o3VeS2Z
d5L0nkzrVK8/a59rrB9ynIfRlaK7qtGTC3FsNXcm9I3daFeK6oJtCWLUix/IjvDv
zKn221rSYN6/w5B5NTDnxAd5ymFdHJCKzHekavh9IckIaTLfx5Gxp24StVhrJ13d
vFGgqLEKJ31WSetDqeHJUosbwco9mT5iYiABBdqTL1JTvdO995WWdPkH7C0Gmdrw
z4uxM5Q26khZjN52oR5yBqXSwK9+V5FxkdIq0RF+eu/uWTwl47qMBWFFN0FI/zkS
khu/eHxQ3K54+CKSKhTX1uWpUNQb4m5Dr4Pl/hTdLyUsyg2aa9MngBL2sy/WRktI
los49jVF7E91OzlSTkddxn0uaFTZV2dyllfuFHuZ5SMZSDwM/Qa5cwMHTMQAo6FY
j1ccftqjYa/jq4wTSrWsTdbrzLEjWuoiasYyFEpPAqMB8g/lLhe975EGYcBb0abB
kRRU5nlTMqxMbWDdf8deWa8ByQLLsc0XsclwD7pDREsqoCWtvSxOym0KQMtdh2og
1W5fUooxJhejhdbrsQZp2WCj7yFncucwUHW1k6gL1rwjU5KNvMAhGf34bXYSEaVY
tClC9rm4lHbSXxa7A+BQWfvAEUGcs0/S9r6qAcVwuLfVqf9ITvonGruSOxDRO2G0
DtvVCZiqkN749PFZv9mEAxiDHwiVbdmtwj9DCUq7Z8Vbx65VwZE66wUbfxRhRc9z
QZN0t9BymH+lF67TrIdXzlARkyLX+OBJ1+ikMIedtDfIeF0B9Y6BY6pkUDUFXD+1
UkBtz4hnzq0TcAVzbqoP3wDQ8rv2ZpHvsgpNqqwzyFwLoV9ltWUwY4UuO0mDuEGF
Cjy3juHBOCBXzngMty42qw+D6EDgvFpkDQ5qZIA75fOm5vhWvBJpgHNndUApW1C3
wWfLIvlPxHeCscMRd7mEjOezm46L/8azwsaMILWOVUCuzdOqDO0h1ppARp/+TQCu
l+en6nfJc9yhTUsI9gWiZtvQwus9Eqvq161/UgSlMQgKQIKdW5dNKRtQiCczQZ0n
MdlP0U9FmuGv/h81RMLKSLFU49bpUTdFaFsPkYBONsuvYIbDBPUAV207VX0U8QxQ
2BTy44M/zKvNI28nPsvCt3lwfUNaxE4ueCrDHBAanp/SXtQnocGE5tnpw6jd7d6x
o9cM18vPT48YHO7dJntJ8aJZLaozu3ugwByEJgXceJ+bnlO+CCRIWK7CLlV/+eVP
TtKzV2CqqxcSybk/R2WYTyeUCyPfU3+82DJ+hqDUKD3Sy8CWlfF0rZrydcmtFqiu
r3lD712M4+QY+Cs8HntQ41b2c7SWwVOX2KxvnGnEsIvIsTPP4+Setxx3prn6jAZZ
/zdMSj8KjCWAoOOqiPG+3stlobGtlqcUlruUuI0YQFIMdjGOndnGkwhCUgToIoT+
tGFgtuGpG03+G+eVvCYL2FuxImCojVTZzTyDTwACKyuW4MD5p4FNftKONYBjoW2U
GcZ6RFbD8JSKJPz1SSEK1Inqmvjv5JWPWZIA9lMnW8+g4Knt0vVUBBvjmlm4uSa8
KWqX5agNRU0AksUBRc8q43jpNY9lScQ+gXZbmyxJp3p+6S45Wo9zYE4xkCCCinCa
v37zot9wkxP+w1cO8CTRvp5SX1kO9BVCWzzuK1SNk07ACWy74JmYfqaDw253AHFG
9UwMcVa3z9y+bgz1IjYgU1AIR0ya0PeIUIjJc22loKkR0gUSnT6+M7vZtDed/Ss9
USOarD+aoKgx/38h/i/vj9asC624pcj/qIQyB7ZvJFssfrwClmCXkw1i31Rd7QEU
iIK6mvqRuG6sIf33LF6hMGQjFVxv6qOyhvfdYy1viJ+pBsV+OxGcRIqnF2R1u2/g
UGyix53VrQ9Usc3j6Up/SR76KdxeGfaIPcU01GorRID3IyEambebRZY4aDct8aiB
H6SLbOF0GzI90XIHf2f+F8COeZYGoC/WFfh23PRhCJf4thaVMrVp4r0u3M6O4l31
lBkYcrmoCt2O0pt6cnf9cO6jqN/NoiDr0S74Qhp3kxMXMVTFC7rZHrx4Jq0fEDml
SFpmgI3RjfGIO5879rqf125ZBkD09Xc2iA/5a9yVgYy/4k40M8FJhSSkLXwbeaZp
Z6V54/AqBvihv2Rdp9YRE3LILUxi/v5tYgjSh7V5fKes8petvrowvx2+ZzP57GPY
7XJLSNMN13bgjwWBkubprK88ebjPqAet0soX8GR+Hp1+cOjjHvXlkdUiRoJ7ZUEd
v74UpYeFux1h9kOiSbujGCYsZrFKDPmmSEaXf9eqe4Ac65afjpoYvJKUrnX66HwM
uXJQzIfbhCtN/+y+4jMXVVSYCYPnY8hSI96zwHC2PBcEHgmehITaPdI0fXrGHS3V
WY9TJGC683R7JrJki9/T4Mft7pg82Bw+pC2YzrR4M/5Jx3QlVGCc0d0EGgKH7UoH
QJH0KhPRIG4fjIjJQryvEaB/wO9o1Szom9cnt64ZZ7FgLxFwnDnY92RkqZgmcZN8
XY43j4/psp5lgkVW1nSAfwWsIwiTO0hGIVTQckxyI9gCi/jU71K6ew86eazVGs9i
lu584UYLRND3rEsuxvANmC/P2lXg7hnUM6y8sQRRWLAfcFncX5ASNO47lVVXdcQ5
JfxT+rprKWG9UPBjUfrPO8muHDcbL3RPaxp8ccMiJ31mkpTUKI9DeCKh9hvfCWNK
cNz+lKQcjySUt3ZhM2gQmmEinNc+Fi4h8vgpS89yzLj57zJxptgQtixUsEDlv6pG
1jVPbWpxJ6nXhtx0kgCckQAbxuXFU/uMSQzQ+YuPSpIQxVO/HuQfowldJk18cW7O
VucfDtYMDSLMxGZjMRNSUOoY19XO3VkGTk2oL+Poqxdm/bUTl9NyQt36PuYzcNtK
m6OpWC4YJ19xFDBM8BEWzmwOcJWkQN5OYZl2A3OaI+BnZNGdFfq/JpWYSvCzh8zR
Azycqe6WrNgukDb6znT1TgIRjtRbbIg4+QaCVVXHx2V0s/LiPP9IriVIYKaAnRWU
gQBcX0B7Ap45zejq5pm35uPat4z5GTSov0noIF5s8YcIK4s4g5x5LYbMOvi3eZiJ
QXKbjkDsjYMcc5gfTIX3bxdj5osisJCJ3MVPCeblgnd4F81lTdjgzhrFZPb/R6GI
L8rmVn/MYZBB34uMh4hggYct9Pz3H3c7BbtB5+wMKTBPOUTy8MnO1vZJ/LvURmWj
CUN2r2TSxjVsLKYbRrBzk1iH5avhi4pvHtFAq9KMJDE7qoFdezck/ILUQqCZcNYU
7HVXmvtUl8/DNWiJDQoqiHRHI3NUCf9CS368NG0ToqjGDvb9N430FH+RkaO6Od8S
qEdMp5VgrMWvAzlAl0wEKauAZ4qVy9Jfh8p/DK9QeJUTKxJNl3Fop2P2NRM0fIwl
c+TBXV9sg1abmBIS8KMp56pwbi0ELOPHCtaYN/NPNaLTZP00H+BEh4PRdHH/ZSVi
Xz8XKLA52j8E7bUBJYJK37tp3DWFs61YzhbVhBFa9cxWgqSe7eiXXjL8FbHu1f9+
ytINum08L36/TUlFLqe3k9ygFf6JaofkN3BLSkKOyuTMgXkDtjRDPHFi2NQ2R00r
zlrlf3zq7ghKpEW0tejjWjKekWCAD0DLL3Aws9ZnIezQbWyKRDu94hn1NmUhsaOG
7hmwxPGsGUiQ4adnXkbst3wHevuMzC5RXYsIAIpADnfC60FipdQWFCCCulxjxhuX
j9dGu+T5NEcmlUfLCOH8LmoX78W298Fkbdq/wvi3a21PmYxHXjxp0h+Coox20TNG
1USgBg53mZBjtdpel0dpdZlqu7Jr8Z2qHibWtA/QK4nQtny0gc1t0CpqJuNdg7Ai
ydTmYLc2IK/9+StoZEZRE0B+zByaLFBBShQU7PUFCPiZ/dTlx8ydKloVWiiCjCg6
N1vX13gOeyglfPmr20I3rzCe6Fr/Hdeqdace8gkAFHrB4c7ryyqRNBLmD+RmtmKX
deUWK/6kPXTDmO2KL1Osias34qClxQYBP7c4uwJHp/biRvMxpTQW+k9eraV9ozKw
oeHfu2m6bRuBJnEAUG4ynq5nGgevB8ziLcDLr2RjVQgerBO/0eC89yAMhOnvs6O0
hti0iofVTkvMy/LDRg3JzzfXtgkvCcDBZDonR+iXQndNxK/X9oEcYj/qHWKA4pIH
gxeA1RDJgPS255/UEMtjY2ZBuEONRNgyHCjIx+FqdcqkAN6oH3js5ibKkbdpwKqW
0dNLODQZYbJPCYwt67cN0eQUlhi4v0Oc1r0z07gkHiuFioTrRiOD+FoZlHmlhWlZ
ZSZTZqnXveV8YzQ8v+a0LjVv3KV2/4ZmLkSFK4WXaxYMoTEZ5+JkAsF2oShlS5PV
4LDcGar49DLQGnF18nqZd6gwGUSBIeQBlWMxERCltUcm2szDH0rphsvq+NzYqNNM
BeUo9mjjzXP4lfvgToqYHS5eDqUgx5cbvMYBdr0x55zr5VFqCwRiE8CG2bXWmO5r
9JCE6xX7HgAIs5aH0vrBMzoweh6HmMx4Foo8ssxtys7onJH+b6TT0KQqD7+Ir+2r
fNkdHYKjwJbeYxov05ewMf8G5eDARdnUNOewEitE3IYDmikvCl6mxdmrx4+nSi+L
aK+IsEmSsqkpAigss8AElRTfIRFSjXAm8Us6ZLLqigZlrMpjDFg+ARZQIaf7cIF7
cvdtfY582vmCJez/dPjPX1b+KfZAHT1R4rQu1MwObVNznwBrYwQ8Fai9HL+GR13Z
ekzStt4fkpLEWCaSkq9uzBqo3dAw3F57XCjC6DhAIt4VK+NagFWYYjy+oIoEMZUs
VYrhaQn7YaIL7dBZLlVAif/n1a89FGZqmAJlowsq+umEV0Ly7UgvbQO0wuG3eyYr
+Rji+CBcaPYFm9n5eTDmDEvaWS9eLePunwJT7iv8pdktJjIBlRHY3MadyQfEqS4O
fr47WwPKdlHDwq/luqo7wd6d/jgpArEIVaoQhhA+x2jGWNQW146ZspEGnEWJBTWx
3lpcPE5apuwNYaqse6V/ioruBV6GUQivgW3uNdt54xOSdxf91EWqK/lFwr6el+uS
/9yA4OVp97KCXfY2auh+JbScnH9qiO9KBemHu8eGB7Bq+wPCkBX20lAskh2+sBKn
e88yOl6dpI7wYqIvMxeQITJFEuZQcrfYqALEMQda+O0IurgNuUY1TjOeud66em4I
GVe6WNWVZdKO9bEHwHpq9VGEH4toVpDZgkSvAZ4pAUN/XiLJUdzw1ShhpWUSzgyv
kIfSAl/THES/sJ4YuEPHKSEBV4SYLj091303dUAd2ryKcAtklT4xccP3ocq6ClJz
Zj6pCWGmtrqsxpnulnIhJObpM9zZpM0D80CNf/jV6RVOHjdRNblP9a2f7JN4Eu7p
y4He++J7unfl6ExXePixBV32V4+v2s9F5t2xOU9e/arD3z1SdTneLw+cGiV5/kHO
3NSnsWiU4u71RFHsrD7MZ/FDpuDTyEiRm3SFxW+HR0Se95eaTU98bqV6A1dbB0Fx
LAH3L27MKE9hE9mmzqVzqHSNciSnv9cAgsOsM9NZx51CboHpp9aUah3JzxL7/xNK
qFPWrWmdXdJ3Swyr8JRaUnAIXOgyItDsw+16mUe2ior29E0fHvvccuhtgCXU5sVI
XjhgWDcVJWLpu8Ta0bIpnIJ/r3raVglm/gJJODv51pgFjokoUg6rR8eG5OMIT/+3
UDF3TvjNr3tOpu8vK1zVwEY6rrbzzCT2Kglff00RrYbGBL1V6j/LpqMZXaCO6v3q
khU6h4F/B3+AMG2KbcimuWq8ITzt+5s8+Z4ySe8jbXYTPQX1q2Qe6TRrZK/9B7Je
prpvMEg77P2hyMER/673ChTxnOQM2aVU9f7wf0XnmPfh2BV356hMzwAsykJzOPvk
GwSSc5fcq+3IZmmYMIsoVZtU3TXtiO4oMlP+4oWyRQ+HKCRIHzqyXROZlgK06QmH
p+AKOncyGY/kuJ63WVMokeSm/y93SwFMA8Mp5oCmqQT/TnLs+GfCsrLJ/Sd4hCX2
qzp+5wxuoMT4YCM04XH5hsJur6++R85Iu/kxKfpPhf9+II6GsB2Wk+W4RtQ+xNhS
U70j2z7XuzNNIrKuUaAKP+llHFyXnUSUyKeooMdU5933Jyu2Pow2pAIkl/kvUv3w
Yp0dUNzHtvHcqEjnG9/Ru8Xd+5zlIVRhxj6PdUaZRuniEJGvKI0SsNfBW577ZYj2
ONGtP+2UswrAtEsnLXW57yNplqYhgcswCRR7HBG5PstvdlQaPbvFibNN+ZI4qlf7
SLEiIe4xJcfwW2344PrUy9XvZn3Ii/Y1kZ8iI/8/sv35VUw/lKbdjtz76GsulUkO
GHIrGXowZSMWqi1eeE1XoQYM0y0DwBCQ5/Nft8qBwnMEsq0CkEwR5/QfRG3XTm/C
UckI65iYhu+QXKLbV7Gu1DOI0VSULKLIAkgwcrZZVEIcgGIIKIFEXeVsiFLCxxlr
z87E1Tgivqguye2ENdZ0n0lQDEP3UY4QlGzeuiQr10DrIuq+nrhZC9SlimlO5TlE
29reoa01wXQLtUIkZ4TMfVmkGpAW+UqO/m1Z/wIk8WjgY78rN2z9a4Lz3+9wVloH
mFJhUJ5+LhsF4dX6dobWYW1/7LO1DjlAeWmID1e8FbpYG4vwmVmWkZxmMVmmjP5r
2zVpLv1fn0RVG3u3MI3Eb4n3fL9oGGde0Q4qqrODr5im+kx4mo4PWk/Ks3sWAjjV
3uS64zMwgp2/88MTywWKJwEZe33vAwzTAcQV5qUJKaPDOP+sxEnzO+cWyZX4BToI
pSKxOu4D7z8CpKTphOnLfKaM7lunw1sE8R+hyZYJlw1p7q2GOc/yYbFG8Ecc1PjG
YjTQDwU8aIZo/5M7XDS9aCMw+Z53moYw46AsmqBkHBiesnBG1LyXODO43d2KKXGX
uoHkkVrsvrT+0MlZOccwOCMhd2FICyjiZ5xjGLl+JjoBbSacz8LFQPbb/TCb9AEa
6x68qaK1Tdz3NfUj/9rrQJ+5Sp/JBGHGSrnsyxMB21/vfPj1B/zP8psOURUCkCrG
q9tzPCcQ3/TliFmkh9pYHTff++xbR+/Uj1x8s7hsjSMpPYW9AhSW/5eElrV2F6uN
Wwd8bB1fK1GFSnEfyLnDyeQ+wZlNxNVUZ4mwzwu7oF+RpvjUR10YwNUNsXckVBFW
YKQ55nqmKg4tEkUlhpeWSFyOP4d6bnTVmHodPU2wTVKNvuLT2fgSfn54KurfG+Hl
DXsHCXpl6H0IoB1t0J8a78e20e78KFaR67lxIy0qgeXL0DfgwGigx/+F2HIJ5Gee
bI1deMue1IW/lCqmgjMR+YyQSA7ZwD34zdDaA495HKo+vXRU/O2kocmvoPIUMhD7
FwM6gWrnU/59tAS3nd8T7D2WFHqYLjV+xbKKXRRQw8VXXtDFku3bMCUBF8FDPIMp
Iu9zGdjoA+CRMOyJHqvAM8reWTKcpmn3OTaLghTIP8IgA4B1GkEBB1W+BNQ4sxYD
y5W9xJ6QjqqTzu8oTDQcpq0mt8qk/sUxRlj3yZPo2DBZ2XM3GprfqHY16hvIlY3T
SnBFbeRuLmi9a2qdswMhuutTQMfvAICK6DPdVL3KgipFaVYq5H9BuMh4jeU2IvDR
Khcr30RMBxELXnfazRRpXF1YGmGH1ArITw/KCcLf9FsVggfeOvo/G9YTqI/zTMei
NnAa2djFAxP96MpNpwmbjouZvavsnNTQq46CXzosVT37Qm/v0sB2rf95jNlW3/JG
dyyhdwkFGI0xnSEKiqMq1wlaMNEVf+d/a+3Kr5DXQhkyA4nGRVpFCdWu/EYgv+ZD
2ukeAfDRi2IHQrR9JrmKaGOn7Ikyr4PXGlNdIQFH7+GaC4p2VAXXDOF1cBBf3KUy
eIGLTbSWxYFfjVMAKS6+XnSk0oZXjdUTgYO5wIG/CPBuypuy+X6XoJUiYeI9OwXG
Ti11xqN6PK0TLjI1zXHklvKIkcZFYwH72OpALgJLw60AvRrz9Nr4frLdX9YYP8P/
yC/4S4u0PmbnpbP8ztOxXC//b6+7KjERnxZCV+Zq+CNkphSLrbnzxP3dIpyllFyo
8yB9wbZ4CHkXOgZi8yB81vJjO/X2aTLNMjW8tNLQtB23UYXQzv7BZRdZPKkXLUvJ
1S7nSIxBRL5PuUBuKChhK2DsjIYjvFTNNnx7lfwd+F4W4UjCdeIXU/QBiCvsBJP9
+ti3UnaPJxky07TrdjyfOzVM05LgVENi5R+cJpurAZrQA1yZ1Ho/Djn8NNiOeevi
MpAGlA7t2HsUR4S0Pw7bE+Fdnekk0iteTO2jb1blqPljMOOXf03S4TvrxJfHKo3f
oniO7VpYaUYBgzylmjQsED4adoc1YnRMfBUt1ClJTXQ=
`protect end_protected