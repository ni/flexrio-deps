`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Jm2uGAVYfY7w9Y5qKstopObZuZAEY3b/Io3MSEcWLhjjnKulVhCBBYAEQrAzzGsT
vMbffkdZgjdXQUg8jOLJXSHZ0Dgbnob2vlppjZs3bgyHCF7MoJ35E+LOsaLimUA7
hlqStcK49hR1hdeBPr/OwfT3UeVrRtQyq0eJXQ1UksinX1G9Pz3/CmcGfTZ/C72x
p9icpt0bkY4/1I4GBvNCsA6FFKH947JqH27OPACiQQRW/K7JToQn+1uhWr3LA1od
lbVrWu8PdZi7zW9gK3jiW5GaPjwbYQGqeGFs3bTKBILjb7sYHxfxw7eDLVMAIu5D
W+OTIN4JiHiE1gCnNEvkSQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="pm+c2fYA/4JT1uhlJGVUubML8hZi8lME4xPobg/m8uM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
nBaXksR//iZ9fraC7WMJWWSrjqRXHxmM1Y0+KKN3b10NElDzVNMlR76DLrcnamFd
2n7uzsxWqhhJR5LBl98SXO3Y90J6BMbw+OBG/MFM/zUulxh2Si5YK5G9GCrG9gvZ
5JomxuZFDu9CzlWGTuRUt6FsE4Lr6sOL1P+hraQDpMk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="M8TXDiNa0BVMX1P60yIvW2WA9jKGGy8GtbuPknDnC9I="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
/5TNZvs8Nu0G+mfp7M8H+iVAGG3Mh5DYZ0Gn3rRNhV8b5CcJKgjQajrRoGl/gSxp
rBAhtT8Vd5eelHgtvBjpvFBA/EBUrRH6CG6pqRt9r2qUDt4UernbZbxC3BC14KYF
7oZRrPJAnF1VRQm36Ql889MrNNGAIscEBYeH87yDXl0c668Eswg2HbM5lBJ9cNav
w8ekrulvcOImsET18l/Ssj19Vdr/EeD+RI3HXl+IWwgFmHPnc+z8S8QKAeMwTDGk
d4gbhuEZu+hKeN4SJcOmnSrayOezP4cCMDfd29bVTjOF/f3NHtyNjhn5nHZenXTm
T/egZVcjVeGX+aFjzjX2gWX9cEvnpYoy5UwoeDRQr4XsNEKqP0OAyIP5WozK9WXE
O7JwTyJW07qj7cFcWvneFK3gjM7b6gvUYsTZJCqwp0S+cK/4H9m0XaMeCjDriqDf
3pfkKIF2pU3UFvWKpi9IpctUuIUa5aihAcEUM9sp4j2/15NGFA4oe+6e/3W49cO0
53A80RQdZjm7Eg6MnSH2gQWWK4AVkpgwz7mpQz3xS0DE/V6P2IJaXvv6h81aH4Lx
r+vGJ1YYbjjX0V0OJJHk+KxFlteMPQD+BogbFf+YtqFdPlSxV5Ef+MdpIcwURg8K
wsro9ChmbI1r1oJivc0/+xG9OyplqLP2WwlDUBY+N2s/oKS1mhbH/BBnZ+Y7Sjez
t6aAYXW0q6lW+3rFYvtckdEbPnBVpV8FtVlwYmFHfP4VxRRFixEmvn2vFPObPdLU
B7wUCSQtp428VqRWNB7UNZ5oi6L6twIpmr/bUHMMzHIW3ZHTLTYJ1qM43cIxdnUp
wGcl86GjvQigRAXwlffuwO8BtnugxQ5khzLL9e/zHjF2SgrCBG8uAQtESF0mu3y3
MmDnx9xqm1CTTciWReWqfG3AAGdqK7k5FpLpYvlPGjyKGseyFCsVs24T79DLD4Wf
uZE9tjCCeNR/u+TgpauCIWKW/522osCpnRS2FfcYzKXyT+cCDql85fw0+F05vZTw
Si2CUbghqpmpqkeyaTuaGseZ/E3vL6WCIHeToSSpJpkreYLT3Qlf0FShqr1wu+dE
v+HClg7SvG2AHmkxMyjwytVIbYK4WAjBDQ8iJBh4Ocw1+tXRwhycPko+8SseWkBI
hZs54RRL0OzHtm49ghx9/uCToaf0xj8A4bdDtPGlrvYS+24Few43llP3m7UdKcw0
1EShSxPwLhbj90h+nyfmhcmkAdjdun1mFZssKD8ZcanLRyBNE49iRe+i5WaVFkjL
l6lRep0vQcSoyNo8FcMJvDNp1VBXOmr9nt0ia55KBdzxE/WFm+IUVDMdLE2PET+6
TJo3+SLYBE9TxWVea3UYgA9+lDF7O3Xr5nxhkHoKmqKciPF+VN6RUD6f7F2MRiqg
Iptota38lHhQWZ7NrmNNdxS6M7tSIwrv6zyVw6ikZd8b5P8294lEIwTNg03RnHz9
osL8B/BNJKA1AkPK9wo4aNoXZOC6ASP3Qsan2Ha4RNuL0zTpkLAo21Xl1Ge1YTRq
XO+hZQ3xAhyd2WDICPfKo2cV8Nh9CtuzepEoBhltiiReUWyIL97tsCHiO87k5yAe
Kwhe8g+3r7wj5CY7CdSATJaRsKW+kke8cMJ+gDvzv81O3vxSHW0DgeRjG3XYeSmL
DvlSj/+pZZyFYETBKr1ut3Of1v7mYxQJgy7e9uKbAWA2weO6bxttFUe9i4iIIpRH
h0xUiU8+5Ui2Znni41zcdPONn97J+rfj5hNCOJxQLPmR3TVLieK6PRGngFpLyheN
ai1jJh1G5GbITO39S+Ya3H8iVvwAcAWaJzx42nlgfNVa0PtqTjx3KhV0y+gVuFq1
IQApqMpzuJLHTekGMbx8mZPmuMn5jHtoVcnakF668IftPj1KwFGIeP24MtIwGB4F
qaQBVGFGTigJ1cT0Q1vhUUuTYmLUTuE9+Xqk/B4UM82NAxAnD+5FQDSSjQsCtfbb
YU46OZwF7Z9NUydIWc4ROtmVVpo9ivTHR+afIxKRhzVK8cNKZ85Aq6s43wXeCsHQ
4/fZwTr+IwoVPLR5N9imHgQ4yBd6G1U7MpfO5DWO8Vu5j8KlN1zvRdRodFxa1Kgn
abEhrQ/iedDOEFPcIX/x7LaLR2IPZSD5sVZOZX4qK7X9eQrqbDI+HS2IpcIn4kCS
ejCN7hCOtMVu7ZeBznTTUEAmu+Iqs2usLz400Gxe9oHD0gsSzYthJS18AJEjAyAq
Kle7HGf1M3lIc89Xvra8V2DEfi/NINqXVB2AnKSApB4UbcJx3Nav28XIfDXcKZEz
S2EnCW6/SQ8vbt0dZY7x+QrgzBfKNMkYhFcpDI9GitrliaqNyGIc/v/y6ng0IPK9
7BnOi0FFHir+uXePsCmcO0BTBTw+YuLK05/eDQvXZ9v1/VenJ6ZEBrO1uN6UJ0tq
WrSuzfhZDzxIvqMuPVogHeBlrejsTdArHTUTbwcOBXvcfXD/6+v/nP685CBpkOu1
XewxMw1ZoGXkPKDLBFyFj5XHqPLSho+/ADMvjcfvGWEpBIpThQG7KNlf0vDqtmLu
XAR4qUlttBRRjx6CXnnsRE7rFpqQz+7+NqD9wlsSEEXijnEd0z06DY5DQmkxfHm6
CTJVjniYLpGANW3aBG+4LQOomtWpIYcwJbbhRAhsAfnOXLWQa4HjX0OkA/ZQpnpY
`protect end_protected