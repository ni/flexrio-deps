`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 17440 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIbuvaxEZn5HptvewZy87nWpqS4xYF1fvDTCdnsnixmLFC
mPgeP/Bto9J0Q3ObgRHhHAYdXn25uMFlt1WDSBkPY7uVMkUmkoMJlMhf/0HYMdv7
xk6uu3tg7XX5CczzyPd0uuzkzVxHxDQY0O1JlieOO2EWV0WKnUz99VCrsftKD2Vm
CVBBLSKqIGPgBzOtoNHGfdpNS83Zve9GJGg9vdfApcldp054WRHtpaZ1VKSTpEBP
lsFKLOFpCrTcju9ihakA/2003IyxNYRbXJ6s3FCoqesaJRw9KRFOGE7Tjk2uxQ1s
6GvCf/xbR296E9XfJsuAIT1VDtV+ekOEUOX9E+10JWz8PNozARWDkTu+o1Sz5ND4
51VuQ0NzyQBMjVxQN89vToIpVrorGnHFuk05TaGl2ufmgixTOyAlkxU2+4NFEAn4
chtw4YWt2GKfxncGOWDlCSzxG8JX0G9g1N9ak4Lb/2Dlt0DfD+H16Xs36wQ/6XE7
34fK+nABp3xQHBay6FNRwZBNGovbBFCFOQMkeRebYK100K+mW01w4tYCNmJirT3m
F72MV8t7pmLGlQPyqk3H0tIWwjTH7f+BdulQQrQSr9Q5CQOxkNbmeGiF4ZLgvz+S
Oka/s9UpzMAUPGmKdp19+zoEh6BnQrUhjAyvGsoouSnKMNQYIJhDWazbV5Ywv1Tk
N8j6bVHw+woDaWXkTJjOtsMeBHgs6LR0gTpT7395XJC43b54VseSDuuqe8m/wUPo
1lnVS7GlArotYwkY8P5hZmyZ4CULZ96Q4vvNGVmbVLSy/l657/kOKt9D/krsusCt
OCRyFBLW20lzV0fUVcQXTSjoxVXaMXHrrWBKvMApcCMev66aeuIqwYTu4zB+2G8s
UCC1NYyG/X6oB6YD0OMCxhRbF0/GEGXjdujdnScDrRjo4ROSJt5uHxeeQWfYczzj
bqQDKQJcXHW9YpdP9x3JrSXZlAvcuzZ9jhmQxtsgkP9MpoLyxGfgotUV71AWAXpx
vflMQyPjUpidGKKjWDc9GMIn9vIPbQYADIUfghyOL5ckXhZnPw9J26bezzBQ7/AZ
8+Xu8azfx7cY+l4JbXZBIxkwsxBR07FEjKoaj+BYQeTcuA8FwF4xLqRFfppYg9nT
V/EM7sph0wk/B56YZZOgXQ3vJLeZAr8uOqTSoA3qHD+nbTUlMrgO1CF20n7/qnrX
SIPGZr6GLYFz8/FJ7YCLGdnnH97eFMW/Z9txExq56MYQYHyafx+tEhdggyxVtqgO
2x6X9qiowUqMKfOxITe9cVL/DyslaxWctBJi6YLXk33FxBuTbyVS6HdOO2sWEsbn
Se76VOmFDKhO7Ohunefrlia6J+ncBd7194ZE+HK9/VhWvXxDAMV7fUmO0q8uCLJ7
rlFdi4Tzl0Xd7FC8No0mHHiuRRLddCbZq2bDaOVc8WaEyvUPZwkQRng1ii2yaLwY
K+hbkP+fMCQb4yfbJ1+lsMf+0n+wgi9Pmoq4bOEGBOhLMvqfyQMKb8rPpEWaKFAG
S2MGX5OAHNutZ2z85OG4N+FYD96HRgJ5J4wgQlfDqCdocJbka7aorUe8zqnYbrpy
zxbtan0wzWEEOKFYXXL8leIwj/pbp87YgtcmWs7Ompf9Gtu5JRm1S7qWo5ek66mV
ZzMdBDRVAjQ7zq4u/eV+qsGK/ILZDEa08DuW5aq2M2fqiHQNIimpLU8rVELzR7hK
Q/V3+JLewTc8X4XEZ2LBb2PAydwXz45iQ/LpEy9HQ8wG8Qy1WrLLRGUzxs2FEZxS
RsNti7LWOtk7GB+lKLEJzhJuiuKvvBOMmoRihiE7L0xkqIO19W4zRHo7XcMZPIm7
Oag4vF7drFbTF6r29G2oei5YD9D43FN3XoFpL7nPAuLWcJEsmRirbKUb143GSUrv
qnbCdU80SrQh0X9szurCaT23peyi8pqu2riU6+BCft64ANE/VD6jc5zYWL2RRDvM
4IxFgN7mzxhIE2tOhqvwAbF0w3GbEwQ3XPYmeCKz/7GyK2aszCHM9z4WuutTAKel
c5d9d2Le2T/ggGaiGPvWbavGO/WfX7q8xFvkBHqfYFrb6PzZmLyou+qKGxpHRp16
I1fu0AG7KB5dc19t+pOP/HIUQ6O8fV+lUzW2DvK+7VjDTB7LhgwgRDxgkfneyLPj
G1Y5z5UEBizrF9PMQk7rHPfMW/ECJ80lq85nD7xr1kQ/fUUWSFY7JfagFVE8I+p0
06LtlA7Aeyu/FtLHEuMrzCCUvRXqDKZZyGcfm9O9yYFM6MeIiNC4OwgQh1sXjhED
Rwa8oIGpU0Ohvgq8dyXn8EaekUKK+wsYzWSq8z+ACEKfaAJ0JEyFRtgEf1S4uFMP
W/BemUrvUj4sxtvzeo6Wmh++Q33XPa7kymjXFjScB2KIeTCZTFFQcvmSklBTcxjO
XCzQFJuSJFOcSuHlErvzhhjfcWoWwQyihKgQdglVQdL+82w6GD1WvWkSSwF/OaSi
xrZS9ivewgpLkje2JoLBy/JirxGWC6RVh43fXDyOhKvjJDRXyI4hlJVrBwYDeH98
1NXyLl9JVNdu8RzTIRzLQ5OekpIiog8QnDSkaFSaMEog5/MDXKLmlJnOdBY5KONM
mAzrtXlwmiMowfofHjY0jOO8P8SAArcAVTm/tu7wdv31AOjNvpsmcV5vpEwmMO7F
2uI9W26n03r5CXmtK6cNtXBG0OnR32KMrjJ/UUmh1AFerT1DRODzZIDtehbfVE36
E++oWoX5xTxt2vSxHS0oK61hBqZuZ8D7Kh/76CPoUxOb1/h+8P5m5xLTqzVeCaPE
NhNWxSMxzy7uHIMGsJuI0zs34YvXjiDZGhYyPVVpQ4XnYVglhr2uGMM9ushplE0s
xmqj4w8czbjlo6za1wLK13O/R/rrYz6VsiUjeQlinEqFOSHIGSgqWRvfk9JaxeJX
yw5GZLRbb3rISAoTReyn/eLBUerAeqQGK3QOqVl0oR4/l+TUvOWotZwgQcoeitJ0
/E82VgRP7ZjCOuaY5dV08XF4wa974uusGo1/HZacDzunbSe0Q2SEt8Qj/2D0/PPr
zeUyBHGvK8T/qqcZXmcir0aadYMrjstt5kmohaiNaxBvarl81cngSXR57ymaYt1D
sN2ubeIKPNqgs3VOvyOoAPUpUjSSXEhkiOQFdhCZ/yd93sQO8DgG7Vsk8y+EkS75
ZUVqp/zdeHVh1MdpNPfsg5di3TxekgaR2xK9RHvkNe6p81D0VzLBy388/BYyS5DN
CfU2bpjVy/KF66moCvRx4mKOThUzjSvxyIyvbWqaax25d8taNZXyZGn4mG4u23AC
JaJYO6RoKypxoTraNRLF4HIRGmteTsdPgBQykUlL0ME+urBY0jktPKSyjoCSgR/C
R0PPAdHujIzHUKKFokNjOUL5IArIPD8Ej4pnojolTIKyKx4rgxVn/K2IOa8Ifzih
UMCkFYIi1tHz3ODf+rBbT9Lp61ns+1HHjE6mWO+VyrmiZp22IwGB9IYHDz+uYnIQ
sBnFPgWUqvqHuAwCbn/aMqGNzunBJabifzQWh4oO40LoIGScpRc5HWVNOfNPMDfV
VIdyOn49ZyTTn/0UCuTKXezeXbzyfjg7H6cn8AXtsCwAtY8jE3eSOcDi8p0lfp+s
WiLttPNIbsWi52gLWs/WcaVAmHL44+kSYfcBveCx6tQypVvUDLYmeKaxN81PEJmM
H3Ia9Ulbue6DO3hSJSeuaLn0m5/WYSa09FrCtcAcrqfqESeyKU4CcItiDtcb+zzr
g1n90KQaFZDTLjtju98NW+LLFafs1YKonfpm9QWkpMR9stta15jrpxrbpIwQUsTQ
IexxI4Spq1vD6+Y6NMseZFTvnD9wyhWEWp7RXKzRWtzCcy0PQbMALToKBJxDjgwg
l8+rokn7SWlx2/EDZvUqQKfhtmusuj6axG7bhhHCI7qZxJDFLgmNClddj63I2Mnc
7pUIliZ7HkEJk6icTqfhti8peTqKB2nYnQlSuKuj+qGQWcrbAJ7pGIdNQhu9FOZC
SJiBUEwpzsHbWqg6WszJmMzeFUp6LVRBBgmZEzjkSrXCx2LIdEiOzD38iLDua8zZ
ZrQWqoL2+LDDky8zjayYlPME5fuMULBWrExELkos6ZS++S/eBUQzbbc1cxR5zWT8
m2rVjaZgBtpDsKPPGm6XFZMs2jt4+4w1bTGwL68oJbCj7Sxs3sNo/yCy/wpD+Fsy
Ifo5JJitEETMPpRliQ/FvhcGZjp3QF/8kliHwAQiYNDfhEJMbIEZ4hsYQbkQY2iW
iQTeKbrxKawhjb4bJJh065e5Fopzq146vrENNRZqCa0p5Y6HPeuS74XTis1PBDkq
j1vSTmEZPMjsz1IGQRfz+S2rLEkAYOkDthtR7hbd5vCnuwc437DYq4rTnjArLSIV
qSmYLLgc1kS0aob9EITx44mCGojGB8z8hL15MzeehBIYQ2Ul+Fdgscybdzfalcna
5iwm5kxK/a9iYV5BwHwPrFaTmINYwNihMa7xouzT6d11I3J8nVBEf9go5PpSeINw
/RhQ2efsL1/L7ziZZkxruCU74uWMXxmcnwofgBFNlpao7DNKYZd53PKUbYC8mm2k
3TcabOA6DcmwOrXXsP4gtPi96B/eM+XEuPjs9pEjMnJlj0/OaBBdOY3F/9GU2pmL
43yyq1C7KaXfU70sQgECh0EXoe+NHIQ7e74bJPYWzjoDx9Gg0ozwzsfneEes/tS0
b0vZhu3e8fUbK+OlX8V3FOuVMlyRwbf3517EYzQxHdM7UWbBm3K7AW04QJ8Nj9wN
aBJ9iAIRZnPqL78bvVObPqNojdMMGh/oPIdaGZejUy943ygFkZEboxXvdN23gOe1
Lrx5uVdSiFeqiTsLXYIQFRxj/6HH0HZNqJqpM9mWsmdLie5yI/+RIbO8rLHvKsby
/N4AgYvnMkUX8f0SF5OOU5LZ2eVMT3iRbH1aTbWX7q6seEdeO4Ofl0vyTe4C4LrZ
2vEjpapt1vxoUE+sfLbgboKybjikn5cfLfqvb3bk9Y6gcCmXIyjIIjS3Kh8vHnGa
uf4u47ZusMs4z+PbffEB4WQ+trE8BON/AhiWKH6nZoly5lHo+CV4UPruGlpSyDdO
xFvEjv7LMwzJR55C2Xzh2rjhq12SGiT/v/ST7oBCAPiY1e/WXRfH4w/unARJTUtG
r9XqeqvkEPSRAiVsDPqOIfqxsdg6u6TpgPqAf89QZ/QYJk1kHNi4stPGQmT0srXT
CKrckYkrO4bkcQpcsa8r3jGHvPop61DsppgpKwv3CS3NHd9z4hdswrjW0PknJ6Cf
Os2NP6Ry3vl1WSGKkl5L6DRLEYvKm+Z5OK0eftktOBj8/ymA2HSGUichOBBQZoYV
F7OtRnuMEH06ZrGxCAZYW8v5WYQuab+ULGhq7ho1sszXohv+P5oxjapKgwUBlu1g
gzTDPyUJfikbTL/+zX+XlsLcrGVd8UUtkipYbxo7X8bnPwf8B9aWF5H0BzpR1Pqr
Wkg9buGDFd79xfbK8nTHTqJOmm4inqs8rnrBTxhIxCE/URN6W7lubGvosxZaYzgx
cIJQY93u4Knn0dfDgCx9fqxhXV8+zTfN5Ok8LSHaPovXYa1Gf8a56WtVl/e6w2rh
rHirQwqZybYRB9KnbX8kTCNbeELrlr6D3KKgQ9d+i2N2QveS4ITeCzAUgX6C3con
ttPE5nwr3ZPwyybLc3rYTO5eeag40CVVf7TTABEx98ClVSnmHVxmJ5vEeU12CRri
vD2K3dN3QJUD5w+HPpcVCgLc8TOYKQU4WlhK2QyiZO3RwKqRTxr2vV1IRLIgnj7p
rXy4JuZH7gTaOzknS1/I1LwxRWyaZx21lrUIIsgiacKmHrT2tqymjJZXoBPZr4BM
lXGoBpEeUOupw4hmOwO9vyDl1KKp/ZFTQQKYK828mmJxedhU6FLymgDedy2/t5yo
jiAJ00WumNdhuQFZ3TWidFUCkdvZLMxF2JDpA0o3aoQ5ZN1Agmss58BbJOW15YMt
JEe3lhvnvX6sGI/Yj71R7K3ELMM2biZFKyeQ8ZJQLhqKfx7XoE7GHZwD2kHz6G9f
dLGFQNG/rHokOe42LOIt+YPNAWwXbSXPGxp7eqmTAJrotneWyo/p85yZ6s59/bQR
tKxLY5gAGdEA4l7pUhB/FlNN55ROFkGiaZYjm5K72FOdtDedEgfiC4ZIftzssq6n
frLcm++UdTQ+jbhXjkPme0TkqJLwfWd1126AVKcGi1WRJ9i06AeNzv+jvegquz2t
fVRQgjvcULB3hP082jQOltVHh56SOkcPJOhMbfAFOxcJ/qFCj6F3bGx1IavTmpZz
b77IslvYNQRGyqm0fzm5C/BgVae+FQEb5qnWuwV9S+wICwGZAHAOIXsHS/WntI/J
xaCi21XqqLlYYYBZJuCIYxS8sibO/PXM+UN1LSS8CXVvfPGgUTte9hbrTGSxxZoy
eW02m3KeQcfpdzXqawz+MzbMEkvsUr/iNUnswPpivdg6N0GDAIRFmDaiUwrecOa6
CJl2UnH9pqK57ynWo0JRB+s34lLuQrkPxXkl3GTV8tE2FRMhbcotTYlnwqN50jLE
fmuRHf5I0CP4DFS4SS8SeLkKifVrWwSB0hE6bWoIu2ayiW7JKhOOXDWOFJEys1ZN
x5oRtjH9P4QBJdwsw9Fql7Q8XnQHHWGl1kT+ieA+LY7nLh/K1+QVQ0iSHjldbWgI
KEi75ZoY4ZnKPID+l+rXhcRafsrUEtDBh1fedHyxZptcCGVfvfzznCMKP8gtV+fy
j11zGVa0cSP69nCOxfBTUR0NombRS1LDYJx+IRH7TXSjenN7CDjZ8qiUetfF+IJG
PtVexzHwR63XUutPc1mdpHGZyWRm31gl80rOvTZWgJR1lxcJYu3dSCOooQ+l9kqR
dx3rZ2N5K0h0nSthaAIMiXj/Sa8VMa9oc3IKU8IKVZ6dkXGQQjjfaM5/MpP9wNFb
BWpeC9RbqOBZya4Fj2T7b2S6BAiNZdWQxjzG/dTXvWXZ6nBcbO5AxUApV8Od/OUq
Xmx25eppx0YnOhs1ahg48xWgxVdnoHWKW9rSeH/yVKsRU+WhAIARE07ul05HJ39a
UlWhHxO7hkP+R73Qq5Vxb0eAbpo+fIx2yFYC36YCSlneMzSCsxIsw6m3EulBJ7Xo
4LBkCYUirtORVhPuuTI5wiM8uVgSwFUcbrvsCVibpGCOR05NcO/BRe7Nkh3w/N5Z
O1NxSLCnHPOtAyfnfNYuQ9LcZDP5pGWEiGSXVE7/nRAxrVvO05BswYHRVZrc+TYZ
F6pGatV1XD6KQr1TE3r4j6BaLl4EyffMuSTHGS4/mlbKFVjlaf/72k/mKHrLHE0W
hC0RTcGVpPM9+EAC1Ezngj7uBshtH12yxmSbDIVZjTr1riWsI6q9bqD4zsXkVSv5
GLe3LvnPRDuRCxsWjoLXMgn5oghTq8EPayFjmIQ1ok+zPaRuBuY2q2YikK4o2NCL
z8tqP0WKCXsSRLhn8Mp5xo+zoLYtTMeeabkhu9ewWIOrvutlLkHNAZLrdY/yuqSr
v1phxSik0zVMtDt0SM9oKxnmrmpk4sP8NvSmSmWt+oKn/QZTCM8SoxtaTzaWbEgu
FZUiHeRD01Yz7IRyFa8qL6u2yZ3fwRPVdObGgBa5iyg2xGt0MxNbtQzIggeYbvyR
of4JLOumiUZTHwuzgptWcHAFPHBXCdYjD1Xo9lJ+PxkvKBFxurd+AeGlIKzR2n2o
1yp4R+rGqB8z6Tfh/HqnhvLgbae+zdfX4hIw8VNIOaaVG26jvCQGkV7cwpxYEyRZ
tkThaNgztmfVIhuRPxpebPcCe1Ng19pTXKNHO8I3olwrsLbA5s295G/Bu7cLmwjb
adnJhcKmyfbu1exSqj6MnxoFtV6uPD4gNVLpTMWQoe/9A6613/nSetD4t3427aiG
LRf++ginc7On3B4PklKZhBP+XPbasKyTdzGfJSsQVc8khSYID9I/NAYvzaNN9VCb
gdIw/2lsV6W6t4paKb2I5I8sZ2TSvUTWVn4awGirOsxmFEMGz5dIUsw4qpTYyRB0
PHO36HzW0pPqiw9/ms+saD3QUA84N7VRzeWVG6n3HaOPg0e3gJx13Aycy0n7S6pi
fKaLAD8qW3H9duMJJoCNHpuHKQqVZC076kbgRVVTDYTsrTUWitnIrLmqmsgYxfbw
shjSrr7mEiqmIRi80PU2ad40CKur7ob8erZJ1VmeZ96pPPyv0RPXYw2PjIISGPCf
UpDnkPlAOI9mhbe9lg5er7jzDSjKCnTIWfEeksWeiayiMvvfoN42KtW285fg8FRQ
aCYZdErwyqzeGAkEZf+tOYW2OWJm10eWY2or+k2sthmYYsv1oNRxAOd1bf6PMtan
XPVW9bvj+ZfRm+PtkiaE1gvDSV6G5fZoHOh4OuhBSQeqwqWLs/pX0WkrF/kpIfsA
7WimSLsKIWnkY1VkEkvSHHOxjM9SV8YMlOmVk+epMDIchhBBmsMje3E2GgozIrJR
urdSUWicpaSyHUVSGRuI3mV+nRflj7IV7InvVEu0OeKLCHNuGRduWrd3rnIe9KEp
UY4t3xc6r4Lh5ktKFvHprmb+f00Encrjd/2vMl15axxNoJ6hSXh1uPv46rMx7f0l
9bdCY4bbMIon62wPAdlQ9z3pZkvf/kcbSsz/zumISpxRJeSfKUjGdcroLK2XHwae
ujSKqLZb4/VMCbFpzzhXCnDvIUVrOMqsOLafzNPHAzzdOF/QuirXyhAUYu1KjV56
q6kvplBYl7+zXmpWmtnsGQc9Tsx0wf9YUNM6fwQRlgWhyf4dvOPBY+RayXjwczFG
8myytI8MQmS4VEnaoPfMcB2GsdS1SICeEOzSzyADmD7IK9zLAIH1n+t/g9E/NqdI
FfwJ0j9wS+Fq45+u2hO6glAUypfDIasEC4GqcmpbvtWoGjnLKAmmG8Gzmymqyjrq
XVY5/Muqpm39kpvkB+P/GFQ7MoXBc9GdN4JALUqCwKdjkRbfpcWWmYRUhNO6bQCs
pXfKhWCSinR6/tLYhp15fwbgF0YEli3VisSBNIMWdfNtKZPYP1wSn3h68PmeZh/Z
CZnl+vaJ5eCtWw4qfZt+c1m5fIj29e1V/6cMW5bAvl9ob/aagTeR1ArpmGqLzU22
mxB7ZnnEFi16/WM8T8ljKosI07GDb5ZzozXFkioDVIAzig6ssuxFl+z07+dDWVE6
/Ghpmq6GqFQS2sFmWkLNEkfQVByT1wUYb0sArQeWSZTFxLZj5bhi7xpK1mXzPNgV
8qAfXkmJoj9U/F9uaUE4AAnXKvGEk0ct2RRoBB5daOXLmzGQbZ4RCWYBUxqZkeIe
0aQnSDSj9ae+8QvZ2VSCIDBmKf708O5Q/q9/JK4HYfvk4biSnum4mP3mFdX/4YDh
5Va8Qzp7Gb7ZVHCmK20TUq9eF8f1GWrUNvHxWd9mNzSYUC921LAysOE11eiyrn9h
K9yiJ1EMEUHQrg+mAJFYQCtRwBKUfYsebM4fGfnzPyC24COWfwk8PfidAXd8T0Ya
BZosR98eXuSSWwXYm33jZA9C0T+5ExKJnB2xNZXOQr67qFaZz0vq9CjrF5pZP6lV
IN13Zh3al0WjvQyOPUGOrlV/q611lmvFpcQlNSvBlOH8MHBZapKGEc/L92rAZonL
CCjhVUGaVr4g1o8r0RBphYE5h6QMBQu2t22YfMbGlAQIQYhxDXCbT6jKTBKI11zk
rOGkZSMnnp6bp9QVjDAqfv/PzM817kuE38CgKydsubuO2ZiJVC5NMfrJeYwY72hs
Q5RxYDQG+rel/+fYTYT6v7RpepZ9ygoBubzLKPkBsIxtxZQ7tb4pz0gz9WDtjGF8
azJIDtlzyz35bXqjUvmyrDuTXpSIwnmWKpr3DQuj0XmVBuRFXymstykPBBYuK4qi
HUPqWwJiiO3TAhkNo/P+3bmUNmm6LuGZETDyC+9OtlI9uNSFCyAfkkbyFnI0VGP0
w/MAhQbR1F7QpkUf1ZaQjdLZp9sUnuyefwPoRtBnhbRNh33Llt8roLRT+2i4R60c
qTtEBS3FZ34/WYNyBKHNPWieVxjmrflV2MtwN63wQ3Yday9TwY9mHXvrn8IPhN6F
lzgwVn1q55MajznjkRWaKnZu7ZeHCOE0EUrDQgmG3UtjIj48oe3pNXLVGWWmAdr8
TRLMDkjGeKHgLDrQVZlSKHyQtBtVqiCZFnNFK3tey4iHI8HntH6vi0J5FcAhNDIL
jnM6PfkC2yPZWTZMRRdO20An59cQ2Bjezhyru8KZIlw/3LOidRw0AVGfeMN6SD7N
ZAJQrwS1qxjc4dDGbcx+PTCucwd6KjxA4Eh/xn0hM7xAwlh6IkXjoPJY6WqKJg6D
M3n3v9TcxtAPJ6KXQZrD0b/usycZM7WiUaU2vkVmatle6+iDl7vDYRVQmgJA/3DF
leT6FAIaIZfBXcknQYywwrOWAMrwJUU2LmPE4/yRPR6UT4Pz2B1i6KX4i5hDXmFF
vr+TWFQIwplFHBENPaByWFq9aTejdGwUbznOOxxRRUideJFoM4VL3O7Fv9z7i3st
ZLW/vcUha7HP5smJrQ9HgiM8jiRkCF8ksGpEleWwWVIvTuQDPxYwdyfRXfml4QcT
vA1NWRzMbeNAScJlE5l4NyH8ye2rOegXlbl/b1heX08V9ldZb+knIfYrvQcDV5yK
Pqbx1nR7nSdS/yqeXaUDLp6sX9XNjQZEXvjoxKfkQtuBPO8m+ig8CfHQ+XmGhZwf
KAaHstI3a4wHQOajnjVSov6usMDPqgfP0GAjbX9dtf4Bcq4JaNMlI1P/XkQR2aSC
uI2O7svcQMpWrum8rqr+HT4OAcVgzygbB1J7mU3VekwPcTF9ZV8WADtScVbmgJP8
lR2d7F9eG26ROvrK/ZtX0mAYQbS6R9AoZgE6tjRO9PwdkfS+vMvPdjeDC5Ax1U/v
NVVjLo2icn++rQ4FJD3Yyg/BDSx+1Jc56DUH4WUGWtrgF4Z2Ou6w5S0D9fkG+DIM
SxPZiqd7icm2LN0n4nSp4mqGgL4lvHYa7wXeB51lMc7Jyaw99yKCTC3FBgHfjtHK
X97qSQ5HjAdUdf9q3SZdN9iWPBtsnsRVmd4dmzDQKkTpTekhm0waQur7K21CNdq2
qoqH0QVO+O5oyIyvoF40QK+cz1b2XHM1OWCL7GbE1GWBjVe7NTxc3gRqIIGB60VZ
TE7SN5qNz8i+EJwdR/OU+0MGgaR1/jg0TMcF3ihBsibh3UVThEyskgfftAeTk8pU
sMqS+zoVKj6dPhJi3xL/KHYwmENWcqOrsdg7wn/R1jll73cIeuyfR3QSGKMx0dSS
kbx7AkK/dEjuEfaeGAqIKLrmBXcIeOzjWJVrWyePUNbjIYlui03XCVhjPk4mVQHh
p6ZtL9MrufNKyUK4WYRgACbFslTkU+TsbFmw2mF2JUum8v1KHJGCh2JMdkl+S+Nx
4mmcIL4HY8977pakx8/56WVgakZTEoYeRRZ3OKvRrRY8yRUE4XlR1wCE3wABxape
w6QYkJ+29PCv6LMz1Am9rI32lN0/QC/GjdHPpGD+jLaj7WbrJ/DqdfmGT/QbZlDa
T+tihxqgiS6BFKhYyy7frSqUPRBflNIcxouvOK8KSH1tLuf0OIaZcOOsCDJHgSKh
uDcd+hLtu8IEhIJp/49pRGw9UhTs4c8d437SNG4DmtxKvIaukPIdzd+LotgWfsIc
yfo2vwUaidC7nImZueAlRejjc/uxLa8SsOkQGiwPsap2W7Mw28VbKvhWSIJkT/VT
qNjCsYkZ5cupEJ3YOqMJsDqGyKuNE0IQ2OHhCDUqi3oupAMwid6UVe6FVqV/uYvp
keMICjG/2EL7QMJAJM0PpVbej46UEcdY86v3zf4xMttEjpvRLU/E+Gj3GEBxaNpV
Zk/wRXY3je835ODdQFHdF1Mha3nYo0ntTU0xbOtBN+ml0fsE/G4BScmmDJl4kDXZ
64oECVxWyfPkAZOOBRkSDqJFrB+5dCeE59V1gxlp12o+Ytu16mw0LgaCHLOiwsMO
A8V0opzvydwNYBeOCBy+9rAhwuryV2CsE/OEEMMOD3U5MaxKSdK0DL0TFwalNytB
tu1UQRyrOlRQZd/c49j+b2o34Or6JcvhAoS+1hjswknbpAhx/QGhGtVlD8gNSzri
QM0t6yz5uBDFkdFxcQ7/H5TAJnq+7zs2vFpSH+nnCsB4vQ4Lka2sx8yzTmtOpUUG
hi2hc5F5Tg3i5mDeYZo2yUADAYooW+kfszfEBRbIwL7tkLRBJLsObEqji3PUfEqq
0Gv6whFOqTJlFfOJk4M3zmd1/D9JLX24VvQwjBGdA9/pN+Ph8xDCK9bdWxRkUAYq
2RXSBZWXL4az3z0eLgZeu+MPgWFPvXS8VdyStHFmedICFeqpysSqUGHeGKnJw2Yn
0btgUs1gpS/0h8a0frZfeDjJhK+/xOdJP4zzVbJuIuqqrJClL7Lt4o++M4UrCLZ2
pBoG4NmAiwblk16FZvqlSJ6NptcZJUdAz/8FYdXbomIV8hfhdJtjRugCNtble1+2
UY8x16DvP/MBWZVD47OzjENEgU3K10aJv9Q3XUA1+gbyrkx5cBMqSUGyioihUc+z
Cpz+elCuhogvcuWJ6Iu4y1LwotibyXrnxb1VJfdxxZft7aqkWj6YB+aP2ZQjSuF4
cLh4iH0ZaQ9kLsLIv99CXlfPWTm0FqCE0umVKpnFd9hRUpMA2zMkIeD9YKVHmQlu
f+DFq/FNkb+xcNaHU2g0Yp0nQYlzd4+XZY8k9v9qxiEwrFcA1Dp7SjOxJl2e9Skr
dLuwjTscztrfBFEXk6ehjwDlREQjXIm48ROJ0hInr5nVRQHaeZ4IIloxw5qKtoPT
X+sCP7kMTnU6uLRtyuIp/ZymVhmuKrnN4UcOFx8qOTsVTCMjp4+rzZfrKeFLjuX6
dwubspS5pc7eb7xZt7N4wGuHH6oKcaeAPdv6LiqMxlC06bxUwyIkk65EjVZcWsES
yjBX4b5H7YHw8u5KrKxAkB5cd2MlJiu3Fqx5P4SJbPIsrKYK4oIj7Zy/68sAm+OW
u0yodp+8g15Nsx31eElZ0CjOVJZWMAI7gs6u3IZaSDYJ68+2glwIEtYRNB7Wgc4T
dydgPeJff6TRxN2JviEj65Pune2i4MEwZx/JlBIuUsLmbbBBkXoA0O80eswj/A3q
8FY7ogqKdSUH8VQvpZjyfeOgQpWgU5+oXD++UHTcRQ4MlEuz5bYf0vwqsN3IfDo9
C/KYco1c3QwHhh7VnGgHDeSrsk4139/bWwlVbj0iiA7UMF3L4a7TgzBmnJ6VdcZF
kItWMW9HJUv5TYbkIA6fr+Yjr2S1fcf7ZhM7fJgx8WEr1xp6t1gW2+LTvwnWqlG7
SaIO6dtsZaMyFXCaX/SXswz3u099aOr1rXU/kSaulTwZbYc+ROquYs6H0kOPO2cb
eXRA6UOBKMbdrR9x6i/avVxGKoJelHIot7cj4fSwuZGJSDBhDUatn9ex4pFpQCqR
jo49xWXHQ9ItT0xOmJZotIoWRZW0vBhF30T2m78EtRi4Be+DIF0+Ga4ZPrgOVyNd
ZXnkXDSHNIpQO0+esEXhkCvwvPoo75z9Y3V5VmGOIJx6OZd8asu+fpKwjDpbA2kI
VzPHbfwW6SFskJLBJETVOb0iyswtAQwUt0GSRBggbkIedo1Gf7UeM0H4pxcmML8m
1xXKUflVEQqMCporYcAoa7JnQqEnSPKjebQm+OBFY2r+ymIfFBHVVnAno/WpADYZ
csyxU8XPd1VBMl0YzUoURgpTof5EnupJaLUO8hUMYWHlqovRVNC4S3JsvOowceH4
x8Fezv0KgPOv03y/4nExyCu5yO2QFGDdLAzMXD5WvhVSDYsQScdLNpsOUf1YGI2E
yiIKdkItqbh3F+FXLLFWo9ADYJB6+LUrCWQIlgtivPjjn7HiFyhEzfvfESb7VudI
XcG7uhN3GfrAfy5SNL9/Ag1BgvYFaZh5d6jrlGHUunqv6QR+OtKox8tUEXf3KNgM
4qb+yXpdDa/H83di6oQwx0tMGUmPD0D35nGnmtJaOTWkRagAVXjftU/r1WQQ1B60
sEefoKV1uqODgu65c8rv6c4Tg0PZEg9vAQrTnwncwvX+zdsWPbZs4Jfz37vijba7
Gjqx0l1U0/CC05USrSFKfWQyYkVQtb4FVJ75n6N3KspKJnlpQnVMLLxvH1NKe3V4
/4dSsSBq8w+Kbg0RSQONhHVC1U7oGfbZLEAqig+QHgV17f8zYaibeUzzUEqBmmei
IxpTAPEhJo5U/MR95bUYHmNb21akxZdbOFfljk6W2OpZgtnMvGJrEskR99BHOSAo
XgTBcBV79zhWVgvk8dvKkPbFCffk9/iy6TMcVejVU+7aOUWpQHxKq4QavM0mwOsT
6Udht/DfxGMDjQojWFEwm+dgmt/tLfHg/ZGffd5dbQRwLEnl/tGg1wkvskl9gtYX
dbed9M/sWPIsmyxfoQyIuDRzhKx/yLN3nTEwzm2G4CoMb0efYW4emZDOemOQJoKI
VTlQEnXI0BwdXWsdWbZdLgGHOltR096mxPDBnwJO+MEjjEFVBhUlxwz8x5Q76XhW
zu3ajyCi7Y3arv6xN/G46Wfz7AHW67SrzyT1BaIZpuQ9MNw0aiJZ4SseCMAjsr6m
UShkw5BWwKj90B40jPjx4VzYObPcUg/FjzAv1cskvX9AtDmbS9gU9xEM2/bGS9zO
R7SXembzdguOnt+qwmf1qxXNtfKgBGkIrFtOEdTvYToZ7P2R0DSTwjjL5Whtrxes
xW+B8/+O2GAwsIXOP7VMEmDOi8rXrvO6GPNrgayq5rsK5fjwJmpFH+aDmQS4oJZA
Se7TspMZdWTHz6J4dlEigmYgIGlQaSsjZ6Ufs733JmQj921RAJ1PbSS0sH7mvLnz
6YzRDiaHlOxwa9exPRZZEnJTnIx1pLiv11SoQ/wwZEYCkcv2w2rY36OHdxGWZ2Eq
bppTmBHTHH8TZjIXlL8gQ4HGLQRsD2uxsQLqGViq1Bp+Vqe6iUfBWyqGxVbSws6s
B1qlzFOXyjeOjHvoXwafekYvE/OTgGf88/oN4LuT4p9bD5iu4EULgXhuznCxYURT
EDlSZwYZG30vstAncmDXQQ+VSp/ZltNZS9VcowRLokga187KcmsRcVObrXYyts9V
zqHXichwOwk7pbfKY7k1rjA17/BsoAVcjFF6L45t4augdR+c6W0iOkiryrnzhwXs
7X7XrGQ3I1bXNelx01IMJf19tx6zCOA59sjH925VMcgc1pjhzMyZSVEfL118vtQz
Y5Nr6eSifNuY4rZd6cYXc4Kn60g87HnHMrkULpFEXNZM39l7VftbrFc4AdX5zvNV
zKOQhchAJ6ZhfIBEhwA63zf+CV85eOsRRKiHmYtozDTyr4eEyweqEDHgO8z1eMVn
fLCm1hVD2zN+w55dKT9esSc0qRDEdMrD4LWxDYMl4H/74WlmzYlzPuDj/JKShj82
86mO1wqUYGB6VEn4tV8yE3n1eW1U/Zj8GUiS/Gt+5QKUIUQQwZ3mSVvUv8uW4ZB8
RT+vFhbvRnLEuVei2nDVXj7OxwvKH9hovRdUAWVoahsNkzaxc21ywVDUujaleo9w
rh97CSwaj6U4YVNfwi7NJqlt1BlNhl68wp9XOG45IkXMBconnKyeGXtDtBoWl/0S
pj1K5tx+5u7xWdTUCrBMuJ+/ifEEc+MexMMGUwVXMVN7NCg74eAegAAdAmfcy5Uf
vsrez4D5ydJZJXOAIitBug4S7ZkLBPXMwe4bz/1G194fg9nhAdL7woXYWDUNOhda
YsMReUjn3N+xCm574FVyxI/gQeQyyjLWv4ibthTYRUlVonsqLmhBt2xwe7vwkXBZ
U4sN/Corzr/n8uNhb9i4wLZUZECDzh4nAQxHAG6RMs46xSABfVkS5zctylZ89M5J
yrd8y4y3r77zmtGIJ4ufyM+F+ETXbQQEHL/NMZxoFxpOGSdVVW/nIspI/bOpZv+8
QbupqySYrcknIzRSPExC9m1dxW85cyjkBdxcrG7lkIi9XY3dHCtMcPClpnzuHAiE
AVRDMN1c40DJZkOQtrcjkDCrN/E2nWet0TKx5BM8dBjWD+mZffh8Njj1I93wVG69
BNrFKiFaHHG540oKVZXmNIXkV4rJ2sfRqiK34qsoD2lL11eHoMyRr4jzLCAE8CqQ
hpZjPSwBtATguypl0W9q5PxZl9A+DM3yAzxxsYEPK1eJ6GKPNl1YHhld46fSlbrR
iphPcgMcePb596w04XUJLCp13wf4Mei1gQCMszeblp97Gu/Rz1W+/vPDTmgFJ12U
hvgzmOFUvpM2I9lO+mKdD0+q4sMdyUmhmVKbptwqwtw5nUtteXFocxwx/xgB1bqO
fFMV5B+8FCUTtHwr3QN5BPoRwRlEdh02wQX1p1YdxehesQepuVs/PHwGHXlrr6lm
niE9Lox9FZoRO7uLurmrfklewF4BNDcHB0WA5HHw24aPV2zOHp1MNApG+UDnyIjO
Vl1ALAWCChf1WIS5/mXdKecXrtNcu3cJnsAni8PdS+EMwStygnAkv5CiHSr0qDvx
DEQdIbCvSmldwCUZB0hqMksDsqI8KZuB3sQ1osjguroeAlxpseeGZ6mkXvnvoqjO
b6b23GzmpQUiG1GMCGX8+C3jygZyx1Q+5jitNPVfOTBLRD2oN9uQCRNfGpPZxPgz
SLyU4w3GLCdVikcx8dIrpTW6pm2MEsWxueWMcToNEq4287sbHxBKuyJa2XcAQqAR
Z4HKoAL0aMoatbL5RMmn/8sUntWjs+BSwoxHJbS6ZG/2SiV1YZ5xC/hlZHPn+5mu
GU2qntu18aalLrcef2Zux7sriVXNMtbJuPqv8iMJFlcIdWAd14jth1PSyI/3d/Xe
BcoPiaUmqfCyWjqpTQbjlB3YKU9P5Q0Edr+HejhichleevB6ivvIF0T7EMqGAqbv
rvw3M1vvTxGDSKkq5N2VJKG9Din+8imgmQb3Yn21EZ0lAJ0l5w+kNyVOSEeCXjCe
JG/lSzFOcadtXif22AJRZGN4ypi/5WRC4jCzp0PjthAsIr59tfE3jOZ8yv5kGFyS
9Tjs3n/bWc+3zC2VGf0XvbFz2iNMhuEDhbEwc2t5CbWvfMH0yE49ti5/kzOCEi3y
BXHUFyDnckQr81f6s9pUX95TPg1Z+lIH9HDwg5K/Nek6evske9ueoJu67fvE49WI
80M6BT2D/vKRr6+h1EEp9eD59Y115q/f6x/nFRizmTY9AsGmvaW2yyyn1o0/fS4y
caKuSei2LxQm0yxvddQLKezl4sBoVn2UMwUFvjIdSa3BapH/6mht0wr0hylFlp/S
TnkNPyXJscuF5SYuMzmn2HpM8zqUSSs9ciOFB7osKFMY6G6vJepzpp+7OTuTAcWB
0fbvUQAL7nWAMkvy88dowSfT6a1A/VhDcFEqqW7wx5a0wZUSp3Szj3eAcb75EXOq
6lCaUV0RJBKaR2+Wx8rNfAIZhhBa3uSSp6DNYmsZPfQ7Jj5lrBxiN7wTZvBPoCSm
08rH718wuMGNozw4x17bN3gy48M/B7+maiZBg4fCfvPpcDog3yBs3YX2AbWUEnCB
MyjfZC/du8uaONF9JA+4meOXuTcSaPaVoeYbq7M3/M3uB7ou1GDpq0NAg5wHYK+6
qNlO9uEYqW/qRcCVS6WniQVGtdIPsP44zSSo8rblGyraPOZtkwzgisWrM/lFLYZW
QClYbLjiQvAuBvUevHQx2LHebBZBoOMhGZIltJZOMdu0fPmFXetcdY3tO4JONCpO
UoSVqNYfZNdpovy3rbEHEWSuLbHOWA5sH8XcHaZpcsXLQ+89uWKDQf4oIWUZSW+G
m1pqs+o5FV8cjPSsI2DQ1IcKqezulkvzWnW0tI1IkVakjyHEMBnHWR7PoRsvGA4b
DX2wNHcCL2GY9TdtPW0QpWQF0aQRaD13tJbphzNezjANdGqJajcJ6dd8slgNhn0K
V3pJ+RAR2UVFSO0zhdRY1G6godOH+G2p2aMTTcb2VHskvBROHzF3hkRSivhZI+9T
JWdmvu9p8XSe96eg+bzKQ016q4cm2J3oCCxVLjqwaN0Yx72nUqwyjmThvIVEwvVi
dsud6gm3MSbg1bJ7+0wZfPZ9nB48nC3RtKQch6UJ8TtfiKYfxuLfpYfNNF9sq9eU
/wD6vMSnFolu3P42U8tcR+MF+qoPPXIn8oxPgyU9NuJtXaqhYwJxnBIkxvUUllFa
kRBahAGfj4L0q9OvAxoqnszWbX/ymDvDPYR4RN1GI/BMkdqhY/olie5wEeNbkCIm
E858olH1G4yxnn8LCRKmD1/XuHrpkl6CKiJ8peg6xEVqCTkYtZQJwukZXTaXEAXV
41wiGd2R2idl5s8xYAbDOx/fKg1wZnNC8nrL0x0tVxpxDBnBCMMFYbUMVMaeyaeS
RGnKbUNXPUlS4SRRWAB/uo8uBrkaG++uNsleP7YO/YoqaN9fqyxvnYOgx0QMg2eW
5YBlKhiL78yTxRiNhsxjhvsruy+ogUFdhqX1QTr52fbX/OCh7opghbmrHFrZSHdP
L4WaGsIye3efWYuZ+/X6pLj5vRlu/MOHotOWozaW/MPlao8dT2Mxxdgily21IZt5
NSe8cji2F5pwlzBe84n5jT7QboJPyf3eCpfLi0MD4pE41+BD0LKcd8garwnBiosB
VIVZ3QZjheeH/6LdLlxy2O8Fr+9SDPlTOuqZCkcfvseHnlLByVFV9Lz9hth8xVyd
87ZG7W7B5XZCrgabcI8+gwwSVgqGBGmfVEwinCo838wfZ+6RMSjKa5pnQoPAQ9S8
A7q6ZSC1Zd272b1cwSlYcrz1FCVSQ5ATIiLrJ/yoK9HTgagGL6rDEAPkyt9xDZyk
Z1HoYweztHGe6mCbWOS4fn8I2lhJx8Q2J2qNe3IDb/HMhlJkIB9jt6LnDbju3DDz
yRJTSOvQ68eHVURq2rOTqWG+M8aU61dkwSy0TcEZDxpw4xMtjSL+5qPNAaWhGbGj
FuR7w1LM52x7QM8skSbQQNk/0TfUy9t7UPYydkWfEFAaotJupyQ3CT8BjhFSyeZ/
ON5ZaPEMtFrltGkQrZX7tCtra3t4debAo/wfcUt1C7dQb57xuSESlRnbWMihuZZG
Zxxc7D+LljV3aho+CN1CF1T7fxvASHkFvJsslSQDR+G2sNh1lMKa2HwquARfnSh9
WJins4KcPSDTtxhw3M/me0qZigipTF4pS1Rqz0CmC4roEzaTa+yEX0SyGx+XXAxA
0yYzexXERt9HjQYe66xV5TBD394xW7nQw7HirrjeCpPTFP290FI+Xeo8UfdwOxpd
Iofx18340HNu9xCcp1Oia5rcBBL338JAdKo52Ra02aSVvwwAWuMWgEuqKXifBh4h
YVx8SIWtBoW6wKAs45FyTJ9jKzKr0jXUuPAXkYjTS9UGxlirC0KvzkIVE5ioh0zw
iLamrT+veEwZhIe0XymQTYlHmEchc2rnlLwRalUZ5lQb3eMFHzHAcmstGV7MReOR
gXeg0pWbz0cBLtkI7gtunzxLMawBTZOdQBNRH6nKyi8lmvxoVUrWah2yvOTiG/Xy
N1z74AYoG1iP6fNiEncxlBOF1X0LnmPqWhV5yNwHiL2LE76qNp0IahmJJXExspo7
lUdpOm54mmv1NpPqtU+6O4cRxdyiuPb26Q3/JyGGLX/o7TpZz/R9E/KZUxjEK7jO
JUwJ4IGFV2YyHh4prpeCsM15E3uIdA/uPcaKv6vj73W5A2vwDWbnCks9Kwj17ZWy
V0LjjkajhI0/IlGxHMk8gxK3Wv7EQ0jcycVKKv2iFRoi8jNU5LnccpnfXC6vPxzK
NkhVzG6R2KPaIFmn5iKpOJOVoFic9oo0B0jblTre88W8V7nNvexG7ArBUM/2lGaR
AeGqFQsF2HH69SFuahASyNcv9OaAEIn4GXsbeMQQxFbT4bcRWeEcH4+zgI7aCbSN
lLR8LwYnYm+6iSdBXu+b5xr03pxj3ozBkaIBXokV20J7ymhRenNRvqDoMh03q06V
WuKXHM6+Z4nTklypIf9xwQJCg89cCOBF/9QFyA6r9cbr56VleK6lYzEOPOuY15z2
a/mS64md4M+hV/dy7R/FMpsT97wqxbDLofrBdJCppjC86iALIuDn5HDpFV6q72I1
pQAKIObk2kNs2cylC8rzsf2mruuFtMGryPolbFIoJDkdf+BedoGMaVOaytp0DIU+
l5KEJ2J8Hs6IraXsoVvBJ9NqJq5Tb7VYEj9sJYDRXsMWJbAa9oNKUZC+GewqqRdy
o0pKUzNvyWKibT92cVs71wxKA+NFYGxlOVRRKLdqqSyzWFQ+9QD7YHrRpSDpkKqq
lco1CJY8WE8DjoV2uTKTRBz4Q92xJZYYeVErfgD6ubBsF3Cv2Az+7ABLEpUUXueH
ODeAE7fd6PH1vPc1xeJat4vCb/Pqq8n4B/TbRV/SQyLyk6UOKwKNIdDJl95bYoib
hKYSCDI2TrS9BoeHEFc8UHK4B90UMWkaU5vE7Whyo+NMhLPkq6TNfGzww3kjgttF
l3wpdt7CH7viQ8yWLozxsDYvl4bQOyZsOdaMjCBV6aSDle5Qd+nXR9AnplDVEMNC
R5e8pGdW37hcUjBdK2EW707HJ9h5zgxzg7m/8PkR0nXRMK3609V7fRbyKaKK8GWH
wbAE5CH8ZRDevg8Aw+ocmWxeGBdLj0aVzmadgRJZbFxh4lHrEeO5l0sAYfMq4ek1
twvEogF57i51UjZ7VQj7GWwkT5kIii7dqZkMrn1wVLMISnj0JsdHnvemB7evH87v
ziqxobAxh39HKa1K+hCcXepSWLK4gPGuSXDzxsVdlaxBMFIw3ATdDiu1CektzA7I
oP1g73IqlEJaA9mI5n6OQv77Q8UGDnzN8QA3snsLP41RAy5w2A38BUBSYSuzGzTK
kQO2E4EBDR89bbnqDk412IhvADlkBvPJ4VYhXMlDx95IjRXzREdJZAVngaRGXhGA
iktFMBJfLR/92cIaMjqZ/yZGhtKrPATQt2aSGdGK/hNmHlBGy61R5U7SHH9hON9e
yd74KxceGXNCn7cFNgwn127Lui/jJjwJ8o/A2a8VHmJxpfub5ssS1MFRpYjLUTHd
5KbKaSX6PmmW2RXQhe3wFwLVpmQ0XiqknSBI222yfuaeUK3vKDamiizG1P2uv3n9
W9mlj0HQteEuGnxiM+SLZ4W4nPg3Hkxo8PxPNcwPIZEB0wy5oNPH/wjcOE4+y4bS
MOrhoJ1kQQ+8s9p14xg8ZDMH6x0zr/TliLK6SzTbbytVDmfhdU3V4rAR+I4st83M
fs5g3550OIb/05lD/LdaNz8JeA0PbNoBtvrVb2iG1kwCMrVrGf1RybH4KB23LJZ6
iJb5tNhjd9jabzX/Wjf+lbc4yh8mopiJmUIOmyC/QC4ewb24wgLSOaS3vaoz/P6p
lUGSWJ7h/Ns5pKII9Ex6Jh4by+6EOY/t7BAKQdiz/N2stjbLBQX9hh5Tj08q3Fsm
EB62jCQ2ENBlOcAF6SoQhE89zpiPeGzAEGkmV95RB/P6BBjkB4R2qEZ/BR7l8OlU
mj3DH7A3Zki01HoNDWAJndzPoVTXDmzUcNL3trvgk8QPy8lnO0Q9J/uModDjXXqH
zlV/woKJ57jJmqB7iWR3VCBhc9i9CM19trt6W4cTs8W+iSvYA7I0zCtLub0NpeoU
HvadnlvZC5sB5u5BuLjCGocLCrk1vYtkhn3Wi8K0xNAjTYXJBkS+6WHFqTh73dFr
6JgHG/NWtYrwZ+/YgnFMsLBibdYg+TVWqATNQ3E12aS7rcL0GN5YrKOZdeJcjQ7B
Pp6TnmmlP6HhDJye31gqVN1xFVXeHGuaF0fV/pg9kh1PW7vvqYe1w0niHbkK5q4o
qegjzDPa0krKW2dqGWAXgECFRUb1E/T1SB3FlF5hbvbs4rfP0bzsD4olfWCSq3AZ
NI2Ylb7icJcQIu8bO5IKK5bkWtZXNzBJpbYrf8tP14MHi9npKDLX10vun7fk2xfQ
QQkTmjAjSF4XB3vfpiRQ8q77IGKHtm1iJA8wI34ODUzMxt5MM5lNIdl3rF4HmGZ4
AIrC46PDAT9g6zEsypFTQ54Dhv7RcY4o1Xq8GcB9y/16Ws17DCspcHiZIaGFhoKA
0Nj/arTREwUgXrAA/bmW7waeIziTD4huiWkkyqXhaLlrse8IUu4TsCn7Nmr/kmFU
xjaWhocGWYZ3GPvZ8dZvJnkxKKHyae65OGjF6hUp+oRYOkq4Ya8C8NTXDbRQ+NfG
s2T/ZBlaBmwFzTMyHOvdF8CQizn6gKYTiKkGObgn2EgqGQYUqM2n42OYqtZHeM0N
y21jEaNK0qpHV1AT9rXRj1lWoWi04bpY1pe3ZCVjv77yH5xg48E7DN5fxKnu5Y1M
eYTBGiS53hyMT9ArpFY41FazwNtxRKYxMkh5z9nHHf66kiY5h40S4mY7xHTw/VF8
uaSVtsC8RJjwl7CsxCnXAksqoiJ6rEgtXPkyOrw4c62YHFlRqVoLwcYxdyxCfCt7
DC+Xm3eKJzVtd65ey/0W7pMVhTmpSYBd0wFXi3omdbPmhXN96xn5KAUkwmj47qHq
GySsv2qBOQ4Z4T6BxGjacX7Dn3ooBqzMauyIZspbmz5NcxpUzEQpDxHdXqfpBpbC
97uz21D6/lmEd3n+WCwhvDelzbbAtKoyV6wtjqZh0L9v+1jSX7ROp5gXlp2C66J6
4PgwtPmmjvQnhMLULwaTRrXrvG1F54z+yKif7+0cBzlzCmzADuLhXiIDXTh6NxdG
yIXxBi2VYnb2RHSmEIrwSCSn64vfXh5m4gwPFbn5I+lGMdOQOStYqCrkHRQaRMur
PzZ2ShHalD6vPPPPcnGBkvLJs+RDzY/7tcIlubsVHXDfYJ4nPmVzwZZdETZF84Q/
CEca/gx+qX+GU+HSItT+8gkQJVo4iuWI5KUIxnzoJMHbO3ci73HBL8bFNnJpuOgy
XrHD4A5yf3VKiQOdD4mDlxqVrwURDECWl0b4nWd76zIa9ULqfgYcxQZ+D2EWieOh
cViF4FjKcqc8a0Wr5G015ym3IEAbXs1eK5aXiFs2J3+tyQU6CzlVGyiwQV1Yx2oX
B/cP99fcyuWxWg5hB1IsHA==
`protect end_protected