`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8432 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/anaBVTumwtXp6e/AWaEdufvljN4ptt0xyy75lxJe06P
SJ0pReMo748kEZBEZKlhr7BdfgQ2q894dtzhl4Vay9AM5o57MqVmi35SsdbPozbe
YHaZr/D26BQwmJoH8YlAuC6iiCQPAkM34y3Mpzqd+BgMTnQmmO7d4gTeI99PwavA
URvCqijyz1rv1jmg8fq8J7W2GWwK0tNrKo26Cw4E7yPPtyYMHIdbaWIgtmpgHkYg
EUR7K+A+sriNRwgK52TyP3QEDVQYwsXElAZzq0zNFBuh7pNETHZSubSKoNryBZH/
57JnfADKnTU5ug++Ag91rq2jaUedOm0t667PG4wH/EkJmKTlxUBVeHBgDk5xel2m
m3wVV884UnDSNlWRXFMQKD9uHBasN0KNMQCr/JfGeBXXb53rTxTDiEs2m6YhTL7W
m7ZgOCILyIrjrpbCT8KYo02dv9KH5cfl237vUo7fV2GF0qrpwPuTixc6SB3GuP94
1w5ijoWht7+6iOd5qgSfcNTa+qdBmfVirSATR6GOUd0ApXzIjZei2sl3X6dPy51V
H97tTyhwkf/jqioeTlOHqosXvP42OnPajLRYLiUGCYe97FtJ5spEa1z6xtDyoR62
EzkwezHR/GZ69jR1stZ3j0z5zVIDGKkokSZhg0tkeSuxq73tS0Dtf8fpEH1FJqkW
iyfx12QraMCbaoWDysYInkt0t0T8lwzrtLc0F/94ON4/pGajSmf+k772N5PJNYyd
+Yb1mgBWn5wp5U1UUEvgkYn6ocaSMq4+45ACF4n8TiOi+HjlbS8FC8iGCIM6AG3A
L/IhI8nu4E26qxdO53LK8N9wdR1VRSYFdFGCMo03Ol4vFWn20+EGk1a/wF6i3WOV
8+x4of7gevNFmnhrltH2qYHAZy8dPVJSxI3ss46Es+oz/kvmZJ/zVS2V4X44N8uy
UorNgKgXsCcyWhztbEmZaAkLf6d75J/giSzicBNGjPqf4mBgVL9RizDRTNiAQw3I
3Z+m7Z07TxUGC2BRW4rc0WO3c3dDyY0gVKIsDsyBZSkj4A3BlcdsUhYgiAfxJuE/
QYWOqnJO3kt1US5hsUXjbNsfJaCc65r6yQWGb5yCAP2XSJcgrZ7tINp7GWewJOsP
XUD/CXAblwM/k0tRV/BHtGPaeuHwml3VqLUGWQGldgRA/P32VBkiFMvolqCB0EGd
yR1dM8I8MBPf+uloAl0DFntlq1A9/uiRIRa3Ap7q+CnGAMY53r2ZVev/23V5Q6Nc
r4dQL194H3drescFy7SRkkbJaG09MKE9LNORijMk1Zc621bAVgqRs3roA62JvCm8
ifbAyX8WlQLpPEPcUYUdk6hKNtUtPGRd+ZdI+RuCA39kNZZ1Zp2zfdUbTBdKfqJ9
0OgaMdQz7TE2faRX+sHSVsY0gF33Xb3brEKlbUCTzMOgpyvvk09vBeREM26N4ynI
jtq38jG0tfUMO5sbInufh8Lza0B4FG2i8gPfReH3fGQF/EyX+XuQmckj/mE9s+jj
0OY1JLeAsrt8zWE/0dH6vJAHejZkiy4dKfuIRO9dsPmfwhCvMQek8OY4mdxpl3WB
Xi7Zx9fzeRVOvFQmlcUxrz6H4ZgMVRcZQgIpsx7KK3oy4v9wthDcyKimcYsW3D+U
RSoSUc/cF5rNm86226FefCLe9U1Eblqofvg8ibnhKO8ESv8y0fUGAZvlWRe3SNsr
xmRGpcHVVII1nyVwmoYwEHtFuj9KCM49Gy8fvHMfTAa+CnW5cvUXvgVIRXLDAB/P
lOryYL2nzP1jAQeDi3928v5zg7r/7Bow7dH47ww2FG+WD+X6//fJYLFtkanXWs59
3mR5JcVOuNXA25++vLPEjbZwlaL3r/HmFKv63cUdHttLQs7U3v35DZGNyjtB3+7x
p/nto54U2Npp0VjyYJkLt4CqQiPX6Ho+LOcRFm5+JcWowTM+mhgWPAR0VEI0iQ34
IJ7RG04EoYcTuAVBNfPKRCaCYWe1YOm6RHmdwxUFekMAN+0B0Fh6iYP+IAxMIdFZ
5WaaRzkaS8WlxGqF1GF0NXeMD1ZiiKna3qwHtqPyshzgaK8QoeTK9WSpzmhJQeeR
eelPJ6YhlyL+GmFETqA9xrSXMHGV4Z/P4lY4By7N66Yt8crx7k3KjDw1j4qr6Ux0
P79YDNFTcagUMQDUoCQ806+1AojnTdfGoG4WRwK5/VmBveS+Sm4rbNpnMjQqj1Kr
wOKsw4taHTC2zKGOZ38AL+WnH5lRCaiW9EzHgRicQWkxARahX2GO/s4bLEob4qf/
CBhJWtLHjo+ciD84YOYcn3vTGsPxqHK1q4+H1Ngw6bQD+7S7EGiztFN5eexDC0P1
r2T6ujkOPj6o7IZaFnoxgmedKFV4pjM7uS4p4cosLyDF/LsAm6HJpGGQ50RO9F93
BScnBxMvM/KoiW2yB+fnFQwl40xaFRi3LaCAqQaaooUUY/iFkCqFYrmItKQHT1Oo
iRAwxiiEzDbAzIsqZyrTIkK3liw0wvtVeIQC8HyqxeQgHGyRi508ZvQDiiKXmnYZ
TgHkGo0YHbljf/eonB0y8FjpSTtp5QYzL6CBo0wIxkWGgIFCJwp1aXKvanvSQhIC
OtU59IaIhAOV6gs10egSBdZZcRTuID4DiUhXRQPE5BtmOYfYSOOytcuNsbGDtwp7
fV0L1ZvY5Iyixw4X1dfBUTaAZKZEGxHm2PturVG8Rwl6GifGXXC/IGTvi/ptX/mk
x41XxVPxAfTQH1LRSmU5i7KYenoKTYEEJgugJ4S7xA3I1liG31+k2hJwJy5YFDW+
6VjZ2HOayn9MVVaLE8sQ7+h2sUsnSLUmLHBikjwWy58bDwfmDBh3WtlQHXPQrjMI
oq/0KFwTx+23SbZSkr7JaXzbLMObmuO9Ub8N5/XxzR124St3MWeh6/bkOqE0pVy7
uLkJthyCkm7CnEU2l81eDWzd/qcNVY4KHGnsqA4FzBgfGOJlzhuUGxtasw/+bBIx
22MP8tXEAyQKiZatbkAKhF/8mXtgxC4p7bS9x5u/Q8SJDYXHoZpiTOfgBk9ntj2V
FhTP6qPSK4UMyQ1oxbYip25JGDgUh4kkRXCq7j6RpOYu69x9keBsXdwUozugVrqJ
JDtf6eCP39EL0/LTltndILMH2s/dqFGN5qQExludC1UI0vBmfANm0iPsG+oH2pvl
jsD4mBTKqZctYueOxY/C4MhWcE1eCF4QOlS7pmC7DaH5NLLxLHhiwtNLmj5myl6V
UKstDv/nur9MSLQkAGJL23F8JkZh4Q4sTvYU0VFAgq4SO9qEODbqecyvTXxdOGRr
1N0MtrO639CxX1/vSHMQkRXT9PZUFl9lxOH/t/PMuVNNPjkw6ux7yGrppHoIYTYX
jgCMimq/PWraxmktCGfCuX6Sx1qDAcxk/4vFrPu5DtvZVmn8VDIev8b5J9h3Np+g
nhFrCFC4ufzufZ6QfGFv2KwvvHvosvUNy19BefbR6kw0OaPSo10eY98G6riK05gt
1gvfO488nB+S+zC0PslCLNi0uXOsindSYGBiFZKoLGn34YYozFlRS94MJoK06VUC
LTnmBErii6TLPSbFaJbTY5YexwJ7edg9GVBvkmlwN6+pcYmXBSNLLcmxtmBf+5iz
JYCjAF35WHgxRFVcFb3F020RQpsuK+0xE590Q0R7QoRRuwOCQyHdnV8u7soG7ha6
7L3LUIxvn8E5OPw4wnqk0zrIatq010AqFr7cPEdBY8Sj4+gcSnt+nZGaqQYcUYgD
JfHHmQW0hEbkwvdN7evQjwTcbzRii58y5OzF9IFQPkBqwLvWVfiRvP2JtddlmbNt
Y0NA9mwMByTNulYkAbHRWy2NxuUK3xS/I89WEXLocQEgl4ghyog57/XnwuVSY7O/
4U7mre2SxyLW6aXXjxMWRla917uq45jJyIpdYWBTjc/5lJmTbErmO7x5fm/Y8Nib
h3Ja1c9+URqtRQXDOts2YuweClYZvcPOy87vH6UHXPTL1UizI44xA4tUCa8Y8d4C
8WFCKHhhzW2fgC7oqeecnFFymnKfzFKeOTDzVrSzJs/ZOndzSg5k4x7QgUOnO/C1
dURZS7tKyDflcHPoahh+ehw3hCY4YwxI/IiBJBR+YOJ+SK1zDb69s8pS+MiXjTXp
9zmGjhLW2AAnvEc8hmvYnKnJSFzhzzAju5il1IZVw9J4bC5IffRdesUL4wadZbS/
YlYgqPyBmHb0yhPDapGXe9xFwMIlc1pcVhxhDZpmVPO01SgIJpXwywUIlVeRV+P/
yAvplbTDdjui6YCkcMgNA50YOQZ4XHhHuUmxG6SVcMfwUuLp80wwpyw193o1F4va
l0SWPFe5DLhdiQzQy45gYz1WQFGVjexfJkfHPOgfsIYsLwbvu6yRVVaisAn/+/xP
eo8lIRdgikZpgYj0jIBLOPmbG6HJTvnq+OlFgMTn+orGJafHb4bOUWQ/DTnfAZ+B
O46V9qTaUif4zdhEqUGFsbG8tIRp7Yd9CBKnWXv2C251C+u/Ix42dlxcGmX300HB
zDieGtQiFtpQNffdDL94Wfk/vXwpKGdJbLm6v+LaBCK8oYV4wYHnPG7BfHXBQXqZ
93vxLzWdrw5KaD6YZuwfgWlKbmWkcEuGSmVpOc7waU2AX7o6av3ZLSP2PCCD5PPP
lEAOB8CKD/7nZbGidq44OWyaFHfWOCflH48pw1AQzYyWxqHFQ0c+oXBX6cYfEOYx
DiVNOck1XXLA8fMxMlNruEHYkYGmWxIzW5V3ubVBiTLHPgTwwxFMbWoVrVS6IERm
khPXeQcLwepIYbgYRsM1809a2gGYGQVKtR2fVXK3ryelPBZjfMoAkhfWl8xtZoac
mpJz9DCLwE6HHLm04exSMFKVTAuHQidu/LM83+LTpSPQv4HRGNIiLy/ZYKzqKh/c
qxy50T5nmVDPpYDQSsOXTmBC5ubwfsiRNrPrWxdtOBLBC674BvTPtm1IZLMu5hoP
EsvZH6oAy2MOQX72u/k8hdh9jT++p1zaq0kELXEHib7nTQpAl+COHxHMPwf0CPul
8Yrd4UaTP59QVfh9AEKF5CiZKDvcDl3AkZiX9hOpwg6iPDznzv3GesNNlS69ILmL
KiWZ/z8wk12jIAaqyB5/7Ej+MOJqE1eNmL9HpSx+FOAKk76KCyU1ad3fzel8AzVM
HXfGvaDqfUg7VqLx8rDiHHakAC53UK3w/SjiHolawgJkaCuNBvd4xJQwWymSeKYe
Eul6SlNpljDeyK8gG3pXcEXBe6GrhXV8CEg3CYGhJGV4hIOro+LRN5UD7PPum2Ft
lS5YG8jL3n03YLvkt7+dkQz+DJLWM42R9bmCiWQV9/p8Ok0zbdaL+a14BPXCF8p7
2xXrtrgGi3WQjO24o3Dw+QWfqMlSAHLdUca1r6Lv5rZpAp54ln9ycsqi1TQqj2gN
k6emYqwsWq3SagoXjiujprOPMAk9yDqCcWzLX83baey11XQn+gYTYVhEAYDeKQyu
A20psDc876gjJsyqvKOKP+WoF3YPdXfX206fm+VfNECzYBf9o5ApIySZpwd42FpJ
treMbznIgUgnuZB4GxMRtYj1kJ+ChjIaUfhwgSa5GEbmGFeBh062XlHBGaiFFQxj
S9P5kW/fLOWk7LjCAkUh/ctfdNHFPSjMCnMdQtJ/Gdg3823JrnbFkDzs9czxvj0T
2nhDTaQTF08xN0ody4l9d1d241jbnsnlkisqm2heTgYrt2eeQYPYUZlsoq8TBjyP
M54cBo9unbwrDBXyWKWKp4EAZ/qpaDv+//jRhBQo/6D3x/ZDfN8DL5ekale1yuab
jWdhxScNRDlOMTrVnjE8aJBQUBcI3SEGzqrYASHQnxgp3OkTrEfByA988iSMZTZP
4SqfhrBJq/UJ64EH/l28mr2BUpaWcdKvysek1T2S50ron6JgBldZ+DAzoBhFkVXJ
V9nTuxCeMKrTw31EMzPubej3A/PRimXCrNQvMJExff5d+tx5DgbccmTBljq7mhmg
o0xRWP7RdHOIcjYFiBXk/KHJLEQz8h7ewIk9n5HyLpax+8Qkm00ahRqGzlLMFIad
p5R2SD2q3FouQZ4eWRn1eI6j+lIbVxIma3PwcbTvt0qeSpd46iU8diiRJATlic3S
hiXLmdlxezgrsS2PnUVo7oPz3LG9FYqn8NKw4ZuqTSPJjPuOT7+vNqkFJgJtnsIY
n5jHW3Tx6D4FY2yQIYw6eZdkX+WlgcFyUH1FhsJvtnoKW1gNLlj6a4C8cD5+KwTK
Ros3LenIqI5Ra3zwe+Lz8BHZcaUdi2I8cWOTcVPrGoXqf3T7miilFGrFvsC6hpnk
xqHyOGD0V1y9cJiXOPJr7s1NGQzDrR9yKWMSZajH4tn5U6BWwzP+srlo5eQAsKOb
nhkmFbJ/vtj7H/Bh8kyAaHmLxuNZvgum55A/9NO/CP0aLYrmBa+oj4BPNBlGhDWx
NeQ9e5cyUYe+62oEVZjP6k/xP5ly0obETS8S6rVUHN4eKtylEoXbRjcnxuVRDcYE
A/XfIwnEH0t0/mz+m3NJjVEP2B8cWHjimobKJezvpuB5Cf1hZEl7mWMP60yiAyPn
nC9NudIpIZVP+HsUboUc7R+Y1qwHmawCVtOmOOW1eFd1MFCEHVHrGPYFMcZJ0pw/
iL1qe6v624C3IgjMgqWjV2ARUK9EUjN3nS9UUHGg6ZUT6nflE29XtL5PoMZkBjzK
WkonHKeYSOomc7NbId63IdsAuBRrobfC53j0KquKhTS3q2CrPhRRpZmXvFTgXnCp
nI+kmi1uybA7t2knFTZa8gTHCl8lHQ31ZnC9CEln2ukrByBg+WqZ+7ac0eYW2LMo
vcZLF9negOOobAn9uATSAlTlqHWbR8PeIIP2EPvQAcKhep3gseijIiIvEg0a1Ujz
akiXIR81ysNbjIRzoEIsRYFP+GawxhN984nUgz1LwkTrq+r+3xCKyZbmdwhW7VUi
ZYaUAnf6CkT0p4DEOgfedunuzM17O048axcfigEEZOmWbOEmD/eh5JxiqoJ1nprz
6M4knbVEyavZpr0iesq0jLChjupI5FiFbmvOgdkoDIhv9sV4u0ipHb5reiezCGgU
osipIH3FufYu21k01KOWpyhreXFoGRvVvqlRtj8rk5mVx9+1Hl6iKskPYwcFFrti
ePpJKrerB+EjxbW0Rnf1cSCwssxmufnIGjzjtfSmZmCl6/wZZfioUIbgiABMJ3Pr
xhQp/vAvwOzWAiSFSDO669AuGFfKoy1dNIngXEd+6seSWd/D96w/mP2mXwvBYPDt
csIonWq+HZVSCcTWS5B57bskALZg7i1jQyq1uwp1Rgf5+NrWLibd5BkXKfdzgrAa
dyG0SQrGrz5goObNOd/GuRJHxqJcY+AwMhJLFfTzu0mW3AGLOu3opSbr8fBU5PbW
AE0r2xJkUjnt7RdnJVLuGu0T84U57BiF5EPcATCKPh4C+Or34JQVGZfcyZdEL9r+
Zdl+ba6thYrZnATYDo+K8JmnfCpG9TPMSvMpv4qLUj4k+2KYifuFOHYvSwh8aTRt
bDokr9xWWxPphX4DD63x7Wc75DXhxZlDKmJGPnBonudrZ4x6/sEZhFU5zxh1OgFP
4jcacrYfmZKmnFAnc++SYMCJ7sar1I4zX+MDMel7kr4oi4m4OFDNGCuCzPHBlo1p
pnv5SXqr6MF4G6m9NJtM7rVcvI8jmq78/oLVdwBLYm18+VYUqVftXePS+8NsiKvF
l7ae9vm6q0ijP37JeVY4FQ6EfkON19k7DeZH5qllInSOYHXp6cCuKUux7ENJLZVb
8uuf3kU1xuA/fpQNEL/aq0hFpJNRKS7cgM62OktPIaqGLgkHJMNWbih6ZGo03DsO
nCFotoLfzU+z9xFPAq4Ij5E84czoozuFaFGRfABV0mZ1WuMp3jrgxlf0pqWFgxOx
gqVS31SYeS0bN23BgDuLfNEDJL5WWvYoUhpv6GJbpRvk0Nvq8OGJcvyUQA9c4w3t
we/KvyS4m+N6bnlcMC4WSDXxmI3Iiy6Rn4jzzoTMurmQTMuhHnw+HOvfvoFx1/o+
nGFPIDuFoL6g1c/44jEo89KGhxB9PGN3/ffKIQrpvOXyMvaVMcxd5mfNAZg/hE7W
lkT6/WIy7VPsDPCkbrrGkQYgEdM0xGm/BsgW8bu5naEoBWtgxIkKynvX3fmzRxKv
OWCKBPXIvaBZ2uJa2PVmh2xSQLqGTG4VuCVhJ6+feMlKUFC2qbM0TA2MazHpK2Ys
1x9HJVo+PAE/NNz6N2vdAm5Zlu74E1z74uwSDtHdZOvY4UbTW6Qeh7wQzFteV0Ve
pJpGjPHWAOnNBSryU1bpyyEuCjq5GMJ5/10PlyHwsMekI2/TVFdDZ7erEz9EAgLO
pD7GdSgjwczSnjPHzZjKJrnoNQpLdOqr+SeSVW7Yhqkv6B0UNOZz/Ydo2rDZvx2U
mmjEc7g/Vnh+sLfyi1wLWHMGE3pYgVeqtOwYhJc5C868948fN6Yb730Fq2DzlL/R
8RuDfBT8QknWpZeqavYIgFLY2bFbnTzYeh5e3+CD9WxVPr89sBssgGur6l324hUg
zheuxq25EQV+4haYbq4PsrfvygRJyXLEb+cSqEcLwOoZgu4BXDNABtYWoy9vwSdQ
qgSOttxSsyUpqMwjReJc1i9ynHziJ154KmHfB5WDXYHUH46iS9KHLR9Dn9IKANWt
6t9nebkm9+RK8+GlVMwTu9Wo3+jOiCF0Fd6IY37cdQgxl5iV2jxEhkYzm4HSdYE5
ohzOoRWsbDXCGlADJ/v7PxiXETeflZ8zGeLZd8pkADpngpz9YhbSs8yCUuX0VHOV
jygM40v5if6MKJX8L+rBa4AkgM1JfrWxkmEoVG2gWZ/Ek1g7zyZinygb4nhc0vs3
OX/DfYnDExIH0Pa6FcDdGnFr6+XuW404HqvtpovqAq99b8obZ5x/NSaJyekHPOSX
hh/hF+kCU31f/YlIUh37l0z7OD3bIPlsSELqPjQbW/Dhed6fu6siov1mbKn6QBle
HUmF6dqP14vAL6lYYJWW1j0v677ijIgAgzF1N8p1Hc4jz7CpDBzsR9Lx8jBVvRfx
SJbC8ANH62yfXJHOstUl5QWCliwf+KiAYfXErH3Kgh56wSdu7ZG9QYr8cBFXPInx
UV83nmdKYXXnDsiszbtLgoEoFC+QfqX7ksRIzpq5vl0M1wCOUedZtcAxPu4ACy3O
Vv+pTWdRwJ8pVkb7zf08ZQteYFnwF2XqouJq6bS/5pjyFRi4I2OLr9zLT7hHFQb3
qPCz7alP3Y7Dd6dD7Vt+hePehFdTSVddt9hGRP6x/Cu9G9Cy8p50eszSyUZRMJY3
PWZuiIkPcFTpAME/ihqH08FuscSEX8kKVWLoeSGdwUyt0O1cRqpMA+EGNO1is1SW
vJYOlUw//ngibCz1ikDyHYG+RInaNiGTeUmb5MVOLFsofBu2xqh13/Xd4tojvN7b
/dlRFDF791NhTxcD7yGy+dg22scDU9tgScYb+vWUtaLCtA71S5HEZsC+clm/yIat
s3uVgbVhzSf/2XIhxp0COBUBmuodlCkljXluXb+zCxdfuoqItAdGRjoxeqKVPw2c
E4LSiw3Jr6kn9ljDLGpM7I+mx4pgKLJ+bGI9Kh2lq1Sy0E1CiJXD+yjRNdEj2ePT
vTheNnlHke4nz/VN8mit3E4wkWN2gjVntiK510arVEYpeLSDQaLUK1Ym3G7jRssw
WKE2JbCdk+jXy3LWESXnpW8eF4deetvcKWyy9Z9Qfbeog1ct7qL6Zc7FKpJKdRz+
qsT+dF/7EBBkN1bTZeIRD9dwqLolKQXWEqfTlztZm1K0mtQZm0Miz9TfPNs9R2Kc
5NCW0Q5OL1H78QFQ+3onZhWD3VVddUzlE9ovpj0ficeC3fH7XP141ugMKxnoYJqa
tyFOuGhIZ8Yn0nK/m5hDQ5XBJl20+R4NvDQhM/vN7cAzqLt0Dwn1hSVpAl0sFhPr
0k58FaqtldiFZgOtASEZRp80ba2mTI/OfJxpHFzRZVQYZF9IbOY1EFL29OM9T6Ju
JcpcRRj8Nh+yvEcfTA/a3hR12yuQugCTe50Zg1GZYUCqg8JXSqguJCgPjppDwJZE
GeQ2lZOxn87G0ijn+vMyfJtvCESsmXJI5KZ/3TaMFtJdNw4hWVty9ADveq8M7k6o
08ImkceRNHTdQFBVxMy4y825CkOAZ8p4e8DjZxHwEa8o+rowMeri3fzu9HzhgWMO
Y6KtGIMbXcVISWPyEONIpVlVmuTqp84ibMxWhtYvYab3Bg7o6i8Yf7ivIua/SN6i
4Qo1LkB6S0/d6DBXyPuEfQ/PRmDJd0hNblouCUqRH+nKFwr0N6Nh2PiXTVPCuKdT
wVNgr2/OK0BAljhui5tzXJIU2X3D6U4ZXrK3XKnphbzmj394eXfYk78SBpfjsiPo
NgQhnwd4aFW2Q7dfCJXDBCHVlX6roPzBzB+pkIr2zkBuZciAy+ulm0LVEvIW2OgF
x1EM5rONSv+vTKunt+7oEwurOEK5l93wvXxhSVxQvoXAf1gfmeNGK8236GBabmQT
IsyOtjhLWyxeDmYq7N6rNeqzEN5F4AlPXSVmLFxkTikE79TSpIsOk3l2Mz4bhE2j
NVWS4L+XbKXhd28M/uBt4oIdAsBogqAmhdB121vkMOnfi4e2dqNDdsqBiPZul2Dp
/0m5HgekXKxBE3CyKeH5hd8AOJKckFgsIj0XiM3FgfjM9Zgvj4eGiRuGnrOKiSlr
jUMXbCZQk/9E4OjOKTCxlQ5LrNEfboLaXlcqOsLjeymEY8C7QoB9wFa+GCAa/LnI
6wiMkzH5pDjksJ25oDVQ2MskUMhpw15V4ftWguWrWQBXYR+1T+yGgPqL8CdSdWgr
tsnYXIWhgGbSSiSp/LUhuXeR2vF5YUFNty9fFmt+jIdOOrsohAqYrTX9KfdpIOi1
6UPiJPypbRzBRv2J4oPaekRN20JFyNjR/xXAMwiTiPYuJR0+F0gz8XIoPsNqMh2z
c6bRBeiwJ1FXuhKNwjr1T3jqNT114/f3jsmIODog5+i3Bj7YlCZV4U1O0NNokBdt
GXX0sKL3jOpBwPufAokKQWm80fqXCQIxOhsTWQza/AM=
`protect end_protected