<<<<<<< HEAD:flexrio_deps/PkgSwitchedChinch.vhd
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 43504 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
093PKSQTlIpLKOLa9A382RrHnn9NN2HzKYpA1RVc+G2TQFlO6eEgyAaqIQ+BDPlD
HClqKi3GGfzc1lrBkPONZU9l00qotx6lX8A2/6IMkn0gBn3o+EoPrgg+3GxxYfQD
OrkVBZl2+bSoUc2Y63XoAIP3uoqMIL9mHQV4zgnv1exvBbtxo0CPzwWhqEEUTyFX
7CXtx9Svv9YVxCy1iAFhRekDdsgdbttjaBo6Eyevj0erL4k1GYEr1dCFrw2oMofE
vHKvh0UzRqnUH61rRJDkBHU5SYrngwLN2D3neoOgT5JQ7xGdMwb1APvDRAkkEd8H
g6BkKa7mPTYxarQ2aqQYOp0VcWb531jZ5Hri1DE2LqrDyPc8m3AUKC3zCk5gmOLn
ZyQ97bXh3eh/K24Oe2q+bSxIy3vaQ93O5PVC+L+oSx5NmjNFEUHIk+Y/GJwVhbvO
CZ+Qms6QS/G1auzUfNpulrOCq2Uctz2KlKR6wmcqlyLvwXkC4jqXFouUXIhlh/Wp
jFFtnIhDN+h6qO4OqAVLv94ESjEgJ6jwuiDBHGfdea7UgGv2tJjVsByIZBVuiHuX
CmxMLR6dZb04A0oeKB6C4pUQA/wlHcqOOBTZyGbTdaPBGi+FpydlDTwdYtLhD9jd
29XhwVDaBuasrGbl6DopzzoDocs9F4FN6yWALzFW6ZhU7Z/lYoMWwn5DJBedN+vC
wciDFXGLnNWiNr9/9eTY3TOxxUkM10CVVUeuLCkjy6gZxBMvZskh8uKEkvA1ouey
bqjnLztI+lvvtYVUs5Izz7e9xG+gAKd06Eg0Vyzgr43e6KNvE/ehb+ZKaZQj7Pak
4OfP9EZmR0fuNUdjPqaUgLbkvFoHQFOhfPvTw4a8VEflthg+crbz/wHXqNVNRZn8
R75m7eoUBMNa5lOjxmt0bT0Tjy1wGN1uLiXrKw1Ei+62HYrkZlM7IK6946cGnuDB
TeGWYB1BDIAQW7ImI6pX63PwtFD46KCFz8BIuNxP2En3oN3XyhvIRxzXB7SxxyZz
rWaXhPQa3dDN4vuENHyFzQGFPmI2xrjx78uVovskz3wBNOGIWswQ2l5SoTNps8Jd
e4i4jnjudjjRSpFOhtiehSZvfNz6yAppbLqLxd6vdHvcVb+MqdN2ASzxKUiAy5+V
vx1JUzuGWCkJdfeYK03mq7gvjHvU8MibKLH8apbya8lEYV3qMcupNgPxQTC8t3Vx
kpIYUDUbr43F15NiRJTsBFQgkQ8frpHkz8RSx8fGZBRcWTX1i/ygGlwmR9AgCd2H
Cv5kLpUqYc2OLEi2VuQeGMM/i+7GIwjbrX7fC9FADbFISJrb+qXETJFL+rtwcNsa
E4crpqfY3IDodhOb9qb8gDrok2N0DScy0AiLAcrcKSae3HlMtCsRtdYQS5DSXWdU
0bOrFPX+f6Rcmu5VXPXLdwZptGgXtAfeIsUlmT05DTo1yNJzVVLclAWgZGMsYHxe
3tCS8mfQzYs8LO4/szyDkt0TcJPp5/m5a/UdXgiqZB5PlQynngg7JRDsmDVgqEW3
TaTVqFwE1LYYMow2WCl1vTqR1eMw544s+3ht67POEyt42Zj4FI/LAjoWQnDT/DIo
fWjA+mRamV0ew5lCG4RrlgEtAd15lI60yiAXizxGhkYa6guGSxMnqFyMyolMl7V3
CT4qMCYmTVwd2hCHrrCF4ULM24O1Sb/RcOPD2+qa7LkRjYcfpgupZVm5H0D0h/uS
pSv4MACesgEI9f0ANxdR81JZPvbJE1LmPjx08k3be/TJDkhhejh1DgnLoW+Co1Zw
yAlzupZqxbiH8xjlnlwpbjKP86yrwZWcgi2IjZQmHe36pmvh8DmUJ1hoWBFQFF+6
MiSLWmvXwBIW2VOi6eQvTdTzznrv40zYPuFuV6lvxJll419BxlHDg04B2HE7Yc0R
BVebw+bYN4Do9X83d4QHXPSGJ+slA3A+0noT2RrLJhmTa6ZfNmqLoJETPrkB7jO4
+N4cUB5VEant5k+jzVgSTmcbjkj5SAiZRYJNI5xtltJ8aiXx7bCc/R5P2ro1syvb
JHSTr9PN5Lvljwz6fnsn8Jy6kWh5s52WC4Vg1dnynJst/3VRDxvDH/plAlGGyYd/
Ef61d0IwzxHYgELK8DmlkDSZua1Xa7EBqvieib1jY34/BjlCCIWZobqCG8m6alGA
z+rs7bhlvrUM53knwKUpP2uooRZC1saWIz036Zic1u/StvDsbKJSZnmQFY5cJ2ZB
fEOwgQpmuoe2xkSGGPLl4WRDmFULntrRCU89AWpFu7UwILry1/mLPBcujWn/kKsl
znVh+1ANmsD95wI2Zf/tsy1WFEgQ9RbDpAM6m3+FtcONxvcmFxxpIgkGji+/7CM/
JsIuF1zJSeypWl++RxoTB0c0PaVSG3AdFo0kVbBZ0Z25vbLBJ1y+71Ri/3vniYqb
nRSGg5czINUmSBw6vAjKBUeVjcCcNa6TiW6T+vtbk29ePZnFIfrlx06k+PF03uTY
3z18w/FIldu6dzBeyQxmr7yllhtcyJjRznBmcnZ3TM6JQz+46BSIyvve+GuRFiGz
kyvo7rMYad40gW2kMfWJIQI81Qx90DttecfpBF2i5E4HizJFqq+j+z+lRk74e6DF
ywwajfysyGYjJQbHR1N0IbtURiQhOnyEP0GgvUq0RUHM/nc2eU9NdnAk6QB8VDOV
wCRwVrDq8vq/u2x1ADGCCkwbipGRa7JT2uoIAxzQe5dGYSvfo2i9uP6sLyCB+MzN
7gBdzSXSZTAkVCMLYV6joa0INfVMp9gfa/830sRqnIn6dIL2i7MiTpGraBF37gde
jPyEdwGjv8Yx1IrbMijdQorf80UuVeWIyIrcfVFF7EUwYW2gWAFBCr13XEapTrPR
GqPm2yvso3mbbsNXzuZk9C9kf4evDgBVoriA4FThi62p/RL8YlJb9+7pMi7qGaVW
IftgiNVvuXXqP6yQubYMSeRqu76PBdf9ZVE4umyMDvBnmP9neJDCbR9hZTuv50PL
BM/cjqPLu8e7USKknT82nplb/rJZB8DOkPz/1xfrCHuHczOmNcfwNs8Yt4z/u3rY
4EEDMLi4ynTRyW5e3LgeCmMGNwVKbIWdfGVs5UlCe5p2zHjnEuqeOO8CYRYdIMqb
R7YDmJQoUk+rLopiYRJO7uWj7M4CLsvZ74hBVG2RlIQvj9IpIpYNJKzS/kZPuimK
l2opG9oT3z1cAm6wI47Jg/cKh7XPI/LIEnHyQVX3zwOv/x3xWE/+IYNBS9lcS4it
P163mgutlMs5eejYbs9CWxAlsuaN9fGbowXXa/tJNxZbpJCgVkdZTM/0M1q3p2lU
QPpwK129psTEJKLVjp6PuTwVCLAES0zzidqOBOUoYPWFlPy6zVvVJ4AbwsBpzUtk
W5l2gLlQOEZU0Xz+eHJb0Eka+fxH/EQebI49O+C0QKjlqMPpRp9/Z9AhmtHAGbq0
pRBLdE2sbNkue4yqpp1/S+G9d25JJ8uWMHuOgBk7SendYuZ14eASNUSgF/HpOCgu
91gKp59uUTSERnomtT9kfPX0dn/Ktgdc/VsXY6Zp5nNT8XMnv736hC8HL1yR1+rN
8Mwiv+orSw7P6YUBGVSmBlLe9i+4q5zy2TZq5r3wSF3atbEcJyyL259bf711a/gL
RjYBMEqzfQgxTUTeHO+EDT4Aw/LLak5ffUiJR7c1G5MyrGd6rNR9W7ECZahznPY1
948gydxCc5Cd/Hw3PB93mUxR5MQvCcjgqkHRvmXT1TttX8YGr2oP+7Fx5Umd9Mi8
q+batFHm1ME2DV0rd3caZs05Wx5crusGTPF8DPG73PELXsFzCj9blOFR1zc9NCFp
WCnSy47ENsEqNntDMXXH4yK80Oa+BHk7bVAalvMn6rGMsRAbOKxyi047zNklLc83
uldHLNvvb4FPnPgi37frthXFqQ6lM3jfJSq7gHtVK9Mz8heimk+mx8bfyuwxD5N+
TRNpeeVwhyVnr2Fn8o50mlXtpJC49sQ/On5RsEVG5FeH9VgxbE98nObX2njChFAP
w3zkU+LJMHKAC/dmu3yf+I8BVZP21HsO7pqPZ4KMEpTmrX6EHdkFcdvHT4aAvkPY
Y9gcKwrr/r643SwTf3TDuYQgBkM3WGgI5RIXVn16R5O1ERI1wKYcBleSv7vb57py
cKwh78jLwWvnEqLZihDPI2jlqrGwnwGEbEr9NkNeGzRwFed0a33RB9h2Kp5xmT+D
Bvx3KAA5PJZxTgXpJzT6I4vw+2b/x8Xvpi5jAk7Ir5NavydnKy3nCXZQOdM1d3Ou
geiKhDdcOvAOXpfRASHmEazOHVnZe/pgaZgsbD6VupO7AthnphcyzvW9LKsENWjS
CkoandBxV5beObb9GbsdjtUUbWrgZAr1LvJfcaA6XggKXwqpT2fWdPhW8qSZcAox
NS4ZseX+MsPehLtI5/+TitK/lCwl8p1W3TMjFw1RYHI/C39ODj7s6+vdSOTbZuvI
kBIaC0mpZSj/d7GnD451XRSEJJHmsX0Yu6+PdxC0fQ9Fxd8dveQRMFcXrG1eYTAs
WPSkKq8NU9lkhuFiPaqYsdfodacIL4w37D3uu4zmy21XWBFuE6OcrZFWs1+tBxO3
OroGO9iP4dA0Pv2ccFqJ8GvUruUXurIBIQ1mX8T8G10NnO3iJQGZAGw3m+B73X3Q
o2itawbSCnCyLPc488Safa4R0Yf2f9kf9t9HlZXvJsrSpsoxzJvKQ4GTmqHTiLox
haCiINSpwin4UeqlofYTgtKtKivHxk3I+JN8q0LWLsceFLvYy2OqrNyjGn1clHHp
1a5w1/Um185wtWVATVHVH7gaD2yT5m/zfBQV5O4Z733lMDtO/nCcxLa4l1DvL2Gf
LGrSqg18kO3YL9FK4Ph2SVLqQSwzvlaRejk6wRxsDNEeUhwLrLiCuUsGXPLUy3Pb
YuyiwEFI+j7wsYoJblHGRP2UW28fOKFw4QceGwxIag5TISKoMvyKRZ26erc4jb/4
cbNRRIU0tZirLN2QDY+SyAji3BT6nCUVLTiOXIyoJ8ZtK+dFDxUo44NJphcORLmJ
pGej5dzQ+ISp78aLZspaRcOMjFRnm8dkRCmn/opygAmnb1NHxJFf5DzlNP9C+uih
vxbhTGFqtf/eHtEgzaDbcSyleSfBP74OJ/dE3+uc+FIii+cM8bgE09AUEC/fILtT
YyL3on4A9pGe1ONViUKECTauu6hWBGASY7WRKmb4uK1AnVKRJTmgWBTLQxOrQ8ck
o1LVzybKbssnaXlSc/k83LSUKXABVpsI3sZBTX1ArF2kvnbN/bCRlp+ufyUttzzg
pTEE1MbJBLGSR+e9b2wyfj9UhDWMa92nPpVuPB0gMuCdKSSyxlk6iSSx1oNtJ6Wt
CuUDvGOsJcuIUBYV/Uwf4sR02s/3vOxa73wbV77jFo9V0NwtUNlWCtTwyAztXFbR
UsJ1fHd0Wp5pQgpX/WKTzYRYnGAu4gepiItWnCqw9hwqfcK2FQMt03FB3O9o7Evs
lpPhK/Nwf5mO4YMQ1R6AGsm6HpE6+ch2oqzuubExEUlycJq97lxOYGYB0joTKki+
8siBMBBwJXNM9oCIQqGHhnd0NJUHpWZL6QtU2NFY56hv6aIGyfliH9G9Oagi+57X
addTAlTlwhP+qvdKjXHC1bU2De6zwosMldtnzMtxzcavkI/cjuwiLojaKUAd+uYi
jU6P5ZpcSYFeR3C/LYKEECY08W4mnTYofrSO2gwxaWcdOkeEPtmPkBAOg1LhBnZG
vUPEMP3Upku3TpoAfNjSpu8shaVP5VK6quKvCDD7HV7Uq/MTLy5/WfTNt8m6rwFi
JR54DqwXlztOOP3bP3JvI6ki/DO1Zk/8UebuVA3G80om17+vb6SrJV49wdgrBRhH
gROeL8slIdcHmP+EiErMzOBK1zQ81nQ7P45Dek2/5mB9ilCJ3uXGHCUUkFs9zuSP
kTRkViMbIIdSN6ET0G/LpcjpmsIyi0mjGvS35AT2yEyCph3ONtjY6iZvXTmaMoVw
BLotB5s4JURIkyNSJF8FJK8fc4Gduv+6xJL5yDEaFiTugdOrpI/uElPNI+Xp0QDt
gqOMNCTjxXMLbgdxWtP74ntVgJEpYFqYSyvO4IRNSmLP0HPffVWWN3jQOmy6SVxM
oHj7DD4mBkju7J8+CCijbNdwqYUZNujQBO/b+bBicwB0KoeJc7E6n81CTjUFtAmm
1vWO5Jv0A4oGuVfVwReNxL6poC+reqpbSv9c/4yDcFNJgRnhVACOHgHU0TEO8LRm
FfwLXY6X9Uy3ibh1Rmo8Eebn3eeeyso+Bb1HHBgIUEodtZ58z1k0d0Xejvb5JZv0
/QHwqCf4o9/FlEPHah3XLcAoG8NqVmFspfeqIdGL/SYwtmQGF84IQoUEfY3s9X1f
99rQ92snTRKpLKknDLTi10uGRTfEjpRiNCQ481zKA+tgj+c71xtWIo7FCULcM1+y
FgULKEg7k6tUloIwNr9TSYR3lHE/HLLLv0uRvamQT8eo7ysnzrGsJE4GBSesrRst
VDNaiWBYcybSWu6dFu8RRT0ywNoIZR+7p7QE9AGXVqpXUve95NNoiOXN9/zY2FRL
Bwe9aBHhNw547KlDEnacG5u9XhLP6EuNjYKhyKd88E5iW2tG+gtFl545RnSokSBO
kIojioHYXm4WfbRxAm1fBAp+x71yHkiAwzMKzqT3HC0Xj63UX/8T8BneVfB1lVDL
WBDP7ziqmzOGdBak28uRwu3FXIARE4g6DTLqgOUJZoOwRpWsnMZR4+c2QD+oL5jd
60PJ6rSA5LHMpSJ9SlT+CccFsbQhd+jPMzZGEJO0roa4wddk7DoNiaDaU1UufStW
xqq4X+nw4RrdjnNacsY2GMPFbDW2/U0Q67+Q1KztDsBUlZ2a5DpxQDAOXcQ/E2gu
zdqGPvE7N18MrOTBnS+U8HT3Q2V1TuM6UjSY8t9RaEHXxtilnz6L01C0sDLRo/oC
7td4QiK/s4tgjL/Tyy8rBt/yyMzVso5Tc5uBLAE+X7GzD1RnOw9NgOx+hX/a0b2g
dZ9JlZguYQlPfd49NhlNPQTFM9LOvq75WdN4ZBXQCC6bywnB35aTZAtLhhje+rOS
cvECeVPW2WMm5Mgrh00deCZwUwTmPAqc0hhrmgvRBkOMeVQO/A0R9eu/ajASHWLW
C23P0pv8vLDoGpWLNRGblhhLqiPerGpOymJszen8yFP2hG22tYZ21hT/gbuaasXd
NrprSc/bxW0vLLntib++yD5umldgmuEaDgM0rpn+vVHe+ALhb1Aii9eqUr3VICCY
oJZ1YbVc48TmvJIenTdludAdFbk9R0kUMyTou+2GgeH4/+e8LjAcGK+jX207tnT/
TlsD4c2aoccBABzTd5tFh3S4mFWAcGFZAXdgDLhSLCJGGQ+qM1oltg1eIA5qCjQ4
nb7pvtIaAfnxHwYFmky8WG/AZhUnDKuhPshFXZXOy3ZLKVarfgVoHzXanfz4+HlH
B3ZC3kUq3BB44aAwGQdJAiigcs/cLtU9hlCTgiOEMaBKAyR2wP362QA1QB1+O75k
FtRN63C8B4iRY2lXIO9gYzWctvo9vyAjJdutxYX/+GYBebHR3YtAk5wkwttcKdxi
4FbLPV+r8GAlo6S9DxOdyACB5S2luso2uriu4NZxkCZGT4XlPvp8y1CJegtqP70t
y0Ti/dWKwPzZaL5P/xwTGCLD+5Owd1242OPtRycX4UGI9OK3Sz40EVhLGl+xTNNl
Sxdkz3w1lI8+fxO89Kqnpitp6b/hmuHWiBII+zc92peYwb0NCfzfR2uq41aL4QcV
zmtW5S6tvcxYqFf71jMfUWLWTeW8khCpdBEg/xPi7ySVyinopa9qBPVyPfOOs7mL
iVKPohnVrk3jfw0bsUsCqHgkUSL++5SFhOMgKp0ZXv3j7/JOrXLwaC3o4E1K+Xce
TKC5wYeQp2mngw0IshDyv2yCo0fkkyYARRSApWiYz4Uw/Yfp9L3edghkZFWjQaKV
0N22sKtorrTuDuEnoRAatt25sA6QyqJtfaiGMmS2TASdV7v4yGS4FFrMPfzudF3c
l5EEuw/UeFj6Fc0ttw6WRQq5zA0/vcLA2ZWtivjYhL0KD85W6ms8xIxhWLKqyxgZ
CeKgT/7754IhGSLmsvPFyGqa879fm2lxGn92mz71EwC11RkrtuKyoG9Dnurl4H8u
IlRClUpofJT7IoS+DpLwx1b8c+Sh9rKU1oXK4OB3bvtSHmFrtPJ/u4DoN524+wwL
4oiq+6OGD+GikI65c93TdCb3SJJDrLjKBL8gNLrhzu18blU9LoueA81wRzr8gy9M
n6vU6oLYec7fUz+hNTL797G4lg1me+svUURA970mUxxeFPh6dyZ7knWpMT6HiEFl
w4BIRbHeqh7KSQ8KgO8b4drV2O3q2Pn1y5/Svw5FgNT+2yHQGdwmxuDGWcj0dcKN
8jYNZ0ndApxG/ELsKfvgyUZenle9chUflMFG/z35LFGbB6BuT0z4moENywHJ4Quo
WRSaZrO6+dcUhuK9xKdXgudp0BwRBWd3XGAZ5ayudHfDXW3FQzvnbPn3zIBvZ3Ed
XPnjK36fkQq0WjYsm2lBTN9CRTpYJp98ycmo9vVz0VV1TzPyIet8+5RZgug1F129
AaETCRz4GTnJMocQjauALjt2Q3bdKLno4KBRciI3Mji1+HH9O89C14tUBu9cuYss
sPjng9gy8EmsSJ/2EgdogYaa+dAEGo2iOYlwG3EWMxc0XERNa23W6JAVOeb9qpLf
6ySSe/ZIwQQRYn9uij/zSvOSwjyHl7j2OeIjAb+RZuwVNCNi9VkfWZO1V6KyNrT+
zHM9OiadmyCaxBQR4M+13QGUW/PRYGWQYstQOI4oD2uS8/VMbn6hJGfouPPDPpUP
ENPW24nuIkjdLLb+/40/nk+C4J7nKQJjnPItF+SnPkxXJKuJ2fpJ9EymUaPfliDy
4wgdsxtq9JFygaw8f0LaDf73l87sEHduKR5Ua7O8rbVpyP3KeVvpGB7WDtMnwZ8L
Jtliwk47MkQK3UKxIJ9w952RiogumTEwCno/+zCwhglm+zSvmTSr2JdZk9qeVGcf
dwSdeo/rLJNsIf1ArsLuu6U2iUInx2EWepDCoeMiY29xb35SS5HiP+ZKkqrMk6HH
i33kbJEPFi9MQgWwcu+fEnAbYR+cXILML9sdZ2hUS/ucSl2+evEuhMZI+wfmq4KH
Aur+O8wGCVWgNj/LoMnCHHV+eo8W6S6ByvQbWuz8kfx84AiykkMyAACCYesgHMxG
4Qgs1v0sncQjBPSaWkwFrfrfm0setZF7zGW+PyU35U3CEzZqpT2tCDMliZ30jS5L
xtD9WtTmN6ThJ1vJdu4HWnzuX9uk8VH8eAW5oI6Yz5fTvQXy6JjYViObPrNav8CA
cdrgtvXP4t7ecOIUp+6zHMd+3SB/QJ9xNdeNktCHk8BAbIxWCnPmIYRdsoNaX8KQ
rh35/eVPaFo0oinXVG4IaSBQAXUg7bAbPDH7DoWJCDGikhY0i4ahGpWpng0VbkBN
tCLPUft69Fy4jEh/cjd6vt5Jk4RWRJXTLofhy0yjK9zevW52NOEwSVoI5ePbGXIi
7UHAMnFh5hKuXBYodMNqDXJAchKF1TJDHwmAhaoeBjyVhckUe97XAq6gx1e0I3Os
cxD+V/hB0Dwg8WNs7t/lPmEw+vGePlMMio3jkD54IIYgNxQY/6rYafO1CCrp1KVE
N0F1MBKDvK/tGFQt7/yr8/8jdWisSadxiY+xy78e9Xt8IeA0ghZVSOG8uKyK89+K
mfADGoTgPmMEtkvR4b9Us4fVNxgBASiXhuKwVrVrgQ48p7za/ckvgjffm4UgyJ/f
2AtrevtQauVl2bx86EuBXQz05MPMd0r1PsR4O0a86boYX7XX8Nl2rJPRfqaqXDbZ
mVMuExD0cFBN639faXz7lSKq/DIlc+pAGU9cChAf10TvqUoqVyu/Uzk3Eokx4eWh
Q4dtyPNsls7/Al42RfJIhwOTJOhalpGQJ7wL3qUvGvJLAGOsRVkMuf1cL9cFaA+d
2+MSKjPBr4EGOLK7EM1nobjq/Ia3zPrrRCJ4zcSwDNKhbP6tKpwnS0qlyEBhwdzk
AuQZQ1dVmdBYDr3M+XMQZ6X3WxOVlDKZu9vHfBWHKKISMJEDuDjhrGdbKgr0RBVR
mcxs+fnTJnBpXNHbMxYaQxAD6/jTrJsI63nmD9KRXLwrZ/QYwVWPv/vHkcV/nWJt
S2ZjNSUQ98JwfsqrHfgxf+a/9CozY1p15VQXbnOLbmfbLiFfF5Um4NRp0y7YJmGw
ctkrgtxr0fwh5KL7bZro7NfIF+LCX7D+v0Ibgg423H3EZ/Gs5YTPTnNKyY8YUIMO
W68hfNezCB8vMNDgmDm1FHFgzAE8fe4FxBfM8TSDds1zeUgUUzXWrWjOKumJBEyx
f4sO1a+4oF1EKiYAG4pJaNL5TrHonZ3IYuGn/EXc9HBy4rVoqgUEwp//HkiTaJnN
ScOy8wbAc+mrglSiWboXQE+MDgLqOPfg5QoJo3rTv4v80RN/Zhe2cpVGJ1STAsSr
yfzbDJn/dzE62E0egT1xIMmRpmx+yGFh7V9YK82ZM6n5RGJJkjClPO4+T/1VVCtz
X1PJcaQfbWrCQka+nQr36LR4yoM/8F6GqmKCA1vb4KmvVhNGB0CE9/WAXi2HLlXp
ZtlgAomR0pGOXI7W7IpQozYZ79fV7Llu9HZthAc4UN/t2vR1KTyjGASgmnGzplLB
x6kEhwPAPHTasfqLmgkknrXZzAfVOQbwo+syi/AT8+A/h3GMlOHJzv3d9OZDqXHH
uLE+t7bPAmBYAUHe97prr143vGYgkSfuWHhUeMK555xWeGuCaXQw/hfy3cRhrpS6
V3TCfHZ/jVCbRnAYm51SXKV0JTg0GhEPnJ34Zuc0aKXhkvg7e0WKqalC7+91Qtn2
cVf9sgGILL0hgzIhX+Pf2oURIzQUS9LqTSQaXScPHNRw+zofzI9o77EHLv6bhiJD
MIrlpD6rmUOQkkrZ3QwMvIfYVxRcaV22twqDfxibOghw0QthZQCxb/Yx2lrdpb7g
s+0aUXvuxyZl9Q7RLPi44SkkSTPhFknoG0TLhg61MBxMHrNblnzJ8MyZ0uTmWJW+
L8Nd1waRR07I8XbMB4hs+bewSakjzKFOSCjGjogQsdNTYpjctUcX2sEN0ygCD20S
Okb79RQ2zJJRd0gGbdmOgSJ9u9UWqhTsbaQBdjrlKNGdfff6sTnmWyQ3gwzYAw1i
7Jrgfg1Kv6RfiR2Aq3tTMbGWudi8zJOWFjumFlCp4LEpCAX2nujCpdlKEvwoEFCB
9UASmFLFP1JdbX4rrQGIRYryOkLKSjlzf7LybS9v/cITzZk0s439r/KQdtVIZoTl
neFGKEfxVzHlagPJkhlnYLz3x7lSuLq91bu4d6PWPkSkYkedO5zAbum9cFFkGl2W
N7NSrDtp/Gtj0TLSoPrvUMOsplEX9IsSBemgYuxdXVgjgm3sXR7NY0u1EXV2S96+
qJQ4QMvl4CsZLVpNM53wV/QzLmMqxzfesD8RhFFSk8uEaRN8rQOHMEHNrI4vIoYe
SB1TU8Ne2cuxa3oQTqpnHzMMuDpHCvWinPBW0DWVa+AZTtLofLxvS+NEx1zj47+3
TKZ533lP1xAdUj+42YxlDzVOP5+n99RYR/5O48eANGVncMYHDjU0OnE2lZpye9Et
Ui4zLjREWYMZwaeomQ9X7ctiqaOTsYA5vAt21q1CEL+hgfC3AmNovP2IViws85kg
xJ0xgoQf/tTpRlel+cQzEDquV51F4Dxr3PswNlR1bIBMvvXcUTc2CzHfUt2stypE
ir4zPNKbQRGCV+868qG+KWt1pFDmU7VlJQH1OZjPU64SRJ1af06W3zHybb78qk1W
FSxl0H7yCTqtc1iAHFy7rZSFgm2IC+nNxn1Nd28q179yLVFpyf8AuTI5vciMybI9
s1Rpe/2MJeuw4ICK+HWFqm5m4QpFga8Hi6fBQeAiLXfbGRPE9gE3WmZvYAzSe4mr
vLrVYGomnVPsHNSPU4llRRE5+twqH0QzjRzZKm1qKnPAfBNMqoVXG4wlbK+//nq+
bpgpWUF4RQBdZGY/tJbmKWVMIM0fGVDRsp0oN35VTG/K+xSDMDWS7a4p+ckqAvqX
Upi1JYcsyvkVbh9mupKDt7BFJdg3VvNBiT9KqOk/c+0ZNGKXZ5iyBDI+c1IWKier
yXsK2tkE4hhKD7yjteNV7vBMWYSTpPaUjOEG5DT5m+IqRD/2N/FG3WIR3e05M/8a
wplV8i7UjwsAKegE9TA4JstDMvx0HjE1n2sR1SfqCW0vz6lN7zqQk5LeyuGI0+KM
D63xB3y0d4ZGO/qy/ZLpIYdTarcXj7fdrGprrpIkgK0iuRRFaM/6HTSFzhOGxBvO
7JLIkZC3bEY38MTc8AfRe+b8ee4c8XJYLEKFmhQFaVwZ64wM2KnVmwx2H0dPQxv9
QEAthPwewCaGZIpHRxzqIVYD6ASfvuLmHIMlQyqsqm61rVjFlgtLzHTzKrm+gNNq
OONJ1DcYDSpuy7XDVbIOVh5kvM2qM0TJ6PcM+i9LGchFyxPKBMtI4vKRaF4NcGhX
oDMpLflfuZozM7ILIcTWEDMMZbv7H+bAwoAj5zBBHn+7c6qko3t8YXE44tLhUEo1
RRxO1SVkfvXCbG53W1QFpjCkou79omMkUfNtTHVpr8KHhkD4wK0AqgC9AAnfUnwr
j0t5lPtP+1iJPjIcADEzbNC3vM/njsxAhqe4kcDy57Nk6YYdGiErR2I2Bmtw96vo
DPFHFatqnX8baiE8NNyk8dzmgbZ93y9hjzql2b+PREy1Rx0DUgSFSRwXaRtMJW1b
DElVWCG+nywIj96lie64dF0pepUHVegCxYCiOwGn13xv0SrZgG2y6M56aDJ7fVMg
uNKoygaTM7t4iZIHYblvLpnHdVsRy0jX+T0nN2YkbJqgo0NiM1zMwiBPsQkeXbWx
7FzG34jcXEIBkKpaG/FJfcrxRoWUN5GnOF3qXHJVR7o6QuFgPUFZ1WMoyHRudTTA
LLrqeOTaWVwahK+hoPsGu12LKRg1KULhpfJhaEYnTk/8PuIRulpmIVdAt92JT66l
EDi3KFV2FoGDz+lESVaVqkTQiLWRDIJrL7SvKRe55i/g2AeWJri1VmCrwONhSq34
IT2bUc5YM+iy3r6rYbb76bMY5juqJodhyEBvNQnxdrHrrw0J1ZqBqiDE1o9A3AXm
6ExmTVf0rDYKRTpY7maAF+lwA+/TueX2emZ5iUfI5Zad1oGB/9Ir6gAGgXtngn9F
WZH+2aII2788wWUI4gIuuENk6/ZLaphE093gpcuYIp1btGjdreTE1DZWdVGU3IDB
j+du6ikWgvduWsvTCsE9hgSTzlfeES2STdDc8dQeVWRiG6ieXMbLfvnn0RUS0eSd
HAZPRH5+4Le9cCRjExXTBLyamQnIdXhJ4D7ljp6j8x7lUObTuGUtyaDcVBOp2csx
NCQiJv6e2USHrVRo3RFcC93++gf8B6Rr8V+2IVWKc0SlbPI1xAVZkrQl6AUEv2Zi
tmvEbjXFr6EB6On/DrwYdhRa8rbrXg7omz2o3aI9/96poh6rT0vKjmYgSHEp/XHn
mqn2tP9aHi8/2qQUWtpn/9OpE6pzlaaqSH/tUiYYuWUiHC5wFSV9JvOxMJqlCxr+
D9M9SxhAQVHHKyocCKOepu4ei0ubmKadPuOsdgoh2c+KUyiP7lUzpSkPxhR4+Nxt
aadb0M4FUH2Msl5GMhpLT/T7trWI24e/ZhvewGgrC6SyjAZ4dvLIGugl3R7C4BH7
08yGPbEsGK7ZHXlzfaumlz6mvlb3pcNawQ/w+jNCiN8o027D8lMpqSgN1t2N0X7U
JbCWZZyQm9WbzB9foTggZ6ARaUmAEIxVoXHe/Wz6xJ4gMdtCMCR2ld49Sn+I/N2m
KoRr4ng0dM1of8coF8CHJ8Afz2X3eH9p6iAXzW/bpD/CVmpLxC+W6VhQmq46k7qU
sCloOieWMmj6kjfkS79vsxwCshpwcLAh/Z6XVNmvm9jzVzl/qkfO8Gvq63oOYx//
NBERChwl2ncAyP8oXGrNVWKY8OnIO0XO3BL+4n8AKrBzWs4q8/zsTQtg64DRacey
cuVVc8GnEjVZVvPas3UumVU3LqCUQAbXm8KFxQLut1fZzktmfyD1zMcxwgRB0fgQ
T/N9qss7vzPKXo/9XXVya25C3P13WstCSGcLrM86yezr1mUAWc3rAmZ0J4f685iv
qS3LqVLedbLOanL/2mxuRo8W6YGcrCfpD/QZqh/B0sltkP8NO2R6jOjVcfxV3VjE
A8420QvJPJEx2O2SMJMQWyQLsKDrdyD97pAHHNTKZ4uBZadYMWR/+S8qJ9NIUx0e
QlF3Ul4GetpXCtkxs8i/71LZZOo/N79hBuZvqd8dHO+yHeosCOhlTi0p04r1QMWp
YpV64/1ppeyK6pJuNmp6pXyWwl21QjIhWV00B5fvWE+c8vQjE1eL2HSYHW/qeH0h
uEh6P0eGGCiPK0AQxVTlRDhVdnf4i2Oapt4nbJOkXzmiOI8xFJVcdOExRqEog0XY
4qA/H/RfJCQnq9bGZCbmaveDBeo+4YmE2M76ZJnUDRDopC74eckXcPQqna9zpRJh
aSEiPnAxVLgYCNfug7joFo14YCdXs4iQLfwadREr6Kmf0SIqV5MJ0Xp4fD8FckSR
LSbNViJUn+ciOK1yjYFMTs0B/tghwv7vy5OyMPXHQ2GBVJgjTRa6Y5fxB1w/hEEW
wM+sfsCP40oD6FWxmXi5lrLFDxfhCOgjeqfG3knSVgm/eFJWCbJDhorw1gwCtfON
VuBjVQCn/uareRZCYZfgypTrcClgHcrBkkJIhUgqDJijYtH0FxiNn4ZweB5zlO7G
H5mjoyaaSBnLp3OEMG6a9htO3UfWYEkKOAZxkmQk1OuqU4cfOuRshA1nwmQI/X6M
oUsPDX0cU0gECULfylnqqrwD3ZO1+UuJNzZERbqCZlAMB/foggGEYfyn2MZBezHx
NY4lgftnCmCYSD9QXwlZ3czx8P12FRU748guxVyyk8bBjWevW4NDp8B4KZkfqOVd
7LXOQ7Bn0QH/qdpHgJiqT7jYR0Ibx8LpHHJwzmHrvJRFnN2IoZnf0sqoG8nvk8p2
TDz/8hpa1rWcLvtNTmxg7/PSS21QK31RNA9xtoe9AIzJXyVdWhSBie80QWA9NTIo
rSOR6OBlPFJW+U67p5YYe0qD3tjXFzpr0v5wdV7BJe3THsLrHsXXam1cJ7dqjFY1
hasNPFiylBRBUBpjrEy7hDIi8nhJ+Uqf1XmvqjvzWlV/9EBq6s1YswYeQUP8rmsC
x/0TH0mmOhrL0W3XUBTxMWUGj5k0tDVWFeqW8NPTFfugLQkiBFcAEN2K/TxtQ60r
org7RlVzR4E1BdTXyEGXJwAPNxE9Cd3bPZtDKq2mHbyg61pscHAejRR8fRbQ2LjK
plgUp9nDU3DrPOD6vUzTzR+rl8y0UwbaE5nlSZQKE/+LFVxv7p70CGMrmCoj6sPl
CmXGEjHxfKZVUOcJ05ZiVcd8uIc+rqm/ozPkiqHBenWmKts+gH8tqoX32Bwdx44M
Ce2dtlFzyt1FgZYJihRg89l4kn7MbQR/JuX0HFYdspVRydS96BHOtjVpurVzqkGX
5QvWO0F/xqxwVHtSYFBAK1JJrpLXJOh/T/GSjlidQXY7KXKYDgaAR+VB6GzWeV+O
FmR+kKiaPPoSKdWJh6pwU3KQkFak2WVLkCDosPRMW4X8O7mVwXI/xDPufbjZJ4HA
GWpnrRoEEmEi28cehKzkgYnwHSIMCQ3n+94mS5i9laTUGP7K8glRXWhwVl8dFyPB
mPHS2GSLeDzms5jx0ju6f+v+vOAxjsvmJ7gPqCszMZAEESlnUgQcIkCPmRvrmVxf
686fCUl4oX/BZ3G7CNyimQERHfcG9+NNbswyDr1KYTtUsZWhPED4SAQuDDKw+/OR
OsMpc4GVZYcXRfIIkRgLueMAKqtk2VCEhvJndr1zlWftLbOGxt4VGWqlEdaPk9QT
7tlWu8bHRxMQaCJzjAKx0GR1SRupVYs8wXeJ3N/7uXO287YTftfHDRmSqm4LEYMh
w6tEL4O7MQKAdIO4KB1AV1CpPR232+O/mte/taFhVIh3ILpc8MQbqRnY4PDvK9co
+UlmdbYKTK2/y23Ve+96EJmXA+Cdq8d6X+ayQxhoFYdU3+eiYSqGLUe/kSuHAk/y
ITXeWoJcYhBchVXcL1bjkXwHcKhICUGLpmSAn/1xdtZVgWSG5RVts0UgP3GwGmgO
CyDM1ltk+ot3SFhhGzQMYZmu3bF7hBaRkO1MXz6kxf362XhINbvXZPmop8+lixv0
aesGJ7w3NhvotdpR1TDPkw1wfPaJibDvfVrVoZdTlOGnFaY5A9deWekKaiUrG2BQ
8/vPAm9Ce1oq8qcCXChCRwotmZNMgmEeSiRgmbc1TxIQL63Ih243+wePIwJxyzU9
GUCdMG/lzZQ1Fn1BVtmwLMHI1TTyXnJbSOmle/En6fapQVqOnIthGHa9YVwyidmj
CW47eajU1j5LVkgzdMylYw79i5fitgksgHhVLR5RqMJTeZfeoxdq6vzanuqZPgMn
oIQJInhOCSzoxG+uAzyNXXw2QGLoI1q1hScW1J3E3T1UZDw2Kn/vwJkiqimx0dFx
q0Wa1OJrf0hgNPlVgW7yEvlvvwY8rDDedemdeDF1QDDc3u3aMj024kN5ieCdF6YO
ssVRLvZfzggn/2qflISF9vByTdvpb27xyJvth9gVfXinXEKjJK+LjOYk4Nvmy6u8
Qysf+BCEu2k4eI+1mFkdVrxXcmujXizevpGm5zHvb8ne5PwckhJwxgpq0op0kq+2
s/+FFeLwDJVf6ZTiXQhXOTrn2d2HoFeLLFhXYq52LYvOw+3YRawilf7nF90i1/dV
K1XVHUjoPkLr9dub2ad31O5AkENOvUkB9k1qMaPlu43ByhjDrLrJqFmCpq0UlRpr
le+K0wqNG3S2wfSPdwg6I4Mjg2uOB9RbTTqbbyjOgCNV+r2idRhfCLxMq+KPTUCo
TAS0UebfDwyGRufkvONHrAmLaciwsnRl3Ih3ZkY5UHyhdNCyX18fQUURe7yXGra0
7aj+DrhXYho8pO7wmAFymj3ZUBE1xeKbiGFCJttbp32pkHIu+Zwe00Oik3e7Lqeg
HJlJ+4nCpThKF0DpB9qehcn8aqFQugP4ILNzZJY416u6VEuqCpLIy6jo5QGFSPj0
0H/Oci1v8Z3C5PuPzzJR4CgZalhWA6bD8BXa2cTO140SGVHO9aFbRm6YyswsWI1H
1SKliBZsZUtbc8mEBYh3TzbQuZ1gLmglpS5ki1e7yJrAM4oVV8GlDPMb8P4oZlJE
AMfQvyAR6KzEgmOmnsPABNotIQFz+/SVOLpcdhUOGyPwSI8uTPFBbBif1bxx7VHF
7rG8cL4MnGduGfex3NEnzV/LVUHehE6+scQd/63tXGTYzTv0jhjdUjtzLAnSUATO
3DRpPfwvg8X8UCxSyFpasyKoyNtCmVG16lrJmx+bsi+X5/8XXWfWzwu3BLMRiaKN
x+LuE6IEEYGj7ryZt1ju1oQANtxjBVtudPK2QHHn4PZC4U0K6dBtGpLv/qGPUL6i
WLN/nDmRN8kJfbtnyqPLBRXYAZ0COiOdvsgkBjeHxNesidp6r4ei59YLNcUt2YkS
1yY1Wnvd8xJA37XkihL+sdaImFfUFkJT4v1/HvU0cZvyOacXi1bs3UgPaUhttNK3
F4fYkJI99OR3EJDfyu+AUNGTjrTCrcXQuBdVsk3coO2U3MkKK45H8C0Ryj6q0yxz
tjg0Q6DAnAaEP7mJSUep929Xew7Nuo8Zh00evvmjN/5ptjMnYcAi0bPLD3LrRdZo
DROTE3Ax0OBmn6bV5/WClq3NpXZiImJXzN7bX2NCa1diFEKFijrSxOz63hMe90mQ
rOFCT+ulmC1D8K+V4TiwRYzWMevdv/bCeQjSi0KMwUBTWDm11UXDI5m0eMc1mohZ
Fsw8JLDi3BcmZ7/KNV61W6wcwVcSYN2cM7Q2Hlhuffg8NrjpdXYR0/r3yUiS9Yt3
FQhK5uqKouI52Vp66plZYr6vzMNTJMThtzIfljgvvB9v3SMV/GKeP5rDuCQvFvDJ
i/xh1F4eDovAUzX0mu8KtCmK02mCdGyxtTdsxE6rwgr4gv3oUGp4jg/DnInhe93E
pCo8fVPhE5+yYxKkIW8NX8d4HKIDjHGk/yQrmDv6kcE8tX+zULSOt1cyrA3CWtKY
P5Yp4cEYlJLsCgMZms241oIsiNY4naa2Q1mmGym4d6VzetZxRIevR5YZm6/hBEpV
EjSnUTo3/QZNriS/EuTVOitUIbeQs2xuMSKjNi3NBaN15QD4REIjYF+Nqyb5cYhQ
vImAuJTUMlm8MoD20Me/aVSxE9/JLJFCOxVtheBcUOwl/KSFJ0kZkgsOj5vK2CMn
svJDD4KvFsVfc32Qwh8Yu2hCsS81PQTWwl9cfR/33FAKtVrmg9TYkglsKlbgLDxd
0kFfQnzz2Kfwe3ZuRX88awrYQDboVzNjJcnDCK0Hg3jmkHThRwTENYl9rzNPopPb
B766VEXQGHxr2j04be2h1D6euprRn7JwSq5LXndijouYyELKvjG3CfJaYC16DGIP
WjR1w9cuYMDsTAQRzZ7oXR/ZeQ6W3y0O0wScec7Zk0QCvsBwHSMqDncofwD2vHnJ
ej18kgP6ddbEDljCgdcigRRaCtN2PLNk3gklszskEvx8YYQdJFm9K6syLSCtbx6T
O/CRYFNYKv+XGKjeJVRrNk5e7YDLogT7dRDWU7BOFA56SG1wWKD6oy0UN2NDv/Jx
v2TxGis7tGOAbYSIVtO08fSzz3Ycrnm1VUZ03RnqPz+oJFHsBcxlGcHtkXVtRx0Y
oPM76Wmb1gZAVJbjYDynFk7GWp0LM0Pw0BLeJZvbdBMuiwxdfh5k6O5/cI/DWUpS
gxujsd8+/RdHz3FfXoyUp3DSmdTVaaC6cN3ZUXbFfrTmQy5eNnd3ty286Wrv7I0W
lv3vJ62Mg0zqcZdbolKnQBDKMC6as7a/E4c74X6c2rKPgzRJk4Lymdu4XxZBYTyR
rMplcJhDTDkyqjg6o5Ek2G3tXMRV2iLZbrqKg3NUenfE5rx3AkwBQ0j02m6OqFap
dRGBI7rAd3yPu5OlUHnhvNiJBwZ/tj2ZZ1L7WpuOoTxO8enmfSSetLDBIqK/Z3+R
cS6zHwAZU+8zcz9aexTEN1/3zeOVzu6C1/pnHNE1FBP3lvBawUxC88VAqtLDfPj5
zgmj3nz27Ur47OFbKCyVWT/PkyWniA722axy8n3On8cw1VwzxbqTuiZ2MU2L5vnq
nbBtVMIUeYNsOAP9N1I7CJyiZ3zyeze552MYRVa3AcXCj5V20f7i5E9tszRQt1ye
VuEJFM4J7PSJ4YzTlZS+DnR6u63dhhmKSh3j7pV4JnAhLCvddJjfmxGtaZoCsfnm
g/K9Awyj2lKOq49KO9hrnAY7HYUv1gprdo4yhU/BpkmtP9wk32goxd/sqUJ0k2sX
lJzeDVGR0gxdB00EQ2LUQbJhDaJeNlpUr9BWDX3xu3ea05F42Ez1BLdAMloISEaf
KTspdu1CJrBid10ZepORHxvMaDMYaYSNjiuT5z/NPzNDU0HjWZs5GSp5iGEZ6EBb
BVN71eM/0C/1bcMIUODpHlVXQE/9FfMZ+9hqBALTt0XhTk2txQPyPQhTm9qtBh3V
bQZCvCzy/hFp+oO/UzT9q3avJ/hKge0vxQZmm3IM8A6FtCouzwa8VIgVQYdUD9iX
8TEUT+Xa7aW/7jwrsascuwvX+Ijmfer6tYstWH04KpntQrmOo1e7O6wtXcQiYPXy
KjzeuCUXZyJo+hV5tzlzceG6fRPJ42oHKOszdGbl9uXOjYsV/sjm0LmS+7iXpfO+
/ZHkNx+rS10W8yKPqoojBEB1gcQMpIRzH95++JQlrmKC/Ipr61zu1KPxj/f4zLrm
WntdKxT9fRzAyJ2dNkFbtG323h0wPX5eUq/Ms5SYWTTK24DuOrU3Walwh9Ic2rh8
wH+CgAw95IERbUoXv9/VOgChp4tyXUgXyRU8k7n27grJdIqHUozeKrXDZz4r1mAo
P2brSAtE/04cBrHiE4m9cQWLy+1SyWhqe+e2Gnr1/M2JQ/3oc2j53yTYZpEuG7yj
bcHXJkN+OxMOTazjEu66OHwQyd6L8z628p3EtK5kS9e8v7VYHxFqQT4B5q1hRFid
ZcUvAigAuf+/3zzr6dqwGBuia2Di8SXn7XqjC9m+O4+soLcW8Ve77sjCDfdVL1S/
tZbI5Sd/avZOEKzN0gEtUKkC64smFeO6gJcq8BJGUnO+0Ib1S+H6HJw8GPCOhvB3
p8zZV4hpjx2s6IXj2QyneGmu3VMODPELWoig1VoVvYr8GJcL8DsiCywem4JHHOLc
y5005S9iC3H0Y1ZlFwSXoBQh1ve6TKdcSskzCeW6J3NHjZC9yeojUGrpmwp2RAHb
xdwFSXJ8aykAoj6qLfO3TudYAsQqZH3ACQg5ayg84nsAgPvSlPhGwlCyhmGytFgh
9ATnALTn3ws2bzxCt3y2qou+cuoYXpKhTvVHCZ4rWpDgWR5e1Ka+j/GEvXAyn+Fz
N3MwpUjQ7coNOtFyUxxgNyCS807NNh7ljfYuEf+1sosndj3x1fOQzdlpvdJjlova
MPU9fZAMiSD5POlonzNZ5zdwPcrSrpHYTEXk0pnDa6p6HUokzpfD6R0i2KAx8Nt8
2gJGW7nPocuyEhkcYnDM/4858fYpWYcvdGDxr5VggsVsy0v0hEd5GBL1zSzHkq4h
k5lj27hhMfryLrXyelU+8Z6zMo2B3BXzq1d/gUy2kBBupVs+w7ZSgN70aXbJMKMY
0j95epuDrJB+Jv+9E7kpN+6nqhOx1nP1m3YvEgqSBh0SNS8ikCSSX5m91fzOHKQk
Z9VN45rS3aKBkj2qAnez3sjDchim9THwnUlBfDFat2J5tvuDYP1LvR3RR8Y6NZDI
LmI9x0TMb+hJoA+c5zfdyJ1Cpne2OTQsPjIZzzyYW7yfl993qEW74NqpkSuwE8jV
mpeLqeNwdiovkuB6XtfOJtuk8E99wjehm1R9W4gsCVaG9nM7Ic81IwjneIJ9Bo15
lLU1XvolJ0gWoWH1C3xVFdINN5Qa5VcNJWfSkSlt5ZEsnDD7qmc/PBU/NFc0TKEx
arzmjgrPo0c3ghJU5cD0cRkokdxVUzml5deAoiwawfQLCdL4SsV54CU990Qpbn2l
yg2Qws5OsVhv/xr5n/U/lVGR/IuEKdqigSWWIGfbc/W2EG/N7eMTGAA5ulcHSqKX
8QPjJdT/HSzUsAysHhgB97qiBnxjs+L1+ztPR3oL80NDfnVUTwl21IYlv3xmUvVk
rZDDwictG38OftSQJgX+wl2bpfMMD1LaBcmn59kKNXAOa7KJS8705R7zf1pDBsZR
gFg+GYPYhn/Q22qLmlVmDcINdWyUwcRMYjunesGfGsRhpCVolUPjAILRuScEMQKQ
gHowh61JRc5kZqlmM902I3aHPIA6J5iF48bq1fNptUvyVMDIZryqlRgSNL9aCYt0
op74iGF5zv+n3S7QUdRcS3l9hpO3NlGKRSkJnMFaQ1aPkp+1FaARP1ezmoorXx1j
GqHTKwtSD3WeUZ0DUe93/H1HwsqR1aEUZCYGEJDDSRvqMQBkCz8yMtyV6h7qYic+
8ZDYiGMlN4h7LoO8VvAf0H2ttQcj535mpN9drSmpJTtUoBVX+6c5CO/JbSNKTbHt
i0ZdqfvQnSKsKVtz5pXSa+c00uA9iV2zViGN5DSrjzBQHDzz9FWyxTp4AG/FLtcj
PcjSnaGzhYHb6RroksYdraiocn51qsiltHGsgTGU0JFSAU1IYMz+LLoffd81vka/
uMV8H/uhl9ZI16p1egWEeWXXX5kStcasJOK02espmRS9LG27gsK2aHpO2Z8jdetR
my7mr24VVXU7ZaLO4m/E80hxdFcyrr6z9KVfV99swHW5s+HeLRyKQ8Y4Es0E3ySm
EoxrcEY/vQj8vuod5Jrn5yagwobzy7nlCmIRgEBgrBSP5FJSmImLo3ovngU1E7md
DmgS388rMu7Q2bgBXHsGe1e15ugD3KUTq5bo0O27G1ShYg2vRr47OnA1pP+TQn+H
nzzwbqP6Ooy6WwNimXmpTyMw6TubA+I8epU07VyQ0KCCvEwAMy7lV4r3ODBMJRzl
wQ6+W7kvbXMuYUnRFmo+Wxpu2G5xzDeVmz9gNUdolJFvW0Nvr+ASt2WV0LqAtUav
CbBqdbxMjzL7qnXpVeYK/2uRdI3TID195a4Dtu2CsEnH6BonQG+VKeBSstrLb/W0
u0lfDx8lNHLqBSJmeCOE5rPlDMH5YkupQo0Tm/M4r1UkDwgI+P+ztiCfuidht1do
X8lqzsPsPoQEMOjeITyXswW2UH/Md4Q5bzLB4MY0K19Iv+P2tkpt5M8weXq6+Y36
hZXFf48aKyZ2scd+NPo/roQmbjXCvjf2pK5rXXfRuFz+C+fglsTAWxNPaaTV2N06
6dVw+AJpkwWqpWyxSQr87nKBBVjSqrjHOoQl8QGFGffhMPT3I81MWnZ1DtXfmHih
5qdL7/TEBb9F96w2fdoIyIIcv6Jbv0IFIXqv1gdTGlRyJitqXGUPhJxWxtXZGnOy
s3mMFaJwtLIJhj6cxx1jhI9TmKUtvG5qUCc0Ck8gqTpTb94/Sy7Hv+yG8+7dQNgF
CzQmNFO0TbiZ9sKtlESCXZCxgGIDVEvaeGk4TKJcanz1sKru1p8J41QP2k8tzxhU
oItE+nUNvDKyEXd61zRFWxNlR+ZTm1tBaEpLkq/If/zaNWSwQovPGUkdJHJWrWhd
w9cDzkm/Kq3vgicxVPICJZxU9KxR7KYB/HzsinnwSJW4rwoqxPF3d7tk8NhrbCTX
TJy1yhEfTQvVPHybEvnTzxXCLjyvs0LZsaxuhsLEw9ZyO12fRDrFxzvaj5R7I+6y
tMUce2slzNB5Sjz3j3hWPHsjT3rJALREOIZmlJbWSzeG08+qvsrRkUYsKgBkUCyk
Oy5a1t5RiIIeJSOpWFX/XriOQDlclzSwAqclPj6kEs36TYl1kG4kF5228yj+ltgR
8oQK9AxavQMIkNgHFV9Ws21uZk6VLqGzNpAmXa38W+k81q1AR2YlJMevtusXrkrA
xB7sT3O2SMVMsdP+cl2FPR1km2xPLF08zOosD7Ay3cMbwZYwURNR23nUECLbUGne
C9syp/HJBHWKrUW+6NHqB76LspmRDLUK/TK3kowhrAk7Fshmt+KoV7gWk68zOihZ
SsIA1LYXGhsZzUDQSDrfNCrhzE+toRdZ2f1kHAQbhGI8a0j9e67tgXrwyiaxd50p
3i54LvGPJG0VODPp07rLWabCV1l73U2V+9R6ZaXIziCREL1J+YsCRT4+lnSrR0jH
4Xe36p74AHNVcADGiSgoq2M8s+dtAokJynafFfsNarUX8WSIGoFXH4doYGb+g33H
C5zydGwC2m6mf3tQipgia38zcv+nXShGj0eRQb6lTeAN1+km1ySoruM3PLQbI57j
qYEyue9xJhSf15r0xPwRE+CVMorWw0jKz9exdR+/Chl7voDYQ4UbHkC6jMPcUYzo
+rzbCZixm6/xdpG2+AkLE93wnfwebTtNhJXMJ603Ow7+A4DXFRmRkdTTWtwyASOn
AKxQww0BI36im32PgcP8H9O8vR6OWnTQWwKECO+AmqAqqYBzNSWaiG/bN0/S3YzZ
ksU5BhmV9uRSmFa47xOD2GPCe50fgbJ3suK3BUeI0C97dLaLALVlxzvQNPcK+LMg
F+V2UETr4D9w4mXYcJJGL001tRjFDIV/7XclTyOZFYlqH2g1XVsGKAUAZKFXXtqV
pmPyP6YZ6hT/640kiw41x3qH/pWKuWD5r+QOjBogwF/fT9MH+kCgv5Xiwe8tGM9W
iIzkCsQMbDYADQpQY3aB8BLnKfP/QhbT3aPWqs01do3sjcyq5F5UBRetqP6Y3YUL
SazvT01690MgCwy8QAPltoV/OcfqhXSgUQvX2zPUlz1NaAOhDnZVNFYVk19a38pO
5k5HutbRAYCSJkbNwFPpMBJ5ws4Ljipd4PPUXVdoin7bU8ARpqE0W1NgjNjgLbiQ
mUKO6UqCr3xcAaoH+vypQoBB35vAw9IGTjfAWRx1BaWTEDZ1fWXlNd/KoblgUM9r
frEnyOQ0irshG/UjKW/FPS6RyDVQWQLmp+m41GSZPeSMllPOuJUONEE29ryX3edA
CNufEeEabxbgoq0Pw6dEv5B/v+iEykUfqJ++Ps2TkVQ5FpuaV+RRqwODTsOOCCB4
wg5pj7qU9ROWS+qZY1rdhWoAxn7o7wY4FL8pa5D3PmTbeLRuEbJXR5TXyI+DWyQU
iF/WUWB0my0rMAj3FQI22aIaLnkskX++DLYDpxBTOvV0inWkqTJLJLjDU6UVl0Fe
tdfH9/BhWMc/IO2KhyhAtY2wK32/QI1a9tDEkm7gnNp5NgtAUgwbD6VCHwQOMZbq
lkJY7EjfhVuN69Oy5jNcsnd+j5+xMS4N1NglWYcWMqDScMhYwbSe2rMBX4i8iGOp
mRaiTV2UrH6HkyTsSZ17gmjdcHDm56GfXNyeSwd+P8QcqasLugdoYwwKlTc3tC/o
ilGHNT6Yd5IKUfD24DUwMWwZhSpJ5gAXif0dqzUN8qBFG2D+y1MsJJD8FN23WOXW
Ev3hac9TkRy6WZiAQ02fb29O6H9xnQwTWjfnWS6T0lqae+ynIynJ+uMwjbrhAt2N
j9WSKGZoUBXUIzcQPzuzAZLNcczNzGe7jJ4MPelglMY8byhk7XGpgElSjMz2nw8v
QtQP1k1cEghVZaboqP7FpahNdnhLR6LIGyDB5IJqPTgTVSGisgX64Pt+LY0V/lSe
aVYyTI2AbN+ZI3OURumG0dMiyPeS2KKc0FhOdDfyrskWgnAalRecbPp7TJQmqz3h
90I6AkMVxKcIniJGxqFDWttic/qS1a28uYIrKqjJu0Vij1IBtrjCtqvdVTcY9eXw
HD/fE4R+fRuOK0yLfesebQu3KJJS+IN7jWQ1eFYZbLpdsWcc2h7Qj/rMq4OieuwJ
wIKnmlix/O/KriJYAw/QdhxmoE2B4apcJ6We20Xkx+dtP/sEws+Kudoh8NVS8/R2
1eLnqv9bE0WydX6izMhjmEfoB7+3fXESzpbdsa4o944aLXOxWhCuVpQQYx943ehp
1zUXSWgZyGJV4KF0TGbFSNvYwCB5xFxLUpqg08/AKP7fUCfTkEyCJbppMLgyfpKb
y8FcFHTbB8rAomiabCzHygtcE2jAcM+iDNAwEpgBxEXP06BCvl/i9TqSSi3S5sqa
PoD75a4kdlFVe9XXB9GWRLfW36ncdTXMXu4r46Q/HQ13+sRK/eD8MUszM+HKmF11
Sz6V8oQARqxWMu2fTbZfp/DZykE8HqolwlLhBCkLjGMTJoyknh0BoQm1vBsFu5CG
b3QE2nejL4HSgxpmVVyFbTLT57rYpdZk+UrHL036KV5X5smlxBY4XQMpEsiFleeJ
U17lDPocuJ68qz4Cx6PStStfIcEsVcdoJtucsLX46X4/o5Qx9wVssYPgBfoI9o3k
4qQE4pISwsv7o6+QBJOdQ1nLAW5zhKPWUwQH7noeyWJtC0qmRB2zmImaHwM47q81
9W0cIMNjdb9ftYoIrAc2lvkQEwj6Oe6jmDPAgARo0KzuTPie6vz63aH1XhT0l21K
kdd22hB5jcOznHH0O0Bh/BHs16eN7KPYjIH+YaN0YvzDkZnh606Pq/FVJgfqoG/i
MaDA4olB5PoHS7Po2zUOmZKj5poDnTQAgGCdzjuaASK1gp2ss6u3Q36J5jRulI6b
yYTxSZLUjcOzvw6vTIP7jCPgH6qMnU8yQnKO/FDEj0L/JenGejthYOlGw7hsI71f
4pl3wMd3zFXhI5PRSnFyU+9QFbcbG11SJfFY7YdCncpLicSEfbpywdix+0GdOROZ
h91k97DXY8PeHBSk03ro0Y1JKxuB1umzxrwAc3Ag/Dv+ie4Y5lr2RVCEFqwRuGgn
by4SsOUzU2OZCb+r/oEhjXiznYoCBTHdfs0pk3aA2fu8v0Ysu97VaPQ1C7bSoA2g
F0ONx/tLll12C0mgCRv96qQldDEM7F6YCcfnInXqketa92QRvcw9rALfODP72BmD
tdr4/bUS0dPuS9vn8VkBH7bcqmYcmxvNiDG0TmWUIXsQLmJiB0MRSyDMJIiZu8hv
CA6lxbZUKvyjnUSGijKrJHxhTH+prY/4V8O703ga4Offeu6fp7ta9uXzVh1AeCRw
4vNm0QoXEMiNGQjQO+vzPusGaemxxzqh7xOisqE12mno5ERgViQZTHV6l/oJFEbR
2V1RweT8bY8QhTJwxvMJOUWylYpjE5roA7Tn5t54p+nTUvXhGmv+NQfQKLpN8MVs
jP3b6+ORPGXYeB37XkyFQmhApyBOIkULOFzMC1i3HLdCClQFqrALmJeszqlLa5BG
a8kIfAEMJTsSueZdtbTiIgdvn+O0X7XgYzBD8BNl8SB4tMpGuGai1d+i8M0nVcNb
V1IZbpmuezgA0pjAz5NcNVdxw5/hOVf2QaoK+OIuQ0R8tQqCTkSyAXdewrm7iFps
WrMDcgXqwLuujB9dtFiAusMgmdyC9KA1nqB56ZKKfYaaASruah45dgMrhRAs9VmI
/BLomyKL0xd8e0anTSKf4O0kHVfJy/p4tXMd4eHrr4Qgcy49mG0cZP9p/82fEsFq
3C9Yn13nOihEaCOv1oqOZZ5K/KJl/VKCv6ggV8C/GkyYygy9mqqeBLY3Q1sWZW0Y
zz4SJNJ2aTFYVNJy3rQc6+ktRYSpQLS/kb7dqhVuvLStzAoTVr0FKjQMNfEYfBdJ
NtYTrcFCPqvd5hxIIUa0eOAR1GCNCK1pUuhN/cfgyG0OyF9RWQObYo3N2nQJiYfq
gBTaBqVyc1hcG2ckXi7x3bryppwuE+Z8Lb7cA20JhIGEXvLVa32kJsQ+6Ew7Ff9a
IyNajK4km4C3YISmPclklGd++hshg0M2z8lz3QgRh7kqC9LRvqvSNEbJYRJVENYw
+a2XWSq3MdnrpKDqFzb3oiK9NseejzBNySd6DMcp4Fhh0s+ntkUhjbNwh0IX8ryo
fWf19Zbsw56DKs+mmcCLRLrMfqMY66paKlySHzfdVMd2rnhVb7BGKPeVlAZvUIDS
JiWjQ+5NTwktXQKXktmPVALfAQrRQLuJWFYfRXAab7Jgc37cDoSbwybEFYDN4+XB
x+4KWs6+tA0xvv8p0w3vEIKxVl6atVpG1/dCgDe5hLUqWXMkicObUfwb7jit5cVw
tNtaIHNS32v8e5mWF2UBlQysmRpIa0jAFobiNgeyouPLNz804GIpXOsl9KIN+u4S
EMSNdlKGne/lmWnzhd21ayrqqjPTvSYBhBj3eT2i68gFAYKstAX2S/pzGu4UY8X/
6b2P8T64eFHZsmfPdux7hLcCAHq9NqrJxGMTt9AgqAeF5EPcmXYHcoXfEl9WXbNg
26PL7WAK8RfgnXD8phLjjWKze7Eg2NCrzi4W5kXHGRUbb4fHpiEP4liugkFqJpAT
3T35dSoeS8eT3njr1z29nS1pLbNsgwBRFkpC/7zD9LRkNbxO3A5tinSdGhQ80Vu5
DHhwevjyhKAu5F0NiqRyf2Vn1+pwAkB+hAH/ChBv5E2zITiGSV4TnLdW4kczIBFT
011PkeNaVZClQxn1A8D5CcwEnNCETj3ihop+KG38raOyqMrgLopxY1KKEizFhJ2T
KQfenbbWdEuFOFKmoSfup8sr8AiSZceKjkvTq/e/MotUrnYw3/uVJgX2Mo6o+u8f
vlqUdxZlWSeRpaakMJ2/qNbpWl2ZA4M8GyPz7fNcLQzM4/4cqN20SqfpEx2qJJRL
qpFveSZoxCUbya9O69PVZNMDvatr+rCAP9xyqzRUAb6mEMh3bqT76qpuUVXUlGdv
092rIh/SS7K22cPofxzPmMb/yJxDDKOgjY7oqKa4YM2xoYJjnAz7kc+2d/sDMNyL
jiUxkwnA0YO+aB4nwSgnALKiPYlk6Y8+jBflGZCl6HVDfXPNCzuw1ZMbul74kPnO
CFl2/qG4+ypLMCd8394PUv8nrPQwEWe8T1ktDyUsngH9omBbLDJoaGOqpmHjcQGj
3/ZYrIHWNnFX8XhcCg11WodMb2OdvdrGyYGeyVRT5/zkQsCFcL4GE3aNajQZaVFr
C6NBtWzKBF545DSC6w+RL8MY+3MD9cJtAJvCvOqkgaJ5ljvkoADxR4ybeCanfAt3
sJby3Imz22HZLtwK1eA7zW5wbH4qO+t+o2C4KVhG9JSkB2D6S4riEQpkPLmOXcZj
q1qx3WPY2PZtDYd5DeBt28EhhPuCxD+u8a8aWXKCQuOXU93JIpL4zibzjmtyxORt
xga/Z5TwOwlR6+qnYdKM9qPOq2IQp/Cb5iald9VrG+SBT2eTFJFhcOQjilYZ1eTa
R5KoyUP3/sTx6N4S2W8bqIdn94L+D+w+P05RoZe+zJLJ+dIGhvMmMBbKQrLL6akg
HMLJ8ibe7BJgeQT2dQ+DzlnP4tjuwoaf6KnSaI+QvBdKvq5vPm3V0ZTpnWzL+KkT
dVowOdnd4nCkGR0jWBeid9Wev+Am6uFHBPFB5+/RjtqzxSlaoT/iosN/0FxGDj4u
I1vsLPjkx2HiksjpMbSMOXi226s0MIH9JM+K1TM1WzcpklBblSx85Ah3y5JtjMGa
/nMrdJXawKJQbuzGcRkNwqx8ohboTwq/h938ppOtoJJD7q06xFU949FEtkjmtRzw
gwjjwlahNjtuBqj2ZWc/Xpizs8vtfWJciPLsoRa54bjURAIZjlLYwOBOibmIe+xH
EFLP0EKUoVyJFiczVXgrRRREws53B8o18Cu8+90LUYAp9InUdE/XL/xPPFfC5INx
K7jX90Grk8y/V2Ir2jHHqjAKBjU/lm5t5TM+s9by/QdVa5QMAEQt8bdyjr/mz0Vz
VJK+6iNFn695BwXJGY4px4WS94pKqGGu5mTxj6IKEv4OGfVfZSqL0/EKcf3NvD/s
lEJ50C4U80meyLZ4QlqJo7XZGvxjsluysG9F9og81c8h1XYoDvyDdHXUG2jDwVZx
diFCyql64n3JUIwbCegdb5wVjaigtBFEXSJ0m/i1flWQtL0SEHdlMbuEh2ZwuGNh
Csma7KjZ6p7c3O4YgfQ3J4XBMf+Hplb+rcWVDZuT1IqODO2eh6wk42YPmVrOEQnE
huu+dRvUl+wbqTtS1zwWmS+zQP9oNUZhi3qzLsQG40/j+4f16nNmtG4P3PJFaJvd
8wTDMEFbmQosaI0z8mck6ISCwuNsojgRQCGpYXwXkDfXmvBzjpkGMMHz60IJQNvL
/zRVao+/i3/25lTxkSgZiaOG2nl9Ii3Wj4750Wq594Rqdlirbi+B4Oq8pJqIU2y5
mZT8wjOfUrUbp/ojpm5gXluF/6MAOW7T2BLfKIn2MCJgdJzvZT96g8R8K2GwX18L
49w2PFlqkIM6uwUeo6UoNNpz2cYesZS7wltDmwH9cjJrlhaITL4KcjPxldiuwAX4
de7kppj9KXkEy5Q55Bp2bWYKd4gokzyVtgVOAUjCemNpg3ESxdMGsRjLYt4E/sZx
/sWqp+JpyEiZ3yINniWG68PZtuMXkLXsAoCT7a0ZgqlZSbI/JPPCiV8B2gP9zeOD
2e5WRw/p564uDc+n6DKjQc3+c9PSRwta3Tm1VcaYmsnaLB5FyjKFdRVfthZGBVHi
lGLwpODrTw7m4JWNtHSWd3VvUESMnl2lFRqW5T2+OnNbAXJGu5cwobOMFpfnNBIw
7QAX5h7KyOIQ5C/vdASFgSOZ5Bc56jpcZsr945o06aQD0+beilR38Ax5KS0Di2lO
uQsLaUQsoghu5WFRkvB5nvKAD2TCki6VzZ7BGG2eCnoiuWCEnKyocIvmkl0wQuDC
4gM5y9O1XrP3s3w5nO75rQcBzywfjpaxO5ThcfX8Ovnpu5w1rhS9i6JAxIdRzWh1
btG0quvXhnPm6re/pJSb5yvfNfv/9KuwxMF/Px4i2EpCtj5Lte0fCnrgYEgUmHZj
OR9BsrA0kb7NhvEjjP2FuCP17n5DrHaGNP/L8C13SrBkGxGFak6fznSmU45Dr51e
iVG3rMFRjDchRWfFfB9Y/SHKf80i0GJwA+WX/tTbYyB2BUmAG2MMWMRsN3rk9TZ+
9WCbaO663LO+lj4O/dE/W/jqId6uwI9REgYwNPK+10OnmmXRMAifseCQDu0ITk+M
Ub8RMO4LuhZ5OBse5eYDv7XNPss4oYeeHL4Fx+IGTpUUtRkUKpLv+xNlaf7Ze01J
5eQHp1zWLmnSZjptk+f8epN20A3QmSw4AmAvlVDSUUKDewO4/dC3xpH01kMqcDG5
4neJOY/lpqMadVZ5/FGLBOaUasyAFoO5iJINxJd2UNIylvlSjN7FYXP9l9Av3iDt
A5HwnCWkZ7e0woRgVrSTGaGJy0AXdYhYhS+qWoXMIwJhMkZ5Cmtq60XInPC+LETA
4aFJOmVvc4p1q1XuqKOkivsVJY8gjwZmz8HSLmy5UPWoVCB9GXCwKn4q3CABAzzb
pQcSZPOqOrlh/79aBEJHzfKsfyyN9Q3+Py8Sd9BpfvTExhUQ3ShZxM77S3X5kFIw
WWTKr5j33r6G9nAIQNMwXuDlk4EK6MroSgPaSnzYUZZApoOosdsY7EbVyYMQl7/E
iX1c3ZPWHI24WA+bFCNdWaY6x1N7JPq5tBfm4E43WckCfheMDHJFwBnGg3cqd/tX
HjDS7TgLBq6ayUhUYajTeFCx/mwkGQJ1+w/4J+lk3ngS/TTkEVnmZhOiphNsShVK
qWfWf/LupwcX6yO9BqALwt5idrB1JiVJaXdnsvPo4qCU2zx+/DO3/WB4/66eEXSq
uLN7GOZT1EbtpoclIqq3vC/QY1kUqjl/31cq8qQjVVvDHeKvwhdhWTxya0KKoLP4
gH4mBAs6Bk9G/zlwvuqtJevosLum3KPL11UKDwBdQNh6duk+MNk6gSexu0fMtD28
bCwA6UEC7JYChWxpM+f5XX8N00LrW6v0NfQq9DUKCeWNFtz4IgfZDeUD3wO056nr
Co97/4W9xo1X/fpozkQR0tjvFslyQTltolfkeGLBVmHei5GqjuGyOtAJWNkMQpD2
mVWaKK1LqtstoUI6KRBzyteY///0gwvJz3rSixa31TBILfOJvrMklkwk/kh9meie
NZPoaHZry5vyu2d4P09YGb+AxKb2wzE/ghBAUwjlsskM9SChbqKVJI/UtBN+3okV
XPUzqTw238bN2Eh6/r/FXUssbpu/vAlahVKQD/hya4zz7Av0J3EK6+zhX7ybHy0Y
5E2ynpMlRtvTQGk0++EdGpu67chAxxIN7swcW8HDPoU6/h5F0ZRZs2oqKCodYeGC
4JIfdGRGoMoZNG8Oavwk0VeX3mS6CJvifHqYHO95oUHRJp3Cu+W+IPhVTs0j9IuJ
s7IOddYhuN+UMLgPsf8EY2JpNF7CnaYQoJOliHVnbkh4njZwvUSPjgalHTLLTWS3
8ouCI+eU4cCWw8fRytQPetYhovFyR3zVVrshbCh2GQenZu6PmeMIOirZHDvMuR1N
aHuFlrw0IwPE/hlqJTSp/Q5Z4o5ThjP9/YNsqjPd0C1tFUAX4tr1EVDizXM6ak0D
20Fqan57e9xfIMiqBn0QBUQ18TOAtObgiE8jtzX881K78//g3iisSZ0C3yR+bDHe
jOEVq/HvCGy2SOWJi/OR5f2kBi2CjnpVUPnWva7XRtS5iBcTvF/GNchS+CTBD5Xx
7mn6p/XaUqILXGfqpbrMHU0PebOBtUYraYOTo0ANKxmwF5xMAvuqv3CtUWqzKpmw
M7EIAmgXDlBuY/VEVUo0PpvdWOIAAHPzYNhkLjP/ZSLLTA3vg8IPsSmCi+KqdENz
2itocv0vlW/EvddmUV2V+wJZtJ55e8fuSAedJAgbBG2yylkrNTdzC27UhfG4mqBQ
S7RW/VbVyOMuoq+LTwgyZhBSf5gqDPDt+yLaZc4WfxH82LM8EGMYhtkTOtJC/B0U
XoIBXJgdSSMasE7v9m+4LAEAtZYb6JpJSxFC7fKNzM8W/9OxNjFITQ3A7joi5pYl
y1cwrmerRqgd8fzn9W+karJMT1YQSGgIbmMrWO8ZtJHMbSRQ6LSvZp/FRg2tSr4A
16/oWNLOB5tsaGdfcltP/IeIKeBdcuaXTcKiYGK4VzQCtlyZg2+79u0gsYHk2BLq
wMmh8xh9li9nq76RdzQWmznbUszRgRbirnitGP4mJ5tKpjoLJVt2WpXhozRNRQaI
u+RDz8DWe5p/xEUq5zb7DireGynTbNm1qitiMHJdmIjz8xtgkGLZ7UybBxmzzBTL
wwRi8wkBQVCAeJvHVMRdPsqHqEfG08nHZYItr5vfmG9eNcVBTxa8ynm3X4EI5lSr
96lv++w/JuIobj+4hr1KzSX7QAtjkfdENezNFhc1Sciv3ZgqTNsRokTEAb7N6Rvi
q4rkEVXC0vx5E3adJNrFhgp9xQ93D/kvy2oOlucDM9SDVywIm8PKb2yzy8SwIzl1
hfoIbYoEzsJgfp97t0X6RdEZF/gz03ZPIE5uovGlHp+RuM01FLte0mbx15SuQEl2
XRyY3l9ezrnP/eeNz6oDqnjidOauni6aJ9WNZmIeCMr0a91tpD2QWM23W4CG8TTE
sOkjhdt1VMNUf3P0w91b9tX+F5OFE6o0FqZmt0PheQTx4MZ9wyLF3T5j7M4LiQnH
aEj5YU4Y0rJ9ZJROi3lbwfqflLyqAGyTtXP7R2KDCYWkE1DmvjYalBi+Lj9IxN3r
NGAi3B0Rol8SaKnxt4VaHQtXZmutKXhCOj19n9ehDZLwQOWbEzFDNnCBr8q9+lLP
qoJtFKUbF+h4RCSPIQQ5L/Ks4EiLUsdvjlB6hyPYw1NPDO2A7QVxo+MWnkgkqe9y
S8hqjRbgksDuJneu3zpKvLmtuW1SxxupfyJzWNx1/1+xfQqeFIalgxB9uvUJcwiJ
l5WGe9llnD01GfxxKWU8dajmMOosExmyasSuBO9GryPph4X+GEk+BfLpX7P/vAMA
tCbS0ImPn0Je61uuJWbKcg/xB1SIjOaqxINg5CAT4F5cGHJY8rskYPyGw66bE3Nl
/cDGBYB1ge8AUBAKGJtza+ylIxkJAY/phuaH8HW3F1KUWxSYGHHayBE1kwWGzaSD
qjgBg8kS7qesRcWw8xGLKBC8pCIYTlcy3qzPfhLuKBsV8epVeaWp/WjdOaDWNMWf
PVySvDFDKNih+9KIOk2XQayP3APC0EUeTVPbEkFoUW9Sp2Ic8ykl41VW/WDvwxSU
xdbAa0vf5PEvSirCtWzW2CzKRyCVtjMXjwS9NYxSYV0KgG8rH1/qj0Dj5yECUSbR
XxaLWJ612xwO7nwf3j4MHSkRHFUe5iCC7/g0/Y/EdLS6Vuc0uBPcZ3PC1Xj79i+c
L3bAA7PUGKBWCwMy8NhCHEI1o6x2w+m6UPr8LQMjvnwIWKtOD/u6+uYGJWWXV6ze
cGP+UdDUNvFHuzpGcjLSwcy8k7/hYWZxEY0jOI41jSdoLF4Hr0RRb1VHVozil9gp
h9/dwPrep2W14ccNYsxmzdnasvHC9ZT80IhWtnhGWzc6KSzvocDsGGv41neMn9FS
oxToaYECb8yZHkA48eNKGeXsnoEuMWKXpQftQiu9G5qMcGrhdar1WUcJxG8MFfqy
R8Gr1+DZo3mrqw13oyIQU50mX6RDy/uuR4YuYbVr2CZX27GOdZ8Oqp2oEW+6hEv8
/DLINGcmt0iMze0G/uKdzbWg5lwibNuCge8z8hXo4ojPNCIbRNLlGidx4zZuulJb
luIKMAnY+7k0Xkxw+kOuSuqYwMTbVbHogXpm8X89Ps9udNklEiigmXUuOphI1WMj
5dMFwi00Omyt/6FA1shkABjiPR2RFU1lB9E3KvnfOFV9F6BwITeiE/K4pNbgUOnB
OSp8ncvcFhTa/7zt0DIllFtXSoVLE0F7uLRw2V+d0JDkeJse6YTelnIyH1LBVP7z
TugCDy5ybeiuu4JZtkP2NQfq+Pi1wGifJlXAECdHs8H7poT6R/HKT+1YAlge6j11
IjviQsa5wy/x4GVkWq2ColXBB9Xlc3y5qslMX5s1NhgoiSKh0mZqYVbGUxK0QB3h
I6eub8/vmM+36yEmNP6zU6MOOpfbyVeqruYOhifiU+yg3aMUcqK8zpUOgZHWMHf9
fxBn/6al0In30h9s+qBY/OqIhafcZUtUT3zAf8MHIwApNCzrNGcXV14H+76xMyVd
x28EVKIJxodNHL2goWwtblIlmkEftETG8R7RWlkTKw6560OLLY91ZjioOeJ9HHDm
JRYaeE1WDQcdwuiAu0mtPgKYUtI67yLFKwBsfQodU4YNRAU7xzUv/sgfIG7O5eT7
7XYERSsnJQoi8SFaby+VqOcSdJRo66XsUTdgjKytpPCmZGGY/QjkqOPQ33P8H8Gc
yxmRe3XAdvCdQpS9aomd2ygkkPBnC+NvjPnZpvRpoS2aDE8JG4kXDuahBFGonSVO
19kgTout2EsJFZNHKdWTDqERclVDhuUyhwPWXMFkxhoD2eh0IKstQZT/bGkSk2PX
va9M9iXVGnhjIceMuLYJfyrKQZl5ya/sCPiJABkI+KmnU76Gb3Iybj6H2UMYum/w
kU54NeboucRqEm1fEjUn6KPjcuQCNU8hPbDqcZ+WU3eB3oM37ZHzFN2uKfuigG3N
KserO/cDFgCw9GE203oSDONBYEFVYhTcfojz4iI0xLZSg36KDMZsn8bbPYrdAd1f
VmoZukr153Befd6YXZs8fx2OBwZJ4a9HcU7Oj92x7JougXIkv8sf36Eq0J0ezxbX
yOogm/viHIx4BIzSFvKfaxiZw931/uhW8KOkv18UeLhS0l9dAVp7nqWq98majVp8
IKO4rBEw5giuBGXiKbvcUY3lMbFSx0m1Dq7DPr0a0cuGyeGDH4USL2G07BUDq2Ai
NLr9pJ2qJ+9SI4AI8TB6FMHrOp9F5aJYWP6KtTY/InhRdQ7jCMQlVsDwIW86qxWC
TIGcbim+7azKeKM4ipNYfhd9Rdf9wbMBkAHuX0YkoKFM5Cso3IHaLRJj28Y+Ha30
xGU4EPYUpFcJC8MU4Fr5LiSq2P3XaQYhbHIRnjdrlrSv/yNXE5pMojf5ckO5+wqt
KQjwXGVAqgW9sebj7SBuLbMTEgTJFhpZNyFIYNMZvPdWX06Qz6cQVe7s9g+ULJsm
fHk5Gt0nhbbgbUhyPj2nR4asm5SLW9j/tSIs4wlk0H7fBv3v9ZCX2TEjFeYIzqqG
YsH9IUiu82EVIob+uOIXqOLRa0cHZYzsiMJcdNiqxy5RnKISYhSmta1Bz8p+Jo20
Au9VmgTwFEoYPESyJHXjudLeEdyWcmDgSdnmg4oPTpEZpbznHL+rMR59P27ypU90
lRx612hncF7otqKzSbBLGuE2u3Zsw7GQnAUCMs4J/OEdeGMkZynLBiotpYkoaek4
J9YTcOqzXWYg5JQvANPxf1eqCiItws9Pi8A4iNN1TkUQNMDi9qXM0t/1qD7u5Eeg
6xx4EvWMYnw4jxwJjrac3d5pwwTj14XT5sRA5QC7iOi1gmJRujDeN+DBW27Swwd4
JMnTDJZJgy6QhUBjZOGYxcLxh472cb/o3UITjHmR+4r3EfH2FhPr5wZMxBG270TJ
SOB1blworDSmANAP8m3Mr1DE38Y8ujlecrExC0BhDe9ejZROo588KB4G08fJKOrr
J7VULTa00OpJV06lZLtNJxkqDQ+l26jVRsZSLFQFxmql1kJPs2cLb6ZqZkvlbO+L
rlzvEMmLl5c332u/qdbIs8x2Dnc3EeBl5P9KudT0wbOn+nhZo3jYDmmA7CAEv6yu
ZtM/38s2KUrJrxtfMdg7WVKHDcCfqTlFXXdeO2g9sF4id86Mk5fe25PV6b81+HIR
rsD2NTVd1mpkaBU9nQ0/f3Nw8z0CMFtcQQn90bSQ6glnvZCKOHpnXBoxEo2Ol2jU
NkcFd1TmGDB8MpvfT1emReNlGFlyng2lVjMxJuekZbLuzOO1AQxK5w1akylqIeFV
Xz2m0OYO4YXh1nyHSeVuopbzRQktPDYAoo6skZAMbUSzK6OwkqUEG3jqUEMPs14y
n7B/Jt1EhU2conWsqdVei5Ha9iBWKvb9olNwD5FMJmIPpZRAvgGrsyH1KT/H7eMD
Rg1FK7My4U4sjCWjsPVwQX9q2AiOWCI4opk+UcbXSgTPfp+Bqh5kqMX3fkNLJDUx
8cXfrbW2bBR1YeZvi8dYF1igrvYK0ROGM7kU1IVLB6CIWF/QQelMUyge13CdPN2K
HaOHbex8DfFYJLzxhnfc9aDXYY2QmRcVGwRShrLCc6dz5/zOaJLKZMH6SQrLiBH7
geaiAZKsznJVPyMXkGl+Iec35fq6CR/pHMDo+6LIMYRum1OCVgf5l0Vzmm/rG7UT
d8ixVHC/D6djnT2lZBKMWZk0QU4hmeSgqeC4+LgKtXEiWbB0BtjQfPWyI29o5c9m
EtFC0oVa5LRoM4n4cGhvp6fjco23nGNCrIykqNtI4ZpVjk/1z6o56RtOqCTn/NhI
uSlnQyu89Mf/Z9NUcx3Ak/MrIwIjsgka+bUi/uLNHCRvLRWYYg1Ef+qyeagN5QRc
80TJDrtwu44fMY4YASQqyjAjlPP7F8TI56fTvsskn+Fw049SZ/gvvhErGU8uyuTP
/s/yTq1MvM0tG5Hqo0XjGP71Gvffgt8DkSxSQVOrkIONOG4uZgq6mtO1Pq7jmb1j
kTf1zJ3TO8J+qf/C7ebperOFMc/G2ss1f0wfB/aqspu7Z5nYvvFCvTrdlLuR2ipF
/ZhzDAUG1WISSs2vLH/Q4ObBC5z7Vb7OVhA7lMScpYv4MUCtxeCIKjJhQ5OL//eJ
V6jkSDV6+mFi06Uu23nsf+KhjKCDHE1duIT76qcYALQFtyKL/08ZCZBHKvgNLFlS
3v5nQZAu3Xn/hQwnHGEUPAiGbap307Oye2qVjb9UvBW8+RR96SJxnA1DDpOPV/Hw
58tRxVajJy/ZW+cxBN1f0R0AYwWAZKQbH2AnOteD2TG4jT+WgEl3SgLeJd7/69af
Z7SF7/MRzzq9SCcl7m9srxSct8NkQL2INNjvb01BS2XVJeWJP51nsNFBK8Vx9hho
kfm+RJkabZGTAbCW977N4yXmdkT1DndYp9pa57SvPfQykl8mvnMppx9VtYlfQqZX
REYSNRvZIeoVE/f0AN4YXIkPNtbWfY7tIw56EmiQy/u6Lid7NvfDDfAu4tTSk+cK
X5JGg+aHkwRW0e5V+6kVUVTYXlOV5FoupbEthx73sHy1IkC0BeDHxBPP3G1NkB19
wFZEYwfOnso0U0ifHn00Rk7HYH27U+0kcMyDnLYhxCbs42MoxDCC2bauDo7TwjC5
FPbd3u+PNlWXQlL84Q3E6OngfgCUwBJpJeKid5LbKPoDd0a9NfAhuKHX3ReaOuaq
RnouVgFBwjGzj8gJX12wGDjTb0FSHeVoAvBQuEZolFNLhyBcDGon3v9eBQbWg1y1
ijnoFiLlhdr292JI9y4sT5WrbfntmF5wKUFIJCDPQdqdPx095Ho2v3Z2NNSF+t7E
F+Wwff48fdjy+jA3Sy2PH/a3wKF6U4gXyd1FiMSjII8E1aqtaNav9ubTjbsIPGQt
B7eejm1mIvBHO8ZJUJNhlwdOpz3fJ8R1NkfNHse5v/73iBhDCWXqT0zdoBbYFGPJ
g7Mc8IcpTj6JoT5ughglt6gACjAVJQbb+9s4datIExCGVB3Il3f/+8vBs/oZOTbp
5U9AxcQWFt2oFjFwAE2XxPk1jL5lh9Vq1P0bc1CEsNnJXb1JgDsFOzg0viGQ6ilw
XWpo/qvvRCvD/OOIMZI2vaBttZq8HemaG3zCpfFcWncNHJWdVt3t4S26/rzGPjTr
itljDPz6Fiz3Ulr22XvkbM/IpFeewBPLVPFhiMs1ug9EREoqlOdcoEXDFcm2aBb/
JSssn/OcNMuR9B9Xg9RHZ4ZoX0x3HQL5EqcpdNzp360iCJIlFjSKbGzDAmpouLUm
r+jTErNzg6IND8aOMLTZgbk2RwfrM88NIg0HTgPg/pydjrrXoXfM1LsMXDWulNB/
Of0LtY8SFF4PEIGt9/NEqqFq7HKss4jVrbouh4ry7TSy8JWD8AF8WhQ/5AtOa3xR
vcsV1NuKq0FmScyiILBAvpes01oq7smDOuLLRbKmVXVadJP4atl855fgbfnpFLnK
ocg7hhKD7d0ow/PZDfvCNpGE3S/6glRsBU6yIk5epVtKyLs9XaqoZF9KkM3vE5zo
nInvjhPhY+SERtrEnU5jvbI3m+9JpTMcRXKCy1nIi8u/3FaeBossjWnXHYsWwOFf
QQZpy8uGShakjd3C0HEs3ju2hIJGruquXe1+anBEMHmK0awvXfsT28HUykMQoR62
zfywiKlKgc3Anq87e1Srux3QAaLqtsJ+IbZrkfgaoo1MrAhV6Tx5bom7O6ubF5c6
gRaMCjlf7Jz7wv9veV3o/i0q0JamtTB/i8N7v0jR2wfgc5oCwkf4vi2cC3qmQHIX
RLJ68zBl2uLE9n+1phk4LQro25+v9bsubSMb3f9irFIk0iTOgrPq5gdDhrsL9NjF
TLyIr1BNnEM/hoP8GEBJqWDym6dHK8104wdf1K3SnRkiKcFd5vyy2n+vmXfxxeMr
0bTlMmCYuywYzGeywtgTW6fhMLPOxhBJGEqfvz/j/KMCS4PCXwOa8JQfslK25pEl
AUrYvgNIPdAJpjVVNAYJOdB6n3qGytqdhFmr4hG/xDRRVXe/xHSy69J7othR8Veo
wZSCzeTZglvIXYmWCm7SOeqMo5GnURL55O0u6xMyc3w8vNy/E+DMuOgOxnHO46DD
ubMELmJrl2Ek53r+QGJVexLPicwNYEjtIF2TDSVagSHjtWfnFmiAeq9Cdw0byq/8
NAaJN9Dqxn8sTS4qn7e28R2dBgPzu92yD6scg2jmRcoeuRqEwCuqz6aAIafxOes/
o5fnCUIPq9hA5BDuUDRVWHC+/5ZHW3KFo4pk10mwq2ylD83dBGAR9SgAPxUyPyXG
31/iyl6wNHoiGodtaSM73FfNLvFNn1T6HkXasK2FYw1FeMFEnJqGAXtPisXTZing
vkV3O9Ik/IehlRAHraiJPpJNpc28OkboISysaEd7hyEiubEhgIxw4uV+sxpR9Tad
WjcCALCMhUjaXzU3EWkVusPSNuai02RrZckir6L6c+B+bc06OvMnsbbT6WX2sc7e
9yaWFkDvz/5EVWejOapBtsmfsUB6mJtgFqB5vj5BR4sLGFttvbi5IeAbsgLazKZ8
wjsVp2j2uOScTLZKY+LyrFZToJRXIYZjPLsoSGrcSyleEwK7lgOVq3e84ZLVahLR
mvfqG5AyxLXj9tgwUmbgWIyH2zma9ZZchiAH4qEmS6KKGcA+G9EqmBazzXCpsTNc
jFB+pjOUcz+9Rfgc5qn+OSResw3euVAmBzPW/D0S/ll27pxKHgvKi9X58lEhlyG/
zmveRtqG3OPGnUKssQHpCDvJtryojHstVu0ynpodP1cgctJXlzeMWt2sSZBblGkJ
KsUaacWXhiOh2U79/TSL4EgKnG1Lo/otYrPn440i3uVy6gUEYUXQsUNd5npomDmp
SVhmdDYxwO1jBVmzdLrOJnpifD7sIzjlIAOt0QS3iW/K3VKKDJ0RcUr+5b5pA5t5
WDCjn4ITwD4AuLfcEMi12LOzKCZnhEThEoeqQqF1U7RleUWULV3CZuRA8kjIEWgQ
M3kMsG8K5A9N5QqB12tljEXgUR3r34gHAAyvTaDvJDUWr8jW/o5TrsKIH3bx6ojU
2+alIC2hkKDfUCXQqDUBB9BX4qfKBNC8nThJny0wEte/q2n9jTcsQ6fsXjqJODP6
lu8wZieNQZzcPQ6RcgMr1K19WuDIAxlbUF9LUphE9vd5rjrVBWoOPvsIZ2bPo1xG
FTpvqHRcPXekMGFvrE+0y/6Vhcf52IfTkZCOAtrdr41Lvqf+w5/cfSB1U5Yr/o/M
A3mj5s5V72Zq/8F7fzogKwFmuptuiq5/iRKV4gETlVXRk50+hDSbiuK1L6hlR4bR
IHl/KwUs6iAlUzqJ0w/YzJyCyajo1aESFu8z80bTrLZGsJJzHWrQR8be6LeZ2tz4
OWxV0RaCk8n28NZ9RjBZ+GOOM6TlTUidQaBqk4a7Q4p6SL991wOh7jTZsNxRiqb7
ZZeJ5Em9EpOyQmje66LUQnjBn7MHGZ/vHLUEpAxbuTy9VBrzr5qv7KWv7HMzgz5W
wIoW5mIdGClC0Kpted16kgElue7oi6/li6hgYsDpZ75KWlcxbufFiMi4tyG63N14
zehITEoiYiSXdITd3PkP9mBEoUgjuAWU/3uy1YX/wO4whLtWXaABK9Nru91UldXx
O7d5Yv3sua8Tyirm3IuM8G/ppaO1cASX3F1AnMsq+PKAoobaKETyO9ckyE80ywiD
TwebQ8YIGFjLRFH/ach0aibnIgLVo6QqSWSmITi199usZIozCrZ77AMwujhX2QW+
G2QlsFrG/WSleIrHPsPrvbZ3s3VkAoGH7OM+Y5i/CtwBmGxK/Q/E1zW7aUd8wy2i
4sb78Y4/cJydS3wp1dTeN2tHFj1Fz4lFNNqdPFpUm9DOhCjybzIqyJ3wI9SnuoK/
SxREQfpdwUTro2oqq2bZBykv9xzXJeYe51mIz44SD4VwKwp7i2d/SpdsX2yw5SED
1bdu9Sssg6tCRDTpCsNeJdle2BsZvJeUxsgZd5YiOXgXLX60Kp++P2Ooo/SQUzie
7/1+5KXC6czKUZOO0M0IjbCvrT2QfETQ14l5XGYckkOV3GVFn4GQIXu7GbjOoMPm
5xpEXNTFZFGglpgn3n6I2sVjJsTKTgZiRXxxGXFiWsNqBE1Yf7wt9JxbmJDWD/PD
ettQ1EMg4M6h7WEZh5kV/vnZdATyHen1p7pAOB/tvnrQ5dWJI+/ZOEC1DD/Hy180
Z2mKsL5bxIIvRX8pla7BeF27w1++7fCRSGhVka3AX7clWh+526zXdq3YxAuVUzAv
lgQI0+Db/IKzElUL8ZD2V92aupD2jI7NIuXU9q2hDociv7PSkKykBLjLuqZhtKgH
Tsh6ML6rzqK3zH5+gZ1+61ZNNFQfrRt+nfqY8TFoqp6uA3Xf+UUCsD6WrjilA19m
XOtTvZ7hDlFPC8jj1aEK2vh4r6NbCR1mo590h7cFC+odhslGlsW8Y7Nb2Sx/khAQ
IBF1tUqhJPtljGwqEVowEzMyDr+v2xNELOz0z5VxzVJuUfEwFDaUjR5v2Hrn5G+P
Nh2UuYgElrIuLUl/I/glse2PtTjfVAtm/GJCBubRZ+srC2ki7NlXBguGfoFRUE79
FqGFjXrGb6hFjf04VYAfO49rTYo0wPd2Lk46XwZ0xaXfV4PUQIgNOOCkdrFuU2Pw
JObSXIUs0p1GiaOP01c+X9L+gt2W4y84ZLPly8mblDPNm/onQ6COktpVa6fQTXnZ
qFG2xnbmq1GeCPOju42N73DOAVMoEAZhRAJKIaW8LA0E3oTlBDrHrZLxlwX+IW6P
8aPQYqZNLqJP7apo2t7PIZcjquEt8HFk5psoJXq0lec9Hnjd/lp8C10L2epwfC3m
N49j3GmKcLBysNaDcS3Va0AHR1Zw5nLTshf/KwgW3HQD2f+Q8dWU5bIloFxBIJ0U
4/1FqcSGH6daB9UzO/L4tN7txtMSlnh//6Ebn1M0JsnHznh0ZtwiTYnNAMO2HraC
j/QIDvJ0tt1hQME+CUlXfAc+zRjoS+cP2rSRdQbpQALsTnz3Usm71612XiJqu6Ff
y3wcopaIKykOUZdWDnnpOq51swBo2tiRKurMU3P/NMt1OFwIbXgQQwH+KhpSap7m
AFGv0SdCcCa/tpRU6iIAGRIezCM5pc+iqLv3iy9lwIdVwpPXV5YDiyGWbedQiOoC
sJfVXMnFAQDWGpZmdFem2g7i3N4yjAEdk0V3hi7orgihyF31SDM7J7iC+3z/nX/k
S7U/HJL28R8z7ax6ROAXrFHF2ATZ02T/oSLoj4/M2EPFfo2s7kbZgexAHBRgf9pK
UgO0T9T9z3BWJntB1cMUcgIZX1RjvoXuFAFYcopZU/eDw4S3TKVDN9+om5TJGTEz
Pdwggf1YKhErfXnwzN4tD53uxDe0J2R7I7wkNZT4dMAqRafwnKPTZSHJ0T1+GQQr
KSSO85aO9Y7fHdb6Dz9ezLgu7FjPq3c9p0Jz0UHa5ojZJFN38ELxQy84Zx/TBoYJ
5oP1/qF9ynyHmriVTG8NL2gF9GzGioR2r2dlcGDbpIVYSzmfmahYySPH25iJj2iu
eXECfMqBG4ddTjk938tl5KwiCm51zytkvDb8rFL5VueaMrlCu1Ms7RqCrgu/pwTQ
iYczVOy7LrfTdMpw23Jumfg2VFTK8wBrusEJHFkCafZv9tvq6txb4oSvnfxjrLWo
EPqU+c/e9mRXop9xNmQJcJel1VBCOQ9Q9m56C/CDNoMqRplWBImuU+BgmxpEzGK7
8GGv1ussNh/o1e0RLODcMjUpFAzC1Xyk13GATdcJ4OAx7yq7z3/gmM8cO6tA85n1
bYUS2j5ecPblXTlfQZY5Bvyki9UJ1Q+tLA6bn6M4EbPt89mAQz5mw9X4naWd6tOv
TWPWpirvSXwbnG9plFjZPWnQfMkzTzFrpbQsYYyiQuKyr/SfkeDmuDZuZeXsxKI9
eY2V6h4Ev8XiKGzJN6pWDP7Ht/O6w4hdRijTBTqJo7TkB0csUNOq05kztm0Q/zA0
NbfklavVKxGiI+wgWAbJzpOTuoL2a+S0CMJhvvfbGCSw0G/CLD4/xuaPdd2r5E+2
4bQWZkoBL/i+RDxYPqWN/sH5fbBQXV0ZhpMmeJc0YnLWklCG55EX69uGWYwtKo49
XGK/CtsF0cLkJfC3fxPwqEHInpDeqA01MuzivhBPOxzDMllLEG5TvnpEI6MD45yS
ou3GdloVg18LbXyDWOwtsbmX4OwpSt7l7iK4QaxJdIvrhKfyxAQhaAruzCrIYr/i
sRAlm1yD2OijjKcTU6jHqQYB2KW2aneNUzDr95VlxLAV23Gobr4BK3dDImqykr4B
QP9XbWP04jYWPgiuh3F6bfnUIFVOrOrCPkrY4f+o6d1xA0nzvjlLiwKPGVvd2qDE
AVOKw085dy18Bl3kE0UU3qH83IXAJo5WFt2O2GxzW7GFP0lwR5fQhAVVD+DXvOAb
6yCQ/4iH6HPLpPzrTQ02pTAkD+pNgHCfZcooBa1y/o0nrqpmMrEPAMph1UAKabmM
MT7uW5lurFoDA5N8qq6PYE27CguyBQEjK8Dzt59Td83jXmKpOyv/ZCZajipj/xw5
nD6mY9IqCZdUmrSUA2Eb9utlxpCM2zb0GqRG9sFlJyKVi9QVkosB0R0FOoo+rIw8
XOv5Y0EaOohGh+8mRE/kqAMTZwhcbDJmQ7sBx3w27cfbxG0PvF6isZDgG/VsTSuW
pqDHZLgytTScOxw6Q/N3e02cl6bM/X09L/UrGLvIE3q3+Z+A4CIKgHq7XiO6L79z
WG3zDYp62HTcqhgR+l5Viel6yR8g/wqAPdVB67CzYI2de3CWXG+TrF3kN+UHWt/m
CuFcYBelgo47EEhsG9UvsKgXBNNYAMOda4EV104Jbbi6uUmpp1e+Gns5/QGdaaim
hWo8Tkxgi0xPhyTcYkz4qFkKuFjcDiNLj7fDeP2fke6TsHt2jEMxCueM/fj/gORu
00+U4owU0LI3pZYhcqYXE4PY+iMWuM+3XPAqsYwwjB54IXVJ9fPF1ThZqY19Q/pr
l76OFnvaq+liKDpon4wFn4rpbwmzmsIqGGAjWGI4FEJgfCbg9mhzS2axyBZaVWJY
eI3G5viE5p4adHcaj/mvh+femnwIgku5lOqKfQRBFRv2vF16UAtCBd6YiuH9Bc9T
awkklpypk+UksRn0kbD/oz9MQrm+8/VceT48+6ZFbDTPfu42Y1lvrfvRo/1CCZWa
gioHAyu/hkKoeJSn2u19Zj4niOINdNCrM3NidxYBNqAnX4l/WpXJtIaEcgOsZ9lI
J1e5toEOwSRhIaSYNr+R4uyoP6U42n+KmB3YzkPGSl7fWchl0+CDLtTR5QDgOZ58
hmtMOhkW+K1/m8WFeI7jWC3FUeYu+w5vCHnivVC/8s7I2zsFeeUdM+0NCOY4kkvo
YYCUFRPuui/6tX4/Mz33oobR7VgotfM67dgY3qx/uDQ3/yzZFfpnd75cZRe2lNSn
D53UBGWOn91tb1pce04NPMWcWp6F0ovYnVociInxIxMCyuPnITeDYyj7sW2LScOC
KDWvUfluLeB1YdzsX4+u088kMMylfZGkH3iEMIVaC6yMdMsWFw5AL3TZZXKKPHHt
2jdJ4tTGAPmdewu1ZpvJrpgfVdvWRUEBp+2Dl6cOpAz7k9xpYTYsCLrll97mnhw6
ppd5r/vMw18ILaoEeZ3xd7bOiWjFj7vcUVhMIX1X73FBwgisqpDQkvnLdZSzfUbG
wwq757s6J5mtOM6O9tf/6nuIch2DmMN8cGrozT5R1d5ycubJHH/WLG/dhXK7SgdQ
gKO/bh2Q7G9Io7oUswnL7xACHX+fG716wnhtD2bzJwaePfL+9bB+JKjq3KR8mRgI
/Ql18Ji+W8duf71gYM7cR1JgFdJ6Gmc/jX74NNWd0JUtL3Ib0O4/eHfGE3Ik15KY
woG1uKUcllFpsOk1xYvNSir+LRhrzbvepJAC5DEomG80WYHosJjzODE7/WdJTGAl
9lZ+idOuUdMfFh/ldVCggNGU5hEcwd+DwdgaLatLLPzsKKICH91bh0dCXu3U4tTI
BGAeDfvV2K5+Xc0rN2AtLkxjAwmIhAKLu23Cgyf+Sz3N9xdHy46c9rQZ7chqPrvT
b1EXgKAOESKJr1+/qSd7by340a3xsCQT2IDh6s0tJfBre++DNhN/PxiYalC5rGdA
dgXN3fxTrdbttEB1+I8Ckh5d/HJzUhKvLiArbEya2pHrtWAiUlKd7tovf9fpGpba
fswwsPQqVz6r0/150t9LPmHmzKD84/P9fZkuEEDyMvCvnh2NI1+Yv9qPKrAUzcWx
adt4NQURvI+S3t8wYlTP3rfNhPwJb6rDSio6C2hCi9ouNqw1yoZ7q/sKnszywIH0
YItkvKwi6TAtKt8pXc+FbxbDSNviK/54f6jImZGz7+xK8pH7xOM5h1W+5byZokUk
MAuX8tXfcLhNAtN0m3zgkV7VDdhuY5jIJTDgJVFGTZR0YYjNHDmp+eJnDdCjv9ZH
z6zQnTZfrZaAX/R8QIzM+QDirNkFMWcsqBvYI2GsXAV21jL7RFymPwkfJFuoLG6p
MOciBnAB3jJR3QvqIQbwAvmrM1FyLGzIjX0BByB08JFRJXEY4HoJZrfmden9IuIU
feYcnqnVwIi03yJvmY/z9TIU98lkGiKXoyAaKxuXy+ZzYo7/o7a6JsIgs9CS2Tih
2BW0/CFbCgkxACod2vj4cEQQTuaaNv3RAGhb2XmeS6deRyB7i0xsqGMxW7xy5rPs
KiE0DvYo/H6mzVlDpDuIKbMAKQ/ZOwfoiXJn7muOkpop4gE9lj1Pfgfai7XAv8bG
chiR8ydVlS9le/qOD4NDXsGKZnxxJCfDEs9ZGOxDTea9cd3PFPA/CW/Il7zhzX4s
IxDJkB1GEQGcQZpesVwddj+jrt4FEBh3bWiTtYaWKphe61DjXsalCSLm+nmFEmrw
hzb6xM9Je7aKOSdJwnkfy5+ohUTk5F2Q6Ioj4TD+L/7WaKMPYoHsBSVpjmvo/1Em
v8TTqpYiZD0Y7ZyjtrRyz3XZc5sxD6sRHjj93FJ2uuhXSGNEDkBjNxbw0UMf/Sp3
vphd+3mn+hf7kpe4NJQr+KpDVzyaHEewhMJBdLfJxj7CojGA31W+dOUz572sbS1J
Li9Hs8lBa5fSvRbZ5uc5Op6u7GhOwX3bAAAbkGkccD1uL9+606x8TvD0swZomMAl
UKI9lrYtzcjb8wyQrIQRnh1ECF2aAbJv1OOVqJqrxqvPAk0TqX4C7CseD8ECjQtk
IvhCK9Fre0+oFU5sYM3iRa9flRuxVOqTMvDffo8yjFiGsVnyuAWuHXjLQIztGV2T
4plFfpW/HK37F72GBWY4DhR+Ds2MLVemwGsl9KByiI45eJTUjzmTUcebZe6d7RG5
88ps8keRttNRZ0Gqm5dCL/CWrG/V6Eu08XfZ0MhsaDIAJ3qyT4et/g8X1ZgE4ji/
3Hf3M719mtD1gafHTEVRGdZzR1FW0PfWPp4ZmIQdl9lmyMBDPsceR4/SWiJJND6Y
s3DSyrMNXrX5F1tORRH0VQ3XWR5nAqRW02pHXW1wk6xwIsnneDejgOGLhZxRqCUV
IHjAcYOsHClXZt4dr9ZSxabulyRe0D6mjxaexc+/iN8FG7SvKA4ncnf4CJcra09z
koA5ViyUE2v+PeLtCHAbmPvaIYD5ZqWZI/JfbXUcL//FU1QmE/UFtgZ8VaXRkyMw
OBNLODfh0EMUHJUzz1rqYdPUw01yUB4HLYQiF8Tbn/YLHL72zDKCtB5qm3+SGgY5
0T8unUmKeTyZWGIA10o3if2YkB32bcy3D7ELurl/XStrnc02ds3b2Z5zYxumajpZ
jOGzpuJUauEKE+oYY/qoFc4sh8WRPP6LG0OQBAE6OS1tT+WgJoZABU4fUCCIXb3Q
4ZJVemIQzSJA+PffYucudu558R0JGA8Wy7QFz7PlUNlFUrrv2EQVhiOGPz2M7Dop
lP+yZMrCKuAUaU6ZGaa6GF1YxRtZ5CDU95hzPzT+zIRaA7s8MT3uyDKNvuFcwhuo
ux9KbuKhBrrKRfUynhmQYkfwak9+StzhcZK07KI9BDRvL4EjwW3Kk5XTALa3Uhok
DWQW74J2ihL74MmPCr94jkfIsR49a+/jzfhVmzEYqVQNGUo25BO+6BkgLrRifxhT
phr+wUMC9zA8Vxbx1cYME9R6EvnrtpeYDKWMJmciJYmuZKCTmbEfyHrOphVCnQMt
EYfMpGJiTfPa//Kg7DRrUYHe5I1746q8hUBCZeWMgzdJCxMZDJPwLDxt3XySdYNM
jkuyYSsiImRLFQlj0MzXwyz9u0eTfLHRI5dzf8i1Dhnj9yhOSH7TMu+4K9q0f2n9
e68UaIrUcjTCyP3T4IYUSKUs+9NKiShznC8kyQ+ghVxxajFUsaeWZ/VIBICpBCHU
m5NJtF8lSrsFmP4BV5zFf/T0CztG5widb0KELME90YaXsg03+zOrMYc+JPslP2FR
ZSLxvbylGVgisfR9DHsQ3brFtrqWzvON5z1gYImBodLapCZaGlscoc0jROIz8A5l
VQRwzpftNY/OmOJxiYBNU0J69unkLDTFLinnCAIANr6zGCmI97mnH3Iv9ZW0uj57
v5V0T/AjyZ1BEqUReN1uLbkK4yqHt9YUgvNQ+fObtAMsyfAincW67zqQ1Zyk8ycp
IUBSQVpfAhEoXNyaqmfAGed9FKPvMaT92yqfpmo4xNyxRkmBIoSDudwkW/+FZuZR
7BlqCxa/iwm1glYvgWUDIjhqrcA4qom2tIbl/JmwXH/qRBCxPTwN3z8YA2Te3Uui
PgVA4d4aQEcm9HSM3JJB0tksAZU1xknnmptFlU2brj5KR12y3z+6YEFsv1jP/Tna
TIDKMxi84MQRrFh+ZJZLoVULH7MNzOnxjjg2Kgv3+dzgOGvmWIMvJWD2yIEY3AYZ
88y9zqPK2r07QTfAwEQ7+d6hNm7vCg91r/RFUsTv3QqNfL/UdH/MyTKoKT8uPN8I
7NvvtjSY1ONBsEtDNjRsI3M1sGvosXNHDORDdX3VdfS1wVwEm94QUPhgYjanBoUY
82LelNQ3PCysngXBPwYP7mB7LEXLnXng4eF0LfmK3NYXN86TUyaClxgJ3pdrl8G7
eL9v8KaIJS4wrvc2MCC0IqmOyUfi5KZrzv42tyDNMARkTMaR7Y4tSmQaC6XhVWcV
gj32iKoFKQJj+/s0uOQlh49LLmFkes70+w/6nZA+RqX5O0Of1tvpD7+acr4qVPUf
yjx5ux0yLOx0XAeXDhlidoGrNb3mKnF9kCpzqnxM34RUg9eZeIbougiMHrSnWgUc
8KFkIFm5EfH5fAFcnl4EouYZJbWMpZzeF5MxM/dGdbd0CVfPtsO/tduyipQmyE5c
p7qvcbGONvgW8vBuMLWAJ0VeLX+9QhNbxVsAs8y9s4xin9qQxASvwidbrbp20lav
4QomPFvMk2zgCxro7ceLZ7E0KwD+zOjmvV73bIujeBaapjfX6RzbFTObUC3/b+QY
PH1hsxEnA0SrsKmA+VgdDVS19unOZeSbrtyLDY6sMXi8727n/bt685NZL1UDF7H2
EahnIEM/VDzDX44zy0HE5rUfkgAfyNFJ2ZSOICIReMU5cASRjfiankzWGKOSZX3E
8R5tIhP9FW77SvRaAGCJOiYEa0PY4ll1e/8NyEHTiVlJ6bjHgprEiyi3PVzq3HRU
DuN/zHZKkeF7foKLiJdqPWkY2IKKhmbkw42+YIpmGk7KKGMeJw8xoSTKmhbTj4PE
6msNTM/kHWv1nmpwYid7f2knwlqMujT7xhq4kSgpfbzpz502if1k//oGhQ3ef2Zc
1sk3Q0xwMEoamkMXERkzY8ebaorqxyGLlErPBtfwvZ/GWLGrEowoh4wlnzFfNui4
BClB5OoGFM3oIdjA+0RiOwyf+iSnGTBf1I6xjm/qn+LOoWv2zMdwENK6vyg+4Y/U
nfV1Iybz5jrfWawgY4QxQm8LCOq0nGuuV4uayGJCYdgoXdgC2X7Yr7BmsO0KUBrt
LeYUPTbBx6oAtmH9NzJhMJrOh3hxC7z5UfM756RuISHSDVPuH/RdI0E+A9KEErjf
sfqb95+n0tnYM0nx2QPtJSqRJTahDvmDljVOHlk24dqPsRpOTkisZqXulPzYOFx6
QV26m6bsw/Vf5qKyODk/xkdhT/jPxTviPf+KcB6PQaoGm6bhp7CQcIX4f7+qHaPA
TetIg0sZK6KF0yjBhPLyvrEqruRVT8+3d0RzwtSx2/CPs0/iNk9uZlCbWvbhnDk2
QX58TaD+d0oKIuVTmZeLNSWF4MGUOTBhSww2UzmAQclHzxjfppvDgSQTeol6RJxv
YOulMJ6ZZOYWpZEf+r8TaALgGQQvRhfto1EtNf74eM5CCZ2h6suLcHhXWua+wbQt
QqfXLOtVMs7nsoPXzk3eT4c7BGhZocw/byZLKkyGj0NDq3OeRvA3qrWNY86Fs5ob
GKa/C0sbAxu4yhbqMcVAo9Yy/Rrk7YjWQmxh1rIbrp5vT0THVECqUBp7Sh81kbKV
ISvyZy04Dj3HQuj18virDRhoxHz0MBTCrUMdxKDEXirs5PWc7ynJTrA8GkoJ+jHF
m9OTFTNdAv4FBZsOrdh5OVrYYMQyTol6Ni0BJY9v2+2ik4Z45E2oXTDajxv+87qI
RwFGsiUOVJYLrp0SYBHojSmTcOklccR2e4Dbea+IlEWSuGW/ni6XLmPWq8FTdbtz
Sq8NOpCfWxIhuz/sA30Rg6XysOlKpAc+6hOcPtfekA/xOE8LfGyLXCur+q8kS5EN
wx2OCv2KJRSI4/Dyl3VmMe2T0TtqF6MlDVByB2jtAFFYSyUFJncGlmM66Te/2ZHM
KgtJHIGgZOSAEgvZgBFAUVmBDH5a0bP9uKYlhxZinILak1q9AA8Q87K0H2tT1p2f
fdtwdusfkEgKN8YlnpHiqUMot3BEO0Yt0+lTmrqhsxzicWKIO4nLSC6mQNfenaDo
mSirtujDQV8tvpHGZw4LntXsFuF+z2ijg0VTBaA0Zufx6/muDPEIWLMdtHBqr7sM
ytWk+Uj2gtOY8//6HIREBUgdDino0PZ1nnU2VurqUovJsKy7GuoWrPONneduOOlA
ld8CpZcLhkNUBmckfUpyrlcm9flqNdpzgJFCawGlKr0+Tln7irPhqqg2W0EVjrF6
lL82BSYKZ8p+OXTSNR1cwWEGlMqkDof6kcNyLtRfSnTe/7pdiNtGxzSy4+3qu3WJ
qcdCiEn+9Xi8tIdsHfI8r8J7LCPLxYFI5sNJIC+pgRj27sfXuC4pw3UnTmHDE9Pd
cCQGs6l4nalLGf6Mw3r7C4wMjeH/xY4BZ/WiPF+wnieYbzmD1lo35Y+JMJ42zsA5
phEQxtGUbuccJcrdIrNqmOi5VDlaNzBamQRRqE79dTppof6y2cjQruqHbPSXHBgT
irDyT2yWaDB8jhqRU2VuF3s0cY0QafXHOOzIBe8GV0O+g+59pNaXNBRzlZv6oVxd
VH0F46KCSrMLPVIhmp6m8BmNPe9Pgz//QND5ppWv+kxar4a8XrCmhUnpkqTrurYP
x4s1xCA0VDmiowJWHUJq/Gpco5Vw11iLBQGOOomF8QQ/6qvxxXTE4wcVUFMc/2Gq
XbSUFThf5DRJo6mywEG3Mx2V8F/VPu5zAY632lCvEvzkVxdI1EQrwo+NLrwFCJQP
NUK28UJjB3Tw2iU4auSy6FMLm0ZJ1Idxc3ncUBQFX0mGapXFRE4DsKUfEFtSkt11
z3rIn1xQyNngb8r5rZudo6JcIWYHBsy3gMlI6Afm4usshcconEWZBkDmocmfp5XT
ji/LrVl4nmXHEKM8ffzSfwnHyBlp64Ny97JyjT+39r49fQxOR7rPCP88BIUnau56
A7FkWcdJiwtfqP+54FyAZxehU1dN8zOgjAjtTNUDFPpYX/Nnk9HSqDFOAEMqyfgh
B8sAFkpRZntLuPy+9eHLYyWun7CDizh5eJRUYFMbeJGBV30oSCHSuJFzpBr5oKWv
TWICcAU5ZzQYVnOTXIPNUcya5lA0H9XOmnH9P2NepGH1NuhFNcVIcaCBr9kr3Nnm
pQzERuzg72d4yXtDBZwdQe9/BuVDkHH5bE3ID7mx3S3eiLmL+Mu224UZq8fu57Do
c0GRpQdO7eYvqIdRK/0+GTQe4Rj4Y639oJ5DlgaOTHv6pFgWn/b2KVvnuxTyhS1L
5m5jezbmigWRzFPQ5n4XtARl+QeoW4gg9AEDeYwzla6IWJqUyeiFl3HWMG1KKB2I
08BJ6ijeAwTXu2tinjpRUlmZ3ubdUWDOCBdRReFXDKsFsNTagH0HOx0byCqa0QPL
jkTYrIzxYDTHmW1ZyBYkSEv8SGV1RIMIr9iW6SwZ8bovQvrcNTIjZrQQHB750Sp6
+1RUvw38DG7OrdpkONfGe0QrmXfxbYWBQPqU/pxO6IQk7FZQRujX0FxL89lV6AYq
wCvAp3DG8qXTkkFHMuxqWTj04yy8DyOsbksh+jLgvMGOA3oxmcYadQaNKqpENgzl
/qxeyLZbC/XWh6Bjx5nhku9QWcw8bH69O99mRtto8wScdJeei8a3vaHDtLq8XTec
KR+S5wW02ysz1BH8ZGV/KD0oIBP2UuQ3hIk5ewZW2ihQo2duGDOzDAThyKvuGaJI
5DzLNr+u33NP+GYlosf1+weGcOrc1MEl7MY+Jh6eq7sAzx/t8cC14JgH2ECKzk5c
1lf8eR5NEUQbEs+MZjOsApT5IHpDBlLk+VQENm5yX9HhOCa33SG6dz17o579X0bg
dzFKGKZtSvf14tf4GELPxhdhmCbG347J/n62iVwbvHnlzfoYknEoWscEARaVwvcq
NPbEkipg96o0akN1aU1NwTmUsgJFcAg3GdmYZPzseKJhJ7itjBS37DSu2GxqAiMc
rwvUf2bBnMiRgtjp84gv13UtZ24wlH4T0hy5hG2UJdTM0Nx592fAh/KvEmBUHF6Q
ywOjWAS1mdsRTmfjlp4UrgfyrtDpsVKxFM0BfAI1HNaeT/n0vfCJqPIfkSTG7KC3
+pcaQFLUQvNfs26oefIyMvzcPnKsgvmi3QxlLXhHKM4WokT9re6w8h6T+O24oGn6
PjiH0nqOqrS4K1FnQ8r9MS9MA/AvKb7v9vBnbwPTXwhFuYXt3ymbbCCfin665+Ej
oYGPB2TzTojHKOEdB9Me5uShQt1ffJSWNR9a5MgclGcLs+8yXeB9ALnyM3y7Y4hv
Nnh/IyHTVi9i5bL0wDvBRFy9By+TCJGlndiB6hqL6Avv3oUDCbXwbPQn/8NJQv+s
J0/z+wGiv46JCWb8GYd89vCrV7x2roXXj3pUNHd+HwdW+OZp5qF4pnWa1W2bgBrP
LerKv6QGgTPSHgWXEqtP9krZE0XmYeV2v4p+vA13JX32RdvOgl/qANOJXYDGRupR
ZURVlrwrdDGIeq6UR08uZcI+qWYmrNUUkNPHZX3uX+ROx0eJ8xxiXHxscsguLmBW
bXE5q+YU4ZlrT/TnKEO2GOrrzu7kUrLtDdr9AgIlfNbwDyhyLmomsETu8zFGK8rP
wQmE+r63pEzB3PWEVZrpjEQCHLpPzgFOepj3UUTF22kaKAGAzlCGXSpwaFRscDXQ
ohQL68J1GhJ4qc9iEk0j7YFNO3xag44+5gQa64NSy634HLStd5lKaaizUxbgJ5gm
DyF1rn/ZCuvD0ICwLwTy6mnrgecEjjVVMi99B+8EkV/R7EpLCyl45dsrqRbE7DDu
f8ga/BOX2MSZ8wGVQIj2hmuErS/W9Xj41+6A2fnD1mVqXFNktl7mVN5gSIJJldty
te99biFLIZzoZbaDQocxZi4k2VgZ0ijCIGrgfiVMT61B65wvoZ5q7AkzVFWcx7W+
pFBPsHiS11QpoESqiUU3d8uzRlnWDkGhm8RWYLCs1cwKeEq6vhvu70kTxFOv4sBk
Z69e6LeVd1FxZLzkMUumc/YaQFw/oB4xA0EXNm7KVkscjCK1RyjQT4Z4lGjV+b1L
gDjt4uy73ePC8FgZpxxwhIo+FlEb823MZUrZFPfZDae0jFxo3jYS9OVaN+2AjS/L
+EsTIVqPkryUJB4ttu+I/RuFbpfbTBPCoadVZKzWweA7EpkyyTwagyrARiu+3TrS
Vsn4bu9I7PwGO0L5ePX0YNl/weKJzx8SvMvzhgg++BO2aX7nMKpVlP1PwPxsa1bq
XZivBSOIwTBcqor58TGv8WRpJ9RYRKi4KUI1R4+z1pCn+a+bJ62OwzQXB1nH1hHv
kgcrlVd3N/PtAwVmfGMJp4tn+HwmJsCl70Gxg+AYCPLpRO6JkZzo3Yh8JGMAkx8i
QnH5gNxHHcRR/t73it2YTqkXavthwr8q7P7tCF3sxKq9/77RdxKRfk0yPGhmCKVo
FTai5JZ9JMXQbFSwS4I7+eOQiVlE4i72AdWqNtL8h8uK4IXLWJbKj3dwk9dq28xZ
VH9weI1qJEqrDlDjWsHF14fNX/79zHazoJnSV52E2lz9+AtxeUxuONcLaSagzhsX
OZaNiBw9w54HeJaZs0Xa6Z0RoA7AWAONfL74dvhHXhnLNWY2PiSshBoUP2zvWt4r
u5WPrvDcN5ks4ICd3SrlicFJjfmvVZqRQ2t90qJ2+oK1c4qWPkGLC/0q1PTZ7PSJ
2wLGrghw5ZlXLjFjaJG6kEA+PVVGnfn6n5/pg21KEgPWyMBFQ1i+T1PLfOPyJ5Q8
ti4bVQpSdVu9pnEAtIJpv2qeHM8H4ZygqlVmKjAlumleukGigCFMXxal1AJukWlc
ZW5JaPcDEspjXH9AqkJ9VUxt8KP3FRXfjpgiv2bDh99Ozm2UXjQ+AtjicCSfIu5I
96DfkxzbqCnIPC2U54XPoMyZ1I1GLsKt6Kv6Kh4Pe7n8QcRpusdPfCYNfPPDXFYS
vphBziGkwdU5RRAGJCVHIxWmOStaovQFV0XaHwuj+u45ynuJjvvfkpYxgKAHfhfg
b++dfsRLkoARJNurqnqATUiujibM/WQ7BxReplPhH5SVfVZZl4ePSK0oX57O97vb
cKmgR2B2X4PR5j/jx0FqdeGS/3iG4EGd4HC5ABz/+q/dCg3e3sqsILvw7kHgCw+y
I8zslkKO8ok1r1N+KklOz5uRrucngShefnlaNQZ7gZ8y5l+VXoaYRuJ9YLYo4Rqg
Nm+X9/ABuYiCZzWM2nzTTfD3d+RMqHLiPEZTei48KTBEfdlB++hxenqautmOYqhp
qXlJMHmHcjuTTAPi/u7h/95RipPmhRtQEc34CqS/6tkoGOCTMqYiUPKDgaWDB7bF
17ztw85Jdag+2l5J+4Rd5Nyg0kFbo7h+Sp1leFCi+X261NCwVR9RgzE9iar3x6Cm
EKjyxClfX1w8NJIOU2qmeJ5KT7ur5fi+e1zQ7pvkgL9PdM9fWPJ7GCFo42/chfDN
8PnGj2zBFYBuUbJUqsRBeccoFCQYW97hwj9P71kWQdIuf0pdzCwQ9w0QC9ZVJLSv
I7wg989E3kwN22jJ/vbYLITf83oajH2Pc9v69wBZmR5x21Pi34zwbiiM86RMFPjw
ITb9FWVKNwduPm98BInIhdtw2d39x4GdqqW8wXtPWBKck4y6JzG39hPoDt5LvfgK
syVocU/pQkvM4pkjl60D6Dt1t5SU1l3IVquNleGkaZjgM3oxgZMDoFqXYOP9CSuS
SjixYMO5H9dhfbJxV5rKtFQZdRmvtXvbgFj+mBsKNGCBH4Zgql0us3J19Yg/FsGN
qT4bQ5QDba3mkx9t8pG+YdSNiUAMt58cMi7CEXPt3TYwPSOtE9iYj4STvbZZhNlm
xiTzEBtOuBuh+FPSI4OQYdRLAZZADxeENE5t0rBRUrenIIkb6Tk9ToX6AZB6cw4V
KL3WJF4VZOkiWBZAr4JXv5NNftVmjBrB+ByYeg+TiByPragGGGrzpjcgppZruLWo
/u/Y7NV1IhID7+pYafgWtSfeXu3gtMeEIhtyHnbsHcFpaOzyWSGZ+nR96DFJMGI9
Jr19Yipuu3oJMIwyXlN/i2fR7Z0h/XVmEdQ4IgzKHJXnoEhNHXPd1iGrOe2NoM88
3GZJxAcYrvl3KNkVUBhMci5CjcwI/upcgIK72VroR5gpYhS1uTjPukovfzFFNI39
MCXgHB8E6TRAldKi5WHsFkP+NUPAdmryi7DtNdU1oswvPG4rQZYt9Q8QC3ewpw+y
gCzN/6x8xf8X29smlXYyzLv7/ZQQ1Jh+oEGx71w+iEHihuVu0010jf3J3TdWBOkn
tirHy9pk5H1KGS6cuzFt5zba0rR1gEcCn9JbdkS55VKWJ2F6DmvlqxvNvqul4b4q
1xaD/0m3PPC9eTYKg1zKX6TO3LAxeAys2pQV2PfvrpMzBmC37oB8uhajfasog9pW
c5K1pdz8U/5rOUMxJCoh+5WOH5wkkpMHN+kaqSMMVpzSRYVak1clnleDCcMwcXug
CQY+DF2KcniwspDqY86aehvpCpzPiqaS4hrxxgQCMqh9uNS88UAPlZHkCVvu+Ecv
4z2c4G3ytf6lFQrBTTlR5c8gV8e6FgMegPjPAjm9hym4Sq1bFfAWHTiawkyOweZm
1Ic+Bhn58vRYF6seiXdoAS0s2tAZropUvdR2PZbk5h7VlJyB0Erz7UKmXTRf4ier
ZoaM1FwWBgA7ccwPBmmAsB4z4hs5oFEuY9HF92OJb1cn7dqJoFtDdGIGSC6c6ImU
8jT20OJgzDXjF/Fc+7kfEhdsF2c/idrFbzqM1HNhqZOvZLLRYk8HdrvWA1UYgWAY
CTHWnCSJME7dMOccQUQOMldjLdbwyN2t2fTAzhWLAWboPHBJoIACu/GqnjoWuHLF
VFMqOiUb3UjLqhvOuefwi9gOesa1ygcPfCrxcyBBM5xC0Bq92H1d+T4BLKZBaCOw
aqRc5XTEFXXnHU3nBVj8T8vlkfqrRH78CHfkDO/h48Wuzxx0gaj5U+TpQqIUbsCb
1TdLDt7v2ImaO5fapXQTGyOJHl/B9MpXJzgsy6E6cuZdghwSwrf/mtpFPY09lavj
nBNSAKHc9oaheVkSAELYMGNxynQOfkuUsfLUzZkF4gKlBf4XhQJw8NzjyZpiCLPp
xXf7BgtTLSw2diGnJpONBT7k+PvMfaMqRBO1V9jGEqHkvHIAkAX57SpIYFPhvvdz
sH8lK1DMd/8lqvXaBzGbKblAnFW8kS0gkEBilFd/c1zYXsD7PAxPx2Xhcw+GVBUd
6Axa8JPnf2xlf4TmMkxguTeAHY2tLaLWCwVabkM4CPwqGpmL5mpjeNXiDOGRteVa
fY6cC0OhF+nnEHIirz6jVYht/yv0a6soq/PJmEpnk9rS35bhsNrKbLVgoKzAOQLx
jcA03AUuiSFU5QoPiWdvapwFXNyVASDY2H6greJi92YthBg6cP/+jZqybop5cr+F
39EjM4mJ2ccGDB+xhEgkyzFV403C0hYv0XwqzpYbLumF+DmsjLiEgGbecOUA28a4
FLsFq70nKCKATR8XzLSQ7PX0jTzMxtq0dM+E5RqYpH7ohU+vFfKUh7sFkZnNforc
e8P+qebQ/S1jdF1tW8ZoIFGXQamzcYsRxqrU0rvlFGxTauMYWsVDFPD+GLJ/7XgC
EZWFYGiFFcRvgkZPRyguAs2oeTng33xjCheP6TIWlWNFXjK3fH31KoNtSt66yD1Z
F9R0lEKrvaajPBwkt2ZU5ehcCvOetk1qVspTMVINuzGyp9w4UOK2/GZAnJEXYB9z
DEoV4MqO+3/HTi0pobYB2xIz8Amn/mVcBig6cmdGDJBuzvqG4x/5QKPQALL09/55
S152ZTz53vfMrl5R8OObhXE2KRDlHWbnUBGiPojF+Mh6+TZKPC1CK7wq8ZTM/sm9
GGxHplbb4/yEGE7wnYOCvD8Ao3bjfacU7elLLhsDRw9XW/fVYRFOxnRyjjid0j0q
rA3LmfX4i1yFRjO+TaeCnWfmUxVeoPTmBz+uunF0lPIdmRFIc5nOstITPna0/Zrz
ImSaZu1E8RArlmIRD0m/CSFqK8kj3YE9w7qaLk+gXre/AW2EGRzPcamKZ97B3shD
2dialfkZ+AzxUQe/uqI7YzNFEnTVUeALWInOgl7qxsajmEK1Y6vSzyIlzX42zmE0
2ZuVvUsQWZY4nrEGYr7BvRN9JMtXV5ih54VvcH4xVwPuUt4n9HGV4625rap9WQJf
K60AWNxOJD+xiXmMJZcGI//eAWxgb5OV7MBM+NXBBU71TpAmXwIx8eUnE/7RSElo
nh8gLSfGxLKCsZlWx1QOiumwbagL/iqrUaDYdKQ+HXjlPmmaLbb+PcJAR/xsWoNX
9L9nXd/9Jm7eWjocoGWzjGpvG8Av+0hkfcgxnqVvU2YxZpAMCVL28+WcVyewi1Dx
CYFjvz9vc66HCSw/I/v9aKYDENLhNEpIfmuJUpks0S9vW0QKHuXyjLJId/RLxISp
Fy3lJjPXp+oLLnLHE9a5DgW4GC04NU19bWs3PW18F21mFqeDie2ws5lhrSefaZ6L
oWZNWnfI5ZnoQn6vkK60zRRckSFM9tPLvf8icAJWJ56MgPsBdzrAcL2Nwwkg4LNg
S7UEGA1ERjgG8WNRW8LL3P9gR7WAQd/W84JNy5bYhmFHwwTKRHhIxbIZRAL8IZLD
kE5f9kSFbSV9fjQHH1/GwCuf/4M//QBMK/RjISziveXN/fQROVxoo6tPJvauubfj
gOMFOmXjT5XtR/aSqnksjr7TPfaEy28SrkHUoXKjyTmspuu/cAt+cGzHDqczmLWm
pfhvpTkRFIJH6B1DU4sbidAkddUDvL+TRU/m1L1CYZziIo9j5yxenC+x5AegtfwR
xzbzV61qtWPd2YaKPpvhEAsd7Re7G+EnQvLFHMYF81zFZRtyewObmOT3fc1Nh3rV
mTPowe0j75ZCqqy/KCGFD3Qg9qmTxVkzkakFyDfidBqR15JSONpHSW4xizz5lMlU
mR4gTKavA6huqrVHWooD75VGAZt117Bw3u5sqhsl6ib7qgv2fvowf8VQKXjxNN2M
V6TzP51sDMuA3SwX/BhJNg==
=======
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 43504 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
u6n3zq+imfgUTXW1Q5t5Cp+ZBwoXgs0ONrt+a69r8W2+DVVKd5Y0rNS4DSjoPx0A
Ulzdz1kdB4F3Gh3NUsnYH9SL4yenSHgmNDWMnNnO2IRi8VtZKXFlhd2zbMyg+IjI
Glgvr99wsp9KkWQ0FQogJEn/Fypn1Q57mSuAgK8+pxFTGjhCU/n7lsZOsTdXpIi8
FxuAkMXPL6+7t6Ofv86PLzhKcOt2Qu3m5HU2RWOJJ0PuM9+939t43aNtJoFMUEh3
uNZ/BBxL28eT9Hc1NbuaX/Ua3eOZhQJqvSTSAQBPUMYpwzBbA9A9CIDEEP4tn6FS
+HLAapqKH7g7jN3wiTXaQF8SgYv5/oBkxN/BQ5WOzxnJm5s+1A1Hz5I4pvpXpRlq
2uY8uEN/bLjj6OR1BB5sq/4L4boSjSWpPnOyFKH3cnXx3tVq0VZkN6XY0kWlqGav
s4G7XGAsbttzUP5WgJzEteqbKN7KrUVbHCjt19x3j+imd1Nb7rV/4pLZEVtxmeY+
1BafaeWkupT9ilcgK7YEIg8aDKrvGviisAulBEVa5KSzuQUsBggIopHbu9/yYC4e
6Nq5mbaeDL4Tmhc1GiamOuCeRFR5dNuQqdN20EhKMBrOy8ew6Ev6d07FB6DSIOml
Bvc/ZH9QDFfi+XlsJClfMGyp9RyeMHRuiVE7sQal0FJCkSHP2dBFnGBBTJjtJadY
rDKMYrMVGOAimkPVp0nIh2fInjKlkU5hFNZZouJmo86tW8FCvhEapd5PldhRuliT
AWWCiJNZ+J6N4AhW+IfjV4orpP8uF6FdiYO7iC8KiUjHIigMSwf/YAB1ElUb/JE4
80d5Nso+jlMhAZkkHdtOEGVCV7z5UHHlLFrTYhhz7nHAFL8KeJI5OPstoFgJgqXx
pBVgpK21Dw+/IiyRIS7i0c+iSOhflZBebvZbPWmvunOXR8cV6DVLTK6d3up2Kz6K
JqL4jcYe/SR8LHsKt0IqEVEomUlfbQyV749pgMImqFBU0eCibz1MCno5hJglTxFQ
EwvNdOkFFf5molzf21lbubtaVohvYS5vyxR1jxp2gfAPfj5VC3JNo9THZiQavbwO
HYtsyNIXSbOB7wjgkeD/BNxdzRREX3Sf8/xVBEI7JSvjdFfj3eD2BkCGl5Mq3C62
Y4yumLV/SRhVcj3xfIzPvdLSmoz0vKlfDCeYijKqhumixbCzhUrN3Jkmn0dbArBw
Z6uKGYpn5sff5PIuODD7frCuDt3sCkr15xrB5C4hVhpj3oFSnAHAfCPr4Qvu2uvP
xnzEO3nA7KwyC4iLFp2no7CLRdEWa5SYNiB7fHxfeWho2bIORzrvvBIyevLt5waW
OhTfn53Nc6Wq5I7kSmMu3Z+VSQscrhpH7NleaPb2nQX10XAzVCOQee/N8HUxMArU
aLWxheenNfB1jKY4pNVZiqkOHBmkn386AcgrZ21zu9sCqlMoeFAsu0NUJZVZ9Uqf
KH0YbP0M6jqm9k33OYMeHms+81rudM2dRTx7UJXFRUrMrTa6vCKbx0sc9BfR9fRT
PcpHPGElP0TFPKVP6j11p/Fi99dALlXKRiVxlw7fgoq9BiHi4J7GVFt9Et5orp3m
L2QumLL/+56vi7yWnVqI3XhxD5pUS+1HKr49n0r2WfecKWCwEhBzojlREdkuF+4a
vdjf9dLFGoXMheDoM+71EtzCkRqKPt/PybjwiYYDnaiqg6o5E3ps/ugDWGm143h2
+Qt61T90/13ZrDKAU7iXXe3OlsavkjI0hD9Y8rvjtwIvZPWnnJcArcmmbR6nphC2
gs/vB+2s9l0k0UP5VmBWjuJEaa1ZXzjPipJU2XPgDdxvUI85vbgn/bPXI94hJFPj
mwS2Y/wL3gpVX7kQc+Tveoo78ViWaFgL4O1WKuBrEaBcGqKkHaK3CiK9m8whNAqY
pYlG6STF5/GQmUqbW/qn/ljTfhqgT1Aay99Vx+wERuUsDbAgP4N+U2yeD0s6ruzj
4on+WwC8gfzzKc5dqQiPpue7VXY13p2QfRh1+RZpnG7PXj45MK9Yodb7cOKNkbCQ
tmX5SMdQFO3IfB7G/v4v1IoLBxmhxW2ULw1ZO0azwK6wYk0pOe6oDjxTcswuXkUf
h84Eo3HWouEua6HWOCmHUw9z/DVPLl5Fh/lo5G8BVFV9RCPpsH23AovpRmjDZkQQ
bDeTh79OkjMnD3NYTEZKXDgzVngA//6CxU94HoeIj5JBrup/JoiyVxCE2LiMwwhD
lRSe4oDNvsS9bTPPzaQUXD6JfmBWmmvdmm74t96m08bgk3+9iqLDcdKHTmgAgZJD
Ls9B2vqWJvoNkqDSLbxyiZmyb+oTGD45XjmN5WVKW9nss6SqMShi4HTYiOG0UGoO
/kP9iM/Ck/8/MRX/cXFuSzfOmlKGaUWirIHupX5SWWUSf93H/FTzrSxuxO5ATxP7
5ovyL6lPzO4H+rAzLgACsdkICg1IZLISbsCFuBLhz+bNAr1fox0jTcPePMy19wkF
d5IsQrIs7L5Q2LiQ17+MUsPQqJfZ/DF82QzjcYRBhOVg43nwFIpM5lwMZxzVqJMz
KmxaAK5uMAJFCBhly05HCPcPn4ASHiUHQvaiwJHC7PwuWNcPK9j++W5VjA5WbqSM
f6GzvbgiIyw8xDQXGK2TYVTrbzGOnI5pNMEJ4HewT41uJep4A308K//R5LGEOjmr
a/QfScD7Atk/aNl0dGSajAcjilVZor8QOCr5leMyxsOzQF4LyCTm+eGz3qHVCSV/
ymS13Oe4XOvtD+illfbtozNdEyj8agbJBhddw5FJRvsei7RK3NXQ123sV7s7ptUG
A1Jx2DBzcCJ2I+W963jvRnuCcgbPLaoT+8hi18pgDEjdeTMfcYnxsrB/eLLsMPsj
goo7G/KG7WCGcXGea4Xt+K5nWX1FWl/oijDCTGyqcnO65ZbhXcM8L+ZTyMfnFHlA
/FUEyMf91uK4EhLIw5503Z5Tjdtql5GWBUjt8pXTYGf0ShgycLtMmTMh2Qf/Zf/b
mHhTfTWS3txyX9X7AkzoRLPHEUX4MR0aFFwFeyFbyS9yOM7hHehzNUdW3Q+N9JBN
9mOZMtcpVN8DPqn3XGPKVC/RtzCW5yGpmKXzQgc9ekyB0rYLsZA9nZCilPkQiNCK
QciViV6kvlBD215DHCbOzYuZjVtLGDZ/qjdUTN9RWtONI8OaeoyIzhnF0zIYlnZN
P/Vf6EeVNz/Mb/iBL3VnyzBnHXRjvn49xN6o8d6JDZ/1vg+1zr/Vmkv3a+RFi1g4
I/Oy+gWUt/i9x0VfFKDxGk/NXO47SiG6Gw58vON10cSHK57BjvrEFcKBjNnj9dds
Wv/vX8qHU8wOJifx2zVmmL0Z0H3aWhvhRW5/s7LqAJ2F5AUhEnRtyjcQIjdeAjLc
lLA2QxuSJFi5VXQsDCFOl7WPUkV2FpoMfOTkOjnx1WNsXsPOPA2ZZqIOM+EDdbts
NsN2MuX2HuLNBiPoj8vUz/jq+YGXQWWk++2wIHGDo/oGRviR1H7gl6rkGHHtzQKV
f2S/HUBoh/dnhP0CK7GXcvPDwW57J3ydS6MR0yC+WhhdNeAq9oMyYzPvn57PYeLv
kG2iEEWn1OQ2dvKRX+Vkt7QyT7V8K0hiCkuRpx99tnCZXQ++x0ksZx7DE4VEGMFT
IkK6/IAZeeumFs9G40/mV5N9Spx70rrSTe3ZUC9v2EsVNz6KID4p+itMDpr1Rj/6
9BY4IYikqlExN3MFEBcnHSbX+Wr04CX4JNjZT/ySdYetTMj/uOihpXR8hNaHmLk+
rMTagnoiA9EmyS6ImA4Dt2PT+uUNp5z3VG1jyhPU61p03IYvUVnNe1CXTd299EnB
7Rn5UOX4EFgcEAxmcjcowhHjwLGh1M01TxkoxXrS5+jvcOar88FasCiMmPpn7jZD
1O0c3KY56y1crvzzVmfYA2tDrrO0gsVtKF8DqVnpIveL7r/fF86Xle/LgtIPvVEo
0BfaO28HdKt52yqkf9vFzxgoeFpdIA2zjr9fGbFKw/81/omR1h8cZG0zWKYl6NKx
E2AmIB0hY8Fsx5hFKClFA2llfD6x+06SRCkmvm6HWfxv/RqWrKY7VCh1Nqgd2xQm
+cHayjJJSFFbAtboloyFDPq+zqYJJmbWYpo7aNlWP9BFdxtw8G9HSddIVd4nQsVq
GKCBZWwO93dIbhMX3sxGvbFBXXf0J6El1Ind6CvOajkPbeJ6neQfEAIQUSoGu+EH
Gid94/SxMldTEwHICuyYQe/nUOwm0cNTKQAVTwdd9K81SDnX8ocqvSaTBh6/ZBAL
//b8jHtq6TaKiQEscY093ZSpeHkeGLZhk0DTI153+rEcJ8aPz0E1P8x+D35VSgt/
RdlbvgZyXQvReiL0UCynPusilviZmy22ZySk4K4qcSrt8u/RzZ0Vi4kBvb1dtq3y
sV8OB2+VhBtY/Maf76da/k5Gij3ZRdwTULCSJw9K8xNGo8v/Z7pz/yZth7r1NpvG
bWhhVu+VwSAQQ9KYB7e8arYkwtTs/Gt5ra56vOQ62G1YSm6CKZP5hEtw/2XN3AMC
3Fa3P9V6e7Dqur6MGT1sfimX36gSgfT38KWJO0LNDDMNCTGJgoWmH9BnbZmJTMe9
E7Cs7McHDNF+X7EC2a3d+vs4vq9ReqPS70tpfVK8xscrmJGBrgqxGYl6F/ll9elR
ZLJFLYhUTeUqtdAOQmz0Twr3SCRP8y3rvnmOa4HzdYq4yebKWFpoN4vodKq3v+gB
X2f9C9fLwCZhfH3/OBEncWjplP/GQJs7ZBoHCneY/3oDKm2T+ZxNZAlBjLboz3DB
VjLRgw4RL1lwxxnsniAMOZfQwTpFzILythl7pCEtiSsXi5K2ln/X2ZrCWWbuj5lL
RbJVIoSSwl7yXVXENXiQGkcnFX3FC0ix/kA9d1AGwOT2ruV81lkPTqxnZQkEDpqB
wqgXUIq5EsQa8gUmlFDjfEZJMYRvVObbf8MsGWUJ14lBesVoEtJWTKB2gNsl9ZMd
YIbpqtQuSmuAJLfKbaVqivAJrYnQhr0+WWXXqKArQj3QR0FkvQLg5+aYHmJZq6+A
uj0hrCBOykynqWm2K0OBKqJJT91xwZP+0a1zHCrqZZ3rnyH6VRDwGY5Hr5l0C59h
UyyLH+3+RkL3CHwRn1X8UBUlbYYo7bpDl/Z14dw88oiNktAjaiENBzMIq8XKOUvN
63KDRYWG9YULsV/95d+1JVNiUBA5XLp6nndJvPLFN9wBazZntqDDjn+fzR29w/NA
O/z0LfT7paHgQbc61ZQy2/AMNqFh8n1tKMFUM4W3hP8dNq+RUiqZa2TrpcFrJz49
gON0rTYZGvS+/SrLSK34MvpcTJgzxOOf5PqXoIF7WHzW6S+C6ZZQl0OAMftKR/t8
ennmVkJJO0GtRtCHopcjY+dwQB5ooDN/Iu3l5V4I5YinUxsWQiHXswKKl7TJiUMr
2LpNrdjB0WXwOPjpAtFI1rFsKcJdLAawS4h6Fi578++TH4OkVrdK49QGI3Nlpv0a
vEbAfMitws39iX2urihyRpmYZ1ChF67GpRPlRYovvUmylWREgYDcHHks6w99vukn
29hxnmRPZPJ5DDgVae6QNhPr+2uTtUSmSSU+5im7CcSEXb7RgydDPSj8XldmYmHR
eJLL+0wSTcLTEvKrt4JlaUEL1lAn24uR+q1o42FVrgZv67YuRAYepxP6LRHAmOHz
A3ZV/ItoF6BSkkEIgyFh+v+3zfudkinD4+oqxeye3qrGQs1q6quxt2ieg1wyvsB/
VOmabnKd1C72Vzda5cdzBuCs7Lk9F1SNJmAmN7qxZta47SJXpfNKyI7nIPhmQ+xh
FejR5c3x5ZOzJnb7NfRm7EHz7RwPsQiOZYCiE2KR44H42+rWuqJEpfH1xfqv6pjm
gCXg21ogt9NVTgZfpmo4PWXsPzvyHmsN9FvKwVMkUvsWyQI/kQ1b6E1Err4urYn2
XuVXQJa9XX6zJjJ8jZ+1qPO+Zfw68Oexy8IJMoXPa3TgY6Dcr7bSmOjGGKJ0ed55
jap4p8i6W4fpzKFezCfmt1RhuRida5jG0qpLgcQw4SrhdV7z4PQvfgCOgcTYqOwu
kMFgaSdcDE/9UqHHvObzjrKs47nW6H+2UAvzBa+zO29EsnwqFGGiZAY8Nfsw/dC+
ugihAYJ7R1LWJT5fzucveoWu8/LaawzKerdO6U5/YgeE8rKlH0T26XLT31xi55WC
YBf+iwbEu+/SgsBY03nruvD+Fbm9mngnoR/MiZPguj7Zov9EIJ/iJETlDPZE0M8n
eIlUVI5oFHeEE9j6X5JnMeeIDVAMvzQmoCV4x0bXEnRYg/NKBFCOWv2jhrUZJot3
QtTra99Y1fU2a9GmazlLcqc96ntvBQDnNdC5QsWCfFGc9HyBXdwYzjGZKudgZyw6
3yydMK2Zpj1TfKDxNjoDtYEtXOtoyMXl34iOQFK1TjIOR51XlqWZZEtFpSZK0fnX
JEo7HS/YFxCM8g6NsTG+ecTAFYdqjxpyKRTtpwV9qJrHRRBpDD3ocEMLuNUsu20b
8sUWAkNo4JkyoQ+SbqOuLM+FdYVtQgJTQWHyCUjj+hdVYGtNTXo+pVmXMhtA/ICg
ei6jziXaw8inkKUYITLTZg8xSgbLECrAm/+52pMHVGGX9jDSg6bCDR8seHowPZZN
mVlQIObvLgb7KWnBaYvCef+i4RSV6x0c+5S7DbVTowabEtnnDtqd0NhIXc5kjoeY
5yROo3h3mevsCBpaw/KvEw/8FGBA04Mbob9kUtIHozvg9aapRJJX7+4a19GxdI9U
AjnNVCa3ZqKpo3U8eUxMDDj3jrU0uxxtVuGQF2NP3EOMC3ohDuJu7knqBZFvinFO
UElvYpTGwIUFSpyULe8MykR+A1ImQ1YjTgIF/4xv6yLhsDKXiEnbHvWFkpxFqzxE
3WRJkFgZVzQHnNNr1lW7ljKpIyXRjC3FwHH1ZB8xVIKrKLv6feVxys9WVF1CAP3F
FqG5R+ZryzQYxJGa8oNcfbTK54J8Y/k97PEhv7lepbI6CGf8HAnXueMiUwK66T/X
ZRywzB1MHdck5ukyD3Y7Y6R/N+gnCi5kfEYWk2IfSfxVS3XPPiaHb2Uz+/1CDyci
y0YMQxvNd+04SS73i5Wo3OVFCnRfYv+srkwA01EweT7PlehON3jCZUslQvohKKj0
w3r5kLQ2Dkw/vcVigNcCtN+GZ++5LGZwbSeJQrrmxsU8yJ2nu7XhjhYu/6oT3Uc6
cUXEc+Gb2TwNVuYQvCLe5S8H7c28RH6wNTZWrvKdrzp+7ky8BIxYGfK96xu0d+Vt
sh4KJZx6gZosonOCp9x2graN33GOVjWIvoyGU6AmsiasaYh/yrvZrGSXSiBj2AAl
yhOlOejP1eKjvzU6W2lu+qujlbZsjkG6u0y4dda6t324N6pv/TZJKsRzrh2wYlBs
4Wz2bWPsPR2Q971te5UfLKqPW4UhcfFTD66G/pb+utKZTp39s8LslhB6zjfukDtC
Al78GwQ7yCjwlZtH4TlObyRFnAuYSLxHKSC3+7iZ0YkvAqWzl98M6vRrlITlEHPy
3s4IywqEop5860rKO/J5fDN+o4muMA7+6BoST4nc07dduhFBZvljVKK5JDiqM3+x
4rqA0sDt9Sl0Tl752Oby8htCKTf22Weh0HaGOWi+gYcCFa4Hciss+WNvZ0yK8EIL
hTm0zf0J10+gDc6mPlMhJCt/dzAn3FSYJ1WLf8eSIdU970Tq3BnMv5KqKreuXvB1
T9ZsKmfYAenBvakbosMT0oCCRv2hVKqteKMzSjKAbTw7Wd1ivbz1Wu/Gc2mmDa4o
oe2PJHt5de0Pjsdq9dfQN4+kZx/S0ZwOoGfU6/690+Zo2cFoV5b+dta066/6a5+B
8KUZS1AJa9brdpWH+npVzjbSxmBt28ylTEDRccUau2jRuvQBzHK4q/LzhQQPI+Q4
kgWYcC6fsnfBaFDu51kkGnPZubXIqOOAHpPEelZqUv3YFHHhL/bYuhXGY0aTZi/9
nYkgtmHEbvZ5yeNjh1fOEVPhGq7Xne5hUSB2hi4bJCLXAbIysuQns2Q3QAV+mjLg
6d7f+P+GDX+r2McxzxqY+N9N/nk7iX7RMQMGp104wqCB+R5t8ce1UUOVPfHIn4ko
PTSc+cW4PKFwB1/8MGYPJC2arcmdPjF5LtCVtHFvis03GUxSH7aoiipRi1jvbIfs
dUrhn073mt6dT9oNP8fYmt+IAClF2AlrH4RPtyLxUOnvuxfNEWtGMsRmI+qfTjKW
YrIB41n61lo7SIJ2/910+jy9urVs4b3G4j7ZGbbjMlImgKaSW4cY5JvtzRnL0NdS
y76PsvT7ri/YK9sPEtp008rUKfl1RhlbPwxfisc2AtKD48gM8HuQF9f7jIH5af09
rUZ7tp6Y6aqvAGcvIdLxfAlJP8y7+TZtb+i6M+33a8Dgnj/mOTOPum7aVkwQwIKB
u0TOJgpMOSF2+kdaIGZXk4GEITTzNu0e6i8ClCkGWIyJbiC46vnSlVodEk76rrcf
y77WPHBQhdyoiL4W/Abo88uHrPAxR6pNf/q7g2mnlTd6MNHlk+JXN4s+X8LiOWHE
pdl5LZRelSfrRKPHOjIzybwhImtrvuLejID4Io1u/1rwgKyznrWHMoaUasu14PrF
nRyMIyWRIfknorakXsulL8Ikqi4EeZnH9+FT5tDYdYg2jz435hXpo08+hgBlRpjJ
vED33QJnYeoLG1+ftg85dXhAjgw5F21mj6pz8Lv6Ppp9813tHNJ9sGCeW5Js/iKS
xDRfCvqMEP6M8zfwHJDbvFmV/ZI11dQnZPUkQ3FDf/ifJvJTP3/bUh7QbWD8vXAm
tjrRhc/u2o1bu3eg5U4D2gHjeTuXH3UV1peWRx0HcqgEUsIWIWf8q1tgo5s5TAS9
0v3eIsL9zuQ6/fIxsIQV2d2UgLjAk6FwcxgiqG3EVhhssGm8XvNmkohCYCgks+IR
wtFgnPyDkr2ux0VrOlrsg7lw5iVXs+Tk5I/xGFZwAhKUlaOQ7M9poQo87HHHp3N6
kfVv8wJM58hkiwa7cUQ46kLY/SPPSQjGSqx4wWRHLwwVFtytmAvIYpwWz+tvZ2/T
dFELZuJ588nvVzYW4nrxfyR4G4nh4pWi+Fi0tNsc0ruwfDa5foODgExKNngHPD7e
M7rKcTTLOM4+EWlYCdiDwMP3HCjW7hXxuIbVeWPnXzH/l/ErWTID7VFa/MXas8K/
/Vz8bn0in5zEwF4S3ejqn+7iAWAeQC/u93g0wFWcpYV5YiMC6zhf1yEhMWLY8j8M
rvBwbIWV1lUEycZ/QgpHERP9tIQtPJuyoZ5E5LEpOIAwKNq2W9GT3fIARcI68dgy
wqRo5s0+YfeCQb2KO16iAj3uw6Io2b8XPhOf3D+N+lrhDVT6hlycFpTiOTU2XJrJ
a0V/GL/iRMe7BLGuuxSvRH8vJ61p/KFv11HNLE02jwEde0pQBZYj4nynmlwehsyz
/qol1YZARmw7PLb98i+USxWElcCAhJJN3FTIHZPgiCiiXWC4uQVLM/IPLTtQO1FD
hfmITNSXxcUTC5VVrV1WLIJlkXLHteK1L5OjGb/a5deUQs0mNo0BgbESjYOE6Fg6
zbKwnOpR7g71aFeuTgKpdIdaepRtd5YkSNFqEY4DnHvj8MYmzIBx+DukEvevxcXa
2pt9BBrPCWWDBjdFxW3/IByNb/K/zdlLS0pI0TyDrJzo9mks79oricLQPBrTRQsc
OiSEFyf+9LO9DtnKPIMzb6T/ajMF6Uj1NFgOX2pemM5vds1rew70dtEBniTNxxC5
h/ugMgnRp9pCDK8MI5KcPC2x5pk0Ifj9i6bS6m6ET6fVRYwDCKOvsw2itlFCv6td
D+tAPMqWsUFwNCXfo+FLd8dJ35Tj2cVVId5P/bkg72EmtTz810hnAuU4Cw802wMZ
WbF5jtK4065kEkvCqgComfjSFmpGvXyhCt0+bbIAnwdWXQke6IWKpJR4An1mVKUJ
hgFvdFxbEsuxOEnmUhsSL4sosXQYIohgQud6q7hGVR6Y5HUJKeZjcgni8g06aZB7
M0Tnd2YQgaPl3oYJzbmSCjXU9BBG91epgVBEpgq45cmf47nW6jmfs9GniTdsegJb
1TZWxDAb/99Rjr+AdQgn6PrAPyRa+vApFihGUOicwBO2mBfVBfQXzYELcdWqGF//
4SX84s1bxtzgoP94uCslc+Ix7x67UfmS6fEVSmLU6woiWSLfv0FwhcK4OWr8zk56
l2ZJlyYl4Cra4W8x33Pld5fWyCmxWpEaGrWYsPPdKUvXi6k4opNGlA9lSa/rMQY4
a51fCe2ao8VSoxHvgzojPPB79yZs41rJ0Nbd+yKcCYBcEPBwTpyy6gYc3FSwN/6B
tUZ1G96a+Kq0R5B5qMcLE3l1WN2GDrBelpLZVONFrmDoaQiaWAq3Iy9AnmQ5tiJw
SLYTaof/AvEeho6aopWEa1chabVDumeS40SEbObBE14FmH0DtPtgDUVP0dg7mUQF
A10vzSP1XuJICxKdS1o2+v6/E6QuUQUGW07JjUkzRf8dyaHplzXR37hAfQcDyMTp
X4EUrzvcIJBSrOLjQQLwOdFgycjGkrwUZJf7ANayL/2fcCz60rk53377LELXP0xc
6URgt/QtuUX19/Gk+DL7vtljGD4RHj/BPFrShtKj9Qr7kgdPMu+nhbVyV2Ix1d7W
fDJ4v712qcs8H7DKMbsKZ0S9H31PBuq0NJw0EnCNNI0XuLGzHbnsy11zGyPBUJnQ
S62XN/NmkBh0J1blRT1UG3hrkC2FBy1DAG0aWIH/80B4lw8RJeCY8xXu3bnEv1Zp
QoIZbCfv6gp7jLsuycV+8K8f3fGPLaxy3ZVYsnMz+QQFJRIIgQRQQFPmdZJsC6yg
QsbLdgDMnFXVpkdc1DATRH2WMdxO0ansFIVKYqlktCcO6iIwdI/jTG47BOViKdiI
pxxDiFZQyeToMusT6II5vQDGeBBhxbUxh6rFbN0gUPxPMmYYd+lgRpR606e+PSB0
dEYWw3wdQubioaqiU0uq+eFKJJY3jFsIBGPRREG5t+k/UrpDZIjhq9/ePlI+7GQ7
clEOSMv3oZ8Eor74mActn2gS/j9ql4Cpf5Et5AI6YWevKYLwjv6DOq5/T0MjPiN4
fFaITHFzjXhM1W9FJueEsa5elaxPaPA2D4Zpyf3jeswA0NDmrXynu2EmzD/p8hnj
dXppIlfwvViG4b8wJVN66OoHRRQgHWdmnvZFUXlAQgt8UdUFWX60ix1i0QTxCIdh
m6H3cd87i48o6ZLW+3fRatSpv8FyP8ne4cZBZ1i3QCtKT22WCTksqm9HFQhTsI3D
KJx2HEyNqGBFVVRN+w192tLQhmJEeUQwA6FBz6inaG1m+c2huFI+BelydnH9S9uZ
XuGJH7ycYYYZprtdPYUuLAX+sSnT3fo9Q55OWGWhR/Ugsv+t1PCqXiOn3+8vI7gZ
bR5KPM8NvhHg9kSDJ6DASo05yLIb7oeFioUHpx00i534jYve7q/wSHynO5kksIQI
GZ7wn/1iDmsKeAg0H96oLWOFy2F6XsNqN9lApRkol2/wMWf2IMaOUYaDPrX+BSw3
vTnV5zgJ9e1zkmduKtbeORhlOQqY0zqE+I+2hSarVJzNgyzqpNF+wCMBfx7oeN+G
6LpNa3izBQm1fUEv+g8Mn/xOuMInW/7flc7fo9w/KLGWnGIGGXuhEGh9S6eTCW5X
IyuBxTQCLtHB94ayT6a9iUwtD9IlQgAk7yTRWMYfwO4GJmjn9VSADNsOMPFgDTsR
3I4FmIVbqTYopNcWcjnjZ0Xy/ADFXNdHKp4/d2NjXuvnfIJWWCC0jzOMSpXvsnZ2
CMmf1XtptCxrQp+tDMOuMWCoQATntoznz9sPlp+Yj2I9Ipkhs+B1AHzHY95BchGn
2NGFj6pJgbXAChDCbDyFLhRH1Fa87nx8bj+YZQSJndMUDnkAe34J1b5cdUqsWqt8
Pkw23MwKGFG+/OXL7wL+u04/olMORlcoj2EY2cOKmq+5Hee+ItHUdy5gLeviNgTk
4C0k0nM8GfOoAYkTir2Ma8f8J4bthGX/XcPjEUFg9fZYJIFuBI12zqkNrjRjyxsT
lHVE/z/di0aqujXVuNzFCyoDPtP/RF0IXbpy1Zv9cKXe4i6dsHYEwPA+lBizV+2A
3oGLwkyEZAbEeYiLBTfoJV5Le7pwAGOGhXUyVZVN1/7VRYqJp2lkqZEM08sOGr2D
uT6XcajYFfNlrbHlX/2NqAPIyFnrcoXCrK8jLziwC63lsjH1rv++Z4xruL16VjRF
rYNwgPg0889DHVtLuP2vrSeNsSKk7+B3xi+aCkp4cN/ip7UU15aWegesS1z7mTtF
IETtHOrD6yUGtIM/iLpwBgwLT212uorTNkgP1uy6n7u4pj0AO8kO6IP2WuQ6Pkzc
PeHUndp+z+S+C8pUu/i9GqkKaDPKyECOcBtYRpSTlvBncR18ePd++IvDfuUvfpsE
iKpd5Ld/edWMrKEQ5gIxJoKqy66/Xasg4Eu71tmeWRDkdyQ6SGTng5fknhIIMzA8
qRkrLthyDK6E6gIABmstcKj7YCkiTnPqms4Msu1TXK4EccpF5zwEEB/IISwoMHYq
3HE5lHTLQWd7oRrpCdWvGH2B6YswP3u+cJKYn95UeEzDJPMyz8aYpr6B6znwU9lE
ntiVAUdtfi9o5FuqybPZmAtrIAjLWn0ZzBEONOnCT3eqUNfJT2oQhvdoRwXQ14x1
0/119boitcV4RRfUDqGUX7XDy2GrCTUPPyZj4CrxMsJuJppAGX9E0vEbOat0Y11G
vCRNGdkl6xRrKvJcJxaCURLxXJpCrfgOosZ6qRPP9kazH6KxbM/a1Grdw/q5YCkz
xkJcAKeqEh/yVTx3Ugsp1d2Ue3PgAr2STQx/8ycUodmzBU82TLq42lyGm1ChIGyz
h5z9gcbd2d4XQtIOoiLbDbIcYiKAPNoo7YKd33HFe73cIZJGeaNRYryEbo8fNUTY
rBXjTFX64dMthqkXRw9sT5YB3z/DCoybPNlYH3S4pwhb6xWwHvrugdVRKVrG8CjK
prO2YgIxNpLQcFB4XhAgZlNslEYM6FtveoHVeXPTPyAm9z+vno7vBNfaW/tRa9+r
cqLO68bUudLQpADHpHuLkGzJJa84R5OIz15+OtImtkSbwF7Q0TPbqIyqgauOAJY0
OMa1NSClKEIgbFwuW1/3+FQBhC4ZtqNGtbtQhURF8BKvz8mzQjuEzLc+sko+kSh5
+a2Ko3KXdUbkdVxC9jzzIgeeonzoArqfDymXTctjtPEscfHCg3fbDHhpH+267N5J
ZJh/1gZARfva4VCLKYaVkVnxeNOqzUNmshHM2MS23p6E8qLYHORoa7+KbP097ocr
NSNls4wu/F4umyY1FQoteIQDzuSbe5MPQWMxpiPg9PSALHJll7CoqQRh2QefH+VM
y8qv/5ntip1aOoJnOem9xJsQpNosV3WrCneyz+ZPR76XHzCbia9/2dwiv58X9xcR
k3bGuHy/Dl5d8U6t8JwiuaBAU4LGV8BH779bO7V6H/RKujg8z8lrUoHDRQEPqZrg
q5NYbduzPc2AuXU9ndDRkUsyO6+rezZHu0C2vREXer8hD6qKAsNuKwh/rW+BqutT
i/FY4V2Y1Ts00l8w/jKNwY/hXSvXPS339dZVBxZi/dhKt2p27YDHleq2WOYMYBGI
kFi91YxibjbRiRff/aPTbyK/XqPf+OuGvU7kT+iDLJnacRHWlPrhxqrTJLxbSe25
87Ztf30tMeW5hvMPXgz4Q9/3odwwB5nRtVDIhM0wvQ3uBXmCkPYrlG5kCeHOPtnx
Xh3B0Rtkda2shdKlIEvEklH4LiXv1n4lzV9wB3akm04IR4NAPRYwX8GzQr7HfeBf
alWxJO9e7FjLj7DZbuHzBPhLUtplLcopDtPobhk6Udns/kTAznIpzsK9OuzOTZbW
aa8cdRxVMQT6R37sXNkdfjP4O7bwcN7oxh6rcmt6zfk+yZCY2iBnki4aOag61V5Y
FjOfxrUPJmb5nJRjMpGILVv5TzPUq3oxXh0VYEpl0Dvpz+FRWSsolgQs7nNSfwpi
J9hbru/GmJzQytACq76XINFJiATx9olgA+DdkqKBOpFtn/UExZ+vY3HVB5NnJgph
Ir3oFQALYaxgn3AOAQH7CInbnk9VfkP/UyHj72jSAhqRGvZ9O8dFwcW9dLyeLTd5
U76F1Hd/eC9KVznsXQ6Hc30dST+9scZJ7MboDDtuMpVksL5IETagVUTiMFYo0/+m
UdGOkz5EHTurk9uDfNR5vN9nZs8VkzBJnE3SSNlKj8GURIF5a5Ti0gE0cEgWmvnh
g5Cv/Qq73VEmNPNCudMi86y9yVO8jr+7BFMJMgrZsrpC4yURtp1+u5Cn5JDssNto
OWZ4ispqFI+pGXV9OalcXChxOHYfT0vD4hMcv3szFaFvEpi5gK6z5Kh46zQsRbHv
CrWwiFZvXoXzuywB8BDH5R47uPbgxUrtb6ioeqhq033yqNmU8oItB30wepqoZ5ll
TYIgO1G/jr//wqDCJuzMwxtpPcn1HPtGZ8InFdoi/ijdn8OYsekye1ZEOLN2v0Ku
rSGa9RRug40baM8aksKEDasrfKY90xGnc0WeB9nOpr/tHdUFOf+cD43Ex8BRbvB4
Jfvc2Puui/hqRyzWpPka8cC1EdCeo0LpYC+mHzNAAHccTS2k2wZIFr2ip3XDJX73
kpt24hx0ZceTJxk8S+zRoKN9pg6TtvHJFdyXohZ4vMiIsQupyCMh8m37Am4r9wMP
AGL02s9IKtceZ/Yy/FGdlrhn9v5iPw1LFVOTREI9X4EhfJgEvfDz5+zIdDGUsZ//
N3bHai/bQDC24OrSJ02P8D2v0+fJO1PCyQWpSwnP/6wve7gLulpgXDWELXIx7Kvv
jpraigaxCqZtAFOH8rb4tIL84tpsCwP4xxBMQXFrulD1V13gOSmkql+QMY88h/CE
bz8lkpnMcc73SJuUA2cXLGLh0LjrP0vz7EMpkJor3qlMy0Wu69uWHOTViAl08KAR
j4kqMLZzToP/onRJ6P5oKHIVqZiftQJyETJTmiLlrIatvxJiNG4jesvPNLSn/xuv
Gi5NG2uzeQlvOoaBHsj39YyLU3VsWU1WXWlXF/QYudcnsXtJO49uDl882FFc4t6g
uvHVxSHKrSScBQ5nBWGasnUxSlInYG59DxfcjW22wBwjKUq6vVkETj0VmHa7MOpy
HevC2g7KjRJ7lY9RG1guhaEyjHW+m8tv2XqT4EIy70JXlK+sOs6W9J9s7cvdmTO5
cmMER6hHpT3etxB/btYw4VbHrERMTBQvn6V6CMEc36cuDzKTaSE5aaNN6Xd52f0H
hlyJi11LC43Di6/7WUZFdC/foToCnHbjR0R441I/VR0980q2BMrNaDJIPSkHmWph
+2UkfkIdpdf+Pk7bR8TqMQXDtU3vXRZGqF8rYTodi2cdwG5CBO+1/KBiYE9IKLnN
+g69VrJlN9jUtOoe+5hG3WPXllWxes8cXe/b7jDWpejz8ZNcwyLBzRhkyWWeedwn
B3OKnCHQ57DHZXRN/zG7Inn/ZmS3AUXaOkyZw6v1NvYJEuW0Dng0QRSyLT7/3AQQ
AwE9v3UuwyXw9nt18ck3z2B8P19uEg15z8rz90JfO2g0Y2AMvUCMLUj5SSFY/gEM
aGEtTbXj3rT0zLX7X2iEkRkrP43zU0RnTZKeWVaigrP9OGOenIAgqtSU7sOiINpD
ADLv4yFHnryxExngAtZexwyq7YHkkhKj8BCPysAysWiY/3h9QXaCoTw5EMn899Hj
CBEqhGGanvm3+Rn50EVEDaA/WRRpEOAIrRWPnicZ6z7mhhz8/aWhsN4rXbSQsc8U
WRO6RFFeRuwgueJclbB/CVjLTFCLS+xtfCOQGmqBSAEyxfB7Us1ERoPPgcSrei08
HuaGcthvxO/7Ac1wxWTK43E9wSMGTdio19OBtCi1ZAuR28ga7n28jc4GhKK18bvt
+eBStqFVvTuM37jG3alvvlZywgTuq37DQG7BCabiJ5/SxhkFByiQErpRwUPCTxi2
GZE3ZDk8/puZWoHg4QnO/b1gRfA8iYXXvytt74Vt7XYXkwvMX/PZ4UMMBsDDjQv1
lDYmt3EAlL/ceWfSgi9MTEv+sG29/gbx50z6UyDDkoq8hbun7Kct0ruX0KfFG4X9
e6G4VCaw++UmO/c/CKvR25HdhWDsyMCbofv6UuODcWrL4wYc61pFyDL8VtmoxRmQ
awA8lKQdLhlRUg5wGjQq++asm6PBxtBhngvz6/jKwU65K/Mt3HpuDfOMad2nNrcp
QIZkwh1UhyVBjC4qM8Eg636+6WfU6bbZpon5tlNKBPe5jozFE9SZZDpk1ApVEAGF
dFC2MjMwvylo4GOyeO6EIOaUtK3b4ygUe0g8SIJxZ0qEjvFJLX3d15xaU8RmzPTh
c7hVzkAZqBcds73FClOyTzGYjzglbhd1tGlwa31Bz+rF+msUkU7+caQNGgYMe2K4
3+s4U1+SkOqwCxVAo0d/daTVKjb2bkTkkyVfPfcYZyKdu4SPyiyxoyIZwVU67z8x
hbfZ2V3k9OIjAXbGNY4sBK8PApgwG8zzJ+YEnqjtH6YntCU2MDEqGWAd8r6f8d9W
Ssn/V7e5JohRK6FXUu+af4mhSJXK0r3xxTp9YRX3/vQ2SjMjY8Y3reOs7R2dRtT5
dpq9ETkZHfoM2a7KJkR+Gu9L3Ay9hmRb+C2rNaT1D6DXz2diBgoYaQOx/nY939Ez
ytEU4lbFbOpQdZw3YyVHeqXJjyiW0fWl8V2j1HwlHiTPRhK38svl442vlbN9Um6E
SKAPQgc6zxmknpc01qH4TRVLVdnWhOZRvm7P4uCda2VTC71mgtmmauAUf68Dq4Hd
l41/c0Q+GTLp1YSkC6qP3hBEEJ9x4tWO0T2XwaashNGak5gcc1afp3K9PjS+Td8Z
Wk7W0kxTXLv++DUjRU8O6mCEWaCrrxLKgtWceal8Xa2DxK9SrcxYFqj0FKKGOUW1
8y3emwjnjJPNaeeFDMynSbQ5uoxfQnHsDimBJKamj7jawgDkHXxTIsPff9us7V6r
+bY9Y9v4gwTOquxNlnpnF4iw4yBFSBaV72k6wHnROI/9wvU6b5aup7+ioCc9xIee
T+iwMnXeX3hTyYLjh5BbYa6IxBHdRMw3eXxVvTIz7//7sTjIgR36iOTaq186KxEO
TTiiJZhuROOuPlQC18A3EpH0Ne27jBGe7svHHMvjKf9+yqXdfvpgR5oGDZ/X/Cam
TxrPSmh4tlUn/nL2/iU4gLf5D8+GgRTGxuHVoaWr8IRvKexGSCQMQ13l3NJMXRLH
IwCfBmWGaih+SC0HsbYQSP7LEV6FsKl7eNN0U/hWGz79PfnjdfmS9gc3D4syO0s6
FGkO30RpOZ0FvSmmFMrjOfG4v9p5ALjKtHa63fCdCLT2juT9T1qHZlIYExo2GCTv
PyWiPK26wj9OYZrtPGBcs437WD6GX8AvI22DCi0RC/8tBy08LQ+p12CzQOprve2U
r0WXEZMGmWk65wA2OJhEor4NbZqlQu/nkQkLBCeNDOkbejBUtcGyqharBHizKDPs
tqzmN+3jBY+OfLtyF1oL6V2ZdfeGpByn+cb1sszEjDgCgMdvP8AgDBm3nyYIAh27
dJlRCK4Lni7lRlMPdpBfIpy6mrSeN5n5Hjf2vmEc4DKVvzpZMp7DDziKHjpYNYJS
uIWH4XKUIrFx6U8yvF39lLZEwylIdRN/dVR9Sqc2Ggk+DNC7ms5wQW6wgJudbaT8
gIHVLc/f8XFBeOGQGGzJZmob5F4OHKzNqiWyIhwp4+u1PSI5tDDlWqhdsNOXXn5U
BDz9nkR+X6hMJkbzp450ooyjXYEE5vRAmp9hZEQsfXtnbnMEl+F8mJymf0C9WLfm
cRh6D8ezgjs97C2k1RXiPArmrQ2ncEs98p2J9h4vO+nuKRmBcLI19rDPXjkavLH8
rgu6MluJh+hCUBOakPqsd+FpaubX5IdsS9a8g9jxpupYzkfziyk1dictkcZ7tU4P
Cvht183R/P7fl8AnnJTptVJYOqw8zASjelpBSBteOvDlFDmDSV3dt7NVT8d71avx
gAkCvkK1aGXSlSt4K8HSvWVR0liyP9hMbj4sCNAbOSAAE32cnkASiCLsDout7FzA
S6AhJiO5Ae1pNAbwCrHyXG9vlIJTAFCi4yCuHuTaIYhLm19KaABFae9IwMGJHRrI
ENjP8SlghqOMnpC3E2l4lsAC39CJJsf68bHN3aLRofnRz0XSz55SK4bRX1bdJ5Gv
Z5ZqX/BMKCLNM9gvUJWjBWiKZpdd/8839yQ+5MbRy/NKP9gmbKi7cyS75hcpyApA
W3KcufNSmkLWkFJqZ3j9m69snLJcnKH2ICJy8efNw0tbcOhajSZcmbcrHAsS04OX
xBkMyKgqnjuPyIIVb40+MN1vVrz13eY4p2+9JLWAOvoH/QERIk7/nKgmHOtzguSe
+oylrgZozO4P6pLIV0jwOkSADsmA328g7K448Wn12TQDTSimVBGlxSSdRtaEVXvF
XBFNnjeZnE7izTy/sapE3sxvMgASnKSzQviq8vrJV1yDYWGeaxAcIEFDgPtNackC
6wpYSt18G3FBOs/ThRYmtlBSLtPOgdI3akKRsj48K1ti/NyKqvMYLoZiQAONBINs
VGDzoj3UrbQqtRPIFDd3JPxz3/PakzbiblJgajJsabhhlgTmYkcdiRAuqNuNKCCv
Vy9DX96qpovYnjedtUUzEkNLenjs3nQLPgFtwUIz1oJ6H8k6b0Vk5TegjrOlrPs2
jhbgl987wcj6NlxzKBx+P8+aBkRiN63jz3Z84mI+kEfg1l8ygJbBmgUia/qcXij0
XzitWiVX9B1ZtFJWtmfjwauOUsCqLHIS0fNB8sP2Ltqk3DTN4z7gOQtoPzrLejcY
jZNpKdzLpqrqoQ+j1X8OeXepgHoNhSi7D/aHq/sX0AzSKiHOhAxmCn9D9hbhLMjQ
7mLlMObgPPvdfcnrfNuZVPdy951fd+vO/RZuqZNrx9D7Pl4PyxCzMkkSwueL84aP
ZPv7UgV2AxtsShkE0wOzEusGN7XqUPZg3lhRS25gzf5KIM2Dyx0dIgwZaw2ScvIB
IXrxAZirUcpEEjtDaa9X9/unKPIIGftmA1YBn6jQbccsjwPk2vH+xjfTCJ/CRTaH
ViEVFtpxMgExYtNTqd3nIz+qRVCC3Q9authtuO4Dp/0nji1iSEPNJI55XwuziVwV
6XztPYA2FJqh4LdLfi9+jDNNxdFL5QE1Et8wY1CoSwmshfiOme/ljyN2/v6ZLNge
ilesWBllNd5Xa2Qpfk1SfCRC+uuiwv39/ZdYSIm0blPGEuNZv0fvi+SgvncEI/yV
EaWovR1g+QmJajyAglaNT/J1t8Ppq6Ng4Ve3AmgdK0W7kKFR4ORNhiVQH4gWvTOZ
fRic65xWQCojFLRIgbrZcM91VTfWs7hNgcP87R6gy8RS3UT7RatvXh/+d8wEdzCY
3sEWVLW11YuTLi+2d8NzpsntHmUZXB7GdWNh29OCqYsbAlwkDNMgziAx93cFKV4z
YGH17W8vj8T/j65N9Qt3p7YSsAJAyfZwWE8V5Pc6RkUQ2efkZ8Ghj5IntD+uZQws
k09ReemiHL0ezcEzIrRI7+2Th/Eo6FjBnPtPFn20R8h8yAkTDX90kduY9lzqkiJR
6qd94eZk7q2yj+K8qWqBL+Ive33E22/zPed+YhYhYvp94ZyRkCZdHdFHihapBt0K
xbu/9qGssUl44YUImfSCQhxBEtM4w06zxvy6xghZPZI1z/UBPapixw7z5wBgMP4G
7GaNrH6X3Ul4A38IBFSCVK+assXK0JipFE2lloxgILiegT4cXL883jRE8rIMkQ7l
PUINYslTe9wiAtxPPT2Ef7L/VUEs2Ou1PE5JjheUogZN1dif/0nSn9Y/Y2zcmtUO
Btug4nWtY9TvhZdvvxpKeNnvOc67Mz5Gs3pqnsVOnz5l37Cv2MK6loTSKZYdFYSh
mJRFPQJ3hbONZl4MNKR2ZjIdcD/txBtLpqnZOXRkJ7chFytIKreUU8sUkkQxscAE
QdwtTPopEvXeDzPF1CQKM/LPsGReccdJXogxLEvsD/Wa+xKtE1ShSzA0zmC9uCHL
LY7LYnV+9rB0O1lOwWa2mSXUsJs46YeCol4+9GVusA+vHscsA26D37znViU4phAj
LhJujxnFJl4scodlLoENa4Ug1dfrudJvlN1sgcxCMmsbZKuEVx2Dce4FcNrNcsKY
mQkepjERJdWpKTAYGHbKh+y9hZ/rSPrKQ8d3t+v07Ve87MY0oJTrd/oeALfzuZ8t
vzK1P81ixGrq/8WnAidnRFypXqidlXJObW0Pm5ozBv195X2XGYPpw0t6769N1GRx
DTqyZrpFlosb2gs7oF5HliNaB/dYBP8HTtXTQVm4JbsQBHAr3xQMRgO4SAMil6RG
YFSRBMLJT+0EbnOE5vPneZb6fb5pWxp0z+Y/3zluZvGx7jlirI8iS18DGVsGMkiz
HUUwyy/RqTR8wbGkf1hVWC16rXH64FRwqHoif/u1pRFICgskPDf/bpNwlrpxsuxV
F/nkBBKlX2VNs9OF1+7JYztl4SoeSaUYiQKW9ervQW4TkgJpgXX+isaehUbL1lk/
S7n5DGQxlT46Y9U1XQgraEFpg5R2qWRaEmDXUSjLU4DZ6/em7ynQi6WUJfY5SWbi
NpJXERuXOsyoQsMbNQbvpEkQJqgzlsDn4AZ1QYEbzZSLxmIsblzy4aL/3HI/tafh
XancOHiqUZdwPgJ4p6TigFPmN3jXaIwNQINmsyTZeveI5xt5kvM8RrUgqC++01vV
Ek+p4anVpYoBOUxZp+MGasSuSA0uuLY/Zxga/3uIBSm8aICz7kXFUkq7YEvKAI9C
qcfS2qlBwsyJ8Dw2deoUzp58qPEkDCfkmZJpyi8DHjqDrBlKp+SgAftTkQn+EQe8
E93VjoSDJ7tpERew9ZZSbuwkOU3jb3CYaEDqFYYCHYFaQBSYei6+Cch2Oa1dAU4j
6uOzT2dgSAmvFl2pCKrNajhFclj4m+O+erXqcLLqB/8HxujdCvd777XM9yVfCqqB
zlYQv09OrBJPZNKkhjxN5TRFZOfyLdSjas89Zs/y7R0ukxQZDIjnJ3cTT8ZfECgR
xbJzVsYmmloKay1A6gINzX2WZ1F3nqskf3Ka6hbH9gfEK+MXguU4nTnzTGvLvHN7
ih2ItuZqMqEGle7sDemBuEp1nkjcM7iBh31DORA5oug5My6KKaykTrTv/E0R0J/Z
44qgPQ2/8k16i7JZqdEWwYWY73s0wDZLU4K//gdV/9ETjLn2rwActjMTeouYCUME
WFil4wN8LZLjdinU39UfvQb2aLodMpySda8XawqqHrbSKghqOqobvB2hhi5TG1j+
5WUtx+634Bv0WY3i4s5v/nf5MRnUrryUADZBRR/ZzUKq9sTlz41H4NSzGKosI7aF
dxepBnRS2UylAX2RyCWY5Tx6enyP+fi+bZXh9+BRgCoa1M2xoMOErRSuvH+2+7wD
OS/17u7bG3LvlN5TCGLl6FvPgwOSDBQ6ygf9I90UktNllXZGeb9svE998ge49RGn
Z5zMOXxgkhHc88YQTMwuGwwXm5Ch6xKpPQuXW/4bDWICW5eiGWEaT226eTEiAl0V
Ll67m+dMLDjE0IRZuJKXZ0XVjocaTaCxl8k5h516oZxP5q5M82q35VrClJfxZ7O6
8rcdDQ/k9kdSc3UGSoD268y/cpFa4D4iTDe7PDH0p8ks4VCTctFkHRVkXgDvjWQI
5o6oSAXNIobKYuUFk2sReKaer4PdEoQhIWyXJsUTnAOsUb83MZ4z+wuBn/emTvu/
s+oFoqkLO/ZncvQSpYUxLIpO6ezvQOA1XWapga9+bOiQh4ED83im2JNUdRDubtRK
pHqzmEipSdqJhRrAL5pDR44USSWvWmW/0YTgCFNUkK5MvOaDIJMyK3lYPg0yS/fX
veu0Y58Q1qn9vMNrRJSypmlr302m2wFjlyVMI3b7hyiOJ8foMQ7QTxE4oxPwqWDG
+VWcggMQCYZnlR/Rxs9qlIVkblSVd5P2/RMyC3Jt2z7RUPzeF7eLx57ldZsWMqhC
bPvJCaci5kasApo3x+nfFtNQKsZ1Odaxn7M4xGkl1Q86jwmqvFW2/PgUW5ts0LpC
0rcOQLz40OzUEHFrCSZBB5scPr6JtYp7+nTP1hTmNQgsUekRtRs7PjxwkKePLLlD
lgrP4fMs7UpO5BLwctCeVA0gp+qkZOU6c9XUBL+g4kb5aet9CZoAJStAG6FaDSZA
J1lT45c5ppbWvAbt0CHiiqr+Q2gMoeoyDn6nAQ/BKr7GZyBJKxqHecyng7S5IAiw
s3g7pNSy93TEIfsTMH35iEnze3uE2JfO2gPJXnlGjBXRrhJitX/zjj+LHQZ6CktC
3rN/BEZhwAbJfijaYUY+JxmaGYgYjrypcg5fIunWlntSri1gamVsFOJGhh1yqdkg
l5iFhdgFjkbjZJdGMIZ+4N7/ndJhsbKW1Iglohjus+H4nvW1VkH7LjqYg5dtR10f
U6tQMvhdxs6sqhcurB4aNS8YuUCaSWHGzdvYoZxfuKHXmzv1GaAZc+vVO58zFv87
eYOl6ECL2bQYqbi7wqasdwt7X1gHbqjUSu8hw+taiQSsY7pabTqoGqrZJEs04+5g
VuxM93ORXcRkFzWfcANpLaLtb89BortXQMIr0X8vo4LT7y53xzxhNMRPAt4oVGZy
r1Wtt/EtZLn4C3u8HYGotO68EeZqC5JrlY6UjnsedP4n5IzaqR2HllHKCMOi9t/b
fNGQxncm4GzuSbFxt6MYpl+X6hM4BZAbBuhUDtnYisR+uxywSjVN1TmpEfK2b4Zq
/KORfHhV/FkBB3bxBnWogsXKGV7lVfe+k0Lc1yWxlzkwg8p1qQR9aONSa8z25JiR
Bk0MMoGqo7JROq603c3nMYAKncsoSfgnufEcodmetCu4My7gZB2h84T57u3Ak1ad
7aOguQb3ChDD/ZIePBaccgIXykvM0wP1FzjPuD/NGm2YqbQDrd799FD9Pc7mhQsm
SiprKZDs0ZudLtNzxVXg15PdS9q5hhTfyM+3ePM3+IA+u11ZuVpfgcWtS7bsWuSS
VsZ+yGGst7kuK3Va4HG17a0+MjnLHw0TlSj8mObjqPxg0otWo9LsMWZabg+9d6aD
W0AFoQMkA8REMV5jfTV5y4Kd00Hu3+FRt+l0tqm0msKGrtRD3hbH5JnPbvjw15xx
xj/E+kZgiRqZ5J+qFmPnj66s/ZL8fYkZnyMg/I+iR/t61CdS0IA5oxv3k7VBghtA
kZ/nifcM2Nu187q1Y3zTpmorpb5J/P26+Mt02WyU/92eoRfIVY7+brruUuskQ66u
3hLXwwowmoSAsMwfugd5Uid2GNQWe3MxjWNzAl2MnvHaSdHueAAs5RRzPIDi5JYX
wgaY8b8q4cC88/6wc672eilg4qJEYKMSqIuCUdbBtAIG2nseMnRI2+RnyU/LljCU
+h8Slt/Mbjl4eeerFtW5ek1QIBA16ynmYp3aSmEWLq/+iNpSK450P6WnUHLrbG52
M2C5zLvKkCCS+xEo+kYccluparoz1PALppf1iLgSQp6RzDs1epYBygoKDe2jEkt3
sxUNTDSun3lfTiQB508xwHpnrWEJqa/+oV+y0qt8BNIaJA7Lz0lmM6c/J2fAn+ke
/iNrtdGjsewmBkU3zPw4ek+cBqyHkWB3rSc/7eXAAolT0gV6HUchaVWltgN0O5cF
RiTyMiP/pGt+BqrKMTA0SFtzHdbzWVIDVo5T7csIsURtJ7aRzmZz8oW+e+o2rWmn
jWLYjghdQ1ZLhM4qwdkO93dBo+NOv0ZakNLleij62splsOjAg4ktTxy+gFDfth7y
m4H46M9lj3mhEfLVrbTpmN0T5B1/DYuSsw7UVr2Bs4qjYdQTaXLF1/SI8oEjwzPS
ZJCYONntzYbW1w/OpV8EPqJ+xO4QvzcZfooOXeiSiI6u5w5U1sr34Hbw0SOI3A58
ALVZk/MYmk4NEXvmSt/3FMpsR0HjKJMRAeQO8fw8aOseTNhtJe+8ectyAKArr/Lv
qJ1XLK1qaRSu2+0WZNse7o/cziJjNRjxBcCdeO+Qr8r+cTlqyTRqAIeCz0S6/JRP
9g1CpIDipE1QKVzYjkdPUJ6x7P3djNHMzBTQBvlz8fq4HpvFI9N4hhp+YxAlsimV
aLyQ3b3eQGuk8URgecPmyp36c7BrUl09bvw9gNwf2NU5iYLMiLfNJo+Dv8N2wVjS
shpKdAjtQfTmdY23P8yGkXK8qqkB9qXhCuQ23cUvdWUdxmisgmzZkxz0s4tqG/IS
Oc8KnAy+DsKSmYG6Rp4rYCCslM0VGOpQryUkwyyqF5DUYHtOfDiWn872a+6Q70Lh
BG9Rm+SqTkvYnJZOttYGDnAvZl26Z0C4cZwnZsO9XuGGeUFuJNfgd+6aHOHRnD1U
2P2f2BMjChEyy4ClJis+TSUAWoe4Tm4VefQ1+7FMAM7W/pHGFVRlOZ9yQFZf5uQm
Xpq6JJQPhg/d32mCBislO9awx7MWKfRqDWJwT3qINWkXkfo9HqGuspnXTpjTq49t
kEuBKLP22JF5n1AkQmi/PedFEC2NLg5LMnzBSJUy0ga0C6Z1UK0kge2PeyhsNs/s
jmnEBXyH1oFjwA0h7Kd8G8VUznOfk8LKA0rGy8jSrSj4sSNxKh4cfS2uUTT2+qu9
JnEMVIiaI8zrpR+DBG//9vFU8yUZbEX6c7rFs2cjdIUzeeVrSPGSQweDL3BlucI9
Cu5kM54HktIstAsCrm1DXzE2/vQCCOM9yo77eBeK1/+e7BjAFwQzcXRDbaqYtiv8
I0Fm49kzAFBJNQsnDWIOuc3r7AV6/YKKeVcOPl1MtBOG8Muh65NCPETiYDNLeHNU
MY10SkgXx/JyiEr1LArWX5dcu3rMWk41zDKGuR4T+O6RaQrAKgxzc8695RCFaV+O
CPhbf6IgqWB2l9Yw6D9t0RBdm9lOix99SHy6lkoL1/uW3omr6Gc2XPZV6jLUQo42
ecO8Lvgd44ZStdjS+qGp+03RB1JC1OO5RtQpo51H/fG9mBR6mFTUL/hYB3scv6Gj
jfiikmZYSqjzN7TZYdqUKvQPKq+mfHPSq+xB2RIXtsy0gEqQevdMdmCsiQLXeawr
wVuyBYOoALVJr/RF/9i3Eq6YgDFn2fFnHma2UISEsXdGXGBxr6p/oxq8SMqAujbV
T6dBcakxTSkfLqIPyiNVVWC9IxP+KQaorHmpl/mlT0V343FAMlSzYtxMkcXKfBhP
RJ/shzrvnMexryuGoXUX03rZBWDCnkj8V/z3XKQ3Sp7pwQ9YOP/Qiq8z/BJoUh+u
xq5POtrIWxqwybsW+Qc/Ys5B4MYbBUerG16IT/bomcXwJOuUoGsPi5PDzcNp4z7X
bp5nDQkVfb2MgQQVHilURI51W+e4h30bcX0TjFCeOKX9E+9RWizavRZfjg2HiHQN
LgI3pP7i6eVdSkgm5qGyqX8mImEKBmsN2crUpUL3qf6ktZreDHj6Ms6CLAPHFl21
4xTH7sz3SwFBLDgbxFKnMsld+q0LpIFYk56B8ft1tRyQ1cbLtGvG3NqbmpdjsHBR
teGq1UeqkQlkZA2lF71fiqtkqpO7dFzjNqwJvQoG8P/EHZhBXX3Y/TG2SuBBoPth
IsvF96pF+M7x426huTFsUyts64VNdKHAhUs7LhaCrctuQO87wDyOZIYSIRrDsIij
I8oT367CSqgoiN8506HQtdott7xQOei9qDw2tthN4IXXylVcZFApB7SQLxk7sLHx
AwO6mMBV19FmnCKurioL7b3Ryxy7lhCVmDgfzNR2/g0k/aJz914VeGi3M/CqCmEj
8MecLc+22klaJ/JPsPEeJ+ZcpYTaGjbIm5YgFGFKMULzmO3mZ8U3lzm+OaWsGRzA
9GJflVlwnVQzmaT+yyAVrqjfVtDz0pbiMiSRlC73p1uV5jNJjxAUz6ChmSAtrsvC
eoUd2VDm1SQ38WLbxcwSynEDAnx6KKtKHDpmx4DVG6GwmataNl6X2pfHrh051w/i
bATHsXOixmreEQkVnYcOgFkYZCZDR23QtY+0f2k8TiyjdWSlQge6NnJBSlxKdeM8
4xWbEl/zRB60L0eyUbiR6coni4aEFCKxg+7QVMbqc3zEiNNPROJSEo++pDjg4Chu
Jct0Kmf7LlK/46Y927QQgB5mVEz3EQVWdC2GFGVxwuNVnTJx8m6IuNqGP2sJ9Ugp
qRE9gXWvL6PCXys1JxVjBKWQRyHTJ+aXyWTJ5+tJ4ExYAuoEuw7W692Ij/yI1GCc
SYCY2nqzBtTC+OS2toemn5uzRFm555p3HWmSPqDDec2Aw7RfrsPuxj5mqIZG/9HB
ee8+swiQkPZHUC627PNsri7JCC+dW1C1Nw01ceXwr355QQf8AyZfF35nWMfL3ROz
+zZvhiP6rB6OU1tuA1JVDKPCZKrOUWrk58mGwfZex9Zf0og7f5MAsdMzK0lf6HLM
vT/7H9LOirG+radrkQx8gasjfxPkIq1n+9gIufb3MqU7gQStl4mcMM6FcQRmW+XK
ZPiUCQPQhjMVVldDMZ2V4Igm1MtzRAoU/HZ4R3uQ4XsmL3Oa+Zm2210PNY2hJXXn
zTu0BrcRb2KOeUsYMm5DwIYCJkOGn56cENlIxRSg3spDNH0UEquh9GK3GH7kR0Ue
/S5hVC/QxEm5jhSsFxd2YxjIygMgkE7cx1OWjL9rFHAELTOzsEdqvkshdX570CDM
9DZyywLLGR6ElmcLHmRhAKUVxVi2Rb2gfZdtrx456P55zxDZfhwAfgJ0c/fInflp
CmHSOGFH2Uw5rAilLJHoi1DTP/qVBz07avQKEowxkXwjpQvjIpS2U/yBRIvLddzL
rQt3yOgOHl43N07hsni8y9BSa1D3kmDwGlyU9jGWGX0mfeVpbRqrh0LCDJDHZJTi
S0GWmXNCQU1fo88mJIlOzV1wCSX4QyYkv2fQJpV4pCI/vRWtPcrAXWQiE+GrHKSJ
fwJcSBi5G9HPE8NsxZboj860WgicZ2XApf4dqqwo3Z/eE/nFGi8NWCQQ2/6p8BbV
YnanV/yiD4T0hfU4JgVSW1MNPRSqXr/kpVDyBIcDmQ71ge3LAFPpdmbb2sAtRZM4
ViOwTGzDFwEPldwLHMLTyI6sKcn0UcgHsyTGO11RbuofoSjiueT4kHVLenocRgEe
QFgOGaMMUqcfrsjg2NbbtHm0SaGsCsa9X+jhy6/SolcfYeCmX0clQivR4MLVPdwz
5xDXTZkFNAVB92G0CW5Aidk3jiUUT5vQxFvopX+PnIzv4ZFE7oWuBAKe7GmbFFdA
MUv/j8yjqbQgtp6PgRzFqV6Lj4JYyv0kOl2bwtfFgrUYXxOzcycDOP5xJB9YIptu
CVMqQztJCJ2447MSOQ0ex5qKjAa0vb4QQ9F4NSOXpJGfbPKGZnpRj38o6ap21QHL
ZoWsy5tGF2RWB6+PCp+XgwXUQnE6zdX6PKid+AwVJENFdbfdEJrbftzmZGPSR08t
l5lhUvU+ebqR6Fkd7CefsVCUDyw/hGS1OOyxDkUNPS7Zhc5o0JPd+zQWqV+ZE2mI
415h2Xd62q18JD5AVoEoYW9y3uc1RiW/cVhNfpZ1kMxr5RFjk99ZQPiJC0KZlSnT
8wf8GSg47wDhkCJasu9Ceb1z8KssfqLbnvW6Bqqbl/U8GBb3E7Oj3qI4kJKt7VaD
biPcefJDWxNTekZZ93N0v2X9717QmYY4/l1JB2BegFsPcNRe6BZuE6Xini64mHRs
k8nSkznG9mrWOl3IFdXOKClm2waCqIrttiNeE9p0R4zoZb1HgSzCeuVokbaFNZwx
BFmt4w5ptSrZlGyhc+oz7804acFNApnWBEffTT6N65QLxT5lqDWET09LVI+yX4q3
9qox4SY9B1JJOfvFgVZNeVVu5L+Vn+tTrXAjWnCT45EVAsZKJoZlWTZsGcNEdI/4
YsNevtRZLjXsaniQ+hkxB2QWInZ2tTRsuk1FKGl+nNUUrITEjj/Zqz1qp4o/3Ouf
7mYEYgOkqIdo16BARVYRPaqE9YKxpHJ4TiTQjFUWrzCtW+hzrObz2u97WFmetjy4
iwchn1+udxEonqZQNc8mlRW+45mIQ+NqjizBKZU//nT3Pv/V0+XaD95gAHGMCjGj
zGk1sduiD2yxB+LaP/wfuZu1Lu6ILxA1ub4sHwSe4F+kfLg4hGrQeckE2ks/u2CQ
Z1yVD+dYVDjJw9R/pE3u7YyIkZKEJK4LQNVRRoQP/sjt7ksVnG2vcvAtjCzsQxtL
pVWjisYJ8JNesdDq9dku6HOsA4d8IGsp70EeS+teBAHiLx6iekwLVuXE5CqhgY6k
2kOi0bKudLHoxDO4OxVVzqJ6SPy/GRRGuUOMuKbdR3GSCyq/EAQ4Mhp8YGIVaO1I
CIyOO1NqG6krOFT/RMlHCx0UrChEXhS55+i+ZBwAqbKkUvJ8S0oWua71Ke+j6vm3
zNVNO1kv25ih5HarOa1oTjans/wphKWEh9ueiQ5ViW6u0zeMcpbdmvuXV5MbIHuL
Zla/ZBHaBo7KiqrmIL9DJz/qCmzUqUM+2BhxYYtHUmCz/ZctlE0odWAXQeqaBTh2
Hd3387zdZuDUGuFddd6blqy819BTzxXLCXWxTcQMUD+FPDU3smYddgEqiGUTbAPZ
fRgTx5rrshIVGqEZ7ZLsqfCc/5sneok53omVR8HyAQEVAnjMqINMnLs46u1Cz/iB
CSGBZf3Kh08Ir5lkq4i11GouCNuh1nby2fbiNKaJqa8VTNq5+gmme8vGNyVi53h+
xWPh827/wHdAfkVxeH9cDRrvZd0QZ3TaFG5/WJi52HT7f7VcWS8jZWkZs6JW14Yf
eC1cyUWX2YoUfeK5vuEaM7PjxTm4v8nhnigboN4p6vq27IZ7PxjdcQwf64YmOzry
n70JMEW5Vt4OcHF9teovNWFuNp29PPAEm96/2BLLvejFAKMj9bs7amx5rsKQTMrW
pZeAvFm/lPXxCFwnnuyFrjlOmzeRg7iTmEhO1SbvAAiUpCfvtwsLkQtexRQXdjRb
ZTptwnCeERGofaTsg7wiuyno9w39VMWwTbkQCKIuPDQCQhbiLHrv7P0qC5uMI+jf
8KlLm17BbiRPBy523/kkvJV/is8FLY5QNikAKvCCGO27XFUsq5IL8/hVspIvlRNL
kZfwPSdfXBINjE2yW21TH4GROqVFid0W+/8b6U3ioKR+hBKgieGA6oFEQnoXcJhJ
qz5KHqFPTI0gunFjtFaoyiPFWryhxcsT/7DOLt9jSkj6L48nlnjBSqrP1eusWH0O
tYVJvd785LguYdRjwhyqVqs+5blnQniLnlT7G6bodRyBu3oPlCJ1Ek5aTXzYytjo
fO0WZVAnnIlFSv3bphdE36ecqIFm3K2VoWJJnsQOSTBjedHTnHq3DH8gOhAuMMLk
bsxFxk1ownTHxH7gJsAz6wanGIGSOQpEcnQhOvIkFC624GVpmqouBRaee+pZb2zz
X4lGt4f0HYIaNOj2qkHWkMutdqq7dg9HYv5y794eJ/+YMWrbbvxgL4hh9LeHTED0
t2dsrpjgxwuMZm62TNq+OSefa/U2HfCeoHlW/dUw1+InrycFtCKXnQ3c6CuQJf/H
oK8+k8omL/os/ZFgFR5+veThPTevHqDvw+/BOGq5NtyeKwRXgWjp0A3D8ClCGCSS
+7K5CBYnVSytWu1wS9G0gRPRIIeBKkhiZe1i699F2hbn0J+zarTlTvwEP8PoZdrA
JUy00zLrz0tYZOkpgQfozudN1HTU6CcdUFtnhvGs+WzQ19kRsRvWkHNIbN9MYxVe
s1y1I7Txr6lqJrWocH48LkLAaIAwhUlg861gX/a70BHyUEYqFNhaof5zvcBidraT
IgtM+59YI3x7GjSHOjIWA2nX6IHfL/jk+aASyhvFBYnstmty3u2BQZrn7NR8KVt9
KZ3syQfNqdjnFzvVjiQCeYgVci5mGWAwBDbITvRhU4xgak2JfN/mranVYHeBISya
NOtE/F+WSs7Srs0YrDDCSEI0mIbGuzIbUzXmikBa4Pqab5YW1LDWYGYfch7FYvcC
fkiSYzfVucb5s2nGsOjcp2lwj11Mu/bXjq/ssVdq/MKQ61x0/yFglxd51FVTBruc
lFlWTYSpbNTmQLL7uLdtkAsIe0noXSUBxINQML1IhtmcwZtMXb+HkOOGMDi0Z9mv
oy/odch87xNq3/E5IRFgcKPMHcPRdPgF71Rt2Vpfk004OKk+3WwcrIIE46v8scXZ
CRtpnu++dCYRRCRDbFTOIsrkCfdgiLIywLcfmLD95g5IP+fek22DDHPT1PdHwJLO
+Rv77d0CeeNVDN06bFmVZ85ibIE2wtbEJ1P2kRNRPUP5tCY34q7rGCbBAv9NxZmj
KFHbaHIBEO+E2E5Jw+tyNII8IUvBqHaBEt6vx2TJmHa3qgug7yOk1uyFGc02z7uN
DZmcKXGAJ9oGgUFp1U1yXXxW+PzPBnfeV5qJV/nOpMHEsBUFGatzjN4PvafaYXo/
EgNb38HAdjNlp1J4m8HgCyVBdBuoK16D62GxSLOUF6w3nDyazPRPafWOC09IueWL
qHbsHpHtFwgUBebpee/D8LndVU8tyyT6Rq+pucOB0B50TbtXOYOC4b0iWCKDRS27
ptFJyuXkcGKdj+/m4qYI/0shFAMYO2SVfkkTPviGX8pXSBsbDHvzZXL7i3bWHdLz
lKKl0DCbJ7zpbN14X9t5Ff3viVTk69gdDYUtYWE/UI/vMkZmkPKCKktVJ4KvzeJ8
xQMT7H9mXrqQtIh+x1ItdwS9eKDIJWzg6hlyUD6C30RpvzbXQiW8Q/kcveaoF14o
s2Zd+tRBHEiVs1Oqn4hw0TaMx05Yov/gy/gVfnR2q7Lwm/AcIO6QzTCOP8RFRv+B
y6Phsb+tcKEPjMhC5cVyzEW3+FAqxWbNQXkFL7TOks6W8Fat2r5vWZRQjtP99kd/
Vo/eRakSgcIVfR5sbPYpDgX//Fail4l11xda0mLeYtwz2cisxIftCbnJ6ZLlf08J
vMpcpkOisrnKBF6+T1HTnRCZvF77PHeZl2OUzrq3znTyGftdZsjbvaK6yVxa9Z2J
1HihUXXTNcA6BkXakZKgRnkPobFib+/akZGP3GqaZ3iDNmsZn+7U8qV6FNBG/k37
W7e6ai7ASMr3rzwvmOFnOWN/aHtQSdfq487o+BamI9jB6N+/ve4IYtDa2ytUbxAq
zLCczT+POxWZPgILOiIwAAtn7a1kKM1GFnmqmv2sh1S68D6BknJMGtN1Gmp+PhQm
9HtTLHoXiRG8Ooz5uNY57YkrRWS25AA5auh3Dq91F6UJkwe76tGnp/DEbf72qMt2
+v+MD2nEzp7xbJNuRhDNqvjwURf3w7XCLDVnBwdYWn7U9XMEX1lrd8ftjBNZOtc5
QI9BbLCdL7HNHOcH5PkmnTpW+HWKvZH7ijUdXoCxrBD163MvA76UdF0NLiSgv0MY
WyDtF6kbpQWRPWoCVXX0idzDIp4Rol5+1TtTmXIVnbDWJgUBxOBP2cV9dJLbcZzD
1Qw3oTz7khbhMjgms0eWVLOrZbId6FIWsmQsVqbj+q64pJ0ntoCQ2TZl2hGRgoJr
dPZ3R1qEQm1SzzMSh5UZzS4LN8Om12xSXDLxr0/Bn4aqFfZ5verdWYtMvdG1OApC
/566bRsqi0vWINWmiRvB9qPA6/XcHEaYyyE3AhMHqtnzkY3JMK6ahCXOOqCU0Ke5
iXwjQVn9qfI9fe7VGXFd34kpkf4NnTmVEGzdHTHb/7PLgrKkO4tC7Cf5cflefALD
3eu+L0kksAMcTvr0BA15uFn+ZJ46XmtKwWBwIYwKsM+Gx1juvGiljM3FEjTTvlh9
sIYohdzpy98z9V8h1qkp8lY6o0TOk6FO2XHyIfHomq3I2cZyqgh+OR4MIKMERaNv
LPozj0EX3yQlBMKqed2UgXMLWnmAFE2i5g4YFXYUKd3QYL7STra0SmG/1WAP61cc
YTQuYB2HJqdv07pWubL6KBvbTfZstTWxkK+evwQldn29oTvyTafG4bfrm5bf9rSD
Jd1eYsj1Fkb2zhKFfcEIZSnPwXJMunIu21STqnkYYJQm2WXGCku+MZuHxRthOKaT
W//6zNk/nEAC8ZFuEtc2O+QRvIWfnl4m3wXPJ08yepy8XXO+8lZTCnRjSZ6j5Oc+
+/K6efLf+vsRAfk4o9ihVPijhH2xdeLzPBtso9+VzvJkhOnlMbv7JsntmGQoSvTh
bdsEKKaOuXmz3r3x2jfQ9Mpie+VtaclI7OBQqOXBG5wSzrcgFKqqr0HBkbAZYKk3
cXuRngN1nrMYENbNsIUKDeywnHT0rseQUqH/RKea4k3fy7pvDjK6PvswmQI6y5Oa
bD3g00FqLuCiA9QKT8murDx3e09cpOCBx6xi+juC1srsvCFrWS2EgDb8FMe4J3e0
vlJkWE7nhMrJBy5CilKZPEjTfFUBBKKwj1p6r3DWpgO4ULW9nLje/Lyz6xkWH2zx
gIDvC252WUQCRgfMSyC/XHIdb/9Jjc2x3Lu4ZoxlnoxC9j0S19aqLqzKEseZuJYj
Ax9qQpmHa8IuoSXmAhWa8EpCgb0yneybpxMw/1cWVamGDv0osWWLAOn1OOt7TV/R
FHYUoEKi5m4Fg08XaA+n2XSlQB1SXlui8KVcrO05amptLv3tRKNneFzI0lNuX1T8
rK+6Yh8cG3j7pFBHQBECssleV/hTo3KBerhoM1KmO0b7wtXJpBxKBxIlhpAEgoS6
GRTV0y+wdJ+3DMaKYK3Cs5LBtDk2CMjCR7zqTZqt/fWMo6uuwdUMi3fh2kkYTsL9
2311APZxeoFV5iTR0Z5zIXHA7YeudMlBiG9lLBsq4Ty97g8/1D2oBEgXwTewQ0iB
vNDjiKOjGCSmMhBQJWqlZZqmWEVpCOIMJFnlbF2SujZxAPPy21xB3Thowap4y9xW
0asH2tHNHZ6Acxe4AVM/8eievJqiEHhUGdSzKqN6V6Xfnjr/6ntNjtIb5KShlH22
kPH4MdnFKExFjY/FlLvV4C+ib/v+O10QJuxI4mvSfAfMghMP+Iujsva9AeP711x6
+4QFyrOJQfMTsJCmRcEGKdfYKTbOJ2ZTdVRHxHDAY1gi+xXQ/chlQK6by1Yj9q/L
K28R78v0eQVj6T93nfVU+olGpFIuLoweAdbV2OtPKVz40jlHaStXT799IaGqA8bo
uEyYQpCOqqSkrEjfcbsHwm0ijRNMcnST+sBGg46W56PavkwIYMXcD7u1Q2Q4uRll
K3qzaqqnc/NHuzCnwo29itQF36X48PM88yLrfY1MRzdq+i/KAAvTLnTPs+5co8a6
V92bTbdP81xRarEnWsFTsweya6O0kiIlHXOhJktNLt3HmxA8OlvpNqjiJmUP8zsD
qBk+Qa9nFz2lOlHw/piIkGiTAU9ftPyg1klSQIJYZkY2KAkORWI1bRwvalyrzuJO
xyFAdhu73qx1nuGx5g2wtid9US0JnIeOIfk48HqzQE4839H0Bo7HrcWxy8wmkr1R
ukvIeUWa60udPa0K9Wp79xY9y0kNyHv40Jmfk13AFw+4D0mvi4o3xS1S68NdmOXn
XeehgsgOeb6wK+ewu1SmDYF5Cphclo5qEsmvgHyNuIqDNbdCA/uj9ROqSrJBtyMj
xp9JXepi2uPUa2q9057rRHUPHv3FCBlzq741PpjIBENMkfHwkFb+dQ8FlohHTRxZ
oULauykXo0hPNwhKhwVUDCLuQomuOI+r3Am9MZaqR6zxS4qxaib3bVbmri5MXssH
9zK7GBsKxoscY5GgnavLZV7ZyriHSltG9tdpWxAsPB6VgTohVqs/CfVwe9qmatL6
VRO2WkN9HIip9p5ZWuzw0xMsm3vXFLBdP7oeAYmpi6ocWV+u+NWIMafS0FHAxuYz
WKmrdqHuh+4XT3w0/y4SQrMu8ZBW4ol6UgOqY+ngxo9P2wRLlwTB8kNyHh58Hr11
twgSmodgK7U/jOgeNX6W6QdnzsBxzjowQKc84PvamY3g0ZJlrCP8mZfDxi70M9bp
nOY5bTf3oYR/WXZZOs53eSHKq4MCzBhL17JRlxkj2oeGsHUlR77ECF8KO0kL6C4Q
Ze1peFBJEg2vTeyuihGzmmfTcdiHaf3txjm9DJQW6at1qiQXd2kTKvAjN+kKxquJ
Yn94Mu693HvlivrtgwPQP0iL1z5v5qSwlplIjXL748Hv61A0dBC3ivapgBC4nVTG
WgMmlnFBLcAiHJu8kvqMLfDEZ0Hjnk5tt6MngXUuHGEokSvaC2cF8bN1eEpod8Pm
DYpOzjxhTw9zoXSlOWi1bVaNcv5Z9aQBQ8C+f3pknLfH/5U9Kh5yHxb7VCPB1Mvw
5UNMoVuMNxY50O/5GeoRqDnQPDzuV0rcel9zh5J+uT7HYhYQPgVgRVDtICzUPKLN
g0OUNrFQX5UTCMKIFxZmZHtP7FdexBorR6q/NvtIuj6WyiVjP2QcDrV/RnBmCnwj
WsiOtzJsa235Kx1GxGmcwczl55e0syrJzGyxAZ9/6HM6kOjHgg0n58+DzS2EjAO+
OQyyUc0Ofpkj5oxKj4Qj9ZHd7z1rS8FNYJpLG4JGK8XfCUhkhoCwI4H9ae4SpqM+
uwQjhtXNe9+cEpB9YxsiD24wFHaGce6IsoRUbaYGfyODzDhLnWVzfuYKJGCA1LVy
eDy1oSH/W8bOKiGO2fIFTN6+jAcfcbxIW9vc5XX8z64pxVh0ISDn75yQ2twEdZEU
CNi+sY91ThYdoJz7MU8t5BuP9TAxsEwxgJoFA15Onqhubi2/ZSmZX9b/5ffX3p+U
LoEqzzpuOVtLkWkMoTtk1I9YKnW4NPSg9VQPljUuvBGUgp38O9Xyh96XcdMsDcQ0
NDkcRWVHKMnCOvWBVMLJSjmhrxJZM4CcPNUYvgd5zNfd/hsbra+JjURepSgqUDQj
9szbI4v3Wc3NDM2L7vgpo5FQ0Ud4tIca+rI0wZc/oPCs8Yu3y+8XFzK/Mweuvkja
/BrfIZoxfgn4I3pF5IJnFDwVHZ/cskGVazV/qZ7NzAYomaxvxdPT7Uz6/DhI+r53
sLM3Oo4WN2b+7oPW4/8/6qVKaFipAhdOcZvQ3sOimPZov3xarTcwMdpyhraGyWD+
QH+Rz43BVJsoOQKMYLScVFcjdVbVXTjoiHc5+wUIKGgPErd1t5k9eOGe6rCXYA/P
msEqtxfAsuN2uvTD+iJZxy63JbEhTS7YubWImP2XeoSpiTfHJ+3XqLiXEHGucmC5
miKRETAS4qn/U55DyN9u76TmGfjGPCcVIF3wwC49UoneOcGVL88Q0PGASLWeyTDS
lSlafwGeG5hZur2vaoSc3foJgPxcvQvwaJvb8pV2C9OQOuXUVQJZxkZK25b4jMim
paLgfhsaFXmqtbONmdGeH0rqIPnWdSnMp7rDOsYlfucfxo48Ge1DT4aKLiSr3pHF
D48zl3Zs1kTd4Tzm5U762mP91lVX56ufM/jaw3LAt94CoKEVDJuTTHe3gpLJYHIr
tBqvcbM5E4BVhcRvpvA/XInb12R2zuBHj1NV4ohT0jQCRFreoCtDSLunOOVbpkJ2
wVL2Rg+az8QVjyGPu75Sy8mwQoQM7MNS56h/amJ1L0H5+mrmP9N0ox3uvq1/eVU1
KPjA4/j4g4aDkRPP/clnoN3kL6JPLu7OL3/3AcBlDsBC1muYmwV+OjxvhUPWVFj8
8MGrfUVqq+9IpWdGjJmC11ywFp2B5gD4yfmEZKpxTxHNEG0lPhYszPEWtf+RrCs/
jsHOOPzLEPUfSYjfL4TW/9p2QohiMM+MpJbB7Y8gFSOCbCu6U/Nhn8+4fwtmCUgh
VCLe+D0/AdV9HxEVUoky8mCnYKBnOKfkRGyDAkfHqN7hbXAwI5xZ5iPqrp6tZgIP
Ls2CDUp7hH55QDWZIfeNSk2tlmQ5Jjg3x3jmLDbGXxoDj8BPTU9+hJs6kFthn237
omnXj5nfECTOM5L/O65Ock0NibArulZ6KeEre1Bjf0tEgCr1gm73mh8Z2vINW85r
S2kNgqvNJPp8D0E+az7ISpn1Y35t2mJCur0aZwbO9f9O1G/H5EyI3Uxqd1Z+B5L3
X+cHHhcWW48fXfG3S0Dl3dVXJFXiawNkwsa4g3hRot74xHsNDITGowA5L61fcLcA
5/fDs76LqDHIuwSZ6kt8s/arYFrpbykBK5lKKzAoxNtEizlQQWHwnTIyJM3eQYy9
lIQ+vr46zh9hwQZAdhGRA53ydpx6RKB5lylcQiDm5Dafh6q781CTCf/VtiLTxLiG
0kBGzCIGXN5K2wXzUmK0cCMjXtoCVeWqG0YnYKbKL4sQqnlvV8Hqr48siIMy7AJM
/CsNBTlbRo7QxvFFYcQiHI0HeYZAj4t/EibwKMzYTJbZ8WlAuuyNJI2oaAlnCw8E
8QuNQVcvory8SIr8O4nUy8u/hgpJVBXYrSsmH2Jo2Sh6kA6Vhgaf21ihaepdcrA1
jaCfcT/ziwTPzVn3ZXzOCmFBaDCUk26DK8mCk8HWCbIjllzEEcN7mEawp5yf/YBE
+LW6CHH/djPmDPVM1lrIqhx98+I6ucp29Qy54ukEuS8fajq4E4F7/rtUuhKjAwF4
r20cg73PKvl2l3F30mji7VVP0+UeAIyaYrnIf8QdFYoE2wnGexNuL5tl24sQwLdi
fpuEt3uRKJ4mOc7einAWicwSJwSjIjVe8HnXKPMY+5U4VetoIQUs3mcIVav6G8W8
v/TKCRB3clYIkvTR6gZFg/42yGy+52rrvKxbio+LBVcmmZM7ZX119d9gWkmb75wI
J3uZ2Xy9Q7xoo87lA/wISmVH9aSK0aX+yPSMuPdxj9b0sOuSMmTtjXxb/4T1ogtJ
TXGDkr6EYeLnvvTk0QaMf7EeZJv8bZiifrnz2aAr45BbS4hi5NVd4XXdKhiYSjL4
cJipUeruaQjr3+gxojH4FmiVvJVHH1tIRZb2sQgepkc6tss2Pq5fd8+d08jwRobN
+igc929TdnpvKxX0yJuQ9v0KJGHUnOeUQlGoKe6354YQ1aAsAfZ58cnP49gzDJbp
XWQ30R2AcUwP7zX+mSXpwwOx8bSMwc/Bcfon1jS+BBQXcvFHGjL2pReizrBZq5WE
SLFbeDl933qFJPffvH91F/lH1A7E4IFPk3dce6/7grqA5PaACV8aXRIUi4KBubgx
sJy/NKN1Ic/DUmYkPqqcU8JXMpInBljlesU6C6b1NPR5pSjKmi/SLJ7BVpFIqWSG
C50azsgLAz69QwnsQjzTsvE6H6p9B7NNubTKbTGAoosyN1dYkg8NVYNbrAu+AZOI
L5VTVJFK0uiDMl/YHeyTW+maabWLD5XgbaedFjInMdg5Djg3RCNOsVcz4V5zllMU
39ZdUTWXCz3F+2dRTUFw+rlh6yUA30H5wSt3ChKF8uUtjXrl+ntnGIbFJY+vNXbY
pJ7f9clPmqvdF3nLt4toUMfTMMrsed8UD/BGIPbM9c3Hx6Vuw+3SiiOlJpCXYTWi
zcITmySP/IEb2YX+Cuu+UZ/pNKUPLQLsyxjmYHp4OwQ5dB7ZEf1pN8Jqdw8MVVPD
0kKde2q0i6uKt12yZVAglrWT1Q2OvAvsHaprcDKkbd9Cf/etBb8on3mX+A8ZI/Hw
aB9rJR5cnFQjV9IZKKMmrG/Zz+wepc6bJMeLff1LyjnTGsbvzyS0NFW+ZTl2u38K
G4WpotThiFFisd4GEo1Nov9ombmV+fg9wgjVvikApTVE8W2TFrLhDZxOXUG+BOjW
stC0OJi/af+Uxa7rXYETUFZYnU1meqW9Ff71IBz+l/larz1oFcBEnaHQKpi/MYcF
HTBVoy+kJS7aGItWgVpfgSYqkTQE5O8r0p64mDBzt3gf5+DSDqbdYvXsqDjiAkCQ
VQzAduFPhjzyLqea+DlPeRnTWXqSv0E0ioRqQHOSdHAqeg0VDtLi+I4KusE2VBit
bRPqLZpjZkXu9qkk+sAXsDgcrXsK/gliMC7W3RtooATRQhzZOwkH0Qpuasb0zZ14
4CS+uZ8DO9+PlqjXodIM2pLC2Qdbkir9bmiTKmVXhF0Jx9p7xmYVCzLLz7LzFUsT
Jx8/OZIuFpsuZEzD+rvWC8qqeeniu0gAcedEdgvhCJYnhDhvz42UYFiCG8X4V0M2
Pbc6PA5FA68KPSUvG/qCs5xtfGNazpaNohTOobMuXTebjJibR6EaL50OymoZ8cXs
KUPDBf7oztItj6YBMDRk0dVl/xqFZkOs4+gVJKmHkO3kLQylAmzLOky02S2UB8DM
mTEi0JJ5PPAYvNrCvy/U3WTR6jnYT22ulEuH0lwhVUtdlG1NA0tQjd4sAqUl4VSB
4neW+jVMnnEvL9iWg4bsNUuoS2yT5jyCaLbcdOOCD9q3t6fgKJhtyFjwMNUxUyhx
BC/b5COjsu+XSL+TMOwi6Nfh30KfpZ+1p8DXzt1UDbjGsLCRmoh7zkR5iPPUR3r0
pkOEwJKKqKz/uxrVbmpQTBeViyVeX9rNANLiDa2ntdBkG2ta+leB84WYoS6L8rCJ
v8kbR14Su+VHhS5n+NEhThijaqeUr+mnANQTEgX9BJP6x67q6AXApGEP7V9YJU0O
d4JVB2pEaaiO3OGCfwggLYfn6RO9VVLQYZj0GrJAwCfvAfX4YP2yq9xd4YIToyuJ
Khuo2qvKV7TKRxcbr6UFxigzIPcpEJzXujaxR4USeXkCAcN4/8FSqyqkvxWlJYh/
1RkZ1vPka+/COaJpZ+tmYgNtEE7tJs/6yrapbdTpRma2KBDw9i6Nxq0bNW7EXQWh
kMzvinaSRi/3hSyJOkUxBuDgfZNjY4+c5RODPn8xNWDiRNtjYlS6S3ZhlG/itzef
N+I7bOkVQxd4CQMRnG3uAgiafZcLXoGrzahjSJK/kREIjx6Ngn03wGzEvL3GtkjR
CczTKFVa7theJH0hbnekO7CSolxuKkkdNcfa1/6GdFX7C+mHiJ4DDhoik8qSjZFA
EaokS0WA1c8ULbt7+rDheOS32cLahlNoaQCyPOi22OmyWctQGiMbyTdWo0REXj40
2pFN7NkSGW8/e+uHt+OT1rO6nOda2MW4vvBAY0dxDpsbc9b0jgLAfdOBUFeFlYpz
63QKqNbCsA+SsL7/B6SkN+Cq2NCn+OT6HmXgVMNZRsWgCibzq0tvHCcKN++VDNgi
1jBHQ36OC5loxZtm8/XjLkNN+WaftOAiz1VxaxccqeJcs0/HU4fKTSmmq8hcJDYj
1oxyOc1KqMsIYE/ydM+SiAJO+HadmPW9gcvTKVfGU0CgO2s2igqbEH0ROaUuB5Kp
RU7AQtNGD2N4Dkd0YbVSdn90OYOGTq7LWFjTvVF2FHsRfFqu8l4Mnqsv6D1MtpWT
Do8YjiQhZ2fXlPFjinqHVC63yFwMHnMHwnB9IhaNTHcq7PhaHQ5HW5vBzSssdQgP
xIygs9gMgU4HrniDu5v8LuYpLwU/pGvFoQXtw6v1h36UFrOM/ix+1XnCNpxPOTnw
8lIii/zdAZYPZ13eSjUeUeFs9uHTeNL6BBrw8AHgDBmeK6wPZKYJC5HOfnHavHj5
brcUaMDV8ZuFsjbZ9PsramGmsxSIB2BKCitaW//CncaB8AL/jRTj2fr/ozi3CsZk
hgxQDzUx6sZtGEJWQ0yMXbaJvCl1XQ67uT+qre3RkzojlFTEir/jahl7XQwZSpcN
YNJ6mWH6NLEWmSZ7icZCqCC1VZhWorE9LIoiPCLV+830I+1CZn2VmAGJ50ixlYSm
nrldWnDatG1jYE+rO3IvoKtTWEemuVfXVtyU7FaYb0rGwXyc/9s9EGtSkEWacYSu
Wv2yEJ1SJr6yIxvW7vYdLzHCPSz1iEbDiCrC763eKAHfFdIMAP7L9s/+taGQedBs
6YFqOnMNi09FkY1vLavu1JTpCBN7sjJibeDwSSujI8s8X3vjI+dGUhdZLfwTG9M/
R39HgMuS3VtV6LEgpp9b7vQTBSQI87iu/VG6sKawG86l9JJ2I2jdFvuwZikL0wWm
qSLdoRPCMv/JjP3/IoqD7CN+7ZGqQ7UrLF0VUCbnweCVMrIwMKK5TJjzJwcXUnLA
K5/kNPYml3SVahL4D/Md8CYWNsFoFygge+siQ4V42gPT9i5Z9g/M6UoaGVCp6f7N
DEZ7O+EMelEavwgDL08IC3yMEc/p0a5OsngL+SYgu9SKiFAVLQuaE3iOOik552wl
csdGP3DVraiXMwYepjdZo1CxheBH0TqDQnn03Ub4NyJA6EmGRkv89QBA09oqX5Nf
fXupQn2jQrJ827AJRFgmeBwCXn1Fq456teYgpsPjb1uKekw+6XrYrxBFrNxgS/RL
bVajzzMEHYMV4cKisr3YfwM4EZ59vnvWpzb1KBlvkfP8QKnkslfrpdxUzLdreAHy
mGI+RaDlFs5B+x4m8lwQyxBOXShMFKgr3+2dQwTjpF0YOE06WTtcxhvoDS30adwG
0cvo7WVD1j3ZlDcv6gxJltGQBbQRvBxSR6+wfWtKyj/rtChq0pzL39/HdJ2ogwHP
rZ6PhAvUYnjTLziMJrw10Ynpn/CEbvsotRuVubkMVT8+xZ5kEjrLsxYISUfCtrfL
hIqXz/Drg8uv679nOmqSuxI8fVoWAcDkV3YYqrVEMmCwp5Yek8RdWCgslG2T3gk+
GpupD1lqJi1GjqBbueuL5uuZB0tFnJCbOeo4UUOmV89SI4Oj/Zi7NPzl9/n5yq4O
gpqqu61+IpvgqO6a9jjK82YfJCqwAtzPOsfxDTZ799IScdzLP4F2H0XFSXszXIr+
2F7qG9fpyolIpsFWGiFC2ubNAcSs6PPL7Skg2oun0iAB+cqThzT/4pYSm5kQqaxL
WGpvdIdsGc9dfePa7wVDIVmEy8Tv7sxJjishA5p+UeHd+9xhQOdY+Qn1zZbmZolr
nSOfFFiy/0JB1KOrUOK5dC1fDKfoYj3+nSuE/PBZ7KBjOiehIs4WkO3dCjAdiOvN
VjyccPVNRphfPbMeadg1ELe0n0HpHvg8pF5+KaLjhygL5KQVhZob/XVh/CiIfG7e
4D1XADeasdTL2ULWDwYhBoLkxhVpMjJIptU+5LapaF59kZQa3jlGyuoWHAs2Ttuu
+ry244O9zcFcuk4oMaxJhtJjVyWwB4Njd/oca9ldRdXcgcF1tuThfLABjVLa1E5A
YfglOmRNBgRO0r7YjEortzOrW0hN8iVZiahKdiz9Z+xovLK6ww+UNSQW7DrRKhyi
JLbPSGDl8+d5ubruYbP9P+I4UlxHSks2HTfoD2AnzhaK+9FhYayS/tCrarxZ2WM/
OSwRQeH1dCql1KvBwNJzGKYA4FplfSjO2T2zSxMEbSKHvRmebo2wloA0bInweVmG
wkqfOduezca8U3mh0cSl7djjCZasLLFy5zDiuJ/8TgCTwN+Oe4eAUAzfTjGp0/NM
OqaaPTVW0KfNNPwXaM4hkW1PQ/iqef0bM0ToAetX6XSc+/LZy9isEZ0GQKpbGxKj
qjL6JlfnPp3O0HZrfMh6hCOFrRzCcUygmNzbSz3yzgBTiXfHAhbsuDvl5P+gNqjk
e9lLc1ku+NS9Wk3Y6zdWwXmBL4LfO4astWvimtsY0f0QyV/Kdio83A1+QIqHlhFC
QuQCgXk7XxFHJL/29APalPsSzMVf/15IkmyGLCQfuXBfBz5C86R9IO7C6l4VdvLW
eS610ADEhtQagTDr4IUkLtabjU+ihxiMH3M+i9dT6+gPmFYztVKyRD5IvtJ3B86J
er5epolbi/hp0IvXeROzoNR2GefYdnGiW5XG8lvV0mKAkXtJE55RnOqyUtnAhQSR
Sz3DTsQnigv6cY3QSPRLCEerBx0TyHoBFppIBxeHb6Bs5c1jBCV8N1Ja8s/Tj+5g
b0Q4JhAuSPjvyh8TVqEpXMe3+J/+dJ1kQSXEmtci6xi7LsDAOCYWDZpw+ikNd8Mg
DFCwNjZoxDMFvup7WjEWewrOT4/Zbg2L1iwbDaXNm7v8/Ulx+nd73ys9PTLoKxBb
FGfdn6t8ipALeEq8w9gPAY5Sa4G9k7whEbrWpFkUsdd6bt3iQMWLKmv9kBZQxIL7
iD1plxjIz4xcfOmVde4uALHuYadtHFV4DfFqeFTC0JOMphLQ+X/TZchYHKH86I7o
X80C5MpcbzLWHuaoDgcIrCIVhYcMUpMfJkfsGa+dfT1iEy9c6gHtvSORekLbsJML
Osku89EyYF507QZl2Zxk94seRNptn8AqJ7ZNk3nQAFu9V15HkPhJiWwz+xt9BZLm
jSDZY+9GtEg+YrnoFsPr8GZ1vea9B/sap0ehObUKGkMpv84PX655gD0+h0uHdYTn
I0sCTkutsRHyK4ld/WlNTPOSHXNrJvKf1w1qWiLx+e6fWSXcUt9JKlctF852eoQo
JcqLCeKA1/W7Up2/+ryqstoDHw2eadLFoCZeRJTnDeJVPxmHyzvY9U+b1EaGpMor
DznxlJSa+DuA+Y5kpBzGJkUaXjznHMFJX50K6SIEh05AZwtwNG6jgWbE3lTkjN5Q
ypapK01JH8yOD/HQqaGc6MZXmliUZ3HhbJ6toIZv5AwFZADVsg0xUJrQNqL4B2j1
5EcakNbmL1xM+1s9q6N9NPd3B3MTti51U6aCiyets81V9fxg1GD9CyQBHgn7/ibK
hix/lvcgKHNwPZn/xb9p/FnaPwRrcDqRA01mTtw3ILrHNjbC2nybFsrRlYFaCZIl
qxoZU2++/L3YxoV/BEEGcPHaWdPN7OcgjAvjj2uu5ypfqJ1Eo5lUrp+d8F1Vmm+c
8j16aAlR+XsiD4Ca7mcK0WU0Lysw6zJWMTkODDCdsRRApJFHInozCMiYcqCUr9um
xiMk4BLcpewcpSnmzJsv6rz2pOVcjKNl4p/OmzkHrzh21ameoeKI1XivvSkTZqCr
E4rafuzVstZ90+PeiI7xyHYj2lHVPMth3Hk+G8/towJ+gR4wE08UzlMgDZuyDlOR
j/IL8hyoIqiBYAukB+UEjlFeA5Vgp7oSJH5G0CudlUB+LWK4zq/Vzx8kFkgwzECt
OLXRWPdzqIto5ks6l9aRPpcdjOVCxMqPnW89124ESgh43LhXPEiNKpR6l6Ir95TY
gGdR+hazID98A5OEwEYnbw50t2PvaR3asg7ky8Mlk3iAlz98O8ifTXmAMuwg0Yd2
6mFoQd+a3NolNvHewMZjE9QWKY5f+d17hQB6j58tLMBu4aX9Emrv8TbdXyYqdARS
jaoq8GiC0U51EKgvvifZti7Tg0DMz5VjCW+/ACQj9DKkqqxNGR4n4N/BeQQdN0GD
U6m0pTvEFy/f2fXn0exxMwfLB7MmQxM7+2MJzC0qaHpqS5/ed4lMPYyEMI5JjEaX
0oVj1sx1U+EjAh63TnsHz/IoBM0D14YtxxhG4P3q5PzCujFn3hkXTSYfcLydq5uR
9syPrh//xWIJXN3pN0IBQib+1yXxcig4Q5brrieHXNFlC0LiAKkSjK07cBcfuoc8
V5Mlqnu27iXWMB+XtiyBy4KCDHGPSkWuVf2ewMJLT73aQjntso7Bx6pGvvX83QCe
gKo9E9SoJBj5zXUik9CRFNtPorcf6+r5JfP4v/xrAxjAtCPKYW9JmeY1dN5/0AOG
ARL8gaRcS97zoOujql7m++Dv+Ad4jcHAk9NVA1qAjURTt85GtvFr2c65Negra3yc
3w0GUFsaSKfw1uKa280BxUMvIxpwy7a1YNrMG9Au+YkU4uULzhqpWsxCpPBO9AEa
EPQ6PZzhMP4cI9qLgHHWmJVlKoWjCyO6kTMmToChJCEeouNUPcWYYIwRzr+ICTOS
XJ8KjTRA13OdynC0/1FPsowIOEQyB9HK9xjXVbkMvH3jI8S+uAkHbP8a+u8/PT2E
xSZFihmHtkv7rfmdh7BnPfKNlsOtE3YifXQcCnAd2NSPhGDo9hYvqrCBdCs41IuR
4sTAB9hwCcexCEothOzTRbjkb7W1pX0r7blUtSXKdopw0CPw2O1UGLYlTfwm0rF2
ury7qUy8zxFJWJoBaATDJLa9LeM8Sq/B8wyiG6a4NXdYb8bZMpwgMw2Cbm+vzE+p
QEvXDS35iRx8j32M42Q4kZP0NkTv4gDrAcsZBiyP42+/IGI7uoMgbQh9dID1rsbj
uGL2Y19nzyAMtaiRlofINJWGDfB+fcAx4KScCgoiswySgK5hslLsOULuVCEJnll+
AMJNGOdCNBWlhfBex+COtBODByDDeM99FcxwRjZFWjrrBcMIov+p1pL+fR3a1QM6
K2bHRYRKDKyn1GqcWjaqQLLl8ju1ErMyEVCB+l9kuCd33oq7jbohXlNCX7P/4G6e
tg7RX3yt9DhepU3IDLXR09ZRxfqYXt877qHFdwCxCXU2ysEpV5/Jc0lvDrLphUa3
qHxxiAFQjBjwrv+ENihMZITyVzimRadexRnKtXhaLPpQjawyGY5OEke2xKWdbgM+
B/zyWU5tiAFwZgHHFhdTN98qEuXuL89gHfT3p4rbUOI7kxcd+Nc1ZhfzX/Fb2v1U
RF1T4vtAjHuC686m3cEMn01aGNGF1VEaxkVNWq5Kn4H19WgyXYpuskdPtFkaURuU
WwgkoNqGf/ucMdISapYaXH2+Dt/q/kUVx1FAL67C3VHJY7fF7/IVx+QaeKsUjVw8
cXV6GqSKeO/RX7RpKLxBx7sfy2cBFDUhrRpR+h7r7eqzPNQjpJ+fKp0hQtpqz+7k
9j+rsxIAFzypPLwSrLpr1eRfYMM9P8/ZAcsyEg9N2IA9fE+1Nvr0xr0FYng9O8+e
ICdT+veAK/iReCTsAtF2IGQsu9QCZhI8UEwCStlgLOqstHUC4yGrugz8oYhAUJuJ
9bhS0NhMEypg6Pv/4AJcihqWZckRI+d5MKfrb0D+Jmim7GoZPDA6q8XWLRIaqEDE
tPDuQl1nEF6aNYtE4MLZfQE/mGe66B2SF51f2pXDujnnKYtVXkujBJlS61IwOY6V
60SM5FB6I/zJy8PQ9Uo2T6e5Cckn8gEuZBVkaPEUzKrI6bdEYQ2vr2rITNqh3eTg
Ls8uHCo/qAhfcOYwYylXZsh6SsbO1kKrPdZcEz4CF93shZjBy+d/tncQ6xq7WmYd
WTNdiSnKYefmX/bqxsRZ/xJy669birU87pH1pj/H27jACOlmWb+794EsPYtrx86D
yucZi2ozFTJbjdyudNwDt0SvK2EEEn3bLk1aXk7KL7MQti3tIeWalbtq+URofA4T
/I4eoFjyCIPuyvhxIl9dipHbXd0zzcT3FNn2WNj84uE+gqoNUVQ/NHuOHW8Gq1uC
A4h9+xs2tsOHs7ltvOBBA/tdztTU9Y2bf+v7EuVUJ6IEo3sLh0tiYefYk3UugoBP
jMB0ihPlxtFQemR1N3BOnqxz/8YQxQv57O20fNbDKzVUfhhuehpIAvSDZKKW3mnP
Sghb6OO/PsF4B+1Wg4oBh/WNeD594HwvcT47zcfin2RCtQhGoTuNhGMk6dbrw/sk
PeyZcbEjyYgKwKnoGben3e0pE9ihNpmROrpn9tyXaV5K5ER0evBWcbkKDDPQhFdd
JxclgniWRd13LglMeJ4LkB3R9No0EUKeHoppnIfRbltx2Uszl8FmXk+KPjMsGFMP
lweyG8ZA+W9w5BPHhZCgtGQJ/uvpWZIXlzGfDePcGBOp3fCWKLiLA3xVKXWlhj0o
9HVoupwamPA8qd/OYhS4jiRLZWRtCYxD6OtmbKcf0ehLfmCNPmYbukcMx7YtZne5
aPuG5mpjpxBXNijQYbkvyadLLw1wTAM8dkODhbgtWTkodZXx1YdCH30WmesiV80r
3V1Jg0VTmrxc4t0fJ8dBVoZcDArYONZfADJ/Ek2suDtiArMd+S71ERIGNIIz3mUq
g+sVNAdEIxZbMEV3AYI2MFJbD6TX7gLE985ViHIyTzxDSTp2T5LVM1zJJPcQfUjH
xNhqYmN7CXoEfMuEA9ilqCim4gNepJh/W8H5kLUBdEIv7nVcAWgux7EjvpGP7sCG
y/gHMz7Ccc8+dJv/Clr8GoyVhXpRRfxWCCSsEVtC39bQ3PSnPytYz2NBGTmCaW4x
3vhgpbaz0UdOmWBHlNV6CQ3qAHmPrN5bzuGrwPuM3XA5pI8b/KN1/HQvf3yh4Sg0
uoLfSLYsPO4V//h72sZXQ8ARkzMgrcG7s365DfpYzbeOa0YrKf8gzpCqbvuRORjX
pl5pRuoYUKk1lEagR2Yc8J4WEkIv0ZSWXOW/6FPLn7wo60qKAOX+/glpOlylZcTG
bnbNUZziWfWM1ShTPGHyrkCcVRkk7w184maLLlxtVvc+9A2Ph7fQfG8SHVpDo0Rz
R1Wv8oYUG4oEkmdgtsBO8HoWkQc4/GAB93Z8nbo2kz2AMDz3b0KDMMz/1f3Fpx9h
UZLOq0lG736ykey2dmS4FXsAMizBJlK94dDeCWG3+AJXFwOJ6aHO72JfcxgV1zll
r+fReXN0zbeqejsDdrVS9WtsxV6SDA2lyGi0O54swyhR+AHyoPhy3yhwu1gIpjv6
jhNGWPbZSLl6eooPt3j9q7C0fEshizyYzP1WRvgHi0wm7Gy35xMpWnCW7trcxgEb
kncjj48EJXen/VTalJTsbCqVGne+gURIwgFXa2XNOfRRHhjSOVFKBgKYG7pMnxQU
t0G9R1fy8D4SQpwfX6EmTRgKh8CM/12hLzuqvs0U8RBt8759GAObF6YMM0ych64x
63zHHGL0WohET4prnhEIigQaLpb/N46yV9ttyoon85YrN2uqQ3lM850Sr1/ygiKN
DB0H2CrFXkdMBSgDB4Hnjgpj8uNsvjQJa8cKVwepEHP1e3Y324D+Fkfurc2SAV/t
36N/IRF3iLw+lOJO3pLCXJCiBvCI4OnpCdavJOw0pGZQRC2SnEn+DOXNzuOXSyur
93R8+1C35TFO0VvGQubIJ/14lz9SSEp2p6R6zmUJ98/W3ThfUV4oFE3OjymMczSK
go5ZFU4SFdJ0JZUJpuBzcWUxuJBEI77JhDW3w1R0b2eD1G0SbZRdjFMy0Zm2J+Fk
LXL/hajyQuH7dYz6htJtu2dn2gX1PiFizSk8JAhhzoN0+26cCgMyWGC55f9kOwS3
zTUGdDE4SwvmaFbQZbFvPT4EFSmG/hepbKZxmgVn+HsDq6v1iYh4osBc/w0ai6zX
V8XMXTdVoj3d9vgtLdDiPjreve82DA+RE8ydL6yKUnZFKqxZBZgcRU5zg5RdTOhb
BHzRto/doexUTfQPWTrNaYnT/zJGr1C+UpnQZY9L/7Iv1jKPDE8Rlg9zrAiu+laZ
YJbEw+6b8CZ4A1X4W+g51gWUngsPCu/Hmu+Rn9HSIoX1UdGDH362hBDJLBtZg41V
dU9YIhw/CpuXdP2ZbmRfhK9xvUipRinGrGrVSgxYU9Eg3y7NdWSguvOgd6N6YW5w
aUEhfpQBZNgLrO41aHTVlnv+8cJI+gemJx/m17j3i+1/BnSS5tFLBKDfB7cldaew
Tl3d4WCBfCMpMMyFb3g+HO1cM1aPbG7hL5pmKJlK8oF1/XaInaew/fcGsBLsBU4i
jXV8KQn5SKoSGBh7WypyrL7sSz8yUcq9buiCl+t54oZJ1aK5OljE0OxPqz/FCUu6
1qlco2NmVdzXOTcYl7zRk6R7cx5gJ0neOjBjlUInHuB154+j7t2/PoPqzHlCqh+K
ZTeHW2zcCJOOZg5dtIW6++uo9DrhixVZvlve4nqyc+UIT/rxr0rAfY7yWzsHlqvD
nFJPH5UMo1S+DYqYjLQ3fA6TXOWUqjlNpx00lAGtjVmqT6NuSK9MdI5Kyp5iL04v
8w+GYxp2SGuh4uOY3keHU/boSzfb6m464PTYrpW6WPZfwhz3j+nziIfWPWeaeTXj
a/UKEfzFRU6BXPQMeWInwbZ5mq9mcYxPMsPYdQtKX0HXNPvRuG9AVfO5qAXJBoWA
68qCHpIdpm1P2Rf5jLD4SdnXtW2V44AwJHVg7+D0S/oLAtIWxtvQxybVaLyiEdUD
YEQ7Y/sawSfQYz3BUsxDY73pMlaVfMLo+0k+fgU1BHgIMDp3haRAuQFa0886xRHn
MhHqwLi/m06x43NoSoDjHxhwY1op0ES/MgLFA5wlgSRUI4ntt+uTKtb5EdBgjnWd
54dE1EOQDnfnBdV6zcm9zDKv5woNt3AwBIiRCOWfD68srY6lVIrai7IBEUv29DZl
9WX1CdhpniFcU9rRjT3Xm0UTxSaFgUblUCjUD+Q86TgJtVvZcKSXVp8OVtd3aaxO
UuvxetwpmmyvaA/5YKPdOGke40zXNDgMEFzmV52fWxvLybLoDHFupQlqxZyNbpT3
jeNmAbsqeQ/ebW+tguMte8Lx09yFUrek7Arh1vWrr3atwwS/nsrSt4WCckWU+kqy
OIZWpe2ssytqjdZFFgT0vK5lcZzx5U6eEDxRQ7j0MeqYxPNJv6URVdDUIvhsDLkQ
NdHvh+9UPsPCelfZcNB5eWr0Mha5FpeBP/UHwmtfSqoZsks8HcAB0GgegHFwBJ4U
8HyfORbJ9U/JwGh95+QyOagczHIkwNWOgWo2eGOvGrzA2GbXpW7Ph+3Mq3o56KOu
izXcJ1tT5xTuPNY05u6yXfZEEDXeUf01TnK1dHtycYa3CuQBAX4Q6x8GNqX3in+U
OnvQIyVMdXt96ZzE98so/jj/4+7j6geFEdwzMJ+ExJQtSNGBdSL3gQTnXUwsHSc/
bJEWiowVTQlbdu/xE4FCOJ8H+FV9GReFlKkf70dVs+/AaGeE+RHdkmkNVkCyQTL+
l2PqBm0mACW92LxIzSA7tmSdoCGyfys3rw+AK1RPPXvfaQLjf8KODkCbz4oUdrZa
g2e37rq6ARlzaDGrN05AUfUtmdArVNKtJ7HTfJhVry+THYLQumHh7Yj7xYrjZVC1
v9tHpzsfTD35t1Yn18+UmIPeU4v6M3E//zRcoWJkfbwCGx4o9+H2WwVV+sN7fShA
EuP4dczFfWthl5oB57wbvCDk2nzcE8CHJaN0StEH7VX+WIFcSMHIxGp6abseGQl1
7ZJIwMaOOSZ6KgBbtiviFCps3wP2o1eH/l+jc/wR277dUKG+ArOXx+PogfeCVoSN
9R2mbjP2RpqQB4uP/Jri4YrVvlT8bsxw6n2U0rsq946v2JTnAmjkqLH5xnmcuoiJ
hYdXY7HLwGu1Y/KMkdWorOimbH2yvf27ciz1bWEqk+dwn5iLzIErJ0LRG2RhTfDJ
5BvbQ6Lt4wNFbHL049PHXo8EaZXpuLtmYz9hEp5eorjdFF9j4zRKSlbJTEMwwBd7
dE4YlzQit3WiQVAfa6hLf02y0Ep0qToMgri48PGJcJsaW8g1K3LsR/JxYSRSoFa8
Mg1cTnubj2DJVWbgTRdaknlmmkqFYJqtS83OVL2pAlc0WWWeC0sHOW6TRwHIlaXL
TkPQkVP7AO51befLhJO+I/FSsDsI7PfGCSI+/NkyV3gJflq05ndHAe7Jb2IwXHo6
IRCjQZHXi3+GGQCghRltnIe5qNFJ12M9gl5OTYmHp/AR513sgv8lvYDwvyvb4QBE
Kz5+uJabh7gWchQCiTu2etn1dmheZULMejtjlvB7UJdoIbtK01UHg3y7BlkkK6b9
G9N6HLnkAqiySQ0K/KsTwwAMkY8yFbVofAPouxJ99DNJGlurN1yYi6wf98UlIoWg
FJlAGUy4M2YzB2X3eiYLcmrlhyEDZuvEMOy3xftdUne2oI3+EsAVPdi2UA8mWwkZ
YEgdj3keCoqhgUWhQuB3RCEwQMPePI3fETsVTo0fSsI4V4F1k1frFTPbWSQSd0vB
nWTI5ciL/1cqUGdz5QLNuCW9MU0FYft0BtTtnOjaOy4EoNAs8xInge03HS2xofTt
VqHV9aQwvft6Ov7WYcr9kWMjkocUmz5wC1ntfo7cDIT3wQ+iwTaX0F2z2YdUi4Za
MRa5LOyUA4hrSkkI4OZNtPo+E/VkEvNsI7bgSp6cqlXKOyEuLntNy4TGpFill7wE
OHefL8YknT4lluXujdo5z2ztUNCq8iloiujMXC3e/EFF9mhyDiou8DXf+LrZAWRw
sWnEff70t9mq9443nGfsDMA6b8RakePC+69SciG84KjPIsjiVD7bRTWTeySF/fbw
WvwZuFTfLWPWzIJCnuV0gY+pF9s0NAvnmQYR7T0oN3p89FrihGAPiMfroiaSDoHa
PTsWe2JkeCX3d+S8941hyXyXTDFrYQbD64p8IAX7mYEMd/QtDo0mwJhCzbtrkzRV
uCL8+0yvcvYdBedilvMP9CsL/bSHRwcFxThs030Z3c9Ax8imCBddrTGTwuLaG+Js
0ZnDe2PN3tPqTG8UhP/zIHYit/jCj730D25fWUY7Mubzd4BjbtJDsRX0RS4kVifn
1ZVJO3qvA5iFvigTmgRJwv+YoZsXn1ZAK0q04/0uub4+sfKxg1BizDR597QEKTC1
SHNpOfXKtAZGz3AkqFHo72SU9iKFnoYVklYIM6nyxfQv/jmbGs4jkbtU62XQVkng
Dzcd8Gv9shIAl4Zg7VUkF5Ah+GaBrQ2TvUw8uFkKivAGTmfi1APbdaykEbAtka1I
MIfGzL8yynsYT4O+blXKwP5LkYJP1qFERqJxCB6DycsrkhO/yoG3BIlw19FHusIr
5SVzHOAWRJWH0CDyAg8KsTyDXQksc0Qgam2HBD+q9ExcAenlfe1wJFBTXEXJuZlA
Dl0CNn5NG4cswjoZoZht2tbrggvmoZ5mcPd1tJSX+WVpK+JRmYwI9EEekFPHln9u
v3n2uTeNBSDyL4vB4WlKq0hg8kWRQYaUc9UOvtpGFUVfkMTGo6RWBALQZG87bBX1
4tX/MHbEl0l5rxYtO9UmXl5XRIQezd/h893x/ONZGUMVVUwxfeKjVvcW2TuQjNmo
KVxfHmYm411l1lf0ee9KguETUoYzSS9Hjxhbz9DuGvdFIBImEiPIEjiqQPmvckeK
JwVIaYMxPboxqBXkNOjjMbHc0rGLexpr3AaZPJmSV/zpFX3gIeVWNeHuA3CWWL6a
ybtw36x0xJq7slAXrSTPv1cn9v/06JL9q+pfu5wf88ayGL79ZFx58KpEmb2I8sWW
8PNYqm3hOwnTP83KW9ih8sqSYJfFxZ4cIAD+Q+I/dl4nSpC5U7MZ92iD2FwoED04
iOT6U51PywctYluiChpZfKH8R93sipGkvyaMd/u9+R+1hP7hnt/9ehBoS8EBZ2LZ
C2ewnWL6cfpk8IdCy41onyymzSHxK+3TfbYuaOL6p4A9gqA89BCSaw1BdVUocr6k
BYHO260GlsINLe+mq8ojPe5+nxYcjvM+Oa7bVCmjAG1dXb0TLKwWRisQpKoEM0b7
l0/Ru5ATaM/1fDj9FOGXln3v/DHDJy5a1spoJovtLR4+6KNrCVCZVcKL5O4nqt+A
UgqCJhDdiNwKQEdsAA4TLoXOpreZ76BBmRjukSAHydP1PT/ONLSSDYpSbtbuyErP
wIO+zI3ErUm8D7idvihQG81mwlpnP6fSuh1cLrhbbd1FeIRy/peNgO/tJ4Cq2YnH
qvQkH4OZe1xx+qhE+RhOIPuxahUwtY8PjoCz+FQiIIe0xKe9hrVQH84ZP3d/DQNW
H+h0AQbwuT0Ty+KADXOJeP3kfi4zwiob8jarrCklXzTvXPHx2kVN1YEBnv0AZLXb
mA0gDqVlNaFXTEMKotaLzSfVK76KKYdPvwfYv4jrh9pQGUnO4g716Db9kVOg2m1y
9UR+C+FPnLYnwARzh7MgUnAVMM6o9Nea24ggAvTZx+XNKn1P2571aniOHfHWQ5jR
/GSoz6kDMstZ2tcuZHRl17CfvkqNvvKYAJjct2UWMx5lR4NZomddJAqdAEcF+HFt
6kSdy/EcxkiSKfkhispZjDAnNu2mzyY/M831gtSwGMSu61MBHSmGO+Q/ugsMad6t
mSCql80UVjuxw5SC94qK0uWaxgkvyR03RgFtgx+6tJBSF7FXzbT/S9x5RHXgB/EY
VsB1aJyDfqdkSkcNeYqksdTrSqqCRzJhswg16d0oTDneRgT0mP6eSYIgcOe8Qmbn
pfk98eHe1hnK4PG1Txh/MPkS8EcUJlLwrSrDsbOrtEfSToIk3Yxhs0hMnqYKsRt7
rktVvmGsB9Ntw1ckug7V3ev3GM1TD64f3RAzWz0Q1PVOGMg5Ycr1Fb7vWefRYfP+
INzalmvL1OwryhK+DBrccLBbVT5VJ0XV8HhDYpNdepPWY90KeT7BQHf5ES0ZmeWr
5VcUTdLv1DjMFkloO9H+WbJVfvxEg63Ftc+mQdgWdAWsZuxKSP0ahn91aWq47HAh
6nhpusMcvlO6Lt01L5HOZTcQuPH0ztVobkXauRQ+jAAotoe0TuHALIwr+oCkBx0S
YY46ZK16iPQsXiQ9hl1SW7xc60H33SOB0aUi2qCGygBt4oFGC4EoRKgMSUa84X6I
QIlJYQna1YAhbwYNZ+1d53tE4MSKpP151BqmRwNKpnHNYzCS+mS2BMDob4zQVA8n
ebv4x6l7Sni8XSg29SU/rAKeFpMRb+NrKMxMyggmJwWx/qf/pv4Wv0FkHR1NudK9
sORRaeuHWmd9ValkAfDSqhE3LpDxcIMUucr6P4KrRMu6z+jbdo5Hw6nqjKYr3E0o
hJbccNGTWl7OwncK56s1nrqchsZ2rv707a0p0jmpAYuLh+ufMEeIfLEn7bKaQNXF
KqOCq/kIQfK2oIHLNg0PgdM8h8f2i7MIpfeQaeIEhVzTUb8SAay4h3twb8PQR2Ch
9tG1nXMtdXIRsO6lx3HGyii1k3lGOCaF6miNJBNlUvfFlf9unRNe3WSYD3scb0Wc
QK8aXmDgslgpfqYYTcRgJNh9tDQhC7jJ95ICuzWC3PCs4Rjysq1ktNFunel2ScqF
0iK4P6Arl9HEOii1XMV8HLhe74CAutoivkup5yVtmCTXnXe4X3XtqTkeGSxZWYts
pMKwW3slRVnKKBKUuEekErMMkJ5fJOYVBHInVNrMTR+QETXQd0xmdWLKPxhyjEwi
bQ0m8y91vAFlJYRgTQmgzuN5SFsysiW95mCOYrgl2eDkLYoU5dberGVhACEeE2V6
d0u3VLTugIH93PK+Xk5aZT+IzV4ESzGYHSJ+6bWzSMOx64/HgTQ6ZJCiTT0o/6Lv
Zdx9vdEV2cZfb29TEkORqQd8GEnwU9JnBwr23L8cau6TfkDnOM6A9Ppw2xlpd/R2
CtUVYTdBPbD4epiqGCauxOi8ww7W9CHWNScxncf/BIGWj6QuufZ5Fy5R2ed24CAt
fZjDhwXUY9HYabuKAsdqWOfoqAjQyxE9UfUUMyEs4Tzp1M4zAiSw7wWW6RYM+tqX
VNArg1uOoaSsPQfNvuOBxuIcSjBKH11jyOEndp7WMMN6cK9is5txatL9X5vDti1K
FKkTMjanrFlYfqvSEoKXnCjPpY/fo6Fj+r5mblW7Q6hujQ1PmVGrkliAh07WgSqt
bcHMPW6lqygb/8Ho+J5vM8jWO7djhABgUe4euAh4LDOSm9X//L+JL9lrFCP58L+u
EppfOb+E7gZLY+vcOsKIGpqTvWhUAbH689x47Wq0uVnz0Xs2gtmzRh81MV6hYk2N
ZmeNZnaHg7c6U6b7yDlWxOkr/vk+lEdDmgXhwZpkpinIDPQF0fF/9rKLEh+pSOVc
svN8hbeFZxR1rSd3SGA6Po7bxmDv2Ge+qz4lJmXKcgW4F/wg+FwLfQ382mnjIrdf
o8Kor9ebSyzqxVXxNZvYnur1j3YnpvwlUTH1jc/dZMefcuccSEay6Z60isT87P2u
gXyQtKpQzeZfTFI4z09xz3vatGYoS+firL3lwfpKtlWe8go+Fgq9Maw1KTgalFrj
QoHGG8kdoKA9lwk1p4BYykEdJ6+Ho9cWHENEdgkBCIkhP30uOAEbDthtZl4XmLLD
OROJpRAYwplpqkj1arUjxuBdMMzn7G0oePdaGa2ya4joxUztO5nptn4YoxoPAcqa
I9N4IglRHnDwQQ4qyTWyN9JHf19EpUpqUIfGPfaIQHGcFXp7dig267ExoJTJ0r0h
HSQmVlIAWD5KFMW6bPIFgjOfTcQDyv/GCLDcnAEWChyG790JiMNz+hsxxp0s7BBE
s8VoTrZIEaHh0zMy5SLsdwtjryiJAgU7tPg+PELfYUtZZ0MOZZvB7eL0NZLXQY9T
uUfD4uT4lMGCBXhTTo8ccRHr3LK6LYelr5vnFilKEqyVbCGmg8E8Z3jSIlKdAivZ
PXmNbX5SF+PSGyoFOwNhTnNuJ9frO2lK5J4gH2czr2tAvfDabp4vUXDi81SGk5FP
nBcxgtG7GECZC7oVWf4AsgJJtrRrxsB69YzAaf+JKkWqGAFYRvTWtl2GpBx06BDy
RuVPYf3rapKmz4w/+IMKt+AzRBZPpukVgf1SDp1FGDiXjYpys4oDdQ0Yf0QwGSid
uph7hsEPlRDZhR86dnky5h32yxSPJTjFMwcx7E2RB3Ur+pI4kqEP/fnnX8ztxsDS
SNdHhMJblLhuzYOV+uyYc6GYb8hXqAeW9VMyj+aoVmIMQzkXzpxEAANhvnDuClxX
CR9QLwHj6QNj3egfN4CTSY59tooofRzSBsZ1ASgzQki0STTey4dvny5FbmxwNwqV
/kSN4f8qFGKGfprYXLZz2Xi/gS0IS7lip4YBCrrruHbQ0IwhtFPkLAdprxkkAxZe
Rnq7TID84/tUXShAcI+NxTqhy/JjnFijeSRqLYQd2EHg8W6TDSPjvanRcNU3t5T5
X1asvWqcSnYOi5pK6XKJ/xBkglmcGhwi+NRhtRD6+CfLMs5tmSZfR5zykDkr1sHM
FLG6DYbQ8Palu3rPA5M/4XtPfahatErcbif/Sdc+f+dvyp7srAbEwy/ZIjb++BVN
ezvtkCMqgY71jDjJzk5J4RY0zqHO9wP8exBRUvVApjaHixazLyasVHt6+uISgH9F
cfsTqOQ94sKePKOJnT6t1pwJmJvDhAWN+nqvdeMWUvl4OqkbEI9U1z55d1Ztv8cu
cfKaBvoLEnP7b4xemhsqTXhWSa5vur44ORIjZ3bWms/yg9F6jO1j6GDd1bhgrvFC
MJWqy6sTNcX+owyuYLLZJUNiJS0yRgHlVMjBAvXzYsxj2Cf1QU9Sk6sjTLw9tdkf
FZm6d3wgc3D44GzoLEbAXvWxdAyoA2UleE30p32quhtk23CFBtb9Pjli/8iSBVFz
IXGhdyQRBAL2aIfwuNdwbRnhB5rE1hCEmiStkJrcebxaPZqWHnlVL0jmWr8G96E4
IBshoZ4/e3GcGxjQe8wcGHTJXvREHYuNsOQZNuFrmH7gs4VkJR4r6QNBEeBWARTZ
lqt6266HiWo73ImUj8h+ANi8aePIJdr1sl/6NZQGIHytnimF6Ba8Ip5fP/Xw8PAT
H8smGB9NVdBL6WV0DQUmD+y+Q4yg1Ly/pL/BfNlAKWALkwGSA0YxRlkBnhJ7ao3h
ThrtkZDGMfg7/HAUKUDzynkzgJXr6JWd6bGZe5X89dq6ciEShzcArElfdoPvPi2/
sLK0LWfo2qjFc0bwu6iWb/ykskVImbSoUSNJmrpjWDDHVrlyPD+66ZMGOUco9PnN
rQeUEcXIRdXMBcsSz+MvoPkXw6Fr7/YHPVKu9G+FydM2XByd1kdpPVZx/BaBoPbw
t3vwKRBCeuif38zctFZZ/z1NMfwgLiaHPh1CQ75F4Qq1J4yAeO7+7RvNUtSRunFt
QHKJEqAQ3cnjwu2cyo9riii/VeCjlNr4Qq4ZUVVZY+ws9XoYMHEN7OuIhWCMfNed
cnqZx8rqMVlotTNMT/gH5lSrXsIALhXIzX8/o5YQ6ujL8xyKtiIA91XWvFairptv
JwImy1BrhTMuSkbRJKbqs3T5L/syyvzKxIzHNwspLS1FeUduJ6+3Ku2f1LdzjKOw
MN7J6msi1ZX9DlXWO2mEQe81LjhufhMVs7pkpRcJG6crxuBrZCL2KABOEmEhJLus
JxFX/ByO/Pto5Hj0zUqvszmaX/1oQEjHBpA3lQMVzXz76uOR0sKHyFvtXlnJAlOr
QVUT6Vovha/4BlhmrFFahnuLsJhjp02RTbeoLLOl8qzAKHz6+ivkvBYL5TWTpix6
wq4Ed7qqYL7y+W9mkaRaQY1MWN2DO+rGsVF8ttnTZGc8F1qZu+N/iCxYdWAvmk4U
a29eEh0ZchePglHOts37qo+xJpt/jfGhdWPJ+s5G+dqR2duolNMug59R0+i0Lsyv
+3oDFxcDOgVNKpQFGJV0RiXRaf/R97mLwwBK7MoqCWMqUvfcA/ejPsKZvC9kLN/3
QDpfhL85IHpbjSUC08dzCXyXixnsGfsRxdx6/XXnz5F77wagvZCnNFdQ+XKFBPjl
bmOskFIeYDrNs/EKACxFWJEenh9yH2GY6dE7Q8Btj87J38rmde9RV8qtToPlVqot
SZTwDX+PM+TfTxr51bkhfN/YCPQdVVfy+GFn5Fx8WEEf6+K5ORD6FRgsTYo2NEhC
GjUcaYcfTDIGpGkyZw95jJ8UefscDkysJ1CIVilfHF2qV103cSEZqywSDdTLHb+5
IsE11q87W4dnFOq3ZlHdAOXkd6bg7x4aH1uD0CAVp2ufsEtQqGOFUJue1uSShzmN
c79F3R63wH1Yn51Jf4RsnZs7lKzl9+oPkXHpDandzXGAQy4JpVUOs6xc1g/MSFQn
4cinVqNpIJkJAO2021Xk/QPPD24l0DOBupxnpuycz/14GcsBblSP+J/q8XDd4B6Z
6ePGH9mZ2sUbj17eE2lKlhwwI/vAGbggw0G4xjvp+HhRnNhogFPSMZbMAyilysvn
gq3lIseDrPYSHLMrO6UPtLQPFT2qhiEj7jl37wFHJgjDdqqGX82FM/DMzNpOl1Oj
Eq4IBwm0WdLLRM57KYjyW4z5LNqCChnW+O3dhf4Kr1S2M8Tp4GckfQbDZqpEWalS
sEH5pUNVrB7QZd3iAxmwJ3IjWT51NuHA2s50R7/vzjh7cxfwcpvs6SASJy3z//yH
Ygb0D/F0wYwzvba5kPptvqLMDJAQicyGNEcg9kiB4zsMaAMfs97tLZKaWFezV3vW
gDiszPpxxv7mldsc0SqjIfA2Pe3CYUGfS2hECFl0vwvrBhkqo+M5JUy6mdgHBf8D
SscV+npkHfiErZnQZJQF5e+CFdVoPoHJZnSEB89W5rKY4JhdL9P/13aRBLtrcSva
AckD/quAwd4NmJyrGg6wO+NN0tMpWUd98KqKdKyRIkvWyRNP97qdoSDz84hJ6w+9
2BIvK62IWZYgTOW6dBRzLd3reJ32AmtcqtiqUL4GivninkZcBAQmwfSNYPv9I+/K
yQz4H1VDp8Xz3KfpofCTiNVAEeJvRtMJOcIiquMlQNVxbwLRp+TSLL0/1Umq1ZMZ
RLOHTvlsyBLX/Kcbc2uIBFs3dgHiYKNS/uqIgcb+mNoDf+Kopt3jFxU6Kza4zeKE
MZZNuYrUSkSLQ6wnhaL1o87CMzTC2NxRsgXw4sZo7Chb6PuaejZWGpy9YXjXcoqr
cnybqeA9/n3EK8j8U6C+m9wtFoAO08HSeifOsSkUuh6N1ZS7VCqPF7KC/8W1/8pd
mq5zEH4mVnsCemZ7cIWILpV6DpnjfJZiRL/cNgowqFr3IAUqqB79Ejs6FuPbm3jY
olj5+nmE1aqOfqWBNTwRxbsOJFPIt4dLFP3qFxISkrYlETvwmSVD2X0albHXQmRH
rLWUtMsTzz89GQAUrvMwACcNernWcDRTf0S010oXV5y8Uwz+3nFzzUX7I3A3Kjpv
f38fTRTDJIwTzJ/HyARdgjSuMtUEzpgDXhB6/FXFjdOcz7ev9ayYfpVpq4k7Be5V
vFerQEfBr08L09+qjKKDu97HHUpZ6fp57/i6/eCWU28dAiiXqn9CsSNktXGbRIwH
fww2bo1luKbvAnZiBVvGtQ==
>>>>>>> 426889eb8ce467b9c9a9f74dd4af433c5046285c:deps/flexrio_deps/PkgSwitchedChinch.vhd
`protect end_protected