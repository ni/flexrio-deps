`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4128 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
8gCk0uzRa924DW4s3mkpFB9Zo4o0LPiWONArfl44+s0lWqEq3/XcZRfZRHT7ZxGr
rNa4O7E3ildhwZniJbd8BI6DvRt1YHotqC+e9jtXJOFiQPI0z3XxZwjwr8U1rnE+
bxhf2+FoA0+o3vkdhE5AhtfF1b8NSTjnfxuIC63vtOkn6oAp8bqvGUHn4dFSIVC2
R5bl25QjKX5kKVk48jMCyMnQkH/GlSOVxlHwM2Tct9dDet+t9DX52ULDCBL6Hzj+
+EkBTI3mezmcYUBNPrE8vkwP24lSyFK+admvpQx7KFtLeT6l+0R9h9tj0z1Kra+e
0YuyPqvueiSJb+zpmhnIVeip/FCWR4FOfY5qwaAlbqbDctVIHN14cytK01Ku7XgE
ycMwIdvMBFZopUKtSLqGv3QHgnLagVpxdpMtauZAqatoZ41JFQj4hEWXKvo6Ioy0
V/PrdpmONJeuji3CuLXno4m4OAg8KBFn2In5Zk0zTY7cxYjn8+rAI1sTZ/9LBbEF
Si/a+pfgzcfO+cY/FZaKTbAnYTR1NO6k5Ssl1A10QFjRen78xR4vqNLYW5KYRV2C
8Vb/Y7wFJErsPQ5MEb1W0zwTnrH83L4B8nqYSMFXfLR9tLil9Ayt1so3skI14O95
eE7WNcUhZ+/7yboARppx4ADJEONrgnhFYCwdIrXEk8igIJKKwfI63rwfQugpOkFu
UabkOugBDvmmKm9i/vnTz0RZOiAPx9XqYZHZ1yqWXHg94JeMqouFjtcqzifAY2Pf
4pC1oV7Z+fI77yLnQWk8Xpf3LF7ZCxf/1WThslXa/vMmUPfXoTI43TRCiPlLFAi6
LodHFBbl7vhv32yvByKZlwEQa0EAnktW1vy0bu0ySXMMd8OlNUbP81VEqre1y2+7
ZE8Q52A2sSUqzW2rOfizXTHGFhO4SbaHz5HU6yPYTXLTJ3NpJHfTP7qrjjpvrTq3
5xcjYDKatt5NILcGst+BrhDN57iTL7fit0jCYHVzP3o8Xs16h9td3HNwRnGRQbpy
Zxvw+T5AnNrgKnO5gg9XPGnPOKHxHhrSXAothHgeinHgAmax0Do/fz0m6d4dWf1G
qp4T0Wie1fd41C8lPO0AkMMI9U58/bH6zu0LdiNQRas+ArdO1HR1ZDfd+PBvvyW/
bdSCl3fF+6i5AQOokchngAM3TUhwSQCyOvvY6nubsc2265n8WC4bnR6jAAJ91e1j
IABRvULKsZRLuqfPT/Wu7l6PetnZ3E0Trj9K2G6gvKfGaNybpTySNC1S34N5641S
rWq874pYv1OvstXcXroHwMxKiBTipHtIVHX5inDgd7nv4WgKTuoTjq2neSPN/yi6
eIgnBdx6G4QzQ6hYMoQAdh/L9hKq+vyGEkL72FOHedu9GPhZORkd2A8wEaC59pRX
wUcPV2vJku6CAVYhxYijC5amP58n8Mf6D0/dPyn3Im9caSJZmBSH1N+QpRcTOhZd
fUKWH3fHufkdYcQEzdlT2Hym8MwCwiz86G9uLX7NwDYZYVJSl6Dxct1nxSRksDWf
lnZ5kTMhzXi3hR2nbMpNsSrDqNrJYUh4CUdMmNFcZxPHBPu0+8Jdz5GV0R7U0mjG
hOxsI8OJJDG4x12goYs7jMdWvLq9pNj5qjXilaObqfj0oSxYSx+irBwFtmCkTzn1
K2mMqDzwVjrN60YSXh7pBpcIkmdP3kAMiGBy5GNCUZgKByi4L6qYKzpLbDFnx91r
ZGc+VuchlaqWcu762b6M1UqD/rIkk2+sUAYNr6SvSLwrtZ5dCG+g9+tW9SLtGR7a
3oJiJRmh612pkPI4T35vnxxRKZzI0BRYXu2KfbwQOSJZLKloCtRMd8CPMSjxnnuh
rhTcJ5+PJo6ooVMNjOCVgmOLckeHsRXtml3U4ozjJM7hfCyTJu2FrZuxDzLlLv/u
73wnZPAUZyNojqSQlmb1/HFW5skJ2qPc+z+L0HpsqRsIQrYpkBvP20IJtJWmx1F+
U5AY/QwBEMTuDE0IQFLvSW3bJwAVJOsoxSEdJRP14rMBURWlwykVi0SGb6wx8B1w
1D0tBetgvJQoXlj2LgBVI0cBmhoabDQILTpu8XsO+Hm5WKkuBo41OmQyQcOaSrnP
uZXbeb8I82pm4jXZL3PB+AdG6onj+sVqWYqR5CW2KnZR2wAWkp/RsGyDcvWWWVKi
SJK1s/MT879qUjOOgt2ha+3d/x8SsgjORJ1YRWtz4k49WyyQNAmwnLkyoyYb8dyV
0G6SY4trbqO5ztSys2cQ2r3OGLsZqsucpu9tXgCoETnby2uTB5CyoTDRoClXfLPt
gEK/kBn8vHLyzvr/S47RiPxoW8D24zgmRRPDfiEDhaxjzIycvoalv0unE4EwDASD
IdiOCDT3za72LYJ0r/GGylh10qPFiVM4WK4IxQ7m4qRfRUlcLTJPagAdaRqBMzAC
vWBq/P3rkT1pFgMTZ9Awu+cUn1bz+/NH/VP1mNMpHzl+E1hQzBEWJDthHCJCpiT+
Ieib6VyFoL3A76CO/GEU5pGY7syI+tTNvIjR805n398weUd/rWdkELfD/htPxpkC
cirMC2kP01A4IWAlQ0IoHX9RD6p+m97IVhSlmIhgLcljhmN3ERBhjVdroBCZCLAq
8lDQk4nuJvJk7G1VghAl6r7rFv1XGjo8IVosxpc+rDvOQGNqLKhRyfnyRzj8iTBE
1FQfbpz1+10bCNuNQXqi+HPNNWnXzTOAKH4M3nwbJIxP0iRhZSxkDqRHmZMVO0Tr
J6cbVmY4p7zQqd+MtVc4sgKlkUaSi5MdWoOVtrMSRRu85eZWdDaVt6KobESWGigz
IaxIeN1JSN/fGt2miICu2e3NdQH+u1jMOjf21p6xz5dYwCt7/rukWLiSeREUyW7i
RcxZZ2QWGnuCeSz8INhc0m+e8+mVC8YBv2qOHizgttiMEUkkmKYm92igAmTXpLkV
aS3PmNIScrfG3Nau759sR1iuVoXGkeR3/SbxMGkqFFV7+DbTyyYS0N7Th5E01/zp
aM5bDvCStaMLRt+HEtDejcOPZZRB8to4joBDqZ9eaw/EZq+t6vuHkEygyt9ZG40S
DiqRTRXJxMq7/ld7nd/I6WFfHizTHPE6+ldB4ewkHfjFnLQLxy3S3uvObaSjiuB1
+CMIZMmCLODEiGT7CjJthMQmfNqglAS6YIpOyMj4u7NfYCjud1kQ5ecc/MERWAYU
uG8h4YV30rcP1tc7Cs0k9qY+npcOq02HQnqQX2NJxm/nGq1DqbTIn1Kl9XPnLusw
pNJFEIk+tV+e5TNRvYVY9xJGROsAyMwJDt9J0bDqlVC1/VquzvVYChbb6NsgdOjg
LLz09wha2Q29Bfqi1ATBzjG7YKzA6IlelAZHS96DsvlkptjZj9LCurT+gahtPPsZ
Xh5QC/YgUeoAmQbYhVgUNvZrGmS+ik+ss+okLXofeZzpQ178xGPf0v2SfKyBlDOe
MvYIW7MFzjdAPFeAWrFgwG9g0Q21DvHsa119C2Mr69/7lgoWkZgVMjs37CjGr1p8
suSHyy6AUqfoig24ceodEooN/EPedquwB7pGGZ2k8c5mwTMujqaU4hpsdv4pq33n
mLCzQs2eW1C00WroRZem4RuqZQwN90ITmZW12+dnR7VO+Av98d6D0AkqrbDN93Wp
/57VOfSlLgFx7XFWkCYjqd7GjbkTM0soVNyeZeZeO6usGWEIqUbwBQ3YvlUvYSbG
aojLPgaq4JtEu/FKcXnvdT6fOKHZi2f+epWR+/Z5AtemE8JLTKJUlmUFREPHe2WP
9F4gdi+i6TS4EgVh+E1fQnuxh0qvsB4lQdSOsCek6UT1ncRNZ2XwrULc39fw+dES
9yFlfNIS4URaDN3UlkWTTPrWsxXuWy1TYdkuQPWYNk6//n73jtc8Wc0xI/Ob6Wzv
F/FfkBvbsUVoilzvWTgmUl2XZJUw25OVJD1g0ZD/zy/NEiSeUCHprDPpI6h+0TqO
kZZRT/op+fHyKl1wVWXf5lPUn3wHXs7UERvxYWfpsoCGJMF+Gtyp+XXY+Ns2eE8+
JfH0jOR3l/zBy1dtR3IeGvAw/Qy9s8QC109PJWh7cH2ea/TG3L/Af6QqG54TaUd6
2zcjYgmQa3F0VfzIn6P572xWzYQmBsrlXoMqrqqUJAYygj9ofsQbCvBLiAuZaof6
iw6w3Zb2iP15WYUktnDgKZXgPMcTt62CVFMaDCutdHNPtaicayTEcukRTcMd3IM8
Rn9hTLqzXG25O6nAsYRQF84YB/75Jon9AAfJNQOSl7PCmBdquOrhboHEpIVA0WFb
nTrfu/ARlpCbSTZhKQxhIVk+4hd5AUDCUr8hhKAKhay6z4tgpTmbl2eQ6+mXGXc5
cfGKaPrIUaT1tNPKN8JaxtHY47Lutn9OwsuL1gwWZyMheu8c+Sgoakppw61kaAvF
ZP1et1kgV6Cvnz08J+QYukygqepYn3vXCXe5ZUy8PyygVJk4b7vcYyafo3gdyvzR
z4z+hIvcR8Q3nU0ZLe15w3hBBVp043TL0Etfh/m63z/dlICvJ5kjGG9/vaSDzSIw
QRYHa0tZikeCSozGpn3bWhvvD9PrNQEmhw2C+a+e5mIcV7/bwM0W9UXQ+n2z42oJ
8KrgcKFGOuT2jwXIsZtZXYd4g4DOyJmd0F+AyFe2km6PW6t2YjZ4BEFERyXbGqZm
4qfFWP0RSd6uwCMi/pyepu4E9xknnyk5HTjPiBDosramn6M6zY6FzwKMnPdUIpBb
imGMiDwjIgQtqrz7hQ6pwtnQwtWCkMIccEctB+FaX/I1HAAa5ZSz4RI4iUTrtsGf
ylqTM3f6m3YEM/79S1RFI2CIr/wd7vaNjNqM9KQ6hE2FEDy0oE3imTozDTOK0Ji0
vGSuxDXn4dRce/O/MR3cyyoptEzcz0c1yw4OJzRf3ybvwsZnu/N4nOq0xYdmjj/7
XYsT1Ac6+gzxcjp+/55tzmdIjj71icslLfj7QjPWdnjJYOnuYjryBMhjA0BoH4Yg
8ZAuR9sNy23LYV1FLCtlLHFXyduyECHpImsn0LlMaJXJy4S7G+MIfT/GuL5qF0Ip
iXBVQbYpV2OKyKF6Zh8QQlSs3vE0J87QnFw1b9ep0k1N5S0Pdzf/KqtCAumBxx1X
u3cpj0DWOPTHzjqOezYzif8w72vnJk99yUVjBm1CgmG4KGRUu3xEX4IJxokbEtv6
bLbSuUieZqMnoId5dhSfFNtSym7SSBKu/BZ9XSNEdgS7kofBanfowG+i6fjSvPx8
2LWkJNr8zfYrityhWeKuZ/EbrEVBDIbk1AHsB6J7R1HDJ0hSvvbNYAbJz72YPGWk
/W3HH5quOoBLaszE3g/V4Blm9C5oBm8PP1Jvz7uNiI9ri6GZdewIUGJkkkk8CoZw
`protect end_protected