`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1952 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
XDmUU01KuyTGZ0KfD/yCU+56Kg/rGyT/tvh1G6yhmTk8AaEUPoaJaNtOEyj6LZWj
xY2wIL9e0IB1rCG8OAawRN8+O5jXdFQ75PncSNmYEzGlNyg/dxfiRaNqm664liGV
2gpp73Y6u64aMWkTrnMCaw65nm8tizKk+/vrczmO1JkZjUv42uv19tCnXDVb7lr1
Y4CxCFFgRWiLXyrv50eghnq+L1phB+QRXx2ZLIitwsWiseEMlEYemRG6NkaaiAzD
ijp8dgJ/j/L61iY3wxefbWq3qZfsamrSj5xnqIapgld8zLY1goMIQSZXg8XAke6n
RiQYuxAGpWMo4Bh+VaPfseugZ0jL4os0sR++3Mw3gVXelKnBBL/FluLEwcj8/91i
H4c6vbhYMcutC64/aOYkcYMlNFEpfjYfFPYTShUAW6Ozguw20SZajmxZybxtFwX3
9wiIwXRSJO13FTfulkg8cUytyQyd/bxJRdha4QTfnwbMTxrrPeuDZOtlmxeyAi65
AVM1uK/G4ZVIKydYD8S+Gcpswkt1TxY7VC6h2MiSaRk/1Y+ToUG9BHhxC79gxMG2
9XWFMLKck7l3tyzPuMkbEIyyU7TLCLNMtQIYnKF7eBcqf3SzF8NZFMUI5FG+KUXL
5oFx9QbBfIq9iPsVg8qKX7y5JYr6sj2iAhOkbNGmeUGLEpT0p+YzS6wM6ZltA0N4
5gtnaZ3khrXuxm4osSYF9FqIkarm1Fd4Zz/HDhrMwFfFlxzksLuqUYLhMBLurY8S
q9bcQBw/ByCHUlcm0DFnD8tyxOjxcxR94tvXqAUqSJlQZBkvxrEo2O2zCsKZaAox
S/kLXt6aNEZn8JykvfXwFjoBz2UL/HUWtgyF8ifvhpFGtBXENoW4LfwG0IWU1xgK
2uT9uB2/wx1ZvB1H2TB+rCc9dQDoLTOKzI6/Fn+8UVG/XcrJ5xMG5py4V4gPUxVn
6KiKwvRxvsFJfuRG4+1dXoVcyiBzKCaQTZKq2R+geoqkbVsF9oe+VyhOotfbLVGa
MP7Kze/FSjWLJVXy0oF1MLMh7wEOYCbflYTRkwc/9h8fKptyp1ttgkI9R3n0kihW
HoUYGAI4q79HG6dO6IH5SLsr5rtMtNvZF/h42kaXhiPV6aTnSIgWQEVOenEwI9AV
7hsb/uhasaw2UxwmkvUR2Nz4VwgmSlWR5hEHzvW/4wCO2KrYTjrvJ/Fn12OizbnM
DejvMP9RB7Q6XHoIM6qljFeTxvO2sjcLJmY3o/zsoR1Qlig+lmt8Sa1GmWi78WRA
FB2Y5BzWb5z00TremEZgAPzI6MnTeVfkP+feUh1sTe7ewpkquFJaKPXM0Ngtitl1
cm0A54qm8G/+Ew22Y7+gHGTNsDcauR9ZlsZz5bSubZzjqY0ypeVk7fKGNa7cv7Kl
aOBqwcJjxeIAhoITu7XKO+dyFOjBo6XU7caW26pd1GKCxKMy0w86RI0wK43CwRN4
eb05Ugb7KcUflS7o5yVnfDHeTDGeKbYl4RNI6qOSdSNpTfW4ESjHt4CpP2zwF45S
o0ZZEK5wqwO6G4QKNGF7ljABy1hAnVLq/3tTqLLLC4sBU7J05w3aOuwH+snR33U5
MFxzoxNjZ8FMkplcmtiRbX0hLMRCrbhF1exTEP5hCQe8zuQnMH+zuxyMNXlvSP67
nEZFkV64bWBIor1YXumabfjfbh0VyisBVvF+qMxJZW480oEs3Q2EwUQaGdbX8nUC
TWUylss2C6/L1K5DVtHM950FW229AT7N78LtwQ+a6YUmIpJYl+lzy1qGwSvLYvOX
xISL1BBS+g87oYbZQ8+/714WbvTTnX+E/45dbEOIrG4dfzHESDmVuTzZnXa8Ypr5
9M9vLb0/gkIs9snAk/x/ziWJFPz0Jom5Zz7nkTa4uld/1uPaeTN1+0dUb0RNzIuy
3mmH/yF3xjIXdx1gs0twEUZwfy597XWYKNciJaTL0m0vJkqYC0TndTd+Ytqrbg/G
26Pn2N3n0HGUS01oKGzOi+K1zeQQeE7uDO+CJ5u1ZmHoFciTK5G2pKzQOXhtAxZE
yz+9vLG1fhG5nuy+kRbBt8R/nyYyDN/08hf14P5r5O6AOCOeQUMCHW1Dx5vCWA7l
i86OtY6RXhE+7Ds/5+rFLleW6jO78r5zHHBlZgzxxZhJsoH1EUD2nd8iIAKIeso/
Zx/UYEkSUXfIGhm0dhWajyM6hmh7MPpnLC1X/FN/uk4jifGmpiqytIPPmKoXUyir
4qfdI0/fjsJOpenn+4pvY1NONlthPsPRHQdn0WrAVeM/SWGUyvbhumXdWdZ5feGQ
Hq61dnHUV2lMS5ryot+/kLXhgjbNV7D4KqlF39GZPLPMTeUmiaUuzl+LWikSvEyL
NzQLZ6E2E04SPunhclBfMjnbafSjtvnXKK1j0+5HIDxtKVwLO80AQAWVcIFs/uVx
ndSoDrQHYkxwf2gPhGOfBoo73umzOGtfvqISUF8goMI=
`protect end_protected