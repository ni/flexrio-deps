`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
j9eMmSPGcKCWAR9PvkqZ1R001FU8QKTyJzFqNLn+qur6INyYDE1AI8LWcxAzfnTc
IpZG7ua3uuk5/kQKKQx8ZIPLfmv6H3t3eWjki8YIAtY/d5E7Gq8Z5mNxMYRzGGTg
TCMm6oOrOTVYlCXHE0X9AW696Z7UGfWirVibl8hs19hrFdeZKGiGht4r09vHR+Gl
FQQmSObM5aSK5wu5KOrK5ZUKGHyBhjnIQO5NnittDjOwxV/57nHVg0pdG6JUqyvm
tEgmCY36RCMRGWN7sekPtNHjqpZkmYrVX1T9QF3h73+8ZekZYd2xY2hpHHGYYeWA
t3+Fmb/6NUmoP8+Pt2hI6g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="wX+NBVcG/A5ruHK3pkDqG8ZVPdOz9TJPJ5saXZYSeQ4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
j/hqWUoxjK88VtH4QmjIrexFOSwtsLKOZ/LCP4cmrqgzmR/e71apdtoL+o8nlfy6
eZxDZMmrZmJGoazz2oK6kz7xJU85UCwNc4cxAsVxNdCP19vZxph/nCYZQ9lUFkLH
uLBkOeFP15CD3jG5/dp945fHP13J9SzB/L9PWvDC/gY=
`protect rights_digest_method = "sha256"
`protect end_toolblock="sqDZkaglKf+bDjC7VKm3lOELrT2Jlynh4UhPg2J0Q70="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
f9kZDbPp4NLiAOFOgATj9W35i3s4a7wbt9jeHjHVcJxMoXY8rb8laqS5bNUhXGW/
MOc7UNc1VwolqhkS7G27SLamkGClZZtXSbRcN1N+5kZpEaBEj1343vVznnU2Dre/
bKlbmouB09/BfSaq9uUVg27ZN5X13uRhftg52zTbjyCmi+BN5qjrnDo/1OCtsjsy
6VsfonBTv1MJpIIW0NCrY9ab8JUfXBlTk+sIwdZJKyaGwCaFunV4IhvCyz77l4xA
9aF5MMTyUhvVHrW5rCOJIs1BruoktmUhIWmIOuqIlqAqQyN5ph5zZ+GozOE+naJm
UTcr9kbeAd9LqDlFXNI7Rx3EaAItMFlHDQH23KrLSYAF59pGMKhbcF47UqNVjcBu
W9nCg3xDn/dXdRGwJzCS/VVyfgsYkYs+pF0t2JxRK1b/zYRpUwDgVfbexOD9ddas
lTsj6wGvcKy6XvYj0GgClSJMuPcM8Og67KlqGMA1vwzXh/3LGLfcTjJR70VvA3LE
/pAI9oV1rrHFffidMgpJzHhh71OoeDFwtJWZj+E3p4jRA2sUCZJYK+ip4SyjTTVa
iAyd+hN045nZs2QnmZaa6/LWiSvZC0Hp3o5U1nZDsAryZd48MdCy3fr8vrM1Tatl
+QFVpBqerg+IUuhv14qjsmawxt+d6lzBuO1vaqRrpkz3Rcd2vv7bOH9g+iMj4cG6
JkDFjOQp4sDichgcUynhoYu7nJWiOvqzvghhmqHIyaTQanVRjkwr9rIYsb2OOX86
eQo7pNMrNzx41VGKSNXSmqgN0ctAgkOtgXfQ+H+s/O4242ZECfh7gag9TBpTZEar
IyqCj9wIsLJRqnhRhJWKHuiXO2u1ZxWe9FBalz9/9BmYgOV3EO5IxsEP3aXHOwR1
Pq7dpvucovOq473cYO41yvAanimuFHROVDlx6JzzkgJWo5YuhT+oXHQ9oNh8OVmF
36cZzhrKfB9E9dU4URaEhoa1FqAJ7okuy4WKpCoGyq2Qzh+GI0fkdaMaQTTSpriX
BNcaqU6JPmRXww38uKGxlfm53/Ln7LflsyrPHmqum8PnS/n0Q4arUdMtBTVrarir
0J88T0fYRKD6bDZjPOcGv1niXvOMx+dL0H+PfhHkUeRTOdnhdW5KqpFwOeIegTFd
5gfsJeGTtDmI7veXblLd7CkDK9o/zyCYw3s8iGa+B2LTx4M2xfbxhr5c3/FMGKTt
VyuFMHukKnFnePDM+3NDQ9SoUiitKxENWh3ryPj23zRXCYZ3SvvQUB95ZRubXQzW
l99nkrngLyswwZVS32HRIBa/cZZoGkF8PuiBXl1cfMmy1vfwioGGrEqtISlDQWvt
SqqFBGsRunkjSnj2URqFk4mTtj5YHS77YdxWBioIOVap+bnLH0VwLLKh9lRGX17e
vVWOf9kdJervt8MEHgBy3byArp3vVCzqWG1QX4pnGJhT9GOoi6Ea6zz6JqqnqULW
uKgM4nADe7RyFCwGWV+3gfF0B9zot54vJ6DwaWS5CfCPMDHkXSCqqqwmKROUog2l
+NLUlMlwmKOxWVLg05wpgeJZQtFBsWWnnApuptPzMqs0G0Dzj7OCDqn67p4XCqwn
Rskk98mt7y/+jKVZ0dNb+rqibzxzJ7uj02m/yp2EEvvuxkRXJEWRm3SM20FZ5B3T
u1tVVVCTiTPTZ37NpUPdpqcG/btir5spsA3ex3OdvUQtgZD9slQu7yJTWCUQvP8t
uYsWvrT/MharAjBeyFdUCYIhQJZNdwWkPesBhsDQmRJWPHv/Yc0RhOz/gcGxz4dW
5oKqplZSFmnD1zQN9LrmBCeVJEeijbW8D5DxkWojvooSudXnX0HIWlIWABTFX0zM
ecpuHSenE/dfjAvIGxGGA2NHNKxj3WCXVMOYxsNB3InL2wNp4DNrdkggHzFAxVen
wn6BGTl4yskSZOnqIzUk5QCrLXcS3YVTQT2gLTTvtPYpNwrlGz+/q7JfdAd3Ea8M
LnhAIV108ZGxOFwNrWIeMKP79AOv4hys00fMr0eL0d2CgZQIz1YeFCt0iCqpEYig
dZ09IbVb5qHb/bmNCHArNTiO0o7zG2KyGR4lZUZvD75+FX9rAGHwxacK5Qhx94di
0fDYuu7ql4INqLwNN9QFifIWLqSbpYkd+akjo38wRsznygJgxHLGzceod7kMqZsv
ExiKwkN4XRXBu4MRr/XLItjBRLB8zvcBrWsS8n889V8z8gmOLmYZP0sJo2EMDexk
8dEEj7YJ8c6tYUZywernoLOG8jKPrIibNYytH072gV6zMieYKwglypMt+YNP/n9X
Cqlt5sdiOiSLIEhO2E+eYO8SFoEEyRhxcN33dSerjzsfuTIsjBycpSLBYHnv1KCS
sbawjNQxghH+L5EDuvlQKvXlj7X9uk1J583Yzqw7VKVUtiayifDrPFEXVZhWed0F
y5/4zxlLzfFvld0BeAgdoik85ot9L/Bfj+zD894IYslaLnnOG+1etZHO1L/C2e+M
69lMs6kPFHPyv37q0qpmRcJVJlHHk+HDEVlk4F8xzvoUzj1POqbzKewJQfEtHAm4
enVIkJbREZ38QNuqMYlTzGwt0sFX+qHoe9vc7x9XIFyDbz/7iHpruck9ZrU6Eyqx
QBeBSxffq9mFplxsOx1nLvsnMEMoE0E4pe7CkEI0cOtSkD7XjEUrYV2eVpsvXTer
`protect end_protected