`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1456 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
oDqealYugrOC+OIsTtIIFHfAp/+IR7cKlGJbRRt0fryLNHvnRtq4J0HUX60vIm2c
clNEq4FxExA9CeAgDdrQyjLkfohxKablXvyxycwljsfDuDZwn1ya5OyCo1mY2+56
mv6nuqySxJyAfXKjaYF1vi8zpyceFQmufABeE9NMMoPM5nE6sSXvr3j1MEELtkvr
mYyQTUjLE3ZlBjqeJ67GVln+j4wIwfJzERyLHXElao+O2sLDOlOfzqRHvKNxr4TF
geYofpM3yr1O9+TVkIFZwcxfZ3us7dvhuiuMG8HzCZg/u3PdHftjMRtHivj+k1zx
ot4x3ezFwm/GlB/h+QsCzFtNHWfSmkh/foy39RIlf7fMz8dF+DEuUHaGF6FqrEyw
J2Xv8ZivQCxh+dOqobpGyAlDrGhlIi+e/oQQaHORC+8MH6k6LsfBp4iUWMcppwgY
RbVW399B36Un99Wzb0+sMqsCZnF//HZ9Agdx57Vk40eFZCaDUEhn2pnLgDT1sCfF
qYWWVKbyiw4ot70V7AaHo8k4a0MhVSci+3AaAW4YDbwBGsu6fA16aXstgTsf0Q6J
4hfEykO+MeVmMDh9UA8AGvMPNZrudjIpnor1bhEik5x5jvtBstzxxE+Z20AMJOuB
/3bl6dwND2g/cP36kaw+JuQnnaO58g8Ma/9wLybYEGBlzFnFudfJjeyxP1Oji3+O
FstKKoIDdXkxX4FZViX7lAslcDmFLjYsRIvTuHm1WC+KFuWhY4qlUGnVOl01Ibbs
yuAI9PT8F9quLAvwzDqKlIJOYrn88xB4Qdf7fYj177KmESqsR5DOrT0sYNbCdnw7
CHWKhRPQTHn5J4sPI98Aat+RxSaEyJdNsGy6fmx1UFuDR2IVYlNGRC1HiumFf+vf
IWYAkUB7DrEyVdQOZ8c80xl5crALbGPoex4WraeHTF7BrrxKjgkdq2C2841p3u0p
j+rLN1jJKYtNgX+/QtwwJKs7L5nJVMo6t1ET2RtiPjxMgvBdNyUzYB5hr2WsEIfB
/a7WdgYQiZEfzoD2JEOmh/xIrkTQ5AlpkTJ+wQXxGv3aMiN3fybcZO1RNHHs7UHA
S3KfkqdzL8MW/1NkBz6tWsQKtkDAGMW7cLrsNNvKhmlZBsdEfJcxJn95s39B5H3h
81U2zulJntu6U6P70q+LCcSVsavfbVf+bOf4WjGu2dPA7lPr1sCPOAG822vY7Sl0
fSnljPgkDDvlKml9df1SfLxSsbgRidf2SbnMeKtSAUzyt4RxGruE/KJRzQRJa26I
MVq53jBK6JRc3g3fzJmmJ+7KIzDk++uA2rEqHRZP+Lguao5EFM+OIWZPGv5QEqaH
rZx+MD8YJEDX1vEwZ/qlVoCGPdtrzXlG7yOmn26YpCvxMHfDteM0N9Ko5mbnIu5y
YTcQ/enYhRf48ggEA0yGjH/UMkYDNI/tQPl9GttI/lcgRcR6dM80iTys6osHrZAn
Trcku7SnibVqAaavFNoSA0hxCFqTo/qBf9CSCeuQSXFZw/RMstauDKtk6uBf4plw
CDZGnrl5nw3U9bIIQ5l/L0I48zG40Fpk+Ftnam3nWums6tAJMIHcGeuld6atmSuM
9RTYoqKc0bu7NmX4vYST4WMjUwD497NSHenZTZhc8mrALCyANJq8OeLjpw2FGqS5
sHvI5YzlVbVtN11jfWylTootBu5qipv28xdhjCEEZ6Ni2RFO+w9fDyLU/cBGMI42
XWoG6EpFOiSuKcwON1eDXi0U+igOX1NXGa2CHwqJS9Mhe0u7whvKeVdAH/xjCJiI
/Aj85t6HdouoISrRom2rWg==
`protect end_protected