`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Jm2uGAVYfY7w9Y5qKstopObZuZAEY3b/Io3MSEcWLhjjnKulVhCBBYAEQrAzzGsT
vMbffkdZgjdXQUg8jOLJXSHZ0Dgbnob2vlppjZs3bgyHCF7MoJ35E+LOsaLimUA7
hlqStcK49hR1hdeBPr/OwfT3UeVrRtQyq0eJXQ1UksinX1G9Pz3/CmcGfTZ/C72x
p9icpt0bkY4/1I4GBvNCsA6FFKH947JqH27OPACiQQRW/K7JToQn+1uhWr3LA1od
lbVrWu8PdZi7zW9gK3jiW5GaPjwbYQGqeGFs3bTKBILjb7sYHxfxw7eDLVMAIu5D
W+OTIN4JiHiE1gCnNEvkSQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="pm+c2fYA/4JT1uhlJGVUubML8hZi8lME4xPobg/m8uM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
nBaXksR//iZ9fraC7WMJWWSrjqRXHxmM1Y0+KKN3b10NElDzVNMlR76DLrcnamFd
2n7uzsxWqhhJR5LBl98SXO3Y90J6BMbw+OBG/MFM/zUulxh2Si5YK5G9GCrG9gvZ
5JomxuZFDu9CzlWGTuRUt6FsE4Lr6sOL1P+hraQDpMk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="M8TXDiNa0BVMX1P60yIvW2WA9jKGGy8GtbuPknDnC9I="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 33072 )
`protect data_block
/5TNZvs8Nu0G+mfp7M8H+iVAGG3Mh5DYZ0Gn3rRNhV8b5CcJKgjQajrRoGl/gSxp
rBAhtT8Vd5eelHgtvBjpvFBA/EBUrRH6CG6pqRt9r2qUDt4UernbZbxC3BC14KYF
+nUFsqc9K1YQwskh0vG3u3RJluVXu7h9yhJ7g3NYsOLcTm6GtYXo3b1jSwa3CJ1l
VBdvLpvRwRR5ozoEqVhJ7n6mMOuP79PeM+69v1cybJSY8FPFDvFGzvXiVQHN7YM9
FlKc3Z0wUNCGsH1BigzyY06r/NhemFBALaujeGPT8q9KA7kk7MCye6vYVgHe0vNi
UygngLzQDoo3wL0y7Tx0TDJyd87HInZzYz4ZGhMpY1W0lEzuiekY4vUKmqTPmW0k
FIAmz89FGEOcQpvyr0uFHEDM6J+pB9wJvWAGOIUHaX6FgyUg7klrZ2upMz1rWXRo
0H2bYE7VLYyoA4GX2dknANgiczQb/lwDYq+jH7gqFjb/PPeE71BPoCYY5xJMibRA
zNMXEWXTeNahoRCe1a33gmzlkHcjw5XjSCvo0lDG514WFXByuG48hy4OUoksLc69
k8WOleMfh1fRhTJz9dfPxMahf43AVGbP+hgcjiyTB7uBAP0QnHESkweNsfaxb6u/
716j+76TsH/0a0ju3sT+7z1W7Q/hdI5zk2mc6RcVYsGVkvPKtItIMHmGeNWF+Sex
km0M241QTCXoVRn7XTCF/45tbZIctHW7Dmt3TS9W6LWL8RLMvXW/f9WHTeND2mfk
/zB/trdWEHgxLFbHDAjozA25r/QtF9VKTKppd2MwsjGBCqcHHSMU55BHme1gwYG0
VfPFMjV+umvTGm3Gwr1DeJ09AdiNUnJqJq8w+PnavMfuH2jP9Ah268g7gDVIK6ip
2vFF69wkTEWe3mNBbf3N9WN+iQuhWNlX67uHKNqtA6YtGAjaBr2EaZU98VvW9QHa
vmCDjGH45a39WQCaFjXq7UWEcCrYJ8WoQCQJ1CesXGDYIbZB6tCEM59MzhNVKHKx
db79pVDyHv6TO/PsvLeJOaAF4UibqMffQODJ5zMQFrcBxYoUPoFxEUoHjSstgwgO
iNV7CTrTV1cNIQmppmkZG+Oq6Qzzcr4nDyu7nNjEG7DmwNG0Vu3CQeAgq8hi6Pde
3VeU1R45+n6icu+bTT+VFuyOz5uFS3UQ6UKM7JjFz8tNBBSy7f+p8/AShbresZ24
LGhep//B3GQkZT4dUwEKcxjqlc6VhTDB8vQVmwGmUMNy791QtmHQJF3S1ixXim1u
oLeFm1Sn+v9OOhjRslCMYSSS9j2sLY6UtFSl4w/28BZ32KLSId8PAbeDgfIbOpoR
gzIFJfXi3yMsWGPTAuSK+oVQnObiRjY/x6K+YnJzn31eOJICl9bPC10KUzFpoOAP
1vFWl5eiP0GBWXP/eNWl+uaBSwQUcrZxFIgBbUtEFGluIKLOzP1fVy6lfD7DMJ6r
8w1ov+4Hxgp8cQlOE6QlTJWXlxnXnMbdpIc5hFWstdTo4/C42Ey8td4/fThLDHHO
tAplNBIkmNpz/9Cxo/XpJT9JYe9EoG/qrl/E5dWQVSVLe7fYOZ7PJmtdloW2Cv0h
SOUhqbrg2KldthAmbuaiLdiIVnrqIjdMNfYLKkVySUwoNXvbfeiWHg8iUXR6pC4f
GMJcH4nGoxIkHXneMJYavdRRZHGNW17evqOgXo5ZeAneoUENaPlLwhsrFUD5fz9o
peSlIodX46bJ1DIF7d+wsgIvGjXiT7Xyt4y0CQs5a20YrSEEeqsiL6g8V0bKbSTI
FyHmTY8RHXEke5LrVwVfmO/GSL/MYhUANDnPC3hYUSh5Hm6vyqVz9qyeelGlqHKC
Qcgaov+pQ5cfFknL2pqYY7mObk2VpDY9XWDVKllosJ/o0MFlcFnlml0+9dGh3yPF
rthB6WXl2iMi2kQ/jWvC76y0cEdgRp8J+/saIlVlmQoOc+Se9SEVvjuVfL9OerNk
bM6eFAvRlpW3UggAjGT7bKYxBF+TSTeOnsHffvfxFU4YiOC92tbu0fNbwX5FsCen
HHiOOcuEaHJKPrMXLKI7Y8w9wdbXo3MCmZNjKEIpqRrxmqT+CXbYPz9Iuv08Zcng
5uqO62CzWl1aMvhTThbHOrf9rMYt+gOfnFVClsIPq7XA1V+xsI3c06iqkY+6LA1p
1W8Ttw3lgbaU3ZBGvML17AkHF5p78wygmtR09N9EKg7uP+P3+gUeZtlDYupDyEsW
RT14Zz8GNc8IgV+fKllHSUiZ/mpcGa//eNeM1LHHHQs7UHQ/zWdQaxbfXhKFdSvE
dei23Zi9IL28hk6i1EwmP7do6MTmDHPSxONj6tDAjmn64PADXlQnocHjWyKSAjl6
DEy+uEiZM2MQMPVPcMFSVCo3dl6avqG4JcMsuP92JYrke8vY90X+WZ5ilut7ypH2
oRk4deU1R+EAQxnowSvzLLa0LTpXrVZyVvRYhK/y42hZwlLjRwJW+m3Fi7xrMXvt
8K5slhSS3oZ+zQg0mph5euBJQWd+viPwHNgu5GGQ/kcvoVqOn1IgSirAC/a35sdF
3qOjp/zLlziFalJIrs69rBfSKGtUgUfjZxKECXpi8STAS5Z88ozkhJ4Vd0WMcHI8
KILfoB+AnwgAj7HE9WwF0WwBlDWB6uIPygnzVcG5Olt+WVKTbGzMFxabo4lVbWLT
FLfFjXM/79wG+FCMg5zjJxYyG3/WYzLIeUSOs9I3NXlYTcK6iC4PGxH0wEeNkvmm
WOl0zn81M+vpH+T1vAY2i6LlmPa2vnOLMkeIAzm6hV6rKmf4smSQzJbZlMGDXcqq
2+lh2mq8ZLzqqGeA4//OqriUMI+tXudVH/4mTl52XAIXJaFgF1Ss0AK9SybjXuZp
S/T7KnP0+syXMo0OAp36FLUGhGGzFCxnyDY9j8ay71bm1lK8xQatRQ59x+3cQvGJ
coC6EQQE0Qu7/w2n1nmOYgCHS16gzvvuXswIZiaUWjmDIHi3KQ5L+7i15N9k5kSJ
cVTv5YFF1w/7lJf5C4AdBr+/elB6IjsJEF5gux6TgP/aUUO3sR1fmhWBB2CzdH0Y
fsRLQza0uSzPWPL42skBNME5j/gFqEhS2ccsNQk2OccQOeU2WfW16RB55xhrGOKn
MeL14tgtfS9WN40Q3Zir++bAx4ALGmN8tg4GWWClMJSZvgbdWa1F2xOogfiuowYh
Qp3g3n8zR0tXhKSOaMpe//nxlYUYkB2CczemI0PDSv9i3iWpCQBM9G7BRZrdIonI
sdCo4vZje4spsuo1J2IpQfOiUTU3U4Ic6ywuM5sKFHV4d0+PkzjZjEZkXtLDFRyP
k4ksyDaNogbQMDKOrs6amGCjrkwOInpCE4ysYGRfF+sSJ02mah6npifQju1APQwH
EHDSp40D+ZVzMobqtauv1RPszPkRa1G3uyroF1aiCGwXoSUFhqOIiatXNQzMTSm9
do5E3BlZW4GRCNb8UB38m56BtGb5xwDqsja7DVXZckJk+VSEfB2W9l9DpU1INsXL
7WXJsJaVXnvwhOMIlHA0Z0G0x1ufsAIRPeeog+wP0xuqHIFp8W/2fjsP5LIHQfR+
+ky9dtfGGUKeAe1oU9NmW3x9HZ9WOkTXsoP4L/sSSBzJgZD23Rnrnmo5OUG0FYhK
ZmI82KbE7hWR4h/n2QEkuTUZ7uEHqRJi/TnGWes2X9rG4soNeD1fdWu3YC/ta5Wp
a0cvLm6bSGaSGjJMbBCIi3KVlGTNn1pDT+hNA6CnRjDjm/IoOsBFCYkQ9nKHzpvh
VNTNXoP56VwweyS3Ne7HnNJlYa2vPZZrwM9k5VZERSsC9MSEPU+LgfukN11cYziJ
2LbQ2/bP4Op34pNLne9xjtQGTifq6c0M98PQruuGRcO54L1tOHe7j3DpL6s1SMw3
p9U5hEyaiFZwwIld0h8i2qaJKZXeATtHooEuyGieCMTMqOO+7rMG5/Dvv3gPYKbE
ZWJCSL9CKfsOWGvfyLfZ837W0dxz3TyK5wbPXH4NLOEVfIaYZHW0t6CFWhnJg7bS
MnqovM7JR+klVQPwJKnw3ifprnPQy6ao1/RoCO+acpUdofPYZZcu3xCOcQ7lP4Ke
aBSf1Lva8pxhgDKXgpiLpH2bagRZbNFXHfmsVFbK8ZMITHBfzPtm4pjl0TkS31fJ
abrOBJ8Dux11nB33kRxyc2jF6sNnLG6v+jUlY2wokBt8e5V/dGxq3f874dZ38hK/
nbIOdlONI79JHlUq5/kBreO2wGRqaSjL3LDSATKfqSSxnV57taMPocpupiLXqD4H
rNV1DjT5Zjw0PQWLnlmm+3gd/nZ1+pD7Cyrxki7snnSK9lFWoG70lJM3VRMdbnx8
6ZQR6nyoM6Qb6pznbtZp8XuudbqJEQ1INvP9lqx4lJCm7CmwadLn6PRrY8Bfsa22
0VrjwKxIleBYSkWcJXbXc7Fp6reDsGMEdJ5W2/Lzj6hSNZqYzKTi519eLSIsowA5
nAsCzB1sZAJGfBahMEPt2kFFOHy9revjVgyCZN9q/8P+bOi9oT6tjPnHefF4eFpp
tLsPZOmyjX2/NjB+8dqX94+dLvcYOAcC9OJYYSHBrvxpe68xplHlzQvNM6XXtXOL
KtjOHlFuj5YZ09SeY/tOs9uA8iqLmb2ZSTH01OVqiBiRPrGnx6KPgPHP6VkQLIpR
2qlQHEls/yuXttZCA1ceSyzigiy5wC7VRo54O76XgnOw5A0JhkseEY/pyr1mlwAJ
5xP8CplmWQwWcPq/h1lpTp+5bKbvsmJIyTV6n2+X+UpgiSCxBYayb1r+CRLv7KS3
rQD3GlQyreQKZ06kd2IkDRwBVzi6KR8P1daTzJ2OsBZ3/0aJoYJ1Jyh8lwNoUpB3
GnNgG1CRIk9PZYNdyh5OPz2ZKs038q9l+pHCwZ+wk0IERumCw1jHXacqPEq9PSTI
pnMRQmfnkGxgduaYl2DO5pX8mZr33zLMeBT9cLxxFJ+Wu0yrekGGRCl4KS4A+KNQ
CwpNN4uXx0bVN5BfgSXaNqTvzwwk9+nXERYfK3YpxSbdzjjeIjxD0Ywh5hLn8O3F
FW8gyLSeZ+zU+Y+XuupdVV4PgWKt+vCoVttLsejEiSslhWXuFh5xo4Wc3EMmQuFi
Py4U20yCyKXCSG7KCX0CjVgrFFnZKsw7JONhQY/DBjW+0qbmgsFEvqJ+t1cqZL94
5oOosOx88XHCBI3ZBnodptIxBaqHutFxyFn11Uy8MbXMeTS0xNpKyEbMX/EVOIT1
v8o35KGiUsHaiLS3TyaGOrDs0MJnQxbL3sSQp8wC3ENLt6EcSnJX8jEk+MqjhWl1
w+6MwSXKpM3cYuyozlzmJkk/k+aMxs9t36qr2EqH6MPHsG40aL4H9TZSQjNYf9mm
HV5Ep8lGTFfgMKG2OLktLodw2CDlOS/pk3SIUHrsDGTF/6K3vbiLjW30Kco+J2+C
UlkCa9NEBu8CokTo6kgvfP65pLrweGsZ7QaUAN0wlIGm9WZnPPwG4AaN3SLAbUzj
z3g/4E4foKwvR9dfe+7c7pbacnu7lUfxplHrKqu3utt5/v8eZzSd4WbJenchG21L
L0QfNcA/CFntXlJGmggN+S0Muav26V03vJ6B+kHPMR4Six09VTHlKqqDfnHDXFTS
8DjVapF0rTup6RteOF841eJ5B35ufoIobTGbeIxBt2XOBau75SLhkf90WLttkREP
luouy4k88srLGhGM5I8Omvx34+3gk1hPuoN4jJFe23QqJOuOx/QAwlDNB7EnNe1Y
lwbNm8Iqb9HcD9Ml8v+87jziCMSw8SS1tt5Wex6U0AB6NEf/fBZxi19MJUtuRSu1
KzYe8o0v48n+laZLA2Q+cGzg+J/ctJfGN5E+Pd9yZRVasYFSJF9P4gvgsebZhRiV
4XsiBeAs+oQxAmuTj+kFu81Szn2MJ2hJRy2rWjtcitlQ0yHOZlo3bOp1/2ZXvPYO
HDPqKncrTRcVH5hs1Sx94smK6y5pQsd2/wszPlEdI+hhK9dDA+SRTyFDyhBS5l0J
fyz27nh51re4M8jR6YYZOHwMSyKyposqBVLzeiCxYTfLX/6e0mFaO/IS57k3nDfO
8TMcrpnFJegpP139/qG9NxRQZ+ad+NZT7meDVosOzIpDQp9CQfPasetwVFoBQiQT
/jEq3yB1jKCNm+9E3vmJlGS26EawJTb3l6BmF4qBzKPGiWqpLVr1fagvwdip3klW
4ibazWzlvmwZJsrc6SbzRDgyXMu4qe75rUIqPf40pFdVROTgYTK9oY9xqb1q0tB8
/J02x1quL9bXmiR0AendBgYHuwROtlrEFcX0uANtp0yX9jmLcqJ0/QOKo/wS3l+0
IHpWkzgDQw2GtlfmtmAn4Ip+hTF0ZnwthoWeepEFCtTE6SPPB9RsL8od3+0FvtQ7
esYJVV5gBF95zscix6EmKYZ6YR8DpsiYj/2T44AtV/KI0ddVUIZ8/7eqnXImFFuZ
o0TB62FQaBEQsUy/cbX+wWtC2+JtqHGeRpIS7wub2qSgntH2DsNpCBPqfvWF9lnH
zdrwmcrBwP0uZ3jabJbTs1VjXldUiqujGz/n8DeCzajsPHlo+fkSM1k9JKkpCWIB
mxZnmxPUzJiSk/yRoRet4TjHWufLNFtbmNEBAJi+dKjLnRenbz85ZoLZAUhFGX9a
6QaNXV6UOONuNLWmZjdyHfhHCu3U3FkV+X1cssdLO/2IoFSGJy/eSnoH/nJAfDy+
rMkfsvvWpojGYZQXYCPCj9nXepApFUpnM97WWZ/0YyTrYWZzrGEULMq/vOLMWORl
vWHqRDzXd1nERKOAFLvgNZtmSQbBxLtl1xyZJRpuCnkz/nugQg7bN+IWtu/q/Pvk
LPc3Ha9BoZbdcFzKM9fqM9gMXeeOs8p6Lp3zos8g+4RrwLE5NI3rzMjN2VSpCRB7
9Vapsk1ggxcZDoilfdxC5hahtCkt6WosNOKcJ933g2ejAkPASvd/Ke2GWofRwnnv
UAXuvvFTSs93YH2NJSB6vlOBuVdDONcy0rSJEldkBmxZY38aPfnRqla09R63xZpC
CWhODnR08bhtq2HBFT5BksdcR0gWUtBBLj+r7ebXpMIA5YLZ4o7W9Gz5NJRwfR9L
MT5lJK9yOmOe/go60Loljw7NYdceR8w4uxOA7UNOM57l8dszQIKXawZjw3fdH1s9
x2G3MnFJNYAD+BJg+VALZqXo6uxcZoCHwC46p9+s9pKYVinH9fwb6p2Jkh4lXf8E
SIb4HubxuaDDcWp/RS4arz+dTlUTjPjaWRH29jVu0RMLlRxC6K8746X+gziQMe2/
+RRWL42khZ8GraJHUk7f7R+e3OdO+8HlQgKJDEQvGITXCTOwUGfRtmSN87AKpfC1
fc6VE1oRcGEOk0uUfe7H6zaJEGnO144+++R4lZftt0tywZWVOjC2740zAXDqgmhP
SuYOqmYGarKGMnBs+o5keHgt9Cs1JDSVgSvi2ROljbLAhAnrhO3Mr7a7DuUg1o6v
Cam6hbxYiRBjZf9PVGRT57oPKIqYQ6tw7z7awcDTaDjaClbRlpnVaBz2gIQ22FWy
AGT6bJ/M1IDa1XigUFXnm1cz+7L2zr1O8xLm9rxTzQYH8gJ6j2cPctVdngU57CB/
xIdpzcy6AiaDgrjXed7WK8mMRsJBQCWfjzub4l1zHdBsgYs/lzJdUyYWu9cVT/Gn
1uEjtCXCiriBclgnTkSluG9Cf4kgB+SCUkdTc7pWtRVBrTK7b2s9BqXJT060IYdc
eKHPaEgZeFa1DS8oMvYyE5TRifxWoO+QhvWqSZrBV+4iO8oI7cQ6fpvPb3wRNlnn
zSgp4F0b5w5XYE7/zzu5S8lW5QxqTUYumqWejn7b+J8f63Oy0KOWbPUxVjN42pwp
WGDTGoQN8WLlKP36szpoaw6+HC5w73xkq6OhCXJ/YcM80Vzg5YkjvAB/SNM6RPBZ
WPz80hJPzb/fpg7Ag2nCacg+f6hwEatnQ/d6lz1AOniw4opW/pMdtlFDK7zWe+ys
D2OHJKKcwUe5wHnSMpuRC8Mk3Lk0TMALHNgEtlchceCyZRUhDlPQBlJCNQLrgEj+
6hl1WNmAFWaBPxg9jb/sbMuMAnHt9wYwK2+UROUL3x3hmOTwqAnH9eZKpnc8/571
w/i+xNbRISxcF+9lSSJOHbIYb6jWWr2uSqs5ONOEdNpVup8/9u2DZUI2hNXezBnY
SPAWR0JjKvfnrhVmjErB7Y7m+CehaTr6fuSiBG7lE7veAs+9K1uKFOCvgeaRmlrT
zcKP7ephTYVL8dly+MjC3Rp9CStYk58u/EMpo+e8E8sjjdaa6NNJGqxK4SndjnQc
GiyFbgzNGm2Q8s4HwzMiMuf3G9etJ5ZbHJj9c6M71x4/vo2a1sD9RJfvIb07nYk/
EiSL3g4UKzM57+LzvT7cL8zQQGDnuBEhyotG2CLH7G2JEocc4VdAfoQg5IvX4/UV
vTZkOAlk7CFJCNdz9M/UUNGwHGiFR3aR9aSOMyUQqZA8wnNiG5R9S/opbOuiEt0t
trbDKHj1YRlzLnKvzNZvC70cmmPm7z6WeZXzua9NOnw/8v0HoDoKRk4OXVr7Rh+L
7F/aENpEygkrAxnE4EZ82geTLREOOaZ2Dj+kvHkiBzIRELYKiuQGMgtP4A6s6HpA
U7DPGWTAGyGTKa2qxleAyMSlM1jPOnBp62r26R2OjS3FuYUOmnZe+K3z6TLIIbDz
t8pZrsDSG3nq2cPLXY/slDNDbBOAJRF7j+w3adeFEDKUVOfNiqAlQ9JdtkVdjEz0
QoA4tvau2r9lnYEapRKmCJAmb+9+dhCsmnoI5RzXL+p7tOPVpCM5gB3QSLKskU13
q0EhwAxe7cxocPSglJ0D59kXvsjCLHLvUybR15M07FT7osXzG3MVzUf7OtLAQRK9
FhjgA7xb0NE/zOgHpz4tvQ2L8fnJZux47vitSFnjedadTw3PtQk8v1BKpzn+9zLK
1UkHMMyOOkNro7sS7HEs/BCpfZJbnVithA8te99fp9G/8tBkkwLUtPOwlZlim1sB
gLAdyKdlKXblK3Jbqk+xqO0Z188rQkZZ8JDT/L5ut+wGWZDZJwSNxHA3BfEqC3IS
LxcizblcpKUkKcMqjwYga8dl+DJv7B+hRWhxkALnjcSpv3A9E093LvGy1JKWBzuV
2/5E/4rTScHnif8WPtL6/nHSPfyuEYa0VL0JlG3xpQ05fKPH43aKi1S3hV7jgoCw
54Psyk1xjcL5CCJoKH9HNFaqqLtO9QsB7kQljjNjW03EvkP6gGnrnsddsIkpfpSI
YajV5LHEaezYwaFO2s519nDliVJedmMmhm1c81d58ie3ck8vX6JOMRvTleLi7kdp
oyp1jBWszU2U+B9EHnZibRX2luZ85hYWeszi+6IYF1Ix6Znne+e2in2e+nk++MT6
Ll+7GxtlbCGsU6r6OJ0sq6pWZzkKoyjnpZx4q2iYsukhCeMG7PMPqL/zfSJzSYqt
0aI2HDScnpYeEFy5XO6ZveBxajjpEM4fkfqGKM0cXMptAbz/PcnI0nxf2U8r4RgU
1xEkHsXfcrVQAl6MTJKDudAoQcNgaF1Dllek/oQ5jx3LU1X7x8naGJK2SSyjNfNK
vEcKaJFaEPV7jc9+yZSltgtRiO4vqUZ9Nx9Sovy0HWIzHyrAexIGNEDdndTy19kR
iMQ6qRcljY3buUaPSNkDZvTO21SaNz+OnM9KA+ego3kUjDXX3AkPBfvTd9z12jZv
JaWCmTnG9CkSVSWvqZDEjk81022K6WMGWki8oLMRQnMIXo9MMjy+CN7BNxCcY1Xt
AX9NLlh4nLLywedGZUwpZCAR+l4dMzhkj+6r9cN9oTQg8kBr3hp9JkcXxyUcL6Gj
1foD1er/gNYE+jqXIgCabla7PvaHf7oCljPblMCnBbVLRJTM7oWhV8mLO6moewEt
VC3vV7T4Ng4DLi4yuMkZFsLjXPN7/ku31MGxmKfsaaQXBRrx4MqKsi/edSE/vOZh
y2i6rp2Ao4QIkyZyvGgmKlYwZf8TtsJ3unPgdJkudUw9OERqhdFncpaE5SC2fOiN
n+b8tTVCkpBnOFhGOBG9b1crqGCYptYzynRSNZSklRBPluRip16QVXoGWYK/fNlA
VgUHEF/ZkHu6Um3qm3Y3WsseUxMJVv23IYPLwIk0MfhJ+K5gVwKhIiAwvrTHZ/7X
GadInK0xPh+Gne7yp+yc1DF21c6gUcaZRZhSP2SM2Lt/G9ACf7O1mAZlL5dwDgP5
VtCP3fDEGYK0QrytqPMHP/htic8nE3wsUF4QwdlkEBLmxAWl9Ld/oE2IuHMltyLX
WEBUSRI4KZhupDGSRh9uP26P2CDUbydrzUi7AYpkYqMXGAvSkTIHz+V4DlIFWBvb
BrHsvXqLJyqkVIRFaczT4R4k8vS6kmSqmE6A3QSXQLHYx4qWSbe7iqAj7Yap9Dsm
bh7TuW/iHshLp9vjpumxoVhUoHRrdPD6oweHo1qP039uNaklxJdbXsbTa+LCkRYy
46Ku9RISZoHAS2LsWnN+P+QDxf++A9wdnnc/vfGvrhEvcmHp7x216b/OJkwJ68EO
yuuyK04e8tMZ64VkOwkbDb3yELK7AKoR+mLz7kWLWFKha7jFUDI2hB7udNx8m/IY
QFvhlUHocf+NvsZeIkuEw9ELzaclfdWWwYD/aR4kEz3nhX5HTcxFMqfI4mA6c3JF
QCwXMrsopwPQzo38ohIuWdAnMXNd+SHloHwG6sADKotEa/glBPZQ2cIX4ikq0Z/n
o1j8rgPbnfdwKxrD/lgmC3nKjjCWEryX0mwrQzxLYo1MgwDCO7QArbAxO4WKjzmh
0uhlhyBgWqXAANcOgj3DUZhINyzzPhGiILIAtvmjL67JOfFtxWnySUe8KZ9Uvcgz
jc2Z2IXa9JmS3r2mhv8j7LUeaBQK6SGZjXSCSs9IvF9ERkJWLmkAEZ4n/B4zK74T
93Zrb5b8pxR+3x+mfjBKsHalDPH3laqjwjQJMJIr4SUGai455ezoFh0RPvOwQIar
EelU0ekgx/0pbkyYMISI+qD7mpvZcw4M2tAmd4DOU4OuVOEutddNgn/iyvknbt5F
H1Reea9iD55JBX96uqnP3vYZiBEgvGlXlZ/cdvg6LdsE6ioK3ugfH7M+O54Q/OEI
XG2YXtp5TlU5R8p+0QLghMUD0KvXvS3ZPJFjW5+ivYMhdArr7+8JhEKfRhQIBUlq
DdyI3GRfuaI6FCsJyBuSCcnGVtf/HTnIp2Nckde2+S6G3RXbW9TNvIfYgWB/O3sr
vmHYkRQ1n3Q+01+1/sRnHNY6VRxOMxPvCmxqLUEaFuCkj1Pa88P1BgHPg7nIeb4P
C9+9DQ1Mzostw6K2kzrMWAyiH2umqBCBr/Vq0gGWu5wmZ/Z+jTaNNe6bFLDDkLaH
k/vni8E055c5zE04jQRq4mQUHj8jYERNmmnVAXeo7QyOwZZMoVDFO8XkbBYXk5j0
uJ2NNDhFz5s9EJazMFRQiCQ/axHncAcJWJtNNRrLtvNTZS4S69z8e+jluVHGuzHU
WmWL0fPcmILptgRgeeT5Vxvl/ksHLSYw2COZHlM7hxuJyi9zR2WVT3jWYVhCRb00
W9vJ7jF2m1LkTCBNJtyy37YlzBrLemjdCVl3ux050pKAdD0yp+Q5b1EJkoot3vSZ
GJKXmiAATWQFTAVCy6hiNnw0upJGK1upAWg25ruW4t8wJg7BKHotQ9nmLRe7UGTT
QxhVm5rKrL0iX8GEmMxHRnYUaM9OGnmAoiSjysaib1wuRSTeDM8D0rbjLyFHvasQ
VBU+o7LCuSA4tmd0zjiIPEReg5oSrtRSYuHU/z862nlrIdpQt5wyuj5w5s+47qkb
mfC3ZbVVJ/bQtGekW1hsYx9Q2rBwmkfzcjsKVZsQl2jpy90Y9JXG6pG4okPkAwrO
8jzvnDAXP9SNQIjRIYRdFjrK53jgNvUNwdrmM9yPvvJ243IOkYzrpcx71yL0dH4a
yf0xrCkFr1+sWG/RVz3v8OWqAA+yXlwNCdgpUfxiH72VyKJ7T+baQ9c3zpYZQiQv
de5b1GrKvbpoQ+BGDIHqpWjvhEAKVPogI9HtOdhJL6PGOdUsd4mVOwh2RZNVYXCe
F5bh6oXWOKfMgHxkSbXPeKJ4L83kkAu34rNblbyK0QY59NwgeKsRJNYxLDfLbmpe
sJVWcRd7l7D7veMWovRg6KQpNWKkCF1MVj4bAQoIhZIp8yZDggAwTO+bUbZi0TXf
IKD62HQUgVsF+vyBGHgD2dTgU1BVJGEkFkYV36Yyk0XRiVrUR3vZt7ldSUXEDTyr
iefQpUC7bMTR9PkBNJEh7bIuCTGMDIMGYs82102QRaLaRd4lSJPzHwUvDSDlo3MT
6Il4rCu34unTmozKkBP3Rf0+ro2gcQDZ9zWn/huwOGLf9FNLrIlAKjeFL3PsvLk4
xDIXUqxjEaphFNq1G2BncewpYVD2g3m5TSXHbDTYKRcAGTOK8FMh11xnA24azAVF
VuMZxXFjAdi3BqhkdZsv6fprOvfnZupfL4vynB1Y4njd4S8NC1e7peDT7BGQDJo4
Ye2cv+jRR+ANxCT403uih3ZRKiTBvQADfe70iZpPqNA9gZtXH3KLbKDNvjZlkliy
kLYnlZV/1wGuLbjNncGAnN8o2ROV29Q/3kQ9DOZGI3uVKtaH7jU7mw8yxM3Ft3qP
Rt7tcb7IprD/uRhTmf/5nlHEszKwpLtlRx0yvm/KdoANkhzYnO7WTaFzB78QFMkY
X4kvDXtem1coEWXSakuKB4+pyFQxWTvtgnUZaCROWR0MN/DU4PkJcPqglq1By+RV
euqsBGByT3d7zBqx1YJTip/iO7u+q5AZ9/Md2Her6VYo1SbYLme5t4d6xXiflgnI
/mObA0pcmemX38moK7CpCkBjjU5f+loG//X6pl+9QXtSHBeVFHvV7z5PGrI5EVbO
6pZTdHDgyZaxL1uC4k+DeBo1q4Ryq4YBDP988dm0vCWx25MkzUkWn5Ayf3z+nbmt
2QuDCBaQzZYeLqkI2Q9EekhCignLbhA0K7lmHH7DasdMB4/9neiEzlmB66snexci
BN8ibNU1wRfg7+mJO9DzE+Gv9DJwEwNnPjiN0qBx67by9NsSsJBom2JRvyRnBGBU
7sxADrHtWrPHaDDE7+DwkIH98MSEh9TcuxtafBjvVWp7dwchdmcoWkRIhdjZdXaq
jDOAo1fAujpqcLiiezcWOJHT021iccix07DU4O0SUV5NHAOlJY4tCP4gu03FnR0u
NZydcAfbt5ximHN4av4oH2F+56Hw2ozSPsMpKUqek8OpwyD7rb/9swIBJF1XJ/5x
k0bR8P9IwnR6mEVxiWkIRVJbD3wwTvv48EA+9lahZ/CFuR7xvOUHa0YMtMZjsW5A
pXalENcylsIEKoGXuLE/7mLfc0AUNTTYQdw9Cd1YdRLghFejJ+W+cKjbg89LUWTd
dDZTLqNwsUWUxF7x7RrLylVUTr9dtBD4SrmWVQTavpwvym0cLR+Ndr2fOm88T4Q8
AQNfjQUtF01plqcS3s6np0dgp4uVfj4AlfubEu3xxFxKUPiy2waBrRhY6BZw5+Yc
5lQG9iTEwp5QRZ6LeG8IyyoFiluxkvJKcIEf0bAtMbE4z1uFWwSuNbp65tJtvYbO
TvvLiwXc38wdU/9jpECFdgdboqVzCeTDztUul9xQdNKeZ0Wts9BWVm3EEbwwS8vd
FOMbYT+KqqHacqRUXCDxs86+mKM6RlaX9tsKrGMTynDt35OR1zTGmgEQFSa+P3Zj
STGyl6ZSET58gKFAFWrYmJWGXzKmbFemOjtgJVozuzHcurvo1+HtNy3Dnut3hk+N
OlFs68Ip7bGAHfCjv7weQJL7VB/qiqxvvTYQ1U9pZUxBsF2GG2ZBW7YFOCcwwW0J
1gChO+Hi4tC89OamlN8lxbhnbiXlPglIULIDwJzhYUF1cXak4vgxiMUigEEhHuOK
4ng1VBFmpj5loDWGoMkjlFsgw+ePjEbr4TYZ1omcQlvAOtYbo7uYAuBCVAuEt2wm
snZDqqOVQupWOdf6EOcpSUtJ08KGwyyfuvKV1ytDzyLN0SEdqEdKOEAhSJ3IMn36
/68tei1KxEMO6aZS/c7WJE4ZXrc/nEhlBkipZRh0IziOBV2oGvmIBiFRtEhhnhZ1
mIqgj+/CsrcEOqjGBQGO8LJwDWxouMdwBHZk6PXmrNJgktiLhVS3vq/Ff8ZuVRxH
jEmZ1fjTEHckGiF1R02igyeO9CvAQWfbtPcvpE2Ki7uRVC+d+7l7r22TaOSxV/YN
AeZuEocc5X4zebryCOg/W9Q+xnrOVLOm9eBu0djTVodftdXptHBycjNzBeNVO1jz
/DSZsJYi8P6d/gmIPHT3Vt3zoqnzYIhLO7O0ud1thFcNPkuE4lRf66pnk9cNFVvA
6q5PHrkFF7Go9prnj0sb/1UOM7KGhnm5fEscgkc22rHJe9xGuN3T5PZlpJtvaH1D
YMypqnJnXfXUf4iNw6fpzN5IciYtIhhg/PHdTCA7aTWzDTsc6FifIFPJUHFomROo
Ag0z70SAzu6VWRrpcRoe69Z1ucDHLCAuz6+t0MEycaepsI+x5LkWkXXvBFksBk+v
e/z+FAil243AWB3zRTgE+m1+HOCzGJwLdvKWxfIpQZQgfo/ILDc/pw5+P6V2I517
t0DIzRGO8Nm7cYiYXgbUko6OR8LIRWV+f7gKlxpq73IcNsyVjjI2W/tzT/RRrK7h
wx8wqgAkCLwhyjAY6hpk4OciR9+ZPaCIS7CtfjXLAaS1hI8D64F7jhrSgMzQo5tb
+aFkTNpMRZr+Uuo1zvrQBQr6/0y5AfKRnYDxrqP7OtS8hDUw3/wDVRkzeCOj19UW
einvaLoOW7R97CN7mp6HxosOcAAnCzvn+kBE6f7enILs6C42sLNrSws8tHrFTJ6m
Tw1mam9D0scC8ws7dB8j57ndT3CRO69DEcXSr1fBlWTe2bGGOMaYcsdMZ4124hAZ
Gyy8Y7yuEANPf1k7BINHFBF1iWESu9ZCParoUgt9jCWU1iXrLH4gX8wyyRLMJGKm
NNsE18pywIxmQ/1hmGk59uFjZ/zqWD07rwoFt1ZI02G8bn2lsVTCXrc0wF9KYhfm
EpwIhS/Y9q4nPvMdSQ8xDpKdzGfwARaMMOyAVJLVyiZwckCwJ56gRQxlOK6cDBxs
gkFau9NoctlPYZvS9zQtqbIOZ1M8TRMeChBJk8R77fngNKtLIehq+jQxw6117Eij
ZE09+ZVNkcihYUrQxn1kZS+h8Wx0JTkDzff2yUL41d3v3WMSishApru8IrZCeNSk
JNPpvOwvv4euMhW5eHXMYDbs0X5/PGTMqHHGyn6/NzjlNmnQIYfqfLb95C3MXk9f
7feCWFywEvQajshQgxTKv2wQw1df7SY918v/0xwEdseQ2G9yZpndWI0/3gnmVpuQ
uBy+f9/SQn8LsuIy+S6voGGs0fiw4xhooHQCxNnRmuhjK0z9FLKdTZ9sWhIFaE04
nLjXLWTrW7bekOtiyNrCE0wIjCTVIS1q1WeE9NxKVR2i+Cxqk1pk2qYplJZEGx62
Wwk2N3tkq0PFStPOqqGB0lKMhWoSox7yjVkzLk18enL+vN7iG0v3mWUaCsKzgsz8
8/85TEBcei9paUYjz9ymh2LP6CI2PTkNZ1orCaqFrQh3XXApaH9og8lsfsjH15aD
UvkJgzYdud+OG4lpCO7f9hK9Nx8r+p1DkzuGZRAgkbGvsd/zuqB6K9N11UKgVQ4/
OVjADjsvFJ5t0azdxvHi8ygpiyAm/09NE1hHqQodUELOy6weojaXxEixX7R2x/hV
oyi4+qE+IzPMc0WB5GO97jLz6QCJS3URXAOf4++9N+0aXFV869z5H1CWYH7MqtEk
wBlIWuR2GXMbuv7NO1eDfmGwchuIWJV1a6ppQVtmQNI5o6t9KyJEu2Bu241myPLX
1akaEh5k88UYnraNRuhvEiCcW9EneEsspHlhSN8yqOoZSiYfC8b2oBWB/ZfjzjRF
XuDZbXFUUB8gdCPHHATSTMtBPEsZRLRKdT+uEHqlb4M/+6082e44SERxrmUFureO
M7/homRoZu5Nj89n0oeTU2Q92FAV6nMPKXucIf6mhUp+cqVa5uv9e2y9WjTiF2QG
sxINwivvbzbE0KTYsu2uEvGBKyvgMkve45WY63J7OOQLsLVK062EUTk/NHGD87Su
c2v1o5pcEsAEfnsP/sGj0pvBAI78z40LZYEIPMu0MW8OAWHZ4PZbvQ01IOFQZa4g
maC8kAnDhfV7TP7gN0FvjOvFFDZ1m85i5MyWDi6cfBKbufauP7zaK/8aP9EM0yyj
Ft6yqkFt1uCGQpNcCgoPsn5mzfZ58xAGNEHObs7hu8sa+pQyHVtU/znBqBlKFUES
6pZhPr2GJ/Iq8lYqjpyFgPGEWC3nrfnFrGiOkLvMkMjs9V4UheaS618NMoe5IhDk
9Toz4PpuQdd+c3tPQxouhmtiIbg1Y8Da2IshM2h4YWxQHBCuTAP1cFeE0F9j5LPf
1V5d2/isgg7PR1NVYTtquDJFL3jVaV3iSkeSRAU/8be9fqlZdQWS7u9TF5gvNrR4
CQMd0CQ193yc2k8ugXJsl7YkSoRXQKf7fFb3Bh0OGq0vdrPblXfHN6qwQLcq39xg
IM8HmPY+2z+RtfhePHxfgNIbJRyAleSYas+V6FcfA7B9ulWepF2I74SHFC4CKw+W
RybffHhjvGtRmBB5m5eLfbi4eE06JhKWjepSLlglgB9Ird8zy5KyK9/FwSeKsU+a
vFL5sXDjCVjPBPrCAjyMuvqR5B2t7qUW34rMz3IBpFr7Lkj+qjL4fQvOCYgVFTtP
NlC+EXpq2Yl3VLlBCXdkOWkfpFzhKwZT3LkxmAVxNeH4i4IcX1p8D3imRRp7ouax
3AHole4Hvtb/TXyR4cp3AwNa2w3daytXU8A8BqSXw5FS8/YauQykXg5dh5RzxvQ3
dVufDBHi1Fea2IGwbCEntjpF5vUjHLvb/p1OXojr4DO018prpW+8hlIg/v9pV4GD
GI6dVl2OGvzOkYxyouKJFeq0aYC8kb5p7r+MenyXnwjLi5I43HiNiaJENXH3GaaR
w6h9d5rD6dJ6BbZlBF+4iYsKgoxhKDN1xILGwe7KxXrQEsfHuia8o5zJJqIZWDAc
uu9SdzBzpZFtO+8hfpRGRsdEiuh3aTJdMFVcunCpWUjs/wTOq3TBSsGoOFR9p6te
Dnk3fWxjpSmjFNoJ2PhROfkV2ePR3n4+XvEUTcaN0j+Db/o/7Q50ZP0f29uqu2Up
lJ4J+VhncpI6zFoGleHgFIqMyMIL7wv6EWdTudk6tBecDRuZvMvw64C8BrEn1vco
peTpqNT7l2rpFuKTsrg4IXS9OXxZVkKRwKwP+RWqr/21i9lirmucUGf3pO1mAYQj
DOla8q7TItg6ETp1Ky81LsbkAout2QTZoZ4mcflJv+wEaG+TfL8F033MweMF2lZU
RzUCkWHs2gtiVoXSWqte3fvJgfqTwWKmmBXACr2epItvjYQazJ8h5GhSh1e/26pK
jZVRw+r0QKMe7gehtZzp9YH5MmOVUdmpiluTp42t50nRiSoDk1AnrzmER0BzAwgd
Hzxv9nA16f/bLnWt9dTnqYvqVNhUAWGhZ8oGzYW5n9az96LV0PXPOesRczVg047q
lkvz+VtW3g2JIPzWBCSBoQV7opDEWrEGDy601fYzjWm7gPuxqWIOo3iGZW/hW41D
9U5jW81OGuBd/f942bDR3JtYsSDhDBexVwR7uskah1JVl1flIwSRSB8b/8QbnoNW
lGLmu4n6pkGcvAyjA6NnWGSR7SPGAD2rOgv0vmEUh59SLODmy7Bhx9iJ2ZhLTSCy
a2tJXVvxSYVyXgSWSghPO5lBVRdN2L8/uWcse+AB5Rfr0K/06umzdYQdiD7Rhdjz
L4VV9tUdKr2u4NbEu615FmMnvxrcMql6gh6kehbh7nkKddf3XRPltU1/O+S7EQW2
ShiXM4CD+u8nq/BS5vTxKqzy2Dk8cXQj1RPl6qXaHue7g/w97qtpNeH1ni9zOkbQ
1U8nejEW64COh5Z/CUrm/3ImYQMfcum0IrAtfbk6/syu1mbz4c2iAVkat0z5c5F8
hVxb8rDUHQ+zNCiKLguTMVZ7KsQH1+UTxEE8GCJqvHx+851iUGGeStCIaPKQjF8Z
N5TFwbPgmNIx7gY+x+cmZr78YkmScC9sZys7wYBKJa1iLyW/cts3mTuw4LB1SWxd
82CkyMy/SzCWMcWuQAs9l1IP6yiiD6Agt+LaVx7zFt+dwSK3kd5TwjLR5OVlvZIZ
1kyd4bpaHxTUMJ8DYXaMKS/zHqZJetbsJWp5w/Do4Ow9b17TVw3T9ERaUHDbdHNP
xHmU7tTCu6Hr5sjhjxL1znkJxiYX6uF2ACd0HA5EVeE7HX2BFMk7dbMOJlo7jq4G
PWNw6XmJPPyIkSoKl45O5CEFpTOFEhyixaoqAVUzyVqxJ9KtsTKwnT169guqJhvh
PgI5N7Jwi6xamwmN2Tfcx+slUv1tWBy3THqIe3HAqXX9oNX7OblPHKmBerTGep+P
r4S7iYs8XpH74O8AXDENd+YU9CesCMhb6aIStslRHKOtV4jHjV/YYvfmY06D3XUO
dc9NeXPDaSOVmsxCInciDOGCkQ1mKE6ftx1abwKAnsKyMggU8Bzwxrz+1uEGW9l9
G6tisLCs0K9B1XfizEQ06kHw9s/YdX9ufK9adiCmqudj4GqJXzmsVtndFTCVDzEj
I4FRTy2fqv4dyedNgCZ4Cl4PF7bw16jJOZdTsBYwHtizGbXbCSO/zI3YK/ZM2IHP
CoVNQvCERJd7Gr/7bgrcJLCsRDDjQQp2iHuUGWbKxNRoktTy2OAtxirA47lo2EKi
T+xs9G4R5SpPxTQsR+ovVzgK9Z28dnVSBavQARYtsDjdWNgLnf9Xjp0JWI8G2GMW
ajjBmLIk4oK2jMuWP6LmOgevfFNiqF6RCVVdpuY9vhKpRdY4ejHyEiR2cS1NA4x/
1M7EKSo/V/OMf6RxGFIc6DDc8n0QhZq/8uX+MQKX0PPqLsCt18z5IXXmrj4aQlk4
uQsvRZQSWFzFUuCn1qa1+kWOSv8jvXZAP19u9bBvZUnqEUi6rrkZRfBB0jnGHtWF
54Ey8P5lF/CmZlsBaD4PcG160SocyXI1jLJzggXmT5I1G5Yy36OZ1hOjx8E+KoM4
XBnPUWcox/JskKF/cEZpET+QvRn54KQbFHcMzDCc1KCQ/vKcYOjH9qpBgjvwJpje
VchrWUrNDV+8q38tG6OULh0jm7d9wOd0ldVFBqubKd+yatwmfbUNgKa/QkTFR1cJ
ozlxHu9uMPmUt3KWN6AkKFSOeK4IlXDsCqEq/Uto/ZtP4Qcw5Ow3/mIJBj5ABtdb
gA/rOJLA4oo5+rR6CjEla7eUajD9mj56OjKZ2CxY5syBaAbKUgmRRCCag6HnFzYd
xMEvJ77hPjXwwKNoP/wr1keS+faRRDFrwjUU0FMPI+2MGatcP0gsDwNiyLWL99kC
EEw5+Br5CRTqyJLFWQkCWJvwQct4gT6tJs0JzwZ66ewqqysBFeNQ18KDmJtQbSh4
Z8d3Cakg1bzfKtl2mcdlErRFlGkkacO48H0ghV5MCKmI4Le+lJbLdRoJxb/PXEFe
Zd9x+obnN4EvNaAWW2dxXhAJ7OSSdLOoGqniIvSXesQrEPGSbGU8Vq+/z1PzZi1p
NGaC2k21z9mvPMDvOW9PZkCD6yb2Ep9w665uo+zRYKm6YepEolCAFn+poC7x+VUv
q3JFI91P8fRwMGpPSrXnZ2Mk0baHUQ6K8iCoRR/uvs5KkYHb2S+WYzi+iZ+HuOIu
1AP9ABMbfsJTO1FtveLDu9VT4qsKe5bl2WESH+Ml5e0mBcC9Nixvxis4FZh1rHGq
2eVz5YKQsORklUPaKs4CS5e2gsjBSYC0ncBdauDddkqLJFVaihS+TM3bayqQ8sH2
VKgQQsvVoZ6t50RFW7sx1eeymc554EFpBbwBrTL78kxcs+7sGjOFfY3GNEfqCRrF
VTulKDcXBnM+xbZsdtVPU1S9AHT4hZ01PTTzXN+Oh3pBc5Kuepr8HMKyJoqge9zf
h4gac0oqCCe+NyMgF8QDgycmYjx9EEoVuu1CoBUnoRHN5lPP6KaA/MplkJaxV2bz
tI1XD0MLNhm9IqLgxUY+Yb3NaGFCsKhQZYf0MxkiN+N6UEO74kFJmQIq306tFsgL
8ltxYVFbFcEYd01Y4GqUkdylnJUI1+fLzJz5i0DvuJzUaLyGZUB2TUDyooOcAiFj
vg0pWQGc3s5CubFtnlZ6gFMCTn05ZTN3AU2wzbTXQImByLP6Bru1tDCGvZW6A5fr
qQKv7BVB3Bzj2NiEfbkVihfqoRFXqB2C1Zy46J4s92sKy1qobwTnok8RYzncguB5
tOfHmdpAFAKhA25IJUCGH8ama11BPhFZn81xUUcHCPPaNZmU5Xcf2Qx64uQpvvJE
VO/nWwq/1n6ZH/zIxR1LPxHKoWwqwXU7nMcxIYcLopiEaOLpBByXlLytgviM4qJl
0yi8B7zrttK56a2pTIpFqi1sdI2QUYDHwEymdjR75f7IJYO32TXBQOKkbcQz/oiJ
VhDQ3fGkSozUMD5YGNeIcDdyaFlll4CeZ8Ljsd5rJ70nSEWzxk/PXKMK73hr60a2
Z3LDQe6zqaXkbqXMm80wnYKYnrPZcG/vtWbS0nn8TB1EhDq5H6xXQZRL73yAiSvh
NEkQ6BwD9V3BgFNTwNn1x3tJOpgsd1LeM2sVE6KcEcNqmSAj9eLgUq3XHQ9tJ4yf
EvIQCQ5aCKPpbvyOfMdyPpzdqqNYzXeK703HYufZSnuA68Cw4yGSt5CUDukti1AA
+YWog/b7L7E7U/GozmmDxVqEp9z2bXOarI3k2lSCwmd6WyyY9FpFOmpcUlJuFyEC
uktdxJdZiCKEZiB6BpZnyWudUHGRBV6MLJmMUznX+jHSQf6OIVDYq8T9g8Jo+t7b
NjLbLH7xrlLTcZWo1CX3K43bAPGMY6svNF6jDUhcJEcG+h1QBxqkxLrjbBXfePXk
P3YDj/mZh5Nin/Epr1YrfDU0k8ephnMaPTkn3UGE6AJ4KrKDSK1hvYpRFfoAIvsX
TAHp4mptNN83sAI0h1M6NoIKHYw/FB4wET9UfEkMCiGNl3WPruESHzESVD26749H
6MAtde8+FWVnb4JLOQrqzlL3waVeaM5rEhdE5+psdaIjCOuVCRHbtz9A6TRhZgqc
dW1GVs1mx5CxJq+O+ak1mdO9lPRx17taB9PCuOf27Wb7UYb/uWzJRPtLKIvsB+AA
M1apLn3Qo38dXIYYHA0jyT/hrx32PK52ZB1AOdyudQ60jt/eGzgju8R9l06cfxD9
5kHlUQu3ehRCc4Wv02Zox6+V3cqSLYUvdUCSwC84bt7SJ0Y9pDjZTqWWrLcFhdex
lBylX7fYDgXwoyK13IWdFrZ0lPRTqnV/GXoFcE1YZ+j7pYh0ZwQK26HphaRdrmaH
utm/v6n6O70SNY7rDvry9NQlkyOCZbPTUbcn29oL6Dpmnes/6FULu6CuR/RZM1c4
ZHyBsZWdkSq6hWzo/kH2sVJy2y6nLlxT1f4Q8wzhZHHg7Rc5hI8c8Jyj9eUV8gPR
8BixoRpUkoTXHte8Q71e2rQwCZaHxh5BcSFQz8GU/9F5o5mqvr9xmz4I/rlZze2t
qBGCZ2Lqs6yQeNGg1d1ROsvtdIesqD2qqZ6oFvKkLzn1wMcSQP9wrrEAybDNwHbP
MKOG1jHbIfolinqU7oJBDcucoDAVzEC4YYMlHXG6bciNFSMs1quda2lYiTwBZbIr
+jPhiQLXMfkaJsTtesifW5SU6vLDCbUSiOK+nLuQa3G/KqmCHaH1TAtUgZfgFkCu
bCsvLKVXmL1QmL9VlkrCwAGCrM/aAkwN9EAaaFMfI0d/qJtJE4sdpuz5cSHMbzlK
mpxyxtE+JUKt/7yrIQ6MmZNAQFFRYnhkMsHTAzsreFA7Kg0qPLLmGOJFzJnLfiHs
S+QyWda4QbuzWMMQq8vOQWhc2DOGf8gOYJebQmoNLHFd0MkVJ/HDl+W+Wb15yFb6
CzpkeYwl6FZmVhtBOjOmFpESXn7q5bYQuUva2aLM44peKSUsDylnfgCraa++B3GI
q1XIkX0oRWbXQlsLmLD/HZHp2EV4TWJrcJsZDgYMXzePDmDFwVF+gtvYBRb7q++E
1sTMB1Baxk9wvjeQbwhgf5p940FsdE2wz6KNlhE+/62FtB/0aOTKuFWkXeMcQtrT
tMkyRQ8gajRoqgsNZlX7+7s+MiIg9tQmdG/wqGD1fHxbR0y46H8pUveALNI2L3FW
HyozfriPIFSN7xG+r5paT6uei8vHc3dRLDoQx01grFUKFUTo7kHZln0as+zYNkAA
s8ZYxuSmRK/0eZYBrspeg4EtGjtv2NP1eTlQV5CItm7VzicoW1a7LeeOJCllQoTa
BFDeIe0UR0vHXSj7mgaxXOCo9m5QXuG2Hzil1Ak8kkypWg1C45+foCoFTpIIYNG9
+0ZZNGfFRx58mWk4My5SzLEh17V+L7tXiMNDc6p/6wDgzooWVZsIPDRVhH5fG42D
FqbtrJ8FQyHfu3ZkVoHAfDcw5LtayIyvVgTvXKJg4lSz2X3ylnVGPdnPgm1vPxUp
2/yirqEAfQHbtiMwMNMQHdtm9YtscJho8NVrtNEoFfAEqJLYmE7zSpLn7kAAPK75
YER+mlnrUD5UH1yPZMfz2vq6I+f8uOh5i05HSUZS47FihDq1H8W3AJ73L3MB6C6C
rd3gReb8Ji78p7T5xbHL0Rf+GSNuRg5qqkU8M206yjm6KdlF7B99mJrF6iAbijq/
WG7v9Mg6TG0D+AdNGnZ4m0n6l1k8ZjCBYF0rGNRWF3x97NUHdGioKh4EWfYR0RAD
yXU+Fiz2USxKXnhMYyBcdG3oYxmBdMo4bqy7dBS/igmhrzoMpEV65uQ9HoijYQ7M
avKDdpm6jpFx/vB9zAREiDZEjQeO+tIhhc2/SH/Key+9+7Wsyqq54AtmW2q9fq0R
9+PCoAok1I24n6/WYxm85p34hDM/i/XFmTFDoWSC4mJTG3hoenta1qTiFZ3sNpuA
5WjthsdpOLAQ54nHOxqgBnqqKV/dvXTUjlRjTnNpnoSLvgRUv5gZUAgVo7Gprm10
VkOnpHRJwddEG7Z/o139FpYjMWXg526flVXPGmMPkFI6dK063Y+8zJzypgmqx33c
1HeGjH3t8gJiBaRoP38tAAnpr0tEb8ep6Fe4tx7/yCy5qyjWJK0XkSrRGAWMwoOn
+6Ng3Mth6DxoBeaHbQgsu6WD2ivq0PmFWdZBLrDTnlw2PHIIvddVkmlNeYyWAIsy
CPBbs9g0nDHS2GOzPYeMp4WNQczsQabF1Jg0d3MPjjWdC0tZsb82HKvES3dVkCrx
xz2L7HpbIT3DyaBl7oxYrchh84NhGniXNbsTRxf1pFMvyF1ngwJSHjB5DOWNrKnz
1DkGXJ+LdyHuu84btQR5Txd4/zUxncQ7ph3n//fK6HX78jZ+TtNXPr4VbB6wJLrE
fvGgJBsuj/Ib86hBAhK+s5S+rp2kInzLrAEKyrn+S9Bk22tD32+l9GcvqiR142OH
N3CfHVpk0eC12AKOVl56IbDjcvTOlBudcxmuqMPmMn6UsozVyvj5M69cFWGboXBZ
APFPRsihHDQV7Pr18Ssvleqo0IP0FM9SWK/2tpxJrwnh0VYqATSscJWQuIXfWL7N
0KpKKT/z4Zv/rsTGeSBqtQlVOr+CHcoPJpde6AKaJd6kcN4v471WYNe7pN+VUYiC
up2x/Ht6easDVRSlroI1+jmr3ptyx1ExgY38teFPlVwUZxak1k7e/0mG10qxXFUY
dL6tsDuPr7O3NUlVNBNGInA7hg1ik3866/zRiasIODKQdfQAhWA9jSgwJ8GjlXV3
v1Hzh+CB3aF6Zhyrj4nzqyH4YMLmt4RgdoA+IT9Zz0qSMIc0hQPUzm6bwBinBDIq
r+Uyn97EjEDDpaBzIXr2cc6j8ly82CcBREzLENS0HTHoEzfTBWRNDC5W0pyK8muo
xQ3MomUs0Oy+zTmmEINJF4x/E17XSlo/htb8UQ3ToKIql6AmrtTpJNB2fVURT8au
OGGRggsHPSymAotEb82XnYm9VSKZzs7YeJAjh8p/AdMBo1BZYM+pQEmcHThJU9xC
u2yDTH+yLUFnM1VyZGoDyGL2ADlYq2JiPQSbfRocHHECez3+XaRvZr2j8HH4hhOF
DmrMvQYSwF/rrWekqEhSRQFcBJKP0ZU5gcZSsJ0YjKKte20rysMMds+HeT4Zjxa1
hJZSYDjwfXQVp8gDjiq2OQ50CD4SN8hj9MT6n1ZOBPOP9eIMkseR3Pj66kCcGsqF
ueoXGGxKzjvAJg258VhsBQ1c73+t8IN7VKls7pS0/Gy12irLOcOtWtXCeZc8jw9i
n7NYuNbnSxvT3g7GLs4omyNHPXzh1FKlVVaqCByFzwiELTU4wrxvlsiWLyckh+oe
pgFI6qSJCQb33jtprEhS9M3d/1zkKlaUljWRPXaoDpFZANLzlrjrOio/4ubIgh/4
XTm/Llh3bYPJ6dFpxDe8eWN5IZUU4H7G92/uJChFIM4PhMoK4icfyZpJGUR8CgCC
AyCBY4TdLUW4sT3om8r0xL4IcDjW97+QQUSDupVWeSbl8u+hPF9m8JAyAgLNeOZY
ZOitc6xxWlSr0QhX/wCAFMWLL2+eCTFCgTz0Ou84NHpJcYo1WGPR8CJLMfuM9gmi
4YUHflTewD8y+8xzCcyB+0exqAe74DElE7SYHlsyGofU+EHnPkLpZ3DdWVL6FYnD
e9PKBi+XvLgTDDngAjPrYNaCV0K/9rxtsfCUt8mtylp59nlAoP8FrNP80HFCo3I2
dj6dVIcQgLkP+KymsFi2UW49iw104DqdAYR5EVSy2X/dcXTaxO5KyuWaalob6O3O
BvOClTIlGeLTWfT0DuCweDRu5hgWkZOHDy5g7LVZvc0lzh1yjT/y2YQ1Wze0W1YQ
MNrvIAjSvllqaB9JWx+zx7AuxrMSC/nJlpI5czK8XgHhp9nJHWbPKb5F9nxvd41Z
fMjy0+udZd+4nhpEkMasRf+RnyMw9ChZJgMvjpR8HE4p+vjfOyQzZXOiE3OffMF2
jplAXhIvHR80+NTvGle3XQRVtfLX11hw24d+G/GPk9+BgEtE8b9yTNWraYw6tXnc
H/8VSYnxGPSt+VOO3RdEitkjEns9zo6p1e/eM2LXTXfau65rSAUtNsKjeTff4kr9
Kad79bkbenELkiuIUz7wdaDgO6Htu6C4+3UFhauslcz5mTzl9pnO5ihwzLZlwwMn
gE3QymiJjZlWWAWdUhfqJrcFg4xWC/sRSE5tcgfAb+tvgrrGyYGX7yB5RxcZO/xo
dep2O9sDi2ceEwsdd6m+3YOgvuAFdpBypDuR3rcw7UI55Y0N5mFGGfRsR/4Wc36f
1SAoKY3ojVPxJ6IxQZkKVpjxPper6irDhfjcHdYNx1eKiJWhMORv5LepkR9pucS0
uv1U2p4BqJ+kcPEsKYE5945Qd9yQSTXugOu/QT5Qx/j6gLGq53k/yNOtv1+hwW10
Ayi3i3OW53bI5kZvrqX8GtfHuRgwhxYp1pLWHvZDma0T01kYXEOa1waO/g3ol25A
rMmf/iJnrYhlUNuSOLo/ZcBXKnuBCOlYsWYuQdPqglDxlIFO90YiMJZAMcKrO4M1
vWc28dj00VXcGrRvQN765s/FKXSpBUefbn/WzPqcs8XyH9LlpiqANSIjY4pJJmZp
PZdHeTz+0fCxl7bhHXiIb8/DMzgIgtyYuFgHYPp9027WPt3usM1wD3h5aUQukrQm
vK3YrBK+7/1DovL6SOsA4Smw91KZutfui++KpGwKzUn0GCmBRjBJZQQJW8ss0F82
3w61AMePUDdqSxRXM2SkWqFip2Ao9QnMVvD0uJH3BP42IcdotYRJrfcztOUf52CQ
nGbwUPz7WGulcP2GFksx7WQdGLn1rwxjTGDMeuRZkKt9fD9hruD7jcFa2K54VY7V
axINwG2/ApZ7X9kh43l9f+f57c37cRFa8peWZ2oeB1oAT0GBBCBuuosd6w1NTbkB
nmecTWv9iTV2/dKF4w+Gh9QO0Kn9G+1mNQtmljZHfocV4qxPLyz30SjRmRgfKEjh
X7tdXYaWMIncJSdCT1p25h8Kcdi3PkA9JmGomm28FqOy0ZLz2vYgPmBgAMIGKPf3
SDBxWgcpLalMyYa8imdlCBloljah78aaPgvAxekW6xkUrOp5W8fPZqaAtMESsMYo
e2gjjU5oakFTcZv3PnnVcl4xe/wkAyCZEbW3B6JpmEmutx6ABC6+81miPBEHEBw6
8N6Jb29z48PjMAbDBZLCMrAf4WH+NlPvGBlbJ4JvvF/PEGwAY+YjBrCTWC+8nMt7
8fM0KgYbkoeOn316tJ3yp8e2dwq1n6rvpdYnIS94tQQtapTZqvy/h9W0i5dwiwlF
/WMxTcqr8bqC+t/L3px3pjMGVF1nDGUla1rgJGLOkZSM3+65ekMUoUkv54d6IpCW
CaexA2+KInW8WvmygxW1W4CwbgXfhKUp80j8fjbyeo6QwRNXMEKdsyXcSeyjgMRO
VZDCCElAptiMytRYsOYK/QfAKPavhVZ/fEJt/ps4H/iWKJoDrIzDU7q97/rBz6pE
1L9MrHkUEfMT2+dMYAsMfVQzfeXWGwX0xatOorU4dUqZSmBGgC56EiwWB7UowHdo
QAZ9CHRd+yl4KdOCAKVeyHHozlLBKsSpzg9KWskwZuwLOaYCJRezwvnl8dc8+YvV
djm3Nm+76XoQbNp7S83e/KkX490VISAZ9Y0CpSfKvVr/Q9X5Kcn/UmZddqA/c+if
NVKGdJ0cCD/lZ9yYBYz8ttnoCJVbpvkTNhPzLZCruWh69F1yHIyd9a4ADW8bmGMU
YyDDr6ivHiJlIadtMWhGqN2VZdnp2wcF2hio6uj/E7lP7BxwT1CmI2HngYm2TnIr
eD0v8QQopv2YbmDNYcgt+2SQcG862oXqTGA7+r9GXXRqKTqx7guxTm9M0S2gA4+i
O0q6ZyQYwRD+MpvOy1FTpG2Uc7gOoUWzg6uPu9rUPj46foTW6QsnI7mZSILD6N20
1PvQsk+SDopM4pCb2AZmYQxjOxN/5ClcSOsIUt7/xS86UI3JBvOw19pkwPG+JJOO
o8qB7TNb3SUs+g5VI5oQ3ZFfhdVf5LMlxpVFTAQeNudNWQs+b+C0k+d6aSiBIiuK
VBxH+BpGMPM+KR3qJMZsVz6g/Ci7ntPsenUoHgqMDCXELHsla8DmFJbis/ZBKLrz
LCWHtGXIS7SmcJGzmpQpVUKvy69CL/gNwNZaHHEeuDgZiRi7dY9Q/5wDupulD5O0
XzqzL8vXzIBIF4DpBpUAHETQfEZc78CENj5V7DoP0iAlWIHqeHheyzSvYK1D7Pr1
RIvh47CWo6goo1vTEnREi+bC0SxNMouxGvXbHs9qX+HYHs0lkwgBmhTBP4osQfka
zJSQ7O+VCUzA6KKzzzKyvQNCUemlvJQ1icJ7QNkLy5B8+6/dF8wHGVMTS5DeXYtr
1CKpEEo8YATFlyCnDfbwEhQTMrpDeukqUHJOfgFMoDLGJJLzfe3+RT0TKjjpQl4E
hJNWqcdZX4VdaaiUn54eXX/gpp637yqlz1LnBQrrXzSMXSejBSa4ZKJi8m9lCQUK
UNntOm+/zECJPnf4H84vWQ0dl+/9ofOMZONDqusfqQINPpM2uzutzS6IrsE8bggE
Vzejo/NRYHe1W62Zfu8hoVevP/baIDhEbz+eAFO+HzKCDjaGHr4WNqs9HxrxxhbK
rHGgrbpOWdExe921ydDyweeU8IQisaviAzxPJKik3UtRoKnZvyD2Bvj705yHz0Ig
BBdX4RQ9xqehaxpdJ4Fj/dcLUfD7dWDzPnzCoVcLl/BJKW5aTTKQFrRc4wpIfsGd
NNGnojjbwmiWpOFHTSIBjBSVKBa2QPES2sSdYTFyBTZ4ExxhZA91FvSmPYCI36RH
FEUIq0nWVaO73F0FeRFFFX4zloeK+8usKYH3ezKXJL9zPX7gUxOzbWPsEDN9w9DN
3UBqHkIpBrBkl1WMLGt6wdZ4uCHCpvHukQGuWlvM77XLN+g1LkAeyVLkcJR96pAw
DMCnSAfWUlypcOrFZEQZzCSvn1mhq1vkXl2QmWaJEGQweLj8k2UySbyqOYQH+GQu
X1Cir/7wbeV5yP3RE9zape9BMcckXZrBVlRFS2M14P/ia6MBw+dbLjiTZjv6VJVI
8TwEkWjoiovxD5n7flrYa19a4gAE264Z41fCVZTKobwTU4VCmAC6v6UJgCZKJnaP
/XWYPYCuucmR+D3JH/sACOPbxonyL3aXygE20AN10pT6O21hJNtNg50uF8BtoRce
Kvhmgf9YIGKPyCzs1eTbT+BmxR9wHBORXgeDr7xaXbjtbBE+QLgjJzZh9oM5YnkU
vJw6zvKUJbBPRsNVOnPN4xrjnYI6Q+znMM4beDo/PQbbHtBvEUmfacPJA8FmlYYD
IuSsliHoA+JlklesnWqm3b228mZFWrmjuSB9IlWSL3MYFxEKZPbeWEAExXCHYk0n
d2twb76eHbJq6uIMD+vbqxRIXLqS1dLrogmE8EvqGZKkBrFHHzw93dFsd7RYEJPm
+9F4kvLx1Thp0GwNWtWCjTPCQImiIZYsjlma030fBuzf0yz5IPt5mn/rGgvX/PAd
G/ZXa5QC1NeqFYCwFq19fyQDyvRLKwkYLssnEjIIJvptTRfjrUeQkTj+XsR7u/0v
DvnEBQtJtbA7lmZE9DbhZLeyygNq6dG8psgVXwnCfVbhaKUSQBD+gcrv3/ueksn8
nWcZ/LODcEMpHrE3/05KUFuWzqMzS12GFpTD0rvTHQPFslmamK5t/u73nXN5/KEC
xGc+dNnv8yL5j78YG7vLdJn+xKWmBlk6YxdEK31r55mkOgvseMwciswp+IFGkyCX
PzD0OG4t8nmlSkPqGjO4bJzqofMUyDWJrMoeiqvc2mD1TKiqVwefc7QGTHx3cB5r
GXmg1XTPdg0w5L7CF3HXgsjhn9CISZoLYQi56LslKpBhWqGPboMZTfJG2rrLCYQp
IlKNpoZQz8pOqOACDHtauDxC4/JaIShNyFBxNqr8lCL+dcD3bMSOAqyc95YJXR5y
agHjYnMABT1p7Wx+MNUCLaQGz4RkNRl6Er63YkpId+mODOpSesCy1F6pbCLpyLcl
/CDotLFN9Kf8twQylwmphc7tkCQ5AdykMY+nwJ3aeBxNb0xsI2pslx8kmqFXOixk
zVF57zuTEXZjybZWfTGNlGSfco/6J9XgxXCbgTv/O/2XFP0yd20rtt1cv3q299Rq
q/WzfV9SaY+qUzEGNX3GiZ3uyBP0dNjUQ6QY69feyRQf7D7yWpmX33D8f2NyO6If
7VwY30WpsGKX2DgMJdva3hyNmWQY6H78Toawm5oz6jgrGvPggqpad+Fbi4rXbLGS
x6VcoJhKA6pUeQkxw6pZ4IkNLyEWQ629FpFR3cntYkeH3CyrcPAEC6U36Mu5+v8h
E2CFUAR1u0pdEni+vOQfRhLGI1J6K32Khu+KEPzEXxyNrneQlTycwHua31WwCT1U
RuD8YwGxYuFgc7cKOrx2Av0la7TgVXGtg+PjFUpFDoJpLx2G7IJoEKZLsq7fIJZ4
+x4KgQ/c2K5prGb7wsLmwbxN2V+E4go2GJYOxl/Z/x28ROZ62ozuvtv+Rce9qzlq
qHzi+lOgUPb0PDYlPei+xsL97gqoGXjIjhu7sxdHqbh322pFqc/tDqgfTuuQhgdT
jVXjXbvi3BKOPHIoieRw7kt0h8rodqlgChV+oCj3KRkneCsRZonqP5WsYc346cIq
eWiwNMMW+nTebmEWf+NUjKUjJRhClYB0XuVRlKK7udgPr8F8uHWqJ3kuIfw9Ck8G
UeDkXxor3OV4sOyjljZj6nmV0CmIlq6mLVk143OLg5wqqpeVHQC0dIflSwfjtbOk
25JB1Snz/XBQAfO+rB6W+p61jsG9RHugM/+V89mUYiev0us61mqfZBRx9aGGYLaD
JHv8wU/Q+9Pd8vq7Do3uoX+cs5npGGjyjGOpMtA+1EGgFMvqyXfaSvpL4uplZMwH
Mi20sW73VPkwYG/m77duFXAnE3By7fnQeU0biSAxpzrWtbm1heU915NSvLNFkuwJ
EoKhqn04Fjn1HXQ3SdX0lmgGrznxU9gHNjOxlg+ErFibwId952ZnLZfI9pn36yCM
ZE/DgPWjoRaMOo8WLGYKA+cAgCMwoqDew5mcg36Yw9D9Jan/lMwYePiclsSyihIG
BHOfopOHpSn7IccONbjHRCLlEs0JOjzIuILgd6o0RbRYLUpVFQtCxaxOpCqljRGo
eZe+IX4SBFrhtrHIfR1SCVUSzSlFb3RGxSbUel7TodYCECl04ICjgTJBmzsR2XtN
EKmglKK0i5XhRNhvGVWKgCbInqRumume44b61HDcc3Yr4ScjqwGQGsDY4USyWQOq
P0aRwdrfJqhPBNGp8lxg8mOMPdsprB1FjttJE9rwA6KJ34/Mz099FF2B/fZTMAil
RmBIFk+HJx0/idsqIdLDvx1IitkPgs/gop9n0OZnVfb97gG/Nwos6xeNfdW4HnWj
VguE4LnuNEKi562UDoIeFY31aBrt+O1AFgtGFCabvpKrBRSc+OI7c/QJpN5FKxLn
+6ueVuogRdl79mhIqzyRVETKKUTNc5G3LYd9x+8V1ZkyW3P6aDYG3sPZ7GdH+GaD
SkwmQvzLNU05w2qd0e4JeKcHOUq4tkoDojEfN7Ayy12iqjwm2dTBoHslFMYW0qS/
KYnIQr8tcvqB7hpfRR7+AMoyUcxpWilUVdThAsb9xfDttw6jr1qir49PC3EUge44
28x2G9AMyenK7u2iIEkNi4GUZ1z56SdE21JLmM+qSaNYT81KbSU5C1yrnsJnjFJC
3+dBeQCl7z0LTwBChIN3YTASqP+3Agy2h3eAeHjZZik0XvOL/l61sHupohc+diYJ
yIM0Vo6BoaGAGgumnYgnKYVpA1mlseVHnu1O+o9ddgWX5YCV9Y1giDtd4OF9OvGI
VKdfHBI1chy5PjCVCc/hT30pwNg/gY9fhKi/FdFvDrdEei4we+xRv6AV0pw9lvSI
ULsZ8MH/ycRnqw7zjawjKnXPEbDLPF7TtbU2bVOhvblPdNGwnaGp4QKMjDpnHeiR
PU7Oi9EBszBEVMQpxbu2P9Qv+6wEBLg5SJm7aoDfla/ipZicXvsMRdS0yneGYsxe
jSxYsKc2B8C/33DmXwXGM9MaduKVctPRvtfmzCTyfjspyXEsVHVEg2lGAF83PRVZ
hBI3yZQW7mih7s8oE48Ufo2dJnezZv9fSzZ7E8HoqMg2rRRaaxOF3cGexmbGu+7f
TeAFgtAytukyiqffE51VDOG4IXmGwa4qTHHgm+/DG7Jm+w6OMgL/Jwu+6YW/hX9t
XnK4JP6bCypmgO+HmDd0PMVNU2Qvg3GKn/D8+clkwpc+RCizbnxu1ZVP4LdAlCof
UW5TYs+rQM4ElgM8L7d5UnXbyPHUPBpcd0ksXsOBLs8jz9wYrJw56z86GlMQ9D+y
tQjZrUMarjc+oIHylxk6jkesCbYgWxo+Z4AR7RjAreFXyjY9OSnBROL2xJE6SJ9I
9yI5Usr+l8qE3UdYFkVibhtqXFoa17kMbOK6KizQs6s25beTw6a2UXk/Qm/da/Tk
1I1N4Kk/nFLArp5j/k+LxomLPRKlQrp2zSEiaPsQ5kOzEaKEzFpek6SYSFtXDHjy
O2o4Qm4Xk8ayJXlKoxKHZQhTGHQuX5fiy4O36vPjdFRKur1ldjTTxka4CxivLbkd
974qoMjTAQgn6ZZP76k2ea12+qC8ktg9KMUKwHrGsTQYVnr9ShmfrZEilOKViN55
4RlYz6G4Rg6cEywGPfe4MLBH7bi0bh3G8y5BAYoqXky/eR7F9KmEgtgSzhS+cVve
vCK8bUsPlsBBxObmdc4AyqqtFZNwT9PP1q2V/6LzdZuRSISH/rmBrp78gzXg1a0B
460tS94gGw9WM1K/vo5oRwJqWWzfNqnYgIgGW+kavHo6aKgVuNaW77ZUwAhKWDe/
v4oCz5wNB9ppQEx5+dCQNVAD7k9ze5DJj/xM9RgoyXR5PKa1dip/99+c/t5ZXv8+
bjLnNd5b5isEkWRl8aMhHB/z/VU16n7mrz7isInaOcoBiNvB4DUx33jJ+xu0jYN0
4BFE/L4Q8x02xmOwe4x/A/6X99fBSZsY3ccY8aIbe2V1m8FYZtdxw57nZCYiUJU4
vP1+OkHPA9vF3/M0hE8uUyCqt7oFt5fJDG0Xo8WidogHmnd57VHOdJPOhCHoPoTc
df6FG46+TKAb6YR4yWUCNmNkKwwlaAaaro0Opgxf5ZnHv7u40KKAxEfSe+lR0DIz
d4uI0uKRfVNqo8J39iGsJUqulPeJ/GytggpySGhevdtmERXVw8UD0vPhdDuBW8UT
ycw33KfaGLqoSQkkT3aR99E00/qs1/I4HvbSvi56gXui+5xC1Lp7L9UnRBrlzrMc
GGUsAaWb9v0NcacP9DRdCG7FHmTg3ujYPPe8t1ENbe3AANSWXBy2K+IHfm2+aHOY
MJTNciWoOWRCo5SBI7EX2WNrIw2qXXodhPa5+KymIrM8ZpiccsKudVnQ0ANktVyo
k91AF2yR9/PoO0dzuB6u5Mb+ioxBwCS4uDjd59zuoyiLgy6/abFnBqStmnIdntPt
moP0f/Sj5dWl3VCtdm53LOYmOSsE2TWc8TtFgqdJP6A3eB8lY8V1bHQdoP50hFz9
4y03eF+hgR0e/U00rWyL/V8ZVtWDTGwF5e+/wl5BvAjZYCd5ZVreZUEgzI+BIp4Z
42hSWYIxgayhXk/Trez3CIJT8IFjjV3zAWbG3/dxe0nf+IZ1FfmJYAOT+WrM3tNJ
54ULfxV89Nh+fe+jfoXAD8RQ1mKDR4b5v/8KYyhPgSFipXnYv4wGWXYL3QslN2hz
NciDV+iwY29cnzxk3F1dmged/o4q/t24X2pNgpE+5S6/LFFIUrt2uBDtwZleTqhh
7oEV6c+hCBTE0OzFWYCFX9YiGaWw0B0EeTQ/TGgpcejU8l30y++QZu9PkmOp2RQ6
bHgxaBzaFJd9Gv8tKvS9xpfAp7qKCRdhCzDbOimULX7+WHiMf0NHGMNJZnCOJek/
fy2m/LtFVvfuGi25U11co1Z/wxAak7z2Fr3tZS+YxPBIl+qtNf51SncS53A7DK8e
2/OCtXa4TE8BahlxHRXPvidsAb/RiHG1oy5ioOyUvh2HnPn1o/9OlaMK1TCgXC8C
KX3an8yzMO60tXq+jsGSQMpu8MrzFVq0A9ymoHNJJG2JyT2cZp9kfAESHZVqCh6r
VehYH/3tKtufdaufQIPDMDjJC1Xtow7Hz8czc11Qlk8JRFPrefEqGuAlpmgsYgdW
a3xK7Pnm/ZHpOaqwhJoCTZZzmE9PDNDq2BH8RcOkShlGZJ2NzmS7aSwiugtxp5pP
DrJmLoGhgQld1ZtFv1AJnQSrfjsI7P4SpbncvTgQcqy63ms0/6+veXoEzSlqyN41
FPiYOdOyekVGzzdhHiYO9f5SXspUkTPxXu47smt3QWHCje/nDHMQ78w2I+5OWJu3
oP5EObjrky0i2uekuNCXGBZdbwMTYV3ephIrNmSQp8BOFomnsatfbLhOF76+hRUU
bC7ITaz2hfLp0tvAaNo3f24IIO2CBhCTLTaNS/vcxbomHTYfkJOeWQCUIbZfHOx9
BHHKgDK5CjakxFVAy/ZAKlggQRmRQzPrPrDCGwqgvCrZiUWMFPipyS20wkZB59Gm
coezPeh4BnzcU22TpRoqLAnorBLXFXaQpKkJYVnXRIPanSJweLaKvwBDMjGkKAis
uZ75plDpnFvFBuEzFMSVfT7Bzcq7t7Mzw56y7vvM5QEPGkfGSOlwWSN4vwH/kUqw
MwN76CP5OxZ6AQcx0WNGgbMnKMUAaGOQM+lnqsTsY7pHNu0y3tYYqlBSIx2l9mTi
kkFLofdk4I9zQKMftbQiDi+Ld8imf1givOr3kVD5RYUsbgp4fwGoK/fAme8+Uc3T
h7YquYkBFdSgq6RSMGGwwmW6/ECFj2wNHCnL/u3uLhpKaxnNZQN121Ojm0mBh4Ll
ZgiREkulWBurl853uleS48Gk+KXSEHEFXpf4OzVklvBpQanxxb6UU1Sz2b14QR4p
mOE9HoLSWq0A92jbGYtxsHAvNAU/vV9oFeQfZtn+D3bmte65AhHlmZryzBge8ZKm
xv3JekaUPFotLLKEUPxsxVduojVPThzg5toZoRbsHWDtpM3xXvg49plipGVuwdXP
XoUlsl6l5JqdnAzHEDrZy3UFBsPTplT4xTb8i74i2iczdVvUbH2KkuAHMSnFRpof
qexdtAsALhPVaT7xsJSISSkZtzuc16EM1CNAJii8hToACvfJIp0RCjSOISvvIOLz
jPq+rwMjmfYxwB/re7XfHMWz02O49SPpbTBQDlG7P/kUIY+k7Wf9nXCYsRizawja
GiB+6feBzmvL1y5lZsOUrE9I7Pmtsezd2CKa8wTOsxtKR9UOMf4/G1F3O63LOtCR
BaHfUplx92n8oPEtbwMuhXV2wTQSTwMteYQ12ROtcn/H/JQnziCFFYsf5eAbEGhE
VpwJRrYSeSPHQq/Jp34NwhY4/Ngrnr7DQ6dn+VmuRpwfgOXQX5pmIXBL7L9U8Qyc
x46VDVHtuRqzfRzQ5cyCF+HkSZ6UdDlrV/fwcfLV3y2Z1+1Xvr62i23mbG9Ekhix
cyXDVwlvYBnK6udm36/UajVKDSeku94Ky3nylsLKj7wQLDbqE9rr6ars7dF1BrXS
5CUSoHRfTDfQ7dwPUQ7GJZJHyFymcro7i+RNbWvqgO3+VEImtB3rEHL+sCZYoo/c
DpB0UGbth5bSNcXaBiCFLcKlmB4zN6Wd8OPa0NT3F3DQgdmXOUEsMWnAv280xbmx
rRJ61ATuPhMVCJRPhv/px2/zKwa9mwkgbfVEzqVXJZKT9qD91wjD6G+EsZQ17jR6
Xke6a0MMKk7y7bLbfB3aKCAle/oruLW4eG/Mdh4BK7b2kNkMvOyBWAth3kAVdtTE
8C8JjsdUMvonggtZD0HLivbrfXh/0vsu/q2+Ss0Li7bYQ81aYRuCALRWJ93ORISq
BQhhNVV9QaSbieJmx/Fb0MSQEIkxHiB6HBgHTyP5E1cOXmq34xelkBMrEvP9ld6+
BNY9RogOr8v1K+JSGZaSvS1Davm5RqoxVSW3fNsDKs8Y1kySwLz0RaTswwEdx638
gYQHGvo4ImEG4w72cPZv2LbObaAplog0DHVz/FS1lffIic93GQqJ0leUWypeSwrI
14v51s4XQxT6gAZsPR7qduh6E597LhJDGr0MCv4lubp+XiQvz2FjeuVdESK9jKCN
CoRsstpQ/ySzAa2cPyFH5KlgoXShbLQbuymVSIh34cqI1KVmN6ywr7zteh44V1np
oHg/v/WX8cs+QLiHjqp55tGaDoH9F67tTVCa97hQg455+5uVqkk/g77C5j7XbcDW
08bKZ7QfHa5dUmrAzO6H0mgVRk2R/OcP0s9X+TJgx1JYeEReEajLMAMd5pwZrECh
K7ahjr2qk3KRbenA7G7jsaOAfPw52ZpzDhoo73l2TBZ7fa+UZ08TDnYGLmRtjzM5
MiqKjcPHuBhcUPS5GNhX808XX2EOEbHdAdpLit5r3+CyRkrwogBlxGplG52P1Dh8
XwJkFPMLUJmVS7juB7/JkfPk2+OvNHB1hw9HIGFjO+Sq1PrB+ABJTV9BHGxrE0IZ
fXDdSh9w0Da9qDGh805V1nPETHnTfxD/vKnzNPOBw4YCIffDn5IZaeiW5zjUc+G0
2rxmhVbw1s6AOX/9lrJ9TXTrHncyaBLdvlIhnVRsevp58CII5/VRGrtXei205qiv
6litJJiH62Zqd6KXMMQ3rSFtU3Fyn9TL5rVQvhkEhfCDO0l+687djpIDCAU2Dyd9
AdULDl1rcModYAi/Kc/VV2r/WoTcOSD15UlBtIpaMSLm93/3X1Ye8KxWyLoDCYue
t0MAXuOQqkPspjLEO3U3qP1YBa3MNslb419BhbPQImUeWOYCoQ/t0Q9o04fZszYI
IRZOfe4hTYsC/D0GMIuiNb0aEmrzGAnoz2P6f1T8JsnKmSIb+YX5TsEOD+xnc2ah
sKUgjkuivGq1cmJZdol99z5xZjLkMgJp3tfNlkc1n/p2U72CgoWdfQy8zUlEgp3q
Kmnbd0vn3J3I+08nhmVsvz/YVxbWc4kRj8k7gZBDQt4w5iyEzhJAWHzCkS/l0lT7
eI0LynhF5t/AbT71Xkb57FG5dfF0D6EOOYE8n1yDn0sqDTp24owcBJhoxc9iQQ+y
VRYFU0XQyWspHu/G1vjg4kSTTO+x+X4C7SgYhRuIwjyqOOWQCQ4fqGJeU1dlbG5l
gjSuxBmOfkZNpiX4oC2wf7Dy8Xx0RW1crQdo5Az6ZPfiBqr6HpidMd+0qiW3XqmY
ENtdPSIgywTtHL3QvX+6hix9ykQgih45kJ3DwcXQUyzXkOrEzRp16tduylhJEDyA
mt/hG8oDeIGoFuBaxvVHwMi24BfRKN+w2Qa70v4A+ATz3lEBozz+eV6TmfxTpuzr
L8kZ9+sVC7WS7UMs2LLfAMNIbvebuSyv6UZRLKfUyC/uQ6kAUj7n3BPgTL6JvTlW
/+M1J1balm/cHZr46GbIU8tdp9wcvjKae0QMCGw8+kG0zQ7m+gRmjST2Jw5mCCzS
XAwlbw/+d9eGr6ltib28qYdOgqb7BGIlMe8I8WyPgr5903KowU+kgqQYPGwpCFQk
rxOwfJ0qXfQraXHCgnPRgLz3F8sqMBcsrzMHCIN5jCKRKgy1cXP+2HB0OhjSoYCo
9WrymZIdi/hqZpl7W01kz1Krv9YFoKn/HRIwl7kU/ZpWXvU8CtGedWQ1UjEyQHfI
QFfDDhLahEpVmFuH1rC3onQ9WYZthGfCU7cKfNdd0Cu0wV++wqy3WWGE2sBMVT98
o9LvSVIbTgNrxKiJJ4PkePswcyInFyg+1qY5oz1RCO61bL1W5kskSr8dSH00NVSr
cwPmt0OHMGOa38F/0ATjSnYwp5vIkEBC/aCZMCTZZRAUr9tj/syjliCBkBW6hCrA
z7XrcQWxcdktaIT+gp8e6lt5E2rRs+vOzC/vFRwtkWbFBSv5KoPiOBUR01gTEr26
0Pnk7cOs75XW7fHFwGOajW/TcDHC70PGaZ1lN/Ch7M7s9sXWOKIxDRS/hfAT6YVw
8GDufPGVXF7nJJzZsob/JXG3gBRPDaHq9xzB6AFmWfXX4VRkVSEWB4XjBj6Org6V
s05rmjBolGOxpaCCfcKJWdOz6gcDmKwiMvCB8MRaFLwuwYZ7avrtbJcBePX+Pw12
tlCHQJLGyYR6vVIoPiMtB30S0Woir6QiATOzoq8um5cVufF5oTCvyQy0MgGwMvX1
QyeZ3t3TT84VWKaox6q7EvBGBcZ0oTKSt49l5vhpzNqFwV96TW9XVIa2voSPfSGa
EL+uVGB25820onKA3nV+OuwnCcACJN7eimxMb0uaAT3pX7NKoVfpyThi6p/SGcEM
c0T2bNJG7CmU0kDkIlUfSxwCF8uaiu1lXkakRoQLvGJOdeSL5YT/DLT3LDmNadzT
V1s+yk4A0YYHBCB4tXcyLj3cAVfx2kg0UZrPRhbrXC//gfqRKuvJagdZlhuJHd3V
gsfYen/UdXXPFJixOOatOraVdczi9QMr/zWYvdq48G0WoOTND7OgFtge6p/gEgGD
OyxawNV8m3ixCb/sa6FUJM6TOU2ArSAxFb2QA2UZwgK+pcD2tZaWSO/WPJRrxJeR
HKc+OHsvQiMY6FuLNtbZ13VkRihNsTKax5zk/5WJpJv7c8IA5rjC+hp/T/JN5XZW
7ObkbXiuVXrb4gbJ9fH+hmRBMXod+zrtMIinzreACBBU6/jFP3q6t6SM2J+5Bbpp
4gbuQ1hpWP5uzXEr68dpOXFGa+wS7vVa/zvnnYYPe6cNhNYs2AnL5Ag9rcadfm0q
k317/VwB83TkiSCDXo0ENjyUPizVCD6ATZKY6H7dI0aPoJp99V4am/TVFg+2qisq
FNm/THXwg9GyIc3inwYSszCcFmydvEdi1KeRYyH0Xasfaexqrnw+D/yGvCaigDdB
fkRPuPhSsTolrHuFSnd77i0Ox1huyDWYBEUWitcYqafIfSSWdN3XQmvKh4BHw8R8
XIwV3PEzxLRr1MJkdKHWjIAZVuvxcQTOAbWiBY/89uHq/+in/3avrkdaaOrAOqSZ
2yHoCZ8m/gN8tfMpAkfsqSy/5jfhHURP7+A4ust89BhWmh289zv2RjQnR0MpoI2C
LcC5O86cq8KpuXUJDhSnUfEaHQCaMJ8/wPpd3b8VJ1WpXuUg/vCnB2GoA8TpRzJz
ln0HxwpbIuRVj7ndA7BUmreeeL9ZhjC1jJjHswFMeKcUdhQlCChAfOH544uwQzQG
gi/OkX2Hu+nqKRff3UV6/gAj0UCkwl/c3lDfaamgonF1ulaEufqb1erHYBzeO21a
yV9ojvO0EgEVKZEOHOXScLlDV1Ia7Y3FPzxzFU5paESYp/5qzoTFAFTxsdF9GLgA
45G2h83Wy3yLt4HxNdp1j1I/2XPbLYicXvxhdQJjvHpeGPPwaq1IzRfB2Omgcuij
K90AjLkwIv3F9dcGSeZg/lVMmsvjciVMR6oFXhSQb0LDk0OcMkOCtAs6iArV3M5k
okjsJHEfetm7T/t9QTyJ1EQcdXUGWsahFGotcgtn/t0fP7QA2QVriE52AZFFFAag
BckbkbydDr4b6CjXAGl1hhGyVZbl1JNpFMwEy7B15krUxHrvfWbIhi9fn3ltGZKj
m/d0UGgK3IXW07EWKGcGbMe2vfUVA0F/YhcDMFReVOdfsktY4zVlOdQnt3zPySMh
WjgGfzk7HWoAaJFP5a6hX5bPD+keiNghjWnDUQm1ZYlPv0yOQ6T6fNSJEahYDgJo
JAnQT5lF6uv0u5y6HETo9PFuLGXsp82vM0zRxI5kH3E0ZewrgpJ6/X1jpNdWBl79
K/v7jK9o3EXbZdKIXjF+yK4Ips/9YkjJPtS7cPEMAwvrcXSjPbc0bsgUtH6JZ9EH
8WZ6SthuqOuq26P0geeUx3CX/CQKtwP8NE3PLYIZFe4Jg9jOkEGz0MPyTsn+HguB
gmXs3cV3aa0FJMzAxHzcjA4t5JmwPaTb9m9FHlht1uN9a+4XW5/xw9nCYBnUfLKO
TxI9fq8m54HY1bkh5zx9TJpR2ycMWju7n35BMzZEbk9rNu24CZiOBjy640cU+viE
mFyXAUygx92V0PZvSKHK442d7o/5j0RVgV1iCj1JELd1nq0764XQo2yZ4l2j3vo4
DPnyuTFf7pHtBVY+jWVU4yMSbMaOeJ5wnBzZk7VlFnQtNLZ92WORQFoSyttRbgMo
sh5IZBbFLjy81yhg5K61cbwjpCm8W0+zypoKiJwdNaeNdXbePb88LQuCNwXrovnR
7gY+2Bwz/GOY9CX/7SL9+xqL8UPD/rtUbsayn1lCuE6Ejtat7PdVakpqHRaF8zGY
G3EkasbwP7U39/sD8TW88j+V66qJgDMRN6XZSfhchXJKnqpsCp4VBslnBJeU1xCA
YkQA1MtAH9w2yxo/TNteHUk2l5Hx7sE7r3xqy/E8yxOm8nQe2WzTeWl4cNAvZ3I4
h1Bb5Oyb7fUh1T86eJAcVmP0cNjzIGh2HhhjB8lsAQFxw+U2ew7n5e+DMn+cnAZa
Jvv9oRq+gNKeJS6PtbLos6qaCjwPYE+3F5bW5x0WA/BNKCQP2u7mnkyLE7ew4h/I
jziMtoR/XrU0pMIESsh7eq/TAZKxAtOr8MbvC8cjI2rH800E+Zxx9mg2mq42p1EZ
GTcMhNfLsBYxWVbkpJllWYDvRnf1dfQkGrnQ/ABe3iy8+LNHXEUKgGoVkBpxfjGD
9+piH9W/ZmuR3d+yLiN8uNRBE9rwXJLNquA5SqJ9ZBjO5oGpyhfZrd4JFMjfA9Jz
nRqH3ERWmvHr5zVM0/gnZ509+bguMTZx8uFHdFy7ypuhHsfMO7fBRFnDquhGrGqD
b2H3YWvDPxq12LBC8X8CE3CaiHBNyORLDjmXphB4rPgr1FuO/slSkdiec3v0e/hR
esrAe8E8ZgfZxM0rzykB06AHqdjI0ub4ePtD151YNAASioUZuNx4ifVZmW2k+Q3d
lhFp3AxIt9EvGYEl33XdC4qXObJkc9Ws3WIL0t5fJWbbicpxQuMYb3/Okq4UACee
AeGICIl8uw+CxD9EccQxQsHn7tnSXPsaa88ZhLWKr6Qxtlr8EXuEfl+Chfmz6kTH
nt8NYjmZXNhT1UXLEi2Qlf7oLVUqZHFQGXYBwdsn7r4fukbemzXCPeWgjag7S2Ow
ifSjZMj+RD5KjkCppiUMf4xfbRc4zb0wUmm4mX8/YJdvQlnLuSDHX3w0DqWcOKPa
ZscBki2MZdt5GR0l0oLOAsvUVPidfRI9UaAbFKcu2yFPqoGl5Z1t3zfLWt8LL+Yz
IIJoHeHvqZeZNqJGEJwSVXJlal+UVaMJfYISetQLxOP+unj03ZwoNa4onOZzdz1G
ywaA7zQ5hYDTGLMFzgscwFrVoDDF+5/68W9hwDzh6n+1Hg7gYLDh43asrMxD3f7+
UUfOKbeSx65D9k5IAFosVQC4Nf9a0BR8aMRLAxMDM0N8x2W7jaqLbxHixImW8tFP
HLfk1ILsBjUAqFnzZ0lvl/dyHsblYplgQ/9ELkEr3HyPTXRG775qUPSwX5Y6g1vG
83DIf+Edz7O4Q+h/ULTsW/NibdwLv+aeVc7HHKgMCQP65tTSZdh/pPjOw5wFKS6Z
akRYToGnYz+mYogX2SxkWrwdwCwrRUrVmxdLltn9WIlPYH4kkm1ASePusZJezaAG
pYSzYX1UE9vpJQA6APSyb+LZa2l6OSU7J0hdybZHRWj6mBBdiSsIDtVSv+evktcY
B0E0wnm+TB+WCZwLXSjTaogq8I0zqm8O1L28YkZEN8QwruzCMXclmRwTHI73TsRW
aOnJ2ZHvNIhN8/Ay4rgfb1cDLyU+O+7nP/J8PjneKTE1MvegN5k41CrilMeeZSu6
k6MlgYjwR4beTrIHG8PD4NClFkuDaTPITdE6VGLirPO+rIpR1gFOx+jBosS9E4bN
gf20486CdGT15srVsDzKmFRulwSWF5xmfLfthU4JRNecOqdQGumgSb9gftlzl5Wi
9ptwPkLD/IXZ+dVuWE0IEB5ttelda3CmNdTuJZo6ABzg+BYo170va/ilkpQVOVUW
JQjaH0mABJBS7SeAUj7tzY/diXZqMwOSp5VTrKoaLcA4HyN+UvIJyehR+0X37DZY
Nx3IF1iHwdK9zhi6L15j3vogYDWEZDV02YO18X76WFwUtH5sUsaW3D/1pkwwl+eF
p3c4wkWuBUsm2gMu0yinqJu/Wf48HEpcxJ2+hhfQr5IExCqc/daN3ohtKN9bXXt/
SS5YPQPQmoKlasyOheKkl3m4MCrF9njuMQzVuM6zmW/xglTO6yHZHyg+PuHkdykt
kx5O5Dtrja8BpN69+N/gFvGdgYbIyf2fYPRjWRivelnUENBev49Pk7oA52llJmK6
glCZGTB196Kp2inMq7PxJNaGqCfO2QUGfDYPeAkP1jKeT9c7r4IxvemSrUV1tLI6
2dPAi13U3f/o6IAQueKyXtkkR+NcdHItvt/4x7eR1USXzyX3vXqZYdBKYP0q76Qe
MTBEBkpcBO/BoA4wXJTe9G7f6nVUSqoglaetXjfbiUeGdKiS9oGHUygux+EV/xVM
r4qH2ttuX4YybJqLOctRURIVAcXVfujQXDfU1x7nBcl5Q5ggNUEt6EY39E6iNH21
Lbi7QX7C0QnwrCw5q2SADq4oFmaoTWNdSPKinMa/wKozQYc+O+RgvL0PujxInKco
kLgR7xUUQUEdo+kcrF0WEJg5PmV7Z9iwfaG83Odam/yzzY2SibLitr4ldb9KVO9L
IH1c8EabKOTWWNkzNA63gIFBTZurLlRL+t1qWXiKWF8aAftbaVm+lShirMLiZxn1
6wkbAE/2MJc/qATdtNlBLNm5LK9oLyKG3dJJ/zD62jCFvxc6pSn0Ggee8HvRTRlx
xr44XyO7byxY1ZqWapXYKu7aFCdFGOetoY5fMrimIXRvVHzce+E7RV635TkKgDPy
liTDnzW7iSC2KRXoMhvUjp0WPzCa9q1TM5p7x3Y93HQ6t3ldf1wCWZsCrmR+KqtT
7EY9xvGrNJ0HYCjIr3keco/8eTKr0kNbnILNsG+YQHdt8SJxGwm/WuZuIGs7ZHn4
WgZYFuU82BUTiztz5OyXoE9oB+63lfNxAZOM0ceVdJZQkp43nxjEgzCGKpnl2LK7
IXL4aOP8ipw+8eAimEXgseOOZGi9GRveAPc8h+gZjhdlI04H8hVaz4hajX3BAPdF
3Vc1nD9pQZ0intPf7XWNZTcsNhCLiASkay2t+tcYWI1X/ka/8iolrjVWJu2fSes5
awVMqpJeXKNOVqSP8rkMzMbZtOSiuDhkYisz6QJdU4teLo7EtLIJaFvdx2qtlKvo
cl5W88fz27eDnjrow51O7hbq+ziU1PcRqfVvykpZnMwiYiVenV6uODbzzDudpEHp
BKdoVwHD0cCEK2a7ln423hcFlFqTCFUSF3BYs5+4R+Myn39aYeNTqAM9MWf/wERe
9fLxVkVS/ZlJNd23xqQH1IkQOBU3vIR9AYBjjRtlYqBk37K7a1+h968b601YmXbS
Vfkq1oemOjD6o87QG4wdwHXtuixlw2bQQSRIyfCZftcyo+issTM9Tn5L5pLeIML7
zeTPNCXyBqzhpRYoCXLjoDBO9PSA2fHLa3ItPnG44XRkJX3UDNS955eo2KW7fPtk
EXUSV5l0o8hwl8nvfsT+L6cOEPp2mXpMAfs92DOcH1Wr/o8XUy+dcFGpWKeq4oY2
6VF/05O8GB/P07uI7paEqrrUK5nDkjuVFojELm5+OdaIOkrfPR04pH6HaUm1QSYf
/I8PcZ5Q9mqjIKUPPvcXRyvHatzrf1YJBuMrRfGcn3kRCkKkQjcG3/dzmUY2R/Z3
o8oF3dBjGxAl5tcJWqW/zBMK0ISELVRm9QsUDGTSvJpU6nHEz0LUuhugj4owUu8H
M6dm08ywJy68x+5WRrxDrQoli7HyQ38LfPAuGtsSCsOEhvPktsjEEajsBikxc4Bj
ntDf/h3uXK4Fg9Xvp/E/7VyhNHA1+dE89ESPIbcgTbwfgj54hegVa4qd99blX+BX
ia7eenrMEWkhcNMqvMM8/wPZzbPl99SS5pp+5rtxpANMgZLYcSJsyEbJzmoQ9bYT
fkeDlOcCR3385R+U8hO+27RIpWH2cpP6Se8Y5wNvQFExREAdMTDXTlZQXAnCBabh
YmIEuIa7EMKJxEYMOHA7xUBevpW647gE2vL22nJgwhpViFei53B9DBSzFldp3tkl
7kW+hkoEOgd0g4hAQGsKAMJyIWDEp+ATheoBLm9Pz4GpGCNLw9iQbf7Sa1dRzNJq
WvNrMMChmua+cARCvy0D1VV1cHadt+7V8Sjk+JtqKVWzpKowGcHzdPnVcA6RcDxa
NN7vgOREg7ozYZ/kXW1xwrC3DYwEyDEYeV9IsMWxklWYgdlPY6bgNOjWBMiZCSCO
ZP8QTSqn8/ec6HWBJE5u06bhJOHXnz5fL0u3JFvTUu73uMnfTKXISZ9LhNRFRf2k
sHEbO1mhzYGGlqnMq6zdzyVuSn99GjaonqJyyu3Tjfn1kRDesk0ccBeTeGadF8wS
IQVeLJt7TmsIpE0pg+0XS61WWfU19H9nx//7M+QIyg7Ww/8sG2pqslS//LJkiYig
5KMcDDHI/OuUuhO8olF4bWowL1bb13lQ2K6qAOZDEhF2WEZ4sN2DXtfIls90hjBq
J6Soyua9rkdPI0O5WsFeQcRymMmVFF2EBYCE/kMGUlCmrWxoHRyYlQuGiXfoG96c
wgXkGTJ2vnsRztOoGoUx3chzDOtbSDt+O0IO6FRJ/do4ywwdxqgvdG1d7YOh+3QG
`protect end_protected