`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2128 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
h3mPGhLvpV4xDnoJxCkEpOu2JeOIfJyLEsE10MXC9aid57oJznYb0X2tHzZ8lNAF
/f4ahGCkvLv7sY9g5k7eO13IpJDKdaVKx+TpFRqzLupDbBzMiWoLyewsF2wuB4n4
OnSSu1fur9F3wel9beNLURTmPSmwED3jpWCobPR6STirCiw+SHQmUkGbI1sdBFil
nRRLFmqR8PBHz6kHc7P769au40IPhUJR+33l2q2LGynpC18v18Tg+do+aopQuIbE
AS2pPbpx+79bMv5GlNe6jhRQIwXQnpLiPBzBdqrnrN9BEPsaYKWYyetenBi++w4M
eA/W23GFmrrKlq/6E9RTJG/um33ZbQsk9EBxRbdG/G4y1pTYoqa3XzAOvKA+cwCL
sjzFLpMGHXnz8BB8OwkPHVu7ygX5BWNBcoaEpd04844Qo0MlVEUcs0YZwhpaPOTP
lTaG+j95H44HPsBtiGXzvqxscPQU2NAgreOdIFms5UUr4oaCchkAdNmuChdfSrZi
Ve2tY0hLGrZwRk/LRNcBHVohxxpDaYdZJdyx3zX1Wya7KlL1X5iEY3C8/WeQL80+
vMMHn2rPXfRSXcKBksNQOfWBOzx2skjbKO6rO4c0O7++Nq0zteaCoCZ8hIkeNkRg
Kp1UqoG6nnALCgBlUaRt/7mdzq1ja7iTGw2BpbcDh4AvZmjnYQ0Jp57zSc3lbr+M
kkGUuyLsjkMCy5lf5c0ggnjqgTS4p4A4VtwhHuGhoMtfMP7mohhQxSadWmmwdBTw
xzaTO6YMTPHwiMmM7lUS/L9rbOB5Zd3lantlht0X5uDw/XjkUGbFCk4fdXOF1Yuo
FzpgYSUtvoXOWoHgN9sAFIESNS2ucKc86WGwobNBO11K7MuCR9acl0MljxllcjxL
Na7Hza3/aptV6p5Km9c50FK5EfXdsaRJrrR/Tjl16jEjJ/ZgMu2CsPjyfTZokEBj
9QIHlMIorg7nEDgyDTCiQ4xLAsCTHSNVo16e9hkktD+6hOrsx40jnub27OQJtB+Z
8knD5UP1O0E92UBTlkLXchH4RNWntY+nXmRqPtK8PSLy/Dwr82hpZ4YmP8eFgIO9
eYToroScvKQfGROcymajHY7IJJDpjeoXXDotP0iy/tUEq+CmA0r3oLqtjUp1UrP5
HSc2jJLQ5oThh191F6yAe+wQH85WVkQ+VU9p85fSOGE57TIlWD1nRfAmpr9kGIJV
SQkIjU2dg84vgNBciPxmjkpM4l6sOyU66A8jTSaiGTk68N5/1Yr1uAMyqhjP0PGo
1cDt1S80eqs1Ysdfs+Kk3EoGabKczzDYGVS2tW9XcXDFQW01WeFC1PNBW4eOEjlz
9QNQSVjPLOQztz7XFgQ9psc+bDZplzY/ftYir1lVJ++PiV1IQBj9fFWtY3N4lWQa
AzTKnOUhdyTil+rPgnJOAytffLUWZbjpl35us0ErDUQzxtU+M4q/2qJTgX9yKj5/
KHripi60orctLVUY6TOKvsINZPI+uSov4PnJmb7cLxHb+NO3+dTBjqQ9qWVyU41+
0n+D0Gzcc+vwlUUQ/wlX6Xa9VsBhUX9kBwrLeCx8otEBl4tXIv9Bq9P66l2SlzO7
4+0Jzp44Q+jWOD3hs6/mPVq0idl0cOE7YtD4eP3QHBSWXgqRcnYqczdgK6O2PoQx
QDhKp1R+6U/mG9LyGvv3cUV0ADl8AncfOy9b0tGa3d1LsL62zXNtqlcUq1ndMARw
+YAxKVbRIxQjGL6N2i2sOWYWQGk07LE4tSXnxfVASSdbr/ZvjK23vD6vsKqu3smt
7YM4UjWC07qKXZHXTs79SmIEM7ho4KaeHMjUHkfgODUyWzTRtPGtXPw481iI5cua
dM5Gw8vjQgSlTUqGN1RUwCH1Z5n1ZS6OVvuJiuqFU8qDpoSzVpo1k5qEMLLt6L0S
E6jVlF25fhwwpmNkGnKNoWEWkK2TO31Wya2mamTTOy+utxtrSKA7hC58566QO99V
3IdOjaRzAgMwaCP2M/bANz6wNS7gzOqswHLxjfiBrfvvPlXHWD9DsYQJZTMdbVAu
wmyi+QzmMQ/VMH86K5bSI42yfQ/519i+yegkbcTLx1McNblQwrIumFtAg89WOZVT
Wld9ww/zS6VwxH1DMC+jAGR40yOSyoQjjmwo/MSQ6Yvu0rT6nwQWP3WvUYnaRZdH
2+HUQiM+SY2ot8xl60jt8LzNKIbOIhA28hoeYfrqV/H1TUIwQkjVsQyE84+YQq4l
3UUspL2rdm3iyIB3e7GbvpE7Lzb5m+YsReanV0sC0WmK2kCaGhpd5FdMcpa1snsj
OCbZFbWeL+3ZVxmTRJ/z09u8xFm2b+84CGk9kqUgSshSKJGpieKiPmp7rceXgF/c
rR7b8L3hPJAkA03DOKPq4JxV/74zFU6FELUrtpcHl7hy+oOpeQcrDZDgomXra8wU
JQwWaRXGVlESXCT3lLgxt5FLH6kDuqKHjGg0QN/Dc00Nl09lHpjn1mkeVzX1ZvQf
807QqZHxwwOe08x+h1M6wAprZ7eBQjh8gfVXYsFZIN2oj7BKLI6iKorsoWGQ7Lcj
nsewM9JKMPOvT1w5sZvep9kiTXmBP9IX7sxcsEMBlQAsD8v8kzWoTmgJ6jIwIeS7
bFm48eUhEWSsGYqhT9nEZTiO76lENQ6fxcee1FePAe4pzr68SgWLAPvgqzn/8l+V
t3D6V4cgcc5peGR9K5WVgg==
`protect end_protected