`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4128 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
qsE8RajP9HKljDY6ykP5IPzU5Y3kHMrP6Nsv92RcCuhuWN7pxkdxCg4Za9rc79/Z
QO9oNlzSva/+6Yg9yTRhx8CDz6KnfbJCyn8UHe0ennekiT2OWgb2uxQA6om8uAhP
PHjjqMx7F+AJoW0n5Xyr6cVzqig9i/UhFkOaay8zWCzjNOuLWdjBZUo4Z5xDsauh
x7+sA7kVqD1aorx8xxKVImL/FZT5XQ0DxFBex5RnWHKoyh9o774CbrJ5vFK7K23/
zFE7JuCdrkIhsaXQt8rpGYaUc6tKWMYd5NWB0qPihiFQTOpvKi6kHtC1WPGNwHAD
j1+lrBHpOUdQIjXrHkc68lxxL1GxP+N+IcMGwg4s/+oGdAIpO4ZBh4lANP/6Yv3I
bMVKaPFXJ1Xe5gHOIBUe3jl2KP0MfH1ppfEYCUiV6SlMzOD0adg4BWnaXcoDJgIX
64aNlqdU7jZfKNbFZoXrXm0lQprH6q8wJrkOXWXvvvmt3T45OQFqPOHhmOCZns1g
jLlQVg9FRcJ88TF9DrihyqIjhZwuzwVlKOcPKpOCxpGxPfDJ0Y0kNvZiePW060z8
0KNVTvdYJKj+20iv62zvGRkiPb7I+8NpOBJSQsP21GTcx6yhGfM+AQxdQmcP47OO
tbfnU2gFIs0TpFHJftHzF/bLZuDy3RkKF5rOGdKuefB4IW2liMJuWiQchyAdtizf
C1eJRIQIf2ne3DiZ9C4o9QaBiXU8V1bCTTEPiEMjl6jQZHroCio7tUD/QB1VS/L9
SZLsNH4iOgE6mJXQ9oT3ycs1crpfrAMWk9+G41JyavYP63nnRsjdChRdr3LGzDHE
b5WlOfG6OGhKbfpSNcdiPnww9Gr/PFvhkmNNy/rx8aCvGm4ja81Hpn9V4ft7QKXE
NcKQq56wdkiSRpIthN/uP2IqniGpT9Es3Z9qLFlifQUyblOkmqwV/UwS0/zaJDKc
pKfjCoD4GsnGqhh0fAwc/HwesezEjvDWEPJVhAmW93BsgWe34xrDiRwoT9GmZdiz
wxw7KDAGumLjoQj/x4K+t89rTqAszj1Hg31SceGwtZcp9dqrvgibqojKnTcliWvB
qQSf3axpfT+S9IcYiQBga5T5nn7wJN4srGACFlzOgDyFY6HFxThJCX+n+NXQoxoR
O814k+yWlHeVwPvarSq34g9GMwX93B85ADvzFD5dqz3LmQK0OydKvqWWi4wp5Sd/
RMR5j/jIS1I45IYFck6flItQSS1aUQiFEMN8MdaBCkGqAbDmHFY88HbAc1st1i4b
cpT0zSkqqqN0eax4N7CF2/I60lD3RHNGPyD7M8GmI1Sy2VLjiC8gk0/AwKjLCpHo
3KFvRb/3wf14ZDe9Kza1HUnG5uVTkvbmv1l09qHzqVujk6cZA3jfDRGy5F2r5DzJ
nVVJkNpXd+aA85uz3Tp6Y3uLxTbun+bURD67tgMtf6ay0WoVeu39NsrddiPsMHDJ
0Sou4oEkLFNLjT4BKaow8f8PlwlEmd6bedXqs7D1uRu6l4sto7JOM9YTAzdqmjWO
xYaF3ZPKAyJVnaCcHMIwu8KPmAlIV98Zj3qKz6orq32BZMW1hEqbVVjbICD22LLo
/1QDCsUmu+j71teCQducPEYJCCX9zMkc1G56cKUojSfWDNd0f6mkGaNLpLK+jVWl
r2KcANhQ/DwKofd+XkJxF86Yl9cWpnXHY5TkUlL2czgLzU3mKyELotE2fI7NtRTY
jMOSMr6Vtj4R6S7fKaYMKIa7CjZrDZ9zgyzuH7jEav+xfdF65f89GXv8LEua1mON
CqBQ+Sss6HbWzrwXQy9K0Cy3LN5BP8uugsR06QP/StrB12t0LDkFcP+wA6sI+zJZ
Ja8INcTlytQKurCIUOKChUyDCq18BFrlHu7MsTH4P6xl7Qngrd/20ri3SLveht2w
M3W+Yn+lNydbEvyOHX30RyeOC0AMY7Q4twsRBymy8v16iU1NLICZqtp/2WP5Jl+v
Aj5n3Qd+vfQRLgn6fW/swfxT4kb/KYf4TPy7J1Bb/h96gRYQpLkqmUTXULyBJm90
hSxeXsMwMjxkZolujXTvviGg6zHcfrZ/3Rz0Lf/Bybny1MfDmRJBGCjSLzRGko0J
CxdhMm87FAEXgT96nMTXURNVNhJjS0EofjIX9htdqUcSref01O+wjwkMuERNuSqy
WJCbP0aUGq33j+mE98ka9reNAwZTC/6QWBQQxuQSZcjFe0vadG+jKLlolzuPRvnN
q0Kzh6hAYiTrr7tVjYg+gIL+E7PftICTmnYW373b4Y46go2SlmMFUxjCWSm6kjFS
k6O+/ECWxwNtE0NxHu5CToeFXZXIQctfKO0brDnTj0i9rrBd+RhbWy56yyQbCGeP
0AJGR0BMi++nCVxy6WQh71HML/xwYfxkHqYRu5IbM75otofDccNzfZ/OlAzKKCsX
QBD+Unk8l5lHlH5SvCtspGr87nNm0Pb2caWb2PA7okO651PtiaeJh4WV1MdCPfFC
Udqc6nMk0FozhP9Bqf08GNcu6zD0QD4cgTsEcwHBsmvsDfxboy71UTaONsKtZV0b
NumRarzntxyJ8oiLNX4qEr4Lo/2/tLXPbYzi28XZj7FisZc2w/0B+8fjGN1vNoFQ
uEcoAcXPViyMkzTa9j17M/hwo0CBjq3b/KsMZewYMhfsWh1ns23vcwSgQ4edz/B4
w2CimS9SBWHAR3DimdxrjBax3cjagZWUBQk+ygJhjGiQCA2tG/9VYXKLOFn2hVYq
9IyRzs0x9/ZKAERgn1flCWMiZQiLz5rl/W59RL3F1O6us1MA2qmzBZRFd9kx8zs8
DfWPKJf7dCJswYytWW7hI5mmU5rC+N+adyDpCHpYjQasfwm0AfB+hGeGb0341x8u
/P8bi0nIbD0dTIYP4kwmtTdJWf9tAPfut71pMONv2aPgzUVxOxl1tZ2MlhxlN/zp
lsj2MTPWMbm3N1C5wk2SW2vdr8ekKvtwsrdFzVFTSXIsaoHrTDhPaFIBzSScMh2Q
WUNhxhsQnE+mmThz0WgIf53/4uKGWc9DMkVSYOEEU6ERu4Sr/u0Q0wXutTMWdpYi
Nj1Z4zzwaUq2GXMApp4wNvJsj9AeJcTDvtRD71Qu2xi19WI0NctXmn4Z10MFnZ46
TAserHtz+oLQfn9OMS/gL+OBP93uPFuFIR2ydWhZcE/pzHLeOzhLYuKnzXnATEaO
V9IeEoTqU6bnbWSSbxhhqp6eyyBcpM7/egrpqjdui+VkJuNsK4MCxWKf1qSRVDB6
12ID5Vc4UMtJ8dnXPC/WsT1Sf/VEwrSqrpE/PIiD6RkKt27vbL18YWXLLUsSrzRG
ba4An6jduFBEIj0aMknjvOIm0VwwaWtRs6D7IbViEBW7YLBmCo2WGvu9zHtVa2gi
hkDtbO8usEdGIoaGiiOiZc8K6dZxUXjqc7v4LjJdNiFxZyQYQdN+M6pAkCaYknpA
OVZI28v8hpvFvpo/7bvfv6q2VAIulLnDCtoj9NsZjEQThYmZHFAFAmOzMBfD3/Tw
hgp7VHp3nSYYcP0pr1mfd3m9RC+G5N7HrpWuNd8LVXgdveO0xQ357adiADq/vtIv
mVDoYf5/IIHmo9nj/1bHvsvJmzrUv9uj0aaU6vd4Oczj5b64BDgenUAb/+fBHBU1
7TqJg/FSl1F/yQae1nNvs+6FrG7xME4gxtbL506TbRxl4MwXIKKpF20vsSAZAlKC
xQJXBRF+uWrlD9ZIEzTbsgbFSextL3jxPh7l+QuGG/a8dI1eg7oLZfczoHxK2KC0
vXzbn92MADuLecRpVnsN0rnCx5HXDQJf0MwfYJL2S47hJ5epL4nKl+WF//lJuL/f
o0c2NMks7A/ikVTHKMXhRwNLc+ORONphDFyxifna9COaMU7XOU9t1D/ewq2nJTN/
qLfvms0bBhZn+gDjUO9d2ufMu0oneTl1oaS/RtKR+Yilbwkcnqx7RaL+4GxClzfB
6OzXnENRVPdoLu3/gNsXXGYnGlKNapniqYq5Mqi5Yqr4XlsY2CO+RijEBTDjqqvY
daYIr2NAQXbntiMi/wv2rRNWfrs7hrGEPIoDMyIY28T4Ux2rgigqhyap9Pbu5P54
iaxJBWJQ26Dx0XiuhH4PhtCnefYG40F3dvDxArlZyzQ3CjA/WGQMhre1TQUbUDw8
eCxKdVJd2MPw6z+e/Evsu3vn0rR/vghtQbAe5aUoKe7Tf5I0OdwavmmvQHWckkgv
KZ/0dktW9wCNvrydPFbeqxm1IKRZkFIuYD9Ck9DTYo9j1F9vxO1BEu/+bOi/Ip+q
tpo0kt+Bt6HCSkWqDQmOhTUW1OKtxeMrq87xlXLBX1Nd5c8XFzwvHFQE5nhpbTah
6/NRbMeqQLd1uT2PnxpJm8X5OVe8p4zEvjFIjIlZZpFAHN1V43BOKqYzcfAD0oBg
Cf3XXS2k1sKckhoRTWMWKo41mmpWBo62ok5Oc0XN8aA+X3t0Hld57ko+Ui32lNHk
5519DkKhQ1iRmajn11jNfyWkx6EKR9cGWF0iHPbduwDXIvrvdf6klH5jicj0mwDz
SDXgFSBrNceH/DoIQ+JZ0J36iJ4WLipfUr0typL6Afjp150eITu37yRO7Rj4NbXc
vYw0z2O9AafjR92/FdSKTk3qR6NG0oC+t0BflHbgRY+WonSLFj/TlQ9MnyCyKzLb
sUlIQb8U3U4O39bzpLSFQHucD+LoxEoKFpkL2D64rHrT/uFw79LxhwE5fOedzpJF
wAWI1KteVbTjr/CXr4cf1/2rH552i0PBMVsHv7CuKzyfqELM0BD5uHZL/8GQ//te
mhEMVccU997yngXGhf9y9Z3JhvlFzUrHGPrpNq/Uyd/uN6cF+fGDBmt7ylvpNkaq
SF6uesvcWdjnTvmBbOlHfFYkVJ0AGax1RHR1Ku71OKrnm4zjyz5+dyMDJBJVqbBw
1SkcNWefeqH+fp03/6f/TihyPYPVy+878Tz8fEd5Zhw696IHfUr9aIDJCkuXAcE2
sOpCHzOQ31fszdlZtqr6jLJJHIC8IRHeuP+70RFwRhs+3ZAOfobqxdzKpalZKeWX
c74kJuBSm7yTfC1m+Y5Xl96YDpP0yMXAaJz78xefoRpgevpotOn4rhTlt1M4/Vj3
9M/cK8hWYJyKVAPR0UsBcLb1y3qaenrQBZ3DYAsjIy4kWEqKeWj9SFVZRcmyCQ4e
3Ar+edrtXsvZK4E8jOrkbB4Jj8zesYmQkCT/RKLmQXxpppJE/W0Pw08Z1lG4qPR/
aZ3/Z+0AQIPI5DH7stcoqlEw0XEWYjLU1fxK9LL5GVd2kQstlzoNtWgB02v1Hb4D
cSnq/homPsvguLPo6MQzypWagVeyFB4ZUEtDUwd53RdGwG3k2Aut5BUEEAEMJfIq
`protect end_protected