`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2096 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
OyGGrfLtuV/iB6oXYN0vYEmEIq5tvrx2MQQr2Jj5pPSXU/a72of/uvED9qXpBIho
EGre95ENWx3PsTlZiAMt4O+oLZ8bA9Vjeg1lujdSGS6sUR8waZi6i8V6JU3vOhEk
o6WM4zqvK2edGX+nm70B9e/KY+WWUejM+S/0dWZW0QlbSU4NgxSxqWXk2QJ0u/zC
jftsUy6Ac7Kenj/WzxqYh9TCgiKs2UkTb3PY86INMzd/Wc+r1FrGCMdxQVa9eGu9
5gWza/N1JrORz1oUJD0Upt1U64ZJ5LDNb5cHsQ8mCcZ+EC7XJ+tWrT6RvQo6fVMb
8xLP4YGYd9Pm9Tlm/Y4+HhiBRZhkXz6tvQh2Mxa89K8JNuFJZ9iL2hyoLVsuUySO
tu52eg3KzAQRwcN/ZxVFhjxrNz0jcJdgGoiSrQ5YnR0726jLisor1D2J0ExcHjq0
8QleC/jxI3AFXnSozFFv1i1rTNuuElLxfhh5mUhRsWIk01CS7msGQjMy8yFXcxUd
VpmEDbsobDgF6mg+dfuN87Ql+PU23RPU13nJg48RcVwx6gNO4tG/ZTfDdSoMtfXm
YNqVxBAsKMpxU05Io9fraU0XjXxFq2YCe/KMR/q0xoKmmnST2dTnVnvz+leuwSSX
Uti6xgFJD0jKr47H14QiaG3Mrkdu/Hf7jrNNO/mOMC/kVXjE/AOy4cFMFhWRGLIA
W+NstzjElmm/do5da7NW4bB7oqdi/WTuWgm8JlRfN/KMjT9TFQiD9XpvfmoA1aCe
8B4G7itYs74KHIjX6o/G5sg9/+/PNpa2ynK6BhjMtwYCZ6x5B5A7dTkV/YpYGc9u
Y+7yjEQREOa1fmKfPmlDwtUEkv1j/F7+J+ow6xsNwI2cOBm6zuadVoieOAQNIha0
LZ4lA1Y+W1ozZH10I4pnJJF8L77oe5Q1tK/fPWeEKA+z3SqEBv2qCovoxTQeKGav
+2j0adzQm+2tVcQv7/KC4WnHhf2QqnO1GWpLU2eXjcRJMbm3Ab/FAZ4YcYIw5DqU
MB2IfsMe4dbx+jmtZayHcVnswteK9LQ4C6eTkhhouM/e7EbkA1ltt+vAbLchwS8V
UrnCbYRArbOwq+2n0rN/QlQDrlsXt2rzOTxC/e+QMFoZVadooocedynurnWn+z/E
wkhbzaRyvn5/ko9dpWyq3CuRHADRb5hAjMMUbmT43pXyr6V5OYT8VXruWnr+PvWn
JMQcxwhEk3BMMvYxSjTlZDYSCSSDIDSmeVFDh4Iz96Q/BudgrM2SEDr9qHcj+WY+
XLOjtbDjC5BxbO9p99ojyemxGFrIJJVMEjKOQebPxbmR+i0VW7ltepflbFSgRWt0
Q4yecBbutyIy9b2aOuvYnYTPXmr/AMQbgZ7+QXBVskzAE5iWWG+Q5BDRfdtizSI+
xmehZKwttn3jMkpNny374lut4bG76B+3uqlwXipUHZlCYbAzM93wMmTcSBsf+R5A
Jl+5T2x2sPjra9LAKkjn4DS8gA71EWrDeDid5b666y+sYPxg6fk2vgDrN9d7NX4b
W7VMSfoZ28DeBnuqjAX7szBWoDsA691a6elguKr54yLsEFi2982JURYYgHief280
99o+GPT+cTvRbczS97UgGpo0TQAIV0m0HC8llFVIAa/cgHz9gThd5VRKxPcabix3
VN6YJEJHqSXOxActWLuZGitjEKTQ63uyF2BNBkx7Z7iNmQjqy7n/VlbXY8bOQ6MQ
6HTnbjbP0id1HFMX8uB6bujSfcHz+aTdcqzXBr9I3xMKfq8Co4ICOVheorBCZtFn
3IYkSMBpJqV5YlEO6oOmdua6xJyv10bbOEVgiTsSbwQB3JA2mXvNUWH+7tUgLVmd
kHwS9o0isa87uphS/J/wyaHzrVHe+WnL0iNxVO1AJdvolWcgd2uRHeI+fUVUt9Ci
7PLRKNLGNfboMuQS6pbsnilT4Un3PxRj2q6NBhFwJw+qBcVPPixFEQ6LGHSvJDzR
8WQSglIvISn3nhM4R4LwI15XjAHDSd1xJAHqtrRKmAK1ra25B9OTY3tRUn1DcDkA
c1DonXK3puF3cFsrp6J8+9wU1njxa7d8yvetM7Ag+Jv3EXQ331+VZKy/8s+utsCv
OIauQSYJ2UY+ghGVHdlZZZDZlsfhsO7bBCTqnxleaeJC2EaULm8fHjRPADmhcLZy
MZdCp48YLQ0kdjBLp3imT3D1JFY2SA2q2qGQz8P2KhS6g44shEPKwQHfZI3wtwZf
Xraa7ErZd7zTWDPrbMCfiubNy5gYHWWPSyFA3ocv98YIY9H5FR9HKH2FxWTfBo9T
wkFJBdemmTlcPD7tTV10T992KEbstbl/EVv603hXzce5f/tJZ2P8hHYH/5joO7fi
R+BvGm4oP9QzD5X3GyENfkcQlRRtC2zkB1qnSkfahz3TM/r9sGIjJxze2GumNKA0
dmQxwCf/JLv6EPDaoydug75uWdpufEB5G/5pGFUCifQPvJBx745oRxS3ctepoJ8I
v7KMNeL1s86sRsT1P4LLJG/oyhRZ/wYuVyjpZjsvlYAkvXlB1DU642f1JDkQMhbv
MHj1AQF3jxnwCsiseEOgx1nptVZRhtubK/nW8b7WPEFMNB5JYK5e+Kim/UzMFpgp
7KHUl6VZSBejm5V2yyYgqUnbnRwxZwK8cKbvwBCzxs4=
`protect end_protected