`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9776 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
HdytKcppDjja7VfYQkCqvErsQFgfl5rfcGO6C2E2kNFDrsbvZyG0b+Nizs+4OZdO
ok7H9x7sYyGV92a3vQK6FaMyjEGMWRX5gI8dOSp0Sd9uJKQ45HyYBmQu9arUwAZl
I7Q41f4Hs1MlFi0B2EJfAx23O4/K4+JiTWUo+7CwIGPdvDM+JSQZ9LauhBzgNekS
8XZCC8lpnvItmUwnA6PrKqyX13Ktyk5KfRl/Psokv0aAmoA7rc2jpVzaqx0RzoBH
5nxY/7OyNlnFi+QDGlr1eXyKtZHcEcM1VJvTKInAKMetXo81jmQw9M3I8GluuTu2
mbq1zowqhjuGyJCKVk6MRHVpx5j3UqMw8/ZlzBrwRG3zF93pQOUrJp+G7lUkvU+a
lrz1He9xXm+ymXy6jc29XQnpBnZT2ihi/Oq+lU0CzhsI7PVE8N7bwZDi/rHGFHeC
mR3wAcwmDwcVH4YwfTiqDEMrhRaenOvXvCulHZz8jEdShznZv04LH1LfO4ow+s0J
whYRlbiVcW8nh2DxBT2+xRQNr7aN1h36JTC5d68eGJGpfR5qygmGzAENc7LGxj7d
MsPVEvVS8v6QH7MnHPxBcO2XWBgbLDZSwthUMjxMyH73LzyKds4uHf5sG/i08asT
cgKbA1zmbdiSkVys6YQcqLK23ouw2ocpM3qZY49xyBY0MNZlYInNNz5CvgTn1za4
p+ykmUbpqw6tGXM5doIrYXIu2dCS3FiOMPDmXeKuuuMkupP6sGjY6/duDvbWAt3h
aUunLm9KsX1QyfkBqRlThFafSlAyU1pvM/ZDLeeST9mvcOKJEVU2jNL+UV9sPpn8
6Tf8v+DX+eI658t4s5sW0lSGV5Jat7fjp4lSA03SMV19rE1zmwFXiNRD/aJTBMKG
6tENTL1Y6JBc5RdmLSXYdxywMvw6XRWWf1krrglfPj/qfKxBh0QYuOjJH8ekVWtJ
TddK/d5QXd5oJ62htqA0mhysZk2X5hAVIjxyPL98lSppUOB5XdRuUqzmOZmQJOWL
ii4o5WLGbwdC0mRLQepf4q+p3Q+PTYa0irKX/9gOcIaavuzKlIGDyMtXgPEL7Aaw
lE/1/xIsRcklYXMIBl6ycRDxxv6w4V0gYXG6msGBnA4XKapBBpJMMmWC15OFmc2m
miIZ1fa7gHKn1d0qTD3HLhJ+3GbOqlReKB8uybn+Sd9T7en3ZKlltFxfolev3VPt
nGbx5aBTn60HmqLbh21lKixTqkL+7dJHoDJ7i/09Orxil7dIlE8MQhMz9oRIuE+N
/flS3k/KxkASv0cAMlVrLLfeP6B4DG2EahfZ248749LvRRhHWZ16OGtCk2Yaa4a+
STJ89CFd2Z+zk/38jN4yAoTyqtGspN1HD7U7bpL80ljfmmq4gGJSnZBWMlzUabFf
v+h9ZhIFjIUenQKimcufHcYhazb0azdwJHMOOY2aomk/8kOaZPoCl72b4mNfRNhL
MtzIzInZ+9U1+cJ2CJye94+RsQ/WAODnjKNYabVFHkCdjWJn7Z1BhFxnyM44DBvn
MpxqKuUPZE/BZqIvXsbuVH+JaNww+9uq/XtYJULKUZDdto7MsfdPBRrdnTz9Q8+l
onSC/F69gRkFsEJalJ0tHwfFpzSQhLsYugFbuUsEsqEGuOMUw469ag+vr5x3Daca
f6HOVEgZ+Jgf6lGAJMheNZ0ER+Z1JQyXITXsYz54tm336NNR901R8KAqXRKJXLUz
FA3MTMhxTZcRp1snIIAYun2Rb+5YjBz3mnaNuHzpv4RPaQp6TqihAiSLtXlWvi+0
t9bKcMDvs8l4CRXaRLCaBpAmLdYt8fSZlV26K0y5B9ct1lDkON2W9/2LhhAo1yyu
RCreqw16Kqs7MGHd81rVV8GP83soYXlfWVGBg/bQpJ1Qvpst3rbHVMX8gb73CXQW
jZtUqC3bYIP5C3AqCarHW3m+aZiCGQGix6ThvrYtJsoSrzbn/tkzsipZGtwFRxIG
ZgnwQT/aXuv5FOrJJAjLkpkBCjb+jEG0nMIIHT0ZJSvHR/V056o1yll+la9PzUhq
J9U4ZzuB6pXVZJ+LIRE7atZD+kKdFL7Mo/G0OFAHyqkuzhuMaBdcVJR/Luv4135T
0ujbHNCrqlVdgqXa1GnNFH9ZCfiePj3/S1CzFtxcAfEu1Hsfcu7tBd00A+HDM7Pq
oO49NdCuroX8jwvGbKjdnR9C6Mh68EXWNKNkyXmQZ/1kiNE0tM1D9Z/0tzBkUlpu
zuJfcPXUw0oZb+Ma6RekiSLVaHGhpcHT6WJsMOVlSKj5vhZRxBb8PL2rfTBfWea8
DIWbnO+INR//iipqTbqC/cesS+CeTdNMiZ3MqEUFq80AlVx6eQ9eNbPLYMcJ1dSS
duJdTzOZ5lCALiUFpzwafORFcNB12Y0mNtnMIjDEBTdtI/j1Si/PbgiDH9aT/Hru
PQQsTy+Y30ao+8U/19qL/+LhfAY28fJMHUvmm2N60pckXrfxxRhCjMwaw7r3dijq
Xis/3k8fxMCB+DfH8L2LkHTSP3cwzdm+d06X3twiZVy/HVULXi8Ybtl8Lvn/JAsp
lqgZumZYQsqgfszPtrij+h+U6NjJjglembs2coHGKIVD5EzoDCFhEOg/QtrFzMsu
dBIqUVzkm75K9xpqBHa2h7tjpbzRrJjNNRAHW5QpZqDgxJB5mZQcQn7Rrnqw5zRF
0P48p8AKfKgVgCoKtDRrjSm05+7RldBZ2nrdfLEyxXb3vrkFjIxvtVbz8mOxOs2b
j3kvBTNw6eDs+NQ90lWUaqU8fUZbKXBdGp2DBNueG/HmckAKXjxP/l06dRQ+qMoB
grA8dRtCz8bw52Wa5kG6SOcOyb022far3L0M1Lnkn9U/c7AOHh6E7+54pmKJWsjP
jta0CGshJ+v1vTuvymDR5FAU2xT+hMBEhmNNL0hufW+sy453D8WDepbulN5ZnMmd
rOmmEDZ2C2qNHF8FTy14DJTn2yuuUHEAqOlMvJRWtNuoaQ7VgiTgwcdLzx4lqLn/
4faa17jWbv9/TSjasspd3bgsMAin7ZHk3qE4dPBFd6oc9Kfrx1j8CmgmKpfshWfA
KwVeC76zLDFZkznlswipWKQsRkWEpBTbugJM7noPwQUS0DkZNNz8BvpMnXV19keP
yXGI42CGBHRfSmYAUicM6lTZpLoAEYrKFqPrCyWRMBINKMCpS9JcjbUWsOhTkhPw
V55Kg3TyyNI9djhRtb77mPtxwrQEG6v0lu/K91SLC9XdjjCdISLM4CPd3I5ff09G
laQhdIibZmDYtxYuh9O1CdDx8J2a6650ZLYfq3vmhcR48iF20KKJe0LCwKRZDOmv
svqZv1+gPCUwyHALd3ORy1dkXopEWWEIbz2hzoXi6mB4aO8xmkKBCemMCXEGS4Yd
i2c5erw08/i6ZEdZS5Xe22GkrN/I6Aiyv1xu5K3v6QRBTfYFMIvib+yiMvGS8MEg
eLh4AcM4sxXzpuydoarHRl7g/CHv4iXJ3vHqCX/hPz/NZSpR+JZrKmNy58t8Raq+
ki5GH8K5ljrxAd8TFEzBht4L4ZDnX+FixZkJBUg1CSpho5bqtLLBwfUui+Ub3JfZ
OwM6vlso/Ot/WzR1svy7F4YgjOIlzLpLBehDAaoF0S2XZyH3tIKR940hytpxi/hY
gS5LFiZWLuiMClGlvippWV1NrQAuyRv9TgDd+K8RJExDNUwT9IVAQBt/MJbHhPa6
+oH+CsEv5U8Y6s/3bFoeKCC7+16bJaY18kCLaamyXzS0UKT0CGuTOhISEAUfMyF2
iSKV76oXeyDF5EU9WWT4kF9ttHp0ChEhnupIhek1ftIlJG290+E4iocjb2I9fw8I
HiATCB2vKEbDHjyzj9YqH7Mhkr36/Ff1zOtP/EfEBmZuPRCvK5ro7njJzo3sFMxY
PEP9hCr2Tuu9StaxbA46+J+9BaoLMjihVMoUcqLteQXTifmi3Jv3s82qshWbyvie
Q8QROTG0n7F6xPBk4Mjvot+jJmsMC1U8tWyG7O3mQPeWoHSANzARoqLnJ1OTpoZM
3DpJ3JWw+i2FAHeNRRgJH9WemvOOCyczJYaOl5pihjW6lKGJt2EeK1zlnfnD/gdb
oTLAPeG489JnjEqjGI9/iig6TRYHkoR+5M+c5M5b1i9viWdVxdbfN1+46l1T+rof
rY04126n/fLvw5xCFSvaDzzmZo+YFqCs8N+DLVJ2iQZyWDUcRgbc12ZzER6y5ahp
Ij0LbNlPb3ryRuEj1e9XnsqdRG4fgq0X2JZP5ds8WFcZhLfI9TDbHOAUA9bQ1ARJ
GCbVE5YfPeBT+EBSjUQ24NddwZGEg2Qe63tscRIXnRP0d+AvXHRsPBTmBjuWdCBz
p7QRLy/ZnTMylVTzpZWRhj+hBaNiIalZDIlZ2ELzzjFj4hHO+jZ7QGczeZeOMWu2
J+FC37F0aS9lo8cSaHJ4pbhx55YLgWCwQH+b5B9Ye9FItYghoeqTFQB0w9m0xmSV
r70qSnxSgbgkfVQuPJ0jpfsTcfp47IpsFGC/P7T4TenbiTw1SVNBTHWM4KDYmqZR
4ViQQ5B3gHsm1/RVcPcAjFpyXRyGbllgHHykxlgYpUUOKsROliWKDoOCy9u+G5wj
2RND1uVUup8IVjNW8Ao5Rj4x8E5J8Zau8bYaZcRxr5Vl3d/tpJOR69VwQYP9NqFn
zvUJ7rX6EVXhCoxFUYH4RXgU27pPXnIXLTOgqLxCPs7FTiHBHrml+8CS2be/sXAm
LOgLEyJTBt3oZO0IezsyEmvRc8fb/0KHlBeG5aqdgnG9ZkbVvbjioTqwkJyu9Qz5
Qz1eYW0yG5RuEK6GnfsEpvvpCOuBQ/EHvw0VFUb+GYQQY03KAqn+k4kCJcg7+K+w
T6EjTPL5IZK9qCDPD9ax66W3JswJpYWOT2d6DjxDxMuUkPWBN+ai+dC9qOdlxjJl
ysJ2zX2GOav1xgdeVKr7uFq16a1fgWm7J4x+W+loNpX6bGJT0VaWzeP8xmcc5mDf
eptRljiBo1HgV7BdkHCuwNa50AtzISMVI8ZsNo7WnGrcQEnHGFH9VF8ePf9HbnLR
9qSq8RMN8MI+TvSSGsVKRY6Mbp5Z3Hr8O/f8YtrEQMwwxU69yhtQlMCi1ArZkjEO
yCPo61C4lLOfsXOmy7YJVns0NIozRxuFbkyibc3911HCD5JEgRFbAhb7pWm2jlpV
r2EjLQUZqWgdW83WtrPX0PO9vQgj2Nuo+qoQ8UY7Y1yiz9F/VYLcCPelWqLu5rPK
xkWbJqo9p0mMAykuw8m3AiRfhCBR76MZh/RW/yqTWaA/aSSxa/vN3e3SsDfalI/a
Mp9qFKO9Vj+4SB00LIkGtk+mxdWjlF/CfR9c4IjCCI+eWghnFIlt8ihxetQSayak
gmLkBH9vHCvJZ43dVUd7p3UCdPEdxSbktl7Vn/KWzjpOUzI9urcY4o4AABrSi9wH
LkekmTey26aV8pGpALFqxWX8NkQr7XPw2BjPbcbRuGwet4y7D5eBeSwvoSqRBShE
yU5SEGRYE0xDipmakN+ALJMNzv5u63EH9sogPywE0Jr2Tx4PGIqqx3ZomuwuuHnB
idSgpm6mF9hfEocvX+eUEZyNZ3HsvFAqzKUVaOgqhRT+w6owyLj2V2flQcCqPyMc
XoP+KPxosIo4HNc8lTBVc0cB0MaEse70KubHrzTSz6offLVYn6zVmal5kZBCXXlM
g4xlnFPFyoPKRDpzcHXZ/MZPiTJF8bJY0XrRj9TuIMGWw5nt5oBzh4z0qtQ4fqc5
kNYy3+b3SIFoyXIlb+G7/RsTE5uIdlY4hqI6PlioABftoNg0Ez4GA1Ng3tCWcmEK
nWOQTFPY7NpyUPyMFNM0xCC9pjzKXkKROY2ZoPvOmd6KMiiVT0ZA0I9aL6vcNe/T
8du6G0Wa4P+md6qQiub9YEw5sU64n1U+mH77D3dMRPijGxQMclGTA/GhEjmdNJfT
2hAAu6pR7iGHZiHduKcvORS+7rFsLQ5BO+o5J7AFE2pFIKvDSs8C+r+kuXf5UsRK
IL92TzERzX1wkmQ0hQAswq5RkikoJBNmob0ht19spjSaDHgUZK/f6uaZQiDdlYp4
qgCFUfy5yF/V264N7gydpQVyymrs4w50PFjGlJmMy7WoOHvEc4KPW2jW5S3v8iWj
OuJIPPnkwmcYMNnnUEmSFuZb2c0kveaGh8xr7318cGzzn8AFDrCFCzVz2ZyEVTCN
RYxN8Nx7yaHlkjiaLU6g/JKFZW51U2aqCh6NrPQHvyxl8fL1yGg8WUzuBX1mINr0
D0eTK6sg5gqqfBMz+nfXN3cldRj80jWVlLnobxBC/enBNCSbAWGw3leA0J/6Btsq
afPEWmgDHXApUyJadreRks6WZnePaxisc9Ys10E+8UdmiUY6mlOO0aYsGJPw0+e0
wsWW8C8n63n8wMjUeyeJ3IsUaUiQR8fCISf2DZfYS6D4+Sf9Etl05SX3HgRsdRXc
X6RJGs2CKGRpLugJyTbpnzcI+hTsYycxXzzSgWHvEjdKjwRbBVL/LzLVCXJgZIAm
QdXZkQJ2mISLLJ98P5ANz4WINrxWZJWkadvjRZLBHSXSZJkmhk86zfh73LJKHTPm
Ya0z9jF4unssW0k35Lfb+D74n8Ra8dMHkEsISoArVDYA1EGYHaspL9svrr9Vlinn
PKKlveOw+iMpVznwZ7sfTy7TAvZaHYW07Pg/Q+IMUbJlMMnxfpAzJGSGX3WMefwR
m+BlgmiJHwTD3je8McH4sGRx4/DtQx091sqjKdXjCTpl49VSAvPlPeJ7YDZeRWTx
18EKixjaI7DDcyEd858hqUHh4zgCi8X20Kz+9oboSzG6lyw+Ze2Z6Co5+4AuLSEx
hirpYyXtTABTSPZeA/t4SvlZVYNhNHXv6wCTNyfgPJ4CgdK8JFZGiI3q2uMW9pdJ
1/XHx1ArKfK9mZgb/AeB7mHbnAl4EzufzxVK5qiIFgeNsIqXtO7y/KF2NuqgSl+i
bVA+hPz1awsWm04Vyifo/8O8Z5HN4BhMRf5tq/2O70a2AXaJOwwdvrQTZb0wUMdB
d6LA40nOnY4BC/LbMAuFW2fYBXZqWuV95bat7IGd6viYATxdbbLtGtnmw8L4lwZT
o+AkeZAg9pRF0EGE7u4ekdnj0Oyeqmg+SZlRXL3Z5zlWDpRneRvSJ79hzmlBHl/9
SC8xjO8g4BKpUNVsMopA4jRFXuIEx0hHMalVFmoiMcOWh3ZuwSDE7ZqzrOcf7VHv
A/BHchSCF0RXOGlnDWo2Pummgee1mHk75MGFOVvHcG97PIeaSSJ7+ScfzI2zNgLi
5dSWk8mkJ/ygyUr+A22jNSKh8z9AycaKoLY3ZsG5UnwGGgKTXjDZdFHT3V+1d0nk
9FC7yIGZmvugbamsrNy7O+gyX6Ceund0i/QmcPofp/bh17aI8e6cCIBa4aj8J0qT
Hw9p2C4Menq4VY0JFnlq5j5QND7SHM3sqDKDIRfaRxAfHHqCLE0t6WCL1A09VfYf
OqNrJnIST2d+KNlqxl6j0tYQ6w2VtLP8z1r7PFzkx9lW0LteqXIBc2wwYiU5jB3P
KVyzOwJ5zA23Qet+aoS3LJjD3UsKp46NqLHsf3CNeNdEEcNLWIaW1qQxsXA+eCN7
EpEBpHldGFKWQRv3j/0Hqa1BM0i3D8IbRuOf4yygRp/iQisxUVd/QZUmVkBP/19H
sBq1FbtlN7RRTktOxiviLARjEjHMDAiaqJ6k3qoYfl+XqcIosqZ09yuWMRpTL8rm
WSb4H085AhtB3xqIlL1FqC/E70zDsGDH6PGe/hUuZ+faTqcy6owaPkG6iox6scmG
pGtBjVzNL/M5nYcTdoHRcb5Y2arkrHKfZ3FX0RtwxhvDdH5frF8Q78bC3SKPobzh
qn1LnOztwkhT8sSNFV8z1+Ry2rlV4CiIM3ubEx9eaDEr0ndCe8d7djvmf7H/eSrE
9kMVS5ldfarW+67r1bybXip5crvzeDzU+ErJTQM9G11w9pdEoYmivBoeXLLfA0P9
lD+lL7EjyrNxUSNYD/nBMOs81/YFbSRc6s87V7PGlMkTdgc1EK9PdItmOd+DnWbH
lCjCD+7YVEqdHbCQSZRY5J4N2JKwvV0dRFtJzSbluBxRRYr6NlUaBOfGrfr6WVO7
xGZoZxdD8Jiwg2WuiN8hKshFJY0yVu2LFhkfqir/BxJ0qlV/DpoIFmetkdlkWV+a
a3aCGsO50frpKG1wrnyuyTWZ2QPgU702wC+VEbbW948Ib+258MVTDLxKL7tUVX+j
srMmuS+D8jKs/zCZRDQ77L5UFzYSCuQFyHAcpRzf12gLEJKoHl/22+kDbpK9noAb
SG5G/+URka7uNPQFQV15WyLk4qsVxzq9RgSCSrIqoqetBoN2SJdsmgPXDR+M63Mo
8/rvqE4h1+J2C2LMryeOv8aQQCsj40GYs37MrZ/twSLAkdthrRGI6r8szBpwYHU9
EmC+ColeQ/7M3QlPAJxV6sI2s7oE+DAJj0VcWzWx4SGdcLyT3MIxDDPaUZaIMNNt
Po0lf7qIJzS8u02efhqPBiUYAftI95ry0qQLxIPZEeNVSti0BshNplX+ysl7ODJi
OCDMPuKhwT0/tZFXYrhaZaG2kEveYgphOV/D8ZCsxygV2826Duu7R3aZwXR4G59r
g5tVlyCdYCiEmEvicx9r6AxJcXoHrBZM94ggXGckEV5C0BhHYB68plcOkwR+kGWF
WPn9/FHP74fMSXv/7iPAys8JyDS9OubCBxRielQ8zq1LG+R9voDxT7IU0Km83BA0
blEJis5Bpnuvra0tMlx9Ctsc8jvIVRrpuj8sieLNzXEx89RL2NFP67f/bigJFI/j
OR6suEkWtfT1y7waf56XwurJh4/r2kOQvYbVG90zVAYLGQysC3uklA6Hl5Veuotu
Y9VpvUmZz3XYxgIcbeOw8LZIP96eQsGlqQb0teDBuYjfjoEgwuoFZl9sZ26+bpAO
TBxvaGQLcwELGabtCjnDmQPDxoES8B8xpaaSh1koEwH1IYzDN9V2LdXx1kfw8SbS
pZJNuSC5xQeV96MFM3yt1LaJPBW70ednRSdLoBqlxHvpgwHPQj+rwJKIowtsHqbs
Ivz9zohzkCbtyTwtb2A4tL864Fvd/HSP+nx02BdPyEJ/wyg4gKuby8I1q5b6+Bv9
fHpz4eGlBGnBjCujy66FOTV4+SJB8MVx5hl/gW5bNcZXIJA6RZJbGaynm5bH/pIp
1DHpJKqPUevaGj9Pj4aS2dagTdjl0nRk07UqakdoVbq4ot0KcOTsKtubT5or4jI6
8FI6tGukEKMTV5yWTPw3aOJ/tfkeLyXCSrIW3gdBe37Lua2ma7aT6UQicu7fI7VB
pRCNFLrymN9SiOIB+ZQvsNMuMtaIJlWDQVp2psujUGOmMS/qpWpMc1r0TvVagU2m
lPxiSNjLQwnh+Bu19fxaeQ8hPlyBvhlHl2dL99baAnpABW4WSKu29CAxU7NDTRIL
EYcLXZvE3WmS0UxsmcLz6pIbpBjSrwLZMBPBgGxIbX7X7rdG3M7oILhwZwSqEgSS
IrTABlKTBptc6Kdkol0z66xKY2RyFf8uaaVDTa+qcHwpHh6t/9vBg8raL6NOcWFY
Ox3k5MjyM6PDlHe2CzObxUV5rFCo2k7oyPAb0E+sqYOeXDZyZyqtvhI0vZQXElnz
AG0g5UMsSjSjlvSzciGnJ3MkGW7h609YgldKz83mtw7osCUrRz2hHYcXSmBLtwuB
7rL7vTsltxKVSj8Ev+zou61AkGNZ2rQt4xr/7GTXp9/e/UsPFyuc3bEmkFRjxv9W
1dEj1sSHTS/aqHAsMBK8nntyED4ivyMX1rOhzBx2lV4emwFYAm4B0+yLTiRDbAu9
Lt621s3OS1e3oOXMlzy0A4NkZrfSCkyMD2wvZ4kjO+f8PaLBYf70S8gJaxUU7ioJ
TKPaac0YIDLTA+cTqfJBvIvQNotLsx2yc8Vor9n+jHob7lrSFfbP+4I+6we5GGYo
mHsqcTK7xin9Bpf4Ws9okJ6EQJ4eX3O/4bEkUSKJklE8gOjbg3Rh2/Jkv2NN1ViZ
SG+/9z+YGqkvVVNEjh+SVpYuHTWi2ND/V7+4CQjHJWbZNA+xjpDFPMel+FF2qyi2
4KQB7X+z9523M5Gh+Ez7d8DkPbJ2BGIQxyRfg/RYQLmCF4JKWVB3b1lp9L1OLXfo
Vik9n4GUvl0ftexG49tYOgb3o6hDkjaogOWumHpz2Zl1f3tRtioH5Ltrve34Gp+Q
6QWzD9r6v0H9J2b56cF1fR5zfV/oopQCiwhuAj5B7TB8uBwLdTwMr4KBa947q6OG
U9RzDmGtmxeRQ6NetgZlDHZbCe3k7xG1btDQO4MArNcSYRhS1fRC26CiogHg1wFk
srFefoaYa8UGBuf0FWrWMWYtI03K/yYLQICTRKJPK6EnaDsxK9ftUan73G99ufaD
uxnGLPedi3oybPrubHK0LTtN1aSuSwG7tC+IBUTUAQTVoVEwDUIojRdKXZ962Qki
xdL9CeHWlUa7QL5/w5bKLsxzYUYw3foCVC2G4JDVI1D3Q1tfsfajRWZCHQ613BGJ
uzyMv1MP7mXAUGiSXem2s69VK7Q/TdFpjJiAvsb+wd2/dEkCTZ9IKrXAyzuasFLg
HFsPQ3vrGEaKcw99OfluD8RpTpuBNRSUe/AlRR/Y2y5NTW00q4E94/jF/LiMDEuA
JxcfVxEvEJ3kJ/yNG0cHUvnL7dGUrj94FIMhr/9m8kbV7vnGXtcGAvJTOd43Algi
C3QvR5iCyB84ixyV5kDYmpVG6ejkjSs+HBjzdDqflyVgs+GCJh+1P8TF2CfdakZZ
TQG87VZt10IFAggowDlK17czwwWUBjoLeErsQQzZAWzEvnp9l90Mlmh3WpH+CgRp
ZUrCl8MMwlYQaYFyUhluaQ4lA2LRkyGJ9GSo8kqluotHBfPwWR9qJAlfQIsb8a7a
EkIkTxZEoOW8YTBCttGINsJN3hbVVVh6TKkow34RgweYvyKrTOb1NB5Me/4Qio6/
vP6OT8HkyF0hrYvbebEmHDkKc1tvZMR6jADSXP9y+RqgP8CJhK0rHeik/7fwRe/E
3YwC+JVJY7ljcgWw54fGmfuNI+9A3iuBo/ArJXBBucfiHouif6ossUg49m8wG3VJ
Hno9ij4fcXRHhdMwibWUM7odAvu2rjqbddwpPk3gquZD2qeVG7bBQjTqt+K+ecr1
dVX1enSyCvTYeKp8Vzfm15PWjAIhyrRG67+0xecWFefH6obRp2hHOUCKrOCp2hOc
l0Jvxtfh2Q0mEV7HCKBLQK1hi/hQoYxXx4GAepNL3H7KiwGUXXI/cP3clXmCtCkI
xYj0nUQGokpKnaQEHTD/mdpIX79jwlWCcVVfcLO2CYtz7J9+h2NDLbhlc6mUT4m2
XEfDqhwhbJzwo0xZjK4QQye/DAjzNfGFKIMcpo4PCD1XRiUnkPB2WZ9jbdPuQuAg
Gme+KJAD8kMR/VRcmVPE/rmII47xjBEsOEby5qQYiKn+zh00TpyLPzsxwOiMlLfO
uTQqcQh8nbiSSBluJ3M2l6Lw22B/9Tuw440J5qNDJBy7wGSCAfnFC98afRyp2EJg
9tdMSDJOWsvg7Sn6bAWEsD5hm1IocHrfnTvZ5L3oDkmCa7IXOv0G2bDjEMizpHLZ
7jlKWweCvtI7C9aA5ME50kj2CZU/cyVsTdZ0hlq+Huuadt5ku9QfkS4mOp1eQ9nV
D0z6H3wwlyhBn173VCpowEjwN/ICDhH3tpdaniPZhoggEScjyNK8hj/VYjFOdtij
CwIARxmUrm8j7iUhnYz0l+5O82i7jptHhSxbi2D6VSstTfTKzbWgJ7WtYlnLPlUn
+CqpgHF1cel0bO+9vgPMB+prVXRi+z1VUuf4IFpPFcNHCUdjfEIb+STQQBxwb2jE
4Sq+PCJ+ji1o41bX36iYxaFzFH36HNp62aMnA0Kkihorj94JUVHbFswNkdn+9wuy
Aew8v01lIWmjwa2+Aa7dPdbjIpLgHvpC3Oy4tglCtQB10PxZJAvJx6XF2krFWLd0
Xp8BNc3HZyGsvPKmMB1FwMiJFlrhr0IGxsfi2LaP+SZssiAELCiPqOeUxKSErs5x
Uu8uSZnmPOnWnx7WMIvo/srI5MRSHR/RuWaHwBArx6Y5umscYhcL5css7+dDcVhS
bwqdyQUSnD6pPMNlCdRlVWH71YGbrKP9kF4Ui51cIp3q3D1kcB/Lp6K4abLsTrK4
De/H5WStBJKtlynNXg+ZOR5ggmo7BeKIltWuXigMCQj6c4wDm/9D6oZiGAUPx2Yj
7K4x5IqwoZJex9PbDKsWB1SHYt8H/ww8ngShWpEZuEMvM2+HrfpGFve9sEjaxsUb
s23Q3k7DObWHfJXAktie7yT9s+av5MEq1JvRpkCfMZSI3bQu4i418GwnEvszejm3
mtZ+PEc3k50twpWw6B8s9YVf8nFToP4wFln/eZbCHkMkWrnHpz1GWlr7JHaBkJEA
VhmUp3bD9KUhpIEVwCjbvYbVKwxTSkx61LSKGiWwaPNqCiOOwnfwRXc7pl/Dq/Pa
Wp84wCA81qPjnWRA71K3tEhD+SnJOGzda5AWlVCPCKsvSDpOWYGwite0685milhf
qnCHwXrUMj6gAff8Y2y6U2AoFIsJaTjUJZloxGKajfh3aElfaFgM27/U1uczZotF
5U4BihXIh0liAUKAe1ZvMUPhPYZGCx4ohfzmow8N36GBZ/BzK2Fx9RjUqF4P02k7
WkvxuYxaHghJ0ccS2Zbu39AwYazYwm/UbQF4rXtuwmrRkB2eiSufURjTOZoLxPZe
CzWLsF4AqSOkpD6nYrfbULrxJLCTQQ3BiwuyH43AcYUPv3ZOEhjFiicg5c/sTBXj
7Tc3Kr4qFrD7APEzM8F0LL1SLjvKPchtKCJbvqc736Y=
`protect end_protected