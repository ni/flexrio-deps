`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15664 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10FbFDoYe9P0I/fePN4jRvNwCFWBa2odqRIPouNJODFqa
MtAuiR6BISUevSNVuTT3xIGarRQfTFO+d7nSFxQEq9pqFZMsJAVdy+b2Q0MjIOJs
BCiMWHAd5Qf6xK/epBWtFtlSoCofEY9p4qRWtJBPKljvdvxgmJezXRHaBV+i2CVQ
j8RsHlL/ZKDwnq6RB31MSsiGeKa3nZHCPS6KYd33cNqUmvRx0bXu2LEfuYoYver3
DTZIz0+mx4Ds4KCAxGF3UGnpxkmM1x3U4jeyHhbfrAzpZEcphKYsCc7f3/M2o7el
Nzr105mpQYhnzF/8syak0CYfdakzNnEd5V5Imp74zH1weXY5sKLJKPUMNLR7A2qo
5OsDpHlJ327c876Tzm4HTZsxrML75UBTcJk3R0Z+f8hERcWsNeEDBWPkkBi7C1DB
EN5YcCdlTaqqsqkPY7KLMnqHmZkALw0ci3heHjLnGQCg30hwZeIzTYCisIGDUfST
zw/M/lIul1KkzgnPjbplXy2hq3QrWMP8prOsisjBUQgI3Z4x+B7NBp5zEMWDpWwA
i+Wuy+duS62cAFSwwakrSBOzfQXedPjlPH2W6i/4461c5cNf2lpaCuweEnG1LUh1
buYdZZfKOaA/orKlw90HnV0xEymVg/iKaJ/FwG3El5lYmqMpTCIv4nYB84TrT8dm
k62g84h9RxYzo0huuwS14qA97IyxjKVOMFjoraHmPQFQv8C4r5Nm4T+9fiNbt3vO
zfWWvEn12WQNAkXOj//yPS3czgqHE0BSXilm0U/IJlh8NqpkuU2UujyUHDA3+tx7
9Dxbd2G3GXkxVcPgLpRh8TcpGtXkiwdLKQ8b4AkqMSsv4OAQVkU2gj8rR1tzT0ac
pY5tdsJL9qBGa0qG/ApygFV367WR/M0lnUvxWGX74Iz8bbzigul4CH8ZoMnkwK7J
zQIKNEW9qEeBRhpGZhoc7UEeI9iQKaes3y5ehdli3etmdHAd8JNJReErzhlGSfUU
4pOL4EZpn7A2QJOrCPvaJMP/8fU0qjCFzESHxCxYwfTd/ECtVVqLl7q/NpSnq+n7
uF4xpBKGC/GoB9qw5A/1EQJSJT6KdL8eQepZz3dleWY82zW8UDslcax9YeB161dk
R7jW/dIY9SsoXxhAmqMASmVT+uKU8b9WjG+DdtHGufFGMeZHE22hdwAcsQwf5CVS
fxoUiNsJu5e68X/vjlweuaBYtl50KCrZPzs6aik/kbJImusCeA0X6/03VC3s2oAf
qvkq89P5YNKy6dJeYWxCBY//O9CU444g086D2yRGs05VI4YfzI4Xc9dMHa5lnjBg
1Bgcph4EuA1NUpOga/EScMZLgaTRQAjac2v9EiPHSk01U1zk5YCPtj0J9kTtDGjv
S2rTBKwD+1lPvY7JJb+Pu6OCLy8zgIn8hZeqdN2EC46dWYJuF5959hZoT2NHFj5D
3s7rvjISALiq9jG1rvPXyHadgk+Qx9Rmiz6ikUNBYoZC+W8rGokVhUskR06siwHH
QjisqV2BKGqXdfK/ireFOLgqQPbbR3cF4cvTNK6jwf9aDatRa9+S15bt50Dr9M1e
OsFkVmRg8GB/OrWfcR/EvHdTWq3GL+0tBGEsOvYgPZG9uyRAltv8wxOynhD6IvhH
e852KxCxyFkx9fXvVL1T8bmAU6GwmNaxbGLHb/pntQQogUfmUBDT5yvoafBDzsBg
MODqkF58wBLA8PEix5JuQ2itn/QaQuYK4KdjwX/JGN+m39Riu0mTQnPtje5dqiZo
NBioo8Yj8uGCexLuw9UorwiEz9ysP1THVG6OQvSZjwStzHTgK58FARimP3dU2uk8
zGJwpNivaUSC29yOfH7AyrebANvG7HuCMOBopt6ysluLNz7yoEsba5snqjzfXLIB
YlSVbwxlsq935dH2vxLUMhrqMJs37dFKIPdhw+ZqYYuc+aUl78o/2oTsjNHX9ZD0
m5kw2OpK0/veKYLRMRbqUeM2cKuwjlnX/T5+bkhrJX14VLN+WdEU9b0JZA8Rgpo7
WWpjnuPJB2TeBTmXKqyjxrVpnMy7DtBqVjRhiz5xjeQ+Nhmo6wiKs0BMS2cTcYOY
chZ4U7B9G6ROVhiZuISP08ky3Rmj2Q5qTMDca2w3YtRODFn4zrsdv3Wub87I0MSn
l1KnuJKqh+2/PcEhIR3pHFOdxxxW4X0DDnYimvZYLCyHtLhY01pBSMWqda6vpEiM
1MJrSCFbMJp0FIG4aaR0V8xIJNqREgNr5ch1WY7/tgBAdI4dtRGuJ280cloDlS87
BOCnjTm0hIIzUS/rx+EoPbhGYNcWf8XxkUJnWPFHcHW+8g11WvRcvpos/ZPpuGaj
9TqDazqO1cydJGrObrEX9Q4bdoQhlweW+7Vgr5P+Ob/lqy5HxgEu2jIj1VsT8nA7
4vAQtVl7Fa1iKkUG1DQBEkqbny996kAmf6dS68nHsstSZJh8QJagj76sE3Db6LuI
1ajen6mDbqo8dhrVtJsgXvj6RobonabX6spH1HNwbdF4KG+J1VbC7DiVFRXZA41f
8HeH1yjShrLTHAX1kDz5Aa1mUA+lGyMP3w1VL16e+kOVIO/bkkIhY396eR8+ihRU
kxk3Xh9es5i25FEI1tGV0+FyBDUhu3ap1TSNdS5X8UsGvShIxdi3hiyU07sHr+TO
hUC03ZPZTbckqIYHB64HADRtuHzb7mDR5+6LNjNwRGLVs+lEYahE/KgeXN4TuEMh
Ioh3uH4vwIWbpT57LM2bNx+SSMCZ4qNts3P3zzFtsPfHSp65KIDdb0OOeEwVejuY
6jxCbpP1YT+K44rS2jdyNLrJz5o4/b7tBLqjd5gVzQriA4va9HZ4vwvajTjZeZJJ
7j7e7LR6uByVT8JGff2uxMMbN6cDYyAZiuq9A/PPfjNLaOSeo0NRq9NvSgd9YZKj
cpLmkdS3AW4UgY9oYjjq9S7zeh0oBh5m5G6QBjGKqt2/8CRtW2zD1SeaUnaKdVvp
zs/Xlt9F/48fR4cTpTje2DgpCW8VjAQd0K8tjrqu2OAi/ohvJPi5aXxG0achIeYt
G7iMJkv4A8f9SS7ywL7UowETsFHQV8yVd/4SYZuqE/IS+p51rha0yy7bKu/Bkics
yYCxGGng+dZzqm08hJlgbvFODmT/qlg9i3UBq9JXT4vD6zeWvx3tkHSWCHa6U5Fj
bZAdR8m6/9epOHAQV47Drx4/o+kljGDbWPJtzQI7DtuFr2C/21CMlQGa+Bi+XCs5
FKxZR7odgSOT3QTrf6JmSZobW22gOhxuefNPriSuBwHFwJjZmJ8mI7pe6edD2eN1
LljI3Nno9zfBwCnnlIEEfSzvt+k6wJAPhIy33z41FXV9M/E2BQjaTAFoiM3p+ZJr
Tgyu8uZjbG8VUwW3tB0Ku+uNQzHxYOxsdlK2ISpl3A+p9BvEAEsztdz3oOmzdvGM
FZuWGVMgFth8QS/6asOJU5CbxkbppPmm0YtBgpbqx7BQ7e6Kf+by6iUY2y9HMs5r
FdYF3OWbNBeDLMfPcoPfiVyTvutJlVPJJUKRZHEFRha8aeUVgeDjkSGvVlPqGrnT
gVmNsprr/QRCxRjli/G2rC43aHGyktJNpodXIJQazmBCzFx9gyL0rzWbg9D8tNna
CiqCF/uvSKuuOAsxEJTHSUNb3EvtWHtxml2JtoAS1qbV7NqrFF/kOgNn2vyaw+/+
V28Yq9tum455vAp6gt79OC7uIO8kdYnSbaPwKmw9reI7bJuM0/aVDomBrJAOpL2e
Ei4DEJPzNvta3J3ri3FNmNk4ENRWYSpuQ9oSKGyCxPdKDZlLaChaG9LDV8R1dgrQ
Q2mBMZQaYy5w8U+gNgOjdJ6uen3qOs3I0aIwnqwJM67Ca3204ySdyrwqysDE9PpG
SpXKygzzPEEog2q9bqo+i7cWvPMyWG4O15qjb3DSLc4zszHTfIxOhMyLmVXwkJoi
0vktEDriHL5KloRJ0vq/wjcBO9PW98eGFmaZDhspWORbYGXGdxjfE38F5l5Q1MW+
Oz6DHthSVa4Q/CLlgfzu6rFVp/gsfmgFn6G40riUclw26FwQmoecwDzZFolWM8Y0
2ggAZUS2bLjB+cryxfCTIgoMtNjWcSw00mn1NoYiIL7R5xvsSrBPyZ3PTBR6DWVl
GD0wF82WAd8R+snvJtLawEd39T6eYP2pDhqbzUUWHVS1/nfnjQk0vl2FzG8XVb02
H7Zsi6CC0z+e3+h1dG8WzEy92/boikCiay0PIKl+GsbGrsxTdIOKfxcFNJJYQZg4
ckYt8OgZ4KqV98NBCbquN4MIUYXI50Uj1z2lrYW246EdplfBDWm/dqr8Q9hO3yUb
FlAGK1YlkIX7Uz5txjdAdgbDaxDiOlmgJy5OipCQjJy3vy3r3+wkKiGfBDf43HPB
31msGBS81NvNe//Z7VEVwHhseurL7GfsyYsdaj5CbtJaB1zqmQp3iY5yUWSVub6A
tNwyWirzFWzzgaP02Z9W923xsad7v0vBlRekPrs0Lt8YdaQdZo/TyFLwrJUWlywz
Ta51yy8WLbBrYjm/ZGMyGh1I1iHzFldoxkFhmChv3Mi8bnKDKoVzp37N2P0tpEfP
ZmZ0cKZTWFOZwmbGXknFodhyuVZAasz6T+J/ZVwDgBlwowe30YfdBVhTsnIwTRbh
OmcqRHB9BQQyX6y34SuQlKMwu9fpSIjtuX1ZXlNKgX5ECikHCUdTaTY6ME7g4ZB/
KSjJP+f3t3Xp1Kvvmfh1ZfjZsf9ojXZ41ee/efaeS6Q4r5iacq24H8TXERuTSlXR
w9OMmh56u9tisBtAtJ8lRrwJvCUH+Zbrcad+vQoCLyYXmXao/u4GfIyqatkxb6h1
k7lxRhNOsbLDomTAQ/FH6AWWX+Cw8Tw64+MEBimR/A6mZW6PD0GgGXr23WsO2qK1
yROaXfJt1YHBSUql/DE+YbOebidQNwisel/rSEZOxMpgVayCUhBB8KRKXHhB8FWM
MnTrepblhP/F+G+lVikJ4loWj6zXHPHm0sSojjWlSWV2BMHlp5bI0lc0I0lplO9Z
LHI4w/lkOv1QotvIg5tLk3B3cxSKIe9Ae7k74hujxTY/KZCvYaVImQuJw5L6cDhe
Y+ZNqz57VpDP+wy0/J0/5fitJkcltAIVXI4lOKnjONiz7LJsuFCiXV9nq2E31vqY
OoAESyLNMTPMeCh+00EORftHHkzBAAtltMF6CWtnMMvgF4RXqW3jNz5h+MrrPxzI
WxrL2XJYR+jjoFtgW6kwSQ60V9kdRHLIUd4zJiDLr2Eh1W/b13/KC+4laWMWAuvw
wYqZ9HCvH4Q8OSvl8bO/+S0iOlG/GcRZ7dWOOC5wlNPIubb5l9oPXHHFurYMRdhS
QObPnAAsoMU2rdzS9jdZ7uRxew0dZkO4qO/mLU0ItaQaT/q3NCBbmeyZPivzhG3W
DdYARnSSeCPB6nYRJjaCDmyyD+xwXTzx6AwcjT9UGO7cfPhT75jb5vxgIcJV7YAX
kJnofqL9O0KFLye6ZHMZPwLli5adPQDNFG9gZGxVbWNaZ3fU4RxyC5nES1nKezXG
2u0p7XFOr6jFc8kdPhTW/cE1IOMWV4T4Sm8eYgf0tOme/zU5vmfwfSIy6PqNjbv8
QEu7phFp9JuB0yJE7WZJcm5tTUyea08WtqyHOCscrQ2vZjFGlFudBUHIfsyU0KBt
9pbtKTPzQcDjqcFhTP8wvp1TgRh1hM+AjDnwGvrBf6m+1VvgrBG+bAmNdn4hmu1U
/Phj1IvCc2pEK3+uBAERHWm+/cPi5jzD8j1FCu3X8skc2pvWG4+33IXWMoiSdZFL
CpG2QmP4F7sePUfMoymvd56tHjFGGzPRnZWKH5V91GLGXq2pe5KL4XibL1ELFJsX
PVxsigVXFdnXiTTifycQUBnJqj09klNyd8aEWj6dJuib6mUDRw2q/f0Tq68wHoUL
TpBdSYrQEMyxyV0RLvfEUINRhC9tLo89vb5ZQ3LUKv1rm2AZXkQRlCwbntWkHJK9
og9teGYviCedfkY+P7cTdBbwl3qOS/rsrkyABfsYAQ7/INf81+sW3GfqSZFRIOSW
szM72VUj/g5i6uaJBfiVLE4CJ2Q++6K8Ub40G/WzjUlQnGUTk2pDR+BF9hLFTOX6
EflN9HS1jFnfygB6MWb4uXbDBzkzcqkTQWvL9KaIJ2wC85aYdu22qbdpuFZuBdzz
FH64VkixKpURFc3qBkGzJXZJ5eXFt369adJD396o5er8g+st8Xhj6kvyRRuZrlqB
kKX4vATlTEEflE40GuCmvhkKDvgzYhM0Ejl/Rqq5G0d9GGFOliBrt8thfkkyyYee
gtl8nfxGlJiFcszSGg7Uh2FNi43MRdVhij/CMWKOi5z8SYkxuOwyu+ifidjevWQ+
2UTggWfj5Ofa9QGKOpmNzAnBrMGaVc8H8GGZ9g4ZnU9veXG6WIINeBkCeUfANxLC
FREQyuHywZeVo3hwuBsCisYjgifHDMEoknx8wSsKbq5BGB8xHjNn7hV+UaW8oaek
ULna/8O9qlafIXcwjukBsoGLczNsota48ubAwaTr3/cMrLzpOsHtzSUnm33Gc14v
plFjBgTfpDzu18+9VjPL04d5kBDWPl8wIUCAZ4CO1SpTXal4hHtgB2ScWqK4DdVa
cfIDRnd6QJWqxQzg3QRgxt+HAqHO2mTMo9Gpgue3wiktnrF4YiLhAZr9UhnT63fl
Iatag1LguaEl4QBCip9jvRUjy3cHv6gJaYDf+P4YqwLaLTqnJdm+9U56A2vhG65E
iStDw2wJit5R7Y8lew+TtiWoeZmPFuuBMckoTTvhYsHSAGuKFxZkDBiD+wY00/HE
mHcQdkzNwf4ZnVbMG6ztdXkc7nZy8YJq1x5o5z87ddrKvNiWwKvco2L+okX0XqEW
jxt1Z3QDNDNZ/qQf3Fo7k7CN21nw10jy3VHP+dkASvsXAPc4vf26fwzSlI/YV9/1
99bLoM2po+cfOYyLAJgCoRUbkjeawXxqJ0UUOzXZgTQiIYN4Stev/cXATrxbvcUk
925qha3oTKXtvc+b33SH4cX0eKDCvr0V8kSjgNA5kt9b717sBHXXzXhj0oxLGCWn
59mxYftXwoPe0KsyPE/DW2gNt1NS7BnOQERyoyJnBOVco5/RQoQm+e8++3ruMSr8
QpM0oSYf4cW6e99Dmf3Nf/1HAJZgVa+bWQqtCTK8b+paaWmBUO9yuFTHpu80ptvg
g/0/RQjkI4WQjmgqDQSxzfclL66xF8YQTqcWg3+NlV8xHdwuFSHzYYfeGeFqYE/k
SuDqMfXiw2Jl8YKbu4U69+0VNJ5lwqhvKu84jVuqT7DKjvq/Nh0lJV1+r2e+3pfK
rzkG+UwD297miqAbg5U4WPVcLMIHRoOeONY75DCh3asSGQz1APToZsnrHU+rD90d
tpczoWulwT2UEO6bOcFtERudfhvmBrlyrB/EWj4sQ/JNMv10+LSmczkbXe6stszk
rCnjMXmnBn819oXxfhLxAxCHzg6HgePh35/vhg+RepOFpUd/AopC3PS037heYnfR
FBK3a2UWWD4Yyz7+kQTizQ90CwxLetbrjP07JPGU2IteInE41kgW+Mr+GGyCTiKD
MhwQv4ecLwuOdeuQ+dWb2op2RkyRhD//vpjJQ0DRwLkeQp7UAjNMrFbLWuzm7YE5
p93PREXGMlq/BT1C/fVkacOMikFe8IOIAaL5X/aaG2NV5c8g2pTLhidqLqBS/cxy
L//9jzgAdkvfGpIyBQIVblCZXjnwSsZq9tX/n3RTIXiUPeNOKMv88/E9x2IPOlIo
nwIwlKqICUQ2FwNHvJd9S/wZlzuhQpCBYhMCtQmXQjJJl1fIiZWGDcT39Wi6pFXY
W44sBFIuf+LwXW7js7Rpqu67NM4yp1+DzrloORX1jOLUXDUOSxOKan8V2NSFrH4c
mCMEFAm04lEZ/1TF/MBmygEbEUt4Mm6+TT7hSwHWd8EPyi6ILkJciNki4S09KRmM
2YjqKyW5yKDnczK5Qm4sz+BP/XjXdb0y/ne7uhXVSzqSzruQoNhapDYR20lTphPy
F5OF/qARynwMOcAGlWFCq+erIY5SFrfohmElDc/uHcTCeOwBZ2+8RPrZeGMYSD9y
bQsc35+dCECL0XjZdd4MTuXZno+qXmoUhMzelHFG3D0PPIGYJDTEDiWEZdl9B20L
T5xcmurGHqT5vrqP16VfTSF8KgQjKpMF7LBPO61xTDl56VqSjJ2jyXF79sNCkfKh
l2Nuk2BetSr7dBE5adlGWLi8gx/jphvt85EEz1b5W+QzMWc61pFxYsSlj6ZkEJqR
yzrxWqhS3U0UrAd4F1zHImlvE3m9up4c8OFcQ7pFxTUEaz/GOkMUV2I3DeLAQuog
mLoqThlkUlePlYAwnLiUCk6ImzEgCXVaQEIaltQEi1bAuG4iJ57jM54dkcX+QrAi
7FtaeFBoAJp/1D/y04Gke63gBqZvT5quSY8uIFggwzWzmVzH4OafUEQENtPCWRLg
V9VHciWDzdMUZYFKdomoVsrwUVuJUgX9C1EbDnPIVN9VCWWk2ZG6M2CVy3J7ufIM
K6KHyUrINMEwMtlIeWwBZl5hvWEx0gNABqmYooZxao8RLhz6lMVOVp6qm21XDYh8
5g2ubNDx1nJoMLvnM7yy/AiBC8kKiOiD2tRNbbTtcjnj1N+oeZ42axbLVDnRXn0Y
p/bSXMtIIGoXosdjhKyW/vsvwjBtlIXrLgz1Sgx8dOwlIin9naQSoeVW9LOGjYvK
yNs/K8her49miFOMjywOZCfZslUPPB5fKWot2AcnTJtAPjf6l8Qj+0XvTUJ0Srv7
CKEGd+/S9Y+ahgIodqumy3+jJlxQd2HV+zZr0WTM53mOyiFNRNCJ9kmJsVqGFGxF
7E7ay3+L+2R1Pz0hLuAgGsF9W5cGzu8TJwiz4gNXd7ndVf5z+9fGNL6qTL55jVZ6
hz148/F050+LaA30Ww3VLFCD0V99S9FX3WbDqbIlUtJGlKoKc0JXWNwLp1d2SpsD
hjs/kPnrMfdiOvuKGnRHpkZhI8LRoWMmLzXAniyJT/kn3GTZlMaJjO0Pr94QNaSq
BYMWnmEgJq1+UeexWrmhlbK198dXjyaorC47Ye/9ARoblbVirCExON6Bqm0AfmGE
r5FWj3aqvPoV8wNvFzNbtb8dSs7x6cmUNtZY+mwSV1EnYkJHI//xVYJewyqtgVmX
vBSEOi2hOSTr/kD4brGJTRi/qrzWoNUgvrZnpv7DWCWLJxutmQzK7JP+Tx3YO37o
iZiRa/VmItQm8DPZIb54C+gKsMC1+v7zh/uRzNVKUBaiQuxe6BH3dXXRQ7VFfWcK
QeTqzM9gi5ZN0WMnWT3DlgLtwKn0RNOvT0Q2WzN0yv+B7jN0nof8xCO8qANwKj2c
nNVjpFw4OofVuvId0amicTKY3E0kwkeX2UsxZXS+46MApi1aqGaJ1pUS85mY8IvS
MPNjfwlg6oqp1+8jaj55qN/QKgsCNA2QZ7SJ71LSFf2+GVCpinNKuBgTKCQ79JHP
PM4OfmuG9ZFCdNBk3rW/iWZVO1sOkx1thEpb87T6Qo1618aaMFwKPWO4nQKsIbjE
PIO0OqC+nk+OmnY9E2VulIRu7fydbaDDZu/EEGmbTKwkZmgVBxKDBtOteVK4wY+H
2eLnpryhRjKOmBbafkcOE0CKMcOts1VU7ogAG2qmdoR79NrZEVLFkSEN1YZajejt
VI8fzSN1mOPot43fmEtN57A9s/Fp/B8IedpRUSPbYbnhhbTQchKzEUK16AnG/Im9
/DhyBgVKtVIY+fbmzAktYXXLZbSyIHHfpc3siS4qn9A7cYnD+FZ01AwdgOwACeHO
atF3PtY0dErd5pohQVpDVKIm/tNGNBeGXGWLAH5/45e4THGS6wr3UJNZ0VUqfLNg
FMLakW5eZKz4ZzR1DYYbpeCKL+61e+NP8RaXhm7zmgRi/Nz2C0d6swkcSSdnr0ml
LSvg8YvVv0U0FbFp0F7UdNVecoaP3zjKJ9saUygn58g2uDSpuzghPWU/nwPrSmze
QHKKruOOAl39GcscuUivWoIikZD8xXnbiDMd5CTUzhsTCo/2c9xilcgdYqF05nou
W8vUpVPF9xI+7ZOKg1r6bgY/OofHMSzcSLi3b+guYhBOcX7+PDqElkOGH0u06nn1
slN0Zxvcoibp9b0VtbGhY/ox/ZgC0zXOY3FIlblEYprpEYRlT0VSsCzOEJrlNeQA
cd/bYjy4wJrsKSMUh129/1j/UOO5R1pIp5sb+QJie9+s4EFVqyElGbn1wKvn3rQM
twZANcUuLgLb3vykiDzMX5s0esiw9o+MrMxu798Vg3M9mgPCFFsf6QabrytYYgIy
5yA5e5GRp8/MokAYYeLj41IGlxudqtHeQN0BqVQkmvRAsLZiunk4IMzCfmi1RJER
4tQ4kxYLK7BiCERY3grEAubk81Cof2HFJ3coH5g89vyAeRTpJtf5kMO03dl5m1mE
jDENuJG7M9oWL1WCfF7A9cyjS5u27FO1G19SF+jFeLeUv2v44DGXZE9G4MtwoZXf
pGqpR05ClksjQVrizcUEilCIAm3XR9zGZsn2CMcr1LMsxtnakd+uXUE0LC4S4IDw
mFAJl+/0ogoNSmKdUmdP2uSl+zwUvpsafxL8d4KwJQ39hsTYQ58+ql5abjjeU4ln
6jBFCJUC7PAlPKm+TMFqHicqD1IYgIxPHfXX2RkFedA3rkjF2x77GSessxZ5ai3x
mJmNvVV/kMMxMRXGQAk4/R0SnoFnMrFzRhM05mhK4itV6zHd+1tK+SMXdXxY4ptU
26MoVNl+SgwqSloWLS4uBxUtMkwje/nV6XP08O4bdamlUDRrgi/uHJfFBRZQTzhP
W58SAq6j7iUF+qZw8EC5+JLqekOmW4Vy6iUlVbaZIGEnN3OR4OnkHJpNT1fFs4TG
zabKhcFn54U743eDuax0/leIp0FhPAMnza7iWJbyMjo3FnUIGdMve7+xG4zB1Hzm
YvxeIVW76DjCp2lMwE2KTf+FDcxmhRmglhTPZEYPFfMbbyu+hqhT4h9UbluFSnt+
diClapTvZkpH6mRkiv00Wn3yR+Dve/wBaqFT86OIzXQj+kFB8Q5mD6BWf5sqNX0c
6vVtpaSIx6BaL1Xe95mwJXnmcersgrbe/u+Wp25ffeYZ4bU3l64TxIvSK48N8Fej
aBZsB9CRJHxoF8/TKbkBzu5T6hJ3govx9AL5DzsUclTqV3Xt9t1et1xXuRi7dMWV
A7m31nMiQZ+GZrF63+vrbai5tGV0T2XcWlvv5zRfT0Uu3OBzesrK/4I2AZRJJLYu
JmVPsRbabk820jtD+SIEFWmnGqHDBp0ge8D+JLVhXtwV5oVxDMi+TwvwqDas+AiO
N9CxVmI8DFtcseLd/AeF6ybGhsfZeSkm/f9DruLRRFN6neJGI8PLt5xDm/aqDzjM
x4oZR5FC+rJ3HNtApfKpe2/gmmrL3I4L6xZG3PHBRmfbbL4pCj0FsH+uIx2XQG6Y
9tnBbuVwnpOuJxodNG4nOIyy3hv2MAY34NY7AD5i0xMUJGcD57dj63AFlxJYU+18
gvExqwCYJleASuWnq1bFOoMZEwsNjTbq/InMoXSteibV0QEczhGZ3dmBLZoyNew/
pfkxjmdKx3nMUDnLpyjvoJ7NW+DSp4J6pP/KgIE6pUnZ+HUtLYWpTX2orYRl6cad
7ZTjnurPU5Ox3aZYSIaJTBYjXmXjfs275dYc4Ywji809F6e6mZZkwBLM9+akSaNK
y8MHadOwu4nc1pbutu6sM9Cms/4xURW42QEnIYpKQBcKnT2hcaghU7E43QAlXI22
zrTjyvtPf7tvqczOaS9tBRqdBbUcyzOX7hvwDcIlGjQwz5Yo6SFU0dBDX/oz9uk0
6+AR9kJ+7GZnDJ9uYtHBOAqsvhuLV9V7H9HazEXhRx02g2NeTm+cnXE0z5pnoPm1
sm2VPhIpDCjUFivTymJa8omr3DyMTsvI4LVp9k1kpjUJImycAVOeYb6XYzU/k5zC
AhKBUoyTRNzM0zj/JaqNNOx1NkNSKKnwWGeXMIu7BfFvGXy3bIGvYqz7RT+4UQo2
h6SS9XJ1jx0fdl24FmCxdQEB9QpJypWaEEeFRrApqh5m9BAxEiC4/CVMRC3/bdIO
aa9PlcbCUtFwO/kAts6SgYoHVnwll/PWO9nrgpX2XW4iM7a0s1oYaQEBLp2U85hS
kvQCxGSL2B8jXb2vWtoCgbFhUvK7oktEUib6QKbWVY8GAq/507V0HXWtIvX3o5U0
kmEWqv56XyXYZej7Sz6nl6197xxQ/JJ/fppkDT4BVzkrMyGnrtsFGLvF05f/7C47
qB24St5CZFqDgR7Di+Zw3smbdIwiWGQhdSlMK72OOt6FryeCPU6zfNgY1FdlxFGN
WiBZ4IcYKu+jlIO4KAqx3HRfkM8ryqIThfV8Aa9NNEUPiA2bvGGvgt4oeB0awLDq
WXFFa7GI9WzvfaMQvx8PqrLvNcvTgstjHLWEGAoeoi+OMC+z8/MuNc0aAopYHwG1
+GM4lh+pqljLWeUzguJg4CKWrOzfKGnhk4O2yppgUtD5IOtNO9kCsX40tea8zQbv
5LTgrYLNgRovmOY0inQgePZySERKffQmh7dlCU2ERyWcAOIte5ogzL0X0c1aH0n9
GDqXhCUy3Kt9Hdz+RYdF+bYf6X8OMBkclI8zvPXBW0AS/KFyX/KCdggsp6nGlvbG
LsJisi9HlPAwjHrjgroeEqSnc9JhiUfqUwGVTo1/QPcV+lhRL1PJQxPgFr9wBC8H
KJVVpvvhS8nUXcUMX1t5qXOCMoXi/25/iGjRh5yu3OUj7BEhkeBgIknOrjhQySZQ
oQS4seeVoADqLSHXm18KLad4ZPvcKFaaObVrT5PSSvYxM3h7ovwifFmB3ZP0OYYM
gjopLxqEpe7kbmLF5sn4GdvoBNKVIQVgZ2CD1y6yNds6L/O9AKU/8oMf8Ydz44Pg
r8qso1o0pnjrStvjzW7qv5T9/LFXo46Y1m7WKDZZi8W1rmdVGEzg269C3le6227g
JkhmAxrMrwybnRtCpU0RhhjiLUEIDX3i6+SVn7Jr1GeC6HxKyCnEA5Y+Sqd2E7um
cSu+z733LwaeSa2PfMgK1cFXRpSsV/ZSCoHpa7PMp7e4j7lEjacLoqWYuhZiHih+
ZawlKSZULt4p4xafyTJ7sfGmZXpTRpzJScex8fqQZcxwAyEjTgaH7qv/28eXshab
LKspz3GB0OYD32+5R4JBxV07mVrz60ZpuMWayLufq/utTIkYqiijII76N8j6IgO8
tw0yMEql/9ON+NLbzukAzwNQb9zSaLuNW/pgeJDRT2Uga/tlYoAYm8ghZHYQBGb1
5o28F6Zi1EgyWVr5u9oXUfymDBhvf1MYBASi7phKNDMEgsaDey3DUkXQIde0NFU9
4f7JeYD0jfwmM68gTbX1AVS//uw+8IFKJFHDzyrZYlyv3nJKLqg3ypQZuNuutbbX
N1Bg6Huxxq5wOD0bceZKUD7W1zNZXWgSVPZJrKsNO6Ek0llip93qm2LXVNjT63Cv
Gk+5wLi+ZXKW+xydbCJj7bH7RKsSOCmm2V9kVPmswKDiPtQB+OGTIUYxujY6tXEA
HHQVwv3C3/CJlsNJvsu89g/+Gu5LfuQdAr2La7eNEnG458wiEX0StjK6mxB7Ia7W
EHFn1q/EnOtcc3Y/2azlhqMgUleNkUfwSaomWU4BWiRVEF7z7N0DGjnSInfOdN3q
YXssD39GXHVZOomybV8s6KZDDglkRNlb4EDxwPqhaqC6HopugTNnnE+ndQpxiebU
jiURaWTu3DKDWla6DL4J2/lFQsrDKNLJjvCWOiSO9fGYCsYYTpLOJGoY25djZdo9
d69jqd/+LYDCo2fi04OCnZrN+SHG5C8iDBVrlyNh1up02QWpNBEsecRy5l4ddjWa
GpuyZa3w5Lqxte/QpFqZzKvRn5w8UinnTrR2AzM80qLpqwSajvEoa1WEUs7uavVW
T+shW5hTW9dE+jw7rfPrpx2y2yFk87Av3NouYOllQ46z4GVbBXTH4kUCT9JAVZiW
qmek1+WUthzMD4Px9qt7gjx2bDRqKO3HdymbgHqcFT+MT9q4LNm0sVII+81S6cxg
u1bIB5pIjbKffsZOQrAUmqIETRg9cG/qdJkS2z3egJpHafih3tpdSdeiCeV6EPFk
FFWLxaGt/awFlKwixZKffozDJuFXV6Xj+y40qGn/6tA/42V53HMv54nTQ4Q2vzHv
0SRE4OMAloKU9uzxRDotmQxo5QOWodQVDH+bXOpdR2RBgpaEbvkm/00nuXvOdsKI
z0w2FAuly34ASv4Zcy9dd8m4U5oNSSI3jgDxh0pwcosMpqOOTvIJpaar9s1okTl/
WXsGfIIiOTcJSqOHceuJRqNBvZ4TFD2FfQLkdufryQ1RvGQ5kkSrl6036G/iTZeu
VxTfzC+G0qCZgvQWSQc67BhBjRWy7h5fWGkyzyFQ8LRRyK/1zBQ43g7eGMiZoG+n
KEUX8sZgUHIgj3VGhN5TQ1c0ahLdzYGR7kGKkwySh9dwM2YQerG6JXELMZXfqwkm
UjmnmYORsv+GIjO1/UHJgCwmIV7XeNLy4mvVMq3mIUD9v4Ysb12DvUxeNJtgHLvZ
UDGkve71HbJnzyS6VqdgEQpWcZH3aBOCa8cKx/uU5WUvKV3BvQ1snpx3hBzbiv4G
x93QotKsSkdZWsTyuuD0zI85BanCDgpQQauIRRNbterRBwcUd80fizqS8EpVFS+O
GgWhmtL8vwK7N6tYBpEbd0VvE9JGNvu5RMa/I3hFg19y/5uPvtLSHVlaTUmoQEZZ
JfiKsXU10mKCb+WebHfwtx888a2FJ5vw1ALvMex3dJ6DNRpcxpNvmSRKVpWZirM4
3WH2oeh5/Te6J/B3BfxpO8uoZCblnqUON8OmBTQAPVkgSI2TD/8JiF3b3zj9SmnV
WCHpnlXE7ol1oJ+ecMSNTTRrr9UfDBXXco5fznhYEk2YR3ZMEpzL1qDBc94snfjo
4CjkT9L+C4v+nF/vZ97TTaM6VFe6e8QdSxJKr+Lxthu9ZbL7yMytcxfT0CrUFDGW
ljzqGY5eRPjwd+y4+tHgf6ffOcJilf+fm52bKMDGLfzNngx1yLjquTQvc0DVX5Ej
9wORYPbeKh/WUEpwfZZNZDoFPxb0yefKB7vwdyU4AbtnrABOxMqKRzPdOnI02GhE
mcDteROSjXC+SsZzQ343H0KfCaLrcLdV2HY81tWyxBBrCZimn4i6ysj3YgRfes8U
1lJelDUeWMhhM/EDx6RNKWpFaqR2doRm/7F2rNcJqs9RezvvZ/wTIbxnGGEgM6GN
Ul5Go8Z/kUG1YiIV/M3YLSsEA9ly4nB+o2nhcHqra1TaQPUD3jZ6WaaCS7RwQO7Z
iqlEeLofeonLzTNdYG9p8wTUruRC6LJZp851AIgsY9+vOXNMSh0e5PGQTytpLpz3
6cTO4S8ndmBA7WdjldAmeTn2Q0o/67t78p11729PW6j/qWcxu6H22/YWgLhJGRba
EiahruhJOkoeBawnGd8K2xUE9zKcf/yrnvg9N+erVIoL1bOYDzLdCl1ET2SmJXZS
m98VY5GJ+zJL3nEPV+meot8ZmAmNEDlNK3QMNZ7yGcslvutHi10NLIDAeIc5QBYd
MDbSiMv2NLOUDX6KuKn3+gQnmAQD6iXAgqIwU+A1vfv1aJsLD541VK2FAVQYPKBA
spyIU7uBh5TxkHD1FtZUDNJxL+E3wsSb8H4DirsBK7GFr2UBLM4+lQWJulUwbUdW
wMTPMaeK6KVmbgQJDqdTVg21Mz4Uz8lK1bFWnYqB5/VWwz8vFp7A5p24vllKWSbJ
hqg3pTBIdKB1OTd58L3zkapmYWlsQdKHgVAhqDt0nIvedBQ6W996d4+yyC+qzfUR
viesJ/8LTh5ZLSkRRT4jHuRymEfH+juh7TUFRjpfj1b+aS7mxn/0Paw2kxXuriQL
nlfPhoJ7d1Mv7os/Ld1Srkh9djYqDFaHUj6XSkTe8kmvuBYIu+r5zAPxj25ezL2k
XuZvhyyGICGLCjGqr5Ago4CxfIWEFjTXNSKtoo6W4pwoa/SIFCDKUAvEf2cbUafn
5DZbmhfA47kGJbhK66zrd1pTLHX+rLAmnJndohp6mjbQoZZozloQjHClxVp8JLZ1
MIWC9fiMxSqjNdRmRz8rjy+3wffSwtXxHGkewaSHybb5XVq5EbeFRarXqdguXlb1
07ObS3xmNl+407qLRuffGfpBPUkdMSZkQH+EB9vndpn2hAGOvNJIePTEMgf7ZEfI
kOZSMAJFyOuNTdqL28eKsq9mJZV0n7KdljRYng+n7VVylQ53le2z556oes1qshHA
hFs1Zx/YFUCCemwGhZ17FhlOmULX26ZZgb/e3MiY8IF1teBy1Z+N2mkMzyKP4+Yr
SUkxhEEmGU77xunIvmRGlSvW9fO87auUiMYUEO+lSJ6DQumcOEdR4wchfD/tkvNX
QwTNZRSuYDp1DwfqmntGKGHQhQfTG5bP2EdUz36B71XT9hGGn2iK/dS8a8SRwY2R
y3i61jpsx7FuIPPS858YQJxwJ5Tr2d/nc1heqb1NWO4HIX3EvwuaT00H0jen+Y8L
oSacuOFf5vQxE3rkig+KJ7rgeyJxrmGycLjrDFcWI70E6ktPhueK8FY+HaRmj7+3
fLuPq2E4zR5wtkhYdhVP55N6ytTEcppkkKH58AmGOiillzA4WZm06VEUs691ikYW
Teji/IYJ2WGBfQN6XpqgA0mtVRxtvJdquiPCONkQLMj/nweAqRuEBgBFDh5mc3dZ
r8WzcRalws1igyT4Aqh10LnLyNWy4aG4qeMoOPfs9AC1iBXwpiiaXZ90EzhmbOq7
9KPrCCdB1IxGFdKcNR4szFvMxqzKY13zzz+LUq4z6a9SgfS/l8P8g+AMhIHFaiP+
8wxd28KFftrDpTJfWFG1S38zamBQ7paFGNfC/x07sBvCt/15llZloRcK6lXrN8lU
3GEu5aS7zNk7hucviN0b4Mk73DOiNpzRMKUYsEy4J1PUWvdizmJ3o/1QTu9zcaRd
0ro5AovNZRwH09c+36k/ooVw7PNIB3j6mbXixF1jq4x8Ds5Gy4YKNl5v95BtfXWI
/C6PauD2d2xrh3uHQV+iC0x+yY6scA1wW2bAU4gcxEW96ReryvRim39PywGd3011
dlbVS7vvdTJ6vqo6rTWqUsSUv8xcTUzzpPL8Mn/5QK4GJXz4et7YBkbRbErlRA8P
zFRUhvjAYHL3xKEchRMcHOK1iLc4tXA/GHdvPzt2lh9yOvryh8Gh4JvqiH2n4vva
8RDmq+k4v9LBMFa8RSD9ClwSVYUSTM6qkS8ZlKFOjpxPE7xE9U/wOawwYon8/x0o
//jmZzBkJyGq8Q3lx9CXO2a9qN/oMbeDd2u70CMwsyvvh+pEL9Dp7mBrSSZ93prL
IZmQf7lTcqP246AEbl8ER178dk7i8wIOySHgnt9mzhRY690rHrwrlLenaWSfS51k
7+5Zt7nVlUvF+tOXB566wiUmTKwtV7kvZNm3DEPtKRkd6oO84ZR08U4REje3U+8P
rgYO/hrMQon1+76XEDmAlhR0DDGMnuShsw5S/VB3rrR2L2cpGJeL2UWJ7ksTPDG/
oYn4idPbUSEmNB6YnsRTlSb3VTI89ReN6iWAimNdL0muZzazbJhMISu+Z/AqaVig
FFSaE1fmqCE35jviGJ05N8m37tBrdlkChQa8f+HUYuu1opK+WRHGxy4stXUk/XS1
a1AzdqG4ZQlKbNfoa0i2icNALfHlegLCRuJ7lCkVUI8DAr6qOJ6ymTwWZdHt5FJd
+NtybO4z4oFokD0bk8O+N0n/EvingaoTb6ZuQPGPFzLhYo+N/YbKaWmW/hxtkb88
l9BN1jamxRUf03AHvqRndUue1UFS+aB0wFYArPKZYIRZNbQG3l6r243quI9HDkEn
LafhI0brrpvUeUfxUdRxVuC6z7orPzTvj0oh5vnbYvribSG0asvxGrPE0EcJubAz
c9hvG7zxa/bA1F+Mu/GUkx0PGj9bxarQkpbcusuqBYQS7SP5wUepjMmqu4rsvuUo
sR25bvMR6ke4Y0EyKMZPswAMMdQ/8zJYuArwosCrNPGLs0oaYies6FtfNRF12o68
gK9RAgXf2nYP+D0L5GkH2mibTLBBwVces+m10ktSH5JaHbqGYfvSIEKt2B2JqW3v
gXO+Vsvfl4WpBNNTkx5MSsK8NsXg4WuD1PsPtWQtQEFZ6CyRCyrPBvXdtihRDv4k
c2xT1n6iO1AC7VPOxy2L9cH7OMKQNGGrPtA8DjXtBYAJgyzS2yuJ0BdVylU6nh2m
ZtqDoyLAuwiOETcTwsIatwigesQxGOIluVQ3MjuARL0no491NmQ6K/TTz5ZwTHC6
w065KB4XRmj5EZY/+vvoCyCTSuqT8IDCLsPaC+0kOOar7+4iuyhsXC7j2UU3HTKq
ExuTRaVVl54/ZQBGEmubZqWE2e72Qx1TeWDAkL7BvrRMxz6aV5jlpBimJXFyXTDS
lZ0E2NYuertn/WeRkZvhd+VTB4SNpakyxUWLP3yJhOwkaMjE2R+sdhUF32saVG+3
3HeJQ9Kno7RDkWKuCkbDuNDCJ8wWyVm2BivEHAQBTt4h8afE1oKUq0gYkatisdKD
VUrhXW9Qj9zBAExzMN83OdRW3lt2vm/W5JV8yD7FopVFa98HKndsBNdL/6KWTo6G
6idv43bu7raLv6fKKD4FSRrkObtMCHx3MkKgudTkZWC25MXDQLg03udWflV4NPd+
2qVJFGoHhP7lcCww2jhe+qdmHYVrWOoA0AGS6E9kQ/eSNA1BQoFg2wn6Zz+rtu5K
Vz+fELMxEwdoXk4mzXHMOJDzrAF9wjQve/VhR449zhgwIrmr+bv2BfUQzfcUbXW9
JAcECEMkvoxawndLaBiIjnnA1G2MWusTopHuwgG9GhGCB+/jTjwH4FP77biq3G09
zARDptH1o/gW8p/pk2mLNYza0fBOukuesV/z3v2M4dgBKaSa00DVjFW/RdUPQhMh
pSG4R4XyPMkJR3Qswxbnr/cCHrBlbVKY/kP0t8zdJmIbEa6auu9y1CpyfyH5btdM
WLZEvM9E2kIaaFkLE2OfVFj14diKgXzZU/2Uph4j57w5O9mGoVcDuVBO701Pk/uM
7UlzbrPKfWFIRuTI0dqY0azMDfzyEHDluoJb6QF4XFa8aCv7Byr4b0er8/b15yUi
HEQveJ8QCFSaPsQK7gsfCRJyfFEPgaTXvc0XGNFMbQtRuk0u/KG7lCYIkvEc8R1D
rFGMTAOtMh0pCrltz+NUDnq+o6MLtFUXcOqu7SmQknCaXFwwsGr1Wr6WWoTGxMUg
TqFCx0AjO4wXNBWqMvdGwMl186nKyUIJw9FFiWvNqK99/m0IyTV/IqxGz/vRdkOm
qYvoP4HrULoseXuCFw0EHvlcaQFrFxTdapaVfAH8XAiU+0RN6MhvHQhl8UzlQUuJ
6Z3/MvLwY1SjV9AZTePSLgnFMA/sIniJbC+XwUNdkR65y0/L2CPbsu2+jf2NlcEB
8NNhpl2pT4aMcyFIw9ZSSgp32IfyfKcVcB0crID9h5GnI8Y7o0i6UQipeftWXnuE
9KnEjPyzDgT9NrDPEO0fSuaGhXomzNKApqXGUqvSAr3bV5Dp9LZFyS9B5SASpI+D
4SVdAuhXuM6YXnWGsFgjOEQTaI+FYIiq4Y97m9SyMmT+9mjtOBW/a05jfs5fhIGw
IIRI7t1A0aNDEKonn9wFZECbxcVo+skDM5O4Vqzfwl/nLx/3HtqW6pIoCHDTxU0n
3nCqPWTlfSGJiCGosQioqi7fAQ3BsfusTt6413Y6kAN67ClKM/1a6KrlA3k7PR5c
NAOQJrypVca/X9l6817974pZ0RSS9W5Y51lNjmBfBx1Z/uTKOBKwf5e+75VQZQ9A
O5wfSsRGBsLXAcPoxGGY9CjpUv1gue068sKSK50q4UCFDAYVv91wWKlPGtbFPaq6
0CXcxiWTIu+Uvhm1rbi1P9X7f2LmN87og/cMVMHHTX967K7+zpmwwkF2WuYnt7YP
Tc4nKJGkMM7GOqDK+3wwWfVE+bdBTiesrFwKhCZM6kDTeCvl/qYxpgMgHZFh7ii0
ZTyx2+dkfg++0CbBCCmc3a8JVgC4DMwA16HVvKy6R388YG0ILN1D8Aai+pg0mcmn
Z92oTxVFg5m0KxSimN4+3ObAnevAcsND9nf7puHs+rtqHE2g15Sje7BclKrrQeMF
dCYdCOhVOP7x+8AK7fmJPjnuSmSLJhTs5LpuHoYOs8jnpJeinm8iyCQ/bNdeIfdF
7Kn4RoXHEshpuuMwPsVGuap3O3etNk79BybI6y+YyPpJrnlb02i6OsgmqnzP+k7N
chN/QvwTm3+dObCFs3a916TsmIcz/wGNi0ue0VcjxjSO0My4YVBrQZrsOX5hMplU
Nq+4Rf7OQmJcb+P+ricGhfQMD/qj+BwclsN6+bBKOY9iC+1URE3g5qCsgB/Kkumr
LTfLOERGCSMbQAa9gAdSXqv4T8DQYgREQjkrwmvZSshy1lOJerh40GZw+bMG1I3G
c1KoKAev9b7Cpo86CBeiPhZLTLL8xOki99mKmgEQOTc9CenetYE35Mrh9MApqD9u
PVv7gdt2MGgL/YPH5mKMJ43vg/nn223TWiq0Re2rEbX2hcPj0oVJtUx2di+/vk2M
wjjLnRErkZFDVgZEgOaqhA==
`protect end_protected