`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11328 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3b6eMZvf+eQ8z14wALfTJHs
q3E8aWgVMNpEXpVH8GIRPzdig6RQTDao0E7IF050lcnDGBUuo8smSU3lxCVMCwZI
D73pqLhh3mNnD2tU8PLH6Hxw73vdtpUi9EfNfbSppKm/b1TIE1ZEKeCsC+1f8ii8
O+BDX+JaR2Um3PrP2AL1EgUIxQ8WX4+kuZDtp5uJdYwYy7VJFYjH4x84Mebx89wB
hNIEbVZO8f3CETn78Wc/r1Qnqh/1eH7C93gMFkHIPyYbhlXSCGOH8gz/DMeD52PO
VOMq8qYu6d+UO23xAzxD3kw7MV5ip3XIX6YQMdsi8MSeYJqtdhW9CovkLAVAlE2f
mnPCxZHKjQ5zFU/TA6ucs2gnxGm6MDwy85fu1Pi/vADchelvq2TIZgXfDKvos6KF
pppsM0n6koQ1bB1btgX6PB2T/myRs9sMIQkG0GQ+TjQJ1Fr/DQ7PNjqlFgofgWyp
L0ZT3cKKApjdPlvZ/LaAjJMZG4wzhsIqx4s/dtw7BiyYWSsXnASpiEE5iMBSrZ45
fI7Yk6XYkG4VGbrFWrPQ2LCwO1nwTZGGuycTarHaX5/FghFDerFW0qVbZmpMpPid
gLeyZjObsOxkoig/bJTqqkWz5McC5pFHhDiS7kToeMef76CMge1H6JskVDeOGUNm
dJDffDeJyqcnTTc0Ix++6iLiM4VffZgem/i8EPqMcB2Z3zHMC6eTRtDdQEeoWKMa
gaHImrAPMkF5hWWqepdOM1wVKGIkWIA6j3Rq15wpVqHz8MAAtk4ffdMSVaHmn5wf
LahXeuLZXnaiPqkeV/NHtYg466aIfXFJvzpJlKNzbit24Wpp7H7aBk3TkwDqO0eg
xS3Ywec+GfXUsetnx6bTI5A+RaabgewGNo3H514Mr7VlIr0vusyMAHfBDe4hY30E
kMR6CnQlF4vXL7Hs3p5gcwzigd97u+GI00924utek3iaRO9tY5POXgkzmD/FH1ot
NZQjnf7xfyzfbP8UI8necNI9rXYbt+2Uu8Kla1OZZG+JE+uJSotbnIUfmZaxXTWY
xvmXhnQmDinzwGc2kYX2VuBShIQXwJNqVaue1S3QCBqiMgxNkmfnm656ibNl3+aH
MMM/M7ejzR7sajhv6TRtQ/3KasPmU5Ez30A0LW2E3wCTACPEfG+zPLgeLRh3FV72
PTy825wPK2hNgS5vOA7ehyGl/1oxaUkK54RQtjJYwQ8FjR7C/8jxU/wIxw2VlPON
8ZkcTDM1ddQpvynj4xn28d/1v8gH28FgnoDSjl34K0RGZcyAQCVs0BNj9CDLg/p2
OMrnZ3mKiHM6nq5kaZ2kvPggE64ryUkHNyQ3LkXQBy70O8zM753VK3K3rdmsXSIO
RiUbyS7PmyBJwn3Ko/rGC7nuAr85ySZ26sb7JP2gO957Z/YeBmvVlw+/pkY+RLRT
P/R5DPosq40eeJSEQO3n8FhdOGTuS8w0i563QK66y+2U9uTAMRXDBU/jpZT5U20O
LkHH8Mw+mdnwhAp+6G4fEXOqEGJecVWg1RygY4L+B5nXOpmbpNlObpIJkx5BMVKr
jAhk6IFVPmFSSlyI1kVOHwypSwLTNfBGvUBtcKwZ6c97ZOVukL5z14kIhlKJCDws
9GoMcaKUWs776cDxu0LfvcO9lylXGBHbtOcRLFLVGJaX+QC4fTcgFX2XJL3Sy9zz
dBG1LSitxiUDPw1ncw2NP/F9Jv0zegL3vKdSCQhBkDaGI0IB9k8zhRsmP4QaDGrQ
3hMhv8aVnpP57YVVuRsnumkxuCeXa6XNC/JzGFZ8vqvG2RMIFMbg4dQxvMcnGtEL
3crF4/25iTH5M0v/aeO9XAnXUMvsg3q3/ieQ8FaIAQCLBTi8A2NKJxgJIANC070n
ZpyAXMxRqHC/Vomz5aeYcuMqXZisC93+Cf7h3k5c+PcBvoCLs8QVWl46EH6eF8rL
ztAhdo0X7xM1qcfL9JzmpJH270pmxTY+eXRfmsrBcmxzZseQNPZkVJVAXST77I3w
0P09S812cOxRjPEpo2L9KmzQzM2NRifJ7ka4qNBk2GzMXJiPukQDdhU83dPRLUzp
ukGBnrJnyhSRtJglalfoMGIlaN/mlYkRfn5+E7Ip0P1l5Q0sXak9bE5EQxfko7sw
T3LlZjo4rOANrxGJAh6IF2oR0XNFlLhQIYIlOVMkZjUX5xITyc1otFJpd4IB5CJ4
MfMNOvxfCLivD+SlZGBvnkDfP07CV7NUC7dbFTjhcfn/ORRrCsG3EjhmmatZgkSo
t7Mtk+/tM8fvV/nLwSloo+OcoBnfcgCkBlrneWSboaG+SOQ+AtSPEvwyeqQZc/3y
8thFFsEzKwlSVCQqwGqpMkL2Xhd3xVaLBuZzOudz5Jp7ae70gJavxeYEhVPdShWw
lfG1CaLnHDYRBs+HFkJKn/mXjGjeopsYvE9fGuf0yIWoM0NrEzBXUlgXxfGWWgnu
399Un1kjjdmbBuc99uHKF61r6/P369G1kKEGU+mGyjXWKryrykdHsayH69fO9g4u
tthMnfiQQl4NFrRtcZdTvNwbrHPBNHoMJeMFyV3CfmU1ModMzhYdND0pCBLBEfNt
uC8fhIF4efLch+WeOz88MEES73x++gzqZlE0s2475w2aAIZIwiVRFitdZyuZAWzo
OUz5cuOLk70o8CDBuQY7a/BmE3ufxy7lcQyjdby84RQO66rFvU7aR37wedDM8PC2
yDwQDyxVtoNfBhAg4JPQqu2vrsVFW6Zmju9AHBrSr+PxVNPwn+pQ8JzLU6ekgZcl
sho/MOJ93WvzKc4gOJVLw77ZDyRihXlIdiPthdUr6mCHjKeOZ4XfFIoJ8citekMI
IZwlczzRaA/OqrVvm6HlJzhIiUyREWPg+2+EfsWTbxAjvUg9b5QLcHQIC2lnl9/I
nge6uIPC6N/n47KbPV7rJcD00ZZgxjtKKswNAKWpy4DpQxXpiZnwOeIgeChoowaN
P7r9Xar7DWuP2ACikkPbyBMBQHed1glpJv8dNN9d6YkbAV3MPztbhecYLjw3yfci
EKgsD11rdwVlL07LXvwyHBZlqFBZw4ld6OwObulVHujwZhj4e051CQkBo75vPOAV
e1TUDe/1Js3NxPXNVRHY2nNkdYNqx6KUXa5ExvYQVq3SD6DKNwcMDFxNgNTjMJyn
wMdqTaoQV8jeNvYUMg8cxud8MXZyk6qLcYOBFosu9R0OC/qzrKPRkOkw4WdXzEUx
NRMMlnroC9/R78w30pe0jd1fQOcE9fSFgEleQajVHPwMZgrcHdWfALJhFUuwCtD8
6RzVpaOCCrGt0BYg++PaZ2eSvrLnqYDV17aKQS/+lQF1fp78al3ME7367OWs/1PG
qSn5MOwclcU7Pr67NKh3Y+cLiPpeVJ3/fvC3rvb5IddCalayenVZhMmBnZvQ73su
EjVYeIdWi0KnJhCixDi5RFqF6K7iNrI3Kr5vAHHu9fikw+fM7xmzwArQj3k6TAQZ
tWQbY7QUuwMrsK4nkSvfk82u/LHjch4O5UOWN2b9XFp2L3HS6zcBJKCT6lJhAt0g
1qj12Lo1S1AcIihOTFm04BFkfkIpUHjgaGTL9CT9/rZ/EUvVWhvPIjgf48kOQGxL
isPo574P5yz7fMJB1nCip2dGKJkUrK91/1rdhoiPSHzAnjZX91x2A0qACF+x1QPa
suTVUwZPAZ2x5gls/kCMFzEPqScnHmyrsUGXzD0d3x7RgZ8HGzgUK0mTAS00f9fT
PDVS9nMXkcJ0ecz8BPHOpRk2cfLAcpE+LeiRhoi7G9OHUslu6V14JQaC5CGS0TSI
G/tge3L8pzUgo0ghwOuqifRRzNcjmIhdNHwedp7dWLVmDMgCVjCtS1O39C949QZw
pB804D9jhGJB+bqESEAjGKnPZSnVTMCIg+QnV5hwnfPudWAl6wFSn6dp9/dDlxX3
SnKFqHJE56PxDuTT/A96fkj2rK9aTEvavGsLm+BRnOIx2So8anPAfcY8TV8xTZ0g
CN10qOvmq/U8gF951DTDH0s2xEZgi9wG3SpfL9cTqvA6fElnEcPxiY/dJsFT27sn
RgVshTwU82BVX+4gKI4pMguveQIkB+k8OL6CUpdWakHs9mCz9MRFzvUq0JiInRXp
aSzdFFH/nzgEJn8jvjRZva0hCRAEmOHOhBubunhwsZekenvARQTpp77fJL/V/ypm
3GhlCCTOyxtv34f5XwUwiiyn1bLhrIBZxBQuye23gKbIaIEptjinaQcNpHVOTDMO
COgRT6tpSTUgPVVIclAeDtwUxJdQiqJE/IMbkptY4u4jO/slyzAFYfUNzYUgOn5B
/yo2QegW/q8K8P9ilvMw67MScL1e2EWBxm7cG3BQlXV3Gqtb3Q2jZ5wzrRplSMSl
8MMYg2YOUOI5orr1q8cvsNeB0hHj1mWXCfdXl7UzXSkrCraWDjLmsG78Rc+M/Brs
Ph2rcnOd2q+e/CqwXwIck9ll5s+MmPDO9KMRBCh8msuKFmAJ4YAbFTDYMuNJUwfJ
7giHQ+IlacUGOp+VR1BNINd/3GEcAf/9pg+sLZVsQj7g/sBWjzFCU8e/LlTYHkLK
vLYaJdM88Pw3+R9xIsw3V3qp/9owwVOxbisZyGT1LdK+cb9y2GLfJ72/n4Lep7tN
O1kaRj3jJUF9KsCU2Kf79N/oT+NihVkenOf01d1Xztaos3AG918dFv5txGuCNh1k
KRX6W9eSIDFz/tqFEbDjWlFdVH0ewzOleHLBgsumDmid2tZhhu/43AELrpuCr4bb
5P/XNOXDMVQQrXwrEmJe0jL+xcI0aKRkkaYSzKjbp/w8ZoQbTI7WF0a7QkSCRuo+
f7LPfpaVxuxHiRJzqZXjalc9Mjdac4icIKUj7DPpPfZT+nc+pHEjsGCTfToQBcST
zSldE27vCxs4DOe+5L11U2GDi2V0TF1jwkD9WoTDfS0a0manGxkn173fdEt1+etF
4JWuIoqm41pea2jq8U3wrsrYIS4lp5ct2TMlwVqFRzq8Nud0vNftcI/Ak4Jy3Ak0
8n8evMAcpqcvRjA2wEqcCOhWNXrW1jKlPynTgRu4jwyvEHuLiO3Gp7nXddoKMI+s
mSSzq5K+jzsIWsGqLes1ubmnehnIQKx2kBdJlg6ldTrufl5+EYrqv+bN6hjXr4H7
Bc8yKjaZmhBxqtGBU258vthoE6JUJBHnF0cd9T8J4gs5cHzxl2MytFRcCmjDvGpJ
6hM4GZU+rbVYSI9mDAceHCMSo/2hACAh+Vyenb+yXyYe6xIsguwhbN1y8NYM+NZk
4ZdxxPDZPrYA/LzwKwW4TfAdAROTuPIsyIK20L61/HiIb8HPlrDLlusB+T5KI7sV
FPH52CefiZQm28d0wsInN16lGooE7VRxwUhGLVkHxFvxQ+1/SlVhUVWL+QtIbBE1
Qc7Kf/xzJw96Z+o1O2cXXLseqk/MIKTEMejorgXrxY6oEs9u1pW/OdP58TohG1dD
BLSCibnm6uK1HdMWUWI7jKfTpaVMzuOokOO0ytctpUS6zHjf10WZzpu6pFSeNwC5
2+C6HY/E7vU/ARAySfO2DCWNGBd31vX738FQnUe00IAYfC8xGAoSPiTl5H3EVoMF
35CoBg+yAPUta2X12SzBJvGkoqEkYTZBU5NK3mEGgCijgoTpaZ65LP7CWYRYsf7R
2WEGegkLqmCbOh5AWEOMUdyIlPyxp94ODsvlJHGhUCOcX5GTbRPr16HJhCcIy6NG
tx3PkjRnv1NB9cLb46Q/3d4PCFOnLicLK7NZ/CCwzfgYPSFV/28GM610nNPDwrN0
XjyZf6vZm139BT7RCoIJBlhuWx72VKDKZHI9wOO+XsLb3MOdBnkcP7C1hJqHb9hU
XWMnbweemzpzohCWa9e/F2GrHTp4xmSB84kkrQQP+qYeuc5H6Mi4514pG1mZQ4XA
kcN7UB8DTCtCzuJViKtgcHXtxiaWXLY9loNeZ/I5+XkwcEpCPu0usmw/lwiMMUu5
XubJib+o6TVX+sso/wnRLyo/v80nNamMd59kAjat+aByE/zYd2wcKSFHqmQ+SmeP
c5v3jZyCg2iBjYFobjFTeVDZ03BckSerLRVBWSNMisKU2HIoGK6p2I1b0M14oiS+
1S+S+77GTILW5ECeWxTVVHZK7Z2/9Yis11kyGi7aD2B7oXEpa35GGVIn80q715pC
iRwCc3HRukBvwRv6Wfmjs6t6AtIyXClyM15q//rlckiktmD6jWNPthGcFiqbP9WA
gIvFkSmM4+A5UCXp7rHn9ePnq7DdPkhFqBsg2ttBoXTjmNFHbrA0/xnbPfaJGsH4
xG0VJoH/IVv2YianOM3X0haPNANTwC0sSLL87t/Vq6yRgqABtiP6V4Xc17zBZff4
RHNgXUHERkqkmdRlsmwhCZtFMwaThmgorKrmBykhe1ZvMDydDOm5n7W28WfmulJM
bX2tO3ahuZIhkNzUP59oAgsCiqZiQJooB8z6ysdlO7ZinSGsDXosR40dSGPPkp9G
Od4PQgTN8rAMzol1/hpk5pCEVcoJZ2sKdOTjwVUmGc0bDAoCDAqrZE4zwXY8SOt1
wXvO4eogSvam1zqIY2HfVh0nh28xs7yqMDPWwG4q1AHLnt4g9EWuAVd5tnsWsqtX
NP8pV1IxgfqjipNeFnn/SMJimNsng6aURTIbkUgsSPYM7aTKr1FppIYnlazUQOhx
OYkFeJXg54wDxwpZIdkeGNMQKBDmEtvv+U8St3D/9WKKZAXP83loEgP37ZSeozs4
x8BwxSh9HXC+MGjZAxyLsjVKkRJ4dmhmM+ncYSc9kWBs3IAnngWYgpbf2ySzM6x5
4nFnYsZdTe4DfyKE/ZOFmkDYkMElpFIp70JuQ1XV72CWBXk7OYbTip7muI2qghTg
FdQ2GlASd0ClY7deFTbjfKkrsiczDdgJiaO0+O55/tUNl3+zem7RZ4Vx/xRncuJA
cA7PCMZ1MNl81yo3jSwaDNzpfYDUFwN7UFKsbcNSw/66Hj2Arh5eXsYeGcYE5Voo
QpRTe17qUzcefdTGt4FSbBe+lmpJ8seRzNvbdIXxIbaqvLKUg9OjcmMqWs6tHqgm
qVvzwBah1iOdSPHRw9D/xxGjTBH5/NA2BfMPyEXaR4wQ7QSjGZHuqStQiSPiousX
hSJ5BdtS+t6ia0Sr1K1UeUm/M6/gDNBp9caQ0miW2tS/Vi2yqUkEIjmUa2BhAUjc
FZDI5GZuOIt9oK34g0ZsJXD7MJeMVgG0xwxjOXk8cEIiR2QGwa6JE0MoalW3ID0f
E58Qo8GKMCJRGY2dwGQzCFRg0fUY0Qvq9Nat1d2I8qXO2rjJ9/jCi5Y3xdFLjtkk
QwVEal1ttbJOr9tZ+QTsQ28Zc5UjUTL5NRcb7uU+SfzAB5UCeyOFjPAuzDbDRSpe
1gT5SKVFFUcr9KqaEnVT16qt1ThdXw6pEQHTXcGm4pYv+C1G3cs6JP1LEo75B+Wu
VChaFS62TwhN4Yxx13PIkgrJzxntF7t74QrF6l6RZwd//oZzYafMthy88fHPAYc+
Wmmm0DgBuZibPdkXhH4nUfdJ8iPg5184R/ce4nKeiz+u48JdNqD+w1bjqwH7OBBl
65cih1oYObpr3EvI6dFeWyecOwuoC3ymkQFUqWBIyOCSrYxPJscWvXOj0YrCEGfQ
6QxZgDCJbo7gHj09B0SP/ZjbpjW/QqLZp6WRuXlNCANOp4AtwbXMQUcbT/AKbX2a
jmKheix8IVWcxLv5GlxUiWZbM1tfCq31WDKs2K3Oe17IXbDv3JG5LtXhp23Hr0h1
31+MA1jIV/POv3E0EilqthrJXikOLVxPJTS1/XHnrBMim+Nnq+M2iGa4LD4JluE9
m+moXhcjwgASHtPJAWj28Lvu6bivggO7+StAD/WDL2mmKcWazTAZQ5ldx1hw0R9e
sYdIHPkNCr8My1oJF7nff/Vdl28nb/whlyrRJTLgPfz80M0V1sZJdCJDnNYm+TwI
CPgV5sB+9OITYroU9i+Mtzp9/+WIXJ4zFixHasu176RlSuAxHQWoxLGWpa6kuJrL
ygO571isNlu9jDbt+GBi8l3Wz/j0XxEpGrLU0C5ltaLTtVO4kVrDAEQ9dpwJ27cC
YUwGaMp+6o4ncXHqEpulteG7zxKYIDTlllPbvycURoBiYmCD9CpRgADnAKGiADMK
XQvmSsL0zKNiAhqjtkfSRjevchPZBo3RVGk1dzvQUJT/FxAUShD6/RGO/jDJ2qz8
u5qkEwdJkjmOvyvdr/0H837bfxLBBH6LxPxivQGbeDABmzVBxYU+6CB8acvdDS75
SdmKFDUVGn80aJAxo16hJJJxL6bVyor1eRgwBQ8/rLC3ruRTrsjYb+utUAK+atRZ
SvZdDZ5r6waxW2Fna9o3zLuaQvFE5O0Ox7R+CnIT+oZoGBiS3Ni1fFxXwPsItsmn
ftv7KLrc7W9u2aiQouG7tiEFEgToyBSt//NJrsc9HACJ55suAgBnj2DWr2MB1JoP
EOpF7gV2IK/c2sgTuruejKAJuEct6ItOc3Jj1vl4n0dVoEScfLywUW2gD1j4Eqy7
DsvRRVG1WufEDaPgUYcLwonCMFZ0FsxnEJ7R2kM0dNEj2n07hcX0vIHhU2sDxxyv
TOrU4WBvxap2Aw48VM/mS+/+F+07S/yy/tL0BWaAjG34oGhXkY0Cbbwpxa+T947J
Dq87IX/4fNPQTlYKd1/ZhYNqzkZxpi33jGoRri1g0alO5lrKZS26eCqnPGzyzn9p
loo0Hka4bvY075RjIvAV91u1sc/7Ttr9NNqvy46SKMdoZ90FCFEAOm8HsHWys7Lw
FneXNQRjAkxUmK92xvKibGei2PBviTDWzHjxxavHEZYzrNCBleALpXaM+KhS1t4D
XF2OEkQAX5QeUU+cvraFWZZrJGUBXFsm0AFCpLh3rJidowyz5JKcSQ5Cg1YluvqU
RENagG6/jmxlOXUEUNTjvjjF99KGmyEJW1ZDFnYrumLgK5NCrw7K9OP8kbkg/SFj
k6sUiHiQVsgLPuhY4SogUQdoH+/QZ2hg2b8R2Bte1HByT2p9+FtGNRBDDruUfrGP
7UKxAb4DJApVhq0qe782AYs/NhRQgIAdKwLxxQLD/CesksJyi+3KUFSUvUMswsqC
ct0wLuBNJ0KJ5+5oomtJaTlENUAtmpHouhR5yLjrJrd3mIFAH7ib3PCWCpfkyfVA
nM+lvZ/6aUZ9dLbT7pYVjxZrIM9xliFPUy9KiPvHxMsr4epe8cgC6+xSgKemhWYT
CYO0uxh220AqomDQjkD6/eaEpgyikjWwasBPelFwKX7JH/Z65yt2USTcJY3kSxdY
UGJSvwGxKl/uKMgiygP20TYojlgICNOqXtroRfHUEktaKsipOQa+WGBsy/y85VT4
kQdUWQ2hH9M+FmrvMBRR7yGEshDqC2DeSBDskLIJ4aerswh16k+yud0zPCxq/ajA
Xld7B9l7MHuHs21eUFkfg0DJ1lWiBRoj+stb3vKoSiigdrT0z5m42wPIg5GRPIqJ
TI/UgipcobZwfoORYGNplD/wgJGlNX12soj4z28zb1pdIeivXV/E45Vi1r+xjLXX
OP7ozKp+ug/aZMGCVbvSYilkUsF2an10gacQS7aPcUiTpN5qyUnG78mIEkoC7SJr
aH9VGNNl/VTopaZS1IZnSD2aNFj1uVk4DWhn//R/Qvu5PdN/ZsFFGv6OEzftgjy0
nM7j+IPSxzELlA+Tow0qTIX9od9zKixcRHsyR2AeEIJSxR0iKLwE2XbaQzJyqsdf
RsRdJE5Q69pJfrRYcTrjYgVURX2uBoIUjavvQs/mGfgQauiYwbRIHaJkEDE0ctDv
P+KmQUty4OmZdrzlV6E0brgcm/scCOrCBvEqv7PoS6yH8W1hKy1L9aDArTC4RlVz
DTV8jPC2uaITvBw1/VPCv+S5YipBA5qEjfWRJakIBUoxBOzZY6qQdEV5bwy7rqVW
Xb8q1UkjYaFw1/uOzAmy4rVwZisa5BWyivcd5g1qvnYIBnJoc1PPC43r0+13lBCl
aRi6yp260xC4B5uwar1ReE260GtEFmf++p7ZcPBH0o7uKgKGwHk7TQYhTUIz1OFR
JVVb5cO04hVVEwbNNNIQhmQrVXxzt/91m4UxYk06RHa8C6JGlH/rO6PY5XRYySkV
WcIqke7jr3ozUZsdHed4FxCidHhA2OoblVWMD4AX71Gm+AR29LjdPrXKc01hiW3z
oVsN/g+AseeIUCo7sUzHSEATi5aydcHrzLQ+R2ObgV5Hd3SaLAqvAjHg+b0waQVn
yNI+1lSdEtUtjjv4eWGy8IesJ+5+r1Q2vr1lpM75U+osrJomDMvIJy3OgB/ICn8C
w99BPtgHdDaNV5+GDs8IAhI+Z9FvEVHrgR587T63WXxdmvyOC4VxP5opeVkA/cNJ
gFGw1pCrPIJz4EIr1EW4cTssl4vyZ/U0JYATTNxn7bJsszDdICGJ4Z8DviRhiHHo
t1c537xTDQp0PsdRi53ds9R8StosKWCSAoFY23IAzhhvsqnAFzJ0zqIm7oGYURSf
w6BpZAaa/9ludceyUP5CRo+vPNp8DmwweGAX7ukMT428eke9Fca6jChY/27ssTZI
+n+dlzI7fWZyeo/YgfEdSAicJXXsrQ6530Wm504dL6ErDgxkmDTt7HUsUJ8F1jW8
JjC547OiQa4hKeuswJ78h5uSasUUstKUMuM8I1vJAorBNVdiYO/DNvfkfhJscx62
1ittup11UgWnQebaLwg/spc4j8B5wJPMtnocZMRvg1QuPDDAHRcHUhfwKbSTs4ol
niRCoLxM3GbocOFxi5H5d4kgFSceIv0LEYUCR5q6dzaR+0xfK50r/H+luwGRAzX4
55yXWRDwnwoHApl/py2YqvCW2tobsLVnHGpV/6XNFLw5R3htkw/WEFmtnMVTfr5C
9zEHc6y13ZL/an6VpaqghhIHtsP6sClnrSYuXOQTPvaB6dL/ZpvlYSDo/ne0jWv/
dOaqDt/M24oKCn1wVOvMbB3YBg3jUrNfxINyEkUO6RREboFvxjLp+aqcgymJgVle
OnDylXZalArjIpwcSi6nQrnF9maR/TBR2Ftb14MMzjnrQshObYoM68Ew7lWajgAp
etYkKsJt0rmziVYM76fm8SRFT5WpTyAcdX3tesbj6PPFjyygZyPMbsP3R+zhUSEU
lASWq6JXxw/q63BFKfycM0LV3UbvMfgad6GMvxMu4buXTbLDRJs2R+GWCxgOZ6yd
jxYbC9Mc8Yvj0uMQwrEqbCINcwm9HUnt5B8YuEysGJTh4cAU/JfpjJeU4xO79gKq
zy8vCUyG5EDHdXEuQc4T3rD066yZvC0AGizyZ3EHKDvv2HpTmISQPcijVJwu92Kg
oeonxZahKRfJ6JV03uuprpch1MgfXut4OGzgc5pJDYjQs4nXh71H5YRpJZGdJjUl
slHycWBkv0pCSsdHrMIKLDY28s+96wqQNOXW9ho4UWxJ/ld5aYvy5PMSFRnHsrea
jAtJC+x9El2jO1r1HoICe/Y5GzDDDV8pa8Yk0hw+kgYHWClKekEjc8RbzA1ikBHe
/qZkwju1lcPERvzYcnAjUjBDnNUWPegNE91lrQEFVCq19Ika1Lvdi0E663hzRlcx
Duu1+nNMJdZM2MkadDO5ib1+/nfIFcIg9KvgoFJnPuED/DbZ9rfXu6FbhUSDkhL2
e1kVPeHB8nnIML8Y6vNj+5WXR9JSqRKh8gWdugskqnvTgbTMVuwbeOZ/FsVbaJSR
ivYpb72XzWXdLcdNMzu3Ll1ZZ6XZioLhhMQ698bxcY0H+L22WTAa66RUb8njCBEC
4DyNlsDaMcWqiXPlXSyfWeKFU2d0A1Mc3K9542pjHmBHSV8Zs7TzGAw7TZnBD8u+
5xKPgGhFYqJaGHZ4mDOyARClrJT2376Fv7q1n8tkcx/04RBUvjCK3hBX8qLUrs3D
4EGCupXT8zcWFr+DCOCrBqzSkThEz7m4T3tsJoj0siu70bCEZKUVEGRivlBnS1Rg
qfBOouXoHTjOIlSYihmq4kVRdOqngjdveeOLX+n5mfyAscnyt4RhHoU0iZxGlA7S
SIAbuDAtr7vLhUnPJASMrmswyAtotmIhYQu2Fy98pHsUa9cZyTMkp8C6m2DR5kVK
um4urYRQ7kenXZLCU4bPvUMcr8pyeT/bn5MtBaS1yMJdw7shspuvFonaTlC22TDn
1P3aaDN0M3iA16J2tBrQbhrXqtxi0/3hGDgh8xA0alxA4s6Jurq4kGPTHvjz4JTU
Yt4sx2KcHBks5ORUMMuMBFDyPIZagiZIW1nmjMglzKzLbtsD+xzP/9A28XNhIUlA
YZYYotAobWjxUbcHTCnwBKlND/p2qq0Jm89z6z2R/jpm7I79nU0ckis+T4amDCUO
91Hr/zWmDFDqA7lWoMoPsWcO9S7D3AFCharjZPlYzmJpGlkA39G406lJsITwK/zH
RyDupXIRd5Gv4hVuQ8fL7IuQ8ehYaGgPyZnDPIrsR3bHX8Dvyxl+tojVygex16uy
O6gIA9Ur54J2E61iwATHUgr4Od/D3IRW+XPkjbv958ueM3NUK9SUw/SccgUgJG7o
wUf02HdCmozO5x4ZDjWbSkOGmda0PJ/s8iUL5dYc+dEoR52XC19SECIPaEhOgLab
Y/H4YsWJoLYDqK65/KPvTvaW1hSDtyDS5+8t+8Z1JqwFmG/hRZb2QAEY/TPK9MzC
KA3H8zCtHMlAjYdpRkEI4grm6L9MXBJMgBQYhxQ4AZL3HWzZSzD8fOfCttLXfy/l
Z8vRTHjyvko378+RUUTdgrhXK47ZzO6GH1dFE/bm2/KmocAMZkeTL7Osc17R87vk
DlFsQChRM7AQaZcEHrPxBvjr+wEAhk0jLyv2c5pB/5ENCuDv3tg6nfDAt1ZeLGCu
29u0+FXg19yQ2H/Lb17LjcCUYUXaMjfAw2gmjJiVwR5+4Op2DLW2TnqPfPqHSTx+
lng3yotrYHTNaNyWam6nVdXD5Twc5A4+x4KMDZyKitfStp5oEtEYjEXps7d7ieIU
YrzZp8UAOm7mlpnLEI4cXaUH43VfUx6MjdRu28Jg/+vPVEicN9uG+Xbu8aFhTeOw
PYige+S5fhdggvFtQadT2SmTcpivNEU+khzlTFHH30MNXt9/Yddqv1R8FkxLJ00I
T7tU+5q4L/e+sSRyAMlEippaNSVRX4IKEpyV01OC104wXFJ5EQnU5HYjIaefiqff
EzYwbq8t8Q83tsD8b3kea0kOkL9VAy3WNlpomcNH8Kim5alVuEzQ8QZBoYqFLfU0
VHYry8zvXY6ckvAQL+EWI5BKF+5+3WODze4eS31jQz4ratzXrbslgH4O5wFKoKkC
fNNNEVIlsCwz29r+QyaPz2JeHZ59vlvWqg+md9pEZg4rbLzCjS3xU+Dok43SbKoO
F+3jJFSey6P8O0myjAFsQuzM00oyOdgqXSjK1yUjNeJT3wENyolio5EK+8LnQrrb
rdMUeRdBzkvcwLRgauFtkP40/oVZyKL0HSrLh0DVPgA1AxaGjgxBr9eVti/q5x/U
GCg08WPbKs87vpjmYgsbWZPTJgtqs84pmsKskGV/dP/OmF92LQFezXo8PIQdGa7D
o3KM8E5gNT786AuoS5gVpXLqOvjDp2ejdZMKwVzHruHKxcsqL8Cfd6g6VNzue/Je
U6QIhvoQw1KuAGOYIJEFjscKBQGtVENs8HOyAaQPmAMsoU2+/vxAR+i0Nk3SpniW
wj0BZmLhUmrPy+EvwI+1fCXLvRhDWZ8XTwW1us0ArsTe+Od9der1DAbg4Qncx6S2
fBA9gXl2/W5SAJ8Cwf/AncucqKIH+0G6R5rkeAmsKY3/TdP+YU8E/TDtZHePY5zH
rP6DJXkPK1VmZTOygfXTO9wef1LnUnZla6fNdaA51nAaLDKS43FXvmFhM/cTPmyE
6LD2TgNyu4eveA1AQNac2tufGSph4DhVOD6xq95CglAN6ifEXo8e1uEC3oFYBjLq
/I5CYs1hOFznTg6wnnCXntPbUm5kXjFP/pp/CyFj4viQXdTQPhYkWn7nh29mv+5j
nBH4cXOlGMpPtBqZef9no4sWXGNYEWkcdBARbNSxM/KEzoJD2lYP0eJfBQ+5KziB
2uCsDiJf6GrUtzOwg72XbTS+bZJSJ4OBfJlBF69Dz+fLVBCEdSmbwSg7rrO0c3kr
dw572DGm63Wh95KisN8lo+3M9jtpmcNIkxDZAFkrqjcDqZdA52u12uLVEmI7yD7u
G+NQqLI59oqm6iu+8ycS9nE0vVN8olXbog0idj6cVXVtO2MQwjtojTAtNeBRowIE
ZLKbq9u6azLUqvDF/dVESQn+usu3WapG93CYEpGh2wCM0G369Qcbdx0CbwuzOZWq
LUVozpBqD0JP5HGeVbYKpLOCPViJXVmwczecykxR441rzbEmHkQchZrx+UinpUjr
BOvqkDunrbbZTxXdmyTeUsHs6RU7Qg1i+8LLuBJFBeU5/X8bNGSjRiHwtSg880hk
Gl+955y4mZs4aiu+jnnQih/9y/6rv9bmwogFgy6JlqbGVnOOYckL6cxKG/fz1fKp
ipBtuvTNxtXFOBAXTro8CACiUuFytnca7cIdFqpS6kB9ZuLk6Sn/r7NaSN3XSn0d
Tl5ME3R87JJOVW9Ub2iK1KBzQ8+9Owg0IPDwXQmRA+M4WlFnRk/pd5QbF4xJhZQA
QSF3e8s+8+K+4FbS7GP73GuO38YcHFTrJa8g4B73xABhrLoGLysxM6hqfIqNxMqi
MYpvB3jiUmLkVNrcwiYi+2t+ZVojDQLG6K1oIiRadp3xe6IzrSkxFBVvW8w2Xq9d
XjKCT+ldWX3kVOIJYpL4U5Vjs8ooL/tMFfSNYpp50wIuhcfpPSCcaeQGAMfKEcBm
iqAkNYnoEhhf4l2t8QyziArTPKWyw/J3/Vy0x7CBY20l0Vsxi/Iu8AFI7aYEuz2V
2U2F9OrFMn68mcMrY7/3wUhcJ6nHKWkb9knMx9vNDdigvcyDPoexF0Q3Y9i9vhcU
`protect end_protected