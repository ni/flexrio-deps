`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
GgG2UXwpbWAyDgGIJC8iiCaxXP/V0pyn8LdO+bWRy4epJkeHudCpSbKgrb7R/dzr
eMPRl97SkH2ReCPct8Pud0iGzA6MwP8/EkWOHMcIm+4z9n88oHeX5gCn2nEkyM0t
spGkfy7J2UwoLbX45/Snwj8t+PYeU3BYlpGnYzY11ad02AZnPa4IgYmwdFXoJTxq
F5mWvubueD0dUlUXyhfeF0wQRfgF9N/6pAE4hNU3/cLamjfoKZE3CSxSB9cTHv2w
x0D0rxJTkoaBCJC//XLC8GjmwvNmBlhh172H/omMf7y48jxT9vKLaqYlsGwfXY4g
f6bBiSKMuVu7Hq+Ag8fQHejL0SSV5OfQaQNsod6Da7/IueXYGbgwlaUgJE2aqx12
L7GzEmBeoyjiA8BXLjQObUEyiKK49FHDWkjENIgj/moreLpUS3s5mPPL0zXkiTT4
XHSaxL3zs4Q72kbCub/i0pOqGd+SczgoemVtFhSgp2B6NhaUmupDDAPQ0N7/8Qw7
AK/CZ+GTvxQWt7rAT7DpKgZpl4KowLQPt4bdO8stsr12+4YPEwk1KvjQBj/yAlJI
Fs2erWJdVaZjNL6sNGukmIEQ6a3Gtjlz3AskZwC7HsfipYND1J3uBqkPVcPQaGpU
jzrXY5NA+cd5/ltGEXpB6fKIvZZ241ohb5ZeCyMBjzLpotV3WUsehZjiediiMgEl
TdYiRrIWsg3T5W5AMgu3hK3nGmmEyI3RjC2xdbS4UCLk6j1K3s70ne+fBFVaYH7e
xwjuJESTwfFRtG5z5/bakVeMtn2engRMVu975FgduiHDY0NetxLlnuzrN+wJzmLD
8VmbizxA/CKX5D6qRlPejU4qjjxT928S5oJ2diX14ppv6L1a9RuFQ3avAnO18ISE
521B64XCyNMRKZktykzTuYGQYKde4UGU4ghs5+OJStNkvBz3SlvMidjB4lkWy/Vo
xVkhzfo/Er818vvB8Rmo5fn+aCraN3BvSj2cTc00DVmPeZ5J/0VPkxor5lkDOFLL
Hzq1Uqe13e5e7NgeLsGNi3511Ali0snz23zRWaVshuE6ynf4O2s2BI888vILcixO
S8dfZsA9Ot/+qlJJA1eHRrdEkxtYy0SJse96jN5oM+VmczHIa79yhq2uGa6lWqzb
ugwGKpm8O6yv6H6A4DW/EeGy5yub/F1nXFwkcZdiAcVrkwwaeM7evqyjrlXmbbW7
Q7YbCfPOaZyyWKRFecgJ6jFsKLDOZMhVyYcvm3b2LwrojFWubaGCGSrflVf3tb3Z
oF6sANogWuEApLP69z50CxCUcEYDVnNDih1KFfqvMXMEvei5H1IlaZqo7ho3MyaY
AQWhpL0qEvqRvyJciNJk3QTiw/HUp3A0tMeD3ETItOgpDNErCPy3yJRVHp9xxgNo
OOtg3xR+NJMLAfWO/FzCgWX1gaMorYJM6qRDmQlIcgiARvHriqPblfW8mBZdQf3Z
2DQr93qp3JyXCnTkPVQ6xc84GbCjl58yoTNBa4gO/YeHjegxIRAEJkdK5Yok3dGy
0hPs4Fr8Iuwkb3RIJl/REMPehyjYBmERPEM7NOTbQZX6Pbghg5ecg7IrZybJ8dtF
JkWaG6SjNY9i2WGLwi1q4TYLhe1tuzEu34Vfs+FL7EHTVgCgAsCGO4IxOanjIvyX
J2rbXBFD1xusddOOFSnceYLVkiK0+1IOylT8Pid1ROq8fjjhLzFQCf9BCbSWhnMo
49zRZb87O5CB7MbolOcHZpRlHf2Z4ex+9PFUVZmo/bG8EhOrfFY3GR1911Jvm/j6
4uzSwzudWrsKMoApIHPmug1WLtsuZjAGzHYPSUMiBqQthVnaud9RYTj4ri4DWsOR
uhUlgtSwXIM+ORmttyH8RI3xbQFgKQD8NGKxicCTl73LczWzcC4uOMkawEgA9Bv+
d0H2t2icpn/bx6PGPJXwC7OYQOsQFwA4EFEYweuzQGYcVCPIyPiqcSaDjB6fHJ+v
pbMzZ+jjtrr6ScJvZvvnCW1fwPG5YDfWHAtstsGqwSF7cJJ5fM71hmC+D3WRm4C8
QHS0/2WJYZyN9LfEgqA6hCTvspJzY0BUf75sTOJ43u022xCDkD0P3AKLM2+vYic+
NgIRNXlINePb6xxqer7qaO/gfGzqtjETXRx8O9+zRSRJL0+TiuPlZxQkp+BH8xwL
1a5vuRZ/DepBkqKCqsN0iDaQ5mR+jEx4/Kw1j9HN22L4C6VmS5ORhSiGNrz4z/C4
UX2qmPK6qX9yGRdCUTs3p3rtGxBs+IWdzuRUxZyd4AX78F8Wxj4jmSKAYvxPfrOw
aZ4NXiDYR++cUGhWsHPsFUMWBoXb+s/FU4q/HdYgck4DVlCw6yFEjpJB45xGovcG
rU3B/JVYQCXNAOkkTlRmhK/hV2IqX2XM206rw7nUbqYS6PcgN3JQv3OqouTNywTb
8p1B929gXFhKbQovGjbgfYkhqp1lOmrjoFURd4E4YJvNAjvZYWPsSP6Icy3TjpYB
fq6qmil+kPXltHneGxVc8lUoHelIDTa3g8ffuVV7fq1nuCXjWvwR38Ll2EYxw4P8
iyCJM/y8RKsTkld42FsMb0mnTDqC7mnKj2YiVRvptq7/AM4dUHD6O79u/NAXVYiU
1WUq/rkpKwXAGA97eg5FlGBUkTDv0EWXU2W1X4i5huWsvJNdO+LWLzIqDLzP2pFD
kStzM42Y4Ioz7pOdVsf9H8L6754EDN6tJttRzlb0udcK47HMrZngWWNYo7qySF/a
1bA/OUjo25ynKEpCxAdzQB1wKHAem223jQ2QwFpOv7H1I9zOqi//3bWfhTHJ7u2m
xFqAZNhWFsLf+ptpFpdrnKcoqIOj4WOAz/pgBbT2m4Kjn5djCvukaj+WbbWt8Ea4
KQUX3IRHA4afrfOtcQQeq+vIvbED85VY5wtwcG0cPXiY1VZHurHxVgcHQMaqvOX4
2R8nmLtWkzMDURUsAPzX88iGVWyTgujon4hZc1nj3R8kAzjYp/k03vE+qrHWLnAM
7JxTgZ8PNmBRTEeI39Cvw5LFeiC8WIt0PKWqLeyPebH2lhKy9eJluOXpOaImec2f
L1v4VZWu7nA6hSTXpBO5vm7CHTP/5mSJveM12KTWdtIlgPQlQ/RYGOPkbvq7+cD2
1T8kQdHRXdp6l6uS45PTqILkC/fdysjUlzn7/U/uYNfWFcwxNl1L1EVZdAtIWAry
xgRCw0Bj/lg/m+uX5UpefTXjYcMUWvZmy5tbCao2Iw/aT1RA4vBsWeRkZsSJJUot
4LaD6T3uOfHfbbTeKUXIAGro9LxoAAjTmvG+00wOh7+yLFm6Ll2RbDSkC2slnntb
SNsmqUXMXGSLF2m8rrdE81cyRfXs0HCLzQSokClBE8HYGtIFTUQ+yNUc+PgKa4z4
HLIiEoebx8fyhkEHtbVNA57ejPrXK44EAAL6lYJIsMRGX2SyCSqT3vt6EYLW0PPk
/wJ+s/VbmZFCcFWJbMLAeO4ijMuPuZHEJqeTNxbVjAG62a3bnPyN7jXLCKr3QzxX
Kibj2ik709UZB4meJ0WmLJ448qKlRsMMdL9c5J3HeafvuWBGDhcMSy98OUOWnyQC
WKzrfiBjd9jb6aFxqsglDXcs3y4nHVc2Rqh+X4nPJ9IyVUuapZTUHpzNfvMbDKK2
PPmQKafffu2Y8T1uTrkqANWxXNV1PyorbuWhlwkYZcXRFwyHW0OOiGxl2fXRuW9n
/2T9wckVYlDdEPWZ0NjoMvLFfMkzgKzavzTfP62kbvfbggSFgR6MMCcdAcl1ZUWu
IWcvr5JXRqB3LVsifHSaXs+2YFLs5nd+/ianVayt61jHBTKTBdSSRMEAqM0x1TUR
oWWMF+qJFxETTaYKIE+Jwz5leEUKkd9Asuquu6MiyttQna0E5TOJBs5n9VxdfZNg
ZylH32o7W6KlE66cmXZAwoTBqx5J2fEJw64HNE+Hu+CE1yp6eXV+HYQJT2Vei3lI
Ps4g1Ovon+ziEhyJ+HIkqKK/f7hJiVrdX/qwWxR+sIZERvYPWX9dTPeuLXIO27PM
4p3Imq5iqkSIbwV2Xg9ZgeHPjSuTbPo48fKCj2SqqbZwX2t6HYbHcUkLKVpGbnjn
yYnGeNCJbWOx4x8esn2hWcKgTrwo/ShP+UZiH5ULJoclqPrnsiwR3eCq4ZzXUedl
oE0GB8tLGf/yoslAJ2GdbRtxV/oG1f0R8OKt311OqQy1rdHgS9CPYBbgkG/hUdzj
RkIP0zsomqyU21wJpQFrlW++AKN/RDjkXUdJ3KU8kbcEETuOHMtkYL8GKchwMiWk
xtd43ChDL40i48sfn0lFJRZQJzner1ObnNiNyKqAXbeFTyndouT45uyy6hElinxZ
iWy/Rb+Zbbi27kRJNElZlt8BUTOw5pOXbxzTovRBQ/FPdpt5E9R1z2IOCCce8MkA
dvIZMnLuLvV61usqx0cZcOs0otb60aTxUjDjTvXapc7/EekkgVIQsgSq5xHirOZe
GqjcDCT5k4Fzw063A4ts0Er5qRivDN6KHmmHvl+7yiGmAjPEsekW1yB9v8irQkPC
CYN0gcnlobxrYeAAYcJNXIaY63eVlzZF+oLLjqTrRlFlXqnvSyghCYfd5G0BLwLU
+zmgn6iA9XgOAZvt18QLjwC1mYhfY77mdwsD1hrOPy7J8gMBz/8LLMnJzXL6R2C8
2xqZaFOgJx1cdZXDPOIyPg59b0l4kfivMvW1ocEzdTH/jseqRRR3/NkxefcCLOi/
qwlFwLN6FuC3DlToIwOqlmb89WipHaSVkzwTszLI++SFg93leeG+sc1YZIaX0Ixb
ZNTxXRZwpbEfsAg5Yyq6RyRHUsM40kTle1nYwRyVVutpoZIz+FTeoPrwN4zBC/lR
Te4hoVSTItEwYOmhrlOYSapYazj6zAt2CYRpflWSRNxaI0cSBeFeztjWiMbHezC0
MqXZabIcTWwNiFVzyOxyjiIaLNO3q8aapCnk714H0CIU344H0rQrtcG2ImSs3fwI
fT2v7+hF/gj9OY81MHug9DregEcyAjKdx/zyvoqL8JYEz64GilXGKkfaNNnynnhX
GMfb/jfkaiOzbE3KNb0HtU5F1YzygzrJaL4dU1v/NYR0JdZm3CM9tozslJzJWhh4
yaZM6lQ/h+5YGCBoccTgGs9957wDEhTe40Er9FPNEZuxYe9Us+NcfQdUONR5Z9uF
83iTiCAwTcnn5ddqS0IPb+XB4g+00xXWv2ivwTTycskBpWhzUwvfimoxxPupFlnb
ibHsBZ5XhKoJiWTMgcwVxdYH6ddbcVkiTDeC0XFjbmDxhi3EXse2YXgMA+0g8yh5
ZR+TH476pHvh7EnuUQTz4k22AC3j21XaULJ1jcCWNPq5d8lj15MI7TN7gYycL7Vk
FI7Oq+kE1y4EWF3zz/wFNYvpA34frAMxI1Cx0AQca5a6zLJ7vPx99vOyA01ruQOb
KRY8JvNa+USyF9MT502PQuswpeW1o10A3l+2pnYtJr53dbxhrmTL+S1XtJWxOG6G
2pBrFy4FJtmxhz3LyVcB/q+oXYGzxkKtTxFZRvZK3gPPjyyJmeikaVeo82vmtKFN
l4onDD40e6n/XoEveZA5LJHkcMZ0xOs5P64pfCsqJ/86XXHwEQqbUT5khFB6aykk
C+K2f2WTsdhLoQKoWCSJocdutxUtH0yi7l7QkF0mSm+StaMX89YosiOos47fvSQL
jv7Lrl/VLj805LvbECrcs0h54bgyLlNSYhQSu2lc/2PeROOpphYGy0G4fRIubZF3
I/S62goOZ5aNgQIGqDJPHLgRh/1H3g2uQLP1sFgXdTru1KstEL7HepKoPd7AqUlv
/uXYeKOSThIEIA7y7QyVqd7XaIA45zkvrE9dzHTZcHj2DfGvQbZey5rYsge1xuIL
iSdtbs2lB/5UGGZTMit+ozwBsFhhtPMIPwCL25tkVsdwtg+/p9IOhZ0jrzvz9UCs
KgflpNfWqXbVsYHYg76zMpWda3PIlDfiiAXr1IiseYxtTwvoDN9PjX7NwzYohYqF
1pJoYZ9fRXUv41EYK6RNdv1zNr6TG2dIQwLzleM0TzivfbaG2Ddcr6plz3TB2y2D
X5TXiJn+FWQO2csoefUGETm0Izju8DBL40gu/JATNDJli32dhvpRnOfSYzQD+I6O
FcsDzLsBUq6OsuULV+TOf+0lbU1a5CLrVlNTDVGMyjEiyt+6gf07NVNI6Y8btMpd
CaCPYwPceyHxlpvHByIypOilmhrheTbt/DjYjvBVIVgAGWIX8B8x97ZmzxBdOANi
cKlusM2DxS5k9XGGapgNTsF2ssEaponuRZ9vAxTsyt7DLe5iSvT7f3jn/9XToclr
jjjZjQkHTan7hUmONaKtWH0YxqCavZTOltQOod9X7LmdjoNGZP/pckc+HccAJTSI
NNhnWf0/cR51emJUMlDd1z59ycNpsfqTWJqVkYeWeI9DiJ8s3Ftwq82CXvAlodiY
DNkPvEexxh53cvsr2ZCuC8bUwTBVi856Lr0CVPTwAEwHRGk41srpJgOVOkHmvX4b
N8jumcXRjyHky85Haofl97en93gr0hl/lH389Cjuf53NMKoAIBrYvEvwtSPTgWNv
AfU8Ao8t3y81bOXWStLMER83QvmKTMbL/YOyoIDiodSZ21yosKKCdJiLeaLKOKiZ
8O/6EDyGYBlSpDdJiGmSjtifRTO8SchmTmRayP5s+Ii7dSSV8zD0WadKx7V3CpxU
MjK8ZuEQj9OMYyVQo6yww4Ib45PTRmDTpyMZim+AqZomLSyq9yEoDE73Wh6bohg+
x108ks9bvB3BqnAbyavlCe2RgyYQ0vMcL8G67n9+rAfaAuLcioat5vGIN5qIYXNz
z0n9AEc1AeomU0OtQoq98DLPt9oHR3F5fLrMV4h/S6xoZqCmsvd+BnMT5h/xKT8J
fo5+RQAkrMxEG/OMYcGpfQttIzdx4TVWDBNlov53pfQDY3Tx7RJepoyfPiv1DQf6
Abgrim2SMp9l5+j2Rt1Zo1nqpvG7mvMq4XAbfFM3AwmVTSbcTsoE7c94IMhb9qVL
lrEj/qEH+pMxXgsqSZPU7gD7WsZMWEJKho5qzWk7pYqPaiBmMGNQ4U4VWipGJ/L4
f3TLc3KOaSLCxPbJigdL8u9qP8Lk/BK7/QZme/SL8avQdvIJlvhR4ai9g2rB0bnR
IxCB5BAbydNI41xLl1572FvWaivyY/8PdXtUKA6tpv6GiM579ZIBc7ARN+4SrjLs
4qGWN2Fx8eEMm4g24xZYfUqI+28nnmExMlSItKEqVfTDSHBd7bRplZvuUgnIFrz2
MnIJ4IQob8SOFKg2kuDfslG5L3hgwuzm86mvM7vSYftUgkYaDHbVztOzCWwhlllb
QAAaiJwdwvBi66JuoxNkM2NC4sCoBRwLrx4uCKAarJhX5TSL9h1a+mCmAD96afSW
z8du8w4jkerhVNQ1gM6PlcKsmRkit8Vmnut19Eo/J1xV08N2ZXGuKI1FldpoJ44v
BJyFDpiteLOiTB9Rp0SkTHxffqFCjmV/qo+GLuWuEP9PIa695W8uIdcqBXyihBfS
MoOZhHT6iehPjUetXRAVWuSnA/9EB1rd09rvM3ztodQfdb9ZxYY5K1xISx4zJ4AH
dnUv5PFPvHYnNKqQOAg0we1D7JzyvNSFjG93hseI3wfJ/bpY5hguA1BwjDYp3DdV
nvepfxCviuLW4F4cNmjYmwhTAPIFaRxkmPvaoripnpBIzMpkUfAWmGIAjFaHohPB
XxoWiBlMjUoQpNLdp8/u42vr6luKvCpa9YOX8fH0DsAZ4ZcwWXDRvnmlC5uErKoP
ybLTwXGJKc+KkmUNumbkTcihXHJsgbbUM98scUU5Qcb3Xnr+ToIRNIElR3wkujTl
ZKkwzvLujEewRfkPnPfnpZFEc5qrdNaYzXKQUumKxfww4+dzybrDAhNcngy4bDyb
zscjgo1kPdSyVGhfBUneCQX65M0AmhGJonm+B7Ul9Ag9bPfedkI5El6Ds/+RHSTF
p3FagaVKLHNK2D0ATSTMRcERnsXS7HqFtWPNpPipO2M9iqs3CYEpktYOuCjrNesT
D8KIGm8GvM9n2byGRCw++Kw1ts59/L41VuLeqkGBdGWm4BQxL22LslqZLkTJXz5U
oEFFrDrQ2ItONfUzW6oNx+w+GSmAJuiWZgL9+rEKZEqQAv/aoNzosDPvBBlo48sU
g6qjcAzSTRS8q5BHLx3zPTrHtr8C2X/aldlgK3sJMSNMX4TOmc8pesDLAKPUgXvb
Y++dEcpa1bcZS+r2wiJKWHH+MxIwlYthk7YvIJqaHqW8LAEg/5YmBjfyuAuSvyuG
bmz5xDsBzmxnCoTz1lODP+rxfdDVydIJyTN3ieKTr3q3BcnesQj+n56hcdTfQToq
v7O7hX4t1rlhlpKvW22yKwdgWuInSfz8ma1Ex6oNsFkzF4+wSDyXXLEhBKfqvxMh
GRXgLuVA8d7DT090K/f/gXEV+n4L8CWuq9WQyPB5BhbEm45Vzmilx9R9yaSY0SRn
0a2+ZwUV/EYK16bffrc/shwpWnd6ioiaLi5pVUlTGRtvjov+vGVQ/S6+RqZh8MiV
0fS7fDGlPotF1rExJhQaAtIzAJYsNoLIulLJzhibtefcxBuCDMF0ewaz28ubJ82v
l78bYXq8Ljl33IYvEpb6nTLMeLFq8cjTwKAb1N8/F0b9V6/BOGXIjJ3DsvHEe4Op
02BYQXIeYacOUhNaQgkpYuWjst4bBsFLwHJ/iFU1AA+Lg8QdjJnbve+jjQzawtul
quyGynj8xNmiVnsyPZ14NcLBwawrEjl2VqoZhsMQj8alej2jiJtyOLDus7RFCYJg
xuklywjXHRUj2D1qsPm1SToW26xIcCifbAmvHbcZXA5Y/pqS0v1vhOG9RWCP8wph
oEOVpeRe1lrX5Oy19k2Jz1cXFKBpJqwFGvTn7jjd982vWrWUvV/QrmEN0CpKYvbN
f3OiTyRezZT+Xi6fPo/pc//jILY+Vw0cO45X3Y7UsGzK9PiD9hHxOyHQ1yLpZrVR
w6lWM7Z1ynTTcXeVUVlnNXgaQOmxzqRu3x/5KPLto+snxE6aF0A67rIKPEvQjemW
sjUrNqlhxEUvKfPfYG0TgvGNkr+ePnxLgPoFB/oGLjAhB8hibxUyBwlNr3Jiwd9j
gwVxdwQMM07IEWrv5Pco3Lae5qQwOey37o7zyYPsUu8hEa3+YZW24796xoT+FjSk
jlP/ieHOE8tAtIIHKlv5ofx4saGpTlJ/W+NtdKNVl9Sa06/4nAfTEyTVyLfU1Wv5
iutofyEcV7QCJSDr+tEPgSkqmzcyB8KfZBYxEDBRB2sP9yj+eU+01UQjnCGiI8tk
okX+fiqheM2pp71YSitG+V6lHS6NivI2nI7B+UdvMUT00+muu1AeT9lBspmEmvwG
0BuNY6WEmdqihpzgomSZiPC+mnpx9VoTNBWvlwZQlRibSZiUNsrt6hOuaHNYsgz2
oDO9s94voIr4Kirl84Cr5fic/IPbO80Anpb5Ds5Atkxpf6gkRH+q6mP5uCk1/c8F
HQSrtpfLY22tsDwmzHS5rrl/4p6EzKZHb9xoWflf1b+ZjJpcUbBQTm//0xDRGtYq
nyoCqeXoAI7ygYJpPRLRXP7MJPmUn/+qbEJ8L8tky7bzE1toV+0qqsEDJ7ylfpuj
zMZXhtnKP4d6m6E5MmCfxf7lO/6l0giP+8uhv1ZcodE5HgIQtv6Lxk4noIfOrVDC
p4Zaa35T43s0kiAJm1abgUIhXnyE9DSJUXF+BA23b3eUywA7dOoIPpV+Bf4lghEK
V+qfQ7XGZkEkVo1gUOfQGfmobQuSokr9jx9BDVZUjaCH17qFgaQZXJfxznkBPG8H
QxW0jK27sPYTF9L/ZJVx9eqMEj8L6vfsgzPlAjg0D2HLG5z/Q8ujrVULi98HFLLG
udAe4RC6qf9+BmTeXLZGpqMQALmFU6qqIkuyobZOpG3CH8we/hpo3zrWXl5iciV8
hQkOml3d3dJp4YTMlJVrLEL4RQmsZiKNMqgffYgHLIurFWG28yrdq4dmKtIR6xNP
25+EHBaCfaOrxzqxpD4Jm+QwMVsHf4MfCJsT5+76Ojwx+zcJGQAGtCyus8/QaUsz
FI1fU4JGosKzPOat+6hEXaxTm505I5zXpWR5WrvogAdQDLAQvVuHNzJi7rxP1Wh9
ZGGJXAcO43WnR/mMt+5yMIO7BY33wpSlTJWhZJ7JPlZome1YQD7g7UFMAMNCwjFL
nOFWsODLwPK+YcDTg3+o9Tz0d81VMbOGHoOgQtszjh8sJyHAQetbmO8fJCyJu23R
crD83Wl0S9cs5/vDqLzLq8EKdz9HbTB68nkfku8cOQVdBP1AtfiKHqUbIT7YwWoI
b11j3aKTDaYwW9E4rUdhoXm3CLBAaS0GFjiECwcD5tcYYwe0iaBEtoSf5CiNn1Gv
B3VBzhefipV1kO7h5COlE70g41WdfH3Y5OotNImNQOCQvU4rtVXLwNJbCZbU/aDU
wQRfrCEglcd4yvjGlgW4mUH/tjaQcprzvkbLNZC5ywCMy+GGdJjAS7tj9r/nn+nr
yTYLeDWipJRo+FrqHGxtq/jZEU+274OF95ehqxAn2CaD55yt1MmMSOh9yXU0Zak+
eWPCAbY9A4baFpEUZHtXv2GDHrd5CZEimwvinCME8VAt9BCuwo9NLNx86csvvpGe
ycrPqMX76kXVwItQpAJts7cuDyj/lmzX83WuvV93EQQvzLYNSIPBoQoS0l3IRpIM
qg7pHFN5ud7aP998O2VAzH4HwFdVc6HVoqTCUXLanZwPuq2jCOJlwA2Yy5hNxMjz
xhEijNHqSACuUXZNZmoI60b+NmhwaEi5qagqs0itw0/e07z5u426QrwWW10nJ4uS
JKO5cK2F8mVTA2xTAldqgpYNYRqSxmzKOo3yJqrSQ3fCfcL6lMBydXjzxjv7k1wN
0c0XDVPrg9NB1zqHACvm4TUj8v5Xuiyprp9i9RLVzfUJfCzNrdHTkO/A/067xufh
P8SjoPxviHT2AqtGEMabKxN5qg9Wb27HfzL35oFY7PpLYgnH7caSWf45nxpqO23H
+/5/1awwDDeIXjsm5i5jiGdD1QiBLyHithQRYZ1uT9Y1pXLHkbEaNuFq37923JXR
jA9tls24L1iC6D2fTm6tnLxpkMczkRlsyz7E+RvIl2vtUuXjSb6e9rSDt6pK+HdW
V/APMYvNG5F3b3FSZIpLd1AcaOB0x5ZfBYtlPc8Ni33i55cbTF7ItRU/704UQGK6
C/2of3K9bH9SUhJW6HCC8LYH1nLEvOL9vJX27gELZd4es7Ab8ZoVRU/N93/iibv8
KFJlL4Ju3iZEKj3v3iZ6Ou/hFysLmjOX+8DRTHKQJkcFIBLi/ozKedcquAhVN4pz
f88s8IzRDbhMLJycsd+Jhzv5/ZKhMAf+pFuCBP75B3ED2JrKlhLl5Csr41EqKzsB
BpYExwMGmKw6AqAJlqZT2czPXpCg71N3u7HrU6Y0Z4PHJaYsC456/PnHlC15UX6v
zOI+ObQUBk4XsrKix3vT8n/LdwgV09YNot8J9/IJMsqByJvo8nWfUGFrkEYV+rcO
VD7NkrTM9VaP0FmrdhbGz+8ODheuGeqGjFzo4KsBBW2oh4wEuQIq6iCaTSQWk+0n
Vdhrw76/OPNb7kl5ARoDmrD1sS1o6aU/TojNrTbT+JUUTzkt+3RYg4GRd0Ft+Nmc
9Ko60v8a9f/uf57ySapoKTqqDMV36zdtT0j7wzDqtO0vQh3h3UG6bNKo0MlnYvVu
qRujIli3Joy4Z54bz5gsxILmZSuYaZb1bCkYkivpA7zFxy6WoGG0BHwwuE3kVgbb
u6oF4uMDCw51hitJwEC+3WLAye3reM432XfDObEwVHw7wcjWMil9KGR2TL79Sw1l
IoaK+Y6F+393jeDziKeAoMjeSRFkna5EtLr/NAjTHc30H7exies92Z7vvJdWRVvx
87evRMxd9IY7YfV95Ua0RTzirZFgtBcHWS3LEXAeKA0KkVBK4CVQCYwOd7yacZQV
Rr+C4ojnIc+NEtHmDkg3HM24iW0hGW8GN179DR/2/ZAVPh6bpme6soIWCyFuH2Mi
eCdB6YkucI/rAV3mJBYe+wjTF+V+SVGpigCWxRDbEo1AO97gwA+NicafJkt60JAG
Zw63UGCl3RK4Pe9wqk2y5sabXvq0CsPeTaL0ZDnDQXBjhA6z2VPFfVswX/yhoul2
pS+a7ZD8OHN13LczfocIWmWhdMZwwxJAQykm91IJoxTVzbrFb9Av3aXiM2sbHEbN
u7O8OXJXFtKhZ0k8TTHqO7SSu7bK2IBLLvbwMDfpgCM5TP6RysG99wwmWzdjnBWl
pJ19b8u5/2JVeSJLBOKuJzRGFjJ2SIyPMHq01Es8wr/8CNSleZjZZ4zyslx8VCOT
P8I1UVO5bcOYLSjcd4nN5aDmsKViEagKcWEvnd36fNERg8akAdfnLWrGWqnWEqlD
OwV89+BibJLsQlzpu8UwupsUG7R71y7XeL4Rxe3sdgPc3mPC+ejhq44RayWVVCaS
FBU/y1IvTSICx8N3Dcpk4myWEboAtN0FodPA74AYdSTwEtnhH8WYE6QJLFX8Kal5
CSr+HQN5r3VmTnlgrmmaV6T1U8ImL8Vz0N24wFalpydsxGVznt1zNcvhLVr51buE
ANZKT4D1KVXgMiwKXLKK40kWczZVGyGBKzYinZSMz2YOCejxH5n41gtzVEaWuvtf
g1V4nhn1HftWQu75iFPu01rfPTSqBvQa2g4PH2NGi/dosCRju6CkKqa5DEbXUWZF
SrUIyISnQdtxYZ6U7Cgf21tn9kAl7u30O1LoNzF2Yy6/FbTtDuDttM6zVSEvLAhL
N+xB1FkQH4UT7sWG7Saby3g62EWTaYdvfC75WLd8/3ofDmC4s33B+5XE1gkd9sMR
4uuXvaO01LkyGDC4+3NpU8qpyv0nwyX6bhswVb1T2Y/WednoiPi0B9ITFUqaJdNt
aZpRM+DJGj3+Jj01f1e4WfbkaA/ubKihQKaGaERMa0IVmBp2AKuyT5yO7Bg/viiu
iNj+2C862R0wR2gJRo2UeP6WnliF20drnFwh+U2m2KA+wEdPmMofLQF1Zrp9RoI3
U4FA3JKdOkzWFzeh27Q6/pyY3vnTOORESXSqSrtXy9NqVRkLh2IBPxd6OoA8zL8l
zP9koZV0WVfMvws+2ZwLX9Gbwbd18e6/r1VIYS+qykZiOru8dqyhGmufwAppFgNS
BIPzpKYfHEZznDFky2/xiJd/FlwU9C8/vbJkipdxp3ETdE8N+ouiJkoCgPOHvF7y
Yzm17m0OZKzFZDYswsGU3Q+Q9yv1Hn1LcE3Kqt3nGTK+hxxqjqmYl3Vj4GOINl7V
BifMKZN8sIiKp2dIJvVBCkvMEB5wQI3qWBqD3cpn35UFIrfGrNas4pWjsW9zJGnI
X5PUx4w5Ln5Mqi+g+m2bbL2BTIDQQhe93UnkknTeTwuatKxjsN70GPOvAVFoj1gb
MBju2b19a4G1G4vfUNh+tAZCULnEvdvGPeykyYnDauUh2mcXXuv+l20Uw78vSFNS
tZV2KbIYRjjBoA+WbtogUdYIadVg12rzda0gIc8E1FtMm7r6qf5aTu43bo5J343x
tw1s4iKHiSptc5YtiH6MznhbvxaugpHQAs7TWqDFnTs9uBJ4zD1Ue9JvZCtO76fX
so7m2wsgIhad+PBl4l873BUXwzKMdTPEomgiwjJNL8f4x8BphmljCfT93IwsRR26
/DO6legzbOAuN3gL/8VrtQM/XuM+sC9Ffu1Zk5JxygePFtTZnYO2T6dr7SHIuBe8
Tl/frJSYAs8sbSu++4TO80LLzpmt2ppfr+/gsNwaqsO5JQWBApahvglWL3/33ulH
nIUr4FEk9cDRgZEumoD+OSKUf+IqvaS888OADhhy/X1gOgSIhxJix1s04EQRGnmf
uueBfduOBGH+tDkAPFtlB+mXrthAP2tY9I9sMUgxKZbsPXkR6C0Bei2knJwPD6E9
HRd0+X1mfaIlb8bb5R29AuqS57lXpkcXpgg1SYT6mjFN529uwXAYjGyTXGyRuwlx
HYn+h6tX5lQK7ZQy7NvHGcsR6glgGjv9xGI0yz0jVf7boQNO7EmyK61MTXtzHHDe
r87ZFFHpgkWojhhst7MNOanFUxRviNJbonByMbivesVS4H/aELt+YnjUtpnnZYS9
kkrOmQh0NYUsSp+hglAvR42Bevbur4lhOcrjLuI/FoT27CrN7tM90jiXUrBJ9Eqj
9PMlJXW6G8xTBF0oJRZ4TjQYn1Q55lRYK8sb672/ZyfwEQippp3x0N2SrqRlkv4q
AaMzJEngto6w0BUrvKF9Vnxk5EX0mhM50CPrmLL5Q/xINMSGOlx6d8n08QE07Kam
MMDR86olfoLrz3f6IFOvC0Jwc+K6/ceNr/xVGsNoaeCL3P1xc5RKDP9vPNjy2ff/
h3NSSeowJAvhXZE1DgA/jBqKmg76yx8VVDSFTh0hsYMn1YZzg8MEw1QT+L7wiSUj
O1DOACDuh/Vc6vjS7xxu2m++W5tH2htJUf/llnpDELGMvHN7ZcVhC0ZnlgaRC3R+
LJl1O8I4fpzgm8+dv4ZhK9cYaAYJpDp3I8T7zX90iMa+saX1MnRKRiXhd6gyExHB
KN1irbmZ+xlVOIXWv2NJdUYV1Imm4xXJ2rqtKCa8hTC0TeOXjQY7cMhe1T24iGHj
Iuf6rDnKm4HaflRmLauMsPD2cnUPR81ScHaNNsbb2tj67qrdBrTAKCzwspOdudnf
3JQ2Tt3uc8ir84SkVu9r+NE9HjHM5HJHWt4X9TNVIEP+6JT582X8J+Sjxky+rkx5
KEVNxoC5OpPlOftwo+j+v6wARxvYkPUShjmvY1tb7MbwRgvt9BR/36+GjeuC0r+V
q8DzyV0mv65QVrJSzOBZAfspTeeXX/NywsxoLrBtResiytUn/X3itPadGKfGJhGu
ahbJh+pk+wa/Q4JB/s/1FqdPjc3oAsOSgr7ROfzx76vvDpSuGNV9MBdBq6DFFTyu
PR22CQIF5v79PsdNz4HYbRaojdK4dqHU16TgPL40KsIcFlKmMMMTg3Z041KkhJtU
8mCVeJROyGTf+3h/FBEFyISBb+/JhmRTG+eGP2miPJj8sJRHBqGldi1aYwceionS
vLoX5jLLMDf0MxaS/JUfNreaWhdEKbTxNDaRgm2D/sT94QtzChcmbg6grno+FsxG
SzFOf5Bv7ygDxGjezpKfPX+ZkVW7iCh+1+lCfd+ath9+CpTNjkdXw+UWCtHanneB
5owsgr3I6RSQ1mEG+LSClbFjLhnssWU0iJj0c9G106NbM6mi1pEhvO9Sg8cXHsD6
sMTlBGrHHVp99TYEA3u00lbNv/AjYSP5MImeFN/cx6rzakt7dFNxeMRv0R7qFDDw
4zJz6C0Ao/T3h0NyB7TYIDuLUAV1+E7D0ue3wU3plkzK3QgqU5bHNrucJd/C2GOx
rVlu5TzPB/1xt+yUaXL7S4ZJi12mg5VuRguDyb2dcUGNvHGC8xXEbc20pKFTWXhB
JlU+qAwLjLVmbrXyJdEC1n9QWIx12BhmhxgKWXGa9uF9aefppLsZXthnFnzJ8xxq
wGl6zGvh73QRBnUye0UFbyNqj9mPR2/v4oc0C8Q2m+LrHk3XquQxAfW+aFAGwc3+
3tm6xxnepZuyRdkXTKdHOOwQDVtTBU6XAJDwMpuW3cZt+5VNeHyWpIQn0ULtt1vH
O1J69M7VJyHQvpQlxTqsXnhQX1jE4CzVVnfcicDnIIgBli+ALq7kDLvg7THb/K2A
uv1/5TKMt9hnn2u5hu9BmEKCSebsPPEu3VjrFO8rfc8PbJ2L7b/KluAsYqlHkajK
cgyB4JmPFbqFqStRRx3O3oq2p+6XsDmp7F4oMu9lw0xLeNMIQE1FzTji9uTvPQdf
z4IlXMtujgyqYFSKV6IbwuhmxIo/QpewTzczolQa5eJ10DPhKN2fm7/mnFkep3ec
NulsAox8xMkklmQgu6+iq1o0DaAoOwuJErF8S8RqUUytnQeqN4un5wWj+xQt7wyH
IL/I3giINutG006Oy3byB3FCB2fbQ3+HVnUDAFttBAkGDo1SBS+5xq3xGiK12dlA
gpFoGUowZwSwbvgzwR/0uXvLawy89LdRVOVPnT6Rt0qoYdYIqczMJIR4wL1GmXu0
jS4YdYts5FwkyXQLf9SHxx2WBBB1st2L2ZjiN40dkqzlU7dNiYPvmKCDhPIuuSq1
7VuecKA8Tkl1SCdQQrw3WSdql0rIP95Z4rkd4eMdCMWwQC6OGvDUhduTa3AFgoWm
a4YRZG1PgpFvPUI06NofUQroeYr+Bdu9ybKZGCAHQQf2BxbX12zj+UI81+QE/i/a
y7RlXINWsjv6uE2BrlCsaBgRPxGq6uoFFcJD7x+x5uJtJg7ENchuAK/hEuc3UDYu
5wkvJ2qhyg2yWJSjAHQlMNjSVOOxACzY4whEvWoNYUjEhKOTU4zO5DE05ia2LbuH
ZHR7Btb7WjX+Dk0sxPf+ACrT/TuNZnWtRp5+dTIAFF1qEkG6D0zgkNC6QJtEvbkb
4E09/ms2p2kaafINPzHlGvTHJJrvBncCcFnas671mE2lsLGSJDUrCj11pylFvqMO
p7VoVNKw/ZI63Z/7B0Bd1jU28M+wbFa3QvGu0eeBMlmDJNrN5ezbClvYWHG8+zuq
lEd2KYsSI1pGEA5z66BkoKVO3PR53oys6+q40+maMaYNBw0263O1SA4IJrOO1UNG
7Q3uD0pd26KcZiFR63SO38RszpKc2Anu2RvxOhMTEY3rhrnmUrGEw/6lhB+tL9Nb
AR1AOqVYOQEdMUB6x1Em4YXlEERtLuT2PvRLIMwttBtUJRiT5XdIfcEptjUMcRLr
6nYCAnU9PwQ+n2jA2xWd/rG/aj7AaRwL80SseqWB3N0umKTjbwoQCDkuVkDf3kAR
Airs89Leo1hPOP60LawkIed7kTAhwgBFZhoNoy+vGKMcYZqEECitxdpKhYBzDjym
jO0fC0AC+R+C7Dnn8e+Nb3fjkGKAY/z4SeRId2vAe+CmTKj9HFZsATh+63r33hEZ
NiSj/cPTVyVGM3ch+lx4DM8sijb7AJ+Wqi4cDkVnk6X9i1vX2z5WJ7GwKqnXucCt
+5WMrafafScLj75YqtdCfw/FT8znmVYVT57fVo6rWjlqoNeI/jIbuYz9XCfCA/bU
9ZrFaMdw+RKxCOHCIo5zCmMsBibd6Qyo/ILCFmGYL/hNi2NJc5URNSlsSbaHhQE4
pBZrcSonYtJSSvXxl29kZbGgvcyzD/qGTXBIKMRwgpGGT4EtmKx0wcmJ40rWXuhc
PtlR7BH81SsJU4plnU31kZz5tPLxU/KvjpNYtoeXPpR0M2uEKy0sWobv1uHFZgyt
OucPlm3ab0t5jSgZYvq1nE7T3Q1vMufZhv2Hcv0+M+mytk2clUsMfQckmZV7S/bf
ddITQCXAhDUoqdhOLCuBXp2pfux5+kml54hrHuk2vcHcz91OU6Tk6oVia8dnFCtD
4ke6UwUrYkMimMLa1wx1AoAk+K+p14sTb0qfFkDRhCwGsfzZ9/5hgUkk6AGsJDa4
7fZZe/PXjzHrBRYnKTkcsSyMmnrmGz3olK3YZDgWSbOB0jt+jBJIIyRzMg5/He2h
i5elHW2L3shP1yiKuE0N5ELLQIb4lokMgdBX8NRoML6vwst9UujE4Tw1CAAOpcNj
nDDK5XbqibXqwnIlwcHpU8bchmqEpodNFefgUR5sU6SB4Ua4EJsTdARL6+VmvnIA
l4E0lnP4v5LRyUyiYaBvoxJ09hXeNMD52YvhwZPifIUWJhCsZrD8bK+uKraRalC+
xKTi458kchSBsDPvJLnFbwQuWlessTtp+HPyA7+D2t6v92bnwoDZq/t7q/mag3Yj
DNqtDQD/JJ2kBLVqM9v2tWPQKp1KerIF6dBg1u9vUgj62/mr/onoFr8cqTtZdZoj
xOdzXMQT2DZQjkjj39927qF4ypxTbDpwy79YlXLGTq8/pu5loa0db4H6CEKCV0a6
k6ijGKoBsgjElDMtfl3iaGRf59miIZRdMOlRbZ4Fr35+6useS5P9YZW8FNUJRM63
wwK/Uv8xARKm4Vv6Mad08jgoy9fAc+8oIyC68OZ4qmyUhrIulvMD9+Kb6yBJn+fV
ZwyUBKw0YOikUU4V62UQmJrDF598s1jfAC3+VL+rls/dGuXWTwvja0L5V3zs+RAU
r+BQ+UDxCAJssqGTijfnq5lgS0g0vZ5+7Myl3hKF7vroAByUBDACWSLpE6lHjj3L
WuX2uQbQffiT9dx6vN6/UdJwHeohfgx9I8h7eJPVLIspx32yjYLZsScEHe6VrCRN
SFARH2PQJ6FhL0N3FL8DL9OfwQX4hWXY4ueFDbXkJFlIvZJST5+UhfjRozhwiorP
8jBwruG1VCqDq/QW2wkEDnFeYRtms7ZqHGuxLWCV8KG6CM+LMB7woKnL0+jIiIU7
WpSp9kenIYJfzvtvNd2AsBdHsbPCJJcR/oG1eLitbVsOYZKOqrQXtROJ4WTqKaJB
GPfKzDGY3jNjPU6W8Lkl5CNUI0yitkjn291HWeivCpxgdAsP5/qndbM0UYlXmCc/
PPJpGsgrnefeUBFl+NTrs64GFfV3dXQwUOPSY9Jp498Tnpi/IpIFFB7x4OPy3Hds
xLS8B7j+8WszREt/3tfxqyhhmB6TpBCCzy7G5A2xfhX/IV+BPaq/ibvKDGrbhXVV
VtPKasTrN0zcGTj10pA8eRv0wXUf3m344yr++CCT9PpqrkCX7v0rFGyAOsCDWLBc
OIpvZjRSIrxUbxA2AZF5IRpJOe68/vll8mNdMcPlQn8R4kbO3okCYqx6190nOXm1
P6VmBTxaSvPzN/6A0FbnhRQ6sHehFbs++36R95W1zQksw33uIJgYh4w5OTCdKjLn
2+6aXjqDAjrf/tElEn/LxDeYJVU+vMa2aQRp+viBhVNZPN0TMDTUfuPw5e+u6wAm
oqtsAYC2QDwqNZaBUUqa6r7PXrTjybXuh/A9/NEP8cv71umOYYdYYvvooGJI3CC0
GW2QdQG5xIQIMBDeaP5eO2m7R9abn9ZZyxfrWfeHkMpsE2xVSjQMO+bmcYjzER8h
8UzNGWvUvdhF8T+zjMcsumeim65QvPEkLSHRfWHSmy8+4IRocb2yN86mmmISZD+r
vzvJvZRz0ZzDHH/St3Zn16U0CULpLM1vo+58mRIg/3CiqcjKEgDv/nvSeomHCK/L
gBaFlpf2mVTXiMydFuzJhknpdl8dnoDx/UK7LQHRK+6T8mTN/CvOk+8KkM/2quOP
M4mxB8fzQrS3kdEh8m77ywMMZzt/GOr3NVzrj0ZLi1QNHYyqn5wdc6vOyYIvh/cR
KrhoUBQtev80l/D6wPaasGTeOLuHDM3rYQVhan0z+nlo4y/u+mDRXLSG9zEgzLtW
z28YB/d26NulZj00QXmsxhY8tNHRN/dza24DskNK3n6kHM0nlVzbJpkI0i0H6wxS
RidxI6Phcdr+PNIVJMJ67qsLYBc2NGJWmRd2WEvSs0utQu/jTMUGuF2/m4LUvs1J
SQyDfKLTcxMz2tddABRgOpPrrjFr1+XZEk85UhDf5/MjDjt1Kliol02ZFynR8ge0
Bbj8nnrKP/2HirI1kYXYpGb+a7uMFSjnrFsOZgR+exk45/eNytUgcoupw5tywwKq
i4HtxkBzTL7l7r1XjbusC1ochcPHNInynLW8uuuo5QymruLiB8ePEsYM1EL47aaS
UIX9fvnmEoPEa3nFaGUn5w+Ac0iECJ6l4nvo+2s/+vwifU6u652OyD7QIgF5S7Au
20vRxyn4c6u9YX2czurawIAOqQh7pvZiq8JIRqMB8UbO8OoUlNajf0aQy0HBypPp
EEs9/tr+IRqgltUX4snYE6B3Okk8rYqgbZrh307TNc8cMmG/tWxv8k29KqRSiBsa
4vllFwI7d5tdLpceOGc88pmZ9xxmCR+RH9i3QS/ZdXdNAe/Gbpczv2LXuBrrBRT9
iBCd1gQ20fRbqLuY78quxPv2QNe1wQPFWgFLT59hkrckiJzAffsTAsdRkOS8ONAu
llOWbgxqQwJ6tXTsVr8+P1Xewk7yZJta0Uu2Aj6bJZuGRDsyjHfySQtVt38SFa9+
IGI+x++2Vc/6+313qH93QxaZkrF0zfdnIa9MSToQodzYhNoUy1MLSv4mZmFrHdn1
XjCoSS5ObMQ9MI8G4xT2FSL4qmOkf+awbI7jMrluU4rFB4ZLPwLzLOgEEhDBGnd1
ZLX2UzO6zuX9l6JHT+D3mBaF44DQPW0QrQqwEl0sEJqnx3wf4YxTg7KASebaxPIT
sHdoFeaOHmEndPOQw9ph2JnYQf9dv1ZHbwg1p6a0pdsnog7XtvG168tSSSocfNZK
/6a9VHfuHkt/EHn9hkfJLQ1jAv4LM5w28D5pJeBy63yHYlJYFtcyvsFrL9sZZvRR
9lgFnzBVZ0hVvfKI8JcQqHloFqYKO/S4YDA1GDL00XUaM/0kiW2Hso88RrugEFOu
BjwG6QHKRj2yt8vsx8kBl6rYNiZ4jguTFqeuY6/hiSzPpIDV6nDWLrEBuo2BvI6r
XSbqyj4BrtZdpi5yFWSkoCZSDss6ZUminMmGq3Xh91HSgeGlaGTyo6T7C4uFTCXI
8qe2ZrclrXJFBuWxar6R6lwUv6g5g+476S88Yhbk4Wrn8nILn4ap/MTLi/TZSgal
SMY/CqT9e2ZvknAA3EuAhN5tbyf2aWNUZWgMDqUiFWE2mlw2MCre6TKyaBQs0dI2
lYQ+ioPMAcrU9pggXtxvAF19DBSPphRWYuUkI83CXnr1qLMSi6oxE3XDLCwdZnmW
xpnThZhYcboYyWdB8FQxhI2R1dsjOMIdopSECSDXspADbBXJUq1xOSiSwHEBLqpa
7OHlxCCqHlnG8mf7Py35oRd54Cjh/dHG6ET2Rx8EksiVS7jgFLghYLxN5g2ETXf9
JLfAJr9OenX+duB72TJCg5DMyiIBtPTe/6FcYlujMU0nhH+3y6qqaODoIEomnre2
cGiCf4FAu3SGd9OuVlwWqCRfBwnC2VM6/o7l9pvwv/T7Xk3q0wPNtkX6qlhjQn18
KeYX8f8FDlWcRRYBcd/Nqdo52232Q+fcrFErtHI5gY7xj+CDml8CQTJ5df296dW2
gcP0lbkRtGnIfzdoJF7tpfIjm2+1h9zPjkF8XdUXflknhUATlVtJsipQw3ArJcu7
wM5wNEGu45VThFy6i9ZqnQ90Sta2DU2lfcRXibrmdq53lfFBG8f/7qEqJJ3fvUla
qyCynKoTMIHQAxFfmMx29xD3E007hIEIJoqxySCV3eJekSPA1XTTQT1lMBMQJrBc
iYPkQoEEZON0973/G4jGQ6/VbBp/mmPUbRRl4s9gzPGR4TQAMHGITPaVxpI9ubbG
CcYEaYbDlpDl6d17L3duBj+QveBzC/IGNUDMc+2g0k5xKaTk0+EhJ+MYJ+XNLDjV
BApDkwR8snQd1ZI0ew3FLuVxL3lj4HtV9aFHvta1XYY2d3vBpTRoMEkB8FCosk82
mj7JbzpxZOolc9rkYLEAd5cv6/lc9h/VZ4Hb6u80ytEhGSG0PjmKVAHpq7qL5P4G
wIGvjOIX4hYqF29eXlPgWEmQ7Wl9Wa4VE4+jMfJazJtwhzi9WWzIfJORVLN2Vi5Y
brlv8SWPXa0UH88fKbB5AACSGEDjwP1DU7axBpbuFGwvTJfKxVGimTka0trre+Ue
vvcfN3jtohdsCNVsJmlJ9YNbI/lAnGosk/BqkY+hs8lHcxiyuY9nvDe7x4bRkDIA
bQ/ng9y84WAkyOZ8tTxyw2RlOZPabOkPpIIdyYSHw8Xzo2XSlGpVXF8e6bPBVhKf
AfJ1FRK950FeF5f4ElIi1pQesr3V9v1kQg+VeDSFw6fG1czRI+PpvIuz9pHZOMXC
3YR4n/vpBxF+lshMZi/yz55jEHRl8xMC0DxReGZt0eHiq3/o+7cRh2jjgW7cm1ol
nd6qEfUX7sZGup5ajs35t+yjE8EosZqfQciSVqe5Tn2MZx47sTT+aYIxyU4ec5c6
JAHZCdz2luRiHpQ68cRZneag0RLYUHm6J2VFmuyAGkYgBblvLUlTEFWtB4sqR3BW
OMkLvytqrTm23w3AX9WXiBwAQlFCfwPrMmDw6bd56CJxI/VAhYD/FcRLhaFyYKPG
WvrrptcE6Xt+3GP83QkGBNJuUyqjUp9hWIxuSbdUpdholzcFklPrRPsFQp9CFhV4
bA/zXKX9PJt3rlI4/O8+FAAfncRg9jnwYEZXWvEiZ8Hj65IPdA25HZBKVCDr3qul
Ph5TsBcBEPbjWpaLb+eL6MOSUBDmK0SezpakhAsrF0aHuD/v1pNxuff2vVrAq3OS
/+yqhv0nG2kb9H4NbJPlTo5rZ6RIFNGQIjWwtmk/wA7CuLAbkw63iaala8PSg5FM
qkfLHQALA2m7KcAlY3xuXbBcg9TVHUZS0BuRseUI3mS/IgMYnG6f3AOFCQdtbW5Z
f2L0VLCGNSlWXXWJKPg2whU4e1MimqZ3uGKFukDKKPwSOMCljD50KPtiFOxNmcaU
/7hxycWyqB6HzvbhcpJcubouY1t+pcVVHD4aIEM8MjhF+09popBfnkeBan4/Y9LQ
R1luCTf0QkGoPPt6TGqI8Xts6B0CkppEmCiOAwYHWMAT7lGDKq+96DAVdfJP/tQ4
eHGZiJwUrlOzUz8nuQaIIc/mFZr5eF3R8m6UywU9Sl+nntKcPGpCq1fGkWcJT4rs
K1oYYT/VAKxLSGyz0M9bDseU2bgGfVHNFWfTMnbKS0y1hJGLCyp2I7w9qZpDONCA
FmmLe7FwIdiTdNRaKO8Sq8JrPjSLh/9250DEGNMKwrX18HHcxkLuUftgyYk9Ci9H
D+kDd5QGfQB38i36qRp0HQqQ5+EH7sywNDoKx3v5mmvofo/f1Brc9CaM8ZaZ6Vr0
dSC4mbdZzul+VZGIb8AOzObIbRW6U9zjjb8FFt36BlQOQIGXXctAojuH+FE1SvuS
hKI4FerO165kZPa3mAWaeymSn/QTx3MlY4MwYymgs7MTsMse04nJri9uUWYpyvQ+
IHw3L7u1mPibyRz5z9izAVcQ8W5Tl49fQ79U63rizlYhykrk9VMCltp3lvFhQoK8
9u0qR/HO5cWNnvxu7pWs7y08isgg40cU9xSL+TEOKMFaj4UdP75jNIDEKY0N3YtE
0tVqVTkxV0bsytkdVjU5wsxF6eHXe7PI+8SXvmYUT7HsWFjZNFhjOdr95sh0EGvt
45bFf7xd2Bk6qY0vMX/1xOfklujn3uiMh8+QiCmZIHKvvl/sbwYMdrdsTu9twq7y
dOadccRp8gA8GeKmimKmYkv4D+3DDvlW23hoGo1cTg7U6A3/3cL8y3/2T1uPd0XB
2XUKNIm8qBdIz8Lk+XC8ybgN5HLy9qYLtuppmZzF49jdOFr5iqd6RqqlPdGzgc0k
cFhyCrhc5x7tpgUis9gizegrswryBOLALEdCIcwfOQIM6cLEIbLf1EU/lGN9F7lz
I94nhelSGTBhmgkCPZ0SKZZ5Pr1jjedS9efFq0axCvvkouASe9UenzYButb70WqM
/WMlMLonQnlk0nrbL6TNJo0zHgKry2u8n03aYSCvp4z7MoqLIL+teFbA9Di6LmK+
G2OvOmeAGqEh992+jKgLnc53ap5IQZ+77PA+JnAP83PkWhlfYbt1aenlDDuP06jk
ju+l3hZdUa7HeiaJyAhl0fIEFwy4s7zZRxeOc4boEhnLpM9jpBXpL4D6KHTvXIRI
dOev5AHJlkPVTCHujt9RWJ784z0ZpbMHcStddVVPTl/XSVqFL1MnE+RV4VUeEGKf
U1Wu6yUQZ8Acd7yV/iq0SwuItYvGflQjWoFIZqP4OlzH7eIcecCHsJ6SgJ7vB/5s
gmebGGZVeoe6h0MIEfYyzMCEr5twiOw+IxOl3xfAp9x1tYjDlBM4becA7106E+li
V+ljP9erVEkUeK+cQ3Vc9X37UQH+rRiYbc/C5CTLkj4H9CVZho/TZSOj21jyrqPD
vZYl0Nm/kcGBYPf0cQ4HtM03irKKrykh2okp/jiLEgJ6cwZVPiujF9ltM1Do+gmu
KTaJblIOxWRjq0affkv6S0XLD1PKEKdDUHqjWjTp1ZAsJeOJzGVtrp4zKwEXleW3
kKuVJKY8NPRyA+1Yb0J9j10S7oqciMzjBLKOdm1lrNNYB7b6Gf4KZ1Ovm6TPhZeY
9IQR9nJ3TJtk12X8cB9Jl7ex9nTErk98eZNst5OL0XmK6mMfZ1S516hsWZCQ5VGe
4NuF3P11t9dMgw4sAmioyAKh+Sk/Agy/q7yphXT3BwXDdSnd9RK+sfoB56yw2E8X
SkGoNuS3PyNhmWopm1I0vZyTGSd4syGeuJ36PG5Ffm3WcnXqxTTManXfAyibV26H
eYLA1y7I5+Vn/+fpSYLCjjQ58NBiPFOoeN9H7ZuOtWljFOvW9pQBGRie8y41kw59
s13THQDf+aIWEqpygLxpJAZXMJoV4JuokG3VACQP9rf1LnP37hAe8aVIEAsWBNvg
N6YTG29LM0EJl4VbsIjq0N8O9KVXVljA5dBt0eFN+mzjTm2HiaYgWokgyYXCeXTZ
czHiDtfeub565NyskAW0zOazUirmWcIO5mA2+/aNeIRIyYAkXHhDCk7gIrqjW5pF
QI4GsfT9uld1onF61uVhehfIQuW8im4KDeHHjNPWezz3SMAWW30LWoD7vAluXzc2
nSTj89K6Y3JRcjJGh5QRZc5wl1LOGWyT4LcpWXtMIZiVmyDWRMfWn13Xk+oJ8waS
qO5oMYe1mP1nq+6zPLUn6b1yWTJbwrsyIuM5EsGPqsfG0ZZSwExfnNAtsznJY68T
ujD7f0YDa+THFSGvMs2Gyf3G3HHyMsB7OpqwkQ2ZGefKsrR2AAYcMPrlB3eLCxOb
PfZ3NKphi8DOfqdKKfbtPbV829dnHFBVc97yUcrEga9p8EilWmqmxldjmsukvUkx
Gt5nzAJ/khiN1zTqAiY9PHfqZY2LN3730Y3Weqoto7xpBLEg/q40DRXq0yYawVt1
hXYIM7F3deG038WQgnOxGofhg8mnYECQHbompThE8n9WSycKAV14HUtxxgIRKFmn
6WXM/Xh/dQDnECa1JMLY3NTDd/ADRPZHEsJWs7q+Dvcmpf3JsDnEXyiTCVdD9t4N
3gb6NK63b2nrWAVl69zsp//YoMiiVWqLW13efmUrUM9hEHaVPfIlaRi3bcx7n7f/
4mKARYp/5zlS/ykat8YRrAKAUaKkvSp/NtHWSnYY6cx/rGzuv5RV7WZ+K7EticMD
eyFsA02f2nfc+Nh1aosRKQAJOkkBv6T8MkK4/0FGZf4Ebcs2VQc9oLNMV6o8VO5Z
TRutmH8tbqUtVHfxukFgIrjxf1iaqdAmGA6GQPqYJstnpHOcsrphGnfXqqclKwne
XRNdCRLQAHVmK0hWDpfJoXasQx1OJCHB0k5rVospBkhR4PmxsO/5NLPz2p4g5lVx
NV44EriVtBCiDM+i9/8ND09fswoaBXjgGEbyVgDWM6P5hNMRdOf51fNwHfpR8vF6
3TKe8wjAhMQw0IVQpxdEsjOnTrVl6wOOOf0CxtqTFxtBg8mPZFDcx35IBZJ3f0BV
To7E+qEdmZBn56CrAMf2Blrf4M+Y3AcdTfDrom1yHf0WjMQrcVd5YY72JyCzWO5V
gFKPzFkIUq2kdtXKwSgYlsj0Qs42Nu8oEsXEKsIJ8uNbZdjWq5infTE7KApG1Pvd
S1uRRi1Wez9pRgNEGtVjt9XgVu4fZyAyhA2g7kTDqcQ1QPaAdw6YD3q90YNkvDoX
eNMBh7Xij8BSNfu3knM3zSDk1vnDEr+uRSi1Zq26Yz15FekM9O7kwKssAA7mDkrF
olh7itV8gymd1I7gNdnQYHBWHtpX7UmGoMYcMdza/OIvcdF3bw8y8/fzkNdG+a24
ZORZn72GnOWIwUAyZA8aF/5gYkNxt/mQf/zrVJvjNccaAq9cYkhDLvKa105HIG0J
hP0C+e70Zh4R62sRtlgsmyu26Pr4aztANQQTX0G6FqVLc3gmfIqIkDMXjHf6uiZT
YNVgVezyYdK4vokABxOzsKTifCUt/+i70FPDKEnJ/bgwbInDwSWCNMzR0bNjBNkp
t6Nc3NiwquW99EjG29ZbK3Sc4TbUBXUvRhI9T5ZpqAuW9gBTjGEDEZg2ya/RjVGH
yw2hjluMU+mn3jd3JpQ8xxqP73WULjwLLYoh27NAsaufLVSV8ggYd9L1hkFsTK9y
Pl9urPGbQHMVAr2R7IYRY/EIkF0tcuUmVliyT5Gt4x3ch9TUM+iQei0hwh1A2BDt
xzkAHdsQdNoHmxgVWb0dNQQHY9mf9aKPGC6ZYJS2GfG2BFHfbM9q+U7JEnktqV0X
t/MlNFfa8Q+oRHcSWusmI7aQyXliDpCWPm35n/7iJu+AzKyDViVlCuKwSaUKhFyq
+aW2IN0tdBp/oIJM/inAxjT/XaboIb8yiPoM8/gH61y58Si+ngr2RCPSU3326Wsd
u+SJHOoE0du+2SHh6PJv+TiG50fxKc5oDhPC1YlsRf+GCmsDM41SeaYuwVxuaXnz
Ot1m2ZrG8DG1zxxDB0F7xSvpDN3be9iRyFBi1cfS0L/AfPj3FHTeLPXn2Xr/jEb3
7ASPDneeV98y6CjrORcLOR48QwC49z2BC1kisJxN/x9WsuS14D3YmY3fOhFqYhMf
03jcY7QiVSTRYo81eRhIzuBLAnNWSmOqFsLEu1Jevebx7PGhFn56Cx0wY8ffoC5n
2JW9BB8JG46uJqpxTGnfan3+SOrDdOJ9j8Neg/JbD4PT9a+Qz/A+4mf2aC+1tGSL
uEeP+R69AI+ifIHd9+CLggQ8DYyfQYVP9Wu71oKPd5/0/m5JjFeNDk+a2Kcreixg
24ov0lXaPr6/wYf7y7k1Ofjb5BQr6KiYNJ9yj8NodkGDUKC3gTBYm0T3Si1Mmd4O
7qk3cc8CRbX61YodUCsOF4y7+g26R21fNjyIHr1zzDIOWrCUniyR+2nP0OfCX8a5
QvCAEnA8vDzEVlXH1+jAB9uNxIOY7/WLh/is1MjY/TS38teWljRKegimYs2gEXOn
wzNgZe8mQqxs8QNSyFBLJ1zW/G7yncVbydUzwwlYHancNSGFTAQ6e6YP324EoZZw
GBGo2j4uN+6gLYDW4pXMUEymPK50rTB3ttiOgHZDFSrshpPmfbuljdy3BrHJIIJh
IMCpB3ZwtZP8lDk0RCaiQjL84TwAAI4C/+RaYTBg2MODk+9ucTuiJracE3IVK+hA
fmnuummh/ThV3y08nINEPH+OZchDIoJ0dNz1OPj7hDpsOH7xyy/9ywCZ91OWRCGQ
6utWmdcP3zDLdM6KAZaefznmNuXzev9r0/g9CJzMdesdogKpb3h9GK4pb8UFI2J2
NBnxnKTyMnhKeb5fTctV/HGjI/njYqzy+Wqah3vmCbeE/gBj270yTwBP6+wyJlCZ
JXKXOCiqrphynUZmiy7loef1/5/6y/JQ7f3/SHlJPiWhwIeK/denC/DAt7JyfwZi
4Qh9TuGxhwQ4br4p4XTDJISglVY4+Rx2tqbh8ndYYn/lMYoi+Dvt03yTMY3j+VT8
cfEzjiE0ql3o24UPdBoTZ02sFid4aCXI15AB8tEnA8Mcss8RPQ4b5fSZKSpvgaua
IrsBBt1k8hMCiT6jfl4f5E9AoMJfWjzew7GrdI0y1LaufEgtoORdr5pqFAvGgp++
n6HtbOSjSDNlr/bkdzPoM3Jfws52PSkVV2IXLKcVSG3AmrZEKNx5mbbpdsWJTRpV
0AhgV+PF6pBWda+hnUw9n/MONqdTYwlrgVeTKonsdHG5BqDbeLTxZG/VrTY/o8PW
SzmBXWGA7F8gcq62rITZ+r1rF8dIjlem2jKdsZj2x0O2j8z+g572ZoKK4+FAi7KD
zcaLyJ1KrxVZkK+yu11ZEt6QLWySBei6iNOoduNwslc9Ki76JNiaSUy4T4vA1DYV
+1YvSLMvE2ZGI12ZWxSMQKK0yXN/xHy/P9/XK6mkJ1ZNF9bkJzZ6AVDoUnKX0lOj
FAn6c10mjlR0VeeY3soReWN2rE9MKn9vsGZHQJAe8GCz6xBxpgXoimaG/+f0CA/1
4mYd4bykDBMcxZTKwrUa4m5dHKm1dAeoNFLOss2uz5hbtaz2D3NYQCtwN9L8xl8t
glQVSU1GSrETEYHeQl/3UpJwF988YDd4Lwznylf1eA4TrtDt2AEAjegOHzZhLZQS
kfF/VSwuY3HVX7sEASIlUBP1ATxeLSrnLOge+jjrdGtpCabI8vqrrsRaJSS7vsoT
I67ZbnDVUjubiiAjzevILsj7vmDenCACCrO7gTgM8e4TDVhdM/1CYpUVV2swfMNm
dvwz/9j56PKa82WY80hJqQaW/rgICtH1V7O5k5GZSBmOtOg33Qe+8WJ2MhGH63Zm
/sv9+XPflnyUwaCP7I/4k4BmCnQ5ORcGRgmpbYMqGto0Rj3pm9pyKp/pH1vS9pfc
qCdyEvWIvYR3ZHS4G1Ebm+pOrWBsNn4GjEmJSBy3ZatJvGI1qqLatzAYxECZ8uIB
f4cbwcFn/q+QP0cZ64gEAp+zlNYAy+BT4ZuwKpb249LZikGXji2JhWdJZxPTIQsU
/aeP0hf6S81KuKuOkgTIJXAWe5mzs9rRxbun9btxhDylg+FhpWVJ86lSOZxCrgvY
dTaiaEQa3yFMEx8WVwN9yPu/S5v1x1W0e0hoUTiCdcgMUJtU5lWFtTKHSFhsJDpK
uMFznF24JS1rdljhBk8TJrbqxtug7vndUX8IkND/L94sFSALlj3E7y8Wn68UPNd+
1jTVazeloNrE0rSFPOoC6pvsFkzKItdB8M7LwnqXh0vOKz0o6Qm/ZnbaiextbtIQ
QgE7ZaD/RJzT0jTIpmLuzu2JsG/litpd3w249VcePWINI4jAwZ370jFp0XjNy3B5
Lz2+Y5K92nQgGXfke2uAgHMPhCor2oPOU1cO6zrrj5sSqO/cbXTMhQbNhrWY4A6I
NwqtREpj07pQ5mx+3wAmMavmQvYft3tjNZk0Mb0+ZaXwF0oslt7DiylYH172UmYP
vcpsMCv9BFJpyfyVVggATZq2C5km+jKD1HhdYDorKdVlwPsuKUoIMAh1N8BwHrgH
Bwoeq2O7jrvcfb3srvtai/TSqx0k5v0Ax66w/7k/k8BK3R6MWFayddW+8NOFzFpk
VzAuc7G6ydfbaXZFGO/lsd8EwpEDGAdxi1XbBYkVfVE1YR5s5YwO/8oupwFl91cP
tbB5QkdV1uY6r+Uqz3O9PVD+siec8O7/Y1PSbXGfOilw/ErNjYSDQqE8z/VRlDC/
YQQ3OF5aaDWHTUVd5qtDDF9ZiHRov7InY3ScPN05j4YEx1y2arFsJ1Ch+DMFOQwN
fbGnafWMHsKZwDrtRG/+ci1Jpr7oj8GRU3nPxJc334GsFf1W/ue/rh8S1qx1qRl6
HPDWoF1v3cTzx6RGJDOH8uoGlUUdTRt9pgNjz06lMZ7YSkXaFJWAWrGpfiHpMJak
0pdXq/3tnU+2OLJSgVIA74TpOYbnIdNhpEkyRy6VrAAYK1ynS3bSQqE0WBRzp56S
22++CNzyS4Yie2haW/ikrn8xpOmQ/UWffP6n6eb9U2K/a3imB13UZ5O+Vt9pZImw
IuvSwYcIAiY26uZbDJR7YLjniWLBRKEGsCjSGTHWWvHsLls1b1sQic4aKauQfT3z
JFsPC93Ap27AvQZxUg9gc09ApYsccuZSel8agUP55tb2AEwTZlIZavSmXHkFaQs7
nZDEi/n8OdP9indiEW30VJcewAQe41ljBswE50XfFIiRBO7KkD7w0ZOQwsMp4Qm+
WUEjnRJCpXjjNxHxi/MOxgkjMRRoJCuLcA1nSkftM+1zrBg/1yRCVILuA2wwMOw0
g+f4bu5ShCGNZw315EaiagE/4+bSVWxasbCF8H5XFaY2rncvNX0E3eqkPl7UpNTZ
Qq1voxRg7B/ot81lPIqq/3DogNjAQvIir+sZXKjJCNfi0IlGqqZHOC785EzCaXUm
/0vVkGSlOcXpMA7ot+5XUTHP5eSbproGmsdL3Kte7Y91K6/GSM8F5GddZwxah3AU
5urt+4/Rmx8JooCPZitoZ2q/cmVDOZ4Y2o6tdpzJY5y2Jaej96bxM19pgrie6we3
Paz5ZCb5v/weTgWodVSTgk1vusz+WQZrHY+Asar5tRduvykXbpFibpkPD1LfrjjG
o971vPfNqO/Xwsno5NZof/r/gNz0TxgX0fvyG2Lg8dPPiGVdAveoQxevRPM/hpBB
eEHR0Ct30pkFj+mhpjvDh+wpEU1ZUiHaR1hCzedTxUlUHvLdToBXoQAup8J1H0Rc
6z3wCKFg7QjkU68l4JVrIqSDp55mdH3gBjDyh722yQ6apxZD3yBGWr4lkGwBVFn6
HZHnedR9sqOU/CgOQ6kvweaTJbDwxjc32OhcGHJ9VSx/kcG961kkM4RUgPcnem4y
m24GNnt1GwHv6nDuCWg/rJXJ9QCx31rCPBkGIzoJIponDgc1XJibt/lAdSZEdI75
dl2ZxrZ+VbHJous1qKQ1SUjM89WYwfzuz06RVdbbrLL8t2HD0sePJF78ZJb9I4r/
ayCjTFHPXGJSXq9uAiQe+NEbKKS0TnSsiDoo09xzl7jE8sSK+Ir336ukelfKeTe9
rCTayele6GO3FT0bH+V3v7a/3CVSjfNq6mnB396n/65pUfNzmJrs690EOeqfEJ60
8qmJOZJe96Ut2jUlZihQwR9NMzyEj1WtDwC2e2UwvliaSPaUdVubRrOtxHn2Sf4w
5MwQ0uyKH2W5tM2FdzIELCEN7RXVrqfOsmOJJ6KM2cytY/KjNOCz9nDgzU2GbZsh
n9cMlqMRPRuCGknps+tRmRZ6DvlMzNFGl5Xf8cqXo94iNmaUqdAPFduTtGNPJm/+
bizvkG9bODD2UKt6jDw1EIn8NaefQ+pA6RsdV3YbmPKe8iwOBtHBzX4hh3rv3onz
JabDHmI6f1J4j7NKzwxBLVlOrfkL49OXb46CHF9O/0FSfp5WXaxvfODEQhAzrUph
IbBWpPIgivF7Hdg7Irke8A0VtrFs5nON0jxc+VxkPYgZFUMlfq65AjmAmtWM0ZmU
uLdgPZz7v8QVJCxkcd0NHUBOAq5M3QYPgj0Yb4v2WmKx/eeKq42k5MGH/WmfJzKy
0T1t2YUkRd0RhlCJk6CnM1AdQJS643P6DrvXrJqZVy2qd5dUHaeNNiNIAtBaD7E8
gM9yRS2cEEMFe/hOlyI2L5L01xZamNmlOAzC+ahzQY6uHksTi3yDFpZNeqgTEi3w
BZ+ftmXM6ztGGZU5+5TxpkMNkFDJkBNQcX9VOL0zFWG4YJBzat4yPy4hwTav/bL8
BvNIWl2BwTG2BnINAhlJhDo+KSM9CiCtluSnYFRKDhIa5ArgC0184116Jd5IBs7M
T3P7xyvSiy+5e7uBuQC9Ydc1Kn+XuYUGH6l9TScKh3cdFJh/CB8igWUHCQHNN9LG
fbeGSLdTeSQXzt7HPAc1s1wuG7xrRTM6b6xvVJmioRJ/gOju8xdacok5ZjWFl8Wq
0H4gZYz75BBKLvMc8+RjVwsvgymKomBz9YsfQyWPdbFi7a294hAXZ+H33LmiJsHW
FzO7HGMU+dCAmdfO5Q5JN0PtRiSCU8P3vTMb7bvDXnCCWVWIKL0ilTVs6sUmD5HP
URQqeBgiAB0C8hWBpCn9EmKDCvszMewF2cvCE4CADkEOuU3/J8T/ZpIkiGyEye4w
DFoeic47Cf385LTsAOOOH/MBZW38owWO1H/WxQRvJZpgR+eQ5zLsiH41fGePrhUU
X/2DzNUCBXdH01++XFmCGBhiT7bB1yaNiExrXSVxpjXKrsjSGW47NhT8Hh7e21Fy
+2XAiE3gYXcscIk9TImTNcmUOGFnyD02TwoGwpS/uhk9N21RTI73uy3DARnrzcNu
h87KXN3SfKV9+WNz2NvmfFKdGmXkMa5rerVb6cP5Kq1s4gjbjHA+suy9iRzNivbm
R5TYiPYs5f9wNI3nzflMoHgS2k0QoLCeR6/D07spafVNnIHCxspKDHtD2mkYfm2N
pVawJc676cbg8o/gD2B42HA7EntB1wCyaMnTihaBMTc=
`protect end_protected