`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8672 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
sTHDbAcNdRVMi738hx0vzk9mekMmthT2izIcLQovogG0HDV5PBooJW4QOfsTby/J
rwpTevE3BBVT1en9HL3WOAA2EqvyKI4bH53UslnAokUJF2ZrsYqTu0M+SEjXqLTI
WHVmrlUSOoFZMMHue4evuuiX7VtmKOT9ZMVlswLWyeCd7HYf/e/39N+7MD42Ftns
kDP5ZSbY8+MBrR3X9+ZEWZw+Bv9ITHZkNChchC11IltB2q4caT0OZqF5x/RNo+mw
FIvGo6q5CUAESK4Q/DZTaPqFl1ZoN3PHBKzGqdOw6S1Y1QG+JV71Y72Csrdxh1Nq
eslDmTZd7sxLzZNYZ3KrfFD+UdUcRdwUkr0Qtzg4mQ0s7JwN4yd9B9Gyj86oebod
MZeEOKOjYFBM3TaXSsmUaLVVtxXPXrfURHgRSlUDlbTEFqiGFPx7uKA2TMpufqVg
qAhCrdfUqnT6ks4erQU9XlOSi3SeRRnc54xqoeaqvGvCMfC348+a2C/7PemAriOf
pAA6ijlDZW/ylgcYjInRYhaiOMyr+FsUpjKDpinXZ2mWKzARFZILmXi9CrjjdnQr
OtZR03TMpht43xIuCWve1WUWGPx46FtIdC4SbnLPYyCc4eyPcb8CI4PIva1r3jID
Y7gXLJvLbvdIVkUToeJlfPPejpYtjIy6CamcMDnIJJBiFkmia+fmzeKsz7PB0zKr
uGORyL1gLVVA5MKixvWNFdcLlbK5hf+VnvMZgtMMZNKOtZm10OC/oTtFZ8hG4uVq
8wxSHgqKwDdX86T4EiL19pmdMKmN8lBUUyo/AajulZTJEKN+skGLjOioTLqfKZjK
Muxtlk84xtzH8UOj5XT3MxxRFnlkOZVm2Vud149oxc5wcwFcZi2OdhhlWEqwW7BN
ZSzQCE6MU63re4zQfs07KpBN7nEyNZ2HFIHBb3+tBf6yV37m7RPnQCFusICuRB4A
F72ExhYE16aFn0y3L5mKA7GK2TeZAXMOrw4AzbkECp5zSIoYNi2nJY07B69tMidd
yn3N31QjvGXuza7WRo+M3ItsakrrvZV0DGveknugg4ivihN5ERuv1unrl/l55GeY
lzeYMUvlQab8Sru/Ult6oj6IuuyBfDc6s6w6axXRqNbdxhdbr91X7vHaQLVXVHYk
9y1aYwnUWU7UOInAN5NO92L+68Y5odRGPOMRkyA/qkVauSwQViZxYzUe0RSh+wfZ
fnIaA76VjHY2HmSHzQnCR9bVdHOUVE4R+MrAVj+xJAHM8oihRV4skmh/lwVd8ED4
I86LB6UHyspe1HtX/Gha3i1xQjFb2guMz+3mPppY31riiINmGbsIhfQnnuVEeu+Y
WyjRWPTL+68tvHeMDZB+s/xol2MZDdDWSJCZp0/AdE7xO75QXAE1xZFTWuot+i96
0KFg9p19FJR/bTPPjlOM7vy9caQ0L+RVyFAFfMLWEQ4yhTg9l8U6pt/mKQgLJgEF
9R9klV7g96oI0nBbJHm1dgrKHM78Os88x6Pv1XTEaiNWE7DkMPxUxeHjoZEJocms
/vefr4jwOdfPPef47pv+UdTY8sl7h3QzK23UwuN1OBnEVrKDGYdoCSBNuR3HydZH
LL+QN3tFotsF8TF5TfI3bYDxnzEvtjB6ek27L8FF+Xe1at4sNUlyQ0CeBj20lp5z
E4ntHZJdHDMtil/vXFNGzE3+GWjiMhk9fax8wVR3FaUjl2WUtcUhloEX2c56ftc3
4loMWldGIzC/W/mnPqSLqES2CXdb6cX92y9Ho1yPA8XMI791aLuPGqQA33MbAZId
KPI/Jncv50CSxgdRDFqsCYAhajV+as1LerJgZuZbDQVybYpq5PBMSK6IbE2sRAgO
/MjJnApnZR6RqXhS98eW/vGl/Vl2poRypxH7e0/VshZopUWukL98pIryj1g9Ar0J
ImmW19Yua2l+pAzVKX/OOMovccTaA7K69JQ6bfFI/RKLerP9vWwfbpdfvXhbVwLf
Jnfl0+7jKT+lvfcpZtTsDNDul0GjT7zvJoxqENhwdfwlB3rEMOwZsuFZ9P++up6N
VOvRPrAOFv1h1+k9GVe+Ri/p+c5fSzQVMkmpLigQVDudsKzlogTtSDqc7WUBY3Jx
NVfvuRZgtOR77nIQWjR2/xuxKHcpskVeDmE0Kx6+W/rjT9xAxkyzycGsYA0YE7y0
XU8QDCqsjDHuExX8QALdGITdx3q/3QY7ht0syhfZYXy3cURa8bw9C7MX9LI7nvTJ
JJ9WAPK+UWRiEcxgHhsyQ+fzxIWC9g+Y/cFp22WpuGgtjjE8YtIg/zK1KesXUgv1
C+lUNMl8FrvPmmIgEszxH6Ed5unTeZJLMXEkIzmsiQo180/4I5hoNKe7hcC6g396
jv033rgcTp3H24pl55ow371gG2gV/YQVIDcyQ8sYqh+DTA7GpmtwtMfqQVR3m6lz
TCeEx8IgY2bukVrAQ+9cd8k5VA62fIKGpFoPyr9M9BfpQbGwIjquYwD/aeO/dKIG
0AwgHzwJWD6y1Njzu9qGFLGyPn1ioxjl4cNZk+tCsoC829BJ5hi85L1SuHnUXjSA
4XeXCPqp7HU5NUPCeFexrWnqsjHIccgcTKEJ4fMrb6xaVDzjYcZMvY8Yyq0Nn61b
eIQFtHHJw7FAXzUPTHhxuICIaMI9O5exa/SH+ruGdrxkXosSdivtPP/93b/vAkPo
av9kibtBoamO7voHcLIPINenU5N4fFa6g9UZthQ83NiKXnZm83Iu+HUz5/DM3s0K
rmSzVp6eVsLj/vvjvrMCZ3cSuVt+NxIsWZ3R9WJrPnzErygYRR88DwNJWCpbbxp6
G3YSkryoWghcnchzsqUmXAxMVasn0sH+uI2VhOd8Vc27Bm50TW6ejQeWe51ojMCm
wGeoQboPC3/zuNgYPdIskZMFvuELZZaxqaghWmg5SnKBZcHnE1uCgQZG3igx/Yup
qIbbPvazF3DdNWwpZgiLYsYJret+aQwApTAF73pynXIJyNy+p6XilNqE2XIA4fmf
zO/IqbgrM+ulKdLO6niNirWkBxLJHtFuE9OFKIZnRIQRodZXmTSJHZ1AchjGAPti
b01zzZx3LfXhVXRf3MPbYdM97qtlN1L6BelvuZcYkYRCN5kQLl+urzLZ19kLzdOw
3tcrDeZMklRM5NHipN5rzAJ0Ld2swZICMzUcJykrEJqCUYQWFJvKgnnO2F7WelsH
hx6rbe9GWhAXHsHT8OApdZHh7URp/yFkL51J6+aGCrWVN07xUjexCj/CG/JCEED0
dlqAcCb2AjxwlKS5f/qMwXkHazEaVLdvj1gZU4UwS3eXF/DM+YBzSrl6ILUTziUj
hAWv8awVevAiFl0WTKOWbQkYtklXjTstqq41riLbObyI992M3DylIE/9QIPgSNpE
KVt/MQv7SS3pDWmxsNAR8UTxDmetkNbpNsH5fytFGjg1vB8NZsGq+fkmixyXqONP
5Fq9CYe8FWxQP3WqZ/A2TwvvEcSehM/W6BBmhp9bB74xqERuTJ62Bv+V+8qLQti2
9WSKWdoPdwjokNBxLSRRMrQZCAHIC/uiHE+tom0jdfb8bfx83o8+HxZtOXRYU/Jm
cAWMoxzsNEiW/e9hKk+BLnRyWN0CBaHskiMpiW70TX5PSttGbsr4yECoK7qNGhvX
qQu1xRV78/bEXD7leyVJgDR+0IaxGMgkZ7gsusPOIAWDbTb3/TfkLR/LcKG0vueE
hjwfVe12C38PD8FLz2SbONmRZIc9H++Vd4pH2QfDqC+qBs1/hV9fuo0mc/Y+w6VI
r72OSBhYmetGY6VKKcFq1KnpqF9Pu+Nhhj9VFqYfTHa51Ua62b3ejYI4W3JExHUQ
yHr5bTf6A6dokyh7ceIJBKY8TUSx1ELahHnuenJAqr7HIAggPKTetiGsgUrgNl5L
RMBjpbxJMC17moiGZortZacosAVFm9LkTpUFPm/AQEzbISHZcuTi0IBNROqG2V1J
AVQ7Cqy8jdS3MLZ9jBl7KhUd/Eay/6pIG2iIHmPzvquY0A1q17nHOgC/TTzm4/f4
M8lYzzMdXv5bhgWidYfYdCxEbbIrm++KYeDT3N+1wtpx3swxdQ7REF9jPaRtg6Qe
K1YcmfCzwmEwSjkr5h3bhRjZkFfZU6Eyk6XDv+AslhJ6Wm8d0SgUN19tLKh79Xk1
/gwtcJu45YBRQsgqzbwPtiizFKzxmywn7RgfOzI5EMXG03yf5tusau/VJhEmo5N5
U9OOC8iM/vhrlkwDLYxHvRYPfsn1jLKSA3qoSg8XDTPK4JImP+WaeebGz3ZKzLnX
MWKGZ85ZNgaTpQ4+GGYCFIW1kRtunVojYqiTVbyvgl8+m7QBa4QYF+QdOJfhQuSU
hz4PPCw4f7jmR71yPhlAGOVXfzZCcnBofU0FMyYZ/QhXaahpZv1hErYjAOvrrFHG
+jTEnF3fCuAk6RKbYnK3XPvk1ujBhT6zddJYOvr3cQM/7HNlgwNUzUgd/j/VX77N
UC4XIqJ0xY1VEAIab/xnT3xQn+9WoEpwMTMP6onkGKseLmfwSklylOd2yMFGBYtm
X9EWsgN8WmXb1WhZFVnQqyo/Z9ypbfb2rUau8lhCgC565Kbc4EheObzXcm/fKUkx
0tV3UXMJDqy3wxHDToYWjNESm8V/UbOfO5VBQUlg5htKgqrqwXvcRwAl07iiYTkT
YBqaxBZUNzZU3Y12JGNNW8Uh2hizKk4zVYXQLzAy9wktLsMAi9TMjkXS9Ggc0gTz
lHQz69itw5X4NGRKM1BLv7RvCHur2YtB8nNbm4fGkBCyZsBoH8Zu8lX7J+m5lofX
iETzrkfV3A13c8BHoV2zyIN8U4xoTM9EGhI7tLxVPjOPcbLTTSzqoOnjBmKBe1Q6
gsntcDmxp6HWNecjMK7Xv0njhRfe4jkAGRhi2UOFAPdVBerfV+BXKMQNz7jQQgfc
fz3/0tMFzBALqHG98u2Ac3fKtil9dggbiFlMNENfkn8jQ2Go0wyFrIel4xFZEdhx
e8BXNXJ9bvCIJAe2iz7qFSc1FGhiHihhH+o6lFHedIJ5vYYwefgEQKmXtxv2Az0i
u/pk21FnyXHvSUZdjGvt2vvk+Js4C+6yntBxE+X7/XHX2uyB1SZYhsL/wrnRfG7q
0pw6NEdOV+vKLh7+rtIc3vYUHtu471RMP1M/lWHPJk/Ey0G1U8AUJmdSd9xPVVo4
0aC9gXzcnxnr8yeMdt3xWlxza5y0ED+5XlG8klL5JlMh5RgCf1iDiygy28lt5T6S
TS7Gtm2z3yl8usONqAhQZgPut6o4+hib/uHwkJGN5Thta7eWMIJwObfiu5b4Iupj
DQsFMx++Cp6wc63BWVuniCVR46AjC+xwBMpZFsLAq0E5O7WGbLslA8URF9D/Fw26
vRa9a9/OfwWr51OVwKDekTi4xFwA5iXW7/XOARV78+M+/jGZ2uBUeKHnK9R3fgI2
bMisvn5J7592iPkXaGiotyJVSXWxjhtR0xLjuG91cfEZnDWJJ8aX+A8c6IiGy0je
tEeHXt965mcTKucQbq8d7vk31auQoSduIc5xibAa85vrycl3umzBGjDDkMLCXRkv
p3UPfHg/AcVKA7az8/9SyHVvIwoQlCjISL9Kkktfy5Jm6JWPDbA6s4oeG0JnXVsI
6rQMyVHxgW6EiXViQXaA1a9YDBBnfUarFgT5CSZfdHm8G2URffweLpJL4Iyi0Stp
ta2j9R22n/boTrLgFciG5y1pq1emBtMxCw7JruG66I8wUP+HnqikYWfheMiGJ3qG
umoJ4vdAyFBMQGhcM6siyZqVtRO6GrRN6pbW1kw2Mzshy+RB23pHsyPbaAwRCwL4
oUsMGgSkoy73+ORXw7cLvp5uLSRVwl5ksUfMrRsfKNpzTAC+mFyR3uvRsA05fhkt
n0LJ0MzMQSlV6XmdzzKt4uTAZ0Fw2Wv1zqbxT0yqOXW/wdmqSQo2j0fZUDqLdOLE
H7W5E/muHd62HsdvjW8qYy9taIqmF7VkHbzZIbTmtr4cDo4oxhMIvNu2aekrgMoL
YsSxSFA0ScZqyD6vfc+T2NpAl33MNYN97B1PhQNzh63zk1hWAFLN+GYYla6KpJQ+
C2KBp1z4nRK+yFRIlG8q8ckJmcVrNA3RhKkGnvmLmWSc92vbUkw01zdPqMRoYIDd
9a67BnQkbloIfBtNeCLiQARJvOUq2/ENyD5Yko75NDGi7cl6uUN/pKuKmUqQOAG3
emSh8sdCIwoZA/SGmaEVp7eZUiuq29kijZOuRQ0txk+RPM41VLfEZhNPlqRgsfo1
UK47Ae8AJWKMh4vnV4YwD+vs1LjRPChiiJ+oAQScC1odFUDwdzwEKUZaPAZoFMKO
zUoWtPrF+JK/25DV2PM3H95agw8bmXpATOCKW6aEu48v2+laQbBeROIsPrTM21rC
DEJ0q12Mi7KAQgNdLiYmNWBcltWCEoN8TaoPNzVtg6H7eKuCIwj/+6FWNP1pDbuF
Xa45DTGWFppqiTQ6MPf7i4APz33AkTwAC8UJ/mK/PcQ+MWIm9RU8xcTROWIGe1/r
DGivbZZ6OuWsjtSVHtAFvCpUDwJAav6QRBmCdAE+UvWpaNsZFQ1XyjnC62frz0Xf
dMGV0KXqKtohTH2ICvf18NY+bkaIJv+FgPCa2OJK7wuQ8OOyu8g35InZDgp7DmcE
UT59FZfL+hi/ZnlbWWkv0hXbfCkwPWUdAXnJxphyLXbOqzVaCMoEg6FF7EgGHJI/
/xvDfXapY+FITlulPhk9ogfiykn90LeN1nMdEwFw7cWb3Ys0QLwZMa807zrwj73i
hZzE00UmR46Y1Dvnj0+OVbIVlGjswpbwtV16z8By//vlspfcaCYpRM6QbKZ/FNGT
uDHSOtCTDstI18rkXKl6xuZ+LJpbsIXFDQ2fPlZU+/Ok+mLfEfo5sJ2LBNtMLtPT
tvmqSs992X1uwQJrRwrjVFzAtEc8MVaNewtc11mSPR+Gx1g1cIwO5TXdOXE+/zOl
x0zLzZUL+hAer9zBGSuWr4Fh/e8Hk6nJGyf3Bj+QbsPONFkLcbKtnLXBTAlkTDxf
8ssq3svn7YpzEcb7Z7XfUJb8/P6RUuYnB0AxcnZk0dyAngxehYi936r1mrIg8Ist
TFwSTisyd352iq9xrb9S5VCiP8pBk/HIMHw+jTFLxA2d0lVUTmwAjBxtQh7OqTZi
41utlbmPGCJ64JB6qu1YvWr2quDvFz26U2xCgGpAA/GWiGZJO5SJX3dGwn7P59Cf
FZGvNocGV3ZjwMIcZ7DI13r0KzCEjGEf+EC7oE5pvxvW98bZDztKHFpXh2mykM/X
QwkELJLtaVjgXeOIKYLtCt0O3ChcGnYHVZctq81O6yBANmTQvEAKCZPaGzAZUbjh
fMvrZybsbQbFgOWRP/0DqQ4L+aGvos1VdX5N6Nk1LK2WOStrtbBSGDyBOg87w3VU
1huMWrQvxBi6W2bK2nRsXuuRx1Q+ca0KHWrz8oR//GkMhgoS8L7roXeCSOWifs2z
qKsk6qJRK081ltCcfy4ck46tFbJjAj8zF6/10+T/vhGOet9x7zXieTyAbedWT6vt
SHGFb4xANuZwktV26L6zbAYIor3DRV+MWfAzpDNUKLBMwCb9imjj79gBLTmQP3t3
80eFsrSWRArezFiSMQRtgtNDjw/bGq34C9a3CoWf18fkay48+zPfOz7U4aHzrBGR
0BvNbZ6PwYmNSDyfREv97ccvuHAhyrCr6I2A6uXyNxuqHsWfDPj+MMoDJDShF8vt
BOsQndWhZN5aPlGrqkm19O5YHOm6EvCJrIi2jMY18GXUGLDinV4aApYTl7wiDLZd
JJx2uPFcc0/wdAo6zDznzRyCT63B+x+0hiFI9U0fNDkno1cyMy2Lz+ygmHygMoVa
hxXU7hDAoY++693fzFx+C3K+clfC7yjEcu+fyTdjDdDDnmwWRz+Toi+IvGP7w4le
+hSWPily+jj2XCtbmVJmQhTRu2h6WSew6ju1OgPCUPMww/tvDBLJ5t7b2gozXqA0
gnrCXIQLrJXNnFrWY4O2OVYJQHBf0AcEP63hmcd0Fy9q8ETuSNiQdS1F9bOZQ2DA
gX4oCNoc1/+/f+g6r/QVZ4Z/cmiQPmElEFdMTtLWa1ugZ8aHdTGU/anfKkWG3edy
Xw/TeoQmoIxAVA+KaA1k4V2e8YzGXF8AEfyWxlGoZe7sQCyC9Sp5amm5S/6NSsq5
zRVMfSFaIikPTO9eXUmtcXPk7eJqmQf2GXG6mYX83cMRAzKTiiaT0Ah1ttGynXBS
Twj3+SZItk/KQmVi6xMQju2VCdK+KhlyWjkbYSoFsEE8VbbxmpyKQfoInGiY0M6a
2TBuSQVldaH6ZI+m6eL5kDgvu5EKSmaLAdwAm1TuPeKbVKnuo8LfZb7/awXU5DiL
N5XBJoIEMKe5rHeaiVvwrbFuA0hvIY5qrgTZTQnIcDcjJnZO52wR2DPQb79fMPZd
kOcnwMX7BvxgDALIyDtogIlmXGukvgCjzPnMFHYrGrUvl1ZSj+Oq5DGeYjeeuAiz
TeVp1ZA4M47kW/S5vL3rs8xV0p7pyVAOo3xqPHpVGE+fvHnWJKBviz3CnK7DoSl5
dzUzHRzaSNU9Weuc8xnxhnDfWalccZvAXYkFC1xwa0XlOSEL1ftgYPmssjl54EGT
ibz0Rfmuzvo/jkU7NUdkZ01CcCaw6sdhbnqU+7MaT9OILaZwnD+utlr5zzPjcU4o
VS1hw3WvPGDDdC5jNl2GHoILfwWAY8KrYhlptxVL3XvJDP53SIA1nE68peancxHN
h0vfMfk/LtXwINUZjnixHq2njIKCQZJkk4ZgByPXP/hqmXgnz2RUtwEkwUxoLhLU
BKtY47PmEMeKEKL14er1BboOEpe4Qj8AxmkYa111YKcF+jPnT9nDcNnPLLvBPe/S
Q+AnFlLkg9+4t9uD6qycSOPxIRXpd8REHRh3cvZbHvqBrHk5E35b+Lld5hf6bvD4
+6meWwehrqcfMeZHAoOD42WrXxQ7wS5Oty478ZqswT/Ifnn0zpaMx9iUYUwogp4A
uvKGZ7KgYp46ZrIFShfIpQDfTnHBNoAvPVh6zwER2FgJTuJnNNWHxy6XXy1NJJKM
MSajKkEFHkIjInza0catbKl/o/D47o1Im9tYxANqarmc6XSPBSRzkRo6llJLHz3i
50X5jplF+jfcnWKoRu2vc7TXgm+GnyfDK6PurcQg5fhcmEIoFliJC3DXh0wXVacm
5id8x+v64Mr5R98WrftTh9xvucqL/UO5UIFxCvywKTL4Wg/HTPFwgM+Ss+Vrfb40
UKGT4+9vptEDmwxcIkwPW6REoJGD8k0BXLy1clxrQ0xrvyZahwPSgbPxNba8YwrQ
reMPalHuv7Y6owED6QXkixkpK2e+q+AtQAqs4oeECY9yrCv3m5NbmMepim6x8GPf
fTCbH3nuUtZwehnfqJz1tVrO2tpGiddMCFK3uR1F1FGHK5/I/+pvQkBciu2bnFsQ
kCcdx5SOfGBxPGN79EQW9GU1ix6W8m/wLHapUNOEI5m2e8uElZmitw73TmQM2s1k
LwaMGvPn2PRKywkyyIKWMSpQdtFjmaidctaYzp45KLEzVWJzZtZnSPsxnWBkTL6R
5KtMwFDKlku36MbINlVcFiY046NZCuM1sFBscQtAMgosSdaPejOlhdqVD8vnVP4F
fm5EMQAZVUZUIq0hMXQdvaMIy4C3pKpBehvm8sBWlawKVWNy2dodHJvZTFGwMExB
XeglClmo8Ips0r5fqan5f8b0vM/ElFR5TOaeXFKJIjNwoH+VEfijc0f5sfpH8Kv2
U56QS888DydCD7d0hei+MxhTdJMlOD2d9tgcRwL5rdEnaBew+BtJhu6M0HGbvh6Q
15GyIbWi+KUNOLzXu2Spm64t7VADl5//jFgtnHV2wpqmaRnmZ5aytQ3TLd7k+hIU
pOgmilan8fEEIOwf3T0w5Atka5zTHuMaLPVx/l0HmoIcmUcvJ8+Lm1nZYxD6W4RC
/Ru5RET7Npa1Nk5+ND0CuBtg5HEwseYMa1d+dCtzhdbcqRErP7LZP73mJSyE+wMB
4Aqf6HR/UTZ7FkEsSlMyJTKBHOajf5v/8xfEQ1nnujgFXqL00XcKj+i/s/SwjKX9
TpJzaZzv3lLdhPKhjdiphe+69rZdk1zPUfwyNCCNVTwVqX2Q3wH68M60+I8ftP5j
Iwb+u/v3OUFuBImnrOgo1JNlBdIA/dkj7BUK3QsfUKE8ygRSD6yf0CL+9amVQd6H
2P00dErUwIbfGjXlWQGn51M5wdEHSA9i4JD8EsSbtDyYdWWrLPHgseG/FizzP64V
DWsWbx0itRWg/LUAaQ9avbpx84rPCTguDeLjmPTqMuxTkPV6/dDR5k3bn5q/MzQD
1UQLhyGajncbX/M0ZXmif7TBmfOi4euFKAyFXgiKC4eXVwH2Q01gXhzm+lOn9QEW
ccZ00CgZQoRAUWexNfAX/8KfW++lKJpC38AZzdUcMODkrsM27BtQ5MiL83p58itr
icGAbfNhd3e+dsSO52Wb1XgaY2+VVbcI4wzrPkwSJX0sx5R/PQKSAuioM1QwRpq7
UnFAQpTJNQLsUvvoUH4m6GULcA3PxLfKgTW8ZOex0sXagEehm8DOCKUiDARPgMUC
C8ejHqfAKN2CdEzt68NhnIt0RHZzPdmxHqqcLNEISnw6xHa9zaw4mRnkr4j2d2/Q
TGOuD6k/nS/PvIw5iZ4QYyZJgjZ+7WQrdh241UFPIWameGjkSTvzplBYh8u7rnbp
rgHinRMQCsxbuDZrBiql+MegP/x4OYJhCtkKNHtkR8+eBHoSJ6i8DyL1oFQvIaTi
dC/QbOv+DPj+Px4vJ48e9q70zzX26g24uRFp3rvRkCX6HkdKt/WXKru2pbRNllGR
OmV22tyNi2jPqeRc/a2BYvlooaWZ+H/Dw3Op1DvE77t7fP/h8BX1jnvec+0imS5g
jHJE/QI/30PssQakYkyfzHbixc0l1XAdpdTrSG9GezOONdaJi1pR0zDToxvbwRSQ
ftRXO+U0QrXnNT6kDXqRJV5LOuAFsHm0O8wJTYDu+AhnTcKKRRKeiYHgh3qoexhL
4flsoMraq/aGHkSMcwyER8vQEJ2sQ6yFcannPB8jCWIgMl/IP70jY1vrsG647is6
D0RlMnXa7FCcma6R2EVfG7WYvkN/JLC56nfuIO62CY0D1nSsDoFMwggwRqDj8iv5
t/PRwaNRRTX6i1Vh6snM0j8vx7telT7plVySHEHpHhxc8ROJVk41nfvOTtEN8tUS
MQ4YwkjNqk7o9+zR26KXPi/OYVHTWe9maM1Ntl/pknSPVl+8i14GVf5AyyQEDO/8
/2qjBuWRdx59Z+loPMiWtQWZwfOtsDnv1yis7fx3N5cp94/i4i9p1ifoodwLHhy+
yiQWhQPAz2ElXkRliePsQ8IFFND4scQEcJEUqPqnfV8=
`protect end_protected