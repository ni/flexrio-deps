`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2864 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIbmFR1WQwtULqkXJtzR1e2c11btviVuCKGlt87LcOa059
t6MT2WoTIeILWv777lI9wINyx9X2IDKTy5jwwZWJnJJU1LaXILnN0avb6rlc9EhK
XgGcOKwrM6Z0XkaMwXlgwzEZLI/cZSrsNblf662CBYQ7C+8PAc20EYz1bTAr2fYT
bNzHPERVs1o2g+UKggdXfOqpUr0hcSqhKJ0oJ7JBjBYQIUOftwIUFKJmRcziABSf
0WI998QXCax4ekCh1kGok4gVlGMgGV74brIlBgAFHngfRXWYGFrRB8RTxykUhmK3
ZQMLgWHd2JIQdrfIaovKQqhCgZjLFx7SR0p7Fx8VQkBVpE00CXoZ/yFmclxCaUBD
jbBQDqfGYffrYKJE6KLPgOgDhQFxIqC+JWlM6eUR8BBTCmYl1RLvrQpqoL0YFkqB
JfP8yXFVmVUN428Jl+k8+XbKmQythoBI/ZADqBg6djOWZm3lL+5TH19qDakwtdft
S3oTEFE0raPNOpVDgYRCWGNAniaYQXW5ghWVzlst2452wu/bb8edRk+8wZvC7Ycy
q6iBh5czOy4+eHmIv0SlaJ2V5Dw3jD7o0QPNWep5hw7CcfqW2/9mpogvIm3Tdk+S
GneINfgxvoXkArp2tZ4xetL1loz02dvNz0HWhDbruP57JTlSS8PeCk7WGOLluwNx
jgJcM34TErUmOKbdIAe6KgYpEYCFnf2T4bNNsYbs/EnkEMDbQ5wtg9NvsjLtt9Tj
BN2f7KkP1oktlX+L5mGLlMCjzL82kiv9FxwdEOR8nuiLrgX9Rp3orak8Ezkaqeni
I9qi2RGwqYDZLnY/SX75bp2m0SBQRtCvdSIyH46qDBvn9djHT9KIwO/g66WJ73el
UWU/s97vHcwdZ7OW95PMMRj1TUt5igLS/q6v0end9rVpnDnYMw96xlgUaQBzGVlQ
HiHL+J8E/emxeImg1fAzfbIKSdX+CtWDw/FEzIfvPTOE+SbZtSrUWHBPqwId5GFL
X1n/K9KKXgZoBQ5xOYrj/hWY0WXthcNNZtuYnlEEnE1Tahm+ZlX4MVuMZEFxfEAc
M118O9K87lYpQTJUPi0b6X6I83tt4xQQSroJQUG+KDuSY3oRbiWdAlFRHL2dIMzg
pKL28gZElkz0HvEEzop80e7kUdQrcK2eV/U4HFow5MsC4NSTwn01U4BQhTbLoVXj
FDQtHkHcgCU3RY+9rzN2P3fWzABx2EofV8e1iqvK4sr2aMAhAZ8bOaR3asELDo1Q
Az9oDYyF4ZUuLDZST5nsdJx3QPf+OJOR/Mebj6eN65ToX4Gb9wV3yFbyuujcFJhn
0/kLNeYVe0SuXrYDJeVXU4YnJGEmZ4tp830pivchasnTx+jxxseR+EWgPWSD6SzU
RvS4RLzCrMhLcw5XT7FCVJs71gwns1zZdWLrAo6hRBi1Hny3V+vHtpPwSf6c8PVm
ovcgq94+k1IvZx+SLj+DctmfheMUjbDAtMxi1enr1bRi7cfOZLaagfbgA3lyfuJn
puAI/enivSqzVkR9SqMAqQ9xCVRNce2+Dbnqmne/rRQpjATN5B02w01DeWNJtXpk
Hra4EYD/EqqE7bUfOG4WdBhoOiCAtOHw/6CKZ6op0MZjwkTlUmQ0uCSGwF9KMLak
y+de4PEu3F45GSDZDnjBxUBVMKZfKflYx/FCuLOAeFV5LJqG1Qp7cPj9l0KL8j0d
jMDxUopKXOqL/lqWXgpnujGOWuxgrd/7SarFFn9B7CFoJcfNzzliDaOHxKYqwVlG
vCyw8Zp9NYVSg04ec9sVkruvtefjxUavqncVrmW2g6s2UDjrEJ/v6VZEcSLdlBFX
znDrEUX50DOogXqENO2RerWzhL89UxGgkvvOTgTOK5+JErk/T0a6XosSgELMfwtv
g60fXDfJNbthADAu7daNR2uKcAFP/9x50tJyLUANnEjlkjK9r/0+3vA2Wvdc5xRh
iUxN5K1g2M+s6ojuAVzShGsVrz3QZglmPOhBJVOKS6pahJhK5pwhdFlQzIRSFOT6
eDxkrdCvApooceg5WrUAMFQcJr9NGjgHO0LhhZRPKNQ98/CRzRiQyZqXcfUGgC9M
jVt9mdCRNtNelhGXT3urm0MnOazX8s/ZflBVOh6rYg5kJxJtQCjRy91WUTX5CrZe
XGjVz9uz6M72v+f0jbrKZggGak02DiFsgsjiHCPUWRCbvAH50AoLAwrINtTUqsqv
uA2s+37CBBi14G23fBDDLp+g7s3ZE5q58O9gr8jIyskbhvWT7rpSHgsCNiaLMFTu
UgkgNnmrOzk7ZFpus+XfxB/HKKphvp5mJaubiBSHEhDKXXDRZ3VKlXYub6t8by+O
TatMbZhqZ/zQnkHz3clBkqBWVzzcNV7etBM61EkondNkBOAOGq8QtKkcL7MpAox2
3KfFsrHi5Y2ErnGKiMEz+v+66ilBc0GMqp6vZPFfpm8/4VBFBWxb7rEM5AyQhaEZ
mp+TDuTAKjQaxnLcnzshEPz24TUpDM9J5IY84uVibtQYXPKVchDuZpD1ib0JXEWR
KHyYVpfH0y6dvrOq4FxRsufOsy8p9vcW0nmusYghCQA1NbFeMQnoHYjemNdk5NjI
h4AspthzilTaitTv3RLfNrCLPOuuV1NNpE7mfQsXRq/vuWpPEewl7KxBYLqlQckv
7ljP1MHLsak+/BwY5ErRT8JimELtD7syHqc6nmZ7RXmOR/swBurJveUkkHadt2Kw
lY+c5E/pjrJFl4lew5bOmYWHh/5ztWk3gGqx5ifIGBsoVlW9S7FdPGC+gV0fu9W0
wCb3sO9BMMIS39lIRQx5yoBp2mTf0IgsrjXcaM9NZ+cG/2TlbyzAT19kdxKdu2hI
NrsCSwxYLQ/c13zO3UMUZWXo8g9d9jRUo23lYN8xkkpv1yKUzjBcSOkh8B4GXiiI
dqd8U5t0o8e0iYxSEYcP6kNbf9L7L96020pOGCq3yBwAJf5rx74PfZvbvRamNUjB
GzmA9mRbEydzwCyJQrEFy1Gxz6K5xZ70tTcSPSSOPpNrEXM2Kj5J3gcU96Vphro0
MkCWk9uQAPNoceHaOe2REPwJstd8e7xXIQUmGSic2RZR1cyp1wZe9H02upir+GI6
ytDWPYWyQUIwRS9ORaEuc71PIm+BV4088oF62f4B96Vp2rKhfmOk3Tb+IhwT0Aqn
456/UjO6jIndhj3rmlDMBMZ4iFsLiIhP67H0ZgOlOid8v68Q2JNxnxiEdgH/PWt8
i4gcww5N8BgzZ+CNeRLVUe30i/fnRYmnlNrlDKR7xTVNVWdBRyu+Yp8XMzfrrbxl
Ncg5vBKrhnqLIHBWaHJNuNFyQesnLFJwJNDWg0i36WmV5S25e/rN3HYnW014ITZY
gitbnE4eiNo/yvZJmjeXANp+Tx25D5CFBEDEX4uW1oP5yN9flFqv5S2QPI+iEjRG
xLPRyfvmsBNx28SFj+DMeNU5sOz6nx54qgk3uSaF+QijimxiAstYE3RjcOA8SjMS
2WxGEvqDP2YCPIlXMLWY3vzBotFfkKjhDDXKaVLR96LjwNoY1ta837iqyeKK3Uf5
5x02HO37ltj6lbOu5TY/xo8oSMVbcuBWuXgOz6Q9r+4aSDsHjK3elQMim4OA6v/0
DR3wZjvcFSLLyUwIds70XiuoQ9G5sRxGx159TwvKJfA=
`protect end_protected