`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36704 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
yB5UT5oQgw999PzwDg9vErTOh8FvvA/Q4z+JMZ73QjDOPWFIKsfC4lgY5YkXAPGn
LBjSzx6GQfHt35VxgCjVhVJtyPUV4M+UfbJzNB/75gR/fO0ARzwzuSSs7L/0wxgW
ngTLxSIAo0XIHc/alhQ7Sw9fQFTsz3ErAGxkRKDvefyROU/oC0umWKN/myt6/iYo
/SMK06y5nIm/+3ouh0iLBOEcL6rH+J+ayXY63V+6OPDRfciG47B571DB5Z3aIouW
M0CKuP1YYyekv5hX4aewWF5CnNqeqP9jQfu5HPuYMf+mhi8FzYtpmwIsD9tXAImR
tq/0Ywr5tMtLg4oMnx025OHmC1xhLhxry/YUZnNcjHepB0LmjJ8oR+gDMAnru1L0
fSzGjcPuYvZXeA+Og2kVz0ZZQHSnfxyl9U3WzwkpfvIwMEJ4wl+0B+rMIFQOs3xS
AEhAQ09n54q7OElw6jqncc99sP27V6HkB6KLxYtt8B4yBXAQFtusPOA/8oXUkJT2
vrIFUKlv7s6JGy3kfbFQp0ik+Fb+egoBrBeZK5dxfhrl5heO9lV0e/kwDJyqS83s
Mxoyljd/wtnjc9JSxTQunRgQ5N8/n79q05OsBh0tcYo1ulmIwQtwhXprtnlErslk
zGccFE7XOn9TDsOSoM2CKAcllFFaR2Lf9n+/qg+qkLV/U98bX85UAzn7I1VxEmrG
671uvjewAVZ/TLL6pmtL6D6Dld3Ipzl15uNE6gNRckpzGe+Qz/KYuUKKZoyayc7T
AL8qUyPHPCaDA0LBQWFrvC40S489uZmjn+9bGAhLOsPaI3uzXQpucf+nMJImmn0G
vXodThN7SAdSyYknR3xFBGoijlhul5MjbzbfomdSBTpWNA5DJBIYX0TJPnqlIpiY
/OPskblSDKDRe/0lYVVi6hIV842A9TlJQs6jxxGLyoTAmvyegnA5vtYQ41gArqwf
iZzbRuefelgHukNb7/1hUZRDti9xnqVZH4xiGN8RQeHbKoNTBuFh6nj4iXILADV/
gAf1JTJrGSUZQxwEtwWzZHHsCxhtDP6r6tyEMILHhEIQUBAvbWqhDwscGa6/3kqu
/8khhZLI7Oe4gHGgHuw4CKBUhwf0eVhNo2IeLcdd0WxKaUIt+4yCeEAuJ+5bJ63T
hiRcTPfq/AghW/FOW1QhDsV89KHHQ/l+hDjCZzau+LJi3TwFpMqdadcGKmcAJjCj
clzEVfz24UHK1s1RwJr93SNPFY46IJG+DVyVlxIgMJMk2xORQTFIHFVJA+Pg40dy
3PSWwjFvMgjcKzlScD8ZH0klKX3LOkEHGByBVTC4Gppc9m5AGHqvof6kWgtkcOel
wv7kNbqljw0aVqgkz0zdrQS2ua8fG9sBNhSs8PGIbWV3NXiEvJpQKMB6BdTsKDhG
7jKOYCsLhggNhOOBYOX6ZxFkfunJFmVHlW6NKHo5uL5Mow/Sx51rT5L4clrM+NKB
cJlBQkSrXnW9ESrcKLYGqQVHwB1W4l6XqNXe7xW/lNTz6oRWol7C4zTarN2vjgnS
eFbsUDuc3hvUseSBNsxpgWH+EzA8u8shmLZpdGCjG6MF9676WyGXcrbYwdg0suTe
kwQQDXUbEJLQbRqCFZFcdSJ/eeZapqYFlTE+AvhfrXnNKUPhOv7Q+/WyMeS7bdv9
edY49jhTSjovbI9QzpQ3aF0A/OXLzlbG8n0kzO8i4VlcBueJZbmFuFFT01ydBvgn
6hygJqbeyoVgkuv/1NLiXUr2m4PEZ80YoXklEXLtj0nerbsGiORDdrn0U804Fexh
O9HLT/BJIbAOa5Asgd8s35vJankWwgkqH3UQtYV7ybdFm5Q4iycKiAK4UjWie2V5
fo/Y/HbZpuMQgFq7fc7R8a53h2A16a5Zexjcs7VWwiy5yIxECpO0X2FN7nLb9p2U
GqKBP+RX7vl0omzWmgyBo/Ifr3hJaVQMAoEDW/2E6yt9RjtQvY5OsCwvBJOPBxYU
v5r1d6YxnOB7ST0EY0oTSw0IkFY9xxA1Lxn+MxHhst2Kw2IsfDNnNpG8+5rfgIXh
+Xos98oI05ViTKhIi49xzSwobLPs4R9RGOW0fnbfogtGWNo8RxcW3CbVefFZdqKK
J0TpwDxq6un00ozmUdqkCUbf2DsPpfWKIVh59ce0Xg+kkx5u1woOgM5dPeDRpOKq
/o88jKMJtl+3OVaUO8K3cXsdyXLLm5lSSwNpJIltTPrYJxNVinf6/EzsSzvt8BEw
9gwNEVxB5moM57Om9FeHyeA2HnsFveXhhOIX//FsV321MnI+sLDP5I4n7mktVYyA
VvPs6i9BHROVgatKPZhqM06HN41GRXK87mSBDKWQSiSwPAIEGi7geEAVVE8plZuG
BtmNxQNUN/sze53abEd+6DkHzYxzhYNCXRRd3BDKGt8DwT3DU/2/U4Xla4OBE9ZY
pb2jNa0/dWF3RxDBiOiyjfozT9bYrmF8T4yQK4yBHQAw1OiIndtu66aaxsTYgp98
yz5s6JjODf4l9ZhvdjxoU1q/pTtrkLya4DbXRdqrXTrBYMB/vTVns3ybQJUodKR5
UCsaU/VzcSSS2KUX18oNQmU2T395hvQBdqiINXzs8oPQLGc3+7lq/VY2UiFTt+j5
lutOuXkDrjYOMlfYj1YEEShNWLBJY4KY4naQ9bPjSZB9BAMJRt0TDsQdyzhVm+yP
EyqndXcmG92jUO4F+wySsrddEkxPB1IGs5B//Xw7ytnNiIXXEn24r9JeXdpNIn2i
D2QbUtvnAAoZ6KsGHDXsJSgTj8EzklsX3BDIFDBQoeOufjDzpvsyOYUMZfewyUML
MMHeompw48bl77iRpt36RgKOXoPZ4Rjrx/6tQOgyMKsh45uI9XPMY0JPNR7jNtau
WRAj6kUlCdmfxO5f6Eplo6T/mwWXk4xg/+FH0HlfuGbV8OtFdIZVzGO0Uq5HiUCA
xj4w92E44IStkCUJBK5wDp1cd+FV8f6CezsJiUuXCcxAHd5a246L4OVwOMHb19Ac
oIPA3U8o4OXN3j1Nj2UOn1ototsh8v36ZDuH4NWDkrSEVo62bgDKRy6IT53uXspa
1xKzgGJyIg0WaWyfWtKr6qMxXRmhopf5Db7t2yjfuEiRaRPMiRmp/t5v0Gykpf/i
BaCPnLVc+e9BYi6cG+S6me9JEfLWVGBYHbzSTXghLnlzuc9P2/JyA4rxiGEsL25y
GPTjD/XXK8iWzeMpMY+fWdOWNrGBiuTj6c4L2fDd6xF+1qjDFt8XF0Ug6O4IWwkE
3uldaJSaAIECNiHzFl6Oy7b4QhODvXyx1r5IzCGIrhPk79+iPO18gD1uiw9vvKN6
asYfj5E2kFStV6QjlkMmgZdk6nwwHX8pW66/vegpsir4Di8IbpSzCwvvgfrhDSdx
1LhwzbSjCRqTyjCEsuxsN1p8NU7BDuh1l1b12bDKcvDiRig+dx7onKWmb8YN0clW
Z1RooxtaDUjwjXsEe6hxUFAQiQ78I3zN2GEKbyxJ0JOG2msayRpL76bZXBiMMGWo
Xv5pIu4nZorIxgHtrIjbUvO8bc2QIwyxi9HYfp4fpaYnp9yLxCVO91HSUTJy64bo
eQUdfSIYrPmL20EqvkKAEGMFFYK58bWLKCTyIMM0cgxM5bA4RnQVlqVxGY25zf63
fqTmhyl3FIXgK64og0CjgL6XJAKbxzjou+RBoQU9lr40o6luvNbhlVlESHGaxpJy
hRHUWDR3BtSYqzK7A5HbYo0dl2zZPFNhYkYwtJlMMXms/nY5zi1km5MdHOwJm7Rb
9oaNUyrUpZUFQeVlRH048a+TuBEoPCxqGWhV8sA0LSulQWvBiX83Jo/aB11JD4Ly
QwBLtu/FIb73ogbSTtr1GdOGfRS25O8dJNNR0hsolguyxMYW78Cd7PaOsMcVJl7G
UygE0xzoZ/k2PBvXfBnC6eG25aFJ/4ad56UUN4ZTAx5bjQsUktiKkHwYxQxoLpwD
DwMg8sFE+HLvF3npIDE28sx+nQ5RMZtVEre8xatpASaqYCH1w7ADgAURUoAdlaw1
Vk41OqkCDyLSk+BRqVTviUgYpyVZyP+QOHQZ6HykcyhJSHvLNEImNUFP0oRNFL5w
90pymiO9FODR7O7ukKczH/Pa/82mfccAuPEaR9eu90IgWxaVDeUNVvrzTYtnsIFc
lvKoC+dVj2Cmb9kqwnF6eLs9mXEPGKSBeIVk56G5EnZUsvkXvZJ2QpOC/WDuxOQR
EOBQMiAxhZYktWxBnGaeJ0/QteAvaLDNCh6iTgUHh0KpxkCevq8Azj1dDlgYqnCK
efvnbSO9p9NpVKB2lud0ESRVCxeqHrduKSsEe3SaPATGxv7ovV1h7T2Rs/ilGT5a
3Z1Mn/eGLVAOKDyrXgjUiGs0imJpPIknLcaGNAMJkhWjWmA+NtV9rnnfPt48P7zT
n5pwOCedDDw2P1VJVoS3U2UTDQWUl09itLO9ptAezWKhHT7l4yChlWJj3N4r9hoP
8/7dpwNYvQEud1mRGsSnNOiIXnP9wWkdeoLk3iZJmMFakRKwCTbRS/3RuIxYsGyg
7DRke57nEen18K1lVzfU9J8VWev5gJfvDrD8MoQxxKCqlv/LH3s4jB31XAnOqQVt
bHVtAfvfSEbDlz3WmlkWx69z4ujA3s768a6N5ZyozSUYclDVIfEAMSyFL/oWMPeg
Iz2YD2aUE7t/tx0Ff8rTtgokWOsRJ/N/8lkZXHmcBRnwNhrjJufI2toRBsn5foyG
OeIINF2b0g3xpXrg3lEGEbr+vlHYtL4yZJ/7aBwiFpxQuVkvu2EL38VPrzWrXVN1
9o0FvZcnOpqoX6awUuAdgpHA86eeGk94HiIelHLW4DX267SQBiMEc4OyJwdAHf6B
s+zigraXr2o4e/U3k7hIWh6Q/btuo2J/eKqhbgHuKHOAxUFDVyps/rs+pKgI0iD2
4V8JU6KI1v2PytGrE6HiESjDaT31xmz3vbB7IFYn/DU96E00P3vLgfBmY0kx6FXy
rVX4wTi4CW8vwLeryI5aSAQGKrN77Csw7dntELH/B+ttlBT6B17crFbBgiF/VcAY
e5Nvrlxys7mmJmek/IOP8vy7E7UFeBEU8AQF4EjCOLirTbOb81QkXdwPaYfzgJFa
aUbzq232xCCcBGtn0bbv0KbXfJDvAPtHqXLvWsQ1FmGD1f/FRB+a3sKxuTCSuMmM
unMIZzDs8ZrjM0c6RInlPHzRHq+9/sDpmYgf534m8Np/7jd1K1lZJxbzUsWBk5RD
e965aXgfnV4JH/pf1K8iwAaPdZL7szSiBvdrqudoNNGdYXUdkjDy2Epg4ztlJvNl
7XG1g+0IVCs0iLcWx86uBFJ4KFnQFV4AE17VjkdKlI9CWKQqDlLuDUoclz703sBX
Zwu9kh2KewUuCJ+NUEQqO1g5XtYw3yIHy2t4kRKZY4zrdR92dORoBmFeZG+JYTkc
1ZJW+59Z7KuWawQxP4go0Jf5dcgjv1j/tEgNGygrre5zZ6QII27u6lVaDq5eL47U
vuzOgNXJ0UUdjoGV4GiOd5BcCdI/vmqAeNxJC3uHvNICTgmO6OXfMmsMqWkNUfSA
A+80Dz4H/xTUfAJqyfk9U5mHUW8DxSnLDEfySs6ehlOTM1G3k21H1Wt/YvlHBglF
sZkEJdCtPEnDXW4LgLSp7xnlRTsOOGiSwQ0G/8JFYWVrNfhACQmlRaTKnHg1Ue5V
RhiKFmq24T5LcA++TsDh5+RiBLfhIAMyVIpFz1ceC6XS7ibDA5i/gp+4gdjV/rJ7
Dm0aIIJ3VkH8V+aXjVABIqgAHi3a6hFJPWXWbof8lEn/VCwd8/eHI0hmQQGV/wCI
6owNISpw2W2OdrvzZG1iBxW9Z13CCVPRzaJ/0I0pnfi18acbAj5ru3fz4bE3V6PB
fBoId+wuOaeIp+eZC6DQBHFckhjFKwsiKvfgVEFGxofvZo9QOanPf240nSuKInuz
U4nuL7TtjfB0VJ+oTlWnnWzfOwkrr5ZsKk27oenwupajBEGB4mG6isWW1vIKcjOD
lDlPmai8VTZuAacsrJfXFRCAvRHxhJfGvhGNlt4VwfVbsA/unUsFI3DKHyccsxt1
FBNZctOidZpjrxIdDOzSCu+mWMIakJ7Ye/Rmh5GYj3erWiI8bvNZsy5lAFY4Y5wz
59JTrhZDhYotvdJq1a/5T60j5NW90k2YpIzafUMxwgo5RMgQoLCC2ZWia/AD7tAc
XPKa0+OFW9RH+3R09oTTFqFWZvGcitGxDtdJhqXHoQQBkkhR7brVO8Ou2sy11KSb
rdVbJJtaBrRLs0VUPlSMgDdOJBMUAsngNzkGf1l6KraV952AOYojv67NmVUcLbts
fr8f3jYVfgC4pXZpDULgUwkuRddIStQLjAo1sRMuSIEBvASQo4k3pZFwch9tXddW
qpuFxFwwKE9xSJnIADa+PyvrSRRJQBZiWINLegbdUaHH4gzXaim2T+JchGjqcj9W
5MlyJQT3b5JsaPxbLgrycV+1uzvu3cYD1mdveAI437e9SqXF7v3TnfKXWmE+C+Q1
y4HaB6pIyjhALCVGByH3CmrBg//ByqTxGSI5cGcojY2ozmxkIstBtgXp4mpY7zrR
aAo2t3zGXLs0taN6hEJhFzkcKP6P8STtj/YoO/jRXycyoxEbPJnt/rLs/Dda741J
OVyJ/4nS0RWVA1elCyqk7LMnW20SwuP7Or/+zAU21UpLZ6xg50B2CXULVdD3z1m1
3XYytIyGdDVYa+egbT0F1zjoboKrJIAaifFUjTQhGpBtJ/jyVLje821S/Revu0ks
8RXofF/dIancchIVIXjrN1YU/S1nSDpib51ou3lnfVCZyN4B8WJcKI7026GjYUHT
NMafqcUmmlLSK9HvXzvFkEWUni2r/LSsmtO5DocW2CLWOrD6/AKGQo+4DlNAwYQy
8znENF2ga50mLoxB0DEpE/y3Ab9vp4o4ocKUGeClyyWsmLmH1gaN12ALizTxDXMK
gq+z6ugh/fcLsANga2MdBIo2mvXpuIdo9J5VGEbXSSh9UjMTTwp99ZksyBYBenxm
WAiM2nwLNqo6Pt2lVOaMMbbZ+ytQue/J1XIxKYZlONQCuY7ReHfqamjKe6YvmCdK
Kx4ec6xX5Mrs0/NG2iXOw681JmJDR8ThL35eoRCXRoLQWPH77/sdep1DhWi3vR2g
IoT+RS8b5r6+OMXqZaZ9C9q1Gwg6LtfKRGYOkJ8mOxJ+x2O3YLq6LyP4XAOWDTBr
7iUjUV906vLEXhhEd6VSAiRP3ulEL+4eWcl09o/1kz5ocxESfIhEdXbtm8qocYFN
7Uu9lqBc0i5qkGZkLlsHZoK6/WxrQVFkUIYDv3WxXNAL3VlzD7XOgoTLa5MPPo51
/Iic+2MNnsJsxUoZVmYLww+t1/FMYh80561mb7yoH6IOHcLu+tn0+7t8m1CwaH96
6bo448kpJ83H5Rqy+rOAkEEyzWPUwj7RqH96bSJiRsoALTrKxrkxVu8/mO2aC/r5
yPooqos7GoghIBGmY1m5957JdLC4+wN3J+5PcLeJmCJvgjtWFIVu/TkboJlz+xHF
MYhUbw+ycuwPaM+rO9xvJIw3R/f7LY9SYApGhYXLUicMvlSc/iOJQ6VQXggUMMB/
2MZxfeJPyFApdirN4XTPbAeezxQlW05X+osEmVzQxzKQlIPCdw8RH6bFw3cvcIxF
LCnWuqAv8X5jswTvRp8Js2cNqEA57oZ9goSR1HBoHs02t/o4eEOIDBThTNTH3vMl
Me0LyB7T/ObJaw2R1jP7Ozdz7jbHsuqG7Am8tT68M6c8zycdcLXZ7ofQtNAtZvTK
3ECszFQsquTeCYLhfWUKrXmz+7NjIJy8K7LLyY9TN6h4fGWIEdmjHoP5ap9CJbJ2
DLQvZ9+uwIjLg+QGRO+JUUbZBlqJWcEdY9xhqQKNYdG6wAL0Y+VSZ5sywC/R/Xjz
Zkbj2ODDaMYyOvIkTBesE5zwMuTkyKfAMcVnZsEDXPOVwFqkomtEqNIDykYpvTtX
LdE9ZhcFztwgOtVMfXNBZ5SiJbjwDlldYYZeSbvGArQTujU96rWMpJz/Bv7xMTOQ
oqZpjm6Acf25kbxsQ3440TPf5JntZj9UbB5DfFq70Dm5V4NHi2NrbozwuJXXpkyt
vXacOQTdTig5DlHznIOpq7qKbghW9lV7q50G753ycuwvBFmAi5SJ4EXbsMqEKMKO
9thg7HORod/JnwgET2nlhEfQqaasv+cTQK7KiIC3kWjjS0GtM/GsbZ2+xNMLwTMx
SCsnibeFKtz3IGkh2xomaa29azxyi6Zlbawt6K0zGc9DZ3biDrH40x6tzUYlj9ro
105twGF2TjpCD0czW/WS6bezrsHr8GS245vKJXlM8yTiYs5VRs7yDAa+sxhdGeH6
bQk0vDKpLlpBNdcbsf+F7TG43rjVKs/uiCDs/LUCWmBUBJT+lhJP0DBwR+bwUChS
FaSaNN/o/wyZiy9DR5f6sTOtwgo8gyQz96LF1kQU5UycBzeEAzHbiX+a0pH44Zg6
H1VOZ7idPjLz+9V4KchBqySTphzucxXWSJQkJfAAugKVokpaFtqZzqsEVsmS8yG2
noZc6BFt4hpi0jDBFr62xMTcY8s/BL9l+AOiYuNcu/LmBFynMRZasw2hFxdZ7Qzp
f5TdWcWW6PZQ+M47JXRylIEgxAD6udSjrfJUkwjQlx2JW5mGlYznxThRzyLRBNFb
oQsC9ZfPxmTIkyEnZzgGb6VzguHkZOJuMW10q19/OvXpEIeB8cw0HB2/A8yeRASm
tGtQAuQU7j4DYobPyUbflHbTg5ff7/plUB8CPBPRsO/kqswL4r+gS3y5ttusCViF
nTM6KgblInWSbr1DuWKgi2H6tT0emw/tFjDpbY1mb3Yrg+LxXVATHPKztJIoVHvp
0ihdFE1oShefKFB1nWUE9r5ACzWMa8Cvg8zgj6QGBMvdysGIHBiOoIxtFTj31/LS
8tP+9m9eu5D46DKpjHPVCuUz4fzXwRvwCLzwhixo9hRNIqIWgBNmE4kDJ8hff2w0
PmMkjoFZxm06Lz+MIaVl4KtoI6KgXPVhcTYR0eAdCGkiRfnq/Hs7L8uKIEYRSAyj
0dWWjEEPJaElxVUeXuQi8F0qSczMF51INWd+EkVr2eyOMhlIY7ECBW2oUaaQoeQN
889UVWEaPzKamC8jxQEnE8mopIGfyhuaSubaxSd+kjXCJ0INAygVf/lFJGLd6gpv
+VGSWSzqwewil97axNGPFUJmYFqXftmj0GMQS8zXWjCJFsHP+Ie7lI4jEUJ4vt32
EtpnVLH1K+Wv15mkBqOj5+BbNlnR3gqsPyMvscA1jCl1N83jj3JLGoWKXjqqSM/K
5CFSG80gnhGoFcU5+LlXs5MJwDefF4NWy7nCVXo0wKmFNrU1ws+ZnN7YEP8ltsfO
tQdDkgo0xvypdTi1pZRo1uQoU7ert5lvMvuzB3UcSdM3ly9S2Hf0ug6gvoWTAHgU
6i3Lpi5hDNbjr85XWyEpWcb8+BURo0iG9L/j1+wt2turImqjLYOVe1jslxEXxD/X
3Y/KpJMmN8vTm4hh/5O8Jp32k/uEFSoZokLA96X4XdnghWDFNtn0j0LsDUGE/Y/6
cl11J6EJOAs+dNGEKZ/wy31B6nlZmGnDqoSHPdK7z4bE4UxyTEui2cymbBKRem8u
QcTUj6ZBeBj6DB2c+xrN35AEtV3PjjIFYalusFPYiyiBHoqKsspuynkv4bmQGMxL
paukPAIQ9c2wST7SfMPD8EhkoifX4DXU+ajls40eYZ04dl+qg6Q7AwzYa/WfiqsJ
euyBHo1tqQFvrsxWkfMpYx4z0C1HZhbGk/yyZjpsooPHSovw7I0bamyp55XsSu8G
Wx/FrqLDc40hbEU6t/fR2sxQhQerh6/wBGzecng4DC8wruaJpyZ8khBEbmteBme7
/6T60a8/I6a7df/PsSw1YK+7LlA4w87vvSgj5gUtdKtyEHTXw+YrDfYkrOTQJcBZ
u/oKTL7HiKKwXJalEP8pu/ds+zxos1Dj/B2gGmh85kFn0uAzzz3zKC0FmoLMr7Ed
G16ZWYXLCtbP80neNCncPB8uNhhq1CdnwxOLLzuvoeXUE1yS3R2Rn+YA/UVeAPm3
Wn1+rZCwm1Hfr0JlodGAxaVjpDWBtOMhkDw+bgSSKhNIXi8x3ylTyCh3IAlqawzD
aBIrCZcFahDo/ZgWs+whGtiAwZoy2XxfphAEDFiKEfWr4kpuf8DqUVMFOw6JLXkT
WYBpyEVj5jxjYM5o4RDhHBYCXpiRJIX4TCy/rMM/IG+sPhbkp0t9nwPqdIDp1NaM
9rPygU1M0jPPkFnklkOS2DZEreMedewrEwGTFdmsbapCWILO2cc9FJBsM5wsH29r
Jn3DsejTSC9ZhpQWBuFA1zAV77YXeqlVBctNqfG4LtJepyOPpksxOZsTEqx5vAgG
J232BaASVvsbZ8KGIg1qh5c2Y0/017QgtZGVuGStYNtLAEjhXLL3JeLWWYjH0VdK
vdG49tDVz6ppg+1UcDq5PpP73a4Mgc54ofWQdLhJmbHMvxjelWr4gUsZa6HJaW4e
R1cOC8uG+GxhRmhIFktbDpi/W4QgKPdt2teYV5xbajsukhhnNWZkn4Ffz6vtBo24
Zf7EwYboUKuUFI6VzE7k7FCCzZ8RH3GNKo0P1UxwD0EGJO/y5ObuxQMN5kVBOfRn
C71Zd1LsaoyQdN3PmBSCf8/j7RunTKxh1u+p9CHAm98Th/zIWZrNJZk/r7xoFzJX
d8OBgeFVmVviZWHsh/MeN2GsbhrwZmuENZoLXEe24jlSrsSWg5WQfFc8HCBoNCfi
oFkDICN0dwM9hnYjAHidJoW+MP6ryTdxlblrLVovtDYS70z9fXPqx+q63zrHmDpx
w3eke5/JFJY0jctukMqrbwj/cn4ZR51yuNINDpRF+kT/GabfN/Tkp2RXMri+SqBW
mh/XUtTSw6y2lb/jz29kbcBuG5RjsRnLruWs1uwmehth7b5A8P2cocxcL70Ue+MC
wjojfjgylxYgu39bbiS40txdhH+sjx8pnRxnvpJ//S/vH8B8aKG4jIUlsOVeB7B3
B440Ml90lcA2/f+90VUdEdBuAjUmmGYbVCKPX4vJBwqjkcyevl9YgFZ24mK14JQz
LGtaHHdwi1onEp58gaYr79STT7OF9SDO+hHCLdsoLYKIt/F22LT9tLSEqgGbpQSO
7TgYB3l/NTo8VXF2VP+ebAUpXCFeSIRWkl7OX560vPnrXnyoF/0vcFhmrLkGyKni
xjQ7W6oTBGcXcOcc8+39eXBN82rU4/na5fvhVg3ygiXw1moFqAI5jVAfoDfwYJt7
NVRK0W27Aq4F+NpzqnGt853nMI+KgX6pr+M4pOlPlNdarlfwK7gUHNMyTBCSLhYo
GZ2ZmIFJZFDXlDLtI8uw8yPwyeDbO4zYcHHkUT8EOHZB9sx4Bw4jkaS/5OwYmfcw
lcx23mglalTSgI/27Jg1GVdy461T/aPiGKGz28dI/8idGbgWWSsv+zoIUzl2q+sk
1J7yKflfyQIF06xdYwve5M2ims9TGtobPkDMIgK4MA+3l2ieNDXIO1kMJ5nPw9za
lGj0nwzQd4dMDZRlYy8S7hUqpnQFDJSLolBvnMtBiVSs5kJAtR5pSkHkO5aXl87f
nMz5+rrJ8h9cPidAKYcWjXRwXjiJhTQVjwdSSBsR28C72hygKJiBXw3HPKH1lWjb
T//0hktXcs/UP4hap13YgLW96y/QH5JR6gPok3fwmlFIauOqYlLdeelECafFVVdq
ZEzem7avK/4OoH592HL7sPR5g1hdp7KClhkGGe1ndir1m054JJ4JdddBOZKdPYC+
b0qKY/h44YFGdPOnXx92po9Ro6vOkNpgmso155MByUN+FPB8X5iIvsqm9bOS+KQd
YoltcPryyLazmXIXPjLt3U/ywlvHbtWwuymj6m8dR/kLeB+EDy+EVJd3AahXugAQ
h++8j/gmxhQBIQsjLFG6hvi8dVD7+YG04eltvafuMAJeq5YIo5scCRTpPPGP7ubC
tuzKCmtdsIJ7evycrul1WmvbVyCpivWlrHxoUti1ThsWay7liudFAxHk8/cxH1oz
QGgm+8cy0JDvrCHYx2A5gQEtwpFjUPbQbGLapy7JPEMCgc1uJjOD5cj+sZ+XzPw5
adjYCRNOwPD5ZC9ND0uTI0iUc7QVXq1o+hyxw2M9F933vllL9h6XWO1IyG+YGh3N
dMJLflXFy1sKQcu4FEWLD2b8qmRoEuNJCESt0OxwKhsFC3yXAoTh6UQ9WW6/1hto
f5lodoV/5hv71CZOwSJ2EX8w+90ExMF4xzu1ud45Ge/x4PZRGIh7fVBHN/17Bhyf
dLLzBImTiEC8kBW5cuiTBV4NJnPZAk8iTPUsY1UJs9j1A6ioIDOwDgIKTxcY36Kk
uZzKIx6f6VlbMCUqsWvxDtzzEtolsbGYU94qp4OTK5CkYnDdJvW2s2BmJ3Gb4GOu
PvWuhIvMK+8tb88g3+LlQMPflJHtXVqm93GqxU1/Ogd7mzjlYX61Vf2fLBiJvMfz
ti5JVSJarjumDRHBr5W/1nn/kAblqgaRNj5PECPtO6Qdoh1GQJDYY0nfPOVXpV8i
lZ47seZChbUXwoXjDRuZZ84MeI23x41G2W9q1ljG/aA6EcmKqcz5O+lC2KfX5zJX
1R/+D3QfDTlSfN8P7Ou3YdUkyqnAD3rpfcFjatw3KKzypv+Yn4zuyWtKB+CTo5pp
k2P0qg0hIJ2ior2DK5j6GfsrhzGmrr41VHymYEGZQsW5qGBbzIosuu69D6/K2Hgw
QJWEnp3IhfbY3PxcwRG+01hYjtcuC9Kef71sxVFHDA3gjN0c/7UpGBkASBMfyyaE
cd/1lqtM2OID8RuKRlx/iMy6SGgLrkQMCYfCJbqqBsZcSXDDyhp2/5pEU3cOapJU
yFQFj89I+aY9NC/VvxyVRb0Jz5ZjlxG+SGurIELZgue8Om8Gat16wYl8hvORBmCl
DGX5/sr59xPHMAU/3KENPL3hXwEh19obzau0FoinIeUe126QWSCiBQETmdymE7if
xTqNTvFZOuIblnaeI+gP8KSa5GDFdXjP8LmSInO46nvGUtt5LlVeDXZY0T3DKJr/
/u3Cu/puXDNWXo1ToQy3Wvi2q2/Jjf6bKY9AZ4Lcdlexdq7aJ3DdEf0oTxoJoCnU
RYyxPejiAKr2KiWgXDfY7Xbxp5AcZP/QQf5GUCf8yiUcw/sJ4kiA3fHpfUIk/rQi
922BedfKKBtkEImFUbUxxIooWru6/uOyRM/hv6wGxboMrZbB8C70LtbPbBecqp4A
+leri4eQ3b4wohtlkYbOrluBFyMY4D4fqBwZaLQczuwvgSZO7O6veY7JXMSGFcz7
1waLR+s6CE9kLoSAp61qtt0ZmnWYX/HauK0YvT30kYshv2d+Xd4HyRBYGzZlWyax
WYY5eIF955EVT3qPmKaxjvxFGhT+JTzEZXQIug945bK9ItcDiViIF4hOUkUqe3cC
EUcnNxdWiULjHg0kL5Lyt28ioxR6MVSJU4RXY59HxFubU/nQ5TubdBT+CvbM0jKD
wWupCpL5611HjChKWs1fOchLqD1rKzYRNFtmmrYGKiXTNdTuTyk2qGORMuY7Dqgg
QG0YWYOfPu6S97fLo3LDiMKAI7d6RMpAIOtX0rU17TOYmAYvIPHZd2aEuv40THcn
YSeH2rygDIDlK5ryzI61JApsyMlQwzVon06NfsfNFvGSlvgAGOp4SGqFL6B5Bg6u
5YMIJgsjLysAATvHPl7QUY+kry06ozi5tP7KA9mtaYSPOy037n9IsB+TUtdEKfSF
xCy3b8eSwgcuyWs6VADVnHifw5qu6zIKbYZXNkmoKLex5WYZDl40Cv/d1lhAmByq
G0kn7OycwBzUepWvS/JpNmd+pCsOaSv0CiKiENjNcpEJOPzsSaRtvyf3x2X4XRAj
RzzziM7obsPrdLOs/OKfGocNaytCA/PjI1XXL5JUPMyJpbXvm4fag41nci3BJ3jg
w35qmo+lgn54jB8tvDZt1Viq5MHsGDd1Vu0ZlaHr9MRq1VhYQfHqonTiqyQlMRXn
0CJF12sDzJnBVkQtca/muE+k5Pg54I13akCNtzYQS2psYb+1Cr647bTff4YttGvz
w9Pe6FogU/0mApFK3L06UbRI8dEXWJnkQh/3sv7rDjh7i2Wuvf+Qre9bpptjs0oQ
KoL98QipHpq54KfJR+ZJbz9Ap2q589Umc8P0rPWDyXppgFCHIEhDBcJsUl9v9H7s
Wpsrs+Tsxvjk05XgdMxvGlMCHveKxv/pOeDPitsqVldrej4HU6apQJJ2jvxqWCeW
5LMug9aweIiSylHc0s+LzrQtAYT1QczTYQUSNL1vcYm8h6+fY1URuriv2DtDCHQE
uBRcy+Wno+NQJXPaSn60yaw2NIgkvNhyzt0Wp53e/rfAN49BwjYeeVchahylZ0Dw
SrSw3D/mOErQGoAn/GZcmIBOK+mLsqft7cE2RcMFebZiOCPjBD/C7/A1o7JXetJ7
6t03wQRIVRYMa/Q63vv5140gfP5uMn1i+w/RYU9Zx8wCQUm8Kzb2/w8dE0o/PPDf
Ls92T3Adz3hz1hI1TwHDyhF2H6ItzfjMJ5KiTEpobJsltvcEp4Bg9fcJeYXZpEec
8EAH5rUJXXWppPP0WKli7t/OLzL+BRiWAqR9Lzr9/lkPhdPMj0yDRNBg02H3YJ/z
N3Bf3+Pf36SVXN7QQz1xvPT87j4e6CP/u6gCfnaKF/ZGciBjB2B+LVzP+kcTDaz8
iheHIw8TbazVK/ujfERiTRVokL1wJOibsavRoNhqVQLpPHKa1sMPCS3cF7LjNnoc
FqAZ4t2vrMD8pvX1jBN+vfrCxavb+9sKBUmf/opRa/ztc/KJ2PQaiuKY8LUWFS0H
yhBi2yege8f8iIlIADSBa9qpCTkS0JLg5OwocQMGfGlvc0pPhimGPmpGhiTl7gOo
GvGBBTFh3HEJpI4xPiypVLtB1Xwm33Wsn2dzM0sgtE1QoGTg1II581yflCgsA0me
m+JtLeYxblwAbxIixAbzUbVoAIWx9yGKQRDHiSIdwm3o2Z62DSs7ieL+vUdNmhnZ
qiszuEIqnsunxGVSIjIBaLheehQBQsBfi0tXVNf9SeHKeb/0LKgcRlHI4kiVNhOw
7wXOIkYSs6HYyxUG3HSsoaKvTI5PhOJd40TLzbsx6r0bhGW9VwACELI4Vec8P3rR
Fygbnus5wbFjm+BEz1dNVGb/9wmzHCLR6qiaKIgobnv7k9Pmf7+i/ooETq4aNbaX
3i57J3NHVqe6gHqMbnA4s0KUrH03c2exbZRINekZqDE7b45+yJkf9pQEUQoJru4h
3Ird1nbjtCf30os4zcx7gtx6pgcq9d02IsEwVmW08MBpOMol2Qa2BJ5bqBR0T7Ya
zM1SJ1Hjwh8J9sZl0w1txVdrQvLe9omlVzYHRGQkWYqEn2Fw+jAntzKyoX76CbVV
VRLRV7s6Am699kGGNr1tvgDiLmwmtTEgz/q3BjXtOdZKbnMfLXl46n7rncC7L5c3
wWeoW2gNf20m5I5whIYe0jF6s9/JjX3Gn5unVUGyA5QEiQmreTITUser2RNcj6/b
2+BE/+Puq7gEBY8LOfADZdwGsVn41V3y/6QWdcBCmRq9pQiM272KnU3+F6gS/XzH
V1o0ggG096l3xvuEUdWOgpN/RizHjmYyYUJ+O7ueJ4RquXbXZPaizBoeXJW7/Sfj
ZX7ZNT2BQZAqTQWI52OfmW3PBKIyvkoCgEXaSlh3c2tKGxMlmVBWGdQP8co/I5JS
c44OThiqeggQziykYSfaN21ifXePw1QwKl9rsSV8loFxX0OfXR65YXtA5nJ+G/n+
czrF6GCBclc3gOQORCXMlBXZrtbJ34yqLd927MVNaajsatfSFdMV72bUYE9QRe89
m06DtT0rfI3YTa8vuGp8e0guwvZMRWu7HYJkqQkcXadKcrrrvZF5lTFX3uiO3HRA
6JqnP5zk9xZzq1Hue2MvUB6/wnl8NM/rhuReN2xG3nWnrlwHpf1SZRC8j7/rUZvQ
OaaMwwRGCJfd0wsrRrWSC3bnrK0xqiHSefWaxNKnJdFzDR3F097a4GYYsB7Y3Yx2
FGcc9bkoft+Fgp88dAjq31lcx7f6kdfFuPvlgDEjeIIvlTThbpwqT0RhB7EvDVAO
fxob/0yXqqkTkq6M51uxPj11aeYkw7DQESzysKnDQx/kZcxTbGcjWb6WenaoftzR
+bMuth/L+A7Ee1QsY3Zz7DvwFIB02XmAmmp2slW7QA5q7BI/EtCb7RXys73c3LH3
37kS/ZhqgHlBXZPPwGdJkD23gtUANSSgrqf3iYy1vzM9MPDima/IlF3M5gWoyL7y
oPu9FQjKIx/MFmwZEgLjRoj/ro0CJoVnODaFXsI6wzdidc0F85v50cOifkX7L/p/
qr0gns17j/BXBMbdkCSHX0BBkfFBwDFZUa/vHW8HTd7plxSd3zVSDtf61Q1pk5EJ
U/RR9u8g477/F0J14qFLXBFPO8x5d9ahCsVUDEbtPGnkcIE5L+lq8xIjxmLLsv+e
1NWNA5CqSVBQmhrDcNqePaZW64JTCjRt9hBXZsrfLPRQN1RVNFlHW434DpKXN0nK
Gzw5LNit97OBBNYlZNVryb2wxQ40m763PFH/gfN5Uw42h3FH/hpgHMBuCUUKNY6c
W+Kt7bWUHWKMItnQjoYcoreKNJDusVhFaQNXn4th8RuVKV4qcaKQZgltmTU86rpe
noZ8EPd430rpHFRKCjMsukkmW8WqBGaqeY1tjeDOzFWfKbuSalLqOapKUDj6LVvO
vGYqMki+Evx+WXvVCZUaPOOVFxaqG6CPT1DTgJzGJmAac03WoDR8MozMK1bDkLbD
Cv7sbnqXX3IIdpXpCZuotybEVYGMmqT4S1iT+9BMbQbpUm2zv3s0nGw6ezrlpGx6
Qoc9T+qdj8TFJUeSPQBMLIMCl3eGbKVooaKdXNv7kIBYPHQlWgI9XsWdOyR/8NSL
iipl1hfm8gPPC8kM+6BjMIn4ZjPyriCKwWxwDmh1DpsLbHcAAX2HfWYYbAbtjsnx
UR5nzB/oF/aTIVH3eGEiKAQYdv2bUKzgztOMYDmRU0angilvy1MkOyNkZfbMT41C
ApaNszfPEVEmbNJ4ZpqPvEE+hRACIIurYmbIxX2IAYJYUMJyBgAMhVpzBmPqu6JP
nYvCl0n98684i3/HkZ5EgXkN8Rg7m0gm/0uPHGRrWkEdBLtD9XO22siGsFcideZY
ZX8aHSCd05xm1ZQ9+JTdb6fpgQyqmsApPNpeCmGVOK0CT+aSRFOfr2Zn1kfWSIun
3jWkBluzXyAu7Nv8REglC4rq22to8cDAfKmQCSiIBM2zdNznGFM68QuOGB/dI1pR
9QRrEKEw2gLcr6b9s8n9ClYyhL6yytrWwAp/g7/Oq+9vOx6xrqTJel7P1daAT6zo
TXO4RTIqz4cTUzdkEiOmXLhSRUOaEEMQjRCLKRJm9gzWnsoAuu4JvYZZKcxJ/kor
aubL/jr2fvsZYDIvqQg8jiS08VuPH7XN6O3PNdrpBIP5mvIT1lsh3ykulbJvWed/
ELf+vKA1rLOR0qiV/00x+b1SSufnXP7B4EACOQ04Co0zT0tUAY94QRhCxi4TF4X7
kECdc0aLdeypBW10Vaw99XztoWXHxH3A1oqxUOr5OtByEqXMxPefgChfTZOht01K
AXDI9RUZZNCAWQ4KOKMdrBR4czxkDi3kBzdAoT/I1aXyk7wrjWzzO7WBCen0w5yS
9VwM6hiyZhYFfcpJlmS0VwL3El9S8oPYPh1w7PMolf2dUTSENL9x0wXR6WK4E88O
u874e8SShHJu63WGkQhibX0Z/CXFXWDgP/wshqb2Acyd9yV1ocfCCaENiX3lXsM4
Zg69BNBgaUY3whES1eavPg7nwrciLa7IG6yyuu4oPs+6bHqce4OHZV7vGub9oSi0
XqeCCxn9MWK1wKMNAoIJzwySiCn7d0haYR2670vyDuy1VsD0qiBN2dzy7k3KehoM
mpQ1JbveXoBEulmkHdiUl2libOYDVpdWpbr4Lf4pYRqIOYOgRtxTn14lErja093X
R7KXSa/0cmNc9p8Ht2JlxhWhdJ6MZViPoqk8bhAntwmRBU3BPP5dhxuJYZyCgAKQ
6lGh69renXSOuhYE8pvnj3MjsxdcxxSkZYOd0/nHeAoJKf3O295BcdZaE0UeEZon
kTbV+4HmniFIdzaJ1PsEEgZxDlEccq4Jd5RGKmXxvnPA9J7ouconh70Oasko7RbW
/waxK7nADEwg5GyO9itazggjDuJuNsE4Rd0cIXXD/bpzNp3o+oDkr2WGeRc8ZOeq
EeYa4/YXaHSABMg2jwr8WsnW9+pS9UqXo/BkrkMtnbxvyOtMeTY9vY/34iqMwJLR
tOmbRE3ONumzRZYrRGOm5111bqeb4fg0cVej7W8DhyTpTJDrDV0AyUUkfEemZuPa
s8wpvipAMZQuQCtJT0hBrCj0cQlUdSP6g0rZ56MOOmj6Ef86gaFO2SgZd1wDrg/J
kzXAOF7zGZL7DkME9sF5w8m/Z+miV7OZJm0SkjiIdXa0KdiMdCjr9RYV7zO8MmJj
50/PiCA0fRrhOktIaQ3uNFW3Gp+3ozIwNXMYyY6n8mH0UZI8eBAgwPoKh2u2/36f
kWQpc524WU5zT66t9nlJIj7mqtjqDj5p9QDi9O8oRngg2raKFEQMo4e5YqHlkX/H
AIDtkemZuqoA0vCjJa3khL5Slq9kV/kfPUBZbOp4eI81tmW/U87St8vosnx8oSvQ
reOHXX3yDj7muJ9/AzPuUHyIVY4Rs11kU9WYfCkCam61WxhaJI5O2eldKEWO0H3s
lGZvlMCgug7SmjkSZa3qmNWHgNzx6KdELdgoUav7hS1DBUNrSDATxBI8akHYG5q7
JDcP8g3y99akJElPuvjXdBYYvjOx1QPpugGfRR7POqCnAs2sr+NBuyWL9II1HgSb
wDLud9R21eQ6QLMS9ZLtq6Vj/70tWpFayjCYYXdN0yNq5ZINjypBlFSRNuzspLbf
Hp8Z7aAqEpeGX3tpFgJBURvzqCf9tZYbu0zOxYKC4PcROsaTu5ZDYZBuO29eOHic
zKqWGCkmwKUXsHZzutF9+rZkg9yp7PUM4G/u18PRDsaOKfb0je8f5tHbqDj7XpVv
F5CrAgZJScRb4U1auvkWG4OILyPx7h8zFHFo52Z4f+m4K0cC2x2I10oX7gZ1mjmX
cOIP44bbuiTlas6ghScn2LrI/mFhFg8ivdHlRTQWYC4jnt3aUY5MGXMB9nuZUZhh
6jIiyKOUZDxvfWUZk57kY3YXtQFwxlss/PD8UzxqRYb66PdceP6rgMFxm7bUbnI3
Wk2EZD3hUL6gGZNPtagTyYj9EaGgllr6c5qqGlXVgSy0N7EO1o0Fb06NnhAxGcZS
cXtT+j6HhTrbvx41WZ1vLuB6dGfNWhttf7wI0W6QYTgN8yocQDOPuRpJ4LElp4eA
CR9JGMhNbN13O1Yr6SHLwsNG/gZ0+ToB/P5xcLhNx7LM+BKno52oTowqu8Q7tUPK
D7Wh9+yzKLcpl6wszcMNun8tEn6bT/Jeb3b6xVBdRy7uMmV8iqDSalIbTP/dBg9B
DhMoEmDkEgqrctfKyfyPjRbhJehvSOJ7BaH5kmE61O9kJT0TieOMVnKdLB8NK6qc
EPmlkHdOZKdYjt/en86ffBNANrtNeOSG+RSmQ2FzLdM060zCf4kGYexSLsE/7taX
LWe6sqymeme3/m0bqFBNWm58sdaFFexCm8J58btGzASvPaz5E4Ar2YTh0tuhv+FO
sDXh3Zqh8qiF2VK6eVETvbtyfh8pkvMi428x6qoZidYowkdO/z+BmGfpk4uq6jT2
7EcDdMVjxn1UtngVw1NpF5QsJkJ9S7A6eAfmIs8tJfd7AmEP2EYeyEPpCXcb5ue9
a+YAxK+pRtKijWd95KROmLO7EoxUuvR4R/bldoxHWcLh760B1ZTpvS9Ua2auihRq
5fI/AJHSbBz+zr3wwVVq36jtLNtRIfWT9ynL5P0bY7KdjulfvNLOc8Ot3XfgDBAR
I9A+tTZJMeqBLoivJ0SISXlC65VTPdXOaT9wJX0lxysQPZm1gDfWL1TMNmWIHdoR
juFAIZIM6IQJhZ37tTgmX3iSRxuelVCdZq2TnvEda4cqe/AEE8R5yZjY8JwCRhw9
ATvbL1vkgdROZi23eLSvFTd81xOEgly0IQqJ73h1xzkP659eKR2T3Phm7P6oWant
gpcqfYhTO4KSAqGngg7SyNiMkSvDMpfQqmCYUXL5vuhsIMCHBT0KZGo7bUaZd5bc
X74hnrAY4TQ/YukL88p2blUF7MK3EB9DBf+NRgdq96d4iVf/ZsCtBM+uFXHAOrkB
iDu0IBJ8X1ytXkuk20efuArvODxwtsBAVFdMbIKc1tiwJ3OWQkZKN1vifnidGtHM
5ajk2ygY3pIJVTpGwym6PXmxJ/HR4AlJt4bNpAFPlf7utoHyTd+va1K0z2Q2cjOE
pZ1iFfVGn7OM9McYRVTibLQGg8s94w5Sve5GaQPvYBGJyuB+MQoEebDiaXxquGAm
Fh7Tc2we/re+Tp+iLmu/lAtavN8eeSFP2ErSbzrf0orDG2SGELg1/3TvnVMeaQoz
xKKql9k/PImUWpOl0H5sN+9dON9hGCKg37dcWdv652qhq7TYyJVHeFkkIZSewf/N
PcJv3jY3PMDr7JfyN/It1TrXApY7EQQZblr+9pUuZxi5lHSxhos3jgH7x+6vl+aR
6Kf+4jzNHl2FkUuJklGmI9Lshd4TS2KLBUWYu+7LIHzsUSeNMoN9vsZVAgM6ewDt
lG0XcHpwBnFqGBOMpJfk7z6NM9eNnfBn9mVfsU0wfXt4xGR1w6NEtuP0+DKSOEnx
jLEkz/SQhsmSotZMVoHlWLCtGNQ56dr80+4m5n409TUeB0FLSXwTqLSIO9+LkLI9
6nm3CLkoaRtZQnpnw6yWo0MdBPAYaOYUpynlieUDH2dwBxlP/HsRTx6XAgUTaWSW
Kc1+2xWva7ogSpagwEPs+TVmnjCsWY+w7+RYQD1vndj6gwsu64pMAFUnFh+gbYAZ
X2QVcd4GV8RC/gsLja72DlDi0usgCccSH/LAcwoYiS8MAEOJh4oYorV3B4VopUtG
0ibSCCWnvMwKfKWsjaFG2ZzPUoRQN+/IRVqB0lnhRDEeLXPyzc3I5X5LGLN1HzoA
7WOVgVVbueepItxvs9L9bbtysDcWNZBCS0+9/ZrW/4kWBthD3C3Os1i7Fi/gfSfZ
DTAQIH4xxLCMc5IVnbdo/ycu8Lwol2jlA8J9p/mFjCk1k5S+/5DiEAfmVO5sYK5Q
Ry7alSGtRGpy9DDHTDyG/uAeFqCh4n9NW9wfRZ+gDw8DiJz7msDTjNu5MDz7EK8M
cCRhZFoe94gJNJX8zUS+pgQOiJwTiFCwAEnDlBRv9HmLT/lrSwkjiV1ES3i8PXvz
uQSzI4gthkQLxS+UHjARaDc1K34lXfIDRAfd/hbldzzFuEAp0659LewMrKajpKJG
t5GPHZkNzXzk9QzdWTtdI3J2Fydu2GPmPEC4j1JiqePXaBwRqYnPOw59dFXxUp0v
CbiDv4F2TFbB2s1eKw5xwrPJT/zgZj3mFNgOxvghT1gOmVSMnIoEdOtratm/Mp6p
mNGq8YOkBQkh9ZBsNEOLnagJH0kLlDqpwJQb3WAkdwzY0RaxfRNBElZbGlC9OBb2
0wWbjvtVPAxVI3Wrn2a2UhmU44E62694Usz4RvI4YcNsqAO18Hti6ZOTxsxCX0wU
aEZS2WeEaHbj2jMLS9ZWICjFVMr75vD9kicHsSVhAmXGwDhdd/NhlQ+qHP79FENx
K9lysfncEkHjyINpnrs6G31AMpeLbz46xPImXNifYZS8yyLZBtR24LUu6eqVZqbZ
aX6kX3w0v5GFDj7uJqus+RqfeVcxtY4wuGtYzA+Knx1LJAWe/4la15skePJdrrzU
9NuLf6f3jwr+Fyz0fRIn2R7SKhCXCUhw8VqN4eAP4SpMsb6izvwwlL9Vps9BYwWb
A8L+RtqPX13tqSzO9xmIQorekKCieJHHO3Qogv2gT3XJuenGbgO75/CNJniV5dBb
je8f9JJunwYLapLKIOvO1hS4J9oMFIhUKO3OPGlaNe+DeJtb7ltvoENN6cvGu/z2
FUpLnLiht5x7xuiYQ2Awe32iwYbFx6Ol+aeFklw2EuG+miwxQS2TOnTjm+z/Ow84
G6ZtnlevsOEg2oWfTW3nXe8I05dOIbaEH7Q9LtxPkMKOa5TZYSNt5UFurKUzHYjQ
QDtkfhY00zD0lRG8SSCssGT4TAUwrKZ626PO3hs3sCfxABWfmxi91NageoQDTVVQ
735Tr4mznNOTc3P/GnJ0vjumdjaZ3OaV7yuYz7iUVJ7tpvWiZYEohFjGaeny6ub1
S9T9pb6bgbj3G43k/L0D8tm3t7mL4pkPUwxOiJk6rQoIBO6g2pISb7wVFny5z8Uk
KqRKJR+gMLzufYQRNKDqXrKJDWqtFBpysnSvNtIhmv5Ft6+pH1U4+cwYapHzMgig
f8NVZC/4cfjSbXqvSqFMl7Lf3tif/I4kxq4+f6GYmZFDVbxp4LM0Sl+HofouNj3s
+cJXLmS8iuUAuuGU6CVsBHteBW4aWHndG0bZ8fGjQegEta2Idoug9Gkg85YdbFPw
VfAsiB+R6eO2/Dsc7mqniycdJ3jops4em3LSke19YxRfYxHN1UWTxU4/eASVo8Hk
L6KMW65fPyPV6u9nhl0B9kZkcs006vHEy2pU7l8bRw7p/a5eSjkyxzZMYNeJiQT5
7OVqQNS2mujOOnmxIFuH9hpW29HSU8xFfFuJOs/3N6WYcvrNBx3f1Y/mHRJ1a6bk
usySBKy2YBnntC7B+Hx3d5xL73cN2B944TJt/J0VWbnJF1ch3PMiRaYjiGuNfsVQ
Bwct9ZCOm7s7UbuZdq147uIZlDbAb2UGAYZs7K8qki4kwl+5afCa8LN8xqGXbwK8
0J9fD8LP3Rac4WJS+qTjlS08KzepvBeVGu9+WZUOiDZHXIuJ1Et4V4wj+WxlvsNq
w3kLaoaR4mw4azuJNTtE8snXpU+wNql+JPGfHhVrbETgIOAXf6Z3l3tp5t6aLnSQ
RvaiqkcXTN3srjnrnUvd8BxjEcoDoP3khcLquKuSxumahqxsjKxP4bJZieE8CdYr
nFyfKgfrQgm3qsAPqTr8fvqqRZST54Luf4GYPNIWZyS0KBPfhXblSUlue49Ctqwb
SeM7lcIGGTBbFWd56amnx01xAPQmG0Fju4Q7zu/9h0zcaeeUjFKHKMkjyvaVZJAx
oLX0X+1CRMqm3UCyr0a8FG0KZhkrYl/1RG1RyWx5Bsuo6QFO4ntlg+wyM8uEo+Gt
o7TzsdM1w5qfJtLODWZMYPte5Rg4yk8HGIkOlYi7qrCtnhX5Ia42Ruh0zPu7K8s9
7udbbIplsv5AindnGAkJ+ATYkXA7W8MmxqjyZogFm+zrmKXn2v8e0g8TDzMLeuRm
9goNjtxOCf9wjU0ogk4vOGHVaJ7rwEq93Bp/os8EaRvD5JwrblDA3dWm8kX3ZoQn
0NJ54GBm/2YRK6sJuYAaaPbKaQ8/9BU4HGvgH7Lg9+fkiZbgyaamAUFg+2e8Pp8f
keBSBuDtfd1ekT39+EAncmEPooy4KfORGM60SmiQyO2bavyYx15oal+j2Rs4a463
u8+TNINW6Vv4B2+i8v3J1iDFfDKj7hlHZNTRQiOFuadLpvNsUWiJBJGFNb8qehB4
JS6MJVMvgUjmAkFhdNjAHhK+mVeo5moFrUGhd9/LjtAkKiJ080qdzuTjoBhDgvj/
9DoOE8j70qEGWaMtV19WU4ZDmxXC0rjxQ01t7gGXS4OTa38tmrGuj9YyEtG5GB6w
BvN8j0+0rRW1VdpI84mVdVh4EQ6hyfkk7qGrP5IWR1f8So6N+gWYQGxaWsVexv5Y
0RQjibuWa/LRWuVuueTl3d50l/81EvGdNufyiSrRyD33KQlWGMWqLSKMCoUxRRE/
7WnaojsNQaaP4ai5sHXpdODLU83H82CrX+H23/IAg2HIcA5Cm222ki50lGpn4Y9I
5q+tXS9bkPfpCghZ7TB/DUbw+9BwtFpzmkKIw36O866BhJjkQpAfrJXzvnMc5/g4
pg7vVtEOvqniFSzHkgLGnZ3NgjKTD3Zpj8VVJ/va0dCyQ4+iU3iPR7CU6M4MaNZw
45cD4rD/BdQSxOTa5NnVoJ1GMulVI2iTOtmxfexb7HiAsChAqeUy1qPnjtAp2D1D
NWeGlN0350ydjjumAC7z4aZR/HA9xfxlb0uYXcN55Tb3FpLT7WSo34FVOmRPO0e6
yOW+pIzpzfQzGEij+PWWoSj7EVxksuJm1YlHmNoXzriigQkYk3lOnHWm3uWpIdRT
R6mSu802/HVvcCex7tkiFxBt4u9hgCjdb7F4qZA4Sc5opUv6IBeV41sOCtbuzfa7
WEC7NV4aXaIanfHaJJoI2fzpnPJqyFrsZKzIWMepB41SgD1Zi6VaBuTJG70zKf+e
S692h/3lx8A+4PwhWgytvFImLrxE8q4UfXXZ9JIK5cl9nNZMSyLFbnbNJAVc3Udj
TgAxvBvUGxADPBpErFSG9ySLz5Jn0a6n2fcGv/9Ihn3hDPEpThORnxw7MVxSLh9a
0lYHr+0MgCvLs+RPH2zgMlDLq15wnfzjv50r4KzXyyE59+JtozTWlnW+y1eASjHl
e9PV5W1Z+PUawq1hIR+qiq2tdbqkJBzKQFHECEB4iDGWoKBvmgScoJeObQs85FGu
dmKoZohqMyFs5Uo+jiK+7fTYU7O69cei+PMcRvl0WV5JdZmZLcmy5kaMoqbKY26D
DAXyfOBesqnr6MBqpTMxaT/aTIRRvZw3pP01iDVMiVshA2Ft3Ff/Fhx8C2c2sG1q
NAgjO9FRbGiN3FrP7XXK+IPQgMWNOm3Lgb1JvYvy9eE9CM8XoDYom0uYobFQL3Bd
VyRmX7Qfzjm7u1MA8Igaat6zmznYQkMdLdvTQfvL2ISa3XUEtkpn0KkVANum5x3K
HD3RYv+FS3TH8VZEYJHluxkgNnUQAqyhh2AuOiZisEPmoliekg/cCqdmUSVy7KPw
WbHXl9tHZjbqR5FLPBOSzgF4na5vmeRqA0FwtAvdW/e1XXvYRCgphIryCX1XlVWd
6o8o3U+l6hWf2SdYd9iE0eWEG4iGjz8IcxuMZKCqRv0+uGVrpVf+clHio7//n2wt
w5U5M7evOVx0kC59jlhXFfdAUQM9wujajCl2Etpr5dbPHgE473tJF/bxzT+O+0q4
foF8KU2/B7gWTyfsGSFZ95AxKF+D+xsWsXpLbFsEqnEt/RQZ3U6tzntH3AQLRaMv
yX55xhnKmqiRXuFU++5uxt4d0Uq+YPXe1/Xm2dAhMN3lXKGRdRgFM/D7TkkraJLJ
n40vzH8QCoMGuvvvEmwiY3ilVYfyh4e/E0XGmM0KI1uVttBeQl4MApmUEC/55FXw
1Dqam1ASxWeYZLuAoBtPUOPPbL3laq31LqXJIF6Jhs83vmJBOLhatJhqDIdgivAX
Iio6zjsKfgZut4YspSrKaaIzu70GLHWEsmZZ5e0gE83oKe9+wbUrnWILvBox2i8r
zpt8t37iBAu6r1leAT2a0y8l2b7yJRWAIRKBKL/fWcvAhCkkzAYb4ekDXnYBBRBh
a05hOl5jkj4UnFc6bcbE5htx0UJ4oLWDIqs1qYT8299zGNMGpsTdzDc0QDQ5qJKT
R/Fmr41kNwMQPp6HUo5UmW1tRC5Wp+Mc+WrzNN0eqfupZaxnbqIE5OxHke0Wc4f6
Y+oYKEe5nEshzEbFihLCzyIxtRuq8F6ruYq2qvcg9ldSIroIHUVnVTck/d0sX0dP
M87sf5l/Fsa9BOXVBh0zI4Plrgh1HTVi1P7uj9A1ItnFfHy8hljKbQrUDKTBkWVs
oBiSqgO0bjg5hfdzNEWAIeP2QayS759vQqdTJYCd41BSiBDaG/kbdiXia8QfOcgQ
34lxeU8QI/lhmyC48rY5fG6mcg+Rftoi0hUt3RYQ3UkyrSYkRMlA3uVXqWsaSIDi
Nd4AsZoIotdm8Bmj48BH/s6OHT+bK0N7QTqDXZBa9TbPNiIKZjC0Z3HJqII+4GA4
K1toRo17175u2h7vF3IVe7ZoEVqcqtDRJbJWp7k+qrszxTS9MRW2Rd/wT6/UQBdC
cofSCXp97cK1nSPA6d6ih9t9Oww1hmb0lz/xex+erAYSyat1ND120St7+wLqkYbO
DRv10qBEMbblVqzcXro5jEvVxaNAvlipxPXUoOL1WAMTzz5xUzY88ZSDJObqje+k
uxOzUGzpwnUe/dZhtO4xx8fAZI8wdJTdS2HNhgy/9Zacs08XsTs4NBxBVJ3+JDyI
KPjlcSVF/EJKoO7URBr+eNVmsK93v820DmCWhLawbgEHnbibduTRy2coGLDMoilC
UUww6gDpsicfLyfkCsn2HZ3GhAhTBl2fC3D37mO55DHfIk3xi/Mgw0YHbTa7p3yq
ymUnVEdgpWF2A8Q+6zedMlODF0+emFARDYCnCwmXgyMN15yeEfqTxoygxaqaXPPL
bF51s09Y1JhygxPHzRjUlqCWVsJOfbspCqIVauI8oozJoC5zoI57J0q2isEXaW66
r0W3FIEjsMVz8Bqa6QVUWA7P0eJM5SUv7dWCxQHUnF9XJDBku/WHIKX028hOCHje
hyVNHG6z5DzFn3DJTGmQ08RkKlgCwm4l57HE+ulHqp38/CTHdkXFe3bJthUoTF93
TmIKmigbVSDGCROIoZqflK3RiH+GbJ74fr+IzoCPSsKuyH23rBaiLpAciaVBd3oE
x554FUx6sJIc2Ewfq/8/fsCHjX4nhPQxjmIu/rvYNC+yxu9T/sXV6zyzemBeb1qM
CPlcZ9S7PH5cYj5SY4Pe9vJEhXIz5gqF+QFAZNyjWqzspUgCifc7rdIYeoR5V51u
MqyVGh9oo8UH+XYImBXHQcIJCfbpO23V+bHi417Qwd4Z+dhOniFgi5jujxl/Vp9o
M9VLNJokVDmEnhAai5PHvk5o9OufV2voOepSk03gIjedFPhR3gyRg6tritgAx+ud
OTU8qCm5iY1uz3bs80cGZXgWGeX1fl2CMTzq/Ne9vQsyhCH9fqkYMUzgi1gPAPgv
bScazJ2Yyi0JKDGgojaSVKqmWEyO+zebH4mC8kyVVWVLA0FUBE4enN9ZzglJk26f
vxRgI0ra4plK4seMERJDOpTPrZ0pzeMKV/5sq4jlBScj/mNxN1xnry+Pu+lW7EQC
f3gpVIa9R0XQ8j3dwnsC9EbT6ShqkjQfs/m5kmbhKvluymU8P2p9U98CgleQo8qG
jWQ7vzUzVUX4iq/eB8Mb63jYxArQxL1JLHmj4CqOyD9bnBKx1xzbf+BjCDCwZ2jC
PuE7DuUcivV538rMDJaBNerxX6ImG2/Ps+R2A7vSthKX2lvqoaXWgZ4VBaoBcUxA
fwo1sCq857YoL95bCGGeeCTfb9dxhAhQg4+hCDODFTdcwewDSPTrBqjTVtSdMOVC
wjbHRgrr7vdS6EAJFf0V7Ik7Yc3O4XWu3aIkbDaqmtlHPamVgw1c6s9ooswDZ1ao
vERaxwKmWAoAC160j3RBXa9oDHLXlj6jIY0uisvGcDL2yLsQmWAYEu58uxf7PZiY
mCCwGlALEvxZB7QYiwa9cvhRDhyf9YMp21I/aMrsC0JRBlqpxNPjjhE7TX1LXPEP
+Kn7KCJmWB0GF3XNzs8abF5v1m/sp5XUz+rwo5qxicnq1FYiLyCwRQwtID1xrY6c
z61G4GWZDzz+MYKI9eqTomMEj1sdOfv7RVyxquMjl+FNIncR1jFUS0CkUYsFzMOy
T9gPNUlPNmZLSs4n8aiRHXeZ6zJZW+UHIckgErKEw0mU8eKbotV1TSnJuxWrnhzR
TqKS/7IvUxBGxAGM6OXAZyUkKprjoXNHOymJ35/BevnLq537PiYQlyWg2y/GxcF1
nNcXD8l282zPTOtH/OVyZ7fk8gWihKcmQZX1H8gzGJZepcvPjO2OGcdX7UB+Tqs0
Oj1KEGOpvSPfc9weyR+wzSjaWbMYRdKIZCl/jH5ZYoB9k/urFNNi4FJtCUvxzqV7
E59mH/OEoifFkSCyW6Mg/uLDFFIzxWTpGNuqof9dFHvuniP+gXJAxXsRnYDTiAur
aRlT1KO14Hu2Opm8ejZOKpZ4tkPohkCPpHKX2IOVKDWumXU1zUSlqLYCHoi2zW6L
nQwauFyYaNZ75tSiZ/yOKssSQJqqzc7LcRvgOzKTxChdVsYbRYnL9WY7roBghS2N
jKfFnWXlOT4LtGeIuP5V62SUrQMIB0iZldymjXPlPHZso1X4NqGXQIJHTv3+kQ1Y
k/q40Won3u2e44Z/+xcmGrlwMlVv7vXGJy2X0d7jwUfqIe+SRXXd6Lj7CUICPvsP
wkVI3HEz/qd5aKC6Pr0vAxnTh/LkheT1BvuTlNjZU5U5FoheP8Nf03ygh09VNcls
AUfC+ds4hQxBeO/mTzh4W04q5zrh5sJQxTqbtL85pFiaaCydWOqqjJdjCyK2baDN
XRBVD2aYdowzAi1VC6sLZagLFS7skriBhJge2px+0z7mhvIFdSBSZKok7DcgDtO1
L8ySlwJWoR1YpjwJAi0A42cblj7NAaiAzeblU9UIaRfLLd2NKF0oJux3y3yzaKi3
TZz0lXwFdO0M9e8+XOI5tH5nLfNxe/Hyp5VHgZvVmYfyqDCP3ATiiZRjwWcg1hmt
+7iAWolGN4Pq23Wpqw7qra2L1uCb8zsmyuRJH17U/tJpXz2YFSWFOLG5PRq2qqIr
B2R15MTQZZ41WFM//teZ7MWgNJUXLxZjHrTP85yN4QUUZHSw73jIKE6U41GZC8Je
+nzQfX6xQwN31PGvRiRUj6mXehRXOdPIbNLR+5/VWYhd2D3igJXhQ3jVJSCQ5UJE
OHX2zEpoQMa+n1zYBwwg8QCB2xZXZr/yn8Ni8F2BOwglmpwMnOLXMmeS+nlxBfw7
Z2QsVR7il5R0p0rDL4gJ2Z+Cu2Y2xW5XmaJS0rGgqi/p91rLkgiL6MFv2zidMoEL
L5c8DbVAQFBiA/D/RQF5o0EnuigDEw680QA4l1TZGoeMz9YOivOiLe5nVU7FB72e
W9UKEZvqa7x9Vr5hNQu8pKBGtEq4jiS0QZDX6+EicqAjEfSJVyj6je49vSCoXaxO
KpJwmfJNX/1bLtNbHgeHsbhY4xaJA/4sa63uY2EYRE0YHUnsVAeMI6Ui4TVLPGMW
WxqboCcZgGPWiu5pvibaK/12NBJ/jfIrJeHRLQd9J1HVweg335V/zmDosLsMVO8Q
UseSlEMuavFDefYdfoskzMMLvRUaUQcxgnLS5cuY91e4YnkHIPaTFpGyxlI1AgU6
hBNzBtNy3rAU0ChonyMJgQfkoSkzDJrV9MiwRCimBqLvmepCIEXk/RaFeAk+ecmr
4YG2ikzIaF2RE6cXM73KE1QEyKKDW3yWXvPrGU/NngYi4Y98QFksLW1bIsK5jT7O
P9i1Qx18UMPxjVPryLFlxi7KmadrsPHa5JlL3H4/hdRHqDmndmd1LNiZYvq4PWkG
fabObztc4RWXP5y/BSaxtxnh0IlEp8w5Dc+TE/9TN4xjlo0aX4S7qulsjXoBXLxU
ioAomBP9TJDfiyc42YiIR/wBSpozq/WuVcn8RqkbMLDrdbAMjJtbEJ3rRf6hd9J3
8idkCvrighuOrkLEXuCMnUn1bXf9RiSrXjGAm/hWx9mlachxi/d0QJ5jGCHEpjkh
7/TgStsQtvaaSeHEIH1hc8guYFq9J7cFiS/tGXrKhFGU+Bwk0oYkY7kvvy5EDOUU
zQ64DHkZB/tVUbLOa6jJUpih3nKcHt82qi4lAZs8UdgUg9wilIelAjqeL/t0gbV1
RX5hSA7uYeYjcgVmaDaRvbvYKZl6lBZUCEUUcyAqz+cyhQ+EoTWcZ2rPTsJ6nZ57
ukwtMn5KmzDt8V/SMSM2w6Jy6vt7tFeocDI9Db0g7nzP0+G/UQrbMQ3qA4+ephnF
WxRTjIFNACBW8T5soe0IzrOrPpI9wFJ3WTVzBn515ccvH9iGZqS2ssVRMl9vJrZ1
8+cwp06ccQ1JgPmjYLYbzMsk+zalC+CnBydW4qEaxHbVFr3MLLvggx8wsnIc+WG2
0wXfoIPjflnZO3TO9JieHzVmnpYS+7eMPchesuoJ3V0S7hYWQbm2S3BOSu7fgbqm
da8/LnaC6DLj7PDiHiWGJGxKPlA4O6E+MhI1ppEmpR44sEnnCxjdpy7KjH36MUBY
6HL6H/PiGmFKl2P6HvvGJhPE2bJaDFBvvNrT5MWQgfQS+E1LWwSuentTojGcSW8n
t2KiH7WVDTSOhENnvhdBd59JAj9Y+oxraVI57s58c1mLWskxpXztUL4raWBRnh9d
ybegut3zXfNn1tyCt+MHDme67Ic8wpiR1PxinalNWIle9a9RfNyzNN0EuTsKRgov
dEExS4k2C+fAPBNdAzGZbvLPKLJpO355cvQTy6g02HLgC+jjNdAakBcpPy0mXMCe
5P0w42cm6uw6ixAA5QzoppGOZYQxG7hXtZXCxLSEDSU1BZ0xZDkQnaVXsNQpqMpr
Jdrj5FIyNcTbzNJdwt1vLxOCA804yryXaCTXktCr2Ep8Y6OCEiT9YKlC/4ykRz1k
QgVppEUATAIithh9EABlryUnsYeGK57E6Fq1nympKQalAfkxUI47TTqYkuYjRyor
ABOWeIpqczHwNPFt+Cc/iuCqj/wWVC40fAib1O/KrhvQ3dqEpIqzXCa8OmoBKfSt
ZE1FeQmbohbYp+NuRAb5UmsNAMirVSovL4uTrwIal2+e4PlAbvLJ8iazH8wXtMlL
wdJC5vIsLdpApMtnRC4/CwcNvIFPx8EAPgXRa1/FLFg16TJR7M+Hxzdt8O+E1efl
IL1JudncqJ+iqvUq06gQi6bIj00g6+wtmOylrwIU/C+syFKhbm/3IadeqZDjAGDs
3QCQfy4SHCLMHRnHAhx2/YkwoMJLzStNjODveVZOh5z2iq83PjGddRSmeWVYKuUc
gGwXxmPRPIOsEw9atYwCXZ0DcGGtPx95sB2M62jszAPwtEWSR0eiN/sMD5TGd+I6
7VeCnBUtzahslKMD17LORlAvwAt9YOjbDMsbKjMsFLOIlFEFRZNlqyKZZsKJewI1
TlxDEfF70XDQcNwUAkrUhL/pIYe4/7cfAeGP3afxUr3pidgXvWMMuNgzyRMoMvvX
h9Zo8Jrp4+xrWKPKqDjbsorUBu3W14/8rQmvuN0Dc5ZeNVHK0Pab0bgvo7xwJrNX
Ai5/5uLq9UREIlMraDQ8bhi/btghd+BuaiUgT7bIkewqUgJKI/9cgQ1dRXlyNxwi
YVodQMbLgOfSv4IlevWtN79eptd7B0VlUdFYURkhpQbKRXnXIXGC/mkIiCPzfosg
UVWAYb53pBirqzYQfla4HYRC4H4g/tNe3NWih5P9dicIwr+FYr9upzDxQdzY+kzo
UqXXer/jhGR51+uCNS+LJjZANvk4+JE3Va/Ow5tQ4kA1+A/bObnI92QgvnmQHdSj
xFACQX4tlPuQqnO0HI4WvAjbFLEIlzbXNk4gyplXangNP1GO/Im2moG9J1VSbmom
utpuU4ZA3f2U/Qt0a2P2W4WrCDnxrAMey8oDv0LWw6jnBDZQP2rn4dis0YcrLzyF
C7ahwUjMS8xQbm99cSwYwgTvC/y+qLpNaHszR4aSbz1abM/1fRsl35MFzDfXrPJ7
h8j27Jcp9+X0Wu87KcZrApSjAtqP96a9WCUtLODJWYBAqyNFrVWGf8GaeO6silZv
V7MYOw7QLsKALJAtAzIopegZ2bx7cGyB7BBtT4IzgGeSRdTygvfAVWP3ImP1GBDc
LOjAnOvIeT742yFSvQXzUbhDI0IHKDSuoyvIYgEtERGwKXPL8/+BhCpM48wwGeZb
lUyryza3om9kD7+8OuQDEH70g3uoIpdBC5He4GKx3BefM72WBl55nJruSnhR3YxJ
J5LVG3KL91zQ+fERnEB18yFSOfKKD639Y/e83VMV0MseZq1HgTjWzZLOX75YDsvc
VKRLc4jv3xucfjZmBsv6JSw7sKqwjXc5br8HWwQzgKdoSTuBS6ddXHybfrIa4Zcx
eNZBN99XlMtJsgNd1WraO+jhETmR5scwABqYjw2v7HNhHrSKSVpVPS5mowJ2YN8J
DNk5j1o596B6TYw8DPo0w/zfNnHpZaSY2LB1dkjZmAAFwY7vKYXZTi+iyY8j9Eig
fBWWKWIg6VzaU50zqF3ZmM7toQntE6FB4naAVQnGtuOBXucZ++MJxvlw6YceEvUx
EckUmSobngKoxZcxwnKMBIl+r1pQdWxDNclJZRDFK1IE/VNmgpnbEcD275g7/19e
Jn4V5pZplP/AdCVIlpl+IcK9xePfi+hiZ+ZmbeE+ezBzqmetz3igw4qi9CDemXua
jeZVWedE60c3601Rndc9ML2sFjS5S+SCiQgexIOeQb0b7fp6Yul3sutmXztrXQ6c
Xl+z3WjNcWxGi6XYBUhIYFEB6zpw23Ka4ej7Htp48E01QmOXHPbbku7f3iZjuhRA
kwAbjAN2FWlTADoG4vUpAhfIJfa1Y6SGStXKaOzI2UOSp5EjkIAQMM2h4kyyKYs8
8kFS6ObemS1p4h1pReid5qCi55mf0uyb1XmHiSujeI8baKaApw7WysJ0sqQd9dDG
THaRL6DtRm8v0VFiogyUsD/GoDFW/Cc9mtwSuRD1E8c0zzcBcdaZyMZNeC5jRFqs
XHUjNljAvvSPU1Ymi5yDj3lmHGiX1A36PRvcbNqKZX3k+jqO2KOYH8pzhfZJfY80
qMuco7MfqPfQr55rJRwoqGGwmoobceO8M0TlfYHBOjnrwF92cTbVA6x0bEoI+3mO
vWTmGvKFUGosERjbejwlKhIEUC/DIr4XBNacy9j98IgNIsA0IKgy0KpIWtaGzrw1
LbKJDbKyJL2ShxQtT9JxaUQV8Ydnybxqy7r44iEAaLJr3cwuGEyWbVbTo1ViuYoc
OfmxtRPSNenWu9NGMXMgpBWQymjNN0LBLtO2GDdsCnNI5LFicLWj8TgWxNrgYjUW
nU/4Yex40WNQMPiMNuTZ48OE8YDM6EgLjMPiwXp1BiMPvOdKbH4iIB5RRz2xEPfC
Re/ffxWkoUUePjjjpZKU4cPFQ81uMYhBPW8RETkjcPh9RaFIO79d0wrqIYtErICC
YJSiOhd5adzg0VOG5vccAd+yh7GjT0xZk5QeCIg4HWE6ZNmSU1tU2CqVFmKkYvAh
b4GonzXgtgrzHna74AWGfRgH+2M0cklk2LeLJsTFVSbB4TZAJs0RXU4I9n2Snav7
4PfXdUulZBp4oH/QKIafZumc03Ug6VSABqaGs0lLd6HDVNXmj2S1enXWsISW9zyC
b6bWoFCcgGTClB774y3Dg31Zgao2Y1upc5anI8bs+FrgDlRYCtcwbui7Yoq9fU8i
wwhGNtPUImLO4nJjJqBRcPSSXLUVUbHUFNCFktzOXIBcpvfZpmCST1m5bguOseT+
2Pv1xTXi31Ho/8S7H1VQ9yuYZHVg4pMoJf29dYCwR1tvbAjwtORsH/pTn1K/kaCv
ZT6XA+c9UtiRgOt3S92Uhk+5zIr/7x7w5qYKvlGyWKIhj67UzpIgmx1jSXNve+iY
OzmZ54t3r61YKiuTSN2KcdNHHeKLS7DWXI7suPJ0YnvWLrQXQnqEykpdm2V1aPe1
4U3Lu15brJW2yiGrm19c+bqtiCtpODynnQPQXCimM3clGLYzNkbbYutzDf5ldta5
Uz12uLHvNauyoVyjJWuVaNcOuVtSB2O7/5Dr9nI30RUF27UpM+40qTWbQPomzHUA
cTMtxPwVBchu9AdxRKHPwDdbyDJmj1OG2/S9ptuPbzi0PTLH5mZHFDxgOlCtnAHm
nTJHJJv9M+QgTVXFvqW3Z8k8IOauPsS7JOsDVSr9GTEqevhnVCr2ZbGjxHn2xcX6
YkAlXo3BcLNr4DhBTz0tqMai8fMYYdC1EhQe7ONq3rthu5BawgCEc8jGeTawtR+S
Tfdbtaa/Hkp6+5PyZy1cZQNUSo5P2k9DR1WUxl218/Dr9ycy9KuG8XdA2gkP0KQN
EGQu1oAn6f+CBGyt8ADXcnaZOTXgmtIasTf5o3HJjKH8bANdKRVeEDJV+3Nycxw5
41YApF8aAXn7tQZAdD+cCmFbZzGjXP40v+Q4uEgrNsWiTGocG5QAPaZuSsNfLdec
/RN2QOa4Ex3v/uky5K28FSPNo8pLCWXVaOFcSVcMBS9r8Ox/r2ukem5o3L8lhz+H
i25TM8c3w2NUOSIDZN3aMj+sXoky437bn+2BdBDpJi/rVzoAH6A3qEObOamjIt5v
CEtgoZPuE17V8L8j/bLbJqS3xzsiJyTyHH2/rGYofDegETIwP9l+J0Led5kmqsNe
w+UmoZya22b3c9R4YEeruZA/xiKBIikiWaXxsbVkuGpV+DfQEsFutwYeIMBxoQYO
NgopeYfCKrsVgr0T15alQN9Bp7834xUt4uaN3hzI2w7Ml/0BM8G90woZxdHuYb9X
onkVTEq7f0V6PG8Mfn6xAl4QXYTHolwbze9e0WdOSs0sgS2mA8Ftv5mBdOn2Cj1m
zCrUZ18qI5Ug4pnAAmhdxMg0mffvQFcstbZUSlEu06NEn2AQrFFIg/wdF+mTKI3b
QuN+4Fgxz+KLGGgcK3Yy7/y+MWVlZ/Z/cmWqn9nPZuS5uKJ4Q6MCF3xRXwokf2vB
wFGr8c/3MhA+lOkbyUEYvaiwPnRbEXk+QMkrsFqP9KeaBxwq4dGdm8pV8noH9k2s
rXPtthwlIg7CLKiorF6YCdoPZj4ACtO0QZpoVmOZc/BbKBZVM4hj4dYjJAVyGBFQ
72HUgEPidlxgANBoA+UjtOHrEJSs12jPXqIssCneh7JBHwgPINgn73p6z6PkzPMt
bbRVKnk9dF5LhcUWsqCPHW75Npu8tGFABINtCp/u04l8y7zMzWe3DLqXMw3AGneF
pgBHoTvxKqJ2RjWlgjOI01sCq/GZ1KafhCYvHfjYBFWKpa+ZskyFqCNwMiFqFTTK
3pp/5yG1un1ss7+YaFacIQn88J2ZJqoY7F2nllMgSI49XALzkVpTXT1DchqUK2O7
wVn9ZvToBqwTuDMzEJX/pHW6akvXU6EGlRWYlB6E5FohzyMXMEgUcgIgiRZGzHcK
oFveYH/paMEVk5nyg8n1ZQeoKhs3/I1W1DyVjuvb81rqHC+nXTcd48dcrzbiKEmZ
StuDCmZRzUhoRAYQqizhSSlaDnw/ARXl1IdlVi1DU/0f/KpuVrNa7BExzq7U+6S9
6P8lwsCkHVLM2j1fNKEGTiORoMh2dEuVZihjrUxNSFfIGHTBdXSn948L1iZYc5DM
t9P3/PPaIokzjsv1KZMEWSlyLPzgkkBXoTIMzbMDnsX+Oe7BnIZLUX5KOwfcaHi/
s+B6YHAgjBhQ0Hh/sPevlqJ/f4RHvF1OU7blPyGRRsmcRvQKhrKNNTRUPTdEYHWI
sOkLD8GwSMTV6pgFmu1utRHI//C/pFl12bDY7Nu0j7OK8o/b6iPC+EAG/NtAep9K
+rsuYI2Id5lHZo3oquQEhNxjCHAEM88Fxfeydm+yYEN/SuXn4uxtOQVUD0h468a+
LlYJXtYLS/dCTc+uTq7UefyQzjPd/4qMHEgfHetcH62uSfLBzDYWNb6G7Ro/o+hi
ZdbXF/PnxE7Du3tdJDCv9QiYykmd1lvp8WseKA5cGyWR94+XaVoE6j1PN+RTFXXP
aIV+9tc9n/EOv9DLMjpCFCtpUtKJcmDvxNdoH8Z2z9M3UFjEP+yxGBAsSlD417u/
orI8ZJ59ZjaYlfLnHnUTkM7ORgPKLqVTyaI9sp+uULWKDAgshPwAVz/cYkVh3QaH
QM59+06MG5jPap5Nl/misavB7Lc7wnmIRu2aZiOTO0JfBjkpzsuwwXftFjnLmtCd
STxPDcflWk8Toes6ZBYfp0wTsFLSvPg1Zc+dKDUKusfNNyKytd6RDSgUjGCQWF+8
4kDzOE5w2v5RKjguOPeMp+HGFWn7t/XFcM8tdUYvUYFwBh/CdtGM1o6hxcdsUokO
+pJiuxnFSIbW+DYXz08mcG40k8uS15uApqK0GVJUUgJuolaLuTbSMuI4FpVHDcp5
8vqem/IAragMTIMe6CNEwx5/wDQfNZEPE5SPq5xJdD50CYZTMQIcoopxYFYBEG8L
kSsEXMCNtxMbbDqzD+rhlQwREPRLF6uQ5ph4PKppk1uu7qss9wn0ptHkXxOZI/u0
n+3sYlcGb0YzKngAstlL6qM55zxO6sd20SYjy5O883Ghec548atvyZVZpXe9q5AX
2uxn2D6pkwzclKJS4JYyHkKLkjv7gw8t5dSOjUObCaoFTmcPWXdaKIXSS8nN7CZL
OiOIxtfsvLbwSMtn72uu6zkXw9dT9Oxo0SHwty2FYhl26NM1oMrjx+rS4xjLGV4o
nU4eODe6Hkn61/OHd1EIDA+tfXlxVEOfLohId89PsgYtx5ay/Gv4U+56+2ewCBld
cSHrFRB2XRv4wgBUxHtcoPqrtwZqqLLw+yWXPIQc+q5WKjMDaotnOrxssmZzYooO
sOC4IGnmCyODWLJEVFHFXR5f2KcegraUy83XdO2hpE81L9OYCZzp4uA6weec/0nu
7KGAz/aepKcYqKdCnB6X92bJEoTkBLaRH8pEJOAj4lzlNOhzWB+AWGuhoYBmYNsk
Wzz2aX1qoFAvStPAfkDXFBHv76HK0X5i3Iud2S/BtV+wlQjR7PcKq55sPXdoVRyu
e0yjjPlAxrDuNKHq+C7KaR2/CXvRG8Dhva6j5q3lvp5KzPo6Wq0EuOytKnzlZRgL
wYoBRu3H6G39CvLLw7jjC+ZFzIr1BpdryxoWQTP9mCmKTUuEdwHx1OxwJ6oz8/9j
VYdZKO3Utdtefwc4LGdTizq8hF421KIi9hYjz54zaz2w7hzAehKCKaFh6fUIoamF
T+KZF30eZdXy1XtW6l7tiomTJIge1ex5s1BArojtJJnDw75n+4FQJB/4nd152C2A
wHSFbQHmq3dTDXPjX2xTD4oBa5XOO0aBp9qqPtFxmSBqljPXAynnZDxyXHdDrImx
kc6KbCZ3/yFHmsxAdKbzxBeMu4InliJWYQN+bdqbzH4xBJqdoDJIeGwCsj3lJ/+x
nu2U5z7lopgHYHeYH1Ce49mKh4oy5nnplYzCtyInEj7GIX0jLonl8a78KGMMZnVJ
KhMFefeDGKuyvxuZJqG1ioI4Uzck9kX5IyR8uxi/TNtJ8mtC9P2Ps1d5xP0M0TUZ
P0y2X40Njo/gxw4ChqgtM9iszX0HVU/htybBB/3aonkodGKRQjDBWhT/yOJfDgyh
YXyj9MDpC3ys0t5bcxeHZ2rHxREdwewI+qiyFfVYA/jWNEXs24mUYvwYCCMdt8Dj
lkimOPGPgusUtcW/7xxzRY6dO1++WQxKFzr9dUranbzBzW1kEx9UOXxCTS1qeExp
gwjzISA4eDD3qOvx9xOczmMpOI7zb+OLz863iqlSoB/gm6dYy9FAwkkkcyzjUAak
rV7CKMhikRSd0AiR2D20EIC5WEwPe6i3whCOghrFShDHHp3b3Pw0jL3MMJrjYYPl
cWZ1935JPhQ7hOMztYRy9YSyvMTJcjrQtgVUd390C5/ff7hE/m1GjT5V+VFsI2IY
2NLTbwg+4sTGWK0+Q5l/z7d0iApgZCzi1rPjpeM2fVt4Wlc6YA+HZM7vGZC43G15
MAM3/xOsQkrhR3Iwwj37cNC/cB88Wnj74EIoi8p5AGoQeATN72se2qGhR6z6oOXz
9kyORwluDYdrtzlCstGtlMJopHp/J6ClTfau050oCZUvmDTxy/ifEUkStVIv3Zrm
wHZMjoz6wc1V703snm6IvkmGKuMi/YnVsYGYnkndw/Dp3vGkDpZWjDd8fLb6vxrG
gPKxSY58oyabPC9wAGLLPnA/5XwvfI+QRmmiRnVh65GxgEPPTVzsYcwxr5Ovo1b3
9Uuvc2ZUCkez2cWirDSZQep7aU22SqqxoYayeHxXEkYuUIeNhnX9JTp03yP656Bf
LOUetjty8sxXa1GnC7AQpeG7k6G/nAJwnSnACPwlfV6VjnvwLJhesWRqJxnn/SBa
3cds9fuNF3zGeh1gQIHJH43vtN/48HN4sO2TFKNcww3NTvBVIjT7+PugmcxBdEka
4DbfeSD5eEFIBVxWGjOMH/cdhqNdrczqV7c20E4UibbStJa7pZvFDJZ8w42i8wF1
0QoH4n7yOCE7rEbOdrg4afTOVJfc6U7ICmG6WJ+c1b+OyUW3cQRphrT9rDAMIC5g
y1AjiuUiOLs+JIvj1KiR9pK5ReGMnUKhihSlpxD+WZBFt9U9DphHKDdJzANA56wL
Z7Y/jYU8kL2Rs7U5KYbmZ3vX5g7+PWqUbFOB7n3t+7Gq+Pk3XXb34OdsbaGoOm7w
zCa/1iqIdihKrNtoG3G4okDyCMnqDx99XymhYDrjKZzP9KyyjAj7ej8lVx+QMgmj
oOjWcwv0PTeT7zJ2kSbOgLcNagN50LY2KzqdSmITfEWrZ2w1DnxENIEObjW4SuYP
e08hG7xl7VhcBalt+14mMXQxFxKw3uB9Os/SVnOLvk1tCG/ljsASmPqbt5BzWRyZ
yqtbfj77DzIXPTbuvmQcJrol7edA7wW2A2tTQiUrBSGQJ0lX5jczrm4NRo7KJRqI
XOcNFueog9SpaPAyMCn1JG6SWDUprSYbSLtFsLosbdfLncUTNsEyngGnqi92A90S
GvPb62fxhLfET3SYBeFpiYvUpsoZaXQN9bafxlqWEdQZF8oM3v69MThS6eM7mUKv
TZ5sMc+mWm1JTwcsqKFEyZJbWUQcsl07CFPOwZekX4+jwfxoSoA9v73apcYUTPbK
555eEKA3cfZnsOF/tQb6neFyme667XFSNmVkg4dBaWzXhyiGpjSbCeMj3Pkf1K+F
YO4yhnV0fPdSueZiuFTEONMQdZYs5bHCeFpTvhFcNyOa6wzH4ENiGNdNMooPwAEp
qzqGJe8g8G1Y7RlFP/e7pcBSvu07S9UTHr2dWt9O3AfOoI9O/JX2mM7QKDnNXICu
IGbKD+C28yywZVqf26BMN5aYxWz1IP4dBmZTD2bGn8emVq5xzD1Gwu/F8JMbHunm
KcqGlQk0Co87SFIQVcDDgHxEMKrVWOCw3+yUm3SLxutWVP4/9F7++TLaD8H6Q2cS
sKI4wZpssxEk9tBUdL5XQk0YD56vQD0Q/J3vVDhjXqbfTjytBRLvE7TrGr1XPRXK
xX20pH1zS/A3vReGVs3kBzqowpCOVphK5LCc8VHojzjnXenlkNxFfN5qnjxoBlu6
F0iSQ7HBbUHmcj0joI5b+FxSOh1SvZQf/3qARQQA695svQ1MzGWyrHTgo32DrNHF
qLamSr/CzUrukAvB3DuGCQp36WWPbCiPzjPtsK7DSc4GzDDkXxPAaXO1eu+QenCH
KQ7Q9479eoBNK+dpaP400xvtAkhx0fQM+xSgGepTZ7rTEzulESg/RmjPzMhCWBwB
KRxtDCsrt3Yil8G6jNR2SjOwv52IWj2SrMaedIFpRbkLvaDyuIaCQILQjBfTjIVr
VTFIkV3UDpMm1hG8bHqyZjT/9Ynt4RH7FUV5GXJhGeNOXQ8mzuVyBSuY6Yw7nI29
hsBmm1w4qNcYBV1WdPecWxrhByQuL8jnNATf5kq3ZIqvZJqdL8Sa4NKzUGfjiMrF
BPyTHd4IQwORqwtUWCuhyRPTkKti7/JUA1KiVORc8xRRDbwM0WVxF+iUZk8rW/gn
3Vc/7RWF855yvOjaHVFEssFm9ITlWBOdGYFgAFmzztauST1YaT2bpzwCynnYSxsO
nhZDIEZyFVebjctM5Sn0Ho2XBU69ue5UpfDCE7yQ+Ooe8CTNkyixAZpn0MWO6pdY
FVyhbDvPSYNjyz2rBxD8AAr74rr/bbsRdiERj6qACJj1gID1Zd9UId1zZUJ2G2el
ZGrXYOpLZMtVYD53F44cEqzQVbsa86zyfKPzFrGsId0pSZm49gTVszl3zocWUxEZ
br2BGOFvDtMzzOJXnMg2n9zSX5xN0V265UhoqiGNAoS45/1lXqSb528QsQXLsKlA
mqYqFC+SYv9PhACn3B0zeNcKuXjdwiUC+Ovr42ISeDiIGqQ25bqHbteejFX/oHoO
gA/nd2E21WI2gTeatLItgth0vFOK46kKG93L8uM7zNHQq8tj9/2G1XbRi2h5qL3r
GmyUo453fKBTGoOxetlaS1I5g3nSKowsjO4cNK73FoXY0Ki0RB/tFXGZU+jNBR+a
Km/JjtERKaaAyvPEoG1MR0IWMT8E+7fN6FePx0tmrVBfaHGK6npoE0WzY4I2evgU
U8h+qXHmOnuFS+VhCPYsXoZM+zYH7pKrTFnukrnD01nvIrHmumgNz4sZiCPhjrQZ
wGP7DwxJREYXrdXSTJ4ODoA0VFl1rBZzGbe3msKIEcSUNUlHKOZJ+rjovq8e0ZuO
QN/X2h+Dko4zb+I0ebz84X9K7lruo41W5Rh+7V5dJm4rn47y9FLqzdsZpu+JqWc9
NK9afWMAz68JfZlUpHStoj6JgEPhSntIECP0bv+406dsbbW+WWVBe39Qdg8lrcqN
jx2PmOR1Om2Q5cR9+gDkmax/4tM2ImqC0erFYjDFx+dFGJRdl/4yB0oRjtnFgsPl
MR7fAC0upTCDKN4AXPXXz8U8CxmmUrUgLM9rxVMbbvumBSbhZ3PpIts//G8xA2jC
R9IWZB+y/OhNioZZKun0ytALXyXBURFAR5k2ffWLwh/MFJj60kkKcc9AiM7CShgv
h0k7drJimQXJIu98fHtd7uXeF4KKBUvN1DJL5Z3KaunazYAvP27ztZJyfqE6x+fS
bV2LaigHTyVpkxPehyIVO9xsEn1xK09G2wXapt3EC0T27TZP9T6jrIFTIYVzgz27
2UTE287wiC2szGEuCkoXiqaz3OSQC067y3E43cMW02zcfK9aD8m75WAWENRocM+c
urQy0Vh477k+nWwQgomSL9VxCYSGqj8fzGbmqsMzF9qBhlMrrS2HtEhqpzIUsJBY
/0cVG/z5IsQ4UXqBIe2SEw2H72UCX7mw4D9Dh7pOMLn6i1Bo/uRdHOGpOkUG8qPt
epOycSDkccXT5HFeVChJIl45kimrCI0J3x1UVJIfJQPPyZmPeIa5GaZJc68gmrxw
rTKqhHtmh1ZHqxwu1mdvVP5SB0eC2Npypv+M6Z30lQNEkxJIdkFpi262S/FBW3o4
xMqCtYvACJ0aL5vpk5t0RjWQpRLbOh3Ds2ZXb9WaNnhrNEQ0IZ3e5ehqNtf83Blg
L4plFOLe60fIAW1JCQ2tVDodiUjAk/whOZMXy+at8QPXP8oH4dw/p7wT2l38/Tly
5Rxv+6bsxIbX0W8wbk4l7eo3vt6oWOdpoxyZMErdejJnI4BNLv0f+1Hk6vikolhh
Y5uP2R+r09TMxjG4lXVpTGgSC44YmAAFfgbZT4ju5PyuYH1XeGdGpD/TlSbvk+h/
hSv6gN1WtOZ7SM6/4gvN3OprtVIIFBuli2IEMJ0W7JGwGnkOzuVj/HKpH5fssoFT
oPJ5JJsVehr3Nq5StDeGwcNCUx8lxXifGq8YlRCH6ZgQ7fliVpLO91CCfn2YCuj/
2O8ca+NuS8LFppkvdVvyoeqWwMROY4X5mpFDZ84tkjnsZLSBtVmP7PIoT9OcGMbq
xN4AtsgA0UJYvd24SMHc86cHkjqQ4X1uHAWsuOg61FYtF6wq5IR8symoFx7Q3rTq
tDsX+RS5Uuah+GhswRRCDWjLwzIIHlfMt28HbRAR/quAaXTw8B/OXrchNoF1Ce7H
1ye7bpkyp/iEm5aIOUl0JMZlcGbh1cszzziDjAtSfU3nd3KOiugEILKe9VIypQQ6
aBMxffmsyKN+hqHY28qslvqukIBxbBjFhmfH2k33GUNPn0XI0qoDnWgjlKHqgrz+
lcrA0wtZSSWFHUESwi6VUerT/pf6KW1OMVH7LfI3piETQpGiAyUTSx79xkbX+ecG
ihuAbLY0YFEIuXmW/oyQU09CQ5EJSk+m3xge70s1ao8n1hacds3YyQ5QcYUlakg9
VEcdhJ07Be26fWzzKE9plZXOv8NZzhon+230idN2WAfmQC+2ujXyJtRRCnCH45eM
uoOrlm1nWN0/jyhi2VqYKi4dISldSDt/rVHGiYp3ytX9UfmZDxazl6FBa+thRSv0
HmgugZUBNe1Ycubg96hrxDuJELQ3on5LPEhQMwkXRZezr9GcVj8BwfheGQE3yIYl
e6u/s1xdSoD3k+8sjpCO7kbEab0K9ZHsevVt8XitvY03jX58oC7b2/BUZ1GIlS1v
PR0un4xZeCvRKeYnQbJDJAgsVr1XDE8vTGYb3aOV0taXg53r3/SakXNUAhJvVXbf
o6RdpxeiqJvAxDVATijKwv9pMLxo3jJGXKEOFhCpFT7e4WmtXgbdzw+qcHOHjG3p
wOaAOfNiQwE08h3zVi39KOsUPNDbEM/jdTnpkIcuvcyxYuQmNxAAXSOaG6bYz/aD
geyRPsE/bjAPZQTBaow5R31fI9eFHHfIgNAoSvldP20vLF/BLT25Rn07b+qIgdLh
llySDKhDQeuO0wIXFkOhmhlmwK70Nl/+CmEdGnpQNxkLSkbVrIdravwU86ZOO1j0
/sFKBaYtMiQa38B1VALB3I8Jvv56MTdHHoToKZb3HHzLtazj1+0UWS66EAGqc3Yv
j7x6NY5evprruoWLAqUJvGYzedI6KIKzmAkVFUQswCBDg6aBcpR9zA5nlvtViRnw
I3zLs2DcbFjS0C/ME7S9wW3aVURRLu4Uz+CD6drxBzwJhx2rpBow4PEFf0c4Ck9x
ZeZhy3uIqDH0xPAIFF2EKGrjs7YX9PMNUr1IeEQ0snouLBsWRwEtHQnGeiTj1TXe
uMI34B4JXHY2x3784EA0h5gh4ZvqOE3crDL2uXK5DqppE9ruHjkqpz6s/lI67MRQ
rAGuA6tgkiMnQ8b23ynevS5181lKCyjaXI/4HdYWX33W0x8N1O0EChWc2SX/o/iM
nHhH5pnlaR1ksqUGLBVIHf4Lap33GDFKe/JFELWQUxXnR0q5TkB9JrUYteSxGfj/
IK01kRQ/3gHklIHrRGzX6PWsuDkb6BoB1XAn0t6e9bj/by0wC1+4Kdq+v9l3lPOR
X4HLc63m/+lRSYjQwx1L8R/S6LDKd0dJdAsm5LSl4+X8pxILIAZcCBpFPbbpf6vS
SQE/GYxNEc2Iw/Z7RKrRvPuKtjKTD4jAE5fxFO2iFwjeUZJLyhnY5HoydNtDLg6I
1CFKjVQpGreg4VbZ7cYGQ2IfWR9yfMvd29RuVAmyZOrXFHAFjZkOAr+Ayq/shljW
EUYNxkzIqMPSdGTczdw8IyJL8NKw1AGubrMFWn8r8yNSgaHGU2DontvT9NtFgv2/
/UjkIUDXEPYNEyX9WrwkLd2NS5542UVZ2xTd8FsjYUnn4DuJX5AJ9AYrot8qFddg
cm648zb3uHn4FDxpSx/+ZT+jEdUykBvGrscpXw6gTxqvrUEJ29QMxQe7ZVEOy9q5
N+hDdCrVPNdmE2SypYrqr74V37PzorZzvuwa1BCwNHV97MaX7DIDgMNv1qIFqS7N
wb+4Yido41/T1BCKYwXxe2RiXIinXQSBX521X49/30IOEW8HcGLdpC6jLmPofayx
C76GyKunFPfISWRGAfFeQgd557XTrYeOScF1oyfllAxsKz/mP9zawtPUfgXyzNK9
TDPR5YB02uDk/T3ye7A4rlpBVyKT3u8YizJxQKz4ZP1aaY11aBulqKB5wUuwQEhV
Iq6iS51FncjCix8o4urRoUM6lfcSXE4VMdWRTIV8p4a24thpWFlXl9yfbDLE5FQA
UNkMkU9+8eDdy8OX0krV70NwuNnwH2PXkTf1icLj27UPszuC3rINoLo9Sw5QJo74
C/G16ikHv0RqIrVqPyQzNilF65RsYW0ptOBDwDTbIhje38brxLk40J1qZBHtcTsC
UbAOiEXiJmlUrQWSfdTjNxfiyND+e8/QSUihcaSljGCf2wNUN5IqjKZ3l53rUIeB
MwQ7RScwQT891vxrokEw6j8nMw8+hSSm7qUt13EvM1J9lamCa7vFb0Q7rnW5Y9Pf
WZs67ltX0MEk4K4LHzr9QKyf4zqOZ2PhyNXgqMIRadBIIT8KsrILgr7E85Nda6wk
n8bVDsvsB0hDWzVpBaPP/uw1FVtk7gUUnnvJXBqKVh9COlg1+kRWakKiA/b0WoMN
rnxOMCrSG7zXJwnmR73npcbcoN9bV/BZYoXoA5zsIkIzvV3PHi9OepubNhECeiM7
v/NDZjf8no/JS4agMoWvsc8PZ/T2eSzUtsiKqqTAh3bjvSXoLrysCXyKVz19OSWO
n3AtvppxaL2Wso71oSvbZoft4Ovd/TCyg8S5ainZazeosKv0det8skGqToStSEKt
TItsiEvFRgOcAY8c+CMhzU3zcQM5u97uM1+JxZ21YF9QxK3AkeG3fVAwneH20nK1
wfbNIurzlcjAtiTpNsPrML68TVMxa+1YAlZTbNgDeRi59V6LPbwmjMLtvtQnVIxI
t4Bqgmd96cRGmU2MUiyL+NllXAfCbN6POaDnFc4ZjNA3wYWPEIAwWn+AqzMxEoPk
VVps5cKamnVFDAtORTmRbvtmd0sGUSfUMpzZcpXVCg4wCHOSitzvMHjrQZA77yNx
LapyWA5Rokw0i6qzIydnoigNiepz/wkVpR0T2Lua1f+4zibaBe1FrKr/Lsttahw1
HUvQjj9cRTQ5bEhxF8xalaWZiZsgJek+2IpGseRuWrkH5QcyfzjQ4SuFD7j/TMvJ
/yuXFvPJDK5yGPFbixMFNhLUWE4Zc4CIpUouReZCdqSTJd+ORkbDj1I84mVurldA
9HAUxjkD2vXxXYPZ5CLD1I8vUFNhh8OO977c9F5E4Hfv1z2b0YmcF7vmpV1mfebx
tLGwN8g1OXvQY+iiqNdx9qdrJ+StG4q4iHsTwG7gRLeXglyExxOZKXXVtkK/fOfY
pIhyWc4OgMU0p0Z7s6QwINZhK4DTiwz02qMJfp5nOll9ByLqtuOxdQkoVcTH87cv
+DVCltwBer6FrA8AX2Z/9wFb8RswELzy7ozlXy/kYDQpKQchB1MQkYQc571iMCPc
ylcjffgjIzp27TMxKNU0N7BbuapKzLvSrfhyJaYFXY7drO4HwRoW6BhevumkQ4ja
U4xyvfs0PQh91GDV6KkorVLt/M/UWDmFQ2bZ55LtWHlnCKwGO8xQi60Ip/R6ElN1
0pZNkb2Tn9AN/5+E610KB18Y/xbMCkjxolCZyVP7XxLsy9a0JUyrHEftF93MfbRv
W9uIDbs9ezsnMVwwnjF6E/RWKnWD0i1NOMvorfIaD9CE4zkW5RCiSjcJRDrtt/87
wyGL16AEfZ7jfvtSi+aCMGCARnHUIS/Fhq53beV/ZBlFDdJe8ep8G0quEAOdcm3+
pPXw+Urs/FhqrnJLhA2LCahskS2nNsFHkbXVvZDQQJ2/d5rEg8y0L1CGDBo/MS7K
h3j0c0LisvEBQalNEGS+0cO7oRXWQUqAr3w/GlGNv5+CtNqiyTAmaOfn5lOm/hGe
AQlM+wtkCogU5/W2Ed3ItAADRZnm2d7cE0yMmn/YkV0SVvXdw3tPUOiiowdx5qYy
15AiNWHFmVWfFHA5f2IfPVqz6NDFjtLLpHIAHxm+cbyFQxljm8eTTOyWYPacqrOZ
CMnisvoL27TRn4hO4YrUPdgDUa6XzA9/gZP8wC/E3uT1Y6StCZS0Qt1w+7miM/JQ
B8yrJgNS2UVNwk1BjkNj9NrPDOthpIWS7tfFxty1F5ZOKqAK8FTydifhyQ+BEDhK
fCLTpOxDpD+PWQlYT510QSvFSNhBYMFrlJO2O8GqDWMyaswpJD7W6UVuQWnM5Sag
IBKLAPMcl7VGTcw0j6MO14hFkLbtY/CDSXWlq2D23vxtDOpfFOObk/A6S3jSTkRm
1vBBKTa6ym4ADH2096FOLwVi2/WEgyfemJ1f7Qz4qi2A/T1Kytd+H+ZrNIX/uGxc
SDV9Ha1uYDkRa0Vuvt1sV5sas/5edjloQ9ezM0zx7JYnKnhfWJls6rtXJrC4cDYE
LRF+f+WHsXpggYgJ8e8EObUC78q6ydnUBYZJFBQA0ltBQ2xyrxw3SwqYO+0jWkqE
Ym1tbxy4ybaSjJQ88NUylDm7geXQ3wgQzn0zfTAOZI2NDdBIgfoKDrbR95QpygTo
y7fnpUkTNP7o9HAZG5q6139T81ayCDI5gsgH+jZUXaza5yN+hxO7Y0bNcfKe1nUg
EIljpDRIzFC84EYXtf7QK5VEzKutKh5kw3SBo+jvfhdzzqYmE4ubYXFfSlFJLr/D
3qxwVxkJLWye9/ewyW17ZMcf9qUcOK1gENc+CoBsYPcfFWSnBwvo159S8w/wlSyz
AxYxkLagNRRKnCGyk9e2hRXlcFE8alv8mi3jsIdpCbnT3BVMjrPjxflDdWQQvmeU
ZP7mLMnisCR4R6moKjDPTWdjKJxi1Sg+5CbZ9X1fgWJgHT2pXf1U2eAhhO8Yr5nV
Bf78LTD4nHsZaPngM46uqjw/uH6AtqRCtf9AgFUU4yFnJqCE0Fp05ME/kMrfEASf
z1znq8O2IV7F16l8+PGP9hnBevBGqi+IAhO7XIg0Z+6kNuoUEffbSKBMNCy/IsNC
GR9VvYAuX4/qOHoMk7xtwOkI12TvfI+LUav+vEn6rPgMe4Dg+umSncmu2OYXvcfM
fqtHs9Nps7IblW8Fs3xY0cjVut8nXkqRZTVcv2wrVo6Jho128pqy4HAZa6rp4zoh
Tz6gMRKdyqHhquKdnaO3Zy9IQhAKyB5iwicUTA4YrZj3IlZd99NHx08RNWsxJkkR
N64IZzRT14MZf+hPpvNATLSE/XexWvkwAkuUKBkKIZJdtiOzN0PZJzQ8JZaApN/x
19ZCdnYJIWf8XBFYmm7F21M1geKPweqpk/mpRo+wDs9prvk2oJmteezmUtD4riHK
O6V1VjW9LzW788kO21URvlrKP8X4zh2tuhQxwH7H1Jewp9U+YoflOoTF2Z5yfxOL
azC/8pxu7HzBvq2oOVNDaVUtPls/GXHgbSxjP2CNLCyBsAGsiJvYVCEeppxnpfVI
DOUt5DAmdlC1z2OfzWI94qqyt7USZRyZ0j8xzW/wMAqFQ6Sr75Gr2adjnJbXz/Sm
Kmhas+ZzOFZqdEQmCXaB6D4zRqBNQ+QfuJ8SH8oT0sd8ZAlyXoAhCJiduNu55Mm6
HRuD7dHvWczxQuCTDIITTSaBIilj9gxwm9THkGNf9nxRDQc4+bC4/SY6fUhYcGs8
ET8X8fvGFQ1ghaphEoh68weF9vBNlJn9FrphkEKJwwOtKp3OUouTDoF7TxMopoUJ
+Zc1xmYvnHSAD5RAHsK1bz18N8phwAENp/mLQJz1VZOmVc/mIRMuhe5YE1xzqsT1
TwAVExXpW6T5FjCKL7fwmiuUF93ag+Waln9doA266ulxCHJ34oAcnOvH5wWbVM8r
hVNwdmNDlJN/tX4Ge1IwtH01JJ/tHy2TKZ+z/CjF7GK6eJ7li+cHt2qisKSMgupc
/uEzhjokrDw57QcE6Kee/yDgL+GrBpm6Tn2orl2sr933TxnRcL61Lsxeo2ZgR0Mu
KCmde6EBoa2DM+ju0X9BzPDv1zKuR1xJKGPrKcN+C7V1+g0IitJPW0j3y9Z0oRwc
6G2KNi6edNHOzJV0afItCJdH8wAitneV5Uh6oFY3H/PTYyPIEB8VNeP87XCwiE0E
X8VT79SGEwkFPVgJZWf/MWrVaIW1qefjhO50jLQQMp4B7TJhY0ocTUevcD/roIwa
TUEMbqsCjQjXVl/ObrS40o2agHBBG0my9zPAXV811a52DfWo3oOg2CoYN5vmU+D7
MjBDHJeyru+yyZ40YF1ekDX4an/i515by4gQV6f6VPV12rqDtHSXQLuk9ozAQ1Ni
EDhWOjn0maBz8Lyn5c+C8RX8mn6gSLuH91vTkeE3UHeQ61ZAoSVIaocDtMwnkA3I
voCvDFm/ODA6JSmhk/w/89r1nZBqmMioPkspyMocpYTSwGIach4EquSVYocVQgA9
AVbp0XE+a+AjBYiMmhUV44N8+1vgkDE0x2tvAU3eSrSm/4vxms3Xtn0TAwqHP1cm
EAc+cuaTjDVtDR4nQZ6nj0kEnBZEtPFQcurSEr/3NoD1lzGC/QkGClFLEpiptqxj
9wZsBErZpYnDoRsFyzusHlBiGiH5O4tS3zrMyPqWqLpdMndveemaf/jy43rPY2SV
781EeWEsTL7ngH2PfiFc7hWP0bsA66S92gEisfISm8xTrG6lX2mdAUEk7SDkYLj/
IC9sBxo12QIQYGTHIdLNcjZeI4d0zFUU2eZ4K4eOkm/gyZRr7i5rW8yV9IzU8y1g
qy8q3+dLcx0rPolEUpyiBRSCfS3ligIh0ALEn7isECrEa0OwyqiHqnHfxkDdibWs
BvTkJcj3PsQQWCyKqIKmDexnenETmqStp72S3ZJmj/v6quhB7FqQosi8fYNuWzqY
DyIMaqrVWWq1WYiiZeCBputNhT7XsRxt5j+81GwLPWbAjPNpA30+IKvSP4GLd4sM
0M7G5QQr6Wu2A8DuR0LgdKhpNnam2aCT5nV1U+qun3/Joo4GFYzUVPaIPSot0A7E
zGS7FhdHhW1T2RzNnTXGj7dLYpUCc/KHZCnK+ZFYCc8=
`protect end_protected