`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4816 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/anaBVTumwtXp6e/AWaEdufCWLiMeUob4QLvojnfS3Iw
NZsf7fG16hVr7J8DirsiRMEoB+un/YEcTHtIzt0tSBK+4XUZ0DdBN2u4fseAAKs9
celQ0qKTFtalANbj35qDZesykHwqqnsmntmRlUzKkz2q5F9sNtERuDLZX3qD/udz
KJ3QzG4LQSOcLAniVnfLgnJAsQZ0O8Bn6YF4rRs3WNYsvCqBORTtvcNCJjiGWm0x
OJPzcAQwKsrwuVnH2D0ePcOP+80jRh+LAg2gJ/tRigIMb2ugAmaEHHu9fzTARO5d
+eeG+zW6RPo5V6GGw1fp9bF0fgxuhqwIrlr26Ph6Gr+Zj7DdJI1glgJ7xrB68H2Y
hPY+bLJ+jvC6VwQyj4+34WEcsewMiLqhMABvywYumqr+eYFvXLCYhSyXST3wD0Ra
2sit39Jru63vEVehUIGPOqOebx+Dxujn/MxVbJBdPu4C8jZbukiXkIPx5yAE3NbO
ZJ6/xoMmj2J67xl2JH2RLkWqDjV3AC25AHutH1vgBBKp0zpwd7WeeGjD6L++LZx/
2Pnoi+7Pj++Vn/c7ahjzRch17PtEq7iu6+tEyAeT+DFRUQnQnDyLPM76QHvbaYHD
ttPTw5Gywk0r8jzhTkV6697MpFjxW6DJ5uWKX1HiKCXQqHnSytODv1k+UkOu4jlw
leCqUIf6AXRHnSIrfHBm3cRqA5xGl6bQq3pIntDLmG8rKrV8/awmV59/238Z7Xmk
afzGHq+MH25s87/J4FLsj1Z3Usd5r5TW6ZLHxPhmuYtQG/awjvNfa5NFIPay+U/Z
zxKYJoyUoFVfWPGh9PQ7giueYREMGbYfPFxFI39QrJd8DGajzjaCLlLtC95lAjFO
Oo6PQgxnRUVTuZ5hGv0BsQvxVA5QvXD6YJSu0bBvwfmHcG6Bb7oKICZYBJs1ZZ4m
rlyIe9DCsLP1dBaH6AglHofRpb5bPmVuCKL/zaJr8/DNT7XGURPcWtDpRVucHUdy
JhVgCMzIukZpabfT87JSA3vQJPpuuROK8SXpJ98qZP8R7Vkt1nIc+p1/+Q1oo/zU
bZ3gwSW678DZJKrQ6iTmtS5qRWRQUzdhU2Asi02R3cT+m5IviCcUHHwW5EEPUiEP
4zjU9tVbpaxhSuQawK9S5/OoBLUmVHQHDKoIeMcR8Q/c/UCBq8hkC0BhPfPwaVi6
EeANTkQHZXESsf9lwrIZSedYrkNkQUEJw6t5BQXeS1hByeTKdpA7MiPIwyKwjgWs
75QOceZKY5vlndN2F1zYUezLEEBzZqVH3slghYF7CU9eoFbcZkinHq+LYv4BZGLh
rWZ491McKhnVpA1aex8gwt30+GUDfVBAugASn9VG23S9jW0a4Vdmm5nqrj+CjG1A
Pe4RcpBKGwiRLEamYZ58wUP3zFkNEujZ4/bBN+9kDKzTBpDyovovWBCwuV/fRBL1
aOaI7BnbqJJyto5PQ4uGNsbPw9jlH3LN5UdEB5D8seZ3de6wdmQKUR+bKBqKkSGO
5ihFt2SM/zLwm+nkOKCpvXDRnMEaHt1RBoszm34HRSZ5dXtCP0emzuiJGYEQ0lj8
urdERhcGxyAxtT2lNb10P/BTo7GizKI/9hrIugoyDF0+jbEaDcwc03AZAahW//we
MyfP0G7rQO+bn9CHWOyXh2TsoVR3vC+FB2OXryVZXK+xy0GbtD2iaXS6VQZyfX77
69c0EzZVyPNhba+XfU71PACQzWz4CMm+CnxG0SZ26NKqbguqaXn/4OhnSwNJwOQB
GWdQONiNBUvf5qEgxi8qfwxsYrNJ4aG5qrSp+i2iFiSn8M5V9hA08+FbnYdK6m/d
dEEArXk6fNwWkIZdCNmGXFxGGP9yceYeBXXPHGXyKk1xZQkfBw+N4PJc+5aeXblL
dXiEEpgfLbO3naaFSsbyjfNGYsYnXvHZS3G04nBkb6IqWBBXtuF6pWw2tbft2iFp
jW72FLmSq2bfSRvv9UrJtUalBLi0KsPl4tZe2C9JOLuHkFEz4L1T7bIolioxZHa1
LMjAy8hY9R8uL93cM3enuTtSpZh3Y0z3U6gQx8WLDoNOCxl2zEtXTHL+Q23voeh8
GFEELHOxrPkM+J5W/ywuQVseg5xYG6KVvzaAgu3i855DZVP3olYm+sbSLya5asqW
Sd4djUL5QOmWkW/qvBnwYsdX3L9Ygvj3ywp+sS9ACCnJziWJ56sO+5BEnJNgzESQ
AZgE6btIxM74kBt7R3HzrYrNTZFlzDP/QoB2ni2lTj6tzxpmvTx4+c1RYbl+0bju
5HXGMV04XfEX6Q5wgn1HpskGkMYNFg07Hv8MlI63R11TEdYaTFmNcCmskx0/1VxY
dC51Rzq0r2Mu/zmvolmLqtit76AZygrGw2/Fu3DHn/T4KtioHbky1ugymv2Sexaj
IODHLymsgwykjnL/L2bseVP+8Yi2lqcffjnJWlQZ/xPGaM5A1gapUDFUKA8393BX
qEhr7/SR5gA36sQrynaCyoYMTnIZibjfgeWHjh3DyhGGA2zgPluwTZhuCumE5tMt
MXr3l8tXQkVLN/bh7pri24KuOLE4oT48j7FqL1hPLinKt5vq15cvZH4236E7qM+b
pLox9ERFQelPdWVU8unJK4T/SPElSPgksE76DHV7z3Easln0rdnKXR9XgSWmY9hX
2zw6yamnqswg26KtIBcGP0Y4LVePJWGrGiQ6klf0Xaq82RtLmBy6ecxOM64mNxH8
d4FR6JPc8OlKfexBSCs8zMAMptwl9AZXIMVQtfMax2BN8uU+gUCEsrXKX/S5YNBg
LoGAG2f/cxI+SggKwUI+Yvt2e1tQ2WaXJfRaTJuBv2T4rI5hMB29oWLS7gq1jrmZ
tyf1J0uQgIwfc/DRY8ALbNsDUU5bmIZh0UyI4qwi2lyRe93KcGX0BrJTR24IHhwE
pKcSOSyt2hP5PZ7D65FWm7SPWD+V5lsBxcWx73LbUDiGOfu+bVk9MY0/sgCmK0ih
bhkJLOO0SUEqufDxhFFEMPIoXdOS0hDNqKbOqguaR9LgcN2QydvFqvQQXl3mZ6eI
MdVpR9Z7irGnHy8qKksJkx8DpcYN9g0jez87HT5LobOojX6+SCn1616xVWxQLl1m
iamfhlTyw8wxyZrbvegIobNdSAfT7KYT53F9NUc8BtATltYcbwS0MDQCotTreKlO
6QaCVReA5qLNW2vEKPBaWYg/nk2G/oHnRsN0ZuU9Wi2yMwh2GfooSkscPfLQqdFC
frkv6kRpN9kFovthyqp/Fce+mnsuOtkuhOvZhuPI8KmHkNipCVuU1W3YEVQHNAX0
OxXmEhctLL5TIaQNCiPdTNUrU9kvsCmhuFLdYbSHt3afOODPir2+yhYeLX8F3B1I
PqK3C3bxBfz2TqYWrCXxdpDaXLoGoF5VE4TlqYSb5z1xnnvVIS6JvPvdtxZ8pH0a
Iy8wiAIUg2giaKnZTyPQHmKvAJJAlFYBP1uI9piH3SeJBv08wHjZPgfyildpGtzR
HHYvolV2BCwKb2IAKwxpIfpBUJQ7W3RZGbUy1ye9cq1D6XIYr49cHIRcB+UJM2v7
xKDdvfNEpZmYknqRxsFoi5AZ4SoN8tTgedVvLK5cT47wMQiHiZIz2pxFf2bP+j/w
QOsM2zqZYMRJoWhCUIOWAeM+IBluAByGrtE/BDQa3lncsDVcpA1BWzk+2k4Cwb4D
bWaIK742LZdcQmhf518NGWn/08MpzsEm2+4gy8nw3Iu5wrFjC3W6IHHI1OURxRCF
guqzrrtDmDZQG5bLkXINU77PLOVn/yXf6CooqcLNmNyAPpwwsOUiViMkVPpFoYg7
q0DpwnIMdHceayUHMZa4bwb1sOJiVyWNe+P70J82L2st4FJBq+PztHVLIXB6/rC6
F7HgHRxbIC8GzG27d30WW20W0dymw52kTZCPMbGjFlaXKcy7YFNxidVuGmL1yfXL
r3+LZ6K0hLlt1+LycX/Yq2rjTsvQ7O4yyl1UUhU5zYGfDsjrF3K3NKZCawucZquu
A+VFnUu9zpG7YnNT4C8oPHQTNl3k76soDvawM92uaH3bhLpPGyrGfOTum5G/AicI
2yioX+O1dzMjuABguV1ibXMjFLSrJXD5CNuEzhCf7yfB6X7H5Q7J2bnQkTUUuHiW
JLy238QXXc+MkTE3D04SotYoXLzjAX2crdJGWfYek+rQdQFUNARn3GhJ+g/dqSos
bKhEoQjXJRx8RaQwM5oTdjV0n96ZRc3NJ8tS9veI89axQXWOOxL1HYoQNSN+MO9f
RkW8OHynsQGLnlNJszHtPdO6Ru91ubxKt7BLEHMEOYc98lYvRRTxNcf77i3VTJUo
Nc0rgs54t88F4opdXJIsph5odosiax80x5V4SIqPITTEuRBj87DSETqy2zjwSwK9
iEtL3o8IvEbpQyvfCKJO9QJUWQqWS4LkaUOIVljHEtR5/avDoRV7B4TuOmoFuJeo
r3VgwhPQ8rcEMTAw/j9TIlPOSYLxwAyoABXBl33KjbVIxFcSEPo3ErsRWr+eD3S+
f+P8aJd0FUlU0Xx5mSlFM3QY9l74gyb6iSo4FavZzvJVwzGiw8bPANWCRm8nOmNS
vVniWknNeeQQsX3tGD526AxRcEZHjZOE3wSWxg/zO8go8eNHeKllO68waEFv1mEH
cbyMgKrLVEseg/5LdUP8t0RpVRnVAO3qQmuDIrei4lUbF1Tx9sHUKTInD28f+l1J
skXziU3/sqYbMICwrBtRfNW6aVugX2xA51ZzeKYs7Ng+03u02dBiF0fvPZ10wbnw
uUefgxMQqBecNHIchXFjfUdOfUhh+q6Fj8aP/zcbV9EMEYZOwsFwy39KM5UdSJdA
W0o2FO+3tirw342ndlPTIPs2aI53m3gMEH6osSq6mNkJ3p2gBNmexvFlXVMTLnKQ
CV2jVWlIyDFXGbnOx/rROTELiR24GRp/KZQz/BokWBBKS+E+fb09fOwSB3SH9Oce
wyyWFHILhvVMKiVatMq6hUPOZ3g74BB0AhnvOcESlmcwUCH9eiRBP29Hl4jwz5mQ
mC4WFaZoZWMG9Di/r32tNT4jWJkdL/UZPyGkO32Gu+1pLcoI177KnzI94hExurYR
TcnHT51cG1FCfUvGacMOZ5P/BAg0T//AxJ7uZNjDsw2tERExpma9bQCXqfyUgkZp
06/SkA89NVk+O/DcfOMd6wiJ1Vy5co6ShJEzIjjfpZvxfz7yXrlFaCcYOJbTpVk5
csntIvL/393BUD6cgAJjjtJXcSIt+PgmH8CrH8L4l9tY7rVYtIurKyLJGn8uQ55k
0Rn+m9q0lohS56Ce2PxKv2qCAoNm7SmIFHkJ89wFrF2QIvg0jzwzjJ4tPSWK2KnF
/5gzerd4REX9cP7UqTO71G456RThiXEUEzEAR8FJkmHckhSMZUpWB8VMoBxoRJzv
dx8C7FLcODjHU/iJ6KyIMbv6ledbfDepayxefkQJ0/VR0zU7SOqumQXO9vg4kiTq
VyvL+upZLJmT+WU8lORO4c++EUqw5QhIZ0KSeFpSfcaAE7JMNfChJ446XqRwHCXL
Odw12R0lEvmZ723/ghHMs1pU0H+Gthd0dGeZNKiCtAJKEQ9FuPaoUYiI71MmuiOa
mxFRYTmffsTCHCBTlOQ2CKWH/47quR4QwPa0MzmU4K9yHUNczJka3cC0rMPKcCA7
dgQWKZNokPG6HphmAMq7uSfGw3q+XN8c9rZ3easLfYH09oNRcSp0fw3/+E11KW7F
HY2yn3CW/GoKUmYngpKzIVUyR+tH+rd3sWGW6U4toiZQlK7/qf7YQ6cO3G9eVkPv
weZWWaQn7u7htwOOZ7D+KMGwOpBDYLwz9jDXXt4zLQ39CKZahiLh5BhilVHUYH6M
9y2QBeLfjO2cnCGPLFpHA1upCmTlCicmkwe1dkklFqlLTMkCsV6J7DCAyOIws2tS
dpIq1hab9K/2VJY7VUZYBC0XHYOa0GjJMEwznTFpAzbWrojzqD0433WbkHopXQYv
6qO8ve7X/PqhpRr9STs4O3u2DBxufmNVaSkt0bcOjle0Z4RhLpOJ0OOaWzjb4plm
uy3cwgRjPEvaE7llpg/+bQj7JBMGreSLscPl6EsKYyBvGRHknzZgIypXbee87DPN
BUhyMZWON95wsU7Yd7+J9tcy1pzELthjXEc+2ovRN+KBR+MZ6gGJrdWHMvSpGhda
CcAN5ZDkkG2QPhk5+kRKXraA+HglvNXDmzy29M7JSFHmtQD8iyQPKV5ckvOzOp8C
nrtc+SW74i96/E3ZTbM6Jg==
`protect end_protected