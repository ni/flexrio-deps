-- 
-- This file was automatically processed for release on GitHub
-- All comments were removed and this header was added
-- 
-- 
-- (c) 2025 Copyright National Instruments Corporation
-- 
-- SPDX-License-Identifier: MIT
-- 
-- 






























library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

package PkgLinkStorageRamConfig is

  
  
  constant kChunkyLinkSize : natural := 2048;

end package PkgLinkStorageRamConfig;