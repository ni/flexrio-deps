`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 33072 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
0ivLeOT4zMq5S+D+IkEISAGbXovjuQHwtL3OpGyyXYbkYNGwFO7M7kAbU6iEo9XN
/U02e92woUWLyhTwXcv1mLOQxt6waD7nuXRtJr69HjubsW4NCbfGvXWv6VPN7266
RZximzOMcRvgeNy6Lqket7j3ShPfhdENIi1U1KxASmBqbUNYKxuTV0V64S1C+Sgx
jMSRkyLBB0HXjsiLQvKM7p5g9ooVOR8gwLz2OLnz5xMAFprjuPb2YXWO+zbWyHmh
HythInBI56ofzgL5dOXhB8MiNyHbPlHI92vvVTskNzb6OiIgUmwiDeQ6ZU17I8lv
JVMNMg5zz1MwTG6LaLiMrMR5TmKBAcNQ5m/CvHlMCy18TxLIjPT3YVOdUVZbdMES
d13sngHDMSPLrQYSrZcu0pK9PBR+aKXx3eTzpPxDqvrdgDXaFERh8gEjUbVtGAH8
CQWk2nsZ3h0j8Lc4S96mSSTFwWoq9WHeaKdSsOIVrDzFlsuEY86d5tC6tBEBsyKS
8B3UwIFrY9rIzqWiGCmxF6+PNUAdEA9CqI7bxzwc5TqSC0p9COY4N1C0IIULDWKV
19VEau4nH5wn8Hkq3pzzxJy33xQaA59SYuJrTHvCTmFhMbzZ6RsdUf7Dvd3HhhqM
0BoHBNzHSyr4fJ/fW+L3eoOvLYxqs8U9jVz/wHiwFroEiuVY8LP8DpOAW1tEurY0
1CMo2QL7/yyvngBQuxu9uhoc4bVf4ipts2GNOtNuFYNNQX78iK3+PRAN5GGUd4If
MVrwpzgGHg6fLvWwA2shZAvxz/QbOLajNNldBOVytkxxtIY9COnazirZx9SSAeAC
1dUcekE8vpuEhVtZvzfjhNcNpkMaPfE5rYIRzjsyEkMZPl5J3E1fJQSY/5cVp9Uy
AhVKuOl4cHaUVUZ46UPMqyExzpaAFIOZixvj+ULjuS2gF0hvK9IBxapr5oJN9U4G
b1r318oZaSHztlamm+9loK5qqWggxDEXlK2QcjAuHyxQaZw94ZdYUsZCC06ONMZ/
YmBdqLpQ0xqb8LK0vDsfOC9VSlAbI4vQ+2FWjyJzIgMrXrv5gTVMt/PVBJsQnj/E
v+OQTC6wABvbhCJtGuu4ZBCTz2yXssYa7rP9iCg0rZKhGfnxwtrTqbKxo5LidG4H
gDuWj/d62/EYsnIGfpN2xwu1ba3E0tQMgI4v0cftaLInwUzrs4woxgJ7wxAvUhFv
Kvsnxx+w8RLzT3h+H+cxT4RbUdeU50uCwF9PskBAlIWW09egJq+V8kr5/GTjp7tz
nGk2OtOGe5EQrLfyfc6aU3AKZncmJklEEIo9qEAY5CNElfjN20TrnZFTLPfUA9pr
0ttQiROj4KtmR2XftEfmbK8iwMequp5BNB13+tIaR30MydhGLmkzNpJRf6jh/1zy
n1cKMM9hTPaixmlF6eOC8vvYQBvs2X/uwnfgcHyVo7YvtyjCJzkITfaGaKqcqGeB
alOZQR3Tad5aQ/O08b28Eu8RBqpo0cPWp4MHKRmmEbELWvuFqo9UZowS5+1/AHDW
JeRki8JOk1PLTQiMfaxs/WA7FI3Hjp4CD/9jt3TZtJQRcXjTgWRSEKQybKrtuWMf
2FrMTeu1ZfmnibOURpkQonLS5Cgoy3btf3pYMaOEzO1cV+hCmWdqOodB+RVeOxz1
3yLz116btfrQscKbIFObDzN41S8V09FHgy+CLTx/uz9WNu3AunpkUXudJpE+nNHd
Qg02wNOC77+Z+1Qoxe1vDTe2K1q2442jbdx5uJ9yuaaShldUP0kRz/udc6ewLI70
2m4z2BMsaBNiBGMCzaTBnNhdyKHbTkYvpiyEgtGRJZBiZZlawsBmfcX5v3i7Hm96
gP5XRk+GKlaS0u4pxC2gV0+yf3khnnJ0JP5vr+/CCxngOnYhOCs0UfsGyDZ9pH6g
8qc2k/VaNX38OA6cZNrRq25/YseVXr+nE0PlyVXaFsHwnZqEN7MwWKnWKRQodxKz
uVCDC/xphSu5PsB9mP46I4AQTpUxxXrWCoYU8GMdLRzl8sUMilXRE+YCyNoIylkU
IVFvg9xFV1bWQYE+3WAMWkDnzKsfAy82yq0i0iH+5esBMjRIY1LByN0ALyZ/Id3I
shkxpKbn57Vr+jTG/r2fI5RUuKebRC2mD5rM7GhelVHv9B5v7kgWyaA8XpBq7ZiY
0EWfzcTSH21w57TfrrRSkaayYi/nHaBXh8uHlCMk2GvtEYof1eEemv0DGtQKhpLI
cIAXv3JHIpZlXOByemvuDMm2hR+RafBv5h5JI8oG9m1vuGFf+IL845j4mrqOEt5+
Qu77ALjpYkTH+LzF0OKcI5Bq9ImwWTGTUqBk9bD/gvu9nl57S5+ib7YaY7iWfPhw
SIdExghozGK1s5EabHpbQI+RI7B+8xVPMuB2YSP3bAYmQELmjzHKKiA1ldhvTm8S
H3dzO33/feCXorTZ+VoY6WLYv0juP/0o5+nrc6Jp+u/ZPYm/whh98AULqdcReoex
hydXaqGmd3kFJQqhfICvT8yl/UBVP6a1+qrvPwzrGUA0IHk9KVhQDdj6wvN8wGUJ
uJJwWP+Dzk1d0tHcvkrfD+Y74bTeW8jC/0BQS72e3I8R553OLY0ltZE/h4CCbEOY
R6pVJip0bes/00MWnAS7xsGsqwhel9NBGXEEHXOJkkQHGbnEIe1cLUIzE1HOt4I4
5oaPVr4DMYaFzmMqjBziTnyibu6SdL2vC9Y1MNEbef1DLVENwM0X32i/JFsI3Hnw
bnc5RhfxKxvBf8PxLdJPFcPgtoB2HS4FVW6s6MgF+4yDyueAaq5Q04tF5HDXYiE7
il6VnelcAPPWEKX7nvTLeW6xcSAqxDm7WrQ7R7PEsjxKT5MlS9Tz6H30Az1AA32G
H9bVSdyArhiNVG5R6V7Mga62KOplrhf6eg+JBJyhhMme8J+yY0z6OABNwzOoCbko
a+/RNC8PTuLA/xmxIM2PlBeK8GPMmNM9p7N8Oa6De8ootQg/BTj+iXkXmDJmKp49
+g+p53RfWFnRb52CWu1wMTna2dcOdYVF8hWBX0OWBoDBf/a7xNlREIVklgKOIdVh
QLMZiIA/9DBsw1QUR+AACLDxZR9lWpblqQ1AI/4o4xLwNUCYtlSvF8DrAgMj1tLi
bVJm+/VsPrAlrgM+5Shj4nRHwRYcKZokGWOJBWQo1b/wkPBEWqOHcT/R8ZQ/RzEo
iQZC9rCXsNPelYQs/ZlhIGvUNyi8tETWWqO5/o3lMMud5jMIBvO8k5OzpMOHEjFq
FHyFrU4WZLhvv2EDLTx0QOgBxsvMPNAKVdhTz6m3LpgZzreFUimqM6ecGdghuP0k
fkhS3jNmLN9Blrrznbht8mg/B6LffvMNycR2Evitw/JtCZKvke7CeNrg6DU4SMfn
f1Bd6e53ET9QICnmapJKqUxT1w0B4BpkzoIhrT5CjNPZ5WlSvj7Ep3Tyq7eVR0WW
HbetmymUJ2tuz4HNbRJZDzVoKsP2XacCQZVZ4xJO0sJfavCXmxi7+SLpsUIF2nDk
Oo1Z1ymOKq5wX5FFmNv7DwWbeIFl/2U/rhnEwfLCOcSXpY8IwQcuXRjNbWa/7Ljd
5GpkMga77W38fZUsBIo058ZsxKD28k3pwGXE+1XWb3MMzEGpUxQz0XNAl0OBmDYg
y0A53zFMDxW0gnij0POPo04cOWe0bic07K2GXANO/wrw0Z3uS4q/A36wr8tN9itg
2dqAsJpysMq8otwo8Z3Dh13gGCe8dffQ0ubTGXSSdt7PzCGCZFj05OGLQtNb3uIx
BMOmafOwYIAD6AuO+VFtle+EiTomGQeXgl/0Zk5q6031wlMfXISbJwP8h3HWCIZu
QWYF+oKoqAOd1xKinTSoWd/dzepp/a8xFuDyoRnfsjuW5hXUTnPJyDeQQJ38giOQ
xUV32SvBeB1fekVkq2VG4N41gButXxyrMYNo7HwcmiAny6xUVDalQf/NvjBB+yQb
7syLKNxzkmQi33umDED9M5FELGMcvCzH/HPxsF2PrbIzlhu6dtSvz6lh9XbhYruI
XZS6SFSqwc7jDXaezqtToEkZloi54nIVTTTUWworFNQa/UWRNwbXvLfuF0Bf4gea
f+lua/ffXQbpUx6gcRSEbc2Sfaijrt2QG0lEOxkxz97+Dy9tLMisL3buHDmaL2or
i5wbs6Kz52ndySo5IIhblbcM2tC6gR4GDW8d1CJi1lpBB/OWzzxe41rhl0MC2NSs
Fe9IXo0gSQJyNcEusaLoPZv2boKixP8hCMXVP/nSV0G1lh+0PHRnxyd3WCkoqg10
SZCEtqZwFKWc78JV/IM34AtnRSPjTFNN9o0ColHqzETzOTuZI42meUqUSLvCIESV
CZvW2LRgZt/YyLXZl6xRu80GA/zKbV5AshzKqwI97b8pjwXgDa5cSsafv24KSSqx
X/srPrafGydffWetI9nz04I5yAnaIIxGkj+cl2QC6tOhsaz/WiZG0VqSMgluEm9m
Md9nBoZF6YJAWMtutjApUTuSmA3SCtA61syxk+649SjGx/gB4bUJDIf7bLhRvp3t
lkRc2TPb4p2MkRzgYn5FjoYrtKARX8jjGZjza4hUwGW3+DjXx4ORzFzwrtImPPvg
eDhDd0b6D4zrcfjm6rfBudISAFxigNMukXW+wIGKd/QPRCewqYyDED7BZccE5SHf
31YUi6+2GeAi6aa3cBYBL2s5OXXTvOUXleKFr9W8abb4jLTzfAEW8UXZc2e1yY8q
2w3fvCiGBiuycFI+AgZ6qFqEOpXM5dHmSIE9erqwShRqFGAweFJawdVs/q5OcL2b
H/mrANqzSDsClsnD3akIcAGU+ZTnDXbHogEGd2AzG07bvFycFFUoaAIl3HWO4Pe1
oj0f8+ZYNA0c7p0T/8byHZEx6nvAoQHa6+UNXYwWEqG/Tmgdq12teikCFKc8cNmg
fyNLEzVoFsx8tMIHjy+D2qJWrxLafSyvKY9d9w2v9s3bxGGW0VzeR07kniM26wus
HPg04AOHNN+Nekm2j6O29CkM9lwmD4aiJGjgnrxQ1PalPXyKZ/M3iybP7hZbsFQc
PNDfk9P2bO9YsMPEcDOVrSw6Ox+gMQqlXuZ/FBG+UfV/7ytwR12xmJ2Ji9PittIZ
XT9aqB3js8+DR7kA5vtzDIMedqvKr7nKB8hWCblcrSkKTY6rcasY4znmHuw+8yFx
YwA/v/2ioW95XYXC/zEBF7AsPcU06XLfVj5s//xsrIqu7BOfWjRpJgkOWDNx3w9s
urZfAFlkn66A3xC9CHsN4+oyAiAZHL8iaSbHcpu2Nn5ByOPMxBod9iATEbRAKwYz
TM7clbmeAhZT9zXg7JLLRGv+gR6ZRFYQyPk/YAtOORLWhwy7PCMhnu03M1r+J9yI
MI0m3yWdcMHLx9PQn8/APCg6VIMCGoas/w29FPpG79JO51Qrf3jxqQ2ae43QKpM2
QHZwGe1vIjLQbaAHdqsahqwecv9oI5FIFN9WV3rrKEKi+qG766nvR/DzoCR8pAXq
vrZ0KdqqlZZuOtUl6FM03TekWvCp5d/nxkGBswPw3bWtfYd2jkAn57RRepA2/QUU
4pZN/m+wYo2KVHjWd1fP4QPFnvBnAegq7S6C0vc2JpjZi0IDI3MpksSCzbI7CrcN
21IlITQdbNOcot3BSJK/X6XIll4OkzVtiLGWReui2c2Xuq+JiDaT+vEKYOcDshCB
YeslWpk2hdDhCh1jbL6iRk87IGOW1Hy2mK8SjpLAa8N5r/HneaM5cfYxQBbDfw1G
sDRMls9mLuhYx8uYtDzmkFUpBLyq16Wcy1Y6el9nzRIs/SihH6e6tmQiT2gOcMWB
Kh+g+EdVcv/TmB3VoBdkAVVC/S4Tpk9wiNQlAl7KZ/EqUSp7vBuQum5iKpH29+kg
EWpiAvD4orvPA07L9Fyocug7zwZLh2gEcIshZo72e+QwEzaWGp7/AtJrqLAwKfej
eH1IRiG7knDp0qA4DA+q5w/G0xT0W3utQFRXtj1JR11sFr8+n34u/0QJd4Cgz9ry
htWU+0hHZyzMqGcnQEs789ELpJvjlfkTyyKB0wUpDSW+yniTTrq16m3PqUoQwdTY
3vUBoM6Od5ojoqaaa5bSr/I+XkHOcm8DSfpSP8VKpaau8Bsb4vu32+iBIP1KPJta
17fyWUyc6XXhUeJ3SIaKhzXfjplVrkyGOLjBigB6hfGw5tTELTjSqfCrBvRy5Io6
q/ifDNyJ+pJcrPgO1WTcT2EDStFyORB0t3XZsp5WlOSqQrdUdM3a5MChfIUYtOc9
3cx0pcG5CrwWTMRQW3MhrG+L0BxagA5F0BN/W/oAGgJi5ngVqI7mkMAc8AtYmR/f
WlMywaG/48oGFOxgawQLQqkzqEQGxe8mOnDAtiJIzKivmsvXaX3+bq+nM5hS+pmw
43Q9Wa+9dhbGO72WDg0Ga/zpnyWfsVQABqy55D7bywlZ6pry3cYUPpKKjXdW04NG
ZCR3HdeE337K5QfdnhPFs9hElKp5xLyTKp4WyirpvwSFFkjT4Lm1VWRweY3yUWhg
Inz5PtHAM/9XdgXI7a25OUrbM1WlJPKUbyftq6wSw3PQsgWuq7U1+7Ua2RsIZ/QI
xI6on10dASICdudQn6cQQoDfOLTdnKlSdqC9tjcuae1oEWDQFuKBsioTE3dZweRK
XMTMI4AIRAQfZWbBzddotuIxhzz25CmZrUDCLxogccJAl3CB9c9Rm5nUjKmxklBB
gSMUT89A/Mc/lPtqfauAaA15I78PLYliFtxOcwhxDeZwRsIwG7i16/mU4GzFjycM
SPEL1ejrNVZr3l2O0EX+wzdb0Vo22N3cq5feb2Kqu39KPl8v5+dmjmO4u3cQSnC1
D2wD6w3La0HvQnjwJkd8kYpcgy/Vv05kwTv8IOFp25U3QxSThGOfxttdLOJMaClF
gj99eUf0rgRU98MxBNwH3/xYAmDsIRUeX1b0FekhbZFB/xkuHUf2TPNNRAnn0K2N
THC5VAPTH39s6woPFNalL884vNvrQgZGX6d/ApL0TEuN/eCZvfx7mEHaFo59cqYC
+18B3PdoA3W1a4JTBWSnmOUfH57Js885NzQ5LCojvlnDc6QkNOrCSCicP9jR7NAx
JxBx7MdJEnTraukkxhsJtBpHZyQ43V6j9FTqYQPcsNaU5LQg2QET4Ytvh6AeJg1B
caiYH83XaxdqwMYmnDFuRNguajjj37Tg5EY21jOp3PzE625joTfegZtuy3eLYojs
gV/4AJZikTLKPeXQh8yrs+2usadzkGfMEDbu0XGEJ/2bdAMs5igbW67To0SCaQA3
TZ4x7X991KP9ExizHCzygRKyvXBG5otiqOAAPc2vOii0tKU1kpKlUreXIgMknB3L
Di7wzmwfC2BhWcH/AdEBpFKbT4f8DvFZNpzRbhScag0/NIXG0wsEwPeLSanQrBCM
h9NGVgvPyuY70vm00rbg5Ba/stEc8371FK2oPUgfdhnQuJt+dFIllcGn/G7EUVnf
vA7VZJ8ExtKp9n9zWUISg6Bq7EFPMLuERhi2G44+1vbwjXUEfMw02Ny2QeM5OS1/
nfOcDJD5Nr9Fhi4GsaHfYZfSZYHazXX0uHyvwxJWv1z01WwMz5dHoplk/5XaB3r3
bc5Am7zVRMhojGhu6woHQ84GFp2m+EFBytU6+YdZJp5N2OdaOzGkbIRVUDUrOPQt
FJJjrrtvKfqm4e3I0BzY/HvC6R1pC2hPaswxUDete+sNF796/LAR/yP8OL/n0BPo
PMp14OLY4WfxYscM0vUiCgzo9jkh3qHl97GbG5dvc3FJnTHM0PKBBHap5Uiu+EiM
5VdVPi4+IhxkFLLs3FKR6p4ZMIjBjnbooyDbS14GvJ7uupojxtSJxccxbT9tOica
MMwRQxIARF5CEBChK751yEjDGY3G86Oell4HIt/3OfS173BM7xnyRwQZa5AIs1aX
BFl9uy1eyYcdXKjBKKqDwE/huheMYoIVT/4qcWkWQol+qR8/Vx0KqtihZzsTJ/bw
D+/xD1qahU8QW8bh42mCgtfOH7nwsfzR36Z7WWVwRugAZOHES6pbTPkYqknlvV+S
jUrMUcjHqli6yJGpnjeEqxyoHA8R4gRCj4yqkF7He8N32ExLJX3o7PIOntD5H3ka
QhIF8oyO+4v+4XuUS9N3okzKyDU87D4BxBqnBries2EyM/hDDB4aqwTU9s56Kscj
jLFPzaiE2me5qPdV5njT4F+pse3vzyOpn34Ed3RNtAQ4n9GO5VU1Jd/a+mU9K3yy
mV7vvB4vHI84Lch8ShtdWU2/p55a7JwmlTl3MHMIbQ6cAuWK/MAj/LaZTl9cvneZ
7Olpjt4PhOzyl7lTg9vjILfiblgBYa2DSBQSU2NF6UoTEQWAqwrqTt4MXQJ+l2Gg
WCaeTB2TwUnHLY32CGppO3AHEe4txWzI3uKTBysvv3awCn8oTPWRPUihk15QyGsM
aBiT1oIeIN/o6yn5MJp33U/ZLzV+FnGQDhHjj8JXlGpqhSHnLi5z4y6PhQl5o59u
MqyH2in0vUIwJ5sExwLTAhF6CUIgFjdHh6gHy2ZkNU3qssTMuWqTErAKpspc+a4R
Xthy1BucXWToCUlp0Rt3SdwIuAKJsVp02RBYMZOtSmcCk8HYvjEeqCY/09EA+8Id
bA7mQGzIoMMTYRfVVrcZu0u6Yi/+jzCCYSRH71iM3mqi6+qRgG1uA4WKtsQrsZcq
+NXqqjyyUWZ1Lh/6Nw9bDJoG/RN3OFmJqKygeZJmKlpmVLWtOCNfeNCJdODVNs1n
waN5droRy0/PFdScwAyVZ2iQuvQB6ttKwSAJQ3QXxcNUIDK8LwT0xCSpc1RYHHf+
JKWy9/2ZOGwypgQ5cJprJ9tR6pdcxomy5narj5IaI9gCzlEM0w33Tmg6ds7l1mus
i50ayRNXWCJkRuyn1VO46bwdIIEm/wzBMx1sd3ztqdNoaOezDZNsef79YP+uGw74
iu4/KqDVx+8LHRTMHuOTKV1WJG4fbCphi5DxeyHOChT/GNiGPqPeLGlEkm7JBxoi
uMPOaAqkjSbkAw2VJPk+wc+4QG28QaIzDHzE8Bqa9wcovrSgcGDYmzbl6rM6bdXm
1z7KQZWhTUSXSyyzFsOGBJ0iJv5feeUeY00nSFwpweS/eSFAwLesxPrmzgjuHh4k
h2/NJIG2Qs6THlG7ceUtCwNwlepepVPZVtt9JhK8e5T6HmIa6Lyi2iS3gLVXO5Ne
3jKs+J1e/LCWRjmMEFQVEa1iFSL+y3NQ6Q+TFoBCAuSVGuEEWiDIS2sEceBCiETW
znH3gpdYKhwuiGCAALFImtIQqUigb2goWScvcDfvun1CrXVVk+Af8yZcf8rcunyz
wkrQ1AOrhxGYdj/D0jw7/LJ5adwrWga/8exzfKcjfSxB6g/GAG6Lhz+N/HlAzWqX
vF+EeTRUnGDyc46Rjpy2SC109r/GsPLzIthWoRiYvo2Sg7ROnaZJ0gE00g8K0lMZ
61ggKD/s+tn+z2nZN3+TKlEBpX6glDAj0CTnVisVNLTewmvoMTxiSjbPmBrh3e5W
m/UdCDSKlJoOy1cQ4xfnSqn91dbT9Mk2/zZGZG74O0Di+G626/7++Le46wJpVmwJ
wdV1+n8JLUkugwS/RE7Np2wdm9qg+yvcbeexgvqwP1NayYpf6jVgcsAyd2J0jcIj
qTY3Oa+DAfS99edjjsi1aYubyopi+DB/ta+OBHWeb4CHOtbzr++nyGn4QZH32U2a
CD5oS5UdEIDsMuG0ks8OWj/MdJoa1MqS+TaK7Rxk2cyAFCUzosv5AbrlyVVUy33M
adLsKDTsMn7l0Nc9vFzR3GJkATMd9FFsO3VCoSiRYDUt9+MVObM/JuUmXsn2UTZe
QVVAoCp687DsWrzIdBKo9IdEyTxXxxOvRU8f5nV5yxhevee6hDh/sUaW7aH8TyWW
TxRuSktz0nOFntUgB/es8313ZFrUg+gjHGLy5dGZ/Hmv4gB8gvU5ONRJ/72Qb7J6
UgupTny4h4GZFXeOvvVBn62lhM/WYgxC61zuGqn91xf7yfBOi5Ah72yoA2HaxvmG
iszc97JfnU+jRCl6S5odrjxCpvIzLUaP+Jzl+0yvhHYUHXaCRxnwmO1EePR8Taue
wVvM9iPXWyaPPH48dFXUb7VOlQbFDvLLExLGJqwolqOuNsY1P98BS7oHCeL0H7L0
DynXywWPhRy+K4I9EWadlIi05L6qKRq4ZfmQSFrPq7c0jnDTXvQl72fv5G51iTRN
krXY3+13PYKcD0sqcQI0V8emohAyMzDpifE6rCOQfDck41NmXlbt+2uqrvC0G1rO
CKdmbrTmnamr1Q5wwmiYl4OrmTNKkeqyI+inRdNTp6zq6YR66YokE+h/nI01fhmY
YqPvl0+0Yz0AsMSJcyq2Qa+euXPLS+sV0mrQK3nnuVHo0S5UlI9X3OejCPx9sRBu
098qVksbE/QbpVVIz7+QzHg+bSYhTxeUzZLpF38vUhkbjfUt/sl+pUDjY6xFClXl
/6NjObxYdbcdO2dxotcsTkRJ5UUncGpijr6Rw5pxMeNqMbMh7VNPCPVjKHnS601Q
zW2AwDiBPGyK6JvMZUrswip0AoVibHXXqG+7Yd8d3OqOXhko+5oFOFnwfrd4sQHl
LM1izG6IRp5BdH8emuq3Fs/6OuXK6YTSUiP4IF0HYV7cvCt7zsTvKOtaJ03LvgLZ
eRZeXXFSM8DbKnglLK8ITBLnOxlbqTSXvNwKJSlctTk87SgvkVIMFk9RVsTO9H5h
XAW95vdhS+d/WU4IlSZg7bhTPfVf8wvnDz3nheE++0XMJYf9pDT/6SjNiDW+2XXU
C7IDhY3VbrJ2uLVMC/UI1O9LWClO+cWRE3zZI5ApM34QLjK8w09+zcGcHJulp3iy
mc3LBNbh7m9nTuNWHlelsu51Av6Nr2WF6XVuhKbjcOdq68Q9lcaI0Hr1TIgXjNhh
tU/NxTAWYCSvXDxPwxuzi+f/G9/JDFpWNcyZ0S/cjWuhgOrnaZ2feTCPfP3Bd2Ot
47S6Dtj9rCpQpBOiNZUPEnfVeZZHtbuCV40KyRd8w0k8XwO/KdpGMvRQhRopdgEs
ydUQK6Q4eIvykHzArqmdxEC3RBUfiVRb7EFMQzWCqQ7esxQqCwD4k0O5CIl2NnG3
DlZXsnoG9zcmxZp5emY0xpqi8icWHs6ytMxOjn4XEeE4uAZjC347+khHnziHw71a
Ilq7g4/vMLFTICGn27FTv+8ImAszY5OGJ7YcESnJm2OxB7CphV5Z7TcaOzYz3Wcp
U0NUaGnjJq+sxJXCe9FEkAWA1v075Do2UsiEwOuVCfF9bq7e3pO7waKWjsnZxUzc
kRWIncTEy7fqi2whUn3zV0q6h7Tbjm6HdpQ51FAMSpj4gg+ghuvu99v0QyRaxNc9
mMEE8jDz22osM+Xm0e9QssCg0D5NUBiXMLxrFznvqqHTnSXLlMzLqa8avmQp4XCN
8qJrx3HSsxDdcVfuap76p0K6QJjBhSc9yljjKwN8P2jqA3z4Yw6TPOPte/OR+Q4f
C+7MHk1piHRcJ01Vho3Ocw0A8jku3oBW59qeQKQOx+8byMwpfGKzhR79haY6bBvo
7sKfvNVscf0jstK4LMmrDaMn830/RA1tAFC3+NZWo5axKhMSx26K1FrAnGRbzbt/
qUkeYBLsMhKj40OAlTKuL/K1jSApKZIcij5Vz7egrVGcY/zzBhvVExbdUs8PZlBd
uyNeLFkjLSrsYMeaPZXjepWOrSeSERWAk5ewgJzGOp4m9vtYRhrqxlp85d9IT/bH
v8rXwjc+Xv73hHoRomM3j9VxQ/zgBt31WbiaiIb+Z0u0wXjwhdfxrX7Wr7FW65Bf
1XN68eT5uCXDFPTGZYWwKwqMFcvMWYk9TOxiW2+GdVW6DpeCgcr3Lmu+VjLeUZUE
FBZSUTZsu8UQ9+mnNz9u6qIK4Vc7NVGPNqGz1H5HZV82FkmnP6sXy08c8uX+vV/i
9vhMtKzJkroqEfythF9W3UVuhqQo2Ot1BBEO7sX/Ptt3xWQfSq5kGbCHjbngjG0q
zoKLqcMd3KCRG6sLibJ4g84fN9hetooNfQwoQBTh92mNCgY5VmBxixb/q4veplD6
Rrl49N9x/BmFrPK9grY59FlSzM6H4W7TIYfPLzeAq8qScDrMTI3Rqm7hAMladYD6
R0Ct4wAXai1egQiSe0Py/v5DenOaTBRkZIKCrHbIoZevTs77KTL2bqDdG5mHQwz9
f2KIy2QrzACVSKT0mHwTqsF1fB4w9xlJg0P3aT5gG6w+ec+P670kK9ixarQcrMIe
aSprApj/b7qZSFBSH2IyFuPocaAlyUb30apk513UOoOfe8wka17Uj66WNa7QbjlF
uLYe74FGdXOyBCzzP0oqWiTHNVH/uxuEsK/GbDcqnZ7djQJ7hWvKg/LaMn/OXrpA
4QZFSpIP4u0hpShBvU9Y5HZ6qW5LrB0exIp3AQRq/0gwN3zTPYZqvqSNiCnbMxIr
3FdBqMQhOI2Sjnhlu5L1ewsqVTNsiQbuQAOnuigqZvLw+Seu6uwfjw39jAz4SIMk
ap4A467+C//ESwHKdIC8CXxZsTNqEr/GkT4p0oC/85usJ49DsjE9UzjXUtq+hESW
s7sumtJyxlpUmNirpCKC7px++UK3VwpXV/JIQxq6iiu+JCUJHGChqyn8MKrlxThi
u6SMSk6nwwgidrgCcYbIKFnZUo7+fqphFphbXVdbBvRmgJNL5QKbgBuoaAVXWSz0
25ZMnzO4NjcfGbkGZpNg397q7lR12YyuLaFhHMni8fGIneLL2oHmhMJgW4xrqgj1
HPIPVK/aP/enFYjbxfu+Pxvx67hKe38ggzVebyV0Yy9zS+x7o64wIwWZf4l2FUgS
xVGjRcp3tVJAVvYDX8v67uAhjd1RHdSc73rj0xOL1Rm/Hy9gxsDKhGNfmsts2eAn
idGItYHtFFKnIeMpmBZt+7H/mYeFDl0E2sK1s3thSBgFEG1AUSiXnP87tvp1oXHJ
o7Tu0ekDqh+4Nv6AidzRy49oBCFVGD/rBnxbL+Q3ug1eo49YfRtj8TSwmbSSJ5DZ
FHzAu9Qnm+2En/fGvYkLMUV31VX8VP1fbrHU1i4kFcqUNQyGlgCvM9Xq0r68EAvu
H1TFuP5tWGrWwk0dl6f5pAJQWiR1SFapY0z7jE4wAIRZyYsCZFzNSh7BLusLiS8N
YUD5SjuXhCCaTPIeDMC57d1BR4BSrMxZnCmHFDUm2GVH+5C7oRVqEzjterItqCGj
UEsrSIFFct6QofC/Tsl1gZ2gVqZ7+PO8LgHPCStMb+HEszS3gwGX+4BPuNRc+kuQ
iLIhe75fT0Crd7sqlkXpZ5ISKu0+d3KP65aRria9NRUT/MRC8UkgbmcfEtDWmD+S
ThEjC8aILdsqyCR/gV5BhyhpMgZ+Ddl2aWIP1mDYhB1M92sKCfRJX2sUEdeGfXOq
DSDxhvp11UhusISjP9lHG7nXiCkhP6GNDoGXDslWYLgLCJwxPUUnW3RqORynbc8p
bwc8gCmCac/MawoK8eXC7ijxHP60nR64dKIGHn9ZIS3lsV90SyETwwj9yvJV74pW
PAcsTySm0anUYRXGXSdKn+PRfXZRakx3kioWEejiYGcsSGge9ZnYtggB6t1LWZJv
M9LWbDhI85h5nyJGiQMSETi0eZw0Z2BcgaLmqAQswhuW7supdu+VHnUcZ1ubccGo
YIe1MPOCJCGaWnZLBgNa3ITMxojF8rXqoyOgZYZ1njtzVZPabaePyxLWGxZfasxF
2CBB5X5T8v2z8Z4Q9JBpDCLG6JjLGgtOd9iTvJj+f7JcfJ8U7Jb2g5lyu+AJc7H5
bsleIcfY1E+CijFv9SCbDFJ+KdVZBf0n6eqr1315xzYANHBCOSb1HQ1HlmT6/lDX
rUqbwgWD9XxUeiAuQqU0HkSI176ZcJteq1vycflmwJm3/Ob0f6q9PzZgm+Qdz9wm
XNo75o2KTXAuS3RqtShJNVWGTy+U4tNz8yds5V1bIHz+G6kUVZ9Fc/+7FGMnWxyi
iaOSYagHqw4EYegjfMGvrVtovO+zPFFFyOGZAh4P+NPf57MxMMiyrqtmqxFxvQ8J
puqwDdvbKNZ6+MHyDXuGF6LfgH6HPnCzaKCQSm9vTHRkZNN2UN/QaZFQiVOe3Z5U
Nc0jD1itBXfiNcfm8rhSHFziMKvxa9lO9OLlEDKsjOmziwORfxwx3AbYxn1P2+V9
NoQ3qn9MWcdXKIBXxOBu9issQoK2fQv56VGGDmC8TdY4BSpEeW8T9B6/xBB/nDSa
m4yOTTo9L/oLD+5yrHXbDjrkH9IC2Ed5cPndj5R329gBx5uWvkSZg6C5zBuWs7VX
3L+7gULLTsOXuWObUEZB1cja86G0ra1jga3OxBqpkUHdarqlF8RkRPhoMd+i2Yq/
kZLQxPv0Qe+ya26nOwxzFA9t8gQAXWiJH5owZykSTtxWQGGLU5rfBqJuVfHu/s9U
9+4cxPzB+DyqtaYTuvXpofwnlN3qgvsVu5c58HaTKqelmFHPxcZF6RGN5tvrg+ky
khh3fo3tSUVzs1jKesNcEvgr/40Y1zYPdqLxs3OrphDfK9XLUUjUVuaLvUcUBRRy
lousWJaML1ctGjm/6kpMIV6TtnpjajuFdXGl6d7CK4Fug8CNr1Pk8NlAM7qBnALN
wXBlLla+UWFn0CvbMqFw7Mb7f9q09t/NqZ16qHM2aaSfHe0407IsImGp1MJlYGnb
t6jqyo2kvBlwVRZyse6ZGPusFwDjTLxRc9/rSsdMYdAFBtTqaaaOgtz9xqZyAjCU
Ce/jhuU7xOWkJhEcTa6ZSgunKfDV8oU4nnzkDeZDiGmkdXwWXece4FbkitjJ7C1E
CTXXuErS0sl0ULR7GmsL0MfTwf3c2Y/bPCfweVoNuhQBiWTCQrDL/HmxSB/tzgq+
oVl50VUnPv5IS1YqTTbeC6bKhrBynSvelOT/w7hR9hfjWRSwT3KSPg0tAmX+XDt5
7kGnB0NWAIriyqIlrHxNciD2F6e7cpYGuK1Q5QywM7QGYi7PdUVk68eE/BRGbCVI
N8S8dOWBSnij25vmbWfISad9nN1jm5u74GZ5z69cX96PuP9q/pD5uW2C/yVNrf0J
jstoGTd8XYi01xookbU9EHjKlhHry58skLTrs466B8qykdXxwcr9BTmhzR/fzDiC
sxLBiJdK1JJfuWRQ/K/LlojTU7uJSKAbrQU5s7OGds7JKsoevpADyXRy+SR+Fwyv
BdDUCcSgGE3iKVzp1VGINIR112kDqmIb61UchQTnP0GWRdPoACFO3Low/hrKtNQR
R6mRwR1NYSUpfgQT2kA8WE3MxquE/YD85OeqjXLRjs8GtDOWpxbQuVDkNsCEMM/f
+BQCTNGUkHgkUKOeaStUCBlp3MLjmSw72OcH8FdqKk/lrr1bi7cn5/FF7RV9Wv1E
pLn6gQZO3IjZlMFVzTx8nMLnK8gQtNRC5bIWl8TUzu3NMaRvUA3KvHmVIaFT1zZe
URRRDqJSX9Juk5+a+x+F6RHvTwr0tDxybWO7r1x+9sXtXpAVwP2i5FNqIAQf9GXd
W7o6uaTSqc/L1jIME+ok7C+ziH2y9Iu/2dWsSaGR7Ikm6VXvtD123JHorDEHJrN2
BDsPJfaQkpCPPrc6/F7S0tb97jmuqjG9J04RQGHDyH/AcWoy7yL+z7ct9faT3pXU
qcH0rwTloqGPx/G19n19HJXFBJ1b59XXNna3pOAkuCj8M9x6qMTtGPYbh9poI3h0
Yfs+j8bTRspCGSUjolUICZvCWC9PvhtJsebwQm8dJY4ZUrcM9yoJgo90PrrkGLKB
5LN5fEE6+g7FW91gbtMTG4Dte0jMCGJWVJjq+FPlfnevnpAjwT6V8TXw0M6T+WAS
/x3JfG/D/PXG/nha5rLjOmvnu/Ms7v951yXacliJY1TlTQ0+YU1b9Jo3AKwfDU+8
a6B6HJQwXr4neKgxhvLzP5N3EVEH25rY3SuE+ihW3r+qiEbs6uCLqEWsAlVqeQ5E
/CqdPC2L5RPmryVcWdMSJrnSShkNMYlTUHm6fAgz/XEguGR8dtIKE30sN/l0scB6
Chbrgpj6kmZhw7P5if5t1Yv/fowDeNE8hnm5JmwQRIpomLKCFRjGN+rIlkxpM+qQ
afPyTtGOBpWQUjKbCUsYg/u+5mMRWSH8GbweVAPrgLnt0S8xXEaw1Q4tus/2Be8w
XgfxJUk6LsQORzqgYNCZ1xj5n/Bb1QFbTBAD/+zIDJbmUxRF+w6BE8/ZpKof+AMm
23Kq/bs8CWLCjLkEvT1KDgnJ7zpQN4LEmdNptI1m1HsxUHVsPd5BqSzF4iHX+jnp
DeSEZLqfOr9a1oE59wnJ1E+8YPxxQdFkZA+98VkNGkHsQLheYZs86CsJxX0VAqwb
kymRZ53Yyx2Gt+pET+hozS8yu+JelSjaMEo/hSH/pm/6ImRIWnJuEE0qrANaK/xB
GLpJzXB3QjzvJVhpKGL3KEhXy+Zyuuu4quPq/+MoeHJQPyMmXoj1/uM+qJoxl5SY
/Hzk+aYRGIzWo94bGJCKRH4qhyaAJv7AkG4bEr1KjtqpYrhsWluCjI/rdRfm1BUn
9EF9FJGA6PYHQLSwnXTA0En+r1p6+JfQiQCwlCsfOJca8hwIqoQZbxaVVUvKIyH8
m5piZ6ZpvRPN3PY4mz0S3fA7slsrVgu/R+bGYI+Lg4TKa4YdkZXjztG5oa/wg9V8
zUAjtnT3ao7n+Zci/VVSQJ3cZip3aivuVx4iZy88b5wQiyBXBNQOhSu930sQfKq3
e/blIQfoPHmW4LxW53ThY/Tfudk9mXjCcI6aUVGO4VAhsSSsHXqx1VuUfGKh+wOu
oDJjUE00PPxhDWmSPt71xtGL+VDd9RHqBHjz2GIyQjVm5TiPRho5i0v8L0knOVQU
ipV5FIXhe79X+xpQN8S0etaizKQNSOfX+/3re86zIGDNcdPm3DgiOkqJSaU664kK
mM7Fi9rUlZh+7Qi2e0p8f+xa22vy/aD9UH/12jYqeTXomirjjts5XXK7TDrf/R1c
DeoSKCXQbINs71WeC2Nsm2q+p/y8eX6X/qUqPgy7jBpmz8zMYhnC2kTR/FXjAyyy
sfro9YASw2Ayka5swK/Dc0+1ilD+/duo1rezA+Vr8yRnYA1tUCX/5rQsKb7mbXfx
MWv7wytKUvCoYlWF4SSPIcZzwTnLTHKVtZSP5XXurD5rmEhLAb+KuRfDLhNoEZPB
58wbtrq3cUbdrmkBVn8QrIGOKiQTzQtsI5rcVHnMdGfZKSx9873/9TU1wtgCJdUD
n01p/alXpqPAWRNNX3u5d5vazrnWQB+PiBAenCAiElttXN2bgkxPdmimwV7v9K8s
cQ896xwnJYWAK+inhlznHTaiQwjXVIWNQy6tJBBG50So0qHV2jl60FV3fYkBg/AH
GaSfPorUfmE//KyR2BFLQwSPEFoT6a9bPGWcPMiX46LnnsBJDDJsYsNWOmVkoOTU
zRi2vXIJ2CzP6cL5vRGgpASSwAlEeblPNVhB6VO2ZGk6ty1QKpmzPsEEcbVUQZ7b
zBL1I69SIswd10QhpWf3xnDH7/oMwYUB+dbfWy3LtcbhUJ/Myd73r1vDx3N9efbc
O5l0PhCzHZPXGcp7XwVRbX3ZxaqvZgyggYw+p0RxDtMBnj3wFvwGt01kdlGiXhiH
INUIfKlclDyJLe/G2EX3Og7hPIdcxtPyLmyKhjRJat2KYnxsCS02ENLd1m+Uaw13
cCVD3idIJaqLSZVwaS9SbKS/fs1wEyBIcaAqS6aFSu2qU/HxLwh8LDvyhv05j5BF
07Lvb9Kskaa4AAaU/FKDyoNVEQ3Kvks5CIXoEWS58sDlXI2tqyAgOD51ZF6yaCw7
pJangQt8MUU9PYjbIlbh/rD622d2usMGZKRg8b9wq24ErdrPGe0ijbistI4yFQu6
z4lxfn0RslA0tgfDHOQHK3e7BlxolKPVqUtLD8E1sCC4W4cbNuyGdwmLCm0ew4XN
OsVnB0HkRfYx80F4kJvFsYPAWsn7v5WS1hw8d7T8kdqm/Qp5c3LgcUWNZeaHiKGO
TeZms0ymBIffEz9ymscU7/LEESU4h5Y+ReNCguQxFMlIP771j8/xR+pVa8NmJJfD
2fDHslpyLKs+texymQxW4eCM4R122UDyOG08o3iIqwMSlt6GVkGb2kXLyId7B9rD
gjKftc88QCQVs9gNWZelVStqa80vurx00Bn6o5ldx3J+qAKG7OrMpsVvQknB8a1S
hEQvulfUUDgXQbp6NrpCzWGlDZiIAe1Ga/e8NTmCeIQ+82Kq6Gf9G5k8Z7z2Xcay
rTInd0BR8gnw1gWRBXAH9qxi5kUqQct6jY6tbFlNYS+OpjisjONfiAQWcjaaoREn
ia9iB774+xjhvM9K5l/ZMuFd9hMM3HeqQeKUeR8bXGsWbKeQt2PnsIFlZgR8Jo7l
0/Aan8LEuPlfhb7X1/T7H8q9Ec3VhVBQbbYudGHeRLlncL3b/4BLQd5vaCKpr4UR
VyEFT5Kl+Ci420mSLOCnICz43nAygl5LMSkcVLvWoBORbchUThLRYGRGkoD8BtIQ
LuhEn6RH7yv+Gh4Ru4di0pHEemjuaZyyNA0msV++YDAuulgK1pcHxvLicOkbE5Wk
0JnP9Sv4sxXHTJk5+k4gptNULyfK4Th4188XED+YYHj3zlG1L13nanYLH+M+vCWu
SJ+OoD3zUAUmGDnjagMzvwpRao2oIqzrWZloaP0NGWnctt0Od7m2lRVbQiHb4sLd
wdk0zVaKFborszFxpEiqiw6TG1jenTyHxLGpenc9uAg2WH7kX33U/L5UyRJsEx4z
+nOyYApm/i0JD8KPEHTR6D8li2etq4Fs/irOd2qL3Jjyk5o7Ws6Rw7M6vLlsZEIL
+I8SBg3hNlbom8jr65yR4Q9u44O3/jtNSMSTzR0yOjtqqjqCIX4khRaaThE/S62R
EWVr+qL4UXeTAgiBg3s5L+AY5qCjxnJiuZ8dmvefk8O8iDU8Oh0bwe7LyKo2xWSw
H0A3WjD+tY8nA6VaYTRl/fYKwOUsvSCDfYoQtmJVnM5vhojxvfa+50hBDjEiA6hX
vGD+oMjxBEePgBGv3qQvACbBN4vDeOgolLeH4M+a9sHCE7qGV1CcQLoOKL/fWMU5
wtMWbiez38SbHxjhuhj3tRhl7vue6T4xWXd1eidXhntqvRbWxxVQ7k9USALM+Vie
uw4bOVLWR3w4gb68tNFkLRoxUpgZqtb9Ihg5MXERj2O1OoMTkBnsVVgcTOsxF+8X
g1nSN6NxNK2Jp4n1FUqgdgPVzE5Yw7ZPbSMft2ATlBpj0r18LVI0PmUCW0hSN2Rp
LMP9mllqsgeTkirP9M9koBbl5jeCCnuDx4vSW2VSkdH+kK6k17kkxXAcpP3s9vTo
cjWSc0ft9m6r2lAfIRWwgi2qLQyvyvrDRp6TsMW+Eqg8HE6exaTQzym3BOQzpytt
E4m1/2+6qs/HrO+8uk5T6/2GJAhv3cqC+08gq9bv12FNss8IKuPR/DdqaGZLJld6
mqv3j1DBrPUU3Jen2mMBFvtLvBqmiQ7rjiDSg9u2j4xJgsDyuK0EfyOUorW6SY/R
91/VY4slzkrzGGlJRCctlpGBWahCszadNu/nfnGrJJAvtZyazwyf7ueL/Co4Htw8
gZb2c4RriTjtgkESX2VFTcc3b9OuWwDzNkhJ/CZpsc+r+BlFSdkvKi54dTXFnoIa
KGfg+SCD75yPMFzaa7rg1UCifqvKSIEwhHh40VGKTQsb2xHgEsEwiEb9os33i1OG
TV8qahX/JF/hqkyAzi+PwP0gNJnJ2rX37mxl+BapapBNllmVfFmHbMEMJzaYCIYj
BXOPUdeinV6WvzR8FmivDvGSn/Lb0hEabM3hJ1pPjY6ZrlBiNwEf8tESu+z8YR39
gaq3nvztIrGmaOGdycxMXKI8LHYFgYoQPvhTpjnsyoXDAQBslxfBH/HyDCQMqce+
KC/EhOsBh+vmchmyU6iWNOJb6rsoz44Uxk5u7cFXKP8TBV1jBMX/3e6kEGM8Yq0A
HdkAPiDeWNJAVw74zmAd5al+I+UGQskmNObcgVwUS4Ogz7n9LQz4aVLtPqZTZUht
yKt8cpBUyUj07ph3a3+taW2jGQBSGLax1FRu35G2rS8EuF+Mtu1pWmyt3VVjg2Nm
7nmt65pWZfs92bGw9LVfUsPOgTuf+CpjQkAAT+Rhe8oneklR8racPuh8txpmzzeB
kUmyo+HXeKEDqVcG/lnsfaqHy64PTa0gQb13j/kE4U0o1tJT5g6tlGftGkqj+IGC
Z5HjdNnmsWEVSP99gKmbdawJNm6dkQlWq6rkvzljEyYV+s4XEFSZcpvFJntXwnQx
PrwusnplIfujU2TxbRA7q6vgMGp9NCoOEMUyi0GaQ2NAm4CXkX9HTXIsiiryH+6d
z9GbL54jm/mTIj34pYGA9rPkNUqnxz9IHwpAnMrizipglnm72/FkFQ7v0yqRtrZy
tza83GD+7CzzsWn8cn3+rrfd4A7PvpzqyJkoU153x4bG0SjcUqnXrCnu4/G0JDrd
yzcVp2qZlmXajYBGQri4wR2uPRqxX361xBvkwjf3D/kK85f+wfRBaViYv32rePFp
Y5d2CuHv5cNqvtSN2F7uA6eqdZxAuQolUPpBhn2ZM8KgxEs4jBNsr7/UbCqHzyh3
SFs8N5PWcUTEStPE9dJULyXJ42+QkPJe4mw6F2JEuU4l/k5MicLWbbRMHhnds96G
P8KEUZwDDpXXl+jsNFiz+TqXOaCfaIogfQVq0PEwtK9oTOT7wiaEtdWRvs/EOi4E
M87Njl16wIoKjAJpArTKZyFxxI2C/EmCf7B0XUHhyxYGJctac6TqDGGF27QnAtOv
ZNxQbdBqf5hXowMkc0l3ozGk5ZTwEfKUkvGn9+VJ8WdyDJLzI659ZgrHTnEMUTAh
V/P80OeMSnmIIAvq93TI/IQs5QJGL+dsbG0zRm+07vG+PpY+/fvIrAQaOGgMrcnp
SywQHjre+7kBdNJwriyshfnWqDVPY8aVyXf/dRq+3PrpnvwiJDd3isMrnO1k6/sZ
ufosgvqJYntK2h5tYO1G3efPZHy6p6ifE7aFnXcK7MEid+XOje9eTx8uEsq79cG7
HQpZFx93e2TNjBzODUPggtHyTRWAzaEAHdjKRqvlheDkPGWv7w0yq/d/eEt/uRP6
fKvUKu+H56W2Z9gcd12Kfj8XQbvecOtuf+8yFvRZDRKygjJKsUBFA2GCKojPXl2z
46lf8IJ0T6fEJ8+JULcDXgRN524M8+M0SNy9nSW8LiyfVmH1TDNB9VaN4N2lGQbc
OweseI+V1nQHUUnnw79ceR/E7XihEGGLZtVm9sA742UbOVrc+okdBWRHUA4707MQ
Km6MwUdC+EX9yawxm/wMKDO2DC9Xn2zd/nkgIRWxfoiBdwPiQOe0tM6PdKeqThnA
fYSkjq6BD1+U3oDQ2SsZ8LHlVOclQvh4FTPE3pauyqvST4H2XenlbgfgKBxCWp5G
ZMk3NG6PbCBAHPyjyUW7Nwa4HD8hzM0XSrlOvmHB4nyTwASqGwMFDUBOHDe4YqkS
Trr20Db/j//FYn3b0OF0Dr4ETkpbyLG4cZQ8Tom4BBe0YZkPNyM+M8lCpwSG8PLq
sDMKwZE6vR05/1wnHNxGsdmoeHOUXbLxedvmhv/EOqY02hK+IPhyI4NPxyFdKIEk
iTjMET3s/PFXKe3jFpXNO8ZMuhPQBsbrx48/I+2tucJrJZx/4yVkAk0Du6Mh24kU
nkGHpnQoaSWYLgcNMAqyUJvrtUi0cOBP6Mx3mMBkAEyIvBwtZVmp1eTBJc2Jp+aX
w3ozgQIaX/vMf8AH9NWhnX3eD+27wazBy7HL6TiTNhoV83H/Qt+scMV+AHzLHkXg
VSLlh3wzKPJgnBc4dwb7HQVbLZ+noQF0wnitvsGOiGzBQtX97EgF2QTJMxzcRR+E
+hohPdD4APo8KcTZ2oGLlMWeEdNQPtEbEUsM8tA587LqwjrJmltayrfXcLMRaenW
VZ3dkH4Nju5LNxZ7OPmiWle/2U9Ehgx20/1slEjZ3llg9DlHK5ShZCw0NRWMhfl+
H7Yr1WOs+o38K5llDVTgg37GxOcNB9OLvigiUawtnR3OfAu6k1Nvdu5+mMLg6Rbs
v/TLz6LM/by4Kn+RGKRPnp/9WbALXxLGpNpiMKzdIFD08miLlHp7LzYoLMOtQ/QH
udtY+RbPRI6Yc+8ohJuIK3g7GFfAXIcBpbWi/O9tWt1iDj1wG/Hpwc3+9cCMajTI
sIwEuINWKb3gy8yHi8lWAnwfWOE6WHGJ/lfNtcFmh7rnnbZLDAoYUE+vOqm1bhki
veX4UiQvskbebrTZrrq3s2P8DIF83TkqsDTtniwrJh9uJdH+/9ti6bPorFb4IM1w
2NeNxCwdEmuaRYrZFznmHaQvb7L9ZcfYzi/t0kIxJ/eofOwUsG9g+MxPTwpdWLzL
XPfno8CGG6kcxivzJ0SePT6hnXDNixlR9OOC+MI1f5XTNPfOy92xc9/Rs6JiDy18
RQX+9oIc8ze1lr0NI30Uje55Mv8cdgl2JKJopHCQCQzPWs1octIMeHtFp2bgQLDA
nSUMNUcyuNfcn7gcSet163StPNQmY7z6hJCuAvm7jhOAtUs7H7F76AAHh9jj4Gw5
sN5O96ibAFr2IJtnSocVg5aWAHISiR0G5d4bV3eggAN8XebVyBGNAHfmk50Dqv8y
jmTeXEly6B0eFHsd6DiyuqrTuen/0Idb7GIgbrIYxrjZIhyyjNjw2UVgufdNqNKa
O+zQG9YwiQrpEXoSEXkF88YuOOsh/OmFXKWBLblriVlEyjzVk76Q4WY4226kaAOB
Vi3QlPwhkYv0Lv18lio2wf8OcqZL75O/1F2y2bbhVN3Zpl54h5hfU/cbqEqU58/C
298NFlFrN8dosnXRso0oMxu6/KOL3mb5MXSP00fBmLTQuKSiYfmZc6Qgp9GTszNi
IqqJYWd073pSM6NzMmvGJfysLE7c59ZFzSkpNnLvTzCbXXdl9a+42xTF8Hfo1lI2
KrYdmDA0GVfh846HAOT78r4lF8qgn2daSaBR0VFxvWA5VtjT0NWcQSFmoekmwDdQ
vymXYHs34Z/fQTSAFRRQBruNvbHgWsr/bajEu6aK9GjF4dECgnePva48mo0Fl5xA
XJQi1zWRgVG9iNOeC/j+lfRUO7VMDQIeP1RMAH2RChcSfK6fs32sUoGwjJGlGNYr
idwqY4wgDjBSdhKWpH0oQ1DTwNyPjaAeuoeL2G36Pl795CMCMZNjOEWHwUhTk6pC
RSRquh+3quL6OJkRH+7N0lNudWcWRjqLVhdjIBBH3i0ataySL6RUC36GJg/UJOt8
Oz4k0+TDcWTGLNkGlfxsYiLj1vUpRNGJ7kfzNoenYRY4FdRoHBovSJUWBDVHTs3E
m5wROSZZUrtha1M8AZjW1CnkxAfeVy4/uAlw96t5h+IzXLo0yFyKQuQidT15DA2H
CiK1z046wM00b7EahrOvBEgrK+PLg6Hk1HW800PCgkL/wPIK4AWquFZsgA4l1k/l
4wyJgundMNU8e72+dQsor0FR4AbW55b/meIuMr+5O0y8mwuUTyBz2OGwohz9WmPl
89ejQm37z0IYHdaoTiaOb82Mf23KeO5DYcDiyb7qF/lMdRzoC8QTF65DGX79hM1C
/niPT4O2U8eESVeXI3w1FokLGpRR4CvHjGiAUbIxAPbuYAnVCztjNglydyNZhHlL
fJOPSFviQegBU2ZdUNwSNr5GeF5NjvqVBB0CEV7YGCB7QIwJ+KUkkTg1R8DDS0Rh
g+0fLBjQblgmhqgSYXlpZ1Ni+7yBmFBH/b6RBo/km9hIYlTUURkbt92E3KNjBUU7
JamDTShNT4XB0hYDb6inP+wqf7xbAwLZeo6d5fWeHs6N/wkPwr1Yi3a543sEthyW
e235yIvD8ZKVaI2ZJyXr+tA6oCuJeWd532tEmttoQgLxoROFgOmgbPY/2MdXZ1Fg
TM0wNf7qRQAfDGWIXQ37oWpMss43yUXCo+yHrUmHb2X5+RxCWnrL5y84n7MPpbTC
K+rRcrwtQb4U3RLzrjfX0UQ+SZj71kXjlyIs/crOYSbe5Saay+7BgtEzNBv+ofQG
PBKd79ogki3Tyz+K5QhH9xH27yGtgaPaq6fTXfLS5lDRH6uLH0eJ5DOyADUHn4ra
C94vBV08FiTeZRszgmYMLtGv82lYYR8bUUXCJpOSghBHQw3uBA6by01WUFqOdak7
j3Zh0V/bkxZ1LDnsbf1RgUPUg3P+AjQkTFWLjeOZ/KhBqq5D0lz4BxAvn/6/u5wz
t/UwUxEQ3RMFyM35F8APa5kkGsmYgOE54F1Yzo99XvDIsBV49OxcFmG7CiqHcijq
ycc0NqDBEsBlLEbk0Mv2FhIZ5g5IJz/SspPIUH601Em+iLcfJBi5nRSFAa8MIto4
kkfrxxcPxNaCZoQJFiA62eSbDvgeFwM81MmC8TBA1tUEl7nD0gU7hIqI9RLguHPf
vNtNYSmacMEi0RDYpDE0ke9jtZkYA+n3e62mIWPFORDQ7rRuNYvnPaI2nVbHhY84
gPj70YhfhuBa3hk0sQiYLncvwmcyV16m1o2CveuKeQPyU2suEN/dQ4KQQH1R0u1J
NhZYqVnkvFZnXke5W3osyRWqAOqvvuAdgaWsz8iQX/xUavVW3lawZ8aWB/hWnenC
6YGo3YVZsAKHAdnWrc+wpNe5wTDsquuAWD/Ms06X0fQMYAQwm+LvagTpoe8YFtVx
DW+PjyA3pcjJwwRJ0/YLm9J+QgCDeI47nwBmS8n4dHD/J8o32+xvEAU2usBa/vR8
1D6M9ITY6SSPkHQwu9A7rI+FvMs8fzL6ywX/brNG2EueFM8HG6Kr+p8Q1v0voTGl
qe0B2bPsQDtyJKzZKOgvqs+E4I0OTm76Goy1FySSNc6FLkPYxURFmYWXY6rzhUaL
qE+acCB9EUCnbLyJZF0Ci7bn24OPMOUU1xsa17iLMT0kIYcbiQ2SSkBO/r6nc3iu
W4i3ktXPBR+cWRmTLsJZPnbJh57ncd9IV4v3c7q6nI+WmRq3mQb/shUkNT+67Ir3
GQ00OzZfu4mfJ4KcHgkNRC6zgPTcEAx+YZWQfb2S3n0+iVLKlLzhe83Ux1/8LeVU
dAI9IV33aBv7dozvy/uY/O0ueqvQAf8FzNBsMuK0rrClFpI8isBIacR0h9ngBPsO
t3Xwq5TSnLXYe8UP7dLHxVZS3fEMkg2z8pBo8NUt5WkEIKVe9ImHVqyejNB1yk1e
4koJ+pRAv7bJfR/FA8EF3fOuTtrWtFWwjzg0VkAC53G/KRmaFv5smHw0jreA073W
gfSV3ZCuU2ZlvP8aljfdx3ngemzCDmp3DNvsnxHZIaaVM9/Nw4u9WWppkbSCExp/
zXa/Kx/JjVgeIjmjG9h9OqSnMKM2KdAChx7Z8KH5V8Sq/WxhtUc5bJRkmCkxO6w7
dT7mGrgWZveLJXj7rrX5z2hESU/z6Bf+Lgta9uj9IMoSybzlvGC0KJxaRIxUYoeE
m6RZl1TK/pI02mub89/CbLjoXV5wHYgfYuVoEq+qFD0EDpuxjOnaIIPJa5ZsBAmh
zm3bOAX/ePbKAXvv0wMvCLWSLsqa20xk3CrNxkzuzyYi/fGNePT/ZG0xzh9eICg0
qqbpAFqT6L/zwpQ2UNAyJ8KkYhQIVkoyJ2+iQgReC0a8WCM890bJH+RQBYOt2XeQ
UsyO/2tSOYu782TtEpOw+hWVVSIY7yU4JZBEsbB13MXt5E0jqF8gJutIBXmwK6OE
4FetRsece38GxhiJMODy3FVRqMr1Jafwzu0wibV4poj6jn0qxc6WRXO3Zc4fmiCy
FuQN0vTqmcOfOsxkRzCawLnuO3KJh/bSamTpYExk2GVnL3f++NHVXqCQ029z1pjs
VcWQkc0fRc88KMLU42FcZgWiL59H7De6gydq76xplDoYrZXLQXmCpMlxqDT313EZ
ULs3pRJ9rm16j1xH/55bw/+1bNaSxYBnEaaGqSOyMICYD/6hVUCs6exyNPxIVNa/
7X3HoJcLdAP5rKl/hMpMdjFTL8nUM4Lxr2f0Sw3tjrIf+5xwPx7pA+3j5gxbSG1z
diHeL2l//2vPPpNPAOZFCLwU6uuE5YyS1ky3gJ5v39yJNIaCnHe9rzkr9Ncqcntm
bnEQjD1QVee3v52TlukFkaQoWvKqmTQ8HXP5nEgXL9YezCGvsq0f8y9Ynsiu39bU
4e6IfjryP++RZ+kw8kJH5WLnsYDGh4kdek77EdQQLLp9zB9xsJt6zb/Lvf7fOsOT
B4uYeMdu7cfcuAF77Z+3U4yOBhoSjk8OhXAPi+1CsYQYVGTVnoVeE73pf026lLq3
lB0vtF+ESx+SEpEYAD75zhlXn4zdDUVyRiGumYj3Y13Lg9er9gu8XG0z1s2/HmGm
g2pMGqWoxkhTzzZhP7yQeleNWEJ2O8VDMw94L23xs95zdWoetpgJRGD8Jw2ng2rz
45xiOlIxANgmeV7JzPxD63OFO1dMOFUn2HeDLDRCzI/N1Gisf5W/+8g53o/ZS56b
P4swYAl5hKMe7RHBmOOC4xSEQuNqWoMxrYOeB27CGcNba9uma3earUQ8HKwFXvcc
c8H2jj5m8rxRKmK5aoQYZUM0qDjjU+KBR8fNDCXBBFmUP7uRwIHlwmex25XXpmfu
PuMuQqRWjLxOEuUchtrLBMI6s4tyefMfCuqnsAOepOtr1Ftbz2z5YwtxPC/4GxzX
XDAK6r8FCS7+OoHHezDxYuiZh1avMzUJjyWhCcxaJ+NK9KCynj0GzkMGx6SdkeeE
h88MJlLNY0WFxN56I/u+464tzb+agENBYJwdFIMt4/QOTAwednDN64OUcIApQ2/c
sYi4N80sK0cx0SUnSYSDsVjqW9KmQLL18iVZkpXkzn3vjLIj9CWcDtrbJcdWa0OZ
YcXL0B25ZpibXdnUG7mQg4XmNwYBN/SMK92xPqNMbX5h6+nE+/IYcq01pinEOu4Q
b3vTLiY3udAUP/uLRCum6aHP7MUTDOvdlcW3n+XnUYU6YBsKWjFMkI/Pd7oo+tqz
6Vx+KgfJDipAiG2pa+qak8ugJrY8OLnsb4mJZdRZMoXkJjbpxZ8S92D/X2lYR2rN
nMVBiVZcVfhEKY/sWvSHC7X4swYkLvFANdhzWaEl81IAFGDeUzfy304eV0i7F3TK
YfXpJDobd5W6vkTWqcVu0tjcBhPeVQ4xyEbhZ0rSfZBsK8HYBEq/M2bax/cbRG0Q
ySNTg2OOnHTh3TFbcOxb+rTWPY4rFFzW2vtmiwb0xIAZeVtUVl4Otl68Z8t92pFY
Q2Rv/p3C8d3fwD7fwqxX+LZ+hfSV5YpbPsJPxCm/thlbJJG38gkoiBp7ZLghUO48
LTQqrdL+5B/qaDlLn3Gqt3m1Au/YbziYiA6gFix5090j8r5xKCMYlvfXF59bNyU/
pkkfaOJC9az9S7jJl8KWZCyZCeOYs3Lk/f+OAvGCQ8WAdt0FH2v2miNRcgCQBRXN
ydPxrJfpLO8jBoDGCOQGaWPoQpj2XZvRLQ4gmIgAUDmmAXFs+d4kp1Vkk850Ches
Na5zIVeOO0ufTJ7PThltxTPIFO5zI/ujz5zhVSzyqJLEYzmrebfsLDYLFUtR9taT
zKUn7E9gNgbWkDXR4ZFqBYygcYNOKniqezUorT+T/YwRHG4Zw3xf3A98En0XJdlI
gbA11ajBgGgO9N4AeVNH8+L68sBvyBy505akjtqiW5brJE8FzHDNw+j3qmhD3NN+
AkjsS3kxct7nHBVPboBmNvuBzrj4gDkqKh85POVmVKpG3Qaa3cEQwoFtAdpoDnRJ
nzVjqR2cBipcDc6qYu7mL5zhbp2eOdiGmb3db2JX2r1jmuv6RpIHiVBI1i3Th0+x
JNj8neB4snKp6lVoYIsS9CcGFN4BAwrBopbZ2sySqG0fO34FOc2YTK3oa+OHyMzh
1ukVt/0OHkePKc2iSD7p/qAHFKYl7zyEFH72KifHYloBpXvPD8ukGBlWbVU24/8e
5rRY4sz4hxAxbqFLA11ynhy/GoJn3/9Vh6ZeoXFlihL1t0NvPv+hwF5kYdmcrdHi
S/xxUMmYGqONzihf4L5jdnQ68+71nDAj/sVcgH9BBsjrELv1DJFcMWG+qkE00ayo
zF8DyCt7BPC5NsiEXTRxHQhofZKrcRKvSX76Ll6nmWrq9aHpQ6nQY9UwzhD0zJep
bVBVNz2iNi+6X+MH+PGLb5oP+VpPyi4THVGzr/qHblhWVVrNKlaiUCfn5FwqnLGI
gmAm0k4GN6j7+28pc8k0P8dT99s2mwaE9upu11uMd610a/QvSAANLn+kVlihCphh
Y0xVK/E59vuc43XwTzUwJMCVShfr6Fl2/EX3kuzXg8vZaJM6JqHChrDN7gKhaR7H
cInNAmZ+yQs+lDUkDg9ZAZNRbHrn9DnJEtEAZX2oaeB51kZ6BfrFMGo/yaeKo6L6
gsAg3mgi7UWPX+uVjg+yMIcWfF2/suf6BmVYCaj/qWdWqwKFY6RgNCVnknbH0NS7
+PpYk6ARLrRjwQrxRUU8jYAknyj/Wt+Z4sl++Q72Jzf/FiopGoz7lXOQw1VPCAaq
vPqjvDg7hrg5eXeMX+Lm4+gvIJlmqHh7YG5Xbl9jcN0Kmo5mazu53clEsMdO0Q7/
Pv/c/1CjF/7wDT7DrWXaxBW64Bh002sWtBOWeQ4jMq7fqrB+kWnQ7w6Zm8PkwXXJ
En9VzOj/95QKZkPhCifd6OEq6ORC6uSMru6QMO+3u26dbj/AwbLnGOaq72fT+ksM
eLQLdS1lFUTO/n7OeDUwY6xo7WokZWJKU1SGksWJl95EGuqafF6V0dmnvdNFw6Q+
QPXb4UyRTTAKAFMVV5ZaXcKVad8olfAxTZt/6boQyfOvHifUwizoWQOfmfX8Uw0K
mbIs2ok9+yK5XKhJ1eHLU3sV5yy7Ks8l/Gnkp6TvEs1mUwZVJjPGQxEzHpOqgF5n
f6rytk02ykGTVJzO1YOjOB/afQRAlZqAT4KvTqspBU0GleWd37QWr1geRgpVq21/
6GT6j6kDDlsbvU4yp3+JQZgs4ns5r+xBM162h3exbSQAF8iLvlI6XJLzSsdpiRps
AjrhmYDe9JTYbSZyLGoyRja6QpitT2rRzXkDePxrNkjWQQFnJ0Fj0r0AxSX/Nzhq
onYPByMN3Ri9tfIPUrPbF/0lRU03bRfybOWf5LMQkIPxD1XbmKUYbo/EMCTSzmnF
UbqR5lgLZ6c1jZXRatO5gB6b1bMYSGfy7EoRRtjpuuhdVrL/qPx1VwEXdstRUPSe
CPUJ70lIjkHKUxhw67pCrgcHGgJfjM5yokbCj8qCSaYh62YgkPkJWZ33zglXQo5u
Zay7uaaXep4VsD8Yb+0kCo6p1fT1h3arNvhleBg2KaCjQNgBCD+eAS+F0+PmjSHi
BRbHwWxiW6eHySaPmY/+Jv5uIQRTzLDUdKVR00q79TsBvAtQFGsQ7O/HPcGT9qZ4
tJQzzsehNCuv3Qg7BUhDeYUIUKy/9eRUX2HqQ9gvHnha80JZjl052PL7thCXw9db
jyXXgNEWmsGER6mNF7EwwzwUDZ2eLf6+zrCXu3I9/+GOlt+/wGWcz2JV4zEqq8Si
NSAnjhR7Ac33Svlq4qsd5/8QRt4ITNamYbDGoYyU3keIEN5azpQEicY3o/cMbbeF
4fbcuezDm8s2rFBP153aykksiMtTkeig25Vsm4Xy/na93wWnUL9GzjeSzdCYKVl7
bBlHSOKRcPLPdvZ1GP08d9IPEI2DIF5m9za8rPlIMQOjz39xEhafPbalGEwpyOe7
IXINAGjEnpGBsjHpJQPfiAEsvyPz16S/uni+Mm/NXd0B002+UFYaMufqHV4knqRl
2xf7L+xCrMk+dlOfooiauVNrWYAhhCcGJUnmczxXl++L6M0hOP7QTcCKjaaAnGSI
vFK+Xrl90+S2uWz0BT0lLttVLYzEIIBliH4eMogt0g2lMKljhlh/5axAwIwOh9Cf
IyxEpOGvqbH57j46tFwT51qfrjbmqq3YMV6RlnEvt6Imb5Luhw4FkHu5+4YcfUHv
1IyHRHj1PXjUPP+7VbtLBZLhHZ+2oivvms1kGf2hOjxDDnjAj2bx8E9qJvBnYq5O
hlAKck3Ddsi6qitK2GRxr2C/mLHXfBDeaMya1cIEMOKQdA43oG6rA6oXg4T4/X9W
9Q6f93GIS5PXbi7FtY6jdeaNRsr6l3WND0LI6LqxtQt1eSEe+UR/jyMSlZ6AB/LR
pAjMkmK/UuZlOp8JSXLFcG4XvqnZxZErQiQPyIOEGBwi/A7TCcns8VJD1FZpXnEu
CE/bnGE8izoyCC1I3UaRs7ddI2cDTSAofCch+tQJMVUZW9kQOE06z0QNH6BoRgCN
cIlfaw9vzFQak/OYpdopI4VSvZKZ1nAAqXu87LqO4MM2VfteKLJuIzCV4BTBFAHH
fDzJuwO+TDDnaa8w96ZcMhqFkJ8O+FWN/lXyfRuTLv0xS6DEK36dgE/IZDVgvLOl
ibuFEPLsKjbbJJrN3RgFrZ08g1tNxo4XTiwEIIzfJGFLtySRpbF8wGLX5Nefk7gN
3MoZhwVK/KFBgbFdSu+Uccy9JW5ErcFhext/NticIklFwLX0iTx2tX4vfKWHxHov
vJCZCuVI2AxSeg07Jbj8P8S58vJKIERLAFUOCWayJcORnOHnE1ctcA2QucgI1wGk
+iUkInjy6f8PisRKzxOZsQnsHIxOkiux+CAE5ic+ylMRLEZ2IlNsHlIE8UkwoDua
NNGIttEvgPcZxe/NCHB1vzagD7EzTDnRiA/f3Ys0fqDu0xh14W96vc81zrUcx5Vq
gbCEQQ10eOTCCrFQwQNkw5Ntlre3PVUkOSiM0vmwSIZb9dL4NwNZJTyBjJyH411r
ztAosj+v3pMTzICvUSWCHfyAtvEDt7ua0HehIa5759di9frEBowS92BeNe1R4F/W
5H/Ate1aFsZvidJrDKXu0KpO30FyahRsYx/H+WKHAzvzmZVbC3kRSOdQTcnze4vE
XzqhpqL0/EvWTu7edWq4MUuYJlr68SAvpL51MCxtV/Zo0sgcF0v6d3tN+a6VCMbY
5TQ4p4Rgc2ZAHIZLYUX/zHq3iyG7PwzxSEhLuj2GLe1bjEanD6RrM1mujAzboMP/
hrVTqjGRV28PzqmyqmiJAxE65eFo6iTxSiUGAqypNoNNkcf9ZRXgY502YaFZ0JfJ
NAR4r9dbMSVT7F6dkXAAJuoVaXYsEKSVROM/umy10fY5tJLC4hfLxnuumqHav0CI
U8K2BWLlrQQTqROJQbQYcWgeSFnqbHLktOC2V9gE9GQ12G2VoyU+uUgkQF5Xj3oF
Hu8fuTI5byV0yM8noLUjzyYPBTHVH9EHxu60xvBcs4flHk1l62dk3xMKe27vjXzd
fIRewOEuD/mixs5RATz2EfwexK9JuDx4qGC65PWEa9mCaJB8WPoN7E7Nosl7C0lY
YX6rHmI4RFmPCAoG2+lTzxBhK2P6rZt5nLDx3svaXIGICG7y+FUqyiFwBcD91auE
T/nXe+iV900ng7yPnYfTbmgwS+MBe/q7+aJzkkHZwgf43t4tqaWw2HbQNpf3w2lj
Bdv8VhJA3K1YMX5eDspjWsdfUybIhxcWc5xnyF3uR35Az5vhEaXjKPM5pbbAyDmW
dJUmMABavvsivNMAQtZbQfsSLGAWp6e/0CcxUynVBJAXgDRcxTEC84h2Sb2W/eWn
SGb5kb1P8g22aGKM1fcSuViU27obvNJ7BLG8Z/+viCo2/k3HKXQo+cbcKf/L8hZp
Tfujh4oUmeunrb2MdjACLruD2r8IzFt2m3L3lRIibZ/7tb1+YcU7WYCbRzgpZQcB
Sb95H+NfcnCL14doT2AAUNXiqkZG5ER1IoptStVAS7BbBvMxskYzzj+42FoOrJYd
CjIaHJuh5pr2GoCtsK4HZJjrhd4rg6mjcFbCDAYNZremDzTBnL6FXU8c+zaVLWZO
r3sb4klo7LDzgPfzjBKdT6hR4aKd7z+oYc2WmXomHcsPzM0en6teFf0/vXSqB3yW
8s5zzeoL2Ne78v1VW2A7Zi7ZkPCV82/M7vaeW9UFm4AtszjLs4N2CUVv4+ZgK7u9
BwFvM2o3FQsN/pG0Cmzs9ML0lhDruIqyijsLdxtpGA/bt+DN2dHK1BJLlsFW5Fk/
DeeLH3z3N4EwGXittWSigqwBMNe/nINvx3ko51hgHgNqoPFrr1yDiJVx8y9BIivj
xNENP9oBvf0aozLXYKp/DrnRUQ+GFYeSwx2PtHKwbpc93rtrgIjylYJ6A+6MRaBO
ICbTymc+t2f6QINeCmvUFrayRCMAEvFyLWnDdAWprqPbD33Cx3eGylC1lWBH8giT
6iAKXLGWv/ZfLUWQT1Fwyd46EcUx7YPbhYtHT9qTsVQf60XYuBzZnE5v4KNeR4hd
pfqzbhVUEGEVYRgVc/sa6t050b30l2cD1RngmADqd60ej/k7bgMYuPo8hW7inqtE
oNJrefpPzWFCKAvArG3XlGl8KLNTR0O3lXJQ2gexRkIOYIBIlqlC7BKr004vh1XL
P4gVvmx5mLb3eNKaZO6FvfNn/WQBRBMxUc9TrG6j2NNDj/npX0wlr73qmGpsE0RB
6VecL2Rvlcmn7KxNYQhVEGGpuMpEAEsHtuCIiigXaQuApPxwtAvLxws/fQX+sQ+l
18FoQK+HoNpH+bjGMvUA/Qx/4fj9arRbB1R6qWW9lSo9sFukk4U5Yzc+YdBRJdI8
V4hAbSlKOtpQHA/eSC3avtOVoPVAHJU9zVrkRns1xekU6YrQMhvj6w+6pX3PS7zH
njOFCNrmd/MG6vGgJbhi0v3Bmt6f8lX991okyYEzjbKXYg24/fodEzeliPDNXj6U
7vFTLcWfVDdcVjE5olA4/Np+ero/RoSnpgfWhdsAiUcq8akAQQ+dD3QbT8MUT0cH
B9twREqkjSz8myPcS7kJ8z8P9T0v7nGQEKhjCP3rn4cgpSzT1MYecctxTG8i2fsG
ztbHcFTCXWkITUsGT2ADY+K4C3s1iNY0eEvWbjYJ1J6pTb2qt+5QGndss/Et49rc
Zz0JtKybNXkg3nqiMxU/hZVUX2asHnJFwJo33hw7eyn3Ro4RvGIivpQpweuATcz1
R1BRGO+FbaCCWh4mY/SG+6GMVeGSg9YvK9qfi7xvGQqu/54sUOFaTc42XpsdR6n+
iCk074AoFCTVJ98daF1Pycy+xB/OFHE3wACYrAmjhewwfdHL+PGWaftnFd0UWrEF
OHNCiJHntLII/yeDMdheuTGKx6Ms71qC+M5rYqWHGs29kyJ0ZD53V6+LVAOW0XUa
0EI36PED7yw3QHuCQCbRbZALtPEcfrNjEg+w2uJ07sMEeNfwyA1uFjxa4MEcIG7r
leWBT+RbfwCelkAGgQsVtnTr2VxZsrLYykj3W51c1Ypb8mdB8NW1WclPhRlDSzWd
OqSbtBpRK3XoZhUwYzYk9airte4CPPXQRXtjZd9t3B6m5mw7QnuM2k4zfaERfVtX
SawM8iyigl9vrRaGAz1S/lTrwOx7YL/lpffwGtU2H4TNbB5+Agi1iXbmc3lKgImS
hRhzz0uAQqx3wI1j0o1pk0R8KUVU3RJ5tGI7OBc9/0X8b94bZqcvJ1hZ08aX8/Qe
PBu8iYHbBuktmM3bXZn6tNTdHSJmRqYF3On13XvCathfIoKimwk21h5t4G/DTYT1
lsP8jkd9ke3i7SrtK5XVjDV8WVpAqkTNYW//exOU7kgJ6GEok7F8jy8GZpGejz0L
O8+5nsKb0HSiV9gf75VcRevDxkQZ1z/uD1njwvyuYpIQI+E6+HUb4OGMQOw3g+bN
KaJCG39tlVFFiLQBKwoklIQPX6fDVEZeAPjP6DL9kJZWf+fbE1z9eC/1TyZh/6qq
lIAJ4ddUdRVvQaltOsStDPReUdZn9C3TVPCn2smlFuHCsQ8rKKHsGzYmtaRv5uKx
YWo84r4EaH4Td+yhHVA9OqniRjGfc+sfFXTqb2ETDMoEr8mFOUIb7IcDOS7qwCSZ
+cb/ccNXR03xn/oMpEAE7XdRL3GXI1GfnKywrjowcULx7FxxKIttlEHSdACuwYZP
BvAsGsiI88I5C+UojHHTZvAgwVhf6DL2sugWfR5r09vXGDktHiZI5dAw2KG+OjUF
aSakqSNVemHLpH371tu9ZnNtOQWjXRa0KI897shptBW7zKX1Rga8depSeAltBXTj
SrQPJ++ll9rVTHSFb0vSUjUMn1PBcWJocojnUm3G5xlwu/D+t369nzJ+FdVf+jMd
q0OkcdNrZ1QBIUzp4vV9OYduTxB0ydhcyk7IsaGqtLbL2+afk2pCzfyQpJ53rFwC
2rWpqJVwf24EIyaVSA3E2e82ein0lO44sfNszSL6XQhjHjMPLsgDF5dpa3LUHqUk
Ks13cOi4lggmBh3jm+KtZIpxQmwReT8jVcDimQ+kqiv/HNl25aksXXaSQgJvwT5k
XXaiyl4OY9kahveML6ZLTPgkpfsWW7C49JQ6DQQNOk26SjOknRPmolvmpBavCjMP
DPBczLlByMnf9yKcUfHZV3aKL8jyJXY4zGRy1OZvbWazlA7k/1zvUUK3lPv69+HV
cCKM5C0MDq0J2AAxh8uR84s480Bq66/736/vA7S0N30E7ZG6wknoYln4twbipKY7
KsFZbzeR19eE8E86186BEf46vfXQ0QRjA47/dTN0QYetdejq+/Y5mvCwg8VcxDTZ
VbqgkYODC7WZ1hc5hfrteNOH7kxuFVekdnYGxkV+ordvrWzctCdUG2YhsxryfoOn
PwDfuxkLRFPqSw7swCGVhv9RrZOWUNfiskaJFF1QUn1nN+8TIUwNqapYD8kjQHIF
f7zLPkj37eQhGRlhvxOW74cTHeAFZCFTrt1zfLCHMn53nola07+jZxgwB2OL1ePE
7C5R4eStaIjHd6lDRb8IY4soDKFFTZrTrQ0Ur4z6xL4T8OEARNsZT4gtqmU/ps8k
ztKQgIsIPOJUt3E2X0804GkLd1laXWPo+pyFPkc8qIdIURi+xzi52rrj6xEbB7Uq
W50qZfSaGhncstOJTkgJmCXqjGvIMFjEKmezYNQ6hQQ5JLFoTT8ePAq+evqZXKG3
VrTDHyQfDh7E4dJZZ6qhy0guWFJfus5ibhUtUCzlwQYirHA58uQ7h5R8GEA6Hmcn
N4SoyKz2y4g9H/oeTh5H0dfNTISnlBGCsN0ZkL86kkm976QNWkBQdF9unkbW75UZ
tePMZ4+36qjtt2JR7Xvz3wiVlTnYuSyRTeb/+MQtVUai8xlou6sRjt6q7Y8/mbk7
+DvQESDSjCt7TJA7/qn6D/IY7QgbhRKKWDViMNFDFMtuan+e6Fk+7VoJlt2V7eNd
U/bGtDPP7+E7Ax/F5ZeY0WJxia7JP65Aw9EIsaY4SKNk4oJBnplVWejpbM3Ve1Ne
MKQ7uUD2cg1wp4g8YjJH7N+C75oW+vXBz7Lr+VTwXH3BeVuAeiEaE1mwtvjgJN4y
Wk4Er30t1BCnUZ/knU/VH4L4R0WaTkbhih0p8ZK/gzSnxtkVCOvP0ZvS635Jqz1+
OObBXjt+zkIXPx6A8dmLXJY3c2rEurzK7oPdpTRfOB5djzY98zY+chThilT4UeVT
9kZTBs5luEKXHtO/UnhDM4hizj7ZForYRrTLzgajjIC6QA49+SCsvg161kk80K6U
83lhZNM9UJqkk6pfRBqetnCsQvyVV9t0BWr3hPv7RTa90APetVVohG0Zg4kW8GNd
hk5mOW+iCoPNTPDsQcYFhiI+ZZfrLfRrQcvq2O8OgreGXdPGRgJniCPrsYvr+v2E
SI38yHHRNzkhKQbP2WRamm8UWLPzvpv/xEsf2aOoHatH27rRnNQDGsGvPhVaWHA2
T0S5TcR4BQ+W+tXOk+lns1ao7fQFP8n8PcXmaglCr1xCUAOmo2e9aB2zlQy5ZbvB
yHaJlP2QECyhRnjOlUg40vAC9rugU1mmIw/v8ZGGLBvMllhBLIbQXsLOlxA/lJ2k
MOGxHITc4T0Q09+LXFdBo+k7d3fI1Wmji/S41QloYMKB4SOP6t/t4oYwCyQviwjg
HEXCzVaDed5iz1vw/eMgnR98Yg7+Jk14M9R52MpQo5T+eSfI4n76Eo7gHn1JWfJG
z99MovQ5fEGaSxjvDfYMIyHft5PvYzb2z1QDk8cxjuMgBtzFsxJqswwwACjpW708
YUqx9bTbmSPLrb1UhQOpvejY78DsiP4XT4NmpNVusFTxYnmCK5jsCIwZ08X0ifgr
DuEvNEJmw5kTZ57j3t0vRNrE2dkdv1Uis4Wxi3zg027iLhQVKB4kFBHGhDPBhPYb
xjQVEwRoj0vNUPnbpJ/IefUyF0SxJGSEmuNFskYNBEVirVkZqe6wPSQU97w9V5w1
MDuOH9GlkxOYqcLceNSMnEe+SLwvTU3ZbU+2UmvNpKw8sJdiQPjGXXeHP9IubFI3
bf1UWQV0j0hu7LRWZH12oUOCDwT/bIxqou3HWrvQU6RCus8+YYM/UoU4ZEFDIsFm
sqfBPa419Pa3GiZolByI+ElpUT/Jcawt8xZhbkq4Iy+UV9ScWPGmDJyY7ZdcsaJX
3KiN9i3CyelB/PI3xqFHekZAHPrUhKTvn06LgegtduGa5pBIbBLFtMwgcTDoD9Of
QL7si50EVEDNSMOVfaNFwCxl0VwtuA9fJkR/XXvBV3bPsiVlU4k+hOmoGl8XjXxg
z16FLQ3hVcop5nxpsY7EVRXULWrwm9ug4BIzz0k4Yjj0mpfcuWsouiNb8mHliVpl
Iqylzo9KsKqtWJAyxvTXOiBtm7S9IxH7XQYqiSRdStMa54tmXdGC57p+rwM2ITGC
a/FJGWvloJ5ccmrEjTU1KSdGKPlzggCgIbrztED1o+Jb0yIVcHVimVlZE4fVAT9U
zKUJoN7FDEJMXdB1WZGr1d8lIoa3os7TadtTMcfYfWGjfAgs5k3DyejzZ8MBQMkp
bNRKYdNViCTpLkLlY1o2XLgspyAhkwDfFk+svuZX0wSp5UmaWe80FFoA3/uTWQpI
hNjq/cNmsesv9K2SMCdzxXJpIMqL6PPzqPRCCrvM9UEpRlzDajZgOk5l2eMnrhuq
gz0Vq+aFIyOeRkDoxohpmKrzUX1fTDgPF5WL2yE0VQJ27moiX9m5hjj6YXNjxBiT
InbF/ryBqZ1JCOedR6EiupIfEZgKvuL8/p8JZHUuqFC2KoMCTyjRwsYktww4bBNU
M6lO+ArKM1dZ/iq6LxG0uL0Akni5i1fPt6cZ7ag33Plryt1RfBdEghRzGw+UT/pl
2R5LXHdfZDThgyAmj4/YwhxeL/fuxK8TJeOLCq54rZFR8qlyvwiiXgNZeSSR2vDA
iQufCyz0tI1YK6HUgymq7YzUYT1BBa9c0QqCp+P0yjzRf+3jqpYlG+zIuNid8GQq
PYNMsj9IOH+ovRC0fzr/9u3bsUkaXhXSUMlIM+X2VrfsFbArNSdFmyxKRtYKGXd8
7jCJQqcPj08OhwrwoE5viumZszO6naYkGeNEpsA7VsmyEjSnfnVZvZflgsswHFoQ
4poVISrOXpDxn549QQhsy0F6fw0LZQZYcQCcpqgaJWmd6iBT9CY7Yp0BWesmSDTj
sM3n+9jQXT7r+ujPZi8RpIIzEPo5Zio/Nn4RuUkCDDunko+xaw3H2O8nxhmcHQGr
1/O/KmIHoKWzvrM7wcWgNzTo7DCiebqLjoYpgNpKvzq2IlstlUbDfuUwm7juj85S
dimXxIHvci4rCKjvDbh9MA+r/C/XRRG+7kd8Gj4Ep1B7vo8bZy0W4aUdsIaZIjnE
7/D0ESTE5YXbej8VUjujLA+YXS0mwVTKq2t9YOx99rtups7Z5PcH4yKazIFIIZZR
+2hnO6z/j0ykx2fJ2QGeW0bo1OvXTEjDUpcTaXBKjSiwXSfTchs+8T9f3pCdCO4h
+Ol8YXkkXrhRhK/B5BbgNlnnxOl9fL463UqUPz2bVGpycLWsRRRHvS5mLErYWalg
Tcl3f+vSxqGgRD1vw6Wli3wOMy3ObpzeVrB7BbjEDKbuoVB+2+JtJsMlAdrZjVSJ
BeO6U8v0yqpy+E81jNznNqrAfLy9jwbcIoYQCEJ0T5Pt2C95J//ihLoTiF0C8SK2
cP7P5vvrTFPaWEFd7mLn9J3RFqp3gC8e+Pz6UTI4XFOLyWJuVe0O9YAbLfWuWhes
kZo92j2oAbwea0TpuNDGtz/R0v7u5XPJlq2k+J5ZnjLzLI1oBXWxE7Rp/zzNHtHU
klMZ102BSbc8acJyhZw+mmRIR+rbC73o08l/00RfztNLCRoEGBsGKPxsmsS4rfnD
S50z7c+uSRENLZCG7jO6g+uQLGmmXe9rEFVMMMogLcFaFvmB/YJb8epHuZa5SVBj
vnHskf8bH941Wil02ihiDrDZz+JngWZScDOv61Et78fxrXVX513Z7bqmgI/6oBqc
dv6gOjPWdPy45rANTciM/5w6juJ6BsiwsZnwbPpJWvBnePPM/Ebs2KCOjfzeRl3Z
93Txhsur30ffQpvapKlKLP6z84TNWg/cgTHdnSJ/v0+v8JfcZN9RD04MGzP5XmcE
Uw3LeGzDPOzo/HsMGRvu2Ut3CijntLX8mE9QbKIR8PeQl1BgO9QsD6jsakA7d0Pw
jxJI7+l0zMP7bUM1BeFl1apd67WaTr9aeiODeZ45NDlCr2knkBoq83c4J+4XryaB
FpZQVA1xzCLPtNqDv1QWL5DwXH9rDp6nD31kkEMlkDgtAg3Q4HVHbZ8Tq6YSmNDN
1v3TnJ+SlvHFXb6N3k8cW5QBl/ebVEfi9oj/l+Q7XNrGODc+wCjC/mKh8KHkrkgg
pNmRBXlp7o0aKvzumGhhXDtf1m1OuQLvLM6HCjhTJmX9JwijMdtnLsS3moYtKSvm
fS3MOGV3OFtRe4sC2fcdSz7BP2qqvxqQx9cC3W7JnfPezFtqP9uGG1nBJMFrHD1k
rtocLuZFDx8cPQqt0wLd8hCGzrLiQ39bKLH/1JspG5O6hoNXfGImAqRQVCuUtIrd
Fo9TFFoYZAeNOsW3eoihmx5mHMTTI7xkNGxZIOofz3gJKYuMhrEU1Wh3h3c+YWC7
Hv2wFUX0KxNGdlpoje6V6vGr7rOoivf0WPdBBLAZqKmBKmaPjzGrli4DAKSleJXa
2lNxHUyVcjYDXGfVec4z9503FgNFc9+RTtb8FxxJ53bL8LYhLxK90fm3XvpgEeEB
vKLksFd8QEzZZ8wHz/22orH9g/nyJus8vjjMqrBKTlj6qBnFzXGxcvNMMgnPZnev
U0yxkxh7wa5jOwT/Dai+nb2ph7/xqcCP9OqeAbDSyJ0hnrQJ2+AMUPl2MIgGkkdw
Iro870IwETbEA6uJGfFHLhzkV1PtxErmIBCCdEGFv49zcgBKxZtERHveFVaWzUZ6
gYZiGnYaBwuBi8B1MmYN+rrTQ/YD1MULjMh4ssUJhbAc9Au0eZvN2ZXi8rPXXCp/
E4g/5jWsL1M0n2kfi/bmGRpkSUQiE6eF0LG3x4cCooG+NPDXi4wYUvfNUB+NF3Ys
PZRssEjS1hftYEbfNfR+/oYkC8Ut25M8VsRkRtLGlC+cQwL+dCc4ULXpSRKSBmX9
ucM7O05+byzzLax7l/GWzDpyk1GYYQ4/yzGc4JgpW05PdmSFfpK0PrjNhz75ESwW
1JovpTKiqitdD7ZY/++y0MtUeN6rrVGUI9rJJvM9asCBfVH3/B/zV97z511pyHd0
qs4Ygg8Nia5JUfpgmXmCjX+a5AwrBghOisWxUAWIvP2cW0ptSEBjRhiqseQYRgdP
EeiFUg3s7A+/S7BVkMOU393A3DGccx1FR0naxEnZNP6/abeiW/7ZWn/GLF2gBhAJ
pzB8Er25SSnacKTvVrgsJSFKPwsOjM5dbiwY/lnYR9uARKNRGc+pWp8Hdhkh8WBK
SW/bkUn7GFgzQgzzyJEYhBv9gI0pIEg7+H32htdB597ON+Tf972QXE+AMZ3F63NC
73ESwrR3m7LLQCAqvXrgd5nxmJwZT19En930vwedqnmJ3utuIEcqVkUo10u/fKpS
F4MvdGkR4Tk0qrr2nWflL2pDPwGy5r6mFCaGinKFQe8m/6wBBxHlpvFvlzQkb/hN
ojYOEtymQFw7B9HYb9jBIwO2dJtAanBHbE2VPYEMypvbGfz9uvdRErR+48pZilnA
kH9Mx6vx2jP8jDf9rErnXG6Km0oTd8bJ8L5RFZjpJzqIkGO80gEfnb0YhVN6F/xf
JO40pTyz8bR5EMaRh4craIccp90esSlBe1zwG2wthoyQH5OEf0En61Xgim+5ldPS
zhbPGx30yJD0G03Dx0qmIq5EIgzzwZB5x95e0Irryk/afX4EtELdahGR6gHGW7dx
NW43GCaIcEWPVQ39zAYfG6tnN7xOvJm6gF2VeGXoTKY92x6s1vdD0WgYf71d1gdW
TIxZPQEiRytmnunEffCn6lnbjW0r1LZoYN4oiA/yamSED+3XLSxU8I8SXNXP3snP
LnWkyJuJO6arv/a20lzK0q2jENp1d21nKBj9eKESax8Wl17cbYJuPKnQ9aC2x1xB
tIB1MoJ4PV2Cp6GnTyS1k77bzSTHgrDi/qD7UzMaYnChSb0NO8kHOnKOJ1oie587
TombZhD0fdN/Ac+mzcWz2kdwCrV0ox7FyZazyCu2A8J4fBqQJw7QIvvLgsX7AkqX
Mt7GuAxSMBNiPmXVoZDjAADFTCLsnhnyoepHwtuuxlfpSB9+prGu3yfw6BipJV3b
SAxcpQiBnxvXijYml4rY1p7HXniM1bYa8CFFtke5frBcr07aAhQs3qMMpwoBhGZ9
u2tBPqjakE7P/GbIgxB/UX+uRrL7p9n+z1hcifbZnhGY/u0/bKhM9L5HzBK1o3Ee
DSaeRsIgimwi1Klhojb8GR8/aMUvm9ijfxsdBkIUj5wsDdMbwK5J1DkbdcKmjjKz
2Wv7Lr9I5JNbidhL/TENKU8s83MgBiFcoZ3952kqO0cdSmGkirgounNpXHNts0Qx
l0KSoq3KLs3xtBb2TmvfpuR2kV9Ri7owhUY+Ivtai/jAubTIyWyyvSdaVXZns8Zq
cAT3AxRMGcKtLpF5/JJlFOBEsvvD729TltebHiI7hzkPtfAR7uydr4ZrXw4fSlgN
RZkxF87gn27ENhrpavHIG5b7VEjHsrnusRtvxPTUsb45i0UL/ZSZcY+GtMgDBzOE
rRL4Ru81UeqGx+BrUiXCnfrzdaubU5zjllCrQ110Js1JH//qOY252vANtPBlH0RY
+PmthiWZ1iN7MPTv1BsVGWRXwedlTG2mV85aBozJjQfRsDtk8/qXXXcmzSgzjzG7
HWXkZr55iWpbig/hQimOzVF7m21fIyMPbZuJLnDafeG3gtdRFtEQ2bLPiH5VomiQ
U8YetXhxe5E1/X1S8w0XvL5q7W58fssXPxJHY53AhwD9eGHLhCiM02kgtliKxVCb
/Moz0dLTnhbAGkhXQ/71vSSG3EMxAAy7NnQaRn5lcz9cvbtWeC3vYJFq4D5/ITrs
bBneIrfE18yx0ft0UnRtGqnTUPGHAm5uH1uwign0syxgAkPpcXya4iJzR3mF2JxB
9vhDn6l2YeKxF7/BipzAK0AzrIt4eFHoIvMIxSRjw8hy4zPnccA6Ga1MjLsiICKI
PjT9MvTV6eMM/6N4aGEG95z0vsEwh7jTHDY19VwHxv9qiXzEgMdOcAS27l2l4yRF
K6HMAGvh83Y2/VUtYG+ZLftMR6n54EvqsAmj4jR9BLb9J1Li0LGaJBtkoJJ4B/3J
uNK3qmbYNvVo7ZWiOHvYjDjrbqzyfqCqzuMZ1vKUQcY6/ctteMTHeHMwhcQFH0KI
B+CKK5qLmZTNtCvIBeJNf8LNiYiz7pNFYvv4FS00SlBrPVh+NJjYpmT5xzK2YQci
DrIVBp4d5VAYCf0TdKxcGsuXl9B1YUYaKBYPLCFxr+QcsBZhKd5m+IIMm+P2vQAN
ZPKU/4xhrpc+Hi2lvvkF9VXbVuRJKlGvvmJ1NcQmo4l4QFCCiAof9jVi160LYPvH
moXMhrS8L80NzzmfkEeNpjubVb94TPDaiWOEtN9bIDX4Vorou50EmHS0Qt/Tg4+s
JnulHSL3NqcSG0dEWl8kKyLorWMMCSbk5YUEqFmFyel4qmVBFklQLqu8YEUcHorv
Oelo4bzYJeojoBY8pqXhysQnybruJ7RxNfdxZ6SIMUOHrnK6WoAmrLIyGAyZ2Gbc
z1K3YShYRySzT5HMS0CXtqi/g3ung+qFU0jfBkuOaXBwcGfrfZtXRoUdAtX+WX8J
46bPvHpOpneggO+vdR1xuEmkcPc1Auee3z/AcWkrMI7GDpRo5JarHW63Tmbh+g/X
o03RgKP4zeaqi65n/neZoGhr5o+VreQW9r5gg2EtoM//4j8izygFam0lJO5itZr4
imJJx3HhhXhzYTKaQSS/GsBCR7DlMIKb7JijgXmxZ6rLSYFf5YYI2HW2oQBUpavQ
z2E4+G87TE652SNlVp3BZKfqTAgIL3UeuGCKxLtYEQAjzWJit8eHU6zdI4nFEg56
YjeKP+bbSp5qSm5hzJptLhwEEtR0zi7jNQ98vdR3fvRqz/pGfNWWvRMBc/mnAfHp
wMVA+ok3Wi5xHzAsGYxnIZjBW3QchNUTkN+yc/ifsTdPdGkzOZZ0QXqyVCgSdro/
nphBAmqefWdphCzy7yVy9GeXHOuz1BwAB/SN7N6x9Qga5gmHf6tYkyW2TdkoYLV5
J7omdQL5pjP3g7IyvBjpk8qFWiCE0zsuTCJfo3W3MkSBqNXwot5kRlQNlBKvuIE3
3UP+WuQDmioFP+s6XfTH5LTG4eiuGgInJSn8g5NWGJNil4R5lVnddt9MYrJuPhN5
6rERARAROy+4aFU1GVadD4Ee44YtIFbY+WRYQNUuLx7kJ9bNhf+d6BS5alTLsx53
V5Vp9XzCe8Bm5MFA54JP6Eswk0gUGHpusD7VUwW/JDQDP/w0696XkW0A2CGtJu4a
XOMl2iD9nH7mvLk9fVaAzM/BINycfJwzp2TQP0neo6vFksALjzpgJWvMhinV11Jo
xxerwxa0W3czXYjNGTiMvR9OM37DJQ+UGNRXu794onWrevs42f7d4/Aco7Tm+kb8
Shx+6RBicQmCf8g08ZtqxnJwvnqY7yvS6/AseCI3ptsuCfhq6DnUjoKbJaL1Mqck
fgars4lDCTKa0Qmrn5bIipUMHsdj/oBTsOYN8UmJpNvqt6+Knq4xFJuPtgBfgcJy
VfCYRVsiu3WWH+WB+zdiYOro1ECKPaCdQhueD/9E3Am1RPGnNncPySq0VbUAPHo2
Mzn1EeF0mpH+LtDTlz+h9eeemZCwPZ9MfzJB5aRyRACPnTKJDiToXadP87OknEg9
AztZ4w9V5qEPrRLlHV6mtfo7XWHGc5FPpFWYi8/fxfoJxhXIdosxa2BFlkv0Kyh/
gfmDNViDi4/Xj0Vfow5J0Px4gJlnEaZGHWf0lpzuXE98QbW0tB6qIXMVlJe+5vt5
/J2MwNqHCCg17Pn1CaGZjCtV3oJG+DXFom9h52+mDuyenf6l1QjPEJo4GTyPNuyp
t/1jfyEqfMNFGj73H+dEj5viFTygvsBWTqFKnTcWw4IxoTqhVi161tZPsMIOf4Fj
K5rV/TKzFoFv//DrzLfdDIywK3e5kFYtGKAubAEpVXO7+Zc9bnrqi2EcOBAVIoBJ
3J8/QbAgbHxGEuKYyzUgfJsOgyNEnxdYzt4eTHA5UEBmC0cjMGLVmQaerizcgVWi
G3BS/HMM6FdBggq0PAxLBxk1sbkkj5HOu7kXeBGhCEQSp2mTvvyS97pePCnrsyT8
B/DsxARYKAgpp0iuE9WS0NhJdwDuvH9kDp5KfZW48IZb3NgAW2N3f2W8/TelBpz9
AhvIEGgUtNn/5/iHWvtoID+Tu9GcGGveWPp1pVN3dczmkvcY/MYwHSmyIk4Eqr2y
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 33072 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
4NAZGBPmQSC1EoH0Jm8NyN/TQPWVswvUgi7BMpn963R6SE8jk65pLN1GB9+9dedp
45caT5UxFmD/SqfJCVNLL6ga1HqOEx7QLp3bvAZrj++5GoFvkzw54wZkyyCEy2sP
N/3fnNqdJPPKIa1nzUnIDFDn2k0cCD4MEY2h+EOH0GQS0qInIKK/1BjmLbJHors6
TFrPE6U+eP11bnJlBU+CMJX0R1h0b3/cWPfqGuGx9dr7xybwZOO4u8KONZ8uTOJK
UJlAxX29OCF2I3pijBNmvBWZazAGRctpK76h3lzqEYyGF6m5Es58Lw3dCh1Ggu9A
HRER2a8KWO2E7xt6lGXUs+/HW4c/KDy9EWKdgpwKMA/ySRDhyTswyHOOYqsZNhIy
dgREqzQb/POI24yN9iYq4qNZ6pJPsRtq4mjw0U250OXMz1AVYbKVsma9zodQAZl2
tM1MEkOg3mkh+O0sI0RmhAMndZiIGFgXT3rdnmgteuI+yI5c6+HxJ9hjcHDwbbRD
Ro3ArEuk4rvYB+aW5i/kngJ/yCogItfgmk8UlI2JA54uQcVVSF/6XwYtPTAGgaLc
M/wN/e5Hce6nKFyUrmyveIPLe2dnTCqn+CptLx2saVYDzzlAm5DgzI8+IRzwxacS
xF+YWoHroE9KOeLCGstZTuaZy6OdXRGiG81+VNC/QA+75faV2OpoOGDgfbzEMUv3
oinisfkpLVqJDIb73xV2eoznyi0FdTQKVjxqqO1qMDwRTtzf8N2k+OgXgEh1zDUL
aTFu7FJ/EQOJGFQY5KM7rtKESMkZkk0/EmL73/oIjkLJchPVh5+EfjbpSFRQGXD5
ggbev/ztNzvTrvPVv/L/FOusAPq14/T0Lp+V5gwMY7i8dCOlPr+JXdhHivfzy7pK
5Q7q87Y/fT9Xp9oVtNszu1uoe6RAZkbOYkz9b6v1Pc/Hh8vjagEVRCc6t45u0Cr7
jiaJZG9hBtDEiDjJWP/Fcj46SWExkEBrGwzDkg3f5XbwLtO9GhNmycVTYHvmzGZI
0m/OAy5EFqNPq3nGIuB14kdLvTtUnoc6dTJtsApUEBRm4R1/XXIWKCIYAFu1lkF4
QlkVFSv5EV56LdaPxJ000mFIKkd9s7crPDsJDSnJTpJWetd+Q1GcvNLDfBBNrjco
5i3v2FpcMssqOv6nhQNipHUwQZiXAsX/vNjH+32UNP11kFoHnjhXNRMCjIDWpX/y
zSQQQ7yScmn1x/YfikRXB/2lFh3uPbMwZzTUukaXTIqGT1C8WgjG2A2RTJ1p+RGe
hwhJ1Vrp1SH86F20/S/tnZfHLyQlYC01epo5v0UwAyAEPq/IjWvduFCRDQJTIeGa
q/j47Ac0TznRCYhn3bUqTRM427l+uFHCtEXCmRujvZxEFs9BEPPTHCrUSF5KXnpU
dk7EAjmoWHy5J9RDhrVeop2DR3Uty6/DUaLNKGb2eap84Id/3MrkuVkAJdHFFL26
kuBGq/JNpiDXb7YC1R715VXQlhJDuNzLNxD6+cxdbkmmDtwCT5jeUBsg9gkwJ6la
2CNcD9QgPItrsBg6n9m6NHUCfucyrZ0wzVkVNta9kKVVM8X2eHmuXSj+WZ61qhGM
t/qKkDFDEv6Y8gm5IgLk7zs3pa9Nix70x4ZWQK3vl0cq9xdGiBjl3EnEweEuFb5J
7jrH7gsnWyImI7pEPV1rMjDYUtUCBMajYNK27cbVb05qNo803uXrR4uoAsBF7Err
XT+uILTLxOC5vsRmt7pL3A1CnMSWPCDH5uQWijltJ3BFxWJm3e8mOaqbCt7mMcyW
jYKTWcULs+Wh4jd0LsHUaYYP6DvkDZrBQXRuRj1uV71PtcbCRvKg+0HZKg/gMUKw
e7LmTr5w3FsghBdw+HuA+Uk958IuuAQZddB54WWag2BYKqwWjWLmwsJhbe1MdgtB
DiqjLhQizi51nHd52di8tLEcmqcKToFITcUxRd5530P+zmv9fd1m4GrusxNpvTNG
erFlV8KRe5NOYcVaDmZOlfop88lQarFmYBo7Kg1Krsl2YaBB58LDrVKpYnSv06cr
4az844YfECTj01k7sTSmcszxInM2gPabB7PZWq9JbE82qEJhj2oNXSM7og7vJTnZ
WDpA9fHOg8IiaMoxj/sQgUH+rj2JcIeZezUE7lMGQQloSdZfMFBe2NMhojFmYv5Z
3rS20icC6y471K+UlhjDdnED0uuiAB779aSMTucFJML0ti0bFemEwrsZ2eX3r0cT
/kOhGUW3y96B5AVdYxfULXoyjKO8vGxFICT1C5xXnN9dhjgY1vCqoPSDHA4BGLaZ
wEkxGhBnrLiRa3DvdjIgN2hL0z/0flbp7wuEAiOYzxRq9EFrJtn6YDekZ18ZOp2a
0ED6kIxypnBuAGCq74sKXvFFHjUInxLrJP6cNfY0Rk4UnUzrI6Ut8yJkO88rkMp1
UxK1KuYB2VU0xoUr1/9ehfsZf0XB5hVBqAk8gBb4GPWQ9ajt7nrJMz0ncHWQid69
83VPx7pQN1L+M2kRsLEt905jCusVcT+nloKtBLfQZvtVZIfspDMSjuMQYLyMwPKU
OBczk3I0gsnwXxHWS9RzFj1SmE8y+3SqX1H4TCof9NV8Q6bzokzOJKutOIXiUBAP
5d3FsfmEumiaybfl2XkZt5r3uVlL4GoeCJQNHK0m67jWCGYUs/hq5TMdzzpOPST2
BwKoVnpnR81WQ7ZT8NtnrjGRWkEZ1wRy4SvQJsd+B8131kRCeGJzy+DGh3hJW1wc
8oCRP+pc0vVho+zcFJdBGxWMXscn3ewdcs9EnuM4V+tZ1M3/o5MwtDzbMhsYAwBh
FQj2p7L9rZMPoFxzdAtlhBZvKJifxbRFdKAbPsxX1BElS4/uE/wi+3cQK5WCvMOE
0vNnflcMcmvnY49QcZIPGJmULyViEWKd+aD1PlSJ6+7FuY7fZrqL+n6LbulSw/Sx
fd32qtMMuNv/77tpqRfU6bIV2cmxvf3+vnAvkFXquh7/kO+0XR8oDecT59FqXNbd
VvlZAPVLsup/LR8Ny/bgpoMxbsrZ/1XZ6jLUPQS53arPhbQL4c4GsVS0o4rk+KXe
saUGsytjvMsoptfujwN8W8q+qwdxF0a0Hl3WLBzOYhFowU8dH56QAr4DMoHXulSu
4075IWX3efz8II1wjzSOo7gVgj2esuMLrlKO6A6i5Bjs99pN2dai2yLXhSCVhmlE
+Ipxh2/tiiWFsDME5n5xa5J38ixjVqFpYX8kCfuIEEqEEOcThquZUb0q6SIgAbGJ
nboQcQ58cj7A2N5B2Lxy0yrGOb7gnBFGNoi9LdR3UwwqlGnXhho8FIx4wcWHh2sp
MGgKDK510bZBh+FfEqoYdZ2E6XJBIlBLLVInKnWs9UISjlo9egCcBRBQ9QzvwlKI
/9ahPrnH9eAZA6KFGxTrS1XKG7xmMZDWqT/mYQKX65qLJUqMw2XSnwYmLUuFZaWf
vtHl65S1thUuyVnQ9VjB//9xCfycZG8BI14/2m5LM2O+mK0CsLkv4dEG0vIvjEts
n/AEfvFMeUtVEv1Xa9lV0xs1mmsKv+ltdnpQimNVqY6t+33F86SP8PNLIO1PwoFT
1avLs+ze3gwp9ry7RcsaagWgSbw3Omn85E/bdFcmdtSIdBvOwObL64G5PR1wBWf8
5C5W9WXKN3rOO/tGpl8WLZeCkqOtwqzUSkkEs2ma+wndgXXUnehpSzFeZ9ure4aC
v+eQC1A0+GD3kQn0Uu1xno6LGYw8J25WSXUJ6rnjyInR503fYfcKiAIKGdon/IE8
RhUKk2JBiuz8dCQjA+oT2VfsE3gdLtj89hEbq0i/hEJZL62w7aNg0WX0wLOx2wOU
LJJA6xSgDqxeh707KjJ6/cfrO11P+X3Vn98yRktA2iJ7aMQqf7hSqqRJO8Ixkloo
OKZqgYqj8pakQjc1uD5omkw5rezMH6L9+pWMACwA7Kb1YvtWG8Wdm1zvbJ0as7A4
82Wh4jffJyYbK1YYuU/28oydd4yzGrjAabXwwED4mfpcJaW9ZIp5QKhL/Krr+DAC
zYg5TOt/P7hxvBCG9k38/hIhyYR1CiTJ0i5slnO/RyD4YBaziF4vqSFltXLma0t0
XsAnSIdztUcUbubCGaiFdH6LPOOw+EyQZr2o1n6+oiQ9dvhoKm4AqV+lb3j3uZcU
G7tp0po5+KEnKCcyJ+IEnYHY9gr9dddsqWIWkPrcUaYgZimmFjUY/EBqUBTq8zcy
JlPR4zbibl9CpwUL8nwuQq+F9wCHGwowRzlCiCWduIg5qoz6uXpAIBR5zuwHqBZE
f5YPq+5Ut8ZYzYd7faXy2fU56CEUkO3y6Crn1a+qCYxiZN8VBdulrB1uSZNTB92F
h63k4ztBjVAA0YaexRmnbKCFX2OXrjrH55vSKgunKCyXE723Ly4Z8Lv9HHS/ESI3
B6YskC7kBw3WwDCvqI6YYkQiI7pJbR7vA3WoPgKdn1BQMD8pR72shW3An6L+2Lae
ul6bWcN0gXGtess4MRQ6ov/i+UVowsxhdDlvg1UJSOHzh4rpcZdncDAFeyiAP6VN
A8QcbEUpLyACGwPg04f8TTpa3mq0PewYnfl2NmDVspdNzSS+2v+RS+EcL7cCkHsS
TiI/uAFiBE1TsdwIHtEbt4sex5OQH5mzO6M7FNwBkD1cBPeJ+yEv6Kl0/+tXwArE
vPKOB/pzIqI08c26GCPSBOLDXZrUlqV/OKWP77m7I0d3JorI1GQC8gkZhhK/5kdD
NvKTk0u4llI7vt6tN5VCkOmSuw6lUOfAWrqXmRcECpy2pSAcfezxZDbtFaA5oh97
MqXsAL+NY+sZVhsGYvIQy2AGEAf4dld6mD8JdijI0rurfAhU7ArjhkpKX8nrk8ez
j5QmDgyS6y9oqv3SNWe3Z5IOjq7fbrg+HRD58EAhlu/xlhjkE7Tm4hkGbdjyUFiE
Oxyavv6alhCnZO2bJLPsm+SNCmicjD2Gfq4Q4/cBcFeU9utzXNo66TO5o84tqyBk
g0UV15CsKOjJSKGJTWFxuiVYBSG4Rfhp9QosZ6QbgkwyZ+2LCkvtOGS2nT98ysIf
iF8BW35GpTNIQomB+z6F8hhJvEY4QTt3m5qANeESNgtrmJ+fX82B8sUVnfb9deQI
lML6XDlRPL8xSXB0eMSd920GXFmezdprEZ5eN9mWfeGR0P70VJPckxDABrC5oJGp
MzZzK5D3uQ1PPOEYptq6+YD6KhJzOfm6xkqojQPUsj1wUrS9QZA6u7Zo6Bwcn7wK
pegGHn4a3se13mJlsoZ8O+o5WI6hRK1um7l7hzHv/OMxDvEUMsR04X+qsP+63616
WoGgpG/yTziggpPPXyYk+d3A3qH6fQYx39JC0y0/a8VzNVvzJswstkLXxHobxEZ7
FzCGDIAU9uQkBxPEv9rB+/GRr/bijW/C1zAEdyc5l215zrPq1sTa0/GDLKl2PRgr
pKwgAhFiCAWijaSvKm+lg6QNRWaai1Nc8LD1zSH3rnQ9xf7BN778f3Ghvt5KcJAz
u5hShD6DnyJHEeOWrlPwCPvGG+Z00QR59snufJ+4sY/WnBi4aI0XT894A8ACWglF
1fLrQ68L9lwXn66bxJ0fIYnfDlN8tnCq9dr4iT+/C2ytrWjqtwZhYYyPCLdImsPc
rej47E8/JTY0o/MOTZdG5xB0RreUBy+qXeexeQ2m+W4ZnZPx2pxqBgAayY6SGvGH
qu1TgF2PdEUpmIl5HleHDaEgxu9OqagBbAvmPo3UsGQRH9MTdMYnZOBLBsiw0/WK
T2GdD6ybOoxSoKJSqbCGNShDuGtv0FFqSia90PVnmpCkBAj6cunu46QcNFEuefRr
fDrbxzTVKknVfoAfq6YFCvJDzW1XEulXo/Pr1l2g8mkOjY/994UGfr2h1mcDop63
aFL0eAdF6JYqrrTNVSHR6GS5cNUavyp58wi84PT7RX3PXlVifSINuTj2TXm7xDlb
CnQAoi7YEKYu6v96PTskxzS2DxsrmAKOPLCiYF/q3mMWcF1NQBYIiPa4+1J3iRJ2
pnkJePhs4XakSVGf3+BEFcXH/lIy+N/rUiyNozUfM5i1P+2GjkNiBCq5AoMVUoKc
QITkIWbXyWLzFuZ2gmoJ5gFKg72O6cuQDecMqHhQdyfKg8kyttwvgE+LAELrutHn
C0phiAX4+rNVLOMlNekf9N3HNT0yCSBdom7N375KZdqN3zG5FXI9bt+rJBXy85Mj
oE46Rxn3hKF7FyiZDN9QIXCRbul+OOPUrhNUUqelGKjRNJYvYX4KPgGDbUrja2ne
jv3meC0kA39wv1C/KKmmf5p110mPCdDpVIRRMMEHx51ONe7ODNxSkEX9r6YmrbQS
43V0tyUJlP+BA/Wu+Nyi6PCq/1nLlAvb5QELVTds8Z6LVPKeEElM4CYv7h4GGYMm
8RVUMyR2HsBeeH1R+6+NwjRXhqarjLF9ACAyB0DIllY9k0F1ig7pu/m3sEKTxQFu
qlELoO05FRJgqOvaiOx9YEfhknvGRpm1IZJpb6tDU9wdXj5U0vvyIJ3THPr3Pk/i
IgSC+z3awh1AFj7GOz5b3YaRjsYKBOMmG5ORnPadVaSjChJnd8s2A5rJ3p1Zmw+B
FMFHQ8+Qvi+d6+JelE7CFBlbKhelusvTaCaRhtDBOWAPuE9j7IyTuBN0bpT57QT8
8R5bklplyHNT/163cwoU9UFyEJYklwhBrXmD5v+VXozTZAOayqcb/lnuaHjYrD1Q
wZInhTIJKd7ToIetHR/zvlWvyNY4GXuOF22MtKcATdTpUiJXVqgsGI0yQLI7ZCoy
i3ch5zxGCMviNjOe3rbxCU/oAqrOTmOf5onaoBTfspdH500d1hiSUic+te2Fjaw8
iC9l0hA0HX6/lhUO/nO5yeVJ6ywUar4BDXnQlbIXetQ3iz9DXLmErSP4yEWvCC/p
Sf/+dHXs9zw3FtF99Tshk3VIAbsuapRZ3bLeSPFpa1AAAeVQdkotdOo6NhkW1MfF
wKIgj4ov44lJo2FyoWgB1w5flWd4rqw9YOWVqGo2/wryb8zJipoUaOnWfsvV/JYy
wSyqvDKafI33Wm/ZQqUDW4aMYr9emnXW7qmdKPyZz1FoHd7+c64kn3zoMHwwFBJz
u9BrPX6qOh4n40SjsNQBlA1zK5E1vazd4JYxj8mT+WtiC0pIo5bpO7RIL53Q2KWg
Ci5Mpe1X5OKj/hapdJy69fLGPUysJ4FOYLkPANygNg1vU/n9TTSLakCkCO9SgfNn
ov3//bvs5+P+V33WkGwAu/jaqin7MkQaJMXXOk1Fpuhwbm95pgHOFRY+/30DNtfj
zKUqnKOLEF4KuyMggJW4egQX/F4quTNVyQ11no0E8WAWCE7OB6moMXFpZvxe1zV6
Dewas4BobzrZk8eIdKy4P6RNoUOg0kQfUwjfgeylPFXfxrMIEOKxbeIwwkm6HWBe
4rTb3AwIJ0daKy9OjiO9pncmeME5A1t+osJrlQeXeWJqdMxjtt4sHEmQd4Bv30uZ
fBsNYME2f3bmHD4Eb9w1/FFdcAR4Q6IrUCEtnq+VNHxUiYH2PMJNwqF/32CrOexz
bNxC428r153DxqOiB76hBl1WBet+a7PBtyKiHkawSQhhlYDbg2ozi6STZJ8OaFBz
9LQe3O5Fj8o2FdSGAEPdEoEMy7k3v+IMY4O2d+M5J3r4ztiFwTVHhvVDp0SFJlj9
vmRU8eHq5Djv2YN3iGd8NGBIyUb+jHNghtW5G/JK+QHT/XrPypk88zzKEVNjocv0
ogecyUP3cBh2P85Zx7NIt5ktythCaOJCykM1Y6QucbKNcL/nO0PPjAG/ondqpc0Y
bUjaT7ogiInJEEdiyS9dukxNg7E3H/1mEkFaIpiWSRfDel7tFMZhHWIXNl3+DFqH
mSx3Hfvc54C8mEvpqfHqDguHz5DoBoGv/3MW/0bfvKGN630kT2uGHVw10Z9DjZzL
eiNOamUHCXF628b01FnyGTRxQmFalwaF7t6GJ9ihhfoyMhviZfF1oQkL4jx7VXvz
1gVLD9Ouz0iG8FBYO268J+xRW1j2qOOIdYLBoEkM5KLdNjI2mlDsdSyhk55eEydB
gsg3i3Q/EA3B3Q26mur7EvB80wIxpLXh6zfmGVNFb8T/ggTQ6tBuE/5I1I12LuEv
jLzXIUHb4/rRRbZF9Py1Ql7hhlewsAU557lAN2YrXaKPgVVLQF6RwhQD+zlEmxjm
rUtLx5I9Ej4u7k8TGrNB/rTIG9x4rvWR++D/9UofX2b2t952DycWf0J/wxn2cRCU
B61hG03Zg46IhqSHk7FfnO1dOwUp8Wq1WPmGFbfjfBrmb9vpZB3+eo17dEgR2VLf
DwXlE//fFWFF3rDoQGPLrGIbzgtP5XTZS/RrKhGjD0UgZBv9ChTzw7YRIxD26LtE
xTvo/PqxSs19Q1ByYP0JXP8gy0OqK9N3ZyN7qMoEiOwx1Z2CO7VRbXX0UzQqI5GR
EihQmzGFX0J8TwLZXxXaX2o0wJ4mTP2EZ7P/v/UV/uL0gYsAYeQI93shqbcAql5e
raFMTue7mjREuMAzlybL9kFFBu9ROzmAQBzWNB1rs2nCCBW5+X58c9VzK4A5kLg5
C47WS0N3lXXeDJ6JAFsMFc0cOETR3MHIiM98QVmyf3EDADlng12vMbEenlfKvzfk
TuzzKjczLSK79Ox53U9oU0lMO5P9u1tICRXpna6iPuH06AvDTWct+Hg0GtsrWcTo
k0PRMtPQJOjWNy1HMPGOYsDzDuPZgKDARZLXKIzj7Ond2FvFuztDhVjyX/42PQ17
4lyKow4DN3PbOhCYAV8WfUI+Mpl6PihI/cb4yENNeJFmdqaX4zYVe598zGtb6b3a
2QfxRIS8WnDkjUNpEuatno08lvN3sMRdisGpjpyXXv/deD4Grdg/yvnufVzl2ltV
fcjyKexT8zUTN2eyDkuKfv/RcPxcWfW93/1bDJz8w1mRBi7pfqJo9wrsoLUwdDhn
1TUJqhBwlGrvkKZIANeOlFq5w1j3EZX4A97KJdX6iZV0rqhb1TZ8z8RWDf7fsGVF
/Nl0AR3LOa3k/YAXLNlFKUYYN3AoEB6CysRrlfUUB90E9V+9yDhvzoRQc/Sk+0Lm
XxjjzA+YA2qeIx388MubpXrImLlV03OW6I93IhtMlgFjHMYw0t1NMVOvmToNj0ud
KgtF8+V9nHzh29MtuvHXaSYZuvYw/FmRVBIXK6M6l42x0dnKJCPHNNRKQI3YFawp
38kjDF1ogA+rrOC8NLnDZpiNZ77kRubztMjC28FBxmFZoNmIZogrT2JW/0heEBjr
ApCI3mp5z8xqQ/5uezwKM6O0W2IWUIkLXLHSTFx33vQn7eUTleV96rV8S2dfz03v
N8F9GB0Rlcuxy8KMY6XFGCD3HuZgShcpdvfmu4LUskfVEI8FxXdcFxCzUGGNQlHR
NKSqfTnRNuvlmgH2jDL7F5JK0+M1C7jdKQrY04I9dbNifzKpM2EZsXEZSS/BG4f8
9khBhRRNzMpQL8ocGZ3rO5GJRqyZxGsc00tARtTORfI4lNmszfWSh6ED3nHrH5+I
bv9rYPhjZ3P+2hkE5ofPvU+cAxV9V48RYBA3OfRph1VCVfj4i6fWkMegeCEGkjsk
0pWFUTmU1wpTZaFsrvBFBgA7jILd0qD6jN7UC5eTMqa7IlPomHH0vbabAoloYOCC
AEttYJIy30a4v1qBCvkrYHyMMf+oo7JG+rkgg6RJTqjbaKhZzv1RL+kf/5TY9bsV
4Y97+RYM8crSlvRLJSTgElR5ATUigZjmw+bA8KOOwOGDCj2zeMQdYgreBgfC5j34
/cowxgnDvEL94uO4dAUn5QBgJq4uCiDrPx/4AAtGpvzQt9rE/LV7UkmapGE04XP4
uJOL2k2uA4GiAeVHGxbnxLCAvGuDyIkUs85V8OypIuGqy1A9yOpkO+RZIwMTIcJQ
dpI3tm9WB4YIrIU8PXqJGmjVtXgTLlEu7KPwmXiDw0Rmi/MdP9kDsVl20Shk5r17
GnQ9pP7QS79H1NvmhxhJIufKaJLumfL76btxrTHLl9YsoJaZptAYHSb2F7g+L8vl
pBmO4Jf+46QfcDMMhH70xa/Hinlhivvm8hOlPksMAnBgDq1L9pbTt5nk1QkHq7Mo
+/56uVf+LQeKq0pzb7NacPm9EwVseePx2iBlb0uE+Kd31sxlcy3HmQ/oMQYJ/JrP
OZFvkHtTfy8A4qQ8ciZQxYVWScyVGlb/GxqTROEkEbyp+Bb1FiLQ2PNY/EhzJ57+
8gbCEpokMruTxsWWT7s0Wgyc8HSNmZgBcWLynC6/sPw6jKAsTr9+CFW6AJMLo4xh
gQKyiG09TsTtC4I5GP34ybwnksNSM62dofxfCeMkJDB8Rhh/IdFu537Q/kWfoCKZ
BhTLzqQmBadLICD4BsF6fIDVHWkRyEZSnovxOz1B01RTHoDz5ERCpyRM9IoeUtI9
i/bN1Up79iiCGRyubNKPoDV1oSXlMcGV+HGXe9S74ya+OeaRcreVDdyOvUVqkJb+
mQe7yugki9Xkgdiaw93+ln82kBEGc79bSv5/WHFXWSWOPejn6QxSdQ+j/Obwees4
tpmnlOysviRZzIp5+B6dyd5wND9tstKXT+7m88/lNMJXOlI4VtGl2VyrdbEL8nbX
NxCHFobxS+GRH6yC6K6OIdFVY8wA+9rZOoslLZbHVNK+Nr0ytpea4sP155TFH1TZ
wPH+aGgHrAuwfYq/+s8ZG/w/eO3FssMk+USz8UcO94orPmxOnwvLBYgmPJveuybk
47U3DEUQgh+E9tTgTQBB1UJJCUneL9Tt1TX+i++Q1NXI1zaBIz+I9r4XXEh6/YVW
wjIuqMVmbaa2QK2w+phHGwOhirHXojtE3OC6ZyScuGqhQdi0htF9+9rinJgWZ0/0
Uwt4RvyOEk3OQMXnee8kdeOGL1WV3X6nu2Uw82v2/eugaBC51y/5S220CozpsM5r
1NCmTbIuSKP055oBFB7E/HdfHErjsDnuB9kHa/2JWaJxsGAW5c7WB+ZFjwdYyKy+
7MSLx7G+YyH75rdJeERG2KHYyIS5/64A5GeCxLPop8T8d1sBOdp4em3/XnxSGl82
76+bJ8wmO6Q2CZ45gpA8GwJm2YvV6blMl9i9seahTLh7YJ5c1Nfx8wo7GdfkMXAj
z4fT5299WZ3FCe8IdQEXqck907t38JSyxpjIlZplw7PHcumXLVaYIHzkqTGtdqKW
W67FJyN0Pg3w5F3yl0IslDSyxbWYv81nGQ14lxzFQuRMyITUXSmerXReYHIBS8nk
CW1CJj1iID6YDt6v2HANtR0nmbm5Mf9ePbm11MMvqimpt7KxXgGkPsc3buEjeDr6
TjnVkYxrR/5ZSLMx7OQRDOSiimN8FM57kSbghjvfPvyd23W4TCnLcxuxAdI0Ij/m
8XRcMKPl46CanDRYLqFyHctR5hkqjU9aKoFM0EcKmpbMxUXRFv7RS7PVEd9GZSbw
Hn0XALP5ZfEymZGcXhvbrJFZU+UA8VfuAy1z6lCYIX5FNaaB/NCQ+fxIBRukzBfv
ZxFhbtojvUsMtXpsqQ9Jw1X0ksxOYBIEQnrhFlMzO7iEuyESz3Yysm8wnN71jRe9
CbV8xe1Vzq7hHvMesXGaJvtWsHqhG+QCVA9wov7KspxtiOu/PoFplI0jVQjZhq5l
tDrWDJoJpZWWiNfYjOu9a3qHwz3t/WCwUjAcnHR077PWHHB6cq1qIqZPV4HHF6WM
evFVqK2zm4Balvj2u1ikDwC5PpHFoSBY36BDPmx7AjyDqnSXqvpFdfPz4LRmEqkh
VtXgXueL8VlxPb1frt8+VNzMwDTq5UVjbtrN36nVBxofj2E9ktqNB1vD4Un4yHZW
F0lcCMJyBTDo/O68mwm+mVULwE6s+jsrB3lEpNJuRLk9eS4/cBRhxP21scNWv8OH
GqUbsFIsdN0ZJvDvriEPV5bAcmHIU9zEAeUSIj6XGylpCpoKjMnG5y4wEeMgaIUY
nBjeMcbnhnWmqko1/Ua/bSeMLQDQfyhNI8rpTXpGT5DoTD4MeF8ekApWXONB2GAj
kwNWxfC9KjuNiBgnl11Uj7JWuo4hjCQMDoVMMNA2pbXbv9zcjBX22b5oXDRw6vzP
QcqXwACb4CtclpR2iAdzk9r9IiGjPHudoRo0Jiyvfv06MXSS2NyJiiaGh7DOO3NQ
riOCeVHKR3L94RsE9A3mBVn++5vn+xTbmKnNhpKi5tmRif+N0HV8HOhNoxlh+vP9
f8b1u2eoevIvCNtPpUaPep3lFPNQmWhDZoLJnrEX1g26r3o4ZG1B32zQOpgUjoAp
oBO3+fuwxtdcueoEmX88ULH6ibOOusEIXf5Ys+H8JQGj0skfe80f9tj084XRHLFo
+xit9PBGx58hyVPHdenPnxbSFyh5I5npzp2eqpde18265SWGsu1p+NzE3B3Nf66c
TQcFv58rUxIVC2bMeXqHC0UL3O5KBJiGwKy7iDhSSRe22cwgsFdcZPFyq19syKsk
f8TahakKaeSeivAZr2K7p0Y8siBNOTbqQJRmbmOto3p55i1vklGA+/pwePps4Axw
b7pnNlGVBZYrozMsXJmre+PljUFSox2TslthpE2+hwrifDgT/8Fh5Sma8+q8Ca+4
ppgvN1Vli7759xlxJLWh35xLTl1YnCtvesBFOZENBvbmqtHlMeOzhDL2t39jiwqz
4pPRvOcSe2A7UFyv3Lmkt7W71hKyjpnsynLNARTSoXfNnynwxdmkPs1JymC/CrSZ
vEaTSn9GenBaydRrwPFCAhwRNDCyEAczLQ5kFqEqHWzmBN2n7fj+K/lmuiH26/uS
+47Ymd21A0qy1P+1HJQ4PdbQNGUaYGZius+zluDLYEZiSRCjIuZWBx6XYaxMMFkm
b8AecAJWGL4pjsMWaOsZSX8+2GlH4v/cKsDcywS2fB7dwOSPq3Z6JvfG6AFS9muC
U6OQ63MgpI/JYiSww/Jk4vtraGYXibjplN3OwaqOHjnAZc5cPUs69QBBP29+s30v
/Ho9CENZwkqFT8ajwBkeDe5iKtJTrbUo/eYef1zLQC5fvMBXaInYIASgrtFpiR0C
n+6RDNnl0mewQVAJ60W8J9K6x65WouEhq3dkl8Rg0r8DSTRmr9DeONp5podf59Nu
J1Niqp1PgX3pOSxWLTu0nryT4keWX4XjuUnBWGgIca70/AOnqgwVk1G59hBDkDQz
tlzAeJnNJz4da2zIqAlcW1FaIpaGoNWUN6g0d8iaHq+znwYJ5pILiT4RfCee4Dmf
kLKEJDZTHd8t5D2ypc+9fLFUywukCdiciXoJJrRgO9sMVh/SAlWA7Ne0EJZWq847
meEpZeFqwKVYUY6l4U6CL7O0gayZ93B22rBNyvwcPboT5eGvC6tifumlTHNG0z4j
v9VzCa6lSzJym179hHY5hjq4SWbAZmWFjKlUerHbvhSeMIGfMYIPpeK2G74KVSXH
ZuViAaJfSWnwhIc9WZroKWbxb8RmiIveI0Ir8tkF72Xm+goxGiS+VLB4850l5ocW
0xPXI2Jzaf5Gc7ZUWA4peCprEXBnLJva1il0k4+eYTDbRxBzz+3lSugWCXgJKrVY
TQn/dkPhMkOoEQOAeOSG+ioX6va1IHlTUoS1ashLjfNlIRdZ/wTX7ooOorWLBr8y
FDMv+ahH4MPLQ0+SAGUnDjXCUi3dde9sUJ5ylaP8Y69RnwZOvivg88jNLLQYca9I
F/I4B6TwKDgyAwrVF8qrnERZpBTNN46PAOuGWl+V9/HvbyztXBOoPJeTQJ8SrYwt
KzZuZjhFpJFkOgbhUiLLVgWy1w+IFrGS0RH8cCKih+s4tPoPkFKQqLLuqN+wpj2W
1yFaiRJD9ejb+QUL0W2ZEkQhW90mTJ0xnNTob7OhmGurge/dUUpEACVEnlkFkdss
IaxSSjDNA1iTj3daWSS3kV8j0Xa1DMNPton2VR6bRroasKos1p+97HRVVm5MzjFP
Ie3amU1KcSB7/s50xlzrfZq3SPnamlilwHBLLoRbi1/cwBTfrrCCvHZFQacptpQM
TKiYT8Q35Vz/7pzat/zfr1Kh++KfEdFu7u/RnpqSKPSLd8VnjWc4lPx9V0m+plCY
GxcUdPBB4XU22Ame9cty5QXuoDQtSCGcDG5NSSt/WEmyqC5kJvxA1i5VDj9ONA6B
Y9WrUj9+UoGxG2Xxj8c4Wxn4WnNlF620hY3OExlk2a8seyPt5oppAsD/vt4l+l4Z
yggUxF4jLsZok9iDqH6KZqDB/Xx+LPdu0Ewx6K+rwjIpZjyw6/g1B8AM08yH5LLM
lwb4+clCXbCTq2AFv0A4c+GJ5b1lb1joJbMW/+lig1hAjmBt1AUO8FSZgo5K3ONq
JQ96a0+4Fw42AYaSSsWuWIk1+13SK4XFBzkoaDSeC75DAiFG/Fg1PrnD0t0Lhg40
h375u1fsJT2h9vHPu+cx1rQSKmq8+Z5AsJYULSCaU5IoWWBOqSMBSxPYyAhLReHw
vxAAwvfi4uY7x5MjxEoFW+E6lJI7INKsh8CFZPVwFDbbFG2N+wiceCgb9Y9Y6qsA
TtitdL24MW0tWsyM58VHH1NKifyVHsO6UA2MQuT3/hEpIa/A5i75RNGkHfIPHw4v
A87grLUCpzgceuyVKuBDuXD+u29PMWvF/m996ZDkASLF2LnQ7wYYljQLZavk5c5S
VFOu84mo9H7x1JOHsbAZ0a5pVh1owVQwVkwdjPSwolOG7YggMfiQu1yVVZl2TFRb
YULmsx29VdqwzluXH49L5ylaEZ/V1076SjGeQLSo+VP1tnpLFS6OUWgC/YeGIfeu
3X8FBHyRPP4lmtUj3wnnItpMgXpuos49LwG0VL5Bg6Ts9t7z89saMhHQpj4e/yHD
1uTrSZ7pTTQKs3ZhJBdjLottVElyIku2xs5DvgBg5TDl1CbXSjfp4V78TO7Syzp6
yXDA7/X1mFCY3qq4EWG8W+xf7gUhpy9aKHGls/n8w53GY/KciZ/EmAg14mK2dAr1
zyz2IFc/7Q/cO5/AdRsHzA/I4ukMdq+guip31+xAvyUjl4nBQz3V7K1/1+IfZcOO
4KJtlA+aR41sZZMEj3o2afg+b3mZeTTFTRp+wpqQDBFgDKAR2k+Mz27skk5wUq4K
BPg0/431gecTaifCpwg/5Me9JrMyVJ/yKw3thTe47NHvUbEgWUiYtUHFY+s4wALC
9x8p2ZGml9+a/MDbxv10BrFEDrV8Qjr1vgNyAyxtZSfJ21EyKucaLU4nq4FWlBBK
TUtCDqpL+Q+Id8iYpyy/I+3xOGpPwESO4kcOKtO+0V8ESBZYetrCnF7J4dTEr5OC
w1/Nw9xNwsEfqSMweBO1QAJcNIau8HPeugpsXGYN0oa+5TU8hEIsHmvRi4ZT+owq
aEyBH9tYyOb8YL9a1sPKJ4UAhKgJTaFlP60wT8D2lfgd38U2UfLmx7rv5RU7p4aJ
trb8Av8OBPz1poM/1+GphKPfFKiIZDUMy7VvFPfcxjm6N+MYFkBE6gYCrDb+zd6e
Nd3KAaIo8VRI7sst9FGoGsqaz/0g6xVQeaZBr1IxKBgcnD5enWOfng98xb0L9pz3
YI+vwdIU/zgkmrChtj9HGZEdFxQ1eJDMOO+yLVSDq3y/8VaTri3f56j+tE4k5M8m
xwlG9oPNS4FeZfa2lkaPZ9xhoJ/ZZwcYdBlO6gZfZwDeoRMqO62f8bDhxxsm7HE8
MdQKm8CHc1oQ316LBdszIewE6+E6nKblZS2cJjNEraRPo5MSztJLVnZ2VONqUGtp
aXd076D/H7RkIzblQZZ6kNawfK5pkyKFs2SWJ9dA/KOATfe8/eF00XzFc4bQf9xg
c007LpStWLhwkQvyI/dosJmNdeWzpcs6JTACOQ3fQJuPZgQdgSKqJGO9aQcYCSmQ
4O91vhHjsEXq0f4BVp5vZW73Yj2mI4mhCGKCUCDZ57LTb09P1619kKBbKgPRSLk1
rtvZqsoKlYY0HZpDl+osYu/e+39CbhB285LkQONUXn5qmSqvpJRYiegVCmTY3lY/
DAfM/VhqXvmP21qmeADA+4B4RBmcWFzDMRMQ4fKwoam/CbB4B3x1vSkDoX0kVTgw
H0sWFghcRByOVFp3Wm3iw3311pBJ6dqyFlAsYBV8XzA2ufd2Tzr+IlrRwpeNBWxH
zX8VuQdaTSW72yDhpUMuQ0yxeszdM4Z229F+viVby98nqqGR34oRVQ25Ku3rSl1V
6bXYM4batUz4ltrKIxZy1XQLM39+r+DUKiG+LjMbY3dxwZMZKbAAXTTx9WHQ3fTM
R6kRt0bkJNEKR5VSl8VtGI5JRyrBoer4hw464FINkiQH1dC65ZbBGqT6TXvmlTg9
p1SnzLhL3tFbC/vbBLcQS0TzOqPG+F4+xLfVMVJgr1DYSacGhBgwXu3NVmCjSPvc
3FKBuE2GzIszxVy9IuHwAOYFWF3xLgYJWOUHp/4pnU9pFpMtZhuAAOxRqjMCYE4T
3m+qS50kOVYnvAVVeBAo0JagPEusHAgtChSVdkwWgqpMkr+qEcFwtzlf53oVcuc9
PfSwq/VfewiOUmFJGIVkvVIycqgaia+Ugv6dZb54NH+STxG6Xru80slhAOfcf5tR
BZBGDffp182goV27uPdE/CSgk4NsWC9PyuEZTqGhcU85kwo8s5TvVKgxk8JfSlr5
XdH5zTxw0/lYU9wZR5NdeCfgs739NkkQ/FQ7GwV2F0hwMOknezytWzpa5IGMgXRI
Qs/XVbDU7jHxUA07grs1f+/6gVT/1qog4ZNAO1EhQMI8KRxB3zfOXGjq7HzMS9JU
yRo9l4UbLb0PjgK3EJspRGAmMEbUNfbUE0F+szaTl1K3a7F665nB9rqUN4jtmzAo
nH9SKWzOjuMpxJuxkDTuwc7ao9/fHe+MuX9H7ITEfr5GNRa0ja8o6ftEDtiP5A8w
qUOmMFJNVYtubracLCbh+AkJkB5y+buHC94BE/XFcoIytLzjtRNSPdvCWjRHF/3h
B4r8TXzJQiPdzyJEUUjq0ERhkFFKnhPfR5+4IYIbSicf+fIT41sjRtC4cVI0R+e6
Jp6QGPlVHfVnTwRZEQxTj+LDVIe6DXRCOtMSX2XcrvRe3Yr2SH3BccygCoboamKr
NjJzTsJlkSYpEqAyoaqD3efupeQHP6Zg0xPwhoIqvCP0xBbBf33ASMUmKlHiknCl
9n8AMfPPP9RNI8coF+71xfnk80G0UuVWn03qRcFURrjqtuBRS1xT9TosoDq6KGwf
X7oTmPtL/tltA7iA/Ij+Y8FVUwrbmBINZEu+pA8QvhqXflupSbMpwWy6gIy6RkSp
uGMp059uXWPkA7Z/C/jwbwlruT4Eh71FTJQ2R06eTJaR1oXVleR2WJLIyT0aYxwI
qmAG0a2QsJlPPtWljVqaSHbN/i0ZuoX3XLMtKLlfnjPKURWRNAyU1/mP0dvBdAwP
4XFgsp/So0dzFGm3MwYfNoXMGJ/uqtYV/N8i0u1/B++NxmxV4mQKs2Wvwt6xkV/F
htERvrlp6NtuZcGKWFPsQLy3dAcVOIqjsmFNKK0LL0Yp3SitxduVHUortAwTWMlm
jxtarbgWArgxAxbucCmB6kVxXTyeNwknh6pCsvFxxR9GCAlamWQONTE0Li2bPfpm
LnBlwB/mgd8OTkf/dKd1fYWu9O8eI+/4yenwlHBXitt8fd2BbD26Sv2/zdLk+SNG
lX7jm4eFscapeqin8rtUKbTVPH7OhhnIrEkgye6T/kA0P3sfiUcaZ1G2Cc0gJV5r
P1cgrLM8tLtNTAWSzh9fHEh39BanIO/ylgtzhL8NZyCPq2L/UGcV2FrbYOP6foCr
GMyF0cnmuzC9nQ/jykbWUJ1uTW3CL84wXsQzXHOP0eBWQS6mmxRZrx6lAxlryEwE
zYbl9u4rZdrm+uf4Ctti/fAIE5iy8AUdwne2xQjuaK8L47JRlcVsWLZq6PqHO4m4
hj+utXgbUbHEAeYPi/ysCvo/nL9UE7U2zobgcGDeKwSfAGzD9gorNBvpRqRkg4zW
AUVjyNQtbRgVdVGCt+aIqN8clnxoHzVXX+cfcSFVmeCFrOYYTnqgqIR8XJGhH2Cf
6L3fX++XDiESfSSINhW7YrIG2VJW/3enSthgBS0kQbLndfhjB/2kLBwIfVtdBkbL
0KU/u6ACJmGvZTaLH79DndE1O9Jf1zeqRgtjH1WUfrS51KCOdVtlx8TF47UAP0gM
0okqadFM98P77c84GUA7jgD2YVzhVHzO0PBeFuMi5JK3FWRIn8QIqMTNBAL3mt+x
3K9DefHAYnlApWqOmc0xhdxHB+PJNoWD3pdYPejSfulR0dk9AsTbF3bv3ch2KtDY
8CJ/AX79PKCDpheIHSGXVdLyd05AZ/QoVESIc/v8iyiTVcXf3C55frHIucH0B70t
oK1QPdCY5uXRDpYtyKzSHS1RNO5J+HNpTPz3XPxCdVuq6WwePMeIeXkCTzJEU6aQ
lQrFiQ9gJt6h6VT/F6RpX+u6/hSN8+L/CoN9fxskMEoBpLszQGa7aIXfZpX8vSZ2
zT+4b7CPr9HPm4MIznIBpZeKRJp3OqX9VMlftzIxFTKrSf2zS0VmDW9U1Hk2QL2y
3sgzSNh3X9ILAETvXrDrzLi+GlyOsDoESj8we+G17HslYsKe+dfrnwy/xGEvnnAZ
cHqJIeRBxHPGQ3KqTZe9Nf/qbnBTr/ijaNjFtMWKICDgYm/VhZ9+uJlToHuCCgLt
/bAMYa3EnVw9JVPEkNRbhRltepbgB7Q/p5BbsmO2azV8mwcMC05Q1wDjF41ssZ/E
vKu0AEZnvDbAZXhGXTtAHlnc+Nplhg7AKs1rUr2xGymZd8dlU94+NgPr7DWIkWn4
qn02aubAbfOldfNbdPGUqHhBUOFKZQTDgz0eVGrfVkPfPtCO7SgtpagvyXuH8ZXo
pxnJYvsZRX1sBjbRHEBgqPbwYy4ZP+eaYzFbLV9Hq3CWBhY2+VjnuzVaLVBttxlP
pOQPFufxHwzqM6s71D2Ntd+hT68wMVF107uIq37TAy+Jp0+7GrFTNdjNZCrdIBe+
2Rl1PXiQ5FuZ/5U9Lqr7k7090R6ZjVpG+gMc45uIKVEfNuMEPBKJCY4aZ6ZupP6g
3qCklCgAIHGajR0B+17Ma4EO8Bfr6P6QGh5JPXkcw8YCByva5SxwTiq/vLFQ0Irq
MEQOD9B115VbiFMdaZv9hStrRmWXzSKBCZb2+9dXFW687jx0vXlM5H3YZPNmcGuO
D7vgr4mj58a3jfdiMA/YiqHtpbywBrFlpNEfeliHaDTJkcLnB0/skZIgspQLXHHe
I2KMU4NHdnSlRP81VuxWqnNdGFuIpgxAK7cI/ArNCzVE+r9oEaPBquMW6sJdpaZr
mr2vBgElN6p0NP2B2tJJjXdlz7EGZ5W+9unRfAD/FCPCOOGeKXh/ZIhQzqEyu8dR
ddB0VNZXN1cH3SFhMR7DCzbbXrjrle1smPqDzRP3pTcxSn1YXEe/Ks0F92mXHT8T
EF2JmMOeCgOVxnVsLSScu29XCBxFjn073AEKwmfdRz/Engur+HRWxoeIIj40anPQ
UAbiJk0ahZ7dWG2kmilAgV57TmxILZ7NgKCBfQ0AmNWfDs0Slp6LW1TeGT9NQI6y
1jsweT05tbJV1ZjBBlQ9oA/mnH5bVa9D0XrE8/bItj6HtRRA+dFfpE895tLxHihF
BCa6gvifUK4HRux4debicLQkFN00xtRDTEruNUvLbTOEFmXrkDnxgJEQFblzq7Xt
fJKMISVWsAHlWFXWCCN2w/6qJDcuK3k/xOeXQq+9VwMj6JECWatW+bdhePeUdDsg
gJ9maCNEb9S76YhnpLzTqqOhajFqDb/XvWZ+MHWQ5ex3eB23CM/G86927flpTDuH
MrewNjTmX4xosl3QOEdS7RD+3DENMZg3anmfgSX28hdcjXyI3pMgDiWIaue42SYA
dp9f9P9iw3cvAF4dQcUgt9axJwb4ZbgXK7JNF8803RXg1GoodISK8lCVouWrxVFq
vbbD5N/AHmp+7aPTf9a1aszet0S4y1jAFNvm8DXtp3cUIjzML+UvvbfBY6Fa9o24
e6kuU3iBKCoIRSlTzmpUlW6iV62uZMkieREC39SOaWB9dGfi9paSyxhn2Qq+1a2v
IZcG96RnIJ3Ku4IG4wmJtCDvGWo3uT6cEQzdnIQ1cKktzYEmQdiFge6yvZSdw6bM
yxuLhUyzvOSnF9CTrHHkutGwHYUc8FHk1/x4HSW7cVAbBASAEcjdSXIB4wZV+G+D
3nVD/tAzGWCqnxf6XH9/infkJjZ32ry8y2oa2iHrq7CQLWFrXvZ9Rz9Y/Cfq7tw+
PYzL9uFWpKp9spLrZ3spvTWOq+Gw43deRXQdfbguQ5t/aTLeYL/yrj2dgDd4ov7g
IiksDwgsA+K7+wUqrovgG46nANBcB3eY+sGCbK3FJL0eTizN8IYl3+XOaeC9HmZE
0d6zb905KEIRJefaaqNsrEiH8XSCnAWqRvtPgLos+GOgabHQAR0nVa11ORU/Tv0X
Dakgxem0f8PkQ042QTpcD9AXDTFe22p0blwUPJ0DCP/AVJcoMcyRrbnePpY8FS3D
oiI4/Oj8/hh6oAiU+znVyPEdpIljIPbjGPceLt7e+RHnGYipCBlaz/AKrZ1XKoHS
qdhkq7E6O3EeSlgC8AGRb2psYLciDrJJFKHPoc7cqyNHk9cHKBIbM7FUfqDd0FZV
WHidNnLeqhpBP3cSMSNCvp1bte/DgSJCpuUCi8tB3T2MTlhC6bYXnSPWov74ow5j
CfZLdhvSEKJkAeAV41NBNX0liIXw7hoidKSNs5CKPjx4RWjvmGbvjlPh2l+6wJ0R
cIVEGF/O6cQdTmPtbUmerYRHR30SFNwYVV+LvpuoPBrX/YiB63oXjgHCDK5sJfuG
rByC/f9JW8YV3Ie271l8+mISR13AfO7sDc+i7SrNto2fNop9lP/3EcebVJiRJBnp
7wNcnCna6FUGF+CF7S4I4QTIKE7yVGTkdBUzLvpYCQfVbiDCocOxZW5EL9j/m8sP
r2OzYq87sqXaMNL3e6tmMrPqrsPO+d0QwuVE/1X9jLiwgpmRSQvs+nAX/IsCTVH0
wiziPsezI8+qQWAO+RJ2IEynQB9oaT4VFiaRRxl2ErY7utqjxXm0qjBn0TXpjuFc
68ATMnJwU/m30xC49HP0dB5xDMh7d+POM8Z0fsWiXgmBx7X3s5JV4L0fNoKe3YDz
4lFeSczAa31DOPvzbEymOOFgzNmKioTbkPag8iDg+2MeAI7nx+mKm/dBQKtuLOc2
YEP0/qXBO/lb5om/azV5SZE4iPcrDTsm+U0pOVROhIejC/40PfSw+XX2GgPQ7MDs
kEsp8QnEYlPWcO4W59afI/kPKN2NjGkCLxUCqMwZlwIylTY0Ht/dluTP7X/EWtzV
FwO/tGDk7Bf/ik3S7M0Eb3vp0Cqlcqn2IgzVMWJcb9H0sPSx9Gx3zjeZqgnABIlS
Jjh9s/fuiGCg5PtRLPopD7Bp+TO0HkyPgTPYevnUGmvzhuI3MkHtqyOknBVZ//Zo
GEiIPsza4rFb2czp1cAaMrndpZUUs0OPvpCc+U4vbt2IPw5/NNo48KUxwIcWgSK4
WBxgA7sYvhODY5vtWWL0u1uGQj8om2n+91pWDCtIPGJ7KW4RYKsLmdPc40kMVtub
o6eb/EgQTRHhPjSizRIR4oytm2GL2KPQFmG6vwRYqI4mJSSYmcHNJwTtpevkvK38
IbzLx6m9ASN0/ZPXN5zlVzacSBdY6cW3+VlivmJJLCK7gXS0MDtZ4um3ikUmEOR4
jLYlj7BrjiNgwyNgKGdlt6iLT4EmpEjLLacS5h9e3Vk6qWfJBg0Sm3YPG6MKJtFL
nB18ZREFjDN79757mhIUTg9vP9SjlrGJJw+ULy1PKDngADlalIOiC1Uq0zHO1IU9
JhKzI5mXMkzKQfUZZN2F7T3qoKMF1dsStoUgEezPVjW0+Z5OOMvFS7bNo3sFQNYj
m94DGKfeC8KUcbn9A5cOPijwOfVcQxNaZuMLLLug98KmNI60hrPW4xzWrrD0nb6v
I2w+ffQN41xd9Z7tcDSz8gOZGakklyqcoCKghGqf+2U145648D58WQTOF4YaRkSn
0itKpmh15xDoQnYvMEfMesDAFmPayM0ncze2wDkgrz/z2LW6B67T1PjXcHP27obR
MgtrcBIjwLnMGqhSy5u1cTPvtOhwnPjgrKVRK5LSx2WRlKa1mg484nEkHUqyDzMx
Wf4Yfqd09BeMUILd/EbC0zLntUBGycp9KEfLtgrnSWCp61eX1cTw8II2oSxCl04N
8dTAzbfGqwECDHudOgckLN6+swxXbVUesi7ae+iTH49GUrG0YBNdZGHxxG+Ygt0J
Bt1u3lI8pafFUzMAayDxDh785mRMWbiycmccyqy3P5/3vVHCeKcmRcVsauhwlaQW
eGlZrWtbIsQAp5RUV8XfXECJuwbiqYI8KDAF9SSB2Ys/l3DVopTbOa1db7OYSQ3u
jMewRH3GwxJIzdUnlmCkRAlu6IDi5/3HOJampKYP7aYHzQp1czsWqv7tuR7oPQYh
I1aA5IB2LC92yLkOj0JpniMfuL+lWMNFXTkuvVYZVB/jI1xgFFbr84+rOL0d+pw4
SwWvnQi7sg4qcUgWkPWqYKKLGT+KnsyTIZJUxV9lUydkM2VcWyI/MShTI92YZH2t
4Wcvw+MObJtZjl7G+Ca3WFyEtB1LTHk6f1I1r2E1aWXj+kJ9QECjaz0UJD5DNrd1
P3HyB5sg2KU4clcw6wV4Nm6kIhWDxvV5VZMdciGRzsAhb6CLlGz5/X+LdGp+zZYu
NYYKYaueZv9ANH32JA5gaNyMS/Ho5nf9liITK1GCBwt6x2/uk0zkqjVXlDxpV4B3
gFnTpagXHZ7+yNhZvm8efxgL23iK1dja2IsTYnW6oltu3MKlkCoMOqcJy/XW3bVO
Zw8AziVOspwAvKPccTt2huy9RmG8+fu6kNmEWfrhzufhHlKEtfrK0mQjMnj/lQ59
pF3ehuOIqACkmiUgtBJffJ+v9RZXjW9oKTsyixJseDCOXV/p0UrlhLZ6lv3VZSAp
BCtI6pwUwlpWEmM1qi0CRHDwUB8RjSDfahjH1qtrgbhxXrztbaZ4px9VTjoItDbC
HrpJpX4BdhD+b7LqaKX6GKVFUgAU2hzzLbLsx70XRI+Cw6C0GI1AdExd/B2Xy4xX
25y+NjEy7A7OhnYXzFXXYYTA8RC7/KimtVhglOjr6QernT73zTONr8beSPK15adD
odQKpBZKjF0I6qFZ4xWtapYlIlDvJq++8jYzqpX23rdwG2RmVooyuW+YC20lOyNy
oTyUujgV3XupPB3me2B4i9OpAM2k/CC032UFp9niSGBhjfeq21av9fAbQgVKCfA6
HqRDpRST4WGmKNKHHYWCNTXRAaP5ArQeWwsVogcSfn7YBChpjDIzCeUNFHYbSa0h
QNAKIiD3SsJgbW1QhLcXDY77YyA+dLo1QzcFIe4C8S33CQ9dcmsI2SbgCffDvwqn
t4jiXecZAp8HCgI94/+A9t/ORkuJmgwN9fbshetwe/utfaWtZYBSvP1+b25wEbk5
wEzUe6SMjrDGJRam3ogSKBu8+eZfxH+61yuerF1pBWQSh9JZgpUXIDbVPsTwAiMO
KJCJma1+4qyRvEfI0YSspljStHQ0x6UfZgQXvsPZwXwISQfKCwxOVObFDI6fzVTB
FMkcauU962bUCy6ThxZHmAY8GRF2GkASEt3zntDYB7lFretdBwkr2cKQmMNEkFLF
NxeBOvjYLvbd2s+4W6hB3NB1DGpB43ju/m+Nroz+nCICW40huOmjpa9WxiwPysJN
x4eEmz0nMuAaLXNssAn/FXfz6sPsrzi79ThTK5YuG/ft2F6vKqcHss7xA30mT+OV
DjUWygTlLhSXZiMQlFfu8NFkGOg6rqXI8uzUrWAv618mB75oQVVNDZnJQ2mNp89L
IzfWswEn7SMq2+4X9Xp9MQCCKMv0FkoXeBqkwb0ZBDU966cxslFVJg8+N9hFduJi
nHhupuxhbP2qvSX7nbJdDMw7YtADj9IbsTVylWm+H//2gfhZVohDeFjcYOezDCrM
R8UsYu0OpY6SEDkniDkp0H0n6+ZD3Sfo3QGB66WiFBwiaFaIJq9DrSVVpeibaZ4k
KzQARJrAQoKltT84u9tmlOhViAPeZCn1OZQrnv0ebaNbZ9jpYjzhnSnhwMRUKp64
H62TTrIZ6QERkuYPFP8nkel3qxCvsS8qTbk9JJniWjkj5KLCejnQht2TAtWexgSm
G0rg9x3OZ+NwTnOOQwQoVwlFWZRqWQYyuysrXCT1eQgMGqF054YrBcwnz7uli714
I6fJsDogrguWrH0uLe3uHZgfsmtVFFIWRE1L89krmgVxevOvzZrQaOEyOdIvx3Wc
p7mxbXoOUBccN1J90/wnogklIHnJ3kwll13fkEwjVd3gIf3e0oNyDd95pkqjgT+U
1PPd2XbddIiVx4t2tzMSBZD3fO7YlLDCFou+4ikMGIiMmvH2RRqkk7wXZcGqZII0
p4xZEao3HRFAQdC+8B2iIpjm3llS0GBRvuNAAeckirysRW9SYAVmTG1SqmUU0XR/
n9851FaHiVBTQPUxYV1OXZEAx+UthPWLTz50yUSGvuPXffphJQEUc4bQO0bdnEJK
wKwQKnYq0Nmb4aALL5IoaXpS12K1Vo+cvnVHSWXhfMvlxA1/395sKe1w2Zp2Gt9a
6AqEuT0w8yzu4NnGF8HgZCgulSiGEbsqCNQwOVi1dwTjU2TXwn0WOfNMhW99Xujx
akBGtgJoqHbr7UD4mAKIK617aBdewiVZcA/IB2niniGBVIgdFpQDdYWRo0qD8Bp1
T7uhzgb3En2r0dXoID4nHGcHybNV+v1T0i6TdO/48bcX7hdF/P3oKvF0b+uxrKTk
gPui5JO5Vs/OSTX9uve/isgHcOI5fMC4jgKsEdQjdK+ob2kYGry7dBBsYZb3Pwyu
Bf+vVn7aJrCS1oV1DuUIuGvH0OLfuXvW2T3K6vFlagEGFAjUT69vqH+QRM9MY4TU
Y7CE3hbtgW/apNHg7mTP8sljhVQr6dlkJty1OHfNTJi+lOF452IIpDlJWOReFSqd
GG81V0g5ins9OOFyK9LaQ+XPRN/jwv+bf2s2/EDFIAFnA68AerC34wsYS7Wuz0g9
sEI4VYTqyeRmxoem92grI9nNA6TtmjCIW0eZryqSFxK67STYd9BWT0bGlkOhZquR
EUdr+m+Vqdy6xU4BE+GQl578xypUy9CUyOuSP0whkIsxD4/igM6+AWDQPIWc+Ic0
3hN0nkuvNXyw0umFBzBEr/N80bQsUin6gRiNnh0qj4wCdEzJGqxzPMi8ToYpMW9G
JDIAvYbY1fXDZ27vtwl/5xVcsU8f3alkOtMSieNhcTQY4FZYT1/i4EtTiUfLW3gy
tjz784qGPq79F//AIKXBQJyMUQegjwtwa7+dditBQtuapoiAhuAPYbzLxB0YEhaC
mh1EIGc9Wf9ZROHLHNI3p0nGhz0HWJuxQUwYpPU4PRj/mAuU8Qn1hrYQOmAunmTN
v8OeFseYDugDRc3csoNkcZw5zrKdiZt29woSvv2OD6BZ23i2N+7CNx/hBzLkaacJ
+hnIvqUxgAPcFnD7ebgyMXjvdmeT8ZDG7HiPVCfZ0STmLaQAyrHxM1MzDQuOl5Yf
9WEuq7E3+QxQen6fPs1Ay4kImn2Denp7WyRyk0Gu7Zh1b8X4I2sYO7SELcJhyc5N
hcjZ8qtwwPN349C1rZ8gQ/T+l4MaA1vepCJRQ2D5FMpVGTyRpDmEHPzMkWoAy7yo
CB3YgQG+8KNr5hr8aD8rBeppM0sTG4xLp4ZB0N+ISLIHeJRKKvtpURuVhzQUu3VC
KGmFB7RcWAlK93FfBlVfI2fYHRfv6odGZw43uv+UMIW5Z3wI/56/uz8ND8MGw2UU
mxkG2HxE+y9lHtOuzyIvad8+lCpkIZ6NzneLlgtNqraqfKpN/9qQMn2Z/a/OkOQr
SODlqh819op3EcmOR51Ja+wx5mAqDeJQRQ3j3lghCjddRB3k5a2Hp9NPBZuLhaXd
pCX9fpRPpAjx/c6Aq0ES/F5SH+UM2e93gHjLZC2B815vAyjF3f505RrBBTbtsnVj
D8wrfpYQ2nCj1BMdZJjo6yXWVj4nxNuv7wFanFqxxWtBbUvMJb19hQ73m7PoZ64q
KBftHywTbRbdnYSaqxzBEdBAlogkUDncwMOBe346g0JloKdfTQedoMH3j4+425l0
yG1hFgi4r5woQ0kIxv+FoXQvpViQBehJiCtQhASAGLxjs7TpWyiLV1w3TbYN3AJX
jSw3U/mNgLLhFc+MfuTF7GsZ/JMVuN9nuIDvOm182hZx8rLffgzfKMO37mV+xb24
LWbIQOxHI76HwasVJpU9palz+RrUMNIowh5bzPx8gJ5MwOuBw13+5GzBCWFRt0Dj
mh0/DiomRc0J2dtivQxbvlu+KiSF8yEbGh1RlKyBqNmPvJQBps+2/4Iy51wqHsHB
jQEMTW5pFN06WC2HNhtjb9NxnMXoVfFr75bssLAKwBUlSB5WGeeV3T/X9cFsbcgl
dgi9mqoq3cdITAfW3gnfTDYik3Pub8uV6LV6qggOSOgF0c7vRghLln3sO6uyqkkK
4iKW+dubPslKUwVH8GcmI99MKdShgAqHJnYo/EbLRHePf5lqay9xTu3Dv7Rez/5t
Z3+RTEzOnv/AwcUxaLAfnnRMHLqqI4shDygmdIdympEuaS/tb36/QD2oUyNEX9Ui
bkWT7VMAnod+i7zAyP2D4DjBCcRm+KxYs6D6P7cXkkYNKyhQUcwdspiDyrtRynVl
AuMJUZZMf8WetfSvTj88GfaC7B9ap0fxAeWYoKxr5AbP8s+w5FcA8mxSttqaqJKo
ZX4nx5cW4lPOBHrFt9gIQyqzcVLuF6FRLmwUXFpEtCF7V+T1UGJcNeCOorGZ1PN6
KYyq+CArv+75TCJRJOqV+HHGFbmmUVF7LuyNPfhmNxD9MJ4nwjg+YqZzwcQP1Atw
4AV20zKx5+L9SBI8LQSWVE3fuiLF2qn+LxKiceR+obE6Ao8aYwTu86J1ZCBGj+fx
vJ1vaG5w+R7IUIfZspvU72lguYqkEUO+PEnKLtY5VsfsztmvhNWP1JPsS2aYhNJB
EJNGy8cg4wthDdMGs8baMoiTlqYjQ4f+9Hxvc6HIq6zQNx9Xj2Ub6W/WVraf7gui
jQDZu+ZpEtt8K+M8gJIVO8qBZVyl73PAREd66YKemTot48C6aEnfMQGzMbA3wmHS
+4hqAITlQBCVBV1FW0ZqvW62B6n1yVRU0Ch8v0P6dGUyUHa86XFLphcojpnWYO6k
s9tBIw2/mNOf5+SijalBfpvpiFyOGa7h0S1krcYlmfrdKE5nesTM4/vZVmk4bdv7
VUGSkkOHVIpz0oCgv8ISIV9Zxk3bjGmr8nDwZLIhoJqy9o4cXhltD9L2Ntce+Vik
xNi1A/Vwi59hwUFZT6FNM0Zw4oRdvTr6NTvP3gjJFVbOPV+MAqEjGx3SnTcd6MF/
utfSzBHBR6vY4+JmHzDY9vbvovNvBKTup2xOr1RPqzcfUOQqMXSzYyadt0IgyUWk
Bk0DaO2WNzEYTXz/yeHaDQSm2nbTH/IwWvjuRkWb2GybSJyUuu9L8R9lhREQL1wR
Gz3VEBGT6hSCNnTaRDhplxGFMi5hR6tJNYm4MycyJwORM/ex5YJrUVGOzAPEOrUR
vdK3Y9jBJzPzkO1VaacQlJ83OXy7wj/qfdzIxD8TTgl6E4KTwvRFvuH1pIvGqtmk
YtojRhlhHyrf8Sa0RBgU/yZR2hpxvZlwn7xcBFXinNcCMx2jf7Tq+noKdW4Ml3Zv
8VRwX2o5zrRDKweihLRiF1qJqi01xukND+hSfdYWBZyQsv83jlcqqZD4MLcighZH
FwQ1tBAaBoDgRD6a+fg6b7W/P6jwKjJJ0xMQXa0iheq3p2LKdxotNZ6fhYXJiQ6L
NkzTyNKaDAjSv56zsWZExmmLz7FBRcAz5j2Edv3GihE8U7+W6lNBmIHqTSA4TxMT
yARrPIb1ywyDpGLA4zCjZkb+gQGRFJ8q1tSMLzIAG17+tDiRC2YZI86xePyEa4RN
6Hm8Nf2KfChcZSEHm7ykubAxxawgy6ILm4IbzEtDW6eka1pVXl2wmophtA2QIZBh
nKGT/TuHlmq+LaevjdXHZZCwlyhZxrmRvt/JRTaz70J5sg7JT6IQ1aBZEa4tOhjr
PQJ4DwcTBzePv9dRsVDYqxv7AR75N1PvKhs8sWY4Qb14d4WS1HK0vlQ6MFRIOvtV
OqgUWcuZBa1f4+/62o5kUa5obK5w/e2d+OaStOOXrEyxoS4p48NRrevM/DYR/SFe
KDg3bKYzE0hTrprFyRwZZ0NZM4CIdH/cRUNj6kB+Guq2rgTto3LfpiYw6YHpXt4P
VJgCWP3nQyemm3dQLLG01yTLU9yBli0gyctcBs2sjiJa52BSm3rHd5mlci0hSjB0
l19Rb+nWnBuO13bldtDG+FWvnuGUULdK09iw9D6MF00VEgvf4cw+3pZQvhqbeRyu
FYkGPFqnDLKJqHDFHtDxRI518JNUW2qSckxdixRqDNBKW5oIbmUlVFEfDYIyHNWj
l2yOl4ckfxTHPE7n/CaUV/Da8IIl0vbm6UqJ9nZblyTDuyfmMo/IwORVkr1pycZb
YQdiFaAqGjcfEBASWmis7FhgWHIGff2g/dtablotRVrFftBUbLsQHtYE/CCu8lVk
0Q8rlJeeeeMluwxbUQMZkU7sI+xUYyxmOw7kKl7x9Hk87n5oBFSOz9vQE/VFgJnd
RZgExArC53O4BmQ6Qv7FmgCeBN0ARZLBZ0eLc9LPxiAZHDnQRkVjydYcLVZqxM93
EOkdUDLl9MYOrifHySbVCPxVTAFcf8CDk5V5f6Gsb5T3oV6KsAgswdUfLWtjzp93
Wuvr/Z7BTmwzSnX+EFc/xB33Vcg552uRQct4OIU6QULDtgjefw/7SYhKyDM3LJsK
oQH+cxC53srgmywtLZm2zkOeT/RiOFHYr02hJedJqaCj62SToLV4MM790W6mPxJA
E4YYkqH+BFXwRj61pTa89+Oafq9cZZau9gjuahpVlxuiLpMYKr9fjY30OU96SC9K
IDPi6wg4DVT3NEtcYM+CnCOiJY30lFBUZYC4g70pFeJLESSHAZBUiw67h/BCDs0A
kQChNJ/CA14cIuJgC1ZHGqpuISnvHvQnR3p7rFqnecfTdf5lggmH7EHIlW64zg2X
+vaMqy9dQABuudsuzThosjTGH2PgfGTRuB4gLYAYH5oXqqLdRBd0iWNxM2Af+yDf
a5IkAPt/ov04Twf02tISc0erB3kgUEXckVkVKDoJbTWvCbv5Qq3xJ6xjlWa2kTJ4
Hwn4wF5i9kj5ELzQPbkJiFstvqPp8323n4jTLWUleHkj0xW8RsDYe2fzijCANsK+
aPryUw6riq+YsuJ91vSavSvJZaxaNzNOq353OblHzS4KDaChWV9VfzZ65yBz9d2i
vsRrQqIUKEZDw/yvRZGGeMec0i9mPW4Xqr+la9Q7M6ArwF9smlzjPI7AQvxNKph9
sMZaMHfqnBQuYpEYkkSq0oKxfGZTIYqAT17N6uwGbVQcW3pa0WlmxOWRMfhNadph
WQR6u9xnrXXFGkSRwYnGGxMV68F0zfTf7gALuCCMW7F/fWdaqN6G3xlnKqk1kj3F
8TI+5chIcF+lCY0cOH/NQXw6xXHXDRQ/BxD+84Ml/qOwV2XX6wRHBZn8KpXe+6W+
VOMb6D/dp2VZx2asBhNBE81tZXAIbCbvTypUWgap2exgfs8fRIN6WtspYidYAx0c
K+vktM4IjF0WgJmj5YkA+VqTAyVvmInuSsohHAzdtkVpWXfvY/FGiX6mNGmEqvr/
DcAVbHSe4hhxWHQ/8uBR59OWutep+pnrDayPF/jHMy/AW2mHfMZCt9NBXW4ah2kq
f6wOUKT3zirZPzsve665iDaCH2KH6xvfHAQ5vhZPIdlwFoE8BqVscE/BX2iHJrgm
ABcOQYT91NAtQHvtQwNlPlaB2UEV8Bzslad1bZ+kk2MG9C7LRGPlz8ocGb1tFq2G
QkuHlm3mn83ZXLg4W3hADK35HlRAZAo6eI6CVfXdfxA75UinQcEoeQWPpsjgrpCR
9QWTSO7qOk3l5g1nMgvf9Z/9NyfLow3kjjjM6vl1FiOPEhHtoTIwX46B8bUxmub9
MKRCdsIeFdAWYQDGAO8U37QY6klAh8pgSdSRcGZmzSUyUQ1nRsj4B5o1OHDRCcCz
863LwtEJ0sINAZN+G3NhwLWwuZN4kAuC05Ol/de/ulmrDJ/UEPUHYz2SHjectRbh
1yI2/KGhuyB54ZNlc6d2xtqupvaCqemPre/gbEn6aqEtk+qdCIciiCPujaUzEbIH
+meEQs+P0f//K+vuxOQanbwrhBTR9AGhSMHeyFTKAXq/V5axP2meF+JJry3LB3yo
Yz54DRW32/VaBstYS7u58eSWXM/mY7mJBGu7tFg4lncaMti9HajM1lWD2L0Iw5+c
lQhh+np9+qe6kVd2gSBeHotOivqOrCOf3/8dzNIUmsVBFFTJD+vD+UUDyDKQobgj
KkW4qXmafsIPusX9HvlQCISDO2NKdznNAjg0EE7BhlaSa/wew3bL3DLrklthtLnJ
oN7WLvalJGJRJ6cCAbbFyb6v1BiUMLFvq8BgAiNBe19gRf3CE/60TsegjxaL1bR2
Fs4F8XSpHK6J4YzIKwl9KusdDiYAVUN0cFym+hdOymeL9CSrqpBJ4PIHN9TSIzAu
Ahn7RJll8HafqnlAnauzDKP2bDnPQI3j3jO0+xEr65M32PViVM7tGH4wGVyDH3cf
d3hEidVCBgWXRnsAPmuh1/9+1OpU5tkVJ1LwTj22954FGOA2585swJQoz+GYRxef
iURKapBzPHZQMKySBdyLDsRNHdeik7FRNsgRqWR1p2amdfI006CUgD2YxGMWCJRG
kJcJaGKGMLbN3TunR8uuANY6/o8D4hxmE0hQmpweN9E1v2ElPFtYSh3aNls1CMcx
xfMr25sBz/MjP/6kg+LinfX/IM+JMJsm3EQUypHaRCIZbx3khTiEQsa1yrT1HpSd
cePdXX1EKY/BfJ9eQhU/+Dh6pm5IVcO3mcOzgGqB/Kp3cxmh/OrZOdB9+pQw8rpj
UBU/2BTPgja3bCWAHa4jGFW5HbYrIV35pluL4K8tk6dmfp0RmNXF+fvQKhGlFy+u
5+4R5pvk23UNG61pWw0wW795TIHm+zkP2CXeZHBR4bAlLhX2oNmsYESsbB+MF4IK
UBdteTbC2yjqi6TN2jjavHzA+DI9H9cvjEJs60NehdU5C2kOKFeMiw+4AN5M9Hnv
Q7/1XDvMMMYGkYltn7J1aiwLMWG6YTdca6DL5/nD7i9lT3D5E54pF08Xz8IXW8XL
p9eI+eY4c7/+6MNKs5kSr5Z8QCxP83wSty4QWtEOSDDsUW3EQBbDkEy90ZQsgQeW
dKGDkG/Vz9jmDDVWPf0YtxvVCr7UydMad30iUrT1bMbU/3mlSADRGUnrWGPUwb2p
wg8mo0uusmpLWQG/gm2MuEwmapCA5EppLaYdf3qbN82Hf3eXMAbOvZPXj6AcGyL0
AGKiTyACGJMyEQHh5cvHcWcj67YjDWGkcV48MZzqXuxRwhfPm7EPfGK3IIw5x09b
GfTmbUX7o/CQxns1IG1abF/gkHXmmXmWqBI0MRXhJ2X4kI3wEiEaqMnY/OBBHJOA
DOyt+c0q4dvQOFrPPmDQPvN4mlgI7qOhqBtsdTPBhh7QQDu7aqB/l7YBO+GqwkAm
O+jN9HOBWGshrlgQCUQnBuJk9BHECwUZLxF1x87BReo/y7FI7ElEd/GKrrkojos0
J5erKHdaXw/JYnrKbr2Lrw5OunS7AHz1Bql4P5UHIQScvTbmpJWe7Vw52C8sNW5M
3xiKLq/1pxV7Ndb9AgpzkCh4Z/W96IQtqK7n4tbZ0dDVX2cc0OOI+QxG8tKkszG6
ZfJsvXmI1mm7e77vek8SzuAi3SMENU0ffOkjyWEamwPV76hO+j/jgMyPC5ih+Gr4
hLXzVGKR8W7/7mYnMS3wHZgJxOwpOh2V/4yDVGZscJ7Ob3mdsTx8lShwllJcSXG/
c2WkDrOZ8CbE1J5jsUyFbxpeBnAPwrAU/+d+Fb0v6D2JSfHQR4+gMDFbjvuw0eLA
flmVUjPPbAXprMvYAn5hGqpGuJ7GXMQ4AHy5wMAnEvOqMtWG+Y5OiWeRKcTVGKN1
YmTyqXOFvCc+eWdogzMKbppoujt+EnTKuvgVIPtY20SBb4XiBj6EGo+PnEwKpnUQ
C43bsMqSG3TpgoivSKJhKlYOsRfHkokGbrkBn9tdD7Pj/qjkWoSIbjdjPgL1NfyZ
tDRqGJV3NrJmyDcuYaCyd0/cT6vIg2zX954wpGAUqMyFIaCnDPRvOOmsg+2o7Jke
VruGGtoalILnz9SfOpMIVjKA+7wxh+gjE+zSlHzS8NNT9ntZaEa/6hICeTY0SCl0
VSEBY+T28vdy+dVsn5R70Sj2bNKHAjyRL+l5dYrq+FUZWX/ba0U/Jf4yX1IfFzLx
pCqnliSiATNsFF4O5Hl08ZBT29J3mfrYmZUvERbrnxohXGgHsn+GikyKdgsOuM6o
9DP2OVDKtvULUq4Nj3zvY8rUALJxGcUaUdYlQWVrceZNJGp7JZu4J6k4Z3qIUS2C
y/aXEV6FP6lW5ahr3e+9sL+CXxlGKjRNDshlUQfS7ai9MHHG6VsMOdpn0/SlwYQ1
7WBtW1FxsCe7pKiO6etteTGW1pKUWwfltHq13Gsefob9GZTSvN7ZtUdG2PZ1EcY3
ZSW9cflF8uuoyotSBYv0UtJjrsS65EwKD5IOSAkaP4XKaWU8LlitOzmal6Oe92gk
+N10h98tBuks5A5s77gDMw1MBpxxJUHp+FX2xLGwC4IOs7BNAixixNJ8zuCIwM0Y
/EP0kLSqMhPGUUjCEXy712CX6RjvGqcmyb3DGvDDo9xY3AYfJtBlW24WIgLYaFsV
Shk+IoHhkgOtDvO++8bL5WR0xAq40qRUr5wYdEHg7TTMul01+r86+wuUORDs1mZv
mmxhzJeh47gKXx7T62mDmrIUAoR2YeriXkzxzBbSkUCuxt7ykdXix3U8QW3JxHSU
icYCvsnjBNN24XhQCgTVn9LB9jNyEdhdINESEJL6R9QMyf3yXyQbabsxKJsnYDpY
CpFXOvZytyBhp8aroOlM/r4833MzwW4qO5rhBLxKbestI2UCUk+7tuMsGCCo2NCJ
N6KdIc7inC67PWuhG0pnOrpsVz/CqH9SRY1lCSUqIr/T5IfuBYRP2r5qgc+b7iu8
+3kBCGsM5AQURLBXkgV6W832Iwm0NlNRfV0c5D3mjiD1BjPbwfPRvX+GqU/R2Ogf
qdiQUPwasoqbnJJ2oYcUR+R2Rzq+xzs2QPj5KBsoJqSj1Ohfoi40OkoDAZKt7mP9
0X2qMI6AYyCaZLwjLjjKRItsAGK28viQhQGcMjx7ycXckWNoE/ZwKVg8zWE8xDM9
f4UzXdWomWfBZhEe3o10eDeUYK9QjlB0aIJ3kMAtrPEfTL432fwgnPc9CPn/IHE9
t7L6ewKJJBdIU2QKkcUIXOtw8ZIZaIMM2pvyvEZC6F8yzQ2JcUP4iY9U7DRrx6JH
4QHEa2rp+XaeEQnZn9Ft1Z24/77C6lWB9gH7xPPg2ootEjIpN4Tg4nbN8v9+yAUz
wvliYyshCgJkhoxOLA4XG5BZ10aHkeYAXVBVpf9gD01UcgINlksRnptFRCw46I0C
Q2tm5+jCiSGt89SEQ13ozLH7UaioWjWjhkmvN2z611GQQUQCVA61imJGQY6JZdEG
FkQ/Y4VsyIUlR59BiyC1gW+Z4keAdsGoNfE7jGRSQQWDbyI0DD7i7CChuWByzAzD
cRXAgkStBkwk5xFFlZKC0dtXfOkk3Mc+XKDEmpcZNQoKeDhVnpFcZOWaIn2R5PI1
bVmYZiJw6suWKRgK3ffZmx3Oe3IP5PL7J0tP3DP8YJvKIatk/6kHLZoEon7wT1LF
vZZwNLlL1PJl7xoSAfOQaCLR0DV1rM2MLaGgA9WLx35FRaCOoAI+zmfx06S3MtMo
cZtYsi13QkRSwIAShPYgLPd05G+BijnqsLCbGQveVj/9WEV8Y0nNsp6yHUWf2ZH8
zHb/O7sLYffXT/i8oJ4gNQSdaaMc2WMtDjOjZ4qfP6vZ2c0d9F6Pzo4lGAF/4+NI
jTq8p6wwXM/BQu+gIHy+yEYYS6tHNM0ULHGCZunEy8l1f5j6FlvC0wBaRSfNHXoW
/WjDs71A84wMtJDUcZULZCRHwh/KuPclJaCOmPcAuoJ5kHwGrlJ8JuAhbu5pz4mY
XfWiC+XWXTUouxbNgCvypOZQJ9UDso0ZStPcfJJK9SpId/FNnQ070WB4+LcGSU9n
ay/BXrQnIInY6z03quuGQ2SdeEPuV3YVZZ7L4HfRCy5LkCkNCMDlrGAzjYH+h1/p
rufg7mdpCLf1gjGDlvy/KMOtb6vitDTdAuJDdZ7fl4QYmfkQbxikAlisn2SdsU84
/b7nPSaVfVY4y0KywVWfB39rAGsc83oaVVjt4c1C94ahQMsXas+/fVnpVZoan+Ap
fLfzn6E/ez77ZnnPeregpEZFtflkbE3Cwxa0f55l8txVvbxizY3ZQpcAA+Ev0kU4
7yF7u67zwDokYZpi+d4Vmen4WGvhAb4GMTXcTrkNd+1EK1DPb9TV+zwn7oRmDk2S
VoPcTj4GTlz1sNQ5swNRVZhn88qIegnSqK6/aaAL3gi5Gu/TdHlGbfJ5jUVU2E0+
kM+c/WXM8LG9a9VTsg7tU2cv/e1ImLhgQcuYrTbTPot+C+bdyla1SocGqKobnOD9
WRR66hoE/8XJ/HsmwDIcFxuXoQgeiw3FhXtfXfdUKOsh78MwXyAR8EBGzoqU/g7s
oRKve5k62Cdaa775gUz6s/8HM9yr4AhG/mCGLFI/zMfGvi4QSKWRZtF2uYJpwiyJ
Pp6h9p+olJhtl7Sv1Uw4l90PxK1/cCvZLYpNU3L9EhQNPdutR4+Vi0/lZqLzmV8c
h6vvF3/SlJy9DLJAYs4WZrBl3LpcBWM02wkEL7R3igPgqzLZx77wjoonLIB09CIk
eSZmjD8wp5AfW5Mu2xn5/xwVBEwouuSdRZb5Znt6Mq/R1Q+K5Xp/vB7V7vLOr/C5
1bhZqQXbBPhXvhtAx1eXpKegvGuv4ML2nPmNT0Sa5TsQzpvFd/AhfJw2fCxwX0xG
eRdqmpdO/+py6HxRHRszXbhu7iin6P2auAaqvf4iHuuw989V9RdRm2rCk41qkimi
oM9HJQkoeZuDTHCTy73tlJohgRxtaWG3uSSmpgYyyi+IzRzV9nJWFCCyZ7dqO5/L
wxQkTIWLGgffrZTeEV1Ik75Dd/GzOX6G61DjbYFEJQkEf4BbOgbKhbVMvQniGvIg
78t9mUDdlwGAwXYAQKn2BGR4vprqtp2ts7upr6fA7ChLkbWKq0VD8D2AATqIxo8a
zNqnu77xFLz4ohV4yZRnX8Z5nVr1BCinrh+lCeveKTRKZ9kctuzisMi00xcEtqtb
kNcaMjdMPKGh6qRqBc0pLBpk25vXwrXBpd+WnRdcH++H425VbDoL22xmczeVoOjx
fOd34+vUgKnrcianA3hLf91TcoNvoAOjqs9qrl6I7jH5jElauikMoIsKHyFljJNX
duXSGxgP2QM4hzXPjU6ru7fLm2ddqLHDBHParalJMz7Vw0XR1Ck5W5GUnWpWcWKY
ZNllH0zKVsvaudcN/PLHoi1Yp51gXCzQ1xdqK9sFh7UNAD9RVT8gN12AIx/qXu/x
ee7gttDxh4M9S6UEm2sD0/enP70uxbIflFgdJnJGJwrQUcvhAO+pHV+UnQPBdNj2
Sy28mdyB73VW8GGQ9XgXGpRJ82c1P4+5fdzlp6lObqguGMRteP3hTDvSaR5sdkFJ
7kd2qEC4Z1KYSidUTAkonHlbNLtvaz5nQ8Y8F8U70mZ/P0yd9yyTk/o85qdf8n1V
Zt9sBHsedVn1gjOdK9/5ljwRD4pzAio0OybuNjGG4+KfeP84kPOCGYiWp+YQeZXu
1BFXBD5/dkfdOO5HbJMM1Dkro9YSrKAzuOhnL8oAeND6q0658wK3+ODVUmbQjX8G
zWYpbsG/T97WfMzFW6dN0WrWPtCnxdEa+DrHogvWEG6MfUttpgd3IX/75m2Ua7/Z
JjWaCuCeUx/nSS3cSc7dugN2tOPiarJxnfpUI8Nfe7BrkgfEN1olaoUTR32zwN24
CPdV6X5VnuWhcpKb4azcfkuvJMfwc8p7fSNyx5sE/knRIPlOP+xLojJ6kbekkj3b
+cH1teYcCUX0NB1GI296DqZcaS0vz9lIa0IdbPU5maA1mlGlfPdS81/zGVWRzkwG
7kxW3B2hd0OjtsHV5JT5/PDIEJgycQQ0FWVZmY3Zj2PdcWj5p2NHQGnrjJB4umNy
3bxcKCJqkboBq1T8y+eqGIXZN4VP+fY4l3y+gGxE6sWAJLECMl0rT7wzflVk36kb
QkzwfoqoltXzQA5heiMc0ek2+SOFcJr+DAJgNcTqvHbWC1K68xryiKfOzMyhg7zx
rLHmfKUxkOIU6w/TBQYXsnLdWOFfYRu8F2SBcjSBadBj69o7ED0syhEzQa1KxcXv
efUPx49HM16heFlLkC9Rumv6poJ75A+TvA/SXj/b+8sXNRoWhcEUbJUvYomAPCXY
YztY/VxL0CkFjn/K5YQYCCKGFSLhjeL+JpT471wQnT7bwx89upI0X0jh2RTFkP22
ScLNOm29xulRVciZHfsxsN84OtCh7a5wPI/zGtBY5ZdRsN6Vt43Mr53HYyJKmumO
YR5jsNun7eDCLFQN2pq13HsJjrfQ+GpBObv51LKNOGnP81hs7+oHARLTTAs2DDHc
uBFJ/XuJbYIMJmX4Vn+9ecJ5oqvnPdSSR61RIqOHXnajmi497N8d0txly/ufzbTr
FXFoH78JfK5MVx/vVd2WsxR4RylmFuSaqDMtIdfc8LN6y/eBqH66E3k8KVcmMCGA
QUHHznfBU/E7vH3CqRgQC/cHPE2r2QcTrV8oVdMeDete7Yrx3buB+mdtpwBxsVzB
7kRd9YQcbtlFRwgTodsqXhHlmfSRzA/OrelP4+O5QdjDRome5bpXgn+iFzYpAyor
4MvRYdSRoHIkwew8eGJgFMDfZ4NDYbRLFozAG4mSWCMepcvA+rSKevVNT1latfiI
d/g3S+igWhTULzCbl6XeQOfC9pZ70RkoPnu3m7THXhCN1L9K7W1uOnnJ4T26POj5
vNOGs0YfcuDHbR0du2sJCJXaEhIlsz9gZ6QGJA76itxKMXK96feKJ6kGJv77gWRg
fUq5B4zCfALq065363kZ3YDdxY8eh72R4vSUmV3FFflgJGp0WjaDiGyXdDseSu2f
SiRm8969NPv2XzQHt6B8o3AKua/ybUk3bs8TCD9LxG1ql2DcwG4xM3q3Ap8eCkno
obeSFjt9TRTr55ybX88Dtgl96Ixe4KtImCg7IQDAsgx4ireyB+jXHQyL4fctM8bL
i4VG79seBMOI0qaBFqZ/3OO9Y8+8c45YaTSnX8FLOuP4ksJ3HVAqLkP7wF5XaMhH
Gy4UhTUcwfwZSjS7XHziFDr9bTeUFL7X3X6XayvN7q2OjA0IRK4vtri1xeWiZ15N
mklH1gcs+Y5Sli8MTfjgxGd1Itl9aWYT9J27nO0xsqISLX+Z1fgiUcAtFXXnlMai
Rb+G6kGr41d9AjtK3IONU1D2fZgBbmsOin2pdBs40ZA2g3nS9oMECXpmXF+CmSwM
1stVLGR0AiSYMjceLR+LrZKjZvcIV5EjXxY6qYWT+/eiDVjVKLYY8/KwLIa+3Qbc
8KrNEaHQtCErQn7VXc4eNiitqGSj7UQMGm/hXBvQgASWG3A4xI5QzcemZKUh/1WG
Sv/ojFNcqg6WKEm7AG7gP16y5wHalLtLmtz1ujUQ/AEiR9lTCdO4yjtfS+dKh1gl
G3lJPCnaNHhXHEc99jRni4m8zFIakupjW7nWAgbPJpkG8ibC83GyBy6JPb2UDBt9
MIAFdlJdcjolnlWeU6Ukv/sBqPBiB7KGuvnSTW9fEU839MROeUU8tlz3zap2F5dV
A4sKBd1RKqCFxjaL04W4/woYYvMJmbbUXJO5VWPuheGGsNusa13rlRti1KIjYZVh
gtM0OIIAJ9hr3KcKLjx71ZT1AENWB9SfYKhZ7QaXDoW8MCu6+Ho3pB/HWsA2gaQE
e0adAQGtxFfzqQhGIyfwUhl6YcuIztdPUMDS95EqdqaLXlCDz9+YoX52+YDoy3mc
IGJObzfEP6M3HuGX19K4ewOIv1JP/64rDDo0q3voqhkJyMFwNx3vrfMRLLubIOJP
cTviYZhRth6XXgySL4fvL2/C1XLAE0TEyRuyD+lq4IdqvG3uA4LvxejKeUdps51t
9ElurqjtP4aqEDmlWpjXjQG0Lj+t5XwRjKQgEWkuVPYlOqCi4OHOcDDV/D7HCRpj
S70SPlLkhd3AN0SHdYRZqNxV1x2YJSEN/5GUu7l4f7zxRsLpMZCOLVT5OkPaZZtx
7pKcEhxjY0u1JCQyNl/lCAK7IblcKF9asI6MBRjXFG77beqRCULf2WBF4KnmpXJO
z3u7FAx2xxHIfaqo6Apgje8obBREwoyjVLI9LMGVTwiIal1IeQ5Fm2vbt4JWhBu/
eqk9DWZqB+z4ky7O8JOmU+Ad8oN6x+NdiQ8JD3wMbYGDTMio2ENaIKG9761m+N4v
CETaaNeX6DgzhD4da3cDllUucOU+qVSkfVrRzjCX6KUvy1/Lm2B4wk4AkTfDd5T9
CmaenC8+LDgkKYIYjfi8WperQNUC3X/ibICEGGHR6dEAJwp+zmbvtX2ZzeyBfaz8
4l4ifu0R6JKZJmXuCKaQwRA0OGRa1HgKdLkdv/1OStNt2HqsgZuz/ihQMMOCrr9Y
qvSU3r8uJvdFKnAbCLdLElMqcVENyaEC8TC5kXdJ1LTqVQKDffncNKCHJCFDYH9g
aZ+oAof8feMivZqTieQ7tOZ0ZBXvZUGW0sAOkHgusrWQ1ZF7nF99hFvXp1aE0NOl
FOGnoTW9ZeT8km5pKcKmjT2keYqccnY2T1x+araBWONrsrqDs3tB6IYlc2KXfTin
fY/iLEqn63I2S60Ji6O1CjtxuvOweqIc50y/6fBnP+6wBuNjQrjNeSb/nprxZxY0
sN6I+BqO+HZaMOa0SYFtPwcjzRZmk4Botk/knfrIRJTz5394TxnMV6z95DHLJ0aP
YlyHjuH0kvBwaD0Aq8vEDXiGtzPUFUzhvnk8MEZLsitab6u/ywRv8cflsnCPIKsF
tDE740Yi2f71NMPgOTljNc5M9tjw4uc7138w5HTLmz3v058Wv+7dmbr1bwWYita5
nXQN/QlZKsz4JwLTINCvu9ChL+dmPaZDMUbxBAAp8p4r3dIWLT3EfgP5Ro6idNjV
g2aW+whgmJhQ22eVz5ZeJagOxpaVRUGWi0ZDHlx3VVi2EZ9WWP2v8QN3owqaQ/kF
AHN575uLxBH1ds0helkEB9MBUAr9FXjYQmkg91fpSAtLg4qQg6uzpHytbjV7aGA7
Cisrv+dSJPTEOZnB/j4nIBkOOUOEK93vcyPG9GK9n96VcnKBOGnU8hRyAaEwVDcj
X3nvNoLlP52NLr5r2Z+7vfmRdA8+fa7oKHxHvAV2BmimPEqikKzxBkhv7kLjcHxp
UCKQwrjJop3xUtiFDcAhctr+L7KGgDfRflqI/BGnO1vOLT/rNg69bDMtSWvdpilL
1EHcbFwRvTGkexpnuQ4hteBiuXiLbWFO2H6y7zNSo6Y/GvPuudzweDjKwTVnUeK8
x0bYa5ZJA0cTL9XjulK2z0dKcfoybiE5taKuaYReruLiUOBAUyU8ByIzFpp3bMYf
Di78uCKawBlMmWLeJgbNkIE9rovtjmvoezkQR90tiKQmgCnKYBw2695+vGzEUsgX
JHRa8XRP3it7xCEJCc1c5dAbg1+RBuxv5/Fu2GKgoP0TDZl6MqHj6EA5R0GCkXjG
N7X1IUyiqVM9ebGzCucC12jWQlPbPhlEsgGK68hXDsIEH8lHj9kLyxXG0DDScjtz
6JZsfHwQDDKUBTJBFo9ybsqxT0aa0xbsXhwohhoogB3IPkH6H0a5yqADCDlFL5uW
KzYOMmmg4XjhxxQ/ymUTG3bk5Jgd5C3jKtn8J+Adq8yi40fUKURbV/pvI9UlCS7h
Pmc/sDJgGxYaIc8CBLl4/fHjfL7kaAZoLkazfRmTSup1gwaKVPrZpLR7Wk9QH6Db
x60f8LL9quBi/D0ayH075PmoM1CLaftqlhr4Pacy2OHF6uuhgGgT2ome4pF+HU2L
N+mt/DJ4XAytU1HW3BdR06OQghwSEgKklnPNnKVJWDHP4e6cgZjYxhkUnfGzLN9Y
0YepwtpsRRx2YL7R0Jq57nUekLDj/th57hIGKQwNMbCSFzaMR1p0KIWBjf4GKwx8
bRFl+Re854l7vQ4TQMmB3XQGnPkg/dqMrY8t6gwDfOAuRiVkKWzSeovjE3ZazfU9
pmFhnCLciQSypEl+Tzq0tYNrlY88bt4KFElc5G+ChVFVG+Jhf+kvBRgGyyeZVGqZ
MqkdIQ3TmAf76Pu8kBq3jfNFoUfxk7fvmT1NES2okobVjVib5NN0kNZfaLtGcZ9D
du8HDHvHtPLjo5YCFzM3wr4FXKS1wrVQBIe+Lc5/r5kNtmgiD/a/x9w8C9der97z
UFr7ztatjct2glrHDosSCnAZx5lqYuiwETmz8rnJGP7Hfl2Mr9uQ8MBsD8DJXaAI
3AuXnbyhC4Mk3K8WNXixLep2LqqI6dK1tuuA+qXgxZR0ZOY0bIh1wWQ4PhhwsEBd
FF6SXPRSzUOF/DuDOTICA5kIJHpkJzqdyB3gRS2Y245hEvv8Tt7t4CYZ2PrRaSlY
yNTWP/t1/FvVyZjYR7RzMNPkKOvcQcuvgg4Vcw0uG22KdIm5V5LEiJxuhQeQrPKN
Vw41meeJuZ0IUPJ5huTM7yl8+n8vnhDmFS1G8O5Hk4DgwxftZyPj3UtvxdmIE6jn
/EE8hc59oPjLAYnsK38ikO145kBEcYu1rFP/oTCNszRlceIARtVk1csYgbwroQ0u
/MqsqQGXfeEx5Rl3zbU824shxoJPILBlQm8qPw6qnBh3gTLJgMZ9SDq92FRiXXVR
SLMfX3P2zinzFB9lGCwY1mIbAMgwp+cUOH+yD0YvOQxJ8J7KW4960pJknJQaL2pT
alPf8SRoOao38vd5ESoSfMV1KmDWe24F8Ekv+UZd+kKhaVoK2OrKQsbeIHZfK9JT
m4r9mbK5p3sLOrb+Cl8VLVfN+v1gkQRVbNdfuhRO3jeziQ2BWoog9oEpt8RQBjZC
C1MqiQZywYunbQpXYnHsvt5iP5fBP4ROg7GRkUveWC7e1UjQ+eHjSRD+k75KKdXW
EHFOIMCmlQwe4rYwFJqyFL9GQQ62Ik/GhrE94AW790ABo4oZQ3cZimuvR3E6b7zC
ZImO4hFWnJIKL6A4pTpPfM0o2M3hJW4EZ7w/roivchCzTW2Yc1DXqUwwYywOXhYI
lfvPpgfdSzw800c8aPeLZxJjFbjQp/KpnuLvLXnq5DPD2FQ6s6uOxGocKV6ib7Ea
JT+tJwR8IY+p8P6AUUs4Ur3v9zaxd7jKjI/rdKrzUqVjZLgRtZH9sHZDFqzanJjc
VaOF7yU2lsBMFiHD/vUmjGy1xXkQUArzN63L9Rd4nzgHwPVWS1FhKwHG+2S+4IWH
rdnjfZ5kJGWyiYMk7luV68F92dZMr1T2SFxwfx8YEqE2XSTxdM4y0WCIkgFKKef6
dmqj6Qb9gpSatNE8Dric4jRWRMlNvsm1J4nlPCi/7pHC7BMXZy0TbnsWF7UuYt/D
EL70ZROuD3jYJCugHR3STIPdSmKOXdJUl+OhTUR4r3I16LI3tcEQtL2guCjPKjPz
CzWcWmxbDuZLjGiKsVRPjY+d8dAtuNAJB4g9jMnkBVjj3qTf2WUiiHFb/nUM8YWy
h5LKy4gIvX8kGoPs3e2da/qRo6Z+R+r3l5mxAEipRCgmcD3Qzdljba546pB864Zw
PGwFsP6X7jXEKdtDquI4uU6+cFrqPmei9BnXNy7GNpRTSC3v+jiUDzd9IBdjlx13
aO29STzjxtYVUltWDxaLYUQVKmojXR9aXKeeZoFl/GwltqFDz6s2hAq12m/TNjhJ
fKGB8yQ0svnOZ6E+uMb5ALgHfSiwbC+IG6yA61xT1HgEKEihu/s0R7y986/AtnvW
tL8Rz0Vv/vR0+eghAAU9HEnBehjB0dK0GHOasa1oT0HCeWXEZNDWWkaGlJSM3Nhj
S09Y70HM9T+e+k8cgZMocXLv+gxPlsi8KHx1Upwxg2hKLEg00YDEDhfQTpwVdDQX
DpUpBhCET0r73xEuleWoWibRf/LKFjKwAZxh8UQryO9yf1kMYrLY2thtP5lcRvgU
nIf8x8w+pOyxAUSo7KtMMDwXWNnZ6cpMavf5zCK4oPQqIhIzNStY3eCQjipHa2sW
a4255QB+IIIQteXriouJH5Z3q7Ph0ySnXkFwJVbvF7OcaL8221qFLjPEicCShgeH
EBLcdQ2pcQtDvLF+XSKMWhsXgxuZ4B4n0jXzvm14Wu/srkGrIWLevG4Y4QmC7gAx
8qwocrexuZvercWvmA5fhbSDqYs7gnIyP3zSjGiWRrDaJo4Xcoqlk6aihiY1pzJE
UTq1nt4R7KpptsMTMfL9N1zgH16e2kz2cWJDnUFg/cRFQXL4zw4oS4BjlpRhrsHo
hsfCmppTNQIM5ecm2TWc7xPILffzvVOHqPly2Zuje6TpNjtbgFS+3cLPho+WaM+n
UsgMPpDdZZf6rJ18GxKFgmAWG9KYUC7T58XeXsW6pHXl8ck8m4GZ5hMOFrEmaVtt
gsWw/w85DP7tfjF4kJ4G4yrr7A1cBs/8p+ClnDU8sJLmyOUm7wzO8rEDbesFvAI0
P94hw7fimT81MBnK99cFttQnaMKQKmVK0xdOTj0x+D06607j9u9tpMjQ16/de7gV
l+3VQ5GmIWQsxLSL6SDamUf7kxnDr81PlwQxcPrmND+zkJ4kclUqWAWeP7XXj4Lm
jF+4t5M+8Pgklgiclrdfvat8so24kQlFQq7t1Rfd8QCxLYd59MF1p2kZQW8UKqY6
l4/d3OZPNnnFsKqAKg3YH7pgnZB/nMNxb7F5yJpkj4h5yIjc76NvnE9wq/4viKIB
plPyuO5Wmc4Wzea1tTmmsrXbk0d2EbqTTtAH35+jHrsuTWfrVuIAquNZTd9WVd0o
iLIK0XH1DK8wrXnyCl30YfzraP6xT3sl34aO20uKaNFHZRonsvPTDR5lrgVO66A1
ANPp+BRc6sPKdkrd7SNECbYTeJdOFjgmFXxo48Jd+5H5tVO2soXs2tgLcOa6Nidm
F0hyA0Blf7h0f0DrHodh1C4pRyga2iNl2XIwt2gs7ooTgZL2bbijHRD8p4gsNEpy
theJm10BzdjR5HFQlt0yMvkIYAt/VVydDiWFA55DtlnPJjeo9QQAFfDnZT7pvT3B
pGgbwWi0sJ2a3vGlmgw8n5Tbs0rYsRGLJA0TUw+qRGzjw1B7ujhhVhuFCOJBb0yt
krqv7sT1BfZ/fqvFvel7WJKScowa87smYpovge5mNUQoqSNFkLaRFygmnB5oqSNl
2lyvFBr1ppE/iCJY/VTQhnj7+aV76rqRV4Z4yECbpK9BPkzPNyl1Ny5zX5/cmiEM
rltr9J7h2xJAf2BiMmTwqgq1BMqHwRurRHsoXrED9QWUMCCGMwN1oVvCJWU51pue
ZzvwIuP8jcSQhJJBNnhSEjI7N6u1yOHHH9DT6VG9QGnpn/o5MdrpW6K1cztjx5oQ
CK77SIajpTmCaGlx5qHbRfi1IfIgFfEmWUT6KFHahSmc5k6akWtXNKPFWE8wGYf5
>>>>>>> main
`protect end_protected