`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3952 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIbuMvKJdIj3U0+AB1Mzdyg+tFX4rCc6Fk7FGLeZSyUa+m
cApTAlemaGuJQW+t0PHlVTBhC1nkOlhP44kzRN42X8g8xnIKIHSZpqoVwfNxKb7Z
wXNbomaJb+7JPNzScld1/x6igveVW6IcKlPfIIs3bRXYlXzvqT8UEQ9hC6c91oZF
18m+AYyv3ua6YQ8qqWFsPS5DrNt/p7jtNYCJ65oMSruRm8qrArnQZJ6vljaezfRY
FPzseCxy4OQ7y7euQ4bjMmcNN9rNEjnRC8ldksJgx3lnPdSYZJQu21i7Ex94yvFK
2+Qb788wiDgUOckQpLE5VGYyRNmabN4ztb/Bk6mY7WNSfmSR4x5EnyDm/vsIH31o
6+KtH0nu0edqIFHkLXrC6INbeti38yX7EGUypvHID/WkP8VqAeoKrHynDfB6+otI
8ndvBQQSkhawQW+LKqaTFrChB1Tkg3z+MWETf/860IssVB8bcYTrlhBL8BA2I8ju
cibWfGvCxEsQWDmpirfaSJ/UCbEnb82WjJw/AHRcl4ZncWULhAviGzhlsrVTyDMy
AoFabx9OCQT3RydeF0X3OtMviUdsdpy94new709nkbaw6VGfvsQ5OKdCv1xFy1jl
1Jf+CSadcwMiQyVZlw8BUzG7jC7WAgWw2I6wwcZ7a93UV/iQLnkFF+6l8b5zfNmq
lEYg+lccY2x1XXRv1HcSl8oRMXILeM/IpsuVwznwsp3kANY028qGJ6/GXMshqbka
31uA17JISRP+qx2xdPf6Ke+RdTsc08fLQmtJsVsXUpjOey/5VaKeFXBptl9CHx4a
ldpeb4YWt++xz17/j/HHEn+qPsqh2wPLS7VsVHBEcT0rzcjuAinqYRifKREoiPu8
nKgqntD+hvOtVXRZYuFE0eDuDr+2JkpjBVACHbDR4QCWvZIBJbZvRS7DKzvpoDAE
28CkunVKxRbuUsbuRRjEL2APZXVD2U5fIxhepRt+nnC8keZ3kjm6RuSFZp9JNmHq
f+EYMtyjvqHN9eh9n3Bg+xOrWlzfvFE0ng+V+JWGznkOVv4bsCn3Q2+W+lwqJ93H
FJX2gNI1c8vg5IrmSS4nj1QProKv/CqRjJRFM0IwstaAL1kG/s/H66INpFjfExHI
A+5QsMv8dq2cyJzeQeaFwRzKIZBdXVvKE3Qym+cnDSh6rZau6v0dRQLw6k5TA/Ft
DYG0/FXSkM4vejCBcjznlqeFWvjiEpOVXUqNaFaQl7wdZUis6t9OvG7Li974Z0+1
LCZJNxV3ppOGvurA1GH+LUZsZitC7BXxsdl1pLF8PHmYi5MSdSWSHoeUkH75Rfs/
F7CFK8fZ52auRcW3G24mMiUBbCpLuq0+EL4TW8veshKFtPI4G8bZazGKZ/RovBhw
UzALKk9VBOkna2Efe4Pz8YZl9YyAxmZ6CHsXaSbEHIZEVnGxe9tHpvavuKKH0J9R
hw2bCN8qDMyweL5d242AzoQRfFHEGVBxyYbQzfoq2Jo39LKEklqqYK7HaJV+5tPh
WwieQzGwNhHIi83UjcsBsUXrcJJMxjXz1sfolyEq4A94/LNaIBGoaU9ns3XwRWdc
Aln+iKopEjg8h3MAEoiQRRzfunLW8jobvD7Vrhn9ZXGs11x3HWBpnTqIGe9QUJwo
1N7Nq3GY9iZBxGSSJ7Y8mt3DekIYiK8rqcU6K36wXfwHwjbsA8p8seY4SJLgy/nR
3z5rB2T/Yu/Xn5+KS4EIqbHix6fP3FYmXFV2jH6Bwf50cPLTePbJzdvZ5jidXyXe
wFHAeGXhYLsh0qUAYFQYmUGR5stWojXh1QvARsAc0Y/1tXH7KXzzvHQJiom4zz8x
i4lBKr73P0EQhyw6cL1AyIrtyz2bDm0rQ/TyIW+fRH8b7HM4mQ2ektiOChoPPJWP
OIGnmtuIFlOjE8p8SAsrRNhsRV4/r867kyWCpePxxMYXnm9tJLLb9ESF40vgQ/Qx
bgomYtgiRx13xYm4syx5RoE6LQ64CrPEmnNK1zoVQyYlVmMugIzTvKAhjaJDmBg1
6HuUO/YCE+u8eOmIx4fy0UT0hCqWGgUBAdKYeAWLqFuw1wwPx/xWQMOlYDgrCmhJ
Ck/e1e5RPMkbKFArLy0exIqNBH/GUw760FxeTEtuYWctCPRyxuFgMT2A16JaECFT
CC8FusDw8GgKjrG8QqYqh/bxxtV/bI8yB4B7ihz4mbp7U0AmHnWZMH7NrZ9GciA2
cKYcDkT8iiXrnROo1NK6DQEA2bgtAxxPLbH3DxsHcf0wTnL/L5X5u/5HJZRkfOof
F6sCCeEsMbYVJCsV+TRADAmRIroDcSpVMiLTwbUY1Vq78oFtE8OGHNnhPcLuQmWu
rdowPSo+bXsxECSajL1zwBlvX+3qfJOH1Bt3ooi5Cr+qmC+/zAVjRpwDObUGwmMU
B+kY1wAMa0MpR9gz2UnScEiEoEGgJyCFUyzjNhaqP/k0QDchEIG8SBtr1eAPvnEj
bFm4R0d6Z4ttJa0JmzvSr6SMeeKCEpW0MFhgQq0bEn8Ywyk6WbHGd5fhd3JaItJK
rN6bg+rXsuGyxW5L1/SzkKc+gkyT2mMHnIvgwKVHsBust3diLTAwWDI/7YhQopU8
O/JOKXyVipPahvRXbc9ioKC5yRIaS/iTQL7wYVkoHIyvTRvofg1xGQulJezhOMf5
qnIe+pgk7X+1vdfrsEhPCWSSc8f0SkieufmE4lIoVZHPQpWo/GnYscAGZMqLPsRx
XskvJ/91lAx9edrfkwBzc8SQpXPNG4MnaYQqo/AitlEEa10sOuvz3PRMGhrctrtB
S2+Qz4SDZDWTwygkt1JH7ByVvk8+0zRbnE+V2ERTZ9J5ItEN0PgzHc5HodZfT+oV
apUfDUuk1UZqVswobGyfPv0w+dFyeGJD5yRU5PGFXRNB93i/68J0kwJHzka/Q0OJ
2TIzDDIfCTsGtDbo0s26L3t1pzFADCac87aZLn6ATq0LvHyspo0ClVZGewtVot0+
9/Gupald7fX+oupg21plt2tmsXVm+Pczgp9iOqqM0UnGM9A8fE6FAo6OCGlAOtiw
NRb4EFG2TatrPRTZDjCYkX7D1CL7u8hqMk7kHNrOdFdR/A+0pJMFNVB0c7G+7t4j
xgWjyjGQQkoFCH//1iAvQSFDDtXLqnBsBEkbfhRBQBp7RKRsw6cag8vSX87o8FWa
qv9+uV/6CrgDIxawivvBDhSOBr845xcEW4RL4mpTTDvaygrD4n3DJ6hca3/Xrkwb
FLzYOmG1EjzX4AI4VfQSYFEdhPTp1VVlbKkHNi8W0hkMrcTnplWkZlfq1LoYuNfS
YAQ15wSxtJFjXkmPJD7Nr0QDSncwJV94/tNq6cGZcp19c0RJ1sBIZT8xG5Sk2HIY
GzM5/ATxpeEA7dfO53EEWJvy+uQ3DGXFNAIkior4LUPURnd0h0u+bkmBvr58cncu
dYv1MhIwv4hBOlv7gqWf3Y2TtPXZmZ1bmkKUSo0R54PaZrYVRLagZxaAM3e/TwWu
holHzz6SrXL4iEhJ5paowAenqB1MxC1Y7iUJfTRua1HvMcmdXDpIUCoe5nQD6A3r
Eun/88W4htWQIIkidxHYCUclMmes5dYVNxJMQbc5iFjIIyhVdvQzUSt1CusDQw9e
5qiuEiGpuyoKEA76YsSQbVGYezFUb9M1937ktFYwpZaBfx/lcCXqxhLi59pghoQE
yQVcyJYB8SUCB22gW2/FpkWYWVfbFepzCr410amj5IOjffiSwq0mH6G3d5BwXvVh
s8CeNaQDMIUokWz4ljlBlgAIrlHHr7kfLrEdMlh4UCverg2bUh/NjhhmEfBd6Dzw
0UjwwwZOhHX9iaSvtsHI6BIWRHdp1EAUk9xClPQsnjc3BpcO8aXTyTYvqzXONYhO
aLnZaZEnJ5EA4kTegkWzWDyimQg78X0fi9aKFZdfUY8FcKPYSpefNX2azAzrIh7o
zzRZTEuZdzsWUHeFBcrb3Cht8SOP+RFRhU81bN8Dx4/qJQWzqUn8V+0DQVDyLZ6g
SaIe1WNMHrKFYgFs5Rl8Hw8anQ8ruKQx5j1ykHIyaEtN8v6wh52NvAhhhnRRR/AT
fZtSfuv/HXs2ALWsjeeWpMIV8TXB48eTgwYSOYwvGepfE4VfkxrOf7qd+4O8CBEN
3AMQhCcVUWJozLzPr+LOot+CNrJrSuO/QGEoznEEFg88I+yLeF6DopmDvYLU492t
ijyIFdWKzRZflMbkmHOEmzMt//9wUIy+lMcI4wXBWW6FLZOm+X25aEC8e+yBj3Nq
UZg0yJm1BVrpAt7Eggwq9tDi06GTMv11uQL8gYVrDw8c4dXl0Lfc5x5G/n0ET89R
ipaeFoHe+Tvxxfk4gH9YkQnW/zxi3cdwOXUZJpLCLyq84HMSpC4dmJ3yu4rVtubJ
ueUdS5OughIbG88hUZCwm7RAU/964lYgR2Se5B8pzmHhCgpLGSY0oUQg0xj033T5
9Vj9BQoEwuYhMbEIKYERvSrnorza8DlWAVN19BYsYXtm7b6ZEzSeZRkJaDogpGiH
G9pTyytNzYC4Lyz7M8oDP/Oh5Bg3eqttO2hN6qt/OxlsT/BAUpstlxCNR1Wjr/us
NXXWN6EOmAsO+qS9HJEp6smhy2Yt05TbaoMTq9HFqqiToF87HscDdFpnv3ORXQWA
8BZtp+RFSdwS5Al4e1lFXH67tfuo5sT5d7i+Eu38fy051fATTJ4lvOTIyQY4pdsl
V35jN+nPGgW+sIzojDLCqjB/CZFjmQgLfuUeyOFAvE4W+B4BaJdQBiixxUXwdlai
yjhRyUnEDdwwQXzGir4QSfXO1Hx494+r9hYmh8PgOBOiF0nTb2UnXhhiJW3pbZS2
wzuQmpzgY+PkZg8UcN8RP7mlO8KWp6GnmRYiSVrT0JV+a+gKCUbR/koooYiWG5mV
9Nxyiw8sTi17OzXYYS8go9O3ADlK0l/vrNCE7QDpqVg9ynsBlm/PJYvJZepr29jc
2Rm4vvbI7IUBJquFRXZmmO46GzDSzJUgK3v1OIInru/8OJ2YglDntqmrRutrs2Ve
Itt2E/9RT7HBATnCk6BLJJqUxxfeJqyT5PFbY0pczPRc4vDtSzHG76YKcwfgornV
H4GOtWPgycl9+2tJmakYag==
`protect end_protected