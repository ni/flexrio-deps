`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 17440 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JXz1+zHgF4n2s6TEZD4KtuQ
ATkS0e5WlIVeyjNZ91Ns322acCQDUgeDerq6TAJNtXFCocksKdi5WDPoEC8S9T1Z
GV4lMy4PWCYb9y6z3Crf1rXX2irdN64c7cds2jqtyiyNU4B71W5gKlPpQ+zK1nfJ
UAsZKhduPAslKvKO/1a7sC6Y+rc0iyRmh1rQNGqos82XFWTM/BDjlxA7fd6pXUpZ
p8qJp9ci6YmVqrKA0zbFWsN4FFxtrnrj2aTgcmN+rNKSYvEfDEa8GeNw9H+Q8avD
uB5gIm+yJoWmm7LCGVkC2i7IBUekoyA5Lp249CnVVdKkq6kGnAUXEDqLiBtB1zEW
jgij3r4d4ifLhH1w3khFyn47j3sXvnCCMnnYDb8r4XVP5lzNLrCCl2PrkyfXaIU0
FYx5vfaHvS3SKcmc0wyV45IKwrAcf0FRPV4H//S/CD50bl2P2SLBHt9NxKxzGGqc
oMo2DllkPlQCYlNPf7Y7uEklSv5CUilHEloUTx4aXyq0hH/tdXfGy7QDwSQEOsc7
bPwv/7geGG2cHU26tpa6vT/glwvk3FFkeVWTD1DUwex/H38qmF1C50DzpeNrvSt+
O3ewwuLTBLaLnDKVbet9CVepjFA9s91/mg9Z6UJejMzut1CdJkfGAqy09n8BUi08
RL/py4ej6Ic0labWg9OfwDhTmmy1dhgLt7ZQJqp4kCgqmCVd6SAnmQflWYaP/AxR
NPIRnT9Ww/aSgDXMSHqxIEfGoFzFolBEvlJlwDaS8QT6k7zitSO+dH++CEl5BicO
B8aX638SDdYU+iEMhq092KzKZqJLveKmhn/ooKYVbfEZ2RNCCqh4g6U4ZA05UDWM
v+YRI8MMebpg1U/VeJPpZtAfmV0pvAlvTj+yjFrDuM5NexaYfuNvqnYaiR/6TIWn
5zKtsAftgGv18Wt9ErwCS654jsEA/+k7X6/yE86bn2coJT/IfZhu8sorKbG38O0Z
Rei282U0MiFOlDa9Ao23HrkFGo3mev1Z55ks6HmtlwmwH6AgQBqj3ZJoU44MpQqH
YHi1SPX5PERPXZCUuHJkpNkCv2rjGOYSHixTbEVjAOCr+xOMkyNDySdkA4gxMyO5
/KUHfG7qGA81C+y7zwSbW2d6RmhqFSuvIWvB3yedDDt6j8PmO0mY4yKGO4JBjpC7
l6+ZgSCY9/m2WbeTyMcc3zm7r7um1zyCMofwlQnxspMnWxSOKP1utGFE9ScqsbdS
zdpIFLO4phcaNJJjJkUnZ2AhbNNIDxa5ORkR6iW58Oth7GeBv3B5CdMFA9lg//bt
eGIfJySqUWGSjgn8gqiG364X6REkBQzga3jJgAklhTZuwovfaAg2sBJgxqOBRhQp
hIXIiBcS07frOa4bnSFuPA7La4/v37MB+wbLjk/2vT/S+3BNuoYgE573Nt4rFe3I
Dz7FeJ+poRqH9Yqzsl6L2LiyiSn3E92tVtT/J6T7tybLFPjUMVqTZe7yqS8raSLJ
gorLFHMqwQRk1FiiQGRwLFdG7OUIAVOvRaefvttgMszVgOKtPvdJuOgeex4caU7g
AoE1MOjJyY5lcURpr5XZmg+2uEXICiIPHaVg7HRaEkhgpirbeIB80SOLzFCTJyt+
+y+fgrEy/XxdL1ZORkfvJpiZ/rgTLZStiEggOewy8S70cs2t1Hv2+Rs8ncVbgJvm
O32R9bVEVzCk1Pviad9OGh4FmUQa37Y9xbrPrC6qzaxlDqzxbVclWYsmegjdqT+h
B/6JnVP9UITw+3YvWy47Y3JS1CgQO0OyDrsRcAW4RLcUvAmPySYOQ/8S4cWeMi4Q
gA55Iwb94PmQ7HrV9C7dJ9wUjtkpG3n9EFEDRMNQlcdbM0QXxrQZmAu5pqaf7/D2
pXwtAktNpbP4IvSvyA7txhyD9R9U8KUIWVVha0Eq5abwrFDiFHK/jmxEHdd1oJJ1
kwvu0UgZf2XEl3eKlWsO52E0mSDL1joUGo+HgU74avhQpqYDxp7ZvBJHxS/jCDeg
dqZ2Xgj+dFpkkDKwKS4g+ssq3CVTTkMaQVr/ZH+TFFjWerDNDpJ/GyHYb1LCmKom
Dj6ibVci8UTwkvIBk4mgs2b5qbTFg8JxYfLYdBBgdchsv6IIWPXPZuvJjPpn8u21
CT/dMnc8cmQruk5TORJwtmi/kscAthmggbgHTM2tNZ70LWFJmQ3R73GVx/S3u+AZ
uB6uzMzZ586cnkfhXmDe1EQ7U+3zvBO55tUnRCNRkHdadbClsmfMxCNtPE1Vo1J6
hCzfWf+t+eiudCrd/NMfZVHXBOw0qj/zSMvCVNuJrTUgt7H3Sp4HhclQx1xSeWP7
n2RwOSLnSMajRb2wVC4vMzxENNS1KDjvCWQm6b3C3utp3+CDHEDZM91C9WFVIIwu
pfkU9HTchbFhMcMW7ESAaOF0lRs+0cynZ3bxG+iJEuu6OaM9g3TFh8N+tBQKBUtc
zSejnx1bGd0sUadTPkaUrCncjTB8qQ8ijqkrXiLH2a924LqHFcmJvNJmT8lRF6Qc
g8Afu49ZexFv+gU8onEaviFpkUartLs2w8AkJpf+n1MCjJfB+xbu8SPgSXEAiVoq
GezdgJYIUxPw8U1qz6mwltltJZwimfQb4Nmcz9LEkWAQkO04DXYEeQgxWBqmGp/S
eQcejZK/KZo7w0o3KWjgBGZllnAyDv2twq72EcM9sHIz4Pk96z4kGip8jlmsKDK9
jc0pQHF5IXgH2EOI6zHIcGOesO+iRT4IZ/I8fuwcbniHA3PihV1cpTqZy4WTVCpi
7F8fI8aI0VQhCB1zfW1+UWMGsuo6cetHLSyGP8eXES1Je5C2PLxjVy8MNYkDeB2p
b5+GhFxi56Z50nwzvgpsTyLK1rvjwCYkTNBtXeFjcfeaLV6OVkLKHfW9dEg16fz3
yO4Xkp98Lsf9fXapN1+w9PzeXD51851q47utNh1iT+3748HnmwWX656PNREZG227
4G6Nr54hF1MuQB4yi0Kk2SNot+ThJefhVaemcHS7r5zcG0omnRZTlY/U1V4hIt3l
LhPdIaLccC9hNxeRnh1CYb34u9/qF0f5oyIzWQ7oy6WX6Q1m2rzhDLW3wo4olOLj
0Fzos5D7UssAAQkbuxPKY1ItOIkmYMp+BadWwXs/Zn6/VGdpmJwIu/jSm44FFCss
IGyF6z1lVKqulcnxmuF7tIRBuLc/6b52Br39sRaLVIetJrfT3a9ZWEtCcI7vZWr5
a5D5hb4ZJxXOam9K6WHElGP5pE40/v17iTCB3S8VpUPvP+AbFFlg/kh36T3VuZRr
hVP5owUUN1f8PK4RYD4tUFmZTPpmHNGLzOGNz9RXpui3PJJ4YT6S8FgKt/nBQT+w
V+uDDwACdbYe2Xx/Lb/AFrduCWOiypZB1CYzRAoKtQEjMu7dL84yBXYgaJG6SrKL
jJepotSH2u1eGabao4IhhGoec2drHqhlJZRq+/uchAZvD+S8YQXIT0y8NlkRAN0o
Mr4prlLjN9BU1+13YxGRAD1WvTLXjDv6CbVM3/Vpcv66fNzojKtADIyb4gyb70uy
LB/ijbCqrfqdbeiUd4pSqGVKNLuDpCGacatu89nAF35T24wiJxb1eVKA75QwIv6q
tpClvwcOR3rIF76X2lu/KBDQdEvKA4lbOf2z+5kBDPcpPAaGlooVFu45whS9YSyY
X1LirtT/RasaYG7ZHfZdgByGvN+QcsYTgxW7Ju4237aA7bzELPRVIwTyt2AVM98x
iXGpLYHbOLDw6KoD7AJ9PneGnZyZgQ8FOEIDo3WBmiAclZyj3dSs3iktS5PsKQgq
YyMdoPlRmZjtadPa+OxTabv79z0xp+ixxqh8YeLw0FfgcAIGsRbJIItAie0qPAQr
iNwroNoV+SZ5WOlXCVI6Sl1uMOVHUQf1mOsEosKH0mWwSKMXCMQS9fuZ2jw4JFk8
w/hgnLnTTc+GdBsNj4KUxiI36elGc7SiAGz/P8iZZiz2nldFX2fNVCGDOgbbD7En
Q8o+DigQGMU3kurcJ+NwuL2uZWgZyOfeEU7BhuEL0JuEDfSYU6YOazDv6EoObwny
LDeux9GczUEahUyOomcnreRk1bk5rSVvnpY4VYaiFiRw2BD0chESmnZiHQDTiF2Z
uPZxRgt/kQdrtIBNR5Jds4BwtOAiQSKaP7zxuot53PjgEnc0iM8pxN9BjwbUjtg+
hDrXGYHybvOW7PUx/PeowXcpECYUJantKC664sk0+Is4U+IwDUzW7NRZP3T+3qPy
ESiNpJGjDGR3L/7fyZMqI4GT6coheScDsfBf/KVZuLxo7wIdVEfJ6HW6pyUSp7fS
ykoyaG0fiti2NWmefdLgBd6zwcjGOFgjZHB58mZNgkKFOlr6PGEQ4KhI4p2PtbvF
QXldUppYrf+dQoQyva+jxjvf/XKwWxt6VJrS5L2d6aSJReLbR2LQIlFc+UL95xhB
QKjpdNt13+VeeqnrUxGDTTBYrfELBL95MmpvEw4EOF2JqYuWmD9G3gXd/CS75Kz/
rbamDg7Bl257tCFMzYkxv992mW0Va3/csDqmy9PFZeKUwD/DkPw04MRf4VodKB6Z
y386if009mU3sdqI4JEIyKFyRrOB2cZmp6JWjQxOzlgWsJxirgDLXVChTuaO0VCx
Pr9z+DjqxMx3eiWjCuSaEUzbNzrLJ1pZrsN7ubkfq7oR+4HmpH1lhHO1XikKFvR6
2Fz1XZ62hCdODlyAQoe/vtG4uXFtS9/H5RI/wr5/ODTMvzuB4O38ou5cwygvJBPh
fo5sOp0WKZwh1OhVO8YClpxr5IFxyvlhn/VEDEln6mf5oSc7lSwRmSPYUYpaEI07
ye/6459idd1win897UbCEopofIJs0lEi2+AK9mlIPgno6RfcomItWZcgJEBDUJDP
VL5OkyodbYqOhcSoVD1vvTHm7KnN13JioYRxOrGNcjeuhRyHaR4C0sUi9PTuQGaH
0ROamQskSgpXHcRLmhctD2OLJXGsrMpdGk5jeTqshW+kdKCdeCdJK9zeCy4d8myY
YMaQ2x4tkv6Ih8vIcvqDWmvt1oqKqjrLBv/st0FfjsV3CP8qVe6uzYYHBkGkKK07
6Tb979xHiYIHfQuhpPQtO7BUmVT2ZaEf91GMJGeNhYpUBdhzAhx6qfLLgAznJnGU
t37IxeWyKt1gZgnJufQui+Pm1OGStgfhaDjYcKMSu56dznNKoi4OM9YOwUAc6BPb
avh+X7pF5WrXSzOubWAdQrV4upBA61EgFv+2W1cs8lLddwphCLu0ogH6J7naBeKY
Yhdbsc9TsshAXEs29TH9CEucj6/HnN4zkp4D8C5UN6ExvMH+Aftb/Ehg7AO1Ki3H
sXpFuoFCDZQjEnFV/P9pym4BRaPq/V7l6OmpDa6Dkf6pNPsjfM1VHvSYyXSWTqJH
4VeAdq0DFSs1bgAZ3DDcf/+IPdZP0K7Oc766OLl6K1i4bptYYrWWXdXgpBqvl5ur
uXlCv94rIGCp7mdkB+BB3eP25NLrYonBofr0ApRNKXj0UY/1txuaqAh8H8/OMNUz
jcWN9sxP234mclb54D5jcS1DePJjtYCuij8OH3rBWJ8O05ch2AagZ+fAzdAm0Frk
PLDd3XOLmO3/NK3Gz6rIOByD2CRi6+/5eDp0COh+XD6GodBZSRN7Mh28KOYEzmx9
7PVfvWaWwS0Cp9Uijc+d7G2s7Lo/eUJhWyJeffUGy4cuR2NZTyhUMCeYnPjuqm9g
M7H1Wwu19RAmWgX3Vp6s0FutcgjTS0NnRIXVGT7ZuL66PWScrovK2FDCp4RrixlX
e9XXKkpGyBJe89ZUYAmQWPSo1rWxGS0qXprNZyDSfLBzGb/jTFMPOuMju0wZe09M
wuBMN7i0ZBiPyq8cjxDAiD+rlgpSTQDDmIxUyEIeLMn5O+nHLiVq9zY3VLXZ/MTp
FYcJqw/pYaDcaK+VKWEjJ9iChxWDCVDIsOWpll2+h8LBEVgbeLIBvT6sMrYR0SyT
k2rwd0ghs1/h2jm3nSgRENxwDVnjhZ4la4NzEdxF2VRTu1qGayAGFM3M1haHx7sg
4zD6TQQW4OtfsDfUsHIfPeXiOiv9AYg9rKUsCCS4lR/oPJTbaQ1scdxEAbjYytfL
HSMOjUonAcMwBpLL91pqNqn6G4fOA/aKuMkrrp76cTTQuFdyBxO0TEsEDobpD9pm
uknzaUHgKJbbvb33ZfMfeYrmDfx0e0xq1miWdaOjjiVzHFZU1dRjz3WomWt1p4fZ
ILfbNRESI8+tPTfffeZpwGaVXq7iJH+hX1K5kWNPC90Aj7uCyGcZQV/M7C+/JaKl
hzyQNARkhppHixqYxihHTbtYbRvwhP8edAIivjROfRMdobaIu2EJq8cHAJbp0ce7
tmnArKuw/WbwB9XC/aa49JQ0ES7SYJp5oj2nKlQwifPFGl3XIeWzpVYaIyAfymyT
0qVItCuOofqduMYR45zX4hhPVXHqJODw562NyQyaj+e1WSYALq3iRd1ihy3YWwNs
/DxSQoNErMwv9jE1fwPqWJuwCoVIwUbcYAm/V9U4ke70BFiWvp+xbFmZP1diTWf0
ik/lkUHuoxVHt+5ogyVHsBVfBgUslIEEuockh+wGOnfH5wlPSEe8I6gihYA1tagy
MKApsNYuORWncRCzPgEnCXYXZf3SUJO7amN5s8OmAlXM+FHXCbR4fAHm30c1wTAQ
tXnnP7mbEvBUAsNiz8vpoCmuZn2PJZGkPmguL7XYmhYnFN8y8GFgLD9a4A3UEipm
9vwSLxTQRG49AAI/rPcKfSb4/C5bNA0dx/iWQq6AshuzUKP+MG2OdrwpsibnfbbE
nzGu1U1wAT1ohRu+6EjswmsIKQ7dQVuzVrdqp5JYsHMmGZeBL27Vgv/YRORdTg7b
gcpzLxpp+SfirnN3uj6plnNlzfyS33B755NIlCUaFky5mQZLhC8vfPBFbhIjEixd
/Sam5w9ZY5ecSuW1as0iGN4PlpDCNlsofK1vNEuRXYcvFnMNLh8zTkmRT/vJLyiP
m+dttHxLW3VqQHtaOIxEZ1SETifognXK+Z0lzEA3MVqtsFXxg17kpATFjFExbKZ1
o9DpVdvIa/1ZBqlo14MWJvay+YpGYFtw2dcPG6kD4r6gOKi5xz9wU1lIcPlcXuMI
yZvvD17WS/41gD+n66N06dFZamvrB9ShIQDuj3qo2T7NXuIlmEQlXJyG/4Aw5wrm
HHimqC4jqdweHPobt5ptiFbIDLVXsdjy81Z0tcnOslaq+B+O1ffUDkdglBFTUthH
tHyBCcRpM6TBDwoetH0brhbmdj+XT2BrB0wtd9r0yy9Q5fapxbyO9jEV03PkegNT
as0W6Vq6QtoPCaSWBKEQCTUdXR2xbZ6PFjdB/69Z/GK5ah2Q6kglzM6kzznPaD89
A4bqxzulXsnEBkhfHs5P6k5hMabnOOsMDdxjURw3nMcJZsCIx7CSE9LAvmzA2LAT
CRwqeDK7J2beOFCFndUz+FRXLdllm04ozd82IQHk34j6TuVk9kuCEmK9d3Hr03xZ
MXypo/dU1XysDtKaDEpc6GXWg+z5M5asBBIRTc8dqJ75zGkil+JxGuLhPiKkO29B
MBKH5Bboen1H2juy7WlZ4HMuedpPDt0b1lsX+JwIdAHZqWMsRdEsQNQ8GbAnTxUs
aUaqTvQF2jF5qhmHbezZ/rN9ZCVlHiD/AkrFswq7KEtayQ9/jZTDEul6oJoqqqNU
+q9AGfRaf2pXLLG2NFHOZj+wZDORL8V0GUIwmdGTaW0rDFOEypuFhJGOWWUZwrlp
p10k9DoiOqR0eLMdPWf6cvl6yjn9GhwYFoA/n5MNy5lVRBZ4cuJqBQedY7zOyCQ6
aTdrcyaWkiJKcBpzvcTydfI4Imk5yhlFAwALqwDmA4//hJgzKPHwa1zhqbFYbxS/
pwX6VcEdd6jdmNIWCLLnpXEAlC12Nh6PKsTu/15QiiNRaGaQFvY2eruhf6+R4Civ
WO528iQ0dzKB/BpD0PEoBF4Cy9KW5ZCDHuqlU0qDiEJn0/TNzj2/2GyQ0970cgl3
XPagJERkwEgDpfyIMnMxyYZhjmZkgJG8G93NhLMlKBjaCebBYRaOFDWqWoIpTF99
Sqjdn5c98ZF0Ok++M26B0xs3FXV32AcAYHt9SL8VNkoEdXhxXC3MbXmX/LmX7bii
TVp6PwlSxh8/5o9K0P0RMK6Pc1pt/GokdwS3R5lCxmVF2rHAW8yHzdhnsiDKe+KS
8t6K2U1rohk7BOznlG7Fbc4X3oW2mP48u5QxR0DOiQ8hWuuTtJhGzqNW+tlzbu99
pf2d/cPMVrAwtaKq2Joxp/o2h0jT/2qa1GFsT9TRQ/A+FkBfKz32awXdGj5Mj9vR
JBa5dDwDVh4+RT+sUqTCB1n2vydf/0ujC5jdbJsti1JJIfycnUpIT+01bj9Uvne+
nRBcOD/zwxWlgXffnWa+F+4ceAAHXCGKzI52QIcqWkOrcfy2lfEnSsRsjy0e+FrZ
+1ffFAo7eevkOn3nqGGUeStiB2HijvVTcYkvDjqxEYIppD3hm6GTPClCTWJFs/h8
MCSKIYFTkU12MzzhHwyZDz7wu0360yL9AZhXEXZdCo+ErXJSuk/86CrUV5XMNwvo
Tfg1rFexVhmOR0BgF3IMHTJhvLzjKRiFS10TDxaNYKBjuaHeAZreswXDh+zwmKrb
l1aSkooEZ9MIhrUfIjpjWoj2GHVcPWS/kUFoOe3vpr8B2KZW6Yr6ghbF1zI1QUxq
yJUEa/Exq54tIPKk0tguJOEMAa1amgJVAJFrNUcUtTx1ZOA25khszTq2Wuc/5GDc
1lNTHWqqLJSpxG49IVzlhaFlPgZ2oTHepjNBlkHukyzSEtefpWUMGfIljOsNsE4b
L+0vnZnaDR7De6+uAqxzoEOVqrnDNJt261PH0jcTeggvwNi4Swec5YJB3AwgP6K0
LwqrDgvUPdCABWqu4hLLJrB+pbtmrnBtQ3APYeH1x043ksE8Phb48BeR7HXRyqGs
pAJ5bmHC+918ey8QnvjQUNGfHWKZMDy5ujMD9JBGnBy218nYGQDWBkRlKJ+P48gO
kN9pMplzsJuIGbLBa2z/htpDUh9HUtcgNS/l1Z5A7Aw0Ft5WXvBkq+SRy6heCIDj
qnsffHAnJWvEmwPtOdu4IqHCOh7Ai8FTlS8k7p0V9Av6fJAdviuj9HthZHopX2Re
TS5XxexsPum6NOnaomXivBaKopuV5cVFEuhXoY3uzf/w5uKOpGk4kHq93z2C45w8
422P90NoDz/C3LqsP1dPpajOmqU61uQWtS2hpn8FLcGLZ365LkYHeKIn3cEhY+iA
ia6TXgaYwBGFaV4gMgdMQ5IpwEaPWbqo+KUsl6K2GFwybotz24BoN1K8I8ptQiKU
/NL/RH/h67ofwidvHFDGVr+KwCdgvLH979SCZyEHa6+nHEnzSCFhzU6gCdlZHEd5
1hO8AWKNpxrKcCh+LjRBdrxKEnXxUfLMUx5g8fG6QtLSPgJ+kHp9s5B9S/FMwOkq
fY2TA87qQqduKA4m19VuWd+ROo/jiAHlV7lplMjq/aynwPKF7P/Uh5gHI8/TMJ6I
YIcjjGjOhaNUHmD6adkQ6masV2I4xDfycvcCkG9zywZwyL0Cvb7BYt1O6xB4Hzds
pRqYb9WwGNCSQFPl34OJa366RhC1VKwE3ekegiM1WyeT74V5ezKisWNeohN3o0za
arvmYCsjsmQdPNXbYC3k04ZmdZ/Ur0mThea7FLHXENC6qNf5rZPdKLoYSjhOmtOx
P1XIvzeJ3X5XfjLFO+SflmRyJNnh4H+FKJxm/c7i2nBIGxo1Pn7+mrjLvzGZbh6Q
bxa4rvE3G80b/PvpTadZ1o4X6DmyL5gdkQr1iEQpHFchHLH8RWuVJp1npgO2bn/v
WQiprFWKlkvAIuHapDD2RsDU2x8nXfNuWSzKhYTV8El1waeT+xI0pYeGdMK3dGQW
kNbzUoYXaocaH2Sn9WvjpK7DA939selOoCwn/cUYb746QnqRQe0d6vA3P6Y5AcU4
gIb+N7WzC03pZ8qAvoLOFJM3donYFSb0caCUJHqYqR6eYUKyE/Ky0tLXDKNkozPO
UfgbRJ+43/HNztIPOFDdoRjJBrPbLa6npP+TfgU0J/N2I28TlFi+EJJ2lmv6PLhf
Qp+stCdo5tsqp8B000mzUbhTXq6Vp8T1BrIcvjS8e+ZKo8gfZTF/L4VoNnrCjV0K
0JNDxDqh9KRxinrJcLE4JEhETwGa2BlsjqXPWAGZPQYZ70fmM/ufu/RTQyx3iaN5
Z5mMWml8hsrAw5gRvPu5RF2BgwzuPVOeff+w6tjzDX0hH5Hb4Qj62/u7vZiMmGov
2qPzs0mIcTqdqnhnVxzN4XfINibyA2OXSw7DVh5alzPakVLRTd5eA7/YNUlxQLmF
+aQivX2fsbQugJ7CCcyfZSAp0cnnyGFYC69Q7TLP5U5VLrHgoBQV4wbYYGHBg2AX
ELW+/IeB35XMb40PZtgG8Og+5EM5D55yT+Ir1Edv3HUzGSZJsjDG/KonY4eJFz0M
wzBtwrHC6phRiNIZkDXHdrMyqn5lAVczjYXT3AI9T/MVFK2mW3YikYS4utUoyM9e
aLytvXj6ui02l1GQ5S+TDXCHZAXM8l7uvuYajUqlL7IL31F5UkSuVOU88/G6fQVY
OMT5/obILVGnkS1t4FmO0zIrJgJFHGHh7CHT9H9ft1+ZyIYKBhQuw2/x3gdlvo/J
mKsPJFrZ271vc9c7wbzG1j2/PFriySAVTFPBHsGJhHhl00cSjS7vGWA8JRkP9vn8
ONSneYShc+P/4V+BY3uoN4ZIX4gbtneAEevYNC15X+RrDMI6FkyYIV7MBPKwporj
Atr9to8fykPbwNsU1Aa+cesmJnSKpNSmJQB2+G0URQDhU9iF90iwcSUwckzKuJ18
juCApFHgrUgRm9G+UU69Ic2ZmeDwbe0AXmr1dH7Xn0INWkBW6SCxjc5FpWrOILFG
L8/z1FW26x9L/FYLImjkE87O8lgo5ZPFUnpQhu7k4sLzs125zajilp3uiv6pc0Pd
BRjRSnl6IaruCgnPV1kyoCpk7P3WzrO2wT2s9pdHqrPNvIbWm5RlHClLlDIhGQD8
ngGdJq/T8rmzjrNI7iOC64G4XYatzLUtYJGTN+SiYWb0yJnLXzsw2gmWVKlx2a+N
L0ashCooZswEZiA3FLAvH2kR0FdbwQ8r+oJtbnEalQqRUJkSJMRn2+eidvAljL5g
R9NLR7Ve5b66hV0zB0MxdVfltc6VT0M5Qk7zKM+6ArpAwGzoZhz+xjq6XfEpji0F
DgTnZkN8SSCtqVUSXx+R8z0CG9tnMDl9CWgZs27tPA86ydaWbF4ijfLdNGdcqlVK
vveBjLXL8FGZUHeWAtgrd/BfgwSx1P1WdNt6yVQ8HM/RmyzMukRy2NipmeKgzKm7
ZHtNgFFY4PgFcTJWEY87cacCx5z8mwTCQ4o2Bnn0AHqowPVhSq6C2W9YGnmXesS7
cZWIEOKILmG3ToHe5WYwmHBvpOzhViyWKFJ0HAu3ng9s+9Y7TY5FJD0xWnomxrjw
BWR/VjAAH/0pQTGdKq3Ma0RDBJsFjI54mkRbSqmNHDN4rFDg+dWd7ZntOYMKeazH
enI1kv8xv9i3AFYe8RMVCI3JzdRXFm2npEaxmgaJHLcElI8lib1CXQS419uwQnaR
O5mXdZzpH3cVRfuqm5k7trEFcVVtxddND2fgCxC513392/A6ALO/6jQkdzXOFxbZ
P0wDAMo1WCJ1qxFpzudrscOkLjO72qutKEET4BD6NkuiCo36n6iOf91ieVQSHNpd
aHUJKHqN45KYusJRTOYB9cCUVkHI08dpe6j+MFMh4U59udTQMEqRKepOazwjVORO
hSb01y5RJH5T4fGBKWkeAKbVAIWpgA3lj/XczkJgIdmLfGZzjGLwc3HBTPgUVTW8
pLG09vTLDy6ZQMuJPosNnGNrt8np5TjkzIoJcAC8GLHCtooMv9MRBIeQRPtJWTYF
0v+blBcuPBR4KkVemC1Hd3tV0i3vYHEu749WAGnaWrrPgqNa3I+W6B+ZZsvq7Vgf
GzITUSYzMgq+Yp+/vw484SbDOt+okcEYpXoJ4+MOnNEm7fmvVXH1ymbMAJBmB6uM
FI7Qvpg3lqSQ035RjuzmbqFZ5vnZqFnrCRKvjAnk0Jo6paFbnGQiffuMgXBs+n66
n9QMdUcWjYXFaiazzZJorHiK53t0kbEshnWond5LqXHttYTEPZYhaLebe+jO4vEV
zEG6GgCx3tCe3+g7/xuktLjluSAdiv+uSDehfC9ffdGx9uhAUiWAIQbUPWlAC5p7
AZJCQPzrs+Vf/0RNM69Aq+qVY50+AJKuU2p/Qdzx4JG1H0tkB+VYODfVm1InXHc7
nbPazXffVMk1uow/WqLqJjCOZpYfo16+u6D3vJqe0JjQJ8lWB3M2Lq+11zfGa7gZ
EPfGsix90x64B5INhFfsYojywfKtCIAVXiDC8JxhmH53zumUovGT6D3f/yekFkcB
TUQ1tOBQ3QM8uVwnOsTbGDiq9Il20wGuVONxqXDtfLA0ketQY0AdfkfwK1Ju2Vg2
yOaktg/jP0CEILohxrVuR+I5jbRu92XuLB4nV3E+t73t7eMkiXIVWl5/BccEbWM6
w6iw7vIJ6ov74K6P1MsibQczJo1GGyJM9+p1wBFwL038ohheTAfjCcpgmzjtVZhB
GJe0ZN391K392AxZeLFfImkipECz1KkgxfemIqiU6CURFx48XIdxliNd/6DJJ2RU
p1P4UqworhozfZz/QjJ7N0Y+ZY9socEOUzeW2S0vRkZhhim2athaNX7LiOTavBui
u90QT7w0skLOe37jWXX/Ie9Ic61PttvGy4gpmIAswQ+HKJXPdkvdETZvOlnk83AQ
08lHlaXCTkG2BveElTV3uGdnPWZ8TLXullaM0K+6/oruVtAxQDjBUC5FMnlm8TLE
lyin5qhmDwNSQIPAjY3FG1sBcGPkCAAwuSvXJBMIvFBfV7bOpYpxAtb4c8qwZz+Z
2Zjv8XLEh9H94vpLaUmULkYv2ruTopgaGSWOJQuTJfiIJatbRamb28hckYklMTl/
qHzmXlBbEd5OypzIP5ijgxazTe9iQm903W3ZA8wBWqxQ/8UKKbLLqEERIolRBk3r
AD37r7aw6cKtnM0Bw1iKbTfLuY4H3ydXSyvq2v5DJZel/h7B/lkVoEJMqytl1VkU
u3ls3ZQwOHjUKQ5uKqyL7zSiVnV9pmDfQETSvLBpQVXC57WzygvAkgKdi5ODiM5b
9CdUvyHLceLsVA5+CmgUCOhwoMPwDTwOyRhZ6SneMIXy0hINisP1y3SBZ7NHPCqL
1+C9shJEWTSz1yfByNtNKwISTjmhmk8k2GyveZES7i5j/0bUY2HLeZxdWFWqpDwg
TdDgj8QWhsOC2rmWXZYUFWE59k8QRUKUfw02zdUWg7+R+2P8AzOJu92GHyp4HFhK
Te4geQK7E9zt22Ze1n1TNirPPWVtAZZlHG0chxz5P1BUu5rdk9VxuW/jz8y8hYWj
ZppUNgALQwqJXnUjvur+jPdbqCPARM7JNnj81pmpI7eYWjmzdnK8awtktPSgcjca
usrkJPZzKvKoMQcyMLl4Xuj8xdqFubkMquYPG7QcysrhDfX2d9kYywZldM4+2Jv5
b48h9wxavMQZd+S7ccrEQQNU2cwh8K3aWCGgDtSy5T/Rv6lxYm3ITcKneGGDmPzw
kKeiVJz363nYbuTRHE/2P20v6zW0VmTpN4IAXt1CYxcHsVMy8DV12E/ZJfKi5VuO
6fVwE5WbLt+NARXVTGbK/Fbs7HRl5V/C1gig+gKAnaI4K+rKvXt6d0SY+r1E+jSy
E2BeSAFNgEfpxGgHwWDjh3l2dH/ROn8RPCGiaf44yjuCyuxu0slwQ07k3NwQ0CyQ
pxW98uPRFlDrMEAJBY3lvpLNa7MmnFOtL01ZU0ENyN+2TrN72k3kXD4N4Rx6nJcz
dqZY+rE8Xlip8MTQM2p0x3jkd0u9Ro4lFqUfO8IbzfsMihz2nwb9x1Ri0iXmtRfE
aJSKIO6Q2x2ewc8b6yhvgg9M/bIOgkSFiEhZU9kyRjyx3bpaFzreTZLoL4B9w3AQ
QDo8gmI31to/x+AsrpWnWOR6wE/ltrsXRLvqtPhmRdMhA9GQWDHahAYKgR2596/a
RDlo6RFIPKsyDz6op4HKltomdiBV2unuKIilM6PbV5Uj8c3cGN/9z2OChBzN4lum
CDklSwqspj6DqA5EvJcptE+0BLoO3oBl87B1pdaULuc0rjI8r/0N0IE4ByIbPIOB
zOuhkOKc1qFyvmavC7gkjaQcxZBqdloDe1e5wqIri6nfjAg6yNABBEc1QHvDh7c0
/RigF5BwUZRdjo7W8eugRXJGWmn8QqP79lBfDX/gXybW86T2Em2TVSW9DhOUy75j
9uUS3ai64QXZ91/ra3pFBLM7mCo8Jmh1fdTvATqgt5rfZLkk73K6DRwgVRJ4IxU6
TV6o/fjYjxd8130H01NDQ5TVLM/yLPtqWUxDih3fpHNH6JtmiSLrwqdqq01ebgWt
sIV4+dVEbfu8sORWzdBxbl4fcPchRcKzLBJJxCEO9p9nKMa3OySWaqXdODP0ygpW
22hkG4m66BajN+IFVJt1nFSIMWr2TSYO7viyU0P4cfSPW7c4PsbnNpz3EvbPYYyW
M445WHJAjZMsWqlN6G/zZ/F8meFQpXPaz/MDMCJq/rkI4JaMYTQ9+kfRzBFHqSv9
1Fl3sUgr9ZCYXkVZn1G3hh9TVcRN8liFWwYR9C3k/EWNU73+h6ZRhkhoJUgZ7WQ9
wUaxu9kB9s0nYivD00vk0/QDAt2PCVq4jBSKKPRrluv/bhH6b46RyxEYCA61tXhn
A9PDB3yuiZ+nRTlpNqUqnUwzb1jAgAWpfiq2hISPKssf17WyFNf7VjO8reMHV0SE
1zLoHCQ1qL+UQI5IzyBbbwCt4fVTcpy0QMtPO80wwGqw11NIUN1haUbLn3ldMurD
R39SYubf18Nrt2OOoroYqLSEfnL++c55RYwU4luErZ+scqEVFqFDFdn4bJHEJ+9b
BObG/VFGTMXov/lSeouRJ6g6qT33TD5cSg1O/Dsa21vIcr2V1N5tesd3X0cp0H9t
eLEuBAzCRTGwdxibRypS+X123Bq+xozcCq23RvvG6IcFvY6tRd1W2hQ0yXcJFGnT
RMM1Rp0PeVJmfRkHQ4VyFVbQ7akRuMsc7uh6yIZNinqGjOp4bQwE0i5Ka76192Qe
fVG58MuwTFNwdVVIycqUsA/f6UUk+PXvi3ww+XM/aAOcdqsy2PX7bKNXAy+Eq9fu
BW/7GvaDuY2Kar4mqPMsPb0QrRxV/RrD0/p+09ES6UDC94F5DQx8bcAFGC2rbbPG
hSvCcj2kmH0+InHHFfa+FqllzuNL+HMqU18lQuzV09KvITKl1p1XoX2lN159M2bW
6GDeegW4lEQeYeYROGRCy/aai9WMEgPLdTMtaYtbJT1rgL0kvtspehNIz/Ni1f5A
KSt8UTKLk4tR32kjlRGAiXzbCsvfbtVLut+8tdLuBg45f4sr/2dRUw7e/QTt+l3Q
GDiL/R1clGPEFsqjkHoBLX3KUGDBzGNqBZ5wqe8qrezIqSeAagPvPF8Ws9gfwrFU
VNl7/N40LkRh/3yFtBEXXF0jzVQ8iESC4VvBA+ajR+LDO9BhTsv7+3AV1DKyqNs8
9z3QRB9dZMFVMEL39WxNpISzhZ4395Bzdmsj8GEVL2KmEDjqpE6ev1LPr58B1zi/
+Un3cjxo3JPZjDtkqWIQIh2oca7ENNcKmZD+ii0lzk4gE60SEXD+PgxXcXHHcxNS
flUBxYLPvdyfj/PFSvPnyB0LJmc7z3fwgbebJ1SrnE721lr5BZ7dGn6oviduWkwr
Ks07fKhHqJ7512CrbSIGVz7e7xkM3aMZVbW5cBM/AkXIN18kXMKHDLoAU8/DoZ1j
BZnbZoUzIjUSmNaaasRLd+aXKhfyy5uQwOl4WTE5hyc4RoMb3O8vBLKhKvK08HW0
mKbyMBBXBXWwTVhEBAD0DCq78ZnGiS+B5vSznnDmc9+w8MfJIJk58JSRNTPIa/15
ERdyQse5P/eySdETOuifo/zFMu1yXqncpBZ58gsCKW2vpP92VHB+rRwNzKzqsk05
nrzKnHERErxCu7WZZZryS0lnAkuePL7ZT6SD4G6axI8w6mLKVllTqxQNNQD1oVRP
A7y8Aon06NLZ3xU4dcq5Fu/qtZem2yR664vItAWptE/5V4PYUcGyFA0Wgz6sXi7W
m5MDcXXL/PzoKkSu8SQEEzGnMbZD/GonyHQG2AlimsfuFXogXgMA/zgvxG9a6Tgz
uMV757htWdiFKdojEaPDGK9CwsCALyoAzkxdztJ0I1dod+My+R7RU2zOuf5Q8GT/
VDtuV+9OlNjy9QHtiJa9jhzDN8fKb70qxvH5i2IPDKrTwGoUXz+a1KF3w5xhjAlu
VVpS3HyfBcQK1+gg8E9299sx2zE16xj77syeZLMgxpXontrDjJt5x9HlJTRZR4IT
EZy4PFJJ0hwyaUyhf71Eg5zYJKyvfKc+64uMUVoTcVDIRJHAtqVw4MZgvcWtjDCx
pB9UzmSdmnbd8xpJGs8O4Fa+3uGoL2BEWMTxkUofGAOrjjHTZJmF3NkRRdD75XVy
pJs5Nj3QYQJLuvDjUi+2K033Plmo6qrNLZKf3jeIqyyKyGw3ckGgpY8/TyB2JGWT
tVw1oWU/veaxB5YhU1aEUeZ0ZNwjitz3znloUWEURePQAPZbHYVH0/s/tYPOAxwg
e5gL6ytVQsdA3Yh0hpJZscnP7Q0rzYMw1TVNWKxWeG7XQ/z0euX+Ysqpad828YiY
ANTU4kiTXi0hb3Obz7n3Q58HQoV6USt9Br+xe5A1Ex+mTKPHezlaf6AXu9a9h9JV
DUmGPl3zEIqhtSqDRJTfo5bZO3lntOZjSKYHTbH3G407wIC2hpW++aE6mRhotKZR
5rK2PxvHQXpuXeberBXb/JyItrc0yJt0fV4SVMbJNNmRz2bMuPsofkUI5sU1yMlw
iDDJye1I/T+EeWbxMrAx0AVSGRXgQo06ozWB2RADgbKB0TLGhIHIFtk0sNGT/33P
uNCKPaDJR1fYjpAkfG24CpDgcYEgVhw+MiA29pMAcp72STZkueDJOk7IOEFUFa8p
BIjNovtcUYReM62Yp/lwJ0FQdy+BYifm/826LDmw5RhR8TkJ3feA12/7LhiC3XIi
Twt3T1vF2kFrXs6Ndg28E+TyifSRQ8iok5EyOFGqDEJbHki9t8nI7AWffmijv+Uo
LupXFcusma1P9vTPWdSCnbUnPW2ZeijF7LZ611t6APZ8uyofAEwiqBmFjmidVLLa
02nzSZQJLceKV+lOE4PRJmid9SGFLBLCqljWSq8BJ35NLPMiN69LotlOlHYd0I8V
yDVAN6qdZL/GIN80XP+a2qlVX69ef5JD8+ghxBDZElUDv5LwBIj1yvqiiT7tm4fM
iUUfKI8SWAk/ighytd6D8GyrfTyKsaG3QemZSzCarHGoF2TJmtoDEp9vNLbVRfUc
iCqBafU1ygnAtIPqYGfl9sOQfuP6eoMUmuaMi482p91aVJLAgBOh9Ta0MYy/71Me
RRWmjdrMeXwgfE3rpfNURBPusuAUbrDxN9Xru9Tt6t2wneZDGjhlNp5FGXYy/i95
56g/U5hhmJ/S2W/l5zxSw5IMSAbLrzjs5KTOx2e+Yzgtmw4Z347zM2CnAYOzYDtd
b/q62YDX1+pyR99xtdJ0aW0QlkZTsjWlNw3srav2lA4/efBo5oAa3t7Nt+7V2FLc
gTrP0dwTQgMojUrN3dW10zvRn9/Sq6eRPfIW6USB15ScBx+LPcIz+CuaSwg4qbx7
klfRJmEtLbpd3ePx1431hwpDaGAygsgjVdrQBPTWNM36iduaHKRAmTmoyyyWOzQb
IepGh3c2NvPvpeuiVC7g9oXzPVvu3MdEs1Z0J/2obqQRxByPDsgUcrJKr1j37ydC
TqLiqExMBl0r1u2/w8nvUS0NofWS7YGosuULAxzEp6p2wCfEbhb7EPAmYsnrfgIY
jh3JDAKpRJs8PwPFYGzTqY0G0MIK/mYiciADxiiIuLQyIdtlNKB8UAfTXccfSYRL
9duZY1EFhJPNKZDJvDZh4/tXSIDijL3BjHXuNwdEJvXdt5uzD5Hvs2+CF1qn/TaQ
mGyotdokgKwh5kxHaJXL/SC3ebXXepCzmon/GI5IXnDdQDgORowULL9dEeDcCoJ3
DN/7tYL0Z5E6+R8tpRZAba/zfdzX6phpuzvmgDO//tTduBL9aEbN8/HwOu6KYUo3
7tZYIMoVmw6n3XaPVF5rl0MHb3PKOFzabwJSfDCBv0JXpvooYBEa2GFNQTBy4C3I
Sqw29DMzeCNQ78PG8pe5Q1AFTby3bNtiy8VyF6Av8bTQcqhzTrrxEHm1nheWokSX
fOsy4iXumw+TRV/M5MztIkpeIzFrjeLarq2adW+wjbwBAjCYOvx6onzYTECbQvMr
os92MNrPt8E4YsmS9DrxQudHMuh9c/CBy42qdqsgz5lTg1IrNRTFmbm3S1MEj89L
Cz1eaLxwRZ7x7WsMD0b7Nra0ZB4hHjBgh6oLSgjER04vLRNLEXVxK2o1j4VRGvcH
q7H5JZmhSnrhICGUbWcgqE6lOyH9ba3mCei0IE154XgqapRoWi7bbetcpYoY/LXg
BN2SKMzDRD3aup1S0TxioNSE6m0iPHfVtpL+NNJBoxg3AZZA0q8+z+ZZ6uao9iJY
Lftd7t6cZQIjP6+qkOyy7JikdNk5ikko6RBCQKRPRU3+LlUVr2o/b/2b5ij79o7H
xP8CJ7fmlpgPR+GzeuSSwuvtopkDn0xJQ6agQ+cgYI7YEmodGU59RFZmCqcPyEJl
Zbu0McNrPT+c78nsUjq5CSQLKZ65nBuEgUdDwwRLzfPFz6Z94aUi7GG1p51D24vK
VfKnyfP0G9ClmGC9lJNFiecX60Ye0Fgla3oem0CvfzGh4sNCtS0lSsEIT/RdPt4+
CVcYrU70G9oMmqE2AGcN/YBhfcfIttT3D1YcDKO2DJJv3rgl61dunL4/MgsWCJ5A
0Kbjbe5+UHMwZoSK6w2jWaAE/j68uuORfiYmzA+XUlCVKhrI2Sab9dr0+aohKKOt
VQmDsVh+eca89+j6qsHRxqW4Rh2K4kqWRrSYnNJmvILuE9TurpIi6PoeGyfBAUvb
aejbdkePAxLrF0yWLWR2dJI4LF1aLFbj4ZVLWAeCxgjGPISJwny+RWFZR5VCsF/f
eRG5RGU5vked5po9t1sVUBzmZpj+pZemdulBB0DSW9+qdXNPfpPNW/+8Qw4VKZTA
IO2+umW0p6ZgiF8zL6gkGvsMsQrHNk95pjNvjGX+onxUV8ex8fZ1VPO/a3wDGLsR
Sbz/8Ohf/M8ei3x6tELAuOYadOcyDGWElaHn54/BMEcfKff33b7ry90/2tl/K8LE
pytFdQV1SFHe8YKP382SxAI6JAlxCv22aWMIVXgWG+JplAkK4HMbhrvDiZjXp6mz
eYZcsrTYZtZW4ODROd0WptZgZSFack8EJoFDgJwsANJKljQJ+C2tgnCq6k+G1nDi
tO10tI6Q8IpG3lJEt8xYDkCebhitQ//Tv80e3tC/cg/IEQTCHh9H5kw7yY88JKkb
qgACA1ilNAFmPxmQVMF/qCNOODx9x2ykl7OMS11BCMqVxjdf4KjlyW/xvTeFXRVc
LxP3APmfvWo2hx8PmJt5UzUoUpYkprUzBCuzBC5/v/X9xKy3AjeO6R3jY/NZiZ/3
qyXGwiayb9kSRWgnNWW9pYZPZvuvczH29MqUd2x0lEEMqK0J+g/A8bw3agK/sfYp
K7YYiXC+yVTd7bSM7ChGRkLjwMnXXUPGjtFd+vi6wFGjit7KF+7AG+pCW4X+UXqa
V6UFl/9zABcC8UL+O91yMBZUmYbi2HCGZRMdWnQSAq55fLzO02WXBcd2wIrylgMS
jAEqPrgg0mUVMh+iJiG/qhkJ4g6tOmb9nyobcIMnmJy34MuEn90OUG2FrRl1z5+v
2wSteVo7Qa10ieIGEG0ASsRmkvSpk+WP82dV6nipWHWm61M7n4lUyqoGixdsI5/j
++E/8hdW0rlwdtaBpX0+XtqwVHmSMCDMaj/u/bMt7FvnCZbXuK46PhXWiro8U8ON
qwRCQLJ5ZJtmwQMBs5YH5SB8LScnNeOznHjA30cWn6uRbiePaFrUg4ehwMVKdSR4
7HM2vpWNvq+WghxwkcBqInylM01gJ7c1YaCRFvxxGqVG8X2yGn4Rg/H8kxHcIO88
DXdNDPctDTVsYKAN6CluXfYwOLkX75jDDiyJ1Rcpi+ZAEEHZkq8vxcqiqzcQC2Ex
CZVaZk8owNDWVKjzHbpZTiw07SA095Zibeynbz+2RFUjZBO80ViXKLpJ9EDHV7Cc
DA11DZrp66XkpGSYu2VydujRM9o5O4W3e7NNxnKuvgGc/4yA1AsdWC6u6paMdUuG
FG2Xg5XrjXycauCy9JBI1LUy2cbBy3P33g1bgrm5RUFjRq3NcMH9/3kpXphbzeY4
P0QcDlNNfbT4Q3xomJ4BB3JYq97+E+EYW9C0oDG7MOfMhWoRyXvpLppGwA0amvoB
7NZfzQ8RZSiJ+hg+dSzARfsNYLPz1XLrwb2Ag66pNje2Qe+RY/iOdqCwu0y1DCuE
nJQA8y/yYVVx7Wpk0H+hb11C11m9FQY52gEefEI4uE3I0e7yzTUGxmgNKaQHFFCQ
rnIepmYfz+kE9UMRFuu0zUQ9Uch7jcqlkzSXiJ97m+en1xkA9+X64G+7JtM6hAmE
sn5CL6Nhw6gyf0T8kVnLfzYsyqaIWXH2wjJsPAf91NauXStUJ2x9/gK1NbIGMsFu
Ykg1xAquPBxZfSq7fRl3gxqXiNO+eWUvZ7YJvIGJ8LFHEqQCD/viuBEl5soH/IGN
TuwlHEOas5cXepvR5do7gr/5wmTYNn3BapPhBRt2qscIOroYXgAAWWD0T8Yl5yNz
dpaJvM+rDMv8N7K+BK6xC1Wwr/m5Hfdio6eDggtI8wcvesKj89Dn4KVy3dk6ALEL
gOfVjSWyfmX+zv3wnbKf0rKAal5xouDwVif0/yTmWLDwqv5Q/VZVZhptPlHvyMXm
RVCcGan9xw3aHNPRAXKZjYVU/IqUQ43vhK/4H+E7wvOCNsc0wH65oj/1wgKH6vml
Khc6qXehjwAMKB/IYbY7XD47vMJsqTgsHOmo7jPTYRpDwqaCTR8VUWWAjxFFV6ut
iB5hURsh45sP1yALkxDL1PA6jPqJCUuJfQ2Y/wbKNUBoQP9jPIvpVNuFyCQuZ60S
JpWrOLkLS+EwXSSDNA1247h4Xqy9hOMZAmYDOHv+Z/7ZdYOd619at4d5CDwYCqbw
F8sLdEZVxS7OotipHZi6u0nl8VpwoQPjfvU+LLjRF15ERicssh7Bg09kqr0PuO/8
bclr6pQwF1vFIXkRR4XSuqsLt9elod8dCkUdPmyU/hyRlVEp7vBvIQ2sGhmcazlu
yKnyynwsWCK1iHCvTVLC0sAkAN6ZuNcfwgK4+F8QWgHipkt3O/x9J8xquqkDuZV8
LoZBByBoAiFb2nnUWIqhnpshHxwKvxTO3nGvmMAnD3BmCy+1Pd+n3BPXM9TQNlE0
K1dQ/x7le5g+f/ISwcQjmxID3uJ95JBMeyIwliZFYQaY+OrxEHVERLqJduJiL/sv
eFy3+4qwVbxom66OsYx73vyds2gKEPHe5S6uQpW/FzJfOfVmCTlLdrKIK5Kl6o1C
bjI2paSYAS31/TlKVEcAUcS5+jj+1aagRQ6oyvCZGZywdVfcELmX9fG9PHg9Ww+c
ZAUB+u+yZVILb03ZjGo1HwFTQf193ubZ6cX29Jlx3g8nddN+hHWprT+SilqAuEvd
Db29nTv6qnKOFvPyON1HYArxw/AXXsaUKT03fsKOlKkg4z7cYUPpV9ydTZWqlXrS
Bb5mfuVYez5lHK3kCfkL7gS0t1OxHDFMLGpt7MsKI7YCK3oOfLnISw/lvYaPvvTG
/j9NHPtSfrzpWQd0hLR4pF7Z6NfyqCJrPTldIyCvOmodcs2DJLcGbs2E34Le9A22
iPls2Npji7MVJPhxWEX/qfSK0nWSm8Du5g5ARoD7+lg/edvm/IetLSZm3I3FbHzC
HGXnCX7wjtelpuWka1WB2Smxh7Lxoxbr41vA7O/+Th+UaajXw471ItMp+jevmkIv
eUFX5mryznbdDPmQ8I2rQDHRvkrvCkRmbOzzKdnIzp18lOqQ4yHxNPL/eY/Zk3dW
R0DgWlRi87S57S4WIy5QecdXONPzWT6RJk1BS7JAXK87Ke56d0CNOuSDrFysy3kl
qgMsr/9DH5iodjpVoICeSJXtTovqi8sWpogWMpdp1b/jTmNlJlWhrIiV6mrmgGPr
JSprpSr2DdIQyCB0VqiszEE78nBA4+X+pHJ6BSEM6L/zCMjH5Vcx7U00tzYZwWVy
/JIUH1grALRgBrjw9ternSUGrzmr2J0urkbPdx0ZQeKawzDfZ3X8NQ1JcQ7J+Vdo
G92KZcULomKURLmzwmDYeNPmZ44olOL8NW+upZJ7vltCiVl6zQO3FJ+blTqub70B
n2sC51I1J4cJMWX+Hvt9qmKGH7vPIn+XrrggaRId9OsRhW32HVVtCjVrxpqIB4cX
770Jvk0VF1KgfFNeD7xY9n/25Hp+0z2o+JcEOsk2q62SvUFgOMzpHnEmT1zkYzpz
Yz4eKMQfEFXHnljjkl+v5DrvsNbsFySGzSIcZcGSVle+dD587ExvTKv/PYa1SRLr
hJlaB9UocxI4wRlsNmmdsdFNnTkMPU2+Em7yGaTImIFQdw7Qvlm6LbL4KoOtDlAE
kUlK/XUNP3kdMbG9bje+LQfKqL4UUiOcRhD5MdexImxMSBOy5FuUiQ1LwiF25LAa
S8z2/e41e9/xbzovbqEv/DxVFeehvC+B1tLCnhxe7t8vd9/wIszrr11ewW804b6E
0B/A3H8JzlBJlX5UXYpQkBVAQ3chQaBg43ZRMhWIYWBalLKC1rt22nJgK1T04SZV
VyJMY6HgNj+LAHQFJ/gfiMkKmy1NuRvDDYlnAAwPiTOSIVH7XHt/ZnWN0PS4rQ2N
lnBIQYIoNMSk56CTwJRzWg==
`protect end_protected