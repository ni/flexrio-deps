`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7184 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhBNVMbsl6PTB5/ApNH6uD+ABMea5lxpzbviLFCJvUttO
BIcMUyRwD8vshJLkde6WoGDnXl5kkAUCG7eC3nYQpuAvSSF6YZVJbZwlo6POQ4I8
znPuuGUobykC872Ow+D0RwUkzABxcaNqoDSqR/tibmOHVK/zPU1T33rlZe7JqIMU
w1Uzx8I0KCFxp/pO4mKN2YPfc/Gc5SyMF6tGdKddp4D7/B0/y4WnPBHePhYM5II7
hnDSnxPPMWkQncEOByO5df/8KtjKDdeEctWo87a63OJECTd7VRn7fxV/ToU3ex+j
gbCP5Cht58Npj+aQI+yhNmTxGGYdEX6eTzepYLflHO/tGLfhCNqvCvcEdRepwnxO
gB1H1xcT7RL4/fD/IYsd2bwPdh68kq30uQgqn6WOGzrCJKWhNyv/aoIs3rRsTsTx
/Y7H+8CNjZorxqT9UdR11c3Yt4DZ1scp2keCtzMb2+avm7iUSKmWe7cxOmalDn23
rJNyBUm1L4ctPUts6ex0/RYhPW5aR/n1ZjywHAonVBmjC1QPi23XyQM2y1tSzEoV
vgnOX5pbJF2RE5MH8COjAFaGD9f5FPuJyUnxOXc9EB9RXsXjoBm4N4JP/ZkL1A5h
dsVKpL6z98sb1kPSsfLWYlMqx/Le19aOdmT8MtDRWDwkgN0tkqejM3I7Jta9NyFZ
dRXLdrNI9efV4wuJLr+cxf7lj+BvAWt4MMw1Ag1N9yP72YfWHz/4+m+EJpwH883v
Xw+ib1nN6XZlXbQh8Fxy5Qyn1/J18Gi/1MjXSqrAOgH5Ot9Tu6d6rdFUu/dPBYNi
QO3TQSIWwHYxLPCh20HccMjPnsx48STHr++NixN/D2H/cHJFr/X29vmzQxVxY074
M9VZAeT+CBuPTiVsFQRgtC39XwKeDCQjuoLp7cfAZfZS27LeJBp1oLOtaMF6h5Kc
ZGXmJtcbxFuctMvid0n3daPQCLuhX+81QvixOrkE2/3/B6kjIa3AN1vqcZD1UKH0
HqKsCc5m95TtAkdsYdMK4nhNMNx0SZgLTewjYDq0cOr8ZlrWUYpJnPrv7hJWHnT8
Tjs6rp6yhzAMXKUrlToJGfnhcHMNXBWavVgATaU2KJtdObBEbKRiiYgYN8PigeXk
rtCNpwBE6eDKaYOiGS262Bu50EFw5Gcr8nbtajZa8yu9P2NbtmhDdxfHfkCvjWNO
z1OOKKu7bUPCz2WkSbQyV7NxYp6kDAzsQ+RwkiV2CBH1MDYdnb7YEBdyEG8aHHNH
SqxRGTtLzBm7/6kATjNVHOqSmSiAt3CIQPoFeAgdvgmWkNR46MNKTd93Vfdi5yyX
4nqy5XRJol5RfcqtxTXb1JS3cGnQNFy4mbURg2iRRmK/I57CzjFKubQOlkY8rLur
UFFgq3UbZidd4duzCSO6vrF5aEhrlJdstPpqT+tK6IFHjSrn9MK21bT0N1Sx3Eum
Nk8vw7o97/ji8Inm5ZpmYIP0T2CjsfwPM8Nc52fYeDZnNN8r9mQunASRazESGs0c
j2EWw8jC6A0thkA/RHY6Rts+b4MEzTqtJ0qP2YNl1AKe4fi7RNXMK5V+5QPk9EFa
zG/1ZsoU/u8MY+svwCeZC4q9hBJ0IbpgoTUd48W4WlYy+xrSMhdGcAX7WRfg8nG4
mgG6NVUlyh/RuT3MrNegLxfB8uPS9k0UZZKvbr0QsNLX2oU3i6yYGrgiGM97ps9g
yxPbrtgJFm8kwJzNBX8tg9qfvfroM8lJdoNEcCiGF7xT5BuPnBSGXl9/0HhCmAKv
+durS9PcXQSwPpQNW+ApOSFlMWSK6o4jwOgJR+ZpH9yF6e2rVF6m94YWuzguG64f
PGAHUCkIlnPR4eB/DRuPtQdQXioBVcarTpx3JuzU+cwwMB6eiFqqIOBl6GiA4ky7
sK7hyEMp3RT96T42ZWZMFBiy4O1FAUy6UAWhZ9FRKGQUtPmtTU/3w7dOVpwKNCZU
XIklOPfiZEsr9elAq81bd243tdlAYEaTN4wprJK+vNdJK9u7l/yVxJblO1AHo7js
RHiN+W/wRUHK2fUGHg1tfG2cnwdfgCbkJ6Nxmub9Bz8e3iSbmdFcKzcovY5PLpFG
zHVrAe49BLYwZsyEJw7B7GUam6mhawuZIxJqupb8vGuMxeMN2ZrcEz3eTVa1U00j
SAGzba/6F5JlfUyyUFuLBzseuibg2c5FgQWUscmzz79m1sNyas8xpKRK+KDsah6i
NT5oACVnoLBYSX+q0LXfY6IsCCzjXBZG55kAwG3pOZPE1TxYm1SKU6EzeHrKJvHH
G0fSYK9HhWik4sxarI4GtTgZpmlYO3SHi4A1LKqdCxkfWKIShNSg9+sLNez7sBXq
Lc2/TKRJsyguPv8denetk8ELgIIGI23lNBqRRkJlvvZTa2fO1WnTap0biGmEf4p5
xDrgDrByCmuyFOUA9GEBbwYfcEZYZw4HsobUbLXX8V1w4eh2ZRvDzj0jqZFsecIe
8SWxjyRcRtZNzGV6tQww2HOmhuCw8jfnfwimgqcBdw9m6JuNslDOYhs5eHoOtyW8
gIpLKLNL7IlwztJDD29ntZW8worJnIVjCBHhQSttvyizQ72KtxuhQas0asY5suU/
tmFlm+bye3j3hSbe/y3Cfkj9piaKnzMsO+nXU6p+AljE7GIOW8YknQJ7lfd7TmZ8
uj7nBqiu+7hSbKygQzenCSGgLrYraAuDIhtBb+lA6q4Lj2e2fcLu1+KUEbmzdFx2
KpNLoFiPG2pdxdmXiWWqSRqUajDAOsIdxlSSgXFkkJRhRZ3cPWG3/1ZTygbaIYpg
uwHDl0LiSTT97YBhtwhDWqPUy08NHuskCnp/h/y0M1mn5VQ0Tf+nvNGoej5BCaaV
/kXvELBS1LHO9Cpn7L6iFTpIyCm4Qz6TmLMUhIGSnEW8GQlGr1Ab5R9Ie6UGxUeA
KcK+BLb5PQqkeKnAx6KP02oaREz21CFJcA1tsrtTvuA2hwAN95MYW58nw0xSpm3L
jsuDN8XPCBQMtJ3DeSPt8mml6o8GvjOQvTvPEyhRDalf+ctPw8EfPOnPbpoTvzZJ
LEHJ7leZc/LabyJL+MterXQAtlNE4aRlhglEDhPwbOrkTr7aodrvHo9Dz00wPx5E
RGhRqmXyW9EtZfJVYnZySEOFOb686ln09lHCTUzyDJrIPdC0WLVykj4tdDw+tBwB
Jm3h0x1QjxJJb6NoC6aF9LZhYy/ULd0iAIiusvpNIVLlH9w+tQnmlJfg32NlcSVQ
SuEgSV90/YZX3sh3eD6elKCWPmrsYd+S/KSrwZhc2nn6PwZ8Pw3f4f4ytBC2e64W
1nvq0LoGzMgmUlrGPc9+pNzUIchT8jfPJh7ut1o2+ktfP6QF4sYyAfRr1d3so5EB
b0tMJYXwsOm4jpaS8MENXc6Qyscha7ftqYE6bNHXHic3UIAiXZ3Qj7EdJWfX1Tgx
TN57PpN7x0oHqZVHtWNqT0VU0M1+SMBVEIxGPi48JWAAXgjqc7NGmdPPirGS5bYC
6a3RI9lahFHhC2PTTmtnjMPA044hmY/VMdeRQyVYHy1caWK1fK3rY3zlw5OHvqs0
o7TkaX4tuY1+c5Q/xqpD+oETvAqFtH6PcT1cTy50tQEaA3Ag6FV0qzcnP7L9o3x2
AsRJ5i0ExIRvyyMacsS1+psVdGt9DMx6EIxH/Xbkoq4lUVWvXjK5cxImOEcJa89H
tSbngt+HnmpS7ZmjUJWTn9tKWZPkD6gdeYh2gvENHMNNmK/DJvvCfFij2vSKVhIE
VXAFO77jN/OCvsnzkk0Xu1a/kOgTwk5u5v9dzcIDhoIqeo2sQ5AS5Kx7QGaVRAu+
6SUJ2zMtKhLiH1iXKuwe8r6LPfHe4W0U9QPoiT5v2rFTwvT3k3QdLXYuutIf1RuH
xemS5bKM67kY8LWlnlpk1lz9TTp5w9uhfNYI1L97+PDwSLxOxohF2DHBG1kZrVJX
ukSx4N/STix3gujv85gLnVdCF1du7F2Tsq6rhWOEpKW4j3uyx0quIbBeyZ4BUIQo
0CQif4mqEup8Q6WNW2eEQGzAc2AypKa1N2d8HeqNDd09IuaNcrhXY6W3IKOi+13z
PWYEBRldZQP/5bqflirDjasbeRXswPx0avRc7lfNWaLKV2EVALL7ZKNptAj66Osn
waM4HNrEKoFtIRjnSC95fJ/I4m0tLdLq5C0yhA6dZ2BEbWvRRCZJWgj4b9FGE/sS
R33zyLh1v36f0u+39xMCm8WUxVymvOxIMIhE+DSDgSLhmF0lVD7AfF+qyrQnEiQL
1utcRQ1ZN2P5P9R1pWeFHRxZMo2ERV/4ruhz3zKq2mIqc3KHmhhVv8/g7a8w5uuX
TDXFtesNyGqpayQnIGfTJjbotd4jwYb9T1+WYP/n/dq9hbUBOFToTjl0hy0oASfg
mPh+Qd2OsYLijiR4L8Cq3sRDakoChKZsd8wSApnXIKcCONxgASpQ+GRHbnQ61uwr
qyYNdcDC55wzeMrLB/L6i6Uw6l1lNHdGh0N4tKphoM6uJxUyWyUUlAzgZ78wuDh3
RpCsgQsT/CVsXo0oRFP0MaLf5ApjJ1lU+6McUqdVKWnz/0xvQ4n+mhI3/2xAE0I3
lHrqmtYifOrOkK6SX/Sc+kEyKyNjdoSu/4ZMoN0YbSXe9iUi1yKcMwuJ9YvpDoAN
rVgUuIjPnmYjBYcuoz0z4t5NgH+oi5OI+oIzpN3qi/9/Xk/NBI4YnXTliZ/t76J0
nVtiXOWjh9ECHV6c67Lg24mqO9DQ1Bnn1lpNe3GyVwBko176uicz0n88dTJic9ni
vQixSs3wtdyEqRZHjD2X/0h0WKw1IKdNvM0yUqNWRw5mn8pXKkkluro9vY+2L1Of
3l2Nx1sFU71pCch/9gx8VUa1BfHt/66f0K00X6YDhUk9lRVXZgWl5eI699S66fcr
iqPz3N+9Y76FIapIhHmUxZe2w+XMHBnjSAFhvFjeL5JC+7WtmeVXkmXvanvYVLcR
mhzm04/S+x7a9FY9APkS3NUVLAkL85KtzDXBiHwDQDyvleoYXZ1n+LETXnKK7SU8
pGWQ0YFEwRMvcFH3jfbvVUzcaUQs9ZJOsNj4WJJSQp78ooHy+7ekC5QgY6AgHrXC
F49xyucItSMCuUCevYppy01T96d6X4AsmPTrAQjBx3bQUlUFwMHE0WMPpdZpbLmj
+enCfSgPpVQP1bq55MfeQ+XrRcSgZkvDq4MQLIv5/6rpsRmkJyPpc863tj95I1Oo
Sj6Jftwy6zrtSQZE3U/0m5WAV/TwYfvcp5z7qxIGuaC1zhDwmJQWeKL9s02V0aBv
VylabtTW77uYCGGNl/quePqwb5e1MFf/IVh9/iUuV7hwC1I1dFprOOHWs+Sjot1/
dDAKBu9AqvDyzlqK/yPWcItGIWQx2lauwfWVQW8F2fKmTUW5gP1GNJX7Ek0yJ/CN
ehr+K4i+QZ98iPmCjW4mlJEEMEI7eBLurONYIeIU49PP1bzI/P5Dy5XPWWlC10Hk
hwiuXXSan57PthIcmpXvFimQ3ouWAR5DLtC/hXTADq9ikWhNKidNXOOJ9A6ZNn9C
8gkb4mxLxRNHSsKPnnZCO8lXgIFG2f27P+MMq2XjTeBf5gY7NXSeb4+ApeWNV76M
xnjPJD8aXytyY/qwEkUirjV7LjJAbzNszqcqBGzYGvqRLLlBJj1gcm8IR948bsZs
TpIyTTTaTPoy8Ljt0SXmiVTkxBzlBSMMle8PpVkIDwU0dpi0BGwNqZ7zteb3+PpN
rQ603EtRLG+x7Fq0wH4MAtYZxaUPOPcEN1QF9UMOAcRq0kFIPrwwBqabdE93Daud
2Tao1O6ImdxqNpNcBqqp+bW+0Qj6lxMGhn0ka6lRKBFI+C+pickJzS3NF6x0Odlp
udbHOVzV+DCaj24wN/7WJU9iNxbQtf7JHr39SdeSgo3szyMiS2tGt9m327vOwCEv
Owx3qOzTWIDVDfTG+kLFrJKba7LU7WbUTUmDy08+CD61y3YcitBwcrwZKEiY31RW
UsMTMvMS5k9AaFERx/PSAempfu8iIPJk/UXv8Wstt88oWdU3QNPWWb8nBZ3WGxUS
Nn8rBgbV9pGFivdWPg58AbW4Qd+cEkI/n6cFfJX58qXiSxL5qsVfKpOwMLyE01Wq
CRTG7aSQLQ/yHZ3Hh8oA8w1/DVa1xNGfqYrWNn4qYbwcin8ZBXmIiEYkCc6hcxAO
6+7U/0E/9w33XaSS+EpKFTAGVjYS483gGAMU/sX/ijT8WcoEcM++lCiHDL+gCYQp
nXYIO8LO38h/nSxTkLOBZh/gQxBoAgu/yq5z60T0RFgGa4UH7S/2/tGmx0/W4XIh
dXkpt5qi3Gjb76qX77OzF+zmQjhpqAB41hOC8W0aAwS6t0oSpybd6T/uxVE0wFIz
MO41fiVn3cHyAdv4SBhxQJN2RBbvGUK5/fiVKLSRTXDgSn0fZVotofu3ONSdKMrB
ErBFc3AFYQFZuyN7qyYMnfHRnB7VjT8QkjWIN8JcXGN20AB2Lix562vS9CtQJKMA
4ilSQXaHPaZK4zh83Y0b1eVdloDbaDDLSFjGWgb8mSg3Pxlw0Pr5Ydp6qRSZJZt7
xK05I8Ha9Cko60uH6FgJiBhX7ykRsknVKxZJ/HSK/V6mDRHGi031JwPUCJ1Oex6e
1Qx7qCveKTT4NNL3s021xCsY0rb21M1I8u+sdPlWWGVyz/GOQZQJNlXFto5xh15Y
eG6rNPWo/fF7hksIlA3xQdCZJzxThoOfeIoxWMmOBfdOI4n8MQU1oAZdQzV5Oql/
gg4/WPCMP2eI7UmZfzXfX1jgIgilDzGBxQOTDHx9PFFGxYA+iSXmeBgWw4JOW9Ik
yLHRXw3AGaM3YdFV5Wyh6PM1mGIKCCmcCZaVay1KmoWZILAyxhGf88BEEx990y2T
dRRahu4aUSQzOf8QBcs8Tzt9iVonAI2SZycXbqdUY+S5zofskaWMBOOvcl3MxkVk
sAj6eLmlIK+LYNTguLuIyFBWjz8LGYC8g9MDLonK4yZ46PATlaSNVxwT2YcUBpd8
/xflTTZs/xUOf5UvCA+IHaDSaE04TLD8WVRqpbac50D1FAOS6X/IjY96P+Dsky9S
95xUNtzst79utmjmu0S7wqM8R1Ay12zg2ZGpZfNYkwR+AVFS6AZ0Xm5AEyG8a8UH
XCpw5B7vp1FNKDsr/stz+7CHawqs/FkwUWeUt5FSLkbu6nx14GnYw8K8sZBteTVa
jlbzG/V8rkY6yWTs0q7gzgWKFPH1Qu5Ospm1NcZH4rAqZusaZt2ruWiFvTolHW67
10gRICCi8vCPlZmexZtouYghxZaA/NUhULlOlpYVqqQf+4HC48PDfrRixP/wCRh9
ReWY5TWBJQSlyHcICGItGxHpJjV5stdJRH6E6udJxlf79VpNJS6haKZ5NgnkqdNt
Fz/j4fFXOv5RbjfzVcaFFezp2zdHLuajbqHdMr2NM/+ZAkoQ6QFYk3qzhCMdLiZd
s+h4Nei9Na9sDV4KQ/0R93DhjLkezF6D726JREqDVAAxYAcyZiWLejMhr3s9Q9+U
zRvcfE9+NJl492TKLsienf5mFBod/m7JUfDjpI2Un4ckzsmRbfbb0eJhOgti8tLQ
TL7SlsAhOBa5qG4UN7Gc6DJgzIAhNf8WGmPFs0DQdYluM0eU5/k47XDBivDlgA+a
SFd++W/jcJa9q7l+Ht42iGJKpBwj3SIWrbvokg1KLniKI5klWkkErbwNUjKjKbJL
h6eb87dQpRQDmdBe7lLLsW62Qmz8w+YNK3ie+6wyJxRQ4jjtl2ixunR1Reamux8C
s2wfsHvp/br538OG+G10cJLzANNlkmTZh+HB0W8tbzW7XphhYtcfsL1W1Xwj6rKP
49mAxvAvCjx7zecGtt5lOexc3jf7gl42ctXtYB95X6IkpP41kAObJ1fB/uIfjhiO
OnBH/LFUNKiVcTPLAvAewMt1IeU2cZ/shrL2qrFSunhQFfrMc4SxRg+ss1Fj39vE
m1FF001cNa9VhVqNzu+rMPRJ1Aig+WfvL7et26CVrUPcYFNYQ6eOAkDcuCMgrDUa
lQ6CUq7k8UJiC/yI71osqMX9g/r9kRU9ma8BnKfpUUzu2xTppiKkHmOyU6f2rHht
e54pVt7PCc0Nw4XBX7dcf9rDggL97ayiV4d7d4RZRHt4BsFHLIV9RNYeNjdGDimQ
TIuJNkGbia6vX1O0c2fsfHT71rvnEQ2TBX71gsoAsKHrtRjv6sQGGnqgz0tGerhT
rXTIkLNkYX3i0GfVuvPKLHAzSv5IQlxX3pCwuvFqne+I9Y1gRU8VivFbZhS4w+pI
Vyonu7aVKw+bfPcE9tkAKGsJD6LoW5a5LWt2NQ1+Gsf1HEdqNTysuAicW8Su26lt
vbQKVipfBE3jYVRz3fxnqO3eLeM4jmBZEwQLc1QmJN6ny3ZlMSHDUjIlmZJ1qIuk
sFV4KwmLyONRZ+vCeBCboYBjfowK7IqcJE38MG9phi+oFaHCwe3x14kWVauSobDA
jRLlJ6CsPJA+V2OwIQV1mQ+A+g7q4JejHUnwc+o9x+8Mamuqa/2ufmx50UbSJTA6
qZ/2ZvHBOB6HdQw6qNWKKDpbQa5REBRCdaTZ+k7sfcptQoFRe1IrcklKWIgHzn3U
2BPXE7WZzlV2APiKu6+9P50wVsc0jFjXyXu8ONuc79uq7USmfP9/PbBUE2pDxSup
Nh5fspuVur3cR9x6OFiltqxf56qYlLF9+eXjDaAMxBaYYOBXRhSSfkzrqaYJ0iKu
5BEngyjPtkGJQEtL2eryKIjxhPL7suI6Au2ZwDEWEv0jLGmTdjnu59iRNNZEfrKA
sYffYeAmOt3MHczVltUQMEXwC6bxxXju+dD87x+DY1MGN4TvujLXRfCAVEnw8Py8
/AtQIXUtoSC3JQOJAT4IKUU7Z5jx66ZUlXJmOBrSO3Ci44utfDQBZUtmr1x+4ZPK
Fvj99rwMP6dVT/P+5jVX4mRSmr7JQ3I52daEPsbNgbaWtiefQMetTkuN8HuAftEg
OQgHSg9uOSwCKjXOlhljjyItRUXn4VHSJKqdZT1AO1FcefIjy8sUxOs/7HZrTPZB
m0K7DPWio+lYl5a21sprLpaKlNEvn7/CD1FGANRvvFtffD+4jjxcagYOgdWCvqqV
EoqNMonN9SDeUk6WsWSS+bHnr+Y+fdLBgS1mA8oBm8Dp/draAaH61NIBHeC4tRAu
OBr9X4dVypYGc+HoWZ3Vo1KbxiOKgRFm2nGP0Iu4TbnDhMo9vtjw0R0BhE/dMQ+k
X+5qLsMDpaYwiI3buhrqU6w16C29lk+1LLVELApTbSKsJhDSQu560jkRsrhd9Amp
zw204bdcC3YzaViaCyk5+FAHkyFYl630oEKJ9vIbFLZSan1bS1QwGKbNwhZcZgHS
G0TJJ4f2K2T4KJx63B9Qtqosg8fWBQBdOrQX7YaY4Uk=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7184 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl7TOuMe4xzV7rdHsSWg325trfZrlt/zHq38tHZh/un7R
mH4nP19Gt/yOeSNiUZR8ZQpgPyrYjaYNVRz/IkqB5EjSEF4wxkXLOKUtPEHfKCEj
BNgB/AKtQboRp/AVj/INkjBFLlALqLBTUmwsqId202ZkKmFRMUhI+H4TZkwTJbsl
zvsNHL+LyKDQB5fq/6E19EUCAcDs4cGjUzpuoIjAbGUOvLJfecAstSBagNdaaGxw
pGrlvO1Orm/zyod35ohx/WFXQKtn6jxuNPzGAaI/HMf3Pp3BQ+CqYqoIRINBQm6p
/xXRSwWOIJluFgqKyZI59qUkWZ/9Wm+4uEs+akOmgslOEjtYh0l78S9UCCdxRQd4
w/o4lnDKMHmvDLjrf2WafbXX2Kw1VD2TaXGDKc9CcHko24isNEFD19W28dlNG34Z
q9mVuZSzBwsRH6jctVN3Bd5PMv/LKuCer0OK1PfYak2pChOW8s2Mw3U2LuXnZDdS
fJmp4ZI6YOOmWKjXSOOXjF7s2KCOlIg/n3YpnseF8m3aLUcKrJABkH8YHrx429k/
4uNWd+McYQCXfJwNLY8WM61JfQjLZ1kYJaJIiXVcY79ABMyqwCCIOJvDF9oHPIHE
dokVVFut5RLNNzE5DNPGqS0RWhuxIukI1b6Bqni2c3oe+ILOSsbPkRyz4rBJIIzC
2r41CTP0SQCy1i6+rHb/g2CXeHXmdO5kVsOM/nJ6JZxJEAXiW2Hb0csgRC3Hy9v5
BLVGZMLWZV/AcWZN2cwx3Ul1UHkOvnB3aHGzZikruWfrES9ip4ZafevNThEQH72V
wBb77G8fbpdZeD5pMPkmkq1eT9COI3vSpAiE/dyVIHw/6ErYuw5OGxmjI831XVla
fypr3/6ur0sGzMV2asEeFSj9yB5ZkKC0A7htLSVjC+GZBthPZTxx8l4r+iFf7/z/
Z/LproAU+gt0AD7NKY3bEHHW1ZDsn3NJgwAr4yR1mUD2fGI5I2JgddGPnSUeIjiB
iBW2dXtHdyYwsvhacLVgKnLaGbjGyRQFinmIumcGDG6phIl9dL3NEVxWCUo5khFa
6c6RUSLDfpgWhIbsBfPHPlJiJUmvvt3Uyt12PTwwA8/cVi/tmrTBjBZ9exYHw9/o
wtHfa721nFiS2V6N2BX1XV6Fu3B+9E7jnfkZpJi67FffPkBwCImxh8pFqrXdoC35
Y+UgkDybW3XIYQP+KSSR4KfXpQ/JSQcAPnzbfIkSke77TGVOqkceT3bqge5bK3X3
Wv02pG2y4zj60e5Uy3YokFQrhqohIFqwKP3wjNYTmiCnahD4Ku5dl+uB+2i0zjZR
29mA/lhUChNIe4dFWqrXRY94+yhw1aZHIxpC60K5iSUt8BjNwymJaLTljAaO6asl
i1q50e50AQ/AZ8u5NMJrJDY0KYA5XK6uOTXjPK15N2qKSwdMG17CUAB5E5aPwa2x
NVfM903v/lyJz65yPeg/qOrSDnSo0W/ZdMms8+RShlRweQfKdtKi1Dbd4yuXmFBj
W6xBULh/cLqA+PWDI6XkHAIc2bcocR0lVb6deweslxq5RiQhHfMw4vqPp+laPiYD
B9GTs7G0t6d77zBnZuoAa0eOQH9mhk1Rcx6qMOFFZkNRbZETlKGgS+DWdCLl8uwO
627puzrFZh7LhBubnGfv70e+5xjK7szM3xMtHULGPBpXJom93+p7H5PkK1Oa+/QY
+w8y3xjeWj9FU4m37fN6QZXv6W8sZMOHOsz2SfgPqj8h+GHMFx1ghbC+1hd7pSia
b+ONOXiJ0vM2IeHWMw08OKuoPX/KqHK5YFhRAFs0bnInFCNl4PLZttTpUI/NjcJY
apR40szmPCeFXAPXAfyMbYc5mTptQZE0MYA4HgWmMIAcErwAUX2oPXRs8n65VRZV
AYs73qT2S1jIYLkWtNyy9nga9gfhNLoZw2OzOMdf3ccmsLkAHmQ53Ihq5Eg6UbCi
RZRQO31tbIoqqpliamiS0QQU8Q1ATxZUqhkRScg0ZpOf8GJoUDbcEtr9LvQieI4u
ukzSHTRhPT7yaMR9y+b7X8JPdXvdqW4Y5rtxdxzxi8oRcknqxT3hdz+TWkkTQFDa
7tcO86E1u0XngukHSJb2S0nVuDbIsQWBpvwR1OZQihd46oLa83VXGKjYJQ1GcA7P
ycEPMmrr1O63FnweNNw5a+/C02jfzk32B653UstHGEBWytCn+XhweKuYSk2DPhQB
yzZgUtpnUgLxP7PgWKAYcBX7i+HvWsd3D7aMSzNpTttEKpp90N7lqjseTSogxCVE
DBe1C5s41+ZBPGsAtTy3xc/7i/YoGio+7ZBdOc/3zB8BFTbvPU2u1CKBWoKcjxcu
MiO1EzLMoQAZkU7B+34GnRo+BB4psUmTuVKpCovQVOwG8jKeSHGmwSRVnJ9LczO9
GPb5p69yJ5NhcoUIFRYfVaxG61svPDar2qcW16dowqnpJJtYrAgUjgJKm8AfTk9s
n3FtxSrxIYhvi8GmaioI+V45SsM/ETHNTQbh7c60hNFqjM4jGvAtlk6tq9BQQAEn
/DU3TfzaBe4AWy8p/uFO67n5CUkCpK5H5YRHMI0z6iF2XRF1da0yb++WZB/hNh/V
BS9Dkh8WkB0Hf7BfjZAga/gWXsWTpVZpxtli8syCObFrz9y7H+HsTVYahp9vQFaG
06upO+qMP/NIVfRO+jzFmrWG7U4w4wsdzrlm+7VJk4LuwAmsiLyOYrNJ03/kQnPz
TXQiC1IU9lStgmtMESUaf+x/DZ0zWfewBFLfS/67RVEqQ09tPg1BZPa+MCU/LuGZ
QofS/iC41X7b9yL3S7SkkFcgwE8c9a0irf/Aa8kasfLBlyOUh74ZVhdz03Qmt+Rv
FtQzPtpu6tpiASFZna4G0pqM2Ak4E3YILozhSEcApG8qaQKkUw42mNqDxbkVTSiK
rqkZvwdrHeyGzPeAt/OSty/ZMxqTqSnJtK7NTTv5wDD+2Y1KiuPAbIreQCLtZXsP
o4hU6DdSnfgxQIgVB4/moqWjbCmH4TjfhE30Jy8DatZSlKcxTDvY16bKDrt2D9vr
agT8UmCypX7O+9smBb4t/H5LrL6epPyEyaLbcrEgIFWKhILBpOcFxOQzrkYY2Ua7
8Y0S0NWJVx+UjhDbTpXpZYp5O1hG5x6ZZq+EIii4yPsoXeDLOcdFhOmlyXHNYONQ
uxu6HDqdUqXEEwMs+vVu18d7/qk9OuAyHqXxSFmL/+n9ExTWppKsW5tQLiVQjumA
/7iL6coP1319FGB1vmRUmIWiQJt+aR5tFW6pfi0awAXDCkKCcz1P3gbVOM/yOJai
e4LkEqq09heVWKeBeNMCKm3nVhe3D3e7o83tQsXf/s+AmM4JGohHMyehYewIQi7l
1q9O6Y+ndZWro0Dq5ksaNQ1CluPsad4B42iP8X9uohIIvODU453czprq/KNsGI1O
N34iz1RFNloVa4FJX2AVGSHqsGOswpvULYagK44izSWn0+/Bp6RSYY/6MZnknxfu
vOUva/E8DDbRl52qDCQ4dLjeQQc5sFcoP0Jq0/Fa7Wr8uNu0xPX7+XUmxhITDXAB
O79M9qYaBL0Us8f09Obft6TXmf6QNorpLGGadUgjzSh/x2lqRGU5qUebwhaGUCdD
03RyhgiUrnKnRNZ6K98Zn23ruzlAms9zFNOOUxHuEW2hCXXvHkbiBtBBw7+XjpEL
EgIwQIbVlUJ63JATpsU+2/+PKUys2zKycONybMxnY4ezdf8GzDQp0u63Ab1aQD+4
kx6LFqdDIwikneXbz976hfXlPVgjr26zpOkEUEWanOzCHYSK6QSAPxBlOGxbW2AK
suJcCWlOpL1+goOHbRcn0jGowa349AypbvNkTtxdzGMBsj4q9PJzbpu4do8U4GMP
+LP5eNbSWh6fK4oxxWjhwLCy/pgfxBRLHs6yolNn4HIitbBVznUZF8R9TBmkyjeS
Vr44Y1wtpIfYYq39e83aNBWwdt+VgOWo9zngM0d0bymBq56NKlBlKSmvzbTCQpT1
wRKCHhvGTQdCCkx6H/Ltr0lVx1tsyBuP0yxQagWjzLzWayeibuAJbEckjTAlWz5a
RyKVvslT9/J6N2Aalv+LsVG0HxoyeHlQDJFO51+1HNsMmss4lq5Lkqc/X0UXF+o1
TQ8qW7meKiR1jUiNHlmtobFe7bB8kb7cJQeD4U3w226AsGkA+YGoJMfud/WscvYP
idJVyfuMbgvwJQK/TG7Y3vmBhcP+BDvnaA7Jv/StZtEmZC4atJiDXUnVEg1TJrQ+
uvoNxIWsktCL9Kb6J8X3X+zgvDaZEZhXtfYh02eFnWLIY19Fxo2gX9vl5/aMmJ+C
8Hj6GW/2Q5xDB9lb/gRQBw/H0dKLLTvp6IDXIniJDquhi88PUesekoK8KMoflWlk
t4mawPA5PrDkYTKS2DoiTPp1HlepxOPtrrxH+6kpYV14PDTk7qUzHFOpl8VHCBfg
LTQl02POJ97tWGiGXsC1uyZjS8Q3HGwv9UWnM2GVRTz93oTTgRAXlcA6gYARiaJu
CfPnbuSflXczfImC+SP5DYdjngw69GiWmWgM9lmxkZ9vzDSY59KZ0DPBQgLD60TO
7ckJ2UgJlRiT21ZedE4WSPvOfIRpXzHjYJ0JV6PeHkVbxDkIl1xR1FltLdjVZ8Cy
TaOkjsw/3YSM1LtWzJzcsUfBnpMdW3r0NoxiZ1IvnNvEv4DiqppX5GpEpu/1KePY
Bh0vQQXWDDTydT8XrE2xCbexHQ/EXzs4+JGv4UTEuA3/s7UE8uz8PpCZQi0m3YHq
op8ftG21OqeBckbcrkIFdAnVb79XxAMys/jEu+N4g4G5BIVK6DRp6oRAuE4vVLD1
TDY/EnNhs53ihu8rpULnbi2kXyeCggZe9EpvgEuk3mQm+3DaolNLHP3jSwfRDdFF
S1gyNBtGHCUiRQID3z71GEThMZpyGCR2tTZlwmkHhFXAfDddpx8l1rDlP5/flS5b
Ux+l+QKPyMkunMsT5ZD/hYi2iJM+5TwYUQDGEJ/aMCjXAIWAqojQh+98YLpCixEV
IBL++/CNERypaId1VGXIycbsjBzUtQRaNdQm50a5eJ+Oawvx7SpA7XQVIKh8+6GQ
TpeU6i+afjxCl2GwmZAHPoDuPDtWLIIsnj1j3QX68DE4OiAP96qrxgbIbvSMS4Dg
fnlKgT3WbvnEYrpCyDg2NSx61G3c2/hDICiUr1d1DM0n8h7CeuKv9R1DrPbE9jbe
+mesiG/5AzrhgtmKciW8wC0g5U4YDB6XxYkv9PVaMX/dOePKIbk7vDXNFdG/fJWH
QG6qLVMi7iSuixyQ7wVhj+sSMGHgnINLMR0gQ12qM0Vsal1/cGHQ8x2DGhi160Vg
lOGchC/5x6ApL4TlLdtMwQstm9q1adNaHQqVKxAp3Ld54zsNEnsz42vIE4I4FXjy
13OP/soZ+pNLrmNOzvR8WKJfvnSOAAe3RJj1QlQifViV+PAhACWKfvRP6tu3aYTU
0UxJakufAaZH6BH9FThzPkkLqm+u624LIqNN/tmwA7o1CjnsR8paA/st0m5Et/qi
PDw3u/lGvdvRDc98KwBayPkMpB0VN1xZ9ZT72ftNVTbOxzjPmI8rlnw8kK5UVMD3
6LrBIndQSU8cC6wEDR8z9+6XfBXwN9xoVj6gfbzz8mkauh2qVWlppO+zq9QBMnyC
uy//GI5YUiG9LpPt67uGsf/P8lCFG5ZfoXxuf9GE/UHybrGBVVHocKL7JAanh/6v
oGddktVQetkBytYLXEcnE0bTIHB+hdaDWykuRxM0pa70VG2JbXbK/RG6yV4EH0JF
EV3rJSIiOxwoRd9N20jnLNuXNjr1Je4cYlUEln7uhbOWGFoHLRHm7p+LSB9/ZYlL
qPcMbc0v0GZEc1LP7Jo3gxb/hJpD8W3WXlGioK8yhgwxSJwlolFIdQKfB+SwtzBA
SQUaW+AmVGp+WuxQzheJJPWkxlfJRcThwMXTQGVBZR/WF1zFCmiuF8aHMho/42zP
FUNN2S1hVyMKWv6a9mIlfZ6RtO1ths38Ryz2s3OOwvXqsGuKDA4BSlCn6TmvqupP
OIVz0Ij/zg9mTRGdt9NEZNVRik42mXPa4gU1YSW+10NWotOYK7BmxJdYCYJh4iHa
bJ64WiZ3PGgDT5G02oxTLnIHY32lBmmTVyMcp63zOnL8fGQkG2RzO8vT6zRtXCdc
Ke0JoxFwuFJcXTlv7X4uZK+ZwpOgDAijpYfYFjS7rX6fvxSg1Fz971mfT1hfx75b
s9Et3c/XSi18fqI2zc4w6cBWmOMNCfHe9TCxHe8+jyF84YUH2EQYAqPig2UuMuT4
xlrrPqfDbR8TYa7QJ/mxwam0DwDgOY2xtmQWTbn9D7Sr16T4b6Gae0o7u7ZQYN57
g1AHCcnV2OCoN0SyjEOXmrwnFZ1QdRw7w/eYJ0uxSslAfTD4nbydsBf5x0xfxlc/
Be1rUNZKo7476pZWbkD2hg7tTZxzQBDa89uXIcr+S8AMd5f6Jy1/aS0FlBjGc2B3
DeN2V2O79W+6BUR6yOAZlcRH8vogJxdCnn4o0WsNWzmsI6Uehy5AOHULmlEsY51z
yeKZ0bCx9Um+3mdpGWzoiGwhjyxu5dZDBoYM6BBaxqewAa5Si6vbeFp/pNwkDHyb
ZWqFwR3+rQbGEeEIDXudgE9fEJVe+1QJll3NGnXMRt9p0tojVb3ztGoNn9aGKPNT
QgpndIzXiLQr+fBxj9+APwLyIcZKTxQ6iaHReYo++PUr1fcPrbNQS3we/Fn+wMTF
8i2c4uZTJpeVNI5TnSRjUxpquRi0rQGmaVpGOrBysHgIGlasaVliM+RQEIFbc/Qv
E0IkGxfzY57NyBT3UUSfSfqLxcDXwxH/C+0OnDXq0IVogbII33jdfCFFVYFtIEqO
eWR0jcOc1nLNPp9j+lY040Hfj1x9/6jB36UJI3XxD22Ywd6SgzmXUhnW6Ith2nRS
ISWVW+WQyG7BWIELCn8jG/Ae0as7XP18pa7E87BXgFIMe6Yw44Jo+vjbFvEX3nh9
3r4YhEv1nYOiaCsagc8SwQK5J1LcZIObKkgD3gdtKIKfNBpQb9OKB0Hk5p6Jigb6
6GI+VwOTt5XbU2XmI37v28TS6NmVoXnfC/sn0ColUbzWdoaOOPuOJbt3NVgtBbdp
aD0icSDKGpzR+C6BBIHDQtmRSWIhtX/rae+P85H3U9XlhFkod7GrQw8kjo0azB3z
4M0/mhkNi2VoeRsNbqnTVwXZRZRJamzDQfaCzNu9n9w2A1NIyGzbqMH8GGffd2q1
EWvhl3j/JeXxw288kYq/2ZO4yI9aML5tHV3TaxegkRdKtPSYhAdL8lb6TK1CMloX
nrIcozsWAxZ0SpA7vxHnLK5hiPbYwdQnQnomoKGDBrW0bErd2BzmV9MGoqEBVrtN
LNVyNJdQU2fjWjCUlQoDzAToDlqFNKSbNagfoHFtLSom6Ks7SZWlihid+J9OcpEb
8rBTwec4FDMzUsH/8HrqKTZN84kzTWPEwnv2fSS5pKV3ndhMWCZvMjpDGKoCLyOL
TeYY3hja+NsdWk5PSVUAJhHp/5SB84HqcOF7nXd3LtloCYMmaqlW6l5jBt7Y+ZXK
0W0LrgYOgJEcTcSk62sh+FBwsBXUOMvhCiOqlekzVgrJRtB/TeXsDHaMHmRujgyi
wcdzzVKh1bg5uZoLYNrK8q2e+16hnwfmIJJlfdJqXVxbCfM9is8KdkM82iWy3GNN
wxOmBir1e6JNTo78HDMVFy0EKOtwcxxPweD/+wBFAFW8ElJ2wY/XFzzlMS3aKEER
rw0BkGNxL2PDSvci9YBKDcyb0N2WdbvbQJxTO5HaOFRZvMZ28Kt/VHY/mESHn/y4
oL6oA+f9DSPurjjsedI+hS4G4rOUN8GATv3YlXp5rpc8ZtQobRLK46LqgO7li+5F
wlj8yXFlc79oDmB83O9OJLbPISppYZeIC/oqmOSnYiGZ6Du09LueEbsBZFFV+YGV
BDg68Zcb+4dsTkiYP1PcK4goXtFhvvl/Rltw49eLQiuihJCvrQMtN1bpIkn/7qFb
NeGblgpm6ndVyii/ePNLtfpc5eJy1SyvP3HmohCxpDqLLHmL3oFjpLMEaA2C7Upg
D7KGl6oMvuPK8b3qXLZXWyfhFouGCOgV5NtIFmbPNMPpZu0vT9MoUbBcA9EeN2gV
+S5mrSYBHSimAkfxIPhRDtOkTFIJ63Z75hMOKpbBrMdCC8jYUoyC5PbZNlXMjgfQ
KvIP9mWR2F0P7itnN4tV3GN08hHorlVLLDjrfegQ4x/5wyfLKVg9z8wLHYjpYc6P
yIrKfqPsAsXVawx6FZiUmbXIoWBpM68cy+Iei08xMx0SFlYaqfu5q0KL0TSI4Cwd
FbKn/NraPtJbqzJKBnZ7EumiHv98inWmzLjytGHBObTLep8z+dHe8Os0LMUWl/Sh
nccqk+HAbAwUDeyKMq2M2RGWftrw8DTWL+UM1zySwcZ9e/vTWyXeY+MLmQqonPHQ
OqfuJZ6uUH9q+adHPtHyCQDmNYDuIHcJUfQeDckJfytKIfGNb+LsjtSppnAoA2Pa
qNWvjf6xEJ3dmzcM9cu3NT2lxTaXLUnqsLPp1e7ezWeM4vRKkjkicVjqfYXPD94y
6gZ5S4hPe1noFmyk41M0zTa+gx7vXYql8Ofjr5Zez3jUf7YskxkF2AvBT2KDj5G1
QeIH44VA/ZRv4/zFH8CNHioFcw7wo8xZD1JrFJvJgwWenLFWgE9xdQxI/DDNiERG
6pUNsIo/zKJIfOzMNua2xyf6l+ywJI+OQhaVp0ovrR+aO8VSYEGr9KyXzotGy9B2
IiPBbIGfpEoTauJJNoYS+tc4ADq2HKfNfMk07/y2Fq/c7D9bjZbryKbaaq3qzYhS
HE+9+S7f42a3dgZU7X3oP02av4dZ88tL6xdEgHkldpDkP4RJiTWaRr4WLqQz5SZQ
wR5Jc/Psohgg1UxcV0itARst97UAmNoGO3kGzFqoencWDOfaGXL0DObzLt5ZPvuz
Dl6tfnxIC521jQuxCafksON5dsMnBq627+N5H73j0C8YhKJOEWvldshrZzNf9Oxf
E4kmXiDX+wbPZkHTxizSBMNc7oX7p4W2sN49Cc/yAi9nZ+Q+cdO+mZP4D9ZzEgFR
ESw1K0n9PcWrAeGWTJXHxoc1k2ivhVrMkVPjN5ub7cjq5Z0UfFtxUGHDpmwoPKVm
SiHuEAu8Jk0/uQP+DpaDNPmuVN4upWmqvHCnrOWp8+kNbHOYSd2C3pzg/jyCi/4P
8nlx5W9Dur6zeVPITST1BSFx7a9sO9x39J+mPntlI5Hopta0tA7FulrZyUeNhWbE
Vl2xV3DWdBICag27ICl4SVHWToAXWLLw+bCiAAXPoeuTdigvMS6ozpATwMlsd5TD
2pl4hld/qMVGEHdnb/FYi36pM4zRlw7qqz+2KBBV9HE=
>>>>>>> main
`protect end_protected