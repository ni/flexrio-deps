`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23952 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpupmJ1IlVmAI52F7eUhB0KOQzGYVUX+dUm6aHP113Xzeq
rlKo/9sJH9VsDiAJ9QN7MxHhoUIfy/bPIsgg4NcQSh1VytK9pXnRRpJPeJU6n7iI
QPJfRRLU3oE5yG2/BpP+E70/jOKnYJnvyV8Bc+B06aujXmmNNVhJvL8TQTBqIVaP
0bwgL5uB9dcPc1JDJVrPYshomZvwlAaDDuw7MwEUP/T1G9GtCglbXtR2LkuJ5lKA
90p9UcmuFvNbeelOijGEyD8boyXMCn1EzSrr/Fnm3a6ZG7Ealff94JBZdEb/C8jH
PXpSmWeOMqK1t7notc6r6HJILIZ77XVzIiVY0O6UicGMTyvlcm64raKVBv2gFWS2
5IOPSDgXfRkX7/qR5Fu89bofjV9FfPLX2V8tW8KTTPHA/+7zZ2NK4XnFdmJl+952
mDwXkCvET9IgSrnO1Xd5w/hC3UYVgxCPJof47c1jJSe3KQ9pGxwe5Q2RuZLzfi+V
1fs3ua+kDjqP3f1ijJ74DzcbBFLWVuQY1CvF2DT0cakvo5QNBy9W225KXrvwGisO
mf0AFy3rrKppSnCyfwGboVGXN5fEdLkZjeoJYP1Gh81RtE0mfKcIhSYtkTTmUT5O
NkdHjxgoUgAkGmp/Cjn0elinHJrZWw1NDZEz6BE+Ko7+wvClTO8jxjr2aWDvXKnG
8K2kPSEr3qx4Tm4kMs/BaCxnOP7bq5xOQChK8DEK/CsD1MSMTndrfD7i6cpoHGNa
cArQZ6Uv4qLdcGxm4MRKCAYjHFKqAkoS2WxaMpjQv7ACFIE5j4nphw6tfL6TSM8s
LWWjYiJvS3u6M+Ph5gyfEp9AseOmjNNlM2UvO6/weHvFCF4TfKv4eDObS5ID0dOj
YsSkzeWni0HOSc5Tl+Uo2QokSU/NrgJwzAUWfz2nO4LlORcKpZwnM6J8uTBRvzgy
i+ybos+cVb650PGsf+h/JZJaqrc42YNsT/HZDNU5Y+DHYz3yFaBemh82IBn0u9fW
qcreWvaIhPVP24eUxJEENb9Z71RVWYaHqPppr9prjEQO8xBZqqt5kNJkb/faawcp
6uOCGKBXLsIOhNrgSjM4em5W6YDb5s/Euwf+IuDb50q0wVg7WRFF4jx0FetjGvRR
s+nHeHIU/eeLNJGoiLrcetoXbjMDT3TrkL+Mx8sv4bhRcezQVaH4NRjaEG/EfY7J
xrMtqaNqbH3x2oLUw8bB4wBkIb9HozrFXeTzp6o2NQKxlNMQ5l4ghUUhB9VJ/SjB
9Ef3Sc3QYrKKs9LNp2IrFJeWziO345zQtT7GKr2X/A5IVdJCJdy+kWL7eFjYc1xK
nbGp/MWmDGPhKaDen7y946mYZJ/26l6Bvme+qct01VHrhJfPFMxzuTm4OQ64PEjl
3XfUEyWIcKUok+fw6+8ES6LJEeRZgzs+y5OFO/DC8BIEYpLMK9Zrn6gTcr4mHNM5
HUYzf3jF4MCtCJO34dQln00aJhHPTCWUuLXHGCdT7jHlnohQJ+sZD51C/ZJ9w/Rm
82la73pshLDzgKu1qQrOF7La4Y8S0+elQgdanHU12N0D/yzUt5m0MPfgZef1Qnrq
TBoGmk7LjLciAd+stFRSCxKKDvR7TASC8MOyCBocWJhh0p8zHrS/GQEan90cJ1fQ
aLGutfH6oUTukOJmvQmZsJdR5NLsqUftYQAvMkpobxuRk05/To8EnGTIhrdobcfJ
17JOd9HmzOy5qgWYhlp3lbJySKywqqeEJ71032f97gdRJPRX4vAm8IfZb/u4R/qo
zwQ000MGMmuFfZAAkoRTf8b0qrJ7r/XcsY+YakypUxrbFnb/BryZGem/eesYITgP
cQS60o+zdRrC/l39DEfeY2rmNZG66aXPQJOYqHdC/RqNp+nX0/74thVaqarNZQex
ixBnkWzyanzwF2JqmeJAhvWDLZKcwjsdi6YyBpnwicgRjmQMgNn40t1V00FOTBfe
JyBaFONQiDkNwQ947q3toj6TRotIjifvMzxDtttJEadEegTc49VcGtDEm9XvyCHo
5nRUh/mjqe4ZFvv05AdtQ0N1r+ZaQYRG1cNhWCvPYazA+45QnEcsqH5xGte/oBAo
tdZioswSi4rodAwK1529lXRcBB0QRoJsJEtzfwBjhdaK+IvDTPgkzJXdouZcItOy
iF22Zm5WBLzJP7aEKxRRflVlMYSzRfQIvW7e+SoJNKVMRI/w8TI4mFT3xvyx90RV
36za4fGO/z+Jr1KLD87/64pRpeTM6Parv+DpL/x3cIubJqLG4xUhDOHJzs+FoxRj
k0Q+nC1Nr2vUZrwMG9EMxZu2ioNdCPUVT7s+8mAsRlDPcASgrCnwLI6FaKcIeKyv
x+gFxi5PYXYY2oNs1FTAjx7AHwSpbzqG3HQhvasojcX5jrl6hA9MjMYFia2dA8iG
wBntc1oVfbLXGXJtotRvgaKAvA7xXechwydCsHt69PhaASSWRMOqLRc0E3j42AEg
BybnZp1JANL4FVb8MGAFQaprQ9AXX72focGzf/FjzniZghayFe0NugiNOvmuN6YH
qvn4uLBfQVIj3veLRkPigVh6tchKOzvJj8vVAPpzMmHwxq8Tcn0p/5UFUsNcGUrS
jbJX1Eokp3A3Y899iEJj8HV5gPyPTh1PerVJnKZqJHPqptvQ1K/6fgYg4hWlilrL
RQAOBXRdmg795fpMzHHaW+PuEQqN4azNodZnrXDKlvPwXfmq+tXNcDdnUVUirIKB
ZuwilUJbmAdJqhAla207hqQRKXsSGaAZE/Zr5kRSILLF1HdR3+NE2wC9DoKzOgiR
J4i0Vtq0gla+BbgChOI0O8BpZAEB+04TkLmCODKfoqe93sa7JFblAdUmOm2oRY8V
J6FM/MVOMUxEhv0Nrrns/oOBQo71FMrl+Mq4yRX4HeZNxKBpXy9F90W3C853gZnb
FeTX6wkdvE9SbzfFNCzkD7FNdAzS/FXsHate184b0dt5xUWd0bKp3ypE/OpGANPp
DxSNoDnhvXFaExtmowsSAKG2+9UrYqvc6SgeylfZfmrXeLrLtX8m8ciiZNnqG+3T
s8Kolr/o7s1n33iNusXNGj9Ub0k9fk16vvfyKFFFJEOP2jgp40c2ytNfB4+KbQk/
R8cCtn+fQvFj07SXC1z82N8bDj39Orq3bM+P5TxIUDW+dJDgQ4tCXfDOy5TmXsfn
FG2VTJ6snoaaiIcmGXzXSAH0eKm/yWSVhyMIRFdUjaM57r4b8HyIllAz4Kz/PX57
v2uQV4kusxdr8W4Tzl3rqRUFX0KTk6+3w5hCOaqLAQ6S74RrpQRp5LLWpzSt6bvR
+logR/1u49oeRzqNIreSPtYcGJezJYvu8dQ63F47v3gFd8FiqVpui8bh9UYlGoOp
hQSqVvqoBogWXcim2cQD78S5q2dcKOw67Ev0bq+M9oQWqGujwOXoy6wyRRNJ7Pq1
Ou1YYSjyUhOegJh1q52IlV+2DAjwfNZhsawXkPIwLV8UF6jEk6tlm+Rc3lak2L+X
cnRnz54CXLMngrsJcGF496fFSFZ1uBJYphQm5avDaOHoKwKevxg5bAorjLC+VE1O
tHVPSBH9SSt0T5E4DvUIEndop8wEgKQMzzl6HcCUee68V2UvJFF0C4JRrzXSANam
ffoKH+HNt/jliQ7Hq9GG1c71vHksWHGaCoyW4zl5X3C/+oDOehqQ/eJo3Vkn+PoA
4l1dSCcTAPFMa6+ld0M2EPZ1vwBfDICq2oF4RqqufFS5swzVXg+QNM+Mlk0AsJ3j
PSPrUbhQ1NB/K1PKuI59ilz3dlvzuUQyPrf33E0+jiDMI8ZeUUyl2KZw9Se9p56w
VUWOTn3fGZOmHre8GIe0Co0zJKq01eI8nXwWKI0wnBm+3vKbwu3Afxpc3faXk+TB
3F3/dz0ff91VI+8w5EWsu4OL1A+LxscYuglonJ6yYiwiEJx5prOviOnN4V3jmXOf
1LNCbFYLhBZNof+uXXgXJGgcn2qvwCPOaksE0oZK8OhLya/gWGDXhJHwM/ReEJal
OllDp6NUD1STmmA/EyeY8EWiBjARy3pX27l0HRUqsx3V1l3UB8GuY2eUfeRZNUBU
Dj7Eyc/bA6Jb419JFh/zzSsioLTeiyh9RVqpHN2akXaM8qyEGQdX/T+ZZNM947Sq
7LCE2vb9qLMooUaUpjrXW7tBtTOSCTnhVZXhFsYZiY6OAFw4O3Epiy7ukoStOauM
tiIIO36ir6jtDxwlGwfjApYnVgrXbqTDBxE6ULB5onQkR4Ierp1VqDUe+iZdfgSX
SYKbGVSPw9zTpb+93igz8BBEya0JkRQbEm5jq55gBE2tstNTInD/mhjwVJ7hfjbF
gB7q9lgTs65ox5q0d0WEUH/ZQibDndbAO9Z9lylq15JS+OchOmjCMZdNF/f9vEMP
iV928kS/aVBq1ehPmE8RP4Q1ElX8wtDkHBYnl0zxip89zHGAtDxe8rutGpRrojPI
Cb85mPpue7Xf0j9mFvbqBqgRVWVuDLow23xLBeqi8LXhN8uSgL/rVl1M+9LOSbw5
gRl8LffPYxHN+0McnC6B2yGnV03HYOUjAGWQZcfnSSIQ5a0fk/aurNtZdrv9O6MV
z8SH27q7DMmXtCEVWsBjgu6ClgJhhdJ47qIWC5duq4ZW9bH+YUWb2EDkNRshbXNg
UD1yh39ctv/kA42TMLGdKUg7GD0xeRz/CsDtyjBu3IjY+3CpNhHa6QxqGwQ6DDNd
x9ToNyTB1X++FLgb/9KKwk11cnFPuOtrhfcu5lu4p1oyg5zQQOdSMSIHxibsRQed
rfozrPElBdPXXHopeLHciVp+MAXpU/ncbmk4hSw1BH+nJdxa+Wsvx13XkPKt3/oj
CfuCB+Hvji806IEkXVu+/Xn9F7qml125cgGmZaKSLEK+nwY1cRX2PcIVprp6JDPO
KZgCMCblj6f0nReD0oNlRpEwKhennlEXN7tJ/kfg30oT7CJfHWqOv94d3GwOFFdw
IW3xXKEamIakV1isq7aMGzshNNliaVwwBRftqEjxEzP7eNDwpWTovEy4N90Vrl+s
tBMumY5Omimoz45+AoF7HgU0nF4WctATujhsyH0CEoTZVIJ/CkyRe7CXlwc9Olyj
VlLnq3x+w/4pELbD8R++b1/8hvxz8idt/Jb6UXwu+KwoIDw3wzI4i3Wzx/7VrZ36
Bq/OB8LthCYKv70B8SqBCJNNOI0fCwsiGQPoOGwAPOQByAcEQ2GPltUljc0YUwze
oYECnZlqogXgOZhlVjngiDa5L8pYZorlHtgzossgAOomqE5kG9+NCS2a8A3/qgjQ
N6Zbhf7XZ3J8k5KH8feH0WwaIWX3xiekfRsLGz38BY7ZpuzSlO93ayqXNz07Puaz
QmDtll60nOn8njrO5j/F4K2oJAPNmz0+IbwzOq2mnMpiAjXlUa+Q6c81gEwumLdy
upIegyandUEFTQmAdRNEe4Gxh3pYfttRbCBdp4FqKScHFuenM6ZjHB1+yUnl4Pyt
7pDukXyeu/oiSxIHuj0pzS+yJ40/ABf4QtvwG2zQj1Dl9+mWy6C/9+ngGlUFjofF
ynAc9XaqVkpazi5ILeHVviwhxZNIO4LDcsstGAjPVj5E030UkWZzO4zjOLcnAQmL
CqdNPmIt2j3xqoK6zdYEs+8ZMEkFPFhkSUbbEQU+5byIfJObZ5c3Uq9ErWyGM6LU
7cJFBjBPUJZai3DULAQ6jYj95uTjiuBowZ1qvZew7q0ILSqH1Goewju3Ch3W6dk+
lj7L3GeAYfgIL0WvT+zLj0FNfVdWalPI0FJ+XGGKzcb/teBZESQh2I8LoxPfdSd9
itk1C6X9p2OGhRs1PcSEjibTDBQICgUPWNB7u44N8JN4Oi/T/0N/yMSMWfCoEIzV
1r/taFrO4af0yllcwq1bIc6bonyJpF/4flDPT3UvCRMuwv308uYcbWYHWIXl2MsL
2fhl/yl8OtIVXuUjYaoqoxcF+Z2rYOXOknOUjgXCgOKOF5tgdWkG0a9T/mZyCyze
dYssmleJHQdDEb3JWIiqq8j9C59znMpGAqAuqON5akm3jtNLIQ27ijfVTNINUFaF
RDHa55bCs6qG2NBFgvyYIamdDEuh47iTE4Dw4MRZxmHs9etAmbnC05Exr7/loZaN
8eiIWli+K0MbJnhOffbdOuL4EzhC+5laoflECg3f7S9trJe35/L+ldxe6YkhGAIL
WtnXrs7dNzk097bENvxaKWU9jDdaMIVZkRfyhx5wZJDj9LZbaDToKePbjLnlf7Dl
PdpRIAlXac470dBjODEj8RxoAo8UU5gqeiHgvS8xYaOt+nRbUZ5efcMiCJfdBGPk
TA+ANI5CBYdwYeAVrxtWVZ2N2FJvappZTAEJDeewJsoJdu6dtUNbJaxCGhojX3Bl
UTLz1cq8jLKHUH2uayqlDNFU92ZjUqAiGyoQInUbJvsvS2uJCEbGrmVDJNv90Y0E
9f5X7C0ftwGWiB1h8avwH/P2eewREK/knnaW8C3ODX+EnpkXfnCjj+ABWVLuxLnA
alaVFa0AchQTq18yqOrvm5rVtpkin2CpKeqzIxZnMadB1cFtoZKGoVgsg+PyJWwo
B2V4TJ02sQLSpQDcNfC2b2/svDzJttH5sy+GgGl6x4Z+Sxo+n813U+qtNqUq7He8
t+m2485+yYnllY9Qu2p4NWuOQokBhHpPNNc9GKb4keglw7d2yip5bs9V8a4vevCC
VQ4A1vKv6O+La3uGgDrGWdfG2hFp9jVwYHpJ4mpsED7QAduFUaiXR3RIjv+PSAKr
EYG4VpU7tonlgTfcMUUafCmlVukuG+KW+TAZa3nFhpoNQoC4ML8S1+vo8KanBbTF
uPhnSQith8/cYUf9VpVNppgeyhyEiZNjD7RFYxYcPRL33UpKc+eqpBJCMILv/sfJ
39X4igHZlWkhus/3nM6mtL/N1tNi7x2gdz81LoTsVHIat19S/A1i1sI4igBfwNzD
UqzFrCvOubo0BQ7xxsXekTB45AAltdJEdFkdVnQurtt+CLlpf8l7dxbtq5W7JKb7
mDZxA07w/roYkNP0lieUM174xGn5OvyY3jTv/VuOeK7OesD46g/XQO/ZuKuutzNj
Som/uIq/v+edk3COgOhuO2ca6mzfK+Kb1yq19OsjGmuKiTWmb/15zbUXm67HH/TR
EmixOgAuz9CUB70PCV7scSLp6EWdmiSN58bD1UlVM8NZrdrKGv0Z2oourBPk9A0H
7f+zaHa4Qxep2AP8Xmrr1fGRN8/wHZQ9VRTuYdyB6PWK5Z4mu+MWQluKUQu0Nrmh
2z3TblD1MTC+VQRJeyGBqOxo+nnv8Q+XHPlCYRTRHAkvqUsbwr12Lh0ySTZNWSEw
qUoWLno2KLMYUmwCuwhUr7Et0588PeRl58uLpNPXnenvPTbp2xn0EdSIAE/3C1hP
XdPbS+9SbQwlSP/3q/tZMyXnzNUPDmnjIiRiF8TcoYfsSlQmyZInGMD2q1d2Bb5Z
KNqJS9dMdaGxxRWPmmMk1m4KCAjEjFCvtKhJ5QL+DfukPElnFdc8nJks4qBWgvif
bVabg/CZyMLGzTbK1XVabsEx5O6YD8wEJD2/0rnhnyVrk0qBW3qHfzUuvnc3JgfI
mbKsVwQcVKSBAO3HpBY93N0WHztHglDeuvqo8FGRNfYZ1WGBqtSSdgzW1XKt6x0z
Li1vw5DZ8wYR8FjNUj2r4ymY6bumazmA59ibLm+KtCbwtRPTYJFNcp4vNNhHfVXR
u2aCtTHr2vMs3yttUX3zDipqmC6mV95c0o3IQqPoJ4C/zfxzRQJ6MIHj80jLX1ds
y3+WEpyl6HKFhgtYoFDXwwnjSEufN2YwMtGdLCeGkI3XKO/Li8KtmQMFzW+K768c
juwBnGmqfQ9m6+Rh1UOQKqlTVaKQT/MDc2cOZfueYxFFIdW6IK5ON903a6iZXHRq
1x7oM4b0F9cPNuPWu0yr+m2odAdY7BzIiA7k/IslkbhltiftTHkzzVynRBbmu8B7
LupB1OPDsJPcVO5zoDnSCsbacqfniYLHZfLoeTIDBWLO5+QUjc21IAcEqv3AAG3I
sm6zO9OYVGxLmd3R74VOU8UJCjY9fyRQ04Yf0VABhn8QxRA4+tH2+ooryK/EsiM0
OXGLctUaMFAlp+95K0qkQ+R6Opp1YyBTy0PMpxp7k2NjOvKAC+fVqgcnd/S1x4Vp
Do1DXhpismqE/2PmvPjsIj1xVxNy1Wf/BAsLtrXcfyS1JI7MLKGSwrZGN9o4Cv3F
PH3H9PzMXTDE1uWs2UByY0zXPPUKIX8QkvY17icsjbCuTNcWRmEI/s/LnjHILS7B
W8PokD6pTANhON/nr190z3qlNt5H4sWD9gYy8RdHXwmT+Z8u6tTuEIhCGalIJW8E
6/f8j+hgFwQn1Dg84cC/Fp5KP/HxJ7apjAVaBQX3jYaRkxvawiU9NqIuTZe9/biU
tAPRTpNSfOp7X35h7XuQbLa/YTx6lgVziA6QTUNhjAPo8KD+4fPWAKnEFhXKYr9P
1s+Bj8GmzVP6Qedj+PWb4iDBnfOtMmg6wJdLxIBtcrPpxsvbq/re5fEO3zPxW9Sw
IMupfefVa54jtE2Hrp0XjO3915ziaiSU1K7SdMO+/3M4eahWc0QHcdUOZRndtSue
t2Wh4xu1B+tHIE8xmXgv1rewX12VuWp/4P9WxfgAXy8o0fRiLOGZHmxJGtFFEiSm
fpjraYAC1AYTla/LcPwXIFQB0q/Hrh1KJBBon+qlzuOCfU04E0Cr1puUAPQVMUeE
d/B0vsD5hBSyCWg9OyHRzcPoTpQ24TEQ4ZAnhGstk1/EOw9e9MEotVwRnPAJbQKY
b4RQD7OsKJvembXEP/cx8ZbmfWEpFUbj1lyNm+kQ4voqrhyhtSi1TNB9L5OaR3tn
gmH0pfTDIcAs7hHebFk9XE0glBL8nJK97f+LQmnQexFN1CulhkQXd3dYSwsM6igE
AYdy520U0JBoaQlY9FRWi1n4xdAQRtZcmfjiylvMah2vlztKE19bYcV8irVabuZO
I1rMmTG0QUdk3Y26GDrFEajnSVJWgbJBt+umwMmkKRxmljsBFLApLDSxRm9yoDvO
kGXw8sBZpqTRapBE3s3shzQ7pPAjRb1p/E1qv8mQ2ItaVrd5FOcRHrJe8hXLANJC
zd27KHxc/5TE2X/z8/JGkXs9J/w7DX8FXWdqoEnAfgLF81HRx8jUZHZOjsPOFycT
ogTnYEdedWKKkDuJCAWprr+6IoVo+WzgIXzS6Vvt286Zp7aXMDAXvaJNV+r29t22
dONXsbzzOfzxsOO3+wxqtUx2AWcv2unnmFHvwVjm7MoEW5YFgdRFIwaY8sZcOr+J
PXmdqA93XZK+mm0lGZRrPImgzrOZCxg2waTz1v9V+js/tG2C2rdlT362H9O8Qz2R
QqkLJpOe8fZv+NKcbO5gWhuEq+Lr6erBhu+E4/okc1c9/qJT6S80BVe/r8pJkoaL
FcsM8P75jY7OUwSfDf2h0oBCk/94U390C4Vm6p7+GzgD+HrqndC7wAQBjhdubzDw
i4BZdO9QkeTN82ZitHpGtiXwCx+2gpK7xcAPyoLKPAZ5NtetxeGWNPD/mcsS8JYM
uEiyft2y39NI+MXPT3Bg2/10nBRrETGYXgZPiFv2PRlbDwF47zvp38rJXeIuCaRe
Z9S/F/ZfeuzW/iy1N1Zj3TgLz+HHgT8zmIAItyM/20MBHHS+pE/wjt3lcHH2XufW
MgEUE07QPyGyEbDJ382RiylTftonJF1R1OUZTIKYFCeqPJhZHUIYqO8cVHBUlHlE
Vitds2q4rS9LrmoUVsf3cpjcrWFqaq+3dIW3xwL4OW8sS7jXJXiwaqVPVy6gidUl
JXhInLIKcTdrvDkJc2yVHmUfmd7lMQBp7v2C05OFp9mH394/T5JoOYIwio31IneO
KOuDq1cH6lJnl7ilJeO2+XD9WCTuLmHzLAoJaVKyLWUKKBTDPo4ND6bHMeD2dhMB
JUkLJsaHKoy4ua/8bGmfTvHlMXXjylalA3N/ix8ADTS2Xyr+R98BOW6XzFDYvQqm
F09bg185drS+fHS3qf52RBWta8m6uSj0GinauQkwDjaBhSGlaqClQOjSygHQOVKB
9USklfVxGH8NVanHfjLYDkMKiS9nl/R50O6yysQGuQJ0/sBdVAmHP5wvbZjHBJoC
q8yjoC87wKLkJMHwQYGSIwyEIFamNmXe3CJjMVVx+IwOi4MW6Q0LNAMn4UDq1dlu
04Y3XNleUWKwwfZav2nnnFqc6rSqHHQaexAaM3ZCUDdB3QwJvUhB8nqj8J4nQmYp
kUDAuzrn+mJzu/1M5ySxqWk1RRB+JiUzSwRkNv/EYk/WBZZrh6fvhnio6CJ6x3aT
wgmhyHbszJjlV5DedhW8F/Fr6p7Ap7Yj1ozN75c5nlpk+nJLxI4+xYacoX7EdHlS
O0XxlHavmK5phCwbEC0pR4XfKxoYqYG2jbSvs2wneb5YhLVYv+lL1Tvw9M59aDdP
lpYzkrHIRiRUYjJISpd8ydglF4hgdXzMhr+BHGPDrLjEkP2NwkuZeQu+hCcG4E6P
S4Dru7xeNyM2+QQ3PdFdyluLatVN+bWKrQZWfzUpKoOGEyD6aLL5dqaTe/tQBo/2
SqI/iM2Bla474FVfZKMb267rhwhUmnYTGygqcuiezrhqsnpTB6dhjqVv9vH1bMaT
k2yrn/XheLhK++Cfe31Aoi+PhWe/Oqf9rhrRpMQqafnyKCY/QW/6lBSFfZgBg2Rf
WjunOgbDKMxu9Jl5qBLmqieBq/Tgg7NBQ/QawKUe2mpJREELYrolBven4kdx+pQd
SDxVP9Ja69c9KvSXbRLrONt3aFDUFe9AxaVBSslptv1QgY5z7kmDo7JgihpDfZUn
L73xMqZ9LY/jogOMVzwBJvWNVjL9tTtNg7THFCBBS8+DPylvr3oKRPhUv3PFDDJb
9z/aRzPwKO5Lm+tIyPWl5zL0yA1UlqxI/oi2JPrna9Kj2j5vpOx39paFn7eVV8uj
yQXP/A6KT0EWxpzud6JmB/9OHjz3SpHg5wgY7JpkDY+MqbfeW9ssLp5eNnWgMzIf
4v/RJ8p7J6/vTYnD3qLHC5BfFNPMaoQk6BX02Uns7EEGS3SI5cEuhii6i2ICupza
UhQ0lLy5g2RdPzL9WU/PuwSR5U1o/UzUhT3SqYPcBYpP+gagwVWTJCREPUwbeBnT
lYxwgLHl4pSxawB4YsXjymfItiogWhDKeHY2DTv8yZ/GgX/RDQ5BjvEnR7YlbmwJ
txxgzCl5HVV3Oee3/2Qx96NcRfd0qGoaGZAZt7FtYqrti5EFl7ENspSuXQ+y+EcD
F/fiTZLNXMDbOkLQz6nbaMY3JkdgdYG1JZqsd7f6ebeR9vo01YTBsEEVnsWs+VLP
lLuch6UuZL/v6GI6OcF+q/R4k8apoF5CgqPyAuZYh2tJm9PGVX5UfTpXQIJpS2LG
nfUqO7x5LNelJ66C7GCdnk4x4RAbrHHhP2rrfwzwZ60SY+yegN7a4VpK1ad2xIZR
4jmjTTGhbtmn1d4JhlqBK90pIufe2lP6MjylStVMZVNw4E7PeppoWgmfVv4o2oX+
zQDOitdrDlBt52C0lRaQTH8/sz53zibgAG++g7bRAMviCGe4nnqbaf1SGQQWwGrH
lX471xckEjBn803ymtVmtfrFIf6LqAMhjUZwchcyy+gQI6LV1avYEDodHc4GbJV3
BNLSHp6zwHpH+s9c5i+gv+w1twVTywrUaa/7tssM5ZjPxSp50AewFTtT2QgGYgCt
FPqThc1wqoOmeuPWcsb3qLpIsTmB4uplL2MPJ3ty7Tka20nD767tjN4w3lXpNATf
8h5Q7uSi9lT8qVJ3Ad52yXNihhgSZz6CPRZ9vabnFkgV/aSljmWuyhJ1Pira3TEM
imiO61uZY881Avj2jqJ5kHOSjzy1vxA1K24HSmETMj1xDuGZUUvvF9Ml+pQeSXlO
mao7DA3ygy9IbOwOyYlU9u5a9QjsnFXsP3eDz3d3KR7C/2hTD7yq/mrinLufzbrN
I45Sf2FeKWE2y5eYSvWQIu4TT3ALXvvhUUZbkahLB9KkG6xUkNXd61/n3DRD/2A/
Ik9QCKy6TUvfAevAmYjGqAm2KypG9ykgbyWu3PdVe5M4ocEd+GafRt7E+N8lD8JC
ujGkVZ+BvLfMj2fE9D+JY321JItwxTcimhETo/nNjS+qfEDHGT90CK9jzsOfAyBA
LzVSovJUIJhv2whU7IBunWS8vnVdPQkhvU3TUFirjrJjmq2Tm6CzG7fAKgmzgFKe
fK7k+VEoHTuiKFB2X1vk6b+qNEJPkcoCYEqDovzv+mBMRFxDu1TZyx/PjVKNIqou
z9wrUCSFDSjNSVU/xYDvQiFuPb2qvCZ4+t81JvaxuOPi1vzbPgNKRckHQYsKLvxa
LT0ghuCN5RBbGOeLaymC6PW+oJNz/KKhopJLsFoht9nZdLfQrV1J2nhxrQ4yKYk2
9nN5Q+wLvITxVSXVRr6etmFfRPU2B7yBV4apEJSgO3dm8KvgnfJkAIeDVb/u8Ejl
77vnZkLVV/AB1FBpBo3g0CxqIPdEUBn6HVj30EXZLWY4obC5/QNgNarPIx/hDWBd
Bjr/3izPMgK5A65NkYIKLS46ial+RWyzZOP2zZHXxURWClHzq/627oNvZ3qh817i
y0pz9D+rFhLc8oCom6jXSAE3N8OK2Gsl51TrfenyUyuOZ2lxYVIVKrmczhbOh3Lx
XJ8TosI9WJ9lsuSMdqbxC8YPtk5RtnPFx8Zgt0orWcrT6P5xVlUL4O6yQjFJDYVk
bVswlgpZWns8YDgIS5w/AnWK5fNykl+jVkcvlweLBGy/jJxBdV2NsFMs1hMmyE3a
hxTfDBtQ0/RUDerboc3YSnac5P9CJSghrKCIfSLo5XP2XmFfI60kMhClkbSxNFoQ
wEF5S2bRwJO+HYC94csoSXBOxkPvxMVAp3pCREL/GNSnXdLrsZf37jcVV/+llTuO
cVrsMen0xVVqaFPgvyb1KgIrRWGdQyWDdEGUgN5b4IkxpQ8kp9kxD+fv+4BnETc5
FhWzXiwc3qmEVJNxrMH3dEL0EDllUmfNH9c8yb5ClKqDxgXTYPbj5MgpQoAyll49
7SrsHXap1fO3bYv7fl9bF4mko1YnBi/NDLU7apL0Owit9utr6pnYBhlgZgKXcu0R
6vEbTncQB9li1mWW/PU/uSj5vLnyl0v9AJfdixJirt0KnTILsa4l1PTVYlDKg539
EFGvweJrUgudJRmg1kT6x+9/6QaTjGXCzzf2X2st4DUyIjKAhm+DhsRICG8bK2Rq
Fiabo3+ZJQxbRXlNnsl2L8gzsLZvEhbSb+b8zC37xYhClTWtKB2wpIN7o15ZCMWK
8sPxhNUPebvvzkCJYdNrSr6Z3FxE5QYYfw9j8kspyYSOp6Uiqq2PGaZhqKN22F5z
idt1LzR4N2GbiMG44VJPRJ5cDn0xbqaorK66VZx/NvCuDIysG9iylSsCSETMLN2+
DE2n5N0KXhlvnspQrUeKRBWCp9EJJA6SkAVq3AjLGiGOqqyA1647KOwJGVxhmWBX
ntCEtig7Rgzut61skarTDNHJ5FlTyUV8PerwtFGbjuEZaGe7oN6YzPrvpcPFeWTy
DVieUDSZAom44xBo8HdccX3ZXTvQ63S/PhVlIQtrlKL52Mc1SUSAVsKJoHx+sc7X
URebpw/1tmguc4sA6LirAoGDLhymuMbGmShP7nUp9T6bH4fllSNjrr03TqGsf5TB
CBg5FMcmlaK/DOBt73tlvvwOTbjiolyPWTr26kv4EhpLfo5RkMAF0I3HUk4ZOUQC
gQ/egmgF600eavbmRCwQLk/t0GpDWJLeztKdzgY5R89gAZAM0eBCDiiVjb0R58TS
N0inj9aJUrFSspTm5UPIzLztCDbsiR2YJzzTeYjC1T2Sep13137lT18NGK4HaqpC
AiC+a35r2tJU36vXmw0+bxch19PJ4EMFW1eaGP6SJfWvE4ls+tHd/N7GJS0bXO+l
GfXPRsmjNYES2vqfwddFnc8kpSkU5bAZklLyLFankN0on/CIVATb2qY9PvL97+C7
ANaOqMZagKdEMlYyJjvwSvi5iG6LzTCRNs9Dl10Xq/RGfno/N9mCP6x15+rR+AQ/
usBydY/xorf/iWWA75B+egiWIWzgG4J0Td3c23c8rFzeNulLDCbg/CePaszALiFh
uyNYrJgrM7esexmqW+iM88FUWGJ409GUXF1PXWa3bHKTmcUVD6XtCaWQ2V5NVemX
Cxvlui5KbdA9jMTVUq/F8LibweR43Iy+uTo9fKNR9fHHvCvkrflUphdH4IVi7V2w
pYABH0xPFkfkkjUUqq5CwVR1Knx43UVUwNHwD01jYsQKTBjp/R6DYMlWLIuhsPLO
tkPGlyvXSVY1SmBkDS8vA2wbyGF1kODJqCdVubfKe9uGZE7zPIKJYIYm98yUy/d9
f/j9LETVa6/xja5+jzK+Abdf25PU0NlJR1NBEjGKfb/e5f/llUc4S1dSDCa42TL0
5nGi06ZATgm3MEnBAW5J3e6rUix/Apun2lXGPWrht46u8KmMEeRUvTa4qJBWk5Nu
Vl+ZoIt05S09INjlnPbppsMCkPDK8tRJhCrm/IPOnYA7xSAcRa0vbAfY5LHJSvZV
E2HOJgpvY7Twl416Xqub1j+VDyS7ypRW94Fr8UjJLLTNtSD4GSktcN9zGn7wdY+v
dcH/Dyn7ihmecYHQwOnUqWo+LaJ3Z5kdT8hnet5JmxB312ZSJ+cjWCoqARCpYsKH
19jZmyQbpMOaJVtFziY6kkONoUpqLBfZ5XqW/hzwY2JAzX6uBQ/38cRC+EG7SwH4
1Md/gcBB1aDIdpdrdv9ERZrB3zCCzcdosFAWC840hQdFNyXtBLdaTt4aijqDBTNA
sP8CtRvl8KqoHH/cKMYX0r1cSC1ApPE4Z1gspunNgl6ixYC6yCC3M2joDyMmb1pR
Cdkadk7eOkjIxAMUxhginO7jQz/bPm1xGkQDtMmdyUVmySCzKyouQFQJ4uEQqLyM
Xmtpm/sD291QaaIvRNHjqqSI2rCBIO/h14g4YhCs0XWJ3iTGlTiqTAGW2yS4QSuX
2E31MgHPAcur1jMLJjFlKEI6LzkKrn6jdPeirSiN30DPdnb1Gf+VoEZBptOX/Gyj
TWScEh023rgWjcQGhHG+XgnpZ9/9v/bi67IKYreErWGU0PA/71U2PxbFvQ7TzmFw
9xtIkoqh5Y+OjuvVyiZjw+/SaP2rd99Rl7ggJcXvTy5aVKJrsmZkH5adjABF5hUZ
u6U2iPEaXN7dI5u3mjmahTwZyoCHgdJJZElLidDZIde9UYWevJtDVjTeWGtZTjpC
eCLxfMcl+AtLL+ImsUDfHZ4MGoDOYMmSlzpj/QBByBXlfkmJuloBWgJncSYNShmM
lN15JT6FNi4zlG1t+8E+Iv7ESbsZcr29q9SgeB4v07vrpHy5nQIXfoEEvPbmUDCe
BDh9Lz11V51pH3mIV5YVS99x36bFcY0K6TZvzbLN9UZQutrHrgu3fa4kcyseJCNz
XMyro5I3uGsu6e9kwTRHW1dkKo4wpEphYNOd1/xbepM5L7uGk/IrjW85Qt0+rDsX
voQ0e7v5CMaPrp/zQ2qh78Ug6svXYrVOlOfdwqh6FWh3V1lQDNOPzmJyQdBhkESI
ice/fA6mK8xSRTPfYp7KHBM4J1U63+J1VI0Hp+vmhmATBZfTUr2VWB126+qQzG5g
TOkUoF6ORe9UifC+qFRKKLOj2cz0XpSevROXt8oBjdex8QgHUQERJBQ9TYxTjOVm
kMskOcmNFVBqUPM88+MIrELRhKa+O1Z/Rmu49FWNyCIa2gLtY98aDWeCSN2y407j
RStaqMYuBEAcbMD2VKRlbkZPnZpvdhSZ5TFxzuTBepxdWoLBoyA0eYBKrWorTLml
jptOPrGA/qVuUFVKeC0Gf1497IFrY3ZTYEhqXV2Sn6P/c1SmZok6nBYEDcQEy0sS
skvVP9Lz0gri5On1y+2m4HCDlagQBXYdhe0S2b487KWGS0QuayRLWZQz9f9H5521
3UM/wpt/vGQdvWfdz9xBoxSItdcv9pUlLlWjBFnbGgUCGLTk2Sbcyshdw4ALLw65
zyfT3ES2FQyb37TW4J4Cj/Dzj0tI9EM7JdwBuWIctROZcJzzrC5a46wsyoZspWBp
qkrZ8NKTFHYDJ4z6sNiBX2bhOgzF+SNPasoGxAKEB4gx+scBrICTGmNlA+L2dIrP
GnahctV87uLmdKlxkkfwKoCTYfO3MAgAF+CLYzZSiSwKUgz3WpMzuQBDnW8J6GJr
/Xbj9Ovqkwgq2LdleG++AjC/qr139G6euAqrxu4Isku4j3LHB33DB9BcyPN0L+C2
od27VunqvtMRmmmfOYMKpRq7BKWV8LrD9c3IgAy7Wz1BwjCH5K51u5jrORDWFMcE
9+pp0R4R2QkJS3EHp3+z6Quy8Kv0kSXlCr1lpPBcmmKOqgSdy2JzplCecvGx1nga
odU1r9FEbWic7S9v/uSvsbF0ooL2oFsPRcgbnOmNc7+JC03uRMQWowCCYgBu8A1p
sDZr6q7kgfv6+fi+LEhpVf9y1t+lzhGEwzoWafVvW/ZHz3udQ6zq3qslAnlvMrD3
+YzyZhWixyuNz5cOXsyOYXnSYRzfMEle4/cEvSaqMa/ulRoJ1oxkzN9ocTDSVCHk
n87mtk9Xd6RbiVv+kybcijNvULDT9Ca6797+/QqEPSJIra0Mhs5XR3/Apy0CwJPq
kNTQjhMcc4McYZjowEgT920dU0K+EEEpciPc9CAX/vkoHAvZ+P4HS6BE13aSSTTq
jjwdXHBZGESqvlCkmQtevN7U1FqIdoPix/dIWHqMf1r+Vf4eztwlEkssAG/GRI2J
+HKpjToCKl02850n8dnx0RFhhTxAzf3ZpDEl+Y/aTcu1cxxCUVbL5EIsgshzm6wZ
ICdudmtc4iG8VECttbhF+GWu3Spf4lS8VB1fIO+q2JeaUCimQqbPX/XCetK6XAfe
V68pWPwvDj5n5UStFjuwZB5LFUOEu7vZZqaIGojnvTH73wQ1kwcuQH8xT+lXolHH
EjBCT6vClmp/Ehd+i2CAD1hkC8cbvG2KVlStF5Bz1Zge/dcl0yBD6m9ZD8/w8az3
ot+/K1Sc8+P0PpqWIomKE+0ald0c4X6QsaitFFHwtd9rl1+WlvpSKvvrEUjsaUaW
TGIaKcPPlwA18fyuRRnzpj4QMWW4TOJ5JoAkfdGKcNvPQhRzMTAutoZDdKoHn06w
cEhrPYmhzFTJCFd14YHnDTDXHZZAossmo2sGoJWYsK226XzJfBByrwsXJDt+20/F
n9xWbvB3E2XMswMLSsXv2tF8sFNsaI5VZ5GnUCXGNqvjpkKTiwozvl0Ehj7pmp7e
L+GCOqAKTcn+HMQW3aozQs7SmivRd2WcDAdnvEsPf1ccQP5d4deCE+EbvXkivSbD
QABxhFrsiSRKOGv2d2P/yk8+E8TdzJdM7b602O9OFxMRk61N4ulkDJukXK0gQyEp
ectYOMoyuG8reKBODUGZpwz1jIhFRQ7grhAWcQYWOwVpc+EHA2X3H2NJvgzzsHvJ
AfGaCLn9ZuVlp/yGtirjd5KspAaotS3/DZXW43r9BR2tTwZiaaq6VYtUFizeF6rb
usAbjk3hGbtyO1N0+khTxOkb2LJJoW73HlCIQmxilIadR28mVC1qymEaQlHYePCC
GSSPqH/88v1Gd0QJ9NHLBf8G2RHcV+938vOj3p4ikt5x6//pCYsKuW0tz3/7cCNs
XaSAEDLxsWVbu75+odjiF0x6+tDTVV15r1zBTT4fQvo42OntMd17BcOkHLJIyh6B
Ck6npfsQnRGY4L+jurcLYO5wgkvuDZpBO+MYSCXmHGysula37mqrzbBr8m7Dpygz
ZssVR2HzLI69pspUEm5qAw0kCcsQMA88VTHx2XzHLgCBEPVjulQmoV7+75Imtjne
OaAbieF7u25e2ibjeU2tpBGUoyRc/vLSkdmzws/zGsI6euaHSC5njQTJUli1pY9b
49nrsjodPLs/vu11TVEeUGcAYHnZGsqwu9J1Z9K2CM4azH6uHLYVF8/pYl6hroe1
rmjUxxsa+WwjksXPea6kSVeMsAnuicllV2hhSqCmabq+YI7vsgoRoViKTNwcwcNE
K55p/ASG56BTQKgiHu0xYJVc+zCFHrDTLN1mG6qa3wj6llGVuvRuKD/g13RGrZKz
OkByaJn8nJ7e5lma3UnjPk69xQB73wnmAjxxkJsjZydn3ka3kDkN4SBhPGZD/y/2
8uLygfTNbZheuP9+pUpHMv6QEAOLZXy9HQ12hKu7pv/XhXqcnvwAgb7IfW6bXQVK
F/SzqBDBjRqEMmcJ7VUj9aTxbTcV1WxTXOl7KAJkyrDlkcHgpJJ4bggmIN3VHdqc
PXbELzfN3/hwvP8NSEZ8WN/Y1fW2v0MnMvPfgmQ0LqIuSfo2WdWCQ1c9DKeeGv+w
aJXIucPllSme+EEB/7j9eJYX50X+bQQPzkp3QCF29t0daq1fkNX6RMWHU8G0gCbR
nTJe0xO/ykTSFBPxicrTIJxK/By3Zyp2PZKbg+TiuTF5NQVPtwbt5NNrjFkTxh/3
YSAeMvE9Ta3y6bLZO6Ocpyf2TcWV7OGDMSmkhKcmCWOkiEeeEwO3pi88Rjrfa61r
cthML77sOxSPpt5bKtuILIlZnd2OFkT2SBY/T5btyuyhUd+Gxc3yu7dk4RNx5LPU
cfBd26sMfhLi7k6igtt9KhNIk2YR8xNyCTH1XAPbmvgJaBosaFJQvYM5UepbcuIF
1MQPeVCSMTKkImXTF49QUzy39dBbfrbBsDu3IAnvCmff/7Ak9RLl/xiQICikZn5y
UsQGpSmLKciTTlv9Q752M1lQkkB0BLOw2zvYu3ojVRC7TpUOSVqCeWctwFrEbO7j
BGDDnca1LeEemg+foiYBJygdm21IbHHe8ykpgLtsRc5okGfWbjNaGgiCX9es//LH
sZ5DpmZupkaZwXJ/k/IYk5ZFhEEP+nl0eJnQGabtYsB42wEVtNbtfbsSqmxKKpfE
5gyPNSDHXcYgYZcsu/dxxxeD2eVikpnr5RgZHsjb7QtmpEZY1CANhMjft83sd6Cy
Ox4XORFUn1DeWZ+GOgF2edUMMuX+7bV1TphRiP4YO7tPuEEc7sDRNA9AhYhksTvN
giqdAhN5XzTDvt86jMFh9wTChBSf4Gg9DubghD7oX2kq51g3waI6OAs5Xb9VG8PJ
VVB3GL4wyQWhKBw+9HIUI0RQTxyU3uzPOJUvasnWn8eMbn1OVcgRuqGPX5hJckoW
9ezh1lVb6UyLEbXjtI0XkaPGUNV2E43qCHV663TwoZSyE6PRdg8LSgIdEA9PDIj8
92t2Ljt49Gqj0tfH52gTdamvP2M/4X0rSZbeOAlOByUYKBtmByJPk3qsWNzWhXtY
B7UyLRYNJ6ey7ptc1xs2Ki4/+2CvxW4oyVsrOJstpm1IeKRKimpTDHhH1OOdm/IK
+OKYNOUcyK1YohbOtyhpzvBKwwbnBMupuI1nFW8gah9U9vkX6MI3TEGH5YGk66IG
CbO8F7Eq2VRZypV8Kzo0vZh8QvbHAZnTcEIaC/BjLVcymDB0/fZZVeLx90xxA/jb
RQNA+w4DaK8EwhfhgYCT8ILtpXn9O59XdGfdxl9KVdgfEZyV0MsoHw2q1nqqQCtY
MOvKG5YF0cB5M606VYBXjitcBIfUq2slxUXje/uVSn+k6I+unoMmJMca1vxraI8P
K+oY6BdxhompvN8JG/Fh/ihr9M4tzSrAKooLjxzGcKPh+R+jW3fS4cQS9v4CtbNP
uIntSkhJgy87Qj9nZhZVOKNeO0yOXfsUwbUUek9e8hcMZUHIBICJGMdEOOTut+cp
4h0rnm2hVVH0T3AN7eOjPWmDOHsHzpI9HszYCD9saggdOn06Y/VEi3p0v+pCstZS
5pZZwUK1cooTIquSuQcNTou6wwO/pAHar7pRB38Ppcwhp2nJkzLn5Ugph70CFmcx
oAqZvRPNrCPbL3a98QZltH8dIYAE9hxD2WwtLqkMRSFiXGhyFr5IbiGBJaLhskF0
l/9xyO0I3wICZbfsFezpPvYccPRqlVmqPHkDBw9ixFF9jnIZnf6gkbe9irmeVlN6
4elF/i90wj4tEW5pzHZkYwaw+md+SmeJaB/87pyTXRkI+GeBgfdu+NbmaMG4iV1+
SL6/NCl6hIcAqZXYdP0eNCbV4vJ0neI6moiV/ANb9ThGyJJmsD2tOw0YxT8McfXF
+xaXKIE0w6wp3nKTg16ywkhUvQhaCHDbmkpYEpKKIKngd1gdv7BFyCV3gYMMlcOg
aVWQaFcjzRimGH+E2x3FTu4uURU/kqbsVYbfV0Mj/8yPQXvdYfKEH41lpUWCfw3E
7zHL3N7rKPiYTjQaTINitc92R7bwcShmd0vlBVBH+UQlbmWA219l9rz4sEXSdH6o
/XRI4v9f7g+N9WLpoO1+mjmgpsUvPSE/A8CV9D9kHca5zdzUaDnRLF4rQmK3ECXu
Ds0vryww+lVZN29dM9alTe/WuMTFDu/k1TxiVjoKFwfIYN+ykEDhyiiHVJfEi46Y
Lm2j/WsF0gkXpxWEFiqfBCvZ/l6fI/3BXWQ9BvHnLICyIUiD6l/6GIxRQKDQMJpn
MM6bTFhhj39/9CcPx8ZvUoEeRJoStEM5A1fJqGfh+Pe/ET8e/cl8UeQjMz48hBmV
CBdpF72y65HZEevayY0EM/eYLvfrjPuSkPaJyB61DZozBDi1tUfLnFD3Pytk0ZWV
V2zOnxHfl09OcXnz1pQd+YQTOJIkg4spaKRTEhTSiWuzuWAyyWqBFi+1ae0bi8/u
YB6rPqqOoNlTOibi9me6FEzeZLvB2/l/heZ5wswE8z8ek1dNGx9dPNHMWfvKg8ws
x+efNn+QpF+1ceY06aZmDky7E277t4cSU30U6mvDTPzV+GzCFyHPZ6SRXydjo6/I
g9xevCMt4EqFo1i8er9ZfVP3vd3rz7RNf0bHdoxzC0qd9Ke/vyo9nj/EzDmfvXgR
A66XdBfyY5y3ZYeyWtCEBx52SZMpOw4yw8JetbThm1OjU/5HSeU17G5MlGvHqOu1
fCNvcNFb49xsBJg84vaFnyYXBhwlko+NLp0kOKtZY7LUIQTRDUQQKM3INo6W2Gj+
2rqDFlzJrIY1Eq/b7+Tf7eF6cBawwc27QOxF/ftnlSz0nZmGHn0TG7Nehr3eUxgW
IWw+E73kaqLm/Me7BTHmCwwskQaKQARNDnsNOjAZsCLeylCM8DYu2DmOYG9pJT5H
J01ApOA4MhinUMf4kFkgtDWH5IfmSBOxJ5Bf8D+TqrggJ+AEZUPhQWG5oOlqxg2x
0vDXhH5hE+/5l2GhfpYaESnR95qCBikGW8k3ogUcp4++tEuzNjEHq0NLUNKYdyZt
LCCgzfOhYdPwQZvBeL+LvIFIqMhOBKdefnKZS+MLTzQU6sWEP66Kg3+crwIMenPk
O9EpIIkiqSlbMQSzfODDzzQCXkt2679Yyqr1ArazNdFZNJhNZkaSjhQs/sKZ+64f
25Q1XtvoqMSI840yitjauIyaaUvQhBPXwJF5QBp38SuSESEKN6dKy1ucigHa/1yJ
CYyeM9YHmBfuzxoiPFOu+V6+Soankc5PLoma/Wegu6/hSLQ9saB5A4NgujDirsFV
lM3uvo9V3y3H8zr9vmO87Xv5SFQkHScOXdh9itzRwyqZUEO5PRU+4ngXzOpBb/iv
kO6HyuiQj3bcw16XhGZA8XPPJ6GRlJaXp/ohK6jpYQOrrcimYWWDZyfPrcqaidaz
JXOfFGv7Nxu4GIyinwcAitu6lILATCVb0B16Q+l9HC9NbNXFFV2j+8NOgJm+WYHX
yARdRalxG/otx15jowN2MAtxrBSl2tOp/Awrbfq1cn/AFVkaUaU2GbpIIFV/4+0C
Gm6/wAtTBFXoIZ2q3D8UXcbPpgossXqOp5FLPLDcocRjYcnWWrYEmdcMtJkfeHEk
TaCtPcEkjpqbesMK59FyamkYi6xQWutL0ix87yxtrzP9KJSX4aqGv0Ub34ZZo4G+
q4lez9/uA7KPKkdBu3FV9c8QPMIfiI9CJln4UBjlHs1Wd/K1G6lbQblrSqZlZhCU
X2+0NQt60JQLFi8HtvWw1vq63b8sPrQSvxLMqSACCX1R7vJp9BLMhODnFtrmCOLe
oayhAuymfeEdC3Bh0ydNK0heTPU9VaJR34mjU/xfOmcERd4HASc66TOl5CU76vbM
mGkmN6Or76Ju7v4gYyBV8sYbDhUtVKtduD55ymeR4gZRvW3o6yKitbhVHy678cbE
CrfgOcbiB0fBkA6+m1nmpWcL1S4o02+jrBdF9Wx3lNxvhJQM/4xy1zJ8gQhIn14K
jZI64TzoQi3LETpRrty/Ea+Ma0KMFEYmg9YPZqrYx8DIYWB+quKMspm+rBv1Mt6W
wxqFXUSq32tc7rREetPFnzYZICUg2dtIUiG+IwxMhiks4wgPFLvqRN5/hyP71M4+
yYB+oXBNQ7bQ5vaUdVMJ97eF2/BC+SpnvHULmZwlSX6qxKmZJjfohbUGyKD4IsNF
yxRI5ALoF3uPcWLa6uewuKoI5poe6BIrHwBZG+NPx4duQw/lAaaAvOT+WlBbS1Bu
E3V4UX4H2f58QwBUL+dtJCFEwPwduOiIMZbIqSpHFisXtp1vETvnr12hOr5hug4X
7H+j7Qyq2B9yL+ylqUz0M3e/AyLGjeZBOySkM4Rlq59mvHAn7qlGIvF6cNcdvGXQ
l6U5i+g842xf2XGOhzxbEha1P3PXk9LP0KI5kCxYZgbqpjH+gOul1bgeU3F872nB
H/nIsw0s2GyoKypuQpy+5coIP1AiwTbiQLec08JEqkF4TrZWCX2oasyyY6/MwlHH
eae0A2wwJaoJTiRoLht2nS3KHbkStkWQHbsEUutgIxF1r8JO7JAKKWOKlHNlfZWu
YxUpDWYbCkJ1yh0dte59ZjhqidLSAd1dffuFFvnNH2L+vL4pGuG0WBb5ZAvlesbp
64tTm+GYuudhwmrr3wT3IfIRYTKjwAFSbB9vBnD5+V5VDZt8MwBVJ2EqY5b2B0lv
4n88oXpuLsgETy1btGONHwLL8Sx+EgTfhImPgg6R+zKaeitUAX3e4ik7PW0pj3Bo
n+DCbkhOBO4tnRTvaWXvACOgYz/W8cx46iR5FNzfurw1QqgVgmXEH+e9siNEUgWb
Caih/Cro4K/pSXlGd7DMCHWQgvi4URxg1DZuC1W4fjDlo9An+6x16L+cHhvtwIka
5CJPrCLG1vXF78aaQd1jfWzpLkXLlSJZARZu3wEuiAFPz1oLs1WymA1PNmNOjxyg
v2cGPCbV9vCbGTQrGxX7/pGxvIlUJCWoiEvqduCJsdaHS/WCRnhEyekNQ7UGy5Za
nj110nNaKpj6aUD0pdBKyPQ0O7HoQINPQ7r/hLkmQ0FuROXZaXgU32qtTpjlztUe
CGnYnmsBD2CC3RBPPewTF/TuDYxujFXi7UVI27XmjrcKCjltbRWGMuJjxqyhBSra
dO6FfbeIMjSJwTnwjd27k+6oP9itPXfu/J6WUe6K9bahp6Ye8/EzmUpQScFbDIYs
GksDhG8hFlitxT5oWl8ZYswinNxVWXPJvKn7Ir9RQ63B07q/IIN5ieN3y039DJOm
qPFm9wv9l7dUYp1qzllFh0gWaKkaoFsR+JD0OaDsb4xWPq+Gw5eN4DAYp49BhlKC
uJxPlU+qgScVi40lhn0l9SlVDVyouV2HNvqYwocgelgUYjGUyplJpbpIKjRN+lL0
6G4L7pH8IHuB3gC/t1L8nF+IvQmrY2XvHkRlVyZveib/PicN29h8OA9eDyMncrov
UGhw5HONDCJeqVH2/LXnOhLMvKkecjGiDhwnMEhEBirs3iy1Ogr2JqeL5mnzIlJO
dX7o/sPUGGyzelV+dYtdLgX3rpjzU8ztoPizYrPvOkS9Z584EGKkREyuYDZ9812Q
Z18or53JFUBqrwODOqHsucYFHzbjhB2v0NohQp32vf5ISdcAQWnfvkhBpCjZNrNh
sFFxnwpyDzIZoFBThrOWwaCIefmcIb4MfKbGIn3S4sTl2tNlaTUAt3l622lgz+6b
k8V+PRzZJDfr/rMnqvOjN1BSUHDev9OkvDaxUtpVz6jQTNoj1okRIZnj7bBbsS49
PUUKmEgs7JnMH7D5ZyykR2tkk5T2rX8yTUcq1nKk/ZQB7ISGByf5nyhG3TNNcPod
LKO3C7/6FKAUhKgAPIJ15WYt0s/QXWlGd4//ppRo9smylNa5iXaEw/iYQ7ecziwK
mR3BFnAQR5tNJWGU3f9kcVoeNnCaACt7G2Hw3a9tgptMWZZljytOo1bz8UP86w/k
bQ2HzW3TA2AHkqPyK/ED0/Mr4LXkBaXCtuJSNVEvPALJX2og+QgO9bAZy9oMQo2n
PVlo5Z28CArPxkXmv1mMeXcIvW40u+5D7toFuCV/qxrGKL4Q53vjA6XUnJL+p+wD
AzdgOfuun/3bNO/0fTORAK5jU71rSJy78lxZNpXhZOyzC8KkfE8A9FJcBjYNfmTz
hh+QCqb0s/VahlSwPgp8xGVHn+REewqnsG4UcckiYdOjL1xaD6L8hAoYebL/yCHY
kBnSjuw/ymxIZHgnWwuRCBUh6LCVU/02JDntSppfg7dYKHlCh1QaDVR37SZWXjuN
i8pv2Q2RbYFkwu+c2ZlA7vvcKW96gSEeGPaSBWfoI5gu63keWW5mZMQ558zRf2jO
GxWG3jB7i0+xPw4k3nn97asg4lxm1ByQs4I6S38BUWZ/C0dbYWpCUqoyCqLVnJ/e
f5V1DDWkXE2+kgrB7u73Ib+AmahE1jKvNpk7JBMy/hoX3ia7UGLEE1pUFaDZHhQv
Z94FRVr+aemyqREi1R7cDnYMUg6C0RK860omKepUzIbBnXc6m7BPoy2QWWecj0Aa
d5AeVe4oBufVb8sSh/j4u46FWm1iEcjqqwdqZuvaQH2aaZRiRBMyRoUZSvcsbhHf
ZQ1sT5Pi8QcDgslV1HKBKB20LM20oVuv34ZdlF/t+w0zMfhXEoQccB8UlikW4ZqR
kr7QYjQB5m/5x0Kz/i8+HL/cv6Xlxw4eNjsDUqvXgYTdtPZd4rMRrGBm4XIUMqVZ
fTp85NA0SmD4aRN5gjUh4rdJrnjYHU1X3IRAKKPONb5kXe58z5HG+Z6P8KLvysAz
ddxdOfSdcb3xDz0dWhqvkhvyPsVrg0deHOS9wpi3oS0BO/7Lex8z4oCKMPldILEO
q8UPUoDO5aCOLegZ92MNuKCh1gQErFZ7dZ47hJDRZatkOta/gJnO7bP6LzV+jmoD
dFWVi/gfZfWeKe5QwCy5WMvvtn2jusivwRz4Mzi24BfcsBZbZ04WasY2XC26nB3Y
NVZdFqjwlP44/KZZSkml0/ofT4CgQ4LgSmLadwMo5sWg2HiepY3o0m7GwhKd7ono
dLyVOPWS7Z8CJwnu06wNwS1PtDUlVlirBjoB6vvazU4O2SNqeSZ2ju7wMri6H/fO
KP3CRqQ6tC4h+ZrTa0qSH84Y35+NdPk9flbIJbAoiUuwE/JDdMLK73dUhA4n8/3C
xlCUajAGTmlGxpvc7zsMhDUg6+xj3YCX+dE/kswvDvioIkPyHgnmCc8ScKNgh698
+KJsMqsNNQGAvJwpriHog1ycTY+6bj+jfuc3fVyPH2oE3zFbiv6XwBRbcyx44uEw
+sTYKzRxCo2NeBr2ZSlnxHTfmEnsO5MFrYAW8osV9hLfqfu9IOlPqh2UkcgHsda5
uxXkS9zb8x3FXuq1ggb+NjjersQwRVcN0nt5L2NDs761MAJxjiNEtnGHEJIVt5ZF
3a7HruYU9uIQIlJedZhEy+s1YQWzjqjlqwILg4iYXN8v4u3SwT2U1riVowRcjb/t
PWVOTV8aXJAQbqVAxwSqp1AkFr0ITCvRXhM4kxG6Ngjj8v2vOcn6duMGkPL9B8wa
daQXSruCoBeea+MG8lnf4zyUHXp14oRdJifCvluc81Hj3tpWww2K7vHFqtCf2Hpr
93syPbCtkFti+AOONadum8qMLpwJs5Nif6tKOF22X2K/+TICdw3RYSlyafqfgCAa
9pgKFWB6Qj6mqjyXGAEo2QvUGA3yGelOYkoJSzWFmL1EUIC5fLSflBv1GrATgEPi
COeG3/XLsJCM5Hca5ftDT/YaGYME8Yig7Fk/+vhSAxKstiOAXIIOSD7jBwTBqurc
f9i2yCaBmpNvvAl5Rr78YvmxjNcC16+sLPyQ2jHLZyglg4x4qiL/jlcydJYyHN0r
T3IAdOXpeRH+3O3z8IcQcyeb08jmGacs0iXwv8BLC9hapqOEw5J9PXdFCM2Wbk1C
YiYe5IOurUs89GOtoVVEdOL2SagFQOygxsVKjUjT6lZzuzDIpBvmNss9Bx48hBVc
rMjAvxkacnN81L7VxdP9ekjinHApiZmAYn7UoCdpylJswVlhwBt20kDi5b4DhL6i
vr3PUAmlHrB5UIQ6Xk9EdLfdVaZBZF6dUusVIhNq+Pua0kT/GFkCkY/7K+GMGIMy
wKe7MG6zGYllhMNukFmaK5mL/tbkrpzXZXELYH/kWijOzJwthSvNHgGycupAt0tG
gmX3RaWR91/qudyrsC8sol7F+0AABQ3cHJZmuE0yrZXj7iJ+VzM2KrjOErHNpLlC
GgE8B0/U3kcJkPAwdjzq8Uqbvl5jr/79MUmkO59vSVTn5bXSnRsbI5qC2EAQmk2B
9s7trMAIdVFlJ1HH54tjxPg7aYoerWL4E1QDxnj/pOoafqm4Q14jM14KciabFLx0
9R+uKWtQ6YFfjryrzVyrVYUvk83bT/jZVZ6VyMcHiEw7QbvBKeYRjICrBKXqagv0
tkQ1QvYGLhZxEQ9tfQSR7TDRTBRPtHLx4Wbw26EZZ1WAGcPcXK0Qhs/6USTa6sCs
SuavlxvtUD+snPJIdN6XPkTNBMMAQWbAJxpeKbIfJfiGR6NfsjJaZJGPgqJ6lIuM
cYIxFNYGv0ApIxmw2S5a0o4vDQJxI0riTQ1Rbjx3jicJaALjWL8vW3qonxyfQWWY
jC7ve1mvGsE9+HQRy26Ycewwj5Oy/LI4jTs/XY9yLt2sewOlVhqPH/2pwYYyexbB
puNTws5Cx9x9k3IALVUD1udRMe0+gId4YbEoJOC3yxqNEXppZAjcdgzGyow517F2
zEE3A4oBewLeRz7P5e+4xovMqks8R/WCIhZ70dO7MjGydsnoWBiUxgLsS6Lob0sg
sVMgDpO5wiQ27S4C7jqi2DeQoOhDHJUSOdgkFVlgNOZbaNbf8g3bw1HZaVp2LHDZ
rVSlwiLIddPlSWUVv/L5XVu5tdfLYct6oE3fu3O0ad5K3RO2t3aWhTLwOcsDe71j
hENrT3oJTw8J2hHIxdO+yofcdJ+EgZFti5880/XqwGFRZtHzW3u2CwFWsClC3otj
trEQTeckeQWHQE/k1jkF9Gj+Q0r6HWpFnywSv9vAxygHnYvnqa8gnGHB10HHwlDN
6WAIlEArX7BR+/k36ADMYbbl+dTX9fiICiSd5Lqb/2bXYQ4DHPzpVCAYgLB9ITrY
gMIGVOEsuGwHTel0ZP8PmYBlxgNyforgcguD3QJ7i+uZId3OccLeDat2PJlwf9PL
QzFIDXVVCSpb0D/79dlOaZyEATE4CRQW7XX607pqRMVUJB0Cysk+R/qkbmyZAe3b
JDHDjMEgrxwSfiaEli/uOyplAPjfsTQDeobQGh8ENOKD18VWPWn26X8omF8ssTi9
1aBuSmpRqs/mq34BljgsHnWDtR0QvZDRwLdrTorpfnnGBd9OK8RwCHrquh4Y+YKw
1bp2fqCsMD7j5ojngWsLBW763L1SfnCZz5i5DRe987HPpl8SDLHNed0UjCaPDEfj
JcS6yaSBqeyVmfY1gckdQE80suUm+yUe296hIzDHUJmkfqGQ9fywhiVlE5S1n611
GufEtt//IVqWzFdpd6HWTxai5ca4ij2giCRGwjyrXuMaHGIfvURVUHzZc2ZQmhul
BoUqrhTMdX5HNku5T7Xg8e+yGdU8DKzGeqDrf+fa4KkA3TPwYaU9hxBcOwnLjbhe
2DsRAzdWZPEJBwFhe3ApJGzFs/H3MaVH+iin+tVQ8KZyPF7nCJZI3+uUvQ+jyVgG
hnbOWrKITgSyW36bU8RuQKrGL5F92uIarZRowcz3DnhW7G+KtVTe6hgdUZVlIg5n
Y5UkjEdZRBZOBwqOHTlgy6KfWkSg1258VpX58zhf1b/0n4qhvamJEz9r7WuxMBlw
Y+QEIuT0Jip39CfLsI1COD2yf4RBFWjf917QfZyiyzimd0M+LgoP0UupyHvW1jvP
V9FVDW2sKTsPULZR9zyRNL0NozWoFDaihrs+p/UWKcEFl5tLrZ6HZOfsDX5cmvPS
kvnHHBlu2ok/90/p4cUUD68RoJIhtPjU8bUhRUySZnasvygbOB7B1WDfiPzjonJq
h22ksMyq/c5LaZGkILWEdWZ/1RAbkCSFhR4Ep/Lv+9ORpWmrqb6iRlnePouvlXnK
fl2M5nS6/hvYMUkBUFz9kQIcbAHiaLhe1fij22B6Mw780nVfB/eIxnAHzJHNir2b
nRFe61sZhdZguaUWUx5Nqw+UPUNa4rz9BBiMhjj8XfEERD81UEgxnXeeONpiCLlJ
Pc5YUg7jdCTz7io5mb30iC81yIzVwo3kfTFnngR6HlutX37RWn9KS9Zk+iZ6XK8W
jKTsXcFQDMeqHZkEb59W5D5P5XYPua2CGm3+m9j46KmQ0YNrAe+rKVz0LCf67gwL
ZCcwamp5NTC7yBdWBW5ZffPVYisyo1RKhXf/ciNx4hLeQUf1o/HQ3dP9pbD4yt3M
0ynBZ7BXAv9JTOt6JswR5vt9pMSbLj+2LPIgTRv8KgenAtrpZ5xl8yfyDWD+AZ3O
yu0WDIGTJb+sU+zZLNi6OZPI921huzCzfImStWtm+HY3VDbxTJMwGu3VshkWOm7W
7nk+sWI4HHv4lRV+n8HoNFu4MZB6TjTU8rdLwVT0wkTthmy/NJSW6XfBbvQAIT9e
EPTaHBucudonpXQGcBwY/tBdKWIAs2+xX7qG7w9SqncVZTKZqObarnPdiKS/Q/kQ
kQqR1Rpw8POthQPSdw3wSfQoIVDIIYPpf4oxw0wdBu0qfzncjY0aN78bA7IfqioJ
Y8KbSnCojG5oENs14lQqQT//ndN/I0LjHL3qo/TlSnnOTd+rIgKBXW1P2iHCy7Xw
FCvPkpLbsmpb3wGf4P4QcevMvzQqkOpJGxSUMMRlUwAGO+w5Q8vovETk2NMhxl2/
hAC6E4N61smkB2vk+10j0KSbzn1R7bZ43Qt6HI8eKy3KWTR75IzdrFJ+78UumjpF
ZLaWZZOObflQa4OIqIJ0jCkR+5Z+vfGCu1QKu0z07wXAXa8v9v7kmbRm2Kmt72Hy
Sce1S+R3UW5z8wRKZNxiyhhJvPb/wKC+4qDBom9tSTjY62eId3Vx8ahA1W19sx92
lENXlmDmX6E/Hh2gKE+1Kse+ln+nE7EjvIKNEO5rYc6RNoIJrYiKjMqD/9MCup/e
YYcoNW+xiy3oT0oFH2gJ2uDWgPUUd6i3ArOUOgqicxLJ2rrG6Y89pH28pb86VyOG
bUJwkmNbjTb2vw5QJ0qRWrZrYFp3lIQpbsMX+eYc7nrB95mZhF3TkAAk9ki8qIHk
FlqcY1Y+kFVbOCsUghTWVGqoz7abgt4bBYEn2bo5QYesFOkLLTZ/CqPSENOraTkd
4af6A/VFpAHgKuPUhfUT5/kG2bbVj02G8tkFTXXRSZDIUMYW4E1ZUDYsxVODxx3H
q+WXXsLaNWoO/jzKTuKnlqURA6yaeHbIBQfsc/1EUVIYg/G14WQigLjclLOTXBTP
V5tnT5XVa2gh8kRMCfcbowoaTOm0yajDXLlZEc4LyajvbytY72ryrx0vhPFTF+kO
XuiTmxdU5MPu6ffVPx0HRTQfH2cr1Z5vsSGc7+ZMjswK87SRzMzOthgEAdMd+ye/
Yn/fu5ntuFp3kDW6b1Au5NwTBVfbpqSr3FL20LY4JwTER5XTkR4Ec6hCaXPdw46q
Xm7x5Vd0dCFPkQb5J9/Uv8MhFhQFSjc6qxvJ5Lu+LV793lCgJGqWu8JuIJ04wCRv
LJPq0BdBv+GLX9EDrYVLjOHep6sqhAeq9dJ3BPwqrV+QxPRWU7+t9XR1JyzSeTss
xDr9pxi5mu3BUg+KF7oaNtwiAkB4Ze+IBcfZLeEERpOG+cUHXfMvphgB8Acdx5Bl
V40tHK/pNP6RiuLj75rph97lNM6wzZD13jhwQmUddnGfiv9ybCQjdU4mM32aDTPM
QETm3vSehHVRwun8lBaUDpQ4iK8P+tlItaE5p49oC9YEviGcdm+XxP1OGJiQw/K2
cjm8E1EShZ4OpXu8qcq3ladOH05jtMDr9mBiYnPz/9alTNL/sPhTsmtTRgoHVo3f
XvBDqz9RwyiNfn3S6xVygYqxsr8nQszIan0eZT1dYj3D3owWKicGyLpXSLUuny+P
6n7Y/YwPuCyMMqd7A8CePGTRxFgSUFEL+6lPfFIbBsIl2P5U6Ub/Jxb2HG0NKsvH
QF7fVJjwO8GTpKO7JyISgxfHqnzobtASN8ZJaAijrGc3JeFoUaCmISm2qijYPyIl
YGsxOBsi14+IJ/jaNQ///fcJySskU1MbgR/9Tj220Xla0vxuOrauo369jcIuoNtG
bGo4rnEi6F1sLdQKdYgLutbGOPeNATi0pEsISOsRQCpA5N3+xuXMtDsknX1le+U2
H2sVELYOUmoX1xu6TSHoOa1VBcg46fLmcpYZduGXlzum+c7/aQFyrLukai0jsmCI
nAgPHOgxvKz3GdXjZGARl7pNp7kOLWcFBQ0mx2DeZXtiFaZmImmJArIMhl9KTKbY
vK48oOIsAQpJztzyvId+Sky8x5dDwLBlEzmmVxGk33iE/PdxaUck7I5LDSvwUDkX
k9be1fIjQEpL/lCunC5+CFbdUHqh9K5Gy9xMjRwO4VZ8Ow2jyFBrdOe+yB+yNBVU
splSxJs+C0WjIgPcmqT4HBNvy+qZvAlFJzBML53B3zzHjOMPAvuteIpqvfnJopjp
+k2U+WdL3Fzn5JjkE3DBZfef0wknwsGTRE4i1WYyv0WVLb34OzSKNaOa0mCujdaJ
IWtbLtYsrIDRITxOPO0c9A1n2jnMEIxqs9xlut41p5j5jctCEPIzDheuvSBcpZQ3
82Bo1PIYxY5ZayiisFmrD++vY4IjWrzJ66hWcLQjG4WhXRt9kKdkg3WiEJZP7mnh
/omhGe5kR3W/FMB3ubbSHuqgxglgWfzpFBsJiWjdjFPA9wPQqBJC7FRyRe1VpN8d
JxrAPSh77LQozoqtz55u+cj1V2GfJ98lZ2kfv0VIPhQtrWZRNQQmVGvPN5i6gjBC
XUHS5TPcebyj9RLSQXcAFevtJv64xe3RmVacXE9lpXO2QZPs+em3tmNIhBbr6NWn
N+ndD1BOzKLIbOdeNq6HQe9Zxl3n8GklyzDzBFsnOllnfwsJiWBCEYR2lCnbM+6a
DsjL7tCJ5sMa8s7rg0ryU3UsfZe2BHqlatTQEesvVDst94/aHkwS1qhlpAqRgyyI
6awbMPitQ6XEwrwi9eCd1cub6qoYfWONB5o/poAbXK3hBz+D2tQ5NY0ufWuMO4Hx
C2iOitU8ECteIwyLnax3g8ub6ZdOEdR6sfEAIEfFbYCZ63/e8m49YvvSbBOB4hBt
sf3cHbF/KRt+fWZ/07ygaFFJ9zFGgZcnYmk21GKWS7x9YTnUG9zJVN7tO7PkdD5A
`protect end_protected