`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3824 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
Z6yALt3nnSw9nTnZfQBUNY1muufZvtlJ1uGMQLE3CKiUIFxGroeb08GWGgTRzUXh
CWuKjL3G5zs4vB2c6/yXafEhkEuWsoK/9JL1wAM01v7PNvj+BFubUmUGIt0cBsj8
cugLuo3HHiM6Hc8hEjjMaIdx2Wjy4WR1Zkckvx/5BUk2TI/Nhp2q/sKvuyODXKO9
NBAZe28Zx8aBB0wyzsc6rEFP7wbL80ioUFLjJa9WGOcgsj0znV8Jyj/vL7F7fVJ3
G4Zhvsky5CbQ3YKoazX7alwQ0RprQe01aUB46NR20YAymUK/SnNMqaWodNQm8GfK
YlRZlKj8wiouIqwC9JEijTUHty/Wu9t7TgyBpFXbNgMP++HcEnqsgAtQtVAGF52p
V8x9YXTDf3a6kPCk42XttpuihAr5/YMZ/pko4XSB2WVJ4Pyhf1FYGaRdhLvbqiiP
Sfyua5SQrJ4WtgmQPw5k/xjhosiGVAI4cKdO2KdgC4iLnSn8j5e5/gNqu6AElFQM
wBjVkEJm6gWTkspcPT3qB5GKe8w1g0Qg+PJMmj0hfm6Ie0shhFAsWJZ5TnSO58sU
pS/c6Q47RYq2a0fYv5A0muuZvbGoVDGLGgap6jLtsgLwC+Ml5vP5/SlQPr6LoVZm
CMLjIVQV7DvyEReW3bRsFEVDuepSqFhMZW3FOU3HGp1PJQMR9B4rOl6L508CTlgH
vqCqoLUmra2bxYL75+QKFOw2bija1FsPeuGqXEv1JoA5KxAi40cNnXcUB32hYtTM
vJN+ptG6uHJ2cecrnGLlYSaKA7HnfcVTulhFO1lCN7ggUyi0Wc6ZtgdSFBdJ/f+k
F/rOF1DkTtZmMtoPtHJuuSiJYXpvR8fJt72ZanPrJixvquXX16DxMEo7krhcF3ab
P4nQVhiI2yDGM6DhUleWm+LibWsZXmIMnl5xv+moVpWFqaKJi9P/rPxa8TQQFU2z
SPD3pVzX/FzVaSccIikJF7zOIQnuMwWnIIEjCFDfFKmmSzMxNQ5xuWCusrfx3boT
6U4zSbwZimRb0vnoMC4jPAMy0R3DBSw39leWK1ptImjsgdTNTjuy1ZSe2jqWBPSn
J2TCDBd0C5V8aWjSOZwm5l6WCp/ng65DqDr6XYOBLps8WLcjwoU8uLiSBmxcEo+O
Labs/0im6hE9nAsTwM3IBd84KcljK7mN0YhluZKSmARkR8KE61sqOknjo8O626VU
mPkJkud2+gn+sEdKYVxTB7BaV1wk9Ooayz6w31LGM92eEUUIS3KY20lTU/wXTxeN
9OUkD1KsD5SRubtEjo96rw+O145jhFSiGLxRzRRcFrgnHA99vQoAK+DUK+hMv7u5
5ZviJSzUq1RUBm/YbJIe9JYQTFF3U0LSgS2MGg6lHWDCxrj60KvOofY0PPQorT6z
G+H2dbg2AE5qHFGolznAxiEKFvh/aGQYSEGadbo09VikbA6Qw8uO8O0Or9sgimhI
lCHuH0Uj7ZGV2jXwGP10o8A3iqSYClS0ybGxpl4ni0jmakUIgqwTpJSueNevb/ws
f7PEoL4cUVzst8OMaNshV5LQhn9V3PpqdHaKu4pca4QXtEESrLyOkGSjr+R/0dbq
WvkvOZ7MGXrTbq6G+duRXCNYbGCVLzcQ9NE64XYopFqKW91tGTohjNc4KF/UBxJk
CJoFxX5cyruyzlIYyTCazQds5xPpG6J25tTKddgYRmbYpDG8j/Og3YmIpou8iKhT
ll48azlCl+BObaqp5g50ZIcDD+X9glKPnGwkU3jby0eamwclW9NehA1dnID7R9E+
attIzN8iargKLIgNaMfvYR+w0Y12bbwNCpkeMXlMQvIiTIxXzlt5aeuUa787wrb5
wIWyNrrjGcE5KIK+I5JBi1HSeA7rtxMKOfWWJwpuLCMVfoVZAKUtX7c22d1D/rk+
yVsf4AtfcoeG1gv5OmiPkmk6oxkPze+IWxAORz4y9psb9Mp/iTx2uA0+NuBgB1K+
/p1hVJtnWOr1Z0IxnkwxTwRPlDBrLfB9ddxMriTUuN3Z9IOGfNaqMHxDpioNJLDw
VRnm2djtnfSiWpCfaCPU5r6KzFkEE0Y3lyqqxj9tKh0Umo6f80vpL/0u6XqHNPzh
suJKAoFeu+3nZxJ6UvhalNwLT3eg52bHn3YtkelqwwhefSDr3T3sIKa7NZHJ+Fbj
sUXFsiYELafqHIx0mjeNCmUcPUxUYlZoAZ16x1ICDDBBRuZdDDvp+Jhm3WoDbQRe
cqt/2n6njldUwSon+aiQ6m7Z5bAt28Hia+C3bHygQp49kc4uosyYn50v20d+di4l
s5PG3dPvZwXWF4FAq9ZN2zBsStJ1zK27IyfnlJ+sYd66S5qcSSBiElYzvGrqA+VL
g7qlQNo8HTni3taxiEDBCEtTu+i+CqAh+TX7V9ljuUQyHnTgFPHn0zA5wtw2UsT+
ddrdJcYuF11PJ8hd6ysIdEQ//EFGaUVE6icw6fss08lnKSQ36uCueioAnXTH+/t0
JamKQ6VgpErtV5lfPQjTtdxeyvQLaO2rJ6DY1eSArGzzGBBd9GWN3IGfOz2G5ynu
U7yh6NhyUAKThJo6zQ7nQQ31SD2FMERXcqPTGxgnHiL/+c76W7R9ccltCOOYuJOP
gy2zmtaTVcDc2P4SnrzNkEpLjHNXxKa7v6Bc3MKhb30lrFW8Zu99+Nd9ZdIjpkNx
8PCXtjLhMmzGsqbItQ/nDp68IVrnpjK/sIWjsKzUK/JJCQG6QVR0x91aqyvzh0No
7PWBljWj2ujTXbCIcCO0GxdP+WW62TqGbNXRWo1O41wnv62H+7xQQZDn5jm7HYZ3
RJw2xT6g0Whxsgn9XyAcjq9HHyvp02/72djDczYE84OL5xhlvYrrcZ5DeUEsU1l3
TyL29f9ihblKEjpIKp8koIvv1Ki6/2dim/1hjk8aVW+sHPbfrU/QN/B25St1R9eM
2vyFVc+AVbgX3JyK7mrlCnZgvUeXWq+7iVb4s7fE95z/NnPnY29yUusody17vivJ
ME4p4H3gu26XrV3yjbfbvpnOXQj41qRRqDQ5iMRwas26KhZ/5bnUpHclJqnThy7B
8HeTfc5ivvcEAMv3FOKN8npQhXbIu3BK7v11v3GIaB4WwZY4JAeiN9wF3I3ZjkN8
+4lV+LeP2/Rm2vvXvl1ItZ48E9PDRzuj738y7OHTDbcoY/Ci3TpZS4etodBXawHE
igKxlEFNn7vi75sQnVupawlmhnaGYO5P9rQ/Bcy77rSO6Qh5FT8FUxMcZXNll1tR
4zapsHg3iMf8MoPc4k1iTgK0wCpwPgK5pPQx+RXaJVvQ40iGyOOi0UGfSUxTbQEq
N3hwFM5o5bNWP6mhzmv1Amp+IMLuCGBsL5LOSLaFmvA/z7Wg0k3sqxQ0e0lVXkZt
QtdhvEejVTw2W+Cbc0x8C6vkjILGvTCFJ1DKcJEgXlgTGezxeBKdshS0Bjkqy/SA
leSmGHRJGsTYQkJHCV6LH1ktZ7j/hUY3p+6IG29x9yQeMJMJgk33QTFZJmABbgKj
SzPABgbCfowHIRUpsdBM0E4X5dp0n+4lT31TsKqv1KhYGgK8yyp7XY8soz7hOSPO
0TVZ9h+yyC/uN3EauHGatfiS3w/fi2Dj9rDsBy/7JXpk7hUxMlsQ4QZnsjmh5ax6
JGaJ7MPd9vvFWirKX5YhZXcAFhY87J8AipBHaEGhm/vFV8RlJdRh0I0xE9ViRLWN
SlretbBSjZLvDwm2cPGi5IKB6dWb+sMWMsFKetjE+a3DSETYwzjnWjpW4MB9OgYJ
CbTP61hQIQY7pvX37iTSrdsTHMzFh79PVCbcTegPW07H+p2kWGPooquiXa6ZIDE/
JGZxZd5bMhah+iAHs0pJP9R4FZXv2vpKAwMNN0TmkKV71dWsiBZtVhB6/C83QHbq
fTb/ioz2NZx9Hv3/DsODwdTEYsS+YMaPtyYEyOORdnHPpOf5eVW0jADRmqBgbKke
tZsVU9FAU2Wkx3/R2UHy5NE6mWCAndFJST9U56wZgau3W7iOuTvHemThkYB55LDm
qo8k54LpCFv7hmVP1IVTOs3y+Li8fYfUNx6ZjLYxK/u3+h/HMO3SMluL1wTi4hxu
kyc2HBh1ZnSH07/8dTTrQxaoBkuZznaYiG4olIbBmyBrhWhtkDSIkauKvbjE0RWE
I1iPlwz26ayozMtyDMFwgvmI4uHshaf+scSzmlNyAM+N+O6FougefxycPGoeTdtY
r1cmogSK6FRuqkA43DTUmfmMdD7DC7CEuRIjJIAAgPdNvYGxabudXjJ8n744fhdv
vY3NNxUrZYQFmb/EDHRVv7JYQg9MPmghxJWSoWhPFHfWqJdydQb5TBruMmEz7baF
sHhJJNksoYz82VVeJwOlPEbg4MWkpSYdgT7duDe1Rr2VVMoFkyJ3YGXOboMBOdPE
YHaEnqJFpBLYNTvCgWUYkbng5EbAKeYMCFuAB3xCybEY0Vmox6ddXQA0resXSk3Q
PAymkQ8SaKGyvO2TqWJY2pR/d5go2NZktGhKTNez+9hYnvoiR6QybB0yRf0e1gAL
BLruR92VdeEuzbOOcvZaZntkQ6QuwsLElICtj0myeIAJgBXuv+GjmuA+B7R+lakd
9pmi9qdid4JQOMeq8x+kDva195LT8twkZN91cimm+kwGftGZynyT7DygDjdxR1mK
Fyr+xpvcLtrRZvOP/JVzZBifyC/pxFsc6/z313yBwRZUQLi2SL19XKKEZztcRmlG
DYtOSXUoId/JZb5I1H2Xggdr+4zk+S+zsBpALeyIIZKDl4M0t7qbfwedtovi3Twu
lUWoaYpTX8761zw+Mp6yvYeCsIARqXPRoivQVcNV/c+bUkoQECxsWYoYdceOmd7T
ziRC/nV9FNEtIFQKnvrJwzzy8Ku/CyjF6zdjwZJsH/uOyx3X0Nuatr6hMnhwEo9G
fufpLIxrmaumFJT4EBwQx6uIp9+sj9TpSPPAjmRy9a4=
`protect end_protected