`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14608 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JXz1+zHgF4n2s6TEZD4KtuQ
ATkS0e5WlIVeyjNZ91Ns36sZQfrQ9R4SbnYvAtVIyXQby3GVeS9QeIx20R5SLlWy
Mx+H2tZLYu8alGncmTDpSdUU9JntDbm+hlUpHp3NlZmYXw39Ee5Ewx+VQHH6s9of
PRsMxUCDG8wjulCBSNdNiwHhSXbbA2+R2MqmrTtveNdKB/bAGvrxVPKQCaW63joM
hD6tknFIN/pGpKpSq6uPo5nfK7xxD54w9GNRxVMZMKTJ9rogh6hX8GWpE9GtUiJ3
yOTWHAw1GmtW/4lfoGArW8aznhhghwMzV3muzANOWy/XUljpzK8jWFq4mmgOW1uZ
se+cf/ryZwK4S7t55Wy2rMhAoDFq3Des64YL0c3/arw5X/LOgMrQUw7Is6jr+p6w
claEpqv1meXi9KlpUfHj5wHfZvBm/9m+RqR76iEBpnq2JGh7QLtoQuyLPZfSl9pl
/oBrPILdbVMEtGJcz0jkm/4ZRob1gFgcx2JbuxHBl8+4L8jDluUB3xY/P7IARs18
UxYI4A2cBRH5lsVjBMwQkuPldsXT+aP162NlpAQ3JOsjL/eZrWM6C1lTXr2lNded
OgVI1JNEngAu9cMDOWeNrfd4Y89PivIZXIY7qs3WQhRvm5SX9YtsOJjjv5Z9mSr0
Pb0QrMmi2ZPHNjCxxD/wWfYSZm0Xc2wR+tnH6ue7dk2f2roWwyeO8Dk/AyxHnNsg
boZTSOsgPOqDvdfw0qoTcdQD56VcpoUq9ZBCq1/ggXaCvDhygQH+GaAmXbwtUraa
SRcOS4HiJatYDkFeAcXbLOy8efJYauHOWFtsmxUu/cbOB5NjHxbwiCJ6QQqFbTVQ
kkk35Q5jo+5tL+/jAdg2OnonUs/qYLU9N/iKM1X8s1vPyAGEJbhK2OV39Guh7oRG
+0+sjLkHtEoJ/BEI72eM7+eh7rHQq8GQkRrrsKnfxisu1OxPdk7kcdgojwHqfxdd
iw2iLqfVgUxTZ4b2Gtl0Dvf1qTuv/FhgkUDlJFQd0nYJgnJC1BCSrA+2U7fJmPc2
HJFAlEY2os5H4WD58tgIlEUh8fi+L1MDZE0ZVH8x+VmHQUCuLnHdWrwHxqY9jBXV
ozVvWdlkKLb2U5x5ULVpX9VN3QY4Xd9tca4kuEFnfkAqLP4xqTY0AHSTGR/nc2+H
FX6xB3h0D4XiEAjuTXlLObS0uE0mfisVdPRG1FLwov5/i16rmn99IRx+AfZ9Pf86
Ogp+f1plhUyXqTewU4AnPsdz/uJeXq2kubFfSxAw6QbQlvBJ8iIhiYmfyelKx1zY
VjT/R7tYxyX0wDjxy9GSoBBrrU309Jd/X794BK8ue9CZAqLA/tlKsH3xVpgkBXjY
KUCjBGIWjrWOxRjPko6df24Z8zJz+sUD9HCsnzyOPkgHUkeBTo3BhioP6fIsSLyQ
kwD6z3EkUnBAb8fZal3yhs9Y6r5gSqp4oTLI6EiKEM0oUT0pudKQ8mKAXn4hPk9I
YgqlvBeNwUAhMC/3XC23tFLwWjF1urDxsWH7HSPXePco5EapSVAEt+Mrin4CaCLm
W1HEdZijyxs4yL+6AbGxtjOsZxKRxXhzZe86e21PqXwelVVow+fjzg5udKQi67AG
cEZBoo/4bBnLr/Hef8Sr45T2CZTB3EEjAvqY+gh4Bs6fn7rpAbOQvqhnNaEStaWO
Ka5E5bAkqeFQ+D4gNFuv5uKXPWuDiRkALdzantPmxSlNM7TlOmUebWJJZHkZ3vX4
JEdWz6aZmzPF7JQu8TlNDNpI5tndiFh6xN1L/h+BN16t/J/nCc0sdKptJtm9L6hB
WJvyt73u5G8zsaHKT3E44WJcngiiV+FfTEffUuT8Tiq86fsK7Ayxwcu9qnnXhTAf
L4nDNn/y4pGRu+jQsRQHYTBPsedExBbP2VZzmlz5ih4FKzdRYsvZUtv2JlmY7AX8
96Gx8Tuidbc6ilUVzl1+HO0HnEHwO7HxgjfyhXjNeXuxMzZH5GspsCq3gsISgYhw
ZsqN/uGg7EawltMlq6P9nSiPgB9T+v7zuhBCoWkLlxusSdNrldXealvYhbGol3S7
3jgaXUWfQn1cUah6uuoB0HwsqS8AlIQ7IZX2qyNlLrklpDLgcY1UTraQf2I+Egiw
JmG9DO88L4haPmtdQEiN7BiUbCSUn0QI9jG824t9wxPo0sPNS8D/KLiCcxPpuq5m
18iXYZAQaWeAT25WmNRQYxVVnTlbtS+9UZrh15pc0lJ7tD6w/nOiIjjplzCurLv2
KmqOAFUTkYabR+/zr0FGIEPcnKGi4Bcf52k2txikRnKCbYRlbwQxjq2kEAu/GF1q
aYdRGKkTDmVxmcPlGcqMMGoF15IYD7nEx0rU2KS5iQLvZM088OC/nsFx6itjlFDu
IOzR44jQCvNAH7QKGKQ6YKLqBFjcnier6zxCHEIgFES3eHKUAQzaKqg/U9at6OTO
1FLwi55lsOwdYHMris34FILbOpqAuQ/6sPNEG6ZeOUieN4BAjFnupWw+Jk5sfwXd
msehnMif4GXvxp9CdhI4NO6gqFZjjqXV2273QfA0aKZ6mAxqiAC0AZJajuIN+Fe9
Ql772FJyElcrI6PIewm36iA/OC0I7rtH1/IdraYHinmICbZ+DZ8a86WALLMBH5LQ
N9doIYLrV9RzvJmXGbnn1KJpceTXYKoeEunh79/pz/S8qPDDZdRdzQBJ+BvxEiI3
zyThsPxxobLS+3Oro30san2nZHfBXVFv7t2OfR+a/wgPb/rY99w8GWkhSJh8zyKr
DuxMLHy1bLKksN9/qY3hFPdepnhA1nu1a0O63+FCrD3xpMNj7RbtS7cRkDxayQnm
ODXgCUR831fJJ60KQr64zn3OxCni6zY40bpnq5RvaO6q9ktRYY2ecOCcrQy3u/j7
zsDD4xq/GhrTk8aHGBHk7B898+mr9d/JqKTTzCjxBaCwFKyaTZVwVj3T8HCGQ63v
FUf67LMiEnjY6JwJEA+kQPnU6D7Uolura5OXAwfFg0Qht+yop+QzwkYgUqT7yUbJ
ZyMJjQ1pEmh1MChbaDBIPRhpv54zET9uq9IPdZOwOpf/oL2YCL2Tdh5Dc+IxE4P4
lJMJd/TXG+7257huhrtRphX0if0mpy3gMkpA2HX5+mR+gbFt1l0828vPIMDIdriT
RzRAasxTygJdMMmXIRojpDUPApp0jp9ysBNce/8wYysxoBKU33J3BjiDIxEjLXfp
JVXoOFtRqmHUYvIMcrZmKjrjzwzO9jnKh02ThpLkydlk1ujyTRNr3s47iDrORkwN
Iei5W8poejdWj+oGbH4oBkSp7uCTjppabOKC/64jgrCQkdg44XIlYnpWZH4uW0ay
1AAswCMJsoWbta9s4e2mdNk6iILJOAtOQOMGFTVggxK1FjWycvbZKeSAQz8+WHfR
c7VQqR50RDIzo9ZRvKYgZgjkJFBl7J/qzrWOjq1EeaV1WHatag/Puvj2HGRUZ6Gq
HD56a1GnIH9X3rw9XJuevbIOwHfMpJUJW0s5hr18hOdjFXF6PT+RPF0fUUBmH+SC
fwiFTqaqUyT96iY+/niDsC8UOjpm1PmdqPpBFdGHxjYkgI78nhvMAHK2g/sEFlvZ
L2QUPP4MGP4wUo1gTgNKrCJEAQImtIjJnA0+ndDd+4hNvpRNupb2lSIy/k2fHwVw
Fa1iDcAiHctfQWo0IDX0WujknOxnDfUMAySBa9+cafIL1koVWkKLj0QFE4+iVcGa
eKWNNGoT45o0umR14Zha36i88n4R01FGqBIzWlIzYyMXhtOCUJLTfd4eNy2imDIz
qbDrb1QBhVmp8nah4hlPtw1GixP7oKrQN3TC5cNX9MYDj+nSwOZ66CHBnyVS+jgn
FD3N1JCxrM21Lmbdntaq0kndCFGtgiV575b9W5ytzZCahdvDQ2HtXqD3V9orgb95
rmlRHadNMwm3W/jz1S8ozOLGFMe9bu70xXQOmvRaaOz1o4oX/DWwzHAPCBogA1yx
IbDOYdryle6soj2HE9yrGNHSTXRdwh4mscVU31WqloCbnBQ7Sl3PrIQQz6MbYfWX
+fMEVe9kuhKvEM845R/beHpG+lrqBnigewLIcbkokPyJq8L1ndhZNuq8I65UmhQd
Iqp6an1KEMh8HosC/9GTOJya7Gh1MH+KT3xWnxiHgTo0W4+x4GXk0lc/r0pvfO+J
gN084gZrOsB7VWVc+aeN3t+hV66aeIhMJH0YuRRT3WoIGHsgRiBXecj4rfQbYsur
/gFHKpgExy4bAOcN5cePB8jZHky/omMPu3RWE3If/XN2yuywhIdCsTc9fZzpW0T0
BQ0emTfDUNawM7yKpDjf82vNTK6ln4wFea/vhVUEtW/Zvsr59J/rM482GMkFZz1F
Jv8lbr72XdoCYIx0JzebjXWWGK3rLyfV/+ApidUVbgPaq3o1amwjJWS7IVEy0L51
mVFwGEZPTSXD4AbqXiXY843ojpV6MGBAN5V9l5mDx1nX6r4B99urjMh6EpNvQUfa
mdvR21fXasuj/gKXtL7/YW5Zg7reaINwGv6F/FF3/rjEftp9O2R+xTGH/u9DqVgY
irM5v+CoXrTNeKnNn/O1hoizQk0KXLvwJyi5W/JoU3OiWM/1OdAw+9/oDaFsNiNX
arBbmFwOsVYqFYgeiN+r0CkavgBFqaUz9vHQGFd59XR+8AH+dnjmQV5dLaEpEnTi
PZfPLSraSws7K/hHBq/v1WaCoelezQR2NQBvmbhDtHCTPXOk5WoIZN55XS/IpNnF
a87G02hF+tznKqf/57Ti31nKjLxV8O4Zdq3bpK1daUb9WXml8CTRdDR5fEby2zcG
Pow8K42uhGrQ9gQS6DpbYEOfd2sr7czqxlYPslCsWfL8NKduuNuEjahLhGeygfqD
KFQTy5CEE1CgPl2VJ1hd7C1h2aONpxNmkQpYlPyhPuAUbBwliYA4L4cY2IwY7imt
a+uFKlAqbcg2bKVaqVHZdjkY20elRSp5gP8CyZVw19/n/por+cyI0+Q0MwK9B04/
IKT0BJBtBk9p7UdewG/JqLOZGjX747Xxu56rEBwp11snZtpqxEn+prukSVxZAszT
Rfz7NBWLoPE2ov9YEBbg+b7DrFOuWjVV70BSNaQubtlNVN+D/h2xFRjISgTI/owJ
nYQT72DNHt4ZTRVuMTVKl9m5MUourdeqyNmuJ7EEhQGU0g1zt97LbJ3HlTXzfxQf
PJ9Ot41xX74e8rniZSS9iJE+4dOoin9wT6te+GBDU/wOHS0pP2vnyoz7uCUmjQ2P
9w70TQW9TxHLYzhE7byP7rC0A0EXRalYavVae+Ga9hZhtowt58om/Gj5wCW19YNm
4N9RbGYuSFX+R+Yxoe/pB67z+cMd3nrkE8HAWtrmYMv1AuxET8PuNZIjxHyJo4WZ
HQdT/7WK2eW+qr6fMZOAHXNUc1o5nQQZFZuwmy/+nPo0YN6pse3gr6WSL8pNhBl5
KBDywSXB6MAbRoaCu1l5LfiwrosotEji4bwoSoW4+Tn31lox4oH9uMYTcilMJ24x
1l81MwAkIwd/aLJbTz8tmrbZ2SlBs6Q8V1mJBY9sy9wUj5nB91nTcUH9lQJJ7Bvz
+SJSxCdk/t5HaNMkCTLJ9pWDio+5HX0/TAYb7cMLVDm2tj7JTbginpPdlnE2ODOl
aZOZH0+iFONrVa30hW7QKExUVlwZMfdSElGsMu2aRkiL9qlHMLBVwW6OXsH17MRc
rtVOsRgq81lCLNPm9h/DdBXPIXo8lpLf7kZfqXqc8FGl9C/KJRQ74xoUgcXA5jcW
IOHci1Iri2lLNuAkJTbCMR9PQbzqpx5Be71LF3Kbk2y+wPQ2oNMLBwh+BuG5Tnlr
HcjQ/MbJEddrwbgkV+kgM6tQiPp99bbrdh5b7biJQvuHgphUTQ5312H0KexNaoAM
ACC1iwQFDEVBwsKpSew8NE2y0OTM5ee/F2JnjUpAFkX97F9/N1QlHiXGyslnMRQq
F9Vq1KmjC8L1LvKT8kTAzRPGNITx1mN4iuHJdBCVZfM9IY1UJ+8aQN8OIuQsMr81
wHIxCCJ7PG8a6XcbKF+M9tGB5BDktGtQClruj2/GFOcqzvczTIB9wCsUyceKIb8p
DNPSC6yK0pD9iistZFFAvPELNQaMCJxlqebl3svLJ1+Gbw+hbnbQcScPNyI0Fm7T
erm2EW3cMgKOS5B5214cA2IoZNdCypWQ9cZ3GgJoMvB2c/sQ/1g4/AiNHPXSrNYS
GVYcqJND5RIR2piKr95qF3Myzw/DetFiFB1c6/DPn6lhpr8Wnqo0nTrO2ECXx5BE
LEo5u3+2v9/mlxO3Qakm7qHOfPDVgsqdjmiEBSsds+PTEeMYgJ1JgDrMjl24V2yP
9gMt7vbERJYCgqzxr53iXVspsRN2fqzknnINB+CE/Msg3g1euINc01kAgPmenOJ2
x1w0hni1Qcu4sIkczprJ+vK9srY1V93Fwd1iJibSsm3yJjwVKZJcu1TwUItjOFje
riY70sB9rfHZtrR7X2YuD/oG1G36QnUOWCxOjO1xvhONBWEVQnYnb/J+kzLWVMsK
pHWSs3wZzZgchmMCaWpDFqE09i48gnQVuV0Bm6q+dxbCWKdvl6wY9NKRJlpexLop
4t0ORTo3wgQU82V8KHRkpH91B8B0DKSCl4JaFJFdmTpLccktwwDGKU6Om08ODLI1
S+BlYgLb3c6whO5Mtl7dx0Gk/ZH9vMt6MdaLdf6hCKWlSHIG7PZtvjACavXteTTk
vLkFi6ZZuDraznt+ygwQ3UXuN4Mnqzts4k9VGqqGtmxi/P7+lySWGkB8qbwiAAU/
WUiDDq7aRIfyGAoTA6NsQolNazJYED449w/ocy2J6Q2epNGvhMjoQMjZ4NTbJWVw
OuIbM6+QsqL3EQLrra64xeMKw/XjVTYmaJxm1anF6PeUpMJd9uDNqbsOYznHP+u/
ju3OtQHoXOy6I+fbd/5mY50DUqKB/7IEKqw9mT0ey6NSxPYtDjk4EC30y/ElgD4V
SQqz4MQCc+XvU1PHpbtagP1YUWu7EHB8fWL70pceD6h6/Zu9uIuWxALnsg0Ne/Ys
vQo9gjfTDU9Ew92/OmPDj6BLxBTL7BMioKpEvkdrvHL39lC6h21ILLpD6iOddVip
LqeceYQ4xRuSWmxTwKMNVxNwowAgC3jH88dO1zmrobvwU8l2oGW3iLF5RuXxYPYQ
8z5CXq0xsJrxvv5GEAW7ACEWEGW8yJCAS+h9DdDubrVXs0Kt0SRmw1iOALQhMKZi
T8YQPZpqxha4BMIkIOuiaTHzHMGS0lJqqaXjaCWNXg6rMnDiL3pzHKV3i6isdt3U
Xbt4SA5B5BnOKgBy5H78cvGbahnng8nYecR4mwgzwhoYJArQZikzy47ojUPMCfix
7fqoeFfdNklj9RD2TYiJnJEq0Ni8KmFvVgF62nDsCwSSg9phkih47+GBLqOcZ5b4
ik1Q/4fCHyzO12MujRbOW2siImpLOH7pBQHgyH8YbnUbXm1HMRd6SONWMTmkVY8N
L9zyTWnI7iUCCDMYcUrJKlG4UdlfFYDQZboPjwUEpQZOe0BgqeWjmHFIpAhlKtUR
aWHGuLUWAf4lbl0F/MHv29WJUk6XJsUFlmHD12Y3YsaqcQrrY1n7hNiSFgMiNqB7
8F51ZmSdZarxS4G5nLaKqij+g+gaFi4O3BY9bmhvQfMjcRNS/TrcYm74PIIFpqG2
olyColT0GC3vsmz1TadzN3HZXx96M9XbEy1ZFTx2KyOErduCoYAAjHbpjq9PO5ST
JsbldWCJg08Y/CgxN/OW+gSXsMoUWZElNBFD6CP+J/8tnPpceHuB+wz+n5IfCk7X
SyfbGeFh9gNVWAshncgIu73ljWz7wf7dQ16LjlG4WRuVaZk4ju5Nm11eq51vCA/A
rKXoomsP3mvNYzqp+wsSciaV9MHoD4JMcNrrCD2/kiuqJXlH7n8vmj2SUdE132pn
yqPOETy1jU/i5U72HslgMkogN2bMC+wAFga5vNsM2iJg8IkzMF/ANmAAEvnfSfan
bS8Zb/kvuigRTUTydvS4a9OTbpyigq0yiavBFg7bFMfevjEtqn+hO1PQMmsR6OBL
hbP6xORyPmaxYVOJ3Cz5bMTALh0NbihyttolcWI1eM14BtxtWVovzvyYVmSuO8vl
E3l+u6IJ2lv9VWjaAkEVCnaqo5Y9YShgK7tjDflBfmasd5p29ZCR+hYQY8QSz3q9
LMxVu2wKjiOFwaGSEjaD+w/XKlCi69cqL0zr1Iynu+BBwoLD3muNGX7ESSdOQLjU
XADBojkPyIdXMwqyQX5ychfgqme0OWSMxOZ2efAUJGBGngarKwsiiIZ8WckIUoBV
ddPuCb2fCH1kIL9x/oT9JlRYMuiogKB6ZycDB1MgZdPMtL0tXLSm9Pw62rM8TZzn
vlsFqVipcZjJnAX5iynvTWYHmTxtfGTMVeG98FCC63/FnYwfzOodFvf1HbFTYqLu
CGxD13KYp04P+CtxOfRbXql87DxiVxLfEVE5Z0vIywtJwZsST7rfWp6/2H/JG4dB
aRjqja9pwkSbdFFMEtnuFwxwTZaU6TAA25WkZzUqhqgGTJeSCu5Dwaeys1SFrj5A
BsVewPsTiqCQGY/0RuQTaujLTn965h8T5mGJtfP9gRZffbB/ftS5rEEPv8PnAGiH
/ZGdtmJaojhrrOVAZxAVkUCpRQWrZoBNwdxyH/KN+aQUsDAwOwbzaGqH4thZTqNa
s68hr3gf59t3H1ffaRXE+VChYD6AVtFnj36mn+FzkEM0dAQ35kX6QdKQ8x2SVM5x
7qMtN4ggwTZyW+YakKXuaiDPZJAELO8Ypm69QTzjUytPOaJdEc5uAgqN13Xw/OyZ
qP2fJLLQEAT1LZIZvqnTkVC2lS9UecIzC5nP1hjgteHQCBKWLHulQ94ETlncyRlg
FyaB2898SR6NzZ2HvDwxioM2S3b5u6tVeKBV1qxzj1/WljFu8p14lXJyK2nf2s5x
FG0gefyhippKhNimgckyZW/dqFSDAUiEfnkKXiKQU81pP1skAqwHjwVf1sVFeNFE
sYUAftoa9e//GK12Y6sToKYWduhN9ET2lZZz8pA55nl78N4MoyeK4OGIHZJwBi0D
JspMR4HXmznYxLTV/jSgG9dER2dqi7bQoCAGxBBO/ZVrSITJwkYqv7L9JMFJkaUG
xu0EJLAUHVdyuKzD09cK2NemDP7UKBF2jUwBSiicPKqIquygPpd2Iq28BRt7uC4L
tTor02QdgL5Sn0tT3yjJIJWhj9aPLg2oIP9jJhRlgL2RQFfHJQkYTglPb84CEi6a
+wZ2Drm8YiIqCKIHrmWGnObZR/fv3vYsnyMOhLk7actWYJv7SC2aWoZAMu6X5FYV
TJF/Uq1gKisASZdCp5Sxd/s3pB6JziqzeFdkLSGaOqJkCwGm9f6tkkxcATob1gHF
0YTgCGoZ5I0BWYfLRs456zdDPjsxuaPN1nShcxzNuBh2mcQvUhTj8fGNVJrVsRz3
GVWDfgdxX8V5hLEZpwdmr3rTHrwJRA/zV0D3gN9LPAIpy1xxB99Qz4vPHay6FvFP
lsgzlv3HYrnMoGbvMYMkBkLwujE1kD5dB+Defc42p4j5VXIg/8phDU8qaDhH9ecY
Kx3ebzv3dqQdZgWoNK6QPMD6EHFYI+AViPspxziuk0jifb6kyV6uku8S9jbmfjII
ftS6pHNlAaU1xiMkffsooU+gxKGHHdd5Oqmao4g7kCUhi8ukM9CJ9E+Y8VR9bwNC
IDnUrsdLB+gM0AE6DTJooobgreuwYvrzE8myGJhJxHE8pfQqGIcaCCOorRpUJcRm
dL1HBdaFT3PL5aKwZanBEDJ2GxVMIuKuzGcRxzBC0BAHuqX9KFiM8rk1ebdjoYxu
ZmifVmplMzPhnx7ifw1X7tpYwJxEli3zPE+Wpu+JXAaOesf0iHJxWLGw5Qk9CcBh
b1l1bHH/8GitSl7ZwtBfvaEkkrvT2A7qscs3eVt8XsGLhP7pgq6qQiqVpBhXxH9l
deSZ4/2mlWimjveQWXo78WfNekssQ7BY8RVRJyyQUWlMNlfoLNjZgGl1lK8aLtwi
/zhqPOx+jgDk+dWbS0ejqoEjOs9QHoyLs2ONBKnx0ZhLxB9nGs9T0TC1pKE+uxX6
YqER/avzccL9DLUVpAtZAGIrWLvZzONj+W3jeitdpYRq8io64tA6QLtbVUMdpUaw
nH6z9IkXZPSfQBS6eHlJa0F51zYlocIsDeqXah1ByB6oRo7IP3lis7XxtFemSZ4j
bdjvvSHZawTaQNwHkswyms5nAmTLKOGnEmnK1IAL6WFAS2hi6v3ke/VSx0d4262d
moBmAE2AyGNIibNAgEs6GZfODKTF2F731fMOEfqdZDV3mo1bb+B7jARvtX9McVRJ
zmNReHJO1F9StknutE5YwIFRAhaFmhCt6EaQEi/tl+Yn7MNxWhm15x+vFTgcTmsy
yaSIq2he3w22Tf1+7T3v8H3y+dPRan3IkIPJQrhDJwgRtB2jKJ+J7KfMSVOP6k/I
o4+MFMH4U3wyDoHC7OaSRneDUGetjtwwn5XBBRO9f1tzkSD2O5dHpEbf/q39pPcZ
oXj0FRjfn3hTTZEQmBfHCbBSCp5a2uvgB+2Ca6DjrXOyo36dJFmCE7NIIiCHlJWd
yvi2FeS3AOsW166ZAFgsBKV1n9UOfLayNpadJPKGBNUmsdjgtPo+74FMPvStUKtd
3Mf4P4qzmXX5tHz6JEYzvky0/zf4CTnwQCY4bdidEz3KlGeOg1Sr0VPLOS25SrbV
sg5vFO7D6gtxgUCGqx71Xt2B6YsHonKYRFnOncptPth7oOdfJmJq652BfFXiflH2
/tbBAUKj8FqIdTNbcCnfXeJlRS8ExKKL6nIcQX3BvX4qIfRGfW+F/PiX8B1vZHqO
yrNKAGgi5K3lxXMHgu40jdJDPeIteLYVGCMJ5ElOrKrje8hIWyqxVhwiExRUbiHt
9pQW8TOKyfFJjkRByG5Y+tSLASGTfYRijEYhG0vocHa20ctX4W5lr/XJxp0VluLW
kXIPHSYHge1DNxwvQqnreIQswlnbbwbLccS3amNLfGXXXHFcx1AuSmTT6oXpgkK3
VmvVIXpIliAAUGADZhBgmdnwp2gOToJP/zZwbPt5xfFKjlkXC8DjfjAvAAFh6Ugi
ktOB8p3JB0iZ9eRoEGZXQT1u8UWC+lChkSgLrPGGc1IUYfEu1w+kJ07mA4q6m1h2
vPF0viQH1+MM3z0SWWY6Wd6PtM+4K0ILeaCl4U08pJkjZ4LfJEt//FwICIyycmyU
wl2qQWoFWOXfCurBkPM2xegimwrEw+O3wL9EL1JhPugteM3ulLQLoaES4OXG72T8
kVrmGdW8yL2FNJUgQ8OcEhR5PPafXC4LVQa4T7CvvXxpgnlQ3wpe4WYCg7FZwKsK
sVVXA43CHWP/7T5WGyQcZ62xVg7eeYkQMc/veX1+MXvB4mtVFEb4gNDWalEKvcPS
6/VsVms3arQpbFGTJhQJ6yIag9J7JqCxERrJDNngDxwBSBf/Mdj7Pt/ZRXK8ez00
6L+7qvaUSfZm/EcA/W+XilYbtHzdENGZKiJaViCt/Defzmw5NmoWxzo2QIjTLKnZ
c16UqzsfK5oEK4AHLAlDFntkqyQwUvdxkI4BoOzI1VSx0pYP3uv82pR169A3NU8/
Gm2+a23fUk0LlXsgvsx9MoJFVLpsDjWctPGthbqorIwitv0VNFSUdObAbIKKmJ7R
K3T68VGqOgh30I/nBfecWDvm3VpnLA2dnwvA7lFxF/+ToSInhooqyxYOtHhcg4eq
WQufVIi530VvGI3oHwJoNXXixBdvgHvCLHn6OqVwSlsdpkzQJ4B1w4tPV5hjfGUB
qr2MG2bggjBZaPUKTW1z4v4tfOdxMtKA99cSIB6n5t3s1CM1POKUSaqrStef2nfc
EQRX4PR/L4k82rZrnFW/+QvU1sMrnAt3VvYtJuLXunoyBLhNgoXlA99tN0r0Wlh6
ssTnM8zcxUD7zM43gpHNsYEzep4/JOV01TP+TVVNK5CdIpCKILJMzL57kG+c28lx
U0BNQoh44Yh0lJikfTmg0/IMkjXFP1Zri+DhKC6G4usGWswoNWpax35s9visvpbc
D6sSnc/duVH1jB+pyt7bRha7bEHFXegiNBSjfC3EAIGfdhvuFAPjRdaQc6ZhDc85
0QtrwDKtim6RJCmPr2PvYDabNB3Mudn94/hiU2sAvCEbGPWgAyoMlcgVYhMjS6y1
y/38naxAbLBi95cdhov2sd2Stuzh8P97vi923CNohaDUZ5YtDRVXTK5+iO61iCcu
9knkPF3PjTPJz/4UWvxkLbXbYzVMNW2J33rg+/RycVcDPV+v0WE/TnMFTlsHes6R
Kj/Lkq5sVtX1MQuU/N6+eCuWI71TtH9wA3sWMjT7RCegKKPhLo3HcH3Vx16+S5oe
vcAfucXpj7+iBfe8XTDgBYWyo1dgnPY3uz3SbIDkZLBtgzjiMlRVFwtX5SYySNoV
AbYt7eExm65jo1FyOIp9aLeQc0qIJC8h+Tmj1n9UaPPZC1bgMAd4Xy5gt7I/FoDQ
n89bLS6b3XD4wPXES0MTuMuVEy29aC3ftAdtD9ccevkxnRnFQan/zYEQvKa9umy8
l/shGw3tzBuuyoYFQABY5uimEUh6hbpsG0r/dMWqJuHpr0l6GQ4qPb8ZSslMaVL8
HB8tblYwNagOlPhrBzKkQFcKlSMipOpboijCpWS364Mz0D4EmlSR71LRHpm09CDn
ff5m9Uy1AEW3gi5bihtCgxb1ijR8NNPvJZ1QCpJxxYMVsznNfKMacDUQ4p7G0fee
wk5r0x0l3GyTa8Z+QWiNNf5lLR3SpgwzAUNNjqVrGfAwGR1lSbhL53iU+d3P2rVK
xBb7HADcWwkYeOkaloug8ToMybPE3R7uFAhoiB7C6CcQZQWI3gTs0Xl4CYr6ldQY
YwfCGp7bD1TGM0oSPK8clWvR9fe/nuIaD/6dVKldkyBSESIhMz5SfWX2SZSmuVDE
k8d0N8Qk7TkIbw+PkfHc2usARuKBAE3DtkzsHucoNIQo/R/U2b8rPLjjydrz3AMF
gwMlNaDPw7qTPHsWAoss36VlbuH9fvtGFsWVbOMy1c+i1X7oIai7XDKxS0NabUi9
M8idgk63nr05PrtiZwl/rEuWlLwv1HRSETiXgrbSuSwvmfUztq0Ym1nqtVrRlQS2
OgDjQ9RnWKTWtPT543gtMvXASK1lWP8v0ifFg8ElGUJZJRcg/Xe91ajTvrKswOcx
f2mSgJ3mxXkCYin+DI+Ba331sk0OFbGdPgMypCmsY14ls5Kuh8sr56l4w9S0H4O+
8zQPwy3V/gJr3FtaR9iyyrdpzQW9llKRhXqk8/cENRfDfkNgcfhlJ8U0iRus+Piq
D7LSoYVlNGltyvjiuAreT7E772boGLuIQjoZtqAgsAnGhpDdiDx78BTshTvBYofF
ok7vwxNqQy940t58re61uUAsxkPuTtVeW+at/BzZmNnzMrKU1nYjV5KWZ8mhiwfw
OncuaWnxGxOyd/7FoEcxJv4i6idJojq91uTLdkQ9W32RlpkOcUGRMO9TuT8ufmL2
ldBO1cVTlOO8wYCkGUVOeq0l984zxIkLLit5SnXzQPSwxPHPaEtKzZLBKUFzROji
lxPXDYTO2yglRMk8Bnskt0fKVSKszxeJgPWBMDP0qujPj+Z+HqC3vbPC9wO8LaH4
Rd3bkLUAD/LcBsfKoVZ7ce1GxKtVBpnzdL6X7oUQESY/e4AjL8urzbtSxbGq1Iqx
LxCYefAmj85NkjgO1jdLLcUG8dLOc9X4GjT4M2pBrrDkeHp83H/y3qs/w9jvnbdz
ISUzaSw0cm8woVJPhCdtDCTg+m9ENvh3cBDAJ3bFyMJQArgEJjW5OzWyw83nNm0W
LQeO+Iqdg9T2H7ggzmMorJwKvS/NDq+ioEhgYUiwATCXur6u+2IO4gKLSOEcjlYq
EQDt0G6uv1nqTUrbcva5ducpXuMnCodnuK4xdFwutwddDtRDBE1TA748ZdrVYZz8
KBGNW0p6OjVTe+vJc+I/lYl0bzwVJTlZQkupt+fS2/+PVsUDowh47+C4uPHEwM+N
4cz5MHB0CU2MW2lHki1mPSfi6JFrd+CZbAcF5rmlOML3QSEG6VSg68Oq0dd8Dpzn
3Khw5fTTNeCQwTXzraA/DJ3M8sUBDvt77m9klkEN6zyVvck5JoM/rKjK9s6bKwkb
lAOzRG8PnzPDTJigqlN2c+XKQZtSw7FIkghLhZTMCikthUWTCugL2/DpylSRQlYw
rTYIHJ2LZ5sBYoglbxntmxooUBOpe38klzXX3zRnQ7pFW3zMCjrsSsC5p6l0j0MK
0A8WljEx3kSXDNVcytTdU/EwZPKxwwLvb7l/aFFTgZf6P/vchPX2TZb7qownHL0D
9IdFNXpRIZb8KQjrlbgE0KK2LOAb/0QTSPKHc9L6uBIa89pLA+vD6m0lOWYt20Mf
axQuWRJbom7lZh7ovr43NDS9Nk5xOY32LB/TmSyDyvdQ1t34tweBNn1GoLq1bRWt
z7Sv1KAUKVOzXAqSLBF+fhlo/q3nOl11w5eQOOdZIvhIZzpoFFyNtPAbdEdl3D1b
lEl3PKbrRzY5HhmL7NbHUcagOLPg3PMFwRXQHFeCjNgS7GdIbVchDyPEay740P9x
iYe/4lfrb6//4Y4lUd5eZHC/B6+UGNe12Bbp7sNVXMjbejD5Q9X+YM40j2G7Olvh
XKjaVwiBuN7qIEKXLB9tMyLxOWrW5BrmbotysfM0qxwGRx+5o4C9t8YbW8P02ocB
DxPQBFBMbvgc0aRUsE5zyHv84gav6eQIJd3KqH4nhH8UNy9hzn03TflGBcKhD+lF
1eIc0lzbg59JOLu3uUEfhWkP8L6Sv6D9TWJ1h4iaNU9kaCy2TkBg5XCRjPPpddsS
SJTbiuiuQz4W9IpuKDSyKUjqCmWTtWJyFYE8TiKr56osNXsE0bZYMgMj4O7O9qc5
Oi8WkcL+M9IbRvO4Tqk7cQ3U/QD/FpwRAZql51xdmc2l9UqDFZJyYrR3BlXUxAgO
HpHJJiYhh1anF9tH1XcBcvE65yCJIa7AIBuDSWWWrrTiW4ut33rGJcjqqseKh8gw
/XFLvB4cGMb1bvnW5Pv5sYei2XwQhRiDiyEoWJv5MjOQ08Mj8kerpxAc9Dr4kFra
tw5/UG3qu3WGN6AMv86NGZhmoHRQ05IewocPQUoijp1uYG+k4/8Q9+72hU2bdHyh
nhhFibvRK+iqOZFqqi+B6eJlKgy1OBSiYzPKOk8NBCI/uFRvOIjATQUAbQg8PNkS
cxEvfHHEJER0lwkb7NCJCAYz03D1Ie15nWHDi1KWLFahO2LI8lNv97WIswewxiij
g8QoPMrzhjhe+h2PN0NeaaUbnboGz7dnhieXxngyQOfj6+ESRArhD6bR991E+OH7
3FIUXD0uyGFYG9tripuuW9WuQ1xMwwVEfHxAT3BDFElrGEV6Dz7FSKOsHaO9FSEi
7nHTl/WqpmnKlM9UfvLXH422Xaf7yRgijoEmIzKjhjwlH2j0PKSNWD2oWG+IkvY4
D0f7iGWxanCuTU8KZy+I/Nr79uXqjScYeW4XZpZ1WFKXmmtfReGfbxa7Jpahuosb
Nkte4v6yqBDSnki/op84oZt4p/mX5aG8jqBREGXd3GBlGHuqy/u6CYkou9yGQAsv
kcMlKaSo1mXy2rzL7N/c7zvXeaYqf2AS4ROBqewpmMCyCGW210w2YFn6SVT3FpkD
w/ldwa04AYgbaUrF5KSHCRyhDM2a1FSeLEYVNJGf2v5n6QMcg9GPGnm5Mf92Ak+d
6Ck3R2v9azIpWuZG6eXuDghu+ZSK4WEhUIucUDZpFGbO1zCE5ldLuK53Ur+a2Kzn
HN0292PinkG8Ru+6t9p6h/KCP+GtMxObo9FflDz/eRQNJfJ4ZX9Z0WulCPYRnLld
2AShGd42iIofItkQI/jzCPu9mRlArUzzaxCH3Qi72eM+4DYuTFJA0KKQIElShncf
qgqUpDVGgbnA2546R5YdfdRSwXvMGcZniIhFNE41s7vsul/OAtyRvZXBGHccC7Dg
dtN4sMiDJp5jTdzkwa2SgqJkdnlKkhNPH6IpG3NUGMiTnyl+zRJOtech3T8iQ2oK
FC9uCC+kOR/BbwqX6G9G7k2BPItU32RbbJnKsm94Fss4YxksmJvs0j6VldROgG53
X8A8HPwPnMnIT02/Fvyu2Jx5Hqx8YyzV3nbq9fkHxWzL8/7aqu+LhONhVmTZowoc
4fkT9or4A+wyT/sqxuCelc58wsL8pjUr5gHQQnvH9T+Bs69aMLL0L+XWp1ryTYDl
C7XlpTR/RdEL7w1xw3T8AbSoiStJ0m0kvccpOcavmw9zZUCLEPzmgK34QWPRwcRR
AoDrAfT/sNu2erDmQCFYpIEhMChNSaXYODLtVDxWWa6ThqqJI6CJCR4s0JMywf22
MxrzFrtRft5w1OoBhgrLqu9eCO4V9X2D8Dq136gNmQrfL9ht1DD8KgALC1tHxJym
kLT+W1ZKQf15dFirTOe+Yy/yx7TwDu6StlDC+ArY6fBJ7YVvvtA1U7bbN4D9NIjJ
wZklIXuQ6lEqciXuoHi7WxQx+GhAwB3H0cqTqQZU/E+DQHtaOA6c9cBLk2ve2Ao4
t9qhqrWGWyUfdvHdgUTxy1hGYuQAG62kJRgAARdTQeXJbJdDjkcFMQPj0tk34wpc
TLe8FVNoaANai2b4zSz2RdPm6HLGRjW206PuZnnoo3tHYfpccDEo8K2BjpwxX2xa
cOPm0g0x6ekbKayd+kwvzXXxNPbpvQCuWiMcNCqjV8w0a0q9fIpD5kbjh/H4esWQ
LUGAGNBSH+IJA1VoALpASw7TDpV6+QaMBcIy+Jq8bTOyz18lkEHKQW/3MckZjpkZ
rVksMlE5UcyJ2jYnhUaYY7SAbM4jhTTFn2v4ak3zJUiHXc4nXUGt7r3yW9HdpdyH
rH/8flQ0zNWYwwM8r5ldUKSWAMV7rfHQ4j0ZBzhWjKWFTo6Oc5VWe4EcxkrJFIZZ
kLZMLA2FcSsdAV7osKGG795wNEc+RpYBxoH4Y+FDBxJTp3ZgS6djk1rC1F5zD0ch
lIGaDrrWez8X+hMOO9Ik7rOt4mEPBlMTyVPJToVigdNV6Gxzid1L4Ma6xfed1G/Y
j0wAYm8nwzBjTTohS+hQ9IbJ5IzHyWdFqi5JLqYfcmtxK1XH4toKmj4H8ZsCSOtC
kXMJS06Cjy7MH518BxUfmHFZfWc6sKl4B7B1K6aBkYf7Ezyc6dTuNGAAPS/wEHNN
m6e/mad/or3yCq64kR0A+01/N43Kz4pmnZ1n20/8LMfb7nBPyUtYDfV6Q8+3xOYp
+1v14P8WAkoyboe85RyNe4SdrvvoaSHExByVOd87ECeRMZhl6V/Ns1oIccZcOdQQ
5DAmIm/S8S1k5XWcwMR9sCsHqzAbk+86jlZApdwmySEKyKzSSv51rIbuloLwo8fK
uCIw3CvlLdWfXjE1qZ9XoksM/JAmtjLARSQ5oLfBkgG2UgEI9jfOoTMavTC2RExQ
Lgq8dfi5WJPWl58kMB5oh9OA1hIgAIL8uIuJCKwR5NhkjrdkNcMvoOTIciFmXCym
9ltom6PPSU+fS/7VjQRvVXM+bbBQyi3FPEQK7z1mMovJX1TD9Kd+3OMdJT40mC+7
2ZABZc1XZsnVO9jRghf0ZZdBL6D1El62g7gnDRuW0C+MVABH2SZP9qM50Y1C8vE9
Ng+YrcYd5pbcMgAeDkvP2KbjsZLFFFo9h+YmjBu6+F3Rs1RJkK1j8APFZbkFeVhe
CK6k+CQg6ijsOpFOeYz9vmArfmkMGwz54EO3q0be95Yq34whtYC+3MROkRD5yoP7
Cm/v17Ct8hd0VBocJdQ7AufiMC415ty7RA+VGULk3xrLztVjW7inIXHpk9r4ZNbO
1JbILO64ppUtTQkfJ7e71sdvwxyQOaxwP/PDQgKkq592rWkw2wBKJmwGt2R7JEDR
oy9K3IVBAt/w9pDmJ3Dg/lwurWDP52orO/5iHpSUk1j5mzg00HgDoCa6DjdEJV65
r71yhcAuLTrRcLwHlQinYlv2wO+/J3VhdeE7zj3XTVvKi4F7eGlHA99Sa98/dOoF
Anh6/wloA9s2hH7qn+/OU6RoyDYqxrCWNlcpELy6AVu522WnMhGw7V/rndHqsOUO
sbuYgwW4ZFxUTIpWBN5p2UJldDouEwnlkqrVhjqFik3+p5TYFJ1/ZDvewYD9Dibl
Aoj+Urf7sROBdRDbHQIkVxesgyrUk01PtQ/Zkf98yzJedzrhnEk/eRL/fCBlo519
VDuEFsdpLB4Q94we1YrvCO6ECyXAl+1/r7gHzv+gnAxIrcMrZU20BpSeuAVwHhCo
zAa3LPPn/LRr0oGWe6H83pEuRX1WqVSippNOL4y1D3ZNtdb28DHyqRuTXuC017ho
meq/tgSll5SGGm6z57sDjX2nbc/fKtUpcmHpfdtNUTfEvFPLTIKFgc/bU4LFKtuz
/cVxAkyBxg9wn9hIEisi7mkvzdt2VCpfKhpOZc8yEJWkK+xqEocXMie3gqvkBD5Y
FElWcCbAsjzaRmBVdNfsXIfMEgG41V4JFZiLcTmcBRis9fdCvYqAohUl2+N7inoM
6Z/fQiKKg/si1rPTGHQWBhqAcZtKYTOQZkdivHqZgYzafdyUP9e4nBJmGBHit4f2
rCshpLVJ8SAzmndyHegY+h5h2YPSFuAJ1YS5MwNG7IoVoYxdZ1KpDYrp7gJqriTj
juyK3iMR0TKLf7Wi4ZRro173qPuKGLnU4/nEgBAKp9evsxYe4HWdJtHSC79hJ8u2
qEZdGSLZtxDISpfADMobCj7Qqi2o7VwFobHGa/GNE7gJqVxiKNCnpiswSz5riVfY
OLSwrEbXKRFsUVO2fFMYO5b+jXOb/008K3SUs+oEKNFo6AZ2zBa98OSnwgpC6uzB
yK7hsEPvnZz7HpvPJBhrdQoOflnyP37h/FgwfAlvR20MB+jiO6Ci7MnR4mb+IC+5
nNhw5azXBJBS1xYJlEQp5hvUklJDbPzZ4gM041GB9ZUaCEimcjZR5AUc7MHBJnT7
m08ZJvZh9qppqDdeMucjr3JNypJ6GU/l2QmtGMI9Hbz5vwSf/8G/DB+bvJ44nPYT
wPHYHmI6Yw6jBAazG3AD8OcFMv/4XhP+tosw6e9sIqptCfnL6/U2+66kCGgfmQCl
fQUcoASuhWn7IKhj2DqIv/9S62jqD0QPGLjsi+kWFYBJ3UxnGuBqUvgKA2TeGPZD
NaRvh3kCIpiIdQo6FFdKbm/cQGeT04/+7kUIDWflQuT6XI8bByozw4iPXP97G77m
SR0VkEQ9IbLUZzyu26uHhA==
`protect end_protected