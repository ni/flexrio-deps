`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
4NAZGBPmQSC1EoH0Jm8NyCqlPLj/T1x3yGUznZvPJcSDzBAzcFwqXKRpDaH1ZsLt
Vj7PZwMXoCrWz9CTK8Bc3KUzczrghOXYmwC8LOjbmsVXpGI1rGhG/OFRuWiM8K1L
A1bH6M7CQ/hdNmZA2hrnkO1xffHSLWp3sOoRuYuoUzGtqoiLUyU2dmf47X6N/M0r
/KgfS/okM33DGCSRGXD40+FiK206qal0FphOsdNwNyEbIzBpV07uJeFMRpLMhJ6W
LlE0uoYVnK8g5/KsSCy7Tcbm8897hMGLKtFDprC8T0qYZ79dXPaVW1c6VPm6z355
eWat0S0CQ2JS92rxmGytgKmp4/B0UbqBOAA1EKenPxOvgjexd6Oy1Ps6S8NTtk4G
Li7ry1R6b6uEBBDZGHfCFXtThiG+U11YgggfZAp2C3xBojf/buIRcWXrkVm35CIl
qcgpifAt411uA+A7avqiiWoQdKWWdHMSYVAWaGZllv8Zy30ZFl9Qz4nEc0nx3EkR
T5BJ4Fy8ukZ70iariokkxiBXEj8sBskjCO9zYDBYwcDjFcE8IR9fGdRgegDnsQHw
fAfTcRHj9n8o/lrGe5hCv6XaTHwURmHgfaiYC9pl1wm+BA9coyTTgy5fVqMJSD17
ZXPGEZNDaLbkk9KnxvtkfmGhe/t6GWBeRFGN2wnLiAoe1CJB+IbChQfR+KoGSgQm
JIMHOnc3M1oDjpv60ZmM8hZVSEoQg0gtR42paIDHb3fSWtSbBNf0yrAbIoZtUyVj
TgQvXgo3KHe/rlGKbnZqqPEuYSHqY68vdFvQEmLu1G97w+WcYfFfwrlwkTcSSBYa
oFo72/WPGsJu5XP46fuEK7M1YTY9JaxqkNhW0lHN2SkZ+UfF2o1vxVNPoPCxYk6c
PpyZXCPN3fuCvXaxlrFIWKif9VfU/dz51g/cCDob1uFnUm33o6PnOPWv9iJl3x+k
paF6vQvZyxr8apd6/6zBt+n0pIh/7KV6K4KqaqTrePFTRwQOiWW7ACfBO50JHGvv
GRhUQWk++tTctkT4bkxdI2x6imti37uN81PmdrYJjy/anvyfk+oOIhtAPKUjC13p
m0WDY5kLQRyOlQoyUsN2iDJCBLvaNBuitFBOL3H0FaRLIl3qxa8TjZof0dbxm3x5
UN8zFCTCxjrLsArYs0QHo8/+o8kYaFUH7GMMbMXQnLfD236Tz2YHXxBwwpZP3Ycd
EveY3lLO0UXa4w7uAYMuH0b1bPAATNGcgnem94bXHvL8WIYzHPAS92mfBlJiK42r
H6W0ttF6XCXtdLvu0+IZGbc5jiqExSd0xt4JRwcmozoy4DNB/F+gpge2ZQCOQ3Dk
ISKWozDbdaA8+qGkYQ/9bFVdclv2/4fyByMBSSoZf7J49rQX8e64/1Td8aJC6SQL
BW8bWtGoJk3OLWZFgqSt4M1qjTu1hh13XGElbje+Klk9Oit1Rvl8rQai/kwZD5Q3
kMmWmWMERQ6B9gaMo9Z4UBM/ZB3LYn6AQpRtbIHIHoMi8gu6IFfxenBfV/FfpT/s
4Q4Diaov9suB4mSL4vLFnAAKrMfhUogqILqIjPeZQ8/GwpaNAWjspgAgYqmLvDMk
N4EiTuSBo35QXyEbCyHzna1HZObSA62yZxw+uGmzc9owdD63weYj7kYbvax9doAp
9rOrA0EFvVHCF4a0gSy6K8Eh5KNYXILBZgAo1obTBuSRgZslWXgs9KV2FZUVNvP/
9bU7ZNBcR5Z6dttUnN3wHJPTWPfl5oX4qcHAbZYAOCab81UdMa5nIPT+NZvhbcWT
kHlQWGM0DLWJXZ0pVQ13mgNmseEthd23DhRl2DgrqtmuggZ1pUU9hEjGUT/iir/x
o0cndlttjKiinPcmmVXFwKd7pKbCmu8WMb41x8m6xVCSf0AiQV0o1SUWVZwq0y9R
3Y4CgLUTCJMBbjPv2D5f7JdDBc5af82x++hHEG0z+hSx5gnAUNoB4Rf56IsLIo7Q
sOHTSlYY8Eaa8Wr/l2wC3uVHqhfguV8ZfSr5lXfB17N20ACaa4CMgBpPFvLMKM9t
4ERy7Kmd4e3lx8nFNJJP6fMla+1fO5QAMdKVBwg4l3uiAsjiGLTPMf6YmV1iyuJM
21zAKcouYLCZNFOMhnpzxvgNoDbe7CsZotUQu9QLVQyPgqz66CtUQU1P7H1KgLYj
LLayRFNvZC/2PGUzMm6geVQeP53b9yY9PJcj4xrMaIFMJoe/HARBrsLt7N86SYnv
XZVRLfjLBzIgWdcdNjfipvcgpNADJItuRqFXiqA0sbiiGV2+Y7ICObPmSUzvgj1X
CBG4KNriwPOXwTGQRu2SHkhfHOgJncUa9c2pKFpZxUovtvTfjQbBrttycIg9feai
CKO4Gv0WrVO/SMONaOBmz3x5fLEhLp1pFeG/6u9jp4ljM4K2zFTERWoN2EwC4+Eh
bobx0LuiPh4PbkU6A+AlnSyqbAkNDu9lEx5c+LRy3Qd6/DnjgC6LbtlKQwoqhdXO
YbZh+YTTUUGZ350BaiqkUjvSCkzm8DY8clwOpo5znrP5SD2Mgq9ceOUKvOd6yChJ
P3HbywV6akp03pm2Uo+5puiRKATYCVJz/4RJuAzDpuES5v/BwrzLSGRVt5UhvCS/
I2BCA6CetUb0Y9FdWdr3UdHVXdNHwn6oJLitODVQEdchFEEy2R9juGmfn7PdH8rd
N7IpOU3bl38XlToOGOTYHqjPlMTr4+FD9Gu8cQ/r8EDFu/G6Q97NxCF6MsaaUIpu
Jp065XdXu976pHiWkS2uQ8FZz3HTuWeRfXY/yE/67yc0Bj8ZQx4xi/NyB4SmQwJ3
C1UA5dkFiuiOedtdpC1ygr/eVRz1Z9SixY9KbBEuzaEe+urYRtTpMjAJgLbmupay
2aIRoF2MWOldBSzXVWWlCXbQ3UchUWwpZjRIxZzQw3d5OqrfldJSyrMHXovAb+aO
qaoDl+T8Uj/NE9aaWEOn4/tcFrVokAHuPkr+4n3FLuzVnV/W6h+KM6exYi3sdgXf
ozgq6l7irXa2Gi19S9jQopqh3SXlzysebDhTD+2WXUzj87hKZCdfsGLvF256pHnV
OldP7hoJU1/ei5dozGjbF4/MZBC8aKLtlLqtFFnS78w32nde2USmeteCAaT54crv
triiNfzFIwNjU9wTRLdF45Xzj1bz05M6mpH8p1mG8ayThaJU5Zg0l3o8w7mAVKmA
VD9jOGzJO3npW7gDuWJwxNK3ol2L09IXkMHkps6ienB/qcmcRg0pnQF8Fk2+pLJl
cR39FkmcWDCcXK4tFdjTCauUmR7t5FkB+4ccKxLim1hFlV3SUdC00+66qV7oayxy
54jiakmW0xhy+yWreBlTE4F6h0xn3iZRgsFHxefPVlbVahMgdHWoADFVcvctEerF
hkW67vSu5O2Vw/2qXIas0WA3Qnp0wQxkjvlU5Q8NjB1NDxXU403Bm3RzugAFbAbu
mKYkGQGT/GjxZL4NrK8lSD2q5FYKw+/2wOjFMeFjf213IW3z7Fhu4f5UF0cIaCnJ
w76BfU+XyXTxD7706gtuSVqd2lZPROKJWjYDJBU/ASGKrJdDebipsA65r+y6IVvf
JZiGF4tx57jmTbzi3GN692Wiqi3Q25Vl+scaqynIcG+3p+DjpJOMcIHHSw3HA61v
cVe7YQonq8hgr9nN7ghyMncMMJ/wLAm7FbNgZRgKIHWedLoeyC9dzxJxOaVaz6PI
sND0C7/A6rwBgQAJK1k2IwtzUeUI7SD3qY8repGaaKM0v1CRqL95M2KwE1Cind3V
yt01kc+YWN7L1sCqrl780jMfeZwXr/UekuAuUn1Ho/sNMrldxpEdsSZ/IHbEupsh
RCIS1B2MNx29pQHGtCOMXuzvjTAaCOJcsh/AKN463Hq2MxVKrhj/tWW6AE8LzY4B
+QtVAt1yi/S0GDu1mH7IhwUZRJU39jUIYvSzZ9eq4/Dm2xT6u44cWuf8gTmLVd9Z
RXf4FvwYLe/QF8tkjmxFjjiQdGsJif+EWCzUZ6E+T1Bbx+8uFGsBw/qPIViNzR3S
8kKLB3DPHSWSgfhyJ1g6EBaSDz4DVLuO2yNJxhgccQjIh7B+H36rz0hmtyE4t/cV
7UqJAIgs9ak4uWGO/szwI9tmPNqIpsN38MMfV95otnskxNuCFMY+YkKHyDhUp/xf
lIzTLKnhOApTjL7QDKB5hNKXN3mGt85AtBEnNELSOjcfLVVQw5YeKtgrbGZNI17R
PIJzP0YaZFje3aUM070Co9MzsnxTymHt0Naz4HNFgxCUIOYc/yeQjcF/65H8Zuxj
PJxm5FraFGDpkyrbbCHIuIwrrQ8YzZzoCWPalA8oFA7sPuLEv2TdLvbIKSKATx1+
O0idOPW3rHvtMmj0pTwzY5NHzubB5SDIzUM1pVAFhILQirEuCCn6hvi7Q0j6SXOz
NGzpSCav3Hf7AeFc62tIv97TxLq3Yk4IS9ln+vvTZsxzdCe3TR2aljH82bGZJYgt
vEmUfKMoKmtLRSM7HEFWtmgD3eYbyDZdGBUxWPpgAg6cSnvfZuCQK3iTl8Z4IKM3
IpXErUg1ow8K6vZ90G2EgXa/A1ddpMSwZ2yy85/frIIdTNh9lp494TASbwiDMknI
UQg/LzwxB+x7FTFeAblAStW/2QSjbztOW53GIFwkYhtf4t3+AzWo4bKS5ibPS00w
kaezctYAqd7kUoVlY+LRNMZWjAQEefa+UnD4LKs6V35zSmtvwdo16jDuH5yNuS4Z
F2dilOQbsZ1/cZ1gCl6gByhcS+tCDzo6GJFIiNHmveFRP6vyRzyU1ibW/b6Afryy
pIZX0m4tJKXWTa0Ep7GhPJNYYuISBH2hKERAWF7ISJxZzSHE9hA6Ll+vQrFE+Gch
7XKF0MQnrUl14/Lya+fbF/YpcXfEFftUh2P4p/VhRPf75JsvPzuaWpp0FKkjuR5q
xHoXlxIWI/QybaBF3CsrJIvkkWQHwcjnuFJqZpW8o14nrpEX6Wf16aq8608R7FU4
qmStqXQQI6cA9CBdHGD1/G5Js191pfWgHPvx+YFSYMo7436aAokK1RskzgLddDKm
Y4UmTrxBS2AkBxWP2/ZZyph03lXuKgEaWyDBmxoth3OtNW+Uy20MtaaT57DMVgYo
lT6ZNiyBABOmWJJQyBGrJC7Lv7lfcqEZ9Plp2w50xY08TsveXLl8T7SfbXjMAdUA
H30h9XV90oGzmojmENW97V3zI1IxsVxSSuG3/GaaLwCunIT/vpp/Khth9WY2bUWb
+LqNPz7qnyPMwLeJyg8ghxqc2UNeeihISwiONQT65Qet9y6GzfLV1pIplgAxngzA
JNBNO7fXYVT2z7Pv9UhADidSMoeOUAp4WtMVMwQhX0loqPZSel6dSh7H2ryBi9uW
dSz5ZYFZ+jC1DP9YCrbNGhE6huBHpVQ25/buyPmUC5HwVu5n4v+pRh3VXEmy50vZ
UvgPXsFiRtlof9iR0D/Ebth7PJG1R+9io11umDbM/AxI4ny9EMilF3UvNH9bORj6
oIHVYdpilsEZUdXf5c7Ng39nfO1zQTeYlGxC2w346HlZUYf/e7FJaPQDqmLI15OH
wLqBkylxNF2TVSKpXlZl95tHH8DqqdVYRsY5qelC8UOrTz0rc9vC5dVGbzfSVttr
TgvbWoBTI0KlA8MAu/4jqEyfRM31xQSfFGMV0M407ThcU6txXvlaeG30Pt0caDBB
wJ6OnthcqwwbTsPy62wFIf2y1Ubte/Kam/+OkF+VLvYtRqkFbkv7s6h6T6w7lAS6
V5p5YEL9mQ+VOrQO4NQTpUdRkcHpxDjy35YwtuzufA6Sx7nwCwpDaLFI1NElaJFb
969+YBKD0O6cU8kw7k2K1o618VanSg6GXTIsM9tGBNvLN3p5j11sGxJhbvbdWzh6
vwXu26rEuY9GdYUzSe/3s0VUK/F4i2CpCfRULj+PvbLOjKxG8qhQ30D/5ThaQKn2
Fz7wtnv6kblr0FP7/BIqL4UAYEGYnfBAnT+x8+Lcm2mWTqeA3A5YhDGOo0uhADvX
S0XS+lvzmgxCrbbS0gC+y4er+vpOWC6fLBamWD56LuAD5IFOgCtNX65FmRj1Al74
7Fjv0OUw2N3GN5ItdLvpd79Z5OkDgXKsu6DPwW6zArJ7Bfyk5cVq2VfC+N3r0C7T
u1PDlpfxc2AiJeRtkJPaK8TaaJcY3VqJKjd0HQa1j/4eL0KqvY2hdGl2iR4Um6wi
P9sgJUjpG5zuUKxgCZx/nbBRdW2JCdhHlA/el44XHAlMf6RkXuJKjLfqlUuYIHlf
eZaMpGTaZFwYHwVcrGwDtj1pACDp5mcZmTtnEC6hjpnjfwXtdm1fAXXPPP9Ply06
tAfeYlS5GoyRVlG+x67CX4rJfuIl12Sz6YmPR/qATgNKMdX8UVCWR91LmygMd1Lj
oWmPdW1T7YoGR1+cS34LyW1+uvClEGVSySc9bnrAVrllvxcRfTHl7Ms5/k/veFV+
7/r9ELbBT54B5ZothMF4fMVhuNGqINcW+V+nXmvoKuESfNzSKsdoPkTxaWUoienA
FH2h22Xp+PC/HdZb3o8RqS4ImSVjT89uvv8gpR2+h1YRpvir8orsnVn8wjpojtFU
cfdqUj7MKL1SsaPUX2YIGa3Wgg9RPy99hypHCxITd8dWpfMyg4/PWQwAibHeS4gP
S4NfyzolGu4vXUWD4vpETxBMK29QQAaFo1z3K5KHlEt1QSxy2Cu8KIgO05QDhoo9
Ww/ZXbDGPvzz2ng3Q+aizioiD8vUAMa7v5CpndX4sHX9s0SzAOsDAJSpWgNUospJ
iuzObS7sceifhd3jsfF585mVpzYM8RFB+WfmZiqL2a1X4J/4CUUeyh29g+N8o5t5
6wJ0NlQpSsiGAASSaaxaq4GUjWE+4jkJ5aBGT4iuzpPxcRu+0AvGbUOvuvWUXtar
O2oub/smQisGvT8+KfQKRQk/HpMQBBPA0JAJDb5njlm8eqqF4eqIX1UG7Vct9bRf
qgPvwuS+N+Y1tuNvqby7eBw5Z6iFqmy0bBZQ5JEUErue5MiguzIMN2yjO0XXKSyE
wuRlCXzNr+ztqi06aHqMt/EM+nIRt537v3tYSf4ii19zBjNTMZgFVBIXpxccon71
QuPxB2106rLh/qihCzp+8zIDAI9cdEwQTkTqvnywKjRa/upCXpcB2ZE+c5R9la1f
/twAuH7pqhEADcHtPeel0aAfVicjGezKqoecngmwNlqxthRiTePvyfLQX1613hF6
gS+FlrXj08cO3dZ+mmvkZ16fWvs33whWjUnxR812TJA1FNFvC4ah4dGzyaDyQEqV
u0ewd6WmKDNgK+mAeLH2XQuXBcuktms+pSIHKrMjArJH3VjOCbwV1YGFCFjzEYV6
Mab0V2OeGZMHrzt77obxuglRnpnKLSbcKSsUU+nqWqVKDAg+5IZdl3QSCO7eikje
VXWUv0L9m20gKGTo8BS2tL9yneh3qHbuy1PE8plIon8vh+tM3HOMsR70dWdQTw9z
o/XXW13RmrHZGlrqrpfAeXDFeBJg4GGtstc9tF0d8VgU6F4fOBR7hfShA3U77hjh
Uk5gZfdjkdiOqgGExBNRWCG5WqwdNr0jpasB8X+489s2KWpD7jjXXnXUqOSGURWw
geaJmzFd7gvq0ZKlIBA5SUfl8tVNqb90ApNFV2xxnOhFdtjclJFhAbQdkVmdJfPu
CR0VtgXS2BIR+/a6yxI+eMdy8SIYLjs8xly0rFylaB2XLlf+N0DA+rkrFrd0sZVQ
f6rUJGkygVJ/wJ9Wfri/+KBvLGoMfXPkRkwe573bwyvUVJ5k9crncBw/3ew/z2Gg
6B57rv1WlZxzb9g7jta5qZW4xI0XuI1fCwQ4uwe0Qfge+btmkRPGl8ihmXoe8KLn
A5xyx0tz0fPmSXcdDpux+An1Lf+sXch44F6Gc5mHw34HBPAdnDZaJxvNwIMNROZ6
2BLvwNDDoCuCG9b/08UdCjJmJcD4ZRPkufwE8zFSsb1T/nTUAM8HF/TuaYs86ITb
uTTHjBnOQu2gdtTaCbUCg9Fd+2FQ7Ff3vxC88X52NulwSiJa0Y46ZN77OkVq3krx
Qv4rHgMUCkLICadOsaFXsuOgVMdeToFF6H9EIl6BKy6n61BirGW4cfDSqkBVKqqH
e2qgw1mzCusZkh8TzeStAvUt1lhxULTb/GohBuY88W9rTtHZ4DFlV2SEhOIB85hR
jgMreQDhbNQ169ZQzu0Et4+u2kELVCY5UyLsHmFn7BDl83PoAvF8W0GM0rA3Ee60
QGVF6+09RUO/WaAkTaYNXPj2Y0Hxiolw/iRK4aU2/vgVBaikse3KyW0NeQrtfarl
WFp7h5n+i9mZohsTXhlzEQnI2WWbIh/UIlULBi40M/hp22Of/rSBo2u3RTAZHT0H
GmhcRhi8YWFh8PDyDHffnhd5kHfTn+W1r3v8rKeoVO8zDCSYosdoWOY+EdzuYR03
8EWQEOBnEnzyZPJ2+9ShG8hkA28tgIuoIombH3EGRxVeJPLt4xnqJsoSHwezIlQD
MVtiTizEf+BxnKJqD8KBsHBS9S98dFNtmAiHFRnDU2Hb9kfSWMxX8ReuwD/HNIuP
4E4k1yvMxV5kiKeg9V3Px6+n6KptLb1a35AXwVUMo21i8jkeSU1XbKRtDrhzDeB+
e91HIsmw7KEGY1KWmHPJQQNdGLggFWOYIS9hw66r9vQGizWymPqCJEEprioY+I9U
YOaN9XSaYzNqhEgogu6iEV+UyYSGdmI/WjdRxARB3EetHSN8NeID+R9k2qSg2KUp
g4awt2TA2E7mphQjhvpyrFvMMUfmsSiyTDk/yDKsBlcv6xy2GMu72e/QkaiTtfTf
QCuhL1hv8UiFFbZo2aXbX9wQoW2H8MWHxkkyBbIgGnflaDMZG/L7bcVS8sGZBWjP
5sP/wmF8PAS1wCGhiGTVypzIKsHutRS3t7c8u5i6NXyg2DxYbsYrxkRICoqypYdQ
M7TNQ/EjyamKwtouXffRWOW2qjU/6JHmgdkWPSZiLMFioBc/oq3JHYHB1ymmV5w4
RaHYghpk3m9bV8dZPDE1NPeY5SukBZNcYwnJ+By07rm5zX9TLBxzXQWgwMGcHJTJ
MJAOhUgYOjgo3RHSBva7XTUZg7IojkRCcgdRqrP54wnxF0z0wYdWoZz14fE12d3T
N62WU495+swJ+19ykm7sMMPLQLH+JGCnlkEKnTrl11m2X4A/Iex7JO/PaSrNerkY
aLkUdO50UD6CMVnzjcuvWDVhlDL+rG3EM6W9kCxB09TRwUPLrdYN1p72exlJc+aG
qYfnLli9gpP6M45fLzznR9ayL0yNO5uyry9amMJfb0Fywk9+9MrbL8Cdv+GTv+dE
3uHjsH7qfVghk9/lBRdix1SpuJAKHGOBRfrXwZi/Xnek3diV4pdn8LoH8jGZ0Uuj
RzHqwQjvgAo0oaMtsRlvT+w7uEQFuhCBVvIx+HEDCpccJmXS/aQbNZqdHNGNDLxF
arBjOnIFqIRzulPImXAiIHD2/LY0aqLJscp+bgixLPlu4xWt5F8Fj0ozFLk+v6lv
2wj/BLYVkTgcMvnQfHzIUyKJGj2FOQhPrnqR1Q/98ejqioXkhVWWD/BAXqflr88U
SNHv28VZWDO7214Mrfwg8qY16Aw27GQY7if6iU6hEddBUwqGA61TF3wysca5Jf0s
pY4EJnKXvcjusTcRK3YUV6e+WCD7hHRwj4aTbzLpFiyVcHZI8MELb0CRnvDWd611
1EPb6nOSMiiBunWHC+z2GNaSHxuau1U0DUjLfjrBgrev1R+Rs/XkZ2aoQ/90nSJK
vn+PK4236wC9WjlhrvWa73JfVmndOkTZ/j6QGeq5OhcCWvEo1b7coqGo4OfA2st8
b2bJmcHXxfwSqVcSM41w3Tu6iDMD1vByVSduI+cdqTSDk4nUMj5igOCUwi7oN6EZ
29uoGKAtIcrfybOSyNzV6g7DwD3hqSI2n8+C0tItMA0gUguzcXWMeT8vvnC8Orl9
X3Y5/BwEsa2sZt54R6gUk3M+3y1qn3+2C1Vh7qdUnnYPQHci2qjOy7H9z5UUoRkY
mo90Bh2BuENI9PNkEEwFzUh13334+A8ZmI7kbWxivKSRVHK67mgArP+3emxQNR4j
LPsQNL4iDNEU/E0u9kCBqKfcN7FsCXj4LzjMmvSMAoYKebThCrwOVw6YPOjCxqjD
hrpgMf3K49ICnEP0Ab044m52Y5UP6cd7ARnBY5XE8pRUojDwcHKC94G90lHIyTYC
BqCRs06E9V2mB4lTQHJvnUto5WXp/BSwRfkJxQSgzYagKGJbL2eC4ay65JXWrYKv
T9esUxDB6LbQLigbwI0di31xGfkI14RdGWbV4wYwIYxjeYfHgkvxcF5q9m6q0lcn
tXPrxWQQfScAyAy6SR8km9eR6GGD+3swJ5fKB+OE8l7Unhht8bpxoistlL7wNHux
oend3UeVGG6dn2ZFHMzlj/UJDMWvwQQ63S9z/DqHzjzpe4t1qpfWpSTHq80killF
8BlO4g4AYEhuwgyUrOw9xYFziyNj8Kdr/o7DGiHnQu8KskMwwu/4mqzyYucFBF5s
MTSEMtopl3LvQ4FISY2ArND1+hFmjwS9X/t/yRielaIjCWW89TcvkuC2UiE2A/hY
t2q2hYZWHVFCz4qIhbMMwLyhktOhNz9ZjQ5Vs2yYUVtPZ+yNlWmvpZHy5NXIrlus
s3iQ/bhWeXxUAkIvvs1DF57yyA7wmSqB6gkwkkLwveOmFXyUFAwmkIcTuK2oSoR5
Xiupy7xjnYGQwIxnDYtg8sus/UrckY1PzfCk1FqtjI9O4kUBNXPBnZCg3FtTm1eY
72kQ5slre0TIaa1Iz1yDkvZalnsyyvur4MGc1U9CX9l07yk8npGMsWIxrddCzuUH
NA9Ij0XCp2JsSyZHmFvKhf3i8jARdC82FiDckzLx4MOkfXjLGG1KbJySQGYmXofs
fQuBSL524qEtwStD98+8XPZvvcBGf+NWcjXM1Vd/Jv1zLaM8hPQH+PLFi6V+pnRM
Z4tXbY/N/KzAIUZ0UQYxakR3nSpV/PgDjRu51d7kaiAseOWB23keBIEwRHIn08ri
u0j197tlYhOtT8dnUhFmC9qV1Q8xrpEwGIJ+SAph1jCHaoprfTH2s9q7Y6JCQs9f
bL7mUXH8ocLWryqKy5+THwYAj9iYWEwG9cr4GgZCeBfrzcbcTSh0F1rD4bhi8nUk
RVCADz2cPnmgI02nfQ2p1ZUBZ44yPp3qcW1TRjInRePRC3lI/UXg5rnbHV+wtN11
90uBl/KVnzlTIxjmdCbq3ZdHg5Cc+wNSw+4ZK1tUJOASZXWVzRL/bqOU89GKivx9
OJ1oc9gE0kVKYeFT37I6yriXro+bZAC4JZK/bPeVmZXqaQXFlYBiZw9Fu3GN4SPk
YZlFvGvHKFa6SzZKXQsjcP59RKrd6bGPOEbMyXPQHn6yxnV6xodgdZBb8o6nm8W2
oSKv7uyMJCqdb7qeX3/Y3S9esEwyqf1hgm0UbQXeZYMwXeHcJuJcjgjaaAPZv3/t
/MAiLxqsA7GK6GG+N1yqQkCXz7cMahj6OUbTtrUVYQjSbytWxkoHgR2kqUtNfTaJ
Hb0Jdjv8lihZzTJNiKitMxnRwjfEMJld1BteMlPWsR7MNo8h3xb+6XrJKT7aStEB
aEWqNMzef70+VLT49pdJXGQhBViDJA6cuXENogrFbhMRBr6ySdU/7o4Y3ob2e0Xe
7vd+eqz6M7ObJ7jUZDTG+9fOHImx37Jm120gzkI0WG0VHQsJ8JMaTFqV4S9A21vt
3OXQVtmiziLFZi+RcSkeGRTuUoITw0Xe50Lxv/TPAgmg5kltlAx/7ztV3p6jJ8TV
Ti6K/0g97wq9xTGg9Vq5tYHI/jj+EVLkzMAhgX0mBkaLsXisnUdC80MatFz7HAc7
2RXgVWzgVjRymVe4KfBkXpXKSxyCNYOphPMRPJPCcBWnKPR6sP1l47eVQApXdUsX
7OvcYJlxbNViRex7HXNl8eyAUMiXHN2+Ol7DFJpbdCbGBzxp3w0DkVbxVGXb4q43
m78Xy/it5RgyTRYpxT5/D33B+KbkQXHTWaRDpifZOQCwO48UsxyfznUMtY9WDs+y
tYhq3rUx5c2GNECBHTQqsD6I8ZMX0Knc40+XK3uff2Cw6w+yEjLsdM2Fy5CEbMTb
5l2JOeEJ9iURYV0VUc7Y1X6tH+rDWyl5medWeIWjdLDn/T8xezDRT5zZCHg6HtIN
/NvMbVWCYs4+nO2/DSZTXUk6/KCZMbQkoQ1TWQoTWNQDAY7zNGVBySg3effubhYr
oYI1IS0Q2nIeyrffzr0HrMax/YOtTbw8ac6SE31jerpZolQFEfzktyWcQKT1RPbw
n1aeErmaJ9klQQgywdnTYUPVuVs9PT2WwKr2OO/4YGIpW4jR13slWEjHU8h+cprb
GjTrFQQTkU5yss45PATRUTcj29e/XtxRGvBBubkaiHtwMMap3BJcNXSkMpSGpk1X
p+qjXHryslzdf3tjmyr+Qmv8AjbPSXXbJS8Kamaio+6FEey6aaplHVdSbpaeaqq1
yNYoTzub9L+s/V1l9Xfx+sL0gOZhjOnmh6dNdpd3WvNQiUDiUVEhpa//KZ+ZtuzP
HpAPhb5OQ8GjUADNxYiG0x3Ztu6UuD17GCSwVr0xpPF81kyBTiDKoV0XFtQhZtu0
/wYTXHHLZ3iTGGruZ75bsGru2p1IEPrWJQQMiPSVYB2hr9WvCYhjYwGhQBabAlpF
p/hzh9kTAHOYcREJp4iXXAjjavYnnmiJzHK8fN0NjyAR4PLwrebH+UBLJv9zsBR8
me6E47KbLeGzEcNaJui7IhxNuUoMIbe6tyDv/cQeVBGGJaVt+g11m6X6NTHJ7mDP
z99vRCefNk7mHkCZO2/DRYVNn+hYBfE73QagGxK+nN0rBIWW6LHjQox67RkD0eb/
mZPwKTE1Uua/StqyOVzOBhChJhksI7c4r6mRH4SicCXJwtzpGNymUsb99IHY0MGf
+zHQnWYfTwQNTsKlue+UjbKXTzXdBh6sj2pRDfQ2Tyujw+u+9Z6Ab5NUURjTq2Pn
Na4yk32Z2jDhpIJe7PHLaMAg+HkxJk4TG5YRS1GXMHXQDC0IWkELW/eky+YOxZih
dfiv/3+AHJoyMBOzbrzU6fzFel83P1Vr1GF9qp9+lV56z4uvZ5ESZ9+x/QNGTzoU
I4mubEINyDnVh4/nt3U3E8cVDpb0VA55gV1AebWLLt1q069a4pNOVIraZ9fz6ZJ+
kZZMFw0frAS+JInCA9hLJoNK5/UF4QopxabNFgPPCo5YB6dGpu0Xj8q5Pb2c1c6Q
Ja81z57fjmm5nwz4DuNgnGHVweJnh7mT96W3H1Wv9sCcBO7jL581yrPjRIaIzL7l
eBlQrxwe6Ben9LadVu1l4WOGHAZ+frPSVQrItJnJNGZhncbugOWG94VBhepvBiSU
2TsBroe6DKdhZj6T2tS28RHNMnq+IFpqnCNcHhOtzRFaYrU/bDzaVpwJekF9N5sP
So5JbYas7A4tPQbu8qkwKu7ur/94hrcmFUGERxvY3R3ep9DQYPXGTHNUK0V+hwcT
HnunBjjbtGWFKjQZEADmon4CfVJ2cqE9FBeZEWv9YqtqQOCt6BevQJv+P9nbfItj
VIK4CNuaAbhcRnQWfxKpaD0lihIPopGZvQLJxNkBrjXTt55CXjS7MLwhF0BYF0la
U0OwVkEVGwlaw9dNlTVx8G5VIBCpOG73Gw7N8HsvguYSSoDNtc7MyJ5o3Z8azb66
U489qYucSbbN23cT2bUUMShVow/GecRdx7doV0AUfnJNa2dyguFs/da7bmAyO+Zg
F9mdsacHRPJDN8igkg+9yVVKfOZ9XAGx7uLF0QPdLS7ONT+lDqWKXHgfMjClYh3y
qNLx9WAs29A/pRbJHQ4ufM95n0yzVu6eafsL4hIYehYk+gffA71FiSrM17T3zMzw
JnpESoxaQyC+smamdA9thbVj58GVVqks0wgUxMUXXDfLJ/LC3v3oUjSR+/bIKM8Q
gKg4Y6xmP1V2da01+z4/s0phE8XqIQYKDWigvQROpbaUYX4oE9LAI5N7/9qUpDTQ
0YA2LR7DFhXHwTWsu47y8kpYlZpFFTcB6JyFHavxHpx2hPFYBeUc4GXmEqx9RCmJ
tgxcdqWtpWNhrDpLxGVy5SSzw2Co21iMbj9zjlpYxyq2fLZtXHjnJaaspYpRTkyx
esVWERnvBDiPPT6D72qVWpYGA93635yv8BzaUqO3R57h2meQHI1iFuP/D/H2Hgcj
MXkaGYkb0XQtRL3XygKxHii2jYGBv8Pu4CBhxNIaB9YEiCSBq8xtcDBWkB+7gyye
wS8o64jb/GZBQoROdvWWbUz732A7xvzd0fdZmjBkZetsyY03/TIWT8YROk7YyOJb
tdN+OckHLykJBaU/gaa6V+XIXs8KdIs0rRk+95pUATI5gUuLROl87zJEFTONVsh5
rgpLqfmSq4xeFtZlpq+OlZg7r+VdeWH5FwOUYC2VsnvQtolJBpMngiMhI/936Yhi
QiNQ3/hR9DVEM4VMlhow2dH4SN7waFcVKU2ykqSfjAnndfcp4TkxLPvkaLxOJck7
LbrRagcmmBOfbTf1LoROqVrsq2GKJ7XJfKs7MT3dFzI04llqCOx2ZUHDIkiD/TYl
KDgyvPid1+UEQhN1Pk4dSOUUWZE/Frjs//tWKByX7moWjfvif44DzJN6UZWaJGQ2
IexaX+ZtxiKC5qS3w6u9A6EmkedwlGfd9IBeY/f2gkVOalPwMCMnDyK0ngoO1d7H
t8zwsNG0BSCNgITL1V3ob0c5yF0QhDtsK3s+YyUbkT8LneTzsEijcqczqklvhKW5
/y5sEtovogHLEPtXLPROLu4aFGkEq+1ZPqtqlBMHQIjMGo5ldH+/YtUBs1Nx9xMX
J8rxWdKueGMEfEkSVgJ98yCAHM2RKeCo2qPLSPxcylvOaduHWjclDhdJBPYwHoB7
a7x6mmona9bff6ZW8rCFWJjc3xBcMBlfbHrRazI1l5S9ejWjLNL16UZl3o+rvU5U
/bDqi70/V+hHaslA+LW3yajB/WPZXBg8rjk9theDzywxSgTT7qk4L6LkN8OsMMaE
I/IEzKTM65r+mtziZneHOlYdzaM3wG7Cxet7lWHuE0vtlpeoaBr6yB8XuhTQArI1
WZ5qMidkHmPHo90ST1k7CIfly+nPqiZkSft2iW/DylMpCQeVZgLuQ4T1QJuZCxAV
kBC8pUYSu+dpcO354JDif7wdC9S3hCTB5q5qBxJkjZw5C+b6M+DTYZh/IcFJQ907
uW7uBHlR9zHgEIx7Z8srOEoGBMxiVfOmcsBYosAyya1Hckm/shLWqZUuRtj/t6Jr
lDJPTtAXJa+sDPs5jDmB4IoKS0Zlx3pdyNodAbrZAku08qkZ+scAp3j+9JMuYJxZ
AD7PKMPJtPjSYrErGXWdPI3XA+MI48TxQlNdb5Zs7D/UZMcWbUXZg/VZNI4fy8te
fTm72EeWy0WlWW8or3fyMAc7OvAlaIN23ULdbCRc+fH3+BXxaensk29/QQbVUcDA
7nKtPcOzgIFaJcv6cI4KRj3TG12Oe3zZWmTBSAbhO8ouzgtRlPe8s0PxQ+6kYwvq
8ecnxKRynR05U85frwr3uFS2baOwYMPbsFCYh7GPmCQn5Usk8eotKJ10qXiXufvd
kNzPe6DSVo1VBJXMpNjT3UuQsNPDA3jqOOGnnIRtP3+qNQx0Epkq8ndDR4aDBQyo
Q2ubA1JhQ0O3wxHMfBa2ripQDxWD8/8GeeobdEZjFmafl7adJ/hn6o6toApcnHLZ
8mgLa/k7Yc1MIdMY9SElyknZzCN60vYXGtTSLxAeup7x7/MXv92lglZYkbRfV8O0
oTZvHGKFFutjmi5rletjagHhNfsKdWUVNce3u2KjVHKGmUZS6tTNpeKbFUgb0rLV
NGfDVn40fluKJbIg3PobTmaI2o0kq4i1ZKt51pACQLN7kWLlD+0mrebdll3vHS7q
wHnlsPz7b3/b9qlLNwvoaq3vzrYg1If8U6qOHuYRcyiwB9uRuH6p/D2G/LhfP+Rc
aZOBrKTL42ex1VMrgePXs3xKjup4xuM+iIOvQrV1sZSc0uOF196SC5DjkWJwthyI
frTxfVGtWwfde2ddfVZ4MWYXKS2lQdr9PNloRS3BbZr7QMjxIFf25+YMkXk8J91f
kiwbg21M69qb9c8nQiqzUlm24WYVh/qThz7N2AYyYhXAlPqfXMMkTDrS8MWT3ePc
JmwUh010iuU5D882QZk8JOfBuFuCxDHLcFZUlrOcyDnGyb8FecvryvmVXuSu1U+R
6xMh0z59Pgh+q7HDm81lkTUm/RV87RzCvQd61L33NRGzd20ErAGwhKmTlF9C6gDy
YoqdcMDFmQ7/YN7j/HStoRtB17WvDzJkF/DCQhiiPqnVCnvJxrJx5VmyomvGw/2K
gxNLNM80cbRGuUv7RHFpXldkjQyI5mayHm2Jnk16BsOosgIQJlmen1WL3d2Q5TWi
u83ytL1mR4r82Qpt12z2aC3KXplKkpx63Bp1x0WwnsY00zjsJmY6r9pdiJM2Y7G+
L54gM/qlsBlZcDnLCG47uBU6dIMFry7uW/TTdYe9bVRzEEnTpWlsHew+qfu3Cb8/
oObrJVwr1RyQaRgVhtZo9CDhXRP9v9I63PXUvILlW598sYsdSPwyNyHBISngZGmg
cqNbYFZQ7bG6NxbF2i3GaY6R88cm0U5R9emYStkO1Buxnnikyoo5hBpNydRx7i6R
5xa4W1oi2h0zLkMT+mHU2TMKQIYQFFCos3bIiF0fY1uPcYt3O5VJZJgOApkRVYgU
pOEHgw/XpzsHh+6j9CC1CyULk5i/kzDmG9pDtH+dZ8pqXlE/FPG5Cte0F6yTXmuO
XHGZvW/HVDZ+XD2kUoB14quqPYRpoD9ii3Wqjh4iATRtmyPJcJhLr2czUFqIDzws
ASr3Kc81RlbcnbYaQDEwmEZ4j54lVjbqPwjteVbGZlDMywNIa2tGLjgfFAZB8NbP
SLeGi0OZrYZ0lb+WFitOViJMmPsQ6ComGy7fQdJMbaK+LuAtAwKReFIalyeqdtyH
f786ACr6+uXxaHY++XR+bsW+Je173ECoz3U5l4TtPV0+pu7oOZiqEijgYX5FRTd7
9T733FIiqOJ/asC30OBh4diw4U81i39jwaqUy185lbWJsZ4wgDLErdVsCeG1mwTG
7HXkQ6XbaZfPrYV8rhzDaruiZc/4OHyVR3C3G1As3a1kmxb1EggKVpPpLlGciRjN
A75YrToeHRsrarBgP4Uh+VZk5QqNMHf4c/6s2q5LfNgH7Epob3WlbCERzsnuJAAy
T+jjMphVm9GpUQErzbu/5/SE6c8w9acqWfSNOA02H3dTxKH6UkCd741c04E1ynUB
lH2xyJW7m0txX4wxlEmOJQP047IJNF0tw6Yt1w78JMzq4/Iycjv1j3sOh8w0Hk5f
b09yr+x44z2c/23lCbQ3Il5SknseLCpf0E87aHnCNbawQgK4cNNV5BbXtKm1mzkx
MbC7uzv9HHdlwcSfefLiZ7K+q0gzFaiUoBAyjIF+GgX4gewQ16iPfU9OfqR5fikF
e9FjdTpbL9O+xmiLmQcN+RC2IMo/8j2p18s5VnA+rTmsax8v4UORWaEMD1KS3Yh0
nbXwZQJhxrosVCwVJfE4it/WUWdsYiyEmzSw8Bkv/cuuw5kYJAJHw50gsEwmB3Ca
tajFIuhck6i9zVzwOUYQFtryJEaqguVk8onZpj6FrDk9WiZy7RQR+XcZZTXYIZZW
T2HoxgRkDBfciDCorq7XBsZYumwasiqOeUo7KujMeJy9nV9eMUK4bNu+ZVjP5CFp
AWEw+S8yZpLFJ3vqxsuttnqItrecOXfFupJpsPYUxOOEaQQQHsojMi0/rsnH60Z0
D2o3muO60PFkI7jrnhtbYiQlWi3efFNgZmdMrQJQKu5IHjxCpdjzMtKm9k4RlsqP
bNQjOCG4uCOqTx9b++vchHJq+adaTVnZGogHfleCE5jkRCo2QZ+DQAAbKfokd7h1
eiRH+PzVqyjEP2+41d++muIeiphmZ+3TB426j9GCory+d8DDYFgnzIeBmf4TDm6w
hX9X+AoUg5+zXGb6NqTQ0ryAtw8kNzbwkSfd/G5k0ql3IVjO6gL50JgitJXNpfkm
r9H+QhQ8tt09ACBd5Cl61etIBsoOl6GF5UcPSitoYHEU/+0Zhk6WGNI3Ts5Bh3Az
IrHcwo9AOlvs0x/IIAZWFe9YbWEXTbn1Tku/6o408TKB2PMPlEJlyz+ona270zJO
jk4LunccnLqPxY2mttSpLSulFuAYfsrHthpns9x9nAGmW5rV0S2ks7l0h75q7amV
XCyDDRNTpHoZRdf+e97xCuAsSaZF6e1M1Z6CAgI+MHH5gdFSrKaWpjfWCRBJ7uR1
/YjymJC1DjJ5fIVqXcartGAmgQ2MS67AKOKBtujuZIfNlOPVWu3/NNxd8IsxJUSm
N/HFSG+tmHcCC9KutrCe2Ion5zogITGBbA0BSIwm2tSsNFdphbf2DgUlYmDhw60y
bMU3OSrHSdTjR5Zh+roraA1EK4LJ+xHN98/YkBOroj5k7T7tQY83ZE6LNkWpflRz
gUv3aNfBvyZIAZxQYiivo5cbrQ2AhP680oJ1NiGepChi6boPQw0MgQLJ42C5Brzi
AqcDdSvC6jwfgGGItwUjo9CNeVwIjniQCH3j/fmHzzhMnmpALA4/HN5zQiWW7KXA
peGfP2w2mUVSHNDS71JyzInpyq0upvfqOz2RN7lvZDP4ckuOSvgTI1ntUQUWtJTY
ZVvs0hl2RAF7nRlO6OxaXg1g1hzBb02dordkK9A5dmLdZvtgsa+ZCl6isQoppW0u
JPsbeUE86ciRuPK1hDV7WdqDIaRqMbqZc9UDhLxwleGdIy/3RNbXCF7xw4ZJ6vRF
yHaloARW+6E3cgS9NHq4wNY39xakKQN8rgk//LzK2P8+DPPYeUDlxYoDd+lgTMl+
7gPTS1uL3QSM6BdPtEcu7oIQZEf9l1YiapdRuLZlPh0WCB6Pxvxu1+I2gIVWBKaJ
zhYnM4IIms0dke3G2MaGvk6ak63N9P0puOZRhShHQsydTXUK/+ZJ/XtbUBwEom3W
TXEopkxMlwpvW+MWtqD9SwImpgRkUS4t2oFW1MnUTvDDTZYqFvIFlV1V55Zze/BM
V67FHqoH8hMeDfMA2yFalBHo/J+oGx1WulEb/biSwEGEBhkTO2isDTVP09jYQuPy
NYPiCxf4MUG98/cEwwg4nAVf5ie9bbwoYj8JCYZdkEIAXUlz+PGXLjfhBnGcqU05
pmmcqZnFkIYBxFcBV7L01UejFDgmuXItiPGQcvk+LZLHahwmcyHZKPXny0OD5kLG
fqfTcnmBrCixENaP1gSLzFj0la0+a9Sjz5PB1gaUiAq7ABuOQFn64YY7S8Ve1opz
h2iMAHEAHJEYMFQhkvSS0swL5CRswz3sGT4iW35e3H8VF7fqeQOCZqbLbIdAmD09
yNWB3TAfHqzRljUqxVP/cBONFsFBzhu0paBG+3MOBurj+xXF4dxQQXwXMJmg1bha
UQbg63S/AtjytCM5eacyt4fBRTmkgXqm+7qjZkJcEWGKTNNpvobcJBJ9XHxJmOxD
VdEdYWgl/SM3gFagf42Ug59PYfvf5r5tPibSSnE/kWLbdyA/4Rdb5C2psMQ4xJkV
F6Jbdu19wGYT8RfciN6qAVxBNk4eb9KFQwrhctiStFdksk0DAyR519Io/RsJPm+/
Ey27ZudRJ/xJmJNpMPAyN7HE988k6sTmijm0vJY5mmKjVwznLUlmQVpPyqHuckf8
lW238XvaOOZtF413YiqpCWf/Mt3UBrTWVfuRyIrKjxC5wXNFCbYomH4GaPK6Wmce
vAc5xPLJosFRPdHbisvD00YvI4uOUbXAqSfloTEZG+UmE69hSd2IXKzhPJpQJi3p
XM1tq3e0PnH/l2nMqWkSze9qW6KHwlLP8Zas4JObz8Dk1iqDhLDeXNraROBb3jy2
I3fwR27jfyOvw1s2AW4iTET5km78nGT98LvcLKJ1nEW00HibDnzJyLAbEB+wYQdh
+oezMC6bJzv4xE5xxs5QebVRUDenOISroqitAKnKBF0HVLYavmH9Ix8TUZx3a4ZM
nb1k/kq5/54vEA6TuJ2aK+Pm6eO9fO4mh/Hbln0PGO+nR5V03TNLetTXGHtR2Q1H
Yp1Rduc04KEMSna8hm/+91+bH6y6AQY6RMngnnKyqYU0EaZjIRUJhS/VqyymGHWU
bME6TfkC9AYO4duo608nALswylqtJiBouOZSm4bLcRSv18wizjRxxobcgmJ+ct6U
vJ2RlOjVDIB+KX7j/9kk6E6k+EsnH54bqzneGdAwCsIrqC2y06LWzlVEuz2Vv3tD
ydGHEK9r7M8rSFQl5j8Xah0genMd6GnEbkse+sy3QXvBsahjkeXSxTgNAnti4h2i
SMi3BZviVcSMhIqxTqKRA191Fkbn46156wSylhtjJrbw+0icJS5vkGtRHy4bIS07
nVYC67WhPbaCJJBREY0icMHX4vRbiT35V+j0wrTXec3WsF1AunwgX/gg4uIsZnTt
/IYBKfwecdOP+Zl64BTpVhSDGbPj7m1+OTYko3jN3Dkv2XbH7K4e8voDR8Y1qcV9
PTa5WvoTbztfizO2xh8QTs5rHfGnI4/yCt2be2inVYj6excpsgJuq/T4Q+XVx7Xx
Ew2sWwRkHX6KyloBDwd5OCcm+7e16TGUa6zXMi77o4M95oFH/SmKjX3GMapmoFo4
q6T9vKp0YsKkadcgSpKgq5ZCi/3Zu9455wIO9Wkq/0PZvI4JArV9PEzjFIq1Xno5
cJZAy4dR1i8Upb4uwLIZerfLdtgxVlqHCs+RPKB3PvwY9OyuWSBxni2mB6iBSN0u
uKXMgl3hp1g2ocyPrJ8eWzFefgXModvVP8n0sX/LAJdSF55qL4ZHhT7jorlsMAuV
jyDoW1rW6YuWdyUn1bbGTMePXccfIbSFaOlrckNLQ7QbpYf7IMZ6sQcWx1MTtDqy
rzsMqQ8w1PfAfDJ4aZPCuDTnurrKVomOXtTXuIURTN0Fu43yFCHR8yJFlfnmlsz2
NM0mr20zXRfAp1Hy9ef8Y+xFrx35/MoyfrmENCpVQ7+zbO6atOLWVcKTDxeCWPMq
ErunXcSz9a7v54IqbCnX7Agb6BruzJIa4wc9Qh+mqzIS8AYT+YO0397aikOL83Ql
BLVB6o97cibptrrsO7Nur9L5YREHIrDzQWlqL9bEiuSqQ4SaCeNb62Wt3CkYUzXV
Mn6OR2KtrAUqdiIfzWhAqu30qflGVElEUspiFW1PM7o8FHeKPWeNWAYcsrBRmj3g
MVIeCIZGp9WULbTiRTyUYs+RmdOePrT4bserKHIE2/2Rh1+//qc11zexx/gwCjh/
Srra62sOWqI9EKhSrw5OE7BuH5HP1PE2qarZtO6y885IHJ9ekcLkDyOgw1MgoKsU
be518m1n0whi45qoVkM5o1nM/0BevHimHQKNToa2djEn+tBASD2Qo671vcBfhfKN
j0jcajC5dDfZRAN7IU+KnGhLKgcxPXo4JoxWurLpn86cbylLl2IIEy4iNguU9aLr
df7K1VlNTuI79OhLQD5lpYgSEbEOoE4O/ipPiZMLb00BOeXR/THvl2Gzh2gJjxJi
q5fZO+6o1TuXYBtb/y12xWw1O8eEYEgtUDNGRslfuR6Wo/SD1oh651LFsikvCUhj
GJmf06suQKsIeD9Y9/wd5az7xkf5aUckbbVNYo5YyLIfIXKn9P6k/BgVYDm2C+3L
kdHCaqFxWv7NpO8pU/9hFsb1QE4DFZB/eze1nzTNbR7I/o3ahVjqZJhukmIF2LGZ
scYurvOQ2RhqzBLALsHgt/AWy4moA1fbqZbzwT4gGyHYhbt7j9W8yeFSdUpqUplc
uiKdrJlyJRHg04b1iY+CU1czA2gZCjHzfmWgDIsQannVy+KWwWOw4G2AeoO5ke4o
3Bfna//6VckjIs9VoEPl5LPmJeSn4/49j1DbUrDJzoXfOUdOQHU+/TCDsJZDUH8j
3FdRPZlmrdd+/5vqxrwtZxw863eOh/PffjJmo6SpMzdygGHQlmc+e1QUP2n7W9r6
GAVpcI1o2pvH8/jauhLyaJ9GynCY/LtZRRZns+H0XOLoC9CGiA6VrpuCkqHH/UQn
fEqOK50zqe20vKEHazcMDOuRx8ERgHoWGyrYyW83o3J2HQvShlAXpmg8VCY4Giwx
28OPnk/Z/E/5Scjks5ocXNHHr82Gqkkj13m01PDrXo5CEA+G6O8ZpxU9vz3dypWM
0UJVvffDq3zGrs9Aqy6YjqG717HhLzdVJ5jhqeVDNYvcZGtZbdlfXzCV6WQhgGIk
05DWh8vP2S71mOZj8D6vxTP+kwW39xTjZolipRsOk5LjsTiPdQBjpJynVA4B5fcg
CdV1A9zGZeutzb9KPOLLWuCtBDGMN1E20TmqQvm1MjavqC33J9rzrVS9WaO8AXPG
0i8cuOlreyCsI6wEFARudf6SUjoLLS6bAF9dizQaudZpxzxMJIRgq7/tXgdeQ8jI
tTI+oDR0KG4mQqEBUSfxy1VyVi/CzFK8UkTmWh21YZXoUaapoz/vQFED37ZWJXLX
k+x3ioN9FGdbekGrde5+7US0xHRxke8YB0voaBB4QHPjdcUPUhPWyub5fzScrM1x
4aLRQ2UY8qDrJXSrA6LnZouF93KIFLrKA0nxmFIbQSwLcTaZEVhGpWlx8St2L5BQ
OR0uUVPljUDtiXjdwN2PdKYs7WBgYrYPFeEiaoVph9KhcrrWMdrREIIWE/aFcpPQ
P83EBJJOCkuWNn2LF8aXsn8e3kSjbRKVuiZZ+81dLoGKFcuQ82e7seEcxv7t2vx0
RI9liSjVVes4aRE7LkJFNXUCExBb1he+E6p73ROGD96/kRMJ/iGDYPZrI/hi74FO
VfspdaCqdLeHvSSU7lBHAVH/OG8eF9sj/XAAdWH70zt1/ekfehX+Kxzdl3NmZMWJ
PtDPF4lXlL5G1DKxYibW+GMfXazyfm1zIeU1cNNpMTF8ebHi52XHVSyNZ1DTlpOY
q6hnowAFZXbVhRe5WL+IQAkvGa/qSwWuCcB6E9k8OfLXq/j8Bvo2GPyPvNar1uHI
/kGhZMeJF8AIcbuc6kr4hpD0z7OYvZOIVAYP849MF4TPLqMKrvhhMZnVCcmGkSl1
dzbZlPAvEfEWZem2xhtcMfD68QbertByPAHhhELnImJsJSgHK7Wjoja3ILHWI2SV
HA6u/dZ+ThikujsUpnpr658Q1r3i92aJTNYFX1Do40EZ1E6GrxqKLRb8DFSFAhy5
gkwwdJgNMQ1RJEX94oZHT5Ozh0fwCsxUUzV/YC0NXumF22VnQFxyUCMp3BTbnPnN
xN+2GOVGYjalowK4rokIWhAO44HXNRr7XwLEkjuDSKiFD2LKpRRp6UL+LHmLfbOO
j4nV86DKO1V4KNPtFmjs8crFAuHbueDHYx7S3p98vDupbwrfgauAeDQzyhRlGE69
J5KLLoJbOMm3hdc8buKi7L86FbF41XE4sgzxQ6zkjpP+OoaujY9eea5Nyk1G9RGq
DjXAHYaMU9H0s9zE1lWnUtlyE3FSRcRGARw9DqDoLkC8OmXGXyak7S3F1tlYQ1EB
GI9Bs+gvU22DI9Bj49rWIQYWrYbOTobRmzzgPXbd5wBm92x/mHLi7GS3x2+k01ff
y+ti4HHpeW58JS63iS3+u+IWyjnTjr9E/rqGNOyBxzONuvE4B8tgtDX2fUheybWx
FUOReaZK91o95oyi0Xdl9ZGfCcKlaSGt9q+Q15B+64amYVeIWsVLgOyj93NjBxJn
hFqMkA2lvj+XI8Nd1b7GdhFYbNuLEwOOTGKzHh8UgI+KJwfoPZH9lR/HabrtbrWu
37bwUW9ccyAeTwiuQv/q6E62GKvSBlrfF4VKM4L11QdwbqYYW10s0ofioYM5kEm5
xNLeLTHwGmaoVEEKyWigTui2pkUPcZxa7OiA+Jkdr+ya1rzSWCV612bdpzq+zYH4
ed0+LjfrVGe+kE2coNv4T4ppKdwljA8UEOjlQQNH5qNGzbecIAcafvZDeWDhwRyC
2Bl0OXT9/wcDoVHJSTFnqn9UWSh1WDjq9i+jB6MQ59DoHWfJBJ99B7a4g5FePouD
k4uWopp0+aqKxQlYRRwg4Z+KtWulBcx0qnHAzlS96+hz2piH9fYa6YYt8s4Iqpaz
pOvGX730bzb0ZPYdS9o01ZV82IGpajgoFQcjSFjlgeoT6SqlLf3bWKY96UpUnPiu
FdFRx2Z8WRtntfsV62MgDESLG6vsB/TY63sFJfwsjymG7eF17Ufzm6dUvrkT2aZP
1eEc824gjVQWvrYdYmlB2M1zdvhSJcn/gg4Zp11vUXOFz0i+W7oENEHcvr+xg/U2
7L4jVGMAjrUtYxjwrf0sRC7AmVVpn2uVWGbZvTpoEoRUVk61bHarBebqB/qRHUWJ
3HmPrHWj1eUudXWZlXMrGx4Uku4XzL3120l7f6zw8l1G5hPcKK5Sq2z1nMyHcuYv
NIWOA26TKQu/BUtAUQ1qeniimyNZtmFRyqofS1plQSV8H/YRQo9GDZ7/4xTh5JXB
x5Na4slG7xN+muSigkflEV/ekB/hSrJsf2D2AIqeCoTv107iM54EC3Ffx2zQ/0ep
CerQM0fgiaDtNUC7Tc2rtv0qkzMC1DZw53t9Bq+FmUebzauNGa/FDMhkRR7cGKsV
IHIQfkGl8b2xCD1yoJvdopbtVL9bXJmAj7S3ut8TT7+GZ+nyIV7ALhhQtQCy3Gtu
KqMlplUForof7nONAoINIYipeS/MwQMXCGDM7lCgFkZVhr4T7fuQ2nj0GJLSZ0z7
rEF8ubRccCsqi6xuAYnG+tlTnL6fSkAMaSHgyJYKBboWMAQLIYW0gTYrTZskVRRT
8bCrSkrM2arFMX5+JO4JX4oWPIiEug75IehxONlmTvGKvFabPifgyCE6x0FdPI2P
Pbe+ivriV2SwpGSCY1L4BowM5dYtU3enF9NmRKkRO4lriVAUuI9Dz5gcDUvBDJhI
TUe4wmI1RT79a35i54vfIOrKM5lm6Zo79p7LR5+tGxYWaYmLci7LZyqRsg9RVtDx
5Mi3MjE5awBmzxn3KLIgRhX27C4wsn+yLqSFsML6r/1I0CImSco3kJLCzJBDYY3E
vQSe+YE4oYiXRuXjuFS6i7mHpa6EgJQLtJaYWhKHqFAfvGjaukCH8beVsp45qWb/
Vwz4ueaQzOYkFYwRHGE9dAwOQY4J+RtsxiOM4nwZLpkDRB/KVSNWuWDlUFRnO3Fc
Qodx2BDO3jgh6brUIOVHn1fI2r3NP39OglPi/YJ4afh0pBhaNOhkkennv6qW0Hbj
NzNLv2Z8o5tZ8/xV7zAO23i3UabGYosLDbzsT9Zoiaib/x2FPRpd5Ko6OXGz6V83
EQ0M+CcbpqZkzZdg61uxZRehvtObBR5GPxwHrExflsLzSfSVEelRhFmvQFm4xpAg
6A+Xt7J1NY1Hab+AlcXiqwc2wPLzkgdolsYsoMOcHOhhsffYJ2k5Ash80RAF/mr6
eXqIjRp2srNc67P1e6hlPSWbpFO1RXIq5+nyJ8tU9n/Xkq9Kl7MR1mtkpsTW5uG/
nyosWnaEWKO+w0sweFTI17GwsZrpZNya1DTLIOm1shBR9X8R0zTUcCmYs2q69y04
6pDvyGeBOuxyIu75kDd7F5k7l44Rb4D0jIuAofv6rwZs8xH1Ld8JlOtMyJ47sWvK
nHtiIagv7pHysLGeXU8OleFfbTFI8ysZog3n5daj5SFQBcyEUL24QLcHd+D+P/cf
/borBIzi2g2wll7r0aWv0wqLzTmGw5oR/iR8eUne+vnjjrIP47qg5ycTWf214wxK
YrHpqLZSSAlDFbaj37xfbqhXnzQIwKFV7aC9SvUu+UbOhW1EunP46W62gGX+jFb4
5byd35lTZ4cUl1u7nIiUT4ijLMS38w17/3V5Kb41lcL/Ih8s19tOYpYE6QcF8/AM
arl7i4Nmjb+s9vVp1yUQOy0IXkBK8MORwGDo2l0J4nODAxPNtdywW0VuC9lO8tro
XeESDngE85vEuKbWinjmU+K+qEcvPDg+FpAJCttD5ZgiY51Zu+LwFMGd9ePhOkPW
2tvrS9meauAWqlIfK0Cw3nKGdVK6DliiV/qL+uzYYBGxkdUoBOiczmrdK8Z7FtO8
hcZKsT3JpMysbKdwDqH2x9uP5NyUUBX44N0Wckjh1hdjEuATvmXpsOEP46FjjZGh
rCmPoUEjtFJt/4DI26t6SDiSYL3y9/MzyptwIeycOCvaZ0S8aXD72FO5es8IpF8a
aC+RuDWhSQ66h4861Wi+jGFiU7PPabAQQ0QTthZhhGlsV6QZc1nEToVqdQ8sg6h+
At64XWUtWK3ZW8o6RWword0zslMDTYcB4Bb7cyfTY2NgzIDJYyu8eQzignW1T/C4
ZMMy0LBDvUObBHAzAjTfDkI0Zy7TSB8lHHHqrZ0eO3UTS7qS1mcuto4gIT/qG4BK
DnDlyR+4OMEn4gAIbb5v6tfichpL+6uBLCp9/nGznGCZILd1Hq8zUGcwplzWtByG
dkvYyoPD6d3it2lJKGSRJ+8+KfiXo/VGIwB1JkD/p4DQJY4luPdrqNNX5GvfKFSQ
t585ZPcdWhatmS/MuUULvdoJSoztMnjmApHfxsOW71RicT148zPQgBxX5VMOQhH4
bMGwTB7HPnxg00evFTZMLIEEBFLkBY9+Yqjn3MGcNUaskchVgpl0nNRNCZGPRC8c
kMJbxzB6w8DgPdAlRZztHLSG0R/0rrSMRQFCUt+QRUyXkkX4iAY1I8MS46fY0Uk3
IyYMnSpv95J0lUEhqgCizsimO2NI4pddRAuNqJnfOoWh71x84whmqt9DImFEFkrv
qEM+jMWoVXjNXE0hCTBi8ZNql7hnDNSva31bwpma0oM99MSvwdMQNpJ7tUVdAcGD
U9dZlJB9bFtWDucxPB0w/mtxkA7+d25Jpe60149dWpL3WHIHjuGiqTI5bhBG69rP
hRkf9EmjsbDJNM3B0kXne4I0rAvvjaaTEUHyQhsuRhKP4iPdl3MVdyQXOiE7KbFG
dPnYGI+zqOn5PPBq4iEhvi+XWpD4qgLnkjXsU+1IUquojbEe5Sl3BvMi628RAkvS
Ast/xm0OHyMnn236Qgl2aCX6JSSXcpTgO1yFQGNEsYHJL7aqPt8vSq37bPlFf/k2
4PHN3tifNnaSa3CViedZChL8plekMjwx3hDxO58PYdk2v3CYXViLUot5jFlM1F32
TP2VVpmR0iXCnVaKZ/y78tHYkqzY5mgAxu29X7tfZ2IvH73F6gkv/yJBLbWrCxu+
24S0MQU9t/wFCi7P9JfL+HNzILnY00N5i3w7i262jOjh55N+BJjt9WszLDyugSIs
7qk8YzVz4nygsjUR/c9QEacZXkmw2eACii+OdqRduRS7tFb3n0H9kSvh3QOYJ43U
4wQate0g68oif4/JpbUMDHrQxwIHSgvO2pOGgKnPpF22UuBClxCb3kQgJNBCRZEh
H3/MTMqXunyVvHilwrLM0g88AhVv3T1VdWv9YfDFgc1XL8cjSlEbjpXUEQ5PmsZo
V9atkWIAQIBA3Ve+4fAvkdIp8W7WJl6WhFjOZZ+ET+90ccO8goahNx/DfRK61He9
2/Y2JO13Qi3m9cVZHaGqYzfC0PYiUls5WviFyt+dN74cQwYAy+zlvglroAwqaeQc
zaNT+2d/GkjXaJ8q1ibkI5TokBGMLcgu9I2zKDkkUNr2GmB/Bhj5KlGu3S2DworZ
NYpqM8cMmS1VCvlhFEQkFDAfIi5Bi8/FnBL/Ci1u42uoy7T/LYFdrxQ22hgNHwHX
FaN2Hjv+qB4rsQNSaqS/oJbcNwgni5NFT0IHXaV5bx8ldmmGkBfzyT/5qutKfOcn
YbRXomt96/35X5FyOEreGIxh2LnwW/ENlv+uTU/l0xIJ/Ln+7nv38ayRrRP+nADN
oKQehsbKTVSBsQInAWvvCgjZD5/Jh+Dqo8sIV1SIFVmA3UHtqDbwkzTxeZyJtM3P
OGlwpuhd4CqmfDbffC5DUc5pOFf5imzDfmAqjJVjBBPHupOGiDOQ2RQ5jlNZoXfJ
SL8d09VlfkWE6YYTTn3723y6j1RU9Sxpfz4JXjdCNDgrylEa3yhHtAF2m+nh5RBw
bd6nlUFxdWSkiB9AUaCZm+ZgFaTPIqpgwuXyRAZEWNHt+JcmQLz2arUt/W3qXaS2
7i0hyE6CZgZU7h3GoO0MaTVlqBBdRT2W8InMRVbeALyykPg1xN/7+FwPI7WX1VpP
0nCOQb904s4FEl4C2paquETANIINenZ+W2vav6fzEXacSb8U6Bw57ZAurTE8f74B
bOMm+jc5RJEdPP6CTvCqqJ4uCm5EITYzSedYIgUXqKsbBlN8w4JgotpgsM8Aa84o
Il80JHMc94wNrbee6//2rywQrTKpWitTh9K87R2NswUtMX9ePkBwgjXwklEoXIwL
NFnIPvK2iFgCOO+IYc0IESB/m75E7CTGkRAXd4Q1YrswrE7R/YkvCZwHqmt/YSLM
i/DshwLMg6ujzko2PhB+VwxSFM1q7KbCeX/Zm/eeNo54i/XKjGMFFVAnUdLJ7v5o
uzhmwP8fHyExP21G0d1tClO3DRN7TxAV+SwfBs0KiCtJGIDmuv1w3TQ8zLS1Qbgt
tq97vWocoiexetjXQSejjLHXLLiJYrI0HC8Qepn4dTH1RnhC8fe8MJAUjmmz3C+L
QbJHwl5rb5EmfYpDTqAQO+iSltShrUUiYRZMSCXJW+8eHXiT5eP6EqtAtq94gvAN
26aIY3pdd7CDn4ZHIURVSFw9Pt1J+i2h77nE1P+slcshHCx98RspZcbjkBsW5Uqu
BjrRelnOOjZtZsBtlVaGu9SfokaoUIzkLY++QxlrptwYxneDj+V2f+NG9U/EjcW/
uJcV3VU9IXpRdvWNqrcsQALx5HQPIn2QkgU3IkMhvsgynr+tTxZ71N7rZkyZfW8s
5wLrkRwyZ1QohM0C8b0kG7KNFFXdYy5EH5IC4uP2u2ROmIjUgzTHCIHjOEwIlb7Y
PgIdTAm8/RwKe5e6lmlGhchYZThUNH/LpWwa2dWssBWUm+48UO9naJpjFUpRj1XH
MZx3XyeNhc1yRypEnOaW+LgY68NEnxN8WfodV8V6KduQ7dXpg0w2KbGIt3/7BvZr
6+N7fl3IkhyUKaa1Y7Z21nfuls6vuA5hO6CDbOsLixSDTaP7uo5Lv/MHnjUfj6Eu
DT0hyRoAn55L9uE1SyHkt1wvqxnAAo9x6JPW61XgDhGp9XJxEs3dNMjpc3ZpW0jF
ly4HHzaH6SWWx6c2KsDlGc+v2ST+/Os7foVEaDFAej5oGsjwnIJ1cOk8lOmELISS
WOZTkB1jmGBi9fA1z60UG8LB9xCNm0pqUpVOv9W38UeNZk/JHDwtP1l9nTLxr2OT
CERx74SlG6/5J2+Gj0hCaVeWxdyv1AszJTpvXtus1UUayRJnbfDunSv2+qb/Ah0r
7tzrsxU1PGbfa0knSX15dkkkZkF5G2k28gSM+D1CQlKvYPiBv541Q92GK80xNJs1
ICfDhPolAioyYjlpP6VLIM6HLwf8zh4e5P/a97mKbHr5f2taPD2CsewY85h3uLlC
BbiiOidBnzgKbf2fc1G8iK920zYlJFKeICB2tVwEbDYLYrNDwxrdV5JoBsH6ujBm
T84UrsJFbq+airSlyw3IMPKPdPzZKr8bLsMDi2oOxYG6MvW3/wtBEQ+Em94Pm+bN
XzsP0JEDRezQqkaPmePOE0kPGfqIGIyRxjOih0ABGzmvP4H1FORt6dGFb10TCPuO
rqr2D93m9ZH3l40j5Qc5OQSGk2h+OGDO06//gVtVLv/iSfL8Uty+Gs6Jg/c9xE41
Gau33dlhikDg7rt9+UvINHicG/LjxO/y0gO8z/XBAEfWeWpXQRCkEq15MO4pVBS+
DEn3eriAGJROlFA2pJJFQha2W/3cBBfR/N2b8C1VZdWfsYbDwqGZBgK/PmntwNxt
loNOvHC41/MFnSy5DWBeZmg8ay0JNFjIixFf1aMIWSDtsQRwbB6qz1lHDAytpILN
4Fg8PGrY6CFshuD+WFNF6fWbUxMEMnw7A8WM43bBgKKPB/1sP3GiU7bc8PwK/IU+
lHzN/TzC+TWId9RfhKTEJEAzCjuLWEscKpBwsj7fUeYkL73otxfYn6kExSYJ4ckz
MftMfKZcISFe7H6JKEpy3cuUuBkL0u9C8UhGSPeoSv77FAqROVefFLfi7jG9zL0w
YBusnCYPCZkLUCn4GGJM8G60v6j6xTz9I3tKPv4jok4/XMmhAGPCLgiZQ1rc1coe
4lS+a4fsc0s4Jz+2VEPKtQJrXlx76jDEa20PZ6kN96s7npGk3rSiGQEQkqOiSKb+
Hv/P+BSNvbgvnOI8E+fr6adTkcjcdn3F/hoeb0Tn0Ug1FDfyJOgu1rCdxYJGDjRa
Yl+RfeKeLV8uJtGzjxaxBanYB7vipopxAzz6YljUCFLcYidKG6bYI40vC00VtSDq
gpf+d+3WNq3iYQ7GTIVG1oWlvXefS97RZyLaR0TovILRTPWY+7l6ZoG/lAoptNnq
0qhOQlpKSgSGmys1oLjb6EiGPXbLa4CPYjpC0b8o6LjuYcDcZsCk8FkwaEDLqllY
n9uPoblVN6D3lO+HIBaJzVc7Aob5Mnmx7iAzHPNmHX+md+YLgnctoo97o8SLGWGX
heYR9J9KWswwu7exZ0m2ios2c+RrzxKqMHK7fkpYa3kFRKSDFdw7O1PaZOeszudQ
IK/4mqaT6qID1Wy08XzmXG+gmI/8c/8qmEX7COsI629cxJ4TyFcluSGMMCVyZQpa
9WHc3Vazwqe+Lwzq3KhJGvB2w/v2x8vEKCb5sInWfs7pnFMlGPeWPu+nq1Bl504D
VkBSYaDGx0mULUbrtEjl2tenKZttcGvyXvZACmgbbPaYAL+seEJ2R4CwqKdnl1h5
KwAuVrLJIGI9gn8MKubiiVAWWCoo5e+xfxTd69ypRwZ+/udDzhYeAEqfMwWvlTyv
rzCL8zl+fOeUBFQIJqsStu+azdJTbsceNfwAUIRrihoTfJqUYfXU6ZgBKEwWHr+i
iXfBg2zcKVsP/fNc57rVueDDqF+6OYs+1dtwbLWPmoAToh1F9tKP20xNIUV243D8
ZagXom4UfR0hgKyTuFAxVq/daAGfq+6ObBmyceVJpYIrhN7iHWgydeDl/QVn1OP9
BxdjXa8/1EEITDTIfxfHb+05cXu612kqKe9i0uMaukbtfGBMNKGJ3vYcaFEvY7xn
53VJ6EAetxb+lbnp8gyyJPac/rDvRArhwNRTrpfTAigR1yaaInZRLYFxrzmwNQzG
EAOPTiZ7el5QQYTPKpN+d1utLvjYZZJ5dKyT5dD5vqHRt0yOqJibaSHs2SCXx0OC
pRa7UFkwB8osPiudALG9lpE4d4bq4YsSapitaK/sxShzKKkWl8YiYiEdxZt7nf6H
QINozXIOHGyimoj0o66VqyLbggd3HWx6EDIm13m5ONtoifRCNWpAiSL0Ci37GAKE
LWhgcZAcGhM9PWyuGHaE9MsC9mdANTMyXri/Gru8vMGmsKw83Xevw3rN9USUCMdw
wgALIQpmuGmR+CQmF/4wufz1B961ucQepypQgStSYnSmv/CVb80idgSLnc7TY0pS
/G4IOU2wAKrYh2pjMdinll2iTCwoiNDRKk8+CsNN2oYtds8PcgBBon7iKotj0YIG
1MAvlFCvoS2oWZvQDWtKV4nEDIlScBqimDa8nETtALLKZo5zPTjnGQQaRC+8XeFP
GKVAmc7hHMj2girr58bZ1LndQR4nnxeyZvjIhVla09mzkINYFQnpBBBB42w2qIEM
5oFwdv/var2ON5mz3YXuHMActOgz5VisffUY5VJ2Jx5WEid8BL4tqwdmHwYq1QPJ
YSa98pQRFbX0GDI4Z8WuphpN9QdTejwRuxGgCROG3Rw0MAYCRsxwy/sN5MbmiRlj
5GQq0jZxFX9KlshpGnBjUkKopfL4J8aUG+kfwsrzkXiuTp4lLXffSYio8S2dPSZK
154G1Xu95SNepgZ6Ypo2KrWrah6dxAHf1b+7mYPIXvLfBfdcYVlbVsCO4IHya23n
illn9mVqHZZNEadZvNW661WLTMHDkcmU8jCd5JyEJ1G9HCWYRVY789Ccdm6sWQTd
opWs9/whuXDwHatHxIlQ5EHnGE2SJzw1/sQcS/Kk2a+5KmAM/uhT3R9F0P5N1kXJ
P2/sPZoFkp31vReqkLPxLBDaPNhO5E8V/IsipwUNaiiACKVBoLVoX134bQm4qWpR
2WYPfdipTjxHpQCc51wHiNcykLK7d8PuWKcaP6eIOptqF9EU3NlJEUSOyXxtT1TQ
Zf6hrVX6wZQtYmPZDsFCn8cA6BJoYr6OaGFUjgnyJTZEZOI8ptFN5FIP+mnELLhl
3bgiqMS4/eQ4q7nvQ1w618MWSh+Pv5EiS2LMOh8RMxw9ethNmXA4+JY3PvZk/evE
qUpaeqmDKdu6zDvVvK/H9Q6AI2I8iLaFfOoqal1Knd7s6wc7jMmoKzr9P3oumPpR
EbNFXBiq2ni/2H6tufcf3vGdAgUAtIg0cTetftU1FFL2nWD8YQWkmGzg8aoPZ6wy
h7WCcaYeQBUUxkHRdK9hQol7Dx+ey6ywxxIxvgcGeaWpG4Jhnq7PASjmfT4IE+B0
v+2Y/6oheV3mS2+uQT5mzkJDQIKXxbOgcOu+iLGLQ27eNvXJvyndjctGOzfb+9SZ
i85vKsA8juiQ4SgisR+1waDhS8E2fsbv11FXd3yfQl1j9wKln0HoUzVBg/ULm05p
Q/XdUbUEkidxGuGC71jmIVuLM45m8gW6aWPdfxhgpTF27epKtKpAF0hFgWlt3vZV
C8lxLOf57yf0HHwSClrXxWP5R9/X7udRGtuMlgOf4XT37eEKQ47IcJY7UcjZqJyZ
6VZkBGnTztPa/+MXl5WqdEzFRhqzWclPh5rj4USMp+cK16BBkNEhmM72k/DCK7Jc
QueR9DMhaFYgopQAJ9rFEo/HZbnRZp5oFA+lv8QBbutDU61YK6vuetMVRHCstGD5
3rkoDkdQ+OPOTlsosk4eVRniUS7+Gg5JAdVqfEv6U1J/tAaSQnnfj7n81awvF4JA
1Ysd//9iGUNC4Sh46z2dxqsbCimT36Rsm1JwE2374p7l1cwT7nIpQ62bGINwgv7s
cBh0LCuFdg7B0m6lOWmtA2pbxOSJKTALYwCrE/Vo/+0jJjoTXMabROzzVnwyj+BR
E1zyTCdRmrahY7tsTKJS1U30MCAkoKcV08Tfr1RN0/oqn/FsKqXv2GYiYgSMsGyN
b6hzuJ/lfPwE7osDg9Cz6Tb//rtKrnbAv7Up2GP6KH9YKjHIiJYRUuvW9qvT8WE/
RVaCI3Ig7V8yXv5nKmRlowW8m208FLrzRl7p9DwR7rhpiyqx0mTy8WTinCV9Lyu5
t8L7jZ4qNobZS5yc/mkzL4TYg2oV6FlA3DlGBT8fyUY6BW2hJ4W9tF6TCOFF1clL
UF/fZLYfOo6TywU/PJO6NHVdMd1UsEoK3KFHmFQUpMBnjWCG84Lujh/Kb/saQy5F
ZRpvByxw/5GQPR4fJ7KCaRntSEyzn2WyMLbTHLZoG54+5xfjGZ5Ux7y7Tej/G2qy
JuahSvQwX2AjflJ7BkeU+rp2MyFTNlqlhBEdEzHz4P/R5joUeFxmuCV+WbjYLFoC
Y9Uzkbjz21PkMJPdJyxrdTpg0T0+sTfaR1W1zYClohisnQ+9Dp8JVuXFTjqZD1Go
mcHedjNKHuBnFNqBxSzIjQ0H7WLvSOTXW5rJIRh9paxE4zzoGBjYmyLl9iTm1zPB
Q7hcXUu+YLri5vDBjCdtt4+JyljkeQzWaSl3fvkvyVqw6urb8HCREZv3ySHpYCvk
HteLPJctyEIzUYSNP8bqt8mpxjoR+zIv8SpbRO6iy2OHjPxiluI772KYs16fNztu
IMMk3kuMePza8Ep3WcAsg4guj80RHC/RvAf9AWt0gQul5gO9WC3TAZ3UeX4MnjXU
xAmwZGeIPl4miE0qQXg/cFwlvprvuZ0lBl0lYXOQhVE/8auKYjCbESAk+uqcgj1X
KcE/YA2QYUQ2y7rKXv0Js6CNfTuwS09XYyq2V0fLyvq/0NBqq1VqPy7M9cECQnXv
KL6rCTbBEZliGIlj5t4lqsmY5UmvWmReK7vIG8rGxQhYUPrAQCTPdXib+YtVfOEy
8GnUtC8umvirvwBP/iIxF0zf+baPdrx6ep2+IGKQqDuk92SXJAYDOKzkP1RF+BX3
82ft9DLKawNI3w5wzbxc8D+2gaTjR83yh7PGcxsfmitab2+EhgEW7CWKhnknG+Hp
DA1WrAbzlctmWboXuvPk3dOCa7OxqOCJnBOCQqZ7qposoj7k21SklHErBy6msPDe
St7PsnZ0ex/X8IT1AP1zw+mGQFk1ggpDsL+hd2LCaRxW2H0+a9RBq4nVKjWJQXof
2TyrEHlP+INcULI+eRNS3omBzyrsY10GlhofLTVxT8xK1rckXOaa+bPDkeIsoKpn
wIvZa1xIRHjmPM5tBiCnX486uTscLTEnPtvPHyfERXXEIxGNagZz3mGNZ8+wddsr
k+vnlDtzZ5uvl48KhA9ajUah58Yj9SoeNB88dc9WOwsjj4Sr3hKfdqi6fgf3/wI+
NsxxraGK0epoTpnyKsEmOrVaw8A41DM4k4w5wbGtmctu4vwNNg9oxwusxeaH8iwc
M/xuYZ6cp9bdKOWkw5cvB8XMkmbnYaQzoXKFvarDKkU7+u2YgLm2cbHt63tjVqXh
Kt++kG6MFF5zT1NkQa+oFDBB9VMu74laDnODOjGwCL+yN90fZhrGTctmL108Kfr4
pyMj6Md3/IkDf2DISPKiVe+AOi8mcsuAhn982A2Py+es8KS2BYHU3VLMKBzON0x9
3+1kRfsk2tUzcNv1izggc+PKtOrAkJPi7O4LuHHJqwq6yjBdEeDswpe9IQjtKI01
8ryd6cY79T0dMM4cY7TEWJ+T930rXpD1948MuLE895nUfhOpjcF3Z+wt/90l3heu
I+NIFxIBfIGPiOhnnjEsD0EM8RnFbLwQ3vwaVDj7gbYg/UJGZLUZ+PubEYCELeYB
xcn1xBIsRjsyeHN/8W6IycfeUwpxBT8Hu1/W4aRl4IWgGT4dzb0jJPpMHb58I8+r
lvwUV5GFi0dYZHsHR8ePlDKdhd31uZjzbk5TjvE/GnP57vUlSAiEEiLqLi42sKsS
QVkPY8Oa9SRtibW8VQ5E9v9ARWlwGl7oDA18La6jgi2DlXcBXBFe9RaacxAgAb2+
mC2FH/Hdg4wvDwPPQFe2Nbc2AZQYNHwK63RyriRlLa+GmFB0vM1rylqVBifrET73
nGsadh5fBa6+ofYGOFyR2oZY6R0yehBGS5v2ljjNKDk6kKNREpHfquh817iUTmSe
Nctj8F6fgIJB4nrSmo3MtMEvC29jivOXnD02nKYWgCLIFEcGK4qVKgxVpnLH5dsp
Cg2JLIVAeidOXArUQ9xNaD8ply3MLFopIItnrBbnKFPnmj1e3NdF1efzJfzRpPEk
E7elxmsW0MydF0XYX78d8vp2QWv2+RP9Dz9Mifn4Ez18nKtY1LETVM4+rBAerGPc
9YoacXVQICKQm4P+ECIEYRxJr1bTZ2UZcwCa9TwQnYOXOLeRzS8fq2ISvESCtGvc
FodrljnIAocVwaqJ9vFVO67XnrOahuX4AwxbRxCOfrgofhbx+bjhpFQdpr9jjYDb
4dfpBawU1X0Z+/e9xmCDztz/VgzWtFG1xThjcp3CXUefR+dLue/RtqGHO0lZEEPj
203cWdCD921t0wJyJGYNNg+AZaGZeFv9r+OZH7TD3bRLcRh0KLpIIRncxBoHK+1K
divnAyfuPBnJmmyM2gIvE5h1N8D35baT5v6ufNQRJz58XOnvggt5CWUGAnIdefsd
4rpVFLI0cLdj3zUX7wjC7ipem2kDYrbN0kHH5Vmczvdvfa1GfGZePmkXLwOlUm5C
XWS6d18oJIzHmXvPaq0iAjcWArRqPE7z1LZtqWsJyqitl2z2YInmX+0pTWhyUpBk
K1dcJ5PZRy/OaWvUPCxKJlNgKCPK9MVl9bp+25+UPkFWRdydrGzRr/vr0ObDpr1M
4sYji3NlndlfYdbkUZh74D3TzHYkn/Pqj0rm1lDh7jJWEaU4C4Z6kIgGIe1AFAsT
I/fi27oKyUJO3/nhKsisNiwj+4P6rV1b7bv5HQ4W+gTv9HsB1w3U64pgSOyygNsg
KzyA5M6YMlHq7/+LXdQkQMUR1ReAb/SpWWZqzGB/KfPW/6S8+eFlxIDTRwqe4u4r
uA/F0lQ24yYZNcYli/nS+weY0A2vsmzvXzLK2C98eaqiKmizW8S++2foLdfFaJ19
jr8kOf58D1gfhzNI0+09CEp8LQLjz9VC/cvu8/ZjlWxktrmiVZLay5oJGnU1lOAo
MHdUjHpi8JoUshf3d8TqJP47Y+cIbHfbvhhxq3zBK3gKGwEUgMAzKQSQwQxvNtVj
VWbUjWz70NfBQnQVEGIKpygr1fXEVt2uUEFfykSzIFnPeNnuV4Ph3vhBgHYwMG59
U1f6SBVSQADKc5CVukZg4WISou9WQ872w1vFIYJBXYSLJaaJqftSFo1WZJZxARyI
q0aeiwj5DcuafUafRUsBNqsJkfge6tjYRrotE5cunPBwocQFsR9WHF38+d21ieBs
D9xRyoRJYPgRIPUVv9oGiLLpWS/YJXynF5kiCMnI2e2HvQJiAKnrkf8HFmdhaJud
REeemugwKyQS/1LoZQhoKYZSgQxy3ShrgW2gjdnqN3SFM6CUTQ7HTswGhytgCagM
K3/beUilkqIz39ODIebCa/Ds/A03lHcasxk6oPlb7TH+aHiQEx97NHrtBp5WOS/1
TE6Hoc1esuWVpczjvL/M8JR+Q+DAAnQEWkVOhrk4ni2W/beL/jC/ikMXET+xVoXB
I59wREpupGOsfM3lHVrTcNABOeCMc/+nWVBO5paYSxbiI34YT2F9FOqHOSa8PH7E
veRA1JgYy7AuNE6CCGmJiJMjDroH9fO38bAl80y/XEMMtpwsfOlFz0JrRU/7zclb
4uJf7YUyONt+9ib3uMyk39kjvUQDvB1c4/F/983BrObkF9YDIzw/EcJvJb7UQ+iO
9AAqEz4LsO3I8KOzo85Xkro3bvuWsVvFmyToa3M0mDJn0VKj7U27NcDvaLAxPoqo
gkp8jTT8UWC315vySYBSMf5KRHsRTYU8h/cFbNKnNkfylZ9QumhOzhrcFslZIK5J
H9YlVcIAg3QUAA7fRxaPm1ovKmpumDsLy1pnpD0ZErKCPVqjxrBT7P0cyyAzy4in
HfSJBx+DpxsIzIy/xjtWntzCSe8dnJtrN3gOX8Nl4gG826Q+FBCCZUH+lelYkfCv
TDG+iDy6a7SFIiBib1AZmAmET4DRMqqqBgNBrPyeIg4cAyiHbQ67v1m9S0kFa09u
+y79D3Em7bwc+exU3+WmLUz7VBgrX4EUoOCsb5Y4l+1ZLs7mNKt0t9+epM0isPzZ
ygWfl5iL8zssvNQGVSSILTBdGqIjKIbdXcSLf1m62cx/XsuABPt2D2WacxrQCv3d
q5GeoVDvS54mUG2y4eFfzGyuym2tfbu/4OAfyZJMrDvPjvQJkWVu5Ht0ckq1mHBG
hgyMAfR9ME5kwQA/OIe4xPntOPn7nYOaTFv22nowScrHAY3vjMf58Zex19FNsna2
sOjq133lmOhekhz/GjtaDo6hlFGC5z9mYP4KV4t74tGLs1a/EUgJVFhiDKq06spU
2gyFWuISxZoF7Nb+I1Qy5OZfQiyvoZMUVB3Y7vVqW4sld0DMgir/thId3ujCUyVT
6GsuK+sEwjMP0e2cVXIdK3hC/44IxRSGxY3rOKOWAfCc9OGdly8Asr/ON2c6ZTL8
NQ8EXPnDUsQn4u5uY+mPIKt5/Jgqf4nCkx90yw2Kt8UsH74dQ1mH6apLMQNEQsDY
hph0nOTRbNwaQdn1iY5PWc5Be9cu90ohDdhB7jKjvegCc1XMytxqr/ZLbI1gQy4s
2i6C/cN8elpClJFRlL9MA8WC2H4FmWYyyp144j6DJt+kW5vgcXoqjUQth8ihlUXO
5VH45G0O4lrtftMiCxykUVCls5F81SwZ05e9+ttmvCT4BanDCa3xWxkThoAtSUK0
7OeGF8SKk+6iAQVid0ydYaWanYPWE8QFfoKZF8tulCkgZJJOO5uqjR5dxNcoGdKa
Gg0wheHM+chB/zPypTMF6iTjyn7ipi9iU1tCq5H4UPp9yzJYC2Qu6+iAkB/kH1pI
Mnnpnk2KJoIADL7pG1pRbnApZfqFjWXlYCTgGJ4Xw410VLLgvMbQcVwWlJZmoN+h
Q767gBhqDa2DRVs5IXt7GHsyKU9Ilw/w8O+iK7Gq8Rr+X7PMgH7sdMJtyl2XSwuY
13brEGBsxMeS7DSgWyGxBcZDDDLmLbx1EYhSS3MIu0JZBJbT068LyaBWqCTULEK+
KvjlfPfRtuA2+VIqg4qz4CB5rNTPv4CSuQOJjGlJWnZ1hDR0Ztb+6LB18vRcimL8
aSb65v51BoOi+N48FSC9fF663aGWC0FeLvPb/dUsuins3gN3cv6pWJafTIzfCPG8
Eb1cDSqfpeO2G/mb4MsBoswAPloSniJExxV/ZlRuGgNps6LK3fIG+zpfoOuNuGSC
hadRnEch/3v7dXwheCh33c65EjoLCKYEsRj1L31//M1nQKNlHXliqNHsQdPQD5W8
1mYdxxVLVgV6Jc4Ltz/rHrbWXO4u2QMc6PzP6LA1oaP0AVRZGCRkII7NYTpfEs6N
jMqoC66bs+j9mIflwTixqg6O5Hgok4tfrCZK3ARZEqmDjk5Yz3E6QU86yXUfFeVu
sBAacyfvyPx2KfPMYm9yWBdi5WKRPZQqQ8piu+SWLKVd8gu6wLg5hEGqEN8qxToL
s8bCxlnmMeYAGy5z7kFWWACHjuhkhTfL/NnTzscJB4IWkSlhsLD2NrzYwj6TBJa9
etBrqoV5qMEriuv5igM3pgPnURUIzZxEbijvG64Yr1QBKfMnYNS555bOunRu0apc
3dmjkaltwjJK5wdy7ygyhkOhx/UA7txdi3IlxCrXZnBk3D68yfiggPjnki9kHDpq
hkA+azZTRyxp7wTzxWC8qx0DYs6AXG3nE5Wt+JWcng2FGMVLodR8fTPMV2Bv/h0Z
fSHZ7KtOOY2hx6WpgfIY4m2x6Lsl/dfMul9A/0/IFIx0T3j1MoRwJNnUfhvam/Ia
icSMvZjNyhih7i5Iy511lWAFtROyGQ38wM9IjGdhwUJpApb3M4O8TxP0KFFIMpuG
bNaBsA7BFCA9DTyaSG3S/uIe8Cdj4ODS3IOV27u8UDOp3IwhYc09jPsNvr36DZen
idyZ/Ey5z/1aPQt6ztSGPyRRAPi6qiLiGVdcag9bWfJ3mpAoro20vlGVgZXR6hrS
dSEL5WDAJvCEaLFjXhLFSUSKDQ8sMgdCEeB9FIc1bPe7tlWLvQ+vT40nC+XzdMYR
JQMaDdYUmQY/Xk/qbl0D/eAESu3fIzcRis1QOJ99xld82GnDCVZx9qlYYmV8thas
0GXNEsyynQtKRgHRM6v3bXwWFhJynXYe60FcHqjpsZwF30K/WvJ69gAjV2ofONQ3
S5thKiX63F1M6BpQxDFSp7JiTxYoXt1zVX9ysZYDe6a6d1gGUwly+ITcP8PLh2vv
3e/FeeVVHJ4pPSbrZGZWUuOwPW6tjGf+dxjxaoH+cU0J02hV40QmnLmQ7S1eGjXs
W+Rk79T2e0fe7htH/vTP+P8+Mrkext4GeOut+vmOH52I65DGknKxTX5eb9orqSGE
DWKo77PELZCph1HJSA3MmHqA3kAsCnbk0XO50aa71bQzEXGkZG5J3TcQoO6QUGCG
wBzs6fd+/amfV5RtAF0VHQV2L+QfrSHYug9H1pyQ3ExPoL948gXVPzlnLcalvUM4
Euw4IkMfWiD3o9Ck8JDTSVxVfdF65MpE0I1gr7teQ37y6CBN3+zC7ekdzQjBJmcz
eBBaYc+Vi5w7QAgO2i1xVcaJf8z7BehEZSiZ7SBku3r609lrN7HUb0iReoNOvKCe
P+VPjRoZRwu2TzOsKTTdBgxPtCesppalgHIx8+2JbF1vYxA3wiyGG5yslWXC94TA
RPM4FfgW3/4GmhYpmRApFOjRPXvZranC4PVuS5OG5y1hlACDguI3J59PzZi7EBCA
28PI6eU02EF7X749CB/5ktfgfP5kO2c6ApPYsnwNKvYfhcQxXR3z4sWo4x/sbzKw
NVJFecHczMqQJqBi//pHcbP5Xd7PZ536T2QwVasSwDD9qS0ws5mBvBeZpfbOT1jr
0s4OgAw7efhJib6rLCs/l1i/ev7qbW9sZ6Am2CnEWCyMzVmoAlKXIMOENgrFSAjV
wAiVFNWXuufQ/4HgLxu8BP3vj6OjBBj8FNNYkqkmpmBV1n6YrK63CXM0RWeRpspn
OGhkm2i/camsmPBm33OYZJi34xpEaTl+ox2tDTJ+07bE63LtoHtFO7Ai8ZJMe9Y3
4Fb61J9QP8CSzgIRtzNSmfHsTeCAqXXK36oFo81Cz6JlxDJtRAmiUHaAe4H15Xaq
PUUsDYddgaOVONsFEdBNW+R6+dhNGjvvJL8SPRRfPVuNEJ6yd2IczLiOEfv+2Qtd
T9f/LQvJN4SRo5QgsMOhPukIQWdvckK6GNIb5ZYyE1BUq9ZSin1HpIVj+RVbz0D1
LuqkY2wk3QGYfETB2tmb6IbyQuLRlyFZl67g56bKcp9g9kLqaldLoj9c/wuPqabY
D6N2CnAgbVEkOSdkqje80JzJSvARXLRSWOpsudPe7af0BWQGe2dN8TR8W8gY26Y9
6fnccN1CqJhDwDRZhMXSEPgLcKKfup/Ak0etzl9ky5HMiemMLCOrbij9agqRlhzf
DbMDW51nawP61ZpLkiOlEuTlweaD0dxjUSwtF6DOaLhkz5WpMrMAIJdV8UDgChQ7
zu9QQDxYRE/5wbHNlsx7nHyqM93/zgehpNlTp8GkyCfAI/rcU4gd1F0ZcKZZfPKO
wGJdJy/LiSyVlT2X3gTsy5sTfT/DB+H5vf95EdugWet6tHVOPtZBBBLBS9xCel6s
0AoyoZym83X7PH+ZgIMzxDGesV9T10BNEWmTA8j9KBF276mzQh5BZaL/qrrRDWbV
w8Y2LKzqwwroAACUUILnK5WZvzJ17wPD1at9+f2h5NHSNqBr24LTyJn+uYX8Z7VI
IAzrrvPATnsPSb4t+g7bLwUapwSRE3KzhG0UkfL0SNzxU8MgpV/aWah02367AAYv
l9mOlGWvwyHmWzpAz4wfiicnvAog59Yz4Ah7l1SAvSb/o8Ne/wNVeOyloXxyiQ7D
aIlQ2LO8InF8vDeOnHjswPY4Up/4HPbNVGDvU/VI403Z2GPFniwuNdCd6Df0aPSP
A5jsyZLWonZdEA/WESNxTknd6XD7rJqdn+7FjPtoiFG+w8wNg1TUaHoZCDa5RvJP
Ib1woC82xJfOa+24ZJb1rjV1jKxN8H0OiaFNNTqXjVrCYIrXo8zkiIuVSoM2UhLr
fMjkHaELsbee55BVbHRLZddU9Pg69IBtBzIRPvO6R/iT/FKrE4Ujp5tYq7hBFZJD
PIQM6knj9cwtCfinU+JezkHjNPrfmEqVovMCU91fh1YvU4GjA+1/qXr0uV3wnTi+
B/wYuAEj785cMRUYCAzE+72AvWuJq6fgRSIyse98K2eOJ4/irSLuH5WmHxopGuFg
sJrfYNU1S1ogqoMdj5+vcthsL+ceT5ngghZOM22xUkJoZL/LHR3TeVadVfqmxdXo
u8DdOC9wxjLkXW0Q7fDN7cptIxpMy91pBAbkcdTUvf9CvLLA6bwVVBRi1+9HXj+a
4qWKs+OCVpH+qkvkphcLRVWHm3EQ3Ug13wDk/GlrguGKKoZyDymjcPyN7TCH+SdT
QHZm/Ax87ffROBQYFQs3Oq7zZLyfa9NiUqQ/InE+QuztIxpBQiU18awUY/q6ZRFK
a5KyfGBCawM2axAqTkQshYHOc5InsTSENZxUEe5wmqFF9NBdoNXCwXt+Y1UXSb5O
4NjluMWXYHhwnGLqr+NEd36FtYVp6GSrrqafXfCDTK/wPfuWx6v4UeDLgcBix+qY
pDNiMmbmMT1O1C+ibldQS8BRApmDl+ok2nYumfCOVWhmhkrTcnz45AQDt1njYMoY
zcb3uAoUkciYWPOQ9PqilNwwqzU25w8m6d3QSMBo1T+Q5pi6Rub3WL7PhYp4RCqO
bRXP+xvPha60LlCJQ7bD2HXETmjUOAS3/VwXpx8Aht8Hd8YWsrgIoPw8Aw+G3pUG
gzRoV+5vJsE1vpx2V5crlMQ49BLpVoz0V51/rxxcK9ifRVce1198acx+W0Jw2Mje
OTu1BZOoisAlHxeG1kKxECGNgWmbeNLqYu4rnBF/0pCOgYlcpXpD8UapSxn4mdV2
OKjxE1XWVVGD6fCgsvwOHXrJq1eD5GZ8I/NZJFk4KLlytkYinig43rmOLyWoBMJJ
D8AlZ5I0LpeG/2Q9Mk3OGpOFr3Wime/30plj3c16/ouVUKqu9yWOGrDQ65vzpqpV
1eLXt/IGfOx678L7oK7kiVV+pJIe71sNvjmmlhBTG+dycYeHxEiAkE1tJQUTyPS2
FQZtU4y5dHEA4IO13TeAQ1FC+ifrVOhvFvXgWCyIEdJmmih9DIS5UK3e8X2aWR+O
NA6MijMTmvcfplm9GieFFA1n/lYD3IfSD1UDQmGGqn+QkqN6nl5IvLYC8UuTFjoP
CO3jS+JLGzyYYHBvFBJONUcUt3PGpkjeRwpydHN83bO7IhscVO5eyFgyF8SRSUhS
8e4a492L1zD7RBeYAo4Q/xkKF1uN6WXnmAK72kJsY1Y+i+XVUf0Z0xHbyw7ucdJs
RtY50ivr5fCjJkzRZTcSpAhCuT2Of8ewuSmOSB+yiiHejOMs21AzCGeYubAzje7o
nF2uM4uWWBQcVU/aSseHuS8f3GB+ffM4wTk3QjQ8IS6WC4AVIUW3N4s5h+Ze6JKZ
WefoZgjactSJuZU5Y5o+ssY+8y+WpaVBJZhFB7Hq4i+KKVZycKYoVldsxSZXNk6g
6Vw/xKN2cjxmwJRk/bobNNYpcxE67y6cTfwZhk+7yvezM+DYufiFCKPvSVBm7n3l
yR6ftL/Zs87Wrjr1UBun6AtEWw2Bzeww2WpxURXZ9yejlyMpbLPy1KK1e7HLCbhe
+9gqy826HdeoH08Kiyv4IY7J8nNJslrQLIiqnyeO3Wj76p6gjEsDJJlW3spf843O
WJm48EfZKhKoeUH7f9EDgrc0SfEEmp/GycMl3H2oql+AWN0QAInSElVjVjbILspB
IlGJmTntTVDiwFdNg8QaBD3H6KGqKK5D0NmqRE7XjV/1h6KOuLzYihflhsYjGTBY
ZG9JE9Hr64s1smwL6kwiE1oyoD9HyF74/11BdrUuchzeunHoH5bGaEEzzte++QEd
Rbeb4MbEJH06NfHOEy6uRbPg8vuQ2hVIRAutBBuIF1vOfx3HdC7wJpvFl5iUei7J
5XH9XL/Xe7g6vvNPO8/5wp5Bayz+5+MQWU5yzBj6YkHo3kWhM+E7Ip3q36F+jl3N
EtTarNbvq6b7yERIJ+z8n9o9W7MnbOHzmz0Ho3hLHxvQ9O0SoR96Y6rhjUunnB7P
LriHCf2zrmMZkFuhI2lmPve55levYykkWMAro5E9sLoYB7XGdRsu6yf9HCw0xFjd
whlfAS/aG3kBJsMq506KXIgdx32xEKhdktUkcMG5dKeDjbKCO+9aZZP/EzfK3xVx
yqS00TR5F/apY4jQGxvX2J5CB95g/jNgaGODHg+dvnFRT5iOlq+gYN2AX6Ro1Qis
1i22z4nxfc/OGtw3hoVQwsdq0urjUmg9nRmH50ZBRtI8FhQDY2U9zOAFJ9BTLnli
VR+nmjtGmvcHX3m/Ii3gQBPx94Tpz5CjtOVAl9pPmVDyLq8zVQfpTZuDQRTxlH2m
mr0eV8Mmk1SpyPxtXzlpxW7ZlIicv7r1HZ6iwzgpgvXnNjyrxR+entTBGx9beHcn
ytSgzhWUWOCDnwBgbVZ1VLmaILQQDKbLTIyZTHHNBW4FAHXCk/HXuBkmDmeLJBOb
TTsm/mYz1m52YZpPPBeS7c7IbnJeqatJJ5DncZAWEiZKoKn7h4m2yWyCDYdmwVyw
JnFQULRqSRJaqKmLtEom5maT51SC4KdFFz0qcnxM13cuyzrw8N3qEr7e/4qwUU/T
YCBDZFSim5v6DMzF7pqaZPO+TJSZCw8DT5gwck0KVBO54ImK41IdTJNdI0s+JyHq
FzDWjT7Cpuhuj2b3qoVcJKndliAFpZKHwK5aLA9koCTwhm7fSmITSeTv/l4/HAJR
zEdM8DUwWupZjaasIjnJRNLAV47IdSSX/ZFq/hbNo/w9rMIRy4hqjGD4qD+rZcK0
F+Mr4o35bSHxYj3P9QiU9KkYFdmyDeZ2bqeFKrSSRlzq86M7bc4HyTu8e6/IZpFK
UsblnLpetn0GAMi4qL9tAL81PPSCidDugKqk97qwUU2k6ArnALV1tB1r+e4dW5gz
0/SVOXPughEmsL9crNq27mdpzxmL5S6aqI0GKskXQAddAJNfI5uhIp+IrviF9o7M
Dv1Djy4KxsCsmjl5iwJ1XMbuw8sxMPdlZ6D3vWNY6IPgBU5hjshaP4ztzRMtSGWq
0tIRHN8migazzeurMRZJp1c9uGjXV+xA9ZboLtqQ7tINwPkS7A0vs0O5fKaj0xyJ
OR9OHsa33tngIOfaYyUvdcSYrM7Lj3X6+JUCHE89GhIz5TT3Ivs8mNNlFBV8VED+
44SkwG7PSom04y9RLhgvrHAJxfZEI/cl4ixegb4drDS+k5V5E7H8UpK/vjy0/lxY
aEYcfZMF2OaGL2/kYTENDEshy1IBL6t3FdoOA2gOo0/MOpOYtRElyJzjewJeY+zU
4lEv+41jl0Fm9uqHuflD6ebqKykGOE6J0O3ymiXZ7u/VYNw+DNu9GxDMbqkMlMmk
e8Cai5ahZC2jJmc245I7YNPaPjRBw8/4NhQmVnzF171kzo/2DTdahpLKMn7AgbMl
Riyfa1bJS6vEMjRPWwiXweRLyhVtCR45zCwzavzHa5C79m2iWzCR2agBite4yAij
4wHOwWtCX4eiusdlCdJVxmYyqr3iNsQvMNgZ7iQgqWQce717sZbc8aESmTFb0PPc
d13UxN1sZfkIJQQx1Oc36vVbDvXKIRqqGNhPa8NVhgGadXh1NRrJAJ77Eg4yQM4P
LD3xdQsbMZW3vQW51NBXdjWnJy+RTJpJggQAOzMzxPpyoKH86MVapb7kMGrxfvc6
AqYfw1V5xwFsHybMsMkPwDFvvo+Zz5dFvceO/4CqA/Q/dHczQcWyIdOBMDj/BWNa
IiG+7PuXV/GlKhw6MqkEaB+xzRTn4eTLFOCtpnTLnic0tI195jCxjd1RbnuCUR0P
8O4vAHRleC4ZBWIgg2dDsri7hnYt3pHG7DjLv7FE+ANTEF+NZgB9O5ctRyKoUmWo
98SW26oov4gYzNaVyYpXonYBeOUHJ/q2U9ci+AzEPvK5XTOfWoigsk9bZfrRQcEu
ZhWcDzIlXwy6U6PVAsJyaVnVNgAqk02BPqxKBSd+ZtKpRawAgXlXkNAnKr3IOPqY
5TcY4sseKn2mTua7XP9DPuFmQJDz303RuPrDKqIvsAiZmN0Za+jSz2pXV2HjzszD
pSa+W81Zx6NpmqUThwuksVzd11EpXkDYLny8ly1PFDpMmzMjo0Zgy82x6PtwP6/Q
Jfhzava3TlqlA0ww7qRizXO+RX0c5kBtp4w3vvQwMh380EuPOneqAexbUg+37ueq
ptNAGP9aIY9XVdgf0DqqZwnrB5QjtvwC29rFWFUF7h1fZgX2QBRjefkC/8gBW+Jw
yhZiEeNyk7YbHetUzTSRZyyforBVZLCb/qrdpzHEq4cRl/aaKHkBBNeJVdasSicS
0dHgjEmof5ANjZ0jr69f8yWSGmgvEsEkQioWds1kDyctirEBruRgcMpDr7s8OOpb
pjnrqitg+Hag2U2xWML2NvLntvQbNni6bxnd91xK8zB7ZJ8z5phwEI/kifZI4ROk
`protect end_protected