`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2320 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
mGnK8YPdKNkEYt8ET5XrlLr6Sw+mAYZoAw2H5ncGSAp5OfNHUj2h9sDojqTAwfqR
rcVE8tcT/RGJ8T5SeizIzcXZDZOqBQOHi3drDtLg77gPgh51ODNXLS2/kmvobYzZ
tODAzc4+Q/CA6DKcV7UuCrw49n+nLAZVj94A6Q67/e0ubGf79ZRXOAV7Yrf+qVkO
WZUPw0TOAyEdtaS/w1N0J0qxnoBqfI4QRQ4uQt9N30Lymv/xb9KyVSWoh8OW6X8z
ODXhYEFh78yEQXPsEKJQVp0ZkdL/EJ3MI0a2rZK7SEJY2v5xmztDmfW0Iso5j9Ee
OI0KjW9XyKsLfpORJ18FLbMyrp70dZ/RgzAn9Y9etNWGZXuU+OCY31LT+nAl4ho4
kXOU168bA0Vh2+dVZULsE+JWR6V28qT690ySGLZBe1MjKhtCwfYrpZJE/atAHtHY
38HeKu6I7nQZ9EhqrSzzKtDLeSJzQ5QMl3oeQ9mKDJK2C2iLmtenfSFTp5cjh/Jp
YeoSvxz3+2Wl/cRhY1xys9GZ4ZlbVgR3JTzTUmeQHPDokhxw59Nm/W1CFeI72yYs
5jB3ccxahzOgZ/MXHFddlrH1blz3497iBYIn9BD3rw4hzg1qUIJE/Cy97tXdsFcO
GpUxEgXS1AkSZsBP5f3y4uQ/BSVT9BNcNSD81FdRraSjyovc75y5hlWzwi4gpq1D
3SafPTnYtywctwtTGcTK/wvo6KtT+iFldYNbkbMst3HIcBJjxiD99va89MwXmnlR
FbYqGU/H91Wd3EC1Fptew/awym4hKaOx8Ee3YlmE6QKPsANrjkCMibD6ZM56fqbA
CNdwdteVI4G4G0uSXWuPjLw3PYwG+4oq0TVtvrbWwLWhb/7WZuJvizQmGXqX7i3w
h3cH+EUFLlw/1JZfFrzlIn7TvjyxV6hKvjWq34lcC6sXss9K+RoTHcncOT3nWjnQ
Hivw2Ya9RIe/WSClx/fWhxHhSWdz8UL/fKIdk9U7DpUKvW72c6JvPBG0zSX890Rp
A6jrqflpwMJH5uTGlWUwgUWbZogemXioWTiOgAdl0Ff4ofxgl0RGQhXrlvNGsx8e
wggqiVl5OFkY3WLBBi815N4PimQRe6/gA5XkvnRfTdaXYsn51CMjCtOV4g2uYeT0
HJZ3Cgc/j9pWydewEkL+nvtTDeEGwGI/lc7UHIFRBoihtOJXs2+MWN1kqvAJVKTN
SkFz/GtIkLjyQvBoR0kOaIW2nw/Ps/fUdeAeiYKT04TzcZYYHnFVkbjdasaSAvgW
IikOn1ZEg+22+vDK5iY0YvL99u4zzB8Xof1m1bzKh/P4Rz25kQIDWiBvQp3t4cXa
DrCwfECxHPT2umDJJBD9F+aEtXkAipVHK8WezKr2dattvcURECQbJi5lBFB44DQK
366iDkwft1kGYYDZuPkXxkxzTnqh+43UZpIEzSwzHKooe1Nxmj3xyg0kFQ99J8AE
ZIm5H3WiQZTBhZK3Re+UP59IYMOwyykJkb9SI49rsGNsmWVg27LWFul04/cwauEu
M3tXzmCn+HEgjgQV7Q1OWt3j34U2PAeLagEw+cfw6tuWZWQoW7F/EAvvsg1KbItN
aqVMfUuHGUO7uyj65VtwuoSWTZbtkp2tjZaHqQmkxO3x9ZjaQFMwKQ02CFgjCtp9
QxPPj3JmiwtbVFc9rpaH/RgEdZo90f9rwNljht5CHc78pHJw9TrR9eybOUgSIqCS
RDQzrk+qB8ozD20E505ATimxBe7g9NqIiJHyx9mgoS0v2y9ql88dzmozuHQdyaV0
ECnpHldlBrOEKNuHX0pU6hnBk6r9ET4Ls1d+eMueEfCWQga/5Kttsi+ZwqaLGJX9
9eHecNwbNgnPwHkMrA2IXEhizLYApI2pAl6rezCB2y94nXyhLQNCS+ZTEY0eBmEW
ZVHJX4In1EbFjRbhvDJtJ2SZDT5OyCOCUKBWBEoDp7/WVDJHsmVdA3a2UDP41hIE
askSsW1+LtyHMy5pQFMbbBNxZ/3KaEpXaL1KCoRnjj2WJUY+QKMoZyK5yHun9kQ+
sawu3f2nqflHsGLRlRg93NMHj3skr9BMhGtcO2Sx0i1MOnmPlnAlhEevveGinWr+
GS5mC2sw3zsJ8sJS43OSlvJ1u6KAe00G/ho5Ws/FXEseZXDoWlYlsnKOlzTA5AJK
cxyyskdl5Sd/ubq4n/UMohIyDBz5vws3mcjWRD6bcqs54fD8NlEeixd3ACeF0DjS
tutl/43UF+Hxu/3qGM1T04jDwBK+hkgbHBtXCxUThZWBrfPRS7iALKXR8I7RRKUZ
6lTH8yW4zLUVcssY0s6qF82EYdx9G97NTKY4f9pZB4scZZiOdB8cAQw5HvyX1pKZ
yAO099bf45rEKN6dApgmrpXNZ1PERdvwf1xLERQKrZk2SCYRH82JJIQd97f01Kt1
3mYl2LJ2fBXLIcmzC4IhI47oMCdJ/MdigXqe1KE+1yHn4479N4I3afRbEGmmAehM
fcIQMVkQ8nAwK4Amphm68LO3e5wxyujx/srLED3o7Y4fkfAh5OaP4AVax+9eLRlb
BNL2BsnrkT8LbQPymp6+3lQXiuZfeF7cL0CvxpayDToD1+64eaJcMNfz0JBDppPv
AYf9BEqzMn7nllrDiTKSoGsHX34O+Ww2Yhnc8BCiKZaWU3x9ym0Nz+4C93AxTWQx
c9oeO5W+n3/NOYd/SvXzaZsm5SnjBTPgLGhg87f2tYEYZqb1noyPG5to1Z9YeROo
oFEYT7eqDh5Ox/9oI/RDl7yvZa6zS6ZwsgFgzq9/waCESxMBsLPxVOrppeSEpV8D
TWryPPIFmp0awk+nUxr8WYgxmd/Hkt+WCxSzhT/GOrJNUEB3/rBLjLxxGXJP3isA
VF+uBMJLN1hTXyVGCEnnXOg7YnxcztBvx2KiqGyxoh5Wm+rUaRXDIza8/hGXu9AX
fLyRrRVOY+fQuJ5qJygBMQ==
`protect end_protected