`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
K1dgx65eVu6lpj9nEzu2xogy85+H13/M8k4NT7aQKerHb4DtN11h0rLZEeF9nyEz
jw6duha5ai4QsSxfvrIGwIicmDkKMUTqD5yn/4B5r0x+gmjPE1PBEYqY0zUrJ8ke
PIeF0VG6IGSIg1Tat43KQ6MU4ipLhWZIvhOBeX0Nze3Mf3KDI/knHu24Ly531/lx
zR3BwxiU4+NwVDugRIMSl87GI2EtfZc2mfFoDkHCTjb5cVsBzkaruAcpO2U4TE0h
GZSRUgpYA9YhU/dig4w8R2KgXfcpsNz5HJfJ4DURnodBVABy+XVY/Sy6BbB7NfBx
HLpRYIuCp8GxTnDQZqUSsvVgQye6iUZVPZgQN0raugFdFOo9T+3ptj/STs1UmQFB
wKtubgBzPVYH9JKMzKkxO1yeoomT8sU/Gkthm+M0iQIq9/n6Jb5uOkoTVJAh+YAN
sSXDr1R5kxA6J9+ADBUyFYoT+aY6Ix6zAWZ32c9RBDJO76+h2QKDT7AOvzCheuiN
dWdfINf+8Fzt4srWIP/CaXCTcIJ/BRy1Mamimhz2I14V/yVX+VQc+DI31SgibdWW
PTxetN8RRHxzQW2EGYL0AXdM0zV92X0BpnqsidpIjTVsv5JXxHTABEatwXGnbDLv
4UlIeDB+m2JWbvGEuKbh4+NhJB6MFOjsLuOteId2mS7g+Mq3JOILysFCzjbBFQoq
WvBzO1e+eoi0WOnlLvCKh8Vx+UzmzSa+V/s1BPJ/QvDumfk13wk6myj6Aw0gVWUu
pZJuxCC5/8T15GbI6qsM24V6gfpyGF6jWU1J7BsEC1jxIaTv65/hAYcoCQZqDHai
lmi4BEI4yu7BYVcqNZ0CZ5k2sQNxgZQ7QhHfoDag4VUP0jKsG3pIIwYmVJgmzSjY
RVFPCnVsTWovxKDzkrwAgCNzncT8wmHYA5HtYX3mw6Pez2QAxBaOxA+0C1LnMy7j
0ge2efwHPSDRY4KMNAQtCaokhINlyb+RXp8ZpiS5NEmELf85X3K2JuwwxQW41FeQ
3auHG+RkJmvi6LohvbZ4DVWixJKfbhDSclubFaq2bhK+rNbsLggN7DpkI40ohgim
iZkH1NgmCwsOZAHxFvcBhtEc2CmDzJa7hJznyyXDMKbL5Ygq8SoJOp1XXw6w4qfY
pin+2K3C73Qn4dZcmDOaGuywOlEyFz/TNuW7Q/Jsy3orBeGUngo97rICfcN0iyCK
u2KJzDciYogoGUeGd3zKQMQvCv+L/oDpl1EazRbbEPnghQ8Djter9qKGnBm1gmRh
RCHQSPbm9s4BySS6phl5lyYIriHTn0H4cjFzm19sY7dnWOgPXq7WF6QzulCHUtL8
fFcMVPmFsyRS825t5LYNlOcLY7i4RxP/zgRRwr4smdlQXs/4LUW/QsKMyIKkWiI8
CaTsPQoWIpGjRCApOcGvV+CxVCfyIYo944y7CLA1to/wXdtPlBZg2Nxnscjjtycm
abaGQ5dp8vr9zmaHVCxCG0yCuN14zV5jQ0rYUagccoN7+q7MdddLniojc8NIs1E1
LfXQiWDdFUwfE8D6Ev4AV/UhHPZzyY2m/fHPzUZODCv322Ku+FUJoW7a0zL7nwtY
mgmq/A9g3PY2oYfRwIOmK3xbqRBgTG2w00/EOBg9h8YIVMx3DkvxJHakm8McClB1
I7f3MLeVHYkS9r5BG7cWaS7GgU45+yU11Wlc8cDRDtSV0UKJR8Y8WMN/QlL6OXM1
UWaaTQ6OELoURURGpG+U9qrH8ObWPA6miulfgHenGBnrUKvxzBbXYGWehBFf7WTa
5OeZONqn6v/223qVDEVH8y+1ne6f0hcUJ7t7GwuEQcjcCvkmJtr3j0XOLZrNZmhN
ofuCOgsdFCUDvL9g5Ld3dml8GwR9EQRS03n/zf4mZBlHKuLeO/e/c5DiXiqL5Q/5
hQ0hKl/F/daDSppgID7aUE0it0jIbI6YQdaCXi/2ofxT/8ICNQHSzJ3pQamIfGyI
w0V5BhvptJWE9TEac5OA2US3lKcgrFZPJykbwrRfRoM/hglkZy99VgzIxrKIJ2Wa
2mNR33qUmnZYjbR46WznUGzplIIrHUGmTQ6AOhlFd4p7WZDIrfK4Gy6tfn6kpDts
LE/+nWX9NjE0bn51f9ZLPKonJK0kwT4UUiZkXe1+yG6c8OAvAP3o7MU6t0sSZKgL
54FU5fpfhDk4yD5bNLUdY4sOOu4xKiG/1e9e2tCZKqWZi7nfKYAo6Fm1HHO9QONR
sLeoDbzTy4peY4hf4l6HHP12sh/gdv5phUEt1Cj0SdKZRDq84peHOZ2Kp2l96+H1
+3o0co+Se+6hajfUx/igLUic7bxkNB250wVvh9owIn5US0howLYzmv6iwudQsqT+
2BqoNAjwbm182fzkvY7dHb99YfYwivoCRGNwQQEl8UV30ezv0foeP/Sbk1rUZmc6
LKuHhMSiX87Dut2/LnBZlGGnuOGv9RpzrnUdzq7EQzYTKZj0hercrksF2+ilCXeZ
JBuDpOXgz7KoxBRpvk3B281qsVW0qjmaLoRmO6bMZYXEmPDV2tsY+ZsXa1W15s0y
syP+EldRLeERP3ZZ2nlTOK0WsgOhaPa+XdnaOqNiE6N0CP2hdLYQ7iTTHz3qVIzW
nwZXvAa1f9nAfFxKSrUeI/WveaDq69vobREUTQdvP7zSh+d4KvsWfAC7DMIQRXVP
7J426NGOeykKImY7oFJWcFL4BpE7UxctJpGHKnI4OshnEYhieYr9VghugW2kpSIT
7P0iSVYnBUbWHj6B27NSF65dqXQlXf2qga9lXHC6+Wj2UVVseR1j4aFQ4akXIHyg
f3nOiGf1oY5920jfHSUQ1tv9PPb48SSUVS6IcHX5K7DgDFHxp1iIyjGVOR9KbB4u
RAYggpMUUvRvOtTloy6BvkTVzPf2eLFRNHn0/fTDzNZfGYl3yLfdMRHfHWk+T+FL
ywd1nX3aBBncw/Nw79RiB8ZV+HM7pQxKOaqOLVju4I6xW62hsjTi6/e5WqoZrhUB
PQZKzOz6T3R0SmKDvpFME7N2Z4nKNO3naXK40Tg1Y7y9Gr4TjKaYPRCZy8leO6R7
LoYuWDj6A+yS45ObeMY9+muuFn0Jiib/KD2Knd36TJRECiTXaEBLTW4/e2FoTcDS
XWqrvpTggTTljXO2K8e2jVPSBjp1A9leB7ZSzsohcKWtXYH0E4iAhlrh2XnylrDp
IJqDVQ4X9P02egT0u7MUAaZKpXViN6mlAxCYO6Bjivjts8EZUHlqhb6m/vueLwby
hNHRvECyN0iO2RIlnKluV6cWTEROCqllCWbhuFSXwdFKrQfdPTBg9bUBHf0fcCD5
DJFIb6udUDOnpfdXM55F2QKyNU1jmkGfQvRe1WYO51aGZGsr3u9PUTGA8o4DxWpz
682cRvpTN1NO5F9LMEL4kpmfG/EaLaqNHl4833y78vEYcl0wnllNw/LMFE4xKt4k
WrMIc6Pyjju7T4PM8hauHmR83KEcBJEHpYZlz8FBke1TPR1Kpo2WQlEJJcDKT+20
usK2LdEFFJA+oKxVkNk3KVUKU3PBMs8h8THcJvnA+T7hKbzQQIywHApjAmHdi7+7
iALjIvmCCdcwwQy+h/S4FjEdo/J53jsTCKaDf07U4Eu3R9XdQd+TOlUvxH0JDJro
dy8XkS0sfidFEoigVAtZUmFEvT4X/Dqlz6WglRUW2xB8v4FJT45ZCzyZv4mYmsxw
uLygATsJ58SamlqoY/nBKv7y6NKVCO35VqOWqPJyLEs5BT69pFysVn5rzgu6Ca2f
W7ElSWl5Ffm0BC7yiwlfleUrGdYjsWJjK0VrEsR4iebAq3NZobLP8hnwRaPEuJyw
n5a9WhVdmsjfjP8wr5VEyhMGw9erkNzYT6PpRKC0++k7AcESQtgXbXtGHFemmSy7
hegH8mDJp6BoLlLr1wNlzfM4NozsJgkuE+S0wZesqlQecSy3ciKWTgjEI1gL5L5h
AgWhO9DQ+4NC7Da+zdwTvgS+QvtoW7wxZeWJSk11UR31+iHXG0nZqhZtpHj1WJ8q
ZBKdl45GF9mP4SnSu1FQPqxlNpn/B1VD/AEC2ReRGh+qUznSJ+af03JedONL86Yl
+8N2TgpWwSiY6o1etPp4/nYBRxHKKFr55xkYEYdchb+KxKby/maNVXV8ziR1jIKt
Bb1jj3VNOgqlMCklkTG0Q0MHLRt+IB/bDCmzpPji19ciz+cH3TFFlqt51gMyC985
8dSLYwDbYvVntoxnu9oAMLrk98MeOjLKY5v9e6p7vtji4RN2a6rukRIv18+yWCb5
2O1UIce1sVd6SM//4NaEV0nswfscAQx+36wXGgfvzs3pWqP5KLtUvVqLPSYGRoOt
FolBwvUKyjGbQiWihKhvBFfaR+LB5AfEny23CCwbTx/Gr7Vb8lPoCj1AsUCOOgVh
AkYV+z4FiscIzFFCJeguIbYuRiTw0mMLzfZOu72HRHs6IojoZP0lpkRCAWSozn/n
kmcCbwusb01bpssaXMIOR5i2AxS7qhJo73JRz3f6McR7vcDcm3bZjmzejyMJZYJk
Fj/lJGjGYmuin5S3JiyYJRtLnNe5AD7A+MWGntvWFLUWEQzQjTM5QN2t9qNF4mqQ
qAaZSBlYZ/2m6Cu83nzd+6rlJne3Uof1KwSbdzr05Hkmg0Yf6D8KGvecA2yUcpxD
iUWhQP6hDNPzQ4sCnbTPCuDZ4eleoA1S5IygtM8ue4Jb6SvACvT3JQIhOor6sSOD
WuLuDhmdQqw19f7zZxmCWCpGGtPFHnFC8bWE4ZKtFszdB789zssJjs33v2qMWE4X
G+H0Qc7Cmoo48/YWEh+IZobZkQaSswrVS2VNa7wwCEGbqDWibabKiFQB7Qi6KibU
GtFyJWv4hF+VWT8MPOT/RF3vykQuRNuvkvi3ND9Clqp+j6ES69fWgN11ECKAuAmm
i8FYiY0NANtxyGeOEs2SM9Fs6qgLl7HLa5Dx+cAHFYjMfpvjmXwT4X9qGq/CmHTf
Tf4XyI/lJCtdcBKDIzBBrYIFcqn+j6ce5qirK2SVgogmUl8wIZEbxIudMngUFJm1
JbZ6kbVvqKaA7egpkJdNytW+OjcJImO0Ulbmxv0PjdXEcxY0X599An8cB/G4f9rp
OCe97aD9MO4H7shD5Kkyx+gvCv9Jeiz6tubED8zpx2SgkDti5l2gWPK6n9ifIZVQ
XvBP259xrAxiEHTccs9hporQ2wlmtHM26N93zazsUi/rt8vAlXYK/XZSOREG5n0S
iB6a3IjZQrJwfD8sdBDpfEmqwerBWB/NqQEmUS0inwLSmjRM5JTWe8or7LH57rwl
uT3s3xlbIu90+Ok9HHZG5OZf1+0WzLUcJLvjo29BtgkDcviwUEhnOiblhU1p2HWs
4xeRuzcYRT3DdSgdW6OP13+CM4YfhYE6PTabNuc+IWBD2L9/zZuqDy5zSs5CohVG
WCFVpRQQR5VFADGVF36WTsDqH2vreqXao92p5M8Eeey+fLk1zLrucWe5wPc/C0B2
cJ162QsvhIfAy+uHTZtCaX2J2kW//twRqLpryb79N9dH4aorI5iq87J2uyUd6NPD
xaTN9H1LatbVe/d3UlyYuNBQkTrM+UrsLY+Zz2WtbEuU/+tYGPJIMm4SKGqIg2Lz
tOoS03djUNdJo25zeTArv+S9fA/X4y6f+cIoygMSlmv+y3vyYlSRbCm+/z9DokD+
jo6hbEPs+DCqycqFnGPt/DWV1r/ImqzeapLxuD6aX/6LkXRpkBwnLH4bvKzQUVS/
qlNwN0wtY9ZWYrGXhsfnqXmkrYFhdWz8gray6tXF1WFw+3ciewk7PxEdrZRSryWU
n/laPsQAAJJ+x/Ky7L0pj5plsnc9G0XRTjIF7PUQowHLch6IOkxHxuFL5hQcWdS8
ehVS9nUk8a+Zy9RndXOiW7QtdRONoN7SnOfdzdNj+MAT9oXpzbg6yZCjqEF9Y1un
7rBEp9f+L6hTAvvDeg0tphf70cSMTHKt2uHmRBTRvY4g6JBjNCWJqZQfhdQYVKL7
+j72yjVvjd8e7HRcytZFlGfAOXid9X/Oq/olHnad8NjR55NQtFugNnjTQf+AfsxT
aHFZE4BQYPoylaejD2Bbg8FqKqk/Xn8OGTWzhTqCrrAXzen/lgL/IpEAme+7cau3
kbG1P/WP0PzBChX6lZSdMJ5v1bTuJL2OQ5MUblsWTACIW3ZZ8aAuxQqCWV6TtPzp
F/7GMC8lc+BPTHoOvCRkhJdxuTq24PQGLMpvyX1RuYqOTiQONv3ELNVvf9sBrkdR
ScSOzLL4sX8/dZyMDgpOhX0nH/iHnxnKLJ8MqWMhgKdVlJW7iYjx+XDCJEBAPn/E
0ulNxrCY0nBruAkI7jVri+u8UhVoCd6HVuEYugYxim1fRKuUjhEYA4Vyaqv0kLtU
mZjB1IIpeCo6MJMB3pmATFvFyLnkcxGtCbCJMkZzbJXOI4gLPA/NcumOqmfDS6vd
YQy2YQvezmBi3llQsX4hbq9MExsehukhOAKj4Y1CVzDiguIE0evLDKTWdlwz3S8o
zhYG+uUGIGQAhJD0afZGka+XqRfrxiJtNG7Jq+oI2GQoq2M/DWt+0pN/aWKxAAxO
TtSKMaZd7CE2L/nXu8AnWPrEjnMOouLdII3RMN7fLGGt4zepHgei81XrlAbIra1u
3NWI/uTo0olUfisyqw29odXLgdT9FQmlYm1LLM8AErYKssSnkb8/87MtVTWSySDN
eusaC8KDXqR8OcKYneYr4HGS/xzfMaofYatxczz5IIHfwWwOfBlFf7BErcQTudS6
DrmvexqXlvxH0+5mNIN0mu9xTZ6dlYfhbdWwp4kDmEjzqsfDTwNKwvncWkGWdD9j
sJrGSS1prPx6Dln8LtNoej2ksb+mVKxqQrxqKkSipMGj+Cw9/RANZ2I/YCG6Voae
LV8NoBrQc6Bj+SQ0UAd8s8WL6TaNeputJDawP811YCwBeelA3kxPgXgJ0BVNNl6Y
4LtHdkrIjpi7pcDcK2MnKBauhVMHevWJDMUNE0QYiyYe8KhFm2oHE7s0GNEoPRN0
qTsPp2QbSAvAy6IdCFBIimJs2Mgf3MF0iLhcp+kAQz0YizpqCVl+NYtl1mO8PHyL
dvLy+xVb3U+ygGUXxmd5XUzrfTgMSWEI1drcr7NVihZsnsBn3upWjQaje/IcC1wL
w2e9+Gy5BgxKt8zvp9Jyvy45znU/m6OhHvV68NXGSE0NpPjYi1rLpD1RXYcaegQz
1rsnred+PPgiy4lDpOecN4wuh6e8k45ySYcWjEEQymMoK8rG425hUkOmdV+KyZhT
Svefwgstr5eptewB8Ryfs18Szijr1hajp1N61SpKBr8H7CInfayPQF8a57PupEMq
UvyQ3LAt/PWJsCwSmcLiEu81nqtBFw8quwtjJBqhQ16ku3sNuMDFDw6r/xKF5vHj
tygrZn63Zg3t89gnj8xqice38uNzipDhA3vMjdtEf/8dxYjJZeGU6nriUyV0IjoI
fTD7uX8GyXbFO8T3nkkHeZlkjaUZ79hkAV3mN7LRARqic6Bp3cW3ZfMtOQ2iuJFl
LuIA9iigmdBPy7OYuYyLuz1D6Jf7C4PpdEp4Rk7s0+pQSUd0ebz8f0oJphkBnuN8
arxVtNOLhRoa/pX3FpBZ7pIpOwGq/HUOt7xCEadNbDpHgeUF5SCdpsJnMAs2nGs5
9mJUIVhjstouoHOqnLPCIRgMmKXVtsK3FLRuz5+FRquJSFjzMP7aDl6QEWfmhoxK
ql5dxi3D2ZUJz412DAWUprOPBETIl5RD3usje+KDlqU6h6dvt3Y8SC8mQn34c8GR
ncDtRExfS6VYV/27SO4az8EkAuvZDgi+n5NYGmTaOXoWZA7WjNwYsqzQO1fqCXxU
Y6SGo1jkXEHeaOsWUt4NHP/y5Imarh/BYpB9xyz9l9tXHyXMLv22K1VgDPP0wQt7
AonPwFQDcnKeAy9RoF9PFg2n6UZ8eQDKXTUKulfdBpj8f2QmNZV0yq6++X2Ic7EX
mhAuljRg+ti3uN+i3h+IHLJhwfZKVQiuOSQTQLi711Q5b2o2tRbASyonSLAMOtxO
rSw8B6jTzkhOCOuu5AjmYHmw6nGvlCfzlSGq9XYE68CRt3cwufiglBA7QuWvF14i
0GG3OMJIrnom6cPtqF3jyAurZoVwUK5Lbf2UcH7+axu+uoi6ExODggjsDBHYROu1
BVCc0gpL6+y6Ci54Ra9RQ76kDPy/P7bIq0+NcurMKl7jW1XTX0SuafH8p9o6YEd3
NWbR89MpsNHl1uB0xqgyhC29cUkwEQ6jvH5kZh9popdJe+h1+CDS2N/ZeNahQyzm
15KcHFoAj31HSfNaXGQ0e2SOdcXOoIoURo+QnFNVR6GN1KEXZRDIeCv0MYXpVEsl
0cx/nzC5o5/YzbVd+DOv48aXIQ+ndgLnksmp2J8J54UYgesP+aQqVg5xRaCpTkZE
8SG2BCYwkrvbu9XCgs/uywd86PMfLqbM6sVlOIocuoRIW6oxP+Mz+q4IJ/gVqEQn
pKlbIuclJ9i/c75WqkzB2AjdTE+DmiHlJO5YJag0kwJgLvwHhuOn/Dhj1zSKRXBe
UnwAcXJ6kU+MpfXt3EfEOIfFDFqlHOvaSs9X2VAUuxvlmf+KNyh1G6w6F5u3eTwe
3UXmDm2jb+GPA/FJB0y/p4dvyWt7+4TSmBqtR4FvMVLmth6jIke5Z8IeF1hwxWID
0Yt2tRR7p7uyuxGtxHqZ8lup14T8DFdKya0xirhwANIgx15EtL1P81v5+d8aOxfs
HLQGjaQ2XHjoWjxU+gShtE5TXI99JBbGxz2Es8I7Ur+IMdLtvPv31FHizKm7M1uX
25PRGrFHiGsDOJ6TeQtL7JT+9fLeJjlSCY0cB1TdVVADOBctNDmhwfCO7XiP1sSu
s/CfyICXqJhZ/Ir5cTJQbhNqmwUuHs3XAsJO4bTXfGcWqL/ebhTcLSdbaK2C5q/h
h5XsdA5a7lgo+rAJ0NK1ALK05gVQds029dJOmsLrARcpAV4quL+bDL2xnWyA7iHB
/0plZMZ1EM24e5FkrpJXw/nhvA2CjGolZe61++pfTZxAP0/S4fnhpTtsxri5wf6T
W37GhGM2BYPhmer0RN6Q45kyCOlt9/1I3nCXh5GBcZ4W8fTWMCNrFrkPCxhhPGHf
uDW1DBf4M0paCgvk3fXuOF4LMikzOiZFJXjDcZ42jTL3KEtPgeNVJIRlbtgurHE9
9JhBFwnm69IktJyZfva8pZ9J2T1FkhPplOlbRi8fAWhYu+vP0VaCkP0VinJla8OG
w6JwXVR2Pmo/Dh1juCYXR3HTBXTduUYG1tltf9h7rF8xaXxKHR+I1cn7sKj9gBXx
2fkS7/tdaj90si+PTVw6qgjHLGyvpXim4T4qr1Em774SKHtvmqLxXOv1PWmLG0FR
nWLOCiJi0x1LSIZabnHSfrIKgTRHKkHKWkRbBP+d9Kg3GI2rlXrxvkSk5h+tcmxx
hozRDSlYUz2z3FXU3AhMfimKqmFXXyWAeGVv2l1C5lhCOrP5VeiiWmfJDeUw7NmY
0FKeY4izVkApPPTmnI2MDd5gX09Wg0m/BwKpXcVkYyeFeaObe4q0pegEpa6Ogxmy
exeTjGHd5uaXVF7Py0E+N0q5LHRjx2qDbeoCD1368XeIPEuiTwZlOWnH6Pxt8vUh
zPeEq6zOKTFfQ/ozuL15FFW647EcKGR224ZhGn2JKCrCLtkgxp637hT/gDfZrcvx
WWkGk9MT4r1R3N5Gtfept6hETYsOtoNZhU/0/iSOU9NN+s2tU138JJJ7ZYOJ9L6Q
qswwvMjwiMQjgLUG25XvU9qe453ny0a4bRcvEpgfQt5K3gX+6WBoxUIOUW4YTO/4
nZptW+ji/v9Ij6RJ+5pVV97tOd6ap/bDpqqyzNYTG+s0uONBFN7twJiwTQx79J/e
DWxYlOK2nsGAhlEkB/kZdfa2bERqt2e7dqTugjz5cl7yfBy2NA1WBZbczwAE47nI
/OWMEDdTrVXa0Rpd2mEG4vGQFaedcE8ScrfwlaF4aJ9oNtNItmIVRkloRswCzO2b
ZeJkV0myjpMHsRv/1tLQ6bsaGm51Ftkt3cix5cJVcYxvZS5u9BDzWIlxv4UP+Hsl
OLkAPEDUCpN8oTNhZ/mBPGKlCHmvRQwUFhsckXdxeMlZMrkyX2aiSR9tpif/DuD8
sY7/KQ6ax4pkugAZPrVkYYqf5tpxY7wb3PTzb7UqEUsTr0oueXeAeAOBs5DvvIT/
zE0yXhdJmKSJcx7YZu/9A5JLqrR+fs1BWd991c/M6SbSKnhyO0L07P3a8zhEOraj
KdkiSy69WeZOb2Qc501lsjIVTGKaIWMoiw1uxqiVW7ie6tZgPpT6hDDhOsuqFRZX
GR7xOjZsECA2S8bYsUgZEwyC4m2F6zJJvKV4l3ZB2lBWBRXXIYS6mL2YHLBagy+d
0QMIvrLr2+0oGhL8xe2kHn7E+w8LaSmsEHO0pPcbg3itJqFJaLxVrIxV1DkdsiHF
W/0Rbkr3aYezCu1FCJEOSGOnZ0F6zdvZSGJR0uOuOonL0RvTQ7cug5GWlHY68Mep
xb2ZjPlV/2BW+ZJxPcWIaF+9lLNcOqeE4T7Hb0FTsVNkXWahLGB4fLufol7+gDNQ
N6BgYvoISP6Y/kIXuFY8+54rImAeOGHjwbCqpL76vX0tXazJIHFESmF33wOoSNLp
zO6vItHOphFiDVQf4d8dvnG79TbkXGIVo9QdKb2A3pBnHI5t7Gsy5rLSWGBbI+UT
YWP+JFE0u1ga0g3zbt5Ik4jm0y0bHLZkGssFdPnx5Ata/1Uhr1gxjO7JanZtOv7t
Kpe7OcHoLVEYOjp/LftjAQWLK1RXiY/TMkF+lCIZNDzL8Q1RyVKPfiO71wT/Sec6
hjMiIY0exzLm2/r+8SpqdLP/uVWK/P2BxxYCC8rrL+N+q7RyfP30uwureg3xG0JB
4ia+F6rQTUiRIhBHYX03Agq74nA6JPXwD5+wwthiue8YWU0G7VElBgWIHXikGeqh
2UdDO51Zr9T3agJeCRlF1GG01L54muvhSUgWEMmN73pK5HqVwMzFDE8reHdL5Hb0
vKq0iLfu2m5tRpjw++kjvvHQ0D0PLeGLSknIdEe31rkC0J0f5DTFpUO9H0/5cqVp
3AYlDpgYS31y5NVfqYY4DuKsq9Pm12TehFx5eEAYT9JP/vRx+5Io8iezhyCJ486E
T1hNJ97jZemiMyr/U3WusnWpg7OSTEhXLBn7y4NTu+Pm6NCEGgavLaf4UI9ILuGk
+RReKIZ64GApQx3SpkRH1cG+dRL1G8XIouqKgRIg4iHzxc54vT3O6XjNLOk5g1Zk
D/GaCnMWTvgWnsvLRUP3WvmFDBogCorpjxsXePqE+1lE34UOABz68TOfwSFANNlb
bvtnZljW1TXrwEQRs1FKT6FH/PP0SEN9wSkTquwvgOMs4mDJ05T3e3KNzPZvin7C
R72g8/aVFhSDc0oIDS7KzJwH62xqpQlaMcqMbsnzjoH7EuAvJUHYTqzD6M740Rjq
LCIWO1k8jTnahncfMJObxyU+YCHtBiP2Ep80DJsGnR1aSMjk2GDs7fZjAPnrq7Xs
4n63iLoKdyeA6867/RduXpEB4xoofLJoUQxWRTJV/N3/aU3C6UH8j5tCjVxHqDxj
qYHQz9C2opbSOzxMJlUP7Aie7iGhCBMWI8PwHkL9P4zN/xK2KyJuRAgqlUnWMXbx
nitjckoxn4kZENqDdc59E7tNsEoEUGMJPX+HLNx3Zrn7kiKmqT8kPvbdr/reOyAH
rrCYtf1E5OUQOah+Fb9K3Rz8h6MqeeoRwO4rU+Q3/DWgS2DUIPNwbm7Gc80J21XO
xV81SMIAbxQvPZYqGSopPKdSH4+SYICTv5ZV7Gmv//HfYvWl+knRjadLxoLT7qcv
+fltxAYe1jZNLj5QR0+NYsrdoNjdd3qLqgUJY1lkQpPiPnqeDT7FVIuSY/RU8YJt
NOBaQS+z/v7q7jJ1P6cJxzev2cHJe9n3isxmJ95RRaEl+9tcy7vSr2CaSoXOG18B
/o/VsJXZrPdT2D2I+7d2hR0E28NOT3J6NGhxLm3L82xG50SXBOEcK9OJNC+GsrmR
MxUFsxj7unvwtdvUBuD22joXeo4OHQu46PF+2fZr57uU4C8ETkP0Y79HlhEjpZ8k
jbkC0HzS7wrLZNrj8AqK0+iZz9vmvzVlLZlC3TLpcOUvUFeojW8hyCW+JGqhEDA3
sAJJz4l7yrAtNvEfu8KGNg76uKXyjrDS4woklojdu+f0bR7w6W0mP6xuzQfwd49k
vJI2LD0aARxzuDPZX75HkY+fO5Xocu7sQVuOsPnVBAz9y1cw5W1hgDP5p74DXqfx
tO4Sh7G3fOo7YSaFP+6IeLm8/bvqqNtCgmfpO618GvHj2Oydapmeu+JwylCrL5k8
5du59N3X2+AnF22lYQ2ccZCPwBvLtFilj/mJPMcOQwQZFcJo8BJaVLZjCgfNEJmJ
boOGEkoG5cJI+JS8CsIHD86V1U/QN+1o0lEqa/imAgNXe64Zm5celNxhDobn9CC0
+sZFXhuVJ1jczzy/MKVx8ShGXwTRTicXyPUqrEa8HKda+cQrGuzhyR3w5tMeTUwX
eGn+2OY2GSFe8GxH9lsLlB8VXNudEpZzWUVRAIu42P8azYKVOdWc9RNbNU6PIAgz
RoojpYdCAif0B77/QgtXyikoX/mCRR/HvdBuPwDixHGCTEPR/eyeGMbXNu7ufnx+
hrIhsQ+ep0pgDlnKONx7QS7cFGAS+2tBXvgADQtrwbmMZAPVIbti17TDWVYJjnlH
X9tajI0eu5UbjBGjAvuM05IpuYRQV5qIn1dVDV4bE6O2+JYAxfizeclS4FzwQyzw
lr+DhCKGP1NGnUeL8ecMKK7TQso6rhs4hGZHFvGY4N2ferjLvmLWqjx0WlE+3Cge
G3fflyY6/CM6No1JTP70uBeCqZkehR0sWQF5dIagZcIIq1VBMGjLarrWVtxAwjMQ
hxWk7uDZNNgO7n2qJfuovlFx9lG8rJ16vH8TbMEGRVg+IaHRSL3ZCDGkZ0FmgTgO
Vqb19DGr33nKN/hXUBp5pmfqfvHMtgcE63znVAp7rBWG0LLx+jWXApy/2Mvd9Qan
P+4jAHezkmjfW0KFdYmodcdVXwKmdPk5bQF3U2z3GsRrLu/lKIFyjq9nb0Fseebw
VpdVaWED4ME2+K7ea95PAd1AIpNSN5W+Y675DvfO1YTijZrNBj1+YDg+20L7M9AM
Vctc6GD57RJ7wF83i+IFqMDkUaDPNmac1LLpnWTHELMmFWYQxcikINmzi2RDUbgw
nfIaIngZQeX4G8yWNm7BWZ+1jNCCv6CyiM+9UruHqkEPspAGBdV1Z//wY7SRsSJt
RzEj+Tgh6iWlkJAqjGYIabpIa+qR1IxIYFoDiSvVS3+QPO5Ljb5RIOilHMW3ZvRh
NXo+2us9NSrV5DrYb3RjEJjo4zWEAE3lWk8iCgn6k5FmYZASCsyrXYHLqn0zwayX
adx0rcKZu1NLir1git6Xbz/NhdTzyHJeDKxvfM2NYoxzGgapAgGXP2Y3/K9Ukhuh
fJqq8L+SQHVKZXPhqtk+BGoYCfX7/FAvV6gVOHnRZA5ocstPmAzOkxjOGJIX/ctx
YgqmpLnitVHVWdPBed9VVv3y6Q1qFXCa6fZRJK7WARsySZ3nJ/G4Y7D5B70xfpjD
30dU4Rw1a9rF5+GQRIrzw68b7VNJYY7rgZwq67ZSBORbuNGikOlOHd2n0x10WgtE
uhJ1cHUZSZcb4jeOXrvr9rFXq9dYqqG3B5D6q9MMaiS45BGdDD79t/IBCpHInG3+
eB+DEXPjG+g+DvLQ4BukJH3Z/mxoKhJq5DW0R2idNL+ogXSYhyZ75UYslJzzK0o1
uY5i/iiWGU4woj59m15dXBA3aEN2jxBM2w0doyWaZ99ZN45rZ6B54d05FcT22JGa
yeXT8v0SEY2SzEl88CM42cYgi+GV6xpj/pAzkMQ2jN5eMKO7tJA4XQmawE90p+RR
7YUHF+WhoP+hdGEH0jDdHfCBlmNAwVTvn+Mf8E11/98H60Y0NSTSGutc+5STWOQM
8pIUow1nOFSafRLCWOJ2s1dG+0cswIGaNrxU+X4knCdgdxcD5fkwSu2L4nacQtLu
X2F096Yek2BIEoL1ZCW+toiKpMzNBxs+O3SXIId5mIY5p/VvdeqGht+/nhBIqITR
4442hW76YBiad5fDFlVRmMjy0eiOid8IPDL1635Y1fYWRRPMuCYuyD0rtYad0nqf
A0E96K6+R+AtKyGbyaJx59l4GzGHY/6IyfWQDFmo3p5sL8DUFS6tpJau89Flo72W
1qQA+3UgPILVqsv3rUdiDr0wN96kV8T+4BrSRgHiMno7qan5DuaG59g8OnpBBOgq
mO8wtYTw41zF5QfdtK2Gdt+VVZmt07xE6NkvPCSE4At9IVOSxgAxBrUswijaqM42
AaxEmGzw4vniOENMcCJnvu1FcXznebl8YkIe2agvyrBkVYf0SIdXhz0okq+g6C8F
5Mp5b4ciOWdszpunVfMbNSiScGwnBackedHX0gPefu+aNCYEKftXNmr0B1g3MWK2
xvRBKz+0uKv/D1GhcFEv3jOj5Tq6CWT+sr7Mub4cSyIwQLR5iDqW43/UH3j1+ghv
jywQyNdIzPNTLJ4R7fihjlFqlKkm0wi+myHC/0mMm8ItYioaBQYMDhxfLBE6vV/9
DHLLHEa+7CzKXHePp3mIWyveWjRXpDL7jbSfHNbDW0G56RvQMApu6ylV6OBqhO1I
nL5ws0SU4jzJIMe9rTKVUUh28X/h2n4hMUouRBpElzCcIge7WFgAGTcu7sOYfpDx
gpvqZEhpE8+Gyiy6Vr2JK5EFPCEtRwrFaMCF2UpHo6Iw498A24NuMhYcFd5ok4Ha
Vjdxs6qG7nXjmn+z4NykLs5p27/34XpWA88wSG+QzM0uzoTH3JhFuHSHmpPyujAR
JDL8oXdDJdQt86GiNyWq7SyTLz3tCMF2gvm6906fNQ7bmoNyUt/VhRvotQksJdfj
j97BcwRM6Ow1pjphgDyCumkvBQC89xnHlI/Q0fNxJrT3fwYwwSVKt//wtaQgI+ww
KCo0BmIvmFCpVNk7zSnDcMV79rEBsC42YMcrjGrV81wa+8jH/vNsBDTuElcUxrG3
N29+p1CP73NU/ZfWszh7IMsX9Cf/ypomULn1W6Yzla1ejBQm0PGZXEnk8uXOKbhB
rZdA+frFwPR/oEQfNXye9Qsj4xlVlnPgn8t9NI1fktGGvw20NxH6rrI8JVZPUEE/
/37dBybfrZeiqBCe6Feu7R9m2fajitALxDfnFbUgm1BN0SrGjIoU/78uG/ajL3Mk
uvF+4VM7EKkQtY5bv1Rfz547FKRRPvHsdqZlglwfFiAhtqvIKe0qJAP4S+qdUDEb
kxLm2Mdo/5bFfaG/CdJ/14NJm4xE7Y8lLw1xL6lvdGgqp4LtuaSenrVnW2F75jhS
bJ3T73mATqSB3SXPjJsU+B+BDCiYE3G6uS6VC99lkMrP2z4xIAWo8VK7mrRlarpQ
spaXDHhIVso30y0jYFXATV9JxBYGPvlpgzgVB1fb83X8kLr26+vti0x0eijSOxpA
IBtIni0zb5YGvgVzGs0b8y3HN83EbN5MZWUmYbDpujsiRsg00AaoP50WuFo8au8i
DVTLUQoBCCv7sSFlNDZmKT/scKnq0VECLM4sr6jw/A3UdOJDZZnsUFNW8gyW2+7i
3mB8YPuSMGhjwEfi9poyyp5GoMnIoshrRDCJYUcEoNMBlQsKoeyatXf0lkhDTUzs
Ia87daPAzUbw2PZoKHJrIr3BemBdoCFM+WCym4fgKp2EtACkHMFe+l/zZc+I50of
Y1BB0EuKLi3+kPoqFXZeVIliN+B2VA7PQh7UTlMCgPxXLa8xZm2vTuDCA1+wKpML
zkANF9+t5HknOcvz6SznybZEtekTKFWuuMtlhMaKo+7L+Yilnihk8KGF0/glx3HJ
9qKrcJd2KmmR5dnjaLDeePIcvP/T8gikRABwf9I1GheXf9F7SG4Cx205nPYaYdxB
ZKdaKuuyq0QbBteQjYmL80ZzNEHjuUzGj5m3SEGQmq9xzHXoMptOnvqUN63PRano
B4WpMIAAo2/QOpqRuD6BMjkWVmLw+GPITpLgLAW3qABhkJ3zv160Ny733tuHBWyq
o0b6tfSe9t6RLlW9PTEfGHqT/neUWC5AqPRUlqgRuCroXZOXSXeMTuf16a1CDRkj
IyYSmpHvB8Mn07pHI6ROVcKMOguS4d+F+0E7DOpz9c97a6w74y40Nz6hQ8/doytZ
+kSp3XGkgAJ+LJ203kNT94I9865UJC+89/lSd2JJMpv6aM+mpiTEpnasJtV7z1MI
cRlNnElB06Knh9SmUMpxPP843lP3gCzY1GLjlZKw+Xo6tIcXp8IJfe546oCvXFHX
0U2dD1pM4EECrlupDi+AODU7VC9ixi182/YRbZgFGG61rSQ2DMArEii5xjPheY7U
RizpndTRAMrekbVw8BYp8ysgp+quzKHHc5fWP2HdzNjwXWKB8FhZ/4KI5GX25AlQ
URNpzhhhs0rVdKpvv6QKC51za/OYUB8nPDgfEU5VWT3e9sWtVkXpwrPDJr8WR9tc
Csb4Mvt2Y7Pi8TAU50cefnlcfZv7bcaTCNA80F38GnLz9eYqaPdsNVFv57ww19oD
dG/we0oewnuvd8OGnwX+9AouzVtfStsDxksedbjkH84oBlShO+GLcftNH+TuBMa0
U0uTOEFZjyM125jbJ5e78gTYQe2xKPF4NLgf3EtqPEqFsy/v+VCVAA3olTq5W/C1
hxcuN1fjyWcLo+MsbpvZ8f3UzoyM6XmslPNSRYFNXF9vzf7Rk1ezBJR6Tj1gHRTv
R5rvzOA/6CW+lFWoGz2uM/O35bcfQcwww7jfxtcCCJ7dfl+OSGWKhFLxuXjOu5+F
HVYu2w5a83mzClpvvIQovW6kY9YavkLedtlBuDaT6bqAv08TsO3hCt3E/wA8vWYN
CIvvXfAyJPbsYoXD/LffwYc2PeRmQj3ygoI1OKfqNG3b/Xwb5/Ct7LARxtPCODeI
mPSO9FqCjikPRLn4Fw8E/KHl1LuCpVzF2WVTzGNaHao1mwF8F43d/5OQQ0YELwS0
jRFWyWDWFdaoYj9zqxvvSFlpkBotDn0AKnUSMBAveaJJzzgf7KsPkWYNlh/MSTI+
1UjUTUO/iNbaG5gIbVP9DBIgxGYcZSb3T8pcGLSYxCDX/M0OjU+h/3QehHuQDB3O
qeGjBtZUWoPpwrNhrpVZcXZzX8RwpDWyi/qCBZd3EJC5Ay28EUjjZJAd5KXjCFzP
eCZWvyk1xJaGHbUOvr4xdtzOPE2694J/M8xhnDHU0Is920LIa27M1x8pzQKZ2pFv
3wtlgxfIf7p0Q7IbwL1NNtY+TLufCQm0TDBX4XyVzVH0AqrDXY8Yr1H62nxgkvvv
zT+jSwJlCAaEDWEkbniqN+Tvq14Od2GxLDECxt3duJviFOUGxcjCrIJpy2KhQ6wP
hQiG7BMkcN7ppiJnpMzA89Skhu9ruvHtl8qBx2ew4xFiAtKzZDuaxYF5vPEzCkv1
iOGEsnLIWZfVzRSWAt/l6YHr2qTsr5v0OGX8AEuuBQyV45Quz6pJl6L2/PrUm/Rv
ukFcFtrMBbpz0HhYXyWAEjj6SMgnifXj1W3FB7s7IjQITsvBiloxkYBAbOPB4YpW
bt6gIp/Gk4QXWhf+HacTOQA6K4UTUGW57yJ+jYbrV0ylnoOhGxUQmmjI6APPQ9Bf
dnq0hzfMteD1tu4QcY9goNzxMJMQToD4r3GovOgiWyxrkRbrRfnE66BnqGyQKBn/
ciNAppGmI4hbsDVRvJPUELRMuj85L2sPU+vEWGOvzwE4XO3YRa/piGqAQXuM5b25
nJYPGqreST6rGgSQ4Er90uzYDAv+YNqj86DDtEAWAlUF4MwfRqo84Rf5K3aSdgS6
o+28lT1C0OPSaqnUXnCn5musQpsT+HcHsLi2Nax5i3Y8ZH/T98WbxeqbA5Mqo8CD
pjJz9UYThI60B+KCe+5LiLF/kR9a2C2adcEigOGbyVS69JEIzIv0uc96P2oJ8wef
PPH6cxKJpbb53DhnmrhiEFLjBXSWW7Qt16ZTK22NjRjRfIzFlfTkB58M+i0a2TSG
0veQWQ/HtsPHFyktqdrbM9DfNYrHBf+unWuzga4ETOhPJD6DlcGuA8JJPtHk/ztK
FRYVW161/j6P+tUIk00kcDBWyHzpxjwy5z7WeFHZsyGARGYTMu1seqbj7Ct7i/GO
o+Ff5plt5r3AbtI5EussuCLwDIVpXxLZrc5h/aTazyDW9k1UKoSD+LQPjuKFeyPO
ITZHHK0Jzf6xhZ71BUK3BHleI1s/PLQmoY3gMZMgWs+h013rpbymjIzAznwP74BG
u9tcKKprzJ8QVAR9Qcx4vvtlqmHFCk36/YXFmU4EqjyWcVX63P7yy5J+W/Cm9F0P
LpICJDr6qNkHNr1Wn0+15fSC+bGP9X6nwTqjlYr/6L941LgK6yVFt/JieyeRcNsC
zIZMxbZW+STQ8ZgszMHoqxeMRnXdXLSgh2HZnD25ihqJXIU6f9yqxF2AxMLPvoiS
8xs5nOc7YQ2o3x9w2kqy0aWfp3IexL//KLCmOXDaydLcMRf19+W8+PC7hTxcNSnF
JICqejkDWWLR51z5gwtyuG9BDLwFrTWV58lyZ8s4Nh3m5KB24tQVxPi4CgZAsJF2
PDZQG6Z9OyTFDezL1nyFp4r2dRYYuuX6MknzeUtlY0hU7eAot19pySwx3j9ZBa38
zn547+h/Lz3Sb8LlB7pBE6Nx6DCYZ0658QBjhZtxh/bhDeMN257/ztCWv2c1UiNO
7rM/ml86PmBIaaqVEcDiF/VR1OcwWq/V5se0cMC/GQsKwBAWr3CB3KDsnS2XlPrR
VrSqFMdnIgZNN6R59x2n2KIEDm8A4wOrerQ7RR272UC3Cuf0mAWHxeQeUR8pZgkd
2yeA0rmnjTivpNYacwGVvqW+Ar/jB+qs8A1Nsus/aBMKapcszjfcUipo86mwkLRN
siM08TgFf50J5Lo3EUYlmd3a0An6cKPiX/CxPLTvgTtivo9Qgi9oYgNn50O72lym
6cl/7m2vXpcrrZYpC69eI0jAy2LA0oESQrgYiAmtJ2dCAWGQMcM4+hfzaQXFlUj1
K5wB3q6IuCtEGX8AUwBMC/Tnoqq72gClrHk/rjNBV9jyYBGwq8vPHyjduC+0hRhu
Cl+AlMJdtRNkvdjDMHvJmCdVQcQx83X2WqHyu1w6UGB5Pqk1eXLdgQuzi9RAgMw7
qyQg8FciO/hjtdq4W9yATLAdeRpAMEmvUwnde3an7yj9zPsBAarYJyGzvjJNzmXm
mJEBvks6Z5pbj8TOKmreZz+nvNKE9Rxwj2+KbtCn0N+4o4Hl52drUZxaSMtnjmNj
xa0lWvCFwXLJ58RVnU5lQOSop03WFyOMXhNC3lfuWs9DBX+868/o4SeA3AURkrvY
DaFM9TLN7HJ0eB7l78aXhD+IXYbARMrgcbQn3RTefnPqGr+w3xqRoZHnPm8LcWT7
dzaJSlGrSFGRh8W88kwVoYcRFeGnpzO8pf8o0Zl57x/tGzZb3DFcvwgeCn1gC3aj
/6pBhtdD86Mh4+zXn6b+OjZO1YtA7iXM7EXr7p5VvSrNKoPlkxXwP6CbFgVALZqV
FU7iPuhheGlpQUvI+0oiC0jP4sHgBJfAnNMRf976Spsif225OwptPw08D56pmuTl
psL2F6UP2LAlZJYvHTRZcqfhrDBHlTP78Yp0cZAsX8ieblsGu7Q7C0UJ+DzdDxWG
ctGl3ligSjUb6ryzkj3jr1qcIVXwEPObxEl56asnINxPyHDfccB/lfd8mDrt6Y3h
9xkX5tkscUbO73t2BxBO0iZ1dZQy49cib1ms5YpZsgkJja/AajG7pCj/2iuhS/Pv
vSOldPNpwQYCfLObCkuSwVFGytB7xGhNzGUSQRscjT5hpC/4S8IQpLifhCHh3k67
ca53aCy3/ia3P88iLWXy6iop1Cn6oa4E0Ai4+vGd4+JHu/I35YGtjddZ8w/q7IXM
QhG6VZneOeWoXkRlwREk14jDQ85qcyE+3SBL21S7Z/me7McR3SN7F7q5GbGN3e4j
891TrPf0tJVVRZt0Dku8U+lqqFc9XS7hZhxgk/acUFxqNs4OgFyZ2kjrWq0hJiud
G3/tagSr+TS/kh2nFmNLu8QDK1MkMjCWRoo+DCSLke2PNO32Mp1mDfvHHIYeBtop
SK0NSZJmt2BU3MZM1Hyo4mgOXtXlyPQ9U68ZNGSJN+RGFbtuo9bD/jCMO+J1kjr0
VcIA82xJlo7Xux9vO6ZCVu8T19RPUIKeP2ZI6KOsqhs2hSroV1IqkbDs3RoJINtg
x8i5a+sQlSXEyk+W/CpR3d5MnVucmwMMxzz3BB1w+TypXMMCdUk/KttJPXIJZCsk
sG4zNOdSUfko7gT8vYNPMJUvQplo2igSzgQPjLuG/Vjvo74V9gLPRtkA74IAwekV
F3tyq/ep55lG21zi7BAkgb0E9MhBeCixeso90JkkS/FuT9gogA8yPrHI0P7IJDzV
mXC2VRrdmSKfmX/mKWk8A6vcaKSEXfUUtOoc07S39CfKCqYio/we7QddFiJLGep5
IWapqjeUbKZM+nmeDpRJp9ert0IRnUFPUn/pG6pnDIVWxJFUcz8fLZF4L9fEUEqa
mTyja9/DxfPpzF+IK6fUlRx6hYUIgoY90Lau64V+d1X2sKZxVxq6ffHjnKR8qDJz
dXbk+yioNX2vsuu19oCuvgjDoaVRzEHsVc/3yYCNZKpQ+Cby8OuG2WB9vp6P2Opw
A25odkOWNXnSGGm85cZlh7vXoJ6kxlYPX1iTGHADWSAwQm91QKVnZN2f/b42rTo/
OCIXU5UMVlPON5PyLS/+cOgyISBatrnv1Yo7tAcodiXDPxbdvua5a3hFJ0L+lqH1
n+gl6ae60JiDimygofddMdiVt6knRxleFA8C39jRWxeUhTAjnJN5oE2gt1sR7/dy
78SREVnxxcf8nsn1erz9igeTh9k6iBIktUOShN52rLQahjeih+G8k1pD/toTikVv
ZA1qdSKDk0+0SyxdBWSGdwBYqVgLnf3bqxdsSvsguuAPMgloWKmhOOfY7DCLe83P
zFFPr7GPsUkxK3ttEljswN8GhXCZQQWqhb4lJGWs3YQhdCrneOVhRwUmeZMRiYtc
rzJ8VsI+83xH36qpRM3A1iE/4K/WaC/r+UN5X7hsWpcRa7pJ6X5YRUKsBdjcO/99
M0lcuzhWIW44fJ+Jptm1lfoDYntHaXXQ+Yc3bjWwkqhS4luL0vyuCI5G6hNgsn8S
1EHD3bWaDQ348s5aZhCKwpWTveqiR2qW1dPloa/E7Qs0STPf5j+YvFG6Nd87pEKm
5Zxz3+BLcR1D6iRLAY8gU0CvybWafrE/R23wOib5gIbMmlrVXvpGpFKt9hveOw7s
vu3ncvIctbC9QksxbI4JIsH3Ife/VwEITUsphdvVhlvtjBPh/tyqTH28OEtTJmhS
qVJdsgdrgewfU+DJbrBk3vVVcuR2du7j/u6wTWbDVlmRvWwpt7oMQO56OhcM+XLJ
t/Z71As2XvjeATFZzaMNuWRYm1NxBzNtKYGnq0W4jcDh8+jZLuVPAj9r30mKmNCW
3LQhUZRv2BgsdNW8GEQlZAndjqtHdGeVHiwmDmsWYTtF2sr8UUpNrEJxEaq2dy/i
8g49bfRsf45+Wh2AyliXmwiadBNXxSlJeJ9OsmE4fnr7pLVYHhJpjtE2xcTyKCFs
fUCYlheKq6iVbO2ckg0jerop012+9USRLEzswhsozfkTYMC676/3yWrdp55U9yKp
bIkkmmvA969yK8bEumkwDsi3tVLP5eIONhe36Hz38gkXZ32VInzPL/gLHIgAaZE7
QZKeMe9EFgEIivt1KvjexMDJtCnmc61PS9tF8H5jVwVo5abJel+Hn3qVwPSSQzCA
I8L/dMLq+3elFmsjjWyd1kGtkRBCTBxMr8D/JYyHDs0a4Jc+aw7eBOR812+gt4hd
BockRDZrPtV4XjfzKGewNB0Mi9mgW/R3c3sdcP0NctUSOzMXLBMUKWTuojJvmiF8
p9ehOSjNmcuqTl44AHUddSbyp/6iwBDRHf572I/GfFfcxrO8js0+aWKpmoD/kAIR
KW8ekXo6J+1WzMQu1ROsygrVeJSNmLryGTp3s3p4cCr6nNQaGOPyIB85uopex6IE
j3yyl8ZE6+2pBNtTTDzQljpDTvSwoqT2tKH0gcnppkjePjHmzdAIlFCIYvfLXFuA
1e45GwJAu5MGRH2kzLtEDTQ/UTtw3HJQ9msYkyftXe/upzaSBrd/j5XIg5Jsp+Rb
DP4oi1j8M1itcdsb02cvrTyRhTFCr47oozeJfvhlFlWlyLsa5CIuYq9vzBPAIH21
YmBYFL7QdrHTMhRv5sCWlIWwlZLGSTKLAxfbGpSJ5eQyeeBmTbdbATVRLnpdwpr2
i+xxOeIJdO9DWTkIFvW7jaHOI78z4pgrBHr7miWiHku50SkM7zHJx1Gav/lb1cyA
a57a0jy0U13s6DZXig7zdPZJo4bVB54RF9xMe+VAhbYjKvBtifobOQXVwjw3g4vJ
P5+6O6RVX62dJYWLBKjSHriUZWxWkUDeTIXzO4b3DPpUT9NhVnTlmGnQOLOxO00A
6RLRgBfn8wxJr9YFXAV++qx6htKzIIBDAcIhBn406SXq/w1HqMc95O43TlZQqKJB
05YroxVGWCOzpMGltycrelPDHX+MHCoKetXkOFIroVkg+9LipuE2Q/yT1hTN34Na
hLV6tkC/Q9SZIzpV/tdzf2i2slWKIHzLLzIPuL8ycxGOHyRFD0H568gBwkhWj/gN
Nd/WLk9K/NeL6bSV81NaIM/dJRRaTNjseR3Oz+K71IqTG9SLM95yW6JRAoW1CRYm
oSBmvUdLDxpsO43eYZ2y8DMhQH4GJ4wJALtd128dCVbewfr8kGErnE5RUr23/hxD
9CkoOonoTqS2uqA4HwVDMdR+qLcnlj4LN4xnMT0tnubILN1r7dFS6FuuuLTUWM3L
sF2l56L40tkRb82AJ01FFQ9hYfmBKfRtf5coFQslydmuBQjRhipVQ86bJ6GJOJIy
Z8AYNrM+WjAGq9zv/WomGqk0YBbxsRAiMM7FWH0n++HXekPNDUh5o/k5t2ItJTl8
GVkU1w5u7TTMBm7GiVAUQG7vwBLGtER+q8ftQI11XClNtNR9SgHY1OBkLJiUXf4b
8rTbgFAFikedKo7S67nofkjbGIXq4f2hRv6qurQOSjnHwERafC3zIEOjuwsNsI4X
Yqkdizt3WBr5p82FbCkf6NHgJ/RoqbCNs3ay3ab/Lj+GEESCy0SJjYDfC/0MwKyh
7U2hgcZ1iRLZt6pXiB6ZYupF/SsUjTw1MUFcPgyQfW36fPmDKVG/Gok6Qa9JjcD2
KjDj2YX94WCrSh3cS/6lzDXHXAMediTYkUiclysbjlJ4EOVaoqT5gnljmT8DvlKu
rFnEwKS7OZkDM57/R0l/5OieMsbBmX4c5LW5HDMiVlJR3HuhipsjgM3tKXJ6Lwur
fwPdUF+wNReywIGmoue2eeFf9Z/J3+2h6fMx9CwFH8qfpXvq0PIMvXRba8QmgeHg
Io8HaYO7bHuXAaQ+dHHe1KVVi/g9fwAjqThfP2KWPfYzjwULLhPzOWoTC4ebCTBM
iindQiCc6a1rL18YdcPp9gdd3DBorrtvtoV4oEsGp8LOYlrWOHFL8duHVSw9qdns
YQby1qPo6pSQCbIOZbx/1g5m4jfhzCJDx7aBGoN9DjpI0SI/exCuGE9bLd6VwnTu
HAxu9XSwk5kdFAstaZ+SKOpbIJQuZQdVDPk7LfsxajPoqnRkZxmmBzemoMQCN4Jp
7p733qJ/9UpGKMQ7Vn8Ip7cj1U3rQB/nZNHLeJTJXDc1TNbrd5aAt6zmaaBJ7FcD
hBQU7maWCuutmv1AzEBA6jvh+5SK0tcEUfpQQLGfgVc2pziUjDOVhwbyaCeALAKc
EcgfJzfENi20MoNmnTURqL+c21h8rLEzQKdNFQk/hXoxvpGTIgigOz6O6TleOZQ8
EZE5NhITsJC3rFGwo/DKzc+dZ099SanSuvQaih/7KoqRwth5rF0sm20CXQ5mMXUa
zXNDI1ufMTIcUDAKZ41fNBotVCSNVlKznmz0d76UmJ8XB8xKf0xgNqe0U0hPOXQz
urwY8rW6bepnSeyZnK4d6Lq3gplP+eq0V+Na8hdM9KVMQ1v8MKi/DbKKY7QTil5C
7SAGqTaVwk1veNevBXJsKUe2HDPYynodIrWu0snDqdliTwcgHoHZkW46mfYunzdJ
ZfMJYEwIE5RRDaFSg36YZAdzuWT7LON5DIYthka6h0q0mI7pZDT0dMKDoxHIN4p2
SCO0fadj/WiHsnkTPLxqy9i54WGPJm1CspGNXWXx2YWCOUotPmidAZnH/J7ZeVC5
+1D8BtR6GzjHZIF23undjylUx2U/5Z+fXgB+B34+j2SqKbS7yB1oGPD+FwwbpeJy
ZzoMST43Xj2YCQOsH/DZ3H0aoC1plXBIGoqQ97eJL041rful/hohW9gD7JDkIrrk
5fmjO+iuLxSW29JDezP2sZHkpupG7Q1Bj1i7UGRPMazgua3125BwG4jmc3d3cYyp
n5yi19Yxa9b4atEbVnPh19LTQvz3F7SMhmaEpEG13bG0EEvYxRHOI51bYZbpXv80
93afPcA41BggWF4OorVxkD2b/9MVQbIYFanIobCb7IsQ49IAE73UvlKVe1bjOWlM
RggYvQb7GI8WotmnM5Wji/kcNhOrEv/GyYFG/SvuHDqCaCtEqJ/APn1PvlKol3Aa
grP4m9DVQ26KFB8UXD/gJEX7UQx0r3cN38+OYMAp+nLDQPafrCsAORPiXx22dadw
um7SXxuOiAJw2TV01dkWmX3ByxPU9qqz2+Pl7wWDzb6PwuuAWTPnHjE7DB08HYlt
RM4L/l05GImdB/STo2qaq3LoXC9tbdYp6o5WglFbMCBRin0ZoD+1DqX3bWa+x02F
Vd2YQpoqeqN5GIFK2EiOx6MoXwRwTEOBeNxF/4rJ59hrdiB/DbvXRM2hE+kdpiV+
V664M3fIKSoSwajISrQWKyIkkLwh5dVaA/H6vSZ4LeMjXZPFqfwUNOq5y6jPXyC1
l7TedAFLCY5rlgtYQFwgaw4Mky042L8ipPTC6NPX6l/fXLQhpne1EVo0XsAAPhzy
Woyf7iqX6qeLCPxf6WdtiQtg+azPEmF1YOxfZCQYPQvwMTg1xTidm/zWeJNNhEeM
9UxwILpvnCOCfZW2Ue8G0ZthCxPSvQb1eYfR9kKBtx0EBgZs1Y/EUr9BFZwAbFmB
1pMbHVlraD7WtF2gJPDZ5jNA3f0QD/qKG/MUBZhmwphhMppzRu8Ob6rZF0LxXg+s
qlCXY2Xxd88ErjLK+i09lbjfcLtb8bj8ov2/tOOteKLm2VRPYq32S+JdMwPF5kgd
Bm+WhTeF3qa1ED01l385BXM0EqOaNDlcU9gph1ipwyc5IO3cGMh8/yLhm3eaELFi
gv9ynzKe0+HTuIYuSOuptkKWEdRAe7Qo4HmokG/AIbheiSava5KwUjrwb6smIAV8
MU15dJlj5DFyaBoIE4syRT8BBSrqZiesa/t2hID0+Vz1uZHsvuWu7SGjtENn2pJ1
2W57rJt+kvClLF9eHnalUmnP3+E1SL6IpECuYds9JcznZMKjPjJkL7OdVRedhIJH
H/buiCpifts6w8zF6qK09a8PD9iw8Tpuu5J4Ts1zouSjix5o16V5MRPTfpfg4VdM
xL3t2dSorBuOg4TMe5Ao+Q7MraLa/PIWuXkq7+DAD9PmNUrMU8S3ImRYa9GSvQaG
+mmXnlTJ31Z2R4jcx6jKLLJnkUnbr6tRBkT1heu4E2tqpXTiwp69V1icqcqEjiyk
5TDS8fVFYeQ/oJ6PcBL6XEQQwALK0Ca8dx3dOZjKP4NKKVVspk3CKcXd7dd92H/A
cMLuQ4r3x97uAfbmiHIX0W08OPFSZCoosMrPHAXwfQfv7Z14V4RNHHfsrFK7ylO9
zNkPQp9ZWdeihIzUej5ZymEd+P8HFU96pWIPInIfLlO9kUtS0xVeS0Msn51kWL8E
rlH5eEE2CK/CBryTUGsYKxQX+6RoHkuf9jEkieNVXzrvwe5aVrU4n3kA/dQVkk3U
OVVHdb9dIs2mBwQbhgNsaOUeb4hc+d/am5TBqIprZf/pMDk/0/AJePbSgesCsp4T
Gf8ZZ3hqcW7DT0L6GW5inFPR5yIRejKYS73TSfQLZj8t+Z72Q+LUbkVBN+ZSqPQF
/e1SqMo+o09njIRLzak5vCqanepFuolzhDHS6rfu+lkClVNrW7++8r5fX5rO5bL0
3q89ph/D6tvdZtc+WWXDGopoKxkZPVgWIGqI4fltYVoseNDfIpfD5aFNYVdX1hWU
UAKm8IIznU5YW8YmMccd1auxmuFFVQNnl3/enPhDKlVjM6pOFiFA2R0iuOF7TxTI
cxnmLcTQTtyqaWlUgi+Q1K1bTbLVA+xfYC5UiNkYczTFa7ppSIG0IXp+9ljFPZoT
fOCw8eUAhyZhfNiimzIGJ/WvQfpmLEyjALCbboLqpU8vstJVuJ6+L0J2hQ2hYxaQ
08/UqhysR9CjPPPZvS5Lda0n3745vIGZCAEVlGxB8L0Y6fELJzaauI/LlIHbuPjF
LHeBvS6fGiJPURU62ZwOXpbR3kSYVABubFBrtxNmPK7RbhSxuJ/I5zi+AXHxM6ju
e7FRUjjy5vxQvrxByhZz8NqxYk5IdsWsn1kHAaqUUHEnAga8X1BdnceiR0rYbVc1
TlVvlecaWPwRrbDPrsTut1xS/MU/OncLyEDx5FhdxaeLcB4n+uzgQMynpuU2SoUf
f4ZhbZYcUf9enposeEer3xCkIXm2qpWdXPaMAFDZ68u77dxDdkp0AL5M+xzw6bzk
xCDOYJigIXzjTeWb9VgZNHWuJ/mt3Jx2wbY3xMn6J96tIiQfcRxPVHbhZl4EOtli
5Iv2ORWtsmMvJJTwPrZPH7isNnaKkmq+IRqqPqA21YqC+hie/Ig4HC7bQo5hZ+u9
aW5VycAbD0YgpOl0zer5ZJDRM+9fDc5YdRxuSm8weu7fv7pBVTJROJTT9E+K1G4e
cUD0V4Da3JKOF7tLQQ6dXv3i1caH0JcwMEvop2lsPPGn8BTm4enBvwiC7Yo6IUoV
9ydz1wFzNI81DpLLdLqo/VTjZ971rF9Ln/Wcojm5Rok5D8FQZk59NlLvA4uBXb2R
I9YUmh832DPfzqeBbVx3LZVCUk9yBnOGPIi1f/SQPWj93k2821y7gSuRtDAQYTAd
VXGMcgPgpRY/Moa4hY51cFx82q+MaKVmWluVdRyXrFhHiQDf0Oikuvl5WyGJlk0s
6gxSrfP+edwKGHocCEQIBHJ8r+6zSqHirf8sUPqC7isVW7+4DeLEyph7sdnrJh/D
2L93Z3vNvrjvMWAqXBdnX06yKNLrxbe9vMTL6K4ttu9i2uJbbYENXYyikbz6x9L4
z3IJfLtp3LUY2sdSsjmD6r9AR0E6NAf2C9qg42+/wpOnsfFCVxNbdcLn7oqZxV41
PliyP4ZauxkMdsoyI9rlULL0aQFxA7IDa+r/yMXs8vDzvxjsNMe8KZfEjyh1D32Z
l6jmgAaRALxaWdiWjvamZ9q0LphZqejMeBydv2e+nApuZuY/yCpXixo42ggqsXGX
8dPB+6iV/cIxw9qReQaxAzbwJudAvZ6rWzRmFh6CTgwJ85BqJ6XtcWbZvrstBPvp
o64u8DvmelQJ8wrmOeEyRE3kNDg0uHaX0sGVrVgifbZblMdO8KIvSbW7KmKzbI1Y
JABHMDdhVFk3z53KAnC/oyWe/gd/zDa2q+shVXZqhEDTfQQtAB1Kh9K0CW5bnw6k
zk/PQ9qyJMo/qVap8wa9ldS21dSI2wY/oX7qM8FUwt/Tqa/LSblsy5fV622z6QWe
UvLRVKYLShVqJwq/6Zrszv5tGpNJAc2D/c/kDWIAwW3ykx784/B57fiTj0F9q4H3
AXkX0B+RpqfUhGeZMmU0bQTG726vPaffU8AH47j6sgpjwwPeaNfcEUaFeIwree/u
cLZ7mzNyvhVczbA1Hnuhh6f+CeaY45Bs+qVHSuv1if+n+PfGJidnN3UQZqWhQs7O
Jkgk9Ab+tQ5wbTPCbDqszlnvxoj61DPZ3Mi0mgRbDHCsnxdsC6bJKN1W7kLGwLpv
eDA+a4NJsin5nwGCjhvJLm+zb2pAqXIk8V2IqYoxURbCuyMhuBTSUcDDHWeDbWgs
PuHZQuSgEr5FLZNYyFtjPkQ9LBCo9ayQE1RZfjD9TCnUwtqc8d2xRxD7ivv4xD4F
w4zyqLZ9alpQC1Au2yhjjW5kzkDsRnDUeF1oZhZOivww4aDUjyHOtCDCudh8TLpl
jpJvtrZZzjWEA2UkZ0wRXDzajhK0TkTjeycuPrQfabuuqZiCpE7XcsRBf4c8JUBL
rlUwHX8xnhJiQx+0oEKVWXv3Lbvb2n8FNnkDglLyrna8lq3vRV53oKmp9XxJwJ7r
TdvMVwGh74G4By9MbvnigOq0QtUoCzpPh6w096RjIRXXbvmPuzIT05TwU8igzY89
pB3Nx6p8/06pj/bQvfJqSZZBm+40D7VEXpAvoz43tmDGd22b6u6XToFmUFMslYBq
vMpr8MYPbcYQ2H29wRnWzsIsK1fgyls7D2ajo3QscMNY4iUHpOsc/pOoUzsCeiot
3iRc0GlNJPxNAb6rgHIXkY1hA0eTa8KJRcfEDSD99KZRdBFzYpqTJlPCuZg17iVa
rWmlOVAQo+09f9SvaetuApvtieDBcMdM5kr0VSkBZIM2K9jazY+BAQPkqfUHeMgf
H0QEVHEBwghQ47gEkH2JkB1JrbCSHhiHgB/OdpTKmIsKYJuGktheYH9JHYtFqZ9V
CeMI2Pf6QhyYX1X+yGZ+jyayMuY19x/wfE0xvJKqPZPZi8+QkWP2LCOJFFLFNIy3
OHEHa8DZZSOIdZN8tWWICJQDTIDGqHQdQehU/vW4x2tf0ht9SwQTYW9yi/W/LQ6D
0QKOGb8068Nn8S8Zk2J4Xafko8I1jra750f2m5NDDweQL4fdLsCHflCS8C1B2z5f
8WUkJHBPCh7n6riksKu6OkT+mbhJKzs1iJBED6vMrdyes6BZ35fy3cJ07u9it5+3
Rz69lE8yMFqyXkfCiQnrjyVWgyrgzVAnP9iqpqEJCTep5dT08o2omcq72Xwn9Feq
htTy6NuHYD991U9JaB+umMGwcTZd1MdRljFNXyjuHHm5FQ6bfhKpDt196DAKwWOT
Or0v0v9+9Bg5m50nbzG8bSC7ZQUA7y5jXSypLIHrNT67yWTlimirYF/EKl4uvT5q
3JTNTiFjcvZMx8tvICZhSu3ORiTAv2byqRtKDvupFZnPFHSZ4VhtHSs8r6Jcjw5r
4EmEyHkKOijgn6ZwMAG4RAFUnASjlfNdSom58J9ru7BWIOyku0YJiKiJE1x7AFix
nw8NvU1NRyNpaIdIe+FlTZRBucGZwPY/7QdFdGpS4Sj2ho3VAeP8VFNk/RR9ig65
DFvyqsM40l6LYJFOKplOnMj+0f81MZ1mN2zJHoA8Wtvs4QCGzPR+aOcHXCUnq0oX
yt+fPgz8bBr1SVh9/9o4pQlA8RVNeQrgBnJlbUQ0iUiKsF0tuWX4gNz3vWdXAzlX
t4MVm9ibZ+8f97D5da4i3J5s7dLGClQLQTz+IJy4eQcANK10ijm83xo0fwJQQYkN
OS5yyia09qF62kZh2SPDNgcgDaoFRCdA6D0Tz6efHtWBkuZthRCNUDWJaN68M3uP
PO779xyETH31IF+vS6szkkxHlZ+AopddrkgAcH3TQeJx6H12ZSHXYob5m24bpmnR
99CVB9eZH/1oI3DUKYxwVjQ+hGsmwHNEMz6JYE+hoLTcPc4UgzR73i13Rpm+GgzW
5W9ekRawdMX6m8qRoc1BXfyvIKr/C9m7TM2plZd3D+mgLaW6i5RlvedxyGo+QlYD
Q8oIb/pEqWoC6GenSMnA6JjBViabUfeet5mz3q9ltTWYpnmQLeDRQGrFLHJs/Z+/
nEdfO9Al45+cGCPCQP7lhXYePsSEbGlrQEL9xc5VPxl+2oPA3SD64smDIHxfh2qv
6ZHtbvzdAD5WJjxR+yyP95KpzG+kOURCFVUTjxKB9nOVA/E07NeYNh7c8qdOHHH4
pncV5aUJqcC8vaw9nI/Czcn3HJkxlbVTFueH2zC1p3Ged+Fon3QhXxWiPSoH//Xq
MZhDS4UGO+ZmtwY5T03tjZLIwSws4fX5iiuBOvENP7OYjyo8vyw7jAtiRUFwzPvb
hD5qyq8OVD6OZ28+sXPsTFKTU7iFnMnX3gGmxBgr/hGu+c1SBs9iBHOUl7CAfHAN
wefCtP7q1YO1yZN7Cqs0i6j9ykm/molw8xnFDjRBNBXG3YdcvMccknbOELoT8Lvc
5FBNfRuMOaM3KNqg0nhArAvGiXOLO0+SMgK1yRVRzyes7fre/SX4BXSbeQ8Ko/mi
BRy5Iqo4k/7I3qTHFlRvvZE5QRifLtK2Dxf8Ws9l2BGNreHWQk0crTC9O6CS6U6I
tUqUe6lO6QPsyUlBks5QCjS6Xo5oDPTpxL+r5YYZ+IKlFga1Q2a6II8SsSVqBEfH
4ugXV32qUn6bMdPUWLpRa3vuzz6kSWkX+NnWSgbJqdV90eSGI9kohBZSpu45CFog
mWnk3zwOjNBB8Ry0Pp+mfH/Qh0djnjPpkKMR2t80vn2H+saWDrrXPTe8n+SapU8y
jMA5S/MhC9exTaPaJRgxM/elLytcWJOKHPC2ZRYpRhIR+Tv9o7ChpTPKLJm6l8I5
qHQMDJZLhcPeUHQ154EO/OhiPfSpX1Qy30bxy+TgWx9q5AG7EQ24SxiBGA98wxgW
X9X1x4gJCjkCDM7hFaoelzgEt4R3d9/E4mpTiNbHuBDu81ZXRcvuXwcOYtP/TQgE
wI6rzX2K3kHG2OXIxeaeiaGg8mruW0CzuV5PyHSIik4j1uRqXftWQC9vpQHpvke6
ZyaC8itfhHrDwpSu6iqRHU8BbpszAsAh3OXZA0zA4piwrvda8NUkTICsUa3rQxT6
M6RDDupDKzZXrEBBj+czQemVIosiJCUScfZSD8o1claHIaED0ZnOgx9f6YPj8g6q
y5gAeWh4QMh186+9aG9VrUuXGdkUfcak71qztUuNr53H9+ApvztXpD9aPFOY6Ren
ULpJOXhgrHYrr3dRYewMn8wjVoiLn993X+MZtuw33+czIhu/KBBuBoTcSRjPC2Nm
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
+HLGyj50Vlx2V9EGPjlr08cAIudR2TQw4pgjKS/0ANH2nkQUxtrOUP8iGP6nUaaJ
VGh2mamUER8KAuiFsXKEg5EqFufXo2YspdaM6M01ihsvwBQChghJCRDXWz+cPeWh
iRdRiaEicUm/e5022pg8nigUUMRSoV/VKo6asXUmjrvuubTcEqAYuuPoCdA9dFKx
EJL36GGVgDHoMbUnun92684KhngzdiaB/tt9gHFKx/7smPPXQbIXJBVL28z+IbiN
vn9XaDx4qA8V5wsFV7EurlzGsFdHvTtWvBCr6bPYzN6/Nqmyo1y4N5ehgYf5qUmq
qDt53Xx9XYTb+Y5nuPlQr/QgH5fJ4QSUTRTqwcKkunAFsqPX2NKvjzT8qVWjaQZW
dfwuxgA1c9ZmytGsB7k/z+DSEpXwCEAC9CBhJtjuIJsqsBOFBa0Exu3kFK0X3vkS
NnwZzBtfL5a18UgAl0ohzsNMSOEQgGC7f1BumMHefEnoN51XnfSENIQzwvifM2+G
1z5WjsoGlfWtYYYG32kH9w+nihFwWJ1fW+kQ9IiXTp5iijsY0x6qN2dVNi7YqSrh
PhRaGgwwG71tskZQ+oAGkBzBpwbf7Le8OCRI26LbC10t8OkWszx01+r7ENu4dFq9
v5JDTtDoDlXSls9/08peRiByfzw4QmNcXLNRNT3LE+j/dtL42rDNKPSfQZgIw3ZZ
sLoKzEH3+nNeJ4OfWZ/3hpPNdqHraeHe9U7wWtrDXsyHnr1QxGODaZB+lIc+8wy/
caAb4aOhNpuUsOJx0RJQc8ZdBDyQEdvIyOV5tDnCiWb2RskQB1q/QO6eH6aS0tr3
NNfmbvFYd3M1m2dOBjKsnYMvJlxjmaLn1k0c7vzr6yqNQ+J2pOEGjTkpuYWwpJsI
//dUsGM41l4u+AryuhPR2HAnDwsmn+6MvE1+9I3qWFjq+y7Pw5eDS1UkX7fuScEQ
aoA8ihIoWTqrrERUEvfcxD5AhS8PGT5HbbkvEHK/bKmj2ScxQazWheOmeywC5VaE
Pq4oCtbgaOBoky+1/W3VCjirLJTp01I3n7lXy63RouWhm5WZWKv3hnOjdAcOmJ70
9jhXlQLFjT0PFelBU0x0fU3Ty96PtCroq90uUx3wa+xh/cxFChBwnS2GvLoZdRCL
AWLKR9sPYc/HITKQvRb9MX13ZiAZ+XalyjNlZVn/SRoXlczaLNrY93tynBUEIEGd
8OYQ+iABUliMxbT1HBhgKLj+cEbnTP3vPoR0Kh8DpewqO2l3bXZnQ4a/E5vcSIDO
2teMexupeaBd3XCX8Scl0IlLE94HXo7rptFjA84tvPm+nmcXPj2IRxEJlp/JPS+2
Kf0p7SRLTFb1V3v/07w/wZaRiG2h8BlCISZzM23I4oH1tHkSX83j7S0tVw8/mQx8
m1XIP6s0QYLbAz7SOhpHwSJVGSXCCTOqlBBBSVDFWiWHa+eOK5KzZ/Ltf8tdlDfk
tftfZGJrMU1l1/7VmflBb1QEjxiMLWOxzuLcQw2Cr8VByDbVuSnc8xJDGMmcBk+7
NqtHXGbz6h/sf/zKjPqviBEbmMMnDIW9TKXJl6GqaRoSLCBR/1rXy4+s23K2a8I1
K9gILQ4Xs/gSMo5Q5pMi6c4/+MHE7He3lYMGBtr4vxx96PgCOu2h0TCJzMIm2yRO
/PQNOG39yK1c7Mt2eBHluEpDJjjHcSAfg9jLhImEoVQShEQ9cf261Q+zycZ2U1jA
w2JGMs7VALBJAb2znh5qJL79GallRSv4V7GbEluDUBgFVoTR63HIg/Jrod97Pvul
M8hL9o8VqvjqJITGVRmX4qOBVstzmRYBqpu8gtlh/BbZtAzaoZ/Hpwj1JiIinSHk
5SvAkk9/fqVWXHazBy9jM4pU7KpqnBOcKWH6//DL7MIxz+gLYt0It3M5JD0HNhZD
G2HD3IJ655r69c7UWRywRlSwJWvQjpNUsUEkwnSFLe9G2Jhc/nRK3eL7CMfzcka8
Se/ZL4MGkZ0QVg82mrkqAPegBIj593yoQkDC5RQuiwF2BJDGuGe5gLH8OVg9K629
JNf5o9zNN1d/FfK+HsEUurrR3momsZ6qxptYbCjNvVdpGRPBuSedgwR9qMSyDDSu
vCtrbVLjPhZPOQ/UzWeyghvoJhhQwG5RpaDIK+S35jNPaLjg0f5I0FsTIuMjDfRo
ViJx778sqyXz8IUXVEuTN4UC0SUsXsx4aV8eR+H1vwsHx4+BxwihtA2Qk8oCmbJk
TgC+QD2TREfGEPZzpGsGZFIJaPKOPCHxzxY1gFulrkLsW5h9YEsob83NXEVQsDAJ
pCWTzSXP3/WcAm/qr5TU4XCOjAngkYCNi1xhYGSf1UoY1hHPE9jxmn8byCoJjITg
7wmcfqyRPS5LBsLcupoykMQYRVHcdwOlHt4JrbR+pYQkpk6P6rdm2sv4vsGBMaUO
yVUO0JKZ++GYswhU9ExhHMpbN2yHp/PUor9dVq+4EnKSHmbSf1wRFZlb5IwVKBlo
fNeFqLVUeFKBXprzLZ3QFOyj0DbswpL8yl9pZuxZwnILPtr+b+zPT8+qakJdKz6W
FehraSKpE1Dma0tsJ4wlU5+148NjWg4MEtjB1QHCOQ7hkBxmA8iaU5iOqLSPhr99
1ktepW3lTTZx4YBUyTCi/OlQ+8a7CEwjTdRyIAitz7KjYP0sQT3jyKaQQAPW4aWd
XnVXC/OCzFbwoDwcela9FTuyKroUbB1u7hnTtB7MMbuxEJh/hykSobD50c3NCb3O
UOIheSkw0GdCLWnulJUHZ+eUzqLnry8wtbp0aRGWnEG23VXDJ6mqhxps9mAockon
Z3cDnhiwn/X4jRjsP/d5jHJDXqG6OEoDXn74pYlQ7b2juNiCDRnISSnq60ECeEk7
ujG96iq5NMVdp7nwSZPUiv2fBLXNkKzBulGoRGSqEc43VY5WY4WeSECYfKkuWZV4
L1Su7qQMZ1t0KwQbensGmePTxPI/PAIyMdYhKgvuMp5uCskk+WvVRCcBcbXpMVql
lB+oX7EqN1QXamH5uuOxracgEbj+Z9eCYw6MqyCRE9OK8W5/QMEXPBMzH+tBn1My
hQpyTzDYd3+op7SDIxyV7EOS01f6BwlqQNczsCR/ppGaKLIPyzXB8cW+dJ9ibYqy
SbVQ7a4yeYz5mkLrtBw4PgsjqawGPBgL1DTcQeV8i3FqUqKfgbVz9CMS3PPQu7mR
yoFcQmLTz1hAJTJNQMNmxT1B5sQeSYEVTBQiNvkn2nyaRLp986GjzhB2REp4ivQD
9mScvBuom8iicZ+Dp1sNjvaVz+UBDkuq5RZkeB5xn5k++p9rALcQXIvYIxB9HeFZ
Holfx/yB58sT5fHmpfMgGh1/vJ9VOhGUW7//K0slcgsv+Fq4knNeXS2GjPgqJQ7U
swNl0hyZTv31w4m35M3ybEIqSKqdyXcptpz9fOw7lhDi2iB3BHRGGLntxjQEoeeq
XeyqH+1cUw2ymVlpc7gDRqy+5zGluGh8/vLrqgXHGAvx8W+7Wz6EQiiZxM+0rNRT
t3QBIqo32iYR+zRXAu2VCG0iVFtcOh4OZRDrvGldwCKwTXp/OSkSPufBJpARx+/c
b5knlya7dCqpFmw0BNqMsCNd69OP49Si934JrkR7ACVAcnI5B7nE0DwU3pLIrLyb
D6+oYe7q4OAjAHsWKX2PycCeUpmVpHOT06l++UFQjcq3Qfd1kTQsWjsXRwRgyuaT
MPmdtWrS1efN4wb+09utDxGcHSawBX6dbV9E9duFTERuYrT77P1X/hECkYemqymW
UMnAygbg4hd+L8WoYUyR5O3/TQglSICtnfpHEzr3/E27T6LCp8Su1P15qIvEtcR2
Q16H61Ktnv34l8Yk4zcAi+6tpbOrnTwNTf+h8UNiOHrYcwabEIqkJt2cXzLulPuT
OYiUqZXViqJZvwy6DJ1zHX4pp8SjiRDnzDHhCcPVWtCeEPa4iVf+BRh5XPuWsFCf
IEwdCwdcoixw9sJgC6xFSosnKxEUXw+aG7YRkB1Zw30agF6M4TlSnyihdpvufATk
G2keJAT/+zYw6RjBuLvTQhT1NcP/0nIyK5s4D4GaiIJ907cBBXtLvJWF5tCXiDjd
UnC1nF8LS2weaC8+TT6CGnLCVQwnt+cv7APebS8Tyru+4OpdyxL0TBjUkEDHOhY8
tgSWNxqvts8FsE2m5G3zvAHF9oif5GsWHLvzJEwTuBA9NB7bcbQ8rmkvK2Rd2adB
JcH/m7sa2Hyrold4/SP9od/U8vuSWyANd45d+0plTNvUwEjwJxHAOh0y8LYxQRee
3QJWUbKFXQ7RQYMYbxuKpiHho6+jHoYPBRsN5emJMOtMi9B/dh4wLtkIzzZ6sd9O
dlQp/h3+7lw+DH7z0jzl+EQI6rZlUcdT9TyEn+NpEygbGNARvLC7yzVBG5jkvo8N
yrMhMMfLZIM5IiVI2nAClYE0mJzAO01SjLj0GmNqQz7AKdUXsP6Yvmc8VjA/+eGR
66yNAbCKSpG9tRjL8g+ffaiYzk6AutSLMoAmaGoqE3rri2E3vt9hiJeAD8Gtwbvu
Bv2IyGLigI69IP8jqxuNjTz1FS1xkJtvg35HWqDq8ubzGwxIebZSqy1ubFIYoBBd
kveaIAZ4vw/Upzr1xPaSm7UT0S6k+TZhjlgRhBbmEKAPBmu7hVufaBeCR8p3SnIc
TlLArsriTOzqNCA4fsbwj265xYaR8VCcT85NRGQF+js64szvhMCER4EOtpQHdBMJ
1dV2qEttLGDm/txPcHxyv69BsU6NWLdIc44yBqWUXuTQgVd+kf7tmLkIArA3hlW1
/ywvQfilCRYNSTbmh9sPFD8mkPd1inrutd/rf8HTrQkQKRWMyPhctCHTijfjt7up
zy4g6JTDydB/7KBG2vx3Mz/tFOW9oWiIl2pzmhrHzQxJVekxBz7BtrUiqOBPNLyw
glqB3bsovgsgKfDONxsOsXMBqU7MDeF6wsoqrV2S30eT31HxnJirzaTxyrhuIPb/
2YYKSFijw+el4E/1hjshdwX4TGeKIf7K4SkUZITdIqaWPpobwZQFtJUiOavT0IVh
IKJAIYElFJaY3KgjVvH3+FKm+/2A4ItLTMDn468aal6trd3cB9nfdmYINCxMPmWC
PS/vLJixqiKlN7mvybzXGe1q38gzWFUDd1LFeqZ45zMrEjvDiLHUMmnyVrQoCJWR
qmpdsWhyvB0fgEZnzdbNYV4HuvQK/N79ZdEPcPN1i6oeCqLt7Z9pQZuqbKNsyMnY
bHYUS9JswJpSgCtvHWDX5AL/IaPEnZ5+M9A11DEu5WmoY1ZS40E4mclcuyXJMlEn
HztzOcaoqjulxznOjl6HYGFnVQNVRxMPdnxr6AimHjkBoIHN8CAs2ltWefG3GbDY
zdtoH6vgKslLYZmsdlFAnY5JxY+blOexSZlk8BKt6ZWOghx4ILOPyL9DPzVpSgsO
AEzqMkeXd0nFfr+qRjAo80ZG901Bd73VEwj+TvfzPOgBKhmNico8oAi01X+apWY8
kbr1bnmEI4pc6EsUIX2q3Ku/a/rKg7NxpMTj4SBmPeQV1gGOsVyFl6tAVCQFJr8H
iF2H1y7ZGHaWHIITgu34tgRmVqNYp821a+msOlIkMuDy+CfkOBPpLYtlqb8eerhI
Fs4ULcwIILEbwFufJ8FGhyb2Q069n/DsIgXwKdq84V+XBRkucTgoDzx8A572IQKq
CjsdVAf118sD7kNgBpLR13alVEUfGXpSBekK7JBD7QXY4NIfSIe23BQ3powghoH5
mbYSd5PW2fWtIHJAAlMdOQRT/nVDqlgyl96FWEye6rmPVKWO+IXSFkGBHYehvwsM
FBwK2e8t8ns7Vrs17xJSkM3E7+yGcD3ZgaJsYaFjp4ErvWJ3iRoaQRS6WCtsEC41
XkGCk3AtGZoonRQkWDAUZBke0+TPGvaMK6l0IM1J4F6DIbLfu8qsevJnBFg/47bX
s/lJjDAgRDc+hAOoBcdicTL+Dh8rCQq4noPabwlbHNXxHtV049byA8UIhPpQ6I0P
VOCGJN9at7k3XP6nZnzWIsI0pRUV7WXtLZWyG3ZKPTEeID+zFTG06F24ZwfyLT39
nCdxDU6/g4It49p7afwN/iZ03mHOTuFMn9fysyVg90bXBSbKMrJXO0AnDx/4eWeY
E6yd+t0I0L2cU+2tEdrpAbbDR8EZTFLwlz/EaX7nWCKqJk2d0E9yu/0U/mj7ysU9
ao8KJV5wJjUbujuBV3Sw2rTFGz6eyGCauzUDGl2Ac0rWjD2vi4r/7tj9xcFk09UK
RsV1jaCOU4o+S+nL48L7CjMWn7xL/DU4x3lSOZtLVKf7kkN0wv0qoiP0rqMB7hdW
4A0Un/1kzJwK7BDzPB8ayqxjmsyptki56bKhy2evvdIbfuYT4TByLZdHPG8Nrltj
ZJ7nN09Kf6W9k6A/nGHXKgiqUCtkl4Fl0/YvpnVzW9gHqA4hK4C7usLL5vVbqnOQ
yN9YOrygeuQAfMheqP1iOD6+9aWvlu6nRlMN57SmW3e+D/MjBuf3+zaZz1mwjjtB
8JHnDDtLRrdDe8vAOOXWHkdCtCgoauxACxbp4IHHzrOL9/jT3zoNRxoVepOpDGEA
caYfwO9gGFzDfKSlglJ+3pkP4JqK1sUK2xzf1+UPI+f6L2B19eqSj3aoNjh7Ynxa
D6ZI4P9uoWOmMsjh1n2n68CYF5CpTfQhkbp+DnowQ1/z0HCJlaTiwpL6YKeopGzj
QYL+UICOEhBRNQspF2QxO4BV10KDMWHDPG0QsGQRZ2xf/kfi7ZeIHsYf5OnN1zxu
tdHIzMCj7l1MBm0Q9GNJNFhWOOW4CnR/wD/PcINw1bnwLKPvx/6dVZf0N8dfqfpT
t5f+GGpHBweUrqs2JuLZK1aUkJBseBY8vN8RrWDQLw1g9KV1/DcaSiokdEQu/ghJ
qJv+qYiTHUAm1aRBCEtn1MrcF71bAt0WHnof/PiwN7WIAkE7QF3AAAhHEDiAEGec
9vXVokMFusEg8SsmV4hua1vy397ZVWig8BLspu/CHBlVFA7alY0TImqMtXfN7yiq
SRfqeyW7woG+OnfbTcmgclpSPhZvWgw+JcUlKqhG2mXvOr54z3DPE714YoVa1p0i
NGvI2MPtLX+zmIy5C110Nt3J868NRLY9LQSOuZuJxA8ZDOV7hZ4QGGBjXFiXpnEj
jYDbul0PxmUBhF6TdRRAY3bgOtKoOmqu1oqjzLHmrOpBMLjtaOtj+BkY4BSJCp7P
58zsapqEwQKCakWuhItixsQR5ucPd8S+LGraqBynu+LPCAt25AT/f6O4kGtCYSoG
nz464s2W4kbefPsWWlLK6R01lJrrCDKT2piH9oFQG/vM5Uwo4OeQKKdwRSsHwxMD
p37sIr/cDFFqCCWbZa5hZvxX20Osi6YOR74gl4IpWY/wBInDMmjmSWwvoN7kjvGD
6tTK3FP8ZQGXP0jl5ymis5YFWWKoHmc9iB1UrVDufA09yQHKFmDr3pG8Q3gHPG2I
/hBhUBiP/rlIZCOeaDZp2YHEE3xZ59lD/uuae2vU1B8/5zMNoOJLKK9Ix/VcEN6m
xedLEI5+L8ExZC6nMuJNYOYS6qo5XpmdQ8W4TDnimSohrB40YCeh30xNiPqaV+hu
So5wdppZwRQTxLgCq10S4oEw1u5kAPkH+/hK5j9w67gl35IpwLzxsFMN8G4nKNp0
RxzHcy4psZDkrBSzeONtwJFVUuXFcLl/v8MYhC70qBFjWL41aBn0Yredxsgcjh8X
TdqkysuRxg2VY/8QXxj9aoLmELbPJIx55J9ZLbWoBGRjygeexkvSnWwb2z7JXM0x
ecxr7lJKY/9j6n8FkWdbcmTLf4bMMOndH5OTlJ1GPjuOwgQWei9kh9Tat8f8yBIR
5qjBHLrb4HSaK5Ty1o4lSBx6Y7exUf0arZN/EtGvsZUxRgJM02OEbmhVLR8e1Tqv
AZH8AUjPEkHXHcanQJ18wfF/C8gLcFatxdffO9GDq8WomozG6uunWALwq1HjbFga
vgDRvtscDrhjz/K7nvjGSDVD900SQlpZELHsUDqIb0cGKLsR6AAN1MJGTCUnqyRr
iNde69V1ZkjgvOdhMi1iIrWZhCWhRHl0lg+BVXSZuy1eBGL+CelPOWkV5eqNiqoI
8yDcEwWs0aCdwyV76x2fg1JI2BjRxAndCz1vfY5TbsspogLI22CNFcrtiL9lVyxn
EIi2GG1ootD3vkh8nKV9OHAcfCciNPxQ65bH4Vf97opWLORyJ4CWePtXNnwxQ0tX
QYUP+x5SfVtzSTEO6VKFRSUuCjMuA+1dCvxsEOjjZLa85p5hUUf1szCQFKt675GC
qHT2ciEJx3UWHWEGbUUnwL7UgWUdlYxLvMszaJ6xPpeSexwmufUjAoHoFH4g7EXS
p6T1Bky4Xoz7SRdW0eXpNPhFZqRCvn8zjIm3Z0tCTCQ/p8v83j2gAnVLGhNDbEc6
FLxa5nMxrSWKYQYt2n5/jVaZq/vbLcl/ihDRBrQnlx/GOr9/o91m9sNxdavM4AUx
VikQrKmglZ4a5itaj8bP0APT0Har6zHcHr4UTti++a8t7xQlMllXo2S67bwNfkdW
QnXWf2xZ7ZtxmQnMxn9F1vhxYLQ18cPceGCxwUJpLZPZS1jqmO/0+30/Pxw7cZzW
byVYfTxFXoz+ltYouVWUbr5VbQ7zLi3xZyIs3ybKzDZHoUl6Mog9GPI8MNts/2Ul
for/NnCulAFtWQTuZBMQiDhX+qWRVaRglt3geWVK++AbiT28v6oYWGpR9MBTYpe8
XB3QZP7AhHxm+2udE9htpyhFM6XxSHCPJ0zfzl1ILgfDhhCK3r9h9SWyMIZF3hFS
AYepSvPOM4uCyU63sXE6n1IIUn8iKdAYefZu2lkIsAWvNuAJJwkNd9wLb2KRO7Se
4QT+9HFIjIbl1OTQI5ZXGH17CwpaG4AVdk2vgNioC2SWrxB5ph00wqs1M3Y4NSRh
awNy61+KS6hBbOGhyfvH3ezX1db9hn+MosOpD3BZcgbql+gOBgELCIOMuubve5gB
mNjL2QbxAPQ6bUhI8MIkAGy/ziFqamhSNkAfry0axGhx1OUUEESZKFpWuwTX8YC7
8SkHjaqpDQ2wCXhos09mbhUchr2a+j1rJrvzK4c8bkUbylf2ObuQUgtyviHtRRmv
x+EkY/epELLvqopiITpPVGNpl8vV66BLMwpFcSoG8tG4cXL5iZDX6FiE2lhJ/ezp
8ndg7xTh26k90GJk9THoSwgh81KjL7JHvE9IWa+7WH9qcAHHmt+2AIa0hex0Uswc
TOafkp4VsPF6dnWkpi41g1+6ADSHUBY5LUzuMfVINcSX9ngwEnUjUAObLE8/V5uq
cGfHhQzLklCEX5/0KLupKXe4kTfL+vrQKF3N2rGo8ndJ3J45ppMk7DI2LikkSqgY
H/fdl5uHSBa2zw25xlLRopgmo0gR9hbzk/JcfU8wjLeOr16XmKfKKzvf0kkguCoR
9kLZxmZgzs9+u7R+f5YL4qlGTyxoRRZBDq7oF8I9U6cFKGjEQYxhY9mFFAccnu3R
KFoFzRBF7fkpQ9KIC6x+pW3DUuG3dA99lu/pSyEtOR+pzZ9TuEm/3VVMmteXGFeE
ISznJ6lhcSutNU/j6boQeUkUf5FJrpCbmsVV+FlFnfkxPQL1AT/VpcON1AQW3krF
8lwug/NdKvbG83nkgev9AUQR1RZCKpzrFBonrAQlhZr3LdF1TvmbvAZTj1idO6Au
H6oAgQp87PkMIblPGB2VGrpMT+5jZ79wJHn1cKiYV7X58yhq1nrO1r/3S7wKtewc
tIsvx79Lf74FJ52eOLT+NOXPqk5W/g4XSWl9wQxiTmRe2eWAWvBoDG0+5pykjbIB
7CyF9bD3waDeJ7Q2aeE3uzd0/CVNkxTXaNTo7jo4nclcOO1oI4ceIW8l7FBHsjLS
I+Ic0bkpB9AxX6C4L8O1Z7wpwY5w5zwhFDzfFGyvyz37EDZP9O9TSG1jP/5BpypV
MUTVlkVVWRgNew0DD8Dwxouw4Glru9Fqk9JIFNAjYCBTOmMgY9HGhvFS5T+xuUSf
j0GQgoiAihgkTBeI4Am7ur4bDCaa+29iEY1kIHsptZMiyoV8QqcLWsoq/NkTJQjX
izK6H+7OTSjIOutl7c71OHHU8/mdpqniYxf6FUV5ouJcjfDoSuezj/TqhC9o5p9Y
RW4mPmCkUsKZ/Mpd9Ajxg4mZgt60MAAoVbLFFq7dkiAIJHbBb4rx4XMKK0KK8Ftt
Dn2rQo13ueR3aXNjswWg6w5YJdZEXXF3exMPfpeqdimPQ+U9ar5qq6Vbx6iMAPQs
dOSF7tMmA45BHAV9pFgVCum1gNMhKVKJJlY7CLa4+lPY83jx+sx98wMaGHIntSPG
YNpyJhhRWlKv1aL6PXp6ISH+gpHkv0VpY3apIl7GcGG06fT9WxWsj3EZByVZYzAS
/OVChOqbSMjAPxSz+ZsDSYNzgMlJhKiezLZR5g9NM3aNcmbCmsWL4etfR2r5xSdP
J+7vP/U6jyHFo/X2K1nyBDiroXBLqD4myy7yimIXPYM9Nf364RmYMZHdjzPwpInH
zK0CpKPVDXp2f3sdoUsiYeeOM6CaIZT+75bAISU1Ag0x+7qAkRIXsbueIxlv67n+
2E2mA25M+hJm9NMSzqqRrlccQftcP8KDeP7asWARSWVIPPZG/Z+UK9t9NQu5Kvnp
Wt6bmzGXFRh7vV7CYwG8KfcPjRlFTGB97GQqEcbb5bQ90G0piJvo4w77HwTKp2Xz
5nrhkGzwpJaeOw7EWRAAJz/LsSB7FXceL+uvHlGwQadL2MNKMiIOV3Z7bdC+VUkh
/QX6tNbduZ6UIQfw6Rg96nnv3gP5BUkG3ulPd9FUO0dKPyAmSlfmAb+9KbOI9VgY
OKwgwBYJYA+YlufIDFYucUL4aGmrYbz7bRdfUskvv+z/32Indz0wLApw4oat1m7K
UrTdlhbrk69xz4ZIgMnIx9wXQUYfHZfABV+3kmRnZe5uv0f5MPmQhJzO031iqcr4
wQK96FNvUBu4eszOTjwKvAayCFTac35w8QGH/zkBXhtlX4F0aehtrVeQKrskoFsS
9ILSXXgPULR6M5GwgKiKtIM3avZzHpjQ25JPhrkBE7m2ZCCYk6LexZZ4EDA5Hn9N
aITTQWIGa/GyFEKZj8//LAT8f9YjxnHRCHSZVEBK+E+galizOyvonsI8cgnV/+BH
EtF9ksGtocAwP5n2to54cri9JQh03jWpvvqSLcKWTW1kzkcT/i7lOfbAmv1z+N6U
RBI4rBeWE0EjS8dRO1m3Wk3FuQBgByfwPFKKbU44bMfoReNfjX8RXc5kQQ04bLjJ
0B6rfaqyzRgXbrW7kdmmTcJIZW7S9EKlXuZDf8ndie9dsPWa7dbZNj0UR35GP3QW
kLgxzDQ6CcpDqzvkvPt50OJ1rJYtfkLlxkAsKRA/UD2ldT6i12h7ljiNhW2KdYOe
uGfIM3B+tEIGRRiT53cI/yW8TSu0zd+VGcP7tBkoCasPqt1d4EAOCunfINX+F2yB
3Kc60L6lev9v6VVRGyX3E2wqr1nNngyebJagebVostzIo6KUof9ZRihFWy7DgxCb
2QU4MDXzqOnkmvYyCulLK0cipdRR08lhawfvFEpQmJWueZITz7WImEzeuO+CVOqa
OkhwkT8JuI6fzWjlSiy5KmUxs/ui9UaqkXDD56s5g/dz8iyz7Q1GaPQPLrlV/KgB
azsFZFyn+p7nKle0PkIeqh/2xPQ3h9UURQX70JjwvJ4+LJvNd9gkHMarNaYot0FT
IZNA8BcQhbbk/5j0uUZje1vEI6kIe2mDztJ1Gng7ZAsaxAaa9kvM4A7wzOlHVzPD
yZpOn0FImL+9IsdeA8bfFO9p90inOVjKdrgo3SMVOShCaJm1RQSFWBw7Mybyy7e9
yL/c1NEyFXpzymnQZWutw61TzZ6f8xGbHRN1CjNpbrVZkH+1O6UlXVjKubEq4XF6
kGXlwj1qRdFLtjV6I9gLZ6UVoguHj9nv5jWHYER7PFgu/WWAGAXiMrvW3+lA4/cV
EbwQ1jl1TAJtTDvjBcJmAD7VYpnGPlGxZ0SzHidaQKTxyBBohTHbXujnLl8XUDXf
YY9GJOI8j3f8iHy43YXK2lVDFZXfDVLNh+hyeD2CIZgjaqZK86gtkm93Fi0tz14K
pWMPifYjWXpMoQEIw/U/hSvxrbKUHl7v7QuR8jcjdLJZib1ixqdOmRgfI/1a5CGQ
R+0SgUnd01ErSKXr3lpZ9sKRr5uIxsvsIeAlMoEExuea+To/07DO8dIg7c9LZ+vd
R9vSRkNJ2ofS0X68Jr/1LuxXb5KCm0Sd0nXez54ED3L7r1hPqhF2w0uL5nd2fWCl
Iyoe+wUxSbcDDJa5PEUJ4j6aBkz86n8CJVBpONymurHlpi47HHaV5oJItsNrp/1e
uJfG8knrgBFiW1q7vvonjAOOV/rEaiSq1d7dEIf4dl5T+NfWNzqLnfKSwMouk5gq
7C+A2syr8OUf6VVX3J3gb3nipRjMEzBqofaV6DQClv4hkZEvxKB7JhFOipDurZ1h
+xqnMufQr/T3TXJRdXTBeoyK+JtsNQ/EEBgBA2itY4DgjKri/6GnMatps7MU5Ooy
o0gIwovvQQkOJGeIkJeXqvgYCOQLQSqUKENLiWqya3yfTGNrHcewuUk/xxAgWP07
g/I1PRdEtAkb8MKytHvA0hBcGIVPizmGDVkluGnHEwQm4WB8ag9QmEu9U/EfXSmP
t0isi7rbrBqwOW+quZ0uTeyc0kmv7VKt4zs7lmJ5VtDSriVWPexzQGKnxB8BNc3/
dksSXe/3nzxFlslnvzujOkgIh+SO1f1RLxHpuU1IVD+Tkb4TPfUosnc1kbKzx9DV
GYDRBkTJzYwQXLCi3k8NK8pQSCgph+dAqYPg+L9ULSnzXHIwjesDbcdFVykY/olA
PARMbFjDQx0Z+7n/cg1635MBaIGwxUS6KEJDAzsaFF6virqe4tJ71+q4j6n+7r7s
mq5F1wLgkb+2otODPsyqA+4DSPs8Uel33FuhJn9UWtD3wwjigwujNVQ0uwquuf7y
o4oLKtRnTz42K5PAXIC++ZXt59wLPkkR0dxZQD1KC7OQhODvPVvncAZYhd3oUEGL
1SOlZDtRJj8uhecZ2/UxuWZ3rJ+vm4LyWU/A56nbt6S2rcTVvcAdfK8FRpLOE0AS
UUEq/LBWPBFD1lLM8GF1eLxS7FDWPK3f0b7cStdpAnGYUuYgDdaHoYe/JzVyw9xm
inv12qsLAkdnPQ09id3EsYrS2e1EXH2XC10HYKNq2jOrpLE2vB7vsR7YmWIuaKaO
5Isp+ZBaqNmYMIMuxdSFyNLxfjuvAJVRxRglFsAUzU9tBNWKtU3ThMKNpf96Gnfz
MykmC2dott32JQsXyV7gPlxqyUgTf7lqcUgRPq+4F3NswFu/I6fYgQWAZiV3LkCW
SHt5qToiNi1Z518jeW6G11sfMJU4AJgqxO3KmceYFNAbmBLgzNDxbpUda/utYnPd
lAiZC/bBarTjtSAA8rFfdbM3eFfqlYynymHCh2TOcHJ2tJ4cLrhan77vCe/v/fJa
iNUboLPLjFSeq2HOnuJFFLOEPuEZj6R6cQEpc1HGXGwr69oODWCdZbBhtV0OYFZC
Ymsj9McojDky8mWWBb3Mmvu1LWStmrbpfXKTvjMkcZzZYUKUE6T6CJNiakvqiuys
F1jEOhLXTY6+se4DwjsyecgjU35fvcranfdCpUTXanuf86yuNF4IZvMPr4+PBtF4
2XFTuTZtVgnGmMsPR5eA4PLt+hZndgE+wg3+pa0YWqId7natrfmKNNYaVDWX9dcV
Jsv/kQ37Wp4Uku15an2byf+CNp/QKefPhCdci0yQfPJ/Susyo+2VM2cqt7B2x0xL
JC1TCDpVi39ezqVkC2f1h6/M4nRy9UlNiEgO6J0hjHmhEXIcnId+Urew5JijmLkh
LQpmAVrxlnX/7tCpjcjm+aPp/n2PIZXRnm/wQxjYFhQeMve5ph1N9wN6QBRFG5xT
0cU/hFqU9dKY47ag7As08HN8U+gEO/SMdnQOKg/BCBzOwTF4GnzLlAEbFmILnGdL
NTfyLQfTeWepRiIyPLhbfeChOjxtmguvSsFPIS0WfwGOB13Rr0ULZGl7w9V+CKnP
MwfwXNgFJnmZ9Aj2jxzoVnahke/OR7yOJz1wmHDsv1Z7reuwaTjFzZYVSBKUvS4r
etKzjb099OwZ1t4FrECMTrS1f2zp39X7M3MsffctYc4Vo57PN6Qo+TustNEEXXGD
GR8KlNCKDIs8y1GneLMsP8WTnvghn86DswbwnIwXWj2KUuN/Xlf/7+LKWyxDpxCK
PMQ5V+9SLhIyGORjfMiVdOCI8Gv4qIAM1hH+W+wZZ/7aZ3/Lrmx0s9JQ2tRY9AXq
byNuwp3MyFmkVw1/Tl+/ersN9/lu0rWorXifBCkvfN0tYfyhQTbMdJgqtS+C+Y5O
QjBBYCyEWq941OibMUAAKGzP46bYe5jeuNnjVH+Gwa3O2ElNH3hgw24aAhWpRJFM
OZRLx1aFeRsg0L5vl7RXqz2DfThq9YPQHT7V9Ps9iMNtzthlKCxFD4/cH7OBIT1E
qM8V0QnPErIPRKtqgw3224E4Vhxz+F+KsCmDY8AfzApZNUrLzJoozwxPqd55GXgx
pMaD1efP1sCFxbmCaepbdxhBTr5TaNz9/L+5IBTtIJhIHnpuciYDmMslJboYLGep
JkWptNwZBmAFEaF4xqthEigdFSRKhkpUGKgpPh6HA2HlQB11ut7Wz/L5WKwPuFyM
YY15gqukZ74TDik+SCOufBMnkm9XarHhllWMalxBn6rKW1vkt4tYPYd49cxEc0i+
rAtvxiUu88lB5wiIQgnNCFtvDllRXPivKyPJLpPtr8k0jhffY+C91kNbnrpi8NqI
qP8QX2sOMVaeBEpUYsoe2tsvophddxqw99QFZ34jE9UQmNU1GfOOJq1GK9l5AsZp
EXdfCgTHzBS+BClh38Pz07j2NoKjHsLtR5WJhV5I3USAbtr9jw/bRHc18c1npxyq
Ltp6yQoMT+FpwJMvUNlTvKf0vn99H2x4A/Y7TVsh4vmiEfei/WQb1CBjnqxgwIEG
TktXoAY6TMC9V5CdRauq7o2zIGzN0inSEet6gVmMq++5pq46EYqS88zvLsYaSrSJ
gjWwRXvd6FxCxO95YZjGRRkjWrhQaKOSUuLZkvFAQiZJ+Uyhhc91Ixmh11VHnQnN
P4I/LOfLtDZ++LoEiYVLMCsFYeCspgc3oq/F2Sqzguz0WWzLUaByVZf4IN+e31P8
i4VBu1N9FNdUjAaZkcyuu3Wk9zgqjDCymxu1Llvq+50RH4HoI61k7ZgcGxBCWAB6
KH5q/5ozGqyNgUtNGZGrfvxJJWHi8hbhUUVCTyN7+fiemc5MQX1d7E1XNVisc67T
fY4yVQtpS75Ony2xS3r0dTQ0ssiRRoVSx2fIARFzcKdmh24CGMiPKw1/HlsVn/2q
uhnpD4DxkKWFaLW2L3LeA06fakwHuJWB18r4+2mulH3at/Du4BrWriEk424GwYDa
h3tyMm/JarwgclXzQcZCHJeMRCnnyslff+cjR9/9VfTAYeF5mXlPxldVmOdNIoqI
r6A4/FdUhDAFpC8mvGWPt4+X2ARrxpInR7Vq58h0+hMpED/SYsDV0rwfz9FUkwKK
jLXwR4MTFe/HQEpDeSrUKYw17DBTxrEPGmdx4M4pnG3lGJ3+zqZW4nMhiMuDwlYu
kwXYBOKxsjsbV5LlWykqLQA75HSwSPJ32+hZgtLuHngqIFL9OHj/VdsBrhXU3khs
m8FRSO4+cswDSByqOJ5nSVhKo5I/qcJGYL6PspFb7DpDx4F0L8dP+f9iRQvzrz4A
hBq1l/KrXjWmrpACMoYDCyjEW2wBiwlYyNufQ9QJ2EicqKEeBj0/FfsdQTLTG467
vpWNFFAObuODZlHz/JhyYTKa6Qdg81WZDYbL/D17aL/FbPfyEiu2kodMM/udYbyI
eBTW8gXLYEUHhTQlv/p8Q8bSqMdhFRK9e5WCNJFawtKeZ3p/kdViKT77Zs27gdlh
l5q2j7oAt4cCiFmN2F71+/syPkjUqCivvkSw1ciADw5/slEy0rvW9NcIMhQEJaj4
SzUZQGk0RwD/JR8FqCMowA65L/Tp36fOIPzo3SPXUlMeEHC+FoSsx2RYtGw+KnJj
zvweR3GhCdEN+seSVjCm0Dpo7DR1spSndVWOOUv9ZK0Yl0OcksfO6DzJKRtrjPDz
txXwVhQM/B0XJBmzdTZGEa6q398D3eA/em/0+tyjuJz3Ztj8n1dodk0P0slYDesA
5RH6u0iOwXMQAUCJ0yuSgwgtjvFPmQFPmfPQvlRHqKg9zzBomOq9llLWo/NSqEPN
Xdot55SjzS60GoiynunbANvwWRk4eyzZLrm+WZfeR6/yGfpDrKitAxoNML8m4CBW
b+yByYyU6pgJcqz0UsTadculx/0dB2Z1AiIU7COHRtaUoN4dUAorYVl/A/Gb22Wz
FkjuNNz6glm97i54OEaveS7DyLIOSbSiKZbVoRilkbQ6tCtkEJfG4vOTq6lF8QXd
AOMmTOeQbl1Q2h2MOgL3HgB4A3GKtxttkYxalI0itdkmx0k4sJGX9mmfhRBfyb4B
HDxLh/BWxQaQZDfQqLFJNnqg4bYZH+3GUwz+UbAvfPA8H4ouJL9Jjr7pEdYflEPu
6IfmCCc2uNNrThUcAkbkG7gJNyWchwqATRnprLvD+cD4EzVibmD5xyz+VYPzzfS5
Jjum5VX8tbC8hP++uPrWBoYeJ+QePvLJnmXl6bT/9nwYEhn4WbBUOcY5lr9RVczy
XlhsRq6C0Fq9PBLOaEgCKemcAQMn2AklUHVwOl22OhueeDwvMW5BWSmsJVu1pkUL
PbOb7LCgFYKk75oHniZZVMeMxJZ0v7hOsevs7D55TJLBfNYqq/khul1KRi746OO8
o1Scu4vNFxIcfi2cXtKiLdzktTtC7lqkjb8EFK6sYSNaiATmn+2FIdrLUjlLpApw
YjinzSPM2WukZZhOYIP4yMc9jhHgRPc2KN/JKdc9ldHw3N8HiJ+YuVoYaRTPggCn
DgLjNXDzVmTXR0MIXhWTtLWJnFGsU2QaWetIIsEwrWUnjAM4dQLrhyBcEjQHoydX
Onh33MMJZWHUJO28wChZrS+KEhSKtSHG1PzRy/d2AulPbFn5UP5b16iR7mccsdKd
vXj6hDPOto9MYWctmS8tdSr8pfrQl2g9tnKYsjbeAA7lxTwhgryEwGkY23nJ1ZFi
VW9C77QRi2zWC+SqBwKjQYZbjhxlY2Ezjpd3rxQhCqEsD5YZtb/hGqfYYkaxd2ID
SNHhassynnap2NY/IvfKLw/1TE6wTKJsFOfa4ghl8GU3jI0i6a2Wg1ANylUKxfZA
fu5OE1Hw/H1VFy8aILbH2OgGAeGl3p7tqh0wCna2uRCxRuqWA7rBmXdhEULJ86BX
nxC72S3y9IHpgWNgEX5QJVax5ikybQvTUyO6N42CfR0J2rhhMPfPo+a+6eKqPrS4
qmCv9B7dSW2yFH+O+8crENEQSkmMoteRD5UomY1ST6JUTEvPDE3wkoYB6Cf3PI5A
92+IFcllW14EcWBvaJb+H7vagh04UdXkgCFozqw2yPdQXPAWbYbTwwIKoJi3DsKE
ObgwuXrPnjIaoP+G+21ir17uRiCXal9TcfJc19rMy7zB5E3o7dwOJFYwdgVS946T
Zbdfer7HXk8U7z5EV4rXBGwxkAHnMCezq5b1pTDe8ZyGNijCMm2W9Q+6UdmXYO8t
TeQgPE5eNIvdBryeuUOfRrClK9lCPtgiciId9QBUBd92tyLBp1FNxu4MhiPXyvAd
qMmtKo1rh9RSstQ55ttiFtOmIoCCYfU1PVwpwP1WyD19+fZnLxktdBUmP+8VQaDW
jufrBYmIt0MpsWOrF/8oyiV4JRF/9Z0PYN6DwpyJDQN6J1UAq6ActB7lnd8lWKEv
wx8QpBHDy8TfgvaP+3Z6aSenZ4CjsRxZwGFFyBtIHBUeiU0qClKQ3BhuPnFaa3Oq
WYB2LhLBOKscS1GNNjhe6i7MQwp1kzkGMnVtjLF2iu7AGVEd7ECsnPbBz/Xv4bhP
pntEP6jo2ETanAOdJXKbPr7gJkLtu3vC6cA56cSdsV5pJdXwzfKrK7p5y4xk18FU
0GuHsI+s6iAmi10R5D4fD9S+MFkIVvvt54+869yP0Cfnes2XTwLst+Lfw+bPKwZr
vukCQj4lhhMvZ+Cyk1kwIDVxGD2GrPuoSR8gjN5euW0q2rI56uxyz3vZftAikKG9
afvbwsyGThaMgiLtgokw0ARKLThivmMWexpyK2MNi5JLpfafV7tQ9/J3Gjr8KpQb
vwQsBYaL4nHxKiJ5zT2lwF83I7Paqul4WD0xnIbykUct5E+NXjcsdIcOO+ftSBf4
KSZlX2XWxD2sxz97Xp4Oa5Pv7SKzG/qaZFHsddbmbVY4bkyW9NecdEvWLu5VK5/i
cF6ragGdP+v7KRZJUtgMrooPwqv4RdaY/d5gfx35BuyxTVv3/w6KU6EYzX5gbOME
8KxDjozd7dtYBbraoLWCmFfQHFF4Ukfk8lcbioGqV8O/NXD0VzmkAPrKprv5cre4
1UrUnSQJI6sMHPdhCeM9lVD99Gtb8E5o4B9ezuSWQ07/uqA1JXXXW4MHmEe2DfrN
nOtvPt+7n+W3Z1GXLjvF1FHWJ4XpjV/8HtUY8ZcADrytKnVle9IvzM5SR9HxabSK
tPrXyJpEFl5OL1EWfkVU6p5/iXGtKBQk0MisoN3bdCaH7g6oLCMjv9Fe1WgJVs+O
b80aq9EIK9iCe0QQGFvFZ7XLVLyxRO45V2gUAeIgUB2cItPZXkZDbR5ergxl2+E0
83DRSpjhQuA5neVqtSk6QGybc1kPJbE/GaiyucGrJf7NKjHJF8/Dn2PSjpLX2Nty
LYbox5tX3jacqCIYD9vqR3r0zdVPp1FYBZaZ1Vwg5c966gMTyQUQOoRWa3ar4RQd
64NkrlI03sObTpgLLe/6RNt2ET1EAgOgLhfe1wcP+RenFnWWskSCjL66DLZD6hf7
WVl+5Iuy7/1tVPUsIYAsygSH3r4KpN+RgAeUIxpZNjbLRlWdF2Lo8GYnuteB/b57
9hhA5Py+NiHQbXGmiCUCdxJJibws/pJl2Ydt5QHzA8TAj6CCtZ3LzOxfGfMVlfxM
MdsasxZmAy4Izz5/pzAyFBuEXcNaluHkRlvT++/GsRixv8O4xLp66uZ14p44oXd4
0nUjq17dxc4IffnAc7xzE9xMQjpbpQPk1ej5QgOlDk6QnYZjIIIf9y9yy0C+3EFh
6jhWEGdD9bi6JGCkssC+kuAFQBsjrlaJ0fUejFISNVX53/2Tl6eWV4mc2upzgSpp
cY+2iec6tNoZUqNBp4unHACrdt+o2ePlqjMj7DCmma1OyLykd+GQzAMQoBpsJCiB
YHJXUjlqvZSLzw6fQQ3VpC3CWX6Zizb4klhrCAg/C1iKGiapfF9rWOJWVGl6P3sT
a91FiLWjN1S5xYWg51ddeJ9UvPsIcHSzYk6QuMEykBULPtqMpsXFZXXXrhNwWI9f
AaUAzqPmbPhy6Jj+WCJ18knq5b2gSTQ0cfpTG4f7XTIdAaeci5UvW4n/kxUm4IUb
RFDUmbzX3U4QSaDuriB49ZKRZVxAtmcaXZpzmaFSB2TZiEnsOjjNkgQ0UOKsg73U
UrF30bf8ybuvg1sL8rl/lsDhNpKKNE1SqxMA7nIq2cnqrG3k5+GUEoPPcFhEGvWs
6IxlResT2gwJIYeNh5MAs6p5E/ZDlm3t1IXjgWwDnXxyZ1KjtSKDfqtVOj5K1A3s
nTmccjmxXT1iVu5SDS45tg8Nnk9AniFId8JmgWXFyIK7IJkt84ZQE1r/j/+Afbjb
O0BNPk3Mzu1S2oxF1CEm4kVaCXbgvKtzZP+qsVL6WGv1NN1PmnmFZROC9wQ3nNRs
BaxECdTTVEy0oJfbDHJnpmeoshPShTg3HVRk9W0F5pTReXYHbNJviqOaMTWu3pD4
iR47+xWTEDeSIBrHj88mM9ai+s26L3bQ5tyV95w26pbL16soJNVh8uZ/qxqoamKY
ihfE6kFVa7cZU06rb184pE1CEDkFQ/kDgmAix9fGhz9i1CmHYO8XtsgW5lNtETwk
aDO/5GsGY3o3t10qX3pkuEpDktGwuUs8knsAVWdRZDqgVakGTR044Q8By5CEy9sC
Iqe/WtFgEFyrKihgevMpLYFRAAr7jYXMZ9lHCVzfZrZF4Vdde8fTVAlQwmWMSMTy
eKnsLJ7lEbClnOCQgDrZLhVf9c4Wg8tmk0pQ4P6V425IJD+CVdK9P48iiiuuqGwR
m1YeTmn1Evxp5xVUJYcFmTqgoUMGkCKmc0cOmTBFPtyQu4U0VkZNTS4pZrNgMAoG
EsZUb8uAXz7nsrYmrVIuOqtH54+tzlQy8YYxFxvUdtxq0j/TjcCxm3qRlpSeIdyT
Fw+8g/xeY4OwOSP6Q6TxtXErBH6I7O729oTJBmzcWrQFBqLmVdiEOuSLGnql1Gf4
s97Se6odrQ6ZFQz4OfIFGF11+3bP2qV4YRi8bvoC7PqVYs4kyOwX6CvQJC7SFNw/
1GgC6dt2tqWUhe5ih/ob9+1M92XAc+EYGX0+ZBAFSVJWlwTs+hZmf4MGKfiKKNw8
HkySIrSYvjGaRIkp5WN0G6Wg3tQzaGQodtw5g1iXjGIt0WBJnjLkbh3A+hJ5S1YB
7xMXhMXDMOUoRzqBHoRBPN+o43tRE+gXIce+vrWXpB8PAVqWgKdbvoPFNqBZ/yUy
mlEnZoHDWvCLGWYaYIm2aaaDOvRvjjx8I+xjwA30y7KoQmvB1E7MolVavoQHfeH2
D+fIjcBWtGddV2z6doP616pnSMI3nul8m7ZCGtzSOzSy4uVeMa0M7f0NmW29pIS+
8QZti4Ksxqk5ATMPt0ICVG0amMeDqU0+4QfpfAN6ceNXTJhosFjbGXhuY/BKAkUX
5aRv022RSZeTGu5lKyDAheyFgTbdFs1YxdEzFjSj2p0PdBMxqNWLQEV0EdVotZgt
a3hRWBgAOTsQUnO7CoxEzR5a+GPL1Si9yEoHYjUPw8TZKeMpub0SZXe0rBsiQAmf
LXgcaA1C2WktEcBUJ5UjZoaQkjfITwJoxdQHNNnp+eF3NTkUeSuFkDenaUnQiQQK
jQ7aqFo9am0/MMkNfbs5AAq+fAwdKKIQIUIwD+rgDlYK/VUt1BzkigAXw3jagPXv
3eubQQZQdN4iXGvKaIaYBJMpgnxQBb97VLbkc+XUazhTldZgFs0bFYpoFrytdfih
E3cnPgQmiFwrIMKUp0BirTQum9IZLPdztId1/7UHIR8XoMHmlZiv2q6PEBaJaIyb
JJ232xyXWTW0fwVvvFogiSPfmO73/6o/IokD+6+e6m+DYWEpJ7btCjcWPTQW/aHv
ZN1QmmyFYwG8A4Xa4pR1Q2hwuT+W7I5wUNtIiC6e2SeB0ejjYcOYvnXuUOkCPJTp
suQAAt86/vxIRN766uowT9r9iAHbCQ+PHUAT2dIX4hatsiNLk6ZVN5sguQ5xiQok
9sg/JBYyFzCqA02PmJvdvdpKitE+ixD1QWu5axT5k6sD2H2QyMoEPpGczPBC3oG3
YgG4exr1Bz0Sr3DNoUETX0LnFK3aq7mB0VrKhsdH8aBN7oqjdFvqBmUDwsxQvIFP
T+VPfgAifRMJsuq8LH6+NNKieLPLe8sfNtOMlJQECtBQksPYLvkcjuueWr1ntVRH
QxxoKu2epYkDxsJqVRwngijFngt7fm6jILxIZ1gI7DlWmsqiBbwk5KvwratZez1G
c6NNB6L+z61s94cOXjIsCxigtHkuuitBda+2wqV0kVfDGgni1/TPWdWqXWtI0NAl
Ow22bQc0gQ1FPKYUD+Myg1tRF4DqmIOZqo3Sd2rNqeXXNPDyzYz7oCgnRBEgD/H7
S2mS5kn8Ir5Y+/dHlMKjlHcMUJVSQNk6aY27HiaUnYLjdcjdxho+4J0lulVoMFkw
d6k4B6NrCPg1Na0XCof2EeHIcQZEI6TjzReW/qFWI2GIF5yCHhlhRlJ8MI42eIEg
IjuKhMDvUgIRQ0NnwcA443Ju9bNUZAETNEuPXpAXyWweY5luXySMwa+Qe9+2+8zR
l8qT5aLZ0YlWmdnwH3E0jdsRPFRJR48eQ4zqyBXHeY23IjCVxWSCCHVeSAo/sYco
vPZfR2JlRhVoPFGDxEcyU1Ck+qWdhfsiS8KekRff5UN7mKapAovxhkuzkr/FP8o6
L/cQoXe3AzuxR9haOtUzz8zGiV+M3zDukEt3NaJxyqc/3W/lvJsDr8oGs/RrP3W1
dBNoq4zgu76u5wy3LhSU/dYPwmSD+527YofegafjqZM4HNKrvHOtYHTi9RrNEeIw
TQmOHHP5wZfoVNi0xGihDUqm9qqQGr+Dp7etqx/uumWDGMeneya44JCkWL8vrEVi
QsahRNXQNxow3CU+ccp0HNqjDj0tZmJcRMQydtEEUx6QB62ujvNcH2ut0lsZ5MpR
uVDgsIhcMPLSOArCKnJOXmhBLlPCd4p4+jXoJtXcgitTBIXKRB2/uEpC4jWDltDm
VWgwa/eW28Y7qi+ew8u+IBt8AQ69j4CycXRYFthzGhJd0o9ZR+8ann6vvpk03YOG
DlvQUp/vJ7I2CQJAaWZZ62FfowPqAQvlqWLXHl9S3zakpDht5JeUGiIaqD5j5W7v
Ct+F9rSOLFu2NAgACFQq+XiC7vhErosLStAWrG319o/+US1k+SRhBG3BMZ3QKKWX
6MsdEQfUEVY0v7mpfxcAc/a5XVYfur8JgScBNM2m1Stt9n5Jdz+VCOcGO0ixw0rf
oEcd7//WyMuikmymOWRSh11sIOfXNGiVHobuNS4sBzIlBytoIDfB2D2a4aqaLY4M
qe5aFg9oo4nRaApTpWP6P7a6ceNhB8lzR5mNxNkv0rP4o5kIu+Ehx4cfeb2hwKLt
1PrZv2IOrCuA4w1zhyFPOU47AaMS+G/X/1CXkCNXTC3D9dXWGoo4iy6cgxR5zZ+E
xGITNDhG0HByNaHRTgVEy4PwyE4BlTvanU8qoBi0XGo2ietEzzWBMK/XjMPgvQdk
rgIHZ7gHnG4gpZmhcLnyX1pOYfVciFQaowfCz2i0kVfW/m4yA1HeyMpwti1Tahu4
D1gOKuk7NJ425Kn1j4nOY+Q/etCIaRfDEXWe0cvT4oh1wckgD5txLbHDsoSu+Qma
tvO/lGZTIEeLBwmrZ5D72baBR7CFnCBGVxVbBccwQ5nAGfDymeFC+bijuxuo+LiG
N4sNZ3F3FpSrfBAJI6fJJ7FdjJhpawYW1r45tRY2m20dZLnN/Jybq1qry0y/2p/z
01lTQs3k6EvmILEhxGu0Xo4qW31Wjm4yEMTqWLwsJwhXbI7FBPIRGVLHKLaeF1XN
XLrao2LEYpxautcQMTzN7regEcOt9ITZYBlrmBm4AxqmR/M9cRchSpAPoLCno/Qs
PaMZMpfsk4MjG2mV1ojewRCptESTzWVtn3NfCLYd+6crWMofR0AhNT2zyKKpb1tN
RYDZ7OLlDtZa6WIXwUxsIQEdPsbPqBjfyhQl5lKjFvIyt3a2pJInBiWBv3c55qbS
E1Vvk8yK243o8ZyHoC63GKzaSycbnYyn/S5hmvbeXEH59U136nKO8TRLaKaSXVbf
Y+ZRoXEC4fYiqQcRJD94JWGpxfJmmbAFmdSH96B7VGMlY1fmRlCAtG9M/v6yAg1A
3jQIk8KtGLHYh1mcW/HpVIVIYXbMtXLUIlEj3xpmBEmjeYqAtsHTk1A9tMdeO8CE
xER1zVYB/uPLBzTgWZhldrFThkDbesj5FB886Qm4KoZkF8UFlTp4RW0BWMbCxRm5
OuLgUW/U9gkWJWuz3xFsTIaA+NCcp0/CRHVG0h5miT4bp4YJKJZZRwb6wQeq7T2H
DxOurfQxSdG02poMTwjI6oiM2NfaVooFFrViAcHi2xYdS4+tq7E9wMnfswaQgk5F
RhsfNs2ahuXVIPxkmafZb4X4JrSEmufhwFc+n3NVl6ZpaZj7tHD4zEnvLlClmhGI
YBDxvu3XAdAeFODjipKyC8LMS5PVTZBuYFdCVpG8I8lI3BYAH2JdYwqx1h7RoYZx
6o+tOE0EtdoKxg+briFFJYTzMTbHwwl+WZ3CEpTNhKjvHCOuWM6y1W0aXzkAR5BE
jT3dRw+2f4FBArXpogdvXJD/mCY5kNvrt9Dwk30CHCTO7t1X2F8M8v3JLRDLNLWR
k2pikMrPXCJ3JTIpgXslEQ2Ala4S97OhF/F3o0iky+MwJRXISaV1b/Hngq+MVPV6
YsqMp63+n1TAgoSn7EraMPkAIhFd0cwdCt0O3MexSyxk4YrNp2UpJqMwtTns4DgJ
sqIGhx9YE9MHG6ZupOwpWt+PoySWh1369V6vcPsWoYn3ayU0o4YgJFgGjphOMxGL
erfYDdHOSMcBKrKAm/B2peMrPrNqs0aUjHS2KRgXY9+8uYLovW3zu5MMqwdAA/VS
3/gNi5rRTb8E6zfYVGCN9D8vgp5XqSGm756Qfb0DR/Ury42J7ONlNFMS+zfMgIQt
YnajW2neTgqTeHU8ENLZJ+pKEm1oMN0kt3uqPeVUGNsxJhGyiCvX4jVSI0/L6G7/
dtv3Zw42ZvS02Rt0GO797Dt611ewt5OZN/yKyUUy2BdlTgfVFbbTZOkDNx5F8A+w
YnVgoQ1S+6RpOyJt1nJcaT4SOdP8buTll195NwH9I1MimAlGQw+EGV0g2vrHZj7Y
py/MdUJF8c6/es5DhIslxBxSTqIPFQVzCpQP0KWQZTCnmheBf8UpxsmHxqMoN/bk
o060wZSeM4uz/a69j2vEyiB45uht+DMhmTS5HUSYXZAdkDCAhcb0bSedTjIf6dPB
flbkVhCiLjG66v21pSDE+awcGjSrZxT0oDMEhO6YRf/sLrPcm9dVApoDzbh9RY0a
S0/xPQ7SrtQMEjfDxXX1LfT+QcBOBC/ZRy6GqYTuyP0wZX1DSrqdcGx/muCkDw+O
xy6elaBZV485sgUIJ2zC2BexqBto6ZIx5a54w4/fnkj1oZozMNY1h0SJmF44nQ3k
6+LqXk8ftpBaJEL+W+LoDp0oCPnRMPqa3okmeY2c7gbnjNub6s+Ds2VlOFy0ogXP
lf0yB4oT2W3Q/DTf5BKrbPkEBvQC80QZz1UOMjkvy4GNLdO7lSZCbyZR27xUCV2f
39eg+7TkXheRvUJuyNXAnLdB2PVBXjQYGQo7EdutzgfelhDuEgRRm1ANg0FY9XWt
T6DhhFk63pQjZSCPAnScdHwGnvU85Jbc9MgO8UPyy928B2zhUA2J6IzmUJPR9iR4
dTRwsYzioiPX0njOuNXFkGJOfZNw+Lrp7SiDpAB3Jq1dvd3CYBqNI8gSme3R+n/u
ckCrluFG9uLYCUYdiuVcgoRcbeUXgQrGO3HHf/PULvtM0M9DgnXKs2yhhLwbKdIk
F9FkwUgudONeic26YRmHwL/rWkNoow4OXVpuzVDZ6GoAKiykCfygpqblUH0g28rl
LwPwfBKbIagAfcr2BhxgxNN7A7ifII7Sg6fzvERX28YysFBbIv2mTo8B04wKY7dH
5P9tpHRvhBao4iYL8YUlr57Lie+QPPBe6JtL+cxarDXXB5xRijhcox+E4sEdAxNp
N/sVBaOdz9gGssg81o8n/jRe4UnjjwlMF8Sasg9WHgxJoeb723kDQ7pU/C2czf8N
Sj/+pwDFiWLWkdQkWkA7EFGS8dfxuEWqGTGtd4LOdMj8jCf7Bxh7w3WN3qkayjak
zQ6jGlRtxs785VacJZyp80eYSvvtEhxCAuSjNxZApzqbF+W3eu+UBltcErV3Kukk
sFVL75KdNpKrMjkAZJChkLrWVYwgOaC9ykl+xG+f2jGpM8veqB52quGx+qMjV9ZU
tiB1EKLJCcEj6I1Ji1ydblI0Jj/tJ+8O+C6XLaTuA/tJgCT9K3TfRzeoWr/910mB
QeV7PXYDezprn2STefRS+xTIJAYMpZ1b6blYswymR5wn3xDFtkAwORwJuzIp/HPP
snMVLYu/agWvFqUuQsB/GdwF50Q4ogfWRzHMcw3UCpf8aRJBESlrHcKfrDBRKp03
ET6KPFD+9d24MaifYgPIYV0h+FiaZrHrw/S4QXKhx6PMnvAOD5vPyExdE6PhPuMd
BrwT8v//sh8tGf6SSdGDCFvyIbN54hww/M0hTEsPc5mjMJSnpn4SKlEFWPnjRsDN
JYD+wS2neEZ1NN4wFenMoW7LIF5vfTI7zV7GrilmLfNCbjfphf7De0oy1XyTYSqW
8H9DRSiNht220WILEV8eQseI/X2RH7fEFqbSOVkMEYLQ5l2ubBzaQypPKkG4jgQy
XUZ7tWC3e2e4oFrlqr/vft8266ye+pbXeiTbl3e9VXHHr92f+KjTffqgVT3gryPM
2wmBTmcnf8KEgj8g+9f2MrW8h8IwdjC1trYdXPiq0ZOa7h+4k2mWbVHeFmezUpmz
jM78Ub7qxX1doqgBmwMsw+qaO4B5yx4Ou7nz5zlBMHke/Ji/K9uRZakV3CoNtVWF
2RtcybQD2kS8tvyFJHfjjRZ5jB6p6ZwOvqpYbIfzkpJI5E5kJbqsDLuntk3q8DuP
4cAkfI1yK7Bi4dTgpVfrMC0WEm4oxch5CppnLSCW9WvafNO2331RLaIWhT78yYun
GHn5zZqTW0OTIC7vrrR6+9JIUZBtLC8hgpQMhdsx65pqWP71KGZBN+DD7zb99lzZ
Aj6LCpySisOZb/xZSeqdo46T9YPB70JqWAf7oGj/enEj87yGJZt+vDSGS1eDXBgC
TyTQgHSS+rvxgJqgXR0JMZjZV0QIEBo2CeWOIo+baoJvY3LcHY+PwqHLjkkpQoaq
TCtBBl9q7g9OlqNiQByiuhc5ZKK2dooZHdE4Dyjuyas9CHMHAg2Hy5oyDFTPiIfX
lqLeMcTKnvXlWTxpK/oY7zAJA7dxp2Ty+REg0dmCsL0TxmfqPEDmY8BPgn09GJjs
YlZ9kvSebPvbdA6Vgc/j7N+rxlHPRw8W/a0yOBczChWCh6UEFgUxJDvRgHowxvKV
Uq4CDoNdB2UMq8D3STvb8GDBH2g/aAL3/7Stm0/LuN1iBqmiZM1J6LgtiXj8y+3W
oZ4uckTW1/i5WQd0lQoQV1pk399MFQOBAM2dSW+6l4jTOopT7C9YI5fOrRWCXDW9
5t3Uu7D0lSMivqxHLHO7OHCbPwZiAYpjAOHv5aHTStRZik9eRpCRRP0J1bEVyyVs
riIXA/Kip81Hd+gBwNvtMCFP5KwvMXvJQK24Zsfzfua7cL5IgTbdCVx65J33i0dE
Qp09b/B+1fn2Xrxilm0lG0ZowNIoy37kmWngL34NP0uX5MvpopnGKPxLu36Prj5G
xaeacm8LtLqQjWIig5dKWC3CJBv9LKmUNaz+WiwI7Gg7x+BCuo5aIlVPJwYR8lkb
Wd92p1/S9ILVT/5Ctsb1b6uili1hCQz7J1e4bXeqviVVcOysW+aEY1n/w+sTCUpH
tCOj+x8Y1N6V6RkT7xoA/tUNnUaoaIcC/WMCqMYbvYuxeODJ3QubxDgR6OeGVFz2
wgn+KpW9E4WxVhQNC5YQNlPrfuyhbV8HwRiq1RgBzz7RvvVvAbcPpZIsUhCseJ/O
5zGIFr02Uf4nFRHwtBPqyVgh/6v5AFPA3Lu4HEMKXxwsEyAyvj4sqxkHa1OGhOgU
OJtV/ArHE3/vg/U4/ziG1YFTLxkRWLDpEomgoCB+iQyDF7iTorChTrqa36NXbMMp
7V7i3gao7oeSDmwAs9pIj8K2fYI7XksopSvRo6/SIDBWhDaUSki4dzu5/IZS9r1V
Q7KfaeBBMz5R9SJLk/24uXmkneDxma53VucXV8mFkNms6g/MvI3pRy27QtFasOcx
cAhwo6sAxQSYsY8Dktb0WNfltUXyaMM/uDzmecl5yQqfjgew2H+d8fwn4ObGOmpx
XrkKl8N6cczNya09ueMb3yevih+wbjOKA8dX233ieM/OcaPpwtS7MUVvA5gU4iyI
m3pA0Afr5icdCnJNIuQIDb+MS0NjyW/vbsTmAlsy4iUtt3Y9E/jO85wjWW8ZdrRZ
q1KkXM5L3pd2t5fg56PnrPAZ5NOdHouInM1yQMKtZdx0/KFOn0vtdw3PsTOx6Z6+
xXHBJgj6StCOGSJ4Q6+YiJ9fX/+dvzNTuXckxW84hM3vup4cjrG8SRL2syky0LIG
aMXSPA3PGgRJoZfq34UJIvAyaaw9roo331KrR6qDFdkWqivB3maS53OAvGYvlYO4
2k31zDEZdf1FRCYRV7xmd/w9Ct+JJ3CX+b0XqKZMpjz6TObV49CflV1JmMQkfuvB
eacqWckc1AoH+J+FAlr8wcdIq27eWqCvF6IkhJmO7byVohOT7oplnfsNEbfzHapH
8pPG9SLICsRu4QccUxwUoU6v6ltX9KctMBHqVIYoQShyYMskO90dkJEsL82auZ52
rL0HCU7AtFlooT95bVHduh7KKjp+/Ndtdt7eZd47j4B0Exu+ZMIxcXzM3BpV3XSF
fR31J1kPw4amoUf/lVxlLz5rpRYNLTKbNcsEXhXJ76kzcu8kSrAP16rRRSCc1ydT
A/ffNbbITMi55VWHpIh2Ie2Z5werBesrLROSKzVIbH/rBtmf/UQ/+mysHCQd0ZgY
9r3wUA1JfJaR7ng/tgXqZcPdyddo1ExUfIpu7JbmKdwXABpfnjWvGbB1Fl0koQ7P
qW9so7d2ASGZFB0wNOM86ZKipteTlsy/H0hG6MmcZt2i+GUkKduZXjqYQ3GhfLAJ
mkFm708Fqr8qR8o39vRM+5fc4k0/CKV17SgNEeukDg/lr5BF5i2E57wbgA3tEUsy
QYHe8pVmvIIbLR0MYaCEC4YH5J9zmc4Tq0+qdgx10znLP2C5mURbtox62TZlZ0fX
25i7xJownCuc5eEVVJDr0DZqMsWE9elWPpeK9iURgsWJP7e3jfTa2V51OJSqekVo
mNPAiNTLmcIQZmbgokrKQF5B0xVtQ+xDurYMiQK1wcApRXSktGY8ARHoPPvaaCea
ScLNj1ie4aHhPjWyFUEsLzjwUjgRJq4RL122GKFgqUr65D0wzv6cht04AyJeObA6
SotrXMKkPNv4ghq3JhNphYoYE8oElGKZG12d41+/dlCNoco3sLjM1VpNSdWs5WWd
T2f5zw9Ekbfr6mjUJCh06ho5gV21taVWZ64+wQGWwEJ4msv5h3nWGnfL47Ieh2Gc
T6s8sBfm4H30EvqpnqrnYA5yiSKQemnciYuvNi5iCbJPsjPXEzpB6pW2CM9gvSsf
3yIv0qE7oR43J9MxiuKwdQOmv42YUqTWYW3yxXr7PUPxi2YefK3zP76jBigwg5qT
8oV21BC+iZ9HQFxAwELwVcgIBHb3jggft2R+hkWjRTjNhsIS6bnZ9DSqPAg7BGRZ
3mVUHXSDxl1GSJZALvbpwei2BNOf3zFDnkbCSnR1vvKSAa9ezsY4mGt9xlZQY2Tq
4ta64B50N7aCZ3q0HeEz3ACDjSdYPOoYCHoejxjpa3eGcKqjWdq2N3v/GZcNst31
I48oQo57EtekdZOJ6/VkqsC1qTP5kS3M5pvHhQzAf0U4F0MpTiDnSqdz2ytovOSJ
2AgpVn+o+WHNObI1Cv3aeNFqA+a/KgurIayA8ircQcGJL2k1VLk1frFzdc7QPMzi
Ftai8V254umGBteRvFlPzFW6onSTUJ3DAKm47K4g7axNGWjLDAT/w5ZjRk4uaohQ
YXYBTjt4GG6+IHu9z1xAZJBpyT6rDXS03RTuxh0ykkHpR5fwn0VLPM5AAnWUlJDk
HVClBRB2BsGbpwIkbrJqimh0b3LAv+GkYxTJ1jokaP7hke8thVlGBcHpEXCJtUHN
gOTDkvXScPS6MnFFa/QRm9wcs4i8Yc7oDvJgFkCmPR/H4XX5o6xg0JXwwJGYoJWO
wD8SuL86S/s4+CARrZ45sX/Cmp5l6xPJePpnP41WLWJ3zodCwanJSVHz4WbX5FWy
w+EgeXY5gCwWEezrrvMDyfa3kPZfOmVh4ZviYU2J6YXquVNeyLnsHf9dtu/hQJNH
Wi+1kVQKxEGE3T/ch/UxR8kNQ+PXRiG54Eiax6jwlbSqh5NB1q7Tsr6Wczo/ID26
QIE/m25M09f5gY3WeTzvxe9ZYfM9DdO6i4IbDE5boeDU6D+9CSCtBKlPSQs484m1
C1j1uvIZBYJ10gPCzXiIC1joM3o2OobGLUL+zZW8oM3tHI97TKj+KU5v7hWR8VZD
AwQtXaVj2nLSug1G2b8xLqj/epLGFa8hrCmJYG20iL8/6Ta7EXjaQKjbgtQPmzDX
UEJVBaM0f7TClfqIEzF4BPTIPm5KKGcLZWg+eWoxQ8a644bGrJiGTbCfh8EIoj7U
9AgaeGnw98T3KvVw4+ln76VMsqrBN58RG5bNxx9YDeSaS4u7wWipk/Pw0LiH+Vgp
fnaWQzsWUVpX9bxZ7HSIORfE7cEXR6oqKZvw+iYQSTHjgeyWD8ikZkaKz79DGwBz
BW4lK9SVQ/uHowP1/mpAZ/5ZfgNj9VhV4ToykRPX0NUc98+L+6YQ+b5UeKlj5Ps8
kmAtIgZzdEqobSOL900YUBY9oqbu2Zd9oPZF5MfirpKWU+ievZpPMaOiL/awGs70
KiA8bQVeAIomF5P9QDq4HxALV2ZENKG+inBuWQbvzRm2TFxlB2MyoHOdV/Ych/pP
cudqpY1Hhyh0LkJjRlr9NzTkmGnEEFnHUuY7vP8MKE3uRwAX0DvIYKkNH4Iqu3r4
cNSUWVojI72JoGxsRao/s70icnWTfEN5zP/JGYcV60Q98HiXUoXsWAzs+7TlDNkb
/m/eapXCStjCiD47vsJKJfE0jdA8gEYe7dLzvLYu+EueXdSRlShPAsr7Esn0G++v
d3KihFtvnBukATgbfBqsXdBqNLnrVSZVo+bewD2YgwhiQI3j/vxm5D0NXhOG4aO4
ISdQW/WphtwlqB2IeAwKVgs8SdfGc4K6LrQgz2gbv6xyYY86fe8owZGgylON96mq
8Ggb3v776QKsVGz7VXei6VCEqXRlBTWTj/CIdfYrOD1DOp3mF3Z8QOByMz/N0NL0
Aa41zrYbLSgLdilSDnF7850t6u7rWyPKJnUFEAwaqPY5s4kWA0Sjpk+Bl5WAcQ5d
iUNaisgl+BkWQpPLVnu9/bIhns3pij+WR880jkytG6VM4cTbv+tJLeMulBERfG33
HgqJK4bxW5hH9UHhuL5tW2SLvvfl2u84kj40KiIYpvNIs3Hx0f3NT/N85mbloBER
Fa2R0mh42emsAySnqyKqKeyxkbsRUiZVIhGA/hYMk+16seBCsmaX28IL+hicGn76
>>>>>>> main
`protect end_protected