`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 43504 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
5VZyab7crLRA+ZD+A50QcwtKhwHTM4ksT7LVvdUSL44Jy7vqXOKh9RQPT1ji19IX
TZAW3x5aKP/ZPv8PS3ySFiFPpCUZGK2/Ke5ZKo++HF/uAEXyu73MwohWi+M+/Pwi
r5XiU35g5kbDOxeQl2EaH9suDNwDivhzqSUmmR4rz10dsDQu5gP5UEwru9tvBX7Q
d9BeMNZCOcZSo1cCzHyZhTD9z+rXxIogJMDBiV+V21KDyIZ3kkS9yu5bI9U7Tmhj
lV1dQZEMdxQyvcvTwQlO9dwLs/jM/yN13hYiY+MNjD9zj4AZK+2DVECaFGI3k9U7
m9jg3OJqK+EbtgrF+lxOfr9fcl7DmSwj/hoL1yxmoaIskvc6c03NrmBSySXakjGs
pXA3ZxcDkWHENQDiswNGxr6rfgzYIxqdTwTWR6JlLsXl4rS5xf1nlVgyBYfpvl7H
u4mx9zgMQfKpOeT/mnefHulHnUP3KkkrpbIp5z03DMfO2CJ3xqVlDClx8TXm82gz
A6guQtNjwnJFwacw+UUzTH6nC2I9t8bvzmPjmJ9fzloW3Ioeg/NWuFPDUDEyW2C1
vKgvnOXnsD1rrXOmjMqxO+QHvzi6dUku76MFw96Zm5eI31nhb9QUo7e07TFTFnr3
qKNf1Xe2gOsNlWW4eX5AqqR7C7YD4B/joJu0/tHAUHlyd6cuD1U6BWT2CzTsSsgm
1SqtW9twHeBpNAlTT/ZNsnGw/v07q6Dbblwo+GE+6UUctUOjLm2gHOuqAA/85zEz
TEVSe4HSbyrD48zDwJQo+AnJDt6XKKk44Rd9bz/4JKM3Z6tfg7znJNRHhCuNPKP1
ZE4MskAUYT7WH7OxBO14Mccdrrc2c5LMzhn8tVNjpTj4gHNAsaYfn5pkHJRwhLbx
lyyh2LwqH9lAPCv6SRq3TaSBXOCr2S2kZ25m5IFnQ1wjF8uLaLYppNQg0S0NJLzc
6blrpu17v92tzk20TA9oT/mjLyu8EygZq/pZmELXE9GQuIPq+oz4Q+ixculoVZM/
KF2ZJRmXP37D+/VEtOylH9OHFRiCnONefnpgDjFLNYY11Mu4mSU/c6rjMH+oMqsH
zUP7AU6auYzP+XRHMQk2lyRzz/wdi7wl90a21sEqu9DojWZTYBXzKGxLjbRB0cSG
iwBKOjy5cBIzcuCbCEsCo4BBJ8OtLAUbZfi++qdSTuzBjAYPtgUyth+Ou6dHCImV
8loUF+cWERPetZRyHFqO21LMvw1qsDyQAJHcMkDPO8HZgmlUmq13CprFXUKS+QiE
PJsPV9GAXslwR+nNgv+EdvA5vaz+tFgQNRtmF0SsvRxFBOvlNUcyQU5VsAhsMGoe
RrONy3Z77U6UoSsuU8XLSsC4KIcVq1hC9rVii9QTA1KRVa14b+b0QTbN0Eh604s5
eRjrHqDjWuD5T7nww+woSYoUleiLi8yuK++7w5+5FLitKGdSp0+yST/KvA7vXrAb
xdChGPIig1p2wY8ylto1A8BxhOFImJwtGnMK8taTjYyFVkirYPjq5jm33nm5ffeg
QaTyEZXn/hrIUEVbvyJlsR/N8Px6v5pkB+RzdvGNese8Tjug6m2A15YvULFpbEY1
sjQngJnvaxUy0E5N4ByUBePPm63T36WaP1A2FQFb1r+Z7RG/Vg90Z+Yx42eWh02V
/YupYK0COwAKkK4lrGHAtitZBGkUqx3dckbQ1UI+F6RZYOifxJUuQP9VXQVkA9Me
8WB5h2AyH+ysxwvMuvqauQYYHMTwG6NPgCEpnOFCr/XQ4bJnYBuh89+MPC1EBJ4R
QGog73Lq5NjjhtCoVYWc7iALoz7B58HD6VqSHswmzqedyEICx2Gb1zRN11fECyFD
LBRcOUt6HKD1tGoL0tXmU8YeZrKtnK2496YwA4DqfTlaDuosrvoJK3x4LHfdNOSk
JwY1/s+mhj5Pk8MNnHVtR8bRImRWZxnKcXSmjGo4a2rB/Wm3YrVuGDw+4tU9/YL/
x2HLtEaOnli4Q4Y2M9Xhw44Rt+bboirSr8GsesE2mOeH71B8FdhWD7UY2XZNgPEE
mTsH83MniaI5riT8Q/NQhUaPAZANUgvYk8asXFjzKJgfmoX/zGxd7AfyMwfjZCdr
eXyczcRtoUNnzsF/uWUBGLWy6tk9zH5SftGOzgk8pDYxJQiJS4rRt1WkvymBsMrH
JtXf1M8xfBcvWDdYczNXrHrKTGZQT9Vp7hQ6tfxnqHbRrI9AXlOS1MWtFwhzwkE1
1+V/dPdiqrXxYTltfCNJA696ImYQqCV9mVAOqm7DjdbptzogBvu9iLzlXAu9poOV
l2YEnbQB3q344gb31ET7yXiaJEYdsgUfRYpKJi0IRLLIlrFDUmMnYXSV+Hz1vCEo
3YbINa8sphDOByl2QGM6kjNqmSNEkaQx2IfT++NiMONUg8GihOPrGhmBz8ytKIR4
hmRn/LcUAiPZQ+A0LbPkzjldyC4PUrimMxctQToHoqqa/NUTiyqYTHtHDkNDkECF
djLSumQLLvR7tqu9zgdOfV8QUsb12t6KX0pxaHRM7mplK/ELyg5NqQRbHarV5/Ez
YzaD7V/RuFnUWBU2dsyVL9p5Tgp7AzjlbRl2QIvVr7b1/HDIQKbTiXYVg1oYRmiM
O0v6TavDzbVPkWf0bDfZLY4TLthQGH030RWEWE+FQbvoz2xSh13fAfmc17QvAIIE
dFB/MPoyqCP8Ar++br/H9zKwUqo/jJwvGbjkA0ShN6UiTE6Z/Ewq4yZXyl6LQxZ8
X6xdIn8gdFNyvh/htnBTh/5LEY7fcNDsJiP3evbtzFk9+MB0BAK/eZaCkJ3Kd8X8
c2/LvGHZWkmKD7XN0ZJMJ8+an15Vh7HsBkkV0O7l0nPCpIGtqouzl76TlgjZCKvz
Se0+nY/VFYUvojXUsL8vDS+/Hjvf0TBnV5Yflg8OtZ05UKQAuKGAPnIdpA21qYo3
xVPsxQVLlNxfbQWyBo7tNlv676H7N8dTLsYWgxISAVvz/n0YuAdkZneMxIGDCrO+
jK0s15SszeCP0HBhAKqE7igPSdqIHDOao3GwMQbcG9oGJqoNmOr64Y+juU1rJnyP
SKrcITY+3Slj00j50nFT4JCq2X+z0MSM6P+ROc3VmsSn6LO/9/lyNcwngA0CR57x
2Wokq3Kbn+nV8jHp4NIUTmsXqIxf27OrOI3YTlCqcDSYw0IjkYoxVWQjpVi+Ypm9
IrGRrwXQQzGTytzfKObw9FTIfK4z68VoBJZybRkq6HYhuNJWJF5VbIOoZjMKfd/l
lWRnWeJ0qCCb1mgJRFlDdp2rEniLLVnEOpv5uZ5FkpEpATcnUFcFrgwBTwU/AotT
nE0ey447UJl6f5EzM51smQkXK6mXrs3LSv5I8Zxfbta0RLfIMFIeBsK7NPQbyBZL
N68UARicu61951MOQHq29ycEecu2tvV6DqSd5nBJxZ/oMoGnkiwvAnBddje0z7IM
tPyT+MWrj0++qAPOb0+oLrTG0lWb+0Z4KXtRRZW/q2BuCrhZTtc5u1gFwF2SXINq
AMe+kF0OGUPls6p5wZ9kykWDsva/j5pG7XlJQOys5vdlKP/M9gBF8ZZWxzikyCLH
y6V7rfoJDwD3jmlrHAvWQ1vLCSuGYzDz1/IL8ClfUiD/qgMZV4s4EEPDKO/GVdRw
DgunuVb5r3aGlGa+mmy2oOWDHWlhWIRkqExGB6vdft+REN6MDvkv1IcytN14VL01
yJeUCVpkgwF2k2xfO+12FYhaGOMkiFVgOsySEfKCdXtSqvtTYVNVoPEiVAlAr8uD
mOgIcvRbxlOtx89u4CYnkpJeLwT4uhOLh8eylvmwv5S+jLPCOwhYynndbYiqHQ1M
DoqVQGYLTBolgTsw1W/DDCRCIWMXdRoPFLgAQ/XkRCnZte8xRTNo+dkrVvh41/pR
lKOmc43e0DVyE6BTpAd190OZwqa0VWv0GvZuoqHu4BPO1gKc29P4ttF10kRW4FYy
djaKPrZB/y1APl0TZNyXoxAB46W4S523c2ld5kJuumyCtd3VuaN10aX3K4zro8ju
hhO8Yy3IyohjVBdfDwNfJoWSnoUgolfYZr9uYmgQWPQZG9gKJBkVkeSm7SqqfiPG
IjVbFu/I1qKQr17qxIWDGL9NZZTcUsub4UowxCGecjNm87JjnlJpahCyqb7OioBh
Sj5va8FqQRSNKn/fKnZ0HQWxKG/RGKd2Qyjs8Mdpv3inoxnPNT0duhKedhumV3Sv
HKqBpABsPTtbbcLD8zVUITgq/akk5FmxGTzhQ5z3RtFkLnV2txZFnBdK9CIiQD/i
lRS9uuHuTn7jmJhPuJQS7JZDAUbPw6g7v6Yddwj9Sp70rTSDqNv8UxepbO4idbVi
bPzzcAQoTDejaHbzVdQuBsCVQm0w56YnoPMcVfR4JAQSrw77meiV9ZY/tc7JsvHr
9tElSPwH50THdN80mT6mYl/fZ/PoFaKdnIDcNgodixfJapJMSwROfXl/dothkemq
pLDd/r4htSPmNVRTs4NQv03lnTs/Rf5xI1y4YI/czMohtVx9vbLQS8BIs0Wznwui
3s7BRC10hiH7HG8Zo2W5/XXr3Ot+6p1s3nX0LsxZBTwcyWvSKHPuiAkVfBnNb342
1kOOUh3A2azqATRjhewO0IGTFTQKnM2yg1/aOv30qtIK5D4CLjDbtXVpCoBDUhay
+pIrcf/ULuU6yS2GOrQM6uhH/o9FEbpeKAfS/qHDZNfHDcAvworaIz0MLVDAC41N
TWRGUBjbAxXXh4ucNtucY6cNScM1vAnHrD+zQ4COrRuQT27uITl+svsvExKOVrfL
maxOSM+8YsbW1xsYv8MAFX7rrFfdppyWsIHAtXoIjmdb1QMOs6THMLGmRaklaJc4
ynailPleERusFkoJgn6UEEKdmI/8T0j9zmqUGIppYMuUZB+mXMz2UEDnPnIaI8mW
ahXv7oDhSXDg309KRAtjr6hH6Ym88gr0pVJF5kovac1kYqb4zZrBOZ1iu5XL16Oh
WjOV+m+Y7sdt5N+QAqc1KtX1+o1aJEkUo4lJwycWCKcGWDOdRvKv/a8zuFA0F7an
eJh4bKjlJHsgbKhciFevOuYOBtxc1MIXY2/xqYSRKupVePZfdd/FbuWwfH091vH7
p45vylh66iRJbeYXadLv5QgIXa3PkqFPHSacccKlx2rkBnccelOIIKQlIdumakRD
8ILzco2fHaS6faVniMG1nGV9WG2eV5qFIYaZAupDI4H148mMcncz2p+fnj8Rz4sw
lhnkQjilA2OCNmXDp0iBylzuzuiLRuHM31XoQNs6C+YawhJdnjLJaKZVvxRdx/9C
COGEo+PEBXJSUNHgXsCI93aHg8US54sNIxRGJdWuEu4EL2LrADkV/t9n+LCkm6eA
qPkOl5n5l31EWhjAECE8x6QiT7nJS9pk6W2ngQcqfHC1tc7m4Z5rkvKi7Pcg2mKv
iEpUl0ptdcKeyjyZFzu0B/ItuGRnLzSIJDehgkSFnpVa+5lTyDPgmbOZWl4KXQvQ
XSmZNxbi7dCpMg3qYIMzJ8lGYr91nImFqopUSXF7EGEzSISszCH4KeCJCMu8Za6z
6w6LboXgZCPXQ5AZr1x29vGYDdSbqNWirNJaaA7p5cL6yJVnGxuzICVXfzJuRvvZ
KZ9k/orDmcN0Y4X7ZyXEm+kM3qQFVltuCnERxCCPJcHfrp4GBS4heTx7W4Eudcw0
1NdnYYRyinvCvDxrIk7Wv043i3y7VEodP95nBrPqL6LoB2ww+RjREXKQ1dI95mVt
3tpEcGaSjowKt3wA559YiFTWe6zhTtI5Raf7cQNuPEqj7i6iBOeWVwAOr0CfzxzZ
OZdSHjbjfR9Sqjr2Bd/fYCUbLEjCzwASVgtf+9IPJg5kpSwFMMc3cvIgHOOWt/7S
Ly1/psIQTpZUTziNbWQwB+MyGPWee1rJsp4q+v7D5EY9n0dkUITFa8Gy15O67qVi
v7ZvM/Ip89IlxiAB6GHaIMczfSgozxdNHca7rN21fFOI1pxL2Mjubwy7qxj2jK9X
bLyAywUwcu4Dc3XubUZzF7Saf9+QPthm+0qTdfO1aTPMPdoeJINCJMmWGbSggBVz
hCsi2ljZqpU7dzZcvO1bKZNq70NJqB7NSTUq1IP1/1QtJ2CqNTaFijqyFlrhlIHO
2lt+jICQDnFn/mLe7LbrGsSuM27KuR/1uMeaixmSna2hOAnwnZUEGOS0S0fj8JW3
kMNk2JkgZuloUXAxFexuuvrpqHH38Ljdj6pMr/M7RVH4YpCkk5s1sq8NSBH9Yd2z
MzmltOMPRnNykjrtM/k42kOCdYkALHta/Ngzz/U4OaRnFrO7ji26HGZHw1RtdOUm
S2YTHpVEGBYfbIet3f8BV3yGqoRONFwn3SQ5ykz+31iXZ0A42dq8m+q53+7wmuL1
qxr7QMkAqV0JYjDea6RonJsWrI+d1xk8GQrMKQtqX6YaF1jAQxixqUJRNAngXvAU
cSOIzcG0wPZJjk7VAld+y+whkU2kFuRrC5mZhxWgq12+OFiqIG+V1wW0aRwJPMqT
NolNKudCBgwzVFEoHtVfZiU65L5b3VSco8gnoz2F/OhGUOIXcPO4MwQeBlD+zN7A
itPVOPA0/tze4vqbT+TfKpQbtzYdOlFdjgYdGRY7W/ogEcbh03a/dZU9te9FK4TJ
RZyEyJiyiR5ZUr68rYv/J6v9hW6Sj+SdbcfaZjC1Q0W4qDBaeNwaIn0/827urJtR
wydHlM/3MF9qLjZiXeZKVaTBvlCMh+cyFlRwP5dYmY7HeCODgEm6LVlCNKSE1q2z
i/82eBhlCDLmr+Y7bGLQzYTZON5Hw88+WYd2x4lBpFkbayLmrauvqfMnwdK6tJKE
J0G0Gvtu38VOiQVqHR1nwVb1G5bT6tf7ijUkHSgcfzlMakPsyAMV23RihNMqneDm
dVr38IDY0z8nsUpI9wz/NBBjQs6mvELdIr4B/Y6lk46ayBaKyHctW9st6aPYTvAP
ev3nIcjsdzxpi92K01lahzl9zn3qddoNwYCax95zuZ0eRBAFMeiOAHYLBFlCiK1b
6os5sYKjTSTaLshkR/CFX7KRhIt+i5xz9qXRF0nXlLBTyrpdIvuLZi2jYTqsoaPf
vpcrEuUDnXzIpVRg7jbVZiNWAsk72XA84/ZL/C+pgYRhDJpcTCyfOIM3T0UH7Tsq
jeNAhkxQQgL0r/dIs/E7uH1MYKXAcS0icF6YGTQEhWxjwgExlF56skFkYWK9V2F6
uvPZiUepzOxstcEPmbdSjj5Wv+IJFLyhwIxTwHECMs/x8KZr9ntg4Z9jRlZJFGHJ
W/uJ5ZpnQcFM7UOUrN8OdzyCpzLUfnWZvsiBJuYMAaLpwljYTRdhOWWUSTG90tjk
gxux3RB906PS/rM5HlcWJJlG6WBiMIOeHCzrjGlf9Xwhmw1mtjJa0PMA8k2FBRVz
RRSD6yIzQ5RvSFKJU9LemqrEqOPRHITAsLAwcPs9F+Rhep56TD+DvxT332ADFbDe
lnzvX39BawbuZILZoMlhzL8PeOwGOrCWhdB+sLc/r6YDzzHO9DmtXudKUfl4FzTE
oFgO0y5Lopfj4wLOwFWPTWlYG3sYI4r8x1goXjTlREzwbU1cwiR/gq26Ket4+8Kk
a84OApAxexOM75ssxU5YY8Q06A4gTfz+zFDcVSTWhdI9oOUdXvHobVKPz9/pvAz+
zEw833LUvKjS8JLB2hY2sfdnyA08fXyjsI8qhCbkH/ozKh4KTuftY5W6rbj9vCQi
Y1rzgBp27dvi58zAGtjYmo0nSmF9YKqNuGQg2bQr0GiRhruM4IOV70kJbsNbLpRt
f63W55NSBwacd7oUs54JZNO5xlCZVCMyZ4X/EzL3fwC8uFP+aQCoorUz1+htNcqY
7HDZ13+jDKgDtGVGx+q3mrs5hfzunIs7tNyCcoUt7AfvmZdgSfn5+xDBP5JXd+L7
/WA7VJLfcD+dFSH7/BaR5Kgnr53DAArB6lhTxYlsAK+CxZykHMdB7FXhG0yaxg2C
aWSre3GkzbQPWGo5RjsrjosOUw9aAijFE3+jcuW7ehbyjaoqXxYdaJcpE8yVd+4J
ww7CxLSuizM/z2upHrkdhjHJhWZSFvGfl61WOz56ioo9MlIAkibtvJk2ihZrG0/L
sKrPErXf99Ilfow5YmV1HoNArFKwbaNw5TfWOqRkzZf+065183LpPLGsknytydBn
rgYPmAN2xXcwp5gd++q/m6ZcOZTH7ouZL+lXPjCJSf7tTmWEEG075LS/F462p8hU
CJRCDO2qj9aRxMwH44xdlsivRQIIEnJbTBbTde7o3vZ4txRB+H8GaWc2UHjs9bsP
hY1wJsVuwmwIK5OFO2uahAmmk+uzsKYcJIg99oxXOvHbQrXqGduOizYX80qiXyLy
HqTRa9MZwgR0TJguruZHR9h9FqKmx2uJoP+6aBbzvwBSY5+6hZkMRD8k6zk+WmsO
Jrdto9rdfJtEDVnvzpoarf4dn0dup/+jQfFWoZcaNq9hZdMhudsB7YfIsmkFf5o4
EwjQDzgWWxjn6Tuk64bw9Uof03NqZUSDrXyMF3foocQ62g9iXLM0FPcKyBAKJs83
i0IWpFwC5BMerFBDqeoIf1dI1F3m7SPWmRiuolJE9BXB2LYr7vQekbYW3Y63ZRB5
y5dpTCqiM3sTatPTGFcWdhD0p6C2sNUtbrYkr+l8G0curd8Ykz5yfTBwHE/6Q1lR
F8Q4uMeMZeH5Z+x3HM8Z6Ldc+JGZHp29x2pAT/ps0XycJtt7jBmNdudVLSP3939p
JotjJv/6npP4cIMAhcGNgLk2bYrTYRYykT3Cv4MTWAB+6NgQ4PJ0LedjcuSRqcdq
W6Vt7D8NGWnU8rvuKvpNHjC52ItYPXx8ZOF3NZK0P5co4XuXuIAIvw9V9kVkVjsm
iRnvlGr177Ans4GVmdg3OT+Q5vN3R3DRgYmedqefCeKtuunR8IcvasJnMQRnMBuS
HV2b3zvuQ7jVIoUdtsm+VaM4IMnwsDvD8DO8jWRnkS5hQSckXgfwnE47JGZrU4fP
GLQUu1GXDAqy35bSUYUhyA0nh0fb82c/AVziXP8JFsbnauzTplhUpmK+lIVEv9V/
DbDimXqNiGkVCkd5nJZGbQb2hz8BdGHDv2W8uAWu0kaRjaO8kmFQxzCsmCKB9gEf
Bt4NVC/4TyJiqzFFuLSmaDKSs3qYLViPiaS1lPBFiTsrEPkcZzPAL3MIJXNIkVbC
4GWv/OWIOYN6gwBcQnyQEivL1Oy0ShG/9METP7t84ZqEugJ9HKN8wddhjPefRGFK
2rQ7aELUTWSXw4KsG7CYojqUdLEFAO+9z5EBfnQin1RZVd7Zai0LKXs+MA9LYFYN
mb5syImt+ujzCPOQQFjzEIeHcF2hSIFDqIyGaSQvy/dO9NVviV9Mo4C/SsIIlMTp
AqNxtzNTqymqPkucqZaD1tQIvXc5B72VzIHyD6vZ7Ekhxx3VetZYh0HV4ulnatIV
6agSULHVjlFRfhThMoTZ+owxWgJFuZdz2stpZiL3pqEb/pov1Jol39eSV0gUcjmp
rCIJde6BWu/9uwPkzeZNt9jh87SaM8FWw0HRbXVMAgkU6iVl9DZhh99lj1zxAcMi
ypYbSs+gVwmMw1baOatigFLi0dEvICuA6jzVSgW0ReL3/PYJ+qwXOnrWSdRNd2ns
r2vRlHxz8a4p4AVb5ORm+Vu3s9TAlFxhSiHqRw5414kKwEpMGUfzww82+sDBxJlO
xDtQeFW8xawT0JA86K4bv+LXzz2dxtdu6GpskQJjI+qbQtxOhiXkdXx7JsMdkWHz
bgifFTYZDNYzDKMUAw9IMVZWkjcuLSvSr61klvboVimkaFkI5sNesJnSczaoLyDN
cvL1m/hqtn87jOkomglZyNueEnK/Wp9CSvhxtqBInAyP1tU3ujKJ+MG2Yw1P2GSu
gXZRB/xX1uhyBJHOhaBOkPQK9OTW3ynfJtx5H9JH8NenHCt4BJQB9ZRExaJFvkBp
aUDOQKgFd+GcIz048CoqWY/VNvlD0kFY0MFSIrnMG+AMJfUf8YvhCyJErxfSzujp
X/QZiBs1iYlRy3s3F0GrzJXBkvQA4Xv4GThmuc/sAJMXgyHFfFaRt9DZSXnR96cX
MnLsScBMj7eOsCYfUa8F+/fTK85Rvflxj7gJyRnhe5VnrhFaQaqes7KPml9dL9IR
dqU+e26SrlClrGdfp0Kkwzaffedt+HXQ2ydbG9hvCQ9sl+ok/jmEfsf0uJ0rG3oM
Yt5xBX7C93zQTCb5rV8R71yk9o31C25P1FCbCZOTYL/m3eUupY409ctkRpJyzFIs
O7UmE3bXpNlBG9eXp/aAq4aMsnOuvlO94bEslSBQRc9gB6JwNFDGkiqXhqVanm+Q
NyfQvW1ALd73UgjaCl/4llSZNwTa51NlRby4w9w5ffG9dqC/nhnzfL41ZsTQPUer
Hl2cD6nYkr5ntMaORC8DfCcJ0F5+SErRVnZ6zYVMQLb7d1er8vn1CdmqNBSI1xcl
yt+5vGMwOr7Go6BaBlQeTjs/GPxU09aMHjXR2CCniIbVfQV5nYWoeeMOoJC4uUwY
0GaLxqte+ma1cn4H9FT2EGpMzPZvOgBtAkMeJXH0GZ+Pg4ad9iKHQq/edfTqzB+R
Sb8kB+BEj7/31aiGq9qDISXWEnd39bkZRRHkExm4yFhSqyRJ8Qnus12WRX5ITB75
icINoOKF2Yh/fE34Xc6Ed+wLykoxzy920cP5YC7HLSaFBjk1zrAvXlRLU7az5i+p
EvalGZQXdePLJHT0zrsQ7ws0SWpmZ/nO+6zvo+cweBdvChaBOzZoq3ZBNBMl6Qg0
BpmQWTJcjtuL45lUHtVbtjOMFHm9K3h4+Uhguon4bsvmdoR19W4EsV1YXjVzxCgo
I9cobhZDqzA/WsA2Td40wQMkYz7vIFB8W1A8vTA5jC+2rSqxDeDBotWwzav3wypu
x0dkhPag+ISN+Ig52h+fA+eHmo1YCdPELp8r1UdqQWxg3CGVTgLb/zkwuTaAHn6y
CKhT5s1Xsa2lpGrrRaggyx0E7qhN/A0zZ8D8Ojo/RaWwGyDaasLp4H8H8UHNvj6d
rnOzW914X6TG1h3DgH/RzxnfZMDnaJniLSu6qnJbZbMTXZKM5aIhHUe84rfZ+8bI
nVr/seu8WCA1NVCEAcM9T9wTE8M8CsuZ9bSLIiWRBkIZCUCYPx9OUdu774+qvRnc
11mmpjLU0hYQD/jajNpD2l+QynkEOhhyGkzhDuhDyqdEdk4svMtGkHTAl0vi3Idz
BcCEGL//+qXIwD+JpEz8YYThZpMOKqj36X64qsM871pU+Zns14P9OyvQN6dpv3mb
mGG0FlOrJz83Hvl2yHlPRPe4HafdUIU/ar8TNbzahkUINwq06zaMF/Vx7CtlYdvt
dAiQTmGenIWZMAq7hsJbfKCjOKfewXtvPU/dER3wPWmrkk/g+KJ8VSzVl5VS6eGf
4Eatp0dZW+2HZKyLVI4RRNfRu3soH6FPDrN4+sHIbBvY4KojjkaR+/6RTWMiFJd7
t+I09JJD3VCicl9HpGCpHSPsHT433PIH2mEGLLd3J+0OqK95OAS3N94KaOsWRUSX
Gn3zhXCu9EXoAd1fjBY6vxXTkv1Ar6+HOnz6uW3p6fZuia5jJ2JKRlcNkWXSFATu
WmHjumiLBfGB1N1vSx2UpdTRvlENkCbGXt3Cli+4/HXS3ijDvtQn+/7vRIrKcFgG
lfaw00rLQXijvH7CtqQS6NrII3uBixGYCUJTKlHA9t6kR/gs9tiGI4ehw55m3DLp
crU3MHvxV0QKTNkpRIOpz66sIvGRXOf7d4JJzWi/X3InIkxf1FEGUZELCCOW9rJx
OGCrgXVIyjTIDgT75Jyozk+OcKV1dDqPtq/QVzb1+jI7DN2reZr/wu6rYC0oeQeo
3WayguNIA07UkQF2A4U5ibYKjrTnuO5a6Ls6FSNzyKZ+lIhc/BymPqWbKogYO5N9
ReunaJ5LpgNEZ6h/h+u+g+iHWM+7E9Bom3F2SWj0inFcYHg6ZmBA4mK/Ed3Jcuy1
dDr4W3FnImUmjGBsxHVxEhcryeIhnV7vIEZhpsFpfYHWD31x9RUVpKF5Qrr3SwqZ
FyBe1q4XwjvSN6q5RwwEEPnEpn6acPfwxge/Wh9yCcGKrB69+3B6ArC/Wvg+EDVN
CAtbLUNFZqRfnCiQkSPCZCf7h/YaKHoqfiEDChia4jgouZCT2/s+MwBxpnWEWJ54
1JYXEEW2kojtac82uWFiERrFlGlwwUNpruWAKp6UxdiQj3aqkhYL7F1PMIP9uNZw
OD+ymnVQTPDkUAjAVun1du10aCs7rutuNoXTDHxcmrpTOHnd+y5mm+znxHcuIcr4
U0Cz5wZID6L51sTSqbOePucE61TZxIEM+XOuDNJnnEMop5xuG/SM4UBGPPeILxb5
CR68BDmYhPiPogZdOJuQHBzR1z1WZdiXZ38QqlxmXRkbnWbXivXb/GxyoaRVg/tQ
BC0XLIureVxrijPy2Z+JbpcHV4WKn0oQqoXlW/80w3sKeaJ0QsPA6DcPl52RSEF2
g6xIE7KMJRoY+pRmRMTI1RSIxwMPU/tOXTkdXrQ5WW3ikxSZOp+i/gdfHILxE+Ws
imJTwUrxTEMS1obzqR7WB5geLVPdPSZo/oc+0MaFwa3ue23ZsAp956TlXEG69HuF
HB8dSpjHoHsZ3tps/fKggAUiKCJ9uWmWkfAz8mqNbEApiPgeF3EfGdAF4hV4rTzX
fhM3j7IUsed8u0P58Z/BWerSHGwcCwME9OeFM7ZKsELPicNufErUY2M+wVwQ2/KT
Mpaz4+ftee+dLzQp5A02wrur/rVWQsMQVik3kpkSA2mxZDo1421ftOdPtFDoYwgc
iZ7UcFnyYFfGN9qCYOtW4zrYqJv+7P/0qfD8F+Mj7pwWIQXJkn9SXqkrRWUwjCdm
RL7nSiXcQbta71ZK+toybZyjaGi1iAXFz14jL8iV7og7uQ6hh1w2Dlausr7CV7HB
ZUjoSZf9nWj03hWayX2weQvzSE/xdzj87V/QSafliZGhioSZvFY98IeiC0+Zstu9
7a9M8D0OJH/WhCeDvfibi9nlbF/oy+9RxDqhBoXK21+AuHGNL0IMB2WfAJ15oP36
IiA5YKmVEN5y6Gn1f67smuCFq5idXnUSFYwQhzEvmno0VgdeUIMtyzvP4CFCaYAc
nLs9XoxbipMPDMovJFQ8h9pQHtTcLfZNKjXIO44YzKHx7U2s8JRN/6vfIc0TPbBd
cIlNSwaGbX4BrEDPQ0M7Y5tanIKnqberoAMMqXJVR28vlEWQNyz6TsdR0EoRUqhY
ikg4t8dWqsUvneTVSNoxSzVGySpNfoo0/qKRdFtQB8el0YuSBjqa62m5q3bAW6Iy
3SsFW+ckZmk7dutMtHrZ1imoC7R53WEafhWkHvgsQu3xpIheruKU1aveMM4CY+72
zuksS3XmH5AAlk+1TFJpOR7Da3sePBOJgRmXClIWHd09bZgs66cfR2Oemb2iqFjj
GtzUumjCW9OD4Z9o5jVViRO7yhCVFLW0cRqamkxxx4bXNWpKczY+iCcYd9GytkBt
Lfvc27ZElXi4yjjP5uSH3zhTOifVf+TCnlvoYqYKUm+75oBWz0wwQ8B3YCnF0e2+
6Ssjtk3mLHxI2csUlglBOB9jEFFEIR+sZ1hbwXwEm0ZcGbgS971UmfukSCNiiqut
1a0MgHE47/nEVUyNnir1+dF9tT/3PUdujw1BaQLJVsOemQOQfUkpRpxdSwLcqy3q
Hsuv7jW4pO34kYdIYC0buBfIlYH3BBlX4JheLMiEY+WfjmhFg0OW2K2o2myEmUGr
9J4M+ygSWM0vId2amXx+QbmtZiP8gxLyR28gJ+qc9/wOkguoXuGku8MQRaFY19Tf
WBD+zd9yRlVE3hKZlblY7ctWr/VCULK1uwofGAA/1TzhpH8kb5rdOCZScWXbahRw
7aa423PQih8thTMcM6v483dm2U6qoA+0W4H3vx/NgLj84aFYvgPYv51oDLGahQWf
d8raZyjRUj5RbAvoXYnajzJKnduUDWItu45oooeqSbRzUAfg1Tp0zHSYrRnufmBL
YhZ9IICy8KN3KlkpLPsFRe/wwVf6djgJlMybIifraJ4J019HiNa6kWBfNXDCn8Cx
5Eod9u+MO3/LVraEVWzbQE1d2j8tbPL1pTfTUZXBlKxhpiiL6vi+aGzJKk3w+H8l
MGbujGzuHiCrq2pdxp4jk4OKHHd+3cqul9c89nS+u+ydhfRXjgrdFkIJZosQq3Jh
o91mc8pwg6JtU8xK3y4OQw0tbK4U4rpTBGEWGLH0EcIQ9uaTAAmYTM+VcyO6GTzN
T7K1Vs8bqDKOuTiBMeBvIqsPiDAJRWqPJBd0KhHBncuFGxFviWdW8TEwxELTDOnW
8kCoTzOqHeS7Gs8EkY6XTwq0w5LnZszgS7ggdTZ4KmqxEyh2ZySXNalLMQwg6bnI
ZfXbLn92x7izpKnHbxoQOLUuXnsqt9OUNDhxmoKIMKB1XffRpasYjnatKkJSBgcI
8yVU1biXbj8l6nekMSv3kSWsG9lcypYtBLEzPvlen50H2Dt1RrIC3s4aImF9s8gB
VVMhHOdtto2K0YufjfNZ5I9HGoKgLqRmS+vjwk3Lk39zq6vI0XXy0QB8o0l5/XbW
txCo4E6GximP9yzw4+U595Rs74yPo3gX100o/KZknPHk81PRHgPhWxBv6Wl250CS
5h7+OKSZjOBshfmoWK7kKT7uBbZfkbu3RcANIY01okT0UQWKXGyE+/y+hhqyIOwq
5l4tE2zzabW88QQQpNWWVGilXFdOT6uZe1kL+BzouCwT+Fcaq8GE13D9ISegpOQr
m2uomytRsD6Lin/dTfgcpIEGHeJbwLupL9y+2HGamilxgwcCD/BTK3Bm8HjnKsPr
wCAUfvxkQRoG6AxF077jYXiL0SaarbIoF3Fy80HXmV4yh5IuhFCDsNb9z2LM8nXd
ybEQrYLnjX6tRkoZlVp14r4ZZVZla79sbQoamcFMNp5N7pu3BapbOhJrHvpiwHjm
pMfebcFOvWVrjKBwMYlsZ/RrpzR9sQmK5rIQ08dlrFEfUc9GHAwkqubbYOwARfgI
fTdXAOgDw+DFmMTA+MDC/PLsgbaprzBZCw2VF0rvWGPreHmNPzo0N4nZcZnOWTs6
t9+25oOIlngROI+HtMjN+3XpSEvc/SGYObFayff5JFeArFS7AyWzizX+wgu/A2mn
EZwTUI5ryW/oEcXqTsXbr0bWXZfS8tKVF7pML6ERtMfJs6UxydU3+VfhrFPLw2nW
gQImAn/BnEGa9XkJivGAsuVambMw4gs7aBYgaTY/F4+Mi27rdfgWG+yeDGoEox5T
GAkPvmpr+jj1k4Uy0x0BXWY5kskcY1YXOoRpJdJGov398tBhrmqfcYRmx787qPgO
K7F0PwpuiszX2hhMzvE5Vj1gnS0RX2pTwguO0XcYIhF8mFJYM56JbU4DwbrA/Luc
2U4D0x8uwo0Ej8uoBY7ATvdpn1FkeEAiG6AOg95D/VfdE6dz4LZU62qVAJf4jrF6
myhKXZaTadbI9AFoE9Wn+AoREEUAtWyiAEQvXKqA8Lwc1Sebrt1wkjhBKVRVTU3y
NkY/Ldf7AWkK50Z45H5pGK1eRfhpcs7v2kRTYjjs0WYnOALng45AqbrHaSnry4kI
nZSdl5D5NYvbWCXc5EpAKZnozYrBfin1jXgvWFl7TBS8QvMb0y+jRFIrDRbQTvIT
gV/Zk0nz2iJbl79p4eWFjWLCxjS+MnJquK7HYLBseQmzDvm5OJecXMB/Y5K+f3nw
VNzwmFtFC1dozxyC9fZreBPEYZDQnKWgsuHf2ZIuUFQaJFLypvC1WyUteb7skUu6
bVYVjCb+v2qOjV13DAV9W8o03/nlvHVDq51RJVuu+WW6ui4c6rTcXAWuDArhDVOH
+UMPrjgrcMVPHy4N6sZTnYZ2AfwmKP0c25GnlfUHGWInTMJKrYVJ7S1lbCg5+aI8
M8nXrGuVcnlh7FmCQUX+6whJuzem7NstsFJ0XilfqfLI7VWPMjl03uvpGqI6x+pX
4PFdNWJwsbASJ8RnOjAeK7f1WKAEDHQhzSSWeRtUc9/G7N8H09Ags6JK05xmuIAc
Wd8G7ww+hqUQNSrLY9BmRlKnrldlK/ejZpXUbPzdshAorQNap5o/CO/t8lxioKaw
FYdNn87Nnha6asraQdUVU3uzGDIy5mfLECuuK6DF/K6TpOQkFvhupq5qiJdFqWT6
QdDV+XKFumWoNHCc3IQZHiJe+wOUv7/PMWWWhH+zrWtSF9ZfUhjk1jizDyTuP9KA
U42segyzivQ9wyHBPyFOgxYilMFUslFeacv0DAoKPnNEcIUPHHuFF7xohx94Za5+
MSYztTcFVID6faLVzkjJDr7nW6BdwEhvAxLCAlAXIDMWUcuV2ndggccIMHOBIeic
3W4BAQVSf74D9A2yvsDxywjp9xGyLXeUdGUiZYINewgtbVUKDnVqnpcJRbYE0+CQ
cwhpgEN5LZ/9Z15rk1AZpWBYBvtSpIXrrZiSdco/VlYFU2bORIxvkQ6ACaRr9CVu
1VE1QvEqJOpFtxCqgJo6lzv5oeydFEatNb2al3V6I3D99PCEwS4dZdia67lNwqzz
U1MO424UIGqxJbDcKjHLdbJUaaHUTlXJapthAlZtbQP2ziYpnrY1qLqROeVOb30K
4ngQsS9Yopcogw5jCGNsvruaqcL4UWzFtx67rNlabB8Fop5g2EUYLNQ5cWH7l/tW
GhEKi+eoLtoSOyFxEdnFSa/8PzRI1uWYJYWR97vT5wWI5qlYCepjzk2yljI8mB89
xD5FdnCAT9KpxSa60anmCwDaab7C/V3E2klCeV0S9xBEH8e5cwCK04aPCKa8j9ks
CO+8uiaVCHHPhsOd9fazy0gLE4fEZq3LmZRV1POYnuEfHGqNy3RNclq5Qk/RBcUo
+vraIEWeKz1V9WyvRlbzV+rlwr6qvKhXf+qBSIT8/Hm/yuSFN+MAse4hv6e9B/YX
+xUJwowEoaNAgvXuIAE39T2n1Ls3nNOq8PMkRcqNQFpSdiGAu+7xjGGEIMAnU9Ep
viJzx7iQVJgi7Lhw11PEdNr6dUQPbx5QZXsVXx0Dvkm8inKPGiZbL8+qXTA7hKqY
TjKCDkhWWda0I/d5QXp/ijc8C+BpENxCvTpSfbEe7YVA4N8EDPgyU6ZrE/qI+U2Q
0DJN93Ud2o3yxviyjpWmcLmoZVa3iDC2EI8BlUy0/Z25XIijG7UZ2rz65MldyPEG
5Ps35nRq8c+ARv38FD1Y4xWKf+lxeT8HyRGSGyX1+Qko0aR25EnWuUXozjLWDFq5
LmKy8M0wCdg9jWVgCUSL7Y4p1Iyim71v8kIoHRcvJSKEc1md3/KMRQeR8Yc6DBIB
GQbdDFr99Ru9iKnBrfWGPJPgM4cyy55GAEStMkMba9QCPPC8u6mcHf7uClSYrlqD
BCOxTKDNsn0oa6G0X3K6wnWoDWdWhJMx6U91nkJWwKQyATb9M/vqNHdczZRMRP+c
Hhn3JFZZ4JQi0pN1Zma1s9s5gpjFfjwwg3uCtcNnoP49oc9dywcL86YYWxKs6Qmf
6HPNULC+c5dErg0TYT6OysDYiiK2w5Sq7HUX4uFw/GdQgBUNKv2ul7pSlppdb+69
S3EKbljgdqp8br/Hp6IB9IMAi/AkT+beAa2RIhHL+hLzUQ+CglKVInUAwKYbuAOH
bjt7LDQNrZ0LdCYhsuc9cfxFfpGxrHJr+AQo8S1aCQmq7/3cepZkIvTzUuCEoPBU
ZNKSuvkkiw4DJm7AStArRWGfPPvFDn2HV70Qia5Xk9s8FkvtpE2TjbM6Y2a6HT8M
lLZ6HVGy63zZlO6BZDqjtLIGXJlasRKabMRIidp0qACB8PLQsh5LRoq/VP2aeRPJ
ORDBLPvPemHQFI90ckKOuV2rIvSGcWW9c+3b88W8nXhHwzoWe/59RSQ25aIXWflO
4G/GZjpNtC9y9t0YpsXQXjZszvF/I04Kd4zsfLLaSaSruye0U55bSHpMSvPTJnSQ
fP5uGxgK/0U1YlXAx/AR9NLfTbOdOJok1yFoQzYS/n2P6PKZziKLaT1G9uLywpeB
TV259gwQFqcXFRI/c2t6yUhnDClU8DJVm0br+ej8v/r4/d5687hgNvNAep3ZTYYs
oWoMIQro5McUMlyTEyorIeorOKf10yeN0Qn0xpjzh9RgxnDZZPK6i+gvsvR9Fu1h
xtju8TNP1+o9fRcZJiMlcdv13RcCgHt9EuYy3TuIkzlWUC5x4A9pk1UsYLg6N1D4
Q3Y/MiDosap0QcARrBEIS8SG3J5VkOwtYaW7AbO7j1FsppHaLACTkD4ePw7s7DtL
11j29U5hQSQm7cGyw/g/hxBIyiHrVqsm0L0aMymwkTihpAiDVLBOerfSK0oFrPjU
lPwC+dsCRPY1CXt8P3eBQiRof4hd64JQeOufRTkrkNa2OFZX61n2RtpZtMfTdmjd
Aww/fqb5yiA/So+7Ufwa31ciGuyGHbZK8dS3h+YbMMLDW/Kuy7FQRfy9ZnBCmVN4
bxJS0qHFVu9qOP9dNh7MgHz480mrF+RFLisA4IIbgGMtrDLQUu6Pk7oxUCgB3ncC
XwzIK9SBUdaBgAEJxZXJrQkmEivYi66qPnuzD9R3WzWgggs3JSRqlvvyJETE7GKw
BW4fhTaZ0KbxO9HQF8OGKtHGglMXd9/P2KHpbD+zPCMYibFkVdtDAMtxuSYnOkAM
BtgG9M0fhejiEEmUd3KeM0dxix95FA6HgSuDSEufeRLh/5QM50qpjTfI5amOvPPB
K+GglPfoq6BApejExoy/7kVON1e8EyG3kF/12mETpCSY1Ou/hYBuaD2D71zmsAsp
b0ezdrzSgsHuwYm3I3Q++4SQ5zT9LeyVB0ueTHvxXzW6zcSogcKGzBwTM6O70vgu
qeHx/Udq3SGrITOQyNjYhWdWfTqzROTvdWEQH/uI2V2v7sQzWa/qzzkazw3s/G9d
xB8+IdLgocZN6sebGxYA93X8CwZ2avkXA/1P29Vr1p57F53OaJSnJczdnyi9hxUv
SStfaI04W012fLCXTwWi/36XCQOkRdyL7vIwcWU/ZsmzHLjxxnmN5+pR+66UFSEv
SZIgWKGLtgbfJ7ixaOFsql6/B2EFB6X3dvqMOKwxpbV+C9nHAyg/9HGxMlkmeCrx
LcZuJjHD/D8TNl6ftML9bXeahpl5nx1kltVr1nsxyvT+pFmIoRpCFeFCRM68VEHK
O24J/642cAEVS/0tikmeL4WtOq1gT8jk0UBbejbgeUXJlp1nAd+AybtCowYosdpI
H8o1Xtrf62FOzPssv8CykOqoZKOyXNt5k6WgKFSi8bGQbjFtHqRqvptXW9XfLB3f
1ScwGKjaR+w6vEtpj4244QvRr1PpevOd5o1xfjGfjkjl5j/J/bZbqrxXI5y6q6tf
W4aOWhaQmMYRMv+nMXDAbuFbNm9pL6nnabc0f5OgHHSlyJt/Y2gonaUqHlkUHnUw
6Zs2LVzuTgNWBy8JSDPwvDdeRmlZmtU3FTnDA1qkzNBhh1r9NS6T03fyAJUwq1OY
ZPrI247sZTCxe9u//YNN7+pCvQ78QoGKVmxWkYK+b1mm0Aww6oLv/wtJTeuKmSA8
TPntT/Hy4Mq02HnVHppx9lVD6lXGhsONx10ctW2xjcBEY1LEr5m0crCu0b8hzhVS
aH5yE47oe+V9Wrwu/2QkdqkDSoEGLORTvUulmDmBLp7Vos+lPNG9CGxFbMaRgHEw
dg3/gZJCwu7ZP3UAIkotwF5hsLhfYnJKkbNcUWn9/y34nlB3V3bPTXU5+iSsqCe7
eQOBddbVgckZiEZ9Dnzl5LMYcXqAELdubTJR8ZIbBWkPen3Hxwxg+eCKi5kQqVnW
js78rtZG0qlYkQ5zxu/9v0yFR922xvJNkDgGU+GR6Mn2shHY4WZYwAujaqKAOorW
umApQn2nqdCCK7UCiRdwt2IprwZ/4EcvFqg/x9BSR32CZUNFShe9bQH56seSQB2o
SWCkydqaCtAUmvd3F33PTgMrN+jYg6qZr31upSK+RKb9JK5JjFwbND5fwpayImt+
fXfr86+1x2yscGsDLbDbYvGqBMoOUnvqSfcnJi83WWp75csQWIsiSrYXiGRQ1xY9
/9dhlxY10mpPh6MP6kRr4HKJWcfDFCeaysiFlpqVSw5/Ut/qYiRZp6lx++feKU26
b4EvEbRN+rUqhNLn8N8yEyycDisS2VzbSqBjJ7TMte82abJE20XRNX8gv6O0dmhW
9xP3wuY9IBoT/1l1VT4J+C2pVR+HcHovS6N1BTXs34jPT+5W+Xo8Lf4mDcKq61hE
Ax90xvxuXbWKyZYE5pWsIzeh4czmJsYaJHTATLbf/ZEh1s0OpTGKbhyQYXeHQS3/
GpekDnaNwenpyN9y2CjsiN9pbVCoG7B9JnbdkgWVhW0v5UU0bxDou2A2wEzEuQpO
nhdqfvAmxCVVQqvtf8O5pN9RqCWkNqnBBGM++1NJ6A2pTYLOWVB3MtjpD6eHdYDT
XcYqs1PIbFkBuYG0MeAnzdoYSEV+qg+qMwHvPpBcl7wNBz1/SIeHY01hZF9AKg3y
kgM4vFv2isIUxCFRAW+DVtXSVILq65uDWc606TLc/LdJNVzTBK6eMwW+jdClZ1Ww
4owkcDxcWuaP32prLY87dzFetMgAjXROBWchH3Ta3oC3NAx7g0lnhDJkoxjoKgAX
SI9MV5A9pnx7cUSozuF3ojf01s1b8713qUxqGxKIL1TviaRqCFMpMwLNYM3sxZ30
j/X5JBSanRahMaXspYvG0hZOe+1uOgR8h6JfjNAYPKal55/9jvqncoYUQzBRp7/b
6MKRd2Fcr5Z0HxP2QQkC5XcNJk5To3DM5oiPcVLDkYm9JjvHoIolJMPpWwrMUUiE
mDE9uO4NeQzBOYTmDpbO+SgU2J5wSUCioMWsy1cxU6LekVNneNeq8qw+WVC1EcVV
t5rgIj2KJIgf/P0gj4UURWcSpAjdxEaEAkFZtnAnm5c0AA/WshQ+Dyjak9jyBuMo
PiHIfBkSf5mfW7a4uHckPNYR5qub0V/5ZMlxOHxPxqsynnRGTq/thiLDIjimzfiL
yrXa3fM4cmcmGYBDBayp7rWc6/Qu9z9H/2jdLjxFwb++iGcZu3ydnWSWj/UNm7kh
VezoZYOVKkQC+P3UL+Paq69gF94BaAZ126CX5/7DkJnCDmGPSHSvtzLcX5egStU9
E06gNeP/YybC89Fo3sB5i861EO1VXj5fj4KXrMGyjZvEGGvDx3JT2PMA/nvXocWK
5JCYDbjm/qJRakDvONLLLTMiPmuMVfMSOCfoVTBs+g/WwJ3xvot4ZMW4qAW7R6Za
sZNEQpPZro+IqeACzGXttIxYRYXZnalR/gLWibw2uHU5HSNjhD5JBag5n+HQ0kGu
rEvVAHsT3cj1g30zWJ6CNVIH0lxkcU7LJgWhEfnQceJaQJL0eZ/dxXUwNAMOkjm6
yVjd/3x4GAIgr423VZe9QUqPr52rhKuqepub1u2kbRHVUcR7veqpDDOVWhy1elgO
sLc5+RF6KzaUWLtbpIBpFpj78j70I2MC23B/66R+FnfUoZJjMs+22suxrlKWTyZW
EJiO61I5Wlj/ecEMTm2OUBLYRtvvWwyfFVpRZ6Jy+9sW6BTH4ouxocvD1XMjj1iZ
0TndSfH/TZtq6ikhL6zKGltYLBUldf5BUIDXbo2u11823zrjL82Zbq38bK0Dg9jP
a1qABWdY/jf+JWhshojnHjYNsgFKx5i63ijmlBdBP22UFSzw6lmINNrQhnCn9Aij
8Rt40Rd54jqotMWmPjk7LC+xO/yBZqaPkrkFGgjPYAL2p3HEdK65E2ceUNSjK7oj
8pjErrJG65uqhyaio/OzKLIizEB6uc762HhKvNePDXcq8IHeVLjCzzuKwfZ6trfl
zdMNnN88/FeuYQaX8oqBAFzxCoWiVafVzGoXmCbwk6/fkLTsQmytqYmF6oMAYiop
qi8P9kou18hWqFLkjwgF/H5J8+qtKxZ+2E+3LoJ9amMIdgtJNYJfizwe8ompL9lR
vHYSg3aGwavgZRmClbx3KZ7xXCE8EF02QEq5RP805HWHutFoLlWWxVcrHHKM99Wn
O4zv9Hlln6hpvuMUfaNxUnViI+eqrv6nPKGSlU95wDL0UMZh1XZLYhxk4FotEwiR
fHJBv3ha9aQS9vgf0NOnvBy4Ju/1FnrDtcMDeNDSUPFQsUiF2WUgsTqGyNrQ9wYt
k8nbBpGRauC9w15oEP5Ww30nYo+OhGy8NAZX+rlTkqjhUJr8CObrL0uwpb2lMKLl
UTVnuSAPpEzgQMNyoARbf/f0t9cgStciWAt6HLt2Xg/doumOxbmbBE+drUqUCGQ1
7pk2/d2l+tNor/pPeBrsZ4GNUHkn6eOTX/vTdBH088jYlUMOaMXp6VMgNF4W8qd5
j2Am88e1Q/Q4mW3AL6V1S5P2oXQwLU6JUjFh0IHuVksM18r6oEmKIjhqqYUYLYno
AaBgeogl2NFWQAvpwLAZUz/6/C8UCDDMKOPlGvO8xXxSA4XZVKT1Ak8BzyaviuQx
WVz4JpyIejq8TAx3Z605JlKFLEavrc+8sJFHSYVPczJUh0Rt5Wq91tc4jgJ5KNbW
3i+DWURgBH07/2EkBIhIjHDQvfYoq0KsYr4xqQQzi8c2wotT0Q/+wsBrqaMhUqV3
7Ql5mRZN2pseyMIqpoEQcCC0/+CMyAugDvFSCTa++rwahpqy/Ck5NMIxFgsQwt16
A/gPLjvFkF/VLGO5OLweufe7yoTA3AubX2oItslhZdXj2M6O+4/d7nObKE8M+b2V
DrnITZ333LUa4iKYYMq3TYwwuetfvS9eX/V9rrq8Ax56d1Qj6aZKIZKAxqJjjwUl
Rkg0/II6LRohxfsyxLxuPNb9Z/DPWRI6ikgHiaiVRJiTRrmEcRB608KeRwpN9bE5
65E9rU25WvH81Z/ciO+wy3AhD8vRGsf45hKezBv6Hqc1qsRaC/hsfYw1EOfXvIua
1FcBH6kksUNPp9YzxnxkF3vJjpcmnrW5R1dAFjPh4naat/gQFMIqu9FZkCCOEqeH
zXh7PAh+gxQy6Ojq0ZueQe/02c9OpSVTzy+xWQ0cO2j/Xu2brPFqkQM+np5R47n4
ijFMJa7fZkUlAPfgJIt6dgW184ZbHg1/qYEE0t0RiIfJKfsUuUCOMsO6Kd5eDbRU
TShxwbzIxXapQCGZgHFnzRsVWgDS7hA0ps5SUEvXmIc2aoRiqcnd6b5cfTCJr4P9
G7uqkqHQRJpA5d65gDqAxOY38OWpxzFIpR1ZJPSX/PYwXyC5bz5utnCYGqFM1Ghs
BVVgpnP8cBciw9m+LHJHlGdpJbDYgOIv6fNPGyzIpst468m2IsO7d7oV17cMIgJm
8WqTnzipWYzEhgeBmJPD7RLi3q0l+nB5+/bQWr9sSHoo0L5JGkTbQS2s/F5f0ZQA
emhN2l5YbAoT8qgF2XZBgruW76kEHtCBDPQWliMrHPDLp4KDCYOONAkXc4CphDiC
wGOb0KcSxvLJDclgzY7zgBD8ptGbblZsrwqrffZ0TcF/l0d48HBn/nH8KJVAIsJw
si6vFLYzj5DQ3le/oS8g9FxRvVdRsvm6jCxJON9u2xRSZCSRZAbFMgQ9KAZdhlFI
gDwFBNBq6Gk9XOl0CkctShbOVhzlsEZudrMXaAtBPqv9NWI9LSaK28HAzfYinWjW
vj53Mi/7PTeh8mneBFRWNrSbp5sbOL80sY+mAHHwIX6rN43P1HeVTTXBjw7Xf51A
yb5EIJDg0JR4gLkfSTtf6NmW2wfhIjH2bq0xu6UXx/ZCMkfG3goVJFFD1X2glJE8
lsBFhUL4Zel1VuMSDSYq1rfIDtDOsIOsyBSmENhFnpesCWtsDWIwQMotjC5HIyJq
+3d/aYufXDdhNIdWD+f7XzThkidFmtvtYlCCHv9FTdbM3lqxnF3IrGN0SFh3eTVc
YIniqv2avJqBN0OHSIg7oT06OdUgxU/6rqjpgLjk+M86xGjAruWujJ9S97xveat+
VbSlvispIwEqXeaPi5xmG1kt0zCwNtcCkTmjAYWmw+0hzI7L6lFFYSYmQGiowrnz
0Lm2gWl7fLuRepGwqi2ycbxTWbtZSngYzRlGnzpg4HYq++pkMVIKfSFLjJ9uCaDI
T0oM87wrQSoUJHzP7jsQlE5RotGEfe8Ppne44F+oyelYLC1Mk0NhHKKIuyBv2l4y
4MVp7aZR9NQWyH8+2kaaItcRzrbO1Y8DQk6E9h0UpmfledXNDIrnSyBZOWKfSc7V
81HXxHJaB1h+NdLc1bhLPR5KZhGMTLJTCTbJfakFGKXfvV55my09wlVD/BCtvphm
gRUxZr4VgbHHzRhuR0BMa8Bglnv86xCADo4yarevSG9S48uG/h3M2hezpn0gBikW
gz6uXx2bX2GEIMRgTQpT5kkGfwtOXLGcm7rtsf1P/Dhw/6v3EOTqlvussd40PWdT
YMK9VU8NbKKIG0PH7oyoU1gMEzAyiNoXOhMsQZYYk3TX7/24QSUIrEb8eOfwieyy
8OMxabPkeZwVrGDrNJamc8dBt2XkKqRUbHHolea18mbcysYuy9m5fPfi5sdMwJmy
x+xkV3YkOO+/k7g4UFTVDN9TqTss24Im0cmvgqC0gi1oqErLAgRVWDRQma7LJ088
EA+SnltnPw5o6v4fspwxQKG4VXD/twKt4572q3IwGeYTV7GKbVsAKdUzacKyAiZ4
4viTGS/nYNkYTkschdlhbiXdT1jpgqwAKosfuK5db5YD6gcD3jI60+yBqc6IdU5H
fnax9ocFZr7wV0DP/IIuNPdWMWcx42d1xE0sKMO1m0WuXPmcHh5MB+BzYyfBOGM4
n/Soc87xrQfW6f5Ye4WJyK10KQtki3FDhG+h2FHUhwUz4iZTg89fkoPChwEqNNn9
be71DNB9y1ReeehlwMcu9voIyBlCYG5NqCbnvWWnrR3dvitiNF/C4h8Uw+rdh90s
Etlw53fZILHCMPD56BEKEIagPs7lchfBFzwCt6rY7Q34vJO/h4/neVlfZi4d4jF/
12Fjpk6yIx+xINn3vkZIiCgy0oJHXhz/W10hTxSor33yCXnoi1lR+E82uG84DH/h
gmj3knH0zunMfXB0tqpdaNizCEwCgHH3sx/vte9obIEi9+I0I68Hd/+26AeXCjc1
+KSFFAmE5QipVlwjgpD2KXiEPG6GgcMZBPohrnigGkp3sWZsEvWd4N5e6QtQulMe
st4htRfcvi4rIRm+1NogkZeSf1agrxcm0mcM+65obEq1CGztL2cC3ILWHflcL/J4
ebC4F1hozneJoSHKpg3h0I46IFnz+8SHnhcGV+Z6jQBIVxDFTp4xK3/mn3n9bVNM
onoHaYxz61Xk69UmnH9PZMlze/MsgMmsoYVXdS+breBQcUkdrhz+Uy8YWtyYehYi
qcW50Y7OcmtK/LIvAEVknBEqouieRrS4mjnaiGymdov/0Uw4e+Pi6Aqh44zXbQek
ocIciekY8kPfG0l+1ndj1ivyPOAjwPKjsIoSN/aMabuA9XG3Hna4bjKBwUrhb0YI
lTajhgFTl8+Xo0SJxyogj+LX4UgTLvKRmxY3L7i6aQCMUVK9T7ZfAgO+oYmBEcWv
fdP/LdHdMPCfULfjILHPJg3DoR5qJKj17PRL8WFD7sIbnLU158pSYUQnSneYuYY/
92P3KCKXXgRAPQYcMpT8aVS3ndCEgFLyLL28hk8IDVbE+rxTBqaHKqKx4n0QFN2I
3Fx6NzvrQ4pXFXiKpwkdt4HqVT+r0w09GKfvBcYuMbw0w5Tbbf/DKYIaf+/31MtK
zcwDNhTA48hpJMksffzfE+2mzqef98xrhyk3xN/couj5PcK7LVtRyuHPvZPnBIyH
a+vztInhdvxsQqi3ilE0MtoxY8XutTkgReU1JL1opCSdgTXqxEBNiFJFgqPApm3m
T6Tvo3u5w40Mytju03ml+9GSXR7uGk18ySMPdE3PdrFSwo7wkJ8fAlhYRkQwy7Fc
hZiiRJjIDaUdKiChvf1wdrd9U8PgZ/6c//4XzzHdTRZn/JOOXwcw4OG86/GkcwPu
5LM4sLOkSEy/vUQa0/lyumVD7bHNNfl23ni4IIYkqiyOObqRUrC4rXYNbqWT9xLE
bnFsy2c+BVr6RxbPFYwusWh9y5K6jvb/Do2UjU6KrJh1BtMoFzpXpWQtL0qUQA/c
LaoJDgAIZA5IRWIIuW9NHu4WKbJMkfZOhZd8YYOYC4ZcAM0G0yKM4VorzXmv24xv
8LQYf5a5PSnuZDmsRztuSqmQ0sxP9lMBYu0rBFkORjrtTx9t412f9JqKd41QKiso
0BSnwrBgIEQWtO95+hYt6uu/3JkxXL1nSHoE12tBQXl1GAU/QpPH9bUFmPGFbFcS
/Jl5ioDgvsjMgo/RpsCjz/b+ZWEXVb96N0O/k5OM9CliA15A/vfC1VP9Ry4nq5P0
O8NH/ngKeU33UaHC1bG1BTUHoJrn1Q+SLzufiDSu850HC8QRA+WyJAYrmAAS+kM6
6ucD8MNpgBYoyfrGss0IEXnkrlSMhioqx5zDHDABjlCiKoTJyMDNZiHhG02Jr5Ed
gO7G7YwDsVBxpoQe8EruGK8wnWLAyeqV84bbcTEs5vR0JgfMeHL3USTqFhcW+k5v
O3pJrWJpPv3IFntL5KCJ1pGrK4c5dgnarFRyfZ7aeckAN4ZFzX0f8V+pyH7Qan0A
8cjAMI+E6OMw/zAp+ABUjwvlQRsNHGY6PPjS//KUvDCToPF3zhv81Z7QHWpjlRBk
iOoZHkQaO+S3mtRo4y5CfEq6fa84hsxRjcxX52MBlnUZ2svFRwp25NApj8evBVvM
N+HbofDhHcFJuVzqKfiWWp4IzWtKAFc0a49yK4LVmdF/6P4kn6THnAtdRH/XDflQ
fhjS2sNzrbtGowNNC3pWsm4Eca7KByoc/WQkDXeFlqQYEBiMsQy1YF8e8J1or3Ir
AKFCYrP3a5hw6dRF64hPhRSxGX/whSefS5u2qdmWFC9SJCbkH5MnvNuVnOxRJOWW
ROOn9m09BX5g5aMXuWb2c3UqoJ2QZ6zhDfpSh+KP5tizq5cG9CQnJLQNvv3WbBsJ
7S0VDu7lBbRZ3erzJsg1Fq0MjMjugnW6xoXDcoUZCk6GDWYNcS7vnlv9e9ZITeVi
+FGrDBxyEl3ohzX7pfAouynm17FzWKTDJPbMQO9nT7i5y+/Gkhc0nQeYu/zpsX0B
4DvUD2mjZWMKWFgivNT0i3DLuaupfzod/9e1YduvdrNRS3fT/iAXCF+R+mWpSoIn
k2/QH35T2DjlV43SuBk56F4+1vONAe0d1t/v/MF8DvDBr6EcCv42MynMGnFVYdYS
JBM5byE6WOag9wsSdbjtIsrxna/k2042Q7yrtDwIRXmi6Px3Evis0JW/XIu1c7Jz
lieDbh4u9Bnb6AeSejyQ0v27u4vKU36dTurBLceN5wR/TDG9QGgu+JbmkowuPt3X
1nbLyi3VMhMkPfo9Ldhk9t7XIyYq7fo5NoeEznsBlosXnDbVcD3vIJYxfdNqojNs
kBGbTj7Mzn0a9FlXlZ56b1uPkLn/xE949foG3cWSdBnHeipjYSG357Ck5AVlevIz
E8I7c+TYzER5H1G0SsuF75ss3cNVGvod9e2ixY3IXR5ufPijN4htYga7c0ohKc93
lpgIjw28JWqqT3G21AvNVsfmHipA43rONDIn4GK6AnEAi9WwO6iIC4Gq97S0iquI
ezTfQ+JSedf7BZ7PCjSSmTKnq9PwcylMdud15wZsobGYgG56T89AHN5ax02r+g6m
Db3oFyO4vsnOrSmncoBuVXTBKsFlVxlA4CughS92FANax3DS0SeuRkZUGuK2P6LC
RXTz7B3rVgUjIvB3dCMv1KLw09dsh/odYj7x8a8R4IptA5bTe0lEvVsAE7gCP/x2
oZC2kXPvy1TItY9h22ieGELWw6qZZKr+dVlIaJFAYyio3n+UJbzURuNoD7r3Btny
4jfXXFRwpsXF9maD+8MZvL2yhtog0QXmttJZyAc079IS+EIK/6uIYM/GgUxaePza
CbGeDbGa2Bxqyb1xoSrJmPqvvuazumfZYOtk7Y/Q3UC80uNWO1irSAooY3v2n/4i
DvP6MUmoHRajwFeJU43xsmDIG8KHN2RXJSPMHLGzNpcVy9MLclcwuchrc6bXXghU
7kis41QonpXcbtwrNYrcoGg7AwBieUGQLR8Gb+q7g5i5c0PZ5YzfUFmft2wE79jb
9dbw/qIRnNH+oY15JaztFnhkFsKcVc+b5QTReVD7M9Yxa5UrXDs+NyhPg39gOT+E
qbsEwyqtUjn9oSFewm9qWRpTbRDFD3QCAm3TTHnP6zfsKauOctzzHGT5vR5cWsph
svzkNOcjBXf2Cb6EZU4hw/TY8/hAvA5yBm643SQJ6EK1VDWNjA2c1pkLmAHpScyt
785MLqdxLHYORaZ2j6vv+kcnVY+91PSHP2bVJ8SNJl2IGURhzj8pOKxHRepE8OeA
pDfeHIGT6uMvko+ai7JVTV9Tbr4a3Scw93uZT/xZ7ORT+d3Fqnal7bXF4vCbVwS1
bMSC7I2VbsmWodJl41I9FeEJ5jBoqBZjF1mmJd3nl+mdq4IF61mPY+feduPd1s6k
FjN5B16+qi9v/09fkoAUKzqWNOov/iR4S9ioO4JPVnhqSC3QZerC1B6fOrGB9LpN
A+PnMS4O+qjfBIbGEvRmLQ8Zy/VT1Jb6bbvdGE+TH2yNuTiq1pQKZ7eLNew+BS+R
jVL+/rzq/mD4RZgM3cJNJQoionxaxpy6osn/VP63DQwQc1WanHzVaNk13RiEM0uX
AB+i2s6+2fG+R92LiyPODiKRp/o8135UtRxfZwmpHQf9DXIbuVX/c+yhK6lIfkez
47tDsBeQwntQW4he6WIXQWPBDBEnEz7LoLu+bteUTYM+7PQHWCLdFL4rrrnmVzuP
eM1qA0dsVj0qpLql5v9clZ0rsCPkpBuv9OQp7SwREFXYlCcHObzJg994i4UdNdkU
2Wn5rD0QNZCun/KycVBvV1WsurJevE4ccZiPo4g7XtrWRoYY27z0NV0FEdeESR2M
k9QFU3+zdKY9sLyRgABjeMRiL1beFbZi3UyabCB6JkSufin3FYuwuHqbfspFBuRU
+3zezDpXc28ZEZ6ZkSlnliRjpHgBjMGxm/lxy6HFKccdwvTP6WQqzQkLkI8lrxkS
v15I5rbVrLJ/RJUQEqgMjwxs23SBr+4iV/5X6ekr4bjynIfB9Z7yHy49GN6j2ss4
Qtk1onlz4DZf6GxnWXbPsRdPDMzgkgj1i4GtRfX49xwar0fBizYAg0/T1d3AABea
g76wN9w43XRqGKhGecNcvYzF+f8eA4ingTX0ehXyDGf3ZolRwLsmE6WLI5RXQwjH
KhzQa6yBA8qrbxdn9Ldwmb8yTmqBEKJyGHiX81nY+ibrnt4TTFpzPXwQMrJIGsk8
SUKIccmDlYEdl2rRYouf4CRjklRFm6DXri2wXRdUfqSvoy414lDCITZBiPpq0C7i
XdMAZOfWJFQWUU+QPyttscl1GwyOvLKaRrdBY7J1cwRoAq9EbYN9qFo7yR4U0CtF
vQIV8Vw42SNe1q1xQOu3pKhvXnzorFw4ycQFSwX6oaX/c2cf5+z3DxEGupzjvMxV
jiRzY98aG71JokLqczycJNlfrJyG0IhKwPw4nmTvS7h22ZAruQI7jyaDeqkRqNhg
O2eucxIyz3TcCO4b0BKoyX1n7IC4bwCWlwxIShgRbqtXiG0JEcZaDLa4xi2oj/M3
bNfH8YmDMmO9WC7F1jd8BLS2GpQySZnhqSG+xKA7Wdxs7wwlZPkaeqfSiw7lWd72
6b6QD9dtG/a4dG5kP884Zh5wOH/VcF1CXb6Uv6wskiEHxMT7+sQ4XG5+vHYjcncE
A09Dr7R3hQeqvjPzgqI0rHMhEQOVzMns7jrsSoE9Vki8mgGkB6wCmALv/E21Q7a8
3Ipoal6x68pq0aInCSm1+H+RXMcYNpIGtwrsDEKYpFqE9sKuGFaRC54km0/tKwIF
jsWf/vaNlSbvK3/z2EvXvLlCJg3C4APblsXd/1IDyPBCpSCx//K4AgAbxW0mMLIC
gALbvDYtm/Mdzw/rlKd+LMUr1eUuZcELfe6aVh8KtvygoM5x+difSkdKrqpWpxQS
LRQJ9R3Djh+k2laqgd8Bkixt2RZvs8h2CtCRCvN4yFQlJ3a5LWVTtMdNuonZhxSf
aVy6JqPM+s2nRK9APVz5w15UcRnEdMQTCB+cpYxRL91ctf1v08IfzadbiQ1VWreE
GqATfGXrATzLwkK+GkRQBBVCuC348rXhLlx1XkXyuGd9dkjsWH7r0Gc+Qu0m12uI
AKC8p493l+5cpEH4zAfzamIc13NAjtLiomjci06ddSanUtlRPmBRM4Dtz6mWL+YU
k1zRE06tZc7htKQPhOrPTO6zMRP3wneRzdd89RX5Vgd2qjZIPCiMvUJ6qO+PCwJD
GKunTe6/ZYGmvpq9Eu3J0c0jOSouzeFG5l+5WH3xTWNLg9qtrqHJ5R+AGLz0brnl
kBwdr9aMlRrJJQgpvj8hLhVL+R6bhiyXCgXURG1Yafi3SnUEULjDRk5s2CwjaCpj
JIDHWNSZu7/RhcYxDwz8ythrkBGbpfj5Vqp+681QcDDx8EJ2HpdHdICbgH3XOVqh
8cKwGsjO+xGRlZXSutYsI2U10p1zuZmukeO1xbIiqaJPxgF+XjMKMz9AVJoITwZU
OqOqJdl7wfwi7xrOdr7yw2osiboq4Vy/OjWQLZzYjllZLy2eBylVgb6cwWb1Kfn3
UGckn+wAKSBHiOMkG4pHjOUT74Zd9+FKPuHE4XI1yW1/NZFfax+uVF11ZpPGNowr
fnrFtjOBA86TPvQh6vkYK1UEHLm3CAyw9f/dgTn4Y39oD4y9eKuZ7KzLjbRkNWsH
lUOF/Nlg58s5QI9rvwBpYx+/VIsLqRKMRrS89/qlK4LBiEdAYZdltzVSVLbYhkI/
i042kGdGTvTMFqSPKsFvCJVDBiDmTZLdX60tzUgnHAD15u4DaoFBmrXQ1713jHK5
v+LyKQLVR8Q61cz5v0O/VG860lnGgusUT5G/JOWacuAHM+aSsAo13GgutT6aK7BP
AJ8BX1Wd7e8eAoZIs8QHYbBUf5IGn6mCDIdQ8DTsiFNXBzoljsQik5Ryi3dk9URj
GxE0aToD6AvPjXp/ATs38KhZKAR8SwABZaOhuBSrdll9wwXpPyqmIM3TPSrNLSIE
Lno25yxv0Tl1GuUnENC8T7UM2F8FTGRhXdhrRJVx1kF1IkA7PDmVRllrSY//Uo9+
temNrlXlZ2OrdhjWu1FeEf1ghVrryV0FK8DmnWIGCHhINxfb8ekoVvvsZxCWG39S
BgjYtmrmi9ZeWCQoqU2Vk24sztJKlyFEADKcJw/t21IyP5d6pqnvQHKoA8eKjFhk
Gs7YYFOlvuGeWHx2YRmETEhXGmN66MbtOQBo/yRZb7M49tCTo1RVlNkSpKu9Kbtq
Sknd7TTKxtVKpp30cNP7axRqVWB7ldeTtASJ4UQedGry3ZHiQY68VZZb6we2wFHi
NAl/f0OEHmtLdzq/f5Mxo5Y0Nb0u3b6h7XH2lrNStfxIHh2OAKt4taZWP5JJHeeQ
8a/gI1fxGA4Av7sni6x0n3ZpO1qY/01v2Stee0vaz1m+t5wnFMqQUTW4lVHvrz5Z
qW3027ZGAgWR5/VC/u6QeqR6nFGonyMzHSuQYFWZQFYxnubcAo8v72ZwLJoWeoxJ
lq4S3DRREt1Zbt/I2mD0yArjFIkyjSjBbLCFDyRM2lkuFjIruVU6AqseXXuw13ss
9TqRZfs6loAiETHNoyxkh8hrBaugQ0DXrj5Sg2KfooN8VjaSjNNXY4MHi+Kz5n4k
yliX7Mb5kWQKQyizxq//RXrG7eIjLYCwQdE+M/q/WSFoimq1tunTdMHQjWxjWQei
Q89KnUaaTLJp6q1ytL+e3RxSAx24B5x2K9nrX0sgFwzTA4UNMP68/Wsb9UbF6UZy
9/+n58oxyNmQnQJCnBdytG3sXF6v0EnMeEyN3AaGbxpG3E3vZaJVB0IH0oGR+wpQ
dYODuPrqq3ayvV84Rmd6KJGWvxovBlwz2DQEeRlAP+EUIhED0+K1FlIlm2xmNo8i
FlZUQ5Gry8raOQRc8wLQsaw6FSwA2jgBYh/CXG3X48be65reQjyOX6xP7U1Dlq0g
S5GQRCev98NYRRuRyF05PImn2YSR4E8MKZhHfjiOXJTKi5LxNkyLxvQTPc6VrcPg
x+GGdTmSMBP9VEqMSim507PLmIbaon9CQ+Pds679BS8z665ZPcLTOq1ZJJrOzi4C
dJXLjiDN6KKA72YFwCe85g0ecSoJya2Uo3qABFMkMSmmJkqy+XotYCuEqUZgWmGk
Rhh++7c4AFG5+BV3IuBP5+3BW4t36q2YHcbngYeEZota8fmLiuqDopBcdTJa+iXn
mA8uvKN4LWfyPvKyq7kEjGLQ5dNm6JLfFzQuKny229D0VfeHqvrJ3D9bGi0vBLMc
u0xcpQzeg8oLTwwe7vBgKK0ksnqcmqBeCcNzR5enilVJeJbf5yREPVta3LxIFPfh
e1XeRTrIMQdDoWsq2H/PxCToE71HXA+Snvvk+Pvhomg82jYQ2FPcjf5x29C2IBhl
Ngv22ukHsUTrkTnXWuSWMuB1A3adjIuQtmLNdGh7wSwx2bvFVlFdKMdVqHLLGJpN
Pv6U2KXPTWvFbRpTEcnT9KOQzGjbBPnReUF+SbiV9qugA5vVws0XMGWUlR1ANYtM
XgXy54c7MRc1g4lHAy79RWu74SBAc5toc5kMXsT1XLhL+0DMHbqH3yRykmOnxRAH
eg+Mx5xabsIhTSMvoO0d6khHxRxae7E7HDMVCglH07V4gfzgxicQmEMYV9Edy+zz
Hn64zIxB5JeJlz9QSNHi4ymO2JwFKE5jNzHXVu69yJvI7jemV9Z+FbgX2UMmnS3o
Z8ijEvQDrYVBNTYgjALKAfFwaZMPxDIkvJyuoTfWQEHIhtzfuJu7+DHKdMZPwArs
1gpdcCXJCGnTfABujwTFH+y1zVEyaxQ6l0zVqrmw70Snu9StW25HRfJ7DEPUpoEp
qehvT+8tHxiKu9d748NCc+AC+OY85NJ9CnV91xbamTRA1TJipS19/xKghe0Ns09q
hDmw9lBzJjBFuU4TuDqO3dguUlkdXyqaTTjEHVzPNTtddwD5J3BmaGrkRvOZRWy2
vYGriUWpqGQdTAOgEFmmaG0untviqsyYCbA+CIbvJm6X7CofsZvNXauiuHfCchGd
EeEQySpAjMCCdkGJ/KzbM7qT/2Dh0RoJ+i6JAzHtDVNy6UAl9zuWD3psr/8UPMQN
XlAV8VDOB2wP9KgudwofAhkcqpWE6A3qdeKGapdfP6BX+GSX425osPNfMjpo5pDK
FYuTq3hc44j8OcGCwZgvvvy1zU/S7rvNfikPOZiyEEc+EGUjLARE5Bonb3Tpq2M1
LELfVSApjcgDfQKzmKivHZXjiC+pPvE//crEUuPSTTxozi0/FvowbPX9PreRlRqb
itRQ4vtYxC7lmG+dYyLS6+FhzpOt0eJnPRYKQ7JQF+vf/VkMJ98OI8J9GXrjeHna
Z+Mu2fNgXddRb0o3SbBnqZYELWWH3bkus7kGmzbkh8gX4Rcp5xMxhUtO593JwhpT
cypc0IsfaL6Ul3XEeZgL3LaQFraHs5mIXcYfwxosHNmO3vM6JDa3cpgSbCrdV2Sf
zSFhSdunmZXJgU+r53BcYxPaaPOkNg+DQK1++NmhfCenSk06YkAmlHvXa/G1r2G+
MBIIaM7jAiTTFhbRwyN1/EFJMWTMWMxlBeMf3NXaG3yzRKz/xcawbvwdzh96fLqC
Ed4C7MuSpFYj5Nts3FfxPJ99/pSDctq18MJlNm5uIBXFgaKCPxprvJlav9OpLVOb
6hNuqZ59TN0Sljt3J3/0a1NLDpjV74udncbwRataWZoDBsLTb3SfiwcGqjuu5qD2
sw6OEtrRRd++oQ3kDJ9Tj3WvrtAobHyDblsBDnKfTYYRQ/U1QHx8vDDJ4qaLPDM+
p30KDuSqzodSSOxwnWyJqd2rX4RpNqXuxdhOV89tmrUiq5691Y9m+s9ESKyJKK/N
jf4/4BGRZSbxrnglnIToICN7gtTjy3Ca+hg9zkUU/NQ3bCzEWwniiig9+6d295A1
MCjU8cRBNaekfSt4S+T5+loWOQQEDbWwwfX6rUmdI8w95TWp6zICLQLrsNRTvX9B
WbXf3a409OK0qHTEfLi+cM0QgChq6/CZwQaJEyYOg+qnOtOXGNM52saEqwvT7iTw
MYTWEWYmiG4pH7ruySSES/jVuH7g39OknQHSCBhpd8PvNzWF6sSbZ3StquB2sTzP
NDfGdb1DypvOcF5bebphc/SGhpgIR88XI9q2dNXZPDwdDtnb3p5nx7so107FB2T0
0OnpDwhXIUdGxNYYvqDLHkcOo4tczo2iUGzfgIRC51PWe6zQFsxUhIYURwYkT068
ceMf1d7U0Uo77Nqs6zXkW3rBm/gsn08hcFm7IU1FnyAZg1B54DlTNe5vTHm19Vvy
HT7xZf2TgxFKRnjq+NVdCrv+qq348yfX7GrFiOv5NnOq5au66RzrFIPN3a3rNzny
xZx1vcJ7S/tpnCERUeuqa9I6/f7WN9WAYJMLqGEfHJqnM1PgAAksVDy1BGdAasXt
NFfCL1cthRIIINvwc+bpuDCWB86hVLOCU4ckDIJKp1CrIQJceSEVgzo8Q7uTIM4f
6Zxe+qqWHBmOH/crjiV12Zi8fAGrvQ9i6OhTqrRSq7+BY8UEwDdSPQhNopdKe+0r
HS46CoUioXD2+u5aA5abX7N1DeKuSSGAWXIiZuHvH8dVZdTVadXlOfvXJkQp+sUO
MmHwd1BS3eVZved4WB6UaBJ6k1tQGSA6OTeP2YY2ftzr8vs7bfQ5/rp6Pl425ONs
LHYo0mlDY061qfxO9NQ1k6DVA4aTRQ4udhdAgYcW1MQ2+iQ925AVylv1CLzbajZs
OZVQbx7+ZJaLQ9rF9F8EXb+MqJoqK5q16YI/Up+8Ace9tzVUInHVi6WpCQRyoU1V
ir7fPN5bMf0/4oPhxHwVLUQEHrz7b4fEWauRLXk4BUpGaHlsrJmEab4bf7EhLMQv
6NqT2lXh6w99KhO/thePba9CoH455Sr7Uf/WDuSznS+ngrkEQO43xQR7vdDrid7a
E4ME9Pvh6nDo5hACyxJjhy+GaIJEemuJSOd/ec6PgmvcfVv0VTWuY8bsTPn3B3xn
2rYqXKD/OMJWqyjWM9pI/QZAbvbc5jYp/sMZw1BFYHKEsra6LB+fR+kzMED2pF7v
Ot9wWpFGx6zSN/4hNSmO3aavOAlhFKQjEQC1jxBMC513n4GT7Pi3r92xiJOUylOR
k5E0l+PNnPuxThBPQcCVTYYalK3KfFakmzsI0aIUfeEGcdXlRzFkJ4rnGw3DtJMB
rSH+SDwYy9iB2GIup1tJD1r0HAnK1hrrNTTNv0TvSooOqC2WrLizYEmDtkBsn9ad
+MR48CGvXtbsCss3lN0+wP1TjSXuhfriMnLuoDjauozocfbJ6DSVTokVnvuJYJ9N
lUPFFAfxZGdGcLb9QyQSamBr7QxnOyNdaTwqgYXH1BV38a827X+SfdXKzujSheC2
E3vgXI4fxTW7cRqUBvwqTuXkQZQ2b/zhLhAh9jgEdnmLB9Oexj/RaD4rjm0fT6g3
J583m5y6nwo35bdeXL0IRNNCYvAbDWnD/mZdcCyLEyUEsILNkrN3tqyrSoWHgH15
W9y7JVuNs4S6EXhMGnSdKUQCrYdY+s92AHWh/txrGDu0EOd7B0plBXZZpH0Ab9O4
RBveD752a6whWS3aG7iD+gR4rUHJbrbqSMBaToS+Fg4L1jo1OKy6EZFiKqq+kXK3
7GurlC9Y1rNPjUDAuCreBTSPHysDVhVs6qluTBI4UmnfOawpCCUL0dqqeuNESoTy
dFV0Zvp4beKKz03I8lEwesQiXeoz3InD0U/8IL01XSlQduCysmbaS8QxQwklLepn
y790PpYgiVYWq5h6v7JiLL0MCgS2Ti8bPwBq6TxtsKpuVTHmXajVZOf8Zuw37fPK
tgc96LD4dUPsBN+Oar9EhdG5b10kzQv78A8zzMwuwB7Lfx32SOI19dG5yFDYy28N
a6LWRpI5A8IS3s88unw0Px1XnBcrOTTGo1wvW0SXZ1zNv+CDg2Fz/967JOYwgc6t
A+3kCBb3PsNRvdd+iUPHISbGjFB01ogZAh/A1v0L6SZOJ9QqqfjJpf3EYxiTRk1d
fiGneoT3HlmxDSh1sllElqfA5J+/Q8VdhE7ruHmqs+mey+KvRm4nwJEuRzJilGcm
u7CB2LBzkEIIa47MSkpdNGFiJVthqznQQtW0coGsleYc9uzrJ2teD394wy78xjxn
ca3+HrdTrJgVc5EPXDMXyNbIkP1HyCrALnNF819QKAjnsu9u1rMFeVnDqoOufAXP
dpYWuGmb/WE/KETHvQHEIV5walTeEvYN8aqPDuq8QWRvMDq8D7z+h7swMPrHraCh
WPttI02aYXS4hFElExqyXwoT8iFNYMne1NCpna7mcWG/1lN1dJw2A6ZWBig6G5ZL
hDrqlMtru2zgAcfYWZmYfkDswBfJydR7P/33VSCn/x43v8GyQVuWAiXw7otpEpiP
jTJXqjQDhN9lfizjRjpxLCklMFMVwf4TbAT4O1KvxhqGQ5pZv84lCFHe+1UkGap1
Vb/hpqQS+AfdbCw4/HIT4b3zwfBga5GFsWlbQTrnX4CP2s14UKtMorVFjJaKlQ3e
fgTr05mChAkUTVaRtvyhMEdxQjBD58zIlwsXowNRBMAOPGZyJ/jfF7q5NFXQNW1n
Pk8wLG0NoU2DGhV3xgbxWgMQx6mtHVD34GnyZokzgq7TWJdKgyricSgSSiQgSYNF
R2kMMeGoLzLZxpWKUN/d/os4PshXEwvOvwE/b4nVY/5sMwknAjpAuTvEcg2erEn6
pMgsjNDwVGLigTlHBAAGaSoLCCsYEtIix5rdwNBwrUSSexM9zVLtFTKNafoGQbe7
e10kMyHlR20MfpcZl2+vNOZgXJ5eFAHcijfu3JTLwR+q9PISR9E5ldCg8XezS/Ob
FJbFlEfexv4N3d23zplIDL2FY9NYeyrgI226iOyKNS9LeGqoPHLVEeXEAfl2CSSI
0YRLy7U0Iu3+BMQQhYzunzZjb43ezxwMb0MzNANJLBpVQlCiokArGJQOPc5XR+jE
4DM94Nar+OlV47BzedB/2k3E0Fe5HtcmbaiQB+pu3+GU65jNCaptbQbzRaNn2eFy
kUl/q8M5cQQ1kon8cFIZ9Exz7IhNSXQDlxGi9n4AfBy0wWOnfdXEsf8BiU6+G7HG
MjdacTcXx8fjwSs1pXb/x2JJGpeYyjHuNErEfIJn4cAt/+1uRFNReslev0uddcI1
Z7v3nuRKNEIg44a8+97ZUoWJVYPfIYk0aSpgGi61AtenODQHDPSN0DIQKzg0BRoZ
cyW9EFXNkj8wdQD1gKLHKE8dZAH/b16y7Ejl3IhoO8ym6K1ye+h+7sID9B0F+BbN
ZpohDZTE1FywaXHLHCJHKR7cpZWoYl3zwYL63qknLO9ENhsTjtdtgWxMOIyza/ui
yW5fECXy2kX36jNPlG8hGuF3oxeE/EBnQ9lOkFJdo4PMjIh09jQsEtBg2EHQ8YG7
/uKpW8kXEQ/TWBOSINGMxVr2tcVOVzplSyOMQuGzrZLekN3wSLcs5LTBp5bWwaRG
c6wGCNXy8Tl7UGUP/0A9XraqBRbovk98Gx2klw4dnYCfvurmyBo0EM3B3Ow1jAwh
1/RUG9RAHY3P4PmAwP1DpsFwjed2b+FReqhunxvRRzznXw4Fwa8kL6RaSnArcVAa
5YBTNMd8NLJiiKHt5zyBSRXcmNrCBKZG0x0COw2tgF+z9c6ZSu9fuuxj7WvkvJEy
XlRxc6Nnvo1a2viSEEj/TmzXBHcuGWe6/t7Cmp8gvMJGCo8uB9Lv7/HH1bYiXj/w
N9MicCnHkER7/sAtLOIPZSFZIs0neKv6lwJJjXvLqyKmujWWITeBieV/UHu5zHDo
+Yj8i6HKi3RMHEUkwDm4VoMxrcYtoYlPPNKD1sG2UtbO/4YBYTItxaTSlWNvgw2w
Vfm8/H6DCxHUpCaYIdOol/ay8K0ZWnAbQbDRvP3nujVZClxuIABOJUKcGeFOfgz0
Yg0ohcONeniFfmEALm6tKa7nq+moigrLLKJ/2z3CV0ZU10tpqu5coQXKIaz/DjMV
HLcWWgf6LdI34M1hG1hwhFEele8hqNfl/TKMt0PZXyNN8zH3sM6qaIGd5JYUogNP
gBj0ASVI08JJQB5X2v8152M+7dhrczwKeWqwnAmlh87ojDTO1CadmK20U/JYV04I
3Lk0Gnf9p9I35pL16SiIa2/aMHgNsPxCaMyabRhateYUhlIk21aDS2FwQ6j+JQ+J
cZkkuPr3DnfywHpcQXzwnuFIe9FYBRS12pXoZQuAmRPiBqevkQDpKsqDKCArPkJX
GDA64c4sZCeobj745ahsyZBy8eZc85VfeoAPi928oLqOIHCovbfuZNylolPW7mbe
NokAs4CaHitdTYZIP1IYYxrFgwHf3S82utQeDt49nkCITdx8p73GV7K4l47cARvp
w+yDM3yEAuzucHRHI899umMGMMt7N2bQHBR0qHF0//IRWsbBDDnxA+oh0KJ943lN
6rMFF4DhA8X4ju0FRxotCxTU2N9U5+zvNyEakZ6AQIJo7mf2Vi9Bhn6BRR7B1JBY
32c1FRKtEXKaujwcCw4ptgXKZgn623dPauSLkwx1fYxvbiNJqmH8XIxd/D1LDu/g
B36hV1gBMM0Pugp3GxVBSD+3pwnlrLo43fY9k+zH6jcKVkFsD3b61g+7n9Uy0Q07
sQySy4Aa/CVLvACxXfa1lhFkF1z7yoV6ai/O9MEWBs3umAWsGa/fuVXNpFKGEL0M
xItBANJZfEsFbvRnl5l5iV70uT9nCIvJf1E1Wy7enLbO2Itct1W9OSTuZL8LTcu6
e2iYQ6W6dDaMuI9CQwUQXMHy7/u+H9b8CJ7CD76mUO8L2osGRzgc/Jm9HdlSjtCl
SNacKksdsvKzqUWCZi45ZN66aSaoqrP8fTh5NTnzMVYCvnDYREMTikqIneer1s/m
woC2Hfw2yf/iduXVc8V6iAdzeMxElnjeCU2SGvp9dtKjve9XcTPcwcGiKFAD2O/9
cncioZr0jC7IsjEFI8mJqQxePr1puxuxu61BrWWGKmAFWWMuUgAl1ze97yUD5QNA
RVFQ9RpzNYuDNl8ZBIrwfaFZM44pqfxZ3eDHYh+pm5pBnkauenf1ETE21sux8aPN
fZC5O13XnEqvybev50AaN7jYMFnipAguyrZksJFcGBm8MsyHKOqJqGNl49+JnuvO
fhS4k5Cb3/cdvzwR66/qMebsR6j8Ju77iGiiQPVOIJiIi4EpEBJB99ldyn6uEUv+
PXi+nBuORTWekC5jVicoTlWrdQrjPn4e2G/sSa1tFtj2ThPKrAcNa5lq3hX7Yq7i
DkdMqqRt4g/HC6abL8tIitZEh3N6AmqBFSbi8UmBbES0bEAsTFhjNLARAYeuHGmo
62K7mV4dYfaSR+ILi9vfL25qhmgOlOS9wOtuBoJO/4ee2yZL3Y2K9p5+rWJ0X7dr
9I0x7HN1ZZFVMJmYmKCWnCKSA3NXXaModGtgTjUnwrqWka47C0MHkXaofIfEMFaK
1ZBdrXzFF1+e1IUDIgYlOJsk2LoMhVRRyoW7jqqM0xpr3pFOxlEcrsZAnBxWKg6Z
cnNUG0MjhgoYQEAIn/IDg9S4hA/N0YrqYxXS3BL+ely/7u138/NbLAAuRJRXA+TL
PDPuZFge2HU5pZbRuds5ig7DHHl0eUrBwYTx71aZO4WxrfWqSTY22FGK0CPgEzdG
2/FBxoMwzA2YogZMomAdwRl0ACiBmjzLLaD5vqb2EMtsyGSdpJxM86DFDEqKI1nC
5N9pOCU5RmWOa5U5mUU1NBJYcIxjgU2lEVSNVqb4IB0xQEe5VmfrG3bv5v50k03j
jR36Ux1KKZX9egFT7ru1YrTylb7z6SQkrrX0fZU9n7sFhE3/1gZSugZaTj89AW3E
ix4JfmNh8ZLwr4aNgYFMmP/4SfAX8uvVGc0dA12kIDXgQXT3TEE0eH9taRe/eCVE
Q8aMNyNys6OkrcHtTYBYVvXZthuSMcD1pVYJIJUK1IJsTuGjAh5qyEx/h29//y+I
HVMaRPCcBPZ5DYxjFllC68ItalvaBf+Ul22dcVpdlFCdZsEeRfeqrf5dct9I0Mrf
gKnVp0xdTlM9i4A5+BbiUEaBNa7nk8ypYOV0ft1xAvdu4WzNKf30AcAw2bCN+8BQ
xVEngah7HIEqL+fz+Lu0+SirSWbEFF/LXygCDjKk73YaCaBInWLdZ9K7R2mobzut
Jx3YVHCv5cJYVl1HT28HU51KGvQztVckIvaSJcw5WLiJ8/YAGdec0LzZ+5Khswir
Izl5SVoVBchMY98UrXJCqEOC0cjrwwTROhUouFM0yaM1CKk82cA2MhHtdkaDojCI
InIG9GbkwrhbIWMRWZIBdFarsfO03ZF17EwVB8TuU2ZcAHlUPIsIp46+x+MK+VRI
OPJXoJNXOhLlLuzu+WUAn5dqr3sH1FmxWHc8uxayEt8wSMlqNNCtzI/2rHsWUB/F
lTx4Ls1Vq+8vUOWRc69+FZSYoMwB1/+cJ+aDRFRKQGS43U+lZQa+h9YI0LN+qiHK
7UwUGtd8ck6ZPjX3u0UnyDEvJdafO0pZblJsP8PnxXhQJUC3zBDoi6O4GAj6HqTO
2d1UQ7wRxQ6vzuGDVNItLDK143HSrYfcNj4/7HjUL74DrRfluswrO6vGWoVeUqQd
IJYJmB0Axh5QgfIXfb62bIxD2aR/VzMHVHcrSohnJ5Z4VFeHVGs2YNCS8zgN2oun
Gn7VryQ8nk5NiCLnZxClFxX9EU2PVJNgwdwJGJxlfEp4WNeqT3V51M0dVrcfFAiT
SNTQKRg+TLdPTWWicXLxTeqqppK6CpFvuVEtXMofWoPFhSLB4EgLJaGb/vw40nTe
DOqtDgp8XN7i4iDy+wWGz3b6nzg8Xy9jsQHJ0oCiu65ES/7oshb/4Q2cuLPkgYQc
G0i7wVwcDa04Q0BjqJT0xr0Z1YiC6uxI+UdFJQPsIA7AdjrICfFbOe/jhPMmDd30
2LQ+sqUbCJHHU5rtaB3GNEWF1sNcHaQh7Gv3yDE/UNYzdyS4a1WqVMnScUBc+3eJ
fwAT0ndhXtAtbiV7QW1RqqNd9ew9AND5DyzsJbY692ilVFqgDHdsNsE7Sov3uhit
R2PN7X/d89qHc+W1sA9z4X4q3Hv95vaWGWJtm2GFTUa8/5hS82oUeGSfVz2ftvFb
qSx4Gh9r+PPP6Ekn3J+Ie7x9JaB30gR0NzzenuhaPX7TTRhOpNWkZ00NCJaxbkty
p34OEs4xDPZLhRBUIMNvyjcvfQqvfUXg41TswZGJcq9llKMBhyhmiu3G0JzzYVl3
NuJ9h/P8/+lBeEeDU2h+P1ao8V521eD47DONXRjzJGvW68AOY/7h5ZVvgwJfd2rO
wUjBO414pvAx57czKQIvwwM31ks+zALzqlMMgCqdNjPMjart3q5BJSyEoXK2ecXN
uryPnOuAdFNDKzPdMzUr6LVxkUGK0Lv5rvQ9/+R0ZT5jJUCUtyhUmRKMjcYHLXRj
x0bxQdvo6xuzngRaYS7V/uYpNkOTH9bgrqUlXZ/Q6cHL7pm0nYZzrFt5mUcpNXWr
nwpoMiyNPXXCH48cpg7+BM0xz+7Bv2zy6aEefvc/LiKcjq3cdj5cODcr7DaeZ+Tx
oeMlVHe6989cKIKDOuBzzcGrRqE5xZt31uJ3ElgkFeJUPK+gwsQ1EwLgbcwFKtFT
zSnnDlBj+tBBosjygoPzrhAvYf4DiqIubZbnGO+ZibgGseZtAoIrfTdLucTgL9dv
xVsTbTipc3pOJFF9aXHWeBuU5pN7H6pElZD1XfPb7tiZjl+y4OsOhklPnV1qqud3
quWqRocngXgqhR8mS4p1MRh311TuKLb4QHh3OKetSjQYYgtaEfQC7vPVypG+kxwP
PSvKD8/bL7ImTKYKnMG8CdSVeC5Jg8YQu75m2AkRts3xwYmRWbVvOT/BYRy8F171
srfKz6K/MCTVxtLP373mLXbt+ovKHwav/KqdB2Afawyec3BkKxNhVA25EGbohnd9
OgVSN2QY883YG3W+GdWkxf6wB5jmnthMg0gBJH4+MAIosJNL6vOprUeN1CjRlx/s
OzapVRdD4b7eG75n4emvS78p+Uz7/WxohGjAFHpVoJwjGyndDBULDz0NsGQgQio+
KrGLrLByTqRhJcfLCJDt119MUS9kSSDfL7hQ0M1IgCeS/sBIKGsoAeffocFTBrBg
boqH61f0y68WdWkGFce8TioDkXCqXbDKb5Kl6DNZOmeYy5mGPTpFIgpKjaQ33bwT
NaskwJ1CvAO5yX8eozzd6srbSbv+DczD7iW1Gzf4TgsyZQ+5Z83YXKGLf2toOvAc
eYQ9f4AHmY8G5TYUPbOO8hxGv440Oe8/TLjvaJNPXqnZXUUxEDMSOvln0VYO29cr
32fidWpb+YZjWcmOSl7n0y76wi6Zk4OxGB6pcHMV19A7mJIIVRxlkrc3k7RMT27A
ivGN+/PSN+KO6LnNRu40AFJJOp+b7pVWLQnh9QmqgiEaLfY64zfnq8QmVKGcJ1qn
yBOpSTZbo7/O+vN4tjrCNpJXyGb8EchSK3XdGDpOUNmppnpUaO0N5QJSSX/mkTM/
BjLmw/YUe1LQF6RXcrYontLiO8gIibDdI+Hn4OpEyHmAOKTGLbykZVRxtbuyBNH5
O8P4hmLO/HkRztwiu3/inW5vSmZWxNnndi98E25CkNexPqENHY8DQWexu76o/6FS
wd9wSRGk0/WUfmy5fWsJOp9lA2gpmKr8qWu2rIaYyCDzm5CQw/G9IQPBypU1K89n
B+LKcCY8UhQYFzEb11H+muqMIv8zgjD5x1oyv8Jzomnrn4DuRMAmkIayZG68avZZ
4sFaF1wMOLRpvdE+seGjK+giVfc1pxsyntt7B16oWAKgLV0g4HjOyRJes2blyf9z
G/paNVY5XYf120appE2a5Yhihvv6i0La/cniZKjt+UlcKMVG48m/Z1zUjj7cNN5a
WmbL56TG51wAkoJjUY9rgdTD9BP6yJPOervK7it/vGH30avMQtqmRjgefjh6CrFg
+mbtE83FjAUqDICp0NPJ0bJWudTCcUl8eQhPOan8p20eliPxyFpZZMBso4ZaHMd8
VlH6U7msUTobrhj0jbC3GwattkI4rHEApdJTsENXkAjan+22qeZfr8NBnLq5iiSz
koQYo6Sxp4YAU7noM85o1qhi1+PrwCKFRJflv9JlmecA305cwXCDtOsItAnZ72Mm
c6RPd6081PglffDgVPZCSzl3NroTiPbGRf78bN/2peWwapxq0CIxbb/YHbQ5CbFm
bAL++6Cgjk0ecqZk3NWqnpoD42ixSMmiIrOnwTlXaVtFD94yo89RV8vebkzN+HhZ
Nk+Qypm7mXenFTKRNimRoRFwzczjPWz83ka1NhYBhm68/uq3lkhlofISq42Udxe2
UIR47pwmR/sKqGpCqVBYLm2ukgufxzEiZa1uHj5go0rSDMz9BpqexVu4CGNLUQmB
MKXkSEjO8vMu6pRk+8z5vdCXi6hZ02gws3JeYMGEvty8Ns2QCzKm2gf1xyyNBiSU
QbptsPBZ90rtOuxFzdR3KBTqaRRLpYouwKMGEkOVgrV1KjnyU76KRRy/H5o2Qyr6
PVGPfPokXsw20U+aifKjTlXA7nE5gS9GR1EA3akFgnGwIRIDAb/VWTjsdMtnl8So
P4kJITVSX9zhi4JMctsn3BAjvkCavSGIuf2YXOkCtAXwzf51QN1qHmRcNoqny4ur
zKBUQrGyyLO7UM9Sdk0Ph2hASq2RsUq1UjFAEHqKfnyOoYNw74TdA1edMYbDn3Lz
6u0Se1CHAPbmW4Mr7zRcu85TJym37PVCLJ08LneNhzdJ/8G3ZVHEe6TonXKupw1S
RmnBug/xOqQn89eYZ8tLgSmiuh7llYd1SqIo5dwjtI/pCGf8P0lLSCG83rYiLat0
2MML/cBGJfOOABglzN9fxCUimYFlchz7xh4K4DL4QZeJsCh/eqFtNE6IjyvHlJsN
bLA9VxLNp4QJj+nfmdgNnVPwyNVMzWlTMiEZrYSqofxPGnn1sfpRI1kFi94OeH/K
vyimE04L9jXDzB8W2uWwf8tPuBgwOn1Wa5UXFVb18h0ey31Z4tuvj4kFHRJdyDsK
SPpBq5VT9lMvgk6Ajzk0O07HthZD2m8HRYxbjFkdSLznMMCM90z0AW3DTosm3maQ
cyn52cUiGTzbxO7kA/gOx2yA72gQtFC7uWcC/md7zAR3xTN+4GgiljK3XzFBmo3B
cJyoXsVZMBwHh2EhEXP56eu4UK8CcuF3cFqT5OTZ4LdUlgWDbv488NYa9elgNCtJ
2ERWJDQVjk4OsaJDZ2qRdjkv4ErjGMplGJ49iONrq97VUYgpPEOJ1SW1ixQTlLP+
3p1rv3vA2OG6xOS2ejtI2g47dP+T/aSE3rCQ4YySAAEijPqT74x/UrVoUCfCASVR
f/4SIByT8yXxAH439fXUoMSlqFKjALa2TKWNUCjze84w85FEGATCtQTzptnfvnBs
vYHbcZXerzyo4DQI8HmbDJ8vp29POYdClNmVVLCyCV8N5DYhnGOM4bUznuxh0mCo
caMaEHEwZSt2sYmpnqaJ8hFecKU+4hVeYtYIwTreKQxXr/2Wv5hI6bwBk+FSRWSi
BEd5X04vBcnyrWbF0X30f5j9aUBTxhbHtw3qmdSPRyXmCxvTNyAinsjUoW2U2Hk+
gXPytsbXLI9SQYii/LYoXjrgufY1o54G4q0QCe9KhW4KjTwdIRlB+Q4XCb47zyVY
J7WTvtktZxpyl3tueXk8GRxLMRmaafSWNz4S66WPiH6NRa9BBQeHRC3yFj4vVYpI
7wBy48r0NtasUWVI5CRByOzYkxKF/YjmEZwR3RJsuaPbXsfJuG/ejoPWgdy0FnDN
Ova16VN4Cic7v8vqF0iyCl8iXGJZA+efgBABAwZDSfm7r8FFzfPyJGO932mQFd/y
S5WtXqqNyvmoRTk9Tc824LkqHNkd/o+MwQIh3ZqUNdZz2tpYFnsUz2slq7zHqeRO
T+td5WgqH2esiFtVyXa0vlrJnoh2w8BkUdx3V3WtQOr3AwQ3opL92w/Tg3tSTaqA
Wzn1ENK7Vfpwb0Wx46n3l3rPmjiMe7n5kgVthwySPi8VstYCp9I5y8euVgjGFIdF
adzG2qif95veGGLeOLFsR1VXPfDxBCHgy9WZNurDnw09S6bHMvPy1JY1+X7Xe0B2
YxQH43mVtL22GOiN9/yLtlw8vRlSKwMmSu9pTgantbgSaI4FihQAteZzKACLQ7JE
I39/+7j25yhJ2VwXAeXhlBS5bNbsNTlbbBoNAyC52pu0D9lk3S/ZEQ1zlxo/JzmF
jj65lyH+HICaRk6yWEL8wS5oT4pLbh+QbMw3RILk6RCPDaKLurmKFYbVD4iD3l/8
dqktSEAA76i4mlpLIUwa+U4cDfiKzA2yD049P04jeM9Kt4yH8RSI30iMv4rGVOsd
3zkiwmIR3qH9KvUgZiFa3Ib32UTxSWbQZzMcG9kROUnOq4FZKL1HVXU02b6RxCMe
Ls8szOsM/Q8NarZJeIBv3ryv+RQ6Hu3JB/c9gcFSLuQ8tpa2BiG/3N+Go6znAgHk
r+/ZjB0l6GC4Z6GbMPLE5emcnjXPj1bzyLGIo6zYFp17uHi1FFGWRBSZp4J1Uu3X
9VMxznHzG4SGf7h+gb39nCyAfO3NLXse9q1LqBNLwSyfBElcQBDHorqMl6N7DHtG
BBTznvPOKeXkocCJaRL9FdbOa/78/toVat68CmziKxLHZ0oQLbIvQJWXB9qpy22l
W59fVEnFPjd9UWqvhwZJJDKr4BR5fHdRgQmaLVSl30wjCJPUV3RfwlH16u/eDJlU
S66jfnM3vgPB1Q6YM5baUFy7BXlzNo88s0CLdUS8U8r4j07p5d7BdTaYbnkRWOnV
3wXdVKHpqmVRql6kpMUsqKZhcgXAvH0g03obxfzqyA27cG2zBm6lCTL3qqpjARuK
0ZZ1zgFsS7B/WPhaW/0+2tgq7uu/j3FlWfv+ndpIW6gPUN8wjbIYIldfQCISE8Gc
4MFidkM0JoIFOvUhZ6N4UD93dHaclFxuV/4jHPf4Ow6eXqVsiy1st+1mX6moV4m7
jKczvcPhgmnbQYQ41/FtB060rsxNKtSi84PMkTClvCJaA/n60P0kCg7bLspJT8cQ
Cc6e+NB2jvHgdxacIFPhMzgx/xqn1HVbOUAkBU5XjUY9004INEnoiySMAXQUTQwv
uUV3lSWDO5O/AhUlZHKsBwHdO5sUE/tGigcwfbuixjcWnYbo6OqdFzcpzt6S77gY
KdlQaNC24iW3CrEviFC2dwL/nzEbX8hH6sn+yARhnSxmz0ZkaiR38TmeT6LtJemn
iwkmYTF0s/82IIkcabi8/8sojQluOVL3YJvSWs8/EON6HkAD36EUHCUBAR1Ip6S5
Ab5Qg74+M/g/Bq2VKOI4jRNN+3uXenspiY7750iakc4f8v3SKrGXr9VuZ9ayskYt
raqxGr50obVOp58SCId+Kb49Hek5bD44cgGVyrNESBb1fsjZbn+fk3aLx+PQ+EwN
OtatZuxKlQURKp7J/h3D22vqNq6SXEFkS2WmXvKQijJK1ySLLYSWPa6VILho4e6W
3wBOtSSBZuS88d4lsj5Xnk7GwV7BO1nOg2/3l8daNGv4Micvbn2aPeYZ2UvjWwKh
KqIxaB7+FAmmCnz/ZIFxQkl/vW4vGcGPDoUMMxr5vxuoIugQHenk6pPwLqliSjTj
az8Zo79YtLqsIPFSdJudG57pmoUfbOFlzLg3f1sXGpBZQBXKp/m5LNQmgfuV3T6i
nDdS2BAy+7aZVqqfNgSn+CfnVbYJgYT+p+okTAe9poiNAwpfmDQZo/ghLHWVnkQP
97mZU6qq/2APo6znTTCbW7gl5pxtQfMGbuVUFMXCRzH1Ki8sr5s3ebm6xa7KCurR
1ndKHIolxFQMdN/qXs6CYQB38erhf4QUVpsZbx3q4po/60KjKF233p0iavQLt5Ag
F1Mpwot8M3k3v37cP919eiqKs0m2ki6sCAI7gsb6jtVFpyEXm4lfA/f65X+Iu/Um
GlWqiXn+JcAHVwRfVnFzTnL9ScG8g2Ru5A/9wJHmDX1XyYlLBdELo5F6my1Pkvp+
YdsAOrljJTwQKhbPgWeVKaWzmjO7E8OAApzj3l87J9qbbOGcbYfXh7ked3Kkx4tp
nQUyeqT3TejQ6B+Qf0iKnJepv8JpVI17kYcFtE9IBU9P49slCLTz/CjbJ9UUjtSX
1zDoi4qsbWuMVrjNIKZ4YaApumzMzODLV3k/eiUYNWaHfQ2l5GXmotYUgy/e5GWu
nz3QmyhBYKcWINC24p+1GHZB2QiLGylR1ANseUY+E8hYjB5WtAmV7CoUCdMjS8tU
3NSXSg3aSNP1Gl+iz2B0ewb8jhrWlYllog1MffhqhS6qJbRorNHH4b3lj4lfXUuY
JElW84XCFyNMaxoCST7HdE5DkLi7oQWfkfwSmhTP+ZFxljbKaouMAHXL6N3RLehU
wJCUOmm6AZNiUZHpx0bOqer1H0zscgRCR1atSg/6v3B/EodqsusOOGDOb/oUz/zW
ygmrPH+t9t72mMfiFnbdqfSmupj46Yjwi3V9S9ZgWHUrZYNJoNqispMKxzu8niAI
jmY45BrkNryqqIQ8HjX4iUxI61VyQ7tZRB8XnLkQeU2eW0qVgIYKLbtYYt7ZzizL
eE9GfzSV3RhFfksU6MCMmFYMMWASMnT342S/ozXr1aWm5I9qEkZQyKTHHNp81dIa
b0uiRTtOJzwIvA7WJDD+poi3JHEvZSTf4pe1tAvr4VACVqBaTXBZN5UOE4FZKbCd
/Y1M2cw8Oog3QqGFJGcn8yhvyFi458BK7Zfk9H4bpKBDjvxxSUUBiMJkP0JQdZqf
Lq+cfrulNHVYaB2iplBVCfCGP0Vx4Hjtm2AVEfWCUguT3eYTMzr++LZc7IAR9BJc
gVrYharCBNjBHhbLvG6SUhug1caEBVTOo5+mfYInG/NdDrI2iq9MeZQhwWCV1aJe
iOl9FfMoXHbhD/e6DjsdD1B8XGxweKDTxYcp0e8oKkrTpknglzK+FlvwfEPlcP3z
ioWkFI/MNiU9CBfrSuPi8rXs0mutzQ1uLQoIRFg+N0Sily/w4UPZ7FrN78aveSJT
hOM1OCKPf1XRWFxX28HUxDo++2NbUpL6EtrPiV5bu57Wgod5UgwbPXmrv2vFBqR8
lHUuMoYPijAnzR+j2sAlPhcMOeowyeX4Sek2+b4cvTGD+PntnH6CtLlLipTBf9CE
3rpEK9uay3Iugh7twfmTxw0wfvrPeIf/SIgtOplOY6N8J2XGyX0ZG7BUTP7pWErH
2pMvrMruAHKSFt+ci3WgbS/Eh9v5+jRPbNedT8cef8TYti7WywMYOx+0AFefjxXd
99ibtjFueax0fF74VOUccKS9sBd9zw92+iXg+re0jAE3QBzST/3+cVNbpvbSxk/q
jS1z/x5Nt5OE11scdHZeudQtEkK1pnTPTI3DXclRg+ipHnw7qabN+voVXKiX8Bx+
WnmvYp0sKlVgeCX30nl3eKkkyraEmKBJA18k3+hyqugAKPX8mL5Tgc5Sa2Oqav28
J1J+D6+YwU+05oCrtBefkQfTFXufRXUVZ1u0T/NoXmeXDuPZ6nr6dxrdYRVGAW2k
WFjgqNwjuebGfAJv4H2YxwekjHfvPXHF79hZgDCohtWFz5od9NX20aPwYesryS8r
dr2mszXqiB6S7Vd6+xFhhAkGXR4XrU0LPOKQsJcSMWgDLdoCAWm+e2VAtmKAhUkr
WVJQjicZoF+6fvNPrvxk7DyKJhlAedik78+LvTgLyZsyM4oavLnxAqHaF8uEWLiX
0nBNhdhUyxX8hv9+yubOgoORQW38gdtU9Li7e/3FJQGVEJBVzoklHfHUEPCIU5L/
ghpCQc/HrsRspYi5mFrIHrJsEUfobEoBsILkV7/bTohfm1Ji/BcnzvUyxmspOGzG
p0MgHjFf1cgHGXglu0dV9unLRraqI5qQfYKOQwuJKbwPG0tH+nF2HmStFz+2c1/5
5wSoEeCHwSqxb3KW4UqV/zSNVYk71PzrBTldobmB6JbR+vBLOa69obirJWqNC7KP
bkj2cuxHCk7ZZaV83zZ4IoVr1OPLVguaqgVM8YR8TArSlfYsEU1z1YWff4FMU9KF
lQirREPKoJkwhaSM1Ub0UjcGejNTSxnMQHnLzvbJp0bAJs63M6yNhfUVt8PyedzI
VQpLj0Zm7qA2LI9/ZJYqYlv3HidtYzlMJqUrAu5GFPwpl1d+AAb1P9dmu4KiQNQz
VSt5yIznyvTOnctWBriVU3wubbgxR+QymtWNP8AH6QcTdWpGkJYfWKkdk+656cWq
vaYtDXD2GkeO68RopddtyTn+r2bvVR+EHRzrZggnBSe3+cErAFrKIRC3NkQ3qaIk
pxY8jKLMSAs1V7ZxlsQqtl8lF6iNUU8+tmeVhzWqVo/J2eQuGyQNKtTqUsH0lsP5
6dMSG3aW96J5GVcYi0P0aAYzPItqD9Gr7w4g5tj8U1Lx3jgvELHTmZFtJYsv0+Ds
9IWDo/FcRWnHUY5PxBfalTFTVbqvgXXH0mpSNHz/v9KMucsd+GEPOtXL4gAHmrsj
xC+ez9EjsqVq4LNOGCqWYA8lYBs14txpKo71BsOwsEZDoH67893ldeLWNB07Z8pM
Vq177tlcV5PHWPkSb6d5xgL5D541hUkeucJMUIZWq3LCs/eUCGDgkyOa+UpmvmxW
nCXYTqKGN5EZkWOYgRaH1xAjJ3RxxSHtbRl5vr5aMwCfGlCxGQtyXaPwkn8l4KqJ
1kveneiVgTXz4D4tO2oOhy9uFz1HKbrUm/UWQwuKgcQou3vtyyhmH1Sjs+czACvZ
1WDzj0QSrxcTiR8AdUAYOSM0vNV9tqvdR+3aP7kaSHO/z3EKm/VMXO1PaosrSlmA
dHF03gsojLCGmCNBLenrFPIW/l+xWYecydJy7zZ2YXl6iC9iQc8OfQ4+PCdGNCQw
zQ5D+pJbnYtxGjxWFMc7FzW9n9FijSlHpuDqpNWHh/MbhvxsK/vBz5CJzatAXHHQ
iwe4K3Ix+lm9qIXk3DJ8IG2iizs0iEjGKZTI06GY5RZho6bguqVpzsjRZ/AmG7go
GUUJ59Vp+3eTFelvcZqspPRRC7DuPbYl1o4FT498jXKcRVGJHaA6q1sJ69SCt+t5
xv1P2ElfUbtTzhwhjDXt+DpjOfdcQlcAa0AFpZENpmmVfb8yL1+q+UfUiICnF6CO
xSH7CmkJx0GBQI60kFXs3TIJDlYmPxq6ESrxH3V6tLhRZqwCmb0Eo+w4qtHIvOip
b0MFgPMnYElZt+j+WwiWYmnkoheYKAPHQfXFjKeaSH6Bu7kC3XqtG6F8Ujyt5Z57
vZVHAuAnri6lxhxlJubakFGySMZHusLBsmb66vyxuYYBzf/FUxzkXwKdBZ+QgRqk
XxVMGm3+UO1tvV48rA9BRRgeAiy18XJOzrUyphWfedpEbq0ZcNVY4Be06ouzQedZ
kphkHD8U8Ocju+4Xjuvr/zWMumEEPU/XJAcgjD6YMRbNDsenKm8jKdXYJ0KCgqgD
lr8QyK5w0QqTnBXgg/YnDENHJ5v3dGasvvVbDzGJSgVCQNghU0a+3leOZx50z1YQ
Jr8FzQnPSuOl9aphdXiRiSQMr3zkHN+dwJJnaT6xKZOHycSxNddZ0ODby99swSbH
7NHDDjJeonX1oYjR46P9GjeG0m+3wk6G23Nl8kXCE0Dk2eKF0KZf5AAHsNSeGg0o
/r1saFVZ8mvKIH3BDcpwXwN/3HN8XmK6aiNnI75r1T9dtPrkQXbcxPPhzuKGtDM2
wGwLkF94b/ZuBPcqArE+KhXu7Y9VtZCcd0aJHFp4AYkWFcmKq19ceKeQMGorAKgi
QM/s/eO3eiOdEjgPDj3l5xaRr6q8OlrB7c9GTk8/xzKGDKBlXsUpNEIBdnxd9ELj
3T1jGR/dII1JHP6INCbnt0gumo7Tt/iVcwGfIRNBmrLTmqQVWlDMdODnQ9oIVyBv
PCe0LWoO4CtPatcKWNFC5zgouhHP3WOG4orKgfrjMAjqq+yPXOd2R0RZ6WaTtHIO
6I3wepT3Y6m93ev8Ozf+ADoSJLzKWpuHnUMnMUqO9JxkUuwY2Y4pB38N4IOvSCG2
SIbE/yETg4PcFr//Lux/+gJuEvg+vlTaVlev8KRLINa0+2Hs5MVkwGWfOck6aGpj
nLOQ2LADUJnrUj8aNPrPIjKhSMBBGJeVhl4Cct2uSck2JhBwZk3uh229wFmmQJx7
9Xo6sqU8BHGCN8Z6QJvw7XjRBE2YYH7gk7BUKdNhNmQi1NGhJZbCbDLsrrF+Nqhj
qvwjSPzC1Ua8fMje40Q/6i3n4ty4G4HRi4NQNHOLLFyL2jYHeW66mdoD6xctCDlx
eHkGHyfObm4KrJiSsiEQayJOjt8Y8n++tagZDao6ztCioMWTO2ld9nsy0alr2+W2
mZ1Ay9mFvkyCKvkZsjm78cluBwFUswHzR87AL/I+LDh6TZ0U7vgRtEMtTHkiS8kg
zFOsL9Z6wxzpXxUg1+1u3Z/5GIh5EJfaPxzPfB+pQH0ewheJQ/ML8qb7UolpH5AN
lTM2D4z/pBPr0XegfmDV69z3xxT6mDtS1RgmIbGpMJG5hvBdQ4tuJQwklqHW0bbu
2skLxuWri2rZPQNBZ+/3VqZ+uYi0LtCBut4mpBZPBVY1g4846fMZKykwQDw0u3E8
DtKBtjFdulN/A8VcpJfTjfo65V6zMnB5pk/GiyXgQZOrwAHIBi41AzPPWqY0syqa
/UiDgCJFLspuVB4f6jtKnPEtiIO+7+z5WaGihazCLE6me1h/YW7bWkctxbYKVU73
xuJmCrw6h1pgLIafWDpbA21Cfvq+1U4j68GjGEYUfrToAzAUbpNmLsbYHIRubv/3
PVE7S1Z5MtEOJ9lx5O6IrEQ5dqiIDLExcfDkaZCF4fjtrEm5Vehmosur+qY9K4G+
S09m4xzqRc1TrqxkTY2uZuwvcVQ+w1btUt9oGts28mcizwe3Jim2ctfcrWvijV8/
mhVUKEy4AlZnERWCqfXq+Kl6DM1xGAYdZ9vEmZKHJSD/2ro+JmwBYDUkphFFlDjq
OAvn3JHKq+MdlRMe8YLo4FG8PAv4UlHQNZh6NT36Z1XzBx4o5VPt0H3ZaNv3eZ0+
CrUy65L1jxGfmNhE/4nkSMgrMgOpcHPWBIKjSKJPWjpmmtX1duKbVb21u0YPCUFI
fX1V89Dllm4PwI0oL90ikjmXKQvmoQhFv9FWcCUciFPWLMbEJ4WEe6rqn8EElJtU
8ZflRF5+3Kvd5EQFZ2OrOFlbWSCChRioesN1vaFlNdG3hv5bpZZ3i94ykD2cZ2Tl
oJTFADKTh5KI/akE7+MGgB0wtFlZAbpazVebUwxsjR4FQ1ppWc7uI6kbJnEJuJti
zePKIFTUAG6oRRlNLNgVVqH5OD1sn3TFlEUTic+59rZZhkKiK0TgRW6jOP4BWGrC
z8ICVqTEfQLHgo/0No0XCbKoHW+fgIHRgCo/cccD2QJ/btmvUGt/AVxIu5/amnaH
JmxFjuvTTXWu/zPAVgM7kC28nBj/CT3iaE+ub1EEf2XiQ85CvEyBWwUnLFWAvAZ4
AY5D9I1vRcVsPoIg9gJkhEek+eGhkqsIhI+VELRDfSqLhmf6TOA/U9A1GhIiJOgY
m5YtfPHymUBWOzeJ307rsY5L1eFHi6hL1MCMUTlY53UdJ5p5WMu5uTPjrj21nDem
zkqZzcjwmEmBm0qVaOJd8vTFZsc2zE1YA3OWmTJm6jZSAqpL4zSN3BvI2b2ztEuQ
OG7siZtH9PDIohKJcyFkJWpIgtLeHiPgyFr+Ce47Xx9uicH5ZO5Mw30P4YrMpiyv
rdn24W+/bMKsTD3SFR/a4qne05X2rTY3iCWx314DUYpQS8hiAoKkW2/CCOcw+TIB
CY51PWRue8yl6gm8LNcfr6W+GZWLouxnvQaIu2PjMsLnrfnXAN/ryi3ZI4iNalAO
mGefYEinsPk0p4QJzBOvhPA3UTL+ICmn6REliWQ+Q4Jlv8FJMnOTWjzS3Szqgfo7
kehWCCLdZOx2N5nJVwLjiWk0GjTgcLYeh0Zc8encVeyujlhHSy9U/7kTuSdBZzMB
sdTXRfWzMl5BjrkFvV+j2ZkMRAMKEMeX/YjvO42r1CSIyeU3R2nj23P+O/P6eV1/
RA2miy248QUdoWRqN+MgFHNZ6lBJETB1V8x3NpEAgr/G7O+nGim5X1j49n9Ejbqn
ad6agDu/8EEABGurLruFf3GSImol7rj2MJgJC0M+NmqLL88B9HuM+Jf10PzV+jNZ
zHm7/GRfaM/Zyp6rio95HYA3Q5/Kd5NQ9kUOZusBE6KpOvY7fvk7spbhJlLU6/vo
hDKAyJYtvG4T1SdP55zE57NttIRfZenYJRlILbaGWaOnNj4HJc6sVdlbOerPdwjF
zxCaiOYDhgkfA5kfwlq6n3l7wjHUsmKi+S0+2VNFjm+hg34P/C+zjP9eWD+NPle2
VH5/ZEjn63K6r+TR6pQoj1U7+1KHctV2xx/ADd6lOgnd+AI4AQfLJDzh3Jw/vBfk
zR7Gca8RY8DJGBk5hscS5ovo2k+vVBFD/+61gBjlkLCGJHvZzXHKRlm1yFRjtekI
GdUxfe63k/0yWy0FEUvedEaOHf1w8UY9wBgv/5m9zgbfvn+4v3Xy1NvLwwaHx9kM
3VRoUwlHNaLLEaW+NTr4ujZv2W4T4d6K3Z1oE2hmEA2kp3kTKEXyKReyySex1h/u
yAG4VZmzgvagq+IAaV6qvQlQsal8/EA3peyVqtV7J+zUhfgACOr2Bhd4cTdUoxZU
+HJL2ETJuIslxSF2EjG4Lu9vZEHdvdBKPZD47NOkSJ8prrY0hxLe4u8QABikGhJE
Mg2XFoCIdbe8kwCTne8gUOqVuub8Yi8L2xJCPNvkoAkZYFVtAkJz0hKanR4aK2gH
GgR6mC41vNFJCK8TopqKhnbQksysXZGPkb9q+fB2v0ZGmt5DKswEp03MpyU8pfcb
YYnhlz9SZyIULP1gCsep1CGKFu6mcOxkb8Ktup4qPKFa3XzhDI36Ldchm7ahp8uh
uRUanM9SNDcOzj23iGK4CYP4RqhENCsV4qZbFOsX3Wspfb2INS5M9ahCVerBYC2Q
2kGl6Nb58Cs41LwOaCgkK0ZGsPiDcala4phvK1uuZZg2iqH0yjCTsyVRmhG8mcUY
fL2T+phbj9uCfBIqofhCUdvCSH3uCFAiOcgDeUsdiBFM/pBL6wIC6uNnSnMdu6Hf
mnWSw/45JKKc9e9FFYFbiajAUZ7PcYzGX449hHPk0tn245ezUHuglsJuJwe3Iotr
TCF9B88MAKhHZ5QxuCILnsut0b0PuFwi80h3VBYkADYoXMsSe5F+h8shZFFjG1IM
W232z7eo2g6Uejw+SZGQb1pSVEv2oFo9Zt8v0xKTfzGkWe3G+aMyIZZT3NRNfapA
Ksi+uKhASurxWLb6GjQAHvIWtoQ/eeCCJM+fpxeMp7IEDP28tP2KsfPDuKOUf6XH
iU3s4LW3aiisho/EIZjjZCZR23+ofIG1x6unfByneBufxG8QD5yzb318yWyaZpWz
4A+/phaaK1P1mf87hmq/icZUDrR850z+JuVl8cJHm6HoGq8v6TrRHdqiKGL2U7Aq
8grvNNo2q7wYZu/x8i6oZr1hAHHrjFEMJ1HxTtmn6zjmX3HCzfSIQVyxkywNqwrV
jh/EQBgdvYVvwrleQEBLTgz/vYrEae7EkE+jca4j29EDeKLfearrMHGB3+Z2uj9u
ZkoxbwMWqEMye5722Uud5FcoU3mavTScCELXlFsYpfhLzxgek8zR7vmWzkGbANT2
9w/t1Zh4F1sU4R9gb9w+K724aJn7U1yuFdHgPWinDwP0DaehMjHl1F+apxpngX0c
qlIAPCCsi2/CURrrgbv8iE389cHHb372qTiPb9NuACINHunjN/dx5b/Sb1zJ2uMa
mkzuQL0OPvOhKQaTJ7cXp0A+Oyl4Po8PzpkEp35lvtPLo/nSpzjtyIAnt/S7PWh8
mI720rGIyQk8UAfdgLegDJ6vMnM2+dOlyeRTMDFaDmMdmZX103yPNSipAcQeQD5c
uH+uX/KGnpHAqveN0CV5We0uSZYrbd110pGODH/1mgL2D+0DmNsOgwqhD1Fv8dX8
CFTz0i5n9JyoJyzxZ3Xc7NpAQsGjm7+nelBgX4F+pcY0h1HUbgA3Xrissd41UOhM
1OvHDMwMFOelI3g/j5Qti1QCTgD85HGn3MqnwvDKAQthvOUQw/CC/6N8NNeXDZF0
fLrtheJCMn0FYXpU8hRE/hxFfDUwDGpoLU5+fK8r9ogrFbVj+gTTXYs24kf8sbU1
mA0P4ffExsYwtHCfXonfJaUoNjXqu3lhW/h+X5XFEOvLeO+SMw4cU3el1AfIR0vP
sDxuO/WzrTUS09Ahg98bqU4Z0q2vLk85yBuZwdZr4A+9o+2CotAlyuitc7ehxeNP
HE4nFmV6S6C3/Qo9YPgQKECaiQ/PEZp8iGi558kTTh76N0OVwJXqVnZhRcngX36O
34039aM63A3mq0zzj/etgjurgyWn0Zqoodv5HmNlCSgyWlSIxxczocaKqoBgl7xX
FqLyWr2l3eP95l9kMC3k79WidiBKCauzou+YNdnJ7iwhN/rL57p04bBLK3wM8wJE
a7IC/ovO9VaTVKHrHhFDoyegL8k21gaM70RXIoRIbbVIFKNDi9bkla1gXDrE3Lv+
psQE+NM6irxHAqWuoHCGWcNScQ+u26Kkd0YgPCwxciTkPJUnVY73kYbupsk2gsMg
D1aSl0Bz9V2Ux94yn/zOnZMnZt3kw5OI3LSHLl2KQo1z3zOxGT4+Zt3x8q+i8Rpv
ZsoBbxSuuge8dizpICcI/pnfVd0brUFLEEVdvis8ITKjZSHtONAASKcHgQvBfzgr
a0wfml+60cDggXVMPnZkk+O/6ll3KrPjGF6b9RHYhs3LOLOHtj/iZkkJ0v2713or
tS6IPfxp0cT97yOKjpThU7zXI0Wwpo2oXF4NReKuQDMYusXslNsj5Ums9dOdOgol
gSUxjZR44swrAD3nK2+1RjaZydPRqHnACv5to+Z9GdsrYrQA8H8tva+RcVEOpb3N
jJUnMVKIybZ9iyzgIuqx6Tc0q5Gwpq9DgaiSE25AjvC0Spgfl9vQNkkS2mJOr/bS
1gxkxy9okwcdBO8mDRfIiIqd/6CE0hLqfcwoqVPpR6rxqFZZfWAtHIEfcQ6/hFIb
hwZuoad1rWRekzDRUtcW3OBHbLHrwEqpe76KvCgQitTINDgKuqY7VEV0Kt1ukfpA
6Ss6uBy86GMVi2DqMonIxcrxY1PcrHbgRsQp+LAgqnsj+jSsN2KZed2dfdiR4KjW
1eZX+UowbNfjxM4/IKD3YlkZioilIuSnnAPfiAyBgbYuEuAM9HrqIi8yL4ZrSd8F
4akKkyCE3gzHGMcaQVbRmhv33ZKaAwOLr8QZpcMc2GYJQFTbo7roMXRRXlBEz4ta
Izu1GFY1h99iBXZ4Dsvslbd+NmucXya7KRZTC3y0n2ykc2waZjnq6ke3OYx0Qfnt
Fan/wV0Va3QM7sa7aCjqU9936IR2KN11P1iizTYTBqkH3NVAdO0xtPAsZ4XdmWkJ
LFNEfDJUJkTXE3fj54e1/KumIEZRuRgDhElrJGmdzrIVCe5k0dYL0VUttT9ElHHs
yLtz+xe7+Gpbj8t/jU1CG8Luw6GTTNBz+hLd4FzhI3GpUWZRdWj1nKY3quisJyEK
BMYOQIDkff3P8nnjn2KbZagUsLxv7b3ksFgom3SQjDdB5Ofb1i5yDPcKkspPbv7Z
b8S7pZhNq5BegcCDWzn12arm1WTbtgzqkGE0gpd/Je47uWIOvcQ6xu7DzQN9zaIO
ljxfZK/VsMKO0k83oSrfcBFgRJALhCgnn297Fb/4Squ5wyNiQ/65DgqdhiYwotFX
GcyFmlLKq2F9zkuffVKPIF9f1ejFkxhZK6024uj2EjhD1ONQ6V0vrTZibaCXt9oh
H0k41KqyyJzvEAeenfZBT4ZcI//nPAoH2S63JByzgiXRBCvs0RRXl0vtHG5Pkp/w
YtyOTw3ETzMK6yqddjCRNnKjX6SaL35ESSo5ww/q7etFVRQyKFarvWbq51TYK62C
z4h02xtt4lxTxZMSKtQkLiqRGpu6oA8smyxosRIXKcXxZszfTaWpDuHaLqWsiqm7
QolSYilioBHvwfyzDlhY/+uuIw1+Jd1t52lnTUc6B0r3TWFRlP3l5ETrHwFrtpdK
GqYsbQjYduDNfiA93XxG4O3xxW7M9OhGUt3rUbT5OknsvtKRdxMft9niDtxuCaiI
NpYQiY4F9wrRTph8TNY6ixYnPl1WJ9zRj4uCs/pSVNKFKubq5QKHGeoFpSgee++H
9Ca462/9GYzJJyvH9MH8te9sG5KqG+PY07sCIs15ejBTS8CH8jEaRBNqySJoV5/D
2lhlfIjgL03bKlylNY/XNDYF3v+4tPH6OWs64eZ9V9qlSqmArJ7IxfRR90J84Bfy
KTlWh00+euuuNNy/d0j2zg==
`protect end_protected