`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
gMcHP74wBZczB0bB0IzoP2xg5wC5NPjD/GsvSQ6VQgzYAsanETMwwsWi4yhFtJwv
5kY07u0WerSDf8woJ0stqW5xF501W3JLIS8KMiCOd55RHBOnavjYiaaLeu7oUCmB
TtTS1R4sO325rP2zOn9YwRbyyS5Ljn+PzFZZUmkt5xMca3p5NGqKtZW2dV6Babni
5HlLuF20Au601B75m2nv+ZRoGSrpkNElxoTibONmX8gBflpIVE7BehhHwaKSucEF
pp4QQ5zZAZjEC6aplZepouGVggAulz5AahlX5bf4opOVlB1J7IrgyjENtw6ysQ/q
DzybQ+ipztSXBGhmcCVU3A==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="jAI3OJE9Sh00Sic4PtM/KZ4WjwT98XM8AMZrZsQkxWQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hyw9IrFLPQsjvXplweG8O0lkaSLBN9Ijv4B5VdTRt6ipKJT9Kzsb5LxCKvkQyF9n
sGPOd5i74hRHnkHfYISGkfxGJCa55ieOyFShOsqTKRLxclm4oja9vTIey6yFm1BZ
54IDCG9h3PqfDiTD847UCSMRvFssyycwv+BRHQMQlFs=
`protect rights_digest_method = "sha256"
`protect end_toolblock="BnLuc3jxknmZOyxfJK70E5kp9u9O8IQ8cgkXv26kHA8="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 27696 )
`protect data_block
xABArkLxBOK6xG+7CdOOiGu0zbCbHMrEntFfAZEE/xRFxZaAZl1QLkuFI77OC2KL
XxG/mrHJzO3taVHgwRXNLDdc8ePbxbAiQfzV3NJLBO/OTJ0aBvTNnPgPVinF3K9F
vtTh7WTfQzQA1nIFlDFY/+6f5znsukSSn1+QBcTrHWgSeNKb8MwIgMS3lqH+BzdP
YL7zdbd8FKWu3x+KUi4xNG3kLeVJHWeWAUW6daf217YxTXb/Db7uANplrdg+aqLV
Li/XJiDIxns67XBwH3pnyyazrRPArCxAtyDWKB7HNHuuOfM8VTxnpAqeriMsxpSq
FIAHCwmLxoS6EGR0L0R3FCW1IuMLq3JIba74PXl5sYDRRdytKsY2hApklylNeE+/
fDKi0oyv0vXqX2qbYFSosI031V+3Fmxagsugie/t6cfTJWv4FYX74opdAki/h4GQ
YQlsEWboz2emX6p8toFHhU6h0o6mWzfj9uQEVmXX706f3t9zFnY3FD0BiRzN8aR3
vomwN6GfPXTQrchiA44ghVZvJrY4gyL7JPj9xysO84qr0RdXCbrnEvaMs2+YoWpy
FodW0jpTgSwv1QZqK3L8efGAnHv8CJJFU3XRHyKYp8elrrz8XJHJvYk2VuEr/zPV
iQlHlCQVXNseXBRcattOhESxUfMFhgBwOM+pITDiROR+hFrEe8orIz66BorNWQtO
g4+CuJCf4pz5EMcCEOxq4VZR4CqBJHXBzid2HiiMI8SGeTVxXtCZMaI2Fqo/XZpK
QLwSH6XJJ7I2YYnZmjXnAW8p1ax3+1g0DhpcKGC7IBGdVblFt8nNnsCmfWGpgM1x
0ZDd+8BveBzMaRWGsfg2Mb0FFFxPGKd4Ovlw+dK31UvKIptJ+iKBcGtOtVieU5rm
/7fCLexzCBUu2GEgvyriCyLscsBXn805Eju+iVJ0NsTdfiGWnEaTU3BBzZOLp0Sz
QrkteODcMj0qs4v44i2xKJppt3gY6goh7DNgrH9oafCrZ0mhGGCHvdsND1pxpeL9
FfsWS71f7gZ4cwMygIHgNWH0RF47/vmYCKLmfcNRWnPqKp8YjHnOLNmYtjM3vk/0
vzh3xpFUYSJNebh6AyQUY2yR32+GpOGFLJTLeCH8Uo2fZuEzjbNx+p5NyMkDa69Q
peGXy8UD+ZCMtUfX2XeqRK3nVoPkyMGLlXr75KNfHaaFfAjAYvH/dIA+8lpf+SFO
adptQP3cfdNdQC9m1Rbeq8EkmAY3nhRJcmcSJIWCxnjgRLD7S3d3Aj3eJF06pbjX
2FhxPd0/khMnvfrXDOdDEVlJ5MJr3gwZUfU3l575hrvkeFDDddsHi30OlM1V7URc
r2o8IJDenQFFtcKDCDuUWVBq2rXFj3KW+K4LzaLlST84aQxMsfnSj675NKpI1M7E
Ab+8hrcCieVXf6ImEmFZqEfxRdw3RxGPO2inWt51l2iE/iIm2gypWDZ57ZCxU0zl
OaXbb41b51kdTrxpxm2ibE5kNhKEdbcXgtfdTeVhgwD0f39N4xGDElkQuN7hF2BS
FsOrQP8Hy5oPrAAHXmw+tDir1ecm8UzSzf4TISUfndF8d4bltkafXz3zps89rukA
zhOx4sU9kJ3MMYJVTwLgjIqM9CN3VP5J/KBvN1EF7rSSUeLI5mXHOq0mUkui+IbK
sYqRcOwuHSBUt8iQYQH8c3HJa5+CqiGilQj494jB3R26+VniAhQ//5sgFUMZoFiV
KaGvJNqlw7BJ3mpyxp/qR80PXeTbHj9DnMabP4XBrStRXIv9UpxYwd5/ZAj3iBgM
RD0wbzDHvhr4S7FLZ6xlO6zBj73c4fd1JpFq6YiHyCKVd0FKzIhitCA8VIuA6F0E
TzrK6OuWaWvVC+SMmTHhaqptll0fZ8bYNVLMthl1RsMlGsVi0rlF2bDoQUeRJpVs
KtXgayJMJW9o2giBhBPsz8BVU83uJbkdtSk3nuy9lgKkmzKFrJT1j/XFTS6Y1iRH
ENa/zLBQ2ZqQXyif6r7pX4lZVxUS0pg/KvugHjQk5crJ+kvsdknVg90jdb4P94l1
UpsRlqbSAq2+ZIDX97alp3Pvv6sB8Xloub3lzBwJnbh7ufvVSRssvylFmxk/h1zU
v0E0BO0EWTK/rt/GFwsfGu0vrwvf+NLQTe3LsXFYo3YsHDZk3O0nj7NWiWzCq/02
lbAi28LNfbAag6/6DOrIBJNF8P/+BjFBlUFdAkngMVKvESqhdZOK92BqfemDzdgn
UNMgBW1EHCmqxglSVvYgR1ZbMO+Mb56KiH4SKd75owxSeYSEM/oUU/r1zD8n3fV0
v9XmmtwthgsZC4kenuqsJsnbEeIVvdasToMoPn6dnwhPTQ7l6RHhc8qkHbga9Itn
u7ThEPOKNPGabz/d5gIigXPTr4CTr39BOd4nbchSY49VtyKcmPzFWzEfHaqSXtFK
xSYtX6MaTgvPZyDI/RzTjqTr3VcMA+k5ocb32janOdRbHB55dKZlQYhQwu9tGuTO
IJ+O0agUAIJrnyFKibBLeyuod40AZe5dBCvV8WA1HZLtaCRg/PitGJxFodK4pggm
4f+V+uQd6QjfpT2/3CthaDXtIrpz8r62qqRp56MFAop44ONG9reiNrkl/rnxBQLa
i8yEfIMchWvWRDlj3c63NTZMRoHEWkzVoaoJl46sMiXpo32fopO5DMMWMgpPMx8E
U5ezPeMYAVGa4bkIXEDIq1eOVue9h/J9cyXHPulhXTvws/ZaRkaFmH6CRLpeqoOA
AbcPLk3Fv04jEw6x2H4xmjlVsTfptxEHpfz+GyRFhESL50bZLei59ftcA1R7nv1Z
K/Cb6fCXfySP+5vmJcfTh3MUAY5tN7bZBtkFpSdQK5ltj8MMix11URx6W7zo8WkN
CqsgZhngHee5umlYvM5CI/Ye2d0FZwrbt2RxH4+HiGoYcjqYCPWCkERNIsveMaz2
9AVCWjnYqqILPp4B8nV4nJ+PzPX6m42vKlMcsPBNm/uR7JNlwSscxd6yuuzl7tmZ
agtf3fg0wj2d4MUVb4cbT+NgxZKSkI2sYuTsHmYlimUoUos3jrQ7MB/73EXeuYzA
EZ4ew6QpdCeX2lXo8p6BQT5xJpKp+vg7Nz821WfeNnnYJOnvZQITebJft1lO+9j0
/Ret/+B07AUkhhKiqIwh8PhS7qHCHMnrRMt8+z4GaurCBjRwju5cCB0qMvE90W0c
E7sd8qAJeiDdKHS6iLsub/01mAI85DruByu/gXUrS88bsoHXsHOKC8+h/ZgcNJFS
VQcCVTvSS9N1engedBo4lkWGqN4KBxhVA6H77Nm3kxcAN1AdX+IRg/QadYX6g5vq
h0e8oih0SHVfgkpNcRserJxc8q/AAb8ji/9W2tJdNFRaJ8FvuIM7ianY9G19UY1w
7CwsCU1058l+wCTAF7WeK7zx4No/X7/KE44f0YOxfGw1cokvl2u1ESlNBEaLRCi5
odq6wQyopRriU/T0el6qWevaeL3aYY6BbazTs32XXWICHTgOw0bKaSh2lICUqqHL
9ACvmUxfhp9azShb6skMS+Dw1MMHVgihJHAzPagKT90EF7k1rm6tC3b41cbSiHCQ
jMRhCFYga+QRTl+IxQllWMGAn1TjKR2+yg5fwQ5it9UUZv55Poqf5KpnypZPu4Ht
0+XDg3Ls4kfaX1cmBGh3TgAL4acEPzl5bPZANef6brcScTI5p1RS+PGb4Nsb0PLC
DFZhHsqXS6qLfdjw+52FC4XnDw49zKaVSChdKgHG4+0RlQ/b5JN9gxF3UiTNzbKT
o2B4K2KRiXHBmlRPMiwXjCq/dJW8CTIsvVg/511I48x0H/kY5nkwRVyaX7YVdZe2
PcTroChIotBPpylXu1vFcGtwL7i1BPKY4DN6Z+7yp7KSqgzrwS10SulPwg7SXIrj
w6KYH37WpzhwHn8Z28hCNzqC18Ykn9CmbdCkPvTAj9hyUqCQfaRFyETRVxrf3oGI
wpZegDuJE8cYAzSbw3f2qcjLPF/aUYNm2u4aDnWwdjMyn3mOTzQeZUPvQ+4rPJ4X
Xr0CZRK+GHWL3Di3eB0MxasP2uHIhekgZE5glpDZOkbLA3rwfelfNJWdOzoKNfeK
AVWLShxORUZk+rEf6cVSmcVynjerQh8DbUx4U2LvKCupOY8lS7gAowpak/zqSwL8
37+yVrUlladzj+KvHNqlC9n3yJMXaSDUQ30qYpLNaXycZrNC3j+NU4w13CzGNb2Q
71m+t6DeUjIsFUM9iZlSaBiLiFBuPWZKyjZRQNDczvXKvFfX7kRNDaB3Pwcuw/KH
V/3MMTqru4CnI2Aw8P3FVXZ6bb8GRpf5aG5qjShPRFQHbNVt2p4KOT3auRLeeb0F
7PWV0HBcomOiUmsggtZWqILQr4eZHy3n3l8TkzJ9HnYXu32srN8IM9XUGFO1InQJ
EZ/KhL31b7EB1S5Qis0cKBIKtwOT7BkfPK82FYycmfsPadhjV7s/VuEPQEMNFVJ5
J90Q3Fz+0BbzLc3gUVGACAkuFD9M/ynkh0nb7udXp0ogj+j013xLI+/M2LghvEA3
XV/QQUjC7iO9+eUmWBPwhOoimgfqCGamXMLkeD71oggzvxcweUW2+0AFEg6kJOeZ
ojqp5tWeFCv8uB+oedWPsbzAEy1O3C6YNP6ed3jeoijC3Kv4z7h6RvrWXJh5Oxr6
iTGIPmYjb+5PDDZsjKx8HGLzQIB5Kn3OtyDl/L4bE47hH9Uxew2E+wgFKiFR/y1Y
P+LF/Mq6CBszoFEe5ywjPSFHueAOmbaHF4ir8Zo3DZtwPq+GlAUSUBVzY7sDnxHF
6xcTuiFlUjvuJb9MI98v4ePpie0+asmnGdnudBlIqh2OMaKyHQGEUAJI8jy0UQPx
vBf4XcnjDmzAkLu51V8mcbDp7mR6NXOcItFpB5pZfe3yLJXgGswR2EV5WsRmxm9T
8ZlLZVrRHjav8/9f81OhMCMwaVRLfbIQ1Dxxr3YukgF4sIsUyATrzpmvLEc+F+QZ
VX/TFHv5K2P101QUwRmCHo20JGaiG6EUvtojvv3qfpSagEMy3ll04oFjQowrk0g6
OZ7Q/bHL2Favn60xKnUHjdVgACGSQ586nUD8U2rtN4LfBS0ck0Sc2aNWjtVsTsV2
M7sGbXRaHGQ0A120vh0/N8TIzJWjstMB6DI1RtqvXytJOOle/iVa42iwvNyWaf/S
b7JvBt5rSw12ZD2/89IUoG3PBqckkZdUlgGKLA6Q7wlyNhtPrjTFBpiH+ad6o1dw
lQzrfJl4s7Resqjt092gmRZMwmf45HNadPngIzwSYDxyRId4r9TFH0MsJ+2jFNax
G4PkoPDZT2FhS9ELy4YRJCqQYChYi3Kd0DyBFReQUGfjncBu4btFTA/gOm/GuUK9
ga7ylD9TZUTJl+I4YUTLtDwh2LuhEn4dXeTM8hLebrCZCLirE5mf21vVoXsb0NSM
xix7Y4uNYaEWA64ptnzioqfnI1S0C4tRky+3raRA9YlxyGHEJeylUgXdmuaM1EUH
S12BzYxFhgz+9z5116vL/h/Z9Op95FkDtgFADYbx0pSZp8GCN6ZDyWbfRzSkWvN/
dimJkrM8chsp2UQth/aRmm1Trc4HnS6qH5fMi+7Es6xe8dkhjWHjYpgAk6cDHIhh
7i1KlBkmiRoVwhxPzq0hR6eKb6BMuv274x0IwH2rdiAQQYKEp1oJo2bUppn05tnA
+MsBFawzyk6ipMth1wAKjDYA+4LaHL2G5aDAjG1TMN5aqEnPGCmF0yWiN2u6JS2G
nHEKbDvD7md78++swpwKyfaIaZQ0DMaqPHLi1KIwE87xyGLvboKPzoAGgnnhNctn
rdpr68BEmEzXv4uG5Q036V6n/aeQUsvomxSU0DbzM2kDUSbzcC4CctzjZCCp7nJQ
RmWVjM/vuTzECwk9JzSWwHLZjkilXnULhIr+NeNst/gxLafpy34HYWh6hfJBfYSQ
Wxuefd2MGECeo43d+XRMzCwFYiu9RnFM5In4wjall+gmd09KuHUNPOA9DNEoXXgI
1xCRBzqD+YNb+wDMvzlLfj3/kXdYl2YhopQumOCTvs6qRSLDhO4qnebDoEnnO9Yg
s7SWK5i7mcjz5Jji5oY1WReWAfRC7M2C2jMk8xhmLsn3elbDva8Ai/r8VLEq1RtR
m/cBjLKbtNTozi3ywqsxALRVT61ySRre0cYRrnW57WO8opZb5yUq3If8HkoYdx5P
cnraFMsyYc+ron0wqBLmYPe96h8K54CDT6W2lyg7pw+XDPLaczxo9uObqOE6zzbH
Ub5TMNj92VhWiMaUYxz6x6I2xjBVjpYi946M5Rt7SZhnokRGk9cS1wuKLH45xLyV
H+jRDpHzjRGQcRS5/HudiCvP2yyD0kY66h7DVHy7zQZqJ0g7v7/P4KzDPkS15lV/
xEsC83qcdRmnFlKTczWzZFGDNASTPf9I9oZneihGTszaEraYBZmGCuqX6ZG0qwMA
rizBzZkYB1xAXtBbtD+ZGf5LmmYk6jP74+S0LIasplu2lZdwsAcbO7p4BV7yHqat
XHF1MVjRftlc5vQ4YGO7q4HcpH2yE976EnCqaiUaU1nqgHdfCgDMzsDJ+CWzo797
Ox7jZzBrdSEo8yL0wu9RpvmTH6U8X5XgIO5swqRY8zrPpVCLjpXtmMKgxoUepvbB
XpPNLNDSu7Q8k4f5fMbFPU6n3u1q0b1wlQyB4669WPimI8uATQJIErzk8b1SoiDS
kSlnBw+hx4KtyI5gDS9qVkxw+G3mjK0PZy/h1vD6IeJmC0cuXcO/4qpPTK0TlVpf
cmuHE+ykAkDhIbWKQ/93TpYj0rUkfyewWNTttb3iXufOB93hL68RTvzjY0KRnOMY
9BDyyf5A6A0xc+k1UoICtbz6lznbZ8BcD93pvPkEOZbV0ccgsTjAkf4jiG0Z2Z4n
+KxQ9rMrYJKejS5xJ7081Jv6Kq0otnuq7PNaHlNbvlqiH5guqUdTZtgnCVQKA8Uu
j0q7daNXYOTPK8yNxqyDfiM62mzTsYUwSvHKf6BZew08wcxljPXvuRWGi/3DdzdK
vux93idgdo6uCXM2/Kvkwv9HbzLuIa8T6aFnHE+PQOrquEdJg1mZWsaQ7YltXzyo
/hirShZQ5oTTrJTdMUbXA29C7q74WFaQTWwvGRlfifCauplf3zrDMozUWjaIneSz
BFvs2pQjG8216HW9fNxxwmMMyPlgMSeBYll1wn4JvgxBs1xYlJ5IPMWQowCW3Lp5
DnVssz+hQKvbZPlFZ9kuKz1JzJL+bMu6ONYqpmzwdwG9fmV4uQWnERIj6G/ahivn
Ji7Jz6npcraWvxys/7cyECyvDAfg0qp+/fp6O458BmN39iTUdpl1X4OfdEGyAV0Z
MZMfr9Op55KgYS4ncq0Rd41cwf0TZhI+jzwMkHTtYM9sh58ammCSC9ilIQBmS9pu
gVISdC5AuNvOeZ6izm5k+FEzgVW/mZ/dgTRcqzel3EG6L5a88O5LvhKhvn5Nl11a
LZxXvg/8OY1EZdrdpjMs5/reDNlhVuCOVnlQOxmzWnJAq6lur7IirSt3KYBvXB8w
7/ri8FDthiK2iPE6+ItsBMPYD85rI+j1WDADImeUpeGEES+a/EFF4AqNgcVwETs0
7oj1NgJHXYGoW1ihJhRhqhQQx6wO2b5iAhLH6qVh58dVGdpyeuOLZTxbifsRkxtI
R9LZb1PYGxjHUJFzJU62MOxg/jq5aFz7CVgsiVxO+upFP4WFKMMMpyPbm7N4XfYH
I46KQaQpKpIJNWg1kxcH6XhFnUdUXwV6AxPuz0scWQ/B/IiRA4Ht4ueWzRwZ3OMR
ypHbq0I2M6fFcCjkEHNupq8Py3BDUMHj/LqxFn8Bx7FIPC3SblQPk9umOHfEGRAb
xM9P4Prv+d2wxZgJWpkSLc8FMPVnrSInT/sPS0bNQn8IIDkaj9FcotZEmxwq0K7L
J5d2skpWB9yruDiX4qCE49n41O7K+D+CWvAzZdBF3zURl7pRGQ9auZ/nSHV4lK2M
FDbi2YPFpnYg5fRPoozT5vcAeDuviCFmaKz7TbGVpf3ukHfx83rFwpVnBADUweSC
yc4TasDtXXBwYDpxPuuKpFCrCwfkgNSGVd2YGlLhPGkoc8ChIpJKi6NEL62gbB4K
dyshnlwB4yU45bwdTchW99gyRpjS9Byw7/8TWWzJhF7t02J2np7IDB8IbuhXiR0t
sXjlFF87lcvGQtWmgwdpcBAy5t9jzPhLaiIcq3HogMqKLfU02RSVaEL7QSJPuSrv
mtUfTiQf2tJQbyNNDaYQx0FyV0ROKApCx/qve0a6/ya/556Ub7wdfU+tBTHig6mI
MJYn410/D9LwR1NnZfvNwkK+DyDUmn25s9VmByMajyciS8++va0QSWNmV+BH8N5P
FPkZULB6S/Xwln3JsV28XGAxA1RkRrdnmMc8RBR93VFwUrtLqdk/aa4nlsPOg4sn
uEBZVdLfGIR57t/YuSw5SNf5TEtFgDH7x7LN5L3oITCfvBaLeEePKtiTqABeDzLU
tWzTBQBq9SbuupLDTMjywt4SvYsIbWoQd/rkoleBT3B2Du4BzbQo2Tki0SqKGb7B
Ili+wV7lyqWxDgMboO9uCZTJWD51dJiVgBrf8vLg0ko1q6WToZV7cieCvPUevwVS
bn6bbUoKrtAHeAYNbmSYuwGXh6AoWXBtNodUQrbLXtZ8cLP+6NZ2qL8kZzLh3QBU
x9Fti1rcbUtdVU/SIqgMg62ahHsaM0RXAJFOxQc6i6YIK7ClRSWO/8HKT0FmJjRA
739xnE4Fa7Bn03jT9Z6tIAFDczqsBM3iZHMdpIIglnF+XPd3P1fuFbsdKLOsHMnn
UyXR+xFCuN0ZFYiQ8pPq14hGdnVXG4jy1QVm0ggHjBo1lOJX5c2cDxslypmISM6y
0gouIRhlehUZqFLi6JPKgEsnfYZbT8ZlYEv9PK/OK1VAwttXMR9vTrjGbI9hGusm
agNGRcsBUmGp2AZTr550yMbREGCVw5ozodgzOXZcS2OPgFcO3uSyaq7KUlQxVRLI
Gbr7ABWtbd2NiklQNttuPauOtn+sz/WtasYuvE+nR5QQuiz6DYAl00aB/Oj3Ksnj
aclFn5WXSQRVBsRhKTRNxoNtSzGsFBlB+/yLRF2BvJ+hEh2vQhKlACXQPJPNUi1G
6EyuubB8fzpai/Y7pLxvi7zjoJ2L+U8OJ+Anmp9coWIzM6+teLKysA6U55KYPgeD
TqMRKDM7vqBPXMpxvvJmFoVcUfsDbqvIIhN3kmhgyX923zBBiCVmudCw/T08WmK8
4GOZtivRqWS9lmc26QIt96Id7vXPlY6Nd6SRQJbpN1pVhOXHsTAmp96AGQB2yF2n
s1AdacavInGS9xArPlajHtzgjbiFPpXTWnT+46/5rJt9iW6414Brod/+CU+UnVH7
pQY4cFawKrOlG7aHwSVXBS6oZt4gDdnrqr3bWVrqtnT7GomGGaiSz4ajdfRIzEwS
ObT/OV1jTVrGgIwR2q7V0Xzkbt6sTeT36PBojPainUluYA10IGxs7Bs/gV3I0Tjo
jqzvkSoZvuBhoGyIV57Q0zxVSA6dlqgsM2CmJeFUwJcgJUxoS2MNbHfLV+DsMuZH
c+42nQuAmXvCNbDLrhH5pGyaq0FFC9OAJf4XjjFr3D9wvtzEHcyVWNabfIzAr0Xk
DdzczHUBWgjh+/sRpHjHyl8MqWXEqGtsROkyXHnMuWqPgRmeXowa6HIEYgZsZCZu
drJzB06rEoHI3x96Y95rbd+mPDZJlsyAPs19SP9YBXAm8xgg3RFsC3Zf/H6DLTz1
dEukj5iUxyzTO6czEN67tcSdE6GmJLleGe5h4DJkTQO7nPSwstXzMX5UkWjuHbYc
Hpp7n0fEvDF2ZGN1TCrGqbN4g0F3U3FFyErLIF7NW/VTks95vObAW6YSJfE6d+97
VXjcimqyZYs6IOrmTQ23i9RoQjUa39iMQklHGa84jiWhSwqLOTRhH8OIX2ztzdTd
UP8YgKZWnG6ArveX9VUzpHEeeiMs/sc7ShYzfCn8WJBs4UenZmUe0q/WvsnFHgVz
dFxFqgOj9dkWf4gpkkXsC1g3xZNS/jfyNfp/GzUicgnbozBMouuN/2dn+dtPHzrm
ur6kdfsDsNCj25KyDWbCtHz+Q2hAWGMtZNHqLiC4kJ2gAtBUfV7+FYWYyS+0UeXS
0/37MlgETKu23NIMvhJcKgevC4AQjC9S9TA7Oi5XmQ6a8e4CJm1JuZ9KCuy7Zo8F
9UjHCTUkmGyBmN7S+Ats3yLSG9WKm4rWPM88U462ukVqTyP0WyZH4EqOnf8JsnHu
oFK/ycGQNdGVloFH5uwltR/NcRb7yzJ/kDpdqY+oGwhA6cZEp8DGc6brnE7p6Civ
GWd5gJOy1gUkqI+aSX1U+fCLoZz3ZY7+RKEjcI8WRxSGLcRxMq2zUIW650djR1oy
uwXLs0lBkKG29QlEWgKzuM50oJpC+XMWPkN1H/OAIVS5AWaYyJeVxky3ito9FXGH
Jt9knsspOmDSr+bWSX62vw5Rk3yqLP75wfEGgVld7iF2osNcfmAPLm0h0Zh3tVIF
U11LM8wE6lr2RrI3Wk3fKuYkOnXHbwqog/02BKwhkDOlh9YuAQy6OhFDEqtjmn8K
ag0nhN+LXrWL7yzrLYIdFTb/4f/iPGtITRjavXlnrCkVMCU9/h59/Ttsde73oywm
CEdpV3V+x1lJ176n7aSNcLtxhy+q4QLks/Mdmq16q3E704bfVBCQCcp+wQ201BIv
05coM/dgPIHj4Xtm9bZerMjx5acrIT8WBEb0DD+Wz+JO2BF9PZrcZln5iDfldP6H
BJ7gG8Qh5I06ceRfFm0eIGZcChS/JFeED048vmCMNGH7iGzmEW0/JfG2F7foTbSD
FIuhKacsO3RBW5UNTzizDZ+8V50WDoPh5CQ45zw7J5PZ1f/GWXvqUjtNOoViim7b
uAN1iA3DoV5gksCEeaU3Z/6FVyclQnklpo3Etu1ONUQ//tmwvGC5cNlg4RQBknxn
pP643AJK6max088Q2xHO8OL5or5cV7OVs84n0EqDrDP4bxP723tP0cZeg+eKUjDO
kC9RA+JULBp69H9jjE9W0qoCIxKy/6LrPhQKRDMgXYG7YFM5dv5jWW7df50jpggv
rApFyKLVfvesvK0f4b4XiXGKYFdyjCC8+dd2CTNR1hXe/wzIPbjhEpeQYNlo+yvU
D4iHW93trDB//+iDpGn+Dl6g3+pKBWvfc22mEy9gRBf1sFKWs5QiIDGDfQGHbd9n
O92YGh0xxY+NeVg/tb2oi6wA6ng1N9mJXZDm7Yv7zK9HwNNOALcd0RqcA6qxNBSZ
no0zF+p7NR1QIovWfwS8y4gVDYKF+eed/bHuE96kxX13eq3N7kQ4J/y9OnafHF4T
VxC/KzsT1ondOj2VWs/Fd1RM4uS/xdBQQSdGU0YmiQxAZTmZMjvAeeK0twNCl4u0
GWQKBMTJXe2lHltTqa7so3WbmjThTtA68DYfTK1d7+FEYaxP1UVwjOh8RSgSHFp9
6b4m3AFdCDLxR3aoHX4FHCcCVTKnUg6xrK/NFDhzsBRIwj0g+aLvP46AcSeEulr0
8YKT3YXBsUGACmN73LkoHsu8p4k+5dWTYbg9HxjnMZlK5z9iFXTQV+nvr9FbmMB4
ldVcmZdhH96WfS7Fv1wm+WcYoIbfoSDJQgIrSr1GEGdRMVVXngeCFXq3/pqq5a+Z
PdPHfR75F2BKhnVJnwo+jMsHPYJYYt1RCZY6UewxDjlP670it8cOqzA9MEApY4Vr
THsMgv4ytXG1xvdc8JSREdL0w4ZIOfbyMUlb2pw3HoFIOdyqtdIPu5JucilRDJNt
sdA/ManSBlWfuhhD83aivxeI3Nn1KaucvDG44qB1n5tjN4eK2m+UmQjQLPXXC6yc
iDIRkX6v5N0Wennb7QZ4ib/+yCzIsmqFH2iQ5dtuYS4xlSoQVuQgfm0p2Efd2JAS
Tc6TRjur6v7H9N1sBezJNfRrv9/UxPd1v6c8POE3e0xqn3AfxMy8xuhGiF0rCEE8
J/gUxCkibXHUlhqLBoN+vvYerNcjuSlrMj0aSJosF/BVn9yUwLza2aSo11OPp8L+
+zc1sbZ44cBd1p6AGdLEWNhETf/2hhfcQQhzV3dqdSBIpWjQHnQ/FT2Bu76dtSL0
/NwVLZE6IVjio7v6DLBuY3/N6EOAWik3/5/DZxWrqn1V1KWW4b75jHt8nC8IWzsA
yKvyj9Ebod+7hs8ITcEeBFflPQhAHQwKI01PSTVtw3AUAK9g+UFlJt4w+35msvyT
JQeEJpbHSFmvUTRXa8laOD+l7j5llMeDzCtYucHrk0QqNDEZ5szQBT8D61rbNa2j
11GHOlTs8edmmgWRCxhNO83GykqLF4FIdTqrDWkQTpG4D2hHYLVqdlHKDcy48Nww
h/J3brpPzEFqWU4jsPrFHiflohWqL+8YpRguGOPqEc5kckqsw6VVjNdhZWtkoP1H
qa6RsM5Dw9cEfClQnczVPBrcEmu5+HHuj2xjApfzTu71v2GRHCGIJz1l2lkFUbJX
MdoYfElBS/VQBv73xF+hKnFpwIRB7w7hE9pPLkhC6JTKHBOaTgl373T9QNYiS4Ko
58U4Z3Lhjledp3iGlhhtK3ZcGj97oamqZZLpcxUBsi/PA9ZRyoS6AhexQ86JUhqz
bsja1bMZw0+Rom4y1haGJjoW+9oVKcRjqE9u+/Z3qQQV71uPJu4QEq7sIZ9aejW2
xHNPTVDAUjO8Ywa5XUodYTr3bWPYx/cBnmrljciPB1D76ruoA6/BLpeZJE8xPgx9
p8UcS8slxXcXacBl7G0PDDllu8ihycxavWe3BO/yrcUQIvx6HYV4UVzm1wWBmrSh
0niPJmFCoWvfC9A+u/w8b/7IxnfMUAYVgLrjTsHreE7VeoGl9keV/PtnI55Jk9tL
esSen5pWBwuissKvZL2fIXbfkMXQdUZ2q69Wq9VP2Al/d+lZExu1gD6mirLSFMh6
xvvhZoTcF1sOg4qE39Xd3znaH0HdqvVe1Z4DqSBVks+FzaK4t5RKJ9/vdCloazOa
/pqlhDdaaRQm1+h7HZq0bBDmeZR0snzYN1hCydfL1jJikrEWElNdVx59iMQYHMC5
t9gQTommNiPYspG1NXxUSa4IvFXeyyirz1oIMj9xgntTwUkMtWqHCsJtCMlgJ5IN
TTZSYul+kcN2PT8YHbUUNO3T4KwnQeblXpwWZng2DXa8vAUq1oiWo4RBL52g2/lz
BPdZiil1x+4x4JyAzKHcOE2WvOOMnY0CqCmSexNcVThBfaex63qK5kz3W1zyowBo
xmvrrDw8nlizLnk43ep+M6VP4AFFvfwUsxgyojk9snkKvr6amcUKDiaXiS++osG0
0miBrfzSC+QQzdyZm1tui7wNYkXfwG63P9F0oZOrfkmiqp/LF6m+iYc/Xo4xzlwe
dg9R2/MYARRNKiDni7KCbVmV/JMc5y80UNWzfbnfjKnCbLZMEbPWjbpaNXoV/GNa
qwACvawrAVxixU9PFiyb0s8/R3R8pgPbDGtYAyjZHKq3Os8+xkjXFCdoxZy7hK1p
uNWkwKlSay6zEuPM8fw3bANgQFHDVt9Gjod1ucXkg6NREmMzKGz+/PDo4bZ2qP9S
AKZWCyW5mx3MX2TOxdCJ0yyc3DySDYeZCya4Soauzz0ynzdfGYqtEKwlc0Sr9tDM
Db51dDJTYetnVlKRALCu1o+O6sm3Cs7gdequpk3jB72T1bJK3tErJiz6jeOX+tgK
IxfCoTvE/hqYte7U4IfMg9EKwt6oakIWn8hDihPSNkXu32Mq+KDLoXRI4w8AYlyH
GWHMTD3jCZYgMRYgxzhqJK2iqdqUOp9ij6bojqFG9I81CAMj3cu3dXbRf7cN8rmj
oeuHmqyjQ2ppnvgtUIS5nYdXqhtsVwLeujygZ8tey6ZzSYWE1Ppzj5q1u85KcadE
98ghvUxX/fzNhkjdUrgNLcF1rpx/Ts0XVu3jjD7zBCmGIuBpncoqIMQj71f1lNii
aMebB2DGWLadrHjuDJAqZWdKhl7uwplkSkAF8MksETIr/RxPAi2g6j2QCyjgEadJ
3ZWr1SWEV6bE8pqRONPX/rZNwl61eiJGCvLBVXjgaJ044m4fJqQ8hIDsKPv/+DXG
eLw6MEAsu7+/VfmWPAQj0A4pKCzPsyLgkOW04G2oLDo/oeSihIW8Hc7jeCCG0dD/
ujc0u4L21TJZl/rjN1iIDpafDicjV8TPizwObJWqMai13qEyCeQgHGWFuIZTcSw5
dpNhzgjgWi0brK1vg5ADoGHENKd6CrMtGJnxq3VyoA8QhhEyJ+wPOPqgJdn3VPJj
H35bZ7ZknrgnldcacGQf1pTKuWB2ptxDwYb0r19cdUJqRj5GEiNif7NFBoq52mXd
M2c44SmsxTQdDz/OCaVHH4CgQBXwwBsG3bXJABfErTwfrd8/Vf/nPYYhkFScHXHu
L75WkCY6Z0k+TGnye47u2Sg7kcBYI49UZ84uQY1zgLIJfTu9d6+wmtyd6zJmk/CJ
6ECxvXVR61qXW1fSj2dYIdqT2A+uMgsfqfNLcG8pPFf+hIPr1W/EtSHaPV6XIYHN
K8qlnILp7K6azWemJmKB2/tU8NBMnkwvmtcThY2AG7pN7LfnpH0uBA9uaxTf2Cps
8XhvCpchk9c0WkX5Yp1Z3JUwjYJClW4iPKaua3cafvfVJkVb7GgzXlW5Ox2WvI08
mU09KDnMt8JSp0YsIks1iXyrpXXvRdV8vVerIkt4p3LX4v+JktHl/3I5khCuLhXK
48799mvNhzAbqHshBs+u9GZkQUZc2ep5plqoYzUzWZU8AWCkay4HSCdNmhS/0NEn
6LcCXjV1vpgG9lvFewGqTznNnFqVrWnfznW/508P4JQwbd/U7sKxHhBxUaAYDew4
AuGzwXUAVfJukR3tdU1Ef04YrAqULV7C3XjvwMMZ66dFc8++euUaH0rIUNVUhgUM
0o4c9GkfWIPgOW3/mfQabIVCVOr0ND1J0bOjI7HzieD0N+qmK06egnpy5ttPi2r6
ww/cZ+y1EqLAGR3dLXLRgr5Gm+i2ncAQfrSQNa/rblLpe06nogELPrvYYYrPtNUE
l4rvx+o3wbV30ZWmbJJJSdoyW1EwY2kEGFDHx9fmjXu5E5/P/EUmKMj8sir+1wou
0HwxAklyfueE+VEidhvs6d7qFwiplXT7YlrAFrfmCSewrOPHh0r/6bYoFVUW/UkO
hnpKbHpoDXpboM/vjx+5/WH6h4MmX49BEgoFIiglsHfSgRaD2kd3CxT2i0xp2pDz
TGqdvptOmZKixOaI5IS7V7JFlwU8SdL370F0TolkdLGHgFdcFz20pTx0M3ktmXAO
Uc8pyZYRGOtfaMJbdKDX67ZcKFmTCrkHzVRkw+zTafcDFHIm9AI9i1tBL3l7m+Xl
EjrdXSJDeYQrOKvuIS4e1ntwBZ2SZzEmRFhIg98zLkOdkUW09B/MNe6oBJT5jzfd
uw6VRs/W+zZHkJs3TpLxsCe2yo/9mlnO2T4GV3WpMFhWThY84/Z2H5F/Zp+gEL3P
X5g4kXXsG0R1PeTcSSp36sqoRTz3tqUCWtfb/xRFfR32ZL4sa0B30LVrrM48I31e
QV8ige9uZbujawajxnvHK0c9sJKviDXPD4/IhkaShgz1K7sMuT5ZdcTYxj6BN2W2
kMnaCAQj4ziDMl5Ht2/4RphZLZVK0aFk1g9TJM8gzoFHZJKbTmFHLkMtgoM0hoNP
aIunJ+sk/+RWfzVQhp4N8V4uqp9d7gLKXH3e1WmF6nC+bhRLutN4/RnN/LKXRJRf
5eEJ35Eavk44jHgl28p9UeB9kecoNuHpY/suJVYyWhHETTvvjFewrc/+dl0GavsS
RpayklNkK50rX0kW5Q78FrkdZrZMg3ZCu/Xw0tyixkCh+FI+w28lI+abPceRBt7Y
js9VDeZoPFN+xpqA43yl926ZvB2kx9sm2eMMDueqy3zYBvIamOrM2zVXdM4aLVw6
gMReQ/YNp/H5IyLA2mgeL/Zw8LBp+Oowaq0QCKH+pPxTaiJgvwuNL8lkDXF3C4/g
CHrcwn6EnqC6/pyFp40EmyzVUrhs8/9UGe87bRcN1sbtWx4PN7yECFzfwuxKcoAW
MmDMQRblvG0vMDioQMjsjsuuQxhWSVVlrSOzeRe5UeioBySDPo0NeCK2tNtDCUaV
S1OAOVya89DznxcojoPWpXbXyi5vT3EWkALy/kLIO5JYOl2U7HoCqGGLcgkAuGxy
i1hazuBaMcqOvZabDwxcJB4H9jN3xBlGujGAtG6628/+0jUQOktO5WmRNMeO2IH1
6rFhJO8KnhykTKc5tlTOz25hBpafy85Lm5cJ/IVHAh6R9TT2vrdnomwsfRneUYIA
37TOqx2MMFchst6YiUm+2pBKgowOxzubBuMKmVlNBMHt2s4ml6CBKkW54zKK9eZX
gpN2nzTH0l5a7YTsK+dl+sUpJlWNGty3/ehDxw7yEvd+P+Ud6mEzb8qVhIZwO8fg
oPCFOHQU1kz90pEv84RogbDwC7sJxrrPSZ+d9RDucbsZzskZ7ABFWJyHM4bK2uf8
KwL8rd4OKeqaCbkl/R+eq6WQsRXtdklFtNEOPO7YhPIq0EVXyMRzc9OxOr2PSp67
NYRTTvkFTgT9hSzf1lCYeddKk04hquxwEfOsyLDmGAa3MsG+VZ4qobeQw/6cUm1f
TwrH2Nu4X/AfEchrrNTGHWd2hl7PYulEnzznLEKWF3uflB/Clu1OvVJg0ovpX4An
ewXRDBjIROKQbDtpHbWmUznQVJ0Zpni5gnNo2576bYaz1SPja/ypNIoyy7f4ntU2
0+r05t63WX896Nndg3oRLCW+p0rLeSwrnCmC5mDK4oLsNiklLlKPp/i/J/cWtXYe
Ym05HyVvS5Il4ecMde88wd+RWkKd7EBf7yrYfDWj1FUsFyTUPF3a1BLeybB1DU5g
zTEPTsbPw4LsdUZg52NoEJnU/nVBR9FN3sLK2deDtGNOt3jIEQozT3F45JxD5XYW
6KFhheQrwScbFQQCvepn/tvHP9XoxjigJiX4d9qzwfG9r0nOdVm1AHnO2wHVqCSI
nBIyncu5qIiWff7xn59SeCHgWuXW4Ipc6qcqJdmfgYS3VjNUHYzxh7hebnbusq6h
2nrDcZhvzP0fX5Vt9lNMI5zgV2/ZeRgwXqJ4M0OI6hy2eqitoCMP9NwOyIuCRHiv
bupKp+1kwRryNZMiU5XNum+6/ZWge3DcgEhObmCPJKz/HU4tkpn1iXDnOp0FfMmz
sTPewWl3vPYs42vIIpEQQSg0pCzNehscMKBKfQVuYr+1IrhmvUJxQpmb9lzFJfNG
0t+usy1Rd8Rlp7pWBCW84EaOTnTEGvWYvAGE3ZDJCnpJLQdx7qPq7Cf7ZEtn2X/T
ShOu8ZcRm41Be4giI92qXksb2cwwQ1hp+s1eQYdQtJdgaqH6N3wzQEdrN9zgyttd
X/7VoWt9/Xu6PDQ3761tSVBET8af4lW/jSXdbr/sbuAm9gQV91j3BRQ5CU48LtQS
5tkoxaxGcy1Ekp4byFUI07WUcbjxh6Q7FXXfrWKwTiOTx4U2uxnaWNnJhhNuQNxA
1OCTNcYWSK6LTdi0QaIEyF45fChDCtCvBhvIEAxkkBjupr0zL7vXaz5FKzAt0cta
Xc69PFtIOnfd02YFQYzRIffy2kWFJ0ibWVs2dVkm08eNNYWnSEwfKZTUTNAtYq9C
M0Y+JLpSmgGiAZCw9hOLcCRs6I+MhjufxXb/N+GXiGLhIG9fmQBKn4UGWZspl4jG
aQuFnvKNjHYbuFLqz6rjlXKWU7z3wDGn922yUVmGsC0TIrORobXjDB1Ifk39EVHb
xBqTyozNLy6w3kglDABmE8TWQlp/5iDUb6441RbOY8um3k35TyVedWlIl+jvNesp
A/Rk7MSdRtVvLByRLkIW2TGag+7Q+wayPsQsJaF2PmCgB3skJ0wDKSX6OR2baiC8
MBvJsveQfQ84e03ny9jNjobb9yWo+PLtbb/PNY5eEF35GFSWdwnGsPUBIS0g7ZP+
vVf/zTZeV3qfQYOlL6PVnXEYvbN/cns0XlpsHt1qyKXcqzvctyPYUFBtnmCqI90y
M+qrq0Nlrz2UdJPWgbmhP3pVtbBhpyB7m18Wa/4gXAHcNKDr+E2oy/Dw5GgrOdav
Q9DGg6F2e9KOL5hstGUy5n3H7EA0TjacqImEqXHz6bao7Bxa5zwY8N1TJuxAFFjF
B/44PRpEFmu6DeHa9Vp93afXwji28TulxfZh19FdPG0aOuWs3pxIGgYYUewp8VJR
T81/Cf9HFkz2ZZrP2Ii73FgNqWBVCdnajpEaXw5XTLnBWAV/MZEASGv1o5z+eBBL
/zs3am/RFZ8adTqSd+PtVxOQXDYQlzIJzXJoT1TdFh3FXOOda2YkyRaa/SGWIGyG
klvvlRvUJWzNOpUrVoicS9XQW2NWYo4ahwonKRclR7IqbZEYOXfhBoBx22t4E63c
srUIE54pL8gws2pt8yUwGcOPQJon3uWSgRDA4y/E+pCMsYyPK9YY+DcnBTS+x3y9
A08vnIpRfKRm5dzg41Vv2iG4uw0Y1uRnsVK/tfHRy17R6aPkhyWhiF13l89XFedz
6PkvRy18pjfpM7pbIx56GkXVHHNtYQIhWtmGPNgMpi40HATMibnr6pdQNrGuSFWs
ra39BXFubcqpQgNPyb9SKjW0VFP9Gfbafw8MDwSNW5Et0KmbLAygN1fb/StD5Rxh
AxPnnZtdUt+PTHptOnC9X/irpWlhrw8BgMlMTlZm1XR7fIl3Qv2TdGrp7MZOn/7B
b1u//9n0cw6WcpaTCxiutSiW5w1V6qsBqLtsApZF4ufKDzB7gCAYD99ODLs3TWXn
IBXe3C6STzZOejc23w+J9qzhlpoLuuwJmydSkBVUMKPzNQJ2BsUQO6iPEBGvJNav
q/X3pDrdAawuyC8xYnzSLD5YPhce/5tBZc/6jwjitp25NOyuAONA5Me87tb9oD9f
0QJR7rMwxzEzWa4O5TL/7YFfRA5GVjUgzPKZSlNtGCtR1PTrVKS/WfU6+artbh43
eVh7zdZlhiiEq5ZhOM0U4nCJJ4l1iio7NEkQ7V7vii6VZCnZat6sxMzqrWOKtga+
cbrC+Z27N6ILHeTZ7HqziwS3z5meY3TO6+V3pVJw9FUi5bJPSYC+b8H9qrQR3uvF
+q8OiRaKF01x0Ans3SjnFbJGUnUOWCJqkFlHoBQ5qgKkA8yDtUd6Ulj8RXnsAkAs
MnPRd8FdYVq1Q9QUkfuRrb4cZoMgUWwl9qdYVmM21er4ICritRVy7uWztvvgnln9
HLfNQSY5eOrZ9YJRaGdBqaBdmDAtbgP9qWyuqlAN/MqMAbLlYJau6OUxp2r/jrdn
2Y8/DSz71JKiTKUHSkh64MADU0ZSmNnnAU49EYescEeWGbGOGjhmxUWmeoSukxWR
lPMcAhA5EjHsa0GeUbo3By463aK2jwKQCNTdZp4aRlf4rCeuykLOIYcA6tDyhTwV
LNTUKVqL9LIAaS1Oej3Uzakun83WHuekAqU2iHCIOG6MinD4VguGz5eD1MSv9aff
8Ff1UoSzrHyVEghvfPOdxy6hhI2GIk8heqgMnjpjsVU2JTkCvvGYPPaFFRFP5+fQ
oukiBc45jY5z7h47AR952lzGFwdyFS2wJGLOFucvwvuDWdFbdKyXxaFa4puh6Tpl
bmMoFgi6E85nVGqLAA5hmsehm74k183hMFlWAlhqJel2vK2/xtpDoBa5a701Ji+m
AwHm+u3BPgg8DLVaxa6jbRDr2pB4NM3r83RAaNBMjhVmv77CrFabOMZNhsZQQUX4
oEmueISZ5hI3fQkXl7ofe5aUc67/krWDE7DX9PH2clrQkixzPL3+44I1SE/hKZRV
tWTAoJbl0R5u0NodHpvzSByJpLGvqaaSlu9TGbjCIcp6UsQ+Q/1uKjCLfuws3Kn5
aHgIq+kYK/ZsEkMM7HJMginU5XZ+C24C9ZBsGbvTsR71BAc+n1GZTmFxfFJtmTVx
aRUkr15Fb1aXKrtrsVoicve+CptH3ePnERfTwa+Fk0z7TKC91RFYmBqQCHaeFlC7
8fR7Zv2pSP9XiM3oXMd/Z3uwAeXIwdoc5WVsw4TbcJZVTlWIaJ19z7uOxS2cOWZp
WNTZgH1TcoMsU0T0Vg945ULUbPVq1Lvna9MmtBu+vnbT42yKkncTGYZza+7uy15s
ueS95FMXPsSoCHDetzUxVPF117VFofS26nEjGTPj3mmqaWnRbEjEwWANLZjjuM1R
4AIMffL24V0JHRRCtzHps2+TJhFfXjdroyBAK9MTRSsD0FHyaLW/43jUZ+DngYPg
DQDfXozJRYnfPlfQRfLKJD8yqlw1YfrboFwALUw5IjstWNjSpCIU4Bc9muYRRuUd
PWua9biZzPrPNnkeLNXIyHXEmNUYj+FgmR+wzB14RTcYmCkXYpEc2ICLAzrTtdIS
g+XGg2FFhxD2vX58LI4jkXO7Boz3VNlA6ovpj7uyXhgNUnY4Fc9MOmldJWBqC4FL
BWt/iHS3UzWsrIfEnY0JjQhK6qfhwlf8E7VjXbkDQzT7xPHRNI1zkixyIwe+OXRI
53LUoQOCr0wi4r8bKRQw5ckI9951boGxeCHDgRYwS/00uVyimrTESRwve34uR5ZF
qpm9TNqs705v69W3znOVMpbIYn+d4HLLdWHkC1ZWpPAK/bzZMNiDNree4t6W/vp+
87Txvc7NFlf0p058RqG0Gcai3jX4Fx5wHnBIe2RY0AaemCBlsUOiPuD3OTd/N9n0
gDVv8Y3W/k/GZEX9Wy4EkDxpZhhe4jZ5niJa83fxxvh8jtrtNwMvSpvLrDj1YlY2
uH/qsQSJfQ4cVrcSzvWU7BkL0apXe0z5JShTEBfoijVIt/ad0Uhvw0RN3VcpMqXE
89+a20uorIeDw2yGJGTwWcdCnMdUUzK0pcMl0IxO9nz9DY9yB0oH1bbRIXSZa5EU
qrsp7/K28x81sSXTW9waO4yjbtXZ/vslnIGpfTNmNFWv5rRXp0cv8N749zhnp83+
sru3CFiVB3UIVnE2eV8XmNH/GgVHlMcPmD+pWocLHSVja3f+XD7DRZ48yab2ioUE
iim36S/qI7fJ8a5L5GUgpBVa2MR40y0lI2ySdkWHajezADdXbRQxswGLO4pnrZgn
nl3zIvhxPELn7IeIp8WYfErDrJWzixJvOakRrgwR+aS406bn3qkAawCkjHIUAspI
8y+wUpD7L1dzZG9DAl0i5yR5N4VxFdnIhrccVTAtRzOw4aZd5jfQP4c8O1y+V7Su
JXnIRC7bgvE55GctFLTpHUpiI5vSyP+1z/+958mFoMOY4SansAfbe2dCPWBxDwRd
AdGx1UWOcuDwr3gG9Wt9o6h/pOMxkiLgMx+gOfc5NmlQpcVE144Yibx1oawz0VKu
hS/h5mwFpcChlV85cb4e07tP/Nb+bZAAAKX8KLFPLFsxYNtm0g9YwchWP1Q238e5
u1tmcMj8AVrK1ZbzcZNR4T2XFaG3WGekAYCkEG3z/AKO8TtodiRaPxj0h9N8Yjjz
qmKnDe2c+n/yGVh4rGn+dscuhLlY0W9u4K/9V5yZ9HrStv30WMw41HQm9gXB60B5
/IkjePcXSjce8H2hvVmd4MNv9pysM6/OXeHdyXa9sdjgqcdMCA45p1gBbe1uW6mH
98uyino7FO+OlTfH8jbyjwlq2JlHs4HRtzxlkoo9RXiId2YUj/Y3HaG5IX+FVFG+
8nBjH4lU0TTLaeCtdXnDs4O9vk26Ji7ulHFDViHNEmW9vx0QlKS/McnonhBruKZs
kmbocIpydVsU50PJgmly31w+cCEHecoNW2e+rLvw+94xR8NQJgsEH6iv17m4NIFp
JbpWknxvR+ZJi7Ff8oxBzzK65LanqE6cx+A0zP6JBttvCTw3L+dkI1ZzAeSrt1yh
dsSk4DfIuhjKjP3OHOLkYKBlmBV+90zu7yUuSTmm2ofupp+ovbinhsu+6YReXjNT
tKiv/XNkg6E8ld0xrnj6yCvWR9AY+FmwqcDNjYOaTtgnhI6O4pZbn+sG4mhNmWzN
f3vdsWDjr30jjxRQ4Up3uXX1/2Lo/b9n/LyWYmuAhw4n/+K+FSCgCO2aDjknnGE4
xM/ppdnhYZ1Qn16+T+41kXuFm4Tg7Uy0FoHx2NNVKibzUcWSDPDwIeOYdz4ckcGL
j0/Fs1z43K2vm3XhTb41lLmp29NDhlXqIsFu0rJG95xScyKrnvqkxSLiX53FAxej
90Wg7mOk/DbyT0911LmXLIW0j6i9d8fmseYDdzb+571R2N2hK44zyhM44TUY/E4i
3rMwWjRNExpkPouseiJoy5e2FVGWQMva39kp7p0/2QQexM7JsdhJflYighj2zcTO
E6RbCHl0fRPFkv/JhWfAeSHulNQEzAmR8GW1eq2fMoyTFmetdimemvrTiKPwC9hN
ImBId0cU+gVsvgxirJtGGBTUeHxacwSGOvD0oAi85uetUbbm2p5NdgY6stzgQy8F
y2UxDo5bjxco2DSqnz+qlOrq2O4YyDa+kLL1Ng+iJ8UQCXaQWKm8xV5Ez+EeKPZJ
FWo42e3lOQzrwa+DkWgczDnVGd2FD6AP+jrNxphpnuqddIeL0Vq4TLwFjfVNW9V/
2S+EhjHxGre0KCfhHt7xrzQ7TfM2JbHIY8d76HI0zNg7m7HOOkPLf2U94cZzJwtl
URisxegigVAvaCBx1nrA36FLrmrpMkC3rWRAY+CTn2LZvhMUfAuq+zaHaMlsC7yO
9KI3iHq6e+7RwDRkCs+/ezDvlIm/w2/te/bJgJfy1nZIuKTYOfsC9P64Wzl0TJXb
XCncrVM00sdUs8+L5Il2O69MnHFDHk7pBgrXrdTHU5rXzs9CAhNPGEp+M9UWj3ea
ycBI/6P+zrLKczCvpiNXwNTBhUXhae9urbXd7S/fM52+4WMZi2P8Xfxi7xytNu7D
nxH5iosS3qV9ELN7VAiW7+SXwprrWuq+gMUyY3DGobGClJ1riAVUJ2GWIhupD51x
eF4zmOZzIo8JRRaeK451fyiGlWy97ZYGD1w9MpURccHPCN9SgjMdUdEKdRugBLDm
3Zm3L+PMzEOjKZCFeloSyuHIClUH9EcY6pozhT6E+OS4fiQ8mRdRSxiZvhf1gpVT
MKTzXnGJq80srAXRQg/C+40SuWvUWZpF5YsBM8HBc8o1DGoWfENUR8nDAWv18Nmx
24wtFRVRDlv2Dj2CPqxXwsY0urPRT2U0zRnbz4NBJEQSeNpdb3KamW8l/R0KNIfU
jdaNKO8joySHrzPZ41F2yPMoH2kB+7HOwulfCJkN9kTuM3jef2FbITVTjCD1fh3h
BkhoYxC/exps71X6kCJB9O2xH83RF6foo2p+x10JO1wij3PEY5Y1QasbKqAhukN0
Y7xBvWKPlmPmC6UODZLDr/99ag30hlRgt/gZUzYcbrzpZ9BYUD2PsSj6eLpNdzQr
XAKrQq33txejPWTZVfeFqVvy7lZhAtEi/iiSuw1zLu/RARPky4GVxGhcc258QePx
73AxC5DvfYeX4yB6pS2FogVkmtyl5Y2UWThrf18e+pgLxOwbYqMg1unGXA/y/MoK
212QsD6USjm0GCnHmu/3ef4QEXz+ApQkn6aIZAYDr5bAxoRA+UGM6MReAtED0irJ
DEOaPQA0Z+n7NEP/mTaOQo35GLFJpZkiladYVxMQoyWY7y8X4OVC9Phzu1SuV4rp
ay3lZ/YxMWWFbckzQ3nmHpuZ7mwbXLWno9e/5g4AtUDXmhJ1E6JeWDWXVxrPyvSF
5lr0K6KruVyQwTp4tRt+jTWayfY9lNl9kkpFZO2lyv/c4dNY+KawUkEaZHmVxIhK
cyE9f9099I53zPPqD5X1cemgIPfszjEBSCFtjZHyQJHYJjMNdyzelO2gaPnTd80C
71mLBYZYGxf2+/r6OPhLY0tKnaHdaVDeovgj6Zmh9VmyWIuwTBSEffCY6D1BATwL
onhG2yvQzXANBowwUSliqe83qey1VFH0qRTtR3jPQA6hWLzbaGpl1AKo53cA2RGx
RoBzjF2cgHCfI8PvBCe2daLUO0nVn9sIgxgyNR+2T4v7LuUpWcBMDz6ndKOVWo14
2Ov1vDlS4bVOap8pgpJ2FmpIlAebne36NwN7EwwtPejztsv1Me8+HOHb2qy9d7gS
7H6wtCQXzVVp/gTnYdTPHmKHfL2PUTsqj1YmaEO3OGNMb1gEbuIW6wy0vn48Iyik
gmwgtgPucVLWOKY7CPozkI1v6Bv/IgeWc43/QOyeNI/9UnL5HfPL3Xp4gFY/DQPo
ja1Ojaf8ufn9nFr/Y/mEux8do2CbgOt7KQxkgiXwqMDosV1oacU1zI1a7tPVKNCU
B1NVYqM2trId09qgm4bbtINVeY3bbnn6/NRTfUbNcdXVAddvUMb0WNukH7LnmtQW
G9BZ8FKwPOHb890UersgX9JO5DjOC2FLFW0cu/LZRji9768zKLssXE9cnEdg58TH
HZa0NcrXRGkZgv/siM68NBS5gn6wvQJe5FX4+94YUQ2d0r7qdSRHpYqgt/wGqCfE
0+DA+PCLAin0NevZGEBwmAtuAIMDZZTaPq9eNnHG8ZX+eqWZnLfpVHa8gUy+dkHz
USVlGWpyevErbDTBhhEfousZED2hGPjs8loZeDIecG/lM0EdZDCuJW25YW5wN6Jf
A8JPsMMJ+y78FT2k1BSa4vkvclEydkzddvXP+EZwRkteoGBtiVGfQ9gTQ7uN1ggU
bHdB3C6c+UVMN1g0xdBXGPqr3qWsVK9UybodStY73pMwHnCMVeJXXY467UhEyiMK
k2yQPDh0oWsMuAarfg/tPSxSJOJBp36gXLrhK0jO/rAd/mVnaSj5LN4Lvtw61/YI
Dh5GgKtgWpW8epsSgd0fNG/VhHntdl3m9+BpRN/0JzSIwspmcSZqm0R5i95LwkP5
QhoH3GmAt6CXclkkFQvl0MprB0lIoNi+oMitAWUDfjCXFp+Y7CTw2ff/wbt6g0ff
htitenouTaY+DhBQIx4H+ManADiPdUtqQm04W+u/EHne59nIFG+q6VUfSWSSqT2r
CqlFsY7qDJ8KCM4w1LTns3HvkYJjUrqKm8iyHC00zfc/qB53zgp7aJfkEoUUJC0V
o6PR7fdNeEkwn28x9mBk83uRpWnDklIcHRI+V3/yyCRPmOxVIv+6uXQ9wNElu+mt
tWDnUAL9104oy2UzAgw6zqPDlWMDu3/PqyDPJbGWl2+CMKFxeOXqecAOoJf7Q3+A
jwDyAV9UXjeTwszilbqinytzP//8WhwUjbcFG9+4jdHgaGQFL1cGAKJW7U9UUGRK
FLxsqVO1UWisBkWcH/1+sRe9Xco7ZjRV8uiMl3O9g5G1NxsXPE+yKJ/zJYFMXq1y
/dK1Og1VqOFeiCM5kKU8O07kikpTBAIvnjrtYSY9c8iosbaOrfj+rN8fah95Ng00
aodw5jck1FIPOKWBeZZeOt0CGaoxDcif/vAWnCq9UnWPgocvmse6lfxAhqu6tmUA
VAoHsSZ4diuzwdj5uoABhxVl7UQeDyBO14fpMMLk+D5Ni4wPU9oPzSbpxAYqXY0e
ELqxmVR2i59yI6COv8mRS7WBAfoIE/i3eXqa+9vNPQ4Z9wh3Ioxe+R4jiUZDU4gG
I72gzDfB3+hP1Gnl2AmGLZW+NVk/Gs0rxXSFqt6u2XwT2Ht4p0WjuzNUYOvUCMjN
ifspH6uqH7Ncu4krJuiTMk4WZ5YSgcVZeu5ARSJ2L2WBA9PVCG587eacboumRoh/
Mimw/MijgZMfDVfseH/xGgkIsOkZld3zd/Y6v9OCV3vGefKdqj+QmS0Xel7uSLJx
X3ptsCqwlmqHsM7nW+vsOIOTspFw94eyfUp/Yg8kh8aCc3ktKqYRmS6P3Mx0sW9t
kSq4ojHY5rMLICNNNJsv8735fsA+IRyXDcAwNmW5ObIUqeQAKWf1mDXKBR31DSlh
TvS1neXWRbOcLt7rBETq16mVBAH4KkJeMO1JzZCl9sCFuH+w+Em3z5P++5K7kfAp
RtvKFbi/MsbSinFe0wUMkD7g5TnOXQ/rJ36sdZLQqmBnkZ2svai7Lpx6fGvqps/T
ny97G0SA/vn4bM76W2uRTRYQd78lbyIluM0k0TWZXPiVQHhZJ3sDROezA9UHRbzp
ojaQA+eZRpbTczZtDKimn/1SoE0JBCI1tgU/LerkhUISVHSb83ggUPW9sl3Pq79e
f5IMZPaFwIyKv8UyzjAl5SDVR+Ufzsj1sVayW6/9UF1+ogs9OOgM2ccJ98mJPKHo
1p93cM/DpeysmhpB2c71yMlwgjx0W/TNqGSeeJaQJkz/ahyqoyFBmw9BhUs5GYIo
1nmhOH0DuqJJaeU2Q67t9plOclEFqfmnBoEG6qeMHC0DMGP1QCCGciuIpGnVLJqV
6XU0vap2PAnHneHFtGaR2i8KSZtoLNeKJqYEHgBAQsHz8DXMlztxH+povhpwk93x
Wmi9xww7TVZtOzp0fFNrSPWPPrty8T8gRzPlYKDoQAglusA2sbUa6eWbjPD58Zq+
PovTiFic8bZf+8mM1BFyqkIafaBP3IWcC3T8Oxn52pl0bN3tUgV175tJYdYIn35d
dV/40/GgQyI5RXZTf07Y7mwbcYjzJ52QXHL3a2v49DXMlVx3d2Bu45lqwo9HxOU3
+seKS7Dp7yUz7Rz9zK+O98CX93tdvfHpb4qCOEAuQDj8cpEQJFz2+QWYYjmcDy2o
LPOP1lebQXxQXE8hbbyFJ0+qgrzLiSHZSbgBnjoSX+O5hYmrRR8IUUqkF8YG3uMA
s59t+SNSL9S9YAfxw6PCW8avt4+DVKDih8DBD8mbgvPvcoSGSx+RLdpXy43/v+bf
2eK7J/jSv7rk2EEIl8dc+3S9wnZMIIROBwm+5w3pGDVAklhDAr6470LndnIpvTCR
8Z/fqPfb4D8jaLWAszVNNo92sHMEeAExGvt2uq25rFTAUjQ2/RpovLa0h5qQkrGf
XT6653fJ42bvatIW0EN1IUoGSSu+8HmIkayUcMGKhq9qGY0udqeRvgUdHSo2N9dd
FOwMWzG5YlEaZ+XKQPTv0F7KMqditRgga302fRikV4yAyu23/jzNt5fUUtaMpg4K
WdPkXwSzNezv7yJa5ueZVSAAvf1qSam1b2De10/WDAgzEi7vrpjhaGaXxq5ybK5j
9Cw+HaZQ8FoAinRBmdl6lWlxcVtFDzWEbvjL/SUQ9nYn7V2UQXYYum5ocnPbqjIj
o5R6tLGNvuynBoLn9jHvsUzRdR32gPdlruOIAOv75papAn7jNLfrevOxMYtQ1+Ro
C9+PSuKTa0viShQzeuqKkt2PXwizNF5ZSigHsKUJ5O/8r5+YCXqkG/WT2VEs2jDG
kHxAMf85CY8I1ka1lAWPZMFrRpxvk6ezh9CXVv+wvFiwVVmiWCU18E9v7/UxFdiX
VaDwfyWTNcnfkYROyZ1PShAXpAzx5ZECyP6cLxMtaNYhV8t7K3Qxpq+2CGggMHhf
0Cl4I9r4qUaSmCczLwdDDlMWwP9sioRkVDpPAFRbBZPxW1rVXB2CBlg7m4Xny7gG
/51sFAkmENjb+T5U6kxHFPQx0fGevxa2QT5To3cElfVn18rDg+8oMcAtwvDJscCx
HXieA+iUsCvIYHBmAMpxSIPNQD3kpocHBm5cwGBLQBkFIlwbqp4LbgBykRlXMvnt
vvbcWPnZAfrMAp7jiiKbJS/oxud4S42dUFV9YYg0l5gdYpky44D1I/O0BTrAFalE
M7CiIKxCiMO7ZEzW+hzaJZtp7soRxv0uWNRiOODNxojtbsvo/aQdEPMS3DMeBLPK
cH/5YcqR4IgoHQsmtCym+oF6XVPCp5ZWUTdjnkOiX3gFcH3R0E6EOpfuib41cuwD
OLWZqGZfAM4rmZdisHLcFJ9C/XR8tiGDdolxQ/MeW/4x/CjLAOYUU6zUWnfFomz6
MzeYEoVk2um2B7v+9Ka8ocUAVN2SSerGZF/BvCqFRShPc2rnO8xLQzdxjmP8C5eq
63V2Gub1q02TWQk/hNkh9y7gly0QIlhsI9iw+CcV1F6Eik7oqyrSj5WuDY0m3hCp
wfPe2gPp+63ewo8r0hZ7vyL1mZ8Rc9FQzJ1MyBk+JnZSDwWNLCwRR4LzyBThLJLk
aCFISAJCS1CLoFOX6kD5o+PBY1fIYx9IFa9Hl1lhl70KDD6Ws7WYi+c+VoYKsnfo
F6mGwgNMo00G5gnAODBed4AqBMRcaystC18GH/RmkIDcqAxrg6aUW3ttmEA17x1T
VdrB3+YsNTUuB4UpUt7cEHDWobTXWENMGqZgl4CPK+mnPHS8tfVpb4DQCcUbEQpS
0gWy8Guk4am+wzcanIhNigZE49FmPWDqJpm/LqRfVSz7ruvfQbAftwjgk3SV/XuP
yHLFNaXTuYl/L9ia3qyc5yTPeqdLqfjy8EiviH/tsvIJ8M4mXYNlxAvEbgp8uJn6
pODplc1Z5xvEyNM/nctUSgQGWIzKppwAWYu6aZ5Rd/CBCAh1GEtUbU4D5TlPcMxd
z1cQQt2fxdGrUF4yp18Zn+95QSe4iOXIqppHxRXLTsNMbs0AGZIgg/qoN2lUPBFy
L4pdFv7+oweAvl/Mlt8x4mlXaJ6HGHf4BrOKOSwdOHTmsvxM9cAJA2EuiQHumsUl
XZfjhAKVWkBfkObjxUtENH1Z7sR/WaQ+O8aHaZouKkiyvHBPlr2Qbxt8+ibpuZbM
SNWHVsRVbz6c8rLdKYGCz+aAPUDq+g3rJLmjRsSu5+TOsKvxAyn/XAfIF4rLy17C
054s1W9LnP+Le7hh7oLV/VTtgOxZ1t1dJvjrQyviENdu+WC0OIpXBH4zqcc2JHQ3
dPJerKfUvL5CIebdL5UlI51Ws+gs7z+dWoy5H+cbNAb4e3xpNHOQyUPz5y4dPZhE
jC+Uqwf9MNw0RrIqNq1FyxUpJBXFeqYHSNnVH+eaQhW5/mQeIUpDloIeDV29VJmA
mw+HG4VLMK3X788lV2JEezeb9boZFs+gFgRaIEned7TMrVZB1maMp5WNMFuCEXMk
a1PtjnBXTKlGo1lV58o2C7zA+R4Ys+u5tfdpDBWW3u9PfciWXZR8xUKuPQOgIjZC
kyvI0FUT6YbgdmW37KbzXdOzmuD+liIEQAWk4dcUN+10Rz7bWmVi8cLRhlGI+7ZF
ku8lkygxvwAske8petbMe99+kJM5AJGCWTRrddViL90ZXcWoFHej06ndDULAv/e9
TLl3wuY96g/olI5FRqgZpuZaipTm1bf8CwLeYiJal+FzN1KMdggGARfO5wJ51wsv
8BxXaxtFtDYPK6qt7Sohk335veRDY3lXwOZVmtOPL7aXpEv+al0fnIkjZouATrAl
jVcWCEuoRJDrm97jg7+JonRUe+NvAJ4oWoG+fFLhcBt9QMPvB1qpK2tmQlHIYC7M
PwxF947SAixg/lL+gLKADb5Uygb2l7QzIGQhAHqRygktTqtB5eusU79Vh2upZdwO
RRrJYdK2OVzWSw8MAy6qIm45tdcWsBJ3UoWU38BOmD9sQxRjnkNe6OaO2snClD8J
EfcXQWDtwYO05lDlxR8fQeJckVAiM1fERVifc+MlhXeKAovE9hh/LcZhx62VSsGT
SjZ+UYcbcMVz4PlpF7RrBsnCMVd1ZCO4pfR8ytCtntgtggkByWcigKS8q8RhvLzu
BkgT65hfZGB1ymv3kl3Y6J5anGV22Hme7tT604i+B8jBRrtzmZ8/CBIgQOANzy7d
jWJsb+TUPCyVZgoJ77+/7KFl+GRr5u+A56+xtoB/um8C3cHPtL/Srau3FMaH5nvm
Fmitn2fc9zd2JAH4pMlRWYxQ3nFsx0nBTSf2hHxRi01PRmkcNg+WwiBW3V4iaQV3
wZLnYTNE3PcA/6k5LzhcE4Kxl4HQuW+VRNEGSRREvW1cVSY9FgCiUap/yzH9cZCl
NUkwxJPHRe7tqY4gnHShTz24hA4yq8dpaevG57EyK39AV+oUa2zEREMr5Qb2Cu24
AxRSdpYAf/4qC+HjwgB18cbtXYHSAqIdgrADVkWqJHIvuHGU1OlGfuhg47cQRxuo
Wfg1/N6b1dp+n+wBsbVbtMW34kbQICj/yhw7K7JNgmZGonY04rVzQtr1RQ53lVIO
WG4zJG2I1rI65fada2EaCyzIFwGQOqXqZlYs1LroQ3CTsOYLiBchL7AambsEkd3k
4R0qKfeTmAaaRH1My7ftheOE/lxzxSNBkjdt7i3ZAsL9PC+cFUADalnG35qqwhb9
gdlKJ4xGGfW0Ic/pgTTYlSN1B3egln/V605tiGknvTfUa7hIrhsxeSAWqbBUB8tU
OPU1DQfpIMtEzaDr86caC3b9nCvt96Re05vwv1/klTyKUg/iqUNcXe5NJEGJPAJO
TJp7qG61TWbqtlvAUW3vJ35TYWrSHmSItKKwUyX9wekbqXjUECjUDXYhSf7v+RJ7
M/o+/H74L3PpY9ppy70XZuqzppm8MWeoFCLHfRHH7pSe6xRdp8sn6wcdH2vUQqlS
ukpgx/BVXfYy4INb/i3g3eGy+N2hCmGlkQKNbGvo4x7B5CJZEp2sn8Muy2umJYxs
0KBftG7qAOjGXezn+My1WUTtkk4A/5Clv2cvC+OOjIxBHyGWWuAfA+h0AdFth20X
i5mpDWAN2WgkmgBHAEtWZ/mWGo6OYvYobF/RqPubZ/LjysdQAjTSo2EJ5h/VnliA
72NlArayubPsX7Tz5YFAu8Rwtfxwn1abNnZzaL/56/4w0N0UK1mdoo88kt8Z0/Cb
5bu5NfQl4fGxK9Wi/RQw7bHVMuvf6e2clpSa8/MZU9Sed3ZzZc5DzykOdN1es1V0
m4mU6byandIkhHNmVD92thG1edQSsR3aMMwdVfaaNSPG6sReFa1kWYJ+rJrrPPT4
pSI8kR6UuGJAz6B2cfbxDQ7gkeFmYwNN9oiK6EZchrAM1VzghKy0QBKigBgPKZer
C8F5wvq46zE0u14Tu0hU9FeB3bIpe15o2e6FTOFS/QAyX+6WS3QxdKsC4ADJ8LPr
bAzdsvQmaVPhLaJBXfPakD3ukrqCIvLEQ4vTK+WwsfnlIZdakdGKqbnF8De3OI0W
3iBmwA/NmwBSanzKd9FsQfIa/XrgR1Fg+m16R0uSJw/bHIA5XRS5P8fJy+mlV+pc
zgegLcduyi74DJ950bN9IKvemQNUCsG3jpkXYYLwDG8n4XOMPYlz/FMqnqcB5sgz
VFhficYo3b79rUaSxqXUzx9velpxsi3oX2jVW+FuyRlOWrj9nDD/ZXtMRpYSOQOM
AQmIipRXF7ZmqoEPV/XR0255M0dqPNYCqTeeRX9PlJoc30REnAWOO2Xfx+vn9sAK
wSJJOUy3S6tPsOosqCwXuGiLDn1+Vt/aib8oojnseqMHWqf3+wcQTixk21Y7ny9x
J4pK2Ar2NAFMPcn6pkuhxcnWbiPB2YHFfcIi5sAA4y+fo45KQdvy+0lQ9MpFV9WJ
04MfB4cbDs/Rh3wEaUc5+WE7OxxxrFepDe+dKbZkcfaGyLIYAFoa5lxPwIrUStmw
Tlf0b/j9ddEEiVjpKUPhcnNLySitnIb79sjc2KpflKiPhSA8gTv27WGEjsmvbgUw
ROPKIZLa+p9OfP7Xp7Y2Rmozi7IodCWe6hrKFecwsZow/AdlsZPl9cdYEHLFyKXG
BfftJyOzE9LQAD14BPRtXJO7baR6RlJconeJLt9jocRO8yEF3vAMMq2gs7EKqRLZ
v14TvgqXNRiWGLcNqI4878A/KLs47pvqmXHuL2WtwJ5cym6KwZXPGQrA1cC8LRYM
7XZldR54sk0qseLWT7b5uyXkmRw/hbI6ysxr9NSIT9aQCp9kInnH9RgdsfakNOfu
++jq6o4+rDPPM4MwhNhy05LRwxWLTKmadtLAHoQ7zPZef6PUQs3v+i0xKd7WEgH7
9tQS/GGNJI3LlHwsSTyfG92bG8idA7z8L5f6y+e76Qi9viypbrx+3m0XN8ZU0c3A
+9VgDj65OWGkCZRvWT3v4r3QnlFPK/T3VwaRrczpNP+zetVhh6k7nPnQ8oOYMFQE
9RSsSuMwnTvp8Xg7JMSeIm3OQMri2jT+1OblVklx4JGF4Wst7SA6AwbG3Wc+uOUa
8LaGIZ1zroU8UJMyem6sZ5SBjJRbxcO1oiUNcgduzp33CdxIp1jDkZ7n1HqINwxW
cohdnzlsq+Hzj8wCTn7FQIQwZjHkRRUyJFEPUbSdftkyHDQdLLruUCDLbEBX8TBO
lkfHpown2epAjRs5Or2RlIG2ya1l/pecsRMga6dkMXVzIjcotnQDQuqlmT485lpD
mYvhK0Tfcpni+h2tz0wB2TgqJF5eeT6EFFvG68KZ8GhT1+pj2FoGM6eZuuMHOLGR
wWDbP2HTN8rGeBuiXI5JSkVztXN415ZoQ/79P+z1jmyOZLu0g4vf+G46J2deLCS7
vcIfzVAEAqZvhetWDVsqvQSa7cuZPr67pn5HPbo83MBrndSin2QtSkOT7nX3wtMn
RKV4R/FeCwVWQWaxn41B0SNgme/vgdRf1tkoc7GCGj3+jqF4w9EYKeuKtJm+IIVx
dZKp+wsXWL6J6FfsI+cEEgl1LCaw4XMu6ZqVbQ1xA3LcLV8OP4+BftKPBZhQcqtN
RfSDtyFva8wZz7waZW78mr3g+6cc6DdzB9dYCRquyKNRojhI5Z7XPvEm00IgNIBl
FcebyixuQKc9BiYsx/O2n4seks4IZzm3Kg3ZIqTcdZHLgLIusZSFrclBS1AnTmQb
fsMZhqIdUsb+F0lulQkrta0drFlWlnvtB4wXoycpgmrkYjZxqKkULgUnNOySCr7M
uZhE+B15MRgXDja4+ZIJKO4c4B4sxJVsWxFOU0cz8yLsnrLrgqZXySYrAnzZgLBr
f8j1h+K9CuAe0wGBuvGjxXS0VURrBKRzRXPf0Eg3MpWuu7z+VudlWTpKn1kKy5/v
R0UXEperntluq2OsQNtoRQ3dymWwAv9W9Z/k4X7faC9zXNzoGn605jjsAWpQlz3R
9oCPGd/DCI2gYrqNFPF2YQZixg4b7IRqCSPxM2WMjga2Nt5Lf6TLT6zQKAaB+Pgj
TQyOTmxyuQAoOYIvRX4t5WennZcutAwvLMlXD2ona/r9spVY+Ye31jc9ZJjfL449
HvpvgH3a1ArkvsC10VdOA8cS6OiYd9qDDFzyC2qGnhppziLqgRD28N+Bmkbew0Qg
jpXFU0LpZ2jy9MsO5t3xHG9pqoC924kUMuEnDX+biLyQpXFCGNPqITD9knj9Epb0
AtJWURTiFqF+vgCHo4qZ6WxB3VRaVj6k1dJk8AVq+1LpmCB4+V/Zon+Jv5fwaKTJ
qe+5wiooZOQlPu4CSogbmw+gN3V8BrSWqr4a/MDmP+dLEjFp1RlS86B7GVgN9Tdw
TKi6kZN1WmKhxD18RuJR2m5Zz9nQau1n00YE7+wpQXZ9RGWExT6u+Lrnv/heaG0Z
4ZuChIcVgKXp9ExXfQQQXgAJS5IT3zKztHIYD+LURhromB+ZQP02L5TcaOkuJDj5
Y+ytR3k/kd6/oRu9OfDZSx04rPFjo0x+Hsz1hISQ2do17PySUf+59PO+lYfK4Mhn
Nkte6l3++OaADgnMXQ0jJr7pF+a/8K0gTRQbTelSD9vdzYM5V6dO6yOTZYvubj76
dqAvGlie3wFo0acNcuO25+tSwZhe59pufxNQAFxidVVMkBoO9p6lvzU0px77fioT
ftILH4SsPENAEfrAtCkTK7MIP+0eUPZ3HHXoufCh7nUA6UelZGXH2HgEros7x3ss
WYc53+jPRx339cl0AvgH41ICqPTE/8M+jRjRcep5/MxQoFg43psa5it72NG4uiSQ
+0EhzKfHm+Ocp1Dyk22u8QjpnKhY5p+/jY1wAyJ0dft3St1kf63/BzK1zZ+PNalg
uGAT25mGAxCfob9+8p0A1wRwlM5UyfR7xXFBhUA7fTTaeF/7yleBDo835OJIdK0l
pginRUODKZQc9Dh+4KTggptOJMRmFpaPpjTFfJvaQlmH/zYoyAbRekbZZKbIZmD5
Lb9GTbiXEL8tMyZHR8YgK4lvpExXRuShx8bVV2e8UgZmMyN2xOkieRbhwOtxcYSL
AhA/nMi760l6mFRITPaaF0JXhFhVospbbEVGsZ3PJj8U/8ugWMsblB+fUYitXOi5
Lh36qzFMkzK1ffhXkfkcMTPyWyd9oPH4EJ4Hmafz1lCAW91bDCCUexVCK3e6Ekzo
k2e1JVXC5PN584pfEDD1B9y3oQhq1PUAuiw5w/409fz7oZXP0cXgNIdfU+JfDx96
yGg3IOgK3LzEqx7gyhF5IRjhPH5Na4M1bwxvM7kw4E8/p4hDvRpi2FOUf4INfqHK
YARkqSSbn87ihK0PiMdbN7IwwYBbQQp1gz9/Mxth63vkkJuAS6mdbq32t9YCsSGY
EoTfJSaYZqxfBLkgepGUuY6nPZT+x2plzOnd4VJ1lpIXX5XhNqKnBSr3uLEFjjLf
YbgMvzhhAPdviW5Y1tz3Mn+oqsVWBcFZuU+76pVPQS/WJsuwPPg0h1OSx6vb6Ijg
rsbucssqBfWCO5j0DKO580zffQJTXO12XDhlqgPkbuCn6KLnw9n2rlyM00imURJG
CNWt7YtFTcu/9DdO3i8b0ZOBeMawqokPxYwmnuYMqbBK6Y2tdQUUqWt/aU0Bo2pS
IfSOOe2nCnOMn/c4MP92ura3ieF/H3WMpMfEAdQL91jmWmeRb11BOsd7ryAgQOLv
wG5xpnVmwitl8OThG7zBvJ12ghIm8DsnuScl5YRbmV8XUVOLCPHJZc9IvBwRfHh7
2cZmJG2iOkeF1uSs/fkiImh9U7VMNZqbNByoV22/VNC9yNP64TOBR0CeY4rPZANF
OdHH2NuB9sSfrn7yw9WtbtS8kE7cyS/fks4yeq8cd3Q6OZwxtWCz+VPUfY5MdbaP
pqUGkKnbs6gCvgwMUVFWfUcU4/o/vWnOQqr3pJVbfcUmWRB8EZNFdddvtBtoR07L
avndCotmVUnz9iMRnnVrl9XiTZJRJEQQcZRpLEVmbj58RkZUDfQKUd/2a6emErVC
knTmrxhVcyXrAGVRHZHIkXwvfwGPka/ULgYNabp3babRJRYvO/I8j6dMUO0MlOre
siYE49pwaEQKVJGLGSv/RgOkH/vvh/m3LhlL5hHOvXl2Z7983KE1YgoCVykJXE3i
QI9fn8Xu60oJ84/Wvd9MNkfJ02B1CNeXM+LyjBDiaJGgSJa66eOk18L4igXc+Sga
2Z2R3iZnoNyONjylGBaSB/wC/v4r/Ywdt3wfIiF29jCnpW7Ieqbfwy+8W45l2g3x
wTJkd8Mp3sWpBc7zCvNCVrqAw4xURXboCy6rhHM6PzaBShZEdG3SFN6oKEnfN/AW
QyOF9I1NocXKoE2cavHMIWqF7lqopkDO2b5NnKkHrib8/hcOvUTYR2rQw3xemq6W
Gd/BvfXfDs/LK5W8/ioUO03ANrXyX0QtAZS9a3a6Ua7LLZg1Rnd1X2nVam6G548/
a61FFgmb/Uwypb7obkCOhZVYhgYBWNxR/Mon17nwdvpXNTPAMWtAdXEhM7w+5bxt
tBqp7kdQN6/984SgFzLFVbh30Icez24JJaBenpWPoj/5rSAOYJlUkMPQL0J4HMgX
sVrDm6vJCfFtYeGXlgMQCfMMsJzXR2EzgjjEEQZc+xBZxXxezYXBi1CSc73m9x31
l/W/MajRrJxaLtCOt2iPX26hV+DgJw7aWywIDpaqt7gy25+s470RGkagmDXNzNCW
7It36tHvx76W/oUeIQZB4bZjjoDwmlkh7nzcMELq7KfZZuf9OX9YHF73PBV9CRsM
B4H3MV6cJjgu6PLyTzobkbHfXzYAzdP0nJBIID/m8w/4o1O8oht+UKyJMCVRPPdo
G/y1+QvsqksKlIwERuvzdioL7e6twWHTsOTZJ+R6wCtB1cD/DXqMMqS8bQ2W5Lnc
S+PIrQIN8dpG2Fiu+8J7/+sHctjV0j9nMBkyZzfYZVYFVr7rnBVLhDUUS46zJbcD
u2JBdBMCmcSYOQh3w1G676ZilU34qd5IaZs991luudha4eoaUDDpMBQ3+3C3nTHq
iBty8MeevVYB8AaMBqfeZF0nyRL8vqliTH7zsjlfq6Jzan11NaTuVBgPN/m1Ubeh
gLIXm2+uUOTX2Cbj2Ra4CDIsAZj3tjY/YVIeuGFBdbmA/xlRoRBqpL+lC2wagJyF
CNVr4vcGP2NzbQIqJqY3oX2Va2zrqI62wlyHDgTUwWbm5oyMFp0Np+o0w2VUdRDn
mdTZkIZfhZY5YV0s3gr0AetbimLQ0jHYm97aClnus8Mn1mtzOH1ec2gldHOwVJfN
4dFWp1wSgMCkFdviD8LQN4hBRD3g87Yd9rslhgAeN/14OU+ZGg+gj42ypTktKcIX
8Z30NEhPOdq9Ps8+N+lPYmkddbchpfkB7iOamuUbBOdwwmWLczQU02Bhv58Hm3OI
c6LwbdrIpimQZBjW9b2gmDHJmKJc61VbFtzM40pMowJQS5DMHE9sEoqYg3IxjBhv
TLHJabzZ32HpzkRr3oswH/1Kij/o0Jznlpa177nISZF6JgBcFdK3FgSdDqODmVCT
UKWOw1DtcjZrPx66t+5HmKAAs0XGz7kQRQVhqQZL+lUGG82IHL69o7AjuW/j0YjA
m/2XTuBwRZWGFyeuw+gZ+4J9Y/QxDB62TAiRP1zix+6QxYiDsK+wO4BHO70Dypy/
aeCnzi5UrYHnuIRw+ftpP5tCs6+Mgvu4wqRAiVA1oLA2yPS5TUhRzMP+VXgyxOlt
8HJ56U7uY/bQkKkQ10NJBoCgssGvUkDTbe+NyoS3kGnEt60yM4hSeOprXM/21WIH
TBP9ptyvD/U569JBatD8Eu5ZsuacYsuU9Zrr4UNpxCqU7FhHz1z6010/4QDm+AQZ
`protect end_protected