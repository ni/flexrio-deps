`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8496 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10GXbr/0ybS3CmweZF54Xqu03kHEBiampluQJvM5rqyWY
bqzm/agl1dY8diCEIo9hhFYtcCmvSQ56VBR+7UeBqbjdZNv4/O5KYhGH2pOep9XH
DwJK62SXzmle9zw0bgfjZgL98b4AuT/2JCgzgjw0SNPmA1z+x1uwLTXM/F4l1KSr
b2CNk66eZr3++q+qBfQFYDzzV5qkngYXtkXeUGw68ofsqEoSzlDTb5jOJVjfTYCb
3HvN2Zs24QoT5sGpdSBL77FH9fm9SnJoZZ4FCYgruVZafvabkn+2W0gAGyGlEhqh
EVMuW1+lGa5ufyvy9+JTuaHfMgpya7IFnbXIgrazE3c2cNmCfzVk+kDDEbV/K/43
B3FRJQS322isAZzn9UdKy1n3CAJApoTot7Qj6J7D47s69HghWdDdNZ1HuzCU9r3T
B8PGMQ3r9Uvc3ZwZiV6gQ8OeOH6dNZlnIKir/B84nbe82N0qfdKnb50jXPAoCh9V
Ax9IuJaIoZcE5Ml/YU62fxI0WbaIsqHueleSsBlhLtJ92mfgA0lGOkTwplUBq+48
0oxYSkxo+Du2+YH51qXugho/1FGaLKk5/BozfZTd9+4VP70nan/wMqCL7QbO+tww
+fFxZBAWe2eCibXxSL860KIsQN+a1s82wLTl2MfnImoGJaEzCjT0fDizluFv5MSw
3NHC4KgmfKwncEXrqrpXEQvfRsz7qaD5UULrsP0oBGBXku8XVTn1JqujrGzzMEMS
2iqx+VsttdCrj6LsE6ikwmv0Xz1x7hQatZZubHsysNzpMnh7w6UNWo8CJbxGzOSE
j8scC8oYyHQNZi3zmdQy+x1kylw5y6OSagThPko70QVE9T4BeKQDNqo2us07scbq
5kixKCQprGiO4+vRKZR7yuO5R6ToHq1kWspUkigIUenrY5syIPeQXAglcxcAZqhY
Tme0AKDY/JKvSDyaYVOJyUMazWfHGtKoJmHtmM3O5NYrRsfbU6ayfzKSZ4qFSQXt
edXV3xj28x5xFxfCEbslwTAJjfhYWNmluSzKKcaMAuxakCFXdxbfXlVEcKD4XQEi
rmMggbTnk6nvHcXIEdItAhxcsJdjrkbUHotdQAsa1UZvYV9Y2JGhTMQExNWL3Yno
pzcJQkE8mQdzbHHOZ84zA29HJP53jU1EjaSvUaKv+TyprEu3Dpi5JOz71STcHiw5
beaaoDFi6SXi9Xz6Wg/Rbw0gvBStE/k7/PXh4BIzpRus9pgOCMok4Bbf3DHRrYv/
ieq03ckUb7DecH0D5S+NxcZQwNQkr7h/v1iE35pxzlZc/Ob4yply/ZiVnLON65on
2MBW0DgdRDGCbcjXda8KwdEtse4ZTpvvd8N8+dOAOX+03NIjIXX5oYWll3bIM0uf
MA556W39YPFVbWWr0CmZJfpPA1N9wjliMVptS6EET9HtTXC3AL2yftfLMGgllj8R
nZP5MAi80j3G8qIPs2nIOHlocX1mD+gbWA6AzxWzqwPTsOoHVV0e7pR8mHhqHXeH
M5RxfWvy6xcr7dvj+zetdgJWCB4WEqdfB2FlHNKG7dvfr1S+6L4H6XWIghUhEAqd
8I5uEZiJ+IvB5ThVebyp0bX/Kju9AVoUXIRp+8RaCrCPTcWVvZjpYsuuEqOReOQT
42cfIxeSNi0BYYVmH3zwFED7Z/z6ldQmfvtDbBSCCI+APBBwD8JMIJR8iAgbiuxW
9/Fn0rUrnddWFhaAkimR67nqb3ap377oe8OJi5hXN6L/KBxinTlJ1kuCbxWDBpkB
Eg7roJoILKThE0Usk0couquIKCfJgvmOGYww9XQW58XTXlVLs6NYE8nzN9WhS9jE
DCt7zkmiYPDQgv4ynPwU3hd1x1KtPCr0YAtNrUGzLEbtbuApvWikNz5igjnfzJPk
55TEqIXxrMONu99kgsLDc6JYeAVAVGCN5+1vJV3d1cdjA1wcncR3zj0BQrEbbOch
r3V2GTt30nd/hPsyejH8OpcgGbzxvIOFGy11XAYsVr91dl6/0AcAzg5Gx5VWYD3p
V1ykoKSzqogq5W9oO+WSHqSYDfGkrE5D59C7DKyptJ92J5NjRsJssTWDJGFq+v+5
0KQyXM6tWECvj8ApTTJ8H1Bhq0AY6Sr/d8IVVxHNnm5Wc0znK4wr5iUPSxk4Ym7H
G8VRQ632uvfJA40c8iY6qes2cAK1Pm2NhWOFCjvOL0iDVOmitsyxKxE8F8JiPO5c
jk7Zlws0Ciy8vN5AkuVjTqmsuz7VG78sj0cIYCCWYNks0+1gLDOnmi79GlKQWA5g
h/UEMyvh28oqdJwzz+ySMRFWDPhGIK+HvOE+CgsipXJTfoOZIpf8kFN/ZAJXMJIp
0EhKlkKFP6OjexsBtqdnmh+JCQDmLVD2O7J8I6KMVwgWdJOVot8NIt3ZzKsuvZUm
JLHfiZ+VTYv3i9aZrAmWO1K46PyJhFRFTXIsVjasOKXeOFyHpqnbkrXNtdW7drCE
Loyaawwj1FbYvZnA3g4BMT7q9HX6RmsG3kiF4lUc6pyV7HZbzFmjdwIKyzHZSrxz
zHToBYezyaYAkRgaECYUToodDUvuoQqj4t4rtdc2+HT+UsrGuq6Tq2kpKzv4CG2Y
2ZUvX58djcJLFlEcIqsZWXcW4QGCvkXcmWt2C01lkiRDmYV84qn3rTk0X/ynEbYu
1yM3wZeJIAQ25tnzOf35OXYwTcaid5FIzU9hovj5CqQc/zronbbF4C68/APkjC4K
aWqgG1KZytoyL3KrSj4gv30Kte/rT3QAgagEHaaAh4PC2mFJ/OpapxVMPKE3GMdh
fojxjdrtPg2uaR24gTTyFgADjWqJm7d492uD1oiWHrLDwDR/nyeFSUjd74BUwLf2
CRgHVExRAPKojpc/nl1SqkgqEFeVnST09LRx1hn2VBzYzc9MwldDie37eZsHU+9u
k8G/9vl7DGMKxer/Y9fFwI/098t6i2LhbWKGXn0n3WjWmBAmguXEVmzh7lKyfVBU
/zE2owAeLY5dCDxhJ/AVkzJTR7CmoxQYJfn0FMBfzE798k1bKO4NIJbky4GqvYWQ
b+rGQAcOT3vtOxoaD14apCxoRIXna/7oM3ckAZf/DFyLrCi3ezxh8jFGtFWMBrpH
e/5j08dpcgRsMNFhUg6XJhUFzG2QIXWzNZIIFgXenW/ca0nWrgVZ7EzHmi1/MAZE
OzvlK+WaaO4S5F7RR5CDhHVWzRpkeKBiO2oOU74UPX5bz4aLXwpMNlZVOlYpNDsR
Vw8a0dKEnLn29wU4yuLzvIXQiPJjMV+Rarg2VzRhaydj2N3ZK5gJylpXnb8iceCy
LxgJParGqQ9TCVrVgqwSdSRyNuVZLv26OzrKYPaowTYk0Z+8quBxy3i/hVOvLqz6
0sdCyvLWGFF2NCU2G7i6sePL2RoroJ0Sv2jFc5LTaXkP1psNe2ohybmPuF4LI7DO
4v5PIcWhUo/2u8JWzLf+eCSKgskTovcds10bEGoB2Gc9ZR98xAWHS8kxsRbCE61a
XvLI0xeiTpLL+JOjWQ3AjRBWUf/joKwXjIw9lB1UWCDyhuNF2i0z+nH0FLRSv2fE
+0l3ieXeE9V22LGN1UBAHb/n7QfApEuJzJxSuKGSO0Am7ANgEQtEostQ/HF0KOMw
3idC++tvq2zA09SV4K6r2w9AewX5Pk+G+nZlnTAyBFQ4TIk8rTq+qqa6I++8MDER
OCg0YOFJl31DpkuTqZeqffXqIcMSdL7Mu4Mf8/jOrb/mFHYFTY5B7GiDaM8nzjiG
Nq5c4M+dQWuQV5S7PnuID3fbFIZqrxwhRjLuTslxU2bdIOKRjmX/AlpvkW2uHN81
t4f2S2+HTHYc7ek4/GBffaNeE2VSySDHJWbshiVwy2SI81Ek7HkZQt8r7MdFy/Rb
E8UOhxkAKYFwcVFeuEXwl7ffXIhyZXo+GcxLaKNMVogbdh4RV9SdOfm8Lnr8rxRm
fE3UWGykxZ1OEuBdAOFD8c10UMzk9MYbI43dY/XDr5YosjDUFtnk2bXMlUluxB66
DY3VGdaU9vfjcGUT5GtU2I5cdVCh/X5CkqcVdJuF+EBxmQ3d93ztYydqmjxCxLq+
c+pKWFq37SPb8tP6GTQDGjsIQHWlZZoDzEHy8cB/wD8tbGfbbUanIHbmCdNPWsLm
5CzzaICxJ2Fc+JltbLuySKeH8Ck93VFJaAnY2jT76vWNUkxqqnKlsMvPJy9/Ss6J
E3kyHD5/9ihoAS+bnlOWgx15Wdai6bumR+jAslnASdmEcIZDRvGN3MMz9XRbKfjm
Y8IJUrKNgz0pG8yb5aogziSpc0bmIqNc0tFExpL5c8f62MzXUy6x0Vq6nYIthVKc
cqutEOzS2dE+h3WetWtj+lJTx5b0LDkDM+5Gw64xqFjsjWLxFmydIFaDMlWbcwEs
wyrLNsfYHzX/0kqUrx7DGK9n2oVHEOIboiHwpCZPsKLLVjWXG6qHR2je967UeYWX
cOWvLQB8bAoGvYu1RMiqZt3nHN9d+tQAJHCXpLk+xFYQaU6Slrn2kUoU9e90UvbV
GA6c9l6REEjwFy3/vY+FTYy79HrrQbSoVH6vjYL3zdhTSlFcyGlALob1jtD/mY/V
BxU6CwkSzhXQRpNO+NMLNBorKzFP5ELvjHiZL5cHwyk8c82w+qrlU34olXAGCxUl
w4kpUafToVgChNRYmbAHAJ/4r0i2H/y3ZmU7w5We5U9ZZqqo6Hicn3QaVj4jO8Vd
8pElwloL8+NcPr116NWAcElv10QdRevwiFoPMoCmT4PQ67Fj3qJXQwqoX0+E1mqT
8+JordYviGjj98Zr++uDn3TrASkvLJrHl6n88oo8rU2Bw5Y7OtaD0jei7bN9rHfT
VQGO5oqQ0TCKELj2IUTeZif/pPrOjrFCiQZOfYJ+Y0JHDGe54U7pE+CXzQCFXbv8
Wf9utTuTnG1fDnIETqn4Zui/DlH064xyQx+k7CEpPZSaalWpQ3htugZzrZvaWiYX
MgkUuAMq7uNfa51QSp5vRDPjgaVm+FLZXwQBQs1yIqhfC+pP9bbe/Xd0P71ey5gB
wZC2UMfvWOe6Kg/GlJphaBUoCxvNVvPMTVwl1JVjAo1wQrDml78v4N3+z4Jyn5Yi
RQAg3sg3FqoH/OvdGpf6N2QpxEZ0ltxxF7rcMiMl/NMHXVuxJyf/xXyNdsbOxmew
+i/IQSYBRR9q2CsYJObjF/R+umwtqfT1xmeDNl1EYSlXjy2wiRk59RWN6Hbapm5s
SWeBTCANuNnlvs+tsyHcuGJOtU+M1kD8UhhudiIYpESeJqevBDVJXF0kPOe3IcAP
YCWAKIKbX91sLc6rlGQPWM8hIHu8Y+IwrtGMxQOmf9jOjmgBl7QuARHQaBT/E4Z4
FXTyXgTN36qpJcPHOViqVIOenYhFApT+Yju1h+SEONs45kCUxm7NeNuuWzvPT14/
+FfKntAA6DQLcs5OfXmICuHrWu33/+tqLMq5Ixw3oUGN+i1h06D6L1HyLoDrNxAk
OKYh+a0Svq1K6fbEW6sQ3MOuTzmV0xrZk2rJJe78QbRS0knRZXZeIv7cZeAHldJ7
/iUS1n46i3eyKBAzXGTAX3Vg4yPdpOA9z0Oa5AB1Mdr8b9mOn0Qd6jTD/fuJ77mA
7TFLoqA3uqcXjzMsmUD7YM6XNc7skZmQPuw/7tTtIjEQTGIdYagWC81CL6YZ18b/
vkVahDbAJmhgS6c4RV72U9UAJHor20nTEeSs2yqZNSWvchRgGIuVHOcc14AIWkai
yoTzENCcSi6eP5HAflmiT4MU2paT1DUY40ibIulao7fCGc7BscnO3z5UKvyB3ieN
hDSlUdYZlHr44f20iesRhWoCh1S6qKiJU0869Z017J/UZwPBgEAYkCeXCe28YeJ9
/K3EyaBrpuAGTBJS23M9umHHQ7Sq4KH6UP/6F9e2Q7i3FUQFNdFgR2paPwf/UIYE
WLSSMXTIUmZJQsDSj3BkWMkm0kN4ZmF7zzamEonomcQgOcNg2jhBIVlJPYKLr7PD
p25LAWDqt/fVkOXvu1a0dIqs4ZN3zKHI1tHI9OBNImaScwB6PAaFiRUoWEcxW+xT
yzg7vE9XiEcXmKsXXaSG8YLxsmjsff0hqGV1xx7C6dUdlGxDB452XMmNgnHjAwio
r2ZXnm6fTGicPZiqYqk7oa+JegcnQiflFPKx2V6wegmoRb7OWiHK36cwhOaxmlQ5
mjfSEDsIwNNjFQ1/C2FVhhZAKfTzOOxWSkI0YffnaQpW6vjMep3UXYK3w2h84JHm
eVQ+ghxwwphltb1mBAvQh39Y/TIO6Q/BTPaj9a8lHwMrwk5Z5UeLtne8bTD0Y9lM
iW5CZEUFjWc4fb1yvBdV1CG7yd+xgFuk40wHEVSL9/IB6NlOsNwAYMsS9k2oIyyO
mnfbMr+U+4+GZ5rgFUvRY6KGtu8pshA9nAcCFLZEtVP5HrEiOFkOS8yZTV4XGcxY
dfr5XiP/UAekTMZ0HroVOGtnQmMil4l7qyCNRoNXVd7J0QIUaXJqrS1vvWAhQ/54
gWyo1fCQkPPb81Bqoe/lfex4oGXLbCq49tuGQHtlzSWdKogVsXlHqHkbxdAU/1EP
hZpUBcnF2m7XHrCIbVx2XDVp0h9p4tm0OXzXXbVJzfle/zmih5QWA8o+SHHmCN9e
cnhnuuY42XQdoYzBQYStiKsU4AFyVjPUEiot433HEmc3yEG7Xw1ELuiH1aNPrnn/
wMnXwSZWsnRpSvNkYxgwQl3xGrpTnxFpgkBRaSTNOyo+OjLbf3E1/y+db4+D9WQB
PDceNvrxqfQ9MLhtNFNq+6pb48D9RZr5e1FJGALQ2KwDDP67OHROYvH3g5LhZSsL
CGOU+70nawQoFnaOOa9NeZB33YSO4eQt6RvJq11AGNboZt/hw100+06jaBbEtiDz
F8DrOm5AKwFuFTRNNjtj5RgjvhJkqQYqzXThbR+8Hd3IgtgdD7hD7fiWXFL8xx7V
x2ipndSu/HkpO23B3jv2oO9tzZEVw2XOfcIsQs4sq27P2WtjORKbaIlzO1MKGkua
k3cRmSjQb4zaAJAQKTkDpnIpfruc+7F0H8l+Z/EHX7fYLZVXO5NVwhjMdv7pUSsR
0Jx6GyTNIPlqVEj14dfKKQ9pcAmoi6yeHRUcEflPDVafhlzuXhf7ja9XhoVdqQBh
swLwUrmvcWtwyxTySGpQjy9FEEmuE9o4sDpa56YAZWsqAuStNlBTqoZaG5A4W5oH
HJdtuHVa7nqCbWMOEbSNfoNCO7FfcvH/oWtCmy7NmZ87LVb/VfJyl16CtIBKVJFt
xRZBbPRV9AO/+MJUM+bWQwaMFrDzGT4ya4S/ux3FbCyXISYD1re/OJVDMxDoL2mI
mXbkjCziKpeQRX3ilVdViejEyPznXWdGGGJ2f2nvloTi7oQ9ruB4YQ+o8CA8I8vD
Rg0cxepOT+4v8Vzdj3IdwRT5cHAmLZhAFgPbmp52kXIQxOAOmDGzY5QcFuyaDcLW
caXXjOJqL9gl1AoyzbyHDQ6vJWqeW4Eh7JlfFtL8IGEYvm55j42hJwuplckxgPaU
m+zpPz/g3lyKb2u1Z6d/a6/bK++eSVZzPxf+eyj9BL8kuFxyMhU6ow1hl4TG6i+f
r8UOmv3g1yXGNRlOrAuSSt8vKmt5g/tyBza3yU7CIPITHhyXYO3uhsrogrhl/T20
s2GFx2YEIkjNScBBJ1JEHqdwyxH4xo6X2pcqiFhT+rx36acx3TUS7mWohFdoDYE8
FPLG6C1zu5+muRTN8+NpzIQBqrU49e5PdN1MTAFfPVD8VrukPxgRBMiXG0IiTys9
+Va1cGuXu1ZEQ/VdlHK9pY+D+Y0tJyEYLwRHKy7aWbP3LBrI7QY6r2cbAJ+wQMnx
qAID/L98rRYAtNXVn/uOCITx5mg21sO8kHoUdYTYZP800IEiFPLLLHheFEDq4drA
/4S5IFDaLdWR8vO/4+VOmuV0D8q7iG6sZYAojXub2ROcZR0oClrCpdtxAK2m3ZBX
GJH2EPLL8Dl9Zi3m7hR78NVbiU3vMZ5QTKdKJBWNjqyMrx4AuVGLTIe7+R4tNOmv
sWrPhSNJc9btdyBL95Tl2Mn+9/E2MO6PHicWozn3trrrpvF7xQoC3A227Q1VlAyR
RpD4rC7YjZ76EOMnNQZtiUIwgOd3yoiUTrGuXuORyAfhbSekyeP+UGxAvAooKR7R
7wCKij2Sr0SMTA4nuLCrVStp16Fp58615//OrVO/ImEJ0D9qjZY6oBM1KWDAHRlN
GjFUPO3JGZdH1gBKiGbG7m0KPS+o4gYNJgNt8eLp8fnxwa6yqrdlgPGxWf4UklFb
hyyK8Wj7aNOOFs4VzdawzBryoAIkMdbYuBj15YfyWHS6bW9ZF2uwtW36iPAPFPaH
wIWSkyzz5xtJchkgaw3BCsthCfIWQF0JZn32OHLxpv7gg2qdho5rmy4LkGhHG6lX
VDSdYiTMPSMELK63f6Efz7aGf7pEGSd8118jDqsQT9vcLDy2QpFkqhHz7pna0yk0
OVYEXlMyzCEXOd0Wzc3Wvu/MmnNapqiAFgQ0Z8aczBJu2mHUtwmeLr0bDmai9tke
fMLzgGE6fuQjtgLFhS3s/X8BwCQy9mVuLqIAhxurzzShGKeAEKNxecZFKM9lXP4a
q+aaMw9uAk51OuIlPr2CecoEkrHqBRACWn+6qvonXJU7zuuKLCK87hR3sCCoAhFb
CXnf4OK0imq1/u176vW+P0oQmWo/ebvqpPS984Z1qno9wMMwzfX/jlgYpHogPDdS
rb3eaW+kSZM9LJh4hTydmybzYKTgCwSQIf1GCZx8xI3KALn1kjtSufrP9IsftKoy
udHfcchgqaTQhIIstUXLJ5H+f7V0NmLinmjGzE6CiGIpFMoi0MBCNEn/gSE2xSR6
Gv05Cn32kOKaepq4zhcI7cK4/d+Ot3u0e4SrZMDUB2xC5tpaVJHxZH74zqmrrOn9
v3xF1UTITeoDm6rQkEhC5T+qC0B0acM9JvwE5gGCutMlyyYKUHufGLA8PHElr47W
bELnuIFgq5J0Ev8zApAjd9E+c8LQpz69XTvFmYWTvNQyBImb7XgzYL2MuHbTLvYX
K15J36lnKFP9DAiB0SJK+RuOvO+WSSbGWgF7Lscx3UaPX5TqZ2KDSGf03DH7FbGn
oGM+3Iz1pRvRM+4o9awc3tGIy4Azy5qGaxtv/M4Nr0Jn/1LIcFxV0bojok0yE5Sl
CSHFvmcQmLeZ7dyt1d2xDSdElQOTByEhA93bGeUrYiPA9aBOvM0OP8FNfwdNgN/X
2YUoJ0TIeg2wgvk9ST5+/kFMB1FoJyFiZGZFsYfuSRfI5uKKcfbBe5bZyz2RBGh6
0VCEtKFdWHT64w+fUAnyG1KO16XeCHGVWTn/JAEopnUgrRGmA7DlMXUqwicbV4Wt
1nD8pxygWGJLgOnh8mmlg+PiA2vXsWOJLFyIT2XQ07arT+kPIxyl4hK5yZPnB0zw
MatFsSFGWA8UfjkOd4+2mP+q7G2HEJhSgwuMKz+Mc/XCHHNFxh0ukjbTLkHNm9Qt
ncrPmmCRq3QvmKgVXg4IIEY/SnNC+szSlL0NZ5VNRMP6EqMWif4TE0SNZcak/0x1
7y7BIgCKbxx6sUT8hMStWHVicRtE3tX9veg2N6gE5/Yixq+lGPaIoGeCGXY7aVZz
KqjEnaoL4sd8DC5KR4Tv3VOiOFSjz3+swDMitb7t4STb6ti6L4cgs8JevWQCP6xj
Qujme2pNSNqtSrOku54qWMTYM4p89iUHVWSdmjl8VdhTr5m1qpqB6BUPVXEGaoGT
1Xq3Lb6toE7f/gJ1/jrPjvzrnxzFzdXjmyByMAQAUTPyOaeRtjsiWuhzDzJbKWAo
VD1b+XdbdWdkJLplEGdR4Tpx+RawBK8LomV7s/fCJS8lGiQfIrUZIor3wgeaMduh
HmiTEuIXPk/mVDhOXsgLVlSCmc3DV0Quh4wcoBkrdTN0eNcEYNjAueAcjl6Qf9mR
ozgT23vF+uONiv/w6PjQlQIMPkyHOKKbiJGQ4hopTlVuWbOBn9xJaMwHDhsIn2aF
hqbR4FmNzmIsLYnvbU1SMhfjqeUTfCcjnubm2dQNinZS1IVwudN/Cv1ixN76qTfX
ksa3qKUHSxvKK82Q2g9+pU1hMGxj8WFwxYHopqYOlAiP1Sk3hyKWKE214LNhpKBK
d0d7GnOxOk83W/vr3CSOYUULeRvgSp74bs0L9aPZES4zPbXujMrOyLHCNfda9+Ak
sSCHFPTWdtKGfPxru9Ua/YyMzTMfc+BOxuPecnhNFX8rS6lVAAqF7m5m92ohWZgC
w0twUmnq2NU5XFg/TzVw8G8KSjZgaJtc5Hy9K6NWEUQSE8J5QRKnpyAqpH0lkeaH
fJAbDHNhd1XAhkmpA8wilrcZdn9+mYACMwe6wAfpf95Q4VbpbpCZcsfBPMZ0imXR
t1bLDB3DfoKR9h7xcgCu+XKVZdxVGcH4+DIRaCEx/QAiPbnEv9s98t7h4WXTb1Pq
tPKR34bDG8ABkqdDjqAQSQAzNy1vKySqpbtGQDIwXksNr7sCfByZOp2yI3glFYEP
uPsuzpl10iIWUB3I/GA6cbBN5+y1mlUzLOFppwOXsfXYyJ5uL6w3NGrqqX0QaNWU
dzPe26EPbYK2UXFLxSqxCtfZyoJDpm7XrlY2+5J25SOKZISBe1S56o1/MTgn4R/P
GXPy0nmHyuK8nffHQgNKNCTNtDROt5De6YVq0pHRaa77gojztz0EWJKMWGtWzF8L
gKpwdscCTuzbYf/BOhf59uKKVS7iCDy3+Gx2uqRGdZr9xID4w06U2+TC6OEkRP+d
+0twdZDZBEmLfsf9DOpW+5jCANpC9azuDrvKkQkWD6y+9k4MmdznWbLv9mruoXI3
KN0duxBrl3fq4Bv78ev9jZmQdbnk15EQkziJwvsxguH1KrqdDO8uoBqNLMqKktRN
vJsWcrg++5jRzI98RxRaY2eDlPOJROfzJKX05nCj/LxXPtoiEA3RoYtl5qFFfocG
Xr77GkD90rWiN5azSqYIaGWx6ixwEExtueUNZbEFTr80QkSv0S/0RMI3jcSPvic6
LVTaqDfuoTHiKgBS0uuEKIGk/jF6hXgR/EKsherteeFTr2u/czQ2TruXvtpq06bM
+hTqadn/iF1Ck4klaPeh+JBvZ7IvlfuceWIM3dQodL4/t+v4obeUgK9ekZtZhoov
`protect end_protected