`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61520 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
akBpHK9XojjdOyFTP3pOwsesaSjQrMwJY6AOSwj2VzgYj0w1DcS1XKDpkIRUxsBa
2rjRO+ws+P4uHRNV+6MQOvqXr4CGcsF+0n/DqO/fHtnosY+4ag25AnzuwvBfrQDc
IMWgPCLYSjPmftctuzKDJjdSc5nSfP59G8XeRuZZR3rVCUkavOZ5QM9ZSJF4jiJE
t+auKPImO51AeKC9XqAStr/LVt8Q0m2i+GpI/ewj+tT3yjy+DMNDzZkkih5DxiB7
x6GFbrDecFud6mehkuE63mHOgKKIIxybgeqcYW5RkxfX4m9bwZimrNkgmHbd2oRA
u/eyEZ2AK7jjVwbZeMrE2uu0r4wuUK3qSnwxgopjpwC089SI8XEuMLUvFYuMsU7u
sdwICu+1YSmLXrz4cA/0IEnnUanvvhse3dhqv8fbjpuzLi6u9Kwb0vhrq9SZ+io3
YFUywmrAKjaV4sataMMppU7hdpVNQy53xwhEzCWXzSwtNU6V3HKL4v92kpsWkh6T
uhl6vrsq6dqiRNITem8arWKpqrEmH0knkeLKeQBmwX3Hmt/ZHexHlOq9iOiTSZOe
8bwX6f+XrjL+sx79tBfgsrV85+3bjshLRJPyYhRR3vbMlf+uInPRaM/utGKndsXa
nMDAJ5T5mP8/C6PCm40KXogWgMr0t3ITmOw94G/vGwgeh+3f1XzX9n22mXOY9yQ3
NUdAKnhklmS9B359WIJiyfOzy2sAFnONW4zXEcegMpD4AjWhMmTlwGxzmW2Y6Xkb
5c9k64sUuuE5n+cM5f8cf9poV0/Qls+J9HPWZnbjBShigDjsw1hlqD2Lt48Z1MYN
0P0iMUcIDURPuecWGpz2IRLTqL91SUvywLP7d3nELynC8NAcAcrxFr/g4iaNs3GJ
6Uk9LYQbZbybYb9vl/+8n/14B93iQijh2hfjEjgqkcbZf14KyZuJT1Ydgg7pLfnV
SmeieK1GM9jfy92KplbhaJZEfReK9nGftLyGdm3PztlIfhUt1PEH0JZbTVdrY7CM
aHOLOD9jdMgdpALcQm/3XvS9dKGRx2W+t6JLzwI1kN4WxpNRchnG+hBhqpuRS9EJ
UrhQOIedO9jKQOAORNEo4636X8gfs4ODRWCwAHOZWOIT3I8DfikRz4MCpPTfRhbm
UPtPdaO9b7hGCdzukw7hQ9SEXnT7BOzfGASqc9gR1LTRmsAfgWYB4UQM+XP9KuWP
pXUzdWXK6B1qqwemuqBhYeoQYCTZyxrMubYZRUeruoWLHOlKbda+yEiPGxCGufqJ
0fTllnjWCcFdbvkXR31Ko1LvCTWbJkhAhRRCwpyNgyD6O5RuNbQMrsPnMPK71182
YVcQCylxMMljJsKyDwot7R/+HiS8bUYREY0uMTe3y83U+C2C3NKjqsVDWucp3C+z
4NHVY98LvAXIN0TZLd0KR9NKCJCnY2TPzpWM+47gPv9n95TcmC2TYNhj2HPy5a/a
1uf4YUpTFGadTqdjf9Ukxzr2nnFIEfXqW1HutaK0+srLjztlCw2UY8knrZo+lOYc
lT263qSppybD5xGJYVMshA9VhAtULlxiJPHi4PTq6ip7geBe9urpNtMv+HcucM8K
cAabfpPJW35GeqJQWkCIXvgUm+YWJPAlVD9xjHC0FHbifRsLsiLIwjCq8z4/qSb7
HmMildKcjRS88sljXmd08UOShMp0XZr/fYT1/9NIxa2ppzCMhj8NNC62NQ6Cqi2V
v7auVay/BF6N76n5OJ5GGbI9Uy/GReFwbdOIoUESPM/WFsM9L2ST6PfWc3dJQwMS
aP+SFUaHyDHBoEhow9pFkUgwuFrh4vtBex41eNfpW9l3omAsLuHxeVIefQWiMmmT
I+RYSPuq3Gr3RVU46H60KUDiDPJbDevwmpTAJoqR3Mj1mvlzHBLupQUSSohK2fdx
ct4IZLh9ZT81Kl0r7oS5qwPj2yq9PaS+NkemQ8v8DOiCGUk789qX1fMfb3R754Sf
HoLRlSyIfziS9tcv/xOp93T9+QVmwhhkdk03dg1F/5bDIcmaC5IWWwYCa9+Ehk/c
8aIIP7H3vzX6sK2jeaow3vHMA08tQcyNMis1fk+bS1On7BceEzvXjjez6jK9UKRL
hgQpMGJHzTdqJCLGqV1BfAG5CI3QkuBiZaMGxkqWkQFukOQcQr5+C3kOIzgN9jMi
iQzKvNfYWNk3xIERt60BYpUXHIUwhysZ+3ypmg6B7upKaVOwzEX/xbYqZIOpOITI
Ypd4YkHRH0udcJEL6a0Gno2zry2SCof19Qw0SvATfjnFrC9rXro+y+TimzNRrHLK
uNbuDPR5egSTxUg+H9TlVtZXm+k+MovSUZ2T+96FPAwvLmnaSit82OHzoSEJCy77
2qdy7X3o3dI+G98FWLawHSfVQDGF1/ZRZzUGb4IYv8CLZMvxlurLfolBjm1qwwwg
YV1RWASEETbhv5tWXv80q9RbEpsPdgJUTOEyMdt515WQNuT1E9ld4iuQZqqughvG
HepnqgW/VSPqhMDYBOSAYitXng8A98VqJZyLuAUBaF/nNIfRbX0MFK1aq1V5XSyp
1Cjbp+zcpIVta/jyoHnJJT7ysf5ED7EpNYCVoJ6hXhJg2uAPJCpTpaioy0hC9rQA
R+1xjJZEIK78CZkbYndOrtjv6o3TRLn3PE8JUZBqSN4EkbpBB5pK5QoU6wJhUAXx
e46RZdY6E72sTVFP1HYNikg7vqlbM2nirRxsg+xtjtqz41Bg8dplLSI97K28zvwC
LXZoInGI/CsaAVnXKujiSryBhhnfq64nSvKJ0xCb3rP3+MOx5RK6LTX6jPycKTrO
+yNd14B7Ubz4GNv+rJu8+AnZcM7RnwCkroNneF6ZuKbXeShcGSwcAcvIxqaku1af
/XT/Ktk6amf9rIS1aHytHEA0TqTBuYaCC/nJUCOg3gX7nWVd6EWNiNXSD1XKeuA8
bUIQyXUh5heAG2Zt0azc9DJejkz9YCghpJoYhrm9I7d4dDsHmUPBhZXWxozjrcC8
o8GtHErOlR8ZCLYXo4ETsrkAN6/OPUjlC3gsvhSyLUG3V4npXtghWC/yDv4+0MzN
ekOA5tfGE3EzoynIccQYRzi6bEJeISBDaoiGJejzr4O8QtgZiYDn6z1PvT2EaFjx
AeDfYPmIGseLMbc6tc+n0kJDc1atxePIsRBg/vA3sjWwPTiUznf6OuhevwYGguJm
7iwvND5K2ICLHzZMoeSZeYi0Nba21rqh79E33bIqjsJa2wL7EPOpCzfRwIGO0iYU
szLiZ2UsJRSL6fINw6MuF9nSxXbD61GdNJtG6xNdcb7gowv0z0Mud5YgJvojQERi
USlvAnVhIVg7OHvjQUNXsfJKB14Y7OBML7ZMIzqzMq2i5tJGCOk8Z4YvHnXkjtF+
mFSGhRoFe7Xav6llmy57aJycKuQ1+0v+nXsD48QAb6TaCl+4xvQw5k4ztW7sFtSI
3F8SyafvWg9Xl6qA0qGTJlTTttooD6WfXG4/jcW+Q6efIqotS5bhDeBTRAsT4Q6S
GDmHqpIA8bumo+6FlhFNcHZ4J5AF78749OT3g9SYesKWA/98KyxmQEPRNYsWObMF
QTRjd6zGrfTAc2gpDlFxQRx5tTOsnvFVDvCpKa/yqYuGMHY9y8qSU/Edda46n048
ebZ9pgwSn2dZDQxcDiB+XAPuSClDLUeK73JpNWPp3R2VD99aT8OQNYQPUP+c5kBh
vxpot/VPJpbPeszuVjnGxwrLzTZqeFgAPQKRVRZ7DG2yGw+wCc0tt7HXNVjYlVFX
Deav6rmpMtwWJgrNwmnob20YWobUYFJRrAqO1I8Nhlj5NHFUKkR/B7/VyrwGftLD
FOugKvfjWHu9g0KFKs4bej3cRGl12q3163H0l+SeqwLzp2Z+31nIYya2G1waDfgV
YSlRjdMqExXloZRJwQYc+aqWYbRowRyZnzA5qt/NVfC2XJx8MYIgCqbIhF1zoKw0
HHaxa/5V0JrApoRdpObRNzQsNBkqGRPY3I/y31d1LxwxO9aiTDsZk8qGyLGKu5Z1
BLu0g87kD2s9TWrLGXkepk0y/LlBgO2NjsLUgx7eT4XsbLKBZqQ6z3vEItuB6c19
0PlL1qjj+iiWM61i23jtBHkzKqNhmPwFXGIlvZQlzIVC3soL8bks/yt7WUjXNUfx
hXcnpH49MfKpjY7vmqW3cbfMqPJAJK/BZqp7MGvDpjrXN9G5kBmNjukumJF5Y9Ra
87AYSx+gLMAQFbk51Ls4uYf1pLqm8peHW47EmWJrFwLEQgKARk1UMjk2UFlSkNxL
nqleunMRH3Dvl6cTT0H3Txl6SSiQel1n5zhXj/NsvtPLXfu6L7dtwZd7o0trMO02
1Ciuzgj1F0DoQsQBKZOpd/1ufpkZ9tD+K44n74+vOSr2F9BeY4/Gb15MCdgAp1SD
hdkId3TEodoM+fP5Spe27TMoIoJpSFIriBm10aqMLrNzb2kF6bY+CMNA1TY6XMrM
eZ5yjG8mj8rYgZILMtW1nTNGByX4jRHvooQZ89lG//2M+JUYYZOygTgO52m5KXiR
wPIzrqBUxNVWBfMpleL+sshvk7VlYXAsBhg+n8CrNqfJSX+IWZmrcmK93FnXVdrZ
E5ovNtOtwhCSMfVBj08yxdUwHgEk8p9eBBoIbpdPeQfoMSqbWVf/BdRQvTY/7jwC
FwUZgddQkvlW0yFv45+2z0U1a/ey4m/9CWdtNJIkxdIGUYYFk/c8wHDFoHiGOJum
VeV4awxYk/ZrvX0YImDKtCsOj8OP1qpQhJA5NBjfLZdfLPg6VigU6PLr//qrCtNb
uvoQDJK52T7xAU+jEZXYpfhb9cFq0IaERlhS3Ks4wwNmKdktAeFniMnB1R50Atqu
ANSb8axO99KGQOvTnDfcpgc3OAxnm2rWr06HImW0lxc4edTHmbXoAiuCO2GHCA2Q
gpI5b4gOiAfrDaQFIw62T3MbNuxpVg5hRkLy4bK/g47e/NrAKxuEulpEsBI22Mrc
Secq+SSkZzGGfvgoJsDok4MChnLlygECEXKcqfc4JbJQ9dJ71yQ4VZtL2QR9UfzU
55h/tIa+Pmy3uJQltcoLJiG8wT/mMWV2U0yRzPjxI661C2O1GHRO1n/Dt2BWtl4p
MLb+/vmSgk7PN1YnADf8XX9rnGLNXeWvNjASv6tLqAq4xpiJn+qfyExmHYoDzJJJ
+bmWVkHZGvDcimhM1mmDjAK1Pii7TDL/9atlPd+KntQkkwx8rNyyEjx9m3/uxQrN
LHRaOOt3ZiRust8/3aGFt93y0X63kNpnJDirJ/kU8iyKC5F3OQpX8WfmpwzZvYnB
4Dodvw0RBsL6TXkYlZhxhB5PePbDQD0djD9anGohoieUzsprLDAP+WD92E6H8e+w
O9ZjkT0sf3npTS+1urlpEuRwm+AdTl4GAmHgCIL1mE1VkLJeng/+LUFhQ+yxmSf7
orkbqIVOIUC+CWl4PNWA216//2Vz963yFpPwEAhQK5q95v2RA5Zq563Lz8EkE79f
4RFfxmmldpVUOl+j9NZlIusRGsUD8ZHS7qfEUeQNzrmghk1QwZctBV1VVjtc1rYV
Z013gXLmpbi/Sdfm8r0KC+ggp9fN6mCNzYb7r4MnGE4Cf1loK4MPXYN+BMzj12eM
5iByrKBwb5I0IsM5J0YGXdpDBKyhZf5TjF0FynyqU0T1N7n3uCLf5jlG5lfTzX10
Y+X2ouQrwXDS8tKUYVPMEJNpSsC/JpEcfl8f8eZaA3nLNbXt1gv3a40+pp7raZ79
Gz0AROrph3ijesIJmpRF8+Eeq2kxGkvkqMIyFJaJjMS4kdYirRlG2JrmR+Lw0s5b
CtJ1qo8nPN7Rrv0RTOzncAwa+LApuz/+YVpF9qI/EdIK/nhmje2h/5zKF9cUqDCC
mkJGZ19tp2tRBN+7ofd5txxDJcAjYDrLucv5iuvAEK7vYdaa2jOb80sDEel4nHPi
Dyy6BJcP40tpECoSjZm6iWMljmZV4HjRceeGSANa0ba4BhHoYQU6sf+N4bFYixsy
yqtrdsDYMtC4GA8NeR2WJRrbqoOdWi1lT4qjwZwi4W7F/nVEjg4xdVcCGDiczjRj
xC1YoF7Xaqida/5KFLJpHmvLJwAzG9lMqhUPZcKOIh0c8bBRhutc2oObYm8kkaBi
cVaE+IV1EUdO4PAH0tVrGVVwPoG6mCvMezHbbx49IPYgpPM+VZIMWGSjoHP7dGoT
fxWSWGe+muRixnEDYCC5hwftvOqkUQsbg8cfie4CV0CiwPRhyo4Ql4uWLtZQ8/tx
C9yjfJYCgl9+5S/o3dh4U1QRZ5VG7Mndhamu6mf7FpT2cy3u+KuxPVKIzRuu98VQ
VECc3pCOwb+dv1wJR5Gssy1rTlDFkhZ5P/wte36j4ia0WbPYmlRCmIw0FzW5Hqhv
Xl3SnoR6gzDxFRGkSG7YIFLG7oY7mcY++Xw3se1ZN2Borubpy24RFn0JwNitRygq
+qDmZeA7xV0Wb2bSUXWLBTKVRqiKRXVNSR9Vp0s/b/8m3PO28+PDPyw82lR75zQt
N0mBCkU0AG/Qve3c3jZ0jgQzkLbA//wYeymzUdiaGm2AnfQicQJtVCdSnrnruLIZ
I3Gop2ph0tPIlwjpnTDoNQd5q9XWapfAaJPj9pIEfEdl1w4O3hTjuyBW0W1ttJ4/
jOZZPyJPlL2BIdS9Xqtsli3JwHxJL+RZ39ocwZmlWaekxaWl/kLlixyjCgDHjv1B
e7ig3TpbKt5H3kiTHf67tJeHRl4LPmMqpULSmKpYTAdtc9VhbkB7xb6O+7OpO2Kz
sWrelnTMOr7YREVfwWhnzt4v+52YsH3C5jThbaZ2rRJMjoEHgNZZOCLwdwdOsbRs
LQssahTPYF/Vc8li1nHzWclFplgI1f/LrkU/AjjBq9At4Bftxk89AHPlzV0sETFj
NqZyu6G46uNHbvBhsZvInEn2O5Jb9bchbVUceYJLeUdCLRxIqh95HX8dK00cmS8Y
w2UMbAhepZJe62f5ILx7l4hZzBDuEIp174Uqs9EdOGBxXyTueiuoW9VLTlgg8WBy
xx6oXv8Oe43kuHlOufGFRtsoizNLNcD9LSDlyoiPCE/VW43V/GwKeoPR2wBbKHeC
TkVjJAO5/U5bF4U2XJv9lTYiNuFvSGGFCluLQQ6+rNfrjbIGzXoCtcpXp00IZCFg
HrOdIe5zEKaUGpKpwv0twl2ArSEOQyzs71GC9FrCmvYeWxg9P4vDq0Y/8Y1vUZbR
Y0xGpmiKOXEwEmXHWeAuQ/7iORjgrEeheKuZLRqKDuj1iUxcw5n6dGVhA+rl/2RL
0f97hC9koBZKiLCFKnSQjVSoL73XN8SDc3UDOdT3QeY7wvTU6/YR9aMTISJ6+UGi
MWpYcQPJwq/dfoVvK+2S1+YZekb9jTVLuOh8R+T2eN8ra+cow6+23+8OhxPmAmC/
nMDIS9rmMH1nIet/E66d/ggrBBqIxvCHdgqxqXhlB68gnP2kblUNpspwfHcPK0rM
C+u9DsEAQLYgohE5mOImrTJ09QHlHPmO2kUCTVsvJUUi4lkKC9jPISvtq5HDzwXq
W8Txy6lrg9ooqLzL9a7Ugvy8YUqPPD/+EocxOL8NxQS+CPpPSwsIAzOfM/9E8T0O
q+QbcDPgjCguBx28+O0AwIy8kMVZMdF/qbILEIcJ9KJ1sXj/eVMMu3nbcyeFk3rI
nHKEU1mFQ5/dPBOKBsohuyVjcETN/wf4knOaFM58KXNmTx6mWcHkr4XnDjMGujS8
Dg2e2shr1gqrtnFvTGW7hxUY+i8IdGEnRBnb4udxMimaHrLOurEodwzNsunZ1PKT
CPrv4kyjAtJdunU7Hr5LVu/uZ9xjLToRPqvj6FBLQD0jKx7/SkTGCbjZmUzI4SMf
NHz5byCupVVwaY6Dq1DrBdvqlDWHoYvrc7CsSkbxJ8uha+m33PrUq+wkmqYSjgWp
dDHz3Z1LqyF3cem4cuz89JpGSEKnqFasjFqxcX0Afb4oHot/1kjTXmWLf//NtHsV
P7EIN0g6ug71FmobUw/izazUxLKCKwOBULVYilkWWjpiBOkZQh3uiB4t0oveD8BQ
jyQRXy+7XAuVsRP0sz9C1U8gtOP7onL+CIOb2ym/l1vF7mWJn2h+ovPvJS0Cs+Cl
VvN7Kv1QXrr5Jxe1/lsQJhyRWiYBd3opnn2bK5MULxOTL/7FaxtxB2f3gY8QHgnd
k8a4NVM+Px6ra1gdmPyzZcJrAdUCXbjinqcBeTTvz/0TU1ZtynSg/J994koPhpzv
6dmOK1/9aq24hh9wEp90F0YSAj6WH/iKH2zoI4HY9K8H0llgv1J6YfyCISXCNx/F
vr8uW3wNjJUMT/Hbo3Ozn/hYgVKoYMIbwksRgC+vO8Qs3w/uV9P5G5xCaQsvCXqr
K1VLKGTO5x83jGmgXgexj0yod/igpcGenRqNFwLPAlVgd3BccAatoRzPWWV4XhRH
NFy/KAjGEa9DoghAZr1LS8hV2ChdrdtGS55qHIRu9UpvfsbGin7pXjITIr++0asv
24OIU8Apx+eEjycPDjmhJMpG7Qmo8nH0BQwETaerxw/kzewLQnuTOXkMw+7ebYk2
RsJgoKXgqCyBimmAAtLNZTpVPz4P17ABGEYX6Y89bKrWlTUuaR/XTVrKZo9rmYxq
ALF8gjVHYOy3Q7U0UrvIXvFttN2G4NdntiSb49K1gPF3YGk+4geSdt+l+SRvOhUo
9iDlPiQ5gBGF2vqEpkMq0sefb3Yy2nV/FFVqmNILRycPVt4EZRfuFY/2kPojMqst
IwMgBpBnCcrJXoEphGzkt/RMV2xiV6FApL6END4EUGDEmSgqdW+FtEkmx/yp23i2
btQHFvgytY+f8ILZ/PIfphJzJ/LtPGz4RIE7wiEylW6vAzYATzXe4snb+cnLIPxx
On9WSxeILyHLNpasHHXaof3lqXfInVKrRUbvX5nTOuchL/+NTczUl8uZlCGPiAow
5vG40L6oDzsvwhIz1NNfL0byU3pu9CqvVv6gjRdzT+HsExgTucA29cdtMoIUnK+i
2hfttmfIUWkgra3v+0Pg022MwYpe4rPE+/fV2gYDtPhk13gLI6a3V4/bn7eY2r9v
zJr+sFVVHjgMTlLJS1yuY2El3TQCM8tcghB/yzumQl3U5dBNuHm3F+eQUWFfqKwB
M8AXkozXCS7GLRfgJDt8pXtg5iRYQ+LMFGFBllgCrUR/y4Fv+2iMMYVru3OZKQGJ
2WqF3FewpreQwcRD/cm5ODGF36MOH1dSm+u5z5emIycRvAvXEr2IPR7G3MgGFDml
JPQWGHL6cEHzZOkDPbjTYxRSSxnGK/q63r/DOSG9NPyDgd8BDoJRDLnSDvz+AaZb
ws5MSQNOL66Ly9Y9PEAQXMGuSgEyOi16cVXDz/WcdTKW0LPidNKGABBYrUhLL/xN
jTy5sy0n4ugO1oykafRHHdNE6XdD3aaNzm9XR1C+6QboXCI8aXXwMTl/P4jPs8Z5
sidlbyhMYFYTLvldLqrgjTlOAU6UREIPeDoe0jjyXaOVmajXa6DevAZIvzTqtTCY
+0kH8ZyaqApjChE/sAezDAIfB5wF0NIWKDqc2nbGlMqn1+2POw6zYN9sIUOUV0f3
EhaL/JVd7YY/XBk18hAN8rJM6GQmVCz9GoaAh2FwgTunc3AQzv9E491pdUa6ndau
lULeeyNiraoDxu0reCV0of7+km2ZA3F5uyVoIYwRePOkBinFomQ+gb1APts0RIaW
h+X0Jda18SyHJnze5AFMNSB7pxbiSr4l8QXAGQatXGSzUqAyLCRhdO2G4BBy4yfY
jKCC4hWkCCSZNEZ6ss0q9YAaAdZSJ1/0q6X5tqzVVHKkFaqfJMMEniKrbgWdBxH+
T12Cq5I983shNv/o4yQKOVfXNGJ4s6shjoiYRKafA4tZcX0zH/YctG0um/Dfk6mM
kTOoj0dP1w6ae/4vzgjWIE1JmasiNyE9rh9ul0rO6wta2KZMdpTlszoHGLC2nbzt
il++gWsqNifZocn2pWWXjMjYHsJvlSbvcnNJa+gmtumRSVJ4zJkjTsE8yhaPFMEQ
41LGQToJe2/kC5KOKlE2NR+p+2WBhE1KH+GP1QBD5YeehSfyYYBQe+x8++GGbfNN
bsFfgOqX6pFZfYSJ3VD6KNvNy/SwIWiyLvjcpj0Y9TmDf0owAThbjs0Z4Y5A+SW3
4NnJbmHHAKUILttEKarGyxtn/lcV1Pd3VmZC6YlsJ2rc9IbxbNAjuzPU83HCZC/x
B46BA5adMT9xNpqWgwORo17asl/V8SAF3aFK5kch0NLAuCrTDnpd7P66EjbzwuBr
SDxLhMue/R35W+xMJcCer4nHCSxhTT/mU7QnxGLu4Jh2MTzLVRPIIlf4OBDLHWWB
OJAbyiutKLlkAQdhQug0MW3bivGtuuLfwRW0+2d+qn8wxK2wPw/IP2ELBfYA0Zd+
DRkgok5NG9m0QuzPdivhmmDdrAxLqjp59n1DmIFJVEpYgPTcRweF4iBz7N4MrYyQ
qQmGqlancgr4QBHT9/90pLlmd5HGXRSKP4AHBIxeVCTlIJof84jAr12A377FOHCP
U6tfN0oFJSc7iKE5yEA3hv0RXCV5wlr0VhkzZmChjZrrsLWsRhw2nqKtp22x0qUY
goOtSJifUgzLMlAY4iqeqK70GUjYLpyA4urNBjmKd/TDjNXTB3D4Pv+io+s37uBp
EMCT2IRu2KV3nEiW201QpC7mz0ZKvbV+ipkj1JHHZvchfo6LmImLYxGmWbUTbNsL
NqMz+FudTY+QN4ejPyOhnUiouqdGZqpgB3RFmdebsbGQc03ZqdOgC1Ypfzr1loGM
de33/UC4Jm0JS+P54lgnUxafruBUJkVAaB6hfPz2UZh/qWQ6u+3bsDLT9gdLrxNm
42yyWF9cuPuprwuPo6R+O1ELFpQgWtuuB9rBrfKRJ8nFzRGoN6upodfxlsDOTYyN
M4sh2vngwWOO5b4J8DjeeN6qY3CvS2TD8JXpdw5ZD/QUxI8kmRof8rdqFlNdqfG+
e4g0vtmb2ZwEn0A1EzlicKCXC9wlXYUM7lawMuh4ATZokLI5q3oRn+sN9kHeTk0I
w0pLr+Svz3sw/SiplhgikdkZRN364aC8Xz2TXFImeifuT1WEtDTqM5qRbIVSQBOe
dV7tcPnaamxidlqXhIztWqz11+7RilF1buSfO1jHqJyH8DFa/LoxFa4y4TXghCbi
1KM7VMLTons5eYAhDBnJXlZnfgaPDNtr1RvHyE6HcbLGYzKp7tuEO8S9FLOkcs5V
NRvkexg1orehVDxWG9f6P4xpWn19qX6l0mR5vKdUjvd9MzGMMP9LednnvHRXuLZL
0VONsmBAAcudcwZwSpWJtYG7PGYkv6QUvxNW6jsEc3fdgoHV11zaIWbQApSZP2i0
jOhLdjtuEN24ibsn5/+10p/ZzkYyKU75TcAwJImn4BueQk9jULul0OWYrNyJG+NU
JI6BChXKTpXK35Q8oxVk11J7KWgcAK7dr2YIP0kdsQ0pEnEY5vQoBqO9dXRzqaeu
KzX72g7FK1xON9HUtXd/Kv222cICZmIBP7jgwuQwFGACs5eFCJqC3MC2Hydz/0Nt
ny066Y9ZFXrIHmTdBpL9KNjBQU9RL/g2ZI4HZ2RYcCl7ZcA6sd/AZcJVwP5GwdMY
kLoQY/6tDUG+kjnZc6pRJAWzJI0FjazD+B5w5BoE7NOzliHK78ExnvJQ6JLPtnAa
J/C9I2SSUWj2UD/JNOeMbYF+8PYcWJrcL4T5dXKVfjU5KjEcd+IJcVGS3eQhNHhH
QDAO3WEuSY8b5ikoE/dqpdM3f/9Di0xiVOkIPl0GZRgKFLjYWaY7BLSgBkJ9BTr4
eRIuhLzxDahSDuw5Or/D/9RMHJpFGqqWtZYEl/KFXYtDUV2jSS8CmayFSbW33ps1
mZSsrzjbbJhZwmv2mpSntHLoIXGpullhy+Ry+hTx5N/Khq0tYfWbafpK4F4jhEWE
3OSfdYVxOP7CxkEtZHlUecnTeyo6Ws4JbQ6m973SkaLBXb/eSJ4Bf5L8h2PBJujr
d3bxCuYNx/fK/ZmyFADYFPCXn7i3o7OY/sWhsmqd8CsTgEKh+fXVPfl4hpge6oKF
NuCHmlOzXt4WqhRFFpHZikG7mS63TP0y/8jau2d0fCTKglVdtf6BKUqp6Iorwiza
GzxpkvNaYkd8Dk/YYarM/BNKRCOZdD2Q7myCiSKcclWKuSfycOk8eaCmtiY5akhs
LgD0OE2r6TjkAcusQgS2qjZfSNLo4ydp+tOr8bpfjnAzquoLFSHjonYyrIxCOz2T
p3xpBGW9AQpcNVZLf0SyB7A+l2uXFJepE42rUIJqFmUooNdxeVgb18n/whwcevVU
mNUxPGfFptqzQ4ZiiIfHry0Bl1PTwFyb+UFZSVo/Ce5h22GkVK8b1gZALJ8umuSq
8y4krAuKUbZ4cUFAc7c8oFU9Qr1cj/mAga7xAeFrBFvpxMqbqK4gxBtQk6EN6Z7I
I8gY9zWtjtvYY9jm5m38VUg3ykmUNLd4tdjk1+Y+KK7ftnNyGWuERacbDp/0cFSZ
R69y1EYzw41C+jG+s5MfWTP0w9tIW1ffDmN/9dYWGYspR7KfQ2Z5StOkSQhw/I7I
7W6/67M124c8ibFpd5dJhE+u9iKpUqEyiHFBQySqHq3seo06ihFoXQAdlHObScmE
wk5vr7FfQbpVTYoUrQkBCvbKfI25qhyCVVvbQrO721gqxDHEZeS1Wjc93uarGDwB
LYCumRUfdh91ZO8mueUqyNFQpQVE2lD6iE4b3wxu1TfHlfXPpvYn7lDFbfRoz0T/
EO6QcFf/f7BW3oMXFJLXsN6AYkuGnQ49QDAtS12qeJOKw193hYzoYwcFi7xGEEDP
G3ulZjfuyFtoF/6yeoBijf0/hmh/Ek/dF2ZVbgK6OWDe67iyU1GVBkry1/8rZ0/n
7Ch2udOMNK3K86rrmBuduvj8AD+kVntKckRwBX3HgKNh0rbRBGw/2bPWoJ514Z09
WQCiAMojldr8YexqNxS0rKa/svi3buzCe/9+TOb1bgtOy+zqBjcPByKatDGVQ2XK
znOwUs3rg38Af869bpPZeP7Y4dxOJIb0eQScU1XaCRX8vUifOmpKkUV7E1BjGzqa
j4RqRn30KZJsVdJR5uDpOpVO4jueTUqdyegzSJ0DhB5aNQAK9VojcNZe+I/7knAb
E7e2j3lpcQaekbfv8D0xg3MAuD/qrQVmddG2wzR3Gf1jO2ZI8qhAGWqRkaL1dXGQ
1n0GIHLl6N47S6OKKytfABkyX7bIiU7PImk0HmtxEuTYcaFyfiA/Bwii383kED79
gn+9n9Iuk1CFXz9DrIBi5hBoaaTdXfl7V5SCNmQqbq2yQL/f/43UBX90WzSQCx22
H4FuiQ1KOHPdNiSVyzUCRRdzmQqQjP8KV/+JJdiL3Cx2gPJt/RrjRp1n8gyyjfu/
08OzP2IQiwdHLQXaei1B5ozDEMOd6WDzrP3IUi35XJgQ2pyph7yAgkSmGsUN10Mt
MJp6XfFtW9ve2mhK1eDzSpUHo1D06I7mPBK3Ai2nWD7GUXkXcqUOi1Oe8LNwxdw8
NLfjzL5idXIYhtgt0+uvbBhUlfypIQ4uSFFNPK7CsDTI3zhQLRx7jPjRUQLEPjJX
7f9zNLsXwdwPZOGKgdp7GZtiWadxSdR+RuH6aYtVfQql+n5+gdS9MQ2dEaF5TCio
EftKW6m6obRkaQq8YGwZ3hNnIF0LzHqCJO0RVoeq9AOr6PmiSxc35F3XIR0xT82s
CG8ukpHt2aaTALbZoC3LrndKyK2R8D2I+XWOZeZ0l7G2mf12Gdb89ImeQb/NJ2Ck
QU0ByJV8wKTZCIXR7lK341kCBgkRF45p6xOnq9fxWuZZy6znlWfAVD7s4iEyua1E
LJyb9GpczBgXDxh66MIHEs2zTbO7I73+099VCf2I2+fZKj1Kh3C48t4MZlwRIobc
Cb5v3FAsWdHkgR09hziTE8dGtsE11rJj5WY/FOcV8FGr82585W5Sgqt4KY0MbY0u
kNcqzuaLWrgmjtx7ZZEtaNHlLVttC0YOrbS/wPZ+Ffm6OSHi3FiJxhHhOjSGDn0j
YSoyDJ6lXDTyJW6x+ocFwSmme/5xGZvgdFHOA2+qGRg27uqgE0DAJs6gbQ/Zqqqy
/Ev4SFg/3KWhrHc9KldPvvCBIPpxM0YtPz4KY2YyWs5wZ4g7YHSegWEp8rTKMSzR
UdFVX21lG5tikL/o+efS2jwDCNqcTAMHvTkAXnyQsjZDJFMHApRqS4pcrNwj1m2f
Aao4FwZudpZWROIXjg1fjyyjJMR9mOOAY+6NhAwsk4GZtA7zX0KFiMmK4cRQ17X8
wng7CGuE3w4Bt/gz8vngNB3Fbkcz1kCBb7l7hOY6WNRmk/pg+llpw7kMi6uDUuM1
sT/A0cE4An8U7Gewfq9/BI/5HuSLb1UHdzZlKHJSvoZZDRG0/QKjiRRyHtL7oCJQ
FOnQLEQVpnniuBPgagON/drtcUMGwXgcvuPn5cqi1VO9lqrRz6s+A37dDlvw1H+8
6c1iE/n187qX/0yEIEXL0yc/+TAhRxm6EZzantINhUDXye7uuL+kc4Mg25GQ08N0
rLQ4dBtM9Y/IscOlLITheQFMoF4PpCFCCECR1i+3nhXMgEy1gYHaL5hdvz+AX2xW
bU4O9vAp7VCGOSXige/aZrp40TkMnW1ytHtNPma17c2pGNoZiT/bxQEHuWF7+9tK
3cVpZb91iEpnl47dd2HIaXn+08vkDIQ90dzYtoILgJYndqKVR4Eo5pwa2kuPav0M
CT4PAnD9vW/P2zwR16tncgOsXPNZ7sptHDLVDms4BE7FepTcvNq8CpX1mznW9LTM
UWRWDFiBOghngcunagZgCG973xn/giA/deM0GlnnpDtdEdkb4h7Z6wBhXDaQnfXE
w0WjVs6QvADX7IC8F6YW9B9clC//NaxlywNcqKsqFr7Q1I/iB4L+DsV7cnCx3Z5F
rtc1gSAzYgIoymwoR/Be9TKHm6zmX0uCvdYDQM6xjpoAbdbDzDpZ3Iu/s3igtHfo
2EZ471gvOlEvhd1G2v/2kZlQPux866MgR3pB/pRaqvn9X/X+Jc5TOVOTgvy8BkfC
gZuaeS4Uz2kbMb+M/9PTr+642wn0BYsz98g6XjlPCbr1jHLFWlxsaMZEnWUKUHsb
V94txfhok2lV2Sc0pil+BJ4X3MvfQ5jXIZTuNCEYBApyFfiWCwyJrcsq2OnVXoM7
iMR04puFwcVi5Rmvsrvc+oHLsnFKBSO5CQmbrXK1Ahoi/T/TfjhrMOp+n0jwGOIo
QIoqIUNEiAXX7FeTTYIJg6B46ucjpyB5TolwOniuq7dOCjCSGCoI6sGP+WNWKFzj
eC364/l12/DdYp/+94wQuBF2kd/scbYaOoprmrvIzpIiPqTaNOG88gt3nv+Rlrio
AclYLT/ylxmYpx5+qK5AgJZBFt7ji0p8laAi+5cCfttZCdESENvZsmNmdxBWcbtT
tCNp8s0E6Rgu3slYcWCaK4i+IBa1buyK54nBHyvi/9ffURbPLNXb0GX2EsCjCxIF
k0bVKfbVHYz8NCw6UdMHswJcy4TILl3xKUC0ubkCjUgLwProIgvnasrOMuvUE+Xe
XAOZnrXLgVZmPxYiHXrJNiIcoyfXYzciBjLSGj/I6ZUdV5PGWLgrMtiFI4cWZ9Pp
JRwtTPtgq8rVlNvp78yGJIpDOh4j9nO4HHkyNnyhIVUM1aCCa16pjqrmiVUlIcOD
5iZucPENzu814OT1IAoBvtWMhNtgws+V9EnoKdn0ID+tsZHjugSVBNiv/ubFdnhZ
GbIlF3MA6/5JYTPp/Twww1kj2d7aXG5+KLdyurzYaQCf/72GotdvBVvXtUyvgE54
yq5zM6qUKQVs/TxVwYaUjSP/R7frfMkEknuIMBtNZp6/owHctrS5I+KIFEJQH+Vr
+t6kwVDFgA8SHuqyNoWz6xewJg60MQHFp2cwrjItUSsQakCc1bYjAqcDXJP8Gzm6
BcyXuHtYW1+qo/QDqFGgqsbnPbjBrJuCw5aB/tMw5W1NjLLvQrwnjqCUUSIy94S3
4divYBS0Xid29/4uaql8D0Q2xsNQl+4Ce9uGbxo9lMu/yOlJma3nCqzVyROvI7c1
X2RFrV8aFUw2dNabWD3GaufK8vqciy4cy2kjgOwvPBrLChmBSPdq6BPml4koySJl
7hYqOMsWt20+1egG/nWmlgw+aXzBEft5zWLbamgCqTUoDB5GS1Ff967fFADCbdsv
f9g7VTrkrWmSvevim8DH40nVYnVZT9T9kTFALyf+1zeVYbfajeLDnUPJI+9fQ0GD
piRAMomuvD7rv6CCKel1CfwVDzvOBnjsKvutmcjS7+GXLhdyj5WP/i1mMbf+z+BG
OquLPY0rQR9/N7pIrRNaXfKZ90gy/CcK1rbX+zG9fNL51jtQtyzoDTDznxC0b1B2
qAhtVegkXo1oO6/oi7WPpMsWYMM3Vyo1Ww4RLnH6e2b1bBUFLI3UTpSdheaQXpHh
S27SUdox5PxYfeEFdeHTifk4FlvXnd31pY5+04GyeFEFDS4m/pE6uEGEKFDPTqHr
JkQAIB7p3oXlD7GfWtA3CB/CH0wwmYoTJId22zhfrlbOvR18zRsHz2Zbf6Wkp5AP
/h/jqXyQvlCPM3ZVy6gOG1ijf6SsaSuMqZHuQGZduyj5cQTBjlpc7eiefWaoQSPW
WkTpH040r/27u7pEDr8dqELP3wrCamdChhu1uGM95MMgHGHG7O9339VT/BUgG5zd
zONulk4NKFDAashQE6bhMK5thVclbR6vMqTjJybPwoyErj2OKMOeUUWPz+mLpVK0
U938ES8KINtg9HCSS7RLUaVwUHiX7T6MNVWA6o7HIEPBna+LbVSWKnvyn+pRuC+o
AOXrBGvTaBEcDfBsZKUr9wHrVBVaSaWVyWkC8ffJGrdcLI05BnPMQwiRJpPzrgab
SqJUujmSgg4lNmyMcJYh3EiKoPm9Hs1KasLwPKKILjFRNd+4wrdcXBtoIG9r1JIR
/nLKGgj8BpIi/23DUJ9ukXIGsk7uPkYzNIUknfdfJsOQtm9qV1/B9p1M+VW+C8QQ
3jCDynzufbDka789SdJ26ZOMUAGM6y5yMOpjqhS6M4YCN0b2Rjp9dKRb8+2G1ixv
B7SLu15TmSXJfqEK8/pJCGfg1Q16Uk5t3dxUIvmqvDfj3bwgDZwkY3ugMJ4g1UDE
hIbYHgYnayjeW+q11bhl0KENnNuz5AFsZSqZKoQZclpjhmswxfaLnv0A29ui5IBi
b099jgng8pioNdOiZM+C9qXSwChUUzhNSf4mvPGQp5+Hj36gfBAf+cpp1XKYMwMU
8rHiIrzCC2eybJX5pJh9ROQmqK2ov2gxv3eWNsrL7tpIMYWTfEGvQ13+pydTSPVq
mL/fxF9lX3YlZQv5kaf7fH5D+vKrq/ZfX4phstTWyOBUfw2aijBeZeMzGhPQ8ZIz
U+00HA3GlctQA7gpOeYo4TqEPidYMGn6rUYbQjJ8lZnvTew9tLNtFmDaoqCglqIn
XBt/bVWcxRVI6tocWeGkWYi8A2T3c9iJQ2MnrRRFrTolxKt3zZMDjhpGD5EjImTL
dtk/CWJ79o0UNUDMFf8yjagwcwmdmaIqAHuFlVfN3vC5UcYidoVWJ2K+Ah1bzB2r
dBf9RBzLIqW+sqWXRhn1lrsYFfAUfS36syBOcRJf/1pizkT7Zk+EekesNdrO4mMT
m6k1eMzIkw64IV5KICYzVAmsKdetR4a2Fivky+zwgSyyaLvFoshEdGMUH4/vdmHo
3cWqpsKqAMKSsUmFrR1fCNsfZjPHYT1wdSzPpgcdYDkJV7RVA9xYiqzKlLMWXYfY
ptJEDORMv3pkOxgRY88HoIkmX9DaqnABMzd92MBwBVHI77zb1PxIOhdDpvbFSSwG
W55ir0TRnDhNsdXIQmQgHX0G1SdPPnxpe8OLvmQRT7uktS100g0Ic2LdUcyBr+Y2
qW84ieKno3TKwJo0k95M+ZIxFHdIVKiZrxMkm1hQ0JlSesWLnnQegxLfcXgcIKIc
ZhEYKIa3eh/5DHiWqaRGpkr58JWBxJsMPlwtpkGu0A9QGbQIA2Px/P6BzejfKIl9
yJd3Yz6mHx6S0x8b/HL8QuJt8vr7qsE66gz3qzJ3PjZlcI5LxHFfUgemvtfRFjPT
bRlRaYDC7IUYhwRSoMiqQ2f0ot3PHDCCdiqfCDnWLkFiD6r4EgVgdxTYywf8Y9Bn
++PJs+Fu89H8sUgO+olh0U0x7/AggtyrRuc3xDwtdUw3RkOuErWuPUGWKj9l28u4
gLnKCvg2dAu7XsyOmHK9OgBp6rlid4SfQqfFJffy5cydODct5R/smog7qV6zhj79
KgjyB28Ehm+8nX0tzVk+1hqMOB36iy3ixgUsJsSp0tvnaG85/LHSX1ZhjPbb6JMJ
t8qH+Uw/Q899d6oC482ScvDD7pIbmSgAo1hOUkT1Z99ZCBjSePn2CNt64pZODTSs
kAcafreBUab7hVCQbQ0T1gy8GTu3e3ED86OKgX9FvVa82NMscQZU/iEUgmx9zJdt
/v+0c5dw7R3z0NgpKX+pBC3hRZjK6d/UW+IYiA5vUdyVF6IXaG1S34UYuppPhGKd
9v00WBczi3cZMrS4G8UHsyidvprm1CTrMAo/3cZe2dGRFWYwDBbpv7ONFN8bQZY7
DQiNak/PNI69ki3W5kf1fD8zv6QFN3USLh3oJQgCab+qHsCCaYsfOI/iuVKPBo5S
Son+Z5NFQ6UZtAtWozgpNdTAcZyDUSEWkvizz6jf75mO0Oly9YBeGeo+LqsBLNKZ
jFqMYG5V4bMc6dRfSTeGntgkc0EeLvwwnuBz0fjfC32/vsodN86qzmhGqYOq/75S
X5bl/2pHqtfUndIczXuH9cFCmypwTB2JI3PkG8j/jklQSZgdPUWl5No0w4jRGGuH
doiuA8NAXw4Hlbs6nQlHKsP2Va4orSBxNXGK4MwoghMtrH1adpkwi1Rv/Ei/jDwK
xnEu1Qd1al260DDnjJUkUQaWztqo1hSV2X0vZc4oSSnLueI79kmFrAlRt1ZaS1gU
Iprc/06n6fZlXCx5U1EWNAm7tmeHBtU/FYLeIwOA2euNg3vRYQzHyEcI56qPDaPm
Ny9L9DtOacYf+5XmRPj1JHz3n7BRbOJ7Y5ww8SiMatIWlstzmQY8N4xL/4D7JFYc
pG9nq9uG0NVG4miF2Fdl6pbCbfHSIzFSs59rsBBx6TY4tMySnG17wntSScHBXPnS
M1bJaqBsHBbhUulvDJ/jx7KPKnNyzJ9rZW9nRF0PjnSC+aS0e9knEIAvgml0tNfz
Kiju8zUhJ1Jukh1BlB3BhMy7PRWBb333rler6Z3bhDf4CHCOmRsKwjHlKSuRJxx2
mlckhL2152JmxAblxLjpOoBj957ORTWQEzzkTZn2jpGFZyz8QE+fA86ePY1hu8SM
nCOlsBoygHJPG2vjV0+vb+V4Mt2TGKEZN9/gDUvwJwPSvkTLbNGg+AjncP1J5GFn
Rkditn4oqPw9SyGFsvR4YrRswwcl2Sx0yjnCiHAHhV/zNPWvnTvoizYLVk/5GAhp
vsh1y/JtuHtYN8llv8o8MOQdeemy0/fXTJHEX9c0Sh7E9jOtKvUlN1bRyPdmzb2l
wKXH0W0SUXwqmsmhG3xZ78sPluMJN/KBEPceAvrjzLnAAZDZuuB6v+wTXTvYVBDp
K2ApMSglm2GKIbrywEipXoEd5S5CDDGC+U2BEVqMbErLu56YPhueujneqkQjs7zI
DLSr5klVtq42EPW77KV3yU5onrHbvCuw70liTCZMSDC5gzWFQ1qgJnJ0qy4COoQi
1jfxR16fQ51at390tekT7944wfhz0FDc66L9SjZa9q2OsAx0l06PWH7jd+HVE3e5
zo4mKNSkH6+gcGdzB75Yir+DElxsHq1N6NTqCWmi2wy6YrBeXXshRMmUCwSiugWR
trvnOCDWyRP9QCSMhnazgJi6IA8HEYkTXrOt31J3h06VthBAFGGZ++fggY2UKenx
zO3qmup+Sz0n9InATD6ZGzDMOCHHPeo7xjJh26Q7p9pt8C2VAd/QQV62W7ERkfV+
KexRUiL0jrusvSJ1+XfAghn/bzNz/nFtTpdMb0BLEAmgYnHEn2YrJ67fagUtYDqE
ZlVWO7YxHQucelkBhmafJUB6bEACeXsIbQzqTmYA9kMCFF5zRU7TfYUwC79MlSpe
whpQMzdztBFAVRsjguVZfFwgfWadQsR+6S0U5Z/MVx1nOO/AH4MkqOD17aPg7cSc
czePk3vJ+JkxOyPR4lQodoxnt7K57Sa5h2qQUfEo59AcPJOslCx+iVOYQmmvoVuv
oyZcTpcAhwFEWICQCq5pGeYQVikwxZlREr71VR28TdlsKfqrAlozgcQWHEhxw+O9
AcTyrdLsESjYVI16bWoQVCKjQCP5VxAYjVs4m8wQexsD6qhyP7XF/iJgT3UwIxd0
ChOYdouH5R+kkrKPVMPJNgEkl3DFCVNmXp08kKtWLN55iqWs3G85crSFTSPXfgXu
nxw4YaYslf7aor2iy3uE7116ddNEHgP/6XuiuRq1ylu1ieBo45kl0HxXDfljsAAT
SFXiztRd0AyDWtyY441ko3IpMG1R+AlrcsHM01AkhFwDMNhFunzbierO+CeuFAqj
G1fNoql4W+Ew5iFmElDLIqZwu+LrKcr0Pv1x0sxR6KVqd2AwyCIop+Gv9xEF4KTU
ZfnBknwBb3O8xMPjq5y0bbt1Qto8ehqRxUKo8b9jhJKOHF9+IgBsgHgWj6tm0L4D
9HPmVwBMUTZtrkWL76FeIC/JzDprklsQiHQzaLTiGR2OZx3LUExJNu19L2u64yNB
CAC9wo5C1N5JmGy1LGa3E9GOooPP+z1pQgu9mwBpTbVKm54d+uTp2w2+sJeP8801
ZSYMNCUtZkBpRn5ujNyRLIS9oOeFcRIB69WFpSQ31b8JTCjdAyXY+yk6QEZDSVQO
1DF7nxA7D496x1yEcQQKs4xsxzzoX23S/O1O0jhGX1xxacAclMS2+Spc2xQ6ar20
6KZmfk4atkguFuqUtCMESqbIt5b8h+tjZu0N1us04/Ts15C/5XQ8yIDgHqtv+jHd
Js4MeURbK4JVK1Z6img0x50JdEgu6S8Mrdcw0Z8Uh6XQszwSfaOx1ELQpCj1GS6W
kfbeuKvht/vQ2oCxNtUWUd5FeD5CcX2nhcXqZMW0I4/mHzqJzJ4NUBb7T/OI/CTC
YUjlGEp+Rj/w1hmSFKG4BhzDUM7CsQOPCqLRjpxQZYZPm5by1QlqSm23Tvehb9RB
KUoCXLsPuH+f1emlupITZKSCNFF7tyh0pv0DHrlnFQtEDSX6lqJ5LCho9Q5un60+
r5OmnarRTYhuGSbnmR6D2+Jc7DZqpjelCwwCCXleEQ+Yeo+qX0vGObmpVMUE5NJ/
8Wbl7ZCbx/z+kSlZiBRIy3ZMBYiOJXl3PVRS3vRiYqEthC4nsEmuHPDU+cOJYFnq
RC0CQglpw8XxU54CBtKhD9xkC1KViiF9K6af6A98PModKO+rcFJzKkYZ7V1za/EZ
C+2e5mxr3W6wzZPfE0IODDka1AZ0edd+B+VEm6NroNlivdgYiAVUN+uwmGjXK04v
9hXH3yQJ0flLT06FKB5e7XTnApL+RnqHsF2X1p7F/GPzBJpSalPQyGkErcwOeZZb
hg5pXfNVt3qJDk4FuAbDh9DCwOg+Wca8jzXfOE32RtzizR1UCfDXsRjOV44w2hvp
OOycDQXik78B1ReoSDsk00vaxAoiWuf8olnLftV3sLnMUn6QzdL5or27SjNCrXWE
qwgeV0FSkqBRVvQPgcTw2uVoyMBXyqLdk+/1gYzOP1Pw6CjUopQsRwxZ2FMaxPbz
vbmDsPCJLeefocy8a/Uk3Xano65b2Ja+3VFvnAgA9Ktwb4tet3mh+IJYD9XCjO66
nveKMfGmwLRYnZp16aDjiP0yzVLylXZ/bwtX2Wb9hRkitdxCNs7XranWOzH4s9WK
M3XHaI95TgcD5qRTF9W7A/4NiBqU7a6DKIWdHZNC61BWScZ6zQRntT0E7IMJNDas
ljeKfPRr2r0MqNrRN69e045yC4aSXXZaQm8DqQrk3hiOqWOji3oGz9rUmtMXyN5C
6iDtr0LTgp+56rwfbkkTl64l92+vrrZ7fTWm7+jRjx48SdbCkyJeRGtV22PH3JPZ
updZevsNV6qtYfZUUwDJxN2Hf0ZuWZhwEtwgYuVm4/TEf+CJoThw8IANT8/rBumu
rJFK4iO3a4xlb/gbxuVxbZj0hq89/5Tm9HH6EjnASrP4PuMPxwo/qRHFo/pUDuYh
m8zw3V6DFoW6eV9lt75Or5srkd5zRrCgJbhybJ4fz2DTHFqgI/MaZFsZFYWJOEyj
iFuTIlMdK1v3pC9F0tbT/6XzQV/bn5jkC4VjzM+wpHj+yZYSCKFSGjzk1daLI1rG
4KwRFmUtoV+7oYcJt/Y96ruEg0YWLnTRxb2VEtOYtWgAvMAwhtM5nBFnblh913ym
H1rakaFL6zZ7XLsPMOabRMg/Q+d2NZOzmyxnHKMuecqvjD8bix0izP+Iv95zQgN3
MgKvDkDy7nXCjLnUmOvAMHUAY2nAwiTZR6BUuW0aYXMk+9w53f6sk6tApy9vqxV/
zg5W/yYd2r8LkjSsXINlCDiaDA5jnNIOSMrwSwZmXqXm5yc/hn9m//Zzu8i1hmeU
B3wmRdhCEmB+/ItxGeQfwK0owpCA8otPxfHZVRdSrN5kDGtnab6mDc6bPwSVLGar
yx09fF0E1DZlpDnGnsEeRSdqKSvJrYhFPvMBMQUxpLlO7hXbt9UD8gaPa4oRNahV
c82kKhPzqPYuSxnaLPuiU1eVf8oFyijbrZQkobBo6JCI/xmW7C7QcWeA2GstpOwb
qHwx2nOPxRwcNP3vJ2Yl56toe7Qykt2DlL4OkZUbd2LiejgTDUlT1LTaV/5oXMFK
odvyhM0SJW/+FjH7Z/QUYX1731GaA2a7tp/xbzxj1kL2fMf+VOdJNDVV1s9erEkP
ZcHryyDMwFNxtlFWKmV5dXu0KuZbvnViYwijrx3rt7Ck4qWigBANRZLUvj4Cbp8j
U8KeE87NI1JSYLCp13MZlCK8JlrhxobnNdGB08v4jCbh5dF7UaQxwMBxEyhbvTCu
zuOb/iiDHapocIvBuOj04VQe0hdEWqFhsKEOoYLLpp9cpLtFtb5j7Qzm9W8ZSU4E
p1asfmAtuxSl4N0K1I2p5UuicU/zySCkcce2wvwHsH7wmdX6UKS/gEoj4cpEiIOe
FYuD9m4iIkamC/iAVEgd5wnfMpafljFn6Khvei1o2elHvtaS5V7rVj28BOiYRHOg
B6z78V/+2MuHZNAc65aPhhRZDiRFs4kPFTB6A1qMyRCAJAxiHMgPS7eFxmdxYP5H
nNntxjCLHsF8iesU3/amfxp3IZt9IzlPzCY6EUyZibj9b5vKr8AXyQQEFH4hIQVj
uCKSRajgOo6IYch4OEbieN/1bfwbOEx6uNCAWKlE+LFOMCOBSba1kIhhKS4ysvqh
3WYlY0ZtAA7JSfn2ldeNyRrm/MF2/JH2kQpAqEWuOwP0ZZSMFiSKz93bU5yznT3B
X7Mn2xZiyJTVbb6SPcV/G9a2xaz0FcM5wlUqwTtQx1FNYUJBmQ10bABm3neBnCas
ffH7tUvaOkUvNI34Hq23WwiSELhdG8aOXD8kommI95B4wVUnRvoPJ3w/N1pi6g/b
yVU98xohjC5YFM90AGEWdPPhmU0sneiRoc5sxLeFznUJzHIhP5plT0qySZB51h5d
Zm/7LBQfnuinUlL6qDTzm8jF34SOmUB2NptZiFHD9sm5HPD1p3QAw5A3tYLeIwlW
JZxbmTr/qSHJglnpBQqwhDG03wOO2X1FGVH9m2yHfci+FwTCR3S1Zt8FPngteMPM
RjyvQb65VpVZj7s+r4YsWwWaawIGJc/9IdpWQU84XStXEbjl88bTBAe5ccGDMjzy
57IwE2C4T18tfeDaeI2XNrUiAeEVFiYcQ1Q32Y53GpZll1BYH9xc7BPBKQ+sL5ix
WTsbyMtgsAgAb82c+7YzXWGfIoOctAUlL/jpTkUeS/55MQngJVNezAsCDJKzpPy7
0DSSiENJI4Ww7egvWX6EJBRSJ3+2jlBP/7x2Fh5Qh1SmFdwiN1z9403rmrQoWfel
fkbLrcG5mC/G1nUqr8msX4iIhhzrMF0hECrscac7Mm/QHkTPvjEwNy6twprJPS8G
6i3ZAAphw/fA2t9caTKGKbcMdhzczopnYElNFAzyHCBpy5WndeeRIwGFCx1zPKa+
YFj5+trqmCg7x9FqXQiL1eSF7qxKpEgfS1cfwhMNV9AAJ4TTZovH2fdCdnNNXaOf
aMmX8+qQmtzzQgHcNg31MTY57nsgYqnClmT6SFrRo7Q/rGkDS0JqMk+7XpZ4eVz4
vf98yiObSW6UKYoH9e7NrjVEBD0WTyvPVsxtUSAsqDeK8ucC+TXD/RhrDwbWMpnc
/2bHU2Zn0FysXdkJA3BLz/jjT6gC6rNpNioHJ2oe/hojA+a1HpbD22+OESMyyUiz
zBfsJuHup5gGjPKG6vAFP6rfo2Zc82k6k7RU+zvEFYdP8+naBU/nXFMkpBnNiQni
Fdp5fIpgKyTWdEN2SWcKfTvSDSOf3hSPCNaZTLmgXVRIQmeSFN+dVk10jEry1sCO
1V7uWISitmERmk48GdQzENb+5eflULUJSbPAalJRaVsHJxfL+cYxK0CSS16o4LPm
qXXvSsnbHj1cAXV31/jMB/4NAx1Z51S8i8QyMR2iFOT69RUDisn4vbcnUeFSFuDt
NDK3x5dAV57Y7cOsbLb8jd3FqEz0kLnWlvAYcsmhfzW83kdNw4sMB54p0hFTf8xT
x7+b7xt2KqkVdUQw5mgQpjoyBcmUWzOxYACmSphM9zL3Y5sw4s2DLFWfU4ZjP3GU
Ia5SerqxTym92MDLvIBXvGUju8cSmNvzWK+2gLiBpIUHV1j5iwRA0UtswKgTK5hJ
ZdEBhJgluYZwefJf62hbhBndg/0LqVfxFckLu4ZZFbtN0KfX2WlAqWw8pvWRkp9x
zZa8RoKwq2rW0hIzIfLDRRamvTK9r5vpJNEGCcl02w+s/zkEU6RfQ3UrKeKn3YKg
fPHQf+WccxdIq729p/DPXBEfaE/FRtD/cQ3iWk6poWpDH1CUehktsPo9JyTiyWJr
bl0GBseIHVYYscugFbE3ydPTqJczb8Q4joeOjVrJ0DAOMVbRMs3q9uvHkRuMiGuV
dMoKN76ZCOimV4Ufk6O/beYjWsPcRtINemSswSO4V/ufGJXKIXwaW14NbjEbvDlj
OwVGvz2ilg2eTp6N59+2/y6e79knKgoC6TY+OYPCD3NVk3fSxD/tPU+44NrCjye5
uKyh4pEedfeS2k7mTwzOSK2X9blXIfzUbYrsR74OLL3y5Hq21NnYX0f5PtkLeMtA
H2tx1B3YGlox222DI6ZW/EU96tIkih25MHCrMPizB1yUrVXOGv5HflZMWQRoB+GY
U709kJTiiEGX8w5E7ibbqFq7i4f6tds4mtzx1KFZpkLyUKr+VCzKPB+XBCiIf14V
QellBViC1rfQ2U5OxOJbJ+12i9OmZ7jhHkne4KBYycIZ73nFmzNPyHdIlyEiwhNR
a8HyJHzM67dUo8Xhp6LaXL1gnumLUSHtZGEoyi+bHKOtWEBbiMiR28S82+vvr2SC
cjUxZll4XUJkT5qzB7v/YCtwAk21SCiGb+17vA4TqyMJGMFe5B42t9DTNVj8MQ49
JD3WIhWrw8QyCIUKhZgjMuecSgeBvsYc818KxUzG5VkoKjYoOwQjesEBlIhFuBwE
wL0wcrbO13SvQIQvkEoy+yRN2vb3hZ2um/WUdLFJQ8rOTuBl4pfarOAJd6XNfj6V
uZHnWVdLwOsnaflpphkZpvKkmx+Sa1a7BkrkIJ7gmpvtE74PkUty6DGfbpbNmnDD
9RYkP8LrKovHuNHivDKAEb/kcU6vRO21Qg6oWCQeZYU4138H03ri9QxDq8tFQf0u
BvlZzD5HUhmGAKDTT/i3UdF7iwipilLh42fy2jzEZzNPDSzh9lA4tt5tE/aHA+7/
solgY0CRm/F5o6BymDvI2I9oNQNpnzdYacHsJn9IAoK+jddEI745HAx+JWglLrgL
iX4p//ORsPW3DanPPNv4hpMxT3fBSNjLjddt1JaEe5QInRjSzpvymdrBMlw8ejCW
qsNa5NXzciM359x6jN5ooKw+5fLa2e0XXvX0h7r3G2BgGc1V9fzWBEJawodsf7L9
Ac/lya5lGuQqcqfbATix3NgDEIAciZxz/UHz87xMYgJTDwnYbF4fyw+aPTtHM2Rl
ECF4wl3oQv6UzPrYeBoPKOkppJYVNC61flQC3v0xbXeVUtU+wyt87YTs9H3zyKi2
y9cgs2Dln/FYiDhKtDnFfkFsxnukGpS8fOpwnrJvxRiEznPVsLLlIFp06WYBBliz
O/UU+OtiH6UW96ZR4myxMNMjFo3P8ytpZwlIi9FFEtHo2JKs49Wohw1RqzxV5FSg
AOl5OleRZE7Vk7FTWxp+/SNz/O7MLcD1j0tvnAmHYPMDNeTVUhAVuL8a3xuT3wIR
1P8M4Qfshae8fzHgAcoT9S6T/1TgvU4phuXJrtsC3On2TvxNdFxqj/0jLGxUc3AB
1DZBtzXpOYIrO8ep/PY6YdQ5A5u6kEV0+Ds5YLtsPgIiSlz7Ru+IrUtEluye/O4L
TNeX8M6eZGrMyNtwg59ME4o7VCpB37k01q5xcAseg2obawz7nZJaYgRvd3rukliF
6+U1jqeppMWgzzsovvAz4w2cgNIMIpZ+1tkqXvcS6eTlNAJpqfG568P4jRjhzUu9
e0N3RuBa28sufNGV7y82u8bxSbefkeZFNcZRGpYPCzFzoP9RQp8cTmJ3rvodu9Jq
AAcFFI1mIXYJdWA8F0ivbnkofUbdsWNpwJ6c1/B0GKeUAHQbit+xkeyq7IWTPMfQ
hus8gxXOcFxRDE8UgBqLu8hb2tN2xnzV4t42PEuKhiyMXD2bh1sfb1CqSqG0sk4i
6ny074VhASOORl4c0Blottie5JweCHJaTQHklmdNYgyTyFt/pt2efhk/2q3UwkUs
jo5ZZYavKmAyINU3s8qZi7k1gSTbvTdEjiicsfkYUUAd4+exSSmu9f/CWJEATh6S
ZXhFKkIL+1uLZ0uLxhvxAtOBRAWdJ3FD6n3XwfARUsMiF0liduhW9jA10fruGEhY
HGLuGcNZLZRFKho0/fsvTmStH5Rkj69Dwi2mYzezMmkw1UOSCujoJI2bfCupxILM
4ZSpgGn8AKWGCmUYTf+FSDuH/BciWrOoqaPA+Aa0QSyIXqEDs4H+vFA4+GazYmvq
YkWSUHZ5KrshWLz1d7YmerD7L1sZeDuJRnFYelg1pTx92TP+P2YPhYIIoQFE0KNe
YyfjQw9S3OoJxlXC+vyqbNVzw+mEHCueT/1NjAKdNmfS5yMD4U1GvmUCdiHFJy1a
TIx84nkkjlVDS74Onoibw0K+VoODfV9B1NZOmVu7yfAB8g1+l9LEA2Wnq6YnA2Ua
WHebvQkM1N0dUmsxn78zEazj9zw93wG3xQyBV+z/kdLCBbNS134ybnAXpJXLhQuH
nm64h4rp9t/q9r4WLAckCCo1GpLkPQ9ksyywOO+GMVs8o2EWi2MLZ98b0d/HA2kX
khbrsevybQb2MecN1PUMqQzVHH++tkV4Zq8sGW8uNqIo32B+xIOPyQgMrkNhVumc
TYKjFdh7Rg1orpvNrym5v1I1QmBQPLRd0tGtUOZiXJdE5gxT9NXEN/1umLYfsGpp
7gIaON1Jtv8/vQ59H+X1XHVOib9D0NaUQLHRe6YF3QCR6muKgKOKp5MZW49uZmcP
fXcTu3iluX/VaDgS5TlOAnrVaQsJ7C37Hhk1ndeMU5ekwl4HbA3CGLQqqEBbT1OY
+UBMHxyIO4MWo69WOoAggzRWVGlHvUG9GpwuQVclwsJKiCWLNGgphJeLZvsOA61Y
ePNQeyHPhc+hzol0B1RPUyH5MidN7Ytpn3SDekYRIwoIXEWzqSwUYB1xeKdtxHWA
EuuXTDOWz4V1htYTeU3Os77Hn903TxI82Z+xCMplMv6EnnBSfGJkFqNUagWxjw3u
J2X0RcqLjqDbCleKZ+1qQqqanzSlLgCV6nu7tOlfw3jCdvhnjiXSAX+jpPvK84AL
fxE0rTvwvXGsbqUmQgyskNCpj32FUmnSYgamvLmCLLWygpYFgiEn6bzpYkh0gbXt
KllhdBnPlad3CWB8U2l8BLKpN/4KWHbT253evZX6HwSyPx1fS5G8z2nhKRi+px4C
0uxDK/t/IcMCYkoB3B+DccAl2a2dARYNK/FJAYzmTLbE7mHdpOzrhYiEDhuTw5vH
NikazjBchhjcDiVrC6R4MHvp6puvYecF2Aq2Y7ozuCG7z/sphD0dgqKmzdrRfIVF
LI4yANiqOdKHaR0SqTOQlJnCnAAqAAfCdCtoN6Ry+WyNLEuvrQPivY6Y0HiCWCaw
fHqDAYGez3pT12ZrxLSXb0Ao+5T7CSPnjuBoWulKL70xBdGhtv4m7O7G5uF9FzQI
uDEQtMEi6uqN6GW5ur/La8aDRk+7MXlydrv5n+F8FVOgoLX4wMOjgi12dpWHGQl1
OglkWNdoKoTlLWobvzEk5dRbNiqcTqD7N9P165q5yZ2tRybWAEKT7ug4gCa2rEzZ
JeucrMV5RGLKD4A8SojIRFY7PyADTZ/16UpGfXipddpjNFFYI+bzoJw5RqImStVy
CLIn6qoZdnZ5Yo06GK1X0Yx51RgFHv8ovPg9LoRyil/4cNTmFqwCV+etetPuJac1
FaUhboSVOi/McolBA84jPggfPFe52rlUCH7G4bQkLbN3bSnJ2pQGv4a6wRVvGprH
Ev3oGTefdqPwm4EemLYpWaWFr6pjrGbnRwansIBGGhpFyKB02Q+LYmsUIPU42Siz
s4KshvresSof3RuUjcCBUVVmmxjjcsDOdqH6JMe9YVqqYFSgHkl71FzcdKAFSnEh
3Tqq0BuiSZwKJGy5EFRetut6tVAenZCiy7ciwFmzApNSkNV7NfQS0qYUcl2U+a4c
1azqJ09Ica7GvCFUm6jxDs6LFE99nGIH7m/PPyQt4g8aVo/dDN6diLGDD5Ee03w0
j61LryraRqiC+QsS054AHyI8dUny9Pwitt7aNRovud6pCoJ5iYNvlBvaDmw3y9bp
atYWfpyuWEZEtXpBSvIRRkF1xXoYAaOVQLYr7uzD/TeS09psKlredr9KeelvVuxs
VRtQr6lLf1pDDwBUuq9k/OITbg+W6xN1zy3jfY6wnDgY76yVtan31yPxyL6Gt3+K
u39HE6BkfcvmdHxk/i47RZfCRrRL4HfYByfStz89VWlw9Yj2aWuPhXnmPODV+Xw9
KLwWo1fnp6qxYrxsxx9CLG51GT/WPWAvox748AHnYXjTcBmAQ06OFXB8HPW0Gewe
/Oe0s5Z/krEiFzgNEBM8OyBFTKF/7cODihScmnT6SO9h2l7UQJpNk/CZIXnC/fm2
73evxKssE9OBAZsy4O4DBkS7RcWxHnCa1I02DZg7Tv8RRDU/giA71uLo9k2pzMk5
wi5c8tGS8XFdqStWhKPA68O5fp+/oWej0tRNHPBrRA0Pr1RlcPhRAxkdK1CcAHjZ
TuKmZ3rFG6zMuDomDOS9AlbbDJw8b7VQWF/JFTxJJHs2aYse2pjrJzJO/Ecdo3CZ
/LSgLQOVDvxCzKvhT512vCKH2IGtlmry/OROIigH94tXzEqU+GKvc+9HzPqm1+i8
hGWsXPyVwKFhbYtnfa30GB7BRz7luHF9ikqWhsfASAPiq5X79PDCBE8Isu8rvGv5
QJr/0NBgHM2jFJbrxVfwFaVXEGfNlgV0MZGa4lupYJ/LVNVMSiT6umXzvvuzzl8A
WrBw/LSrJ2ylRcRhdi5kQV9V/pMVvbLw1viHjcuOACUea9SWQYGnMH5Z7NTrjeOE
qj4/4H2Ilecw6O3FSqWDRkbIe013b4jOazlEmz+jGCq+rzak1K6Q51PLDWM/RPev
tPpEOCNj1aANVq0amI6PSbiqEMdjnmLuo73UeVhayWDzK9teWBssf1wUD0hYamId
l2qFPdWK/5GsrfTKVaCyzL4fXgSc+mJHAMSbTUyGc0l3IDr5rOoC7DJsTvJq9Pe3
AizL+N5+F3iue2m9oR0J6KU6MF+9FW7DOiRyaCt2vsToTRYZ0Fby1PAyVSwqyEqp
kV/cb05zLr3CuF6K61pzCqZn0xuBOcLA3Da7n9q+laXu7ffVtZhcvBhvxAIAdrBh
dluXcTwYCr29t1V5u9i71fnLah4XlntAsPQhgPJZWozwS2SsSDgUQb+XzgvSoXlq
ZYr/iHkE1DIBPpNIEudBoZKdIh97qoGi4GCxtSQz5DmdqfZhsLYzD9Dac/90yB5a
Iy+ROKvzEBSumYhCNJsrk1Dcr9HHwJY3bucD6rZL8wiaGaJ6PYQOl0/wU5QrRi0N
Jz0HNUdrlwPxmindjZ4tSOUWgPZQuTBakupXaFB6ZI2uLJVKtTddWJmZRxmQVmRR
nvtstJN2oOkgzHikAPAeAjUSoFjJaNrhkzRSHSJSta41dZLvHbYMdnK+u2bvln5w
re2+Eue/LgX4pTHcVEbBg9l3l+gIwdiRWlMQM3ssynfLwTqiid+HVzxXJDVDJtXR
w/M0QuXcnUK/7Ub2A9Eojuk6+wtxJF3fEGTnU2n9HAqmJ0E23t2HVc70w9+LnaC9
Cm1iE+BgeQZCbyX1cWfv61DWWR2t/GcdZP62jNRce5tstFpHyceK8dqhxzjh2gT/
rmTE6P4UjjtA0ayATBQX58ieBkm+HGpND27XKIqMSxZRFNLPv8ql8Yp/ITT5SDyN
Q5NpN7SDquQF/+gZHSfdSYRRHeIWcbQeNTon9NHiitrxdiXTqXjsm1KOWxIu/ajz
2fBrAbwZ4xlwxjM3NS8PuQ2ox+t0IBixjxjH3rBApg5M81r8XGdDYXKWTiPk0dUK
+P+KJXNYjmS9IcK//DFpzgSrc3FFCEAO/9KPFy2aMayMDRmSDUs8itzDbl685XY8
aJ0fKbwbn1MAztCc1dcOkzTae6b9tqJZbjv/QsRL6yDmiU8YPo1nSDWr1yth65FJ
vizWI+KcSmx+l4QU+9dQPHbsFuOQzo0/Gj1d8hluiaEYGw5BvLDD+00rR3p1TPZv
D4rKRSswQttEevWlqwC0RvunGvEtKjyrkvHGzZ5aUnKAlpx8hvpi3Nw1ypn0Pnte
LRmJWQ9qnZ501pPyJyWKJWlBjKs9Nbc6MW93G+6ausEcVpNI1vn12KI2xPSYpTEU
cTPPO14D3rRcr7qCTNJEV6u/zmzBivCpa2pZAwyP5Mc2X50IsoG8PrHiSxkLfB18
CQEYtTdXJp//saibwDWS0bT8m03ObVOAIF36+6bqj0ImmyhCnsac3stAwS84zhaw
53OJorBMZCZk2elt1y6ddI1tcdYK0eMIijjVAcJ+ZFUH+7KiQZ/UCEkB3gnPFarT
F+dCQ4KWdiPl2V5l5qmSYmfpgVyPohnanrbyNOhVr3WLNc1lzD8TGxbh6r+EODQf
tyRTd4tfpKh30w+GxWiaO82SJFcL2ZUPHt6Dk5gNMb0usmr2TOY/bNXERAjd+P7u
rAhG3RA7iuZcxVEk+gd5DkKBhXahA3OKTcdUr9j++yEiwUqp9//HGPUhKL95aRRv
Jv6fC47ZNfJ/s0ZdLbtJwNEbkXAjL29n3nthswfBYsyhPny2nmSwYND6rnxA5df8
vRMTrFtNQr7ZuCJ0EMDoJfrdWQfuLyLM5c8997LPjirVMp/rqkM185O8+ZQehfrR
kUc6uI9r+MeINFVbfGrACUY6v8ZMI+qbqlHJKnRF3jnonEOTjdzHnyWR+T5jQv0B
h66eZGIR4bPgoPil06VgaTpbQWiOxt5mePfN++k7lhGdmdYzMix2QwLt1r15b7vL
CJ4GE9aTnUUH7/+jgPbM4GJxLhilfGI0VeOlRv8Pe0pjuUcX5yYXw/ObA0TkXNEF
jGWQVEqqlepwXYNZHNgQnpIjksFWChKuZkwsWSOhpQeHk+hx+WPl6JujRkNwQsxz
J6OEZ8IOI6HxD6lcj3EhYfJl13yyhuoIL1lRIEI+5DLkYGmLl2vy+3xI5VIAWSrX
bcLGJJIbKw4TPVFAzAp5eKRHgVAKqEotZowMFl0bP8HZXvoZcENaqRE24cKRmBq9
zhAXkH06pfIZ3QDkYqPiF3aQNbdvwI+oavsaPHqGqbnfpkKkpjSsL9PgBpapoWbS
m7O0wTa8UDDyn+TpR1Fcs7YkfRccu0cI00SyxQE9kUhW92vNppfL6lFisGVyqszY
b3vGxqNDZbwVOjOhAzjH11lIJta3TI3gVHsn6P2oJg6m3T4hQxIqMuM23KTTKTxo
zkrciKORYF8ZTB5PakaQjIwPpY0mhCYQ1dF0X4p+/Y1ZnmN4zP65sVL/Vj/ngl4M
OzRs5pqX6el+Hzg9DRW9+qFJITrOa9HF9c1wDXkTS51bFEl5JqXWtTK6Tnx4nLkX
tt6ACJtF1bZQIRw3ABGISbotayB7c2uwPuwFJxYcxGWJcsiN7rLDTYXkpll4q0GE
EP9DxCCFs4kGkkY4s7msy7y9lNrpGkOB+ro92XyTabWfChp+V4CkL0prUGbL4biX
Ycks9Aq3FrTi6ng+SvQmgUAhE+X23t5jpesU8gZNkrA3DgTcKLjH92u74GSww+eT
SqIlXb/kn5MW9kl9KuIhFQhU67rlSPMxuZIqTospMImKOtnrtuqOFAXUg8HUx1uP
tWoRd+iygwg+w8DgK/jard3US0k9/LeOIbTFUT6QtStK3/swQtAizVj4nvQFViOG
D1A8qQA2PH9i38IGmAVRtsI6hb2najYbsrgcP1+09ExTjqqcX2JTox3Q+UUrCIA0
KZ1nfONZlro7ZZo4YJFu0m1yms1GtRPO3HtW87bAzry7HeNKNVJWXiTdRLkoxGio
TKnjwb1gT2pxRHfO7zNKEuXPfWqGIqLoXQGk/LKX6G6rnC2oI8KWPuN6D8ddC6qt
+KrJdlTVojHdSFSAOaNfEbcqnXUG9kZMA4+cEEUMN/9zRiCbErxzAsMVdMgvysb8
xRMIDVlN+/Bjr0kuSXc6ATorTW65tscy3ORROH9AJrvPhizYU1GQNGYQKb6S92sO
AQlGtQM1eiWKb7Y0oWTTprydUq5WAoGRuqnKZgPdb3KCp5BHDfA1Vyxu2xQdWGgK
swZOgcqIAcdIj3xHMFUqqvHNHOrEtO7T7rm2lW1DWLH/9CBupbIsRH8pRHztj7t7
NVADmCSpY8BTXicsk4lF/qAtOvPJEeSXOvNujKjdoMiHcUWp6GZ/pwbrxE1xAP6P
FUQPEe99sraoFi1C3Pu0i1Glsd+Sbj6saQgdboxPA5BnOYC3oITOU5ye0eQGEFsg
mkR5M+fJPVFBnVDcjXkbVrtOBlolH4+nZi0fwB6uSADw/upsqLbvUAgvV2E1muL9
Km5+rJA2lVGl9bVnxsiNDqzMDs83V9MgfMttrnYkXA4qoCAfAx3aGKPG/IBBGx2g
EVqhIfpW5KdJYKx5PN2Jwdn9oazlKNgtTIa85L6A275Xy5PTYt+akcru9JtScBd1
TKbLO8DnUtZvyfxS2orsM8l5CHi/N1iL/76VZ05cL8KkzubdIJnNmOqRyI358mji
5ymCWpYyAgUbgISGR4mtSyQYzENTjHkyFD8/b3S4DR+Pjv4toSSTISDMHFumS+OR
iDb+ql0Q7rxunVEW0TkeW3wGAqTOY0I8aNm96HYFfMILYNDnuoCGGsisJdCdr8WQ
eTYjMAaes9qYU/y+1I3M1t7FZjHbnOFoBkX66OnKGzB5funUFgSaAvhVIUwD+bXb
Q4GKwDn9TU1L33GSrOLq/0Ei21xn5QT9DcS218nK1OAHsN3u1WBxwzj/HVYuk3IW
Gjj12XMVcSwaxmxCk46xhvnM1dKrNToY4azdmW5uHPVBY0Ax7QhPClrEuGjTaWH0
Fqb4lEpENEuwa9qGBzu6mhIk2hPopkTpeWg/7yEOtYI7SCqfVGeZ6+gEB9f/z0Jn
tpLD2woszNG+2i2wEjEToVWiuopczveTeiS7m1CetmeTimy1eRnlkRbCs7BPEQ0t
IJMOo0O5b2g8FtEBEUTxkop+ODEbkm4wTWtdz9m8Wuozn6rs+W5dwja0rCoz7vlJ
YZBcZv7G0iU0ODRPFBLkfiaghmdTefevJfc/RG1ydOLMgkPBMXuCEFqc4K0NBnIs
WjSnjllNOKdNCTKPfyw4rYATHo2nWCyk3rZkD6BpZyOQk2PcWkTmoMcUGkoDwdKu
oLw4b3Sxhr+Fet8RR2/y3tPSv7aNI7JU7iT+vqtjuDbfo1k7LXxSMk+03L1iGtjC
d+qNBPiH24tRmZdSj0e8ZGLq7sWksL4cJVAlTkw79j2N8XUaf00ksABQl7XkPY4J
x8Z1giMQU7kuEKBKuR+Pwujp1cPgjx7osQvXfMwQyiO5V3GzYqPUgK32MdIm89d6
a+HB8hKHygkC34B8GOz3dHgMgs8g90FUdeQU8uffATJWg1sUPZS8Qjpqj2kA4I+p
rS8Zw6vCYmPgQ0HYXQflLvkm88zbjm/C6WlecKAiE8UcRCmm0We/j+R3uWmLgIAD
n7XKiEs4lvrXhahwPWnJ0Qynb4AOW1iHFSE3XJ5D99HMDCeWb5DGEZwdAgY9XOlq
tAq3ZANY+Fx/MYpvAq2ErHO6SYUKyBaSVjtI14WtDFkWRAWTHj5DjExJSYTF8K0Q
yUXScSz6ZfXuo3McSsfmalJBJIVavnNt6tdMmWxg6vXx48ul+KKTCYd0r+VKRR/1
/MdWDdcqPrvGmKnKFuMIWIzMPom6NpE8zpsTSuIXritJtmpWh5wkbhBwGRO8clbQ
qw7bGQKC0LDsZqk+Lo/d7taWPXIB2nyqmgy2gd0Yv9F1FNxTKFJDJTR/DbxohRbw
j6yF4PuU0zZEFVbSd6srhbecX+qtStQfG7W//hV3zm9gL4i689chvyMLaE7pWSUs
k48qfxVtBwQn+vWAQLH7yYdPj6pRfALLxELSJrMRycyL+CzDRhOkweUBzo9ruonH
9EUrah/zj+60BaoaqxoyBltQkejaeK23SdyWIrq4bhQBQY19oxl8WCcdtOW76nYo
IdxWvcpk0Q3dCUFvByffZ4uTRCFSx6QzZpvReuFowsMXU/I4r0M0eCuKKNSJXIOE
JETZLe099RXA03cfXDWf3UJ0sG/Oz5haoZMHeQ68rYP4RpE2jSfyoI0TgrfKJH25
Pi24M5LsIPTzqO6eV9NvcIoYNmvIkY6TL/9RerF6AL0WZUCm5n1Gfz4xEEuad/Gb
hQbhUWQdpA2F/55w939D8Hvrvuk+g1xpGjRMGZkp5G9m6wEFxljJzXW8B7vuGqNe
2J5MzcR1fjkU/lwC+evpVESAuBAm+4sVg0i4KXNAHczYVd/xiEEJkEQSFMNQcJtu
YBgspxLLtuFw7PhEVXbbF69+xzAGL80y0SgCrB6LgGadBKugL2xPLmYkYtKFk2nJ
3buyqZl7l5WdxGqrkrnfP4bd+UyIICwhkmb47lHCJxH/8k0rzmNVnFqANkJjAvQp
yInvOtnfrBw3VXEL4EXYbvNf9HeomhLOskSE7zqPMp3eOQ3onRrDghmvEWWxhlEm
Y+mTA90HUoEI1cBL6TLyg0IYfaSHaB3abySqHr1qXVGdqJtHTtq0TD6c3L9eUaHn
eaRdk1jWM9IgJKhv6YnSZ9jOXyHlbsN2dc60VhcadHLi5QoYUru3Aiow6l5als7y
H+UNZkzv1JESrduacbjj5sC8Y1Cg8gFtQX74NsziZ5izq3wk4CbprntmjgeNiobk
aCCybAn2aDxGmiKquCh5KnhEL/x8o3z+vkqKO8yOumt5fBTadVecjutsXeKyuZLz
q4PbV+stp3s/pC2g9qV0JrOAJAPVaaqNw22CQdAJI4q+F/Udz8IuPb1S+99GQnbL
ipZQ2jHqd61YZuww1Rubmqmx60lZz3Z194tnlpQSuvJ+xAJtiIRJUpIqmuhAtTBy
ttN2ZclZA3hKcBWr2wmQhkL8A5NfcZAHvk/S95raEXRKFMStnqJDXQy8eplUYj+P
9vkEQIpSNRaCB8GtFMFmBNWOcmujCfmmN8P5YMv22IrCrF2B7fd/ZFkvD6RL2OQZ
5TfI8z2Mh0Qg9rKvGJkEINR50ZUn3vmBODQJVYEKHFhD7c6cgSZExb6eeRYw5nc6
bT95zyBeoTzivILDBZcoE/IEhu3xI8jCLmW1BloxhdrFuXrRAZ7TWyUG9MAyL2+o
VIvLw1+NSLpH7Z0rp4IU6rIg7ns25dcQ0WXDmidhTwlbQRkOOkp/INHEfftdw3nS
fGQOoAdMd1hRgN2tJZ5dhneIQkljab2x9BQzU5pktiikB6DImK7WVWvzBLlh5pFi
5ViViTJ5wTG4axzRsmYWhinvYfLXCrsH68l4jUAtlFutWDzF7HMiamhlhsrmBh+L
d3Tn2Okv7pCx2LAKaxLQVbkPGYmYuS0vyYejkUWNDPylZlWg4PJSS1qMFGuaMYb/
yY0dhSQo6IzbP5hczAqi2NRr44icVpDDIGYvJObjX+XdBLqvvEk5Fp6GYJzHtGjj
ju4BDnxLIfAXgpnhzn1mJlqe/+OMn5A0IUfQsv3YMVaprfTwgyuWpbbtG9SURwud
0Hqh8u/Xsd+5wM0JKJ1mdlbVLR1xzKB6FGO17ZJBa5L4qf/GNfBzxQIVnPmDBhbc
42eE0bMbM7tGQ0zzBMV9D4DPEQx3mO2TK03PmniWNbsbPEi+3HATRXc0zjZxAg7G
xaDWHlABNhJ8dF7unKHllwsOEIKb4k2Z2kmeSCOYl6sLlE57w9khYv75mCCl/4mL
n9yWaA/wkQYeOgq1mOyxj87TrkT+lCQxSuxBr0GNB0GVD+dDT30w2KIk2PDm5V+o
eC2jPgwNNIY+ROOCcDa/X7sQ5mDzoPKiBOKNRHt+vtewqctN1/ZtAjKyt492USuo
cmqfb2Tw3etdcwDdsNcRyo9dNWqqgUqJyGTjECgQOnbSx5+IuFH8XPRjHsDJBHfl
V5DJx5KbxKYL/J/Pf4oZnaaS/nB+ZueOiWdqcWzoF7iprBNWCQ/t8EaamUcqeJKO
e8HL7Sd8M7Sp9MVjE5TC06nUbeETT4ASq3ueyshKythkZIvTFAgOu2MRKuRHxan6
RpnEtcrqIp/SfQXMtJWEfaX4bj6Cykthpal5RBEHdv3QOUNzBTd6xdYSw34B1c1E
3xArZGYYvdVZuZ+r15fQcpSzR50dIkrn2N1AG6oaynl+tTS0T8jEiWj1xwfy3tRg
zuhUi6LNCNIpA0r2VTACcG93bdzRnCWKzkwd33AQ2jspy/NETmFnMg4ApKWKcElj
qeXdTnkJobP0HrbLT44JSvYAeUges30FAIRWi+qAc/r1HZ3HiHBtP0s+9ssuwctC
5Id8wbRn/u1Aars4p/TQFVmBmePHTdWiGFXVY4ruaZ75/sxZdMFB/ioNKkqfJMcO
3hyLjuvQImq74mtBrecN2C6t9r4CS4DYdw8RiIfAk0/Plvtypt0gUc28FNkL3e0h
aYAAHaQbyB5wcOER30nKYD26OlFD7917uOWewNZdgFV5cv1KXg0LhhLppdi/PAr9
gn5na93o4cfXLQm7sseMCENDV2ToXRtZX1r0B/1MtoVMVuPhs/cXZ1nzxF2AWcEC
oMut5xT1C8YqSp/LBJAlSdDHud7LU62b1XWQH8GKXkzOoJ7656asC6nl4QWAqUjL
EUeTH5hmbzDWz1QidBo3jV0qLFIEVkOSmhTsxAig7S9pTUF5TMsEXFNcvxsIKdZi
MSbBHuVVHGu1pufVOQBqx/urGx3DVSLu26aOxdYMdkfiuVe5JCT8BFYcfS1e3E68
nGRoAyatY2SO4w/JJWv0ImiQR6QbKC1g7pStaXAYbiREyZ/6mwoq7cWMHAcb7EV6
hLjzuBuzKJtgXYl06I52QfRvz7MfWAh1eyZv56e+QcSqXu14/o0ehQz1uMhXaPAn
ImrHxeRCczUchhEDin0+VJk9f8qzvw8hZ/mGTEaGiPAE6nI3suMnmE/E2Uhhc4NM
00CCiRJ+uRTTkPACJPY87ZpayuYYBlkJFj8xrqx/IO8RuQChgK7HF7m5N2Uqlvx8
GMVJUbGzeBStadceaRu0sVMHYCg1pDRN4ZYMVcYCQfJDnVH5ykW8o3pa3V6ClOLp
OQ2hNQ45erLJNmoqAQUAKT/9CU8C/BOwFfH9eASn57tjaRj75Atm2P80P+/IXMJ+
ll7bdk5e9a6/+OWGQVWGT+c2uMy/bJsln2+oXpsy26r5SOovckJ2bmPioEvU2r8S
vEyO/1mHsPokHBkaf1wLbmPkMoV0j1YEBmUNqc/qleQFKzRM98GxvTPzyJwOdWJy
p3vThnzi2p9rR/u5Y+slWKmrquBIOdV8gIXvQ1y3XjtAwuMYieLOS4jtA4QdBGLq
a2SHO76J7WcJh2Rr3g7b0rgn7IO1eRYTkDEQo/eIYQXz4Dk3o4CFiuRrFTy0BRgp
Rt28Z6LQ0wrmTCpNMb1o5V1kj+REkzs9OuIcPnw2JJ/obrSb4Mirg3f9s29dhMXh
TTtZADbf9blz2CbelX0pq9aScj7sFV+mj2svdiOiDr3Mlp41eM/RrTHX6INcvPv9
63mK+IKTFUZRujWROzoHRkQSifxgXdcscAv9biCeIWpzejFOU9i1besXnPtsj7CN
KrjBK2A4uLDWkgTMoMEG2G7z2ap73x9rmLQ72Mm0qa8iEmGiOP6RWJZ0zpF5FocT
5b8x24QWPPQIw3QdhgB+ohTTCNoDSVgebLo7AXK4Ek3T7XelHPdNhZUl/e8fP/Jx
BmcH2ZOFJCAaEX8PYDbsEdOPv9MUl4PVZ9Qgf2oL4aSBa09tm1ptzC/qCuR2ZFPx
OEfBMxE9M1dqebVNrmj762bWcSUW2FVn3FEH36wxVS2lYalPM/LmPywul+myK6d4
b4u1KrxoHsx5YttDwztVcddI9lMbyOvV9pKr47M5u4GlgXOBrxWPAfnYiGrgrbqf
pqhgf+vBFXHkCbmzPu8e5qaEJ1afd7BSqCJVBMxvyqqmvz8cJsVzY8DaBAI1ZHSn
LAVvu3HloIHIV41NEecqbJ94F9hnF+kx1B5hhOKzonDwgPDzZCaExmbAIP0p5Yo8
D0vvdeQV5j6sy5YsBEs7Aj/BPYfHTL+AfxdkcZNgLUaC6VSm8o6aAb7dUsWGWxbT
ictOqw3Io5F58ri4gBno/5rUy99yQ2UExq/miZsYMPIi0MIK1N5vnykB53lUeiXL
iZXAd4u9QotH/I6ZZhihZwJE8rDdGi3jintHgJGqUgVTFn8KqrK1G7wI9F7rIgqA
S1uwBoBr1AOfAglTewrbTuVGw5hDX92ZVlC6s/eOpZ9KjgCepuxD9i0CoBkUYGxj
yYjB/nK5JOU2WKq3YX4Gmb5DrtOykJt9k5TTnXvWJWh97Wv/gq+AWtvKcrjuhSoJ
38jMoSQ4f4kW+vUpuw1WNwLOiqEo/KNTvf4jFluwf5dk1Ua2XkYxijY115y8OhnZ
zJiGOLhUyOH0vmUPnsTeWQF1/c28APBA7GCDnFzi8HhWz1VdBJhDGw3Z8pBl0KcU
A/zioDzXH6umVSXHSjq9QgMaErf9uk/f7ggbIkOs5wUNa2MBDW2a6gODisjMziCz
2LyCAThU+cO+rQPiZhWX/mAg2o6G7nj+483hgQhkFXJ9xjWHzkCsNBd+pA1gtJ4v
8yi/GrXmTqXX2ugl0fi1Hf4HVIbmFBFOly4g5zeP9xsL8D5YKhpo41i9k8XkSMA4
FWj+MAWcTgl3aUoGRXup1dg/LOhJm8I6GHw+jstDmU04zOZkhoggywoe29xWc2Vu
HiIJ4DQ7rRC2IPpbyk8Y0J42XzNnEDyBc7a6sbzvUpRR5hKHwsL95IMJ3b7xbEwl
FlTL/PCPZzF6A9TXFdHZTjFp0VdSiiSeKY6pJg/U+yVCea/iDrs7NGGNyizumh72
HhfSzh50PBLHLeghH9fZ+x6CZNBSCPoWt1Ahul+VENH+lC9JiHqjZhf6azTxO9fB
i3Mv4UJ1EEhnU7Uycxe9FzSggvmIotSjjVMfXwx0iEM8YbXNATyGwBlaWf6CZ71e
bYkDxED6pWF8zQo6LUJQ+s8n6362sB1J2grZ6KQx/1Nt95HmMbKWb30dBk4IE117
mCHFhKbHwSGDyN72PueXkPUjIFFMt3pUwMPNxj4wj6tnqS+cp/DK3AmnzfbC+3E1
GF0oaWz4LLOoQ/HgsGAIky0U4WEbmQyOLHtXdgNcWlFGJrC7xpmOPpoS+E6gSJuw
6KwuLx+7ri4K/B43VPKYF7Ylfm+cdJXX9YHp1CCjgmfLhzNMGXKYA7Wf3LA95x3C
ZT/vzvKvDFeIm8X9rwY9Ny1SdsU5VVLMnVHPSEEVPyAaOsEm1BBP8oBiS1Yjv07N
ppH1gIdQI/5N66xxErYm7CZNlKHl+Fl/PrL/RUgIDCZry/oyIuKfYRSXzSGl6S3d
F3uQY4wegbtMPcZHn6rLyfwTIlAeDQarHRkDO+9Uy4Nd6SCiesvPK+IYVCJqryAV
5abXT0Wy3aU7xsntUN0cZNlcPTByTCBbn6LFeOEwixNml7+Bk5g4Nd4FfwUKcXN5
lEr05CdnudDkvtX1rEimii06Px07ryoIJ/FUFhNDngxfSZksPmYfsycORA20o2Zg
0GznTmTJJZ6X5DLxJvzxsE/Nq3IPrHIeeVSW6QzxyKdHtcw23ouzVzejRqx6/HSS
qhqvveKFWUn8m5bHBosdd0SvpAPzMoR0dxr6mVnjY6+jQCS4fnHr8s/TpV/erAWU
RwpPSlgI3nr6g8vr8EldAK757r+NUmb+Nqou6EpZvz9aZtQwmCiwpCBFxkhHDfWB
+gjR9xv9xHpTKTOPCKe+Q/adK+6RewV4qBVV022vRg8KcuGTTFZWLfUGp1RW4CnK
bEQOnEiaMUtRacr5z46GhgYan2/KVZqnwGw79Sjhihu6KvVnHma3TO3MzopcJU0w
pN6y5XKI3N8rVMUuxA+JuOPLahPiqlsyy5lpdCeR9LvesRuud+4s89Mzc8jo1BtZ
9uvmkLcCN+LvUJ28FdYr1B6W1sxTMqTVwPQ0JEwOlTfG1Vgm/hA77xOQ7FHUeCXX
xOlaz4H8zqnWdPgUF0fwT+YmIp+sm/NrNnTn3cWdpbpEWG2RdgbA4h04UDV+C59D
T6IGiTme8cg7ikJeM8swHRU2xo5KZ5Gx7CTs8jSKhkXYe/sRynTTbvCWvToDVN6B
6PiypbFWrGRWg2negQQNAH9FASPdg0UgjH0pNB+8CWqiGNTIIcU3H9Ttmk3X9sNN
YtubApwJnelI0HOPOZGUY7xUdLFFUnhceZahItX8Iyvpily7yeGHsTTx3yPluxi7
3EBMwhAqSml8JiEDvHXSOdn7gC7zaP23GaBQCdCKz7gHSxDpoCNSw7qmqKYPfS/H
8O/mjBHPRkK4goquthQe+I+MIrYyqY7UjexylCEm5IfQ0bS8RjhVDFR+Se3q4meU
1DWrqXUPDuzR0GNDiMMgogva7OTkpZAYEZDvm7K5Y3S5RS/ErGy0YCOtmMC4e9u3
inqLNDA1UnPagueztFJ3+onNcIxpmHpgr9eCfQLyXN/mHwtCF/yCLKqAGekVKL1w
LNumNpet6nJNWGEnVrpfnt5ukXUgGsqrcdeRclLp32UKBCdSKx97j1V5HvO/TQq8
KUxi1+QDp0+vIyBE1h731qTm1CVxoY2NLJc4Tx2J6UJoNvglbTAtke9tFPG8ddx8
7yMdK2uJ3Z5+RM8jpFDa9VaSWZy1GLz656cBphfLNos9YoApqwViQervba5N/CcL
ybshYCBh9vMhqCjHPbMwE7GN9mpbnmqr7u+OZXFmGjWknICXtcpOX0Pj1QewYIjo
2kU2sBv2hcMnoAnbDS+gUNzlzl6c+dViQDvLEyxpXVvWzfsuW2vc70I384SE+s2X
5YQzMRzCwoUymFQrx7z9WSQhXLXnJYlue29VRdCuzI1o1RjKqex6n1kIAAU/D7pt
s9GvwIEPNIKEbO5p4hSBTMxzjO7JmZsJwaP8orQ9X9Zb2npAGjLrQhYNYMEcRh5k
FHT2SPe+FJZvBWcK881US+O/8c/P7W/9o7mHVEpLSrimPFobqI83FZd2G3/A1vHe
jmb4xs0dskGNjRk25ZgkrbC1RJAmPAjotPONX17cor/8G7UgNa2INv0h1pdDqWiD
WngVsv8KitusoXzvsAmXyjc1bNqkPW7Exx4C5FH4YxfzlFpTCPt/cSK4kCip7WaC
33VxOe104Glz8FpG90rrKXpZAl/qs3hYDMUzJg5C8Sx9RKFyS0DN+i2nlD/vMLPT
FOOFh22EfCStSf6RtRMMzrhIzj4O5pMk/UeFqkIqq1OOdvKpli8++0OcdYkPvHQS
Z3BBxZZxhw+S53hxCwwSi5zcK+DzCzEwkvq6OTdl2LP1fVBgXayD7SR20OcR2MCQ
jtE55c8eO4P+wM9+ABNKQMzO6K1bYtgwqxAut9MMwJd6bFc4sjK2Q637B7w+uRxD
0zJqUigW4OUxDKVgV6eFr0ZWC9vRYQvw6usS0vG/CVOayBtIpwVdikkgf92QljWq
A8vN3T92p73Wvo86UMj32OCoS7T5d7zIemvV0yW4sLB5lU9Hw1yJ8BCz55fzUFXe
vGz2TzwRdSSX7ZwwCRsEtMaPK9rbRDNS7vXvF7scidQfjLEpMsKOURMjFDz6GNZy
lb3A79EmwHj2qJMDH/MVkX/EXtCXHSQlge6KW3gM+Cboz4w8gWMDrlExSz7K+Txl
JyoC8yO0WR2mqI0K2ANVKs93DXYTjR9wPDrWiqTVCxhAZ3NZNzT53xGXrLy1B9TF
b6xXc4wZ8GS5wCo/UgbLfQuVKCfDo8vEQb6l0wRR/MSXkstpVP+XA5rX4t0xkcvY
lfwizp3gnrcIgZ7Jkn+yXjbi2++0J3Lf45HiUs5zVINL/wi5yhsC9dOOf6JHngG/
o8tWXm4w94ai1FR/LYTW2XPufwqpwAM0mk44GYlSKGOOUnR5j1BW8OdokVUbrdRD
DF33V4XQpZqAAT+4FOSaPEfSNGYKfI4ogiZkAsoAI0nKI53JT16Fjr73mmNTog8x
4nY5l1GopA6O/CMGf097Lqa5k2u3zOIcVnJblbGyrjj50ClupaneEwpSLwDyC0Qf
doqS+VnxlwCRtr5zSZILkBnqiqek1wUkCnzQxTLRvy+IcMjjbsCDHzkEOOMUEM6u
zLwqe9odBhFn0k40k8S6/AoqEqCEcGA61Doqd8/0R9SCLAQzP2s8Fp+WFPVi4uts
O3TE7pyJ9q/e3wTYPdXPdz9sz/BGfBYryueuxTsnTCj/PiXDPpNY46xJNORjoaDk
6WbHTDK3zeD80stKtOEZ5yDPc+nlwdz+J4BrUGr0+ovIsMIqCRaE6aQ5ooSUUqRp
X5EkLumBYCrKJKPHpsEyx9sgrsDJEKNCWrOla4nGKT12zbcUgjFQmAgPhbaIKgK+
iXSN01SLS9GeSxN/v4aYEu0H+VWYUY7/ZsDRMfFsXjmMxD8UdxYpXe9NEFm1eZU0
iwg0kjKb6InjYr+olPr6BHmaZfIUWxEuGTNVNFertQxqP0SqfyH5MZpWs5Se+gFp
2CP9XZtrRRIbMUs/5MGjK+jqIBjvO/l8t/Ba/Mc+2AdgWBNUIn7sdysNwB9PKjZP
EUBOvIydSjVC7/mByQe+B4eUy6jdk8uWP/d54M/UhJMX/Rdd8QBOLS66JEerdFWl
3bpTTJ4HlIS9pexpHqDOwgBdrUlTdUw/sUal9RAJslsnN4RkjxL432jLj+zG039e
WHIEeQUBWMyvy+XRRNmSAYClWlkZi9caeUvDn5RosCgS6IIdnFcWMm+AwdfDK4Ij
8JKiJmGX+ZfJJZHv5VVMgkOd/AO+m0l/yWaadEPWsCQrDI5dVBv68aZoCK+h5ByY
8dAaT2Z6DUVnA8Wumag+KU/bUB3+8xcWj0QYhtbcz1hacVvoAE+XWOK8BGkL4l8G
PG8WpHJQdGpIBvxTCBdBkxd61WT9kH/X2SE1puiU+I1dCpOYJChvczFxe0Tt8I90
zp1sxNJ0tdSaIITZVHprcIauVYjZUvtP+99zU4J7EPb20kQYZu0hbJ2F3F0ecey9
poanHu1J4+w5l5J/2vE0k3BXKAKpxZHfNl53iYv+q731HMhBKWwV7I3+RCoyfMFB
JVByTT4U80ncDFn88qaOQQnPN8a3AvJw9lNZGEcFQnx8uw62aWv42W0qCqpVRimv
KnGPplyy1xCruzK1cxub6rcVvJr7+5DYNf0GzUcO0IcSD36L/DwhvQ5FggrJg4Hh
BdF/wPtUZY3HacOGnCUBzhHcjCrIB3294dm5JOvGTWVr/5rVaCMQbYPgRVivdc7g
B6RhvXS4C7ooZfgSkpN4l+LbtDsW9QYcRGGmeqMkYh7bwLZR22QqsGr81XuOLPpn
oUxGnF0h6W2/0uQtcISEdf/tetCO/3wV4Ltz0IkXZpn5uY36GJroLKJpC7wPcLXo
luqTApFsICO4hXCRyDKH/BUV4CeXiqNlh0RU1XqaEbEpbyPgRtuQr7NKg4nL+MFP
mneVBedlOGH1IfCAo5SXAiXVZSE8o6Z9BPjNAyVCGfvBYK81b807qkqgpIdmkzGB
yX7Tbg4Foq0TzyT4VT2AVyZ0CzeaRiYSJZws2HluOSlZbTZrRZTOUIg8dY0CK/Ul
y2dvXoSwOkrNlP6V8xf9xEXAPoV2LriwlKw3LpcF8qUt20FIJWAk/m88oBKEEn8U
DUdKSgqHmLirt1N91zYu7mmo1GCNulOjx5hexkgO0PVWcrSLzaekUtxr29ZjOG/j
T4fPgYePg4A/5Hu4BRz2LHuOAzw9Q7IflSJirVwGXgcK47Us9aCQO6YQI63/PQ5Q
cUT03+GP7f19MlBdaHQMrhxO37/PTJ2h2VWH5vTHcbg4KVp5f/pBNT+yrjvM9pTk
8zeGHRZJtXrzAz776RZNw0qpr2SOPNzzWeeSKW4L7UrGDzh7fVR2+X+YUYCLmcTy
9X5OWXiJ/cZy74MhTKWTbNEFFPOB3TTD6PDeQEZD/qWf8nrYiq8O0IKlujgpVjBS
ukeytUd+yZAEhEgtTWbGSu3EzumzQCIBhVNj5IJ234Xjs6sYM+ElqXYYhiHk1cvX
MIL6EFg+8z2RAFiz3zcRn0qvmJE8iJz5Lj8bJ5BL2O6eH3a8OZyDATlsCax1/BxJ
8z7L/2ucribf/oFoebn8UbZlnA6ML3i43F3OdtAW/IR+sEtbdWKV/eQbYiuKFyPZ
CGoXN2mgp0npbjqyQmGU7FDZgfw/poxS8VvPFIsToHpYTUmoqcqjwGVbbVtZjz4f
krSxrnLQRZuagcEvf7qXcHVVyspDhGsIG3BLjTNd/YSLC1xzlQ1dQp3VTOWw/g2R
Pn1GG57ouIfP3KX42Ocj7ZyB9Z63WdKiZfRaSLerv9LgwwglUa4mCtUO7fHuMsdN
odcadNuHsl5LKr8yNbApup3KK8rpZORr36Q/GAbfzJXqOsCNtUPTCyti4yWLIdPu
nRRtQofEbvXUkjJp4vJvYivIxhzOOF9n31sLMBSxjbEQ7z0LsD7y39b6dqih+anL
WlW2sw7WNZCF9YlCj3oP4CtZLWyKtv5DUDTKGAe02j4ExjlePe4BlXxafWyGZFRi
foyC4xGwgrRqu+2hRHbnmV77M4kMUFfKFF+mkZUDzlziNqKshvtkKJwXLv87uAGR
G06FvvSOJDhM0ajPgnFqvLr68dyyKscsZYuLi2TKPR4H5yxg2tZ78RrjTdXP5FxG
Ep32dX6eyBYeXQfTbmoLG2Vzboxb+9C/RMWrwIdKe1IrZwINkx4gS9XG1Xm/w12E
czPKzhFXqT886X4ev9wu65/3ywfIAnSWccBiz5mqQVHyWowUyu1ln7zi2yKtXTSE
t0Hv/lpYXesmijCPSCTsYUb10xoWnYricGZArgKaFwPqSdjFucs03RkmEEfJjxxT
woWKVZh+p7w/rN8CO3HKdhFoHRqhFd1yZTl/bJualsHU88dsdBrVROEKDc2TLq2V
rwD3L3qi8J2fnErLmrHuZVipt2Fvs5ouWryYET8dd8YfR3H1MhY77Eqt+r2nvWTP
ciPLPHrcf+lYFMgTdPgPWe5hOQ7s/Lf8DErLMCOrDgpp8Hy3p6eVUfrVfVgyxhRJ
C7HxJSfs4SkGgwecUpCmUcmdRsSqbqQ3P9u32AI3tD6LpS9VHknQcwoEQgYTml3A
jo8Ov/rPdjsQC37VfTYMYBIjdIUT4qw2EAqsEUBqzUEDkmDzyvWjcauGyEmoIFVH
tzul8yusiP0m2OGOtEph+4wDlewV4CxnP8f0PkSua4iZVeiJlMA7M3a7pUvTYjQK
gwVhXkhoRpGWpImS9cWWlL3Hd++M7bKjwLkUL+FxNC1JQjPgcbDE8wtaT8gkkuUB
VjfEKHxdHa88si66xqLtIR1rVXAr8ygrFKz3DlhYidwpGuVc7CtSu1+nFjqQ2JmX
TBKNrplPasAY6DV58OtyJO3LReV+oMkaKzszezygys9mlxfSqe9zGl9+rYUUIzkx
samyCxrEP5AVIGiSC0o3vQz3oewAVkaVcoQpxMSUJlCGPag0BbTGFJCSRXJqrsRj
8AgiTC3EXiBtcK1zx3qvkTVkBqtkp98Tz32GWSgjropSdJeFz/lFtptZNvpHC097
VRR+l1VuwURCX/Hdy1Etj33SKD+UcG20Nxn7WBONG7KaeoFqRLKNRLTzIm18Ekdg
/Oq6taebq84DNoUWNZfT/+aiKd4N67zD46zFguruHH+m6AZrgkGESvKAYsY0kUSe
dXqIMDM43rJPcsSnoU5ods1X7m6OJuh7EAvaa27tZerGms2+bKgGB0UPgnXPfJJt
/qRjwpHaEm+m0/YgEyHxSpSLshZYb1mRyiwFUHXGr75yAEG+7GNLZMvPs3dWUD1G
RonqRK4YAc7e5DuJkoR/QQBcpjst7NbhUkXWZblaCVREMGUw8J4n9pbP7Y/jumK7
M2qFH8IRT6U2x7uB+NiWuiZ595KUmYyI4RSUnm6V/Qbpy8SlIgubxJ5iuR1J6EuT
HrPynhs4Qog/FHLOZBHH2MAOXmWpLjPTEMJHkkHjYs42a5pu4bp8tJbhXbMn+TBh
MCc/iJQ6fCOndlgpFwyZYrD+6dSYdLBLsFcdN1r+UG3PtT7vlKx2yimowDQ3OTVq
gUnSUfhNMR4qbhynLWKzP7LbO726dOqyvNclFY/dlifKIUjBaNJTIvlvWwJbgUmQ
zlxI0lvuzFf2S6ufY4rYofXb2PK4ocoG6jPARVs79p4zDarQZN5DouYg50AYD5Nh
sPfx5GOX044x2lgejDx84eR4aG/WzsdHX2lHdV0j5+fCA5+vcfA1tNGkPAPLIKKd
2PY8Nj7ISlXYcgD8nFTRRHSlaQwxx4aCjAShfK1EomaJ/7kR4DilNk9iNH9CCDRS
I7ugvXm6jc7ZpJqqAdbBSLGETA5VIZKQjG3Mw+fyL7TWtjTwAsHDqBmlwsJlp/MU
dHhO9WE0bQmyqWtAQpCxXXdRWVjvcLmK5+NOsuFxxKFu+z4LvvgzIibH41BTauLr
dzpq3UQkgjKPk5SfiHi9gtJNvkjwj5iZ/pC+/zkD5cT015LAAeBvYzxPvawCTPSa
rKF3/AM4W8wXJoUguPAgfFibSAzgwRZ26AOC2Sl9Ry9cF6BVHLP5NJsuWKXN2BRR
poyvsL3HfGin0DI09JiwSDZvEiI9Uz0PVVCtKNsRg7Rqn1+XnPJH9afqQYMZwiLS
jGaHDHBNcx9Uu6DZeA/wY6IuVhasVl1RXifjnfSao3oMbK5y5JfKdsE6XYYylrn8
biGUWWFDMgnTe3RfaGKhEax49TnhEDusz/LXbbHAFOQacrd7Ucru6oelC6+rCLac
ofIiLvyEPmKsdX7W+tKuUD/PVmq2gMAcJhgjZjH0na8u2tbXAB1V8i9oc+2dg4cJ
bi0NO/156vta5my4yYffwpWUHaJH+0I0xdZKpuMFftqLmu4Mq70/W4M+ezTAzzLy
ywBvZXx9xmdVVl8OvrvHREATEDrA+2URk47dNB02q9PgzMNCS3EEyoGAyrifMjk3
3pVxlZLaov6/ojwqfEj+CBJf6ZEefqbVg6SpNPblUzlrQT5yzlFL/svTt2Rkfnop
psu46186Q+2CZyPCSr8SuIJo0xMe6w+PcT3Ulad2NP43bE0WTuj/YiHKKNObqTSP
sgCbET69tRe9x7fgWEp9UIsigcEtFpbb3/CMlaDbci+CZ+8AxwdtbUlQjLz3c+Pa
qzwcekhsVX1uaSH3/BNweBKIoWs3hekYvoOSj3b2NF6mQgjQSCtks3lghhh8OVUv
gd+UPqy4rxNikCDipVb81IbSKovFDgC76Xj7DBLIdXQ4ACl5D6UcE+pMb1eSl8B/
kpP6bz51CkP9Q7dmAtn4BBvrOFlataL4xXN60LWU86SFBPfBgOIhQ1IhmjvOHOcx
mmA7iXvNFd2bp8y1/JdAQNTnBQAYXI1aYd9by1shi925MEiJXeGSN2r+j1ErxcBV
fuN3DPardC2ZXUqoXzB9obx2Vklef0S0ph0XRxGNyserT69XzH/Q/ujQ/k7qNchv
R60iXrqIQ9HPIPV/Of2AstTkCisb+X+Jidpc2Ah0O7yvm30N9b5RQ/aj1WQFkI4x
0TBzGhbfNsi8i/S8or93X33r1HnYZ6gc16zapYjf6X0tXKJhyz5DGVsZZzE8fMdw
Ncjo5SmBfc2PZ7nMLCq+XpZRJtiMdkyIxMFHpkEvfMz3BZ7I1VopOarTs68xQwFA
Dq1Mnp/TWhz9MUbOPQY5JzQ2hIisKwzh0/Vhf61sSDkCxUv97XM5kj//e9vw4qoP
lypQ4CQIquqKk0ugxPLA8qHaBwHOdPpTPh/AHFZoAbbm/rTlLA+DPZ177J0fkoEI
78Qalt9TtfYRDRUQWg7NBypZ871GugNzOQs0CWDyYlAOoVLuGc71mDFQ9HgseO5i
HAT1ZLXttGyo0bFuZcKrKOkcoSO2jbHF3w1wd9aavvhTynq43CzZSaaGtbj74U8t
xT5uH/8wKgtRktWFwbIkApG9FfuKZ0AvKGyXLMFlV8td5gzzL82XrFpult7quUxw
/hpB0Mf97e2Fo5wE2dkxViIx99d6klY0XVYESCl9DHDl19Rw5yMl+LHvuWEfsnhL
adV9LS6UXKsz/rfc5vi3O2wCF1c9J+iyBL8ncgN2FEfFh6cCJTHB3L/8G5KnTjFG
Yq6z8pHfwJbllW/TRsTaajE7dGna/NXS1haGtR7x58oCzHmkdSYYWTfn10EEhDMA
RihpjXAL61OLEHNwEaJvrZddeAb4B60/OKGr7eEODV/tN5xb/GJMAJoGYCqQHjCr
BjZMEXxjOUgKrIZLqWCU6DvVqB9IT0Bgde7lqaZr0poqgQMAoIJNifjumjnQ3kr5
DSFpllYMhE04a4VE20fCcUa55BvDwBVtq9h7BtDpc9H3GFbzw0MueuEhx/UEFl6S
Q6KXffxT6+nPra9NgKEFg0ilRMZICqQ+wwvSqz5jnJ5k3nuPIF3bSGY4rRmEGsn8
kXOJN2FxDo0YOk3eN0ilKyUIDCD/vZeoShsR9u4OUW7ha83yh+xryVeLVXuQge5l
zW+9DSTtilzUHJSdIJnvFrFm3OS/RvX3FEEo9OTfdqu2EL4HPzrgU33/1lzV0AEj
cM4rbOIFbqzM1E/NP7JFWj8hEm0bJlYt2GLEQXwWv4/t12+HQo/3DyYOyfGyLK/Y
aqKHNdX0az/21f6PpNOPSWZw//poFvYET/ddcyiT6b3/ra5PHdKzJ4xLwCpreF98
UhfgPh0qvNFyM4ETKERCd8uFbmjO+R7Zk+nY54TjW5RE3VQBNCTMP51Lyxk4SVx+
rU696pXRCHilANv6MHIhvAnHbZbfNk7E9/ACXjLZdlFsEQgGrtmm/qlY6sO1P2OD
3tyJSGU5fHhwlGwG/vNngeem00uiURSwkmNDZqjNDVP7xceK7rLyJOrqd+NDqzlA
xmv6UU95MfKJigEcRTUVGTtyf5nv+soG4k2GsftUQPfcQz+sQMdo3qkN32jR3qir
LDCCffMaGhFTaGXzQy8Xaz1UdaiSjLHZFunIezzpsvgKHOe1jENBzN4ZdzBh4B5N
XQJXPCYbXCuOX5DijVg6fd3Kwl8J1hNmXi9HtWzCaAxb/7sVhT+tcn6FC9oK07GG
lym4HcsSD6pHL3YBuXmKrlxoXXXJeJiqj325vniDYbU96rz0bqblG0i1VRG+VgPR
30g4bjNo77awLDiZhNW7PRSBbDQFyKe4Qe+sJvHH/aYN3r02Jzz5/mvWKwsO6Glb
Al3130U3xpTlIuIxR+FFqiFOqNbAALyM/fvd0vGsm/59XXofpMB2IH/bkr1VzTWA
v4KcSEESEsRSMrgC7VotbuCeTKxfyEvdKpkgH6ZbC+9f/WIM6Qn5YyCUz3XGE1j3
VRvkJy/TT0xm1PUlRvFVaQya6aFgrW77V7lVXj6YLytlDswqK3HjtNf6T1SqJTSe
QzmdnCwOdlc6ctfiXUMwE39MGLmo6rSkASRzuKfEnLdArmkJkbMGAnna/QE51UaB
lVM0PH6bR+5FM5IhZK3MDc4Sx6J1r5UQrVCrWPGJ1egqbscSqUoFwMC8SvuolY0/
xHs1Sez6CT3sPfAPk6BkwKuvNw2Wr4Qa5fr8J1/MtVPerbQEGneEu7BHHoZGBg/T
stI1mVbJlNnhioL0jOLhI4vFa29Q5gzPyed0oH54tJXO3CPIGpl2b8ReWo0kul58
M0vxCQIZTt7NVOT8YyGnGoHCoEOJ5rJUulmfbvjkml2IWpfQm10OJoFr9jos0P4j
PpUA2e7fhhyYkUmjfOSYZiBuTGlcWKDJSUuUSwwFBdD1Fk0AlhJYuyiCuWMj1xhp
HMAqmwQHyAYKyhfIOlYT5mR6LCTIE2l0cfRg1Dv4w6UTfMawcxXDT/3vBBNikzKK
IKxbAlcKI9ZivTFTUgk7mC/CjyXI2T1rPe/ZxqBMNP+jmeje+BomCWfRLvIi5h8T
SrOCAjit5FqVCIY86Moxin7EzNHpv2s84FkyugrbP5L34pkCvqmU7R1ceo0T6jNN
NvVNp0qJs7QXgtLW1GocB/KPsl7apO2KKk6ub07WGWzmPcavmHnGz9ZXxddVyZQx
WRBwpLxq/WTPLz+mGzAcK61vFh3M3qCHYGR9RYiXVKCu5kOBtHM9OPXHnCvR/2bp
OTj/0oCaDwpDJ5xZozEAI4bdzghnUlRDEVQyGN75AeQFt8nDIMNmsvaTwtSPRp8+
EaEKqqO7tkZa44LXCmd+kDNk0MuWek/ZB5OY8kCeD0saasZFdHHXz2Z2IkUNY30l
b0AZzcGInxpq9+89OY5E0Wp/Zj+wCWNfFYzkgtug6+Mncn5HhiSLM4ZY+7bq4z2i
8UM4jYjRWctA8waGxBH5yKMUpPVkM8bVMuakUDpLnRANNH9kwWBZEJ4SxilpXd1R
UXiHuwEYrUFU26q/gA8SvuARqXZU5RKKbUZx2/kW8Y6NdvJImbDWAAkpfenOtq0R
oo2Fak4kMkXvr6LG/vA935SAKOr0fIHS4v1+daOjx6KJCDqw4Q0501Tb3gsOxHgO
nYNd5qomSI3C6GPmjefBc7u5QAIDHrQTBjqZ0sqoFs4thKDA2ym65HxzkgIm5giT
PLO+nA0DmkJb5iBB5psBbRSSaUtU5gjsv7ukbj5aL+AxI7Y2o6WNaszas1hU+wu/
MSGNH+hz4nmKdpz3Wpbu0Z167jdE8mZNmTcsm8L7RzLjjftG0hDoOUXkvEDtzxXj
6jc2wzB9bWEWwI+CLV/DiRJXd3vGVvJ9VLIWT7Zwl0twand6xmJaQZWSADFZpSKw
kMsRidHLIdKXLEbwyz9nVNJGkAuPua4mhSCiPE5mM+qmN8MzGl83Zxo5dLJDnknt
r0bSlTakTG5XvOvYDlnovn1jsZquewFJ27jxdZ0Z5ZQnQ+Or10tcvil7+WHKZUfp
zLqSqcsKG5vaLpTzz82NCJSwAV6UexvN9KlMOIcU3Hf2gf660eItCy0NFFwyEmv2
LC8+UBeik/xX63qR6xwaMtKfLjLuo/VpZZc+TIiBq2mW/oOCPM4run4IlVDxpLia
Vi8z0HZyOlqyCk07ZPq1EkpOtJk/9Dxg4R1Ix321e+yhmC4bej83Wpcg6Ig4FdBC
ica7ZdkidN2nukboAB9ZIlLapBTNWmsTTGketwBwKYKW+ZECScbw0UmAddLmMtZw
EcAxvE04LhLo9duAtUeidh6xqUrH+IbScongyEN4Jq2vg+/HgGUnuQEJg2H0b15H
SSRb3B99NpwR4pt1eyV25IynakAYZcxBpTZgU+/NnKv8dxcvo+rIuakRrrEd2m7N
2jnmSP7XVHApqcmsp7FY4/3G0sXHvLU9YZEDkesK68OoWZzFtBBI4WSzU6HaU2+e
kZykN5cNjqCMFFR56A7KReSJ2WPA7XElTGkWRLCS3smTGA6Nxi2jGSUfAhtoMowf
zmEZA7wPc/ZbHw+OBtB8VV5Xb73NlUzjhEiw6sBjECbOVxmmrlz6Ygslr1Vr0Lpr
xfyOrQdRyKAGu2l4P5OxqnuTsh9R8UWSAP/yvAXG3EYLKRT9DTyJsq++wq/aX0Q+
PXuCClk6Ojee6uTI7nn3xO1lI5n+6Lk5b+YffeNJ31Bk68LmoPZ71+JbutVjszA7
i76n2gr5fmDGjfn0yorn4VwgQF5/sUBvfhSVtD7RJgLLvFXcqXmEgsx4JAPDp4+0
BR0JBlQiZx7P0EqT5pvN4fN72AOehk9n/tswhaF5XXuU97Tygkqt0OZU0hJza9NQ
hVty4u/pepxjeOr8CMVpq+xzMkBMfB/wsDircQvvfakMQ/lhJIibOLnfuAhhUVZh
AWQD1VWsTNOryGthqHj4FM184woUiZiLtJ4ubUl1tHuv/dvNjQBKs45LoOrVCoI+
rWTqqlPfa9z8OfQV3Y9am2vn0YDmrM0e4Q+PEunlxIVUzvJowUSzHkrqDugjzONJ
R4P8rAexi1qd2lJ6UGpfr557Vj22P1i6okcb1qBzsDZ07dWGpxQpqEkerqc+aQYL
wGd3taRanuUiRmI08lZPr/W4i4cMHwCrnOUflVAlD3SlrVEmH1GkObhY8fNMMi+3
un/oLdojucLKpUIcgHpl+KheBfjjQYqy9r1lB+dMtzGQ3cWDk9Wei6XgtammbYe6
UK2GlRVel68npVMU0Sg+ou9/nXtdptkiqxjUNYDo2OpEIs1npSjwUrPghFEe/cis
50SvbjJsEb7IF5XzKrUCNew3w3cmKRiYOmT8r+KMixTJVThAtM02mWvZMYdH3e/z
27zmDvPOSF2JKdIsias1Eh0nOC+sqXmqensDbUchpVfQxPJouNb7w0UnKm/mHHTI
BfVErRiSyllt31sxsu7uRSb2eDJeSQ2MzOFk4VxAi8Kw390kFh4tL1hBJG5TZ3eR
CXDIsg59vfMZzqo7S5Zhwgm7xr1qDI+KnXFmtuein11j1zpFdRObU4wupQE+SHDI
ARRMpgOnwJeVM4rYy1inotzjfxUhc4za6nuYMKVLlIB+SD/ka1ouXlRlCOYJhubp
ZhYSVc613YemmM104wT1iy96e/7gsV5lfXI8rPGsY24F6vyvGrGpctlTIlj3V9e/
E71uLecVpw/6/TRfisvjCl/0uUcNbn5d0RGfk4ouLH0zuDiKnW+XBB2VaQ6a5kx0
ky8RtJ/92IyybXapoToGjF/skCQlqE/1f+5SXfnFRHSPcfVBiNfiYQ6Z/MC5D9Yo
CPC9pPq/NXdIHP3oepfdUioYwSNcZe0r6GsbHSE7MMqtUZ/bAGWlyvfUrPey319P
1rNz1hlnNifzRV0+QcOfNHR1L7w/TRgjp3akGGt5ForlztrXoSwpdrHx9WbgYawe
QDUbSdWkH2ggqPp/wmO8f1lqhiU8Oxxs3cYHjShfKmss1x2NuJJYB1bwn42YkQwJ
Zb84uElhxIiiKTmEtDNdMie1uwPWtRDfNzH3xi8/1gMsIjE7dbsT6AHkEXXJPJsr
Fu/Mt8YNl4ixSicOghOOz4Q8B/+LShEElVIm45e2GeSsyGK85Hs6WxLhTTJzrkYk
a6zPlwlzs1p+s4b1WQCkiBuniMSSbyc5+2k7A4myjrXfDTxEjh61VtrduYAq4tTv
NW3ukHZwzx2vKG3BimRsj+Dvu2AAXFVZwiGKs3V0zr/MmHrQbjzCmWxnVztPlCyo
lO9NK9X5xUMA9+FqZ5CCSwmF0TP3FskW+Cp/W3Rqd93Cjp/ePwPSKk7AQPS1Pc9x
hJVjf55/1db5IMuPs2BJ1VG9ojwgrNy3B7AR83SoNY2Ed4ri+7ANW/9Z+qgENknn
QUU2LNpUqCKj1uOBXBPbqzINZO8OsO4A9lzatsZkpeeIgDertHaTwKincseVOBlw
U9utnApCyLoCng55O0Spj2Pk9/YfOk4ql8hXTJ74Pj2ajldpNhzyJZqmqqWzZ0p9
TSRg21zWzPlHlQ/HmBjWPSm373o0ZTdW6X3VtQTaFc1g+loRJo474myuDScvo3GG
BpgUx68jGaw0ZwJ8Q2BxqnOL0FqUhQBBrt8JHn8TTxj7+A14l4o3uJM5EpKqh/T4
RDd8vuyVuJFjfVjpinzg8lMKPnfqWMKXnA3aSwYw3XPipw+egXQ8bRgoriKej2kN
aYduDuHp0SEYZyD8B3DdCd+HtajGzoPdTsTus6c23XBp2DBFbwoe0OL/FL6FWFCK
ia+n473caEQeMGsTWqdOuZmQZfusqc7wrTEBow3r1VyVouyYY26NNZ1QK88s29Jr
8FQq7EKZ4qxChiTZkAnotTjBNUTJgzSJhalotf+wGEsS9kjGXrgz0SxlwDqBnyCn
mVxFmoubLdDIZ0irARao0s5Z+bPd59ScCi35oFuwI3PGmjpJQLHf1TIQjYUhbeMH
WrlsAouw2GRYbEQfoXY2SY/9uSqRktlnYcoGpTyIS8h925E2f3bXqEzwTZMX1E89
homPz+dil71rUDRcMNTY9+F6xAe190PoHh3bKz3iC9F9FG/PwJaD+nBs78G1v/K3
tKtBVQ26+ZW1D2cUpywcjt2CbVLEwmA+UY9QB7Il5ACKFoNAKdwGq/6oJYjp9HSg
znGC3MPNYJ39KPD4IlzKVbN5k/oPeTzvNzOBhEVS/gM7b5AOKnyVq9yyXRpt9rSK
NB+6QneZ80IgAxJrRdpn6N0FBNkdGxc+dguk2vL4I/ey4jtG/vGowrP4xXVydULy
NJtdrUSMDKsDmln3u1xDU+RgC6Tcui59jXFIKVA6Er2V/hcpvzIEYYxyWAHSOpfh
f3rVxlc2AXfOu8TwU6TYVgNpA01EOJdY94gIiJOuB6eG63ppKTPWW6ep5VV6e91o
Dwot9+GkuYGr7vn2qcA0zTlfQkhAgOQ6+D+OjCW6OwBAr/9RihTB1hArWvuc1M1E
UqDGP9v9dHbMuRCzeDFfqIaYrZzr65R5UZTYXrXS4HjKRumiemI33ZdiK28z2M0J
jheDa8029SGUDR5u2diay0oRmdVPov+x0Tw8l6r4YupMimFkiPYjY5BCRqzEhNSs
NKoYERHGunGKiHyZ+qv4wTu5z1e2D3xuZChCqBaLuxVHpvjlYpl2UEYLY8U0+HKn
LpmVbmPfJ6DNmk0kcVpAWwBvS3E8WLLCZUFarOF5UK0ryDLlTz0+00fMzuEAvPOF
W5eWpBK75XsOJfqZzJmEx4gj33HS4SqBv5zMcr/kpCq5joxD5LSkJH5o2SgRO2Um
mxwz6YjLBgTVCTUZZ88jdQl1KLI2WCQw//IyPrZPsoLTC1Tv2LArZEU2IZ7nxqH+
l08ELLJpTg7qvmBFgUWNMbgUdQaLnRS7QXMqXx3exCusTdCxfqmg4U37oYt8nFj6
RXX8w2+PQQZ9HE1Ghc2cY7dAwy+45tmXVQcw4gxXr//FEVNfv1UwQ1mLN4D0v+OA
OqSUNymX9/M43igHtk1aTOWo72T0LOtP/I5R9M87sYhpr/g+ZtMf4lVbpiuSkAvQ
Dlc2JDWUeBrr8dtUxjzLOcwOwXWMZnOtmse2IjQ7kmOO9c/QgGrvqMEUpH8JiQFS
Qk+BFU6A4rDq4vU/hZsqtcCiA6pptKuBMBIagSXbtq8cH1GpZAlqhqmrjdRfvZii
C+n8qR7G7biQZbBJKVg4YGV69q4gOdTtSX7oyHelwYCyn/fxnMUQbeKKRdD6DsR0
P8X0N7lHn72RAlW+OO0IrUDo3qAbWoCB4ew2rxtCW43Dwi3mpiQf/CpUzjPnuoxH
n9wbb0Rb359VgCXHFrDPMZ7CNp6m0o70zGZloI6+s8Eb6LbUjzvqBGRJ3fVqOyMT
mUct9lLP/5qFRd1eTmB3H9PMWGkumXi8WqkJ38nqoyLWh9Xx9A1RBM1HWGU9j3xL
l9JZHlNkorxuruDerBoYwYnAd3ky54FpGl8UxB622zKb5VUKtaUS4oHctj92PVg1
PPRhe5DU0DrXyuugJviCIa5ST9Z+o7L4CGpAWO6cf6uTtLW2dDvhvL+YdWXdW64i
qRTbrE8dXM1sTk1c1eM++3Cw4JV3KWl6pFapHS+yYXbbTi/u9REACn9PUGhOL2KO
+a1YnD8TmCWQQ+eL5Q5TK11zxP2xrMtXMQhGpxyUT2oJkFhCropBZu3D5XhyLrXL
iMCxSJCTOmhD63ZmNSdEBkLsuZNCiQpClgl5Yewei0LezL4Fjr3TVELvmD1AVNcm
HCW6CDImHCQyg0u3cGjtoh0qAmyaP/Ffu6Jhfh6Ec5Sgc/fjicpqSlIhvRkcI6ef
RK8y1dga9uTLVD8TzIbnFC20qFgpJ9joFYGnaFWMdvuD5gQ3P5TALomPo33dbFeS
ztdNaJ5SJGaG7w/UDZtciOIzfU7c3VjGfuKx7ezH5j2+DQg7E5sqQ28l28M7IqD7
9KI0O2XEj1VKwejCCK1XrpSujEWRDdAISwVdYVVKxz5HAKZ1ZMfLSYX3Gy1Se3iR
2HvQT0gLVItPer9oJ964iMomSU4qELrP/anZRwLjclEur37dKDEBJUChx1wCTg/4
DCPsCTP8BxPZf4z/q17XIQXeKYr/UCZYUNfhBHS0F5zVTcuX2TnvNHZLo0QXj1ha
r039PO2ZGABsZgKZMB8RjIsaGmomiJMGPhs8nraCaUjC9KJFmnyphpa3Fvldm4tI
63GbAIhJYEQyQzs2L/zjsBNMC4wPjTpHaj5KpOPaIWJvzJEenzC764PZE8PoXz4d
0GOzAyjuKOi+EyuJ8ztL4Fb+WIjRICL5jvmYVKFveIhXuAOEe2OilrhaKENHkp6g
go7fKGtEXuXXaea8XKr1pxq8OuN9j+w3My2KNr6lPSXAA4igLCRZX8TWw7I3fngz
XmQ+qJ5YZTn8Vrk8tX0DwKFjp14dKG0zgKp0E1L+ssolqeq26sf2LVw2ClQpv5YI
1L2xXnEng/Lrqdot8FoWhchi7HYAjKmSK9USJZUE3Xhwl8QDBb/onynnqIBmYQXk
DRalK+ZUu/FGXVuHTVX3t/LR7A6HuKYYVtADW+R/alYOPk9ugLh0SjLtajM6iMud
vYS6FG03aUN1X+Gf3gEby2J25YwjG8eqhz6KakiEM5l237kAWhLvPjjQ3MWLl2Nq
wsDBaYBbotSeC2SB0qf6jZi0cHO9Ca1dN2c07dgBHzD2GG87R0ymAaoKRlJo2lut
4D2L9kGIxTXVQT61jyAtnow6twdGZsZ2lvKsRzMsV5NWZoO5Mc3onmP8C+Tescjz
UzpqJbAgjnu5WL905NDON2l1m+aR7ZGTH6ubvTjsnLvqE+uoh/VMzi733G0Rhgi1
Hl+0cZc75dW3+nJtXPAsUMsVcm476tdIiTdhsCUKV3wdj6zqTTus2/lKC1CmPge+
MuYVUxvNseOqwc28pG4VGGmgRYlmb3LVLgEpSAZ1bqgjMTK1zHW1kXiKNWjMvR2j
lcGl7titykFI26HUBu0g1ApeO6HW3LASttLiXgVQG5zwiIPhaPnhX7qGUgu5sF2n
wzn1ZMEvJ2MKoY/R54QBLpw4ipMYMcNDxit9hNZYGW5j5S2wL2QVlwQo9/JeN0m7
sBumKVT4TS6bOQWja+MDjTrqbcDRsjj13aFhqGfIXqGKqbb7v9UJPr1LD2OsJjYm
kwwdGuz0UcbKtc3NLX6/3YRuxvmznx89sTxYvWSfIgsj9HOlRaMXqmcrzOSeawwz
SB+bw/72nLBaVR8v7yLHpQhCDxgvchQ04ltsW+omxesHYuQhAKytOJmWE4T0IIyf
KARNJr9s3CTkq9alrlzXmPBe8OQdePhEGMvZGfCHguzvGDJZjbEdTMFHq6pfnJGw
3wbSZWmW2i0R+nNdKlNPFZTkpfxuWPy1D7jOv0r3YAKXSmUY59P+eegTTKnfOuJJ
1ZWzDuXO+omepu1DcJ4TriqZwGemuB8uquXhYbviQh6BC5NwJDKcg2aPv74PcjsB
I995G2EBg1hLsyIOIGBY3ZlVKaETFYq+JZdA/Cr/plbgY54V6ve6qAlcldXTWV6W
/LV17+rbX6V4Zy4dEdktTufm9krZbLF5kBB9GNMRzA9Q8V0HqZFxfhhh4BAJzz/j
Drz8l97pt7ZJNwlAqMclVixl9iY8XegB9FVOncOiTNVk/5mqW0UjexH2t3KtLHtR
FIJ2BO+f/Af+dO8B/vyXcoBAP6TjAGJ0qEVxggCviS+hd0hHHYeBOqahsom4uFTC
F4DNthDIe+nmFPNN4v1xIMHHLmkL8bXCqFdZMj2OXvYChtDJased/eP1axI5s0T8
nibj17IxysOas1hWqAqs7uTxap3Xsdakkk8HnY+Q81AEnvimNxht6viKU0lHjcKM
XU4CtAaHYNGMHSNG8IkskRx/Qs7vncAeC45D2AyUmZtfgwpwQWvQEnHb8eZ5AGrq
VptOiAYxxrR93leQrEhgLUVbZINzOs6qn+jbR6e8eYFtT4SqcsFaTvZiixoA5rse
ghV2REA7OqB2C2gx/USumQ/N0nb/3yv972XJ9wAEczkT/Cd7vlggEj2PM3m+qAhl
A5iQ4qWRczcP83jVIYm7OfutSruUyL2QMa8qewJrBIsAzCdA+Gquf3XHkIpmkO7K
V65JACRoLHFtphZH7YNTpUm5ozRO6VHUCRkF9Rqiq955ZHi/dB84APz8msl3O4OZ
aFXFkoGb3f+NAXvVKcYObibfyYbRfVae91a7KnzZrtPdtU6n85pim4Kyoa9nGK1w
uvQyMWTGdH9A5b89L9FzZYjs04BjNm9bvuv+2t8cIR3H9GeMOnNHDkw/DUFQjRcp
Nge3KVJSdRxUPWfP3mzHUt1R60YGBjCx8NIFIoTmliVFTXhY3GwV9eBn442ZbMAk
WvF62Rf2c211kZ7uD9b/1k6rEAqY0UFn4geVIcl/+ffzB9MucMJAJPTwgywSE5DA
TnG4RFZdGDfPIHV8iRss35Ne5Ch6C7VWNw/QLAuVi1uQn6FRtgFevmnjWnamEMEK
A8AGZHI77zaiJVkO7vmpBRz4pq4FkK3hl7YjjRX9y3/7sWc3JZpUNFJ7FntRkRfO
UKHCquceNv5V59v7+Cri9Ex70SVrgtmUz5YH4RJbMKLfaKJK6jUVNnUtOBGkfq52
fHNijNrdmVie1sVNGasqRl1gF6KBk/R0OXbyaDNKuXPsOV0CAljuAvMi5CfUAMsX
l5zexHCof7NbQvSg23Kj/5yQH9v31n5SFvg7HFJZ7o7H8WYFCgy53Q2EGZYmsFDP
dd6RLemKU5KQBi19HL9EyCXKfk7LkNtAkZU2IgLWKhcM6rGSHnqur57HBuXJLE7f
gASrT+Xam/U9zUnWPm9Z0/DTEijSJrHS9kvwOsqeB+yM1YFLmx8+VwjqA8atyVB3
9N5hW7uIHDhlFsLSEEhJebDpkY0pY425hn8e29ChjOGWd4GK2LFWXkWJc7/JXY6q
+OLovD3fHxJ8/Tq27bFcuAK11VFuYlDPgJcHAFuOB2lmak0dtBU1tQZqDFdA1m5Z
/nLcYd3eBtDeZsFVaLPiQtabuiGJ9zHjR/Gils3UaC6KyWmjQGv9JVfvsWcvykWs
T6Io7RE8hKKTTXbrnz3H1UYueQfL5uWNnOlCr7S3sdhDzl8qjuHnlJYlgiUHOitP
/tdFAFiSwR9aUeuj3+/++bAU4iOnb4zUpWZJIcR062T2a9eQ2ImHpKqZuNl6P6WX
KSPPR8ELV1NKH1RfL+kB/+l0ZTAODNhuHesdMHABiM0e1OdigSEYrOXkNdAchSri
EzUNBngWly0v3ha0qjth3hfa3TPiuEkQWocihHdi7WRqTC7d9lxadfYuK6lUkq+B
UnTD3O65qj2BiDkQLBkLA7MqAEjjqvFy6NB2QRQTDyaVN8oyoMlPE6YaLDJPsaur
y3hM0zjlYwf2LcDHko/HHPXTnb99tR5jasHUX6fbokm1snsGoeAO0BwxN4dnDAT9
fAFk+Jzdst4lk1NCW6301pAkrQWONa9a3FTD5BtYZPlLPwBAIjWGnzyOSjKdiMkg
qLMx28qvfIR/k1UuC8Yyp4QgB38MyvfaGkMoy3UjiQOIIZUjewtg5IfFvfmHBt4D
bmnY+0mTT035AH5s5wshUzC7ObgAKsr6xoJOspy6jY11xXw5a9Bb4U681KwZQEtP
Nn00XEJzPxmAJzPKY/84Qf6mIEV115HCEq6Ww4ATtMx6iYlwup+unGM2XuAiIrzW
fm4tnI9Tjm4P6EI5c5tq5h14rQgI4uOTjJEVB/eqhiUJAvB7Eq4p96XTlNhMQcKl
Y11e4Uq3OkypMDzLh26KVkVvfLZrSVKpPbd9jBw4K4Ee7eK7UTpQc4QOpcZn/Vny
Ce644maLc4KSzNh2U77VCDZac1Gm3rZkOOwpXRgtUevz/veQ0c9TSMNzZBNgEaq8
mhYXGZmpUxKg6lk/SuGfURNy87mwG0vfEgRUEMjHYssGTZjPm/UVO9TWGsKrEPZH
6Z5Jkz2suFnVfMwpYFN37g7HDSdBI3tvy34QLypmPYhXkst6/WGMJ6+YBoAuWtI6
1RbCwwowYQM0XlE/ab0/c8ngJfWoOMS1C75FRX7gZF9xIJb2sYoCLXfWccrPWlZ2
spo7RPNVPN5CbFEJiOUVc10tTRzWiBFW7MsR7NI62DLWjXU2kaEhCMSnQHjKnUY5
5KDfd2hcKu7VvpBZzvj0vUKFgv1X8Px7MnjvlkXlPrnIocWDv/KbD1I3eF/KVIgd
gfHkAF50eQ3kPQFaWSTnAPZfvuHbK4RmeM/FIMMbd22UyplxXFVnmHyhGsC/nmwE
YdQB5BNpJMNc1giq/wtg6nA9qhTVbZ406+WhHKroo7WrdcCtNBkCQMq9O5jTuusr
mCTXTxNGYaJ1mt0qMoNC5pkrsSn37BZlqQ6afGhdDDW5Zg7pbSllIxt7PJqvQ4mV
buABZF58thfXWdWzJDu8RSmNzbaNJdILhKx1tldR53d5/m1/4zcMcvzdsGYH7hze
wWbAXSruL7JcwMSkO0MsIhW/1ck7s3Qepshc3OWxeDBr8jXHajAelNmzIJB0Yqt4
CiWV4pOo4vZZCZ3lEmZwAd7PEHL56QYZ9lZy/lCgPOif0mYG9wu8Eeh2sptbeBb2
VLTyUlq1AkGalrRC8BWyv39celL66cn1ep+hJgTdBX4soB3ip56B4tUGzGQbv3EE
dNUGbUdnDMH+PTqlYqfRh0xF5AHTe+pFG0umQzmf2oM9xmNfJsVx5J/+7XkuTtBT
DTajjINg1qvtbUndlHo24rPWYRuhuO9p0kBCJx+YAYMo9XysZETUmbSWlJUqOv5j
0yheasf6jnFFRAavKVWNM4pE1gIdKobc0ost89Mep1o+cbMwsNvREXGjpXz56/0g
QisQcN6HIU0ZW2pgLdEiAT/Bt3noMLaDu/TgPFHYo7dScpkGRUy70n8m7PBaAyjt
fxPJ66POJfpRCgOy5UYt86gJpl3bmdO/gLzLGI/TRyz5uG49oFzFjyagUIJBYOhJ
6K8Nir2/TNM6eSZ9GQOJLT5jtQJMTW3skI3ghqawOU60cDrIqIVwDMw82tVJXyga
k0kzh6003t9HVn2yZh+q4e16AQeGpaBoHM11RdL2XqXjE8EDpbbeh67nzOiLFw8P
VDQudle9CVURYzdlgBl4dpPfZpcNOr5ymGdm8wVOptr8zVT+1bORJpG1RqIubc9O
oRZa9PQ8L0/o0Y3f29C+lpI9u+viQLMOQcY7Lg5z+M7peD0+l2ddcESL8Dq0Y7+Z
OHxTGTAQ4I1Z6IpNwVdh/FDzGhWxatterF7aeg+9Hxe7JYKMNeM/IibyArnYOOCi
CoadUPSVr/aEhyPzFIyBW1S/HzHL1Z/5rrwH8mZhY3ewNZXCm9qJOK95ns7Epu4v
nT/Cs+tDROkejDI/A95wL87yxecp8Gsc9uTQigzufrjF9k0b5YKS95qFGpAppKtL
QmhJEnZVdF8yGhdrNOijSTiRuQ8bEb33w07CDLAlIlvY7aHS2lW0nrMQ/n3kLh0c
UEO0MGgxTB/mgPS7cLZDgWs0AniVEdk4NDmbfITxEEh7Bnu1duZUOGv0HVUwWnF6
VqbxrrSpw4e25TlssxXGAu3JmW2eGLlwOKUZLAocjv1Axq81dkbYA0ZGxQogk/O3
s5F00+upJWyaLLuoObrmdzT5oc0QbDYetwAbvaTAbANSlp8LKG19Vnk2yjuoXeWQ
nAf2FxbuIc/rBAGRf+5UvAvNX6p0pJhE10rjYnGH3SbIp8MZxXUSvrx7WskTH5zX
iBV8O9Agx2FL/X+tSJqNu8xXEfodkT6ixTavmAgJmwr0nrNwdOSMMl55+Jpq5Z8T
A2TVPAj6gh327NGb01UkekuVvPBqv/vc3sSxfGp4dsODOdJJL/x0s0D7pV1so/fb
ANlfFSaJqMdbrjW0v0q7SenQDyZB8Df/XR4+1qS1idiD5CqusKIK09nsVugmeFEF
klKtVI3wGqmlzBaxbilWdPNQWOg3R8Cj9yV1P8LlVO+y6kXy9/WTGeH75uMwbHHK
HesDD5VUDY5rvzaXlaf2peVQk5n1m4QbSG7BpwzWo75XpqeYsj/uA4PwM3MzFyJD
V9wAk8YjVrXRUJmWYxRs5KfHdEaRheB04LC9Eq0Q/v9Qtb1HoMx+IaZ62SvgFe88
RD/FwnlyHxYSdozV8Zc7Vxx+GiSsulOIR2rH6e7Mf8VA7/Y2eHNqBAKLgwxMp3il
SczWIshuiYZ6URth7TcMXmpVcq0farqcwL9aVBYz5JmCkBwG8Zpceb05lpwhGVxZ
88/9LZ9c6onH/+Cy2YYNPU+sDkEK39kcw3RHquM09Doy1qX+bfRiSl8QDgM2Dc7k
FzR/yxlwNtLnvp01WjQkrnzD3PBNY8xG+E2WwcbCMtVq/Jlmlo97DfagARV54Hwm
Ef2StLSzkTtS1xUw8PGi5K9RwC3ihGfqRzGLiGlcTkT57Hgpvy3/A0Q4zSuD/wVs
lp3yYlKUQc6lbaoZueWgBn7Jv4pjcS27qG3N2Q9gSvRYYBqN1hHKlIGQDrY9FGBc
mG2edH8mZ50KYvYrU6UZ447oPPWP17N7lqb99xKlVv2VwRDEMamqo1RGY/38kg8/
Pi+VwAsCgNOKGHhGuD94gVNRstvLo+TesEfdpjJw3yg5b5S6Bx6mZf0vnnT/juiT
/CpQDfEiw9C8PQmc+uS33LvFeWKd8N0hGXL6Mg0pdgPG8ziRosZWnIgF0vaT1A8z
RC5Ds4AuTQRYC3MgnyWNA7MBLMhT4dR/BN1NtidBlOC8Yuzrf7l3yY1yLW+eKky6
EnJX/IZyzGofi3LNon3WJR66di93rbyJErDEdht2G/xvV6KpE3fzV5Rjjgjb3gi/
DHL2DWcnQGBRVzSW9kELGzoApB27vRMieZJei+1pR7v2PCIihFwVjlKHlw4pW8He
3GD+/EzkPHrk2eIyF1Hl8SuYWbgeqqohpsMjypj8gtW4S7p4uwikD9vAnpHo/WpK
7KDpCR1HVhFAXRuJa98RIswbS72+1psMio++PcKK7hyd5X95wZ7cmTNWO+PLy3E7
sZR3/9uEbKjHVYKDd5SxtPK7xo2yRgWKctSYlMbR4pH0wY2ZtrtQWWr51ZNLP7Ao
xU1szhMNla0qXJSI/HlED8hAAHXPhP4tUZXBfMEc5VIxrberrGxBIzb9cyOE6t72
OO12+BrYjdGwbOga+ypxOqyDamxzEDDFLhB0xhqTLtp5kcvynpsgBKKuzWd3Ym7A
5+FqnBgnB7V5M1JpIzXTnrXq6EEggAM5U3TgAG7GStXwExFeDl+bTxr7wXzcTtRn
NtnOxVGPOL5PXUgfG/BrubzXmTJqfk5UW3IsMMu/pS6ZJxLD92Viz61JHrzMhQNZ
D0AYTmu272P6mReTkYYcs/wx4vGzNbYl5O6UnyAdz2mC95Tb6ONU3R4TRzjjlJsz
LrDQFMtxMkEcOyfJWpUgZlVQagG2158A4I1BjWFHtJAVrSvCeVmj0/7aaP8G5uBH
Ix9wG+afA5+w5bLsaUa5tyzWt0ld427oh0EUGl9RU1OiR51svmNiD3hEbvL/geOy
bMkc4vGglLv+Ef5/A6qAhN6yYgVlVYVHIrILuEB/f0JGNxO4kcVHhHT3lve3KBD6
MiHJF4jLenxkkxAbNS3YHN77OH+TgI5ZC7xbf06lOHqHFII95t6llJukTm4RLIrG
jLax1xeWx/PzF7XHH48IV2Xygl7JSSaB2j6DDjlNSIQ5+BgOUvp7tiKia+gMQ6rR
XmnJl1aR1+iPfnVxMv7v2lSTeuSP8Y4ik0jbWmHIuUY3dOcVrZl50fUcSkDMy+2X
76IcyUxCZKtWo2TFHiWoklUiCHPPc6hM2iV67iwxZe09uAlqoBlAd7rcH8m769L1
fO0tCF4DXXFonCRb+hMVA8dLn6psZr1sBng1pqncY2iWSE5rGNge5d4Lh9KdnItm
ugibF19xt70dtujGQqH4Pysp8wVA3r7z7h9ftQxs9pkEPvj8tHAukN3v0TUemSe3
vaLCAIBiramYyFmeHDIiWdbbLkvhcgA/JvIwd+AAxsk86Ob+33ZQhWGFdz9cwU9j
IU2m75i7pQCLW1F0+XyYQlOOIAkPsLMVIJWTM5cEd2fgPbrUUsAMlzecVe189gSV
UsVTauDfU13nHUiioL7avoOFGwmJS/n4e1ALQzVXK4LrAPOzcLzJfWVJW9IZwEBF
iGQXurgDj4b08vgHU2pSfqAkfPxYpHt6+25NM9/V8aHv09K6/2teJ/aM0PI+wbVU
uHr6WqjJtH1tcnZMu1u8lJR8vgDCyPTZqB0M+9kO/4x2vp86qIHjSR0ly8MYkMUu
Hf0u8UPecB9PBNzeeYQQAgO3aKqX3FVkbGJWqmIEMxwFN4jAKpMPZaiaaTj1rYBl
5JwBLqmgJ+O4FxLNQyFYYZBvHSJf8eitTDDjiGYgJhKERjxd7TBsMdHmd7EgqBay
GG4/qvlwXSWHUhqSs3a3yEg2nHPlYfsCJKGoH8lHCQ6qdJwyc/cD7SNqgRZ1Rwel
NnoR2DcL8NtFOCjhVHb4PIcibTwLZtmSFA2fX7e1afyCjv3V57nLj8fpy4v87aPW
gFRZIzBM/0vVTaeLqZT1ygRidXaunrSvgKZ78uvuC8cRaIGs5rwb40EsqwkvSTNi
rBObyWbHIebhFcyeGpc7vQIA+eV6g1FttxT4M8enCas3BBtEzLhTxcQ5IsamcdmY
ZuU5/wFCYonyVipqUhXTm0SyNT0YcejqDmpO14IMp2YPMRtAp1jhRObrEC53BaQH
hX3dmjwdTcC5fY+Zj3VCeQmUeizOTy32eNsOg/WOSykqmu7FfAfdeLos2ZaQAoFw
iLHUbhMKamIEr03XzxEbNYUkfG4KzIEG4aCsMNoqLFmvZH4Vm6ye3RpEjjRnVaCT
Urww2o/sV+/uYQucHaSnKLplCAgH66gBlWd2D2nA4mS5ppPi9QcwZ1Zqkfl7kP0V
JAnCBLoy9rz7fJja8jKmrRmSwPGcB/rLmU3RTS1SL6/YB1WW9QGXp+aJuEtF6uwM
3JURKTHg4AfVAV1L5RkMhlrMpwubbABcu5LYYIAnD/tZ4zZ4vmemdt7IqKu1hffs
4TwStEm/y9jmTYF+HsszfCpyVwaREhRdQnFJHB2wijmQwqwKs5ROD4QX+amrokkW
4LgmSFG/dGoRhLLoITT8crWNtMg/oEwH8GSboXbyj7DpVJM6OsaG51ZdoJVYe6Yj
CBMjpLRYcol+v0WhU/W9oH1IMvFZey7WrTkhp3oQ02pfuDSvxYVs6J7RRYX9LYfE
V44JTX6IEAwCvFcflHiWkfIYRYG9T0ngt5NWZlIn3nZABKMTOV1/Ow7H019TvCmm
fxceauwcRAf/t203fKNHiaf22ugBwUDxBdKcWe6nEzCfVVe7TWIqJIrLqUj8NJgw
GZaMs82691ZKeeW9yzlFL1Fm9GHm6QFUB0PPkkceTUAq65nyN4gCLhBlCapjDGMB
7hxPKuO8WpP16mYiRnrUGwVOenOKKQQidiCQMo3CV4RLwXJoJ9JbwOOWROjOjf9E
1yXGZZsjCovOwVsaJQigFAmp5v29+24mjGfhc6xW3BPBAc9jIth/nQQOPKulWz/u
pFxGv7HgjpVvlbLPUPHDmGek/q/zcAFju+db4gPsOUj9qulndCxxEBpVE6Qyqy2G
h6BZVjq7y9t/ZHPoMYMO9mg6cxq4AWqLI07fCpG1qTFYgcjPW11H90I/ZuarqlmA
mQmwZa3XyV1WXlFYoXtE5YX7xbRPmM+tMFuCYirytAdJ/VQ636M0jZlItxWWJE6P
8Bh1+J5kP7GEe3dKpAHHd9pfkpOzwveTQ3XmMYSvV8Rd5R+uLWBW85a+clXpI/oJ
Xl9RvZXiDTShO/NH8jLV5id8WUYO8S0ggXDNZby6SNEftPqgABwOvuJObB5IjxUT
8twHmtETYrcbxCL7GLEWzpIJ+RDK2sQydnwqAjXu9K31E0wPYq9WdH4drVEiiiEG
NMjqiuZhX1WUD/4RBuXfFTKleRpsJQjxXjt+ISx8BZoqkPkvjdDINYKz3/mwgdZ2
wv+3Pk1v8qsVd//tNGT4h2J1q4Fq+18q4DQHlmeVcTbZ5jh9wbenz1L/j+WVHeQl
nx4F7d9cCADEoj8Gfa7NI88QgON4zXTdN/8I0aqjpQIrgrERx+ZwlvKhNUlvtQsQ
IrmSb+G+6ctHrqxD/BxFu7HL0o59ZXR4dtv84SzAyjTOELftWujErNaIFSlHsTKh
7QgnNQn88ENwuVpeYHg3eTFAqA3iG7BbRR2O9SdvmjCCxNdrc1jHcIY7EVq47ZHp
iKl/BpxU5xMP6dgsTUZTW0NXkyROVQ4dgpQ6iFBKgc/h2nrH3VK32oTftl1how2g
bamhzVGpq1lC75mccnYpQk3TPXxyiCXCP/CRI1OyGHY3KlgHcJ8sQzHhqc/6zgRs
CKyxVZiqPO9TnhW5nXu9FkRjV/xydDlB1Z0XJX9ujrxDhwx2L31+uBgCFP72V/F3
7M0lXguCAE0V7sYXQEVcLi2B9+x/ON5gYTR/kTcoiUGtPn86w9u26IlfuZyAuxRL
I3pfMX51MX2wGYtinPSX/ObbpDXBZlJ1jXuaTpdKnrRN+O14eguVstczi7ZbTzt4
5bkdw5LP6vMx6H0m8isAqQSTtbHYj3ktdK1BbBvzKGIeDWnJ/np149RnlKXrSZ3K
UQYHiBvlGo6PkXtmkzfqdAawwN1WI+1ZptZjRC85x5QJ4+L9mSOGwRnbXhax93qK
LJs2V8ZFrv81KSYtFvu2yDFYyDrt2oOUOnBbBWYTzPcaU10cH79aK8bix1JaUo31
Jj6/y1NWLhEbEqs45dszqdujnrDbqI9loDwKmimpaf6AWHm4CYvTE8vRNqmHEDxr
Kur/VgZfn8VYmloJK9qeS/PJ1DeIdIXQqqtgzaGxama9qaP0yZfZZQF0kphdh6Ad
4d0S6g1iRo0PNX/dLfmWTjlynvsXvoLrd1J5kvmy8BsC4FzxGk1W4CtO2w/8y0ek
qoFDTRaeaSu7m3shjd9eNDJP88Fqo4uj4fQJ+O18jZAkbRlhOFk+Y9264UkArpDz
kEV/qxybhwVmSJlsEIwigOt3a+qJoo6y/F5Oa+OwlofKvTchsznkA17b8rqaZ/72
6hjpS3bO1Ch04YbI31Cjj8Jn10Ft1L+tZkd4o8lF1stfhlliO66GvxuBZsEcRoru
QqEOHXR46pM4RPC4MMQimOYsv0Gd0kOlXj/9rqB+vTESUJXhuf5a7EoOnSjIWvpj
p24/xOy/YXFKfzOMlvU+ExEeYv+tIl3lzJqjn0F5FJTswBMPPwxK1unvDXwZv6EK
6w30jUaaSH1KSCb7UKK/GHMT23Djh2dwSc0oXNCFU6JQIDt33I2xPTMs24P/3ACN
YhiFB3ofA4WlfedV3QKjIHj+iQMCcF8jh2ZxJIFVHdkZpfkpOziZW+jRdY1eE2Kc
0vRHDasxmJWXFiHs7nMgr8mEuZG4q+BsTShL3yzelFl1v5fV/qMLdOCf7f/yl/sA
9Ft1TLKRPCUZ176p7+kLXX4cbpKNYyR/Ar+bAPMYDFvV8PKtER4i7Zy5HhC14Ksy
DcYV+WtShgKJL3uGBdZvTCKXabHcNAoFoeD0TV2HdALJP7z0vTKetZLufKuu2IQz
DKMNrY25RyHOlxUIeliX5evAtOakgwcfdXck7g6nIlNR7s6+5e3mxfj0P1R2gF7g
MXIBtSkGzREoQqHZ36aWFi7sABBcV9J0o1xH4PRwuEO7BBocohR3SQZlQ4SCdTh7
bjZOZOtb9C3J+2dGNx3BLYFLdUP3OqvI1xdfCus9PTwzIl6508jVI71xqkr3h5tl
vD6mWFLHb8DAYTnrz8S4KH7FbFOGErRlkwn+kQIqZHADbFcbLYZOxg2exPYgz5v0
YxjA3oAJhPvNeY9pwzK3GY5CnOJsf9Mzo5D3ue/xi1y3Q24WfovlYkXncAATlmWj
4jLAh/oREwomyN8Zeu7JQUuZkLHgX3elx5X9YrKUveXTDuVDzXfShHN0uF1FzdPs
DvMugBAhih4rRBC3JPEiWo0ujvSe3zBJvEfmz9ESEGZ+v80LER9weWltSiJYx3yO
2rOnrYWkHGbmaomGCT1n0dEKukSBQXmshlEwZInw4XnIWhv7Akyug+p6l1joVGH3
66kXDFe8s42nrB55SUb5H4bcRSoJqhlLf6u2YFdTsEUuM7aLRgioHAKRgUyc5urw
otC+UX7NUN+96sa2d1ynrN/+0pSQvMUl/QZ6hpD/VHFVjpGbIdEHJ9npMEJZ6AxW
kWtl3iJr/0B9n4+eKlpEcU+P7CX17xRb/dOhP92ORhLeRTTmUD2U3YtA2IfE9tjs
8OXmM999RzSirPrWq21+oMq/2aqTn0haQxbWU34/3+athVjiVWes6Mll7vLCyQWI
HSI1UpyBPMQIdmLxaJAVkphQNDf3KMfQZ/M/CJPbqwSzAcAfy6RC1TV9cfCqXnHy
4clM0064UEcaf7Fw9DtoMaoZHFSFogyTwAYlcaIH1LgrzE2MBDVpJ8vZ/egl5r/r
QKeUdel0vnYVxwHsMhDV/hNkBwVzfyqSt4vzV7TZs3kV60EttYGFDe4ln/j4BHvI
cXADE+CiZ9hAKWhqJlWyxn1EMTBDsrQqAQR60nzu92PzasoN2QiuUGAqExhiqOAm
QcujqGs4e/tf+vqw+q+6md8/BeTmILS3MAqQST9h9KAni55vt/wCqViwsBD9Ifos
x5c4mfpqTNG/thcAQ1wm4Eo6QI5JJky6KQ+6MMCAjpNBL9dWigH3g0XWcXbJ//Qo
zNeDTCbL0dseny6hHBuideYPsYVO3E/9hkLeaDM0ph0GWT7ORmov5FiXRZ1L5vIX
i6WXx0OwRG5q+QeAildrzYsEhqUSMb+dlAN4C+7aL+yUZt5+lI5+K4ERwc36zvEr
feQtiQUHfSg5cLLSfMxgUh5du+eHnIkRN00+w9m46Vc7qgA/KZ6P1XXFaHV0w4yg
skkBh4kVD0sbOoliScFDSpBivhK42oZDTo+Q+nLKJzFwNJY9ZWuQly93YqbO2Wqg
55MT9xAkmkaShGkP8ni+31jBVbJjnrkVQ+c/4U9Y/7d0N61BWu1pSDBabrLFEAop
EZY+H1FgY8mH21TBnaxr+p+2XGSqniezvBq7Sp4JV+vM9Mix/n3bdHrvNZoA6uPq
2sHy1APvDWTZkvGdbKE0aITc5eeIoEhQmbG4nMb1EHPQTgc9cZilwQQRZyEty9mY
YnjvIhDxpSbni0NISIhGWu+FS2LKOMry/HeO88WbedKAHsQWyYl98uB5WqmSG6TB
6o5e2JmrKqvkzpAgXsoBAL8WSGclMvn4rtVVsNThPKCBgy+AKdc9L6FFxsL2qa5A
uKeyxIckuH0m4zBRb24gXjNbtplVypVSi2hUHi1V4hhM5w7ZovXG+qJ4+i26S2ri
NtStYJjougvHYIzpVJRDqSW+wUqdHtcz4dZpOq3PmuUrw45FoUSae53GaBNjhZa3
dq43Qg+azQtClt91OeaahdR9Yx8XK3c1RkQvZ6pLPKAOcM6/oTD9nf9DAntyBC1x
y1Adbju5h/FEGxs19PhY7SlL612IB5+uHm1gf61pMaq8M463RML85sSlhuDv0AO6
3UtpNuGdm3/aQQypFK+ULOP1UK3so+U9cffXY1S2HRQVgpYCKI5jOmNgEqwAe6s1
MgfY2Y7RsEpPFz71lK+/1NQHMIh/Cl85rc23uduHUMnysyI30AZ/Ts/fsM80kkJn
DnTa4eAOrzw5w7NgdLK3IyO6N4GxQkHshRB0C+oe+kPCToeP4mQANvSk9osElps6
3NotTGkj5RmcF2l+e6YO6vXru2ApeTh1I1YmbQKERV2gEwqnLbqwass87VS+l8Ku
xdWhSq1lGIBmS80XHxEGY42hipXDa/mBwAobAnSUwx9ifOxLsLKmqDP1m/N0DfmT
QxpV0uAeQ4FKZNLURaVDytbfX+vzg8XniNeqNyX+hq2QlYR09b3QOdjzbsp7A1mD
hMS3uJlQkSKL1PnCjHokk9RsofwDtRj1ymNiWoZd7rUUvGTlspsRsz+2JSFPbEWk
eRP4Iy6PrEwTH86RaqsCN11XN6poqeREPVhmub8AKxTDE6G74scJGeyrSHoMYoAB
iIBEuhN6uTAoIgUQ9o+f0/0ZUn+botaungxXbn3GpA51W9aXFwA4R3RAyUbGNKwH
9tpHGV0AP6eL8G3DTm/koZDuIlPHvzRsaDsqd+xDx0tnOcY9FzcOjNp3dn3rm2Qp
oyej1UnxJuR0k0g5KXyq07yvE0EK/lbDw/SyOtVFd4uQYYwIg/MuESqg2pzPoMp0
E6yDBUlOKYe4bgMBs/f4kJxM1ItD83xZSnG41tixNLvrFvxlJOGhK1cJMow0aLnp
kYnrV5bB0UACyGpYSTNF4AJGkmtQLdZOB8qUMiIadCt0TK5nfFx0H8Rnc+jMkKp8
FQNZDXp2hbHXljVD8web0OS6EVhcOe0cM1SgjLqXECwAshuLP6V7zKkTzpmfo+UQ
5xg4FDbe1DrnQVER5KlBlzrC+0bDr2TwNLihV467XS0lqAsAv0YLMGYW2SPcMdAI
qOTadV8XYVHr/vZCLaoHBIvP1nABTf4T9el4lxiKdmKVL0Vh82eqSB2SFdUkr31O
2Jr6dAF5g4G4Zy5bbx0IfRlxaVFTEjBwNMCXlX9s6ocQI8EsQnx0TfcQoV1tROFS
FcaXFevQdD218mDOQQp598YY7hQNx/diQ10/ykUiBCZ5AnuL9JMlJTY1Q4OuO+dN
KzjUKdo664ZQvvo7nwA5chsFKmSAsLLEye8h6V3axeAagXLqRQg/e4jbVbxzaKEe
rzWe2nNOXglk03/3UR64h3E6SXQT3dzGTvZdfFhL/oCVngtZPHAlf5ALwdKO4ZQL
ISnz5NUSrSSF56xHk7o1F4De1o12UHaMlkz5NZ7P2b7JHNu1EBPp58mVdyYG8hgi
NScAszKP0hFtJOdpgwLiRnWb4l2bXRzvyAW5whcOnWYyFNQg9h2gSDFJI66ltBIS
G4+mZeY48Ln4IVJvXrJ6YjzJGp/trYbw+eZbzln8GdlGGFeL0oRMdtrhNnJZitli
AusBbC6P5gkSd8qWC8YrpN01xbKKVFcVM+y9I6EKT1T6J8gOjI8DhzeN2mIOWDtk
10paFAKp/BdrUtNUMCTaFMpqKhi2dgpfONk+XEstKEZD2zjQaXSM901BwFOJtdRS
eO0AIm3M0Lq3NlT43BSgWHcRdNyPRjhE64Cj5rzUxTgOzeLA0KtQA/aIbfGSFd5M
9R7jUR2fzkT9f/k/+A8ZS5WknbgS+yNEooobvkVTPdmKolPE8Rn2jo5ONNDOX5/p
58crRq//czHDvsBTHyL//X25mgmyLlfTn/G+OZH5ljZdvVzIw0XgFTq1boXhwQrB
v6Z48MkwWgDeB/bTqDW2QBh8juO6UC6wXgoyPa66QZCShd0D3qeZQItigGAgCzqh
9N+FfH0JkLOofowYZRK9kLQBOZEca1DI7HPfu2JOLYuvP+0DsuqwGqvsS1yAHDZ+
TSA+nsEarGdQdQATGR6scst3gxr6ju6StNSXB8FbjQat5gi99PtmdP8cNtx7SiqW
dl8Imy5ZOeEN8gD2Lm/PAVnGh2Oj1gmVlAIrZ9o9Hw+CLHJ3V6E5Xxe+Pf9pq0nj
B7jm+Vl/kgqfZU4QWe3qC0PxvKqkVjpevuv37D/iHJgzzbxDa8+8seRC2nqdxW6E
XBHXy10w/KZY59cNChImsieZpPkTfB5dlK9HGMV8J1ujRQK+dHdlv+RZBqBqEjiI
vte8vY0CiMs03S1nCtNsdV43qd5fz08ABPyNk1nUXTeOOerPS5zHjAXIHLP0Qj2g
s2VIWc+kKQx/X5YPISRSHSWEtiK4y461U+CcmN3hm9DUgGR90UZW28mItvFH1h+k
3ENMVttX0rTbty4f1uxCPLHxc8qI8V/jCEuHHlI2DLj76R4DQXd0kmnGQvy3XnEB
xnTjdHG34R4VjMCWE/XpXji+fGywRYII78i5BDGodLq1v9oDBx0oMFaOe4nL3MNQ
bJYsRfBilj3MGBFbbKDEuCLtjiejRhHQXjEJR0FTIygNZXVMJiIvhoGhad8s/Lkl
GD7iWDC14Ckod9uvMvnfmlaqYwBuMfCgAnsKaM+BXsLSbVcfeQGcwX6o/jzqchN5
Mb9qVhgHW9zCOY89I0FeuG/Fi3MWJ7dU08TaesegT0ftE9NoprlhLMeVbzZQKCHi
c9CYdj+xgzHCi7dy4tG4mMXvxvmybVxPSGRCpqOmv4xXxJ6bce9HN9BJaNiTLbnW
Nm2QDuldhVOOsjTpXIc5tFV4+qwm+JSIQLO26jMDD6j+IvKYrj3BjfLKB4a8KIO3
R8hX7b95t+4DT+uSaIBRuOU7/bBfGiLJDic3tD/RmKsX/vY9Gozbkr+L5iQoc+Q4
kglE5WBZAkuqLRwopyt1J2JcCIUx7uYYMMlVQXl2zvFpy8VJM1TPb/NfYKiAv5eD
AGcioCBR+TpIu7+FFn1EPE027GnsS5luIWc9mxbWxT61vu2Z6N3I8vLNb5EuyQzh
o/mlWpd4SoALufV2iPfaZYRsIHfPlm1Teoah6XJjrh3oJ0K1mJJT+F0dWqRRcDO3
PiMvepSRbUM6EJ4RvhrfxJ4ejk53WOLHlsK7WyGHjBFGOg8YgOkH1Ik8T3sWNc5P
IpkZZKwN+V//w+SzTBdhHrCs93v05d385g88tL81VW7qCc6XOHy6h12fysFT+9vq
VNXMveDrcOgzyVxEtsgLHidA8K1+5a+H+2I9sn81xIk8l8Q8OlHbbvVTgOaBusww
XV/rfxzFt/463gVY19Nf5YANvzSXKO8MvjvCK2axwEy+FRWovMjSuB+7Ly0H52bD
4KYMBpBmxnFzPYn4l4c/hr83rsqUWpDjjNf/NtxQKDxyye+W/bh61dh/5B4QvCYg
DDSsxyo/57JMzBGVMbqtUXOfZWEa/CwBk9o1guCtb9m2qRT2Jznu9xOSmHhtqF5y
u4OV0/xj8WQgXJQdFEy0hqkqCu3jlfMICmbQ9f6gq6CqBNRyCTDa6A3d+KfHVhmm
ipCtfVaxGaDgLJ1Lbh97EaJbTu6R8xpy4LUKmM5aufHqbADPHGwgNXskuGTw6SmP
SJrc0sI3ZPAPOs1DOLAFwg+4fVEOpsT9LI1yM2UODzUn2jIQqLJa4xdYB+ZzbkbF
Bm0bX5ybTAc7J8JIrc/+kkY4SDgG8frvs4rjDYPK0wlsyx/MfT659mU/FeG+TfCL
DoRorehZy9QU/6HlilQktf7+iWOp08NEIO1Sqzzq2DX9Y3aa/Zjfp7mPzjYfIVk1
N9OiNmuxNUOm1+cRRj39BBvRcj7IrmJMEC3B+xmFRTfixWTaFp2RYLhvAIIaWlOd
ahBm/Ha8aif3kCMv4rH3cnDHaYJu5iXP4quT7GElkgybQJ63AmjdqixS1CH1fLWD
JFuIqsC5EGNfXweq3fumuak0ccH3GsbYlLAVuN1axHn4Mcmw2qDbg/d8DB3ksFHQ
+ACw4CJSDb/K/dhMXJf11TY7Dvo5iS0NrW0oIBZD+AvL/HNKsZ5TIF+s4nQifnua
0VHxVY0wpPeWfU8vflvCMPaFZ/IvMKGfTP+XArqpI1mua+GRoL2Nld2XVhGleXPR
Ll8lOt9+i8AXP+6HuOG2UST86xKTvnVhjg58ROzo2TEUQM5UGSlvJwmAs12MrusW
ONPEqFcT1ANXVzvJS6k9hqqMyUh3dvcio5/+8guC2jJ9jXVXxgKUo6gbEqGPAyPe
/hBEJL72PvcYNJfeJ6P5yT59G7SdyC5iJfvCm9tjmVCM+v4V2vwBTifDjdKRy9TD
P9ZrmQQUZDfy34thNDINExIyT1mqPIUbnETGRIyT4KhxiXC4ZX5rBJ9XGW8uoqm4
9eojYZv6j7NGz1WEk+L8GYGbdYlh+1l8Pnja21I1M1jrPYNFbATOLjZSilZ5vPo0
oreYtkw1wrGrAmaEZ1lm19aBETASfN7+raT+Ty2HEtnO9vzqg2PEhjQiJJx/5EpO
bV1Ijggwi+4XOXmBosxqdmvnGK/r7d2pus5fcm0j+N5MpQM6ayyEHoW4ik9yV59D
c4FXJ27BNYyoQZwXx2USS4H0cvvfQF8ak5807WiPKwyW1lBODgPBba52AaZTF6we
9+2uPXeg214DVAvVHEzsF2bzjUIqjeaLGYDQTu6y/Oe+xVDP5GW5t3G0YVJN0WBE
0HBlkw0nG2/DeNxXFJpctoAH/sSrOD1r5CiBCNOcsEngmiDYL9iHUhktMIUri4j8
3J15sRPpkVco0Md88PpSZ2Co0We9NVNGS9eZI2qdUhEECf89/KrpM8j7Bmp3YabW
JcxIxBHY0XxvcxRaguV07Iew2Firo1H5htWY/Xz/Q0+vvEHeb+uHRJiugRAh+yyX
1823uVCh75vRKP6J7n3zrsSPPMSd9cIsL46nxYAzmFNbI9L4D/f5WIRgEQNZ/pbr
un3+YngNt07cVwJCwiMetHDPqGz5f1SF1maFi15lRN4MaDUd9ay26hGS561unsJs
HyaOfrCdBV8hHu9FSTBFpc2UoEcByxUP6hrbJpKkoSqFSgiI1ph7AU08+U/mr2ds
xxMq0jKwxD/lJjLRyEs+tkDwVzU02g9hvCbmztkerj2ai+VqDhK1S+eY2z5iPPFb
lBz8kDSsvhSbf4Em/GZqFvM4Zepd23HEzw/q6Rt4DxYs/gzGnZp9hUKXqZO7qb32
FAAKE8hz6nhWRv+XWSHbBHlFFY8VuZryYH1qUgt41sZ8mkGHrXINFemCe66LQpmv
GidcKdQ0+ew08zVRCZ2d91VgQ359eyOVJ/bftAUWXVId8M6Lm5dg8XKe2E/NHVQa
iHb66HRmfrzsv31E9VpMKlrYi3VcSr6X32q2efNnG9pRaVuSq6zx92AlDoy53d4Q
bVUNveGMY0EctunPIhaucNyLGv+VsNs6ldY/L3qCXjPTz7tEcIjPcVQZK1odwOaG
C4M+Puw1iBHQ3CxdnmFX9s85W+/E2AMGMXGNg/nQwiqXXc+5n0ycwxstWTXxXhzd
yU7xfYkZFO1jk8V6nEC8b3BXbwzOnRibLfeLXKDULY6gTf+6QuIBVlYV5WMTxIqW
5SJaTxKlfgxKe1tbjtI6MhpUnRMF+PZPDHpc/fSVSPxi6/qTL3EJf10LYPryEOib
IZoK7gkCnjeZz4NM8x5J5Zv41Zg9MKbE91KTPms0DldjETYGU+ku9wYXi7X1mnoR
gKPKx5aAXDY6H3QxdW5kK2kg6UxN6Pisw8eS9Z9fJvxheV/9J0otjSxAfElkpETA
HsF4lNLGmyLAws1XjSQSOChZbB53B69rsl4kRUWYm9KwSHi4frJIA/QHw5WZbQMz
Mjz61NSqFv+fszB3s6gKKTd6fbzjMVmmAkheZuL9mJZMAibbs6a63UNmvy36URJi
ISz3T1l0Aa8zBF7K2qirqh2YEu02IFnY30JspykjM0gEMltx1tphiOMzcMOeRSPO
9empL8xwnnzcWyT0rkqX44b2rdVWQxz6yhlTmwKLovaBkC5qAcXBY1igdoKQweZG
5nM28VbwNAd7/pGbkhnAcGIYJVZbCIhdQ15RzqpbpfFbJUyO1e+ieTB8+UWdKf4y
tTxeUANWL26eY8Gs9gTuExRnEU9mNkBNcvqA+J9h14CjlRTsWWU9uWCSTPVdxwfV
zrmeovNoLf8sHheITbNQmcQf5b+kGzHE7MWfv/1mMhlhegXHtcczM9HcIgAyBeCu
jw0OGcZJvlDa3XDKnClukllOLiE6s0JBMfFU8JLQMSDWM+7pPWFZu0yPsq5HAg/e
q0F9YpIOYjMPS4CuHirnqj5suAfjcJ/hOpXiuc8C02l/c6TQgqJ8yoNUd1SH+HcM
skOEd8ROhAk3oGT8+MfKBK59S37Ah9OcFlEl2wd3F9/EMVmvC2azRedtrhEacewi
bhS8FRfmXsQqBFZXQ2Pv3sGUWcTlrdHw7zpF4SJg8rRAKbM+gOKZ2GV4zeAw7hra
4HYVVbEFCeE8nM0CbiUE1BZ7OxkRQBaJd6BFMvfDOMptgMMMthgNmDvpYK2tX9aj
QD7rnsU+sy2apedAmhHqA/17SzwKkXrsySbfsDeQkAj6J4F8hiZ+ctro6tBH4EXY
PwaZH0CJYVOOdXJ7YPsVfIxpcshe5cADGRCYmV8JLmOvCc3viP7Lktb1vOxsIXZa
t5KLHYity2fwfj4gHX1uIE4CrPsJW3ju8ZZA08pJi1ctxOj6Izb+0cw8U0Jbh1dm
5OWAGuKvR0Cd1vR+viSCiTIr9+X7j5yt5lDcwZ4aQqA5U/VdfI6Qi4PsikL4BlZm
E3+uv1/wfxHboCyMyURGip+bPLQL7AYG3/5nqcYTTY1Is2gtnhUy4/pfHbN94/Zl
VWz5JlBWYcnLA/BAf2utfseRLV2GAz1FwNWt7CT1IzDx/fJEGWyUpSb5pd+wIHUa
O8aL7xpiTi/rc+xyOQWt1ZLRVluKrIxuSvfl6nrVhhNJYH/ofpSe3XgaMYe1VX1p
Rz1DtqOyV2HUHEfQ0SdgWYHNjj9DFA/VxjWVqggP134KF69DEoeQLXkl6NgfFcby
m3mGWhmSX3cPqLCwShKVm0D50xl1UzqKJaS95sZpd+/JIctsksVtGyaUoJKgorKt
/GVa7zyI/i4SogaUNGmNtAjPwt7pyeaxoTnrXA2lx3G7cpB+hQeM8NcMO3+K0u77
zmOGjjaNjFc2DxGAuJGSycVzSz2Ot3sv/+iqYJXbLyyt9c+pSXITUR2ooEpJ1I7Z
80qGj3ZGCFlOs9a8qQgOwiHuwtCQieqVdOR0He1vA2yQ6PaOouJ43ghJM7NCA7/f
pQJxNl0/piP5E18g2116MRnAYdto+eYfY/sCiYdbznVEGCl+jiPjXJP6Dkxhn6tb
KeT1ZsTwUeVXDeaKdBoewT+KFuPgfAInDYyw0ZWAJyaUDHdW7O0SdlTNZGjkKok5
+iLh+knA7U6kdRM+YeHp30Fw59cU62H0XQYKTuMKLAZAe5c1eDCA0YFx9IdY50w5
VyyogS8Tm0N29Aw0iRyzcHlaUamSgBAIMQleq24g5sfX3i6Xa8R5R66bT4yR+foM
Qy/ZWV7fhRXoHVcX0HmAnPoPbYcIm6Uhw2dgoOBYq0pmIWgoEzjGHyzAYn6Z6rRl
w/lifmdHfzIVqHMM9nF8SsysZ0g65iEcQXMN5xBCho2xe14yJ7RAXu9czYCzCdij
Xcqg2JY6IviRdgNm5fGJUdQPBVFyT3aicw6ztC7nKJ825Ce6wHDR0rphEnT8KVbu
lzrTUQrx4gjhy77W6o1GCKMKKzhg0E6VXR9xfpJQRGd6cESABUzRm54rrA1SVN7c
mDUIB+yYpEmLyaanF3hz4hXKLphWrZ4ke6BSDziJfgIe8N1F+wb1bZbsERqbKtIj
HjsICySUa5GJB18CeadkeAgNiTBA9QPDWV4gOJ7gQq5Q13yGCKOEVDFelktLvtWX
qKhm6VtShVXEt8/4c2x4gkzIalbSAyPm6g+88EYPvg9WxfVLEhVG1uGBgGRPjqOP
jVvpnWqoMzWKpVzka7y8O2YyI7KGXzmymDkjrYPsATP1vRZ3oQceHLWCS2RZx4EK
983/Qc4iEcACYq0FTUXK8uHfoooQPstTsSMIkepgp9ZWEiFIoxnz06YR4DVnRCrc
ifGKUYjsdjZNKc43npQklNXi+KZoQHt8rpU5i5D0qn6Sb6+IH7so9ZTe9npSjEkY
75a8tBn/XHRjBMloERzDUV7ke8hstMYukHArByJYvYTtuP7ZqM6eUgDqZM9uHoTq
rAxjOvDLP5qySvB+j+Zi/j1IACCRRHQES2YBhqpEDvOw5Ml3zyD+PT5pKGysTSpd
6nnJ+eb7zflhCXPgM2qGZ2INzvltjN0zIMdap2N4Nsslbc7KbvZ5fNx3OETysOpp
H4Rxp8uL01opOHlA+/GmD/wRQoUZEF9WYthlI01BmUEMXtetH5onQvnJ+OPiBiCn
O17jrI4u/UUhl6e8JcFgVw3mJw2E1df3esF9wc+H8SQhlBPyT9pM39+MEpxhHENv
uIRKVs0DKw7hDtK5NEo2QStCXyXNHAkmowmNJDtLAiOn2bq68QhkoJbUVAQCmBVx
PJ2t7AGXTUczT+nkiVjOu2hpFdJL/k16WeuLL8Qy/oRoco5Lp8qhw/VdAAQJ7DK2
OE7A5yaRMQQR1qeLAexwSqGVgNbvGgQrED5WyuTAA9gALhh9nu0XN/B4IW/su9LK
QWkyxYSE0DTL70JsBflk7nve7SbCllbkOoyww/yxgD/hMHgb2NGAyHl8GLv4DqeM
zp0uhxVUftxh18Lq3oWkmWT/Ktp9NMr4u6AqhefqX73POEVIQn4lAXnuIOC618zl
oGR+IPqY41/BK9XKiEYiUi9xJCUv0a2LC9vSlIITBRiuLSEOWIhGFIhq+zRd6m8x
IX9IpLLK3hvQ5TIG0wdFMKNH0cPW3Xi3+ZhEcgBkJZ3ls3s53G3aNLpmje2sffJL
9y5ZoVfOakoEtE3mzdItuguwNop0tR4Adq8YzoDGq92FtSMIUpn9UbrQX4T5suAB
bQCfbJw+dEsIc2nbPcGsZkF94kfPq3vIbLsbj18m06C+SbINVWiyFVWZaPBPHTuK
5raO2Qld8wCaV5Dh17ArYuaOXiKsE2Vba8NrVw65SX8ETVag10J7v/CZXugX9Lf3
wBG96rJyk/rYHO6Miyimmy7uwgx0t+5tQQ/j2av6d9oDM+SUy6ZGqUFsKbE37hjs
OzD9t5SR1pgIz8z5Ef3x3K9rJzQ/qgfFqDg927LCq1R9wW8biQjAJQgvyy6S1rMl
V8yqWcJBx5vKh0yISrBJ51gLlTUH8EOjS34VI6aIRKsNdB+Ygc5CENQfty7QAs/c
pnyEjUCyrvir6gFExdUsU6YaeqQWmbr5hQpx1Hr5YR/bXodfSUxLKw+CsvWe01PL
smOIPpPEwxtN8+ghXa3wugRnmSPEHzX2/GtGCNU7cISWksiMhIEuNOYpYtHZ3nxU
IgnqOLO2yhDkeSKEsFaWuiMZBB93oJhJsyI23HFcCcU8MI9cgQ7SSFpgjcCM4JiW
kUwXPjAQ16kNNVfmWVuukOXxsusU/u7dhXgjiMW3RWtAljjI9ud/V2P72iF/sJBO
P1zzKbWqz5kfxbW3n0146yVdTkVmwVWdxGUjzjBm0tXbZ74f+4g3DJI0FvxmdFS/
atmU5h5eyGbIT3+699KyNVkm5AIeKyzp2sM71Dxt5mWa/zTtERgmGBfybyqPvMAk
nHbpKKBoR4CSFcDIgpXi2X8cYdeTmh0uO418RAgPBvWkGcaj5iQlQyi+LN0XJ1Nm
nzQl1nBcSqKiBEYOa0ujbCx8B37G/YlKF+6vp1WNpdqvDagV7KbQsOqGMFA917EW
yB3WPGFsACVVNXOtmjpE84wp2Fs6JhhGDPgI3OmM6ysJYdzVED1MC5wRBePp1UPW
jxuTDLk21jSPLiVAsdsk+y1L2D60OrKGrpgghjDoXtmjqrlqmrnryIYfTycjcOAY
Ir9xz+WRIyDDYqy3wgNZYSPy/dNpckR4JMkcQBf2wf6V2K2DGWt2Omfkh6SVpGHD
RjJUmYjX8M0a5SNwiwqHeWcWiX/Oe4jy/pjX8fF+JjvxVazqjlQZ8GZ9QUd7NVkb
1Cx9ByulePtDzijRbcuzNsUw0+KcdccajB9R4kX+pSl0nWV7HjuxiTfgr9pyiONz
232d1vCr5qvyQwCOK6zePA0UL6UCgpKpaVHTQ2qDJmKUH4NFH0DI7613PJWNiK0h
zhlbHdc6dnuj6i36K3xO/rlCoeXlUJfrA/YE/7le9tUyl72hUUL/qXSsWjEGWYBG
7nJWfzScWK/MHwrRfITtwbjAIFrG0RxuJoWTvxlIR00uOM4vESaM9J1dhaWyZ1NB
zVL6ODzUyAA5N7tu3UWEY5+N0DYtjGWWRwGaAitAUXQ4SNTcjR63jpxhg36sUuw4
ZLK15L2BuPghoESgMtQfCWTHL8DK0ROYzp/6pqWkQ3wEXpEJNlcS9T7TwS5ABDLc
BWxrhdGCvjqmUWt71czVq5F9jcCuJ4ns7J4blgb1l9B6QFn3tq/8mFu/v5YPRXj2
zIm8hNqCjWYct7PArMaOc/V7H5rt4KHqscMxJ6zdNtejv4Su9O2ZpCUKdEh3mhHS
p1qTrnz+3JLm/ci4g3Yh7ADDJ7IqW/VjB01XboEXQOjqn2YgMz5v8nJsCApxm9N/
bPXapZaiCQ5T5J+iBZG2uXCvFTMhHTaLgBw73V9lp52vtoH4XPWR547JWYzJJ7Bv
b8safD416cncIgF+TE5s5CnoMOxSchOcJQBOE1xpxz3e0Rv7naxNiXwB83loJhnM
UTBOQ9HweuJ4rsiC8Kxv1yW7ywmcTNEwH1Qirn8NYYraKAYxQMAWAK+ipOfHUAaQ
7bEqBhhgK6wbqp1D0mx/UMnXiJJLIAN7g643uZisAbUP2nUK/CtFKgTh2bwEILxl
AujJgif48e/zVqbcTdx9sXUAG7+8y8yVv0IpvWQKb6/yCk1oo9rcfxDvsDBWzHyQ
UYFvGWBOQaR1VZjO00o6PmDxNHT8vfD7KcBEcazH0mtWCKB4WolsYklJdZQNHDmZ
ddTCZ+j6ia1KvsXGX8eRFoRz9VKM4Z9l1m0bGdlqhkOpHJ/p7I1/S5TsCOkYyTHk
ZwXJk2L/V56XMZFkMsbIpEK/bfWfatpMsja9iU3GywiWfIWwRX+9iefkyOYbz+XT
OyFyxd57PZxFvblN85XqiEhq35wCeB4WJTGLa72+vJw=
`protect end_protected