`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
gMcHP74wBZczB0bB0IzoP2xg5wC5NPjD/GsvSQ6VQgzYAsanETMwwsWi4yhFtJwv
5kY07u0WerSDf8woJ0stqW5xF501W3JLIS8KMiCOd55RHBOnavjYiaaLeu7oUCmB
TtTS1R4sO325rP2zOn9YwRbyyS5Ljn+PzFZZUmkt5xMca3p5NGqKtZW2dV6Babni
5HlLuF20Au601B75m2nv+ZRoGSrpkNElxoTibONmX8gBflpIVE7BehhHwaKSucEF
pp4QQ5zZAZjEC6aplZepouGVggAulz5AahlX5bf4opOVlB1J7IrgyjENtw6ysQ/q
DzybQ+ipztSXBGhmcCVU3A==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="jAI3OJE9Sh00Sic4PtM/KZ4WjwT98XM8AMZrZsQkxWQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hyw9IrFLPQsjvXplweG8O0lkaSLBN9Ijv4B5VdTRt6ipKJT9Kzsb5LxCKvkQyF9n
sGPOd5i74hRHnkHfYISGkfxGJCa55ieOyFShOsqTKRLxclm4oja9vTIey6yFm1BZ
54IDCG9h3PqfDiTD847UCSMRvFssyycwv+BRHQMQlFs=
`protect rights_digest_method = "sha256"
`protect end_toolblock="BnLuc3jxknmZOyxfJK70E5kp9u9O8IQ8cgkXv26kHA8="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 38064 )
`protect data_block
xABArkLxBOK6xG+7CdOOiGu0zbCbHMrEntFfAZEE/xRFxZaAZl1QLkuFI77OC2KL
XxG/mrHJzO3taVHgwRXNLDdc8ePbxbAiQfzV3NJLBO/OTJ0aBvTNnPgPVinF3K9F
vtTh7WTfQzQA1nIFlDFY/+gLU2ja9rmC8ys8aljkG1Z+sUCy6Q54jFzywaZ0VAGT
HxpuDb7YkSltFL7MgpuYmhLsyymk8gCXTt5+p9Gew8jaAB9sFdU7uOgahC+lUv9U
A8OS9MMu3i2npZfJ1F9bkLoCKDwP45s5xstRJFOYiNZHU0O6ck4L8i6bWwkZip6B
9M0Z2b1bhFc/NvL2YSYr4VsyYP+htFCkdoxxgFYy+wf+f5p1vZP3wA3vgwo+oOXQ
A/MY2tdLqg6dcJJEsUAqiw9g9FZa2OP4PQUjCijKmtAqW/25ESYqIxZa9819iKSg
Go52pPtRbh1ZTk8GoXo2bDtUSvxjh/vbTCn6xPVcQxZeoLf41NI/yCrUYAGQvDgy
QjXStzkmHmC6JxnNVlmuSGhfM76nwtJnmHAtGe9QyRmOX6WoNvcXYBcErS9VNy8Z
UtY7dhJHyNvCW7EOtn4cF7gtvqG06XJPSVo0VRZc0AFP4yyb7yCMvNj8liEHYeU1
VQmfeQhPgsEe7pQcIo4ILJfNNbNXOWS7naPVnBUms6CO6RBUMlww+0ReVOyUJhKA
Jy+Z+sEi2c01McrM2Bxs2SyvgvIHxBRPTUTc3A3kPuMvgMjTJz2Rd9gnnpG1HL5x
vxxdeJB3sblgWW6vWzR5gb2eUO05Gu5FUGc3VK68UI9y9ck+WhEcDfFTmVuQi2qD
sIeaDC44+kwo9RpDzgdAgxntUsoIogKafSzAw5AeTZiCa3pkBE4UzyH5ddikuezc
H/lkwVUiDs8YGYqTfb1LqpeZpeCJDLvRZ1wdOKkH42T6FnXC4CYCQLNmjX1M/5Gv
//vmV/OZPHEfpcXSbpnqGSiHQjf6ck7+X4ySNaRNY+Ffqhx3z5K2zNzBWOLw+ngN
SsjzE9fp0Ptw2gwDKfFXbnqhaV+dRK3fTF+jrTDpXcelzVv/M6tdYnKAmj3DKrxM
+t+1gcZjL500GQzy5D+2t9VeFbEEnXESxH2q5XvGEQIeS4apRz1btWot0/ZuMMSy
B6OMzKsjQIYg1siqI7RrFafDTgLtbTM5JsAPbmz1RRh4mBgqErPYhNH0sfFqBIYL
r6on++n4A/Mwn3D8MMVbGRLn0JYWTh/G+IVeBKq6D7NtMb6akFQi7/LN8h2DsJtC
MIBicsmaabqBtjytAtG0jiHJ9lHCUxzA7nbGh2AgOOsEtR3iPK20KOdewI61z16y
GDUhZcDERLxmxGDz+x0UqUJzvyY0CeamX5jY9qr79BZbB5RdAUboXNnaxy4h0uea
RNpR1SalBnTw8WqyhNNzbo14wJwHKo4j85gCaa5NHCF+2IoaIXDIcoGEkSdTtRgO
NTOwnAZvJ3t7oVnwM551TCaAXwJOEzuWlMYD7RRMAy7CD3JPdUg72rKGUo2gvTSH
wXYAeLoFLko8SFZgQR/IRtzUhv3jKD5blV77fQIhfDjTVslXxDYDyAWMR41oNJMv
+cLetGAHT6stnkQL7AnjVrZVgh9LpfMQUl0yUx++u8UXytg3Yv6wZGJmoQMALn6m
osWWI8NRCVtueaAxTdAWPtp4qpB1t4Fhf1F7fXBYRPk2rapUGGsUPmbW5QeWRSAY
aNWsOhgj5uYWTTgwYGKREo7frg6ISzSaFvV8ez40j2Y2wsveH+1zBlnDuemtJ5oW
NV5cgdqlKpFhePE8vo8xENlB2mo5Oue54BTXbUW6ODYrBXbd6q+4TK/YM9m3Ir9G
pb3YFSzeUkisTTbC9NJePnizVOzKZ5voPG8DXPSJCxkFt6jLlDtbANlPRzxsozar
SFL7Zn4bA6JQiStnhfhJjf5SkQ4khJKPnSFbl9auw3ImNaepir4vPyuUTIEdYh15
mn6lMrEfc4XrXu+zq6CbbbWtWcGoktpGgCmsH+dedxWbOEn9N0p27r8TdDlIMrM8
Lj+4tp7UqCVa1cbwhzd8t9oLUov3um+eRYvCXsdBikLV+WOwJEzd6mathNoR4al6
Bd95p1ZC74CFaBCsRmYNohBAQJ6KKvxoVyXy6w0UISAYoXndJxQOLPET3JIsxdrL
8z9ngvVswkmYigbhmk4GvtFaKWcz6uUyK8ZU9osieLvIsHggj6BHXCOixDoAxEdW
bKHkYCpys6gjRGRb8i5RnMPY6+i0GC9fnQWpQmyL0tW8Sc8d7w61Sg5IZhR98Apb
IOun0lp3HGsOw0fQH4Ao8nsjYslEeP/at2t7IC/6L+R1o9OlD82ZIXC97g4V8a7P
4LcO9xOpC8haynTIXda++0JHd/FNtd2VjzyvDe0DaINUw8OCLtHaF+ZtghKCXTdc
scyK//OcMdSVOLUObiT8HQV5mcjENZA6q3iqKvhtdd3sAoqutuqhMuEPruqSjXOD
bSFcYw5Lzg/J8eokzLJqMy9IhtbewP9pqYciutXfTBwR7bollTRys89rY14A/u5d
/r29B3YglFIUQcbAI2VpfIdso7Z/VQpfkhNR8xm3XnAezx/pQp7rbSrd8GOSt6D0
EupW9aFMpMy+n3GutWDQhutd1QqAY+yMccdXUv29QY6N58pAe3VRpjDLOEEIOElG
axQWPekccuGwcGtiMtzLm/XR+s/OKeJ2+jVOtQ8ToreyF0JYPo1FxoEYLBqE2C9s
WbOT5I6CEJ/indMd1sIcjrhf4skC5CiKa9zcVp97GdSkO7WC9Tiq4/7JNjygOI5R
vn+KiG373dUXCK2c1QzJb3F4x24+9vWVKHu9EqPP+NRjPaGplI1apvuFA1S3i4yV
vnf5TNgpI0e4MTOQQG5SIl1PvhSwXp83aEFfZY/xF4azNpo2qPLmfBiPF9cVXXQH
Gs2R5MtHY6TgiqudmwPJiEaDwsiGFjDe3JMU1OfpqzgVBVGS6SXHYhhhqklpIyhO
S+qUUbGgDfTTglsVTAdxUBJqph0sLzNsdNcfXIunrpUi4PxIdHo3FC8CqmQLUSWS
cERaiwm9Id1qGRFTHpE54pdVua6G8tX5Vjwp4+Ty51xlFNO9opFo8q4E4JZjV4Ln
4SkrR2JwuNAUi2Y1bIrP2nyqXtbM8j1tC+0NdrgOFMCUVBX63N7yjxJqQZQuGFI7
UYk5YlSHTPfdXM307lkToXFsz1kFZuhhfwYsSIIKlcFbvQNQfZnAD8KhMZMpjnU0
0A3MgTcVy1ad8x2ZHmjdk89DjCs9qfHZUQNMTATy7EfvRkVI8i7347T2yhJ5pnPL
V2krDDBv8MmHRWda39ZYNDT4UvMOvDGLf3Gnc1AGx8BHCPDJkhy3iTCeDYYaf/oN
HQ6iiAUqLhZjA7Pa1Bcix7v2ff2bTX29VxWFv2pHPswnREgKvsvjV0c9efa7uG8y
mTNmS9LhxkyFjyZ6/jtw7hOQspxH7/28CWnsJakslUTL8r6PxjaqC4h4i8LuCVU3
7jEDjjBFIzUeDseOIIISeJhyEqH+Kn6lQWDk7Lo3Q/AiLTZUKUsHD5UVub/yKE5N
Z5oZS+PiiJ3l4+j3VJ6gwOxKZwxHRlTG4aYJ3rRHfhPQFsfxMwZh3dR3bJwHs24/
STuyLYQwgf6XaB3S2+2mvrLt2VRs/b43Lm9bfVFmOJ/KKSzaxbVdBp/MAAzkCAeF
O7OUZFMuzq/VEkQLUbR2UeXG+lPmVfO6ZCtVW57IO+XIuPTYPES8vHxRDu2K8K5O
C4bErnYzeAEzeAW6JNdmNuOJRLrcc2BHttjxcP6tWAQV3hxX4xf0CRH/htSLZOTw
DoCXhmuxr9FIdRGp5Sdyw3Bkua1pEpeCD/FL81XPRjP5HV4l4LxzG2X1tevZwDXF
ovWzyq+36lojPkDp3i2xIyGQ8ExgYd5q7wj5pzde71pDlcSlERvw2fOoVwdMyUMq
uLpyIvKY9+IAWx1rycz0z++eOrEKT9OVVsww7iHwZzTzH8/2g6Kckd9F92KyL7Y2
U/3cCTlKTYn403Sot4CzDgOpqobvRr43oeAoR/G9cy046nzZKBqnvQcPMgrkXLt1
y3zuaowIw7Lbpq7RU8quHL/tDC8RRSaaxCyJtOpl2FF9c1xOOkcpYFWIXav7nrlJ
4lEcu6DrF7ar86zzrmkqT/lSQtMb6KYCZmcd+t7zPaJyTCnYE0spRhHsagcPOKt4
/ZBr86oOLg0F7XDq0CSCmUs4DY4eXIDwNEp894CKpnW1jbpbQwp7O4z5qPQ4c/Xz
kZyqetdd/MEBn2rVinR2s8uv0vLq/LH8kYwQDAaisRzpooQDoAA600m4Xj7FEen8
1kMRKEwpvT4eVSHgtQEjYPXvcNTp90cpxAehx3Mcc+9fKO/1Eri4rgGNVPHWR4PL
Ham86vvoNGHW0ZcenayYdCIblq266WqBMF4prweJZE3EqPNreVWNFodLd3SHclYx
+m2jT5M1e17rCua0G185VSPobjGucwmSBfrflPIVIlooXwq/6nUc3q44A2ChEsyR
L1RyNV14WqWxWHkwO0MB+prREkBnih0Yd7l2NdX3RuwDhzUKbrlA9t0hhAAVRwNm
Q9LaKH4FGY2hqXSiDFf6kW2qhLU/NDwHPxLGHF6fm1Ebg2RmS+r8ZBtIdmeB7YfU
QR6lTfs0sh5hmMd/gMNkzmzUcfEFuj5vxmcOXrOpVu1yA3z+VC69kdjK9wELjsCp
tyYGYUdgbPRIRp0nZZRNb7v22N9XSEBAAHmxBAZiIuQZ4Nhkto2d61hEtA/cOBb6
JNjlDRg/v3cLWrsniFkWqvgezklXNrBJBksHyy24n5SjdXA8oMA+m7pkX5SzW39w
DbRHo3WSZHKqcBmrPo9SaWsZVvvoKB2Lp8+zpklE/9FgZEq8VtALdRZSj6/LmEJm
Mowk2ZimtcskSWNbpOhwmIse5LMnbC4xo8KXOWLqoa5l/Vl1XMCgyVKDAzKF5Gns
JSlhZqWCFeZCu7OxGjITvmebDrJ3Ejq9ckV7lYmDHzGMB3sTLXESqhH/koh2GPnT
QG/6w3SCq/DIKmCopmGLhq6jIlgxYIoCSLzmAihfj3aer0+vsJ1dWIBVaSMdQ2k+
i0gb9Lj77upOkZKf7KhPj58y0oYVW3D/yrL0xnVGdZAFhupfhVWMSNdVS2edaDii
t0gTDorADo/5Y9RuFqLpw0yVp4BP0y4FNHqh6XU/oeDn7rzvMOXMWLNakYbTRGw6
pjqxeuhdwma4n97Phe9EXrTrQpdFBER1iNWVHw0iyUKJuxX/laarNgLmbJ8gNchR
OXnePYmwsPkbXzNyKtligZsbGIMZ9wC0v36mcbxqrLY4kJrb7244t4WEMvyNykHT
wOQdwYChayH5EpmpQyS278CbuWorINw6sn2m4I3d4GyLsjf7v4WNgtnoBQNh2x4R
jHv8KGHLhuEawbDS7kY7LYJlxchOrCZGGF43elmh6SCLe32bRiy7EWvHs65wqsLY
0oNR8+0AMB3egfwyN3FZc6YBHYxlURh7G3Dh3OBfl81s8B38uK60+cHDvHuCdLdS
jZU//YngEnTa3bPhw3RAQ047FlQGeppHGEP4by/mBODgadjqCiXU78Qmu9+aNu7G
FBRYeCcMAZST+KOXIcVEvtwMlKC9HVQHmM+6UUT7NAtmgLFiUk+keL33FbzRy8sY
DtUS7HKwwlMqymF9f0vvC6RQA3MBU3X/xrRA/hKjdd+c+s+cqvYGhnLAyESY3aGD
yRwnmSRDBdPdxAECLcrT1ORnt7c8QT0qklp7zNzp2dMj1cS4UV+WlC4T0KFUthwV
+CM8zvr7WE+z7qDbVdOUCftOE2gukqzbLde4/XNJ0vI7yYbPUNcrwGhxlJ7vHUZ5
I8Udd5q743h5hhE3z7X9+sEMB39vNHIrAmYsLhLc8SttMwcw8KRaNIvHBx/oD+Rb
VvFO8FYlC7DxRoxXlhKZ6Ka+JhIzp3m5d0rjT6aAzPdOr8FibPulzKrF2DhZDzlN
AQoRnOuprIYdjtTQA6b5upGkGl6006VbpNSU2kiQezF8HIcBG1/z6PpfmKU2u8na
3zl10ui1fRv3VuWpHYWJj4P2tJWRf8k4D7aHU1CS1Vznzlaick5v4W2wIMLdzr4+
KVT4JVppSPhk1A84BQ3Pm6FlnjOP6t+2J3ficMIrsobLb2raCGVHPqvU1K0xk7mI
7J0LkLdPowgzEJASW1+RIgLL3SZBd+9kl+4jzK1LV0k4OijbdCfFRZ6zdFDZSCCd
hWDOYcVTn4csegRxK7t1u4THjC8gAlPqQOe2jIPZki/hBa4f2rDvgI60iLHL6CbE
b/XghJ7WL12vNPn4E33lHOIsk9o9Sy+nOEbT5ww2EbQpUGFFGK8MMinSf5t/ece/
ihKXqbs5ZI6NCiu0yFi7rz/Sm/RckAlDEBabrlEI9+v84nSv1o9oVh+crXqFED1a
HaTiD8eL39zIP2CDl9JJsbGyEDaMTJ+VToRfdcMu69F0xJtMI8JbMHnQyEbtIrD1
zss3QrpWv4zOMIpTpxmF4dHnlLWcTWQgYBmBXNwUPvUsrL9tfOzeGTLOnPNh2+pE
NbwsJ6GdZHF213TzECL1JCa3aTg25ThqvqirM9hi1V9+gZU2yuDftY+GKN1J9veB
degCVqQl8bYxgUMCYW4ume9o+UtcfT+NbAdPncmBOeSn/nAwhEGR7+dxyYJrledh
RDYZRvp2sX0GbYYvmnYFqYxCyNYWFpsGHvsBDm5MdR6KnEq1By+7J4b5xp4ybajP
1w+CGAbuuNTlpn2XhQbj3FR0LPK4c0R17Enm/oKjHkaD+RyX2xqoZy24gyRQDYOm
yrmlTIlvOQK70aU7JWjxmAF9v0J2Tjflcn/jS0qqbHon7ug0HXcxZ7By7Jl1jcrr
lIXrr4KCacgNZSaP6dpesvy8X1fYacavOMSMk7E/Ki7Sf3C/ygn65SKVVNVFQ/lu
Rz4xNeAr+gAA26hSLMrICOAEdbXs5TSHf4iC63b9008jT5T9si6JCsW4FAbsHsL6
u8CsmHtB1ewl6EgoHrrjr3sQDzg76GmOFIGAQY/666b7xaoQqZhKQQlMhhTNdVCr
AVYuXy0A8nCeFj0rzSdRkOBhCtWwVxHeFxpBkDdYMYg+D4KNLbEMI1jaDSpT3E1d
cXBWlg/QszXgyysDe9EmPUXxuGswsm1NS3oTLJhKLk1CmP6WaV5V+ZkED+TY6tMD
f4Ocd88yaaCY+o16jIwELT0Kp3SBeDlJlWNiMAWDWR/tTur9wRWtnr0qn1KEDeUE
DNIxrJGc1aL5BlBXTwZ8Dbghl1EAMK2LcS1wB8z9Iog7pKutxsl5iOVeYtEkBue9
JjPqIQ4ICUYKUzMeAYPKWhotPXNuSFhHhs+bAIP9V+GOvMy+eNOk7uZ4lQhCTTwm
NKlnnVsZ2AYaNYTGlJAaW1my8cBjRqDL8Bv+oyRe9ynlvnw5W9Kev4nXFZPO2PZX
CdY9zI0sW+7ZB1mfKaQcVsp9MvqtSxZc9Ax7DOpJnKZDH4sdv6RRrGN767eDtDwF
OdgzjVg17Rei9Fc4p6ajzvhbzb6pV7DRrS69xYpqcMW2GZpf9i6nKmi/ci6hMcPB
z8YpLu80eYe4/ShDOIbKBFX8AWcJpecNBWonSZJhwCj1YsPtZ8Z0rmUKrNqZ642o
uEOfBpI5LWHdbXselN0RpSXKLGFAI2aTeeOCG+qoCxf72k7hHcGYGYmrE6irTb3N
YOOG0De/+n4c1NBeFpl5cwWfehRUk8ILVYjnc8+f7DiUzsFgvmvGJSy3ZHCr3Nki
ioHf1GUeJmBeCeQWJfCKQLKziB5VDleu196LNFDaB0yfhR/PwcjvP2ntkuQpeD+u
H1oSpHVRsJQNDx2eXr3FCd/KEnCLsdM8FOaZSff4uzQBY8qZxpaTuF7Zw7tLtsfH
tcx77/3LRbRz93Sy1ArWk49A+Oc7kjWKRGOgSEUgmUCq72ScKhWpuaqGKLCH7jNq
P6ZGY28mdunDN5Tv5q/U6p1YDm/7Hy2xGSzt7UNwkALomgZWT70tZt4hHeLp++ir
QLbndYXsdRP6upPGqRD72Xk7WWqkSVZdkqg6krhxCnOUIic6BXPijPF/uAxNVpfk
QsStDJMu13aYd+Nya0UIo9ug+6+g7Xq+mCQxp3mNBLq0eJII7VG1MM2Y6i47P2OR
7BzpfQzZWl1fnxs+cHXYm7bo4RGlokdJIFX7KA8XEFP67ERzJ83S5kEvUPfKkEvG
wRPUH7V8TUY6alqKavbRMpCVnYG2+JXxGy+LXQQTBB9f8Q8p5oOi2nAux0PiphdR
+Iz8AIceQjiJMAgdIZXtMAWy1cl4xqVl3JH4v/hgwHSEe1mRlw0Py++vA78p9ByZ
4Wzz5CafjCQEwImiAQm81rPIcMMq9Xb4Vdh2IF5Fz4VX7J7Hyvb/EvbE8VS4JdBo
STFvF/Z1jwquhCy5yAAa9SRQ/bRXfaUCmIk7a7WjB3jXbbCtZgXR1HOdR6eChq67
m99zCXuFl303HeevhozeKvvw5PTVAbKJ21pFU1nF+dz4gnBLc3kL02QvmFUIYrGR
Z7z+ix4qi6uf0XdkaltRfk+jl3L7ShIeFAUy0gX0rAEP5HaSu/6tBBA+dFFq8pK+
E+QosvhItfcvGkb0TIR8Dic6+hb5SrpIPkrFI/OzyvJEDy2nB0KZTrOmjXBKxDII
6DRRxqF7BzJxVoq2V/VHyiG4CgzeWFjlkbgssu1gz7GC4BfDQgCOO4/Zaqpap8w5
vj8hnJdCPKo7qImW33/iY0hW2+FSdXd+76r8qFwozSGvCxtF+d5aeNIPVlKxsPpv
iVD0/gwA6877dcMiQ7jUZsShvq1JZNHH/nEK814bTOhtuX4wcbMgxynCXsWoIoGY
GzjwLJvsjDp/cnK4cJVqHkRQ0b2St7XKrw3yYG7SWlrgYjdgHWm/985Ht4Ouy9oS
hlpASqGdfC+cNedtfEipmWlpwg3guZmNCgGY5S9ZGF01kx2iITGtnxNWiZD0hXTI
Pgz7ffTUZIvLGTNVrabRUEVe+tL/I/SRU23ib6GxY9g0dBU2nbz+dRH3GKUTVF9t
lWtM+kQicnCZ68MzL6XfEsxZHmJcaFNFlx4V6Yu8IdQV7sVeI5X/k/ZLbdsswwHp
KY/hkHgm56GyhJJr65UOR18dBBlSDpdKG9GVNQWWxUlbPZ9/YdnvBICExlBf92L7
1lHbPbo+TPeuJO/tkIdYmKNSvzD/A/wpcyJ2BLAaQ4lidUi3KnnR2LVvDiPwWw2x
05jKgZaHoH7AeKAz/OwpUqKA4DQ1IsqtxVh+tqr0m+lquZRFHKbCdsHTZM/0Tpy8
CbOn5hLRdsQWx7tWlMlVnOA5pH2RVAiB8LHPwc3y/Wyv/OTrcD5sJTGxhXWgyx/m
DuO4dNKsYmamir2fbn9e7YZlJxVG72q9ru/B9FZ3Gl0bH0gbZNyqFvQAzuU+yPTp
MwO5vGz4naQ3TmvzKGseLkJ1fH/Q/EMU4lc0sht1bMBsfZkRO73XJhLYZ64tPnU6
flweR+ccmleSMGIYyNQ8lmW8SzflmAB80r0fArR6V44a3dH0EiascNozSsUx5ceA
j5wgu5N+GcONXCgqzTJZGBSvxbFCLj98nV1hUhsIRZes9Jvg1dktpTEOhDOP1MsL
UOiopM2FuJv0awQ0uoc17yT6OdjH9nf6X4bWdS4030pSc8EdIfbnshjAtcwjfYyi
1qtxNPnqzod2Wg2+pLo60LpKGjcuB+DCfgtl2RLXF+S0Rb8t75OcSXmUt5Oi4drG
r5bhRgxSSKhV3L46/2RHdlbaOZZmadFI/NjEA/1vkMzBLCE3gx03n++sFmYXiQiN
L/D43caQ5XkYoWKkH/Cei2iJW32FDijqCYZgENr5AvvKJgJKnnAxYN/+T0hjIgWs
IP6GEBkHMF+rL+L482HO9tnQyLkBREJvNT+X0EkrVd5ZkHcTGWWlEBD3lHdVAU6v
S5jXrVyysyp/F7sVmYk6CiNwgDlGwj69BVTC24v8HjiZIDwFpJXd7GGqPN2Gkw9D
o5GRsffN9pWaBM7o5GIUsHxFlfQ+CV2XE9ZBjZTuW4gNRSCmdGtKVkngM4oiEx+V
xsEyxPb5g6bmRj4ObmgdD+1e9eADgpkouGWGbxAW6gMqim2B9r4WXT6zUApGT93Q
ObU7RgLDB+ppt7Vv9KIGB/pOW7VfxEffY009BQ1Ia/X0dpayG6gYpKtMoostl6Jv
a6ApkSrpcY9W6YOM8ILvIFUP8asWiWy8roniMnc8mojbomH98TGej4SrE2GrlTni
IcZ3zZta5vkny55V/8+8jSaE4sjPMs4R4WkBzduMAa6hPZdfVHyLqASfXPumxsNu
hr4XO5EsVYWBcZ/jfCww5GkEMTtUKTSxizOPS1drwwjxIzs4khpHEg9j3NaYrZZd
3Y3fiPX5QrnbfXDmiouNjKM9n01pTQuExLMda34FfuIiXmEBfX8vPrXPwb4l1CKw
Q7db2qHetPJlLTyuHqX2njoawCP3sGfT9DTqX7DPLbi5C8kUG5n22vI84SBF3lHi
bVa+ljcUU0B3ddlPdbWBCky89te9M9dz5wSILV0FVwqtEgh6Cdwenxpx+tf9g4gn
9ysjpQbSdPFdTreYiOou5gvg4eeX5hKUPnk8oEmTZ2X7hJKTuyGN64FQdvFX8RAM
9iUgbjma2vlbumxU+DliYH+eTPahf2rVA6lqMPgYHs2nxCzrjJ4qWwBRqoQVsPPe
aHVBYTGpLcA5JIL0fl7jm5VozYs8WqGLA3P3ZHMKEPsoVrIXDwoaKCGwlYV6OZXj
88OcaOpALmeHsCtXrayKXhjx44/QB2WJDkAhzKu4EuATXAGqewC2Uw8ht0gxAtcL
hrxmvKOm6BeuAgH5YFNNinzhYOfgKGaEM4WB+MtidG/sJEnl5NVc2JcZ02Cno4pa
+QA3CvpEb4lcZsXP4MbrZauPy+01IJ6/K9NUK8AST6TmXAR74LYXVRNV5jDWfnFj
1uyX1xvbV6K69B9xstkn8AP3YW405KAWufhJTvETuNpzIHOlOco3NhoWC9lkT8aw
LeTVAoiKdaQyTs3mpKnlDW+xbyx0vhWB+EvWr7Axl7oam0EDDOMGy5OqHAFv0skJ
JnSoy0RV57tvqPk9ehGy2MPn74enw09hijnG5H5wFFiRaOU1R7fk1DEj/TqF7O22
iHfHalR0t6vd4Y4IAJ3PXKm10dMo+HiQEEM7V0P761sfIqssBPIG2v7c0brigXd+
3D/27nOTcypbe+oWq8GRjXP3D7BVQhSQB1d/nnNyq0rauwzGnapnxdbyF313z2WY
Lq3HKWVFIRQGZhuUu+bq35yy3tUbbmqj6QVYNSn9U7QdeDHQ5BS3cd/UZP/WUi4d
UvwKsMf39SH3cAj5khKc0shL2Pe9Ykv5LiMCd9OQyQtEjHH7Cpavl7s6HEGdeXoU
lH/79hWP1AT1tn9ej/lw5+QFDjqpEhEeHlUpjCdXfw+cXAXSqVwm93i2LBaEM5zK
8btg9PLtrym/8ggZfzgUGc03pkcuFI1+/S/5mNmE15B1Ze077VOHQHHWCGTKQyxj
S0fTgKTbUM+F5Ik6qvst/hgoEWFX6GtSpPWyliuUhpcDNSoJTcZWO+dbnOI/Fioj
CDnw65Brz4TXI/mC85XP7kYB03tGC62BDXLmLabVNrXzeVYT6k9erfB+ZquC8671
GthBqcUDoJU87WpZsq7P3Y7ZqgQmRnQozCGvaz0rt1lBqA01Ey8ytXorRg0OOxte
CF7NxwG1U0OkltVe77V+7nMa6Pjur81q8EmOE0IL5SSa9So0jxgICNCngZ7Qnnhd
o+PdhRbpNJuSmhw8DmKd/nd5I7RNuZVivc8rb/1FvZKcE+ANh7yPJ+tt4L+fHDMT
2tzXPQa0Nxe893wLcMSm0k9wqUFRIQq33KBvv4BBoJYxYvPzgls5YYZ5IDxQ5U2k
Td5IajXHAYLM7dFGH7ol7BJDA8lpB+ihKi27bxsKvNnA1aI9c4xWtlhhX7RG29CX
5kUtPcXLiTdXebQ4HIbWm32mKCWJPZFezXSvxswcBr+PHVQi9NWKbFYvXlkhLP8H
R28a71iLKVh95RWkYII92KzIbHqOSaH4WQ3Eav5lz4HYHrPrZ510bN8gBsgMcYdN
SCNR+edFAHsqJVOqCT7+zBTjKZiFTlxxLZ4nU3QITPri9L8L3mZD8JyYeERW6yZO
u70/zx4IqvtLbgtFy5gs8K6a9uPTueq2h2riUnNLK5FfnFHtZw55Vk6ASEw+kcZC
FSDniM3PgeFc+aomYh3KWUtahi11Xp/yOGINVIluaYv3/RRScPG4hD4v0qOr3k+j
wPQxH14rn3Q4ol8V36W5ljHAW9N90ixzonnsYHaeEzMJ5QhBEIJV7GvpsjD9MGEg
OKsFGwYFP5npQ4F2wp3bd2rhLSriLNBRtdSaZ/ULl6g5I/iSmQXwrf8M1K9mBbQH
teHcmjx1r3Sv6dNarubeSWZY5/b8clJO8p2/iYH+mJJ/lZwK8bIdEZqdh2P1OMD6
cK/YS1v5SCGh1HafvFj91Zzc30WGryRXdoMhusPt/wxprRpmnG72JXSPmuL6RawI
nVoyVHUrbsxGxmOORunTWGKhhzJh74zHk4qkBqfu5RW8qvjvOOfgzhqVE62wVkSA
gpxSmXvR6Wf4b6KmWa1Txy/V6S9jfX+q4W7t0ECOw0A8BhvCkj0OnZrd2+3eQoYQ
xsCJtDtAR/k+K4yrK+aOLGUDBUBywEjraBfawwGRloq1/lPoab4L5p0Pntuawr0w
YGuhyV4GND1BCq8dFNEJTlIOXB/bVHKOABRgHCDFQVKchgqKV12JVC1lwbdZ3p9j
vbrA++wRoGV+oJhYGh2shXJ9Ekm5m1nYMSI3dNp0NeiUD+cLDKiiBpv9jdxQIeGs
0uIUR1J49pLmFoMmsIqhfhlEVhTobPaLuJBzfRVQnfiJ8rdNzWX8nBHwcJ/Q2qIr
kHscuohNPiKfKNMw8oN7PDYuR0NBLRXsWakADaQVluBi1Len751ouuMr0SEEwJ50
RZx26jURkR+5bICPoTe60S+F0EzQ1+XsFF9yR+5btVSs/DkgLdXVpwXQ+UJSPsaP
IkIRpYFzjFOOe7YSGs56D6x5e1E8R9mkhjaJSIQcYQuEW/37dSOAS2VH/uTVoffQ
s1XCaLJT+K7PA3i1TDetWprbC/+zwjktaUA16yk+Kc1R6AVTu+JrFeUUiQUr4ZLE
SBRBJRn3s2vdOu1MMyj2rN6NL7JR8JrSv0XeirhHF2h3b5+Ub7xvk1OPQdBpUNJh
YiCrE9xmuhieejc3mYL+E62DvSEd9kYeFLHEak34F8CFlnvvHw3K5w7ArOhqlNFV
hRwANpFuXrgTFV9ljf9dwOcVjocHaW47BvQ68cfjOSSiBpxnSuXb65qmOj4oEBP+
ceQQ06QX+VTvgK9lgwNTi8jJmQJrYDZavJCDiHBr1zVwt2/ND9aURmhfGoM+ofv+
PfJNABRyghzliWjbEvldg38DhzSqzJ4xtMIRTMy/9z/I2Z8a68/F/Jyohl8bL9Nv
2DLRIbB8xbKPoSbYhYCibjotxa5+D6JqISm+Q6FCOaelEHFZSebWEI6iQ83WPY6C
NkagtDS9p1TbVuuF9/1awyOJzHomQ5hNzVnyL9oPWLwVe2WiQGgwWByecz7J025k
mymOWWgt2qqiEnxc0EOrVmj9lX8YixlzzLi7xTYRTzIsgdAAlWbiBugWrQPB+0fn
fSoLlhRVFaQoIY74nCJg/iVv7hbkYmCT/moa9Spc4lyXBXf5WmiRZg7HgodLfV8a
s7iPs4mXLHPNpWi838L3/Mwte/uG2682KT+DqbfyRyKC5kYrgw/z+AgbdOa2JZ+2
mAXWNBxs4/gsqk0m0vwB4Fa9u5INs/8iR0Hr/T4cmfcxy4pan0Jz1Iq4iNjZWY7c
crhSOuTPh7ckj2dtjt4amlBEi1zfPo8sM3BkGHsyCxSv1V5+MsWCkBDbaHV7YhAO
kmRbayvNVDwXXwLfAchGAh+GHY7cBb0vJhvmiaO3dAW1vveRlq2G8DXEFniJh+0x
wL4OdHy3rXvb2dGYUe755Wbs57NviVKO2Hcg2ZGQ+jTz1jDOBh5CBq3nH5X0LY9r
HGV1pBLR/Yev9xv0t/bo0QZ/0J6ij2lNzksVxkAJszCTSSzG5ZdBuAkayOfD3O87
TaUyhRDcsUAe3obffkCkryWpon2g5RWxjgqvxjdXCpnGz6A/tivY4U9h0NIsKgBt
MnESdo55VGstpQDdAyv+hoRqIgZsFxjx82wDJFj4VF5aL0/ZrSUxx7OmP0YRbWSL
hluTcz7B+OkLXFojoetL752UABxuuwIyTi8Dk+0tN6HCoIfKETlrE8nFjQXsBLrB
3bd5wlOwGRxbpccy/j0mMDK5vfdXyHMitZ2Hulwn4Mff62ZTBPLXe/+faT8vp1Ny
bQVRD3kkFlXGiuQh+Mq8eCIIZEut4e9cUsOExci4bwAZRNpbuZbMPPy2f/51OTZ9
5BChJtC+btB7euLqCgCjnOI+FxKcAeUcf9BycD1tWf2Z8ojnnpINoWqcb6ue9r8d
Qkt/INXTZOWU6X22UaxNYyDqkyhDCpKiAOnj27n2oWYA/YxMuw7akkv7TaQcYT1p
GyRGGlfua7ZObY688SuGbtub+8uu9RJFdUTWnca5HeWM5LUbf7IvctJHr2cOi6ST
LdXsNcHH4/73dEZxAOZHCJhX8ANJw1VDwLQCL6ZttXoHVxkHYUUNrIpfRLFcfBQe
ZE+ah/UEmgWnBu0g6zfXJ6tNh0nDGFo+Mf9UYd7fhZ+BhgDNP+NwH22lmDF/Omwj
8gULeM+XakOtdsAPfpGr7SBrKnIwbQwfJC8jLBcgspcW6ac8POAY6DPVyOkoX/KC
9K4WPSdtuCq0que9z28e+7dUyuxC1UEQQgVGeH8acqwHyX6ohOKgeNr+/aB4+WKc
V084DRtgLZZSUOaYoIGjeddvsaOq4W5PVPs2K4VTX3ElECR/jJqyPISBD4wCn2x1
2q5WHgoqSpK6PlpoZDWWwRQqwcd+Y9PaarpRBNHHoPP6Vhkc2CZwoJEIlAq+k7yv
sZazL/M76VP99+5WEw//EUFw1376sof6571TSrZq9uFqBcGUCwAJ3uIrrk29wCPB
wG4f18P1hk+eYAqEjMeSPg7Xe+ppL/mWhiMOKHIul7iO/S2p99MCJL5NsyXkeOix
+V3styqvtYcektQ8naGSjTJDNve6iZ3f3T4K6ytx1vO5MGFp1gS6nLMci1xHW1KB
xJdFeuTKM9EwOfAN7u4JX37gTEOKBIMFB+VnBWFKWdTnzrLv7TmqHboCGQ3FCkK0
zjujmB7zKSkWQW6tRzx2iuW26UJYeBf9Vb9Rjz1fXyTCbgy0tJvkzsG566ciH4lW
qgHGoCXAofElxx1vmZrfEjSsVCe7h+0ZSPbOnyfDzpix3dV+KeRSCpSlZg8AG612
p7i1cPpOeXrPRlVlqEZV6o2WhtB8Zyd8cmKPBVM8ZHs39Qsbwf/wJBzgMXdWlQ5a
odXzMiUwc7lUFMzePWkYSFTnqp3ugwYoECRqgtJrBHQOVLwbgxgGpnZNKsWBVoG6
z0NnqEuSof/dBi30QHkbYQOfTxZp+N46tblK9bHGeyoHsqDhwpZLG1S+B5LMRwhC
aiNJOFMQfZdckCm5yGlBYk3tK04twH2voZ4Ax43NqcI3OrjdifiOo2aEnSk85FiV
gY5UV7BWmniV8qvhGaRivBmPWB3Z8DaQiue6xHpXLbVK1gzAl3OcL6zDt/N7Xgk2
cIbJ6UzBrsEChD2zpA10ETR9qC1IALpxEeiCFlXFjq1Fs8Z3Sj1wcpy2OahvDAT7
KriWQtzsUyETC8FJUi/+5oIE2NoBDGWCGRKH4mPLhoFQuqkXh4g2+uaSvf9vSpwi
ENlwM5bwDbIv0ns3CeSZsaIFHHt1Gl3P9JuJrfHpWJrPi/1jjV34bipUlrHV89E/
Rc9JrF1u3HTQTCId8pipxELGJzPjM4tu1ojMyQoTeqfHNQbv9J/TScs5yvRqHXf5
1w+IEu7t0vds2eK3sqwVuNHoFkJSzxATrf84C+J1aWCs0mqDLVu9qgDzo1WBi2Y0
GGe9D2SFY7EE/6FE36RTMwY9HYTFWYLyi64wdBTiJb8PZa2/OA8CAQ2cU5oLPx0G
Ll0B8OPDn+fUj02C+sNYmp2pe7r/sFa9nSZpLqqSYWCxg8vAmd7oeD68bl16IuDY
0i5ngr+LWsbkhip4zeVDONuagiYjfAr/umtGl+yDInKmbBsQJkhYiJcdwQ5TjlvH
QwSo08ZcQUSZIwbQbxys4hdl7KuTxL76dsWUyrRL06kiHpjcwlSSzhXEJGLlZyl7
mbJeMIpBn4kREuQEwy5FTA8SeSxt7O7F5gu+Jpmlph4F0hUCIqL90cRX5t92iHHv
thevttI46fzRNyxp/xRDL8/QDZ456f2dzcfhaaCNbj6B32WV5IXbsI4+NZBej5GM
dUqwLeKoiWNMOdJAHp5PnaniJxsdRGDZglmGzuz3ltnRA/y5u0NsraRzI7habJ/A
KlThHg251lFkDTzHhd92+dq5rcRnnvoc3BRw5+dl2F/xLugTXAN7OwPZEx2U+WLR
iSyDD3+O6xTEY3EaDT/LdEYwPlsx2tgb9hxYYTBQ9bjeG8MgtLkHWk8EIZNncGV5
lkAuFcA/z+F7kB04bN5vcOG0iuK7SDf963KITSm6B6+1CLm8/Xy+Y9YhHU0hO68m
NL3fEiXRw4yq07lld+VQcxQksUBNznC5uYvVIlqaBcqzhS6ZgeyLH2nfJz5rQHBK
RD2Q4ALeAH4gf9RFC3JJvfIFzcuPp4M9eVG8Rx9YUBCVqlLChxpMFSJyRZ1uGmXn
t9+5wPc4ql3R2Ulc6SqHF0+xZ1kpKLvUl3D57ZIjjl6i3TANNCnmwX6wAkGjptf7
VZ3p6gSYoj7lcJNSSGxIndu4YPvjuXscxn5UCX5OejNghFN+h8O4hOWQDZLHM6a3
8Ohxn9gCGtkksxX+h+OpeSlJo58br5RVSrlmvwsz6sGMcyNV0IHsdTpUOuqTO3qQ
NdQzAvDADgHHa6aoxo/50JDxUHYqpCiznk7nFxbU9/EcDu6Q4DCMsM2I5ow4AxEY
k3zhCivUSMo5TMMHwtSb+qSjWbYiSz90CS9GYqcpuLTkoYI8fKmWfuZ1oFNw5IgY
fK+anp0Q3abrex1OVWlqRNCbMGIgASS2axuBeEv5e/tOsadQGXKROFTKd+tdDQCg
4pZxSmDSPJdkXxaDOcn2344TYikXYysN8ame8v2ovuFn8LaKG8F64/8ntLQGVHjF
1CDUuQL3koJPwVuOlEsexuPGFB0aAP7EjgI9bhRhSJuj7x11RZf2zW+JqkDxNwh3
3XKt3/T/zQ2fhvQqlpbXz99eI5sxzHuJpMXI5QK1EAF9VO/4RT7QV3XbFAbtjEod
Qp9ZmYFKMh+vq+hxHBTVIhv5mnSZu8rWrY6AZO7580Nrr7Hm9SYuoJjzIEZF6jvp
2cpZwD+RFmLDPeynulXjgWg5bz6CKMJoJs86wVu21NVNR8h7oa1NYfRB9E4y9dFq
b+/UcEYrYqPHgeGzcDESW44u1sVFvoL3bW3kSSkiW1gql3dt45Fq/vnK+RChvfs2
r886fc1rFq1PQFk1RR20J2sxRuBRXi5VEycdoU0s5rjDNZ4Q7K8Dphiypx/Hvkmu
sGkUhy7VEosO8KzWejGxIj82tAkfwqEu/dWZiURa78mosTWVK8uKINNO7p4Qfrdp
FQ6jfYwud/o0aJm/ED3yOTWt7UfAM+1z+gqpaBludtYqHssgk3r4plIvi/9eshX0
6rWofYABMxq+e4ITyjNarO14jkd4uJsZZ1+tdVO3Dixymx0JHvN3ZSsWqvXniRkp
OJqi+OcmzwfYmttMYPI+X3H/sbELCJvh78ZmuzMZ3h2hrPi0G/QRQF4ZS72I0KL0
HIwfk7toBve2oMTpfHnMaQFlSSQ6HxuZOxTqEG5sMdfONfbIp7X/Jl+hXVen4BPj
ZavPoHRuBOdwA+ChDMMiKiQdTgUN5gEpEW84WeFvb2O5ohT6mxVM66Njh1nvWQ69
tr1zWCzbcvyy5oompW/LUi/j0eYi09YhwnjIcdL+xg7oefmtSumXyyIJdXg3WUPJ
OQwXEQI7FEeFyFGQwlQmHEeNvqPO3gWjBEm6ofVQSPWrrhzzWy76UD5uE1Bktlhq
mB5/mQ44GFb9vDVY8x/IYKTR05FskR3I48BybEc4dezPqnKV2ukzYrlFhgafNcEt
jvCEWiG6AiAGBW56ue6JXwLCZZ2cEwhJagg5AeIQvQrbddG1h/Y6rIaQc7IWYjDY
rcH1pmqkyBxFwRWPjX7bOktgKXD9lvAHXV/mIJ5N9dqMkdhJBjU39GusYrCRi9Ru
vWQa34e/lUnUgPEyqdaO5yNY2RmKIpEjGNv1w03K+HT+ylT+hG4EUaKi6t7F4wx+
mU0onaw6dTXqQgFFSE5Xa1ahNNCuhQ6CO0esW9fTkW2sEo9vGBks+twovosZ8M2T
8vXCi3ck0+ExS4ioYAVnHFMyYj4OibJqTukcizST1CzcOlofZFOjHB85QNUkQYnP
+acfD944AiCH2tPUld3a8WVAfGhyvymFemt2qvEJ4NNlCDP8IOhImv0BxSp7pWlU
yF7FfhQ28F5wUcaIajs26keD642IuoXkY/w0pYQTJG7CGyG1ioFmCyvR78VGSw0T
zzLerZ9qdy1fBcfyBUhrG+8PYjUCIXyud9wPBncGy7kQyoPPf2Fs3YEoGq4G7klO
TnRy/Ek3ZM3hlM6ZmzZ1X8JAVS+7NoCfWL2/fpBcPobmaN29wAiquMNy2JMd9/0x
S8g80chpoqP0izrQ/HhLCvLb/WbCqOEFIQ8Wvuoyydp/NoNVloZ7k+7YzUhJzdB2
e/V4XPbo5H0LgpW1TrjJg5WKFh0q46yfqy4VCAZ4zZrk6lR8NMrnr0KlKpzyy7oz
NKNlrvzITdELEZjanqw36cZK5mf5nPh8M8sflld831b3bd3/JLlrQSkdJjXUKj/a
S7VSYm6Y+6NT1bSRMEBAioAXkQYrCg0x5WG0/QQ/+q5f6hsdXTlBULxdaPRp7zuf
nwFSL3AdzyPFvqneTTMEn42k6X1j0Ng75rJc5kWJ1gy1tK5Ui5/K3WDRf6o7wRtX
IA3Zp1XZxiz65GrcmiwlpCl3XZ7PJrmEXf7h8BXxwtw/8iJw1AIo3VVr6hAI81n6
QutM9sXwYRf6zwvZxqx1P3LpfBMxW/fHhb2KvpmWJnDfcZ9ApoGXqQaU65eqRCK1
tKKq0GXNzwzxxPUS8OghjWyqidpT5My+u9zzcjK+F+eLxqHSgzvg4cSzTdeN3gJw
KIm1dsRGGJB1mUMar4covpJJgY9RZQfttOM36RJ4PBr2CJhHS7g3wnq+liACdj9T
jjwZr62vzOSKyOblrpMa8WSyQtfgiCtMwapgXxn/tjWAN/wsa/nQoV0Ps9InoYFi
OwWPJJ+X5hjlT5TiFNcYIdhnLZHSMy/fZy7ZG/g1OCAHgp8JnloxaYDgt+b5quo4
96cZjnMVqBuS1sXRuyzUL2fXnqQMQHw8h5HwyjEoX1sM4XJl2qzBs0qNht+nUbaw
hg+Yslfs9JxVz1KrtmY5I7BoIu0X34osQ0YmywAKljlilHMc9m64J0jBAio6B+t7
wrlM4AkKF+OfzKWH/0g8/z0HNF8wsi8v4MAUwhnk1/AhtqK6f9PIKd9W741vNy7V
O7biZXjf+JKa6pgU5/LgVmUIJpZ0miZQf2GWqjlCsAGJ9CVuPd/FhBL7uGn2OUeF
YuqEvimVpv+/D4UJfEgvEPCNw91GG1ZaR29V+QWQHd1xmzwnag1PXbI+ROp7URlp
KJ6DvM6IO52+lWBbVFJ7Q0m3SG8vhZAEzMb4Y3gooTJBCkMrGy2I2LGLfgdPJxUU
oJU9UB+IHGddQ7lMWaVdhEtzHT6HSbBTzUA6lTPbfCFgkBrMH7SYouDPsbzZSN1b
jpLUnU3vVdgp8wC0RqE/l4AbbVJSN4K2FESpNoBoeyBmaEYVXoGufZ1qng7BD8MN
pnc6nZ+lqpr36W/yVsxHeTD1ZYdzkT71qx3zt07LLLxRmGjo+Scx3wD4RC2/QeQ3
Q9f3Nog2ukmAExrVfcYjICfqTMLVYICm6Wvs/+mwawAeI9K1D6EXyUZoKhuAmKPM
V4a2Km+rtSy4dO+MSwwgbBOF1WMchoaAxBm6mLRmU1pWPHgY/Pcdnp3xjKE3HP75
BOSmh5qZK5hfB36MrGWL2TFzNHqwZpEoZbe82pbUyu6YLe2e9ErsHiny8ng8BMYi
fZYCskCn4WprzCPxpn+mvfFwJl8NrlzgDrXGMl8wWe2bJfaFdUnPwYy/qid3CgWZ
vI0LMm8FJWc7ymjpWm1r5GuNqn6vWPydOp8cWvnQ1wrrKvqv8AA9+jwWOn+aw761
YHpJlA12ncbySfEgN9MqGi6cBp7oLgAUtv9hUlNv7SrT2SMgoL2AG6tSZvgWu33j
gxGrilaecD4DaGdR9/fZnm5sjYSFErlo7wnN/Kro7nqcjkN7JqVa4IdLAb+IAI5z
kwVYFRCP9HkRd9Mt1zk3O2w0TCZaJdnZSjAymi5Ka/7PC1SGg4H7G1PCUNek9wIR
1NUslDaT4sZGaRcAIK6W24Qc4e1gvo6unS3Fakg60rfXUcOIyXalPkuOOoLRN4zu
dLyOV8i+9yPWvMITZXQFCA34flogffqSXSB669iZMs9kCLmiykkmv1ypau+Wh/EA
e2M60S7ooWjP+XWa6i41wkK6GN31yOr3tK9XZ0kROJFMgdigLiy0DbtRyiNQoxuF
T1vL2mgtOkHaLQ6csFIbML3WYxExpc8GRDVfeRtYgYw3GCcq9S2rfv8+Kj5iBSST
CikWNiXh8FItLR8AlsLMtvs8l5DHrc4JXFe1RlRjXBeFkfevLJGxvj2tIztSYLNs
0qsGiOioq91PdYIlu76evc/onMKg0tbDSYgtNmeR4hyvFIbXH/9PWFEzPf2cFmAJ
WzKdpHuvePS7kDF3bq4hvsnDrP49eEEqtoUqII/7Gd3WDFE1z13YwkQ6A9sSGG1z
t/i7WALK65MXy8jYomKVWS3OcKmON8r9GqayHnpNrObouA1n4d5wavQ8nikeiUc9
AZFGog9C4gvlmb0dnBga7k/tsQ29NiZlKE9FPuPDbUYyJcdBk9hQ6zq6jTYBdXrd
J+S6VydaMnWFz/paNg+WyJ4l/Mg0IsDzCWWQqj76XkDBXverCKPhiuV6xUiwv8Ad
Bd3IOFw6e6V7NXZEqJ9UotEzqorIwbhwwccDbApOHuuPf9ABjCF7G7igurjJf6yk
YW7gbST4MZdqnAFQj13pfXnlaaL59blKXbSOkzdu8hten3MZO2v2bu85xE4xh1LX
0I8qElZ2a2qDuctbvAHqQoLrzMFyK+FRrzC6elogARbux6BhqTgyo56Ds7rVhfJz
bvzHE2W2CVVmNKINt5rnZDHf7DR6zZ8DsOP163qqgMxFiGTOO8kR6ycdmAESFiOD
9yEc0nuumQqZn02i4Ftc1qkbTn13PwoZzEijMKjWq8+tJzWOaNBSBHH4bexRL8FE
A2EAfA9XkumkyidLXosBezuHr0BtpziSyGAZz/cgLCX0SKQsmo1NphIcPSDcHvhy
w3hifxN3EiPlSxNzeWxJmf80VrH0PgZy4HgX0FOKA/GLQ6YbVg5vE6v3F6dml6RZ
/RHXxOaSsvvtzFmZDLR2H2FRdLKtdhLva7kl323P9xMWV3OOAVlb5JEikvXUq33A
d1SUCGKVowkebIiVaEVYsU8e4QQUjraQROJXAIC4k83zi7XKJEVnfNEoBcbC0A7c
ADpwpKhY7NXLRyF4c54h4BGNnvnyhpq1O6NhSoPHmOToK7Irqok6cCYDbviTvX39
BHwN4m/I2DNKceWHolICM1xH86LjxwhfK2rR6vS2hkv13T1C/vr/qmf1NgIgCN0m
hFDPxVZfCIVSNGmlL7ponexyC7kujClpy4HvZTBID/noLIiIqwfsJ1XDUZiCtl1a
3Aw8QC4EEfdOJPSD4BYCpv2+yBNcyG69bMLW1w0seM5o0/jc+Suvx3d2ak3adeCC
2SU7IuKkG1CpBeNv3wysdc2eYzfGEXXiiXNcirjqUcPq7fT82FOWJNqWKYPl3r/d
rX1FOa4pLcTR1h6IfE98ODxfWJbG9yi36QgVEaN7CMjfQm3cOxHJXBDQtAHxYwnX
qNsftDFadGK5utCKBnPOCblXrwq30QvotNWhJDj5hnrOQ3vNvbcf7cg8NXXamGXr
RGiREwxCX8D2aZGqiCdWW6i/3GnKa/Ycds1KglIIg8vdrhkAusgV4c+WetLWkUP0
gMfKyxpuvQVNPUvos1h7PgdWLmJwJ3LmGXQH471HQ+wmQrUgy8SEivpuPKeHuooK
HBr0jEg02/aYZDcK8nBhQmDlPnoNt8ZK2CbkHlkGE7PshRjkZJDAGeLsjEkkE8ht
mK/Hm1cIQyPqLkLjLiQbYIqH6T4AZCzQErZJIWfAPx0KMAu9bBVqRXAN8bdGsft7
60RkP6nLlaoUN15Nj2yg6g0eSDOudYmOQ8ZkBb+aY5vdVumgziQVoTNDWt2gfYLg
nbu/F83rrWf5P9Pm3fWpQh4gKJmHsPZqqPkPSuhBePlrMiPZOhSXXTYp5rT1RW9z
sIIJ/S7sMyzR+5dEBczF8d6hbubNm1IbKpZ/mcMuUvP7pykgrQ8J5nRMRnYP1COm
Nzwz4BgEjhWkOdzwsMvnZQ0ndvCb1c/G8XB3coRBEzNJyv9N99ewavpQ6jwT0ZAx
12Vwr/ROpLNSJyD0xrQ+98wzlL6vbGKNiRPb76pnCFozzxYo8I16Ibbrw7OluScE
7p1bVfjM/7mP7clvpZSb8cPE1obFK92f6QUx6mQ6SubFGPCALrdZWLp48N15eKEz
uY1U5bwp8alEr5sj7b2TDtu1Cup6Um37dCL3H1UD7yi4OC+LvCrjFT9B2CeDT3mZ
YsyLdAPFBqDLfjVsDvlnsgVZAHrI/gsj9BxQ5XTJpdlmsb8bZndeaUwJklgXZfZw
PIGQpQIsXmKLwxpuE4ni+vFVTYdpfIZwYUa4DNTecWoMae7p94h+ivxTy209jr7J
wNel7030xeEIDsrntjmBSRgsvyHVUrRRMYpAgASa3X5iZEG1Mzg0FaFoqedFRI+I
Ak0q3quZpPsmsQkbZKTR17eC01Fg127DtsY3TrH0bpwnLsv4ZljAwsx2phToubF8
vda1/ngG1yCt0AEzX1/g0fBfc8bz8UCkCypB41QMdJAXNhT6/+ZzEYJiis4l2RVG
C9FSkzBjuKEJV8/tsuaUZfxSzA+0JGV2OYmGI05bFi5Ycij7zAFOF9N+2eZqEOyr
1a7xZahwI9luFEzNqHzHLyaZ5yHh0B5g57OQEiSWDzwnyR5FHmUgf4boLlHjJQZP
RjiTCxRZEBLhXusRtCi2r2VXdBnVf+OKcESKjiQ8YbkSQQLqS4tLFe65MxskkgPu
lekHJ4Fe/h47aXUmS2M6HjFVsRpEZyQ5wINqAOPopNVrS51voZztX53WWKaTmm7g
jT02wTiR3cbAGtdToiJWABOzJDEfKxcUwuWKDcZsKPpjpEOct2lst7Nf6oUndWsD
Dnu1YII9Xar6M76f+VKP+24+58s/c5sSxMHPGun4ZNn+g8SBuQTr3RMboLsUapV1
03nW8OXJ1OZNMD7VjjuZjkQA7FCaKwgg2wLwPZSluNCDljV/KvR43JhLBUy5Vbes
CyJvcUmLN5mdo2ncIGxVTIWJPxupGx9ZefkZYs+tRq83d0NIuzob5erzpmrsIB38
Wca7BGPMtWTzr0Obc/Zv9+uj4WNHQLFviWlHpYSBdCWJEMv4UYvpVoJ60nAaeHir
b7PUjGBFQI0MaVzqB8qAZKn3GJPJnvt373p6YfG47W+4+yt5wseble7h470B/VWw
ggFh7y8uvGo5IlOfjCWHbpEPCWe0/95jh8o/8Clq3AGqtV3ttzcXyFmaiNCCMnA8
s2LyShMj3HrPuMKJaj/AJTwS/U36p4Pg4ZIqQw6fH/VgHFRwmcYqqjpmNOgkLcZ3
JEbjAuVBj9DJDuX2joTyJVo9REpL+3WNHimAk6ZjMmrjCpxciYFXG+Ajo+k4SAyg
hor4OUDx9zATfAeuYfeXESr1/5hFmUGTyfAsZnWW+6MC4CaX7HvkyqAcLHT+Qmvq
jgYmjrDJ6vUmVs4PyBzLOj0Sk5jHp9HoiKY2ksZe0QICdAKQwTqS4G4Mb4tX3bAz
WXkfIIW8eiSC5ji4H+aJe55hOxaQbAFKiFJsXBv9Up0hm2VgyeZogjrwnCEi32dL
BOQPv3Rcv8sybYrybu6G7Ocp8aSylOM4v1KVBrx5uwi5Q0e4/7VrEK+8iGzmE/tf
3XS1wkM4Sdi+7/3uQD6SZNYhSZZIC/CE5cew9//Vfpo0krF1m/J1kac2EJfeXpL0
98gix3ZqecPwYkV5yc1wDpIge+Wk1wO2yKZD9MABYu8VNpJNBPKUE/VufkVdUUHB
cG71K3Zx8jHM1FC2wJQ7QhcwPmWT1mLchbBj6/WypweyaiAZAwaS0WRwGdyqXQGC
nXp//448/LL4uyUgZRYPbU9oMDA4eLscHP3UwjoKC4R+XKCjnbDYaL4QJwPAKUAj
Sd1jX6N5oXRZX5VT0WrHF9iK8zTWl+G70SKnjqH1dEOTEsZkfO7Qt47SeRsgQa1e
WvywEizPR1YPR6o9EMwSctQObKHaiRfECNA+lDM8jGVs6shOEdhZPN67Jy7zF8zk
B7+eHUsljlwFrq+iM9JMOzXJXWaXU1gw1ITG6QEn0jHcxy6iqOk+wCLhXm3BcB9j
opamnyEZDkM5DAL/3JL4lgpFTuc9MbxEg5yDgBDoLzSE7zy61KvaoevgdPgeruHB
Ps7h+uPP2A9VX9QrTBwwUhDaNMp+XqcaeamwM+nKxxJD1XbuFndn32auRBGVZgyc
Zdk2fD7IZ0WlFCHl3UhbnnfegtQh8Zp51y3hn2CReEioyraDxfVwIwjZK0H4n14F
u/pyCWBkwekTPZsZweuyyWUHCxN368An95gcDGlXFgs33p1cizqTOXdLkNDr0TRH
XULo/eDKCaRT/FhiDvNm7PWGzNtsS3oj/UNuh+PIBgxTsHFSCocjInNQ8UoHDF5N
SuN8hRVtnsY9j8UK2x7HcZxxaz6nhvXwivMSgiOBMODGKGJ0JlDU+Dmcdyy12Vih
HsO0RS1gpPwzLg4F2ZxlFcxmZwpTnc5Zkrx2INkaZysI8Zw5oXowmM3VVQPBfNUq
RUAGYc74/lSGEivBFh9ce99/AB3eIrBfiouVuvEKlsc1N9cq9ayz5SSY3nwH3FbT
fA7ZNjiVrIngoI3MRgoi/Ef/x4QmLIXWTqde0Itt+2Q9WTAhM6RSMxKLRphxEe/P
jWyMg1xPvMCFFHRsUwh/4VV6L/W1UHVOMRjsKDo4hbrx8m8PfWsa+T0+EJqXAkIZ
DRQMz0jfpUP0yZazG9e9+hUs70bhAahPz4duKFHBtgAeZedKiD/rvOWisVHmgO9B
/eN6+4CpeL0nDBoDldA/LBmkD434vybDta8trOKwhmTOmW61lBI8AmrMJS435A8a
PDx6TSYkGs+pcw8BKI9tuj9ELOJChNwc6ofIKwV/nF7rfsl/g+AHfwjUJnxtwX99
y6+Hpfc+fcun9p8NRcc+q87avrWNCfNczIEGSzqngadUh1VfQLDYrQV1zeD3FR+u
uuw5dzFYPdySuJtf4A2KeoBNFL9u4Om2QdCi9MQaAVTUwqFNGqPhr5I58KCOI7Kx
hjmDP50clVouBOYgkLKtirv0VPyihgNM9wl56XBLhWewKCpheKjAMCFZ64W4rXAN
2sCEwPykyKtkyR8FPhwNcEx91SQQ3qQDsSGugrhjyB6ec43fBixeStSMm/cUdAqo
5PNmlbWCU4yx9J4mmdC77hpDsLbFxb+lV/L0snJ0ZyG/MOsJ4Oco8ceJjJg9INTK
iBoKOq+Hd4o36YXuOayLoyNMNN2raJQ7Ob4pGGTGS0G2Zdp5clROrXPbJrl3619h
GXbIsWf6yLtqSQygdgqQoPt15Kg2zHHw9HjgiaMdLiwQoJlqQBa74k9TdXA5U0KO
qC2WDcnSXQW2wmR8ODnDqa/eAoDH8FloTIAlK55nvR4Ub/2V/FuNDCtjZzkSKdXu
agQw+6oF8R/UiZqzRBu3tgYSfl2w9LXcqHahs+bF6M2tBKNXwRvkkVit5dltoKn9
V9Qt77oqhOnHo6E0iGsy/Ju4wYvn3LM9s7eR1LDxCxclslQZmSS6zX9P4LvqeTCw
V3bljs7IDk+ujh9+FimwqEBd0cXiQCj828U8YHu1zfZj6fUoKEzvQzJvBzu2yRgM
uaR7gR7l6UeR71zz9U3ayWIExFd+yoa9NwjNW13TFzgwUl5hdAyVGP397LWaVTiz
rwdqo1CqpkvqOUdnGQRHTHNnMitTPVVZbMNNH06feL/68eQm+861216HfG6EK/8m
PPzBO1oYdsO69OGadQ9vFTgUSJah2vn1inyogD7wfkqifbyuYrIMNE4VGli1x1Uo
1F1jrhAfKk/ipY/JjY2DYb/U/JMcU/7Ksxxp6o9+jnBR4OovnYPMZ/kbOHUzihcX
UGC20JePqw/tKBX12CdrfOq6mzfQSfJhecAIgHCgrzziqNn9v5sRUOVCem6Qc+og
WUlapjDx6xFE5nbElO3IDn5xeqoKraQW4qL5CCAygtCeDwhEXESTHHgFmTLgKc0j
PivwFTJxJw82eggKc0bTfp71RwtqWmCZj6MEHDXxINk/eiI15Tu+u/L7W9PDI1Au
ehLlnIAB183e52Aq+sKikGDxVo//o/lGBOALtO6S14LD6lVVrg5EerR9vTPMqRcM
dO0JJLSeHAhFsZeWwEdSLn6WO4xJ5imnE66LkwV0Ewltxz0HyjFucHffp1SHeERa
PPSIXoKp2oCJfn8A4tNxoBQ4MxFB2M1dW8lirokM8Jp2cnamYey58GUzrKBkkqIU
1jcT5EHXcIrXmLe+9fMa+iufUdxVHvgnFJcEgDbYsL6/Zir4cyPvO0IxgLUaAsRs
HCoiC/K5u5g4FNNdo5ujrdwMYYDlI/SlpSBxcETrVenIQB/8n6+qydS1UB+s8hx4
dBvPw12XZd8AXLOSi7Mr6pUyIbao/kjqZTJf4Lbfzmb158pFkhyokN/rf1usBjJ1
WaQa9cS4i0nKAIX80FGSvtGMD7r/4jNShaIptdceOf2pjtKfEYcMQMI/8Rc3kxcP
cn90Vd+S+UebJME98FGd2hUnN4S+Tyvl6Pi7XNug45QZ6SZ19nV5Rao5sh4U3A+K
j1D5RGVPVvZJ/vfzYt5XcdOd5vXB1K1lmreNSWIbfS5SWXmxnfNRgSBId9nitM3X
yRxdylStSDAC9rTDYvmXIUyja9QxCvp/p2V6eGDT7fyoP4am/Ser6T8dK+cUayJf
ua1UrCdQF6oqo59ZC7JQOuIzHFN11Yf7xXbyT2lnMBI5IfSYnT76EaLDONs1Jmbx
CjGI2plpFl8I6ikqcmYnJ8FptQBtCDeC+GB5Y8uG1FsgOXbEpYIrKmipuMAZtx27
hb2SV0wrbnDxD3VzmKkrF2Uvq3SXzViWy/VdkBkgpjkJ07vyNFEv5l7eSvyX8XqR
JgL3jhY1vn9u15qo+NwZdP43/oZpU8ZXxH/aKFdnkXDOtzm3+PWVp2nHyiyO2E9v
7EAS46Z9a4cQLobe5l8coo7yctKJIyBNlzpJGOIqreDz/gkvMVn4wSYZ6Rxd8EFZ
xrZ2jD3/QtdKqtyjEM1X4RyjuvWo2tgGjBUtRfPHKIz6srH8y5y7y2kgEDg9nLOK
QvSu+IEjhFOXFIpJuLbnEP/flbZ8CrWj3EVfJDmG1hIr5dMZWwV39rD2EDiWuICS
mlTCxI0Q+qn+KnUdejDxZo1QHVA7gWQxwFUl2EGU/CymyM2zU0WUpHYFaYMagUx2
/dd+aXTcPnlQI7plR21l1mDkckD7Inp89pMNvwEtW+U7CdZUaPr1id4GdgN/nLEA
h7Xke59qZFUw/rwgnynbxC6kA8PYop5er8M8HsR9ZrE+xwBncQI8S7FhCm2Cd/YJ
ZkBeKbzdxzrrz+GlyLpdDEx7jHl0O1qEJcaIPyrQdIrlqS44BDDUtUd/FdyNqwLZ
zLToAk6wbCnfQdiF4EraneLvSJ+Xr9HzGb+T8+W8bd6ET3GcFuxSmlMtFC3ew5cE
vsG5ROyy9xH18v3CIzQFKpKoY1ucEaBIiolWG/Vak4covaRVUh4xgFtxog+ZNVPm
DzBu6zE0eDtlqCVvd8H29N/j6nCHzTe4oMjaQZuVV5TqkKWe08hBLsYqbfrMZyLA
fnlURcv4QCAj6MWSoTO34BKx0CxbvnR5H6M5+NAX1mW5qC991TOS2eDddsjXm5Vq
4NVk1d3PE+HEzyO4XS80AjLpHzzwKqYdH8P4u8RAWqyzGNAHKobEvesJAUs30IAU
fRq4dphb3gkiV3+L85n/7Xx5xiOvazRbxaWRRF32iHDrMt7vwDSJ1xO2LjOMrNkz
nop+aM8A6cSsdN355LCYfj55MSFPT2a/A6ij3QHWTUP3M+M44WVowIx2ijdSTFMK
12I1KwKh6Q/ujdBwPeTR4J7IZTFgouFbgvCabXl0OG45q0xR4O6rO9Gedb3S5ZzI
rcDgNI+BPzpwvKgT0R41lgD7FdZ+Pk1S5l5TlSENjQ1Is0i7649i/XB9/y3MUuws
AXuERzuAVacux+hjOcsE/CwEfJQypTm1c+KlZLodAcrTrNy6zjH4oPmOV/iteUDv
Q+XJ12nsF6tUqBXAszJva/qbur1hZJFf6AWw5RVykbb5PVnI663l9dztnNSWW5lV
ubDOe6s/haA2Giw3LwSd+2/+diuDxNkN/IqyzdOQ/0TR8duuAdZtQ8E+YFPf1OFk
5oz1AXXe7DulDDDyS8lTgJkvZvq8AE4kpdA1NWyly78r253P19s9NKGlv9M7Wn/o
XoUSfUnuucTISnb3gW5m6UseaCvVcLbnzddLpE9wzrfNqxtc8YRlzRXF6aoVDrpE
xoZpLcLEGXwoKtmLCgD1dBOcSdQeQYEwoUpc76oCS6AE7m7yPh1j4ncDxyFBLk62
ce44sFPciX1cOK4Tqu6+9H/TYDwczqf566ypA5wSWLCbS/xPuMxn4ldlqOv03XOP
6K23GgBGWK6NMwv0XxwUV8Zbn/yxSOFrj3vpVTQ6NcuaJ3jiX5VTlA2E7yTGFrFu
eyggzkh4oApd710H7CwyYJWjmeZ9qhjgJKnqNxWLWQaXjz6Qt13knxm34mIceh0G
kalr5L+G6eOHciYJN119fL6vz0Pm+UD/ifo9FGx//ACCd+rcX3ltRT0nEwDtmQyR
MAutkA1Nf1iuZG3mkB5YBM+kKg/RVG8nX9wt5ibEtnBDDb3/vN0gzUo0s63oqqwb
Jh9Xua0+Gp2Zd7TzHemIgCIoEwOru55OTvF2+ezRs3FmoVec2f+YycjIg7ad0R27
rEj0hrcKBbRJ9KeVJCio+B9KaP6weMBa2V7mAQzo7B8oeR/1UJZJMqOKDgNJQB7U
BAt4yMKoW5oQ3DlV+RecFKl9wmVNqGz5HlZl97MK90LIm0IZMqVoDk7k7O20zSFS
SfbAt2IxDQ6p24RcSV44Ea7/ChVp9pk6Uaiq5ON3cEVsLX1AIsTgNOmTN5HZjz6E
aK8nV1bK+GahoqaoPLl4nCtRrQZXSMKu7vAMPhXPQnVpWgXjKzjgrsINPNLymBNF
8itZR1mcHteUQlvvC6qQZLFdlwj8rs71xhxV+UBcDgfF1vuGvevHeDqW5lDODqFc
vW6wtxSuOOd43cICLZVIgofT8Nw38XbIdSC/pdH2a0s20WjxUq2PnSvytwdrPTT9
p4HlMkJ9gTsqUiS1PcN/qzHlGfs1Ly1ymXLl3KD1Xbx5OmlFvx3frcngdEABH8OD
ABcZf1cXROX941f+3Fso/1Azg9b5/KZ8awyndxAsO5XDPkQPEuN7uZhfxZlH4px9
z6uOokqE+I4R5MaW9p3bLyNDmi/DP4VI9ap8R6vnHVWpqgDDC60S19YiYhhKDbn8
YLmBdWGLc89HsR4N4K9j2md2XSnvQm5ze+8YnxibSnOLUmMz0PQ10pcM8yBYFlXz
YW1JGMvO61gEgGScnDBaGQClh2TF6Rv6y8CXlHopiM728RnuuffFFTRWusTAAVKL
SzCzmMXRJmynWgv9hdZs0d5+R/M3qIts+vLPRHmjJYCH/xAZ4QWBNFu+3iHOaz7U
uqLX9NUYOTRtC/z03dPQAqsiC+W+T4QnQ2xXk2Jt7ud9Yalx/9ffAkHwn8keLhuM
qXb0KbYipf6LlZW6piF+0CmK8i+hLm+pcRwRtIf4Ogl2izhPXuyiSlX4syDQrRNX
VzBQPx/6zaCreuyfFnxfbxgofVbrh75RffQWXBizNQ1TAqm8rOTytD+18wvnvKbu
maqtC4S8Cn40E0vcwVyxB36QXl84kQZcqVhnv6xGeYPcgOIEnhCEy8wWQY9qo48r
b07o9VoAjfdf5OCyxg8jHdbHTHoAor7iBZdYeUVtsGQs/IdaQnMp73Wm8ln1DSaq
GUE0eTD9ZcZZ1eYpmVziBLAmCwXz6uvPqIvsiI7bpAE7/RZsfILh8bcjQhEhbPv5
VNSIWQ1YFfz1KuMFfZyoWxlHQXSvR/zVgrF+THJrVn1xhwwLZlvlTlg+4vkR6tpd
uqwwruGQfi9x1Zgg5hQ7lpMlx4cNRJjQGrmxTsLET/lUxLJcyo8GGMRY/rBzsOtx
6iEm8RqhbbCt5knhMv44zTu6yXIPxKqikNczb0sJaKxmkBcz9wLQ30Q4sQLbnThk
sJtR0iBMzrAxwoaixU0f32WYtNmJBkfaA3Bc43IQJ7UpiCioCdlC5SiRgw1cMTQp
2P4oas3EvXn3JylhBh3KdTgxTsY6j2X/bqYYAyxefZi3Xx+p9OPUsZR9NgscyS89
nbshyY6qFJpreEblKwFsJb8gHKGZhs5aJyktYxy7MaPp0/hmxn84Zqju9HEoZ+A7
PTrR4bRie0Q5vX2evYhEh3ryP5Pi+h61VRLA9UbyqKw0Ba3eLNv8NXVpTgajBm6R
5xne2Gh7LHw0r54CQZOEqyWZcUz+83+wwjzMeu26Y1gxBvxHsSkqVQrCBb/Zvofc
p6fQuswm0cae2833RYt3Vau7lsv5m1o6Jeye/IaXn70FoP0im3FU+QY12+SCfWUD
FBJmmZMzaUnhM/z7zNE+3Te0vvvyywHwDWxLLs7dpHgv+hRW6KzBY9EFm5wq4/aZ
P4IVzNkCdn0fiSExEM7cvKIJlWeDHEz3PDjxjhNxTSRLBP68+sm7TtWA/KTAhQsV
UJfqsOhGRqFw4l9IR06W96vdJZ9eQGt7EyD0QBzOuIzC1XBKmvWhjqK9Ab8TNour
vvJaqwP5wYL9dRYv3M08hARXihn0NK+AvGRgcZb4jffvRxQzDLGLGSNW8d5FO1+8
qGhvGEpUL3RZpPr9+qWVz0fxR/lqcDyaE4A3N/vfBGZWEIpSD50d/pibNfHTGJCE
a+ZhXtG44rIHvATqD142ZV47arGmDmjFHS1SJ9Bdt4DhuW86z/l6qX5B+nec/+XC
zjAKFLuL+OSfafNoycRI4L65B0akTKhFD+KD+/lJurS26n5E5bXL9mueyAakTt4q
bK2Vbb5yz03d480/yZl8Iyjg0gYQW91pfT9PGfgvIWSpg2ArOl4p4kKB8sQWyyxB
yh7PSfDVKFh/rQrHOetVIt0DJkQSHjyyLPyPFJQvfMjs0RND6J3fUrbbtHuao5I1
2YIYveVhOhnL2PK4XXs7fiYm6nmwjs/GC2b1uhem/nB464ZrrjxV89LVj8Afq0Jf
5c9cIk4SGap4zJgaD1IZ9+t9J3XpyJuVW9IagaeAvkFV056lfvXSwPnEtXcipO4E
tv0E3jBRtmzeQLX4KFKiFps6q8bcVf6dX+e4upOuGpJaucHsG7UYQrA6coz9SL+m
y1NRkKIULt7gjecU/ukL3hhmH7I14BKxQfirS8sdvFxK2fi0EUb/XReCAb4qRh3F
kSR2Q0fEloGhFBcOfL0pl3bIGQEoro8c8elQNyfMi54+Joo8f1+EPNj0N0Q5CLPL
4iSQAWDufUL7PDOszbMqmVVaSMYfWAGV0j5DZKblM5KaQwalUlPpEZ6Rca5QpqxW
6hfzJG7BtKWXOqBS+FU3dG+9Km8ZL0iwakQjfAuWiEp189Zk7Q7lm67Garxq8Kyr
aWL+Gcl16SZJMRbY7zNVdOeOisugilOa5uSyrjmmFHNIi8x+Z26tUGePuBHFxPep
m8BIbFhkLWjEJsDVFHl3cANUVbBmzFiFwKAojvEgl5nVmgd5vEnDfs3hbBVn+god
8Gx9OhIBeyG08ZshB9vYNXKLlE2tPsrGmmb4jA0Sd/fTCgxD1vqW/hVgHYlg06o3
avDKzR+JaVhl1simBZhoVwXk7BxXgnl/X4rHs26Mvhrgb359273eLLEqIRvDee8C
8U1aFPUipTmhFAWAdda1DhXn5MaXtJPRn+b+pHGUk7qgq6ZnWJd3ty82jFf//s2o
z2KHjh7xqn2BrGxdT6CFKilwOEdwHVwQDEsklrFKgVVyAMmiOnxqGmr14r1C+Cup
k5RmgjuEsYzeE/vTcxz9DwU724LEehCiqEHjM4kooXurScZP5w3tNCdK5vDlzOXA
EGWDdKe5ccggBj0ft+ZPgS21ManmMBZMolKzffkthfvGWMDM7XkTa+NkFqsMXKpL
C5rv3wNxctFp8PCL7ibtIl01XgyEPEpRyfzHRPdbWiZG7TnjHqFfzyrXRKVJl8v0
tLljlg4D4sfxVJwe41g9JUG5JrwRBAKDRQZJ8e/gx2wdTe7iztTN0sZLM3FHRkLp
jCEXX8ZoWvhmu3uYu6MpUf5hjSBFsX2fCPNOciTap6igMzi93KyA5ssKkfq4Wp3w
2XIbt3FdRcOjN8LOzuG2dRgi5L8gZliL1JX0qkWpgGpxmLobhJrpW7bisvq+Ct2e
7pIrYo4cji9KHKyvvJGqBg7/n5iOYwb7oTA8BvHYKkUMpDzh6JxhhoowkA5Z3Fkj
Jv3DdNsaidTq2ne9cnTIv/EsugildYGFu18JYlYJq34z3VhJ+qtlvO7R05XE3Vnw
JdVFUC4lP8h0Iijw1dlspARn1NBxmPgUUlBwbCB/wcxK0PAce2gL3JM7bYllS6Sr
igR74kQ3aQ/44TkaD8W/NB7e077DamYzjBoQHp2yyn6qO8ayUYK1roit3W0y72AV
nxtWGmaJ+zlmA2hvIUIlfzs8meWcXxvC+hUdou2c/t8u6W4VV0PVloJoT5MBF+1r
2B6/sCBWFeU08EWT8bNpxfCaxmFKPlzME09k/rYwJBtyNBui6TedKkirwXoPI61v
8vhAneAMAkAwHg2mFro4iYCPpR41QJ6sm7HtrLP1UcMekRoUtcAJB4JdamcbVGfn
+gNfM/5J6mnv4MJwKjNsekl47Yl/3HmBYbsRk6wSxPpittO/W7Uhow0l2RYCdRbU
tm4JK4gWKv1WPQYq+W0uwT3QWGoxl0lEDmwUld6JPpOXWZwG7PnPbOUDK/dstV3F
k9RY9WebL25LyFjc121Bu7fX+sTcKfAZjLFnLeSPFqrmH2H9hosOLP0KiPwXIqJY
hxSybEIKFymKSurt4nNcxJGW3tq+PJEahTatS/RvuUE3WQ/VGqYlprUpnrCVroWY
yEA7ABoWJa/ymjF+PkREOCg97LsMcso0kVi2IrD3PuGbEQPARkde3814fJbI7H89
SG4XTBQFNMkw39VTeRQNdpCVyyTZpwxwbNY1jx7Cr15e6GguFIko5hg6Dq6qL1q3
9+sKmmfwJfHwYUMjQ4peBT6IZCwOaCAmXgYw0tGh1mLXSJHYrbKIzK2Y8ipkMcDo
f7LlUbQufwGc5mCr89SAxP4hkzdhfCFKZ1K2YBJGpokq2mQEcB/WpdnR+fRy+uiy
Ykd+ggw4ikXQ0aupM8N8m/J0Npb4tPQqh/oMb2RRI3Syidafa8a7x0qsrjsQdBUL
SEqb+Wt8Irj8I44jlfM/fxZmzkf5de1zeWSr+dI8WqyoLi2fBU+7/S/1Lygxb2in
/DthAkDGntraJ4PT4Bo/MAhRDnS+dbH3P1f9oj3/Jwc3d3sG63cklwLhhMX5LK+F
CP4lGBeLdE2kiLvVs1VTAbZTGhU+DSSa5foUUl+TKeFzIG11BdfIygVYB1PhU+ci
j00kUvpCjUlXinQO8XwcAo0tRLq7ln4IT2OCt8Kjp3kamDI/0bnQlGzdHDOPPt/X
U3hiSO5ZsW+it8y5cMnWisFclbJ9jvorNt43tXZQpC1A+Ic1G0plqN+lnzH04Egi
je/lOeYsB3pHdmN4xAtGnQcpGL1nNqZ+zJVN+WfCd4MsJTiTcig5Fv8U+Vw9OABj
8b3LGgEbjwgN62pdQUGo696Xx7fk5DitmtB8/IL4Vtwc7xNEurl1YoXRrscWxT63
1rkmg54z7P4wF7wRG7bTtdE5iKbdGo3Cu28HZ80qZzchEzOm00VemPQN5TMqorBs
YhQ+xddWfpDIeOM5nDmpEoYFlIi7HQY+2rdygv1lB2N+FKe3hRHls7w64YWREhpU
rUdIihaJDj1a1AbqakkoaUSo8X4OofioblUPWjAbgqp7obKjNIU58iZqjbMHHA/f
gFc54+wrJnFdzvh5yb6h9rYiK9ZvnfNHpBMnVRgp9lHr6L1d5LMF4Iv0Txp7HU/W
Be8sErVVaks5ixzHLLHXvB4D+oI01eappyI0XMdtBro4YtV3Vsd9vtE2HoURhmn5
xqI/qbrfFw1QBdolrXaCRxpOkEDI2T0BxTEOvBVue96JEyWSLmkWezSqBy2/fhku
XyiZKogp5yvSiF4UU/paC0T6mc3xpEznm1XaG9VxK8LVah0TAAYM8eks5YQoY0fO
rjrCSFxCkexdpN/AiWVliSPZIvB/Hlu70aYDTTyblUGI9h7VY1ae2efVW5V0ah3Y
NYJoWYcHCmbDFL2ib1uOnVo4nKYaw/RhvWeLQ64WfMckNAV2p5WIisvkez+K+6K0
X9V6QxqxkLgOHdWFlPLNDPDHDVpJGej8wOhVbY0wOibnz0NFMCHMYjyZjik1rNSr
KlAg09WUiBOf+BI3GainnSq8pvFZW8RjZgRTfuJpkCl6hczGofVKGReny9x5bfRG
ZK5TSP1bPPjdMDm0ZSeM5edkcD2xYuKKrBuMwHbrjijohMS+gTVLym/uSudvKgH8
uS0yYfT7d1I2vpGZkfaQxa4vkhv9V/2/+HMrWO9VYvHjpHtoyO/rqAgF4TzLxj8E
O2Oqy0uW/iY7NDCMwiPtsq8JoOvna7g7pjdDAAKkvdb8R8If+X7ALJ5Jj9A8d5CZ
N5dsNfNqWES0MPIPJreoDLstsXn8QfRgrcLQLDwUypWpAyjPA8a6s64fDFVx3sPr
SWbLyNqnVo7aq9NPzplnwQK3fKobQiR/rlxuIZQHwAZNjhrXkjWLcG2KV9nN4sG5
E9zEK8IbQrl5J3cq9MlhRdLRsAsQ0rvYS/wh2kj8D+GjQWEW69JHXL4FNVqvl9Z/
KGlwWKxmW3wdNGDOuG0FyK1jN1H+53QLKd7O6mte+s61iLWX3PRATKbcOupEZlGA
EIpN0UBMsqTxTS6bJQq/skSESYaUaRo/z1BNAi/CWqjNSfOt75Z8UVika609GDAs
PRzPqfu7rPKtPXLRsQxoxL5rRgkmiBr+aNvsB7HfSM5P9RPTzX6pLDtxtqxQbOvK
/l2deZvBg5bUCPexhr0Y6hLQm47x77WJYyuHNRTcFQZuN4ZwmO1yIR1CX+LDX70n
X3hTPRCsgsfO94ttVF2ZTZeBbjnf51FAAKCklQKuT9WCM/9BoYuWOTbPVX2mxWx4
DDdJkDdVvYyLWTY2GzmaZ1zAtFn1v272S2T+SA6pru0OjUOhkutJUkbgrYHHC4WP
VorswKrcENG17+dMU9Afel0GFVhNgrzdI0cs7x28QAB45+i5FEfrXYY4/3LUuZqv
IawW6rjCxw+MoN8mGsys+8fzY0C2qlBlXT+sJXsQ5SHNjsScsSeR3jlqCssTxiwQ
Q7YVpxQS35ppZV33X0B8lUe9N/BRI/zVcdc8wrbxNH/redSYgAC9totfUzoeFg0X
f3QprfK9nLN5HpDA20GOQWhdrhMHs827oJB+/UfPpT9uMjwxtQv2btGNMwZP76C2
lysUcny1vC/vKln4T9y+Mlnc9LMuNpgngyyrKPSu91OawO3okHxzdwDrK3vkx1Tt
vFAMHc4txNXpR2uv/ndm2Ye7sRbWvFz5uU9roIbr382aBy2qJcjsvhdIBodXBcQC
aPErNFd2I9McyoSm1sjGe8dTPy8THQI5rjg2zS8Uh4elFq/gYqLUIrKjwmPJOjpo
u3BAVGSTc/hNJ8255b+wHWQNkVwvaZLQPceoi8gxAHSbup5y1HNs0zOtN4MqLZmP
g5QlnqzoE07qC8x655+BwdLkLS3ESgIhKExMFfGeg93IRRrhrHmqfBrO3GHN47IQ
NhKk864IaBaWsaPmxcYH+dIQiZESYoxTo+kAeI7ueXnRUZ9JnFyq86zVqaekfpzv
w59Y7wiWXvD4JWWcchvYIhFIWXqS5z4b7DmZqYyxikxL1iDb2RB8zCplQyl4yNK4
tQO/x81+2RbHFJkQsp9bEVTp00zoq/tc2+uWF/B+n8/GdovmAa4FhyatUc2XPYzs
UEjMFQIJlTPPOda7vty6wnho53BX18kyH3RfwdVYYDU6EgkLW5iz7LtfobxpV+uJ
zu7YyczIV9m4O2R7hWmQBbHDlEp86q4KS3I3bVpQ/RxOIkna36aYNteK5OVPV4ey
AuayVuhIM3Dd2XgmFYldoO1dvRK0xJPoFnRhwl0iEwd0hnpoDo98sKEqHHXaNjue
0XdJ5QkQv/3CYch3RUQ87S/6zTfAnyS0bCCfXxaCNxvaJjIx/cPjmIP4HOZ3Yl0v
HQgqD1780h4GmVIEh6tjUtbXrEFEmCxAAZ7TZO4y9HJG4CzOh7ZPcQUsANmQNo8B
AKSWDtq+GITPZPhw3huhAKdTMNsIhm4akldb+kp1IZD1Y6hlPDNKDdXPk5IUPRjC
3pp4K3eIoQBNgXMk22+3nRKONz/VX2oCEKzRGbJNYaMMQX4/4wJmdhJAmADHp6in
fKHcEBmhqVPB8iM6x5jhekTe2cYP6o1oB6GhYX42aTG/RfhAWRMDqvkFJVnCODiy
S+dB7TNxbvuQWsGRDAvuW/NFBdnoS4rf6QMFRLYu5Xnh43KNoOs1vNf6xwscyiIT
JzYP4ttLLXs+Fc+MGOT1nq/1zOTsPhPysRMx6gTQLWicQfIOx9e/zJC4BCkFypGj
1gpf0FZ1ZC+g5Emm24Wb0Tqpy2odYvTunuWnhrvt+n1AwsjPMFb9n+ho4DjhA8gO
wpzHqzhJ7JlAO5VHlAGp+9ru7ezbfmpBM52387bGqgpXaQuuR1gzDxF2imzkd8vi
hGu/jd/AZr+D6po00C8L/jkEo50N1PwFUug4S+qGrdFYSsZoaLb3y6tpygI9gIi7
lUtuhRVO8EAG1cZvM8uKzowFMe213XForWpgaOq//NzaWMJMOKT3PqIZgpCLzoTB
Uo1DR5WxoKkLWnbyOU7tBR3736vnsn5sB54KxbYVpH5Sr1kkkS323u19owW6QJ3K
HdXouNFC64/fSPKZrpnIW3ayre3EZ6X6r/keHNk1fDedD4yHAI7xO+2+x9jI0aNg
8tinYQH77VrLK+iZTuHd4dFezCvbtjUbCqODdudpwA5XuI1PO0/PGifw0M5QqJ8a
vtNdDRJT9BxHLajTmRFj9gsXDq8TzNpqNnGUT9d2iMbrfjNl95yORCncBJS1OWEg
n6fwcLQb/LCaNXjhOxloV8xVl/NfdB1+Lbzc4hCJZJuHUkAoMhP3apK/LAvHT5kD
l/aS5wgc1J2o9FM0sFZ/VK/rgSGLuoKCFezbtt0HIeXSnlUAOhZUyDomqkXnmBhO
OiAQX0OG2Nd0ojf6rc9BIaKRTlIfTKLIA0FYSVazxAXRbAMh60n5fgLRdDndqs+j
4E2GJwtf1/5OR/6GFlgaDytwcawKlG3xMQCRhvJEQ3ulHvBxiBl21IWCsgOy6iyu
4UEdTZaRNnQtD3JDJR11GlijDXbfoRJkFlibDKwlZS0K6Pow2OFws3zv9eiSqHfP
FNRkaVeGWJdPivwqsiOGwcbHVQIl3V0L724mHlro7UdaSMIF504l+UwyoW+GFHeO
y149pAoL4/VVOUF1A1fX3USxAi0ar7WtzC++X+SflA02Ym7nQ9+DeCPUlh0QMkz6
wWNhGM5JAwxYegPLeUZFxBTX/aOGaSXCKeUJEe/C4xAY13+lUN7F7vFgjQVzcb2M
IiDLN5lY2wD/D8zLpEfFHzWZIJp90Hp3tjsUIsTexYrliYM2GLgrwpldtQTL7l0d
kjvP+0ht2iAQj0TnCk6zzrMWqIF1IMyDUKDT9c1oD0Wipiz1IGCzKB6HmQ0yrQhs
LOejCTtwH5DGSYPXNzM8EHv6fS5cuiMD8FMY9Lum9uUCuA0TzjzK9yDnjR6ylTAR
y6lZqkZjAJZsluVQcJXoh7DKOof+ZcRGd9aZ8dxPZ2wRG1iUAJEBDrOn+b0KshIW
MvQ35kJ1ycFevp8MbZwBb+Zkx5eRofrJmpuAmLnuyM/5qvZaQrwLQVabvW2nrZ1h
FzYPXGpFDAUaPZevzHUx8nu3fSCUUOI43mcnotavNTB0SRs1dthYFhrLTUJpaQW8
tKdKSkcGBWRlnyX+0mBNGGDj0Vz2u5qMKwrOjeR8TRXmpi6qzL5t8noNU9Se0jkw
9AjzJiqo2CJIy3BO6qvvoz7IZVxGxva14ny7vVhMO1iWzcAINpwhaBNd4pDhcR+0
RS+ohG2/ZIvmYo93iXND4IeBVORch8DcI4FpwB13CnsxouTSyK7F5er067Q8ZuRy
WwPf5beSv0HkDziiIpycy4g0ugW21HAP9CGMqLaZkzQIPbWTMaH/KaDIpq50IxYt
JytsX57aAa8tVokIlDjatVSIE2nJJ/hJFqW/6FzCOZ9cKds6QTrPaudSuXpizYxE
rSuM18caywuD4X/xPHULj+Rqx4kitdiBJhB7fZKqwg+up5v3DGPn6YE0C0YeTVkE
D1THIMdorktuXHqkm2XiT/nh93gVMLSUJuEARFswbvAmLJXNKKLlNn/q0m+1YAHf
afVw5Z5xEsBYocoK89hdhAXLogkAj/NYrrlmABcqoZCf1w/DmhGayyOLQiAEKk8G
NTiC1M4dbGL90c3sNbyB49O23X4o6+k7vv4SQB4UFk5JiqjVWBHBZLq6swM0Fv7N
4eL7M/CWlOx/4XYBOMIH0Fu7MZRf1ypiIwDFjeLhW6zXAQ3NgJ1iPDnh/vLmCtEl
IgVFUu4wf9UjGw5Uzts+aDGyRKFpAhac01P3kCljnSRyH6/BCwKcivTp2pSBkNtP
fUn9m1ceIwibwLmsPAqQvgaz98YgwXs0NVnqit5Y/jgp/01cUtSDjBcjJ5vtwwl1
GsS6FrZ+qGsD0GeoRocqgMn18EQxM7egaCklbXjFys3LpXnPLV7y6QxWySLL47yO
LQzBmgZs3m8GECL1KOWkP6EoSLJ70GsuHkUwPM6usFkbAI9I09tRopOsJbzCyvgn
vLeoa4alUofgij7Uj4Nqs4HF/2G39suYX356oSL9ENoex5WIqq16gMIy1VMMyRuM
pEIa2VhMpjfTyhaK/qvvRJEx1hqVcT8e1WLLwHocmrA1LX3gbr7xILakCFAbg7jS
7zdxJduvJp9cQnhRdamX4qegNDp7UBlb6bZy5e30k/qvZs6VwsHtM+lTTkZkJC8/
g2RlrfA+pW4zpMDxJKRZBLtONSUZ9b3PNrR3wKz145ZnaJOvAgJP2Qnt/Cu5wqVv
rafQL1EYOoIIrqmzYxqfaeQYaC2EvAaEjk+IzSFBDciu8+2fqKofFu51E1ea3Mfm
gWTLa77GkpRFzgtrrGNpf03b4mrk9apFigF90UHnOmI3frAISU4x32s3lyj7KMrx
BCEa6naW6ns2W2gz0hsX5FYBlD3CmBy/tKjTUYmIxLSWQk5yGdaGKM/Xj92JTFS7
2DxKPwJEEXpTyVqG9B3PKNd6DAV3f30pyPWrSOybg8gVFGgptq35dR7ypAzDXCby
ksIA/zaC6us6AT3I02XuhEL3ALwR4ApEx52oOCJ9yH+alXQnZz0NVy2T9A4rjNRT
E0kn7gvnQ6e2wHjKg5Ppa8R23gXSCdzgfycnvsI+pU8MJm6UN1DZX95gpOW9Ctb7
X2b1i5L3DxrwAzCh/Lua/zmGs4u2Jmrb+46Zevvh+Ez/6XmM23vE6LlBqBSIWDsD
BlmXQ7kRAjtJoiMTeJ9MhtQIZ4SacBIpIHtXnnWV3/VNRipP3qCggvOCdoOxvfjH
jKkfxoOzPQGbeIO7Q4ML0GOqUIdzxRNhDbHL0403FtkxqbcPUT6Q8qlojJr0KW2Y
Fh0kOuJqiOAV14OqNU5DEh3L0DSbDG86eONyjNOJFYTilqkWtmUwDWpe9HD+a+Rf
zD49EzXXrMKfn0Cxqu1GqzHOKrS6KdkonjFMBwlF3cZN86XZ/c2l2C6YRlKpoU5B
CTtihrBuZnWWxPQptj7xwWG2lUngEuY3UMgOu1Czx1dcQdEYdP2v54O8ArPtKktb
CzhGZctl14Rm6djUncjN0u/ShpvPDQjIOQohpO2pkUYWRx3Q7A6jVYwd1l2hn46f
7Tq114406UA53mCXHdBpZogpuCDfOtatRNAmgwEAcefQ+Pb3CY1Do+2GGOlEWXjD
hGJtP0A06eyKzWP+CBu7PU68pTB8PzFyR5N4xBXzxe7UGccaV2z4xAFiqDwlUOoe
Zh/fC3ZKUAxQQRCy262FE01TDCurQxPc4cBtYqLPCjrqxfMb2+m/eY5clOuGoB1N
aYBqwMQXTwdTOVft0oNz9BbqFSPA3UeoQKWIAlxh52D45p49O0Tm176uICRj65qh
slKQ+dtd3e2TdmBMsPOBHIrQWiRCaAlIjGzIdyYvzZZgpgkj5qxw+3FNq0GQNh8M
W+XT1JSVV+ExkOrnvwWNdqSGXt44YVTqknEbQNgs3VpJbI0LMN8e+qGK9FOjZZQF
jbqgxWl1+8ZXMPQNJCmv5GU8eiZ0HfGSQ15990V5YySiw9uW9kjlS8ChjENwzEkV
bkFtLPrgGzlaT1LdOaGKjxlko9Jd4bHgu/JsD1laWhbG/CeU3y0ePrWm/ifaIdNF
e0J+60JC6+lt6xxIS1z4YQznWOQsIo3bBNGwR5xzQXGcSNKvd6eeSl0kLZT8b/0K
qebSlXfqdszqjB7n7cXZ/cuUBH9pbaVhOaGG6NpqHgQPqOFb+nrXuXx50bFoAb7T
WWuTaIuyezSTKZj6bktGsM4lr+nTbjKGoiB3CiJ1eiIXXPaSSyA1KPogA9ppdCpc
ldI+vOpjYM3ddZ0I7k8yIqfmlJrWDUXYqZwNaK8qKJckM3x2ZXRfvJYm+pBfNeeX
v25/yR+6B+xqp9c1HpfxsUACCSHZbCvm/K+Gw9QCurTWqymwLVzxFX5peRKruCzN
GOop2zU+MZfFQK2uOu+bEvPgO9cCEZ7oVhnkPJicHUCuaLdlrwVPlNXLH1n3i7UO
S8tljBdl3JY+iVJi9cTAXc204w5WmMa9mv/6rx9eROkG3RkI2pGELuG09dHPThyQ
vdBHHKdcao+TpNjQeR0lB8U8nee9MchlwhuTzIKj9rGfWu64XqCOHe/0Zc5KMZQZ
feQBHOZNKmBYbh3KX5aonNRMv6aohaoKkmN0iSATsUR3OYhpWLEKU/awtt6AA9hZ
Hga/24IsgEcQuTE02IXCsWP/p5kDzkyO8Uu+rvwgivhW6VeT7mzeE7SvCiuTm6qX
Zv8q55W+Ev7QjOPma/L8R0rB9xyVdS18G3j+PZa5AQ253G4l405xFXUIbh7EYF2Y
A49+f+DbDnAI5DRhF3TcEjPtO7Z3vF3j2CPMlD3AMD+lt6WIeVLUvrW22JiI9oWe
wAIeUKyvsv86sSSZHqzO/I+5UxNNLjBs2ewZsQFD3ymSZqMUw1ykmpZK8Zr9aPKm
lyykdlDlWh8t29GmYPkgm1b1j+Iqw0dsYGVZG0W73VRVYJXLgvTBcc5vqx3e5HUz
Nvh7MQba7WxWnOIZh2Kw2BugNoWxx0N5Yn93FkeifwMyE22o2QO5TTtjU6+9vaqI
emLlTNzq8VKSC50nA31ggJ/E0HhYXRldpJM4BVBYneZTnR2omsYtt60YQXWou1Lo
hV2Wg0ph67zXl6T6MfucSBkj1FLwLaNp0ez39Z/zuzYeMBe/0CZHNvmr43mQoJrG
F9/ELMFA0YIqPv39JMQhblU/sfWRGPV45jeuR1Y1xU1qUPrtH7cFUiTiHNhIBlzH
TehlfUAOrGwgZ0B86pP6XW9S9HgKwNchoqiRNpbBZ7xVLYAf+Wa65pyl20nJXg1Z
6vzzd3egZrCoRUtUglZCRyz1i0SLweoKJyhzePqkzHn296zaHD1YIph4nR/C8Xbk
nfDfuZn+gcgc61Qo+YhEF/xZk1kgGQS4eIZIEe5XPRjuPF0bryJQIzErpEi2K9tk
LDVJyb4GXjpbjYV/Olfq34CpiyVS9ut0wRYrEi5BIYGCXWMKA3Id5+88QoD33UGx
vjRkvjwEIDXIoShWUvP3ZiuwLYniu/sFpgmPyWglKpK6/7E7P2I0qrzrbHXzsEK5
i2nFz8PoDXJC9CicBgvOFU/Vf5DWhKE7iJ75LyfXkEv1wayNqGnpiazWYwM489pb
WTr4KEHRA4KGzAbzEWVLg4o2FdLXkrMgfDCqbHAzQ8bDSOxM/OBs7+/pbku3XMpa
d5VcONnv0ALa8QZSHUNnXSLWKJHL9ubWgerfEZ0WmbKuWr4qK2s3WJSrP/FTAKG4
r+7tOQYcrXSCtvjBnaaoDqMVW1h46byZBpH6XY0lPEQTrwjVFmUndL7wMfRx4Wg0
XCHSNvRzVmI8jT9yUvYjpyzcSR80R8Mh3X8w+wQyISQtIFlLgXVfr1pmZVKa93gF
GuUtNz8qqaE9fsDJKPBwyAUzJXhXcfTNT5FSf6GyNbcCaYLpxQxjzczPyNPHSe8R
GD8ykZ0+ONeVaVMjN/FaB4nQMykJpjSxx+I1JhlWJEH705Loq7jf+jEXdHPCvJRz
iN3f2nLffIq8gjk+G0i/7DkPScN6oP/fxZfP5YcvvcN60hnpzApb5CufEMz925w8
M4R8FAFH2SSPef79jW91+bJqJ+z+ADe/1NJ7+JZItEDuQSxLYlBIPSTyQF9LoV1u
lHefr7tWbXXO8Vw9xShZgneNB+e0qWYjxc8gGihwiapm2TcUUA0AcGyOk63pP5ld
CKojrZcdQMwi5SY53E7ZFCekvUQPkEBXrSQMmHu2KD0PmkFP98m7wO7lozWmq51p
HBliEN3COkLZGxt9keQVPofKOZEiQfoJs+XZfA1lXkX/CsIakKjxMqx/dEvIMTAW
ZW1HZv99EHGaXZdxPlyOK1bEh1lPSPA7E1CIp/y/OqkFhPHutMcrzU3WxJUNndUA
/h3B5fXjjmKPn7+xhsZPTHROXSJj+Fu3OSozkV+JTFWaDrMJx5RYxYM/6vT7BBzh
efdOl1L64390SVAV9J6sSEzHEivqcyoZ16g2sWAVDZqspWceGXgCPawBOkKcHZH/
49wpfGMOfQOKEID2PhJ4N96LO6P+Ps6qtUWO9e2TPuqXUixnFtMANN9hdcanOWK5
DxnEopBakzRZHDP6Uv1997H0UzrFTf6xXOu3I7mm/S24dfk7FPWbCJdi1DY3IFgi
1O0RUQko/x8EYhYrfx0L1qrut11CAaee7ZPNx4QUmfWg058fS2dUAZHuBAAOPJKb
Jjo60uLAKprcqgK7CgQdf1ZIn3C7L0rD95DJb3UZ4GjA1gBZo0qUjHbp4l7Yyxlj
XO0EQunzLA6Luls+9eu0RmvCyNcjS0XwPNyniOjdkpzgv+m7KahuKbO27NI+SJXg
bW54ZhucQXkJKN2nqUHp2cXTM91B5HGWakK7jnqwWGHqm0++aefLbN+Txn/dBda3
tuhKJDDN55HSlMDpOGfhm2jez5pV6IL7wUsdbfLB/iNJno33eFuSh28X8Duw1eEF
6O21PmAukGNjhge5fyoESNDnS9ZrMD6c9eXI6p/zYKGp45OYp+G0grTOpcz75sJH
fxjogyNIbFl3jNS+TQNoVsWx6tWZaHZNGLIWAcDQLLWY47Twh6AoOe1OPjaaVOtQ
/fmdzRvPnlZ7ozzZvJNl2c2VG+CoaX1Sh94CPJHtCQJSeuNo4+1SaQ8Ql+1IXlQJ
TDaWqHCIJESa5vIbom5CqAPPoSwnFrnqY4IoYgV2ltIR9OIULMd4ELnm3yoRW56k
aWcsRM3gWLJ4QnDgRwcU5jA/JaTy8h7tf6eE6XpmPDuArE+RTGYSoAwxQURLTAFa
6dlOdSXpW8TuXDoLvKIxa8QNZfe5JdCEfknjhFmMLADbsTvmddpEbKZ6J1NFHv1e
Wgx4SLqgklTyyY3VNR5K+kxo2zre6koiVbO3MQZeGsRNM1psG81p17n3JjZX85UI
VxxSUe0KI3qZwk+IFBUc8vLa5IVZGZtwUiROBmUBPZHTuLASKYPZRsjnv5iaVHLU
jDH2glhCafuiaxKJEFTdahft9gdG4mWt3gqg6ztCjcusBqTymZvTeZ5nXinbdt9a
CAgCecwCCEcUXT9N+57OsgxSwQULO3UbxTkjCEhQ+ePIu9Luu3bTIKX4msavLGd3
z3Rlx0R/BbaHk+C58XhTllfncoPw/ltaxj26yZUyPcpCoodWXWTa7U10KNyuP0t5
S5EDelmjIe85cZdnorg1Y1HN58xjr22vjFU3WZae1fGN/zjrdP+sktKu7nYSOpvl
IwgcDm2pWe53/2NKArHBm8sXZT5j/mBlX0BQX5CZykxnROq2+adkjNa9qHs0awrH
FUJRzSuxrXFAXskEjvoA70QP5d7z6QB6xad8Vb/F72uVAW7uijoF3TuwU4BqCo2e
SHtXDsES63lTKuCCvfXd4p+EEfaIwF/CH1Gd56jknPMSUmoyyQIx7n9j5yUFzi73
d4odP/yTxp/zpZ42U/yaYHLRG96qoxaokIE+2jakwm8FlpgQ+N4JqblFzq7iLGX7
Yd+d8VKGDsYL+/WvsBtN5cbY0l6Kie8EV+cwzPk2pnWNHvCD+ZY3/9JRDjzKsaeF
DAf4U3hy6dZk4q4BSsE/6Yqv6W2xT+oWZh1VEq/SXkjFQA+DFH4AfcHjCn4U8igo
JhJ0G5pBVBlPUBqOL3HxDi1yRMjv5kjGxZHpk/olxOPgYHKIEnLG8Je0X/yCs4x8
eArdFoROVRelj9tG8Hgsj2ZYAQyG5YYlZKC9iwwOJ6iQH6OS9JpTiQbYDd62DXtP
Z0Nx+B/vZYyIHccmax8/tae30A/KUBOmczmJa07NyU7GGUE58WJO2FQniJycPgey
WSUmRegnIFb1f2vyUn1GSHsOnN32SsXYy4CvyFpZEXgWzfK7s2nwfAgKlTFNiiqm
yw24YWI9Wuput6eRAg+rrrLy5o6Va+CNFXFa/OEld6CQOIaWiCjFvzqQNgUUPBOG
9pd84d9vz2/NU6lsmJj1lTNSLmtF6SaNPt3ibnMhjmg7BQCUfAreYSi6+51Pa5yn
JPOSkGF8fzaKiOEdJr9yNotYtUcHHUqyYLgPvWoMrvMS8QpQ3tF9G+DVvKYedtZU
1lxkwVice3Zjci5AenhrOATbXJ7F1g4ehcWw7X4VAE+5RDvX1RzeQfC25K6cb7n7
2mdAiqOePOGeoEIk7eNTnV8RmzOD9jW4n27NBGaHjUPG5fF7a1M51byJ8UGv2taE
LGOTGcBpXcVrqsnBBXoZq+36KdSE7jeCbi405fNEROKxv/fj+qwAcn2CYPlAxWmd
CAxUQsoiuzmelVyITeU18RLW6rXTeGp8TjWG5+oWtKaEFAOO15Mom2GP0i+oEazL
iU8+iUwm5H4pdRJq2QvniLyWqR7ek2hwPU27OCMOCg5jXQG3Z1dkh1CVCEDMC0Ga
iA5gum/kgwH5aSscEIpp+I5i2/gd0AAxLUEWYVyQ8yyu6bMmn3vC9nNqB95N9k4i
cBcSIBlrNTQnjIIwWSvX67MHS20ajrqj372TTQAKF52pWsyyPFEQyaFyM5CIuRe/
H1KL6h3IswCtORws5RKQDiFA8kJPOKhYAB7gL78N4jcvjZtaXzz6jL7UikCF3NB/
SiNGcHtUqWqvYjAOv2sJnyySJeNDLuKMiR1YjecSFtt6kygBGlYyay2/dL1UxO3h
u3lk8ht04mxqvkAS9phjgkDTxmiZV2AnC62pVyufyDTe7LNIgOWQDRc2TlzAYAm4
eyhTHftyoex85WepFSDqEFBiROK2vIphB9VH+3/H9xeffU/EtlYZ2EwuBV3cpKxj
RnRCkKooDPsYHuE4qPgzwQnzmMh5qei8kqPlD2YUOVqnGfyUXvsWZb1jxH5iLHwj
OCtANgF0l1O5xjJk6WrG+TVGYnFAX4V2FPmdtpyXuSYoX8gb04ExhebAdhIaJeG/
Pim1JpUt89zBUeU3P87rRv2TIRK71DtwbTiAPZ/jnAGlYY0Ksu3wPjJgY1+bGxbS
uYu7I6Dfho1MpROjvRsz64fnIDrI/+KYLYfNJnCPrQR6LYQWlDcPRfFPWi6BU4e4
dbDFlY3fdPkTICkui8XMS09ZsoKEW4b9d4Eg5DDHVHLcjdL1c12t8Be7E/FTBsUq
7mYPo+cZaZmG1F6m+pgfF2Mj+dIuGZ5/OZutiJOkE3tsw/ekeQ9m6PlbPP6qgd+5
HJ0rLcNaB8EMfPhd4T2BAuSDtIUbZMagwo35qSpxtPLd1/sJMim6IrffWVsegZba
D1YrA/US4/D04x+VFiF/uYJmTLRtF2OY2OAe0y6ZYVLIW709jigFfeJ551SH9Ps7
jC2E+fyANrPJUpoKsfcaImfQagi5QKCiYkSLC1g/6o8Rzuu/MRsCicAbP13vfQCD
b33691jEkVRsBxauNTBA3pbN1axJSXvyTRUM7dc8V5uhUJvFJhSKYOZJm4IUe6EY
4TdGUA7ILPtUtEKtI7NITo5HFdi9pIkTsVBRsmsLv5juH/PRTyY3C1aFEC+H80av
VfSxHehcoptyzSjl6sRO5YSN6Rh5I4+bq+SWxRLACK07t20Mue9aAEs3BY69Viqg
cHARAqMwb59U3XrRvs2NQ7zRNCzoD4dVpaRngdkALLmNbPTxdiM9hWR1iurEmV/J
9JysmuBcdThrNO1oQagEbXgG10uFTx0l/5/OKOgfmwRAbsrA6mY7RLxsuvL/lSRn
iRgSlSZEnfjaM7rTrIhtTVBtYyG2DQLoKd12//d1NSq5MmrPGiAcuWmfp2neWHWL
MRehnx2Dv785zv6bbuRwGmKxu6C8Rtjl/VOgcIvBV2JUHA4ELdyYvoCAEB1n5MIk
uGgL/dGEr6zOphP9N3ij+F4K/YKr6hYZijDl0/+okoBi68aOyj/JEHHBvhOTDyN7
FlNUpT7Vscy9tGOX0gFAtJNsXyXzHn/jdP7omMqZ/1G5j1KG25tATS0I7wPUShlR
wkd/VyAXZk80Bcyx2faPsh/KHzhCGkfi1sdftADNRbKxG0WI4KnNamZIZdj4aIs8
SY1Kxh4yhtmPjN53rg9OeB5lJkp9/cHH26PyfXH4BsFekkuYoFcJi5qK9HnnT+Gf
qVpDccaw8Qykbdr7c4t6q98HLS3Bbq8m0AL2H6wECangnUiNAncWpawia2hsWVyn
oXNyFYotYqZt3tyVz2cyBUBHOuGpSyF2fuchE6PGWTQTmn+ebgp4CBYkm5Azxzrx
BbsXse0sjtBV0eHAfFWbxwxHWLVZip0CjrsvpiEPs9fS3l32CMUvV4QJ2/WMVgae
bvnPGBY56IxXu1Ghyhk/Ys3XwopwrOB/cg/3RnytMPzzjfEkjZK3kaL1otbDUgr1
1/rs8f8AlJ8QZGnay5uROpEPpYeWWuzK4hCQ8f5A5PXfKryezNPvIbQFcjoeObzV
dL4FEHQwPBbpFmyKCD91jnTRBj60DO+PITyDC7p2DC5QELKVF/iVOXT/q0GGCOMB
znY3xqXe0ZUMGoUIAwpHs3UQDCemGgMIyB1RZIBk55tG3bwZVF1sk/xEepyCZt9M
K4kWqT6qarwAPjzxXhwLkMgQlG9ncqWtukVkF3HRLP9nLmK2UwT/UtXF1q+OLLXF
5C8mO2E0vdF+w+B9LWtFG2O6SYGfr/eT0cKUU337NIMgwuy/3kl0I1IfeX6gvmpz
hHyErMnluLK+D2P15ACKVfpRXOo3Dc/fdiUVqUMu4HUoBPJaJ/Olojhp4pGeTpgY
WRLvEP3c88PaXnZP8urazjO0+UJVg+N1rbxOeO5XVccWB9SNHsZ0RbvNk0mtqwlt
TblPXLBqb4w6d0inc11Lx00ignpyVzqGHpk6aQO0tgbvOfs6EkLT1ORGmFCeH+oW
ED8sC69B2s4LOoU4yZLBRIRkdpDSU4BPJvbnPBysOOH4AoljBKJyUlKJFW2dy0vj
B3FuYHR1tNuMb+IM3goe48122QmGrzhPDxFobcvtVlohK/tdjDSxNR4C7mIa1dfT
Ge4oTMfN31OtYPJC2VEbDZopLJe+vfR8vH66LPVUBDc+jOkK208AQ1kHMqiTidYT
EjBuhOnxwkOUHo30BT77ZqCsHKtLLeBSWUHJ5e/omTVFxiIIE2UnVUiGpNYbVK+9
pKRAZRy833+NYtvH6vgWkL1mBzxK1E7lab5Z6bEhdfkIvp1X8EJvjQMFHvE0QQ9L
JcORWUqLXuJp/zHpy8RTTzQYwfthN+icWktnLAz/23QLI/KrFd79VdyGZocXpAhM
uBxfzsyoMeYYjcVhJ5OSaIYX/re78dRlQ/hk0a1P7zZdd4wfmWq+ptQnId5oUays
HVYNUpqHxtOkPxAaDE0ZFzago8Smm0Y94VPLbbTs+pIqNE9rd81W5DmMnVLsDy6E
doep0avdUZmLpxwqj1PEbC4cSlKmpER2D2DP6ZjyP7Rch3y3X8AZrZJiuJcQA8Qa
25XIp+HiP8QBznrLLwznUtdTj+lLug8cfB0RltzzDeKrYvrHh8EiqJP6C21delHQ
+bK47249L3snu0IeDLAUoUssi9PjA6zK0AO8tOqyFYULaqwUj8IhzEoK1qNEmA4r
Q3yObUjy1ow4R/lQ2oPUvC0F0jL8+2uL5Rg7gcMGbp8yMrAJyABatt+HAjmJTX5E
keIQwH41+Bm/bPo2t/shoZjjOAkeYeErby9MGYJyifKIpkqoTUCUUD187ppL0wcb
9mljjbtXARH9yp5wJKdvO5/Sk7H8zcgRLAzSxHMFfLHLSuN89D4H+bvN55abdfZG
ev/r1GDMrTob1129sYmCziS/s6pg4agRBA1TgXDYL3kjYw5V80llUGBxs/HX1G/o
TaQuCsz8B0ymifW38JjMaJrOfDXFVQ208R9sQM3z3LUBHLxhekrc3rS7F+FSfxOB
OzDdKHZodReix22Ndk6JAfisWsPhTzNVHnQkmBZEem60KRCwXI6Do0g4yuLR2KJ7
j9d/xqUHPB/rNgmKyo7foB1I7Z2w2grjaKbrscWORdPZopgRE0riEGBtcbaFy1BV
9D23yUHLNyQZxipI6pTd+3b1SIXLnQwqiQihJPhiUOl63nxscv70UbQykDZLW4y7
y8gxOMslxqphV4qApW+VWjHtKAAIAdCXJoSbincMGlSZWVOCjg3Z4XEWrT64Su3o
0TfiiZJnyt9OuOelJLywKTI22nEZCtT35iYaxux1/3kRXtN9J0g51cqu2o501K7P
BXolFKagjrNeLLFmaHAQTzuQZLHMVNCRjLXZV29Jo69P6U05gG3lXqtlHPL64jM5
Hcm4pjE10iv+9HrQ9w8gXvI7hui0TCYTwcsy5x8xHteAT79CdINwnuwtK5iUQTpJ
eKmwCUrJN5KFwwY5aio9NzCDiGNWoB9tCG+lY6qERcVPDAnLW0zQ8pw9+hAjoou2
ENq4n5xcXhf5lx6yRjkwbdNazCE1lbdMjhzB2r8deXaLc8TBRHbAFmqhghqLdgyp
oeuz/xrTiPJLquWf+I2hvzRyQNaLvVDFvd3zz8K5dnq5Mwglea8OZ2OK6NPns8WU
TNIHVwXQqZrs4v/aIxpd1IHtIX3PLwlUm9UehzKMReP322Kw4G9rsObuVbIWV4Fy
3pfFJ38HQlh4zw/4ZAjqw2S5+EcYxdkf0+6KnCX1igI1w2IKcbS2Sm67hEsxIcmi
9uY9LvtoeE9WlhPXc2g7oy1mQDAuoZN6bSqm6bk+NIf1G3T8ONlJuP4Yx9nFHfue
8rTrLQ33iSS7gQDUarg2a1fHMBBAmHP8MSJBjqpd1xYj/SWEzfNl4e9AymVU35zr
QbYEoq+KaokG5IK64H1LiP9WSNgI0dRBlVQHDETiYzQRdmTRZGmP1Y2kEMo0LJDq
WBJHHX3i41oa+ta5wjKrYT9cybMZdrNXB2a7XZyl3L2mVZ1vueGnBDehYYAmn7pK
vThutbDlIpvNZH3sDNfoD6pcKuugg0CzEysMkWuVFcBbksxOlyJFTJBuv9fWS2o8
6a7omJ7MgR1dzSgvwk/6a29kXUozEcRhh/gOmN8Z2kYWP/etqBUj8puke3yx+0RY
`protect end_protected