`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6912 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
MZ/g83zWCQxCIBtfOHnYyYp3T9H0lMiL1R6zBZ8GwR8TpWnGBwv+4zRuKRulM9+n
Z8fny5vxM1Rm9POuYTnqr5AVxVED86VZHAmsnLNtiY7QiuRMBfEaLaCxVMdAisk2
iaSqf+vYeulS+0swfU6M6wePC/8vjXypkxY8oUGRfV68KR9VAJsy9YHmogm3DbFM
DIX6rSagP+NbuDWNMHbWdLx7QT9i/LLiBHQBWTw5qDEB8tK6EmgrVued0AGqBM5I
ONCVSXM3sOKBqbrwquh1nSt6oWcWEQVTmrQuJOZW4RlpwS+IcXA61mxeSAfkyC/a
erMrDJwhdugef9GotoOX/BA2jDUo97S2dBdWtniT3Dq/vtS2yy9KbbBHCLG0JeYK
R36JHF809TvmZ+oj4ow5z9iTmVmzPRy6Z66v07s8HlmjiBFO+ippqMFfxpx4e1eq
6f613sCBdU3Z95cVn8xjWKUNUXdDfal+IAZwrEIaGDTmj2ZklLSf4LqZB8dVj0CM
2g1Or1ESXf6QpWKxeRZHfX8fmFYaFyY96Dh/V9yVSxpce9Ze7tlvewktU3yCmEbT
DLAXs9SP269TbQX4TZXMkQVQD43Vp6lYUA4p95WSQqSAnVLbjHPxmmZT20x0PzDD
3q38w7HrWwV+oHIhSsfwNE6sAyqb7y3cXo4qKjw+mSD1aVRvazPCLSQRx2wOiV8S
TdGeu/0Fp25Pjuoe3rFQowdZzJmEBYzMtANoUwJh8XVKmg+9LAk0oMwG3vulEPlO
wGGnmwLn/hXql8ZDBrzqGNece3bjOC+slVEQLvUd2jJ7cGrNnvMHk8bJ9XkaaF04
wwTPau59vMbNpcgDq0UH/6c1PDKYfMfEvaYlTLgNmLsea6FikWcj5cX32OxksDdJ
+9LnrvU/b3Qd09MDWoHxgb2ZTpKoEpJ/uPVaiKLm/l9NCYGS6JyqxSPuPux6ju05
mb0p6zylL/MnOeTEv5bnO7PWBUownR44R4rgwvdCd8GZR8znCOBul9Og8AQdTx/a
KwWte/k85Te9gs8AlxZePjCVZnhOqWcy6vGqh340QqSflFNyy9HS5C/ETHS/DH2g
JE+5u2nIrEe+xBO5UpXiT/tJirsvUhrZwIDeJV7Lojb4XWAjyVS6J9xktANFjlad
2MizHYuPluaWH6LSwBPfZjV6pE1aQQkZlzc5p9r4VB8tIsWCAVMulFzrZqxifJbL
c3s4sLnQAyIvSAueMrnCfQb+RuGGPYbjmMVVFDHZ86S3HBDvW2LKVoPa26X2Tb39
fqrarSz/OZLNI4tc1/t9Xh4Ekd5RH8Nnh0IwBg8EkmnUuh1kXOqinahVT9xeFgyF
mcWOCARRflaGpWD6lKy/CD2de5sHEpbAuTPw+ffE9tm8/CuF9PEbM84qY7gXGPJC
IhwF5VZPTz/MQfjalasqxjJctQn9C05gn2cd50daCa712owo4d1ys5e22RpMzRWZ
x63/BtxKe9kp9mAxnYGh2Fo48Wz8SCDS/WtAlwNGPgeRpaoEOHBcse6RcK6YOe7A
2foGU8BYimtrN8lzK55sfD5XmhVFo2/6vGH8THIMfag99qOWPhmKz+MBLyVylXXQ
2jIYylHGS9N6mKLVDy2mhg59DvmGGKDB+Yjpff+QCfJ2P6OUkA4D1CwQ7dIF8cSs
GWZ0wRHWQ7raMrFmrEHHp6RUBkprOgcjxfVHgXxIop3DYGzqKyks0t7EPaaX/hYV
yp+H/dNNQZAJP2VMi4tDaeolvnGEyJBwiXJby3oh8JmKRTjTqb3LnvaeDr5+OlDh
off5DpXcIkoUxsFdHjUAGfZQ94RoLt+6D+K49hfPED5GzFTm/1FpcO5FfKNvmETt
n9eFYAzXrGMt7e3J5fS4At5wgenzGml2Mdk1TG8I1InyJFVf0VylhYptLyzouyiO
Sdm8+qXKrHJweBK4u1LrgoKsRpyDd8wmaPsck6SrNeC/P/wmbepm7FmGvPc0eLoh
vpoIKn4mUJKvHHHVjW6i6Uw+Mq5SOyJBPT5tEdoOPqtrtbuHNv+YwAphEmbIoDN3
OR7ipYHwg6aCXVT3xUo759PrCiZouK7PYmtubo64A/yTcVJigJ5x18UtuZQhFd8d
yRtKvNDBO1VD1Qzl/VpH6tErWw2E5U7RM1/gA+Gr3TgGR4GjiCCF/+m/hpVCQMm4
3hOGnl+FnuX+UKilyilKfugE3oZFxEAbKool3p0wej/QccVDowxszy3MqCoi9hCM
FqJFwkCA/e2dyYd/DBWlSIdKFBntYqLLX3L9yoANJVZ6SKT+Pb6j8eDgRRVcxPdu
QYZnPzYOn20BwKxBQ6m2FLMgfQQ16CLdZpJsifKSenJIK/OMcY4bKIHftFKo8JYy
E7hqDmvHc7DwiPVt53OinDPNFOedj1p9ibHHJmCbjU9tYiuhFnYI4aEG9b34LJ2T
6T3SFDCBc1SUtS5xZKfPPoBqz1vNpSF75NSoNYqB/z7/Fvqsp+J4vxhA1IuLRj3F
+qjF+ssHqBSaYI8oWPcg8Pa0ynPkZNSu1afAVc22fhKwI2jK3CtAUCfT6CsO/fO8
vxAptPnEWNpgr2P1nTF6d0W4rM8YYHZv4dHP+3rOehSotVgQkafasROFbcB99Bd6
5htl9ukmVD5nHTmN4KmlSte8D0dthriP3hJq2w4yeX1rgYPY+Nho779haM2/ML5i
NhoLUWoBuxv0l6/e+03wTBXYey604fY4jDL8DGIZsPw9JoiBXtUqDYICjfKVjwhW
7HPwUgXrpP3jTtIU+3n9tZVnN6TnJ66bHzHi+N8obou86mF9NFqN6M5homZjddEZ
r0tB+2KBmmgR3eceTCW9i44l6UIe1r9zTfugSbA9dGLtitbc88X1MPJb+D+t959p
vHCyG3QjCU2QPZmPV8SU6JLZ4LT1LnbDCN6IAsDFH3inarUDeaJJvB06dTBkCtBn
WH40XmwyfhVRRE0iKBeygfyzqTYR1nJv1GQxuCzbX3bmPoHabugf4y757O+684VK
kK+eSW/R6dENQhoowbp7SL9LxwQC4DDteSibAvL2NEd4VRQHXDNsZqX9CZqjIO4i
uFH/Hmd2hn8qrfCpF5uMGimcfWcxRIUhyea9UfvvQ4ZTlrOWM+51gT5wiDGj8Cc5
V8bYefP9XSd7g/Jsn6RE4fc+jM/rUmN0FIwc2c2hUiCdTHY0UC1ckBYdxq5qUKve
9IZD9kRYns20lhzUwDJK81Tl2d72nEVsLhMiC+DaKcqfjpzo0itz7Ev4yqIrO7+0
AYCv6pNmDSMygm8VWAMKe6ZxTWzUx6rBFWoBaPSKQDVfW3RsX0EOk+EkVWfirV0p
nToFLzFiesBBsJETPyBBoLTTlAgeCeWjijejbT91ANixy5e8Wv3ylt5B6i2vscx4
h8J042q33kyUfanqqa/PTwcDZxnxWdCNfLNLz9BTV0Y5kwrqmeAbHy/BglgR9aZT
fXsUnOi6GI9GNsZrMbgI/O/RzZTLyevjgDk2r/nVw8v6P897jFeoNXXysqFhuEZM
CiemlH3Jyb8yJDKo5qrIgWHEQwzNnfu0Jd4HZVQuS4Mj96xecYpZ1hoHm6XdanjN
viUpbHxF0HBn1fYpajReaEkylyYUrHfloC6V7RoEcfvMOPxVE2gD+gP7LL0Z20O9
EldXybwWwwB4723GWY/+rIaurDGR2GdUFWhMpweXijlkzwJshYLcxWw7GQNQ9Cp/
kvn5wpTEd0/YtKtyWKGwepu6cDf+bMu5q0f0k72/7CsHfbH6hORfvQwNhOfx+EnA
8JpfNqb2jalCsDSpDCV//N5XxHG7TbJYwYCzs7H9MXmVucl/M20n6Omw7scubIXd
r3hprya2S7V/IPm0zq2wppXZn72vFSvO0k4nFva3eNIIF6rsXI6TR4lryw9+I9tx
PItobKudt0ymplgiNe2c62UHiJslVe1cD6NH1lg4a5A++b/cc8Ej1jIE+KTGjhWu
w5JIimgrpXcpuYKpDW+hZI6x6EtveWf23uPOZOLXM6E6IqlwbQJaC21SiPszM1q8
EVrNwPRaoIbBkHwC+Gm7xWytm0rIvJ2FNdZlE55NA5zjrNhV7S1SM/VZa9B7+Bva
AICdtQSTpWS44e9IC8Mu0PLr+i+FslGR8mSOy/pecPRtNedQ5fjlOq18d20dzK+l
TT62epeNgSBpUmLf4Kw8YVAXLpJjdcA1HnvinVJZeAzP1Vi/3Z0ajFkPvSgzqT8E
GuvafuJNLyXMqiA9esLSTbjPBuJdsEf4HYuzUwe91MzypXIwWFfpe5LFuoReTVKz
hj5alssveJvBGfA3oZdW8mojdj+zIWdVX3UQPzU5Ddfsw6rlUu4oeVOelC4Cy64m
ekBDHZ7y4CvlWX1cnXUpdfzxSu2h5A1HKaJzTSvRYjk8rYU1abjhxFu6V2l1C/jx
Y/uAOutSESEq4RIrTs7O+GEGbrmoL2LDh9wRF/4fZX1sX2sWpc3ZGOF6ZiJsQhUO
pkeVRbp8vQL+ftedDwk/vKyQ4WVvfdUtxAtNkRO4Ry94NpkrEBOoZ6pQPXDOL69r
pCNaL0seNrD6pgM0ZDLYYZApQvwlt1HcgSCO/SUZHQq6k1WWeAGwx/2uYcksp/+n
oCKEHGQ9cbTqtelLWqRLp1QKFMUd0/YZKUUgz1YmIOqWfEr1N9P0p6HFTlJfw+ZB
BBkoK5XQxFI8ccBkeXepKEzoD5ss90Cs+a3cHHzBC5//3mD1k23xWEcqZbSzuiU6
JLq3HvrIVn3KZclj6a5qs1jJh0Ngi3CaPBNTW1iL2EKe/SJhlIK84nyKZ5yRI3qR
cGgn/Ia6OJd5dkWABiYFvqCAKSJsIEyHn7zkCN9F24JxLDvZopfR0GGyTK6LD/ll
DGPMRdhSAoofF7IgWHolTrh649/BFH1UulMxvuXCgYbr0W1hxPwjdBU/SmncerJ4
MTvc/kCf1mmAvo4v3I8+yRnj+MoMd6Wdp9Vq54M+jtNeSXdOHL8e4Rs5Y3DDLaSO
3yOx3GfKjQy7Vi0VtfzSPJfSuYeGqcWV6Q5z5IRJuXSh/wyQAXC9tnLzb2nELqut
y+0/DWmcci5n/UlG55GU9Jio3FYZy24NXijASAAK5862GYef8iT+WtZPPU4IrRIK
mN5RSnTNRmpz5opEPV7+yqR49b7mdMJtrlHFpm6NqH4kj+uogtFwJapCMdARdlxv
i919qOQ7+COXjC6ylheQiMFUJIrDvP8xe+X3o4Wb5Moipq6fr4R4efD7Bgpa5SU/
pVCmw+prAcVrfSoAzFxL1/+q1B97xGsqFu3L1Y0S/wmFLYiOwdVsE50M0xM0Jjzm
cfnoPYGDbafS8z3AB4phz0b1LWIrJyKKes7w5YE3z/KsDEMPxywzEvk43+nyKUoS
jEZJck9fBbqoLLijdrHLdfPKxToB1mkmzmVvXDLhzk+zq0UKAW5HoO5wrg1Sn5IV
tm2kwz0Ls35AbT72zItMFQMb5xygahrJ2V0tM++kchO67YNEKhksH3Aez6FJ6b+r
TIMkIcC7hrd1NfoeOuF6wXudLlevSbUpja0nC3WJh8JEmPXqDTCFm/VPlxRk0iL6
h669XnVHjFHAdneur2GikswcrpT+kXZuN+rylOCI5DOnGiDsV0JmjueRxhq+BQPA
XqdL7qoSq++4kkX8B3quN9Y5cg2ExzLY+lj9ClyKWvCIbKtQY5jUz1dNDkOmc0ni
RCT9TKigk9kKElihHnwKn2IxtaU0+gsMXym4E+BwXQRKAMimfNk1O5JiDCHRocDg
iCu9RmkpBYaHsJbz701t3kd10rt5HzTR8V9FP0up5hFsj3A4GifWBbnGb/yl4r1q
YI7ru0hWiplNH5I5BpejcDjVf10Z7YLn1TUplIf4yT5Q+0iIQJgft9bujIqPNZ+U
o9cHlldQmqCxRC3PoX4/DQZOwqYohcsGioXst1VxWdIBi6SZI2u0XGZqIrvEqjyi
Z9f6AZBPJ3a0HoKObcghCBUAGBMXaWyMQb7ql0eHVH7zMSUaupzk0sfcQL8QTwW0
wTW+M5z8wewHMUKsmFW885EkNumqFs9QceG8VANd5Ggz7wBIteEVYBg/+ftuvYNM
bou+sFMSP72yb7YTshELAE7jxbZvwJV3CtRL9Cf6X2rkWluBWO/VSJwt1x3Fg6Rv
bDdoIYLKQXbK8I88PY1JCnB+LQJGuy6R6OC8QiF0CS1XjsrFcAiknHhYV7zLdOAY
htp20w96UZGpb5nKFVfsiJT+ZrvZEmZl7f/C59KiTiJrsRaF4UGkieiM1eQEOCp2
7F5TxvXBTNE0ODI+8PIOosu5VqXb7HvJ3yqbHTJLO7J1OcwMo5JR2oKeHxwYAPfj
Ntd/Mc5XUKHu9TScA3VWNP8EFcHbNaQaRyScQ288wFE4rfHWbCk9DpyMmCw+dVOP
aWFr2EIkWzSItS7lxXbPRAIbmxsrM6Z3MtzJxHiWlcgV0IY9VA9G2mgp0ZFW7mK5
PXQm9RAI8m9q9E+cEu2eyf0Nb9KNqb19sIOADPy40WQKDT6Y+U1Abqkoi9MnLiNF
NyeDv1VtZJMhSQNrHS3f9XWIhWt9CAoWPt+d9qYkRRZl0klMUfDo4FiiZesCd9cb
8hftbpXtNAXrxXeyuWdzb5wu+Z4EOtQr+AKsxSaDR88n6En2EoE9HncRCKFKdyKR
0nAwKxNh/qZV4UG+xbvt1My/gHxmZl50REpS+Oy6Zxuxq0mqcuI7GVNpMCVgfXtH
V0JVSZpJg6auLqIJMZiR4WmE4tbuWZNyo226/eKbsp7gdijyDML4hPvRJHL7bRPA
QG2yit+6zVnCDabhiTOuGHwMllKxOoemjbe0Vt7Js/i4515bPyBNMYhtgRNE+rxX
YQLES0pKpXTOQzggoRi+/SGpyuIOS3Cy6tSoPSW/oMm6SQdRY5fEjr+Jdq8wQ/1o
eLvhRHYrL77sL6S1vu1V5k+2PK4wW3/KQ0k+jrwsUm+wq2UNeNA4x9UU5Bt6XiRn
jMofSRemSaWAIPf9EMkVcljG5pQxHBOwSIapPp/azGGlP60CdupQzb0TE8//qg+R
SQU6Mg0fz8jr8MEG+tvgDv+oCarLd90/eEjNHKXVlvCXupxTua8FcWbjmOwsmh19
IrFcspexnTWxfwD3iiRdOwt2aX3sUjLsUvFdlAJ5zGexSZQN6gu/1xELTXmjOK0F
PCll5QmM4ljZ9T8FwIxs4UOgNh4h4nQQvX5n0k4K9JU69bpD/oFJyrWF8d4HyHaF
YlA2lyK1MG8lHMu8HTA/YjjC7/A/BmCPLfUu7thW1HXoFIO0wR/2LKAlw5I7iSUe
svxEinARILpP9VZIkPM7Oz6qy/K4irJu5FVgKnrlUv/2voqAaqw4sJ1pLXHgl0em
4AG4UGzJ6qJ7m5U9BaSmjfN+b4LXGwP4z2sK4G8tVCOEpwTtNSAOPnERMFBgpAmq
FhS4FvNIFirxhnhZacwuDleIZGPj7QnjYs1H16A0TGeVegkSxhnZA0XTRWpc6HGN
CsXWx73egKo42xmTtWiWjbCx/RbMTO81p8qzI0KM1mzMNpJTqBhiBsYUjYRsZaYc
g2PESSdk6ciyC8fE6Vtkrdw7CzS4P22CLlZIhU9JQRhrU3DDuDmQ7xwlDBpqLbAT
nCDkzzJMiSI33wnmUP04c+F9/Y/Oz8zjdLfs/dZrNNPGUzf7oUgw2rDkqud3SUfz
vBsNNlBb5+bFq+lQKAN+Jnl9y6m6UrPqd1kxX81IBf8vGDKzfhpm8TiOsJl3xZXs
dQVS9Cfgqozro0oPFsTe66dQdchsyuYejGFyz1t0FrFrbmLvwma/lHi0eO8E/QQ+
x/Y2PlaMUiggKXbv5/sICY7gktNCwOCW039fn209GgWQnypBBjjq+XlZAyAoX3nE
7bHWWERMzU5HsBaf3NZPhimiZxi3z7TeHyO6NWjkE3zD8u6ekgQR9Vt8dR9SJAwt
QEpoQ0pLl64CH0k6fPit1bAsMvRZO6i5DVhaUMQ9Yna/TYKpA2fiwaAAV6nb+mRz
pOcgNiAVPE7Vv6s6S4rtRvKFFxaKNbpD3eyosrnZRBrmj5RE5XydqxzHKeZWYovV
jM35+gi8mbpYcwTN5Q+Oh11sUYQGS28TxqcxBJcaByjZwALONd1URD2v5QbGC1vt
bDTX+8+fhwsW3dcAZvuIM+l2Il0pPACyfzTp54cvCqnxkyIlEpfYNEQuQqjM3jsZ
DkGAiopLGF46Ms3YQQ04jgbBUr3tHv8Seuyv8FFtsiviCuRoPpsDfgd56G2B9YF3
PmHC25OKEYrcmFRWUk+tH5503DkTrxyEBIWmLw6izjwFavPg14Q99qtjOQnkc4XX
GjvV7+L8m2KgvHgHH3JZluc1saDnxmgpby3RrkKNnPd7xPyEUf6U3FlWOB4cyGWX
2xpW2ZBxePIrmNlHP0/Jkpjub2ZYgonMAAuLGY5kM/D6KEv7vqIFO27Iv9Y7MXWe
tBvqFK4eJP3xKvC47/6lZ/I1+xDM09tYZ3qhnU8hvmMtothu3yfX7V4QMnL2chgr
jNpEYSgTM0edIYF/nrkWL2+zcqVV5BldEhKMRthUG9HxVN61UTWU9KgGhx3x1wpf
4fMxuWRFb9Sk9Ng1nHHPhS8NSYf8eEfNezm6ZsukNKR+mW3ZHSZ6cNgSvUDmpUXp
ipAx1PNTGlA7ozVzSQnH+sfQc30z2QWzJNxhHmi51pICxRiKRMNXBzfY8Zjfx/Yg
YMCdDyunkABX3CVoSWG160K9MMwsAD8E3HGtBm7DisrFFpiKPG/iDBl8x0KV8frA
pQv7j5utxEBbS6ARit+w1gJOPgsZVRdRHTcilZmuo9ZcTmW+OyK7nh0YgrsOYnB7
2JfCvbMS5q7knosyKamm/kD/P2ia3AROFlzsoOV9DMLRyUeTGuVHK1qLqQlGwsFX
ffiUncwZQqenoAykK5XcNPFDn05Rpu9K3tDX8TVDMuJgctHC1Fy1nogR2xJmxgSf
k3m0yqa1e3hdyz5NeK2wFqTnfhNAe7usxwgulSuJK3gGHHQjS5dYWrN5yTob82eX
D/SK5JOE2H6LpJfwav6Nff+jz4y6jWa0mxkbgBDkHDEu4MKx8Ycu9q15wRNMLbTJ
`protect end_protected