`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 27696 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpOM+H0ygprhIA+aH9bckA3RFqMQzAPcHlHxaMgl8bjo+
/4NsYvDHterdm0pHqy/9GWeoHk+O+LdpFEIomgYkknz4L6OXdZIg3/4HrH8r9DX6
OrzX0vJ+uhnk8x0Xfe8uxzGQz/SVjViGmSORKJdq2OiNlKZOfqyqi+hH3wZdH8DR
n6OK3UNIcLtRmF2INVrjT33prblMI4TAqYY2BzblvN+yvyUv9vWQx7fYpLfaEzAk
2AkzGopwfpq4LxlzIohS25E8/QmgUzaHI8MMr2+umXi6WBAN83W0lUbGQ+7JChyj
7SSg9/GhrTPKQpe1TWFnSpoI63YjOvMqLBMVjQPY4+8GCjsrIbfszNGAVhMr9nFz
i62jgNuA9ig+468mVVh7y0okOaN6VAN0ZIxqGV/Dcuk2XbVvpBvFXdZbpz2oDgtI
O/wxJ7tfKFu0glVVVrsx8Os41i6gFiK0peTR9JuKK173c4NDP4/ENJUB9xBseYbV
zpQElvkRrnYaHKLGUuf2MJJ354cH5bJe6JI5ylkgZV4+yjRbjwea8KlbVJaeZhwk
3U2Kxn4eWY0JkoinbyryvOQ/X5BZQjWTunk1uyvgqQmpZMMAjHLJa1TXl2f+yPmX
XDKcMdCw68dPrzoHXgncjmCHU5rYDYAW8yEBwPIIyAXhS/hhv5CpmS3YxND7xAw+
od3ECxxNDFf6mOCjkWR7NaNY3Xpg4N/v6/4+R+JhQs7wvileBrO3Lp8RuTYPObdf
8NPV9qPBCq9mUCJ5pEFFbemnEAo+YxuIDhrCAjooAKAJOV94SIS5WOdU23DwHKXf
yigjWTueDL6sTTj5HiKfkIXBOve0wAhSR2NicQ5hgB55IKTXRLxA4MYVd51Z6aJV
6jZ2Aa9jADF3+Wtw/vWUfC3/NKb2r9FmEva3rJx/x6f93QCTHpOJSnFiTCd1pEDh
iPfdkd6NhfKfyfML3U9OEY8AEn6T/uhSZxYQza20+SJzEd1pfFhs1DuFeSFcz/+K
Flq5PZIP1IJoQZoek+1T/k3+FM0tWerNbh0KjBZLYm8iOy9ZIYOeTBolna3dr4Y9
rWu+ZAf5GN7iY1VWlAzXcXCGfX1hZpTHpFGOF8AFrFwTVHr8Nb5PKDw/GbdW9KqB
rQWxGO1RQ2ivuWQGLELpis2u3QJKPsfvsPnfhBgIDR9jMYOFpcv2r9brFGP207O3
AweLKUNjA1VLYWvN1NtSe3dD3q+7qzYT35RbQbSvGrhGlNULFOAM/Sbu54Q9qE9n
tbJzLFJiawgd5qIan4tQ7NjkAnKWvrsjyY9UChHzKdjfqHLYTJGIYzZ91mw03MpJ
aGbdASA7ppuh2R2atPsOX9OFSqHM009+vGkJsMq00x4z7365GXxsmQPqXKmviFry
YwZcvh+/hXhWIcI98EO2t+BrocLUaJsMVR7O+E0tFC34BsG5D041XX8cP6pYbTWP
ufCL7uCLRsPe0+1euzN3B3uMsid4o4kE0zKzSC4lMTZuvHvsyd3wZ1KlYIQ6r1st
vKhv9dAFe87DVRxrhrSiwgRULDFXU0XKZ59n1Ob6eTW627etyroAzzcFks+xUH7o
6yQxt1mk4sjR5P3HrWBo9hEvd4kCEx+SUmZL3W8ZnU0sjWWIIGrbCp3X8VIX2apH
7Vk9pjLbz7DMLdyPZr21LLniZXQxo9PQwnmT8D0WFnYhlGWXAp4vWpLEdtXb9czW
eG1RozEU2FY0BMcPhCTN0kZofZm2+uBRatPBHTRIh/xaSZnIGib/mc152SeCHL+c
uy8ayS6xP55IhDrjamBAZ255YGRqmxE7ECTYpUEVGIXR5NhyfRDr2kQbTsTD6eDv
HRPLi2PyoptVl+5L4NfKGvZEl1L0y0aw5xhASORfnpU2PBqT4Dyy2dAPeViv8gyY
LWs3p5fB2oOEIhIc4Nd5Xw5n9ak9P7HR97FjE5cajj1FIGsJgXXXdL3Lj2y/cXqU
j3166/95ABV2eAjA0lY0Yu2AsS/BZoozvZzW63JzeZINWtlRTPUhvWDodEeJ19ue
EDHQSR7XWsCN55UgN9EsMprnBMWC8GLsB81TxeJlLreaJwQpeQ6SikwZova7rG6M
x6kh8F308um7dUM+4xx3HvPqkZv7UJAPA1K9hcDOg2PT3rWlPL8/Yd/Ft9g/MCcZ
VopFYAjugUN5IYtysqj4E8dbYfpIkkaP6GeY0Fhs8FN1rwVdEOPGEaKLLcRezDxD
evAxBkX7NsYCipEkMN65x04vGd+MI59t+l1UHEBBblxB6874P6+jFNEA2GHkMasW
CNU8IUjv+TAOFOPe0veegrtZPONSCtql0uKTGZA+CAuHFahW7oOhK4QWGLzs8Y4p
KHt0AYjg/iBIPOMZhh5joA5gzVFstUSlSEi4g3IytCt3K33PLchTl65ErdM7aBrF
9NbO5/7NJ8VVSpLf96J4q3F6U43znVfDc0WsTmBRrq4l3XF9lqrJQrqTrIR45Iez
I160KXoPU4xw3gggb2Op8V7eqXRyco7snE3hLJhRYy9JxDQt7GVx1UKVASCeM1Gl
MoljUlxcDhnmfYiJah1sOxPKObCM8923FnZAcnaTNQ/H3RNY5mcLudvWz5b49+Hd
MWUD1aaacNcj/dBKGGYdlyq+0iXlTHS7K0F2TWwAxEy14nmwC6Wrml1rM/m95nLr
N54aqtee5QWhHagtOIQKmrK4PJN6dumlsIN0VVQ0NeZGTgtf8baUDu1LDW0kCrVG
+/fXXUwEJ7AmZCxZVkORQxm41zkKfgfYA6ARDi1H045/OfcCtknfOVRl9gCt+yYk
CPivFsgx3LLxmO7SX0QSdzlk/yQEihX71n2bUPS8Df5tdbdE958sD8dBEBfSXEzs
+gv3sVfphR6HSSUYrpxgFTjk5uYL0L/9GZIP0SKLv31ZCCf+svDBf3bhfjUvCRSB
GuWcpMSro/bak/4UD2hxtTa1p4WZUclNAejvzDdv0YPlAORf2r5U6RbJLPNb5c3A
g1dF5wSq6Vj8akeUWeutlANDDWnrDyxi7nlnMJjNFLwiPrqV7+f0ftjilAwkXWyO
cX5bLFDA3Vtu/tsOwp8ocq5EqRgw3SDlQkR5/glNBSR2Gm2vsYtHOGJLQ2FHcV2s
1LOWtqVpPM+oAi+3APDbddeKi+lfeCHyGfaSHvPgdJkkTMJMYiJD2EFD/PIteuLQ
0gHtg/GUZcBkbhhYVnC7U0VsSPgT1tvZStfdixuadbZDbwNTbedKjbP+vn19UVCR
hbTzd2IY0XbydJVm2HfNKrhusWEE+UN/8+WrL7ggGFN9NCfKmF8AmyAD58NcgAzV
BV4Czz/psbz7vl1sQm9IOA7WEGCa6Z3LHHjEY3K9W/G8Ka+6gT/v3RROfLcckdDa
ILEZZtRWH0sDz/n23LxbqHpcHzJ3SKDAbtf+Mrkh7hlLW+RlQHWyNHXkW1WqrWxO
lS29Np/tT7q35dPjId2+QPlWZe5uHPC6UZaAiXwj7oDlq/CdSlYYRH4ZEM8d2eRH
J462iFjzh1vD/Z5c3Cbh0WAn8OUnpJWqaMQi83TPIM9030PBxOTDjb1kqtVyuLxc
xmBeu/BuvsUm9WUp1eWlgMs6sWboC6VY8TyUyYVJigMU6Q6hYDauXy+T1ymKMCfs
+ROPTadnkavqt9fafTTPostQsOs33Gs/sbGenoTRNn2hgLYJkdrAe1PANabo9a7b
dlLsy5k6NU9GM+lreSZhE82PsXO9T8gIL0DGUsf2iWH5Xhce5GvWDGjMK1ATNeVq
HyiQ2sirwh9EyQrWakicOBBJ56T0Acel5EvFYFszEcTC4mjVlV5HYczPprBKltIV
biiXfdVKOkXUT+pF3n7TH81H0V+AyWVXXD7X7njV5nx4tInsz7W9qdrnkHSfZTnr
jRRnLwxeAYDwhdfJMjFIPG7Zd+JTJ/Rq+pK+yXgGLJv7ArcthQbkrEPGNnn4/ck5
PTm+1HUNwEzxmAd8hhHpu+Ri4/fcKa8+29jnMxa7lBaXjbNJoHgeJ7NvIcwg1MNE
it/RhJpR/lIUdULlUAHdzFsXBwuqKqx+CvXcuTRlLq8zJBYwlKaksAhWo3sa6nwv
M/s8aECshLHEr4T8uU65XmvKOhWFYUpwHOk18JoxeDjMNY1dLiWLVvgsOKhLyRcC
x6ARPqHYsYmmRr9f6AR2ilj2c6p4FSSkNKIsO6RiqqJSqx5FLc1t0qPA+iIChtsl
I3UMTLmqHPQNgEULbsuoJGHV6M+QNKmyv30dl1DyTb0qzXKT7UvW++LoQ34/DlTy
08Xi7NnQV9GP6tQHq5gNYm+Gi/nDlnm1BLpBjzi88hkRosMJeWDHTvcjSxKJR6e0
2nwaILG/+xvHi1VoL+wr4jxG9UOEWlvrjbehKRQNBluZNyjJBu0zdXf2zT/jpWux
av/+blZxc5iK9grk9usGCmqShBw6qTqFT1oyfsj35UB1l8jTwV/vRaMXsqN8c9F3
9Hlrbx5O9pbUjshT9BUwCRpRHjBgo6+qKvGqGgkm+/mN/cXMbJTh4w8jOj6QaUov
ZIGJM4B+inW9aUBjyvwQTH36784PTmwMqB9saxHZINkKdIpxYDw8t4X246TB77X3
UjuleYaIv+OSO3cMff5mcycNV8hrF9pKLxnyew0Llb6ZzcwnCak/YzSxRNGC1HuQ
HUnO77/eVuuYarrSLyvEmPyvajealzD0j3wES0gGUeh/LDPxwaJ2NXe+3UEvchoY
1t8h3SgBfAcfwCck3t0vlNrtbdUdkLQFp581JFtEBZ+U0ELAGLvKfovo7oyarQU7
rAaaX74Z7VwVMDZQi591kgMLSgOLWB/KTVZ9YIZW2aBB8bDZW2Z+BzP4hZzskS9J
wJq0lMv4QyMTv2LutCnt+Y+Sa4ShZ7dGXcD9nZOSuZ4gtEO9n68LvopGd7h5dKDa
BNVZf0gbsEp+aJwI6Q+aT2Hv6oN0tX3qIAV+ej3rpGURNnd8zqhaV39uZnaIVsyW
LNc1wEboYn4KcQjjO1uw5QZRvf+qdRfTN/o2F2zR777Q6vQ8jJdOrxXJAB/1UyOG
3Aa3hbKKjT3E1dkWg0LDejYjO5VEudJFD4w17sQHf/nuuMQTSUY7D1miiN/ECuBZ
OAwFSz7AOJP9Ifd9la93O+45/FQTuQt/2tA6OwzAOTbGAs8Mp9iuvJcxpwnl591j
d7XuKiBq6ZKy6jTlayPI4VWxSFlunIdRsrfZLn1FTKmCA3E5uNIG4TV817cE65zN
r5h0OCW8vXi2cqc3GCk3HX8aqH31mCyVDwcBWnariJ8AeRECwECE58eZdK1IcyrA
E9DhWgWR5C7MujBpjHkKAZP67YYyLWrVDGCejviRcbd79FB9aHDdZmyOOytvSNUy
UsMDbo4Fq+Ml/TTZnFeS2k0HexFNF7pbpSUWTL5PFuzfgzI/8MlWpmAWErxQ2XUr
jNlVo2ooVbrH5Lpuxq8TCRzf/Qk/pOVfI3Of6h8AeP39paXjkIugccdLsMlMPMkp
xB57XfqT5Jz0QZnaO0rMJxTuK6+mQNWbjf0ultPhLyRol1O7KD8dM35snP7hcPb3
MGcIh8YkDNUcKqndJSJZHaME1zh9FAyJFbzRi4AZ+thKwGWtU4Wk4yN+KrXknI+C
xEoyZGyF4kBH4qrJzTifGiQFTPBRAVNHgiXwBQHmoer3L6OX8kIM4Sl1bzvJU+hH
0ILs124LX0VWRjOCzeiOKhjG89PDekPNGWTFwEQUrJuVOFGbmaVp0B71VE/8BlpA
/1aM/fsapRJiO7yoUmAFKmCZjxcKlFLDsOpZTTuEOH8eMK3cqvSpptMFvNRjoxET
Ppk77PUoBFakjYAomBeALasoTCQr+ilMfBlJnv5XdL9dA+c+JBjjmfWyvR1/W+Ua
EkRNBiP39dU2OgeSPM8x6AqDDO7Ghx6DLCUjQw+tl3xKqS90buH2Hdw7NGjEWNyz
R+rdSDsJ14SET9Q6i47gDZiP/YWy63SoVFwXYJQ8fNhFCIgD0xhzTeFcN3ikIrp8
WIuef586jSXfl73U9KlkFFK4Y/L2/vqTl3MnjAmyS663xT4h0FXo2sDx3+9bEqlt
sWq4g3mpTngRyyXJeTUsJijlyAUH9msQ5Qp0lZ+kC1N4hGiUULk4s2om/h65FHyu
arlYdbOJ3hcvEsLMMYP4iGh5d6M81T74ZlKBjPaLaynZV4kPaLG4VcCIBsJluDt7
zoB+keRJbD1ytfAjp6czKa1IiNZIlYnuVarxdbSs4pnkRzN5uS4UgdScJIxSsdAm
SRl01bHpG7dpQ7px6im7B58+Jn/zFufWglm1IaKOFu1kCFvLS+biMuYhyojopf7h
yQZWqHqVmlemNkxN4ATBZkVyP6auE8VuC9/dFk9UleCw5SS8SO0q2BFBn3z/OZrb
QqzCXaRhzjEaTTymo9P1jiPAvsCAdwdUNBcakF96c2BB0ziHs+h9yfNVIAD2Mpem
MiGY+BrtyOPuYSBCD2PvOqfcEQpgtuolLGQH5DHD5+62Cq9jYwa9qzEedUY12siU
P7aVSkbbIYxWR0JiazLp6D81lbDN/tMZvs8vBNX1KYtCgTBYSXC0pliYVGXIpv4g
8W7yZb6hHBUhv4TManAYvsHt9fISquxNzM/gevFQdjAKIM4tBScVerAJlmFoYZTG
WM2cOcmnrp8wYO35AbsoAPa7ULkAHl9ShTc/I2Vxwm0+niYRKWzGLfgxR/J6E/4A
ksEMHQHUR5lf9NrEPgI4aeX0Y36VGKUs6zq2X71xRADyjns1zN/4N+0ZXTjTzce4
8CIfwmXmUD9R+Vrt0kz2fpbQRJzpFBuq6JAUNKb1wTDinj9fWziHjDUHFk1B9qYo
b0IYkf5Z0xIqgl3G1a7+yLzbV9ckvGIUmAQPvwImP5D/c8r1HwT+omRULtOkryep
LMgSXfxTVqV76nZihHd7oLveWxYTwkK7DFk8LgDJOPQOslcShUmyU8n++kxD5kpP
x7qh/EyWeGVYZK5cVvKs9Bbbx6MceqrH0aQWC3jE9OHRvq9Ogb8KbvTprr+0Hy0R
P4Nv5HlXiloiiM52uOvCkaKu50fr6JV4uw2zZUqhmCWEWtoUHHnPR60+i47RMJ8m
1xXITrXuoDwm3l2eXkeOy5KyKsugIbCbkgJ0rV0G8rIaTB7V0Az/kh2gb+a1RcaQ
5ktTk+5I2S9i5/Z62ap0cluamAoOuRNmCCI9hoN6DbGGEyBMZmM4VqLF8e0psGMu
cUBXNhkRbTw4lInbEUNn6sZUi0ECFfuEhSIoMbygpob0XEvkBXOA1nTfnkixzHjo
gfjuhYzXHFhgwIHJ42p8In939Ui3ofNxFNf/MlDgsyFISmbz5qhHuDZ6AWryuWPT
eB8Jsk926hnAVoY56movrQGUJT/wCiKd1+MlvwczP0YA3UexSG49QCeMjR/zjTGR
rXolO8REed3hKzxkEkm27fRKnKM1P3o6GPiR47dMn0bXimlEy4yjUUt4mP2m3d/O
oc7aaRNASrYEqIVo2JdNt97occd0Z5KQY+fJvVWDRXWMQBpR2PP3/SjuLMvS3Tx9
P5TgvlmFCBb51lYApvhx7hRHiF0yc+w9clkdxWQRSRZIVi9lgOfw8yHigjRRDB+w
ny1/SLIp0D6Nb8K6X5k3ZnyVeNR7sc7Um0d49NWMweqhRCa5pubLR/FkpJDNRLxv
Jy73q7/tSL+RtuhSem2wlg8t5y5oSm79/IviFHJZBbF+pFlHL+D5vdl6jtmOWCFI
ZoF/bx2F1OiPo0ALwB5cMQbvYb3Ia/VYxLMHXl8lwcCQOIP9nsY6dIrVrs0+oVjL
x5y0KMHOPY06M5n0cw3WgyH0q/x5nMyrRUZb+RXJaYbdiM6bc3hJzcYo7YCIH/6L
LnRmiEOyqd4YJb7nLE8eBHEqmFZFtmTSyIDFmTZaeoapg+7X8ACmvOy5lQ54DcyY
Fbl4iM7QsLBDrG9NuXJRFz0cQlDQAxcILxFehkKUJsdDUBRHwAqmIG4oeqKZXPU9
W/cV/KVAC+BodxKolaUr6rPVDa9ewqIpUhxU0P7GYXepstek2Lcq965pzQGeP2w4
QfOPuPPhKCpw5Xu57E8fkaM0rgCXO9XE4Ai05BxBOiO8KoEKRmQ4Rez13aO9XZNv
4WK9uU5TfVkOpUVgGL1lUbrvyaoNpptLAX0LzzjZHLzgKc+MKVh1hmcsuNdoO5lz
+CFDYux9A5I98m9s1IXzAwNiYDnh+9yFmD8JHVlDvTBqLyUiwwBLQomyxE8g8bDm
tGmpdbB6aloMBuG+7kejhEHmnChQUvoabudFIVC6Q0yzzlGJzvc9zOAKPft/aDEQ
QzBbEr9MOEnb0XBZZH05FIqIzzGarNEwhsEjAqvRILGSOwnGBgXUutJBQr8QoWZ7
gth6Xr8JaBPB7MgNeMfaXiHvdQ/JDUz9EVBkyIxpUskrru5oDeL9873Jpa0DwuWl
agfwGEWiaOsk0R5PFYCmxXElhaVWNBaNHwYek88Rr2Mo8PdIKH6Dg1Kn3aWrqrXo
zobVNucPmIcqmG0YKQfQtL8ETBqK0Jpl4bb8I1HYNoSecR/OjiuQwTTEcW5fqa0c
CEsWkB3I6DUK2S1tPPMDopvmieuW6e/NEN5SvwolaDHFto0icL1DR7V9Qdxirm6h
g1ZmfX8oczN5AKVtT5jllUKYuN5F+j7h2gRCx9gXRPsPx7v54oYM6PA9XXUFlwBy
04hsFx4nw123ofmwO8S62CaM/T3wbs4FtPSE+0xLk0z/qly1cTfcMhPm3q4MoEnL
42sL7WX+DrCUYk2dTUnc+aYvcluugkCp2EWA7XkKOur7NAj3QBxh7t3TB/zWi2zG
t9tOruAUhSzURZuhQpABbMMzzMiO1gVNUy5Q+oI7LoN3pTPi03k1TgZzVsiPqGzm
0hogM1OfMwv8+qfDNK18XWd/jb/Gd/SRWXBCZP0ivhcLTOcNaU/pXxAO7Eze25UZ
fpLV/E+95gitQBAPxp3qqScYfHFsnK+zD+6v3aA9BJbjMK5ujSNmQzFKdQ8yp7xt
zLmLmjWzzx7aIokwKUqAomzZYzzf0gG1A1JDtlCltKm08MlD51p4VUSapwzpGnbi
NI0fFu4wyW/6cm5tOP7YdAQopKh3DgPB8zZTu9XfEjrK4lV5kLh8vn3xYwdluWKm
KY8GzRcbws+YlKm3/TuE1b06pH2BlCWYibRhWvrKWHyvapvLDxBDVy0bMM0HDFNg
MQd5tLU5OnkeljBN2WlSMWL1UHsAEVJdxkUsQv6GcSVxdzbq6z4qLO/6ugBEXeUQ
cnmLTTKh4x78zuPIFazzyX72/EtPIXfopqv86SgQaohjl0vs75fUoTmDtQdN4HO7
RB/X28MvPnXyzoEh2UGy2SrpLqWyA8T//XvtUFz5YBxOiKRV1qhaQPZ2j4eeHf+d
gwbw6bNhr5l02W2nFe4EP8+vauoabMBvIS2aaSz2JEu4Wyirvtb33bKb0dNJoHUH
y5UQKg6xMAy6t20J+mebmxzRgtk4dVHk59WIlDlddivPQs/QViKDqz5avA7rCG5Y
tLp7FrAwh8aGSbvc9VwdeNo9JQQKG7H2DNIB4RNhb7QHcDEAfASUV4CDEFlNImJ5
WVSqrdjimWUw9R+bFKUWgT9LXiPmzm6hVC6n4lHOKlz47RSGqPofQxYZjSmRJ+i3
xM84k5lNq2xnMFegQsoyoC83cVqFD+hcTJCsLq3/msod4nn82Uzp/sawu2QfzWEu
cJCp8j3uzMCmNo5E+JHohAr6VLhZgIytuJ++C8z757PNf4zYqspgKrACV6eJ2/Te
ZY7XIa4+2bTJJeO/C6yygEFCjAAF0JSqpCgtLUqONI/Yywfjkk6UbXQtenAHFGV4
FAWo7OglxKCe+iQ4BOuvEWzkTTo4SURgSbkm1qV2aZAwBNVQzbvDFasRlP+cHm+x
d7Lq4ZSIW8o7o2SwmMw40zvk0/3R2/sDqUiF4PR2T+cISotBi5h53XSLohpmtjR9
wr9JezI4f+maihrPfc0FyHDZn9CAMQ7wGLGvuJCw5eQu/869Yn02fT1lUqd4qB2B
LHmg0rTD3YMFFSl7DeW7+JRLo4JXrX+Dzm9g9o8bh1uDEdH/N5+sGBhbJSQz2q9J
8YZ+jiDs8lh/jX0duwy51VgMlIMqerEjjtKZ5YTlwsKUYW45qu5jYVIfLRnwvSVm
5z7AMLC5tswLxxhFUqaisjlf5gkH61xENiPDQUkgqK9KGGYsiYIdBs7v98F9VZGM
OrfI5mH7SQ9oZyhzdzyPDKBza38qeP9/+C3Bauflia2ox1Iu66hAB4+pekjWznqz
XaKDd4ab8aBN2n+7Aa0r/EFYagoOFpGQfXWEQq3/C93k5RAI7VQsX9J50t3O19Cr
kbPdNPA6pFLMvFAUetAZ/oyZ0SIF79uy/ymvW0oOVwDRgG0jQQMPthcDgQKS/WKY
V6T2lv9F1Nf9eClzwI6agL6xrh3U3v0oWnpG6FFODdzSctK7W9lcDOS5Nre1WTSL
iHYQQzwmul8Ye9AvZ9rQ3QAurOWPKbnlRX/WyBcrZwr/nVXV30b/LTMSM1M412MF
wk/MQjocmqBufximJcnKn7icF/zsNVOHewyBcmc/2WPAnZDEyLJE+kWuUcNb+EJa
Vw+rxorGf1z91vB+xtfA4LBZ+mY1u/w87SiR+4ab1OSemyHqamnluOdoBaHJ2a4Q
pnTKT8CIaz2ietHEdW1hyNgfKrHR/vEm793ETjznB3UHTGZ2LTbAGeUM/aP/waMK
w8XBPrqxbJT+2MI2FhmO73sS6EUEQNtJoRLtUNSJBcyi4361BytMurTlSR4jkRhO
FDfJsj1yH996tbmo6SkhuhAWT6JQSMsFs7DLqac7O6SJZUQyd8orBobdYw2KB19T
a4OiOtOvFOsnA2qJ+tg0NKlG6uUKePQF/2Uun8VpJUBP1juPmBxA9KiHRZgcIJLX
rjLjdEXoG/Wc7saXLz8dNFBYwskp00Zu/n75elcfjv40MjSBBqMDK8KhpZqmceTb
5QDOqUSTa/lbewhG2tbSFDm93vcOMuFIruyJXgf2VpHuHnc25GIGFwWmDfxkJ995
qIaqRIOV34Z2avD/cst9zC02G2yP1olGP6dtnW4JjN6m2YM2P9AuQq/afBtrf46o
oLMPiGUu0kHLq2o5pN/e+dDXGotOuloNxYdmX0wuqJRx+EyB2/LQKjs+g6dofLJZ
wLVZVkqZtaVtPGo/5Y/OQv4Vee6fCumrJhQHe5wsPYztpY0sCkiPGz9IYYhv7r8t
4j5JWCfeBw6ZTRZsM4qIOI73okTjrD+jD+ocDl99MTivKxbjY8ULEqlkYWnvb/az
AECcinEXOObqks/WTmPtug5VipywOwis3RkWQaNAXrxkBNsi65VdvDgiwTsMTM9M
bnci2Kx3gcb9aDEC6QTVDp/jMYPBx7bnWdb8NnJV9lOZLRtSxT49zZ51BemLPmfI
5MwDZCj4rTt+8YD6rdDnbmDhmqayZHZoA4AuCUkp70TQuOFPawl3vJZ7AwrtifMy
kiHL6/ytgnX0FYq/KAagtPEvmF3VYt0F2QOwlMyJ+F2z6su5WpS1xhW2l96P1OWj
W6yPqsXseKIStiFQay3F0xDjp05kHvoHVs4LzDtqpoIPrylNBQwcSTymbzonksry
4HouMs4vbj/Il6u9Sg78aYGeJuEL0bEjIIw/5w4Hgkfidv1HomduHZnTueLIukpq
sR3oormAwPVo1p7lCwupjNawjhfzgq8aIwbA95qIAaAHEX9Y8K9AcWMWxYzHivZY
qYWlKbJ0tsO7IIpZin2xC0k1YfV7B/fA+Requ72qepwQPZL4+k8FqH8zmP09ap4R
b+qeHkVW1K3RdzGxFg7+lqPzziOEmT+j99KXHFX9WUEAgPkLd+29ZfOBQDTZUwvh
YtCSG3K4vKtf2Q5fgg24wASLrefBC6S8pwSUOcgJ/leTj9eyFeJzU0OjG4o0DKD6
e7SNNE9LK3szr0afLlNgZT8S5+8bRLg1Qwww3m7dmOm4lrTMgh6ccfUCozlkFHL1
JILwZDu6/j+2V4l19wJUOR8iGapIFhyBgj6IVEiXefJecGVU3LppTMEplIzHjOWa
w9BtN65bU4mtn/AlJ69xv7ipD7SnrqQz568tZwrOLEI703N8XdBO+B7Ovlez3PvA
TDLX8QSmnD7KX1G5ILWGTT1yr3dBjKJyS1S6M9iOgYLdhAULtUVlN9s0YdAf8eQ1
C35uE17d7iHXqQbELMflMFF0LDpf5UlbYrzEA3TnCsvw1ygOJpi1JzWUq7vzQyI9
bJ7ugZg0Et/Q2WAnDscWMBvXVQyDkHLlRbYLah1awsm5zm/Oag7r2y6QmIjzslnZ
9pfUvVjRioaQbkxeEDEttLkHlWjTcDVnXTxTeWbA/ATaC3R1xVVJzPXUBdjQPg6o
6E34WEpYowu4UCycIGQmd/Hm33pchHG8GiQobImHa9Wjw85910yGZSNC/rCBk0wX
mOjPc3bWxIMYeznxxg2Kl9YTh8tgNGUbCxearTDMDrkuFCNHgDj5XYesS/aJntWX
eJoMUV6sCs8jvnhawqY++NJPSdTxfDEaAJKuHmEDCKv5pD7fs6Sbbeb9jVMhGjW7
oh9sWghFYek/lyiItEC8eh8SSRdrz2PbRYiVAk9lPUXA803jM2fodcr9be04D7O9
T++7QLuLVHocEcB+g2BWMdDHcgk22C9UNEIWxaYtZUu7tWXhf9MdCip6d4aKrdsM
T0ItPoSO80y/K5twyk4l7NBeU9d/XoLBKI2ZAt1ow4P0DJPBwAelT44+lbWgPjra
aI37VGFGG++caKVfcx/zphOIA7Tm5kr7x0NYpxbhanU4j2L8fFflVPSNrFPsg/CM
kceOIyo5hMDFslIwMkkLmrFoswbv6zSSgF/+Axp8MHCROy4XLiK7Kx7HrJpHUC4g
PEDKkU0gr3pF6c7inpoWoA4wM6YtgNhbg8V4AShFLkg3ZiE0AWsSc/4QqwriavdS
q2PVqFz2T1P7K/6tNcCuJEOgTjcpUz/bU0by+OlcOfc/CclZGzAwvxl+z/BjOwZQ
HC80l6lZv1k0qlwOjcYVppb0JvAS03BuaohJqo0Snmhj1khOQRTBO7KpRYkIV9co
v+57VNqH9Zj4Vn0cA128Md6dMBU+20j5EWsHT+iIQQiNq2kkd5c5bHVRucbVKX6f
+9djjUqAETW0E1XhAvb8k9oysgfOM/Tfn6alWTuWwoFT1CNd8/RhDowVtG4nXK9D
aDdsG8ZZhfURDW8wix3y02zntli2buvaLBUPuUG3yqiBFNY2yjcFXfqaemrxZ2gs
r4zfRLMd1ijMx1pSIIP/tpoLJAYxPwNgPAUAQ1i/5s+WnU69seXBH8O8ulWnv+cL
482/fZONQ+jt2PbICfyWnF8tcJrRdMP5BPTwofbnMLrgu+BTcHBySkP4CfF+EHar
4LWLcMR67ShOiihdy7vZceje9Likrzvgd9p4NHa8E4gwXlfxib1xqqiHJS+ybOGV
Gp0gqil+j9WPMZyQ6mt+vdJKWlpD+olW1OihdDxJMgOjrc/XCdiYskmCcxtyC7I1
9Hk3e2hEOFe1or4LSMQhfuFmJhTPUyqf8a9FtMps0F0Pe4MEWKiAEWQq/Cgk5FMw
sdQk2gvVwlydF1o69CEwa5FU9pp/UPJ/qNRCmLNUvMyTeffRkYdHGKfSlB/cjwPm
NdDt7l1R0BX2ugUr/XJCiaJX/uk8GtTazuIDkKdYnIhXLWZxi9RI4gDaxFSdtV2C
XbcXaEMCgPxw0R6z1f4g5iBsYD0OGI3mX0s05WvCPXSCBDesDhPXLPm2c0dRxMf8
3oXLxXijZJ0+RucJGMdLJdZxKjUumGgm5xTSQfawfIufL1S+OkkcCCA9ahlnpKpQ
4B+UfMckSmEZix031i4APHTVhJebgCygKGIoSa8AnIWRgFlAVfJ8nIpqHkbaQ1pA
dQIROOIa0mZWjBMOFFU6RTL2Y6xomMxqlQdc01IIHFclOhSuKxN2OO8iiDGS2COF
YTPurS8usGBQ8nd/bL7ufob6gnf/KHn4WCSoBmB5kBq0zBFaN32vHKZqj2sV2CvM
YCkk/rDJnKtJED/z7p3f8yc54gZYAuJiwBu89tcI3fDvhs101LSOJMrwwDWuJsOE
G9/4pw3AM/XzZL54HoGAPMKvYMx3vmukmyELoIEJeC00I7GsIBzNHMSj3l8CFuNl
S0/GibMMfHIvDGgKck2K5drIZ0COjwfeF+8cJSI8hCpeBJFjkktyCfb4aQO0epLx
20d7sc738B2QhQNI9mJox90MmaC1bJTwqx8aeVHnJNdwmWZr55d+rm64XisN8/Oy
s6dhyk2VZ6RLLDAzG4VmiCR8tlvsAgXS4yE36dQuR5o1d0yhOoDacIRiu4GgLhm5
jGTv9eP1CU9NaccEg0r2dqPP4hG/WOuko/Ve0sq1hfk9zDRtoAezhDFLkPxuexOr
6y2so1Hv84bY53RRTY0aGDuBvwkPkcFqPNNF41Lc6YZ6Sj9j4TkP4p0ysuG/Fsoc
jlXBDlD7tu6Yo9bXRsIuUW/fbdeUxszM0JMhJ/ZshmrPuovkL7cyCKfa97lqNIL/
zekexxW42uA9h5kAfN8qVb3hNVgnwXR3a/du0M8RxnBYbB7lAhu1U6h40hvzZcdG
uOIQPXLUnlQw031mZc6SqF/KUkXYX/Hd2vbeQaLcJ8BJcyJoSNmnc4wmcqhJNyu1
gDBYA8G22hFHfebUFARB/ZPJ9u+T20yDWrxXzWQRT5dbb+ToSi6eTf62jhIalmmY
Ugw1MGy8bPq3i5nK7kOg1tZGXUNYsWanhxSebM706sBqJfg0C5TtAzzl8tDT20Qp
cpj470R9Cn4fvbe3pYsrjGOBZZS2n4oAnslJXtHPAbh20Ehy2u1G4NQqxtCUYIQY
ueQ77iyAORYdQEayqnWkwMeEYL9BkbNhGUM0Ns7gdeXA2Erxv94b3n6zRV0AOobE
DCWB+nfH9KOs57+wDVl0MVRsdH8iIjXWyBSk4Jg8vgPYlmPQfKPQ5zAYUnPNm+Vy
nsTXHQoZRroB3hvdHp4HMMuYB6Q3atQRw8I0ydYVmHQJBqD3asJir+VJLtXa8HPd
WHqijfyaYcPYJ8BMo/nrp6Z/P074w9FikoEVj8IZdD0gy74JE/0omWBFId430op2
jaTaPqhsFpfAgprZUz8EolOVuNS9AtnLYKeo+qRCToWNzW7bD3oUZzJL3ZWVs90C
MfM7K/2jLbQ8OdAluWGJwMiXVC0V98yWdmstXdxrsXbVdm0jJAo2jNC59gM8IGdh
Jid96CT9qv58VPAsUDJgwbxni6A/d2MIlq6qu/GyK+g6I3cQJF2Q+z+MgksfCv3e
IWtT3l8SuXH6J1Pi+VAqKzWfjlV5cYFyGHUfg/XGRMTnciAiedxXmDDjdgEe0UsN
KUjkXPhvA3Fe6Ggca69WcbpaykTUgGxw7cprWTQdtcX+KuD3wrVi4l3TWtL5iZJh
FI5TPNENXgKyv2n1uQmkwbkuBydGjMqpMtFtmdj176q1lVOuUUB3qwX2ia8F/qet
5bKmOPAE4HCg6wvawt7qAMJXo1FS9ijmYQq8RmqdWLvrpgCHk3sX47KHMWUfPDuP
37hZE7/GPYiDCz8qQdiyAfgCT4xxcJdpvCA+rhdcQ1AC9Xm+E28dgFmfuBS0CXKy
qYagqTc3Mqxa8/w5PPXpokPRW538zzaKFc4EaNUb186pAxoOPKoiRaKSYn93YAw+
iezN/SXQ+SAnp0ot8f58njblA5z3xYWFlyRBpRx7JLdj4sGPAeKZhGuzf1VgeDIK
9+GUFq5O0eXegF8B98AUbgfUoGze+rkpL2uaOE+LIynDvt0LoSbUIg03RamtX3Bn
gRZB1zR/4flNAWlKq18VitAFakQMc5+Rzkyg/j7rKybN5PbZf6PLeDKQXV2u6xeZ
1psP2k4y/E2PtHsmtxwtoIidepmraqDdS+Op6Js3PHvInrGE2Vz/cjoZHAEbjCcI
T5iSguh/YkEfiF8CzJeVUZG3UTNkvDQulcbXm4fLfGAwvOsIzQQFRx2B7bR8PlIp
YfwpVfS8HiuiMRx8dM7h6PHK+WJhzDC2ZI1P10zGq/RyNk3TIo0FHvWO1z0nS0q5
GvNur2L8tKLefUm7OfVec21y9hVlvR1IyvC9t+M9OERJJz31gd3RJab9o9sSyYZ0
hZU66gBNQjFQRi5L9KW+0Ra1jL+xjeK2b/AddwOiL18ew+tZ+Jz8MziN18BwpYwq
v+rA+qT6EavY6PjN60VcLLs3ppt1cmIJSuoyblHzcyCBpAxSbK9LwXFoA9skaD7v
7IApzGlkElTCk/Se6rVG34pe7PcfBFa2n0hO+NylZFfTcgomSARByXcXmrX03zOo
1pdT/7OkIg7RA0hZxWLF6IllNXzC/cD0rYHOlJ0zGOV/RufZUOddT7kxIEGOZUFV
lfN9UrnBKRrOeuarSdUKyKlnV0lmyZyVEmCROfxSnktX7y6xzbFDn386s1MRUJTX
OBOvGQakdyFzssphGpq/6SCDgPsIrX/U4aY9WnMgq+R6aYh92B89Z8GUrl0+ACw8
UDfhx5efm9QvUXRrtzwm2JwPlUr3tGX57yYgAFcZKMH62EvLAb7DacraZ5gKkHP2
fuxp5NiEhvDpUhws4HDKGXLHalsDbxpSG/oDdlQsviKBXOcvP0ywBZ2XXxcEYUMI
iyMIkOYMjP70otPL/drQ7qqjPXNKLTwdRXrMC6XgEhwC5w+Iu/UkomfEpWp3g7B3
nn6rUMuJKP2PMjH6rU5TYoj+RMCUHT9ygDZTnP5l9FpJSSEEHLy0eMWrKx0FacFf
k+a8UAfhe4ge/ZFLhRUYoR4AYywNkY2hlymhFQlYzMT3y9fZtoyyt0AvwOafsyYi
3dfkh8A7B/BtGda+AaGQUb/dlvW5+xZrxBEYAMvhhJCe1fnP7l3mN/QhjfPkGK2x
e5KGBJFhuAQhuQAe4A7u5a3juN9EX6PTMWA3ZZqv+L3cG2Abg/934rmI5+4sDvDk
Z0V3yqdSk13+HgkkSAMKtig7ADjK7x2OJXukQo9m/dvP4HlIeU/xer5qECtSanNJ
jHWeb4uyCDcVpYJkgMhX+bd0xCBMN3/IWDe9p9geQpbbAli0TObLyxa9rAwcG2u3
0sjFmsoa3leUT5CI9zBWtrb6rjXr9TOs2VEczWSgGQ2Ujr231gB7pOR+zb52uWRD
b51Jb1/M+FTt7MfkDgtpHrYQ2tBaIZQck02tL/K1BmtINx/9IAXuItf7EHtBgl0d
ydvqOi4igLVynRb7GN/14KbpTTESFM+gHnAV8aCJAZjimrU0UQFnAqBzrSjh8PdP
FxedarGqA/KEBsdtUeG5N8Iv9FwhoVcXldiwRqp8ZQVqidADaddZMH+/jzDbqUH2
ec31tgtAhOf51fRpyaVYqo2Nqxb8lhWZdd/gm4Ghv3OmIesNDHuYMueWbDWoFPQK
E52J9mqnqkYQgoEB/ufvP/6a4I5jaJFsOdL8tiEfdBzOGgx9lr9Toh5UfgfSfnb1
WuMPMCPKsfJ93MlE0o7v9N7Az7rAFfPWnpsrnagg4avOIVnBg5gSYU1h5m96JgyB
R/q5icC1BL3s0OQIhm3jM+U+4LKtKswVg7EVbZa+MvanNzAwkWZTWUBizVLByej3
axq6A72lkRuRdy8g7PatC5Ol6UDVf2R3Ye2W1tbgtwNPCMrX31DaoQ4v3ETfjw7v
gZvBYiZoNpBrdIuk94AQD90WysW/6Z3CGvzsmIShb/3wD1FI+mW7gllNMPtj8HUv
/bG1cW49zmArvAO/LX7l5lxmUc0oVdWgX/gg/xeaf8+wePsmfAsup+tOLN2eWWNN
i68CGOY98XQPBfMQcxvxu2w/8Hyvj4NtodpRpBvaMq1be9ULXhZdjIU9TQrAMINh
rQdyj+F6J2lpFbIybDOWE+colq64eqoPc5vB1rfSLC0VfY5/kZ38LM3aSw5kIboQ
EVPO066wL4tzLJuUYqcFPM5gd1IDHsvcw4vefGwmiLLY9njwcHAr7hG5A4jPUkH/
sHloc6Vo0GWN/tLY1cEtVJxzkDokyJF+tAw5/iUo9LSiS9DOMO/WWIDnHKRvr2Dc
R6Bwk9+BnS0uSYFT/+Zmj2s1luz6zthqNJ5cRg3B+BUWkxOjEb1e4C9sdL6IgahL
ix0Bq8oGl0gobJe8JBuNjbQu3EGaghFekjsEZJFZFW86v9CSszJg6zn008w9ZIGT
gvXwwF2rWdZV45jYVR6VUIIsf1l8J2PJksUg5q/aqw/IJivcoLP2wwGCv/JkSRkg
7O3Ir3qxxZyaJpPhsvTFLeU/+mnEQyKuctPWXqcXWQnfTC4d3C5entkpK465J1RO
jEItXAIum+jr3SzUIXnUaXoAG7GOeK3g0HUrC1vmTbat0mUpTCLltNzLRUBXQljX
1CZkhlENbEPsnwrwywuYKW6cRobJzH8UvwuHDcs/rIZxQwBRqtPczkmRGRXvXKLO
szxUs8jW89MEzrU0mOCqhAE1k9yIp317T7IU1Tw/AG7XztbZjiI5CzMpWyKzq5Ru
9DiZXrxP3DMnj9yfJmwzylrd5eJoeH6tL/Vqfbk4dek23psA7w7/3QEEblXQYypy
RRjvFp0C7zzN0GhJsfOdQP6eT1mvxVMlSLsU+WxgZQGlBUwxxumGFRdhL+18/83S
JQjteOPCVWNxDTfv2aX7NRheli3PzB4QB21DxBANtNIOuRNjFmWHpF5vZRiRekki
Emdi9ujqmR+cx00MpMd7v70vwk+M0+v9Pj4XKfh2sF+iaGQpSfaNpBx5Rt1SMWyb
zHUm0k82YLrEs88JItHcKemTMSZ1AVizO/b+nTojCBuNN4JD7gxz1eo+v8urEBlK
rFTjHWR+LmpSotKT7uI2aNfkE9xeE2YfZnFB0z2948Hl9Lv7vQqMVcjSIYgQVugc
P4ikNfPhem2Pq1/YdnYanfNadbyzgaAQcxczATTqWikOkB8moGQgrzvLtH39E+UA
bdpy4I9nBR9ggM/7U3NmvHUNK+RVeBwXF4vppOkQuGVd42j0z3GFv0JfGUiM1Wea
AGVveMandH7o8IlVBMTOd/N4hKidaKtK8fcgHyMln7mi98aqzBpDmc5S8wK7Gq09
fIUbttbOsk9znVvdJjjnTvbB6YxVYY7n9H/LxUUQGXgclr300L4J8JWKeDU/83wH
omZhwQrEkC2Au7H2OfHScjC8nlSQzFutXOQrJ1mWbJeICaJ94kLtLAKthel66Hgq
ppeI63MTc0ixRk1r7bGubfbSq0ha6OG4xmtKmU5rYQNE+waKy84fhMhiIySdzxom
fBLirXz76Z/EOsgh6N3tPEvB33Ce1dFJjPrOsp5xhVZ3E8pKTKhvJp7t7qWM8W4v
vAraUg2oF0CMAX1s1RpMhUlcoWnOoxtGPXYWQDIfNnMIbKbWFACKwucxmeeJuben
kiP2j6dff7+s4w7fZYDJQGeQc4D+PxQ4CwZK23/+4ifZXvA4pkLgiGzjjmfRtG5d
8rc0+xRIoo2Pgs4Rw3NDR3pIVzdojiZnhsOVuNa8qntYKVtcS4Q3M3Nl2l0tKFS6
7VD7MNH8wljzh9Q9X/ZjozafEFOybDkOzISFaaC2FXX82vBQ2zwhWf11hKeBVfgl
aNaYamEC2RTFuVTGxg5e8/htqW1ajA6mLCPzwqKWrJpA8+S+UXDZGtu0RJFdEaWI
RF2YLs6Ka/x6MhgRYulrQJTz46m+FbuwqqIr2RgkqE70FmEK+oo+p+YzyyMPX9HW
fo2wWUGSVI6j8CHUqI3hif84tiv9B7xDQNAwCzCGJRauta8x1F8MRYTWga0/gbtc
g3F2P2NoeBmxXYYxa0mxDn5wq3ORjdEKY/yc/ffR4LWCJz/0DUpSe3jj2083KQgL
eDy3Lw9cJEs0XrkBPrsjYTBrcDcw0B6ECXye1I88XndOhC3UdNfwliIxgWbIGU8G
xIbSOzr5uTGiyzVWUmt0LCErAyhGGVattWLnS89dhYKr64x8qzec8P/1cncwYhYz
HP556RrGO8efeQhJPbSLblcvMVnrmvwb7U/4mFmApttZtcrgbMwOQyBeNly1P5CE
XuKkV1jVHs7CaYOsICh1l4skq9+L3+u7m9q8dcRe1mS3yXuiR+YWbPWGORL+E8tb
zJm7q9tuHC/3bd1uI7zT4MA7GXlO9WrL4tnUZ7EkQK6aQN5Ham/TX91AP5XkkR3P
p2eOnW3oPmGzcZp7CzlwjSNlRwFTK1mS2u6KXTI4O/mrGLC9QGVzI9xGywiaEOn8
WTxdO5hSYuG0cly44osshLRQB1bUHzu9uqAQWmcRaUDdZta+qi2I/u2t1KxHq50P
mrTvptJFcjTg0/bJ8awMXwp1sh9JBJfhnS6sZKhgG7zAYxmtpLeVfAEVHr9EUaYa
YCgR14Ud5VkEmm+NIdVQuPQoA+5ZcP7ZNhQbNn7S0DTn0wcDjv+R7rDtAz1x8j4q
wL8QoV+BptIr9r4t/6vGH9lE8id6ZY2SXngAJH74OFkvEhchAFnZc/QcVTTP437z
TKnrUGdBXRZKLsTRoqVJb57upG/Itlfq5xSx/yl7qnCpwSo89mEyD+o89ymgM71y
NF2UkA7fSYWaSOl7+JfNRfHXAv7p90l+0ASXa3irWtD/uQ2MiayzrUdtXpqOCBGt
6jU9OFPHVlPimYiGfKufvncKkd+7hDNU6LRHQT3B7YO0T74WOVfnInq9cTdK4ha4
nUB+F6Gz5O6kEVpU/FvCctK0zUUEQpR+mj53Oh2+sFZQweY5rnwZJKIUZn/5NgpV
yPbHWJqlTHyWxEZyKDhUXSuAD30s2q2cqi6BzfqlGxqDdbslDa1Q0j4Rsi3rW4rw
thWgw3rBEP2WtZ95itJ/nZOMGEwLOq2xuKMNkHeljsD63TGDgi6lXCW8NDHN4sM3
eJccdXf6RQ9oBhaIjvqleivOD5WxNDULgQZUnc3e+U9tJ9ZcsMZJgYzCmR/aSwYP
i5b079u08Jakmle9FJU9j1rMjfM8AFgEdh4hkFIUgyVZUhBaUDpjuAEEWLcK6aUd
xI3MciZRDih4cjMXaBMRsml15tLFv+YRaX47uOXIfIrreqrs4Ai29bbBzxcA9iKY
kEuVKhUfN59JM7QbAGicZ8IQTKaW0VH1WHuQRn88IypvaMAddt7yLSUKu9yE4Pnq
v3Xyc7FAbbab19uN6bV+SnvgGJRSWYucboUrzgUYR8O2R2285h6+xRKl1etgTd1H
V1hwJpYqldMa4fkmH3xc7w3k/DgBchVtLWjCWtxahfHm64cB7gGJ+iyU7TiPRYFI
+L9YWPK8dLdyIcHYWIgxQsTjtFNOB5PM4Wfui6JlqNIc3nv0gPCU4lPsABwylWUn
Hx9KoI+WIfoeaYmFpxNDF0CwQHak8YRjItuOUE05q5zsVqZBUM8htNmAu2rnowGQ
EjNz40h3WA7if7ZTKW5NdVj/Zv5B+d6Y3jbu2cfEYPnKrsLxiQKlo+lAd6ClFxgq
nwEynEqAH1dCK4pgrtI+3t2ENaRpOZqj4rTAQodFHyxu+MUhT9wgfm86mEDzloMf
i/X5KLVasabfbuvXmphnHogH1TpqAa0c6sRBGVWwBpo9pKfnjqx1ol/hXedDubk4
rBDeROJ49ZcoZ3yMVfglS4i+JJMgTr5iseOklDUkWOKvoprbnvM4HcEIBXIdxYqW
1Z0IyZ68veTd3vKqzokHazbDRUuA2ntFAS0FtcFqkz5fTLCJ2arUc4YfIMOa6DNJ
zDLVNaDevRajpvZ+L+4Eid7SMRMQmZYyyuw5U47s9QWeZgmVaLrjqfibNijeVI/i
h1ULsUfLVFdpbW3z6RKbLT0FHGBRX7Pa/OSDdYpQ5y0R0EIuGmhnYHd4fiFTbewV
U+gnVXUYnuImKUPq3VhtUGeWb6TYvSlttW7Xp2dWsD/bmCFHC9nWbyXDbb04bvwV
waVaH5bdOu3vdibFTxCppWxxWodk06KSHE8tACbc4EOr28FPGm33S+Bgo7c3219f
AT4w0yxkVSDwdPway5Me1N5Y9f+hujYZQ18zMhlQeysUSWhePldijnEF4ea/uLzP
9n4SOrFZag73Sa7TzL9ztt2C7a8Dfl6UJqwZcv1x+IT7SQncjYyboX0qu4+pXyP9
Cn6G5JuSlZbOsZqmCVTa40qL7Xi1s9d7iZS/miWy+XJAScc5wCMplVzw2SZtf7mE
cLQ9W6bCARJDVbK1kJm0+rDt/eMWKf2BHHKmPxLG0FcBSbbQdPJTDBHFQbN93dlk
jTkc/dt6jphkNfH5vm4at+WBBILjgXeFpoGP97lALh2q6BJZgPScyOkqyBrtSnB0
W4n9JMCAsZDhO0c7OKBV1IlvpMXY5B7T1Dtg7CeUUcoB1WPlYajdnD7qRpnhF38y
yjN9+VIeaoaiqJZn9sclT0zOX69wI4Sdr8k6Te7xuI5z70NpLlBRnyNP55XKomuF
CQo9wD3IHVIL+4a41f3tU6xUDML7g737Q1TDqgyuwsBFSl85ajuX6TBnFKYPsdOf
4K8+c/y886KO6HTRRIl7AIRrL2qIzgBtwu6r49nSEijn/WrDosG17F6haxP8MvyV
zbmiMkevrlmsurkFx/v/I0cvduBMO1S4pN+ihIe21B0GAgi5jBYEJ2anHXIX0e1t
EY3cAg0An3WDK7J1U5q+DEotzn/NEqV9RBVxJVfBSfqlX3Afbk3IeLzp5k6Js6Cy
dCX/a1ghVj90kL+SDTFbiY10vY3xU9XCEPm4X0CW8QmMR9mpGVmyA5GSns0W7CWR
C0CoK62ubMDIt7/GW4NNBEC9/ANOHuNOshMiA6Kuhwig0YRn+cX6/5SxvqvRDD6e
yLv9a8qd+BqQ4E5bYKrIM99L3UU4nu2/CtO2w2QgPQj+eE9R44NGhdxpwQ1IzdcU
sTvPwW9rZ8JMmOM2zIHv/B/yQdrWxgrxAQREet/8RK6/Pu1J8h+N0NRs1o6r8j0v
5KEEXX1lRLA3T5E5ZGjusKsbKqziTTYW3zsAvm1QdFK5Tltql0M74zPWnJ4crwb4
NhzuLblY1BrLTAkeLr/McWmZuuda660R9t5ch866V2hvEcMUj3I8DhkuTEF3zIV6
+UEPqU0K3VooTxnzFM2/CCGkZTl0J4rpOuMvksfTdLDvt+7HkSqRvEn1JzBfZwFp
lm3FxzBk1+ulQX72yRLyQdNEXy6Q/aTNGl7c2A263UYKh5s0BUQRQRY6JEHBv53+
LNagb6D27OYNPpfrbfEC1+WeKA93j7+L6Iw9RAzS5oKhiyZWtgfhjpT+Xon9Hf0S
j0/J4RSshJnscxaV7YTtmbq+KI9+HHybmbl2MrzZvFtbQCY3YrVzXlTU7fhpFWog
YJl4ga4Ey/4B708+yFjpg0Om+789B1NV8IfLYKSRlVrxq1w5YYgVpAk+WfALEyjJ
4gx6L8Scvt+prBvnQVH1mgeJo0OZGPbU/TGyVQshQb/pGgtnqYUTQmRbez6qd98w
0jd3C4daqeS3zmXX7ZnUsy7f9Q83f/ABubBM6tdMH4FpB9zBLw/xdhqPJoZk2JKW
5qOMbJD2oLZAMkARRuwcr4qRmJFDERXkj0vOk7PMClrssSoC0ayJcsnwfodHU3Mc
9ti8oHGX5yWpXXbWZhkmWb7Q3uaI7oeQA4wbGb4EptOrAHNCijrS7W0nbfVpushf
4js0lPSbhdKZDDTGgZBLfCF8flgoz8Es2vKQySjSiSF/FOeLB8WZBUBHi0FbZ8iD
7VymMClTnMAtMUj3hKIcq3lf/PqbvWNiO/lyq24zSUlotnNz2VFaupSBIZbrdxDu
ythGlKTgpilrHMEWrcYXbh0kTeprj7mxOglQDAweiY7p1yz78II79AuUqNv1gX4Y
VhorT+YPSiapK7DOCfD+JfrUEJ5UoSwHhkGhF+CaTnmQGJOUMsl3c+DhIyYRWAtl
YJv779J9+Vb9/Z+MVTW9KgJPSKyR4/Yu/xqHc8vkq+LPWUPJx8d+WYzad2q8WbdI
lQRVAUDvPVROOx1b5CiHEQsqqLPvWzsen1ijHz+ykZTuBpL3mx5v46J5iEJ94puG
2vzvrKsCeqvq75A9KzDhFi873rydmLSQGydTq7DGlN63hhIh7671eBBXXiiezoMa
6REHmTpViogNGqn4Jb9dxtTV+WN/GOc/mSyeAstbOcbvGPy44r8BjShhbdpDihy9
hT7DJRdQ1vf6OIUZsezU5J2C1VYTa+3BmBtTOIu5f+/NjfU7dWZ8ON4uWMZn0f7w
YEMVOE157WwXFqTMu0R+oQhZtxj+Rws+XbVMdf/L1SxxzfB8GpzyvEZIEWfBAEQf
63SsRUXNwgoG/wuo7OoEhQ6MWtTUzjuWnSa3OyM9qJyyr3q8gZWb3Bc37G+mdpnR
33L1VGbCrA7SF7pO3NALY2dXqMTjsCQ+p5y8SzqZ+13oWj5zK/yzbzPjILobpdyE
VPC4FSZ5Y6WQRcndgLR4sjQ7VzyiZd0NNHX6nSYr4rcep7Y8H0lhxruxVrL9PhQn
9TgmSthKjRm9Bc0uFVIzuEAKNAlANCppEHkJU9wr1CTGNe1KXUoEdy32eUYiQFnd
a3KhTf36+tilER8ncXM9CGTqw6z3FJQ5+KgdFrCqmJNHa4iIT8VWutlzx3Rtb46L
9dmkeSIDhzXkt16EFP1zJM79d6UBmNkiIzrYGQr7Tl/90Blhjw4gTm8XxY8+GLwV
MGxkoQMQzu3xCqNNS/knZnLBwCIBefdVRLJ5CtxrJ+Nildinvfk0B5cvRl3/z9yD
6JQcOz2k8UpqgI24aIqpsc7C+Yms3FevX80FWYj15cooJI+Y/rHuR/rj4Z21jkEf
0FXjrZSqM+KETwnUFTuJEl4EhrtydIdy4glqEqRh2tz475ws0RT3hyk/E7SEkPml
0eFCvHk3+waqVQj3XXaXywHLHXyU7/HtYAfMVMnVvw3cnh8Kv/8c2MUkkEFYsZaG
9EAeoDVxdIHYf0dzSs1sHkeEiKytYrz+uGpkhTV4FAsmTmjYguMhG+EuZRl5mtuY
0bI+GEfzpJAFloIqGjOXl6B6ot3mVvhJwH441odwhzQgWOEa9V2ux1w+97orUpek
IZJsA/sXyET/aF3tUwo2dNPF7mdOB7dEYtNntIouin6amliM63u4FLyStFo5j6+w
k6UpOzMNshS0swGVHJpj1VST3s8LpTsaUBoDFdOIr1gpTVv/bJepfKVuFqwI+i7X
NoEXSua4fAX7y8AbIioqeKER9vD9SSDM6OJwjBriEHoUJNlx4g8VhHI1KwdiqHN/
/gRnqahwIahcVItgkC0WBqJk33DrkZwuecdjb9tcU43pV2MkLodHVlqt8DCIQuWj
tKW0/71qyzI3aHF30JV1TJ3LQLM0EuJCB/FgJqzA7A8KwF1ojEELuq/g4BEi/6a+
a7Iz2Vl/stuStGOHq0GnlfxGx4CsyI7KzF6HX/TYCZq8VQRadKh2NB2ewFtU3Dsx
2AYh+8zcBc5YuJfzpGduIQBqSoU0m2wQQw4sc6iIpmuN1Z+Wso7Qf5Ve3My9DRTJ
Jj2xGqvDeNoPByk6+VzuDQv2HYGLArwM+O2dvB1MetIvv7CccXkeHmVhcJfiiY0K
xkWP9BeN/7zC70tPFa9YGSXcZG52Ltm6tpYbwvK/fgaxWXpxkkpGm/3IJ6VrvTgH
ZAKnGDj/hjHBqqZ9HgDzjVkmeqHwru82vF+3nF5MtiZJl8N0mQ/QuutRPIxRD8M4
gotUzYU3EykCq6JspFCO58eCH5GUapoa0KSc1cvsMpsYSvMy7WBho2PbuHA6NOGb
yjNsi8norCUwcz6KLSSx3Hn2PBmJTqwmFeZH5CdaDc17kUeDzzIJ8CfZYk7o1EEh
VL/io3lVIXF5atJ1khyNa6pEMN1McOqNznIWqbrRMF5r1dW/sGZzGMrX0AYJTAan
m/Vn2MvIgzEaAyXUE0ULJnXmiipESrOpNkr0CFl1ILSx5WlmoDTKnvOpw+k29hnm
V2SJjWs0aeVHS9ZcjuHxtYBkqmweR7AxN4I3h7DOPLUjTnn2LHNc2Uw+cJEc9zeM
p2Rys6UqZd+4HlguvxZPeCr1tWH2EgNw28srPInFRhidXOKsj3dloHdVTgV1ukGX
aena6X1cR6DKHXQJ0+Orh5/rV43/5h3TWZsUl0W1FOvZgWyYlt+Ika5bkBAXuS2V
D//x6GT0vmv8+5MyE/GL3ZKEXd0EYfaPSNHtKQBFqx7ZNVyIfuOY5CihKnIHejVw
XFCRYa0N9DdjE9IrNH3fmU7EfUkE/0Sxocqf4dj2cfiObq7WGKLSDc4dsY2hmGkG
9ENXID3q/tUz2FgXq6ZdRiSDpqIAKjdOsongRIr3IpWUvXE27TVe6Ys1/sZY44A+
vtxhlQ1/i4kmcVGxP2P0cXV9qm2Djv+Ye/cle8lEMxFAnmCAzufnK5aa5vt3aVoG
M0OTqPYN2f1xWMtRUCHyOnbBoHpf/STN05dDdNVLx7oYXNtFF1E+malgChWufPo+
qksi8Zk4TRsPEPQqmSc5q33+WuLgiiKIJuRcUZA2wHdjEtUqlLYPQbyxaAz1qxz/
gCg7urnjGcqdlbgWXYu5V3jbXPgQ/h27yMPC4cl5Q+XtlA0Uq4X81jDpfwaagjjt
DWQ0dq5QMXLHB7JBn2ijvd1RY8nqlkK53mF+stHBzsvEppWov8iubGgmgwY2q2L1
qbgDv9jKqk2eEymlrOdJIUJZOzIzxwNNETpvUQTM5ZTTOwWboE0rO5kTyFA7vopc
T4RkaQQi6cbIXLbBFg2bkQD8G3LEMfkQ6GtEg/uSPsuCxZrI7llTy+LF6OBkY3v5
YO/ZxIJyWqolsQkWpy1wgKhrK1Nro4zGQc6bH11GEy2DsApSQmT5r5+BrwG1vdVQ
gBq+gRBBZf9hE2cCFYz0Wskc+14xI76rUQeRxi6op1qukNCuQlbRqIbK34bg+DCk
a2L8azYxUrtm3IqaaivThgPXe6F3OSzMNibOL24PbS1o0Edrgqw3/3V3SHSA/NUR
EC0QJSWlrQJgLi0FVgsbWBbPw92dxRzDa126Ufb2CxHqxDI748thqRWUgbQ2/IcN
zKOwveCsZItvuOGNn5jIBGsSPH6IcW13RWYnzGcxlq5K44HeZzJb0Yodn8SHluFy
zjZIp8errMwOaH8UqfecsFj3bGP6qUT7hveByQQln4aHtBXYFD5oHOLVWMY3ag1l
JwDKybnQmtSEb1brAUarNgMN99bUGGsBTSIhOV/uye3PnmjPiOfyvEm7+UlxnoDW
aERnkfBLZjOyPNS+3CR7ZP2y+kllIsMDxB2czfo5PgQu7M2XtlY3iUXxoLvcxAKR
f2DR4qp5k1O8iRauOa3JqleCSuv5t1gk18meqeRKCwej9Ee10ODUHrtnLG1X5j6n
U3MDY2sCfwcvM4TggeFXUio9suLzyt6SGhXy1R970q7+CSINfSQfNL+Wi6RHGcYW
dUyfihozftiPe++hck6KSBqO0bCkFwloeTPsU5fo7hBf5FfEWQC1hndlgcmMznVs
sCPj7+kyuksHkq+0Qg0BZMYGRGz7LR/rVEcrSeVZbaZuhCHoYI6YQbSpckyRxZco
wqXOHOS+JKDo3+PH0ttqMvOBUFgpKTzpTd9pbN0Otl8EBJViaFyiXv5y2/qjM+5N
3an46tOje/LG7lwV8Y0RvTFwVT8AK/pZ6N5uZL+lnVUsCwin+ZCBmI6/X8gj+nAB
j/VUp0b8vfqH7dNj6Km8SmGH5Ssuhy1/Gc8vwGFAYzZqfx5TH7rAsbqmHCsIWFko
56BGBYmnq3Vbkfvcpoh4d8V9cHMhqGgttKkQ7GaVwFLwkC0LNxB7eMpISXUxnTH5
WxN6LOlDv2BYF2YuE7yBLAYon9DXhns4QrbZvm7jY/6mSl/lwgNNCmtfiB8L41le
h6OkLFkE7jJTyB2Se8279Wn/HuIMjB3oTUK8F/bOlZYgUfVDtqDAkuY98KaBl/XD
OnEfYssWP0f3udddl9MCDGwAV/3t8133gb0jFedWBFYWrLUVJrKu0NMIA+kT5Bet
GDo8oGeqAMOw/rjqXJyoZc2m/nhCYt2LSshCBR3UwM3KmWp+wovqCEnr9XaoS8/6
sftWEMNOsJbONY8BVrkte+ePo+lmvdhHfmSwn4ycMggFrpYYwXQ5Z2l61Gqm+/Rs
GaC3B7kcXTgvYC/WU9V1UT1Qvr7+ao1ZN1JcVfTJd6qnJ5IVfq6pPt0o/iEhwpF+
vauoAPKIFlIlh5lCssGNzEjflimE4WXqpCmpTiF0NnW7qq60AmLPoGF0v5Y7iWsG
b8X1r429y1bLAnsmLxS0/GURjzoOCWqIdqzHWnKeO6rsvsOQW4NhZ05l6Q/eS/NT
BtLoFmNTFTobpsVkGj6KHEBOs+fx5SsDtwF4Mq1Zl68zAD3ORMSzxgWQYoT/S+cf
RFHO8+xm4ZAYj96YhqBl9nlBrCJ79dwRbeVxcELcMaEkbD3/aWpG54xOTfcY/Va4
VAY1k+3apam3xBKpEIm5mYqje8lexYwdPGbY0pZsF7fGAYPRgqCsrRKBAfIl/W+J
MtZeq0VUOqqRQD/6QfpnOP0sSEOhEKzoa/75p3MyM8eSXKkIFVGi/2QOmQRTEN20
Jq/S1OsdtEeYXmcXtCQYI8sv1LW6i4cW4vP7HzaF0G8kp2J1oZnfnHJ21lVxuuF/
RzV+gAa/GosW3k1aLdF1MB3/DwpqSJ+c276JlIT8ZzRJBFdjFdGuRRWoT8a+yoTf
ThLj2E1q5ZvKBaerjJicNQvTPrisohypyKoLakm4VMyWbc5qgItsHLeT07Cu9qB/
BkpbnPGc+dO4vfY4r5zF/IoIHnriolss5jhrLTlDGCyLEZmUaT3DAmDgO0rXM9hf
mPN+TSBoBB2JE2hFDSeO/34XfUGxDUOZQukFNgbGLLevTICeEkUniAc1yL3UuIB4
tYzspvndUtZmwkRpgrar/BDoHb7osiOHNKLA6P89a82vDQhgrH0GZXm+7q3zYYr/
MxCrnXYWsXDkKVXxE2nyvQWuSiJP+Wx6IQWP5JREdPWXluv9Fg2tkY/9/JSVB1rK
ejwDvj9OQTKhCYYHb9oWo0y4VQz5a4a1ZhsaaRqC4uB/YGQ1ccI7h2NYZ023Apae
kZcn83e5gOVUbHyxhgwz1J8QHWNxkDAvt+58A6zztFpOPuXjbL6SDPLWCCRb76AR
nvekVsbD18PNIm2yJu12E/qy7TtkUiHqXkq+km8qfndnnnRo6Y1bQtwL2DDSPxgE
36qzBxqQWpETLYPFEDcgR/yXXqpjWmAjOgy47OouBxQfHaHVM4BfO9exFKLkuASk
WAmUfMY+ZDeXE0ewvHiWHJA9ZIonhIDNiRViKdPokkLW+oTMapGyiOB7aMIfV+QU
Xo31IClL1ln2McMSt2l+OOVBCFISzovT26REy+XLYq+nUcazlFC5BnNaw3Wy6z95
YouX4zt13mhQIL4EEKgPolYELlCw673LkxqDXxYKUyX0/tmzOxrmJR4va5cWrt3C
lnMfSy4JgK9DNPJLiiHE5p20AeP68s0ZyBtyWwZBqfusMX8a2VG641tjO9OXhdFt
uwwwTdRut0j8XYQuTa85hZNV1fdVA2UdUBYW7S6z+Bw32/R0iAOXty+vJMYqcqYU
uSt1Xet//l36xnwr3uEzGYzLpV2xQ+qINpNXuPDabzOkgUGZoW7XprIaKnCWWxWj
he501aLDngUKqaFWK4QvqD6TECdSYZmQ7a9NtRBgHIvbMp/WclYjMWWgBnNE1TIX
jj2/BIAotPw9bYBckgx5VhCMGNK6QmcRc4BXJEvH0YqTUiqGt0+8LacKFIWg12Ar
7vSN+cuIkLyVfnJUJ7v3w9jXuuXyGGM1BgbTQre3HO/nx0Jl1WG/ZQOCBGbmmU67
JEbI1t9tSb1zWQl16S8h/t9Jaoif3tm4j9I2aMFeuWAgrcry5GCv5hK5S+Cqs6ei
azQ6WZOU+SKhXde851RZO7GjNmbCA3wZo5xSSvPjYyybD2dyffQCuJ5Km7Wz2gFc
IJ0vvv2T+MNDvonJjviyX9UzASPIKdVs8E3VSkxBKTDHIILqNpCRH/ObfAfufVUp
Hpxs0geeACGcb7njQH2zg5KhKK+TS4jcX6L/LpfDT4UMnnYJXWgxCPDLZxICLUz3
Z6Zg6fGCSFY4RUv7kPNxx9WufN00qxAp/iJ0+lpSRoAVUf0fUppFQB5RL08BakS+
NhTsHAjSm0kXgujSJGUof4ymN7iNwS3Oo/jcI2Z7yKFClfaRJWkaUSOgS63nbHOi
1ehAKU6A9iU0ItWXgab+F6kgOE/MMrbHTpN9oVhq1Y90YkqQyZO3lCLfQxixP05F
Vmo1uNF+YGkw+n8QP+8pCLib02/3zSd9uiC6WwYE6xyS2f5MNC24uwD8R6SntmXv
M6kU1O/BtsDZ0bnd9ZscjdeHgG+7XQnrPfKiONx3HT7lPbeFx6xptxjmsTwyAtPo
hl5IV4qByVySs4ZW618LmuvTTKWVe4DpXubFuNnSmsAOmu1JJNrlR2GMTzMFdS9u
S99XPYLgKKvpA9c7oBLpNhJrwbpNH5s1xslh0RSlovAeTO9eJvhnJUjDK4hOfZPq
tV9xNapu2fnsXMCUhw7J/a1RY12RSCO3RnCO5Lok65skGYmY0ECd3uVqZadC9d4c
gYOkFmLaS3g7UsEpj71lTj0VlQPuU2LtP384D2KbbTsty7VL1V7onMBdeNfC6np2
Z+xN7aBXIpyb856W+0ZGOPbCeFcg6+FpvI6UFPToX91QhH5Ush0A+EgWB1icnD7t
Q5wX62e6Vht95f8Fu8fvAxxetOVsTdwYkTfNIMO1WYE75FP06YBPVVnxuYmX0VFr
IBeqlpvLjrYtH5WllHO6BhygbLrLXcwusA2bkkKjKAoBV0TE5qWh5ikSroHCYJpr
8OjhujP/Lz6AeyY30OoyBvPtYncawvrKOaZ9oIR3zhom6k99aNx/xWl3INbItU61
VqWMy3NtocQKm/7sg/5y20ftcukmwt0Da2vmtpPLgYqJNgPBkKnXNjqJpNcYN5eU
E/uxeD4zVaynbxSjDSprdxbbMtTUzNsPPaq1TLzXSssgf2uO7aFZFiyt82k1kGNd
5cEX1NcoktjymjSr+bE5/PVpfs2frOSj01XI/hyRmkOIBrMg6A1UtWBHsME/UkXR
NT6dIXdlg9ygdlNR+xiz6ZCBnqMZsa6cslKuYw61Aj1wxFa64nYqAYK4rLV9G1DH
Xd30Ztul877tjLq78UEfC1os+Ya6BAaOzfYPlndjtPPH1cgLcDE/VPTNWazjETHs
x47aQvUBaWb1XymLR83lQeesvZpZ1l9Q1oh48VmXWvYuhA6IKL+Wifs8b+lbBAlY
fO2o2Nx1Up2Ho8wzC4XPCDDd96KzKt3I7Qj4IJK+g2+wtbAvTwRcEUkzQ6zPs9fG
6NIVb5xntRz87lwmsTmtZxrIeFJns95EW358gis8mN3h3sxL6ksfSkrAGfjOz/lJ
sFmQWSLUXOYhPCfGE5YV3VkXAutZiKrQXbn4BdEF133PuMjfg/sUzkRwzrmiZl0f
6XBG982cjQhXO23A3xh62R/cgkOXLAyrobQ9O86kvsfcmZvvB7kuxQtfNCUhVtmQ
lyMbwpJNy1A2eO1QeRjCajQNgknIfbxHP2B+/FB+kwYfj98CQP2xAfizJCzbC21C
CRIOhf/TxxROKhnTCs54K8mUyuM/s2AjvWp8LpCFocokuXMHyysX1x7qWcSh55fC
BsFvUUJGE3RpaOJbcUKvAHEbow9Tl9Kii7T44A5ZLrDDlPs3+pb29LOTFvCHDKgd
9sz1hA+Npoj5aksXoyTSzEvcZVbMBqkPEmC6xd4VHOgZuwXMv/x0YtAtB2dgvxM4
rod7YBbdjzvjw1Bg8fUB9me4FiutLNazNeJfKwxBKtChl5d6kzsmP4wVOe1eM6PK
RCNDcAcep/rHF9b2Cpvl5C/NKF6CLM3b2eZ+JncDOluiX9ZPhJRO4K2tUBJiyoaQ
Xf3yz+Z5SA8qbR8bDB0Jkcl9XRkySnM16KBxS1YJ0k+LLrCmpOCOxKvgmTngHP6P
meODw/8TBUEnpHt8/5d3Q8snRCcbVDX0Y4v/f/qZhnJcv2zNQlOyYyDsOSo3rXJs
hb5H6fx8wt89Vu2VjqU453Cv/ymwkaZn2U7Knj33KT8geNr9fVyYH8QJEl5LKcRL
9nv7KSlONjwxOHFhqNb0dJ3s4xCFnLbxiX0g8fd6/1ocs5kN/mkppX5oS5VXnYI0
NeskqPGtMFD3gMLiUZjXvx8IfbkDmxfzCsOa/8f5K+r6dSIhHdRe/JH9LpMCjlLv
SrlF5YXplgXvdCjM8RKxgTGKTbKoJ744S5ccxQAzI2RedXNZxLWEBZs55tpSZTOP
S1GsBfvebmR45BkOO0t9Nlv8gQoVBKS/x3+OP23CiKBjHe3F0UqNlgrNSNbzoLZQ
li0rswM9wSKmeFF2wDKtoa4IfhzOUhUHKyVVjdPIWElW1Q7zeXIW2celNji7Z4+u
FIUdFFhBVNEBJS/eoOqLhLtD+C8Gvtcinpw2l1/EoAs7E+4XBrDlrZx/okjlTs0j
ZhY25VyMe6TNB5WBF92PP93Gc6LtZajsXZ42C9Qq0jzXmq+k/9MpnySSd/JzT7qm
Zt/G6/Bx2a5H8wAet5wSBabcJtBzEn+lEvqAsh0aWCtFuwMLuyIXEge26iOjQaPM
qXx94wvDEulR+3b4SbruF/XKJF44VsLPu8qtNzi4JI6lCFuDr2HqK4cbXZsm0fwt
+wnPcZFb/6bjXR6Ucv4u+xxqA1iJUXxSh1F/icj050/mVMRxZeVCcgL2A5RzPyhh
70vspFnN3mdy08dKSMKEK+alVEnvPq1jNuYRGxiEarzu/rPtB5NP1NVddUEjivy/
Nt4Z3zYTITqJilI3lvE/U5wktEIbhSudA9BLrOTvLmL5FnDYqMpbMIBVcZiMgIvH
h/ouOJcDG8GpgoqoK8aNxiXVJFsANNPhu1MEtf3AXg3eSZaAzvCKtqAvLARPVnD3
D2b+Cje5oIted4hfDn0Pbx8CeQpPN4cSCd00rZrD/4+Tf+LzF8Y3QpVUKoinyT73
cs0vme/XuagOEWHrUBApEX0io9/ddnnBmne6BOMvxU+oQfpa3B5UcwAS7i0VwCKw
vbMNZCR8Msgl9N9EaKlBv0K5vPrjNCE661IMD9JIhhcqBWWb22fK4FA34G0nyGTU
fKtUSsCK+31eKuRPlFv91D/6TFOTmtk8oTlV4bKmbEl6Gk1Pl/vAe2CxzI1BbjpF
T8XbHiWZjnTqKTAVA4pK08dfXWAGlFDS8CaazLzskU73G4UCgtZtGiULdYdL49Oq
51aRACuUSjxWXaXF9L8x8p6B6eC71Mz2BTdR37KgNNsAw+vzj0XthsrxgCNHxaiZ
+sZvjv7x0IBGxbXxIMGh2jkWcasgxnTHmYAdQW9dVzgxtvX/q//vrPODN+bPfkvR
gzT4Q40eWzXl9u43PrS4SMpfbAYGT0Z11TMGDvFGXdaEtJvoWOTtaxMyUDL6U2As
YxzKkPe3onjFze+AHEs6PjOMVo3gt5xStfFsMZrRMb57e4hO8JEmt5L/8ra6f46J
40O8WIqpn5sXpFKmnxdyD9RHBdurYa7c+Bue77yhfXIUTC2QuJbIc0VpgGHfWiK4
9dFnkjh7HbZEeJ07tb3zUBMU0l/dDhlMQhoiic4BHGn7ldKPLEATccvKYjLoOUSd
HeGzwM31vxlMd3AR7vnQg2uo9V2P2gCp4hheT0eCoijh4kOTIgNEpGvRL+c399e8
inf01hyz2JHB0uP5IWRqWHTOKqCbOD3NF52ViCwDzhO0kptb+KmkcVR7bOe6xyJZ
LWC2vtW8J8+h2gzRQ/BtqhVu9oAvm0lELDUeBY4F6ojSGe23hobQnFZoZX4vbq9f
FXW5UMAvqSFucyrwfP/FGOAu6zdImolWtdxb7q5EPPrMaqLiJukxELz1bYoZX+oE
ue5shX3BKjoTGe5CYkKuiRswPRwiK/ebBm9Rfu9Auft2gDX/ME6oNndT3STScesy
v3uuSe+pILAseYlkcS/QANJZntZfdqYQa/Gbc1jeY+QWYodJV0IkTsmwTJh5ixfv
hddUE9L7J0oZKDOjcRPDKzAa5D0i99MVlOTy+u+wtXKTiIJrGataEjaPYb8xXfDG
DVLvOu/ciQnj8tSPjSzC32PyLRt6bywrh7OSyiXhhGe60DJF/R9nQfThWinqFbm4
94ideDzYdcKhRVgdkMDGAjYs71VuzFWEdvpyeuOSV7S4OaTO9tBEL45mSpL711U3
AtliXHu4mDgALISz4ynstMiokL0cLVAhmzbZT8sOHGzJoY18+NI3gWRbS4dCGGva
Yt5hEqHRa7J6peycTcVP8dewepyWJiTxDTUW0vujZwOaZWVdqRUIJ7n9ClUKuJf9
8TF4h38E8acyzmcLrMsLrAufzny2IL9Lx8fH6Zl022VwlmRlo9gUElCKi/PA1STX
MkMFY1YSHckuFFvQlSxPfW3DKQSQFovTbmTTtPTIL5TJc/rxtnavTR+RGgbkJ4h+
w3mF5xRtozDxwFdXrwaWjgZQPK8rkC82wRzinX9m3jfkntDHLEIQdKlsrS4RTOii
AZ34Wwilvol4Zr7A3kQs2cctON3Z/7Xf0kDsrOb+oR89Q1nUcF33UXlTPuygAJz2
FONdkWuL1ilZ3t2n66iqCXKRFa7iUkdcpxg5/3csBz5mPqNnW315VzsAttegwShy
SOT92KpoGBC++ovFnXrqywyQkNVbKY6ca2l3AjxZqby/BT7UTBknTN64MlgU96XG
gTm0mAHgj5SB7R7Oqp5oofQ/61Aav8y5bGpdV8IOy5KYsfWNdNOoWhDIByJCN9TR
jNHsi80PZZx9ItxYAUbUbBXmBaA1CESHxkFZT2LDGMMvONGykZO+wO/vQGDecmZq
xddYiIKRRJb4u+dMC4YaRoz76KySQB/6iKLfsnvwd7GqRP+p6V0/qGukt7ut3SVt
6VFfTXpDPTW351C77g4pj/sPN31DpcStbrRtfIY1hHe1oZJ/TyIKasDLejA9azk4
GQObUOC4TWjIpedYkiR3NA8rp6zXkr5kgeP4kHSprBdlEZiU2dwRUnz7TXpgb2+e
RZxCgeVvwelyKLvb+lteIEUlAkJgZkmyGjLFaStYJhpat2u3tk/IH9ne0+z8mLVh
U4Q0gkg1Wq6r5v6NVt51zsB8gh/GdPVeKaOYX33sJuTbSkRSfycnafRFShI1QYON
U+emITIeBdtIzUGQrlSvv9zKJ6NO1Kvs1FwJl44eNXZTfddHIUzyVBdNGdDuNVeI
sjl+ydPcarkeJAP1fstiv2m1lw12eQwmMybUPgVYoetPRhLGfj1TLQCga9XW3iRa
1yaBCZ2UDg7ZLvS3vTAtMb9L+R5UytAjAO+TAuvI3I3VnX5PNo5INQKeHviS9a3y
WL5w029AMJaCJZnyATku+H4nh7A8l56qyXlqN4EQb/A36rV/8wEydQ43YHeZHrId
xNwpbVC9QDE/aUZKBhXRHcta+Vze/whlsCxFOyhP51Qb3783ZWXRZRZyD88iqtcJ
TeqjbP1kZbRN67dIoGeClaZoVK97tWcqf3Y+cV1GR+WuwsDCtVuKvuYKhU8B0L/n
F9/NOxnMNWw+nJHirdsefi96+fCX1vOT5Km54HSCYhvikJj7Vx6LXOmjvMfev7wm
BgJNbrmQI0DFSjd9dQup3aRotDILKh/nH20uNUs2MaRDGYvfHc5YBQllKd1k5hoI
rJqhweJltJWYoG5FGbSSLfbfRxRcPaW6R1UJ2r1mT0omkHiU7DNMdNNGTttqA9ZG
u5dNEQ3c6eJzird2LO16ouGWQCsO5YkzYOF6b0PXu+PrlOrhRLbP5m9xMA3qnv4W
LyF/x8WpWlfifqsOQrV/oJWqGN3tg36/9M+9/bN/CX24GAiNfGzKXeRtITvqMv9+
i/JlUzh4wL9xKmsWSammqvbmR+uk05FKQBhZEWHdDSToe+QpZWQ0g2Gh7DzBmji0
04ertVdtRnHdnLLu7ApP/rkEdBJNb5yqyW9euODdz4+w3lLxcXv3bqGpyhWuP/r7
YlftbSTQnWbrTmOoLxRbNGRvqV5BjCFo5tDEVAeWNTdhWbDTyakOuiMEW6my/u8B
NZrD1HErzzPWn9SsnBUXpGjUTbkHMiyFwvage2pkWmO04So4WRqPGhv89Wy5i8Q8
7OxLRAMoLlGv2my1A1Wk/sWKfXc0k75LugkyiYRutzSY+NzxMzt9r/uB3VMnAOTQ
1bA7DOpssuLNgZ4nXfiwKFpQC9K711/YEgmtDf6yA2PzvvSV0b1OE/Gk14ygpfgR
Ci/tBe02O+hA5E38E92FJKPfH5geXohQbriVYzyJEb9682inOjP9CauWhrDFgi35
W3Y26DOJz9c4qvn3/M4f4yjHwRDDH/8Li7JclzIUxk/LWgRan5pyMKg2FegnDdSD
o4grr/G3bfC6LR5CziFP7Cx9Hdzzj9OIATdxQAmyZhFhgVS2V+UwHbMsZDnctMiy
QMOWscnO3itFcegtg6Wpie29200c70qAtDcNWRWzP21Bmr7mkPHXGK+mar1GVxRS
OMN9iw0VXSa3rQVPUPOLtEGlr2YUCt0ROwG8+K5e5gToeTjMlQf2d1EwbF8uoA77
jWnNXJNDO8ATIbwm6r065EWPGHRe5F2ANvE7+6nyC2cv4HUOsYg37xO/JZkzIcLa
UcWBGgVtr3yVxEV9e4xlgQwUzoW8s95TsUecZ3jSJP3hBqr0bFz0QLedXhC11YWL
`protect end_protected