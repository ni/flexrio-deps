`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10128 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
akBpHK9XojjdOyFTP3pOwlnrEYb4p1f4MxzHqe2QQTtBX16HzmuscfeOI56veF7n
C5b2iTKFP5rXPafmWjoFzmeR3Wvjx6Ha/QBBB6X1sc/VKfz6fyQrgFXL4qdrw6GF
kJol5LiA5dp/DSLVkDN/xkTVqEqv01o84ZSwpU9m+jOp45bBJm1ZGzX1imU9b0py
cACCsofODO2Qr76cfeEwtDB+KkkF/xnxjY4hQRxA6QIWaWRULDAHe2Vc/KzZ42e5
qhkSpiApFt9w4FqKjBBtzxEaOrMks5vwJNYj1oZwzK7N11gZUeLZp02OVXUMilhp
SRAspjvtan9uxkOsVEEE6/n/yoXFxSibrBpzE2v6jXn7Wy1Nd6uHmO619Ux+i8y0
pBmByM6girpxFSrtsoDFAWiJ6++wuuL/aA8vTwHQPv2ifDP0WCU6oE7Wcz4ohOA/
WOg+DjRa/0s1fa01c3zBYYhIKbQU7DyYE1gVNZQ8s2jn2onRDs2HQiXwrZPhKX5l
dPx/wLl56mNmwZKDZ1VRopZIxxLfx8sn0Z7cgJjP81Lfeyfbffl88futTb/bgIsQ
lhim2TMWKlLfegF8ugZOzgwF4oR/pup64K3EomA3Dx4mZx0Lee18nVqqU6ugaABg
lwY8QdlBFFSjMc+tcFAvdFLIgyHrI02sUD8rKoLjzGPxmThpU0iVOr3J39IH3zmK
h+BUUjnF+uGokFGdeAhB1772H030db8indVaSX8z/kaEU9+F5+yP3Cbo3tHc4x99
kFm6TeLApr0fC9ZuBw7aa7wpiHtYXGv9o/lRIaTqt6xzV3axBlDKBh8UXEtNulHH
KCNBxsTgFJyL6Ih5CY+YjKulCfa9lPNJoYpJEai20PJ8wFuwiMgUb+//vqPPZqKj
3USi6lR9XCFu7qD2RGxhGftP8WEN5HGdRoIpZY9jbYzp6N8YWJ+BRI6yqu5VFWUI
dcC6ljiRlnkMfkjeaQWiAG9I2wZWkV6NqxaLwzGXFKSNsZYBzo1xrWm/k5ReKIYK
f5hQxdiLZEOTlvz3VaEC7bQu5sy4DMigg2nfQ+JaoMkUgrjJ6EuFkwn3Z88r1hKu
Jk9dREjuBfbiFaIDkplyYUM9jXRZG8kH2yzdJGtAr/ktA++x9X458A/Q4Nu8YREo
HBnl7rrUfZXho0iT2Yy3oF/5XhzmEBrgmlzdGOA3bxsPvtEiw/+ZazeL/OziEoYM
t3FviG7A+Vk8vNvrQ3+CW7nP07EExtPUbmKGX9vmOcSgjQvBaxcDqLIzEVqVxUHo
OGvgjhnNrGNZyDoWqORN3yPwk5ShYpYfI7TaapEc7b0U/V/q1hogUjTJeGnF/WTi
B085chmIqxXol3Js307vjpAVzUVS1fUkGSsEszWsJDLdu4xVMZUz5Tdw7ZTxbxIi
KKwS74brePu0Cnf5wmrh8ecdtdYRQADl729RthesthT4raT2KyAdgZcAWGmF6WFp
phiGKyCBzt/fVKdQZwsuCcQhROuDq8rhOxjUieYTvNBs7phocFME2k5ni+KdUZ1t
NUwBFuMD4kZIjT6VY/KflDwODGt4EXbNetn/rcL+vFYMVSSGEzBkfqW7bXIFkRUR
79kb9qXLha8Z6tT0WxIQVXC/CvAatn9eqe6/vmLjMrpo8sTFvbisLNWVTIsUfSj0
IwJs0VdzvvsKT1S4XGAe1BljYSQopLbiwmLNcMZ5ImkgAT28AG333Z6zdIu9aSJB
8vn1hVkDZmr7ZU0R7NGRxJJXXNaRcPQMjHTjL374t5DANPQnzh1iElAmGlFZeUoK
5f1RJGbVfGaJw3VKZuquU7Gn9neIKusIQCWY21veAcLH5Bh+WHV1LGE2j/VyJeOU
inG4OK/yaZ74Dt0xJGocr4nnZxzqj5FM8m+qGK7nlSeIj7OfrN2UT6YmK4/jjCXq
yiuMMHAb7ApXX8iY4iZFDj0Ac9tVBcTq24PSe1ub6H9VTCCHnVaaKgDkUMNxV5xJ
uKjUJbfQvS1HtW4xUPXTzmLwbxN7Navk3vt+rI6HqFMMyy/gQQWpcp8nOoWrEqlD
Bx0KZ7EgMGe1g2LTEs59UUuC8YjKGZ1HZPEuR+fqNpPtS8kSbquUcyIWhGe2hxKg
C78JjfhgZ8O4gvXOHMnkjjIJgIA+IOLbeSQWBpN7Co/0ixd6KJ9mDTygMLXDDXEf
4vfPf5upBm1sBtTK6ZmGPUv1fWYME2ZLwXIrQusRj3u8a9mIH/UBr+oPMlgbA9W1
sUxHg1PpsR3JoGdt4VJfU48if8XXRr2LnMLBKo1POhABBsSEmucnpsVS7mmjRqc+
qWmxMfFr7ad542xCZ8TYDbSFe247I8MqshGYOzHvwEu/QIu+820PG53G6/+W2nF9
Egw0KgDEEZZjarwJkXuFKTUdKrH5QysbhPxbD9037mESNw8YYcO6W1UxqsezCUtp
7XESOFr8oUQgMX/PuM92fOVp/kYb+E8aKI3r/g1Dv+06cBxM3gkYS0gyekyshflV
H4q/k6o8AQDCli7kPkumjfsePL89RlaiAOvzhmqRRxN/d/lBC5VPLw6FLDUEOSYt
CUv0b2c6P/RmlzbgWg7VtGtPj7TPBeZpKKIrZ/wr1aD6xgfx7dwtZwzuOZhvj+k8
FhjuF5DDsgWMrJ9g+8NVqDO+9yIW7+WBlt2SobVbg9klHZuSqtTh2spWIfODYjf3
3SMMBofnmkeW2d7bCBq98Ch+XWsHMu2gtEuJZLTKCVDTMlUOKaOa6uFD+7KA4oeY
2u/fvpfrGQrhDHsPti/9hQO+kN+FbJlloTbEU37Lh/BynYcAMk5U/AJH+Y04pIu5
Am2y23cF8NulbsP7Ad51mzVLiwBaddeIsFYy3DJNt4bqLt+vMDAb4q++u1sZyfhJ
7CHWVsXEkOs2wb4aAL1Bm4WtD7Wep4Axok4+uJAG5ELWneDXaoUld6vytfa734Wg
CPMtz+h45REl7IU7f+B4IxQIlDeAeUPLfc95JYbN8MvcZikDCJBWQOl84QeE6UPX
RkeRAR/rNTzKQKjZ84VEEVzNs+6Huut1dnFcXizqPp+ejPlTF5pD5XHjA5mSOEWW
KHn9n+P3p+/fjW7Qqzx2Sg1w/7CNnfGSJjcEM9+53D8l4isbX9RmuK18vQQVGIQV
zXwXGjQLQTTZHp28hRdsqHRMklEigUxA4x9Qtg5z2EVAzZ/9pN96S4x2eGLegd/f
ZqjSigXR6QugXSi5gXATSzSj2EiVcZyi6YrQyXMAHJ6UrAqFh8N7ZydX6WNzj8Cr
T06gwSgCXRMUe8+DZS5CXC3y9H2+ByxHQ+mMbaiiC9Wt2a8g3ImhJJFbNBdmDiF5
VWKqMQS5cM932KFvzDv5SMEF9O8TeUi43i/L3Z+EcG9d6F3Ge1+ThSo7S7lxdmGu
UexMjgfKybgVGn0Hi70mdQwDOj50ePeeAuTgtz7DuWiAy5YWyqKWfN9oEzbOvpb0
vU4mknMWRTh93DZdpo1EkoLxM9WXeMWrV6IXscq5UW1/b46wpO1ZMCoZb8V/0VjU
QYJCp31bx9O4pnGh4Lz51Zvq9wv77Io3P4SoVsHOa9RfWHzNL8JvuwzWApayjWty
8rIlnyuHOw9t3XTLIbLJ5ZyU3RoaSB0oCZtL7wbfRQz7PFBCJdl2qyZke+0fEhbA
z6vYQjBkt1p9+pwp/6DR5cC+aYqn2dYN2uwdPuELQGwpx/bUtMntIlhp6L3O7Qn8
TU36RKZcb26fhspF3pEFAcUxRIrs3MAzgdnIkzXWy9ACy28gddyc7WETgfF6VstY
vwWHcCHw6bFcgB3u44jRMS/QODsUqD4wVEeK6q9N4TmdJxtKEhDD5P8tqcHS/JW8
Nl7DGsPH59FLndN8h8o/wFw1zx6A2WL0NSMnh0UGDyzOxv8ZpepL9ZCuq0k6BwVx
vIk+qv/kFL8iBVxK1F3r51Pg9JH3a6JxmapAwq/YP786J3nHU+HImIKu6dcxVTwy
aZY2oZz2ApbrFOwnxL85d2O37gxIAebuUtvaxeVbiMI7cRdMAihhF0Q72jUI5/iU
hA4x3OH87R+Oi0XHoQFnds15i82GtlabeukHCiL9nAeLJT9S7HtqVXG/lmfTU6TO
JsUeatTH9ph/YiXWzrlYx5MxFLclkVsAjtowzTIVeoWVdbJR5FPcN2DHjqnm3g7e
ecklEYOwEl0LDf53eMrLVH5AEs1M97ogfwHENzmm4FKP7WUTTDSzUsh8JYFnhGRn
q/27JFx2WhIanMHKVC9P6u48Bt7FwmRmHBU3DR6O/rvn9x3FTZ2r52P9AVgi21Dq
+6JA+KZEJNRqPvZ/GVcpd/EXHYAYtGsrc0DliTRbZBdcD/AGA2p5FSntD7XE/Cqm
d+1RJsskhV84mi5pp1lNAwZz3bnfom0q75T719czsTHFVuZnBOO7cGYOw8FvqRbL
Q/26KK+X/J/hT33UQ3YzCrOY3m8PtA1SQSxKFwQntUe3yd42GpRGn25KmKDlRghY
wcpIT+sQLRr2ANyvumYPk121mwwjJK9uA6GCz/mykEpqq35mTAXro34mjfvVYnxh
wfKuOc18XKssyQC9ZLs0EMYUrVP2/Kg++J6aASHTcmh2zO5rFmITLU23F4+r6DWg
g0UWoo7E6OlmLGlYGL4saUnEuimDJiitR6763g+XEsyYOif4MyZnDfh363qwuG9k
gxhCFghxrDaLIfncYWC7D2DNs4b5+cAJnGspr1b0bX+SdPbrjTjUr9WIYavirJAt
w8krHCNYwQSOP9Uz0+EVawuuwfpeO8Oql3s6Lg3pRhaWDDvhEgr+lXe2Aebvq/fk
le5vjXWt95/h4hDIcvFFpU+7TonFXT7BwSuhpIYdFrew0QIn97HScuLZrrNihKCm
3KQQcn96e1nhPAVGXX0GBS1mp6++sKV+5iiaK7QOlIsWR48Aq87QvAthKgvxrMQb
pKjDX//KNyEV89ZYYoRcfdLdWmOIsuaNDFW2+/h9ZGpX/N07T2A5cV/z1KmZNSIq
o06uDWyxpcsRNWjErcZIsaaKjS6dyh3KSv0PKTInQOwjzxxBZ8FMy9yTvfBa0pJH
/iKyahB9PEoonVbzVIDwyN/YDaMgGI5VTu4EoAaHqznNgO1v+/WLo7343br9X1k7
RSLZJ1pqiHFAILVEihWRUyJI8vgnIEE9tZrbs3JQGHnMj7Ouyh/ISHZkrDy0mD74
dKEK3Hj7TagkhTUG+JkD/6uc6EUgT0QHpi5qm/Q2d7G+Gw8HTruwPV0iArjlZdVn
vJIBs3iQgUZLhAaqPvUs8heGbuw3h44rUN2L2tJXEtDK7x+9xStoicExuU7DEiNd
Ryafg5vqvDB4EJzqeGDTXcsUa9u2JlFOP3aF/q/02K1D5Oa+aiI2LrLo3YSqxHYQ
b/buaSMLDJaH44O5nJPg/rlfOV/OqVxqD3U0J/q3nICvUHcmoPWppkDzO2GQdmcr
FPN2O/9EtVL4SltK5gVl45/7rqxCCTdvEuEI1yyBtCiCs0mBF94dNdZwHP9gqFrN
CQ0n8OmPigoaTcnENbnEABPR9iWSFpsa8np3PVssaW5Ph7t7O1WF27ETHttqopCE
tax6kTtKMmb7VlrnK/mytGxEngUkguSE7CqeWjfEklKASyBstcOgy/5E5hjs4G9Y
BbSGwk8IAxtIaypJe1Si21UV+o0vXHJmCAGrKYGsN0DT4wLWkbGwWC256kMcskkX
eH+rbE7qfnLm6Swi+c5n+uhoOstpTAEiyU76L1m6nsmgW20s16USBjNZ8m0YK1bv
u3x8KituycY5S4nKjh3M7Kul3vIbeRnD6uAYGq+JiUVwjVLIQLKIir5w7+S+DYZJ
/GAA7d+/oHhYzcCqUI0xtvN85rWJw+eOfLlFlDqyBL6//BTa0P4BipH1Qulvbbgu
2iF9yvgwD0clOPjKWUvBZnDFIlCM5wh6isDyWOWwCbTQT23y0hVAI4e6EDWVH7vD
W2s2KiefTdsjtsV0xAYcTVaFgl76mvexNM9SbGttwGAOAx02QKS5L12BD0EWtuZY
Yen6H4qW9yh/vERT3L2G8qGs5kX5LveM54IgWfJ+/Vrj770dFILZx2s2AyLxgRNz
YcZ7cGpFmKa1L7dUYqrReuwNVI5x7Hnfo4sLiuK6cn5t7TvWTI23dnjldpwywWWs
5pWXwxyIR/Q4vZvy8kltLTWmczSDgFy1gy1ojo7VRsx4X8fpZgOC8BUu37MTTDN0
hLTQrezfkiv/O0kFqjY2MuRC+DtkbbmbOB2BrIK9WfO9kXt/yvktErXqZIraxDAq
54xSg0Rs3TERsIIiRxpKvaimLoVjhsT15tltHk+6/D+WZERSvZuu1EZ5Jd80AtjH
2baSE1z3qoocpUbT5T3WTB1A5k2XJpYY01LjKGdhJeGZYKS4XOg3RwKW4+128UsA
vLk6q37zfErfFPiezfzloQntuRt0hVE+v5NTpo5LMhL1xMFlw1TdRszxr8LWP0/o
DF+D4BS1OnqVsd4jr4kneq4eZ1VfBUWX8eZE3DUCWAjmuE+N25HPpfVulS9ACv8k
HAJXZfppqEuo7+numJeyZKnUK+/xByV5NreHKIf7m/kKI/rVaLYiV56rwe9mf0nl
lu+aPvWD8hfrYX5T2L5SGyHOcme2ChUbuRiRaJoAFCoq3CPWdzJWeV7QhFilEumG
3+0TUPLRRunzMnOQN/Yo+HEfTY4MdHnfylP8rVTQ0WNfJD9dJq3pGhdW64E/EfIS
V+NaRSUhJ+UeceeEelJcIiFBH0Spse+dyVERphR8IL0KowyDSXr29PF7bspc7zvF
DTM6Q6CbQ9lcOF92TCvAXSRCnSFXfsHnykOquOetu8N259FcwWefuAmHQ8JmMJGS
p8CB+wK5K15ngiaBIC/3WcacihdEL4/dyVEGU4ADCjP/xtlJSry1oNgjjRTe9O6f
ZyATTV6i0zJZSPM2xxkClLw4pkF7go+K/Lm+LdLUsmhkAK7MmqFkuqMwmKyMN+Ti
YZEnGMnlm2UnEPSiw05hgZ3PqE9LIpRsxgZSxXe5WW+PuFypLLgFeVY/Jr2ysAAp
RS1igtdY7FcxTe43z1wkulzLlQSr31n/j0tMTIKDZxhjyO8T5WjvULk1aflY1BR6
g22Yxy5zLjA6FaOd9yxv6G1e9ub8fZ+ZKPnp8rtohiuwHXt78Dtm1eJDoQaleeYX
pDmp1ieqDfpJy1444iIEzkvhOrLy08YbQnpjsm0U7WkE1gZxSn00mj8ftvxS1jxP
Tt+FPOJ8xcLWjiKw/qV1f8GvFc/d1vAb2CE9WH70s/UDBw5NmfCm4qjmxTfhEbJl
Lap9kGOrJeImQp8jXpoPOH+iZbhog7sApzR88YTgeLDiHWgjuM1u5HD1cvHcIOhx
XeZPpP8u3//9CCifsIw5Mt7FUAJ1RmJxb54Ec337jh/qlBSVnDXYkHhW1JXTtMoU
en5N0M8fWPxJqUkHOl2skFuIJdFHlXEq3oQmHIvU6dslD7hVYiAreMBgCPRHN2b/
H8OB3qJDId/36zacSu2A8NmSGTD+UMjKhNBt1Z7IxOowqYlTXAHfLjaupIYGxoiZ
WnLhdmofS6TSj342qfej5Vq9zkb9KOVi8x1BfJ1Ewh0UzTuJ3HlznaagjVkhsz8w
A2Pw36B/zi1tNn8fDroTrThj9wnIy8yDAtb1Xlkz4q9AJHsACrCicCdiFJKW2XY5
OIhN7K24pZBg6cen9iE4N8tGq1udqtXY5NsYi0stYdE67xr0lcmnrhn/MWLx3rNR
VtkUXIL4ccuuF9V2sL7MmcSdFi+d70qzBDjZisNydHbJpG97eruTMh9Aaqownsqd
Bizumhrkxx3RXEwWcEWWCtauAJgyBhGENxfqatst4KJlz5atj0BT9ki65ycsimvP
XTBNvtoFVNrfid/sZZK9elE6xOsOX6WIa+PT5H2qOyTAAlP/Vaclf7R+lGS84/Im
dquHrJ4vHLcfHuu3oCP1FyT4BQsVaj5SnGsl9cpEa+TWkU0wAur331GkZHWz5E9d
zV6IfYU3Q8AqVTDEgLlKkIMDuvrWAObzuhhOPrSNvvjsWQbwL31xpsByhYlp6EoR
l9DO3OKzDPa4uxRd/gZ05H2d9/jRKNWVS/LXop078xUYfKnzpC4MHxWbtf87XtI7
lwHOp8ittG7RhcXms9O5UIRlGBWPTIJh3AHfSgCCRGEB8jsn1QtrD5X77firgd2y
l2bHy252730Tmf7ZKa+aNJPO8AraKTKnEVHXzTzY2A/bIb97DTACJVnP6We/X/Zs
hYhGPgKku3msUAlh5m5fbzGrPGCfWhx7756v9+XDbJCVfaCX8H/8VsNWY10NkzF6
K5tu8CdzL66tvK3MZGC1o67uuRJlejo+NU6Yl5p6O69Njmw0KmuKGXFK32jjFubH
iMAnw/psrjcIMHbiS3eXa4XuZjfaEE/yjzHyOkDP3DqS4J6zp/Su9cjh423uIl1q
VUPfeDgQ1u2lcO3FocVxrdzWqyB8d7iJtlnt6giZIAJyWWp4ZLOKQ9EJ6a8REF87
Gl25GAjeIgms36vm+EQBFr0+lcsb2MDbnijnE6zyMDIrBEBybW46RhdZub6AvJCF
UlaBVFFzo4g2X941Y7kL4Bi19mH6UuCeHDs7tbLJ4BpDvkC11Q/Av59meAFyLgzF
Z9EN1OqleoEYTIv5VBYaYksz6RNZWrXlKduQWxkKlS6WP8xKFJ8gxXHLJ1MMskIq
GHinlxxRY3KZHbJ2zDcLsnvQS2ZzUizJJvA+kuFpnOGxcfefFVbZRZus+aVaw4Xo
RMNWitAbGWLbMrpBVKROJnbhUpxT+mPE3dSiTO0RNyM2RFrslmKl7S4qzuogNj9J
K4rp8S0X6yEhk+SY5GHl5255obqaurfu4a70DON+b1cvWI3nqjK2MKWHrEXhgvUJ
rYLN+/3tvxuUJJMW1qGrc+IIdUzizz5eiyAvWMiuFqTJwVdfM6yItq3VKgbZtulL
taklRec7mVzTtB8rFwqcSnDM7CHCjqQi61DLTHTU0KRWUaP1vEj5yYEL1+8fYBbf
y1OGG8w4evjzgO82gLO04pR6hJBIwNle8OEK7L6Sf0bVu2jdCYwhxj8Cl2Gdd/1P
gqDDqLRUSjjI1rhkzUL2O/wkGSN7hz2HBNza4ixOVoTlB7fAvEzdYM+kqkscBLLd
EsAa2j7YZZaMwRQvZ9a6yvi3EJjL45cjW1fF/dZRQpYA32zL+MEZ4eqb//YCLgPt
yznR0IL+A3BO678GgWLkD/vNcXamQgKZyrF4uLYBKz5jCUZvTzSKIbQ/7vzpTNUZ
hjU4pQTbGKWoxWwPrDZmBIM2Sn49Cs9cav+JGvulpq2a/uPxvGT6l/wGkpqdqaZG
f4HEvZc+YKukUOQO/d2coI9jdSFvZI0LBe50j0H/jtm0jP7tiVqm9VJ7UslCmzVA
sG9HFePd8n4o4gjdo0NCSXnQ3CFOM6irmT4vKBrid0tUnnQ/4wVh5QexMMUgY4jY
P1H7ZPa6AaUlQOehCe/7zrnT0sxO2CwBcTD9wTrI7pHfmXBOXcskJAnVzxauFuW8
A0s6TL0HgmFg0YJk1RRjfaZ552cEuWMTVeMx4Oz0iNt5QRBDPemfZTOU8xGnj6FP
fY3FGNLXJJdbH8WVBr5upHfL6N6CfOqAtsPuYhY4cFAtnx/C5IDlUg59PWxwLnhQ
VxR0OJySfhxDy4X+rlqpT99UOqLX5QLCe8ab0i0hmuoKfJJxFeRz36UL/ttY3byE
DrGKSBaNf9hyE/LfKH/19wWuSb4mz8OHzNFPGQ9JkCuv3l59wSVbFS6GQnRVtkVi
kl7GPl79vEv87R7sVPp6HKnVAsZu/whUyNj5AanqsIGSbHXMDFdzUomZQ8UHHM0E
+cdZzkG1CyLHVDXxsb/jvE9Hax5ipRcEtKgbj9N4rmfxATqCrg944Ds3XElugoBI
2TSUKObEO8wVFSrdpY1+b6BkhYf5qWeX02QbaurOYVmTD8woiEKN2YuijxzQDa63
K1hzMlOofBfAQYaN4o1Y0QjHRjxBoIyL5kFc52Is4etbX62mvCqAKpBzKIsX6Gde
cvvv6yHm/YkwTkR5T/1DrRhDESQQFjCPvUeyZ+0eofY74KM34bADhY+PKX8eFfi3
6bVJxTC3O16GihRbBc5kq3jODiIszo3eB8LkGJlobVGaD5TzQiN0yOK9Me+bOGzh
KrZqXamMpuuxIeiysuYIfV/FOO8qvMdcYWa2lujV3SRZsmnWauBVAUkqgfVGBWwU
ZA+2Y2kFrqSPwEGNHwvb+7qVN9nTc9KhzehPHlness1Djznl4soAIbCggdSiccT+
cyPhGmPDMdmVX3H62uKOLzLXuvLIB+h1aqYcluQxAsrinOzPxRGW6KhKun1SblH1
46O8zsNjgzHPp6vl2ZG30R9ZMi3Njd0aSv9ldXCR/ZxYum3A8goljMAI6QieIIsl
AN04/pMIhIRyN6z3jQMMRLEWmNwKElZ6Vkl6Asj87O9EHOR0Mcj2uX1/1iGjPzEd
tLkLlQWESqSx+ebCWKCakgeI3mQLYRXt6zcycrNTJPab3spoNCR2D5aSO3/LkTlW
aABIGJiWDpA/nB9iNlti41KKyhvIBICPHL836OBPpDQ1oR2q+5xeblEvthgq2ioM
3rer14y/jz7fa51bBWuAPQ/IxCDJ7PGrgOyABxyUakY0vWmbKcTzsLs10ugR1Poh
JJY2jpgzu670HgGuTqjginv4bbNiuF5w4jQbIdAA6pUt0m1ECtLo3jYOpf8subZa
FAIUfKZsRjPIu3pY3Z7c8MsxLSl1b3eSgUTu++2meAMz/UxG5Y9TSHi10tJobHE2
4VEcLJ94uPlLcEk9rg0Q1YnEXgjumlwQf6L/rY9Z3mSAK+fyTejKdYwGS3o5+paJ
Ppj6ugnX3K8wEwoti4wXcKpsk80jyA8+UgtzZ5dzPdsJYSzcviKhHkgZ9BXCcyrU
jpFE6q5M5joBnkinCC+4un5MCE2U6azjvx2MQP2giLvXhkL8w7sl1imdL7fDyB4U
99Fu86mBzxvrJOTqTN9rcij//Lp5HCC8whYGw8Tbtm5dev4CcKB3GT56Ym2Hg2oy
dx5h30Jj4UvlJbvXKRWD2Jbo+23YuJmVbip/Nzk4KbUq8AvR5fmH3fMdgMb+tgC5
RLmseyKU3SjmJliOuL0prdQ+Mv2pJaR3/TbnZJ3H6gSlQhr6ifgFm2XGIXf+gpSC
HNHeayt3bfrkMv2QbpKEPoBk8xQtGVoCoNGyS6s3Xhftni8fQ/kN/EH4wrYcU2i9
ayzT45lODf/x0/J5xZA1jiBWB0fXfQV5ke9couRV15tslcIKDIq9NgwfoGn88sWx
5weIFLgP29xUn5b6n+YU72DLmfZ0qixbEnHcTc2k9oyAaxJ9AShmPCqx2a0KANpz
hqOPAgaxLUZBIzSubJROnlYVJToiBhwJvOc6xsw1bFksa8oZcUxG/qadxDGpbq5H
FIRSBHcosb+Ax6b68j3CV1PJWagsAeZ/NCLE83WUw7g1XwO23H29tut9l4e9uTuR
b5kGBuFmQudePOgJ1pTAd4hva7is/fMqk1I+o4yPYv1XZlcZWCjzeTupe7dnnGkU
MilbQnZZmJBI8Pu066Bp49qqfw4U0zzBdughfalHy0y2xls7XFgefmI4G7KjLXId
Nh8dInM1xIMd4Rer0dz4VtUFjmxP6fcsqpPnTF1hjHU2xXuKPjFkdXOYGx7jGvXm
R//5Supw0PvA/ft6PQIyLWXYSeL7Jht/1hZIB7bWLP4YstcL6+YRD4aSb63iez/r
ZboCRqgeEF7smxmpA9s6/UU/IRFjeDY+/ch0AbyiHpOdMNGmosa2sYDXiqBo+poa
LTHHWQxiixNgwCH51+Szf2kYZP79nwZ1DQOXEOixyyMbtKXbvKRfOZ72EKD465FH
qGPEceYxGxX07TEXgm8YeId2PAIOaEGmFA23MplxPhZCad3ORFoDlA7tHATy1IqJ
fsPrdrtvpUwBeLHlCWluwYIFIZBc/RkeL/Oaus+C9I/pfVTCIgNvOMvkPp1DbJHu
zfmELhJyeEUNAXpGUmu03BttDGbzltksgdFBTYEccZyaI2kVUYkMVaBRoNh7Voj3
StIl2ner5rP5rd/8278cpC79CuQigRFUpHKRenOaaZmyQQWUa0IGKq5obBydtq9a
cGjnxBFMhUaXPQzjzTp54lcMXP7pufpEnkTLlraHt9HoOKd8ZmhoMoO9ibiD3weq
oKiWoloXceTffcuJF2vP1GeuKSEYx/oqJK41eCHstRz5EyGj7dzv69yljimm+VRU
tpc690Dqtv/M6iAbgz+QtBVq/5XKOjkHpIMFGCKTb6x2tuUP/xioroKgcNON7fBy
EoplhMfXlEVStC+R+8egBkecqwwp6KvdHSOjRxo24fb86aSFsv27ots8y/7YfO7k
6QEUQfhOePATuT8oI7PkOwPw2bJ9JxKDWBf/i5ECKAlPlKGXrDG3HqBHBGpyWFzV
Y/JbLAHiaF0UFeB3LPeVhNFiO4hL+yXX/uZcp7RVkBO/eaX05npB4FrlA/yUf4RY
+e71eEDhCwmn0VNHWY/sLXu8koXCGfx2u8Dx1GTOzJ0iqgUlBF+L/Y2xMbYAN+9q
RXhdEi1K41WjSV+2HazmprzFYdul06CUXAOurzVmYYXwxy4HKGIxd21AhLGgVdCW
w4vo6gFOwxqKoSPkQVJjHtg2VhAiEC/xUIdCgJ6qLF6uEd1go//F4vkhScrHS9Ij
wzUBEo3F74LpgALnfTFN1j947kSQMUi0zZma5ewpjnIQN8shDx78ujINIFqQVjTT
93w/eC5yKU/H0DzWlP4cK2W/2WIu0BtixBP32fXI9b5SZlyXMhp/lAxAYpEza2sr
fxWNCpfilatvXB7KBfeQYG7B1z7b16bx+HsszbpHWofctEGqhlToONmdv1yGX1zA
xvWLJ1EMJ8M9aw+0kgOHEQZyXZj4eMeo/1TP1psQO06P+xmAIr7z9G3DiRDP1bLt
jy9k43S970K2jaPKnK3kThOZGUuJrsI/OO+egQngJqrdi9FX7gRgUP9byiQ4dcDt
P9q8DusYcpv8WGsxpPqYSAgNzS3MkT6h0yuNxbgSbVI4AomnpTjuOJ9TNRwpLuAb
S4HPPaY3/LSRthIJCrGhajzK6xKq3j7KB6UtaAe+NY6+sbmLWdfmHzE3/zjIBX2d
sItbkw/Mx/unuGFbg1xyClTThVS4YTEM1kMVn3q/udv3YJ6UB2cfDgr3LsyxEp/U
OJ3jJKTKSuTDokSt0u0Slk/RCNqSVBWg0bb+Zq0KLEFAdZsFfXucks2O10MG101s
/aHwQ/MHAt6JBmcf9GJkqNARqtLN8mCdc+HQwBRjS6YM8SC1HDizsfZfJlUXdR2F
`protect end_protected