`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6912 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
cnmYCVpqoAjvPlHjUQ7k1SvzGrKQPSUIJuD3zQatZs9DoV6xY+crtB1yO0FrEqTl
1LPrjlftHrz8uVSeKcP7+M4232aqa2UyGggRxZkzWQ7tEKWZ6IsN2RAtylSZLtqc
Bp4dQuRBjFcTCJhnq9YQfeAWD+L9GgvrJ56mI8k02adx5iM55DM3Q2eQgZ19eGqr
OW3KKPV+VNDWCbJ9c95GhKinWJ3KjBLfLxC3WNnCLtIVP1aWVhkiedrF82kA9g8z
LUcipMvlpqCQhl3tIzpb9tzSFW2+rRp4Y7XkOx16V/PGBWec+xSX5nyzdbg3Hp2t
5G0riyTkp71/D/sL9/oBaSXHXIQrdB40GISlHeirbqTNRwtNpo5EVS3kKq2eIlpx
4VoUG6TsY+K4NvVK4rZn0PiOXPRMT4+nulApz5WHow9vqqUnHYb+svFXerG9rXSk
tJoNchwY0tY5x5eP5N48S0ZqhWbexCfkuO5otR/AOcW/AJBiyTc/t0DOKKpDoFU8
tyxV83+oFAdXIWK/gp5l3/gyYblL5SlCHCUVexg0SPAxyKxXpADSfX9E+ANhRzhR
yejdJE5Z72h4eXyt5ekIsyRYx30Q7z9ffYprSsmSoD3+ybobsffImAbj530PaCcC
dJEWQhgae6Ij/h1EKaGnAp6INMb44fJpDriY9cusBmgOxtUyOc4SOKxMkbKC7G/i
av1xePU/HAa/262h1KshYDoZijJbdVV7PmzBpGncCNoxwA0Dm13sUUW3sa6Jxklw
ralq+Oh2aXmbVIaydhZ+SglpqKmjIVrjk1MDmRupRBwTu79RhjcZ1lSEdV4oWDGd
Gt9v7NmRrewqClESNJpW+B2KHAs+VNflcKujIf1Fql4jopU/IUZU3oUBHzAeByGG
pGwLjRSN+4420G2wnRS8NA/Lrs0NV5D9mqHDdQDRyOijJT8T2ppGjYC4yrlbaCTk
vBxnF5d3IupxHpzfbx0GMxvqD17bOkfrkA7I4OpQn0CTZLk4KzDIJLLnosvCJExU
n6081a47n6qR8/oCqK2qZCkenHwi3B4wryRr2QaeNLGWNyIK5DY5bIxYirPMAIVv
Cj288G6O7mx3HJ6m/ZjDdfIkudGvMgUZw/xBTURP5YyqiCG7k0hi69S5HJw2AtL/
H5qHXzGO9X/YgsqfkVC/AWwK7jJD5YvJ16mYNJ5AkQ0vzpgBbG79lSsRY94q5X75
82WWebRnHF6+tXibwNuT4oXa2/ZtsMzmV2zGPxk/n47WcKt/N6906XhG+84e66kj
BvgAebAEFfZ0liLqdJxrkMRj7zce1S8FdTcqNTHCyxiVKuxLWlyK5BFalNknBT4L
gM9hZluhIPdLUFd7SCCd3dq67/ROb7A8g8JIHjQ5rS4eZqmLnGUM6m5i1J8W58mZ
vd3kEpJc/wV5vKnKQWlbwPDaRL4FkqDopypeLa9hzgt1Bn0CIICVTT5w7v+oI66D
KNaVBW2Ckz1IOu/oP/s0CHb9kwzHOLbsUS5hI8eUMvd/CH4WyQsyptbGmf46k4fo
NUpvASWj6FGy7DaqrcKRocwBaRXMPx6/YF+1pYcjlzghACCcz+K0d5SytswYOjsO
fuI4uCt79gIbXA5aSg/NkSIQwxvI4B6JXlUH94Sbda3VIOZZtfChnFMuC/htfRHJ
cMujlD6dag4aLkU4e17FnNdoMI8piAVy28XBHsjybPIVOhcjLEbG8GfAFELFQxFK
WyYn+rnh5AM1AKZiK9JzY4pUk8dF6QJKmKnrtDwSW9k/QJ8MCdGVfF1FIc6TdGe+
WUXllzAPIZPAzMNm8CH13gWSnUpGOo/FQHOsvtUQxJGCZyJe8KTbThzLy68oXUKI
s36mjuMh96oETnQcHPrfRsf/qGJex/zYIk3Pq4SZu06b4dnQbgyRfHR4jBXP/sNw
yoeJ1l7dzkPr002Ha6JghhqoCjGsb2JzCZ7xdlFA74AgCNLlYtrQvn9KKcmbmnwT
kKYlMXODbEM5BlSfFGvRGi791ydlAcg26e+H85nQJhwA7euvJk1gmafM+hzOyiHW
1XNfBAGMVLNss7K38PQqqsRNP1k1rxYt1rbE+USRDuegr0Z1jWR0I/OdGxTpWSWB
e0TGDIRGCIcGELh9/flKP69Ul1+At1J4tgkZkyKGVCKLmlRy/qOlwCFaTvHxOfKa
QuZXZR+S5PhaucHKLXl/4mJfhOsegwzGzOdl4VoOjP82nUAUJDlSCs+I1ewMKeiQ
h0AAjcTuDzyVvQBH8eMQGKIGzOeXX4x3IzFfFfJG4I2j3Q7dsB7Rn7n3TgFNxywP
nXNiuRmwwH1Km40adhCtWNZ0y2FyYDKjwMYCwaC9ZUNt1VWB8ICXJzmDD9GRP2o6
p4Mz3+c+r2tkRiT8mkOAoR/1vcNANXMlLEF0IsStKCyTo8LRZ1rNQQbra8dYkuzi
pm5lU7tcnKZY2PLnasSQQR+g64nQ20nGgZlYFTl/7oxkUkk2SctMtcxeLZbfkhjy
xGj2RvJl3PIoVxcVUg1jrUG2zzV2i7oo3EpjzGCUdGqpAtaGlI1V77hCtbIAC63P
Gw1RMBBaCe7gTrKWlOUH9H2ENx6bB8gp0SbowGleUVVVo8jAohSEs5LzjJtujsEw
FZQNGGgW7AwX0xX2nsouDob3Ofa9Qd4I/Ah/g6AXn6ZFwbiWwuVR0G0A5ENm+6IA
/4wjbLL65/1AWyF8Vn9/QyxVIgWDXoAHnruXHIFsoHr4D1FBQfvza+UVXODjZRgS
sSE+vd1qbr+kSVnizY+fSWrQ9yUTIIU9TPTYya1xDbQMe2FfJ/40H3f0oJI3PgGY
+7110hYopLdFwg/8jxa62yqpi/RUP/tI5TsYdMtzTqlhpn76Ll6YnbjogFtbG9e2
wUO5fQJfN2KhdYu2iH9jgxKFzOh2D3ItkwpdACV3YCHpPeSst6ali28E7gVOApgR
H8k8OALPljIkOQ+Uu879uzEMkzqgDz256SSAeHoZmnsIInRKXdCQo6v9L2DQHXNf
Jg1bf2BnW4Kvataa2GvwZkwkTjz0ujxcWxGJoZ0EJGu99mFG7oNlKmlCBN2cwnQR
BLNyexAXfCCcsy6lldgEVb7itITCaxpUHLTU/+jhp9KZMVDZNZvcW5Yu3b0jgwWs
oS4svAcWOtacx7z2YCRn5xJygYvTQ6cj64VIW9fk/Ez4tPVBvUxULMVhLG21jG5F
a9iYwhNj1pCeKo9B+p+eNuHfT6+SzOADOdSJ0PTdiGVj3Yokb+t9kGoS39zLyvsC
l5wgfH0fgetbV2kBr+IFNufqGArV3VDCwm2bv/4GrWqkkYXEbwLcICwenUDQxYI+
5CoGpYAkf5HGod4mYcKc9BTFICDKPl/Lr17OVqq6c0UgeqXPl7MsvATjo6mS4A/Q
Tj7M0z8VGkDirQkzfgOL/dNhM19bueb6hO/4AFEBcLzQpz7wJYxIGHYHGUwNF1bf
W3Z+0IMYJ7NI1FxOLSWXcNToa2aM9aeGOMzGg+9bhxeVv0O4ttKELIqGmdLhIHVY
9Ho/DS0D9AbdP7aRIRqOniCnpxW0LwjofeFh4jGEAMeaDwGLS2ITz8pZziutXKCA
ERMJ8a9nwehxINoGDHJHzGIOQZpEmF1+LFVRdfcH6YFZdvTuSUqdAR1JVpZZvirY
Tkjutu3Ocf0gjPod2ZXjWLz7cwc/SvL3pccvjHqKIDqLeYa+qXnTstXwUh6exEAE
r6f15X9IDhzVw5XYqwXQT49ROHk5kHLouvSXV10U5KVz/tu0xXZoBC5dcIy/nVRX
N5I8icko4j+5nIOLvnpT3jP1PwKUcV0ySeDv3EfZvsVz9mj7vzwRlXWPCvNT1wwX
h8JomN/Fb+jx/XPk+PxteMDeuYAjv58nm9JXhnvJy/5ONdsEuFk2mFF7OMmDmhmK
Eug4AkvQzmMvLhDp9OC6HNw4lnv7L+4OqzGKzdfAgvhqCerP6TymU9NautdpVhOo
6lJWlOmOoa3hk0b72WdDOmC3D5zDlpjMQULL5E05Gzs6bVlzCGk2skIm/qNUGACw
o57RAOMpaqGtsn1vw6g6PprtXO9TDPXTpCJiNibhvtBZFxgtVW49+nFkuLVZg6yQ
G87hNZSIZ0QhIt1HXu2IGYcPDGYaoEiCtceAFDArizf1ouFykWlurepJOpHGTRU4
UxNzC5AsAvev9SB2ue/6Lrw52/Q+Su9P1qWTqqK5nWu5VzkluRFLhL5wix5/B9j6
xvKh4rfU3MdlfygnL74uL3Ldqi57iMkc5SY7bTKz4mXChO81zsJX62n2zJ0DxHaO
ohm23LaKy0ipe0gd8AfbeOCBv1N3Lqo5i9E9S+z5U5lK0mUSUxhPo6+kpub6hvTJ
jjjYN3gxO7Piz91Pt4fEvycJ18lqMjfYQiJj7Z/bQ1Jw5+HeUmLn+qd6zVLFfPGx
l1vG0jQyGyNgvLuTqrK8N0xA5Rio/8a7fWbUw2Vu2dFPe0cVPfxLTc+2GNADGKtf
qBEH0bRIrZQV9BQkgRcrE40MIfubTFEjfGwJKeErvHaF70g/R8ngIuWJbKEh2epW
eapKDov7lfy2BOwUTRXlfCMWenZdBEfnYnWXrAYais/W9TkhJoYNrFjwdSYu2M63
IJuLI5EpnoMXBVL3C7h/vvx3VrqkBSY2obyNzjRu89DpUnqYsWKnrBSYsdSvSJ4t
uyr8hBXoUILFXNfB0wttYjEvrlIcuNNJdZ22evHsFJQ/Aix1m8EChp++yDWhn/V6
oZ6ys2mTrKjh4joVhxNOC0IPZN3TCi1clvUBub8YWBpZ1nR/lx2T/mvKbcQv7YCr
H9yjDRlLDwTls57Knk7j15Okybt6uNOl5KiEGK5f78XS4fJMQGPI5O5ldJkDuOyC
/WVETV44KaOpXy/fMO4rQ8DVnHdEOtN8IJHbc0CQYK1BbmA/86sbcZGqWwrX58x7
FH/Ep69IoyU5wN7RbThZ3P3R49k4ehTOL2b1XADq7NafDAX/kQFlaeWCBGItGmlW
ShEjrnqiw3aBTDpEoQs6yOYeXCH4RaYldePuqtIb/Yv7mn6P5nndAYkXtivB8pkk
Up+C5oqDCXE1kfGMoBud8q0YWkkoudtsSbGx0SD1HaYDhaG5MzhOMu90XEOdiakQ
MZywlTk45pIEh1vL/yCG2pR07bYAB5WbvEdV9M5U+eBU6zIgJ2H8jvsZ11pAk0qf
YqGctGvFXpQNHU+UDuMuaqjutcKkd3UuG2iTGOuaa7gE1hkDjkAoidffYlqEOF2A
Ixa2f17E3V9/XboTG7DOI81UPgKpqiO4Kh+JoRG5akilcViqsIAFdpPDM/7cX3tT
Y9lJeVxHiJXlYzOsoZekE41BnN9c5JCQfjggNnqoi3qTpQO7FuKoHsablZB6bpZu
C8uoccVfIVZubkGTR5IXTj3cWLVvRVTKtlWFklSh1wOzRmHBCZaIFcwaXHlhxfTP
227suHggQcuzN9QqYxhHrQDUoWVKQX3nCVZykdF4l5BkPiqzOerCeByeIt2IkB5i
NaoPWW1KX8tMebaEyGeeqyZCtDnfsRleF1wMcoJGcP7Jlg3uzx1nklnN4tj0k6By
eyfZfcGbDgUFoTow2Koj3h/FcYskfIcUFX5So+csJjqUd8dBLIlnvylJ4hMFbGNU
wU8snm3PlP1rGazTeTvKI3Nph3WzhqPYr3rc0A6X00j3kAm0EqhIU8kb3pzcqY53
RXMIEMd8DuAzOi2kGdHlwJlm8lxqzFP0ghObW8jAsu7EB/pxq2z+Y/xwNXXkze2/
zXDZJOUcGvs9IcyNtR3BJf2hIOCvgwgv/06KrDf2sN0yLOKCfQ1eQafc+tMsuUm5
Xuj1iueQ46/Iv4hf7msASrH/UKxqltzmQBKzErwjdTXkr/EaieBkSSOQkpyflkze
FRqTzfTWQ9XnjQ/4w5u998xn59I+tsQ/MEdQDHGCxeiAKGq/xlVq/s3yOWJasF91
lDfQeH8RWw001zeo+VfM+2u4XqyT1AqpbQmdd6apqh+58x4pnjJwfAM45Cz1MWxM
EOdtNpO6QFwZ5WojlykmZVdzL5KbR9iXPelEN0FXTkE1UdOPnRRN67zieze2I8rL
wlwWZiudBLZ7BodiEZvNpOiDOPNqvj26xZ6xk25bMRy/MgOFVX8506O4F7OzTV1Z
c4wF9/HvSxhQbErg6M1z0o/N3Cnv35jFEYsIAOz9EnNLahgIffsA3v/e3dxgoNFs
tS2ZiBtfUKMa+bLfAZF3P9oNjY8JUBAFxgLy1gk2UzDKg12qdAnq4XD3ceBVw/Ay
uLUuE6LwNI5VOijbj0c5TDkYTXgOnFyeOt0mY4t4XlDHv+eHqaGQNWj57kyEIJ68
5COz6uBSNitY/BXEgwPQia9BX9dmOGOw564+A5s5KvDvS/ddbNxkyD2JYFmFvbkC
EyYPckDSYF+L0hpWBKetTCzOVTz9IfalBH7GCNIH7VV8jL+RDcVXjG+ywdNEsxps
PMhrJBcQp2q0oRWSGb6wrVl/rYGPq1T7jY+WdpibWs0JrtTUqQ/sUxEzsdZEXU9T
st0ipmL2BqTaSZYhl2ctvBO5YintITr3toRCOyIReIgX6UgnjzvSZ+XLZmoqBfMh
Of1XpdfauwvaTke8fB0nLERka0XqiNXDpsJ7WtUAAUC+pBQ6/npeouJp3TLPTnrZ
Mm0XqbUgZqCXURnqgi/m9O5k9fUEu6Jc0UgQ0NdK3cn4y7sYGyjP+vm9C33Oe4xG
VUTqNBJQfKd9nTCmwkiSG9vTwAPxrVTxBW7+BwHjGLJ35Dm3JebMGCWO+JKldwBV
8Bty/F1gMLsHydBuuIKxQUSkgVBtYJRGzurPLr0VnmT0jZ1Gvcww0o9QCDvwES+7
qne/mIArvPa8ysaqQMNGC9JpOnXdooYdTEaPPLJOlMlbPL+8mWJYHGZn4AFNI6ph
1Xc2Cj7yRKUH9qCWByMfUfUIMimtgj+k/RpJphY5znoaFGck4q3soENFM4JZXtb6
Lp/xHvjYkYVr5rCaRRARc+VJMsdcvrFrZRN5wyMMx19hHmQ5D/gJl/PiaGiRLOiE
Yu3Fk7UUtmXZj/ZVFH/lVHy7AtAgTL2q1OGcHmbJ2JRdJpEvj7xNs1KhbsFGG+ju
6WdZVnSJQGuBKO2Nr0rYVmzf5z+suujAWXxqVQ5bVkM0MXjIciR38SLVAHiSFSPF
av02yXUiUabgLTt1iqqwuMgXPTtlZ3wCeSPoQGc/ppU0FuWUFPEYjKAQMGDBAPPy
OaSPYypK5+nRTub84ONe6tDFkd0xGBbFF7BSRNC//nYgllO9DbmZLtzBSWVNNDkW
WLDGxrL3uiwsKYmzlXtO+Om1lpDfG4aOfR3w44NHc4YL1nS90eFwYrNAcJNvzbHe
ZYMgi65via2YnFnJ1wBfExSqha35/RB0AAP5w0xxVn1bu0qTNXG6dzsXrOE1OFto
9pIOcYZNCKuYSKKhYgda8fvZhTRrR72KMz/BVH/I+Ci0Uu2ZebMO4FRUBwmbpQmG
kgJD5lZ6jiwlO7lX1NxCobp48OTDAli2rWAxFHadK25Sz7LfZbMv59va5NLUzz3F
8YNFS9OPnAP2a8Ux2nFv4EMj3qLrP5YpipjBH12gXIl9Ot2ScYXPtNxGw7S6lSyj
Fd47XkCur6i+lp4ACKHa2f1Cp2uKrmq0GZS7Ul15spvYfEva7Kn4zkK+BJ3ZMXTh
nlc/z3daNjErOYXG7xMhNCrxWwhYi/Gv73N5FnsK1PHjvpfO2HKgJWo67bVCITMC
cncgNyFaePWHXT3fo23E5bAA3QkNcVqcDUQTPKtPjAXEJJrpiBihU+t0Gmp2hCxo
htZEtsOjTbbU5W8NdxYhQQ8Glv2rfelFxLp+cRwjIYwCpJI2bKBVXst54QFdjPuA
0X55LscipIyRFOVQty9+gwYkDXa/7sFhIZHbDbiU9o5iX7plYIdzQ7AwTX2B+hFR
FupZbEjq6bw1wKOc/Dg/LzLU3GGy6L85OXW8UF6YzKhnKQsaBcDxXHsUlOxzCu5P
+lfoyv0leBYQEh0yun0Hs7O5+z+ZWbb/3bbqWsUvY57d5sUxtYHZ8HVZBHYEsPL4
9+t9ka0Fr+5q9iHSInLM+B1fWSd9zAG2PYGM7kg52IeHMdVBM8xZ9G2gI5kAoHxT
IUjAaT7BxVNBFcgchYaJu/L9VcQou6tNLGMkoAH1iME8r0GEzh7xBN3XjCleapBI
AfxMRMBubxlompGLS++UROZ7G7DGyyCsyZd5nRTUJozr1JdGxcfoYtfD0p2Li7KR
bI2fhyAJkFZwKv+BdsmYixsuE2LQrtOD4QDAT4/1OYDojNkekPllXbO1gWRwqYmT
gTXc53c1bSLORtUPVof0Uyrfk8mn/VjKedYttcuodPRZtWZMtKT/cxkTMYxt+7Eo
L/aDxMhGd1pjvSNofUTHZjQECSwLDhU7duOeZAeBJafrKQDQjiDJ/vsIWTYHFZ9i
963QQZ+HCOQ1lQs8fsATLDrQwjFjKk22DOmyoddCNPwsomyb1c9805v8/P5O1weM
zGR7ukzBbqem5GvBfkAcFLi6sr016tgz0H6/L5ZUvJyRhusz9DBAh6MArqLWdA1r
Sj17w7NM7YrRayvCoEXsulGzG+kRUDlinwhLQDYAllK8iPMhlomjgngXxJGR6qtr
UWJQkw2QB5GEi/vSDiJaG/CgKXXa25ZEUVUPsEiFfdKtkPjS5v+VISll2jpX3QP0
HXm2klGeJLIfbfTYxqiFkALwLWRBxuIhpAWxtkLtVLLhRWGLjYfXzqY+z4izyvR+
mf1Ig9kX08V/oLOp2DAxCxviWUQ+WcD6X3TviOL4xubyXb22eALHLxxA8HVvKUwK
GPkEp3PKoOW7t4Yl3+3sBGwOlogPV6EQfpoPQNcQICkBsIBKUnFsWhgrsLRb8ERQ
EMzgn0PSmVRgrTq3PkZ9rXhDQXMkOAXJKingPhSuYtm0XHG9BDJJ77TfR7ShDUMa
UkQDRcbcVGnNsF2n0X1dG9yLnoWV4TGxtVh2AiWT4asO9ZDDG1LmIB5GWqwOGcfT
7rtb1fPU3DCuivVJZY6CrCuWmfiDsBZyN87g1YxQKDSNjz+o7ljDp0xDVosAVv9Y
`protect end_protected