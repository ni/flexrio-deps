`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24384 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
VKWNRQF+vfUNEEp7apOJObSd69Rk35NeQZCpjlcDdqSb0vnNGdqH//t2LGPmMZXt
YArnSgMKTMVmCZuffFKodrSkmU3hPKQyuW4uv7NGIPf7RxKlVeMyoC7VSCBKLwiZ
lmobsUekprFLfbhFuGuoLuJ7JvRu14Ge98fPxetcuSskAdd0RkvnEFYZ8tnfAIV1
kQafHAeZdrp8/vaGxJ+RA/g2pkgFf4Wm2+8MlDRFQ0nHuE/UYR2UStzhnRTKSu+D
CwKk9AEl758dEYmQ2IVEzMsCwL/t9NJT6lzJzjog2cU7J2WbjLWBKznMd4JD2BNX
l/QtFAdeQPG7IR9pzraFofxekG47xfCYno5E5WsPzk88No58maSraupefpQiPCtN
78ykNt2rI4nGSf96AlmGjdftKykf1bSOYXaCD7u7fOr8Jzv7kbwIV4KxCFwZcHBr
SnpulCriigfHploKDWWfBIt+DuCvFntjP4I45An6VwGAJWE5qUaByCc0hLjS94g1
qwKXYgh/FvQeclk6qEU6vhVK1z0WBRSKAVMvJ7dg1w85OdkIszJGctGC7aTH7koQ
EZhl0+u3jL3Ul3u0IcsU9bEAvzBQ0ZKXDqKdXgP2ylGqlegP0briCEFN5aLHbnyO
qu5ts63HTihAtAJIO2gr4WLPHeTwF2KR+RWV4ektktacMOwbX4vkq3YfszCMdpYZ
i5+2m6aP60IrvrcpXiV2ol90iI8ucQjyfJy06QH7e4N40/kQtyzHEUWDVkK8Mds4
gvmyR8IZBBCUBAHEJ7uTMblnm9A3sKYao+PWIWtf8mwUH0PWjRMouJlFNXdDzMGf
bW+jlS7RPHuHC1/TnpzVqsAT8hrwAFZ0sFycOWUUOHJajOCHKx/08MuIrjxr9uL5
3R0wfJb+mHKWTTcJkThN4a8w2Y6UkApWr89VvOjqb9bzXy5a8luRy4XecEvdS/L+
T+GgymQK3yuBfoi0bT2UbNqVFUxzOSRVO7SegDODqSEWAwspPfWOVqdtHS5M55W2
3I+7wVFfbwg1yF1gcCQwWZTi2XF6wt3Y+qin8nZMuYidKCSlJxYemzn3Cih7vuj5
Ag5JrjGVUC0m3gXm1+NUu/W0oaBXjFwAcC65AihQaw5LpUtAtUhPNQaOWNnHZTP/
2J9Stw2lRWufRQKvyx8Xih9d7rY62vqJxEXoN1R/qA1jl/Im9BamNviHQUrIQeRf
tzxMiFTH5fg12oL9WdRYupyJ3utRpvuVKIV2vMWDeYVRcX89XlvIQs4QhbzkDE/b
n/xaLjkaUkwjb/iiCCl31FYYEkId2bzv8zJAZN2pN2DY0GfchIQDTz78aBQu9/PB
D9in6diq1+r8720Zs8w7iruQyvI+i2uAd4EXYvXuWHe8qXOTnp2abD4WHP4O7T40
Z21W78StZj27N10KToZa6sXk4XL+Dm99l5/ONHsTmtqc57iZcFPG16zKWEWuXzIN
4+CIEmjY1aqU/USvLQ4Dv5TG3g4UMzd5OIUi7ls3vEgd+8SFxxIebaSdLdsTdJ5B
oNhGu9eUtXJZGfgT5Wp+GDsHg/O6Wr+8WNMdsEx3ODOxJ3wuoym/plFvdYEJ/VnI
Nn50yMgqlvL3Kh1LtoQ2p4L1N6CcX9h9ot8aCEK0B8ezLpQvqlJigZz1RkcPcCJq
QFwwnECgyrItrh1HdwsDOHN0jinBJVvTb1eqSG9LWxYD+jMZsIdxwUJlBlSdWAlT
Omp60mt0FNINDp/dNSIxbb3yIL754rpxtaUmIYGkijsO2dz7D0AVEaF8e9QHzjX/
YydsUx/eubjFAmnFyqav0dvcPHgTtK8Z4leluDWfIt9x07G4Z75Jh6KYsrPoH3uV
6uAmnRKRdVov/AlTeJy9fjy/5ldgIopwO+TffL6TxeFJw9m5EEiiHk2tnA76DO56
LQie1l4fvdWl81yJIB8xwQd1TZx2xYtOCelDiHUuD2C7Dnxd4HYsweqw28LCp1NN
lG7KHQQ/hLBkf0ApZMAEBFr1x4ZaryMqM+WSFpccKh3UIceRb52R3p8RsLHydcBO
koQPpn6UYkTrXQ09i9HbbDz8hpdDCPZYxJaplcQNF6vCbzhOE3ObA8BzLxG5VE7f
uDXR3Go2LtCDz39fMvi+86J8zM6YeI4whb1CPJq8diblko/R42C7kgmbXUq7GeJv
1M8ToVfRBLftiCWRtxOaxVkqoM5IlDnuGULKsTo9dnw/b3Wg5t/IX9/BmiwIBHnq
vZV3rOiI/peXoynnb/ReR23LGSapytiTcq6uA3M6QzQrxo35RfwbeuieFXqBRlEs
Ps6vrUvtxdbbYC+ieEXK2Zy93lUbnuanODC/qTDD3utLGWiWn6JoGK0xDN/kZR4/
y5CbHAXNFCqXNViGPTwxUeiLZCIxlmn5k5+z6CJZJ+a8xK9gu5rdbWFuOW+zM6of
vlcsMUZ/ztN1f5+GY8oUxuY8iynM1tuWx/GOhfqphj073k0/X5ysQkB1K5c+BteM
sfoRQiP28YUuegvKJ6aietOW7+lhlCUMfNSaGo+Q1FW0l7R6mei4pU8gIqwSz65+
mCSvkoT0piCSfSrsi3QlwF1qT8xEZE98WzCjtwcE9wxxOPG6bOTkE+FTko34rotr
0HBsYdfnkwOTV16OvwKewXOg3Fi7JaD6zfzZrOAKG/N0DFUlhaYzYe+JUoDzWG4L
Lvmafu1xeUa6Auv5ABOen+ETGsrOD4M/azN0YjNipwUX65BFFRgPzAO+TSKYYiDx
IGssf3PTTYMBUmMxZEIn6ydlnMZJULbqY3ZHiDER6sEYpnMSLjX15A8Jb3xEDPOP
HsDEsdWDjWEKcxBJfRcicrDWLx+Y/IfNHTbAcTG3k1ZDMlDWrUA95b3cmCRXShzz
vHIsheQy1/KEBuA/7VoybMSOvhkcZ4UHwdMzxMhbsyRpDdUNBc1hYZkHusGs2OFj
gwEyqmao2obo3O9EMfKgba4Uy5kiVCuEy7UMkN3hqKyuYPn0HkHroEU5QH7Ngt4T
0NJUIo5dBt2LazobcnFpYCVyb35qEXV8sK9Olj1BLa65g/jy3xnwiFWCO0Yv7MRz
YcMH4vQGwpj7h0oCelb48NWrxQgZUriP/UCOk1MmDOlgczKvncLhxxk74BpLJxWk
PY+i7Z3Un7Vea6+O42ZRsbEYHnxFBAzt3tDJYKyKQJMk421EJ51ASHvGtFZ9kxqm
p6l61+gY8WVX8xllXTRQ8sDknhKKDiR0Y4EwuvVfh2l3gUWAkI8OKCCTTxg76O5/
gm6oObYWQZ21Lf3D/7HVvNxI6dBknzx8YFGep3xLNaBUQgMFik9sdphu++oY0gPc
0sMd4BvyiHVppsXWb7Ce+sg/8w9WDEpq7K9oSZKH/RSQKE9A6dJANO+2FNxnijyD
eIolbyy0y4NHa0phjjiEb4+YzYYD33OGKNbeGSZ/HOXvj4oHcmft5OGX5MaPcxvM
MwvlKTq4yoCFFgHQfoLHa4egbzVL9yoEhx8SPxPexoA9YkASuiaJ9K4i6iwFmQhA
hcDa3MDKIzQjYBV+bRjW82+yPK4qxTugWS1cu9HCmb9vM7zc/xlD45VFtJmeEdz3
obJs6rNXzHRMeFUJkyxeipx3Ri2E/MCxHW+vkCLA17XGD8Yj1AaPqq4qpSeqPo9i
nJU9xbw9h9/0t8Yjwe5UInhX6foCouvjIYw5nIVlTEHY4bEnSBx8BKCkeoY4+WGy
Ua19Ckb/FIMUFDYxJ2lxx5GWLv4WCR3V4UHlEQcydV+d1S7RFSjrjsrrCSqEzneT
Kd7n9hON/F/fTsslqK+wjNXnWh+wp4wLxJRILgHmRWMtr9/9fKnD7O6bedCWWaZN
C2yFqmdHIQL2/NiNNUkZcD7HikG+m315UFRw9lA1vkAriIeSbjrjNM+xqo+cHQV1
WjhQNYlHrkJsKIVuHlcLwWeCMV/3wfDrW+XM+Y7JOhIV/kaoRbV/Ld3UpLzSrokw
qKPA/zB5IzCzlUm4cVBZu+04Nj/VZCsUpM9aGH4J/L7eAxEXvVKF8hxF1+waft7P
/WyAEYOWICge9iwmQWXkfPOS3HmN/5ApMWySFb2Sjz0iXj5ILVbfUTbO9XOhKqMj
ZAU1En4rV7RNBdtcovxVV4rLpO0dkKS98dDdbnTP2suxRd8/dIXNUdophSub8Vz0
3tY+GXh1dx+oRPIuoco44ohlAgyJXXg/QC5h1NlXP3ppTL+CviPZUTDRfIGhA5kM
SsBtGcUz71klHN1SdW6v095Uec/cnNrT9EPHyes8I4SwGs98ZRn3b0+hKSZh6bTC
yyw6aBZu+uRwdQw1VWxKNSte3nYV1/p209dVYkGvcZztGv6D/PkWPp3L8FptOG94
jBGWD2CscwPFRXkR2Xy9SjCm5H2U26S0JNhwsQFc/S6R3rsG8Ao9PRmQUkTj43Ot
Eu91k3BbbUirnjhP87sPgoS+IsVb5lFjvPLU+Vcuv0y2MSP6T68pZ/O5jYfe3e3O
z2RS99+puWZ5y7Uim1Nx8GpdMF7QlSjRVwjyxIoVt/6KQmOMiJEF73fWDrn4RnhY
eDHxFWhqYkvZ7B2PXrkLe2RyuVszhkq5/BUylNL9yEiknEzReSl0gYZMo9F1Hwxg
zYR57y66miZ22nXdunXcKPhVi4takCe64IE0Zm7vwQ01+Eyao7X9a8U8Nk4zzxhc
YfpgQkz4YKgQ4LmL7hQPCPparIeMvs6FvwWevFcdMwlBJ8lB4NFSm9t7g2Q7JOJY
T8CM+0itIRAPfNcUn62BTiz4TpsZeWkb3zXvLenui2LdirWfjIr/JYSeisscEjdo
yhT55bH2ms4W3yvj7kbApL1UG0aouTdIche9Ex7zMTIsilHSUl3kIIIdt1SuwHJx
a6VplVSvhPnwOZBxAV8zZ1P6dwJ5JLYlQSr2dgW8nuw2I7jWYUu3eoLgF1OnTkFs
ZvDvb39gyyh0qQKSZ3jUjLtLlxzHUo3CJS283Up6bFq8dFlzPZXxcFErfqk/pNw0
kn0qAyLWVUhzdAQ7vagd5XygINNEyDfsvRgb4YfJ0uucEsmtZ8OYYkaLIrBTZ9Lo
RMo1IDerdCcy/DgCrgBkw59PW3ugDSzWMOuPY78ivNXESA3jK3+aq3kJGlMA3iBx
5vE5ornujtmo0O4WFpAl1nzfdM4/3wsNqd/UILx+i+IqZUt8NkphJe6Aw3jmX8np
NzFijYZa1uvqWkfNFjgKFxeVy3XjwqlR+cTCrQMfvzdP1bAMDHJZp8YkgBBB6wxc
WTBLZYG8CcPj7sP1jshJMpCTbKTIJAE+3Xp3twgznJJooOg+ofxdNPPWD/yLpsZA
jBTXk4OQznpa2ctcx5tUVhzhxXVMv+wuQFkeTRL+ZMySL0aqeuM3kzEYINqPJ9DS
TWeeGsgvpz2QUQ60dE0JyBd+h6yP5A2Ltpq7BkfiM0xBoKWcSro5zk2WogVaoa6J
Fitc590gMWzhflyP9L7eZXfPuWURCt9zL1WhEz0WXA/h9P8siAjOZE/uML3zLmRL
clLzp7KnzkcfmwSXa3Z350cm6wc+a5D0AL7IGoC2S13jd0PUj7PDN69aoVp/7Hz5
1itXSCNGUJ1j0NL/AvfOAjHIgTtKW88MOvQkH6LWMjifrrazyA73a++Z/NJ3ATEC
kRzo7WpbhCUjBHKbGmkF4r9MSKEGPpAZw0jstpYiGwzAPWO1dUdZFxreUWkWu4fO
08auQMm01HNzdWBfqjrNAPeJuC5KiggA/9cmi71LWqhQ9XVKKeuu5uWdGwqZWzCb
MfepigYaUMwWocaxnpDJx/lfBsx1IdBTrTCDDzdK9srMASgoHZ+p+AjpfpNc7+78
h5NBYnHKBYbIuDsOKjydy4wUEP/D70C2D/8Bl3EFyffhU73MMx2w1ayG7CQzPdik
Tqwwn3XE5JF72pJ11oio/z+HYT2n5lAx5GvE2f3SXvJwn9DWAV1G6IyW6w0xgAoK
9wW1xKIUyp0Zw0jUIzAOyEnopzoYXxGJFzYHvxlrG7rYt6Sd0WaXGgBHxwYGRaSI
9X/6b5agTGBQfY3Z27dhCfdqZoGq75RM/yKrLcifdrDEEEyBpqfENgHXmPCvVP0U
465HooeM5Ex6x+2/nL9XrWNkFvEURoglBrWMUJKGISb1b1YkWsL51Y9ZK1yIF2na
k7MApC5N7P0Oo3wHFohiu044KAq4FSX284F7ZREixhkSqJIolhOk74qPSb10FTxW
HSgQ4u4taIppsTkgAM6iQnq3TbqfpqcLrQw22YVNfqOkr0rVQOw1F2ccgUJ0X25W
MlFR+BVfQhyLrd++QoVUj1HNp0eSAHflKWNh8mM51cPMx6SIvu0csAMPiUf8X5Ym
XR9OWM9wc/fS9w9GDHdj63pmkOtFzbW+lt/r2SRXZ7LwdcJH7d+0gpuxK93Eqawq
Y+Sq8nqGSGSkN8ba9PVvFBeCbMil4J9o+rhdaH5VWIRisDAcnhi/ELGt8OFydF3W
yja2YxCmswu9mN3buOg4GfkFyKCYUPdjsTcHG11jddHgGSnbxXux62ReyJeXfSwy
EsTmBx9rnyx6lCoBCSACvdqFIQIbSgshM2kFwIfZkG+Vle1yiyWy8niuv6HKELJI
6EI3uXFNDthoA1+AeWueolde1CYjgh8xHgPb2Bh9lpZtXmHcMngzRnSyuoGH8wEN
L+dxqOQ03zRf0akWvmF5i+HnIlwi5Js/1NWRymhba/KQSK6alGfAbLjnbJXr0BQ+
pXyrsOZGpB4YRPJPxVhfYRZR76GENgE9GqniFkI3570x17uLarsEImASIrNsWFoT
AGqW12ZTXQhkBXu7YQt3PCndgb/1WSBvQ0jAzc+Lu/Y0EX2O4gFDRetQV4HiaS4B
5iOL0VF5Gt4af/iiHJNdgvMaMoFNassuLtniTmWi8BKzn/Cw7a+/A3KNPHwlubR+
zWJthgA/OT8tKuXDvpfoDPXXtAfPpTi6eBOf6GjHGh6c0tuRjkMprBzK22dQBNgK
OUrRQY/e4Yas6kpm0BKfwe9/TdPtrWLjmBj5H3HDwySzvoaTNSNJZpd7eX4wob4V
214FJNAq9FSIot0t9R8aNGMNtJeOjW1UChRHROZ+hB1jq+uocWBmi9TzNStnl5e6
I5mc9XT3DYjdFFvnGlRqHkzG7Nr68JH+fJ1JrYbfkvG147qtPV1/8WAAlLmpw54L
M1b5Wfalj4V9UJOzgldOhqGiDRiLoaRVz1wDw4v5GZ4Q+C/GtM29FfQ31S29XP9g
eh+GqxJOMPlMZDXvWthCmiWHVGJhkTCg1TZHTUEYD8+BsecHk4G1qX7/EBZvtoCY
uMqwvm/zQIO+DbZFAa+uUbJlAkzq6UtuM+6BekjO/tarhPg/TWDazrtyJIPE25A7
ZNGTMqe0mxfi9tzF/Da/j3cnIPepsvBa2jysRvQIzVVWTwsg/xBVHOHh2WE/yX4m
dwbI5pSta1n94PCerMNUYdaCbXA7AHrhkDb+F4Q8q90PhbiepiGOWshQ8M7Rw9xP
eremqZ0djJxGkqLa9e7c7P4vz3Jzh5ahZtUdPNGt9JV/rM3NE3hKJbxauOD77FFK
ND2ae1MLx+lcxBVW0FcUzfizI3yawMKPR0xtuOyQyoJ6qQADDnebyE2ttfyG19pW
sV4eD7tN1z2cgOXdibEXbanHq6UzIwspG6U5fJxciy4KvwOn7fJmm0+GZo5H5/Tj
yOuKcFcKTZ2gDHcjPA9lLvvv8zwd6kPj71gjr743ye+BnEjU58E18OTEFjN425/I
a+2sZQ037YnJ0YjrcBZsN4bJkEoBTw+zWz8dyKXgkpRJJ6DxMfsa9np92/6yKSyt
/UKScCfp5CI060RCIkgW6xenBpvykSSiN5xuOEcXQvZwoedL7BIYuDFHACFHZ8Et
EAP/07hiZHKm75vS1niSZvoly+iTbA6iOO2nvC9gKBWUV0pJZQ+5yu/UQFs1cwP9
7oeAziz/KfV42ZWPqUN3bJTFMdxU184g9TTgXWu6W0/sHyIXLlLt8GyKKnCaJScx
I2k4qp5BMFO5Q72lDThtAcKw1yHAN3dv1Bvfm/dFhd4pmvOvoRuaQsz/48yQnS3F
mc6FzH8ss+x/3LZsWczoc/1o0hl1GOVfyhWRafpI9EBSN/Uv6y5IqUO9npVCE4Yx
rwFIDzYQ7dEvlJUfNvtQHI77v0pphYuJY6EkKan4BaXKgwTbQWcxrsC7bgq3isoV
gKpmCLff96UtBxKxSVMR6T6tQ+KF2y4s7BeCCyFHwafLVXuNT5aGjrlfghwIAJH0
ScKGH7eJCTn98Sm+0U5f2AlwM9bGfkOVqb+DjXLdbjaMeWDAg0+zjVUnz6SD+Kro
+Ic1w1ygVaamjbVaIpbyUAZGVjh8gGqw/lDvJFyb25BYcOBrDwnn/kBLKOWN7Rn8
CUBZUR7ujKGjCpAURywEnxX0FCL2Z8kWnYruc3orWR0zXTSaxevmvrQWMSyl0pxQ
Sd9oRhyivcEKKgVY82MMDp8PxlEbwGx+tHY/gf/IR+D0BLZz+Y5dN5OVXxYS1U9A
pb+gK0wSb95jpJKdBKzv8VR5oNMVHehNXafejrAoZ3tl+ANsvB4NZSuR9A2EzTjg
L0v1E7lI8M2+ru3EXOofSq+kZ3YZ+4XNsIEAt9oQ+1Ats2v7H98HqwO2gatBAClK
YzvrMET6/CsQoJiOgHzy8gs2i/jpDnyvJM28pdAoHI0oCPHFyBxmIodVLWQ1PecY
Y9yLJDv2EYfXull12GuXYpvVfSI0jL362IHlXz7b/qw2FH+OBcoqYFhIheJJfnIB
fTEcwCk/lrrxdOvBbQ1AG4aePpG1rnH0SEwWf+dYjBGvhhISw+JqDixNGlqDNfSy
lzzjCxhtcz6JwY3g1O0vdmHAyrcFB4X3ssc22HcQh7r5RmDZsfysd253qUsQ2TFi
f2DaukeuV3P+FpP6zoK0bVikn3ENmvten9kYpd5C2LZphq9eVwt8cUaWKNaq8ZW5
RP+Lc4+TUzSdD+az5E5BEAXuy8qphFf/gBxdFkWOJL+iLPt+kTq/KwrZBSbgySEK
Rsv/6zx3OrTSQdqwulxyZFwHRIAonfUewhLARg8raMR0IiTFtoKa8e4GFH8EY3Ux
fnR8mr1jLfKtR6ctLtHdcemVwRu6/JfVNq65RwF8WIouCSf0Z2EuGxkDPVdjhAJZ
amxmo7GbLrMLQ8so1G6eF+PL77Xdoi9dhj2BzmLkO1B02mjdQ8hDHZleQiqce/sw
kLit/7V20NWFNM3JJdhdOZ4EqxAyJqF1PJg3AuuL0Frposjk0aGFvrPVVOk3msSy
9gJoMqzYevq7fVherSjESODag9NXyk210F4ZrVewwSxyskNgu5PiD7zuew05SHpj
ioDHoyy2E39i3bqVHrUQgZ4iR+xdyZC2S9GLim8vzHojy3ALH3fHHeFWKc2xwhCP
6ZDBcz1qXS1sxFSm4TNrmhwzKQw+er7L61sqEeXqRcG7vNWcuUnh9b4bTYZLDXjq
e4CuL8LCssGXXLNjAbyV8kLm4jeEg10ctDzRrho5g7xeZvZdQCj2v4PqHUM2ePC1
wvmEO7ECgdgsI+8c92+9DJzL09MkTqx+ZhJaFdf3g1HNGEIzfTwl8Os18d5oLUVH
vqXf7p30q431QHf/PSE5H/+Pf7nJJZtkEayZiRIVKZ9N7emtr5QdOaJDTGvhAwNT
ia/oeEMzuwG9h/E+dQARYe2Xi0ZM6O10CAnYh/bjIK5z51rWGTCwqRdQx9/zkq67
kQNvWdT6R3g6gkXHA1794hbuHte78iMqcUTAa4WuGpNRAOQ0FYQ8xncgUgo5b8CT
PX0LeCBSTHwPZcUwTpFxrcsIIHTueHizYMhTvj2fN3fdb8E0eR9o0lyVF8JF9Uka
gXd5QpxrSvpXwcDk1RRvWOUjRynI6Hf0AxmVCbO81nyOPeaW5vyhNeyOAirRL0/r
yj3WBY5/+4S6L6fu+aH70kratf/c5X7k/ZS0j5Gucj9Ly9t+rETZTKCRrqcF8n6R
3f+mzMKjJGYSVHR5DF/2jzin3ewvoEPQX5iAbHS9Bx/OKabk3pgJWJduOy+5+hDU
ISqQ3zCfGgEnjJSuMZNt7ka9pQomvvymEykzRYz2rUwFe5VsS132YDCtvdYtEDk8
nlv8oSakexwGGqR38LumbxMMt7Ak6qfncMxuHkpXDg2fPt7jpbw0IqiOnwxvcVdC
/mAvD6c0d77ecZwiduXmeIoRzysJX1dwyzLEkrXL1uloR5e993c5oL61wkn+cHxK
vzkv5196nTvCnHTRSi5W4FeMRUR1+XvoJvzw2V1nBiTDC+9rTcUyK1dX1dTRSCzz
CcK5LJZhh2qiGilO50OBy9ssDOmtIERQjyZVyiFB/Rg11yBKY8oh+cUxhMZWk2o4
Co/KDun76TAlK631JC6PBXWjoyr6ER99033snsO363y6bifecERt4wWbwEP8WIDl
AgvtcZ8yCj6NLw8icI1freeHpSKuqiO1q9KoqPL+ZwanbKceENSBGVO1NyqDrICS
798vNfdaJPaLnIjgt2pfd4THuLmTkV79MwdUlbGB3cA3G7HszY0jY96ODOVhvhwe
yHZ5GkN+avBJ3yHsb6wEfaRotSXAPpXqMr7WiVVB8UEi3OBt16nKC3wqZ4ipGIbg
Qz8D7TcaLtigCUSsPNj0XHyQQjYn6yDNNay0mz2W0vnFgKR5ixENu66NRmQ50TJx
d5GM0QAcR7kB55NHVsTTo3AiCng5w0FhmnoHdku55m5JNBNv8HPRyBdfhT4lsD+b
W7YjBQNJkM9SUaQfdbSCnZKStmTUvBwoiT+PZhyUcg/xp2JOZou/t8mRkKop99K4
yKHEoW+vGRww8sl40hd94AtQ9ytbZRJudzSSGvuyj4ctNT9KODwCGienk6IiSW2x
zp+qo9F8zme7YeHfoF4DNzuOIvFZjgLJB+/ZodtAejtO5kqe9vXbqU7L+gKWR3HJ
9QlywvmyQVsF8eIPJX4Fz+uqsmNr408/bmNRFuaxDXdzGXMsiUA/EaZ1MUyIW37W
aXW/7tMkX2JyQu6DcLyEDr2YmzSnXqTakJ7lt8mJoAFeGhntmb7bVAZd2/38hSbd
8dYNHOTRNkUIQb9uwghCGDXOWOch7v5hXlKP0yGOVGhIG6GEDFDqWnwfO5GsVPQB
zy2yFwlzETvHucFvnyjCV7XzI1SsCYu7BXj28O2cLhi8oVHtodxE5keK6kGt9cbx
wCRvl6pPBkMj6i1diPt40uIgh2FrnrbVPF46kCaHVHjZ0EJp3QTpy9tcS6usuxe/
1HuxidY9NTVSU4/6YVBpkOZMFgT0yoXBh7TIpKJPX+afk+FDi0uDNkqbgNF8MHyJ
2n4XIA4iFKhEOVS5PlrYPPxdMZzraqnNdiAi+0XtSxX+oOfvkfmUeIf6bcAARkFs
16zMOX/UHLMhDUGvPpPFVf/LBxxMEca2xMsAXJG3rVCBNRJzyaPigAZ6hRX7hYGN
G7IUa++2F6niOb2fhSk8lD/vUYwPK3QFM2Zbjy11xaG5LyKYy0XRDCuA7mhuE9vJ
W40gzoBADmL4v+J9VTV4jseWqG3rheLr6au8F364hGKZRdOjsXsWzVU+rFDdUO/i
WlSfeqdiG4KwCSSCuVRx/8xFcG6a0g7ai7KvfI4ozrLms3/b6AiqpebVKTXmWJCI
vvmSHeaWXHR+4mauQfo34pNo9/vjapQGelE4juB6ZgjjHoujyyX9B4MXRJc76Kjb
FQUtVisJC5spfasc2Xzxewmit0oafoAADMvIrrKMT1eLUTGOoGIE0xE3mJkfYW1s
1alU/o6Jyvpyg95H4lFxLbI1J0MoxjG2GTONELl30hAP3CzS4KP0q3gZDMbQGa1/
+rel5OY5hAw8WexWT6DbPYPvvlH6wGUcYP55NaOMmOv3Z7QAEdppqImi2y5nWKwh
AS8TjVDhkPNqpes/keFMjVSWSJotxl8oN6SHKOzgunflnX2YDg5zb1CCF1DLclb7
1ncTJlFEEOKsThuGcyO2rYB86iUpydzD4QVLfwjTRMCjLEs/UWgpp1fX8LeNqvEX
aZHiq1w2L8CBbd2MimzFA3NNCGhTgm1R3+Zd/YAlGOZAY/ttyWUa88ru2aegBjuh
xBmujEZNRFIdShmfawKM5Qn80LA7PdkyppaI06nzc38MQhmFH2n7taxo7q2baXrs
VzNY+Mkg1SyFzPa7STf4ZdotxqSCRHyyV9y3+XndVrK/0quTcn7WMBWbAskcJv9G
gH57hTxkiETLDFI9lyT7CBATSIsnvUnWsrvdYX+hpyixPtl+6EkkvdHVr8sKVHqV
fcVcFqqqe1+SqN1fkswpbiVb+H/GVqUnM4S1uFodH/w1IkyYykdFZN02FAZNPOri
0h0eKdFP07xRWLdlzsp7+cS+efWDQ4ID43rioEr/7g+80wcoZMnMKIxbCIwNNy+A
IQmg6vMJD/MlsaHncY7IOzPQfzxako5WGRcAvQU9sXWUCMgT0jp75ObrqjA0cwEr
Q45pCxF82CXicnVqM8og5+7BfTD5m9uB+TZETgsCYbv5KUHWAnKBZ9f3IjczJz9z
YIk2dLGY4pS4s3d6ZdtjAzeYalTvxriSyOfTi9ZcjTiT8iCMuz7ZU0H9HIIVoU3z
X6c0/EXhd82rdxdH4TGAM7kw2NJ3oRN68f20tm5ZlI+WYOH1yu2EoKVI6Ln/0RRM
vwHcEycski8gwR/TBM+QOTTac3hBrpgg7VqoN3OIjazLlsDvpfBzKgFm8vjuURDo
I3cdIFh5VTOH1RoQnfgm4XrqN5DVgVOPeczgB63BovJ/r4W/Og4ArHbTXEPnxUJR
5HfbdCq7cE/CcY9vICGUqHVIPU0h2xy0gt9m33yeKlgiMWZV2p8GatMhfjVxbXoY
gz9rF/GzKFlFI2tk/7XVt366M/vdoiMcEM1RRGskYoYSnHCWcA3BSmiz/1itzeAe
hNdKvLG6m2ZrHEIaefVL453d87qGrU0+ke6MllKQROD7ZbzQz202JrYpRuhTHNn3
Mr1KdPPYIep9kEVMza6yi5+ws22SASA7LWmpFYfFFdxUCNMK8QDgHh22OVMJKAiE
f25iUCdwK5DULxeQfAVYM7B62jFV4wTKXT3q7sudmemgfWmioQk6Ae2P7+rOPSRu
CwR+qMlDyheEz7OQCa5ZsWrDfmm7KhFq1KLkp4r4slka4E5Hxh3/ivwZXaM9DwO3
fU1Ahbfai53PUKKSeN05CjVbVam18dgBxo9ANL6SvWyspUmnZiGTJVt/TI+gQDAg
krQO6tELvxYTCPS4xKzhKpIRxlviW1F3I8c1lomKUYXJW44HdSkpBhWTkuP3fvkQ
1KebhV+FbPlhsgrSJ5jD1goNQriq8Kibiqv+A0hMQeKoAs0gT3ctixI5BwC3Kxoy
Zn+BjAKBEQv3P7gdzWyN5TTQiIe8WEkyLWAQ/pGpW0HjMelFrLmjbZIqfywYfJ8h
C9NtZU8c8uWtmiorwFnO9XFtj0W5rJjous+5WOhNv4mCU8lrWg1G41T8og5t5rvR
MGf7wZO0oPQxC3067cwk2bkaKxJOdpblsjtyHLQts9qbC4nFsX/jxRqPKTBPw+gw
2hMBTmqJN9o2BgpEIWHAFs0FV19VpOyT8iGffjwMPSPDIA6HhvbtcLvsw/eCXyz3
YfqPvnFb8+27NsXqjIK9yXPWxuH8KjkaNnMdlxvd8Vq5VlXDkGTsdu7sebw6yTOb
k/8hSJ3bCZB/UtbWM+JtfDukOsO/Knn9F8/PWpkPOoGBR4N+MTEwJIwZYs2whCv3
yl1RDw23uzSORFxz51F+8eWYztrtbKbtpklinbWGERDuYiXEHUY60RP7iJ/A+I0l
2h+NWe3jawCZZYC2V8wBoHUndv+/a4guS1cGIpQlpMMNhtYVpyttlOnkDaTEkUix
dDz1BDnrHjGcnX9o7foCeNFPl3BAJlF59MOIU89OJeAuiw18OwY/nZk+CLW70exV
lOSzojk+/mUEyJsY9KcqgXojyPvCuaCHI/8tniZCvjeSBO4Vf3BNRRmTFGYDsBKP
KNI5s9EuZUwQQGkCh/CbNkveChn/TbZoKxUwTW23+cSN5day4LZG1ZzGCAXLf7a0
387FY3KKQOnf3J3ugx2Tut+urXWmqjWnDJR/raE65bRExCzSzBR3wMYZ6KR5eIjq
Ps6AVPidt/MdanAMefyp3lrmPnF0dAhPb1dOxKsjSfwlMlh02Khd6nNO4trcfM6I
hML+kK66BoOsvNd8ZCkEhNCI+gqOdx90j/c2hWTkIz5HaPwMPh727GI1e1LerD8n
L9DuPx+Ij4ihVeDG28Ex+S8SXGkWHr0DmgW51eppxEVJw0YJ1ehg3cy+jMV4FG/Q
Yivydj5awGMyQmiSB6NphhpS2h1cFK+/oGn4s3zHBhpXaZnI1vphEfAyU+dLc4ae
HQPOe1ruSoUoYtsh6RHjqf+jjg1HSJjgvofD0u6sGjJ6fVESZg4r7W33jKby826P
xgnNE2yDoG9qrfubqqPNm5p/M1OxSqvkcxp7nU+g5wU6A1iXgZ6OUIPCpjaf39D9
zzLbkXfq5KDP5/1GldtjoqfDNm2oh/EK9xXp75LevqEvgJ/eWsbuDG+EHF63TQxY
LLNPvhx+jtmzuf66RybM9z2lBWO4m7Uys6TeRhvwstNsw0yLNQ+nuYR34kMDinfN
PwXbOJpgUVpI8BgE07K5bufB46MWhmJ8elNnCE20jyBbhb3m7Xs0E+zbrqncVSdg
Xtdw3Aq6FPd0sKsVFQ2vre8rlWOXoZcAMtssMcbG/J5kQQ7j5efJWv7Wa2AIvZVt
DwedJDCEAv82cxuVRr2L6TQ73IO4HNu/5ZdNTdKm4OvYWgYfPm0Xw8fnv4oG7YlJ
bq4324FPMOmtaZm+Ovx/LaIcTrkI+PG3JatrTHtCtim7dFveWsIjI08yC5aZLQqA
jRzCB08XZIw22I+QSgy+7PspotZ3+5fGAktIPXe35Jz8TYa7FHPV4bqcBVPISnzu
fcsgfZ61gnYV++l3kllNI8lUdnthySwbXQyct2jn72fZdGryY9NIuY5Hw8sztEE7
frxMOMhvpvQ3hyJ+6QUJRETe2zkb19gj+d9FkYdPANnneKZw3hc/NVhShzKhgSAE
mvkOW4RsY8aJ58FSKMH/jug1ktyXr54inEWXjYDdqJ7NccRwqY36Hcy7ej2i1aIX
YqqKysq20qMkOQ47Hmnsl+GrjWvufv/cz0Chdstvk4iHRyNHLIgknKf/Ls0WuSge
Xvjq4Jbb49L9AK4Ba5T0s38YKy1ykpIrIahzYpaFIJaLtejXwwI/amzJhIBtadth
2AYG2byfdb/WufqIROzyPHtgwhGkSD5I5l4gJOcQMJtkr1PhGhXHbC1whGKyjXam
laGqLyKpqWhJXsZgSo8bvxosCaZBPKTpdo7EmefAU3NtMYVvVE7hz4cu94ePHJoU
EyxzjlpKw5yr08F0g83gVfuvzeNsXrWVaP+D+IQ2D1TRKCGhNmi5W64pFOaF3hem
XsVV38UKLbLJIdYBCRmSAHB+UkZJLXIf+sjL9nlJFJRu7alU249U18lWQlf20wlK
zK+aj/2tJ64Z0qQPTX6M+TMxUu9r2U6s4uEFkSIXw/0mvoo2s+12uCx03sl+Q0lZ
D5X6+R9EFKgQlOVS6TS2ehO0e0lkokHM6lzOnm2D+WgbkUOyBHmxiHzVR0Q5DHVf
Ct03tr8x/iDQJULb9LV7TUUJghSNVBwY7AB3JMgPN7fZLpfSZyzgHGIdmKOrTZv0
t+AI7w5FRjHLui/8zT7XZdGf2yhtdJe9kx6Ggu35D4pNy2hl+afk8JgdVesq73Cc
/ilYSgWAHARmnBxqCOfxkEIy6aMi1FYLIHkthA3Qhsn2cqsZStS5Qn12VjHrzDtD
EHF0h1WghYrRijp90bJ1H4tpxc3D1F9KCDbTEd1b1p8ptTKF1FyeFPHLqj0seUAV
DFWhE400pfB7GmbraYUrweDjF4M4DuFNnfbnyAl5fwzS6IDMXD+saXKptdUJNe/+
G3zaqXPGeRXK8dbdFSMSgZEoEUoNHivNok6S1UmhoXeexSDqDP/YAo7Eq+fvqhxz
Vgf6iIgy2x9Io1etQ8tgxKyiGyhkLqsxwfDud0yIJO7t3r/BYMnm+t4rSzGVqXrq
fJaM7b5b7D4OV8DDG1BHxyhfaTdR+h718Bszrf+KhS7Gfdu0jbUdFqxYv9n7qfP4
b2sGXSOHSwqO9A8lNAbwSUgIgjCc1vBoAnboFvzVPVoTCohh8p+3w84M/jHfsi3I
wGEp9WpDGJJdVVhPzZs5MIm51IABQbKzrrkc6QW8UgXSKIPMA0olJLs3WrN1JFn3
WYoXhrvsB5GA9v8BxBkxyWlavYkSMc5h6adVwEa//tU3NRtRoh2FaOy1ADRWs8BA
onnrBZxaSJxHjGYkM9oUr0Gl9FGBQQCUDQtb2dJ6tsLAHukQwwQShCj0Cl2piN5o
Ec18vt17wQaM77Wsmx7s5ILIjiAG4zMKrXpQJtmfsNK3v8Fzwdvb5CZjLcYQ+nk6
ll2aHw9pF3fA9ebp5udFOWll2XxEFpfbXSFAuC/9vCoecSxwJ908eqcMSr05w+fN
nDgR6+TlwGgxMQWfwsxfZ9lBhMNzrDlwSTfueTpSmlaO5thht33ol3mMZK6cWK3/
1sFLIVnZ2ULUCRofs1RVx+VVMGWJVa7CsMRI1ESOpvX070dNlEBt36NzXXUOPm/X
t+6GpBqd7bmBVj24bo39fOvlKZKa3IWi/p1gW4qPQtCt9ex5B8Re3USz+OGZrmwV
nK6HQgvbxyDFZuE/K9JyhW4nbte8G6jGM0cApOSqViAsWREiS1Gyq/nqXfQdnzcg
4/QGLae4HawDGDaAqMtpwcG2ekMVITNG5jKUyyt4rlGtXLAC3yacuFv+bSQRNrQE
XDQXYJmiIDmMeTbv35CN3bbwTeuZQPgfLRws+yZJ5ZIFH0xBK0Le9AP8ZG+6cfHC
TawfwQJ4UehxqqKhG5ZbBRX5qECSENEoGt0blCg4LA37ljelCJk0oxfev+TygvTD
I6CgTrHncRnk7TOEC7Rj2YJKrqbOaCrY9SQn29snKC+ok3u3Lwj9bb7g/LhhcQL3
jxpvGAvkOOKggazQLlh4sajrfGO04wZlTwS+G+P6IU2muzYoCNUvFzLgCJUKZHuN
BJ1wx6LGOdL5xnR1A4aaAVBjd2OFFoi0upxzl7OQeQOa+bZiRlqEHk0YIm1+hZgL
y85qPSRIvX4yQgujdheaXUcE0fq1Dqq9G2QRAsc1BKDb2ijL4Nax8UjQOKtsFE6m
17uZoElRHuoYvnyhp5+E17hsKHrDQUzwkuue/K7gXZPV5GB7cUvEoYRFhJIFaRwV
RY1MAAeBfQsegdYthUJeCXHNU4R6+SQK/TB8wddZBSO+4ec+ILRXt2yvwNVgESNP
jHyH6OfI1Qlk3+mt8jAHahAVpF57DjQij42eymZA7gEcO1sfXz0LTr7F6LDtc5GV
3tzFO5hJeflL8gx9kPNCiYhkG2uE7HGng2p47LY+n8US0jA5L/WoZ6c782BBMqKj
8xxjxB6Xtiu4gOXqyY2TIRolC9icHw7hIYA56HCBYdv9ArXXijoxzqtYS9RzR8rk
i8PnEDZFaL8s3qnep3S5agvqgnA+cNwkkJB1ZuhxPOuZ1XjkJlSPXpVwSPR/15aQ
bkxdKC2HTWHtYsackKXrwSajQf+vlj0Rz8GpmUyyQ9hcxyBWbmhYTKqMT/xt8Ob4
VljiJfr7fr+e7rbWRL43El7okDIlDAnAZjWCmdSEl2YjJuMQdj4tUeBKOzKWz0be
fypwhdtUbQke8Qiye8Zr1OgI32hQU0zB1aaTKSr0X/z6JYgKtDOlCxZsNW+fGsqp
ZocMd3INzgODKEPq49Wpk5jugV/9mXFL2MAfCJ/7RZQ63oLBnpiRVTkAm6Ah8Nrc
/VSvwv6R55GeMev7yf3OPcXzu+6IUHkeCP4WsOuYAegHY/BCgO02DKXs/7uAN0Dp
kv0kmAz9S6EDj9R2WSsvEQrFkkvZ4IW046vTGmw4ZebdUsSm4nby4/Y/+oq/liMq
/E7uxTeU9T1kPeMT1jweXOiNU1R2er6KdUeiu97lJrFSy0tQN6os2Dx2QXwB19Rd
rwhRTnuWx/Zb54HHIgyHP9VA2pBlJQyyva02LDxd3nkIKrVD/vLs6jAcqOsoMVf+
dM4isp5Rh4+vrqKTrBBhwReGXQf+qdgLKq+VZKFT4sye2rc115+w27LCHLsP8sga
HvX6V+Md2gyJtmo5dtlMeFRWI0BdP/M0s+s5dZmqc6xnl/BmzDzyBOi13GxfFqAF
53zWCZkgmeujUQKhrGC7sgWX4VoMVya19h+wCfoTXyD4Pn9ZVOwf5CgXpfeyy0rD
U7QT+4d64WLMS5fNXCm4mUz/fFhPdvlZIIPSBJ7vOOVlzsYwZISRzeU/oFaAzXKZ
34/5v5QHMhB6kZrKdKx09gXMC+qE293gkGgXDFmjen2MZMmZoZ/04m+5zStHanFZ
55UxGdGYHAFtXDR+s71E1AxwCVTgn0vz7jgG6rGfJdPldj02XKTURk24xJc8iaOj
+OoFWUVS6avjdbwZtnzte+CPwYprSx9qnde7wmC5hSZd476FHdivphQGzgQ/ayrD
63afjXgxol7nTwjdflcWz+QCTXlkd2qBBhaeGOgNHUpv1KPl8Ys1lBEhYsc0uIIG
6NI5R7PLKZzg80+8hvGWC2q1xx9JddxTWqWFQI+Ij+6EzZjWEIE62sN3UQawTgXF
Kb4hj8KSLyaeda4X3ed5bkSu0GEIgVElAK6Uvrpco9wlNo+h86a8bS0TxfO+fMB7
7u9mAMviFPHZEvgi7Ucj0U20lIcVnL4oDGSI+sx+5hLfpeNug4vPOlRvWxDque5d
s6VJwkbT0ogZb4TuI5JxTEBIwc9H/qJPTgCkGdrzCYsgq8X9xu6ENFnh3YI5/D95
YVWJr97wO+kgMQt/OkDAQGlzTJzqo9P5Dfo0i0/er4b1lqR2FS4MYTwnDnFdviHO
qecT3sn+0EFWyMFJIQSGhNx/tR+53SNP/TryKD6v6Hn06Pep8KDCdtWVENnyQYE/
iFn0/AeWZyCTYv5N7P8ViDQ4esHqw6QowEjaRXFlgeFIsQVC/3tyKCNDgvdfksxY
qhaGrGLymWAoaD1kDcXGGP3i0STSziZ3ZZeuDk4/HmPfpyy02LcPQ7e1FqV8qtBZ
Raeu4aJ27vShw3JpMVDneahGJr5rzMrVkuD1Fkn152S1NqotfbleJ8dgQRWcZkvW
FMIa0tpj8u/dPwfh5Twp/TmFrd9v/Ow8zk7xJa60xyEop6/8Ks1ZkOwJB0ULupOr
GaJajXM2zzxIDeLkDUAaNVvzRQmroKkXDSPfSkoYnmBZBI773PWFCnO0fSNaSNfO
DJdjBIl4Ui+MMKVSeU+ULulfoSshA5sAjAd1FB4YxtrcPazOe1/T/NVIBWQD2Cki
7w0pw/fGsaSmVi3Q8Rhib4wymPuNe20NTIarNSQlZ/VDO1SSpto14cIilc+O+tDO
jgKpfFoevBFDnaFyikEgeH3PwJu0wwTE9GPy+6gmaUHHjzu4xfe78larAG2thrC8
ndxroBw8DhQn/wCXLZysmCSNxezbxFKjjvqRKgRLs0YCcmiT0zzHjX3+Hp4Nyr79
WXbVkkOIlfCEtqvqKLw+XLxAAevdjHUdm8cH+fsuzvdecNXw22glkVt6PlJMRWYq
oNX0TgkYa/pLluZYhl6q7yTShqJpbY27IBghQTzjKLLMn9fjviHz8vxSovAq1lE6
ArCba3nU4aq85v00smpscgnwXc8RJj+jmNXpJuDP/Hu7HlaBcCXoxzorioY2/5tS
6gLVRuilJcWcBUy85jg61t0PV0+CXN50qxJdJtfmfgKYqwiksImMIaGK5l3Zl18p
1jqSzXMYazzGcPNrOU4WWqE1D16pCtMU81eqNKH9ptIEPtSV4AuYk/UWwNFNss+m
D6CTTmFiKoOYX3qRNAO46mOEA46WWZqLD3BLYJEeT+h2pjZ9LkPuYOa3GjmrOqXl
BpZUqkP1ldbQi0kVs1HnYXv7uHrmF6pZ/ga8oRzsTdo6o1CFVl4BmcnmSwc8APfF
oKNe/80YHpR4mIE0P+XwTvTJaDkyDJ37dTO2PRY1uIYyjhxuCDEEcrd1Fly3yNQb
DW3Eec8gnSvQbgLOolRoMbvKVWonp6KIQda3VRelTzQocz1UVjKDTjv8ZPtKKGWL
2cfQf7BsB+XLQd/LCPOn5DlW74C9jVwLAVUNHpA7tAAZYHwpXHTcK4iVFZlOrqVj
tkwCUj89zc0/uvTKoWEbMhZjzBugMRKQcYGDiktw5HAncxkJsttraHqbyFrwpasg
jjeQ33iqgV8FS8hbhL4MeCdK/ibYeMX+ceRvPhTOy6qhZcOXtskBxA88QHZwX2sM
t8N+nHY5I1bbplGN/wTH/5qF1v5kE08jE4UIhM4Lc2iNTcVsIbdsJUaFmSSf1va6
Q+JZ0j5kj8UxclmDgHfPSCzbogsfWipT8G4+q2wIna/IsBjxi55bW1BPBIyYqrNz
Yj361SRaCPEOU3ZHcmso3C1Tk1IZvd0m9cDeH4PVHmZP+gjfGEMyUTCYs5I01eMl
mNswSrrNsiLmaRbdSgjIjoe2/gcV8mTYa2j+WI4OSMnuogMT3xmX/ACnprIbET+i
noiYVQhvGA8hYTGCkib1w1jO9rvn+W/LX9Y56LXIVEMUoLbvfxTyndP6ImBJuhOX
GNNqwzomWtUEhO6cfFs17o6sOyPMLPPhoDA5ngSXqByShqZfNxnHM6Xaoqf9Wfaq
Qsrhe/9MiL+ncFvZW8X+fs3wD4jOjkzZGHqCrmfZMPX4dmoD3brlQYgK6gtiaAMt
ZwlsS1Zq949M45Gi3/XTb9420g2W3F56hvcudWwD7kB5Tglxw/TO6SfMnhZKCIyc
uDgVQW/y5cMIsTFzXF3oa/lvt8ZaF3YFdEesF9ptFQ/18NhabPO+TZKfmWyUyHLA
iS5H4ECzCogk++GXApWHUfLCrQTvTUf7OAvmEaXfiJwASGUoOVvR4syBg01VMMj8
CE+iQJ48Tk1UgAxDbRkApZF3bekThUuhdGsmXMw5ZnYfrQhkdVk+4UeRk8qg+BoU
IGAVeS5EMZpmjxHqHRCnUtlOYQzKv2WiD2odFiI5sNN9PwZIjPGhsn0KimO5IS6W
XST7wwWtJZZWNMJYgWD3Dvf9cBDhwfuOxah6pqQD3UO10bjx7g4ICsQxKIIa00fJ
cvyaLjQJuyJn+j/IUq1ONMEjnur5OlQbMLbSDyqm52hcag44/hJjF4PjGoTNKs4w
X9gvkIN4MFPL+IOW1gU84No8ik4HBvm+bYUOd9ptTvlvEf+CGlyDubhkq27UGd7I
gXC8o0pyUaEvO7Sm9xaKBUJbmfqtInIjxEKpZ0rbUFtnauSNVZYvd8srPTigRr5o
xpjM8GYhXsILFtLDktl0Hxa6khU5oq7u7ydJHPwFJ3XyQTd4d/9+laRJQM2ojJQL
TsqvmedlB56ha4+R5vZ8uhpJq7pUI1KU0npWhVTD7h+XskVR/uesWYAOv0B+6+dj
m6OLkMpHTLCd1ri1wORfOLPRcGSvwXZ0wnInjs+vsa9NZDo0yqHlm78gf+mR2YPG
RTGqBsHPJMwc9WgUskCysiszRECwzyXdzuJ3tYboAIK2ixNHsw/6KZkEb5iwZhZQ
VSqlWpp3+qfGlyNG/w/ea4C3uUm3jUjBebIgxySxg6mqcUwNoLeM/jN9GsP3YvQa
YGKUpTeFY4x0VcR3RSux3acM72gOaDIsJ8yUjMS9ATA/JYxzI4KQrP7g1b9g9dZq
o9L9x/myjeM4NWvPTNPMSHIsjf573h2DkgcV4O7w+TYvXJIpeiXLC/ZSwc+qrZoi
dDK9y32924n8ssc2FUc/emrG5hj0ebyUcBqm3cXaRwkKPWSurQraRnhkOli+pkYw
lrZpFkWsH0ERuW/8dtLOeepoCrD4g7cbZX5O9Z0TwiatAbHf8gdIW260IdSbKSTq
F9tsML12D5UrlFNLtOCWs+gaulkd3D6vPU8b9S8DLuluAa1zMLugugo6xNmqOBeR
wdKvjKMW9f3UsU19FWqruNofv4kRGcONCbUP+oARuuNVngmeC/mmCZM6ihT9IuZY
WJegH9dmHrPiccYdsJw9ZaavxXd8yaC3dNcnumIrq7OM4/hU+69ghRAe4kGYqbW2
/uNdQnOrNPrUFFKNiEG97MPD4tHnFPMFmJpcGyKePs7rIFeZQgROPE5a43DS7evF
0FcFJF9qoq5RDkuTTJIvr3KH5KY039idpW29EK5qYSUcgza9NgWI7ZbrT/wGCZhF
zYlgHtWvw9XoHUfazrlIIHzOEQNHlF4QQnGGUzt+Umbf4vIxiBsWRa9u+xp7DGlZ
LUKCcNS4LzzwW8q7+KdNU5vrZpZp0xaL4GHP6pHu7xtxrkbVgzjBsoVSmsthMvuw
Y3L2+1i1R4XxgY5iqgvHH5IFj/30YCcNxrba053GBHfM/Zw4shX7yJRO06lG+Xcp
J0dwl7JQTO8+rFxdONj3yEWJc+MomePE7ZxVHlbyS4QzvsYcroNJGEcYxhuofKGm
KaVcUrwFNBog2UTmO8ErARZpDhAzz+zm1yIFsqwjrDIDuDC7bTfxy5T+3TQC9eI4
NUrzIMskEWnXMOcK3kCLUQlLXfiMOW0PNINDo+VZd8/JQ8PXlpkV48i0CuHqsKhA
PJt0g6EInaI4czjLb8NKC9seAK+2F/k/txEt8Hm5ajyIEmJ4axbmNNFEpfbdzOsF
pJabo2dqp0RKUX8MC5sWHz2lyffgsojC8JJhfJhsf/nBP4yJS2WnrqLcoNoImPqS
3fh2BqZGxB0l1Q3L9FdZdJY38Awg2Kpza4ziXceRI6Qa0J4WkX1tDsrWfkpkftSF
dJWeMsoOkgaUkizUXVIm4Gox5rcB0oO10PkZGR0QH2FMU/GFDYKP4wlHuFSh4nJ/
wfc+ICxd3RnCgYglcE51NQsx3GZs1oViRLV2hAWnZK2c9/xIxuwyGeby2qgHIMAv
OYRhJPPuHpImmyTT4IOxHV7A95iMF2lLyGz5T94XQ4UL7XpFw8T5IjkmyrUdu0Nh
oqH0Mkssk2AVimOAyX4yG1MXmAGiCGBjlU3yZYk9RJuX5aLRseD8iGrHVRdrRW9A
Icrl0l/+knQtrudCS5jGSBPLcNNCoNqFo8100QZVca7aFCMj+NCd2UjrXu7eqnB7
MA7XpayIBGM6lfMSkqnxHODrLp/oiho+yNlMNijUJfp4plyoO1811gwRZ6hb+DUd
mCn42Lcpkj2WMeAg1GYdj1Tsz2HYki2L7Umwv5AVVEoJk0KR2yAr9TskIi70aZol
oJk4VZovE93J7uSh6vywAgtD6fo4NUBKRMkbc0Z+2hnoEEv38rHFRV5kJ2sD3Frl
2QcmOhpAE90P1hI015KPc2kMh/rPgPJjlODJ8JMEZgFR5U8k9XVbZjfPmHntRtOB
hCcPRSvT9Q34Mx3yhLcnQIkHSLzMFr722IuMw11Tbqxhwiquc/OAPuMnkE2RjSZr
qHqTXDBfWdHCa9pkEYVFhUIfAD5NxaBoObqX1Fkv6b8Out16AaQZ2ffELxMh7cMu
pdWVOFpYsVbGZtP6rsROGJzmj8jqkycgSHHI0tbK+TdAQuK3wCnjOk83bTQIvJnE
wYT7H4gk+J9PMBpFZOTJ//kUaZ2pnkVrupUGiA65N4UrVSC2hDs+AlX1zzsv/Q4y
6Pw7IYEVHsYBdA8Db/h963iOg8CZ2MiWAppLiPDHC8Axws55DQyC5b5XotsC9wOK
kxI3Fhz2y4KPxH0pHn1Hx7xOCXRUyiUOkeQpC1mYeKxT9z8Wr/iKnMdYOOw4n8H7
LiZmozpPnQ+z4tvlSH6Cqm4P3ehcxgPxe0fIDrVftzqSqecdtELP0J3JrgsjGgDa
9rnyvtGzEKy9LkgV7gcPsGjHna8kaTzL5iKTw1GL62vRu0A08Mrm5Tfe8oIY+BwN
yk15JIKFoLWQ5lIUUsFuu+vcR4mHmxh8EJpzr+LQivWqDCSX8IcURv9d9HdEgb8G
kuigPfoDtAgeE+OspmGUJnJNv1obkpcfKYamZB1EdK/kR2uryi58sAdvYg6HtEYu
T6RSLQhkZFXatLxL+01mBlOwpE7CYORqCpWrEo4QoTxfVsk+FhlZRiNEadiKEoL/
QsP6SB9ZIbMDZVbXkd5U50uhnr2PNQl3+dggp5Ki0eh6MGulaQEVYSLWzAuwOazG
ch1w0gyRe4doIyaGfsgO3LlUG7P5ELNZLNpwKj4zgBYNxkgiVZ61UyhWsj257JmK
urtBddzrMA4UPv1IzjGRDgJdERDW5//zmWhVyPSFl02cO5GOUYCwmbAqwzBCDocu
JPWdlzz3QVvT9xiPyXZcVDbjeraOETocIathRXEGR6bvgSamuj1T7NBOsNC1Bq7K
n7Izw/9UiKgEJlKQ98rTLtC/jRB3meqBq7MUZRgx/cbMHHWGeKHtjEXzw3aNJXgf
3EpN6b4nIkDV2EdieI9z+yr7KB5havA/ngbG9KCfPLkAJRo3QR4Q5P0+lF+l4Myb
neiyZhm21uOLXX4vuM8geed7ur6ArPc2OfHBW2CArTCXu3933RzPw/Hq0lwLelUV
n2ne39XEeC86r82jByT+C8mZifTmefpLTOu+xGmeKf/LnW/Y0BdrtXZo1sp0wlDV
RyI0bZNdIynh7IS/qlRNbBLRxLbxTHJr6UU2LLrdOPp/8BFBERZbU+hCixHFkqfD
Ia2NpN3X5dCCvvUv4KvYoxHT2ViZ5x66GOl9x8CsPb6lmGFFglGNOF8bwq01cu5I
B24O5E/AdsXK/GMCuaXO2X3rsxQrCqTw+acw56oE2ZpU3nVMj+SYx0sJUpybGRIV
h1CwNfaPw2CPm+wCsqfvye3DJY6jgvxpS03H+tngrzVnvnCm3uBsxTByotQ9SVtj
e9RcmuQgwRAidpYisQ2hWUXp/j9JjhBo1OHKqoWtg2AM4JO/Z+eERBU8c0I1JF+s
UbmxB8AVC3MF04uGBL7Nj5g4IJrBHDLSILcxZbGTmUjU5u6QU0otz2FCLLBguHQM
o9zBAYtv6G72d5qZwnLwxCJyyr30LHw9G9i4zqXKZVMl6QWhD7Szk9DNouu2P00z
NOnxF3FKjba3uB+gYn8tW88TkjHY2bo7ZAPiZNMqPuZOqFBRU+6LwqIGMxDiT2g2
tMd9wyyCV4m+RFt+C5iB1JhbmkzXV/Tgf6NEpyX02JON3umK7BfXi7RFPIm/GAC2
kdhzdQN08V5xd1zg1VrkLx+loxl4tbvs/kggk4K2fqY47mXjkZTgRIGnlh8iO6Pi
IyIA2jrA7u7r1HrtvUN0gN3YFICP+snZ/Xtw4U6DXQyRx6vNHASRAlHQk93xib8D
3QHY9ul1GnLTGc9GsltkiR62LQD0yOvTnFajktKFcvqpmKmwID6iCBdnvNi8p84x
6ud9hNdwQT8sYI9gKsBTOdCiT7J2Iu7oN2P6p8hx8Konur2KZhjQB6zNk2ZWAwh7
yELtBbzlBoUDEh9Xl1NC6xiHGpnDuQqqW/+is5UtLZ3EL4izPn2SeSH0qKxMDsId
4BD7ZeBDGF4F4ZsFdh8nud/bJqzr91A3GCrjfX/o5cw2pczSM/mRPtIkszwPdkuL
gGB3X/tH3c30sGVthiBd/L5X46A/qqXXzd8cm02UDvw1yXtYXc13CBgE+MAF3WNR
Y3BG079I49WUnwi8q8AiNf3MyJezQd7e4qpA8WgRqa9UUrHaPxafSdjYT+L7dCwr
82b8jCNIru8u2x7ml3945Os1QMH2jEub3JB+vJHfFDMHg3p6J2hvEXI57ibouw07
ZBN9PdJw6NDunYgexQ4tAv/8YJ0UYRQ68Lw8ezYHtFHsylXXBe+Nmk1yyCCGYfCT
sqYV81UAc4SSnPp2wnXa8s0pTq3jyYTrXeiNrPOY8D66HKyQasMeLvd5Ng8aMym6
DTFEyzmmLvyFddmw5YpPVUQbYv5S6gWhxMZBwojxdLG4kvKEOqRQCiOJ6Qwh/9mx
goEMFX8xbKpp+UJCC9MiKU5Mne+J5pPEEeDxYC9qAw8H7Cz4wZm+eRgCHPAJG2AZ
4Bt0hLiCIRzyB3VMc34zS6Yb1yHXDTx0ZFaV2mmpcfrX8QqyV4nUeMsZURfNnlVR
t+14Hm+KTitBYZ2tJb7vjMSSmUvkl8KqXXHzkiQJXB6uftvTxXYbdOakrU69+ODh
4RLX2oiqRUQ9TvuiZ0hFfkDefDW9QTuf99IWQkM+DWrvnxZjbP2Afm/S+RCWqb0p
TTwvaUQl+NVopEto7TclEbJTdDNN0FHCalG4hFzjqOJlmHRNqWOCAInE03Dhee5W
rzd5HHXZXqk0mSSlMvaz86mQPzYp5GdB6JKPK0gmzeo57x+HMOQCIBcLYusKyDZ6
4A+dIEq3XGUUD0anbTznlG521qfJPLB3/OWwgAHBpxyaM5NweVN2tJEPOjPSeWtD
+0Nk5lADwzfUvnXt9pv0bOGDnQkySwwcIjS2dbSIFLyvmCIr69wQYo2EHz45s/+i
CD1if++SDPPKgHjU/ievBGWSdX9dWPqPR+QZgIrz6WGDV03wy1t7WgWUj1dA7Unh
lPg+c9mbMK3zckiOhvx1S9UtDcnxSuAu0vwACKtKacgDsAKCaXwHDVJ03mE0rgAR
tSA5pyjWhxrV4o4kzC9TV59xNGLXWLN5sh6itJLRfqzyoFLwmRh5PdE0bJZwdfR2
hAeBRox7QKJ6gJLt1AK0M4eT8SuVKwoYevdcplUhFPd0EaxrsjzQtqylz56w83U7
xaErMdJz8SRMDTZ4W4+/pGz6wX0G9+Myq+AO8s7Ij1dowEeigVPQ5M+jpnPDzYUp
LFkaEMigEWibODX44v9ez/k8y7/pveGasacGo1azXRcsUY+ZGzNZH+YHKsDd9wQN
q2kAiqwTsFCvhENc8SV1HJSmlgwj/QWjnC7M9374w/D5Sy2tHWPhruTCiVFHdJBj
h2ndHtbCqKzk760tFC+Cv/yuOkCA0cuq+vgfA3JpM51nCkLlsrhwip1AIenA8C/p
6//s+NwTFjInOpNPMN/24oIAeFkNyx16aauY7tAM8t2E+2XEQzWI7byBUS66x5iH
cXT4x5XoClW14cFt3vz9C1QGVWc6KwjtJWCQV1T62PcBfUDGZC8az1Rm/bQ9jgAl
t1Flbaqh751uyXZq9PlhmcQ8xw4OF+mp4fEjko5nBneCtKqK2SjySt+q+UtDnRs5
hM9zhtaZU41k5fM1phMxjbcSRj6dHtweIW8ZOiJs6NuKSLmrax7jGs6Se5OQqstw
bI6dYbJjPliTr5bfTdMlT7jCRemMyktlqhd6BakaXIOZKPasw3co9CzP650PXnYi
AkzeyG+F2S32HrAF/+iklBcJmRUPLVw5lStZymiel5WP23KwWDqX5Ask978TWG7h
12qXgtFqvHSSMwuqbfW+ZImcBBLXgOMWVd78HX8VpZqJ04FRo6ZoYIzp/sQ9RElz
lroVErppbrPe5Cxs4iVXFFuPsRX4bAccMGPWJPlCy5rroc1BwCLuGy17RyhgKmzX
re5dNputzDqpLPdg9f2QoVY5YnsXoJ4K/ES05GY9BBwlgon7UGmrOsCAwvBsiad8
jcJaKgrNZgGuDAblIqd21qYl7Q0ObVSKqPI13wbsTlt4mYuVMWy4fF3QBwQqtXU8
46NEj5UzNflUsQpudgnEOvdUlZBP4BTZY2wQvnk+LYymiZyPeHzK1aNpebjhF6OA
qLnINhKmFaLUwKln4G3DAxbX2C0DnOPHJnAHk9aQeza4mAPl77eDR0MA/IUm7Bgv
t1pgVComDOb2m4EiqzJ0HJGC1vbKMxeoH4KvUyUtgNZ0nETqMQR4OcQAIcpK9Q7H
9ODAEwqPtibuJtRI4krTrbplJji2ADMa4qKZoGUv6GA+75niIh8e0J2sxdwUFk7f
J3I381mu0LTkrvX26mJ5uew2n1Fwx1c/fkli+MhTvwv8oiN8Akmys0rHyYcRsrjl
lgyJJpZkCSxz9GQwsduf8oqgSKVTiebVF2V5JTjTmXtoQn7Ped1FkPAmx2zaxw33
ijBY/CrRT+tkMqzqSaQwYQAbQ96IvBRWhBdGmBKyFuiwmZ8bzjzhxUvtOG1C4PFd
g8tsM+dLd6PTMxfzVbbGBUh6W6SgDb8Qn+mCTKArNYMGeCg/e5n7N0FpgdoV7cxC
5L67RHX668jSZ3tXsSKpDzB5k7HVvbBtUNBAZafSqLKIZRKiJ6AEIJE+siW1LejZ
JIjp8TLg+fRjGhC8tf3x3pQZNjU94Kn0hvZuXmRLUJK6iVZgSXm8N4Wn/Txt83V+
EWYH7PvUht8sES0cnr4Z5R/DegCdXMDwpEVMHGgdvnnLbWVpiSKKT5ajA3kTpoEx
yniUi3y/b1bSYDjgttcxeOTYAWx5FdYl8P4wrMSzjXJ/0PKGUWrFDHDFncgPFj9S
waCR5pnPloKp0X8gh+6fr3LpwhyjUwTpzEaeYDXf+GcqBZGq7SLDDtTBfv4Kv/4Z
1IUjPJtqOMke2m1x6C21521o9Df26zZ+lBhep218sBrGhmcDK1PtZjb/+nIA9bMD
HKTDX6wJKSqPePhcbB3j3cDCDggXVSuPESQFvhk4LP7m/ofZiBsYr4kfPzj6x3eI
m4nAQ7hZwaoh4zrMavs9m7Mt8A9kWwmtZt4OU7mIatlWRhocRFNc/pB8KL4PYfXq
r9Z95LJCUQG04VZDmmFePA3DiSZPTjujJl6PfLwp3KeKRhT9As5eDRqesodWV4rd
9Gek9MZEYv2BsGFeKUM8HAljz28bWM15UL7FZijcHG6DXHf2QCQ/cW2eYMHaS1cn
K27nVxNA//e57db7U3DKVQEJVBDOxVF0nXBlSCFFQliz4VonKQ6VKyjcUo20ttaI
n9/+MZG0/5uOtGThuahZkJamaBFN9jeaGsxCbV7XU0yOnBMgVRaB1K1QDWWYRAGW
NDloMqKG7UPd60Hk+U0LcU2cCIZ4pGu0rzFIcZHEE+pqVsW3sE6MFP3h+mCyX+Z1
hChmqFJflJV5nQLeD47OQjGT4ZKTX8PfIeABXGGEQn2PW64bHI75dwAxRXm1Yno5
k3BKA9G1WbJqRkKh64T8d0mr5sZz3PL8CZIpl3ifBb4Pc+T/04Wgs9tOO3vsmG0M
CKaeAqRjQTUsqWUlKtOjMnj/rW4Mt0tSaGmnwAvObio334mv2tN6qrYuCR+ClRh/
IvN9dse6xXjrpFJ0s/ukik83vO1rzr2WQ6WCqCWhelQYdsEUUq+lkxE5nY6zApZo
zREdXDYY0K8IlttlRAeHdpX0h5TTWHoSrdTF5uTH1IhnSKH6tjye4ypy0LMRGxiS
2/tTSEJ95++ZxNZDXE+Ka8/L1VSEZZoWn7dF97fA2JHfzXDTaPIoTooHKuuU7O4v
Nqtum0yn6kaeWrdUX+w7GVUNVqhUBoK6JLGdv90rygIVSXXCwUWL8aJsDYA3GiYj
MF+IFUlO1n2jl9sl0g0aqotJ7bRGJBqO6vFBmu8WPXEzN1gBKXnMwSq7xekV8e41
GHqZ32sxnFq7k3GSKLyT8lJ7I6OKDjCxIMxBcJzpsoS/l11uQyBc99SZ9m5CgMxL
L4c9M3/fZC8dVceOWFgo/pL+Zg1aYzCcBfrqvJPofM0RB+nUuj6QFvxh1/tBxTnu
CnyWMDCdmlWI71yoNuP5EcrvK+trP1z5PdZ69Q7b2orDu7E/r2+hs5+WxtLkrVLl
8C/4zOH2F4X7CiEqMvKFpXB84K8bIWgxTJs8Ivp0wqjrKx9livLbIWiO4xJA9z5q
UYBpBBX/q6HUGpFLFpZieryndYKGuGwSoJkvBOsJLNbu6JvBy/WQb//0eBZUbZOI
PP0Sp9l+hAZwsHo40zIEFqEMYeZJAkHz/4N7bEqHTn7S2IdF3jDMxKjx+GQ/G8Li
q6zA8hvUkxgvAnK4z/Q7HBZ2tw383GMulEDY3deuERp1NvD9kGXTDfunHhVBYeGb
aHKPofaWY2gOhG4I9wV8OSlzYr4qon6v0LD6BlTBSBIV7Fw3VuovdfZZpxO8q6EY
Ca1JRh8s6m6oE51Q6JsadfVCN2hQMT9C/gASrRcN6GCBDJA3k3UQiuQFxo9Afx09
ZxIOlKXAyBsmr7KzUE25tGn7cWe67mtGrsYQYu8gi/95IyAzTyPb83E2vXYefsws
62AuwdFVaGDga3B1t2PIKcqjwtSE23s/ax328VFA3MZaYKKoIy9D87ymUOwbCWwM
q6w9yAA3k8j0nq6bzcuwqCGOHqd6PmdMgJlpehnc9bU7TKqBzC9SPlnuwlj9hKjl
hR56WxO112+nvgxzCKVxvpQ463VfMRTA55o0HV2FWOQdTk0WA+9nz+efoRoroud1
emph5HQ5OcW7wcQn+JUdovHFtzCXTZTS1/p5qn1cZDUa2k9/w7cGAEFE6qbNwiki
lq7IizY3obz3xLmpf4dJKGiCx9P1qe+F2lQQBLQ60aXwit9ZwrdSz9e2hVa8MQyd
82kbOSOqZzIPNGBjbY1C5DmNTu4HBCvx7ENAhJfm7Tt+KBi9Hgl1CI2mWBsXlfFS
U6JQbQeLMVtWGFMne9uqZB1ZUBEQrLKZn/xT5+f82nQlL++fqkdVghIXVviGHWms
NGOnFpRWuNXGlMZDV5ezO1eOd/boD6YOxx+L98dXHfelQ3RX7trIrVlagyz0r0Bh
Hcx53y73XEPQhwV7zam7mQDYrqM+MNKfQUU6Q8OfE/BBAZeO7o5vXNTynKm5KTOq
8XmKB19QpCrRaZQ6UFMWwc6kZIDKoC4wuTbInE3ej1FtrjhpyejeR4SpNKdqyP3i
ScWETHxt3yCNKtFRrs/9wWbTIYpDaGE6FUEsL0EiL1HB3YP+EpUxMDM4nnB+C0dE
Uly+GqqRCB7q8KIOmqdRbpckFdde/Vd+Oc3RM0/hHGj0y0xl8J5ByRYYaabLK04A
zjeILJPNRLv+b0IGo8ggKNzjsCkDJb/tBHJ8RmkwpBCfgcTeM6Y54S5/aSrbZX7z
gclxZd1yoYQDe79Zj1dMzuvZNg1cvSc9MzPUwn6y0aeh17OMr6q1gsf/pIQi8ftg
zzjMKcY867UlR4hCwG7QfSjME4G/E7q36ndHNjnXnTm0h7QZ/6goH5GptA3oJJzl
op3i7efN19EPDiG0kQvbSladM19oy8ySMqnlp49uWDF91zwIeI5ukY/T5sbZ3tkD
XthlqEjpXQHoZFjYMS6Y5ooueEbEhrdWWBHsV5KNngs6Wusw9sdREht/2jP4+Gsx
M2jAZZzgOS0lvxrjMPiQoDQEJz7nq+zLH3/2sgcEWLQbHq0KlAc4/jJaDctSqTfc
CMsYt/BiIUjJDGAmpQb6IQe6q7/IgVfFLXWwzU9vxgJmvVo28XDQ5uenR5Gl5n3P
y8I7GOpFb0t/V1tRd9mudenbG/H7u//HpwRHhJLznRThTg+iedDh2Wqzluka9+ZK
gWTN0mpUUwAr4dRxvK0F4ET4OOkuKNg4R0/JGwL6vhtbsJLF4nbpE0loFfw3nB19
bdigXkgzgeg1ngDMJsVTJXVGUmKr4pTkPMvKUVxwlYVgpkes5zRxErVpu+l1WeIQ
R+/mkhUiQmcMOyJhIjsHX9QWQaYJvxfgx0JVBb3Zxl8B7ZNkSrIINNBQdEU5r73X
hYkanbc3VtEWJumVycA6p7G0xi5c0LSfSH4QVL63yASdKu3f2oUh8fJKcuE8V0ED
5kKmmyY2BtccU4tyNEj0Xzdc/EpRt30cNBZH4m4Fm8q/4tLlOhb5st5y9NE9bhoq
Asp6Zl2HoPweKXXosYGQoLMPMv5X13phON6eT4S+mjW/ImhGldyWnU2sKK2+wznL
S2/RbL8Bs/33SKK1Bb+BA5wNGsCL1FQAC9qVNFQfzs9XE7oJN7T/UqpI4N5QPqvX
VzRkYB2ppwzK5oF4v6NcTHGJ6nwKecBELq6eHZ10QcsqfSeLrV8j4/WrddwJAAE/
4FwT4+e+/VpDqw+zal65mGpDLaTRp6FbfYxdoSVLgzlHQZBUpZUXjAPWPLM//USV
kTL98cuhxyKLTlmVxEOfacMqlCoGJQE/Il8v48KAr/3Oz6JzskM0OidVUAT2aZ0T
LhVo5u7DQjgCR+NL0u9bcCgfVG50olPr2q+lec86lqXon8+PKeTIKVobqlrKxGVZ
tLyRzQMQ9UXVml68ur0ld28rjze4WGqW23+fwerIwRsLp4b4JFDcvpj3EGLp7xTm
RKh7XahhYvdP8DrJPL5uVYMUGkftd/SOkBCLzdFvS1xyWE4kSfAO+27ZRqTqzw/3
H6GBz3sAtk2WwAGHsvmMMTvQKditzDx1O7BvgTnUFfc8F/5iqx6QgfEEWaazt8tI
`protect end_protected