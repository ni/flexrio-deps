`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4368 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
akBpHK9XojjdOyFTP3pOwpjY7YH1jjjkBYghEISQ8ElD6OhGEaCwUyq2fWSViGnz
liaSVoHzMIZHyGBB2IXbJWZR+EfuRXLqgtlRKbJzwqr/6Iq4YK4Cwf8AnH2UIsmm
3c5hihLsgzYjA6l+ec1p2zbAVuEpOyAMREgXim8X1lOVVirPnKVDXb7grghDj+GX
54nJHSNrsCIgqoGhLzq1enQftcxm7QeyH+R3aBWdC5KdA7sHKeClOPolyCnRkUjG
alGo2SSatsyV6VW6mPggPpomb9qZZ4J/Y0ftgiXD9qJprvr9SP3ki7fpOIsbZvLO
Wm6n+qgzZihNX9gBSGSDP+fyPI5f8nKPULsMdvHLeVz2WNLCGNC4fp3igofb+pf6
XYGgL4cUojLo2ZVV+39682WhkY9H330Ny+zq6pgxGU3N2LVTm2c24WxBU0+qBZ6T
KLnlOvww48SzwvVLfaF/SjVxYMMRQRiht+Qf1mpjq19u1ayDI/QEj0xrj+y/MNQe
qfWTipBRHqxHICsvCtM2n13Mv0pq46r+a4ljCJBYCjFru5h6P4uaNnyvXmSzzDM2
uykMx1PGDtq7bYV81OW/hz7o9kY63A4o4Lqr59FjiM/+0JSQTF+XXyTtke+KWw3i
Bg0lAtsQVc4rVDBLukk6/K29b4t7f8e7KlTicrXmrZYBDlj5MMfZEgfDXqHFTbVt
6MDGZhDFQK4hWEDDBPQObmrYz5Pi+HZz/Y5BicM7M1MAw23B96FGUu/IMINwncey
hCDFgjSf+kggopiGXGu03al+PDgyCT2ksHSwSti4Kvmd7OO0c+7vFhn400ECs6Kp
P2iIArBhmCW3JtQG/+ZrYx4rVtWzMs713e/Q+vVPCE7h7uuG3cAovGk1mXN/Obzx
9fEveM0E6XOhCrlpSRlV+b901TyOSKBmi1x2v41c5O/KcQp5fK7Tzf3B8XBcIkuP
NZS4Dfa4AzlRHX86UBERFEM+KraspfdYbP1MXc25GIPxQoQErpxYUkELYsFyKZiS
KIdgsQtj0jRV5dJmzACLb2Flm1uxPJ4n3M7UuCcQuHU4Tm0svWFWCA4xMlmkJrkp
K2rVxdh1E91tKMNL7iZXW4CHIYqSSb/jTfSDz5uusUaSxGNP5esRFZD2eEeNALAF
h5cmuFU+fz7dqYXIXnQziwh6qm+VR4Y9BbrcX9JT+iI4PlsNCOAiEfwZrw05QXKN
KDJtMateIlwoB4kKNomQ8KZKYfcuDXgQlYt1wfyLUtXXAWrosZX3ph6aRcqNetHD
Ys1GNiNb9jJyEaYeDu52F52Z4kQadLASabdbJn5Dgzc1qfWY16OEAjVYW2QCIHrO
Pmqmu4vydCrIZBV77b1k1H6wXPkAOxGdLUKVxj0j2or3CpGNJXNjpVrlwySiFsZk
6G2HZyM6qsGK1HfyIStKKamI5DMju+0XMa+SBxz1VL0jDvDNrpx4G5aiMWkdQTeW
7tPlDEAa7c/LKD2bKxdwgtqbSu6IvXPjDbiiLYKTTQ07t1GwPgWZbX/V4WR6AdKy
NYsEqfRzq/zV+BrAAo4MrD/eu6kdcej/nlWp/TNHaq0+fjm7cLlGk3VGG7yzJqvj
pqN4V4d8mvcr1t+ex31hwDCs43Hg8S07Gy9rLM1eX0wlJgvo5lGTf/x7mEa6P5LN
lptM8gqbITQDT6bpAQFnJ8WvNmAO173I3umNqRu053AIE6Wty074cJ38KJ72DnVg
Yh6zgErkk0YQmgjJO8pfB9Yn9uDni494VVAkbHBB2E+0fqiuA/P+5DNxRBNcAM9B
H47i8NdEXvUEDKQL90+uq8jp4wiih0HgYB693YWLi77uherkCR+GGu4VYX5zwdg1
+OwmoWCdFcctK/dY84aUEFcgfurEkeB3b/DgkwZkKf9YPm1I88hqeBziYgEq9+qv
4cHnlmQjgC5Q7gYlgJ6SW69T298UXdAqQ2j4npJH0va527FKQkxc5RV8yMYEme+j
oaXAsO5ZUZ9BEdqXOjCeil8Kz40F2Dne64WenZqnUngmErz1533ZureC3RFu5nXI
lnudOiC9jPgUW03KxElFjwkRWFHyzSh0b2dR2VXKFgNO4kWLpf7cteNHVDS5dfCM
Hiwe0bauMaYt7QGIcgrzVtpo5IFfCgrqPcI/wqFethtR5BR/KjPvglw03aYOxS27
5EuPL8tKuem+yV4E+wEyNzaKXaDHufV7/cHHZtydUohAbcoGPP3nJGFAfB/Uoi80
dzxFaSIcwhW2j7NdOlDpwuDSh8BKAHcJLbOvgHXe57ioYgZYFRlcMzCLwaXJ5F3o
OnJCByptNVC9Y6bTi4ELSPqLUjNNNMw4fsqanRWNVh3ilG+jxJvjjCTIJYnU3EZr
KtCKdfICrfadwGRv3sEKB0Ib80HTGTY23dcrAhTNucE08jlyuFgCkpgb02MDKjE+
9QVEoZCiZ3jDw/d+YMxPS463ng6YOlQG6EPteICqAvinYFgIalKnOqXYMzvUDA1q
NZO1RjXylIIeB9HlKCcyIX4j4Npj6i4U0iG1w+dNcgk5RjsIoQaS3rE6XzzKjfII
550mR6BQOGYN6BEY4T9oQVdLpyh0DMAHWmmL6/KKrqvMvuqb1/48qkuhTAct1R9g
bM3YfVCpSlPnvBoeeZUkNLk+o61tWohG+G/J6F60T0GSDzx9jUVQDlawJs+FVZXR
BpQq3paj18Or7gowXk6yqbwfJFprxHYQ2GUQvs1G9xca9FdCLQFEdRJGMvwea2uu
Wee7cig744ROLbvPWe3XcgjXQMw2Udol6FyCvqCXligzuSw9beD7yr3bu5w1v6bG
u8PK1IVulJKo5zNlQ0UdsPD5pVYTndyTgOxOTrKT8ZdJhjCGjHIXq9EXMhPOA2oh
nIgVUSmUlpQFGeQgHaKoUS9qxSTyj4ihX0Ph8t4D2BZUz5FaLpVRsMgTDjdgZHWz
FU4EvF1PzmufT/mi4f60XHgwpgZGUYgRr/Za9pfO1v+4E3T0JqGqS4WVOF6J0WRV
dNUK/hp5QODSX/9MIHyNzeaEFs1+F1okufOzG5bdTz2nS4CT07RWUl1vzd8HtDLg
ByxHNHh4I0P5IKZTPquQh4EyojYCwDZ6ISsoIivsQnRJoLGf3UzzOHWjJ+jb70FK
lGNGPuCncegc5HM/NQFdZLyF4AiQxUfLnrZKaAN7J3ssw6Bk8bhaxrSRD3kM4FAg
jjmjb52WvtXRWiIj4pwAZSQ9caPjugISF2C7Lavg1eRcXHJi6Y62k4dmLFa8+L/m
0Sy34x0NZylzP8w96HlR5IL/rl2Z69zJ3HwavCIcN5BrrXSPdJiE8Cu+XjYd9nA5
EyeJ7zY9lo4fBBN9rVAkfr45pkOxAxCPEZte1678U/Uotn1+KkUZ7Pm5daQ+QBIZ
FtC7Y4Jp61jjC9ludNI4Ni2CzZiFUA9dmMNunUG4JEHMIKDrgbR4jBY/wAfAa42u
0JVE66Pl5nBhYnvuA+yHAGN8OrzDek6BElrTfTOuUnW7aFCdO9uQgShgbBpFQNr1
RWGRyaWR4YwYuuAAJRhJoXuywxfY/+H/F2k/0ni6jglE3Bpte7ADx0CIxGmF+oIk
Lt4Zh55ng0XBUoXx31+5/ZqcLfXp93+9MXJgY9CY46naUmZbsakjirr0FbNltVnX
sBhUxtY2wKw26BvY/fEGC0MR8Pza0B0LDUDadTOyuwu3OeT+A6GCxNMtXvD0NTJz
SRVQc6qipAQAySqvfsIHLb26rYxWMKkepfHq1tdboPdppcL+gKieMteOsj1Z/TXM
z9qorp0BphLO11FbLLNVi6jzqPHYCpvmeviqDQ4oaZmIdvLAHwykRsU+uhD4xj6H
4xQafU5rNi1hcnPldsZT16St5NJN+0hPJ2BLGKvX0eeFaraLgHBuY4gdrHIMAvDl
VIq/wtbPrQI5CbbsrPKTIFw03lssCOf56aj1heX8x/+NPkv3mwvkanCH/vPnO6lC
YI6JD4x2TLjo3/zVZgVXOCQJP5wfnHT4++cJaD2DqB7HQWa26o2RoEpzytPXT/0e
sgSQcmP79PGJJZlkHl34uV+bAcoz6gv/mAYzRN4kJFsgGWsriT9Am5LEao7ia4HD
ZaWSF0yWlQR4ZpuhKYO3eJNv8DkQTGhgl02koQYpYH+VdHg5Eunboe4E7tSzKosI
P48bPs6DBFq3ymGEVIM2OqHClRtDMWAAQP4qMy9ZSMjeKZwy5OPw9TLQeFWWCKti
R7vWv2NjEZmGyCCd9Rc2qVX0ddVsZBWLa1Gl1FAIcEOB5L8bupLOp1Er0HT0+Kz2
SJDMIVRE529SOIK6yNc8EOxMRfS6A+Z4adA1E9iu7dFq+9Q3xEN/PxYTbUPpgm+p
ElCXR3cA4UMHHNveGkRnFfP1vilPxLSq/kDlQsjXLxfYwbN3tvDyTWQB1oxl3G0I
145gFE3nOs1936XjvgzIO3+zFp26uErQDK4xKfFHxRcshUjyzXSoPt8QHRAGVFsd
Z/r61Tc64RHpSZ0jmvTXgvpxbq6wvEIEAJRD0Z2IysoR6W0L2Ja5JoGbqjPZC1st
L5On49R1UDaQasGFcpuqKF8dezX6El2T80M6CA+euglJXSjhmcV/3SvVPJ715SyP
xrFT0nGdiN3/1oaqoh+CPPAUrU906rbswvll7NUdF0um+0TG/vBnFWLunvZOH6rP
Ohkj1/49rmjYgvD+UVtESMe/g2gdH1gk0fnEP/4iey8q3IoLxd9mwbZ8WDknWZG8
8sMDcjMRt+q5Ve5gOsUEf0P9yvLqYsnphOqC8pLAOxWUFy6QU765XTHd8phrbfJ5
EIfPuw0osnvsozDqdkprxp//ijZOggmU4+0sxddNpI+nDQQLN21VSBbrVAY7DkSN
26RtXlCeJi+6Y9P25n9TOGVqSgteB170x9a/v6DJ0bJaPf9jHY+MtBve8+fFPBDk
5a0QkB1Jl8JJNa7RAv3LjgzNenImsZInRu4va1jaJti1pQlowRLrACcSzKYxdIoo
3ztIz7U29R9Z2ZWurw0BrEeT2qV9v/yz95GtbKJVl1uACCWZ5fxS9eTJqlOkGVn/
mzkY/FoOlIQ5KXNO2fXyFNItCK3SVhyTFLVhmPXjruCCoCjwH0AKYQtHhVfRn41/
kJwXMWlXTU21fIfStK/206rUyuqDGTFzsnYI9Cf9c35jcZPy5mqhdQT41K1Tg4nk
3mzz6NaYewb1zEIHw29clJfdikgcbIt8f8Hx5qPF0mO8WnLRvN490LAAPkIeqOX9
JC7i7yqnDgILPYsCGXPxP5+xm6/hNlcqnkSD8DvKOna3KwrIFHHAaQriEU+0pJ5H
7idexhMMmW1FghqIC3mfrvlCE+6Pv+hPBJTfIS6fS3Km4vG56GXOjt1RwResZKbb
UKMx1si66Eek4cMYFZy4pYV9IKp/eLgYA+7f1WKsbm19DFqT9hRLTzYD1fn6Ralj
aUie3eMHjijPlRkEUR5SQy7Q9rpzii4P1GsQJu2x22HAtIiwWqbYwZO5dPbXztIR
+Mfhgr6qOqBMB9ue6LpAgrGy/AlYCR4oDg89QHrCSY5idSn0r6QBezlpLxu4AL2t
I6c+pZ00BoNsytKMoGwchAbG7LE+dqFDjVjB+cLp6mhJcmj21BPh0+YXqlEGKK+A
W3EXAW7GzEcEIz4+mPCjSZMjXs4mBIC29EcLCtsSZ68tcywLAIw1yu9onPX9XeX8
`protect end_protected