`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2128 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
2n+M/KhW/CoPvt8soGKLVmd3tYsw3c2bNhYvAFbDiUYUoIwxXtL2vYt60VV8XL0a
GttlpnOclQTVbnSSnMT20pKuiiOafdxiK6epp6rO2wCZ2yGisK35Y1O1dveX6kLL
2v97AhshsWYf65EIQTvyCob+feMCX3/NJg4guuleTuFLVibHyewwjb45VfUJJefI
FegSaAOUZkepScci+D9b25wJqgEtd27Txz9xE9yt29moZ/RUA0rhDQNsoQmoQ79d
jhdjnIT3rlLcaaBn/Hi7PvNnQ4dHSRM6boLoF+sygfGPz3BkxsQq2P2fhgKxTXdz
UKfydab7lWtX7j/5Kto0uLJRalbtSDSmWal0H9e1hm6Xlo4zxxiDVeIienkDzTKt
Qp6QHjNttYsNS710YeFvbY+Vusvzg1xGpEjtsboDfuWRAIRDF8Y9H3lqe2o1viWT
hipoX+SHX8AlqhbSHmwuB59vMQ+zbsi5NLnNb3D9hTpSgbrcU4f6NjYvdNc/NgoF
gkQ/Z4MKzlh+6KySnnFviamFJAYHImVzUrOFabSrBk83oxTzKoFjDrMKEew3UM9b
z+r/BpSXpdoHZTs1XaNeBDMtise6nfDaWBKRH+2ARDFgnxeIzGwYu/EqOWhhJS0c
Yb9AsOv0bwNAbxkKvHQ3koqDfFsmDSldiHs6cR7NlNfpKkKtZqUxoMGMv4sv+AQ4
5u0iqBHDSosjo6VoTgJwQZ42NHFURluCIhbZSngI5/RpEVJAPL2fzCcrZIPs/O43
9Oe3PLBeNzfppdfhobRqiKRBE7orRteMA1uRTg4SJ60YS0OlrifC6X/qV+LGCJgg
OmAluAfy1QARkboKxbm0ttbo1zJEw75wa5jwdVdUFnk5uBwmnx3DjbmVGoP3l0mZ
cjsq4pRpAF7ahdClv5zybEeP+pXYfNRQm5hS17TEZwnPzobCwO+QxfGIU9T+iaiy
sNHkKI6uddGcgJL2CCwRE2Wd9vPKCOIzSx5qOAA+BM5kFL4vy1S+Ei/lP0fXHiSw
endzoZR6f0yZJ4KFyG9bZt/Hx2G7QXqA0tUj+sKwnJIMOZaeOfat150SNC97Ev+W
p23KHur2fKOAkijmpFf2G/zNYIRxap4R1AkAxn1acV0rTqDmj97mH5VfninGJwWf
9YP4/MWx9Fm/Kff28xQfNKbeyU9Of3ZOAmlz9fkmt8GRJHt8CL/FCqGJf9WC9/69
AL8vI9LbcwqHAZEkXi866qR6vogXa6hGCXRL4F9FO22KVCPWCky9ZDHpn6whbIg2
17dq3IEg/uGpuKFEy5V77TYc9lFw+UNBLxkB/YgnCo0SkOBV0KScMvKuo3e2p2//
NuWJfcCLiIPxfu/3dtGCWn3bsrkz/RMofbab/tiDrdcVECv5iumvzlaqfql8gpyM
hIOtsZrSBMNDtT8MKmUVIYEvIjM1is31QR+775HUVWs7TnHbaJrjDGh37NWtj9lQ
JMefo1TWWkkUKIzs6VNCc1T4UDNa/aHKHGgKiWN/UogTfiJLrnGGAuTVZXubhbSY
mxJHvc0O3qztZOjUhoPIY/4giokgLWz732Mgy4uu1ty9PyAlLoLq5ErMCqHJhMt1
utFa5Ab/NttG5pSkJFO1PtbGo2Ru4uTR5u3suBQqdgyyFqjGJx5FHSRFwf0iAnYx
+Ib1DU30KLhg/WnL3/FXGIBwDrPXNErUg8hN/tTveRItIlH+v0g7k6NFE4n7cRbW
jkgMOxD7r6LRNmaQIl9n3Dy3rZlSgCzgV5TwLo72FBTa0ABLXACm1GBM2ISgEClR
5r1hNnEJA6VThEHOKkBXrTF7MPjU1fRymMORXmIcidDHBhpFS90LEt53QdTqWo4L
LGYudZNLdk2qxQK4it9dnua+OhpjBRPyOTDIq94hNElhSkeDvKLx6T31uuVwsEAi
m6mLQrI4nU4veTVbnVXDFfoQIaG6VyMnwtqWjMSxMddV/CeXBnL5Q60G8ifIMm5Q
WznOTLm69KGTz76ely/O62qPKv1zbgf3dv/iUbIR7fD2bIXvGZ/7ibeC/c5MIJrR
TCsnPetnEcof61N9kN28wM/px+EG05m6z+Yb07jyVOtbyL65XOMY4hwF0N5b2xkA
yp55Aqh2cYcgchM6WXwHNd9i4H/G09V8nluR3A9Zkgvb8ebr10p0BbC+0phsdU8s
5s61kYOSty8wdP/w0td8DUKSOnRTPCPDgI4o7dSxMgl7/HT8lAT2v+QypgZwoxKA
iucgMiH1ReCvNcW3XCU/yaAseV7973epW5s6rAdUPfHfLlr6Lwk2SxNo+EDeWsiB
jcqBm2bAbiVQ5Jfa6Rb/QSTK4ZER9stqmYa9HF1ZQ0VSUzP7BjpQtRD3O0H1OWAS
49yZIxziJ5pkEN496qoe7yJEkCYqg1JX3/A86yC/sVinIC7tZM3PM9zPjl+vycPU
mx+NNorkULo46SYAlaArUDF1OIYg8pP1gk7TODsJ4qaXEO/gPv/nDhc+1h6aWTIt
GcAphBfYTebTg1mVSEgj6XWt6zePbS7mX98vLlP52FXZQREqfI3k3dbf6I9c9zL7
JKvbPFhoTTZpUBAxT0H/KEbn8GCBr+VTBMTlCrjL4b58SBS9O2NL2oFQE91OPRKB
14F7jJeyvKFItsKBncuodGlWD3bPWj2C+X6s37Mnh8CzsLQuaA8jilIsAKSsTBl6
VIaiGT8ivDV9z+4sw9LuGQ==
`protect end_protected