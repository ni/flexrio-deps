`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7152 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JXz1+zHgF4n2s6TEZD4KtuQ
ATkS0e5WlIVeyjNZ91Ns36sZQfrQ9R4SbnYvAtVIyXSebV8YuzTAxVu5cSEQTk61
5n2r5/JhhTkuVyXS/x9FWMaYUuX0r6c5fOIIpcYX/N2Il+0Kfi+w78MoFgt+jC+g
Y+B8G+/LYC7PboHsDcQKNQwAEHPexPG5fMomsxrgSINO7D6yb3aIpDYx2ZJLCVKf
5167YFW+t07c2OUezhPKRx//lZW7IHnRHo396Qfz9y8Egad1OyDICc2zzeIewYH1
l2cK+jPjd4++s1T/IWLG2bo08NqzgjrDPwK7K5D0/iECv0gGclRBL/p6nk9fiLPO
N8v1ruFupVpkunNwuuqsYFKMy/w3hvCa5x9obH/BcuQSA0+k0IVje2xkxJ5fpMLi
ZA29lGACuqSANOY9jD6YFBDZZyKurjxZlaOf+B4BLDd8b0FW1l+bFUPtEnFP3+6V
Ys8u738/NfIWZxcdoM9qVWyZ+iM8SVveRbvB28ukKdBLeJR+mJ7etNQBL+GRYwPy
/UAcPV2a4JB6wGMe6NHzZnxOIzHf2WYLBZTLrt9xGbZrrBWYOoRqJn8fT/KhkZN8
ApEYWzdAiVNBFunf6xZJoMOfmUlFKSLhWmeKnw+EDRFPCuPb17WMxNr6DA54lPl+
cRP83Tofyj0PVJ9yJGxUPbnQ2urj1lGaIn+3+Q/YOf44wFCv5xoz32MvjgF+Od0q
sKxjjg8z5LDm3Na4U5TkmiJCAPN7QekpQn4xiJVLb1SthL9zaA9G6emYzQli++BR
B7j78bVzOIQ+GcIwHVaxQfp1fnmSZgsI12eaJePZMSZx8KlixaT292VZ3jpWaQrq
Q12bXKUu2Dry47DZowVl+WipKoSBtvrS67w3POE+Ql80RnXcgr3oog/Q6vXVIawu
Yw9mmzZKRrYT7ZFAPwyO/681cYvBqfuGLqPaKitrMfQZQEeBx6OKUpzqgFwgVSiA
aq9TUD/5RU668Bb0i4znLRDVdIMGpLVC/UxlcVBxlIhQkPzhaQ4rfrNoc6mgzqgg
1Rhf4stA4bGGIL3eDJg7daCjxbU7Pjx4DZjO3HFs/NskpMkeQyTcsESrOjOxlPaf
ebOXpGi/+HjdEVYQxKnIi0YtJocCKSA2qLgZ5Q7YeW+u+NmJYCgnVutOibBq/J1M
zLZ+0iyZKdLL33lPahahzt+gfmrfq8aFYJsMKLDtNFTEuOvYsbJvnz1nsxb1DNuQ
+Ukg7D5Psln++/soe9FfIidqTSmB67VcqZrtoz0+z9unE7LI6odaB75+VT48pzN9
LOeNXBTRiNtmO1IRssdk6xrrirt36A9/4sMv3IJWSzvpw1Dz6AbpfOmsDg29ZQN1
mCmTOb+hUKQlxi3+u0gVe/w93WvSSdqH09DyuAlBUwhptXAkUCaqESrqZeA9/XAf
sTvIiMBqlmAR6KxZgkK9JEGh52RVQdVuY1t00drPysBa1eIpdLjqJUKIvWZq+WZw
KJY/aY6I1FtUGKF06p1LztLXZzOXS/7PtjWPixWdiA90rOViMJd9rTIEBGGKIaQO
HYV3ayAoK2QNudHwsA31qD0sw3NEwmEUMr4bQtGnCM6V1e3rbDWzT22d9OrDVEkj
XADHm89xox1j5uu3BuR8+kpYqIgehTu9D/lc8U7Gi+py47sCgPCS7Xe1MxUJfxyY
y6GPWZ/6IvE9Hic1ptJu01zcOMVpE9Kf1ioiNHCBZBn3idReqKC5Ur47MTFyYP1Y
1bpH1aoOXhWbf+P/wn55yMu7ex28mNYSWOcpmHuND89DYTqf71YyfUa9DsuOMiZs
zuh53KPzBnYPv7y4mBtLiaS5AA87D3kHcrFQD6BnOKCGKQm5FPV404tGdK9s8iAe
9s/uAmKKd5U1tV59SbU+bESWcgMz384UYKJ/UkSwnJ+YpVn3KBd91UkE+uRqBQh2
PGBpZLm+zgcNrq+U86SfxDnLNVpAQPspINdyvMrWhDMTIOLzhfgc7h/wi+g+Rd+A
daWIcFffZtlLyIfUQatEaZxm72eiePbSpCf6v/DiIZY4h22acmchn4L3F4b/QLf6
jq5Z6DcXmYHz3xG4k70oouaC4OVHBUPSxcdphxtFQ/1y1zVT6LhiAluSTEQSbbK7
n6LCO+RE/2xshjE/VPKlk4jWqFZeb9jqOs8B9Tyb/BLjPuXwKRM1StjRFPKT9RH2
naLZmd9eX8paP2I0jT6t5JOSMZ2nOQbO4zOvPWAtdNSegsEhP8gt90Sd9GLo+4jN
xNXTWK8HgM2x88LzKWN4gZdO76eAAxQZPKr2TkTTV/lFRjyHtkgUDGmei7IDTyO+
RlkfzoIbw2xqvyICKVi/AaVFifbp8gQRVay2gt+pCVEnQ9z/qvyW27rKUvNetVIe
kPLb2taMkerNMuCCip6zo8D4a5Ek5idB1sjaaFT3VHsCjViWWIkaIfJlBz5UbpLT
MNh8EXYaXpb1OQgOxuRVKVl/t3Db8iSI5mNd2pIYOqNiayFp1nYiQPkHQVorKT75
8ZSSmeZfgQGF7AVb5QinrjZBZiz99Pud8AgUomguvX+nNplJg+AynlH2VGjvFY51
86nkcnyunEaM/GkseofVow0oW/Visi0mr+QkDLY/npm5asVZyK/yTWfgu1dFPKIv
Jvn5OMfQ2MeSqZxUsv3GTB1RBv7sEsB8dKTYEbEPFwlVpTse//0YIl6m1qoXcfwW
//wp88HtPYCKGWqHXChZcBUAA5Y71b9J9cIzcNF+D2Rh75jR8JvFYshoLmzb/ARH
EaZ4GqiurttOt1cdjsMSr5i/ov3MHYQ+le4z5ySc0fpTBdvWPXKHZnWwmgNHpvfu
ryKPfwIzP8QMeNrqrpR1AwdIMzlK9n+wVhHiiOYcWIfLU2wGt7OIdIGzP3rmGoM7
7BO8Hc1jmDLhzVt1aQKDe2j0PM4Mg4VWMlHlmIZkJg9WK4TsdShQIVXEPE6PO+sQ
nUysLpGkokTo4nD/ppES6MI9wcBqKk4E1IHbtoPkSERUhYIKEb503M9Trn9o4CHi
KzHn+DYu4DL9k2D7RR77IKVC2B0gNsoBF/kgPxDDoesokSIJFEt1ws1t5qAFwzgf
/606xlwuaLDyrm8j7NOHyzDVfhQ4HP1Oux97zzaMIhti5ssvveh6riYMVqQj0B4p
UtbpnqNUQXOQWMrfYw789kCcLWzqOilauSzaQMDKXiFNHwvnXQ4myjhfnDZ1yWi7
bQxpuo/R7YvNlJ1XE+MKfYqYGqAn4RcJ8G6OKS2idaL3cLWkCE1GuhrneR/9U/Ux
WRhreQYazHboExaH74m9+jS+slSNeAhWthPj9PVvTIHCbkHJMScTDHsGVkhLCgjV
mLO2sK/RViLfdBE57jrLzVQOD1EoU3n0M9EvSnoG4Cb/EWrDCHJH+3a3eRHui0Od
jmySqswAn/maawhqobm2sIYlRVbx04TzzfK3cszMIHHv3TDGHYmEzXVIQtp6uX02
MLeAIDo49eTGZMLlK1qPb5JISpf7jZkGCqznJJyFMXZoZWYVFqE/j7x4f2lqCbbI
pVlwUmvckm7cJ4T8wI2MXfq+F9iNvnLI+5F9hFDEqx3le8JgMfNAirvzFIZrHtkl
Mq/Lwd3ourwXsSpfdnOktoybQ1hjYO5jdiMmK/4gnEUfgQgPKxG0aOr9zSD8F/VU
x/7nXkv5fkEu7SMYtyS33rO/fTbj1rZn3xp6YpANYrVRcGOGoUO0rEPPRp+/rFLu
p36OG0wbRVsCIJY9C8NAKOp92DSOWWbz+lDGeFQcwQE5tYLHditJ4T2iKlfxe4b9
UR0Uz8sjmm8lPhp6GzpDNI6jxOPxzz0FZBvrS2PCmzPyBPuCCNfTwqStKwfu/EZ/
PegEtqkm6cmE0jSJ1DNA7hG3VMBhKi1eLL/QVKslqKnDNmF751oERGuDglHDgYZJ
gt2lS1c8et7jkx8nLob7RnhE/Kp/e5rBdwcxvyAayddPYKM+sT3GSa1d2427AhEs
PJR4jD9pAbYXFundLze7efS1GyhkNmnykuA1LFMGVOkaed2ScePCAgHj2g79sYDS
y7yvKXGNqP0wrO80nE2lNTvTqShZleOFYAao7xSE1Y1eZbXxgzRUB6grISB953Cl
kfEOxP/XJpK2SfCvirps+hlwqBbxHCyP6/5x++yoMdY4VIZzBdlgPYv0al5KFT6M
q9zISv+n1y04MXSHQhSOKMTPnruveGWiCdT7zx5tXvnzSMYahOtcQKYxkjQWI4/u
LRsX7+pcQQGRGXqqI7Y7DX34MOX/uaLRXXaOoCa4/SkkZjjPckxgGczyXRzlDuqO
Kl48N7hRtdX95BZCih/UOCCx7f6aHC9HtbHrYaRiP3f5UNu9R7S04P9x0IXQjYbj
0adXHxTBEidee+2ldqM5AyzrQRM8MZ+AB7Pf9oytgutToUMFz1dkynZH03dHpK/5
2F+8p8EwEgEo3IMWzO05YJLLZisgvilpiVzje9/PhTKVZTgbHevqChvwsc9Rq07z
tBDWpn8pjtmF7Whzz1hT/BGEYNZjgqFj1oSfRApK+i6Hp6oPIurxmAe2YZr4hXxX
QGH/GUh9mmjcu4NlsWM/9ow6bF9Ea8HrDTYhGbgdXY1FH1hzzmYWBnIvapbzgJwB
Jwdp6wRFb8gTZT2YE7vHvz/gjbU8b3cLJv7OEuzQUZQSr3SWMwkBxZ2Wi5IfVvaH
WREP5zIyxHJUz9ekY5uO/MgpWc0OIEjmTeBZOrG3cAhhb3ocfg1kRStO3v9N4lCy
ZtszL9Jivydle8+drOuHL5yZ5nvYLwf8FfUdGqx24dPXFfJha3ZevxYzFBb7BXOS
wXNc8//3z9d/AuWOMeBf7VVWzPt72qGwl7tSsaxXwrlisQ4lIIniab7m0JaN2Pt6
6Lb8myc0vfy1qxpYN83WGNg9nEkMWicDILWzUCiBJvaYLpP7aRbHx1RfqpIiaLZx
LxugWgO+9GxdO8kNhht17qNW/kr/sV0Rdd4LouP7O38DnR9KSrfz5e0oeZgZwSoF
GJt38G8BL7NfDe70XBmR93ddUoEk/elpFIpyEUtcidARhTztQH+FIS3+URH0V9/H
R6N1DJopzBhHkm1mDjLBwZJcuPh5360mlqXv8dn5ePk3t6xP/5zw4gJvV4TWPuf8
2HKI/qE8pXZLgJlY9PIKtOy0SUH72ceuXjj82firPquhW/T26T0jYdhv5/JiGElN
fyd67bUm17FskwyIqMcMco4ILAVAbVzVxCzXXfi1NclSTeOYV/5m3+ISV1aGWQ8d
yw02ZTk4riQN+Ye71XR2fhFGmwSZ+/9TGl3W1YYVAq8qBdAzB+DlyOPlFNROkfam
UPJ7WKgaN81DPoxe+2PY0aBaikS914pFQCoARpMYUzMaKDOGRt9A8UAhx1Pn/yD8
DdXsWChnnhoZV7lbThbsA/ukhKuCdAZ9RpU+swPKUqHqUNDF3CY4m7W8hqXLz5HN
XynjQSqsLdsKZV464zzWC3vIwVv4j1IXomvWDprAPfdZtcCsJCR+U7zsXuxWGTuc
hVvDw4HlUo1zIBd67lPTV3VJTpm2MpK534Dc540C/zUSFD5bONMtR12BUPBGTUCe
LEZjJQs0qI9HVsNmw3aHDsdHTqRTxUMhOj4kPQsmNOd+Ry1EAQqe8wWtPkBPkIQ2
wQZGDWxK97HX2zHVCqxsc4bKiRZm2+e4hMg/TYea8awEKhAlSe1yIEOPqpV09tmy
5uPQfkZgWXEFI2ZoHS3l3Y5HFXu95V2fqPWevqGdYCO4XGzU83NqzIKwq2Db5H3X
BtnnZtSFlis3M8kf0b5b2G5qxsIIn6PxblC9Lt5K7fPiwLPECApJluLsqAm/Nq/S
Ob+5VVcfZ/I5t4TfxLh7a0ZnzQHaD9Pj1Siu6tXE0l89hNDiYilgKdR0zzA8V0/9
JP9z3op4JGPVlOzYLJn7LLyA3RigWSw6wnt12anV42Sl90h9l5plmS7k3XEh+L8z
82b68cCezWxdpBXh1inLfhNEaf9rAsy/G7S23Nyr7XmQbuNalwSlVcVhKadqDTQ/
fIOc7Q39Vw6B++zLJWvobB66/IUFOcsiMl+AZSdg/hDyqF4A6Qphhs4eqRgZI8/4
PxgxQ7AcGiq4bC6g65GAydriDXQLsrNGWnlgTgcZNRaKN5y+Oc7EjInck6R8ULr4
RqugQmoc/JPCrregpiJ+8FyQUQGhQ2FdUJw8/0vuM3QAthyb/hXTvc6OaEuh7Z2Q
ZMBGRldcRBFU08NeuM4la636zaDhtfT3wdx8PSfZckMOeIcFgOTIHZaGExMDpkoG
AYZhbq5hscjSWuS9luvGEZIvy2G5dMSdnGXRWN/QYdEjgFpgtHeTBesv6HiayX1u
iPhaWcz5yrE4Vwf4WTmqQClRHZgNvFJTlV32MGCcc7D3lgmArkqewXN6aRt9bZwI
ivY3fKxFMg79pcobWXAQ99dRbN7uoi/W8VC6LGeXB+BJ4uuKfgpCBhrSZKzfwaqY
Y+SLYl5gAL4Ki1aSOYBN/9g4XfFVQGcUGU9noJu5eA+3LGMCDowE/kvmBbAl8AJz
VcInQqB1JUHwBAPWaa5W/gc8ClCMSSW7DR8g22W7V4QaeEJoA9et1KL/wrjxWfid
4G2+FrEAp2MCYMdPfqoNTZNGMlM8BctivW9dU4sfz8i6nPS7kFXIlZ/9o7pY+0KL
7aIo6lmbKIaPSNbaNXO7vusantmGhgvW92+mCEMvsCZ/cOpfojjZjeVGQXQdTMcv
S2NVSXN4rMU4w/Tmoj5Z9B8QSL7lA54rqIUuhraoUvquvYqojZzYwDIT5V7gqQZc
kp9+SOjy0oqhnCOmnsQc6X7bk+YJTk7gEaFxhqXcKLrS8ZosAp1J7y3IFx9gt+en
w4b9nASa8KDdHKaqjyT9lus4hFeX5p3DrL2xGCHLNCzHghFHssRMM5T7ni+S5AkE
NEDKEOsbkOOTDmDTUV+Nop7Wh25ckDNXHx/M64jBZ4ngnH/P44NkYGlvSE6yJWwv
p4bmGsygn+MbmO4EtAnInGNpuXKOviZC64JMo01cG7+CF1k3bFNLfUZtUJiZbiht
nKOmbCzYVQeacHKAMCQMGdHimlug6TdsCsa7B7Gmkn9o/eY+YA4RqUu3t4pexjKp
TUuarWBabruOmjt1N2QsCQ+Fa5xLNRK1L6a2SeL/1U+SxJUQeAerikI590Gm4kI3
P28wTyO4xC4MZ71tbIihq5pTPmtYcAt0HAk5TIhyb/CCFFvFxbnb8AJgTY+XE31k
xd5rsVhgdA0Rg+gXg61dCXilo2CBaW53MyjHWlRJSiVSsgyaGxTReY9lHqb4a7+e
ojZ1/HduKlGrtA6FaoTN+mvugsk++h3H3TPf1fONWhW0S/jJpXXWXyPnuKaPlffK
DP35ARBoEB0WPlUatPc6QYE7sCOsFYZKuDQt5v/zpdRnW7ZJAPxJ3wPNYB2WLXwe
1HiTDMKsCWbW9ILgweEqk8jjenH2SKYHNPmaoGjday/r82vDqZToX0TBN6ZYnDHm
YLyvT2ZSFvQBZn1oEOVsDyBz6mQTt7LBI8BAKxqsp7/zPSEALCd4Wu1BsRGPwh9w
SrKSwF8lhYWy0p8jvBWuraRB1Eq66L74B6sNpDo/6FilQINXKB7u33XkeoA7Cg2B
qo4mfkpV+knegxGDIALHnKlW0g66g83eUKIU/neEWUV1H1jHtIxUUU1VzssGmR5v
66GY3COIw3gAIC5VAl/wDlYrtGPsIg4yYNj6JpKYEG+o2+YVXO4s1ys7fSu1DgH8
qPBy6ocfWNSNyR7qGNH/rQVFsMUkbn5sPMzysYt4Pm0gOX5xqO0kPQhikwYxrSn2
beEKuZd3iBXkQA4SCgr1kQWbnOVSYqVQXu7HFz+sk3sxeIOtpoP8359EvAepSIIU
ApCysq6FToVgcyOoe5Fx3J1mBhu0L1ySjp+ZM6G2cryJ7PIKpqmL6aXOHY+a5hzP
A6zIezFoH/GmZh3m+BSGW7/K4Wc8MRpfiehfXAme4wm2u3IrSounaSlpBlnfRuTv
4wXis0rC+de+g6mFwCbunKolyyS5JLFia0BpyiwItgq1M2Y8I8uT1NfckacgHxvG
XJ4EVqRtd7IxSllqRt1eCJeHmj49qSamz7hBslJldpDrnvtbh/k9slqD/ILJirWc
OVq8mx3KlhagHIs39y7A5BzL8gb9er2rSa9fo5vwJjCwjoevSNl+mNzr9L4nqPhj
TUPjqTK1/EJUmY3Fpxp7KTrHmoF78bTZo+MgctpLpl8kQ4R0sIT9PYGCesE/662U
FZRwGkOLit7bO3Cy3JYfgxyt4MNoy9Ze3sxoLnFZ4/d3NJWKYzWga6wgzfVau5NN
rw8wTgTx+0LpFrJUG9pxTd++qD7TIKW6Fz1YQOZO5PFYoIKx0Yr9SPBhfRNcDvFM
srs/PaqBJvnO+rkl4lNxkixXiyIr3OTDMuM+VwLBybu8GNwJG/2vugKVUMg0kdBC
nprFzhe2WPjIG6USh3s7xrjDDo02RD6gAi6Mihb3Q7Kfk9g8O2xdi7hQ44HJlZUn
QQ67OO95qMM4NJJSvFngcnw8ckioRE7MyDp0qx1fTjXp8SEzfwNBzBQJjbpSxekU
YGCjfQUFyfFyOd/qEhcmz7/kPZ99MTpeJJ2Q17zZXvnct33U3OzrNxsUoPh/sS3A
RpV5TqN04ui4AHUvdE0UpLVqTC1B2ZWmKqRhGL9t4AFA8SZh1GrHR3VrevK8yYj0
TwzJLCkP1Hb0QwKnlpsoZXMQutSB8PVQt1hTTsEN8Gbay02HdnOSX/Ew4jegQI82
V2VrmRfR7dRhDfK0dOI1QOD/DId780b4qEYfbB1HreU+xcP/xC1k9hbLf9qtQ/mh
EwDg6JBEi+mMUnY8ZEv6EinymnD9jRq7XCsaz3e2CfRvEGaLqihC9NYCLdR0eP5J
dHMuttAK+W0ExuCvffIO2Jap5LWS6/NWI9msvUHdE2r/KSBMIswBq37wKC3Jpcbh
mdWISWTUzsSzOENTw+vb4LYInCSTDmJyt2f7YhQ9dI7TgqEN5lEunRwQr2+qtfTt
WvZMArifoym2gxacbRHz7SuYAsshO5eOO2Pf4L1jXQjz8khSPIbcrKF2Y175BZos
VpyFjHb3uyOtzslLOv6B2f9I0HLGmcIf0/UBAnj6AZmEl9d0xqrWzum5H1s2kucM
WIOAScvdxtdNFTOouUSLji0sbnGZcRjX8tw2m6fYUdTAkHmuAwqQdm/LkloQAg4h
OyFzLxcJkztFZxkht6pmPlFBhAODOp92o0nYVh0wzn/dvKHpnoGaUEshfFLAMQFz
ST8CyTJvxiWE9rlMNtv4EUFD1aBTmENrAcrU9jZk9XgLEvKOoKTmsHnY/gvCWHLB
M6hqAE/oZoJmrU3ELOsh4MpfsG8MLXpnXoIqvv+QtUMR7NzZ3Q7uw0SExG+MhCSl
`protect end_protected