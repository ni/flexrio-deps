`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8496 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpulo5ukDc/tRQVITd5MlhjyJ5QFOkWkILPYsM0VQPyfck
7MosXKRUIFuN4mhpqKZaP+5ePH0HAYAsCq4KbKDMNyACMPEO8SMAFMxKH0NN9blG
wPLdh52FGWENsveomzOQB9jr1kuZr6mBqhtnsNlkimcRroC6rikbP+asELwyaXxv
Qpooh5VKL0WEgdXxhqQI9F0rGBD/DwRNVIF/p2bInNDt11nz+PzqZd9PX7e6kJAT
iIV5xJtAkQQgn4EvTTF/yumLM8fvRDKvx8CYpHZaXEMT4x4dpozS5m+LksToS9dx
/ovDxuZ9NGCuGpcK5zuo1n6sdn5Cn96DSuiPRp+3maSiJKT0QwmJTIdwgpPyTKdi
xFUOF+Vdd5Gf9kLkXdUtJKi1Xvf96sdsCVh3bC6PCeUDRNS742T65j05sl3x9/Dl
xSzEaqSNG2IiukQM0Eyl4ueyeMx8EqPMIa3ztm8hVggeKLkox8SeynEqgCUCNGsd
72eDCbRVSb0VZCztXg6/DiCRtxbaF1GXfRmN6B/arTuzjorFRGPqtYFObY8etCf+
NO8cCyxwaq4SZPtRandnySWJBohpvyokoMeYjskgzegcI3gZzAFZCxLQPKHLGLFM
4DPhrrn0dD9l2FDx76VoTvf7EUZEEBwrB8OG0RqVmZJIEWx4HbbPNc64adpGPfHH
zevNbyo0NJigMiHrlsQajFOyYabKyxWYVXd43tWQ2JNreaHTz+rlAuQ+8jJldg3Y
agzJTrNv87mh4SS8/T5NMtYtCL81auqBO4eNjYyHAMzuI8k7679mJfHm+9uQHoyy
tLNedJP5A5tdsbstaSfu8zkEyJUAuUSR37qsYXQdAmF3c8aBYDynJKUmncJOV7pf
bZO562d6VYbxdE39CcqKLKj0FD6GlmUo1iK/9rU4OvehwaydGGKIPOQkJ+2YiVr6
V7rW/oMomW3U3o/mOwBx66V/NE4S0WFpQBpF/8OLHCo33ROHefKLtvvw1Uq6yt/k
wyZpvIXYdh3QOsDG+Rdad738LcaCm3VI1mISX0XnOvANFHWoZxDjCG4KsFsDfSUO
6pue8Ojbij6lk95lNpEyMEVFo1qPgudcTdYQVECVMCYTzpy9ouI8+KHY3WPHRt0U
KyQxL2BYFBT17ecTK4n7SqFj1e+L3UYp+M7TvsaDBgiz5apSrq5SGw7qSkBNPbgQ
3X8fapn+PECxVjGMwfEfzgnBpeWoAng1jwzm3EUezh6aznPZrP4jToCIOzbPikWF
XyDdauCt5uaS5ensNutF8Gtsm5sN7VGFTxWRLSxNek5CiagxfQbvGaBN9E5XORhy
raovxWYKs5zMiNp5VI3w603+QDF65vJ3CkSN9dILEzuXuOOdl4c8C+Ej0w8+ApsO
/KAFG7dw5nUE9zzeY2ID2rewvJuPykeW82AnuxESnYVB2bzrkSa9Y8jbuSi/qw6L
oJBnMJbnhZ7AEziCs577w2XIgrof+boRoNk59375vxP6vjlmpR9uujcCaoyfgFRD
jTP1Ym56/qxPYcxt2zowbG0ZqP/5sQB1Byu5ZpobAOkgJtV9QJgAUHrBKT1BqKSe
RY4PAOYGbSyGfy42PQXRuo1VyF1YX86pxuPBgEy9QyTR45jYntuLVlFfuu83Ew3b
zOgMacRq/SHoOtQqKOYuxHdxEYJCoKBLgJ3ArxkVMtsmYT+L2yg51Bi4LAKa4/ft
H3cIBaSXnBcTtqRE4Z91OxpF4XxPPmbnS46DElNKBsrv1SpK0oUgwIzBRGmPnVzn
0cgjSgealPmarGjcVTyqaRgOU0AMhDvw91redRMrXa7WQ2rro7xy5Nu276CEiiwE
/bf88VVBgN+ClLYNzniIQVRKESsc72Y0zofX3HPsAusR/uxnvfg2NxXMzNWKylVB
xu2n5PVKDR8esjBI8Js9UzBYyWlChjKaprG46kE9ceTtx1VDRZ0W+w16N6juQI9M
xXAbdIvlhlxftRfcNzZ6p6WvikGLG3ppVMPg5qlRjUPtCr5j84m3gL+vb54JWMJY
oxnYi2ANGUKpBLjltIx8UKmcuMUUnADQ/eaT7rIROF/IgEfqJF9OPfdmq6HjT1aG
rSbpW66Ykd1SP8BXolTNsTkMB/BIur4oPVvjUcpvgsi0OdNtJoYL4k4RKglZJ3CW
iJ9I/s6DvfRnniGFWXNZ6ZlT8m+YBAWBPWomTBTgC5ETzZZYWn9dcFQq1f4j+bJe
ccF3xHRwyLvaWhTps2w7Ks+CsrTJ/2BxFK7EA/5ms0OGQ07ptpTL7OvWAPaKVfCl
1+f8uf+5YKxcgH0PdxDq6w3a6OT5X4FyC8LkxlJ85HFVHV/TPU+H1kyhi0C3oI+J
k0w31gPqe1AA5y+KeZdAgEAf/TZAhUdqyo2tl+bVfajDbZBfbfPlU1QP03D2oueN
91QOWs+a3m9xXOn2NahPKnTNaDrEnhwYfa8xJ2IdO5433PB3dbYBUh1IOP7ZSEXj
un+gxiQZ5lpiUsQ1nsfDv2ptv5nym60uSslRKOVEjyu4K+oG32yQG8UlRcFltI1e
4Y65F7nL+Djy6hkNsrlBiorv436/LtGLyhw2QrbgPuEXFChgIHRkSEwt/O+CU0Xz
Qh8U0dtSpcFkTjqWrTYGAmYyjxi4U0ImYV/a5UVVKtvnkf4ozx1EUFisDCLNAuGV
MvsgFM5zmYMcIBlH6zz0KoAc6JTzQKXqDv+dPO1Fe3I7enoEOoq05z3Rx/Crj3Vd
OQdRpNKD4xg1++J9d0/edMC+OuEzlPKJgcxA/gTLG3W2t54CtN4ACQumOAmiiAHd
BUpDfABTHFkKljb0UPME3u1xqjlV3YOBz9lth6CHiujtABsI7iH1M75va9ueKOpJ
l48VNMvo/EZm079nI/UA834dqIN+w8/IsYPPpQ6TnSP3iS0g6+J4AR4QBhPrmrZr
zabegLA7oommpc6iyIGzThpQ0aGHoupWmt3GAr/bzwOoxQh5Nbhoh0JMpzqPqN+Q
3Nd1D3UAyuBdgi9YyBUcg8gJLQpJat61N6GHxgIuIOo59UAolMLopOZvcHQPZhpC
GWQqkBx/i32P7vvhPLtGy27lqbagoGGp6Po0BAbwGYXGqyiFHIc1VCK5nr6rtsS7
cT50B1NJmev1puEO89xl1FzM8TgIbMD+H3cbr1uk2n6CyAjO6cVyL9zUv0Noedhj
8n34AWM8kAY4oWHem0QgoOfIWhszMDG1RPHxGURYDwrY7yI4sqPP5D9/g0XUclqI
kh3iMI2yfJbJDtB9TnXAYvxiHR1hXlYcPVJ19KZYj0IDcYJEHn72hQFbGiDOeL93
Ydcs+YPISjVXgRTbzrG/Mtr41bCgV5SNY0soIR4yYlhESjCGuqASvkY4kdCOqAvm
WwxZqVFHNdh8eGvjoK+HUEWH6obKDoDOr0TX8RIDUbLAdV7ZGGLBBlPbU8G7nCYR
M/F9YzhmlKqwXR7OLKd5oHgEjM1xhRWre5+jrm+W5dRlJwz4WXi611CPxpyj3YD5
uKzbZmpHFDKT9p6GT8ydFe8FVeSryX875Q9XWh9esDRqdlXGIkEnh7nSXcTfJLWC
NTG+/ftZ1k7/J5okfpVjWbD3zkdw+SbB/RtTUlgeENEtZlgN94TwhWgQgC4gql4R
Ru12hO9VCGiSlPk8Ct2Uvh8I2P9F7hVB5fNG/UWJ+RXWKPVzPKS7K3Zq5uM72Myg
bWB49xBVqPWzkznuvfCcxUl+qmg0Jgk172hgqoD3jdnNOJnUWc9hEoO50QFTpZYT
LUUi9xmdsuBmRWgF6BMf/WeiXdg/Y8dkMh5PoQADQwef+meKQ8lPiNbmhf8L9zPm
1vuBZIvCUeccH1ax9Vygk7M9MX112Xm17nwIgDKx3ZeS+3n5lSLFbdMjjp6R63te
h/Z6J6NthtlJ7pVxFGYkPRgtv7bSgsuUSgcr1O5yyqU3IUbbdqMRRjbYcXDDSj83
pPq7Pv+sOYHvBSsl73sgxL21iTP0Hpi/T7P8c3JCedsa+6SzlasDwxaF6vRxAB6t
rcm5qAVOHcridwYhmMi/67VbtmwdCOkuRQ3rYvS/ezxJcQMM9994MjmpKL216dNb
extZ6liW3Mq1v7rgIoisQyKPIDfk16vO6RIFmYkF8G20RPxZzEn0m2tdUk/WZ3ss
GP722IzGGR0mH8mitretko22XLNgQnOeFiEdhxObCWEAsi3+g0hKfHfEX81j0Z6B
bWWqliYc59+eM9mAn36GGngpWV4hnNCrxKBQNNQmFt7A+bWgTOI3RuwHlD00fyQY
CLK6GJco4NNnMyjmmV5Jqhe+vahkaxCJ4BLW30IjiP9H2I/j59hIm1O+s0/pzQx2
4fJiCfFIEaTuJKo8p8mGgzpjBud+080AAN2yt/AQmE/IG+fWhYn6XZx7J/4lp29y
TsbV0cZ1C9Cg+W/YptTwk9KM8/nMWmH8xmxLiBx8z1PbqjVJyIgF2J5k0HfXhJf9
vz7dJ59wp+ggZQ10Wg4GHRhH273IZJp6PGCkOPOCr4eG9hZ149e+doh51eHvad1a
yQQe6Pm4FZ+OnUI5WaKczXpiGwhBk0Fz0gCAK4oQ00EW5M39/EyRCMrqJogGErMP
P6cPn5ixQ9L/JZARq39zInNzvqTPTYKxgaGFwTD2V69YiDWOkqSNEgARCj+UwqZl
cZlgcthMejnG4oPAa4yifT5fiSXOI5wNUj4tN2z8LwcEzXwfn9oJz/7HZXGNyeI6
gNA7cB9cW0Zf8zi2Z8VpSYOumgtU7J3+vLLhcCdKpEHpHXBksWQ42MWzcBa4BiuR
vF+KacsrXGNLZoUiEf062q3/Wo1NdfF4qb1cNzWunbjiXYPElfnaLOhWXh96hUo5
IN6FrYEg4O5YFe1L36vCOzzplB7xTA8yBJNicHOFEweNVtraLnEjJ032kFn5jPpn
/U39KC2n6IT6hCWdq8exYI1rsnwutWfQ90kO7jJGY7I7o2b+lJLf/5rQhT53Ahs+
luiZPPspf7U29VkEAOat+2OfUCKpfcYQJop6x40t8GlQDDyBWGr9t8TC5OUybXFR
pHNnhQD4Y1vQVMJ/+zV4wENTcRbqoYH7XRQjKBxXSjsoHAy7s1uImdi/aj1WVac5
C4EayUYUDObjJtgzqPk6IBW4k/cKZvMTUQjSQ/FfW2naLu7+SiSkENe0PgXN9eW+
1ZwdsbehtfOIHqtrHF+N4+2qcfwCZK8lNibbPabglXNn6crdHKKiG3JrPOkPkOsA
iFBD1Gk+ND62XfEIwU2i68Y8qYC9zbK+RxDMxdhKTm1GGxMkDbVaijrljCP6h9XT
JBH//v5PLkr7g0xnVgibJIEr6K4BPm6m5y28AcDM4Jw9Yr+dyEigTxOLD5bJ/VZy
Gyl7KK++Nmy9wvj6+YGDE6B0774OsTzK+q8GTZN9CJEQ8BSICN40MTVhelXw+0gH
/cMnzkY1KODVOVcUK1IWrVgQkNcIj427qC1zLgETQqRdsHMNqAZPVZi44LtLqfDF
++XBz6nsloHyeYW8/OamB4d5VqMo6vzWOiwozUQsP5wIrCtq3EHEg1kvdL0l3YDN
jRtMt0xa1Hsv6GO++3P04CuAyGKSbMX94NVQRT8nIiBc2fD/HNkbm+X8iM7omvRo
ctMSGyiyac3cfaz55RLI6dYEtRhBzk4mDCt5lo9kvRC4mHl+Xuk9SZG3wdvlhQ/d
Mp7jHXj9uviLqoTAmBDQD1M4M1xpEp0ogt8v54zjRwNGwQ+bDCD+N5wu7E2UqEKW
8FObZ35UzZ6obh2GAMGVPoK0gcbB89PrHssmSDmdT5XaQfqK1qZMFlI0ywg+40ZU
Dkr54xHpyMiBiRo2DgUhi+Ay8usWQsLDd/21W4Io+8U0vwRhMhNMKbB7GHYpyACb
PGSVwmnYLxiH8xX6si/2B1+IZvm2HIn0rgaM2wn+C1yquorWHiQEiB1sfs4nN2e0
WKdfVAZf/gwsTFKOP3qiqIGFSxxM/vuELTSVAraYd3AqwNISx3dGkbkmtW4wV1IB
ju61Vxq1fqpRtrodAqmNjGVbr3JwIAdzsvLHWWuDPZt6jvwn40neHqROevEcp3Wi
W6K/A0nbw+WyJPsHmdfitskEdbqzS+QsBajt5WSTIaR+ywEpehbG7Rgkhg+59Ks9
U+jfmfuhT9wIavEm+ApxWjLkljfSKir7/7fDZF4KOajtcc2WVYUwkWLxeyDNcyHi
MunSNYpGDKRXokDh0Oj9b0i2RyFlia7gkYgtZs1anuzjB9gi3mk+2iTLDdTN4ATR
xRmDnEVMgYrBrnuqyAsC3i3tf/P4ifwjcwysmjwyug/KpSUzSoZ7Czngc1HBmJjM
FrVFh5UcN3rIDzO5NTtvY7zu/rLqcuYUpv5O6o57V/XMzPzI/TX8KI+UR4zuUzSR
FO5L2iJPk9RfnGBkJzoLc/p6AaVQEwesvsxnY+kFNMvfI7EqGKOLWRTnGO/Lyb8H
aFDNm7Ba1ygabATPb95e8iJSz/IXgQIy1HkFgO7O0u9Drecf5fuqhAs9yPX668Z6
uOQKnB5/pZe4Bv8AENazi/wUWpsJFnx+GqEzYJYsy9/19jpX0PMaVlxf7GGV4SRr
hNXmbrQOj/Wb9mby1Y4rhvXL1VpOG+piOCtxKuvfbc+iVRtaN4ZT2MyQLrDCiCyt
iUG97teh/yC4YQQRXa5DuD23Re8l6XY5rs6E3BGaAocoJ8ybLKTBP9GnJ4axPtw4
3KuSLhBbUmaX67YBwjqJW4NnrVNyrbmpwXTIsXXhSAHXO8k1QBusc41exhIoH5wV
aFZwTGhb72n9KD/MG8dhn3L+H+923j3XyWAQETAVeF9ZkBbzOVpJRZbR10W8+VqO
cVnms2OrRfyCthw85+Ywcit/ADokyrjU//c1J99lPUB2mJUj04Qn1KNTLoR/O8KC
xiVyI+VcUr9IGURsHoEx2xOPMOhbPJYMJfojj9VDWOvG3NNR09B2OVjupmC6Mwv6
4qhnfm0us72ANnXgnPQ9LwEUgbF9IfUXWaEUGIHOo/by7uiitcuu9Fnqi9YfSbGM
xKs5r02Hy9fb5+vbemY79PzuFdDV7lKVXOB3px06FPR4TygMnFp4f5ep5fYRzv/d
uesL7Z1+4jxePGwQHUe7Xxgb9i9PEJh+X7MnugAS2qoi70oizvQDMGynQr2RYWCb
rqB24jMPleBLjyH1Gz5tLU3x8UjXfAQE2i9MckvMbqu2/cIdHWP/mj3zd6aHaGJS
6W8kmBx8dxaN7fVE/FdKOLHjW5/J1BmicZtpM7jXBXX5ijhZdSesuC5jIKpkvgt9
WPVjt1Lz31Ppf/2kMyft+F8+dgdGOXH4d6H2SKsBqfMMjXT0M7SmTr4n57Rleaws
2i8Kv/qJcLYHD3SBchWhlKMwLr38A9UtaVSNOQ18mKLChfptXnMthXbZQx7V9zgi
/HwrTyyD2Btk4l5AICZke08DOMINN8wTHGf6/rtE9HSueF+9cHKMjKImZ0JKaCHf
UUTn76pZ4pEYi00zq/9n4h2pCpcMC/DeGeWpQvgHTFkh//a+wILGEqAAs44fFa1h
Tdyfc6R6ZY6t4P9XPU8tV5y0mEQagl0k3znd4sd6NlQTuzLUMQX2X5jIJzK3GlGa
MxTcfA6ffnrHdroagjZKfol1G7KvVJmWy7e9/gGyr1urjscWuySUd2HPC8u6Vn5p
EjjPAwnDrWltpQYs0mrYz9HFBeL320Dod4F7desjqTn49cEep+0BcBfEtYziLawv
scMaY/lmHIgwi3OIpgQI6bKZq62LALNfPbEhlQTHScnV36x1LKCtWCTjSgstmesG
RJePZSV7iudzoozaTscQpvAR5wOScP8BTULsK9W6W1HSViRzUPxZuAR1QzOSe3yz
eCBCfXw5ZOHJQ17/lHYliURsL9YVfYQyWn6p3i3BtEPAKQG0ekLU0bazSkGmXzXB
o1/wRL7sk9Z78EMQHk3KPyNc7mC5NgIJ0VQBror53ulUGdwR/ZlFjpoUWjLvitu5
qTN2ft5Zt2tWK6m+Pt99LFor0fPzJKm61unXi5gZVKhoBdc377ovtDJgR0mD7NCW
idBsnKMXjP43iN5Y7F+O7Ujjj7Qozhk+Ak7bpZi+Yy+ZyqavJhw75WEuw8/B2o3D
8B0orNF14t/nsJOJG+uGO9vdttV5vanFKCTZuOXnbu/M/yBzerTAIyA9SbwwBvnH
oSsYAcq5EhVcO6KukS3Q/a8my3y4j1pZWmcN7rLnZk+2m7mX3x9h/ehU9AAneopB
MfgxvMM4WGHEp7Jqy0CjpFjXUjOKMtFc697JCa1jokJJUPiz12iyzTM6WmQPNlyl
UZaRzc0HaXo6XFs2i5y67ZOsBtnZqUkLVN8h90s6Dk4NU1VQ7Xc7XycuekfKYmoq
YwHkz6bYCVIjOTN/eImRcLIIRMRZOs63bERY7pILPpEbLb2Wsh9l1BwYCHkF4AG4
QaRqMQnlmpNddFyvrmAosSfhzluFWPof39gAn4+RbMAs1rPWvO1HlaYLBoiNN7ha
7iiETwoPgK7RkZba0DVnsD8RgD582bKEo085GZnJwuAs9JseV7NhhqtY7dQHnlKz
b2YlkeFzmpH60BojiFXyODDGuddfzoa3p2zxIJ5OQYZQfpDlig5vIgomwDvvlPqW
fU4TDevxcZ6QlXirMkN3x3KvvXzyO5CkO7KBaN3V+4Ecv2rGQ8Us412oUOiz0s/+
SLzm/eL3p66sMw+3+CyjBNDRJokmXkiqCObSG+nca95KyolksHrnXE/KXKludxBa
36nQo9+4fywkRtXRNDGI7dITS+qFrbv8nbowsS8flOYl5kJMMV/9cQE45yRVtHPN
Roms1oVRRS62iNwByHlA+IkXq+NzlUgKJpNMyEwYpqaw1aTfE7WhHodcioELrs73
p3q/PtPG4VROkZsvNcf/UkOyfRKkYddHRki2JZMLul+b04egXZziQ4gWLZvAb7kl
Ow/B3sgzXiRyU+uanICaJ8il2C3FicE/t/LuGGDlvcHhIpPaGH/bxi6FXA7XCpBX
mbHPdwPM9XChlACSy+obknePl23FR8n7cjE+yx2CQ1BsFl7kvCFSNTnIPMEqVsMF
09NySk5owRj8txBv2ypuSYbxuHFXTrWMai3c1c3tf4LngMmvR87l4vvUkQoITRvk
8kPCgWRweCItDaGqe+hTfbChNzwLshHTHZNlqKS+tSSndpDnMyr5isqCW7LaFxaM
YzljraMYNgKRKOH58YfT1yKGbFY5DOjQpUjmTb2VzVrK6iFzB9g1SWQcYtJqG8V7
3xIONnVaUb60HkRFfyVZKY6kOCwAMxvCEAEwNCLALwXRsJabF/s8zdQBbTHjxFHI
n9CsgKIz5YEMteOHYvfbbofzSoHYXH1eFn/27QHpnvvRe5YJ20SrO26+TXK7Rg2J
lkYp/09HNHe8zIE54s7hp4vGEx/WZUX1asYMzA7toa5cPO9f1h7s0OdSPaG6JYgD
EMNXOLqWj9/e4dGao/DcndxAfun4dLle8uhZHAqQ6vFnlJ5gh4F4rnaL8ThCvaw5
/0k3vHoR4beAtguAVb5Z0YRo9VN3dbLWzEZ0gDzwmkj081kwhhwMsyFZWO5NIKiR
edq7oAHgH3hmA6Bbm//pN+bVk6/WaY/m4eZIQZitusBp9VLdAT+xXhW+cqWnQSBS
E6clr2HNX6AZaE58R0/pmQZGBbbVFfxsP3A2sDQU2EGkS7Zv0+YsnW9dyWwsiuIo
sBnA82bl3eOYT2Jc/Asd0rABt+JKXH5UOLx3hZAtqUyC382SyzxlQ3Pw9MP9E9N+
H7BJ9bF377E15eYw0gsMl56YbytAS0o3K0QW7e7klfwzJt7qutB7HdcKyIcYXwXI
e3ryC17nACES4TPRLMxgTVNg8Iy6xLx6yPzJBAVTNFtv4hFtp3RnJyoi0et3Eynh
AEk4U9je5CyDuacrvTtFUOHTtJAtKLoqDicfBRuJdIJVdkL2CVE1m7DmaK2H/cua
2vziIkmopF/w8v7/ROH3jNPQ4L4kC+4dbFrCtj2SavGZmAvcOmuYV1+vh9ESw03w
wihTdOZOOQs/z9qlqicOBzyexyYkniL9jFLgCtDBt6BAyBT9nmO4mf1sVicxbnUC
WW5jKJK4w9w2aHjlmPBNso47WwcLelN/F+QCknkfLhgenx+H+dJuJUhPRmNRrIru
yIDZt9UgJd6+s6N5LwvE8epsyTDAutugwwD22+ESj/Nlt8vvUD6vGdNYmlfIJfte
ai7IRwQDWcHTBFpeMEpcjOEf4iMeTt6iSaV5ZzPCHWYKdLeloMf61WRC9IbJL1sH
npxivHYqMwe2hWQKYIeSb0ImXeKrxgxhK1Ga4t2cN/N67ZYRiQg6ahuUBiCcLmOk
X3sGP8mzoXDabxPK6VsTokvtJNUwtwVSGE4Z5JmnpVbABvTejCrYxrQVtAEleisa
pCLe58iZRlSQiSSS1APGsMT5vxyUKG5YbWefE0sEagl4zcNshMUj5Io9cjyseZQJ
NePQilPj1/RsDfUKMdGQ2YXDN0zvTQwMiQAWlw2AUrCSLVqEFM/lnNjYPxV9DSd9
L3dvnyeuf0+/m/68mwLHsM0TJmjx/OUOLHcNpjjM9+UCR32zOs5P91RXOOx+MmXL
ozl6zTDwtw82/NxmE+Pug9v1Z5YUC/31eo/ULVASHfT6oy/S3WJKbk69dvfQ4GWD
syS3VSOxDvNzL8B/iyFhUj/rZ6rurk+QWeINL6Kp1n6O45GntX71BviHNAUzkm5S
lk4BXbQYsCQoi/lW4mvSLVvQVweIU+98t3QdrhLbR8VYGsArZijR7TqeQi2jWMx/
m+13V03Mw3mCLMlFfbI1G90bkpxo01p9wCbLKQVZLyO8ZF4BsV2rJp5vJMmqmSR5
b1zM36Vr150Gi1xzGq1e64j1/Ti2RdLjw9thfIWVGQBhXuvyNLELqXVH7uxAXM4I
JShC7BQUGFSdrgQegHA6/8KI0KbGyUpQjfrtHHdm2MjdJr9hNcdgs3sANun3q5xo
c7nvsoBNjTWqiDTmhNrEipzuPU8IEzhzOl8g0wnGTP2QywAJVSXwLIphDmSVh6wJ
OkvHND7kZDUIY8jFGMPKGUeuvp6MJHoolQ1EpX+DhlPH5X8CrbftmvF6WPgn24Ol
kMpTQ02wJfQHJVSzTpM3zV1Hv/5GZMYQ6I9NsFbNBJjtT4aPLepXodulJcZcryKv
`protect end_protected