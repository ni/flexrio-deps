`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1872 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIbpmYfLOJnRGfzVwv2SxRIe1z6iYyUz1btnTX1HZ/yzcY
hPz40E9y5d9kUPVtTSmTMfmDarzRo0F/4+zULt0sHRj6upKmAqGrO2gSBjkDV7fo
L9APTzEwQrq7T6Ae8M969YAB9UTuIuwEiw6IPp9Ev9s+4K45/eakwVq9ySGwXJp1
7QprgQbD+A9pIEDgFxgJAs+5Peh1r1ddOnHrd+Eyc5pgc7UGiGDtd9CIpaY3cvkX
YPHmCTY7uQ+NYYCr/7xXKTM5thMRZF0VKrLWzdbDSVBvKkJD6jzwpr6Lt+Av06r5
M2aYQHMKn3elKs8C1ZKnPkPQ1wgXSHIkloUtC+C1rda7PD4019CZdGpIlxrwFbfF
/5TT7YkdmasVzMatYhZFwrHxMTjxN1elg/x8YeQqFPxkjNmUVfD5qWz6k6GC9lzT
4hThSP13io8KH4p8viAMUiZGFFPSr0vTvOtIrrIer8P81jswZGMb+4J5KpUJLeDx
5nYpqIbuPhrYvB4SkatLnnaboLso0hvluTEYMJ9R7hhUA8/r/5Az3Irarxks/ZQE
7o0UBImDuXOqeD9PGVcbZZhTo2TPTwgM3peckzCxQI2vOgzY8OzCtFPMuk2YJ9rF
ue6vpv0s8Eq3QV5eLcMRifxIuAHFoyv6HEahtk23es7tc2yMpP/RlAcdHBB2gHXZ
Z3OO0NKs9tbGjRiQPq4jnXA4DNxS6OXUEBDAnuEAg0GtD1pSIqxh8qxFqur0R8LZ
UUUJCyBh7k7dmnQ9cNyrLPDz73QCq13QYmJdon37qo16be5ZRkXiYHTqiHMqSYwk
9LtYz1alJ6KLquqYLUPbq0JYKTXbi6P0PnnwT8fflnlbIYwO5I/myESP7/GBkJRH
IKP7GQkcLOHVu/2aBUKEgl/1mUP7Uq3u91k8kYkvM1S2XHcwinqay+9CyKrPRKyz
SeX5EFdDEjIzX5RbQk5WVg4gg6rp70gy5QYlGVMBpPTO0S4UWyniaFLAxOCxTCU3
zCCfNeWnOQOFrA6ZgJqyVvJFKUsWssYok4GbbEpdEnka9zbkWMKUWxwzyxlqHDA0
8ZsxtoQlGZL85XPl6UU0CewAyvV/4Melxc4DPFTReZmmKFzSTwEE8Yku5pVn5ZXx
ica9JhR8rG1eZm2p/kqPMunNh9ncoOfV8xPonfTGGVs4r/iC3NZBwMvlB/Sg/phC
InsoNhp0dclTiaXf6rDwu+P1eoDp2jhacNsujgLiSvwG69Of7pXcb6gjkd4MR9xN
JaDDake9WLZaDh+1VYPTjW/LsjYzVkeZ0HhKLE81QRv30tfOtGRKY3ybduIz1rl2
lYJKwAD4pbgMWLe3rhrnxHVaQatfBXmCbNn5l1KS3H/3uEjm/btOQ0mOpjnVBfuG
1iTuQlDw50G1AgI3uvWb4Lt1VYIqos+VWas6GflyobXvD0CyI7kPc4dC7mFxIr/T
cs9e9OKWerewLWUygH0/aWd2UshsrJ02fXBIg8aGmoWNXKLp67lO0lChqhSOFCZD
ZF1/gdbzxGtgXKgrPHxn5PCfpA8V2XhvV5eTt/7Ct3apJ0KIkVpRISp9Xj+wm27d
ggDwM3khqjdy47z7FZUXS25zk3Gz0LQK4P9o95JmG6BwQguNpDmbauFKEbTnxESP
8bfEOUaXYAz0CcDkmFt+e4LyUbSWaDKuuqgju1B79SRaEszHvg/KqL+MWn8UqZDo
M4R6d/HrlctSYPcRGsR/zS71S1HFbYc+FfFDeuWBseYgFqhtqOgwVrKXoPaMcbCu
dFwQTIa8Xjh9ytwe+ChfXHc1RiHHnvnLrgDvnDGbHDsWCrbsNDUtx9nF3Y9dVYyv
Kj/4wWiU8/guO4B6vPS/Vwykf/N7wKCF6SYyuaRSmCCMy9PWh4e35Ye2CgsENr7k
1Gf+yre8nMGRV5dc9Dv1tRXn4oA8xTFP5n9g0mANddaxjNbhpCqpvCwtQqw4gzR9
6FSUQXo+YMtYOOOOqJaPX7mOl20kDjXxThqd5jqwBwERf2u8lv1x8j8BovRjoyoI
56kUgknMwJH2s8aJCfUp6jm7MAIjyzsupoqtpzs1BeEWcoQctsKfRN9juBH922vV
vF9htCoM64GH/IjtlezIyY/lEAxaxsGNdoewDAZ6ExS5PpqDnW0iKCIXsXJFX3xu
i62nSGgsNNCtbrE0BsQ5dqtn2ikqdU3R4fgXufnBjzVpPBCU47ZQF8/7tzPBfoD8
iKwe+JRCNXIdq/M62cHRFylA4025eLC408FauBU6vBemXGWlw/E0CAMXV8BV+A5j
q/ZXZdT6KbRA+k3rPchSb0Fu13krhk7UgRr9vMT1ENo6HSKlgaZ7MdooOcP866QK
`protect end_protected