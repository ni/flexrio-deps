`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21376 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JXz1+zHgF4n2s6TEZD4KtuQ
ATkS0e5WlIVeyjNZ91Ns36sZQfrQ9R4SbnYvAtVIyXT+yyNt/4VBW+6AXiYLBtjI
zZWpsDIlMr3WW2xApDVyUJ+BV0yyGYfi2I+NWKxktoe6A1qwmwHxLoE8bkMHiu7g
dhqnqSME8c9Ag4dJY4VTuuRJ4DZf33E8JcAAt2X/YNTHWWChyfBEA5mNYh4ZJsHb
hR/DNUeUGv7yym19HmnXs3z9AQY9ZprtTzFUv3nBrIYkieaq2b/uAY3HEBT4zI1A
rHH7E+pLM4XWlsUIACzFPv8lhUg+4ezoKp7wZsRynAf7lB9Ogaed8/H0ySKQknWq
CBJxIamHbMQRiB7uSgT9/3CjowWCQEaqeqaEYHWoCpN81b/hpVv0iP9hWGbQU0Ig
nWVmjFnTKYaVLQWpkCBzrQViMt9SBsRpQn9abKFF7sU22RRLyrTWj4oCBkQXFVZS
hNQJq6Avay94NLVf/2CA9fmydSIL6IgQrSd7kylcNd06EtJCxeSkayBvSbCpQh4z
bmR155VgyoNMhG7jQMq+qVe6/dWgxVKWwtZ7Edy00WeMT7stzv4DgQtuCmg7HMtc
1c/koEsr78jTh4QXiiLWClJE4qGbSJ+TJURRdR/ydCiUNT/4es5j2fQHYF+83LGs
e45Jr4voUM8SSk4eecrgQtS+d5qPvzR0tFR4G96uttFe+Nv1U/3uK4iv8nmwSct3
LUjR1Epcx+ziZvPRfLMXQJOVj0vNwP38phk/lEmoX/mUOcpgpYQXXUkkwd7RUhdL
qPTeXyQqpA98ix/X0Kv/+wpjPm4ZduMekb+WfJuXHoy/CwT+2PCWUmjq/wd20PBz
+017ciAxRpaL6DJtgUW19ZdrjkeDtnF32b+4/+KDIA45yisHkeLbZ+s9qIW+8MO6
XEo4qC/Sq521f1if1Xca7fBMz+U4plyVLxKoETED6i1DTJP0toy/moBm1aZegdFl
+LNlBEHL5lRQpYX/wMZyk4qQBEch/M14VwPXAmncbhvM+dJ7VJgkyjTKSow4F7ks
4vBCv3nuLbhIKy1ZFp/8LBu4umQHBddeo2wLezo4qD8B5t080SEcrKsiiGtMh+h3
n3FYI7hgAywdsrLoR8hANDgufgyeZe3+IrlTCWFHwgbI/d4knKDFAgX0+2ziW0lm
xXHACuo8Z5VIcw9jFC/x4dYCPGUxv0JULaG5VPZw4Rv45yDu7UNBjnMzM+yqbTaI
XkxNiLjnxKOTJ5er04cFJDoKuVBEfyUCGYcU3WrfmwZghPPku+JglLqiW1rbOVwy
DoBuydg+miDaPDrjHMAx5PgSddr6TVmcminbEwL/OUtCc37hJ3DiXq0L4pDsj0CC
bWEWPjTXWqVYIRAcd8ZXMiitMaNSJB1ze4rHVsG22X+pAjqFxof+P3LQ5mvbzix6
o0lrUoW0dpjthc8kEaXZ2rEuraCLjTkQd7wp/VI9sevh7QdmnxQwgHfIas0dGq3s
XD6O3sFKND8uVAleoJZgayO4zgtBZa9dFaKSkaAjeEH567x1G+LSHw/dWqFgR0Tg
iL6H9o6TGHwgKKBomfyVhFlQ6DFOq/K9P0Vj6enyHODq6Szg+fkAEyhTbEd8eGcX
p9jP9oNoy/ZiXyrbSolFlTiuOKBMBpPlXsqV0U4EwayYejkITzMh1GqsTsWtUt/D
HryQEbKa3W65mli4Az3CKPnbBkluyYFy9C3qGsTe0v62CC9AQhQpMegkIITwEP+T
TjBoT2VuS+Z8G9pPcHPQi10wTukmFc0qQjqmop/HgX40sBjAJvFNs3Vd4mEIZ/1R
u0l86WMeX7/YGW3U3sXAghLtBOyt6GYN48KqgA02gQxGOtWJggaliJusCRSUMpdV
NsakfwE1HpvEtQAQEcAYJ85v+eX68B2Zd9YJDVQcgem0ZGjhjHRGN7yeoi6Ixdlq
IWXCpbYO6BxSwPSwRTrQqmtSOY+SVg8f53wUBZ+APlxAMcJ6bAg+/b6WvgmUhGwP
8HFT3oMhLoa91YXKNiiVP+Xb2xi1jvsMqDrep+BeIBhRQYE5UTuK2ZCi5A/jt88K
gozf4/CbJ/q1lYNlCzTCM/VY8lTjdfQ05zcpp0MJlc8Pz5ku+zHsE9H0jSqMtayt
TME3JWXERaa46wH74OaqTO63MV1N6CJFh9HvdhLn3EDiSIfo/CiQDrIw4hkNwEGs
91k3uXW2XiqE3+pxbJaokleSQ+p5/7GjFstx80wmq+sBDEgww5/b5vgSSK4UknPs
8SvKGDatwnPNkVcqKYXPmYKnGlFZbCBsZUFOv1driqI0GqG8NUfqwi4tgmMDu+Cw
Bgyks6yEZ9HKnaIiD5LpzLWW1J0O8/V/Um+VLocUvROLuyqSqlhcCg7IE1yRxf8s
ol7Doiu/1Jm0uumN8ih9PVYK3uHD1Okn3sL+9OEceDVWFVtFOg5kBoCPOkKgAsg5
imbBXSlGTIfC3dBpLMJ11P3IK8uWO+a34tt10tLANxhhJPzWu1TLzHHRFS+rC8N/
z4JLxWHsvkX/H9Dyud9JuUNutzN5nGIx/EbTQauVSfCHRrlg8+jqy4BEev4/Uehl
zRzV6J67Ob4W3nJzpb1lEISq1/1aHBtKhxWHpv8VW7W58ozrvRorRdmIwpS4bM4k
fx6xStxqPpaReHRLasrcQ1alhNoLYtzbJeF4uvFvB1pIEt9bc881T9u7p4R3sLa3
tNf5ILI5njY/403+5kAjiyqvbjOPqNzaTleEyYziIyxLoRDsHaBMwCb6CdBtQRJo
JqbJU9qZ7/ieJkO3A9JYkRr3L1GwIjNcCUi52ivJ8JY7kEwX0A586bvyTrvo8Ndt
YrsdCdxkAcOeJfcN1LgmGsIqFqiB49CB7Im6XuynROd4khuIz7e5Umagk9y5wp2k
yQb2l2ShcT9WMsvp6oF4NYgrM5mC7NTxJENIOgiwj5hWupy6tP5dVirR70kywBT+
BwoTixfLLMMEetBuCVbs/zz3Ctudr1QddXbf8lxMz5Qk7gwoAwuhjeEfPdC/Bj9r
j6mljrk6b+y/es+sXSEZlPGl0K/LzNS6RPrCMNt+d9sR+1kmz2JIaV+8o2ALeeHt
Undz3Y8eAY/Y3Zg6+Gv25MlCgoVmBuGELbe5eTo0eOPuBoictPT8CVc9xajyxfl7
uiRjdj8+uUdvDzdXVa3yEnV2SBCnD8I+I4FTZ+7OmrFGVNfust1llJ7J6pa8tOBF
tpVjP2nAvdJZzZijhmllDs10+QbO/98sP94mE0H5n0ZmhijAw5zXo3LqCCnvUqZu
AVZBQGqUfQ3iIIRgUkOziJiOkVZ/meiOlOm3ugtJR8xq2w2XGaQuPpqNTh3ABgG7
PzfQh5ieF///I2vWDdlNBUCoeOuWp8s1H//Vhw4BWNB9VULlXEH791DTDOHhsh2D
lhxAabPzYrmCOsJQLzBwqQAm6vGV9Djym2wBZoTsHSO9z1msF9ToRMqmPRqAcsXg
35HyCtmWHpJ/Nhe83gJ435bfHnkXnCXZGzXDnFCQUE2Q7Pk27sOdd7Y/PPRimxxI
/IlLp1fGH0N2HUEVnOI0ebQNmHnQf0ZtpxRCUuMFAzEOrWkxFPci410HbjpX3Nm2
Dr5nLKPrM8rYnBPD56F9a/4FNpnEfg51PesmbCz2MWYlwvS4z1Q830tWFrplbWa6
lEvSX7qdDFIrK/NNySvujw9tS4fudB8hbW0o5Mpqg6qKj4kL9fy/vk98xi3GoTkY
EtJ+PfhbsmtZMqCiDseTGLxCxXF6QEaCBMM1qI58FILvmDgvLG0CXGGF4H5v6IFi
se0y8BF51xRNdlGzHZZNWlOGYfXFWyEK1iLMimGYvRZluU//8auKlLVY/cFSQoBQ
R/gvXsyJZUKcXs9eacqJLoWc78nW6vZ6jU6xxHsT4XptbeL39jv4Do/jRgcmNqdu
BQqs+LT9ND9LCv0b0ep2uXXPSzlhB+KR9cEoHeHbT/HT0EA3hBRzGyujUNulXXN2
LgGm0w0reSMDpjY1hpf1tXNpIc6eENH9U5sa3vcO8+BEyF2FVQunUjLPXepzhi7K
GyLPJbRJfEOFSJM/GouoZ6J+QebtLt9Cp1sqlqWgMgcFHoKMlapQ5Q2HUQdblXF1
VhH3I8r5lqcXm31M1SURD32mUTdA0k2b6UEt52Grz4i9QsYt4lWZo/np1jwfhaop
XDILmDud4XSODIMaQ0Ahxtd4DIiwPsVRX/wHOZoMlKVZsXcohTumiMi5blHrzouQ
OrCW0ilXiJwtUaJxNm8wmcZSyt8COt4SuORLIzS9sgt+q38kPhRIejiOcO+F1qcq
8uD+M7+aGh6hJ3K/t/5a1aFtgRZbPM5Ds5OTjoFxMrtuulmhq9q7+kGEKpu4U8ar
Yvv6dz6/CyQSUA5oX3VL2y182YqKQ195BY+8ujavmp1OP5jMdktwUwEqsS4IoVXQ
YO6SaN1EvUA5NuRrhjgKivDgK+Z2cR4Bkbv6HhkE5cdmlHRGZ+f3zJMPQ062EOYy
MNZIicW+aE8mhgrNz9R+t12/PicgsV27M+x65QxWXZf1e5wUeJVUivA3iArDa4Rz
WbZ57OKQ2UGFrTZqy5CCT7iOLXOYjKoh0TkVfj8AUqZ0JD+OvA0fkkVG0QuAVz0C
pEq4i6t5VuTRUiFWOhSyjMHbPOAzp1QP40Nl0cNHidw1GemEiLOcsZNZto8miJgX
ZRLP0+rHpzBEnfEsyEGu/NYDLAdF7j73oEWjt5qrtLVrqctm46Iky/fmVM80Ek/W
8TGnxymMN89Qji6ZZfmD6bUHuFcpboeqyCNa1eBTmMeYTtY59rZPqetg0Fr/lwZo
teyPKM+QN956lEONx+s11IZBmHbmKwbbD+2MwAACjeTwh8qZ3+RrVW7xwrN3H/3z
H/DgTCCyye+1PgvGo8k5ehtClG10VU10smJLl5r/tD1q4IWdctNGaK2cazbygfzf
QgB+jbPpQYD63GJadM5f9IrTP8mUS92kK+ZIug50hMlVF0uW8Iztv7D4de8lHq/a
/yZaHtGXwNml0E9MVwfjwJFNTtyLw+stku9hF69W1RhmVdbHnz/tfDItc435ywhv
ZhUSYOhz8OiIxUE508v1N3FPQh+Y5y+I3ILg2IzINwKCiNGULbCsOg72Al7x/4y+
IpgyNmezEyaNdqYph44yY0zxdTzkC9dadociIdi89RtbQ5du1hpkWKVmAivfOzkn
QluVEu+LCaLpyKELiBNIMFMFl5mqaK58YdeF3ToSepG8goMPktjhv/IvE4YkDJds
ebivuEUpWxDl5f6tQKkn5/OS9Z5yUcHcr4bYJQYvmUZOUf1YAQqgFX+W1MN3wsd4
bjO4QN0qKzhvDB08EMGUFmKa5ymLrXT9hWylmSr3Xbh8nHAejAccT2OSbfBpij85
3TlGl3kWr1mz6RIU7UUf++gHykl8saGYeUZpmXlpJXrNz1O08EFzIBLfd9P+uOkn
o3oCSvzvjg3N4XEel1xbPs8HGrcZvHEMkErgGbAebGrZMkNNYOqCDgYWRff697qa
oBg3W+ofapgVjdj6wlIuawxzLVXeooBU4zQwi2GONMbBe8yE39hooUZFJj89xK5G
hLjUmUHowYqxjCWvRGg+uVvYQjDUufegNLdTaUXVgxSHUEl+K9cGyy/VOCxzqsiA
9uhSufr/ZDfEJu+agpCRDVXsJRaBMUGd+5wzIF0CgyDDi/5N2ANNmEyEEuKjJUcQ
TaG+MUo54i9hfKv2OLPn4Wfy4cecV6bkyA9j15Jg9CnNt8TFhc9UTFiow0nEJ157
NrqQAFGsUzC+/KvLXzq2MRYZkC6AMy9tvbbl4Cs2czKFazUFlq7k6AO+yVcaqohw
SQ9ylmQzPo33HS5N7//PgixaYDo47Dt8RnHunQvCEMR49IVOWC37TYk1k1zEpL2z
2M8tyVySWrn7/0EifoVUmhnqSUxfrfxI+m8IDkt+PuSwGnKXzzXo4UaFGfZuq1t8
NyU6e64u5ROyDAi9sKWp22llUhMm+khYM9OZxvAsUBeLf4LuWr96FaFPjjSTlpXk
CtHSajtRxJ1hvOp8hwB593Ca7izahbUMrYQWGKUsgV68/nH203etC2qMuEjAMgLB
cB9O1G9Fr0LPDfq2PbWgiWsb1GiKtN82X1jqfzRMm+Hf9MQuUnL1EW0qzV6TEc+o
4J5tfmf3inpD/KPdMiBo6f/NMu94WwUF0G0/3geTXrefCNsU2pjI6FGt3zkGXkWa
FpyMGf1jBE4GY4lzVbUUfTA0ZWtUkiRHiXvrhJ2H8n4q0Bx4N8RpxnnfAkKWS7KN
BuYsaSQURXGU/5gSii9Bcda3nXbyNpgDfwp0HXvhyvncP+JDFuy+19HiExVOCiwW
2N/y/CGJFdT/6wDLJUEAxThBGZRX6H9aSCpOtm/x64VQgSWvNIDytkfUvzYF5gSP
gET00vj75vQFvMkOKPMmYrxreJ4In/k/KoN7DVzRdR6cl7yiH/+SVGaIeXWxh+Eh
dc/Vhtp+sBlrFMsWDcF6sZyAv1rIP35cgh83Y4cIzNtcbM22Hn1ZyA0WNyZQfzsz
ohW1daIP4So2e0bVkzJbCQ5kBPfSD8Rvt2QMQWcQlabKSk28xRKq670N/SBQlssZ
2MG0BSacO3nsLwbbK3LiEdzgrjvdRJYiPNlNC77RgNDyA8a+Su6tXGoId95Xq1FM
WhhoD26ohE2ntybi5koqyjA32SNq5gabtzKryDOCUqoT/GZziqgwR1Ete6H9r3HI
w8R6XV0UFUBPFIrMTcfnLld9Ai0maS6JEB7G+Fy+JjWbpf0U4PNdCykbED7TnCOW
YN2dXFHtZkmgSze7GWtGph/p3zW/3ph+tndv2gDhrH7zQyIfYSS/bljMlltt9OR+
si27FhtshRbPoY/LBkUuqaRq+5DJxgTbC6Sdh0bOUd2IIncSXtjfS9ZQI/TTV+Ea
Tr8VjrHy5QA9y3FhnjRMgkLvyvOjUGOUoLKKJx0P0myhBwDBm2j719xDwBTV71Jo
XEK6G7kJXMOSty65i1BbEv5AAyN/KtlX93TopykE2AHr8ml+BjT8of4hxImOxf81
lngTVQSJHP/S2UCN2W8NVtSY1MkGTkLnkKy1T+lb1qZ1Zcczbg+HbcyWcYAjd/XM
QIsIGQtwlIDib71B9gRkPxd0qP2n6LBhk9j3ydtav51IoMeiDIcjLDGtIFgPAYtY
N2zb5NXDR/7XB1G4nS4jriqOcR4F65wN0y4QENUX0bcqbqiRdpE7RlhIiG7r935R
zZqd4fxk8AjyqiAU3w1XKsJQIc9S1Z+4M1EKGs4p1ClMhMiEOSk83bly21QRmfHp
nI2HGK5LmYDu+wN8Q2VeMc5jcTWxwJM0poFIb85b7FzDEopPPr39pfGObe6NfqLC
UZ0SwsbC42HzjcaLWXde7vbeMKyiBY/kbtE06HLXMG/nOO5CA4pvIu2cCzspD3AB
P32PJfFXlpT/3iUHiIjI3NiRkJwIARfnqVq8aN8MM9xvltZSoIqu4yWMcihzMLjI
h4CRxS73sEFMwMxWKBQWdAvBLC4BrxpUzpDLGRpux835S4GP78pNi327yfajrlB4
RXgUgz/oh6432CFna4i4YkGNnd+1eaDeQTvGFFkg1OqAt3HY7kPC9JDXh7oUPUPE
RslxQZwJvXES29NsGpT66gk8MLSem4zjPlF8InebB/2j5ClhI3b8IF4gD2NV7OjC
sS8iRyKF8p8F08OYoNBIR45vfVoDEZLjol6qJmYiwWX8iZfhXC4OXbruPOzk1Lof
bl4gt9/vpsKAdhXufrlLj2Fb8bM9R2+gz6ArtcFjCtIKodipQfXE/nNmlkEZiIuB
3kd2mV29IJSZAP02fgei5G0WVeHXXIWWjeuzM3dU2Zhd7rDrN0Qs6PAqsIrgcUr1
cQFIROKySyy2QGgTBdDGYSYvqLnS4OIXGO2FQbMfbF2UFC111musudlYvvWzBgPq
GlTSHT/egTO1byr8fcjEIuVD8g0oPlCWRGCZflqAqoVVOqp1+z845FQI7zuhMvDQ
nqrW/iLG+Ewma+MR+sAupmslOOpAU29LRdfg1eyCsxGAcaTGG3th4U7L+O8waKth
I83ijugA8XDpyNp/UKNM2Xg1VUjyLPRELPfXMGtALgoQDyiIibtD4Z7ohD8COFMB
GQiYeMDjcbM1bxoC9yeNYmHuuFo+xR2soroyC04DsyfrBpbcfjGZMoXPG599HJKB
DBQuqbVshAiRKy8R037HYHHtY93j++ZRBAQZQ/MNwZHMbsaJ1zoBtJ0Jrn2ZMjW4
q9Z+pP8Jca8TCvf72pVLc/UxmNM+6R/GcW3J640hUwNNShdWB0CvWPRIR4E8U//R
SHiucih/AD1VEsF+clrrRsnL+eAstgXTTpuock/GhSZn2bra29K23iIGl1qA9XCu
zKTf6vHJ9JVM3FWk2aQmIp5b0efB1KW1i+5bhDd9Lj2JphTpUujzFZpEWCBlj47d
JuBDF9bKzz0HEr/kQgt+971WQzRQKSH+tAfVwtctltH9uAIlRbjv2WfnZUOxWg4R
YT3OyUjn6LY/b9x5oCqf3V0h9+fnCJDthesMC2CLy0I/eja5a+LcTqWS/0bgJJFA
OTUM3A1qcBl5Z7UMP0IS87bLSNa0YFaVTbh2jJ2o1ykNc8phBu4puGRCbBvZiiih
zAMvg7gZmpjkbk0qNQQ/+470chA6iwFbQZCzRREOyriFZZpesqXsaYsoxhVmZxcc
3ki0xNV/voCxWlGtSXzYPFKJDVCDOxFZqk2uuX4bJGo6/9FzoMSI8gfW1KFFwl9I
b5l7jHCDcJwNQWcQw4FrxPP+7UyTJ/jjOpSyFyG8yPQod/bn/gAWOS7d8P/74Sig
4vsRZ3waL1fipzM74+DavZ9SoOMeEHIixTObjUTo1ltwCh5ryXQkGSe/Ck3qgN+z
5Zp1p6xLGzgUFDSiuG8C4MuLsRZVq5LBGVCHYY7TIqLVLkLwplkEc/bylzGVyK1g
uztPZKKARHbASsy1Nd5YN+es+GIhkAPjl4yWx4VM/BznknpoupNZNV0KmBKuoGgJ
haM4Lve2oLjMCPAWeZS7Jl8U6gJLqdd0ZGgpWKYDeqF1437vXq/52Ij4wkNDt6xO
9JWhEzkkZ2FzP9lxodt6etmNHaY2GkuNR9K/RatkVS3mQVrrlSsqgYOg/RLL1m3a
BndENz0H0gYXNutdWFkyb9kBjpnrujj6HFmaboA9c7G6Ht6piKhGAw7M7vpBNpQp
pAXgwTtvfSe4exTtWA9m23vQcBh+wktrnWeUI4bxC2BfypJebfFt5N0pR1nnC8Bf
iK/h1DAglKfeRFJzg1GYI8Lr8++TAEQ8tCh6QpNAWKUE8R6QRnmEs7t3Gna6aX9B
qt7ZAt/jXQoufQk6Vmkc6i8Mu27lPUTkFs0IShWshvDuh3kgQImCsgMyTtHAtzid
4cXvvx23fPqw9rIj4W8nUiX2zykGcN7hloo9QWQMiX+Tsopu7rvQUXdKi1ODDgCb
NwYdELEvCvbZ9aw7ae86I7xSMlCerhGyBT3GIlSKXbIPlqVrUsIY41oJv4q4DMw4
AXGRPeqHS4/xeaPcLdubmdyApVMZtwDeHzEFzNeJrel3Rb7senHTALT/wTci43BZ
DdK4pM4X4HPhHbdge/AKjc4CR5HQq5M/qywzYpc7FcnrU1+s7XhMvbBefYeHEAZV
39s/rJ5ExXdeSk/4g83Vl9/TMbGI8GGOxOX+dRCfH+7Syax1y/xX612AQuY80Vbm
kaArjhLKmw5Low4IW7OaXUb4z+tDPwV1KyO72QHsq/ZW8MsTvx2aTgY8DP3tfTT+
amP6luilMPmqCKJucZ9/d0r3FkT+zX+YqGWkIE1xMF7gT+8laynsNLLfAvjoRuuE
x1DOKP/3u8EzALR294wMswS0oV26bD8BnWMQs1l0nVK80L3I5Kc7pvFN2Htx4Uh0
zpp54hMrIGHkv0W78n5Il/jHrexnOUR7NOFQ0sXoQQAU/EDrBTpi1/7SKqKiCYy/
W8yh5zvK6g9BB0TecJe/KzaAgRd8FcM3FWz+WbHOwzbtpoeMK+aLNQfS3eGHKVt+
PY7Lk4+CU2koSM3e/rjDqljzs6C4DyZ7a/F4Zj1rIW32i/zR/E28dxqif7fPCPKX
apdyz+VhAsnx3gS3az+QdwyK5l/OdRiLvzqJkb3GJwR/fDopmyeAPfywX8KUODR/
ygMd8S5zaLhCH9eahmoY09Q4fDTwDc8mMFbLTbBnkoa6IPOXXHweTKic/+bqwXg6
kis+6wDwqb7YE3Q8aDIpz8/zJC3K2Tmme7HMmRGRWDCFpEDRK42dAPqemPDvDhk4
b+y1MWc5Ws29H7l7QqIeHMhC2qpaH6XIXJPHffJ/ya6o6gEGQtJDg81ZzEV6sCNS
136CodfmrEXbPvXoW8DLjk9zfl9/M3sWOnaWsPT4kYJo9zOxEDbZnxVRb/en0d2N
XtIffYeGjx1ZfzXhZJgDMSeZwArPp627qSIBwifZKYwTV82LTNXPl1bFVVFN3AQj
ZgZf9EwGjRM8rGII5H0wNhSGPG8tCA95/z629w0Jy7ggYppi8RD+xundB1c+uwf9
9YAgfQKqT0z2E9FqrefePrl4SHhQ2Xy011K6s1K8sC3lKmBkcYmsVR0JB0gAGKRC
ffzK5oJur0dfnuFl3B96gPDcr/Vxcu+4h/JFpE19g72PtYXfMsPOKfwZHzIL5uNM
c6TgopBhNMQlNB0LTPfaxoBSh0XzzcEsvVZ+JagDSpt8FYzvkbeHII36OdZM2CF2
zfFatIIqAweG9ZnLXh8PjZCKAsoQ/eILxM8fuKPI2C9qepsjzccD1PDAun6F35jT
Lz8vRFf3foLT45AcjBZIg2TRWAexsfSp0w8Tey/d/FLDZPjJCW5RMdR2qSxds4gE
MiuWZHEEY15gTgeRZqMoLG6CNPbU5ebP7RD4iD+DxgfHvdHZIcJSu2EloaQ8Dctu
7DemAWxXClP5VfIMbpQanIXr7klAYNwVj0uUMS22VvgouE+NfH56S9joYuIVwDj0
xuBvC8OyuVTD32rOaoimQrdCWdIHsI1PZs6Cbb5JSaNanwuNmQqYGxcW06Hndf16
FWBInMvXpMV8Gbxs/G3rdzAYce6iAcLeV6r6uVLl1vKzX6CwqvcytXWY+pUqDpk9
+G0DbiGYadPUiB4ufhqHlJ7wuzXi2adnf83WwLw7rW91C1jJ0Q0APypzDBSgSbne
zHwfAyUjt9MtU3cmNldwWs21yvVm3SZB5Gusu7W1ys5bHZmfByEPwt70zNll+0Yk
z4JWNEAXNgJYA0/89hBYptxtBBun2lUUCPNVe7oIi1xOSrMpP7gk6K6dd3B+gEJi
fQUYme8SeLLXoukID1FDBzBOsfa2FvKyOGJgz3+1nfb5awLdM1pwrSss88EyNiQc
JLrD4EEkB+51uhkBAFp68Hh2L/nDga5oN0zMs3hCz21a31npMvEb5A4D+gegwb8a
FtrCSEsT3XyRbnow4R4zKW9cPIUMLW/ItRG2Uu+pPCxQPxvKieBCzwwygY9S+Rtq
UWlTyXdAkJpQzXLLTLBDTFVif6o2jYkPXm6qNqhI/Lrk/VTsRDqZADIlSeRugz+0
GlNDpfNPdwDZgOfY1LqxwlElVh4ogvQy71pQJ15e7JqzDdIjaMNEoJHWKtqJYjlk
QsNV1bLZyzulce5EV+N1Q2ckZs5u5uUkwTwt173FZLBg49h74CTxmtc2+DD/UhRz
ve2TGqoYB2MWtJGXKRVJum4ROlKpbAQl1VvWy+/hEMFiQbjxCxHvTozEiVKkaGrh
YKYeDg566mPNFBDBSYs/+mkQzSF3PLqV82ImXjdvU6afq0Dv5WIN3RXX69PrDHbp
qvddmeV6PMhrhI1LVK4FzOe+BbwM6sSTXS44FVF+BEK0e+9vpWqrP6upp1xwAGJ2
+U5tJTWA+0fS9loPxqf2xvFjZnNJne9Y4vm1Ph1ESEKZfnvdF+5a6C9h7tM3yE2Z
7YmLFAJ77QnS/1uvk8Q9kX6rgErQK1EyL5rHouF5AS2+D27fiRWPlIhP90TzEzu3
Pdv+J9UJa2qxazLYmpt9xO8V/QCA3/4kg4EMRdXFWqKo8lA5Df22+pguJu7G6Q+g
udAWuG8kzOXitJ5se1LvWJhRHhMPAFNN8FoD43pUvHj9jYDRNexbuXfVKTIuCzlq
WwyGvh2zvV+F2yB/YJAaBtC5Lbk4aIw/5iyeKwaEXbCAAjOK91XMMzbBGS/rO1NL
7F0R8+Dc7H90YS/ifx9BZcaqUVRP5S7m97YRLO4V/V1P9E+WMA71sdYfSi77uVaM
BHkMhkUzOSiZwhBBs4gPk2B8YdUxNe1ZTYIhx6y+WkO0LKCKeLGHN5FcU1PfadaG
Fs7kM9Ys88ZSMpNY8emU8z7sPQJReFjmFErYpMpP5ndYXgsvspT3K0D7bX1X5yeF
j6X1PgMBkuCFAwujYOY1LXma1jEs0h8i+ujSJskZyvBnSuTyd67rHU5JKM+1rjn5
hRqLZMfuTzloqfUb9BRNXYQQ3l5smL2vYX8YkB8GUN7Q8CL2J+KPhfhjFje9wut4
lpVwa1a26Hoj3jfj9KRp9OsZg0+wWYGV/03bru7TxTCPxp/3NssCdPAQsM/td/ev
/zHq3CR9CqgwtyC1Y/BkK0bhYOBGGISZ7dVNLp0D361G8dyu+k4cyiz+jbPSFV2V
CNXvycI5B/oST2HNvZSNwKhDMtBHGkFLD+s81NgmmS+mXfTLvGhZ0NU/jJHzrHmI
G9BIwGK9tOqXvU0xjzfNf6ydnXbua/uv8b4cLTAZdLz0v6Z0AmvoEUNkusAAlDiM
nasF3lSiEaFvDM+CDvp2jTdsfRSnzuTSKEz8ECYdplPShW3m3wtGY+RGwBNwipLD
Rtx4nsUtJZ6ioSjwtsu0jm5kRb+JJV5fDfR3tVRIi9s1pOqt6lzatIAYC9svsyE1
GW52e8GvXsY93GzZcqSK6rTwmhR+qn59HcJh6Ro6SykOA3bHJ0AfZCMoJAnu5AGo
6ZkH1xJc+gEYC2Vv9STWskKa1m2ndsibcBaT92UXNNKqpPbV63SYy1+D4Pqg0tF9
HVqjFpKZXBKv3kRknxoTFf4VkqUQEpkI+9mf5yVmR8PVNI3fui4+netjeb+fEr2a
dG1xipErhr5PEnN9kl3JShKykpUAdGFvA1CQMmS1vrXNJcPpAVDZCW7eWqmHc3nq
61WAp0hRK2AoJOpANfgKFN5/kvF8jeBkxMi9QiOG6AUV8vZaIenfB3HlVhkbMIRm
Q58dCJKxygT5vX7i2Q10eBqXbIUNQ6+fLvWuI4uy6AllScfoACOsS87Hr3IwywHN
b3fNwOJumEVfb30oU61SIV1FA/Fd9h0cbxC13I6BoIC+8W0IwYwEcyigmxyfuzCd
b/zTHtZy4EzSn6BwqMK2qRe1T6szkJqPlo+UThWGRKm3Cf4o3ij8PeIo8bi9EQWU
B1n5UUso3MdaD1GjgofswKSJ4+5vyIJWSuz5CJ73gcWvTWJxr45x3UKbJ0dTWv/k
gzMZUx53FnVwzH3JVRhLiAZU+uIBUJJUf6ySU/0Sv/EaDxRAyKNHId+wWLkeLKti
as1ji7dI35xjMotsZb4/h3k63iL+Bu/vnWCxtvcEg337qnM5BpLDWIALWbXpXPd5
jFtNXC5DUwn+iyVGtUI6cZ02e0XDcdytUZ1igjPYTitihwQJjP/NxD//Q0knryd2
iqx1KOEHabBz6mj+MAX08XvKv9erfXc6XRdAZWwXYbdxCnXeILxmVznX6/VesGLB
WKUtnjYkjQSeGBs7glW9qDS+vymfh4lxJVSIla1d+yBrSivc0zC0sJmrYV6fh3X5
+moEp3WJakjj88IB2AP0KnvH+3cLXTBixNFvg4jNY8RmqqrF3Et841rU3T7b7+hv
yTqLCRL7RI45undfrQgU6DOlHHrrUFNoIv8h7H70SstF57CWrQQwZKhJ5EynTyMZ
q2KwBXexjef3FZkOTzpcHXNfH2Vb2uUKZi7olBpDLymbs6MvA4UoqwSbCRKwY+0a
BXpcarYR5Klk+2QpANty15lLEB8WJdckY7gYul2HOhY0uKx1PQJhrBjudOhg1Kz8
jFFSlAZ6AQTOocB29nYJBb93ePPBMkIb+3+1Qu62/jPhwUBhu4CvATetmLV4fF/y
oGotsbM1KQ0BZvcvEBGQ9MOYFKuwJ/yCXAuqrd3AEx9+iyilOYnAgeQKdBUNIn32
hutofSTsR/rcxet9FKHxFsg/jpQ4CPsMgo2VpnqEot4lxtA7S81vDM1smf61u0TJ
xTlOgEdTH3Y4D73LpOrVAM1C/KRmHOEEzzgxPUl/WBtiqjt6nusIyO6KWO6Hnxqk
kNH4YQPbT8M/zzQ1sBGv4Y5sUANIlflY2KbrEqG+mKQxknQrboOSzXH2HpyDexMf
vLjYSZAt6cLDfVnIxzmQO/XLbdAgvSSMuk8Mk5GIh+SZvCH2LNcUk+gfeSUWnvWr
BXAFlxY6eRoZgbMCGdLabAcK8oYLVIh5Eka1aOyQSD/tyEJmSpak1G6rdzTlGVah
s3scslt3uTMDy2q8gUh1goqZIXNb0v7PpZ8tUxfhMzpSOL5j1SlvddtXlX5EfaI9
OxahmGLywou2GRDlomy6HnYUkKvGjLQwbk6FRNHdyudC91KOw8ex2ExEVbn7Lffi
BYwOKwQPaNL8PNCf9crQiAkrB1Hngh7ZtkZFaPBSiKkfgONKNF+Sodyaoyz6bceI
U/qzJrr9G26HKK591Sw837cn8p76m26PZ5wWgdDeQlGgZ3/nVYttPVffj/syVrYc
QsNu5DqQdau3vhgyEZcRZQC5Hi97ydHwgpN5o3Dvn4rphtbUaEO0DWxRBpUhku+u
B/2xE+gWdoIzc6ofFrXVXekDNHOAXfcjFsDfXT7J1TlyzjRUcC9P7DgpdLeFxMxr
+EndcMzCBiNnSUFim+wkuqfe+Cg/8xODn5kWG+cU5c33zcArItDTIztiD3a2GvNf
d91fSc9V3tHPdtedv1uf6P6N+Ykp18Qq6KnyGS2ffpECX9FREQDE4hE19ODNUZ6F
83C/p0m8cD2tuud0OyKbtpe9j2s06Q5CisL1H3/blQuD+WoOJjRQSb5KXOocaOxX
xFvhZ4l4I1w9dkHluIidclhOdADl0CTn1iTMbCtFxllPqpTobu74Ba3OHhAk0rz3
U0v4bDEUJmXkjnTJOxyiLho/lz+1+TT+BGYUgR/C4JUlbls5ZaRu3z6ckKmIuMKZ
HyHLVBB//dxVwird1IYcm93R6wZOgh7sL6SPA+3iSoBbOF9JF4I03jPxWT7vNGTA
KczYIxqfFJT/aPaevINh5hSNUlD9A/dkN8tE6bYzaXfmaIZOWDvbZ/6M0ITNPHNT
alQ3X7e04kwrHwfhTrWeIQLzfVD+lKoAbvrjGxm8e9g93lSnqxpJBSXLGcI1acUF
xuVvJ1c4UW14rwZU39MJ9f3s0I2HPi0RomNQfifcqMD4ZKCWYCHZ/iOTQwK6znkt
xxnDnzSsPklTx04hvAdS558fGQZ0I3D0NEz7JsY9Kq1bDHqt5Hu0PtVmlxm4fSXi
NkA4teC0+4y1KQEqjAhPPGwUFa2oyI8rLu1zEJY5LHgcLlHYT7Bzd2evw6tMdp68
eZ+Ukob8/0p+3d9sSYB4nULzeuDRHYvBmgwciSyElq/jJXh0h0TSk21eqaW8IxZC
cPCk+ocV6qVFnkTCEHj87ZRNMuUHIQH0DlBRgJmk2ib9DCRMoRXrSL7oWTFxNq46
TyVhSGLzhwXX7zAku/VxYBxFanZ695TKkqlTaDwmicxzTMlbSwYMmrhJvgSRDly+
ckOm6/dm6CmevhferCGo7QH/4/sIHMR9SjsrVTs/YmZ71P+oOpNfwoOd9ZXT61Pg
g3845YZCp0V1BnvfQcey6n620UVglt0q5NRUkgkFKwlRhtbCEfO5vTRQneXFvrHu
XOgz+GJdd5EiJ58f+r5IJ45/ygwQE5Pn2Dfv1NL3AfzCNJtbeVmvDoNmDoG5hj1l
k04HLx7DOgi9iesdNPysFzsjw6HlLc70wqPJKPcKFtlvDFb8wZsuEp1dwSZYnaCK
kjR/qzJNYlwNS6s7IYtGrUmPi4z+92Xk2PkhKu/iafTctkDJH0dghcTLrpM+H9xD
EU+5iYnIPZ/vd64KNjz97Uy1ewIg8n0I4Ws6XMEgtxOeld8MA+FX+Tro+HbVu4Ht
wElIH68/3VE3LE9m+z59Ee+a8llFZJi6rp6F2LC+JxwWYLyXDbF+S6BRMU9wU9DJ
RSCiornxCwGu8yjhr66KT+hfWru+C+0SbwWOP1gEfYLwa6WP7RKIMiKA2w5mhODk
xXaSKi+DPspBZq0B/HpU+zeUrv8Wx4J/I3sAIwmUZ7doKQYGrEa5Fd1cICDBT/47
Z+Tai+UMsndHE0Xhz3Jq/KzWhuRSb6zz28SQW+/64rY2g8b40rjq8mFZgFhH6Iet
DQGQu4/SE9d+/TULM6N+gLnwGvGcMGee6agPnnyQ9wIb7FC89sMuI2cy31mlzaHJ
xPUWoQsA10HVwXrbnBnqJ4n24Vnc///7E6tSVUm6u84o0BSONAGJ7xXTfQ1AyKlm
FSOVwvbYuI9KDEZpyw8kUsSCjXeArONXs266rOHWJALmlwiZnaM+1GuxYtWLjR20
BpVuin4WvC4c5pvFdt3j/ECU+GLggTC1FwJWhWqaVntuL/8Qbr6w0R8nqj/SSQ7K
APxQeXPhLI77c7Td8dHKc9GbQIPfhjrasj52JFmsTZyhTdZywki5UslqVVcxiueT
D1CFf6NXAoH+FfYdSQQYs79axjLtAppiqrtISe2aBl0YQehJkZDRs0qmyyXrKkkZ
Otyz/pFXn04ycZfq/gZSnHB+S21/4SrR4oKWbMQ1y050zfcHq3SStA5QyXTduxZp
1f4uQVWviRvKGmPV4+MRHKVTt+v7SQGgcVpYJO1rO3NMGCTu3wsNpBRzqTKZJd4C
LAL07hV4hnC2hVsfR3n39oCW5V/3FLdcSpESlA/oXKiQB18r/2IB/v9wxmdFzRPH
jVZ9VP0ma7D+EaIdG11nhqz9nQOMbuiK5KaZeEH8lNbC2MpzH5XmhqLUOctWJj24
9fMWpCvgdM/vuR+L40CEgaxqIDhzHMDhTskvTVXdqsera6AiqWRd67DE9NK6r+PJ
2ZJUbp6K5jmFsbxd8fJLnXLQoQ8o6thOfmhNEAVL7uV/G1zl9LjTLRQKzWPnltTd
E7Hq9Vm3J681oV+M9Bbg5wJWazCs8dojh1Ww7LkhSOEEbTJkbcEEMrkOgizxMzOV
oeDQaAXbRV4Ts8ydqHaoX1X0ryU6cCgwTQQEYnPCMf7zA0LSr0x3jqgfuOBqbkWp
3HmM6BYTyPNWezoKiu3xb8FTsYDFvRUQpV32U3AFu8y/1Et2qldH/DokwVV0EpyI
3vWYyvyfePF87sCOP203+mgs8QszTG3acWtB13yjEQ1cBRkMlYCPJthnhEtu0jYt
Jqnw0kRha9Q/eNpSX3ZWxFUSSIeGI/Z9U/fd9lFGBEY519FkEu3qEc2bMluQGlgD
GZvatt23TEX+QEVQ5V6E+pZmPrleC7N6NZJ7ouaA6RV2wN6U9VWZ7dGbUxglw5zc
9aE8LwFwQbBs/iuDzokgDVnWTPgw9xrf+JO76tlUKBrmFJ/YmeZnBRlGlBXbiVaE
FuVILFKeTfADJbLnpZvCrDLgLrWvUFrTsVMqXU7JNkeOg142GZg2AQYHiNGoQPpb
PLDAqiHHUCwlXmfNIqta13Por9HOMBdweFjHP/xQoU/j9JJr0yLy0xG0/pShB06u
VkpYVdfumQg/iExKcogQj0W0ZQ3Xgt3/GjcIv0hAFE3ZQmVlM5mmwSvH+nzJn/s1
2neNeiJ4EFeZk6391QqpH1Ab5img26CY2cAH1u4rur6y78Z2HFy/eVcQe3zs34N6
xI+xAWLCKCqi6o5e4NWkzNiWkW110c2/mDJKsZqyzZ+BD/3tKbbZrQEeLzSrk+Pd
NrjyUuqmoCPHzAW0ETFyRlFL8NNfdk+MLxaiWOC5XYvwevKKagM9VWai0RxGi8Jv
KUrCt6VKNC1aXj3eeP94cSOk5lpOKlDiZIVFcQ3gJnbqzAb9PacfadRfr+i43HDI
WpJL4AfGkw35AjGItO1vVHj3hXpyfmZbHBw3LfL96Ve8f/V6/rSowDkjwQqxNE92
RcblntPdq0uGRIG+SuMjYG1uLcv14BH/cg0szVMB0NJpZmTY+3GLjotR1M+W3cFt
1nMj7EedO47bC34a/I8XIgdcuNvvGOcg+b8tMjTsSE5juRgf5o9f3gecbZwqVL7w
Ns+i2J2kKTMHCEyFMZNTqQiFfSOSUvoPyYre8RUE1B6IXsvwSfj+u8sQKAFxmAH2
W1d5r1onmhKkjHTWeFsBzprxfX2wOADEksj9EhxSYcaLe0ram9EjEakrilX7j4rz
UkJCLMnF266Yfy1Yha2E1s2rOilgM/SFF9s3gXe7MaC5AFhSKg3JYxB9tuA2BU07
eYqoWn9KDK5FZsMi1his2vvxc54/aM1Fvyv3a3G1mftCdNansWmQqS6YvGml3BED
tG/J/1yVDSn0HOlUlNFsY8ZBG/nwOzM+9p8wNDG6bJY6rBsl3w/TozGGzziUOSVV
wepoDE0+2fT3DvniMh1Z/qfvbJhl2/45o5kWpxWHUuoBhNQ41+2euOUUgxeHQ8ye
Yp1b1C2hCinn2ZBfho57ZBASS1rYYV640tn+EEVRWCM/BotFSlBkn1xmui7c1Pto
rJKG3ISShVPFAIDzS3oiaen3y/a8HPc/fTx5l3YLmuyt8WUSLhPnkCjEOsvbKnkx
HHj3Yh6GomwF3TXQbGLyyPu5LMqraBH/TvAxsGdbRj9kSDuNSvBXdicEM2IzivX2
St+O7UeIZtrarDuWIfr82n0ZtXJi2w3hnKvTQtUhU7hmT5QjBSxWMC16DdiNfTz+
AA+QJToyiPcr8LvYhECtugO5uEYlLNx8obJRuhnzIokCSMmwQLCprd/xP50NBQly
2VTiHYvoVukiBxbfJMwQIxGVBdu8eVNnlcgaVA4j35ipJCjECbt7k4NtbR0ta+vn
xDJHp+khvu+iaAK3Oerp1ebK2ZF1CTf+Vu4EqtRHMe7VPoL/QQbtiiyrNqwaSUcX
b41Deh0iXWDqgs6Li6LlwiZNdlfXW7HYls1IS/oygvJ7S7p0Q8A8archRYkSTdZv
L7gnF3lbweqI8IESlyC3YS7eI2/58u0VSp6kTicZB0v6jfDob6nrK0eZVTbgkIi+
dAvTLItRdAXijyh7qkjo7bPZvTVVoJSCa5N7p9FwagkuOzULTMfEXXPsl43r382f
pDbcgnANo6REeHi+T2ONkT6O+Ug23ah1uLCwg+iewoO4amQWy2Dnny1CDZ1Ae4m9
Vze8qkvnnrwZz+cHDonoTZZ6lqj6OZY2JjoPzXwwIUNaErbua7gx2YUAArhpWKgz
jgcqqC4LY+7S5G9G5hTrULWJyAnm7+2XK+J+rT8d+4uq7vA0szoo5LlKHMW6Vi8m
u5BU/KDrIMmu3X3mUxgH6h0Hc644+EfUJswyGbsniR8fQZZoHLiThMKJxJx9JECY
d86/g4AnOUWgIPq/uOh3UMmzxnFDgRii6Q52eUEBIC/MOCmSZHPReDFgK0UDCs/c
iVXsw4vk5MftH3r+zd0uZS4b7DhtxsxeD0OhjB9rTOUHK7UlD6mcvg72UOZY9o7A
ZPG3GsLgsVnNyN0NbWqhRR9SHEumpAeUtBsdgu8bF8S/Jltnxo4VHImTLv1knMgL
817uKYSuL7GdnFSuCKFhpWWRcaNgrOxSLdh058RUwYZd8PZIF9OlVc88OL8W6NlC
rWMHt4WVJikTlz3n4Gvvf37OyLRz159K9s3vY+iu6mLzq0BMNsaISB4vYESFBvVE
OPMsxK4ZwdyP6+aVkfIxzi1xdbrJBO4rIqUWJB95WHwgKDYoGUgueQ05hKxfTXJb
vivplo6U+bJVio0xnbZXyoOULbVAM4YvdhENCm8iZtRCXVfb4qY5HxD1UZzcvh7M
PdCDSitrWfTYVmF0d3uqqFpXuYtNQrGhQHGCAgtfWr+Wn09RiE/x8DR27YbSk2ay
lPqhD7F8QT6JWFO21N6aC/ISBzIYQslTHSW3KHzM7fRzDSYdroCwA3gDDsHUCZ+D
MkxzTEqywWnAqFo8hxyIl/COTAR4TdQI3DfTwKc2wne6m+q1lDWxf8ZA2n38o7IH
Afb2towwkBPHM/LD4pgz186r5w4IFrZYLCa7+KyIMrQ4XCGJ1nPPaU2NU0GBIvX7
pL33pjzvxZwK07dOX3KcvoZGDTSNdMwCn4oYJv+Hn1F6qllg1VDD9OfTT9gll4Xd
+48L2gypMYMm/FlKZaR2iY25wfQ4uxh74C2A5VQaAJi84IjvIvB/mrv6L6GMl7E/
QShJGV5bRJInDxrum85RfnLm69kxcZw1isnMgVVWNokMfz/hswMN5EcM4Ax3SAee
B6Xr/bYb9zMtSjt4nTuPYgIIsXrRkutw+NKW1aOruXK6Z4aEVS0Yb4MaoEDoe9cw
ubXe8aOPJVMX0vGNDSYIsC+lOiWnzoZ6urE8PxLurTZy74DlkCtIM3ix/oTdVYF5
asXB0I+zrCyQohtrg/CdRKhmJBxx6u0DX+swCU1hBbSZK2uMAJFirhGUI+0HV19l
LAOo+sq3YMi810miLH+eXLaOtHDDHZ/h0lpflZ9jCdKcHSOXbDrKbYKO5HUaSsiU
nxjKcMCp102Ssr5zsi+kKJadDW6+jEqRr6AM+ddntNJpmHIqoow/aJCIZ1tNCGvt
pe20QEvQ9l4fLtXR2XqU+9i+NtspqtbIr9IN1q/TqikGXG+pNjyuhGIAdh+GPxqS
GjCBZEa2mBKiQImlkNtpyamqWnVEiZbXBs7mUPKzrYyDQDk/4UHhEswcmFEEBEMm
6mO/26ZTE7/5hl2HYeZpp/mRUZhbNekyns1z7wZM15UrGiaLWkebjngZ3Ltl5C1p
lM+JGDvS3rn08G2HrMYEX60RBOEI00DaoTM3blhDcVduOBK4q7xu7XjH7AohKJgv
BFKtI/dmJe/JB5lZKoA2oC7eMUBI4brZcHBmwStSgZUYgciw7P9zDKh7wyHjtpvh
5q/Xj4Y/iz6q8DAjcMO2NyIvpsP5rGZVjI6TogzCqfqAEBTDZEpg1lfhGVqftizB
V1ztC8zw5jdUe5lmQ5f1T9NczoADfl2MKtq/NW4M+4nTO+8XSt6VbEPurWtEu2VU
R3e/+xPQbZOO5mketebBt7+qgzmoun3rmRrejK4zTI6okz2MVHu9R1s6RwXbht+v
0SrUzbAmyXY/kI8fc7QqyTcbqHwUxpcjU57SO6Ula3s49eGRZhHBSEqdoWgFffxS
jqFXXXJq/fAn8PEH6m49t9a7woBz69VTv818MRvYz8z03uThpQDVHygnmCRvyycm
reM9nAKtYOhYCvug1b9TClX4fOaSup0xEpoIuAAjz2azAwXAGqrhZEqt9x2AC20E
hpj26slNU/QfRI+9L4j9jUJj7bHjYgyjJrBoR1QBemNYh1QdaVd5OCF9t+pNpTxE
ZE2UOuqGBp60iZbXBuutcJ16VvqU8QLdSP3PQlCnCevj26KkeV9QaxfhkvCwscRn
QSJXLN1BSmjX8zAownRC2cMWvruqORRxbv2vWA8oAwo0+XvKoxBwNrrcomLEouJs
L0SChzDd5pp/l0J8g7V35wBKaKf8v9HKimz44FxmGf2YF6SpvspX7ttzlSD0i8Wk
RNjkddvS2g3rlLxK6Lgk98Gb7AtK32JgeNe7nJpL7pD9t7LaFEC+oNRmHgGzjxRT
RcO82TfTOGFtiEQuwt2TwT8xnrbN9ea86K/0ALrCgtgTX8QBD/Hk+7IuI/zgxvYe
2Vsn5r3XHJTRIgftGroVrngpwCXqjLEA0zcarY6m5PddoO1/55xttQAdZ/g682//
OivGhP4MNUXo0DcvLQ1Qh8ifDmrFQ8dou/zjfAruBaaeVmShhgyhorvLgWYquCJX
DIl6aYW0lwQEZqzH48+FcHK1zLLjaOItrdwMEaSb1OJw6kZsGzjAepQ4HkIYzDT6
C4iN/Rgxnaad2nKG2hPYXpzOr+aK9Esu/FgsEnWE5oyEA7RqqTnNkHhzMELxY+IX
uFtSN0tn9f4hdXGeZTtFKv9ILexnxvxSlSJRkdFkxNG7R3GezcMa40vXPgs316r+
Fo4YYd30P55H6mnr49TlFMBmrB3RPmKGbW9gmBLmrT+1T0GDzH9QD0UEYegF08PD
/lOilXVPGK2ddf7fMCTcFT8ZiKtgKOtL6+xsH785nbIr6YyM5nHzuS7N732opAT+
TRwrV5Ckdw2Ru//CsGFloFFPTIiyKdBXK8R5EyTQKNvWqTRir1nF7VBA07xL06nc
xHWHMcqjjtgxzxaSUkimSg/Bt4D/IQZt50phZ+om+uRGEH0MYpoRjisizkp/xupb
HjgHOBLg8FbXLfffnePDhIU4Jpuw4Fy6q74P4boATxazcq6+tqmQhbMoQuj6AmbV
GkfNanoTmrOW4Ug+fGXOfZeQ5PorGNX4J5uxRl3NxU1gSww2fWT6OchqrnREZxFk
jAnJdXuM8wavL2drHz4h6mgth3aZ1xaVBRoPyZR7Au9/aWjAG0pUUTAQRkaTALI8
D7edGjWf/heQOCyZ6B6zZFxUogTMWrCh4Q15ovuFxHvGNia1krKRZzrQX/ZgSra/
//BrsTCZBIYnlSKsF4cijyqaey5cdOeU+2mBw13mC52a0IxLwBmql9MVph/tYEIH
qCz2+QDZ17oiCDBBDomLNAdATS/jXIQF0NukTD+yXCH7MH02SFbtgtkO7J3+rcic
cARfr6V+3+mxcfmtKY/DktbEdG123nTQIQkPo3HxtAGaIx1V+7vgEB6W6vwLdpp7
lPNMe1UhaPvPB/FDCvOsGZYUz9qmbr0j8XmxyACgEahL5SUn9asfGRg1H55aQcOh
J8/9fXw3ppg5d6SeGKp+cYf8ZxEUlwrsfcXDKEvDPnc7OfERprGPAwMYV+tawyOV
ZJUif2TT0MzMjD341Ec2ow+8/kq/4Q/W8h49dDy/yhonKP60xCY4eSZ6Yi8htJzO
3bu36WjPUROorw6Cz2zbw0oWWJGLfNbI88gP38tM0TULiIBnDZiNUKnah3jnw4U2
MawPk4KHjyzEbtRi7LEi9V1RXQQsC4Me5vtWxkjbMoN2asLGWWMFj/oZlh8TUAsf
612maTZE/7CXGneQenDPf2s3rjibMCn2dT8MYNOmYeBBkULxe4NEXtMFYYA86Rh+
Nqm7EJ50jBBWOCNzAoIJFF4PdzG38b40edac2U45nxXie1UgW1MeBFyh0eXGSmFq
qs8tmQ3DJvnRcVyuJlKIjY2SWHiEdaEtZ0wFEBHfiQ/HJA1ofs9CWvwJiK/tHhue
NVSp9kYBOtByQgPjwzE3vSRJznXFumi+jY/CuiGkwQUriAbWNmC3qPjuSchteO7W
S73gdmJn7VbaLiQdQ3uSMIsLyqcBEcmgABoS4Q5fIDkEFlbbOxQ/FXL0bBuyC82X
rkpZyI9ez01RCP24XfqQzv9tgT6Rda/rpbI1HEpI3BCFPXqD+bVzkWmK1ZpUTRBu
pKZNXuvj27UBelgt2MgepEN9fLqZtw0u7li2pkXOPcPo1UGSSTKmhYLnd+xM2gSc
YQjYNvUvCI3cl0iIq+KAQFn6wbXIeQ92ls/LDtuyEHJBr7BN0yoCfQ1p7NDtJd6N
ryS8+HEJk+5zGiedG9Y5dnGZdhTHWZ1S+Rthub85X6wnV2zrlcCtJriZ1VXReluo
SGdNECWNTbKju6EzYuQb/kqrp/ZzBG4GrEU1JCeN8gU6jscT7y4ys0xE3oW/yfh3
7z/yWdDcbQ/cGfqGKE+5YESIrSLFcx84ClTnQgj5Xuo/cPhyUJEpL77E2JUwg7T0
hiVc7d1aEZRfjfwQKImOg0D9pbDXvl4K5rSbOOxrMMZSWw6WspFaUjhNyphZfwCb
ndsk0YCfAXQLXF/SBPUlhljE0ev8C1d2Ln9tRdqF7OLHwLMhJEsx6A7vlIcEwucE
wtH1/Jx5aFJyKhvHk6byA52Bj0iVEzM2bSWxM7KUzQBDZcbt7NbxuF6nHFKSXuSl
TexV+gODAejXqwPjBA5AgLY8IRFm0vju/UAhez83Ex0v/KeIGpPWpwtTHY95oeZu
aAtKJPJjw0F4h5RQQncXLCnTsqsIW+qAom8p4wYjHRlZqqT8wQlnYUHSUTYGzcvB
Umh1vnJlQdmIU1OyzjLMTNQVRUB0vNfZlWkrY1pbZbDgO5dQmPck0mMbuzfsciSR
lPq0uQBV6NwEby6B+F1XQ1v27MbBKOj9AxjDzqdagrPsNQWT6u9XtBcsKET2vz0y
SSvmmKDGzcLjQL9cN2/Uej+9bHNKjIXRGPFu+9LLCXEkGrpKGk3N0kvxDj9AjiPi
nQHurGhS0z/A9QpVVvP4R55yHQAHaS5Fks6GQJWxifKeMoKK8NBvhlJTyuTdkS7r
mbUkj7G1Y3vsCVD31VZ4vy9m38C4XZ+VODPP5dIuG1YbeyOsEj/rz6mdBZan/+eZ
Zg7hPDUms2Teej3S0gBNPRpLbREtLMjTyhk49AzNw0YAW41OjnmpmOEYx78Gb2jQ
NsdJ+OvgjOOlub8VAkRBBxOmUwNiqfrp66P89wzrpB8xYgOsyS7B70Zs4GoHZoUZ
DNF1R5w66uMzvpJYx7ebU4mpIMOul4Od/lL2VZnn+JarNJvHmpSVmwJU5sxwHF3l
+zHqkowMqqzFIx19tllRbG4PnsWQEINBrkpbcDicfVOTiqQgMOpyV+MwM5335S06
4yzDIedxZULk3w6+lTOJFJJetxV2l9nNbeu4MRynVonV4ufuSd8sZpZNjrdA9ksZ
QyRRfSBo+LM0JMUAzNTOVpjRM8HM0VFMWA7l5wL8dWZpG5MbiMxkhvcnvFZHsUam
B+SzfnQ2X3dgkm3THptBpDoCnlk+ACyRCGdfh8Ot5jvdQqHXfXgN8IfCNOR3MReK
yGIR5REOX8tPUoeWaOz5tcugBQLXMXNNoVgexzfccS2ZlmTis+eZ1MT5H+OX6yz6
iOAdcon6Jb0Gpb9api8A0zcl+G5MWb/B57mbnaf0vAtTpOTgviXu0j2oL6kIPtSD
C3Nh0Q1dpOS36nqMH2wA+BJUnvdqjyqUXj+q9+GtKW9I5f2dKaDn2Rtf4S8/HhH+
HuoDtcvUfuQBzkYE5ZtWOc47EcPwXxd28cbVuJncTeTYE7UUVgWzRExufVE97ENP
wd2fsWYvuW7gbmirJ0Is1Xu+RwjpGFnaMJdkKyUVYezwk8I5d1HQLr5GtQeW07lZ
nmAqG9U4HlRJCgCpPMpTqdmzvyi6+FxcCDNHmaqMhTYm9wOjC9yZ33Jl4CO9OULG
4TlhVPzCV5Cjw+foMH5WB5fAkfMHlmp9GmHkv22nC1oUhW9rZq20wlTfQ7wTvVLU
oIRlYQNIZKXIjVd5R7ttotCVW77BUU0s2eBFcIJTtd4Ak62zESloYs6B14TPM6CF
8yfDdhb3mDb3Kh6fdJgKPN2e2G661SwV5Aqc5RlEXOwZ4DixdXsyez5xggs1+DFK
qbz7yLpschsk5R9LibnVNLrOHbY+a7X+Yg/wNkgpRUezy8v6lbh1dz5XZVqidusy
hmdIp/7DsPd4NgalPbfhYdHyc7QCBmqutFSVZGUtMEVmEUrTiDb08Ws8paEU4HEV
2MG2oVUxCotZWAYmDXnHbd5AedvcsuQet24lwawkQMOxy5IPoArvSfNUncYAV7FZ
y0S5yk1dEdxFNd2gdx8hhfuBtcp3kKq+lt6XtXFzKU1mGhmZi9g9kq2Dr2cV3Eh+
rhLnemwMf9aWL62kD+XFLLkzi4QUkPPKBw3kYI9Lpt/cjbXrm+g2H7plKq3CngZ6
ocxK0P/9+6gOvZxkumB1lyljxqv146zEy17vJtHy6l+Kh7aBUVyViMNZaqXq3vAG
Dxfbvju3zC00T8EC1hrwdr/UEe4y0AHExA8mjZw6AZ3DUYISMVPrC2lEvS9N5LYV
WDVB+Qj/O/YKf7FdGJIv2ad32umVs4eDOj/aabbfOES/SOvT2+NMNe4pNafpr+jH
i7gGTvXdTxTQwZOfKxv4NIZGtxpxx5/0Q4SISYJtbNkXT7dYcZChALq0PO1WM5B9
8IpHfVZyIjnO3kq/0I39Bdr419DxuwrGjSsiT6v7kZBRSjpJMUoDEiAtu1IEPrk/
zD48AyTl46pV64IzU/MOCHY49Z1jlRHcp/ecMFaAUcCfJF/Pbse9lwbvv69nNbXJ
Rw5grqj2553YE0Y5ploXWlo8tg2qqn5HMVXJzMzM7xZpx50g824ThiD0HtSNE+A/
gtEp5aWBQ1nnoZ7gxSQQYuBpY5N6PRekUjCO5mw2WwS3RkZxXYHU6hJKIvgp65LP
yT64W1lfmB9ItBVn81ppMFko0tmMUaoSRqGc0ACQ1q+82q7ihg9PHI493ACzuvyB
D14zH8mdSmDYhcWwcpA4ds/5QBmU8g5nZpTnYtD/7c6YkkiAQnIfQAxdN80wKlT/
dOSUsgQauRdtOfqHaC3mRNEel9I1K/jlDxpp85pnUp7oC/8yYrjHs4EYWL1roGFf
7eZWBsNODwKE15x2xWBAKnIrE3VZgK0EBLo+P1BUgyOgu0+NpRCLJbOMM4Gvf5RX
TKKwMmGuCSmIYKxZtGE1S6t/ZZPSjZWTKFKufk1wHXXXgPc3ArghuhfqhfTurKKM
LhPDRoeGE47Eow7yJErjfHU6ZBDWRQEqPX7hmnk4un51YlljFboiP3/Kz6tiB8BD
UTkHJSXE0eT3HV7GZMTx6sLJd25CRPJhsTL+rLA6soZdV9gvx04olSovURQD37ll
ppray5cO/HJpj3Up63Dao799DC2avIcYDnNr9gaTKTZAbISID+YqX7bjNWXnXbB+
p+jPXAQgNVKEP2gtzY9VZChwdZOHxO276+cznnwbsd/QLgbUwI1SJJgfAP1+9XvY
wB5Yh8fSDu6bZXTtGmXeubPwqqK2v30IHpH/awoY8lfO/H5uR7uc2U/lO4au5u0a
qo8uldczyRpoeIB9MnodyASqJS+0eBys5DdFoiha6oMuG+gSyYyRGUqoZHxu+Tpv
hfhQpDFdwLpE+bRUQTeyhr/qqyDdcGeV4c4chQ5+wb2cUygTeNhC874wYhMLFETo
o7G+RyFBGGRD2dLgDLvaaJm1q1jTGaMA7WAKiuYQ9PjC5g1O9OVECQBm3I9bv9+s
grmfCQlSMMp3Ze0sZfAJyLh1FRgbgGCjnqBwpJ5UIcq+4s5GLxf9FLLwSvtCmTeA
f48PJatAPP/fuLmtWDYeEo+yQPhwSRJT7aTUsG08iC6U0+KPd3BwMEQKlF0/+kPz
Dy7UCV0F8KJXij6tMSLBO+744DTOw0o1nGRE8dVploWpm1ohk8SLlk09BGcjvQki
ThO4jstWmOtFGjGXa1npnoWQv4OcYEQKGdE/Oe4ECBWPK8By29bNyJbtNYIDBh3D
dmE9HvuSluGdAtuZFFTN7D9HLFsj/nFnUjNFJAila7KJg5S3/VG07QTpX+IHCM9a
e5mXoX+/Nul9hQcWShvgTfiTsKX4569755CuU2ptvvCvbmExhTsF7YqkefWhw6N3
cWC68pzW/sMnLdNkFVo6aZCjyQ7qO3y5ENOG8f2x11/uDwlz5BF6WDHM3D7eK+MZ
oEp37tuHG5O+MI4bdXG3gQ4iAq9FJwCnsCKfq9G8RSehztj2UAbt+3jEpJo2/GNr
+J/vLydErO5k7WNP+WW3oqIsYHZ2QzNlwelmZ/gJ9nfoDRrwNkLIpXZXI1rSpmkq
C7vW/3PwFrNSsRpAgI9YPMBdugMRaoEOzh4Ow/PD8LwLLG2WCc8xQoR/hIoxZ0Pt
iBAMj0K610WoI5FG820YvGuAQTnv2sFlVGY/kSakvgxKmx/39IQJ+sQd1d6aSUoX
JAhAc4hegxNR6fKwRyXISs5nWyRFyVXAJT0+h61RCJwgN0qr+Q78OAj5q8Xfrtlj
+YbAz+ISI52lh5dcF6KHmgiYYUDnCHinNIJwc+TVgqhPhvtQC1vhgly/VeAIF40v
y2D7RvvRBywOeXLxS9v40ywym55cZHH2/13y7NvTPSZE6OUHpK4xsdD4OkzbcZ5A
dN15NJ1WAiKBrZI+evqLKr/5Kgr9dXZF0VNMHBvNdc59Zo0ioVF6DbgTzBB3Ys93
RDSsCs2Q988H6Zo8FU38+oIpaAwiQPB2bop3hTiBMqrp6cksIqctoIBUyD+gZAag
ida0Wj8ejJW4tiCXIPVu55k8ZDIEgblwFJgO6R57X3LkPTV4rvBUizSyb+12qxYR
DM4WQL4eaE9FXcgdwiDLAQ==
`protect end_protected