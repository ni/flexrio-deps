`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14192 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRvp3o8+RItkxKTewZIo7szbhVt+X2UhePTL3ONuIIS6B
jS4QTIDES1AAvoCrVfQXjH/RAVW4q81cCPWznEhaUUNEa/sFuNrFRae0h7FffBzX
RUch+C5EskNektRcixlp39svVqE/rLFNHC+eCm9cPbUMIyMqtGqIX0OvfSF175Ko
HjF7yrXs/PQj8A5rLPW2FPKbB6GmQZk3M7FKncgi8DmAuDArhW07UeymrNYudH8T
6iQ2USvmovAP5/2F5XmTqqpxw59SS4NPSZz1+bDL7NnKWoibn60M7GT3j4A6sLyf
ZHzZQbRyTGPBbV4ELivNycviEvjmcht2xlXD5UuXh8P6UFZwmL8uIDAxvb9Xelj/
dbWYVRPOeT0uNzIVGqzoFZZ19NQCmzkjMA4u9YhRccXZEVeLOJk+3UdfOkmLqZKD
tjP7GDtk+w+mcvfH9ESDZpURuc/BW0waK8i9JD3gQ89V+Xc9oT4UNkNDNnWl+Xu0
qhjiXmeCv4ZwIgMUnj9gyGd1pUgbPCW0stU7cuoLcelFTD8jKMzYS20bNJBADaam
GWAnOh+PmlYsMuwcHRVC7oXbYX/S/JgcIan6JWUBTuW5SC2UqGCZjW3QW131qive
s1K/SsrEEwmVmnYBUuFIsEy0WgXKT+5MhdudDm+H25L/mvGtgmML6ck5dgSJIIhO
RbroVr4OUg8oTkF9VFXLvlo1kcbBmoHp4bJP35JfgSA6oO5z09ugnS/oaAfKRUy3
9EnAr/1hmFhA5KQAG1IeYna2NCukxbgdMom7/tF7ws68qIpYJtHXIvgJZN2YSI3j
YDHJ6ccoPOozJ21yT9ioAwKxvvze9jH0vVNZJu/UigVpBkk0h9obKzyyZften5aI
yLCSkk8oODYq0iotszfxmXYmPcloixEPzqEh1cJy1p+u+zppqpDZXKfIZet4/zLW
SiI67trpXdZGGBRSJR0gQUt5Ie5aUJqmrwJ4BEY64jyoefNvBSKo8jjoWYV/+h7N
lQQY56q0NCKnyKV0fsx++CCElJtjvyTZK9gNMoBIzTdzplFvKeZ3X8+a8XpQGjDG
ISrLZhlByTexfEW2BO0l38yfIfOh8poImhM0d79pJn0iDfWCq4DJ8n6yx52DBouz
QtVihXkzLhHtoBwW5RUfzVl9rGOy0JImZ1id0ZPR7a4/AuVue8hiux1Jm5VgdgPv
ZMrI8pQBkdY3xHUJNav+VfHeEYFHbaLju8SjiQMxq0ac/McqSVL1PrXDePIzGxvj
BQvX5FD1NGYI8myBYdCSa1v/Y18GwGvdxTYm03MToGB9iKVXHCksGcA1FWf6h38Z
c5RkG0v6HgT6Qvfc3QQB0GBds9ftBfdrYLv8gxokYMzYQ2adpEdoffLk5bdsshgi
+iXY2QlqgGT/WSJI8tAKZgFFG/ZgFG41WqRaNQRTxc2Ghh48LZDmJVgzn+Yn46Od
Es/gzZ3vU+HtXeQeV1N0XruJJ+/P9jDUHgP4MVDbVwIq3qRfEeDJ/9aRz23PqjKd
5dMc3ajf4V/+1JOrMv09FQlRyKqB1p7tGm1oz5av+ASbgQu8mCgLo8W8Q+YpUTh7
6uUz+R70y13IIIgn/rahAFdH2lw2qwfhwnUL7xGQJLAde/3A8X/ooJL2nKTWA2Qr
P6Mk42eHS9Opcq6Iu8insk40LFCq7ebMoCOMcZHTBGagMWAlus4ABIsR3WJulxqa
OQql2YhHgxLrG7tMqtY/yAsj5upaBsMBJOvF+0eqbfqlei+tJaFwyOt5BN1O5l3g
mfhJrouCxgnkkUF3ftRpdcn2XQXGmRakDuwKqx5Dd13yzzxPGj8z2R5jJz3T91SE
UedsQ4CEFX/pO05RBo0hdc4wuk1Z2iIKHGfw3XxXDwf1DNXSmfnxQqKANbYZHwkC
D4lqJ8FNnSEqeIC7QZyeao8pakOx+itcDwd59uWixWDwJAPxFL/ft9asCNDY4nDr
OtpFCbM2Fo8eeVe1GhUykN8sdedqHNNdHDrDiz//YVONNKD1JHMAedkhNXwLpfx7
BjRRGIKyZRXb/SeDSDiRFQXjrVLHimB6HI4x6ltfcnjvKbfz6WsiYGxSJboSZDA8
bVel6k/51DQxZYseUlkFBHVQcxSYcQHV6E7VQDFs0k4mZFu+vfYZCZqqRY+Rqrz+
YyxRiHW1NbU0gJR5SuyBMlxwNpwaBasKA8gujd8YBi1RYIHeOczy0gVtUU/SL1DX
W3D69tEFHPfAT1lZCQxRyP9cbERR3hYNPpkoeXervH1kFiqoE8Ax//PFH6aVh724
bxHLq+m/YwIwSBkLkLykghqcMntkO7Fr/+e3uhTiR8+lRhyXDxw7y6k8uNhtkPIT
jw/JHF2Rtd/iCAH3Uxh06EegZ4duUc31y6EztMYjnz9ElcinoOXNQqyylaOnhZLc
GNgjpnfvVlmV911h0wFnG9bZQlDUHFuw5hkMB8vw9o/AaW9CvQLt+KsLyhW9deWc
kcVTAEWg5tDqQXf8xdfISetgt+jDO42vVtp8nxhlfR5ofGagMxrO5YtJ6qSFgzGy
gO720jGmzHJfvs5InI3jSmc333C9D1ltxY4/XzhBr87T8w64BxYK8nt6bjLd+K3s
9X6zwZc5xuQ7gTri5loy+I1BP2gKlH9MbqpiHAj6mBLRLgaaSaQZODGBgaOkQvHP
ReMZCTByH+meu3Ig2PFqC3zWjB6f9dHwovLXzqF9J+gfIgDWuFy9mw01qgLFAd/g
WJ7w6lUpllbj2OGegm8tF8EFpj0mGLk4ncwLo3C00A0UBZzEHVN0TCD76FMVVSiv
pKCJM4IMiH+vmrIULHmae9xMfRnr3v4hv5he9vZKzNfhTGQkxNlBU88Qk5cn+WYM
blI9WP1W/eaFobKXqQ3s5bHkfmpUd701aEtoL090TUjVPNdpRD7aKeZ3POAUZuho
oJMdGWiwCsupxWnMOdNlh3O7r78IkNGKgVzjjdvlSGCel2czjCqHZR3hVDneEgCr
VW99HctQCg/Sje4AZwhABottDFm2uc6jFGMe8mkf6AlZosbe0l0+4rWPva6k7VGx
naYzw84s++9JXeNIB0R5z1hbOO8MNaK3ey/E5pLt6ImqnvQ/V9IcgeCfDqkDT4Yf
DwcfyKRMrVas2If/44UzGfmZmo//biEaaQFdMXkVWANt/HaajjhmQUqR5tPoTUMI
rhUE0WDNKJWQ0DxRWrvVPBYIv6wszTNjZmspqFng4iyMNy8E2S0oREM6aCWT8q1d
O0D/qiKiaWsAoo3tfULr7QZ1YvSeoTryS5P/unOJj57NNb4UXD/egqRk+P/RVkgy
bOsj7Fl5qukYDjiauzFsUqtIPdt9KrFYFP/UlOPaJB/uMi5XRDyyY+Vw7JjEsqjR
/Xfw4ZZQZK/GJIGu6D/dJfVwPe6wrSxfmy3FKDXkGnKqYqXXfKeZYUl6TD4nvXqV
ftJNp2eJJtiGUPkX/gNB7VnDQ70MNbym6od0X6K9s/L4U92ZgahJ8Vn6SN4XozaT
DLqMZNsMdnjeTDQjD6uN8BLs4Oq6coVNVpXLL9ziadMMGFY2Hwb98v4LRech037w
mtg6Ki4zoRp7R61PSAhFuXZdzNfaEFYB/rgDj/D6iiGuKQRUOEu0s7x7cPViVF/q
zP+WFosy/qYgvX5SVo/8nPp+wYOJxQZ50QYii5SaAAFG7K3bqkuI9e/svgrtGuV5
11LKNx6+K8i8FP3DZw5NG+R47/vtSlmFbB9Nt+iavLYMc9GzQVlNDAapIL1dGxxx
Bzryu71rBRYSOIPVcchBNPdDYPazzirSP/CJm9HyGfeBM7vRJ2KSgjIfSz424tjx
kBNQLocsLsA0K4i8AVhJjO8tmvwAA7fl0sqz0Fgrcmbn41Sk1t6+QDpaZRBGcupB
m7UQrSF/+PH8wfjn5iHDJ8KZlVE5Upf0tMEOqnb6h+T5FqCp6Vmw9Gn77GD6FliV
CptNxzPWiglucsGN+JM6OB6uvyZ1psz/opU9UWDa7XhuKNPSxUvPTQv3DWdamxY8
1Y2xKtUKdPjD2gXFKnTVxGuPcrsg+TI6fLnYGhNevf7t79nwxhy2vWuhg88a307X
+aYktDqrLOLEWd9FpZLjwQ/RlqmmGRilI3N7GsT5BkvoJtedk9E1G+J7o/lQln5o
fhmAp+f5EDlsQrWdT9p589EzJQYIHzwOPsugefyy5ryUCk0LKe0691cngFV0wn0G
ui71Bh7rGPrmUmNu/O02Y5PlkDogDyIIb2J+hLnadtYQqWmIdEoOz+pAEizTh7YF
Vb2I/USm16+rfPmsYNGg+nV36CfQnGrqczLQIeluCc63nQ2bp7xW8/++gLZG62/8
Psp+Y5PJAMKPGnyBnySUpLAipq+/0u9SojSVqawHdengVkH7W3YDYEsfptTIMNKG
ESaHx+FB/4MfyRGBk+2hcfJFayRwcH4WGoSdKIgbdUvYwfbca9WYuHkhLoSOp4er
lKixB6WQgHllqJVcVSkYT2ZsbFlU2aMOHJgpVBXs0PpQiYRjLS1qYkv0UYPDvD8t
Bqg97dr0LRXZhzNvj1yYtILnuX9cnLPatP8A2HuPA8F1FJSVHPyAEAxNIRD2X6V9
hoAE3keEFN3GSy2krDcAH1z6QBNzhO8yKeM6rMiyiUYCpIu7cgUGUCUDZL2Rixr9
1ExRpEBc+rI8AQmOK+kPHpz+SO9dhOQPm7zAgAws8UPTBC47aUhxf0Z8EhsFZeAI
AF/WrFyg+vVbA/x0X+uswjwf+cohLSuRa+3dGEEKxwFVz/+FN2RJ4fA+NutmXHUM
ycGTdpPgzmsIU0KjkFE0HoaF2ZBeFy72aQJZmfroiqViRZ8BgO75U9PP6v0u//bm
oUEepu0/QhmuXyaRFpjS1c447vCW/SbjmVf318yQdYeOEEvgXKgQu06IM5+xyz3G
46mHNzblbtfPSnvWdC5F2mEKagXVV1LMtyD/zNvbwpRzlqEqk3p8q4f1z/hvg7J9
D1Ip0CcIj6OWHdAn0RQhCfN4sJODTlSxINTtXyg9+7IiI0J0f5ZOI2+PLlkRNHpa
/jspR5e5TmbYGeghaN3nwvulUpIFkZbrjI0lCy0HdMdcUCGBGnvW1uL6VMExNsfZ
nBIEgoAAlbEQ19sb2rVyjSJ0mjo7HmSq06kUYtT0514eRYryZsQD+5V2jocJJmX8
XwxjOS4HSnfL8gEFKp7bWwNBJMXFgv9IGXNsLPYNexplOL1uCMrPsaVydX4FtfIi
QorSB2vBet1cEmbCso/vGjpmNpkm6TN2VqnChf+fAgsc64mI6a20qLV0bwwN2mx4
ITbh9OtF+1GsZxRn6hl7k9UNHTKEjosTa73PjWrywJUb7FdzwkRYDhix8kY3k0rx
aX5CIIExNqjauub1q+OMsz3zatchX4QbgDFvm27YHsEI9N9JubuPXwazWQlM3f3i
K7O9p3DfP3g7OPXn5Voxkq+kAb+X8fFBr5RVaW+DacuQkzBnnUDdPvxsNDwM/KvI
7/425LvYX/7AID6VHuooo+pDlFI4OVu2Nnxm9p8fO8cAqXPTfQzcLeZerdEGg4oA
TzOREc76Qoil9bZ5B+kmxGZYbAGvxeH5oTPlw0OzSO7ssCpWS+/MGT7A/UHd/w3U
jIi2eC1a+koPPxXtafrGLMEawkcSWMPC3NCGpcc/egT3beLdZreheJXMoaBRTbZ/
yylqPSExGTmxwfTFuEcw0FFv7jB4QXa7oMJMTU5QBkQI4tQe20Jl/8RMuEh6iUdj
bnwpphMP4eWg6FG5PW5pY+ekxtB9iQhLeCXAlfvgnrhu1bUScTg6EbNL1O55jd1U
2vkHrUPNYdDcbUlEC3ru3l7Zzp8vGoT/rjSshbb1Dj9LuaG79TyUHUhas2cycn7g
aSKIOt+Rhp9r0PsvxxerNW8cap9eC5+neIs8ZS1WlulZ7JeOfkhnfU2AFXLnrtyr
unqH0jOPyxxZ27i0x8KsEhr2IhGUHRLepj6JkrAzGALQxbXIbx9iAVPuRMvBTyhc
i/l0XlGmFawnr9kautt/QkU7gb6DvAT6g5t1cOah8BLd1tDX+KV8EQxDnutbbps3
Dzx21mbsdxpMQGAmgoYkqMV5HUhDygrEVFMpKA8Cm2KvmzqtsvD7hd8fb7hEYoX+
9ZwuvKOvt0Rnz2z8mmqZQumMZGkNn1MtHbLJnBLRpbVFxUdoBNviPkBqGlCwn5L6
7Fd+gaJDkNJ4mMRjOTYDrUsDVtWsqQS9KKllomnglwIBvU05D6hSJHCd4XwjWwJN
yNDwnt7otO2VmDkprMjcvePmZw4yiunQcMSNTTLcknWMB4+mCsbSu81BiGtRDmxj
4m6yTCz0UUWuHp40tHXTeGYPXHA6yJQBEyR9+mlPofA77qgtPIHhJJ0LPxQ8BwxY
fSv+OG9kiUmGrlNTvlbF96tUyZPOr2zhpRji+G3b12swVrVgPSf5a1BK0sq4uWzm
I3yb7zeacuTT4xOPpM1giyBH6LcYZkILRgp8tnvF7opgGxJdMCJvUjaXXIjkCKos
+VMgU5Gwy9iaCzavAau1rFm2/cy8yaut37f8hQB8S7YNS7C+cs3BqkWyOr8pHlk0
2/x2lukP4AO93IAaJmggumxHDPU2F1c6UbZe94CO/u1+cu1UHnQMx8xBoKooxGqr
f6FDwxQfsapimRFk2sLIVkya1DyRBH+56te8lKatr9ZIvq48Hs71w0sSO3DEQkv0
RIIzGn0r6nFvtGq+RC+82TMUb+B82kyvb2rcT5rwU9y01TMQSuCF/6L94onCQjfu
WkDj5migtK/n0avaqwF8ZBMDHhPYNVijlng4L1anBijCcU7gkNTLYYVJKZ/qTboF
XBlEgN6HC9ghIstmbCjnGm0vC4LUTGN9lMv1RN4bA9a9iZeYzJOgpd1h+pvBGqwd
rWZQy4ac4VT848uR1YCoAEKy6DJrJiSUqC5/958BrEKTH8Peo796yD2awolqq2pq
OkwMVu2dqAtih9roT0WPP8a/l7Z0dB/wY5HAjO/P4025yFG2jUimGB41Vjro6/b3
7fLSKvRI1uKciFsng40V1H/n35pzHXQY5xbZdoQtfag0pVVPj/kRTRlQ44TfZjEN
6fZNfnEVHLOpdINHsscYF/Z0jkfUjuYhV0ZI2l/22Gvx8flhSIJseNjF559aCJMd
3iXmrbQuOde5METdh0x5f8bSgNtLGje418quPN29J7Eo3n8m8YtiBFlDLinVKJ1p
KCPUGuBT+hBMbtgZfgI2d8uRa7f6HeVoWT719Khtwp9CAKPyWPhxIi8gSjo2e+7U
JEM7W46XjTu9G5/LJzsx0tKhgR6cCbukXOdhpWr4Q19yxx0Ed4ZnQcyMZ0KS6wOF
pT9ljeXs7gNY/ODHV2NuuWKKkoSc6uBL3D5YXRq3fLfiL/V86V9aHlvcoUEltO39
Lcz9L20q+uwn2BqvgHXYNxTUAGInxCIM09BhlN14RyubnhFyRFeOFsvsdsYXVCxj
yXbn+YbkTjFPoRV29eN5/CODXVEiUUPbbyM7rJHq7m13FM5uvzHFAa/B1ES87RZN
MSFs31+otwJlH+bA5489mzZCEnLqVfRw8fvFu/tmMGizeGFFn3Scv4HlE2FgbRt0
PONxOcShBTbsAVnGZi4lgke47lyHEP74F+e/LkLAVeISGhgRP9whtTMr4QHTxTAj
qikyV62VED7IhGm0aZQJT8o/ORl0arrqvpVoXNCF7qKqiLILU41qWGko3J4JFfuo
swroUtXLXWBsL+rRF26iIL9a4Lflk5lcvMwnbD2xey1rzIXrdF2a4X688SksPfCX
8sG6btqsMqj6QyJSHaCCEmc+t6CTpqC7+BY4/jDmF/EX5Nl/zXnM8DF2Oy/3A6CA
7kuu5MkmYHVQZvtvd0cA2WqOo4KBM+vEkcrY1wgPz2KB/SrLKH/MDEnD9oyamVbM
a5NfqRsOCN2jAE3dF42hv/Dfd0anJ77ijIrZMUWhxQVnBSmmVeDop3JBtlqotxzj
/fyJ1tNm8o1yd+/Q2scpB/aHuClC/GBGr9NabLF85vMrnruT0kiqZo713Awpt6Vu
lRyVoY3/HIAVpjRmAp89lexuUOjVsxkLMQFDHFOiBBU7L/TzRHHmb/bgkK/4UPDj
uUM/gXOgoDADmGlpWoe04CyXUo8wxTixtbH56T6mA7d0qsbUquM5EhbcHuwBRIXp
a/ppGNXzKPpG+ppmayeihXNg6qoWZu5LezYwHfSC/0EGansHTdfPpBlYRB1DZFFK
EqK5u4PDWCZWFcONHu8kcHJ7ficUC80FygxrmpjQMNpnRqpaYBDLAjBbRRb+7vOs
FoeqSsJ25Ux3VjZT8G7RC9hABxMqjIE+wKdTgo7RVN3AJF64v8y9AqGDz587fN3M
9sI7ly3SGBREQAMX3wxdavUotBNNODYU6HZN1cDksHw9SD4qHz5hsxntx8+Xmz9d
vnm7EFfAdAU5WEBPNjWCOaumydQhRm9Sjy5qvylfIFHg1jnA14t+TnAWq2hj1kUG
OnvfMBt5yYoFgYlTinAX8GTQeLZ0fUcTHo5fsz9F7kWjc3MKcaGkh0WCBGTt2P7B
/RddRXcVQj+T/npHfLPPRL8q+YsHtV7WrxjKwRDrDTEoczijNE0+/a+GjYxDArt8
TRnA8jzA9+Rzmn4Okh2wlpp76u8Xw+z60HditKDxzqn8b7rD6qWimbaQ94knoET5
UoDy8vyohYuObtDkKujW4mD1D+i4o6VAIC1rtMiLVvyunA6o+wyru/vUFmfbZq3Q
D3XY9GLkwcrCezEasHUk4N8pAYf6y2oYh0iLYge1eLtopOh4jHsdG0Ldxo7KVuR0
ETBor0F57Ih9rhnKdo6NKBZkLObAXft81s74etEyuRiOqo3oku2kxR/UgZZhO4SY
qJ14pn0HdEiR+CdSS/IbdkG18ztnoqR1DHcBgtO+R8pxMYAVT1LUCzXbd/CqMQG9
g5muJXi97xrBq1EW8tj6DlMZbVK8fFLftucItAvFklenm6AYyfIbbSQybPQcYM4F
kc83AML0oz6UPtdWuuWfoyFSF+QyOWWYhMC7Hlpa9/wxiE3YRm8LoHY6c3NmlfK5
oof/CzsihJuZU6M5+LbeDCKChBAae6H8RCLn2xRkgz1d3+x/2K2VB57qBgCFrQ2e
3V0/09CGuij1oW9YYoO7Bmf774i8WbN80ikjOsxF2ngZ8N+rE9h5p3ZbcGGc8T3H
4JzexBq8vBNgFqjDoQVaqzpyww45lkbRQkhhxi0sqY3bvD8ly3kkc/jykIYJt9eS
vp5IGnAhWzIAF6+pBDCWq69LhgiICvW8zykswOVkVrlGOq6Bpi/DRgB1OxfYIVCB
FRWv5sxFKkwEDs5NFs01u7Rcee3803fJBtnuS/zvgyIOfixTdmK4FBN5Wz+E6XBN
rn5PEpfPqAQ1qAWux60dP2fYlDQeLchUjuAddqtzc9Dsto4C88uNMA5Ik6FQf0ju
JMNUMp8gwk/JFXsI+gESppYrPrwdxAwn2JdKnN7Q57m0wFHWqanvhCAR/RUrTA/M
g4C8bFgmf690iO6BbCxaBoWTKRlIqyj560WtxPRCopUj3vOApikI/Q+RYUCJHBei
77KQCf+P1vqvqSb+tv/PmM4LdDc8cM2QvcYhjd0HljRw1EDL7ZN7ckosY/wF+SA5
vlUGMK7I1jyhtBytZPk4nyo0k2CxOgkkzVdk+S4GCska2KPxY7eozwVnqIXSCdlk
F+0HT733F6it/tQsM40iycY4SGPDoxf9wa7BAbXp0Dgem+3NBEgYzi0LuedasrUY
V3akGyOxEPU+LNQrhx0/baURzbqKcyZ3SQajUdAcmdXwemBOoG3v7pIG7VQgwS1h
3zlKFRrJaAKfPAsHC2RtvnQJ1kYEV3LpZdF9QBAicMRYHLRc+KrZooCev2fUIxQ+
GtqAHlyBBu9uO5Aq4FRxeyJ9BkUKa3gpH/xY2x2Oyz7ajU7pEeLf4Kh0bH270Bo5
Su8SHgYG6oAEeoycuzfBIOCmkLps4Vuu08mMB+6iQ6okB9d+nON1aGXZj3oFsLlF
iXr0X2+c+iRbnbQqw9GGL7B/p2Jp9uPWBK0+ZywacpTTosswcChUjF/e0Jj509ay
8FiqXaJrVP7dr6wRHHPcX6Bqs7vEqDBy35O5Nxf6uW9brLP5AvxRqe/87EwuEd8u
Couvw3oeFN3RUsgOL2lxMytjdcdIQfHPPw/AZ837SofkNgkDU7+duKm+WtDj7nD+
Sv9/6dI1oMyTe0VgGWf2KTwb8cC9c3/9Fm5UcVIjbZo1OcY2lFBZyK5l6D5j5TqA
gD/HKN2EcrDi+aM57RkJRUAy6zVy+SgJt3E3d4d5JQ/LdGxC8mIbEkFmHO+6Csrm
p4lGYYfygvDDqZ27IDc499QsGbnCsuGDAJjX//X67gK2bSGoMf7j44IGSgPcns3o
qpjwKSIcQk7jHJ3tDwHQqVkVRtxpKX/LTc2kntriSPLXFO0OjaIifez8yuo8HeFu
wrgz/h1rYDw0dATQHq5VYufXKKz5oFlb7L4ZLwGa5tEODaAENvzqjywuNlXcHKt/
+8s193Is/Y0v6/accG1YWbiWod6tqQVelfbxekBV6XUu5B68+jt43q6exBbj3h+X
EzpfriA8Zp9FtUj1d4Yyg6UG9vubE11adzgJQfIA11A80ljaFvi5KMroLLOGiI1y
Bgry4+ocfccsLbrZJrkZB5jEeSRAWsbvv2wjA245TKWREaNdvbBEayYqyKV7leNW
1eop6rI1fJAfm0F7KDmLl9Hv8eOCU4LsdQvImAJfERAv/P42jFk42QS9xkLSrtdw
0XsHtyLPf9l8iDgpayPixAvP0+COQE8+Lda1pQ+AcfsjTCYn7EALdPUFv5CphN7e
EosXteS7AlvFe2DdSaw6JwZ86eu0IpeBtX8R5yzIHVDz2CyVNkRswmAck7lm9X4p
h4wW1sj37KbqNXMdoO/Pl1jfxFEJ8O2sJdFOR1/Qy79xas+qKnP2sLgrimEKDSBI
mmCRozjjgR5Kq0Sd/Aai7sB+SZ5SC6u0CFkegmbDEecdHsET39YYQmzDNe52h3R8
d1DUtG+kMzXK7nMvacehhLlm0v98WxrdY79BAcLnPisLx22vvHx21Ses7mkGk7bC
VCJZb0k83gYv9BFGS8tluRD3nDtbXphhcFsbT/eohbZJxikVgN9vL4nrR/XYlb6a
WcNQifx1ZXgkl/zq+1wACjLitwb9oGIBKpeOWF1IE4K3Vke572lTSlsf9iT3utGa
HQrIIM6Sin4R4R24af6O/GEjlJv0fJTIcZCMtaDGUyRjOjs+4z44Q7R7xkWbdiUJ
r3derVvu70F7wKTs2zi7ySJuoycwzGdBzXfBIUfWXjw22sDNvE6/xFbqdG0pSgMT
tlB0S73/n+u3Id9JT39u7SZyje9p18ThmcFMohDLOtMFfGeenipN9HZlssy6+evs
LxJkEaOLTuFg6kKNIYxliG/V7Uvw+4HFdZwTZdwwjI3/M3ci5IkFPuNvBB+Mal6h
RZv0uRmsKwKJtd9PXjFinMTzw0z0VLI1QEuZcNGwokMd3hy8/hIDQyDuVF1QNdej
3pCtYcrYx2d8bHUV4vYVJxH4VFKQg5dLX2AF14l7nV15mUUw7XcoJON77sikChcn
uf7fm4QDYVNsu0YKaZU+1KkxtHVsQsavf39u0uJ4zPFBfEgnYHxOjHqbc3W3FNRI
rAJo5fhhfwUYNzjkqI3gEkUmRXQ6r3d0IPPdJmClaE7GWthRTgYKcJiIyNre5w6g
XuvOBKXLmfGZzpAKBnnMT44eXdUBARZ57DWmzbZvWfmHGNfH59tMl4M5BbbSYXQt
eojX6aJR2rEXdfnEZOOYboTcXkCrOC7eYQYVOOJlM7LAmCqd28aXmkkQoSef2Dhg
/3h5Eu5Wj1/o29dEcoyh0YeHl/pmlibUj3cUF07vTo+i0e5UWAUiTndjTtTReTou
jJAgjT7Vs/XPoCqfZCmEE3Xj40P0aGKKs8pbbPtfTefiWrpBYRDnB0r6gWdlI9jw
feMC8MeCBKZ2n2f1DGfAlZ1Uksyw7l+iPfbIT1V8kHcIyFhvyRR28se7uT0h3QB5
GBbBkfjuZE1lhLLhLHbfOXmYkPEKiXoYNTd5yRCyFoPlnHC1Cn+jAGwslyQIRQvq
lFcKQazAXxEsFCd3jEt2XQqULWADu5O7+49z8O1oM4p1nJYXLEjr9YpOJyEJ9rjI
bxo378wjiLxdtbrF9re1lQ4nz/1S67rC9Byv+eQY61vNO/cSja0jes7BH4aaUCfV
08pgW9QnkcKQBD27YYqCADjtVqcgiHL0T0xYtFMUqs58zyA/kK2COVcrzhndPM2x
w2U5J6G90A/PJjPqN0w/TRcXDjkkj0FmYNAWMcqFOZUKToctagh9e0QUa9+Ik0il
I7iCTX+cIcKfNepW3fiIh87J8Um5gwBbPwFfj1qvugtpsI8dd/3c5H8sBawfrPYr
N7T0iEi0Yyg8VWWlPhG9DBSE+GLqs7X43Ihi/PUjSgIkKLyoJd30Y7I+pS1paMsS
736KJGmJCdeB1MxGSSoS7HJL5YLoLD7rTR/2NFlRlZIhYt6aOPpq9yZ8A5dM4QUD
fWQSaqG1MPXPt5IFYkK+oTtKjej4XoulwCX/Cs2bloHWwNt2yMrfRKn+G7CPrLhr
H0B2m35x+6zktR64viFRl2dUijtKuGMd+nJRb1Fi9vbxwGvSN45dt0cRAMDVtlUW
R9pTec3C4fa+YdMFCZtvybr1PdXNwWmlJFUK/PrWxsvoTscaOm5prpfUN3J8rBT4
wXXDxAZ09eeTLGZC3mACEvysILmLMrvfc94U50pqKPSQNcSXRJymCj7IMFalt6A7
ijDVA+HzYRvey1lY2hIxKFbTJicxZZPi3rX+a6ppzbdsup+GighBakpwwdbLgpiD
CiP+LTVSh6aeyYBhOtJyxKKcYhTfKCZ7bRnb8RF0eMXJXgkxGt1P48jvVwyvIILI
R2VXBMnVMgDD5QdWaOPF2TIpplbieTDcLwzyTHQFb6fzzjoB2Q6KAm5JNdM04doO
EKHI80K+YtRjkplYJDOX5q5T8Mm8zgvi3FI/4PQHZpPxLXOJzUyFohNg27JHKiYV
AeBKWvY208bm6jDI0niAEwtA8eF5tzTT08BYmD5SqvTR0qo5V4SkitPrfKajN2Nn
0YwDIXoO0MYsMIl+j12i9o7ON4xtKXROGrIMZrKQJdEKmLEuXDX0mNDy3CpilIo7
7xsyEg2/uczD123l02aIK4njEJ3VaCY93RU1fSQ6dlPr6+iJY2NcT+3LvILd51hP
2MgyR/FEt4ca6avM2Dmeg8JHnfvWgGe3rjCPfwbAm/DI1JtM8FRjj19vIStikfXh
R743NhSk7TyC4oM7zD8UoAPOqfVSwhf6oLGNlEEEzZDrdffyaD50vi+ZYY7X31qX
1EbeBT2wrLjeGXp549J5JwzE9j4ADVitzKBlQL0eZVmB7S98lvytHLhV53QjEAn4
pRJyBk3ZJMJmlKKg2W+VWU7BiEQSPC0JnJT2VR+fGRuPM5ZdSk5Ty61IcxO0gNtJ
EQI2e9Ygp9+XiWQrj5blWdx1FfQUdu+wmYdPz22j96iMrWnkAG7eN2fflAqrdL9A
kN2GjNOSuhCP94SLvs+i7OPELeSbYdiO/15zX4OLyUlr/DChIqB1kdbLbcuvBb7w
O4WByd62JMn6s8q/Cse98lv8jytpdpon1a2szgQLeIDTcRDfPqtlz6b5A07g6/xc
9vkawYuFC8ecTn5AZX5SpEjeaZG4EB/CJFUIBTUtsD4B09ou4WodXGbvlee6xU+E
qmmjTwHb1vo3udOS+OOE3PDqWD+L4ZzrYl2LWD74Jrh7lK29QAUSeWZ9ef8NG8Jb
uZYKhjjb8J7E3Y77hybXPLiU/jmBX76+EvT8dECjQmlZBfO15GWZhHp3YyQhrtEk
lmfjzdmf76YrlUCSwLBCBlpMH5vGR8DIr70QOSe3xpz4a+JIobai9lg1dYhVfNoy
RpZMkAjAitswFcEWmzfARvqpJIsalvgS1bukJIrOPeHACCoV8ZnJMUNJ6j/4oFji
ig+pJ62IXY72pmBExI/ni4fnQL0N01iyrg9yRqfsLhBFI3JX/nT7Jm31LcD/jPy8
BQaOKkqhd0r32E5uEpUmUkU02+hrieJgVWd0ZHmsQVf8gIdt+jyM/q39jLCq46j1
2crlvH6H6oJ0EuyRMIvdU8/UFbOxGK/ig0vBZmD5Ubh3klcIact5l456rqUw4VDu
2x5Oq/U731Y+zhkX70VOO7gsAgFLOdEge559HcuXKuxi+E75KpFdnOEe1vAMTUuy
9+p3hDq74ZhY1ytUyFYQgiSfK+ypX6HcFmTLNIbvHBw8xmMV/KhBcUgrzcP4Jsx7
TLal9pjkpoPaklMtPv+DBGcxadTyZg4eGxgW5Tt+jQkHk/DHsAOqfMQ8N5lZMOo7
kV2G15rDDdvkKRiZ9LB0s9y9ih0ePGZNEkh9o2nmPpAp5CTPrs2tUMfe/t2+lGsL
cxIHgVIzioZEvn+VS8/XpRgq5/XsqXxrnHSs6Jlo0CL+8YgHS0TbSgrs1Xu7ZJVP
5TWCx5VxQLD9acNS/po0TJ9sMwwd59JWQwIOmoKQeHOvTvbFYcKFZqF4/YQjcrix
KuPxwTu387KFBRPmETCQZmKAW3XNQbEk62Fp24ftpNyTRqKxw4xcNyZEd/bVKmay
iufMM55ggvQVIh5VZPXVv4wIO7w2+tcidEv8QRYoEZJ93+wIO6zewFhyc5nkiMTK
pJ9tty3jl1xrDnUa6+hUrhuJGSRT76KbnlwgkQnyOrYYuISzjR2EYVUe6TYPgEaj
K0nbDZoJl4LqRWdEWINbpPRRhtZOuL7oBGPt80n23OmX1faJ489d48cMZTDdxICq
R7Ff3w0jnETJrIz5aw3LScrtLd3E8hKaHHyc7jwTH6L9GOi5s3J6g+jFksduDRqz
ckv90+qpjiFqOBq0HpK0SQXWHuTwXeB3Cx/w/t3vvOPVOl7eQVuG82g1+z04ATq1
WsMq4blJcsxCaHXq8oVkQBCc+j8YJ6tWNxobuMjUJ9nBmHQXq0CUch73yNp7VPnl
03RkPmSktht7UNj6RXOhDIbHQ4EsoxFJiiHl13CPZyOQustSekMdiuMtL52FfLIB
PSOOLQL3KIFPDqkeb07upYgzuSfvCyblE/iK8FGFLaWDR9szYGVXudzavUvjmVqT
HQyYDwX0j0gRzEhIBOIxEJ+OTW5Cr+j1bz0lQf6JBanz1YHatQ9TtZTbbcxnWk5/
SsxEz9Ld0/b4CKZ8Aa/qt1kTez7aHYI6bljXqouwaWEGT+JgTf3fv7rQzr9wZDZa
1eIZmtXtY4TnBCyAMt4uzd/7POFxdsT56MKiZt1l18sbwkZvT5jlxjfpDRz9pdJ2
ReBUS9Xf+TIOAT3Zet6QSuoC9yGt1S11+N0sj+DM+PLrmZlJDffG5WXtV3yAt81g
pGW5leuhPjBfrvZRn9DhW17CREkZAvun1OcpbOsApy9K5O6gpZeYbvnlNEII2Ydm
0F5qM2A2TS1Tf/14THCk/7/B6LCT1E7mG85oTyrAoke9BU7tMx1mmAGJEOjgzP/V
oPGYs043UzX28Nd+nBfTUUCk1jRTGoSNqzw+VeXO2XYVd1TKlRsmh45Q49afPd/7
/G99emjfUoUPty784xUFgvBxHeEgZnLAye5RvQJn1DTv0XXxtPVMP78FYNiLMHU/
8JDfkyKztZn3EpbLo0vnmXBplwk9HOUFrwsHzGY/bwfH85oy7ijA9evcKCNKCJpE
9B+BRzcKTsipyO6jUsXbNlGrT/yXspix3InjriTDFAjN0PWNkiyWT1R5eIj6T9z7
ZOQUT+QRsspnjtSEkMKd+sATdJfjbylD9tAh4rATTJDFIT9FRWvdd3FU3LDP3RBy
axC6wo5jn4q+aXLXARO2fUNJpM0Qf1+pns8Ccne4T+dYh+AT10MHlQBRpSBUSiKS
nhRj3MmDhvOvDtBIeasAWUi3SmLoZcXP78yT2iDhryzJvc+a9uLKHorKJeHouhJ+
9MM7AQhJa/4x+N9XcAUkF2awZbbgH8sGDjUzQhP47jP/wSac38UiZi1F20+QBbmE
JuAOcbhacFpRkXJLQyJhjSDc+5CQkee4H4Sx/5UofxmxthLciABtdnl8Tk0uGUZE
Xt0TZY6gl7qV/x7FpL0i+hQCwGjjiyU+VJZrPZ6n5ycOs2FKG9UNlT7VbwvozXGA
O8VffljSpeK11OIBpT4ZPKIdkdynPEDHhUhHxpCN/EnC5LGn0dOEennx6c3UsflN
bY8dO0ZiSTo3HQdCZRF5EViODkz3Mn505a5q8mMo8CMP0su3pyd2uuWkr0wBKaLo
B14tEiTVSJQ/LNnhrHoy5/+F4VWz8zEzlAWlKfmk/pNSRStcXBEjBjAghkYSu+Ar
mHqF+Sh7gqLTL5UcvlTRwWiEJDAzkin8ue7Fc3JQ7KZ0/BRTekuiCYy3lM3RwmyM
GeDFMn7AMrd9Rgm0XVSgseezwmFN5SF5EyJAWAykthvFivrOShbKW87kWxZdsgiC
1NVPT4kyCtRmQ//F6aGAs7ml321rmIpIeRic7r5iybs2S7+dHlN+9qxSQQ1joW9+
4d9jfsEO3HW1vp50+aYpG+tna+NvkIR8yFmP8mgtSHrYlTySu3D1l7H00YRPfvIi
fUKYT49YroMVfEB/jih+r/llc6RQFGdsaDKgMuO7ciN4jut9o5VrjQHpNP5/UQLF
LoIZ9FMq2xPrknp0g0QpauK3A7xnM5TK4c6XVog3BzsDfr+PoBrZIxnNQQoa23fI
qr9LfDuiLCeIUH6xkhalK4VLGGOGd//kzh1q/jLP8/X+FAuScQQyLmgpOaCn4epW
x8mVGnIXFCht3N1A/aiNzPoXgP/HI4icCrufaIixwsNCrxqnZghxSLiAmIgZbNYc
NHQPsvCpcSzgMcUyHHx6EYoF6FqvttAs3n9suetH/iMzVdED0AufsvrL8EztiCX3
/fkc5cK5nfUR6+x83QZsSphACPDQp5yi/W/R1gNO4ZeDGu5Ir1RxmKj3g1EVwgVW
LmcrqHXMED4VnkbR+mMYb5l6RZfs9pRUN028aOPiCO3vRJb8dIS0x2uFeFrCf7IG
L/ChgLVr2MkxqDdTdloNDkyPLYbnk065x5+dJ+WFoTRxHQ5Z2RoW2BKrZ2SlnC+F
3tjwred/bLM9I5vYbM1EMpOIqkSsr+ZlO9yklDHple7MzSz0mgFKPXOmzenuSj0x
5jwlWayujA1dBZERxIRWoFptX4xytF2CBWNlOBy2Z0LnnRWQVXhtdsq9jO9zrkbf
zBCKY0w2YRZgOiEteX6ZFs5ILxygSn2KkXS3n7IPkEYZNddCpzZIB2Z3PAXPk504
PtQDc/xGGPOrsrFNBnCAqX8wH+Amv50e1Aiu39RZuordhVk5rxuEqkxqFzf/mCYF
GOro0IA01MpXYxAz9yc/I8lnuen5jSqE2Gv20VHQva8lTy24M1oSXemrj3S6N2lC
Frwb3ORgherXFtAeGd1HeVJYDxilPJUNf+r9Qev9UT0+KMTlq2l7hy7FLYMbnEGm
BQp5EA8gdSuvgeG05QOJlaNnTMxzV9e1YLb2MXmJi+mQBzPZvoM+jjUGcAQl+/nL
a3kizRPHhlwPLCbw8hLeSxlMnCsFP5rFLnHQbyO/ZdqIs6Q3Bac35N5/g3aR15ba
KEaBi8nIgvK/wIh4QFCCcKD7JyuSaCIRHcA2X13wS4LWhak+LxOa/HVzziOXKpOi
4IkWifP8qMlKkuIG0wd4s66K9d74RCmglDczdujwFvraMOFYVDvzpCaHvgpLpmFq
ta2uFBH+eVVg9c5x8JNi3ihPSFqhCkwGec1BOYKq/liWzSA5ChtHRPoSnKFTM1/Y
Je3d5N/zaXfyJSqPzFk9fLwJtyOYQf3ZdDtXIfgozAEahFqBQXITUikydDgKLM1t
0j4azrbmAJnP3nbPytCWkby4oq5/faWjOiRb68fbwNfn6+IJIg7gEWfroZtVp+ki
k8OX2TVVYU521t1XFVqV5xxx1+38D8Gra85eHSzbXu4Zy4eJTY+7pbot4JIxXZfR
HPOdGnYbjxAW8VoMbnN1IvCECSapy6v0aILDlBIclnSAjvt+xcgGl7CIWtrM5BIL
ViDnATyJ6EBymqjSUHnvSTebkFQV1yfJhKFPOi6dbco984gTWB7JfTtNETT+dhmR
ENz2RLmSqEgd5CgtVHNVQmHH3ryL9vYZJSFxqQUtY7EYU8+Tj2ajpuX9ByreAIEC
F/qAW9QSAKxSui0S4/iU72P/wieOuGEBeOfp6qm58+POVd5X307Hf1cx+RVZacjl
z4iLiULDqBK4thNRcDjo+ofLieYj2O/bdH2wr0BGfRrcbVg1HR706DgICM4mlD2H
4VoNi1QGlY0XOBvxSsxRGByaVQ9/8wMmeogelKQ45GKw6TUN9sQNvdd/ZcJqkvNr
eeZwwDpvkFhTh7JgmqhGPvASUEpRFONTEghOU1v0W5p0kxhQNA813KYmgrnZsPb/
9S6WDLIW+HuhnyeCWwjIYaBz/aRetIsRf/o/Xcu/aixdmecqKjCPrUeR5snQYYUM
0mdQ+lWXDMzzss5YYcK/ybRvZw5TM/QKc3toaSyUOX70H2kcMFWqbwDdKsIrcr0l
z5kqnjyNPa9rxOASpxBRJ9m66ZHTGqRSCZ6Lj7r9SJJRydxiOXLVTav/NCsK4fH0
QHnhU3FyCbvLBWaXba0DRJo744QOrAdRONSMBwGk5eA=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14192 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1adJXUyNzEKX18xw111ld7mXgoypzN796waDHH0d4t1T5
I0lGFFIMz5EjngSWtbSUSqbOim2MT+8xeQRUqtSqVBkORvEee546C4FX06Q3xoQq
zrRC+FDRsJGzBquCS0nDs762a21RX8JibExeo6hmoah9+gB0ElvhUXzn7Nb4IzNB
+jqBfwMOMPmzddQRg0+B9lcYFIK1WmxgV4/v1AO1zWPPtlhVAa+8UV6CsaZe6bAX
0pl3sLZODCHyOH85GfWINakofraDTw8tjUjJ1GKjcu8oNJq3SaXdD36cMhd4Y7jI
HO5MhbuhZdVU9iSqjVmeTeROBhEvXPlm4kBmAFkNStx6uGPVRXZISl+81r08V5uL
nk55MpqhwJUvAgrjVh3bYuJ+LqJ9mORI+g7NHtz7h9XsjmvcpnULnqeuprlr7Crz
ReVZweKMlOVA/AFk4h6vLf7tJEo9QqcIyVsQlKTNsNz2uTkKp6C64eObHgpctQH6
SyHol2zmvyKKtSLtIRZpo3J1d78ZpvYswY8kse3EwXZhJEQ73HdqHfDXqSnK6Xko
orrnwSdx73gnlf0lKI4Zg8DxLKTtoYtcVo+8kXlCFnWFoWw8l8fnNWe0/WIdvh/T
43qLNYGMYUYp5vsncjE9B9KBc0yWGE5QSRmJUq8pzoam/pNj2zP0iZTbnt0VXhTm
uxPg2vIz49glVQjNVTwl9nYt3ByTbfrGEmXlzHdxyW7UPdggCL2cr+ZGfikVDe09
BL0G2al3ZRlK0xqECDup6u6/w/neDg+MhwpfSKheh/jonBmxRoSS8uVXG1vYa/as
AoKLwYl74KOPE4/WRTZFSa5PmKvyfwDB+gBHf7XnP1Rm9j+nF/XpPWxr0MQygg/g
udFBgvS/Tk8rjULKgj6QW81eQyi1v9N6EkiVUcK2yS7Fm5W208ypQmL9O/122hHN
54TxEJ6hkoBF96mXggoDTVVhvYpaZPWGpRKAyoqPiesRVSP5rA0wlpo2yGCjiyni
rFo/FTeuwtXLUCkYCF6sjbxglcYQxw89WH8w9blZmup/lWDdNJosVoNiV3F10SeC
c3EzXmD93Nj4yP0h6PtmfP6Tb0bvyzptp0Z+Tan2NmY+FCuQrUJTo+Djch2UiSR6
DABtsf8DFh62224NjRJD9RSIo6dzyNccaKXV9NAiX0bhc6TrcJznMZZa1LkoH7lz
n4EvlT8lJX12yEoodpz7D7Aq1vNpNs4ujSfjYDy24KlUVfhD4qplSO72x0GiuKH0
x0ySgNRhn4QOlw32gyHXu9a4V1SM7w2B+bAnUrwwbhS8BXqKgeGzhmBDpjvUVWc2
y8c0DOeKyQeFqa9B0Du7diQaRHsH6hRHv0DcERncxrKaLieraBh8IX2c9gelE+6L
P3tYZDT+GbAwzfAI0tJekgrvTVBwqJDbaFXKPY8nAt995HFPzZUnlb/co42cWs/6
ZnLREQuRVH6Ew2ZRZjKLyGZ9X3YPiRzJpupAoArvCzcxDEGzDr/k1ZUZ07SbtB0P
UsPhvu10p2neE9igMPG4rHQYtddAelJ+dJ1+s6v9B/Sza/gZM1zvwgMKVzbAj3gB
AKsfHknweJZ3wdwKa1tLUEpBRlCA6ChXxDM7IHHui88SwEFGH3ahZ+sTIsb5h2AL
epGTqHJQLZlyBl2ZW2+7nZREvTxht6R8dRBmkwgYRK3jzzUGsdeqqnzRt3h/fmv7
KP9dXbqBCc82fB4vYCnc7CCGr8BYbEHY4DFUgzLDD55p4I/ytwxTvUypvQ/LIXCT
qEt5PSd07CbYz2P0T/1GGbhkXFbU7Wg7qaaD3MR4E+Hqf/V65ncqaPXstQzlzDtv
44R+ymG+vIdy4BAEjlsP+UOWdSHG3n89e+TS3GtTY7nIJCwA2QQLm3ATmtdU4aAR
NnT1C1jKDIWp98rqxizBNnDqZFbKPMHaFPScxjf1efS3c7zv8IKKsgrUxQdywO5+
x4hfTOxRcqFinzKYngkCdm86UGCme8bEnBIk8wNKAOp9GnxCo/eNHq6h/WsTJARZ
bEJquzuAQrK+84PvmpC4Mzu3lS58eCoihJZ7gri+Llp8hBvQTBLYv//CCLsC73WP
q/cZ/9CHFVD6xvqk8nqBJj57pCSCOsarwIRvWxxhqGJpEzFVJMmnjuTwsxwzSn/v
5iFqnC+QhsKEiQLPu4QCw1cDU4Sdk4tumj8mTCWWkyJJSsGcKuXztFjZMCDl0hwL
1RgTksrTN1iC6j75Gh5dvIuuyBUEFiT2c2tTTyRgPra0L5I1F0QKIpCXjrevOzsa
ejQl/dv0sYWifGLLhZSoSF6D7McYzl9dzrSt0jYcVQR2PSmaxznoQhek/vV3x2Ff
hcMMTY7x2wCraKW+LjvZ8hUYgQlCLfRcviH48CmEGoJVgwm08HmLCE5ha9zoSb81
ayWeKXHlIOudwohJm2BKuPC+vSn0xaQ3WxWesa9OdG/kOz5cnOXFIgvmPptWFSG0
DNAEfcLbyu2B8wj6rdwyZthoBSrn56+2rkTtEznsVcx4CYllMDUU8UJx7hxoEu+o
H9521R9e9/FBSw4xUtv7v0v3gBA/aKEf7igcSWDroA8tes8oq+SovLO47wlFJcfc
uvSfSce27mppaMR5y4CY64POJquii3bIBnOc2ghmvTlZD5PeGfiVixjgsNXpyQGL
6WTh5ijp2g8MTXcSXW0emC88rzKYc3hrqfEwfKIiA4xIZDXBLdQmDxTzYc17aKXI
9QX3TkaVcmssOfv/HslItF0GUy5Nc1tkimAM9yCX//82W3TOXOLSqt4dGA2214WN
zI2/8qo1g3aU7olZO3rgH/o0SL+NzI0bOc9tqTnVTPEyubhy23WO09SRyw3c5hpe
+TaU82FubvcSi2yDyKS4SFvXbxWDHCUH7WJK9HWeMrrzqJklJwCpVudMvaZeGg4Z
q8b0zMsqJ6Q9OsKYoHE6RdypoL6hL/QbLjWnxHfXrYN3SVz9ou9WLfQ+uP5cUsgP
+1yDRB3n7fo77tSyZp4uSVOSI3Ei9XgskWK9F+NDCUfFka663UZWxzmSCv63yP6J
DRoCD22JhO6jOUaj+1g0XA0W+A8tutEQv0UPcmCIyWnH479MjvU1PAQc5NBpCq5i
/lQD50cBFu/EJ325H0mcfC5ptpx8eA/SA+ZeRIdCkTAeifVbQtk22WxmoRbBxCQG
0jzCyhQeBZj4TvikjqYtrtcUm9lpLftg2hKGuG/MtCaRXaxRSxauubY0RpXugQaC
mUItWKFpMUo2LnErpp+VwGzFaFltRlZK0S4KP35qx0yX7wetzWIkTN9zjQSUBLZQ
SvPCHKIlUJwav/U6ELqKdMVBF7MY9DVJEtquLHwFVqTwBZigD11pS3ej88J2c9wo
YMJfzNicLnVd1eypVmcma64SzOGO2fzLKt/m7E34NGQN4afcYpTGD7Uqm1Q5ycq3
Uv1b9kXSkKLWUlW3oJUj8FowUe+EIVcUqT7l/vcnCInlvPKYgXJSI3CyKjbHF9c5
aZadG+ZxHomLFsx6Xpyf7feN1wE+0tjjJCD3hLCFetg8QTl5MpUKuHbfhiJxVHVM
8BY4u2OoRTkRgvt8VxypAZJV5yDWp6W1FI6H2D6k2jthIPQ3AQ21b3RMf0l/ZZHU
OR50TVwn1cfwQJ2fwtVcl1djcRRwCGnBRXE/1ev3hg0bTta5KC8MQ0Wh53N7MVNh
taA3hLAB3H4eZAFXANMjdQMM4p5IWCrbSJyOrX/Djn2JAcSecYHVql3vgnXEeuUc
ZJZGH8glZZ0aPKJ1PzLzN7nzdBFrXmAKi08WL8gA3/co8u8Oq4N913d5OAyNvc6J
hCPJLRZjSHexmPAS/E2tYbwtB1cFSiqbHbladR9xmEtYvl7BMmu8xPoyfK4uwRSK
vtzkC9eKvTCWN7uhtO1ru5tjEnlYVQqEepXlQu6Mya6WtWLsZvP/Afzf58wCjrm+
rtWa7MM/kcHHJK1QkAgklN1OzKn21MFo3ZpyWnHRQuf+IibEOtzZ97+b5OWT1eOv
ZZr7SjyJrPnfeyVc5n8i3I/ZQk+qjuBCpoVRwHuRHdxeA+yl+geopn1KW08RdHbR
lE6ZWI/tZTZpgkt92wkb6jbuB9W3+lTDoit5BUgJpoCVwGhRGpPdmNZzYpijAVOr
7CZPvZzrCAMom05l7WekMw5krEn8QIe4/EqBqCTdnitvV8f2VIGL6pNk+PeJiukk
mtl81jiiUhQiXWvdJ2cqwZhtW0RAujrOrp9QTZiWornC08I9YZYaC0YL91exkbW1
cJ2IwqFbVvZ3U1qAhJM7EXxo8yay0spBxI2ihvgqVLzEkIs0Rj424pPivMJNSV6W
VyFhfBp8j75mh9TDMq4D1pd1o3zE+eCTfE5QE2ydCzTedPydBdOpdGC7Sw36UbT2
slyWYZNsAbLkmeUHXNoLnvxUxGlJsAgz7OPB3C6f3MtpM5LS18I7RDYyqc7eUVeI
UM5BeLIVWr5O65Ye9Le5/bu268aPUW6obeh1WFNo5aT7TBlLX5E4HWPOsNwNL/wI
AovNr1dLPWR50NrFHUx1saladHgxzLipnb0Ft1/UA8xBNDCcexArhr7M0egrEXzQ
614kxNi3TCdETOLHSZH5EgLF9iiKmQ7RbEe7Dqcz1mIuALT0GCnQ7FB6M8JxO0Yu
vJgmUj7uL+Zxfe4OxIZeB92K/LIQsbolRKBKcL915WL7ymSAOuHdFrE+1lHNHyMa
uzcwYez26lxqDPfqQsbn2bPdzdy+l1HWNSuCtzXrQRiF3WNEAM9Y2jlnIXrSGVOF
qGQEJtm4l+jyhbFQ/VIkS5hjmrf4DoOKQlxT7rF2KBzd3pMbh9Ez7mV+HL1s1Byh
vkNoq332wzko3hQGqxBo8i0FNdfOHTt1AHhIxKDWwiGys1iP5NEKCw+cdUTCMW3R
mjRR13yYmTDeIV7jVkBQWqfE5hWWTVYOd6ZxYJekQk/S0aeXvh11UTzFWvsoTnRT
gP9SfCPbLJbFG+hTjWbarYosPJZrwqFqEBn0o+Xt9F/T9gbapwqQkDKXkCdTc9GB
ZynznBSIwXPiQyo8h+hlw6X58vT9CSLcJNbLqRVCxh2T70Ydzhyvpv/xjciByzjX
6jnm2/Yb9oRRXz/5r4eUoHVLmb1ryo3rG6SugHV2RIe6gmpfjGTaZvd6RIjY9iuP
IYel0jWpbue2N18hijXDokq5WFgAXfzua9nlcmk1rH45WHz19dsFY9rqyIgdbPXY
cLj9kYCRXFoEqDiVIpt0dUpdxcMAWl/aqIQyyIOReTvQt9+iO76EiPQd9LmACIk6
xLfLcq51jvvBcslEcDyrzIon/RtgbWrhKbwZNlNUHI+uyZeFNDSm32sR+/r6p1x9
lsEC/qehS5rfRjp+26EAC3iXUJZswg9+kC2/myj6TiRdJocO7+beF5tzU94bldhx
8WHpKNgJ5oIJJbMmevbuEIjhU8y4eScq7SaQ+g/wARN+mswUBzLWlWqvPKQv5ANP
qfE3h7x6i/myAtCDeIKMql+F6oXHW8c/4ffhe6t5qX/XuLu4Ni4HDWf1V41xjRAA
4/bvkVYn5NRBME1s0tfmXGSy1uGqZwmIeVzfaXKQWKvWLyXxQd+VOHACqPbWYeKo
L0G9oNxk4gyZ1w/q9BRupWVGV1XN00I39csMU1vEQNZiZyQykCO5YB+hItFTTrEI
jtzjCC4D9T00a4KSkI1yl9B44ELy6SMutLr2MuYdaKtlAD7zOoc1R0/Rhu0JJFXK
G9qXCt6kXAManxIDNnYqNUycH6WWHd0zCWtDTztcJDL1Ty5RR6lcDItAKNsXq+Cm
XOyN0ZslH8QFAHZT6lI7pWt3f6vRTBrUB2xUFqJ2cnDMYDSo6Vn7HarNgAQIroKE
2zMPsuEPh/3UKYX4e8iyLCSXdfJG+Uqg7/02DT7ZwvUFgdAeLcnoY2baqaW9q+et
pOVMao48hqaDk1CHa3DUgpD+GUKhjkVJAPluuMT/C1NU7cvOnPHgMP8ISFdQMz8i
89a05FVbsr8vCcq57+WTTJINzrLINRu/pV6mb7IOeFj9OReUz49/tTeVfWmrQWSQ
AoBHMpbvlimH/fJA0xRF9kx9IDr7ao02LF3ar6jxFwQkNXOEKuosWwlS2wlrwjQY
7y6CBoy/k4EmC2RBKdFm5aH8xtAZPnF7NDgZy4SXhS7KM8o9Mx8UKB/0ozyxjRRS
YAnvTgk/ZMCEKg+oL3DGvjOOR8324+vOMVzwrNT32aCoYf17xpKE5lZKb7pzl1e2
6aUh1pwe2J9iXiCyV28e+RCrst6DI01bMuljqJlkdX3JDh/sDXP3eBER0/evy19n
JRNQ3djmQWBDasP8U+vCYxM3IU2USbRLA0jG1ZYmdPbpnqCc6JMEhQUw+kwddO4t
coL5KjWZ8ZWELYJJCQpMHCQt3/zxqXH9Z3MiJBXZ0dH/MLMAjgol9OVIWx6wwOyG
DqZj8JmN89FtrSi2xYfnW4gB+26RXriaIbQam31azbQ4lduX3D5FyKOVsE07a6WO
gkWw2meQIjUYFNgbfi2Mq/y4/Rkeu/mOxlNNoXcrjGc6lIS1XGrjQE858V08yOfK
2WM/hRt3DABAQsv6DyJoxgoQ6VtyboaDzJTD//7r/NcgYf/09YMy2vRjcLJ70J15
wLXF25J+Y1Eqswqmfy8FoIkYVfl9nVo5qRAAYlM47wg7E3QZ2R9nTP25HyEmec76
d6gTznidvSGYlnpsGAeQQmSq9TH98uqkqbStO4Xjq/8Lq0hinwtW2/Obe0TGE8nA
9w4smPDy90AiPfADC+k6fupoM/cSOtP4JcYJwbgt+SN4CLLeHLVYAmkuxMrD7is4
WZkKNkkemXY7zTco2GYJriY+kXp2lU50l8HfUvSv+ZaxActrbUQszfh3qAhOETBD
PkpVVFAYQQ1TCfujUvuu+tm72XWWs4XG8XKtwOx8MQnsNQ99VNcY3f/1UYky99ab
tB42+R9LX7dgd/tFnQUJa9HRfsElspcI6+fGEU4Uk9mylfQdkTrXGQbmXYN4Rnbw
+vxvjoW3t8FDf/LBqwtE4Q2zq3Yqhw7Z9blIXp56Zxb8SdqLpArUGb8mf8Z2/DT9
27TQio12gwfmCIxYv9IkZlw9Sfc+1+gsBZUwEcis1uvujWNkLjKCs1fZXVM70C+A
/DUfRvBBOz5FvDXu50R9RYDnwDRI8QFWpJHP+lgd5e0ClV6EN0JqhA/WaItQJk2p
eLGcyOoY224bUEIxEi7JWhi0Jw12NgJG7UfiQlJgnP1pTiirIIkM5C2OzfiWwWt/
CAdfsNQokh4z0rQrfoEfPkJmKm2M/WySvvlKD/XAb3S5FSnm5AR7+Mnx0767s352
d1J8l2iqsERR//eBetVO5DOqZruPHsldZvZFdX2/LJgb30/gAEN+5O6u9A0hM1Ni
qVzwoqtquiLygQmWO7LlQXc2hdOFGbrevFl7gbPHnsbUhKryGcVc2q3Jl8w9d8d0
sNK4pJYWH+j4ckX1Ior7SlblT1aegAFljLOSdfXolqSn6OSn/uC1v15rPtApJzS7
Lz4Xl1msc9QHCi4uhnlY14sLQcVa5LMogubJJBzg5cMduzeSfFETTZcTC69K0Lly
ayudLPfbxy/CN4SVmfVmchD7cMW+KymbUANvfRY3h2Y63TcFrs9bqQ8Gg49SRxWX
a9xEG69p/UKFyboqgLZIms1ZQQ7qRyJfh9++2hzbNRuhm1vVPiVWFppGQwtGIQlI
jhqNE1BdYYgrL8OyJ3z0o2B6Zhe3xHTNqrXSwZ1I8D4Qma1GKAQ2eAiR2ByPsaGy
JNd8ExT7VoosGQfV8r9J1e0RrShlnJ5R2TNp0LLsRZU0C7V3uzsIIMx5irrB2vX5
d1+lUyTMhKx0yufE2PjEvQw/3Qrse1RyU0TSRMV0yJaBsGgaUGLElxbBWOwgfjXP
uYsyzhTLnCJO/ivuojrWivXfTLL/N3ONR66AkoRI9QoTNE3pUVP0RcIDvyfOeLrU
dZrbGDUjU6qXjzKdvIdPyKTF9/KRnFNh+dG1qBOhuMrL1pMOws6CHS7X3BH4H5KR
ObZejtSFgsD4lKkGJr2FmsNCVs8omlcjURet3vCPBqyhlljQrbOKBRlN/LxDsrM+
cHKZ7Qawh+Ah1tls9WsbUVRaU0ceUjeH/24t1RiWneN/MwUJ0rkGFZiM+tf9CSyQ
8rQsVLqZeMaG0Xpmfl2PHKr9X5WTI6bnjJMaNWb6ENknvNE2yYLfMtJR5oEDs0D4
TJZ9IZGCCuf2Hq0zeUh4RPC2iZjUkRQVBNLcBXGF2BW+Qc012W0B+R02WEn5p1l3
eL9EInLRTk0ecoxFyG6Znmc+kiFrfCsIhggflP/UiVtSY7H8UHv5MfOlNKhHoGz0
FVULUIQTL2WXGpiJBFktw2rvHOWTibi+YDByZOcYcdM0E9gTC8mF51GMnB1WOPan
v9kv1WTPQLbJ86EjcTmzEl4JOm2osbuiH7fiK+cS+TKqVB4LHHpeh0WMJvNE216K
r4k7UalT9sUzRdUfUG0jjg7ppqXcOVthAY6pmbKNPuEIMVdu6UflIwPaiaMwYLmd
IJacniT+rSpvaCVuDQKf4+Krw1nRwLJ19JdRXvhu6eNWYuOgza3lfREx8e5bu6CI
fTV86ezOX8kJNyS3fECbieBJDoVXb4UgBN3t50//PYmBx1M6R28A++1HF+mCiifW
NOAIIn4Ie41ghkWFIyvp1ctuHe6kTPza2q1SEFT16D+E6lVMeUAvcSGnJxIGMwEF
yo6nbNCeLJp3EMy+6VskMjP/TVa5ZbtkpxEyo8/Ok3b9AWPtrG9UuiBFXSOgYPaI
7kkJMn8ahct8xP4mxyspQbiUPqbekTwUddmpS6tl+WYklgL8TVSEJrspFikaQrMv
Z9pI78OMCg8xdmE7FEqYbo20sH7hH0Urvcu9GQEvYP0R9IL97serzbVJae/lMQkR
BOr1CZProhN6fcqoaetgMnHkImHf+FJSvE86NlniQRMmLBuLTYWgf7tUFLS64evY
dk0zlImOpb/dACujjdID1KPJtrlrODJbVs3uxhdOMuJBryp0qwn1iYHNWYUKcIzL
hZQo3LZzy6lXl0aKY2Wb03rJtDlGRSb37eKu0oKXVxyE/nAPVMvUmUgMudf+F6DS
klsk1PZabg8yJSAkVK3JjEHsN2iWoBYAtLbqYO7CN3IgnbqsSub3hAWxCy+vPSqA
DWPEFxJ7o4m9P/NIrGdpoD9b4MpRbLAG1qjVCe+T+sRUqEw8ZlKE2CzT7m6cPJTA
i8t4ogXa0zDFMluwopm54j4oAorTvsIAShtV8aSHuMVSQ7gz7q7s1px55nNnLuY4
qR8VeQ5pLc/WE0OWnfNKLq9BjdRlZPyr6bIzZn2jVke2s55ypjFCvL+90W9IhPbh
TbesbIrH2yv+Q8+AhEDJ/0GD31eX1Bh5uuT7TJT+rnphm/lBOOpmtrOuoBVIIN4c
beKDwAwuLss1zP9lXcNeeLn7w/tCH2eQ6FkREv3gzfitO/fsqzF5CfZJawc0St9h
BVW485ToLRvaBZ36kZ4gGNFQG9UlaTIoO58I72carKF7zxBDZK2cfe10lyGFBJqV
XfRXiroilhkeDXwHi9eNi3G3XI3A/ZxDko+VDSdh2GALaV88MbWMqbwT0xNtvphr
0B3nGuTadxZBHTsLZD+iejOVRtZsIeDpVIS15+lAuULeUYtEiwHCw37JhD4SNPS6
fX/j7JUnGRuBhoILF79LIn2N6Jw3s95WHc+08wPNkNQ+mEW2yqsVS2usC+1NEcEY
msORO6blIPOdFWuIgafg49737idCqPr7wDspdZOYGouGviwjC7IkF58dc/cCgVIL
PXzwutBo1AxDCxoCqfIGdRNv3yUMfryMcMdfMqZUK31vAvFjKYeWNKQzT03RnFZI
+nU5XqFtn5BxcAMFHKk9AsqhDnN5Og6R6YNdOza+QEBTlH3LljlFNUV8tX3LzLyK
zVv3yipowGbyEI07AgzarKQK60IZqoQwwY+y+7MlSrryq/vjJ6tzWZwos3x8jIcP
a6wm7LprgdPu/AT9pS/Kq37roIm4uP4esb+8vJWJXQ2iu2AznNNC6+hSyFVmu3Re
F6cprLLZgp50NOvBOrGRRlTefyQ8LpiCPnFMZEltJXDhh16d7OK5U05fwnAROyde
6t31WOM/Q/t/88ySEtxGwbc+8qWBwrYGPcceaFjDC7cAUQDtvWHp3Eqgqjde+lLD
xWrCRFLqowkfEcU7sIFiGHjpptxf7xWhXpkfKtUyNRgKnXSCZTs3mm6uirlmogat
35UnfxU5DcaJ5FpGOoquzl7+pWhJ/mzeX3o9RtyR0jjLnzKmqBw56jhjFuVB6dnc
cOFzorhQrMf6K8UnLo7HkEOjhbxsblvz9AhZC4+fW4+tJ1oUb5uEwlFd+EvNWr1e
y51tk2asxur00aCBy0RkwvCKw4jdD/09xF3ndtCWGmF++Fg09J1O3Ngb2l4Wawf6
8mKqm4SXlgqWcp5xTXnlc/0lHmEo1GgJ7dtz4OGQhQw3mIQKL7/VcJDdJPvWONOC
MJYjOjWrkSbxIncd5m7saSKszOwGqVAqbC26FUdAmMyknp9nmS728r3SEubIkGQz
JUwLxRQq6bA3IM6Xel+j4CkYky/kK9wO9Ugu8umPah3lvZnrztbza+2t9PhU1FFj
dzPZEaObW9WlRDC8aEq0ctEFGXFdA20Y+wCLa1pFJUgzsSpykJJxLXad399Uf+sl
4ncyTwOSEYQnSoctgdHCTvor9jPrHoCpUVOE2avQya3SMEiLa/Fo1Sw1q3EeWdLG
RMyVIznfsce/+iX24ZWU7+8s7mNo7ffEh99rKEpFQhIZY/fJPckwRjydGteTwiHT
snW/q7rAoJC5zsM1pZbfEG6FeE91LxQG3LGvZ0S+rATJIbeVrAUYVaeVS9a7RbLv
LbpkIxzoGlKIaEX0rY6i0Qbve+JNLalpDZr6yPxgmSviJ4PsrmkmATdk+FbZZ2gc
HqgIVB4iVvHir+0NvvJskZSWGoUkjtCIxJEwNFkImjKzAouWTra3EyJnCsjJhREe
najEZQcE7EkjBCCrfIikVlY1fhmoqLT3Uix/t75eouxDafeW4PxXnAy/0IMsZ+oI
zI3adGRh1evR/ePSg1heHwoR7Z2akBkkCL7SzZZ/MPuwmfF48d5NhMow00wJhvXz
WiUZ0F0/xqO/+X6mm4udDrhfIvYkUVgUycugkK1F1J1Sc4Mw03uVmWRttwcqv+HT
1gqqE+9Rllk+gKoVWtSttf/FO16H4Pk88sietFtEyoQdFkAOc9muJVVUSExfzidn
FzyqamjiLkaLfF3E5wpT9CI+q5vamo3KWSvhvrQTfZ2uTdjs7c2CB4w5uybNc8cJ
3ULhXjLxc/xMJK3YrmribtwfhxXw4q+43K0bmy9r55rb0aW3s5hlifFQIF5hL8gr
5W+mAsunUpFNxHc5PwlYyCAr4/P8gMTwus83vyDzqd6QRGItPSQClaDj+C1tZc4R
xm+JKyhvzDSc/9XJz9VhapAcrGMVC9y4sOKAMl5VP2T1/1AdKCPEgnDDTjwm88Lm
7OkBqo8rueEJHcWiugDBGDzC/uwglTs40siURg3/ruEb4OTh0w0GyUcozTVthUDA
cLpFbwpDZYi3xyioSlPw/EkAonbG0ShICKGJNY3eeMx4Ir7brAC1/SAj0FxeH3K4
wezOp0ACI7s2dSR7ismZSUyCfskz7O5WzNtzasWYSdd8HikfryS2f/SSbEKRaVKw
uofs5kvLY/ltc0eBolKrUcPdp3dpCx/hvAfGWTJ4I8n4JgxjcmBHyWlhYOIUpDsV
CO+xG7XI5w+0JzngoavMbnIO6ZlA8gWwr5rsDEtiV/6F/O08TMNLB4WxXU6t+EWs
Baqw+HWMHpCyu1ssGurLpRMHbqsl4a0mM1tNf7t6MdVRQDC1RStq4CtI+dbPDXl3
g2/Y74zZ3PiDOoWUaNri80M+BODDzvo8egG65pdRGrlTWJ/ZbjLPYTzH1sVuAvzk
fLV0zFSd6H3nDOFImhNwRh8RFj4UOQp6Bb6CEvQ2A+rOUdH7Ft1XQa/Oi3ATmoM2
keMHmuLIkS4vx6vAexPwAZdxmHsCgVxbaOju3C98mDhRKSwqQz1+h6gPFCZxDdqS
B0sN4DFKyuOxkciNq0lIZv7m6NLBEMcuLfoNOKeMby06E2nFKy/CyPv0z00wlJVG
dOXtaeGf5PwIESErlGvzC8j+bO2y5SLf47lJ4JTBm71HqkzDXoBa32wk/gbCtC0o
CSt65GbCH2eseO5Xdcza69oSvYtDJvg2xwOHq9mc2eFj18ztg1wXAPq3LhHx9htz
xJv4ZdVOVinoO8EKZQhwQhI9O3jbTLeM8eCh0zSCLnYmu70kI3AVmDXhWfNV6Gco
XJaoW7eYxlakzEbOFk0YD3mbucBmIq7J87aiAcU0gXgZNUbcRxk0qRb5ltvoFOhz
EQW9tsHMnaLaQAU1pB4GpwXaD9yk/FHY2xevFIezVcx+WOCugHBpqOThjihC6tjS
TPLyH0/eoxEPpGMqDnyI3N9PwxGPt63NWyjBmZ2qgiCbyxaDDVl1GInW4vN8zGaD
XlnK7TB/PiYdl7V1qr7jmhR8MHa7dliygR1NI8qt9EZ0/ytqoZ70VQLrO6ni0/J9
phlToPBhBiZUKnfXEWWPTGU6N4LSFeqxNzVqwkwey6ympqWib/Fs8AQohgR7/7NC
Jm30D42m/6PivfoCPphXb8hlkAqqSiZ1XXsIYyv/d5K/C4SIvsi25IkK0H/6bh4/
2fpwqPIsX01vHqxxIob6QZ/PblkZmyT9AHXxzA3/vqvpC9eN8lK3QgqAfm6OMFLp
wCanNGlNvBHviMlhYZDJPxUfqOoLhAdGs6/uljoKWHzrCMrWtidzRUx0vLTwfk/i
wezBdtHr/yqZWKltI45o/cmTY1uEfo5s1uBpYHtzSabp/LopjrEQV1i+cpWhTS8R
2yE7xmRWqm+/4lWvHf10f6HvocGY/U98ZaxX8ZT2SE6CPqzDXBK0Af68MkmUkYS/
OC8UvEC8dWp9fxFvQU+BzCp6fagHTj/26vu6KtAq6YMdIt1Coc6+MHYinfJRWZ5t
ySHZXiUXchdGwz05wCgBjh6sBUNVHwhxZyy7IZyaLREvRJ0NdGPkwevDqSR7lM30
Gy2QFIh4woo4sVlfR4FSsJW/BsE1Zq+NmM6ERb1/DU9DVmWSEOxWmWRLsrYnAj4r
Ia33OLx0SVtb8X88M9vYtWoD7Fiv0XiZ4w2WTT7nd6DiWkJPhKMpo66Pk/51HX8y
J6gyTLyvP57Y1VRseobS9C8k08cKN/to+tqH6ilNPY7l16T8YIx1B4ig+8Bb4pXH
qFc/1jJfly/rsPd38jBr4fD8yKmHOwtB9l6eEenuNFeDxDPuULPOPxQK7qgSAqL2
WEYZzyixQMBSU/2TLlGYbK1uHlHS9oLEzrSVWPcMczcb4XDiAfSBm1OOooh5jSe1
baCjtuGGd9OvhimwetLniKhAoZOh48Vvo/r6fFtdQkPIqB4Av2H9RMxuCK2N4lC4
pOzvQ7qvUmRCVNgJXkVO7vvh8hqFeJicRZaQVJoydpyUnYm7V9ZT3D71lwVpbbfn
bKhN+yP40YU6Iy7bN14oOTC5yoU+y65y5MZsJQl2e/Kas5saoQ90bOfIWXRDIMH5
851MpOQ8kYnKeHg4Mwj/QwYtTl7WIk3daa+KqXfYgZVnzN2Cn95ngheTTSViJukK
IoPdoSIBWYdIXxZ4G5RSK2NxIAH+v9OyGq9/ljmatF7yg82f5ow0uF5eIrg1CF3E
KxsLLdejeK/T6cK8/oXB3mg71onFN+04yNs3j++RXiSC75swQgRcdBTczUUTVPxT
ZbPsk/h36EYrhy2cWQarMbCny9vDvHPJaTi2FgR0ZfDzNuuQxFZdSYAXUE+WKC5c
lyli465PvYy95GGFiOkfzoEv56oxyyCVgV5AKBmBU40QR016FkPSHbgInOuaQInA
nBtxato1pDXWQ/HLV5lsyVlpa0RXKbdy7ZPh7HQbfx701Vcvd6a/+yIE0R4yH0vD
NPcLMaB0sMrN68Wqk2cFnIYpsVacoXVe7F5tT91fVDxib0qDWFkoCY26gHpXOXy4
S2O6pclrcxWHyzXaFfAPQHKxurxBX3T7znVbxLUOOw27dQbPoIB7jWXQ7uwrcxgX
ZMHHCoMjljIn+KU+27M1GG7YQwObGCoN/x0xcQuUElpBK9HkoqNbvmSwgUHi1FDX
7mqEyZPREoz9dE4RZbYdQWraZEO/Eg0OfTcvkvp1h0sBSnC/2moyjyC22R9gHwtz
1cRCYxDK3KIByL6TLnDDgN+OCosEilGiWcitOhRGCEl6R+2f2fCDSJBt3mFKrI3s
XjI761Y1cRzKjgXsaAHI8JMsLVbsXerYNJ/9110WCBpwmSOTYPu+IAdEzuRHvMm+
FLPkj18/U4M8w77rlTPaisbNXKEeu7elBTqA9TpMGYbyxd6UxCBj5sxBSBpqiY+A
RCVBJVLEWS+yodbwyV+KrcdvBXsod87K3dDGS0wTx1rl+FTW+xdJJ3EXhkPVhDVR
x9JB1dtLkEkljq9LfwCM5g7nXkk72whkA3wr10nRrXz2m5oFl2FZCnBvfvl4Bc2u
iJG8qg05YHXaiIbMJXzX67hL+23KS6hxkONA8xERKUXqOo4Y+AIXXtbRyCa5Eg+h
ljaOFpoJc57jfptcFYsKVy/EpgVYfk3TpuEUr5yFSG81+pON7Xon73KUzTStJ1Wb
r/pVZQiavKhZxQL1kWXnbkYKArZki3kewATN+LxCRa6fZAUwPUrnOCrwDDiVH3ss
74tUjZ7U8tGEtgcpmvoIeuxVGk/zpuECS3i/3Wmj67YSAjtzKwAYnrWPke0OTzTQ
xXsk9xninP08e2cxAKwj9jZRzVWAJIf6wv2W38lBvoYze04C0bPVHI81kHkHi+fU
IKXg9ebXcrSqCMvjg8auymb9M907Nq/qUVSNKGtkugl85hk5xK51WF8tXs7nwk1H
g6FdctfqWyZw9TykFMeJGPymjw5QKjhy3frhKCBHwkB49osdGDWv33k01sVGfsOF
ZJreRiXSvLNvUJP4YDlMwt5d1Gax7bYelf9p2ECAyWW+1Hbk4sN95VzSoaC/0FdW
P9BMaUEvWOmW4D0HJ+Nu1+Ng0jnvQU4UH7eMZv3HMayH7hHIynnaRQ+F716h7Hxx
XF3L7RqBUgsTrKzAfTXiVg3MEWTLIf0kckoWAA52jB2jZEG289DzOepr35s7LHGH
WGiv3t62Pu5BVw1dNX4Vw1TPa/kNkEuKfx5o63UbtwXaUJkttm4vIPqidzQwXEZO
9jvamJGxiR5CHkXEmUUunPAy8DVbR22tM/UNcGXrIE/8+K59C3rl/LYeeVX7J5I2
B0x6BCuHjeCPOb7ENx03Njw9OS9fY0U8/wsZUUP1/P/n4z/A4usIu6JAnLKLhvRS
RbGO2HjZU/9nqayqI3PkohkJN5yGWNmcbVrPvHpq3irirkwgTbZl5ebUfctgalpu
NPvT+h469ugQo22oRh67dvpz3YZ0WSXW6C2MWl4eU1XEkTBq+76h4ZHc0DFNpvUz
+4gPf83j4UZpDfp0Pp94clr7hlAEfIJuMAttOUqQew9y1yIE4Shb3EluLnK76zy5
iKQwxVjhNKVUz5NWaOER77o+0913a1b/utbhHcWGlkULxgJ+DPDlzl/3jo7Yk/SV
+MjS50QOr8WMmvKirFhcN/05BPck678YCTj15GII3lh66rc2+lpmpJUlgTbpr97a
eLc/Prq5lthPLfxyKToSnWD4Es3vd5/ZljkobdzgPz5xNcYHyfYgd3RHWu7+HT7w
41euY8xz7zWxKs52bVjBFJiMV+Smrpcz+v8sLkFb/5vXit5VJAKUjK1C3hTPFvry
y310+OiYY5rWm4+9n57lfx4ufr0ECVfV5vmhEdfopHB/n0cv/mtthETN3T9u4uYC
/3n8mhZhaOWzwsW9N4ytJCmpgMvFbqTbudzIsAWkWbIzeMP2FRCL47o6AWC16J4r
7mP7xihuY8VzObhHfgDCxY2XTWi9NJmAu0cuDJLdkQXSM19sCatRpAEiL32QGsn1
imcf7NvlytV7QiqIXX5769qmDGLAn9wSGwS+V/vZ+Yme6jqLMPCc9KtMGClwBDDk
Le1TeWKcFBrBrWvj6HfuqJ0v7BQVD1Dj+5zxIQxLU71uoyN9HKVsMkh5YR3RRXyG
9CQqtF8GI8c4q3zw189c8inJg5VYbjH1HH7dvnlPJN5NmINHiMVGjanDu/skr+gv
PeHq9QLX7b5R6FyTb59lrGDeCYwv46gi3t8/rQ1ER4CjeiQbceV6nOYBnvnhpY7F
9RGBYb7tJ+Cef4oh3RdW4rfxP0eeJjaH+UKUJskcOFgYHH717t4fdBjHvqeYN0Si
IHXOK+vPqNTYqdEcayZ35Vt0cKh88ByRvgLrx1od/LHME7P3VzZ9JMNW77nc+CxF
ASXE52fprwH5p3ysn+ChcITOSTmW10bunOQbEvgb0bwO5zcXac8ic1nnNa6+CgwN
o1/exvuVjlGkTysBk2uiOOvc35Rf+Iq4ZbdLDu2d8JEM+Svjoqvqxup1UT80+AEs
H9pL3em3VhxwJTSMQe9RM1Iz9xPyRXqw2NYVdwHAnZMp4I8rp024XpspMByuZ0Da
n2iPU0nAE1iJUmwtgBM62mHAt8DyyPpS3RupMa0x9RCAu9nfPcroj8C5uN/iDfSD
gVb7YMRjQkdYUdrzFPFSIh7EDT2qb/9X+uWOCWk84GdtzPwL6sva80o7yuSa1m4n
0sBjN66kCM+w2Oou6LpxnTtX4/vJ0eYAfGuvUSJDROFTRaCp3Ak98MyDvochA2mk
/0fLjEQuYHmhr/3rbew6i3uerxRH2xCfM8uOcIXPQraVzZ0uv1J/QaKCzMB1n4Mm
iDgbdpEIUOSGM/PMKC9Mpkt9hLVyP3/nPDEetYxmZCgPqhpVY9kcDGSBAjVQymzh
ap2PNQxvs7rUfcwnF/tY12RdFyyVdlnPs0pl8tn8MQxkSgrUrPWTuTU7iwRddfoP
E48uxNUrUeaOH0jwYJIUXlt95pavmYzSLepPVLfcAzJH6vfEzvfWfo8AU70YsHek
UAFNoPR1hzx9N30I+AlcApeZnrQCBhSC3vO7/SpDn0pBiDR1JDeWC4W13MC2mJUw
vdwbrUPn9IQnomlq8boiJ7jShuDEj10NrBChqjaHTWYPDCIj+kQdu9C9qFwsq3Mc
7YB/QHgEftGMQeWRihi7KWdbn0tqWdfKKD05HqFUZThN3safdG5Vnxf2d7VY79V6
cMpdzpsajOkZWu/7SQWUH29Epncg+rwefiJPsaDsv5JSEMZgZN1onrLm4vYy6H3C
QyTNM9bGlCpLoeIV+42l9/vLq8mtvsSYo28TOFbZ/37RQCAn45ttAAGCyw1OGbno
Y+AK6EEq3EyuTC4wdWaRgCIp6SXulOEyA8Vh3lPP7ZKolchabtojUGeyImpBjEqK
oIB3/i4IJzLAUm2iU+dPCjlk4dhpyt7Py1EWD7kut6isfasYO89eNvDNWQSGAAYN
zQVmFyaSurSpgZZQCPPXu/fcEmrngo6m7mOaZLErObVTKCfXzGwSoEBlPkZqWWON
DU7bcdOx3lPSFhCnQhb1u51rCFDDAznapjZWrogmEKrMCE2StR9O8Q6nkQAdvdNU
DhbQsR9o9VhSeQDaGifV+KY4mQeghvsQfH1hk4Ycf+ah1hA3vbT8DQD5+n5Tfxi/
OxEgMMerXoXoFq6jvgw4X1b0puYpM3U8plQJ+GJkH38h/OP7VSP5EjPf7A6N9cJU
t62ouiMYTko9ak4DcKNf3cyd/8J6ZZiBywjgITfltxEgPar9cWpGftcexwwfIRjV
b/tCReAd40E+1fQgxgARUmnTwknLj88hi8E0ZDiYuba4Kgm0pHoyFph1Y2IcgnGA
ZCfAirQ5CfEplCEfUasISlu0HM3+Rgeyx0CYLHpz6WRuoklSq0xTolaVev+qvnJf
Z24iTu9b/Leb0kfWU6f5wKuVTzN6q/dH5ih+mbSW+CNqlpqWuJsEM9AFn/qbgGYE
gv9w6/mctQ7yvxU+f2zndmSpC/UwzK0GJ01HhJ6jyGgfa9QoY9DBuy6npABUlyTO
f3A6My1+xgPIcHwSJm4NCveUE4Ofmik+6MTR8p3rglgGowtGrEidIhGicdyz7P9E
DzZMYNLjYB2PxgmSyb/3gOPnfHKcZJMQd/9O+Kb80rRda3W8HLP4tj6/f3i6D5Y8
TAKTZh1XaiJ75y9yc56DxWDCND0Ci/JnPfLWzByt8vh1T2ku1gNLd7hupHGnyUzN
2+KGfs96XMxNnJLVu9PyP593kTS26JDgo3/OkvhYVRjzzm3N+IqLEls5C14IkD+D
DE3e0OdWa65vIPeUaLGmxjrycnrAtO4F/LuBoJ1fwfe8YiafZev0uDXPf7Dxqbfx
lrAOMEPzuXact3PZIRiIsUxmPLWjYaUg1pum02+A6sNIsxbJkKrbw6Sn7nYLo6U4
BcxEkMccNp/nkZGtKCFo7m0QTz4oMvzuD/nJ03cuzYdtmilkC1gRJ/nfIHsKcTNc
HWlEdBekqeCp73aFFY36iKPjvBieqADQnpeJ6va/ZaWp4rukMr5ks8L2I65YEHDi
BeSSR5dTMALebVt1mDBIoqRMNOEoqPfRqiXrwmO94wOyZalyWHmskZbywp62gQ0c
sZSCm2Cx4NRGYSITlg2TuvwKqSGBJQ3qLzLpLrt04ko=
>>>>>>> main
`protect end_protected