`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 35344 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
LfLaKOw3utJqtz02pVdKf2iSjdThvHkeLtBEZ188g39XUfhi562igqDgA7t2Q9jv
sWIxnLRFcgi2FYxmXAKlQ4w7x/fOJqQJ0RlUuyjD48r92xvysHc8+9m/enPtTLiL
Ab2Gcx9uzrnVYIuZosm0boIcNZ0U1BaG2MGaSpYTS/qh4opVD7f6B3tlB7hC0TS7
HS+QNCL5o/+tZIPLeGYV40iEsV/9bc/U9pYgjJOfslDmPk5sr7yx7MHX06UZPRgF
b8vsCQ9UasVvwIMgJlbQhB3v2B6l9dg+R/ZKm9S3dGGvOgvm7MRLD1iNEt8sjXVC
l/WsZx9XXQdYEaC/rmz5C+B2NdwRXVRbTqCh6GNWZ7NjQkJiiekc9LG2jtYX+Xi5
EP8t6FSa0NC3LZehR5EvJb8x0I4c5t6p4OjF1La4qPtmPY36tEj07PyXuVppzVdh
w/IBEMV0AgRHKzjx7PzaoEIXZVe4zysQx2VTGAxrwb3Q3PJpoyc0mg7sPw2bglQo
JWf2VnTD+pcOl52j3xYS1EBYgFSaCwjKRJVCWnAA3aSsoIj7Q4/ATK8/kX1BYGLL
3wiSdZEvGppdknTPi4tQi83I+9dycBIAlB9srl0ouCNmwvyvck76KvvTmo+QIOmZ
QB2Hu/aS6nVxrFD5tg3p1ye9OQgcJl+6MPdirZZII2oX5rNXm1xYs+LsJq1Kq/vz
2AH/meoqk/yVGmq+vtl+46YylFZKpNh/g/08xbDhq79J4jceDdnIqcJkE29CfyBB
+Y3wbQw/W0Pl1cZ71f1gfbadrYmrzI8FKWZJV6wfYcAd8aoQwVvE7DsMMBSXe5N8
ku26mGe61ub6CuQFc1Msaj7IM+2GRi4ov+oyx+b5S1U0d4n2I9EmijApluTCekcU
gCpFIIJU2zIUOuIaXGdGpXlrTVgukBm6U7nxACumnb9/jYJ1+f6TxnMaQGerRIbM
sstsVcpWy6wMXhCRKuMwSwHVzl5Gk8ziBZTWgGU7iwmkUv5YLkv8q0UJeMWYpBsa
/sp7CQmuxEDT94NvKnVjDuA6wS7ZAL0C7XDgyVBT6nhid4Xa1uA3Pih3VHtUTozl
I8rngz27Z8kh6h7uiPZoJWj3NT+xQSPRh7qmJHKtZFiL3EeQPVtyS1L4jf8W9ZZM
W8ediH1s89ujqasXwvGaP1tMJnhAkb46Y0KOTIGLdFSMCox/mhyIjIysx9jWVC+O
4R9lmh7sXePgx/M/AcUNdxPd6DW7YqpXYalTWKm3WL3WbPy6lgbPGhCOLqlttMIr
vJb0GzGUKWld2akzfT+Gd+syIfJbqFuYE1Ry+aChBjAfmhyfvZv3xssp+pRMZTKo
IuzdH+dFbrM8envX3zTIVQpv3knvXKrYCvz6Ldkv2WUvA96AMSlkALwFDGKx5hrt
Q5mxLD+r1ZIoZ2OXyIdJER9IYe+kSZnwg9f/Dp+ox/CMSnpoWR7l9fax4AnQV8c2
o8qpGE/1Vl2Z8AOA2D3/IlqUyxor7/uSZujmU6M4W0z4atq3CdGe8NxCMBaQBbBd
wiANBMTrviiqOD/lW/JtXxc6cCFYaf0MrEFuJi3LGQxjyc5sVzd9/KgxL/hE4fUG
dC2iLrX/byvjFmv0fjWBPs7YO0LDR1cZPcI4gGHOHQwyTQ9NJ3RF7O08B1XmZY+J
IEk5BHEd/5MQ6klnfUd6SP/lHVP6Wam1os2FPAg1K3daWcah0mFWecci36BbithO
5LErH/SRM+gPRpub7VMS0Hn/DGMq1N+ePJV3D4DevQ9OrdXQpo37j0OHhxbUpEJ2
yuSq/ooQB4hhLUUriu+fhhB6zAKeTaCX8S5dLuKsv+rGh1QiCL3O0I740OYgEJX6
2WbkkVn1qcQTQUGuPMHQau2vifbeKBRGXujKwAkwZJKG93s+QIJ6I02e3xRja1mx
CTF5LYF0pj6CXUaGqgSjlv2G0elmfbnXpjYvtBOK60vRot6C6thD9BjSkgKNj3P+
uUD8ZpejIDlpcuFOMmEw9F0JU/hN/EzM1ryNhG06OAdCgW9MgZcB9qG8ECVj5uKx
OunhfhTfUBTbG9ZelZxnRVC9ws1yACp9e/3XCsKuZU/2K8bd6KztBm7zUZGWriaL
HmLT2/a6nwDXzqLDSK0SbJizGkZu6qd96TKzzUd1eXlmpo6sinhqb3Nbq1Q0Koz5
vHgS63mvDB3hmZfkuCGuQx+ykwbx0F7cDdw1ZlO07XAGLgY3NIbrGnc5tk9udGmo
b89Naaf8tzyRdN2kPQVI1fh8L7tEvSQS5A5AWhIE+QHRD7rKfCO2N8AdjJE3KhvK
LOGMwOqp7+zhT7kJ8FytkmRireJKHoMArJ/jyLMh6j+ijU2Q6HLj0SCpia85L4Zz
omJJYJEAmIdgbDbz5MShslifuh5HvwHGEhkpPlPNNugN7UMG8K6GPvH6LpvnKzil
cd+Bb/DFj6XTE7m+WFvqE+dG1VoYiau/Gnu+6jhi+mv1P8gHBucyrfq3KVQzFv2y
f+EDTXq5JBm3sVHsnDRATSCMVD+2Bka4sT+Wu4U6Y+7nmJ05+GRdvyxH7v46JAH3
HwAiWGoCYBIBzCzYE5wQsamr6t5c1jVRMeT5HAC4HvEaz3tOq9KusVliwJmt2QUe
vizO5WgbgTtmGAniWL86vfxzXDgqEL2avkzxu3G6arIexGCA1ppJH1xJYlZ+OIhZ
/HOO/jQCoouT6wDkwdbUhIk96HCgBVZ63Z7kqpoDluQXrG6tlk9vo6awY5qKM7S/
FCcOOGmTKMo3FVSFZyB+tchOUK09cmEFhNUnFM6gI9olJbktOBWqupsd8YauHsuS
3sJ1kNuD7Fle2hM88weryDw8yGgYVgBnZio00A0/moudnjjh5vxKP0GBLEyOYQg2
+6lgWTzxj+vSmoGEKODQVEdLpC4dpk7TPy7ouHxOXpjtsgFK+rrgF5ZDJ4XDYosd
RPpjlRIfILIYwV0wdk01u091OrLcrUuT8JwA4mrrwMCkq9GG8bxI6TCAYgtXzNu/
kfo/NVqBZbOZcUak4DEDLYBiZS4u45gHikaF8n9lvTkwehO36BsT4TddvipQt8lT
KaA0qL5i1hNjmpKYsIHNALawjKcUvAqjQSw5TRxJz959U/GgP7U39Kcwu/UzzzxX
9e08iQ1T1I3YZvCzB/Kx9PbEyuWzXEhRMeebXEoVUbwz4nGY54HYEcJtrIE/Ct7E
FqdyNUZFFGrh2epRcietuD8za680fAuA9mbWeYO9QE4TGaJiyhpgi7D8wOvmbviE
ggjixqxM9Ok0uH/JTUprF8HWYRoKHUCY7JydnmYrauE6tZXLJ67m5UzDiS0NrTMp
0fXN9MHhB/PMwwgrJI0P7lR3Edk7OQH+v75Nb/RS3U1Y/CIkNQ+icGS6ZobKKisO
S1uhbVzQ19sSMhjseEPXnpAXG/VPqUw3Od8X7nJB6qg0cwda1VFYnxBXk+e7wNcm
UQCLwXWCKzyuZqJbavXyEPYsQz31qO+LlxYrpJmFZJAUjwn6585YLnzmmnjYSDLw
+8OLQ8XeG7p4CHUk6ch0aIUN2MzuhnEB1C/7Ml5trusdLGuhwaDtG24e1H00bMgQ
hL/zIK78tA9hIvtMQVY4/HTdRMe0QpFJp4DfTVn+nB5kWvJOX4TdGCO/r6q7Frvv
VMEvSiRc9mKmLX6MKUfP8/Exjx3LauL+Z3UGacAg5dD03MGZbgqu1lTnZmAhqQjx
2Qx/3r+oMQLr8Nv2amcA+C1kQuFLW2pS3Xo0EPfPiL7sVlnieIbu/bLNborusLby
Fl9JgtwnrkF+BK/H5h+rkwAKFSihlJsr5+jFUeWU+smOfWtcHJWUYACBeeuzU/wV
NswEjgsfqWgptCSDf+khuxMMirnOeA1kjkx1cFfGp4KbnzDYVlt+PLAbqErhEUjV
zJ2rPqWa+eKQZylODzvXhg1G1Wc8y5Xd8Or86FvucdVXPyNCJm1MdC82unsGwCLe
LY3xgW/JwMXWqbIHWBybZWKgb6Kx5x5+GfEteSlZe1HQW1GLY7uZOEwYfkLbO+X1
1I27FSmpCz1Rwj875asJqaCWGj2msHv5M/ReSHtp1i+QF3HRxCSNCjJwkuil326Y
MhknF4Ifyywg2JT9cr/cgYsNO8lMuOb6KqvIKGeSV3u+s8zlcjI7P0wgt5BRl9vp
SfwRKK8KDvgLGVcURd48HfWufeXZPaGmSl+rrppOx/clfc8PhgZP8XZUH4lKHcg9
gLqZBvQkZwPgE/+vWPwRhILMDpHdoZ3gfWnka5CQohRQ72380TrIpJKVpDWB4+/l
Xsjp5QNeBM0KAaPepxpn727DSjHeCJSzZauxLKAOw5Mg64rDFELIfRcpZEKukTog
gibn4MWI0tUTIrYKGvZKPZJ4FATmS9v3Gtwpf1S1F2NNj/R6GPG5xFk7KDsrRzvg
36ZqD4IqEdJT78EOS8/UYrhrM5IcgRv2q2h4CF7D2JpmTik7jwew1yjEEQAY5Rnt
AmVYJnaNISZ/4cR+hEdY4jZPnqcPlsa29VyAksxv/K7TFlnXKzraBYMH3TO6TzoE
fDigt7zg81h19ha2ZTt+yzt85ZeT/IsmLt6XlniOdFKzU8Fiou8hFRDdp3yYbkjG
8O0NxGY7LfkRL5r5jKhMwDKJj+P4kMfqC6sJrD2FN4L11Ycvzn/UclRwcBcrbOyE
DSFvtO+QsNMc0aHfVelhjcICKB/l4L3TESAQc8HS5L/PhTj8khrAt42e/5jMGtCx
8Tef9gPowaIZ6P5j45tu0DL2IroC8XBvcReXDqKGv/pLVEfBeBnG/UYegjnDHc8M
w2Y7yGlvvw47DzQ+0Vildv+s+M2OjbC3hJbg/asUky99By/dDTGz9CDeI3n+II0p
JiGgaBDr7hXrprl5kTJENzQL5aNtKGuUPSX2Gwix3fZFKmBx/E/rV/odTJz7u22K
208wKIZ4CDC9wFeZI5+Mo5zgMrh5Hdr7pEN9XQvahiVyt6mjIaxyJ5WaY9K0/6M6
lxhXkBIEkNgnCmi7aTphWJxIBngPxB+jfPtO/ja49TwISVag42JkdnHQaGthlpKK
GQ0B4nBzrAOg5ckhNG2bRqaS+3BaaaenVnbCr55oW10mljym94a4MwVHfQ91lK4R
y9YuF/MmFDGOwmkxmR/RzK39wxtpfFZuldZEFOR6P2qUrCDG2K9TE1EvkzMonI8v
0YtJBnu2rbZbTlDzOo10lJz+sD+lG/7FvPJdr5C3Ue9ZDJcJ9mSvz8RRpW+5lNjS
WBktwwPm493rEGrAivH5yAwbSd+cQCIVaMDLBoE7+EIZaZyCka90nL0ig6gKzeb2
09W3RZEnJzcHe+J8qYnH70XzJCj+BbMuQpT6TSe/R6GjterNB3qeRdLDyLQJv8qo
kVka28jIj8VMBXcErDYRrKY0YGqAAY7uMXmdSy78aoGrijCwoSXk7bLIHF4LZg86
/aUZ0C4dnXQF7J4KNJ5TQUUzLhWCyBC59g09Q9iBYMJ3zfEfbQ2lS/kDxfkcMRot
YTNbFb0MSiQRLJLU66mW4yR0aaBUscEiPDekLnCDx1s2s+7eL3JwKagreOfiBGKI
0bK08BdWMAOoV4QjXjRYw6EP8Z0zBdNyTkr03Hk9ORBfdEGhhtALmI6mptBde7FW
cpNIfSF7QPswHj6ymZOVw5f549dTf0+2Rx8DoEKnseo1G0C/vAJo+rLmwPULYdF/
4OVmMj91vS+vMhKyKLYu+U1PgS1EOzCgoTFApQmRH8lsECWVZQLbRoS9QhLaIwSc
v0y82q5gszbOs9dPYuuBD9SM7Yy2VBiL+TTjQQLW/NzigfnARJ+PUtT5ezOK1RXw
iGYBuQ08pVNnce2ZSKk1fqH8LGmfvnzLaI6jeib6rgccubdFlOUYAwkfHBM6OhJn
5Wv4aj6+l3kor0gz111EPRZTmH5t4OSpMIzWSkP4SJHTnVM+71WNZ4A9zs+IouZr
7MMpxl3opHp0z+1UE9ko5o6ju1FVTjroCis8s6RamP6mQL+IXxrf4xeRygYYqdFi
Bg5wY208d0bcxPl+cs43djWEs/UBbQS7QQPMquUlNtf0/NQzxyexGazgxMso11js
Dh3KOBbBaWaaoe/6A5qh7qLZYD/P/Wcv4ZJ7Krhd0HQcAOHFviCxmCRl8hwAMak/
P9g2FgVzcWYmhup+48GOtu8q18uX0d+JE7oMLbQp0J9CRAF4HAoM5jFtgc+EpqUr
EyTjL0GszPN55WgSBVBkl0hmHqpnBNR5sNl+I4ZK+Nrpmtfv0MYm1bLJEBijs1lf
SMmD8Dm38tvFypa8Bsc71YUnShADkZkUQozbQ3wtipPD3ehMwU4Wp3ZPncH1G2xR
/lIoH67yzgEmeBOvfzER7zFmVIRSeqeqM8KtW9lydHNoh8KDdf7RhFXTBIs83eel
o0iSNIvvtZltqyHfISlCBTenxIrI9DKEK5LU0BddxpDtmsR58oXlABU+pw+1jX/E
Nbwj1p4ivUNcvx41tlwuo9HsEp8381LYVrqm9TF7gqYO4aHW1y5ihkoVKbZtJSkm
y7Q1zHENSMfJ5WqiksUFn9XjBVsiy1ab6i3nwgibl8276AYpK9iF7IaT4G+JnQcU
xsz9eWewy0ia//WDrjDFaBB6aGJf/nl1G1IVmyI/cDozYZ7rkWGe2FcMlyFZA+HH
WwYhtW3hB1en584PmGu1SLA/b4s92W0uzc9rHLGw6PMeyD03NzXY3q0By/HlPiiG
t2c/zFFs39EFSQVSmKTbFfBA+7Ojc5hMJApppIup0ZrDCbzbuSNAEBlNPCW/9sEJ
4B5sL1EpjkzT7FUQ0o98gh3gLtyaubxjr1EjHOpG1q8I9r7FMpTUGHi0KYoIzYk1
5E1PVw4kdExTfboICPsMEqGLc87lFt0RZAkOFBVLkRXKGIYic5LOcInXc9lSc04J
x5WHPjeDcd2Lm49EBfrHvQri4Td64TBxRpjgUk4us3pr3NZeCOf0G0/hba7aS+Nu
yJYP7V/F/MRKbMp8M64HKeL/KCSh8BTMSMQ7QM/gUxgY/Xlt+zHF+cW1g+tIcD9i
kgnM1c0TkwOQ2xjsPeEF++CFITOLPJs1dfrbnXxYmIoEjMYeCBv9MMFW5gFuAFEJ
f4Esd9fP6Jt/tqpbcA1U+9oibMJPbUzp0JXbx/N0YPVsciotrym7Ez3ABcBnyPLn
porRaphuvKCe12M0EFhL35U81cwssfG9bWTDdHe3/U3j20KiWYMXSj6GJfuyxtdH
JtvYEDMgxOwAYWP6YlNY8gYZvmRU+ZTnOn6tQlfmpZrwDkieuJ6v9yFp/2fS50e5
zfzOvByGa+BOcrS2mDFV9hzQq0KCKSx9liU0ys9WrXEpubhfZjkhoK6fRKAS8Qan
wNuV3pA/5LCfTfayOReR06qad+UOi0AmSzbhTuhEym6BZIH1o1xpVkQUJgI1GUcA
YkX2nnzfM47Qp3FrpIWA0nlGhBhBtAoBACrd4iFuusydIruV20h1P5bFJGvfYeIv
di5C9AQOanKEGNxGh4H3jYgql8ZCo1Wq+iqHNnbvXnGtOP3Fusb/MEEvskDJ/fZe
Pfx2vHGCz49di25BeSTXptP5Yc8zDcseqWpc4IzNwkCcGi3jCUnqWg+XRcEIvRXv
h7difuDCrPGL72dsoWcWarLLP6h719pkhzLwcFNtqsfClMthBMrEA6fTQBEx/Ayr
qslcJ4eAgb23mVge1oFQsv4YIAz+1tbPS47z8wofGXH9bJUxgn1b9Ky6kxkJJDSI
akTQr/J3KYEiPRf+pEvCbgH1NXhp//i040DwhK2v0ZgypfHMiiXjCKXAuEjqOkNA
YosuSa0twPdSNFgTI8Qg5eZgOk3lHhzWjMdKF6l+0JwuqhLsxIjNoZArBIlRo+89
U45LLWLq8UcK5LJU53vydozKsbeObt+rGuA1yOAlM47K4VW4W2owDTSDilnBLbWj
6/i1zl6wabMvlp4iR9PYzkzOK95TDdjSy1abXTJ1MMlO0Gp+R1tpSOaXrRFk4fCr
ycsMqELBe6VNrZjgekYZPMER/alTIBz6mazBVz3HHCoNhxcBmki6qT05sC4LKQVP
guxnSabhOH2rPy8rWWVbtR9k0N/hSet8Hfg+eDtZkwbl6rObzbuFrfb6MDJiAfci
wMZrwuc1ysQqXfB2J6Im2CbR/fzIQEGoHNfuj5R/A5gyhEOZZSOa9UVQuOOtGjzx
3bW4Xky9ApNBBOIbe37y7aEQnM6VB7QCBlNWdGEv//9SIX6VZHCcsoG0RCZX/WvV
mSM2YaWVDlT0Rma5gYd96a7KtUdKJ/XeElq+ZCrjGg7NJ8Pt+d+gC7ctQ6XgbiS3
peV/F/lkrCIjs5M7eNO8uIofdbXBbq5WEwsuhxcwDSJfhq9RBmHhe3tPL2SeAbLz
Yd65rrVK2WBnw3TMgAhK/80i/rGFGfzlMW06nMo8B6h12RbqNTzBjdv/lc9HRREx
Ie+mqCBMqasVHcuQWiPmSlmRh2oYun1iEM8++rPWUSPH1fBP9YFlwX/0gSw53uO/
od6/Ed3dOw+IfIXVe3PjEHTz0FmHqAjm5Wbf22TCu4HWEcl0c2y2PLdDZY3c2lDp
t7F2Cq5zZ2PJjA63zzgBvvLW7k1TaTM01HXB4nKkdoGNhFSXZpaETG9NNZ/Xq9K9
QOifvxSPzDpkmjCRirlKa7/lt4/WFARNPQC/gR7B/cqLA4EnDJBnxP7hmBYyKmTk
3qchhOUORdSDwRq8h22p1FfxS7XnbOqJAdLLepec6e1iIjKv+VPbFSlO6xWL70iS
W5+ApPnBcWrtPVHDr1IkO86X5CEhbBYb73GfV2lmEnjzmwV6/fWoDjrecAguN8NO
D6c0g2fj9PSbHwGFCzcTaIuwhWZIAw8DpgxpOognrwwQCifyd+8iq+zT/z1cool/
rMTOtbe/m7r5E4TMOrVMKNPT/0iBkr3BI/rZw4R/zlifNk2yX0bxiIRAbLVxO0Qs
5tBcdIwr3tw97crXPmsVXuYPiWxYdNtCeS0mfa4ojaNOff9h75mKB3wTo09IJfHI
J3Q7BGMfyaCGzxo4fZVgF2LqOxq/1SIm3DD/M4VfcVRA3jEZsdRpp8gZI0c0kt2w
YYIB86u4JBfjc7BhZmMx1aZ+3urHpvU9deE/X0A0Iei3dUCLHVpJt8VynmWLw9bY
K6HngQ+kcxSkE3UVd+YgxEEgmaFM4ECwql+m4qPikNJH1rV+eKd9sIzlHG9eHAcx
GuvbXnveAoyGepHjCAYXSvbJqCJkTcgPPXNn2dio7XaaHLnTtE8i7/FaA80htEFT
RcYLrUO9wGx2RPpE13XNe/wHwdiV3QqkhlJ5UQ8RgSvHJJhV0o6vkjPFLpGZ0IMJ
7DNuL8ewxqmSuCsdxIddYX5QbgQyEF4RDlLZUA3PphsWI5o60MExTDCUHVlNzD8s
8xhpkH18xt1JHkQJE1K9KULxfUTiB1T9lpuPh9CKQXvPagPwJs7PrMJR8bpiqZc3
IWqZbghr/AOxrIZYTuiY1rB+pC+0lGO0ThDxyaSSC/8y5ilWRkclXn2htdHL3TJH
ayZT2jpp2wArRlKDXJnTPD0nTDfybmQ4mE2VBRedAIsKp7Zu2+ZrCpt4UJmAeUzH
sk8+0B1CuEwI6XB3Wrw9U1rmdsoyWtkkbZfzLcpf/c6HXv8eBRNbkLfQuGFzpt1H
Bsd4EeA9+2R7L7buTKr7P2R3SqwwUVPTMu9RGO/2xLqQiSmNUFHEGrIIa/kyrdyd
D1TaBiAL6z47KY3fNEcOaa0g8/y5RyijG5bemz3BeHhDhccw1ASY6qNXbsK3rxg0
q/gl72BW0UmgG0h6Z+9nagUktggE1bZcAt1j51+psmIDx2h3wSAWyj5xVzJj/wtA
igWL1zYpFM+e4BC/4WjuWiYyt1R9LR12PfJRQ1WOt5mp3/wNFilHb7iwDozqRQ0h
f7AmRe0VaYupCbHxhCOW5rG1yI37nfh/BSJjuomtWjm4Wij8/648XhtEc6/s7vVT
lvfP+xMlYQAjXfz0ukkgr0lqYTMB2uMaCq/s0GFxSxgii1SnY6RwdGdLFkR9wcNC
9/SHc8BRERVlLwBo05kd/zQQuxZ1r74jrX3OKZPVDb1dnfl/JMZbv3MP87UyUY36
tfCF18Th8YQTmn6vknTWTVn4IUeMYicjokUDl8WAncvJcrHdI+pMNFaLVrwl9nQM
IQN2n6qDK8goxb+tAuX5TsnYKyOjAnvcwGJv44rmzvHfP1W0Cn7U565lfa+GFT6p
tv9wRXiHokxEQLRtQLSEH2Xy0V5ttsjJqIGRYmKyRE4O1COWrNn1IVSZq9RjJOsu
pX5YMKc0WTjaE3jyXxGGoKLmNIQvvJ5BJAGpl4rT1UYhXCpJs9rg4otmFhglf0z6
htyngTq8KGlwxpWKdxZiaFR56B1aN71/4BL+Z3hXH+iNsZWpTWVYx/0U9RXb5zHa
FkDwCdvgT9+FyzcKVlNpl5LFbpugp/IZWn3m865FoSAAyGgKURHczgcMRSpgaMm0
1mg79CWfk/upFXJ+iAft/dJpWbuc+aHQXa8Uk5hlC2SSKuzGWmZvhmRE1Gk6yjLk
mUDK0aU/nEJzajUoqQH42JiyUFS3chBKSnldccsd8CR2Z9lw6bcjvD3/0vNaLkLV
pLyii2gc+GLliJf1c4gHJZqSSjdPp8P+QGTHcfYlnKlExR3Zhp5a6YO64jsHWUSo
S+38wgrYk5//Lwx/dqx1YcvZU7mLLigvvSF1AT3PQKIrSq3mNvddYwprJMMzMjwK
O5PMbzOP2jhn4vkjcdY2C6vQ0Ws1+CU7qUsrqjXbwJ4Ou9Au6TlT8qNqEXjcEi81
LPTGePowiBv7wfFVvmZUNTdwI8eIg6PdUfpoaCJ+7xseuSV4hA+Z5S6Cj8/TyC9N
8WIOeEZAZ5gPOZN9SAiM9GoQcbwUVMo4dkNJv14tSnvVraCYhNv+U95jTQ3M2O9b
yGKNapt01BfSWKXLMszfNofW5ePAZEqTkT/BJWwTR5rbIhlN89Qes+c62ejGyCUY
z4wIoeB4LhFXihEcBherPfUw6rQoW07HCE9rDuYPhlGUmIRjXHke0vqq+t+nNCJO
A0EX+k/hmUD1dqP2VEU9WkqmTnbzrcdIEUm+SviFB7kj3I9ch4W0HMRbWZFsXzBX
erBVBVOjl3/Bkfvjbji6coRfQ4RYhQ0ifs/Y0SwCZhLpfd60FItDoxWpDWUvPPwl
GNwiHv2X5P167dLnC29iJGfONLRl6TNTmWL3xguH+HiESXViIlKTVVVaS+PyrUNp
8BcnORW6ZinqAwpiLwyp4vT5klXlzWSk382LBudaoQtUoLo/yZJqbbnWfQ8aDg5Q
jjAzWf9KzXmzN7ruB7+wP4fAylZA05+xkSJj+CoZD/6I0WDKS6gpYUFmt155/vy6
V7ZYM3lcEs6NVjlFo4AyAC0Yt0B4YFaLywK17BYjZOxOZCZGU2PydJ/j5Mk9FcIq
mh113pJ57qcokxg73mixnoIfl2c6X5U+mukjUub45MCtjlWN/apfoKj3a7w0fICY
Np9kmnuIL5cdJG5mrUv/o1Ra3KlZUVVcem5iqnmpQhmoQXFF7hf6IWTm+TDaMqWw
zAmq410f1wlV0Tcba5AfWs7p506j8Xk0ygEMBXZIiBs1oL6RZ9j5UuiQ4YLy1xcK
bW3+OyOdNXmIZjRcZ0gSV9tMfjoW9tooHs893zQEiY4+Thwa9ScEXvvd05nLMTRB
focsfDsfMDaxVL+YYkGn4dV3MK443NIftnWYPShMqFNUDjYw+F3i0hA6YpP0dyXL
EuF33eHu4tW3oMKlqR9c/E05Owl7uU8q3jQ9SJkoNbdM+NBscU8HRUYnGc7yDFZB
Ym7qiA4RUeTOqVu4XxdXCZUuj2R9FYv/30GPS/3Z/F0naqV7/80nlZnnTZC0n9oR
cE1x1JI6dqOu3wCGXPoxRdlI2pQPF9HSYR9QBxM+CHjaO1gAI6wt+s5wu2Le8rHg
vM5ndF8cie6nex4VAzEPvKWNorCGuZGXWODK7FHHRRvAuCB0PVcrv6NEF9eF9INR
Aew/Ifw0lKjr1gksmNIyvGkPDv4X8T2DMw3eNatgUCCUr3MKdc5vKrRPgAiGW7M+
c4AuyksM1nuoqBnTWCd0EV3NYoLHPcAMvH9BEq8DMdyw4y62WUAP9GJA3rmYXQI4
lp6CexkfRJ+Oa4sTwLPzhXgJmqP/sM084w9j66mdpF3dTwiHhUpR8FuOJg+NgOYl
4kEfeqhJLkeOC3SsNxnDRixarHeEKw8vCzLRdYkvwPORuXaD9LbwPMqwP8dZsh1V
QpKrKbLVw0GxVLUnVcOJVQ7esGQG/yr8PRfACY9q1pa2ijCm0LfuZ7JwjpRRoxom
y9BdPo5SpOcU79hfzU96jRS8z2Bk4VlWNkYqlYDCa6eYjGe54AH+iSva7hRkwiv/
U8mZrj0mIHyj8UKdVcvC9MQRcCtVfma1d7mO12qVfEPjaDOjaQ2p5hvA9c3AbCI7
l08hw3sMhXk5gd79o5Y7bOhLpBmWbry9vz8S4BjWzkYB5xu//ecXFKZR/2i1f8/V
bu30YMYak2eE7Q8TaXA9DYKaTM5DbxbYmkVGhZUFKwyJD0jcb269j2yn0gUlx9ex
H/pvn7UIZiRsiYyl52nl+Eci2CoYcBlTlbaAzhHGf2K08W5UqLQe4PCrYbLusD1S
bWWGfVzZmVodUVOocIKNyG9eS4f6A4BcHjmyPAJyIFpwzjl5UwIp/MPWQlz9wXe2
RMJDYr0KAT5RAbnW6glUjrLnaE22U9ZtPWkUe5nZkr0y3rkveDn5xG8vVqNYQqPz
3XBXFGETgogCUnV8y/U0y8UkcLKQBRS3i8d3RikVMfnAAuQoAkUV/5AtEI9ePc4+
RGIwYBAlQ5eDw/ZsLXgGNS886LKZsuZUiRZG01m4HzXE6RQ0+96BBfBWD0ZGwq00
pVmgmnbkUXmMPYX1sWFwy2GLNDTiIeSErnJxPwspbXbGOOCJdzj6w6lB+2tr7sho
qurFIvqLNikdbL+5vXFm58pUI3ICsBh600KfNP7KlJ8XvasfBgruD6WPvPa6L+H8
JTtuynRhX65nY/d8OxMq8bQifqcWkhSYFZmvhII/RrItuNAfthqvgBLehe5WCyeA
lDnoMJ3+JYk8z3UIvJ4H0JVYuAJNjIzCzhNdF2rMe3Niq8Yh9LRh5kLXL7Mw+bPH
Lo4i6Y5g6FGN7glKB4sdZMJlRh/wV4Ouro6xwVVUgZkXnZew4LtdFR7NQ54MiwuU
TdWwVfznWFJ3+FjMtG9f0anx4o0DYpResDF03fZbenILsHWsd4KbIb+wf8BHx2KY
jUpJZW7e0redJzxt8Ep7RP2w7XQqMzgn9YgXPNNf0aZVrYFhyiCGZCp5C33l2PFM
6NyE2VVGasneI1UZFQhrhD2pwXCX5yYS/SLvw4vtxf1be5j85TqS2i40xnHzmx3r
15IeHq4oKaSPhayk7g87Eh/1PtvdT+eLW2CYH5EHL6r79bWRugvsEOUn711rQR6q
gzwAWMqJJi0nUznOztwUZshBJZ2rfUWKIunQ0dD0z5JRD9g177I3v7XyiuOhYRw7
zurTS5WMOp+nyNksb6eA+PtIsidtp0NsIF+4hF6RvLIvMfBeuC39Isp0YX86q3qO
lJtReiKFUy05BqgkVdmaiGGbvSXNaUac/ISflYRo/z5vxS3grQEstZzfkEHAOSee
rpuVjYtJTr04828gMbhtAFaKhJyX8ozSfV9BTBveS0hHi/8V1BKCCA+NnPuAHsRP
c/S2mWqaxnpaqUcTmp03d2SZhZ2/a0RiT9vKcugKrdNOxasGFuApXICBMDsxyyXy
Ir066tuSppZ5uRXlZgp+3XhESzeqRS8OcyQdfmjoo/cUniF5OuQt0aJ7gPoBG8J2
gmFS4eCE+hAR4PcGAR4voS7/eYV6iLL3bpFy+wuOf+VHsp1cctWF7LTh+Jd6w3x2
VAF688MtE18PpJotDXjXR/j/uSjsEwQBHkTwMb7vwYElPU4kBWo2jlHpyiNEToGV
/jL2iUda2nwY/ZhDLbnJjoOX9cR7EGRNixg/HtUPKDbKlJLSmFgl6zUtzTLO2xeJ
Y6z1MRgDwDP6zDkXUnNsARciKsZlyQGLDxFnY19e0qfg5y7Ye43a4OkY1m6depDL
mVmuGne4RmMhOTpCgo6WIOkBx9l/3lI3v9SDyNQHK8HfnVVbkU2DTvm0KIAKsc0b
xiWxGhiqsGmu/dZBmsDuxbtkjydpHuXT6sILTK90zdiUDOsWCAjyNR5uv29eT0s/
zvZ1ml8qayPI2HbRJubL4vVFBxCqzuBqpPongaP+QC4ou7vzM6CbIR4+C6ZANH8V
WRD4ZYWnMfLg+blobeFowViE+vL1MtjG1S1oBNxmxepnk1sasOrHVs75WCkLx3RA
JxBunuogbdBLrZfuZ0cXawDHewnW4NOulUTGQ+nO9htuTgu516eEK8yYQ01m+U9f
6laMmgTifcgEsfaMQkmFRpiGOHuAecX9cZU4nQjAP881VVgtjnl0RK4bOWTgPLli
qLOP9CCo+Nr8ENz/b09SzPrWBgQo2yP/pj+0G/Cw/LoU0w/FbkJEKxquU1mpbW3N
Y3bptTu/1Es2UCYWnhZavG6jT5TGfiFYfVSPw+k6t4/+RB3lzcPyrTlWqiRfv01c
eTPvw9cZlcJ6+rALiGL6NVjoucVxJ0xJSeoi1/LAWfo0fdN/4HHLdpW8z0P7CBB4
trNTV34IU6EEQRO2tFlCJ+Vf0YsCz4PL7PfHe2UBwpBpzhXLjfnRmC6qNhZpSjOu
SnqKBfE51yCYOlLDJAfINrysERbPKESgRjT5Uma+IdNoflH/maJG0HG1293AYlKB
waXEKrcUAbLCYkd8egFM/EeaT1J5ctQ2UG7ZbD4W8TZcPs91SM1JsX5L9DZvCba6
G3ENCokeLuJYlqh3oTtb9vCqZjKWZk5o7tuBUTN11uADPsYj++b2eVE9RbQ2fRFP
ZqC3QkC1iC/hsriU64Xt0Lj35dtSp97ze+gXCvrofwMKlH2YZd2DNlMRYBoNo7SX
g0K/dyE2LO3Ht+v6M6AyeV1j8hKTS4PAdzLduZNx/Ezc/hZm1oLI7+l70FuaFEH2
ANDwQdfE4Ek43gKyKnQtt8EtD8L5gmTVCcnNhoAdgcOOiyPHl2IRCB18ARsHvRcy
Ux44dUl+HFfNNMBoKWxQf4x/olMFhg86DHEI0F3b0+0OC4sPK85SGvZxO1PXPPVO
yvsyODaynO4nK+JMcLdB2Th/RVeUmAoasbaHO9/9GLixnpNpM9FmG5FdzyPE2WER
hX4rEnj8sjSRCu6zVbVnm5NGbms/4UUJoHKRpcaIziTH+0VuZ+Mvr7nCUYjqqa43
fq57M7r1h74861aL2I1WgVfM9AZ8mF04+xAj0EUl3SUGdsxJ+Qd5/YNzbJ65jGUS
Qjp0kJWHPZ1WrX/+4jwb2hFTuw3S1SmKGFHP/sT+iVrIWsuVQzC7mipOAeMtcVs2
6kVxu8+K6R0gujp3QZoJNKo6mP0XpLE2lBN/By2pYVtoSraZPgVQCmRTg6FnNfAP
ncFj4GDYWaI3jbfKW/Kmqw+rpGC1ZO42IHmLBz3v28gnos4aL3wn+wPdhKPYPG/E
pVMaHZTDE3yK0ZPDEb82HJMk67WtOvrFApKiN4ivFi8MMEur6w/7YPYmyI23bG2D
h+tb7pPQCaqmJSSGAzSafTmH0qF4a4xddenUFuBXUtyBVfUDYElFZ4CFLiThUrG4
QBV13EpyzcsDOWDbmUuFoNPng7k6xHoOLkQzIfrFN1yN3NUjtITQPwvXOXf9IHL1
sIIQwCTTROODEM7jM/5Lk6d84A/9L2un2i4WdM1QvE6ZxZtx44BtyQ+JieQXQ+/L
YoSyA8CVglFiuUmu8bbD4CzvYPvwYaOrEZmLwSv7iJc7xuhBCKwt1kIcqVTKHssT
h0UTtCUbgEaLybkoj2MhlQYMHc6XCgUVF7QyO/mX7Z4TPId1o1HGozo341lS1po4
aMUJRZFyVEpeWvLg9AkORXPcDPVpiptZzODHEtK6u1HvZBuXmqX1HoTemAsiNcwP
f6TUh1IzbcSvXN9PljjCNsqVdPwl+6aBczAt+DOlMHqPnWsbWLNpQkaxErQj5Hfq
SgmrD/JKluwgeTNsMHRZtbeniLJ9huGJOxw8U+3gmMZwMEyRkk45MocObbyljoUI
4UAtzF4+UqpZQf3HH1fALXZ5qNOTA6dtcKeeC8aY0O8yhfndjSQbjxn7g722ndUm
HxagtHVZ6jfMd4oOy9jiuJluqT4NN7EKNOvpcjtrzwfZhRXFYAIOe0I5BK4pVDbh
c841TJkXA/pE2CIy8Tbsn3sM/Nkjg0GELp2tBRelmoXOE+RmrprTfpmL10toll4x
uJ430JdVQEW4m5R/sYjx8Q4VCNJfwLXu7DTkp7c384EHYYCbl219H5s0tmHSg/i+
tcsc8l+U3WClniivCnNuWGdQhr/C3uYPqDrzVKdt9tZNi0t9Pb0bHRM6LRAOhyb+
qIBgV3IgP2Sn/w2KkB907Ye9sQQkxgv4/+F6wU5a/Ocfd+AhbGHrhs0SJbGoSNCb
t23TdfjKrzjR9mMsBAd8HhyLjaisNKdb5H6w7iAAbf9xESOBUObtUS0EbKyRl7hz
Yebyax0I00myEzBimKeXYmosV9VQVkej9LnG4kCC/bsAIk8Gu6O32rERX9t5j90W
EhL7KGV5Z4GdvUfhq3tnvXoZ/3uuf5CAhtnLofIUdtDf3uxanVbt5b9oZBYbX3JT
YmnuMXBJWeqwlen3BN3mttNiJP79DmbbgHEEiwwgc7SFEaByIM6XTpY8P/KuG7Y4
kig+Lba5rwJpsC7Mz4hdoDPi0M+LVQEh0koG1SmyIhHrfBnYPBagJAwu2KwpbQuf
p04661mVWbJ/Yh718xgQA/6EamYFKa0cJnpOXNlBKN/sBW4Ax7uoTbULjZv1J3aG
XJ1+JgfUAEr4cWth0a5CDYbrT8AfZMAEmMNGatPpIUMullDl6GeCpC/xUKqHl3TK
UTVgd8fkNdy3J5AG+wdXaDR8WobPhpw/hEgvReE9NQa4fc9ee1ZrZhzfEzuraGof
T5Uzh+J6rWqlGjgPBXwfbWGdRigC5LPsR9f8xB74tdb5Gs862ylJbNZ14aV5PZNm
KM6ecLUeicOf0y4FGDBfl9ic1cFE1T1HXgVrZpwwqRNgFMmJ63fxvTQyJ+tusXKw
LJcsbB9VjFMEoevYnOFF7I3s+ViNdCufbubOum6a0FUieCSE1+/DTbLE7VUclu9H
p2hrFCu/WlLjJBOq1goOoEIFadEQup9Bg02mR/B0b3bmIDsZJoxhL7/wrRZhjCr+
FUz6Lbn2tRZXUeMjXOK4+MowSf/NXuX2/z5dmRoESn0TJHxJdYVzJ2i19uTy2Ce8
lw3h3B9T6lKiwGYvt6o6wP7/Wsip4QwnWHVpCK2GGHNbZvJ0e3UIONALStJm95Ic
Zl5M/JGHiit3N6bETSHCMUzAdHMxjaxkJm2/1pQSIEznJvwnMpI4ovril7C/u9kX
xKfKSaCau7g/74am5Ot0lrpUrkiSLVN7V0w9rf3pQmqyubACBGBpkaNfee1PGFKu
ZSQdNeCA4q6lk/MaQNgwZp0A2Yqr9YljG6nw6bpUNQZQzWteAJKGi6PCQ0LW93c5
sKpYWNhgVOCr3QFYCQPo+fmBE6qcIEMySWJnzVoE0v0T+6v02+rdVaQ+IfqNZU1n
0z/T1kvEwDnTdRf7MZe8fBlUncvHzjg1cm6QB9pKCLUjbSepng1e3ZEeEArsC8Ov
p9R4LzWGTPo8zmqfbXW+TXlXonwW+6DJDS6T8jZFey4ooG+5A++Am0k+SqivIjtS
7JD2b4VppJ68iVmApLlDPKdlomvZ4bbNaGAFV6Vce3chTQwB5ed8nVBqGfG4Tt/2
fJqPtq/W/HhuTBqnj+cjkD42OpbWhpxxt7dC8BQuUH56iV8RuYJfMnp3ywQUZc7x
nupP8CWU0r4OckY5nkNY/kMAi8soTEvGCG/YEjr/cSHTt0/+uPY1FOx31SDR0HDX
dKMpjoEPFTgTmj7FsbB4xISR9TOTBGWSbH8N2vjtAKJkfrdsXAogU4VXRFB54Pmd
MwSHBPYpWB/SIs91st9ioM2smBjxLhGhHR2NYKJzsIOCuGlfjdrLVg5DhWr2wEq9
uUUw/7I3oSYSUBzKwPfx2dUR85CysG+k3TlGHfKXqFL/Nm1pQNc7v+wRHwJK3E3h
aRVs840YAzpam8VcoFlJpULh3+x7VbtYRj+ZkrrwIx9xsoXGz2DbZdASWNDPQ+Em
C0wLUFXJZzvyJbu+/tSkAaszNJwSxxiW3QAeVuN4GqPPQsul+0icFLK7ZcC6HgXn
eFVdCqujhU7HdXfjokW4Hs/oVlUWGsv+kh0o5bGMQzI7zUfI0PjvLrJrprWUXnb1
ltL3G8ccEHWRkUVPMTfEadKtIOjCFBVzBTc0tUMwVn1R6V49Ihq93KV7XH8Y6Cvu
cFslv/CjwMMfyrxKgZtl9y3ftbuDQRslg9QLFeUnsuvYGzu96O6/HSaEEyDyvD6X
1w+SJRpetGJpc2ZtLgYpmOBMIumfR2SP+tQx6xFuXI2cuNvdRavU/XNUn+W56NAf
CgWSkNc64TUEUeAdvTD+WiWORba+k3gAkyrFIczPjFMIj8NyZdtF9YxWQv9ajyn9
p3z3CzE3e12dR3IhWUkIgg0vh2CoaU2rK38Ab9RQGLf7f7RcxLPsEczMrlZXAhQP
o5H6fSboA1XqUAxczhLNrfV7P7NJ4tJNMPmelEOs9ew3fNrUT8TpkuPVRRAZ/LFY
vmXhz2Mw+dCzkMYjdVCEcOrutuC7UJ7M5KrwISvvJQ6uVKQlZbcyXNf9+vEjsZ2V
e0Y8R0Wm6WDLYEVF3sHHeEcPTR1eC237eTI+OqE6Q8z0Hp4n6rOZPabXzlgYg9TP
vW0jPMns80PgfkVMHBIUPjh7LNXcXUN7fUHdoZUssQmFe+IkrjStgaAHJwVCHBPb
PtexMd0LdlAkdCLtLXqWU5elCHaofosmxuPcmwyqNguFjTejYL40f1tXgR9TFMBV
v0crmC9dWqGWm3haA9Kw7TqcPor5okd1nYKubqeX/jOTsC2HiqU3ZNFw2SgKaXfG
KwCEzznW1B0OsxVy30zRakttIvwvBWGapYNMcln22fvKSUQhsTkjj8OqC9+7U9jt
1JfPhJAzV6faHe0prszgwAg6mG8QlVQCZAtkQdhissRs4WYazhYsgHHtnX8dTVmx
VULSNof03PoXPls2QKr+a/ClSCDL/mjpJohSmQVDDWah2Fdyca6H4SmgOKxUNVJ1
fwk+n9aUQ7/d3rFiZLTnY39FKhuRBpNbEwNi31vdWO+80YzSJZpq0c1zcT3PbEaY
SQuQw0OXVd+l0bnargIcw3XwMh1t23iUmABFbttUlTPnrtuUJJH6jxiUA4+8IrOT
axtcBQ92s+ekpnzkNtPpyCks0acu2Wvher+L4txbWSAA7UTCcqKJRjSarRwBvRV9
KRkLu3HpQBiAcZCluRg/AbJZ/2dsT/tZK+Ke7tnDSevtf8OGqru3igKt1GxjXtEt
W4soR6Y5/uY2bRKMpzzuggyVs/Z7MqsZr9Foml8go3Y9pps4uyxA+rceDBA2JXxL
oS5JmARGXHBA091dKTV0CeIRqR9TwF8sUI77IDgaC6ZyMy+8715gR2dCWgfADakH
YUsToBXgJ4Gd6AbPKDki5zczce7NC/PGOvQr22OyigDxUSCoAbXMnuoVjtdY9OX3
HYkA0JmSA14zGHOLHqhnrg/+f0YL0B80O2EBIq0/pRQ1SzFzi4JtjkHzbAeEpY0G
U/NqhQQd0qLCgyjpL9lijl5I49bGtruJ3ytW5nl5VHBCX0swxpPGAT6LYGAQF+Ki
ICPhrZI7/uVUy7fPPxEWG/NSk9N8phibpI7KuV8giFZ2gF6n5SlG4hHGh8zcM4v+
5bTIgrNPDM5OvDk3xj4hGGsXZa0kQEaTmclp9bf88nzLoMSU/GIjxVc61jGOC2sA
p4O+Q2L/Vz4QxOBYkL1UGFzB19vdLzN2txPKI3aUnkQHN0GcecQGeOfoMaziPz4Y
btnr1NtmF4r+TheNaljd+1EFIvF2C4Iyj/WyXbgURv502VMMUKz/I3SxAPaA06Yd
TZSri1xngb+ae2Y6xtAwMz87zwdOafwAL3GBEnxhzTIJ/5XFgreLbJ3W843Ngygy
MAPkJS1x5rjz86NuGYHOieQd0QH+aNnRY55lgftzh5nIEvJEnUUe0aI/8CpR5Gja
glHfgUVRSsTjDHG4lxvUbE3I/1PCx7/G212gHcNBSLsaXaQUJ7uwHQwOjyXDuFIi
SFU5bAGXPKcJclUU9QS4tMcay90hFovne/UOMOb1Imljfi0GWdGz4wf+m7YkFOiB
uGYfnbWNhmy6GEw9491O1934lT2OOkXLtvrehfnSyS2GIVOAzEerR4PTI20Mc9gw
yO+8rSBxjRgjABpmaMpDRL43OUYDH5jLghSCxqa7ksRrkSh/TlEPbE48XOl61oST
zxrW+8FnhmHxuyXnQ6mvuKp3CR4PEszv2k77XYRksUcBl7uiiTY03agYXfnafPyE
nZQ0X8AR8jpR4G4Fr8V6Iq8vjnvtT7dWISxTq2+Mq/1BM9zWloQNrn/DRXypGoCp
pNgysR98CO7gEvPy4jdABIQHmruPEf21ae9bCkxraFYii9LJVWJajqh7fQ3W0wC4
q0io76DKozmiNid1zHQo1JjUbMkCmJHrfG2Qsv78zbvUVJ1SZcP4Elq4KbP+WMZl
Q31l0jzUtDhjYE688JHD6KX0No6cQ4uMDeMAEycuLhPVFKcGnQ6mx8814pYkirqV
3KOrcI7gHcKvqRCkwj5svV3uyf72ijNG7eX1IcfzdCJsCyB+DXXSSzgQY5bPAFjt
KjSzeHJizGnsGE/h55b0dMksrox4Kej83tS2aaPCHoqhKARSuf79I5xodJe6bSgs
iqX9CF23ZCbpPNdvJ2X2qxuWA9M2vrZ4s2oegslwwxrFvfYq5kgpX5WdoV9oI0Up
0si7EWy/gsLz3z2frmLJoLbxbbofELlCm8yGg9ryzq3QzQQYKiNuMrqV79mrjqw/
OwU22OEiaCDSOiIM1S29u+Xq1OLonXhbow58oSZ2U6joL3uNuC4nRh5sjrtKTphA
P/vYlwFlm6DgrY4zD26+5gkiHOvVJ7zNnFLKH0DSJn1N5NHYfN23dLtrBJyU8Zb+
dAVzBaY+B43Ae3OZR8u70o9rOEYRoifAu5IAi5Fj+HsaUL1IKEmbRpuxZKcEjA6O
TkLN13SOAaPLXuvi+ZrbAaNqjKFmQHhKHSiJdC7giTduWu6E3kXLD68hppRMUD37
VRogN4EYwQ2OQ/5xzcGnpqx6H4gAfPQz7UFDu9n5JEElFHPQuN3Snse11HWRcxvk
wBbrvUUzLaClFbFntLO59uoeDM2RDK+sVafrMoJnzP2O67/QwIJYMhOsE5/XBEZ4
Cfvso4ZU16rCm1xK51VVTjgpotS0CeImyKWApyU4vkE2NXGyjIiyqo26MfK2ZR1J
NsAqwmWswRQBXIT5pQH5A5RuPIQmR8+WVy2M2xthkoPYwiC2IDH+BVhj+zBnDm2I
fCWrvIfWvLVXuVBtRbj7Bw8yErJ/BSubfa3D5a/lGgmtpTPvpAvNBGXygutz5DB7
LTkqvS06S2Jl69qAhoA6wCHfsY+Mr5CuCR/MTsySO7WCtahTdEzo6d+uy5s6eZGu
Euv1gOWpFMsu2LnRMH+WoOPf0LtxTu2GZhU+EPfjM4BqdO2y8tw5pRb+3yQT59av
vfUE8pNaRSeE4pv842/9NFFCw9uHbog0YTGzHRXtuZFtk/Ecsr6DqB6mGSavItyL
byGnjZ+aZdptzyveadKxYTGIuz4p/wNFV5bf9aHr8ZAs8JQAWoMVPjE687mxLrDZ
NQiiSpg7psf8NcyyYiUUf0WLA/Wcp4xx+SVagVtYh9p5B8irRjUQb4dyTGouQQL0
CBo9lgvTg59KDOaAxU/WGmv05ydwJ49spmT31ainxWlhPfb3tvD5QL0zI14Wzp20
jS5NN9xc7Io5ezmr7QhdH7IbH7zQZtzYZq6piLgmD1FJOHlKshTnhWTtAGWTNZJk
0U2xlTKrZedJOHxwKc7OhCGqErEkUnuhp7IV1FZ65Ss2TljAJfwD4wS4uHeD0U2i
EOQ5ve2EEL6O2DAlTR+NZ+QAe1qnZGvfaHWpy/11DCk5Odfk94spSCWAWuOiBk3R
w13KqYfMRtqqttq/wFKA1olUT7txXJE7rpt7f+ABGqp8zpPX0CzWgzk8EWmF4/zn
jQe7yYkaDcOeiewow7J3Cz4FtmcZAmCP9WC8Sx9ScYZgrRxaxIq/lasbDu/uUEWt
EruYGcldWfPenJIGUn7J7bwSMpsIB6CJSP+m7S+uB4bXvO5gjdmCGM2Q3rqLcfJD
HiTXVMdmHYAAPEHTU+QEpMtMP/xqQic9O9HodR4871ljwY6QU7p2cm08CyA9AQYv
6thVmLMYgg3xlDWdzQULax5x11pWUjPEHLCtn60E6SquEB/bBek23ULWrHPJOKSR
EZUocb4yAYcFQYPhjUoCYmI6q7HMaENinV7xsEhWJeRMP5mI2BJTyz8qF56jkvYS
zWZ4uF0l/jPUMpP3vCndxTVtHUh/ZUmYMi/Syqdr0pazwqhiwVODeU08v2cndEmK
/XxRPN9LX/dAqwuOwJ4Q9LOWfYcmvmw935ft3XQF+5sVcqB56j8NJ3CvwmKthb3p
fXnWHlbe+Ao6Yuui8MHrEQDolyerE6CF7Q9UJuVOq0TOJYD1zLBaWG8tYmTUpbaH
7Fp/g/1286+BMMp8G3eQnwSChplk+CwsO3VKrUkngvaJv4jhgWHJTj/F7om/qSoR
Y0R0mogxAr6hikxLXyYKR5gQOLUd+baTH7nZJ2/7tB6ZVphM/O7DC7SOzMMnPkbj
QHdZbOuoqhr2osAWw1FVjkk/Xg+YZ7c6iTzV413SN5eOc69FK88Brgq6fnCP3juQ
A0wNbeW2vAn5Y8U8DwuTudH4xUi8TVT2bukHLu8PiK4u2viJj0osb1DQsVYGogFo
uuPQgow7ZlrnnEytn9pkhgP0myvU32C0v+AvGy+4GtSYKQc9lJVRdKmFwJFxnn6L
MehtgzQauZfqf7zeuppwHhK+e6QxvMpN3CZGoMosFduCw2U0AAub66NyVTP9EbaY
PzfC07OWzeOSltUc++VhEuXYW+Gvh5suI/Tf8PndeMMSQQZNc8LOcM+0cgtBDKJX
mQF4ADFNrYyMnMcSSxX7nn6o0jQHEER2r0AbhYcOxZboVLx1OEbQ32Bm4BotvPGv
uc5RvbaZJGvSZRvovY36NJgRUpeZgkTiyhREtwv1nmOnVF9nvJGXDFJJr21zk7lu
zmsVYwOSHL2VybI/Fz5kZcB0gcULcwgkDCXRyXVy1NVQW4Ucy7xOUu+VXKQLdz2a
Kh5NKWho6xdSr59Jqn9NPE65jLcNTpPlL2bl2tr9ec1q21L36BvTEbh7abSAJ+Qq
jWrmC7SSC5tak9/pCepAGa1w7b4uvUbyajeA1pY4woqVc9pgaTX3an6m8eGEQbM7
rory/AuqjIgN3I7y3aXyQ2Y1TdlVtmZYeeqUGRmEjkVkRBH0uNW+WvHW3ZD0msun
NCZ1s39rWhyiT1cKZX0h1Vtls+bzSexhYfhaMterQB3y7Niygp/jWzO5wiPVxo+S
/wcG7jt5NIcCO0vLNzCW8x9wxyIlokMbutAPb39av+EaLqEltsL1tIsSkGWtX8Pw
DGLUFMb7DkV8ZZBHRPhi+10dk9twQEcvVdY6VfpjQCAWhB0Mt5DJt2/7LDP+mlHs
fd+8LJrlGvb0S/aAD84K1zqT92PWnjqM+PZAVv1LRoHCeMMdG1jVQiXAnVpyz6Yw
/sfk863FPccU78J15cKfiFxNlAAbRENsC5zTFYYv/XmWZYWIkxn5tunQld7fOMtX
k4cBLEjgVmKX0NobG/H8hN/3I7xaS42xuWVGYkdWeEmnJSbIMERKPzx3Vk/cZecs
1rs7lS0BkIJ9XLduAUaxAnnWx+U6JDhS5juKwNSP5Gri60gRtARe/zzeNMVxVgp2
31/G3LSvuEiTIyLUxNrEBipyiEN2XU9rNi236vuwodyrD8YMmnAyglNqiUzdl2n5
821KSVkGN1TEU0HHkPl4/rPwymGG8T1XXmkrg/vsD0lkXM2EVYdbyFndWTWRBIHK
5DC7IlO8Mc1gA4swibbvKGcEiz/gVGGnXTIvDFxZEMYOBota8Flaa8cZ6VzWLTNF
O+qgklpVCMBck69Pyet06aHV2jPh7EPFZMYeS8ZtOl2ZdbfshvGWYoHq/zKWLyp7
V58RhHQecZx4Zc5PBa81URI6UPEsWGNUTlT/b533w987J8yWm4qRltc+xs+70VzT
Gi99whOz+P6c9KQL5dXvkIAmkidv/M5t7osT/NCm6+GiptYUDR12+3GUJikO06+Z
qfDRNmKMIW7AMVkXbue/FfQvFCbbct1X9uwAFBppIeZmJZrjPD5N7nwYLNaKBX1l
yeSxJubikBW1qwfjyLf+/3OZMoL2kmG7Rp12XZ9e7HaKeKMAA+770MiEY01QHZlN
Wa+2VS2to8MQQ07s0SjHyUu6EQAwHVZCpfRmZutyH/CP2WGmggVpYwaZWLyOtLzS
jQPi4dUb9E1Z4yIhML4ZkCYnyYHtasD3hbGsj0EWckjqcN2wa2aF4UhXVGDeB+Ds
Xpx9WOvYiXo4SRHTQCkZrDogccT79P4nY/7Y/dM6CKdewdBubUNUIBxCrWMl3j6y
dhC3cFEN5/dTJql4S+ouS4JWM1iHAj7gJiqBYZaVNZrpS31Ep2CC69kzk+KYqzIP
sAfJ0UWKhyJfcHuGvAeuqSySnt33mRmuO9UCHyoIJ8tyJPUre0k4dBK1UDuZz+pU
/CTAnCBWwCNHtQK3YSV0od5FO0cwBnQ1hM2nav48/BMgkwaL5mInu0aQfPsz6OtF
pkJdTnrdu29V6IYdLLlBDgV0HA99AgdCUelShHz+RniXkrAXzWfhbKY6JkXk8h4F
EkaKuVMmAnDzCEHnKDPKwNVbZ9sHDGstBOAmlYOpxqwIgVC57QKamPKMQomuqDCj
67Ebne7ZesKmI+rE5myTIM6wJ9vPoI7wOcupQ1Xvq2S2+R0oLjZLGUIj2HOaJVjX
nrClXB61KUOqM7GGUrfJol+Bnhm/U9IcZhVh7/Cg5hgfDp3aiu7HPJrk1XQPnvXN
40Wnw+zR0wxecFgSW1+CSpBoLofF43/jfbFkYQkzDotuIu2+L+p4yzflClYXv4Hp
spesI1maB8Y7q67cPOoIgDd9bwHX3gZzTwnYJuTdGlLVdM4TIRw+qHhICmuE7Tz6
FoRWITBtPtoPW1MzEq4Ba35h2wk1zlEKYD+KGQ2H420r7N0ASNF65INkhfmo7Ax5
oXwkf7ffLo32qyiOJ61TVFjcGJfX59Y0hOg0RuhRV7tjE8ULu6aNnluB/SLYgK3L
mYDiwdPgUvoziMQObVZrHyPAs5S1sPlYfe8+fig3CAbPvlH8xsAkuLDQ0+0KZ71R
a3qL63GNV6hOrJVKbcB8NnhbSNfMOl5n7eTWfUFoogzMSZvUBxrQmZJS0wN249/y
I8Sy+kcUHhrbjGUJFEhZ1J0uKPSCDUeHgB4YdxbZ0a6CfjSoOdgjiu9F4QsAJ5IH
DScvmJTukJ3UbAZOC18gPT2WabhSISJ9mcEkHaOkSTqmehcTg/6ejwApz+iaMBZX
YsWEhyXWQ/+ANqqUXv2zHJyVpi8ZZzCGiuiJFikkTRjrL4I9+/X+qZaNyj8L6Tan
tvfiqjctI7ivgQK3IvYH5VnjylcJ7b0WKKzDFSaRjrZGd2BJPWGSbmk4xG4H3WDH
5Q18LgDM3yzH4rSaS96SHaouCaIk9A1OTG+t6b8gm1KgUy/sS9e3Tc6/mhGIArcK
oAcdnr7zrCFN5Zx9EMbUBf4hrjuwv4wK7JQNUJaRw8A+xfBF1dqoiYBeod7Dg5jZ
rUVkpYOpSNrmrXHRZ15NQW+1OSb7xNqR9cdQc+R9wnpe/nsJSatEFh0I2YVmmkBN
bjVGW7pHqNgnAZc3oz+YKchYR082TFhyizXqJ7edETS23Yz564hv1GidIuXzHgLG
UUTi7AZtDBlAJqKLQKPnGppUmnMoX9/iAZY8+1zhCOAszKzHF2QEFK3gNonENaUD
/AOSMO0chkVYK3TInF3y0/yhzCTNhsIo8p8HoDJEv2RGQCKAZfx69rIZxqNrM4Zq
YwRo6U7pbvDFH+2k5jEAN0kWDioCWTHhYNNt6yi3JhJ4I636Ljgf+riB0Ouif7QT
BmNhOKcWmCy0fiKX69S80zsXD7DP01nI0LL1AZ/ddn2frrEUkrJOYdV8W2LGvlXe
a2zKaApI0XB2gMWmPaIibG5hILhrKDGzzpo2VTwBYpGEZJ2saDUYwBFAvKoXTURN
V1k+cZ61J4Ehu6c0haVjFLgyHhUCc82k1zQQj3tiam0OdgstQAmhJrkcvFFvZ8wq
XkYwKHuMoY26e7P4yv/SjnQv0G4dhNqSXSRH2q6gnBWF+XmdqKDcRCTRkyl/kCmJ
U2PYHJ21bChOURE6d/qCdt1xP/CoOTd+n8w/f6qfN69dlkDC+EShNeIWQwHVR/FQ
VHzzyIYQmY/QLMY1RjgGXsDDlPbAKGoWh5PfS3LPLmZwPORIfvoxCBr+m4fmg+Rk
3dS1Ak12bwRtSgAV1FRaoVKSa2aouK9GGWovHGHGT8+Qo8pkqUORObz55BRZoxIK
w5GEBGZSrEbch8RoDq6ErJBLTnY2hmlcXOi4hnDjD2ub5GdCYhMv2KYckkRvXWgR
tsfB6WbqWvBrTE8bXQDjXtWj+IvOHe4HiE7uZ5l5xQOsZL4zJPPraJZ6dtkCBKGa
WiID18HS9+zCvaCD0ln98xezO0tT1dIQ8IhHE1HOi7gsQh9SoL0oeeTYJ20+IGc9
/n3UdUYs9IQ4wurPWbtWWtarxVTKDGpvVyMV3ogcXlTp6ueaBB7GGVrHYYZ7/OIU
ZdBDLxz0TGwbiYzrOPU+PtRcUQpj46jYqZP5qdfvywQf1Rk3CCysXqhI14SubFxq
KcDQHXZ04uT1sKjk9PS9yAj6CC1wLJr983LsEK2U2tHttc3PmleGJGEXLxXyI70Z
XDwz6TyQ9xEcFcwV8qzZJ1eiG19lJ7yMlkS5S5ql5JBxhQ4OKm5AZeeq8srs9QHK
w0gqw1nOZhoxAO2sNL5RdwL2baj3PCAQU3yx86zN2GAVC/A1+TQXy597SEyjCk72
jCnTR1PCj/eWcflLbTXcjTsfbfKXzpf63DuJEEx7qemJ2tg/m4f7d89PYGpPlst3
3tGCfcy+npC7fNkLSyidRdHYZa+PXrt5ctRf7TB3YDDu+hl70z5x2kpVoPgwveiD
H34Z4ZCUgPWys/67hyzZBBYbqWkJ3K26GY/X5WxhGj5+QB55A9IrjiVixGVDyhXP
Dk2lLVV0dzZoDFUe99lbU+KHN8rnW7UN9BEbRv7PUMNhU81KkCmL/LdHUlyBAFL9
diZnH8wxw5ah2p8z89oRNWQVeCCcphRYyTvNiy0eFR9DdG+hi4hir/dd4L5StLgi
vJKAJ7/6UqZetwcv+WNhlNv2/Hcb4YbA/nO6lNvp9SIGwioa69iBFHrulnwmaB5z
7dl1SoHO8VmCLVdF7DxlMjZyNYuXhcgcJni+JB39QlP0iMi0xtrfx/fWSUtBUc1i
S5ui4u2fuHWGSVBDGqLXuczy5cffQWHf+tmhZg960Pu1NTcelW/GqOrrk//vfFAo
27aFNf2ePE49LV033KykefbE8RdfJIvnmNJkX7l2z1w/Preo1ihu8NE42THDIZWb
qCec7GCWVjnMjw3YudcioG9yQ21X5Yumz964oSJ46kICqWLJuwB2+sYhoBviXNOw
vhd5VKOKhM1yVlhhW0yZjHik/Al6oWwklgBvEBG0WYoBGj7rI9m4Z8FOH2XNzRfe
d2B5SnTr+Hr1mBXPOcc1g6JwgrfkKTysl/Z+dfGKYpKiDkscT27B2YaHa+Y0+vAc
ZqAhLiFPJ8lGbiBfd9rHqUXy7dI+2bETnUdOVdInIJIkiGetW0o4BfQZ6GlpQX2g
j3gj0wSWlUMLcomyRccBfGEdqkUuMPhF/gC4ZopjT5Z4HIevn6aWzA6lMB1RTwIz
jyQKQ4bIK2pDLA34M9tJeRddCjB9D/Vk3jLPo0CcRUqGCKqXHrRNYRoXXxU1Qcc4
v9tmlNWrEIlwWUS0wKBtbKvhvHFRKiKb1RPsGVoiDpwBQal7MkpsQptzccYeniMI
3mJYChYAVH6143WJ3b9zYnRzz8E0RLQ3yg/3KiS9LsH3x+ze5gRdUC45KK0OuXWt
C1pYEVADX31T8aLByIIfoAAPQ82iKTCYH66+7Y79Ht5qlOKAfdjcd1oH4Xs6bgr5
F3Ymce6BljOMrnlP5jKzXOkmwr9K6a48fV4anqN5Ldiz0BQgfSWm8AeaHzPfEhuf
ZD1ZXZonpUxh2gl4ccfgUH/ySRCH/Xp3xTYUNvVP3oadZciJHDrDAnrR3vFO4HLO
A3VbDm8bkDPEN8CYVNuARg72Oc9nAc0Ma7ia9cM3TJZTrDeL8BU0s0tTTQPODosf
ZnWkOzpNHoyf+/MK2vSxm0XWlgOLfZcOAoU6LDVVc+84jrZtOihsubAW96ZnRhwi
kWH9okDtC7YybmMyebtItm1jeCAn2SJ7ajEEBrw7C5nJ2zcv8FiYH8qX/hMTNOw4
ysyd8MegBnPOTKU5tr842qrp6db40DMc257k6hajTAteCW7PUufYx83AxbczYMsy
AEMXBwggQQRnWlHi7SF9YhDZ/As49YiD5lE7B7TADUrL1tT1ubXtRhtmOXP8OYSF
z/ypPAiw+Jr2p5L2m1OYSM4jNS9ipE+JERCw4KwHjDw6333fS5oLaaoRLAiY9fY+
R2mDvRboA1iJbXIzFJEC26lZlTFAUR9IhdY5kXysWruOoeHIaC4CkbF2gRafzztX
b6qDOZ2rUoMH68ru1ovmXcmG+XY+9uhhtnPxwRRaZijbSykjg6ggOmSjr/ay20Bl
c99822fHCPM9+/AvmsEmkM1TJYMYu9hgOLQnDBpxXS8cNDeMBdMOqKtblgd0ZkEz
S37d0SDkAHOwja2ZTAQ8I2QKtsQz08pCfxbRcjvYE8DOBh33IZuCmt6RpHz2Tx+c
0LKXtlCZnpNn6HC98TMg9Eyh2MXO9+ucgPxCM+BAEqfX96C8v2EXwhXNXprfF6YR
uIVtaxtt+0WaDkexMQkkMoS9R2lSjiU17nLQX2zRoXHlmP6KSiOEPPETmcFBVNHR
0Ynl//3/kvtK2g8rYqc/VD45TpBD25LK8XdskWC1ttPdX7n8PDcYbSOoTf+Il1T7
nRcrhqnvb572Mzrdli8JXJTrq3bs7P2ZDtcn/oTbvYQKseonCgWix0cCMOjQNdE2
gEyn8ALFxie4egBtVdqQ06JAFB86vsJln5G+sKQo0+JIIZ2vH31P2NqbL/z7//n8
+VeNLJXM1AddapZH8qlL1lyR9e+ZSfJUTrQ3Bt1UmMtzORC9uWCMBwdR9OJ3KX9E
pv/tnrdNjRThyyjF8rhWZ9jk0Rk4dv/rs2k/CfCX33KM6vv5J83Sydii1ihgQJcW
twlWhIxzmlhE/VmciA1bCoideGwAH5YlgHC/Z6tZM99ItSj3zsAo+N8igBB51Y/O
e3/FxBn++7Q1rQdogqlsCdmogwOSb6SSY3dbod3/W2tTQrNuCcM7Qjbq+pk6nPtO
2wqC9x2ZcMNOOEMhJo+HbdzheDUyROtzDBMvs65ogKt+TSyumCAMXTQcHuV3vYbU
3ShL28hFPM9PlfWCLlZPqH/cNHW5OH8y5B5O178wrQ7KbRiuIHCQZjJlnUuPdawA
mPqaPR665yADj4jKvAY2wOMLH3QqIg9z/ZNDm91+w0W7M9gxy8vbH7LdMNKvjewI
hbgr8gG8PC01AAiAmycLtRuze+JzHQ2uHz3V5AvHWLFok5yBD4lZHoRCetn3Fn4t
83n+7FI2+82iTOG9ccU1L1/WnlkpPQqp2NDyuOYmbNS4c3oaQHOqD3bGafJifuUZ
RIV6YaC0bYHfE7jFxn0+YwYzx5qD1h/3A4Xu7oHQkgR9nF30YlJc265q3AfBo5iC
qxJh6/8QooX3iFa234NXftDO7/GmEGZwDY4gJCH+zKA5NDZ/9V95PQpWszWef6ar
kRi5UQNrFBsuzif8CeBkBMUO/DXCTGmKGHXdDfrxrFO/Qx3kUGQ69BrmLgvSwT9m
G4uCttKbGXVINmiJCgA1wTio5SczykNqUee2JQbcmO42HxavrXX70VzRrwIpVH1C
vf8s3ibOpOZ0xhluPLDo3hoGs6+CA4DujaO1hXhmI1qJ/W8UPBNst92AaZ//rC6C
SJQibL2m87ifIKFQgf0XNdYJ+CbJdCIfeotLEyelCbiBJLqYvXByN3hse6WuGM52
Dr3nK46afSMk6jeIgg2fmvnJoIwxBVNeA/hrIyMyKU3Lz+Ei6IHJl5qkabRxKcaB
w1mdSNi9x95H+Sy+UMAoxrU4SFuIxeXVwWeYNKETWgBalnu/y1g1s+6EBbihGrkN
5rgTv0DoHMI2Xhty6WLyM/WXidNSGCr3o1tIEc7LDP810/lia3Qns+P9W58xZcjP
SPNPQ0VeU2M9GqssWxeUqLfmho35+5qjlnkBN8IzEcOSsytzheBLMWJwgCptC7RP
jqPP363EJEc8q9iVa7EvlWM0zwb82a8eLRocU+tPRmD6fcJzucaqSwGLdlRwzk/p
RejfIvuaC/daC2SRu0b+1dIjpW08T32Fcu+4jao2QWGjjsjr1TY6ghXfwavWkTYq
i3MCCDx3TOuYqkq3WqCQl4Z/N0tcfeUggGBcSj77anvHPeRGuzyNi07gCP7nzJR7
Hwn64mIMRm3uF1ZEKQFzmZb90IPI8l/uGL4qL+wv/qTpkN6GeIswWckxjKhMS4yl
694cnFL0VXc7/1seMFXLziBJ8Q6hQXjM0yKroTd2DAzjNulX4MOZC1mU95XPrpyg
5Wsfh9ns/NKY75/rsMZS36Gy01B7oLX2ZkKYTG4oU48OoV4E1/ItZAIxkj8fkqQJ
35dxL10tpJrFiIVLfXkMqZRw1JV3meK9ePWgBRkO8wo5yTt8gpb5K2oPjVFY4Mra
o1hH25aCksIuwCtYe5RwPjY8DZMFAU1j+i3bCvex+aibC8tWS0phKLDr4UZtVyav
1GoB44g9gO25o5RxAAI/XmsAKRqwSybQY1RW2balw9xoUfh2q0GGXfxABOe1ojB4
wenGolRnU9OMrDedsjZ+00mZ3gUmhcyUVJCGwhphvNf+ag5MExbcvvh6nwzSmrV7
DuK2mttAV6dGE5wVRK5DdxUM4S5FHKtCgyA0SEaquOuC+Lhygxwd2qNsg1LsQRhA
0W7m2kgKP6k8hQ6MlGkGsVH7zS3oqBCP2saxgI681R9U201r3CxCruE76pHCd7gp
0/bjkWKvMGQM2w6x+PLDH6gF0tJo18Jz80nZgBjKkmvw+kXZgaf80PFTAZljPYXl
6nw3EA7e5slF/N5jrF47d3C5gx/UhHMHCT9HiwzJ8LPs75Gh6ja4x5FmhHabKtBw
qA9kW+2NTXmJyAUuiDsNGMDDjpX6I0T/w5NHISzKsV2V4DJzaNaNtcWv94396N5M
gt8Xpb4F5bpZd07vzsl9QMUnB7B3go+z/EqCp29TRH574y8r11X5k0RUDeGV5FCW
F5BFY5umQjEyQ+8R0mj54IBUnAhr8TSOzNSmGHaidCgnN2KvXpVdIWcwBOdcvNuz
3t6aE24a3SkxD1W6Ql+SZIb7WI4N5QOImFBSW3dZ983u9dS7Sy0DHsVDaAVJKrc/
NsmI5rvO9ue4bmOJvUKzUydXx91G7lpiU+v6bA9yGHohdDxIkbfAljhhUe2AOpDJ
cLp+jZFWCNZeAPmLak71JbEuuFNNtJZlzolGNNfjS70fDIcY4mVHNVUo+U0s0105
wlYCO7P8P1Tb/1aOzx+AH51x+yEKSQx00MQGn9ZY+AQX0wqKOwUSjzg3H3ENUdXX
Y5CB3h467TtBGgj4P1WBLL2nLrF4P/hd/RLdDehUmswy13LcWDr+o+EyyQqsWdgL
4YKAWWxc5S6IWaLSAfueEBQKyr9F3SlaEt4aH16K5rbhr2z8LfJfYJ+V06B/+2ZG
Ya0vlj8Hx3rwPVfPS3OYbwxhduMRPK1lBGXrEBUBwiNjF6eBLziN6eyr0pas+s2D
7vR/IHV6csFpHO7B13JTNLXG2nvjblma2LMn7rXh/iUPLhZyS5+RgESK1zXTdqYh
JCTWkbrNlrYGtJG+cucMK4HSvZpCgZNtUPvRk6k1IdP4MYaqcFObIPHl8MIZlEWM
CAVsubGl5bnlTvV+1fpQ9GZAl2gK1k9uG68Gbjdyo3+TISzycyvaW1943TEH+eaH
0mJRoQ4Kp7x5KEA9IYvEe7RzknrbeJ+tpHrO11rupzLlUBiRD+6a7Qkj8OFqZp9C
I4q4OBueZnsHw7VE2q1Y55qFgnzhcTWuy7l5jfIY4TyFm3LTiMg9eS9qpSh6vrx4
ku2L7ATAkPiGWTTDcEd+C6Tmg8ZYi+LTs+ilVloOvgBjg99phY3+D4sv5QrINGbu
LkmzBU53YPCuGyukzDGePnRZiCIUrAuFlagYdP7DfSHrezdIegbBhCHZje1f09op
dUXFab3B1GsRvf5YQmB6dYKOI8qpuJtiLk/dSx6uik1t5WtDMJWL707D7x3htrfe
NHFTj/Nz/iIRoieMCfToYGBDqqHHGRH1htf3uXTRvRpuPEGljRNvf6IzXtPGMoMG
q8o+Dp1rdIjzRuDYPc9xPORFlSM+NRu3+sVoxLrETxRWFePQFLPfR38gtpfXHXHp
qjNUMqcWYhBxkPp7ZXVzAnuIF2jgDE3nEuPY4xuPkgLjRX/+7GXnkEVLlxIDx2IB
qH8QuOV9ll8UZQTOxVHDHFncvaPzw1hx/wisWYLQNzMEwXpEemzODKTOIPEcWDM2
OtTM9HC9IM/Jmc8S8us48AqY5WUSjqPQad2kdWB3bfSLSwMxnugrIcAFGrZliMxS
b8tnkvpWeeM5Ks5hxqjI+hoLBJ9wcMOSP32dMJ54kH7NQ/7MpVz8olgSAwofhXBA
/KWe1gsCJBpZM7yyMvKhr8IOVlCGsOL57ew3AVe2ATIXHQTgtv3yQKi8EvAw+daJ
QD6QxMO9xxASbh2pvzOSJi92fF9/5NBe6lUzNXyaMKjJFroh3f4GnPN1ZtyVyMzn
E+W9xZ7EqDr+H6/4PNG3ZdIu9U1eV41LYNHpctVVjYHMlZNBR7dKzGGAbMxFGt5s
vuzv0mZQvizWTLkbtgT5JTaUqfZl5Njh3JCpFL93vpI9zSW59NsuJ20wkoU65sPC
RA3QXNVsZ96vAI9K48ffSR6GdQ2/eB4mixC4sOrVmPZUWT6M6l3kVO01w9Z29NwH
rIgqFc4IjcvH0idTT7i92sHGYIVbW67oJgqYBIbUi0MKkArwU9xMQ7GbDAJYwVfn
nMh9kzIw19w4g0BJ2aPY7Mb7pjGHlepHLZgGXx9N8ZhvuDzv5+9cXLcmhxXiWh5h
kA2yOpblogw/eTTGZY/K7031Wwg3UUeBe35C/KfQJ8XsglNX1CjVzUxLlOg5y42F
IC6u5o+QxSyYYNSWTy1v/5P1hEtVi43n7OMq1sCaNvDr7ftHwVnvMTEPdKoqjPxO
l/opESRcErIHQkqjrjMAXgDetlhQB55cCbnylVWar49z5KJmu5GO3RwrNuGZsX+M
GeFbpWG0aNvhaeQk4+/SoPxYVy7L62r1fRlcSKGMRxtWDmCBlwJxrK+Ev5fA2NBC
+vBDloDjZJ/eSoRpCrDcb2M823ON81iAgUFCRqtFEK93kPLH9o8PeyWYXLWDQYwM
ckXA8SBh5iQ1IPY/FrwSELEyxSHih8uIkCzPbW9x8/0sKlJG7Yj6Rj/cj0+IkRLb
VyJARkL/WLH8KdCwUS9Eu7AGQwe1iszG2gRMNzku8l4I1B6fmz+xB/ZeT4lgTjRJ
okafw6gvBz9FKpdKD6q5zYrg+3/W+cA3e3MVhaibcYsrJPMzgzXpDljC6M303cTn
03pecmlfWc8Pq4EH+kKGJ8TdR3g4aPhTMaiNbnfQUYjmT12EU7ktTkkxbs0ISAzu
HmMEDNa+3DRZO5159r2PbjECiod0grBWalyWjwAayEtxJPvKGDWQuPkogy2QH3On
A8CcgIIO6jcTqhNKzMTFCZfJwxwMgyZyjrCKWvVRiCLzywS2Bjm+y0dnBkHef5dF
Fv+pGgNV6xdnY0mvRb6JggW13bw3pwEHYAKLEtZEFQxWNzP7TP8x9Fb5dvZ4sVCt
zSeZkTxN8ByVQHmxd5LnQSRy0ApYMxv4qROcIWug/ul2naP1F3swCs9XprjctVYu
+CvfR9pMtnooFwA2M5i5MN/yUIpXKfa+MJwFgmHti1U8XEL4GJcmyakXuTjQppkA
EIuz1saUO30ivmuKKFK2ysxF7yH718jio920GD3wtiFJCMuHdduCg5j8u5cMULL3
ZbpTCuDQ0hdIKtPL/DTCeqbdHh5gbQr9M7tA5ZcVLZcxneyilPHBDsmHRr6qLsSu
EatuGH+Hr9wyBhWQyIXEzoDUjBmUjeQwOWmYX0KuE0ECuUxFhWbuvXA0gxNqfZYx
luvIbDpeNxvG6gphdV4EJrXUSjYirjWTGP6++Iq1h0nS2bkdMJwhDSiaM7huUvtu
vRDCbG6hKSz3KgtIkL7BIWo1SV2RrcmK/h838ODKbEoezKYY3YIAqjwVT3r0ZEiz
rUf9G8CRy5HAD4mypU/iNHNmyOFoc039WUvpDsN6OUgYKLTofqpBmhWdjyvRLMOe
HtCOgPEWq4B8HHQVTcnsVqkEGo8PAAkh64yKOVqUtCbak5JLAWBAhlRY68EKuYiQ
84dsCXUTPv3xpdDmcKEtWKrIXRKZKqRRH2BuP3uLad0FKhHK/cj8YyRuyMaFaKFN
UkJD5Jp8Woe8mISgYBhoEFLqHOlMN+4QTENoX9Uevp5cyYSaWtmteVY6/ciPV0gf
/OemPjHbwLNJTS4P5mcHFrE6s/BtCDCTElM05shPTH7r5tb9Q8iSR9aspHfYMma0
VQK00FL5+F3zWr9S2hz6B+DV8J6ShMnWsyPLjh9cZyipMORQdQwMJMNT4qL53bXC
vR5IL4aGwGywmId9278x30XwA0q+WQIcQ/GYUd7PqS9O1EqR31OEmaimC5Qt1Q8F
7TxSvNdgMn1RKYhrl7Dof+VzofnqRRG+C1ZgD/LyTbgfGS7473EXj+gayjXOLzVy
jmKW/eiepNeoqtInVO/q9q4xowNtKB4Ax6tEj71rdW47xAU5gucGmlCf4yA96wD1
//pyxSExQ+SLplXWXPeJ81NQKbeJrbnjA5w97WKkA1P2l912HZp7akd9pyfvz1Yl
pO+480n9d2pjAudYwG5o4fqC+g0ErTl1S+ITzqEyFdAOn/GfWRMWSOmwetstgKtQ
Q+Fy/qESFcuDGpUKZDK7hlHum8QA3tZ0rEeyeMBJrI53aL65ZEVz1XWi5Zn2lUlX
I+ZlaxLUz6Q+5r/wxIJ4qdNWk2x7wwSyDYpodFXd00cls8Iz79ThJHF+RyqjQmfM
tjPdmfveoPEoBnanppkekhLwKCw6HLwvHoEJ4MMcp1TVr96at5/+yotmItoAMY0G
PxLNqYBHfaS1S8dy81bwWy6bJ/UcXTOHnhqvbXoLqR4e5Mbiu+Se82HrY7sjdxWN
eTGV6UmsWcBLG+A4t5VQD4gSO9+icreQVfsVW+CKJMmtnRcatdko2wehRXFt06CO
j6C1DtlQGbPh4ibbpJIRvqYhsGdPlqJohYQTB6CnR//0zsJyaJqJrMmX4R8sxySX
6pP7QShmt3ufhMa7njaVtYa1K1nZb8LmJLhe3eynMjcLtGH8RcPcZlGek1wrpX5r
qdb+7m4LgKVKp4PeHRsCk8PrNLwkiUoLtaIEbdM/GXJfMEpbsPNsIy/YONqCpWkC
vME8NpgzRgw3v6Iac621TCKPE1Uug6ZRMfQFwZgBQrahV1AQXOXJBao49GH4QCK3
LhgVXNNuVOdDAlY2FqKLzFjAahqPrRWAlpo/4Tka3ZUiYbIhaPalQd1Mcgn8PKHG
ntRz8rs9QnvNQ+9sA+soTnAtaoXa1tghhtIk4dXIf3PMd3Pma9ostRFEnLRUszr9
AICzQtibnRMrGgCiIYCiChhbz1k1zppQqk9TbuCfOPm38gLkBPIE02lK2F/dskNY
6H9kgdiynYlJTWx5OZ1TSKbJnbwt8YKW4DjDqpZMlMNzT6BDNNVVvJFfG2oidOa6
N7jsz5NaHkCHYd6n/cLnsZo5UF82ZIPfItO38+qs7QBncHblftFm9eaoreeuA4h+
/PVg5SafUaSeiVXS6YPt3rk+0LbiH/q0yAo7K+xNqvJ+06gaq7PxbQ/Nrmf+Mvw1
ECeanXZHy4DsmYc/0ASDIkBlHrylBWp+AmIRBeBNCMlR10yjXJLygNqCdYTV5+jP
M/5zNlCJs62g3UY4EMVjpyQYik8e7GdV6PH1QSZH7G0CuDCfhYy18rfSq/3Ya48O
xaRZNRXjfiq7ItCSUoo7JcKHjwdPiMb6TWKr+tP6+A4MHfpLqFcXUM8mShb1lxzY
pIRZb0EMKm7O7+QnVNvcgo/fD+4yjzppk1/ri2rW/iL9RGYUWrpe8yjckknJQ40i
x7st2lyUJaRcbJ+RkUXwQiN311WAbj36NnK6aLpX/EmE++PQWlLEorWY4+V/C/q4
AzLwyCLbLhJCdIDyRFI8DXBnfcy5C+oBZWR9u9Dg9T1v/s4iLAO4EOMmC+2laa5E
yzWER3PSDOD9QNsZtGWExZrAtdak8aMYGnMCqBvHZNCbPb4JDwpoLmiD/a76aymd
tn5cvZfGLfdi9tZPyUrLwaIFlorSBGUkPiF3fmUU+Gzbc6xUgxIEg5DNUCHGY9FR
g2zbvk4wHOA7HQou7wQSZabLOikQ9+r1sVXgPOuEhsSjqrIbRve4hHs9klNbyq7l
qbj75ono1DZDUgK88dDZTaUmMyojQsjTybVfaWRaUG2HFmUCBXgK0JxxqL2dcsvG
BLlvm9nXQ3Wy8zYUNIfxS10f0hb8p2peTDYypeOhynPXdtHozDkByg97jlaqePeZ
javPRvfwSOUoVlza5+YG75FmCufZedSyfP6dLSzQsRZcVEcEflbIzAa+mxtw1RC7
d0hbcmBqzZOXxy2+jHtML0p5d0wdlYaOp14PNUaOULgHrYbe8nvSKjIoNqC96Hsa
MfoccgwHD3Yt0cFaD87dU4FPc8DQrILV14gA3l62BxC0/nG8jCuEZF8KzKKROq5C
bfOPchSU8zmrE27DeffvZpKQL44BdUMKK/76yU2OASav068JK1S3hHUXHrzxbpdm
9JPdcTxw++a+fZPwmXaUF7DVDxEI3/+3XKYm3kjPj1iOU+KzQfyl5PrdxJXg3nlK
HVswTTJu1tEAAahncx0OIuKcVAmIdiV6SIHuumqOrDNo1Kvwv0BJGz2gsdDkgfhL
d16Y+KiAfVJrrx7vr86pJ3vQleLjFCvCEb1oJ63gTw0mzrYKPl38mH2lomJpsnMs
2zX62Q4oP94H6163zRHeNiVrO6vdaufpBei9hT7sVpuVZzGRfeWTF8ZhnJcSUCAM
cFA1h6KZoqfQnBWFFDVjjGDEX6eUdjrP4iRQR6Sy1CfNB3yuJEy6uapu7RqF/ict
5a/dZTvwS38EW5idvlm2EmvXbG5LOIqEn8CRV4i6D+Pvy/gQV+sdCve1oyFwhgF4
2IVMubnSPCLeX14NN3Qs/FaeuAaR0Tu6yJ8rdF1ZJIazQSmgqki5nq8eJPm/3ast
LDuhbPFptSFs3LxVYBRM/O2HgmyC5WZQiiOvGgD8ZAeT1OB6od3ushZJyGONxqml
pFnHxWXVEkp6ht/Q708kDyQWjp1rDYghUgE31FkWlHwSVKCtaLMr4zpZRt+x0HN4
anedta1T9l2FJRnwPjRL2Lf3Dba7YAexM6F/XU+LywObsQr8DWtukoRIx+EPMtCU
1mgjTFI7+xEJcAoslSxn2kAYdrYuYKnN55gCjZbhTBRwYIKsbE8O70mJZ61BQt2O
BYjGSbJv7jF69jXnl1f7Ve23o0mU24ULoKDMR6/+lc4qa1jCwap62KRqbPhfxzIL
Z6nzmrm5DPcZ54U6Lu1jKP8qIurF+HheTvPCsjaRgmrt3Fqi1fjXMB22eiEv3YSq
mVirVkmBkTCU4rABV1m87hHsqbovCoyZvM768yvov89FLCJtaLYmvz1ARDSGbt5C
WIZTnV9WjaRma3Xid8qAob6qZ/Ely/PypCL5cFBVYSb4bqIwfJr0PPslhbHMAgGz
BPLcMS2RhyNdF7/J5mlXKecW0eC0j1LwwtAJ6LfcnA6Ezr5MXWruby3eYMPNd4Jv
z9u+wk0ZdLXDn6rGtD0Z4wfyKjhn++8eQZySa5sk1/+RfJqVJBJxCWuOhHPWxSik
fsyEOYztRG9VmmsSoWiDYYltO43WsfJE+SZWezEFMDePTJ7kGIRwg7h+MQJ+ieJx
F5qc7gnsEEjNtT2acrTzmvSyBgpOKEWSxn1eBRdf3Rvih26UTpmaYiR7qErseRl+
k7Apq1ofqbpyz7nksVDJgRHFKY2bYJBt6wCxYhkg2ZSmDMnUsMRtRyZs0QW4OQs8
pxtMXu9+qwA7a1Ffw80pkJvvBh/ujT+wO/hEsTSzDSHTocQMRo0vziFDW+czjxBv
P30Rt/faXJjBFEpjtrPe06XORwVJNQgUrI93oTH1Ice1ckvHwWBIY+ZzGS6VPtHS
QwJ3MPf72fB6Itk3LN2ExepizU8Ukk5JEgwCxPnMIhowvavF4p8kr0AMl/OPyFk/
TrRydly29rpSUzBXHghUHmSMcDBsJ7x/cxl2Bed/fnet0WCRnukOxXZiVQ2khg0f
cFsKWEYMO3zfRIBEqJ5TNJCxXtb1nUWoZRgaJnka0NpoDQEOvMqZut2Ak5BizVPE
j5pXexYfnyNH5hMSgzlwja/5vb+aD0gd1k+nrRwosEzq4FAM3hDQzI3W38e0jA5O
JxgoGbJJuYfZltLcHEb+mjw4jHtHCkPtFr5dcqkTKD6vAQwj1viVUzy4eTsAnDD2
sfjTRN4ZTjqZBcEbBMluzXrKo5RuY1DGMc291dQdjcxRSMn0YOinTelg2Lq2jsTI
H/O7AxHpmBfs59DV69rzIh+qb+aMAGwhdpYjNxqKyV438wlJe5Tj9SZ2kbnzTRqx
S/xrRxf74HglNZtcDhnb3eGiZ1wACk6uxOCMUd/bbeDMFCVzG/vI+VQjvSigCYQZ
vXEcy4JUsx8DLGW3uBeEw0leVR4175E38bUnb+P4S7+c2Se0lk9JMh5ankbSReuJ
kaRQ3350Lq6tvESftCwRL8V6qPj1BuoE8BM2ySmim6BfVdfQLBI5m5J6pcGVtR5y
O5lWrFnO7Lw586dkh4CxGICiNpJJNqOUHnvwxu0U/FsDg6uliFEYfjiLz5RdEWFx
EBnrHYedEwThanugDexVymXL5gMeNrHKC6qNxTFIMfDv+aK1Ke2xOn5VaBVYRtUw
Opgd/bcPu889Js9mlsM/xi8OOa95XyTUWF/zQ645oNpO9fJHWJcLVqg/fp93V++M
bqVzIl7eSEdhseYRQddBNNhSyG0cQSsDITYLH6ghrZmnMZ+PfBqUQUmcljWcL+5m
+UScJN9F+F5/dOuIorSBdBH6bB8a29TtgoR3X5YaVZmDEF+3HLSGDrs947NlX683
OHTfXrEuwHv3dsAZWTieQLUmkG54Ld6/nWZ3IG3GmQrYaoZSvJ9EEcnwBMG4+QN1
YhEgrU9StV9nR6WQUctIfzyn5yB+sMKbfi39p2QHe3pFl5itRHegVZxd1DoGlE28
xxpxYyy03/6x3E4gBay34LcKqIHPwsVfjt2czSTNxccxX8qMMGVKZdvAqkcuYfZc
rHK26l5CM7xszDZkc5ejFkg/OCI7qdvWJsbZLDR97i02A/+FzrHiHiwiE8eDe5PT
U2e7SGGW8J+H8AKi9jBV7lFgqHZku8t5LxvXW3TvlRf6xYWTaL7rzXgRYAqyznAf
FRiyWVfvr56EX/8If8lpKyi0y3fTGRqyFwCe6Lc5Cp+zAFVueBi5utbbFSraiieq
mQABmTJr5AqGvteIxgIgKbr2IBab8cj54EtuSfPBohPA4alxc62l6IM/KbmEsmnl
YV9zGmw7A8YzJ3NJgaH+TKojDKgKNDqy45jmYbsL22bNKjghxYb1voE/C5p+8fZT
mjQa9vuJPfNwi0mH3oFBRZXWiBZXlUA8YZRup2rZC6gcrHGDH8Z6K8LWp9GpBLW9
X1qwiT7rxbkXIpydjIvcAoSOpVCVf/g+OuDrpkyPiiO0WQ6yEWtuq87ZOH2HnYAX
72WdsAwR+VPB1/2tC2trH79JRIukHxwuqpe5oHRU0/tuO/gO0yt3zlEUuWoNvvYy
1wY+z9lY2oci2+sKeJy7dMzAeWa1IY/2k/FrvP8t6w1X9TmPxWstpnzdkJUn9lrB
lD2dGygk/HNR7IsHMMPjK1lo17c28DI4E36w/tR3PXYjVAofw3/dkaQqpjHKCzdg
yPnwSztJ9bS401mYo8PExtH4UDbtzHuYFoQrk1zPeymm9wd3IwgqLRtzo8gCtPzI
09bxKoMtz2P2K9dxeJLkxeZatwtChgVAoegoDC5mSv6kF6ZK4NYP0vq7loPb/Fxg
wkzj5mBza4AUaDAoNsn3QLsp5Yl3h1aVD6W1s8W1M+VjQC85I21p2gQTe0uRCEd9
rVRjjJ5PuH+ueGxUkqdh4i2cnXY++etwiXPqQ5zu1KHNBCngKsYWGwB9xVyIHpij
zu6Zu47i/qR1W+1nRv+C2RZaJiFwbF49stnpp3uzH2pt3P5C2EQORJqtQ0S4v12q
++MZNltbV0Vp7y0TYRoRxb278mcqLO0cX1YEkpVe3b4F6RkSf/CPnmt2DKYTSyW+
SuY9OMEa5UhPwwDxwOXvnFreVz14j+RU9SY66IyBEbBXc/4pylRGjYQIQC7E5HiD
ttMiRQjPbtXmx+oQhBxpGaxT/RmZLhSPgmEMRgKhLEucWEq1s70O2KtZuNrtqjAB
7R3ocBSsVlMBKRkfnvXPJwZ1OmevCyYmobpRAC3CORP10uQ9fGSax3yvJMBtknkp
DAiIQenACXIpECVcBLzQHIKEpUDqgCpsQHY7DB5muOobgGgD0za+wxOr6FSE2vq8
3cwXWpmDmSqeVpgwtrEbQQdmCjZglafUXIMvYOfTXPh8tOEIXxRfON7RiWukAZD6
aIvKRqxzd2eI1ZQ1vPcs4kQ/Fhrh7VkrEKZCIDl9IdN/6eWrx9ZQknQaqBWu+VUC
L4n5iiv8EgpanRMwS1qN3J68nLOgv/eYlEc8QKi38ouWaOti0uYzN8BkSIM4WfO6
Qz+1Grr65nazRW2hcGBS4dM57+UiFUQlj510NjV7yssI4EN03cKYVovjoJknXij8
Vejc+qhZ461eBMrmy8O9o9IW5wqYpOHPp8Xwi6JBO4o08q9Uq0SLROkAWBn849lY
lBfWS9fRvL+ajyRkkvUoHWSVbKHwVQr5KFRFaCHmlK3O1b5FueQ2zt8J5oKYaq8i
RenyUOrI+QK2bpoB46Hd0ff72NSWQsJ6JxSsorBE7Unp4Y4mdap9ZwPe3GjRMoLS
88l5ImDSkujw7oSsC/Ir/dM1sotTAPP2QcLXZfDtDcShS45eEFBvSz+m8gBPgGnm
5GHSLVEwUoRQ6tRXXn/+Ud9aQ3QhedCBuF5rXt90kgoij/WxnkrFz8iGL5NNngMU
c5a5ZoqL9Y6GGG55VDy1Szub6u/tiJ9TnA4AXCvMCwC8bMpmwMDgFddIatlgxTdA
mtJtGl0nPoytZ0HLP/l9EFRHdJZIA6hgLfTYtHtCO0po/TPZQV+uFPvQPKmkFHuQ
LCHHUNCy9FwqsQEpzSLMvnwtghWSLJRiw/V4ha/ZjkZ1VY7gK/rpPN3AiwZXAeSn
x/0enIcuok1e9nJ0fyiAoGETWX/r9ombH66XTKhS9owQv2CCZFHKRJa130a/MSA9
CxHUXrT7Jj31qKP+A6C6q4x9QzSPzclx+MN0GTWLBzsYvoB3HHLe6EqejY+Gr4PO
CsQHedzaICpgbc05a7ZIXpW49ltezdC9u92e4+R11Yusj0xTL7UKgn5p/fpjAl9s
Z69zkBbKPpq8IGqYyk77rRxlEElfgVhMEatf8KAWkD+etA6uubH4PZzQzp/nRLOT
sA5fQe0u1DYuFrTpU1moIRYJkOttX+BgfQU1wX9kOv8jQRWS8htIJE9hHFtc8J04
odEi24OTMUwKydK4N24hHMUhFAFMFkA2tkWHNk1L9OkdEchAwjH+DpGUUHQGQnfJ
6noH+18Ygqn2x2V2rL+FyqVsWRrTEenRj9L7H5zEIewCxVJhYFd7cx0sisYxX09x
AeXa9hJUSZ102UyeRZhznNcQp8GpvAtKAQqgX4t9qeLNOv97bgtC+Mbfc5aZyniE
1Slu2Q4kSmR1Nmaa8NS1h0svzynnVbFfa0wovrV+NcVfuUcKte2JlRmiOpWrrpBS
0FKBOotKESQ9mFCsve13N0IPgjVeUxil5fKVgT4+oIa7YnSsIrcQ75KUaVxj+hSq
nYT5MpZVNjpry8yTyBDZtemU4xwouRhUStq0y5duU44BLCGiwvIyB8P3lOmhhrUw
Oa/nZcA0iSWwOmvLk32gR0RFEPY3kJOXOCKb3+9/gLqpZkXYgnJQuPiOPF2GEmFo
7C9iru2xZswyW4/W7/cnC4ogv2HR0d/iHIEhlkV1phvy5akq9zJIfFBd0pjT+z0z
TBlzKBRBnY0ninCf/tgop/v+JTIOScDxposAcdBrmur2sZK6qV6LPYSdQtNeQdf1
BhiAKCLRrR0AQI7HS/qap2PA4zi7qfBPj23esjbY4YCE0Jj5aujrhHhhwsbyw2yu
4nFAtQIhFlHvsZ62UBq0hvZG9yPblcxmKXgwi9i2P6A7Z2e7kFEpCKOkO8Cdv271
PxPlx/Rhiq/ULfaIoQFPyf6mPu5+0ILu3nQRf3bE7Rlblak0R80LRCZev4xiJNum
DsMwXWUlI60WsB7QMsemzQrE12XkySu8DGZSYa8h9cMzwxeaZ2nIWI4LAUexUzbn
g6A8FHb0WlvTJnsUvQH1ymD1ZWOF4+cE4HlC6GDpSZoKCNkbr5anz6Azo5qHj6vW
WenonE/Ryp/YICf/eD4HB6OFB+FH/fnLgBilTFAYOWXu3dbieqGDBNVGXnruXqHG
2U8SNzDGi7Hp3nq23JIMOYqNIxPtyulvMi2gupmsa8HvzSGR3vcJn1DqdG+0Jd0u
P2zhpiFjf2wbzKRoE0vxwZLda8Hdc42MQSw2q9+fYk5LYmwG/V9PyxwnDd5LcAzD
EUz4UefE4K/auyd55WFwIyH5/6zER/PDJH+JLB+0+vup9CzU6H4MeeT8gWkjuy0X
58iCdjCGdSKn/o743/PgqsHBwmxr4/n7bXsSdvnmMuEswNHC8OLSU6wqsJYNNPiL
N9/TWcgEMvdAQGLQ11+I4oGIM6LVLpk0Ta0GO/IChruTBxvgomlhSSvrHDi9R1Xq
zSzCcmjbrDs1SwxH0JdnKrJBClVb9Wq+6u/o6fww8bTRv1mldSAO/08iPcFuCBI3
8SyMSb+TwwW7cJA6SZ1IWBDgfxdsdnUnbH6RMXBGPi3DmAlOFe7/oqBZRPIfa8yB
DVMEiHpbPcvNjZxbDGb06amyQBppD39MtTI5eSww+yDgjdj0+7VVCWJnpKsXe3Om
zXnF+vD5zofMKvASV53lxKDubrGBR6w4lvxWtrLi4O2Ri+GD1NvDKRpsnTzL8qEY
Vz223VR3MoHgar2svRZG33uk5uaiNkzAuzL+gvYOx8BRK5FnRVWptWVcRVgk5m/a
UytG4Sx/T+1H+nNTNkvCTKd+CGbdQHegDP/OVvmYmS2A68Rc9gVUruMYve96zXQc
SZY5Ne51+Z9E9/RfQjWo+exJbzVpY+aLDzJaNfkjxXpVPKRlxpLcuu/F7cXg7Dy4
irCXt8EFNz9T5oUEXh+njKjyUUyHFyrec2giEstYlVV2DsuVeCDkpXaQK3a0+L4k
Wkr7oAiCjauZ8GbGnUGd8RYQQ5d3+ihOcqnMyIm0fjpTGJBs9QdZceVGBp7cI5hX
7SWSt6DLWGTEUf1wyeXf9U2yRC0/7FUv+VQ3paPoCE+aDspo3mcW3EvxA2qKkDRn
eXIJq8uxjdDx7GkIz/527SrvUahsXwXXHUYn5uFbPdD0ou6kWxz2nhYchKsrrtwY
HMx9/QGQACrNYgrf4WVumelC/3gy5r5SRzCrS/ry6q6B7WA1EvtWiDorrTXkX+lO
pdyb6ZnfbzHgdYYXKUX/J4wy7UatlAWfm+PzhS6rDa+1c86tTGZafnXLHWtJTQwM
QTwQ0GEJp5YOxroq4D5t4U6PnsQGVkwmzO5M9RZ/soJDGyowCPb09EPn0DZm0o9k
xmTrhY2D5c7NHfWBcA58u/ZcoWBwxbbVeZr7ULWMtsenYM/zeXtrgFyl6fWRQq5y
Cz6AXCDFPVJmVJA2TWte57uuuiOK136qEKbVYNym4d2F1M7DdS+4bqvtXfLZluH7
tTPAE+SsphtXlYRS03hZy0XH0eYv0jn1/IQHdkyv/UmM/OSc5u1RATmdSOzxd68H
iw3iiyBLEtqwnUOWFgAERbFK9kdzlE60OUzlKEdvZW/CnC1I3pqbKVzXZlIrb3Cp
mLwTMUde3sgSwzdfFaoSETAdyuiNMaqihg2Ni80wFNoB/+qF1qj0F23/XP/dMBo0
XJR77DImuO1AURKkF2WZwdLwd2yUABMU+ucxR5lD824gVPadtFyXv42dh3iK5dKv
bRMqAri44OV3bwyE9kFsYBeLx5AsgwALe2vU3GLtLnN2hPaTC2q6QoPn0oHoHwxT
K0/f0KmD7ZWPiWyWsy21l61eqPTHxEhnRPBbJYumLkOrcTfjloZLMkkODxTvVTdO
yO7bnUIx6H+KKk0hG5ripxpvOrM/Q9k7JOXiXi4srL28nn0Ev7rL1VRNOuGIhebi
hWgBNkENjgnOuH+h2oajaPinoTJsrmQncP/GPxg+r7Ty2Xxzv/klheAxtLUzxnFP
i9WsO2lgkNrJ3fifdwrSHQMp0iXhouMo7jHaw+pKS7fcLv0LvP0pitqp5H95PF1H
AlkZJTYEVb9/11CePMpENMhN7sdwVuIO0UEzY52LD0DWGNob7KG6lO7HATIEoUQm
9EIdyfabQUZwUvAJNKOPZu5KkFEAnXCy+6DoSe4tXqjqADgi4anl5sBcR9XTGN8p
CeDH40kyKrKII9DsuG4nA5uIrjza12KjLcQtW1p9efcNxF9VUaZzc0zIGjlDGDb7
P+WPHbthpSqfTHAhNYS5k9vCFFsJVuI9ffjUUlju+bglEv1/99fNQIYx3iJRNTbd
2OhNydLOCuAhOdFyY/JYacd5sUc9+4Xv/k35CSW2PWPDbcxQ9Bylr8ER+7DUtnbj
NbepveqFypp4qknK1yP+doFUeeUIUdarf+rXm/7yQi59hcq2CZjfrrHrQ/gmH17C
maOQFB2C08VddQks67y2TGtbqWJUtlRjxD4TGlS6bfO7CpKHfe4DSruP25S87Xb0
zBaNCLNHUF1ePZNkCzEtw7YotuIjHVJjft+fjGMRWEwTOv3bJFbD1uhH3nqe/mH5
T9iinfFKTVXKa6wJSXtWBkCLsUnW5+Bh6it8ItlyPbmhH8f+M1dgZRHoHGdSUuza
ZB5i9ZfxPnjU4FuRuoRw1GaTFLOzoHJY4Lkffzm1lRgpan/KgKa3MkK2AhHoaRRd
euuw5MFlYUsRw9TY0tMIuTfbQ8fw5r0Pwjp7sOrsVQKMaRCZt03SJ+VddWdNZqpc
I7LW8IV9W4mHAXvAmzrrmvFvKEumacpctqDJYwvH4wl2sVHKCipaWiO6dTRk40VB
PB5D2flqB2sb6ZamMvYEc4xW9IMoe5EZDLNqDCH5zlzmXG0azLKheUiPK9fgua4W
kdrYKR4Clua1xaEtknlSFjlW1rd1+YfGi2nNKnLbsNup/KT38mYDikSJrw/giHwn
yrijUrBWSbab6MipZ55jP4gUKRlK0nedgwP+juAUP27pBOWPepCcaryhxik89C/L
SJ5e9S7zyTt5RI8trPePmriKpXlPA0S7LXkn9VAG655PVHw46cCVGJJxtKtiTkNu
MAY9dCyy75H6nz00+94LR5HZIbR3VQjHUPeHNZtE4hwzCUgzyinfb8Rt4XMwms7p
1QY2vCz04mceR1nubL0rYW0sT/HopgY+ag9d5sln/tjb9WogeuYi7/aDsOxdqekV
aHebpPb3oHgieG0sXFhJnC1AwspRDIrzLR1h5Cwlsm41IJH/oCQV3W12N7utqlD5
eHKYfXTU2DRBnQrEQQyMGUa9nPHrZeIRn5LAV5wJbXV8YOmh7smgmQ7CJDv6ychG
Sx5OlX/dIh+uoTB/qXb4at5kFZqFFF1sFmBBzYhNbcOCQtHgtTxfOfHRT6Je9rWq
LBhx/a3bogWirw1S3/EXXedqCl53xI+p4vx72ngs9er7BC2ILRJ9gvTxv5uztthn
9KNHB+E12fRI/jDKVCkpL1BsJViK/ESf+80lvoELGOoP2jtgTnWDbAB0B6qvJ3cJ
//y2VjoJxzEDfMEAL1Eqfi+Nw+waXkkG2Lb52awxxoDqB18mPMZSreFLWQg/mRSN
6fzbf3orJ7+VRC9IjqQYwZwGLdnUmAZ/sfq8ksrx3cHLixodwJ3iALcNZoY6ODRj
OKyNTb2Jm73lJKcJh8PY1iUtmSdNYj41+HLYbUAMFa1jX0NEEa6qmlFTuopFJUD1
yvKj77LJUe5uiLFR0P2F8w==
`protect end_protected