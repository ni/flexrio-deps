`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4368 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10CeaOEXBiLhDCSNU2a59EqJ8j66PzdYNtXJ0o0ns3Wl0
BBCOCEvk8ygAfN7rhrEuoNq1NaHWkieehidwQ1mbjhsTsEz7xMN8aXJLFoH0sulL
OPHSq/xR9t3uXPHGA2GzKs1PlbpWiCbWtrABM+dSvAd5RBMtH/KTuunjNp8M7MEZ
XtPVFsK+tivzixh0FHD7bXn38YbH+r5MgxxZaCYY4WQfVzwc0WFy65WWdGZ/3WTT
4z96uCMYqistzlCFybX55n/Ouqwe+pqFf2B+u/o0cNRRb1YJ0+ah30VzN9Hn/oOP
ETlDb/zdMWShSEYAa0gGKB7JjH1+0tAsZt2BRCGnywpBZXHGHxHqZMWzC6/KRHGq
VSfaOvOwphj3knwG/iYkr90E8pYEJG1XPTlx6gZEFn7rKc5wQHc2p01ABW34IgSg
riwVTjolVNk2jpuOoM605hrKRU5RmMGCxTlDzSAnZk3/ToJ6QrS4dkUgB63oqLVS
3dNqZ5ZMP5MEVTKxajSc+nkZdPhg+DZ+HLUNjKVn287jak0gGi6xGPepaCToXwu4
dcJl2gEdUEs5CdPHD6JmXQcAYsJ8P1+ZxlTg3sPvEA97Ha7PUz4UVSJrdvbDKazk
K7/LjYOL0qGx5w7cqIBYcYpE1p6DiZxVwldGIaASr6TdznM+J+yaIvRHHs5IA3Hx
FW8zapdzGQfncbBsmPqcgooccOjeOgZoSksSeSm4ZrrK7DwIsics3XyAyM5wT+3Y
XSsyn/GXdSPZTvKhIsG6sMifFBqov8r9WheHUA3a9fPP/tn38a/FGJGZgvuLhLAD
XW/pHcCrSvi3MCnDso9c/ipB/YaLJ001yHSzvrkpBYsuh6wUnv1XmZR9J5sdC2rg
sI7BKgmXmdvmf6bOMmB2sl+g1iI4ZRJkFerovPVnoQAO0d8x5wd5/sVl48Rj0lgv
gCkmAGQstBMA4+8SnsB7Xotif9FqIuK46uTAM7W/k2rzJRpAXwoiBss/AwVJt20U
gjkJ0L6U2+cNNGI3rm+sRZmuWp1HtbLOQTOEGQu1L12BQq7xeS4KbiEd/zL2ljkt
im0JQzhcO9jhry6xJRegoaS0yWT8gez7qnd91B4J4yTAi5S+5dyYU62n78X3yk9/
kg8vkEtXeX8qdKLNCB4KHkzBr7btFiZLH/Zh7Hwa0iToe1nFXcEuerGoVlyhA3D2
jyCJbvrEMGWtYF9IVUqsDZ3ggk7KXl8/zdlI25yTqUaUcKPHqpCmHDxOfqwpAg6L
fvfxzEcZq8Oc6xLZRkl1gscHWXEPINtwHaJ99jws6GuSIn9+inCFF/9N9EgoRVBm
+jyFBmAASMJv26wJPHZkp0JIKGC+LbcKRc68tXxWOhiQPBMv4LfnuPAXkvhT49Gk
vCxyCmOmbVzcqbaXnVFeJ2Ya8Tmo56CRmUGMWLEYD8U3lLWGiZdtXawRs0/DO9Yk
efMzRQRBd++ljeV5XfgCiojcHk304mIe1ShRweBImMkU68obUpqnTTfo4HbdeAZg
6k6QdeVZn56we6d2JIR0vvQEmYrXC03UoVhHzh31OxTovCR+t9FQK0P129F6e+av
4rfAGsXWgSO068QOEW0rMELJ6K2CLY5gLTnsrSEBNjjfOa0AIxiNVM9OR5SU+McJ
m2/9a+bu8OtgE05C9bNAgS8q0fjKYYRN8L8mmABRQjhWbnNYc8ufXv0b7GRDVr7e
RbneJj8TxbgSzFvTucVWSfX6SmSGpt4ouC6+0hcFPViZVLduZCxws0QyElR2/Dj0
pmPwKnI7PQVxqWtIrn6qBtGoNHYBW/UxWfqPKudiq7C82/n2aDPen5L1L3C8jJJf
nQVqE+fdxMhZ589ptB5T5+lyrXq5Pw6Zq0nTtj1snZA0AOjH1R0sSrlw5sgF+LZi
o04KhbCSwHBEYxlGqyXyB/hQ3tnFNlbD4vJHPhqOw1bOCtLVjzFCBN8JaqHPFi+C
ktht3STXw30l/KzIoskRSItOkkXyR7u5pM/yazHDLFhgjjtPBgUvjEmVBajCqB26
gwU6pG+dJZPPYF1iilbW0vWb5i180qH821psarANTIr9ClB37yT75acJSanaC8lG
FzEt0+WGESbAQflRFWdaSNpwgeJ75rvQHPEmPf/nyAvHY85J/J/zIvlFIM8ioyBm
MsRbLYqi+chgbcv1vmPG8CdbxBq6uDg4zJAO+yda2j/l4AZuXnXDXcA9YcOwLf7U
eATrIJPVA4qW9CNKym9MIFIZ5eDClxZrKm1TUaTSw5E+H2OQmWjJm5fe+lLFoCae
UMZIofNOoWT+ttdWYlsTIWN0Lyp0nOinC2Vk7Q0UKQNeoDDL9nOc8jTJwwLMwpbC
ebiRmMHeMYhYpcG89C/rfxWIW+YQ2JNK5J6wU5lzTZpX+ySpp0sogC1T7VjJikhs
mu3XX88dLLeB36tJiWrwNYp+ClV9SevxY51HYgxO9YU8jUG5nWpZ7Xu4xmhNZe+j
bZUUk90z4Nh+kycYVArCv65g+qa+g6aD7cBdyp6Ae1sQqToVpU/e+H1WtFVI3Zkn
TJ5Mw5X1qdGB4dHFYTpzy/trqyNYSXsXiqK/jNbcR76JEa/Abf/ythyPYxBY0M3I
f0P4wnUn37oJHqXEihbiqGg2GGGMMFSPmZhwtHNH+83K5oPwhOdpvBcMxSmRlVHb
E5X5a/oGxZJCFKa16MBBhHVS47QVRxCMXWG7h2865fW8Il/zFVbbsono0kuhEyPA
NsPhe/WEbCvbHImVv9t5B2usIwjesDD+SqV9ifCE20J+OM07C4BfZb8Z85dC05BJ
mJAazHHiytxCCoxbqAGbyYrnzn7qZSlYWjnxDMpfdy3x8exwltEk+4K2T0RLMFKZ
nUID41EFDyaSo4ZwW31swVcW8O/Cb+XY07jgL6JQRLK3haWnDGDH5TaefYNCOUvj
eW2TlwdH9O8GQIPyayJtoYHnJaYmxYatPeW1xUIzTm1kMvHbOpv71Sok7o22vzZS
2KrS+VU/E+WIJ794GE22l25l6NwTvDmUJF4zKzXSBM8SaNWbWpK+FqdyhWBLOvQi
9j9nKLO5rMssEa8mf9j+dYmdNgiaFd4muHb8+VmwBNLGFQhcycnViDFsJaGmiJYC
vb0X31GehrV1tYRnMLCgPy1DjKR9n3/V89fOlSGud5H42pZprUyubn8Rx+RuvkHG
wJV0D9rvYjQmJPYah3L7EzpNtbaF+e7JH595LrKGp/wehcyuiZxToPoIEvJPdwfL
5K+lB3qU02Z67zLows1OX2lEmzk15ZdTol44rqk14IumnOIwsu7vAHg17lim6/mV
EMMex7iXD8m4bW+vmGsLR/D0HpzVl4DDgiCh+2ZVxZVnG+3yo8ClDp5Bmpvtks7O
sF9lCexV1wmPsitMnuVzP2YiE0ImVrN5KPZhWSQhdPwW/aa+snIcefDfurotrpM4
4EjBdQrly0XyVL9o3ufrJA3Rt7UUHUsHH332hs9yheWgi+BubYNND0ApatvzRyxg
fh+91Q/mn1MHYK+ie3cyKLBWAvObzh5TY3E7F6LH+HmmUO2NZy6Xa3W9OF4LOE/A
CeCw/0P8zPcPW+GuGpNiv+NZm84mepzMON0h0EfeJ4/wicZQWfqK5n0e0yIDEkLz
JPRwuUXLKi5QKsB/SFWdNKm0i/ddOBJrc8D16f6CoLsBJsiYbytrni+lohLDPD83
k1FtjXzYmht6yEOGyjiJvE+uxU5gY+qsEQqUMksWVjI2bSOq68Nr4EKVwaHvlyMV
GIGfHeXQaulcw1aco/oKVySO5aFpovvqqMkftkJF1T4kK3XmmztYJSdcodP0m72n
59ci+omestamDwLmNuN4ItZmO+Gkb7ZbQOO0CB7IOkxwLX6Sf0Vrve6eiHAMLp97
mS9kj9AZgFy3ahlaXV1zD6PpC15aeXrxPbtyjV8LQLQi0lZjp6uy0BwabtjUqIeP
YVyQqKQ6vXnVuMSzWuvmJ5BPWVAx5+CvzycmGmbmlH2XOEQv8k6pQRz4449yMt0C
9kXV84LS330XXJuPp47ryAw1rIWwY3h/k8jddMDLw2x2pQY47P5U0U0mjjwSn9uE
B5QME3vB2wdrZsPNudOy010pKtBEAu3YS3zj7QajeISOqaH3JG//X+4bk38IlqdT
CDrcBfNSZ1zD10b62moyweWljKn1FY6wPPLJolW/hpG96/540bXMtZiXtiIqK+GF
II67JEHSWGKBKhI/jeyCpoTk72tyUgMGvkE7yd5U4IlzAwR0d1rjQnRqoHG18G+J
O7x1rRvSJ2nCtu0AVY/gCOHyoYcQSmY9WrYVhuHCvyzrXL96FC3falqtujwmp1Pk
0wKLkHWQpKcmuAuz/i8EM4+3BzVcJOegWQUf3dyYW6BUL5eM6B16Vt+e7sT52wci
xPlVOWfjMvo914M9vQckNo3wNbVBN2mWhRSeYOyC4uXN3rsXmtHY7T25+xFVvwjf
vAdDcwpYN4BF5Ap0eKS13/UHdu/sKuB/nvwHaS1kcWzXcUxcLBZXLMb5zcVfHdzQ
Y7FmGGs0nL0qmOz0GyTjveZJ/ZGJ3JCcEsoCtG8rQbRohxrdn9QpLhqmpF4eSH5X
X5Xe84jMvwUKvVog4EqXcrub9BSev6dts44/kkJyd0mxu9JLMI+3hHQwhkEBsvKk
sIp9WLGIwQNQeWnK4vBf793KRXo2Q/Ve8qVY8rJu/SU8gXKrIhVzE3FOtrmEtsER
xgTO9NqpNGHGsheXEzxbQehhGFd3xyZ+LNlEszuiHQPrJMtUm+nzAl7byu85uIed
mv3j7p/T6V9flLsXmeVksCSsFe3V2bCdEk3kMpXJr3kS1Nau7Fd7nQghugHKUFXQ
/2uzHrHYmpevhf/EjwCEUHznHIHtTedjYV8BeeR6CyzEMq84/8yGoLBKZcYsAVQc
SocaV95n6w81U3C6PybcBuWGgL8S0GI5knCxnKC4UOtvKaDNKvZzzqEJay32tE9E
1maq+8tb1Z1HbzWp92eX+LkCviZDdD8apWJgRvdbtYyWo1rAes7FdD47NgDh3TSc
fJKERpbDrA2AmRjduQPqxQZXEkU4DbIIUTqxdL2Z9f5Zg4EEN0l195IVWF5hYfCk
XmPrRz/ScuA/WOBT/R7ag/CP82VlTTTxf8q8SD000BTILh8FMfTDxdB8CMM2jm3r
+8YjLf+I3fj1HofdWtuLAV5SMFEtzXRhP+UlYkIS8EvTngXl0mxmbVwFOIrxW+F4
8iVBNHnklOBpRvBEqc6EbNuO9PDwoghK15ru7dP+lhCa0nDhEjyZfMZWcwwoYIEv
dHuaS7MKI7tGaMvbdaXwSVji2zsmjk7wyvqKp5vAFqQKX4JJU09FT29YcY7q+dHB
C58Wi+J1SK7H8S0x6G5UiNztT4KUeTNd9PlyFLzFy/LPIIbYosA7ox3rlnB0gJfE
VcdqF9o3OrLS23tFn2FLOIY0bgGVwdhxc1vrGiFo9rsxdljLDtakD3n2y/7KCy3h
aOE2g8biAf1fiBDIqqBXosCY7hHWa9gTLvaSs2B7s+sSsH+h7R91GBZR9nDfR5Ri
K4mHhlKQWcmzR+EwxxjQ02Zw+HYjFZKWFL+SYOlpp6sYIfVR4X2BfeVc8If42/f2
T3XXCMVX0QxNcZRb5GM7TVvbBqNSu1O2UtDUOyurxC0vCcQ4g+jfWh42Htt3k5U+
`protect end_protected