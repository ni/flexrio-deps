`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 17440 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmWdo24EC1SLhDeUV9o12ewQ
ulXp2xSZ5P2RSggIKJUy/d/PAk+ktwStKTwvmBN+fVwn2w/pNqh6PaGI6VWUMPRh
IS69mRUy4Av9hwa7ZOQSYTvaaF670RD+cDvNT7KGUL3H0A/wP7cmE7yAQu7QsuJL
gEHnkCeJMH5nH5XMOf80zMrnuDKGFehRnaVoqpEnlS/Hr63QWv2o8G9aT0ql0u5f
s/BV7O6heFxA3U73DvrStyDx5GcHjN77Wp3zpWrZroZoEkCUf4Gviq3GNLDMuBEb
Ui+dQuDSTtpy874ReWmIOO+2pcwaaKQIAFpliuyf7PxnpnHLsLl6gK6LAV6i3adr
Ph5+LXUaF2xtDp77xAqII9MomDsuM8eaxC9vAf8y9PNyGIB7qmB9L5v98JeA6IXh
E4VD0AcgYRY0RKFj8LbgulSGOKAyMC11MOsNYfayGCTVGf4+hK1YYAEs3kqFKlwQ
NhxFZv1EcttxXYP23JW2iG6oU+R0/niEXt8wcDmZUm9fi0Km4uo5ARuyg+pFmSXl
rbDCOd0mRLdEUvCQyGiCkmk3DzxGowGoJSrhP3QU0MLI/EGz3lqAhsBkaIAtcxbd
4tupV09O58YQB/bEVMviEYbjtOvx8jVvFnyv8Rk7lobz7CA+kvfDIicPs1LvGDin
OkWTlMNld6F/7x4znHZBIZyuSc3LUAdR/zx5eDHlHLSId0Rq1O8lrjmV2JCviXAa
QmSDAP3yCGQWW05FGzrJrG62fo9iO1gNMKYKc+WF7kBG5//Eu6LmsFgrnT2bnI1u
MfrZQMMza0LMzWbcx6E1d/x7stwuQk55Aq3Kn5Zm1pYzDpM3dSZnSwplrLI3EBy5
/OuGNCwrEGaazz2cdOC1lfOJ+vVyv/WsDHp0igKlxS24EDfxIjebvzVNAl5nNsYb
Kv32hD+lny8991wE4T9tCmIm6I4dbV4DPZ4akVy1mZZ6ELEmKJ+GOCpPvScHabNM
PFXHbWVVb42Ul3jxVHTgeOBGyNd0MRYM9ocxpR24BE3Z5w1VD5QowRneNfxh5dlA
0fp9Hgq+dmbR43ZcjoYBSAJvTKKcQRjK717+VRb1yRRETp0VddaMDnm8rZaW43r1
2d+KKcfkgpPuRhaBf1Rvhrn2JXjGnSpGdNphhU3xmu/Pf/QqdRTFcSF7HCgt4qS7
S6hCKaFg/r1TBAYg1axRObxX2qlj/UckHuCgam3VoNbgn43zOJATgAdEVQwlIeJI
jzB9wGhYOPnVJUcBc3Qn+Y2+QTabu+o2KsaYLehoiStBzT921N+Sv2Mv0eOqSD+X
Yxbl/wzCNjLVXMGk7cE+030V/KKSRhopYmmpM5/GQNlwtpew5Hwk9Vg0aZ5XSbQs
Oq12TIjvnePqODsWDsa4k3gbnH9SzB+k98erhcA1b4n2mtaMhmp3U0IFt4VI1hgq
xcpbq/npyMw8rgEDfeHzFW5i9+jZ0oX7fymXbdRxIODhZfDqXCkL+NcmKO0AFabn
tniFbrtk9EwcADeottoG+W99SfPm50TzBIDnfJBOotb8iTuPiltZZCpyEyXK2sUP
1GbmB0SQ//drn4rR+gkn7L9lIt8ZuzrgUM9hudkrqG6XOZCqRtCTsB2ViN/9iYXF
JoXarnd6SuTMUG14+gMWvlBbJhfRBF2KRzUlk0CCG7U8905k6F37rJY3KtZ7R2cQ
h+ZWJUV0msPQJ6Io4B1Km6iYl8GZgh3JOEIFAgKFTrEnR5huLqeyZioY7nliGOug
RF83iQVmLKq4RAqcTXqB0SJjUVD74k42nmDb8b4gwRnVhvJHP2ByVy9MdNFOl6ft
VQolzXKRy7HIRYkcUjiWIgMsfqozLqOg1/sf8WbhXuZcHCesurKl2+KHwzNrqhOK
rM76d17Yoic66utNoiSsumy8ZP35016jwrP9ddBcNaLasEzdjWubK7SB/7wROfdn
6mkZ+3pEuV46B4APo2ixWNWtwfBuKWH3t524PW3SNh5N7SkKJR2hUOhRa1/xLyND
qQBFcbuURtDWCEmEoJdBb+JjCoF5YytVjJc0LGSn+ciCVb3slMqUBVU3jbO6k0Uo
JQCuW0pSdHrJlj25vNuTGAPKocaH0IkM3eU0Ve85Rq9sc7sHcJTC1XLIEhDn+TQF
v2ktFcNCi6iYZ6aHFqDVjMYH759nESFjxOOErJuTeyYiUx4NXhC3rkhZumOBozV0
LoE2qqHwpu42dHjhesz161BsmgowVAWX9FnGyoiFn+74vyJiVJj8Xe2SjXgIOArj
PhxHuzcYmer8SnHO4BfyFD/iSHmSdxuIZYA5ZXe7EEN7dV84rsTC26JDXA2JD8fq
ybgI68fRzE+SrVuf8q4s18czSzP0YEKquLmAXtF6fjM2VbJpO1feK3TWRP9zF89y
NlMe2uFb9QLYE1FeSF7wvuyU/33TgRGglwkoMNtHG6La1vsNjvLE7gV5CNYAdTfs
YfIjlwqXKmnDV5bcM7WT6Me+llaI7PIerGilhZ8dWi+xlEvCcNTqA8RXeFeHAEhW
mqLNlHOQjGCIUgb8Tl5wgtThxYTKFH95C6w/8slmqC3kdIynQ4pCPe4iSzledguB
r/vpl0uUrV4tg12qjyfdZM++kCihTaZf6+8QpQ8g+Mv6UXU4eU5fxX/1DWwKPwsn
kRBs+AcoettTWeQ3IPfi94yxGZQUD1s7MhKqTOFynE3w78ROYGY93doNO9VBYScv
5Keg0H23npXfYyEhmsETABU85bwF7MJLbB76ULyWsbFeFtZVPPOqJfgxalgA9Y0X
g5ORoVfAJQIXL8ugPO0QJGo8Aq3Ixd6fyKTyBhbOPApP2+/2DDeQf3HzsCyjD/AB
gJR3tS8sdU30lBt5wH6gXxjU6DNrTofIQgOFlN958+5+WxDaB3ccu/BKq4aMKZFn
YcHicPAqLyA5ufpmeHAxZfedJ9HggGj/TmrOWQEf/XeP4p3AOM/A6t9b8+QH7Jah
AA8SxHtazevID7JNTW38L3OmzVbqGKfFLmPhHyvaXvj9Q3f1i930DJ9jmxk4HYUb
T+gTpe/XphaktmwSS7gDGqL1tBPESwfj0KzzouSfQHCIJyWDk8EnGpTuMHDVb6p9
TPtU6HizoqKaXq0y2XCB72ELr6QPZyxWqFur7OuH9q4P++m86mfIkteGAd8+ogkz
sgA9qeR9NlgegITQtJCmgzlHDQ9LjWgdeAkIQPEnIXhVO2dj/e+6vwIfqjKg4vYv
tobIZb2ltsYoDrMGRUi+GOoCvWKyFLCxjjXdl4bDR8eaz5b2txeimdi90g+XZxEn
5ZqHKMYTJUvdX6h/Fp7rVKF3oILdFjOonhjELCSw9ibIwANvlrXhOdFE6g2d/dB3
u5BBQzUDzv/6tln5gfmpuBo62ctzOlhDSrAIst2P8Jk02FErsaK4/RAtuttMHMh4
1pqjVuGF9eoGDKVQfNmWoeWZ+LpmnMk33a0O4SKZ614SLE8cIskwNvCWvIPBVRpY
mz9FjR1RXWaQMmfycT/mq+pAoHUMSc7YrkJnXWW6AZexrzZNdkM/Os0GeHi+MQD2
UoDCcVQLTbmibzazzmVCGYkmH+jCd79gHderiF6+StYberuZzJKs98FnLlvYIth5
hAtT03/j9R97vqIjCbcWw04DCsIXroBq8Lj5ZzpMFDcxB2hCf/vVqzS5+MVOo1Zd
fPvi7sXymjCysK2FvzkCrCfSGWOFRZHKVM3twr5ha3Q9IbELnECKAG4yibt9GbwN
UZDZbDU8Ch+mGEN4D299xScBbMeoB6SsOHUnduJmCmKFRPmKB/ey/G/SsAuOyQi1
txZ+ZeF4OURcCEZT1SlPdIP3GtUIJzECp6iimoHxjqOhSfx7+tANWDQf3eNuKTiL
E8rTD9MdcuSijXc5sh4LTmn5ThGDREYabdff0z5QKZ5ezUirhfdMQ11ApOMPUHgV
WI9i3xK1DUesq5KE3TA9yLdcnSTRnFqSfefMW40ZvbFQt4zxfRws/oBtEh1pj9w0
VLJYQjXBcnIdPD4eIgvz/SGeLtyrFhbpRA7B0jLayXpASDHIIKsl9RvWgbEf4eyJ
jw8N8WRgsPY/Os3XpZIwrUBl5VbseL2TaKdTi0VtSyA5wXlu8JHxyuXaIxqS0oh+
rDF8gCJOrCKBcFJFwgXUjlkHg9uM3r6MlhYbhC9Ub+6jvdjkD8IJ6wmVmFXiZNQC
7iupInt0sz7LC6OJQlgdtdJxmq36Qa1Q2mAZ0Q6iOF0EvWOoyXC+z6BOb7Ll7w0V
V8aNEpa7UxQWt4qUjnQDLJfm8Jy0HwkSyrhD2E9eXA+XfZKwSSIcKe5H04rF5u9z
PHdCaHZtSwxNsTiJdp05NDwal08N7oQko3qbl8uoVA8IpBJtWo1Ci7ofhbGCUVPD
SEtfgeT03kASJb7pG6hfgIVrdB5nzGqSCgR9Ti0TmpnyZI2PdcRSyrWeBXXTcNDa
2jj+AW3FYFuBuTVP/bLrxqOVMDJVMzd6fY0/cd8jconqAbmlxgg4PMq0m4NCI1sF
WXSVoC9MQchyR85rzLkGxrL/OAF2jx9ZBd/H2hmeRAUPUZDn+QnWLdlOUNfmvHP1
oYXhSNkF8PKNUz6uZ0fUl0IrfHeYZVpiXuwiGNre3j4KBqpF5G17xk12piRZBxsI
L8dtCjwmbSwHYbNoHG513ZEis+zNR5KTFXOBUReQR2PFSgNV2cItjCDwG5iSeTBu
zlPQHyb41ig5RWUU51jmVpBme+o2cE181ZZwydwz4yUPcz3kyXrMk0OkCghMvtqj
SbTmliYjQ8fW3poatkPGl+pJ4962edLvMDX0NajgUnvEUZIMUTpo5GJUUgeILV4W
0AoUUVsNNmsJCFh6dpzlrGwTKlOUcpmwdWtxWyVu23L1EMVZM8k0FMBgW4hehtwL
bbQYWyrmN0N+GB9y2jTTOw8R4FtdviwaTp89sNvdPvP4Cz9+E5AdRgdMeIXV+w9H
6y716bhQC8W2CY6ARxmK1OZE8L5JPsxJkfFvFOib1P4iaMQNnbLjyfLvBrtksP5H
HIV6GnWQTQLYFbSrNLXF/QYHELNAB7uZdLrByxpReX0vJBvxRk2WzUR/hVhul66J
ykfNdCEWFoWVHGx3TEyUtxilw9zY9GPkOnWglXerVn5Ltrz+3fyaGAfkN3Lk3ZUq
XDJeBWmY1maqJgsSUh4Hj46fEgAX/pi0jBQailgaRMLfwVkSopdfb+NEMs5zaWsm
9hbsQr0LJheWmVUy4ykI7vsmgdladS9Jk9O6hOTAeBYp9Mf0/GX+ll15P08PvD8n
XE7qz842eBPUE7HPm343wDMKGQh/3vmQ3e6i/Njp/JAapISDdfXkVVwOfFQr8BiE
cWH9l8vagwfO97BYgX++cpT/XDLEC6XT+ohy5n8SXD0NyzGHBjuYX/eLGltVEFJo
1ezZ04NXI5uuhWXiMaMFOrCeXGONnpwJEb95utR6/ZTlu8FO+IlX1dIalzKIuFt4
MRIK3rtBJzduCH8ZUWvWIVoZpDPWvBxnvmkehOHkTReSVhJ2fZ4Fy/E3/LEZ1SiO
E3MHPNYZknX79DeVYYtPdw3sHOhfU4NZPL71K9rgcwo2OFIEGqYHfnvVtug1JPNl
WgwXoHSftU5QwV/RS0XIyyUIJoryq6+I+RkbY+QdsaAAY7f9xX7Ob5pbwM7eytwG
56EbyP4b+k/FnfdSIXL05sVHzwSPZabzU3aEUWSUCPSIFWR5BIFp5Je3dHpKhgCs
JN4Qjx+ghDgDvnNi+GzYsOKVt8SudnSwPJYCft5YwDvUjqzocECMhxADQFdB6wNG
0GVTU5ZAoxAoU/J+PlqZs6wZo1AAp0dSA9Xghcw5EtV+eB09xwB3xN1kGY6O2VfB
nFHqyGZVP1aaftwU0Xhhh9J4/0cUFhDjU9Gd5KI+g1J2P2YOhEtEFcNX0jM7Mf5U
m2PYnjEP9g7RHN/UiWKT+6Ybd6vgUtjuOo3vUl5iVu3oEqN+e19KA1g2MaW8W88X
bea64tj1NWXsTl9gjNTx3vvQvn9BA9/hqKb3rJStzyI/1tyUpkDn6xELhl8vjt0J
omxiRvIrbXVq2rmCSWN4+xjuM6V0kmNgaD+1rv8CxpTrX3OW4wpaL26P1oUDWm/m
UX8yE/Ui7F1TrBcGhUrVCFFZ5Bnl6Ku5TIeY0saZSoepZ9uiwEZET7Z8ds/adB9V
MCT8UAIH7Nb5YOIC6bZym+BWMNGjaTX8j9YSNrLWxjcPqpj26M35q80i4nNYX06Q
VsgPrfKTPwVDVvMJsF27uknjZc/1rVaCzA2neTg3nuLgLjOBCF8RtzF40y2TRiiW
flHYzy3Da0k20joDO+WWMutGhGtoLsrlLul09iAy4BYsW9wdNt2Xi5Tah4MwaYxY
11S32ToGH6CbnkL7X+I/4tQuQ9yNts6phApnuxIoCwG6JNCk1vamwb/29+CytEzQ
7Lg5a6vqPUqAEna9t7CmA+mzBljnoCg9HYld6yre09qNOLj9ka/7xYShVJbW9VOl
XsIVS9B/V9dbgayS5reRMKI3ULgTWo3u/+NVGoQ9U3pIuPfgcx0Nonv2U43aB47y
v09Q4hzpoWmLXGXgYTheLPIjedZCzFHI9/e4/YagZuxDLoljMsNn0MFK3ZfhGJ6K
i/ZaSEQE5le5rGOccdImBfq8VZ2xAiVEGl+rAiSgrpWgpCMm5VZVzf+DVHns6VOR
FUTnVMl4Fj88P2fegsbj7q23Vw3NqA41fd8uxNir2B86W66TC/MmRRhTge2owXQc
2IWRNLMjnlMSPL7NRwKY+BqXKpuXs/4jKkHvQSIkKEHGLZzHV7kWz+B8HY5O3rrB
GrNztwCrkgzAZSkXFJHEr/4m/2Mpg4Car01S/6V6Nzi+cZ/xCdw4b3sfZLubHh4m
i7imFJ8euafw1ON+MMAuZNlLPgOzvWQCs5e4moGkQUF7tlq9M10vfYV5r+6Qc+Xe
PSQAOwUAzBDchRTInUxms1qtaRbYfYrBtdtM3NXgEQNXda2ZBy6cg2ZW/i5VoP/W
HhHzZpzMyuynJs4YxWTNe/yTGpynVM/F0dpKisjN8EJy6mZz0KSLK73YvdAZPCKT
iUVTgKkDy1gTyyifRonZJcrinlo6qhQwXcrvRe37LlMQSBBFOL903nIUx3sKyoZ/
V3cbunpUhaa+srEWNm8b0MUAX4P4VBP1JceouEkM+8Gg+YPpppiYOfp84TyEI8A2
EgSzWE16qMUAVvVZDo/iAB5BzDMRQE2DGwrSHjCxRWboCZQ2wOBOsa65bUwVJ4FW
jaLYUo578tQVlT09SWwGkl/M0MDixtFpGxMDFWQ17jIRvotI6QObOTUnWMvi8Sz0
QMxdGiwwyCWoXzSOdpYYME0LjUXn3VQKb2/O3DBtyhQ/xcGB3qAR379YtWm6bl2j
XkGZMmVRsVVUF5Vj/jYN8U3JiGn0roMbYRxg8dPbgGK/APpYCbdXSEUA0rI8VJEK
Nl/dom404a+kKd41N3Am4ogAF3xpxQ3V1djHcJ3UMe/Hmq/EOm5DV5aQKKB5mPFp
+1H0iYEeBR5VLTP+khHk2tVVByT1ihuSwV1f15zG0eQYN1YlikwvyMWhR1FyNins
DBTejyPpWB2jkD98RvSTHEIqEGysXUjp0eI900DzTOZ+lQQND+d8jwtrLSkAteBf
DYr6XTkEjn/5yWUnN56l0jF7L4pzYyzC0WPoQepr4EugOIjjfRG6i0KoOsrfmHmV
W/2s1pFkR5GovgWlG7JcHVJVbL1fQGsNk4zwt1g4ZxBmz+PbD11P4ZUiBPmfq3BW
kgCs4u/+OW0HuVBPSEPTj0vw3OSXR35/Et8FielfzWvR8/e7DRI95724ERs0tkT4
m2Zs6jEwlHVWvqip1i6tm3FDJli1g9mWO8Zmp1Zeh4Gn35o+rHKQvJtKwuQmApqv
3gQsx9HTK22r1aR8HTi7NTdArCHMYdcAfGgZzh1mAurCu9ti+HWMKvFToM/UeT4u
8ts+UmRpcxRCsCr+CsH5COtz9TAOP+w/EM96/mytDYaqj0PbQhE8KwQaa0tS3Fs9
xJ3aeYxLH90DLk5oxFWyzuIm3NEVGk3xbtWQZ7vLcAVlMYwNoXP9b8/SC2h3T5an
znuJ+EMxxhdAwuj7PmBAlJygGFV0EcCMkWjGG5MexiEVS+wfXfy1UHVGMKF5FOXa
NEExzlCuAgUr//oxzLYTgdyEVQvSOa/TEUDvwz00qkcIpS+AWHp1ZzUooee8nDT4
mBH0mlUd6bBw/iguGiHXC9ylGM2I6KQdN5g0aoXvDJv4REMNEqcTmLbgA1fK9ZhI
G33SL0cphUAHC+HnazFNJdjCJWkRxPui1cnr/5QHEbZvLC8aU/iENh78rHdM+4M3
8rfZuIYlgewDgmJLXMaOGaxwXuvVLEnmorHgC0LYmcEaPgPOPku6otqyFLKdrc2+
aBP4wCivAJPrr9Me0Ar6XO5S7JcHtu7geSzMJROoIMskzAApYHHeLqcSkMQ3zQEX
fUbaApD57dGfy0dKjjXhFYynkzUACkY5przhOHepnuTLRL1KpmoezTcPqa78p7ij
1SFCVB43YTiQpSEsvq+BUGN3o3vLuT7D7mfMFhF2qLC+QuNpeAjnh285FfhvrpLQ
pg3IP8CtAd/hUgXHw1f28sKWZUfIrX1AZaMvh32+NYXzhlSjTwh8r6lAuzLvuN2t
B1k324wYnCMxArnokgTR5wy0hVucBpsPGznZ15CTUHDODjRBbjzzfm3ITBdeG2Ao
0CPW06BKJyGUIjLdwws6E4u9G51cdpVxnVi/+l0I07MijKTXxt5YdC2x09vhsI0n
rQF2pQGCaUPG9fNHxiFkq3ssNzcQ9/DQWrYLsnQlcLNjtNhIA+wtdMnFIbfhpWCw
7eIbzEtT9OxWqI4UgX1qjOXBQ25uENWL+Dy3quLq7h1dVW/ptfr9Nv/wEFTnT7KN
16f+ncMh9NPZx8qOhDEQ9BVtX11yhtgLzv4wqwh+D1YNORp4k+B+sFsT6UPuhJYa
Dll3e+/tlzvB0bkPWgP/V8dc6fx7TNJwud8PXIpPIfyINdGml9vkS1KAzsk0sD/x
RmCbuXvyKNLNMrTQKo89gvGVHyeGcjJUnqJHD2bPpvQutbq+pYQO8UssvCkTzdVp
NlzYyE9XbMXf5uegKv5FKDxwSzE+WNILkJH9Kcyhatj5G3LFAooDRVReZ3I9TnwV
yls+uEYZqkcetN/zPKCGn0xv/rCCaZ+Nql9z49fscSfRFk5I9VgF8fDKYTBW05Cf
A1EHbx59AciYl/n0YyZiArzl+JbzCtf7dSk1PnYXqJsma/8EHX31WK9kbZ1YxnB/
/cH1rYzgiq/7vAIAoIxTCJB0nx1neFyCkl02Wv2xgsM0pY3j7Wl3rFrwSKy7yout
oVw95uoElku+zvvb/bPQgpaNUhE1/V2y2/wh//yrCFDtU369xNZKvN687+QX2ylt
D1KVVfQeAYYW0alUEJAyVAWVD7JFfFB9kfEi4NpWbnJMuXgNBeeH9YGQnA60iIrp
yVJ5R7z2K5RZBjlsoplgCLTYKUZ1GR/6yqHZM/BA8EqJakYbQ9GO9tVhucih59or
lB7gfLe7hdEv3XkGXSbw6gZ5a/Wul6QMokdlceaAOFp7/dLhbMLRPz+X6HPBGl7i
m7RkETZG34OJlLjM3srcgnUK2W1z7JaUGLOgnWMehQsOoExWbXoQufR+B0sjGpg7
p6cF1pr2OTg1kYqZp6t8x1IkeXSFLTvuG6pTwCanAo8rGpKXd+C+kibSIVKnOwy5
sSIwhSx+4cu3qffXslvehhFWG5vlRXgMg2Dr+Pa2fxCcSsP1Utd4f8uXGOGLgHyq
Iqbaa89RnXZTVEIac21oupdXva65A+MP4YKTN1Za5ARZo2D7K3f66sw2r9+pIP02
OZWsdGnUJ3eanwu4itFJumHDzfXpYqQBbOta0LxKB+oncTfTQwzMFYZiimQHtL5g
EOmCfiYWQSwV51+iuYAMxGYEsBhAdw43xUcGfm2k87/oUTHuHR5L8acKcsrJVm3I
DWJF6Sws7d/Ve9J42NoN8BBlEJkt1SYk+Cr7duAb9MFleMTumikE5h2m97RHfg2q
+V/pcAVgMZq53TTWsqdIPOXksqZvJUBH8AYgTh740RSbzcOiZpqZqOQdUQdBUmGy
f7edQZ8wlOJascywElVQGv7TCY7r/YiGgj3j/6CbGbn1Mi2OBLajAjoxCI1rH1hx
rpJ6543VOaLwdWsY/OYtv3jxf2GD9P1x219wi+MedkPEFZJuyyCvPNtmim0Xie8V
TUtinx0bzPPPe9+6UJasqDzDwi55sOX/d6sTm9LTftpBFc2pdfhCJr/0ctr3zC1K
tQzS7kJwkz/y7AaD8AfLiO3ApdHzAZvg7zInocOjVdPlQztqzkpJgpG3GGCPTOWS
ggea3e1koFlrpYXwrAFQfsjEtGXSiHTHUkeqZWWVeqFmYkCVbqkwU4U0yoMRIxQ1
kHAl9hrQGA1Bs3cfdjJJAtQSNe5TVblHzfteueFJtZpExMNSN2nT819UVYES1W26
DVll8uIJM5cAL1w8gkPuaqZr0teEsRemEJaU9nY8JhXS1e2RyFYBNWfyttkLsiGj
beyXMjODPk4mrYVXYk+zvQU+WG141j754cPLbk4R3Jk+KuiG4H/c2azWVjsovKAv
Ni4oFQMhLOaDVxd8+3Ev4JnnQEZTI6s0SDB5nJdylXl9pNvhN7dJiJ5qJgFYmDkh
nfUzEMSsHTYrvmkNnXRcyACaNCfqhxacUuqLbgqm/cJfnPzA3QpG/F4O4v8I5oUS
Dg3ISIQUTbexre649YUcFTv1M6zNRw1hYXv5gstAodspt/t913cH7xbesxz8ukmS
GLk8+CWLZ57A+JNWB+P5wBO+Vm/fcIWGKaiyJlZFfnXhE7lh2LXXSZ2SqOQtjs2F
huQ7jZ+zD1oFuWkNmDsb8D7w4Ev6ihHyc0ac8QtevjEeU4CkcmPEnmCOOaf+RaL7
zE/XA6tiBMHl04lgZADunY+0WO1y4DrDxVQpMfFivFMC2UKvwPEEVMlN8Nhej3dp
ZmyedaZ+KfB/k4vU38Wrwt2uTLTOsOEth9M330dvg9QSQ/jKMsMGiX077GdEXePI
Ah55lG3PfooiWyqalgts1R93ldM/uEFG75J/JK1xRQRV3BcWExd74yjo6KZEEcj7
pLnimAHmnFNMMVbqLftA8BIdJ5ldMr/V9hF8sZKWysMp95I5ZRCTd2Dvdxt6/Al9
7qLH9nNi2maqGp8yUIPf3rx4vFoAg0LPHnplJGZcx32ExnOsA0Rd+qh9ThfOuCc4
RbnqBOw2rkORc1rZOzrtoe11akWUr+TD+M0EtvqPvQz2pda+1BsM+AmTSbyEPalc
F3OMJ7bZWB0uUxnlRboSWBgoqnFKUoQI3oPuiK9Sw0CFN0m6yWCTASoaLE7xK28S
yPwpKwk6mB7KcNknT/VV4Q+sxQ+C18cEHDGLjLK4WXhKkgZXA/Qvs2wbSLIbrW2K
Dg02vtZThRxlXrP6wipWVDP0xfvsu4/+9uo/5AKiPXQpz4S5q7lvk7x8AYoTsBbM
sHdXivVAf1qw/K8+btYRCsHQ0MBLm0y0WIr74Tk4iszHPmTgGX7rPms0endqxdhK
c0liQ8lNeI3kqZ9aRavZ5BTmunUL2NJ8L+5d4jz/k6mCkG3GRmgrpZkqk5S+tOFE
Zv174a3Jwmwt9Pc5t/giKYK9JLDCX8s97Y2IlbpFlsErKpYjvkFmqHNQjpkUMz1B
zlFMfy3ovXC1XcOcccqm3AFo7ow1zzowtthQ+xIo413HxfLJb5ke3HrTnR0ypvD3
DedWTNNsBYuiPFzKwHdMDIg4csolY+cVount3h9Q6a9gDgVtSuK+MOXVSGbE7o5L
xoqD3Ox7nS2RaqHtHpqUcK0oMgsK7wsciPFt8pTV/upZEPZ9e69AFn3i1cezQPF8
iEobSlfzipeuQ5JsTt2zsOa024GP2Xobp09KwbrvFCQ/44j4hLCeFlSXCYXJB96+
BkA+S/LzjtUOhpdm0eSYt8q0X1wuogcCjKEw4nnIDBQxt57ttANGsjFrPNWyGtTZ
OPJtfjm7Ss1x+Nrkb48Q1qIBvy/q2hmK7/Zwiag3aNM43h2iQnC61rB5U3UdttfT
pesL4y0bgHhlnP/p4T3onphQCNY0aU8ZqCflrFXl+b/seVjmtopAmNBMy07sRg1S
gbJnmA11stX+H/kdmp6v+yc8xvcqVo2Mits47GOZf1zWXF8wgetUAX5o7d5SpyFo
h2wHa2IOgV1a4NRIu6prkAoEoZS/YysLjXmcd6rt9bm9ZusRWNolhTGCMsunVpXH
LCZhWWNWeEiy1TbiXrCIAP45OVZIb1LrNLiXtabbHk8/k0XsBpUVLBpB2UwlCZ3p
A5OikVTMN6P4hvmQUK/lZCsMmJeEvMkydVsdpJMry9dZZbxNYHz3NMO19EItNlCb
S4Z/rxEBvTSnz7GHSGK4fPe2YQY8upYkI2YV6wrPiJg1436WzAtB07UFOO1le5eS
RRbF9/Q4TdiLLdHktrCRioyepCrt7M3YX2BNwIWIc5tdXHiGaO6vsN5bKYZ2uN7l
eVQngg6Qhfh1/4WZVrbxoLuHRc5SXhAxAbtgkT34q5UcVAMPUBF99sByN8REuK7G
EqDqLes2bWXQuJnp33naQdpKjJoqQgFsq83U3qgqV+zFlwPP53KhOZTDq0uq5xwj
5EoSuoNLFxqSz2VmrpGXOujQVWV2GXZVm4MShf772O+XaVDw6wcab8AdOUtNd/wm
jSNTu0q/tGBTG1vxLWMSDawvUIWlCYGZttwjpns9lz2Iu76sq0BTQ60TysZ55e4m
Vw9PVyUn1FysAmcbRIc1bspaQFXeskVQOuG2asF+1HOrOUFxuL+dYcRCRS+AzNAh
todP9CoVf1pFm5TWonu52fhGQ2mAeg7ua/9ezTzFe0M+ZFrB4hkFH3ZmUUIxjIPI
fa2NkL0muUyWQkrPBwefvty3iU/VZl+hvoSNNR7GrhiqlCR9+5VEE6e1on0axWa8
fDl/L5uudeWButFc95uNzPp7eMNYlwFYrcfI22jeg+d9CjmOlYVVJsLaWqBLhNgA
xMtKbxGSDZCM8hDY3OKoHeBayVvT+zSkVs2ngNsdXlV4WXAZHRGpTL2WCS7CU3hq
l9Iss93v+6jRLnwBzsVmgIJPBJv8yOO1b2764wCp4TIcWl78BZFvVarnHe8jV/bl
VkMsieO8eFI9UbdejAI1nt1b3WxL+ti/pX8cx1Ega3y96qMu0SlnwLI6I0SEIwvP
haNUxj34whnUCTkP9bEeJAqp+b+49Xi0J/yXFITnueW3uzk8VIAmYGWvzj/7nWJa
NYCq2jC5Tc5l6AX8PPPIIRUJJhEA/M1smEl9eSNqIwnJFmYc65uWaOp7PEtTVbJ/
o8Axb6mfUXR+9Z8lMZJ0kxVmZQINRqUVVSBBWQmI8HVPiJs1E412xT4wadO8tdVj
X3ZFpOY/rZmRH6VtSZxrXefWnChcbpA7RJXYON54o+jj/yhFI0lD5qKzWm90ycel
ibf1QisHr7RXuoWeigaejEMYIC/fCrgPmgzo9+i0ARbD5c1+xOFvNZ5I6U48ZyzC
7Q3Wq94z8qGBtHrcSlJeej6UWFRzSRSdoqbjdhVDR3TE/qkd1eOVmG78+N3r2xu2
J0JP6sSuNaNahQESSvClnFdIzimPGY6LpCkkXz24NMSilXIRXM2vSc3MTSyZsI8y
qJtL2FkwqWYouGXE2YFUcXjuhsjORgaBamPycMrUsw0S8b8TZuV02ybBtCaGq3PS
NUTrJ8JROUru9GPHYB3uc4fuo675dWlfnYalV0Itpm3+XTogYM/LAeQRtRFAlya+
EsQ57BVopf6QTQRp4olkxvxbTmJYvE3HACS7ENYJJe++Hr59RkqdIJ1ZcVzBoubx
BwfJOZSE4SI3LW+A2UbwWSkXSqCbwo1n1A7wR++4ZoZuvKdCgVLOisLKVv1FwSsb
WM7oJkUPHvcdiq0QVinlOY4jgX+VFN4aJTTg9CYNR3rsTebihSJtXx9tzkSf4VKr
KAqBQZDRlxORk2W2vmiW39MCSZzDhtwM7nNVcfNIbxrYXdVuANG/wXL+hFzHqf9z
l7GYbVJbN6IDsZFAe+8/SXwtvfZatfPeMHE57HD5ddG7yHrNxTSSdiIOFb7jX/1R
Z7gPTLXWY9VU36DiSw6Q4jbcmYLLHO+pAebdBI/So54m+HaIc9RMULyyoclo/RT+
SnT1E7K+yJkqVNj1F/PGr8v/pj2p5Yt4l8QtWjNMr5CjUfhwA+NFTXvGO2gPgPXs
EPkfR5L+HksBzRmDQBD/q5E8FmaQv33J92jyZLkwBXL0Sfi4kAunPgV14GfyD2o1
olBqujbCF/HxZptbm7MX08hk2oBcrVi+s/frEYh8nA9Z9U8ErxqgFgTYSDxvtpAa
Yyy68KPg4l++f0uhMUfUOTRpsQPDtd+kEtbqtvxDS8eR11QxFeBUx1BwF2uu7Rbd
Mqyv2P9EA4lQHF7EqiaLUxdRaDVsDLdMStcNzcQwkeSMRmKv2GTqmhvEuzJuhJ6W
N+XB7EszPELto1TAz5tW922PIZ0reKCH+6XxmiqvEYsMxGuWHyBIJ0tHrBqy9nKv
uT1UVcBT0M6Ha8dr+4Vb3ff+vzcPlF6AjtohUL+aouteD9oL4Ve5mqUGdl6zrTZu
U4M1InKuqcCVkqFgdByyEZHEfyXOTnnxhyem9rejkUn+U3IlOTwoGs5AfN6cASh6
hUSWQkJXk81JkEdw5tKubUO2tYawVW8Gqt9Gqf0RtxyXTKx0W0OddDfUmqJVRxIY
OmV6+6GuWuIlJdWYkWKVWaGaAIocc+9OH6/tbPFqI/UxNkhIS8y8oRTT492kHFhW
VhEPPS+ifDXi3GYlVMsAOQwl/7f1fGQk1WflGQHlQH6ijtGXbCSn2SkwYI1GBPl5
Es+ujMcR2EV3gP8ScwWQXraLDUVf0isL/8pMBynrkEVLm5oUzUZXwIcNxfBKey47
GPSxdJ7608ZEqVI+E/r/E619Ib4kg6pcVOIsjtAa6NuyJLj35hbAQnJzOHmtg8hI
d+KY44lv2aRS2sVQiP5Yb/2w2SaWIZg2XIIRAeuVFJ/AH5mLJK9/M3SxRtQnsgmq
TFmYTbQHAtgW8uNGOrHoft6T7yxb9+uF4EHzJZ5QVkqWDHOJQ/h5Yq3vi3fnAICk
PhhQdeMOxe1AF7GVRlFpmbmL2FLTgQ9hGpRLPsAmEei8UMIrKI0QJB0T1aub+Ksq
BZl2iXeSyECFmv3aLE4FCLRI90olCmuNZoMWF62YE321q+ST/9gp15nq9grZ+H1J
x3d0FD9RiwIRxlmXyyNmtu1Ae/XBo4nT3GAOvS6OPPS5yAFdkRTE4i2syaVetl4o
szze8g6ZbZ9YF8mKNLAV+78C3zFxhtvz3h7+xlFaT9Fmvd7jAmdQiXP1NczW1Vui
Ep/JpjhMLnnBEzLNfxIs5WLHN06GNTtUDCG0HcFDYGg4Szm6Q/y4J6h0UI6RMHE9
oWnfDzdObL8cnTSrXScNuteyfx/NORCGdQ6m08ouyuDFPQv11Q9X26ywXrtWR6IV
cWUdZBS6WZWfn4kFnpivd5cRlDtuxLbgZafT3ehRqLg1OXfKhXVwGb1PcjVmv5tI
Ga/SUH6lkx/oDOSSiP/0f9VhkHFgPcE9YSv8phQH3ZS6wCZs19SlINT4uFbViDwe
J0bwH4MoXgUo7iU2cl1vLJ9rOCL5MKmO/vJ8jUDUyM/ZAMktb8CKZHqtXpcmwr/J
psvFa94VEldofXzPur1TnG11bRJKWlvqTFy+NqfSCabkNbQ2HeqZsn2zIJJYgbqh
XkjLQRBiCvazM5S74RhxkHSWDkSGY8sHqnZdnSMgOX+N22pD4KFMrT2NtgFZhhi0
XiC/LU5cKUxAuFAmGutmiY728qa+XxpZyvEvqxjFQQ0mh4I5pbtn6ngifk7bVZxS
e0Oqyl8WI9+dhm5AfuxKw9ROgt0SJC/bz9c577Zd0EOQ6qOyuMuCbRaaNLQkmmwy
LbnMqYdbVzw/ZuHZzcKSx4Xb+jn3MMgTLocQSq470rU38H9/DPBBcVGigzDcCFB8
LcY8dRTigCEzkZGnG6uqBz6wzjic7+nsFg0nLtulXJJP81AFVU+DxfCaZ8YlDKRI
RtBZgmlDIE2yZucg46jeHV1aFiz2lyq4Xg/wDZydveJQSzh28JTuwWOL50Z6+Km/
fhtyKo7EZvNhhGC+1l0MxSJCEX+jtt/448Tfd6nWVQ0N5ZGSmVWs2mIbCxAsYx2A
s9ov1fPnBXLChbcpk1rbR1tESChozNaXck/gB6SNV3IXDplQ6f+wcJCRo+88BZT9
cuD6IXqXpcXiBu43OOk7jOnbmlPTaIQs5qwaVDhOiKUSlJlYaOPTfvVdnTUU5EKm
8BwQda6cEpJWbuLq9Hwvi2FqjxFO6lou3BqO3cNwUhPAtPHBU6mg/EC0KNRZmtnJ
hoA8+DxVfz9fjZiTilmrVtLwjKe7tJhqc/COtQck1aIvWbnMT4ebiP6SFqzzJS3z
SJ71D/0tsg8i1zwVyKBrSoj93JT0iW7d1oqlLEugjUvqAzDVMC/I6t6TZ6xnWCrN
a/HgwTWrcvYe3hhb6YxfyEoDrY6I8/NkfaxP9EtR9TUCXMSQDoFGtwlKFn5c8zF2
gorW/b+f0MHQw/t3wTWT2eqMb7VFydhX9pbTBXwk2MC1BqBysMEQcxIvH3ubedYh
hmlrhXwA5j4f66SMZ9PnHMS370yXrZEOzc9GzoV7jkFBYCaUXda2bxQf21QUGRZY
jNECSfF2qYHOEPwpbizSKHp2EGh4flolz+q4HhYD0h1eh8qcHzRdigZpxphOsdme
qxp9hEhgG6newi0cgVqFyawoFNLZMLpzzV424K8icCoSMDwex1Zc4mkHkAJCChpI
vnY2HwDQ+T+aWQeU5+40A2uYwgtH91f/zELif9AZykRPVIiR0zoyQqjxzXhbpUC3
I+D9c7/sF5d+oRmhqYFR1/06SQGz3Ik0sH07lVqoYqbCa/i5yE9k/RsTc80QSMLB
qO/Ma+/kr7oz+HM6uWOxrzvp6zzZOEtl7+KHFW3NIZgpqEbTChdi2uxDroNy6cDk
3Uan6z1J0ILwigAjIr2gCayvu9m1TGnU/C0YS/J45Mhp7fMS+qOx7XoH8l/PeYGW
lP2pAKMIMFtdYU6v+nlrpW4MBE5Q+JCrgYSwKTNmBuF8+J2AQmcN5Ll/lyJ7wUaq
iVvxMseyLWuaVWqGaucJ29m+bRvQcMic8zVRFmKnm7NWEM/LTfqQ3+Fcrgq9AOdK
nfi8w+3pIM3tBJ7bFc5704jAvKZA84otuR9UYrC+gcaL+BV8KeHrI1swUtit+N25
1eRB0EkjN9NeTOqgDlxd+lXTLBBNLR1g9NHyaGuWbz+hhgtR6gUFruhGbsA+UVNS
U0lbjGTDUx/ZB5p6dGD1XrnFBksAU+FXcKFJS9jY/To1eGN9+othIXl49Nc0L0k3
557IlY32YMC+wiohnAAKltbBF4xI6AGPDDsoa9Wk69FN2WehKPgDg8HdYka0fOK2
WQrbxE1o8IBP2hOqrk8hI3NrP0n/U/O14LG7a8f/tvTMMN8heTfHDEyAjmqJUpPH
MdJ41IBBD+7mtb3kuk1Y03ZE1fjm2G/t4sxaTMoLeqAPC0dQO1l3PozwZ1FdlXPH
7tazO+9ntw/6eZ9dmWvGLNuRbS3AwIA2IjDDDb0r42RAI8X+rY9rhkaCIXuvMmSO
TLjNFUu8UeKcHsotLWo98Clbt5Y6ZUvwH92b62iuL6X+NqVQVMauKM1i5BBwOdlj
tQ801rJkAakIUzfZjHd1v30TZ00OgGlQGlPyNUbKZNEVkxy2NTYkvzJWW18bXg7a
xlojF8vdFE7qyZ8Xp0C/hsBiW20vqU/IKL86Ke3ITOcjhYeS5uV0FRzf8r6RDK2Q
NX36is0NYH7Zf5axF6niv/+cvKekdMjcg6OOwK4jhE58b69cidocUxXM5S18qeVF
UdCA4TKp+olUyIPHaQrgoxtB71dHFXuVtsgp6ZL5kZ7L5vYtNFg+ZKGFQJDEa2Po
fCA+7whQqS8zavC8FF2nCGstdxws2g82c+axmsR0rw/UmSexuPLNSqxWQj5gX5IN
eS+pDyt5EljeC1wno18h1AgCXA6dkr3VACTmiOQNwoi4q9fGkSnsPpt4AFxKShSB
iztAT7j9h5HPCTouCMJMI8yetzrWjfPJyOxjCR9IRbEzo9lAXAVQJgyack4xck3B
TzHK8W0iMjkPD0/uINvmHOrAv2/lVT9cwlEgNy9KMlsC9TQUstdjBKeXX7C6++lF
wfkhiIyguFOmIRzjD6jaSDH9ui4KKJ8irwnQK+Esqnk/cIukEK3KB/zplVM3WDq6
qu45j1W84XNlEXhSBD6JSlNSOqzEw19PzbjBH3jpUvQxm6o0+EydxTm2TXGRbUGg
Z+43BsJMUhQomcJ9XgcxY2+faHLp08zy4Y5U077fStwl/ez+GxR6Ua0w/FoWjkb8
kK7M9z6ilQh4E8QU9M51APMcv3Ic5xz1yr/5zTFdxFXXvUfQ/gZPdpcMZNG9yV9O
qCNPMPOgadtPmC00J7kfF1VllHDs8yeSNzz8P7zn3D+fLn98/5z7oTw00MBQAB7N
GGHx//Hx+gF/H+UNClBjKgJazphl99QW4g2Q6F3F45vf+sQPjU1mEoMS9E+H9uID
rBdvMqnHlvvOSmJQ7DCy0Mk2/aaAoAlhGE/8z8dlvY3ToyAoRR4G3ERknga+dNy7
aT7pzaa+laxNybvouyy1b3bvPWmT8eDoc8K8uwMVMRcdRVcDeHtWoT0DIPsH4gvk
8MzM0uJdD+4ANxT50K7hYmgK+cSFglnnaxtCh3snQRlGUwtdEi7VkJFrvsDqQOzJ
cBJFDSaKZc8es0rL86ueUeTSsMCU1vNf58JhAM14mTP+w2Gg7rS/dn30FaDSiara
896MphnErYSXAurWASdv5zXfE08Fqs+sbhIXqF00hijqSUiQwdL1fyvNm359v3ei
Qx+1536P5ZKhV7HrKhUM1CwLhdPPfaHZc0COVLjqXnAcg30WjYehi/LgyVT3eFBz
cQjIaPZQiZeJSO8nt+ZA7RA/Ih5zkNEITDrTeqfETjgsAOXTo7Y7Enp5sIa6FDNh
o2FO/30T3Rz/ujOH+qB8l6/lLRWW/RiooAWFJ+qjuuvOaxcOwAoT9jbCR2d7kn94
QG+vx7FZpQTJYgIsb6UQVp/gcniLaIP8JCB9u1ZmQoV1d3M919TjG2zQ5gFqO2cQ
tCex/z5sMn1du5708cLm4KcFNPefYk7T2MaWoCncBlF9zIB0EOW4w/Y5GoXFoevB
6dCLYrVQz/41hjcC9XUk0js9jcDwqNIieAvkVn1bHMHDBUYknrCCwtg4YSAitUTX
RPuHYAgRH2kAoaVELBlI85T0TvUshBHwtWlBbzBYrfIevGtfHEDw8tWb8eLI5LW4
JQIJLPxxZ+Z559XmLv9N/WzCtFBgpuZMHEAM1MyByVQd7UD8HUGdLq/U3tAZkXAY
FIEGNUwULOxu0reTnhDLECQUtABjMo+NfEX2kmpLnBHUA49fiO5Pik02hzNx9ZSt
8sfbtZo96t7RG4h/d5l2QhjYUPFJzpjlBP1QYGZjM8aP0DzHA7AMItWx9kTsRnUg
a8eCQdyED5/rVy4dBg4z94IYtCvCK065sPdWrh2B6F5zNQZKnXVHoquVE1WxR3s+
x2QabKhkWS3bPpc6cda/CPYreBHf8XFWz8HBkPT439C7hBfUD+LdxY2bUkQ7Rsp5
3JoOeQHnPTLb/Zk2OxSekfhn3r+DI5uHQ9Nd7bwwatzXXR7qIvzvI0mOPYjny/6O
0ER14FKsQfoXb/AmOhFOH+4YWKMan9Osj0KBal3r6Pb+8k69QP2RGVi3k2QV8fzR
rYL3cJNpH8D2c2Mac7aw5w9fJ0Y/V6Aj85lk/Aznf3epBC0JWjAS8+LPhR6MbfEQ
Nr/b+9erR+TNxOh3OHgrUdF+3fYu7jVczsij9NZsgnIe0aSMWYi2zuXQNm8Z01eu
XVlxuOXBmAVanUG0L1wNtVgVokzqJOlC8CAPvmxmtV9Ovq0VK1grU0mvVcS3b4YS
MEgU+dj9lakwjqMYCo4zwY+cvjVYm/D96FPWB+dVEE3XY4oggkMahns3I0uXe9+l
yTbFOeEuPx4vmfROBBPf6PIK2YSr4SR31I8RcYWRxjo2ogSmRd9hndlH9jJBgzja
5/fffz45zW1ASTqEnqMRT19Fu0hwgpe8hFogcxg9+17hh4pdbgQY3vGadZLVxWVB
K0qoHotlesywX2LCGwwkXSkijaMgn/nj5/Tw8a3/lHo76OROvuzAfpk4JrcqgxQR
hqB3oJg6pkJjHFun+gKnuKfLbFEeMuT/URnYEx5a3ojAnmwH6B6r0EcS7wIA3Ixz
n7sHk9UPeeTEvHQLzvgXVqhfWfAXdMxW913Ok6DM7gAMCm7S9F2/X7kzoGzyM2qC
dGKlZpZKC/fV4Trg1RFpdQgM2QKSBCYBW6BkrW3lE1bN5F4XDHwQovLkfsk2+EVo
64vizgtoVOXaKip8GO0lCV+4060GYa7jgOFyl3S2k8bsMGdMjvWlDwXHHtNaKGd9
qGOgVcZs91hot3pVTT5IbLqekDKs9Qbo9DB783dUv3F88/vHP471imx674sdUhPQ
cVhjZaOUP+CdGB7DFVCqQjsoBGCRRwsAFKtOFyBq0bxCL9iO772njrB38p9vNE4J
PgSPdOBe90fqqE0agPGohhyITcODVfxd/mmvYkpe8GwDfbEAf/kU44S2n/a09a5S
JEnJGdcOZPjdnohSt7UyD4NNK+RAnzRP70mjKwq0pVHcFBd1dWRgde3j/rnYA+8t
e7wJO7/uOwHyQge0SDLga/0uaiK8tVZH3IRECTt2OPJHYQ5ihnA1HGPfoxBLV/yB
yNw/PEq3mRGxgWSo5CfnITtxhmSAqf+wU+y3Cy96g5CTK5RnRU2kyhPxol2vaCWD
yDs9u1H3QABVfrg3og/EZQVPRZFlHkiBEyJrtb4uORHZ6NjD4eCNyNaqcMnwIaz5
j+ffQ79n9Txk4iqvsSimo48MuJTa6F48AvSRmf7jxclrtMWkBgOI8OUabzW3H4Uv
WKszEOFEgy9qBZbzf8/zetOZRYWC2GmrFl/Pq1bDQYmEAMgbdCizTa6VjCLv0YaA
KmIvq88ROJ5vwlm8QTwvuzieV7Hmp5BrGZOtNpn2GD9382m2kX8XZv5OQRJXRN8w
Ba3n4KrEw+cfH6XOVERb3iFwyfrUxPtMZ+T1IYitj5DcIo2bZ8DALPE+lt3Vtryu
ab+a4qen06Qfa4VIbaPKSet5MugROigG1Om5qFhLK38qguJa4M+TTl0Et+jqDpFd
4c3b9On9LEXAvHhOM5Sisjf0vRMZS/EG60e/xsgdtXCfMqpAv17F5Fi+EAbamhoV
wS4enh9n2xFHSDybqYWDF6wjKJcmNFs5iQlPstEpSOip3HEv4V9BNJZ1Fniu71NM
njx9g6YM5JE0SGei+AHGTe1DdzpYFM3NBITnBVZ8vQK1vEuvnJ98SVCSiT9uKY74
UJswiqNMewubP1rAqDoVB+0e+PSI9v+TSu8YvbqTyzxwYJDIebYLlU8yE3sV+i/B
aQYAA7R1VpOUjzh0Lpctg97dnE8r8VHPNvyXh4+sYKrY9x1EI966enAv+CTcGHWp
7z+ozjx5tUc/9D3/6C1azs6m8WRUsgms7u+ie3jGhVxETmv6iC1RfgQSkykTUnNh
b2/arOrHx0i2v8jdOl82LwKJjvBSWlzxNjmEheEvNOF1cqII961xBAxgHFIH/tbW
SWW99l5QCDYY+bqbc+k43/5eYtp2W2T6wKXdPioqj5vw28lp+XTDWQ+wsATa5Vmi
RERiUzIG1JPWnlgix3DwdahTRA7bWbug/Cqu99XLehDDWt+HCPO9HOWUo3fc4Qmp
YUbeaV+CXyOwmywDkK0bZ70MzWfU9WqAH8iKc7y9+vaemt2Dc0mserZfgbrX/Oxx
g1pcRzhDh9TDFFo9BsOXr/05anrjN8728wuHyC4PJO+hszYqnEDWLvvdzPGD9MhJ
36PCnmmxjinm6JFK0Zf4ptiS+3mP/fuULXY/FRYIh3Ls6yKHSAhsGoiVcZu8noTf
ka/Ia/jd2/d+4odknCKCLtcSFDqzB12VWv7EZnXX6ZK9co1p690xkxkPXaH4lUwn
9HE1EZmAKPZ5X1ke3kVuS9+ouGUP6mIFQ9XPO1jy8fWYQQMZlmVH9RxD+e/y5iJE
G+1RxTZRenngxmoaxE1TkM3OJCsh+6stsQMIaG1cm/7cwQteIPaZt9YajHZ5ouA/
pSL+twejrBct34ijXQedubNCHI+ZvFae40h/CDxMqj3VuxjswNuiBwr8za7SyNbj
nxUfgNk2qYLUjEDsSlvO+SoLEaF/pI1vLB1wyH9sIFamkbltw855DCqWpOH5UDZ3
nfMHTNHwH2CsvmjXNTxaJQJbTGahcIqF/cL45StzxzPoil++kLw6bO1oPP2/m6EV
EJyUPFLQEvnpzrZAwH8PcR1vGqKNKcNUmZ/2MAy0Z8K6NrT9laomQXPqMNtJtVIh
sM8ZFpv3JWBcFfW8Zq1sN0mm9M5iRtp9IKDe3NfQ6WGwch910ph5mQfuGLJygfiC
kaiPnYllQLeeX1sqhSQ5Aia9BUVqOYvAy/cKv+vlmvsgQZZ8aixdIQZiAUojEc67
SAZW3CWFoOyvYQeHILAHm2hdgYQE2t9g7sarZR/lT4bv1FLM9xsOE6I+gn5DStHl
TWs9iknjS7iUlaHVkDjP55GqwfEeOLZLCaaNH7ltVoXhzAdbf2zZs8wPjyRsaAnL
blndSR+IYetOgllrRfHKMvIOsebaMPb4ohUnzuusR/KMDC7ntzSN2n72rpDxKlRP
wxwzo/4burILlyZgRa36zOpiyiHdN8Bp/SINLEUEYmfcn7CsPkFA1sjt3iHMocN8
YDW+LNw09C5q0nEjBZvX82bNFQdvZ/k9ClU1RzAj4Z1Ly/jbh/IQh9Nq8SkGuKBV
+H8xLS5EIuz3vzmdbUcBGzTTvVJ8iZzAIP3ahqOYlHwcW9nT63dkjBQcWV2UoQ9+
y/4onG7L3zUSRvTj+AtDaw==
`protect end_protected