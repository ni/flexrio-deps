`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1952 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
lzUdb3s9JuxfBG/gbheUITCbaknzqCnAakXBQN2JkkH8pFi8Z/060rZGKS7AErOK
ZcEo0KicktbfQ78J2O49ShAtQCap6+bVo5JuoFKe81aKu3gQFlrq1POvktCKUn8k
DPwQ7FD3/6CCvKvPuVZtRO5/dfS4haouPzSelG/izftElBn/znIjOXGjE5ZiaX5E
eTkn4wWoWQf8Q9ODoKJ6FVpOACGuzzutTfYaIn1bjAlNtZeZFLAhw4uzkdaoiE/g
2iQfpucmiTcCY2LAgy/AS4ANjFJKtP8hqrL4tduSOe0iiimBNZuPGTYI68xo0iCj
kEQfUFcgH6QXcijLgfwGfYRgj0BUS4dfyO4ilplNm9sbBv5Rb84g9wWztPw1r9ty
BGbnoVFkgN3yMSFAvugdX4OwpYN9ObornhOUJmJaIP7wiyNsolS96x6leHSgBlaI
zEOsp3EBzsx9ZV5IXKa2bQL8OHCN66qRIJ09aXqZGevWkVoOMRW9wubQF+lLkXa9
9YRowPX6ekNPQnj4w05C/VQIqrxON8wxKacWF+1EwWXau02/weAsnPzjv4JUGQcv
NMAV5ZLijjVVwVnsQgIl+IXy5uXMs7EjCSiX7DlZRKrM/8ooJPDvoc6wd8PcIBSj
JRrdSmnpwkEYo+qIYJBiBEhCOBWdnvqY/B3biDOz3ECi0Y5gpnHAXw9gnm8KdWW/
nEvs452JKoaUHXzPMjx50suxrbdLnY0/2QGS4j+0csMnBP/fS6P41VI3Hn9TmQpP
3/SujYi6Ozoi8sCBDEnzhqQWH3yGVNl3be24AD6bcV8AJkTVVbw+Pz349/re1hDH
SzO4ElC7d2TtRJTRmrw7hrk8fne9IO7bu6RL7ydnqshf0tkglixOAViKJYP1CZSW
EFDvAiTgT/Yj4Rc613rRHdJHM1u50dVcoo5HiOLADXKNHkfc3Vb2Rrsu3OvuXnm5
hzpTn2OksB2QCt+23fLUjWSSsWAygkSauFtmFRAty+jLmtrY+FFZpFzNGlDDbeGi
no0N95V8IohMJ8ffp9giTWQX2dW8MI8CYa9BCkgbA0mB2JC/YcX4vNWTkukwkJe3
/IQ6w2aHNAf7I1+evpYNrdyn8G3HMjEBbri46JOijLEtX/shGpdxTtYa0fwXaHMJ
dDNbHMZfyyDF25FFahM5tQBnJyH4pLb+AXIxJ/vd+8TKW4gK4MXxmcw49Lski+Zr
BribDSvhDbK5O33SuCwWhhHS2p9XgXbz1emz4ypSDjdn5XuVPxCceqlq9mrobBr9
tWNl8hR8DhYgwvHKry++nQd9mWVp2KWaOjPO28Nk+BECKEqXt0WQyoeD/WKPYLeC
HawIcTvD+yuMLYI6i6gNeVyrPOkWsUiuqLdwL7aVbJJDQGiN1AjJxPIwlOOLeVTs
KTKaHWR8cSNVRaEFoTBSL6wAPpWp7BVYr1PkvtLWxE44r9rE2r5Uobkc8PoHqt8U
LaeXyohFX7RkhCyGvn9oCtZxAtMesPCzMVg/laEVcfz0AbVrbaWOFdw1HKcr8LqM
vp2Yke0Th03+UKy8QtxUVlzl50eBWwQxjBgnfXRCnmq4sHtqNIRuF5QijoeBj8KT
wgkd448vOYBqy3Rt+OVmCkDtgXIOj1s9OMuXRXFAfxegS/71uPZBDLGUSiO9AF8r
q7kGvmnDGyCyFjfo7dm00K5Hh5EW33QCsCXeBSCS12pmdu3kUFODn/FG+klvaRYF
t9feXUrtlSwPCkzXvN6kTS7HOhXjfIXsBOIDuEfzYXOpmb53iUFMn5vvDU4PsjLn
JWDsJpi1f5CSZMSyB3bx1wTDtmei54RHo2/ybaYW+Vgz/Jq6N9VYjKTin3rfOv2m
8miknPj16aXXkd2vuVL753coa3N1VjKCufPtI9PoZciMfXPkVaZc63MODVE6UI8z
+IjAjTc109LG/PqfXca7x/2XFQlKlY6Y5sCVlbipY14yy9+v6CHqABeiLU72gKqh
SUfA1kOzlGB3X5jqpKSt39+tdsJ3y3EPZykNtMAVOABcFZ8reQbopvHbS52TdBcb
2bQLI1eZhtcNOPdAwaJhZLqvDcjMvEtWosuWcTbCgpGERiNbrspxOK+Hy0l5l6fZ
XtVp2022HQu2CSAkaBpW4tslKEHtbwJujifYwP0DX13nLvXvNk3FMKiQ6SA7vLhW
df3kiU85GU5yGNkYJBnyVMhNP/8eB9QziwKuR+4Ewp5qI7c6CSx3/RS1Hv67qK6w
6oCHpAPv0/xJPii5vDmB/Akaq1wtg7sBk7ptuhBtMnax3DxQZZGp/tEIUWVLyuqR
GiGF1VF4bwW3IXisml6WxgMfJzgjIa51WjAi6kQNA5VoKKPeGhPumExrD8QLWTJS
r7TrbhaDb/ElPg7Rcp9oc5j8OgzVmxyK0ucLio+ZNDaP/Z/x+fk9xqP3uyFkkBKy
h0mNGSHsxhZT6GsJyRRV6qX62ApVTEvHqNLOtjlLUbA=
`protect end_protected