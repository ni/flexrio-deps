`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
gMcHP74wBZczB0bB0IzoP2xg5wC5NPjD/GsvSQ6VQgzYAsanETMwwsWi4yhFtJwv
5kY07u0WerSDf8woJ0stqW5xF501W3JLIS8KMiCOd55RHBOnavjYiaaLeu7oUCmB
TtTS1R4sO325rP2zOn9YwRbyyS5Ljn+PzFZZUmkt5xMca3p5NGqKtZW2dV6Babni
5HlLuF20Au601B75m2nv+ZRoGSrpkNElxoTibONmX8gBflpIVE7BehhHwaKSucEF
pp4QQ5zZAZjEC6aplZepouGVggAulz5AahlX5bf4opOVlB1J7IrgyjENtw6ysQ/q
DzybQ+ipztSXBGhmcCVU3A==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="jAI3OJE9Sh00Sic4PtM/KZ4WjwT98XM8AMZrZsQkxWQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hyw9IrFLPQsjvXplweG8O0lkaSLBN9Ijv4B5VdTRt6ipKJT9Kzsb5LxCKvkQyF9n
sGPOd5i74hRHnkHfYISGkfxGJCa55ieOyFShOsqTKRLxclm4oja9vTIey6yFm1BZ
54IDCG9h3PqfDiTD847UCSMRvFssyycwv+BRHQMQlFs=
`protect rights_digest_method = "sha256"
`protect end_toolblock="BnLuc3jxknmZOyxfJK70E5kp9u9O8IQ8cgkXv26kHA8="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 57664 )
`protect data_block
xABArkLxBOK6xG+7CdOOiGu0zbCbHMrEntFfAZEE/xRFxZaAZl1QLkuFI77OC2KL
XxG/mrHJzO3taVHgwRXNLDdc8ePbxbAiQfzV3NJLBO+gsBjmIymaCa480cPNpHLx
lR5W1Dv56y/sDQszohSaAdOFh8yS4TnBMvsTY6OZMGHszBFPGwQ/bs96DgLDz/oC
3b/JPBw1gOXom4Zi7+dr3d2ipccdSD4+sFQEkpfEmOL17UBtmKqj8nqqJLqp9ulU
E8beIB6hmPTsb46oqjDF9ibYQ3N6Gh9PG1i1u5fObvL3SJYZdipYYA7kAVW7/3fz
idWK4T1zE3DAPK3jRULs14e0GDKI56aCJN4dkoDr3oMA0/FHMqazkeOuBq4AOkDr
mSueoCf9mVtroI0/HVYKqhH41GP9qV7VqZJwNQfI718S3RpZJCtNgDQnCzWnTtM4
TUyxBApuPkOCMoU7gFpMQZNB6B4eZWbLwbcSeRdfj78oPPU9uzZccbPeNBBrxEn5
NZUEZrnro/Pz2ta7xRTYizszBX5VpPTZmt+Us+BWzCeBCrBaDtSdAUDvKHiv2Ymo
RzfcHCibEq4XgUm9DoXezrQclAIxryc0e3WaNt+jTEIEF0kJyjo5SGnIkvXlxR4n
wsuJMAk5uowHYMglrHa9Jib0QB4d4eLTawlW0d8pj8YdMXdVwDHezWfCOvOvtVBw
qkG8B+qzwVRl2PBe/oxMiryYxRFUhyYmRcAOFowPfOaURVLeTIE7zOwclmL4ASwL
0SO96hwm08uQKbg1gjxZr9WlyrZIjbeCXDQ8TGG+IJfTeFx6b2SuFie/OOugYUpS
ASd9asky4BY5x+55jUa2DRpJoZuj5pELuvqpKShOwUJbprOBWu0JuAc2XKfbCcRl
uVvSz/4mjOZHIlC27fVkizlVbzk2a7zvc2Lr4K2lg/k21u6Stn/yY5+69tsA+1AP
mECe/zz/WDSis71MXJ2mlFoUgnhyLaEoqb9o8H3qE62doBMQdqcx8TsWcRB33+0K
H+g0MUe9AWsjeCr7XwZb/1cQ6qxS3AGkituzSjpagyG4oSRCtsmDk7n4OKaoSC49
KwQPUzJiOD3eSojT9bjA9xtgjVoeTejoSbMD0kJLQQ1bndxF2esV2VsLh6kleO2/
SvP/WktMicS2d0OFE0fn2HpFFXKkDCbMcv/ZdNSqEPmWAf3Jt11N/LylonEtnyKe
pYeX3nzuW0muplArHCGqUWUZNu6kSN4ZVk/Tj+Shtk4of7c3UYh+RCui1yP6W/3U
Zr37uynK0ys25mWL+wBcRLwt+GUCB75m6MZIi2nrwZLKNIz8JVCtxVOllHcNjOGE
nFltosHiFh+X2OwEn7CZXrQkEEJeKwHctd3ZCkKB9nDFsRNT2IXwanG1VHG/G1gc
btRcnt6Ad09RbaJE10FmfC835AkHt/Vk2Dz7jQ1mVQ5xOkMNnamz8Dqj/whIuePB
eIAp+QiERq9JAhydgEDdBA0+op1IRndPchf+ivpjBtnyIeoWqoIPQHfVilyK6jKj
fWEmw0930LaO9mvbfQAccjZWVLXXJ6yKTl/LOxKRQiEsw+gqr/4v8ewPwSNw49BM
gIIYGpLJ3aEcvNsW1UCj0muyiYt7hF58c+ja7hDQba3WVvA9Pdugikdw5WzMgSG9
wDBFw6w/XMDgXiveaAt+5lIaGECQuxXBAe3q1zmJwQTzZ/0ccN2oFghJAxTSSoLs
OqNEMUPL0XRsvsBXK9r58/s5n2IuDB+Ek6jiErT8FfN0tM77ibqa+cIo6qSWtgVw
l7rpbSpBCi21jcKzvoo5YWmsC7/86GTIYLHrGR8T8cb1U5VhB/C8WW0TAyTJbpdx
XMrePyA5w6olmb4ZL7Odc15N62mYEjh1A6JXqcVrBTi8iqmkPeVsGDTvyyBex9Ac
ceqXFfLYR/Px+EPakvIJQZjg1prRcfe/YodQOkKm+iMT9iDLIyo+xEHdAHxnWSq2
w82WKQWXMgN7gwGwwYFEKWR1hMiS0gk5j0cUA37m+5lZZeSbp8Gg45hh7c2JHwOe
+qlyZkhOWqVqa8kogxzSb1TV3+c2EQtOXzaptyF7rNKLfpvg4gUhRUBc5u2pAmx9
woPZl1tZOW11Eq8TXUNtVzPMLz97D7rPSFMeFak3GBjMkAYbyUAnhtd/kM6FPLfr
fZ+w/cIcj62ltljda6yXWZyLZSXTIRfpoHxEKgkCja6JSqEkoFBFg4qUB2zzgEnS
VctaQVCnjtf85pY0FN21NEzq58QXmrcuyzFEX7DeXGOEPyjEfWkJAOhqtKenBVjY
+HDpIxvkr4ArcAdLIvI+pK4vIZBsza3nUeapmpWPVra3VuXObp2Ul6EoVwJRMa1h
b0Mu4AVfJy8GpLsvtsBVIoSWzi55RBRGJwE3YLgz+YTzAGJF2z4q1uXcXuIZjUim
2rhRdmTOjeuadfU2MeNZF5Jciv99lT11j/Nn9W8V0MYIiRFuYj2U9nsjB/sdK5w+
M9GLc0dCaxbboyoNf9peaICba94oR5lw2eU1MmfAIOSWnt8MnPhdMU2czlJHcm5d
eiPT8KuEwEPy0bWqgUh3+Gw2bLEVxzXFxQaIekXQoij92CuQp4OmY9dQZW0abbhj
wWIwxkhFxZeSPjprnidYtZxQTHQjY9SsQ0rG5z7gvSFYiXsvGGgmBONKdYcSJHoI
SgxteHNFBIT6pSaxVR2F93cA4NkylhWNTv/DEFf0zT3KQG78ggRs01sKQpE0xKwW
YC3EiKs25HsuMdkIV47DiR+sv0CAkDmPL8G3e78mtjejocqZxuskWxbBnt+nm0fL
Sdgt/tWIQT31Ed+r0bGafjlIE8BEaQMKgN6UFj5wEYkZAlWiUW1qC5szYREPtdQH
qi72dyLjByI5DWnVgkGP7Ftb4VJLiZevCEure5pYvXgYvrx2za2JCIbSmD4gXqVR
p7ZxLDPk1H3626wKCcIX7jIuQHbguWO7AMRCR3wgT7jiB+RUDNJba2cSbZhVjAP3
0c8tMth1EfCqf4fB2EnRSOlY0VIeNuqJ3zznYjOBLqMrsPa/J2c/l1wAIPET6VZj
yMw6T3AoIRxnKe+QDnWN+c8JSHNm+wiy8TRVjvSNVQDNxSQJm/siTJH5GpAkog2Q
uBfwpZ9yy721Y45b6PAvFw38fpOntKrMi7+9Xs4Z615xF3lPZak5VYzuWjcAOkUz
3NTclrg6rCV8fWjev4oozhiatKTq1U/mcDOL/H8N62ixmGOc8OOyyK0c8BJrr/i+
OqqYge6pHWu7DBEWH+Kod6mCeyCbabtmVDdCxpNIZOmLQrKSe5bwQHNav+BU2Ksx
x+uoPKBDDEBLqGTXoHzzCVQ1Cg8WceRDv42jkH2EYYWaX5OlV7trKvbylXx2zk0H
TGHs3fWg3o554kjCNeqXyn3LyESY/ktfdPFMXEbh7tY0liWolCjpEcj/i7gknbab
M4RCo1TXQboh+jRPjho7lFRSoNDMTNmmb5IWXUmsaHFwxD2Bshxo89l2ml/Z1uI7
O7JL52EzelbG+DBrX5D6Sw49wFHSQOdQ5H47Rc89MJF5NXZbqHwwnLKBdnkAJ4Uq
yS81zC5Y/5A7/efZgftyRL2kmkhI5VhvsyEtZz2ny/1vPDAk8TQWNzT5+9uH72FQ
vzYAp4QAL/iB020efwCtksJaKmjEdG2W4654/Iiz9hcJfCLkD8EoDCqj7sNMDM1L
bpWmFJlc1Cu8ivH0u74LXnroGX8ZY/LyUx6EZFMpW8u9DQ6av2zO+kw/Oc92g0Ob
XoSuMb1jTmHNHzW9sLKGybjdiEjyIbvUwtbSIJ5sjs/yRbLC7FsfkLtQyz7wO5xd
cl6zaulgTVWI6Fy5S1t5GWPzPWeHa+7T/u/1CyUaPBtKGWMJtdir7VArDAqQ3/wE
swKQk/pDS65flX1cP8PTZUFEJ/ToKcVvwpK+7+bWvGo2q7RY7JAxXrmKMt50o9mc
UTMDyJfOXoYCGdEn3jhvBthnfWe+9/7rXSBt1GduoU4hJ/471/GVjTMSE1CIZr4z
TuKkcRT7Z2ygKc71Crt3exBLLVzgzOxgX2q2ABcFU33tWSWyBIz6LsFXN9Buz8G/
/uItO11/aBmuZ2DhKE+y647O1yN0eMUBtukJb6XK5utGlCcZWCzg0tjg+DwtgNDf
pe5IrtEUhEvAwHLvybDJvR/iJZTkSO3ei767wmZ/Mfthb18vp5C1Q7zH1QyK3Ml8
Tgpsz53+xOi8lIPCLHxHsT6eed8NwaUX810J1yicbKaw6UOHNrlkJP6UPQq5iKvA
qyRCpNpxnHBnvUaV5xTfJym3NKGCpRrnBqvn/k+fS38bLWpgF6sP5U1OYy9EDdry
3jI5M0+Set+2OQzzndZAUiyb7PiwBFQw/aCQnTbrbVjHCzSfZGPPpqQhEQlMamWK
N6XRxk3D5qogsw/1QzuagaztCRd71UcbHj2z3GQtuqx+LEbV1by53D2Xb/frW05L
NpywFkStNHNxBmaYmbDsTYBSRvEyYlDLGIaMMVvp4yBAJPgRWRlQqJyJo1eaSXBI
Q4C+D0mAiep2/KKryBg8/q1gJqbetpkuWJCL+Dm2PYsrJh/mzraVe/05U0h/K6l3
ICmWBBrl6cAwQZUI3kPejiIkd1yNkCpyKTm97Ya7IoLPnOXCV+51gVcuvmDNkMev
exocLSlv77Z2vXhdwEaK+OsH/EnyrE9r03w9TC43q0RdY/u8JjybwUQmgnD9+ieQ
ZRl0SRk40ArMbEhNJtht89t12K2+6p9ojE5SO/XZaJdYaSYFxcPj/EjNQQ/A9qR6
xVzpjWGV4nNaNpNYzQNdrzJaUpGXXT3Vb5ujSoKt8EebiEydUfqL9mGUSiirDxPm
Xmg5GTZAqWXyC1xT8V0ai2bhzBu5EdBbHPAFwRs15dY6bTsamsQX9qLVyWpJjWDc
FG471M0vNbjfn//n48q97Wb+pqWoTqvrXCx9QvXZA3BkYNuMCNMIogonDuEnodzK
3QqRbohh+sN8G2Dw64A0091goujAAjkozg4BdFX+XN3ciGYxZsGxt83BDnH7wY8v
3WESclGTF6vQtUChYog6/+pJHdKbaRYIFzgPBr8esT4Q+NME9PIEqW0P3ICEGNTa
V+EKa3mfgWO01OfxY0iTZYXo20HOR3N7IdwPnD8D/WjQH175/5sLEHG6+XqdU18P
NcM9sh+B44jOabmQxeXhLA5h+XV9DNBETXWSS/PldpaIcIQuE7HXq7ysgYa9mxXk
eFEtzTHihJDlJDw1taOiecRoCT900vtfDTgV73rRVZSYvZIFkjbYaINLBQcIU3MO
X5db2mkCWccsctWiCaUmAJ1z7mV+BxxDTb+cD46w9KG6ggG+LmPCCyREyqgGCqz8
IbuDjC2XH99O+sSm5VQqT7L4TONdH4miNmsl+lbxVsIpS5YWLJhX04dhxHxm7zTX
GPsdNqWkmU+kye4uqMsnATdNxHPRLCnNEEGlcSqUQaRY75URDdl0TFsNkVFbAI+X
VgNFkPdNQsRuzC2XNtP+X2dq0We0anYFd89S/S29NqFlZ6JPh4H8pSPNR+KplfpR
89+iKhvqB/IzzR1Lp9TE64NJJ0OiziaaYkM8pSvZm8NVjSbbw0IySuFFkSu2Id7U
EbUEIlgohTtBzC3tDkxKby2MB072HJpnjz+Nmge4aVSJVJtAOs8q0gNrichqwU1D
+p5EBgKEig3vl7FxwLMHf96O/M2dxeN+UC9h1Ladjf57Cj7Jo/ZwB7/s2fSAoUCn
Qgrk5lc81FiDmLKT1eG4KX5VBB/eutzIn3t57raBMXrYyIgk4kH3Bfm5b6lH19GY
y1+6tRN/Fkxv9uM6UT0iDCpLHn7ifBpou5i5/NCd98R7rrk95W0mhiFKUFxP0oSV
Z8L+75dVuDbAIMbCKcEUH0UpUUapNlwBdcNp73lhYNqXfqAudBV2APz9c2RJOwae
M9LAx2EkhrszNEELt+n9jlKN5Ct44qPysffJ+XVI59px9KcOmNWnRdwXGDxHBDuP
t/Vo5Rq6TUf9D6sjRryLokkpNtkDo8luyme8UmGXd2+5kOc2iLQKMgNiHwgjSo2L
VFq6I47jKzNM88xhy5TwdeQzse/vPIfFtvW9ZFB5r/bjSStRdYYmZdNcYjqInj2P
ew1+fBgEv4FCm4tGUklgARQxt3lah9fCm41wtxfu+fEOtHGhRb8Y4FXbWRb1tRiQ
quliz+AJwV8vYe2rSwUWsxcVwea5b7LzHX4r+XansgC97Pk1g98d0iN3//cAMXqc
4kLxfPXytk4xqtef7fQSjwMh6ANYOsXrAiNSyRUl/jlIbSSwHwf/WWumfujYxd8n
IHkMChNsdpzvELiHTd/eC7c8v8f23C/ljMpPozIhNqUouf2H9VkFIncYllXDpmkv
1W6Drthx+/TE1fPhCdDZYKXxk9F/Of54Ag2pEmBzQiwxtWBlKDZvzN+BRHp6CVpJ
NuAJQxvCGx5hkV/R9BgFI7fY2XAhn/nvzccHRNfl+Z8iFm+p/ttIoizDqZvB2BY6
MrU9olc8ugbviLYdoIkFiXczmRxZyHhvrSve9omeZK7b+5B0sDMHeWld/7h4R+LA
MHudGuFdKMVKsi7k7rHXQi6k/lJGFeRk5ZK7LMJBd9FSAjONr2sLK7YJt2mb0R4b
l9i5/xGx12a4fwKzv0wt4XcxCOgEWPBuvy6H+1+tAAY5UxT/JPNdYJMcOfq9Fvta
xbscmgsUOXQ4nEpTHRSJu4h5UrQcgr9RIz9FmP3hL6GycQaoLm6G9OxGEYginvKF
Q9kRwbKcJ0I3K+0hB+qffyUHlOSfNcz7mxiNPopSiteAygA3UtuRT/xd1f5o1kor
+OefyUW6M0MhSLqI8SJH14PN4w4nqy5M2/r6/wYZOvu5LQhFLxQEI19Nov9qJyu1
2ejEe7Q7bL9If1hq0I6htuN8bOqOkhtmpe8SIlX/Ka/0nJ/3p19GAa9+bKrhLwBM
1XWRum2lYFsa6CSvS2dczXjm8ddic7aLfr1bUnkBNa2BglOafgtmTi+IboS0mDss
dPWemFdb35UgGhoxZT9CfdwvCkgh514qXNpUJ6EGagtSTC9r0sGg9bgDqkE6xqKp
EkDHPv70i0IpGgvl1RG/2JipBU2IXv7dy8Xa0jiXiKyX0V9vSEmUjjJUNt0bg3K5
LJJfWqPm9Aiy0DRTclkeHMNG2HD2iy79vVRGLsUOoXYJpt0vwkSQna0L/Zi2cfTa
Hsr5H0iIAk7cAlAhzZeDo9Ozq0OxLoX4UIdYbMAehizkG74OAqriFrO+Fb/6L9t0
trtKUh4Vjq64fjJ4Q51n6+9eD9aVoUFlBw6Ejp+uzvnvQKkt7t7PfWYrPrOZIARY
dZ3Opa0taIUvC/DvzaU3ee1j6+JnmHF12sfEfUS2/9EfEuYIGv4y8teYt7cb5llx
JVjYcsyPCSFADjWeA6STd3vqCuYzdjA2tKcx+6xm4zsOY3/vRtV+dfFF6gXm48vB
JsVGBdTTenyPDORYxORt3mfeSZPDRF+q2HmoeGgyyoosLLauCe0yeN6TMCFX0E/U
iEZoZWVmXSkoeCjfmIbapfV+q1Ha5gzNWVxG46Q5ujvq/vC7FEZTK2007zYgFypz
kWS65HgMvPLpv+wBp7A81HH2SedZQZ9Z8u3M3Ml7oMz/0Kkl7DTtSxhOeQG8Yu9X
GkjoZKcSzqiB0d6EKZRxJn4N9bCJ1dEiYiTSEQP2Yr4jj3omeHvHIUwnTZN6QwG8
aGhKNdc2sK+svz9W88izdvK5NawcgV6tFjvWAXywGW3YS44jGMH04Rin4x4nCdqW
N30h2L9/wLy1kn9Q2B445JZ32U1s+dhvHuwcxbru7atdBGwsiEvK/H4rq1/zuZY+
IeqdZpbJ1P+iVZ/8OdO1xsS4troxHvG6YCv9MRJ0Aj8B1iCZ9Qxop5wflBYZfdVi
cwF6yb5RPoGDyTLqykk8XVChrwFeVKJVeUKHkb+qYGlfbxGwdzn6LwvJnM+bvJzg
owkiLgC2ALLiW8rVVpDFriQUIzn9YIqeRRXf0SMtlolcP6oFNYzwY33uDokNMq1B
EnmNkeLwCN8g0EsZtvNXRtbThJ48GyIwrGdf2JOXEIwciW5dBsDqO7/qfW+n2RvU
fIEHJiaPbgjXLIFtSFDGjg352n4J8asWSbsP4ODHcMpTKfhWn7nzIY0YcyFr9hPU
dN8vvxFFFBl0lh1rqZcH3xa9EUrmQbA/+OeGcnAHn2WRquZizVHTChQZAAWfA8+b
qcYFW6htokKUO7vhb0hBfZi6BpNjGhh9CZrQ9Jf7mIF93iC8p+B79GboFh1EUKEJ
sSuhasykGt3xeNQ4mRk5hf/vGbrkTc93tfOMgiwtLUIqb+PqBls3FvUAH6A/z2se
wW61wj4GgbU6rmdlBmyD5EqGxtadFZl5dNQkHUCJ7ycTGl8ihnqOXU7xAyFz3Jmp
dM/cUI+Lc4XTsuv+wjAI1H1s84TcrFtARU7Ya2ZBVhkvswroN8hujMnOZ52fLTuD
vpKKori+Dn7yo/TYG4J9ltgIgA5JAuiWDReKCDQsJEJjifHT7sUjX20ak6/5xJd9
NqaVmLVWKQ3Z8vzpK3ANY3jifQHu3xRpUo+FnSxIyemAZs/quZFtNp6hbUTfXz2m
DMu02jNn+ffsU2uk5X9dLFjgQAm9r81VV81rC0ZIhrv/dlaWLtRl0J7t4IdcRLZp
H0ndIDgbILQVNXWZPj4f94ZjNY5Hz8uUlTP7tjetRLgZseB+9bwPm6bMM2UwIas9
Lj9Q1aNBsKb02qb519g4IUlWccVMe8zGyjEJr+WXIdubN5h1XFSm5Sk47i111KIT
/2g6xGMs3UKoYUC4EZSDBIxLCerFzJli2cdzvu6ld4hcsyl1ZaSmRyJ96WvumfNr
dfFyXzTHDQ82hKVsFEWFoaWB9zPg7wo2YgMKEgHAbHgLx9YquWN2PZf/HLRutECW
hbFi5xg5qmtl21SNJZYKf0Kzf87vDWre02i1QCeMRbidItvxIUeYd0b3nyWQ5lAD
La+aaILkgOARwghg30NRWfOxrcl00GVVdjic2L3dU+V6N+pA4jasqG27yHIuOZK3
iv+rAhNaCQ88e2rrw4hTDVucEt4TNYsoRIGkIYF2NAHu24coNO05ordu8RAqV4BS
jEtUJ1VrQOSS8A0ql1hd9p9EaCjwgOD6vi/1A8STdhrhwdrq0+Q/4A7FJWYD21rK
fEp0gofOzAnDkw99R6eHhRaO0vO8fFAek8mefdtbO5tXY9S/UGal82GVYmeVphJI
hzQcd4jaHvw19OeKZ4O5jcuTtneuSdgVnBd3jDVXcWtX66uAkuiuVAYQmuob3yiz
MU94hKozMdWOQ59an+172MbCmE7qAyc5pgtmXzqniGiDzefM48eALrcDp0o8TQLW
fEVf4wPV1Drp3DlpjvmF0fth+aWOgJ8zG6hXxW8w7/ID9dLiCGRQ2C6s7kOLBR5o
T59gnXCqhDXZfwfCTcNfJmQi9WPB+G2iza20idom9Ptsq0cW0CXgF8lLaQiAKqtG
1/RZssogdK/K/T0dBgd5Ce274teEUhFv+N9hQFSLlIVLHBaj5m9UnKEbpXkVoASL
wcUp7mWrxHe0qRfoXRZwq1dvCkrf/NmsqZpg+s2segBpSJ4nT3M7hREbJe+VHQFB
xj852A2bDhiEtQpGXUKV+E4VE3A7S9S8sdGgGjiIiojIY1Eb2HvShBE+VXhcvYdc
jd8M4SITUFWUIDr7J32nf499ZyRnQFColUaI8mXkyplqmOxuGFq4bkOZgnGF/sjv
FlGFk7Mw9TdeaKD8pvNjc5EatPQ35Dl29J4mRk0mvtCZlGOzjCScMZeUekPILNkV
MtWyUoIx81/NjyPnb7k7VUp+7OOHU8ksVLOkLC3eKBA69RllOnrIjJ3F2QGN+evy
2URv/KRWXmsMmxOTHu6CHalbqZbESkQlFZLLxUX46xbWbV18DB6H7ZTjSCDR+HAv
cKAUXSTnAM5Sbe/crFlpr9vA5cWnC+44SCqN5sim91I/tTBQAMi7qhC4YCXX0Ra7
N8wMPAcM6NF23p9/bt1ZAzqGpsocthWKLfPxw0ZnjzHt5VqWkBeGN+xUHtoWr42m
bkApMvn0wuDGSGnn7uBU7+x5GE3R9DxIwYSWDuMd1BhjNYjnQupkiUr+tyJW6dwb
2p8+ZHli8LJg3jVoscunaL1AyFrFzSe/RptJSoi70UiAm23Os/zeKkIC0fyZzsun
fksqlzICLjW5mEvMMr6DqpMIxWhdgZy6GDYBWtmXqmLxMumc5/So1km5MKAWoz2k
ZG/5c8eN/AhfGznkR9KhRcMX3YK/kpUBdhwS1M9AB0E/elVK8DYmoKCgNerPsFAd
rTQxzq1J5XwrZSjn4Dsfo7TuGcB/FiHhdrfY8tkoRumXtjH5qrmaQiqpNAferHCZ
rKinJwTlqwDw1i5SSe5bkLgUnInzWk4EfKlQxAO12oG5Au1c0RIlKZyvGJB38WqF
1HfQxu7gV09YYgjxIsvkoLktS4on/d5pKy0or9NF8UKNezixRqBcckG/njLR0yMl
HVZqPt+hj+7pRDdyMXluRYH9ktouuZhXVMILnEW+NDsjItjCfv4z0nHjRJZZ2d/U
n9pdgsskYCA1/1zKzQ03xQ0LnJSdOQ4MFtOatmo8cEzMfdJdsEjnFO1uPIeyQj9y
NCv1T6EBk0VVHzqKyFEFdCvw/A6bQ/xHKd51BLT7erntQGpGFGkjen9Yj04rddpO
WDd3sLB97Rg7zz7W8SNPG9g8zNJ/uKTT0+RAzhoh8EddpcUxLpsl27+M1QMmm79B
fBWHt1En0ABYSiYCQuRG5BSmLqnlLHy9Lkx5mLeVcJ82BxVNx99yqgi5y2yK0G31
y0/smuUH/iUCt7m1ZOc+TSU+k6UILXWE/g8Srs4t5qH3NwYuCJthbTvNiTmT0OsI
e9+yhVwhVmpe5d+kf4ZAuYEcW/JUwFmLtJngtS2JsJrQuR4us1llJgW2Evhfh0Mk
a8ivr3GhlJngtN0Ovk1uM1Oc70oQJ7/NolQE/8fF0vaciOpi0oiopkh9eZ052jx2
SFCATr9d0kQUzX2iRFENnPWm7f6kTESs9vPneAqAmd2dXcC14LsWhTGJyEuuea3f
DwmZqwh68KtBw5qKu9AfHUcJzx+EUGIQFNubACNSDrEhmW6QGuGGBWMOVE1R+z2w
g+a9pnNDjQ4Hbny/djvU3xdOx48Cg12qSM+YCnexuF8ier0rYFM5GFjLKJcevHRq
+/RyWa4W4e5xOPsnyJ76Pe5bAGrHBKLnnOH0JS85Opv53zp3IEIjwsM134L5KHmA
16mATd2+jvvM7PJRzOtidI8PJnVHwFBPF1j3vdIja2gORThrrS2ce83PXkFiXg0z
RlWyrNgmMDum3/77hksVhLVE9Lo5N3ETY7kiNfXxvDosb0Favvn0Yh2Ud5VQfBJQ
MGIEZNiScyGsiysRNn4XaJ4F4Nu5Xbm5xUeqersaaUlKIa2Y+5ZAINd+8wW5XxQu
b0Gct8OZJgohEJgrw5Xl0706xvQp5wmp+aY08rlMOlwEzQgLp8Fb24xVd7UUiqqh
vbGDO+8Ibq5BNrwMxSufLLpPhsj3LideBnSJG8pAvE6p9gYo8kKoFdHYWnvov7nO
ToO8q0Sz5t/BtveZmTriSCt/JLMVXeccA1HCdsC5pnqll3uM1sdDHT1LXAu+Snv0
ttE4eVwQC1ntD3WQpO5iJwmjr53LYmOUHbXp/ovnrxyVlZ4AbGmN3qMOhA3UrXkS
UjHWc8SC6/7C9+k+AlkljvgBi6oltQo1fg5+1ouJQzlEmIT9BeoKPvXP13GZHiAv
zLCUIli/h/DhTl2F+gnpPEbltuXztwF5ZZWRFqzHqwi02M4Y245KB6WHeIU24psT
C2l1io18CDxZhnFGD1gGwho96wvaf5LuhZDgh5vCMJNZYccIH1SX5lUPJuTtpYTo
TbtvZy44QC0O3VRRAxMCXVxNM82TK61ab3AUR4vT+tLzmCCQq57CpMxR2xmOWwsJ
nQl8LUBpZR1WUPDm/yCupZ3cp/67sG+BO5yIj1N87C7f2FiEt5xJ7hOCRlkuDCd0
W6rbxXjetlphmI5/Zsc+8UH7qOH2SWzJzdRHbNUxvcPqtSBEMTIlgELLa8iX/EYK
Gxkgon090dsZda+nW66puB0ACj/pdte0VzVxk4IkwzNHQGMTxgWHojgFxO+Fe2My
bYJEOvfgeWibKdkTk3o54xM7JLd9UDn9oS8MsS0LShLpOe3NpWox8wN30Klv+0RY
0O/n2U7aQvhqULdfn+QpNehZTlC21SjBtNaQSGNlzhjfawVnP/HzIm2soCUNJk3r
bWABXk/RFbvVT1ne//5vXuLV8qaAGc8evN3gG6yD2ukRCC0uBf2EqXh3W3Cf4gZW
VDfRvDmcv6e+71SuowNEbc9R8xs/gnJugO4ta24rjfGvatsSfAfunhhyJv88Naj8
9SScooleQS4pCjM5XqBsbUGVXmk5ECqyV33pvJgebmelWWEoaMs5q3gTSDOzHBLH
BfvQqxIf2FDCfJbpmniHjbqyq2rFbm3T4p45V8qG281e32re8FykH0nX1xib9kam
AdtKf7K88M9UajXZ8d/iT6oBFAur6m0A0phtcbRYXMvzbxwZpfJcKxr01GoCH7Xi
d7eZV871jHZxgSHiMNfAaMWt+U7YXArxxYoY7T1Fhwe3gdjnbRvmmtJdZvJG7fZi
RwWwLWPzSMvNonFR0j18RkTcGAk3I8oP0SJo+NY4/yQ2nP9Aljw/g8FqbNohOs+l
tzpNkA/zJ5dSeRtm1pc/Pqleo3H0Hh2ThTMh8zOFqh/EPVXXPji5mz9hFGT7eocd
MEMdrCsQimFhrI0qi2KfTHuEUBbuomGSNPYLiIDhbM/Y5LQqFGzRwhGC8ePKVtfF
NZhL2YxVt//DhO8F0aHSicmkyS6SACEgZhdJqu8+eCEsZ3c4jh1CBwuSffCz5QkJ
pi5IOKLNkfjHAXRZc4BR/Mepzxe3CNuoIpM42ttrNTktU+Q+RcBFS1ekTsYTSEbJ
PpfCW4a7aq5LHBQ2CZkY87i0L5q1Kp3CPTlFGpE84iBGzGhePcteWS0GwKn/mIOl
irlgSipSh4hvxGWR5fMncYpjvJ5A21VzYJiKaO5EJfhXvu2VmkpX9wQSRY7vMiJp
DcqD1e0grcSf/IHpvBkOhFIADtZ2k523efhzmGxIrJFuXgHnEEJ8q4CXkigrDSO8
kgMuJyfIfkzF0P1VN7paEsFnws8RDOe11V8jfKAIi93ozhg6YsI0nSfAti9lPzi6
tzcE/tv1E1PF5SdwCbLpWQtPgW/OL7ucXEf60Uh+C1oZjD+S6scGU/3Yk2Zu/zQx
p7av0dwj6jUBMcQAG2NQau7cQQXR22WHOPeNXkY0+mVrSc74gp/+WyOjjKkSnApA
ttyvJHuiE8y+dHCKxeOGee5PdBuBraYBt2gEJyLGVRhBTFMMRj7dbthJiGw7aP90
85lcqJOVFujmgdM7dsHXmmJHvmsQanaVzZRSnyOh1CoDwEnR5R7ziTfzzXIGcEc5
Z7Eri7OFL0RHJHp9pLw4xtFUoniNWzgSCjYZUv0PGq2ZsQ3nnJlpsCwGjpzWsNlQ
2Xs8nGIDfc+hJJTIONTszEJiu+TpLzA4dPDUniINjqmHU3NZtP4N4XONJGQ64fpD
kLpWBRXqYbKiyFi81znMcjT585lMmbJlRjwQSv+zqiPgHhYl+4zZ4xH9jPt3tHro
k2leYzrXxLyKT/bwKhNCQmVHM/Q8n8Hf53OsB2rOnrJ/DH7jtlQwElT0hZSrRERv
9nQp2XT/sI3pP1TLRWBROXUq2AZZ3h7OZ6KlCe2IJyh75dki3pMLmmHQp8PyS0t9
Ty0PumYp1zWto9tAR9eTkPSxDTu9OLMnP9O+LKhF4EPXPBnGIBhl1HXpGCn2bF0D
1t/Rg5HTwyhkQ6c1wP/uY08t5CdtVv7JWLQciPEooUJIBwDw8HfYAIQhjSKViFcf
kUE6Or6Z1L01smpWoTI4Qeo62O7nnSbLz2SbXnv+NKG1jdqQ6f8TmauL3zlsXUO9
TdZ7yNesw5wBPupgfWl0ZpnCW6Y4cbeNaHSDk8FO3cB9mEHiJrL3vJi+NJlFWQGb
Zl99G8J8Mxec5lwZLszgklTy80/muVDlHG4LsiHK3EngbpgAGiUv5a17/pb5VOmc
M781AiAEAuwlNQ9Ypj60t23tQY1AleIynl3K27rbg4DjpsCan3GLM9sEdjf9MHSy
gRoubdj7cWQsYdULkpT6JMK9yQ8fMOT0XMfzsmPLktvgaKWhQZVzzsr0DGwpB2uv
lhuHTMxNhoYkkCHBs0TuyzzIN4XMD9O43eqhmgYy7ZgKpZF4SjKRhZzY9W/iD8Rw
Zklsy1idYQbOpIqCgFLMMhi8OTqiyqwp4B7rrvbxpajHLZQVV6rkyjBMjHU1wjnw
EZ3n8LgXaUu10Wo8wDbIpTPfu3PXLWCG/8qLy/7+ghYpsjlsLbUIM5owcGRIaMr2
JRDMeX5cJEumJFmtH26YvYaQtsH8pNy+0h2fe8hlgk2HobUxBzhMXKjgPYRhiOF2
hYbzWxLEWDT4NA+0SoDorVr26iQ54JuKhNIZ+ehq79IlVaMWJN283nXPzaWjQbSV
8Ww9+rJa8mriE6/WFKqjozDVM4MjswH2Fm/IE7HRJXHx9TkXDjmwRRjlCkfzQwE+
LHLzMK9Ntj2YXEuL/mU4N0rpRlBx7rZsaPQC1Y4j3XeiRnxDs+KXDrRoaSfmDYTq
xlXuYoh3pn8wmW8/PWhc/vliompa/BNb6OH/r1L2VYhDW1ApoJszEF2qVIA1OVfz
j71Rfsi8riMDnX0PcOX5oLe4KjwI2RuAl5e97okVdHwHMspu6FR4oQhzKwlcU6yj
vsyb5D09Kf5efjIzZ46vlh+2szSOCurZyvvmXv7zX+pn1qQDsHqrJq7GqIT2SCHj
RjBLgwJ7Hdok4SnYI8sS4XMK09rIPo57cEL5tShGbuVMAPoyvqQ0qf0wrrRKMJt/
XUd5H9CX24ECaPV2x6qugHQBNR6BpHWpfrENTq9eqL/rQKaPEA9NOduPYwFl0F1y
6lf+qSfNpBCslIo3QNiY/pQ3ivcYUaMBvKGO6pWz0M/bT5Elc9l5wgdgNdMKSCVf
zTLDQmGY76B078PnGDzM7AWnBpCzmfNfKGPRIETFhiURin6pUoZxeULUEcZAL450
mPn5yRMS4TD551JIAdwfFJPKpJSDsZu71JkDjlBEzSC2MQI6VzP5dyX8iApyJ8Jg
AtqdGuhx80THrtpcDkiXTy9iKdmYFpdRLLcO02Cs1c44CbN+e+9d/HRHj7TM/UVb
bWqOuX1pTsJqNUwmk9YakcfrUC1wzbR0Q2GRX7mfMw7qAb8br8Gikf6x5zEvB78W
2iSgJ29iXIkTwGC2LLxa0qMLMG17V9X81q0T9oqaYjmPiGzgEdNlz6ABHI11BJ0N
lDPk5z8mjJRLLlk8yL1cLXcUdau+JGn1x8uDwTSKT1yPjS+LymL7N0ezN+Yfr97y
K1MoNDtVt7g064WGIoqu2KQ4fV1JMwT3XiNCxOjdxAYlO4F9zB07u5AALDigBauk
QdsFDbt7uuaVUCoard6tosopbdgW+m0v9w0mePEUVNYIWnWzCmKINdc78RmDw03g
BhM/XqBMbAaYFI11bNo70JrbKO+GKfsJI2tM13noIsK1TM8wWWFsTnLVLv1sRKbo
jYTp0e9RKhO21lFXbx748M8wtejKTmT7015xtJ2gw5nlQZh5bsCpvgqa998V4Iv7
EZaIDL1Ff3Tpc2PJD2BgD0uGRH/7Mm85CIv+eldL168kkeJvSWAmREPhpxZHMQnu
QuDWzhRkTlA8cI+vJXeNSoKaz1UxjVWRpyp/yY5PpkYd8cObBcjHnR7zlOOJuxZg
qgPQ2Bub5DHh0kl0FdbwiQJW21OfH3syq4Be2GVtUfQp4deYk2jPfPF+NX/GsC2z
u+fBp4L9a+SB1FXH8hBySHua3bUQa/jowbaWBabAXXOEmWNz51NIZWcTVgz8SSFv
eUzhFLZcdFIbYWItwuNMQ+cIZmWI2Cl1GB/i847P2zdctSYorluqSBIW72lXIPCr
hrsVZsENlSImLTLv9X+1Bo2O5g2UPReAGw5cmpUyIxHFttddAVnHxw7a5MBy7IX8
yBPig0uXMFOMxiPgmp4wqkhZCyEz5fgYGBG8izcL01jsggNTiKEE3d5ItlitLpN1
CFLXwOwELdWjipDMD1e1KkEoFyoYhvBgdGE/Uxm81IL84wVzazrD8o72fd0zYrdk
g8iXCAOVyJC3hfemSUMwEQEqNBvh839NZ8dKGHu/lBPPINW+SPxir9OcLI/PVDMv
LjvUHIyc29vsJfk0HTsalunsUWRNeUisqXLB/oNubMtWZeMt8w+EFSwTetCE4CqL
h1AKK6nkyeQlFaTSiXOgu/+FehA9xeYJP22MPd+YTcXxsJIDcPT9SeyzQqJA10/W
I9MkUbVAXBmqvMm722mPQoXWZ2PPt4nLRwLKqVrkGJlw1xqkwLd+WvH6O3WCnYVy
9QEI4pENhhknRjEa2BKK7NAnAAC2YHRJUAC+gDlfup+gnQacDXBFwBCjr2mmR29A
jT1jDlYwnN8yEvKL9YHpbwjNieh5+YJzkUpE/EMRcrzgEcAPOCSJqn5nq5xi+oBm
qps1wvnEP6s7i6uhkANq7NFh+iearT84pIYLLgN/kzGd4Er+u21dLLLy0PCwI/6Q
fgjrdypkvnzmTOHx05dUBMEMa9G0URmkjoSi81jymDmCRLdfeLApDeT8gxY69naU
72CKg1rGVdpuMACCsjQpfo4SDjfpNVSDkOSQ967wJW4mvMSAff+kdFxjT1kN9e5F
5BVsZHJLRQ/meOcO9AvEa14zDreXQsKckwv7+1/kgBoW6dwZ1pIe+seHwvBiVrAc
F7WPwpEKXrCtzcPqSFFj/MWtwta2IHF90AVecs1B3xriEdVZNKDcVpW3+GMrHc/H
pDULTiqxBRbvR5wcVuLtrF7m4cvZ4jWPHbWZYqS4yiIKRE9pLxkwmaVC1equKhv8
YzkU//Xs3O22j2E+rYjGSm7NX/Oy/Jnb8UM6tMjYDDSqq6QxKDiGJLI8h6nF4jbg
smzG2aVnlcWafEg5z4v7JXbhQewWgo5t22Nx/I9vTL58sYtZmj1Q8ZUI407BhVDH
L2MPIib1Gckw7uCGVGkcbCeb28GA/Ld4RqL9xf0psSFKT+cNDBDA6jhhCI4SxJFK
hGDzrcpE8VuW5wB5qmTdM/nzhhzvkRiVg3z7GXLBn3dbqHtlfGMPq5mFk1GWwFEo
yVO1v9abGwehkcF1VdYNaIaAnloEBr6yIjrUXnK2NBYQdCFjjyd6VAmCCaVvibs5
ikpEzoi2m/Yt+B5L8BxguXL75Lf440xiFigYnSahW9S0a1+pdKYx6H+XQQKfEyNA
EBiLef0DqWD47d5IO+Q/OI+Mxp4YPcAqYYFKl4twuUKpkPcDdHBEVBOPy2tY/f6k
u7MP3VrUKtn5hd26gaHYLdj6mMOQl2ZwbK3IhHZGQRjqCeDllxngFdDPnF58lEdu
w8FmJqqSL5fH87j0j/Rc1y/vmNsRW9/9aVbF8yc/rH7EjxtcrIPcvM4I3sUyYJqX
tpvyEJxOOukWocTVQUBLApHqyFLBnObYM4S1wfjwwbw8gxnSJkb+dYScxr5qtr0d
+F+3oV5Wh88LdrVemk8h/+a09uYzOipWFY9dzG0pnjJLZaFG8hF0UvGcBJKk60AG
rypJNWOynIvQwYEbR7SaqTUu8V8HxeJ8OEDYWHZcUuZncN6Z9PZ3Gi+jOdeh0HXp
/DqZziTevDbfl8wiKuBSi+7KUa2h56iVCgc/zkUWcqnefgOs3t4+jibEtPmLCFQ6
FIMFBhAt5xeU4DhgfhU+ZcVOQc+eKOcqxVK2Bu3uMav0RU1PRmapDKag8kdYEsQ/
GZwSHezNRZYHynmO9/E57tzeBRSUd52LkgugivLahi69rQVHk7SBKugHrTD0lWJL
5l+YN+DEWuj80M1sfr0Ajq37DFzTy2VSNrHR76/8CugNxJVdtAHSk7ygCR6lvjsy
+4vSNxkdhU5utv3o+ITHp1o+xdcBqA6OXT3GPYqBuAzcRLEczeJhrOTmzVnvXaVF
c3uWAuFv3UeHuk+ffx0fTpju50zvNRCkKyrbUSxEzP+YsbrwlOGlAei63N7fWgPf
rStz2CDj6AU9xJnh4fqE70ZH2k2yFLv/0bY+RICzbkMigxb6dlLcav+JvzgG9gx0
cEsEFQioB+G3N7wVNTSwWeA7tsrgNiT2cwlp3tzgKlbeDG5bOsLkd1ZpB+7NqlMs
CI1btletTsdBqewObOLwy2IhBSEfUW4+Hwx/Q5HNt0cQbNZNDLVvL85m8PCfRLL4
FQmBw9tUkuRtDHpf7m1ifTbcowb4He0L37OncQrDu5Y0AkRTkd/wYSTQSVDiB2D6
pdgBD5LPxjUir1dImCQl4unA7Z7WVQ5w++llgA7ul5Qnnh3c2yS5bdAiCcswtE+G
Z117qr45mCRibgGOXCRMgT3T/gxEy3npfteyQaCM/CsgrBSn69r73w45FhqE03V4
ypP6ifXHRgP5VnLiVk6ulEltny5osrHLSDijRjsebCMCTY/ewfkqSHn1ewGUBXpQ
YeKSZubohiTYE3iGL4GiV0KdP7tmKDdg84Osk+3EMdn2JZZQ+4QiqSI7I0x9BC56
eJ3EZhc9FWeDOUhN/vXKUck0v3eywKhwfozyzqD9Pj3hWzv/uEBkvH2W9X1Yrh3M
wDCesvvn6k3YOTY3zoqcudnQNxfp747MF4j37qr03iUYHJOmZ9bGR2lkWUro39Qf
b2DGxAGjNfPdppQWfgzr06dohzRcfm+caHzcyGeqm8yquKk7nZbBmZsDSG47x8Lf
KB1c+/p9jsfu9ULWiwI8RGoM/SEYJSpM5zDHt1NzKviK0NLOjWy5LpFekWzniUj7
5gniy1OxKoAVHi2e45NtMqATQoAQyv0gX8CnxywWIWjmnMICfzmXajVfDZofgtXA
ZD4Ti0WMNsOGHmh4/0u0nUXxUDtFBcOn4qrtL2VU1FESTAClNWaGKFdXLzT7F+3E
xe9oeJW8ug27/vw0bA6IsnzFUzHipxHc8cfVJ6kAgtNjH6N/A3MCd58ggio7Fram
oWPhNfujzLUPSl4DkA6xzcd7vPotyE3CgegO1RbsCnBevE25oW9Mbg3TQ5qd90GF
dCWaTyhr8ekfcQWijdOr6NJX9z0V5/fhALAgMlqeT/ylFs7D2yA7FRW5qzfSdvPA
zmYpAbvQpXcB4PM/1V6g8LB6M13wdTOlf966XA8yUBE0cOucg1nxUJCPDBDOjLQD
59b9XA6dJ/LGKQ3ERESKBJxvuT4G4ad8+LGUu/MTeWOaxGt5zQV2P8t7IU6XNt63
JZoOh0so8hMTTOwFRfWBQmVcRqSrMZQtTxCKGhl17WUgIyU1xwMxsGq4Bdcg79Fh
XLVzG03ltupXvwZvrCgXjf4x16B/rTOKXGvwac044sEZrEY9Jh7ijZ/y/as7AJ2O
IpDrcVqLwFEJs/fzsPYXDP0pIo/you9yuB1scJ9MQ5yUnkwDSsJMusoSMmmwRCtz
Dh0uifRrEeH0OVr4PrmkEBTHSBndWXNfMMkk/VRN3yEUeqbfhbHrMidEX17dhTEG
VKmMuUZlQvnUkTbaihgb5BbFPDNXymCZtjQ0Y9b+SCQDytJ328b9Dp5SbT82Kup4
Lciz8QLZpjzhcyrDjp7VmfIlGJy28cKPN3VCD4RxhG6N9jMKrJcSe4OTxK/XUNxq
RSMvuVKKUOFuZwv7qwyQiUVczntNikcfZlHaSmpPjcqMIp6KQ95VV7ywzAAskEpv
29WS1KhgnQE8dXlDUBQeY8kjO2M/3BgkKnOhwV6iankKV0VWAU4d/sY5L0U7hb8B
eN26aA16b36Bnwa6Ky9Z5aDGo0U1Q17Bwst7C1k/9gJLDtBEPjsH2plAT5Qge2j6
AIYRBvXzoa0zsqvKoGvGNB4kpdzlLZxUPuEGwD+gifY2h0HWU+FLndhF3vZ7DpTr
I62hntdnP+u4XKPgltFD7rTfK2coqWs1lat6ka23C+eeNqCYb8A6vkKcaWpc/80L
W1oGJcFSPEZXy39YVaHgkpPtmsDXUcrieVR7vJQuIXyl5C0K9pqIiaJJ7tk3TwVU
/3VxIgnMS0SA0pHNpLSBDaa+L+/CC8WF/nAtg3jXbQ05MjnZ+iSq+UYG0f0ptsP4
sd06a4tu46fPhE8/TFT2M1NwqlZmTLFzLEvevxaITMujORu4ZKfuXRHHngLkki0y
8Ww3h3qbCdzL89XeID+ILnwctyFN0v50rlaWQiCd8pLVcwKRKqRtI/+fMmAr3HaU
CV+EkewfLBMOYWeZjW8RCbsgBAM8UsKMb2KfsZT2xJVwGUuhANUBltOXAG0lIiAD
Yx9b+gTlUx4aOXzelmJZZ1mHxtC0vkItFZqZ5kMWahFNLCkInWmuVHVE3m6929pO
xuwb16FpkwGsMBSMTgC9XuxXyNdhWWnfcRZDjUcOqPTaDCaHi6vhRICBWET9jcud
5KGFR1ZwqG1o1g/2r5g4uMC7gnJkQW6VCd5Z1ULxtni1Ge86b1+6M6Y3Mblk2XjD
EQBtbgC1EXa881dNuxm5CbloZYb9rLekJlBosFxQRuCrJKZV3JsmsCWFW4hGw3sM
Y8csHjEQzHbbQNNQCR4/Dk6Nd9okr0Seumq2iPFTJJF9DDP6o+/kesnugLEisqVX
3p2ugZVwhamKdlGf3lIzHprCsO4kPjQ18RvEoSFIhoK2Xm4vGzzbxjrD49+Cd/2i
K19LqlmmDKrvfWsQRgB2fgnFtstpeRiX2chiq/xPzmT8Lfw0VFGPg5Fmiz6ziWd+
WD1/MRVpeZg/xlD+ZRI9XPX+GeWJgAl+jEoZ9yWPX/t8FH63V66G+A6SYBx6l4c8
4Hs3/d+fpnI3oQa6XGVPAhGb+S7hgzYO/6okIJnSI9w7S9i5yopcRboaJqVyCIUL
jwrINkFAVBBacGeKSB/tSUXxDjcXtKMSrRBk1ZPKqOz6wUMtHOALcbsIc9GB+uBm
W00FJgTpsIDzOhKByTcnEuf7j8qzqbJJZLSfok9Gu4eXzNA+oBZzwKi4wtVhNm6X
JboeMj1Q6mxrIXQRvVE0VJzL5+XN4OHe4wmEMSsKMqfKOhKPeNm/xQ36aD822E+W
pzYsC80r2w42XDsAarpYR9Op31bphXnw7EWIXiPIGI8euYuE2wGctB+ZOUxXiTKY
dZhh9a1QKij6nT+tFgFMJ/QKBjgfrZ8XAfzyPQ6EkBq3ZM6yCkVHXgXFgj9a6RbD
3arhLRNSzR8O51C+jNBxLphWcFd8BxjLzbyledLphuQwqQYI/IMJNGHS/6wUg20Y
AOJMqB6k3PDmkt9PMaC0Sngkp5r8lNFA0Jz6uvYf+VJjdXTUWqzZrL1Wl1SZ7yjU
6hKeMvM0KBKReZ7BGaMePmilDgcY5by36GlZ0P6pDo7iPjJyFoo72F47ytoBNeO/
nV2NPquWe2+d8HkdfNcC1yL7xW1PUBDTRa1zcSho4KefydifES+zUYrZfcJYL0Xs
hKK0Cju7Ax3BfrlXEqJDIczROwldxZ+W6pNLe4vNUTo/ZMYxR9cPLFsPNsn0fI+G
QEM0DUccyDdl+zTCrfZiqIEIvQAvDkC6Dmw5s8YHVPxpmGfMFRVr9w03vePePfcw
qha7f59YCYwhyJ43+opN170FZLJ2Nz/iQ5MFrPiOeyZg+prWXov1TI0UsKSDrhSz
ieXSSMdf8mXob/rPNKx3IWEX1UC6BuwVkpw0xlRyP3A3L0WR6unMXqCznrDUBqfH
20eLX8t4gN4KjqxL3BgC8+Pzmtap4KxYaI1oYU86udq80OeRUBZjQiNt6FfHaqWx
XrVMDxyPjP7RqzXft01Ro8NGwCXzhMWujGUSjPUYv09KfnPEq2A9plvqDmmMAP3r
u6GyjOLSG8ZEL2pdXOckVElLR9VlGxYyWKMzaJEukSQbQifwIRvfCKI3EN3M9XCR
z3dPqOYhpmrKxwDQ6dN+gS8SwxlGGkVvkh9WNezDUnUhrB9F5XLYu2RZIm6zL47g
k25ya4qPsbYg0S69XR3ygwfTsTM8cjOWIyBbiQIiIitp4PycE8Jdf0Ir/kFsE6WA
caaQWM/gVpoUpAgr3YBDSSRtmf9UNraUSz/IWOV13LRtsAs8VSOF7hjxML/amBDG
sTNJjkpnw4ZV8AhI91dG6/SX7QvG4R1nAYXJlAjneGjK4mWUD53s5gl81XtkA82G
EUINyV7SGX+EfvubDOkoC8h/LKfqMxXJQ6f5jjVlyEyvKE/en7JtaCD0TqRpFR2d
QybmfsE2qSEquUYF1Zu7hadDkhRcXIvp5Lk9oz6iJnX3KqLFD0VIrrSu+TZGo3Fp
4V8XB7J3mIgJW6wGT6MSlDC23HwK8p9yHLfZqZb3HSQZgEuvakGPrhCsOn4Hld4+
WnmrALfLp/xqCdymxlWGzp4XtiU8VwwRuQ8xgapjH2yOwsU2hkVpZ3NIPPC64b/Q
T/Bs0zaBf1dn1vda6f41WBF2Uf6UKjSW3rPk4ycT6wW/yhafpO2WoZ6a4LMmyMKn
wL5ayMuC306pq0yy0uvouWgHC+otKTEqNSPVfnN/AFKu3nghRZb2+82uly4pMQ2a
2OFuyxe62QEET6kCqhqtgW3rVaunHX+4fE5Z2PJ7CukRJf2sA7Bo16J6rdxxILG0
4mzjAQ5gu/Np1vB+QM9LKlV90ieIb/S5Wga8cotyLTmDIevYMX1oflNKDbdsHrlW
04GeRSHQJz7HSablbN3iekqoejYE+Z/vYF3yTb2Xjb4UbCE/4YKzorFLG1J955K7
BZ4MiLB4snGDkkjIkG7G2xJzDAmGKf4XDbnzAJW1oyqaiKQ6Wq9LsguR5liN1bZn
MSITjtksO26cLxg+93+hBgRHuJOZVUGKZTA8ZwQEztOQdm0TGS+2zyD5Dy1pC1vI
wb72CqjC6WPSs+AmCvsC2CKB4DmCEf1RUDUhXTvYUpwFWgjcN5MI9T0ctt7lGuku
3N8XpeDDrhVDwSUCEAJNyDfeq1GV81gR3UYUduvD7cWuo4gGGqmdLBaZvmStAlOe
Zypr19Nz4pBF4hI3TV5FFSJaYmtQ/XwCLOPLpnDiq4dqMj6Q/fyiN3yztzJT2Hfc
oVr1yvi6niqjLPq52XXb21HgDV5ee1DUPAj6Uw4onm3wC5SlHjb6/SXsMfMvQxqC
uAKH96SyT4/9xo/nHVnS/Bijap5J2WThrBYpJ5jIe8jhRQukFZU2P1y66/iScX2b
IIhhSNUVYJvnsRMTi3/XisuXDYalcseKEkwc7Gnms325BW7/t6Di8sPvOmM4laHk
FMKxLr+xvqYrocKQ9k+UU9H0o1mZNCPksWYcM7QyvHxj10o/wJMwefJdPnjVf1xC
e2U0SscJNRdTmviFFL0ksNpS5rIEzDx9pPybpFR4HFeluGkNle40WUGDx72ky3/U
osKYIqHZZB1xL85KUFoiME/RPkXyBBuwsc07ogzTbXwJdwi7uVXsHVrXphZHiufg
5SU5bS2Lhv07vMrGfoBNdO841BNxmIzXfm4DHRcvwPOlXD6Iay5MfN6f7o/GqHsI
lGtdfrgWIInxLmRhK+SqwaKj/zhuOdA4OA5qZNXsBUXVtjGeSJPZ9ghgIzPTat80
QkALu5CwY7d+2LNFvbJ6yCbVGpJrekmVGu+olNdyl09i5Jqo8PS3LdvRedeKCvhc
wtqzYZqzJQBJluFteNUcJCNhxpZguC9mklelA5WsXdFMjAshQ6GA1qH3pB8afDLO
2Xk6Wq8Gve1Cj/L1Agtzdby8pCPkmvbCTwE+fiuiM9Y13UiQMfDzkTJ3bDNzJoaW
6DlHDXbwaThY9KoxHtY5JO+dUs6YmSZBa2HwPJd80FFT8SG5+DKpTSC2aJ711yqH
5fApmbJPmoHoAWVUwv0sj6LrulAigejLEEuB6fLjt5WxXjJHp3HSBDg3Ox9c23UC
1BusiWJN3JQTCa3nj7qOsg6Q7vivO0ZYMTFKxKt1zpTSJ2U4c4EBHrqn9XcvuEUC
bLBGrfia6rk3feHH7gkMatftV6itNLTsbWpfWsK2qGJw88AkSAAYVMzQnOrtjcYX
jpxdmkueIZj/bXj43jrnTZvN425GF+5H2FXoJQ9Z/TRg+SwdlImgyYZuLy/B0juO
k5nSyuY/Jg/EdcRRlTGQs7KgXngBwxhSFNqqu4xe9n07BehcGTQfhvyfBHizL+bX
ckBFETg5a+0wtKx/ZwD0dBIWTfH8ZnafosyARpJPhYyqUdvTlX4gm5lw0EuZXPHz
CSM8hWztq+MTK2F/2jTXL94LHAZqTGu6HD8BAvkYDFUn6b2ah0M2fWF8BXBocR2O
IXjjaz62YwSc8XmyRA08iSU0YvS4tTt6JjonZtxozsnIPt4tlrbimk+kE6Qs9FN2
RIRVaX2JHgWetOH4D9qis3oE+hjmSOA6MQ+YtXHghql5J5s7Y7G+20CJ/iAhedxY
vdyJE795I4GxNYF2iZMsMkaMTGtwm73EMryzUM5ypPXz+L9TP6m3u9YkHtZjb4Gz
jGOK3TAcx58TPEtbdgzn9zR5uopOt7cNfWNSTN83HDAdVS+hYobbLBDMK27GxXko
A0/Ltl/sWmEBloS+ao+n+VrgsAryt8RbCZtZpYDW9tsmqKDFWNI56I0rdGrw8llK
dQT8z/N3LfI9znL2lb1hxROIj/9bm7VGF22uXfz/tpuZGOC2nHG/X84VhtvHyB1C
nlQ5rrbTG7OKHjr99TisoVs5urKsjz399X50VOB+yE1sSR6NtvGMUqbtgiumpBkl
EkK1XvFRoJS0R1ZynwR9udfuABCVm2+ijIKs/cS9SIZcu4srrHYdyPckav2XaUZK
ZwszqAVsevG+504nSRJQrEZI6CzuzAbGh2zLzeHjklbijqW4gJeITLDtS/btp9pp
M2N/WwsY8UgwiHGdRhYzT75z8AzyYuK9dQLT5f3L3C/vxsIMzGnReJgDBdTORmJ3
S4noTCyHkEVPiVWeWNPuCPQEfKScAZuxZ00IV6QXJMxr6O6hMPBuNTA1VOfqROYj
r6IDkU/BATEuUcuJmoBfvwyVB0llps9Wj2ycLM3S7XKgLDkVKXVyijHCd/lai9yn
fhSf3TWYr8kfULH/i2byyUyBPr+MH9h7VcVDrIOJhpbqG0ivMreI2bBWV2nA+h6Y
JsTOnu71Psf+dOLxHzsx0fi/hNbGF3Lwk4WaT2DjmqIhWW+ZuL9T2T5Z1LTjOf6f
I3TU2/HY1tk2VkoLzFcJenO3gqG/ezCSGZlcsDKDgYtO3Pw0+/ae62PCyzGq6Nva
y2GkaHvhGmU2xVbYinuUqA0UweKZK3tDmZaeGEh9SQDaFtiN20OPOY5RdpGIFPe1
7pMuxX34rm8lD/ad/7aUvaW6yUc2azSVmLza3gFKaCWykjhRAs37ZkiQcZrf6gzC
OH1JUP09F1A2E1AiKxPFIXhibhORChty49BQwRZp7cAObefHge1InMwInTXvZ+I7
dsN2sUDwMUoulPo2gDm31ZZ30QnZuZ/nHKg7PbUZ36LsXRBbav0dtn+HVcJJnvsd
jhkYlu4uL6kpu9bKo2yfpE3QE92DAep8XepxJOdrRLbD8cJyPfS7KbKWzJsMVw0n
DBqthVl3UQi4E+C2oehVg+vBKEw28rxP2w098Cb1oIfEJZ4lcw/sumQMov6iztNx
xUXjhymNyovfdopTb/KOeHHxH5pSdhT0NQNf+jU6f/J6zCAecGwkfhX048Q+unW3
KGL4G08K1LmaDVEcnBZcCL9WHscjtfc5jVkxfD5jvZkb+dKZDaDgzOFxQnfTVQXH
dFtKwn3LmAGjX8iy60GTcBGlMEEeCGQ1BoGpGqQ9oUq3Cpj44oZLx4dnQdfO25gq
CjVjUBkIlfMvSw7AXAMKtReEQqMZdsYrNeYEBLTdYTAehk2XJBpQZym5cdvdn3Bu
QiV+MeclTQW1RNyub+QvLpEIOZNgQnDwkkp8sZdnAV5dynXAYnXePY0MT3zbq5YD
poUT2IRpUMiOGz/6aeH4IMlemG63qxeVypySUXVYEuJg2GPXVhQjJuOx9g12wbtT
JcrLujk4dWp63W+HVhTHffH9cIlBbrG8w5rnuyIE0+9le9fQBQ9SkqAadHikzhHz
eZjswYcoMySe8UJ5jCAlOeCY1ynK2s+d1usWBgxUP8FC/bnqOPM/9efbBExT/Bmm
rzSnCPvM+bwoEzEPcDtgwrpQoZypnRTWB2fsiYcPJU4gJa54c97D9esaByCpaspp
uTqCV23EgX20yZzPo+68xUFpWPLsb27vx9e0B148c/geP8+qzVbAzckxNoI2snTV
zI1teJN7FV0dp095SojtnMVK7bxgQgBfOf07bOYP+n6wwDxGgb4a7wRnGmV4N7JR
OMNPeqKZEyTptOywFV1btRWJkhd/SiAcr+tvPsY9yf3NSQBuLkvSchcRgszvXEAw
HUqzHC7u5/YV+C5k+wQDN6z18FUGq+ZnelR5pVi1AUroH63wHbkfX5+/6Ic4i1eJ
3mbLvHBObHkglC6WIO+1qd3Gsb68Jt4prNTOadVX+ASw9j8JPrn+hXVOhRsyeG+1
BT/ZAyu3qw7RopJhBUVcIqW5YwcspokNmugjiW/+naVRroS80zWi5JpY4FfkGOod
qhcmDzeXFpxlXLKy9Z9TuZQ/RaN/mAJN9S6EFsSFtYUQy1Kl6bGivWJemQmnxWc1
xhxaUELTz4aGRDRZSsS5nWjPqtVvlgYj08BA2KUqJd6OfWONwQ0BA3nRDZwHizDL
8ysJhC/1zsrS2ZQSVzCln3Td75YkjHG3LbSJ0aFM9PquLQj+qLUJAX7/P9VlXZHL
J+kJV6ZFdRy3/qqp9Dvz/DafutUa0+UQ63sPzZgJpPGYgTBcyo+RrsvOwNt0GiPw
ql0xTZvsL6ZGiNuUONErUYAHpOcU1wv5r+wbcnNaHyJrc6WoH0f0tEW8gXlBAh40
VzHqIpaNYm4pFvOwdY8TN+hQh3DXpnKcxGggs2ai0IPDwkW0oEB0X9vcNXYkKgng
3+5oP5/9oU4QFPVj6CW5Ou/UZAy0CKEqGJWgwu6+ZXxuP43dwX/Nvwap6yy8+KQs
gCrIRnOHQcf+HrNCaYFhD5X9ZoEA1cGFl7JQFtnznU6STuloGCv7opRI/WJ71JZy
vQq/1AC6e2ipq3V7H998pg/H7BXV6fzHZ6M+oRciCAdiDSjFRlOM4c/aywRwFTxy
ALUVtSfwnCivxAPIsD6xL0065ZOwNhEh5yTLbO8PRG6s0ZOGZZafAneva/ICXG1Y
1mRSShaQuTqOYwUhOHNCGI604oV6g110TUVJUyJ641w2cPH9qpG1uPQFOqn2r/G1
ZQFPJ5pk3607JcF49XNU02IleDV6dDLp2HNEE4QneSrdfzIkyYu6ekWOzcFbe+xi
Lpka3o3b+B1S90LePPXb0BHfyvf3yU/SBk3AVg4vTXq1t15hSVvSAdBt5in8dvTM
5Sv5pTvWOxTwdrmioa8MmfAnn8W7EewuVDFVqnHjh6dHeNeXOv6Lhn79jSchD5nU
PYLXREGVGevCxlAMGrqU2yvgwvgbf4BC4X9f1x8d89E2NpLt/yydhp/VSUmcLisB
LD3fel2ycO+hFJNhihbzO2cIPTedlycLr7i20XLo270Lf5Hm/7hdF1t4EO2tzxU4
T2LP0urUk0IaTxDqgOMs5BeXKoPt/JLXl6AiTIfRvFstfmzAcXBtIBEF+2tSesHr
GwEOIHey67PolgFk9kzNVJAI/OsHQolEVbtribD4G96MbdhUSwQ4sOujtX9OQUau
hiIrK0BGX5fZPgQkKTnx9cYqxOhi/jo7fcr+NNaF2x6dua8iR+hxk5UJhUlZ7Non
t7Ca57RIO7P4Lpg0wbK240831B6whnpTeOaYMcO18doJJsohtV05kgAeCA2Dt7PC
TkHP1y9eiuU26oAj3DsXR0uO3R5K4nlRDCqbGXAhIgd+G5KzYbSj00oBrpkJMRbz
ECy9PR6Dda7iUhC8fbCZQzai/CcDrgCCHXh9u54ahOXVJzUhMxQf+IzrVFAQOtyz
BDwAJbSmRqyBTmjrGJCLHGTRkdBVcRdMhnHriZquokthqdPiHywAtC/j9hNt3pJp
ZG8QHSO0TnKfITabUAxH9O+Nt4Nwdv3zb4W0H2zFfwN7Q9NFP5VbPvauvPu5R0Vy
05L6OG/FL7gs9tRq/5oUbd4pb02i50IRk4OVG5mDn5O0RROelFwxKeAb4bk1gYC6
93n2lElD4B61O1PQ6ppdg0/pfQuG4oUnWWfmVDWKrKRRzLJ043JUrDHnoA/1PcZC
Oe41MtG5V6haxi+LOZoSVrDZsoYQQLp69ZWvtGIwL3wACnnMnNYftxArZUbd9O9v
M22VnGo98vNJsdDGvG3RofcgB3Bj41loT2yEMZeotpiB8vtSCow50f0ZMnzAdadJ
GUGjh0SQCGlhHQUfzwkcBGaCw9/tZXeWIqZAOQdx9lpNhfH+fahGU4vYR5HfMjg4
EDnCx2q3nDut3QFwTtyh3pPPCD54h3/Q5PuxwgNEA1B8E05/TUOOuWyB4nq7KRJK
u4WNe/xXvCHX6NVHhG1s4nlkpw7a6cZNfyIf17XQjC7JTCE+ozeQm4BbRJZNeww5
bvdGRKJlK8+g8K7NDoqj1E+bWaqDBuaon2ES7oe4qv9BfsLn49Zau9HQKNjyi+BX
o7zQ090pp+rLXTE0xjZeqjnGEsZmiGjI9OZomraQkn/Fq7MtVFE5ZcbN9prd9aeT
5CO/GuAZdXCEnSjXj0yacplIHl2anIh1BoTIZ0M2ciHM8R5K/+scovO2kW7uTU4J
sdJ2+BTCoEM6irJ1e9kMASQSK1+//WTvNRJT55Ggc66bX5EoFYKk+VIV0eMn48MB
5bitvY86uddnn50eZXb4/5A8KWmAhOEZajo+etzMdpBN+3ovUdYncM/nOgRjWOYq
CcoONy6FQZjVqq5f/vXzx/aRwt2WIcDih8tgH+txmYk7zB/mUfv14eAYr6OziCAV
9X4s8TfUKfn1urAeHw/owEsyeOJq3ZHDLp3c9VMzd+Mjw1GK0TBvUTIQIqyzJWan
koeOX+9FLCgd1p/AcJD7WxxO+Wi3eAglGzYRQRdq1TnJZVoTwLSEaT7a6xSo0Y/L
blZzZW4/flbyms2jv2DuVvxxA8ExBnLlsUuDGPMVxUcvwYPo3VGCSM4kethOE2jV
r4y7UorHAfasL0cnOkpLSDk6KbY1pHE4nf/Lk5PE71YAuZFLfVwQsTole7UXyTqo
jUlEbIoAza6gA26OY5arHu0rY8dPpub07orC5wzIFPXqW4wNTKwn8z33SLMgdr9G
jKV3uCUIB7Oe5pvkMZOOUkfjPJzKFpMS5/YbbZG/lQuHWv4zzbU8Ywxx/TEQOXFx
0Hoe5wRTad8jC4guUrVatk8n6KPBPICBg9d1hjLQLWYEKjCoqeyZfM8hdZWJGDQ/
adeRQA4ghv8h9UwmcnoIgOIXxGOawBVBziw1B7yNb4sNcHxXkEDjY7X6/6QcaoKN
071NVWWbny1mJWnjfe+gPpCt0yzcRbxk80HDoWH2uHN+Fr9SkQxBDq/zZfNyz0f0
QXDPUe7IhRCSGdNq8ms1VzQLbAyBcoDeaYMCvl8BkDtFmxUCqji3P9FLv7VyMnd/
l4ALWF0okNruBrvu8JFQru1I+b06auC49b6BhPIrEZPRLBDVBPPWApPlldRgQjdC
jU6PzrJUiqyZ2pLJQ2qAoeHuKssavqOPrMpdS6IOJO3AFRHODmLaDBEAi8MiFg5e
LY+/Hq3s2buu5S8Y2KKKjjDCHdSOI0bZiJCSFdxgTOoowjD91flpBvJzRei5OuMH
l7LcYZwavLP3QuSOAWoeO8G8fvokI+s4WXIYcOVmergxu3uF7c3gP4gHwXEbpbBj
HEgwNQ6lbo/PJXbddCmHJ6ArqkfRVvqFzsYGOFfS4/bm0OfWfN5IcUKqjNzaPkY2
/iJ+y+LfIWjSvqNecWF8Mqf2Mh1quqbIitcVUIwiPZL9FgGKs3YYfdnlA+8V1073
Wd5WoXTD63B5KdxrUPpWUHVb+FxAM5LvaMLIGrjp1TLFnta4xx/zENIK5sUnmSpS
t7+sBhSxrjUM3REmQr+slVUmTVcmZzhV/t3negeZT2tn7N6pyvYmATqmFvI0IBTW
2MIFfaXIMqgTCx7VoVdt8pi+qhKsj1EMX2ERKOeM7YP4+42f8xgsniBnhf41+Xxn
v1kKQg+Pzjstyowt87LWStag+D42+9IxnLuNsbsLPWibDQ5Z8ucHrHxSZNzD2xbi
xiXqHygxK5dzBcLb0BtU+LNvBXU3LlhsZbqRzU/CK6a/FLWf445h0MQMQL2pBz9w
Hc4C8uzjnfvtAoSDPicByzxxsX9PzA54pXRD+dDlMrZZ7G5RnNbiPHRBHvN9Wl52
fJ3Tua8gywsQv77SZdQA4Et1IBaKdnE1/FU6SCHZRoaj7wyORK/bb4MUy0oL0S3V
TnLBe74ZLVaSueWAa024qH4kTDJ2KAmmaPyFQsVztxZosAlcLGxmFByDo+oQOwwW
IVCr70lpJxOnr0wvv7mMCI8CA5BRy5dL7MIm+DL6iWlgXc1ubc65cGxR4uNbcXak
gH7n5t8JbUtrnlOGCmnD8Jof3oXyGFCTwZbfnb5S18gzMFRr0krAa5dyCaI6pX3C
s6RDyL2v7NhSrFpbcqA5+Obyohg9azM/XoGkuPJQmjyw5GFd6F5dtteuIeu77Yu3
wT1SaeTpZNOzMvGFfXlUZBdK27YbzkpV8vWJgAH4FgjxkGW3kWDqTO2xQYyqcz69
NAFZhpz3G/x4P1se71Kn5nUm569YbJITraBBAr/3Jv9Q/pEz+9Kx3gTD6JDemFAI
qBVFOCxDkpUul8L/SDbXfUb1v/aaxybJxeiVkwsQOIXr5a09O06cW2REbJhKn66k
ROHP6YLRyXzPUCU/YO0TougpFLnhyEu8wLBZ45u7+KKqFOxwp/UccCa+R1xkxwHt
lZ6y6rhdRvdeKy2kKQI3SFcLmbtW8sETxWPOtiqzvomH609D5FO174fHYrCaiW1L
1fb5mkAjsHOVayOoL+VKF0giGrLW2sJr3vw7A6I0gxjaRxqtMdG0LJrgh6rYPOha
nNO2Yq2NbkyV/i+n/HaT2wlK3yQ4I3VIZJ8tY6m3v+veLTN70jyNYOk4803VCFtI
Y8RB/HdJOmdpx2nPzReyJrz0n+2n0wIdbPmgGUbDMbe9FlmEsjkxgZ4TkSkVNmCK
1ehh9p2ZkJCTwb8udUOg24uP9d7WV8SLpG/ZUrzK2TXa1vQrcJUkm2I9eVEsuPQA
sSFB1Xi+1ETiThmxWSWdyC2q+EzNMzyUB+C6XXtLlVjF9Zg+WHP170+W2zHbx0Bd
CIVyJv4qOi4ARPBbrpCyZPqbyd7IsxgtpU8JXSzHBNpmUADzFZb8NKw5Kbz7h2Nn
iIq5VjZ76fIs0SwoVmYE8Xo8cR6Izs+WvrWweX6HkZKN2ytF1I7kD5kaeSjXg4iu
GJ4ngNigOy7Z7cT6ZjO6llRM/g9SGGEPfKuBsEsbjNV4uiZukYUwR6YQESMlsPcA
WVWjc6dEi8KE6MrMbql0bGpvAJzeufUgsm2WU2KdS7o9sCqbsYm+o8rLk3VDWPCT
FNGeQ/fwZlvvRedEcm/ZPNtfDR89WS4EWehX9B1+9nsmumtzyLOMtBHk4786PrNl
QrInQ7o2GPGt89OId1Yj44aoxHOse4CC61fYYfiRLP3QMqSrk613Ak5nZl+H1LPj
S9VLSB3SI0aPRsYVPNzLB7uvBY9d1fDd/DLnw7ECasm6R09sw8Ij+0DXAC+vAtdZ
z9o2K0m36tiOooFt9W1BEWlGZEKDZCvNzKiTkflVtvGSRuYiUESmENZsIqwC1zEi
btY9IqKfxPFZc51CmNR2DAEkbcw+GCRZLclq023Ieb5zSuNDVhIHq7UTdOR7uDsB
fnfDzTpeWa13Wl8x9OBUWIRc/sbri7PRQ8Q9dFvx7K1vINdNRsj0Ma1yQ4zCc9+O
5TgoWUB0DfkW/gdgtjVDC2dSGtrMtKdNdqAQeYC3WvmWewQJBiChfgybefIyDN/j
SvOADeZ5TcNixz4EJIn/wn8A5YQY1kxT+fEvcEf4YFXsNfUiY2xW0tH2bEpKCAp4
v+FTO94TJ4GL9B7wP1+K+1ZlFhavKA+PzvtGfqN+IVSiEUxVioVWsv9IaQjp0P9I
6baJxD/CGNPkBN2EnXOJwNN4cGeqnImTDRIaTnYG1P8Nr7DpbH1b4/EbMFUI/xnu
B3jzLA4tesf2NVMFz2WOP1yB91krT52nIyFFpKJuFUOcbkvzN2PWYsSSzz+RQJpK
O69TKdzBXA8yD79loakj+Yjo0Ewie/8+8z6AUEaaFYA/AFXmDPmUTNHsO5YVa/7f
jPZOyFFH7loyGc9xY2OAApgoip6Puq6lmoXIKmHRN08zRkjWwMmoMLQtzxdGen2u
alGgYxsJmLfOC36TjLLX3wBWlX9MFZiT9Tny3oB3c+wBSdPktIGkEhcWdz38XokH
1T3moeCHPp7p0y4WFK93ABMFIxyjvokXx+8Qj94li93EuQebaZjRliFwuWlFOFNt
+aburOL/xHLIpmG2uV5s4PSWd1EN2DmKEdlrVg0/EEADZWju5IktKX5cVrhQF1Ly
rEN99/63k3Fn2MS1j7O62uJ31FbBpcSOs2xmNS7ihSN43gFKvOoaFtVkpeAFMmHj
3EEwHvX4yJ0dpe2LG8bqBme8fachpW9yygvPAQt4zqemTRJH/dT/G5eQGX2PNRa7
/QVr8GO58VD9uMFwY3HYxZ6R5urYnCv96+cAnyG2WaAjdAXM+tT+wBj6iF3EiBxC
Jonbs50MyfoRYNpJYNuJ/mGDIGI7xKf1fQ1/CSAzOrbzuGSmeP7lkcB1snVPnglv
AB4YcajqU4zgcEuqi4vA4ie1pf+2bClQIffaAHVi/ivVr5kViVGnsEUYRz0MZoZ4
g1Sbk88uQhtrkDRiagvZGEYsXP9vL+3gsChhTOJY6rIpR6ijUg/9JjLa+6cckubE
9XDWlbcVhFhvlDApaMcuIWdoNAOnyD7lBDw/9qGEe++aFFE35cPVVztwJB/jJzg3
ASiu5ljN4kvQwoYCcM17ABaeDRRIaS+hLReYcaf5b+KzA0kyn1Wbsk6Ei+W72ZT2
DrC8NOVKmCltE0+d62Pa8xsnjwQXaXUMlvym7zrsPbuNsThXTOjJ+/GqcdXl30iH
lwS+BCBfWHORFaYN+LIl/VaOvZ0PpqYQL3RWLgYSz9YuZZiw0U4kZXAueGZ6TLEb
jn1Qu+KcygqhOGkMr1/kp99Vjq90WWUIzFgU3+ncefJfrunz+kuFMADV5xLbq/sv
3CTmBB/er9AHt0lnt25YFTRxA0Q5WboShRk/UBJsiyso62t1U6lbSSi4I7FKa5SO
k+pHM5y1baA3hnNK54SKaXIkeUqjZgAsVmPeAJajDCVD600ZlPR7XUZ9APfbc/vK
SssRF6znB5mnfEpDKZzMx3A35K51jw4P18i+nNiRi4QV7q6kLaFNmJfjaAPvdzX1
d3wqSr2VcmlJ1r+UIp2siA1MlWLXEtWxs71zKvKL2G+sZWxEg11Fxr0J3cVpDllK
WzLum+laJniuilklX20wkOsR7r1qUct7DO9nQqXKee6MLybfk+KcTzbqLuNFWA0C
qIRu3evA2Hh6Gy8SjX4Nh1nt69lmDq/pFvmWDjOemFuhDcfUU0HLqdDzfsAMvSRB
R04XRiYsOvKlj5kTLv+yaTapay0umve6JHzFUZ18QOylxMv2CvWNN/oSnifMKHhy
0Mscvg8lOUChJjmKZz4O58YBzR8q43oc/C3kGAdPmRHUAH5BvO4acBODVZbQ+Zgt
zws0sqHDwsDJt0G+KBdc/Wvdnba6oEOgk3yuUkCsJxc+Acu4GoXy/dtOz9H2y7R1
KPFZJ6gKPPsMLMa2RICfiP0IuVP2HhlQguVp7zIT1OhB7xBeQfhoBzKx7fW7dWue
wwHHByQYU1Fe7SWBIwJxQB2tytMsrz4c1ceVn9eY4l+ec64qLSkCU4WJpKghCKUU
WtQW5N67m0VqKNTo1kySkddS7CQHG0cTo1bB0oZqlNXR7MMe2cWHP1IUiNogokBW
ssxMxw/wx0SEMV5zkEC9sQFUkNO1P1Xh6AuwTApQfg8IeP4K03YhJ28WUC6WMRb3
JpPyGdfHZBjtvOyDUBqiwyO5pD4TsS+XlZVlvTHh7q2IurqPT08v0Hm5opHSmolQ
V789+KbIfqfxbitOFEN6ww0HuqxSXrAZEA2g+8VMYqEF62u95kCRNKyMGtkN+7rg
i9niMqtHLQtDk6xj3a7lBgqp7m6T+JA33A0Nii6xLoTi3IsNDxqiOBK9VpJId1r3
n7IxR8BTf2y3Ow0CdBC/18uHv1dqBwyh43cP7+IJCS7wfNXpUF+EJ89MEuxljpad
4taQG8iLjjbhWXwhD+9WHMgjXyyoMZOiWIGelteWh9fMpoWfshYyNdeH5hIFNoKr
qz9Hrg5JoH0oL4swmBTWhtTaq0HmkocZPH6xB1979DGIS7lrsR1XsIZNyEY7/afU
CpQKk1dL1CqnyngP8ELBi7uv3KXBkC1MCrinfDhx1Cw3/Lt8k3zFCicaD9cYxZW4
W2c33XUHddxZKli76DHC5bGGKT4OncXt93bXYQXExOm2iOnL6Eq0AJQzSjAzGJm+
OWeuntplda+1NNhVcykHgf7JYlAzSlFXm78thEPP8ifP7fu7pxpmLoZtkhwGoBD5
9wSrUOEEKIEH4+SLpIWcwv/8pXCm2j7jJ5+u47DLWeQxbMB2BopO9Gmh743bAAvZ
O8IB5h7DNy0vh3vNsTYs9pyLRdyxF/55uMRhrmIeFh8TVm2VezSdyfiIfwZPyP5l
hVxk0SUpNdwZp5PztQRTUG9V1u/pZ9z8repkBpUQRCwy7TJO9nq05R+IN+GhRJbI
qBIkUPSxF7zpUIpL1gcXaYX28d7Q1KN3Ntn91OMbSW7svKDWadukO0Pfor6ABNu9
v3xVaw+G0mEry+YWjEcqwSYF2H15ziEYO6RsJUSQnzMXyfuwEPBxfneNOzw2Q62Y
cqYDVfzi+HKbXGGJ3w9Nce1tEMyTvJ9566OymVKmHKWQo+kZmSFCKYjdOIFC9vuC
XKP4e9LY+4sXIamgzt/fDEkhTG1dyssmXa59vb9DOBo7vtDUVuqR6sFUyW+uwYKL
Yt+sGRGSZgSHEk7FQJr02qezv88gw5NdOFk5bHQKj+aEmz8Uiv/A5jiNWVU80BaD
lxcJc1ihgJ9wT6qsAO5FS+5kiDE/Wde9ewr9gePqOwKMUpy7es0Etz0mIF0/Nxbh
ku3XClQHjPlSN7boczOLSvumSzk5MJGvLvE/FcSy3GKZYnEY5jpl33jEFXrMbvMK
SX+y1KTODBSjbwuiS6xLfqd4ghv7s6Ju/PaN4Hgaxm+2jFVwRxvBt5VXDiyR2Lah
omcknWf/tfAUlYLBxeI5qvtgOJ0Ku5AOMYInB66gXMOJvFx+ZDvU9P2O2ZFnKpbr
AwarL3sxhQKkZtiA5H7nF3M9wagL+oG8W2/IuJR1SHi/OaUgR6rUBHSiynOB8iHK
rjFUzj3bAnGHvBB6Uig0kM1J1kfjMkcZ2/SRAl2FoFgzXaxmOodywKK9b546gjo8
dYoBGMhVwIDla8WHFDdjJT26qj8CyAAM6XsIhwEbNaTugjQ9L9t2n6VLXK0P7gxr
wRyxjWHfvA9Ym1gqtPDvu8BM6XSziaX4mFnnJx+7Hzg3cuxsmGFD1rXwaan24RgZ
Vjv7/rDQOPjlZdpZriefheKpjA8wCqGaK7ynW2cE6B/2vk1RnyCzNq1MiNj3u7p/
wEYO1p4veF9Z6xxBpJGmjvclrWuEMHAYAgXp6wnl5Pc9Of29Ywn6dreOiAgnV3VH
x2p8R29ejz9V667gAngBiYZ+UGrVXbzIjpBurDnx5neukdhbjPp8Hmu/4Rku4VcZ
5FU2pDtvuZZZySqBLO4H4fX6XxvfgA4tr5hn26lr11ksDN2hjzAcmEDPx8HBL0fZ
osdL7cEcfDAUlZWcmVZAYcOBxDf7JW1clc/2uwhZ7d3bQm5UkFRLsu4QQOf5P4jR
vn6bsP1BoBFd5je6lOLvX0/UmMVtoM+FmnsE9PIG9MV8WrEKqQxb6BXY5NyJfOE9
PS3fA7WKamhvBGeE7OnkJT2K24TXm5F8OCNEMt3jJGSP9ARNw3p9U1Mvaz2ZOoqH
yCoNbfCxwnCwcAwTn2ZWKuEZ5YYMg45P/cUh2Xnr3je713HvUhhicKnc5IIqt54U
5+ZQGYJeOEFcY+f9AjFD9+scL7WFF4uvOg5JZFBw8ayqhQX9Jwokje8GPGWqmB1+
Pr8l0cXikPZLPjGe5JCRLqkEtRV1BiGmpG6xEZ/iP4Ht9lGHMN0tEUDs5zctVHcN
lSlfKTRkzF2sHbnHPXbtE2eqx0lJkCZn2OGpreq+n6rCfJctwVIIwfBaGBq4sCU5
a2WFkrwAAXP9IrO3+RKWKjZjviAWVc2o5TvVJH6ATn5KKuMZxd6XtpiKaZQe3prz
WlJUkjizG6ZGzTRXvQjpxwn9CibcA5r+G0wsL5yMyAmYfZJ0qq7zwq0rigLLqH17
GQuJOS3B9lUJQ3vLIhMe5OqK+dviy3xVHwdw/VWpt17zJLnlXZ6++m613d3PMjzk
Dch4amfm8YUxlRBnGMlvNOoiJ6a+CbFR/BfqZDc37BjmkWkzgsJZ/N5SLc+9HlN2
NeM3wIOTvFV+1/KdWzLzwsOLFYwImKDkrfFFqhpCltU07tvSdH/PFxbpKEVhc/9J
rUmrKfVR6sT5ErOaZQHpUjYsH56twQD7/RNZS43caNDG84jpXVO/j4P2WcJENIUw
rR32XtH/ggsz47reLl+hoVAieS4qvQanN1wGxdGemWvb2NvVz4LwKz489+PTobzp
6e7k+ozPUwFjJ2p0ZlwM5K8SYUd+ULLEIATvHt130oC2n06o8ckVagNeWPPY2MnD
Zr0vPsrNNB7GqoJQ8ocJy8/vsk7+KUy4IEXTSqRc/r5JAbeV1IQeGoHEjCx8INoH
GAiMsiTjc3GIVUdWMK4+/DmbabNGo7X4+MhxGkJ7HA97vyDUYAaNeeWg8zx39v0p
u4gB8TO2ackMW4aUjE1S06Lf1PzyHlHhyYfg3B8JNOx+7juRkQdIvpY/Dz+OxGR3
scisRChp2qLO0yKrky3wMVn7CuMRXvcGOuYlJvuivc4zAYdZjOsTvWwsq9GQcNfR
rzOuuFr9Z1A6p91l5hF3Xobh8YmC/nxBUd8uWrqM5ihThMyAGIZqNcT5sO7tQ7J3
kyRlusJJVivKCEXO0bNztEbkAkHNTQGwnqT4cxRK3GIX8aMI2kTiErQTmvp+9ptS
OjbAEIp46YTZ5qg9ZNCUY0skKxupRkoZ7+p6NtRJOGVnMP7q5+nBukzd15As79Id
2q4REo1qNN8eWYHxiC17gfqIyME+CSlzbPMS/x5foohCkTzO6U3KqdU2FyzjXitG
xKjMkunaZD7gWymZhaQfaTvUqEucdHiUZCgdRuRPkcpq1Bko/AtOu6J64cqvakxM
18qqx/OKTW95McDJxPZCCWkJgohPFv4dUHw5NtOOlYAt2KzOUvy/V5T7zbJLkc+4
QXy2KHdFdx5RYInwXvXvW5Z6YgZPuIQxdsTlXfJm279ye6l73jeL/baRhK8fYast
0lJI7JG9wya18E7F2cg+ePhR7IcQXHEwhC7TE7iVic6PgC4H5FgIYL+HygeW1tEN
doO21ioi+lFWQT1O/0DAtKKZ6r2zvBF8WmOGUP4aISfr6b4K+t2tgXc1SfBxk/Sm
lPcY7AfXy7PMfn5gZSQFDWHu8gVBDLHBaxsSp6pGZDNKlGioZ/Dwq6Id3iBhkRhB
YUaTJfjJybeKg2/Hf8Rzz0gXnneHfYFQbu1MpHV2PdEI2GizMXhVJkEudzSpXCgQ
atHUDNLoV6E4jp7+QOQDuVh37vOqG9cWWS6z1LUiqEN2i0NQqkL5K33QBX7D3eYp
TjqwUg06t0E+B+757+sWP9ruPawza6UuhkbHU4258H7avjvCElNb1LJlbAbuIDts
r1b0vwh5Mc9OUQU6cJp17PUi8mpjtYun6E12E70H3BoEhDdeemTbmZ/GQzP+YGiN
tIhnNUPPYdF+2S94uH9AMeI66PJ6xBBqPf4GAaRQAMZTNQhTl40/v4VT3bdeaId1
ThAgynMcj0HxoCEIe6dN3t7zNZN/HnmNI7o7f+8TUK1dQnVlD+JVyvegGSx6yXAt
JgfX1GyHNvkHjuSxRNGHBt8KJpjdeJWsuBHt8IsGzVyw5HNu9Eygan4QjFeawCg1
NPPUWvwWiCD5tYiSeEkmtciUUo6R/1IZjRanawrHsLygLoyhRD3VbLLt8G805DEK
sJcWpxsqpv02A8ejPQdrvFpBiAcq8oYbOZm5RYuoJdUvQ5C2mBcLpWbdT0EJWHv1
NblqYxfK5ZdcYzaM0Sqr6AeII5vz3FGw+Dq8siaG4b/TkmYnjSEFp9Y9xgvm4fKT
I8ZDYchbLqLdWy7nm6zjimzjnbyAmrdOoDm8FrtWXsrGkSQz6usbYHLp94Ej6amM
tGa07T8NIycHG8gb7WCQR+3nnnMDS2BtoJkuhlN4ILHWN8yc8VYDgmFoO1BbvJIR
Tv+ZXZshRgH4aNP3EgXyVHreadp4BULDrMsXUEq3BNBCNwaEm7mhhUnYe7rgbKXN
1iTjGwox3DEUsyqHOHOZij8G1SP1tE0eJLryVA8RH9Oipy/gGpLOVY1kj54sCFVl
vvURcwOiOOEBOpnpursX0VQoYEukw35k760Q8CXE6eziV+tPbtW6MzjNhOyzP5/q
1tfodGtvJx2OOx1t72yycRd5TcT5AdH5g3+wSgSIYBEN5FnLMk1ZFjGL7yU+NdGe
vdz57tLCA4pgj6yzV94gjsXhWpRCvgUKsrNIFNZ9oYyqJPOVoNtWnYZwvVgRFK2q
dJk4SIdUtXIYNC/fGv73M0XeQAPt18DzNcf48D6TXenqAukndeENEc8pGmjspi6P
mF+pVFKRkJ4bW4IBw4VhgiuPrKIuCyEZ+/JKdZ+Btm3RhWOnsOeO2TPBasvGwqaR
cSHpPP3SS+eHmjKilPYVAx6/7gKEo9zExCZ8znQj4hg12JoqraG1zmark1kl4ZCl
utztA7JsLdAp3SXV5lxLg+tn+VK433Pgd9kAeOvfCd7/uT+RYx56ft5pUHSHELJw
EgwBUwmd7qElUrLqlOcM9rqzIVYJY1k3JfOrJUtyjAz/a1tFe0HAtPfrh1Exm5Nt
2YBMw+/FM15D/LgiKUkkWdvH/tz5pV/2nSWJzviLBxPQxEb1IxfGR3wOmIHf8Hrs
l6FXNLwFsyMF3rj2QBgOOhTlS2GJIFXuf4f8SM/mO4XwGpfkwUZ3xhe2TlyHwc8Q
tz46DHdeiVa9u+OjXn4Ihi+Q4oPaOMGpo/oNbCKnNN2XCjLQrMQ0VduZv2QjA+yz
1BLpIqvPhpnM/HSbwNbt2gj4P+lWyo9MaSY3TRKScOsCvIouEWN7TR4A3pjHi63M
J/R+RsLcJ5jZbePESq8p8fIkIWtgjhA2zQ/EWFapHp7fbEiT/jyLw17T4S/e9iTy
vYH0q/3ZDfJjytZVaQjNd48HuwHkn4Wb/Bp1NAdFCt6I5Sz6fvNUqt/DQjewUgSu
wZ+AmP4Awza1Q0u0h4xdSyVUutzF1lFBjKGjf54ff+GLmXl55tEuYeaIlV2cpClE
R4Ys64lGl4I5HqBwROxs1SCBFN8oG20z3KZGGvMZ8XN3KJct5oG6VKZbqybFjbzY
M5ncXRclfujAQ3f/UyuIyPLh1aFI4CZyDuaC/QPrLIjMEZ3/iDoe5sJJ423rPoMd
4MZrdJ9szf/c+Fo9GYgeMHh8hBEtu2TxSxofQsFZp8f7OFcbiPwp+cH8DU6183ts
IPSz9uQeWJUyRA1juVPs0guSaL/KX41jmRR7il+FWU2PczoxzCGwce/CaVhnLkf7
v07GNj1Gsmn3CkVrJ5KbEtTC/2yNbuSlJA3XgkeNRDN/aTuRvj84RjsbO6Zfm4c1
UO18aKCJmRwLR0mepD8485hyIgEIxXo2k20pZdxXgMIOl2g0c8IKHrWnHtc3NawJ
y761Q9FB8vFulNZeo1v++siTHC/zQUoFykahXcJbk06WaKNj3P0a6Y9PVo9Q92uD
QTgxcp6PLCxwhKIog5kFKTFKTSqwnNKfhsprzJxKCyYyLR4EMPk3ysGtFSG4ffte
2gzz8KyRXgMZngTAmgXJ3R/uahiGX31FSU1L06T+F1SSQUK12a/yz7C3Adw0XiLP
AyRbOBPDoD7UkiZHXxONYuWeoGz7hN8fx9Z+r8UaCe9ph8In8YXpHl+yTvv5mIqq
mJun4rEq8Amxf0IcEii9a6X67/O3ZRkXZkanrxDsBz429eSko1/Ty4i4HUYWY1A9
7f9DLgYrP8sWMke7tOywKWa/YOy2BBlPdJbIn/lmNR/X7Jk5O0SlFvDe01449Bec
VW9G0N76bv+wVwkYEDy/bRhc2ls2LS9Ro8bq8PmoG/EyO6IfBg0qpnxQ/vCDt6KR
nOhPhncxVV9Mg/gIHV69xfYU240oggHqNWxsKDkg0hZTEFKX0GBCKPWUeuFxHsps
BbKUJ3wpvpIt9mveELs9ejxIqi0OJe/cgrZgflRuI3Sycj/z+xV+uwaDsO4NkdBF
nu1SyGsKGasc5DeiRhuyLNIaX/eieNNZghTWav4OkRKDUGaTG42UCJYIbR2zP/ec
oKrKLq0wjeEwrEFVBaYatqIxXfpDelv4NUd7E78C6xKEPquDak228ilHZpoQ4it3
vscGUq44V97mf+ZaTbrTeTfMgI5DplV/DmJda3ZQPYxEXqQsgJfCS+hwfmRL3UYf
BD13eOqnoiRn4WyuYHM4gcC+lhetUtJochHsopH4hR9qFgMDKT+ekVw7/9mBvF0q
PVZQHOHDwVH234TTWYsvrpi/9IiDQGvWTAck6MnGp+9+fztV7rBqat8OrRMTzMcu
X0f+xFqlniL1ahSLDcZ4qGFLc2E+HZMrIq2gobQVaDtuMABWZHOgI/T/qN7BJEvL
ZvgJNN1LpWZG8VJ0nMkFwcTa4omLSUG42NmaURmzesP1Xmd0RnlEnTWvN9aq75kM
PE9MFe9LLyqJY8s1Hn7K6P2ivLiZ8PSoRkjg9Najs4jB6fpzPzyb3OvoNVJKvalC
vSokHddmtMkImY5g4K9t+JeQkLf3W1KcUOPOj0Kf9qMsSr4Ks/aB9QnMKmdUSKV9
zRHxNZBIcvZxja5OcSUUfKY5BXoyD8cYMjhHsSI4Sxi54NW1wz0IOlidqhfhCc3z
WcPtYje8y0xMvKojl1Y7GfmEck/Ul41zWi3FBWupJ7eK3H/bvH681PwanXlv18R6
eInv1lAgRABgZLcoBFdY2IJXVZ7UPe0BSh6wFLnHTEaHVWCArDKSUl91eResA9wb
U59AWEgBkHsz0RFFVMb0b4gownhGGO+fDkKHGGhgDZ8s33NvUkTTpNYug30rWjDT
kS8J+3WBLy5LOxYl4LpqcTUYmVX2cpMGRZxgR5AmWydb8+/rvoCYFnlkp/OGyFdc
6lRs+yU46FMx1GqKPsoGOjvgBIiSMzsPWyvKmhdcAti3Kt1owcTvPy1TibtBA0F4
XzBSQlg5WMTzvSqHwg4P2IMAQ3altbNeDe9dhoxz2WNsjbJ62cM4A5Jo+JenP30o
xTF1V/eFU+yeC8BPiY8vQTJkCJeqLm719f3GSAADTdgjLoL2cvjZ1o/7Z3zmoLI9
Wjs7rU+etG9wwOtZmYFwrzNeUtlUglSncC6ea/mMdfu49Sb1wXAhGp7j3Y0FDWga
a4V9AkRtXjhrddEnUku7WzYuFydGhDPiDcfwGZONJeMyg67EdAWRLj/BbUkM21fP
t1zBhLzVMYox6jXyfTpahcGxm2nNpACzS+njyk9msj4mtPQ5/D8e2SoE6K1bXrnv
28hYSdUdxE+Cwwwf7+KIiG/7VyntkBrAmLxJ+h19XjtITw2Cs6fQvGqeuFa+grbb
5iyZC3dL24PwUkkHHoVoZ8pW/xo8di5f9VJwV0BiPjYFIc1xAcx+8A/CqCnISq+Z
T45i26ITQYZNyG2l6jlhEvKP6msHA/28ej5pjdejj7QhPir4vHaiJ4jCYx3693a0
EEu8Ltc1+AdYQbA9zGLuYy5L4UTWlLrrw0jM9pJsTXMpvuvbUWNZtVFRcJNCQuyv
6z6qwqAmHIb0KSgCAW+9N5HBgyMoj8B/N+NZdwqEYMFziV2BiPdMrz+Py9GYVcvh
GnbYjc3S/m4FJBdzJT9wlmTkGjNgKRWv7lKODm6tRfTvO7XkdMvv6uE4dOxZvGCV
ZJ5oE2LcGHeLAV3qEe9HLbA9x8otSRQgugJar/HmPFjVFhCusmM1t0RAf/9lxE/U
h/XobRqWUffutn+UsWYU4wj3JeB6vGebWJ9HKEd1i5jgtX9HmpZ/nzY//2hp/dlW
pu2EVLRMEcYBMWNgC9f432E/W/Pol4180ounkid0jy737bdiSwg9VncMIFobQObS
+5D6m4CV2QedLLvWDuWYcQfC0KvmC9Gks6bRWbr4rxpeou9e1+sGgqDkxwSAItDH
8StUg4tnCSBbPnVEeFx8g8PqlwOIm20YJ8uALKXPYkF0j0huhXDc5bTB7uigWQzo
7gFt5pUWiKfDbuYElIvVS1gz23rkkzB72Co7zjlGyhEdEu+CARJtkT8TE8UzpDxu
wLr1TRP5ZK+rA53nKobtcQH7LSo+mJXV0jqd2u/l6amEP7/QVINC3ZhicyWvcfib
xJhKaI0zm3l6Dtk6iDMAFlJSp24v9PwmPcF41UlZ2BBQZ+uUoMo0ONyCc/9850P3
nCkeojJhsU4CbprDcLirixxS85kEG3AKkc8sFYoVgiURt+W/PmbFb1WhgPqRQbV+
8F9ozeOmNt2d+BqhQ1NT0wdZNBrL6BIlkPdU0tTGvQDT9FhfYYG73kKRzg9pDWme
W2SBisqTvyVO6oBaXu9SjPbPT6D77soiEzl0PuWs5pvimJz2uCAle7OiYIH+Y7y4
apgSxLMRw9ee6cWhMQWkhpQlnWjZsx8I6sdE990iJ90iIKNOIxqIKzRf+8vGqQOz
iHESMNk8ekx61EfrUpt3wEl+qfWYx82D7WxrGHwIjlPLtsIlY9DbwIOTURg2jFdN
pEx/1MmMZ6QjQR3qpGlAE/yTjMZRiBTqKHSMVjKQTxOAB9iUeOQC/Bikbothg2Xq
kH2xwIAlN+VilF77vVA9DEuZqAW25TpJ5rveTjvSwRxbD2epJUv5/NJuiTWeWJLF
oTeUUP3IU9Fw+5uPi3eCfsmi2mAevHvNQBN30R4uvESdriJsn84nxjGFWKTl/wAT
uVzTc5HPELDfKuQSFRhJ6Fyl70qE+4FIrJHUnDzXo9D0j6TjqM2AlhRwuZcEU30q
AX8FBa3ua4s+fb+l+cVq7jChBFNjtw1RDNAgYgb2Bu3FZBU6YgVxdH8ULWjv3z8Q
uIf7zfKE8NxJTKC7267CBe+zjeWLk5InH590fcy92z+crWExFMotmJxx8wwxtQTM
ykO7YrKmv/SyVolIR33pzemwv/noMbCcwM3phk8UXXdaH6e8Z5LfLYxTrceMyr3P
CHrqMOrM5W1jrX5xgAdWXMULN+C+UsU++iqD3M9by0DJ2jBVn2GnJTwT4SHsx6F1
smMYI1JZ4nKx1lkQlHakAH8KoZ08wK+qKY9/RGfciyl9284ZLao5j4WFSLkEnyHr
GwuHirzpbzWEuxCou6sftDkckoofLj7ju1/X145igpUBo+Kd5KXd3Fq1dWAgDmD5
vYXwK4sazHP+dt5tkSi4omW2xT1tCkWFPPkCcupgI5JjEslZxsAijjJ0KusnOb/R
O9Ho/tjWiTovVZ7erhPw6FbnhBvD3mqSD+vMhhHAojM5tcev/l95aba3BMezUYE4
V3RSwQZ+IFNDxG9XBGFJD++E/Z3rp/+D5HAuwPD+jyWc6bYK8v1t6LL6ooI8n1BA
UbpBw6TnY9fftehcgxyWPUVcujs7SE3eDD/f7Ay0RmtI63hNilN/12cZHG7cHSdW
Ol9QubT83MXZg5kEFS+bt9fCzVo+LlQTEo4ZnxxvY+d8Sj/8tLCtp8N/MOZwqFYF
k5BntOuXl0eXkb/2bMHA5YV3+pJfP0i1v+IA9N34nVeslvPMDwxZ6l/bQjdNogV9
nf13vRPDWFLyTaFxgL7yjmGuTiagPGKjLLdd6De/Tn30C8GHUgBY4IHMJRXpdFEM
J/XogkwPY0s/Ye+BHcxmCSPIICexjgUh9hZXkxUgx1FBzkYo4oOuxgMvDWmZ1ONE
OMT1Iexkz+ca3XkfUH3xFHqwkIfsOmdaAOe1Y8gcEAw9N66yDkgY6ACZzmgXWSNo
++NG7JV0Ns84sVr8hK1rP9Zf24FDXOlbatIiei08ci+kW37RNokFsbZ522ndHnnb
ZCkfVyMMDErknFa1zSq1W0Zfb8r9Ma98qADsavCons4Mpnck4dm2e7kP6F6LaXiR
ZmKWWwC28VJL1yAITR0Ng6UKm7BrZL54HDLBG9N/NSX4Mdcdg7qRjjgA8f4sD1O+
8H0b01x0ksOO/RGmf2VeBdohiepL7zyka23Wlz/QO0Ut625pKqlSDLMH+UuxmaZM
7n1Oa5qwxpT4/MUjcSX/aFUVCm2SvuI93eg0V8OU2CuM1z690SLTkD59htJq3rTV
MzhLMaeKuFmzEDtF+OSLUH9ZRiYmUelrm57ARL135c5nGRY4wejmkBk7+u4bfufs
52CibxSFvdFd6z35dosv+aaUsm298uQxddgmVhp7vqQOP6Vh+u7Xdp3l+VV6xkOL
6b+IPuiuIX89Xccy3qXqezyyBKcwGU+ynF8uwpc1ErO3dsiH6IODMD7i79gYmqhj
h+AjOupkkVwjJ/FpcO9Cg7+5gW8aXKA8oZ4Be7qNImLnucHR7MI+g7IQSDTgRXfm
1+j0tlSMDyqYh7BZKEnqPNQo0DuIe8r0BaYjsE3L4FWJnk9z7s13dtC4ONnnqIUp
UTzqjkKKw9QRzhwjwWHD04DouUFYKOhZouqiNv919q8UbIhnX5NiAt3E+AURKHPQ
3tMO4EzslR9DkFdS0CgHzNQk9kcJGe472EakxpUfgpxBefKHjW741P4aeXq0DymR
Fk4xo/I6ESccTBu8Vvr0gKzvcs2iB7nwb3IQY25CdxUv6VVJzO8zZjQGNAqJ2tB1
OeQX6xH68MhtLY2OoCwZfcSTpBbDhEIksuElpuhGPYgsGzjeP8t0XfSiyq0YB3FN
+CpcadTXl46LVVIIOjUyDkLiOevc6ZjkjDyqvAMN9fMgTqHY+fYbxpnhaA8zSwRU
VhIS615YcxX06pTXkTGpxMLLe7X6UTUkbczF6Y6kuiM+ADQ1XJ752Omm7h51pn+l
RokCW7iMfJy84gxDbpusEqcXXdlnITOHKopTCdXvIZV1t/KGiRBaNRVKyb6M4MfD
foAW7l+KY3AIVBrWtnthfT6KVccM1QIJLqPGqw7xExtVfJXYgPbka+XewsteQNkA
eP65Xii9r5r2GVcgu8sdNshFDsKjxgOti6q5VTVoNK2albPTafcVsxWXkDIMLQtf
8ePsrFt/FfrW8x53tUlaHPxCUbc6cWcF8vBihx8TMdmpd+Uh5fX0bga1bnGKeBSI
KqUiHWAZq9w3fLz4wFPCDqztmAnB71LmY5rfi8Nlj/pDRFQcnrgXo5G+Bspb6yB+
IPOsN+iZrccFKzKX1UPL9TcMUcBO4V+BiSYUjXmP01ApYrijqIWbmp0AQng1aXX2
a/Bu4TEX07LwXOFIdRn9qsbTVGqdl2ZgTRQlkZl7A0eU1v2A+IvXlky651Ag0l0A
NSb5CB7gef5WVAbCaeHit62MYquV7st2HGhC12qwr2v1DFIU21vaGwiM/LoXPP9D
nO1BgTBYO7PvA+i0QY5RyKqI0kPpo/VZ4SPGkMn9fjkwzVQij5ye9cbE+mPnyoel
9Jv2hCbXStd2LVAxewTqt809YRGH5SCPdUXNlDf8S8sO9decmd6NDKJTt1YmrJG6
85VaqcuzpBrDNZbcJS3igAjaz98Lm5z0/d88FFd+5fxDbvE+z1Gde3e0lB4m6Wf+
hqzzQbTkjIshE/x5HmUl73cC9rlVRZCLNtfDItfn7ZkVrmgC8V/ESHOBfE2sHpSD
R478v/JJSqRVInF9m5WFEAZnntOSyBqAGNjiV80rGwlX0A0K8vjoUPhYGGiK7sGV
5yP0BNrzDTFY3ochoP7WMk4gs1wnOuqggn0JAinmYPi1CjrI5VOSeSWgfout4BnU
Pwr1I2jPEgCWAzCmC5IIKWkECaIHUmB2+GgC/t+28PxHS19GlQoPPND8liHZrbCV
VFgqT/wPX2TeIVr0N/eEcRKH5D/XVwC6IHtHeqx+tQr4fJpyFGiN7fZ087A//BAj
x7VTgwj78Hpbu4Kili0jxXiTo0Xi3bYAGUnaPNszygBTiOy3phBAR/2fCBm+dK1B
zJ2oSvBhsflic+QQtIx3sjq0NOTzN8HZsBuLR7u1KPy+/rCoXv2Dwy7M1OHF0nRX
WV5lHj374BWGSOA6j92rnLq7+GxXaL/Ul77pGiQeXeypkGO0K7i2Ijpnf4DBQ5yP
V3Ka9EBDwwTzt47zCHyYEvMvexVO3aKk+WgAJD+P3ATdTQMNutq80EM1GPWdptDh
qDeacye6cPKbWRz7NtbihY+x8eliV1fHjtgFD/8aVQYL4U/o//MeApi3xMDQkULO
966k4HRlivK+XVFkj7ktF3BHDqgcftQ+Gkb0/7MzdsrfsaUEZJyRm87ERgY/UUES
ZtdC8ZL2gdBNf1F3U5KHpF9Gx/SEKrlIcnExS9Uh2FI3JMXpgDWSJPOj8p8uNZfk
10jov71bsfDGQiKWIG2aCspRiWelOE4RkE5IP5OY/3Qm8T7v7u9RCN/BuYiUg4Te
zCsXe4wBgcgzkL/jRFbVhj6TZv+M19tbk7HUVK1oZWcEP7XO2jUDJIoN8bdraLL0
+IpPrEXKNas8Ylf9ZqEUPPBk5q95U//xnRvNWcz1wwW/2mM21EZoRLxrVpvye7me
fldp0i84O3R/hljbSOREhPpjhN6SCNVg31x/Lk0DNQ9zueRyfPiUEJet8RivIzdC
tK/1VgF34P6H1dM2K6ZY5SSPhqnkOwu/EKWH2KDikLtQ4ixqW4aPbf4aSaEGSC3V
RM8gDHT7ibXmZf1+ZwrKA2BbyrG1e+LgA5txfZSwmpPiB7LHJDeqI/5qQqwk9zJ8
Q4Su1j2NyRnF+qhaoaeQGwe4uc+2U+QDfY2/xeFVLWCruPZyzKkCsjymWfnDh94c
6b3ZqVDDZeCfA2BoEBlsMZbkh5/ZRF80UNxViNVCXjIeHMkuS1ZN1IpVq4kYsAoY
YWRzz4MucCyoDms13/AIE5Ys0ZJc5Sa4KRYEsV/ZMyxq5QsA3ilBAJnEHlohWPwf
ztyX6SWkedghh0DzyryrI6VaRWOPCIyrK/sDnVBpGQ0E/6Xg4b873bQRWCIPH2zO
sFtphaiNKCS8BTzqNgr6LnWnedw7Wl9DG13JmF6tOg2axa+3xF46iqBMHY5HIP78
JPikXz38dSGOq+sktTGSiNeQOr1ejjWb9ScC/jFzUhq420isM88WQH5RAvD1/0Ro
yilswHlOLMKzkfnpNuwpiZ8n79Sjb9TuC0/0r33Qwi5kfTcY6BBYwYHX3akdL30p
hSzFciSGTqE8s+GiGO5liettUODiyd2Wd8+t/NiHNOeqnQuDiPnVkn8skby+s5D+
zvp+wp1fk6kIHW6WBkvQk7FFbVeSpULghejvJoFF+NyMy+EAOTW7LnYSkZNrlvYf
onNeamoeVo8a1lvkkH0v4km6kgsBRYvFSUEjVFBtoairlpysolBEsqshPhgVlAxk
PtwjCN8xmuaJop39KKMyxj+tVg3qVITHQLuzlAQu2GjtaVQ6mOUU3bsqQMcqIQFw
Y5eIrsQEW+hB4v4E29eq31zNmR8XnuQtvqh7p4uL6PkOwSG/xgzVrTV11MgIkWnu
veRS0KLi9BU3Gcf3ayUDP4XgYWAoKLMId9E1NpubarTFbWkK61WJRUq/aQ67vpqE
JxRtuDP+zui6MWl3ZJ7w39OrmSSj7Mq4Rv96ytmC3Bd+SxkC/CVi9lZooQRVhnWU
N+GBFUPRYMzETsTEOjsRMJqRsnsPoobKiY84fX4dpfeH3svpoExcNv8G0GEcNOu+
ZNUXPgr4fB+QVq4zWyTLNTkDhMCWh+lY3hrJJ+q3GTrRKX8U1WOth5lggGKXnA9k
HNWPaORpUnXoPqlxuEDPZN1ZbVNLfbht0NgBKlj5CujzZDzNpFJ3SMThLIXdbLNp
P2G7JkpWK4Nzckb6Fhw7GT4/1f1fLlPUQPBac8ZDOdjmU6LSGpPuDnGkQeX0lhV0
gBTwv1W3ruh34s4bxTPc4VGRPEt94XKe0lM6LPLQYiZK8mfBZ4Lk7LlYrgsy3DTV
5Zp6LgQ6jZqcJupSo3R4oTCF/ZJL1LDaG5an+w8XqPNYTRJMSggFMsWggHDdKdDZ
flIFyKmQuzKxodX4AFF6m1bJgOjDnSxiclFcc6RQ8sknYEPHqsEw9FFp/QiRG1hX
hfjgeoLXphk9rI2Je8Wd0WoQpji9gJiq8v/LNyRUPxWjlOdqb3bJhidpGG92hMUj
Yv5QNCytKwJofAScL1nBNBDHo1A+X4pH+A4Xy5+iNfdWbISfERJVM1PpH4B3Yom+
7WRE2+LRFXSAt8Y6yGDcUzKe2b0I8aozidLwe3pVaTuh1uGALulhqqEX3Bedg1kp
TbmI9CH3ielrYD0Q1FRcvbuWGKqHr1X+2SfPCBTGt95txpXR1R5b+hsfb1CTKp5U
RjnpgsPe+RivPrrWFwWSagTL6tWdTabE8U+ktkE6ZP3abX9YXzpef7aglxgwt9SU
8n1G6VdfshUHraVvWxobEY+emfasR6uUaxVSl4RpWO4Yaf8vKS2mJ63vM43rNmVU
NDgtD22Vb99UO5W7LhUOrYESSGtstYtfmkJ9r238un/SbbcldyuCSSdyI1qjqeRt
jCyb7wtWKL0NTozy1cJluhSUYEFFt6D9GlsAksco3DJBmmi6GFVQGCQi2r5l5kCs
wIH4cFnEmyKVwOc2ZHSMNoe4AYXvV8U4cduFulQCtxVe5ZGW+WPNgSBaucih9Lay
eN5kgM0SSpD5Svnr0uTzvWwXRZ4WpO8LzGEgZnk8UBpcafVflF+a9vth3SR1ehnr
909pRvntxeK0F4XqWm2sugW0sAqvx9Z9sbuiW+BNyKgUOtdfhydigPzKhK0TbplZ
JyesdeyfeakcxFAWyqde2U4AJDedPG9vL3I8+jiLUOZW1/6Nk4Ey1efkwwptQsU6
auV6WYyZd5uRq78Od0lXL+/miNSEdkGlGiWvgtcacyEkkbhvw6IgbBz78TzD8nhI
/CrPuBhnxfUj5xkKqgtNgB4SFqJY3MU3WoaowkBl1iMOtIaOrMcRVHewu8gM9wRX
Hj1y7+zfZui+Hzl6LwbEhUFlNIKvcF2+ssOfoq965dr3TX00v+5ovKwz/q+V+ZNL
qKScAyJYI0dZD1XsqRxQt1cnp6E3CZduuk05wUkj5h9dz56kKnaafvubOf0ZkkGg
P98lcZ3E9BSX2tPfwvuj7Hd8cvM8wg4ALo9BtXPGJ4kkNmTal2cVg5j0hqetqK81
WVjuXMQqBOkkkg8W1W7FrWnB1Vdc5ryqr01VZF2NZIxyTye0iQ8Tu5b675Zmk5xH
q24BCH5EJKRevzU3jy6AUeiyRuIPxlNANrvi9BfXV+PAKgfSStUY3ZWci3djRKJs
c2BxdkWzSLjImcDlJSdeZduUWfuT6YpsdISNeXpXDWU4UhBO+bAbGo2VzMtYc13q
yvPT45Mn/RgFNyum1XFshd7mRSOAvrxvZ4pfApEUwR03FQMzEQHj4baUYI2V5axA
SXawZBpEmAl+xyy/QH8xxUBN1zcvUZ3zvsi+zKWd8d29d4h7gf3ev9JeY7EupYRs
5V4j0R8HlXC7LJ4esB09Y4U9nEVS5VXWA0te84ghL8Yvjt3nUdLXbb8Qp5HVlxOR
7Rxnuwla4SEMjwbrYEKnJmp7CwwVLEkJu7dGbNfgAUzDwWS2Ny8wd7Nf4ZCuqMbf
El+HFN9LWlQJs5PaeC/TS8xa5PdSpnXgM3QbDV6+b3sxgkZn+rWthBI4+e8dVptq
HDIXqEKhmkwpFDyaU19+rbHBZu6UAgjwGPuAx/UU8LLx4JDwaBtukldAN6ABFJkG
hMic1jQwQGm0w4WZKRpCkazgIm6jJDsxqhJ+yoy1mddEW+FpCAmDgKp7QWuD68IH
7OdUD0OAtgg1d7nR3f164ba3Z5gM9fToEWNS3jxolWmNB9W8qazhIV32k+r7nihI
GWOowHDz7TeeKtq5pD9A0NpmHyAiW4kbAnwsDoQy5Ffb/M/lK8CADnSc2wA/5RR4
io4tIIx4HUaGIYp/ISwdZ4C7j2uESZZTpdlzJCA03gxWK85rFAH643Q39zCis2Az
oEyuldyF8CJxrCkGunchaSCiFZeYpxoRzbpga8EPtwMREK0wuMNi5bp/ouZaHnfq
R44NTa5jhFNauE1J8fxahKH/J8vqRxjzsTtxWoY/SJjgCxF1fRuEKzYSq4Yef4Qs
+IXw5HJtOaHwgGeI/6S0yVPqcGVTiLCAsVLXof6Ooi2jyRXo3frEBxNSje6IsVml
X6bIL4fqbVVl2xJC6qpx8hmuqHHgf+Y0uzeZtGYUd7DqlbHO/fXVA1CtYwBYop9o
GDD55MUfuqbPnQrowe3YuCfmfhllv6+Q+pgrUtOGUwQNnMHKftPeNCIvGbA+Y1Xt
FtN0y5pU+UzcY3IpFpnmmMZcEfMYcpoUBYtSlPYcx0MN62qgEwTTZJiW6BEl66ky
vi9Ud8SstIXKJdpiznANMO52oDkzsCUSMOJZlni7Jos8E6MXGjOcfs5dZOxv8GVC
rBzxDOepio6AlgVRmNS6MSwP1aMCE/ouSVzOgdX/okQFf22AdYkf+igE41bWrVJ0
aPNBDS4zZ/RFlqlzesY79eS1fdo0HoYbq3UbgfBtgQ0CiPVm55BvTtTuXBUd5wdC
62ZPjcHd0uXJSyudbVweDCdDBVpOkwwV4ZeejusVEPquv8T+LNSiLnf08ajipVji
chn5KB4tgZOHmWxvSkkcFCmygv7VmYbEpmfIHVqcD6r/iz4GH1EXpj+Ow4LEloQ3
cwU2U1tqQ/kLc+XYfV1xxR9HEGqvvtgaa8w4PBPgXnKlMO5+NSRrUq87tmr1WgTh
WylMeHyMINxIuw9p7sG1xRxtzmwXRnoog5jBkhuth/dVYZ43mPCUQkNx6dVD7Wnb
7gZ1hItvSOrCoiA70tLI06PVXpKj66wXjdUjijHbB9T00+p5ncdyjvzrlVq9b97a
5o52D8Yf6ttYwEA/MH5OpDG1BO5+5Tfy8b5EOoJVPW4k0Itcho6NxiKoHHfdP7Kp
UVQqn1lx5jc7XacABfbJS+1onFgxzDDFK6EL9NEQycWCxMZ+ggKRzpo5emIReUv8
zuWyFHmK2XVinPzlM898PddsUaKeYBgC6rLXZH3Yp9lvdAfbhgK2xmcjOGW07Gi7
jJqZTIHoXlsCFGpiQCU4tGHnOqHryx6z4cV8hGI/Gm+5gF6juNmHoqTpVCOEm/tG
mX5C4H/HIuogmtGZo059LID74vmMl6sge8CpjzfdrrTOCHtzxQjk08fQCqZQ+LT1
cMUfWD8YJPmN4K9I68zDuyNMc2Ct6bJqsOaosktsZnRv3yAGyg/QRSExMe6wcPf+
FXw131ZLi7z7sINTrr2+g9giMNTuTsWdN7UBJ0tAYMW4JoeTTpw8Bg5tbQWQGLpi
AUTqEoVRC/j2kxC6URRQEy1U0BFpyiPtm/C1iiM7ZOWApzcgqS7VS0NHl0a4A1PZ
WXf/fsiy1cEjnIsH5rBGgCbs2hADOkjoSL/d+ubgVpuHaWFsGUXGw/0kGye385/p
otg+szKNEuzKMtjlYnz0oO0K5KTrv4k3OHaoeV54upMXzjsWqPmNgKVZFgHI74hu
7P8/0nlVorm22fCCjEN2KPq344ZJjb26oXLCrNyTTAjnB50fg7VkFvk9lQ9mvO8V
KxKV8EOjjwGeShxM7bRpJz4DCsQz9BCK2816tRgdT9jGKqSey5bdE9afnWlpRND6
87yzt2hd5jePh1WtMB1hX51U0EVT6fkrIGgne1LKSp12nBn8XtwBX44f96Hc3i8Q
d+W3E6lN2dCL/jG0b6KtZ5y8/mfLDAXcqmpb7AybPMUxkai3kxCS8hmtNS+PWuXW
CVl/GYYfxWKhiV1tMnxsY/BbIGQ3XugToiEqnXPtl6++Xv8B52dQyyqL+Dx4PdU/
SRd5V4ZDIKqrMi8s0uk5F+ziUHoxMHDdcdJ3z9E29k7gMo0SgZsdHAujcvJdfvdj
NQPPeMTfomnP0D687mpzuI9w49UC945gKTwjGU6oVUsi/rxWMD6RnNmOzbkxwvLD
llXx1E0XD41pVslbb4uZSCSj2TJ8gxpovTFdMlpY8IYJnFz+43Ku3o5mSn8jANua
KjqsnCVGQ8C/FWi+HTFsTYXPfIUmSH7OFpQcuJMhk6Dfs/XKVx8B+RuSMYllUG/+
L3Yv4hQF4kDwV0xhDbNxBr9RHl1IXWEpWEISfGWn4GY0dDzQRfXmBedsEvdqU+S7
KbQbISlKLaRdscIhsr3wctYj/gtVMV5/iOivYx6psDT7ji+UDiXvffHvtR/HgVnz
dcAZ6EvCNDaHebIYzBfMIpZJLMrgReUb+ufTdszrgSPNIkL/bAmPvblRske068MD
g1CWKjtUQaDIpkX4daNgnqYLJYXBf6caIbI/haSrYxn9TRUMRx/iFFQMqwlehQAU
stjnxibBFXKrhqZMttRQilKcWuq5YNHpVziz4LaM9kAuNXiVXKMdC3rPPHzSAmbl
uprxNJ5c8m40oVaaR7sILhWg2c8YDiBcdWKfokjqE1ga42OaUQpRimxg+tDsesEz
LTiCIxD9fLKMxAsghoXDXDadBhQZNYmj9MSXV/6xho2/0gPB/UhWBvEUNlgZdi9H
nj0sb+5jbP+9oZbZquWNIoeFYLW+kffiY18i03cxK+CtAZd1cqko+deEvR7AWkUK
ZJs5++k0yHsHCoQTvG80gvinpeVnF+w2zEz5ba+KlydRDh2IgY95EKQmsvqZygg/
FwFT9WvlBPgE0LP9tcYJxIMmogpF9bHcTuzSIu7Gm5tNvqTKIkw+5QZ4juGAXpv5
SvVkcQfClHjU1eEpG6SzzqAhaT/h4+ChDs0lqyF/nns9tX6yOL04z7WqvDw0k6WT
IMmmPsso1ovhG6lWPXnBJORsL3DLA6lnSiracei51MvdqZyXkGyd9TmsbG2ruDvk
44dJST5B19ddFw/591LidX27gxX0gVhfH4IqULQJE4vCpsymi9uvRQ3s/yOpMDp6
o6THWPBasubmnZuMd5duM5jXYdK1mwWeugmUAwxeG4NuuYsiEg6pEf/uUefO/6r4
GiIBR2oXUroFGMiQ21Kr6BDXcCpbpvZztC4PvxxV7Wa1ixNgzmgAzChZ2zTB/1I7
CNf8uG9sG8yFQTV3WydP6RCWyBummVar68JBUpnYnzABum0Z1J3/hJn+j4MeOtQC
WHRffFY5OAirJ5tpUdi8iTTy3sq68kS8DFV6OG0Vy5xU7NNUpvPcjXL9y82V4Ezz
koBT86T61qlrDx8ONIy2EyihNznGEQn9LoAbvYeTDgL5pUYE6J8JeWINtSHVylCI
2QU0p5lJxpWkjNFhXwd90cZiMGnhhEIk25SqCsT1u0y80GU21xrYd9dHMJze01c0
R1suTCVoBUR3lgF7BQNUqp9numT/VA3W1wS/RUDGpY24pL26zoGqs5wrGewFF16j
s9v+gNSWM8jupGQIkjIqsLHPwI4UjYuSCIpvPXYLZzpiJzO7kEGLmqkSI7bvcORB
hwRODym5A9LUHHYgRlzk4gIy6Jizvy24zD71Yk+h6l9R4LuQoeaz8X96wDT1Fr/j
Qf7uyRZBg02CRwiZx5qdXrw6qtyvEWz6hxkIPcgbUJpAbDuTiYEY9L0kg2We3Dqk
k54Z2OTZWtU9lJdnNe6ctiHWehiWKYKqP3Q9reykaPG90tL3XIjytmZr3FakeGM2
nwnNjmZmsHIPGQZ3QVwuePsK/6Xz/n4bw9kD4pEQBgfaUYDX7B9to6M9URwdyejw
Voq2HdNWB2pAKb5Mxw1KgMElXjc7W4rjn+C5IPE2WJTCq6wlpRlZx2LsumgFiVtl
lXRHYV2/PYT8hu8cCuVQHijLl0QbmwVdyepZOU7k8xo6bbyuugho/ihPbtu+1NTe
EiOJDORhSYXeweqMT4p6/UPL4DX2TYfON5a7lkmecXL0RHq/PQ7H8OUhvCdAvqyz
1sPIeY+RmjdIfJ1cGbWrhn8wYZ5/R10VnJiKfko2KnT4ZHgwL0G7PJcQAq2IUr/7
5hmHgsmP/vMHIoSC9AU8gNsyk/pvTF4GU5Ngho/+CQhEPtdVUBaXCWyN1L8P+Aav
LF1+23mGDL6kUrpl/D5mKay5m8FK6i+lXYYhALNblw9s5G8uzELU/7Ugs4Fv+A8+
N3vnBhqrdUQS5nis7+vqDpePQz+B1+LZjbxNqdRbPaFZ3XnN5gha+LdjOWN+WnCj
d3bC64gBCu7ClXUXWnHgDPJGdiM7PpdkGJvbE1L2sIen4I8GfF3Tsf7jFYmVL4sa
Ji0T+GlFm3zv1ciDookRSfd233mxmNOroLrwlQdlfqNgt/h9pnkMClghfKdJly/4
55U173usSQHK0Zavx30Yz5tVxtxlQnLQ4tbvzr335zq2MFPdzLBmcL6AYKb0HOjt
88ayvN76UY0qBA5vT8O++U2g3CX9l6osF42D16ONvy8lUsFzno+IQDkmN94nT++I
QjXekXrGAdC4UfrmL/xJrguabvKrGoHQzObz9KceMwrTYseTeJ2YiszZ4FzPSPJb
2qKVqfWHBTvRpJvbYiTgxbwLmx4IY+U8WnBj72GL+jEb70qG997EGH9XUjw8VV0+
dCMoODaQPiyupuo7llINFx35s2QB954yRbaFxTOrgB9eYzuzf5CLC8SWT2ycnGpR
LQcWmkSu5L6ZLJB5CRXi4/vLGm52u+zJ6Nz5VxQM3R55MSigIgC8FcCtcCJXYtDE
76H5JHVWjg/ZF0Uff2e9smfYvUi75uIW2KjPnLV22orV0w9byKicvhfM9FOknka3
tVtTszfVnWtwfe0+MnrkgTrf5hWkumwuYNiKDu9HJRmwC0Tn3bkq22IJP5P2yxrC
Uh6/KdX46nsNAwCBWeB9x2wBbF6uki0wAjHPkWzY9Z08XzkJO6JjuQDid9/x7NvH
XFqwC3XLs234n/xt+b3p1hOFEOOifkQJAUfFSrUtsrlBuE4TdiZdA8fRHjiYA1JW
zHfJla42IIR2nELju7afC4fB8Zuw7zii/sA7qvgUuI9AW8djn9JiKjdS843U3SUQ
NRqbB0jLucl64F2OEaAlRxqkmfqZKhTxoXOPT2ncZ9MD1+aPT6eb6B5Epkc0NZE6
zeb3u4UBmkgPMH3MomXCqz8/kjLY8mKVsflKn3ZLYc/QpnfFrE972AgtKQactKX+
71KiLUNCbCLVBb/HyG4HGzfhQrKetngBYDBIjlCP6EfTYhi3Mon0HJialH6nXqk0
QEYFuBSqYlFA49nNJ5zDYDqW19WmvYNaOLj0fIcBhtTNr89srZw/pKFwlv6Qoh2T
Z0yNUFTEDCtSFyU6KIVtTf/BqW0SMrXdvWTF4DAPjvyrfC87GomhIA98WDGhU5aw
7V/NVN2ReKWEO2dZ7PGMC9J7VkmzKjtWF64Lb3FVKqsHmOMhdHsYI80dNFJfgSD7
Z/d1SB/4WoaxxZkiiVbBq+jEmu+g/C6t0Ft7fndOj6IGkt1zdfzrvhEvfEsg+VkT
kHpoMnlywqi+dlW1VxftXtfotP7kKGSRAuCIlXic3b/m1wMSZxZzXKNFGaO3rlao
PllN0Tq4oKWaY6TB7Xb86HZJWHxnFbdp8ypz+tdV4zWoLMOWsSZ88oVLPCLSf0od
UUTIWAKiIni9JWeDHF0elgSQJ38g4IZY17G+1TOv1Zea1V12A6eeF8CUdsP20DJC
a5zrrKUy4KD/bgLxca2wwG6RRQLfbFHXQ85kZ/qFbtZTGnVbgzBoRwr8wAy1K5l7
FPRQ4b6nKwvpC16MToCTytH8WKRZdeuhmf/VDSWNlni7n5FuN97T1HEbDIPbKoGY
M4ZhRh60+w8z+1ubqyZAnex9xxf3li8PU+afEDECTjN9r3FCqj4V1JDwjH1hOWVV
eAlwb5oBt+Uz/ab1LVOnmjab2GFLda8I7a6o4Jm1BrlnfiWsSOHFtGvwfblzzJDY
6yhl4QhVwtG7vUwQ/MOptxhQZOpw02+IpEKQCXuQ9lVJCtM1R1AwnZSjO2602cu3
rCTIup5NqWwLriKW8twVnyJwuN86HGXICbMC9h1mCXPGKEORH0tyebci5YiVhLvC
zFUW/GTI4i0n3IoZ0EkUH3eqrZxfC/kSRT/4k/6TU/TR7ejg0XXfxQlUQynF5S0p
Atgs+xKjMb1sqCREIUXeLh6D3xE0Ykhp4u86+MFRvIo/l2LI6akIaj5tRgblwYrL
vDqjesvOoW7R9xYhWGW6ZmgsH4WNRzMjPpOYeJFxbKtPcibE5UdQxiBzl8v0Gdkq
SzZ4rIQMzbm5TDF9TD8CqndfvdYxk1x3AUG+0UeM9Ls4ikxhVcZVUmf2b8nviqbn
6FctBFLZkHGa13vL+P021vdQoXDNz/3IhuIutcGEg2mdzTHXJCcuv2m7e5PfT+TB
KUNq8o78yM54DxCv9dHJEZp1L93P1tnlmtUpsj0/iMdC6puT5AJZn1xsgcmYIFbP
+rruhccFOPTJxQCayn0VjKacLC0ScwD87dKUbSyGkSQqSXhGmc8OrPOXWXI4aNcw
XvTBm0EE8gyRxPK7iT64UnRuE+TVFlIlVGr3IDaOIRpq1kWa4EIErYCe/i+EvDy/
a3z4eBo+cbgwBabEgmZjajTEkuEgTVBHXcY1vCuyhARDK+rPNUApk8jPLkPGxPs4
sNVEdM4o8XMWsePQulbNYW4Fa3lG1txIv0c+/ssqiObbCJgOGo3aTOK5mPoM4xJd
rhUHGgqET6CMK4+JMTql85H0Zo9sLzCTfA1Fv7t84S+CGt4GyX5sZXLnu5apqE2H
hCShrnY365VGSVSc7ecYL6Oxjv3DmXHOlsitfkX1uamXxDEqsLqtKrx3+EXU6zzV
rPzUrHrjFOqGIfPsehfqRWrlU9c7jLLTi7sKo84lBKiTkUDTJP34/lDOFhtHKVLW
KEmp3geEttBSzWtlF/dPsrWOEdzLoIONOBM7ukxUkPCM5L4S7wjW+vBve4yr5sEG
65ibj4sAEmn8u/4D3CKzG59jFI4FqMA1ckbbM0KIA0lloUEHvNWWFuGIBS/44Ad4
uydEeQrBgKt4RjPzdcJqWjUdH98ixVVK1OP0kdjfl83Nk5LnQm262lYMuWYHlsC6
tzls6xwWDKIUI7068WJGNRNiJvT26fzCSL3lDpdnS24kgZtdN8R/IJhRSs0HOKFy
TdofuIBT0lfQg9VxDNlaw7KEdQmhsbS3w/HHR89dlzdeX0WUsOozpJgC0WAqZ5kg
DyJxg7pqhCp64idTflM02Uhi9hzwSnjYK0mjEk7areMItoSGyiWKsd8TdHcSh3Vf
2nIoQt7EpK2lGmLH31TolSRTFGcxLJG8X3+Akiu9mag2V2SvN6SIpdVyrDBIa2z8
qfeZ11OrIpGYEWBFZBRrhpXiCMxjlClR0kTCF7eG1dbnptxnugUPRigFim2ISInj
d6qXX33MtGxk2t7oNsU+2tDYVyHrhvKJlZHE4YqcKZkOCU7sHx4CYfmPmLxTE7eG
eyWO/SiUAIfkSYqsq1LgHfwV00UZTx57+NvVc3RcnIXi6y4goqSKr8upwHkGtueK
uTXAzqveDny8u6+8QHSJ/YgQZojSwoHup11+kRZWGMPM6f6Ubs7BRCKVbBu0RWiF
Obqi/eM2LwbkU5xp5UnPfmeoqFQJj4+hAz40/sbuKAihr5FdLEki9LRnxjwzo/uQ
BFZHRQqnZymemgIx4QRRO6BEFFCF5F+zdln9oWzAscSjI26dt63m5Ni0bGILd9l6
ZGUBDhSqFmLLgikscj1VD568j/lgWY9HEh50fBItdanJp79SenPsCSgFFWeq77pC
OsAAw2hyLZYsOZS2oTYBUAd0teHK2KFpkz6rtzCAjLBPP3ndq7iJevC3PjmTOObh
urtOnoRLOaB4/wGN0T9IlXf/gR/xxS9QjhqPgF5woWFlOD2bx0A9G/Z++Xusw5sF
jUo9yfI18nOY5fsIhRcLyVYF341Mfr7O36YiEONAmEk+02XQwTiaSlZr8yrGwjP1
sgD66Y95fS7KDVQzGUsQz3JyDm1DI9+6ULifLvpe9J1at9KWKPRT9ZKMHIopbZUL
emz6Ppumh4MjaoEpRNGGl6lhJ9OowgdTsYmzcd3U3vi2cCuko3mWGMSXtKtWWF/1
WmGWawXWyqQpF9VTuAnF6vMJVTD9MqwhIMvilq0sszXW9sYgK363rjPNoQgNrDEh
pZs86mwWsMMw5Ar3gT7IHddv0C6XtNtXz4I/OZoI9/qt+ZojzDVD9OnXO8P5XcY9
Yu1ErPIUSeq1lsiEl0pvx27vD5SC5XK3gvG946N/64C/1/flJx0Vml/UebPhsJmw
cUib+7dfGzO2dQIct5zEbQyTYK6f50MYyoVjq3vVgRdqXa7h92HYD0gNerFus2j9
oK+C0wdw2huta7WJVZLwpeXx+KGb4UjHbpb77bTASGrrhrzQ47d9dcIebpwuoO8B
lO0SDmQGB6FtbKoARZUqug6MUM0zCrEaQbklY/PWxSb7N0T/8hq6LuYgSs6dXki2
BqOsFtxxr/J0vZG3N+/g8Bc46lRNcDh0yrWco80LDhCnSWeSbj6riO4ZeVIQAI6w
7iFCbioVk/ZygMREnu9cVC4qSnK4uiLdButqb3EbD8AsV7DAizFeGLklFtN3GCc6
PNRYgXuYo5UXNUVQ1UXVXBBx2w9vPyvLyPxAS80jPm8WQpc7umYqFcTdS0g86x41
bHQssxinxwdwQJej5Y9x+gDfUERrXQ7jPQu0zBJ19M4hHyHAXcgiYyQpanU7Wjku
lBm7YSSqeeMbCPeHdNg/HTqqaOC9GxGiwS3zU/1EGfmNwvoD6xGxVhCwRXVLQu4J
yQJ9vhr+JCaYXRtBhVHob0WvHSDZO9i8RhHpTUs2yKbBcgHGg4S+Ou6R9Qn4+9iR
2McXB/dYka2UaWOpAwA7FsWviba6WE958JVgzYJXUWg/g+scGJF4BLtLQytJhJ6g
WV61NlWCywzRsvECNSgc/p3xiSvRGYbK/Vliwn2OpllByMocqTi16DQ6gQIftdSZ
h7kUMXJBfVGpWBBl+POQKXTYlcoATXlhjaWsezxLQW/yyrNk3KMvYpWECnzIu/S/
l1vh09SAh0xU65+SHzL3mogzcqNVlkfnTYvyuq9j/M80OGJu0TG1suM5zp5krGRO
bPRihe+/SRgoMpFqgxiNFDpWj4Wk9fQj7ibEfi9J5/eFpyq/wjOK4oDqNntMZS+7
LVq/GSkno/RbD8AhM9rezgPI93Cvm3bvW0EoWX5cvrxxsDQlLTcg/mHVMUwR1Y5C
KF7SP40yzCHduHy1zRQ4zTS9H1SamTYoI2Jq74EO8WaSokOFLmP/6Nrk2rI+F4d1
cHki2nAS0QnSwvGPACr80J46MO+H2j3QEOH6+mkLLVfiGmQ2PGkVOF+hNDAHmWjb
yVyALb9CCMGQuw+fQlr3v6Gw5t1PZ5IXvsiTPZW6yBbAN7UpoMCT24jUX0r029iu
0OJ27l102KbRsTlKRqK2A+c9Poyg/5fEw03RX8pgKc/nFJsLYqoNxZ8mHpJhmPe8
NyxwknqJZO9bxWO7DHpYETWvWACgOBVH4RAnbTeiPqcPGiMoJl8irlJSMmmJQ3cD
HIN7zWjifdZypWpbMvYdYZyaz6ThVukC71/emPryBA/zH7VuWz8Y+WMyog/5FbaO
o0MdEj41WRwug/+2BL3GLYMZ9emgnLNb0WV5NWM5OkbJ4tkvTISff0XQP/WrLvmR
JEWArikgy0DK3qs1k+xWrJZsO4E3TYkKKz+VGzNXIsy4bXh8xDt3nVJhiNavoQBK
/jgpUdH6AcqCYYDtf/euG2YlZIgQoLV0w0SwxIMY94F5ItxEzc4l1jiLOAQFKGaI
DLLSH/+F/LZ5+hK5LVeITbHz8ePkxjPzFoeSkqyWPctavIxVVeqxSTiC6ag2gmD8
3n+oY2W3FMzU2FALzmcnGOyCMvcQ/66NTLIHZmWz87IzU8X6Y5AuR9Dz7dF8Mvel
WVKZTd/OUU0QXKBL/0wzrUZVoM96VeOBGj27DYL/L4D5rlKvpOO9MlsrrBx17jYM
znguMgeMXJW2qR1g3G+w5VWpu3YSXxwAfPTBlyQqX2omuwvcjyeoK+D2L1YxY07U
EfASLYXRkO+KlaX3VJ/tgnk7S2LCWO0ofkSSQY+YG9mqK+YltwBlYasnFKK+NBDf
ROg0fYaSXQ7LERjjXijBDh49uDmW1FEI8j08xPB6qaDwhjROvgLl8ACMe4awkVFh
4FSKMKC+cSigyyqISs5ZHd7MA/WFRKyv7QeX2EenmCnnhKzuZC1gZvrFO/K/WB4m
dkXxQSQl61ESJuuAqP5ZaWpo1LBlcXeoiyGdmZBgHciOyrkHC+YstS8NxMwx4e58
qsIioB11h8aBlQEaF+7xN539/0tuWI/+MmzUfNDy+ARvx0CSSh+U6WfY1YRgmAgw
TqtnxK1fl+SxE97Lm3E+XSJ82g0PxNs5u/S96f7I8JuJNZ/Sc8n8STdSa+J/D32K
0iTkA7lvtSZ5DjrqX1WQvMwz2ktxCWKmRFnZ/ZHzZl2FsXncUMVfsZ+oVXn28hiG
YEe5jtYNzYqI0CWVJegfNkqA0K270+wHr/PXl5iKd3Bnl8Ac/FfdTFLkshZZADfM
jjOhLwwfKJeXqqst2sXt0CyundIQYJX2st7NEONdE0Tb5FQVsWJs231i9/kH/omh
3rQ+cI229N07vzofneseb5G5KW3UWBWe9VUjdM/mAnpNzk87oJ59oVuDd1upHZrb
O1kpdX/I1fRv555gm5YtzZRd9PEeihY6g1y/6uJrEffJOQ08uq5xNACLeNMHeXIO
ekz8STMubl9w6rAGSXdSaIlUUPZsg4zR9mXb9bKRUkcVKmmxZJTcgBEuHw4Yw1Qq
ekyzFOI9icr4U+RL5ZjG+RIvXTLAINC7++qSPx7OO4ty3MmVvYB2IWxy6WEIEMNe
S3XuC0ktkjLEKg50ZtXYSqA4Nn7ppUsxNGrg83i1BNX8zKSANwFLxV7OIIVRmYcA
EjL/fO2/Jl8UeLvfRDMuqY5bBQm/xsfuu6NVzKIL7KHe628/YDgipLvn/cv6oh7f
8fVAvqaduN5DHVAPReLv+ZBk/J8pEZxUmd2v0HHM0g8iOgln//dVPui5k6XGPiLN
cjQIo0Eah99azlC2AmJ9KgVbwnyD8YPMybC/6TQ5tHKPrBM8tsWmfaTj0emYGnMA
hGcdat0VlAx9I0KAVqFeVA6jKXvqumbcqd5nfFS4/Sx1wf12c8xIvUH4byQQhG3r
u+B3LW7CErK5fMqvHFSuagZ/UBTLmo03QWIapFk4+48BfVLlXNltGwiW7nwEoZy2
JuviAE4CP8h+xS7+uIxk3Q1Q5Rhn1aE1vwTIFXSipttjxsU+FaUqTrcaS+m/J0RT
fv0S7cHNNTB6gOh3+2AXU57w2ymwZMJIfAJO8CbtLr7ZdJyQFe9iEQkCLPpzYQef
DIBPdj/sAGnheYdV7xwrxvKYT9aXlbnPCjzFv19jG/cd2uAy9YdfO2CnsQ/9iLWI
3HNdjiqG3dWxR6qjS16JnEi8uJkXRFlBBQvAV2e/38KeOGt91hgWCAxrviwHJXyK
neWLCEedttaq8znn3PLb0labi069BWSPAS2FFtNXYTt8PMloEz3/RbqeOg47SGbF
ngetCxaDjufgDmvFXaNEiKfgGO0sMKi9UVrSklHapjRaG76s/Dxkwe7Pv4qHtHj2
zSqI/Dgr0kZqMaCHtEdu17RLuKyPGbz2A9ysHHxWjt91jvIsBoHytKxQ2w12zhp6
Lv9/rV1e8vvNdiD/ddqgigJWvrgCqih1yytHugKET1BBMWkn56yKS8+40Dv1NGpA
VNpt8ADxQaoRKco5z0s67gNkbF0qbHGFskf2A/gKco2G7L2NVAxJhLXvogotLhsX
1RDSVJS4H326MWfPhOggfzEYAaKNyRoXhzlW6Z5U0WivUWBh+WF5VgBLaHsucXre
V3kleWdT4TdK89IoCH5xi7hxI6EQ34NXU5nl9hPPK7TvkhewPhc63z1g7YG0sCQd
kdsWQtJYoQG8peBnh9zZZaEdR/GYFLm1FfGyr6jss538IqdJ06ysmysFDK6ZFjQc
uqFEk/Zt+bv5KOSqRYOskLPUtULBtR2MbCUIwBsCUi0E41qpISf+15S7LKk9f+iN
jIUXA2ldv7SJWYLc/hcAA8k1tKiV31/GyVjYSMTxg5S9Pr9pmHu5RwkWqhpkOhrH
vKzs3KwPEF8+VmnzS2bXLIqa9y3P/zpYc/ymrd3+OkQgxysyMigHbEgVwoEzKoFA
JL5/lDgUP6RB5zjXPrVNm/JWrzQ0rae4xiGaGu207bSFNOMsP8Y2iIVK8jXPkVYR
pliMBHKPz4tGdYqlvUeV+XDVZ/seJsypf++ZrkYkt7/84kEe9pGK5nEYZT2yIH5b
dPveMUZBiqHU4gij38Hgpes5D/qcG/6x/hc7xYHy0NeIrRY/onfypZ3qDdisJkN2
r7vVsKWbeZLLU1Xn8z0rH8hpw1IngwMxTgxoOWtD3C0MjiNC7x7Af+qrym1Gk7Mj
fNlnNZ/tlKBuowcXkqkDkZiHOXUGJ6J1oZmMMSK4D9oHmB7ggxOZp2hkm3UZMwqB
uAsx3juV1iD6c4KB9tZ7SwwM4LkOMxsfFZSMeyOS6R7X/u/xwN1GXQV/12EoT0fZ
JtL/tUeZyd4k3MJ/Xtf9xl5EHvJ1bfOUyWp4SQyWZ5mo4gjs769midoNvKm8R6d4
HeVMByiz4kBTWV7rojsKrudfVktfxttm5ovTOJjH7xNDGuddLDq628S0zM7hSuYs
DCG14hDyC4uiNta+KGzhkCv5WX62HOj7eATy6Nm1uOuwTv70JiyMSUFETZRVJ8mF
+0Om8ZfEe9PpvZC10nPygIiKgaDCQmoO4HjUGLpRQszNb0UsI7xSdMO4xQbr5TuI
+zfI4QPcjVnXDLR+j77UFfe3iLyY+Imn9W9lW5psuC7fo/gGp2DiKvGgBZyejvki
J90E3LcF5hLDBsBpwBM5hycLO2jHiInwbZcdBLXd0srM+qI3QQ5HGQ3tMXOXeqK7
Fta2ddtyHoha5F1TtOn2MEVB9A5Q3W8jvzHlLr6qQ8D7tXtb+H/yLmZ8LfVXwrhQ
vRlOg5KS12Lq1VZrNc2Ghsf+JRcioJU/p1enCKFW/+lhg1TeNvg106TRgkRo9HBH
jhXLmPXT3vd5C4lE0IljEbrtbTlzZbK9gFCFp6icniOFgcTcQX0NeSdPu1BC8r2T
MfeP8zcA8Djy2wSTXPziho9XHp8JfDgCDjmak+WIlxrS/gaycPdQjPiqwS9ExI3p
/stij7JHXnINRGkDYexna8TW5223+wLCVhQtZN+798qhGBSrgEmdXxACNjeII1H1
+9Ph8BAOG6XNAvqv0fSsuzgJ78bXa4iVcuZS8krJ5nP4Sd+Yxnq8jpJ7Dwll+pF8
OFCXKL0utNbswhkYkfpEZa9zEWD7hTy/gBciOnGNfGBuS3wHS/o7v2pZiZhFvIrg
TTTfSCX1TJ+K92u0hUVqpBd8ibBeu5qNi9YZHL4iMe13sTW54JseS7auQqV8ikio
wah1TkTA/w5u6TFkdbHS7/fnTX4BZlR5fRb+XprVDJS7mOHFhUCbtowTRcSrNvdD
Z21pWvoDGM+E1oOLxaBr634GVQcA7rZpEJmXSbhYUbScjoztfXmHpEgisKADWDQK
3HqgOYqHnwRABhSdJ6Z+zMUYdkEOPFwQA24RcQC5ejAy73lwLvCQ/Qbp+IMtTyJq
EBYe77c89emwrybHqpp2rEx+BG9/NJCyBEFgTdYITVApIj8gGR46UtkMMTE+eys1
qJx/nfxvdv8khb18TtusHcsJfnkVF8sNdoFW6KBzljQz0qOjLcFi6OzsWfyYzijv
gk98aSPU8bo8Y2S1VQgzEtr43m05yMs35eCD1wQzORBJSVC8mbuEIz1EQtwE0jlN
odD4p4Qi1uZlRGkm9IPoqrnxJR5MHy2YE4mQUU9kjBlt6nBDHrYPNVvK5sse9MRd
FUW5PaVb6sKFETTYRJiRV7rbiQnTzzk/YxvXvwVUoXoINscq/PldvwZwQDn6tICO
6szEcYvaG7oYpbM8XajCA4NOaoHzPNq5ZMFjSKaTMj6fBugq/YM9vfeRig5PM/b3
oT3pwqxQ6knnNkxH5mYnQcNyomzczAkDkLcB411MUovVHPwzIDXmMr4rl8TrCucW
WxkF9pS5tUcneOAFIJ7LPYrKp2uGrtsK5T8cfIgIQqcgFX2CBM2JtwOQHmQsNEUS
T9/bGIoS4f/KqFIYDjgh2SIhZbm8Day4tIp7Q3TmUJMkebwIWlqDar+MA8oIV4nu
HM2r/HKOaZZaZiUEjmbU6yOBDI4OOBZHVYkWQQg2gFwGAIMY/xF62foVW4rSiskU
qzjfr1m3ysd01NyyC8KmcksR2nNDzc90VRDy5n37teNirRFDVXHDlE3YmP/YzYGo
YroEJw7aAPnEZ7+AaSMSwXBUjErhVnhkvacU9Imurwte1Atr2eKvfeOROs00po5x
kwmlbhUfB5xZEffNNBAHKQa3B1bvTPf7ipyrCP5EwfdpLgHlnwBlNDAwByXvW6CL
SdBVRHiKF87IG21sifAj9OzenWSKYXQNsL1R/jGfKcJOBgrSnmoD4odsEyyfpGEg
2sP5gK65ICQwx6K2nqkFRrYfpkXuHfEOZZ6T0G2Nbm2QMvECtUP3Z2gQ+od19Lxa
txhGn1X7nbqjDfN9VZf4ae764VWFNxDSJziySpve+WDjiSnaCdX47zkCcDLJ/HGh
CeRR8BLnTgiCmhCflogt2k7osV1NOK3qfbc/rDFstwaCaInOOpzkXu2L0S/BPKwn
05BMcktH9vMmaueRItCtw1y0sqRPGwULt+HWD85o1mweoQcAYpckzvewbmR5xvzh
m8UEu4L4X/Jl2A6dWoRCYiV8L72MjUU3boJF6AupKPBepG/adZV8tqdFD3n6YaK4
L0Da9AhZkk901hHLv0KyYYk6QWoswhPG4qcfy8mkxifPsw8UKjfs5102eoiHdTLY
O09JNjlGGIlzWLB9Bqr/giR1mdXsdohTBH0Pnn23rbTKyC/fiweigVHw4FzqDuEU
Nxz9wipc5gK25wChOGAGDRNq7h7Shk6IP8yOQbqrujvQ/3CL8pRkuVunvSt/AhEr
/bvf1iBUw4Tf4MpSddXSRUvzCeXJQ1kK9Gd76uebijTHFFz21S4ZDbGCBjmE73vF
yPq0z6T/cDwHX3pM5QWszdsm7JJJxTJjsNbYz+bhsmDJwxg8gVjfryUWAnQuqL2X
ggA7SJFGf98OwNNrUjumAGS9Vq53b5eFRXaZfC+QcpHVCcz0JxWaH7RPCkQinkvY
fxoEZL4tEDzeIAdG3DLK4aBVMNxYe5F1VyEzwj52/BZ21280RjympNiWluYIdgIE
l90Uwn4fUtAQsG8BCKycc0ckE3JXyjTcFKBb7RdbE16GfdlVi0p2i4iaFHD/ub1j
ar1KaXu096vuWhQqazwp9UnTW2t621JhTBKyeJvj3drj5w0FnPy/cpQa3/HRO8rN
vNQMyrNQr68e/VYUNtGt00THMCDe1ojDeECkWUboCT6X8k0ul/yLlClgGb8gaXIv
Hh7UyV6T43S5ms48goqwF/+ZGnDPfZaC/A9gE/Zq9I+1WB8m5wSEHl6j0JNOxxa4
KBoXmhTAF1AincI+ecvBCLJ/zvXiootDMcakngQTWVxs3pYp4Zjd6t1Ao7+mUBJN
oVlG8k56Y7BHbQRCc/AKHH5POIHvASmUXuYXgHnP+szC3JnmYmle+exsrlmxEvmw
72IS9BFTgqSe4yVT0W+LbEux+vWAt/0tlNyQMMav1MSCT7OEAwHcXKKCw4+uupcX
TLzkrIfedC1VHG80MT0/UtVr/0KegnAk4rS0LgCWKidVJQ8EoeEXzgqFwBb1Ow4l
pm6Dmd9sxZ74v0jD8WLPzgeWgwA6CuvpKHNNeJeuC/sqrV1V3au1x/GfAQzE2q/2
IUt48M0cbyhqm5sWIOqZeMhH1Anw+M3YDQmo+wIQ7ag7nhRCeT2wDRuMrbW/8Hab
+D+qaG9KRtFrihLYhmGrrcSxTjiFD4XegoxIpO8o6KAnbVS5HwPZuhi+t30VBRq/
/F5piTL6iKdCUq5Hsn0lh+X3R0cQAP9DkAI8NsthvnmsrK21YFTRJ8W03Qu4NmNj
akgwAbgqFJfJSnnxH4Esazbwriz39Q1FEs+y8XToWh3EVmj8hmhRsRIYU6GlhKAD
oV5MIuZxDIfyM4tQq1YiRB3yPKYiwSCQL3rmqKZOKXkf+pv2Nj/k9waSGrrO+IyZ
Lfzei99aIQH7MTW1kEABIr9QtFfQuxqpYiR+hKNiFsJisgA++dUIHHxNxiVP0/5+
Zza243Gq43Zm96o5liEX/k1rG+1k0djZQDYk8ympAnFa4l97MjwfMWKxlLPWtSG7
YUGYwz1sl5Veqc9lz/8sS3qSqSKfBZiEvf8BIR2uuRj4QvM8mIIQxLm9YqcIbXTV
pwChCjIeG4vjXaDAs8qsTHkJHql/hIRsrlv/QHdL9ybJKi4AKC9U1NvTU8wNh6W7
frLK5a98mh5OzVjD3W6f/QfOh11bZlX0f3tTPPMeP2Ly1jBvLMdUPb8w+u8Xafbx
GYmcb3E8FTFSb/tf5tSZQ3oZ7rr3NLPJOEKVvJRegkTrPw+rG685+ejp0QK0delF
MD4RM2q7YxYcV1+WiOcWb8lwCUZ3NxNmlh/RO/tBfnW04sSdx7v7kKZnc98c7o/e
CH72scx4n3Kp8MrVyaCXOjQNhr35dqf3k8pHge9rYzfzcRB0b3XHKJjaQIvY5uP8
xtGNcpjFCC2cRCOb/E0tQs2wHcAMxoJMPuAFPXwp4GYICSWgO8TaSnlbmZUUfW55
jbySJWT7wf03hi7eB2QA7iGYcNI5nTogwD3isarcGdlomPMzi0r9GJGeJwqa7qTf
4SHiCNGkCQy41WasPmCW3VNFfcs4Ue3XtXr4UeCeNxdgDtOd+hW1TEMQ7aQpoqLU
Xz3rZutzgqxUBsg3qDfPT9QTf9UV9RK9bW91OXv1A5faAckVmKo4RPO7E93Wv6D9
rPkqXWqqelg2fPx+fLBKxERc/3L/TZ/hKLZDKTF4ytHU2aHuNMmkxbVuI8Iz2i9o
rPS3Y2eK7WQBdn9UPK1/o0KRlEVk9pgT3AQwJlkNXfTtiaM+zJkNstOLq2jvf5IY
5BsH5C0cxfTVI9SSau361WwmHzPRaml/H0yYzSlOVABqMoEpnveu75Q7vma6MhTj
oGx0TUIYtLWlkrkza2fsChxWITkRKCijHb9h5St6ggpnAVZv+/JSRlKMPQkLRD4z
1f9eVM1GUF0q9CqUOLcDiNuXvI2Xk+f0X+MdTq5YzxM7EFSg8TD4ic4LQVf5aLIf
+QT4wBpUGa21usqECCTPim3sOmo4fxGsH+ptwtLTbJFyi7rd2+FwcLZ8OGZiKimK
s6bHyaU+HLMIbk2T9ZWc6BeiI9uhwSCCHaRPJCmtYrPLnpCfZx5ZUnBnBXzvbGcJ
dsSPCorqHjOibB78PVn64/Ny7/KidVIOL0okTPixQJNCnwOeYLWEDDKMJ2bvZH8f
s0V6L9jPJgEN6ohW0aZUOYj6AOVSaa7HepKWKHuxjr/ZYdiCV0zCSzSSBpSTHpU1
lD1xuozN2n+HD75yvF4WpublKsiqrkbnkSM6dsg4C0yy3X4ttVlpNnKoTv+nexvl
TLaQfEf4IUoVRhVkSauVvlDb6qNhYPkYpGYNycBimlANGg6A1NKy0biUGnLul24q
52qDIPL50C/F678EHS4Lha6qs5zMxyOCw2WQJmbrmTfcK6OE1rO74hhH0xHWJkys
6LLwSApKnksWllpTsbdKtvy7w0JWo9bEuKq5E2jtjABoI1VPYJWb8x0+QcqvmFBF
yERs5Omr1W7g3y//L/0XfpqVAYtE/K0MCCEpuMgcVhirPFyYL5ZrUNVr9BiATNL1
/NJ2T1LgFjWE6J/0fbnBbbwK8E3tSZWqSuXEXPWGx5IWBjXqCUbhNmF+2K620e7g
44K9bGTbqTK4aprp7g7JrwrgwYpEhd50l+zS1MQNEn6CKOhT83LOaeZCZH+tuUpY
xw+P+Z8cOafgZYmmbwpIdLslnnlzBucMqCDmbBmi6peZQsZoTplD9JaZooiyRf23
EpjyGYV7mQgs506TavdKDzEkfiIqy3us4yDLw4dCHKK5/4g1V2x8dKD/2of4Bj/y
SXS8U48vI4V0p+fmr/ZFHYsb7Bwgv554Zx3tpe3w8pe9DumXRKTeZPdQOmRS6JuR
UGR0rpl6Xeik4g/GDzRXI4abr+zf0OkY+gPrnOXpGzsDxyZQtwHMoWxiacI/sIEk
QyxDgW9Gm4hBrAk7HWtGjpW7fxyMG/NAcAsigRBtrYWRx3G/TwG1MAOZF/mD+H6A
tm5dFc0P40SHmjOXs5RGkkB4hhWqHO7YwO8M0uyhPlbipvXzxtPwCsupmDPmsmjS
uh2ag3WYRM377RjFZCNFBl/7JK/o8p78LiQtcqm3GBCNP4QhFzAqjJ67ifPLkQSk
7zWTZuD0fQZSw7ya/tH5D9WfCXbbj1fMBK0HsXD9Q/RS8rKRd9zte9xXL23ydAlE
l6rlhLadE4ln1u8wsRvYBbYdKwvTisyjhKpgpyEYHbDDZw2cyqyOs77ZYWni7YDR
0PxowKg3+rZuTtG6ckdFpd21uz2KOCQLhgRAzbdUZydFBSBvTQPG8BzS+DZAnIOq
kxhecWkg6xtHdlVUfjRQ1LoUIMDc48f9CdTBXR5MP7XXRaIOPy+n4gPCQjFkVYqj
wUhO/QTPxj7G9oxaLvyj2bvxl0xA+aYYIPtldoad+xyhicdAelnK9r04XKChqZwV
TdGqJTqh8l4QOaUPVJN7pnPH9A+mGGNCOrlR0MiS5LDhjv2KuqQrj3doNY9/L93/
hW6luFPskNfdalmdbUZdmkQfT1TOa9Dvyf5Fw6XSBuW4QD2DjFHcR4RHDKn2CcgR
qVSI9JEnPPlZ4zkHrj6H5f/aXYcaeO9RRRj02GJU1x2MxASq0XlLNyzDPcBkopTq
5VuDgA8E8gz5sy6eMnuvWm9ZrFBJtwW1O1DXbyMHcm+ofLLC62FTX2H4C9hEY2XK
i0UzoWde6jnz/ePtI0F/cghHV7lk9natdJBvLGJD7jYoG5DiXl4BDSWlc+MSkNDn
CvyQznfszOL+45W9HCcthdZ/x7nhxkxiwMDGfRQ8Nn//k7hmdIPFAIeqr2nvF72o
3GWphYjuwFxoWcRA8UnRq/oAhduvXn3SX+F2CcJ/cOnizZZiSNHfw18nABXtDt0/
UgNcmQCkQkJK4SQVbRiOmOEWAl624cxSA3fe8Hd27tqRlA0tIQqPcx5PnqtqEY7A
K1h16Vkjb6ZYIZ0DIW4sYGmi65gXhr7KyA7iV6IEY1ZUBaqpkhkxvzfuBwcOTkm/
+h32hl4no+2RKirs2wgmSM3OPbjliwFAVAe9ofs+uxdRkwwTzuBs5DGqsb7nq3hL
NkbkQm85xZpM1pSekvZZ+Z97WhHgc4oKB2653Yz60a1m7eAizn1dC6/oX5orCKR5
GmKl59cfhpdbKQyvqYEakGrLv5i2PFSklPXgTCLbgUrG0DmiIlLdciUqc6mIrLNB
uY6a+Hqq2RS6OIqR0Nr/JHDXq4596r3FhDbmdPxE1mVMTzTcgAlk8yR9GvYgC9pn
9ZukM2CGx+gBH0ooYozm/B/4SyOeO+U4zpamRQJEceiFoT7btOX0VmXbU2mb7782
7HLCZDvf6nQRNcyl1N83uyeYrpo5NtlTpMzNDLzugCMtpnPozkw81pFryHgF93Jg
QZyftUPk+fR3hVF2JDOJayc+0K3yo02Ckw1b3jXeN3wNfaBaWkm4g/SguemawfRH
xT5XdtNn2kh7dvHLEA/kySsV8SwxNbuI7CnFwQasdFpKfECCZRLtH8639cN+RjAv
KkkXp7vzHnHzMpKtm03tb9AT9QfMsjGnxOTPyBKo7BPFdUSD0Cy8dX6MLiZzLggj
+6FS0FV9x4VCxWZQr7CnMil+iWCgv0XDt3pEFSu5rzukDXt8vTvQrCIlVQfWxXYz
vDH24rb4u4NfDXat7IgKDHFJjoLbETAPPdO3Me9wzxr+ZJRek48jjT7HyBl6lNvV
9ZY7Iq2qF6w9tPTl5ZhfkzD7CzvNgioWvfrT620H42+bX5w3GRJjnnVl32liFfH0
siD8rhuF+px6zn96eCibEre1GyEnjrr5vvN57VgbzcK3qaNe7uAT2GTEgVIbjnTs
G6F/Vk2rfsxobfqEv1rpdoxtEynFTVLBdo3SbAkjlG0abBseZKGEY8x5H/SIXOV5
kzxrd3g/ffmm3E+uNxNd7WZ26FLSAfLe1UYLAees5VghE/AbiAtL0s2jMhdqS+8A
fvF8Ud23BVTsiA6Qz00fA01y3gcdWxJrqg54CcFKZHAjnnurW5O6sSUYtTHh7QE+
s8Un0SiBIa8nTxGpCUPGBb7n3CUN12cNvz1984fUdqEDi0dK3T/xne8qBCPS/jdE
PIy6P2cmU8FQtHLByl6BXE+VIv+0A/1vBwhoDllm/EV8A4Srtfu8MjxGj/MjKw0Z
6wNlaAUfjyxD34wMeZ2GctRNazB5//PhSePtQ43CL6bb4Upc2q9EgjwEH+1SRQDN
UY/98KZD9HTR7ROr9udAZ6O2/u7Jt7YSUkfZ5+ffQsDkcJPiPnITKXTTrP2nW0Lh
bfGejBPV2/xMYIgxibycPdqVk7HndcogVNmLj7S6G1hPmKxI0tIVIbjVDUzLNfkg
ms9B63eFH0NAiLr8CJFizSSMyjNoZ2CQC4YU8VZh3/Huc6xdpPVGRAbAjf1x8Fc5
rgk/tpEwq43ZJvG7P1gGJKm3MRNS9h01YUF75F+GEcjp7K0s8Z7ThLULowvK3+hS
MMvPtAwNqPThFGEG/+htSpimWcCD+p8jBtaaQTxxLWKyCalHX9fEaiZ6krhNo+GC
1IOGZ5OmHzGIzmjKmFDqe6j/Qsu9aY3sq0CQmsU61XV/U1gd8c+7H8HoOlP/slfY
AZe/PSATGyMC+KLBhpsCcONJDWiQiT8bIqkOZWwh+tdrb1eQwMXBAIoNSwtkHrMG
DH01BUZefciiVGCnI4y7s6uTsfHhDQe/QhMBoc9USWKcsYYHa9IaVhUohURXYCS2
NMgGAnrbzxNI1D+71gy1Cb+lXPGSYH4NW4KRyFZndmtFi76vrl3o/YMx2qwjOXME
lsKzrBwHQ/WBsC4nTVse2uG/swBGjDEh/8mTAGiMMfxy9QCrIWx5yOsGZRb3PCm/
wNkVUATg4B+efJtmWiu9wpHHYiEULaqH1+K2N9JLF9Ms08uuQB78ol9DOeozaCW0
nyQdB+A05ggNU1OVP6Uci2J9T6djBJ1u+SMmAKS7TvZ6WyLqxojpDQmusBjLlfEc
1qLCVcZvCGx4qGzLp5lGf8fSWe/KLcUzb5WeFIWhsqMMA5KyuSa9FZeAAXFG+zqr
NpHrVWhIMgGcK9Mdm8qFWJAadqaWe+eYnPALF/gpf+msEssmF3AgIki7WGrr63CG
gLFFyLeoQTwCGx5GXPXm2QrKPp+a29v2xkA4Ys8FqAO3owsv3rIZQfbXv/2Weaz5
7yEUG7rcfrcTf0YhYUEzrc7A9h5vXdGrNV96jvmFR7Dsv6kT0dReprdora/vjH/J
nEi5KvsJgdz/IOfu5djcAc6G48LHU2M5U2zKc9Elg1yiAkU/eFyIxSgWSFPQLnFc
v/GyJ0woBgWq2UUeSo8pGtKRa9Cad7iBwS/lYwK7yTunoO8vazUQk9drMm4afYbg
Sub8uLdSfGK8i45FHIT+jmF4EcgGAxcP/gSTBXMQwfdiJIxgtvz68V1GEVfsD4kn
SIpFblTBtmJKVrJ4knWzqLC4sbfUX9ODAdBzO3+BVps/OTwc55AvEWlqd2klTj4p
pudVOrP2MNvEPAxyRYw4n6PEhp1dmo10DdcqTToGq7EvcLvx68B70grNWA0Wdrfw
r7w7NkI2NEFXDXv0Szm5Pkd6FK16EznQAjllAB7UVdMmXzOxINDOmPG5/9FyAWL5
01eAHBgOzlsD1fsHdmmBtdBFEu9W2yYjQNV6Jq7R3oKcDq2X/YrGfvwEJ81/+IMy
FvSsH0R9zmfzH6zj44sd5Gyco2O+WDh5+63C6psnU0xe17tpFJNIiI2u4NuC/3hm
jAr0Vt0Q0EvL3j+0XfB2STBojBiydQzf80tDBM2BZdXVwLElNS3eC4JkOrN11hkj
zhZcAKwEzqf7Fu2nMsfiKTIArPwNFIN2cZyrVSLlkB01dxG3g43bnnYKrp06lGWp
YUb3Q6WxWPObUJodYz+RrwFjy3nCG2kvJQQQld5T9wXpd4gFxo/oBuweKnZYgtKy
U1fzqTZXa6S+DCn4oIwQ7++9wCbaMnAG0WqA4Z4QqTuFF/WlZbPaeufmdjobxOEt
EMiDSBOW3/BvLaPG0VuBZoeGkUp2gro5DgSfW33hei7HHrVu8Ks04Jm6WZYfrtfk
gw//TL8NCpmHmEEWor+yPKsDr6daOUH/QzWAJylCKUU13naicdpldVWKzSWdBfXy
25TZfEdFs3hU8b6XCQwnjUG8/Kaoo2q4VkdSdXAGawRIiuUE7XlSIXANccjVz6Sj
v3/w4i55Emj0Nkn1drvJfCKOrScEa8Gw5IkJZIgay4B1iQU7pukcn29V8PTIePAW
u3J4EEgalFqRkYRdIDNE7rNICg2ZZPPwY6tOOCv2cP1oWU7AdVL5fRifNh2tCIvG
PjOczMDD+KDyKdE0gM4mzbGwb+vUUiRueIcrvgEJL0FZMGXFkDlWh/GlerhdP9Ss
W7K0ltGryEowHIMYHIqfC0EdNKNGOAw2zJn/1W5FngobtQc1cSyfSmbX0xFvGsdW
q1nPmr+Axrz76bNV4stKEdeM1hRr8SNmFuYepkA5rjtUX8d2GK2nv7zj5YlNOhRi
6tpyuX0l+1C6rHX5rc7B0ms2vEZMPSTW8mrTgSN5ZIF9P5/Wjs98YZvOR12+Rslx
qwkUSfN5ElSU4gZzZDhVHrmYuKaQXGteicnkkL/WfiaGY3mj3mXMvWb7IjwUoBhs
k3+TequcMeCUdoBF+OZA0dfULBtcINy4ShpBc0WGvkng2wKvnG5dfMLsGd1PS9za
XGXLHlKl+9gdGkOGoi75pDUMFYRxGdhOFSHwgcV3UBHYcAnOHyo6vjg571OjDFOh
Yc5Lm1VRtuaT5KoS22y0FH5bpfnxeFJA+2m1YUl/p3YlYuPaqAiJRHnESXk4MoQP
pYAQoucziSeiTkXEu2KPQ5HTPUL9ydCNqMiuZ9+kGZzl6s0/V5OPp8zrOUPUdpzv
pPBsTwpsUtCiYr6N0+5ImaBRj0F8zHlV7BuCHJveaBoYhfnFUE6Ij3guzH5n8eIv
6+7zwMgCaln2j9rvGbRgExKO5ehSdIX8TD5hNhjaL36WbMAEWvNIJzQsZFyvzsbO
CFknVwN8MCXHMiVF/Jn+jtnnBXVzMSUNiAM38txdUk5ougnPk3hQf8G6Te5uJHBt
B+9aEgIPtvh/MGhB+c5OHsvdc5fNeIbHiyVh7oGwijK2GTZnS05c/IbzBNb41EA6
IjM8WgSxc1i0HrpZuTh1M69BE/8SkXOBwIUdJKwRTpR5cNGyUMTFv5cilUA+HXQH
eB0p0V06Uxs8NbUF4Dc/fav7v1/yxqoOdjC/KFYtIXzEohfCFzPVdKJwwU1qRzbF
zfiadY82dFEYPGQJVFAFkB9GQ7aC8GvwwvLxLD32ik3y6UQE5F145/zpmO8JG1gr
kSr9K50cD69g/TduT+fJ5QQoL0nSjfpk4F2BFxu05mvqWrco3OlVCnNG/9mF7363
RbE8Qyj76RyKn88u6SPS2dG2MsiwsXHVX37S09t3e/FYfbV6d+0+rfaINP+qUXZW
fCgycwW+p2PBeWQIrRnIREOI5G4hmBIR/o/Yh4gKWWkhgwlnPcb3uKiW7MaGIBBQ
DJBBPGlEXU9YOt+Ef1Iw8/jc3fmDA6gsqc5qAY4iTlGSPTKpTJBk8M7ApB7bvJ9G
+xvgwFH+WDprpNmhLE5PQxAoVLN+TGa9vQUBNIj4WtlJu+yugn+jayMBSmnw95oT
lnn4iAcBzk1mCCTYmP9PNBY5jU76F9wO/wV81DmXOdoIwqMhyWadNhZrM8xPLWLw
3/a1A69e7ebO8L+MfQEXMN3JW9/eajKXk+X5vZ1MePgOyGnCZTAj4tIMwCT/P9NK
ZUh85Z4VnbyfYX77H9yflv2rP6prXbgzY5XKYehXZFW2mF+1TP9uHXc7+KFa0wIj
fdKq8P2WYOUdHOLPsVWiulHl8P7vnHoL9/gofqoZihNufxSLdoHqF6ZJMpDT0PWg
NW6Y14PDDi5nUQyzO5OiflgeRfUk06Dux/qS+amxOcE5c7yZ1posVb7W/Ds/HIUm
PjabsoM0SIIuUxeQ2SWkSnZiCSW91+ey4zFFTJonnr7QJTWaTJfpnwf889fLD/RZ
FDsxKuxrmckFwrIO1W1wiiWs17b0CVW2HU4WfyOyC4SrYowzwwsItzLSjLDk97Af
WCgBHGcz95yPk6IiGozRM5wO9PxCx/BxennWGJNiubj9QN5x6L5z+8hkLbj5wZUZ
e5kljaP/ozGURai3Qsf6ffMXU5gIjLcQB6VLo1uG2u/w2Xjr9nt+b3cWGkFJGCQN
sVrhEhdtESwdkRsSDdlw9VThbOMwG7N1CrR4pCVuOIrbxiyMWM+sos6iy+moje2G
KL/stcAnz2WsFRE0OtDwE/3ZMO1lX33+s5RzvtCSjBg5UEvNNeE4GLfDlka/RD2p
TaeOCNKw4DSBR3KG1CDeW7gg/naIJQ7VplCP9d9Dv3XMLwELP3AV3l3OH3Mh6j0B
ZWndn6tuZFneLMgRnpdsfuxBnGRr0qvuDHOfnevkyF6R46ZvBTmds6fsO84e0AnP
AzJWHjbRQLoVdOd23SwungUEY2K0fFEmONrPIb7Zh1EtoYENNYmCyjeUGT7xHF38
m3tkr4wXINrIh6/aulm19RHoM3m8L0iPwn2bzcqqCh77BIDeCUFkJhx/2ScV72ia
me5kbn9pwoTmsPG+mWjQpJhobUAcoptRNlFxCr/sRfsFTeKL8imGaq66oOzyIxFK
2rmgguR0WT6Lr3U5JvomMW817l9Q2EpH1dYeNh5yaTvCxIcAKSVzB0eWX7RNgJwb
go6PGrto2LAYLZPvml3A1JacZ2qIqMC3WTBPCWqJ10duNCe3DAXoAVEO9wtsAurQ
d889/NQ7N0BtLps7r8KfuvtSXlUJvFP/pWsYAjy8CEKHxi1yutk3O4tVGkDT0+/u
C4SVwKPCuN8aAxhEwSawELJhx+wEm74NfRS2GINL6QLvJGAm4T1adg1wr5d7zp1p
dsVi+kYhR56gh04+9kAcpXAMsT0ErBliJ3f9OHaBD6AhsRGlFBRg9lrNjX30rF+d
jSuwlVDex82peeOzsCVUDsJ4LJkVYQdFexmTkJ/naSb1F7jB1O23c8eHug/mq3zo
pkC/OIA0R0ebtEhKbpVj5j0GYDXbJQ4Lm50UiXx+6NfUgmfQOEDe/xOI3/4+hu+J
8JUIvgPd3F0I/vN4YAgYapOuBb6gIokqx+es+9TDWKNfbNKBBer6pjQv1BWWSit1
4dXU2xPC+pusmqcL0RXU+3m4hKTa8HSwiGAPUorgVH0/JeNxx3fP4uCmVl94kQM3
Z0jY5/+b5jbZ8hdFPXhjMxSrveK2RScRqLPISh1VnBA3zi048CRABowc4rWoVMb3
ME1TWB2m9UrI7SkocgKB3SSLHE+FaaygssSvrqBJJ2Uv6qB8IVSc3yJu0qdAA18z
Lo4zEHh9CiaNgaObRnRiZMlkNY64KvxTBgLuOPh736/DUDWfe6dxQlHIwJmMvGjU
RMsA9yMTH/X30HTcfstGLK7OZp0BZoBDJT6CcTLqtc0F5FPsxEbFNEAeHujE7Y1U
AMWSentvqh7qQ00huzEuFlsuFjkM0PrPZ5Nigl1AL4icz37f6raS7fkdGxCB2WhI
2Bkwk63fWqoiWHMcfP5eIFjFz08AzItf7ujBihkWV2Ylj7iVX97CuTiXrshvFPqM
GXIn0d8AmgoBfNtXMPv3K1ku3Zs/ASzZHUjcytRkqS7qOEVWfcW2/dNP79quzSde
ajGJFZynI6BY09m27w0vrp/9fR2MQDOVjA9Ox7s+IMt23E8KEB/+ULfhidzx/GH5
pceJBMEAfrXD4//YhUeKGg==
`protect end_protected