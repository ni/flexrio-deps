`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20704 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
dnVBOIGMhMFpJZXzCENQ2C4zQeA7ThBtRChFyTpiOgLnYObK5IG9mwBzUaQiIULy
Mx/7aH91cWrdMiDoeBFn01HHvt+r+LnNoCN+kxNXeKsYJqiaRCGBPvfrduItL9+O
O2Zjd5uJgZe+SjfCaaMZc9sxK3Lu9yYJp1A5PosAhw7pGWsrCSVOeev+/BwlAUqu
Jw7BOJO8NacrFHH7q0APy4LyW8PjaWp4cY5fzc6Rm4YGdoPn07y2I5ZPckIfcScg
3RuKJSuBtuztGJOUqp+uqKCHXaSgXLUh/ahljZ3b5g6TyvvCJARmFCHCFSSWLSqA
PIyKNLLyPQkE+hLENnJtOSjTO0AATdkm2rNEpzGYAloSSDpupsv+hTWmycZFPtTR
qaisWVgMGAomAIuNay4sbF7jxhH6SWgx2/86jd+hrR0C+WYvoFnAqktuMbS8Nged
VbogkgrKQjN47M07COJYxaBiF3NBtNolE7iOvP+jQt5gL5QWF18dbS1HlE5tYFGh
/n6dLBnLB2IP7yofC9VazgTJJuvUA3sJG91f9TU6PlxGBHqkVsAM4UrvIwrOkvVX
BjG1BJOGTynClTFUHav485AilKhg9u1WD6FjJB2BoulZbmBJsPXl3rin9YpgqSVg
sclfDOEMZMgQOiE/8haNatqY07FluAst8zmYr/zadILhQ/ANdVNIkWez6AMQMYE1
wXsyS4ZkgHjA0b9VBq2bLaSCZiJhfOhKC5k0i/PwQ++ujYqttTvEZCgxm5P2Zrdz
taf54GbmnJ3IXdRPBDuCDo3GawUrICPFxc1z0yDvV7ZjIsI2nJvfNB2mwDWSo+zw
csG8g//ZBL7VbNd4hnVUoT4ueyanfV5m/fgZxQuIJjGULj6+C4YSwG0T4NTKv+ME
H50Jai/DUQcU3/bH10IzEjOV1OCf24JaaA6bOyOIREnehsUrJmv3WNqCr+vkBKOb
9VyzcLcvNUJ+G/AQI5tLftLE6wpPv94zjf5ITQQAqKuk6Cc1XmFETXsKmMBak2w3
xDtYgIAIt6MwNI9ZzxaWBAQlZPGd8G63MMbAIOpvFiY7E17Pj7YfXdw9qwb7sL+i
96lpEU9CyQHwzRaWR3YSCfsmiNZ0ybOy+yk0Og8e0UkziadFN38ecLinJIjqcY/c
hOEcZyvequawn2L4W8QGVPk7S89IXBS2HSW8/vx1jUHHL9M6eESnZzyP+1fxz57a
XAfRFKPb6qxJWm14Zd/h6jAMd7WlJppsNgfByiJp0AxsVkie2fT14M7Sl4tYDDr/
ruRCIqRqPbXvqHlPUpeMNmt3HY/NdQuy11TX/r8vvLog25XVNggPzr7QCvnun2pv
NJj8+BivdUR6S+CK9ElQARNGzkjmlTtGutL71jXusNogjeEdJInn5XYJfff1bdiT
JqaDm8MZFRqOZQOjJ6shoC1BRImF3SjATigiwGDVHA+Tx3+rDBSdPhMlAldy/wqS
a/81zSFtxeHEXa/ZPekyf6477bSrXT5jEKeL1+CfHGoCQHjyiTdL9WrsuAGPcIqJ
O0lOePARhVeHJW9esoZqeM8qVyidTqPo3XfRNul45ErIiqXy8ESXYquam5wZRHk3
b2llYZMwLT7l07BPG9y7YNS6xljphkE2ybSM3DmMJb8uUGGIgTsJI3C+AhkUJNMH
r2HdPdyOJOtFmQtuyey3tlZBqdN8aCGig23mikITLgoJfRKw38A5wumewvQvXMc+
WgtXtXYQGwjDTbK2dc5E+wG9rIsHBx6E+xCaJC/B9m7hEnm2tegmRTrBOu7L/4Gn
uc0VHwpdkC6FL8HchQ8aS+wH66XTGcN0zziFauSQU8phczoeGYONDVZwXSp5rCad
y4E2r+6S7jT2U+jS6Js4g31goKhK8xJw84Swmtk9CR82dz8/T9tNQ/hOsU15Mm5l
qnlUNwDMyF3VBMnNdcbSnImL+ZlU9ygHd39X9p/UVOe/JUr2CXhXBPsA425T92+A
FDQ1dfDCDOKCel5+ZMG00WfXGrT1Kgz6BNQebZqEUUOXDwfRnGf+iAOJX8Czn4N+
04WsvgO7D7qba6jL2asEj078ETq3866rT54wCedWC1A13OGuUjrVxg0s70vPbbO4
RhajzSGAi6uLFeiesNET3IFELxTMRBBSrePOxfM9fzZ0E4RUf66yc5r8jXQQj1wq
OWYJwzJmjGo1RuqBpduq0IXImmXxrcfndBBw/H1Hh34gj3CwOMAxQg4Fmo+gXmvN
EV+HqbJwKcfclxomwMMnJmFEXY+IkJwmqbKnI/9LckmEerSX45VY+dWihLUOVIo6
UWcOqXCNUJFYRsbN5YAs+WGBO8TqFBnwurddtAdgtvKJTvtPpZlGXZqIdWxKdwti
SZomTuJ7c+/lzAV1/Ny58wDjGwmu0jUmIHYiYncle6Vh0DHNJ34BfpX8IO4uhfIS
dIUrX3LsrSb6n8m4x7a7mw3UXdfSw8JXQq6UxFSus/vUKwcB7AlEC0FBPJ5oum+b
dX2uZwYj9hUse1AmFurIzv3PvYnRnEcM1hn2fWiHRr61DJ/NbM3EGrocFhfZMIOf
mfZC5o5y1lAV0PU8XCfuMJeRXj6AFvLSZs6zk3dPa+YqCNK4N5zbtTNrRGUPDFUP
gclX20+LNooULTiMB0WkgL8cEa9+z5c6uTdHo2tAv3pLT1Csuu76J4SnDLMg+6CJ
4O8VJ99y/Ra8Itm0b5hFtfcga4E7uFBJbj5eiOJ1ceZFdvW4Z2CCfjZClBaU5Til
4/dJRaE0dfv7HrajISSemnIAROKCrCjSNu4Ettr8KQ2yyQs5ujjMQgoJe5Qw+wXZ
SiZtDKYtaOtxzHWKtNutd0zINzFEQ8H5P+P0t5K57Q/agGqQpVmwsz4zz5UCYRay
mX8UGyZQ7wsJ9XRZ/6iko6WisAq0BugmM6Hlrld+A8lS4a4ECP0cJ8+2s9UHWslK
VGS65Kvn0mmZzEV5arou6PHxTmEejfKrMKu200/0TnKyYGIy+wXzIRWhIthJfbTw
55Tkdu+nWjEjHpp/10c+xIfozVoAOynd/6blTVelOzO5CDBnEwxPiTZ28a030mGo
jSZXMyDADnn7Ve4Z/Bl5tPECpJqP2DvUxlwDsuDQ+1QqsF3QGsYvtP9xXyL+CXka
felhLm/UsIucfoxyQo+qPseP7lbi4oNK1lPCVSAJshiBhfI9RyHpSxbHC2r+ga1N
u3mYDpvH5fhJ00bYigDpT8P7A9cbMWmxCAS++j+9VbJr6e4o9Fe8QFueMx9czvnn
PTRa+eMS4aFC+SzEeoxWTH6UyYTXWrIV4ZY3gjPIx6nwW39VzRkdnWjrxGfksOFA
BT7GFSJ7okzi5qPXR2+ILoWSFEM9i0c2nnX4O1j6TILF5lBjYtN7SKwk3Xv7kSoC
RVt9EiqNYigNHjcLZG+xaSGumYwIYCgUfRpjGlqxM6GhNzfu8ssSV3LFJVD099k8
Jodg0Av0jv1kdjNITGhbJFhjpiGh8kqjm0Sqbqvgpm+QFpzzqDFf6Z5fPGCTgXIF
oe3jg8UVtsLubNMOvyes5DD6GA0+bPPF8bB1cfvz/VjZhmPdJv5bBQLVLRP5WG8f
vEqMMwEI6J2/OWfZinq9iAxmm22OHFFAb5fZBf+3QLoxu3TUgmu5kDHAh0SnmuUf
RuVpjURa0EpXG5IeRSxshANfjwrB+znmMS0j9bn9ayFqbcf3otdvUWUZpFIiK3Go
2WhjbWsNCEgC0EO/e6B0cILcbBl2QL35nNUrshB7ytqNlBsnbiEcM6LSDEWdnFHf
1Trr69btNJW1Cod4P7R9wXTTurVM7R90qe3YfcJlyEE1xf7G0cb8Mg8lWN8E0GrM
+fBxu3LY/ZQxBjcayW8opEy8HCdQ1bAnRBsMn1lq/cWq3n7yep/+UIeNn4ANfxK+
LoeTirs53+MzAdye6HLlEhRFV3o+RODyRcUQisBCba6uFd3xa10C6WzqSr0gvyCK
BtPPbADyXYeOjvtceresfsXpk1L1PABPMoCIc6Ku9ms7udbrlLdMKZt2tly1M+mS
pH6u2w2lfb6SIZgRjhpzE8V7VIvgSDuMw2tDg5kl1ldxTdU+0x2ZpYEo0KnhZxgO
qZs77uJzzSKRHU06iT/5rFp2fkNh5xVop/biZeYO7fdyUViuPriwz3X0v37nXUBh
bc+9cda5SiFDSQfRCLiX0wQpD6/8SLrWtkRS8q29ych7Q4BWIVZ7pEFsx5AmAQom
YjHJJ58quUBXQhtb9MoiRd7NFPx3d11zuJnIU8WBNm8FP+VaOT6rRESpLPvlRmMO
frgwc2cJmeTX9UfQP3yYkj/podiwx+CI159b18GbAyhubvTGnk/H03sSt3Ht7ycY
SlLaz6eoBhjfaB1WVcBpcAI01dhdqfBzoaruYkr57s9aMjVCNUAcDooBcPNvMM/C
WWaapJjYziZlisvZGI/Fx5kspYMKAz5RldpP7F59dAQ8+OiqZvQTKuJRQB6QDIcw
InkxwU7HLRhq61jVmQOQVlQf+buiy1A97y9xvt21aU6vp9YZxkjTE9BnQ8uT9LvS
taNKYXsHGmsqLWqkRtS3FjTflBhZ4RSB4fuFmjuK7gdKxED+0fVAgq0pNSmhW6/i
8oyWSGJeQ+a/0/8ciUa5Ekl/5PLbNZSLsO7L0Kg2fiSjyQXECuGumo0HjOOhlCZ+
yfXqNcfH9DiRdKOP1ug5kwi+zf8IzCNK30p3oyXtWPt7BSmogXlKniZYzmPOYJww
Mbl7t18nEhKe9GgODR5BEJ8puYjZ552gb3GaVwollEKIaHG5sDkRmoVjkDHZWokS
5eZck9Bw6v0tpWljXxps6FL+0CqRV1eXx38/X6ZKkFYnUQ4VZ872CHLYkHQEqNDA
7oGyBRtyTV7LO0kyq9dP/zF15nX6UCsbNYitwq7fEQ6ETP+zhVBZdYSh1jp6Cp8b
z+qFeiU5x+qKJXYlwSJVWOo21u00Sf56keWGvibq4QCQfl25r0wyhjgPVbFsqVza
oQmMarCmVNoRUvoxKOa9Tf3m1PeUq6ibXcBf7/2kw2osDzR6rHzbv9WJPu8fALa4
SxNK4HuSdYsikLZnUPsvnvwml+PBI6xkaKlqv0abDvN9+YIGq8wvoJ/r1/Z4L+ML
+u7+1MG/mrloW20WnUZkwiFXC7lOsLaaJUW+s8UVtMKOJkAKsbpWjvy9l85gJ+Sy
qJJHv7bEOsDdrl2orM8KFoLBDgQHyZsYFpLF3yPrx2tz7WDpg1jKR+w0Lg5A8bnQ
7FhwcpqHvZR7xeeiwXrZlccx4cnTrggHb55IMu4f9QHuwEGN8hCMrKpgErx6F1j+
0YWTU6P6gKtUhVtz5nuvbpoDRU8tkKlcFgX4/1sXOp4WjJzYtuX3tkN33cQINl+K
3Mp4+gj8MNp/Fivg/iRzygm5c3UMNJtrf7JB8SMubg21OAfzkOUwdcxYnUkue39l
jtOF6U7W0viwBmZbJA8mgyxUji5O1XxZdkAfTfcuHX5dbvZdUjB4Qq2Z+ZxdGPL9
zikedPSXiJM5PuQ+PR3FCpu1XN8SbaTjSggIu1CWEicot+ZfJo+I8d2M14zP32O7
BctmkOfObh8FKxDZOKaNqGvOqyjfghBY4LGGaQBQE2MflVNz8Q7x3ZSiPyaRR/05
PAyLGV4lQl0s/YvqGRMjH1CpB/h5Z5jDkCkOtkkMYp5ViPCEqXEDldZ/yW0LWQLd
e2YPtOx2Bdz5DYmnVL3DOS291IOgdksnFaJFgO8f6fh1KtU8WzEj+SeGsndWVq47
dp2RZ1FIzxRjWGAWMuoejT/dxXO0bpvCRp4RKAsiu6zLeFY4W5KLu4Glvz4hYcP3
Oxnj+XI8hVhS7li99UlABKgCCCQgDnyEuIagl43QlSfxOBQzWhOT8KQEG7Cnweif
UZdNs/Blk8da5CI+7memoTANm/6bcSqoogmUBlpcXxYm2zkIq5byDf/1vGHiwOCo
XQ6LXbJ4lXpgMG61UtQpsTYOmuUAfFivDhrAwmc5ij/wE7HnKp6jReQjMOy0DuzE
1QoPkIu/X3Tjr8xQWhfgDQkXMhIm6q7W+yP8PaCwaf3dhO09dknM+LC6qBZvD2ac
eYEXTto5WDmGkkwG8Zil/sdoW2tbs0F9CbRMlQUMbhIQBEL9J18VNyoOcVYuTsXA
346O/Vyx+lXh9wuFJVimdQnrHnArfk3uhPPpQ7RsLBfKjT1gW/4rVK7Lfnf0js4X
y2dM/woD569w/WPt9Oa2r+jDhmV2hDH51Yj2oiuUfdsX0HVv8tE1wPKdAcuSPLJ4
UwfVPnczucL2wd3S41IQWgzEjHmdqegP47/PBK0CP5Ph16WOnMtXh+H19ZizD1sh
C9l/DptJqLBGIjc2YB43mc1mZOqixkYkm9mx2gZ1yfGvxX+7Igtpg7thRUeEVJZH
K+GF7UYaw4Qghlvr3m8GyQpUtwR2a5DTZRsNrLf6H0HFLI6vIPec8s2+gI1rxdY7
tY56sW84RA1CBGc/exyMQjs5kc29LS9wzUCPRlKuVkiVHlxm6zFlmXjlIXbwMjdh
R2vFowVdgM6EIwfQReW9TRuiVjNql2QSliQRK3Vl09L/8Z5e4K6UkCA4SoNBJNGN
0zHRP2Scu7cF3kD0W8P28M97pXSp09tCrtyy47kSUBX0fcHVbrSeG67JiXI5+r6f
ACIhOEmqUmeO4UinQZYY11J7c0xAvM5jf6n5L4difZcQFiS6r2UUJ8godFgb0h5z
fkb6d9Gr3/jHQGNI28rNb9wT6+iyHQ0fGeMtwoE/ReqtS/evVMGE4vdvK0GjmOVi
o28KUzugmblVh1eb45H7Tiz8amiq87X/TsuBjDZArFuUPTTe6Nxr0YQoqyneoaaY
0ZFFM2uQg1JjuGhPUI095gBHo8NeSWbeHNkoYRG5WD0Y/mbX+O67dSh/Bv3aImt9
AArIJJlrUbhZvU8pIOOOisDfSSEK7pHxODA6uUfatB619xmWL8zcqoraPxtOQgnQ
Wpga07aF2YIqXtDUzfhxiAdathBE1ic+wlaDHRXGZFJbmbSNbANPJVPZq7O9NCB/
/WHiUWbdFCgMu54qxq3poObLJo5wHMTFpcIVGOzCutdWKl6MHGsSo8fZkO7wPHTO
ttIbYvvIGH6J5quWuasX29L3D/6uodGotNq9j0By/Od99t3mhC0mhD/niWkOAPL+
ddD0u7yuDOV9g27oUJRSQjm8age6iQfy9NqWubY0+J7ttH8riReWgyTvSIWSaElh
cO2djUkg0Jz8z8B+T8eSXd2ylSseEhx6Xo0DyHv39J8+gL4Xds29Ho8hoXKtheHY
o7KoOLz9Z6Wj/+aJylYw3J3X12ew09J/N9XyGW0C8P2nuF1vqxtWCz39cop34tqU
b7QcwDhwsFYg8bxjUMQyl21iBltgXyk4Z6fYLYe1PfTvzRvesONTakAWgmMgg2oS
Qx7NTIRG56xPWbbO7xj9OMGH/ct3WlkM/5KvIgiXKnxxT6P8L6O6eWmVRbnNHyyz
eqNmalIGFIEm3YdWGjKVfQuPQjnvUWvfkeV0QZ4/Ln4u3WoBTARkBaC7XVEkrR/b
9Lk+/mJMg/Day7odbG5Q7bdJAMjy6eOFahUydvec4p6IgCePV6o9eDiKFRqpe/g9
dO6JWOZONHftE4gNL3mFK2GV8YDamUv9Q4+EmdXhZlS7p1zM+vJQlcPnU7ROFDA1
56ADsdZEhRvlbcSNnaZX56VAeKPenp/A4OQd2QQZAFjiq/UKXEr3bdTHqXd+rh7F
gAubRR9emn4vuuMchycYdF8JwYwxmuwLpznT8X3++hRMnkpfxHngwX9LMDwNt43Z
OjIj8frD//ugegsPzcH8zbqxMDxnrDHVzEkp+FKaPfnn/5bcNbX3UwEnrWztmJYH
JLOGqbAxXWISVZpCpYQKfoJyM6/klwqiVJ0AG5zBiVjITqmTjY0xT/bAdQpjLdZT
aQJjdDiWeQzb94AkOQunMkZb3Qi+7iUmL8sqhj865EqU6bqW3sB398BR5vEoQHtL
yNn9tz0tWIW2Fy2fSnShyafjcq1N6v8migCOEt2kY/ExtgB2QcuyOKrkOa8XE7uj
mMHEz5O2W2ym6cHEdvnU9oezj4gmfA6uxTk6plGGYflRWA+2ae+3/xI2pWBDj4jL
y4FLHb+8VVvKSpGwWH+B8DdKxnEBSJOZewpjpfBlAKmo4Jt9KqSbO+IRHz5QquP4
5ocUO4R0NwgAYPjO7lzVa1zSw/MjkHVkBDxe5uIzKsLWy3Ik0YJ2/15YLVHh/XmW
tpSxW5he5vi4vwUAz6pT2KwF64CKj/9FGpbAaDyNx/l83OL+84dBicp5QkMixGNZ
Npu5aKMZ4L00CwPTe26btpPQFYtvkLwokmOm6G/K6Exp9/Db7sB3b0bcMTNEb/J/
/ajUjkQcOxpwI0vNtXTTY92Ls83Q2jc/GztZ+Xg/Pzs1WRvVaf8+AHUmfKAQMHG/
38zyBvcZ0onHImnHKsekjss6hWEwT+GPSm4Rq/B7HPteGVHf5NE+GLcVhvM2vALZ
YizIrdjgM1MswFZtFv/pmBjKTP5nS2spyYIGWj0swITEmgQ8wTQqFK5f5hTRXaLU
qghZ2CdYw0DpVA6uGT5baFJdalur/F7j7NTLppoLSt2b268K35MVahkS5lLHDy/D
XU1n2eLPo09m8Vqn50Bf8rY0mwDx3jE65LjEFaji69C/vYpY4tFZrDgnOc5jhUWp
jvCksMO7dlKGUYZzEbnfIifbvAbYfarkkvQpUOsjzjsJsUsrZhOXDv61wlSAbCwa
Q6giKny0TQNPjYjgCjLP/hbf1FnjdsIaiv4bI2ovl5nE5He9lhzeyW49phnWoKB8
kCu6ci5DWBM7PzMXJG3jmt10Iic+18q6CyXQhLtKRw4+nIHcs+kZcs1eoe1Xa3DW
u9frBvkExyFGrXvfKFxs4kOhSz+ZeueQb338S+MdAFm2JZy2rtw+iE8vqy9lYtmc
YKwQ1Dcqi0ZoygMWJF2bUezLSX3ow+U5wFEXSTO+81AQEuwEmWpKkB+enkuksTki
F/joDrYg4meBDspUXFil0r+AGqEEE0GOZaQD1QHhxFmSWCuq8JrEZab0TLcGgr4O
ZuhKhz72FsVLfDY5a/xSHjCB0vmGEM6ypETdhX51ePLs6Ao9x87wiLlhnavMCnol
QY64DvxkHIMfoZyHOqgXzKhQlvfAZq9n6/yGVv6HjIb4ds2GEGh4N07y22GR5TVJ
Et6Ly2Xi1o4Tv5Opbj6r7N66ON0aLNs3YqplpXj2JM100uaAfKbq6+UmAMy0HSGg
n98gFIThJYsf+Mz2K5MJE5gRxSWr4BcydV6vrfsc2mcc4P1TjeYJnPXNVbipoaYF
kCujY4EgDkUJU35X5s4o6TNUuVbH5DpHHMNePLZXU3uAM9UN6ObKqRr6o0ViZnvo
b95L8CM9R2L7SzBUn3W0rev59dZEdLUKe4jRkazE6mitHZ2u7ytLrOEIgfuRHcFb
yBa8xM5W3QpRh+9lRujVXQmBDRIU2RWAbfm3zQzOY96wAHz2pEVnN+Fw+g0/lsbh
CX6EDn4ksERZ48Y94LABLLsBCMmJH2UQDuoOqQaYjUQog0JotguoC1XgP34b6b4E
S16Iw8qF1ZKsGFwmoRTM1aNnq5BPx/QpnNgCXAFpftu098vApGvJ06Z0Qc7arBJp
OL9AHTN8uUKimk6EAyJEDZUF0vsVAdbX7/pzSyl0L1ejkGb4Zx5buV7WDFFlVj8U
bR69SEc+LfdnkzQLLwsbJdI7oPH2f47082bdunYr9wC2C5QXqT2vvIN+sB6kzjuQ
T9XoDHMRYEYl7oCn93qu78R+be1/OfQQ7byixfZkDkfRZaXZ2MoD5GqoWCyr2g4T
TkJFaxAr4TaJUGspy0b0SmNwryYbrR/hUVNHF64sbtO2i3GfiwZehk6LbtJmPZVv
+gL4WqGbzu5X7yKiOH4+HZNAhvMMxuwJi4kSj/Y4CDW3VeACooKRyLX4l1g902rt
5kn1+zZW20KZlmqmG97DFdEYJPXPEcrIaJxRNXxoBehUJe4CyRVFT3ngoEIUQeCG
k0mVB6aakU2R+IZz0uem3AjehvnHt0xKzSNEkNSucLsFiMyqD1sRg8bnqZvegbaR
PZjbZ5ASIHWadZ7ravpav1qv0Ga1S2amiTCBln84JefrpjTGRgyt7TeGEdEfmIda
L6gPw8mNXOyQWPm9N3nAw4MhBcxfI9omB/xHUwYO6/SvjrQLSC3wLWQhZtogdkJU
rOf8iep4NwUiilBjvRSaBiyO37kinCzWpkYlKx6UxlILIZ11v6kuwxf8vm6Qszto
5ALewPa33RTP2PM/j5mkEuiUn1neUAXOUp3jSrOlnuga4f5jA1vNsB8psJshP5rI
ZrjhQYJ5UEMa3nmfIDFMi/VWSsocR/0CmdVNLfYvu3QTVGkYZbgfX3u2Gg7tCCnW
fUtBMBTFNDRQ2JeLTKkFPhOm49pwzMhzp8/yS5wsn9N1Kxt84OWqcor/zitsEMs7
lfS0oykpo9G5Ftvu21Nk/XtxSlRWU4lZiBCRa2jJcMiYU5uoT0k2OswX5HXW2oJf
Tn12mf4tchzg8ALu1Fa994CeqdYAMVirJvseP1eQZgegzX/yYzAJljK2feaJlt/3
XrcwyK26hqzFQ2bcJuXW/CpqL3FhzfDgMo4A5YLkUP4pIZebudh1XZzzx+1d7jVI
TNslb28fDKK1xewqHCuSeagEnxP2JTCU66Lu6/vBBXpuISw//KMH+HJ1493mKy5V
3RZ3Q2oSri04kCcjKVCAcSuCITI2nMbnv/Adk2aBdWbqEw4S7IshoEgvUbIZ14aJ
TYQb8yww+qqmv52170E4OKyULkMd1IXj2wlwbRDN4XPg8B+34Ihzh6ZqysbzImw6
8pUZqrMZVqwKCZbw7NzkccaGlCcNt+3nKjR6zDX6gkXewcPbk1oMAp2Sek6zys2P
wWQRfJVj3sit0tkZYMArEHrmX11RAJ7OjuFMExwWko56KqnZ8kOd+QxVyGXRqHEJ
7FG+GG/x1JUQ4+4u3BhFmG+aI/j3FoFa0xwA2HIYbxSwlur7qeVbABUKiiORp2BX
5Y/477H/nE/bVQoLoBCVr3eQwRPybvNYk3aOEXPe9bHGQ2wl1jwjom93qzxGWj+r
9EOYLm0WKRvQT8IuJ2tU0jP7ylfOukdEWtGZMLtt7T6Bxe7kfwOgcFsbBxuxdOc3
uV0UUuAzAfKSsj+0JitCh/LYNII7+S40VAzSzpStHFA71Dsu/MAljTJwIqlgtgRN
yLfFzexqWw8UoFBNZLZXG+zzWyzpWt3kWgyFjqSx5YG0qdERyX8xlkpZrF1Ex3N4
k9XHydQmwFO1/81QUZaXK8HYK5d+t3UxKosE4/YX/1YK+JL+cPlA29VCXb2QXcaE
oIAinig8MafMmYQ/pLhPHBsKSPjxwX8OGj+jbR9Rk/cerr+N1dmdy9SKnLnchwe8
eMrpNSlf/LhosYHVzGItaTZh1R8H2+Qe+EnqiSu1TCSMJ9zw0Uf8nOMY2xk8pMbE
tdCEOK4V8gTPxuhKkOMoWcPQyV77XUhbm+L4kMH3lYPUKqLn9VeCdjDujegG5VOY
XpWP3d08dPJFBwWXCbJrDeqhjjZiZWsPlMsYhrU7Drk1HKHVkRvv9W2XraCrd1Np
DHTEURvi2KajJ7s9FP3dNK6W2Lj6+vXFmZtFf+c6mXsfUJgQIx73bQIyysVQwkO8
WugSHxqkYskQEcbQjD3AqwCZNx1+IgooHNcsbQF7SBwfNkEU1ZZoLLWjykNASEMa
KhemovKCjvn2Y3j3grnThNzN02p3FLMzoRNqganesmZMYC70BPQRTYjAs4rT5FQT
J1N7dKxXAqdjbzdwhLUr37Q3DUy8Cey67ktBPfzc/lxSYgtvleT98fKODxOl1Xiu
mCTWT5JvbNKoBwtdwd042NG5v1oCBR9IIXh3IOsGXOQ5PHb2SYttFtRDWbw1LZdF
5zWaL1M5ScItNAYP5/bc22H7dPIxX4yhWlK9tmzPwigdXHIsannu9vAJB9tO7xON
6QdauLIMGDEEJ1Sn2REMJA2tfhID6kTH3Jo/NpOlV3xx/6oE75hGdrH7JuvkY8b2
tED/VzQlwQMfcJYBBIOtD7ZoERYaOUO+1FApKLZ0W3wvTn/6yI8tVtlw9S+ExSW0
/HTyiU3voKyXmXUh06EK7acdbXiBLWAfmNdB1TsaLT0Mz6MWOyGapumeirLi0+ZK
uK3eJ4zDRKVjFVL7ycsflDMbNpka0VG9iFwpbgIqc+XhgU73wNnoJm4++W1IYHjP
L65l+v61cyNgZBDNJyCXQzuthk1ATyou0gsyMzMgua+GoNbhkxtd54lUf2wTQED3
siQOIFAlYJWUmTYbVKJzEwo8IEn1QBEDfWyG0sPtRQeh/8eUJjWyZAoB//4fa3Gl
/8/h4v02ToYboIQcurFuIvL0Z9dFLhAMgzgcZ98Im/D6HRGHGZI8G/DNonlpiEZE
R/2GZRsyyw3XtvLucYsJiHn/HPt/y0SPyBpBAorYC3VADm30ca669wh55I6uFfm/
eWjuWdnx0q8LpxWoLgR7e6oz1WkIIaVhm+Sasa2m16gkSkcETXjHtPnjYlKiROEL
ZJAdYgy1Ztbw1gAHBqzYZnb7LRjvU0y2WUIhLahe9MrybqCHoGT5cRx+0F6FEfws
Mg4TRA9V9LRMUj4Us911wWDXs7942Li3VVUqDP85Y1VnsfNFZeIXVTKEL9uPqy28
TDZYboGjhAtJOy29fOGqZt7y9+ZCxO2KMUURY0p1G/F089Hrhs6R/4owOc/nRKPZ
eej6lPg0WAiLmmAwIm+UEMEaR3xF1Wu5BMB0g5/h0qd/9iJ6QZ4Y0dp46Dq6E6Vd
pW/5kz+dtujCMNxw4d0fwmbAyz0A+t2zlEvVPwwamYWHoVhvxVMhC7IZr9hc1x3f
p6tNapRX4llmmJem2mNPzYc6o76d3aiyc8LvyqHRrRfaS/5+hTuYkgytaBp9qiRm
MERqH8lZbqHC0tinCrdeZjQOM+0+CsJ4JJ4qSfmOGpg7IyZRUT/+Cbw5mU8LnHSp
9FQzHjdSlAKvyKk2/zqQC4OEq4kLhvFaBYYE5zsXNLU6hWU1zagRhxd4E2asSrfb
MkOo6t9ZgsIkl8/y2qBNNNmel8847ma1aj68Lmt5JUGgJQGlev2VuBUWjz87b/QN
DTFKnfovfoifruKNqM+K3cT0l5Jd8WunIFKcR1vPtdRBSTHf44DTrZUD+orYJRFy
I4dBc8re/JVJSKYNGKNU4C695LwJNpQ+CpRNKQWRRJrSg63BJrahL2ebh0ZrOHpx
tc2FtDVhBHhT2CrOJAGPtiUGF8daiciAJfYPbsVKhzRd+t0kK4W3qYGsT901Xvvf
SCldkyBywAuzTc84JXipW11kX+rNEXiDTSwZtauJf0NkqXz6V5anyy1e3gNOhl9v
wt/DLJy3o1gAseWj+9qCta0TBuE9vxhVQFsdj7pmBoNDzPp306CAOiqQQLAE+xxp
Cqmbc5DsuFSrrHXKg+6uAle4j+Y3c3DA3987hjcX0/uytkHYzAy7nmOrgnbXIoXd
9VCT2iJqjhYvnll1Tjr+8y9iiTv3GWK4t1U5Amg0iVbFHPscGHbbDlQbCF358pJ9
ze65MxkdPJJea73A1/1+/ZpZ4fbRq64TTxzbYZmb3zGLKWdV9COn3XCtsvVTE113
R0nW/bamce7bAARLjGwMq3Ljcztr+c7MeO6A+k5uzPiKwlcXg8hux0KQ9qaaOxKf
icX6NQ16QRB7U4se0SZml68yPSbSrLW4OnVJua2UfPxz5qYhYGJsB6E8L7iNJUne
952ClqjmSSb1jbishElfw6uLzWGjvozuwy8TzuxdcyJ9tKKyh4whngv7qkYgwwwd
7XnVSKfqfSWMRWERm310BvfyQNngjaml+Eyi+YQBepgm5Pkot4VWfsyz5tFqrT2l
DwlvIXyrjaUDAC4CQU7iE+lbSeB4hPcXlNQUKD582Vjah04G+NuQEG1My/DZ/x1a
+NoyeZ3pNgPwEP4yJMLAdvKkLn1T4etPmJpn4UwiEpXA9v374BFT4QNDcZ4a0rLD
hdhTcfwQz1j4NJ0l98AuixlQUY0tZ7N4m0yPRcfQrKeWJ3ePy/dxl3nFTMGC7Ytl
nEH3XWQZELH+W/VAdcyo1enGyaJ47E/relcFlC/CFgG+fNyK1Mii5kJUHN/SIiIF
5Ygp7eSaYJwQskZLIzAwuKpHj1IderW7tC3D7r53hS3N8CEg3Zz29X+yPNTP3Jpm
ZpoCSB4gtpDCqPHJaSN5g/9sP67rwI3dzHy1Xnk3ASDGbfSCQib3oYoQnil2hZ91
owPAdO8rLjxXadWaSzZ7O+HzB7op5Fo5EB/mxzvkKPSd7zpwugpL+C/ZxifQ9pLw
F3APpcdi6wKC1IycmHXiBEFrwSR2MrxEb7+GMcYHq7DGzco94y9VNrH6eb7Z1/C6
7wGOmAi6DpKzfc6X7VtV5y7tqL85f8znfl5xzdEvAu/BQmbQ5qHvIOB39di5KwzQ
4NvEBjACFMtrylRX9nn96r4gw2V1FFCe2rspTfG8fyQ6f+/0/eC+CBBONsA0uiGB
R5vzLxpOSGVbp/hIWxATcXScX0PNMTxyZ+D3Kx14WOqUnSDdDrbsAUXF21/XGMQQ
AbCeOjKh/+Xj9QeLUv1C65r/VyoerZgVAJIsBm9yjxTDMqUavyPwVcZc85Z4qMRf
PTAm6grn9ZEMqLaDpAn/bZGV6vtAOX7Fv/39Lz1BW6RBxTXj4b7TyWXKflHG6aOo
EVd3X7wuSep3RsjaVJHkn+GebPuZfG33VlDQD0nMqLRCslCoGYUrUOJpo+uschwz
cqjgfE0M25lfwLZBBoZbp2N6XXu7EAmWmdFGBMoQjGI9X81Iyi63zsfh0JVaWj6W
OKLInnu2P4Qb0bJbl85BbOQ56n9zhMiy6htES1yN57YMUmvzHgn9D5bAGNrkNmjf
VDiik3m2/VcBYhkxC9xEgPn0QeQ4+h9+AkWiqDVr/UBgjK4W6A68318sXNFefffW
SAEhsBpdoAn41bF25809/DwuNTEo/MWbROcIBxv52Djwg96ZbJrXo9VM9lg9qd4n
KRveC4msSInULgGdLBwsFI8nG0/bvecTJBpsEeWeVGs4N1ZXdXpjE2/Bxe8xeLa/
4GQJBOp88UA/oLc9LwYvYRaz7CeFdc2DOorsIPzsohMLpVHlYPXxvOGjap3ovEUL
KVnminxWxvwqSYO/ovensqccv8VIb2xo5mjqINKBcfTXHaLoJCVW12aPeoqpZB5I
OVrvU1uVI3NmJzdEPNsYJsk5X2cYKIHQslCVYUFzpt7E2xFq9lnNuk99fWpgsfBf
BuVG4AUNZD0ekPYAWJus/m39xg0LrQTuSqY8pF76nL0YH1qr3piUuaIVv2e9tleS
1+K/kn1ll6URZDGKnWpzrUFBYbg6OXil6JF2HdnePskzodLbPCx1XjGqwyRMsnGe
MzoT3omh9URzGo33twZ7ApbRHn1xhCPHEgXmYl4ddX0nYYCu9LXfYGPVjMtUa5EA
644WADG/WqP59HBkPdQX0dy8EUJrH24uHWTFiU8c0FvYp5Q16kkjoXTGZXP1pvyq
OsuQp8sjy7ydmY1MaN3mjIjnBOuMWvuj7SPLlDoDdXEB3GCO6+2zTTS8nJCGVvu4
gZCayRYOFTCqwh5/n0m5rmDeKlze5YucFPcQZp6jky2dQGxNziJ+4Z+6mbQNN2mG
lW8InUSKD4wWT4zdY4+7biA56e7v8bIrrSiWzryZ8eucZPYzzCnNXxOX3JxOYjOS
7+N/GhShVG8d58MjtJH2iISyY40qxGSLjQ9CZ/y5HVTRdJVIy7ZrqOB50vBXkS+R
D2/s1AHnSDwNGeahIAGtDryvizsNKD8t6IVDmkBk+WpphYTpjDq/pjyiU5ns9Wz8
bNxrSkFxgb3GSTYRFZW1zAU+jvQpKcYOkuhwxrP2VaMeaulJ34IlSNCMbCjYbbQh
BEN9YypmqhBaR4/flxJs3e0wdVzWoV4mYpRCamZ51OntYYUqJgcCQt2WD/7ti0c9
xsH3jZPWea3RPG+b8Tj2wp+8nqNiqSp5W8//YwgZohcn8Q3cE5rRKYW6dTpWKca4
kzHG4ZVF8dfNSzk0e/qIVfVDiroy+1M2ZigbhJqEJsWa/6SDtcKE/ojYwlr07cR7
rJ2G5xVFJlSPBrUivygKAx3j7iPm2hCFU4fN0a2fpDXWoHZeCRyRpHHKc7dYJWnS
3QYeiOlK3wL6uq1jz3dnf5Q3QF1sEE3s6A37PVDusb5YvIHx3a3JwHqDpH35/mH5
aF8WXBhepV8C5ID/CjYYp4aAhRCC9Jgh+3V34HWSxdY1BOOPVwCNKWhtCzpZXmys
cYj7VRQ/EfBSu8QnrTvzqY4lUlfXJUFEjAW2QHQYax7i9oQrk9HtlZccgAWPg2+S
8WeT8pFZ2GPizMbQQtRHtW/PXCxY57R+SVZeXfBBiecR/oxeBdT4jxz0GLHIibq/
lZBiURxkPfQxiOsjBxINFJUdoDC2uL3WA2JR6L/TNYNgz/WNIzKS/y8Nlki4mjpc
HFo8t71t4kvc/Ze88GrqS8ZXhExQoSM9Wba9MUFTSkbscihTMazhrzO/H1GGHCjI
IyFroemrC5DCcXFQSKH4m6ksKHjPOw2kexUT1zJxidZuIIZKEeCVNIcJKqihapoC
PU6sgak5io6CkfbJJ0AEFRmeC4lNILRJYgPYpewfqtcnNE4NlYVN9nqzqw62o+Mu
jyTNNsFIDj3YjikA3yiUvkChP+7xhU121zP9ht9BG+wlkz3laDPoA8qB6IiTm5c2
XkCDjxBS6breRA7LwYC2TECoBhKmXY3ltyMcbGQxZD8oY6l13Nj/HyKKrg8ofVa2
5avcLFliOs4yhJJRDFQsWYFzs0369BvpGz2YGXLoqQ54r8Hmqm+WMY5n1doJzBO0
ECcZ1nKQFKqGTe91Yx99qIivsuu+CjdSIYdeQ1lPjz3r0WdM6ZMTPNbEVPz70gH5
gkKkKNQQAnv4Dc60+5YG2ULTnN8DbO1g/pobr+0BWncbEOM0n9DHoETx8FoeOw0F
agv4I2su6lvlpykz1IHFgc8bt03oT6C9vblH7TY2pRZ+zvi/MrRLnV1t4gDvvNsN
08NLd7nF915j8OFHyIh1OStgTK+u6xDtn8hP9ThAd8pGQhDIUBZt5/mPL3bdSHfC
87p7YwTk/y71JbNJ6ObGyXiTurBTuGpIn0WlSZ/16OtFA5+/jtqnl3l2SQj+2abk
kfr0ONkURrwG7+3jWH0xnxw2andrnHdROypFkkmF7zf12OJJOYpxUmSsQP0u/wrX
DOOsyx0Pi5P4a1xwuQlfUN5HFcLAQTPlB9AJpeT3ayeIHHd5/dnZl9A4UcfahNL2
e+iQcJ+sS/63oOaf/garynu5smHfPrjbUHAoDP9gPDj9Pq5poQs+U+0JhDs4L5de
M6YmKDVje3mdNfkjbp9hD+OPts6DIFHPuG+r3pA6IG5BgRDBerK2NjCTvdu6TsDG
PfOUis2SgQ5kxRGmB4eURU29jZm8+6Vi4br/iDPGfgLFj6+ZEroRPEMx5/oGTD00
7FlyBcslH/6c3B6iC9hy0yQZJqEOEL75MPimvUB1cZ/Ecn2yv6qNhjOb+LeUDNzx
SA0QsfqEkG5TU5DQqeYVt3QzRAHdeLWdH7zPUiRowDQPkQ/JMj0eHjmXGdobCmMT
7RfQ1BFqUgJ0MPF3gnwLWyGnO8vZdoVo5PSjQmHQjOkYU2i+HyODXByJIW+BGPMk
DEvPBZgiXG5eT9Vhq9wFzAISHUNb+vGnnoOPdbQgJ21qov5yo6d8G5/FRDlPb/1Z
t40KqlnQYKoI6hH+89Z9FHFwGgCFcQOX5bJfRJskGOsfKAY9Qw1AEo+VUjrb5nsL
43ssmL6kQZXe7TFpdYqmet9pJdR19bwaWPc0laxfhQHdY1tmipH9T6IqjGqfS5Tn
wB8OvMAHK35X1WKLeleW4k4l/RZ6Y8QlJdL5PFz2QVDo9+mtiTVe5Z1iD1CigSLU
PCPgFAkp2i5iOARuRbuAqq0W7BSvfp6V0FVpHTkTsfYCYa6dm5PH/xFbpIquHcAC
8zuaDWmY64bvReSio+/3fDLK61gbD8pRhBOMBH4Gs0JIQbQVC3Ziwih865K+AZe1
UZtDse/seKOifL8DiF6BslY9T46do5TZkLqa4aNcyPLxIm4uQNpqopsWskboerKJ
NMywS1Qs5N6M7gwL7iXW4EoykKQ/T93Q6DM9lAbeX0VUtzCziIItxhwCG/CvOQba
1iFbc/6jeWKb1O5xcHuK6zauDHpZiL/qFs8YvzAgN/t00rOo8h3QNFYfMw5LlMd7
lmYTGDx+ceC62z87RVy3T97UtowoSw0j6Je6KNQemcMA1bRZuPmLF1n4opaP2wfL
oq2tDswuu26HyB8kGUG+9lnMVp1+dYODjtKG4ZphAQwV05tCfYTVRJj9S1LSW+tL
9uch+vqexmqhnQ8HbS4nYZMYZvqY595wPJT8ZjTetSIy0HwfnGZoVFl1eWnS14jL
jzoRwxjRKFbfQrAxeZgCct6ieeS2CvQNE9usib9qsJd/aUrnBQyCTZ94/KUEEjji
VVAOESTBZL1MS2ksW2ZkKm9xh365kJGHj2ba3q2+nY0LTGPo5bRzZ6XjsnEW49nk
M8dIH+KcrhAQGshWRDa7cB1HHc0pkndoXdKwpLNlg1YUdKpybL/o6q9vC//vnskB
wlv9e/KwFzTld4T+M3B0RSKAph6PK8wzMfrp5NbN38OfHWdsw8Z+LvOyUkoK0j0q
7fgJ4CzrN36qVMs/xT5iCfs2JotC/Kf5a+px5Y+KlQb4FmXN/Khp77A+412OEiNf
0Mk4UhbkDcRpwBQrhpWCP2FQBCjt2/HDKusoSGlUflJDLOdWEWY/pPFG4DIOKnMX
W88N5iClpnNvTD7du96GHuVsEBIPy9+f5TRU8RcQbPEY1mWRf8eOVUkXqG0aZ6/H
yDi8ba5gI7PmZSG6g0EwMbyumHDnt7092/7PmcEnGAIMhPZWHr6bD6fNCrdZfibR
WuNZQkxEuoW2Ayw8RZO/YCgt2nCfxU6F1wotf9AWgrCurJe38DTkua45ocJvgG1y
l8nzPYuY6YhGjyXuKZUd2ffMB754ZYZ8eKzgPjfaOdRErAH4zWXXy+qmE+TC8OMu
WIlD9O4YfYPliFRNKoqEZ1UIu5Xfg9SQW4NkdJFwB0vHR+NWR5YIdOrBEok1aTHx
zM3q12ah8B0A7T39MCY80pLa3PSwajDc6Fb++uhewFnFRKF5emgy/tNWbGgsGHja
5I53GVyfPc5st8uyOh+XDYoRuUndv1vKn1QMiBJIhUtcZZIOvHDhnR76hyWIvWtR
J21cUnsbL3fsXfMHCUqahP8NYwNTSyO9oOBCT4eUMY8t5uGCvjuWxa9jAAC6/4Q5
hHojI3huDExCgYhWUsxlATsmERW6Bj0TGcP+8XznraM0TrcVuX/Oft3KEP6aH0Fx
5f9ev6OZgX+odA11sX9t5MLzLiOBS2b78uYWFqWshjQ+6EPeqQswO/2y4mNozM/a
9wFKWCqnB3LqyS9eQKRgxPxnCn961a+osSOQVroH1C5KiegEAw/cavZLF+BC04ny
8VKBGv0eth/4WD9UhBANQMShoyE/O5z1bP0IsedkN/xFcvJ8uHyC6cq/CqSfqXFC
+30zZxSivBmlu4l24lFFJR1pnmvmLDno/dd3S9ngLsPwKlYAjm2K405C4RinnG+g
IrtZEQoQ+NEddhw1+eRoUUOqlwXSLesLVS0GOT7RyP7JpQIKbk7xaMuShRA50S75
tcMwos6/F86dZ6vCN93P8dJbn9YtOKrobOXF2gB8+WcGNhwWVrnwZsoUXIj0xWhZ
/9gphSdV0OjJfjQew6+i/CJUpCumnF3jxyWZ3Uviu2Rl3fWt8a21EFv66fIQ26yA
gKxx1Kb2ryS3eLRSpWxlM2d5FyWTES9Ps2YCR5zNZZ1/D9/5DBJVEuqRxlgxi9x7
kSFb4jfue1tTSmARw+t4OAU8c6yefnOGwCgdmriUp3iWiw6X4oP2ozQk+4EBfGva
SlJ5VaneaSmohR7AxzdIrAuFnFT2XCsGSa14y6ZjBzXBRn+vZdfs/ZRTfykKuQpz
5b0VnTTetWMYpz+obp5FrmqYrzoXjFcrDvMyarV3M+hwz8oDcyc2rmKfOi6PYoF0
zja4MZrvDs1sljN1mMefhg2JrCkjEMcmp0lihYTOCuhIdAuIOm6Y2lyPI3JfLddC
VMiapKiA8IMAc/ynvFGvLcYxWqXyk3Myt3xFBcTNaHTNjvAORqVvwYUOTu2TTbEY
pH4reaaluo4IJGTnOzEtQ2WLYOTbl+Gl1S2xab12Hx0wyDtvKAZIxlGxredWJif5
/73Iy425/L3g+N6qQW/EVz4tuKNWU1fjWJb/Ml+FkCWQBbsdOC5dIOf5E2l0W2vZ
mRhhA+piq51ekgvH9TqQwcTgLb2w/iN/nj+KRETOiR28+GZ7zWwm2Y7TebRRvHTI
oIvbhSRAxzdLcj7rDjWH+0tcdTzIG3E091llQufvZpAunFSiAvrnGPSRLRCd5rs8
viJS8KRP1iqFH0BOq76f/srFthzvVxVTLINizYnCCrNn6XR/7vecy0G4XWdOPjll
zp3O6XBkdIKxa780J2y9GvSAOQivTj9PTXqeqCYov3hGtGt0s6RzprklKMOlE/vk
BWroMq1orNsY/TkDi6FTV5siI3pYWxkMJcdDc7EGIYKt4NyKLIFLFk2vzpU1ZCEj
BjiP1KCW9nrqmUKZGT9JklOo6ZE0d388lHea/cHlHeAAjWV1+1wEqLcgxTQi1jn3
gBs7HhduiuR5R5wlXtCfVRfhOKkCwji76+2JvAq9tl+TU5h8I9ItvF+XSioCOqFl
9qXWHrtUST6j/EyC8LxEvGEoSyz6eZpXvRqlSgqx0tEV1h4dtrlvwg6CWp3I+Ux/
gz1gdcbG9iPAv5j1bzVWVm2oIC3VB4jv4KYrYL7rEsnZa74oCJ1fHywJul6Ngz0d
919XviNZaTOysom4gPDfklaYHgVDUZGOke2qvfAHpX0PtK8Si4HJdc3et0VztRw0
a2c2tOzfaYkDOGUbXCwfmLv8QboxrAem0JUQytTQnp3cBghIe3JA/VW/U34SAuSg
T7WHfKko2TifR0JbHiy5dB3/YKRQEQT2UVMHOrdKWpVGL/5Jzs0jfFwfolRCnxuj
3hAeQFPvgGgJLFsBnXrMQjYAxnSUn4/zJYHWDab5BV9MDqk+MgphKJDKfzKGrhY6
6SCgsW7iSMhf4aAbx0SVrkSOY+Cu7ehQPB44/7DV+9HoylS8WURcNVcGY+rN1w+0
aX13G5R637CibiZxeiYrATXXo7u+mIm0HieB7PiHUZyPnf1yYkuqsEqRpQyswbdm
NxU9lWGbS4r7uJu4SPsGKQD5zcsH3C9p4+UbNN+aG62XWEFjEQojFwa7yf1L1VPv
F6heSYtZgckh9jZLa37/s80/FzGD6lpNMKV0T5PQALOhy+YOinuvJzdXanKdSLSN
xftzP/VsB45DAZMddTm0hhF75A2nX0z/hTJIvFHsa4qNWCXI1kFlKOJQEX9qOMkq
CsQdHl1EZh+bB4Da2+W5uJnGcYxcv3tUGEmEbNquiu8eZFlNMne+5ABFc42gr4bY
Na3K3YEElwTPAKzzeWkqousQvBfkRZkCc+DzLKqu/DR2gM8672zgS72JdnDI5nhE
c3QOjJW1RumHotabz7kzeuBq4HYYCGQ+/X5AAOSQG2+VDDFy8BMySUttkJQLf5Xw
qJanvOYUk2V5+FWRyKHBQsFwd2072OuYtpIRVtpF5uxjJp4u1/auRkYNxFc2/4HF
El82FO3YuiD+H0zyLc90gYWKYhGB53f+wneEPk3iWFHaewykP+xo0rsxUvKLxXdQ
ElSA2gco2pPok5wR11AUdcEYMFFqDcLzgacguITqGFkh+1qJcSqQWIqbnQzZvS3i
h0OZpU6wGL6ky1kVJ8hoAWIp/jNnjE0SInnoHGOSyHgIyMzSXN2DParkoIh/scVW
nJ+ZxYbDKNpwzEQav6MTnTE6N9obsHP2OGuUhpKirnamFolQo1FPP3ZgNLIDfnuh
+GOk9gGknByKv5cHIx8t7CLpBbRPQI/OApy0pqR5AbnTPJ+mCHUSULOlfGak8U9E
0Q63EzEveEyUdOhouOxxONXzp71lvqD2lTX3NoSAPGKUJo1VcnHrLOdpRqJgMUq6
+GtU07ZVTvXzjyRARiYNgXWGOMDLTlP4ty+r5gZUICVPzgOKlmsioJZFsmSSms02
Y6VOd7UPo9uruN1yY3t770SHpnR8WFQaSOgbwkifk27dbdvw88lX6413+h8oXaxB
AH6DXWpXuReptq2b9h2aziXBS9ptbAMl/9e524PoTLE0IgKnGQ+nRFZ9dC9c1P6x
54kCaMenng2UAMk0DylwfvjlwWNLWh3RKQlq90akbwLRptnDP7JyOAQHTr1L4KEN
AykTbtyILbqsnlgIJ/rYU/NIw7uiG0zCMD6Cb9qoi4Qt0+i8HpKyTMOzxFV9i7SV
RPdR0FI+2NxbQqqMsyYhViCl4zs5Z6PZDC6xoXXptpbu+0ZMJkTDZ3Xv9bduuOc9
d0wOKajKQ3iOsB6lmbJEcxsI01ckiNfYRS7lBhpTAxz2VwfCuVdWH5dBBH1/xeVO
RF9SfrQb5bGABbS5bt7geiv20aDqs5UWpHtu2eZ46sz8Qyg/jIo4LPtWotyCRZY9
5ZoXhIiTwXKSApbVlP6maGFCiopuC76VDfkw8cwZTfjcWW4YH2ADh7u+H/O4oWHm
R4WGXddeVJsCle5AfXu1JNGWW/zM3w7TFhdaDBLbib9Pk5dyIVA2V9t4F8N1gkxz
IOUuYHn3KMTGVvSaMk8i1+jBlzMntqlI77v91AoTPdq0F+QJOVPSERrzB3kgIMY6
vJY0z7lO1OdkqGfv6rnIrAO+IBVpaJTZRerBeX6mWYMC6tjLI5RfLd9VhQoSpJ0T
LPQhc6IB8NTG/50gDo/tm/uc+Y4vwJybuXiFQU7CR4yfVRSljSi1LeBzp5u8qcIh
cqeXNexMUavAWFvG3MP5Rc8iOsmXd2YPcQ2rEGsJDX3857mc/mydS7hQZnEatCkP
Pz9Yp1sQ1wRIOGA8mJHmn/Iu6h9oQzYk/+szR4ae+6pyOfphhZPu+C1jI7N963dS
KhVDE/UEGiutjRWAhZ7Qu+Yg0TW7zMSdXKDZDLZ2oBMT0zJFB2v2Y1yjZmQmn60o
YgP+dCyQdJfJwBQA1cA2CaEemHtBleJWSA6XMompmXfhLrnDfJ3EMeMNnOy2jskK
6ocKvnYxwR2ILzb0NXaiDSca6ZA8L61sddW2NRT7I2BrUokZ+45aggG9uIe1Xeue
Dy9Ln/yf/Nge0nm17l8VoI8gpa3nObDwZVAj4KvMiJkOija+r0V+YfI20YhtejLm
5BUHQLHcf0OJwgtQCQU0YUppwmaEuR1hs7MxjDxKT7S0FfsHm8edYNauK/1Ge1E4
Up/gnSSELBfF3eXdDTscQavOe5FC79vi4H7DQXCMwGjBsFZcIGnkpHk3KsZuBU7p
3KtUXwc+rXsbgCdlYFfFkdyq0ptlzGvwFpYCFKNnRnN55fekQr8qAMU/qHTKnr5A
g4UoOokqZ68Bv0Sa/2rwXsf4uICOhuRXJ6FfbHNuwZ3DhxaVat6ZDVr7nKO7n8fJ
N1qpqvvBpbn+FI2aQ5xBDKPvofOIuersOYizdSJZapGMvxYLoxnwq9R5ZAHmdgjl
4+2DDuIMcIGqR7equU5dyWiC9Pun9oOVigtNEOjnwmX8vUhC0p/wrZt1WKPvx+eZ
+tn/MVDDcNlVN+xdYUh0PpRGdLvRQH8W+LoKVtmhkb5tqRfUin2aZdMMxCD7T3ae
n5BwW0s20kgadzdDYI6CFEDcEAouTkuWi6MW13BWWX/qw+Tp0Jj6F4vavx3dCGkC
Wr1YtW3c+n5S4I/bWl8MROxwP7M9yFGyzUvoqyoiOyYLInKqUT7zLyZPN2+XXSXQ
34t/uBcfBc3kgECCd4Bs5AvrwZgQZB53nSxx4JCMKQwPRX7mYHm8R4PFVEG4Li8Y
IXDIY1T01WrOBlwCC59KB6XmqwWVs0XWyyLtlJg8tibrzHU/mUWLbXecwv6SiJIa
sTgupuaPKzcO2HGrciKxkgdNtYYngQiFPbdvli4p3K2tjdisobpaF0H/0jdRNiyV
laoqMXLKNXvG5g2qUbOABH45pX9Dy6+2XSOcZ+daotZ/KYOueG89Vd7OG4ctC0JL
y0pEobkpVSImKwV/b9URbFs/DPv+kLKmaiaoAPtjP+OsIv6ByOEx1po2+OO+fI/w
Sjk6xBkulIQEeAS5NHqulqa9M8+Sd9T4vqY8pGCO41IbHJptPlSnrqMyLEhJJFjs
/YrE4DljhcLjFBAW65DaVZkpNwOrI0zGseggAYOQuNUgNP5x6lk9LFulDrojaWhU
ssJvcsECZuTNucLvyIK6w+gEsd5ebMY8Xw8wj4SxdBGIbroh/R/4e2E4YwDvQL94
WF10dtSPPhsAg9eMfUAAjRCh5hyXfRr0/UHpU/WA6682osy0KggoRZjjKO8at+FL
8ssN6tzBdT03YXci96Q8YKglXSKbuK/Q2B9rEECUxUENNN9Dt7/POPXgGJzCwLbp
DxPMKjOTH1TB1HHOfc0PSMQWWe9ijlUKNuVH38ohb9ELdPfZI+rHwY7I9FrASItl
RJ+umYKHmSJYjoIZXJTW428D+s9/kXNNWPEhSAFVmlJusXfpyOZWqGLjXhWpLMGG
bOwnIPpsHmITs4moWuOXIoTAvnS04ARCL2kRz7RE8UwJDNYU/NTQCO715gpeGcWK
fm9N3JNU7tA2v+ssGSq7mujMIBFK0VnkyuH5BFrecP4OCSLgipo3PIf792JjqwPq
sgW+7CvQvObRmj1wxU/9e38SrTKC6slpqLf1hkN3EeVH2YbcCmYiH7o3rnawXBg7
Le0KMBcGgfYy96aejeIWn/OOMJXSYe3ze8guXGA8YbYb2KltjwTOKv4ZBip+Hfr/
TOnojV3VMmNOqjqDciWGKuTE5wDnJ271MinuxoCM2ppbkEYeTJGFGbbdGV48ppbf
aisRX1VqCI5XXsX2rooGPU9ypGtL3cKVZ3WZgrmN+c6iasqiaNI3S1VwX4ptmfZ8
9JRT/PGwbaRy+v1XosyzYTY43UmkTRkEiZHkPkXouVz/n42KfYXekD+oyDnGC6uZ
iXguY9m5nKLLqbjJ4ZYUYjoiFcLZV+5DvP2QUMKiZxxaruzIkFmDw4DxRBF6l4mJ
cPdE3CGB0CWVYyedLRiTxhbcrR7vowa/kV6R3PcavN9mHijRuCqoHG4zTzWDyIwR
R95EQwwCFE5r3V/L7x+fpMhuQHpilV4z+oubKtU14mguIjMZo8b/U0KYMOhR1xFQ
P7YFDxuvmGItXgvvEad2qh2agRCVrqt3nvLCyjSaKhIz3KrqRlEokSR7DGmB54I8
s7f9btT4oHBJy9Io3hlpLteuTLgBIG1vw5DmTSnLRYHK1T7lM/66MhLWfGAnlW0W
wLSoH7cVsiltAAEsAU7OO3/tGC+Lo+MsnC3kc0v78DZAVM+vv9zhi9Iyf59OzZbz
W0y9eDf7GZwGZVDyIpWQJ2fo55Vw0eCWetD7wMkwY2gMleHEmEC80lzudAtX2urV
C8i9GhyLgZpF+d500b2d/eRFFB/IDTXLv+NqPzuSDcQKlbsf1A0Ykb9lsN8U1sVr
HIXBD9MjSbIbV9vhjMVAGOg0xgpldmaBN39RyDwudeTJY2kYWT++1uDtrm4jLTAO
h5M2o+Acv/JwooWkCMhV//Vo3/mmpH8LjTfiq/hc74mlq5Ch25P2HifVSQlMqydg
Xb9lnXj7mbdJbLnVzHWfB+GvXiHamQU3x0uuhlVV1TdgjMIdvZmicn1YKsnDAqrT
MSFAngbPbZnEa1h4XPbCmRZ2ilyLTd87xHWlMJ1NDSfgYPjIv0kKsLzzeHuSZpZf
gi/5v+nk2goqsoAGAmJ/uU3cmBtWUq4vwXsQh8rZPwM8ue88GeMhy8lufYpiSFqY
jYbt/+UM5sl5J4CUXzMXVBTFlUq8b7L6KJ1Yr5kH3KUluHiCCpJMdgWrcM+TXksY
fyKDvUtlPhr27HkEtijbHHySA7Om4NyOgecNBLkt9rHL0VH3iy2FjVxzr3NFS3dp
2c2jgkE6bGh99j8EvkII0VUOpeI4s/Fx/+vhVZa1NAiqdx57DDSoSr6jzYjIG5Kf
egNh69dcu9H/mqfltMLujBnNnmG2pQF9VVodxSYqchgDTwWnvcGaGP2ztGL4xUpa
76OM3UQX2WfBNIXEnYbB9brOXM0WCwjkaJD5selrNacuUkO57XeLs1XaKJr0Z/Hy
JT9y5qplQuw+dPRE69jl2JC8Kr05QHNtklc8BrVRHF7v1Sm/FzMj5FlDT/sA8IT3
pAI9p8cXZSeJukUnMcQHGOQtADlMMWErZLDvMyhoThHCcFKY60Bp47hhlj6sRQnC
PG0H17/LBBCrn8MQC3e6rVRUl/s5tWgkCoGqvu5HQ26EIIon6lYZZ5saBAhfhqgy
2pDttLnmSC5ZMEoQkuUxbzHxO7ikoUmEvpuss432iOY2FUSAK6ul8o1ujxu3xAIY
b2O5vo0X9pNvx+mQwiHMVYSrXSqznJHG+oWxx0OUFqAfwPitsPqeXU9UbqQ3Qs/P
Jt+hwsYjXbhHtseo4RZvBpLGAo+9uG1kLEStxroEem1zg9OX7QKltR9VE6764pG0
ez+Td3m2OjGyULUIHJhCwPShRNYjWkp9znxOTwlVLXXrhF+AfLHhYu79NxWSS5v6
NDU+rJvqfu1MU9xHY2PqYTyGsfEiTQ5ydRjqr2bMse1f9mJSNjN2LnRCHs/dEmt7
DjoDEue/fFpcasqQ5vjNs1kE4UlpQ3+EHHNOhkhvMCjEo4IJrzRdJH6k9A3xH4Qk
58hUmAULmeN+cVvCohvRF/NFMRu07StxD7wYheOj4p+5KZA4G/EEc90PUH3a3jCG
+h5vkUtNSat0EAy01mCkVjElWTJ+CKzm9ylTOlHf4nxxrxb3pYufZlW3CczNdaQ3
KYnc7Iajit7kb41qjZZFX5DpGfC0D356/QRyqJZLyv4JOPeV0NtrrPKK8CMuw/V8
zu7esqj9SHAawzMF872F+srC28YlOWciZKhqai6/JH02zPFtH0menAGmVpYzNM3Z
gCAaLvX86ZvE43YxzSexEdSYRydgkI12WFK0hCTeM+Ht3/YVV4I7v7NMqkTYJCPt
b14hoXk85VlV6t4w6CoWWdtvwOuHp0xo10BGqWtNJYYxCEyqjWZGi/6T8T0CX0Jf
Vp4aGBCvYRTzWmspdEHRXM+XU9NLE+Esw+084MAH5ejjSnVLKA/yoEfAG0yAEKey
Fin/pYeAjZ/e917+2hK8Rg==
`protect end_protected