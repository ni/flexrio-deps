`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 45040 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
0ivLeOT4zMq5S+D+IkEISP6ghVrxgZ2wRM7mZFGMs28OKNzh8wzSofPquIRF7Z3e
6jofza2dGmf4j0CDWIKkcpDb7YdlRCYjLml2mpuZNFOI655tEIn4DNhIO82rylHE
9bhM2VzxWC3Fu/59ojXYezeI2XQJwUjAI8/6YBXef3TPCswzpebU3obMG8/taBUt
DsGKBHcRQXcT80FYk7u3+RiVbswviaSQQE4nhKNVA8dsUN4vOCAcYa7C6qkz+XYv
YFcLtt5AjyYpWUdUCPdGnOb8kcKDt7u6WVhuuXebNLwoR7ozydQWsg3Oxw3U+e8d
pBAXDS9YPTg2QlMx8cLMupGfs7RN+3oBA9jXXSmgYmGkupURw47edN1eKU3RHQw6
iOeFtXygvKNdiLYP+7dpbSJsZn+AwqhgAirrTwviTIJuozruXKpM6wYnCvp9pt05
Vsk5aKR+lvuYv3GJPSPvjq3DD5zICgo6680IT6hcLjIdR4Ws8Y7qsbR0+x9RT8FY
nxkHi/jJFEnYWtqZNQitwpmGkbQL0MFecGefLfFd4vSEDLY1X9MhrlBV0FN83Jjq
7smY0szf4j9vAPwEMHprT5+5hcaRSXQQnmGGlor6sClgLvlSnpOJX5wriJV/5Fva
asTcm5BFBHo8rPCNSoaaCjGIzB7emHzHpaMWt6qnUDFsYHH7/84r6JBWDgvSEE9i
ykn7GiJu5W+x8MAWJJULE7xFNMtOK9+QNTG0CoRFijhK2NwINRoQzhp1rgjOENZn
Dwb72pifAqotNmEDYJWBywokzQ0q/+B8dDDW534DFybCBdMurfR8AieC3rvJxzsH
FcfGv8cc13rcP3nrw2MrZ9awrkZ4ukeT9+eWEp3x/iCiEPKxkcHxw1btR12K8Nf1
rvBlJyY7+/HbWhiXHdcW+oDDuMDJ9zrB9UxdDtR1NXuQJGPtwxTh2tjsg4vxJq/G
VSzYiyIhACIg3cCskmkyUnCaUe35KcZIxSZ+7oLEzR+iKALuwQCTD6E9C9dU7QR3
AMlDuVdku7c/rGbfAQ1oZQgcSOrkwoT00ZZTLOe0lk4WmPD5DlwAjL+1IKco8UYL
jcVivMFJU/2tiumPOwKyV7p1J0c9PtYstxLtxo8plhPs5CVHlGycaBhjSkxvvIfC
0svdWWt3SioR23RQf/HZ/QzI6Bny8AhIH5UOHjpgK0WPl1Qm/iBz7sZPlDtitnDd
yb6eGvgag7+C5aRC3z+35/EErOzd3rFjXSWJkzv4DUiIbdqxyN8KFfNn45J4QAOX
NKVaHE6PRjHlKrK3Ppya8FbFrER9lOMvJko0Tw2W7LhOtC+bij9aqEW6feF6ThRZ
8mg/CrIBlAK8rgAMOuj23v3C5EfLGQ32kc1Kn3RqXpcSSgnMHGYH4bOAUyWWtHbo
eXqnaHT5t+MgCUN9osQPeAwTHaC7mHxNuOA1KiZmnsWxkIC/SdgSxNGM67DwEMVZ
3EEIlQUBgP/TtfJ+qRtiQWZ3fNSavXH9nvteGcP9qYANZB3n36gMMUxEUU13YT+4
D2TW9NSp1b544KSG5fKO00irK30r1AyNveepOFNraZ36JuUVVWDNOaovDZol2nti
HAcQ9kHuVElBMiCGlCOC7FgIn8B/koCNfhO1iw+XUJltzfG2u+nT0jJrGR2WH/5x
LMSUEo5FzeuYAxi+SO0ZoWRDCukmJdrSf75mJjwV6EPuDIg8VTqSJkbpCqtPeaar
/CWlixZyLcKNginrfK6XyXTrIzEKo7vDuSqbFm0/skr47Wn/2T61IUyBeiU9c1TE
9JDRwZ5pwtxEoszqOJYrXo3H7aVAlh1Ri+YyOmPkZ7BH7ZWw9XM64dTkrlcv0tRa
CYwa5OigD2M/COetx678Ks78t92bvUNsXDlEoOjsCZ+A+Ow1Y3JPu+S2MaP8idT5
TpPeOqsCsGBCH8IhPq29J/TOInbTwhJjzwV4Fujg+mIwAzsXiyskXon3ESm49ItT
1e7CQ6OM6Y/4VvyTl+D31GWIvhbcoCBb0XyF5kCIxM51tUUtORnFC+1hNtYijGUS
6ukVAq7kKkfVhmG2t+8p7Cnc3ACuMQdvMQumNE6pV/qx0R5kmo6Rj3Psmdz1Y1M1
TNvj/iKX1DOFbxxhXJh+AhkGkzhV8nxWk4QNK/WtKZJC67v7N6aSLEAhbYiu+Vln
PF7x6vqaPgmdXAJXA3fnYyMhDpXfatZKqpSd1n1WseVC57Itdl7FCNb1fohW6ANp
MvKli34gqXaY8vj/MkR7nDZJE5HyQ1aBXAskub16Kvp7f80YOAZHvUhcT6dm6sBz
qhLScxKppvgmr8bUOBnThhlsoSwR/4wt1CZkmbLI1nvGliqBGK84wNOSOpTF/ebz
PHLoupv9NU1OoQswEEXlmGEzPVgUypsYA1mRSs7Bh617edSNzOiwIfnw/j0sS4rH
+qawlqkgbg4n1BnSRHKBLw98lYVFoATRMoOGpWBTWu2uS4NR8dgfzyUrsWnZEbRK
eAIdErTpTyipo6W4szY6v4bDDx7W/GkVc8OhmSyHurXCoZj3pDbHaESe9T5QZLjz
h65UcQj7LJAFiNJ9atmPYbkQBnzx4vz/nETa0mOH4MSf1GIbzsFFdXbOqoLrhrc7
dgY3X2WegL3tQ0B1njstYK0VtN+3gTr9qJSNiz8AodiwX8xqhWvZ7hq+fWnM6kNq
k1c4JckezDiqF6lhaZhgz5GqIZ2/ovoTQQWBFe5deor9G4PVoz6SbTX4X/t9JzEK
ui5yScJjY0vj0u6kpiAQj0qt8a9dNQ8/sQWHGI+4nO4vPh+75h79524CPxbS6a8b
zXBF2DRbhVOCIyK23Nz2W7XuTpP0LP8rPTYAz2fHETdnVSDI5VBtu9IRBl5itECy
V3x/FvOPq6wxhbyhc3L9sDUrNFaWXfGNz8wmXi9H6x7GuXRrMUk2nOIJ+Q1uU5yF
uWUTbkvTkB5eF4M4wE4rvuRZPbt3q1xHa/F+f62KBFHQ7KQLnFZYRa2SLsx/M9/c
qVXIpduoc6s/nHMfDI0HadWKB4nsT6S8NoIjkzAmXhMVXLu8lCWrO0TqQWRCiKbl
o4dtTprnOYSy4pra2gv2mii9j1FkBY0FpBGuofJzdcUso2B7WnpfjGCiYuXAh+0i
CorKD5fYMLz0zwHg0njQU3f5dldYH4DNdYf0YKMWupZGd3ePaulSw8FRYBssbY87
pcVbUgbE7rv1v33JrCqS/lgPPXSkIweRX/A4Wf369OV66WUu4aoAdjWdL0/0I8+q
gWStQFxXY31WPLBo6zcFitY9ALSNs9ji1VquunYgOUy8tpMBGAzJJqgjVUZhvq6v
Nb0pvP77F9hZGr5j3uDfLgRXI/xXWKJQSGDSrynyFr8+4sG4enibU0yCrvJ+IB81
TQx5IuE+/kD4VC+8gA72l2DEo8rUCoqKr7hxv3CZWWNVA6m+GlERUSTKzQzcjkpE
L5yX80AVXqFNDi+bjd1YszpfoHzXtamYhH81afYBKFdmXPoz1im0czeybHrmoUdD
yE0OfeGHacyERas/WX1WeozDql/PutreXxnRLtIrldWqAwP0jvHJe+NHx5Q2M0n2
BGF4sS6/dDqYNm7F70uZIio/nZn6dL7Hdxa7XuXz5//piW7CDjuf1N7AuPLtkvNt
PpyFCBCU5g/nqW+ZjQndio4zoq2AORSx0Dxcz63rXKVxcENVEG1rk9gZnorjTgif
SqBX35fQ/D/d07THrWhD5OhPB039u16Y1K56LAgUS3qfhtjp2XfhbqkJyMF6ITA0
zAM6Pg46EgLXltuAnQCk1RKsGfiYFVTWl855ZEjCAXsCIdVn60WC+4Kevz2sO76z
Utmp218gWf+YaAOIDDFRP/UQU1kQrxrdLEP0S3hhDc9MSq03vCX+GOZY0n8i6fpj
K7WaGzxyl4d3AdUZb24JOGk5ATshF1RoJPXhiemuGkDjxecHIS3qeA9Pfi7mJWEB
6FflX878+yLbSzRI0pTvIrZZf16gLTEXDbAF+53zSfDnhugI3gcRdAvzaN5UBxFd
+/cnTNJr622bK0r6V9QVL/SYclwEiM4XfIHva1OY2TmxDJo3JtkoflqKCyvKlosC
YdQuKx/nuQUpcakF6G6DFcrZvIeJznt2HNufMkYFVnZYvEHSedGeWSqj7MpOaPRl
n2UvSPVqpXrMrJeR4flLAm6vQHBK1bS2vcrirbucVEAcluoZiJwzCwBGE8uDNybC
MR3WlBYGRoh2ItzLjSpglkTMFuelxdkI1RATYy3sKcO8RHYN3aW0VHKbdecNsrnx
lRiz+MKetoTTBcbar1KxCAdF2K5bxizOngePXBKMeTJxdUBzGegLJwAKJg3AusCu
RnEy/ap3sJfTEawdpzszTxzhHF4qf6ESBqmuaejYylhzf5OvhdLVUFF9paDHLUKJ
syOT6BLtugCPneaI4TpN9KhgfgfQXkVyaYJcON2Kv8kAUf0pO4EZqtQVz4OZVzyF
+332eb+MOftpAcXvNAz3Rs5ae8UCe6Y2r/dovy1wN+HN0nE7X42Zjes6JT9eYtK5
9k1ad/4lxJiCJvtKFGkQiTG0eQVm3Vy33MJ1cBGmRNak1CJsN21tQ2bOYJjZ6FYZ
WBYinUJ4ybZDzKZ/ntg8Hy2D++JGpmJRwOxCTy3ZianJgiYI8Cccphdgpabfz8Fr
ztuWcVICQs4hCZ3mP3g27hrHwoKX/D6njtrGby6T9DC+iGbDhOpgsd2JBj3G3t2T
W1e8nWgXl22SgNaxpsGkK2SvkS/qW9L3bCNnpxjagjxTQ9VxLfjBhjgU0ZhPWQZr
kTYtbUKrKsz89zqtAK714Bk0M+ixuOPsXbqCiFIvN7ihtRkqzm9udGzW6/bt3pQD
wzeqb4mJ2lzd2Sc0sz/o88Qt5umlQ28n1G+ya91Z3vtVR/E3vrirDZ6grhEQiJ01
EP/5VKJ2kSxrDfQ09VM+X+l9l8EB85KgTGDtsmK7kbqgYmGylMV7u79JVS8U5jim
AKZ+dCO/ICVdo9LdLYm9BoqNs46Y6Rqk2CBlg0p5vsl60faF6Yk7B9N9Ns2St17Z
3tO4QlRg1vKOQH8xZQKS2juFoJE0p8oqehOzjyvZC6xq9f2+ZEI6MRar/n5jHsbe
ZV9aql4lacguhuefJeOHPNuHkPjKqmzq5nZCQ1A4xgaJKv3g+oWPF1ZhmThKorLY
KIRKGKybTPn2PXlJK2ZxSgEwEbzrIM/9wVbI/ARSuyTMXkhvYA+90DWA4YnWlS75
CbAMo+T62D429AeGAuumgjSntyE8WYk2FJHsWk2SdSgZztpReO9wrMCjsDov3Dd9
Co9YBug1S3wgvuO8VPHjq5IOwlkzpV2jtPWiSNoWz6pF+9Ni555/modWkAR94EXY
q/jA1x/mWuc04iH+48Vppls37s7dS/XrRc6PSkKw/PQFyx4nZOevE7GXXQ+Vob/M
0TTYSu5Sa67OwrL579sUrqTBe8WzlOX/+ADNr5eXHRxky6QGPZssFnnjqYU94Uo9
+5IxcIsHpH+rDmdNMdSr+OAPZf1StI1i4T5cn7cI57XmzGFjWcdQb1auFLPbY18a
qOkATxtclvE2BVGXkdGOkj9esaJt35MuqSKpR8ILEi2JGj4h5fJzCCgXK+VhRVgn
fZESUx7a4tYtQrTYYjp0qyICOYwDfqTDmOtOkHFwx2q4xn39WhIuMsI8pH8pkrx3
UiCoMacIRk0PIzZhRBnBlMb6ZRoBlEXdbnU95rkvzvVtAw+5VZnRahZwQf8TMTpz
88zAkL8c3YZt9/TFcSHjB5gSVS9STkxK8AJS/3Rs7OOsbuGUaijBHk1jaFA9jlju
QY3FtVOfjjS+SWLE3sYb+A+xuHXCBb3VM6qNibFan5XWuTk0k9v3p2KS8kAYztuq
RtfSye2DtktSH/3DIIdHr70vCpbVtmfzYeS9cDTZPCU90qPb7CacPG/DO/50WB5Z
/9Wp8VY9PXxR4GIlUQXhaWDfnzHZzGkuXpVwjZfcXsHZjL9KgwdasTsIcwvR8hy3
JGNutlVS1TJ6vBcZKmch7CSdc0fsN/+HDY2DxTTAnpUoT5jQu+BeOUqfCWW/WbZI
Yc6ze0JtfFcpsS2yA8b3eutwzoGqZnizk0fA/gKGH/FpIHkOv2lRiVACsCLKvuLk
5cuIbMHmngINKMKzeaLjZdOlWzdiXgMeaPZjnlzfgT5mgUs+7vLlH5ojXEwXU2bA
Umd+YLYQVwptW5A5O1Kz0DpyBC6IalE97bZRjpI7jXu1T7vHwoj1L8vXtsavckf+
pirmFhX+3agAFmZs6a8RSAggbdL1IXdR0W56viJe2Uyzp+DV+BXEccdQyEDVWEsr
eHf2/lpXNWadQde7Sik3YHrgaGiqmTOt26OBAROshyxIwWajUfDEbDQFiIdi576o
WMzyjlY6G7kWaeDFBEHFknTz1E0SFwyNThaEhKjA9We1mtopvsjPP2FzhtLapSRs
03DlxeXc/ZWV9iPLnCLJNxVGO7wDj+qDpmOLAyjmBwUDILhPUrQYzedXcNKoq0U2
oqlbWW/9oKnYbd2YWzamHISGG5LPrn0ybSp8qxmucB7lVfzSlv1grpbCTswEDiW5
ijVQ4hL4Fz8aeiKTKnGvPheWUWMd5kFqrSlr9oFVUTTsLu4F/m3ePvRQNDKJVhFA
Y7TSx7MEuYUKPA96NVajN1EmlMU8ZTlOQVGEHjE/8dtuU2S6/mln79MqYz5dBI5Y
ednDgA9V19d8+9uZJAwnfn2ztdhQQXQd+XBqAs0YCq8Hxy1TlCYmJdf5h8AsoFuH
srE3+ipKFoX76uVKW3oyWiWo+lpd7fcRBlvh/e+ARCehkCrxfXcUwZRoMsmaHNIw
/Wpk6lr173AQkwSuJ0ks1H+FVeXa12uVjrCTRcBDSOHVmJEJuTXsYm3MC7eM3JRX
ziSII4pV03O8D/eB9gnuINU+K02lB+Z9eiAUYHAHTw3n0q8Ir6h7EG2SVdMD3fUQ
sYlicbwHVchcebu9OJTTG/w3FoVQedHDRfCWRutPsNq9MVfWiDqDWfvH5DwRNJaA
pqJ6wiQEJf/WKKOVxvUJW+t0XK/Z3pelneTv8GXSkTR67JHw7av2E24I9TlLY7f/
1ZHrdBx50VrUDKHXwir/ve4ooUvitNJuzTqtgbXxDmrCubZ/FA9OziNu7AnMZ8e0
KtwsCc4P1wRCajgYuNc4wZlp2H9iJdgrA9UsOgoe/u4dsVyRwRpKT2JVLEu+bPgJ
hIHXVOmLK3fHHp33MjpdvvY2dNVgJSBeedT/FhvgSxMyg6IBpbkL/SkaPC152F7v
wpnR+tCktXmT4lwqTicO6SmFeGCwVAW7I+xy3BGUtNTNOk7YkIlyhiWMsmE59TXK
kq2ks3Rzumh0e1f3CWadi+qyayyHBaoby9hM7EQDvN9w1sXzSHAN9TnjVIm9uQRm
sNU5DK7kTpJpRuQLFuYEo99uHT8nbzIT9SVXVrvsivA+EQg3ivSCL+9fVsDEYLa9
I68i0iwnB/u8zbmibCM6gzyXhNM33MWg+q+I8yL+SgC9WV7TfCZ6MTFw7Wbfr4Oi
0fMbHKNlBIFuQRQAgBPibeOC97CpkjP/uwkWD/CCjSy18qumLYMw6Zc5xEhFSx4q
y+gWn9p/o0qAjR22Dr/mHFcy+eJ/ed5PE0ApTFwKohBqrdK/10ZOVFhtXf4XXssM
qlBY2f4WjsAbuX5PJ5T4A1OgjBsjwHbs/Be27xhfCQSR0DvIg6IofbCYVxTabcUV
Mo79x3crGvupn680mYsU9oPDZOpycNGw81YvHgBfuH+Py2J7cq1PdnOEOlgISOl2
yZGHAn1bECEFeqHIAY2Bql+G6mSwhYIXNwyx1/bMqSkiamxBtXwWGpx1i9FTvsty
YYgR/87IoJmgX94O/AFTRJ1pfvKnIjrDdb+jVVabvSLLsW2YkNSo9oatjwaABFj+
GzbaCV3YNQdetDOeSH+sBqH+USXCX/iDLOWf3N5ozO6QHC4DSceqdwVlv0R7YCh9
kgnyIfkdhwbr8he0OYhG4yFcPvoB5azyB3ddRRLXSgnUTZzfTm5IXAwMLLzxy0q5
Q2yWhRKSkBL+he18v0GPY6u4fIVaSm4Aln27BSv6KhyNDhhXaFByTqhIkXJSgNgr
6m5mL/n7kzv4E5MydclDVv5emmmWNxhS7sWIhlXBCXsN3oTxV/nI4flLUc/kEcaA
OHv3uHTWtw/Az1THq0aYxQp5ln8hGhw5oJuacVSLJzBHTFWpKzlHBp4M91fTYQe4
LMeGvWYJRuLgPRMEtCvtcO7+UkueO4uiDhw2FipJ/htTanUG5O/IWhjC6GtILfaf
qDFQiFswW8Fm2IoL4AcrHnu/8qk8mmsBR7V8U4s//srVLTGCP7ghoq1Pa6YKIVcx
7rPMIMEcRkBtdN55IQAK1lg3zZ0buekTEG48smWD19kH6zSYhZ2R6GFNN9TVkufP
ClYGA3Y5FyKb4ogg6wZJEfgDQFJKuC4MO8hZsHV/PgYWc1syJlJ3ZIEQpwp3Njmt
392Byw6OouurxThhXpOSUPo92UY0ZMgdEbC/uWrulWr8Ey7DFLRiABkwpmZ23zeU
oRf5Xv/26FfuyqS1cNPFRG5Aw4V30Xjv1qkUpK9zPYEDOpPqjJRx4cJA0TZt/uUa
GSWb3oszRE5FLASGnOQ5i0PSSIh0j2Iwx6bg1OZAKQQPAp8gO4erHI6sYnFo370w
vHcbqj+N8oXK9OOHnt2sPjtqqY0BBIYR6kvUrMAqPvL6r3S9E+KmPSrTbS+1Wy3Y
Qhr14ICKo51kaDGy8bEflFW7C6bbkJENxDDZpWctnkIVfmhYHZaMgEgRdIlYnWIV
JJDhWEzE846Xm8W7hd1zn2cPNFFsDebc8I06DWQUlK/gwpDih7smn9mt16Guf3q3
hXJlCLoV49I2KSSMSGsEqP/KVz6AFAjP3Xr1ytttCku6EWCqIKg00sGekLVnjv4G
asqJC4OORK8sYwBvZMK1F5v56awCIF0kqbuWggFYT89NU7flj1Hg2CbSCX4NVIsY
9P/LSQqKLm24yD6qrMVp4lBv5AO/79n94I06nKrelwdd+AtAnUfL6pw6JbD5JNGL
F5Z9MIHvN5UBFoewP53Yy0XFy6InaDRUfETIRB9UZ3M8tGbZMGrf5bzP6s5AiUbE
/dBSsXx83v86j1RcY8/MDuZVD5X52rRVRa/fIhnrQSxivFDnce7xnw6dmI01hAtj
+DOKyIlMQe/H33IhXZes9kc9sOFN+ql+t4BzYNkQKhwpQeOIuqC51Ecoim0szyRW
7efeaqM1oVFUVgj1MUN2T7B8PQcYI0uuzPHA1MMPDjNkkqpcaV2ieXH18msRv0qJ
BCdvUR9d8vISYdzbAu/RcM3ZmKc+M1Lynuy2lcz01Laduhyltr39cGs65t9DxT/O
nGTN9GRYC3gqjYdHngWn5+//B+ZYCNKhL4QtN8FSqD2e4B6+fdP0BtWFVQiaOxMh
PhE0aHorpGgPtufGSvfNQ8vlPtPpxSUlBIKk9zZq6TMfAeIJhyHHQ73Bpb/oyMpB
ftvPcWeuMVfY5IKLFvNJ0j48/CN+EyEQvbGZbjI7LdTP4pie9WVIyPgXXF++Mbd8
Q8piyiY0T4g21gtI+bsmQZleSpUI5m+GDTPKlgkPtFWRq0EUNAwH0Amzjkz5Zcl7
DhNfwb+vL7GAWnSi3ctfojFcstJE40yBmVs3F60YazIKu+sjlvGXUQFX1lS/Cn0g
IMPhjFwEKr/QaK/om4Pm659VkDCc2beId3ANJZMTP8BhlVkR4HF1GnmsfiQlmaXR
0BiUGN07NnywNOaK3qGcrNBlWg+BIhpCjXIYk2RyQSz3J9eJuG9sJsRTG8Hdiway
KoVv5pwCg6Bg1zKJrgJqB7w5akXuHO8UCAczDuU4v1GP+71UvgZWmbNb+TZBjjUT
vvxWZ5tJdvXSJ5Ag9YD8gVofnOJJZENvAlhEX4Xf78+ESdRjDDOQggZ+Ve1CSo5n
dFXGPbrB/IQb1kVHHJ4ezrSoRy5yPK1JY6W5zrVnriF6FjbBXefMutuga/9NPAfU
yFMTAz5ege/RIkGSKmXmNXmLnghrMR9SEPpBji9+2FOO/J5SAFHENGSV89MI2b85
jhjSx1GiTBWTRDz/N0uz3Tnqx61tQ5ScbImw+fA/SfK0dNRhY74tTjKyVs3JcSRL
pi99UVu3ywROKNS0+bHZ7/u6eXgCPUsp9XXdjsz0qQDD/7C/V72EG0Uys1/FxgIe
DktAvqsQbnskppyY+J+W3G1yHELj4hcOxK4bkKarKKEKWqC7ugqhUlW2PDZ9mHOF
jhwryQ6bplY6SC3bqgf3PH2807eVCT6bzrHKQSyyi90+iH79eyWQkJ8blHAzIsoz
oGvbmJZ8pwyNp76k/K1ApSCjPHZTAGDpwN7O70FlEiGD1W7EEkDnmx9ChqID/z1l
6tgHa9DyvsK6WkUUKbGoCICvwhSSxBiV0jzD1V4hIe4eHMTl2+VoFrkPjuE5Aw6J
zO5wNQEHXpArnJa5dnbZx/p2OxUXdTmdvgnk4dCSIqaB20u3KPclDshwmEpJT61D
U3+MJqEElFY9PDoSeYv2MaCn7Nmtga2ht0EjSMg485RutOoo4pWsBQqwD7Uo/T/6
iaYLb/xlIKeVABMGoELxzaz1lW06jX4H1/oliya6o69OEG5M01452LH53uYVntv8
2EAnzcNJQrivDPsl55bhWIC4x35CebI9pprd1Be/HrrJkcNVPk9D2NOqhAz73y9U
FMoxPmPV7QUw80C/ibnxjsn56Iv69L7xn2Hwv4Ckcc1t3SlAwWFgsfdFngWWeVEO
lhGxHVABtVvspCQhTJ0F/YUXQBQiw/I6AzxvOSEiFuQbjGAIv2x5lXjsXkC3csHs
OjFX9LeUgMZHRUExPxqTM2szBfDNjg3G8p0/5QCyF4CVJpSM55tkbg5vlpF8zCTB
RiToOZKt+R1t54CuKKmOjd7SYklQMNFluCxNAEOYnU3jtLVE4bDH35sr3RAj1wSq
BTFAiBWmfPkfhFD4y5SZdUF7sQEpiyyE/7d4CWkoaqvRkAaFBcLz4DhTDyjsILFe
QMgikuEJIl9aN1kQ66lD74D5CK4toe3Ocew0Wpy3TVOfboZOHWKRy9WcYLojEbnS
TeMfy+Y3+VE2FaVtNJnoxXnRZk8cCt6Fm1Qg3VojGqNBfvpyXgBd9I7ChLX1WBx/
Bb460FBpBtm4s9UJzxWaCqAlTpRGS6atzbw0hEh7BFf+cdZW7CxK/OsiZvL/T9im
KhCL63vy8jvOJvw2n2TFAFu28QlXEOQdo3ZcauQkQqZXgkFiTVmT58MTOxr0DOV/
wXiNrb0qsbe0e4SnhsE3+T4LnxCxhwYQO1tk7joVKBwiB/w9T/4DlRF4bqrxNc/n
wAGI2agZWe5vstbwBim3cmqKhKd6vcNPkHvW88ga+gAP5QMQvuSVYL66MXgd9VcR
exC/3U2/hZWgph7PZwvtYmooikuXqfTz/0EIID3M6BDn7hRDlgRhZHdcFYGbBLqE
vH9+c35dX3wWmi1xpCuWLfXci7ZOaN/SX2X3dQ5sQ/UrYWcRxZC1M6Q8Ul/MQoGq
G+bOSvDd18OYlI2Qr4VJB8DFErOs8wE1Yrbhq5NxhyAgkWDmCm4TT/kz6r2YTnnP
/4IyLUgfxZ4R+nRffOrOB4QX6n8WyO7OHKn7lMI5bMBWtKkOFLaxhmvPdFUBikKe
IEM9q1eXV9S7EAWC6Df1neKZLZraPWbQHdR2D1vfnmIfwSQYVWX+xa/1t9wruZeK
UpKlnY8YsEy01lGmCcw//V7HK+2E9sS02w0Sm7p9harVcka5snnqKO90FvHJdtvf
fUcomEwTfNNzJCb+cb3EhyJQm56ET9jXerX79v3Wb5N39mT2Tps9LB5ZJwc1NA3v
VFUwAHU6Miu8APcg8idXkXuSAo0TxLQMwk79C0g42H5hp43Tgzkvzp4j9G6g9fdj
Fh1Hx6WxrmRdQnnE1gTrrtFBAJMB42kbvKT3evClzDd4DeXzyyATyJrnco+gt3Bz
ItZRfmzeCYmfc+bvUsFDpfpASNaSzskWeB/dcknMO4Xf+9UP9Kp8cpK/BVJdyD0g
G+zRnGd5wPCRW0otGsHVhacpQMgVyFPKHhBQnYcP+ohfIJSt+Ilm1QOo5STJnGkl
C76BRAM7YPFo0EUtpPVJC3xMfzXd/nM/q2ykHFzuUO0R27X8vWmoWHp36rfSXsho
kUhQ9Eiqzi9kPnjUvMQlnfTELunHIxqgkyoBf7sODxg+hEJOI9FRbom9ebtWDAkD
RvVpyN7eKNF/DbQVgXV2V7PCLCCDegc+1qBABUNTfNqTKGx2VnEiWps0Yi0U9fOs
kbwMu8qHpbK+tltmPPVTs6MS3M1RW+nYnakf5Ys7Dnue8L1bjlwzuNgsO8U/enAS
J2oAqFg+QO9Dy042bVwsA6MvWihKCOpC7Y+Lyyat/6/9AVTJIoHlK+sD6aeCzceW
Fv0+DGBsnsmQHJFvHq65dgZaFze0AGYvrcm4omqe6y4uLouecWryrApi+8dEbIXG
lO85tL+M8FZZ6AL2OQXLmRntPMt0qG024NlMYYpWpf6fVv5EGvQGN6VS7vxopiHN
sn7NgA0rXaA+KKyYmDRZzLt8VyeO6JwN2dwp0RsHBLxhkeVP4RFw1mpjXqXV+R6I
rw488SWKFu1Vja6TWYJ0xhLPBZ/rzZkaQpZME5oPsW96hBnMQcNomo7EM6i/Upva
abTbLi+xPcvHlNGLpS5aPafSE0T27ksYk80M9TRWJdFrebDGjb/xis3NrY8BAhkc
pD0hiiLva3Bc6LOil44fQm+YZoLd80/EFjRO932NhsnKj6BWfSQiyt9SRYxiEKgV
SzLqt/+kDC4k0tFwXNRgQXAnAO3NyUXetBHo2TQ2aH2PLfNmwyqp9fmuLAJJP3WZ
LQ5WuAy+XZIkMXO3PvI7RnLHDYlRSaPOjgU2MQtPBeSFYCRfdaKCNO3q58oP1rxp
CDPd4BZbZMXHUbtefnNwJS4N5LPvDnThZd2Nem5DXNNljt/2msW6oCvRS6m+bRsw
DcEPQP/myaW+Mdt2WPDBVyK6ZnCgaKTaHs22P5B6LfGt+qZIbfgHRngBOXaX8L8w
EBOrk80nZMfucpLk26rWF94NxTGEzZJ3mIp6VGz4zUMMntRH+81inW1KDttm5SvI
5Do9MFf+XNpoKrIfW+5VGYCHl71X1KpqI5sXeONBw9lmuhMLQ9NXwoH5j5mhZNfe
uITinqAynIEylmE+35KYeNNkDKUuMJiD+S2p7G5ZQXIkICz4EqvTKosO2BhFH1MG
00vOUgoviSHCDlf4KZ9RbHaISei3U13rBWRDuDo8+2vGEOIFCHBRVTx1/FPqGFHd
BmUcth3OiWLQuAGvuSiYH01HILxF0nVz9OwhB2aHYe33HYdr0gMG6vAeM/eaTtPf
ndX4dXp4eCs6BbL5z126IDWI73p43mARVN+YFZFPb2+CD21fbKOMKOypd6hKHW7O
98R1e9ftZsn14ZEEUVQoqUGu3ifixxrESBxpeHts1qUsNAThVwLCLOSqwphPBbcA
JL/0VXZ+N0YQ9/SCnJfnbHaLdu0fZXWD0IjEV6UTHYynLmwa38gdxKD8nyCMwkMb
bsbVStvoV5kwdqgYFwiWzFJfEaMCSAHf5ng9XBYcn2RxH6U0sPprD1ya/+SSvMrK
2quvSONdUOYskivNVuK0axN60N19D5QTabeivylQAOqLztNODA6C0fufR8Q9LyKh
LM0PS8S0HxWrh8ex3op3Sqk0jNmDYrTKLBBOYbja09fWzo95LLgENuNYaHPXAkk3
Tpda2PQb7de061l6zSGN7KJJoJkimuyHMlzD8O4r4TyuiUq3PlePfs7OHrZf6lBW
ep7xHZ5e7qkRF1oufZ7bBOjLu0v4NBeSJLfQTS6PSA6w6a0js8OGT51KH3/rGytI
Yx8qICzVIvx5RsGbgcuEtG9UZDlOz6hsovxWFH7EUTlDkW872fNPSzYTHp5onCmD
YRIMxmvk5ACH1fYFr75pHeI1VdQHAV+2naDlmUIJrhm8y6tMacmqgVHotv82ZiFM
egkRxcNEIhI8iUbvqM9qtE1UY4GcWxZ1TEzl2asKeXLd/onLwMDg/tODIlg5z+Ea
udOaR9Y2uM1EnLhM+RbRjh45ttgs6l/BC5+4aHS9quKRhbTRoYVidw7O59QttJhd
h2dT/a5gXBJrVOBSoOwjbUsZN65eBfWtUuxXQRA5Y/G8/6zi2MDOd5uxBcb7n4ks
ZlJOuNwEj4MU0SiX9DhIY6hEXSth8BOYhjfMuGEF4ehESGBhhJmzCXPw2KbDSkSY
msXiQtoaWz/C4oD+CVVtgJN4dMrC9QsI+hSSAaCWu/9wabXOkTCxhr7v607FuprL
PG5eYNyWCgWQ9GxmRCkSiqjJgm6q3nGIIKecYY8xoRLo09jeGVnQjdpeG6DoaUof
H0Ibf+vVnNUO6sVNOiceklYli7ktxyG/2achlkYFK244NkJ3metBsumwx+seJ5XH
QkUlIu6Eb5kPu9cnbwmCT8ghMMnEdDVpP3RG1ptTfpzcc4zJsEfM4OfQBwridSxu
GIFBXvHlp6IUuq9SDfeM260ly4JBYjNZISlgTLji5g6l/D1U6kuWoHAhuSCPmskI
1W/GWAF8LcqAkGJi0HJ7fAFIAb/6kjVOXrflNzfPk2mie77CwMWlBVaoKA+bgK3t
a9K7x5LhE6EMPBeMoPowU53pm0aokzoD9nTZA1roDw1eejcNcfzKjE8qtnmZwx/T
SXzc5PCSK0crNn73ZkJZwuMyAIMy0ihzeR4bxh3Apbx1AEOAZR78mXtdHMa7b0NZ
4o4AQnPysCx/MegcvMeQnen/Hs0Rip6jHePOIC3q5RjPfPfvwdZuPloM/kq6o81/
NVdYh6LvF3xmdol6AdjHG2A+4NkvHhQcc1iU3Uvx7s4b3S6IQ82KhHUeQ//ywAjf
9/ekoDRaD1RloewV3El7c3WkY1PIANyMyrPBZbWLFTYR7gs5cus9T86SSuWMs7gx
yzdKZVJvTQzotx5gioITI7YsuTua5SOCtI79Xd8DNmcyHzI3l+DSPmUpMDwTX9Rx
z0+3sCN80xvdFAlc7fOh6QwxnbwSpLwzfKZuIjo8PTpMJuJ0SDCiTWhk8nUDboDV
o3qgmRJeUP8WX/s+6qT9m+WA20tzdsxyTzalujYXwdrIAGaJVKlY9VqtN5l/SxI2
4dr5B8zM+GiUeIg4SX93sXPpGwuj0pXdxDkcM5OLYQcR+gv5Ae3fIXvakwnBdoyn
o6nhE4luzxrc4vEV06kOX+/jt5EnQ+kwaYV6Pj1kKvWBJBBtXw6hjZxnBdrmrY/V
5o8wnRB3bbwYkMvPXiASJnB7hKbXY5unTnnJb8S4kbYUNmgLo8eMN/mouCEV/YlA
VOYvWC9ZXXMSaXlTztNEFOxi3tUEu8oo3XQv1BEILcy3X7Rbm78FRM8APLJw6+P6
ohNb+jHlaECOl1RDHr8a6JTh3KeFUuu64ZD8E6Opm/1vqGulYJIUyRQeyzdkb3mt
X9FOE7L04kJhnc7tDgB2JR/paQaER/71m83cXYV8yEdiV6S31opxZmlzTZQMN+bo
Antl4oxpN9XD++Hf1QGXKREBMaSYgOKo4KlfDNCuqSkWobv3tJDkqAKdC9Uw6ao4
V1ONcgemCCbDUJwBg61efKGpE/T+pUVXgcg5KJ1suqWpwX4BVAFeEewDT6laT7jz
uAdx0psQfH8fYjuMLi80wFNZTigDyvKNJ30a8ZrQHHBuV7fYWE9/vk7Kv2GKXdMi
i22W2XCpXyW88lmdKPBxmYnwFdWJ6daWpTtywiIy09P3D5IqMhmW1uE45mlB3z1P
QFIQiQxSZZa5jpxx0ZZRaQYw8+XjDAb9QNuaJz+ce5JuNeY70ZPOqfel6LNomBG4
hU+OmknRyogOrJrn0uBGgRCoBFOA5kICIU5qkQAZFn6KBCGXNNInIDbfC/wfjefQ
gKLtTGQySRoTB5/MuMoJJ8PcQcgkcXzUCq43aTuv+RtlprKkcFRRjR9VD1D7BULk
xsXk3r5PIw8VWFKxvEqcR1CA5Pxj42ehb1RD7P2383PDGjJyhsqq+izZYzNpFjgK
UJIGTeCelJrFQ/2ZM9ZufSoi2W6RIkgL+cGJUH+kS2LfPrd/tDFKq4XhtJr+W1+R
EP8TZIr5MerfoO/5Qb5Ezb/+c9AkLEcUY+kMBwgP3eT2RMM8uPWRnSO1GZ0ki2bM
zIcuXtmmEhAVn7vhQGiJ3pnq/8wA+4bPdkgIehw5i8o+GVVnqJJfniwJm1YkAPyO
5tpKEv4e0UFfQZ2UTbzV5pkppnyx0thI8qFex+I1V23Nl0CeiuYwP/l2vytH5p99
FMvsqlzG2wMtAXFO5FaQfnh2zW7D00iAtzyZiW2+vv5CZ8c+1AvLhoDvAg3r8HW3
QjJnwBw21t+FH8ExI6S73Iy4kLJ4ukvFjg3yeEAlGOW6Prh9O8YndqmYlQRHSbki
rBEQk0wU6ldg29UOq/mY1H7NquDNjH1Hx1gye+kvbZ6e6x9V9TnCMfZV7CQKku4m
WakSOTYXunYFnrOr7ldrsEXC5TRfU33SAD8Uy9FEgHag34yRQQ3VGiUgB92u9EyQ
tALyT5rhnnHY4Kmd9Pr2k8LjP5/BwGUUrIppoIxTbD8VNeMp+eHstU7MSR7++Ub6
rbpJYPXeJDTf3GGQTkH7cnAE2X8Dsh/dA+VIK5L1x22Z4ssgpTaTbc21/6TNPCZF
0RTgnyBg2aWl602Zw0ardtEd4DsztumDw9cZ6CdDDrbsEFgKnVA1GhwqbxK53yyC
wEIHLW5+d+/yvTfEu0U8n1YiTmwdk4JlchsHO1yhaF6Ml5Eq4B9cAFZkVM1vs/qm
9ReMLgC+QUUUIzJyUxq95npNP9BypGmVFJVhd61/pvBJFYrPWnM4+biAGP8cTbVF
NCsCQyw/ewQWJw4E17wtXXnLK1FRuRDyANPRbIBW4WEVnv4VkEAiqB1mU4w7boOY
p5qP0rJdkbaFAKjNtbmVP8d777ipLO//tPv1DUx02afRDEAJSSP508yU9PFh5jn+
KUdvJW3LlfixtqlsmtnM5pqHrHn3rj4Dp40OwwS3FtGXtwHV/a7MP4MpjdWKV4hu
wYwKOJWLREbOkfrYbJ0XNSf1oydNbd8v8Q4gkemRDpz/ZfICYzGH2boL20bgFoB2
a5d7OPRZPtnf+NZwHpD/5gGQDEdfG0gEjhPoQfvevT5zbLsOv42Lajy807tSGnVW
YsE+1Z5VQ9P1sPviL/IHCQosgXiMOmga8FgDJGfBbUEVyRXA1hXE76k2tzfTddHL
9pxftZiVieAwWqPupdqSX3YBAp0o3d5AfIAqzgXjC+875wppMvtngcUxtLDVNiix
1NgGXx95sqLo5TfnSoUWgo/cWnnT7LVMNaUYdBbIYlTRV9+dptSrU3NoX8l3BsET
w89ndae0kouDYZG9HCz+LAzC5aHJoLCtKdETkX15vzi97VPC5VgSaP4cyiB62QOM
bcZAJb7pND7ipYfkXA6a/fWysgxJ/I24YnVZbfEJbdaTT+Wxr3wJKDtOr2SBmiHR
t410t6zAB0p9jYzBbs0IHu6Nu+h5JG851+C91ePAEvUmeY/mHM4bwrpLKJjANaV/
LgOB4A1L2+WRPy1Ygd1wMGw60OvHlPwtnvlahJ1EyRshkJ9vZfWwENeDi05BV7ZA
MdAVC/zUzT1ox2RrR2MNC5b0ZcgqF20imjZifn6ztu0FTKURaXqlpzDcwOjHxfas
//BRY/RktFbbpeke03xn7zvk3LF7hA/OIVgPupdgitR1cCo18X3xgGk2D8jNTFNq
nuc2Fddm9o2dNQ1chbzRO01HtlLnW+63dPLFTDG6JfyPPVvRQ0P69nkEfzuCagxw
R/jgsaKAisCMoRA0v/zOEZdb9HOlK5mbgbcyJKMr2q/A3gwIo2+a+qOp1qXnFFzo
UONa1TZJIoXBBE/Qn7jEfBptwDDag/dUdlz7CpSE4+H5dP19brOEGpj4wFn3DARI
Mhr+7JFDU43i9NhieZB7weCxv7MFiQrj1AbcuHlI4kPQwvsemr0wHA9H7xjJAey2
xTBbu6Z8dcSi902qZtt2MFEW1YiDFYN2c7vVXvXAx1DJlhtMbyDjKBmM3DauvDIE
01wSwN6mnH25AMzVQ/RpSIYiLAEzCiebMhYJ0xHA4LYb9N7awYzF1nkubp/bsja/
n7Sd57K/ECfrV87mFYjncgygxrYDOX3ckJMd5tOHugthXNfzVOneZI+I86ARa29d
EjkWyvShnoH164XFDCkx3CjGsYUubTEcqVSz24GNq1JGmhRmt4w0aUfLZ9N972Un
Lcdtdq1QfEyMY110wo/nLeP7YV6yV5gaJLBZwLL8k2+N/cGcmlVbC0wDUigboObO
oeEYCh5Ko8QENfPKWlNr2J9rTUMP6+A843dOkEvw8HI9Q5MOuIZcqFjCu9AB0+fG
CZnyHbag8PtScbZUhCyZRorzzNX4sFeLyEZy3I1f47sUZLu3wk6e+6kEtylgqyCX
WngiFApQ6bwb2RIqEnfQNNb0nEdnoh6W8Zn6+g/tTyuu1JIUP+Ghh/aBd4NpmiR0
TpRK4VY/AqzvR1hkVlPp9/PdXJetMF0FTHXzjdgSojl5OJE91wsoCj189yO6Ysw6
mM/A3gwVzoIVZG3G0HSDznMS4enT169y+WpVRbiKzWZaWrcF7Zw4u5XpXq20Xv6t
eFnAkYHhGjd5wTatL0fzUIRnNeLQFboH5MB0syQdmXZobTUoZYfyyQ8GP5lYTofE
flsSMhWTbaRai+gwZGoJwa61aBFvF/CHzVexUPrqujxPGKguybQJ5d6OEfBW6fWO
95SAyqTQ8KLOHMGTagt3rvHmnOF6pbbSTYA0CYw+KhCfMTZ79aZ+kDarxmwoJ2c+
IiyjMwHKs3gmHwEf31Da/jtPRJN9K5BFH8Yo8QcZHWCN1+iFvSuZVCzMeX5s/0mj
FUiCBDdGJvf/ftQu3XQo6OcVoeVurxUYKiYospoj6JAHoOg5eYr6UImRtJHb5YA8
lhd/safPzcz1i19GaO9GjDSD/RcGo1K2WfWgzYYX1IxB3pJ4De/qsjkSTK79JZVs
/VFbVgGQQrE/9VKE3r68CjsAnHg84+sLRoNOELQBEjRkUeM/4YkXuD2/5qndIjue
D7qcAYDhCipWdPmW9UN4iLoldjCjcQJpyaLNFOgXXDc3oVgi1mWZ710tmjQSyhhv
GkYJyihFIltIcSPHOpYV9vJJy2A/5++LZY6AU2s+i6yIfJCZbimRPTO/zrm9zYlm
U/JLMvuvXrFa1CMdsCJCLt/Uyuh2nVBwvdBQDkDZMQNuPnfrxBOaNjSUCisHdPgM
AZdBxPpoTWuJxVm9vDvM8movnRPbSX5koceczhnxjab4Lz8XfEft6moIJWnYWRhO
ew1TFUjRVvFmahOKjrsm00H80ZVU9QU1P9Emw59hC5YKfXvIlVqeaoL0wlY8Cos2
hK2JeoJx3EXxM6u+73UrBbQKNqJTVbarLOO5atZ1zEeHfOU7QjiT0BFCrBRvDJ0c
DlreanieZA1HIi2EMrGydzrgfGFlwv6ILeP+uSt+mCBJlULSOmo5kUdt9KqnjDDc
QsFBnIWYWmCyVrxjezBdGgue/Ph9jnf9oXdD0huMY6Sbz63GaBSszun+HjeILK1k
B3jemEE9utgIPreXYvWTjNoERRlNIi8CvLECoOQBOz4mkVecaR7+UWbIWVbc8hVc
ACl9xNRa4xKspj/TmM/+iwMCRemVj9wpANO1WLrmgMKbP9//H54XSXLwnPR6xK4a
gIXoskBcGuKof2YIp9gkL7rmKl9dODnETGQgAMtfVgT6yQrZSVgBkYv/m4OR5cyp
hi+JMtRhQ0D8SyIMCi+hQhdDxI+a7ioMqnyo7MZ85JCqWfECHYPWG+p2DFJGsA8q
YbYljlohr8UNjJODEeCPQYpruZy1mOlVuLpKsWCX0sfTpi83oHZqXHVc2cG+OXqd
MbLxPLok7AOpIWlbkfd7IiGICLKmYzWWqONAYGijbFMRKaJtVspW+rJheZbSi0Qu
k4ob8MF7unulbUdRwTfsKrPZ1oIgioxZohh3/+CYYSmPcIgYd2S4M4Q1kLVSDlYa
Dq4AoLAETSO0TeAqa53rIhCqqWWd1P6G/2CORqnypsgr7II9SvfeY7+L8NVfRmG3
NlIvlKmhazQh1AnUWQY4vxbN3RKSYSN897cnZkqyB5E4Iw0+xmHJMRujNKhSR3v7
lG2DMpAPp706AJDClrK8/5nySW0ZWk2df3U/7yh/JIhanYZxl6+BOg+1SDHHCJXw
61bE5JZ+h0YUkN1ZNdrD5keXkmx8V5gPfAE/iASFp3aluz04aQ8jlRqoS+dy45iG
CUYt4A32uE/2ARHkSAQoR2EhcRRLdRk5sAvfBvRnB3gpJiLD9qu0q3Rm2TfzTggj
seQgXG9RtPR9FTdf6jp5CuxvvflbfxNwnrRJPKRjjL88SfGojeUOeUszITYEFNxp
7XHgQQaTRF/LsaXjhtIcOGmzsAU/2YsZCaHL4gVYLD/7IVT6Rcqoi8z8uddRDGiW
9BwB7uzSBA/EAFfjtEr2O35agMqzYO5/cTr1wtN4RtG1TVtaD2IqGShZfJIwbRVp
sMjRlCnXg7aWrX0ogrPIjDG4d/ooiurejwrGWtMqUTjVW1pMSYzRjpAnabYpNx4M
57krTiVkKu++aHxE4qLfvge8PjOAUJOfVZszb1MZPy5nI5z+J/FD/0T3/zA7qN98
eHB7u1W4o8g2cH+9Lv2ixiYarNFyXZNvcY3hPjrbEt58MS7TuVZsHSFiQbBfjNUr
R4FqgR1eFSK/qarsSdvXtxGLe+O8p13R+ijs6/J142Bdd8VjOhS8pEZyxPuztGH1
dRZ35mCVWFP4LgOYxbt8x6GhDdx+HMHDAH7XJqb0ao0HGaHMx9Kc9Jty86dhv+B6
Nh+BdTtrOQGJL6/7Rk1MU0oY1dwpT5uBm/UuEAjSxy9Ojtlt7lVsHX2LEz04cdW1
BQHQX4B1sKPnsLm6BjIwmAlxsztQ17xA0ldHh1DcEcH9Q7ezkZPxxsF0CK1dXZAE
thDHooKJrpKXEkNsatF/tUSjw6LvpkpHimyTC3KQ4smmk5L4AxBeayUQe07pYCPD
rpwxX8O8Mb6IPHuvVZBrRHKzUQy2HK+oPtqQiJW6ASqWAVURzM/UHGocUlZ4xTVG
wl2zQzUyIBy0NleChMbJbummnpRB+jLWCxvgx8nFv02BoVkeUFVGqWwBHItaigX8
UhO0VYDz34K9Tnj4kUqln31ztPZfPJY65X8K1W46jE7fcfb6YMfeVTvj+kHLdA0k
BJUzdVRiJNKkudN7xatwbGCpZS8FO/rK47l1XFS06HpVu5sFuztx8r49YexNvsg5
LEQofmycW3bRb9sfEt859HGbbN3WDPmb1jIJqx2lhy0Xdpq/6F/3EXRhg7rHLUgI
OxA128HTpzIe+ARIh7ORZl2Wb61pPZgtBV4ULtJul3MV5NYosGweYq5oCRM3j3Ba
kIcxONSESpfRxM0anhe2B1by/fu8AHxg/qxTZEuVIMq/zbKViJvVHboGaOweIWIT
2EJRoKvrHa9Hfsw8u3uao2Gu8au47FDuHHfsRmwObngbaCiufZlVV+1wwkVtvo14
O0rgqnLRPQtODEnyKiDGp9odOFEEnVBWS3eAXdotHwBL2K+yyxf59/uOgTjFHjsr
UwZtLnLiJTpo28fo3JL2d4j7IuQSum2fVHNMgaUCQalGlQQ0KUw536Q/IJ1xiv5z
S4/uH9pnfkcz7Zm5z6gSlbJhEc5BbCVXwa8Js7Iw0rW1ulPUv0AcS8yQUFRjrXin
RHgE7mKGxYTvpP6kbyp9WIz11ZSxeMf8wnC3sp3eYLIKlprqck1V+Q0A73t59oAY
ksqaed9DlRaTmQCZi/CgyGvuLJmFJWNbGcPPxpqgPmoJXEVddqE4tgKaEgZ4GXl7
RA1a1B5uUOh8G3n3hVa3SRiEuCjs53F/M4/U3mCanrGIAwurwol7xx9zANoq+3nI
ELfOSeuo8GKvxySwptjJH29JtYx9QUgmsKQZ4exVP+ulkdsVD2/bLeSfn0fE01wB
C+A9F3HeF/gvlqnArJHRL95ibKsq/tmFsSQLXFOWPq52J51gtwsS9oa44wFd2Fu1
pqs8YI/ZT+R746+tuUTI5kSeTc5hl7Yr1A7GGTZy3AoD+bKO+JNflcOWAIjY84Av
DsBk0ANSMwFr1Zc4sSloQapEsqgPilnZE6TUgfatfzU2qNKQa43MV1LB+h47IU9N
FayWyKJOZKZnT+SwtrEYnUfUJyKKxgKkRi9hb5zlnP9WIjPI5fo/+mWtxTYso5G3
4/aI6KrNa0P7+8lEMDx/HSGvHOQBDCtKCbqeA200DSgLQg6wcr2zx8sqQ5IHKp9D
2RO7t2X+H2oHnPFiGm+2+tWsMF+4i1UDmWA2AaR/CzpP5+bCpr67963iuQfnaeca
5MsvIuS+WYzQi8PfgTJTC+OOuv93gq27yI1HXeH4Mfodqy4qbkJahN23/DKIjwWv
0AoA+One2XV7lkw58zoFDjMtAt4XbvnY862XPaLoloWbXVVJnTQVysld3lZRfKlM
nbu/pqcvBTCNUuM2/IdbS8XxgheyYWaIM/fefg1lkSXz0HSvEY/kyTZp/j17exjE
BLPyiTtxrYliSWVq66AczFa3bZw+srSeTbrnkHJZ90XOfBDTv4/YsbEViDPAKmXh
veh99VL4K0suX/Zm/itL9lLXid0/GNdR67z2RP46llrcrD0Tm04kHra0TBawHYiK
iokBdG6BJqH8xhTdB4lBX/OskIu2QfzRm7UUaCLZr5Ge36qSLzPXoEI0W0A0qMC6
7uztaJ2IRLj7wFbvlSgebieKHCarwIWnI8ztLpuEbr1f9hmfWk6OgIIvl0ljeMjZ
wfMvFIvcEOdCgOAcqFGAla9ZJZyWDY6x3su98KohsCNjF7hAUYf+mhr0GZ9/6Yst
bvfJPwpC0AvqaMqIJFIa2If0jJBcFOaLZ7Sx8zDI9RKxaT33pKViXNIoKpLx1os3
Z0OaPnWmdukAqLUveVoNoo3YQthbDuqmKlc/RaMitek6WDxEIQQruDqP6gsGOS66
fFjdYmqGorPsRIBHGeihZkN9JKX43Ue7FYBYSMbdPnQfGhLEyCzlGxIib4ikXtYS
2F/GzUWAhF2KydUn/tzA1tUn04tNHAFEIkCechORSLDiUtN+iPC95WTsS+5zxX8t
F0h7uavXxG2bG5w+GveKU7h8xA0uGzm2/Lj1ty+2dR2iMbnBrUDNNy5u1fRJ9oSz
7+/Xq202/rfOZnT/3HyXJCumYVKmnOMiyTigOZ0u2nptUgjvep/XdaQkYUc3cLQ2
CpFXmO7LxRgnzAmaiN/4tVnphSpRVIHSuI2+NlrSEnex1OOcnDZQa3E4BQoGhsu3
NaMSJfZxBU9hcOVT4HiTHvEU0rlKCQmVkm1S9UuKZVg+vsWC4DXbb/E/5xYbdGrg
hherF3xEaNcZj+Lx0mZlwiHJqnQq3cb0R4F3bK5TjUA5QvgiFmavAhObE5jLXy8z
R5Nk/HAnib+9u8ztWWGKmdX2O0ChG7uINMyCO2BmD+tIjKQEHhdDmZejCm85KZ3l
5KYU7pfHQ7qngzgBQgWqX/j2imx4YgF+Iqx8YtQMYg30Mji48h01dq8s08QcO+aT
JMPjnUgmrjRw3KMCLE57T3+TCRMUPLda+G+VnCvclt47GhDDrScmMTVbbE+4GkL/
+sc08o7XrZai74OWwkaR8qc2MXKUPLjiGerZZDIGjffj/bD1dJ5O5b0AQ7+Hj0Of
G0sprdyIawMdUwJYbYiYUoxhdV4QW6cwlrz6OclCofZ6TqSNQdhGAEYT2/lYrUsJ
GN4L+0PIfNetj6PUWo9ESDyfkURIUXGZqhMOaihe2yphVNfK8eU0N3h6Q46hMXRa
N/y8O4SoXaqY3rIm8drp8KJYcggHddPNguK7pFHYH4JphE925Jvq4qGAqRwJXCkF
x86lzZ3Jxuiy2etevAEwL0icHcDpZ1ZYY50mEl6Sba6wTNQlliC8RmrS/UwrDD7N
gDyAdtJGSsimMbJUhiRpoqdQsiyxNDMz00LP/zOX85JWA6dWwiEOZR/3sxtch6zV
314Ykp96+z1LPjFH2vKGx8N8WTyrsJY9bFIm4R3XZhlJjTtqerstwJhhuNItoDd7
layZl43/HQpM9WVdguD+uh3WhzRzua3R/fLco3UYGsWfV1Pd8BZdF/EjO2OxnhFu
7XHbHlbtO2gVXTXGvVYfk9JA6lD7N/V0myoSK8q64m/uKfnveWFa2MTjX4KQCTeB
PI/YJh9cNB+MslCnn0jjwxfy0pJ6VqMBxeYjMK05gquPghovX487aQUdX65zPuQz
LzImzCfi/7/DzavGOKlJTxmgGrPUixCzGHKF/Ot+nagCVkSJIYHTvhol/ABPdzle
/2/pebWI1zp5Zo9h7wGHE9I2whMc88/rJfuO4tGH5v4BFFhgskYUlafxyQn4YK/b
yWLKKhN9OGmyu90cCqbCxlf8npY5F+7DQDPpQpR4YoTFqJsKk6oNCeYSPOcYdXO7
pyU5ePKDjWwUrKlYFmLaK/D4fV1iV7VrAfV/hnon0o/n625r7I3vbna3GZIrgTya
rj+KhbRJKhBRflAcB+Y8F1PlCtZKKyklY0oJTWiyLegg5m4nTCNWf0Rs3Qc9kQGe
1LhPr2ZGyALG6NmI044ufZEhLA1qmHfd867qzICBPewRahxXyS3A0+fTbTn4SF7M
/RbcSJ8cz63MKkom6kgoPqZgBx6tirTLQH8CKsdnZvNJ38q5GgbJueVxDQh7TGFA
y7PtLkrYnM1GbWZlaT3M5c386ih/KDdcnsZh29n4ee2PU/hY1pTEYyjRlNCTdXZ/
/SnQRXpIbYW3IE4Cb7Gz54Wm1lw2Q0/MLzINODfsH/Nqiqou1fx0TGIGebUekLbQ
Xw13y+7HrskWhOOFXGmOc7QHffwyOxw0c4ZxtKaEQB/QmYFTbTfBqvpzfg+R1Z1e
kfQOGsp44naYiqmlFEoNKEBnHrr0fqFKTUGnfBGJLwvB7ZqTc0SYkQWx8M2bNjpG
UEj+Wvf7d8yZanbEzkQcA3FqVbZWyk/Spg7Ojb2XlkIMG2JFLMKZF/flWSXJ4Zp4
m9MwoE98knpjMFgcTAczbtofKQyGrTAkAbEh/479tzYMBWpHuQWK9kxN6V/0itfD
AYU8/1RcYHx6qdZn5SYzM43YZDgoL2GrwSAfyVF7sXBbk44TLSHOdBZjXGAfgntw
T3oQvHvcwJdCgdF4IEwW5h1zsCiv/24t4NadKp6+ZUVxRc7B8JVLz7ZEzYec0KHG
PlAKEZ1p6j8eyfHtgpxWeK/UhD52sxHR7+33XmYmJfpP/YB/vAk5cJiMrD3doldR
7NFCorAisBaiDjGsVQvIPZTldbI0QRlloUafCohspRuyk/tmnnL4LhZbmrxwmquX
MHvydFj4apOy25+wauxpxrLyOvSjGBe/Eik3rvEURhOOcXVHeF++2vYzs7ccfy0L
CAEaCfg3TuVbZbf5s9kyYfq8+6BbzPgat67vaImA3Tnd2XIvV1y1jq9cv0S1P+3r
dYbPl0HYmVA/UQnId6cgVhPOpt8ob13/1t1+5RxGYYeXN8Pw0+7IsFtd3DD9Uott
K5Z22f+6ORyfj+cKyA/D1HICp+n4gKSzPWcYnrymZM0bFC1DF8D6WhMw3K6QzLNX
Vk49M9uxz4phZ96hJEQ7FSpwYFaE+UBVweBQHCC5YCio6lkBRw0uvCCATfXyC1Hl
23nE9npzSXVnKZx7NpbHAKN0qMRB/bv51yOyO1FCaVU+2KR9JiCbTezc0aB26jcz
GitCJM914j2ch0Emy6nIbXSg/zebGVmroCEbOlAb0ASBJpbN4wT7Bj8FfUzz/Lad
FeifzlpUeuwwvioYpNZ+wxTA7t8A04XFCgNbB9whEW/JMG4rJr4goDAVNzTVUe+c
AGe0COoB6QvGZTkkPjib8XWQuFNsunfquWKWPPp1PMz6P3lcxM1bxzeZ1Hd2B05E
EhP+t63npxwBm9c2jQR0B+4nlsJ4bpizPT0ovvdjRq6KMorLABsqwjmPYjgUNC1j
E2JsHafGRc1IpgkykFdBJqRFrFrmpzE/gxxamh6OBPrkpPsedXz2/vLbvN8+G5HL
GRd6jzkkfP0dDP4bV3NisG78cyG5C1sKPRKfQ5QlOYgDYf380w5MXv/P10RKeifF
cqxI0F9rNeK83Q4PYZ5fD5XW2Z0KHH1x/jW1EeKNki7WzY2rIkWMktmdygxOgCdm
C64yvV0gwJQ/ezx7rG+HK94AEQE07w8VTDYIMMoft9JC+ee4JHVAOEPqa6HckS41
dVbr1JbfO4aJ0i9IgrsJUex80sfC4t6ckaGArA7ntGDrbxMktk+14LtwmCIpHm4V
kPXUY5Oi5fJ0fs93Aukw4cpLt2iQBVwwgFTmaqZwdGt5l3U64Zkmq/kR0+yjgFRN
KZ9bAl5b1K6nKlYW2dWIapKHleQFYZ+ezjnsf9ZtzoViO/7CphIAEIYQda4W7y5s
NUc/RnzJrDkWJbiuYnGqkGYb+0QKYYDr2qHX6ADEBOugzMkdn9vOJMXjHZqSPb5p
D0oqYGf8PkedOp4oJtNue4FhHOAITgs/hzB6pxnn5Jk12WJWXgxNSaxrkKuPEh8r
4xkwxsHFjROuqhHPRg5m/32+ejxEj6ywM66pIy6nSjyoSq9mgdEmwh/j56b9zgon
ryihGfSE++tbCc1LJfnhJMwBPEmf6lO6/wiT5fQ6ffYdChMIlUk36GQv8QUdNvHk
8QNW3v5yBbaPmj46hcu2FCtAlQY8eaGKVuJRRkdRouhTaAR3meM+ugScDRLecWpK
w5cfOYGe5uQYzatZ6w7owQcix4gPsLHX4xYwmUJfvxt5E4txtjl5G2y2LNOlbLHL
CX7j/qqBrfc87QsZdbYqgW5/BH1wS6rQh3ojrQ8vYov3zrXyOJtrV/aC5TOY7C5i
RzK3QHWCr1zPM8YEQtL+djb48GOD9DUpaNLrRToZWaxCZFun/eNeZyGSdQp4qzm7
ztHqKM0/6JZH3xQf/L+bxV5BgWbUVhDkMtAb87/FPDRdRINHnvmSF2M1diZ57MO8
4rRTJud/5FWfPjqQH2fDLGJysQK8Ft4XncLIB64V5HPkzNMleAlt/YzKJ7GWo9eF
2inm0sp/Nz7JVOKj2hL9Fige2Z/H1g2YSeWYQKkennw/QuEpYVuHM2rPHd2bny8Y
MHw9lq4/kseP9uT6ZSEBbHshdTK5W2bUgZQiDBtPvMz6JYwauEqliNTMuBgCxvzq
wJADHXvYVgnpy5UBykeklW7xUG4Ua+AlqboRwj8Ny/jqt2e5M8767g+PXEnrB57C
QRekpzcIxV1crqGMJuy/1Tu4mZe8wD4pn1VnxBG7Uhc28t6ycidI5t23ZnXcCvyU
zezDXIzPXjdknEgypFiHgCRQtoRwiiXd0Rk7zozFSHSldPyl90KVGYatCV4BTBgR
DSWs28xrbTAnZk5neYgC8zFQrr/Pg8/ip282AfKJav8opm9imocFnfsPO1LZ75eP
JC5/9X3vb/Pfrb7IIyhvV3Jp2JFJbHsxDQrRUrTwizJ7pWfUaNF2UD6olxqXDWOp
7oTrHtCExaQHxqnT55MJ5SMhvQWukic+6tU5/jDQXi56fZTZW43ApdgsiJ5zIxWT
yije+0tLehPNVQMirk5u1Ecdr1CHbvS77d/4j3edAXryeTD073wjL1UEaEVsEZzM
gOt74Uxtovndf0xF/kAakC0IJn8uApbrT/DLumPsxzvn5Sat92G9/Q5QF6GJfwgl
a1Tko9TYl7qcTzxk27N5aZj93fXZZ5qQBfN/HqdGEkThR/VWaCCPLcCInneBiE/V
MdoUsE95ZVNF5izWc7Tav5bqAAl0+G0PbC5c11eUVLCuv/H/NnvQBY6HtFtsrL6z
FxvAkn/WVRAhYCPUxCZvD6mJrYYqjJaSB2Onz5RyBmF8492F2WxUYZLcGq11rT73
pEB6f7OvfjjcfCMP6JoMAGrqL49F7NdMbTlu9j1bcZ8d0KMqZAFG8hNuiZjywSkd
tD5NbSxUw1A5KcecHwtpBEbjCCGtdgq+OUWrILz0algId4B1PXyI72da7E80Tj/w
C0DohM1Anx9TH0EKiVZfxcfRdWh9mPdHwFdiEphszqjTmLiNEXhnzey4M/Qmq1+k
eNLmoxIKpfmfuKCzGh9TOKdxHhdZoxUma1d3tSxSmU4GvYk1XKZapDXgqUZ3Yluh
GiTyM2to6GpRWC7eQnIHjMHgqmuAqZXmhSdQTWPfk6dW7iE72xREUEV93Uu1oiKy
5+FOxJ3IEjeivnDCJb44Ca7/9KmDoE21tMQiIBNlALAy5PEX1bbpkRl1y0r9srFL
A2LdUaDWuvkhzJSWFyteYcOTu05MWNei15vaFy9NWirg5DnqNcZJh5Vg8+jdfxWz
GcWcchG3WGlnX6WKIMxwtqU5PO1fYBaLITprqyLd3PXQh7FrdNmLz2bDEz6ZpRre
zpBVWcw8vm34M2XhNFZPjdGkffs6myOh+J08oLLo9XLuFeRl9alnfb/9YK96OQeQ
zLd7SV8jZGKaecZUsg73Wu82FEhZ5EP7o6yRHEtUHvtOl8ah/8C7b7CwfmyxAVot
aZ1PwZ0FvEQY1KFfNnXuWsu5E84pnp/92/V/QnKtAKJZPuc5IdR26oGra5ji8mZr
Zls5GJ2P4d+Dr86xK5r52RI/5n/v7xQhAY87LXz5TZy7vqhWRBvTvLDVuM5emIWk
BhgZl0H16NCPm5RWWfwOWIKwuvZyTGALqlmOoyBt5TydQgARvs2z2RJKO94StTbv
kdbp+Xd4/bxbKL6eyU/osZGarZxYLBsW+iPOz790H2DBSvrYHK722GTrex/CoBNu
CNNF9hHoImuPKDSQGomy/54+r/mpPNGbH8a9clUo5nlil919RlGQdASE11UMbQwd
Z2Cd+hciJUrFo9BvqKLdKjILEzwo3nnW2KLDu2RLOMoiVjIJUrLE7BBkiDSu2OlL
7YvLRhazhuz8f+TvFxyRPNfZ2Ibtl4xMZqOHuGdunLjC3GMMGWc89oxu/xOFghnd
KvkkTxZKx4taAptH4kn/PMDMwBDMBexu9rugUWYdm9nKtHlUnZvelC/52DBSNo+x
EzuMAFzAaFY2SBU9hzjwLsG7vWUINzO7pdY+SOlpq9k6901sn8TWBbwqgMHtj52M
SdnAaQ1ICJ91AHwVLFUiSVTQSYJfiNyDuAx0y7kY3RxgVjs7rNm4ymLaEmY28Uwm
y7eoMx1/jQYnYw+BmOT2ADq+ybMFVZPbYIuJIdV1yerMs+AXqR1G/0TCnRJ3Ieyz
B1Srw703sVOyyvlLFMNhhLcpR23ZQsrQwSoUzO4CBk4RgEGYitMoIRcKegtFKDBZ
AUI1nIp1mkwwBrrsKibqAzlj2KnAIgV5tf3W5QLrmE+2NRs9pwJgoOaO8szytpvV
7CpzYE8aoO3AgKh7OP1/b9L2QoUmIw2bZk8Q2pqjkMyJuvEwKKSZQXK3m05PSkDJ
jEgfd8tM/jf7lXBjinfgu+09+4xBkBfb37DlyutwMacNoLqJ2WewazDseMS3QvBu
X4FYYfPW5GLg3shTASu6QslDhQwopHYea6DUeMNvsNatHTRTKdKGGc0EqklNk4GE
BIhxc9nkjCKEMR34fJg7hR+a/LACwtCuXGwdNLPYKwm2DwgeOMcGOqAXGSCbaSBA
hEFb8Eu7yitWDv4pj0H8o3jMwICgCcnrlHSBs1UZs4fpMWsq8yUe/BFybtosV26R
PsKPDNrW5QxsDD2lxsyjEjlrQWQT0Uvkj59WcJNs1DqqyzmCsrVeBU6xk3/atdZs
vKZzt084LDPR0hn/nlEt9TdkFlgoOFOz4iHRwYH0tUSKq7V1t1wB3sJTdEuLzjAa
dN29/d+58hhM9Ull6kFcKbZVVdx9xsOcxI5KeokIj8htIFkilTV63TIt560lLdRp
Pitcxc34ELKt454h9+q7XAYqFE6zOP+EzzcbW6hOVks3J9ImDnI9ye3ukJsickrQ
ju/9IdX4TMiOTaiI5RHskLJwMCs4NRVBpTC8mPAmrRgVS3qLgdop0AFAyFc5BRYH
KuqL2us3HwX+g/WIF0b9zdeKaltAyx6XdYkQpLlch7OxhJMp/hvkIp7PEQOADK+y
2mowYHEG8VKH18c0NfIAVC3pUmszDFsXH8KHUEOuUCzL7EWdR9WxjL0rkIXg1CIy
OaHa99UQcuJk/ykf7Q64ULvLmWPcVJ2MqS/i+NOZwyGRlfhwI0LwlETHiFI6zX9+
J3cieFmB5oXfagPIG6Sqw8eiBX2Szk40Pm8KqqN/0+d2m+gpwzmv2+osRn0bCb7P
N97eyliIqOewJUYYfv0jHuGeIB/Sk4MfK7SVmO8Me0gHQGie+GyHgdNU56O1ZeA6
FlcsL1RWSsLf6UIEWQOaSweYbjbO0VjQLGZM2V9z6h1j4BxKesJRYcuFaS9WBh5B
h+akEgPbm/ggwcum0c0vjAfTQ5Y4YkUNTnWmEUo43Odk9Ag/CNFwvyMkAmo6JY7U
wyYJKws+0SyzQKkYOjqbbwFirapDhssOPin9iAioExslaJxmWmLwY3+ZcVSRDRhB
FzFnihyiNqX+JXk8SisOdM25a40dhTyG1QIGbUndld0xyGPA3QJFOmeu9VraKOMl
EKLyYTfydsRBz8jyo6xrzGQGxMAUllsA4bLT7b+ItQRzIwjdj4ePj/dfx7LFo/ek
wDVjdoUChmj03IhEjcvcNFCWACTT5nfahcTLTYP3EOXOrrBI8PwqDLu83tlTbY1i
dxmJt3fJ34OWfPxQDKnzbagX4TkVTNOWcIkqiojImFeMkioULwXKUdgmIptE6PIX
Ji+SdzhzhQ4Ila9q2O6KS9yNvvV/5XefbnvE9xYt8N28/cpdt4xuPjgVuijrJ31N
Sd+yzqzajBoxaVP8SGyocaivb4OVcLX1cIHai4LqSWaU3QASquhIscaYnR7Lu8RH
D946jLFtrRCv3QxR9cq2XemHEgN+rBDhx0goJtK3btEkkztL5jMqbm+HgGR/PFEK
nGSMCaArnlMDbUDmrZw3vmxUwy/SquoM9F52dXQGnOpS6b5XOqRPdv1Hj+/et2B4
J8VLRySFYLzlEWwacjJAeqkbXU+Wg46A0pop1c0EU6RwIRHTMlC9ZHgu/65GuGmz
BHbZ5i6J7jef88RKRGbqwq2WLlCpFkRPNAUDtG9QvBmc0HxMjUmeGiwi0wGsP4Py
2qtaCHrz57NuNJdkldpm9R+8zY8pBZK5tP+x6qy8r+OhH1aJo9mPyRkfXWeB2SA2
29xBMnL6QBY8A1SdXDfpuEvcRxmpl5fBQDCoMUUixlpKUE/J9FtyXZNUyXjbPZg2
OVK9cZktc9+p6d8zU6Xw9A4w/rksvetkAXI/tCn9sTaseMTwg0BLp4MDuVFvuwGZ
YsDzd7wYj9dj6Z2bvGmAeTXogfLy7TJ2a31JygHYne8HtB5OH7UJVQZYCOd3zT54
RrdID68LMBJLODxIoGSsApjV6MTYS0Ys83MHejfi3OLdcpUMwPo9QAGcNXOOFKiT
ihIWaBj7PXeGSZz3pGzqqhj/OD8ueUczLyodlS4rvXzjLibQdwDcrUHLFn62L42G
7qtKRcG0cU+OY9+q1WznpogkFsuoOraEwZlzU78fonLlYd/ZVNcUogGoch8Pu0Si
osOzZdvlK/uC+SufI+Fq1Y+HHJ73MZO2JDrb0xbJB2PjmcMMFLWQLUqhfukywM54
dSVV0ElEe7HILX2mxW67N1oXP6z4Bb+p6diehDz8wzjO74pUwU5ssmluh+lctBni
2DkCkxL3LcxeWTBpkQJWtU/YzXQtgI7TKyMIFNyL6mnKgTASHfpN0EWodjadGeb9
TuYq15CZeRV5jsvftpOLdjn4dJ7kE4QcU0QT9JSI7bfGtF4ObWKNQFN9IH6SEIyC
GTqDO3lHqPNKTFM5SFtNtDXeAsk0w1VWZcNu6Wku/lunHn53nKwAx5Gm2BxccF73
h9xdGJPVN9eW0KQCvILid9f58P6keO4QpLHNtQtfo5oqav2gQoHClczvnO6FBW64
hlhOOiyluASrdZoCLh9pMpM2TT1YG4gKLGpNZit/Y3XhRkSuOu0TSoBMdZk7k1xC
aNRGjT1u2qvZbMg0x+aV61jB9paR1xqTclPrVBsdxQXyszzxhO5x3ph0OyjkVe3d
EflGoHjGiJYELz8q4JhOuL1JEKfkx0A0Z6A44QzfSOBhL/d83rdoDS0nwHi+A60x
FfkgWrLekqkX232AZ3eAJj2I+wiY07HZaA2HmiDHD+Pm1kGHnS8QQWMtIBTxOdJj
h44H/A/v0dgfM8JECkp9GCODpxcqU0hiY0q2El5D4gr1PW6Y1MfQQaHJ9XIroef6
FMm7ZMqiSBMR6Ar+SfBC7yZs6wH5b5EQIPo5Blrp8MjtAkwkMgnr1KC7DyB1U2pS
Sjb1SF3G0LwC0mU76wmvUWh4jpycCZ9RtcvPVuBpcMQQswLy5gcuAh0HPXMd/45f
VZbEjUIqUq9Prz/RGRxAKFiV0WHqPDJFqvnmx1hhL3hHtTFPp3Qr6ZoeThrTqeqC
610AZtLDO0l6SSIZ26oDga52bLdrr/IMWON0Ln9yXsCAvgSADPDK+n9U2WeREaRN
O09ET53CwcNuKFbzy/qhLHHnsMcWDx/Vvf1o5LXvm63qKdyreUyqJiUu/y96QS1O
B6s0sHnPkQl90Svd/fqX+aqXLqZYvxgWWiTbv0A5FCH3lXwO6GOvhEGvor1fiQkJ
A+OlCWxTudgPMHE/mmidlH6oHAIHam4lChaR42gvWy8tKZse+sCJYHJSec+yDnSB
laBtVSRPe9VsZg+v9nBwOsFejNH8EMFMBk7zacCqca6duhBY9SfMBIccEFlUpBJp
hbZa5Ly06wVQLliI9FWj1rX4FkXSVLBJJw7G7RnXnqWzWAm1qpcTLKuwdhRO2HCH
zzWfc+R1pvHzhxQ5tKas9SlGml5RRdwwA/6vw3QJkSQM5+uKt1uV035kX/a4LY87
ab5gQArdy9gfzpS9z4VEPVk+ZaWnG7bg6FiIuaEq6o72VjRhO+ddzMEXLPGN1RVP
1ws/hScZlVJlhqx21tmgupfEHIByLis4Dv9fj7A+mAd0oe9NSisE5e1YkL24qet3
H2v16HUrPqh/Inmrl7g+jaNmBaebbzoQFokFtU3IUxqfBI1rHd/9/swtY1aciJeJ
kYACwadQx95fntftv1RR1ho3Ugl23RLAnNZEjBdp9mpoZfl9xh5HZHKo0cYCPVju
5RfTHnzTR7TMIhm/SS6xibH/3t3Tn9ul1eUbnU/KpFUDULWgrNaidxd7+4kNRi8G
JoVqtc/Yh0smURL6Te73SKVXeOwwqXD8v+5w1xTYprnrDH2OFBIa/JFAJAgBDnVD
iZqNlEA5GLlnmRXWpQAmcMhTiYNRCaTQlSvqS2wjdzd/vDC3vAYuqtaHqO83lssl
Arb7heZSr0fJQCJY2BLE/AVdvZ5hogDPWb8mhyms7Df3OzlUWPIvj13CNXiCGhVj
u7XIh6N8KemJExY7iryKGPzT4zG7P6o37IFs8xmkelQv+HHbKJV/kNToQZ+uGF7H
8QPADCPagK5bz1c9SAsB9aufyAXAy44Hss/+y4gl5JKXvcVK/LqpWS3JtecZxizF
eyJeazMgsjDadUKjFZQrBZrKhOP+IF2Mb6Uy6ZAlQb8ASSskyHTCuj4MDPfrEi6U
6x/4jiyyhpFAV0qJ4mvyFG4IRnVvkeb3R6+/IPcR7syok9o3m7reteFfMajNHpcA
CIP0L29bb5CCGH3HdV5r0Hi3dC7QImAALAvFda7zotUmhO7/b70O4EMm6U1bkip1
MmPWSpKVNjYhU4nYJSLlx56m9ziWGOcEkc2qAIxzhq4rUByY5NN8wov5HBZV+YGo
kFHcjCAuoNg14TBn+V6CWn3o/7MsCRUWY3BnjZeGr7apHzYtVWFwjERXWEv3k/WQ
V8W2EDLTdMR3mzRmh6Qec+hsDcU8KZbsgxJaSuz713xZ2kL7DVOeRLPr1GPZzJaV
4vghg6/ZT4Y8VTGc7VNREe+nzATWkZB+fPfxsoGwg/0u/46EiWcX+WDbEOoIm2DN
mZi/d3sFvKDL7Y/gtKjssOkjfk+c1hQptjRtS1fRsFNwlJS8G2KkABaEb1ZEUcV1
JvwqQeEY8OO4cLPSfV7IpASWQdipf9AD4x2wgC5hfVtyW9QCeoulckOGtByE9IKz
mfN8iaoouGxwByuF7Lau+1DXMwz3MMwiGCHQ772r7tInKusspLUgccTqIoko0nu5
ktDkAs5ahJTPKBpfLl8sj2FFbZpwW48EuNUJbA1lc7MyKEUnM130UeC7pNPaypMP
rBfGjxfefjC0SZRXm97SjqoZBQ8RLe31cMXc6qYzPxmZehZiiIkIL2yXfCYC/RtY
uaqUOi+0yvXDpVJwdRmj+doy/80y0q86SDxeDw+coPKUis50QzON3gpS6sJEcI2D
9t6aR4g+hw33u6VdcAy/gIq4b1WE6rStxmwb+ZjYZB83bm8sFvVEJDOoOGE18vrh
6N1v5WIHfafACNWdkKI6FEgInuJVLQ8fID1GQgIUf0H3APZ4rwFjQWIrnteJZYNW
kREPCY7YoSX6iIHuIofQCju7qtnG3MYBAlXsgWGHDLRa/QFaEOjW7agIwjq1/LFu
JXiCuvXGoqrEwf6RY3G8pxWmPV0/sT8RSBB3uHR8e6Lu+vgdgpRJRIxe/JNmLWat
27RxrueGw43j/phJDAwbfjZX0QGQjdPiIEo4tYe8MKn/ustywcS2QvtKCsf2Q/q8
XnrEPPHKsoaP7FXWGVAHo+ECwH1laMJJCruhC+uhiFxt0pP58I9O+keNDTFOWEPE
ithxV/AiZ6CqOuPSE5U+lf3FvUdd+r6EXExjXug4NTQPqdR3X4lqYebkoqk5YVZO
K71oFFyQWKV1DPiRloZ53SUUoI1sEsdN+mVVlu1WZb6YPZhdPASo/ANcw7ZXhaWt
/ViI8bSuscq9J8Tf8OXs6SXXov63leFfh8vk+F5Wlb/lcb9F39fV6bIu4qluOtgx
Ew9xMRkFi6VUSrQ/tc+Ie1KKuyiqhwUW4IvM09CPqn9j3nJ/3Fiuf8qlBxj5hIqR
xQ6vY3Q4FN4yTGTkjyUA1L5HCg09ZC61MEBby1ic0uikxqjmMxRJxiPDaaBnxZ+8
PpBT1mQu21RZzoJbyb/gfWHomCQDsjA81FTJI/mN35ojuTeL+3MnBJO1Jq8lyT8q
N0kRi2dyfNKUGFRtB/oxEEk0WovvJL6chCmgFcNffjLGVG1cbOHlrAyi10vvdssf
b6XLsFikaRBiI09INhQY6LIH3JUQfgltx2WfXoUTx6RXEhmBbeevdaP+MjlxtXIv
+dAvxnB0MgCJ6tbsektXTPOgLq59SeeoLMnTX0ignKj3jaAyIvAfdOV3SKk9lemj
UalWOnS/2DcZwv7Z/jNaDaElct39l+S4ektzPRe6YpPAnSLqwJxX5kxTZ83TNC9x
mL/4SmPGxfY0MYJ3TZOZCA9l8UN7q777X4bTsKQu6XSsUOHMAcLbkmWcBpBJyUTS
hUAC8A1fh3epVdizcQxIQjd1D2XIjvC548pfAfHvav1pPq0WfkYzTypmA6yVdbVM
axNKzFG48JnDv/cSNrjzFbWAm5z3FRHelNxN0mCO8/uuCFIv9aEe4xEOFqdk1bbg
wxnL/SRbCNFezdO/8vzTKSiSH+81VEQUWwzpP4EaePt7WHYOs7pIEkQ4MvzVcxki
hMlWrp+geg9STDLjuVYrP9CyJcSofHx3PDFP9zQDLJ5ufC5ldlWIv+EWPnnCRGbi
JpICiF26u8ge+GATBphWwIGw/v7fZ3F5mkfTspX80aMtKCXVjht/I2CNUCMt2UM8
XuIu+N7jAPCo+uUEXDrHAW4XYwHjz5p8+qrb8bys/Hgc5zI/aIeN+OC4N4WCvs5R
s/DNSIh36CqpNcPoTyWRAKoTmMTN+TIAT1338QroBuoMtDzL0LlvxxQoUzvbeJ8/
mPZp6CXOhBFSU48lCOVkxqgVjsPSclItM3bw8L32E47ZvonXoizEcGn0DjyxaVG7
2IvrTUAEh5aYPIWl2fG/m3zR2aKqw8fcNVDpnsL201NYwl8+lKmI8qpOKkV/A9gy
CI5eI477ntVGvg7MdGMgjmaVbyMHThohdGqNRRxGe9BFsE4lbO5XHqiNKgXZowbI
jXcu4kCzHUEC4NbJXc21gneEXqXHR6nkILZD4FkBtTVNm2Kd3uUytsuZLEM2Qsv/
yawe8Z9jfzZQ1R4m2AczGZhuadeZSmlfZG4CH9hK0BLBJuZCnheTHkd3ZaZBbNIv
seNwRlfvJ38dhbgtEsRcoJX9CFQ8Yr5PtTQQ7lXAaTHJxYvrTREZ28FkJrogYTpS
qca3mCGcU8VjpX+NuPs1zciOmtHVZC1Al+8SF0EhDj0g5otXHnyBOeg3CYiVIxDd
HfKfpWbHSLJTSKILGPdS5gcrkG5QPVPZwItgU0W9C6I87ICYNvtS66QAeR/NovTe
cye2f6SfKJT6X2Mu0sulH14TEMidinlPaqTV95vHSC0aNrW/39Hv0SyMysoCtLDF
zy/nZYrllpRvL7EiVvpe5uCtEgpNRBAEaAtn2i1OgnCLE+03Fe/C3riMCDNvF/4L
nPCTxn2rFWPQgC3zZI/otizh8Dh8LNmM1g8gOL6Xm3FN/PZTx2vg+xE/+qFk0yG8
wDXu9udK13ENlkxeQ6iFkkSBVXH4dyn9UdtbWR0j5WQxha2da/dUlTkc7YATc5fC
O0NjpGdVCpqjXClnCVixKi70zJ2qOMUyYbHo/xkVeQAV26v36ng2bSUzxXyHZwml
9IfjisXjK+4cXtVoIPnj2dP+FQWAwoQY5P712xNbLgIWlqq517pVmroes8GjxWvj
Q1+hJRbxZ6gCf0cHGJptmoyRCd4e7lSChEjkgxm45lAgEOrnedCUu9Or8XJqj9Kg
sW7Zrd2PJSyv/nUW8xXmv8+6DGPlcfk73jtuCNJCB7YfKEsKGLNIATexmgS+E6xA
y9XuxT5gIrdVFhO+wILv1N2xvgGcVMdswbD95mjHJofsi3kOBMqKHHf0zOnVciVo
HoJhPiFArXdq+GLfEkzLR1wyWhVHHFY+aDo45ZjPiJtHpZFzSmruceOx7GWAMDiy
BGbFZgz2iFZHr5f5R62QvDfu8aWKra37qjJmnKK+dRpx6i11vLO1sKBjlCul0eWa
YH30a38u5XCJ9U5wILP6w7KGFijOM0PhLRrpo9nTiK97UnHvws9PELE+nt3hmK/2
sGYTO/SDMmJTvxOQOSv4tkcTC4b8OmwRqXsSX6mA3lpI69w8ziR/XdVKzHSBPvAA
A+uXf8WIDxgcaJLfoiqRjIAmdJnUgxWt2hSmYOmmbF66XtOGqORWYy766ixK25Fs
b0HZJ5LGErLUgTuIP+Yf3sfT+uIux6FX+twQZbV/sZz6WH7DoZbCndoGRFBoGZkX
oAvUYDMptgJpr+Z5BjApif3OghSZTG+bQlmJj2w7uygpTboYM+xjtnInNCxXT5Sw
5qAtxBXyM6z4lENRjWoI/ZVkM5EhLFE2a9SNSPhrVtmGJ5e3nwBikG7HHgj+qlw9
zJpCBorezx5ktaToD8Pr/gt9siOMTgGQ87JYU5rFaBT5o7RV0TmpeYxsaKGBbGix
fF1g+4+7TGZmSUmslCcWhIc9C795MdedAgVnmhvJogHrh3hAUp47CheOnkulG1Ye
/dli4BII9BOFOrHImW/JSojxoE+0HA2mjph921+5IjH+fgu09nRki4uS/E9rhOGS
vAw+9JnUmfiYKjM6zdHyBZqWm2YZXvu51xf6Ox6ZX52qXSmGr09H1yF1DfzFNCP6
7MY7L1OKmcrRJBJloE7hlND9xOaMK+8vuCAuDXhSQojv4viQP40FsJYp9CxTnaPf
QG1hOxj080mFNm1PgJvjcOAsL6nOjvrGQchkKeUSeZMw3KTQu2dEkZf7tutVnR2J
1Xc9fuK8ImwQZgRjGWHcADkb+x16sjaNY8e5jShk8514BWyMD7fEPYuBsTQOLtWf
QjKsKNsQGDV1nKj42TsZsXlKy7HvWhddZF+tPn1Dt0sVr3R/Po4Q5bnKvSfj54S5
at0PDgPriwyAzuqymt8OZPupD6LkdWKlIvv1nAE26ONODZeuDgj9sz64b5rPmwDE
LXMIDgJJqUfVOXv2BI13rOAvmseGRz79FQuZIobCLoEMwWr4KuNFLyE/2rdndDPO
lLpJmmooCbDCvehJ7ZTu3IQc683j3Q3B4MjP9WWkFWhzR6382JjNr3T94lEAfn23
nyp71Vc0AiIfULsLCTeoH+Mx16oOn5P3TyiFRZQM7iIdsykwwxJO7qohbPzqKTK4
I5jbt74rUFB3p1PoLel3NViEYjUpudA5KMwUdkE1JDu7QQ2qemc7eRhllv9psw9V
wEEFGzmOWsUKHI5hAYFOOXJKg7djV8sa9hac5IbU66wcAVFxIEK5/qm+UL5cCEAe
LYSm3algyl2U9GkOxJusYQ9VaZ/Q8+IFIpoXqwNcWCP+MPCEke2Msf+8GM2hi5eT
2hCl9cqr+8TfjSUDbeIFXLt7LfX5A4fOlniWR6q1Pc28pdjNuzYfWQ2rbPN/Ttsv
AZKzDEmBYncXqiBmVUAsqqry/RkKJwaC7IQ6w571GyluLks1KO4wqMI02hniT9Jn
Xj66r6O0mKRG6ci420JKu691M02YvM1eo1rVzpl+oidxTtLZKKdmQ8YRqtSBfj/j
gl9fNVjVV0y9txPSugaJxhfLVwzdbBtDGjeFs9un1PHCBuKgJuKK/k26RhrwQV8y
QS+QvAePE37yo539Wg4dTL+aPBKJziE3bt6SeHiemRyQnaSk06I7ws/MbZSHxEHb
8PiJLXZEbJm6zyTnmksOXcRf5hYdTbI2JSS32q5O6r82qz+ZjbQYcQyZRuWX69hg
jhccjXsjvF6GZ/e2orvXwqlie8J+Mq5aHQcRZa2ywScF3aaD2bjj4rc87A0LU/uj
3fswLmciPsgiTdsEAjZKKHL0jTdzR0cgLI+pVaCuuSE/ZAsujYhjymhONecsGhq5
MHkvNHhEeKavcjvgJsQfzgY9i4B6jJegykT31lj9pflPlQqLtiBB3BKi9rv0hY63
32F5f+roG9DPEcBnqWRLCs76kOJK6V08QNcjS1sr/svOnkY+MgUqmDdQ/s81SbO5
qTNrweaJk7tUN5X4DcioKjFTzloIpMtPnb3bGZgLzbHMGub1L4oHfYWSS64XheZX
/Ep7xAhljAetOn+UHKRTVgQO+S8jl4JAWnkNroAWYJpmoFzR4IsE4ntP/OBrzqfu
ICvRt11/96zEXn+0+h/XK2J3mr9p/L3dn9wm16NdeQsaGmZeSZ5eQ/lX6ejc1d45
RqqoXva1gbHXtyH16EM2LCAAYhmMfbrQLKYasiYK5XblTo8gxWB2MjzoA7KxNtEx
L8UiZgkYEqMLcZMfmyGDPDv65LxavUEKeDzcdwamL3pZjKWzsiW80+9W9upp18b9
iS6psfb87KjgePaAt4LmgyIytEifEWuEKMj67qKRHtTt5mq6csJKcKrIrCiNGrFb
nz1FKpiZkrcZcvnXDv5WvF/ffwhjqB1iKxtFQY2Rn8OHvtvsjCcLaQ+Gi9kMqeeE
vc/qkJWWbqdmSK/KQmeNk+6+FEkMrtr6ZIVdRG57nEPulatN4Dhi+SPVvgs2v+kU
uXXCp1YGAZFS7FNhuedPdXnGxH2MdTnhhwtDlJoEvb974ZXEwVGUju82Jzu2jdFW
tV1fM7LBtmlmBYFsPhE3w7NGuAcPRLkpcSIdlGU+Gb0CtWnJfwTZNq3Mbm/5QW0Y
1LEw/ackINP0iAoUZ1n/j1BVAaYX0N2+Z90SlJfZvnPCOtrlvIjJJiaiir+FHaC3
QStu5ubCgFdmVkiy4jSghGVDZ0Gj8GPtrevE4w1VBD1UrpbyoGu7You8SAkxusQQ
oAjXM1DA0PGRc5mT6wge+5bFz3+IAc4FZ3BmcIWTm9ZjxxgQVYwqVYt5SHzRlsB3
4CS9ZNUC19grZ2KRMLb2rQ3S2RflWiYZZf8mcro3NT4Tt1jQaVQPZs1WJ4LfYNrB
+wkPBo+4EGVG35bFEB9d46+BBxUiye3ZQS4GnaE03OzNMbnzEEwN2dawvMf6QQRh
8z3cArlnFWwSTMwhkUUUj7+1nY/ksvvlkrU9d0uGPB4s3M1egl05sv8ZwicBJt7T
cPbjxovqeruW5vItMdnWc29aAkhUtscqJNlJyounjESDVVW1o5eiM+cCvY8lhOt9
zQvujkMuvRLV7qyw5O8fW8GUQC5Ulr8yzJy7SaZZcrrU76wxgtVXUfu1A7CDO/2R
aFbmm4cJBaq2Sz4564DJWfho//smyBKPWIO+t50amEPwdbup15iEiHjyWvjC9Njf
RoresK0GdDURCyXa4bZwa1KAExf6WxqfwusjNtD5tAfJEGTqb5gQm7Ba0RbIsmZY
WHewi7t0PwxilETvG6tqEqOVPlgCpXTm03FkqYbDIf21stdm+SEFIdNUhCeOMb8p
t3wD3eEmYM1lA0Bk5ZZeaklhS0coY00U/+Ww8+TK2uXndH4dhueyl9epBLtNoFiK
tPRbIX8Bv1s7/T3XIFQy73uq4cV/9Et1m9jT3KJvb86TJRxuV//wZjftJclpOBNu
qRbfd0xMkIEaPwlPfx2q08mpaeK8gKlJwHa5xZR1OOlJPOfVtBscIHe67Ln4cayo
5eGGpMNRINfCKPVVT3Frw6doeTRA4OfOkad1OdqXg0BTNOOe5hLjish+UyYkyH6f
F41DgSfl4GkhQ22DFPjBATvb6d0w1W9rNrcHpkeJrTooht5hoXfhgKcMagr5W5cR
X3wLyra5hR0K01EjBkwL6OCQr+XP6rkvXoZ3NdqJNZpa2s2QlmqB19NQ9OCm+1l1
WSH7Xw1ui+36tJahZTg3OvALAf/rd6MQYxiVTcacVggG2+9MqdgCv5Fyx+ZX03k2
qk5wDLo8hK2DpRHaKZ5XI+6lOTNO8L2B5MkmQcYIQJH4MgJd3ep1VH10obZ/i/IM
eKu06teG5dBROWf7OoaT2B3k+0L3RS5+cDH8hwVJ1YlEublL+pV2pcMRrraEkB5K
4ma5M+hY8PgduamYCrFs4Vnb3CFJTKhhPnmV6ZkKrPiq0nPOrFTNwalia1hirlaF
5PPaihT0K8LXOSlLAG8JUiWKO0hIHkXSdcwwvxLNi1VLsXCb55QdX99WkmV/A7Tq
/QrQWQXya2hiKYoRmK2u0BrGrLfIRVkGeLO0uGjIEpeFv0SbrGc6UGVK4mTNHQQy
qJzfvDSvo+Z2eTaoS7QfMet2YYNqBQk07AA1qt8vY9fi6pMhmft2g1kJDzd/FKrm
e701/JzSP/0Tyj0ZjBp4q05jRp5wTgIbpBGHoBWobqIwzIigZB6lHq0y9/FELkwe
UjUpXwgTpM/7mUoVcovnTApiClW8AzZqNtXEyg6+/ng24F8JLh0oU/FjM2xc0Rrf
VAm4fX79b2iW/pYKBJqFqUPwPjoFP7vaFHIlDy0mSwHYHh47Sx/gBmSCg4ZCkUz9
g628AslnCMqhurkX70sPtY7w+PIgJgmvhRuSYQ4Z/oasmlJNjWajj8JKchJnocrG
X88WuatGgEWMFYtl8jQ/tHwCHHI64PueprcDplXRLxp1RfkF7Vl+G9bxp3NqXIaK
hIsobRE+br4pC1BP4Y0uuCIgjWN2F9vUE08JymdutfrumwczHQmkD4rpNg7mDA/C
d7yqwh5J7wrh32tjNxPGZKeHbLjzml5LQQMbGKgVq0aEmk7cyzgFniszHmwUIZLU
FQmlhU64LDYcHQtfMafN05kDorwpFXrkJCpztqNDUdEM8BEaUiMf7QXeJXfc/rmN
sv30BGamUA0pFIlq9iVZasqAa5zmOyG7CsiHI0fQu2c0pXrLu85lD4i1ehTDdylc
9GCOiQ+UH57Q/3pdiPGjDz40tBaiLbHmK00n1xxt7im1JEotsbvUjDog/zxLzaJw
2NO1uytxscvBKR77sUmxKOX4W6O8JeaMgbU4H72FoZDmcDL1E4HdeflBTYgotxzv
SA0BCE3Ktd8qjk0OcjOM7sHK4rlmHC0v5Ax/9SwfUimWcazNj74/jqCGymbn9Jsq
NPmP2kRkEVC3n+ZonfyoGFa0X/Qw10TxO3MHCtlP95GFZj9QHFLjgnXmLfVWBG1J
S/uMUuyi7TKKWZ4LN3auyHFpEffNbAGg4aS0hjwOAUkFt+nEyEHa9gpV10btDxKo
pO4+GPahcWPtAHLvYtNstTNtDc4gnrtN8Ue7sj3WA5+RXsVRkJZZ1zlxfu3RHfG0
iAkB9xVshTtGjCvgSJ/G/3DdefeAYX/qgrPSPcz9VyPDxI5aBgBeY++gIYwMG/VP
Kg9Jn8/vQpBv/jMrlYB2NFUArck9e7Wm3BAkX88wXcexCmK6O5UpibHWhGDgB93i
phhFoH/nYWG8UCsYlODmxZ1u27xJ+VzuTcIryZMOZgQdijK7V5hl+RyGSDgJdCtY
6+UA5CoK2P6k1mIt7LHlJPLiKPmfj9BJEXaq2VG2xs4shywfFQSyVnNE8+il90Tt
ma+UmrkriT1eiu3aEOgk3GmLBL4NKbr1wdqbpJeUGNRfPQMyHRlEHoJBYapJKehl
Vnm6owhftfY6L6mcxFcmeSGnVCiZoWdXguV9mDK2v1qFyY+t8XyPWQpGukijrd/z
FWEocCpr14iejqzMdXTvlwaM3a8U9MmYWsv2MeBjQlybQWzo91kMPl9zLEsijDk9
noPY3TB3Y7zKnF7vu69Zd4d0azpMsrHztLnb1jr8ydwTXZ1IkTtzkZ3caLmkxR3f
yeNEgcNYL9lfj9ZnaCwnM2kNStte1pZNHKLRfTrcZQXEDj94FX4RxUUAYVLEfy3I
/GHto8MN7EyVBsvsh3+82Uy3Q8WEsBaZvkh2JZjtfL0iNXzKIdo0UoO600NBPi3S
BDgD1z20zqDkDoIy360EzRfRYYnBNqkeVdBGh2tZgS8Z4c6pIqmoSfkPe6EAuO4l
clMyOlOP8thz9N/0s/NIge1xCWNpx30h2NJawkqH+rRHONSX37+9TGGJkbU8WtJy
uqWSf/ooQcDd8E75B/lpJX6kzJ0OV6/i0eJw3NJVScryELCUioo4Q51yRqX7hh6A
Q8HNXJGwiQsbYiBz/p17D/5caiUdt8Q87xlcokKzsp1cJQVXjcHEcD6KSF/hWnEM
Kzwl8nzbuLC/FCzC+bA38TaP9T+U70QA2fncIAqOezhlmfntM2jSglcT104kMcud
CtC3IJgSBmuty4QZgKR+nqZDOAxYzVPuGIIuIvWhX4425IKA41KtRJXipwqYgY/k
Y6wyuTuXxiQvdUvMuK14wm8erXv1hWTdvwY/UjPLU3jeETlMS4DmufII8yHS/Yxu
TniwP/q4hJRsXxx2svtt5Y3iHnOQ+iVjNg16WCvABVuHo0S3Oqyqoe9SFqyoTKSL
oImFswontzbvZpxtM3OkRjlbFYeQAzndZ+7pGrnMVFF4bYDNFFAPA4DeMYiZxC/5
cYI7qHBfxxNfhBsB8//VJp0iBbaxg1qZMwLZhY4GXFY7F2Z2FdLtkVBfipUQWjH6
UwD6Az/N/AjwKACwqCEnD6YMiruzfvp/lPq6/XmTZHzndHLEGSfeFoYmrF5723aa
ORNCMIxS11AEQGL7k73Dxc4L6iY13QQEsiG+dzJu4Gj2Yzrx1TrmQysM3TS8PjuX
rjrR0kwLmvNt5+94O99q24RJUoYVtj+s3CXqVfjpOcU2yjq4fhAtJxvYe8twhhd7
Vbfi2vglj6VczG918JgOEsxyJFIaXx25huY5DU2V/oVYrP8NSa84aVRraY6QQTAA
DcymOkjrEEYkGz3hILwZJjZviqBZIV3r6TGvHjXl/7S3pY7pvtBZSroholk4A7Df
TQDMH/U8P/Of1M1nE4ykTPBLbHA+oAmvCKgxzsW+C4HGUYlA1HdcSptnXXd/MErg
tXsRrA1NTnrwkxQ9kb5JsRaE/1+IWjw0/cx91QF4MqQxtT/DZgAdL4x3yruaVcmk
WRG+QrGg1a9zeQs1kcijqcEf6hlVPDkTOmXGcOqRHLfu04a7J0wxE/VTNPXj2W7k
avGt2t5gUl0RyNwatEcpn8CS92y1t9IcWEx5Ovs3rUlWW2CvVS81MRyCzrmLobz7
GvVnY/L1uYhTimfhmeFAim6c50SnF57NNyeXx8Z0ISJDe2swxGtTCtLVxzf6x6db
vkxbiyfVAewfIRW+RsQuIa6nytso2jABSJJudJ9eCPaG8EYe+p+RJoCUsErgyw7p
zgxv0UMwjbJ8s3c1RsHg46PRx/01Rr0n+eyGx3q6ThYsfwYcdqIwCw2wJVLl+zD/
UWwjpR7/RE5EZXhVyxBpq5FjnudeybnRJQBfcGbKVPX0jOGwy+WuCTJ/o6Eo6gX5
OfIg5s5Z9Ik7hFY6VvYkt1Qqy1yLncVNnLKhLqEzaX59/AcmgrLs4QPy5P3PSHxf
JXapGxwgRiSdI9MvTFYZvS1SXHqE97lxtB19i+2EzXCfwb02jn5WmgdmKTy0xpj1
wZJKXoSYUjSqQ0HC1QHFQZHpiFhSnmWME3g8ic9+kJ7cFofA+UAmT/0EWoiwtuxl
wyXm1Fk47lO0DjviduRQ639FEzvbzRq/WHIm6q3MWukYXRXVwbB2glAENRF/1XuB
IYKWBCZFDr+/JERCcoUF9HN2e93UYdKzRNlaidlS2CxZfv08ss0hdJvdQd3r+S28
p4d6HvrhWWdqObPvDterI9ARx3srsPeCfbu/STUPodNv56pKdwKDEDiqgLeia1bm
t7BauAR8+ZTpInFAVIHekSqQt65dGFwFkKyHQEuZ1MCdEjG0QoqgQsT/D4eOgZLl
8r6jjb8Nns84CnjYvWyLifCRzDSBEW1TUuZs0ztzS8KjN2fqQzVp1yahluOP4jsG
gjY1upQ0Hwn6VbuAcH7EUiYDHxodLdxPLBrxafIZiktZaqiWrwrILLYaHb5DgGIc
BfR4yrlnDn9cEWukFRVfeXyizOGSfNdX9Bj00tuUsN/TuO1vF2Mho+zZ0HgICH9b
0dVOMRvlKEUk5hqq4RIR8SLC+gbHDA+zi+Xrz6r5prGiYDjYGRaAH384hseORu12
iR+b6MbN28PsXafbHL4fcVTvX6Pu5FWZ8l/bgifF1WpTDfffvHJW8vSUje+XxRzH
DYMTu/lfSBeyrheFAkURfsoq/RCtPgXbNQMpKJXAUdwrKhvcvKe3frNcV4M39HbT
NM3yFFVYaLc697jQO2rUdHRuY+BawVoV6dpOr/Hd7TvWv/amJJQbK07LBImZD/BR
1QQR8lBMvqMWleTY/PMTi5YAJUqGw1G9pN/9PVj0g57OYXGsoNhx+DaJpjGciPPp
+HTjQSHWIOtgzBOTmQbz8eZpmNX2TbjD03byt++lcgnGsubKzVLVlXotELQLZVtq
JJkF6ElRLp9vzP01Ago+F0Bs8hZrSTp++0aLCL+4o3RgCxpNCQkIYmLwg7TBMrao
mQO8tOEonQpqpWTM1lqGpw0kBdYLc4grztCe8rZAs02cS/LSN6RqOrfdDoEy5Ya5
stFbVK3Nt7Ver44kdfjqFf9+NRTgIKOY/QDUuq5Vm2cS0FSJSP21nDHG/YaEB86V
y8Qej/GiP6xJpTomwy3g2ptsJLAzHn3Aecb/EA7oiG4P2ARo9jKRpM5d4WthUqE3
LJwSIBIrRlpzi+RL6NbWxIlpJ+S+FiJK7zq6qY9dQKrueuSh2I/VRt8y5+3Wcqo0
KJIeNo7+7yM4B04nO/u8P6tqBCNo8DZiyfwFVoE2pNHWYr+4t98eHhR6TeWL6obw
UHZQI7Vk54g3xReZ/6YtKti0DH0J3aZErO0mt/Qg7Q38t4ESmhGQmHbtaaEst7u4
ZfGEeSRHD/f8/mq5OjjTb4gA9Mhz3v0MGevufrAfHhTO+xyOW6BTlqyuQALWs7rs
8quMirlh8OOOXjwVgdV0DUc/GaQf+QTbLEgnFEvE/AjJAg+l60bkgDwGeJNArXqI
RJmBoMd5LtdTW4rYmMZtwBfEG9RQLqY0gNO9FdLkRCXdYSmjBP7hgXJZigGmsJXO
1rQcPD5XQj7B7LQE9OX9HivUkUUUoc/BchXDTQtdf2qSjLfHFHgTE+h2f9RmHQ1d
JDa2AsqunNK2TGE7isck1Cf92Jbcfe5O4ZPpMioQBMRxnvRJbQpa7Vc7fz6C0bQd
H1iiu3oMQ3ASqAamqTTdIshw8cHqyWVgBwRwpEnS938N3J7Y0BJOrvrZgfEsDDe2
rupMC2P6eaiAD5YULI7k5yoo8QDCVZQE84GjFjmIhAaSgbB0VHACZvQqZ1KuhOW8
yU5WHlVBncXT/9ojA1cEa/jNgrZVmDMMtD+tNukbEtfNXSxT9/pH/sjIUiDYQ5uy
AlcZXLOIVEIB5Cv8iyn+8IoU0uKGHscUOZCDEydMLOtzkz1FY+j/wAnaL0D7YKor
W+qIYMwMa4mWfRnBAkCagGxFTFFAchodeEz+x4IX0AYtiUQH76KmUtH2HG26Fdpe
SxDZo84DtX79D9qpttJvE76w5QUzztDjRRObMQxfg8v0vmQJSyjZPa5UL0egqMi3
j9i7TZSMuOJkeLwwwpsZsi8gCenyrkq3kvrQOpwJY5xty8T9g32H7xD8WF7FTn83
ep5a1u7AZK3h8v91S9jPuHm1DyAB9Gy/9+OXaKRiNt1x7rBc7cqG0VUGwr1BgYzG
kAIHXrN36Iw418y3zJVKZSFlDgGuxUDe0NWboNRE3doHR8mESkKH0FP3oJoA8wS6
KKekt3mmKQqnKZutJpJAhnxBSofoUvj+clBC6YMzdceBTkQrLu8B2Lco5ppc8fI/
ka0l3J5D3F0l60vVCG6DirdBpr/WNtxv2DVj/2Tdxx5jpCqMzSbTfJuVlkzC9dv7
HF0S1GtC0wmdfjA5w/6Ivs3vvJ4I4dfwxMF9/XgZZUcluEQQE9zhoEbo/JUWcw2U
NIkShNb7X+4qJ/9gYfjZRlq2otGw/2RKhKuPnzlkFtvVZ0y54KabyvtrhaZD9EFt
XTsZi77xm2QRf0N7zj8hSqgG72BJxm/Ma3ks5HuFwxmv26CGQco3r11+WDQVpmcS
Yl7a1TRA9NyrrE1pZ8UySx/nxJvD9zoNm4zJZkyw+euoGYdIRqKgYyt+tLJb+MLl
WOrfYxBSF4tkx9Nz06qRc7MdfTYbQlDnWVXCKF5BHNe4OoKAC32BSK8hJDZEzKDV
Y/uZ0pukIyqOsKRqReN1kIZWCMU8Ave8uHtlkG4XNjA/XB0afcSR+sFuykUF6hnr
OYMWquIv8NOo4zUCUcsKwd6YUxw6EIaJqNNBpLj3nz97HimFQjj6TJk4yZOtKdEU
MTTbQf7zb9iNA0NQUnHCvHhdts7PEsrADee5d4DaZTCsYOlehvVwGXQP7eMq9cG8
30VUjOOm0RasR85FYfZdDfLdT9mMYhCV/kt9d9L9CbXOlz46Lhiz8H4ei3sFU9R7
j65t5EJNLtLdqd/barnuHq1H8+7pHTctD7I5IFnkzWnZuYf1oAzu0fkzfZ+M5KlP
LaQLmpVpuku/3EoGUHaNKb6UeXhFLWBohHFaPAphRhrJ94s8aIL/mZ+o+I3fAhFf
VpLnZXi1/fPp1cySIFUqx9OILfd9bY7cY3r0KNxZ0MvZ8iwBVXBq1PKt48wA8g05
fHvVK2JrNH9BVpTaOqCN02gExnkOVviNyU4JGhJh8t/zO/BFMVXoDHWFzCHi4kXC
uAMrJ/1f5qbeyGSK4qBQ8GLqn/YYfTt1o/fQWFaQ27rRRX8qN7LFcBP+bOAwa34G
VDhybjf8xXM4RfnE+vfgKGMcdLPITFtgw1Sg1BSE8xIw5gPkXatvEywNTdSkUyOd
sni6b2mXt+TJdNQdVIH0R5j6zZ8A1YG8g3VWJ5YDxSbBYdl+1wraqDx2d/RgE6mU
+x9yr6yQ+gi7efh1qgEEl6KFQOXJ02RzNuUwXn+1rsnt+SNfMLOHaw3K2mKyqKvB
cPk1cP/i9isxRUlVN/FWaCAPMqappn2Y7mQ7khyfvlaqIAUCsRra2Yp+34mAyWVV
wgsfHRMZdomTPMi4cmGzg6UXqy2cBEO5ym8y4zrAW1VCKRWosK30NWAvb8Ea4w2j
xXA/GsGOXgzBUu21ockw9ryMdq5SWyNqjDULPkP7XV82Som0NXch3uCJcQfGhdoa
ISP8I+ZMIlAzyQd5860jOGOWoFzBLKLCFvDcm+uTaNSNz8XSykUAvgFibLrDLcHo
Jg3+VhuTyfhiOzK7k1Ma3ONBILRHSvxzNMJMA9swQjwb3atO6mw5xl2yPSqik15u
riyFzUCSMiaQVY9N1JniF5VtaH1CDOuS1nxMLk1N6HZD1Qs1D2bkxSYIjP829BTE
21LpAsdGgewCI9G2blJZ2Kr6NuO2XpVJRWpgvOWTYn/N7tPq20DgbENGVHqP2YvM
ZHaaKDM/gAgzdk02mDdPDuseyYiJB6MxLG/bs/ns4R5KvyTIxizyvie1FjuEBC6R
+nyoWHXkRzvwGTHXnMVSrFiZ6FwjPBku1Ah+QrjiXWL9EcE2EcZGeL7HvxdsreVg
tKUOJqWcOicjzT8oJEOsVdCfP5OQxUicJFjuZ6bOvX5osE4UgrW/5OQZlC3qwevk
q1zjvgZ3mZUQ8O6aecBfu6aZcTLk5SuiJ2+hPAHQO0O0fZge0eaC7bHGPzRshrR/
cSTuV2eojpw1MBDVeSeK2xQI0+YsNS9KmQ3F5Zo1UiRRuugHEPilaWT9kBwBs0aV
AaffFO/nMm1iejykxEmoAGOevt1cpJ173N6jZe+G9jsxu9sISPPs2r8+Q7JBC0eA
IXctMvbrSdwPKjua0iYAQhPWbLE7b1kLcyL3r1LPU7JrAL9om8An+9XSy8OipdZH
O6OAOUEcaAaMXrYy4xDqxuzvlMrJVAR1xb5YQNNmD3hUvqMrfvwQO4YGMLg9iACv
TregzoQ70F7avBCzFwwwDsmphHyVx5pTps6I8/sxUJid+rlnyuifCrEdjaCVdF4d
1DIh5qGZZBEwpJqzEhDYLKrJWTwOIc784KHykH+A2o3GdwiJlzQHGiMCPNUrIdxT
R8C8cGbnRKmT2whN2kfxIn5aH8gfblZIxwlL29we52UsnfuixNRMv03dL7O9hF5s
McYspTDH0tVbKf8cPFYHMWQdPB7CHdb3nb//u+fZYDB2KGhLrFxsor/GmPPUE/pc
ZxX5ClWhahFWOrY+4aO4zNp3PGa49nbim5oczFPTxKF0PtW+WUYNGqE1m9xxZ/+n
ntSh9NJDR+KRwooBQGz0WPekSApluzQWHVkxB3bduHDZkBVA+xjq50hqA0blXdJt
M2F3x2YaphppyH+o1AGeJZqn8wW0MR7nDCtN2yzkHt5bCanB8/6ItdMRIP62owv9
cxT0esLsUqn4QAT02HM4qnarlEQsuxV4wpPZweHRamF58FE1HMxbbdu6qH3jYY3c
BZvVhd3ujgCBAqOXLP4WcJ6Eqgl4eP7gqmlHWGgNuSYFijwCGzL4fE14ZGif15Ck
av7xiv8kImcQvbjhli6829HBTRuORNPMDSHjnk/ZvNBsqebttd4pNE+Q/mjKzv9G
znpgVUSjJGTBVHpql4OeNTSYkIlhtxMSv+iMNUFiqY/iOLlba0DVUBa0vqjZe30J
tLWa7UKRB3X8KGfRqJ9pOTN6qNLln1+oemdkBgI6UFXXPVx1Pz5urwR95TLgl4Uj
7XLvOkUxNyeeh+KqbuOyLumybvlapqPxoX4hqMfITpukZtoEomVERAtSmWS61Bi/
FbxPE2jHRKcgZmlwUOyCPN0wpVutMFgppYVp0/nPHK5/MrGh5mzcpDIq1oJFhVtT
WHVo1/lHmEI4wcuGY7W9IgnK50jz+qI3S1SjzmzrpLCTeMOUsidXpQ3WxbxJa3di
3VqKcYtxhOqJAxubDqFo1LTEkOOU8usifFw5JHKlzMNox6DWFi/KlPAGs27cHjGY
q1OaGJUQTnrE3/nw4JPXDckp6mB2R/a/sceCnW7p5HBPcl8n7n/NkYKUiEIpxC30
qM7lbVlIY7J3kxBZw8lvgnPvUStqF3cOosfXl+ojwURwoO6J0LhK8/vWG4zslozY
Rhwnn+cenC4sGXuoPPjeh/ZusiB6oLvaHQoMXLNwg59IlPtv1p/rdXaxPEyI3EjO
1jsqPz8i7bHinsfBujGB3au9YEnBqY999pWY3YVQxuhGD7E4Re9Z5uDvB7xkE8+a
fCZJ4J+6CrOgaijhvaLLa/vIcz6QgvrvndS6pUVmCodV1PFbm+z3NZB/a+AWH9dc
U+OoTig6RdBc5sfWburO8RDzqIc5qe9gjE8C3cdYuoH3N0pqlYMaGXVHm7eBcTYH
pWminF+9W/SYwQ6H1I8f0EVdX+iOstg3SAqbMnc8ZXCMxkGRI8GG9O2WlhTpQuKD
vRHS3dDWLO2TW6gdz8Nxl0HnX9oAru7AS3AEKyPAkZKLgIX6p966Ms0RfS790M4w
l8F98vEoQXeBtSaAW4bXMNOZsB5mcTPyu044VanmRHDJ5v2TWnJdjVGPiA7sT9EA
JtAL1ZKbnNAmu06rgB6iEDbtcMjly5Eo0lgnSZZLkunJk+4V1JsJN0lY6b2yp5Hq
FMB/m1Xtw6OqnvYZSXiP56OY7oifhyhTFgSQ6c1mhZiX2rtTC5z6uxbnMUX3j5Cc
0dcKwd/07CizIBDzQNpS6pvqEhhubgzSh6TdrNFeN94w19UsnBEXgqLS8w7hXvrJ
J1wPtAghdOHgRp3IVxFnpmVE0GBlPoULrtu5y7RlaHEBHE87aDLsksxlSP0LV/RR
3Evg4N8HX2TE//BKS9nFViM0eUOP4dzn9QFW1NxCnKHMrXJnFjttzhyVChQ5d/m5
o3FB7OiRNoowp+cVO7uyqpPb0KqNI7PP1tr20fMZhL8Ku0V7gLdJDM/vMIKnjGO5
fn9sByx7ld1BMRcq5UifxK29olrnTFBxL86bHHpqGXh9ZGrUAMBMSIVwZloY5luO
IQDYKcVdrteVIR+KUE+U3WszOxpmwuv2jHFSinV0ga/QFGGULg+cqHZu1MXKA0pE
/73DLTLLOpWqPEWLjz8LsT5OyxJzZs110zD8n/g9StgOoW3PTmEPEu4vFrtcFgV/
NBLTOS89sBcdyf6Aj533pSJqa8mCrTLsSi/ZirFhuvkEC1zvhK0PVKBecf45kTb9
gvd7QPHe+80EMK498Q8ZoAKqrdRUbxZ3x6fW5r1ic6PWoFZtAxD8GcuppWZIAtsT
rOaDYEUPLyxMp0HUHceglW2yG1ODp0+7EhUMGiNL+PM01c1phlX4oQebSbetc/UX
7JCi9G1SBSNSb6elI795jyh1k4jkJ8Bxyi8xrWP6OuLkgSJNGNwqqtT8v4g5FIq9
i8fj3WuP8L+1f0lZemhkk4anRkizfejgb40ehkjSrG6nKlZyBzyLfMXruKgMwgft
ncbSM4D57NbHmx1B/R8LbMf+kxt66rMmYzr8WafFVOGmoJcYf6pSv4VjfZdudany
c+MwNxQx0aNQ4QkRg0ZPycXG3CPfkWp16a3iUjVjc9jd8GDy4V1KmjwJsChffZ+V
7crz8rNrnCP1BaKRNtpeeGKKVHlqrjDyPmkT5MhrTE2AMGFArtkMBlxcgCea9E4j
Y9UwnrVaazNTjOZ8XkmNS1mCbqnWO2wX/QhXMuv5nsoewDERVioFg47H3TrxmzP6
q95+OSL4SeQXYdSsww9qc8qAzagosJlOBkENzI+sSWWcUijgH3AXpP3jaz6h+4r9
7mIA84aTRLVN5O4aEoFhEPoNi973hnAtrj7phcw8uQcWz8VZUCqX28QZCahIj2W1
PYMowMKsrdu7nJBVeYkByfbQE5cMh8PsIonO9tlv+Bt1RgYnLFymucM4NW6J1Rsf
lHT6XCjKNu242sZvwjjhurb+dDXAYFgPUvHllyjG2SzQtDUhw0XL0LpDRuaq+4y+
V3UnUoDEI0ck4reca1jFhWIR7Klq9ZoiCWtPe9r7bGw9ZR5VAylpBn+RQd0d70YG
JqOdLcS6RHWr4oTFvVxHsHc25rT9gdVoZph0FrUdkwWpm1ADctUvHYem00eIAY2G
Em9KZKZL8DsQJjsjlDDicZorIbZ/2flbGIj/y2XWGc/TN7YufMk+xOPO87aSOUM2
PMKz3Z4Ts8z0XmMI6jEHcA4VLpzWdOLG5zdbz9HI42NJ0guWnux5S/EKD1viohfo
IGJ+pNUM5pI0+dFhZ+KND/parrkRuTv+RjxwWZgBcm3y2o+XOZYqT+DpTqRsKgo2
0/PoJIlFOMTkjEWWEH9GHrsaJpi6zNq1+w3YcYirfMnrl/mG65ABufPGlb4LBzfs
kzk274wrdof02yvmKhx5IkeKX5na735c0FXmxWJeFjm0VtXZaq9JkdYzjDPzBaUY
w02wLaJiOslqjDE12nNXiu1UMQQtS2HxCE1pXlAT7hcp3ShBurndMufvHPJGxcfS
agBhLxnFo0w9YnG1kaJZbhzmYllazYqmnU7+rSRXX8cnjcgHECZ/wYVuh0JtoN15
9P0vJoKSJuwdVygGzmx4YubFJzNXXkSp7o//akFdWrWxlapWuUreburVG9fL3a7C
kQQbkAeGgEvIUweW55Eh73EOANSpblsciDm8dFNzxtc0lXVGJggrIbxxzOJX1e8r
YTHa9GCMO53ufvIF6669r3W6wEdNyxXJr0XsitTNjyt5rb3bT7zmr5HzKQnYGNnz
8LX7UWFlEzYj6hpO0fFQZ2Rujw3W7NcFI4/vbuAsgGNbOKeTQujricqSHJLbaNlz
yX+pvfuhTxidJKmv7EPBbdOpgxwxKhH0fLMCO9Hxfp3cMSWcmplmZQo4nGfUIjCP
qvjUqN2CLVPDtwVFVvQW34h82Hbl8xTAOJANSQ4M4oO0gybp5w6HdqE8tavrNe4t
gYYiH56aX5iF6qhCDohbbL4xRfQrso9Cw25oVD1YYrlU5oz9lksIGCHMz0vYgr2X
fKzrGmTovzQSnylTf5i2hV5Xs/wm6bryRCPnxTtTo9u5Q1nhWhLhm5HRgRjlZX0S
7FcwgSgmhkLfulo93jKiuxwtcy4WY557pz+FVSZoxilSj/p7htD4LixF9usb3SYF
wCcfS0GazhxunN8usWGi37/YsBYjgWVdAXzaviEQdP1B7gP1FhkT6G+YyO02T+od
O45yrFaWQwxWJXyahonUYCjMqgNPJtcokOY0EZ3/jl/Rgs5kHvEvHE3yjJ+PBZ5X
m0ExIqyZCiC6Btr/EfcWtkYGjuBnjaU6oBSexskU3TuUfCTro8AI7tAl5N0yi7/0
A4g7FsZFH6ppjxBKxi2MkrvIdjMiF+HyrBrXoJptmfbu2RQRNPzrGJidTVPBKdQD
gOZB6Vw9JzUg+rdJGsc94vCqQQ76lOtAqOtwZ7UdqB8ArwfsdliO5m5cfkWA91iw
5BLUtJ8o1K6gJm1okE8e/lVVAt1qq+HKu0csuMlJAXtz8nmo5TXFOym9cOS3z12s
olsZ33XPRx9rmV4DXM4EgStfzlTQrr2Z3uCKdiF2zl23bm669rF8TYoqmb+nECWU
34X37I1zTo62uKrhlA/63DN33uq8Sxu7zywJpmRtQH8GY3fdY/m2ZxhB2OOty2Vp
6Y+QRb8Y6WO/EoJrjZG1Q17fXfx6odg+ADrbN9iQKFOy9N8hcVIhOKat9cknan5/
ahOthT7PKHPSVp0DgXGyYklkujuClwhISLyBWpgtBKKs9pd5kytb+rpbodWU4Z5r
+HRAJouorapr+p/Ya7pqE+FmryFrH0HzbJ6N89t5ediAp7I31DOFNIIsUqRLpuQp
uOfOKsHWvESTl8lC84djNUSD3R2UFNIxzFQJvcSBF6c1nX7yAKGMV6UNX9wKiAX3
EZv9d3zQa7vY/nx2dmZgJmEUxBdcSWm0/jXjTxO7LAf5S7OjkR+Npi6XLtIQVn7K
Lj+vPNeS2g+Bl3PC5hSJ5trsPThT8XdtlnE3PYYl+E3U49siYq6PImEzixoyKb5U
UcMOedHpmvJa6m2linxWVzfqDORFLME1twr1Q3KzNt/G692gncoYm/zLwsmyzF8F
PHwWCkcWD7wBcw8x7CQY7IrugBq6liuw6hr75x6cNfhpYZCBRNXb53yVSvntljwE
GaY4bkj9aBPU/oROYmPZ8cD9h6ScxvWRrpiv+ChyrZ9JcgPY6V+gD1uxDGt9AxLd
t6vZir0XeDq11FNBwERdeQnBD0nDSLFAIS0wtAjxxk5oJwIAU80YjqIpC8kLOcsf
QxShtwt75mATeK6B1/XhvfTsjQvRiFd1MV6eQLmc/0qFv3crT84TV3o9Mx46clUX
8JoHR7uyx57tDbjEqQ8sgbObV4yDm909hNtPAsMD8sF0hUtJtAL71lb2pxkQjbGo
D2H8rt+JXhoAPDB6Rzb6/d99BHwkKla9EJeL/wZRhzeLMLB0at4JjWMHrbD66kx6
+C1eNe4ixLmNyHmr05uW3k7wTOWEExQ1sSnQDrgynXZ+gZoUa7esZuZmnXNdu3l+
maHQtr8cGJFiPSvzrxiAZyPUs89Ev1v9WL+MSbRp7c5aMHSAxn+tQbTdTKrtbVhL
BOxOTUOUz04ZWSEeXS7qyZGSm3X9khoT8J8DhwxQPmOm1LLFKO1/lL7HAj+u4lh4
IkgdDE5WqPqm5hNDqBkwbUmH4SOfRkazbrkfRghBXzTjhKH2bjvZeyePrxpr7WbZ
FawlQiAtpSOl4KAyXwfKExGxfG7WsvWNVyajskuGvwxjjoVp2kbxDd0apY6Zr8Ay
dFQOnDSdFbk73X0npd0x74QNnW3ZH189N0Zu8y1pYyQnzE0H1EhBpOSaOY03N8v5
UtTpRpztKPhyRfQIrEvvfhatwf+LaQYxAvd6bhC9b330ne3eQq7qooA0LUFzhhB8
7AnLW6nYeVefvA+FwYI1FqzvlPP8enHS792tNhfbmMdzQ7nezcQwy9GPYUrRu3Su
Hm+SQMbZzWaoO2PDYDmR2aN4Xf6uU2nlK3MCgf7PTUnX1ty8bjlvlCsz2doKTr/l
Bi/b/A5oEt4dMvU++3PG5eSCxJ1WreirtHML596YSFLm5+OrtH9v6wH+o3YmwjGP
NWeIezobrz7aTyxAPgiyl39r5xW00CKDW9zUHgiHCUY50WQoGrupWkAksk/52fiB
GZqagzorfjtCcZf9/tfpUiiZgqOkQlILI6OqTciP/jq5hy4xOK5zJ1Wq4BF18qFh
9p3aqkTsVl3lXQRl6/VVe5wJmm1FKiXVUGqtstPyVAmd2y9Zyayox7DRmrMZCakA
OMiE5w/ltspGaiDYHI409OamrAYUB4ugK9F3h2NeT4fq+T6bCunGs8XJQN65qi0X
9sz3+3hO1h1ORlOwyRYrDANPIF5+oEGT4B7AhhfKLVXMok9ZuH/tEEne4VFcHH4g
VARkfFOWuaHfI36lW1YIgUBRRSIk1pduFcbNMxdgtLTIQKbgGTCti96X6gz5jrOA
H06fRsosE0cg6vT+WsvShc1VizKYrBUnN07KDssMCpiFOAacHN1JQ7gGOksOAdvX
tAPQiewxTYsiT35FdMX8wUN5kigkVN7FyvKp19VrXPPI7T8HeYbQtjwnh9T7AViY
P5qBWNFsrUAdVqMIos7iPgCS1V9gDQiNr/tokt5BbXmiLGuZjju4vn3JLOMivR3b
IJphMvQzFFVeme2D8q0EJ/qucwg9XlfVmLCkngLbc4w+e3p4HdtX/GQWyqlmZfkO
0+qACouEGTADYtTlpT/N29+s7t5kXPjPyGIWU8Y1q0BNKUzO+edYazSZUwoyPuvv
Mk8QboT8r8RjiwoGMX1LlP/4svvAiN2sg7rWA534iNo9Y5FRpBkHb4UGWGnN2PHX
/173csEtbV8JDa0e2erZSgcgksDBG19wG7Se63cLdVk9Z0MUgNDVbJPYju6XuDvu
aHiCrZJLpB8Y0BFYmbsRQBm0AI5DsT/xC1pYcUt3CquJKvjQGYrmQo177YbK/pZb
gZY5sqKvxs1K1c1pI2KTg3kVdWOF0rj/fwsDSvAx7D07PmQigXkQxh8MZV39a5tz
mvizPstluWOqDV58mnsn0RdzXMae/pzgA4JwYnjIDGmvbpBsOg4+1/wJXiRxjcXZ
mdH2R6y919kNh9EeVN/50cM3zHwew3/4BD+P2s0QpX6cdSXNZeg3OFNtTkNBH1XB
wgWtqvosfXujMNmjPpYg3nJyKG1QdwSonLt1+wOoX3oRQ97x3PjCIDrXmhiojaNB
KB3VfTJ7KhNoWrMUVfKirdcv3401hLCAVP1euti8E/tRNJb11QEHeX83ojWMZceZ
ITZgA2RsIQgM1jwZ/Mui9Y6bFvTckKd33SlN+hlOF6JIU+GgoD36x3DE56XD28++
s6VfBYw2U/JKeRzXUkuJwbXtsGFGQGKP5dPePJY9F5jM3MIeoRZrogau9qzJJcuE
L0bRBE1HiEEIvqaB/66xp695+4+Jx/jGJR0ssRn5UUU3a+bWbmx39rfxAjvKgbCU
kqw19vH96MUVDpr6HfN81/HaQyj5IxFgmGcne7sS6jGoGX095ajK1hrz9ZWQFLy9
m/Bs8ZFEJbNrypp0i6vJJKpQVgKfgKqtdDwa4D0daPP6au3WHLo6MVHco8o34e6V
OedhUn36AwdvmwPFPdgBaGBVJg0h50aAHxn0ceaONiiN8Bupm73wjM4yONYINT+l
ZAYuQnlLbgfQmq7sN+veUNe2oVN8ijv05Y6DT+GvhFrfgT/CC0k6G6rizf8RPX9/
Hc8umoxJt34FK+pdGJvX4u5nUFqq63m0pf6FKeWoUNrl9FAcd+Vh3sW+FkPs4u/D
aoTOzol4SCvWEEk7Rgl2GD17c7SgEPo8gMHmOMLMvlRU6ARJI4zH76A+GEMz09rY
jn4bS7WUafXsNYKNXpIpURdCkO1dKK0Abax18eO/hm0coAuqGRnFPVkWQATGpCzy
R052QqzP0uZjk8jpvLeG+rQRfbD4+CJuJOnleXdng79OIjC7rbz/0KmrU5WW8HEZ
HqWvfMGmKHqW46bQwdplJl95bcVWd9rSKaD5GQtN/QP1XQJGCsOVUE0kUaJMiAxl
iX1zGvedDeYi5WgEORwvmaKGwOLIm8uKmwBqfckFrJPvzqUFQEUg1ibgrTSOKsnf
pNcWYxA5wtL2UyammlcuOkB9aGKIutmF5eEmABIwTJnd/pN3gV9v44duzC7vYp7U
Oapuj46p1QeOSgc+kuLOUI+LNHdcpiFxT4FObLIiwgBHzLdCjXvMt/i8NCSg0his
s/pQ6zDO1jXkIlyZPV9wK4U+eoPzumCX1GvkP//GykKPHP57Ltogalz1IblPR4jR
DoVRvPPjQRnXUSSYCDZwaeRnE7Irgd+fm/YDemOH1PKqAQDhQOqBYHXlKgiS5gRt
tymfyUfGgrcpaitw/ft8nPl6J4p9sP5lHA3aG2AJGX6Aq6EaTOZPsW0DmNnyP9/Z
I++ypa7vgGHwi4pHXhK0UJKhlBm+ruO8SFTawyY1rKjNV8HJL2/OajSRsDdKfxwL
D+Qb3WgUm1IdfD0/NCRpm6njGXj6y4HGOtoujSmaQpXojei4zbGp53MOFWVgdJ38
ek5JGIhxIaCeiq3euxFQN1jSe5lKq3f3C9JH38t83Fa4pzXI0i2Dz+/27/jxXQwK
ukHCr6E/zMWpfDpAsgNEgvdrdxRj7rkMtbDjgTfVhTF18FEeEdHneSU9L/FjQfUZ
ZYG+2rdbNr52VQyscVPLk8OGZznvBlxLGfplghpZQSZN0i3+i2EzfujBp9ekTx1G
Ci2+T4VnfO96stBUK2zeXS+a8QMn5kDZYHtyPcvbbTCAd8fLxwn2Lu/T3+Yo4u3I
IX6TVK7KVQuqEJ8i9nwasKZpFuw1KdWJlEMIb4qEUclV/OGWDghFOXNlAqLl6K2a
CMM9lx7zebYP0JbJVMGuo75jAlLZhjB7/TfBX7NYRaPlWAfYHAQoFQRijfr0dQYk
vYg2YIoY0JtWcBtaOIXbRcnJTFjTdzRps/QNofekuOjUYIzR6cJ7oVjjRoVKC1mr
v0XBr6ZBeVuBblmeXZCyPG3OGd3CCbv+M1MjgI/x63sOmle1AWtWdVocHvWJ/FF0
y5cQPAzqCC+Ysm7kCiFV0ToJ5uMbY3MP7AgSIr60cAvinuKc+HM0KxjQuQRWOvvo
wclV7G/87nyBT0bpKs3TveCOqaxgEZKnpYhH9SryBtjGkprMQNBXa+RFIK10mzTp
cP/QqIF+srwKxzOr2tj2f8NUp5AQCt0vB2+oOYmkhG2vVv4DigHSjHHccF8MI6b2
qhKRfQkQ2QuQL57yaafDIBQqADjxzQEvR4JTzYbRv+9zDfeE1tI0HuSNfslpa9MI
qrFrALHd+dMCrm+32/SKHdpJNbO+Wmp4KyjFRWcqmfN+hDlNJabndVIoaOjEfNyJ
TkiW/6g/C8wRak3iP5V0dtsd+aBKNVPSRW63mtagdY/Xw7cAODa2zFi8tZZIT1Mg
jLmSAVhHQy4q7D1hOPP8Vbqt3lky0AQTR2L2FOKn2ZS/110+ltomnlXF+RLNCIvk
7gTUJvesYtCiR66sX74kHTrBYl21DkM79P1F3oqNln1yml8Ob55DbOg32qgN/TZG
H3aeprmKB3fETPKJxI6BpdXADov6oR/97SVRbGuZErE6FpVALsTMHhX/N63Q5d0P
9ARxIlnL6Etj6mx+M8W2WwEe890HCbl9IwP+AVIkVb0upcz+e0ngg6JViMdpdvEf
T7jSFHGw85VZ1zzB4yo37dWMlLDYARqkWSgiYXBueGR00lr+lJ8qB1z8SyU9eSiT
DPIKVa5T5b+akLKY9TcmfhNZCMdnL66V5/qW4G3XOyPHobWNfUs9CxArr+/VUWiq
HVFu920XgSInNQbLq52n6XceNlAD7CdIPXVxjgmID768UMGd63W92KYLUrK/F11E
2N00TA3WkM813NaG9/zzitZe3GsDUoanXxSxU6ItVo2fLUDZB3NHFXhUGJdJx44J
ODtsvN7H/wiqogBIWVIeAU0z2zp3BWH6C6rZ640bnFIhwU+3qOVfh99rQVi0CPSw
sHV5c9rTrYG74zVGcdW8LsXycgXCDWS67nV/ahykeNX9zK8hpAMKdrm/XRbEv8b/
Y1cWuui/qDe2Jsk7Xjm1ZwsRoYejpIZAz0hCbqTdwJiyPddtBkLKX+Puegjx9GuU
hJN39XcADG7WMCkaq8PXLbsJD7kYCN//ABx3YLSMV0AGjX1qK/oUiUcWpz/yfMer
CYd/LtEAcITHy+cuHPo4WEjjoRIgBirzNYEHJXVX2xnh6+coY9LDQ/n8M/NYtZ/g
1DZFROqw5BL6XbyhPBT1aDo82WuvIgTJWWDU3dVtNCqASureE7jhysVFgEKWCwgl
NsYJ2Ai8m33BnsfJeLfuraUwbyGGlSJhFTxC1SKSn1cGioXPXKQJ/QD3hGb8YXAZ
S5oWUSX+Z2byU2IiIi53HsmzUQbUqWztInJFY6IEa1dNpvRV7Y2jbj8XRdHmLEdW
GAU6lenHh6LeOntQOd0K0omF/xnQ4R5V3xmVHY9O2sTh9nR+0mGPt7QBc/cORecO
BSsSK2DjEeoGTpRA/BwQt9FaMDjQiubyiTRex0ebJijG7ukB1UFu3xBT6IrOvC83
JFy8wMr4XS6c3eE5HnMzveNQ3gT5+3K33MCmKJ9qp11t7PS23b7lAw4naqWojURo
fR1ira4++rXAK9gDc1WcgQ==
`protect end_protected