`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9056 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
iOS4T16637ogvUHHJHvO1E9zWyekqR6gJIEqoyePTeigwKwItOKg5Yr0rj/Xb/KN
NqLEezaf4d+DCVXhQkBpFfScZmRppd22VWzSl9I1tx2o8e0EX5yw2MBFtCCkx7Ma
KK6yKD6OkVxSJj2YWMIRj1yn+kM1ifpzJ3mgPDSvnhjDwjFBU7sJoqcKGRs9o/w7
7ICfuxlTb1dsi/hcINBfDcoAfrgOVozJQdxl0pY1dwka07EQ9UhZ2dR6SRBv4bM9
im3zEAr4MeYacvpdsBC0MlgVAYNNpvTi5Pq5VqrSGpEKbDVYKJBOhTPSUGuu6FIY
WHddtpdPBnNWJFyDlHnU6AIDIFaueOLrMmprsHMdBDcHPmeFo29dLhdHprz0Gukk
zfGB++5J04C3nWgYtU6JAwZ46qWhzosMiSRCiM4liH03tk/WrnoLHG1099Hh1Omx
n/9fxV9brkDA+ikHEb5D1l3ncqQtzaAr0JoZGDbvBjOpc8RClrHQM8rVUJy4xauo
xzkboZKznW6OKaAGdC2+7omg2cJE7PcDsfdwIgxEuDTUKxdsqf9zYI257Mfyy2FA
0WuynrUFRY9H8uUaBDs3FgeDa6NZYCbsN2krqPAfViC91YR0rNxiUe2wjAmCPRpb
+cajABjQZeCRVfIsovmOfjA/OLH38/3mmiFScSMRHW5zucRUZJ6xTCqNcRHTr9RC
TeaTtLMlONS8MuJDLwl1KVGDN3qh/Qd9UoWj4pxbuUv+YEBZwB1Zizvkuoalhte9
X7v9/FwSVZB4blPd/qArFBRneqCNRThwn7plReiH32l7zAQQmqJeLsi8jO3dHDQb
C5vdaWaamI/h3hm35aURU0sSxXucDRmkr+bJh0oGu0IBXte7cXx7tgHSu+UGUevT
tTj+ZtR2whrEh0C/DutWFVS2c2HK1Yx5o9BWHz/8USOg+JNJNl6NeJfVu12M/4uN
4UQY7RPB339Ntbf17oyunJxCbBtW5UqC/Vi92Za5XUUkp7YEvrvL6YBSvH9A8HMK
qumZkIQ5pKL8Aw3VaUzTEyl/oZXAck5JYEkTnVtl73AHRe8DeZeQMY+iDSy57VQz
csB1SsgxCa9bpdT5XF0L63Rav7YYjB4WrZxjfZFWJdCGZm0SKAiocStjkxBiZMuE
FmUioHJGJEux2+2coqS+rnnP48TrhxDvnQLus4bQdevjEXWiKUN5+tpjT7175UCJ
KuP+SgwCxmbwvWIEtXPSaKW/lWkREnx5k3tFnjZY7TaPCNNf9h7iz/XlmqgsjHOp
ajs3BN2L5ryRsdQPH/jI2vDpTM2C2RnAYC2hX97FuvKl3MFPcPPv4DGgHpA6LVsQ
aMIVC5MjnwjrVadTh1s3lthazPBzriXPKRWJYevYEpZ8DEYZ7hio9b1y7R0YtKzB
3no/WRP4RaQezwbclSy9EYmaruXakN9q6N9kpO/5Flq/FaJwf3qprebr5GPQHo8F
y9Q8+qXYtPH6KTOZN9ri7ES4F3/lAenZxo4mCOshCOokjgfsSdoOUSBpSQNyvdk4
/2w9iHNGuFhx9R8DtoY8KvRUvEU+kvlzvqPCSy6FGCy0TmBHYOLPbe59T/qaNT1o
Vi9g3D2hevV15c3W/on3qGFoyMhdyiCvFHFNj+3rPUCkdBSh23uFP23nu6VE1+Xy
ipGxpfBmYbExDVwmwRUwHwX7cbV4ho8Li8QbQfA+rgwEElG154O+8pnhxvA1Wjzg
lBaOo5YjBBcrdCRW8DxCXTHH23eeC2VOcWtvJF4+lSshSbpX67IhtL+VrbvNcp44
Kq7h7FY8ABpEHixnBQY3NQivwh4yHxYwPbYJ4rsqWZI0dOev0tBlSTAOUWJOEjNT
DFK0ieTX3DOtXhTLAlMzSjykcLYT9Y6z/PJNMYEuPY09q6rsKrZIB7PtJFBG3vpi
GdXMacz+Ri9rWNr6tOUI6cLKV0DafkjTlzmiXUfpAyYlvW2YVpThX9Vh490fgBOZ
gPS0gSne9B3OEcxBlCD4ZmnnA+R1vei8Q31TMmjQgsv2qHyRecFZQ+S3WJCy+tiH
2zMznirGAvNTu0S12XdjqllyU+Z9dUy99iPX0vrW6pexvGNkd55YegGC/AkwHDx0
WhhDCDeNbt+zaXmV2QaGNStEpu7d/wOYdsgV6orLL4DstuQN8jY9B+TljKqk1kRu
a2yusXI/1FqE+RxeRJfecgm2mHaFqjKG0rB8cRF0RQf+diZFIjrZe7fxfy1yjfSN
VA2fOOVb0Xy6YUGYAPR14GbaJKfkflHGXxuOlfn3aIO8h2iBQIXvP53BO577cgzz
lO3QmydAXcgG7AsIgOY7J+6zMrOgpeD4fsUcaAwLg0aMi9VA6Db6fGEY7GFnExkA
1H2ohXztqalWUfwXOO/KACZDHO7ZOVKl0B/txEs4lgl+qUcHE1YF4hCislHjuhiy
ptROBDDZzgdCPsSZqd3HWIB2J67UjD0KtWSKqoCdrbpRQnHUvcJogoJP/8GCgMDN
Cz6Ek6TQg0q0fQVxI7psYBcVofb2EWmlTs87+QKjPLl4IPKVJSBPyhjoRfasZbdR
DWigFtdCCLJZuXgEobRWu6E9SP9T1jZ8k9tk1zNQue7allYAmGuVxlIA7XU8QJtA
oLFGmvLF9otnO+JHnjCeFU+Bwmy5lZOpVvPpzLOe+ZfoLIV4TO9KGlGXMr4nRWG5
MVY4BPvY/Og2Z84bQSNj9fqo4/H4ZKyM/2LyccZerLO4V4L7eH8c186zyB17FOVw
gx4W2bUCTYxnpsYEmD96TmyO0i9NWM+axarOnipB3RmZWEs0J7eEoqvaGU3m0+6M
pCz72JAe8YvmZ4lFkY7u6a9p6Lumo20Gu2t1XkhXPJpDTS2KUORIidwcA2iFLio4
gABiVjrbP7B6zMBb+ZnQ0N+Br+fdv9Vq51ni+dd8WEU4LilHXNV2c6yLagV71Z/N
GtpZuH245fp8147oEwYLGL3nylhP9ajbuwBU/yX+NQjnykIUzcM/dIy8Fn4v3Xii
Sa1QoH9Cx+jr6j7canJ3xL2aDt5BqrO+zjMww7xBjniIposWiV/j0B/+Ui3tyc3c
qgLtY2M2rbcWAPQ8c9gqsTR7AOyVfg4vS1jAG/lJb+3ymz1iV8MnvSyeNypFirGs
+Q7rpNrtpbbTlrhFbXOHV7CVFz7gvU4s/G3dD8jdDWv1tIHSvOeZPhDqXz+iEjed
YWrRxfodcKFE6wWxvvf7PauKZrKYdcL6r2RPgasI2iDtmg+i4WbNiWZHAHQIcHIw
qUACTE+vAKhwTMaqQEMwRXCqnqTst5Hjgwua8nAauCoq7gqFGzNdAJY8LuA1jFXW
DdUnb0CNB+43NwMGy8YNdmpOFr+XFC0PXaJ2Mup5EKrUJCBPCa9Z4JEPyWLM3JB4
6+F3kjszhHl5vai7wC8L+Ho2GNkwSpyujM0mvWCEY9J8o5RU9CELx7pEoxlfjhMj
3Bt3bJR7XthLhdeOPilYBGStNMlOHAuZPmgx7dFDeAzu3dvkRuKRjG7RzumR2078
I+tSAFzQ01SbL2DqhET1zlCIFDtXv681p6bVS1j/9W4OMHse9ClWqS0B5WR4WVFb
hRk001PxWNkPAtbT8z3J6fd0uJhUQ1FCTtkRy9mUoL/wHsm0eGf5a+wc3i68C2+8
wPXGoBBJXIKQ2xo5XnLl70zhyQGUHo7plPrW47RuYM/8iNQzKjjCIfF6ILhwrar5
n6aojDqS5lEH4YFjdj7ECq7GoADoluPEnLuobGMsG1gl32EXZfBDE6eZVzi5QlNE
jCeO0CPY0qA6WZkjCJltpBVMy3OsPHH5QiXLvTg2DunKEeB88JwJFux1otTvAA2y
JEbdMlHYC1OMdz8Yz9ESTBpc/7g0XAAhtt9++HbIGwVa4kyLBJzWCjN3Ux1K06xp
PJTQSB6fEvxjw6TOjxNgpwUsUyw2nTWrbXDzZxQO7EZ1QTu4rVXAwyikuO0zUNPu
2zVUEpmkA0EJXbJtsPrpbepZAvW4zF0OTR6UZ/13Xv94nqIFfCEhcPKqzWsWLBMs
QrrR3uW8d+pAVGygn7RWgHTzm2iQtGRgeZwBW4C5vrN6PsPo1WvTGrLBh4y0e1vt
nEtIx9wbUOI0kCF+Xhsik20K2KPkr88TlVJH4gh4vC7arJAJNGSzKyD0349Myl4t
PiXeUYMe3/WxXaGLTvA81dblhQSm4Ma+9YN1ALaDY4JW2mPWcN12xznd3IKwPDl6
OUe3yYn4YA68TluJJgDXCcZNuHLMuLqZ59x/XIldsKH370NHSsz0i2iEap8Xz1bX
+fvjjDX1KfqMnh9JdSRSGH+h/9fczvgDJZP/hU5aRhCONXbu3qxk2ZLKcp+5OSy2
KceRNZ+4PLfUi5EjQPTGH5UhuB0UFHhdq7Ne8Va0k8LJQdsrrX7na+sFrRn1whb7
uRaB6rN4KTTQQizQPZhS1z6WjIFK0NtGcikHGL335soPmgy7tBTvC/ldZIY3O9mF
nJcGo94CmfOApxnQQkB1PXx1xy6zHYxFR0Ywe9h92xgsoVV4BVW7KXg0YsyTSvf9
gRos34jf3XSoCpFqYaJRLLlfpk8tjztmp6ddEGvX5vNVUPZrcuvYZjWo1jSUV8m7
C50J3NQ8jW5mZ2rMlo/0U2ffltbRBDUtJ3qHDYp4Cpw7AAbuQ5I+0xaSJqcwTnun
Jk5BELkuvV3Zc0Mfe/1YnQsDbZuUDXj1tqYBlRvyXcTURETWGhDYSnfwutLriJiE
xp0G5cpHr5WsZQote/nr5qnCNJtKMjOT2dCX+JpqpoMbK5lb/YnO4hFkPaXXGXQF
iPvRfTZ+Ls+OMdRu5kc5yHsTjqjChUgwYXzCXKf2temt0blCXijNbAA5hJiHkeQt
WFORbr/36qDyDY1lN9II6zv6y5wfvv59Ns779znnfocr48oDIYAXCEs/r76as4CE
XUTvt6c1UWG+dnwKXt4RXc/yqduLk1EDIfm+3WBsmHBbFFxQ1pL32clKsTYaDNoq
wMqUqo2sLvBIY0atsj8Q+PNjQo/R5UB7X6N4qPFx/FSGmWFF00PsBxJWpaCoXCQ5
tdjxUR1DiIVwd3mOMe2DnL5IXuTfbAQNqKswM3OT/DLkZ8G3hKueCk7n59skdJFj
mXBkPAt8hZQli1kPNoWxAs195KvU+GjU9F5p1lQUWcNxXM/DscB+DJ1Hu5iAe7//
at50o/YbdSudsQso0W5ZsBMv9v1MeLHhuNO84XqeeQ5QfjntOwXo+p1ZroUc59B4
hVAqAnYb24PwAgi18PFJsXniA4yBaqPeIUjRRsz6zx6+jAo8OqatDKS7C7+YNJ7V
Txyc2UFVF7DBkpD5zoOLfvkIpoURueX9fhpnW5YzfwuHfEco/PJ7Hsy9qUOopHmu
KGiMBDbNIgZ+SDZ6KlLW+vO5ZJyCNovXGgGkvDviCb3Br7+CmpHhiXEeKbOlg1F2
aSBC0LNI+BimIvlYR7J3XFQDLDf7/kOtnVDclCnP/6YODvAH3uqYSUbx+GRhk2Np
OzUpmzc7LxuByTWCd+kpAXtbDtEVLnx2lIBE7Q+BwEF7e2LsmR0cbEaSu+xuYXJ/
i8EIQxvCpqO4oz5n5bN4v1bJLAPhX7G2a5P8O04qf8BgbwdXZ0aV8CcvXRiID3YV
eA8vk15T4bRo639x74bVKzszRzriH95r/IrXJKqFfVfoAsYGbrLqVWHYZ1MLGPf1
1GsoViajTaIuO0fYTgh1yoQtsuKrCbYFWrRg4y3uXASJ3NUM9ONtxI+D2AWxLbzk
m81ZdLAnY14ut339K+3sJIl+1vTUaHrclc4/B0N5X4WyCNAJwsbaKHaZOaGyMU5n
xOx5li8kGDHyjYYuvB6fFN8zT3ugFMHIjpVPIXdj6bHzKyBwOASVDbyfnRl95iDS
jPDvbT9uVW6SzH0ZqwCp5UqhCF1//d//fpbkNYbeTwUKCAj2YISnFbXAvl9DCLbv
Yz8bI3cHRKKo3ROiS+AvMf2PwJLQkBCKGrQM3qomSCcv5sS6nS7iL7qRqqbL6jd9
WSp4jg+SAjQWBpn5hWZ226gaKTNkm9DRxDMVaR+pdV+1tTTXGHoeTHVEBmxe/uUQ
3glF1ZzNGoAT2hJDxSAhJkp0aQnuEHVPled01a8rOGhpXU3U9YwTOnMv+2XKZPOI
IQSUB0dT/ptiIPo1wVrCH2HzPaDNYajSn0rrMa8SGz13hekiUOVAVAP6A/cKjaU5
40gUSjEQwgVTUUtHENMEspMaheh8DiIZvxPg1/0dWu/ShNsU3CTxoeOcdnHW/sqn
MzE/qYoYj/Q5GYSrWyOS+Mc6G6EEvSjAwjM8Ib4iwfa5eQ6MRsEyDn35fDmWYWqr
AD86wEWtLvGlYy/ex6bStJLcG2owpyLjNe/iGJ/flRdGbcRVsZ6XQIKrFLyPhpF1
tlYOSn7kKSBrJXcaDjyHTkCNqrvhYzvXYNKQl/4qcocG64dvuzNb1gkUkJrDdIwt
ULIR5QM0ZrKNTkXHIAJEcNqs2HAuOT26qcDmSaCgg7wQaIoJMJpUEH5/QnWOFA01
KfZmQ8YhbrNOyrsp/C0b4dB6Ot31c6xjClcJTERNd43VyTyMcnbx9G9P/TET9DiX
sMm79m2SmTL629Ksdb/1fmdZtNkIRi3c8rO/DeHI9aKYJIgO+SGZee7unruvgGof
EkqY5bEkXfEAMdO62P2ASE8Y82bmBj8Qbrez201DA6ESaoxdJ+NL0p/3UgtDtrDA
yTUqqOaH91oPKSsM79WPAxqQyzlDDc8KRJq/PVtm3MgkDb1lgO0EzojONJ/1I4jZ
E3RG6E0peFIDYB+7wh2h3nZXh5PIWTPzg2C5repHwTtIS5FBB8YMIp0q2DSpwPw7
3Wj6SZwLqNKItsv+kPuyWesEqPN+Pt/fua3VtY0KqOYjxQgTNDgqtYn29wyQtto4
eZBQ3F9UPEiIBTwI9in3y9zSX9ADX0f60wpFIR/yWGlpBwDoucr823Tn07z2Ok08
sKEnDr9J+ePSeXrMFwQs3dTCSU9IshGby5ekYVjAxFiTNN3hjlaFzJIz2CgXzlCV
K/3TLvWDCZnFdGwqGEAPIiQ3Mh8U79FfPsx50h4/nf3Njfdw7qFK0Xf2iCSiaZaG
NCIBIXPy9XTiqj+JtutV0phM1ygTiQvkeUYHAUBnFplcBawc3/9K4BQko3F5tDyg
7YAd6zHtk3QldNi2obNsSMoCDAorObxIgk1P/yHxoyD1szZsh/XMZEwGioCkx7h/
5SAsJDYEZtQC7IkVIBoO2isLvl1fLwteY7ywzStZ32/ggCaPabsFKC4wqUK0cSxK
CFRGTIyqV7t6LXG/Z6htzTEdjTgpeSMwuze8i1Y9BlpovUN1HB1fLAVK1a08bxGa
hhlAcPV53JI+c5BRICnDWfFUOY9kgtA0k19YSLl2FnpPpVXbJ2qm97Ztm3lq3dUP
J7sAbmwmgdDYJxalEqV5jmBU/74BJHDPpnuboVK569mQecrO8HmRIVhBxqn9X1lW
FxXFRAyMWz60VdqFrv9vI2aUVM+6fBYmXqljwptvNr2QFP7yMEgVc9eDI1mmXaCX
YppXhh+lveapmI0DdLao3RV1foNAqyuAzWH6eUaKlftj5tI6z42o/XrIvVMA05yX
MXTdilx5m0mRlmm7p6wYVYeT5QNt9F4g6hrfgq+m8RRmMKvWlFkV8EpH/p5u3zWy
na9fTuF3p1AT6vsIvLSx6Xo8wwO/4AmE4Wp0DM4IqM/h+XRsecJhpfNptuUd3g0l
CeOsn2zcqV0xAUpvRh9Ynwv6fceWTjI4Z0hOWuIFGBCRuiJyZjqbgXJJ9FcyIneS
D8tewb0eU2f8o9J7t5Gy36maYA5h0TH1tjrM2x2Wd4YP0RbKTvfULQvdrYo3Acvh
j4bxR7cDXhFFm/URg/RwOFBkwWzv+2ktN45OaaTAxenz2PWlW5ERKLV4P28L3Gx6
H8vfjMWltEQA5skN9ZMlFBXDe4rfMqB30C24kJboPH264QcUEEKzxJTF4S1od1HH
53HTgb/VU9egPWT680LaAuHq2IPh2q7dJV02mq3WYh4fWdffJb14Ywnzus+9VPR8
s8Q4Wr3hAXrjKCLo/GB1G6gTJXrBWVZ+giISOtUwwcpeNDvv7nSipQ3lqI5TO9/U
AxgycSkLVdOx5C3Ls3w7XDjAKYRO5X4XnqSanL++vz1KYXeayKIVqtbZjQl6ICyr
fvxSVvMcT54iHTfOy9HXD1bPvyPdrfjn1WrJEhdxDQMiCwXa1VQjLT1+TPmij8HV
Z5vf6mxBHmhPQ9g8fub/5Z0VTt6w5xyEaSVFBHh7zSi32geRqOiAT54Es1zapE5F
aTGEbF11UFcS0nH+Yn3YrqgF9MoPVEe+0CPb1QtDFxWtu01pgaSDhCrQCdjnie14
txHAWqn4SP74i9+CnPoF/bIWlWuIzselqM3v6j/BuDeJrWvGWg6UuPt0OpGzxjPh
Zk12B3WV0gD8juiamdA0q4HioIC7JBiq5olXtnP4lkj4eQmYGbY2ByJcZTkl+Y60
7iLaEIApVg3TXcnvZ1BPJcxWqTFWeWMJ17bqcyIkjyPQqrBrwCZ2S5nIq77GPM5q
15IbU1Zr2L5rnNwC+Lj/Ad1cfO9gQkISmB7gr6GyQnr0TRvlQgLLl9lFBI7Rp0Jk
DNkYNzOF98jNQVLkPP4tFc0WxYYbeK8DYRjKCiLXA91yRFNwPnWAXBkYH3ViO9yP
3HlF/OTXcZTK+4dVnqTLRzOW/KbPDIb1HHP+kNevrqoErbMZW3a8dxJrT6IZ4YXc
inGJ+Cm+YMezsZ08zgCKLVJl3IY2N2StBs0yZ2ppVIPBThsfGZ2Lbyd5XoNx4xml
jZnlTI5XmRhCgPbW/0OzxgzSpmWpVp0uYTMezkdywKkJyhT9yj8tYkgsit7UCajW
YEui1+IIR+rxYONGM+BJagun7zGfiKqAMONWAm73Txhqp8w218dfd2TGnRWtNJGt
ElgBG4loacWI2eiLFKwLv28n+rbJit7i8zdZlzx9cu7yBnFVQagIO0pavP2iUTyj
319E2Jr+V3KrKfJ0nPBqSKRcIa96BXFMwIEsGUDghcZiGS5O982zvbrR7Ec20BdX
JVYKYgm6itAdxDjeMfewNg6ykfVP/SRxE9D68F7Mft8dUeRuZ/gR8qLiyowe0YXx
VFeftk0zKtGeOrXvlWJmdXnikVQ+5CrPuV+2XbZzz0DJ4nQ7wKl8lrU5tZZued/I
vpToHLHHAJJDMvyiTZH1CX6qKxWQNFHhGCJyAhcdLORHiMhREwVBi5Uphmab6H8y
epxs+fBs0rEsooGw/H14OeTU2vMPjUSBgsVvHd4KrngsfwNzxHR4A82i80M1o9Lj
C5JuEA6BAfpRP22W3kYGD1/CQmcZ47cPSC1llFQacHUpm6I5SVzHbAEkCSllGLsa
eUZD0l6hr4OAuBH9yL3xZrKmBWioUG592AB2rf9W8IghmdQLHmCn+krIpfmVmm/Z
WWG99tmOGOHXActjOwd93KqwBZHcID/4fWGP97KOJg1LmBHwURAlO864afKHNrfr
BJ9BxYGTADQKdYJakNNrMteSnAAYcEqIo8nNcEkSNpwkigqKMNVklnFcqzb3OEWH
QRcZQWKVd+3//yZPb7gyCYSwEQkFkdaQ1NjcmDpdWq2kucmPW7c+Pyy1GLc3ua5q
VKJiIP+6/xfEKfiXTJ64uBY/zcIMzTLfw3YJFHuBJGDRxJUaj9thV1grsOdC+MZC
CqBzBIPvonBarb08f51iDJU8fA1N3y2abKc+L57rndG//PPUz7ojDlDJf9UWiifb
GIiLMX4GLnfE8wuEWTG7y/yuw4upFdv24TAfSP1UiA0ENz0eJW1KjKTxAiIuOLna
7szKQ/TILsKjszKFk+OcdtiuJBk9joj5cWkjQ5KMfPKkAK1tREGN/Ch2Z8PY95uS
se9YKocNrFRYm9E6cgRmU9fwZwFykGda/rCHRqq6TCUcfaF1Ec861i/mk9CBxSHE
1su/1gV5KvIfW3/u6LB6cp12HQU2mc0w/K+a9sSgOGqjk+9ePSlymw+0s2C/S45L
5AIpUcb+pZF0Wtm6UEaCfOA7llF0PHgfeUu6T0PwyhkFiaSredy6unuWEWlygIFX
KeL1dxslGNIX8y43q/qkrCOpXfc2dAmuSbW5WRLt3EZ9nFoziCyIL57D0TIieGVo
M90I4U/3jshQvz0kCfdflJA3Ae/q1VChfTjthZKRWRRg1I3i5u2ImBejr0/KrGsv
l1pOFvl/0n1eeVIZ+ymqBUQB37ifANNWZkxYpL8BPNGIgMfzlK7GXTlYwlCSaXix
OM/Px4yVdwDkmROZJnwEl1eCz/IYdGDm6nQP22B6snsupLaiqR/HF/RmlWkKH9jt
JX56jCujDWJgFmo5HcrJNB8z+nQMbpg5Xwj5TNMMhhsz51ipfoQHhw42rxtrGz+W
FD50yx6Lk7adH2XyNh+Lei6YZMk04vW/+G+X2DSbN25ciY3HMypOTT/3W/vJ0IWS
ziglceCDqrsSpyXZT+rnVmUwc0YPzTN8ethQw0Dol3sIr5dpoeOjHpsC6GJ+x6pW
letzlnfCc2q7+yLVFvyxM/xA+6jmV9ukJlgqlACrpzwPEhfEEWb9xEcxEAEkQl+A
Nzsjj13/I39suc1zLU7+SGZgpb1JpDy5z4JMK74IOzRcOoaEq6RtaDeGpo7LkC5C
f8GMA4AJXQEQ6iRplwDVwnId2g33GrMc7uvl9wN9hF0E/Y9c8hflzWNyj430TsOa
c65pRfCP/nVn0HuyP2ToXbRGACoE9NG6emWa59mmbYWW+4vQadUUyVegn2YQ0Mjt
Zc4HWw1dnQy0dKJ8YO0Fu1n0ZIqbT2HhlAum5fysgP+WcXJz49J4fpOlSHSJh5Qh
4uEKCQJMSXK3p2wdcNTZQrQcsZLx7lBPYAMh00MErzBaApSHzU6WnqJPh3yDDPiS
+8xoVEi5/lw2HNZSiPh1Svu/2cfHKlGFp/TEw+crfxS98MrzlcPzzW7Qy+eFnWNl
3iNx1JV8xpM3fYx9fnleNzLg3aU/MMQIloUPRUI0uZLV04YX7fzhBCUNRuA8O1BU
D5wnMGo7jz+UFSdi9xG471YPQZ/RMrnx5wrVYQ0dU2Z1TyafuOmySC7wFFVmsjFI
t4lebJc+0/GfM04yPbgvW2QcLDhpjpZZErD6jS6uVwFXSNbUeDHSUSRjfoD8qdef
QRQdXJwGXAknB9mSdLsErlmZkK0P8pG1aL+N53+DCOBE9w65KXB+qhXsFd90XiWC
hmtgyK51MJdMDZJl8ZG05L+i3t8MST6Lk80O9coJbb5eoAn0FUst+J5vaVbAdECn
F6d/IEmj8YiPMYFSgqZ6M04LH5VuKeCrQwzxBvPiOHeCwCitx63syznTVeqBTNdo
rcndJywzLjCOYJZPlM5qDzrRu1jeaqQX6BbGsESC6gDs6k8zrPIvKOHCu0VO5jhY
95ZuG/+7E1BLPxP6Ryc/VQarsPZdSvAHvmosNzFPASgUFTq0YW/CbJGhba5kwRgc
FPTGJ1+ZKE359D5UmGK5eg67uqaocmW5NJhhkJjF8rJLR84QwXatq/vxJsVCY6Oz
INZZo1lw2dPxxseDatKcn2iv9Fs/o6SJX7BVWEsLxCgRRU9HrqDt++gEN2X0azlJ
Vq4IgLm6Va2B1d0fNwBdDYDAkwpgwEVQvf27s3UYyzNYl2+czKYf0UCgD6gDh+42
2POHMmIwxrWU0sH4U0MmFb86PWR43Xs/QzxNPv4J0qM+bICkKZZJ6/EZQIHFPR80
RZZuVoUept+hU6Aest0vreeppXGzgqZrRjRRHVZip1SjD5Yru6rzTavFqVBSi3aT
oRsFefL1cczX43DPYWZQ7VlBu1xTGE2T9fVN2mw8IShGgw0UN4RjGPEpUWFuyTis
aSoNeFjND3XLSVOpiARcwJUZSZMkWb5mgNdInibqexc=
`protect end_protected