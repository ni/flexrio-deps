`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5040 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
3urUxeojDObSx2NGJ45J625QLt4lNhFslIZ0bh45quC8TamlHCpLZOpZQxVAbon4
GNr9KS6EU0vh2LY+rUMSw19Hv6jH2SIDAId9rROPn7K0gHOUGUXhjOMYtFBZMAe/
ivTobsep0bTxHkOUkbGA94gidfKYr427T4FqNqrMgJpTf3IiAyPo+sJCL0rZzIth
JoxC+X6SnjFEkzUXWkXEPvtujJmM+oD02JWlMZoX4/9J1Wqhna/k7Xv6xCDTw35w
iomfnhi6hm72lnEmbKTJO2NuV7XRY5b0qKnGJgaMzJapkJJ6vs4OzLQQzvSof2mA
Pho+Afx8zOIc9SgDWIbZUh/XTgTCZk4v+Zz0QLMJNrKfPWQTCBknPXUyhDZyg5/I
ijFMi0RoSyfGBwVtOBF+vw4xEFjcqzPnBklzpWyv+1+fhktFjBrlOEVnDRzXR4Do
/sTZCQuWTWivYfCnGLWX2jj4zcWR1/m+owBcdqNd9y5H8np4OR4X2YMOo5R9tMNn
BIWUAAR8AN2lRVLZbDpn9GIeE9wpKa9yFzZI6fJFhqUfqNOtVc3hehkVbd+vgNDo
e1O+UYdeW97Jb1nHSTruq00bPvaeplWGCtL4czOCSkODbJP5ezFByXLYWM/4TYmG
qxkxiQ5LKAZBSXJNIk4EGyG2+CJ5cQqNwic4nMDMLYA5m1jsBALb3VDXqdSMH1jm
r1bW9Nbmj1cOdJi53+09NvHhzEPBeTdzjW6XQeoSZNvu8ulX+BL4LsY1p9kozO1m
C8qO2ktH6yIkZ0AGDtVupEaKLc/+x5nyRX+lEHjSbCHTddEEyGF2rbXqiNfLDZNQ
LfFbhZz4uZqi0W3ZpPC0eKnBjiiRFBfxagIQivI27AFW3t4JYhq9c8GcfitVqrSV
yD69C0iYzC3DGePmlkeJsU6HFoSAZnnkLs+KyQMeuWrlzIpuxoIUl89NqMbugMoS
uyhXQ5QTSU8J4AjtLLkFoM3XO96Hd45e/KmTeEdZxBpTgKMdyiDrUxxDSxL6hSYE
K7zGi2AI40kkelu7MWKgluaIV6nVhnqBqiotwzeaGFxgf0w/5VIR2qeH1c4SCLCd
nrwUT0efVvMD7eGK27c0WMlayBUSD4cQc9tOrxf1QPimy/OIR5uy9BdXoVIzkZlc
qPmjtoLOMwaIT8gPbuL52G17lol1vJXC2Fnkrvjw4I24P25RzfT5D1MU45Mw0oMl
Md1Ttb2zC8XfPd09/OsKLjZXyxWTkur10NUnB2V4FFj1bEU4IjoTfOV74F2ClK/x
fBDjpD9VP7QIr5BTlwSL5B28e7eOQZmB+39VnquG4G9gCqoEebPlPZRpH6ysUbM/
gT6eN9SmlbtDklaxGfJC2w9BE/+oIkS+02RPVmhCqE3UP7gYx68q82U5qiT0sHQg
Yql7O8jBHX9n9LDpmutk2lp+711wEeh0LtxEHx44NjxIvRSOaWnLwNDx8EQSiKf9
BuJTmw1m7L18TPfBZ7jvoH6ANZwSlgZUy+MaMXZUYTRV6Bjb4yTOVF6rZbJrqONB
EalJrOjgPNcRlwWE3Zwg8CnZkMqiMK+aH/cLxPvOTsrqCwYXOR3NKfXiYM9txVBO
9ttHcuvZQazw+gdssI6yK/2HTaDE/XxngXQKnHuKHaCF+GU7HOIHehdR3B9M0G0V
pM/9eNIR/ogL5E5IvlnBopnPN59h7SZG2FEUgBqUlTPacxAzQ3jkuJKaaG3LrO0e
/dGggr0ZAKlXl84EIjFBu7uThKalhH41N4uQXja5taj1fHK1ao7krKbh2dflI/d3
bJFB0jBhUmQPI/rYEf5gFK8T9Ngip/bRG/aloEIGVClrWMv5FN0mHGreHAp1RfTR
adUdNg12cv2jYksxWdpNXmwWt00OtKb8xaJCGkYt9bw6usrV49s+jzdgtP2Cyaex
JZPIb44koY8mDLcp8/V8c+xVVA8EH0SMMVLd/34XJo2i4uczPElPyT7X7xvSda8/
L+LF7dsbuOBPAWNHlBA3mcVQQ9QZ3gAu+ztbMZnFsRrVaE+f69bjzTFgMfzrr811
CB0ryA+S/B3ZQCuxKi+YGbHwbuNEM+2ZEVUJUXdHiX5pfFLKXOyfU5TJXLhcN7w6
q0iM7wRBZSzv7kDmNaw4sh2HXjCDT8949AfWVzoTdfuaDLR1fzcUiZ2wNK3T22J4
IqXzsjo6N4/NphfNE6vHiMutp8UDI0slQ2woD7ew+zrhlVAVfidHs+jgkb3MHW9A
S4XBgrn+IhD7jnSqeDmFQ3bDow3Rmv63tHeMZ8/lXaIt2mzuAcS1Wp7fzBsC+AFL
K5jx611hmJJmSmEjLQmq7msNqVIBiamAkaL7GcDlzyfp4F4co281+ZeZIOFSPD4O
H8S8jLFpVb5e6n+tmpu/5FApY+aKQKR7ejiN1if3RpZ0thIHK4YVbM7Z1jlqZn51
iV+zUrsZnrUYFcixN0pcL+qSCAU40N0Fx/DdXN7STrWf91pDbazBPzPKHgcCszul
1WNQGigHtzGNZsJwXUr3u6ws+vDXqVeQKoQ98AWnziPb6oOmvrTL8+iSvhpwKcZM
2rxYBmOXbrTDX3mCeqb0Pf8uCOxkh57S3gBmJvabhT5Iee/Ih4hgdfBt8yIX3q2N
MuDkOvOtN9WTAh2FG88LizwHWKWW6fvkXkBc+yPTD6WFK44DzqH0a3P3BjNIh4so
SpouyM48Ys8RHa4dp1YhMvahORXzbJWyn5QiYPbDeS58NoaOS2TAZ1W0ik/Z4SO1
y7F4oIuUL0NQ3p+5OmfTDy5CWzLevsSGUD1iAth7xd08H8L+DpJqX667X40IYo+e
DXyOpAdL0jHFpPPGbBVZW4YkNyuh+TRe7v0CtwSWUULk9/q6yQyeN6lpYwoSpZF4
9UAyFjdKO+/qfJ16jC7fcqc9sqkTRh3Ef6OR0zbfXYes0oGAP5gjLDbPyfsrodPe
Q1/YjgPS/p2FlPs1vaBDiat0PcDM9f37GvU+6U/Mh5HD2e2AJUQapVc1iF+vH5vR
s4cqIYQQjfi2B60RwxiPfr+N282sNm6fiaTtciC+fXa4rBo7Tawi+/Uk52nvI7Ap
sGgC69BQ9X/xRCdUq2dQn+PabQy4ZPgi+Ocn83Zzunuf1P+luhFu0Jzd2bMat2/s
e+5YZe4lzqLFEWFz3VEQH+TJHcQtE4b9UdGkOE39KuEl3cF3K2FEszDomZsyVuRJ
72MCYbMznqCZtRC+M1FyZhZjlkgnI/bboSuYTuZzfOSccKK91347xtPc/2K3fzkT
46yFFSVEfS5nHkE8OP+5YIiH7dwPWk4DoPP84yhJ2QOa8qVtfF4wuDA6ybVyvKfs
IESwUeNQt0Pfgz4r/dk4c3BaL+KboHNvAsG1UpqsKsfSdhp2m68pX9BMZWqALzNl
CRpO7tkZFTXzyl9G2q4vJvpM0axUj1bAJVxF0JkvQL2ykFPLC0U909rzLk0aQbmd
hozA8H4E5ODQfb0cZcAdor2raXo5Adbsv4ax1klbNeYHOITkSLd09Zvrlv1yxHE5
jp6RVegpCevLqJMnHwy9Fgz/eCT2UJoJGYAVAGRn616C4yQZqsR5CxlG2+IF5oxl
6vLQSgCLVJSEZ2pGoszIBoFW/KFFzDJ+IRrhyiSNJgqGun4VUOExiqOEBRfwvHi+
+pyToOAmyVb/QIIbw5Th7YBXA9qhWkPO/tvvakjqEy4Z27yRG55CqsZ59ZB0xoWT
51SbYr7UtbsubRUTEP4quh8bw2svQhlt1JKJ+0ROhg2pE+PfxkR8OmcgMmOIri99
UEaL7cDQeow0AeMTc1pVfjWdjKDYvvP94uUVdgyglDuuAOxo6o12gGI+pKc9osX3
Wljt2stHINSF48uaCIKtM3TtaFp+hoV48R1JajUGAcgW9DUgRCYT/8B0j0Yhwo1a
0Z8dwwYMMM6dGIzRk8ARZCXsUzVAuGgANdtu6IfbfdqrfcfuxNV6uq6STJHb2KOp
yg9TQRYj/NWDTrVMHs6B6RLU/QM2I8T8vsLKekFqvxX1VBPydy+jyRW/kaIPhrD/
7m5uMy19VN2PUjpRWzdZtw+xnWDd3KGhXopvKHfhMOEc1H43wppbGC0IgLAEbu+E
wX/G3Ll0qmq3UcSGDpM8PpM2V+hDwFRt9ksKJOH4OLcMZ/wGRoSNSFwrusitP4w0
/dqCQN/GrA0WeIPJfttbiBgSV7vIjWOtQw9kdXQJpsSJBULk4bqXs1QGm/p4+ajK
KGQq9xt2v1RtPg4GBan7G95Rm+pK+/DxYNlYzZPZXmKY9ZthFo22UKTCg78Ex0Rj
j7lGAD2Af8yP3J/Y4AEj7ZCpehFc+ESMCqRMHKpdAsc+L6dNm0BtdjXD6txClLsf
Az52Li7WnZ4g3pyrbnj6Pwm/NhaI7HRCG5Cc5IzuC1HF183WDKOWDTU7+mSLSeJn
wJIx/k+ncElnwlEVeg7rg1ds+oY8J7bm+xJvhtZfu8M7C4ylyp+9N7awtNxDktd9
Muu7P562thIZULQcEGBSZuZSiqVNd8IJZML5Id5nD0zAB19sfiCPjeWGmCf7Pb4f
3dY74dKj4oxlJB/3FL47gXVd8Ep6jp3zZMk1Ef8bY9oVH0Rfvn7dCbT+Gkqikj7L
gGH3KZNPOY8kInL0l2fkb/Ef/pF8PstvJP+PDstNGioXw6m1JsTr35cJpBe+Fam5
uoO8O3vG6E+z0tntlGOTRdE04g0DvMU71yausglrJyy6krWijLzPWZO3uUv2CDG8
73XdpiwvUs/t8O51jOAj+5LDfvCl/iug19vOEB1WoOJDLDjmE+vBGv3XvXUMjAtX
cbvaK+3elBNaUeGmMFdPNxAuqUqAZYkSDwOKMyRMCMW/bgAyHiYxRq2sScYsOJsf
GygNkamLrWIiN50aoS0Q29wGMHYdTcSAHDqRGIIpZIdd2k/oKKXQJEI40d4B2kyS
1E6qGQtTy9iqPo3PxnHABrQ67XUFCklXL28+Cyw5sWyB+J0qERL5TEy2RDPgrNHh
bADzKXKJTFUOI2Ishl8vcY7XmIfdzV2DNzr5TrkCOvVHCaLjxkGZDzxiRrMK4IRV
UhQ02hz/Yxny1ONhn3w+az9vk1pT49jjUmNUMBfmI4Pt6vEt7LYUTjpVO0U51N8V
LuExNhByP1vRo3yqS/YBlyl8v2HY8BHgdhEXTa32V4zXN5vgTIIRM5aEcRFMwb/G
vlIfxdrkEpqluZ0orQ0ykXT9fX2NiEkSB8ytXOag4LLVcsaKJGEHRJvV4Jlte9pE
biWhIfrYOPypdrLmLeq3uQxoyx4OTI2obV73/47/WOZPG47McHkiP8N6SRGyLIst
JumGpA/03PQQenokI/15tWNZicUVuMA9sTpLrd6mQJz2ouJuyMu+BOLl/Eztddn+
0DmNt3o44rN+7+80oKyepKJIe50ewoMAc517UjtvmS5pHh0lu0drAb95+4ApzETq
bcPr44hiQO0zaMJCBmylPSK5lOZjqPw+NuyhSiD3lXaAYV2qfE5ywA70Ep6IFo4z
38e3fA2dvLveBZ2qLTfyVCbztZIUx3hUkLoKdLd+egG37U6TQx8DeSLV1lF/ryZ0
DBr58a5dRBRP7hZfjY+MEPP6jTEXjoMQHLFKh7pandt+OEFgA7secgYGpPe8M0RF
oEkr3MiEG9Zmaw0M8ZpBBRnZqp0K7NEC3j1Q13OdrP842AMfpihDb2x8j6jFejFk
Gi9+Eyskrvmq+qhJF2vNLPtoXk9zeVwPkKRlPpTTQdkPiNSq07ZWkvV3B86jN6wP
M0GfCeZbuXnJbJq4yvoHX2g4SZcd4Yzn5852xdnv0fGpZimvKiSsxdpuwNKWIOTc
p1youNoiD7faj9zwgBnNsKzsPGoHbERxXgD3dw/3Psmh5+tHYJBTD9fdIX8Yq6LQ
rNs8hoc7W/bmoTwpheE0EnsM/d4N+IlfZReq0XsOZz/xQYf/MwPjL2OoD1JNswO8
s1/AjkuRPNW2M1Z1oDR7hXViMLvo64z/V4pyASbhCmRL1X2CazFkHs2g1qVwFoz/
n71LEdZIlxkn3aLXysxzxzA4blFmVlw00vjDC5DeezmKazMqMkRgTDpoTj7NEjh3
9IGKgwBPdSDn4Sfa5b7LO94o8Ky9uQ854vmNpB+Ih8lFIM0zn9ZciNDHCBFbtlty
Z7degBg74Fq6bNoG/ki1pCbv5IGUh4Ti7q6u2+eXdq8iorHoTdYHoV0cRbNhIwQ9
MhBCjkWjd+UvMZ7Lkz9vBKL1kFb5b1fvd8Vk2X6zJNfXTAU663mirEg3QTtNdq/r
dU+0jtGjzohFKovNCCVbpzthfZQ/xvhPZaB+kuY2ts5Dx28D3BmV6EFRjtJZ1Fyl
UwXw4w2BfC93XtLGU0Glu5enlImvSPBAIrgOwbQ7vq8eRRPIql/wIEDv2CaGcBGZ
jo+P8EaQQOF0IUBhEnw3zyUhC4HWhQMmXIIkWrpaEcVYwcT0spUiu2Bt6smYIQe0
RHLwT6c1IboFUdtx7j6Qc1mmKDGofom/5Pa2OtpDKveSrrtFvEhUgw0tMHQXDYDK
+ux3x7sQLAXRIMYk2h7Rpa9UySdma2xib03LluzqlKpVAJEgbvNlOPI+acAadmTm
`protect end_protected