`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
hVdJHWSfELCmA4ds+csnOQAALbB3ps7EiTSHEDd//nts1r+JQrRE4d3bDPRJpiX2
Sl8d+xAK9BIi4i+3ruAzYvB6kuD7r+gs02Jsvd/1kn7JYK4xBxCjtdDFjVHOTEl1
sSh1oNiYUwLuwR1yKfP+xBhqxD2Dv6pCKhH1NdGilpJQ6cvivGkSunAu0tzP76T0
4x1pB179E7uIeRplfHWX03KzEBF+eVtfgXVp2W1BGjfAe43y1pCvNYZOh1+TY62g
EgAFgbo7pAujZxZy/YSiZjUr2mGp7o83qMXyusx8+rQ41D3X6rxfuP0RiId2pOpC
6oq5Dfkx04a1dk4s8w8cVg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="Sm9DkM+kBxuxXCFA+l3fFkxuSWV4xqRc4Nn7Ji3ukao="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
m2emGBqRy4AuduN4dffN8194qYvc9UXRqiQc56IrQYMiIVQPyh59I8SYabcDdspI
7AFHnvKD5YaF6tQfxWm+mlcmMEk2Y//aUjxeiGGs+RkKgbHitJF/K7nqg1dmKvDg
a/GaBCq4Bqh0EehlN4ntP5HxM4qcvSfh5m/Coe3drc4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uG91daMWA1mGkhgP3oZKMYye3UAomMWgG80HuuXg2E0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 29664 )
`protect data_block
c9NqBF2D1wSep1rW7utzHsk2j40aow1MnrccxUTvKej2Q1cyeDDbgAml4eTSXI8z
QYgCADtWi7S8BeChdv4B2VxKcS7CMq/DaQrOy1MKTfQzfAlK0iubmlTkljLy0Rwd
Xim13c6uwpYSg2ONMAUgYeHKHZ37vGnuCkHlsekuFyy9ydIEO0VRbM/oVvO6kZvG
oa/qEu9YBlmV3Zck9OjN5f+3XSlUeL4Hk/FNwGUaTpgi531PJ55JZcFAPEoBxUIm
hmOB0q3zlHihiLnWQ9hGvJXyDZO/RTsUSnzv6FFp9hIbX44tZP0atK304cYs/qPi
9tenm867GMKinP/aecSQL0Ay9i4e2iBDZq4Gjo2yORyYmyUYakpfhKPxjbA3wxOs
RXTIxwo00fVhbZIjezyEn2iMNVbfMl5Mi3xOQpAi0lNJeXxQQIxJWoMVG44CPkWz
4cQMBILRB2QrZdpnctenyt9J9DBPzIHu6wv6rZmKhP3p43eWnIu9Hu5RW7maeq2U
iahiToEoKSg/a4AKUTK/otXbUY5zx92/BSp6R2vusaUuG5kOCZTogJLRfjme0A/m
Ph09Hs0ZjVSMo3Ht6VzayC0GO9j03zAKeXMInSn5xhopQluVs5sRL00xDjEKXpP/
dPSJOz1UQsx09AUBo7nxojto1NxOtmUw060dXUpeWYNi/6z86exFrMbKS3NCfFei
tBVu2oMOaRfJQezr8C7JAnLUN8CGFTL1hlvA8EmAEzM0gtSsoDyqGvwK4lCX8elY
A4Iv3XHRnIaAGOFnpAW/YMUYHbbCkuEylkL9fcYcTEXHeMrAnBZCFZfc8Y6VAbaA
Z/7IAOwNvasG+pB2YYkCnWBQ4I+O4MJ7FlZ581pNgvik8c+DrakZ4TvIhzj+dlUG
BIT9uGMKo/gWbU8Fp7DhHQqTSB6EbCVkrHsMD/ishjVAKDeHLn8g1RUP+TGvEn8A
39luPzK7WJAN3gReF3v/k8Mq4t6DkvafREY9e2ZD3XBFmXlYjRCv3eg7Iike6e5P
RNjev+0XP8fgOExVbEL20R3PbjeOg/wpSUhjY/plXrO2za4/U8LXuhRRTJOP9DPB
zDGS1U1R5L28WDSAB/fXQFQspwU3mbdEhvKFDYLar6uO2OuEQWevjxuTFCgXtn+n
/+XQA8vr/xffBMudpRJyU1rCppuOF5HC5Z0HWeCVGRlkDqNPo3FAFzXVToLspNoE
nyUruFwE2glE2en6Jhu3+jgR2YUd9r6D4/KeTmaBtZJ767boDrDIaZD9aQMjCL7W
ClChGw6Kox0WnPKdH9sHwyCRM5/s1W6zW5N+E2EZ7msSNkVP/3qqL86GGKB1iFZW
rwZQZq1x2KWNOyERGLN+0MYA1+QyG7x6WigBL0Pug877ZCSnCZtFrI6YNnOiJZap
hruB4crtWMd4pOE55x1NolLI7Ytm2S/cqGnxOJSlY4wWPFJO2hNMrtxSeJk11CBR
j/2mwtieR3eW+zncZUrtsAmOoSWav1STGlnEf7TzRxBsvkqEfo0KDRYrpmIJzPkf
xwwLdrzth755C2QgaUtfVxUoRVqxQp8fBhXrkwraayUXFef0H+kVOvaYAQyk9uwK
7IOVZeqOyj95n020DLkmEF4eSCY+e4r2Pc27dhMuiYDCtXOb3sd03qT2GNrCuXw5
LRiITfUe4vTbPVc2KQ4Ab9NtQQnJwWQuQVfh6twHhShT6UX7kqbXYTWOuHi8BtxK
HohqK8t02R3zsMKSzwp4U720nMqUIGwBYJb4G0ELQ3EBYAZjoAveK5b3j5I7oAIv
KY2HngidZ5lZ0iG3Mf7r2wl/IBOY+XkbhMPrb73Aj7KlVBc6wL5Ltf4GRZXd0FRT
ihcpvmIDHG8yfH2VEvx37YBnLGTUmqAoazM9qjyVe9nnYuOW4fPCcOsmy1aafvD5
kNZnY5CYmEb89kfJQZYUGVQBUdhd3aj9pY6GS/4ik12ZOYgDecr0hlpvCs56PhEk
jku028a2dIKXHgEO8oHYx6buikNGoQR2//VF+7o5rQi0NV/VRPlgoURXbgKOd1UP
ZI+3azbRw+LpL6nXApl0SD/aZERIbI4TR3NMx2KjciIi7oB8Aysmw8tVg2F+re4F
ODj7F1c+6aQPWvhtKuXvBF2VucsWrLJGTU8wvuM2mnQtTu9/Z/w0BLUajNK4CvN/
nels+IxD8x1FTez7wQCVfjHXl/eBzGxlIWZxjaPBzXRheH0Ei04dOiGvvcs7upnZ
I8jeLp+MiPaYtKvcNOS+FCiTIfpJHLm82J4Y1SkFs5Z8sXoxuuedAO13otdrW4g+
Kt19iFHrwfTEsfyijskHQ42h2YosrOilxeANa7qN2c+hRE7h2vOGkwCmBH9LYKAM
bZoN5xQH8gK19WiHphrXnkyeW5prf50YK3CROMPBerpj2PbQx4JLwjy7TNOy3m4K
75MqfVXZVb/s2h5yLz75pmjjtvrqfjpneVt4HIs5JHlE9ssTBFa6dw551sMBMQgJ
u7IXHK/VmVcR0NPhzET4UOckreW1XxkcX5groE6jHMsrde6UQEclPiO8Cz6KIX9Q
Od932u0nZ5BUJ3AQS1nJaKDisJJtoNlbPW+kuwNXTNwQrAu9ZVmDKIC+wjDMAll5
jxhUtM9/INOsoW8ZKdjbGBx0JepAiQLXUDuR2dN1OU5kfZgcQ+gNi30INOq8pgv6
/n4J/MJ1tkmuUVk6Ysp3GwV/fIvTIPl2kcDUcvlcTNonMJq4ejxa8G6f4wKMX1/3
X0OxNv4YMM3iVzZFbZISzUwj/rneoxR71cgCbUzSg6/rBuELE1NU2kld09XBN2VL
h5U0MAJMBL3+IRow7/qb0sJAOnhOv+pFlrTRA9z9Mi81jawVyhx5FEk4mGatVnjc
COxVMdRl6RgLIIFjF51A3TtIhsmnClisQ8tUmovEBqM67ciWWjdURjmrkBeDFQ1h
XHFOE0oeeVb91clPU9c9uhCa+75gFnsBPVDQityx+3TeCED6Wtkmw0UogAxgnl4p
AJ3jF4T0Ullx9hfvWQ5PFZ+DrP6SnzSoryeZnerkQc2L4SXiy5Myupw11eo4qDsi
txQO4dOoy18uXc1aTGcE3Gt3EJkt5k5bEQcm+rtIgzpW7WBO80EAZMtzHdvh52+i
ET0oqmxKNaLLlrUbSKDe+BckrIhNir5k+ufR/8quuFxNVAf/cNk2nA96STeuhr7V
fzS1cU1V1gxKfKiFgPQJ8kg6W2XcziDuAxj+52a+nyKFkeUQB6GIIeGflNpvvNgd
P2blo0jRq5cuXLcPm3Ecd9T/IgpwzmFwSDhcUmrZQIHnH9GATdSvfWHPt7A2kHrc
PsETECq4JRky7Vnwx/suoKhBVT+bs5h0PWQp058QQwayuqZYIYiufds3ZrXEHTus
xruCYfQIEtPRTeIEvXxnHG5FbQcSte1wj3KsSGE0r6PsiSMW0LNNjTvcJkV/IqkL
LV+Fj8hhseXwd/x4stOsTz8qh7E+Wwpm5hlC4dOQ/ZvjccVoXgCNTin8HxKkycF3
k+STaj5uiCdEEdgWJm3prDs4lYQMXCEUlbkJpVB+QiNhjcrxaKw65fMHOpOoDNR1
wmpRkuLMlEswiDQ+eBVvgVPp76AhqdmP0cv2RBNWsLpcqm4+FTuOoHfEJt3lZD+F
q67uzN6cMwmY4kArUzaJt6lh0qRU+oycNHPi/bn6eCm3IKtyr7b0qxZ8bqQP0ZpV
MBH4+Rb5dRxWjfkEIu11lCiKIdih4GT1/gCbrOQhNTocQi5pXDsnYvVzwYU4ibLg
Qs2b5m7bP03+qVbcfdXjSaiP7mzuFE/Nqv62Vk7UN3d0PLiSxFNKYrUEXp2rplE3
b2V/lhOWBrfvgKsYlVNbyn4grrGO1BClVfPHf6Bh9f1wmc+9adUUPfrHNUHRcAkU
czPiSNIA2nP98xULfzIupHWHIdiTobgetZGLpDidt/LYOsM2lNMpppn4oAkZE57L
6PpUjG655KToGbSrkLu5VjuPvCfM7nD4spadn6oHc28o0xMD/mDwrT1Rl9I9e/qa
qhEUBYx6mTAMJcs7eNS5m0FCyotC1p8ZTB/MGCGNF3UGrJhfsHOr33RcIlbEl8T4
6wFghDQO0+I1T8zSF/WEbgYbyElThHiM/HktdTdP7EOgWhlMx7zW7NJ69wpbrwaW
sfyFeWQc9suUh5QiB+vcweC++Vv4iCgmwYXouOC7ZADTRIhpjccaSMjsYKtkOV7k
245j9punOxVknNk5pP/YApcIt3BPU96jhlGmrzxsM0uiaJCzaQbRYZe+EBtWhfgI
wRFKmxkZKbntBRoj6Ua0OSOn/6/gte2SBDcbU+7wxS4r4Emzu0t3ugcFI9oJ7lnr
fpFPX66+0FqIHgGT6xK9gygVVbXjVQt2uQHjE4qOC0ZI7TCYxB07snj7MBqCHhRA
fiw668T6LF8/6hkNhU9mZUoAKL9weHz1F5GiyTSjCC6pPobhGHP9QbArH653o6cr
/KVdzh7gF2Z0xeYBj/XtL+pnzQazwuQ8tZ1v3/njyar7lhXISwCPSlK1ESqEIda9
gVG8VTL2ms0gVStrSDCmIlcCTXgGshEgK97KAGRdHA96ty92tT3/gYFgUGChyQPu
731pjGMhcSX3KNHwmZSafIVyNvjxngipq73cbMFcPuVxUDPOCA5sg+8DRFOi3E3F
yAxQKfmc5FQVCElAKPUjpGLtJ5Y4DUYwRmIZ5bezv0TDQWrzJc5wVP4Rux5m28EB
fzYiW2Y6VItA2O03Qur60cSnLY4aJzrIRlIkEqtVuVdmuUmWfA3UkfQhh6ucI/89
FBk/UK9noC1PkdOwnS72RKx4kSgP94IGZ64KSWger/hYqO/W/6dN/Rynly21iGOG
mM7UyCIgdguCCUHJtF/REaVsnJNv7qudcBCzJlAPOgwiIIPDSAec1jkmm6NBAYCh
c6FpLQsRH4Sz07qOz1hFKdxeQ+cpu4pCakfALj/tx5Ef96ezkgf7WCfk2fW6R7Me
ldkT8BFCCx+69mEjcdTTMctHiV+FY224Ik/zptX3ougN6uRtREFq7WwpzUNQ/OhG
Z7AlPL6N1MiZwa9gMi2G6DlC1DOzVzjeGZDvJ0UBR9zue+kdDTanr6+qOQ3KtBvF
HcuEox3/3tAIRHa5VEJmmI/Xhn6SYromw7yuAGyH0HJzim6cOlC2cT9vXY1v15x6
VAX7GvmMXj1Yf1S3+0HgsP6uL4flSm9SaiOrnv8LMZnPVn/bKb57bYxgejurAJtV
+EewZzqPnSTon70V1hZy1CZmY29PlBKzQ+U34a5jozG2k4JJL2g6Mc4GQgqlNXvt
tk0B2fUhVaxvy2b1j94SUREVyqiAMipuRmqIkZDu4Dm1HBKYm6OQi9cXhbJgHUzF
Bw335UZj0DUxhWOSJ9eUefZk27PDfQP0uvWok1l/z4P1yvcZHD/pKd+t0gJHMRwk
rVAS1lO+nOox5NdOqzyy3Z8gs0DHg3JyzfwUoSWtsmYMPWZpJXuOLPadRU+jEkVY
iYTkKX4xkioNQMFTTuP8PErsTs5TCSWtxqKKmvtnKW0DZaHV0fQsrHOcVT3yxBZ2
SDzYs5oMXGC4pa3cNukSgx/8e6LXSSuKNpAhzDMstoMmVs6piA9C+mdZR6Bc91kP
AC5rV2B49je9PZalOybZ6dxatjF/OiM/WN8zImeqmjTgcs7DdNYdn2pvrm9EuZuL
3letjp23mPBUWmz1FRk0RuT7Cy2qY/YeufqBbhXqWwAob16gPrCAi6kM5dHxS6eC
VKW5XYwLrDEOj/ADeNqpd7FiFyzfsV4fep9r4Mwd20HkIVT0wFgVF889RTS44bXP
13IDC1rkDDwWZQAThDaTsiguIkGuzEPxpwWkRFWEYFi45R3T96+B5sdnlWHKzAVx
deCKdYapRI35781hF35dOFODjvC+vjHNBGu2on8Fr1UqqwHpDoBJ2LRX7zTLggoB
wkcuriDVtLK1rkyDSvTLP0Uq8HcUWe7gqsvhvTdNj6wKEqjrp9uTmn1pEriJ8RXG
tlo+Qh2zUbRis6IW/NlK2Dj0Lr7sEv697GX830GC7ZEL8eDRfUfmLwrb8fYBnBlV
MvZ/gPIzEtB5FAtiXAJA3LjaMlbTJFVIVOE0Odjq2bSwl+yezBwNZmmsPNJlS7Xh
iaDDeIZCC0/zVF3e+b+1G2hG0i2Cph9i3cFyX+aC8u9aQPflxeKRSWrHOdh6ZIl1
eVEh/TsZjGawPh2BwBj9g1t/zTQ/mCf33tWm/lVvBmGIxXgYZev4jDkmaG0jac9p
Wj3WIcMXpB4fGTnBU8u2TQu1H8FtEq+vM695j0Z2PkoyLotR1XN1a/uFxUVXJqtG
csSwlVxQ7nh0oDupWj7BdxXCBbHzeo062Dr+XpujxN76Cecx0ZqYFGCjqWAEXIAn
QqpIQxT5cj2PvIfHwKF3i14XVm3VnQjrRfiYoH4Nt1cWbo/YqqJroa5kjHd/4AyV
4uIX6zjRpM2xWgN5ttLIczVvxMe0AiWEkLyp7CVDh8u+Owo8s/BhicMDw3SYjfh4
KrSuUuczFDfncukqAG9PGWNpG3IPVN3DrMAy4buL0MQxRlFCT0v1hgzDpkjQoN5x
35bTtHuSSccwO58EB2RRJTT5Wbuvv0HaOyGGxcqdiHTSz0RGsmoAFDPG+mlJpuZL
GVXk+8RizF8Bx89UP9UOJgdeHKleF7iVJY5M0XcFdmxS3sLkh1CwJevmRzCHPX8D
V1WAJZZuWdeRTA0Yzy1BD4+veIiWJ4SsnVsF/U+Pmms+v2IXfjDEgfeAAAI5lMCM
OWSXEB2pYLsOsF2dFlZyxnSOX+T3dOoJ5iKxVRbPSyRZAxhIVibDi8xDpJeZd/1t
/GRyoha21mThrotFdvK2gFE45UILpBPZ90lUoOm8vgtrvmMHuUNzwy+XMu0Qm/jD
4tQgre4Dhn+RwyqpqQcqFmlZYBrQKtbtrlS1sFOnyt6T0SF5prvoAkVxnVG5RkPz
o4NcHVwdMbOm8X8wGN8Q4LnTxDWIk9SJKuO8gL5zWo3h37HB66RieVtVjANmS2qO
wVvoaet2QdSL7SMz3GVfZbUeltEMmdhDjDJ8b13kRxjOUq05LOzi1fZER7PO37sX
Nvj8o5NRm9m9xuoED6N6Ol1d5PaP4r4ff3WgP7SpHnSK0bcXp1el1xxX2HgZ0D4E
75/wN1/hfc1znbfyteyVWhryVVZO2MCJT7/u1pQmvSXAoYrdx1/TObzD7UguDFJH
p+lWSa7yhKpviHd7JMDVY5Xf0Bht1FFjqq6/Q4Gi7t+h8dc0vZJXx1mMNNc+7bxS
sGvdfSmUXh3RgQxMcRpDg3e5GRFps2ZeDTf4wt4e71jBnafcuuBOVNgiouhUYqkx
5W5+Qotz0zSmzQfJK1Dbh5KBQ3ESHvAnX6EaLXkslXXA+8WnN4pPU9t3C+mxa5UM
rUyppRxCi0wenD/pnRxYg7ksZg2iR0RAsJOO7oH2rRXbp5tE9cIF+Sj7F5P7kHG2
8Ijz5XDiu/L1DEsp9u6ArE1vHSJF4l1GMKZI7GChYH2r/daAoQxcFFmytOFY5tCW
O8+/N1zK/GAHfsJgCYDjwh0b+TK0yiU7vA6+GvC0RFdZo3tMUINEhUkqe4od6pWW
leS8dK+sfrmLxpPTQ5o4ClcxWjBlMBX7gvcIN2/8yOV0xO2fHnNVwTXb+Iub2ljw
OsOzljRqwOz92S9fltFjPWT95lI1CaOPskUBze1mHNRMZRPQl4JrzkkqPGsh5N5J
SkGJah/jIzSiboPsG0JZVtIVnclqpdnstyQUyczs0w2JwYVgC2camJbJUfKtzFPb
bkSfnco923UHRRD/35OdABs+YH3QJ3yDOKHXbqsDVM3C9iCG6oAzbRTcdAIi3Edj
n812VSeTelUozzwd6+FAY1PYUwT/NGVqQOMmM1jcQky7Pdn+tj+dwciFYrL9sKiy
avq8ShcRUr2TPYjCCIvlQpjGTMEaLP9UVtHlq/TF1r2rMz17OAr1J78KiipzAmHI
hRQ3VeB+3nBw1UC/HcpNNOr28fmiGFBoZGk+EyxCYW8FN8wXUzTCbCFc/nkCX7T7
xVETwBLExwOljuiHPa7BlJtHMsEHGN1dSKt5xyKB1zrXk4sSqiR+MP4ZkaC//y/A
kTNMou63fG/fpKkwgDnn2Dph76bjXTkE0PZXgRTeteQAFv7AwGVkbXpxz7tS7W6V
f8FpuJj5rXdYaUU+hrj3fR9XcOz/FuYQPAfu7HTqLtguoo7IUfbe+EMtRJQlffG6
T7aYmCY/6f+LrJ0GAA36CRDVY3VBrTZ2P/NcZWVDDqq8B0MrIFOZP37M66ez2wX2
oPnUKIgpNWcbD8BK+yoUE1HI5ZO7g0HDEAqqog8OA6EMO5RmsFmrbqGgSL7oadmd
QstV7LFhwS+w8/qSl9zA3wv3uQ91neuYWth/B1/EfJ5NDA32RO61WINZ5PHedqU5
blKDDHLL+ShoMcNtOnIwynyp4Om9r3c0TpMoqxJ3kDXGwL6SW3ly+XWd5wi6saB5
MX6F6smH/5GI8fj6e91W1kF/lpu6OZW/jGmeycsZUj3cKj6bNxJ1tm1mJe0uqp92
01xif1Q11omAXfZv+d3NJ2QuG2N8KhKqwH4Dvdv97yxL4PxroA6Dm11BPpAK5/Yl
FC6g+9hPy/rn5i+9PnqPm/BU6bM/Kh2O3FU0ylxT8LXs7HIUvIlhuXtg/D986lEw
1eNyfaSM05jSnY1O/sl9vvWy+f3fCC/Xt96ZB2InesXZYb/gelm2IKRHWWsgvibQ
umMhZ2O2PXToqaEpFnRFXfIPCVUpbUCcSUpBC1iIz6KV71ATeG3+nt6GHt4dwzKJ
sEb21tQYHLktkX3XMLh8bKin/BKEWsFdBAyDhwAphNR0Os08cRfha5JYLKO1OC/0
N2mop8dbljl7ooaOG0WWidtvJL0+AA0ZUQstA6lHNAg1DD5KAN6L5T4R4MwLB5i6
JURRFTf2QcboecdCXZhnoWReZQaHb4AXsaTBELMf58V5C6u9AgR4IQDGvpMP9X0Z
DujKjdj5B5ZkUtTA9y74XnMD8yz15sJFWMuqAvyLBsVE1nNO5jU8hAb74r/yJoPy
W5RSd7qbyIEh4PRxhqsVRVRdwMZ1wbLC9Vurk6MFDZjm9KmWD6ThUfqnH1q5oAqJ
LF9nhrdmtVplxTbq89y6dS5VGwrBmL9kB+qTZDuex/PMh5m53OB4OB/QGQ4yaCk9
jQYVM2YNw0boQ2WnTalkSObFfN/CtVjI4otZQNHDld1pwa0npcEmX7sSSZcZBETk
aSBhYc7tpyFqkTkrGu2sbaC/5DP2MawNHYZqhNnef9Tm9SFbmmuhU4fNoahBLLsn
+jPs43pMsqQnmAOCHQWwepVobOCpormo7UMxWtjazR6vackIlE68ihOdEEczjutL
/sitveCLm4Ky4nAfpONsHRCD2YRFgX1kO3AWkwkCxbAvds+ez4DciBPQr2OZEoav
F6J9DOfYYNsNvb27JhUEAZV7ygWdnRVkhWNZ4y032o92VT50gdfsoFQ+wxyt6jNv
7BI2+Oy5o858Gj+KCwW5M40Bci3/GDKQwXnDeQbyaDX+eWOyHjR0dFk91UJwko7/
XMsDTCBCJ+jb2clTYH6D0VtMhBsxB4skMgxGWubFuN1hVGPbCf4PFeWWXZyZFuyj
Ye5zHO1zRb6aTIUiVkRe9FwXejN0/zA7EbQ2uiRp+bBNS/emkB/ll6L1/PkBIpHF
xOtCLcRHIhz1d67eKCQ3b1eEqN98qN90hMAI4fUzXWBpRMKW67u8vskt+vQGy7ZK
Fu3iCZjugW89UzE+DryuP0b8DAX5TBOOWQ4UN3YW4JMNeHPDp9soCKV/KFfD7g0/
e4wi6tl7SZW94fwNxzUksJtAAJwEUhzWkvNm3Vu0xfAhLjOmDSq4SxgOqhtv5wAT
ABnGQ+q8FAk2rgoQHtC04MMZdvW203WJKglLQCx4vDk/gU4FV4oIecsaW9rOZMcJ
g1AswgtCXTy6Xi9GGuER3UA8MobjmT1IkGQeZDMlkUcmyKMEjfXdJdnxUHJLv8SL
BHKgpS1OwibLuCBBLvIm2aAiXc6BseY73aJ0zbY+6kngbIl8gfQC4r1FaG4Dvf/c
18k6lXt9loPZS4ycV0HG+mBks7QvxRfNTJZ3FWXoF7k2i8gVFQZm8OsK3LCc4e7H
oFkeaUMZ8o5zRn/W8rAC7hPvtfeDs+kifsFaFOLZ/StasEiyNPjXMqiO8maBkU7J
kudrCpSxT4vHVfURxhrOkej8LqOuLAQUD0T4sWb7MUnVD/h3ait6NBgKdOcaI0Hq
zBxXm60W9yswMd+RwF9ZP7XdcLH/wKx1vuKPINn0KYknWTrbuVmpUcPmTbM61FsC
mJdI0CZ23idN3pt01n9B2feZVCQ3u25qObBJDrb31LKgUctX9+ILAJPxI3E/LdJt
3RjoBqq8OwL//UxQbbWdmlGu+7WUqcyqArcxJLGSlV+I4W29napAjmjUS3KlwUt0
+QKRAcfrXwv9DflLer0dlw1Yc8DL6EQ8tavzvss7wuZfYbdYgHhe2qrANOlwJlTf
eK3hNhghc/VSpbmfRBjhm8UuljLnVTQ1L39NNDp9expnZvz0ySsvxM0I2PwcrmHk
kT2awEg9FtQ4UDBcwsPmU3mD1nmCCpCDMpYt9LjcHuOt8DvFyEeMdiuljr//5kJI
3QTxDF+LVIDMPD1nbVNADAxQpuuqzRVSt/5xpAt2NZL1r8u2EqmfW9Z5fVwU3/ej
CovPF3U2JQzDPoAadkCFqY5fzCZzuyOYs6AZKQXw3YcuDa0OZ3Ta6XNj3czFrUXd
YRoMi8D9g74uyGuSIICjD3mb891KoHwouJqpcOcRpcLVV79B+C+Q6fS+UbuS4abA
duqLsWufC2yAipPX67Rht3WvpuAeQWsCATrLDD2ip553Xnj7HYYwqQKS78ZRg7hf
QDRA8dL3SZ3sP33PZ8WhTp/BJaHrn/bl6K9eUsqEYXbHOSQVAv/oMv3eEnilLYYh
H0g2KEVRzq/EP6jYBoYqvv+qcbKb5+d1sK9onkEsOjR5ywIES093hNn+5G9iPLGM
7UWucJAdheYPJlhi+MoSk/HQiacpJbqtjHPBOnUldZyP2chdy6bPe03fDIZmdIDI
hY0wUjd/ySDsveBct62NOIxErrSYNvZFXpDSay88Q0XNsZkxrffy959MI3CzGTrR
0Y2oSQeAVVPkSP/ZDg/LAQv/MuZnCXiMC/93eswV0RcznwvADpzP8+YTZddJyNRT
pxuxeiCFT8luEgFaQIuQbAZ6/iyEU0YBjVl2XeFhWjur79HNJrazNspSXKazYDmW
UzeF7PR60SRr0BqOtja9NDYdkwKwwzZq6hw3SfJ2PvOt4/xAF8QnmW2b+LJPx885
z4RHTrnHDfCaZJ9u8ueASV9rk637LX/rTwB7R+EiF+CyMc4d11HhaYfEbH6mlj61
X2zqkqoNN6pT5X2PUbhYsLXPkH54Wgi4+YZhx8hCJtENbBefpBDR/va/OfdLXW53
enwZ3adWA4RUNUMhhkz83Lq1lxeg2uUpwlwjMqD3XB43Hqa90oP9vLnsKTAOYmgi
Y+dJRr8Kz3L7J6DXSkIXuvFSNPZfOMdXQdgGst2s72q9nTajEr4pszZ6Rp8wrc5v
G1ivxr3PQd1BLYrAK7JTZBb5bqYBD0Jqulv9RbKLHVUme+6ILSlUuJFAKcNIQGmD
f/f2fONiiBO6Y8XcXUmPjdJthUy3/0MuHBK4Vpj4CRF2NaHCv68BalrLJ7eI8gCE
z1obijAsGfMIz91ijkU+BS07Cp1MFsVc6LOOXCKxwsBbY4iQtg92a8gcQgwUWBUq
hmNLncqa3ihrj1X5VdP8GallCCB9pE616+k7eQIHIM8LIUff4tmO5iOMFno3RQO2
Z7y1RHQBbXrr2IDzu6G5BLjhTGO64kd9E7UeJjdTlCaEkGTIheWy5cBbTl9Wl9al
RJoPt8dFPA+DQHEGvzLytS3PiQDGbsrQZNULb16gCoeP8+ODSDYZ3LO0mcV5h+jN
wmzh1vEkal9dLiwCWIOutTqa4fGHFW52+YEYOLNbYo0/KJtZzcZ3ntFoj1HkjiVS
Pxp9AnPpUiQLrtuwQp5mCPKQhtkpIUs0/JkItNFA1Ss9O2sHNAyvuWeaFVNvVvBS
XlKJdiNKaHtngCGWRObC7TzPBiBJ/1kqTMXNkCQLtOwI1odliphIRiAQmtjpTXJl
qfiKtZY1Q/FOtneJuGUv3kMt/pxyXXlVYWFA9uEm8c0tDa1N9+8Nt0VGOheW5WAr
5ztCRxxNAPeWl2NyqXs0KFuuEuVoAcy+uM1+Awu5uf7o0TmDioo1sw0XGBqP0kLv
i2nLOUxXq/h1sfJy7GPL86z07VmeBXJ2EJywiroZ4Be6upBswGvLOWtsT5AQ+F3l
2GQjD6UDu9d/RYdmEpwFkm1DP+1Xcpwo9CMPCh3lxkkR+1HjjeHC0K++bPzleEiL
4oRlI2aQhu2SIadzhGkTyd0UVpQ5UJoc7eWm8mYWZLieIyopv1C36waw/8UPXknI
kEQHJYrJ6/YBC8+k14RrwYn0ChPNNF0JQKmXkNNRYyWvD/w/VceymMM25MluddXz
NyAgLyKnEiW469ogWLzNBRKGWVrsay4xR/8EWVqvcRhLj2iozcdWlUcooun7zymV
ZHnrrpbgHglgAGgonLebVK+YgdIl4N7bIBMlEVWiQEBoTIRmWQ+gf9POXTRJqRzJ
o6X3UNgBbETjBHdnhu6eYitJ7VfBcbqrEdoQfN2pVMpSAQeR/svOIR6CAtisliaI
40fWLaxPE4IVIzyGPTFQJTmB5w5DIg64iUs6moNigzLs29YdCR+ujIWqhv3mWsFy
1ABPG9PbJqhBDpBhR18xlFpO8L01ojHeWom9LXNbiBN0F6ixxis2qkRuXVVWs9S+
lTHKuu4P0OPFPlUPI91B1uMD1ss+JmlpJzxBp7DY83c0bnO1FRHoXbENXU4wOhaR
fjiY0Lh+g8EPYCaCoUcO7vBtdwtkPX4ZLnC5M2dlJoeJN7x+TCVv1A5hFaoUjzSg
VCbjZLBIlp1I3yUyGCO5+DHIeQ3mJn604Ym3h2ubkrptuI1Rz/ocswvdtNyl7J7B
oEeoPUKTuHpJJvYtPEl2gOSQsUn0bVDWB3/1ov1ly+62AaoQnV1x947wvYb3kCGI
VssCKCWLaKHpHotBR0n/cxJtDkQfZOiPV3jELz1Ntz0gLIOiHdJ4xu7wPrIl7Qkn
ZFiD4wvgW/hfAjgpfBd/SzqD24QCi3M3nm23QoVKRmbLX3gnRqXiNmvCVcR3hS0O
IAsv3DlDVQkDUXO84BgP+G7/IPEjsWv/XYQtrgHJx0UcvERHXkZaaJliHssyoNON
F4K4asSHnMR3Ot+15stVL4rVZaVjvOTuew181YWS7vewgUa3SJV0VAoysIpYhTD9
JGoei1chvs+dmIqn8kwMjDL4UAlvPrxLk20+7F3maLKmHuGAXGvgQkcKImfzaNtM
coRQ6VSmfsNDZc7jCBf6Tihs4WVNnO0SzwQvNfgzPw4HH/SHX63IOAqY9UNB5oEC
o6UUOXtnXUuLQgZR4iCpoF2afU2h/me2YxFVeZcevDmHrW7k3LuAIi19g/u5HANz
WvHVycC0vQiPZ56AnHJzet1w+258A1bDriQTGIy7dMZWku0bu9O8+ENHNCtMlQ3B
dVgAUZqMeQ4BN+8pdv6Rbi23JJgxCiYzOgO5GScFUtGQcw33ie8YQdwEce6rQFhp
nN7ihQ67Itbee3UnCkbv1ltglkOtooj6qJH9AGnBYTFN0HmO0wgMTiPzMyOmTT+f
DxnVTBr/K6owC+Vol3d/a8U24T+QA6Vd2oDFdZeALiR0RU1Z9LNuedwWlMVXXUvq
FYYEt3WzjEfbijE2j8IiKWAgy2aBT390yRsigyRXNq99PyI/ZekrPn5xwVfARIKG
ZgxiepKCXZVcZc+uNdP3D97bDDVxjDkBKSXbsw/BDCaulFZaipwDxvDTbRDwATlf
7RJaDbXBIPuMibr6DZf2IRBrN+r2HTG16SrI0B3CBOT5Jrm3WGZIf4ugftA9/3Z6
8x9IUHEpgUA+kqAHc78LSG+mkKZXYPUKm5pyNFBa/W/tZ/ZPcNCWSUege1wlZuxF
ewi0sVqvso4uSrr0c5FOwyY40Cb9LkeuJf+k0g0v3SRzcJ+QC+xv4+927t7lvXDM
ZMjUOe8xaAdP3PP5t0tmvBx5/eM4xE9Nf+1dxqSo7x1aJjS2ecoDTG1EpicD58tk
Madu80o+jCUUax78AfIo0808XAqo3s5fphnsRA46NEsuazIqZHtj4/UbmQur21pJ
LbwQeW10hSD1CU9MrN1uqm1PBMxX0MC/rRoujwaoyin7i4AZDbiFTIDc1zOVj4Du
d5GiVqhDIRiXrQpkmU92wrzr4EWXgCL+BccE5K/u1Q5p5S7eLvwEGCObRRfktHQb
O1HSv5hnLxRHxM5ExqhRpdS6rShFdnC3xLIjdagn/QgWEwskGbmprdtpv368PPnu
oBRJUri5de7pMKyzqOEEqJbyV8D4JDWZ4Id/dbAEJlOiCyvE+djl+o4ft4HZ8AYQ
LkGiN9+IRAM702x+ITShmWmDHl3eb3Fj2rIcwDHoURuVd5H+234WriImrdXQJzxA
C1IVWCO8fh+9CiQ5kUSb0WMPP5wf0K5m97/WXoBYV2Rd3RTYF7J48z2VwhB30GfL
uo390XtW/Bv+4JXkywD0kvpZVgZ5FQu23uOJq7CsBdgL2FTbbBdiaygTpve0KT+b
TFhxwQw9vWDjyKa4Ibrh09DDhokD9cnuzfanWuCAk+z5cmFssS+UXgxlzGOMYUJm
oP0syUlqWgHFBBtWNurVlqcIf1rtbbp/LEGoKR7Mq2unsVjMgPN2nQUeW7fDnIeS
17eFYkz/OX8v5Iz+F4SQ30EVsbDga+lCGvNxSikJWTr4OKSxdQqQ8fTf/xwjoFVD
HhQ4warIkGM6jenexibBvXvLy16qJe2n5E4ApAYsg81Ocs4dOiLLRwO2Oghmwu90
jpZOvx7lm6AagTy6JYLySyAiKC3qI13ZEDOTRR9zVbc5DI7rbcT7yX8lq6bT2/Ik
VhMM4gNtKsxPrBVLWp4BU608tSffcRrdD6qbQ9zhMUoa3Y8nCOUeKuLCPf/AcoJ1
9Kz/KOliJy8EQyK7Dn7XKAs+sU+Q2WSRxpQqRBAsWN3eCJA0FLAVFW0qUlMElqHU
ciqj8t5dWtCkSbPWrreJIOBRwVDZ8pJQd4rKyvoxD8m5ssm4dGboII/UYmZrzYma
AGQXMNkVHpxTL/+LqRjYbjSd6IjgOhX6K42rjVImrnpRty5y2S1+volfAcSwMHM4
q9wd6DKVldnJXuyc1lH8CwOf0C4Yo5pA93s8Y6d6JcOAD0vln65Xa5u3n0O3tP0B
xWwTA3/oI6S9sGfDJoU8C1cEyXnyGsseWuz66ZdystEDrMbDqbC+1zgEO6V/RK3x
dq5KNS2Up+70/sMwITlvg55CEhvpHXD0fA2tQNoYbjxxQlIea4vjIDOyxmQP8EFz
k90GWjOhbxsC3WihndGGV1P4e+yWThWWYdKaId7VT0Wz1x7/8OdZLKqxuI9yoryP
OEgnj89vvbZyUOgxJq+OHao5CB9jVvaBxT82UAXHWY+gurkIquQnGaAASPhBzJjt
8loC1DZCrd9I0k3rBioB1pC0Sq5Ra+4LXghXdlzuxrtBSrAJbd0SwzzA6RDlYRKC
0O+6zMOdnidAC5WUfymnLn9pl1t1l6gvFHfAskaViLNVuEckrayVhrKokga0thfA
fIWZUmc4Wnd7XKUJg5Qfs1X1kBsc6W8ICOI+Uu/nv5OL6I3Wi89Cxlum/+yCjHRx
nrhOLHtZKi4vWM+1XBAC4ZAn5hA6fPPLjjsr/lu8O7fttAGDM/e2/aBB610x/DqO
hftX9euERbJpv4kBTTmRBXGtUcc0cqItwiyLC1HpGLIVRv06ZxUnSVjdiBxBbbEb
kzrHj9rySgOqjhZW4Ikl0qpCYPQBylI8ahqDo3KDLRv+n6kVbz34mHJ3Xvp0ZoAY
cXkyG2xR/KMdP0kXoO4hor4E3SUqMyCZN5vtnmzK2YS4NAL/qsy/2LadKHHWkwMV
ESGLVg1yEdD8TKeM2c0otBY7vFr0sYHsMYcH39D//Mu3mNQOjkeumwN+pJ2t92x0
UkQloYE75iO9EEhQUgFEIW4bOC8QmpPutFBa/KzawRV/AGgB9mOLQiW0F/2npais
bcVZRMob5nqgSmiVAEKsaXq1+KkkKD120dcVi/ohueVJjrcBNZJ/79bwpbi8ycFn
94iQeizWkrG2w2y7ssGc3YaCDlhNI3kB7jE9FDrrmxWLYyq4qBonme1jQtxSa/Wr
xo/+mqRB7g26IZXGeLDOO6oCQDe3Yrrm5BneDTCmHolfHw/gPW5Y8lGoUSkgQwEN
3B1XMky8hYjQfYkqGYEBwykiYonXA5VmhFsZWL4liYyYNBvoL4x6jq9jTtcxOrCq
hD2eaX0NZNFtskZXGXHrET8VlInQzw7T8IRUTM/P3LOa6QHDAyisTIi8IgwhDQpV
Rb0gebJ/O5yK94s819dc6mQ5Jn1qdYrmkscLUTiRrV1Sql4khXH82cvasNzBjYTl
PW3d0Cx4GMW5cAY/3fjUdb8MV/yJqjPxV5pUNoHlw//YAHGXUi1cgAehPuDLzCVp
xyUxvYy67MR9Z9/8v2Yr6TYN3rtpjhxwTf3mwssmn/eLPIKhovbwtYj8r44I9o3n
2znrjjsd1yIjLMMdoCHywcnpgRyUrim1yIVblcTgSprq5fuzf5K7wmuXWmaQwnb/
JFiQyf1XYmTgh69B4bngM3pHOEjG4Z8u+jY7VkQ7KKyqcS/Tv5SSF7epIkj2o4+E
85Znnw0fCevaHwzf++DucHH35cTKD71Yxh05Mqyj4kdpcZp0cGhdfu2CfN8Fx4hs
VuYel5lpgGuLY86Bpn9k9U7obrogZai7UbR+/7TweaZwRffrQDleWy/pcR2yrJH/
MbhMlaJSveYbR2LILmk/PrM2KMQwKXBjLKUrg3dGGWJMw8Hkm857RHQt7bKbEe2N
yHqecwnk+rhgVSmGjSqyD5fpP6O63cFt4khA4vx5ft1qlIEoDHikkFxGgeFunlsy
Wc9LfG2dl0CD2h+6PK94d049Te5nDJMfhh1WyP9jzF7hsTlCLpQYpoKS3oVtJLYE
oYoF/7+lSY3sU0yhCOqsN+ss3/6YQi2/Maj1MUo+JvngTj4IlBwcuc0VNNscQhDv
ZfqUOZFRgxql6qQNu8l28enL6TvRwSjeS/8grsU5za4YVBBivfLN67U9l5ku2PxG
r+1dM8D7jmaGqh6AAfs/A3YJ0khzCMY8rMaMkx2Wvo4Z0Pd8BSMkG7pWnuSpJhQG
vbC2eW4xjo2l07RmwZVq+C8ccAUPxoCgsPpjp0JsyJIjDzKmVL12+ejmjX3S3yTB
JtmbekGKIXjycco8/Z3r890zECep+kigfPdzYybg5MCf45tdzpJMAro18gWVI/7/
6Oqkn170qrUtM4XVZmzvMhZfIhnpX457I4SUpy4WxCXCzIam9COFlr3l3o3U0Bdm
VGfzc8MQVLV3ohu+8JsW5Wi24+tbkhNK12CRyNnx9uKCfQRf5HTpyHXil/ySgz7A
ipKPn8ecbQKjTnFUN0Db2MbKUoOb71NcDW4PxuCTWiBaTGelrxiMTLOz8XCp8Na0
4cmapK9vAwYnZlfZ9wxuCSr7EXwggPBlI+ptf5JEErRwKCdmNCOMkuIBSliyxdEr
bhC2WmdR7V23GJVXbsXcwNcuHMGNUKhjjlHSvVPk46gpBoCkwYC9fz5zDypaUsC0
Hb77gjMX4qhCFu/XrcoJ62OVkyd7vL1zXQbq/fw39gKVAJEHIZs/Mx5o0Zno6p4e
Q/AmYH1xpDxwwyssN5C+Raxx3Ifq2J/3wAxT2bEnp41TJdNeBTh/JWhuHvio2vX6
MfaCBhBF39BwzEyeQaIaXSwOaPBvY8KAVmoa3wM7jx/YzCMRzDp7VN2KX4Lu5HZK
Q68O2M8i7osJk/uoOjOs4s/+tbL2fnnSDK+5QsUAkmK5RA8s99S2tf8wqJHlRLGa
298AH4Cl6vFFseyHNWhDxCIwh/b1FdRl4sZupE+iUcXnyyJk5IJDupjetLSzaM1M
2SBf/9f0DkK7jCOzsY3mjPI/muVV/DD4MaqWB4BTAko3Zaq5ppZj3tvBscOKhmFp
cEyzmsIlQy2Tmir7kahMLjagi6YsQLu/IQUaSj4bqS9uR7VQNmDIAZIHYqVJ5h10
kTOwjfBipYzRiliBOfaI0iPMkXLTuj4jB+frMS8jaAtCe6qhQQbAxnluoZ8BxTzs
GdZRzB3M+aGy7XF8sg7PinHbrT971yw4DnVtEuvKZeXBfT0clFjK4+AQB2u4dYo8
RcKyqvgHbfHEoviOZ0UP7wfarkgEPBsveOoRVbgxJU7+FczY846s4c7XRMGDV2js
iuJQawg+ox9obTNqpBgk9I5E2n5+q0hJrB2Cwe07sthHGc/JiRL7JXf/CkLz4RcA
6C6Iv9PDDSZx42aAncyaibZ92KOAytikaMxsEJcx0abzTG3B340bCFS24J0N5uuU
PfS1s5dYoQ3Y3MOdSW5F3dPVXGTZtKkYCinBLp+nqeFw1kX9ZzNrT7ueVf28ehMi
SvYeX4SA6mqXHos+LjGIwmlSq+sT0+p789tWQ3RGRps6zqCQChmjGkuBTFsubzT2
Y6ueB1RAbFgbcO86P3WZ7ty84RmHhp8FfiXcWZEemtnVFAKWDmxMG+hw3nEbt7jq
qcrBDLBsLop74SO/zu2dqazO+kp1pQBhhCuJ3ibfyMQl8O4m5tkvafICSR3rXXaf
MBOOwJqYL9JZH+6HvkVvJyImxy7Y8gPTY4azsHw1Qs+o5ba/1KnD2c1eru3I9rSs
EQaxMc4L29h7BENuUPgswsw0OJJFTsTOJyFFwEJfGEV4hwo8qIDWEtF2mvpyoCkb
drk0+BejFok+5oX+28cB/CF3H7F4pR4kHP7Nw68KJS+Vlj/iYtCgZA1kZXzQXu5V
5Fq3ZbRcAeqxPQl01bXHo4X3yWTdxdxScu786Hyg2xE/buCWTqBSpKRyJ0a16y9u
9rWj98ncSP/ZNcFLSw5TJJmq6QmdBLP7j1C/J9YploPFltmWjdXxkhIB1RkDSILW
ypz7RJq9PuFSNFSvsfRFOEoqYvEydH3knOtt5tD0YeVYnIYCkd4VeU/p8wkdJMrZ
2RKC3p8xHiocit2TLtlIHuGJHu721hqLUDKrQBSEAJBYbuJmf1jAM2IVUsCYtJQV
PEBRlDHVZT1QZ3Aglf1UwKSlB/MGP6EdIW8kK2Ik9MPmflfG/Hx7qAbafn39YWSG
/Mb2lc0baNt0Ma3MhNK+sqR3pqCdh+/o1SjV6F6HTVVa8DIudPgc/VVqaUbVlFC2
MASCXJlLcZ8t1qDfvAHZUgqj1RMFm+o6RneMikDJH9faXT51GrntLU7IDHDnnS8H
wjxX/uFtYTe9qY+LY8zVGJobKB8r9ag2sfKvzujddjHYvqJzxwwnrrkzg3JdemnB
YZu6SIUtcT9VOG8CFAQH/eheLzV3zlFIcgPDVtlQvS9YgrHpCokU7Gd8OzwK6RI7
OGg2y0vGWIv9idJRh/foel6+eLSEN4N0MCaHjzWsXVtdtWEOPFAF3jgAuz5Qsj2H
L3l3jgfQbY+3apQtxqjaaVEdoPh7/iI6ciIZYw/02eLYsodMMIcQtnwOF/SdqCu6
02KDhuCThCow2K9jZ1Vd5gbgkWyraULpe4G614o6cIBrzHD0YQYG5eLnMuUEm+Bv
85OnZR6rfiN/pO6ndm8k01/9RWOJzJJp510xVH8iYTFOKZ/AMZraNZWNZ4c3R8/u
teTZI7esVr6ZhprFOO7f/MtT5fSq7et4FngFhGAeVONMgkdHiIH5ZPuh0etQ6x+R
GWbqSCZ8Gm6Pl6YBXPWhFxjLYTSv4fBG6rrVPkJLZrYV5Yp8qv53HK+fb9c1UQhE
IXAwUdoNTgmZD418dA49wrkrzkZQR2h994/UwCaI7IQuF4YY6SXXywOCACRBo/TH
aS1FnCuoc8evwchAV70ZnqeeN4pDMw68r8LyTmB/tODrwg8ki0fT0yUezqdye8SD
X7w/j/ghtGb63zGBWXSTswEFFA8TDSWcf5IB0BpRq61lbjOcpzWMbOEVbvHegFnX
PufwwQ13ReWpYtKBnzRMNupNOKGaho5O8qGyIWiIemjqD0YtKWYGp8l2znW1HjtB
3d7gQ8DdJXupW8zUnh7v8Ub9COWKi4dKpd8Laz/WyXSnnZnM36hsvccYrpeyf4Oe
0r/pkWhv2upGH0pNP5wpT1UegO7nMncviHCFSVUt0VhtkWj07aZDKCQDMw13+jzZ
OI4GAo3pdkTEpdOCBL9DSBiIM9gX8FRDSDRA0RkQaic1GSTgjweQAXeMYV29HQnL
eAsQwfGzuoOawaHORZfwTO4anjwqBhtefC+eMbhJkz81DdnBqPcgcmzI83p7hFHC
rXEaIPWk+pnbThnt01nHucZELlVy2EQF4HhjpmKw8V88ZLXjqiKYKOAMh+EfPRvV
1uGypzLNFIxt3KbGEr8ERvSYeIJ+z8YtsL7zNEGDQ3gvtXO+8cW/vsHsGjKQvwLK
CaFm+9j5vxvurdLrgsxfgVR0FUttBoX45dFeSY/tQyY3GlDEToPjZr9rhgkt8iq8
j3oY6n7Hxq5i05hSzPP7Kn9rZUxa0vX88W9NdWn/FHF6P/sXhrMkiPhlg1IWBZFX
NybXdr/vrJrqy1/MoNw6v3yg0MhsOXAr6POnSZnbOefoH78TnN98F4hiGkEwGI8l
h5bCzBYWIREjNZxo+vg8o276zR9uVZFkTfy/v/ZozCQRZVqzmmYU9DxGQEr0axjD
7eVEQ6YepX1DqjOLzMuYLyQZw9eY/BkoPE0hBEX7RCjDDUz47HCtEZJ7668sIR+r
u15cTO1BS7w/ui8cSShFW+jTroxwPiZjnLnLxDSsnFdgDPZpQEZ4mRw2W39/I8fZ
UERi2+8DcCIhI+9gll0wdNnpCfe8Z5PwBP1qkZZ4tWVGyttJ+DTC5x5RZpNOcfTh
0lzv3y3vwDnqBXHKMDzZbSe2cJHO4YaYCDUubuEbCv+8KUmsYEeD4GIZGdproT6s
NTEZORBW4znf2vyjVbbqS65OFIhY8p7/tS1QWoTS13Z3AhWXdWEjJnT7NF/fsoRD
lIQRXiy3kiL2eYY4VK01/5xKJi1pJX2+N1DFcyeTdyDnTP0nGnIukWOuHKZpbdVn
sUknx8tcQx+N1wiBwHHhkfoz59Kftx5gbU0jMQdpl21LLOf7vk/T3Noi8BNXKhbz
r2Rl2h8o3Z1YXAVPUeCNBTshZjarh3l7nqbqMufLfPW2zur0baRPXhGnFV5Lblx4
HDLJ6gXC6NaqVes13Lr61J5BadOooNejFyOShn9oBZ7enM1FEupJSF3ptqrxli+I
S0hogWmeCCQ6ODNZ4j9ZtZeflW8I+6nldp/kcivf1P5gKaw8V0cyk5Iiiz0IFkmH
srXkzWAPHLkx5FnHf/rPm78NFBCQ9SM8/ye7YdafJ+niKOZKG6EwL5Ok8EAXHDBO
/2HQvqwAer5KELaBArVRxqZkiw2rtYDfxX4J5gXxnbgzy2Bck7ceHXuKcxXIqnKR
ZfiFXUaAUcZ4xj5/keVC4wU3Ey+eNhZz/jwn/kq09zDaEyFRydX7htZRBB2v+rIt
FmPcTwoU7Pq6sTESxh59y9hRryN0a7JDaVgN24dj4/NaaaHc6rZThOYEoAbSx3y9
/X/HjHm329m2U9OG/Ye1b5r0gLvjioQ/meGOq7a6OAsMuWpjroaBWJLGcQp0dYWt
85TYyKGVP+J5G4iy2tppV+kR6aWFAh1ejf/Wy9oMDEttz3uIF4zD9dbW56He/qTz
NayjJm5JjHtXaDuCfWdiOBzSYvOrxBrc34pN/mhhDcjMNHtrg5+B8sFURi9ZDV87
AHaGC1ehL0OskA2ZNagWoreCBtFhoCeFRvZ2bX8MQ8VDTmB4osw6Fa8BQPaWetIj
3Vny+PsTM0r2IGM1lckvx3BurpmnPeEeFNIS2LRRfaUmNJk772hVyyQbOakUoiAJ
6flM54Oytn+fTLI8y0M6Wu/Za7wvjywCEUPwqIRoIoY/xJJQCr9k7rUH9CwwtapO
JpeKdYMCiunEG19RmdUp0vH6r0kynxi6E06sbq5rhqsYGN09mnOhbzkLhPyxrLEy
sBN43rVOFchOKF8MfmTQvgKymrXIMXmCg51mUOX/bIkpkkaKzveKyu3Q/uI5q1pA
KUxJw5ME1YQLDCmk4uAJtf+YMq/FwUx8wb1FyLuza2tAeAgt65zJ4gozNQ2XticI
Lq7yUkSWn58/4FboVOCs+eHtTi7qpDg4dNVgjUPqAnkaTFhNetktKteutcr77rHd
X7YJWaRxEQ+xy4eGubWxCN8qxTIVxUq0hn3tIT8ri7MZE+MgCK8Ra4AkAyf88e3o
cx+UN0VTrekq1hBug2CPoDgLTwlhpcfu/l57tX/eMlfDACjVZ+S0hQjO4lhLzzUP
T5ou8A/l81+AyGiS/FQPmi/fPhELkLlVBUFU6aUWkjJii3KyT9+L+CjBCSLetfaL
TQz3YX3AHThJ0Pv8JLvlUXeypVk6WgpIRRFqChe3thW29CB1x3lrlSdsUReRIu2C
jGeQ5H+ufPBugQDjE30kCcyUHDslPfaTuw1f8pdAwfUzG/WN48VZl7kyw9jGKOT6
V+o+iPc0cVA/Lfm4l3fImNSrGauzmCXHKwGT3Dr2UxFH3f8tbMm408hSwOkqFB7x
8khNWSCU+xEe+nTe8JMbBgTTA3UwfC3qnd67eoPKtyNZLUoESactFhuq0ZsEbYV0
3SHENZxqd2R0XxQRd8ixYTtZudIRSrpWXA8n9wCw1JAc98S5EbAREm6oOPl+zqzK
ETehFJ0xJPqaTBDiecQaYBKwQ1t8f2S0ETfmHO2Uj2xwVXWhbw2s+haDZy+ZUwk0
JUaZXNXObBSeNOhMdrytxHj1LCcvoThZsGjF+inPOhG9Zrt9hFZacxPJgGP4Eqwo
oGHPQaW6gUHNTP8uQh4po3JTQQCir7F8QoABJLtnRLVS0RSAiEc/D0mBCbsWK7GM
bkOr5UAjp0AlQ8VygeB9ULFoEnH+JcuYtNGkBGZ+lMBPx2mZy9D+VRrhxvCzyw0i
pMnBB9cIGonMptF2omVO8XFHLKsrd9ZvTCOVf1kqxwq/QisCRywDtm+eaoiRmGtD
csW8xA2Cj7u49nNCuBCnl4ijt/965qSoBMbHnWh/7FIDuyOkFSvORG4lJacLb/ZL
F0DUn5djOWozK6BsL3piW2yjjbUlriMugjT3w4W/Is2P04RnLyt4uIrdameermKf
oN3kODmc9MgRAMN2fZX/2cuO4BHYVwDIYEoia9y620brsBzHnOc8wUoDyOnUN13Q
5Ju0Q6Gten72nb4oSgFzhQCP0Qw+U0GCtEA7Lcr/fBlTHdxxu0QT8wNMeV8Waeh1
tHjCOe54DFbxVzYUgdaNHUv2ynlgkOtmo0h/kNuEwR20vG1ME4nXC41PDb4ZUXbu
u0w5DdcM0HJqVStdkt7l4orhU58fop16CaRUcSns9YWMyZVQpzvUzr2RM47mZxpp
ak8Mp7xN7qFfDkTddgE9ozyJdOjUt6WozvuifGrRf2mSBI5LknnrZhuMsUtLAhBE
ouS8rA+50vyKmx5qfnyEj4K6tP/fFYK2ajzP191MtR1vjzkse9I7A0RZq+nYNbMn
1jj/ZYdxw205JuBxS+R6bfY1aKysbx8YTfyZG1yEb0/3/gDmR7+tqOUb0LxegvJq
djtOUc6ka5a4/J7yQ9UHpN5qaR9rnrrE5RuepneYvcXcDstDZnsDrF4BLYXgaCan
H0LSichEyKUARI2IsdwjVWVS/E5M8cKXh5l1NZyjP92GyjLk3MmcpQ6r5f9/M0Bi
FpH29sdSW18yQ+ITEWzZyaxwBW9I6tVc1toznJMnB0nqioBrUT1zRf0SYAyL8if+
jKN9TTATdLEgLYwkPHbob7+OxZqFvd+PzUn2KF0TkuN1KlP44Pifpi8Xw+IKU8Rx
5qocgE6888YcEGRwuWqdZNz3I0XZBCTGDaq9rYrq3hnT6x2TYP+E3kzYJnzhv1Wl
BoAsKEMl+IfJTk2oc2bxFXExFEMANB11VoXhH7CIifTDExCr5ZriyDotQuMidMXI
TBbw5VRDdhAPwO/u3fvGQTDVbaDwAHQIG9gyPBmsyNyAY+kDNmCbT9bC1dR/SIoT
0jK65pKReJNVl9Or0luqfg4P5H6kxllj6icTqmWDkIHW9XCIBQdhznestnoG4CJW
yzIrxGblFHnb9ddLUjptCidwVoYA4cBzSmZdkyb7dpbclHutpKdFdClSz/iOiUm1
kATCfkdDwXjufxde0xQl0nhd67UzrgCiEbZ04Yyf0jC/WtEwpEkXNe5n7bNdxhzk
waXRayVc4Ayfsli3Q517Qt2pbHjrJLGkKqM+IUkbv7HTUCB0CQU7QWL/SCqD9vui
M7ysdZJD4uYNY5IRqphqlDoXbiGdFy28XHk/kyWp2ZY6k5qamv+2QGMOSEtza/rL
mKQ4hI0VTFh/OkEgUvyQTA4d8yKviwoLKGp9qOD5F9lr9Oito1cuSwVMwzeMEjRa
C9xYTUK/jnLZQFcuoaA5Lh7LapY7rplUrvOeu7VxJe7ufzlXWksVG8WR/8DTXdvD
DWeL5sqowGeOcDtreBrhHie1JFkAKbWxQseJHQa38J1GgvAALDeM6EU6Sbz5id67
I2/dc99MbnTToSe0rLsCyMhHCGOPII2UltJHi6Xf2AsVpCm4kjTPMu+2yiOTqRfc
mgt04sT1x4a1Zb9qOhZdsDzGzQo1sH+35zj2g1ZlkCgsVdyU5w0ldvLd19+AHX0/
jfE2yg2z8dhWLQ2OJW2OH03u0udvgjbQyPSgkOH05GVE9wL8QTILvBgDVbg5SgE1
YLmAYcxSLtQ3+pPa7sbR4DoMemo4/Mnhub5MqV8fE7w9q/0w/Lt6VYpG8ws5g8Lb
IN1FUqvhmide3Ph2Dy51P5/sRbMUfpkk81uknucCG0tOrhSPeG1CDDKAruQ3kx1w
KxtAX+7TJF64ltkX+tvjjzRQTEaICZpU1VMHYNg+7X2NLbJXJUG4al1Retx7IoTk
hIE42nmG8JdL8fMv+KdxtjnMSCifBNMpO3HEe+9kIULLgmGfL2nU5Kksy5bVHwqw
2cEyTBCyCUEI/QfBCZ+gL+l6/8QMl33djh75MMhCeDvnh/GfFYkZZVxIi1mR/Caq
qYHRM+NTtjapZyyJ6RFqp7W7Qv5Zuxu3fY8mjom8T14JSRqJ3n83LGG2N2dJqen1
oT79SRHYdrmMarOpmmJ523Pe6H2l4/BpbTBtQielkvjI0LI2DhA/ucuPzUyUBIF2
zPvT+Trecs8Y07/ljkQVywIDyoDxvofPxb3zZTMPzeWoPH0DCqCDBuDpKD2W9Tkp
Y8rHYgeu/iLaO7t7g7252uWU1POTeChXQdd56z5B/QXuITX3Ps9FEpk5PGBdf1k8
LisafC7c68iiRHmiyyPcSgmghbnKrLyjjPb6AXnGjkTkbFrMsJPBr5euafFpfzvd
j7tksyjrcLkzR5HRvehmQMt9QOCaTQFjye8imYcLZ3x6njqGQjPXGnskt+/HUd7I
Kso7MYVdronNNefCDqcDomV6KYlCA536NG+QCGr7jYWCKVJkB8LK6uaBrp5YhFkM
9pZdOfJInEjfUApbO+vqXI8UFB/zJM1d/vIawL3Yoo0IZfqo/yOqJQWXf3J430VN
XUE/OdPEaMSAob9U2zAPgJtewCMPzFXg97jUvxIO/FEGF4Yo9a3Q1qdy0fy5VwLp
OQ9q+sCG9CCR4E2A8DPiCBbN4CUDYLoL0QEg87OwuClSlC+OACHZlyf2ek46a0aA
mB/CVN0JSGT6/Sedb4E0Y4yM769gzcdkprZXZIDHVXrCMHEO3bAqtlmJ2YD8bDWZ
EM57O0r4cVpO4nXgfFzYp7DnO7ySKWfhrmDhhedlE7DQq/kNQpuUSvF6J4bGqWMO
ipWkSE2DZcGpq/G5Tx3CFsaO/eJUjVNDmLTez2lVErZXquSSv106X9BXzQim4Sjk
dORVZMqYFka+ibgHGGm0iFJBc+VaOdqVTSObJfP0lehDN1YjNvfCQlBh5DJGZFj2
iZnshyvSUeEpOHMSA7/TpIPT1pxkqOumrVneU3mmIJ99qI9vzpRHTNJzSMNkn+/8
h9PE9w2qkjYuUqQDDIw8VOScLmhAJ4ZVYF/9jp+n63/CnuqjXh+VYdp2mfLkeFmT
5rjSxBfgwxSEyFb0crWFy7Uzr0ob+4LkpGj6rcWX8roROK9llzD2rRaHLNzX2e1E
xEQrkopoP/uAcscbB24t8rzHXiZwS47w3WWnDfShmm15UbZWZrcLmvcBBAAQh16j
GRhAjpcUesO8FA4uVo2aB58A5zFtPi8rJEgYpdZOefKDTqR6pEUD1xTG4Ki8nFWH
Yb48ybp87nybkQCPYV/Qi3JIm/4qWIgcOci7LdTTTvTpTGjgiyJXKfpmZNnxTFyX
Ui7WURcGfjatdf9JJiUyW79KB4vuilUzxqoh9CsEiReHtDXnyg0DziOYY03pKWE3
pcpucKv+qjB4cwA0hzrTSvTx9SPPC6ieNTAcQLae9SDUB1dfXyXIxrlRKP51IuMi
IZ0nKHZYv3UJLEHzdaXEk/ZExtwqWtH6LhooHLql5TN2NAK5jUho/n5gCBvDI6e2
Wb0rraKSeaZWMig1D8YjrfORU4jt7zcP9saOjgzyYNVowjSyLMzvpW6UWbuXvksm
SP6fdaUxYgJ9wZzAJZC7XcplF4hPajiZfdkeBhj2q5BfiTawI0m8gPo8SMpq4W2K
zZedXQVa4ebHHp/J8EM1reYr/utd1171j44GrQVF4Xv/Ns4Yw8789O6ZBxAHk1pu
g4Y7oOZM9PF7yI6u+yxPgX+j3K5S2lJWxGVubayuZ3mJWduYFqj5E+uE0J0r6+Ka
hpuKYM/RIbkqUzIPZD8bZRxbTR42+WxCWhGy5RP+6EtsgGLp5NPC2lL7adueQl3o
Vl4MIhJ823VPsKuqfOpReJNCYtfMMTQtlI7V+luHXVjEw3REvZ5TdQMSCAR/wy5G
QpGSN1WH3fZAxeLki1FRascYtXP1wgEoYVK9WR5ja5qZY1rwQ/uwYlzKM8LHXumO
7WFhzaWWlTPRFa0jbrwQuo8wcpOKPN9sEc8LHzkYVoZ40OkrdQ2ZduRxjR+9n5ZZ
Xm5pZe2wEdvORh9EGp+Pxp+rQsDyktVoUPHh4Y7kGcmooiiArTTHUUih7ZlNcFKp
uq4ghQcFZZdTXUSKVv7F4hw42RFcWLprLNAmw99eWMfPlQQ/J5Kp03WgpkvicbWT
ITGX+zjBAwyKLxQHSoZsgePfjS55v6q9tk4bGGR9xF9IkmIGle/msDtD8JmWgLbu
jMJewZA21b40wFn2tQgBS4Pvyoa7Uphg0RC2nCpIMRmsZcA1YZjgdCdikz6h5RKA
6YWHufRm443FoZS6Nunex0MEHAeguuQt9Pb9ykknHPsuwabsoUOhDUVlUDZVGMIf
spQCrRe5gp6Cy95w6adFXiegKm1UW+i+Vl0xSuH5WoQobEpePofudayNqSytFYId
izD1eaA5A5hMC6dZqhuJ4pj1qyV+8CQM1bUxrcSnTBjKcpaDwfybz/5aVQ/05TGe
0jrCTlJVvWpDArBPGI0WHqRjK7wjTuPO3jvJrroenoP+ZRz1TZkiPIS/4M3sqss+
AEuyitFIptuS1NNMvQxVMXFI+s28PmqxpmljJU6hjY98jlIF8/zXgZvVH0MSnqLP
FN17Qv6IPFcHDYFyvSltedePe9q1YQBtDW9MUZ7YLiWpkgVISZAhebO4pni7pUJr
+rVcoj9dENw07kB9h8EzE1yT5xiXWvpWUh3+qXCt/uO/hK5zwuGTCfQz3rjyxEGX
dY8MAk7QdujX/z+Gw8zA6r866iWW/YOCx4HP6ZrEtx8mnYaATcV/oeShgn/BVm2J
xf4zvSY4r1gxp91f/HXd+IEh29Pf3BEOUaboEg3faz+256dlAJAwivoXnJRoiMH0
EjnnD1lxGo00imimDVd3kHDluJQATpXg2HVbxt9/6+BdqqoFTe6Sz9UWsVJv6jM2
RibmyN2ae4yUZXh+pmXarDN2yToP+D1ERaXXbfh7dFd0WowjZm66NmGJ/nOWgIh/
aM85LG4VI4/18FXGdMfY9BzLtSSxNrXNBxMg1swJm9bEJIYyBWFeSs/DJO+ci1j8
JNi6ctpCn52bIYxuBQw2Mvr99syUdcwN3dT9NQoXQcvHxVYk9MfTd1ZCg6ODwYnF
ELcmKp7OzQDwrSTt4D1BS430AEnNYVJVz46eGnEKtpsw+VyjZDt2xMIENj3K8Ljt
988Q7CwRJ0dZwtU0P40fE9eWD3XQDMWkE7B8inOHNqY7Bmg5qs3+V1JSQv5ViMy0
42c8CsRl7VZwC/J/bxBfWz4436edaeBzxF+i51RFb8Wkp05vGvafXs5b12+A15F+
YBU6zqMorRs100MPniqF0jMcf2PqeQl0o5F/v+OWO9lK/0iM9WjXJn5mS71zzcGU
BSUZ/bQvlsehkl+y4O6TEx8VYxq8C1bsgD556f2P+3zYB1K0BgeiETCD5pI4Zwj1
yACa8HKBNUaEmgf37ZPP7kWY7mMZy9KxpzEHT2f4rk+sXu/Jf1Gz+K0mmVhjGsWN
aMV+IqJKPvFVzwGUc7dMZj8lMEE6ek1VbIS0MVvkJQrDAgGBcENyO1dhIaWXRuD9
/UUL+sxNSzY6VzW+6V79P959olqiHZUMYzpGNDRKWX4bnu6wjik+FB2BTzhF16Wt
R8E6uhl27T202NsWUoSOpKq1xXgMOTe8dCxLkr5R+bNG+uWhEF2gmktPUma/aU2y
s1PVOpqOmiR6qSEZWA2yfxQKiCqp2FHIa5+q1UxaHe22W9wtu4mlAbq23OQAYQxZ
YnU0oQyK/xOeAF6XtKhPPID/SdthCfuoOP8qzFdrNX/nbvDBhLiSPsQXfna6Ung3
fpJ440YTe2irUxivfbHbCzOhlQ9/tAn5sfOluOJlEwy2FA8fKGiWXSyf/aea3shL
j5W8NJwTFfWE24x/VQA5GeDHUcXR+u8uauLbuHfgXMOoN5lsNrnE9bjAN2QQ9Oqn
kVgS5ai+V0SeuLuSTvsjEae+wBYWiTOrN2iZY8+X/8fW+/9O4g6ClNu1+Ys7VTyv
TMrcpYRlejfSNmTne3kksEgFbamaCEIcZoFNVExGH8ygM6MLUpexs3ajDqLhEe1c
upvX+MDnoQS5EU7dWXYmwlIni4n6wrawokxK55CYkQT6FkGnuASaj8sXU3LSRf6s
C7reBejBMj5PWGs1dYjWxt+LTZhgq4dq6s/0QM04OJx+LDMPJpi4IRHkmWVrXMjl
S8hfBVNqUjWQzgL1VDIs8buq8RQdT50uCBRz7qyk36JqQNaaxKRXkeNnP9MGJFxV
3SdRjizRbCxttb9eskSPkwEKA8ANv2hXSylZXUZ2EcjifrVQf/7MKl9fpq678aP6
VvdDeaA89SUJoPFvIIlMD+m/PY+J+A/FruewJXbLlT6RGrtLnRfEzmocd7hYcJQJ
lZ/QekufrRryX2mP8jKHB81uOu0rpYo6OwnpdNu2pUTioZ5TKZsfUTNq/4jP8nse
iB+UnLzEKY/FA3E8NH+CFYC0Y+7xhwH11QdH1Dp/hrBjYqzcTyviKJ2Tbm17hzsA
Y0PMeD23dp8uxQ5+7pwWmMqa6WWLjOnjz1Vuv4xWFepR9OpO06OMTeF1aXTkp0eb
SbfLl9HmPjHHRy8hr+U1qZIsckAaEQUqLylg13l6tkqtQtagYMf9K/8jwqOANs2l
Qau7F6NO92nJSsopGv8DNMaUa4ucyKxgykzyNuprPNY0/5j+LFgdP5nJcK5MBsVh
fkc4pqtxEGLLQMAxpj/SoTvKpinE9YVL8NxNPdRsD7Yj4kYuu6aezPYXyedH/Z2u
IF8qyXiUMU5ruhVD+drYBuP9LRJO2nxOA5TJXkW0xHQqLZSLN3J6SIrAmZw0ErCT
GlINRXGt0pXl+aNbunxCfCDTGo3zy+AdQFCcXbmD8Qoalv8a7b1bPEDHRyjfdvEC
NMJ7C7TrvLQC9RMvzM6o52RPabad1EC/+RSkVVEJCc4DI7G7YP1ZoLUQMfBn5+3A
+Ud8sCBJrKx1qy4AHD2VEjlBPnoFOA+iEdArXd39ZKYGXpYySrHhRo4QNm9p2FoU
adMSCpUoNxegP/iEUn0rNc7s05LyPUL8k8cIaZWAkl/upVlHX9nYUk0RrOgpGErc
lEKi7LW7/DpBjQ8rxhNLXCIdIqX+/EPBY+56hdRsV5o5L6tzMgm8CuqOWsuvmjh9
UH8A6UhsL+yYlPnqZGu83l+W+mmHdurhUo17Bn6po2ZJjBbIzd9U+XBr2OyUtTSF
fFQHZyA1A+7mqIv7I2l0eApkd01KcbHSOjrDroYCGCM/k8iOM/6kZq1jMjc/5w35
TUQPLc/jxIjzRcrr1JE21tfwliNoQ69qEbmggKCHRcaqX9Oear7A5o+KuPO4LFBz
MGZ4UfYurPLpJOmoD7i4vRNs6cI4yKb8Z+a19Hn/WMQmZ08VGCJzHhe5VPKirGp4
FEoo28NCScTszZVJyYyP1lUsxTZVC/dinoveZPDqilDA/EbtO0F3SbzJNtmHM6NE
xa9fllw4HDnLBjPO3JSQFjxcIePir/is9jWMl1NiTbmDq8qaFUr8cqo9YId1NQq7
2o/Hdk5nmudohJgJJidCHnCMrQn+4q5urz91fk9rgMShsB9IRhddvtPv1zEdV+C4
uvoyuE4XmfUjs7viGZ/wfBfPIiusz/+SB4i4eYcZBa6DxwpVqrJzwi8tB53tBkNv
mMitZ7gCdu3ZDNFs3MEK+UtWZpvAdnkLuZpTweukOmMzJMCY1i1wUDkEqNcJrvIm
bdmd4bqMF3moCya5PKmlQOaIAH6A6pleXZ/w7Qs+hDqkXJq3/gzJT1vJ1ZJyaVw2
9QMo+y5tkWxY6XpNfgKrW0E7rOo3HOMfVFa7bb2oCPMzr8XsqRkmDSuvdAcwZpbH
pZXoGJrXXWZGiyJNfWMl0lKTGCPS9UxWEOAxPiGHS1G+IrjWz8OGEUGRHT3TMqzI
U0mRuiDoOR/MwH9OuK4PeYe4dFk2gs0Qi7u4XxLmnaZ3IYxbyw5IqzLP14OHA7l8
tGuhtYhRNQsVTVSQOSTkiA5FIWD5eY83mfP/e/rCWSOvEAp6w0h9eH8OYgxVtYS+
ShQ3L8KY7NPG8fufjS1mMOoV8GEgxeo8XGZXI9ocEKDbuwL4MGaoaOqwE7djh8Cn
lw95fzVGoa1fPf2L+IYGqc8Um1ONyJ3abClRS8/IKMKAgdjabURXkrAJzr65lyM8
rVHmHfXxkxWpzbfGEOzkv9c8N33J46BnOolYETClTsS1dXS4pQtkmpJXUehoUFxU
KHwWtsBcVFzgZJMKrT1to/yPOkHnPHvVTPiEGluhBSdPVuhtNE81Khj9PP5DZpj2
fNt3nIIxsMzhCVN+seXmTe7Kh5IYIyJGBNwWzKLwY4bjoo8VBlYsCGg4fOOZXiKi
xM0X2xk98YDWmrjrgjnlioc9jRKurY7Gd+jWtGsd7uA2VcBgFOjsCK+4L8IpNk49
t0fx9O/b2mP2jXqB/GZXDq4TGZ6OsQJGn7PTuL2HxaGcD6Q7B8eQsEnjA61+2V5F
PiclqV76S9+yTV8xdgcclrkYWY2k2CJCU2Ad79Ib0AtWdKAHaBywamEPvJv65koK
RFN37yieL55s1oncwRv6u2rC3cBxhx/XnwwQ+BE3Oo25pgYpg/g0m3DbL1JEK2hp
uLWwvCn2hiPz1DgR0OA4NAqPnWbA2WRuMXSX6sOkiEaN1MLgMTCrUcej/+TIPRhN
R/izjS2nWihLh9BnMmpeq8R1GSLbZeH6JUZ3QUb1e48LEoJQJpO73s8rcw9GP67e
WWY2ifjoGOgjSLMMpPbQ39ZaBzYMWk99LnBrltue0OcEKh+Gqh+Qg5qAO1MW+pWJ
EmZUIEuberYwH7YBO9fA90jwQQkt55mBOaKFqrH1Z07fOK6G3ZPkNfZZyGpOTUj1
tRTlaq1kWIY+VqI/B7J1jBwwTmVAPSPT/OWDrEXWnbODcwA3G+ilBSyuMmwIJQtU
OAwAECJ9OgH9P5hqsGh0J+aHJVPDmLPEYWlLcSLakTdgXmbx6SMFGhmgyXUsR58n
tKZVnqj8yyWZO/7T8fhvejCABw+cO+FnlQmLWcEbj85hXOwl/NW7OWWp5jmPc4dk
8AlUyzwHXwIjFii7IjRIRuHB5tl955kz6oQoipY11RzamIbZgbs+F5UkMawo3str
BPG3trzMHHPh4cTFRdS5Hh8EDIuAlSGYDPUJF2AqS4DfLUVpMJSo29U9wA8XiR89
q5ytU5Hy3OYf5UtATAykHsK8S6R9njcJ9hnKSfTwWKtkPa1hIHo3NV47Yq1PomXm
+mqnmVfOdtK0AYRGTIVZ9TPDvJ/mbRKUGw3XjVnt9UE+R7ReLsh7mXWQgfqDiWXq
RNq9fNXuK2AolyQe8ZyvorE+LxmuXRGY6vaYE8oYnN+2eRWoPFe+eNzMLufBbAgb
nBO0BdsURh1MFCrVDCDzXzL1DGzgCAVnPKQWIxMBfrgf7TO6T+GIKdCFv69YZyKh
eHxjKfEBR1Y1n2NmBnxugRxYYo+WZN0WQOd4nkuFKNxjqncPSPJKJTo6PN1gkVpi
/Q9yt0TXaj1i02LsXSqRi4nCUAM4OZjH59u6tJml8g+fhUg3NnNSeWcKbwAqYQYi
+4YDv3S8KZ2/FYBAhu9ggwIQcwr2eq1GhsnTwl/MdpaUW55kmFzou2uS1tZhCk2b
gxt40dpmHWsXCF+8MELEEgeoFbIC0yjedfGNw4yyWqSf0HRV7zZ/kxXPmPhWKu8g
ur/WO/nsZbh0VoZKLLEuQ/qT57EUlVQKIZYhoo9HkrY09WFLczG8Gq5Yq1AnlWow
wJFxCWFQnsZNmgNaRnmpg6dYAmzcZfDpMbr6pZKxjdrOfYLOJq5MxEN5ddo7Lxg0
o2dFfXRegPc1X9wwTUJMOjL/vNF0lk7wM8PtHafp1nIjavmrx+z6k157Mw1d1L5w
SyvwWwwLSIIZX561zSfTUzW1Zt2SacPEANXLQt8rKkwp3915+Z7W0xdcq0WySdR5
173Y5ViuR8WzCtmCg1wNKxoX655ngPuHJXKkHMQYLooy3um7v0IjqWNPEf7NCWaW
7FBIxTU5Dzle2GH7IX/i774LNQk1WCjZJaFJP+PUDRwPaxHBsDwdHfPnu5SHXx0n
Vs0wGHg3ir5EtbAJBuDrgVp4MRHiXnOjZPSAIr8tc+aXpp8cEd3gc7DWudzlc49C
/ZB33sdMrlZQb5jt88/gH7n+aoPJEZhqgBEqx6Uz+90nTpXH6d5bKnQg6eOV6kPU
5MyX/5rO0iBLu3dB2pIJ3QV0Nc7NPCnVQz9+lAzp2Z7u+BRLlbvKEe5eAQVrsNo/
+/uE7uLL1ZaxdNxim3D3sHU/1+VpoYr8iGx3BvhwMepxJyrMPzvu/NYzgoSDxsQt
6vd7rXTFXqHerFTX+B2n26wPl4dUXNoZqpPvyWnE56kx6E3qc3zsIWQEO/H8udEc
1GSduYHb9tamSpR/8tfTJ+sfqKigOaU7KbERrrRDdo6UB1FgFbbpDOGXXoVO9cqj
Uv/QWjySQ06jDTpun9nmXtUYx0iTVI8dDByeFg1dgy23ob60qyB4+9rlr82o+3LE
u7k4KKdTaaMBoKBWJbH9qRYAhlhLcBhF0OnRXqO3uGrUDH/afV3nbLL6em6bEJXB
O+qjxmIdwJzH+MSVZMPHbrBJafuN8KOGls2bwSDpLFsfv4aySkj84UjmcZ+fuuvp
McjDFuzcqKncxpPot7kjGUjynI3A5ygc/a2ALeV6HOUq/HSHiEpHqsyIW4LkniME
bZqItLjEG3/CEDp+ZEh7DyEMJnEx+BX+06hD/BFKvIYzmejarpQGaoRq68Oq4thL
4z3WX4TKRoUM2AoGiH+bGoc6XYmCEkPyDk9idowzx2l8otCMkOmsvjV/6t2KcKoq
LvADAjwm0q4hwu/x8M9zQAWkds1qua2eZrbGwCLg/zQtqQA9+uEpaWtgPhEkxG26
QoMlyS/EXYHudZcePY6dOxubFzRrFhinuoxzzyi0Xzh3GOzyp0pWb3w+SmQo1WfS
UrHYW8Igvd/d+dlZfNkpWarntkCwnUMyQTTJmf1dZYK0Dknr6YsW5UgMmmG04Z9W
2PrPES5+yboK51v3osJCuVVf+pXPoJ01Oc4ekMQvMhZmUXOjvqc509EHNObu6q6d
9oMUsXykvQCe06ybXfGcURob+JURlX2oSO+pSjZKzwNubCHXrCM13ABppb95Fkpj
wwjD1YD4H66jAobva7u3IVQzDxtk0cnCpXpLPmigPbq5gVvSItwjp7f3i6gukmte
skGs5XCfJrOEiOfkU3f7a7fqbYuflF/8OWRqhGpz/wNvo41EnnROAS7qFO6bYUq8
pWr766+O5npv4XIjMVMr2tFS0pmUlY9CMn6OH4vMXdyUq2s1Mv+ENLb9OKUoD7lI
VTnH50rejRn8d0YHf/2eroyES8suHwg9aRhWXYJJqJBSabwgXlO/jHJG3D3q4sTc
5dU7IMWXHFaE+8zSfzhJlbdqJr/DI/c1DyRgKujhNu0XzYvKb5RDp6qfX06VjkiU
NKMQ85M6QHWtRBfBQGrHiXvlQZwrIBLWearsR7VgKaT8F4X1W388l6yYm2t+FKmE
mb0mc6I9XDKHM3Jxu8XZC9UpZ12CNN3Q4TzjMNxN32WzMOPYD7eof696dPQh8fXE
9vR/4SZHl3bP5osd3GOEu33LuFE2UQhD/7WcUOTRIwsoeFW4cPvmdM9WS2/yUehL
SeWvXae+ICM9S5EiMxOk3HpCraaCXoDPIgwndFwhsukdLDoKgUA9Ed9F5S64PFEc
sVHUDRTUJurmtKSNws1K6Omodu0UdjVY+XwxTWREXemJt7/a48dY3RiXIdPoyQUO
vS96G45/0TzD/C959t6R8ZWoV9t2NDegA0lklxhEy1ccaiX0VwfnM1BwGwlQ5Jtp
tEAUNFfYSbZ5IjzL30sGf+BvuC8BZpm1HT9ikFeUZDYwQ9z+Op6wwWpA3ehSmGuW
wmIMDvnjLgVKkhQnF33/rDTnq1SdZvX/J0RIwXOOJc4Xyw89ZYAKCnhgqSEWOuI2
KEL/+1x2lUmK6W/QxrqpfpAVhv7WHM/eq9ADdlfK5A0+Ln03sUzFKJA/ZoMh84uV
8iEilWD7D5f3OGAPYrhb0Phcft2ljXsr9NTuTDbZTnOnCmV87LUYQhXyEVquU0xo
IMLGISnjpm8CQZPRhgREolrW5m6kc64EC3+lkTdMURLI0UA0yBobMX+he5yGkShk
qHQz48Jb7td6+H82CKn7XQllvoV8YKvXRze/H0KHDkvcduemMMwU2wfplweU8Yj1
7PzoWF4/+gt0DjYxMCqrij1P0wySqILpVURfZYwvLrZ1AtERyTKd7Sjmmwv1/78J
77CnZqbxSaxGPgpMDRaPxWuWby2WNZG+1zGvTwGQvxH0OTcG2w/VTi1zY7Z28X/d
MRVZRG5fhtRxKhwmnEljduRa4owNlxl7HxkXXU09cDA8jojthYB/+BaD3pztHpUB
qmh7eRi2Rm2TaI6ULoEBvVUmgePr4oXH4QTeRFk6SIs4mqUyAkKpq07pPuwtTGGO
YFHLR89oVJqW+faYyyuwX2dsgOoiPHt+9KaoZzJ5EU4xFyHPDK49dyF7Gr9Dnk/o
+KuZqjn7pw0oJEXEM5Uw/myPCJwa1oHqq94BRnHngSsUO+2vfmw2Y8Ooo5BgDtI2
7unQtaq0gEMVQJuANXiI5qFVxuVPTzRTmGsvqfIt0XBfJYSr4sdd63Zs6irn5rCx
QrPtWKwHIzcJ6lpTFJ0TCDYjGiVOkAEjQ5uHsq6iKOeoIxEi0yplQrdu4vAJwifN
oOkTYk5l8Z7GgqagHARhq2TYtIBWkcrxPzzv7Tv6uE7qVr6lzO0My1jr0Ztv9Oap
Mh4TEpSCips9v4HDo+qrTMOaznYBkrrvRJCFN07kQOnjJxIzKE9lOVAgs/ZpPJS8
KXhzsOBowWQHP1YrcK3ao1la39lGqcrVgp4AHim1LJUeevTmx6BaXJPW4e7Y1oNY
vFKBfVY81YD5bINZ6aV50uH+sI70ZUdmVbl4kMRx1aKz/eqLhrDJgrC4RrBESnvK
YZ33M68X3g1QxclYF0djPrHt9wyf6Y1YduZtdezLX+6egNPC254bvO5EN+UWB2LR
lD/y63JKR0CQLGFbe61kEl3sJBoTM8cMfhpa4MPk53o3Y3xM5suFz7KGzYtmYJCr
8UyBbseZPcVgtW+9plaIjyRzdsSxidj2MLLaJsLT189SZ4a9fe+ihQqg3NeILzxj
a4cuYQxEPQ2oluUOuZKVZIWGkMSv1V8Nxm2GNDJPJkMu0fIigy3mEnbxNY6WxhzS
K3bBCc/JQPTLFe8eewmo33MfcgvcDq6iIduHFB4QMnvDb0yBLQfKWlEo65umtc2h
YFaCvI/qVfFyPjX+rgAsk9gbMGaXdoV1H3s2T8oYEjuFaykx0zwjWx7lV5wD9D7H
ff5QOha2+LvKSaA8NTAFOUzpDst7+N0FyR1OsgPo3X9D0s4kn2gsD51Do8FOUBb2
rE1Fh0d4uu7HBUH3+P/1oLn4a7LvC78EK2HOt1Ns5kDsgZKhIFY00yXSmWkeBRjx
mwewCXOwnfGgI/0MIU8aUvhwfxXZQW+cQIo2LkK9LTZppCfecJobf2YLNcSN2iZm
5Vr5NwZLxIGoF0Yipa8YbFPpLNwxtQX8lALKLSk9nFc6aO9kmaBjSuxOYuLPm6zJ
FKIqd7bKFyXnq1tyc6DL6QdwBcnGTioTDvwulHsD1zpU3BCpkurZJIKb+ubDh+3w
cwS6LS6an7LP3AbkcZaoByilxh/gDRyzjluRZTymPRcNG0rgpG2butSTi6hwqs1g
DGeAkwOBtA/hKPT9ysvfJv6lcqQPE952JWKVMHPc2XcSQyAeXkvNqREa1r67yctt
FxDrf0cupJHwMw4HXLoDTsdmeW2BOlZVVAvrt0R6/Dreb49kuDPrnJYoBx+O+ScS
LuRZaIcR1cYoY+plGR3iZkv/znLKkbEp4IyCzvwkffhdAax1pQMamglylwQ0La3A
kYfX93v5xBq3Xvv80lVhJsdhzcILBiTOeHIk/XZ8U5lhXbCN9tTCfpPobABV157h
g/BJjtKMtXF3yuFE44hNMMwfqQvstMdB5+3rAR+WEZtER8Hf92vLWyRjdb+ECuvy
EA7IIPwyWlgaDepT/ql5Vyu3jUeKu0oQSbWzbDqrUXsvQ7iby/RciTVXTBAdWB8C
t9TTPmhjWQe3qPPUls45Y0KDj1v9sqtKV70Ia8eI3L6l3tEw6qqGiTqJ6E/8sQD4
v42de1W3JmM7oxxJRE4TdZO9ucHZpY4VCx8jV7RSh0gd3QaA48zBSAC7ej2hjAaw
gSyZw7RPOPTxYVO8S31kKIa3IjQCPLvEhgrKPIKYKtssozPQf0C/Csq3/ErbNRcu
grZHRfvmeA/UembmvsSRsGVvQQg/oj9BYBCG3QzTnBt0C6KDOQbhRVHs+MZWQx4F
AC0YIu5Tv/Etw/8X/hUkaKnohh6lx7nXcXGqdM8pcuwMtSJQ0IV3GTHywoo1Fm0h
PAVSMsQVwohADrtdzUt7vs2olRqxy0An7CilUagbLPOgow1A0ObW0SsnaGf2hpnL
caY88k/4zfAib5gHwMZ0u0DG3/jHpulTosd3RBx93zY+pGWJ2FGQ7NF8kqOjq06r
4JPB2DyOph7Px5omQRIgVr3tCx3YFttIbxnvwsl7QST9RlmMz9woHIPVwJ+M9CaI
iiNSL+ZtCQ0dG1mKIXSANxtrnQAsKMghXTOx7phCLyOoJOqQJLXu5JYFdAeahT+w
oiRJAQtGNiHyjt430JptOtUQ8ulMALNxxCWiND9OaEGfDZ8lrbUjnt5m6drHYP6d
uLMl/LltBBVdu512imJmeZyR+ao0TzdjqOvJ34WLG71AqIgrC9SnSlAEZwTFLd2M
YGHg/61vbqq+J3p/8Oer1e+pezayJ3TI81eh987ppN3GDQehDxkWswfgtPLBByYK
XcOUMZ1m3EXItKgE9XpIHSoHhC/TNObAQxEF8/648DNNnboia0P3RFjDOpS8xIuW
pYx8Crvfq8/iVAkzK8S756CXQ8dduzjgafdcMIqPr45wagMX1gYIrIrGG3YSyek+
Ab3D54VIzJ1Rd90daUANV3454OAg8WfBXsdRvH3+ynHLFJLwx1PU4S+x9C7JfP4I
nOhmyNRMAnGaeML1sQ2fWF+DyZ2P8Gxx2HxMEAG2Mu9+QKqArsLIR6dy7oCNtwOD
SRT88xmGVzNoE067XPiNj65eoGYxuJ83B8qcfoC+qpP7Dwftg9Rb5+xzkJovokVi
mkmpp4AEsfdajAQTETBHsfJv1rQ09V60Bo3cdIwgFiebZQwkactXIt0i4X8Alk/K
dqTtYLwZeOYWNQiSM2WE39ooeqgN6eLxq100ANlSYxBnTe7zhg0wrnQcFub7TFFn
9wEGOCFxcRFUIozfkKv7aWHxC/XX0esHsGYXTUyO7x9asHlday/ix44WPlS4th1M
wUQLYzOwAVS2DcZjsDCcHmQPEbvvdP9YgDQm33DBdasmE+nFC13n69BZwEkmPbb8
uXioUm1riZvoeIqcU5FxTbU2jN/+JVrRaWtN3dTfo29rJ0h6PinIboODchH/348F
3UWps+S4cpQzm/vAA3KHtBIE1uahNVnCVPBiopbxS49/BXuw00RP9T/nCol0ZSvL
3MdOZZQUKt6YqJqrXJjMZAm4d7oeqMzaW+dD/+ixNumBiOhyOr3r678Lb8G/kb+k
OiKxAWe6n4gRWr0imKW5S7xOtBQo5s+93sUb31eh4n1ijiclx5Bz8WFebtiAGKel
2oY+OTk0ZltK0j3ui7Me/f+mMCRJpKQnsn4StMYsY4UIYLv2XvKyw7b7QutQnnCC
HSWCEv8UkXy0bAW59S7IXOOzrnUXEK1YjXNLus7XyUsrHCz1vg7av7bteBJ89UfK
PTqzgzLEJOkrMttIC0UTZUQGXHHJ75ml8y8ujsqf6pKtX3pw9ipXcyjinC8mRMP0
L9jH9Cc7zqGvJJ06C8eg8dyUqsaF4CMvd69gU9v4AE2/wssB7YqWVH3OKk1iy5ou
yU2GtpXzOB8J1q9vUHmHd+UrE49FaallJNVS9l9S4w2bU58OKOQXmfFy+HRcouXn
WVS/XYln42+SZZN9u7ZQxC4nD0AzUgHMceMXt+xdsd1U4CrIqFbUubamL677iLpS
AJmdNWyEer33qQRAdlT95xhQmk6as1T920oJ46i6h+5hH4rxEJwWsg6BGyc+lhN+
`protect end_protected