`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7824 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpHC3/QfnGubCjG83+Xjg7QKYIfnQmKYrhnG76Lxp5rWh
Ydpws9ZyjDbMC+Ryua5L0wNZYejsmKfuD16O7X3HCyGNFdzTpjjeHXYuFh4HdZ1D
FIhtU3mr83sCOmze+xcchgGBufX7DMkFDbXx1rcgPCgPoYEUaz03S9wRbC/Hpj3J
E8ZuQDXYg+JFxBqPYTdL0iBfv4sN+aMKZRUDr3NYNbgjxYEmpa4jnWIGdTvCND6u
0PlM3yiqx8vC/AMGJcZx2nT5W2XdTEbwSuGAKC7xU9NCPIcgofBDLmCn4FrV/JeG
B7zFzrscECZrdQPQ9yoB2uD4pyagnVFE1LihBg3zND9B5lkJyOM5Y027uYxcEtPy
O6z+MzYwgpz+JTW1tHyZNdjQW9HV7ZkGnilKPltQabBtTR5G/3bDzrKl6qQcB+iv
7dJ8CqrCX7Kq3axwh/8UsTR9uYCLHD98duYTw6ocPpB3+YYWhNpCn4yrok/Gwqxk
mlpB/kuggY9ErYc3gwFjJu6AlZHBdnXfU7qOIETSqKeHfaw4f6qCECgVJ61xvYWz
db/f9oOQydl63XpePCoYtSvyZQ7d71tErP753QbAQMt6N7Fs8QVHVG0OwVLvk2xQ
dHt/vDujlieX5QS9+Q3KPZd8fqxrTJOezEc0Hu8ZjEDjC2UnizpmF6CIOnxRK4iR
2NUBUyiS1pt5pnWINQjp0HpsdN9FfVsZqFaDU7D/wiM/C1M3oLcvV9SrxJlnzB6i
ltXxaJFOJ0g59507xOXYmlldvyqO2ufsDYmGssMVq00pp6C+jPUecJvedQR6YDz4
uSSJBnTx5SeQ1WW4y2wK9pY6x+MmSYKPdU3pn364CeuKDckXgNN1Svns+niey2Rd
aHk6rjZy8Yt8MQOwTiLumwOOHv/yBGDCInYmWYEDC5ZQ7scwDPtlVHaZdUhriaIj
pTC+nV5mRQBNf8pnVfeSpdpEwqPv1QYzMzBkzLraQZ3GbZrd1yLuHYWkjHnCX2JN
Tk0YrAa0jqk03Gl05VDMfF4VehZMEvNJgXtbV6++OeoQ18TQR265utAOr1avEjkc
bfCAFq2h21O+a7blJ5yYojX3yhdrUUzcY7ILEF8ZQm7UwwRK6Wp3lxm2qYJLWfjJ
PbPfOYa+vDsTAH6PHYM5N1HRbnnyWcYs4f/LWCmzb02rpQEmV3Mcv4c7dodcbpf8
xry8hmWLA54ieWMQOEHghHjrRLIb4i7ks2NliQ0rjIJPkGGJ40PMUIKipirKesZi
4EBOl7Ortz3wm+nZ/j9TwP7aw54Mw05GjlUOsLC7Nsuswl2EpKcdC0kJGm718vUX
42/7CBWatWm0vfDyuJpfZv9yGz34qBcNPzFj1to8L/FVnhwKh8QgTdz59+M0iDeO
NCbLn9f9s1HxiD8MPom7fnKvea9dlXKACZwtLA6ERJ8bJmOKSbKqJ1qpBOG5Tgb9
Y3NVpDTarIH5hd75tu2BBE101p2Q1C2twMemxf7zff0JHRfpbHQ0yxE99OafAkvj
RgjgFrRKtVPJmA5N47oxic7+8mMb2c/QCvigzQMICx2Ud3MTKB9xCmiJNfQygy4L
LY9jEMFHDW4GAaRz7xjTmXweEQ5QWm/5XNVNWrhss/BQ6/aRcoIuxCnHLCap10Uk
Th8a0xHC8715ucI2G7QXxgDRVnTC+6+6HEitof94KQ0g5dCljaeEADRQnX1/gGC3
Hg7cpGSIh+Oj8SiV/9zzc5s5U8cIIBmmWccPjlsMa1XCdfKEW/XUocec0RH2LiNq
emyECoN1F1LTqX29tlk2AsO7FiHufVk8kctmfBgaFONq5ZrDgQrlJJyfCiW8qQu+
Ql0Tbxsv1PUyp8dVOVrDNYWsYELeJDOBfU3lOajypkqk5J7EiE18yrk3k2Q5Q8ys
vyFqSl/MUrElS43NiwBFFOq+NJLUGvO04uVN8IqN873qx4odnoszwF5vrPf2Nawe
WwUVk/uS7BNCxLlpBownITgOI8RtjHKVCwL+97GOPrYNECeP9+GD6nsG+Qms1HJj
4tpOHEosTyxjaII+StPjTwIo1926e4rRP1xvENM+FPnnmGZy4iCF2wgjAt6yFnBv
S4Uxbn8CG9f2i+UqpfCtNDV9xf2ZxplvbUjqEsTA/Cu9V3JPXyPo0PDJYDWu0EjI
Hcy5uwOCKkWualM3GVJH526NWQSsfpJlIXmc+MFeRu7fUPJ5YcWImbYQOiPBYCD3
RLS1NFVjYcavSXufLvHQarB0Us+veaTTiNs8IcwjxsO0IAPmZ1JXgwUbemVu4kk7
9oN2RFwkSSbIqMBM4lEWfGCRRAxBmNtjs7a4z28m9PZPOQsW+SUV+bafjwehhUPE
fND+1l39dg7upQSVoDHy/pyghQLwjSwBpS5o4XaC6BA0ou8DJ6Ttc15wa27qUiSv
l1Wg4blPSCQSDi6zxJnoczfXx2L1R69f8HL+QWEEooagiSOE6WlKkkkfYTlsH3/7
gQ9hsNridI9DkwpFH5wB97BIp1R3AVwcejY4vqyif7ckb7ZEk08ljZMW/dp/+LaZ
xmJCLCXWr5NqcqWPfj8RDr/xViRRv4d/CcZ6VIE+WD3SjAEHCGcGKuPCCWJaW8LX
XyvUE5A5J213fgvXaY5CotLKZCL5gC9Fh6RXIgYqGemxiGP2CZNIpVt8sVA+TU6T
+BvrlEVdRerKJ56GXWSTUr0ghvVhTYhiULpxzUmXQ/p/vLBIskqzC4FHhiNZf+sB
949FQFj+8fBG1KuW/RHuMix1WJzywH9HuF4SRPBgOIciApUu+fURsqKiFAbuBNzs
OYvOxHPMCIeDI7lcAKJv/zE/UU7/3lmbSVGEJPUiV99S/J1Q4THb3KmKn6RI2osl
7p8vq3vn8nt5HUllBcmwDs7lgocsynHUjwMlPsNPijBUlPrDPLSkwSBi0CAPfRhm
pXZwKCsMeda1M4OzeFZG5JxBfp5R+miujbS++MmE4C2a8pefAS5JFJKwgsuI33EJ
hIjES+Hdk2IVWCTVXbWhq2rGZGKEceSqgiQyXsCwOW1boYIPKPK9UrR12EDG4FG9
Lm7Ls2SbHvWbpAR5s3GczVhXjcgIiDYAkrQYMQi034iO2Z0rJ6YYLvjWRkkHJ+pq
3mbH9e/PJmaZPmz2FVVGSHwm7YP52WXLHN2iQrMm0sYwXXViSF+YIoBPz71ShSfD
HNSrxFOnutasr1bK1jQcMI49Fz8NxiZyL4X6AaaRASsOOo9YOZMQfIxNXySHxDn2
mjDIVdFHB7aHUN9J+2kKAzQOeqsCTlzyT7zFG1L1Nm2dEPC08E3MxVIybE+boyIt
jE5Ek4z+ZeL+JLa4UccMloX8iCQuaN90xEFdQH1yMdJghqzRkwf38G//xerBj3TS
HCZyRbS0+uAg+4K0eZN0m+/S1DTf5Wmo3iCAHtKLstgxiUv/bOYQRBfnb+13iaej
p7Wgl2mS2Uif/x8NR33EoUVB9qi6+WFRx/NGa3AW04MjhYH+gYFWpdIwsb5+iooN
EEbHwq7NL5YJCSLMd4COnec5hgwY8BwPCk5Y9Q5GeLJv5C1r5rYuikf/TW0dgWQe
yn3SgEicwbs6anIkt8fMhqKi3mHbo2VA97hJxcG6JhAjbGuYRQquGZGnwGdhLR//
ZlcA3M/nuWbge6G8gpSvX5amzs1JQoClb3AFKUVFadnBOq8ymzUUz6+ciuY4dTWl
D6XReq05GCWE7DKOJGaANJqb+xVqCTW89FFN4CeSqtxkZUKXVfpCZmrQKLL63OS4
0sW4KJLfk5DMiaLImADjoVerkriM6dBuHc1z0oqsEuFYAsugT8krYYzSdccKK4+B
QlPzxC+LyLS3HF39m9sK+/90v6ngnXDOhQeFmuOnfRfG6gIXQfs0aoURvmNGMXWB
gjxLxR5pp6lTyJoeic+HKHSZ/zxU/fM4WjoMeFssFStrrA5/8aa33fBwsq892zrT
Cb9faBquAsXQG2KRo5LIND8kF02L8xbRo9wCG78Lbxy+8/u5990G5y43kpa5Uk9C
/Ss4U8huCcDRoBZ8cCPAJvhBWBYxrKctc/P72LWk4LU95et2IGBIKVfYllmwgGGA
Nn0SsgJLcommV/CyTSzut+bcxQxhNSHl2FkvgXPcOHzeq8uft12PDgjDxvVeEOgt
LvexJ5OtWEj8od4/RpHrdnNgMEjEr9ST1XetiF9DYBd+zQErYFYKgDL+VtithU3E
v+fbysdSGPPE6Rc5quwRXHK74daC/Yr1smPQhqvfLZ01LZkckQNEsrWrvcWU+5Yz
IzZlnLfg4UWk3aw9jTV/ZaYRNj8NgcBjdots2LWOUudFgdu42EHtydt3kOsc5/pP
XgyHHDcWVudxOdr8TLvrERzB5cu4kolQn1gfv3irSsy57ig09RVy1GdDHqTChfI1
+AWLxLdw8tpGOUVW9JrAUAidtHfz+k351iM5i/sOnNRaGYHntymcpLJ+C89F2VZ1
70SCqmmvEq6b1t4gyk1emiv1u/jEkKjP0qrjPweppUDyeaU0gs8hoUcFPHEfCfEA
iOrETCDKd5amHUwIscuR2MMAk4jJO39/GS2j+OU3zGuuvo8yk/nh/mSv0VBDvDXd
ZIWi7gjyVfrb0+Ac5c88OwspJ7us67yrW6N4lHR+ZJcAE2GW/kGff2VRK6M/w6P/
/K9C4w+PyFPkzNLHm5H5CXNcq+kScoYQWdebUmWfO1LFKErgN/+CFlRlwaT6z3yW
rb2XMy2+8Fm6faCmbclc3l9cIFfrv5CqiXCEjgbKu9Ih7zB/We0ZyyicI6TIOqjn
ktDWBS6VcLWKDpfze/VJLAbe9vrq96wiRj3ddKm2VUxi8WPWjHrMRmbiuJnI2Vl8
0qwumiWS2FuGHvcBRMIIG8i3T9HiQk2da2RNAHQHJhoy9/Ye/8emSStJY7PGaQ9G
jERlcFEuBACjsY+89M56K5rRkNnvGrtdrc7b+UmTH2LBg7XKBHCnJIzrogGpN0gy
blLyqkYTEQf56EUc/5T59Xfh+2iIiM/chmvD+nLPYdrj33kSpDHNkTpGXxBk2zhM
p6iHfn24lKjR3aNtDdphE8v6mi2SGiNYDfkBqoeTPZf1n9XYe8+DeeYkv26EW607
SyaoW+9v8pbnWwcpoXnki94SjqFXYHJDJAHWkcji20qYIiX2weQlUkeBYLrpjfcy
p/31Nh9va+hEG7hAs4cQvc/D4DdhDEzcVIVggZdU4Vq+QzfsqgZ8xFNEAU4cgNz5
eOZx1eTNbjRTJNKA4UeBssGAittdp+bGV2UInwuuLP+Y0VJd6C28ZBIwkalCK5zu
oPBsBGRuxOTNdYFzFHA7msG2aJ06BsEVe6C6Cb/b4m2/x1hbyxZrphtGi08/vktt
9rJ75mBUfmdE2i2glpv/UONbFX2ft0oDW5i052HDFVqCkcBAt86RUO4KYB7RN3J4
8EPW/PFW6bCGg7j+ZXgWefc8symVWGhU7WCBfNQqBj+8iP+u3y0CjvxtX17nWFnp
/gYMo6Fu1sP4YuFG6BCy219vwObq00/IHlICyEG2+gjcq3KoSAfGdToRiA/LDSXS
B4HSJaEZNW67CQqRrjW+gJ8NTYPdimmzV6Qf98JU03+VuOkdO2o8I1lDcjFEPCCR
cTlxA5xaQv7qXF67mIxOaEKMX1pDJWEypPmDS13AIzC+g0+oroCIZKD9ViP+x7yG
ewjzM318GJDvTx78qI/yj64mjMf9mYiJPytqCljA25ctQ8XhYMTA4Z3Ww/tLIau6
v06+hxwBb7zDOvUB4nkHpxnHN2A2+bG6xVPb9h9WUr8DgD0MezZEZO2Ya598mHNk
1diCbdRLQh6OjgEvQrTxyR6BO0JDAAcjPQ79o/3QFD8zFMmyYiAsPH7ONM55kfc4
/IuEil9GpLOSMnUSuYZ7LwQURiBQA0WO187wSgsZzQowph84ZVocMe470c+F18qN
is9we6UvbP/S7MEjijtBvpofHqFS9y7s51kyqMKG7JjgzzAo4MY5G4G0jogEiDte
lA1ulLPBnIo2rDBdhEmIJnIaPHpzVgLh0gPAn3F0DDtjDMT6ADmAzi2Glues0P4/
6AqbAKor2yfK22e+AF5RI3f4oshgGoO/XWAbLjITHgXpFh7nyq9MEuP7rBhD4FnZ
g6iTMgBv2ZEWiO+vjuJFndbwp6v/NNVh7q/rK0pFcOLHNPukBj62kOGAxOSCpVn5
6yTkC8fSSeGINOuVFuASrM1alRx7nbVkvo14TNXn09yQ3SmePGia58lgjApYNyLW
fUgY7QCb6uowFAPGQFI8KZQb9GuBokK+Ef97qkq3T9QImP6r0arxGJ4l1vUxURP1
l05vnXHO94dQ+PZBZofKx+7N5dLdX0p9gBsFw+HHh4CQnLY26Bzgh+kQeMNIXURc
+WjRGWHcX63+L0Bmvwp0lJgB9HcYQn5MIjBNPgnFbLg07q/AxavjCZleofGsfhs1
T84p6Se70wVcjMm45J6WutAR0JsWy1Zf65a3zOMzqQTryy0DTyLjmsAbtORgicz9
nap+L4FV+YJMKigS8yQE+op1dtCg/OqkRy5s9lWTWpnag0NF2OsKl63Txv5weWxu
0B1yZN0bUy+o9IDOo8um1IOpwZ40ykkrvFIgtekk23Bp8dV4VanfunyPQusMzEGf
dKFgwOgY1Em1S3k6HfG+ovYefDhWKyipznXWBZv4ulfOiOuaNOMSOhWMOqsP4tAN
WW2teG9hzixdcU4phGhxsH1f4o4aySfECYRGHhVKY3aQly0fJr/vWX4wyMJ6hGCl
0mQHing9wY4F6o08BhSPqjxM4TJHxM9SFsa0v4fHOmJWoeL3An/ZNN4AFGMRWHk7
HLDL2aXRegF0TzCC3THPXfkrGXwGgIezCWi7fjT/tXN5DOh30LMu/9gJ/AZLHy95
UHLlUAqtqaqTpuz3dgbOHfaX2od7zmiDoZXHL1eFrPuauhJyZhobIXu+eDxJC1Cm
WCs+sXRa34oncaIjhGOUcB8/2rUmmDU/O42jf9W/dMlZz4yrMIOf8ZQCNHpsX1xy
p17zntkfC7gcG99LVLuVgdUij5y40m4gzekWPaPREDzXgJU3+JuC6WaFNjmEyPgw
qe/ZemlE+2HtKccKPCPmlOq7Vo02/l+fACW8In9bcHhFEOM2HBfiJyB2yYvCJz+4
JbBxZR0SAJlOMKmMatGvIUY1gSk/sLgGgE035WyigLpGO1icKq11yx9B+//Oi1mq
SCv0bZCvB42EuhwL5leUuNJSNKWJThoOZf+6uRfv5yEdvpz355dtCo3UzeEBzXcM
vsRwyvwZ42+ees9BCmymQF+ZoRR9XnSCtjb3hHs53qDCMtJhuEcdLeoum74orn71
scJWXsL6H6W9Mhlcv5R0Hxpx6gC9RJg8y69N0JxTnj7nyiUAYFVq+hIjTL0ktCjP
tN+K4ZybJL8ICfuwlGOzdaVezB2lF+L2mBeJ7UxCE68P0NpNbEZQ8zWY2KqsgVYd
6nXnoDpnqFdBdGGoxN8344p9hfAwfUg+TXNfHgtX5OG8yu+uqiIYWZ+at3AR+x3Z
Xxpq8sUVRxDNHkPMXe6etJH1TXoovVAkwZ6oyKZ1chyA++m8pxRbrxMQIpKF/B3D
+9tTMtuQiCYmj0QW3TEotGaRT8QhgMDvs6aF8h96vtukgDC3J57IPvkW7Q7AdoKu
fZhIjMqyo3dlovm9r/UVcDtSWGcBYnl8HsGSgfhy5F+fDWvaZtX60KsuMxkeMX5b
Z2xbWefltoa4kD2JrgODryoRe/66+O6jSmmis7knYub+wcXq6bzawveJcYNv2zSY
AELwPz+wWkl8BvHDX9tPZ7rs2QTunNuJvINeVtBniLdMj9EW+bzkrmPGvYCPSmjl
2G1JJbs709wDXqlVywss4CEPS3t9O6oWhwNQPrc0izMnWlrxgRUsZSxShOD0CEbo
EZx87+9GnoJHwpRROxQaeY5Uaq5t4Gk48IEIjNNfqSxIm6pVqwkWU1hIOxkVL0q+
yl2XeaDOgUZEpNfrdiGa1dMKmwiB1MGVeVFipA1kInxVlr+EsSgvofIbP2fKiGQE
afbCvfif1nvJQjEFQKYYBYJtpCqxJ/RzDmNWuER/2DrWsYNQDt/obCTfi5RbDz4w
KD5iXUCgWyawDQWh7yksY3Ewtrb69SZnE3b77futuNaYipLq7dpkBy3/nGh+AOvg
OXOIPdpgFEi/k+Cecddf3Q7xqqJCLhAxdAVxwoVmUrSguDK04Eb06Qp0yF8ZFUZ8
36lOUdPRNnl7qKLVgCORdxnZARGWQxTP11fJPhNsddKlwt+z1bqny1yojIFbjg8g
21HNWcR90nb8kyhbeqpLb42Iu+SAD1tDDrP60fOhWAMcNaZ97TxcZV0K/F894ZQU
L4fJvqxuPPri+MHWVti4kzf4C/YrxNRyghkA8f0kWAEL+srtGQayoybCcrZJSZLG
dRQSh312nrxfVZPOY5HOZRybrorwO/1oJcgMjKmFacE3MDOI25qKkHw21jXcBBGE
G/ZiE0eGPodV25dYuSt2WNk5/+XxqVAQ3djq3fiLf9dzqYAUGaG7gwRNZKFeMYan
UKN/TB5+JXJ8BXpZZOO+t388hjoFqE/LpVLIPX11tvbgSavg8+t8SuT0G2MVCs0J
bOoxJdMaOMQtDKt3CwCcB9GwVMGBOQ2Kh6S+Qy74qq4AyiWmoGxR05CHcXy7i623
HiJp6HGk/c7mf+NLa77uuPi51e0D26Cugx6SsJ2rpRFGIQ5L+GB9LfhLIruu3PRJ
/gWZm7/0XoD/+9ulYVn34Je9x3SyZxE4GFtb0pJ7OKTDvpy4EvtSmEqBbD3GE9Jt
XAv+0kzNdy8NDnuEh5l+zK3XQpAKZP49MUGPI7AgICtb61U5syo0v276ME/kvyap
RBX1gWyiDwIUK6qm8U1U9v2C46S2VUFTt9/b9EYOgFIevZskD0sQwbk4F8XV0ob5
6EMZjZ0v6aichOZSYLcNIftUL+weL4mHdsxxC/goWhkRxBfajPXFpVVLvx/mT17K
nowqAYWc5dTURVbr9P47b3D6gl9gbOcYHIeJhvVu1ScA1V1pC7OqmQRQ4PdT1jq0
ydcyt37DDbkB2o/Qlu87tkUZTYo2DkPaZrS85yBbzfYIej4h2q3F/YejxFVsYH7X
OG3jXKJXp8eE/5vzgWK/fbIQWkGG4f3geFmK7RVaNt+kZc/grU7q7I/FaYj0q5Wx
dYIzkHz+2jT/PLygN/51QmmnXTYEi54fY+YxaZ5WVFTFadzdhqUTg/PjoO4QWNSy
nloL8HqVioYXAfGE+hJAaV2W/0YYqPJ7V0+C9KjoD+8HL2Ypv2vWzQdo2Ub1FGJr
RB0BEujPwHJCahS3Lbh8aSYh6ZmnPYVM2dfAoRZyx8mQabDfEmkGp+YUPEaJAgXA
HrhvSX30g9JhwsJ63sjgjdmqRF1xwiopGXsnI5d7VdggH8UkO+sl9O+ZEKz6UJrJ
btAeVPMuNwK7xZACfNhyS5ganxJgCSKkWOboV3/aGL40dvsbOfc7p32HjRL1vu4R
YdyqmPIPVVpomWMpyZ2acvwFTvZr/a6AZmIkXjqQCyoKYGVouWZa+yrHgtWeQ4uo
G3JoCKIi1p/4WlwF+Ec1/YKYgUIHRqwx3ewWcfRYX3cZEi+LzNgy/evp65fH7UrA
6KEo1tJd3kO+wDuRJH8IVGWQbGOjqEJLSf9gd6mtC8K7TuNywei85a8srIZxkxIT
RMhm6I7Xa/YMKnyfZBo5AaS1nl8avS5+gbw3gRZMasdorQj2PwKstOC/pG0zUHBS
Vef3+Rt63k7EK/CATnyqsgUrSfnpKHd8yrTCtiptar4uq1IEIoqDOK08+UFwjXiH
OiXBtrzr/kphGyVvMsUuhV8u7lgPweBK6Pxkl1JIpbdZzot49m7C8Fq8l5nhgjic
p6+Uer3u0HOpDhTqOFpgjkZ+ev1ye/lfa/NkNEwtmmEWpquWIun9uBOSjVCwLLoS
ZhW8jzGfZCXhTpKiYmuaLrSAjXzBpIpwxgO3muL6lZBfVAZwc8V8Ylf0jdhc6fgR
ZzAg9SPVSMeJhYNcfXmXfiCkfgWKGwxSE3Lucipm52OCOj07/qGRi+oI5rkJC+eW
u8HZvHAgD4HfSaEoMOiSohJ5Y5H/qdfCxXvaoEbDQqB0/oITAOILtQkSzT2ZpvJe
OL9KClS5R97q5vwJDJyRVPAxucyU/oC6AkUwe5R1OtdVDBXlq1bP0CBpXwLZptGk
iZT9ZHTrvPD757zGK4G0/JC2tItqrmBoR4NDxMqLsiTZKbLMSIEAPAV8LWwVbuEZ
`protect end_protected