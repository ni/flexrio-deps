`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7296 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
ijmWZQe4sPvaU04iZFvn8H+fk4c8D7xRaSSnbgUkoMc7hVhgsnzD4n4T87Na5p9+
PauP3nK9naWZ9d2jlrB0c1TajgtrxVEKWMfMIuK6Ug9fe0Q/lYhuWurYd1D4CUrx
YCaK3AMS0clB7pwtZGfaO1KqlpWFwCAHapcKnsXQOY3ansm0V9bw4w1NeIUZF0E2
BMjp1LBOBTWyt9wv8XwzlawhwEq159x4CdItQswip5SGLe7XqB3Ts1K6jXu/UnrQ
CBCgO3kWrjaBhfz7Ky6+NxHzylwEJhMSJAwQQeixB8HsOrxrgIW1k+5OwzB9mg1t
zfCgjUKpcCv09vC+6Q3cj3Y5FD0fDNO927/Kv///uqWA8xRpxuL+ZCfPN5+R3VpM
h6/jTHoPtJ5QQWu+liZCkfgytwzv3T4psTWF+ncgGB8RARiR2EBsyqfnMWRd9fFZ
UfZtusi0JdrKh4dBBI756m938kSXpqApWneiErDsP4tuIxLwFxUohzHRMlEKTtzS
K8iknH58K6Pjq1Cjs6kPzWbPjtHqjuTxskVIL6loAU1kv60xhhEjGHnRL2bJ/yfb
0N3RWfvjgPDxlOu5SF6Ut0o3uW2ITSi1VQ602nrBSVGF1n4hT/8MQYGUJyzRB/1t
sAw4BD4Vl5KYJB9I7qAj38boTfwtgiCvazw5Fgp+ddzwTmqR1xIKiEUcpE/HoS38
M1RWjgfzQZLUb4yCSacEPTAisXgWVU/Ul1KPzKxy6Di5Dn3VMmbpmpzuJW+PV9w0
l8XvD258QMk77uxJZAnlqn1hTNk+pjU971PbLiPnbWbHbMHO9RubdL9gfRI2P/+9
e8oN8i87ouNn8P3UxINXFYcwEotLOoLaAL3BKLc30v+QNNL7CnehT0o5CsE6PTdP
f0hc8aPEBbHqVKIzNuWEAi5ZUVTLkQgmC9oY3ZxLJBk0RZ6iUJlzVH9QhKzYBuh3
kmyQhOq1hROUAWB3E8l/cVoPSivKCX/ZG/I9Ic6yfByzoGW2uTzdvQCO/21FhctD
7KySsRbuosf5u11H/ibkLGRmkPdgcIsTtQ2YoZ4fRnmuglgM+aTIowYAJooHbWfu
VOYI9zWmxtXxxr5xbr+hJFF8/KZzQ2c7dbuuOEz81KUTKZBdFv9CfSmZERRJj9D4
VqDRIsfUrlpm9uyhXM752pZVAP74JhAT3EBtizYGn+1RHOaXoK3ymyhDhZqAfxXy
NaYYgN5VQ7R+Pgk2gM8eDrlLcTRhk8Pj8opYQEqUuScbuECCkNTEKTsf3f7Srj/w
xPP7xYXRvZeBvu91fKJqeQY2gp1a7rMLWkVfZuXnrev88mDpWyAfzizx0Ol5tlpk
xB+QvIoAU8eLXVyQZQdAvwsG497B50Kwev3CjsgLi4uz7l7eGz64I+Freb+Q6M3w
wlVqQpx8EZStn+BwN2a2tjWg0hH9awqOIKUmBc+JkKRHbhT1+7cAjvu1lYvSue4o
ixulFNsdMhHfhC9Tqy/HFzwlqk4645oMVDrbJ6RTRZHl161GyljyjnzSUtM77IRR
xPuNVMyEMGO10JhGWc9Xhuvgh0ZbstVzju+O0pfWDl47EAHp9njbE8Ef3x02Fl/i
DUKIkMVJ+H7saqzzg5gYItiKz8tnpcBgvEpOmQoFHuTQfQdYdgKfH2HZyTP1EYef
cVgUg8OtsbW+C5Tgd38XUR+4YH4NaYg/jpJ0gJBa1mdb5VwMdI4Da6YyGGEbtwlS
SP5QNJrG6cOGN42pmjdBaaXBrCf8rXEjW0xLPrkNc3L7SRv4iFHy2ZgzhbhT/ANf
Uep0pFxplgOiikavgmYk8EqutoV+Ucojk1TppcjZCrt97JS9DVBtcZzom78Iwvrh
sT7DAKTCI+xbyZQIDEXVTl7ecuhOSVRhdimwKA+JQLA9rvVmBQ6qBnM91e161N/l
D/rFvxlc5eMJEN9FdClKuPzLpWkiVSnUvbI2V5Ej6yyfAHEojMBYmLAvhPaiEGa9
UxX9Ypt8AiIVu6yns1H16zNxfo1GVgXAuc3AQZHs9JnjC7DMSEYCfp0ZJElJVuR3
MT4XVoEFkgdiCGzr3eFfV3JYJDY67NryWkdpe6AkEy+Udj4xtx6U8KebzAOmKBjN
lmk6BoDHbVFNW0z6WCmAeWvfDBM8ZV6rQa2bzeOdTP1trtJjlxo6x5qSnSRZBgZK
MZdFjV7jGp678E6yhXcsskyIVdthD/3ckLhxnnP7KMJ+b0cGc9bg6pUsx1eKQLpf
VEpOC7HHTNTWsN/WvMkhsru0ZKhdzcc/wuuHRZSXKzbLBVsm4PrDLs6Y5lXklCAW
07VDT6MKDABlXOJkoG2ZAhouC9ULoZi3ojxRL8WG0F2ADWN4MpWzvzFp3hq/UncV
CfkkOq+mRWmBmutapPozp/HvK5IsMNEDAIbzH/cwx8Y3OY6ygy9zL5mSXvi/EcJT
1zbc9yEhPE1jk9NBmm71qFJHmL08DWDmJYWnYIflxwDDV9glZU2kHzxKO54lj7E/
iKAx1QgbuGyMi3MQBHemFNBIhCOXM/g1F+ajyHIMKEFu/J84hFRSuFPnmPau+yPV
d3wMrNNLibuo2g4Dbd0wrjYjeZLzBIJFu3xPaYMYZH4TC7Zh6WOZLMta5VGr6Z2S
rB0qMep1A2f+ebH+otsiWkdr37HSiaFPvjuO66BYG+toFcWrksTckQ7nNDiUpCQF
VuktB0tr+GLG7l5FvGfZhJX90Ulzkar30NbF48EDSOT+4Hb+TxZKEdfF0AUZQXsG
3potuBuLKZ3tMGJxtbxBJSMk864cnV4WkKMlkWeY+nJRhzGXr+YEfFSZmPh7FgZ/
el3nSKTRHO+YM8BEKQM+o706V5YG1gylQvYx7QC8QLeugUFB7zIxjMOKZD4NqnBo
i8UGtXarcU4M2sXNFLDFlkZo12Bjg7VpZ8NMtS2oCYGiX55A8bWXGjp1acb4SPaA
m+8i5R//A3ln7JmdSSSGiGMkRpBkACDB7cDRIkU2s96zWtL5u93/I29j3ntnODW0
02JEvRU7fsJwXbp/uHkE80BKwJdzFpiWPiFH92BHGAc5M7TQVLazRtM286BgSPWJ
oF1InERFUj4C5XEEy7x9MYvChctrTCHDlYt/UQhhFJgMyH4C2aN1kGU+l/dEZ/I+
PQPUCW0OBgLpxBGz7Svu+fF2Q4ZSUWhem9qOUUn/325hWdkkqfE9VefWebeKo1VP
YSBhwg3TU7uVDE6tCFsZW3Zgm+0c2Mhum7BnxSIXHJdbWoTQwWgjUwTtBPBAVfjL
u/q+Fy0V0RQXlDdXsEEe5whSafY2St90FRFd/trguRdv1rrvl+Gd2ENRAGepvPy6
exDyfNgSe7kGxAx4V0UUX95x1zhMZyysoy0RLBeKrUuLs6ZBo3pnzZ/wD/6ezbxs
SUSkhPMAtguNVS4BfGrmUbDylIHv6I9htTslpfK9TFS0ABdy/IzL5Yu+Fe7rdvsd
rurhULz8BjfY1IL5mTjAH0dm6tlkbAIA5xbdQavkANj2k9sne+otbSUOaCq7ZbBD
Rpn9cDemXUP9WusI/E3+vNf4JmaoI5uUPazh4bV+EzPdE5wdajDd0WcXr2j4M8sg
svkF36MElnmA/Y/Um9C+65ehx18uvMdmiX84MyZ86jzgA3GSftuvphm4z/lqmeFG
Xb6e7LlOpvxXpjm6sJao3wwOyfqkdn7Sy00REiIWu6xmR85FUCt+rLLIoPn3d7V5
p5o3dAFfhLflj7CvCyCZPslEH0Skqb/FA4w6FbOeVpRYuu7UVOp4c3g9gACg5S13
gnJp6uM4gHzPc0p10Jlf0veGxgVExSlOjK4hqKLVRWe4Ly2irg0L3lzYqEkQGhzG
JbzgRnZHtOqqy4z02bdISxcN9tCNqEy9t+j5j42G8D0fYdzGrJFW1faLx6yA2q2q
fW9r8Z4+twet7b+wcrwmxcaL03jYKICPgDtcnrac6/pepmgo0ZI1x7k4WUc2U+5W
1DSYR0Q9No0/TWB/WyEtGXQFouax+Z4nH74AdFUClol/+ciPW1S5Kyz6TqIQMOIm
AvQTi4fGSEMRgXjr6BFkWr0A7LEvVSnfGbusV82HIL2jLjNXsU1O6/K/qOQZEUpC
g/LR0j21EzxAseuzG7l+y36Ql8V+rS931alIc7AtXwD6lzksZVrsVWI9m+eYzlZs
f3KfX2zp07mtpegtr4FB18gWg8/WDhXK2WAFayUuXWSPRIXzudLKnOm5DUp25H04
eSSKuOy0W5cLqvBCxTFd4gBuOW2MuoHD780pXhD6hXI/ejaNmyi3+XwJ0rjwBABl
dkItP1880XyhDOdJwYFphvRbxHmYvAcR6M5EV/a+KHygv5lGt82KmNcAG+0XfvOs
5SzRHXn2ypnjMKZy37dWCYtVpovDgDPsxgr6Pd4+JUxOPg/xtDV6YqRVhDW2ATwA
8V0PQKgoAlMBP0dGWDJ0JSPrhQAjQD5t7vnrAvom3M+sK7+M6p37hocFBqtV55+J
3JWXC0tKRxqsA5UduaR5J2WMVBTtaG83P4fFom39e/a2MQbxMeeMooZd6xXfTjgN
/rucnpvbECChDOJisr7zaru49wpchtCw5eKAQfpJhhVirj2SYcZ/b2t6ZdUIhI+N
RsfqroiPYtomrYNzG9SE0vL1CLpaQffjsrXgRYn8vo1/X/9lUn3BxoIZSy1p3gjX
G9A/kXHPxzSZI56xCse7bee0YxdWk0CjXoKndVhvbdmkWvqUyEcs3dSgwexb6D74
EuUIfflhwQWWSUQKWtvnLXiXLN2FwkYh873vlOQ1iQ6Bki+pl4oo84qBGBDldTkU
5r+/GC+F/P8c7795oCF8Qa1CVWX1VLwHGHAhonMIZBd7UFC8RauGVeDxGAUafaKD
uD4wTNDsknauhYb9MGswpWXlCQXerVu8igWN/Hypu9dSXX8Jk0UjVT/12JGfu+dD
pmGUmYC/tg0bixYd9K+K4D4IaSk9r4NOube09AMtZH8Y/ci5g0mUztA//EMMnZG/
LdAVG5GJ9fXqKFnV/s3p3k8SU9bkrVaCDdE9tn4PvHQxM/lYmTulNG6yYHrUoj9P
X7bP7zfXxmarxF1yTbo4J+AeJNo/qbD2yvyemtGnALSwBOWm4KeyoJY5jN+PgSZx
/Z390npo7VOgpaemqbqkX5Z0ZS9pk37AN1rn16hij0a8w7VpW3iulTLbHESe81Qw
FV33ZgBH4/8vJrZC+y312XtCy9kGKK6BvWfnOZexCYeeFpFJoXBEoT8n7v8zzD/G
ons7LvZucY6yTHuxW6ML8lr+Rs1oDgz5YPrGvAdCA8dAyfW3XEeTguQY+NssHlfv
3a99435N0Z4QI9GiYq0shCifSU7RwRV6pxY7SFhxUxJiHZXGY2KxP5q7RSTlhokL
wzIvA/jQ2ae1qOLKSbbOrFCLDuK/WICMwPIvigV3fAnMcJBA2oSJxOBPBw4v5QfI
Oo0TL0p6z6yeAXD5ceDiW5UbFTbpSgmT4127yLeLxqJrlTj1k8Sl3HU7FyHg1JwY
WBTPdRK50zW9Eh5hRF5WYYnNpb1KzoYp9bbDLgFWrSqphuivU73Eukp1sPMBHycW
rxK8plUAHfUnjRW2MVP3vewQPUFNYdXShH5OKlFMkAuLW3I9JFxf01jAKfLlvefR
H6KQQ0xOnEBYEzLIlY86bb2imDHYwoDxYTpssHSKu4803WSZecOEDKxf6anFUYYJ
FZyf/fzoU1LNJdOx8/k9+2Q9H/7EA2YfDvCFypTiMIktyH5mjrg14RMBRlyTc34t
TbmOmNVJCxCn7fFxCPRaSJ3Q7AMuhr6+xSg5SYavqdgeb8CnLaUklojcJizvPKsN
NekkFG+pwSf8PUqgXEfbgzXZDhjIRVnQVT3CrfFXlTlvFFxFxYlJBkGb9xotSmmW
yTEKK1FlYekP6qRiedbM51JhUFpgqgqwGqiNamSrmb7HWFbvxu0RhBc7jPMVtqac
blhN/iB6ozXaUccAplcxAyn4cXGrIAl4UnrBHuD6RAtT76YujpKzO4dcLFzP6HwG
Kvgpz6Oexu+UZ2PFim/gha56sHTBS8NeoTagBrtuX6h10eYVYN3Vkq4n+G8Nzpuy
+P8gfclCf8YH9uK8LM3qJvs72RIjtMdWmo891qXWeRp4zLR4jVG99mdAEah2PrV9
oS1SD5jfI1/eatj7Wj6Gf9NR/pmO1HMuJU6bIgbqVvZ/Tju7zdIBJ+aXYqfsqkru
RB78+H3XR9HLfwdrGvcnSOHJK1jll72+J7pTCSaFEvYH+sLJI96PQsJg4EulRUHk
S7nNA9UprDPizECiOYlSVpyOB3k6SgHtzNcxoXGGfeL/xAXBCewHCbUzMAFikgjK
Ak/sD3JMbyAjqx39giyrX8ZKWyJ+NQ5peQNP/xvWL5C2cmW5kdvhNaxgUy3C931j
py+Qr5eLFxIwHWrP6HzcpGRMDdH8pLdfqU/YZesOlU7Z5IAHusUERrGMBv9+EIJl
+fXySbMmIm3nOLnrXcoEO9QkADB8FZaNH0x6Sl2dIwztUVME3fjTPf4YV3RCoKJa
8h5/k8Yk35M/INFHLBGYoPccKkRpMtY0Eset9dLpDrDt3XygWp2pROu5vhUtzcF9
JRlHnfQd56LouhH/TckCyjxOtiDkCzbdQ3vwYygnk6+q9+Hvty3JzE0ZjD8Cg10z
zhUXfL4wPpw9Jkv3Is6WQe+7ZUGAGlJmTDwi4bKK7YaLGVlwEJByuq3TSgxzCZRq
EqxbHiXRePO+FH1YD4Ww92KBoi/SiJI/1hE5/jA9XcRR/cLDLM9vqTGwfMe275Zf
3mCSk44pEEq+NN5RiJ9P2lJIM9kZPVP21Krh3LVyzz4jMCG2dmh+iZtK1/UE2pj2
mz9yB6BYAXjFoS81vdnufD1s4e3zj9Lk9D9mLDa3gsuLePz1oskOrQkkUE7Djn8F
l/TwSbym3/kY96nIjQS6hue0B6GHjiU80ZKAsBy8sGy0l/lcLzWWr78VEW43N9An
ep4vQdDQz/j7C22yaiYds/7cTKOD0+c2vvI2AiLfvD4Mz/AIoL9F898ykJ/ZoxCf
EAhhmbxIkR46WaRU1+WrIIXvH8gHQwa7O/ppJ/OhitRWFeX4bWMcLYXQ2w46k9K6
eyPy4f2IvEULM0LjW77i2jzu33dabdYJHrClTYMeunQNkbaYK+Qs+e4PBxtzWNR1
p8quYNaS+ok0BQ/F13StBrVIM6oz4Gbv4nT16Bhc4MkJEw9j9tQOcod0xKTXAt89
kUlwP593KkXx+aJLBJ/Ox4yhdZ37WK0jb6e9fFuKL9DOe0wvwc429bwbtJDPm6kR
LLdjvQgfPksB1yo85YmeG2Fs4f+KPykNEAofBC41e5BsKWuUsX+K+wWvTFxBaGuK
/ZXINQg6Bs9ITQ50RWa6J7iEKNjmisI6aU0sCMGp13eOa68jAI30MNFbB/pQSu/5
Fkp+/kmiKYAPYJl1t6d2Q14Jc/L3sxyc+dKMxmQOtC8WIv9bd3V619NgH2OPwnhi
Z6elwqztIM5/5q/LL9kRenj0HExT/ZHBNM1fCLb0/N/2uLbIiANnHAiNfxf8qV06
AEPaEnL28EZLoQGqCt3DCSbTSYJEBqfV8+ikENKWdY4wcjkf8gQVhoInJJJqCk4O
f46hPEmDma6+SAljAYId6lQWEUKD/5oWIPpaD6U84GwGh9cpCg3ljhmLbETUQKln
7r1vN2WoX3P/nHSCloGN8zZhvp8pvCR/4S+gJrWBjkl6BXmuDel23ugNhva6uAGe
dmshcPA3XjDvoH6h6ml/UHA5PGz9nL4SxMtXmhQDjGWBMzqHoKdnSz9ACpy0VlFC
cAeGjzECXx+1Uyd89WDyQ6IufDwpTkOpJYumUwJS+BJSbBTJ53B9uDjiHOl0l7QD
jWnQWzpnDvkRBK4MDt5N2Ff5HhFkaerP5DrvocMiJTftBUAjGAWF3B2iXj5uiTUk
o+Z3Cq0qEmieM3XmolxRXoLGjR8Oni4LPx5H/WO50uyKkgSgAGiCzEqLA6LbxmiI
8ZkI40GVo+7evanXxWifwnu3mBS02TmnHWxJ78a3N7GVtrSNiFdDZPofhaG3MB7b
ed+3mnVQRPzMwrDW7wGECngP6gmqGeXA9aG4VnmNvzwiou1CuYZydFosxBj0rf86
LIyrqigW0AM1n24/WdqHxiI5IpQID4n3QAHciw28HIOc6V0dXSPPvIzk3UTJokEq
HS9GSXdiuWyejGhQbSBsyjNQ5cRdU56xyj+WdE/K3UYsF0iWXQ/71FWhYDwVEMmS
cVL9gl+Yio+cPwMib0z9mb9BJ2JH2OQ4k1lD0dahwVZjFhjZMQEHDb6yHcI7xpo4
Z5v7G7JcEidbW7RNT6rFgVL2U1uiQkuTqmCoY8v6KoxHET+rCq3Ht9rtxFwxHVfl
eh4KN7VFsaYzB+ep2cATO4cXGpVpt44+bANyYohWUTpPHrh6T0rogyLAzsgdzEmw
tOzwJ5MkO3k7fngpX9HNFIGcBlr2N1j5jHD+JWM1MjDujMcnwA22XAd1WaLojy1D
+W5ZiMLyWQjYTBbGpGweC+taQWRDu+NVW9GBjg7eIdLXoSWG0TCExYdaVtVSA4DS
JMvmSRMK99S8XRLT71AFyYDdhLDH333O29BHhG7EyUulzo8eSGG+apDkrBurtTHf
c8K9hu03fQs/sDp24WvvIAGiCGaaRI1mJ3b9ZJlQbRM5SRYgSBmDxmBaKYt4fJxS
0GrCKlpFtatj2lJE8N0+ssTP45jgvVGCxL/vVDVW9x/bFQXeGdhZVxCqKBhEujoj
pTuSJhWyi2lJYZKWDz/YMAEsT7tObvoUjPcNYCx7SiSp8y2WtKYhgbnpb7gbmZQe
X13n+0eDmYh+SnfmGn/yc6jlICi+H8MII3XsKslyKJHxb1GvfSnVNKnq1etRPpqa
6hHdWuBtNDSpmHxHuI0CXMINHtMbNv5HSoGF6GJJNaAAiONRsCShzgoNlnzG8KRS
Pg0oUB/gjBvVp1wY6LHkKNoR/sn/gYd/M0rdZ+G8YjYkF0GtmSogHb2+yrT26q9N
tVJ5ZJkgDeu79YbB9Wb5/+ZyYFytRTUZqo0ktYeramMpDbu2/oXQq+Kt4R//6yiL
8P3idBHpEXm0djGawx6z5YmU0ht+jBGT9OJqYf0PIqY8fKIBKU2ctbHSK2lDK/Xu
q+uHhVMl9NMYeRmUPM9JGsB5fPnBjaR7kJ73FaZYWESRfE679Ptn0qn9reHM6eGK
87ExoBOz5NIqT2Aw7T77UIk9jKlO80lNpXhNJI7/L20U0hPVKBdD413SihvRGHup
hK/SAVQ1uPagtnZI1nqgN6xVIc0byYGy5i/KT5Uyu1U95IHqCnsE83BOnLU1bL1/
02FlqVuyKuU7mRuJ4NkXY2J8WjnZy3KZ2hhFW4XyJXu5nGWU5/vg0yiHSWDAUKZA
WZ1DgtlBKSsqHpGw2m+l4+quD6/ErKImedsNqrS6gpr560/NZE5esXPn4egHSXoF
BKGNsUs2r0KRLxvU9jZSLl6cBi4IRP7OBpq7hyb44VnUT18GOjM2z6b5SVasBGHe
lNs2aGRGoqeF4U5vZ39O34x2qHZsq4eX4Ms5kFpKHEALZl60/tTmw5KW5ODm2C20
`protect end_protected