`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10080 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmUFVhi5mMoX3yB3JgBuKJm/
sz33zlo19iGE0uYXRzR37Y94yhJAImqfE65axpS+WNRC+2ADB7mor9zS+LBJTzw7
cAfIiHx1wWhPi/R4C8jCifePj+Bi9M139hQHgXvr/TMdaTvtrFQlykumYT4bUAmo
rdsivp1OiYZJ6MztTzHpPixmyqMyRC66olqIURHLyZbJw7J3/wJkHOUV1oYqHHa0
35vhl9X6ZRPCJ5FmQua0LZzNB3PawmFBZClaAmUWJVEvljAImDLAiV+b4YXdZed2
Q0s0WjN9xbOwwgZa1mrkj9h+p21ZvjM4cef9WargBqJS50HLtxQ7lnTeUw1nISNy
eodMN/jTLP4lakCIm0GButAnxZ1vZxyhNr17jHkXEqozJyg6HuPlpKzDF5vCzXrW
cxm6LcVyJcOpG9kRUg1Fn5lPxkI/MEtSRsNkXcMAzHC6Ab4kd1W5DoLRuz5H7w+P
otC+VV4oD4AzA//cLUHfBcJU8Yz3dS0GdTWTU867BEGbaxvGnfnidpqcA9vNiB3R
gYdu7VX+kUZM5JfRTrOdt+OKo4m4SUwM35Mhx3TWnBGcwHEbdvUgoTiGy+Vd5SFR
znJlqs2t09e8Q/Be/oPn6PLhAWPIcdr1Zci4iir2ejk6QWBuvZEybgAWdkMtoFru
aC2iseniRubahKACLuvgv31kIJaibXqlVg0NmIRGObqyGl1+6/IUBNbBW7QWwxMH
/wxiyfnSWxNvnB3m36jvNyC94o8Xgrf34Vzfi0pIwiU/hJpRhj6XakL7/VUhoXIl
B8ZYfADyObyFGyb6U6DLHzYykK7JQ+9X3NS/BmCTStYVD9fpOAFpeaSIhlaU3z3F
QyHdrUqLvMf7poIaWhBB/SL3TforANFBMk/3nIG5vnuIikGa3zdgKOLBPUdootxx
T0XF9nNSJNO64v1kaQVEfISirGGV639/0eFCTc5adQF4dN8qXYcsbJCrlPUxgljz
QFGzJAJhdxl9aeXzPCC6YA6d+JO8IbGyBs4QcPHjjKCxJA53CYyF3DYGLUYYwxKh
cfgypKdvmdTW2ms1mRSnPDbo0DdHU0rZcDe1PazEIJiQtk4XGv7YoZT34sz++qnm
GBZApCvW/CUP4u3/5WQXoEpoGYAVnbNxslU6zJ1hP7R/nAAUtikPCconaCs/RI+W
e8zfoMdSTKlf0l+hGQ5TUoI9Ed4xBmOc/76OZ2wlzzsU+6rRjLm2LyqiZbrwguhN
Eu/oxko5qVXboXBAAaBpA7gC/fBFPW4FAIqIicsNqrtzLxbH/mnexk9cxCSatB5/
/n9W4r6GdAgNvYR2YVEs/gz+IrAc+Q+dYnBQyp8BSN18CPu38g4o2q0RP5LSJRpa
mW+lGDz6JmAAx7AeI8hV8NnfvJcy1skgAXLz+csJSI9yjFVj0fbW0DBPNV2JLDgH
Ihhhqpovcg0xx3wj2t/2idO3gULzWVGmAkHcdynz1KVDXv3nrTenB8wmn5Tm5+mn
PQdw1Sst9XzV95ZwNpPJ6hvDVQnwt1PCuIIlyqNELM4ojLGwHYdELcq7CPATtvXg
mCkS/MTbTMbRtMWzaGYE89sdNmoDv7vRd80akQVy/vtv4cMJcn2txqoqxDrLiNZH
l7w+pyoSGUXB0oOkQpF8Waxkm4FB9231clOoPevSjTunadoc5Q7Q4gydkCG9TEyp
AydSWSMZlyAFQ+ga3F4iChST6GPnsXaGmq0o4uqSGK1dN8s1BFcnVdOB58Z3Kkcy
DfX3iSD/lvIIzMXq87SGee9iynRgDHkz+z/0CA0OXS0q9EFaJDZuOBR1Mq5ox6xt
s2DNpavUP7T82OTLZ7lkJw5iLKBXOGS7SpBd4LNw98vxvySnOh88xRQD/2bHOYjM
wwrIBQqvPdxa+ary2QmKC1eJCh7HuP1160VdGgyApztli/Ydl6Bwmq+amS1nu4/t
3Q1PQaXm96kaPVnzMPuRO0t5K4YpWph60WT49sTgyQLZXIN8Df9J2omxguDAlAvD
ErOUn12HIcar8qsEAnakjPWPjJK33YlaNw+KQJAVdqOV4P6F8sjsYT7ckSb7JRpf
3R9k8hPfjCSZpTXl0goje2IgJH9I0wgsVeuVZnW2trHHc6GRrY2Wbjx/yldGA+sy
TaDlvOA0YQCMQawA02ZyaOJlAi5h5sSCfH74OuTOFb6tNZyZW/GcXeINQmJaRVHC
fQxEDXurJHRrmOdiuZoy9We9fDKBDoZCQ+fthbbQVQ3STDfYldImugRFgSI/2lse
TnhKiO4Qtmz1p+K+keWYaIlqIBjT7vcP6UdbTHrRyHo0pErIkJCexDhdtWR2MEEQ
BL7BenLq+X1TvCSgut24YNVvVuH7B+LrMqaut0SiSDjUNlprfHAmCLdLZi9ntEEC
v5fMAaww70YdpcqSzrJ3fC6tCMqw0iDgoGz/jA9QE91kkETH8/CjQvsPdd1gHuCc
qROFgjNVbVx7munPsbS8hlifVtHzk5786rXgU/OzcyZBwUEihuFsu1VwI5Hqph9c
9+048QceriRbMHQPmu8lvQ5ogbKz6e7MKd6r58n3iG9xWnPKRbMeQItheHkTjnwy
DteKEgVGfS4CRPWoP98MT3iiCWopNmVrgm/DNT3SA8wsRljqu93TmjLRUNRDTWtE
SWA2L/xeIqSxisJpfIKlQ1F5IIhn0DF+ezNoAXWXuppqVVVLhsrL601BXnV/6/AE
5pSQ1IbEzF0AfJGPMmpEhGA94BSb2N3SStLpUa4X/DEFQLZelAz2iFEmuy5QwExn
6vCFa6IBFWKUJpAJP54WOBDtGQLH3ht2O6iQ9OG6yWiqGKfSdFe/9FgFl1PCTRje
w1ixt9zPS02lCW1f3NBoWia71fjJS4AyaWJzFrGsblh/qk4+aG5gpK8DW/hhtYEc
xOrMzEPCVrbUhYTgMW81Au442wcac1hKJ1NTu7e+9RXLU+J627xLsg6c1rwQrhuQ
ByySKXyTwzsJvF5P4hAgt0KCK6l6UAmNS+6vHG8m6NL1RD1da6m7NBva0OWUJVa6
m2D1AAaaKuOZt3vE4IueyvZHYV0ihPBuyHAJ137p5PdQMJk3Z3vs8AHYOVRG4Gmw
KJhP7xY7pWPHGeoNo+5CQSCGGoixI3jFwRLc8LSPy3KACQiQcQmWBrdyNoYXqeZU
Q+CDgrPN70t3HsO5LI1M4b1qSTTP/nzuL+rJmtFhV9MuiFDXQl/G+Azd94TYOVrM
IKPIcNdmH/7u9Awxumba6OOpn/J1JNBV3TuQBD2zqahdlQ39uILGCWEuB1zSBi3W
rCUYG0+ljWhJ+WnBQwcIJ8+Jqu3I9FpnEzgeQSxVKOVDB2d6qVaYVC+c4cIqVts2
JWk8grO/ZVJ+oJpdlxMgbW/slmLLDRfzOSts+pZEDHeWPxN09e5jQiQG4TVKT6Dw
XaTJP9XyVDsvXStUn/0acvgGo9bvdWvy12sGlRMtm+lZsriM4mGyK9tJlajjze5T
JIYc2VHSgv6Ddd7XVedfuGg2L6PUnqTCNq5KkG/JIJP9CYl2FdTRfqkn0ji5P4UK
kRbXYC+PUkWv6Mz5ps9xr/ueQdSScLs4cM7rhmHdOZHDpI8H+YM1xlgLr4Z8xDcS
qnMbDUm9tT6rsI6JLfHUTv8FW1ODoCN8DuMu3yZACEc7nZ+mS8WU3LqEST1S+nwv
FtgGAscbWCVCY1YwoUPuETGa9Yj4xjlzmlqvz3TvhGi7FWXEz+lD3SBDKwT0Q5AX
YU+jQw6Lu/uIVxp4MLVO1ldTE4iy7F37axiJb5cScyd5gCSUlQShC1+NjMW5SuAJ
avGxBZCvzcbZTgJPdDL8W97HGA/6fVDk9mzheJDw17EmLqYClcFFaY7SvHjqV5aT
/xL3Ln0X6MzghsvOqFtAzwtzaALUXw64rgjhv5YmcqwUdQsL4ZYQS4EzFGNNEqwW
MAMIgoB3e2PYrs9tKAHeigWRSXaPtwpAPtSvVrvu//9HQNxmVAO5Ni2rqy5rGLsd
asN0ctWYUbUS+MNghSFZuWRtu7jz0o5gnX3N6qHBKspHU72iwf/kNx5K1oP6P7AT
5AEmW2Tne8bVQSlWymvTXNso82Ze4ncIZbIkLYfNoBy4wgCyDQGIlmy4tWi7v6i9
EdA/6NOCk14MruY7cNynd8UKZD+2XxigKOYWHPHxtlrQqhyoyYasnMSN0ISiqaTL
146ldKp7Ka1tdTlpE6AyQwSqe4bQPEfmEMo6m8D5tsRli++NQ8gOWJgdRrhPivhP
QCx+GdXicC9L2IAraYHzJNB7+i7d0Bcl9nDRwd+UXR2V/7q0EONvtx3iy1hnxB2j
BnXl3RrTqECEjr6AoKAL6V6fbCZtsSsPxebaCXakTLiZt7pIOcLivfwBEKB9fDqu
/xhGUaKN6hGOTKznSHKbS3UMXvbWICiO2hqMfY8qFC3AMVb2HzVjyDbvezY7ve+L
LYWFBOaTjnotaFY3deE+/vnI8Pqn42WD8l+qXDNuyUO/j25knqOe5oy7uosbruXs
iPeCw7sFrHTmXcYc3l8Ut0AtYy4L+ZrR5jRfNYpB/jYek1lwee8V5ePsQdO/4pJL
40dgIH7Zh19rhIft24DuPXtdIzdt7YWzh5SoViAdy8XA+WIxKZPnIw4zcQ/bpibz
6RaTl1yWfVwvlX2BC/Ja81pmMb52WinBlPPYNbE8xWdmv2pVbRjHEhQMRYRhVV+1
cFYzptLJpQYJZ8i8P1dMu00yb/EnAA43/IV9YRLvnR9ZRVXE2hXx9+S2oDAdQSCZ
OEK/U+a7wcn7FW7zvSLIOkZopG4mBC3kYy7uCnK0NFyjeGQyf162+uyvrbZmx3RH
CRnaLi8SZ/CF6Vz4J120FBAqD1IqeoDKrfNvtz6kmba0qgegFPyWJi6HROz04uMG
W3WIDyjvVqMpEk1jPEkpEYC/aKgoZ34GufcAc8f6ZjX6EYOqqm1y+OAW0rF/xYJ5
BpWfsvmPbDML84OaK1M8M4PECRX1QISJR2gqX3ns4RstHa5Vabtv8tFH+RITHOqz
zC9mHXxBeFHjr6SWhJAinmx+P2IUbOvyTdX97q4mwcVaq27XG8oSaSvJx9tm5pz/
cBkQoMFNqIh3xsDanVFMXe82i8A35WknXuIO33uxGFQDe7rRiPCFD71Mt2bAi+of
oFIJzZGYfkiW2HHqxLbx9S+8XZ1H+j/jnni1VMGpPpRd+CWYQ05k5VoslANlMswg
K0sZDGnq6EfqPTvLJldVqfV9t6tOPfYDQ2cswsdgTvftPW5KfPhpYkcIhhIAowpA
5sR5NLu03cGna5xj11Zex0VrUdHiMitTdIkF7Pmu8dxVLrIP6v2EuUacJ3vgt9wE
ZZwSX9WzFJpVSfsc9k4AvT0xCwaFmpaR/a771HgkhV07Cv1PK966/BYFVNurewKT
Gxmrur2ZCmd5/OLgRNkq0ipuWMNSThDMlU34i8X4GXiUwaUa4vei+QIs/FryQ1TD
/O0n/m4Hb3WNp+GfIPfcn98xsV+J/qTCTPhQgNeRC1y09bChq/vNB43Fz80eMNPM
NvTyIPK9kapwnVLfaZe/OcA65p+2rOGmquWUh7IoEwwkzYAEfveemBEBc6Szaj9a
Bc2AmEof/TkAshY2jbJyF/jFblKMqVgiSkjGWTMhykalMDJaPoV6nUFP3fsq8Mfr
TsfaU6XmZcOR3MuQiIx62QPeHwFuUWnF8o3rqy4iXRHgjUcTHOVC6T2bV5kim5N6
FQXZOKs0qAR0EtnMR/5qSWv5jut5tnzo84npC0dZUlNXbzFTr98+F63rNYr/a5Ou
Vx3dEI6NqQ2rGAO3+5fu1PTPLuaeKpY8SR5bOvSoE59HFuqd8iFEEyKt8Es5eC22
AtCZFffAsDwG/60MLUnfU2BjvIe9qTlg4igZGmZXuit4h2CHJ8d5fpqj9mKSFC8D
/UB7N87pevu9g+mqYuhbvqXNTJd8baI6CtGm77srFKim3r8iQTr27UPzE9ooZTfz
QvhgEKwtIYfeECkxGosji9RH+lWcHc5iGh3zX7l5YzUMzzq3cGl4LHLxdY3LvtdD
XKKzr44PDr3JBPp6n7MHYtudQ5mbXBMxs7QbKFoZex2bbTa50Ai/WBog6cVX0Zq2
dXbgkKyjbuy02DHmELjgFdvZaWcJu9W0gilqrRGz86cliF2SEWlXQemxDUAUhiUU
DAcyFbft/v84Ul1OHz8snI9WO5PsjHUr31Nl8l7WQZT9yqLA/WnZ135wqwgcrAcj
YwEH08F91nxIdAGGeQ217d6IAZPk0HRRN8zZCdAA+FL/vKip2cw1kl/hzjhbyw/N
n+y+B7wzscL/f2vXIIMfvVxqQ9UORIuoa0kzD5wk67W/NPs1gT1M+yaaH/Ryf1KI
dhq+3CbOjtiwM+Q5y7jA1fNtRhz3Mp7mX/WEIfWkPp62WYDlL5VpJizZ+EaFz9py
9NE0zh731aznBwjkpcuFvMuqDvKdZLjJCp6kttVQHVcKn2dCEZE2Pf4BjnIc9jMD
d32VfawQIX9dCXRMj8VDGn2cutZyBS19dUxV0kCgU8XyumduLTgfMM4Gmnmu1stl
Go+LhQ0IMAhOp4zJRtX9Oq43blTN2ZF4KDfrSfaQlcoODQbQfbxwn/Y3VmIrtcCX
ZH1b25H2OnMfS6B51iqKgxqSBAGngvWt1WtCf/KbNPudmj8jGFBGugH1t9Cyfwis
4DfjFpH+2aiZCLIW0qXHMux9NWSuSh2j9xTfPLwK2uivYXRMXJlwaBrc4HdOjwEy
q9jrSs12h5lIn+vDidUZLkYiGRzWYby+c7b11yWbbiThRePMJbAQMDe09Nb/aSss
VkwYzVYkFYRjpYXqxgRXnp/i4R1uoNaNn+XRhlq6DA1gKlEpEklkcRT+Fdt2HJOs
8vBzVXQ6yEoQNhTodBuLI0ON9W5ipFQPv5MQNg9M9ojjrqLQhC3zb1aC/EL2wlAm
J6CTgMrtsLLCjtQYLUWunwxBLZDj7J6hlg9zLIpcNUg7YaqPI/4wj5z6r0ZfPLCR
y2fTKu5E5f2eeFVbCoLmFL3WbUo/PJT86ViK8ZQd5GOzvwNLkkGqJn5DTO5Cys31
x5MYUlgAt0a8lvJcKwVzTq4uEN2XeWRIYG+ZoFPz7Qd4wca8itOCgqoQNK2jw441
pibSsSeBojP7OtvjXnCU3hsT/8zMXmwn56j/SKoTCP4gtDXitTcr6QXq2IY8LJRj
xg92PMTx1t6wUUH6y6bZtiNwptKMHHZoYfbbhUN96mD0diBI2UFnix/M95ubVOkU
rYIPMtqrUGMky9+mUv+1kG3C0WTQUmLIzijs14EzuQWIS/sFFz1Y77dr4U/ap3je
IhTdLEhvYugyevvstDIVs0537hKX91bzW5nP1RumFjzZpsNQGFZ+WYjYukkGEMxx
eqgAojzIZhBV5Q9aAIIg1AG80R9/wf/0LDE+FttwaXAvxV2SgCtf8dMbyysXZ593
1prn2wPiNtvWDqP+wH5AcHLbB7xTcjOF4AcDDtfle5ZlMaQeCGzJcqTxRx9b6q6V
BMxpJgJ0y+aBAJ6dF+LPTzCBZi37g0VPlK59mbPJzLbPY85KJCv0uKlyoOCpN/b6
e8Gn11nD4Of1KZA4wSTRgGx0syG+GHE+iXVo8Iwl1XS1YdLBwWKRqI0QbsObvVPx
EW8LaPzxw823SCbBuTdU7Co4Yqu3McnxT58/dxNSF2XkbOwlqLSJR7SAhEvFsFvy
rOrGsuV8ljeSjmRf5bYYnlZ2J8Moq1H4DU4dmpnZtJkOGzgAFGU/3j2LWOl9ymzo
uMEREiidwZJqSrIRDiBg7vD00QJgKMhLlHysYnDm3T4dsFcOLte7qG5nJDST24r5
6CvZDhAktsAkCSVP84fRy0DRYYUkTIKq8SNbNu50l5qYypOZV/i3g0Edw2ZHCKv/
IE5yL1bwIrXo+Cvtd4cf5jp/JPgfEUXvPvzdKfJ9sauQOlPBv5GdWEYrg/rxxWWN
G9qYXjVzne2BGnHwVl14gluddIVfrK6xHDI0bHTQZdu1mSb0JBSt+v5s1uhBOOKn
LQ4uOc0Ht9eheg6bJPElqcKpyfwHmZKERCjOW7u9wGlGrJMhyt8s7QIgQcZmRwz7
haLbTFUi0fiJuKJQyIXd87bO5ODbsQZX5Gl9iT9GJvAEJQgjTn9KHyMJd1sDXBPy
S4IUJIc7nXt6RZJ+9FinJihs6hE9MVaetb8nIqXnXqovYGHBEgs5ikjSAmWxEyqG
WzXhfF+IBHZr8uK+RrXX8RVIKFNy5u0raY/h+OUCaGhxLjF/1pvQke30MiMckIWz
EOXUmYarCSTI3jr96peB6Yz4ANk6LydLl6VNfcCmpZAg5jQYFFWpfmPVD9hbGtW4
y9vTVG8mrybbdrm/EEPekU8/4YLjvGclfD6/ndyRTfE8fmzU1eMI6/HbTZsoJWwR
no5wdVup4GJPWfJLy2NI/hiumqZCxWMYwYIGmALpurSxH8ksvpFgFTtoGOIfzarr
/6lEEUDRhVSphjeyRUkgola23DrLud1SbxA4CQIbfq8YmAV2A6ffCl/N+g/uOTV9
ceJEgDOxlh6SYVxBK7uW+pRhR6aC0vU/yDjFiqDqovJe67AhPTe76723DKH6hPv1
60pBYhr+X4g9ILFZeGnMM5oAiESEFd9aaOlhRJM4pYzxPonRK/zxz5za2nMg1a+0
zKtxIfYyk9uR8YU9Gnj/O5ffnu0mVjMCE4Byi2myw/y5kCDLZ96DTfoi8XcQ6HJq
aeWC8gpY5nme1Q8iplw73q6SzA2IJh/A4rxIPJqbdSrOLDJnyMSlMOPIajuohli8
mZRdgcxsfSEpbbOFp7fcyRwIgYxD6rxBsYocapnHRfPllh1DYCRBpmXJBZtb2VqL
Nseqnog50OjR3V79XYiHwjvf5S4xSh0olQuomaf7jE99qhyQQEfhN+4j+Zhze373
e7wwIszmWCJwR54J9K4imM2GloyRQwftJ0SHmbYjEcyTg/VLNIb18Fh35xSYlcWX
3mNJSl0vkFEi92QVnY12X3NqLgof3Xjlyl/1URsnibBc7337QzPySacV25htwl6I
h6mb4ZBCDktKl8wWHJhPcFMmRPxULLJ4KPJv8sYTiXAPCbNTP0NX0m3jl93MAmQo
4JDZjluPiMLUFmm4CPuXHqjfrukADcNKKxYGjRZAPqETfia9hN54/Qe86G8YSFOS
oqVCMW0G4Fuz6EHxpKSyBqFXFq88ueTsAG/vrilnV/Ht3NFJA47IT8IPauEVfcTa
p2npeOGgiHqR2e4HsOyJ19Ea1nroBxKCPYTU+aIiKBEAokNSI9H+gvzdfR17Ig1W
BZxVU9fUax+4bzkp/hx4eYZLV8BtPiZJvhXlNsNm9ycbwRcMDdtLz3N11hUkwff3
ro9F+gGiHJi/Fk0hvcuxIPJubmlmVhmGCW8Znu5Ls1VooTbpryH3CYOANF5FrqhR
i9CRWtYeZrGI5rNcnArOenys4z8oJBifNr2zPbWzqCQ0Py0EQQpyxTXYsLyDE2iJ
B3IiwNKUNTgaI4cRwYocVSAuV144V55z4rUB/7HCcKx0tzHN0AKvn7MStXEVYH+U
e7Z9EBgd7qsBcXXTw5nCPOVZmgPYZSuOLISY2yn4dEWrpcP9/UwYf+ZHyLOahEKC
+LdGHeQMpPkxr5+3Nxh7NHlrnEsEboBNYban+dm4/qSE4nu4XSy8E0gk3icFyTOR
WPcywKeWmGc3EbLGsfSDp0Bi+p6dNo6xkF2nOU4l9rXAl6wKCpBb5VWwP+Y7RYhQ
N3LzId1ZnoWOgDEoa+yq2++ZPJXL2NpXgG/sU8x6Nt0yuRVtz2RhlHDERBSdPFDe
XsaDbeF1NnlDXafcN7T+J3bO7P9I9QWjIIFJ3x4Ts5+KsIDPzFQkSpqhcG6ycY/y
6VNgpcIIV9p5N+vM/h9d7KV0cr13nYQl86jhdvvqHkZ6QmFKtYocE5fV9K64/AwV
BzuL6rf8wKDOyxGpMk184GlyDF+0v1JvOvuYEJs6CFDc+OLGp4nyengO8jEJea1l
bZt9Wa2/9B/ht547Gfi4QiAa+tV6wJpBwdC5QPmHrr4BmOHPnrG1ydSI3WNtNDK2
o0eLIWUwY4ed6WTkARJZ2l3ZFVM4jPsrkQbTpLR4rxRWk1ogJ8otcKbeVbT+P8Bc
ozhnjq4zU2ND2+rROu46h+KYJ+Z9OqYGuav3v/QSe0SY9YCWj3vocFfoZCeKGsSh
PoYfrsDome03XYhPgH3/7OD2FChsxY4b/Fk8dJUFg8p5ObenVZ83OCTEyIlfQ8Z6
gJxCbgnJUe3nSj5hhA+VbTklGQVs/T20M4SdAE6j6gsObEdehozxdFjgSotKtn1u
FQBIm16HPUPk7qKUOaavZ5FiXTfwIQq4+97PfuyKU02YmsvO5HcmQ8c5B1hkksDT
MA9DShbo396PSBoFJnjxh8J6G2x9PyG8Ze9f4HcaZEqm5U6uyYd0W8Dk8lxdGcyK
ZE82MhGSptywZ1498vXARphB6GaE55/nK6THlKxXCTB6ewRtsTMHMcd21Abe6isx
4C76Q5+uCgjTvwIlxWynhx/94rqa9FvC8OxNjG0/vT17NFHGXm5S16oHK+4yAa/c
6P0mWoMJowN7kA2t8GrX8dInLJ0rzgLzHN1J90ruM7wzT15VKc7tzWSSgfCUcAXs
GbIz+fCjlBOo/C0Ts0rDnqui4SQthKxMkhyVAF5yXamx0l5kmvprbkzUXfO08jiz
jXLlgvDQWM6x5FLj/+qy5UluUwdkt9f1B3cq3cVwgRTXLgMWNZARolJPjXzfc4jR
fR3DYXBGrzK/dy1CKc0dzfikyRsouZEk6ZkSAzF4/hDkSd8Kz7pyw/TcTvg41IwG
Vg8hacL3SWut2UNraLN6gzvVdAH73Ar/WDx22cwOoDpwV6Cyw7kbk81tw1JopI8u
ZrXfJMTT+ssKvnzO509a7tziuWC+W85mnGMu5rkdWJIvANurA9b6GyZNovEHbkxK
ezE9pPJM2FhS7JU/NK54TBBClMwGnutOVnZ3Yymr5tjoA6PiCrk8wEebZBJaOQXw
1zK/I16YDloaqUi7PfGFO6GGDrE7MBMC3a5a4ousnl/UtQlQL+zlSgqei8Uku87m
N28TwG1hPIdwU0QWsaq3QPR4eNxuZQuOrxdYQQTVawI8kmTUomTrLRunmkAJId/7
kZ2Cvmu8QiGsB52kctJQ84PdR3dgD/FIeZw7P3qZAXI7+KHzxCY9UPMV9pL62yVe
JLth5BtMhYhSP7thKAxlAbQEuZ73qaTIf+IiKHE/+HwLp8lUu3LPf2gWS0BVXcR2
l6Ee0dOB7Q1qnRVewy1NkqrzwZmIA8FZ9plu0Qrtm8dbmbvsdSFz2cv+4OBlyYzs
eVF8pD+Z8PFVyruWlQ+slS4+7dh857DkrnvCQBQtH2SnVTTlC/2/2aVDbA3/ubX3
cj39YugCpZILVCR3gamRGkn4Ck/3b+Jctd2nW0EYsKP+YpjCfKr3MINNOWVUegfV
kKXdCNREjLQt1NliEKG5w126fcDQ51cj2zIBJXvW4GscF+4RStDWpAOsZlQp4f6M
HiE6zy2FaXqI6Uyu5dh1PHzRMONrI3n48KWs1g8zQwuWMuNyEzknrG7BKFqP6rys
DZt1bCzyvbuaRcEBFApVVBhwLMVF71zfzm59gprRWePfCshogkIxoM62jjLprNtY
KOwZQWEXGqeJAMzWmEBCXBXYli/2nLZw/0pTk6daUiv4rJRo6/5KEMEyp5QIdgnc
u1sTXoXixZylwvBC3uEZBDo0XuFr/JRObtwnDpHRXQJxmuckFjQcATfuaeWFsHxq
o5QmvLgpoeih/0OI7mUX/lamtE6fmyP2gy7cAlTHwgtvXwBGQl1VNmZ771HOT7ZW
Ybz7BYxrO1F+XVGb1Kbd+gQoSaEhXCQr71bXby7bWLBWNu7lgQf0kIPc1gGv0DZK
UCs/REm4EZjztARQnRHhoFXrGIeSLqupPmWRZm8BmtrBbE/wt2zdU3Lef8quWR0w
qbqhB+izPcyCXbiy3aN6TPFsZ0dNGqJO1oPSsReO8gAs+7ME5plkVFxQGU5r8uEC
dWmdBgZWILSPY2tglQGoKpKZkjWiAvIC2mJ/UGOfrrnlUUvgdYv3udfmrnkfjzWe
2O3b1N9BYsixAAqbWdkE3ETusqsoobDJujqQUX36lIFsAgOVDk0GS3DOzBUUihca
uvbr6t3beYn3wlpOZURLRW49wilSr5uHJrTxiFQRbrYuqbJegI6fc873VmiGOCHj
Ai1h3CDbtp2n1dkO0uR3b8d9yrjkj8hu2JxIjOUwXLEonnbybSfUuBUcEEK6f8Qg
n1LdmK4KM/UeESzRpKBcuTlKCluEB1M2KAt+KKCJ0ZMcTc3k3LN3eHeOvsdNP0VY
6fj7dzW6kkU+1VD8U9EMMBqDUkZ6sIbcDRi37NZCQpGRP1wZcjgmMQUwyCte1WbJ
MRiJkiY8U5GldU0tcezH8VrLdhtRCeqpLvTWmHajx8zs38Z2uqBSnX31qhtWj0ew
MOihddyUvQVcY4gy0mYyVODeSK3nOaFwPyvG9rMDQTThxIF/6AGiQKbag/HLQFgz
I54z5j8oMBv/QR6H6LgJCm0bSesGn4whEtLbhDx5vpBq8IvmkGs2mMoTNwa5IeQD
wbrUsjKpI3EcAL4h5wPxIVQOVttQdN9NzDu1xwhQ1wwTtMgBrVQ3WccpoHimP7ll
LPCquqma469eLSAdxmeatyDG4pAV4JbfuWeI4pmMIFsEwrxwWapPM4Im37jb4xd2
SVv4VUnqpvphDsS+BaRb6zoAtg4OXcWEHEkFfUmkJwuYSSJdGQMnCb4VaKZb+wx/
OBzCJtqf+YCdkrxys1ioA3s7Hl97TcmmwD1ecwKsmSfaUH7khC6fRLb4JSiYj+e9
8hMUuQrptMqwEj0vMfaweXhCSAqNQu1iyVB+bpKSHW7P6cCy0m4LOS28cUqrV8yy
U2RauTkfLAj23RJdDW+SM4gGWE9rvALJHzTIHcaStqTC0r8lMAPEm1wd7S6/2YHw
eHMffp0kBqLcNQNES3jRfkisoeddH0HOKv8+4nBWgijSRmZV+LJ8JYWBct5LbbUA
zYhJHxWeD2di+FkF7uZo7agu9lbgjGKwPN7OwWTFOajzB5cqaqWeCqtBMZI6dOuf
T4TxEtS2MccDyFyfozsto5vOD3WyoG7D9B9Hgv/X5je2tV66oWlBGfL2Oi7yzVYJ
vHS4QGuJ0nVWfglTcnn4aFV8KoPIyRCY1vd2E2jIwgBi2kI8omWYyes8GVRsDnUa
qAl+FvYt8OjI1Emadb25ooG1bmiq0m24zJLvqYB/vFU2b8W1Lsk2Q8uN7Dq904MG
`protect end_protected