`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 22016 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRpv2xRODiJMNLGiSdcH6P4QhuDRbVm+q8/H6fw52YOaN
Lm5QfnT4GNzUn0LF+8OS9XEiaZxa3ti/7GB0G0D6gwSMGaV00+FHbeznhqJR0n78
G1hZAh4aaiQ3WupFCMaCOJHDLUrxTZJqLQDjuau0019lGLK3FE6OZPF9VQG2u9fh
XDEi5Up6SJr287yKvJ2WHC0WBoDcqUmKcBoRmwxGRU8/JioGkZOgooIxD7zCo/TS
I+QtzBToFqEk7UdK5QaSeoIJyzuHDyTH5FcbwgZjIrfUPNAg2IWR8yVeXH5AEZU8
Nfaa4if4oSVR6K1OvyU/cKwklDMg8RRxKZAUud4589JXayF0GJyxKDl2rKOgiY+I
f/GVPH1Mn3VMRgUJCxutTI5gjVUiZhdPC/OS/WEmA0Qla87G7TAsvxYVzQbEKJvI
DoTMkYpjPfNe2cm+039Qkpu9mTb22CHKdappsV5EQ2BfytHoNIFOdDB7Oa1O4s7+
8Ck4jyJxwtjPNlABSkybiJ982+PYIGH2Zt+VCAT5bSK1Qh8uhixw4jYATwlC2Qpu
Ebi1yM2th6XuPOgrlIt9c9zWaGctOM9CW4JGZPMloi8ltUMrS0qcaFFCYv6ic/Bh
knY9TajuUQduoRpyh7r3TWEicDvAYvjPnOnwF0Mr6U1lw6VK4t2UU+XmeFabtavi
wZDnwglVLkFzDGlJrfPUZM8PsTP+QKKCzKWgBXwLuLfel+EA9ldo50lcUZljZwG/
JCyTaKcwNSwqhNP6jfAxB41JE44A97ZaGHS0P55ckIN5gZvS1ywcZO8Ev06Bz4qy
rz9DV+B0HnKTLKQ3pypNHtL1cBJ7fatbum0qi1xIt8Y3EOhT91CUtYNQF+d2RITi
t9x6eCPW79dWdr2qJ8PfUwLlNf0lMqqY0TnHFBCsekUdg2SAXghn/9CB+Ro5x7QA
+ynnfexDTvB5HXEzRamk96tei5Yxr6kJEUwrCjdXKBAnUuCIvuhFtxlIG9IW7zKU
LkVQsQ0ZHubZtxERx6WGgjKcZ6zytO0l7jFVDO5F6l4rGGFnuIr9Go649sQoUNLx
Ew5/8WYo0rR9+bmYLRJNYqtBNuypfTlmQwqzVaXvYukDKPaYBzTc2Ap2MZLYlW1g
/ecqxowRVSZvh6sRtyIlMEe/3/xD+nEQseTHICx2bc/M+skiCpaZRkMPiZqHEfeZ
GQZWwNqUlC0vjj6OApji0m0Yd0/lwAO8w0ukH4I4l6S/CMS8f7Id9VwrxivtHJRo
mxWVy2JABWplyUUeppzjVT6Te1KEBsA/HSdAXYLQgeqK++ZRRlgoC7bstNIU+0wT
GY+F0YvhsmNohy3jO5Yxa0gssOEFDoddiGKObThcd93lDYmdPXhRwtn0/zkZpoxJ
q4+jJ5lT/nm/ntAjsG9/IcyXMRPu+QEIAGuX/vEdoXygmK4fQXDzL/fB5YtRkCsF
8zEU8yo49etKjLe6Vovj9F+kfzPbvSc5MMgTHAKIq0TaRSb9Bn4zCHe2u8YBYU1y
prTV+1SN2fcy/q7ek1PrCO863FiCUfAnHPbhMBIe6ieaE6etKr8Q4506KcUk+F3V
l0hlbETZnq3FDySb934LsSnw7asaQCnOyWccCUk4z/Q7uhdQRPVbA9SRcs2EZb8Z
oFK9amFEiAJnkK0O8+8OeDbYE7e5ct+yHya+7JFMzXOrw4F6Va7LR9PYgbrTjUjK
wgOkJZCVNmnn+xzPw1YR1x9IiX2w4TCtxMU3hXNerqirvDrZY/3Mn+10amYkj7Ob
Tg5v132Ud7jK3lobSAZG1oxmfJTAuwE+fmaFIzRH0sYwM1dCkaZaVBa/XRAx0sGa
dtUoCtBWwp+qswwgqSCgXDpWFS9Cq+l5sR5fpXAzFuI4PGQ4nBrlRiCNHofnuG4U
zKlXkAEa42hH1ZHBWq4q+GRvI9RhBOVWHfjOXWU4+UkqdkzforFxlszCeWGAqbkg
Gd/FzbsMfm+mOxIrQelTQ7HDEd/gk4OQtLd1ODGCreYkyvzjEMb0WOfZI4LUUD+J
iof0PxwcGf1AoyMom6S1yGUUB58NVZ10oQVjRgXhMdlbCGhYuzSXr6CJowcGNyo5
GIaS+B7XzljiFFtWyIIrQNxUVI3Pu1Ok3C36uZuMhfsGftFuGgL5q2VEHFnZzHK1
R1nJWeaVfn+LH0j+33hX/xmMvnx5tSk5DJgkqT93sYlkRKSUgNC5zPVxsVY81SnO
q0tdmq7J5SXvyXPjAUmi8ig2/19Ec8Sr48ToBjgGU5U5Mq7HyqLPC2jxQmnuXNR9
GVSliZ3K+4C2cqHx1iJUAduwsjyCSKhXCkP+gzAdGkcqU6IHwCKV8Iu+RdV7OYgp
wokv6aeX+gCUDnEQj+Kno9L/Y/gxdbgu6PNQ23OdvL2IgnlrYVoZkReVbYzSPk2q
PoyisGRULRjQKzB06ZhAvl0aO8V5bfq3oi96G7/re/fJm4jdfG/Mkr3+89XOBD2D
uYnA6+XTD4mO6b9Zsx6ZdzkD3C2DTJmYkmciZ6cW09412YDQd4QOjlOEquAUsfKX
ZuEQ4NkF/xZHC1rsDsCibqEt/U7rq3JPz0L/rufTscPili8dDpqxcfD2ynniNPXJ
MaDdOVLHYK3jXOA3HY0evalaLTgGcItYfo6RkqfqhaxN/yVm/ROmkGDnrORJPcgM
JOzMk4X+0ONlUUh0Sd8uI7BoMnX9j/+EuUWBRr++scrsImhXwpv3FwYYMZnWS6t+
5S1Ywxylbdy8MIvWrzZX08Isqd4biv5EFcNLFbblc1xilWdtRf8lp74b06Wda8q1
ZTJq2Y/Acl2xSZICmYn/47m0NxKk/UPZgMQa5dbohXfKYj9rm/amY5YYjgYDbWU8
DqlC83Yx1l9fzxZku/v1MNoK01HNtuLwqp0wd0hGPYuykGFo7mHm+En1QBXYrdkk
zhOAKeNnaKqFtY1i9Ua2z6HBMol0+xyqYhCeVW6QcyjqeFRRBet3ZSK/Ma603u+U
fipfgAz2AFFp7LSfRX6PQRvVlhZO1rHDR+4MAeSpNZ2c5y/3XbqzEmGrNgC1yUrH
A9DbEl3XFTtbGs4vp9byucRe6clcmlUUf0iNSsob31apU8CPjO+i1FLHfWmyUQQD
tN0VpexA39pGlW8aUNe+EzL0OF6orAgVmxOboaKrRapKmFY+uvwolSI5awiWf/NU
NYJpAd2BPuqNV5egqC4Th+UOudMtxPvK2OgofhcMposmH/ArTFLovZQ5sDVTVBFs
OtLIFJv1reo7n78nb4Ojx3ZB33Pkj43c3eYUmB1+iAnnXipiLo4MLk4cshRjYc09
Yxz0Ex2jw89V/jlfPoD3MYyQ90C0fHKFaTAjegJ4pte0uGZmxtmUS5wXEUrWJ7ap
WY37oOGTXxgRH09eNFB8KCB4qPXtajyn4AhCwBbfA6Tlg2hnRej5dowMuFSRkqej
5jL8daSfFgSjDk0EuuKhzhsQiuA7/WBLXAzHThrubx4K2GrM0tmqT6rjoIEayyKC
Ln8Ek1IAnzT4+rVTDMLfJdZR695a3i9k7HtKOnaSx+gyDXyayeOc5y1ZexHPypXR
mCWvfLKw+Uixcw8l09uMTdaqx67sXiWcDvKcBu2lT0SHfNLWdie5nllmoLvVq2JS
dGloTd02WrL8plTwxhhCOp7zQOw3W0xJ1WbxBBkgbDi3KfwrgR+DNZphe/w2KqHY
pCR/iIF/yoNKrs/mP4dq7XVEFxwBBFuF12/3fle5KDXvIkvnhQGu1XRfIn0Y2W//
QPBwWOQw6AfwnZkX5PKpIcVWS+eTKFONNKse3XJpOth7Xz20TCNfFUF9MCQgIXvk
WVDbSbZTAHCuuVAU9Fy0HQ83mlkGJC5RlzAzVsdHv72vUZw/rD5MzGv1OBesJI4j
rRdXUkBboeB9Yl8aq4u7c+X8qD+FG96NiJt+CBKdqFOxt5v3CKwyFvrNC/8dlW8O
ymM/xUIry+PM/lEFPG8eEllADh+Izn24uvXwu4dTQEGUs9aIA4FU7KJLYGU6ZDD4
3OOpAV19A+St/kDl3qiHGiVR9X3PBjgrpD54s36hU9FxZUsC5eV17v2m5TYRrYtb
TYpYwd1LGVDX+ZsZ9T293fLGhY24m6WBToLZgwPWhD0tfdjG+DA1ZJUvOfrTeuTe
Qe9tqCkt5WDfs24VA7P3MNKSnMOCleyVmBYJ5HPbHCDqAvS1m/DTCzZwWyPgoENW
6seahkwDtUJE1iQhNfgdA0lVUHV8TRs3fYD/y3t6+N5Ip93K5ORnjUXoQcHaPzFZ
elO7aHmnnU/TUqTmuKoUNfq9o87wSWl/bTDhr+7B3sUwyX1IX5zvTYyXWbjP4YXr
tnkiM9VD9vOQu3TLKg5FVYh/h4M7kYGGFJto9MunQLgpgCEZWMk3jaIQfl/w1Xcu
t+nRR0+NnDS1qI4R+XGsHyZls/AHNYWouRWy2FpVBzBcDEJlyYBE/jq0xzofK/rK
ircTOFNnJU237WNakTHX3zssa0lvxgX9pUqzX9DJJuA/OXLg0R4h84L3JkuOY4y/
0vx4Re5nbkOjto9ZylSiJaKi32zEwVW875GXje7u12lui/71OGH6WEQfZvWsvgub
hT+LaDzz1Uvdkj50+s8XdI5tV6ILAo0BjTR7NBfiORkLkdvFmvlfKV9rU2kV65oH
dhupcAU6B2IY5yvqq8mgR6X98qvuEkkQ9L+6wrfI1qi5g/k7xFPjm1Hxt2un1GNb
VI9C8G7Wyv3V3xhgJDxH7k6rkzp0/cEgDhqOY3yagJZblYr1pKKe5XyBzFYEhmwp
FYaqSp4a2PodRX3sK+7+3u09WQTrmrOQUlFLshc/vAO+HTHxuGVzM3wShR3xS6op
JRraEdQRdhr+fs15wHOI7YuGexhPEcvbAnQNrqK1yOGEdyzK8ZUQ/uTBnJxbu1LG
6Q5dbvSRist3E0x+KCXCnKQJdOS7keLg6E8Mk1GewAjTuHrzsuFB9bYaqFTW8B10
HakXhYYb+w++5RIx5Gwaw47Ix06Jjh3tEe8Lrc34VLEnczVkLCADDMTjZyi/ycpC
H0rTOleBzq9TEfoY3InA9W8vUS74E//wf6x0uMCQPtHjcYdHvKhhRYRiAKyUIKGB
H35qt/eY9ieGjWG7ZkJFc+xcIyS3sInOF5D5W+K07bBS2AxYhL3vtFGZC4KL71PL
qwTjZYxTiNT6GqTVaV4CQO/Lq83eFbIYkZ5cgnN6TJgjtgRnudbNmCaPZbnh8Bdk
nlVJIDOZJsHXCnwrZuWcoukR48fd9wUOmN/T9jjLYQ62i3x1TSotac23M4OKKJBR
ybh8aZVleUBzwq7s40jwbuwpCwcLpuGXmL60CoiX+UYRxlD5GsXdNKJBdWrzfKnk
MTUETa/CJ+Uc54EtQ1S970n8dt6zDl8Amu5Nr7N361ZVEKgJLOmg9UF6ec39zMxh
uPQeOeLu2ALrrghIdXkqPK3Q7n9xRvjsfeJZMpEsSdsK4xcuiv6zwUEmMvip0UCW
BjxAL1dFeyH2Q7JAiWSmfUSffLBiKrT+qd6iId8bjIAqUYq4TG/YdCD3RjaJMvDt
p3deQMfr7Pqh7Zia8G8fRIxB5QCVkVOS1t3J35g/E055AQmvOwkTp7BAcpS8R8qt
RbEJX/QDCNAsdSnoyriVKMLcqqH4Z4kKa20ENEQbcuiWya5OdWE86Rxag+rK7B2C
RKb74QxizWPqoQGxyloOyiJ2jSarfJ+VlgAKRqTShwTpwIlOTieb2f7j9neSamiF
u2q3uax3VF73PG2lwpsAAeEEYh7AHs8g4sqPLfMRQBZTg/6ki53d92bo64oG/Qyt
CX2CUa/mnwenZGPqYqxqf58XDWmxsNdTjxbL0rwuThyckf1v/Xm30PnJDyD5cG3g
9RkbZoztIyOuFvGxYI61cnBwd41PvQUxFkYOR2sUzu7EI3ELN5JZGp+u/veQAYXN
ujMMUxQr6tkJacdUHE7vbS1Rg1pLw4I7Xd4AMk26fTaEJY32auxy58m7cOp0ZV3i
1+WsSmUAyTYouNdgzRyDTppPaaotgzoZbd3zeiILK6xTAuLFr+sBGZKv8J4KTq/X
NIr5PuWqzXulnE6VqUTjMEUZThrcSWLNSThkEurkXE2GAATFXNtAcUHyRyVuHS/8
5SPpODMGsVOOEGBgn19eRL3KYfhkM2gnpgPAW4+6uaXwyvwL0W7ThHU4i/UmRNIC
UOH2Q37KNdv3D7a07ogG2J+cO4YLZJCsz9HWO5WhjFXUDFUb7IPYHNcKliIc6vSY
AuyF4569g5gycn1Q3KFBTI0IwwGD+80gUKoGbtmBPAu5bAr2gLNGALsEv3HDLBEH
x6OSeAbMPa3GZmG4bbUhW16bGqO7KJ/jn5eGpOvDJvrBYeEe8V8n/a4Gq3gAluW+
eXQZp6iu+qEQbjTwkEtNZZIoKnDp0lMu3rXyHRBdJs3iBGebRlEACu9mQtOumhoY
1OuGsXwTWYbjkUcvVfG+HgIhFlTWiYlV/5/1fRwtTUT5/p0+kuWBI1MA/E5tUjsT
iBtxZBznmRb+B8y1L9nsBWO5tin1fzK/R0jBMTQxtqkbO6d/qa1PezQKdwTCxiq7
nOAK2MHrhgE+Cm6dgGqVeuf83tJqngUtaPSw7WtJgi7Zfx4/u73Kd0TmASg0VgEG
vKBlsvsCIFGy60ccKxBUk+8F9N0rrNmM6zk8RRIcDT8A3oGpauQCmEFIdZ2MdasL
35w/duLvP1PBle08sJIcOwqQDecQAsd8kN1qzXFY0oIFKmWUihtddYPeksU3hL1E
aVS4sTFeXWpl6C69ZO8WbxfmsGZ8exMw/IMiw/PazVrvxRiQdsSJqgSQ3OrRhvjo
mZkyvhK/8sss28KuXxvMN5ImQcF5pWexOmSz1oRXZuxvOQBLBRDP+hcrlFekbRVT
dK8cGXIF1e0BOPXt/2eLL67cO6O4/rvQ/uh5rHYGANZx2vUhtl1Dme5rmb87jxwh
fjrIJTDXlNI1zXKx8/uVK/jz6WX3TRDLMx4bzPniu4b6AzB01A/GFQtI48uOImOL
ZuWeSiskZLGGU/4dzMSnaaGep8rraDSZ4YLFnS9a+yHeYr+Fzq83U9diFq8zP6Aq
Ouj7Z5MK3PvFxdOsV53hh7YwDua5orJP94iddVumgGcq2efy3/HiXPQpE40sWzKj
VkrFZEg1O+iyklrRWudCS/GUAEWs7gcMf5T3Hnfbwl0dbLCkCHNJU4UyQvLQbVa8
qMAPHW3/rSSs+i8EWxMYnDjhwP98TX/e2BuDTs20oSVRcDucb0zbnLzr3F06kfq8
RNM8/G1R/Lg7CeycyKX7dPnpqsqwX9qEYa/pbhf0hrFzUT8oc0Ao1u/GU8IDcitE
PlqISfBGJXUYjF0L2SunRfCR+oRWx5Q+KdC6Bwb1sBSF5I4UCAGoMAB3Q4koQDxe
WBNx8dTGD0FfATWl7IHlVz4wsPcP9WX+6d6uuCTixT543xq35pTM7sMAZUtqeu2x
2qZSoYuyrh87KoOQfNP6hiEN1YajyrvblZjJFMr7oNm0pnySL5UTwxBNkqLSsalH
oIGFqievD9WUupOCPT9/WzixQ3uy0N1EyCWyWxt8Lhti2VhUrRabbvRUFsXkGOeK
1VbWXmwHohn8+kIjbkluTYVH4CUz/jvj7/NYBHwVRtfx+1pgJaXibNGJ2vWW2xar
A8dLE6ujlCTZHyc1dGH9xknI4xLchtaHs/gXJJSBgVZU7F5l+qmPPMrmLvyMsZox
6FK8X9ryfgGtyagsQfdQD8N/nwIF1mlw0ihPop9N942SBzE3xx1CbpdmpF79F3dc
gYnHfo7cOUEztD/KMdJVu8iIaIj/GqnMzGoIn3JmdugIMyoBB1kqeGi57Yrg/Vy3
3BrEIp/8UM+MUyhW3L2uJz3nsn/Neev08JSSpHQBfYNc7Dw7wtxReKGzZZePLIns
EG2vcw/SvBjNd/63ZCJM6TkqLRlB2De8la3IyHktGy1AOVmGy8MSYMpwgTsMX2OF
WBCavV71quuanjD9ovkeF4hg2hoaE7nVo1lwiAZrqvey1lhB77ohNwkHcz9CAQ1m
Ytrc9psIauhmUG1POSGv4/6b7t4jt2k0dyQ+mi34DZ6GlqdYcF+Zsn+Pg3IC52hW
ukC/5rZpK5L45ARCFs/e3q0UpMDFbhlaIftyvzj1w8tkUaRYJIC4PpLZYIHmh8Mf
5aTofBa7c0/TpMm2n7ZmksGNSPFJz2P7fO0SXg477gjWbZNymEOdpU8vhLqLOof2
vjoudGaOHUzO8tJS+giOxbpFUgDjWFgvU6iqNypIiI3PpwX1sq4gyJlKYfdxyTta
v9HhNO+uLLpbflEYjraB/Bnz9qB/tYFQSY2rsbPytwQL/5N4RdSCia/eBzObD0+p
VIGTgnE3JuBwmBnGxugBu9GaeO+vcrxx4r/BTKMZ39hO3wGDVnidLvFJN9O/Qa5g
iOqLi315mikSQku3GUhVfDMjzJO22OrcVxs+tp6AX+cP5LppjCNCCbGWnNv4plTH
xgu4qBl3pFr4MB8RQGdhNM/kP2wI0dpbrJrt85jGXmR1qocZtSYY1EHubfqPs1WJ
uwNhVtIHBMFgjW2mpJonPe4lYWCe/c06i2mB0PiPe8WL47AdblcIswIIFETFQRCv
cbvzbxJwJitUqVtG0DY0IpOIxRMBfbhpaEvRwyJFh2NQAyd+R8DiTxwDi/cAnK+4
4GYmBN303Y6nufV0wKfKw/rIijgZJAEkCRgiVefDG3c9wu+EmAR6v40WB8KjW7mb
iYH5Vwb5sxl7nrwJsxc19mdpNhDWrcEDhNatlTwzpp2WHCSKVXyEzTHLYFZtF4x4
OFVRCkb46cRHtw1O+mGWIUyLAlTWC2weW8r35Hikm+vHQmiKD8loD7dzyBHvCmfW
rsveEWwivybXIPekbM8mCXho/++nIvqKQnQQbodOtGb0P3pzGqlYw/pB7LGD44XB
A5RXikh/rp2JzAkjRWzAPWvTskVhKgmJtnZ98YwxZlg3CnQaG26JFMWbfAG3VFav
ez8tCvhZiqilWGJI6D8CxQOiVeJX53VlAx/gw0G7BALz6i4CrDiqIQcofWgahgDZ
OV2GOz4CwExvkb1lbu3L05WNI6nCHZxFlvHXjr97doldzihqxZCHOrmzvhfgg0Cc
9eKlKoJ1On/bqurI/lUJeG40JGOQtmCuh4Z6lZ9dw9SXzwHDfnw/+oDg7BQRmgx0
eHsQ3ydJWXv0SyMf+x+nBHa+PK56xZ6L7eysJe5nSNBN8+1GGAZPXsnnOBzlIdmK
8cnRzz7BsdJU6fpkqVjAmhxLVEJmm8GNQqg2oAfE4HxOqzlTQS3PmfXhxRdMPC6W
tjBupjVpqnZHsvk5l9yQUAZNKR3HMSsvlcskbVpPkG4+iCUXMSYjuOgeH7TiyA2W
ro0Vt0TA5ujYT8gRgjM9RIV6LhrfqNx9cHcTkB+pAm+HGafkE+Zn27vp1WmUoasN
MthGqoA8kf52cWcreqH9HRBRXKfKenxpHXqe2MDu4nxgzi+4do4vkwLB8SrcDlJs
0v9btpk4xPAGu/qo7O+6auSM0yKHlL1yvkpgFpG+/z9EL2WwzWMLjEcWnGYfwAat
iOijtC8YHnOeJNeZG49BTwnjvcu5aJkwl6mh68ap5vYs/oMPRNBIdSMStxa3KDDP
PsYkipwENPyuVMSFM3MxO4zHxLAUaQPMRCfohPJuu5nCr/UlfkTtUqEGR/Ghw0w0
bboRWI1sq1zOSncjJyclpAA+rSM88OefCAIyiOIfaqaQV7NpPiXhXZknSu/WgYOU
Aw5OaD3rcfSXF59uaxLv6HtIgYiYEqna1KsKNrwRnyFk+FzgFyINR0hxjWkx100a
3GXD7dyqqNd3OLeFXZm00fnWe9NT6Xo44eHNuwySDRy1RKAv6WSDSyc3+uUrYg7p
EUd2vBDK801lcxLuH/ix30ck5i9Q+iUzsZ6jWL9L7Dg2TJa75BuN6PWEGR8Y/Sgx
Ep4Rg+MI0MOf2sJ96F8RKFhTlUYE1uJe48A4LaMJwc9CGd50jam+frDimerQ1vfs
BSGs8xGpqSa2GwDsCazhkg6N5yfJAoPuaGFMecHWz28wxBNM5Cvlkj1O+ts2KNKV
cQ5bLsYLHjwIcgK0cgR9FyQmuW1hVqX9h5Ca8QzCTm/i/wx+32WiQa9C1zQcHSrM
wabSQWPGNMZv6FGYzymAOASYo9WtD/Uu0bgbN4GWwY+SjSL0MqeOsbiGpDDPlXMk
VSIuSP3WwU2T54H4JyHY/adHy71241KHTa8iE2Xjvb2BQsRBJf5jktG8FrGFhgGD
CXrbxNhYDM36vUFM9szNcEbo0a9Qaj4TKL0VuPDTXgNNFPKdGjlO/lkaB13yEjXC
c28/eJ96EgqYeVVnbfXKr5lBGIaqZnRGULkrXJThQSf7YPd/9TP6vfJVL+v3BpG0
JKk212E3km6T86as0LnDMsxnvZwCwCcXW68NoSLfylHWm9BYJjlkicQ6ghA4SKBa
l47iZUJB7TMY0paE4ev96KCWmZzMqdkU0yAbbhy80lfeP+4yAWOwyfBDW+fh3qjM
SZa6S6/yjuYtZtkLfeOd7eViuBJX2mkdaNhAih66ahZuWX5kII7EcX5Mm3fTUX5k
5gSioErUHUO7GGDCLKjzQmRsvrYjkzb0TdIF3nGuLDK3ho789I6NsSjTOI2HqnmK
o7ZFSPOPTR0MDiDOyW4OjN2JjT9XjcEVrrOit38O+nZYYp+FFT34iTFvYX7Mhx0a
YU78LdGtDXyBGpAjvbHRFfr+DPVGFaGRJomM9gcdpcZV4Ha/toMTN5uga4bR022z
UFH5kDhNs/wk/T8uQdvPri1rOoIHpMpn2f2VL3KioM1nZKQpna9P4JTscKI0VH8i
QdGUY4KuV+jRdzaf38B1ztdomb7LIC6s1QEc+Rn8Q7eyfpN3CUfCZyMO/AyCHurO
gYEBCLF6cGoyuCk0eftZZQ+xgE7fKhSSi0cSpUdu1Eh6P2MxW2IxuOcXeBCwhERK
MRWJQAA9shuXIDRG1xUxVlXh9Ayn3H/A2oHL7Wwn9EaO1Gk/WZEmuQoT6uT2c3+j
e/K9SaUzFhR1Wb1kEQEAczGrlyAY2uJm5Edhu+KBBgh4oll4MYq+jZd/aXjJB8BW
qkr/qhlr7ph7+uHTk/46v/JJO9U9CCvycvCyF0nVK20m3nPf6cxnHW/+fpo6l9m4
GnEzawI1QuioCY+QsQ0heSL6ZhQMXlIKn94yZ8pBWczRTxQSh+jaxBMTGs3YxqAz
+lYEimGIoU/H8SGgMXTZ1kHHb1JBiczCTxuqbm3Fbwy8Cxy8AI9Mf66avt5uer6D
AZusDL/ttNKadp8gVty6uKwnMsZPnHaU+wXH2+7qTrXKMyi9QD56kOX9dnaX0F7o
cAmGpuRWtfwLk/hN4zEh/aBXYHMii3nBxvmoaP9+Nui+WMC1RZ3GJkgLI7hQQnCQ
HGS2Nkin+GaJcz/rjBNG3Kaf+8p+CmbvnNgFc+69jgO68KQGgRAXsBZVxI58ZyHA
8+pck6iubclqA0/SYqL0AzShu+oxg+nhL18frCd6a62IyW+cW5Un0Ql79k4Wepv9
pZge0GO9NkfqSmdSkJ9TyvYIxRibgBrYMXe+MpUf+aSmezhsT+PxTBVBP7Vifi/t
KTVEZnXC2PCsWmgEvjX8E13ECHNu/weG7hY2bzRJ3p9JIDUE0PNNX72qH1dRkUAw
9LmDxJlrrMCbOYp8Jqs7OTOJvYb0birtZJkfhJetAmiuMRdf7BkbDtP8suBsQ0k0
gNiUBYlc27kEWDsWGFP0n+Faq8OSOrDm1dQRkbySRTU6wNR8IvRepNDIriR7pPYp
ogJglinhAKTiNPjgG6EaYf+sMz2CDCY4Gy5UhxonFpn7SRYO4JWIHpQd/8cCjOVt
WjSjKv90P1AlqfheyVvxHfi1RF4bL+N/zpqfsuC1rG51W5Y4TiCMA4vvum1dFY3u
G4IG4XORna0rhp3arlz4c/vXuFahAVUQ4uj25y08b56uzjNlcAYMDhVXNsFkPPnp
1WxT1s1196F7lMEcrzALGFqARTCfzBIZ24MtyrJgX/U/ZB4t1spVCt4c+B4Blq9u
IdSmPPza7efyL+djHL9NFZtVmTpCVhpiZHqWGaxOSpcHAVGchlkLnYM8B48dPfxD
Ox5QlJtvVjTBc5PuTdyQWel0WS5AYo2W4cu3hvPUyjol5xsHiPJx4TIzYOUg3oAW
Hpb6ePUJ9Nt9GEqKhY3iua5ABWFCdv56A5jcnGcAyKRS7vXGkOnhrtfMSy8es/BA
sYdlEZBbvhVKUcAi5PV3OZvpnF+49yvUC6P63fosD8/iR8DNPH8bpxwhOK2KxucW
sANYDgk2nHDIIjbDJ7Lyg1D39m0/RCeeVzGokv8KzzcSsBHPP8qd8U24tOYl6zuo
eQHj02sVulYZjr7C40rSyIm0WmKGiB2k9NsRYTi6/WAgKdmSca/YP4jtlTN1ALKj
Ad7YL3RB/VcPNq2DbvUJHUZ1ZO5OuCrebk3KlSgchT9hcAIVsji/ULff/8QAGVB7
g67mNEglqCsD1wv0NpQvOMJFQttU+kCwvPK3Ci+J7FPW+Gwdh7+wBo0TsYiQjwIM
eXE9xVhNOQqRPRMAeN8HEu7dWRAKWT1EtWy6jKRP3ndp7vME9AgTQ8NwLNyVeA3I
Gt62I+TFl8QD9hhmHmZFAOiARyeXNYwsEdz+HoeCq1GzjpO2Y3ckPFWDdg6h+5wS
kO2rhDUatylsI9dQkrQFJFFd/Hmy/Dk4KBrscqodgXSVdpSMgpoV7tRrTrukTvqP
6S8fVQ9Uvg6cWnvWyOFiqhFoGOeRHo/o2OPCTJ3T0HK5JQoen12PouWSpiJVLXMp
6QkGTUrFhObcx+fMvVFyUdSvT6UOzWnAWbyd6OnF5SKHKiivlmXJ4RVzMGblMSH7
FjxQeUn1jLmtOwkhBDWJPKoWce0RmrTXZy/K8YoAC0FezJEVvEAel6vWs/n0M3lC
2Z0kXUrttk8UhL0DMUHoLVOjcjz4FH5ftbv7iqQzsVDp7yix5QIIO7mJ5XbsDLPD
PRrkrS+tA3BIs3D/5rN4BjrGDuJuBSCHvzxFUEzjCpPidVWjOSrPnmCy6TmGqiNl
teErIhm6lFKQDTtx7AyvIMOmy7YtDVrVC3wXAproi6FMvKrzgpkqyNsel++c41a2
uVBnKI0lOhQemTdKDzFDfATlGYqkDRzM1eG/GpxU6ORdCrzjoiWXFxh5FP/D3OMU
HbJRWum3W4gEiZrD91QKwI0fPOuqGze22V77//8NQjJS6o9vKsxoz47oHUzbUkNb
fOWdRnuAXG6IlPeDUpaBRs854uXxfx4A6hhFCH1uUUsvK7FGgi0emXFaD8ICNEyQ
7EraXAnsVbUUETxiobmxnzVLmMc7XGGslXg/Rouz8tQ4zTvjsRXFQiPFCCSAsRTz
AK6HgtUyBBfiAQzYy2r8gzjkyyLZJShsAoCBwBRZCqhAnuNB8R34DWQgqRPmkW6T
XIHZKQj1iiXFPtyNfDoF1KzR8Qy5i53mD+7QwsAVD+MHTYma1DzEaKWZ3stOpb/t
P1J6JkzeqZUdoWW3RrUML2+8SGi6V232g3X5iiQnWc+FcOT71ateKPqyKFd9lMGd
8LUIrKyxse5ImS2ARsdE0MmEnMALmzRSxCmR7HvPTKOqrjXZLTgXthkhpGngdCV9
P0fy/pD13b31lF3T+/0OezuJuNG8w/jIkALL95ogGDPfWtHPES7NrP/5udu2GMR4
rvM3/kr6X3DMQKElmb+AI+eHapNPj6kg/yZcX49V8VQMkFPhK/z0bVJu66sdeaR+
Guhw37WKWvkilksq1VCdO35Au0UScsI8Om6DLg5oyJ9WVxTYPg1BJk1ULDZcNpe+
Hb8e0gLbHAeZXJh8BkitLdeGTv0QG7krvEb2nQaU7e8uSz/Clad5vVAo1bGeYpNO
ezrZAY1AUAIS6mj09Lj+RLoGYPcDEYVMzMoZjYfqcVrKNXOKvjEppKjBZ5B7951n
wbtyJNETOS16DIVDzXWhpjk75Rhcy/N/cLibm6JziEAAkMBelqwxcV+CHuxZVB45
pSvWWrmEr/qUsFkTCk65Hl4x9PLq6YohqE3hTyJY6VJ2qIcoax7TnfdIw08YpW1G
oAt/P44tyxKqdpEmV7nbkIrYXh6ymJPNG+7eKwhYpltKYkT17zb90x9EDmvcinaI
swFq7OdobnQ0bRbaHQCgkzI0R8YctL+r2A/LK7ipwMfHki7VkcAFec6TZlvt+COE
m3T44hPGUPO4zJ1ghy8q0HPX7ehLsYIAsJMReTrAa3uQEIamEmJM6boWbA2ioZCP
Rfn5InpWD4OFcnV9cgUBja2NLEzh0zzT0datL7F4tARVTgLK8jcAbfLPc87ISReQ
Cdj4sdarKYbTZYZxhGH141RnVXIjHuju6UeNYt3u3JZVlhtTL38o9XoWn81NMtd2
sa43nD3YGzuaio7rr8tf6KAdly78el/Ilxr8WDfoAFw/zJGjDJeQsoa35ozsQOSJ
da9NidXwVQmJELlRdSffVAhbnRRera1c/UKvMgA0ORIPVHYB6mH78pFqL7Sa2xpu
zHyp5UUHT0oH9B2pl8VdBPyNxc9/Fh7dNdqwxIgMVVg+e5GK76eYlBCvva/HOo4q
8M4QxetvUpsH/UoQn1qQ9MM+0hc0FxcmPWZNNgjabY8g6AgvP/QtCXMgik61MsvO
9OT/8ySWkOJO2aLKQZnEt5aE7DBa72xrcNKFEFGAxpSO9EZKSE5qeib9B48i8ZHk
hOqbiWuxGbvd9bgzVndzZo28i54VxWvtD0Py1ad3EoftPm+2AmVQ72EketB9IKmh
J7jqAe47lrttHVOB+w39U/PTj8E+IKCxEUPkKcrUReQofTb44clX5qRHZFrT4420
21lz0JS10hFjyZmBMc4wjwY2Q3sTwImSBp3gE2m0AFTGSy0nOdJtF3SMdOrkCbTc
h+7sWxeXhr25hARlXgIfdZ4sQFh4FlX2MuPLkj2vxq1UHhZY/LV4204N4E7iwCKh
vrqGNTsoYKL0mF6lCDnJUzx7GiOJfPY4pPiWEA+0TTaQ4UJB8mavs19jefv3ZYR7
FwEUD3DoxogDNgkkgR4AgcshVQXGQR0EvDxSMWpGtZTIOZiWovSW20+lIwchxdzn
0OVfoNF5F4/Z/xBLaQe0aMyzBx14NqwBdXfvzOfu72ffbkBolNKDePXxoXENxP2c
3W1DqQR1xTLjLlatrSw44gqua27+qa2B+o4yF0a6V8z0RxKYnygNDelekICNbphH
erJyIrAbTYo36ZfP4wF7OsuqT2ypERuFlCvdZHDqSImwDKzwQioyDeitbhz825J6
x8fBbXSgDRcX418k87F612Jk+z0w5rZMS1JAvf2d4veis9qZdCPR4HWNvxaq0Jef
ZBOROJs49Og4KlgNL7psS+sZDV3QTLsAW32Rjce0iugYpe0zZvo/gQoUU7qZBvn5
A3XtS8iuwZfbmz1/+5FOMM5qlWkGhus1kAnYqFA5LGjl55sHo4gBULu04TQ0499J
+5lvKAfl1hwcZedvrB5ZZHwda/WPZ5ZdUDxYvoNVNPJAyFoKmnztnZLYo0vWhcqa
6YpJG9nzKAJ3NOdM0x3bY11RYQ0243ftCjh6Z6A6hnmxxqdszMGA0pLu4qwKQ/6G
IAlMUqc4yFaIGzOG0PNngumUtvUJYJtIZ6QJbK88XelyTeS4sBR5CmC2M+VPXR+w
pJ0kuA4oR84+DX6ZI8T3MW44fdS0aGXKTJQ5NqfpnQsMbQOoDI1RMYGsttq3fJfZ
pu/cXjdqTUL/Qj5L8vhlKldnhf91PqEEAB9gLr/vLYjTYnn2MFhXZrjsiQmCRUqG
df3NFAn+ms6rC8J/ZQjtgLdGqDFVzD8V9KmJ2xLGe7259XwHCLC0xibEgQ4CZLkl
K1kCVRTB7yl1KR7uh7o4FweSd3+CWTB51bT5WTvKYjDQsb4PLAIaLyUWf/Jsfr5/
lnPYRy6azQlLiZ78EV6yEY+W5/9w04H2Nm998zyelNq2yEGwOllPja9fG06AktHh
YmY29L9zz+qIIBI+doBDZPG6keUt+2EtymAQeB9OwfPbvhw9HgySv+JE5+H+TTnn
NAdQmzVADBEAzhGG93u90euVD+k9jFaALjz+KJgZealIn6yqsrNq4HaImw0uWf8V
zXZNpyIaHRCycUramBE+elRYBvAQ9UtNz/00JsmTAnPug2iGz+CItRAMz4w6fL8W
zzWMbp+OWaBdWj3Kmt8zczFVaut7gTvSftCl55/l8N41RsEFDP1GgGIaxDWWFJXk
PpVox8wkSJwk7sXw2xwDxlWn1wuVhTccgaDQ0Kh9Fm4leupcJzXfybSksgVkmRKk
pIqMIG7e88hC+Yqvv61J0lVvo8Gb/6EUU8fvNH0cbknrauUOjYhQrHE0ALDn2LFu
l1pEY+d3W7c/x528qNw2ebjJ+oVtgET6KaeFFQQ29OE6vKnxfgdrErv0+Nyc+zaL
YPVpGYsjB+eQqrT6Ol6XH8jY/OHoOh0NG4bSAv80Vu/QrHIRsJCB3NysKoSeeCFO
ho6q6/lN7C778l9KWthHnuLdYNug4L89rEEa+kOpMNy8NSKeQg0TpTd8cwchBJHA
flVyrEJg9KlSrL7Me/iXFNCGj3N0mKFR0so6I8t3sMaz9C3DjO8DmxJ+wkNM64hz
elTK91YJ2iKEe1M8N6GiChi7IVVObgeEeH5oQot6lqChsAt7VTQbKCEJRpEjfCJ2
YhgCB6KJ3Zkc9TBsVovF5r5aAkYKOIhYUxsltKxo9OhvpOXPAX6xlrC3U6puvyx4
AbPSIgZzaXi0h5RR+gRWmu6aOEDwRC8HpPwAlKDagPyHD8e7cmWqMvmPl+oCr/j9
dU68OFaIOMy4UQOvm6nNHtU7RAc9MvZRcmjmr/yJIyOddas4Pt8OQWhaNRvnur31
z+oG25m3G10jxbtmY2imoh54dj3ujGMfgnHQomfQDwb56XSv6efUKqIw1p1gYuyA
Dvx04jzyW7jZHrsbH0lJEXy32z1VqwyAmrL95CyH5kma2uHIMIKNJCV3paIVSnIp
CrADunACs2w6HcncJYmKvbohpS6BQyLsy0q+AXVhfxpvvINdknXb8gnQOH65+dzP
7HzGGCX7xY1q6cf8PQ+NKnlg8n7O4QQRCLq2py03UXPHUB5oPWu1UE9Slu8jcILu
ZZKi9CZ6VDH2FiiD0nYDFsB9zfDaNRr68TcKS+AufGPv5fcJlkN2ndITZp3kq3kC
74ENBGIg8zvTD1sj3gjJlTLTx2ywzltD1TjMdk8hsSselguoi2s8B9IqGVt+61gc
ePs12ZPLM2a5xq3gOCk8qeo1Hss5/q7mpqdwFlHF4qFseVkFhY+oRJJMtxffBGC+
gIRFQQ9ScW4nTlN1SoKtKA9beULWcYrMaKdU2hqrcbBRjolthj37CXEkw6I9pv5f
5ECAwdAGB5L4oZFuYxKNCP3bvaUklVyR5fmFQ1VvixwoSjai7dhlBxteiX4thjZ/
Eisye1c0vmYwP/P7Q7oR3gUuEjBIXy5+ugQxkRWqmzIgVO+rH2IsYe36+QG9OENe
zJpIsXq6zltCII5waYOGFDRfTzGxcuMSAjGDSnFdcGcuYKJrkG+y1D9kNV5eAivQ
BbM545quvjhndVTXJ2WgNuUU9IouYpCDxq7oYIKzjFivW/INfScTRqaXdSPgVXIe
NwLLMDufvJFxioowbYgQHVNk9vakZPMxkOnKPxklXlM7d1pDECFFSRT6JLZjItXf
COJE22Yb1RrpIgLDdpYeouZTCJm3VuPqVNKQXyTR7IXDa/xPM3lemRQYXoaGEi8E
Va7holhruo6OFmQ06U8kgwf8tSnqvkE7TADcX58WGYfs+d94tXo3c7XqtH+JL1ey
4eiJJ7i4wxUJtD3JSUsCawWCmEjTW1pBHLoZTY4HWi9H6vuMuY2nFH8Y+9ZewMlG
afMw5zO0zxkYTojFhdFX13fdgInmLXuFKjsYBnGHlgrXR+lx9+TcobY65OaFU7/z
ysGhyyFjfyFK+sKOJNGXrqq/pQyCWU/9IbiGVXQgFv0eh/PYYJMD8bKVtwnGJ/Lc
4B9d06OKEC7M19CQ4/8qhs+bqgJMBDgNesmYO60iabApmp7fF7ZYD6LZQB2BcvAU
iMCPNpxbL3Yv2Q7Zh7vm3DW9vZn4JrpP/+viH7Y2/nAcEvN5gtz1tf4qKpFjcvrc
hw0Bv89yq0rwrPFSnH+/DqUX147ZC/AHf/y0fcOZ1Wz/Gw3NHwWccSUmrop1aDgS
dnodxrS68a0K8z2cMtcnrA2ppiHqq9nIvNl8xRD52OOaU5g2jm5hssde6cT7OxwG
kJiFC0hjZsdVyt4QYksfvGVJSSZEJTY+X3OlApt4dpJRrfdeaEoZGQr7ZjS6A2cp
NFMSQuhiwS6gdVmmw8PYP2sucrS0u0NoukOEKCi9M0dMCMXE07RwZoO5yAHzBScy
HvbvOm52Ydbs3DUkvMhYGcRgm+YgZ34UqmiihjRJXh8f95Vt3aQSSIg1bIdsB/AQ
G/zUkuCjk+ubkenZ450xKX1uuBnqS+Js92/PaUMAHV9l+HfUAFqEESWcvWSrnkZT
Wv0XDpAl6p76nUnOGoxw5sD535nZZgDVMN8QNnJGrQh1bSUtYld8TwyjbQYFIw0O
pBZKJDWqYvDlTx/6GAjyny7nPhYIyQul+3c9jAlVhdN2+6EoGcZgAUJtUylI85Bq
PX8agc6AGP2KwB2/L1xsGMXIaqERahiAk5A7im2vML+e0gBm8URNNeTDvl2xFyjU
kqDpW1r49huwzrigg5jtDslzYZwI1vIzqtknspdFf8vMIzhks9FJcx73pxIeSaa6
Mg+EHhnTCD/6D1YzBpyd4YobLaJBiX3ar+bHdw9e+e7+kwUUwD7svVVk8Ka2eHbD
niPca04l0M/ddDkRW1rdo1hD4UXtKJ7lR4btgf2EQgwuxu1bbsGVDu2wgCVHElPD
VBwjQCSZa1QizVHByAzrepKBS/rW/+zVxKGkU7OM+bmmi0vld7ZTe17eA8kbHzK1
Ubxgh2gZO7nLT26OL6rjqn0B7c9VnssLk5XtiSLs5MK7XFa7Zdc1CVcj+22u0nic
MPVtGEWtMlZGVVcQPWSujGDDl+nwN9dJRBgDesJ1TYRmHJia8dzd0W2sZMq0PnM4
A48D7d0Cj6WXAW3xHFYtJ9bOkosvA2ds+imFlFwAPspzUix7vPZbIjL5zstiKFOr
e6wCOobwSoeE/yvyOkh9wrMoZMsTsSU0oGD3seli6s3kxvWFq4q/VUBgkEJ1xKC+
qv+WJ3R5mkHlhxbAfo84RDIMshFxQuhwhLXFbjGwGkRyf56dxAYF43Y4ktb0VyoJ
UwYACzwjSNqSX2OvJLUcTIi1ynVWGcgphnZDRjXkK6lWhWT8K/jMVcxAfR09p8l1
8D8dKdUQMIRaDlVR1AAYQrWunW2iH3O6SPC9NSAZVsynzp4bH1Z0oxWPN+GJR7PG
pT5B1qO2E6qUgpq++um9YKUnXy/RSupjkcVFGbESRmiBpSppIk8TOS7JyVIG/HvE
jCP/v/iUi7RIeEtxdNTvuCZx3qGSaFPXPHSKOZN24wtk//8PrYr8RHpE3+AQQO4U
BY/dNp3gi1XGOyoN58z99paaE+I/AOi7UV+KEWFesQQWx6ltCPFfath694ROAQ0P
40NDmNaa8+RIlaHe/s3bkX9uLbDj4UzqbhC8SSErrJbx+95wjgv646TINot5a1tM
Xsx7qNfL5vg/MaTor8FHaJDwRy+kJ7K5EZZWj8wHcmkxoGMJf3l+V1sLT/1qW0ER
befvXfZKTW2noeGRrwdCB0w5g/FQTBawi78psNFDaiJ0iRt7GkJ+qNYo0ACb3CF9
zcY2+9Vyn3RW360GbsNgJRkKYlDL9An9r2svQndIsWaAEJruokEnXXQ52PilVT+1
NdHQJ6BsN98BujxxNvRLPlvjUZwCxaFOyX8xWquC9zZaGyarBQB2TtnwDHA3zV0k
AMvRTbkcT684NAWA5mbRQkZtsPnkzuP4qRzH+DAnrSjFckq+Vzx9CrUyOXAe4OAK
voEqxvLhWdH7wz52+ItzuQow8J5lAnGnjKGDboZAPpx1pbYtodKoon4bMSvqIVyR
2iKHnyTHgbwFxEZ+AZcN+PnIhgMfX0BSFQws0DKUxBQfyvG6ffBDqPiow+blCgPu
w4fn75JepqZ5JoBeyjkukUfy1wGukWZezDqlUy0aUicJl0jGlZWzrsdKJj23ZAj1
cp/MUjWg1yPg5pTdUH5ZpE2YsBVHMnM1T3GXOx30lxQfCjCk6IHFUaBMafA56FRh
husk1joY+8Lu+APVY57kzKXfTGjfxzCj7HoimAuKZoKcLTtu9innvu//khbTwWS4
ig59Q4rfyFWGYXABd7gKkWqBfR6Lrc/xyZe4FOB2U4sVFZG/D7LEylY5A3dkXYuk
oFGO0dOcBGiu+r63Wf2hB/twqdSCz287OfGNyNjgPWBIawu8fcVMU1GldMqSnO9Y
fvosOx6iz5jHzPhcLDIGx4MhII8sje1EkLR7QC6TYFam3dzoz7n3NMEvq+lNFZ/k
af4yzxoE/Nrlrjr5NzNl7vpgWgxTOKnB4UCFOB6aGe9HU9qxPP2YWEoTWzcw6+QX
9cuRRQq7oJtfN9R4nNnv1Kw6ILpBvk+jPNpBgepKLF2eqbwRhE+kdBCeD6COOAFe
4gBOlwn3gPfyNeVvgZVnOrvANAbudbn4SLBA4v1QoW4uoUnJBSffwxaiQe6aCj9a
79tTFqVpOPMpGi28CuGXlGAEbAa6UCW6qDR/lckK9MXVK4ea2gyLYKFCdspTZDhS
Y3VJ8RWkDrgAiLHUXEObrYOudCnVulaCKq+IlhZaFLB4sRgm3Xeq5Yy+m/hj9ZaF
wFJefRvzlLh7a9TiuQO+Ki37ubeuNe1nOBsYz3VzPR9s1ziWaA7jsKyvV9Zmu2e7
fglx5XnukXLdV+0EL1FgP+NDTOTeOEqBVPruNqfkIYTu2DIo9dcsxGLaPe1AUmJ3
EOKkfv3AGnbyF29MUIvWsW0m+3e6jErCkdvl/9OvLFJd9P3mt6inKo869vq3X5JY
f5BQitYL0koXwJG+Lp5FplqEDSitsdpYjYVESV9k+m27E5IFcbnFbU8rvSWNO1SB
5OtgkFZOtbc4Vn4XN8bI0tbJqb19iCUolskmVtCirH6EOJQEg2B2fkt2oR4+CWJa
X8H1GGii7jXx2M6JphqV04BsztzNc+kdUdLsRRkgS8dx+aeHcjXVmf7THjhODuLa
ADUXngmFfdn5g7NJ/K9SIMpgt9gPnUcYfGrqkl95MN9ldT0oBFHPUhStQjDW+Kd6
grAdtJiv+3Y0B76HEzcQtRgArc6ZiO94cpNs/RipjHablIn+ZMBDura+JigOxqjW
Xc2dHAQy1eTEyQF5vgnIO0DLE7h0xCeannDIoJst6fpiW3gMvSSg0cHrkCMZ+aPf
1lFCikrnFgMwwyLcjz0+kugRle+j+nWr466xuga8NPGRgnxrj1maYri9Ka83hBJQ
nkCdF3ZUSFuHO6oJsDg0p7Zx0a6l8u5xASQ3y/xY8Zua5qtdw6OWeEyjWNeJH/st
/jg0HjMeZ6Eyc32mvw96f4cygENF8Mx1clY/0MVBMjKFRUNoCTwZkqEA5Rl7r/ab
cAo8+TKBUZi+haQGPRcfIxu96Xwb/9scqQFEwQfa7k0peh/k1+bBmuL6gjrAwQuZ
9SANCrl+EegrnQATTrI3FpW4W1pY5Q5ZqBtcSjXGdRSgwH0oheoEyxw+WWqId8mS
3vPGMovPEmT6LczK8ZibS1Zj9470rU8auKbuih3TzdaCZ5a2Hwk+EMul0/Cqdst3
oBWp+10xf9j3/6AvG9XtgYI/QMr0XyhljnXdN3CXGu1lfd2cb/L/zU435su5T8bh
njkVpEbiQX5OZosqSmLUjA/8QKIHXKVQuy9Kx+H+uZOjuhnPG5hMacpS4WM1AU5+
NMyKywDu4+mZxQp1aeN0uL5w9rXdtWlZKUFKQexbEe+2Y2q1lIRiMRPe31/+Cywx
btUWOtn6igXHrw02fpxsUwb2QO3DOe5aX1dchYFoIaJTqowUleQDzZn0YWNLdtBT
v5UXr2nzYpo7l7wm6B27iL5mEyx8OfC3Nhx3RK/wcjSwxrAITMeNU2lhDVYW5CyZ
qO1STQ+ubJGd+j4SPfJf+fZHua2iIT+GlwfY/6TBksiHMOIODL8IgMY5+38qnkWN
Y7CMBCc9NhyZo2z4JZbhc1IUpQNxuFlvYmpQ1hANPR9rHousqrlMSf6F0DnHWfXw
AKlOs2tQN4aVrxfSI4t9I13t43LyrxnVSu4UwnS4KyLhdJmJqjIvD5Ajs39AiHik
jl/s0dAejeJDJKI1ze+zi9+eUlPdIrwBGhMiTHKV5mDsjSfkqtf/WWVSvEYvdUED
oxEarOEyjuUp1neYhGvOFS4kq44hh9LW6fB/yBLoZiDslstuXNhOUqmPcUGtJjUf
B6wRD0cHhx4iXEElAnZsPZ9OuaRII6XXmo6j/mQFQd5D9nbOfn9K8mlFiaUqKUZ8
96Cx9NDxwbEcG6bSP1c0sNXhuM7Ebojo0cy8ZQbLnjAEH+gEPOuKdVKYyIrDnRWm
FcPIkOsTtpAZm1+EBjZrWIYkTeCTum0e678/1VteoD+CpF3r7nH3jCr7XFh+2MBs
MCMKcZTLEMy7iwhtw4jmcRL/GJMTv9E2c5IlvGtJ4ViZV6YoMmhsz67t8nzIOUqR
eSyN1rGmUTn5xAtSsvhzOCob+JGNdeJSduTGYWa3lXnEZPrf1m+swI9Cf9QLcpgr
dOqfElxMbcDLTqy6oRUzPOdd15UlOBBIE3oX/x80pMLdXFyIEm3KNCyyq+6PsZ3n
PQ85V+N1udVlKF2rAxqa0NX7aB4yhnNabFKUXI5RkdfRuS+hZdM3p3QGMqFOf4v3
EbNi+o7w4TUpaR/dr7eZAfKT5oUp1tfWcV1uWl/YkNucq3hqcM+PhytwS/zDpc/9
whx/f5B0Z+Vphujl8rvW4ip5W1Sy5DZ8//SGA19wlRV1TAmiw9i+P9LcpO+oo2DJ
pUQ5uqlG5xY3WTzox5mDiEwJSzrVHACJm7WBgtv/cEHem6BBP6LY45FJhJ/9qZgW
rgNE95Efbz3GHYefhEqHvsQz0drxzBphnwI3Vj5/I+ha4gEVXyX5KqcA+qnRlY2k
+eB0TER4rFR0/+QnZkNV8uFOBpyykABUThJrcTTBRyWesyP+sqIQHEzeFa+IQFLh
ztfTRQHfhvQxSQaIlQNWfCLKDbfXTshaUhw58sGi3aMN1OMrkAXrcCW9pLhv0Ig/
5JOhyq8mW4VtBFD67NIAEEaJfYv1hAKQWdv89lO44KANmizm1KI1M9EeDDec6ZqV
r5eow/gQf6n4TwPgpemGf7ybyaQbpLLRxpQGiioOffOxC5oReJwBuBrW87LscZvW
bSGFmiQ7sHM8VPqQzdB+Wwtqoo2HYJiVqYbDFE57SNZ/jMOXPBDk8atAvGtwBi0B
hMBpnsiFJ7l+Ay4Q65kSGpBKf1DW5fUTxliLGFYZPF9F1+6ZZdUSEP3dOyrzKpnu
Wc/SqTr3LqEffchf7YCphW37cO25UfO6K5o7ZBOv60CNyfmco/OQVr9BBGVYOz0z
xGs+WiWpv8mP2x0C7uhlyEzLT8AHLSx3QZ6eJaFj2/bDL3tbvKAsk38YmkimhJ18
TsONMwjGN7qkyhNQ7xOT+PkhWCV3v9EUmlge9p0RUCUB5Cerm9+qCK6/q8RgmpCD
lcGjtzBXqhOpoZm/bqTY7ySRfuDGjpdWx9Qkk2Vcv4TPioADOVRKajfQhH5qfnhK
PZjULbC/cCzQ9DEqx7WBfIgxAiEWxzEbABc2fgAA0g4tEe1dyvP+9B1hMc0mZB2w
cyHL+zfgaZSRU7R7axNZM2L2AMdAbuav5Ve8RQsemUF50GFUmgT/rbAN55ngez9j
mCqHHo+C52UZJNM8C4LQjP0TF80odCI35BjaZjI6mN05PhvD1GjmVN85tL0QTaUl
s2qQ8nluKvvjc34iz6AEa8miAGTxSReUvjOzoO/tOzgCLlce4bN5b3sFI2v4caq4
PBXlCDxUWiLpEc9zTxg7GcZVfg0op4qGVb61KyIuUi4Ygpg5HHxVSnTKbD9mE/1O
GaOWevZDllLIjTnq52aHzFlDEmd0BTfymSMpuAe/li5M6Ut7LLKSir1cpxEP7lO4
utqcxI3wfCvAy8IbZqx9oGJU/dWivApZQ64+rKF/oA2CvXQfuOq55Qg9GEHbSmEa
jN6xBU1xOcXSOW7921lQSo0c9WFSbEaN11AYQxg99BsYew/I7cAo9E5Lh4KINVnR
srO+xXaYVoBr6Jw37qYsYaYTNGrC3gLLOuK/KQjGSZeagQmd3OEmSaC2cjzc62nt
ok3wIL0RxD/NJ/M6OzOTVp+HsXGR7lGx1+m74qalBwJTH6Xqgn5bOxixMM575SfK
dB4mvrMl1O5Ri94HQYnZmWY+xEQcEcRM5CYhWBG8uhAXKrYNq8B7DRLIeo6gAXqv
A0sO6uNKsIKs6/NgHKIxtjLyQ9N+959WI/MTOMVL66bC7CT59LEnB0O9lxHt4krt
X676CnVicSxI4VhaXTfsIHQ2ElN2/ePz2nhu1/Js4lXyMM/3dUlkcQ7VSjbKVJgR
rEc3yhyGzyBtreCoUGynEsyxTGx0ZfE7FtFSLNSOXvlYLBgS1cEsEofbaCwC3OUR
fEBpdW4bhObpRBpQXdsmnPt018+vUWtLYpyFcVBr9obK8EqGbdET/QINjJWNaNdC
KbEthuje1a4o/iU9RJAfnlWcsE/lrJyxX3S8gXNmH8cFncWnoa0MB5Z3YAPGhFK6
4QWoXtwbgb/+0My8paNqDom9KzQoLX9Uo1NYMUgTXYnRyG8u9ZRSAWJy3taLu60v
+roYRKKfZsHxoU+55L1yjoj5Us2deslnBedvZEMR2x6nxditBpZauOEeZ6Z8dZoT
H9gLgxbHHeTfuzzbRdP+m/HpEs1/FvtQCJaVRsbARXtrkDAlAm97C/STE7hUDHqi
La0IArOdKxoum5DOc+FuHi4Tj+RdP6P7VQKT+tbTNTbYyCR+086gOBqcU0csy9aC
1L6wqal7EylF1lRottPoTHWPQiuQBxNlR1p+A/TMK9sLGI4+7s7/V2wrCQ9KyoFU
PsXvl9a8w+uiu9rV52tPHySbVWX508l5UMFccpPJf4svyUXisGtu8qasukpSp3a1
38LBGde56wpFt/P3Qrp4hl/wn2ZsLCov/2IKCPrI6boKPSY0VZYs50lYDtkZhhS2
buTCjwQbXjsrRsznSveaagPj7CH7y5adDUobe4yne3GPsGny+bBs1TpXhvM9XuCs
hF3AlNh4kNiyTBoSu3jDZ+Lf6B0rgkAFH1Mvlp6R8YpMtAFksYRaPiDgi5Hy5INy
Vcqo6phCLk93yCSdEPmKrEhwEV8x8IEbq91G8I/o1UukNLVNW3O9S9odRPnQ6skV
wmHQHItICTp7MO+getB5K/pIgIwL4MHXKAoAHdMN4GBbeQy96WBXqfTrS9tZR/gA
Cdh25Iv0nP6fe2GiC/FQW005ExkjQHgkwgqAXw/VJX6uVAguPdt/pgdLniKWxwH1
KsMIU/nDBQZeh+nfXHJFsgKGNASe4rln0e6wlKUmeJBp05WjQ5oMOXdbdd8u06KT
aL35fjL7khAixmOd24JoUbbfmabsJveWAsPRX7eeT3NODuCWN6olX12RaHGUeFPI
YvypVonI8lg5YJBBsjiyRK4bND6lyiSl9XjR36exZIhYejvZVZ0qTfjsyvuiKKPE
9Mw3ZqZJvVudmMMM9HEZFDkU0O/DO+dYyiVW7a36HWfGrS0ok7GDqk8DdRDE8hBQ
AX0JYOr2hprPUpAkFq+MWDCvyA6TxRKSbz1/+CzlT1Fg7hehC77dVAa5tgu8A16y
nTXFxhiCyaQS2X/PWNqBAwQi9KqQAT2pHuFRpgoZCXJQpMKFkoTuStkr7pDeKohS
Gn2SZN6P3p1JB9sdEGEU9hJWzZKTqrI4FpltdcKWlKTG4HN5tA166pQKtkuO06mc
oNB9303nCsQnzG6bR6+eWSk8AzvSTd0utf203vJ0vU2pomYnuCUcSyx/YqCX0ctx
4O9CChANiMW554kQIa01wzrn7Nxjja6I+I6L8xbyajMsijm5opCT3Ft4RPSD/mph
40i70sRmCmH5YTwh2i2heS1EaYdJtH9Zt5IAYjnXaeGijV1Y/Cuuj41wR0Fklvih
4ggTCsd6Ju32YC27K44mohOvnWrhinPSBq91lzT0da1t/2twPrcyAhYs9j3yb5lw
1DhsHzOA9FFLpuaaIc2P8aSII58QJgCk1B3uQta5UasW3tmJatmXHb0JFHpIme/A
PG+p6nlu86v3VQ/Gz7avgjrH+Ef/cvB3MU7vR40w124g1zFqWeuxxu1erTpij8pm
Leeh5BaNQjyZDdVR5t9+Omp8h2VtGAYk+5ceblNE+fE7Oqy3p9zd96LNN1Ol+49P
8IBU0FdfTxq4xBfWelspEcVX348/aWlK64oDkDIr7BB0+7nH1pxN74LJwtQEdar3
zuVjKCwM4PSMWFOEU9dwXmewKuS5ucRQdWG3vcwMcPfQ45mIi9+X6x0cFk/BVNM+
VP+1r/CL1NXibwpr0XZeyVjwGT+fj4y+mZRAT0XVqTgIhlAv20XnuTf/YaZWRKF9
rY79fQlWPecx9Q0aiKxbwF8uiHfg5aZuRbHt91BVK9rJkECICadLxkWDDREAzu2a
M1/EvOwYCefaR+vJyKjbP8ILgNPiupyN0xx2WWsFfYPjQkBpY7SOrYuIpCTEBV6w
xDq/E2WWIzWg4DZdpGVIg04EAEm9BMmZLyn+IhVXnRGaBsBPtXP/+u8FS5dJQd4F
9MHnT41r6YePWRp27ikh2ogFzlCixwFBQMsQYQUIsAx+0AtUQHDBen6F37ux5SJU
NugKDlRlql5xH19axRFP0/x+I0BEdG61xU7Q2Ii1UF8DW37xJwbaQvMCchDsf1vm
PSBWp1VPdfoejQGCk1BIB+04w9ngl9bgvPsj8ocqD5Dns6Arb3uDwVTkBGbY9N10
jtU/MZKHpENYabom7XFuZeMTRA5u4VnJnWsRuQ9HYv4qjlV11H7RwF4lDZp+n2Zg
DJxuz9wQdZHNLrFnh7hOvNdLA0Tiob6dN5FLBPhxRJfdiH52whAH/9UIC0rdI9na
nk8B6Isj6vFztTjpokMPoEAhEMfg1FMWA9ci9RyVt7mcHt6kdknxMD4Hv5+D7cYZ
PYKd9lOuBQfm+hC1QPjLOvrNj/03sxQ2m/SEGWLX1x5LOwHOEOXksVpdKsf7YqUJ
ifL5JAyy13NdcA3tr3OR1VtTyO90PqxkYReODiIuL6HUY3VEOgW5AaSgG+175xNx
dFwLYPoSkiOvP7A2c2IRw6rGnI9e6S3m/Eba+l5W6xQxldVjV7NvwAykRy3GfPs/
nclI4v8G3eBM3nkYkzM6rrsF5ggVhoSG+xVQxOXYO+v+r+PL4jLpgtwSS1UE8jJI
3QQi7nWvbuAyP/1gGTpWmmUlHaq/i54hHjccYiss2VMpPcEJ+efiAz320MUomrQ4
RzMe6l4wm+kNPLmfXNgqQbIVjJB2g92h8CypzuMyD95FyuBEG9wdp24WKjP+4cSZ
4o1f5svtLGPjG8PU2tIndEZWbhyAMAic48nDSawvXxY5J3Ud04qCalBOClZOkbIj
DkVgGnvLvP8XsKUf+vEmz8PsBAHlYMj9r72htCG7rHXh2hT8QXkdrr7J6r9Lxhsd
ex2Uo2e9+Etq7GVlgWJHTcERQB2WDlXaYf+xp15uym1/VV5lww4SLqe86jHQURJn
e9v9+HGRQsveS54NWCJJdUGoXiNHE0o/aarUt+SdleYVBT3tjzD7YfgAKPAtLFsE
Mfo0cCEGn1hKiNGLT6+MpGx8HbDsjoXsMovk2avs00LPbVEyuXMIdNpJjiOB+tX4
YVPiy7Armf1Kj4T/dBcGXqPNrpEta//l8aew1AX9peLB8kHkJDBvrz+2xXBjb0qS
YOogsbPjM7mJvbxznQH06Ecb/DBw1WsSn9V3+F9tE1Z26c5wSSTejG3WlKQf4Vx9
cRLpVJwoAkOteLYZ2ja0Jdzf2+yGaTG7Nt2/gFBQxbjzZXh17ljO+vUY59TYyile
olw/WSLXRrB9Um9Kwtw8tmpJLSb/o5kuzzErHtiUPrzF0Dk1U0XaKHM0zs2BNHgZ
Z4qcHbuGTgpx3Eu+BUya0n8VQI8HsfJzH8OKt4S7vIJM9ga3dHgueFv4lKFNdR9J
nzaVIC38lrkDvMJGIRh7W1PvnAd9byOD+qiF/NmNhVQg+c1/7CMVw1RmW1WYGBcW
aG2cIkLmAXisWTtdaSiq/w3Nlc7dpT76eetucKb3t3wNKskBhu2N8HlB43wG6XSL
IA0Z6U6Bv+MKVDrR+D/CcjtcwMRltLOwF6XSjqonHnfJ/h0U1X4AftjNDsLKnQGN
5Xos7WZMjjyHXR88zgrlZnv+qKJuYreA7jcVhFJkt7T3U95uTJtGpOsoraDoMjxF
JBWiJUPqN/4L+FECaGGpkXQ2TBgkfzmSNhqxzVNWITzjnu+2Eojcv4h2FVXHgRrq
PCdo3y8VwNiQ0mt/AVdXDWo/DLxVv9KO6uAV7jVkAJDTwIVwUmSPLA/htu5amlsR
cyXaz/121UQ7hssh/0pJuBlDHOylXBGYjO7965wfL4Yl+46zrHnrrQUSonbrm5vK
VeGhzzW2yn4CuGK0K5BTWp+S5SXVjqjYmE9NJZ0zqPuRmCUTdi/zXPjF3BZZHKrr
Vr0O3l3vFRJSF4aGjenjpOenwzJ3nDaIB60dZ0uAuO6/CT+zd/tL1vxiupnd8cbj
g2i8PZwuykHdKfwNW+i8BE1ZKhCivvvI+Xp4cFYlQ8nsn/Ho6B+QvOF//ljAAk+2
rga5YaF+uBRcxA13Hf1/7v+pkYUM3ChG7xmwZmq5Ewxunt9Rq2RlVY7adtOYve70
n32e+xybVyJRWo1LjCsUE/iAGo/6Z3Dtk8NS565INSVuFRUrYXwqAunRZkWkXwhS
VNWLd8+6UvHDznyUoBNB82b2lWRReiENZY6+C1Is/QQEtkDyqpm8LD/02kuSLOiU
53Q6pZqH/X3RG6mfgypvJwUNHDJC8tFsBGVuEqrWkCA=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 22016 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aZUBr4JsYgrjEQQYUVE4uP47X9KAQ23Yn1HwBB5gGrp0
YZteGlkNSz4tvoHMt0oz0s2hpcOckPYrlxIrXCVauztmS4Mdhn1/nUH+55ju9RhQ
Qwue5naItmFKZf4AVizQVMWLmXaBgdnJSsa51kE6Hp79oUIaDfUurTJRoHdEfZH7
NXuYDMI+JkPdGIXdlYPV/X8hdjsnn/SCP5k7n4s6qXefH8Vax+xNalutKYEPx768
/JBB6nB8iY+8rsPrC9PrR2ub/R6BQpbSBmJqhWNdDJM5fh0hWJY2CgPE8ZSUStBW
AzcohVqlK4oXdHcJCO6FpspmeLaV+O4iHeYMIohhrbNgwgZiJtE9D/4gmK0WdSvq
4d/vARzyemNV+rnZUsesTcysxxffSbe0i/+27znwXn6dLOwHEUKBHgZWHDQlZFlV
nsxdNt/urQtozW4dBAjWzBKaJk1RNwKhk8mPJT5+9xtTZOGW1BLxsVbGELa93E2V
2cOlvYpND40/AZF3NGE2A4oHKuWZmJvI3nCWdUsExqdVPwqYoEKZWc9IRL5V+3ap
2J7qju32/n/d7WlQNANh4pMya8fW8TwOKSHnvKZanzsUWTiWyg5YjnJS7oz0d1v2
8MbaPg1LWdy2op93Ia1wUrIBwF5RArBp7D06hrm59ZxYdI/1NbEOSNl85jOdVQo7
fKiGYc1xBzRQC0zi7fNvHmdDWxb+oXIpPb7Rh7j5s/gDcIdp3ETKaK8P9nM//rca
GUMjQQngaQhQb6kkEBHZ9TPkORW30NhFHBcCh8vpr8kjBTeVPQKxaj+gfoLfqvgE
16HBKy0Z7xl/WS7zV0O/grz7wAvcUL6x23hqESS5akU2P+WSLo0TKv3twF8RQtob
pGjDUWNMByyegaOSohTo6Ognu2oiaML6hgekbGNCu82iveYuiLT685J0qJ/wyG46
f+XMNk2JAy9HrgDp6ewvOOxqAtufwfaJg3tHdIY37QQWSfqXRf1FLgx5n4cRHxqm
Kg6zgdLeRwflrSP2kWJxOqTAD9U++XUdtG/yvl1Bf0dmsl74u8zD95NPtua+spId
WEv2E+7z06RDjlCh7djOx/mBjELd6mB40oYs9ueohOJ3i2NBFk8UiiqdlPqYue9b
YLOSsk+G3mZUH+lShEj7mthDmA653pACYBqF/0zh3pbtHDE61XnXaK8pA2itZP2L
ar+KRUYk6fbcEkwIxX+jmN0+ycFwM1krQKJgra4TzK3lnEykW+tR2YGjcP03jHv+
sRRQpZxBOHeefwWbwxBej3/5KP6aDKQLxbNDA1N/XL+bHFCZRRF+6Yd0fzirJzhS
vKoYQMCVUp/GziZRYkk124qWT+RSWjL+lstZxvwKG9Z7TTWc/l6GleY0XxvF3ip6
hHlwRveue+ij8JN/UzzT02mSf9WhtrVkUaAEFtXlOjy8aSdIgHuVn4G8E0vOiuYt
IRvW0djO2pheXxdD9j213j2FVtFwxFjNvst88neV8QwnJZaqPAy79xyHL6gk6FVy
6vj5FzoFBfbEYuw9+x3lzkXoZIH/FAOHlxyH2JJi+LacKJVjSIubC7aD3USOz9Ni
j4Q5GoR02Jmf75ulac+6r0dJlEBgesbx71y2m/dfL9ek1RaeAhjjDa/I3f84E0IJ
e9PktvKyWLWWlNCdQeVKsE3FAGRzCnQGJRcfZzG+/07OsN/67q3b1ajgHhJlN16N
wYUO4pCNGt3mRzigFfJWo9Lravi+4qW3mlQD1PnbpRkU60wiyahCh7z5kU9veY8A
ywNvfb1AscMk3cvC7kf6nEI/tGtTlqxhFvGBvw+kBB8XprL5by8nDFzndYL2O61E
ObbRGBINpGf4O9J+rQRQuNfaexDwvZFvk2yRVYWg18dKDcyTHigbKQwG02FnZUkV
FIOoEmHjaeZ6xK333XEhROt8+LMkVZQkOefgraaPiM7mJKCviPB42ImhJ/Ghysfd
/DleYAV0KnnBpyXX6iUGxCSgC1EVKi1hV7wJ5VLb5e/BoCPpvvZz7lvMfg3D8eoR
SE3JOH3RN7mSDpzQNKMPpRJvKVExOGBHnJyynV84WiqoOcgU0/xf4yp+T4wVPfHs
Ze+gFIvfMpKB/CGHlq0whOO8Xndonc60bXkMHHMBlNfQpfm1sDWmGqMtVtmyEmnZ
j3pVgCq5E7ajhw8OqJOaX/I9DFRQAcIYcYlBk0rFqIz0tqwyvGTgdg8ITOYZC1jv
yqAsl3eJ/eNDJOsS48OcGr1rpTnGDqq1B3jkGRkrs4fH0V5qLrNNW90+RrYwQbFT
Cif5xuq9k3JhgugQzY7+kOja10GdJiITKRKU+j4D/1nhT/DfQFz+z4E5cu9TDUHC
lhcFjVznpnn6LOn6cr4JABycnmAhjE1A0I+mcqrvafwjiyL2PWR9lkAd1zcOQ3rk
dn6JGmGgWu5dFJlWE9556y5rmlz1mmGvaoyT0XyNWBF0kbVRDUcdedJrquOelzqC
645EtvBQS1HMfqZ97RTXXrD2P3dDN2jllo8lEOp4SLIhbOzfXw75MYsxIRNxlwxt
amN7YUi8cRYPSaBeKIqRtC1CJR9qUFIxKSylBSECibbh9XrGHwqYehPsYAgwlKSp
PYbQGEaB0YZK0/C4jeSlnEdkxADdBRRfHUIf3RKWwqboFQTIwE61zjS6JLK6zrix
vbHwe9bJkLO/EuzPzJexeZ/JNGIQs7m09GFN/KJjKICGqOtBANyOxNR7P77LjdPO
sX4knGx4vnTUzuGUHAFfkbrVDL/+B71iooGa2fmCz9uNRGLtSoWuh/ppp2f10820
jOVAuhiLdAvw1GbUPFfcKJauXtf9XWvTmVIStWGXW/pT2STRi/ceAIp3DEXwBpyf
LzJxnG9k3ie8XXJApmrpUc68bbXW54tHjBWiT2AXCW20xAOS957ljHY0gtp4Ps65
EGcgFw1dbO9Arj5gKrphuPCxn/z2vYxyVdaiBFGxxAKtUjd5VtCTac15c/IgAcgT
7GzdvmZzaT7UJtc89tIJHx6+OiamgQXTk1FHAEr2Fxt0F70AumR9NltykO+eevM/
UIK1rmHPV3/JgoARVgwaAaxtgAkybNRXbgyP+nSy9xDH6yE5/tvWs7y3JrawMVp8
/FGqY6PiaIVRphO0kgf/hpnh6ax05gYyRdH4M3Ed5rk8JoKGmDoMyqNw6WPCCOxY
9LR/nRGkHUWjscRnsIxr5LeQkhD3o8coDTj92XLz+fekbcuf0IcAzsuFUrCDF7MA
fXK9R5ENAzQ/JTClQ4IC3OOea1iyffitVdMF96DVL4/1Oeldap/DDi+FU8A5GeL4
oXKRFZ7ZxGnZCoJjZ+0pO7Dgd/f9csA+DLEDTHGVZI1G8NLDOm6eK4GvTdCGq9fW
cGYf15fjRRAFOnwKGoQcUcz1HKj3QRFFwH00/yvVamcIIwIj14ZONyLES8jMLNKS
N8kiyksIx7ajmKeBd4yeBy42+1qVvxH7QRnd6CBOCe6J7MkzWkSwKoepYEXM6a8Y
ir/Fs3FXH4Y9ZJldZZ4cJdoXyDjw09ZNOfBJTOnIqNs0DyFyPeTdiYSXrHD6XUU0
elqEmnbIEPiB7daHdy9d8ybm4pexyMk5J6l1tMxxu2DMnpM+oBtuj8vA5CWyceAb
AA00UDAUA0OV6czjDcQ/5P0mv/kgkewD9ygQ8+zyzazmbz7X8pwASMJpWhDjL3Qc
chqtTGmJ7e5Pu9PtrhIFJ0eekjC8QY5wPndRTXnULWx+aejN1YTRgjUlQgOZmyvt
fdeGX95NAnN8ZW3nT0yVYowzczOW8T6z4mlLAnUSABR7fvrzKqfK8IbelpElt3en
XRQFfiXFqUorcHNNL7yOIl68VLMjhFIjeScxMh9E/H9qARTnzFp0oCkbnSGgqOI+
x3Qn6iyK4K73mN5N6CSSZA++8Cqw+WWE4gqjoCS991kBkhsDZMZWXwRN18zbZL2l
opf98Icxc1FyN5B9ruO0A+wzxVmfX9jGK9NpB8P9NdfGXu71+DTqukkoGgkv3NqB
yakmWaCwPfP7w1QX8oJ7nsj5BNVBPX+v6ORKXiXKLsSomZZ53N4MABlVrCXRyHyN
Sns+Xcw+SfPfsEAiBVOYUkdL6OA5VO05BqK2qJNRdvr46iV7XSGsbB1AHNEtmyq4
qPbKn36ajNHwEsL0EQHmbXoaB11cRgugZdZMiS0hImqrbWK4W+ABTLbGLbgfEW5O
PqR8PTPM/QgLPouxqxlHpZ96PMsumQZIsVUqVr5CTMI689kB1nkmzyLSAMCmtLO4
ehdE1b4R+rcIEkzMEV5ZeE8JnfdmV4bykjqCL7MZ56hPun+Yn+7Q1iBffOHJrhVB
X/u2VNHWo89s41meizf/ELFHrEXIXBan6igr5wEud4pZS6zJXDVBShU359IttIjV
EzglzSdhxnUcuDtkeHKcwuzBw6YoFGBM9JhD8BXDKTZpxaA3m1xs/ZDeOLaFnjzJ
Oh75bC9OAzZYBGvAyPeVpGUjQa+vBOt6eHdi5k4rK44TMbnmvsNfvBC+HVq1CGIC
Gkw2OLtXIFerByWCnbD88ah7PX+xnkdIcnJKKLHTv1OZOQ42AAc/kdolrzcdnrtS
JTc3crMGupDb/np5Kzoqxm1tuywvp3D/jZGO75pS5Rl1DoE3Tq5REobTMwdtG4Xr
d3M4U1zb9/eGKdjpwFYNVDKgug4V0c8Y7/o7Xj2qY/k2PexKz0Wav63XNgig31Sz
OXMOBKV9x9x+bH1AKJANXnk6hvWXCqctCvCb24rOeQxjvN3xrNOL5Gh67AFnllR5
3MkMSKFO5gKbT7m4w5Nxra4Inpy+46XCDgK9yObttetRfgBRXLZ2Q3v8bZAmI8Zy
aYtlTg4xwu/PZrS2Dp1TH5rZ4fl7fJjyrIBuJhRi85qqfa0STyYMvrnbv7pSE36x
7jvjr9biFacTYwqD+PHoDEp1f6kVBEYw8I+VjzjqKwmxIUJuiMfS5ZCvpXY7w1qF
8aOj++KUFsnnH2S/l8u+Nhpk/gPp6+1L4IhSSeopNlhdVFTSyMsuC4dMiKNtHE/C
UdRQK61kwN2zCnk9rrAthp6n8WuQ/hsyavYuKWW/o2XnACN+edjcjnbCsAvRSoxi
3SPsfQLN3PofqcKRkfJcPZF4QyHaP3ajYnL7JrxnRnRRg8H6DCvOJuCad+FXWuEK
0KL6J6YWwD+5sUgs2cWQevV08kgbclOkVsza1q9gR5djbqGluaLVoDuE/O4nnu5L
bi1A+rjEOI43l5VwtbXs+nGY0KJw6TPu9YVwr2uFvJRpBbZAsp4IrCAeuuCijMEy
Aa9n3qdDR4Y78MLIH0KpSsP+T/6qJ5cWlv9QBger2ijLLkbIJpF7ALAKgJ3/pSMX
nfwlmvoxn9MAGZFRKJXGziDyrd0t1hJ4odJFHCKkTFKKwMIodRt6lbIDPlTtSnMZ
P//3avHa4wQeN7wtfWJ3YWgdfqgP8psRS8/9cAo/UgfisU99FlMK14mVFz8JB7/m
Wmhhv8hok2x3nwDi7z1ZioJ/HfzzEJo4nwawV3m8O6CO3BkVo35y1eRcn1qhlmtm
lUlq0mYy8TG1zHrO+xFEWYNAGui5BTiBpjbfWchIOVXlsFUm8Brd7kcoeAtgEVp3
fXyNG+dttLlusLR2BInevkRkHLSvaRHVjCDT3uIONpxfU48nqo9asEwVI1QOnf/g
2LPaYb+enl+pQAp4jDkyKcpjO2ErvwsQw4nkvdmU/cz6+CCgQwpdIiCHZf0RRIST
Gr2MwPEtX9av+wwYUVANlQMP+zuOlTMNKNbd9zF9GLMiJyhiWsxbEW3kue6N9Zp3
FMGGigikOx1+0Rxhv3usP8NmKF9wPmKGhGh9zu7Wby0dK6gmovn8QhmWCxtlF4yx
sZymvRr5vG1YvCxkcOO382PDDynLDtx7V9HaJMRZE6wrhDxxu9VhnhywLT7peeom
7/CW9wtS3IdCVPeUIYwjcGjg1zziYjx1ZAixTGaHNktGsQ4hr+mci9Rno9X8fWn3
UeEgGVX9E1Z1wPVCrNHLk0yqFMYbH/8JBiFOZU9mszdU4Z788EwNI0fVGeW50WBD
kBgDpJCN+BkcUvM3QpwasA3ThI5cxLurT0fvNytjbVU42VD3pR4wwiTZrXWmrD+L
D2FMo2jqVCnMzcNELssjE/OTJ5IpuVwuFyt6aYHSUnpPd5aA1n/FJp7HsjG2yrJ6
khSUwKMB8DFENJyz5BDamYOak8lzmwURH6aFGIIXfSkPKBx4+GnL7F5WjT4fQD60
hoJq70Ct7kEaWS+5SuMFXPypCgkTB/4XkvUkuUpgxUzJeZbzULnKK1bBEn50zH8m
0Orbty42wpKNEL8dGQgCMUcOxg8bkRWTZSpSpEFeIUHE0/zgJXNzcfukLsgAJZUD
KdERU7f+Ffp82qkuXKXnLi41kOzIkIVvkRHlPwsdLx+SEiqKPgxFns+pBxxW/RaJ
IN3KSpRSFp8bHIkUWlvvDbsFZCYL86Orr05XXT4Li9aJe2jnXe6i20y8PItnTnmN
h6SDduGRJJAuUoGsiTBmcCQsFWAV1BmVCOgt6JRAM5JcZ42tuIDR5IgweQahj2Yy
HFgrSjgXcH089M2qUShNdTevUVqSFpOR8IfXSeBbo53j5w2RF5Bk3FryMrI/Bwcv
+gaOHT63G4qL/LDlySz6ta+RrPAGkKIhJ5qSHMMkXj7AJZCrpg43ItWnceVCFLs7
JZ8gRzOqju9OUK4BaZnVI2/53DtaMc40Z6UZ/gSRr9+ZYTS152vsebiG/AJKpAqa
rNZ60LCrBZtDZOmhE6RxGOTp5NMIYfN8HvtcifI6YyyZgpoGQ+sJ8QD8PDfgPZZg
Qs9Wa8fxkvtfyrsiOnRFMZLPlfpxv632fOUFJ9iZ2bBIujUvCUvrqXRZHLb1mXIp
waineqAbWhEdM9STCkPa8oeNYtjdhpWnPTLo2QAtAvacND4WY4n1KAdTSgBhs/JU
x5wVdsOQV+sXvWOR7vGC/LtT3YJlGUXP4k650ZT6oja6lDdszpHoQS+A/cY8tkx1
53uwZpNnja1wdjPfrhDjzsIzTK8LZwYm548RYiqZrztFsFRkD0u6FTnxm8bGDVSz
j7+pi4GD3POX7620oTKrzzVstQ83hbiyc9ejhDkgKrMcTySjqeLluljg5xNj8A3m
9evwqC+g2Ws1kSK9JrVEHbVfAzCFrsKLoEoteDh8aVuXzj85PQ3HRG1dyJ5uOj26
QtArtbP0k2ys51/8FypUm43+WThDJzC7kAmx59wwoOvzim3cKv+R4maMVPeeSjoV
A923AxWIyxa/cCaRoTmbEKbSSfSUl6keDVX4JMB0DNCHGbKbPTQhIrRCI02GWc+6
Ir3Zw1Ed6MJvVE617pJMqs+DJ8avr6r/2paw1zilvjq7EmgzxWhp7GPXJrBTXXKr
zQWVlPS/cVBym4Y7/FlHZBH0jI5msdToLKPKDal42BYOahm78t23BLO4SY3oNbqN
eACelJLRFk64eWvvJzsPLZdEBAsGgxnZyNuvbyiFYsCLF1a5W8swM245WVY7ykP1
kE1QgCifc2n7kTFswjdVHvwGzl7InUoDaDoSqu6ovxCPfVAjOlBu41n9fO6eAG0i
dv2M8HWkZZJ1mOj57A1Bpu8GQIcJKyYhOU5ZsrwcB6MJ/OTD2idiAFjntrNrVJhT
T0Ra9NX8J/LKElC92AGRWS8w2fyUV6n5TjzM2bYZ7vvRHueA8OPDf8tbB2yd3hkD
NgfeB5IgFqKiieSVB5wbXgk1x5YP2bHYB0faMgvGxsRf09tsq2w1E56g9tsJKUzA
xlKDDdekyGkd0t+bJ6a1WjiAIEorQ76JBwZH2p7LYhUo03fLYqp1ci9xY65HZ/WK
yaG1qSYjyYGaOFJsC+B6jplAbXtu54VkxzknydcvoG3yKjTS6OtZWLixjFH+rhuP
ED1TUOglO5fZU93aYFRxdw10K31jC5HOz4GoqsRbt+IeD7m8IZkd8VfhAkYe44pv
RQzXaRsMRZbLqnex5hSZk2APK/b//3UTc6SzL/xsRIHBb/lwd1ZLJ4VUJi5m/1EO
+OFXysllrteTUEbpYDR3af9Q1crhgI6llH3uTJ18/gp4SsqfGq8dHgmj59Geciat
Fjh0aMY3qC1kb3l1R1UkhjL2QhCkAriMASx/zmh6opNh8ikDqjgwh4xTqayWWdWM
mVc8j2LbSBlYqB3fH8mCKOg/GN6V6Tbpj+m0fzzoVI0qR2iKwjPHJJh8RByshZVf
XCTjPjal8ytUI1i857Mp1gXN3osqKAt2q9jn+aaaB55l2n4nGCeHFVEOo4EkRsEP
MnEMBdi32lpn27ywXXtJEauNzKqkYlpp7VhW+aPyWdAk7xXZg9jFrk345dpO4iS5
wKW6nPPWLoY7aZmn8AXYekS8OvoXNsamajRjRQMapiwylvKcvcbOhI5H6DUJh/2W
8nm5H8G2bRQCweMVdvQdXTlTgUTqHyG4hzGmUcaH34+/xhF4NPzOT1clpwdMdbaH
NBdOx9awUEbh0AJqkcAxzgBAvwD6yExwix7+YH+/silUk/oPueR7Q+sb08adbibu
6SxQ5EhcScTAYbVTcfa6QLf15lpbViYqdH5aU/YKslFsfkXztyfvBKN5IhF1LXAt
1uhL+bs1Y4+Vef+CGXl7fvwaRh9wrwBNSLtYcYRcBWO3UHMN7fN78vTlIw/3hFlZ
VN/TR+CC0c41kJh9E6qYg5gKG7eOnTrdTv+zEM6EQmKMCqC83d6cQrOCUPlQLecT
UQ6tZS+nlzwX6EZ5A70/xtRDZYZkaekIfDOh0DLV+GKZyFd718VHVd43dfRaBSeO
wdWYtZiVV1wuBgAbTOROfhjBBiCcMJbL5Eac5YgAl4tT6uwW0L9g5Yitb8SXAkty
/ZW+L8h8IyzGaG7zjRsxEywZ3oSm+5disVFVhL+GialoqCaAU08BaZa5jBE5hLzs
zbJf8V68M/2S2KzZj7Y/BSMGyBFOYy111O3t/OBvl/1ptuUFMpDbjVEbtVEQJq9P
WZXd6gZmZUfZfXnPlffC5/rd2Ufb2fqIRnhi5s2VMMG4T3Che92ypnDW6t0YDzFa
662WduOmJkGcXY7+7n/ZZzLe4QsQWy8uepzlusZAtc3j75p857VQ0M6a+wzRJ2wb
vDCl9Lxl+DiDDOIFylz9gM7/w9gSVlebBzGGokNrG+KR7Fq9pdLLrLxnnTb5xLHk
pJRDsgI1+CEVI5IRjHfyef1DZea7/qh17XNPEbrwnvc06HCd1EuNMlu8+6pDqNSR
4TIIm9GVq9m1ydfCE8ssm9iPe2kjPpU5/HlVkyQfL5UZxoWes003dDyFhCUksA9I
lrqznjHgJ/my6roK5p9lApbzdTZhKaaaJiw2WbDdIgYLWhjGZSmJ1KmxbFuW1dyb
YS5LBK2KsuY8/3ILLsmGDkYOJXASTtxp9rv7e11zCFdmj/+da3m3qwb0i0Zgk6zf
Wn8/DdnRRXvQMCEuJze5+LOrrIEgOBLDyc1AdgHdT1t106rFSceJA0SL/RZfwYnq
ZIcH0XnqWNP3AzY+k5Ug5oxrAbSl3IHo+7kcD7kVsONHV5745DvLm35AOHVrroLG
B3bZmrliPSNk54RFZuWt7RwLZWSen1c5wWHofEeuxPXLrGgODNJGuB3X2eoP7Dzs
pZBy41O4iM7QigDRQcSCU12mno2ceRAAhk3HDwSs5NZd9jt/E36oZVz8x19I0Pdv
sREQCXsIa5r85SdFOb9YN7J2k03HSVOPAB6hp0tRhvlWM4fJ/ajLv08QaghRoWZU
EYpcpfjqSW/PbbKDB1mIpK5l0/TRn4kt8t2mxcm2QJLkH+EzA4kGVHqdjT/bbwkJ
0t5Ea5vpa/wm0B9/zhUvnbdAzPLFMSFE45xZQ3apv3BGbVB/z4qo+wjOit9UoxnG
mp1Q2+aQeOpAinYEwwCj1IudhM5eamoQ0HRvM5FQDKw1zEBa/kqFFBk/OfNuWatW
E46GivVW4T4DBawboUV2ejki+o8Z6VANdpN5fnZf7g8kkpIzldJmJ59WKQI6iQHO
o6PAo9kuzaFav1WGImXjUHzci+k6TgTwPLD77yktfU6BaKAj4eUuu22mlhPC+kDd
oclq1GtYqaMxxpKH9VUtiCaxPTHmBEUppb8HM++Pv3fET8Vw6yh4xG4e7xIYFynS
cn4lETgptKSlOwhJWeZNcGa6MJoJelrlC8EVqXReVkiegluN/zpVogyY14JilAB+
8eg5O/R+D5P8v68BCjcIliA7CZ+kAVL4nvhsjTL1c9ebTLMDKgT5OJZsnl8iC619
BQo+nvhhuvvcAe5bZU5k2fCpvY4a2GOCJt3BbnXR7jJUOIztlyvlpL+7wNtdgb+I
K4604uInRBExsxiaLsNMsCgDYL3hRzPmzFP/j7E4DHz3+kcM76HydOe5kMQTaMFi
8H4AiS1ZX+y8HKXIwEgQ9/HjwUS+shLeqhMTEGNHoza7MlP9QvOLfBovTTE5D82+
ShZ7aABnRuKIXnJDo2CqFX5MtjH9p3Yas34PWyPe2SfY7ZaIbHZm+kBVv62iS6/Y
0LpIhYIvPJnag6NC4il+9UZjF++3Y+JUCIFXh51tfXf5XR1YRqW/E/eAvtJtjlNt
ZotH66Ynq2U0MrJmPvoz0hb4n9eZyjBD4bCmG59FGoc7Nxpckx8GIJhgr23NJC+y
nerjE++WPa8U7CW4as452AJfhg466NUyeki//w/r8moNhhxPnmjvIVY2k9Ie9r3U
AnmGCw9U4pMafT6jCDo0OSwInIHapIelqlo4Zu1m9A4WCm/fJa7HocZCR3n/JD7D
isnr6Tm5CaRPfEtD58zcl5tNBsgpNvcv0Qli9Mw6KyDPijfgUgkGSnY6Uc2foK6W
ZknSJNdtr77rn0C1LrFK6g47/TukD2nQ+OOhsEaS7MZtEM991OsgtlYh1gldahHh
zqGflp+xGRJU80XM61OfhPFMLIrD0pwxqNxixCCmLnX2gVGEfI4/zfuR/iDEsoxi
z6o4yW0IEv/3ivg+yS9/OYYFeyoAb2EJkA9oiVvvV31oFP0VzvAGgOIPCtKYbTtA
iLFbb6mOdxOLArZQhm4f/0ZRTaKghXp5jkfpK8RQRbBwvSJSIzltSVK5Bi8OIwX3
pxZ2yMGG1PwFhcjG8UCyEuDqAlIqgTwx96pBgNi1+K0siMxkmFB+fGwCrRewqAB5
W7EDg6JX66mI1R9m3kO9aBi7fPO1DXvohA9ohCcpEljKDmafT+mXbInIe+du6x4t
w1YqDcemlsHQLPigEKxFYElBqWtXfHBKp6AYbT5o8xKE5phSE/d0Ix6uqF7uRaLN
xkAPE8SzEnxtDQQdX7avSLZtKC6Io1coggn0O5TbJ+6wWV8P8iHkwttuJ2RBlz4p
gLsbaQjRq2hUAm9DmByLCMHxSapmn0vMQaSRxKjSSYGhL7nbl0nMaSSEczijFDZx
D4zBLl6Kff/mSrgW7/Z4gPo2P1nlO35N/IwhoG94rvYNPWgqXh403k2N7bY5t211
vftSNhGTStLs+qSw66TlL/si4vvU8l5JPEkw5IUZ9QaxKYUnKXUGYkDfCv1uwYQr
LVTfLXqdykUDe2ismfEhh5y7aS+qjc7CxIkZhnMkuAOpjYLMMOcMkpA3ifIm9ufK
OhLOxYtTbI6jwZKk/DRo1ba2Qrg/3vtIUIwwJvBUHjv1zYlBn2a+TSBJIU+DmYtk
jmGAMYbcTXwUP7Z+DmPJrhrfVjSbkpzmLcZ19T9TtqEb9UCkdZ2HJndKLoaOe14H
ZiXDA7eDsY7uM/uoElSX5h3ckqso9SbsMHOxChZIbn756p74grLvdsH3/HpTRTYG
FBGRkjvrmFmOsvfp03jJc1V4Lg4KoYr1KESWKIOph6qbyX4Iiuldfj8aJBMLnKKu
zFRU5RXZcSktm6HRfiz/LkR1g0wqaUl2UO/n+PRobjU5k8iYUikerIB/CpdLQhOJ
rOqWNjZg9yax+mBnniplmU99MHCdDnma6dSPPVz0kgKZi8jUoEJxNqRN5TYSimNC
g0wji5zjm1WdoBQZ66D6HPBHvyltCnyJR7LdbbihUW2DziQ4p0eZDa420X5monV6
817VHIoK06E38e9v2K8OBp3wburw8jMCmBUd6GMziml05bqYYkRe/RIGqfjYtTPQ
/X4YQ18VKdbypRN/njtDXgB5v1+ulJDSncBWHTlcmqXGFtIEc8NhG+7hOOrLIEf/
w2xJc7339b7vkc09kpHVdEd8OvGZ2RCAUY7bcqzrgcypbn1xy9OVzI77uc97/ZwR
nprbGRWrIXa/rGfg+4yGiBoc0eT8bhhHNKhJZuk/AtkLZbiwXnIcLwLRf7k2FJG3
fLG4tKQ61tR9kapmxs20+qvXDpWNSOT3ciVR8vbhu4XQOhc9jbmZF6QGSuswW6ep
+/AfZvcChTUUBuUiqs1G1MQxBc48RF0hxc3XYsOVzw9B0Olj3Qou6WYNaws+cDFL
qjv4H+lljRPPzDr8kFiYIjpN2kgvDcvrnZ+/bVJturqBHHrBIDIiri9jt79VDugZ
56yQ+JlugrzWDK9GjzmWWi0b+Dywop6ZcY6nflZsZFLBLnSLEkZEGbZc4SvMEKmN
OT8ajpUWGNBcqQVl96S2o8ZCIjRYZ6uvzWCMtYhdOJPnXcqyPcjTTDl145swlhCd
VWO7VXTPggCszFaJAaLqliO8yZ3HsBRlqVj8oT69nUTdeMBLQFSJTYJUbrSZJCtC
aMHWYF+B8wn+YikORjj1R+soen8b85Aq1n8ebEpvdi9n6aJVZtcF3/n6xU4fh0e9
k0TPFLbTxwToOXIlAH9W8s4QLSwGFbbGNijIhjzCatFyPqr7l4n8L46M8bQaJXpD
mzlkJClQ2sEZp1YNSaSnLjDSnPEnTTzfqytqi2dInOPdrySbJ3ReXHnswr7mX+/9
WgCmhva33/NIhxyCq3WrWsYZRUM6mMPtPxLMr6HA75k1SxhpX+mmBjLT+p17yBNH
CRCa50vrtKH+d0A3Ao7NvVZede4j4Vp5T+ASD9VIklE8oH1WDS4QaeGQhsql1QXv
MRNJp4yb/aGLFFzFl4aOPV+lmaDX8MaMaeXLoyQ5axPmYxolhqLvZxFFCjYkeWQ6
Efcz6B2IXZUWUWuNbYkzNtANnNxXEbqqpp0akkCs67swMePES7YNriTo6d4TA4KH
Go1QsM4YCksDbPxZxt311kq3L+HitFhkj0qTZpIM97VDWW7I7/cJAYymh8ltHQGb
phRPSZtiAouyiebXoOS6muNydZv58bLlhZ40LADH+vyNz+XUFAwRkpEgFT8xBjVx
sxunyas2xQK/cQJ4P6xmJF9nggADoU+4fXndmm8+N4J3QJlZBEEqgD3TbIhZWxhX
F4rVrvzkfbW4T+mkgQ/2onEO0Z7dPXVRgPmISkerXILQ0GCAys0Rym6hP7/KkRcj
zJ/fbJpHPmNCPeZhMBHdHqN7A54ZbXsFqj5+NihWiNAORp6L9CK1CaJg+rPiRYRj
MG527+A67mfRXS259ryRUkJvVUELk5QoQcnG+lmEhuJUkebHVYyO5kpYpsdu6E64
7SMQ9AwaiQmGLOneDoRksPMmdPmJUOHonWso+/qakCzZtSgDd6n4wC7kMxCrN99t
UGfGUseDY1mINGaVh/V14mav3MpJRs5/x7RZUcW5LgaeVR6YbSSL1UL0jvPfVT13
RaMfOuZAVNSUmAnYjqegbFz7VjUoBQgYG/Yt1W/BH/hv2UN88DeWsAFcX3htEda9
himKrcR/brZlPOqE9BI3x+FqJp6mDzK5AonYDmHCt8EShUeenREKUKfQEt6KxVfB
9R9zGIipDAxPqjpvXexOiOrc47vdEn5kKrzsSKy4PMBt0nFBwQssHd3vHPmG2XuP
SvaBvDDa/o4GcdH9uAJ2gpS5UGTI4kA5IXJqd2BqhlM4bvQ/z8qRCHAfcDgVchpe
YNvgyWKcMUUZzBvGmcJaj+tP85xjXODz/S6TGK5/RTxG4sXT1EQcl5LSoDnwDJD7
mMXFvwOskWRLbBnvSMKoCbTJANsIFXFsOXv9Ht/+1Ti7WltYwCMU+qH5B+QI5eIT
Bn4fjypr4Lk70MxJu0iww0r0PSkT3u6eDfRAY4qwZIQMBvuo2TnspsqhCmPHsf3f
1S5Bb6H4pQw85vwkK8YEBLtSmbpcAJCKt83DRjdUrvJm8gT78/MkLSFs3MW6ATt0
3NaxVP3gWheXNuXJ/C7AyuORmz45nIooM9aF9V6hbIot8GyYBExRHWUnqLDpec/F
5+UxcLF1kgQPAutEviJ3bKKnpDHC+EK1islWfTNpqbV0vJERZ6t3i42QMCH0uH91
BOtID9nT3v2BgZRpS2CEGBMZGf5YWlhmCCMCRiQZhEM38ECLOEywYAQbo+/hVVi5
O0hGbABD08+0MiihM/wtR00sy0fgOxM0jjU/jYj3kNhyZN6HDZe6PacHhUTR2SW/
7jGpG1BV+5XsVZwA7sqHxetx3KA0bQVioePPvOicDX9eHSz/o8yhQl0b0BmKpuDT
7ja+h33PMllHVBwkOJb+LiwHLapEhcnDLCJvrRL5rRo9bFjeoLRZ/bPQETAidO3h
AgsmR7DanoFY9KcdL4QDSHZ1z4ymYfY6uNyiiykuUY9cFLPoBp4jBaDhhVUWayVa
U4RIgCKzZDWHKEZKgDcafdBD0AMt1N3pafWkNDr6wpmm/XH48wx1+SnlAPbU2etV
BV+STiKX1KxUBTgm0gAhc8LViSa+UmKxZAqQsdS5YDloQ54VNIJ+UX6GW7qWXX54
r0zr0HpaihOPaiKO41ovmlHUtYCxxl0IaPyyUIdGvoSamIMkTm22Yu8J867qxxlJ
+pjOb8xyA86/TKbeTw8FfAbxalbjM6dxoPbG813Tlbd1v6dJHeHtrW0kWXSVe/f2
9L/d4osDStwqZ20Es7HK3SxaYCAjhwEOw/t9jlt57hZfSKFYQUXMFQN61Ps67l4U
/acGxoFkEew+i5ahqLl+mpzi89nM8bECpxNJWirv7alxLd/FBwQgbduVZtI34pI8
yZ0EGwFVb8nppzqdIAdWhoGR0qVC24Epi1FIG5QRomwRs+nAanxKkRvgY5psNPqO
IhWNKJe1j10NULopKV6b1zxDla+vK8fYdxYufzzuRST0SLGZpDdvOtDjM+coQCON
gGAWdiU4apbDM0VGYCIx1eNN6U13wyVgSkF8a82n70mjY6Hg2wLwULRl/Ewlykdn
XH0DmAXv3KW5+TMDUDAouUZhcuPL77utnsk63SHP4Hs+AU5dbQUUUjTNBSyT7wzK
QG/KJFJCIKcv86FlPZfzbcj8mRJ+uRrtkyORPU69Bz1E5L295zPQ6wrUR7iCQogL
Uwv0ecD220zQIqk/BtozTSmwDKg7mCh/dInBEQzBkDT0O3+tpG9A3LGXsVd4Ms7+
fqpn7h7I9HOFTDcXxGJmhzMIR+Q5MoCw2ntBqakmagWeHfHKeFMY0AeFRJYBR2JT
qytUc6X/Jd7qgI1pX/cn+5+1K9KS/djOwNTbm2ZlXOMSjzjEIdQU/BhhXVtReBdD
gRYVDVkiIxTRQ9RVT0ld8qqsWaJecamjLPhrQT47L63HQ1BBfqBOOGUdz2hhgNt3
Jo6wFiZDOy2xkAqBK2nNh6xc4RlV1pqxwetXtnkfPs/57rWZTdy/sJkRbNvs+dBP
6GxOVAqc9Q4B7AGwp0RBIuqGrwtd9+Gml1mAywnCuAqEjLKtiyY4wWFYum8zIXID
aXUvBhKF1U7dmMOUvKF33iYIjdEcT+2JGozo7DcnI+ebzOwvWUj9ySnYZdZQAPvi
R9Vt76ulfWAFIG6sbp+eXXKEdqDR7uP2tqLPyMbWjxc6sRB7LkKhZcU/vc7fyvw2
c1ZaYA/K9t1v0DAJO1nQ9eWg2B7u2XaqV1nUaZBHRXFpYVGnRSOejim7J7FnAP2d
kgQjLIrDNU0LEUSRfEe2m9iRtbzdZm1jYrM5HDgKkZcVGF+0PhWtda5LaTDJsGY7
rbDg8El5iCIjD8VacPZBDyetLjWqdkkaoAuY5SCRjy3PqEPcgN2Z/Un0CW7BhlCu
hIGlphEj+OXaG30Y8RCp/Eg5eR03XILicdcBh9XTaKG5HwYBCH5E7BS6+zV7lpRS
MPeL5JSHSmPtT7tDzND1D+OHtaEryUkFg3UX9W9fmJ3NMo69ayBmJiU68qtY8M2D
hz5LBAxg82vyEBfY7VTSE3p84gpwosQIxYYkQp85n8uxS6p74yyM8c9hIZVFCoyg
OT4FnS9A+Fe+4cMz6wWGnoeOc4mdDcQ0LWsEW1NqwjcwdLIuP6+5YBQif5KCiNiS
GIXhM99QQMfT6nZrm+k37aABNvZzGuBq/LNuRq10HPWmLiJa1VA0DP4TZ6cfp3T/
kOM/FO4l0bxK+sKkY3MBZ+k8YrFM19Y2/uz1HPP2KTRBVr/c9Rh+wB2eeLvFAEcb
9UqDfnjxyJNeZ+56WhNbLyNgyCi4/7biJHmpWjKTBuodSGryjxda1t06Q6nRA9hr
aBVZOHEntLS7nRqcMDKulcl34Qu4UDAhGF7JPAND08/a47ey08xwng8MvUJr80XP
XBI0NnWMJYHOL+iG7Fl5v0OytaSQE90itUK845C132J17D61r9w5lHmHTnMTx+1S
Urrk4lmAXw0UuNpajCk+NKgWLtCTlWGq8X1XurYQO100IWpSPN/ugb8TDL55MOHx
1ZSd4BeeLf+vupnzWjehE1bwTDLbG2CAWVmLJi8TJMbIbwQVDV+mV7Eg6po71IEG
JR2/AmsojiLlDms/dAdRQwEBVqqSGw3EugV/okEF6QCF6swiYZJELtVM6UWyQFa3
gW8ud4d3QnPr2JtRDOHF8XLB8xeLQNfH35DJ9SLQFYU/wHGSi8JmwWG8vFpo+T54
Bs+ejYWB0r2V5+NQyMg5A/Xi10mENX/CK/i0URHWheD8ugPqnhsGie0E02JshItd
zCUs2os/c+YjoDRMMzN88oaDeY7eAsI5qKGlXtiYRDWuslDnwpmhM1qJbmJ/BlpK
gpKWJJa57g6YyNB7jI4BqSW+57RGsPCrKSGszEqKvtN35oB2jgJrggPbQV7+T5GN
1SrP4uVPKrMtiWCLiU85V3qR1eFfnUdwLPt3jCv2F8AIdN8MQBAs7y1lchJsWYzu
ye0B64RKlx5NbBg0JQKyWqYP+SnkRX+J63VlK55PtgmM+osBIAAaO4HUh8Traikn
CwVHk9XHjEmlALmiRV6N2TEnCIt90090XUASqi2yro2FMX5p3LOAyAksdrJekYDd
fHEWVmRvpVSwFNeir6zPULgtm9O4CKABbT0n7eZMkWkaDClNigaY5ZeLTgul4VYI
gTaBxT45soqupQWph9OAcyw+FNSfQ3gF2y+BrNi0trPae8WgcMYOTpV7ZeckInRo
6gdwnA32LoNFE/ysW8CefNTzWeFoAeQpVMdPvDTzP8zAizCEJPamEzFDnMgPt1iW
PAimkvF9WwwHWqjpNp+1DR+RY9axFyKrRWetO5WwE5/wVVmQauf+ORzGLK4w3DVt
BqKsD6ZMOMnJVhIh/DSMm2qKe3z28saRWfiB9IrmzkpJ1u40aRWVakzQyi9J+kX5
Hv/A4KbS+DPOdb2+S+Ci0qXfUn9Q6GsoYntzD+9J71naP3fJLoEmR+XMHP8rL7hB
hd1r/yGN1XrG1+I3HcqOroa2pAFtYxTHSTtHC5NDgl0FqwAQSDQE6DRMguT0meYY
5i0M4jLvcQEc+J3zog6R8mSC7CqcVX0rRb2td1KWc4x20IFQ+oMNuNxF8NSJIv5K
1kYg2RLQQL5A7ET5zDPbjr9TtgsKSV+21Pt60MWl00WH4aXYM2b2OPy6AClRI5Y7
IMQleHvdnp378W132tOpS31C9zOFCApIrCJB5jRiNgnWYTZ7P/gnhQ44mPU2Kv0m
/8C1NkQOcbYTlB4jqeRTlCRio9DfDNe1WjmCL7pThJ/OX714bezKjawpHRghPvax
19MAi2ffOW9ro17rskdMiARrGo28l2afCJiOm5pl6ojefhnPVYgF31cX8vbeCu7n
P6X1VxXPWIvkcwZfEeiK5JdLzV09P8yJFbp/aHIVeYc5TaqrE5KYbngw38o3Qbff
7tRKYynj/GgzRKq2Zy1SA2LjUEIsGtcCTOdynYTAsthCvp9jwwKZiWyimQOBOBmG
NrHzJQ50pUNZPtSOR1SWyvXvT5wI503SVevAidL8X9B1dvA3i8fdTKjQVikM8Pby
mJGsbnriCyqD0mqNAqcoTC2p+joa7cgTVkDwwBUet4F9uEW4rYSmNPMr96jxrUin
TvRNbYjQfNawT2vuHvWDb4vDHttPJb9uiaa/IfgU5naV1rNKpMNnbZupUX5G9XwD
VhYUxnriOTZUg1NRLiPBQzxFQCITV7WZq6/VZtS3mST/BVw1o11hDE2KrY8ghcZm
xVJxzsQ0fThAo8BZLiIqlfVr9Kb3egGAFLXAU+l/VljChy8sQGRC9++GSSSYNu+y
LspGsfTc6NNK/5aTEeiRPLrYSemjy5KKc0rL8Vlsm/leGjswfGohkJOo9bxbcbI/
/BsWAEY/tx1ecteceGus/hIpidtqsVd6Rrl2LjSTQwY+jXrmww/j5MDJ0Oq0yJC7
MeKQ2m4OZCEeh8o92hH1Jjetfpi3k3Du84gsAnbrZw7cNyAg2vrKdbd1+GB2B1iB
/wRq7H8J3d5aF6iFpcHozeJfOQJRJ+d5Y1i7qIlGc1fmNp+ltCpzScz44GnsThee
YIenSPIRxQnrAchCif6U/OaBbyOHqawq/zTX5W5mGotOEcyaYNEQ02YYNs8/BNpE
tFWa3UbMQQvw/hxLyVQct7z2f2wgASCG9hn7BU+UpiGkHjpwdcjFXRjMOa2BZ+uS
dHnuge6EXTy7Te0aFuiSROrzL8wQnpgImzic8B2VZg4yg42KR4k5Q96vCJTzYmya
tTTD7bFNa4rUOlG9Q3SnL04Gh6G3h8TlyY3FKvrNYhPk+jNEJfdVjuGcWdQ3p6Ad
TRcDRfJYvhMww5qUC+y4GHnCuBu50OjN/mlqcTVtiGBxhPHTo4LZ/bG0SCd9RxKC
uL9kZ92vU14qL5bVAPyeDJrDEdHpwxcOfFEmE36Fyjrzws9Kw0CmZD2aAozcS5AG
AW0gV8JiSIV9sexrlXWlNEyHxN22WvwUi5TLM4C9yRYzYhf6Ug+Yj5ZCP2xSjLct
zWPvELY47Py9sv9komo5LqZh1mkWS6vy7c32W5j1AMv5WU4jkkq60PqrrESWdwzt
SPBNtp+j6FK9z5HV51U6zDl91cVL0UZDKzsg0pd3AJl39Ggfh7ueymdpu+mrvGa4
5V+u5AwtYLuSOwkYBGW2DAHLFIDkgLCiEyoZCMaXTFGbgdn4NKUH1/wKew/p++hn
SH4xf+DV8z2zQSK6LaChoqAkAuqpqz67qyufwl1vCVtFsryOClLT89BD9exvG9Zo
lApX+LMJFM5BfwluFHCpkDr1TSgCuyMQ5eXz1kwuhCph6uxtVJ/Gb60jMdLOEKSD
eewqCx4YNl1EiGqdtVPaUR6guzflHSOMbOYd5wYC6zoloNHYMa92pcEwAAcXgFYa
gsKQRfX9Pl1KkH2TUlkRRXMieHm0eYY3fvT6Tj2TELQno6tKkwjFtatVZFbHwscT
3zYQwFZ+Mn00rrYv4leHVijGKPYNThjaP2K39VP+ghkUCOnJPURACOr7grScAono
4qSc7drKRrD2h5hjYaigm0Nua0ozUrOs98ysb0IxMv79STLnNstggwW2wfWH8NLQ
B0g6kwOF+QeUFyYiQrQCicxZkOTtTjmRiPplfwYSpRSHbqF+RWVPEuwA1xiZo07z
HXJQAkY7UTx8cA8/kNgc8iPSwDXYTlV3yv0C3XovmkJimC2C+e04a/sxfOgPk1O9
bOrb+BqHg+W77LkqmBWDtKZZqzAG4pDE0pEruSiQFEozBbzv4FdYzzYGJjq9W/Y4
aHpNFa9SxHAQvmupvcpIdlZss1cffZQtgBLgrRDCbaT/FCW7rYXsrcIEgxLsKIHQ
+Dl0sxkTWtp83emdKvSbIQgFH+8z8EQAan+QssOK5aG5p97BHDSPFszB+WClpgot
SNAYpETzB2SkBf/WMSUUB2rINfVliVT8vTU0NI90g+Eq9hfKMWBoW1/YBpiAKZMD
9eLZaF/nBKN0vDN6h7ag/JP/JsV22PVowY0ivKODBu0Tm46dAG+v+o6EI7hXolaj
LJDsGvKDQCQIQF/R9RAwiD0JjIpeGbo/VHOo+e4PBCMKCaQ0EFCbM08Kgyxgl6cT
v4vb392OnanwnChWGasXLe3He1pLK5EvpHbNbS0b5twiGR92QWEt/7Q3RW/0PN+w
gHRgNXuNXU+Zhb6Z/bwr+23KFUbJ++laS70D+vlid1uAXuMaVJA6Nf9c0IjjZ4L4
g3RABqNBe4dLX20EO3oCUxu8a2lApjtSvMt5SyGQAskgE8A/bl/dyzp0ZnNysmVK
iPwpzNf2F6TMsm+m7TeWg9Lb5u9Bhvso4s2HCEowkvKHAJpg96CZVLo4dv2gbi+I
0rIZVmCLNXXxmROqyE5VzHHnF99L8a7Lq1Ks8dgu8zJmf3/Et/eY5tbUrWTDg7Gn
RkFzxbdi7pqNbST6HYKxay1At96VXW+Se+fHG0UEQupxSj1PXd7eZLY3Bzg8ucFQ
g1sVLmOOsGdEnrQCPe6yVWzkbMS4RBCxbRXSaLSLt1yVb1IdzP8C3QcOfeiuO8a+
RBOiyBhWCDhVaSgBXdbtXKEf0Kgj++HAjAep+s3RaTpuK2LGR/jn99U1vDbgythW
GYH3BAltwcG82/LRY/63Evtf0n0i+Dc7a0SwN1H+uY+IZnvlvCxV9TUQlns40zrl
heDMxFkloLEOPPHHLd6MqVAgXfzLBn+WxC8OLKfsIJGxBVSe5I8hIjGwFV/qYufb
LjjhZRPxcRaVH02aNGjjwJVKRV0tE8gGGw7vruUya/BxG6lQ0R2XIfv5PXcW2AYx
CWlg/NeQLNl+S435xmIhCFKRWyOO6y8hGsTInPDDtwVWxSaDUkR4MK8YUF04ZD67
ANcHCpzAJ4tEJsa73Mbkx8zVvVeqyd/JncwgAAf7JoAKa6BuUaoMCeRxOFl62/7b
+CKET9Wbh1irAsDQG4xSbnDrWjCZn1vD2AsnDC5GKh1uLhjBnnV3ZuH0nt/tAkHt
9+pH0Vh2PjfIbsCtXZgYfq7UMkQWpWD1dTewcMx1CBdqaOcmTZR4GUTEaWpAMAOt
yWxvFaOj5GmRsrRNrk4BhjAjCHV3M/WxCwKqUCr54pHyfOIKbhuT4wKFiFxwS9ni
ljsfIX8G71XRRYkH9HA6zhCs50Z8tp0KHGQO6JzJ3ZQ4ZN01KbZW5SaTZxR8Dhlc
19ViIqFQ+wTkLRX/r/xP/z7pkvSeFLmUozaITWoQ5L09toIOFh6uL63GMzyeOX3h
VVLNrbaZpbbKw7wB2SsvVcpd/rP4zWQY3LwVht0Aa3k6isliPZPHiDqbC5NtCA/0
mKgBRsMv5b4N8TKdDjjQamtMZ8ETSNaAASpIcC18LyocdBL/OHZ8ti138MgMy11u
r13f7XGqpRoFWNijYi+kjCAoQ52ObthED7rvJ+m8T6Wvzc1qp8OG6h3rdXKXAbpp
PunY9JUMfgrbg+pYF1ip/elenbsSzqJ7gZSaL0Iz7+8C9z+EWSfj3VTolV7ZN+UX
Wd7Odxlx+7GMbBoC0RfTtVbiq050ZR2KFMEMvDAiRaQOWPSazup6iUNGAg23nDrr
VHuYNjRd14Cn2Br8ZxYb7YFEmFCNnoXnPwyUfgUDzm0cc/kuUQEjV5kxbbAyDvD+
DkhSxMKcSVeb9rUzrR3Po1gRbr2J5C5zUgrXvxoCsJtcWVa2fcqgj4WSJbE6UhOq
5DFJGYueV5izkMIM0EOV0WMgaiE8YM+LaXv/BdaD1Xy10g448rz6UPFfyUx9grxA
zxo10dYO80OqSUGZMRvKuHxET883SV26NVKY9+1k4v0ionGzhGBeZRg7UdUpctal
ECKRTzrNrNQhZlhp8Au8OdcejOEvgbp7FsiwoGj5uFWHv7rlasLXNX1VGqcAdPWF
4B0d4cEMRUgshtAiWyi7mtBm7DKVXvEnB5FMq79Ou2iNh6BYwy3dR0+HhscI78k0
YadSs9AsSv2SoAGm6c/TWzzi6F7m728WbPdMj85Cr1xhFiVtw9NYuQxCebGgdRm5
kbBEkZGTCODMz+/p0eV3esKXJK1BTPdXN+FEpoYiagS+nq/bQcA0mdUgHBiYOX2Z
BomH3wEeA3XgYEUeE/xVF94wsVdj7MTRvPDac75A3+QgR2w5Go623z/Uys1lrCE4
cS5GSDg5zXSucRlCvNRAxOLXqhMcoxGdEPTMVvO6ElAf6kqe9SwxALw5HTkPMpLu
pvgf40fKM/xq7K5f6PoVZDLI5hapLGipfAQX9noYPXTV20NG0pXBKmYewlvgzWtg
EOdjah5G0AsqbiCY93RFYQV25rRXMVta9uUPuRXtFfREp/DNSRUmJz2OBFdzf7ML
6BgzE1GdZjmPCDO/lWYO7IN0fDPMwqzyuE2EYp1NMsK3jZp5l36VabWsn1PPJRQ2
H4XzjxjfJEDYhuaS5cCG+u6wO8Qv+Uo8htzfIYUU0ocP+4PXzjVDkpiV7NYgYHvJ
w6kh/dknX+UUD+IG+q+bROGu+rt13hfOK0V9flHoH/CSjbA98nYbV8o6zv+SjKry
bxRULO4liVGxFsWgza+/ONIe7Qvh4L3eSzTjjs5O0Ruf4UAUJcz7ICbQgJi3PGSK
EJ34Ho89CZ62w5ubRmI8Rpjy641tjnV8CJBCQZAeTQs0+gGEE8E13vQXCbJLsXJr
MnG7di7UKjzzDiu6INuKlmMfGOQ+rh/gKlPXRR2Cui32Tf6qJJZReLJvnocUmOk1
Iz7Vn6c53nnV57JqQaW520gOo3kShCIh/6Js4fLUEwdarLcqnaBIUmGNbUp6fa4I
Rl+KkfkwToNVWqPargLgapMTNJJnJwaQzp8HSmJetPal1e8w70xTPtfc64tWkMz1
d7R49yn7LXcC3ITOJRaII74JfT9CwIRpUmnVbWZldrwzz731ubaxu1z+Odw7akFa
92gwpi3OmIhnAHpUGBfJ72fF3xYfDSKhhdwxft99TNQYeM6YaoEcHblDU9Jd9oZg
J57ISZ1WUo4DpbakJ3YqqWiEUhiE3ElqlxKPPHxyMWSoWQl4WHfFKM8T+zwMg4Z4
mFRPdtWTC0qKUhLdJV75jML+4mRD/D92vQ3PQFkpOtGrxqTJNlFLBcjjAPfY0uY+
f4tfjC+C2sS57tuFZfSRgbDUu8+CCHD6ID61kPCXFPG0IlPR5Xj+M3c/jhIH8HB7
VJK1AedaEhVxgjzbYin4t2OHjw6kgAWnwAY41V/SaB3+2BrIUCGQTeCRt8Sabgv7
QkOFqzmEoRzH9D5RPDcfFahiRlicry5Qmrh1UjKUduYKHjWU8QUtS0iIDfib7uEf
FkBD3aeWfJIZrDRV0YZwDCO+W88M1ZoJr++NLboNJauqtRxcI/R1gDUqKdzVFz52
HZdbszCsXklQ2Y7KIyMUYwzjqqyHWBquLtQGfJzmc9yURzfsX/4ay3t+aCQgNyiL
BOCSAKwH+kQozpO4B4STz8EQc1dXMag/tbEsZinLd9vR9HLCnQS/b54dkQKppkrs
ncFaLtDqKxiOdXVjk1AQ0x8fiNiIOwr0rT9ePqA+UbGparT4U7qXEUHGMtcCXvsi
clyD07+RXHGircWQWxa/16gf5tROWJlzPvwFhauQTk1F4C/LtaHYx7jDDSofW508
HMoqkbiYADshPAxOV35yIQs6mnAeiFWLB07IwJfvHg5a1zH1tRs/6K64Rapw0f+i
oA+piqdNrCI+H9QLbWCXplcpGs0pavqvigQyJFOLBMIzTXXN/61M7+/W2NSiF18A
JhWjIKla64iyHa7wSORSENIfDaWuksG6yjId8avyp0eCyBw+59jddRgC0csSa/Yo
+p1Hmry0ctzHY5ond9PRYFZdeJuaWK8DwxwA9tikn/frlMFrkXRfCQ3wEv+EXeMl
wF4HQo6D84CVBETaDJ+wLVc2/MxM5zG+fOxqtn7SHl448Cjjtl7pT3w9ni+rrEDG
q28NIQmuI81536RzpzUrk11jAFaMjrXs1+QjtzpN6NKQs37M2uQfri0UUH1IbI98
pgLPdDi4US6A6Flnoan09S2vmqyt+5KfTKT7AcuMtCcm9Zs/WW8XJSUCCTavLuw4
bO367I6nlyno3gAPdqSpJ0uPPa/uWjwQ9IBnwoCFzmdL8v97RMZp5so/nxkFjqhG
khcIe05S1mimDHaAtV2O0KwDiz1jcgowOHthaoRXnJsgCHx+CTek2Cy2TnIzwgJf
VH+WC39xz3Iu2Vhidg3QDB8C/miWcbNGzw/ek3PKSAl61e/jXnxItmm7FsqfHPUJ
E5nCAVFMjuSqz4nwPrroK49SticgaDL7qAqhWTYEcdTPN1qQvy07V477XFJEul72
4N7SlUFpFyPoRSL4JWeM/ytZegKFDIQgxMu9YFlzPfBAjJM9mYhuw9QzbZC3O7HV
ulNyw5/K3RJq0EOQzqwjdLrJjqA2l2/OlMnZU/pHXIPcUKEc3ySubauAf9sriucg
Y0mBiI6N2tftD4Ec8FBDe0j+ulJNN40UQfCFaSpaV8Al5WuA+EdfZqUggTs4EBFu
pawFsbPmzkJGImzX4WMnE338KOriD24jjS4xU4yoIbo819erf1PGgymYU+JgG2wK
Plk4ue9HcN/+19j0GMrnWs2pniKDI7G3vaz0tE49fhwhwTa4M/MLyYxv9l7pfkIT
vIMZ3su/ePGMDqGm+dhv6BVlQ2gxpWRpcNk64YSf4OUhRjY3iRV0fWoE1U9aYwis
WposeKaZ/XU4wBf8QAsAP+eoWj5Qi9YQUbYSO0kMF0I5r/B1U0ImxO2gHVsrEDZZ
sF0lQJc0IaHhjvAEyBrdn775hiBE0MZFKPwjTMJ70exDygnrZjWHE9qVgQ4Tvcew
BzVMzCaxicDkDE0FFandFndbirbLKE7VJkD9ad+vu5/v0TOz5ofaf/x8pQkpn7OD
mlE2epBSNithyWlIut+qTUPzbJrTq7VapTjqPBbfkxYaovvP0LFHGzMFx1kOH5TF
MHy906w8PzdvhEiEQRbP6bLZDp1xNeMUzYny0W9Qrl0pqfvGX/xprDe12sXfomYX
gew6Ul2Ny6ehpjZVrETsX8yMDPKdyNkA+F06ZgeATztzykogRV3K+OMgmd85+s8V
4R8NWTxQUETYjvMqBhzHaV8YBvmhf7Gdewbu3IwehM5lqS7JUvsU1wHZJbcTP2pj
qAu6Ul0+MM8bMVXnxeIUIdMhUF/tLWD/Ftq3ye8yomq4dYRReEzf+V6fatBEZMTW
+uQcfF/3idP4X5EgyazCpps8VmEeo5rERzyq9eog1U8vvRLqYBX6tsadJM1A+0hQ
o4ZajrUC0UnV88L9UhCY9vGcY4IV43fzUtHjOF+tEWUenewrG9Q+cHzU+kQeSwKQ
MyI2LGBBVCrc/66hKd1grPhy7wMWKpd7lxI8sOu21Yx9RHM2No5g0r6TLjJ7ZYBF
Ow2Tjy+tJKTLzywZOxKNG+Kal6y4AIZxFZpLAktkjBpkXt8XNwVfnyQxkTYWuZoU
OxiumcS/XwOJeREtgsNWEMYqrlnpx5ys7bN27lGt98gLEZZBKyvpPDgjQAP7/dFt
W3jQkO2Q9kzb+eNa4G1D4PurM+jGclhxiTC9o85lsKrZ6E1EDHaADFISDNNPpPL4
8Sgog/BiQ8sKJi+qh/nFjnj3O3ToSKGFbcJk7UTJQkeesa4wInAvrYaKneYVluY2
+n3cJtcuL/QSZsaCeGNhEsXT5+xY+LyIxJwo1JcljGY64aesrEV4bjZULRqKnRhv
oIQKvH81VyjX+1RFqKPOi8nRVNMFl7Jtky+AZ0mOWtWjTZ1SRF7nXmodrtvf4nP9
DKfZFLI97elAItPlwIeAVnAEDP3wwuEADcdXPAuZKqGt0U60GGuJG9DZm66AHqU4
1XVMVtyAJGxmghQn63cgm9w8Bvz1K7Y+HM+iiPx3MStCNvtJiNUwJr4PAy0YBSlZ
kD4plT2WIHjxpzP+TWzaAAFV1x4hpMkcU0FDWhVrmGOJV0X2oavYT4YTa3QhM2nI
q3v4/tua0j3ml3TMmBUjGNOhMuPLeweuV5Zs4sdcioFFWETosub9uqqc3hmII1DS
rKTw8LfYyan9Xr7MJI6YfjKWJ/GyHECnQZhEfawHAJ6u2q16AqjAPER+uf2tzZbl
SvGJzEMON1TLuvg+uIacJL+6cXkqLiWbJFcnfvRKuFhIHWsBG3UF3Gkjo5A74CnG
NYW8Mk/0suJ7IzeZBa8XAefSsiZU+IY5fnocciLWGLjRkXJeIbtj42MzpKfJuHOf
EjAEbi9svGe9tWe7prveqQeLszFnYhvuKquyqdYHjuicwMIXyC5Cn4kgi9OGR+g4
uRYz+7xaEqdRTGmhfp9QSh+toS9tXQ3DQGxAWw4GdVRHFVdw/ZoX7rs+z2VReRpe
vRVjipw3t+EzuZ/koTngP+XQfEip7W3xEqjaYqMJ+P8n7Gm3drOd3a2DAmiacfrF
ocPtX65mw3fC8MrX0TuE7lEvs7tW3OG4EhlTiaf0QCh4pkZ1lTtGBpeyfeXlvFxh
51bwqo5klcWnSw3U1x1YhHW2ogNE03c1Q/BgmQPaJdJ0UPXrkMUVyN7vf1tfMkkd
EiiSKRdjR2XURZM+yJ/HvLkz9XuQo/7g3Cczvm4NtUta3jnDTyYJVS5E0bfqPmrV
9flfr1i6gKVVZN3C+YreuWSGqeC8XiC2IW9nXZqjBSq5mMRu9Yh8esob2eKf7tb5
kkqWor7qvNPF4i0aeYxjVwwIPOAOFf3P69DwSHXFrSJkaSCE+nksrYza/HOC+iuu
/svjY06npbuTIm+3pvQTkeeyvOQ5AV8216vJaSeQeN6c87gnCjy6Etx8a993Bn9+
CeZBErk2C3VHXZE1iJsyHumtwICBOaoTwqMDofaG7/l6J2ivH50FrbBLO8sdqY/p
N809m3vTxZXfmTvIfQXXGjj24fSnjBImtjmuHoqxYp/t8qaF4NkSsSSJ45qAduo5
ggWwfwGILUBb8WHh1EvSHXeDgRz+4NfPaG8Ed02md57ULB0HefseRrtFNZJNNQCf
4apWwESJ6llKIGcpMMI6+nZZ5vACKDeC4LCFWlPMhQaTLGKyuw7aEFwnt1ZBDGnG
I3nLPcyJhgdMf6zovSlorshuJNJnhraKmX25ziZqo3wOmfqri4WfOvMzYX4Sa+Kl
SjQheep7igjQWrabIpDUaCKeiusYNEQ88/TnTjvYdmQuVY/MGz5uAmdl/aTfcYRu
59wjw538k0zpJ/gvAVzp3/svEws20yL8JMRvm926NwY0prihx3KQ6ByXJDAxqoPc
rJjtEBUx4GDpQ8+JZ53hOGEDlLRLlY0elc/vFmrukp60Q2qaBJ5vXaUA73kplpq+
auhQpgeUD4NiKSeE8CfUjDRdwmx6lAqgRrhqsDuJ+sdsALJt5BifKviafSf1wqsu
Q+hT5++MafF/WXifCQ1FqY69dOgqK5B7Z1TZaJQ2vzRf/Exnjq8w5HXQ9W1aAOMJ
JIhna5N0qTMQ+8rI3CvK2cy2+zZOven6vwd134wsA2M2iG5hqhcCIHFXQTl9WVgT
2TFSvZWY01APQujAmXMTsPYa+RVykLLzFbE43NKx/QmOd3esTRyKBIjh6tlY55wK
YlB/BNDGOZtOqJRO12btLtjF/3SqmFF96AjPy9OcZNJbegpunWLRPZTxz1t+ypzr
vMfhamvdbj6n8eRndWFP8ndFuS+OU3hxdAZ8Y1d1fAn3VEVmSBfzqsbue2cPKqHj
Yk51ZXhpK/Nu6JcUFXhwHjtHbLamYnBUINPX+tUkrONXriXILSAtfpLfweRbsc/0
ZE/9u5sOhXktVtkBvJLtdmVgMdw9votlym9bRDQF5ongb29RMVlNdTDcfOEvGxhR
3OluxafsXjkAmmkpinvXKD/nR/R38wxrFRAivE/OWeATVsxo174kBCRvOepLcpN/
3ORIMUxswgIZJCCp9050iFW7qoX6a3sUzF2sKz3PLE1bwiHCCEmX3+LrS7ukIYlu
BBvSkKZOJrfU2ZxdXnzMGvbIEl2nTzGwa/jjx/srDepwXyIUvUTqE0Nyh71u6gRw
erBh2buSizwdOts0dCtU8HHApjcB2fX8X+gG14TJqeP15L/PJApf3OFsgCLuwFdP
HKt/TO16X2e+/AFQSSKnUi6pysbqAEEc/RsdudEkkYwy30+uubaL7NsH8AM89doG
SiscENfk5PSd5DfehUHqsTShTej2BA7d+i1a+rYt6PtATUGRotb0tt6e+8Q7o7LO
6mnI5X/yXynvEW7/iPikSs+EDbKHcoUHvr42sSa8reH2Zmx+b9mX0yzW8yYGsN35
UN26TcN4M0YTBMLoO5HHnGWX/cePo+4PrraNp3g+UqjwaOgUMn2fauz7Q8F920wQ
z7vb0C8YqVz9aXyGuCT3NsjZzfC08juRTAzvuhhalUSSeI5K/5iHGtKsjvBu/Ond
yJYAkw5tPDgEzivj3XXkMyD+lbxjzCG3FB8aWpJz4c+3fOy44aGnVwDD+OeEKgbJ
7Ccfd38xcLCDGThmPMsguoI1GXbQvhc+sR2sf/Pby7XSR5/xOfnSvr2eqUs3HWP2
tXLVT5E8LzzpSFULH6Pk8RIYaxCcej14rdKGDZ6erMHLyBYw8NFFpnyFI1fPcXHH
0v5SN4FSYoE71jpcr66uT8HqOfdIUooSW2KAt3QxC7TyoqsxUCPbKgui/wCojs7q
Ev3L6MyCwyE8aCP22sKL9AKSHNwUhHnEfzwEQXQ0lq1ZRFIca6DLtm7+b9tozUjy
69WLa9ogw71e34Ll0O2aWR1HbAyYDtWDfsI1FTw4NO0gdS2kY4I5V5WaFzyDkchQ
E+yWAoS8cbR1Rt8tjLjIz+ZrY7imlNWJYozbq+tA/fOBX2LtS2qllCxkti4+/wRv
/m2qwx3SlOOZQ9TuDxPclDGVAg0tzjInljqYKkdxGRyf4fs3ondF8u/azOd95KA5
qaCEzuK3apwHbIdfN7gBbbX7YZbVk9EDNqB8U+Td1HkL1XrCnhCKoVo9ULNGbIHs
srId1DXgLLPZekVMY1T7xsVoLlJQVSsLdBaS/g2N5g8=
>>>>>>> main
`protect end_protected