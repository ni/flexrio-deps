`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 38064 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0gQgIG1mJzulW1XOK5NnZR8
C8XqDUtXW7uOWTnSVqbIbkDFuPnBV/bx8mCbCZD8vgSrhU6d91HXsMBCmR7AJZPW
JoUqWq+aH61aUGi4mwNo0uBMdtaw3U3beyeZ6gdat9gb9FLNxygjHbyfDg60cvLn
Plajsdvv2WzPXrv+sO3wZRvwj+HA+HDiVDB8AYEElIURz3TizWT0lmzfthW2s9Pz
4W6wxdCgbgr/egJEaEbfEMhiNXtTCL182PtUZePyzdwnxYSO7IFhwv9KooaSPYPs
nPO9qRZASJzMnMV1XR6wjXRXFNRr4lt0zqF2qu9aDFnFeBZNLAqsQAyKb7uRBIs3
QokUjwQGcw05gvD8K3QjgD6eRtfbqOWiu1xjjxF0A4AbtbrBE81X2zDf/rmVbQP0
rMf6d+4F7957VOMw5ZtLMAlnHbSkbWBGkStLsS/Z7Ny3qoKK7x+WyHBeRlMVqqVJ
bI5y1RVo3KMbKgz2FerakXaGTEEaa3o0NZVYid9HnMLUFpbA0VlF3rS6aStWMpQl
oH+L4ZGbTsw37hVL3Ra7RMUiAvp5wnwqZaDd7Ccyhqoiha+NBZvn897hi4PkJqz6
sr9DNpDcXcV+b5+sJU5qg+IdAAFt7srjdMtQD8h1ALyFcaww4EUovTABwpE0kokj
x5ylFMPbGNE90Au5sCDhnxbcTvpwctQ1dpjpS4vh5vvojc3qg3j8/IyrGVHM+NeH
wN13bgRxT3b4nfBYTJj0KzwMbWMjh2RxK5yoes3knUxyUa5UXtRi8hJ2FNX5d5WX
8G69P+WN+IVHfxx7lRU9XletieEiZcIhbEyd/8I1jIG0vXhRWpT8vVTLMYuR9otz
C8nBdPKrCnnvr827CRO5rqHJ5DyGtneEOu2RKpks2L4a6c8nzj81rkott73Uv5Yw
0wL51CRoY5ty2DW3pHPPlIj/0RyU+9N4QNZVD0xxgGwb6+HubcMxSzx/Y93s3wbR
UsswS38uUIAPqJMyByDOEp0Z0SKbZTQRj6NcfQ56hA3FkO/fv3bRSVdwxqpxml9i
kOzBaHda3YkkHzGCJ6b2XhFr9JMG8xHWFiWDrnmPaTjbQhMRjEhWZhnm/QpOWCM6
WRbDNERWkyQ42SAxvD5DeP2m6lQ1iFhX1Sd0mGswqfChzCOQmRqv6fMnRjQvkpiT
XVmh8oI5C0x0SMs9TVC/fq1tXYTYxz6WH/o4k08rlpxAY61yhU8z1FfT2c8fH0hH
lQ3lTsjAVxEnON0MkADFqLThp8W5fXFLVEPtEmDOyiTPv+rGDZd9TCCotkh7eIv8
jQfYFR7JtwDXglfsA9ysngI6rxhnOOzsazcop7o1aHITypITpFpXpYSMhS8qAsrP
V9VezOPvzO60Jz2GOh0+3BTc13P0iR93/AV8PQ54Hpd28gZdVm7e8J28aDMsF26T
HYK28E5DC68xocvb5lyprnUl3fqUJgV94EMp5unSor0GqX7tKz9zVGVt1fnQoia2
A7Pur5AkT8zj48l/GslVzh3HuSeayeaAdZ1DDFi4A9uHbQky7uBKITZxEiAIxeQO
hWC2OurwxG/K5tSTAnClYqlLByWyOidPjTjiFqAYvwYdtdWY6bS1PB62IcvE+6Jr
QlbQxq4DVdt62ZGHQshHXfXi9BGegfS9e1fuumKCrej91VCRS/l9ijQtdbK9uQ1N
eQqCtsIv6fRH08qYixOfZdZWxV65ptntZEOdsnO4iiGTKFRcxEhhXShfBv5J3Q6d
CuIHZyZAE9GIcnJL3/2890+JIAwsbzZJfl//F2xBhajQV7VBIy09Hr1xM4fKdZgM
uy4EZgtTKsdWyhjkbarhsWFx6/2pju9rh5Rw9PVVwU8b2CXdCZQLgB+OmS/2NKeU
eXQHx9nOmLnLBQlBV5Aj1+m9Im7lddB+TmXRYbVSylCkXqWOdgZTYaOdBHdch6L5
tSc/1SNedTvwHuzCIwSz9xoVP+HKTsaqNAX9878vHQ6pQN4/nSO7QBznlH0PSxbu
UViUY2F+v0DQ4kkF0+v6ImJudfMpHIeswHXbYJFAmEqo/gfZVq/dv+rLVODab8wc
MjZBUj0drQ8Ac9+oNFD8E59EcGRp6FedpIjxjs762QZx6IOj4D8ZuHlgM2IKy1dy
2NNDqhLLaCeIHNHutd1r+SMIjtMIXgPXcp+1JVyUfbu54EveAoliHHNT5rSELMdd
kszm027Ht9hMlwi/annXGr6td+xRfo2XCHBe+RmaVsDZsWN4lufrH/ZVeBAe2EQk
8FACGS6NOJ6ZR6aUtGlqSWgtmwa0+OT3ubsmlGGsyi1041FstEapc7XAOYxXR1Nk
7V49SRmgWK7HQoH0T0G8d/Lezmy99ZsFg6CCzOm9vnIqNmOWq9lPJ60A9yzfyk15
S4o1UouZ+eg0uEf03Z5cbdCLnTvIEP+7i2hn4ESgXsXh1/cgA/O8iKnLjVtd0WWm
UwoQJLEqrEo7wTdz8sjquKc4r6P1/DHLOD7CtIpGiUG0EYnwGa2lfpZE1E8NcOS3
SR1Q7D6+csoNGEVm8TiXwMvse8Iiv4MnVgHmcKp6EeQokyHj0wdHPBJgV5NfJu1R
W5uFywWVIEhZ94J1yspJEBysRR9TxwXaDxETH7l4ZD+x2mbeMxUV0GZILJxgqWHd
JGv/71ANK5NC2HWwurO9cVjFjnr1BiwwIzyJ60O/fZc5U7RlgmCQse41u/Hx4crE
e78TyVisaQCQPk9/pnv5Cn30Mt6cUEilCzKnt7QieX8PFeIqroq40fUO8mFEO77Y
zRVl7XlUwiqDOjY4UUoMQJNpvcDa6iEmId7dAZHia5VgYA7dTjybb14uI2qHYOIc
3s80krAg6xs6fmkUimcQGIKMACXb8IUUXQ0LOD/jeqp2UjJUDWiexJE2KvRC5IGX
R/MwTZkxD8sqy3Mp68BksxNJbpln6s/nnnuxq3W3vqKAdHdXFBfxVgHzheSWnjc3
QFg1Ar5Xvczs8Th0M4mX7FC8kbZIZw/ABbwAKS21eVRSfAtoFlJauYB5LKAHv2XH
3uoBR3ViID4cPIgTaUt3nklebCFPaeN2yGsB1fsZmcNtYLbEVCnRw0WUlny8tVID
hLFuOs4/6rYW9irsAuHlNWnsqiOZbYKDTL+2TcBJVv+l6PJkGcimtO/AJyuD7S3x
oYu7DeKaDymTBBl8nmAQJHTwijHVwCI+C0lByo7aKOMnyTBxviERu3LyZmGLT0PB
+4UOp8i2erRxib7+dnR3Nm0rom02/paZODJsPk/IuZCsC4gRWZ6cOUxdSYM8LNQt
HEvvpQn3MHLLuI3BSjXwe+PRGiP7Ud7do6Qm5Yj89RsV0P4F48ohgpcEeJmgqdTa
5WKRGbOphL0PqUOGebrWRa3ATQojxn3iV3LD17U9ORU/d3J9DBUtGYhif4WLDaDY
gV7sv8vtOVjnnokFOWTnp10FVER1cbqmhALwV6qxi9YNM8wVwzSa7uaV0hUxoZSW
fmvseDxZ5yj+dEDSdHblC4fQ71U38gWaMlfLpgcR3DWhw8TuPhq4yyJFWwydIjtj
od180y73EgrbDHGeB/1DxPrn8M5coOnolPrVHpOoewJ/AocpUbywapb0UCoinKTW
ZgF+f8QqG44/z1rrY3NXJEPz8F9AJS8fkQs8hSxfAj4NIke5ERCYjezWfMbduHjb
0MiZ5CZ9WGUDDxeN+qh9dDe6iyIER8x3aHlhej2VZK+SctD44n299f2sPkcTBkOk
wNwWV8k7wzl3kmSe+LOeiNaRbsquMlHDhv9am+KkOOGEFlo1EOZyWdc9GVx+VFwW
29I7CdgC/GBwgjPwApPSmGuuiltPqVFHkPD+ZWO1awA0nRN1lBrquSfDZkz/sQov
0QRl3kN4bgWsEj8F/U3eTbg1gbR0q3fyM3G6B4FAvIRfRCCPX0GwDB1Cwxo7y1Ma
+mSESPaFut5Rto5y3/o5Nfp6rKmVGseMfoN3D4eLxYESNtZdT1hhxqOjpIKZ8B+/
52PInNTHsiz1CyQOIoSSBSARhjpd9IE+P56iUvsqPO8N3xLpNaK9r5NHg/TFnYck
OrM1snWvveUcgB1lC8mF6DwvojpqPJ9cuWC3nYc4qeSF9V3drqE135Qxj5J+x9sw
KNPn85bK8xt00EsE7XU5PNj0Y8AtVhFeES13EuSldq8icV0GXljAGdFLtVMeW/+l
YJMywClUtwjPJuY67H8OepGWGSJwVWTaQtZvvvxrWbJ9NwH2T3kPgkTSHs6z5LNC
Aoaw5CCfYwzFrhGr9pbTbGl0Zfn8tIc5Ekeav8a/FeTew1fItBnFG+eNJAMBiaVK
Uf0a68xaofXf/zDOdQEaEN15/VHsAzPRR2N9BApqULY3zt/O8HklQMR1m+arWokg
jjIceHmqNN0EVIBco9ma+39Oo3K6+1LCebqMAZbyiPbpXA84O18ZSSda15O3+8Nm
ybWrpF4GwohDb64RR8bDMecqkS6KO5sde4JPNehUbjMezO4wbJUc7iYBd814BMGT
Zn0TN3VzQe2jFoY+gmhLn3Kv7STEHvpugEn3ka29bJJn6CQQf99dyuZGEHYrLthr
n9zxuEAkZEKJr2BIv/V+5wASfsPEmp6soEFo62ZXTSqlhVtqEjaGLKexXUBburEG
cRhUiOqzwm5TDYCx9BsWVkYLBJJubljDvsiE3yIDxyb+NqUb7uQAoKnX+7mQd3jk
5jZGqpsjPchRyAK1zyBUp/7+Y+YFPJU1x9kT9psHpLHq5hQZe+jny3Gma8tAFTSY
+pbBKGk0+koexmjmP/HgzlUe5+geHT5wlzD8skLXeAf6B13KLE+RBRF80PnX4w6A
qe1xEUKAb3v5Bb3UmnQuJR/sEe1rvIdmsL8yNcgXRKlITI/WXtk0ob0ZPGRj6CNV
PHdVkzj9cRM8Zs3V9279mJUKlJ2zZJ77DgdFKM/L8op5pwkVRQZC1F2oeqdXrHpJ
miwyYLC/UrQo3KYY/56vROcT5Sgd+cIm1y9GPP0cnmIQphSXKKxXhbJlA5veiyb1
m7DBsuMQy3m4BwTsyUHplnKgnRp7C0AY+bgJz7kyrvhJbViPy1cCUVwbxeGyACIK
MwGuyP0RJmhkEukXgjAUbXwi8yescp5nH+mmDygrmDsnsRNmqIhdEjs9qZQJ2jSr
ogBkuLqfVZwih3H1a5gXTQyEoxgXjCbMAnUrCrOoZ8wp2NNlSU5anE5Pw6OgKMny
RGzciCQqkD7Zb333qz+1SKlBSPKn41FcEwqFwDYHcwPNA9KQZ6Qu1YkVddsrj4VA
jD2gvpvDvwGU/q734FvKsIhZNuusyCTy7L1id+0HJoI55rRojBlVtmtq0KweiY1X
dlxd91GpHQDOnaNIZFxBhcJD8oIXQlX0CGagN32O+ME+ZC7LjsJt05ua6W5rkmEA
GgA3nI4PLGYUi8GM0U2lRnUVKdvWnXm+979fXnZ3zIKeeux4S1i6njBYcSaZ9S1B
1L9NjOSCCBJM2HuVJryxKKiNCOP7LMXJV1HOpifa4Rwz5jeq38NBW3i27ERhdXmL
hirD2Km1+eYcDP2RbfC2Ie1gr3krvrZTSbDdJ46LH7i28nxoNTKlXDWcfpCILF9+
y88z5dPZc+GZ8thu+yTvR3GrCosSslsRrboOLqtrZ2/hlgkY8urH8hTSEPDK4YyY
P+McJEWMYU/eu8fyLutQ1LydONPQnzD3RybjSNxliHpZt8v0D1Q1Nei3OOLuf3fg
MvfsKgbXVVHeDJx/WjIPVBTYlzSZqis4jhhXd6rz40p3v5qEFUiqTgKY/UzeEbOS
aMjgjFrZ6ZP7MGcnKJSJ1r9x1liEn1K75KfkJbWXPAHies51BU+InQk+JbCfTOaK
84DbkR/fgAd9IIA/MMCY7DzvaNra0RDCGr2iZPjjmuME7ogLkuyyeE0MExWFqZKN
H1AFrUoJnyv0VS832N/u5ikjakij3MZqBrlpeZA7IUrjXfshHMcivHSai39/3k4T
R0g4PSnQzpgtdKJoHCk8/jpz0KIpuCNcba6/TfHNLM6VsBd1VM/94Lgf14o8VLr7
c+ykA76xwbWCM3iVGet3tVQYTgQOQgji/9Yhb+YHwa2cUolcBFFHCh/bxCH4FiKM
vGl11mQjNAKSVYvYdbiDKQRsp1lKuG/7XCOC2RBoHEqI+6wDdNLovtE/lnRo9Rs9
ItoMPszbvLgC8jwT2GZj8AyNNxGNM0gCAMlM9loE+rR/WZ74SbDc0kqROd1p5gPl
90XmLipgqDH2A2YvdKYHucE21A0bHwAFcjXoQ2CjlqYG//FTwdLN/WZyNMN3ge7U
gp+GB5O2CQAB1XYHtI3FeN+LDZOsQOcdx+aNX/KE/IsroaKCv5ycQJHtjIrAmUfs
TKYUCOIqXJItSFgqWQD14r40k11tIJID0Yi0kvfOhHz7k4KRe1NmkXR/mx2ez6fV
r7QEcMSjoe4D37FukH5SMFI8kcgXAS8P10NCk4D6M1iZwIIiQwzFdWxx3keh0W7B
3noULvOU/m8t1/p5d+e0Tdvk8jRqQTtxEznc6I8jhkq/WULQrirf7A+si0uFpsyM
b4WrDQhvqVeRYoUrQeVQnZidC4tM0KtFqREeS+P29on00x2+ti8NzkoT2GHdNp/G
VYKhWkKf24SNhoVkA+73PAy+mX1APJIDg7FPazfBgE7I2PxzoWdXGreGbVwCu5V4
bczBrpTEDBlg27hNvD2nEADsfownmL8qzkMzAl1GSXBYxCN527qD/UeqSLFvBVvr
3RXYXEmR8oCq7GR/BZtewzL3orhNaHtXVs0NFd6qheOC+hwOHPzgfQz+zRLqjaLN
zil8aZWna2XCStahVVX7VCBSSepMGz4fqa7sHvhaS6wsPuYGnfV+Rm2RhGfDKti7
cndDEmvM/zFRU+gdx2lJGmx0dUybpvezTxQaa0xQ3rgXMs1hc43EN5SneYM7fxWY
fgrsCU1k1AP0Y+Ohnsge6Z++HPiI6KRjfuEk8tNhgjsv43RoF5EywTnLaMxDIlUf
E47Q7yMujTvKFQITL2lfoCJ+XXTUM3tsrEPmgiTAl1L//fvSWc8hes4hoSZ+Bfyd
MdOJkn4OamOSJU+PVAoevCXrYlM2jCdtMai8hzaovY4yyIdKjC1YG9Bx51aPsOu3
R2nihKaFvLF8b7P4UnNr0EW2GEfDHweEgdvmKzg9pR+LjPFW3PiLKTGxl8QIl4gG
vSjjE/zhUzJ4XnWPohXb02GLt5obxLeX6i1/6cpiPPwpKUeQlZZKfB3kcMoR+5IM
s01dJp/HCm0EjiAU+Ebswtb0qbAnLyvRCLphNIK44Z+SUdy0lx318okLYBUxI/6t
l0GeS5FgeqqBhy34Ke1AfR8lKrcbNZmbX+GGrSkM/UyIHW1NLFXTer1P3CtJDbMZ
UKcgr0NJrzjXFzr0Fn5X3WjELAB8vVnI28Wba2L/NdvkmtibLkFaPhrcPb+qbRqN
sKAFxR3EZhzVZ13uauRikcplhjuDByE3fq4aOvdAQu9/z1V0G0xkSSPgXuLeJBgD
wE99MQZv56eJsHM2iY5ZBCiX1tyL+PUAmNL+cJ5hG1mYgzjl0mhpyZE9Na4tClRk
ehASF9ZgrWk2YcHT0RPqAscRlXR+aT4vTB2UnxvZ0jN2izUVt9VtZU5/+HjOQJuD
MV2LE4a0Xp8xnk5EMGqQeGdlNduuIWq4xdHZNWoWjRMyevWST6kR6UJFqWRxIiTZ
nn3AOvZMPqEjUm8rAoLkrvRCPIOHY1oodNS0bxrwIOTwUHLmo5/PbVcF/kqeYE+k
zA8NnwdbSp0v5Q3R8zGKP1kLX3dgwzhoGwVMKb2UtUAWl1YrJIrZXdlN4evxCORB
LVoXQ0lahOPsW9blijNiIeI50fEd7Rb23/TwO6kWtIoIxo8R1XT9j+SGEWNMW6/i
AH3qpUjl/Yn+1QkjHOvSoUuBRAEmfNGfMWwFdXqhd6FDl+DpHQogNAqy+2bMBp14
EdidqVX1+Hdh58RKt38TkrWBYjFO+IvTPJiQCkCStnCp1TqkJCul7F5pzWbh+XZk
ak/TuXyAbVHrn+TBUDiUFWRasS1EboIeNy5JrbxdKRKWD1GWvqxI39TcawjEnUew
IKw+eRcq9bWU3edJOjRVckDUahUa+c8iTwq8zv1cYFYhzbvNq3+6NOF8y3Lgmz2V
+Fp09razju+zYRKetbraS8Qmk/anLcjX2+leAbIYA1CdZZYUVEi9XNqh8s2UCp1k
+7zst4SkSbGCYN+DC2mR141tt5KSW4VJl/2qp1CFuTm3EYjn9o287LZRFJdbDlLu
I9UMnhdimKh/dInd93oqyAQ6MR+WErWvQiYoXmxVFdr65NtRTDKp2kg5XfemEGQr
72C9jli0LahABwolrVRVaHLQ5UJxYPeIm0tm2C6u/YlZEYSO/MJAQABc5ffbyvVk
7w6fKJIIagdFdUO8ItDp5+WNov/zz2iZwIAXMHaYFeTkGwSh8nTMhZ4XyN7L5OJV
GQUxuPWVguNlRLkSS+XYwU0jGdSbWO6AWIgf7JGGUamOOx2IGYhp3DORYcVkjfiY
gHNRITpkgBWlmwK+fSoXsy/P9jZYr5sXyEmoyUpNMK3ZdNb/+wC3oAZH3vivkFPT
3a0/4z1hqDSjrwX60EE6Gw+E54ZgHkeNecHXEs111YEM0DgZSn4eOjejMvEoGXE0
MhD5oW5/jLPJygyDL3474Ikx4x4523rGxfqMIhGZ19SwwAIN/6anDnCX+2BdsKZQ
OikVjVgvxzBiJHJb3oKpW98HnS48tBdW+RFhAiaRUMsoNkiiq77O5CYHn23JVpdE
/yOpnw+yP5QHhozIUmcAoazOlkeiUULrEpKyy1zPMBq5W9Q9cXnmtEcYGTFLh7Kp
Q+/oK+/P/Lp4rN2vPcfMbrNYi/6bpfleRXhSrovbZlErt4icVK1lgI5cmIKzADPk
UPoojdFxpeaNKC5CgSXyAojx68+cN6cDUxYu+O4+wV0pJWWE9OparToVwGL5OUkW
yPetdwDzlKXPJMGf5oKh30Qfd2YT6zCT+GT3rbL7SeMVMoaiMeWt68GxxeW0F2aZ
WpFDK+GWVX3EyQ0MN6dk6R/DGrIFo45F9xc2o70DHySrHBN1yPF6trDWIUVTMD7x
KDLz0hG1jdymqhEBgzAI2ZFQl92694GAeJDlCqQZ4czfhw179/s8KPlIo8j07YeH
I/2il5ZRuhS6FLWmvfsPKP6YHkGKGnIumQvx0TQJ10nsCu+pKOOkB9NhLb7bHWte
zYRK6N0rSoYd3LYb6BXaC89fvJ8BCvQ6qjR6DSB9dPEUZkCdjzIIbFQ0IZOgum8F
teKjuYqKm92ooaHl5KOXH7c+6m+YS7YwWFhiP7qTkXsO81J3OJN4hpF/pKUTUlDQ
zksvSABxDU71yKKvtZb3bSbWnBzSKvcN1La2PXWs0SNKlvSsBxx8cq5Tnj29Cv6k
/AV1U+CtJd0+hR6YfiBWM1FD15hCIq+uqgpIAemuW9nwLdCK+7ocwF8/bji/3PtP
mi6lL7lQe+bZGRmstdi6OfTfQIpVX0GJehICfyrIfaH4iFfCXWKbU4Br0O3WSPIR
s6tCHLGMH6tXT3hc8nrSbBZqbHOAwIz9RcDt0Ceid/Jj1g1Pk7MBSuRmEWYV3CNN
kovtWlw9KHTVBZFD/nw335pWggUPCdWz6qgdJcRehwPn7kML65OgJahCYPB3rdKi
8RsWfpGQ5A1q8kl/TgGkQIDOPpB52EsHQqLTsZImQTw5b+urqwkpNNPoS3jXfmdH
jpRkG54+5zvXBfC8VcjaGDUEVLYU7u750NmadhjCj8Q4NoVYnHoy2kmgZIQM6ydh
2oCH4lOpiXK9dj3jrsSn8NhjxtC9CDkiK8aWsLe8R29yuGNo1c/x+qCtd2f7aigx
ekfdNiBLbsz56ueljHZn5n+rU7G8Wf2Ph+3YxXcRbxohTb4iwCPtTv9h/VaZU+4V
sDR9CZNk6vtpW+zTEtkABu27N6Q+JN6/7VvaL2I1h6XhPHYx1y7dXzeDEyG39dWo
0NU0G7IlhCTZkH2suMzzd/G0jZzgzbaEWc39Vvp9QddaK0D2gDYsrt9JkAAr+dhS
M9Y70hU9+cG5oHI4XaeIK7epGdXCVkglEI4ANhdOZ9U0R50Pc2dZcVCyDxNiS47j
IVKm6JHBXtQV90E+YfLMZ9BHpOIyUHP+eg1K0BE1nuytdFa0O90KRKErLbbrCNOS
zm1xS66veQVauOd6vsSapZ472jQy5TW/FBbEbaR/ReYJ1ObXG/Zsa4UFkIUCpwnR
ju1UNwGpQwdx3AooSDgUCjRyCLFDkjDB51VYk5ndJn75OuXdYl7n9kRZNB7RriBt
AAsrWs0UvV3JEu8dLcxm636cLSykH0kjokvtgw4hARTH7bV81iyzXCRNAKD/Tqq/
LUAwUOeMzZPc6h+WK+a8RdGpdOAeQjc4ykL4s9A+Y8JdYtnvdUttRyLBD57KrW/M
vJaRL3Gre2MnjsvOFkkVH0wOyXyKokjqqTixSfqR3dFVo9WtNg3RPLym90tCbRHI
x04fmPteCH+JWB8QlW9s+Bg2F99K67U2Ymv6oqlmAXszZrlrKIrQTd9D0DMS1Z7w
GS+4yly3ALbPeP+NskcwKdCBywK6ozt0MkmKouTwa3a+2oG+zwV4S/QQbdLGZ5ks
P1SYmpfuhH9y11En5S0ps3NcMAsSWY22jZkZAjNOHKTGR9nEPddzVVBrbA/DhrGo
aNrw8GfU/4j/cJMdQK3D8F5zU0VSdSEs+xVDppCd+XKT1ZUS5NRctV/Jqyj1R4h/
Xa4B+RURpfc3jJbUTe8Xgelg0fOJ2pCPumnxkrEPgVsYCF1p7PR6+f5awu0BJrcm
iRK7AcYv+0KlMEZWdiZCvBTjyJNwmTVXDmUCPvOhTlP5NHF5cVVQoGykHZ/Pd1uO
mfYAhusK6BnOJ/2unMeseHzaOh78Pd0UUUToVbE+gIwEKa+0H8YmVs2Eaf8WjzHO
jzMOnCLG/0CViyOVZseWJmOKkqef2vWaBBFJbc7eEy6LXKgG+wkQNNSnfFxXjcv5
U284wCkwnJER4X7Evp5GIDuBPpdcUngvFjCcy/6BC3K1udRpa3+ZUX01VKXLCzu3
inmfsnwY7kxUFi8ZpLdVV1juVJ3Utd7GK0ZzJwC+oXgdYoMfLV8ZZkqIb7hVFUiN
AG1GAR1x0TYUXa3DCwvh56blmzHviIk47Q8tiEj5AjKh/OVwp7QxBk/YmPV2Su6K
9ed62QXs+cfd8HZzip3DM2BV5O5+iGSGuFF44eA89quP8+KWuSHSBTxduiZ9FYXM
2gIcpiiDJWJkhCmijWW6MRfxzpPXgGC5FYTk9xtK/QoKOdBkwiga4IeLTsazgiDq
8F8jT2k3gPzMFMrEZv7zCZ4QowlN5upGRltzGGl5qNgkLjNauf4Gljv+6ATCDizC
HG83PODPjIUvAX9UqJEDK1pvnK35KTy/cxmFmjMJFCqCs2cA1c7wi3WTCEKbm3tK
T0cXiqBezwLquVkgI0mg5ZSxU5XLH3aMwY1HpmstIGps6QYdlDQbRpB9ARey96/L
AofGkrS5Swrlq6iFTiN16TvQpyfvn5OCUphhH6+mXQEwhSYVMORoz6Ae49nua/gK
2KUnLhqjzuHiCd0M80Y6JM/te/vikalEIQn/MGOqwf7wp8uFkfJZ/Fd5GevBcx+S
nvfDavyIcjoNEQunqfS6NqobrvlWC3TjM8gWtANDTOCq25x4ciPDOjo34OYZ3+4J
s4yXycD+qpM4lp/TryVh83vsf4q3FetNy473T9/CrZAQX0VzFf3tGARsuzME+LgR
jhALOpNWOjZqvRM7pM5V9667OOc1hksdfgWbnl0Hmr1wHy3Ohx2VOIA+kwPDTmyN
bg/+guoVwmwrRdmW2rGzFlbdybBV25f1PI8IkJWCvtJ/XrEQOy0LlCmZXemm1Zcu
cPBJUa/y8wbw4HiLrbeNvznTmGD1mZkczguwa5S4al8+oXEVMkj3kR/ViG0Z396o
7WGmcYtdIcaJOxe5O2X6szR3AXWd1eVeTbQUCOhra6Of4ymYDpM8oxSW+UEKhiIi
qNHoSnZAIB3HV9zAjS2WLPA5Dwzvx365ka2vrFBnC923sybyQGfocXyHya1hcR8P
/Oaqqm3KZPCLWbICp6XzsP33v7wAjhXdHnjI+Y7WpvA+K+sbGMWzaAKtjyr2MOS+
he27W1ZdTmwwfYtbL6RcJj14EPybKWJb6205GXxbjWzXBizgziL8ltPgInl/+IY9
oVVmmsRv6uKymskgdys9azFKCzMGF/xia/eux0+wj9fTE0Y+cQ1nU7IH5GuKmyGj
qyyz9vT7w3qaLjJyRDrIyC7cPtTdHOBx3HgbKaTe7GyeZ1S/qIDNBQfhwa7mR9IP
xzbdVgWx29UpU8TrwQECH9/19sPHZnIcAzu0GmjHCFN4zjBFMdfZFjNqqbcJ1KZb
zJoGCIM6p+KL1jA/wy1AWqIDDQnfsyajyrkhsNIYaWdVLRlxlqz3I5Pl1GzP5Dxw
2csiWYmqjsC0f4QOKT6MlO6RBmNjR4UU+JVn36aw+3/og9q1+dm5jfkiAVXpKZsx
NU6vdjyI5DhM28XhHeo0DNTRRuRh3/JH/4NGxqzrQnqpRMEYo/qmXoDrZmcyuX/b
k+rJydvPABOBSwnRWO+Z3ByaCOsE0OCdsfmfdkwQ8wt/zlPHT4O+9KTepLT2KZz7
XhimvJWRsuuUbiUfDV91ySZgEPczxw4zIR3W/D9nah0XQosnA14f47+/s93NqtMV
pZJwSmBASIvAMdbpMq7LlIbB2LqGer7lnB5pLAkfAhxM4VzAEXqiu/TdjZf58FAu
kiIq35mY91WQGk5fF37HhmrLDwP3dxOa+Ln5dRXWYXV8EbDmBHjIkD6kqVu8yO4O
b75WTIiu8M8ocQshrKzAhaN2oQbt4HT9g4HMP7LkYocFC7qqL+IwKqoU8ipo686x
4xq0UcFM4LsX8/uCoaOxCy0dqml3/9XfE1beaBE4Vwv8ixxYhr5omZBDbvvaWyWU
KxLOP+xczefyyYafd2e9CBuxgR7ZHZJykByZ7IB6JUt7X8iEpDqDAVO/I9odMZMt
jWA1nteTcob1/Wi2NsoWQ0g1YOC1iaD4Vvvbb7wC9XEUvUDHw9Izn71NpajYqhqe
OJOD0SX6aJ9JhwAVqNM/4TB3qDSduuFMWi9x/bq03f5cw9QmLfS2SwQKe7bcZe+v
VDEvmrxknYvnnpI4oWzRWEbcVbRCNEt8ZYtznI+pYjTQQOc5k0QcGNc17fbimZ6C
TBDUOhekv0hNiQY4oWsHOcbgUClLjzbJd3oZTTw1kAA1SF7caD/qskMIXkblAnec
uCSosdOcWO/ix/9SdRqXsHOsF2kQRL/yrYUiOI/KtbAQ2ef0xG/o2pXzxBcc33iD
QjEfxyqmIEJ8CRXqV5gIhOXFlU9tF4ZX2ir4qGGMQSz1UHTjat7DWuCXJrA21sLy
aO3PGx8kC1u9DjyHSiypqeAGUu2aBqM4nrmtXJ1igumVSRqUCx+MmXLFoyjGN3uk
s3nA82bl5Vff43yV3kMLHacjPLFhEraL3MWlVnxpQa7LjNG+PMvXkiQoDiINHiMY
w6yd0pKKfcudbd/VtTWOCv5Z5fKl4b6xZT9Z7lCRtJW/zIHE3FZfBsmTMr0RVLV9
kruEzwPsE00+L8iqqYdbfMbkZ1xDL50JINbOfGCF4afewUMnYj+5jiHOtvw85mzH
EjmS6E0QQ8hya7KYT6vdpvBkzuMDkxpJoBkqFKSfm7mo5arK1n09eTfHojlo3V5n
qqyCBfhAuDTvV6RWw5PUnR7A7ynPWCOjVai/LWiiS+mQa4fHT2wm8BHuEqrOdty8
v13SZCK3ANJhDc8lJy4wTzzRJxUehlqGjxCcuuJen12XuljU97OOPCFGPx8Ke+Z3
7Rb6md5CEtYj1cnQDtWSD3PjbrdSKdFxrqNiGkB3aNgAMOdcMJYn0AoqcpyIy2jx
SPJY4di6oYTL4VZYe6uVprJVtk5snIJjdmGkDzFq38K2xWTZ43dH9mDgmanUWOuM
njHIsdVRthsv+ZnOIX92OyD6hoGw9L/1wMi0y+hacSOW/UY6pL63OpOQVUNmrH6E
VwRTZxYRRzEjYrfJeWInW6HwNu59LP6Z+kLnGaarniSkOYWcWm2TE3acPijPGsP2
wEcEZSOZcg0P/j+rLBJwprczAUboY+bvOZVpyLQFjBl6jeyHvVP4rLWo6n8iOiim
iZ2m+CAOTKNFwE0DsNp2uS8MVKL+HIL6jQDmSeQyTY9W8MCaIo3xxmRa4H/tj6tq
ZKYue+acT37EbwtdMFJYEduKth4yEG7zs/QnwNgLb27sP/0/HzTbFu1uwpXzh6gK
a4I5ZWYlj+enmExQxS5owdpIGEXjL/XlM7l2lJcL251pUeXran0ZNoG58Ev+64Xi
p+fMg9ngjfokmaZ4mg7TcW+E4+5NDn83IrnWP6TzkVey4W10idJXaZRS4ieoiieP
9GyNKElXd31LkN/VM+77HqZp+BOHYD9JKSDXSfKkMHdDp8h7wRDnJjn0X6Bv2QgJ
cerbmtI73Bmy34btttE0Rafho0K0kU2lAFe4/TJ7QnH3NmM5Ga5SGc8j4pBunqHT
pji/1sTJyzWmdOpQTRG16QMYGhqZ5cR4gNS0uO4eXgBA7YfaoauvmJK+BZTae7b0
xtGXevs7y0mGgfYyYTPr+x3wVIm2gBdekpSGqd/DlIOTI+a2fSeYLdDcVeF1cLA7
pt/i7PTsro3Qb3ELwj6VLAJ19dfAeRZW+54wHUlF2IbSe/ieSCEEOM+sYoV8i81N
qq9yRnD+zv9t2eVpf4TR74MhkQsPf4uQ2hkV7sHDZWfnuakpCTqPOUX89Pkg254R
6QZSJNyn9f1lDBLPa0ShgWBzCQZi+CxQCxkLS98OrYt5/v08IjwYdOLlItRYwBGP
egGU4jUFsrVCdP2cIVcpSLQWj2T7RtyIxl4CXZZIu/CKQL1SWHiQ7nP/WSb8qELF
32hq6iusr9KWDNjAmbV/8psJzbWjFd0j0HGXJuPN9nj+MjYlxf4gD2XN16a91+Aa
ciCmfyGnLsHwmxe+H7AfBtlXxKrTXSwQ9+d8OeC9FujTyL+LjWJvYt/hT+TA0bV+
qji8MTE3gbjmkoZIhxrXhcDehEsiFGhqwmE3lktMnxjWmbPCknDA9mAMjFuvFzi3
ebXdSD8su5/xlALTaysY7vHmlRfaWQQ5DALlEpMsbNABukq2+MQAC7bPyTopoN7v
Zm74jDY5+l+B0IwSLffBeZnEhUGQf+PA1wJrZ+FTFGnnUUYYbNeGPHmt2yPRnuhF
ylgtH3h8OYYEQsF/V7dPj+Q7hFcTFyouKA4giUtvakM++vIGQFN1+gP8y548wOwB
+3ghHRlfc2rOxWgj5eRpEx6KwwHylESh6Iu6rzhB+VowH6Y/3JsaGvQm6QrS/oOR
ifbMYqmE3qoQl+7C+689JV85dQnWW5H2AWfDQbfq3r+Ods2su7dWWJeKdEZzD8io
+4dNS9ri2BUaXyp0WndWu3BLrkIDhtrCTQeEzKdIaykzc2cQvjCmh1SBUKJImzJr
HUyMKIQ9c4fE69+tiKLgiKiOHA0Cr+kRXFlErKMEb1fHLB2WxJYhLLfzkB7lLj3y
L1eeUBaubxS1oaHofofpBR1nNEIrx+FyXheVj/bmBzNhVWV0UU9wm1NaKSYv7CFq
kLVSoW/DQ4U3rlMC19BTUUZjraG2WZD+BOjrNGc073hwQ5Sry9MuOHI3/zeGJTtI
CTjNOKQCECFLSVg3+a1SgmJvkRYYk2bkhWGbWIS2ZfrzxYltnIrXgyw2XemBw7LJ
UIW0QmVzPN6xLHmBJiRuTVM/ISJH1pp0kvU9MFAfRtlhu0zp3YaMAR9Jn9MXhpBu
isM4D+3dCcRPt/EnX0Yu5VsNxoTFo9mnjersPOY2Ec9cdHF2FlPrfw8hMPkYAHBG
6HCUh2fQPUhE8llh3BRLQQ31mkdasN7Ia2ErXfD3dQhjXCN5zUjd9fwG5ToseAaT
Rq/pjZVgIaXw/jyuSZJ6sy6KnwYRXiWnjkr6O8u+gfABSPq24zEHVZqThspWyl7B
HTYqnd8CB/7I1dQevFW587jEUvgYdWIsjU/4fqL/fGsHXsfRryFCgEHlcrqjxiSH
0xCXNwIJo79tO4v9/ZxS3xwz6yy/btJkenUOZQ4TKjZwrBQ4qyPqPN8kXxNuWLFV
bBfkjx1D4ZeynbB/Lsnd6+n9Pec7yoV6MtTc1MSrscAs/cMs4sXnHYH6Q5wU/e2f
jm/n0rnxeO7NNgzqfa+fRuj7G4B9UX4MOw8jm1s7ymbXEQOj9s0UocsFqeXU+DlR
CHkBYFoUsbQQ+qhFu3Z/KtPlzsn2THORpaeqxAp2H83Rw7Ip/O2W4fhLNr7vXgwj
r9dbBU7+NHt6j/5tQ+9Ud+jmKrwd22cvuPoFKVO3YiX5sJlZl3tNBnXfRfhPMXri
icSGpVfORbrYvaN8RakwIaDGFlnOuXooVC+jaFPiUMVoRYV2ZvodVoRxrav1ceZs
aVWk6IbNHXfbOScNlsoJL+4dTRdDvhAGjn4nK4kL1PMu/30GizLVgYmHGIE12G0L
HGbJ6A/n5g1JxsGyPePtu982uQBMEM1BE9/6mf7ZOgTkdImg8Nt2ySjHlJ7WHSa7
fNPoUz3OHD3kjuKvs3sofjBlw6+u1SDUK/KOg/3a2flcSPN+vIKCMFjcHniMwvfO
OEaPDghAkYPYarkQLMWAfbgVotndVFGfd8+ccAIUWYkq8gFer6H0nG9zVU8EWbLV
00KYaSQYABk0Z6VJMNTzpe5pskeDqE5ltBKZS0Guuwucx/Z0RCTfg6e49cc4GE7l
9sBXld7Xae/voGJsgKNhl1iJHdY64JuB1f38OKp97VzlVb/91i5V0Ldrd+meKf9R
hzfBRVM1j5oMJXLc9ruLVzfH8LPNyXo+PFEJ3rEUcYL3bsthxB8aAyCpOz7oTjs5
Fl2mzVuatHS6H24voTJnistPRCnOTRSUQ7n8ehsdjb+By46cGRp9YZ0wdkKACgCh
QX4SMN3skbkinjK0T586Kkkt+iy05YMSH9HAGdW4txqdDuC3MehX+VS7CbiJXZeo
UKez5pMY9N0ml+59VgEtWF2dRHj46UqgubGER7D8e1FIJX5d5Oo++Pv0at8ZvygT
eZBy4SgtyQFQbQirL4vU8DFiRS6NcMw/O9irPAiqQkhBOJbBMy125gRGo8oTwghJ
sFoc8xL4kqaMPFjVXeY2FGeWcj0VMZt3vMab/jrixVhJcPqEkNnBBHuR1oNChSAP
pIY6APYqmIBOtX1atLif8wuYcFijE6akkVFYTeU5l01MHScqBsWLYCDj3OzgebIo
UGq1eDViWghMzgC3LNDLFnNrysMfnlM4yXiBhdWWp/IrGEiPiL8Q1xRUs7YwZWH5
gCfV9Bh85+2HZ7w6fWlFGDWiOfQpMfhPadzbSZBZMGExF0C8waRiQ6ca9V04Q6TT
iS0cs6GJZ82UZCDouADG7j/h2R1r8Kaa8Gv03VX6SKR7X+903fTFV6a0UVGjNsO+
rDGlflAVJnbqu+LR+c3YebwKyVG0rrXN/yuwhvUH0G4CQPlAV4hqfO7wp+uTKaHy
QfIyTK2i0Z+3jPi61nHQ7tr3C0E1y4Pn6YRcLF2eKMGv9NgUI7ZIpRSPcNBjUggz
vCuzMrYW8fO+9qsb1hST0Nbx7CT9c3k9eCYkjFcphqsSs/Bo6BUQKpITnS0dF0DX
UnzyCDJ55z1Ib2IjTzoqUZG9fUrOfi2QolNBrEzJZj92xqCSWXsma6jQuzajq3kA
0Jw/DKlSAnygXWQarfuPS3Tw5mkBHD6iMo1RlrXq7xI2yjD1BWUcx6gHKKiTQ+db
2m4peYoancrDCJNroLt8zDzo+Bv6LQYc6qg3seehETI6DKB1JCpEaSf8VSK5ZSdn
cURjCg7gwbAs67JtXMhqqPGFzXj3L4wgkxjka/gpwfdq8jQ4+S9xxnz4ZqNHQSVb
YjY1OgxLrmth1ABtYcayA4+2jW2/gMN8zTIbTx3wRRYTImar5ea09lYW5XDAtyVt
mWVfBcVI5S1u6QqEG6/ReiiN0E5P7xCxd8gxzoa8aTzK3wG1Fjy6ygUfv6zX4O0a
nFi5mAvJEI4I/cjW1fwhqBAkgYpJ/MqdyriHTwEC34BYxUxqkuKLGnzUm4CGt33L
+QyjS/mCXYjqc/2e7cKbrnX/Gpl6pz9q1L43ijA8UUSvfRvbYVWOFqiYXkcKH/Qd
rB3/9cNw7WY38/P3pVWazRM5bpUXM1vpEmHFDuw1w5esgvIQpljnxcNT5UiC1IPU
n/mYju4Ex4A6yJXJFCnmZRQHoBAUuAkiKXRaWceO+m5N19zYRx7Ls1v/+ppRfBvx
C9z3o0+Wji4xU5nFh0QO/sTJBGMEcHa4lse6Az8+AXyT25n/rqNmPS1UQhjfneyV
6IC3l0ysNex3eg1jpJgHs5okSwwDjTvz8IWaDbvU+sUkQr83F3GIIY10CZy9TLnB
PSzuoOiwCacwcqhTj7vkvHf602fdlYSCvgAhrvAkkuUbV+rjMhUJ2MXqoN4vl6o4
OldgVkpCBZLIRZDFNKJuPrL65Nv4h3yxUYLZwpJk2yUMdLwVTFMuzDIqOYex1Dsv
qaCQBpqC2jBnw96nUte7VwW6MNb68ulJQ9IVxoOSfO8OiRh9pAeK9HqEa7p9iN6f
YNMM2/qnvkHcw0rk7H/skEHHaBYcEKFqOCepjsds++sY1qi8L001R9b9Bj0yHEk1
q6Vvkerg4FcGXcHrDHYylwvlr6Hs55PM7csaDQEAkiLfn+tTvCTUoAIGqjMvac6K
F43zZkfRFVAzNteFSSUy3CpRk+ViAh83B7S/K9P5WMF0qx5m8fZgJ8IlzIAsiNlj
ccA6twpdCNz6FYnqyrUw/H47PyMVFQGl3EB05sRQOgeAeXqGpALC2PAou9QVYUgF
PA1BpetX7thmdobSgMxH8leM72oe2JaSSv2UGj5ybPITnu+wUWLCW0NQlGclgGWw
D/rJyCGBje4LrmIcu51Mr1YhON6AcvW1FIEhdJ/86M3DHPeRGYd3R1m+a2S60fPq
n+LdhGY/Ym+naLgkxiFhucaZg2PVPKqQ3GWgd0P72fY8XXXiqk3w236o7cYN5GLA
DI0qEOu/arDWQJQ4iUhWNItHDZhDv9mcui55izYzKh9HYp9QUwQugbPBTTKdYGcP
ciP0oQydDXI028PVubpe7yBnsc8IEpMK4U/0AVSAWLRRMCXhknrsOSuq8jrdMTE5
EJ3DHVj5perjuM4oaCluhV+7Z4sDpbLIsWTY2xmM05nRnJ6goRmFvDpCfQ44t2XZ
LUKPma3FfwVBEu7dRfyDNoC812dpki9Zk9+QWD+dezpYimSA4xOmsLVqs4LtU8cJ
3rQZBDJoCHtzmnAGs1/rMao89hKDxkjYaVfR4/1DzZ72FYOV04lKyhn57o+vdHnv
3NXBftIYSgFR0+1E9Z2NLcSiMihfP7OBn6Z3kyxSnBjyQqMnqxVTZQnv9WKcORTT
LNFFE4on2QEK7IWzWUKQJjbCKrq+KWbDK0fKz5Xh/JqmzPvZ73vxYbTyib5ElDcr
9fUzFl03ZvGp7jsOQ0UmH5OqlAxad4un/mC048Dfgg8Y6TDAzM4lf3utMhnJjYpU
lakq2RlMrCThG0E7Xx8uwi2MoA4/ooIZxu0Z5dv/BvwuDxlmGx5NvICWk2i1T7qn
YpWlrqF40OgzZmKJun1PKM1MvGgHcVYAv8oStEwZyQQYF7gdvLjdbGE3fTpLvpDK
9kuMZ2Y5OcI76+qI70mP77H/bMrr328P0md1KYNR7MijE87eafzCnhxCMCW+Y7v1
phsOSs5wC0KYs4vdOs232NDd3+Y4UlBZiwZpb9ZUg3xRghDprIw2i7qtXr0yj/r0
QjP6qpUTpytAn4DThP0HmSWhrwfIaMY11uSyq3VxJ8SdASG96EzObO75j2jmWTRy
BkPeb1gy19g46CSQTk/9a3Yn3AjIyCYSLeo+3wnIlsVn6DhSKbwozMm6Dk60bRP1
nmsu1lUGr4JmfkPJqPUP0qjHJfl/RnHU/p2ifCNE2KxgibUOaik9JzNloNQRl4pI
ToenVejuK2VDNqrrrPxlE3rSjYaTyO3SZXvdSLxPoVL7ieUVp5tibuoHB9dl1bgv
aY9NrmOIr7jm0QqWdytQXhzTQXNzg5XjqIc/ulnqu5yvWpMF2RaVolFJcg4Vjit/
PF1iBXvBj1tApGAisMLDgYjja1fkgN3c/oHUlHQxqxbCNyFjOX8/LFT3N5ktZ2Cb
AosCaIFIH1loYXXEC2aDU3RutWaW9QUY7/jdw1+X8UsekhSVt/Mo9nirFKi9K3Qm
8mncd173NAt1FwegCtJAbV2B2MS2whRKvkQJQFl8yqnv9vVEpBe9btAJx4aQ4yge
HPEkMNFj1sehf6mvI9ChWvsblbtLrLQ8C1qRRpwJ1lRgw39+NWp3PTbpyl2BEdKE
DWhKnY86k6VLr+2GurZh9HyUoD68KJauYECoUKDLcnCJqrs/RXIcaqD5riwUM12r
6y55QoEjP//7PLbQ/ZQ+SsOinbdQoPS3+ABhTA7PUQZUPWaZU2vKhm9oHc8Ua61p
6YJQwzmApwTCRo5FVsoLm7F4PtEpqi0y8nN92VZWS9zZN0FPZ8/lmr5GLiIs9lA1
cYPuqdDFRmXR4hyDcsLjvQjlpvtwMpIbVi2iXP97AejbobzTGRryals/eFzE/r9k
Jjy2eyJMkOmuZ7m3RMbs5TiL4iuuQqbeHFcpLpDWmCQ/KAWOY1+RBNA5Cdne5WLF
VtShGjttJjFGXLnUofY5LtojLXCsU8FAqe6tgeKDzgKKM4oYlNFwdii4+1K53I85
uxf8DpC05lMZuXUkc/S7oEQtxQJDfEqi3kqFvHVzbfQrXM/FtJZKFi/h1YqTIr4n
nSTHs2CrzqG80xBJ2dcDXgTcUu0hSf2hlRP/miiZ4lRv+b2yXvE6Fc20/4IgWbKS
SMSc3NwTaJinaCeFv7GoXqcVQu6qa4/KZcAWlUmNv66P2QA33xQ12W1xxvpRqRX5
zgFW1LPeCwCuAldkl/UWwujOpM4PI6Lrx3zZAM4jAEaqtxTmVTmtvqmNexOFvYma
NWjCp4dmsqcwdFCDRMPl58ijUHdW2J7PiQRMqWIrlSLC8fXb/BSx+VdnTTkRM1pP
AwM6U1RYU/44Tq82NDfFIBnPxRoFcYk4qI+b3nmu2/MzaccUr36lLN2pZNm3J47y
yODu0gsNrcjtc0n21Z9UD4ufo5TwFdM/vTEIvj+rLfQogDUBiVACin6q3xe5kOks
RyXvLcKcs+GfHZBua/Aa7OlSu3Jhll3vIl1j6S1UPMsrpLuOZJMmQEQqK67gqiPl
dAD3/7K3Saj3AV8ONJHQMPC5/HwqMHfLCjXEsl7a9BepY6ZXo3EFBkP+wMjVurfj
DoxGQkagYqEDveqlw7clZmfM3EFRwsAd+oV/GNiyjwObPf0ac/Elx4P+C/skijDc
UrRLifqUOzIsOUDwfYcbuNGzHuLaHdgX/7BykBZUV7538lOiYIjxpkaU/ijuOXWw
dLEczOG9Yppy/0GttjHUZlvqPoVwwbeOnJGm/oqP8MQ7mga4JnCj6kaW5EfVuXrY
c8ou14tm1mHq5so9Uryum/XMvJMh2tRCEUvOvTKR2Pekw0Zf+UKl3HluQ92QzBtZ
3JIrYUVGzVmMHngE2ym2q4/lHEvrKs4ZRFmJMdXUVO6zcF6034pD/xIsAtLrofDb
ifzsf+0QzGJbTWLztPXAV2wribcdrKpchM1dYmkjOJ+QBq6HcFYLTzXintzl6vJM
IcVBtR9Axdemq5dsbWQlYUDoYSnbyXQRmS2fl00qc+EjO2vo42P98Vx3He7lbUOW
sdwgFG4jJMCRKtY/ShYH0l5fOzyr0VJRqJ+fE+4F+F0/lVbp+lz+z3sL4Ypqh7Nw
IKzSozDnPObK4tX+IOiIS2Ts/CiENdijFnijFYK2NcdeXhKIpH88ytn/kZYYvwQy
WpZ4jAC+kbysTrMqUmJrwcHlUSoK2JmHbkUupKR3WJ1EZdPv00DrVGAcE7BFAx/u
S+6EC3izFQMRg4TPbeDXvU0rZ/5cd0L5NnmzshII4FrpA5TWgBb2q8+LvqViuN2p
k1qUwiUwBlpO80qhhH7wbd52dmlujtK+X1qwu+OmXS827xO3z0T40LzTjNxMxJs7
kaBoy77mQenojTGc0ETDteb3iVmtzVomN3hSv0vQSdPmIv6RmhCIJxLQKrVkPr2w
99Jz8GTDnCgP89AoH0iNdO9UTfw+waLsZogr8A4C22l8AJ0PGVsHBKz454giOpYg
+N3+ZYhY00duDIHjHOMo71UpyezncT5M3FkN7jnNoBJIRB72jqscZeTqG8XAzwTo
gwi0Y4awNuhYgGFW79diLWQRuuRxtCnZYB6KhJ3nj4b5du3KEK46jGsvPfI/5u/z
h5gJOJMV5P+Jzh31y5gcpevk/3ckTis3kx6R1eVpepTcAU1OCEkg3uS4Pn9TKbb8
4ckv8AVs9iJovGTseInVhb9GjOHvMYntrQE8TaN6NTUFTzHxXuKkEj3NEZ8Nt3hP
i1NSgcshx9RWI5LSqpyamuYLoTABZF8UJzWo/5ub1nzL0jxrH6lcJZC+p2JLosqd
Z0spNfKs9OYT+V9quEJP3U2YqgMSLWgFVB+F6lzQA9ipl+gYgqZ5E4QPYCtXvTiG
OVP4STylkN5pjVIfn7AS8urazAz6rGICEcRAnLz2/n3xQfTqt54ZGHuOpDTcLFzM
17VuwdAJmXccoFNJXJIdhgnxtPivTxh3M4vTIDV/+wWXnFhLl35Wkm+I2tms68Tu
+0ttEg+++0oA2okAr1HGhRF+8RjXdSd/Q8sgC9AISelfQ9E0OsySIU1FWYijm1S+
gQ8xAPb8n2E+/Y0uAKmTtkBwDr+xEDpeC/H1mvgcwmLDjTp5a0yxJ9Fon+kYZWXj
0Xcl6RLZ9DbMqYjmrCl0tf3ia38lrxsfzEd195KfHloTPlyD7jr3k7qR+z/cBiNC
89vlxJ1PmeI1SW3wsGbPdxZydq4DmRWBZhlnintya5lf1tmxXpEXpUMQr1iwMKSx
W8uajww+2mUqx4BGVEwKgaHT0Q+XrJTtNgNBzy9FGLXYL/7pPc3mCLK3AnWf9AWM
Nf8y7kcTD4Q/VeU2R2XyI8IpmJkfnES3Sp4DSrio1qtjYbbhJB+9flSvX6YlEotQ
z4gVbhuR1pN3meUUYpuKccIF2Q0oSnr06MAHazH9y6k1IULsYEE6z/3zFVS6KeNZ
4LrDTvd61TattRWmV5sTzUC0xy24Szj1t3qzuR7/KRK42FnE6zRnrc/O4zW+MMCk
rv9VNg+pJTRYAJMeFac58WaTYUq0xyb8Mt2RghJMg8fH6UMaRnOuXSz0fhNNGbWx
xWIUARroqU0kngtK880uhdJw42yUlsnIV5P3DfuR/L3Xbx14Gk7651U/N5DNrGUn
6Pow67bnySZqL9/tNHIqg3dR/NgvM8nRQTxX50a1urWw5Q5gY4CX/hyFfou07Ixi
IsEyaaIx+vjrmaWqCdwCaJNM+hDvFdbUMJzr+XlxrJTvxKzTkztiy5KmN63SPAdb
QjqrcY8kgDDpeRKsPZ2NrU5ephcmNfyDgoQ92fY6txjrpZXp5bO/sJ5IZM/Cnq/Z
/ZaSIg/QrWuw7CbnRRu4I+GIAimFDyKaZ1QLO6FSIOIbo3ZNDUswccD8VdtnLJDU
QNVt2ggDDICTa0PAlGGy+ZkkSMS9Jc+dZs4ntMC67iqACfeWzipXDU/QddDh7Y2l
oljg0kHWaGH5SSHKkjpAHgE7dPt+nRvUfCb/OxLsNtcbChv6WUYUid41VMfRwFb7
J8Es5Psbzyo3EPyyULGru32iSgqPq58RSfW0+blK6ZNbscnqnw+x8OH4SFLqevcg
kMusXzsDJXm+zUHVJ5e4xsBJz5OJvDm3qmeUEPHvro5B3J/SKjVzIhVQTWfoYayY
TIg4Kp0WNjYd5nXRIDLPx+u3Tu10fWkf4Cbi/albFDlVLEO56/dBQrxlg4DDHDOa
OsRs4EblXKfOIMs/oOe852JW88jwINRhwoDbmHH6cmvhyb3TnyFs0j5jH+ogGsXY
1xxiHdPbNIr1JEiSNNI8Z9ZrlLbmKZHW+3k91Yl/39Fp+s3LQqJOuMWURHqcveCR
CsOuPgVK3AT7q3mQUf8U3wVxlUroVc6TTWDPhRleh8OPf5GrwJ5GS9IYDukkSpWH
mophXxf2rLpcYN+tVxyNCYZHZUmC+xaYYvChhetxmrI1ZyFIs6daSvbTaiqm+SvN
+feA9CWkP2443XvDWiQpPaM2fAU0TGEhEQFdS3OYFqszyD3JxsWnOXZevQAUF3NN
SyHtoVGGMYFfQETbsQZ/sK3fj3EHh9Ykr2uWrb+Oh83OwpwoD3H7wx6yU4hxvfw+
zhRdr+9XioY2klh7UpSje5jVyZOA0gzQGYnbJBQj/cilYnG2iShStoQI5/SnJ8Ig
0s1J59FloFkZgrA+ceoToAu6/HH4ZZpJyUU1/6ihP3CxK/FeevS/pbdmaUZmpV/e
kvZ4QawCo66OzkTu2G7xIzzSrBwocqbsct/Uwzt2rPUPSKgQdiSCeIdE084cIUeg
wNhAiYiP9I4w0f6tK3d8zY3ffmvkUDxkdlX3jYX8Ti8s0c1fkY4sOheqZYbej2qz
YEvrJ9MIkchaPpOGwgHMgl3mDJDD9/G/FigPRT+45lQNB3TeL4PkmcF9QBvD4QzY
lasrL9Plv2+hDo6T19wx4N+bdESxYd272XfyftgnGnIifkfXPvH1rWr/BGXcr40a
5Hqqm3n64N8EDu5T1DaBuHIN1Of8yhTArbpiG0130M77hY+JE6N57UikwWiagWrW
zvavHixX7oMiN4CuyKoaBThj4Ky/KF/ZeDH26DJt7onmg7OB9OYpiZMmHDlf1JSh
yUfkDeEv8AwgB1QGAO0V2KXfDXbLXwizF8guLOhwYJdwK6BoHKBJO04GNncC0Uz5
iwGC//xP/3thraYcox1j4lO7e/JgjzJV+12ik878GEZTU42ccC7XSWI68nobRWiN
gEtdp7nE76yRqmzGxbwoZ3gKVF7WodO8W+RSsGztKQVezzlSyMrA2beDj4szrf0N
Dy5QZu8Bo6PUFTXiavm9ktpgeFCjObgZZGCNLj8ZJbpIdBW4MaPYi4bqRHH/D85H
3bc4v9phN5Jx7LpSFzbf2AIYc+LR24KOfHgC0mcPqdSEBrE760wPjQC7wnx1W6jl
FShM6sVzKq/h6PQQLILctz1ENIWESEW+r9UqQfr4BxBP4RHMPub4qAMX+5nXkMoG
kvUXh0zqwWErf0m8IoO5JkN6lzTR1q28oG1ojbepsX0GK7JhLKSIvZKkTsV1VK7R
0hnjN9FJeddf1UmXVuFzP6e7VUH2fJeM/NL4Dmzt1Ls8+QQeCdgLzJkVvUy5SQT9
07foOlaa8P9psVN8f+Yvy/LEJqwwIKS6kU1WZjpz7BxcGC8kKc9oBT7wW9V0VvKr
pRpOqf5vN94brxh2OODxO+UKBPQ1Tuz7NayGYXUeLYxVfDuGvnlMLbIVBgfwsQaP
RhOH29xDp62gs1G9y57YBvtlINPk+Yw/RCv8m6EV1YAchx4hDK0/ePe1D4IHAIJe
fBJK1v3HGk7d9dFGVm10INFrJi26wdn+40kEl6G+csLNKBRZozidO6rn1XnpHs4Q
qIBpdN+Ijip4dVY3sCwn33BgxIXCDGvfNXgC6h3inECPFuVU9Flxoo34FNsy9k/A
SZeqACkGvGqhQsOeyAgyz7q0AeIRX0vpvGVnDOHvtDPF2rNf6pvvZuy1qf0zbsoh
ZuDG9AKwJr2rCqXyLDvR1Z8EzzHPy/4wTbQAdWlGODWde/Mfr6ioeWcx9cb7B3U/
riNXbYRuS6orEeVcX7D5v8DSJfdG39C7Srywaw8mHtd/XbSAetY7ZJukr8rjn1OM
a4NMp0UqTGchKt1uT9qvpbaLjDHg0LcpFxZumwVoUywzLakVLabv5JVNgz7bkk+R
h2ai+qJJn0NzjfmI+or3djh/gZ6J6t4F7rEm7y+238IlNnzImrIz99R53ogL//Wt
r7dBbVwOX/Jh17H3ai1QPcCaLG+jwdjNY4zgoGHgIdEhJPqehmI3VcrL1rc9p7g/
rZtj0o6/dvv1UCIVDVR1wNY1SV3UYwLGA8xa1ORTg81f4K+AX5RXQq3Xwu+m5PbK
COLOwvZp2MnhN4EjKNRTPlifyCzJcl5C0lBD6Ege5lQFPQZ1KSdK/2wF6bRwE1Js
G844FKKNJ9iNlhrrui+d782jChtQX1ziZxqcy3nJqBhCXVtkgXbbyHX1oQNmz3sM
IIX/gvcfperKwld2rEZfzuh9hLJJTNdmKmWPAcKu9d+vQcGAfKnpO8P49jSQSPBZ
EO1o9Z2mvycnZFleJCuQyavA0AGN25bmA8DVwr/ERIRKn4ABzGITPnagRkJaZgn0
dIq8OUcq8RhLMB6xG4DU4tZCygD6Ld+mXvXHHAgJR5KuS/zgF4HWq0zLivBIfnE4
t966lLQuKQuh3/rpIh9RNHoGcAO6YsxxJbVMHfYXfEfzH+wP2sBPnljzFEDryWGD
Z9ZBe4nFwyxylmK7UVB4r0Q8WpPr8YREk+0jDb1fTULzj05qItzgw+YBKoYoTfQp
ZD+TWmREOP0C/FXpeJT3VNkUbouYn1n+Z7o396udRlmfEdGrIWWAQndpvrfdP0LY
VsUjpPWlU8MJVr3FdLz7os7anI38RFW9UgGbgw826HJOBxKX8yq2wP2fTYatNKRj
tPHsJee4D1u+rbE/H0tts/rRVzobpPKX5pUOxlA3E30OHzPG7H/8GS0ewESYnkAc
0Xn6vAbodktuVFevs948ObSkiAcx+vAFbHRsOLtw9SH3A1dwG8GX9onz1opmydEB
qCDxIwf+rUGXQRpcnrkd2iCkkl4IsSbs0gD/loT+VQU4Yb8MmHsMyEddvXSKAg2p
gokE8sH/MjC8nI0nFZ7lDfdzYRe9ZZCMSZQK677Tll2xEKQIDfpKzchSfTtS5ivQ
vZuGEheOl5T8dYtEMzW4K3Z6418RwAhPkJqM9iJQjmJCCmczHOPRwvXYb8TwOXbh
NPgMsE+e9pD02cDQLrRcsHTbkSes6+FWaEZJWFtyu2r+2Wj1PgKMlrBAOK6C6p+X
41QXpVRMnGxEaVmlwGfsJB+fB9Voj9s0pnlG1yqCYCtKa90blZA5tAPXZGut9hNg
kcUQL2RbgnGoIufZA+39L6LgCd9TyyVrHyYzdcEDjPam5E+Jou5JD3Xul+O5JqWL
23wk9lGsJfZdxP2dBln7PgANBqM8qpOX9ouy0rpn8J5xN7/sYxJAdHCwFZtTiu//
ao7KL9T34ucDdNnuINlzRbbgzQ8DbOmgcD+guABe2e3g3e8xKGu/A/Gr30ngiHwg
f42GGorvXqtBKoHJ8dbTI7gtPuS39Hzzs6HEQ37WVZiTO3e4uhWayg/TVfaIIbOn
Dnf0qPnrY+btPyd3rQUgf3mSB+kbq4OUWz47QPCqVmFehQ5FYuQVm6vTMUtbZFUM
AYxqWeqPWjSANeIUK0xZ3nQqw9n5KU+qTsOb6ckmEitk3UyAQqlKgSMggTWWsU9g
eAxxzdwHmFKVlsFF6VvUdPWJm8aJOXTfOsK3kObidJYhiRwQIqpH5YOh0ZaaViwC
Wpa0L1Q2uJIuP+0o5Mm1Vn0BFRuiyl9tuI0oyIoWM4RZ9egcJuADztixMuE+aM6F
f7fIB3+doruF4dnx4v6I40BtWBNg15w4aZQDRhV1eMTgI17hRZdqr/czeemqQdkw
lboPXzxHuXt0pl4tWj2u/kvpgXpuz7+SdaUXIz8HQei/GxunWaXplnDiNrGud1IQ
AY8lzFsh8tSUEgxILZ0lY5f3aGUP0fupKu9rKTAj3AJUuaEqCxOU492bUcURZ4ve
EJ+Kic27N1ArYD1xsoj88sX6QIDV/3gRVHPjQDukfbi1u0U3kxNzRvv62mJoy8Gc
6qYJnWlxpXX6VUg1RYB7MrVRsLLDLu94nMQxNcWbky7Miy6+Ejlo7GhKhdSGWXX+
WYP4RMG/VPZl98rnVniwerE4RCRvXW/JuWjkeXC0S4m5x5bveRPy+nvs9CV6OhjC
9bHOBrgXDl49as5nNwa6Psps9wHxPQx2OyNx4+KNJ+jlJ3gPDVeDvRjFlfiPuKrw
OuQB0XD/DshI007o3f6oO75TEC8RyaG3XeVwfcNso3/0yp9AyCDFoaGXlmXfja/d
QGUyRFpB0ezcp8jmsUbU3IRpAyCvcLdnv93v0pkvjqC8YoEIHmu0EAzo3m+NZJGG
c+rhz/x7cx4Y0ObrkUVR12UCuXNXcO9xAdftZWjTp3JyAvii7LQfDLkbleAJRj9q
znfoyubKZlYtU6PeBzI9WuWKYnFepOKx4ZPg30siXq4ohBupRHNbqC9JW1xuYQUx
QJZHP212OBktjn4TvaOz2WHEODT5j6D22x211GxhUX3y2xMTjs057L9vcgU8QgxO
A6IInbh955b07YHupoekvGUMWA4HZEQlO1yr+vl3Xy41YC8Vk5D4XQGJ5klqOCyM
uN2ZM+CnZpQaX8Bw1LKgEKX5N1+e3Z6KN77jYuHUs1uRWJA9D9H7RNq61TBCKzna
zR4Gxn2ForIEulsc4pcbydVRmFxRZkHT/0ZKzWvbkJ+UcjEKFB1jbAUFjBQc89gx
tva/fsn/8mdwoZxeKKSGIjFCrSqQxJB0Iae79+hTS4ki+H4tgtFstNEVPlTeVr7y
mRWJ5GwmHObfQwX5+LMDUfLB5snv6YWlYqOTd8o4zksZhlxDlS4M6eFK9Vhuk8AV
WlDEY5dN/HqCh7knqL5gXXnIRDbODencNzanOe0z+5pGDal0+/udveUmlV5qezjG
HmnYb84SkwqCK13NVK4q5KkAtk1gt0DitAhb6zTpjWcpvcebWr8awUcjj9ciYUP5
P2pmK2xlie1rXuivhyoUKorXUeggk9wtSHYgbij+WB/EFxZqbd5ZmaWgpXvOun7H
Fk/9ysgjAjUzhr6k9NEBMB6lHOg21iMB3ofIm5x8zaSxnOOkoSIUX+WQ53YZa2M2
ZO2OsIp0H5TFPZGHYP1sU5+9WVT9d+CdgyWLCR/dNQCGbsaN++U5Eu74NdIcH6wq
0rlLzhabETq4pNR7QpmIWpnSFODV9g9bzWJrgYab/tBb0oP0IPdQJkFwSS9AFbLu
+noAsjDNfiF+dNIIEGB2nMo76eAoBBrObjZTZTjh2z1svIPswIrUMwLN0ddBrCWL
jCphHx+uI7rkOmaGxPH4a/UZ2pMatEcurYZHtUxkGctvWH9d6xQ7TlGR+JKUXopn
CBByub8URHkku8B59nuK8lEb7/v7rIQRflxKS2mYYb3hTSHS7otB+mhFQansuDjK
Ss/BSzpC+knE6HCLpTZINQ3OzToMLg+CLUvsEcjjfz9zwnlJGvIzd3W8bBog8VE4
PPFUg8GfAU/mUrzQCGpRqMqQ0LvqG3ba4/+DtaLcjoY+Pf88ApGiz4JPPyvdVmmI
MrQuEpOfKwJWuNHTDyuZiNRKpf+Bw1lkLqz60jEnVJQguo+WsuEmXuphL21FL5X+
xdv3kCBEPOBH6lqNlGED5sbcsLTfWlgYoL422B3aZcYCl2E1+28VyxZUTNT4EOQW
mCfGBGAHRUaaj9P6b01YmA3R/E5PI6rPOB+d4JzyFU4HjrmDbcG5BL3RaDDP2WsN
ji5hLpfh2CrtCS/kUexvIEFA7pkGWJ1JUYMBsdg5awJyD0/rX6pOE0SHqrtHVibt
eafr2cqtAf60ZrfrowX/r5o7x2YYH0lbj/oTf3/HClWY8pe5k17/Amrv+pCVeGb9
uY+l/Ant08NgL5BmxHRnLDb2/ZXCMjKS8HBwVqNLpxXhXJj9803q+JGuHqYOsCHZ
p/guW9ztGgUPHLgcZfiFmDdMZLvwVwuFdkaVL8Ptac2vNDEYLMPIMmhygG7rayz5
DXC+NNRYtN6ZXkS4XOHkMCoxUH6l7C3PQYY5L/1iftcT8WOIejiingftBRWxEuNe
AWKoNLb3iqHQitKDcWLrrqijDloc8ZH2qq1DfBszbXpL/sZl9Y572kGkj5iBD7wB
rXinx9tiV9G1LANCfm72ZJMqq9AlablvxN8qXTWvjxftOWVnxQvkcsIlY2nB7ahO
co3TtvpiDsBMHPpN21871gDTmfDjvNiNtmAvdwo9G0ZJL+rFTG1q0EmSs/3NhdRg
XbB7MYRVpxDndSpq1O0MG/KtQyiwuIM2fH9e+G6ze2kvXjYjKySp/AQaHf509qP/
9aoAqStDjXUnRDURdP6oVBp3NtVo4KTsvTepZe9umLfSHmDkyAjgzzaxhsnb9zMG
rBg9J4Ptgl2puNTsVLKYEqKt3cSKUNPP5eoGHIYazH9+XnV32w8IF5o7LK2+lKmn
vwngQqoi0gPnQkqbZpo/nTUB7wrw3Ti3X3nwV589/7poVWOTQxUiTXUhOlzm6vYo
bJJIJTcXxEunL2Bzc942GA6VdtPJHJcf8hVyeXf5wzlGOQ4YD4tyjoAD3aKn/Ooi
4+yAG3ZffCINy6Ypy3h6ve1/D+h8ncbPpbow1siWb/X5wDJKA3qn0+L8y8Kw2zwQ
Y4y73JhEjxH9RjHlM3E5VMPNV0RLX74Md+4HZ6nWz4UfJVFpp1kbwyYk/hbuhECu
712W/pKGhXmZU0p0JjNtbTUAh3MBjFEUqphp5sJGRfgW/4eypG3FIlgPLm7U3Qvs
HKMU/Yb36Uq5HDvN0brzt20yZRTE2uVuNE6w6/LQQkIOC6NVZEbNgo6p4y7vTSr3
yRLHn/Gdm3RN9s7D/KzNnNexvCKmlX5Glx+wF35SFANdfSaW6YDtF3CRvJia7yMp
Pd0+omRpw1JxXYe6T9YCvx4Al/vyVx4g2itab8b9YMDd3jwk1UPdc5qsRBo6q/Yz
To2HlDZ4F59+YY04DpezxTBjC/URQJQWuRxT5gPrxl/IgOs6y7SFoBmKfsl+ZPnF
CX53ItT8dnMXnlsfP/G+uvaQGhrtGIzWb5B8YdUkTi16lt+c/kyfzGt4XAe4npRH
nFD5B4qLMZUI5HvCWg+4vMq3DhjBxj8VQBnKkwNRnOhK1WsI4sBdHXrJvll4Qdyj
Ty+6apxBzPaTaMAvuaG0rbQsEbOemJynOf4TGMRByzOVpCAl/0voPSf4UQ8kqpwN
wiZgtSrKFe1NmuXc/FPkuB0NlZ87LqYk5Hd5ZZ+jpQ+9coTLJDYK2r0vjUDSfuLk
cZApCwcURXRmdinNdWaocNqa4PuNA03S7fRnEjIuY0ib/jhdbmM5pi+pbZhPX4zD
nyVG2P0019soGmDpIQIaJ5UaUqMpcVJJyRPAbmGYgPJi4SPJ788so/LXeW8W2M6k
fosaaOtqOGUb9CpjgX0ioJ/zZhbKpMZnhh1PM26Yw41t65oRjvGljCQNYVkEs9P+
SPdih884iTXFK39CsVJG9sUvtNtSFqF+NzT2/niUF7ZUdc5gTWIe0EKxFs/Xd20a
we6fDB4qaD0bZ5137UymiPgkp84Dfpsxt4jY7ewPwuLZMvew5Ks/5UdOBppUJwKy
ix4hHtM+CMynSKMw9KBZQ76QK7QU2/UX87PCYKjwtVaFnuC6F2DswmuCfEGU3/yx
J3nnA6UTYQpszOLNrpPW+PTbRYeD6X34lJFgqrD6LKWJ69piS/Rw1XYKNYTzrnns
lO4C3M6wI6u44xDkzjEN4NlUtBkXogB0XU9XM8tyC2aP/LlLHzw8LG56ZL4mg38o
TK9T/o5IPP38Sb2XyHJFhz4MnsE9kzIFZoh9Cu6BQyzVTU9yBJPcrfScoQfoq34V
PBETUkNiKuuA1JQq1Cb+WrgbHVF1zCkYlASiBQxX/ZyZOm+fVEU6QVdA6sYjosvM
koVRCxVVJIp/x216tWeQIqOLurf9QsoRoAjgRdJvpc/B6MPJ3mA5JOsg4oLKsKC7
3+uFi33jyGde2ylDyY7DQqj2DMF8iOU6ldlGp+t6aMNbiQ/jYSHcONVN2AOeXyLk
g5Ml7gNHx2qikbyp8f03SLcF4lDIePv3071cqGEBpSM5BNNrVkjx7XjyqMrkfxD+
QhHvNP9f2Odngj2uZp1XVRHNd3SBpEMYBuq4/3kVRW5Hj1i0m1C6hGnWfj1eReYn
BSLRpfU95fXMyV5zljxnrHkmHrnq7E20XTHPt+LswsH1XckBc0QOPoNIreyZN4dR
8c/L4w8BWJB8DoLIpa0pQ1/TYJsrlOXg1SqI/SE7pW1m3zbOs1gATpeHwSSLqhE5
wLjPi5rQbfHEj7Q5XFViwYAwHv/WpbJyDgSWF61sui4r800wbKHMURWlMrDAarRd
j0KjRCzur6CuKRTh2J2K3xlr2mKTwbn5ppc6nYozycop6IZSgDi/jfYv0CtllM1W
hDBITEd1zsq0HpeY3RZpQZBgq3s5rf4C92IsFxVhgP/lCpyZ84wi0rFMt1DiVQVQ
OwidyH6u2Dg36u2PcGh91xbLBf0XIH+2mSTHV7s0+TLcKvaSmummF9w+YDFuMGS6
vHzXluWUwMHO73+rmvJoTUi05rIRbhJVgyOAHGRKUw9k0IYmxjWLIx4t5695Q0ds
JdM2ZhKXziP+eImiBUIcnqp9x2eb4VgXNndmwWojXrRRwlauAJnPJ8JSGSXdbMg1
cMdvmfZKs3RKHk1msXwjaZP3VKUNWse4FUMGjz1b1VteNfHv04gaei+7FQzNErCw
8DcKxa8qc3nrGm2BK/XCHaTcfzyr58iRHwkZMD+RcEHlySXwNgzi0U1+Q5Sx4qmX
eYjuT/qtqUmmDX7I42imrcP9P9mQZIuL3Idr2f/l5i8SVS7RmkOOnVAqtjis/rPZ
7EvOBDQBFOgS5CW9HZXqgZ+Mx0xUAgZpwHxQ5ZmfBcwg2ht8bvQjaRZWi9GciFyN
iEE8RUwIwOg8v5h4diVeOllftnA8CS+bq8nqpnhT4KN5mYXTUN6Rlh63U+UE/AVt
Q8ORWyxdsWYEfi029eRPa4GafPSZcenN1l2EapJlLp0A0VsLkdMUdgMYi7CpNRI+
dpA2AIi6Mcbw+TduimJDclzIsX5LegrHdExF2FIL4GvbTrcLpHMnp8l5ueRSLDsJ
L881WKPIHnajzn9ZMXUDIcTqpOznmmatGU+PPRjuQCYhKTiRyz9jNMRc2U6xdl0Z
BhSQ39QqD/HCNULZ3Q1To092fPmz9vw2iJ7HyabyEKMUIOuJOMVdddBYXcAUkzJT
06NKH0cY+dSh1uyU+nopjUE6vLWD17awf1RiZIT+p+mrk10Z+WyO1MF8YgKeAknQ
krz4z53ssRUkw7V1TP0KebEa/2kVG/aQas5BdYpKTVBeLxP2pn1OGXRFWKYuIsjW
jQboEtH9jafQaeYEL6H7hey0seDobYeEyJlmt1lYsQWybhEVAr4HxtYkawuwstcu
acZI6BqANVg7U5VBP8jYzGrZMdaZbkjHrtimYdnsW7OdROuhUh0iqlsYQeAjBK3w
rrtc7izk/Ufz82sWTLAWWmg+499GOY1Z4+rTdNhe//TH0o4ilQqRUqSQjuEpjtsr
AedSbXz/QmpIsbYLG9tfs3ZKjoxikrlATA34DZTs+CgXV1N95Naqk8P7cgaYGiNn
6/EfVDRupZgblOoxGaDFBBCzjrkBGlwdGS2JlbM5xtSR86/YtKmep0U5Mw2M5rz+
P9xUpMf2lC3PgVTEsWU37qQmh9m9V/5LLM1tuIm7dhQzuHHkcSXUZ35WWHkr9N8u
tCbp0yicK9AWa4lOjOEOtgzfLev4mTph7XQDySWEfZBm9k3XA6DYGhMU7KZ+5bh8
GN0lEPQnFGUVOenAA6tLbJdwzoeY5kVq83JFjtsm6yth56mIkiVRplgwtAmarvLb
F9C1PkZM8MjRnuzcIOhSTaR5DUniy2AbZOQJPixSKX+cT3MmfpXMrIuPHFJJAxih
/A/sPIYZFjIRZonnoyJmih/O8wmxzvA8FpODYEIOuQ6DVeVcu71kLGOC/C8sl2kU
nV1yS9VnVrqVjYGa1fcYjvO9C8hl0TIk3BM40OGT5FtaIHhgv+tM5vqbBL2T2TNh
WJJJwsxuPxc+dL1dxa7yn7Tl6dXHDjhXt9ipfXwpwOiJP/6KqVO0Gdm9h5AHDflh
gIa3F/73rQWMBvL5ypr9IR0tjlnlElPCqmJr/gVyUC+M6JrF/+JsQtWF+GOsspfA
omzsAv9/lMGVdYi2mCXRi+hQ0VRFQ3EI9iNBPn/E7AUaQY3pu/55wRuV+ZUc6Tcp
q7uqy2fN8ibM/u8Epoz79p8Rydr77CqbATCs3VQju9opzLnYZVg3MGCFs84K4iYP
6cun2lW1NMTGREI+73rLDNw+qVOJLGO+peB6RgvUGba+DsRG1Qnx2TpdhqBcdsHW
uQHaHO0qMM6XaAub6w1INjRJwte3w6Ch4lIiNuu4odkKjn4kybcKacVoLfe0I1W+
HvxK1uVBaPsF/ux/8QIks0uIWTGPk7rjm+aQUn6ZJa/LqVUJkpSzb0ZtbvNgf85F
opICooK3X9np8Ijln6TVK6tt2ObSm5H2u282uIW+OB40rtgtRyfIiPgFGIueSxM5
pEl7PF7d/aqsZcssO2oiSTAJX7y7XXohanrr/ZG5EwpHZGbxPx4WYo7JdJjIVYN3
px4j+k5tYslKbY47A4pmrlHY4vkK/lPxJQSha5Ku57Lj8AAVBthDIpt+m1Lfaw/M
GEUlCQR2O1MKyGmuZQsFWCsEVIJJ82oOu5vBDXdjEPYRthGnF5IkteuWcH1XeLHi
83m+BfAWAqgIfNBpeL8Biwh7Ce1u285Sferzny6rbHf555fl+yI5dt36k1FrWQj+
jxKhZiZiIVhBAXPGm+L8pGSn1yetXNsUZNU9dy2TJ4sezPfoYbW93pkBuV72z/QB
iphbHUoj2JOLq5e98gpZx8c2Ecf6oZt/8hDbM9XrYK5WW04LfkaLrz5iAjwpc8ho
mn04Iu2r2PxSFV2d/R48yCoAKIRQnlHjAKbI0kXPdijA97TEMK+otz3xvlh4mYhy
TFfzeRLRPFzwhcL6YzAe2FKl9aYlldxNG4UhuKA6fLop8+Zy8B4FGdmbu1T5eTpv
Ipe/XkYnQhDaU3OVgRY0rUXxZrVYGYcp8Zclhz2UNXll/bdX6adEEAS6Uurltval
wDPTFWn4rkpgdq4wAzwVpTv4HPJObXikp0k3LP5yaRDT0fdjFG9KM68Gpu8DPvdT
4RL5lTmMlMsC2st4aMiM/3YR61jzYKSrYDFEO8YoN4vRCGyiq4grMkGBft2QPw4A
WpANnjL/xWdZKZOWvMNLQ7KqjybNIgvYyEJ8Tmy7RIwpEXlAsJpNkikH3bS+BYfC
ar6oyefs4ibW2rYsfUr/yeVhDq1IhdzsoP7MkHp3Nw4jZ8U9ZoeTa6Y/HXWzdHPW
LbTAPo7KjzXfK3jAk2tGIh0AQlDF4xiqbRqr++Z/G4zUwlmkF50mzeKq+W9MDvjo
JtlXhQToU339wl5wqT2qivW/haBJSLukg62k583k9dePaISb1y2Aw8K6+8L80xpn
PuX/cikbf654cmd5rUTf49sHgeKK+0N94anPRrJD4T8cIgppn1MPNxgtfRxpRcnQ
3lP7/qfX1wu9eHCnsDNBO+6fFQ/ZkEF0tZ1L0bpzeIzqsQs7snLHTYrlJlEezoyl
faDBZLJtDssDME8APBDQaL91SqFUmZoCdU0YKuRy89iRduOx6299uvbFRWziB6kn
jVnkX6N8bFcabHxw+LTT0BdejkrsPpCfxPli54lHdRGWEPcqptKkyd3MaXIMOk59
Lv+6bk0Hy/Q3boW9kzVz6A1Iyi5fTuOABPd7/+jzd9PIby9mqm6YrTHxyu/yNJYE
GKOyJNdl7Jg/Pa5cmCUe3TmeLKQfZ8fm6xlv4QrvhHf8zWRW/ua1/JVpxSwwHw8A
Tis/ynIQ7tlhajpPnUwDl3ReE2bvGXvRZLEKFh0UGwdMzKsEFg3JAYFcT1bm73bR
Zo8bOgwJlDmnwsavD5ZiBssPlYozD7/bcWOTx5vCl0QyrPvFWQ3BrOxweANSkVVC
vM2i+oPC33qWOU3rz7/NXeBI91llJWIyoMRB/K/aBN5hpMoQx3B1igW5T5JRxdhs
3YyZpahM7qYTiwn+T2gm436i0QzyCYToDntFnMlEx/MdvHZ3Qde+tClYyGkEzR6V
FeMwhHhHOZGL2XWELKYmMKdCZtLXHmNHJc1Uxw2E7h+yLr9tWsPwso4wOQBqCUw0
i3fkECaj7vqyyMaTJJ5kbYDViPiPeM+T2CyntyVY9orggdYMABYKLrEwvmYwTP8n
w5mgSctVFoATKCe2ljZI1n6c5Vm6dHZobF/ZT6xjgpElOVfQM2qDl3OEligbtqHg
0vn5/53ly1JueexErd4ABApntihkI46xqddjRHG0tXG8bJLDFc/2wuz7WKEHamQl
AXqQRvM5GlLA28YD4WvKIa/UHZee+6ApNl58AQuaJwHrK04U0uiQ7qYREMkEm3Ee
bAtzBA3JBI+ADEgkQhi91Kjf1ZTs/+oSmt3KkozmLk9uYQ5qnLD3cNojeUt2r1TP
ujrfW3DEWAFtXptjCI/zCiwdGyp31lY40/Lv+VDnNgmPRY8/cx2NburSSPM9Ekbx
s5jBmcB+/sL3UQJbFfR0GBJS5z5fx+2v2k4B4cuSSorDCdRsPvSkEXjuifYCI8/h
E4hmFpgnQveEpzFjqc2vTxQPTL7icsR5sHbr3R94aGiCxjiS/XTrB7B3Jg+SC/Dd
od/oDwosxzkzF/MKE1MU26FUh4cz6tecFJpT9Qw2ZgybL2R3gMCy7/UCehMrlFYJ
5Uig3YRDR0QsatJk8CJqEFmstW1awjotXkdXeCOoyWXh/68KPasHdsoHMcBti7U4
dZy5oI3jM8HNspj0jPv+PkGQpS4JpIy42elH+eBp0ai9jZjB8oqqUSUl09A2m8i4
C96MdXpbp/nmGIbXBIEMgq+ablcMJGvRJP/BTcO+xNesW1DTzezNpQlGwOmHZjDl
pH97d7cGogBzkIEgn1U23lsV8r01UVY5NDW+rejBmTxL3iAAzYa+w3nfCy2awoEp
UTVUc7EiuekoXtqwryBsYjZAm5TrXIYfCgmPGzt2n6uDqNYm+x6IJWpEooePPOzw
1G+yupWPfhFCtS438X5gdUpa+H+cMylEupW27cmZu5iKtmep5FCVorJhn40gtADG
qrKRTyvdF4OLO56qiXeSKUZIdy5pK3QgrutJdPJ3qAdnhk3E3EJagDwkcwIH4FAb
4QnXHVwt1HjfV5agFli7qlrK/wa9MsCVLfnFLr1wqhjn/pyM2+UXr6H/FiE38L4e
f8W9LrJpW+rEYOFDDfQOdyIxn0nAQZO9DYJ6TL/tklA/brhIjKnV4H82gUxNKzY1
QvqjaKd8Xas76e4Msh2siUQpiV9qoL//M8Yms5BAqpcEZSnhFKjtw4sG+5WO/45b
7IeRJ2aMjau3q+Vn+fB/pN5ye+cWNOljTW9KSAsJhgPzM6BRvmM0YXz9jDLEv8pv
V0PitrA1s7cPMrTDWzjl83KimYZEJD3C1PSM6bszJ5+P0Kve+Jaod2uiXXdgtlOj
uYaardciOkB7mkyaXZetQjkC3k8QXmtU5hlxsaZRj++YxP1d1PeKrEcEKMQIV5LD
Ls5RKGXdfz2QIkpZ2h5mpwBNTRELHwVY/m1WQyCNB6yfYVaAhOofwn939XbI+9nY
3s+k6q2TeAK3JlMBTkMt9cWijYTh5QIYGnWXDF6CIEdZrDRgjeqwPwkULHOOB0NN
iI8X9QLClt7+j6FZfLUpFmLFu0wFSYn0hjVwvqjl4AHDaQOG4df/1jlr4F0LWPun
9VMJSMJ3DpLr5xmD7H6b2ZB6FftXCy2ieq4dSVL8hySJF8mEljx2uTmj9ne4lBm0
dqtlTskUBvoNkDXQ+R97Zm1frZz+LhtcCt0130VkEz4r32e6nopQUF9Fb9DcUZfl
EZT5WmUmSxqTGbphxvtPVnDOPJur0P0a+KOpd10FO6M/bMVigAU9EPiwPSx7jxW/
XCoutrjNxJ940M6ER7oFkKiYpE3pQO/aDpe4h3WWZTA8MaPOppezQwE64JRe2gPQ
Er25w2/WNGyszH1paTLPoQlmteouQRAMbD4d+2BKf81JTqF4fezgImLhcROzVQpz
mUqFdfLzCoEmu73FJItDgIyEZ7M+0afjfsrjP5P26TVqAVzVY91P+e8+2pHmmmAT
mephJ2gWuyf4b/lqH64P04kD5MUnnGZtD9/ie2KmSiis24b3ATZxpBXHl4oF/IKd
edQ8ft9zlc1olz6U384Df0C2CLbDt/5ZNSp4bhqZ8QbhNxNdo/3q+wwUwJF7WD1L
p+Xqf9jU6L7Mm6JOlDhvMhHS9fJ7MgRq69bTb2eXG2qNIlPOsuE+Kos6t8EpJ4l2
mVVw6zRth0cKe3O/tLDk5GSrBC3waJdk6UzyPFsXFgoXrE7Aoc5mcMyxWP3RIDs4
MdMtk2dlsuZ5+qs9ecSx77Zf4mmP8IdVS34mVyhyHjeQ+Y1CvS7PWbJPrEefedH+
S7UHTSTswheTAYZss7A+lTGW+IW+P81LMkwlTJr5xj7NoLTPcaB4b2hXJmFtNlhA
eXgUXBlvwtT44op3ABcRdTf6o243HKdq6KLxqmOu3zg2QsDaY59kxvqZrbiycZb8
WZFmqw32WI628ZfWFSOrwPhgIuFVjAbPEAEs5LavRM76K4IRt95VMhyhfAuAZfnh
/vXK1zkrN+VcBIf3entN5H/NdJbWAS5ek8TFt4fIrFN0GKfrv7J1dKTcrUZ5fpLp
6zXZpkvq8BkO0yWuFBPpYKmqIH+QTNMhl9HtZuL1PF8maPPp2GhiPty4ftnhUg5h
VFX2TCyAWckFQq5HHn5r0cJMiw3kgG2Hrp//ZoEg82TiBev/yBJEf2AgzzHq2bqz
6W9WBzCzeTZZ9juzL+d6Hv91tMalF6vnDhQYOvzXUt0CcYMEognhoikzH6RaJLno
Kg561C4L5EzpozIrlWZTIS3RhhHrVQhR1FHilCl6F9IDKhmOR/mr5RTb9XJGSg78
PFKEMllCY1xuxa2Xy3HeMQilyd1mKMKpHLLJmD8mdcTkabe1ZLEtOzmN4a//1RwU
AX0ELQ0fvUYxz8/TkzGoxMage7onLZ3D5csEkr2TCaTf8KxlJ+S/YeyJj6dYNEvS
6Wx5dmkb597qItnvOX2Lu5K8fOuuygCuA3Pb3iLcO7TTUJMjWt2AXRm6n5kpGvR/
0KffQr185nCgpjzdB5+0UxSaW3L0u16hJk209vJIdW1ubyWSdjBc5t/lhmfSZ5r5
fwaUW2Ovf9Nb0c4xhVF6vc2jwDyyY4/AcCY4iqsMAtNZN9JpApM2kogki99ACCuN
eV8DmpwVdvLAXRlJUKyngdYmyyKzYGLNntb0EK24eYqcfOgavo7rvSKLbvuTFIJi
g99iglJRgJkS3VL85Nscfh9JNOHZ8YFxHNcbgrtST3RpkM6sglGaCqcpZNkZYMdV
XVjwMa21OBemvT3VVbW+cOYffoRXpA4xLs9TlOONSJP7Xu6Orbg8xoeVKDO6Mz1t
2CrK1Qz2sugwRg+z548kWxpdYvXVOWd4lWuUY1fZDAdxnCZ5AzLZQiCO4X+k3cip
B10xRBXQczUTEfJp8oOCLLntFkaQzbP213r+ktbSJL3o17MhfsR3I48nx1tyc4sx
7B7rxxi3CpAU8WqYv09UJ2XPDIkzv5E3LNsw71YM9C97+c9BCMGmg0ZyPTR6r/7N
P3AYAPUzT2Yi0ME256ypF7/fOQF9b8c7z38WQGe061ZJSVHGZOYEwbRzXVXsluKQ
0A8BUeYUkA8yxxTRXY+yQZ81gg/Us+kiES8Nxn7iCuowpZWit8bwcXsCOIWzN4+5
skQDfunq2T4qO1oqegkziBTHeb+IYFHkY0IxsKZvnhsbnyWAJEAUR3ayA0cRMSHb
i8taQLCijyFJD4p/SNiKPSK8NMcC6meq6BICS4rT+Fi31YAPpvBTFAZh2ah2SOCn
KSSpevzITaypvD9f4PIAhJ4IId6Vd+tLFdCeOYKk0NLaP+cxAbZfjS2q5FY5BYtc
3VaidAiNAwlM3/OBE0T4qlTqkGVE7Tb5V6ZI1tcE747lgsEQGF5gn1d/ryZCcAKL
CzNUM1/9h9ALNlBpdY/SPGsU+sjG9zuJ4aAaFhxQCWJNxpshB2B0eJl5zVkQjSWo
ZfBWgxAqauxktuGPPZzq+8dTPglc7rauxkIVslfCnoudsZrldghTDnepGIJIKlxD
KCYnODVelpteQlWoAXYy1OBB4XYJAn68dDRgtFgLfcDC3PLDMxcTD2Y3pLBps3yY
q0eoU65xSF7kopSeXFHsGeWJAyIUvLQEACby37ihUCn2cL12qquJDNgwmkSXphIJ
bsHeWu2ExFhiB4PEtomPYviSHIwpNjodeUjMF1yWj50OwDOgr8GgcfKjco97ss0Q
PAW0mDCWNN3bkc+/OA8sJLkY5BQx7t8N62LgwgTgExa3Gv3w26GLkrBc0HgwfJwg
RV3qwQKtH+TowtCp6dxCh4D4L6oOla8Vyn9li6zaKj8F8Fj8M8yurJfXYhXaR+dM
U3JkHEHkPPTuw8J/8SDehxPkoYw5xwBJAGakIp/TbkeB+Wa9p0BI/mESKkPqFCyo
SPWAi4cMgEsJ7oD8ocpOWnmW2NXelP3mEPQA+mNZKc8nB/I0T8WoWlLu/PRBTnYb
lxiHvVJXAoStbp2MRNyhLUDKraeJGTPlItG0OCag5EGYQNFZ+Bw0+y44S7y/JUk0
+Eulbr2Vcd2/wzjmX6585HTksoCaZdae7QOjJbF9uB8wsbQG6IEAVq04Hh4hcQlU
qTiqkEjvZA8FMKBXsudyQod1y4EDkY4DXxur/boOTi6jvbpiVbN9c7il95gB+IMs
ZNcKpR9GmE6VaPVHgfHRAsJlQF4JLL4Ln4mSC1lK4FtZjZJ4C1scHwtBiEVFWnzD
Au4vrChqcHQwP7j8B2eS6tKcQYuiOa7igFE/12opvLuAJTLqnvvvnYXwZvMm82rS
mxh7ms7pN73AN4nrJzOeT4/ZIcD0eHN6V7wAAJc6fMjOhQK4BnEIAUo8UccWzdch
2+rJpj4/yp+cet956YQ6TJqkpGTVjzY0hkSXRBlpuY61cw3bywCr7bc/7YzvbXZS
qhTOBJwvLvGcAapff2oGnrkLH9gaP2t/IkHK+N2PljP25JZTyQ46H9G/0R42S0Yw
Hdz3Ot+2Okh1buUCLuIs+xEobrT9EVtO0ewhOBVgg8g+buatVjRuQZcV4V9IhsRT
+XxLjk+4yKbeqj0eGwxbdipZJiRjw0o2f66pmCjgq9HRWWQZWCYD1VOEfSlt0PLF
gBWmO2/rd5sT7DU66CJh8H4N7/OG1TjlZnJ2H3VtomvJNcXIlDm/x3oGphpyjjeZ
K2IuedvGahwxWssSTrQL7pidU4Ma2KDvNtRKn3rnEX0wA/i02YOEhN4tltRHHHpO
o66jzKzpEn5ozFc72YWdozJSPWNbY3Fjn/ku1IMWKc3VjuuWkiewkZ13QljniHBL
9W9rl/vGTYP/9/fSAKkcJHNdHLgV/kcvD3+lmxQ8PapEclaKxj7X6dT+fG1iGGmU
IOpDx548c3uuRedc6Kam2wVnEz3lNpphTpJj4koWyXtR1SSs0HSmsqHK0hyBfGjQ
Gs4lc2f0dNoM7rap3TOEWJWCFNcyM+OnLW+fe6ECNsr2Uocx6aSATLXXGFvW5ufe
rLdgFxB5f9yHmrNTTO/u3p8bD4lf+FM8hxDTky6KX1RAnwkr3DqtKt/ibFpNOFZV
iTdXw02yOf7Yesz+UGRgRwfxSHRUdyIrAKYw7Mn0Zv9rWf5n5FnCnrJ8KE7zDAKS
PjtKbH2MyMUROOaGkfk8eA6bu/bzmvlGQ2BgVC5fSXMMKRKd5abZ9XJ6Osj0Nk1Z
s8r/Pjb3dCWGvuxj6REmQ7TguqNYy+B6LoTZ8wz8t63ksgoIKACWajxY7imO6NOA
mkdVM4vnN/UBZAScNWIItp0ThMXPvp/ESVBo+nJThYlAg4xpJVNRylU3Mc/sGHU0
D9TSPMpy5TR/SOpgSSJZHMh3ob/VLcuC3KkYNsGjd7RxbCiI7sG/vmWDOqeDSDbK
eSZJgpKbC0M2W5PYnz2Svpm9fInmZ04cshxAX+fcfN6fC43wlmh49z/kvid2tBRO
ND4TPi/Ue+GctI75a7L7ci+P2fM0DXaC3kJK1R92pwpkxVv6j5NXA0H4OPzrtyNJ
7pVpJgcsuq7yXzCWonMoDthiFpBJKGi6aLtp9PHvN881oFc4M6hcG3QYndhEh6M9
ihruSfZDU0MRftSgZ1BmlnLNlnFfs9zv6TXOJduBvpr8JoyC2vmnBZPD7J1XoaG/
0ZirDSi40sH0KFvHxdZrXouIFexuHb2hQFPvXnadxp55x/aveVqjt13OcD/NRKUL
UfY60uWyqjOEw9LWIKvV8n/p1Tm+oEJZiYwB9yxHPEFmzAwrwdVP5DfwbcCGEd8K
7yGyFRdoL+1pX2ylzmBrjMObAngfDS3wnIBtYdyF0wCq3Dpu7ZThTT8AX+FUp06o
xhekrKwBJZoVqjIK8PiIJjax5EQbx/2RbCuSaN1IeIQqUty+OEkKxce0CNYFQt/B
8L2txywr+FnL8P0V67isaxLFj9sVL7alaLElPTQdE8elDFdg3qiQUn21pDgw+H9l
MMjsS7EJWt8EGFd9yLxuIGkbr7hqiYxnIo5zuFOg/5UReCEbNA61mF1vDsgbrW0D
iynzcGmoaR1jKHE3/HJSZmAbGKm5YBCKbmPhIo02ypAES2UTH8Rf4YxoNOnoQC74
/JseIWjTwPRm5rcOah91Ghx9qHWPgx619IyFuC+J+b99rASDvR9i96PnO8L3K9Xd
6Hv9LNwhUJCphJUM1L0CxNBeu/B6txXM6YiyUaV8gRGtphnrMMpdTWzLY8OZEENw
wgsPb4rnK/D4K5RXuoPTwK/2MTccc7xxGdWGF+Ob5xW2mkC490yxQKcFwnrfEoPX
no8sjZCMPkdIvmrWBPr7uIJTD2ZnRaWHHJ+6rLAd+RTbrOCP+bRnL4EE6CYyriHF
RMOV056EwM8N9B/wBMNqBgXH1orL7PBcs5svGhp6n3wlo9WB3cQYVhSzRw9g/0rA
PSeH2CbKF251w8XKfutWfZxeuvbyj+TMh8FJljHGDbH9wEwATVumbdmZt/17c/L0
qgZ0ZVqVFh0oFJflVt0/hnv26W5/4p3Qv3bk2BYTMWgT3cDeGHXKUyfOx+Grwd6j
NZhNNwn3GnbT1mNXnyUuUOUt8BrnVLOGimLZC10kQmjuCSm+9PGQFXNtC5Kx1t99
rJrQVrKR6r6xZ7Wy2bpwLNV9eGQ6EoTG8DI3leh4OKF/qB7Xx1uaFHtQL2eIHA5N
V9HdVshHORGq3Nl2zf4bCbfwAFHRhqOFdPlmY9sPv+/2mcub8c3VDkU2ZE7fxPRT
nKTqYq8ofguaPEs5ld17lYD6wugq1xkgcshz8mJ7iuVEL8wx1WQQ0IM0+HssMWfA
+jHWrDktQfnX42V9tt+IEHQJvH9t6kqGZgjgi9krr/rZwtncduYcQivxcQcFh3ZX
GfRirAdXuCgWo/i6rrduE10tsQZNg1RIDe4nlC9T3bfciD+sJgKixOu6ckpdSBZ3
F0AvEMZYZov3kboYFKH9H0bBFx6RrBoaWrJp0P7kgtAssnyDbUVuVVOf2fnEQRiv
rBkS7AH4yRia6aWgiNKHXQJ1XGmDMZyzW9xAmrgeYtANxpKaqfEWmPwvQoO+9/35
wFjSJK+ofe/m4VxkFWAPRQoYPUWWvJFUsGPvldI8DvnoDySHc69OQbmDW7HoQ+7+
ExvZ30rENyHm7LnFOP7S/IsKX4ywRPxZT/0yLWelt/+RMAwq8qJ8CGehKCS0Hy+m
7ETWXN6N0I2qAvXQ5Zu3kE91ThlpC+K7DiftV8TwVtAQhFSq9DTGMgdXjm2qU3s0
RC23QAIlS8qpZuG0ObPxx2quPPJBvBaUnLguW6spUyDLOsw1YjyBWYwCnxTTzn6p
W5v9m+XGCyumOmeAYSYIeSJ5EzW9dMpEO5PzUd2bfRhAFllh316Qhha5RyJ7NGsk
f8cMo45n6M28gSCqgqcVE4NOFZTGNOwjIltI9PZ63kgy83TNTqSvslRVGU7iDPo9
CFXtu5uQnPlLMWtPwlCQ6jN9hxOC6Ew+q/+BUqGiAsYdc2/w2ITZFsfmw2CWlr06
Q96CKRlKM1ZkwKp1cV6Cc5HDWKPOCI0ENJXnJdDq/tjtnidww2za8klPJawsCXRG
YZxRSsS+gycTuZpFsIdg8lKu2CgGA+Kf6P0WiLiyhiwXxC52sROeq1Ecm9gfJ2f/
DbyuB+fPgZD5jn2Ng4G4CrLwbnOH44jW0jqvrAEjeWPGJpZjaQAH58mZueWOmotl
piT15vLNT6qPUiD5FKmcSwOKTzL9IF5nsTvMYrQYfuASN+daEKVlogmyK6Puc9l3
ch1xCBXPEHLKyymKpk/lrLHial2cgdfFvMnpIdQGAibRKaWpMjlpaCaWz99Sfe6k
nKZ53airxKWeqBdGHKhyUHjaEg2eQcD76BvBOFvl3uJcLE+yFbGJ0naoElAyQtL1
iShF9mCFl7Ph1DuyyqtKVWsaffD1ga+mYjm5am9aCf3Rq4grU0Szo0WaQksoHqZt
cYXgFYMbjJIWKTTW9w94gdHA9UFfYhP2uGxeDijyxqwJyyuA7atllPKH3z5FidSo
Kl8bzTOgwT4q0dLq7qRB9FaoGmEu826h2RdnIyeEt9u63/4WTc3Ivjtqn0bL3lTl
dObull42UA950/XSDjsgFCpyMfPJCRvSTwk37Yp/seyQQmDHvTTimYfVGiJVIw07
wygG/jO8vgtFAA7g6iCT6I4Eo5G2Gnz0j6jmkJjxj7dFhjtNSs26x4/Ah7NfarDN
S6L8kC9my49VWALl3Fkr0MzGlMyKrSEsakCgHyV8Ioo84mgzbRIQ80wIUVh9g2D+
nHw0T5ABOcKV70Fkse1uWUBM8/Zm4KVgb9Am0ehSvBMAWoJQ7BIwWhMdx84L7mtU
SYxjVXztUkRH3KGgtVd8fA6R4NU3F4OiV14Lz1DVwXf+MEfyLs7xVom6CfdNn9/N
D2dwuM5jmP49fzHRudiJetj73EpkbhKV0MuGIn0pkBJKm6Wj5J6LqUPODGuppSLj
6PsDo+Ki7cfNWTRkJJ/V5gKrdpn2aNeA2m1XAijWo5wGLaioR54DAG9nN9V9OuqY
4fuh5Xl+D4LtsH08rLg5RKpYPvBMYwg50eK454OyNM979tXHQBa/sdqUAI1G3j2H
swi2oT+2llHTMLFJAl0CaWeeaMPbiPhQPW0DyOIogD0fWaFowNhWDJv3K/QL3nzi
m/5lfo1C/SyDIT0hsdapnoWkiYHYfeH5fCdlVkBEcmREwYTCvGtCo5OyAbqKmWzd
jVs4xxx2+Mplbgkc85G3mkjwEqaysqn9Za5kkC0gjKTqXrnVW1tEX6SRm6wpq7YY
92aa+Ix1JShc1SnjDG7HtaAUK9W6NFgQl2WW4w300HQKXqSkNxWJAG+4xlvf/flM
BBF7apdjJbGoIH29oYMlSN6AJ7u9BUspWNTuou/FSj+gJxRPzNwmEmmPSPQvU1EK
4hvOlv/FPGMWBI5fCQ3SukoraY/G2nrm03RjEjduF5xYwjg3LC7ZED0FSpaNyPIl
Cqizd8ojmADQTcTKyh8rTlVEw2347mpVHjxjRZVD2HMYu7mmQ0kdKz0G9uka9vRv
yTkfd8O1FGY/kPo9A7YCeLaNFhFDhN8IUQXA7a4lWXW1T3rOaVLd6v+yI1TIn5ce
b16ni37eZ5C/cM6szITxVfsYl2YF+Kx8favTarVWgDRThHmhuS3ruXoCjSI170i8
Gd9IGZDBtVe0Pbp5M5FXZQVkhGbaG/JpgsDv+3IH2sMb9PqCm2sH2uE9wRC0Zhv/
fJ2p9QhgGRFO0cvlBvbHcy/nYwj2Vp7YtFowhSWWWzwGTxy4up2spc3v2S9jdAu2
/qCLN4p0hLTDC/cO6BB0Wl6XeSO50Q/6BIiF1MPjInWYVisqYc45Vw7WqA3Iisy5
Zey1PmxxI+0v4zV7FC4nD3vhFstSa1AOrW5itxOscEdcnCJCod5cglww3KClgJie
7jMl0NzwkDG7aUGSOFfg9/IfHmthpzWgKJ6Vrj4W1ODtDYmmb60/CtvUsO5IHeIQ
ZFVFZrsQS5JEMefOmkT+9WDQa4ogDODzI+G15VwtDZ0OEaXpfKDMCLidjWJEPmef
KzdcH+9V/Nb0vqWTjWEhEB0DG13TzCV8C+sjW/HJGXarVKxvLZPMVJ9nuC0uvz+t
1G/O9t/AXXNO8vABKtV/T0Ei7uutmb5eISOTPW0wOSsH1yCB6I6/FFtViKk9DHp7
Uls3WknR696lC07/7wFMzlRJ0moFsjr7v0JabBObjq7tkKTlSYiu/VuTQKcUrjC5
tNLLg+UNmu0wsw7V10aMe6+cV6qaQSJtQwa+OkKUB4bIxom3SXTB1pp2ps62qit7
yVM8jWWv4woidbhFhPcMWKMPdrhCCvuz/2PQcFOPtjcgalY1eWr5zpm34n+vUdbW
/l7Voc1tUSbv1zHNVFOmjd5+qrKQzsJe9eL3XVYUNs2iNTgHgivYMmi2s1E9R6jn
LLX6lpxH6vM8iDscVPm5wkkKV7dilBNah+WYv0NPlm9TE+JU+zaTap94YSWbMQG9
5yEHgsHVjgxHK02A7SJG341MhJCE2uUb+cxBI1tS+H75v6gDA8r4owo4FSuURMBZ
fRc9whUWjxpqAJc9wxWUkynOYGHP/quvUalpgiAakf5qK8SmOG1tByqUZGqePEzj
fPb+DPtdselN/otSDD9W65UREQyHVXT7dhgX/SFxHePYkGMTo8CSd+JvV7QCuUGs
PGEInnq7k8d+TVLMePp4J2m/HpzMWcJGz7k2Acv1sdu86Qns1KFcyxz22SFZGpDv
KnJ3b3Cdp8yopLv1zb8eRZsQ6PdFaNCBXQLudR75QvTrqHOS6Q3gDmJZpyhWtGDD
du2zPRaEh7k1HDMRskxgYd0rbdWgnY1Vb/C64xNCPsReI8HDRvGTEWndbveIFvEM
w4Wv2dNAgUtaP1W/LuMCsniMe0WVx2n9WjNTiOmJVqforovOmvdQJ8Z1dpnb+YSx
YwwzHF6u5gmDYSpoVcGXmNJ2deoT06Wd6Np/Oax7sVC0g8vzXJ52YPvrLH9rHQ4x
Qqt59nq1U+nqIV0HxbhTMNNUwBpT0CSnWRZt/OKtFiH/CSb9u9k/v1YmEJxAHWqr
A+2icQzx8BuntkP+B1Ts+7L7yVFsa7Tfn4i1xX2z2Ugp46ksEKDj0hxAmBpcdnwK
P+fLoXNPuLNpKCovEZOHvbrWTQBmEvyVfctM19ssrLDQXKI76lnl63E8/amr1+8I
6hiJlFvZNfYFRmH1ozaNJU1V8+N1jyisH2/BP9spNnQNppfp6LNcgHaKlyTpZqID
uA5Vh5z1oP4OFk0oCbkGnVH4UsaMeu+ZOVtBp0B1nSIT6OwI5AaFT5LNy27F+eCY
lvnkHg1loMvxzRztzvEfqSntQBt6xXW4DRmFVAkTs8bs2Gxg+cpGiZOE2TMXZwNX
bcVWbFrgjoqHr+xyfZpSmBePZ6GfDqdTe9sBQS4PnYh7MHeCMwTb5s0IsmvoFVoj
YLZPwtgjWiQ0TWuSi6hr/QIHUfO6Pjl96BrjOjkY57ytman08XiaVXzw9v73ArOM
iTTYWfbbCKsFzb1hkLaDthOc6zX+dEsf22mcoDlRUiC9gBOlPU+9hqeMt4VtW4fy
Yz0pZ1fA0vDPEgcnm6FFYC95VL425CKTyPauOJaxKrrrHWCyunsIYkFL58dvNXGh
PB80nxJwnyZxvquXPGbEviky51cqHmTDYQNzNaah/2NpvXwbaEqxArxwms4ul/OB
DsRzdYO3vXJiap+PrwMvuxEis1OAvHH868RLLzANI/Ia9ZPk23d3DyPADX+jmlhu
wvs0NuIqr5NvC+oZMnTA6wAKRcE3hhax5BD+K7duC8vClstWn0jZ+sal5E2vbir0
TPQO/j8xw4wxN3mC2YmGBdGDkRDH8pDRCvaxMU6BYAaX79ALa05ORcriQ7h35I5E
Az/XN/4v0jadB7tNYeriutFKNOsFdfisW+xYjzIpvReDGTItRdA4cbILBUasALHS
39bXu5M6k7whqZ4Ccn3WOuspBDZp+t/lFc9vZpHiJk9cCSQIW/ElHkInm67KCLWs
ohwk9wSve9Y6p4w6pfG7Rf/DEj11FbybXPhDI75AzjC+nPL5RnO5no0sEzSHD/86
pOgKwa5PrwBuUmFty8Hca/ODdooJ6MeZG8vkdn48OTE1TRL5Jjz6gQYJIORkhoeD
hGZC60chNorKbOjpkq8shUCRWTBgp8nSAuk1EKzQDLy2JSB3RHt1/5V4K6v6bA4O
fH7jKvwEyXEKlEw9b2EbsvNs2FsB33yOsUvRSfTe2gQSXjy/pWUclS8oQUZhbv/c
W2pztINfMSo/xN+DdPF2DoW9B8QiiDXpfJDmsA3E/NjYpP+gsSjvwRObjB8v3k16
MZOmpD6YGW9ZxVm5PP0HQNTg7sYS0910wj5r79b2X0zQhBZK07LkCnUF47uvN+rY
xv8jR7SPElDsRToHOxl0sXguy/65L3N7aIgoBPi6SQ4evD2geccMAH0+wOUPGUxb
wyot3Pr/ie1doAgBH3jrLHG51xzLHQ2NC6nvBdl1voch5KABA15afU7uWE2L7RSz
VQJDUTOOV0Pt0lDVcDLjGG77MgQiS41crruxVQ7coouYhM8gengKSZNGvbXaz/or
x+K+CH51IDfI9X8ufNj0MyeiJZgAcTbtV3gXMe77bBE1fLQcfdccATHNBwgv76ro
eQnT6f/nuvaU4bBeWRvnvUbUtZs2szNSmgbBnYMxHxl6eLfN9Mub16ZS/8/Lq5WW
4Z65Tui2wHokQjOqOSyHiQLw1xzW7IzZnOMmt9PAnAJl2zzRkC4QyxPWMrAK3Of1
y3z4/ZrFe4Ro5MGik2+djIHX98BE8WcghOqkGhbZrTKBCConlugliDsU2GcB1kMU
dFEgKxQLuklnrLKQ1nBsNWPpmgvVrjhlr+K7F+NCoKi4Gu2J2ns9nSyd0lWrQ7ZV
gzyIdO8/cIlPozDHUbQY/GdvjZIZONPLIrhinFuB2VBHkMPI5RgdKu5FdPWeb+R2
pIV5+WmOt6BnawhyvJ8DeKev2Qz48QBqwZSAzEQvymYlLJLUtb8G+4Pwk2MG1cTV
UxLH7vLmIt6QAbRtT2SQ2kqZcNp2nVu7p1o76qObT2uXkqb9p3Uwz4WGruGv3jCE
35BzYigKuLAmvHZzMoPGHTlk+0YMEI1aNMtk1cV26QT2M4o/Sbez5reZGaa3AmPo
cSGrkfAMcuPa09pnuhB7Cy14ftLoX6fuEh+CZsLTPeHeYpPFvKfQ+FqhFiL4k6Zw
f+ixGCw5kp6/mruiYpuPC7Ur84Hg+ci98da1nHA9wJ6S5fCATfg1JAabtxNiKGIb
qwDWH64r+5WEMuWlX9bW6YPLR8RRVeSvqZbf/cPCQ0UtvAafDRE9/NqDyyDJXiDy
M6j5W0db2OKMuwTyNn6jLzTHiXr4aw6kbc0ukAybcmnCmk6ull/Zhq5v27Th4+WT
Ryhz/9kPOwCl89ByruSc93fjoMDWWxJDT4DXRH4l1jT2+mQWxlE0CeNtBsjmsZR0
XZr65Xh3tETiIAVeAzKNgC20Un5/HB/J03OVgS5f1pj28S8RDj04VHxQHcb0GYG6
0zwR0UgSy1kCg6sEJmd2vY7urYUvVxrMy8pRh9BjRx6THG7xnSF5nF5lohHFoYvM
foy7xmhi5zZYXE3Z7LS5dxXwxV5uXcm3wmv39Ti5MWV1CpE+EHvhUm4+q1JHnsvy
qCktUKjBiOgffCw0iLX0s5Svdsz+JSyh6hyspfJbm6o1+J75dxf2QVwTJ9Mpa1BQ
Mky/M7Zsa0hKiIc/buNJdXybV3CoEa33LLqfvjf3Klmw0zT9WmxLzYIs0mFhKVA8
f1RmPKY15kSDtEE/hjqU4gElUPwzBvsyOpUjWVLmw6iogPCxUT4rZwnMH+6nULE9
5NoPiA0WtDcHlhHVTvVsEqn2IHKRAmFcLQLOlMsCRVghj929vdPhfW1RRsFlRACo
FIl7vtzJPzP5o57xVIut4nugFUBdxSLnno0+OgIwlsYdTBb2kjwATWsOO2WA8flb
VbjP6Qt1LmrMkXR6OaO8A4cGDVyBS0G/DUNM/qxD4M1Q4/UdMuIr66+byVAaCTB8
Or30YpZUAfKm6L8yytUlmyXycgTSXYn4+WgkV7RVGPnc/DAOC8hlCEtGwxKiptuq
mevZfpqXnUp03cOARYLURqFdFFf2YO0hNVgjTRESSIVLNbuda4uY66glx5BW+FGP
Gez7USNG22NZ62vgcky5KEtji0wtGFDPsc895ayNLKRSsCwjBGt7volb+7bsA01Y
Gciurycznv8Nr89Q52hmXO9pYbsnrKPBExkpUNfE/8sWV3XGAfNM1XtJTYlBccyH
`protect end_protected