`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1456 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
xl+hxsegM9+gPkvRB6CsqR4GKDBdcD+DDxlGEtaJAL1YA+pajBx4Ckz5al2xTQDF
+6QCGqu2c+nhKYTPwm8LYsCwdVLh0zzf2ZkTnrC2F67K6faFjXAwwZGvBdrHGQZ5
/N6UexVGe4Pn7iEO4ryPwXWpcZTnl0prdDRa5DIdOrPdwzeH/tt+yC/Jjg+Pp6hO
Ifqq6E6VmjuY8gztx22/yUyt+Ne1AWF8vzQ9epDmEc2rUHbIoa3U3uYSv9kwlQsl
jiHxD0FIs8CAyMoFbuIawfliLm7ewqgrEhl7hISQW9a0d8HML3IvrjqPnG2nmmMh
6eHOZEi776lHQ2/Xr3iilNyNTGn2MTtwvXTm+NOz/6+cOGEUDvzf3xzYx7BiE+Xy
MboaaIIriuM34gKnm9fh6MvM0x+GuwwYZpsM65xvAoX1+5KEqG3MPQ+S98s14beE
UtdpWtqVTSjHAHqvWWARQzq18y6jpDqLZwfuzYFvZCXTc3h688v074p7hHTapQK8
+MGUl0L4NvbDQfc+T3B05PgQ/wVrmt6nUEoVrwaaJ7w9AzWBVgGAk+JNt/mSYzUy
1fvzoOiZiUDB4i7AJZbE2cPVS1DbfWezIm2+JzQmk4LjyjkAxLpQaHZZVC77KfJW
oqOwdAbz75gPgMgi8bZeUdBx5Bzqj8Miu8Cx0EqO+ha7s1PRrG6dwaSCb0jdG/sx
UInZERF3lOwPoqc5FtxaGdvMNEOZ1hSOYfEuXel7vp6UYPUgFTp37zm/+9NC9OD9
bVEfnUXcUIGC+uc/Xt8YfBrnOg/l651xWhv8f547nIpayYRNiI5qBP30UaW4zGK8
Vq8BDsZU6c6cNQ0DKA5CJncSIg2R8dAyy/A+RKkgyhXL8jLrz9tpQ26v0QzjXIn8
Ep5tyrCZOfzuEP9iNe7mzDExmeVIg0sIr8p3L82sLm/KU9cwuaxz4dB3EKZpWJBD
PtBHx5UT6IwNwJ0EKUt823PaXQEqbb5bYdEqOZOJ2d1XKMnrR24rNFeeEKnsvzpg
rvcMfNF/Sl4MEcatoUsPujzD18MV74GB3rjrEclN6nVCzZoFS3vuiE1Zpj+etahF
K/+L9meBMicgpy2TEcsTtUgWLT/RV+cBUNbqb0rNVTEyX8G8fSaeYxXLv3+M96Sz
aJxOrdWXE3whzR24QwkeNnKT52eSCVSFVa/TNorpkxAoJ3zCdPWKp/gyCmayku18
uGTwGtXW6a/TT+kfeXTwz/Ehq5GD7xEl6nSzzNYQIRXFaVu9oZwanC5tVXocNUZA
CsMgDhtoCpI3kfaH969+vy0p0ZknuwNIIIFswOpPTL3NvFjKGAyxfVIwHtlle0qe
CBJyFX6RxzmT71JYZUZsWcifrh3pMOPAl25D8XKZndaKleu7bG1zjazFNUJbQG2F
MLrW8qxgd6FRC8n2II8csRg3Q0ncQ0n2IWiV+NWUTVSlFWm/ZzUBpigYK04dROnw
Z7GuMEFP3trB7aINxJeY5HTNDvxOGSsw9wCKn429ZLYquAFHtBhPCjZMNuEvNa2z
vvfL48tBMZ0A1KwjhWHbUmK+eC/rD1916azPiFStobS1SByFkYL01HeBcZEc+0Iq
vJS0PCu4hovOaY3Pd4vtFwjG2kNNLEdtu2GXdliaPvuTyAxfzo2spn6eLoQ/o/HB
zYj5kHe95oqKiw1Cj6HCSoL/uRkcr7KaSqQWjuTW9WRx+OZR05xbeGn4SGevP6CD
lE2Lbs0y2VSV46vL4oxgyRCQ12cbUPpgUvVA3w6uiZvbLfzG65ePI6/QZZ2Vk66+
xaCktqOB7zIneaKg7RJ4Dw==
`protect end_protected