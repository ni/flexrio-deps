`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
X02cm7RKp1b59UGd/Qw0lernDa63uZp8Of9QINZf7jA1WbeD+7Av52J3NlUvj/+q
RyoE7C0PbGZzx+iX9P/4iglAeGoJkrjurSM7gzJAFrztSIznJ8A7IVrMFeiquijJ
JF/J07y+vzkpvO6rXVfAuTaqE6CDLgDXlsTP5+CaGqNMpWqR8f2Izt4BPNr7vEGs
8Z0dWixiagBc2+RHCJ6gSQhdN/I/bImYOD5/QFOv6hJFh6+Nq0WTvGf7ahelwFt0
RAKjS5m2jb7i3GqPJAM2ltJsEXGMqlWLF5CELuwji7lxxpi7HEt7U7YF0CKgHEw5
kF/8xsrElaiBWKXpY9L4h0usz+Le6Pykj8YdekGz2n29iASq2CtNvxKAAsC5xV98
jM5dhfT1SX2O0ej/ELsitHkllWfmo8VnpzTgg9EfZJzfTsp5aosneJgZ3yXVP8r/
2RFUAuglltyGqvESUU/vGEQwzjkhF7tpboymt7i8sRJWESdspyoVLkD8kg2vJFLx
XuFUTIfWlFgWL+d0Lex3dCKx7sa+2QngrVtSJTw3V17ArwFA/0FTOEZzNxvhwuOw
DlPMeWFzPeNn1jm5tHN5SCJzXLbLDf43epKfV6rQ82w702/xztkUM+4AdQ3ydLXT
s8MuSqyOlofUpbzQaoLXvjfQdetX4+Q0Qnd6mf+bHFUUvw0UaUXWXHDdpLt5rtLK
QF8ek3ktQpmlEgqWGQqClU1fD5rm/hzpFcq+Vv2n6nCy9tr1qR6bn+TBizu1r9kc
tshRIItSvAF2qnqrp2Am/UzLT+1zWh9wN0w7Jjj0GdebkoV6g8cNde9QydCGWt2K
yGeM7t4X31US7oKkdQfXpTglTqbpikAvTGqxk4xsZpAK1/1oAsxmy+4quEJSukE6
myH5Bfy+rdTbYn3LY2zcUdLMfLE1e1pr+rPtFNWZTEfYi4VIDTf29oM8AE6b8wnO
poayD1gsEbUs96GtBkqPiiqzSM/fOMbkTaOPR+NIlgicH4atw/+oz4K1bGhkoUCY
zFVgvUnTENAfG45KQreoRJQqg3fLLMayc2kE/zFLMatqDoCVdiSWwgI2mXEF5M9z
X9vcgCXSSllTfy58J7dbMJO/pHRaOqGo2PrKDXKDqZ/2p/Par6mMV5yqziBKx9s4
N5T512zQJwTY2TP9L5TYjMWqJTAp9oc+m3zcTcEPjMYJaru885ZmPzOWEykdRVPy
az5hFBreWqolhCKdMEts1CYg+6godGG0Pe3LIIhNm+bcbh/8pbx0to0AzUNvdsFO
lpkiwU6HU9uIKRCmN2oYVIIYB12CkuqtnkDdS6WcYiBMzoWg25rg2ZmiwNao3Oc1
Kwn3l0I3/G8mc4mhG5OAh89UIqAWDMKl9m4hM69oK/YILmeJ+MZ8E1kvY3CPpSpi
78tMETdBmYeK0TczFbW5tQQMtMu+0yCqVAdj9OCCE0Oxdq1XBu+/QxizOgjfCYYO
mfG7APF+/9aVH0JFsnCO1F9ePvIkknljIbj7qgeNpAcLzMybwdMtn7eN1OHYYW9j
KxRDm9Fd/RUpi0VxIJGqce4YY9utaSnjVRoag9HVqR4qtZdkA0ft3SubC1oGSQ3w
eaTVGPfQgjXMSoKKEFhnUfulPxPwDGTIuUMGnlTrG1sU5UXufM6H27wJn4v0rVbZ
r9D+UrA+z0sQSDcelE2UcCazApDIzXIZTpkxMKvFzG5BNOMbP33JS5w8fk8LfyYJ
XfDuK1JWc21plkZb5vARm82bRax+qljAXhnEL/oKGJST9ANeuBO0dtpG+OLRkjr/
74PW1whHLBiAZSJqlL+WZq/RYWii1r9bwj02MOMelk9qR+F+aw3bdPeddu8wQo//
e6HWWZpOfAD24I63EprMi33hiY78XOAFRiKqDOUYXWJR0OkpU+A235yXEHzZxhgo
s9NN6aBcAoGTRiefmzuv2M2dQtxq1vU12MfsXMEmCAuoG0+HzQ4oCmDTsiAl1E2Q
mJKTy7yYmfO41wsAUTnqyz6yY90nQFRXwooGh1wv6f3FixYXIq5BFh+OGEFrLKR/
gZ62K2/AJS6nAAkoVOCoeaNH5z/w2Caonccuu+f/ObwLw7x2G3xp9KErnAa13Dug
vD81JeRh9ujnvV/9XEIPSuoOJYbPONm5YVCVEtM6mzg=
`protect end_protected