`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 55056 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
TDkIdcJUWDKCGvmrQYRemB8U4kX1hPgGoIYMRPYAqcP7S/DyFflj4Ibz11rHftAF
p1drFkj8kymR/BW3shbQAiO9rAuQam2NjzS+rl50Dh5lpeFPkiaxRa3M/Gt7dC8b
MTKsgsESACi3GyrNzKfs0yNCs0gDwlna3Pq9kpp/3Md8085cKz9QeJKcmy1rArpd
kHVMy7yms6UhcSMc0zJUyWnVoKv69JQm5NTTXW80O9Qg+iMhxemrexoUNs9UTjo/
mX8RpAptfGDekYKNVtJd7YqpB4++6eOnFeqc+Dunh/+Jwk3WfF/N4u4avfSkwnv1
7sKncGQytRPoXLYivh+JBxbsPDpI8G5Z4Ekan6f4GBEHl+R+Gz9erz3jIeUDc1V4
dTonGXg9scc1KOblb/fTpgL+fm/TAxL/Pv3XazR1W5MLEsajxtaINNHMuty5wVUP
K1yppUn0sUFj6X1l36hy2wZVCOW0EiNf94PIiasylSMyTQdLcjRHWuki5wYvMl8J
LUA+c/BLyKoKgpFEj3QjwdfXZ7+mOFqvxTnweQ7tgrtMhU0ArIopsJ4eennEhFcL
0tcYlY41smfIbVn54O25WIjiupctx9ndI93b6LEw8+cGU05E7Cqsbro6wHUuWXY5
G3r1/a1ase96Vp1rTeaOKpQwuWqJ4NUdybQv/acRmsEUVq70StlgFGYRXe1kcBAy
Evuze/hQyH70GG0Jfp91/Mi/9iuLl6mjOUCp2Eh3ihPKnyzaZAw40BpBPF2XDZBw
UBeviq/PVOgzoytyUzu4PHkc75pEQ0HRKJoyBimVhb/QUBFXRWx713CHBSR0ug6V
h3Tsw9ZUQ9Nvqkq6P0dVFc4c5JTp9b5U8c6dvjYAaTo4CfHq0EgV7oMI5mEC60CM
gAYbUxRSg0tg7nc82IamHBh6M9WZFB1LdY0Yue0VK010N53bFwdsxoPcM/HUv+b1
O7QMnFl45Kzg0yV/2WCkBAEP2jb20Pq4AP6emFfxsaoajsMTkchF62xn5jHezx+Z
4Q8104MIm72584C6y/w2qyyROvq1ZxDrXfAxkSMW9OG4yvvxLsW9Xq93hP0/5TeD
7loHNNUkvKhTTTebjDW5cTS37zEED5yZvP4O4t58Apw/HKcgSdBXjQgIiFrg1WcY
fNx5PLEBuTjjaj4aMgLiqxyxNzuAT0mZeUaxeNkbnyziwclRKQCb/s3lCEFvbiLR
jkV3wNOUasaHBOg/jhokfVIf3SqECbIdR2tUmp+MGesjULzn5yI/e3clz9wX5ECs
x7iUC+zBgRkoWtIMMiMflsKw2vrijGGMa6TRGYXjbJYXfeA7QZsbpzKEwPdN4YcE
sWgQY0Br6+0zv+Gm+iqlUZt8rj/1qUEHbFADGKvouAYwCKoaOplhos7/sZPLCoOB
8vYCplqe3CDSW6Romiezlo6XWUqCiLvxAJK3i3NvHUth7zpDBIaqAp70Lggurak1
QD8rDEOw/NpfuwUIl1JCApksoUf/f32w5+rjuUwNTRnuCzWlv9uwKTTt44uJxit6
FWyKtcsZ9G+Tc7mcNUq5ejtkJePa6M1eWKdEigb9XzymqxDdSML3ehvfbU9944Ce
4bihmam5K152U8P7q9Nwv291Elq9pAZQIWft0cZgmFu8J7MsmA3D4h6o0rj6ULFi
hZu/+BUs0r3ACoBsx+mIkkoUc6qOLnABIARNAiVmmusHLt1JyO2sY32vrK/NOrqM
XlAO9N1hI0WvYEaQ/B1NNx/ONGsbAb83mMzjNHoIv0kfsoLMU7MmYOuVRmRKDbhA
GxD/SAAYZMjG1qQXPKkghneadkcXzNN4yomnw71YLSHmGAYPvO6JK/y/K/NNG008
lh/9zRnqJgHLsliC+wO91jH/27hejVfmOWPWYRx557pgAVafOSFHnPwnd1fzvYFQ
v67rIp7YqXUUevOHwoF0EJZwOr0yQHs3pH09u/JTRxIjTkd6qQ5UPDLap0mBwf5L
e6KTgsK/qlUnwPuKTt+PuFIa1FDNCknUG5AaUCv7Tz8mUqyrc1YaZ0Ha5IHrdR5h
C/tAGrkQs20ZmTtsLt8CL7PqjOmzeDOLHsfZb8Lhq5do5hZKu7V7bLYtnRuDj9D9
HwO0SkwCsm8LKAPDdPu5Ot6Q+yE1x0B2hphz89bCLwR2fqT4PvjAcbWqqgNQU0sT
mGzOs2To3LjRRZIeF7fbkxmCEZYZ35/50ZpOv9fJe1idBTv8GbSMvySADKeD4pz7
Yufm0ME1q+LAiCeUpMk8uQrYqsxr1TVa0CwrVzQKHqm0Jz4wbsLu7+4hR5FN51Ec
hSSIcD2Wn2YirqmtdmbkvEFD/sQZa5JQIFppQmXBNjzNAXTkaNX7bNy1Xs2oISKC
GZIpk1o8aM8u2dP1IhkrMzsemxCcp7EzMP3NH7NKQ0iOwf11q1Ne7feCcLaQCnMa
x+lFvxN5YRuR/hyoiYhtxGaxstpf4JghOwTscun9cffYO6OH3Gc0y7M4bSMxJwZu
sM9CXF/FXo+vj7sXRMmh00pU4IDQW8OYRBUSKJSFRIgh2z+o87DGrcOcKsB3GFWR
3KxTVdCN7TZykTFi9Dl4ujdJYPjyRZ9r1ykDnrjsilJ0QCeO0vQpa1EMkIA5Y8sR
Q5TqCGoInOcnX/0fV6oZo8AX2bF1xm1bAuN2lCi9teDQIiyoPjRkJvRexupbedSz
QICzd0K/ftYh/GWu8po7IiMeEzLoRBeW4PXzzSJA0JsyTe3lq+cmWFv3KpQrfz4j
I29U9qnCste84gHIdsMxHkRtr5jW0IhMS2S71kKeIJ4hm1c6h6p+Pw6VdPU5xnga
nor1YjuWDyoir8cOHZRIGzpISmNOIOtC3H9/C2RHgUMwm8lZ3aSZms4jY0tR3g07
ZdqfFXDSWV5YlrNO8A3T2n+mdnxAaQsPePz1gIEqpak9c0KYCJetE2PP3wfkLN9f
9G/rIEAIVIeqpHZD12fOMzSmZJWZmBJM9skyyR6zaVXW6xa59X4BPmwcqjSK52ip
BszvAbVcIDuYLXcpiyOk3n+fLFeHNtDJC19jvJDw/SseQBEUs/cdomvup95IAlWR
nZcBIaF2HfgcGRlHqUVVlOmVKF//vnV01L+/Imp+o4d/TpUsDC2sGoN4kTLA9YSt
sC2GbQz8MEhN343cIbUnDD8Dw8niaHIofdRlqaPapFyhlnYECyK/mqkXyrXzibiI
m2nYPOFX49dHHBH2ksUWXofQuSvi7YF1s7DxSiWGdkpdInL9nc4IocD+nTukE2Iq
aguKEQRHCKAIVd0VpZrgdPZYJ974dF0uI8Q+Vj0pVY+LA+KcI4/iUTh02Q3szHvw
OSXLdx/pooeNdlJ4M5vcMeTTRpNnEvByLUSfiZckv46jqFZCOCrB2l5uRNwuT3c0
ST/Dl0251bzzf+2FDRU4NUgv6YHu4CeCEuL+SaqI46R2Rv7aytzoSjLAlVldHB9N
Er2R/36SB20HxsLDA7aaH6d7c0rAZ0P0HrcpTmfvpAzlBkX8ri3aFgH4d8BJqsSG
Ndv/aGR0C5ECM8HXgJ+Grxp8WcI58AOCEhsMlghsiffjLwBChpnkdZbDAXbZqsIs
8sefEmhdsh4ZowNxtc18sY7RVbhdD9do46pu6Hrt9sdYxqFs8bsbv9uwhMZnoSrH
lcgEmi1DF+9wXcVEoFyPKMBdXlRVcG+eY3mzQdcqZc7qCLJPT6Of+BaHcEH3xIOX
Qb4bS0TbKqQij16K4+2fJLCPteU2/tR7KiqMAvctyTTIY5GwC9qA8nE3RW8DvT+d
o78M4c1yGevE7zIsbqzNqIsfWFwbIymM9IUfaXC7mZgl7JbaszgwVG0BkPbIOSRX
F+duvnM0cbox/ah/CHiYMCQ6V3VFiBmaceHPPurKeoQCjmPofQA44hGSnveLQSuR
pVdf2bmVcMvDPj9bzBSgr5zSujxlmBTtUWidTMw3yKzzE1euRUzESCntjrzx4jG4
eAZoZbJ7CukhDeshQkwj/d30ML5s8qy9soACY4bwqr1oFYYe/yLCShX7mfbI7CXT
ScFVviRILWJcFIszrAROIlYdJyjceVSeumIkwy2P3DrYf02yO2neisBbmhghvCjX
9tdNt9m+pWR6zhNU1bILKhbfdsM+anWujk75l2As/UVTUeayFlBchBKT1uyxguJp
YgMpV46wy4LtDvRaAIWxi4zIRoYON29Zmfj4INmkiIuAfkZpIKTXfBUZHucVTAN2
ansHgzrll5M0nefwupagV24Kdl5/scFtYR22ReiNsqCZJd2MK3CuL8JzBitIQUBY
sh0pmIO59GUSFRPJalkaV3uVY1BYWCfKdGDPIg8dBQCk2g6rN25DY6RY5MGUm/iv
oJqy2q0KkOkScOx794Wiq/O7sWYnG9uowgBqKyaoAA4x/6LB5ncGv2J+hsPLhhH5
lVeohO7pNLOP870NqRF5/idApbMpkxoXcczBzH46Il6tW7JHAM4R6H1CSUk8zPsj
VgewRKdnhLqmqTnMlkNSs1Beca7wEPqPCxxv2Xx1tQ8/ygDjC1wt/SKlCXH4+eLc
cAbP4dscmO1oZUEW+z2IXE2yThT/yiHJE+MH4/g/lUb9D4aNFc34L0X+fcJv3YJt
Ts6iMcokiTtt1NrAfDgWFqBnQ4HBwFt3sLo6W/WsfjfNu2xZj4Z39DzKjeRduDF7
owqiP28xMMxsBeYFSpAL7pASAIW/eY2nJiQ5XqB+JnpM4GOfkiF5fuNcBAeOJeaW
57NDvXo/pLuKk8WKSFLi2Odyajrz3RV26YPq816zTZPV1qa7oixNtHmzuJ7tBWMI
CTbb1TMjZW+6+9H1RSn/qo37veMlOcZjMCialys2xhnYH8PsG3GOqD31mTkhQR1d
XZ2b7oiA2FAl0MSfm5+hUA1asAFQo4dGABeT20W+hClcwWwCsfwE3PCkwuJKSWte
PaLL+3U3o3OMqC+rPGfFQnI2mDSbDwznYJ+7ldRpWiz6seXs3r0pxnm1AKiy76MV
eofNxPC1tbBBiPPLJMNVnS0+kidlQdXpVwlids6assAbspzuWqp0xdhc5QMEWiiH
WTJu+UpfbhPsLDPet7gSTPvduwFCjJiMihzR0Sl7RrEExTmhWdg1ft7OE8DWlLBq
/q6U2GuZSC9uS7kKQ3jhF3UnIVSN4ZyCofqnWKPELqMdQuX+pO2ly1duTWBbJN/U
EQT3p+mCa9BYMeCeO/YEiMeos/IF4516nP+324UrGY+cf1DvJ+UVAge5nRLUuUdo
EseSgXfB6J5bZZRQR8kxaELs+StDQANTHZvjYLvhCnyV3cyl/Mm0eEX0vzqNKWs2
SEA3noEcoWieKTjto64z7eAbTZrW3I0z+f+LZg1mTT1iWqNKVwFCagRT+oVIQC7a
mAP2LDmYZ2ak3kOoW0ah4a5Czeeh5tSTImMnbxF6oa6kGFa+fkyCmrUW2a3WzMjA
A44C+11qkLLQLVv2rQgkf4kG9sp4rslS7o+lF1oSL4tpjTOmCRTlyP+LEB1zZ7QY
ObdSIsfCU8AbmiDLcBkhL4ZkaqNMHwC31Gu4l4qr1TLm7CABredJ1Bx999tnDwjJ
DG3IRcC7aqMbS0zKcGsALD+hReeP3/oicSOJgMgpn/uO9fLDT8an0k+BNndm+ePg
FM2VjsRmRx8kaQUaFCq3bdJA7+TrVaMuqokhFcQX/sbiwWsyn8MSBMsNb6dGllQa
ZF3cu/jRKixhILF8pAYdWn/YsdcmRCpEyzyJsNl8D3LCnGQSSh54Aid+HqLsicf2
yffkKXnP6hETV1mngBcU+ixs4cyGKTQN6uIi6QNXBg3vS8aQODHQoH20f54jSxF7
oWRtpJ4fBn6hj5KHf7F632o+ckkpEYi+1cfzlutERAIg7Nt/L1KPbX5OAvctc6Id
GspUqesaHuUVSPiRE4OmVFbaxZvgGRjz6PF/cuYB4rENeICz9zjKssUW6IeXwYZN
mv2nlJsOKN7VVhMuKeAufSfM8n3xpjo1DUo4Qbk8hL0MI8hLBwEwarEmckoZoSQA
BozNSgKBu5eh+Wyo/HrlIYOq5sVAkZhKURLFa0TKvJSqgB+4wUDatgRNCYdbpOkC
tKsw9Y546mRdhFk2I99JiqSfC+iKR3dV1cumOq6p1e1gfDY3kOR7BlDBWkRH5xBL
C0QnZtndDzgDUH+5Mwrng2QZHSjE9esaVIEGqJfxDrBCbDf93Zi7Y1XGzxEhYJ7l
9iNbWDDpCdbVcUvehXsQaNrnVxJ7K8pcuFsO32CCCFEnY6ZtJeQvJmJvZu+LWk6C
doWEDab1Ak8iFK/HjJo0ya/Jxk9ca8KNzBxQJhL/n13UFsTTyzUEXMeKCCY1htAw
QZOkPf49tieGwTbd77UTze08X/CTeXVDjH9Zm2lNIQ80ZZPsUjwkg+mbkr8SIHzi
JTk4MhwNWzPDyNz58LNG/leriisaNSwG8HeHbjrBpDHgG1ONq0U+C8D4mndBqF1M
G2Z66lqTrPD20KmDiK2Chkw7hhvdWW6lIA00UJRUKaPrVURMjFV5T0EZtcZb+qY3
cYq/PYJHzXKqRLpuaa0G5ywMuFQMlTfIJs5C2KbowtIpWJq/QBKMMglnyrqqms0O
nzO3JfUtQbFJMjR238xQzYvIWpK3xdf5Cy/5kiJDCu9ZCZZAnlY/QY94cKnxSnFf
Alw3IuhRq0vLwN8sRm9z8EjYcuZBYM3MB+xpR00rPW85F8zoLWamlutirOHIO7M5
9Rm/lXkQKoHYPMVLyk1cr/XK0Rt5ykRatdyCDMGb3RWaqkCeOCFlCHR825pCeL5K
63GU0omHctBn+yteQMyvCVz/E7ANnCIVD7dajB7nClxwrx3VG1hN9feGfYNy7NRi
JfzR/a1bgITxVCNsH+Y/efQz9spBNUiau3/NRqfz/Jh/r8UtpYzV7fmHdnVYDxuk
YcJ+7hKB9wGeq7MVkmir6r6iyLuCne+lFaanGyiwIq5C1kBPgp/jOyJSrDfOPf2v
zqMDnn5g/BmlWfDY2rWedxStdVc0yUakwcmpqZoPfYl5953oPWyZiz6pz+1qovXF
L2tUpoNAxKh/GMQaUHyCSbcK6Ch+oxD8bzrJV+owrvepIOXaZocwpckinaMZSv4w
N9CuOKEO68J2afr8xY3ykMSb4FGVYglCKhvaZkxs9E28gOv5OnJstPHAbKGEmRia
/DNKTrC6H/tYXPVQ2QBG1EFjgW0XTpsnl9qyd5Q1fz4TLPc0j8Bidf6L2CZ5uYcY
XU2q/Jmp+Q4jwzv1kTC/oFIqO9Guz32i0jC/bg1S/Xo+w+BedtZYqI29KaiHKSuX
rlo4ar8FD44mrbPbAeVgagH224xl7JQPnbe8CQUVy7lre3ls5Legx9MMc7+nuBVq
zI1594NhRyFkLTXW8lUGb7kV2fXrVxkdWKzqfiZ3m0DJOkrM/Z+otL7IGiFsCebS
3ikEw9JPnZp4eH0lkfuDZImCGNhYKlhO0vOYFsMUfnPuzPnIWm06w1O8qANQAvjL
6bxex7wKq8mOhSTl8ktt9LJuwQw2KiAYIiBPJ5wjrfeqhvSdy3VXvlqY44RxRd3T
aUG83zxxhCnrHaf3qqEHO+9EoRmNk9QLsqYS7Tf2R0QttYbcAFGA+/l7rfmP9S9l
X3/4OBRIppLABP5E+kQ+ZVcd4YTn32WP4rcYAKYlSWtvbCZUd8+w9vIt2wdMZnfn
uZ9HdigtSp0oMTC4Mx1reEPiranVl+6EOFHEkMy0TkTgnDBDceVTFV5dfsv7+4bO
IFVrbChXHtmERWo625LZPFGdyjs8sETALQBlRNVR+tFFazIWpO1dgfjG64ubgL4k
eMIEvXjJrNscza6RgX2CHYv5GoJfOr2iJmOmlzfPd6WSjXPN3Yuel2bSi0Vw2vqt
k3XxytNMpg+SB+XN47Z5/t/Jpj1J4N7YztPtBtAwAg9l94msdSKPV69wa5IbE/tH
dx/LE9LcMWj9U0xTmQ7RUGruiF2l3ObFt3O2kEmQnhFFfR9IM8xE/ZK+Jwb9xmL/
aaqJQRvEZP0fJSA/nLDSlaJXqqK+AV5jOIvtBfFHwUVflD0UPKcDLOFTVdlCOSm6
2AJma5lrvKXteG7wv6ew9eYHSbXH9ITDmLdnPgYfIAQ+5X5+97B3bdQgF7p0fU58
H+ews7QW/59EnHvmb5hBKmlEJy01oMyh24nSsv/hXiahjJSJSZzTuzAUYUxX7C1w
xrjNFplFxDgaF9w858q4ggsB7d/MI7bAxQxwr/gd3xUD0FAEaTKwSh44hOAui9EM
K/5s0Ls6L/4VqzgcqmzL00eCIHX1Klz6qB6ciKJercPpn9RaDBpFErmZXmurD1Jo
eY9X7C7IKYmc+d+hFKrr2UCliNggaAna3g3oz7F64tZ3JPdi3uKMTsJOvMiRlQZO
qt+vpCEwcGk423WqL1nAJe7ARLnqj2LyOhGb9Dl6rjfUVsnlonk5A0vLsrcLfPUN
m9bdO1T8eNVX9OWF84WYjRRku1XlOeQwzxckGkEdlKGleiZXlfSam4pc4EJIVum3
Pckrx9NMAN0yBVSZt+idi+m7O+xZTO6eV4Fims0pFK9ic0aV6qT+JbAbLUQcIeuT
GeLsxafUzmHFww6C8crxHnRgfiOYIvLrlPWKHifqle/I4a+x+6/EDt2d5OERODD2
QjmNXlcSjRx9avE8OiVIvI/HTTbnggEdc+mESyXgCkKSDWgA8n3eAUFI3VNp+3/9
1FV1FbkCUiUGtP7Y9F6TM6idOr/q9RPTpUybMgDqfMAaKSsX4b/cIr2S4pfF8M2q
VvISuRBIZGmJmIvohvUwR9L58uBzyKOXomUG4pFRTLrXwetSNfEvhrdkBVaqmpMN
0kwW5QngrZ8seGIrArbIZtGLJAwlmFhf2LTIpte0vARVNH5TULX6sx+phcnEMHU7
AQyfza1dj9MU3G86ZvCDVUDuoNF0OLtmO7CM7BlEK/akAPuyOv4eMqP41ER6G9dw
nVkRRHwI3mWPjM1WNyrAkx+EWQ3IjCdTHy7dFSHFQowIKcdnRWC2+aw8LLVq7w7n
zzKp31IoX1semM8jvxfgT2PJ1BGoT2alBx9a4eJPr6ut2lVUsd51JDB+E8i5YPUH
Q2UEflppkSJKxFD0PBrcs7P93ef+jW21DBY/xdJ/HPXWc95+wzJTDghZRyOdhvfs
lDS3PDv7z6agFfc2KhD2m9G58AFgV3pknyR8p3yL7vKBb6jVQiwfLcfZlhOvxjoW
z8hhqlocckY28Up6A/sMYjERCVOtLkP+bOhUobRp7PeUCmGnNvnfHhRVWuYlzS+m
J93MCrjbAtVPy5vvXcXuqWqqFeJLkTde/m4xf5bjL2lSnm6MIsoZJWSwsYN/H67H
Zlf/xFzEXmc7/XLF2FSGb+mmG0l+zl0wtmdlz7PhAkU3QaA50AiV0oYpUU+Y7/kc
GOTQ/1ukpT5ESECkVC7pchD/XnTcX1MuaUtWDlTdBYU8Zi7kiku2I97f7c59MfT5
j1cQKfJnWleJsDTFYVp1RCu8Oa6Y8vfkNTjE35aZdcg5jJ6jxyf0+Ph5IF3fPlZG
HxU8Rv92WodktV8Qlw4pvgslKx9KxwqfJoq0b248uo7vmz7Cw9SlB78JO+mpG5cQ
dQHrbhJ6VABw0068YCRDA04s7S9ahFra84TlF/+RUwSLy2zVxXrfdPGPFaKEhqGo
6yMK7WQGrqcHGinPSUYcToKmaC7QhgK+6TL1mgqF7Pt9j+J82Tk6VoEmBzL1WhcF
EQcXt/VjrhCNynOPLi/c69JTtHRt+PIkcVHstokHCOEhcmBbL2GPu6EX4PFQQF4d
RhGZLZQ3lIWd9UIdubz8KbfZWzrEp985wAXILusvw5JujKHZWHlkX5cddq3yPHh7
Sb4uyDYiIPn9fIEEmL3mouZ2NTgKLT9M7G9AcmENyoJPaFXIb30sEA9kM/qizDa6
HLWnt1Lnn3dL5IuwPcuSPTBiSbsJADMRuvqlFq/Bea50pgDHfXGYKaC7sruwiJoq
nPZZt5Sw40UiFWzC8zB3sNcHR5B1/phFNPKf0Yql+XNJ90nXQsSg6FnpNjJAMKy6
Gzoy0DoLxFGPyaoUudfnwtHQ6TCf1A+5EcsDm1HuY/osi7PCV1Zep0k7cJiuuObi
fl4k+cNzJw+lY0HMIiFiTDTeRxyk8uy+sz+qnTEDsJMmE1tKU6oy9ychzi7OXzZl
LKT24CooQfUbqDydyDVkU52Xv4TAmrUvu/MMUiALuslQMzH3iYCPw8HQ+v18H6wr
3w7nMBIVWoPOze07ieYqf1fkUtAQ8gkkVcLuw0yqRSn6msQwfRDSEAyiO4SCVYVG
DeDmpbSMcCyLQyGGW7g3/xU6j34ohA6Y0eAYIyArUCSWVLhaimIHDgsGfWJfTMYE
hKeK+jw5TzQeEEOL9GOrhja1XHCEIR9QrrQMIAToqnSDdzpk5H6qAdo0WY2NtxuX
9XsTUZZKd9ZdWqUAXCIdtK9i8KW9cfqeLVS6IARfsUjP3lUuo81mW1df+ed86ea4
gf4Ic2Pgraiw7crfu0xgFqqCroJm/Y0v5Dr+reGydOkFv+RVulQ6HWzS1eQr3p9L
tNgYpLj5ZNs/Ptt8WaXi0ZtFLben2mlUJhTCvmhDO2Sgg7V8pUwLP92KOxgciVmk
6kF8yYwtrPHbK5RqQNL3GWqUfZqivbfM/Pq7tNK8roGRxUznK1X02erwfVS8s7E9
qEvOhVmhna2k1NZSXlE2tBYeUKd1WGtYSApbqxwi9aLeyGOwV9u8c7syPhapOGRL
4WUsIKnhwvd7MlGfDZ8GkP09Vhl3GD449S3ETHLMI648oQQ6mG3gAcnpFU15QKVs
OokjDFRGN+9qaXEGQrL0ZVrrxLQ/N7/wtm2FRi89RyPSbGuDDqy6ESUhdDT8WQ3z
Z8u5GQpvYiftuRHda0s37wubWLOMGzN7q6h++bGoye4xpp+C2X3jnNNOpsOz8PLK
7c7/zdhflrsNctV8u4nlNhKYieB+T2l70LGjIbxYpDB041/knx2B8TDuIc1UoaQ5
Q3r9RRpgwWVoPGlUqgfwkkKWexD5yLUK4goIG28VNfnU8qwPDjQg0M+8axHqb74X
F9+WyCys80BXWgBF3I+usAXDdk2ZA1nt6jiaTHYT50fCg2p2A/Iv8glQ2XxUKNSm
nOXCgvzO6/Vni/rZRZq1GRb2a5HI/9rV+ZB383eBjyRRHidMGwR+ZA/u+GheTRZ9
ArMNEbY/dOAn5gCabcP9wc0SZAETLdmjZzReT0DC5gp/1vdcLHfrqZqsE8zqzmvw
KYnbGQY+Ahb1ldoMlx463vxcmfchdbTNUK/Ysngwmx2pmJUgjYoM5SSTZlOJL5nH
U4DN7rVs2UmvBlSVUoNNblYbpm7z3jiZuXKx9jMaTICU2TVkpalFDoBWsY0H/OGT
n8huDpM2GhC/H1IfiIMwmBKnFPXi9GowMUTxZcEgz9kuRkbJiW9RViCuoc+gcS/u
yOWc9HZGdqzQ3cwYnAcnoHWMmON00HJ1+SQ8BdEqZNYrjBpQcoL8cFqmuSdDSb6k
cna2EYcTEcAQQAPaUmi8l78jkbVg3AJlCZhlkeWP85mIhNFT66CqcRuJWV6rxSif
RZmtFjczIp4KVs+q43fvo/77ksI+n80ZKiw7FWb45LlBFFiXdCBGlzsbcSRaDka8
Uo7JfJZ6OlKvgkYTWhmuGHWIKb4vVLj9sSpP6IxuBB+7X8qNtv8MkTSqmBMJL9ks
8cG1WV98GgtDSQ3ev1b4dj09tEkHbCxjFF7RIWA2PDT850H1FO4XTF/v7hQOaHzB
UDmY6xpffDJQMGTAQz64Ret4Ut2+Et5wGsLMkiIDV5lWOYSOv6CEm2Zmu3U7EzW9
mCFioCpJc+3g5WPI1Z7LVSjzJhTmr2yhMY1qipBOc8Eql3/RF2hCc8LRQVsbPfZt
wr8/ArX6Me7xY9GjU52ypft5aOomFoT1yy9jvOWe8tIIuPho+HRjkS3ahi9Eowqg
66Y2u6Tr4jrpm3NLqKkrbQPUlJuiBIqUpsSp+Ai2oLUtpWRsTYd90KcHBUPG56Ug
VAM4c0CptgPuLFFXAR8DiqAuqjEvlV7+8aaaqJdGpFXtOXCOdHt4rg9T3nAjO8Ob
dol8TW16DpQn/y9O5TlW/PUwL8wGU0sKz/ru7q50FSc1ylhPV6nYh0uC6fUeWh/4
lw5BLnQ9fhkIQWrDjbMU68yOdSuN+iXIHo2CJeifCgIJ22FMRwlmFdIczHWyhmUj
ZpQ0+Yp0UEI19U36wz8kcSRCHCDneh1r22qbaXJh6mR7mt2vPyGb1f8jYZYs684t
MWmyESTZ+xyMs+IJtWaHBbwoSLn4xlEsZ4pVhRdO7efB2xG8xsU3j0Nld8QoY1LQ
sC2jP7dXs5zXPKYH82pFhpHCRyeetsiYJSB547I1vSftWkxDaNlwUBxD7K9xyTrc
QZumq8XfJ8j3SGkkxE6Rm2UHOPUEfGTMLP9w1iN33LWmgjD+4FAQzfREZU+W0RUg
9ExurMw4vhFOUkYgiltsmrbRQDkCP6/bGTLCqShyLUSp3kINGW3PFLtVrLRSMZZE
DA+NhL7lyEAQudVvKjR7ZLnvABRqe1R9AVqGbAqOXMkYKBaEV0HXzY4ZHlV9sQxO
rH9VxPH5MyqYjz/TWMXea05cE9GzbrCGxpa84lgI4Wdua8Y9AsEdIYraviDyThaI
1oQJ+DCXTP0eDNJhI1Ep/wRPpslHKealpl/tUX3hsf4SVVvzqhMd3BvzZkLeHptd
jP0IOPUmEcJsu7QV9wX8pRheAOVVLGxdFmeUNuSR1BKdsvtAjD2M81/Rcd0piqsT
/S8TIArbxcmBWnwZrFkqacwOxLwv1yGZkU43rTLDMdFMXqGQ0JX8RYozlXTQ6Lg4
X3bJ1fu4ST8poBC3u44VbYDp88bfDYUp/i6aMkNYW2mI2JbWdBLniJ3uKUC7EIdK
0qc7fql1VzA1NBEVnI5ho9zgn8y6+QJSY61lHo/ychCTWk1V0F1GwpdzbVurBFDh
GNzKlllzOI88HxIoP2GHjaZRsqFOxtAu+ulHTri5ULxxmCDF7o/NMtH1zIUtoo6+
Pc431TGWFANZnWHAjlrPVR4b2u4SWphEPnfYuFkOGmAS478BRPdwCFr/jQK4T/NY
seSBopFBMrjSrhuD/3T10mV6CYdNJktFXhzKSLYfpTIcnMRsrAIEDWhdB0hLlx4E
jVBuBI9cqB5kspTjaKgFo25585cJWXUwAN+uqq0vJZx5uyUuonqrOw4h4FzJBJar
ei1H3JqwYTh2eC3ncLaMZkXDeIqNEjJNbx3EYRBHrPfxnp/qI7xmRropq2UX5NCZ
CttubfF6uyIwk8peeGiSE3j1ZFLY2p5Lia78ea5H/6AFi+z+aThv18vwny7dUDXX
oNwcc6LNSaNKJReuX9GHjvLlGYIyerTTq2qZsxcqMI6ZIetyGnpDcfzv858WZwOP
fgBPcjAagSKOrMC7GwFAFR//Df3xAM/LbyhaWgikH0g4tULE2pMIzzmbruzgLywz
BXiuOi8zr5cVmPUWHYD4t13aSeM13blgQ0wLF5vZ3nEXMma1xP2G+owiO91ryCyQ
Qu00X5ZgVJLKZBigdT4OulpMxJIwEQNxKYuAnKoGzXD7uErVbP9xFJBBxW0SpUMF
d4M/YQ/qW367G0viF4y7nMzUK0Wcz71EpGsQLrVP1TRlpQfYvpUG9tZ2iOkdS9zY
36OEEJsZZypcGJxM0Yhpur+hMAJTxF0inRQIBFuX5b8pc86euRmb8ud8SJ1iSlsf
hEG+lgOC8F8VYbZMpIjMs6Nk+nhq0KSTo3m55kzt0bGuZ0OWgHVxFIcSbEO0RoFe
kJJGSLGq7mY0/XYAmOv5oxQ4GNBN8j3cZTdRuRPL4S6CwnZfi1U2wSux+ZMxeaoq
1es4CVpKIiTx46DhAxhZMGnTCEB3XVOw4Sc70NdAHk9aSlmSkTA0LKJE6MSnH6fH
YnbKyHIMBRts+QM4uENpsJHJ3z27QGKmvVyt5xTZa6Wecqrk3WS9gSMZQVhbSGOX
/2nniRjwUgF94jjr936BJ123YKWKWiSmoLo45MpN0naYlZ3l0HiA8QVo5SCJdg6z
vWuI5eWlUpsSH3nhsytXrdGEzXap8cncF7TOUtZXQT59YseV6wqumiT6b6yezw2U
OgmhPWbFUQ00c03rwjEFVUQr0EvAcj1WzLfZUcc6rPXB51nCSzs5W5tWRJfQVNeQ
N1jPGUylAXZeOrE1ARQnrbAj0svCNonn3vKKDwXmhkw9Xh4wBDS1Jf66J2pqDs0d
TEHFdsltXcxwKShZprLu80de29nqktN2lbaKx9v2Www/ebFo/RINXGf+NzBPbaiU
0e2tp2u4GVfhomMbfzAtzczXEP7nOQcp/4vI+7Zdnn97h52sMGKurHdNm6fKXQ1Y
43UPvVQcjfepND539xhtg9Pwgnumcw5ugh/FvQA6KtIg6kWYsas2vg6W8mjAR66k
eCsVxmpnGdzc/8DbvgzfnZSxEa3t2HPiYer2KipD6I9hEqRt4zaR6vBVJmw6d+X9
79QeVjCevYZFrkp9fBeteLwJ7wepjL4s59OQsPQ1iNyDlIuYUJHKx3ZO9oYtf+1c
Mvw6O8lZVinJJvq0Orub67bk048SoBghPmqSjdsVgDho5ATLWZgnA54Fqq75cj3U
sgspmbMFOrEncp71ovIsoE6lvbj+IHdPL0UH8O4DAzbVEz8PUG+jzIKBvF2ipWAP
nGOKa5c6u/CJOOHgOChm80VgoqcOtwqYafiDXkHSfTyyNoabt+vOUdNg0Elcl2VO
phqEHgfT/poHS7hRptE13n6j2qPBJJKFuDkKjtSflOT1kartIVb51iCCogBsAi27
ce6pHyOpGoQBjVjScyBeat8abOlyOoSqHiVf8Drgn61IN8s9WtiZ2abK5YECtDOc
nnInaLVBCeg3RtFMA48B5lV/zNXgmX+2brP5zmEhp5du1/e6qlEbSGsHqBGLKb6E
xIiFfyrB+5sLx1NB/JgQy3C31zB6VF97nXAAZTqWVLuq41pN3luIk5PHP9Bb1aUj
FH31vShOav2SnBV9sV8FI8xwISOV0/fakkZeu8jdCTdz/yT8ysNs2a8onG2LvM4x
fUzkiAsDdD065EBWjEr5nui+4fx8Edo19qRIKz+s1JfQWg6YWjlP9XObpNxYW85j
X5fOzt18z4UxyF1ixbaHYzMZA01vBfFAJTHGZkWeT/ergNFEb3u1ObB8iLlllT3u
n6eExtHqS1VLl46WmBN47mY8nCjDvOoCpLFYBsLgOFZZ1pkcAVZWIdXtyqQwNsog
1BTYPWfnqaCxHV0XAkhp7GZEmhxd4BUmc7+VK9Z24VOIbLiuqUHKbYYBcbyOa+9M
ll9FL880M1uEncQWrPmFUhx7DmTjJNWdCiyyHD9I8ORbgxs2/o5uukm5UvbzYB9k
Zc1iSH07DpZ7hmDK8aR8znWovbwBVRLXqFVD7YQj37PCSfQ5RAXThTGAO67BFrjV
PGkKO8ajDutrcfjJUosPn8WUAajNbjzcMzky41RwYzuvWrzKpQvswis4N7XH0fw1
O+j0yf/JDdoF1w+9uz4J2jdfRSPNRT1Oltutd4zQDuQ/ob6qs5zxKp6BrylfEPDi
2q5YD21Q/ALPwH6GlBfTQo7nQV8YOB7ZRwB253gvCmhFdLuZNAvTPiG7WvtBXhc7
fxjuxhhzWMiloUMcnTLDaT0deULTbJUC6XbYxJ9v5Q5hKx023jOTuFYSRRSyI9eO
vXFneZdYW/wlrFChw0QqeuwQdlerVgYM8z9mMDrQWYLm4j9rggBzHNlWb22BrPZA
VphhJ6pjRZtyiqnqLGTm4yYSDdFY6kEScZ403tVpRgQIqPsIdjX0CtgDFmXvMqOa
daII8IeSJCB2wroevWaj6asyrTFaaEXmdbIsVtpuedkzOKOeqA7A9LNQrk16pk9i
jtrL/gQ8p/LZkIXjw9QtUzYqYVGu2qIpg2623j0ovnVNL+61mQscZVsIMZH6honj
UNNnDzNUVDHzTpHGG2TfW0j/OX1PS8DscOZTUrqkPUpTrEIYJEW4PcCu/ksn7Eg9
601XWt1s0hPXjnypaIFtU8C7hAEWRa0CiEsyE0TLRReYY8WNBHk0qOkFFSvyIFZD
CxT46IhMRZ2I1vGmi1FXrrmuS4UMQ2+vukT2ObyoZQssoJLWFSy27v2Uog3g7mgM
3LnXdtzj08ASIhb+jvb1bZE9LOWvCOXNzMGBobtvm+7Ov6WjxyBLMhZ8N17lYGI6
scwJwx6/ceLbvo6OMFttunBgf4o3xMgOlweoXyn2JGZTT4qeZBjQjS9AbmdPo3fo
+huO7HXlA0RMqbm3lFyMKf99jUGBOnSEvxlF0WZiRtRzu79YxbEMnnnF9JMflFfp
hIqF1Sm/E01Qk2oBTMK/zxnOvBv6ZcwL6aQv/dITncAVaP4gN8zBAsCsA8hOTz8D
ClVO6SYM2HKk+mTXtzWrnrhcTkkSh4OZOtPvOPNa+h3wpr/uUtQi7xF9EUgMzc3Q
CpLOIIN/VH0fh5DSSsSrPFB3D6Sm/ReLmwYo/Al+7Xyet647wFLCr3fdhMlMMjPk
64h5vM/Gmheb+b0HYeIhmKufK2id9rW4DB2v/dzkgfXg+mvn9WAzl+88sEdH7gq5
04BRpMiyd/0qS7d03tUhdV3zhSDTwXRLsn+j9W8WEH3wEsUwg/Oq1CwOl20+sDRu
5+4/dMlw2vPJ3PszLgvy1FaIf1xJk/cwsHXPsQiAhczkW3xn4nU2qfEYSMRAnuIO
Qx8kvysfcSuEQkQHNrhkdiFr0Pq2m4ig2NJD8ofeupfmOLNZ91RoufcvBxSUXLQd
BMVbvIj0usz9CxFtU+ovaV8M5NXhuYtX726XU0WyQqU/10Nu2AmmN/5/Z5nnMdkP
4uz8zOHsHXBDAf90FRQzYM5V6vzqegbknwKgSup41hoL02faPCGtxjklmld5lFXv
EkYmkv4H3gQIQZSgZaH6wdcQuUYhxvA3+K5Pv87eArFSscrjNUTrdbgPhOB1Q7TC
9EcGscej5KfcUp3XvTGu5C/pQJ70Lgpt24oYZMfT9dm+DqCcFuRPjt/S8Mv0ej0k
VVWIGEvdf+XV7kTwiNxnKHgbXXwOHgBNGSiRE2qkPFYKBGgg9EGjHUtEWK9fomem
52bYk/iOR5CA3dsrLkb6Ni9HImk/7Rn60b37FjbRgCcKvk+JxN50SM1w0xwbBokP
yMuLw3J1leGTTRz5kg68dsbFusoQbHkKJBreVmOC5CNsUnlHwM7JqMpDaxof/Tws
3WI/laPyuN7YXMpdV2bH9THG5/A2XprtS1i7ul31TjZ835CUWs4wA3fq0ctAPwx3
4r8N/Vzy4IA4LPmxCYzmnzDX0nxFHf+/9q9PJiPSqVRNh057JPSsaCECX+mrqy7c
9ZZtzv2P3DL57JX87lcj+8+mVoUmU3V/2cAL0SCk6UdpwGO/Nkb43rizhCbHOfuK
7kpD4dtiQHuT8EQ3GtdZnrAdbms9e253yk6SR/Z/GyAu4ZF651rIiw27bu0gh83a
R+tt6+WBZwjIKhXJFwjOxg4uYvh1gBmoQihSvNJRHLMjSUVRTub9DGSv9wWYg0WF
tLeYX1lptYO4t2yFc71PGWqxz+rgKG5+zsSST+1D5xeIUadKs3u5M0CeAVAfygse
pcuFuv98RzI3SQ1BY2xvMdKyW/RDPnxc/wOcaaE2c+V49PAd7ZgWdw7Vek8V+gIR
cZ2/CDHccJ2Lah2kcjhvFBlt7DEdl8uIs4sRGETNvaOBRuhQi3NMqZu3RpJvZn+C
6bt24V8UuYkrPqXY0GWwCoGx86nzcA2Zxa6OflS/WDNDzS1E6EhIkcfAOOOnliVI
DIshltkqX40eafauR+IWZSmNHA3xrqjLobAVj0l8IKhB5pPrl2z5Y6qtKHGpSJbN
qOQObRmU15xgwvK7aujkGqm2foB4NPyD8flQt4ewzgDMgVWJftho1MrWMGlciZH1
l1/mX/FLKfIsNaJ9IMyesRUa/F2XhevB4mdx3Z54XnIw+4MgJmQ9fwVclb1lXnpl
k1MeIeDnQLMrRxPnZ9sNPnFcc1bEtxWpdo0oXGGzefEUXuuCgxfPKdHUfDbzFKah
b4J+CjVJdVgzAT3ORafS5ojqOHvPdwpC6vxDM1gvRW+sPdZOEqI4jDxVCBl7/o5t
cxiaYHDB1SIhAYctDdnVd1vbv56OYcMfWzPmRzekR7oxkCpo/M1FCIpGWnZd3Uop
H4YuCIYiyBNLAs2nelhc6wYAF+7hP3myTtICjcfZdo4CVly+9NTmh5jDSxxafvoI
95aSoh55hWcJjnJ+BnE2sG0eI2OdvmHoXVPsfLqhWbXWFrxkCJCBK06IyMHhra6a
M/Kw+P8ko2DwcTNWPwbsdz5SU0hwDZNB/sOH3LRPLPiiP86TfQ309HpMrn3SNDv0
3uM99YIVpxCQZwM6bfTDiQLmgkqLwS5BVYHeNTFZDGzvsYj8Dm4XJALzLisFptK2
J2hG4KUIMh38wP8zVaad10QnYMTuKjIRRC7T9qb8RWeIN2lQpbkQr/pCATkVoRoI
crNJ1VBKzzQxpoJHAq3sdSszgyhLVKcGWf8NMjmDNI0HlqtqeaCQco/+aj3k9/Ve
+dZBA7SHjFfs/CdhLcDIsEiCxYO3uv4zb7+JWHC0OzG9+N+p3Udaw0B+pOY4L2pe
C5X/0a03jSxiyPPD+DZlV+OOBnzhBBR3vvXmlo32fFHtVhzzrA4lsS/R6Q5lWHh0
3scE84oqHkQgKZCz7Qlqtlc501ttPLx9XR2mvHuVCiW1YcRJo0SRcOO5hhsXreVh
FxQ85LVwVhdtMY8ux6H7hJ7UeY48jFz1dbLvgGlssZOAdnwi7raPtn3DfmmZoEmY
pAQSqEb+OvBG1KnlrO87BdDsQ68a7AycML5A+UYtZMGNo8yuTepVwvNht9JlnGEn
0L2Vnsw+BUKAEHPvaTTZvC+g4OLfYVQ6QrDlaJsQ7CVYHEh6KLLWWk6WHY8ZYv2i
QtwgX89VbrxTqekKsuFyVrs86JEIt1jbvgpGjpBTNiYHG4l25w/Mso0+rWX6CM8X
l9DTGlgqfBIOzuHidMuljxDHgXxSsnD6cbqZ1G1y7pWHf9JwllncTTF2UmKJ/uQ0
FNpKrhiEi2/gWRn9NXEbxdxGTkedQ1HpnBIjDfA0Wbar5qoQlq/3JBYccExxqZME
See8yBFLUSyZf6QWTZZRvrBpore5dghiNBw8bxijUc+HOgwntwdd0VsZICnCH+GE
YFQCOjx5lyHK1rK2Akj5Tu+U4CFLb3umym5Ln+0HNZYpi1uoBaTezHoVmLzC7vUw
Hv5oPnaUcIfo4C44CsaM06a2KRxVDFKO55ejQpkbFoRWZjRamkiLPywQr5yr8ucn
80UgRLeHTeBny5bvJveCs7bQHzbSPPH72VFDLD78kAcOXphgv0qubB05RXoTPSoI
IsE6hN7QlnyYqQc6R2JytqAyPTIJlPdaWN9jr0qBbHarD4GUwsK3kRNpMQMf/Q5W
PedQCXC2fxf+iqJl0rdpcof5oNH0IvMqCfndrkizKlcyCItsGJGWEVhQGJTlEuG4
e6xL7a+lC2Wn+SNhX55P1ltY15/EFKICNOmusDmAOIITGziOTU06huRYuln6DHtH
4sbfIR6cbpch8gppJcfbC7o9AR1bGT0TBQvXt64Hcc75s6wcKWQdb3F7aBRz3hXF
YoTxRvC/k8kDEtcq3qScy6vob73BWtyrUtIAwA9Ix9UDjXfxPvmVXltP85zMzLT9
a8Ltbchrl6IPXRHdhhhXtrGt1sGydWpiw5gviL3CEP4o8hsW472bBi+eLyQ+jKZL
ZLQg/0XHSlE0/7/ILNshUqeokuZRQCkfYvHdQIo/CQz6zQq+sVccWpicUgVZtNUD
pZaiSIXZyMUpLI+BPvNwgFy6SaBN6xJj54d0pnumSdaYQVLEymBlEtAYXvFaJXdf
7qfHLGE5IzbsAe4Y+4FyCaeNTcOL23Okr+ehjcDmvj+D6yJdgD++GpeQuNKvc1sR
gVh2nhBgda7Otq8unbuSAlxvukrKdoLwxQYuIga5giypjf27Gdzv3rT+8TxyBK48
gF+c1x5hr4lcxrHpDBnpMgt0bn3Ozg2q3uiepltUYu/Bh8DZrb0+bFPKsBPmD3xW
vVkGLAmDH3NLYGX4Ml6VTXZkng+pogXs9CQ7U8V6GJK/xlCzAoaov+OE5Z/0kNuz
deKrUH/ORtfhRLD0hsWvPvBoflO0aKa6bk/V+nKXccr+yNeqGzFw4GnexaEM4np2
4biuE99cxxxLMfjSbz5bBhb83CJPWe+7LMv7Xsu4ZPI0Fqq1GfAK66tpzkRbKC6s
qk/ZdKYKsfFKmrEfTraUtwga7UDJs267vUZy7rHm+ktA8ZnWdNFtqP4f1ijx3vLl
KOvxEnQPb/XiaafzFLsJZqvaDjv4K5LnUlopjt5Zcz0vKWAXc3Zg8wApSMamRB76
Xvm5EssXnJ1ZsfXQ5sBU61l/6A3QRYU8VpPwFvYC4HoxSDmYqnRc2+Pf+6jU+dO8
JxqgtfpbPDzBVScAlq14n9VUQ5Wca7UqmvRTcSpv1aKQBNIoW31Wa46BtVcs1iOV
mrde1xs1anTdQ4gSyUs02/jTzlqkbaUBzEkmovZ2riV1byg3WOLybtLs7914Zw/M
4zWv2kRtRCFcqvNq9uEtvxD8dxFpJO9GvV1P6ErkZd04J+5QeJUgBV5rgzcp+iD7
7xgIWNVVfQIacKr3/CbCXW4464TK+zO30Ffk4ToK8dtS/udFuvnSWqKRDAIhnt8j
7fv1Kg3RTw0WyAkV9yKWPVZIRJxKoGuv0xP8g7Kf6p1qbQdhHK9XKys4q6JgOh1o
IOh5K4P/liSnet1oKYr5hxa/9/Mrp9AmRJCXVTItB5gRDOjPjP4R7/stb/2tSiki
hto37LzciH0iFBOiuffxCeDo8kxqK0VnJSHsoGWYbItHlFKsKQ42WjA6Yzfv6Es7
zI1uQHtoLXGDZGj5NRFY3Dl3xEhb9WHUqm1eYZI7vjLCgk4GBde1k9y7PPTW9y7M
4DOgpp2uqGyZTaA2udi8y1veGu4HYXiFxuJxIgTckStrki7S4IlumsGFI8doKlt1
yHHDo9+BDvtRDWpN5gpqUScWqGTfbLd5/ampQ5zprWR63yCiQk43EG5DmAcKFgwE
eHeaJ/+XRzlhyB40hDpS1Ars3+7sMPFwO7xw50HQSRNUia+GXXBL9mluetLT0XXr
+PUwhJFlfigSuptQFKGd0Q4oKbi5wqNVwnig2QU0jaVnQvgW8TCEQ60ZHosqsBG3
nEM94hioyE9gUD1NjwU/Ia9xiPli1uvUkaqOLz5tu9lpYnIVWQ89dWTnTFh0x4eQ
0yRy1Ue/Y9k1cGv9SeWGZnxx4DRYbxs7QTC9qA18JTZwcSNIBbxHPxUJ4ddO/MdH
1pReuTPZfD72QCc4N3tY7tvuKsPZ+yCzSITL1H8muvb/qN3Z898VIMuOAg7qYyZ2
2P956GQqrNIprUjQ6C1XADTtOgdl9pFk3+brKFr3zo0JG1KaZFe8ny10BCZ10NWB
0b76JNHB8xNsHIP6Ogd+uNL34z6Rk/saw/NOioqUSJuXyQuSDfXdpe9tKVx3xMFE
3YCrWiQaHkfUhPS95MuLVkxKUlTzvu4CCjlMJWFaTDDT2p91znQOAJSb7L4tLpzM
77PWIVsShWn4oWXFJWlHAQ0jo9NYDlkH7xgITBby+Uyv/Z0u5B/H/7k7QqrmLBn5
RUsTdS+8Nu4nRiOzElcdZHLystIW5ysvEAi2wO+KoxYblj2hMKaMtIjAuP8evZNj
PB8gHMQ5a5bBjiq9340zy66xWdfcR2LDA48wmRivcwVotUKKwXj3CXx6I/MPuIAs
PPnW6R/3u9uHqiNMJv35wechZfiJlyyeWS5kHhmVJlF489yoyxfmHY8gbjpS1v3m
5u1jij/Bp+x1AvbZmzLnTYMKmycUW7pT5xD3lNsAX1l/q24Ueotal3feE1kUsZAi
f5SZVbU8gC+OnypTIlaZDjxf0fn6qDjgWIL4JbgS4UpWEffxPWd9xbqOSDnsPlqL
26Q61ZHbkk7z3g/YlauiSs0uIzm6L1f+fI+lx8fDgVt4O28XtKpGm2Cj2AekszeL
tI5bbC6TI2TfJnsAL5fbezwS84y2Ch64VVvzJ22dtQL0rZOAxXnk76HZG9DIGBIW
s6PRc0RUsyLxT370NxJmHScflqDv9Kd1myCqcMbuY1VoGFbl6na/ht2PVtUudYwd
Zpqa2XtAyfD4gZRrVe3Xo+jSYx5+u6lvMn+5a0e9+vv0vlUIpRpucyNouuNZfR6W
2WTiF/S5HirYVSdfv2rA1/WGBRfP0rDRNvI+cpv6gsLhcZdbo0Ht5L/Lc8id3pR4
rRFveH6PSsDc6g69h7HZzGuIipbRDIQFCe4URO12Y/fcGBdkvJdxiGrnhUFHvaef
OD6zh2F2zHUAh90m7TNN2wyCV+HXszX66kSOb9S3RO4cTQ6d242LfzJcPWzy+xYa
/KZxIzF2labN3XsOmm70wwCD2PWU8jdHQLEw20os7eNxQeRRuXZnvEa9fLBiwzlv
4bWEh+G1OGjr/95PZlEyPHvf4vGyMalOSzyvjyGxcD4EsH1LSWjtzNnAx6W7zPnD
wIP1t5Fkck2/a7UTo+W/JCc2y7+iCzCvn6WoT7ESGXXdI13MN4z4bHPQKMb8O9+J
Vlrbnq1AYM6+KgOmqSyLqmfFOGGPXvDJQb7HEDmlgS+JXVl42cmXkxJTlErzRlAH
JaEIrRGM1xOWSJHTn5vbJa09m7hhUr662Uxe1zsR3yLN8lZfVfcgRoUtU8ECAQVp
Jv5Zqnt7Pm1CuverPvx1f99LPcEsijx0Lw+n68LG2HZD2NmbLQc7svVcMKCMFRF0
IzKtCUgaa692HF5KwBf52vNfnEj1LX77GucjeAXiZ3Exk55dkmTTsgSMQmD8kEx6
JvoSLPohMD0+blTMyMR9c1rCZmNDPIs6NKOQMsIul04IlSLmZbrKHfo3/j0M53Ur
4my/ps5iYVF0MZrruwra2cBrlEhgA5obH5oBHaEka5v+lr7Y+4pMPh+qGK9uNf2V
9hE9cTLXH0Kz0CzK0KJRgk5epvH9F2nrAvcys/kvAFmnaQuMN6S/NMcxzEBNxGzE
+nLqI+H9YzEVpFLEwQbUmyixL4whH0mpYMb9tslrUtqI7v5l9MM0mBY8naMeGesr
lsPfa5QFGSRu0MHPAk0wTnL+YOlW+XYQyLlS6VRcsVsW2Rr+d138njTYDZNrquHq
O3unIPhEcOPE55/lkUgxjk+jw/YJDiKxj29Q/QFjEIYoAu36w11inxkYnScWHsae
+UKIg3tYu262hnkNDbi2n7mtDZSPaldeWUMo0LEj2E67Go+USeK8hmMa+k5G6XA+
4aZCdhcW0Mfvt5tHr0Jz9HtQCgUZNHmeKADUQBddTXgc7czU3mJ5izUftjwqJrjP
bzauyRSz4vIBWnMO9QDrrwmdAgH7fCkNASr/kp8kwd0k4lyNGJhvLJnM8un7r1Bn
7aEM5G3Iq6hWOa/0DI+0bbNfwsBasdG0+wA/he5Mps2cFqWiepKASjyvGBOCTWpR
bD1vorq2qwH7AErcA++fdczysOYAeAxrqIz+DQsm2qi4HFGg0l+X4uyBp2Z5Aa5G
GkUZ5asI7p1kc2vnw5Z2icvksPmMIYQDun+20KrEvk2BXSD+9u+yBVq4vkf5iDjq
iN+9P2I3Vl8pyuEF2MuCIEwsnqEq1+FFZ46bTOQTGtAZlz459p4/I/KrQDQs9br+
ecmClyYhyuOt2e1ixyG7+Q79DHhHnf/y8Tx63VLfG5Nm/SmGoMptTuKUGwi2SvtE
2V15sfoF/aVOg8lcgcVL+3eK+YjBm6AJKHgoSui/t2iTv6+/gEGkYDK/7CvLN2bt
xreOUI45spooMkk9djbqiNd/SW2Un5+irW3FO09+7R2Y+W6IHvoD8wcObiTPHo3z
SsKVi4VKB+wK0hCXx784CFXujBbUfm9iesgg9ZvZY7mAfNSUCjoH4I3++MGOqECF
FBzd4pnUomVnor22XzKdQMnLwr+N0mbk0WPcGhK7IiAnfuzqF2FEju3uITw98QWC
qEkgqWYd/WP+yUGzudx1DGKHqNkspIR6olOBuo9OEl9anZEBwT/Ee8G8E5obifs8
IyWESKe4qS5/HM+3r8EL/hX1c+S625AMmDlCS5lRoR2O9h20wPAAhgAM3KH06lAh
mlgGwo21fRmsDkmTLfJ3jz/0w7/Pfkv/rB8es54O7f4bLEyU9b86rd5fMs1m6Xbo
4orFslDjTnKDVhPYdSpctuu22ClpUndp2fHNIL1ol6n390EQBKAoqKIfRNq9Mrwy
KdCArM1s9bPaeZPyNqe3rZC9xPrelgsgsXJCCvnStqt7PcM1pX9/lnOWpl2Wz2Uq
+ZwWWaX5CExvvg4i5kOVsDzNXgI4wSj4svlWp4wfTLnzDqci1bxeluO9boTBVFjR
Jyd90D2ZtlsT8S7kU+TRbgEmHy3YcHY/iscva84Bp54C1SQxSb2NS6EVkZel0Z5V
WhuIMMK4hUsou+ZM0NMWsuh4kYgHoAhgfKSWJXiy35rEskqloSg3WgD5BR4a/AkQ
atE1YSS04oFRE2qomm0azCUp36joVGhbo09J2BpAvdsvS59i6MuXS3RZqkGj8AQE
7tN3tVL19tIFmTntHifgYiiCzDS1a937dGQif7kl1u3MVOEoHiQSW17E3WAQ/iH5
parJq55XjQj12yOQwjnJaQMtukhAbGnhC3ZSrKlYKlQvA5QdKwdpBi6tF84EvIaV
D5qniDQNnll0A3lNj3d1+fkbxK61UveYrsTBgZF8tBk0jSOC/KJm1PoF6obb/yCs
cmcuJpmm+uVhR5owwsDjb8QbXkmdVsLx2vtBPdxHj9xR1t0Atu8ZYLvpgOSbehCT
eXZpi0R5kogoOFDigsxsSRLgI3oHkCfCy3cQ31pEJmF+y60RxXnpKaFc+OfmOyf+
msAGqET0KWc2RtyAwsPHupVfOgDHmwWh59pOGSqMB+zdvKSvxEeS/c7jdBMo20UI
pajDWp4qKMgrRi4+y09IiUVZqpwHz0EGbW9E0zZRoLO3uYk+vX04cTfGL+1Gs4BN
TSz5SyF4BLcpCS0vrR0CE7UnYtpnNR8x+rjSvmGVUKAm98Uye2A48QOwvMnt4Dgc
mN2k+Hq4yhgAwnGgVJLbyrPWcVOb9Px6NATLQXjBQFTNVsKGcgNsnIcruDPWc/+/
eStPnJmy/231AM9UAqTTK9sOX34eoSOv5JM/9++PG7AVOmGlReODW0SOot3EezZO
CYQIt2o8ceWZxUtcNV8BaxYTDHtZTOWlPEpkaPkbI37JoBCJlddEMA5k4Ei2eqGV
26gn/xWQnitnvX1LCZHOXL34K5kfIrAAhN3yvYRl9RNQ9jYh07yeFy4q6WWi3cIH
6fpWUhJ7/1W4AX+u7D/4Z29vmLLJoikWuHGf/I7/PJDP0oGxrP548eHsW6OQJpVM
Ec2Caoc3e1qy221e8lAZZV/pG3bQNmp0YI/BTlwWAcTit1IilfTJzMVQLgEgaOxK
zYCQlP/J0zELTFwaTl85OABXxYpn9dcpFYGGOWxUKigtVypBRJlduTh7KqqXFtbN
1qcywK8j7wxhMiAxoaAFKlADa+bIKicKtUqnVu+4mo/l79vBpc4ermls3WcWOTiY
0Ofe12J5fB8myBd9sUlCJL3txEso3ujct4SnKhvx5yRorSudQJWcdVTJgrTnl6oU
nfer9qMUWRPtZ80OYcRf5gFQaSxxLJjieCmegw/UpP3WV9mgG+Ews3XdybIm71ry
GnJKLOKssnyDrYsHETC0ze+yKB51SeOoBeaeaHiAgelsyc7czB+VSm0otSJ/hxPp
ti/eEeMYZXY9NqWMM1iJ4kA24SrhDc0dpB5ZZlKYvwjgC2CArcxemzKeW49O+VnG
w9irDeU8xxcONfN+1v8QUIgZ40XwQMwXV1/nt+ljQ1FDIcvlDioLqv1idW/sve8I
siG9EmdzB7FutOPs2RyzMT8NcXS4NqwxkNYxiQr0iAncVfM4Sa3kgfXouyIeSXNG
x9t7OCTbfdfyDWYkY+phTo7cGJq6CoZl2dov6cIKquX6Birtoc4Nim5YBHidF3RC
oaOxYTjWQk7d8FH9W8cbtwD4xdgRrbkR6q9eJxAnf5o370YQmTw7jWOp2sv9O8oz
25dS5kPrHyek2JqaAn0TKJF1VXtvIqmWN5xjoY62IVRQUgxPFsVNdnk3vIKWJqSm
/iClwTtmzNXUSPhj4g8pDhKJ6M1bVT33lbvW6KnCH8FEpKtNJa1qo6yyOZnbmUKr
LZ1SMd/9oA3erS0iJ06t0WdaTqL7tC/DrfudKDL5XSxSBPjPNts1nHTDbPnxQNwM
FIfnCuRMr/fyP3FpfMSytnNoV9DE8Eeq3ikGvGtmTyeCepUbcg3oYl01o63G9++i
IAejVcW6t3Lsm1pewR3Z+RfLBzSUCn/0/m/6JZY9kuI/loLycK3GSrJc8QSPg4ji
v2e+khbiqdUJ/vhq8PXk0w2xYda1V27oSzn2WjnlImIcsgt9NcVdkgEvjRINGGrR
Jtirhi5Tkw5bj1EbEzwyHH2BLf8AqyiwD8KA0u+UcIoEX1wbluczPbbCqzigqTWK
a4ftCpzzxqt4H8LlRSoFxmj2p3A2wPWEiSQ5CCIv755EeqDnJDD5Ne6O55fWEV5h
XXxGOAyFGhjFz3Vvwy/TtS8lEr5fkbqwK6A3cnwnP+ejFkqdTCGafR5uHgajlwOO
rS7BKRxUN+JBuVJmxbZ0F9/U8hpagxRZZH1wJP8ReHyB8GOurorpKT13l9ITbY5o
aP8okbIZkC5s4mf/Bc7hWUzokJ3T30MLzPfek9YJf18odKOT1Ez0mqTD5iVm747D
HbyX4ZO3P6H8IhieMyKk2gXASUQuMhLZGu81FjkHlNzgFivsgoo4ggmRSRKn8meK
Evt/xicmbu+J10+qOkq3u90K4bZfwi5N10nJx1QlTZLTG2SGWRTOUwzJRXkNc+V0
xkQt4CHSFJ0arQrAw86MyJkStZdWARQx+iAzgbc824+22kzUS5qmulG2+18g8+G7
+aHA4LvtubzPy1983eJHTus/TTLq1GYNXGvJwabd+IIyo0BKExx5ORYs5xMdn1Ln
p89eDElwR609B5t7RfLznah0cYX4NH5PdoQ4c+cf7cuxEG/+9b10nXnyqzoeTch0
g0ldPeylGV7NGkEDiwsa3g6can5UDV2YUTxxYtBiZRJ64cC2NYi0dlEKnFu4hLF+
OCDazzaRgjTA7mpWZFfJuObEESWEy1aidme8uDHytgDJNt60H74m/2q/CjrsKG55
DCC/Tux8fTavOJoyFHGFtGybCR23AoLSZ0SiMT4nmElrOqTXLAWFNCs7IAtvFrEq
4CulFOWOEdFFWMbOC6Z/rZicZwvzhcAyUXsVQtNgtpiqW/PT3jTiJrTQSc95dlcT
M+Zrg0RwEvm4w7ln33+rd7qmykND1oJffR3XR0Eg9AtMghx8hWJb9HYtaiT1rv3Y
zjubx8LbWifkejnUb9C1nAJKE+cFExANHL/msZjGw52LsXzjpO1YB0OpfgH7ZV0U
Upqjs4QNAM6iHvYajFUS7tpgsnA3y4cjzFOr/GYuE1F6Hfdb7GUoIJI1jhN+hZkq
lQ6F74voTAyZmQo+GVqJhVLhi6NZ+/TypIcZRt8GnUoqZt8PrS6EoYpujdPVRwvs
JuMZNxR7OpcCtlTxp7KEq975vHp3CIgrETbzD7x1T474b1TKqUz+6l+dJaoTr8r1
yDURmp+0c95fSGyGpTLVUEgYHF06mfdMjzChWki2wwR9qwSPsTZFkV5SRxVV14de
1ak49ZcpM2Gfp6sb5MO5dqCr3tZWjM/uoHrfRpB4TvkWsbN3RLhwaRWd5cv43KZr
qMBoIq5QtmcCnIwMi9PvF5HEyug5XLOq220qft/M11WKlJNh4G9OljPIBQw0dSne
IKs5sV+8H3eAPhHapCDKP21+lOzUOkQJnKbtp9aZbb0oeyxEkxBwD/61HCZkjHvm
FXE73KwdeB1MFojFnFOJA5au/Pvj5HXd6UKMytx+078/2Mtfd8KqJCswB1SmrxIT
B9HMd7FvMs+hKzdy842T58ULbGYRjugEuLyyw3/yzuMe9RCZf6hl6ctVfDaLScCx
2nspRnp4BRDMGVkdkkPP2xIqtZTLPYwSwTwkpnimgWYZd7Y8sYrhx2IXHwsHjf/Y
FzfX2Y09ZRl+5Ks91m/JEXqmMsIBZ7Vr/rCPe/eXb6bPSvfwFRNFLKz7R7HP3/9w
i0J4dlQpO3xVOr+64t64TT6jOgow+dwXQtbZx7bDi0vWLfDVEzwhJOp64zqFa1EW
zNLwOKaXq1JAiZAyo+65iBOa1vhWu6ouGeQ8P6A5oDlPg4xjhtgND9PslJdN+Pg1
fMGthFiY9uJUu+wkg0ICIiHD/IsKuMfoC24WUZ/XGr79YBdbV2kTKL8LhmLBmoPP
OLLg0LgzDOOiBA7TV6SUnqeH/y2Vy9RW7rpsIdHmSdx1cQq4E6NsC8Ac3Xdp4CSd
lHb0WNsStmSiJp47Z+pHG1SJ9XfqxJcNu3FxEmsvbB7ebBtoXyj95dkmsXMNsme2
8QDximqaVXKgSTebiRUOGXlB+Mk+SsaVrOtEyTa/li6o878mEomnACVlv1NSTjRl
W5prdvfpYUXceV/oWRFRSpfAQ5LUQc3q5JXwRY969j22o1aCPaiHr8iOjS4YI2Ik
GDdXkAZGLndCQwcj6qL/8S5V2Csxx/3o8Ie/08+5EFtHoUWmlY8cd46M1W/dZ5wt
3SWCVc8wI7lMs9sjaVewFq88kKO7aAHpAMilZlXgNbYxgmxiJkhggU/C+pGECNOD
a89zXyFdIHm0GKXUg70IpY6g1EIm6Shv2Bxbwyo36asNTyGjVANFwrnvvk2Z0GJd
BN+o2u4w4skjnZf8Nuq69Ib5zrZuokvNwueXvulHnfC8JzKUZD4kcjmKAPdhpGnx
sb0TG83YASlY4o9RavCgINESy8ORjcK3m0AZbR+7iqMCkeh83AMssR0lAzB3HkVr
VR1IKmWQYD93qtWbGzRDvQjyqYyEkzKLx+NnORw7Nrl3ucUEx/CKK3nFM6fMS7Ym
dtxENBxyXqNyHbGLuYaSi2Yukb7LWh2dgbFPHNx2kjUJeH7DgQBbp6CCPyZuuIbk
mIOE31a5p9hv6NdBGqo48IbQdU/T6TKiCHs/O3XLov4P1gqGwM3oEmGRw3/GsmFZ
ByzDRaUV1XKJIzeKQK/BsNKFpEPm06/4pCCe10rNv/gpAxdYsxSZjoGKgHCWvbPd
P//JkfJ4hm+KikPqZ28GtV083iVFuNmClkrMJpPfrK27rpFVc7NxIYkr35h0PJ1y
e5aik4pNBOV6/U1QgMM/Q7Jx5NSgFfyNvzavLM2Fuk9/Mwnd8/A6YSmw9hbhZJWX
JUFIVV8QL49ll0QoibCIK2gdBktDBZkpXID05mjkA1fffmWSesU16TNlrZmBy42C
J69NSks2Ddvf/+tABGnG/8cv6ozgywXcAhDWc59uQ9f/jH7zFCNi6jFuyirbgcdu
MiZch/57qOchH0vJw8G7aQJIGVWfZVdGesuwaLDLnVJjHWNKPiHrsPJGAig+FBY6
+t0yBkRlftbFV4ap/6RUKuF2ZIrZsoRqD1z1B/1nub0SIMv5AU+5quVhu9yC+H6P
5Hk1545fSA2gkteSF525mMCUgmHlLaXEhtJgVX4nuAjiGCzKzo/F6ilI2ma7xKZM
AOkSh5YF3093FIiC1TsS32wZzVXPdtiF7IWsmWtvRTTXhyjqKORKUxp+wRPGgron
0se7ihQGm0rtI0zqgrreALUisTSV61k+n1K/iocV50pWYFuFCFeNJS4Vm9NOQklq
tFZ+H35SlKBaxTVIgePZ+mWS0FnhGOwUMhFpAnUMIxD+xfrEgtAvpRrFLmZo9LiB
auAXmaWfp+uPLMMVeOp5KqaUNQgteFTEQxTKmbZcp4G3xKtASVs/107iMwVRhUC1
Z9uMYE4/GM6nbg3iDBQqaYWIHuowafBOwDlVnfwwCcmC1cNbhAbVN98HiV59PG3q
4/ZWCC87ZrNsYetDFfhBTtM80lsyOqJST0+0twvy0OAROHWbLfxIaZNRm9VTvYIR
cGyJ0EFfCjHcHbmozIP7hPCJbk8C74QjrVVfMJ5xmpItcdmeRjdnCQss2bLaGGM3
9uvOF1BtP+zYRQTjyEFNwEvdC7VT9sVoBCIRLpavSsfPioFgkRAzdC1l4P0mH7y4
uvlMfsjo+09UADZFd4aUmCGepwJhCR0XhdM6xxQmDOu4jYU6u898IymmjRWSbXy0
TDlFc+HJSPrPnQewBLKBkBn4nrmQx8x04DTNbhGzaVxqaesUdD04bON9TrDbcsm0
AXlTEiMf54j4YmhKK+Sg+Gjo2FfR+VOqXZc7okEV0jre/fhZyTiETqI940Vhjb7Q
CJ8geUL+JDNn48eDrBX+OGKy6EYZ0KiO0ERB9e1j9cQYD6/k7JZmwdCkNJoMxzU1
b5vPtvxmbMMVdb8ulR5Ojjsz0JbyXEH331TW1beBz/vDDM/v8eE+ztcd40Kn7jAq
IqE6oYJrbnO0UowPA0EokXJDQ9FnIGbewDwSlmKDVsYNQkVlKe+7GLPLEeZDvR1D
3/tZlv7TBHWb5co9q4Pv+jOYzMmw+iatQJfhSK3KnMlT6cZ9j2V8jLB3mv64XHME
H9Peo+wVpjQk4AOxUIR+EBzfpdUtV0MLRHRu0rvOJy5PA+dZ2UY3Ku+fhEFh3rS5
l5peX+rJz9viJElPu6rJVBAlDxZcciJ9/RKVebEBCWLD7eP8DjIVimpC9g2WjVnH
RgCHhuevsrlAri9HlL18ci8di4aoWU96jVuf8rts2428SmxGB8epWC46Psd9Zqdy
rrvpvEgXO+UTy1rDUsnom/Yzmu4NELKHd3/IOZDkrXLTkKL8C6PaNOPjraknwemH
3XjyNuBQ5HCMQ5TP9UTOn0ju0FXEgteUMO+w34qAtOA/634xQB/j3GnswuP/Rnu4
hM+yS6w55yhPZfYxBOvNeK8WJQeng+Mj9vxQFRP4PvrEEUiGEBuGwvrQHaA6bJXG
bNBUZpSG9VLArc8Sx1bCfg09BDrh7NpZ38rO3RTMUB4AIRluW30lRMu/Iks1ya3a
FmdYEyjv453t5ZyJM8nYViwxO+VXjMsi0M4UjshyiZlkjRBcwdqmOmhCw/FAPhqM
gNHmARraDqH13LI8ETmv8QW6FOdtQYz9r4RPC9xdLVzJVVgFxHXItcThUxf5HGug
hhQo6kL5JX+TEUUDDRhmJ8AwAml9S6Q1K8HTIND1IxWXoa50rd7BYhp/mppQsSZg
zrhMh5T/bSzhg10Ji7NVSqbVKC1C1Md0gciZXpDjXGzZRcyNm6HOSElzArk89i/g
MlzTtPVcEG0SDpAN+kuOr23iHV1v60YjNOa4cG3XhXaWF0aWvWdsrkvunHVzkPQS
HN/25vQHTHajpRhWyqAOAQAwiqEM613XDb+NvXGTRxwsrXmedMSjbQzcoKDE0B8t
rgkf00WBbcYeZPUSspn0VgFWt3j0NyHEmFw+HP2VVWwoVnLXQAWuO1KAJIzJ1QHI
qTK7YXn+X4orUjbDFtxFLIPtmDY3PLUp0B9ucAiONINj8ZHiBXNG6d8VOeqEgEuY
RTRnUv8tzvtyxM9QgbYFFNNSep6DkiB8HZDRyY9f2x/WywuUPCBUgT55QPAdzXVE
ia21jGUt1+8h3cUFz5RnU0kpxf4avABPqTdbMwItlehXcmjxiT4k23yEXa3PoTD7
gyvpsW62JOWI5yoNhDfENck4SEv3Byv2Cdf6FH6npRfGdLKRYUM97ICUC4OwTNvq
EmtTvgStlJNCmgCZv0D2FFpQnD9rCfNaw9QaOPw2guJ1UsICSeqvlZufC99WA/MS
VzjAgpPKGGUMjfkRJwR0FbwpJPCZkqQkLTJouP/wIJp9yMkDTVNx81d0+iNoVNC/
+tVHTonz5CWYVbq8VN02/QI7vTlWcvo8xqhk3xaA8A/JsrkjXk0zTIm40SAChLqX
yblXiiU1BjxupyyBnN7v5g16+6GT0MUo/eISbGyp85huTb/HclXdk7XOwTMhnuOJ
/KcKOyf/02RLy53ssza/zuFOC8sTGX7wORyXxmfZQnDkwlbzTDgyDdVKh/Hx0xXH
k+0i4IcWuOwzeiqtqjIzgcHbK/D7mecUBd2R4qzX/laNGCtcv+2VRJrSP8YcTi+Y
j5DA+ayiMiipPS3qSnjjvjyVsVyg2avflK0XCP/Z5EsarLAeiq+SKBPh6q3/ZYmc
352ARKsF3kzIErZjyAIoWd8sF6Jwwbsc8HXyKQ72cGfMnhHlOwM2iJsXUDY1cB3b
MfNWPHJ6Q9bHCZq0o6i3nA+1mkm0yLGNbPJ2iAz59GfcsMuZ45O82uLo235gnld1
oBo1BfUuhAkAvawNL8gdE+IgZQYAGa3xYoCMR0yqH33aoaEGE8gW06H3uIEiLu0g
MjYnSeBbJB32nvqGHJjQ8hVJieoZmkCPjAQeZ2QhZLJkB1Mw5dPUvtUVedY0Yz79
0aGnELlXl7yQVtPfzwwqz6UmC0Ja+sdJNLGUmsMkC/ipi5+fJDRynUQjKKkkTdQd
h6I/Voj5NM3cLJD2ocUikY4Jhwyy0A47bXTVoRZoCV/MD88L8han7/oHKS1sFokP
FpxykX2q84sccuCH2hGSGpXqgKxuaQGy6kmWxJ0d4TefyII/9xbFd0mqCtVLtURB
xPR763JinYG1KlsSsRdHrvJrNS6SEv4DXKHI+ZxC6wa/1H+Rqv6HhwnnZ6DVOOwz
5owPKcmkpqndRUNE3h2W7vX7UN7zJUCFZtoEALRecuwTUCOapgQnPsSqQo17mn4F
1MH5VcxphBYpZ1Xa838pL7nLUEijjV3vlo1KeDPzhlq9wjlCrE+7Fp61TLgz0M5d
MerOx/uAw9aiooe0FfCLjCpbYaN4iykV7I8LXInX1Bpe8OgHv8k0Nj0FcFsokv5B
fNxmuwYx/hclESR9htr7QDW+XKFwHuEX8dfnDBq76tg/T4ZuLmHgUNhy72Y+UKd0
B0hOOiANpbtO3ExS/v/86CdYs+ywdJNdnDV/4m5vvVYht3Kbq6VCla/rVNRiphCh
JyYFVs9eQ4BwehxE42N0JiEn50ykTMT5U7pvuL7AyPZZLMln1ddYnM9cLyQ4uhkW
wF3RIk6dtcytZK1OK7j1cee2SnnaG7//Lh1wOphyAhpdexrUO8L4zNCEIEkLBtmm
Xdz840uT2w3t8QjzWevM6hPu/GdoOtzOp2hq2UbJ6Fbs3Jy08Ma8B38WuRrEPCc7
sb4CizlCorLofEMLhUqjI2a75NPGQWl4/Na5vE2lYiNxnLtt6U6/n7P8cJ0PA2hE
/nKOn92Owf5IFCJ5HfLTZIKpzz0xtptX1v92zbA9Ik0h5AFVla+NjsoZRXgAYp5b
81bfVXKpRvbJZBVhLSI6VhzmlkHGJ3LSORqIL6Q/dHU8UO3DoBFmxBs5C/LfZJqr
p+B7c4v8XuPurN9wmT5n+inzV1+C/wReXWnELmy0BQDOtyHIydltXj6S8tKupwUh
C1Jg19AT+3odNHsEQw7yyMuXLvemt8v0UYR9lAr9gLvRrHLElZD1k8DFhH3n3+YG
Nxwq1RbBYjYZGAKqslS/D7JCyeKWAXuQbNPWAUTbp0SQ8uFAuLuwJdzGy6UJRHvJ
S2N5IXJs/9ERvjFnrw8c4rwAlxEe8RKrmbTwgrC0xL67AeNQI5LciAhTVlz5PS6a
X93rCyVwrVzBSGTM3YKp78WSd1gdlQwV6mtCukCOUOQ8SUX4/qEyONl6O2+kiXhX
wmIFqkYPevyuaHY9ssWDzBfkvUqTzoX1MvXEN8EDEf/s+0HQvsxCIgIAfmD+SEmQ
rNZmixl0u6IGQE0HCRfwTJPyyz9pFPNnpuQrk2uYT6G2jKNeS6dKe2CfoVAcKgdK
rWU82czKCCyF9aGW3GAJSb53RY6/sCh1/nwMfG+G2Dn77O2JAptnECkOFM/NC8su
j9IGAdyn+/SG5EVkokiCBwJ6YilWW3n164/VVT6aClwSV0y6q7GCarp5g3NNBcz1
cG4rIuN7cDH0NIUHmJxrr5KUi5tRXHuENOe71tSlNF2t3nhxm8pGjmRsg1NrG7j6
bur2bevjJLCQVlFvtZHcO8KhbwNcOLUSwUm08aEiZcgXdUKCGkIyL3Y0jOfB0/VB
RKcjNxe5l234DQ12TCotxLFhOx3+/FdzWV2sheclPcUFx/P3kxP7rGFXGsDPYsqt
AWA0xFVJk8RkM/n1Nic7oP1z3dzt3kCY+kMHZGdsGiH7FdD293aS3E2b0f9s6mhz
ANYsUoGl5b2H8lbJEcnUcuV5X6pgnZmcOxgI4ha6+yYFVPGNNqHt4K9pZT17Y2n6
bQOnLbP+E6OR5oTuEZPe4AMWcMSDr7Y6EZUHlAfC4O3U2aDNmIdSuSi6jbNsinv4
UJfXy5YCN5mvwbAGz5tl79OkV6nD/eHpcuR9AzHNotBRj993RUc3YdDPLO5PJQtR
2McXT4OfVI/jyId3m7uu2j060m8LG0PxZvsAJ2LTy+PYMGC3DBmXobUqkUbyf+1r
A3OXQMzfnaqtGLZAuw4nFgJQRkCONT6XImDGsEI6K4iVM8j6NikTBYRD0/Gu8KW8
SA+7AGkUP+BrxOk8jKtMaEXAE401jVn12aY5u1RXMdSze/0mHyjNR7ZXf/WkAPXy
O39Qz+W9Rxgr26useulXPabrW+FpCkc1p3gbzlUfHk7MvVri4xfh0kVRltKP3HP0
WrpMBXc5UC5Ted2BMEbw4AM+ORgzF8oJ5bLyxG95RPy4CQZCFhIl4wXpiQRmpMu3
bzBUPkn2jVH8QK9rWcnBSQEXeMhm8W1mPS22mCJUiLuM8WvlmC3DF6qPoA7UXk+V
EiCuJxbmpqPrps8MLZxg6TH7l9zChW+junJ2M+B+7wRosl/9ynW9eWgIYait0UNp
qzoTI1WG/cxtG1UVxKphXIpd6NMGcU1ewRPycQPDncwZ+5tXHL/SHkWF4LeTHz4x
/z7JcbRqn6e89v8gJq+jz6Rb2FsVuLh+QqOQmSeGusasJxx1WNSQWU5216hRdyA7
gLvASi8I3iFdTrh707imyDxe9fuq2KrdGx5iNc18Z1MCnUHXffb1p1o8iDOK2FMx
3GSkTtVBivA7leIDkOSCsOcHxCQg6enIypCfyKK0m97F9zHofXPRxXnwm00sz5VH
abQDQQ8TqPiZdEmDZvLBGbDAMyy0MhGYRtz3IDozEa1HqJe0ZK0GT+CPmgWX5veO
iwmbCQOQzm8k1MGZ8nj0ELFyfiByy+UMGq/2a486dTBQ0ex4WkG+W2bvTQxCNBtZ
ZTLsx4owpuWiQN5HT9OiiEw2IrYGbStkwsOys2fvJlwIpDp8eE8wmToSbB2vAvKf
95az1HBjmuwVlGXoPRHH5nFmhlYpx5FNGMZXatlWRHUpydLr279ffcQeu/b3Zr5j
fUo0HxbiquBOh0UANee631gB9P4iB3RcvkcmNmpVfBP6UqT8tYNdfoMJTMfKHv6T
KA7GXgAMIGIKhjVKSodsft1Oyn/+7jItfDu0MGFTzSsRSqQ15JC+qDGKAEYU6pD0
M8PuhyETirDsSFXJuhcQRuHKJs6vCN7PghhNY3jnLmLIAKDN5J1QR+RZJY4hUcBt
b9vF6SIayNKvkjmGhW5X5NoZ/Jx/zfkc30nIrZXpQVGlJOMVMFFVxGzfU9OnFNkS
po5fJ7KF0Qsrdh9kFGwLjhjmal5Cji2JyJZzzglMF8JIGZg1U3ALxtZ/GktkMDjG
KriL4KhX7zl69DSjXS64XwygRwb2/404VJ+oWvqbG3GlReQR8mZlRhe9FHZjLvog
4MYkUtXo85bdQv65AhLv8Qtji8yWhpBnegLRK4B2Bjw5hk/q8baLxYaVpzGRH6cY
q/Oum9er6k4yRmGk8kePzNglWoP4fPM3jtlaTfxFg7NpgswF5Nymj8HZTcxjJsqE
TbIV59xBNAyl6QslKduwFeC8x+wrc0p3NpYZ2FaAVfwPOg4M9F8QSEFWMVnFCI5A
6/PJ48dFaok09pQnJOKSVG8VsdFM6UEodx9fBuml2193bwhCo+FADV0gvBP/N/tx
ewjrP965c83fV52jvCvlWvMJ1ysfOpmhTw/rUkLRpLmu0EMWr0doXQ5g6fxBwBHn
7geawdJi6s+RgCzHMMdcOIXqFMmcp9fqGt7+5foKv0BC7qs53H/B9faiKq6bLrej
oSmGRazIfFPB0dpIJuAp17yZw6am9DPSgRUKn9/a8+8dJHmsDP9LVadZDeSG+Zpl
GQMakDj7J+iHC6ZPFBHf3geO9mqZVDye81CK1xo+FW5Ne8TAkPw8mVJjfgNTo0rc
fAbl9RVw3nNljeQ47G5nbd6kpuKU5hJROoZlkcUPb4qmeEl/7e9VMVc/9k5tT2+A
W8CIfpXfr2eGHF5WCn3Rpby/iThzS/PnhxgWo9jSdj/3gkr8+GdqJJyNUOv4CxhM
N+5GqNP7M2CQvXKUZe3YvZukcngz8MMmpqlCWqlkZiBoHiFqyCXHL9R3lS/3dOA0
FT10FkjnixS3x4oevS79iyy0JAwDGvFvCMIbAyxYhtyHYvdKDrhI2A9YWDISVmi6
5B+k/lGErk1pJzpWgswBJ7tbID+ClMuFWntdCpdnuVNO8H3hmlfRFwXFROxAKKoB
0E84BDLUWnw/fzGuY6LXHjvhDsZdZtEqWf5R7PICfmYA7LNKTER0kQOFGk0IAkYc
T1AGW8H+g5XxEBingkBlnzV8CSIoi8XWYbgGBdlKMmpNnG9WXdYrkDsL03gVZYvJ
K6l5mvvY7x3QPXhF9NyYMXzpPcGHBfIOrTm/AuYDT3pB1viqSmB4ea52uGC3kTIt
eHjKJsyEzSe+8QXS5Z+LplKRLrXGd6ci70H6Exb2BEP019uHsYUt2Olf3RnyK69B
+FW+cEI8uStVSWxnz6FbgqJV+PnQLmWJ6aBkH62dLtdev8v8gpvvyIRHRgP1qhbx
OaH3RFdouw4SLxcF7r9DOLggrqYKOKwya4iOICcF63lJNVEwqkx8E/30qzurtkLI
3q/0kXzL+jxHp5XjJVtDrgTj8opdP4KxnNdvRa5AKcTXjJznDaxMxrd339QMBYMP
FLb/O8RyZ2Q26SigMmCcUFySHSD+nDX+c5V/PYJKW4E8ZjhrqqMpCiIc0iAKB7YV
xr6asCAMTBN1utIwxEq/lxR/0SqxPK7ZQ17iiuukn+WLbp66Z4UJNnPyVgN5mpZb
Du1Iw0XosC0DlTXeYcG0Efn8FO6+2ez7nmICThCrQb2YeZZK4mNwkb4yOF8osfLa
mXIiaKs0cgKgdbRdNCxADc9MypAb6yn3VlNoVIMDAbyjiEcBCg/diQZ+M2Pc5HEe
S5z148Qc1U4y16xhO9AAMbfo6XnihzJWLaK2nLTxYrkq0iN1lafcJVJLyaOqVmP7
VeBRUgOVD+y9yYqZu2Vd+FKccNQmbAgmLu1ZeWzuyDbW4/uO8lqZ/DMJbtZu6ndW
71y8cznp7SFhMfSxfijjyQ2bMq1pXCCeBX7E0UqYBJA9Sw1AaB1l7qQSIimzHkcv
lrgX7G4NgiwvWFBJC6LvBHpkJVRSaPaZHD2nde+jfv8TOhLO7bcLssiMSy1xpW09
SPRO/lruyWStzbNvUkB9l7T0lYhWDJ9+il+eF5qNyTBm+ZeXYiVmWPq3mFYa8G8q
YfDVFFU68KwcBEazL4f7GrjowZ88DD8ljhxEV7c7xs1xuYJumUUqlUqyjYgMpbFU
GrIfpoi2x9KUgh2U3oNSO38cd2X2NLmoSHsXh2+y7kOjafqe1yj1u/GtJySfyQH1
c26vI8aZmu9WN8/nSAPjLJNuMDiFKz3L99QZjh7LFcxWQIxFTwirFKcUNDg9w0Wy
dZKOpLid+r0tfeFcCZnxajM7zRvaWwbH8z3UEHyE//mMX9f/jU+9xmoNJ4Ho2Ijr
+zbHvTwZyFhWYIcP2Dq0hCYF8dF7H/93OOn0xw6+94MejQ8B+PH1eveUhi1YysQO
a+U38el8vpEADSpnDonz6qmJ38Rv0rT8J5fYYBYUXtlV/Jslz07zHaw5vDlWAS1Q
ihtpOx0aItgqEdBEMazVpxlYQBehWaKQNFRMFtECGva54t24kyE88MVgKaoWa4YZ
GLP0DnthsnTigNNgTa0Ajf288Ee3oM3l20VmptMANTPyYGBqCV31IjEPKrbxT5/z
qJlGYZQYES26Kq30tGS2V3D7cQpmviKiroGbsobH3dJVaAjxf+DeKYEyWL2OI7I2
ia01zuYsFdtkqW27STfObutot5Q/UCVA/FC/2pPGJDQYCxZAADTznrtJXeaBEhaw
VK/sFMNap8YtziRa22xCj+jIlgTOoMgGRp4WxnPyR/GiiV/zynPP8XHdAS3zflpA
aSS/0bjosXtS7qdU0FCNE/IjeoVRq+mhS5EJYeVQRDkjdlL70LgQj/LCHAYrn5gf
cZEKWb1ML0v3oXyyeeIeRunT7F3jrCNtcON+I5DY8Ol706UsrmWXE89TzqkuPyl/
YxEsyhdxUTVECQGcV7yJ6aoDwaILnR/PYOwiM7an2pLojft0bbw1niYzFw1i5Ywd
lVyeLo7aSS98427pIIXnN+c+13sfvKUgnqD48u+UPXcMKUYMnt/jD9t3jFF1ma39
/FOuEw4Ygro/7coL//2k7c+RdYLXpx51c+NWr9CeBQ85MD0CkfhuEi2y9FTtvBZz
dPjB7Sj/lBc2irWO18dkiE4xUF5jrSyw4EogzgnOsq0NWXOjMgzwubsTYmoC+X0x
mmoNTITnYc2k8uVJI4YvIc/IJBwszGLJREWJ6d+YbQzX9t5rgxGJl8KTNsQCAaaV
tyHP1p/nBdftN8uOFmFMCVWa45umuiQNWlhg9aTkNSoSPaZoP42N3jluFHf+/FHE
rGDGG/pCjVwapb+QO7P3gbkWxasxNiEBD9oPyeKFLedTGY3SM8olmiU4laSLwujh
Jd+KOfK9vQF1lBrG6dws6G7ZGEcY9tc9+JZVmAo/BZb3E8deRo2Jp9+eXaVy0JEG
eAKf+uSi0sebh199j3laRTyJtXkepMuoMwngxAMlbgDAzxIK+SSZuB9vVnWlhsm6
pqSR1qy9xksAXESRLsAFChVGMRRdhuimj9iahAYyLuQ+iKue8Zj6cqcxUJp93Zma
jOKExK4Y/vc/z2DvbMN7FUF8iOlaXCsS7+nBDvlQcd8EeiMFX5VgF+qu2FpOTjJH
Fg069fmiUD1XjC7DP6t40nBNYpSkVbtv1FrJ+jLfDs5nOk4ztJBiMF/gXFANx/Zw
sGD2s4AJnpjyWjghYUMo5Xu62OO7JL2kZryatq9xKQVO0z7Z1BKlJMzTqj201Hjn
Z6vleNNNPmo3ipVcdB0ZbPXZZw4ShQZxVnr1bHy4UKgtI8m8BgLc7ncGToy67eY0
pkyB+bFo5fZC4nocnu5KURBdQfrptLBSTxz9g4TaH3dioHU1/NatUvDMriJB5wMw
UchPoyb/0dDF6E1B3ad20eG0V+HaRRX/PPBta/iZMBIS+BHRyC2Q4RYbnJCYlJrT
r7E7VjmbkYqA1tNNy3Cd5qIOiZc/3EE4NXsLhr+jv0SLM838Pj6LoRXZGqmPLh0e
t/tjl5AXKcvyak6vLA6Ya6vIsnvcpmLxwFjuZyiElWST4A3cWKOpRPkwrshMyNRu
8tYu3ApT9lWF5xfCD9oMmLEY7E58jra17egvMWjXn2H9+OnMybCwBbLllKqyb73v
t0U8AQKrzX+aJdC1S9vM5vKpDZAAyVw9MJfrDQpnnk9GYQ2S4ssAy/4+vlHBwqnP
wQy6ht8u8fVB/zd/HaTLFMOimrWKf7R+8g/Tq8APw17C8FwCnr4GKCRMAOiGHeb5
2ioa+d9IqN/YVCwXCtWy8r/YdMH5QypyrlSfEcPsTHXbt/9uFUtIXqBL2LO1pwvW
bbGp8mB1eR/btgxq207+vVerDFl/De18Da3jFqHrDBYWWivaz8ZBJGR1rFs/nU78
JfKYiyRz3InThdu6RQh/xz7WtWiLF/j7vjfKwGXydrgSsKDqPeNaAJUnZgyQMkB+
54U3QpGS7pKpvKlE0cHbjXsyBU3qXxBt3gdWe0s17A+MrhIULqgt+mG2pOCl7sxF
LQXtGLyXZGbxPDqqM7Kwp87vrHNLxbQToXeZJ9IqAstpkKKNVEOx8HH5nObko6wT
sZBuPPZDdUPmRWAP19YSpN/5wYVAkbODxV2BUgQO0T4GlmIT0p3klW4XzJGe9V1D
rL2PTer0GNB1NYsaHmghnfDF6nmLGRJB7ArN33TZBXpIvB5CQle9qu25K5M3Ih51
tF6ARJn737bDsePZTq0+iXXS2BUu+Hq4HQZLrScuDiUeDgRyEtrKVOQBcua03tzZ
EdlVshmLgg5G3YVBw3NU6grwEvJc+M2Ynfdl2YJ+fT7jAGYRJG6ODO/WlkwYVaEy
Twb628MH/FlKy7VAx8OqmpVFyZIi+XJblLtULUX8DqeyUKL+ZLAhAbWJCNmUp+9N
jQpZggOYhOg03iGJsKIQfmMjhIfBuKgh/OdrEemxh2z87hjRv60TZXdJcANreLAc
LIeON8N3PYbdycx7i3VEYiZ4GxKRHOQbpYWFR4TPQlcIYKmwgU3EGsgNskLRs85n
sfCXrgRV6stV8pe0A3LBu9PFUIPSXmBi0vtUibwxZbkz8u9edTdU4HrUJw05Oz34
8PY68m9bRgAJZwpqnU7tv9d6cCUOk+Ns8/RXitGctY3CIDu5rvfmYCwYenDf7S5v
ufRBVURS/hP0VZJUzgwsA43D94PwRxR+/JkFoMtPMWQz70H4T6PMpMz12e98Rhgw
QlnCCh4BkrxYEkheQ9+TUzmqOoYuaaOaRtuVQ0/hTbxYAT2G54sHYA59GAgEjmuR
CZfoEByWREkpluP7ohS+iY60GqDC43dZA/v70FAiIJ2S9/B/zrKOAeSR+oKzJUrE
fvpDQInH9P9OQgYIMjkhHlICShSnMBavxZMtLn+q6AWlLksLV0VXOQrRaA3Nhl9m
JV4xfjAREdYEAz3QW7eregdZzNC5e8zRTt/WuQ4gCQ8PyFPBA0sGkyx+/0USiJy7
p+iMGmZm6bOXQZyJOqJ8c4blKrRlxcCV5ufNvjNdnAlytLpkcB2Um+szQ/fF62fe
Ng+0+UPeHVb2JC/bcsmUdwxTWYKd5+Io4VF9cBWyTFql1ilLodMs8RK+Aqu9Ozdo
X+5H03OGh+YZhmZc8T6r6+xYRWKy4JL9JwITY2ILHg8OPFoJDPLc2raSZCFz7OSi
yLGCREhG0NDIyeG7dcP+0UjZ9ZF2NbmNNFsK/SBF8TFbmq84EPVTamT9NtMaNdVv
2VSU2h8KUdMLN6JdWrwEAVLsv+qcykfXsH5/ekuBbaKsHvlVcxiRR7bRGWpd98mr
lTGo9o9E9VWoD6cPi9xc8NNd0VZ5Xvmw/dHQuirmMf3rkm41di+IyXKT7+x+KLSm
pEg+M3n+pLmLW0tIkLjRv+jEjsScuVq3norned3yYGTdvOd7OkK5D9TvaT+AdajO
rEy6rgzSpnXdgl+LJsHlfbOpzSKljXDOzbQr9XgoRp16gQeoBw1zxue3Nd9A3Idg
IUzL1/H3dKTdV/kBDWiemVfKkK440nG74ZtAAflDem7ql1XT+OyavIeZJhrhmbFG
yJ76AwXVpA7MjYq22sObYh6zHuBa6FBqKncD2fSYwqmZts8ru51VhzrrBUbnaNC9
WmgIrvbXKMxzy1uFOR/jzCusXIYEM3rS6UKJ22nqhVcnlV6M/3RyHyCxlLKX5dVX
4D0sGna6TCgYAzqOjNKmMH9gieqyYsSxN36jhqe4QSsoRVLsSwWekHnG0atNIRw5
U22F7gbvH/FTD8dlgj3IV/9II9qBHRU7cmU4J2CL0q8XHHkQSKX++5efNlVa4lVw
mqPcuqH8JFbQQh0FAjtqX9gZppBMFMsEDIlV3ja+de2DmWdADkPQWAOcUFJ/JIMk
EZIiuNhDjCcBBThzq6xRYu3izfhNygjAYL/8hfESVRfYRHniAMrlHO+AfYsaFxgC
Nxq5B+Gf0JPLyMeWVCJ5OaTKPY0FwRE8RU1mXiq85f7HKX7d3COdMJaVmYszEI0K
H4RsNI2P2EGZaTGI6t0az78ivDB9bpMc6/whkNJKFtfQQBG+IlHZ6gQEsEnj9xCd
5Aa+EG44EnosZBAbO8ZNEgYnMF8Zl4SVaSbg/0XUiJLJKbxEkLxohi9zx0A/qRNj
eR3erXuZ7cUigq4PpK6zDe31ZIqbHiWRrlPUpBB7DpcsQek+9YE5MNnEwh5tdoab
G32ixBThEJ2VI61pJ4cIDTT02+PiSQCEP7mXkqNtvA645JXxoD7iwrFvX1uU+J+w
3pFjVm1sNYuH0WmTZE7NCef0C+Yp7N2MonxHBKkLqFtAxhWNc+GUlpmKTlEbIV9f
ALlY0vXhSv0oJaIWksSL4IB0d6mpXma9T4dG2QMMQaE9IY2AWpqi4v2SPICICOyr
Gt2H52NRtX7AqYPcj0Cgaj19D+wluDBp/tuhZ/P+jYX2iBsdXWXzs6iGo7rQ+Rhn
ynzncwxyAb/111iafoJ9HdwIsBoRBIq2JH9zAteH+GI/4Hkuw/RKNms7NoV1Bs9M
gjSTYkC3nc90JZTGCOxHYqQmFfmaGkuoUTB+qE9myaURXMV1n9SbFPI2X2pWFfgv
tklaHQZ/Z3VMxVrbhdshbDu5ADBc2+XPcOghHEkUL24SbEdIVxIDuyuxTLw4gtB7
IBuauCi3LylHJRnG0Cv7SyfOuaqpxI0M1xI48gY++dAW9iBNTc2W81MyDhdsdDJ0
SySyY7swJmOFWK08Kyc4XoUPx0yjeAcJ79lLk3VB7VysVUHvC6HYvWU3PZsUFWb1
6tIzyYwCSPlfzpFQlcUsVEORK6ALZ+KPkDnBdWmENI/xk6VopvZO+DCJvJEZP4zR
0Abv/VNgLuHWwjXEGaJy7v/NLwPMew7reB0l1NIVOCzTGIawLcL2SxMQzHlBwvCn
cMl419WsQJjQBG44zYBpea9K8ubK7lf4ywhATDxcFPmY7Hq70wrU0ikNv0s3cA4u
62XFZkpH/YWQkqGC5GPpZVB/MAfkslyhnQmNmns1i8pjknpb7gMP0uLvZQW2aULx
MhIBY+IZANiz287w2gGbNO+LwB9LFPEEVc6hkC8x3hggQIRseayqex1+tNmO5uEx
gXvrnvSvJJ1d8QFicuYNqcF3BpaHJ2Car9hNKvELnMcEIpkFoWWxhq/Uu4JFfvuA
Ikzvpr7erwq2l0Jckw3mCb4dCsgfJ6pV1b52yqXlU836/zIFpi49cpUzHhV/Ntb0
L0P8QZvGzKztHcafAAGjxZ+vDyOlpDa/dd5U1AD92D2SGQ90x2UmaglGZfJXjxbu
09uJM01TfRXLrkatc7nxJz8pH/xE5EveS6CdPdqBv3EBuhu4flVK0jf33jSlQV0Z
y5IXbZbPM4H8SkzjMN70wuUQOJ0zIoPtllBdlGLwNwWQx7kFfySMeyybqTw/oeD6
GBRZ0OjGXHaQ8y5BWDaxNCVCJIQys3GAyKCXR592gA0Upx/Bqa/FCc2Hhk0BBrv/
lDarNs5hQ+TQ9hWpXb/6i4exjZVTm7IPSR/x857VbPYrLZ72vspTRga3PaSO8Wa3
rWESwRTVLX2ZFxUr1ESbjosoI06IMJRCxIVzGgmMbl47/UQH84BTqE4KhXYz3Evk
Cvg3K3t6BoNFlOlhP1fc0J1jeCqZe3cRwAKcCNwaaqXZfs7NpFWfHocJLlbDfUb0
6LVtlEsgVhXQxG8FFpsLPm9VaKr/aub1pE4xau/wYX0W3QrVXpwA+SDkE7Cl7cK/
Kgb1/pCjZ9C81SzhjNbQvQWbzrXPRdKipIlvfag/zyG9BSBLtLT9Q3Q1pkhQBVkW
mqEOv1pFC5HUwNtm2TNHuj3hkx4AyO9BQkukrUz12pCLOB58mJQnfKNqU7oTzoRc
MKCb/Rnc8vRax3lc90qzDoa0GvdgIAC1gRf6/AD2Pf3FxLt3GO2qpuX5xZf2knBo
cz7AcncpKRrz9h2uSaf2Biwcvfoy+mPdpjiis1TB56NOoao4kMyt1nG4AJ92ulwD
u6C5DK6zfV190c2NScQZhfi3Ip7FEILccDPjkYTa/CwuxESet5XQ2KP6CxKyxcaE
hP/DZFuQUBnHCIXYy9EyRGbfs98wOrydbGESO7v6cf6tMQPebzE1wDxVYoTcOOUF
q6/BNXeovXK94KvKfyzBsGiAR00l17luzJKfibBGft1u8fvLR5wPifAvTGMSwR31
lZXXRf+plb/KxbiA4kvCgRFwOPVoyCO3VgXOJ/tGJQPIt81qUITuYHajhF4uxl7b
gs4zRtaeA0DejwtQQ+f7DhgxnLAKks9WftOOUL02c1Mi4vlWjNSRorKUwSj+zrKq
JUAoT+1KmKpk4TNZKmKkUUWYZvE2JniPyxmE8Tuq9G/kVFh617M5EcLgsFQMz+DJ
EsDnjjPyC2yKIUOruylnTe+1qMcJXS4XuVa1G6hdXqhGB88O2x2teUUx6o5q8Dbo
Y+khIajqmsD93iwN/xYB+EA/fZA2uQUoqU0YJzyS8/nky1rs5Gg7v6lmUkzWbkSN
W8zUTLEPGZzj21JwaNDBcf0wrK9E/yh51XARGfE86lSljlBuRTIfEqCOSVO3xTCm
ZdA9ML1Of+JVkehupDuQLYRGEyjsfYIJO/kLZjsppl9yd1j6BkZLot22/diCfoO8
Wrs9eINjK7cXOgPT5lac4P5df0avI7R1fsAdR/Ad92+M1nbPnKJeoRT624dNM/JO
Y8aPITFyQa7alrbc7bc4DbvY2+WX05MBevS0RnlR3NMPRQwSFBJZ5dNaJ+wXChVj
Vi514EFcZrWIVl3TnIjk0L92vCQYP9jEO7aUtTK0cw9GtgZ7ULm784Gp8mLMNnZ2
aoBJI4GFPR/Ch0+m4sKw3g1JQA1w0Azo4ciGcOoAaeHaDRjyPhSWdsamYNkp74pe
tvq0DLisEQadPX34BRbIYfMHmGVam1ONrmEA8V3+jbNOsDGK4lx9sj5ew8GTcZJp
+l1R8jkJsF1ltUuq/ZH/Dq61wKWDwANSjHWrq8obiCA+Y/HiUJ847rUAbEdOCUyQ
1pL4RlQmwUYiw4I+239y+D6jEM1YLEICdcwtBxHePuNXuFzFvaIZpAIcjXeueMbc
3+DpEgbKeznl0QFzdmOU568L7FO5DwyzQ/gtjsfz1XieHXTP6gagmZqjQCjMaQde
NLfqciYW3/4TuveWPDy5nS5AVIlhaov0CtDYAoHE5iacDqiJJPVuQTWPEEzmmMls
P8RcCw/Op6UlV+mgHw28dgdpgqSRINOIH7dIb/kxNDJvt/NlFk6cwYEmXLxbGNkD
PQJ6eO0cCTdsTYiTLOErOcylXFM1keA5P0bH5mgiQHNSn0AyJKU3yA7HveRTyBMJ
9ULqKlgjFtft/ZjtX7cc0T6BUZjHo416PRQ+2s7L8DIeRKefjoQpMhmYs/zQ43M7
iOk0VJxQP/bJ5UO9BEpwqAL3ZjQXFMa0Fh9ULpoNq9Kd1LaRnUPljYh+9GwTxjGP
PqalrNbTZo5jvYj35lwpb6RLbwj80xpjSsyYFx+dT13sTkDj42BztFPG6lWESHpR
W7gLTajIAaiOr+SZL46INDCRKIDjijfPMYXYHnTdcWOQ1yvmxrq9/8RsRBV1L4XP
ICUvYJ0sEVe8kCGTwni2RstWg4OmVLdc9IHIRRHXHYODEe3dxDIlvANF0RxXKvha
6USCjDRrPufAbkuuxN92Wuri/XxRSX+n01uw3zRHr8Uo+XRXl3Ub9EwbWpDQt43/
figPuysLpMNCRzX89Sog/1kHryDfDEvymBckWp/E1kHZLm1uFfNajzgIMuKztfhi
S1avtEVQFBBohWfavAKdHlXCDlw+zQMxd52jJ0u6LMFaPGwUkLhKtpqoKL8Yv2zB
6pg9eXpnTajNpJIwka1WPXgBrMISg6b5GAjQhqsJyZpVsS0od4SOYqx+chbLCeUu
3e9MfAYe70E981C2hSzvmMioKGwnwiiteWogrfo/yNP9KorWQgfkKiVkv02bve8h
CgcJ0h9GaIVia6dAXa8f4l2pUM1chXf7mWzr69CSiYP8CIgCjelO4VeLiCgw7GEb
/eWxRcPDrh2ANSrCtMuMUsXv+sUnDD+0afQBmPRPk2yh/+002/U0W9yxCgG+jIxS
79OIAonK0eDFWBpdLhsfJnKBfa8n22hF7iNkPstHg2XvQ6dq+cinKlIhu1FB9umT
YrVXGy+rnCTQ9HcSTZ3TY8/jwaj7vAQ33+hA13PWeEdkNnTSE8d35FTcIND9ZAO5
YuPcPdjVGe1Dt9LSzIx84QhVe91wedYtgtVEdR+pHbWOuNbHi0BMAaxcbTvufBGQ
iwTStWJH+7bukPotIzyFeOvKLCJu1auq19ltJFD0RdAYk01n/LKL4jBFT+CHSUVm
wVwHEFo6ek+AxIO7CAaJnJGLRcABaD1AIMhU2SP6qxcz3BBsZngztNlVJbFsf8RT
eDBlQxJxNUxP4oJsyuFk4cKWo9McQ7hlGt+OZQWxFjelKGVzshesHJ7QXPvA4NSD
/IHgxGbyj6L1MOaRGWSJ1eYv1EnWOh8/Vxer76oJmVGS46qKr9sZbSu4oPkHMQq0
osrLwjnCE4g5jYefaETOG9mDtMxJhkhUyCcOHf2mcwvIkj5Vyp/7yrCEZCJyyAoh
2Wyl++U0yyCDbEhrG5+oOwDVHBV1DENVJ5numJ0szekDXHH4ogzU2xwjT0VwAnoC
HQ/lOQ3Kpf8fjoqahNK8Y+ub1B/W8FCdgctBNfVMXwBInGVXXhnj6oKRCzWn0kuy
o8dhrDVyFhOihVxDUsETM140aZwUris0WFnvRwQ+3mUc3LgUZU9kt4Cn2gDIc3tQ
VmTDUPTHUc+jxJmQxjU8KZu+vc85FDKy2hcLlMOFR53QGgzKgJJ/mWmwZDDYYUHJ
I17aA2FF/+MtxLyYu4XnC/DrGex+QCCr8IMh06wYavCzk1VmFjicsZZP/j0IkoXY
wpXA5+P7H631ZXh+fW4is13FYPJ/R1rx90D+/dte6AfVTE4ILeILrD0OC2MG8V/I
3fgXbRlf9a79ZI8XUSj9haTeMsysqoGZBXB4Q0LWC+JA9Znhe+MY3nYxyM/QHtsc
MVTWvlLIRYrlhSjQthvkkqixc0VURlpNpLNqHiZXT5xLTKPH2lISoOI44/jbXZ3x
gNNehCALIgKT3okQfWj8g9qZm1r0V1uaKpj5z3Wu1aoC9ORUZxm9YS1ehCxSXTnG
HjkGXUtIYVVgrNvsFjZaHVr90RoQ4Hw9UHMm+lGI3k98Td9Rufzi/4NlmDU9au2a
wUvYa9347OmR3a9EL3eR7IintD1L0cBjEggiIPPejyk3lFwIyO+WUtXFm8BEAA6O
IFMaeuFb+/KcopRZxvHQhbbwsl1vWnGKMcv1KTav7rKteH039YDLRJGevSD90r0F
J/Cx0qeXihBI+BPDLHwqhdaSTD0NxRDH1cnEooy3fdP4TQ638CsopqRzU3IbS1Ew
assHl5nfFDlpJGt7gqEyKO1o+rDrIXxH6IqibMFJwxvi8G0AV8Nbe1K9XOGBNRb9
S1AOWORxkOtZMXraqdDtmLVhkLb3accnxWUB+XARMkMi787vk6oMtjpb1ssXcIfE
5oqhLmMifel9FjlynWoOEVWjQy68fNcqcUrGIX3SrWwLk8163T0+nWRzEAUy90G8
QIevu8BPfN6OKk+FaLD/7vXRwgRFJ2fqi/WgwS+F8UUW6Y7jCDAK3c7idI/YxysI
qo03an8h1BPGqQQK2+u0eW+GghH/6xKNhs+frRXNUvyVWIiVn2G+Aackyk3r1G3U
srGM8Hrsi03XJUlpzs7f0F3UcEU5Rk9XQrkIl9CPzQeujmAvtaf6CoEauNMRqf1K
iTVlNI1ViFc3kZBPXRVF0pOC2ZzNptI8goDCpT2MJQfMZExvCA0Xu6XannWCALxI
mbtix9yPhfSb2Etws8pSAdZA8gBfE6mtkviUylaCq1ic3uG6gJ+PdbHpYRQu+1if
1lmYsVGOKpnmjzMitvfBUtnTW2lnu3SCnPnxTQEv8THm+msj0uZqqKuRDwXxiZOa
RhlrwZ+adud6+1bN/9Iq85iOS3LTTxoN9zVkIcnq2rD4b8mq03lUeCHCBgRLIhCy
eZB4K6BidhVAFcXd26woxHNMWbSq3RgSq/1SGGJ9PcVLc6eolH5T+VfeRIRSpW/v
ACkmjyV5G4JuvE6MWmutv8aG/YbPKeHQZ5KOw/F9Z5fUX5cllUde87H4N7/Ec5SD
ddD5uwnFuDolTDGFRNLmo2i6hJhV5lIxgQnMR+CLZ7oOYBfapBgiU/gYM1ao1YFL
cbTDw0e1QOcOkkbm7NUMfqhG0UoPzamCBqySllrvPDOd4Rq72bPzbMcKSbX2AOzz
LxmzsQyQCmHbF4hp7jAL9cdJpD/GU6y4J/5iCB/NhyI7rpLaMiQjnHFcrxGizWgA
mWByj+B2U//HKUwtYp8QTuEyV9bvJRofuNmBZSHMLHzhW/WcmF5QONn5MTFSabe7
9Zh/PM4rm+oSx6L3oXaG/ia2LTMg7n1TRY0b2HJ2uxgldg1giOJy89+3e46r9OPy
/vdD9LmQUGGrvDtGiNJKmKHbXeGONjdxe/e+mehjUW+U9Kbo5tYrGL9jN1/t1K3Y
+SCPMQR2VbBQrIvrE0fJJDWxlET4nwMzrJZACW0saIFi4FxIqnA183HA7fYWIiOG
3PE0dEzw6x7y83br3M2fCRbvNCtsemuL+A7zeKHO8CQLdXsOnFHkoraqRb0OA885
YFO8JiO/26WJNbgUhLrFIBsq8Y4EUbmxw+QGFUIHyR+0d0W1IDM7k//MI4StfR0G
EDVkpZavlrn7d2L5JRaA6M4xkhAB/u0ADY/sbB/fHzjts8B7US19t5QCj0y3UCwu
fCtTywwuC0LM/k1y7clZb3tMscIF2lZTTUb7YtgkkmWGq+sSY6Cvla7xsVGRa+eK
PJ3Wvg4ZENuwRR37vQ5ilAZKtx4WUfi+0FeeNKGIbaz+vkCU59vfRmpu/iXMrgr/
swEdtSRTBVgcC+E4WzQ1ITPUEumtfPz8DI/2CD8OfKP4GS16L33P6misJtycK+tk
Azf9aFLqKr1EykOB73FGqv+IH7XpcRfJ/SsTd7JEjnC+hULwGc5yioeQ3Yx7y24o
QHlX3bzRA73xa7PVS8o7B/rKT73/KN+eTViENeBrKEy/3Ic1x9hPvtRJlMK2658I
DA8e+EdZxP6wUfVbSOMfl75wuRj4BBCZbuHiDOe37ZG/D6so0figeuquKxtvZrpI
C4jZHycDuo5fL/VwwClpY7rEq8T6qTvXr8+Lqw/2wbkUSc0A25iY97T1vQtPt/wr
HEJiSj1xQnoarAzNowOPZvYblk9+PFpYUoZy8WOAuurdfsXQoE10BGdAWDCZYAHr
aUul1nyolKNXv0J6ksCHcWSzbF+l2Q+AWdQmlLAGRzQ9PIfLOjY8PYHeEnkzVWjC
dt1HEtPEmu50+XEbNqzOmvDG+8n0ve5R2b2hGJ9y2/x2tTtLxK3O9k2vFJsS9ON0
iIbgEQbVRaGmmsJju8lMdRGfUBlGQK2K97raEYCZ0aBemThXYOs7Qw0uDam98FuW
KgPP/No+vidGKt2K1chFXbWubI3eVOjYFY/sudmoZNn2OsLkawUQiHAY+JbtgIMI
KVUdO7uWFqyma7zGi8rCwgto/JWmdJU9fXM1XvRL/0s0NpLIjHNMOK7b0tRTHz93
AoWvEMVtmGfwmO8K1gveKCvne8rggqYCoxoafGpRMMIb/m+MfdtIjF6xFY/CFrWy
x4aQw3onAGSBmWaSDn3k6+PnWMPV/ZQlyikWz/GT7NeYm7RMmPrME0FV2BstxvwL
u8GhdoPsrXS7U3uKCAvaqrsrPVOIz2qM3qBgKthR14h1Pf4IKgC/RutHhBG8XtXy
wdEJIfkpwYZQh/124eQvinfjMIMoA6WaAfVAy0HXUsU8s3PLVTS/g01lELyyPu7K
7N8vj79E9SKBUTTuEiVJ9GZEApdYabUfYvS55+8Nr1VPHmaqGCHl51M554RNVw/A
sosqzlNErsbjzioNatPFFgUlU6eQ8wNgndxx29mhS21jSajNJ6C/EJFiFJ9Mzs8a
xtLnCBJ5j3APHFmRWbuOyK/NBHiVioip6S7Poi+eg7hj132qg+yQrJgg6mN9lXc0
4B+6hC5P4QxdVwjnQGTuerfd34IkH1YTYHqwkzqOmpDk6vi8ch3vawh9rKZpJmCg
pLHtv+3Vz8z6yhjlQ250JJkjmBfd1qpuLuzjHWBr5q/BnYKsJY1idPwasO8a/BU5
kQezpWqqyDkCHAGlRdSiVsSVO7rYuNjJmg3GG9B2gYgqCjRMtEP4A9Q5B7pL8WiO
w3QGSGfK8RJazqTEHmq5Pzm95E6tm1JkQm3v/2p1lFkQaZPBQIt9+7NcZbwwsrut
0Te+FoeH3iAIbPEz8iynamrsXrGXg+LHHNTBkx7N4w2T9Q5Z56PGcfEvoyWrZ1ss
FyzVC+sEFSUveUmqtRRitPC0AbfK3ji2QUgMwDd8XbQJfBJI+aB8Z4D4DxLSLbZP
E/d+iBtBh6HmCvSUlEjD8ubvJ/8cYBAqWov7xyxzPb9klLcraAEkAPnxv1fp1w9O
g6hmFzAL8umvAcy29LCxp39Xs35XYJE4QsPhYOxxclvYzQzVMtXtpkvMa5AHyCT8
IVaSPLBTCMcEBvcMugpux46LN2A05a6qSbM9/J0x8dzA9OjtZpqCh1RRgL6Y6nMe
Oo3gC8u1mogpoyqyGruWJmb/zfaDoLKZQmFXSfR9LtKAxhZvGUOZaGl3NofikBK8
2uHD/rR6/Dij9y3RA0V7uNUXwyvGJG9uWB1/KCb++C6iDFhBvPqEC+XIkVgPlpTg
2e2TO4EdN49PYJfghNEttlbfp3ol7/Gjs90l0Lv3q6pdZHChJ3PH7mciLsUjnNwb
ZaNaN1Ob+UZASrP2zt+mSMUqfLiWkvjBDQoKRZ8p5nyB8yVqR934aYmqdQ17czA8
ycnhL21mvyxommQ0JFwa3TqWP9T4/7I8dfFsdFThc/7rZ6NriwgbyViDvRqw3soe
LngufmkZEfIVj5q0ro/iH9Z5PK8Am4FQQIMhPwXuwYE1VvCsOnlGK7KfE8QfhKpQ
MAUEufuKEuK9GoMd0uvBoq+JHKvBxvHefGnMs5x741U9YRIDbMSHYIfs5f7jC8FJ
C6UfsFojJU3M7yBacHcaaM5ZqcWp2CjiCUFGLVxaNvUsmqByxyvrB9nuA1E4UrXz
iP2lRMyUeeDY9ZhUFNNVay7VGVDXSBTkUKdx0F4SJPSIHSfToNuDa+dSOe5oT+x2
NOEH3njI0oUHtWmvHuZiK8hgH/YwriDZs7Yzoq/G0C8Qf0M5db2wWsssSZtoS2nf
tGwMQcpzUPMgEL4b6ZSOxq7T1DXCmanq45O/9xQcAqzcbaP2vGrUJ6H+QLIUBCoJ
lT2/inRcHJieMVeGpOjglAGy2+pv6I+q36WK3JKXolYb4N49ouaMvIGSnIS2fyIy
sfdySErQHSYmYEzWKuM+RiFVwMATEm0pytdZDq5a9hmPVlIEXZVRDb96VNlnvoe3
AsIc8VAVSLAHH0u6CO8DxDzRfsyIxU+3GjJNX4Vbd7iIPKfiktR9ULXYXlHEIDJ9
dx3VYNPpLkl0D6i079QKD5zZzrOe7LSpZX91M03J7jvKlgFX2acPXThr9MDts39a
Bq9/TcwgFUW9NWEDzsogf1JN8vXsRd/AtXRGwCAYvNyPPfPbBhVWKSikjdkDrr98
f2nG1CC2a6kPPa4UTy7yNKud5q+NGXHVbAAuVFpXKEtqvz4dZnrUDGHq0Xd+Q2II
7TJl/iih2GJgC1dqsCDH3ZSj8M4pZPzboiOP22fmKpovpabSO7fR4XP3e2OSsdCb
clgCqmx8FC8VoZQF8O1k896rfvrbAi4zzRBFSw+kTdjOGhZMMwN9vrd1HkyeoICd
+K/2h63+mPdVM7/sjrQOdFzIuk2iyzbJJMgUcPhvNb28vjRQ23rR17KpSFZ5FEr7
ddoSyUXts56A/LgLeoVStXLNPWNMa7Hz10L1G9LvgZGgoMzUN3wohANKMH6GmfsO
oH4bgArsyZZgd1u2miEI3U/JAK+xxt06rJbcqVmWbcSMhSuUuFH8HEcbBwiBO0sW
oDIjyMleEduho7V7ZbGcIaOd2LjzoaraWyjFv5MmwDT7xF2C1HA+TKSD5RUHGIAI
8UQBjeSz7ykC6+vJk4v6esvTRK1qILeKz812E8lpXQNla/Uu7k47zhp3P0FQ9cN7
L8aFS1WqzpXNWSFgu0/PIKFCAw3WJiNIUYWNz8Lw1N7379W4LS02KQ4LgLmlazaO
PUfdysE4C9wqDjesHdBAdDwKaAJIXfx+O5XbKAX/Hd2gj9phVRVy8wjSHH/zqOUM
HsOcIiJMRcOUjaq50etRXPGsQgA49c1XhPfzKgcoCRBiUOcVw6i1QK2r37rxze6c
V69QOGfj6NHg/l1iEX1Tks19gEfywJLyY075as1hhD+umbyy1j4WuT1ViDi+X3kU
l/+77jYxFIsoTf1wsTN7fc9wN07YmXcYoyPZE3x/wrU+jmCiF9r/NWfWSjVUgXJq
jR8gdUVsdzb0xgi0/m5nmp0VMrDcR9wzT4djfslBgyikENOf6gD37dK0yqTg40As
/2pWQk57MrLp6OWtQMf5AnCOTrz9c7ekUkWwk/+teDQeasXKxi5ySj7k51IIB0ef
pJYyN9slfNOpRDRM63vooqXJT5yJhxLV9qQV7tq6vnUS4WG5vMuwGIpPOaPBhK+B
e/fB0TYK7OAV2LmIDIpRqmG/NMbdNnah+WpvHU86ZKO7qwEcShff7xGKrWrkesPK
dHFUFhnDGeKKJ6NCT0gVOwbVTjExTuaOPxMoMvjyMX3K9363GYkAFw1rlg/JLQEl
1tpeo4QWAGoBem1c1SsAGZqUgRLZx0i2HS66w6X7Z/4jhe++pWq1tMLX1uHTMHKv
s8dpHvQ8N30jK5jBS4o4jJ91iLnka1XwNYYJbwtQPeiDJTFBI/44ToQYMEf9U4xr
R+r6SOYj4+dZm376nfqLJe2kzwM9wtTAFMu7HE7gmf5n+xLT/uFV6derNp3naMBa
zB+gzyrrD+z7Xd3z4nUFxXgHH8QNVVIjsWXDjkCiGNGga8eqJw9MLSbJPIRBaFQv
tQT6LD7O369kv6PrBy4GPifyLgvLidlze4AXP37UpY6t+j/uVQr1kO2eCyK9/qZO
od48DBo4z07hZb7v8Pft4/Q9qCz8qnkQMxheAyhR9ZNQO9RcDAiyG5VtBpdOnvRj
1udoojbbaL6WbN23QMjADTtZYHNyBphsHb6OWy64lDvcFFtEu5tLNi1zHvuPi83F
NklIvkBOa99vUCBNQmilf9mW6M7/Q8+R0Wx0nAM59QEayFotUalPADCePxGvglwC
ir/9AlCeG3If8UstH57imcXC83pdPsC+ai/tAbsgA4EsVNxhs3vi8HXYxeOurZAE
qnIsEPVkS/o2B13cdqL/PQw+9HWjMivrbyExO5FY6My9+QCLm/CTh0MVks2rnmGR
y3P9vZSCXr1OEAeF5ysymEYn9YiqIcIN+dsFXa0PZiVrV+W9sJPreda7tajKAr4e
tJG6s5lfhoRrb0k9NZOlpJ/0CkhHeobXJ4tcmEkdlXkb5H1Gtg7d6QENihWj0Z7c
JXc3jsEZwH2Uh1w6dbNgs5tJIXns50IeBjQ9gpHv0OHtwIH0SKBg8wB29a5QsAxg
i0CcjeH0X4shUcYKQz6NnKRCM/AD7HjHOi+nzdQQ3Ng27zCSDaQPha9v7uJWWDBY
R1PzbMHvq7Y7m8rXrfNdIRZxq6keRuUZg30hFrJhZYi78R/GHkNApn13Ml6oCn84
xe8y+OjXFeltFqgtP7YybmDhzPmzl7vzP6t5TbwVSebnpxSJolY3tbNkVKkyRhwl
Axht+3nVJem92W3craKDrh4QHtZmh1YFPJm408zv3RAI8RdjkOZYtuVuxrcOfLeu
hrWEJN2Aqvzj85WP8keGaJjGKPeks+e56S5EchVaZMOOyF/LnGnx/kF0QWGEWe6n
Oo61ccLB27YYexELaP+lcSCNFTIz3Vb7z29R1Yxw6qSBphxyfAnHuT9MKaim0elz
I9cKF3Rzr1PbSVTk0GCuI033YbUuTZffDVZJNbG0pUcoiIqE6uItEyB+n9exfGBM
PobPgj0mtzI3B4SYmGx1vZgKUzEWH0RRqDuqjcqL1hTkLlnM7w3JMxuLUim+6soB
Sz8kSjU0y+NkHIkKcvvbDpdVwIORt+77jgYii1keAh3pfW0IDxHlvKr921akvnNo
pTVrkHH40AtmQZeA+3GoSg3ZbImddwkXxpJZbtwmjEj4eOm5UZoYbii6/qk9Y5/+
we1vi8rbfZIsXyKcgun9diZIzchZtYMQOHftx7dPpuXpYqUBhTXuR3DldWLOX3wX
mDD9Y5osveuMQeiA2xZKlSc5uxIhrxXa3PkaP6/fW09m9O6UzuPEj4CahIa8r2uo
kil/+J+yjDKlRB22iW4rKinh9pscd+pc38SsPF4AKbZZl/fs0j+tXHbZag7rCfOS
xOlX3AMIEF/tSaPzxt1GWYl2Zn7D46fS+MGhVChQerBFYbgwoITfjuv/FU+DFKp6
spxHE99IfG+37Cu5Uh5x5+hPA0JmHvDakllzFNTPfPp0ffJeSm4MJYtm+Jbcb4Ff
T2aJksjNKtZ6ohzRKqZb68ohiGQeF3VcMIoemoJGR+ntjyTWeMBFCPMfXyF3JHKb
F67cTYBrCIBXDfhJtcvMcdTc8koTNFieBMBWbRsnYjRFp//QkPWHZymOwza0y1qX
jHkOC03gGZ+/pvfBG8Jf2O9OZREBFxbqLAK1UjknXDDbM/O4eShULnr2EXUIgCEG
0zVnnMnxW3sKsBuu27JRmcJ7ge7DrptwNya8YaJSbHzDr42o+b6bdmOnwYsIyk4K
aLC5kZVh1eYeV/nfGphjqmSW3thBbg6gN4P34JpZ2b2j0DkJ3rnv6v8LH3Y1B7MR
lt4UQPMNks/HqdGs1gLNkEDxVi4egloVZZ28Pv4MJcsIFdL5JjMV56cPtKJYHJav
NQ3NlB4ta23aVOwmz+hmzNq0TNE+qW0i6rKNGGXm8d7FbcHKa/LYo3NATYw4J9ll
gLSGVYRiyZnuSTlyZykUvDDHtaIGplPtnkH3l6tddryHaHEAXRJYDzfAziT7U8ZT
leTMwyUFU0nWzP9s/UYfsZ/8IeFkHVKT6VsvNKB7dclleEKxGdVp4G7MQa1YIliX
nFE0fS2wZ4rUCWfWYGPXbpSIJE2Py324cW9Bq3ZCWB2g5ixpFZHao66FIiTnofPO
8b0gM6IS0IP2uPKEB3VWyDEDizr6/qkCD/4tJOIbA2NQVTYMsoUFTKJyT1hUsyk4
iqkGnwvN6MQg6coC/k+rbPAqvT19SOOmS+r78E8zGUq0yK5Ay6bAKGoIqLAQl3Xt
0/fk1OpahvWK5Zll9L9OAKgRWtHPJG3+R/mjwXKxzUq8iODIPBUlQCSPiNRcv6b4
litTlopZR0F3wyIkOkgxl8ESuaCLE4Zx5niOL6dBeL78ezt9YT3vBySRlTUo4B6E
vamWW8KRfxPYVDVbHXt1iKuz7D9lInIcW0OqMD+eKrYRLCiK1BUPgtTKBEyElyCZ
oE0YXdxWySz7pAOxoEh0WXKLrS4dEJfBVbPuRyntLvn0jWcSZ9EzTkVARNmgYBhK
XYT7EUMBu8aGf0OHBCtRc+q6PR4Y1cGbIoF8v3Vitvi1vJACKftSnLlOR5Pf7UGx
saecQLfu85BDODE+/+OcPeIQL9/QPGTw0ME59OpDn+CVm1OyqgE0Nnln/cagAXR5
l8+P3Pflb53pRihJIOo9dU85pEOwIfL0s8JvkDw84zmNyVg3tiUx+rufzRaFBSy5
qbhWwpX3xDXfCrtrUweNaogAjO4WlW1OqwqyssF6Bt0tZiuDVl4GgXRcvG89wTcc
XdkSWix7sNq19XzIt4lmDPyOtyYkFRfTLDejjpSQxhYnmOS+S57Ml5mDoAW8AbGh
WNhAOx9dr7yM1b0N9A/vBQIgQ2qsgZOMD2Z7PelVs4564ubD5Y7dA69A59YwcaKC
ejch/HXSPPgt9/NxgKhNJ+mSCGUdyeEqfgkTCbczGYz/DKL9mpRxcgwfFYleif0V
zxmFMfEc4842GsggpN3LR7qen4gFXPYYW6hbNGGVlsXYVNK5n3PK+e3aie3f0Rqe
iz/H2j49trfhzinLjFHzD6LwzJAO9u6FXpD9ZJ53E01EIQBljvJehXAVm2NCBYgV
mO8Hc2wlj1Ox/FHnt9Zm7pZq6Ye3QSu06nuQjmgNUb2jsNNFZS9qf0lxNFLgihDm
guPasDk+AH2xuCUnAaUgTlFe2aToN3a7vxRFsCmXRD2rLiUhH77Lx3hbVlwqzqVI
6Kq4oC/xiWXKPBOZJmiYna3MklOQ0vZVG42ePaz1oPsKFtc5jo9c95KTERturmS5
cotirQ3M9Ed1IrmBhsWUroxhgnaU6u6oMA1KtalzDFQ9wc/cQelrufc1FlUejg1a
tHZ0O+yL7EqebGECjefmGOSKs5VBO3+CqImlyAiKpFNdcKV9JEdzP4fYery8XOcB
fYrq0lzdjQksbWTxCEgDJxXXj6cNYqUm2ytrT1rcqj19mUf1j2GqxvSwai1kw4bn
Cg41Ech4dvgy49g90uKCeBtUkonY41X5NuCLzQBadQpxMWIpAaiJ/RHmY7Nwt2oM
4S5hDMa7N8Jb3Bk9CLyW5hlV1rc9LUJeU8O2hg9lBNBQ2bBjAEFjO9E8MwCmnlMD
tANU6nBxE/O15Va+AwnmwlpVqoFGxStkYjbEBPNlg9Vnb8afKh+Debp3olHFIVw/
d8hvufk84pOcPpeiZVWQCHHquYGuCrwbgM9L+ZTCcr/RcEnNvJcKQpCQaPqII03L
qH4/hJDyfJTLpB2FXGSQPI4DdId82wXo6WNnf3sDv7TR/bbnWrDllK2ewj9NkCNw
k3HYdb2MN96pqwJw76eWApWlQD5fSKajq8ToV3uNvhkh6FcFhZaCRkLtHqpZ2rSG
Gzq5Otxu8JZKs2YZx+CVAS7mhP5BSgnXPILoPIRG+qhNcVL1GVj9tnuzPSKspSDx
Oz6MPEVmPwSgHE0szOr6KrtftHD5/QdyeKr0ZhIkMdo1VI6MO1TVryggELSP2Tbm
nfCz9zcMwFh6LAQnDx1fqEUrAMMzGVBbbR4MLgMQNYKkE/mlhF+2UB39HII1TOyV
NJoRovveAk4GC2nzl8Zx3F/z4+Q3W2/PaQzb5VEEdTcKwJwxCOa+IOlLc/W7v+8K
T4ut+KHI4Bp+unSS9XfFKXFhIB+Iv7EKet9KcR2qSgg0nDqeNCCed1dghBD/T9lu
fedYSRAkh6NmEGMnQgJOejdRMAWcBFKEK9LvQk5Y6F11oeodBbgPPb7fXMmce9/9
Wr1erYazE2PtfW/I0NO6AOk4oLvXpgqmMvw22eP0LdhYNHoTXleuSMX762VXW7ug
BAAthv1IaKrcW71T06Qs8Z+5+1tQD+cQK9yIgtgx1m11YhmIcLHjqAMXknQvM4fU
BQvx74NO8xOCx7AYvxPBqJYVqSkbD5U8mndKVvPJQwF+ZHXpUghtPchJG28aPOuV
URArQqbhZPB7DVRTi8G8SfzaNJ/02Jt1E/Sp4ihV8KKWqZbT86nGVCvvf7PBmh17
zHf6VQ+TF0tY0E+1Q6LC0sFrrh2TlKMH16Z3jNXhRpcuqPMrMHHaZ0RYLerWnoQT
wwqs3WVBGb9Szj99AJMZ8xEqDAjm8BKMAwCgCMQ+LyYoak1QrcTxc920bdCVxF3F
499K8ocigQkTNb+HC1Moaa71j/SeDah5cnw+kDl6wIOIePrCpEZUvlGzp/Yl2H62
NDlIUv79T1y6eRYrnVad93QfocRS3GoUiJ+ABmZGZfa6wE/+9P+3TIQN+3BThl/j
cHquCZ67p/eB9PMBPcvsHpjsMT+CxJH1AJVxjzZAr9Sa7OdJv2ikRjObmYEw6KkF
Uq5LMKj6a77bDYB755NSr14bXQ5rBMGuqTYHeH+//Ywut6EHoS297y34pHLPk73c
QcvJLNeM5C3V+M7DiHX3VuB7PxYlnptV4QCou6rAYaStZ8qxSaM8/vlfzdJnZqP0
B7jR4VD1oSJAApPjVAmf4ZOOCdB4zvsUYuZjk93sYXYwsPlzKbskNvAqbnHNwno9
mz44MlhxioD2sWtE6EKsu/PD/W0/ygFg5a0MXcq9cJZMtr1da9pc/TIWPMSnybvv
UEhpaGg99dphULAQnXuRAylz6vnBreLq0K+Hst3MIVy3HD/erRJu/F3mFq2A0vHP
89WifArhLil20bPQ7oYzpLx/CuSdA74guqaGVAf0kfO0I7m7ZBvgccDYNRugEnij
PycKaQKDOIIx0EeLxa2SDBN8Q3bCdlvqoGkdgi/ukZIAQ++a0/pnOBhT7LvlTesN
02nH+6tso1G+hYwXzuhymgwjGrmCcxqAPvoyfUUIu8TD5HWLyvB6x13iJ+edxrvN
9rJZFqrmmiLUHKjAA9CnRPMumn/ULkw4YojGCBgkLirLpCykysY5gSBHG8/XBdDI
9JAHYAtcrYbhGTFpS9aGKnnxPZlpygYEwDmAlH+kbYog9+tanTJ6OFxKXa+ELLyG
gVFHvgTkx9v6FmSkaCRSHGQCj9XaOufb/SxYk3Ti+cK6yBdeygQiUnLm2gq7Jx3f
+F3yPcDqFh1Q2Y5N74kIyEAxChjlNB+oOKU+Vvrxo1yDkLXp0brwaDStvWHjHl+e
2p4WRYay2f86I0zTWfWvvKZ9/lXo/GXyNo5lu7wrREhytaFCCUpCHPi81fXGjlCz
3pnFiilWjLQj9P9Vrn3Q4nU1jCm5FV4X0I3YEFqhzu2jJ4OPoRmXBzAIdm1LUwyD
Iwj3ZvlxeDmEEiAgTxhj/hdMvUUVrRMo0r2SGK2g/sNJFnJqdMsTz6pEuXOLWzKM
GaneWKtJ5UKIEqx3OhlzvbGAdgPkHRFX/3xncjMTR7isnQQXPaa5GQfxaGCoMlMF
0xNdsB9YaDZO5qWKbbpAb5zsQL1EQTV1oePQGxj1KJxqpJfSiN2fbaR4uWPadP4x
bvTTzlu+pS+7apGMBAmiDs2UxQs8R3sSFzI6zIc426lQptHLKz4x53J5qV7p16DR
tEz4f9srpw/4mkUkaGOpTju0mmymtQCimBbRODPC5aPB9PI0lmDEevs2BQstKDAF
hw44gKOkTRveW9w+VAZldXjOd/944I2hPm+nnJrfjQGfo/uG0RJTAxs+GY4xvYR1
unTTCssR4d0NbWT5P8SOBU+fP1yStdxmbGCTXWLAOTCdUTmemyz+UH9Rx+YgZavl
OhJlISnHlowMJhDHM19iCdoGGBOhOZDMLVLFYbCfSefIo5HMGzPXUqLj12uqxDlN
qUWfjshSCCjQg/P6iXum8QNsCPFl/tZTaR1mdRJ94z47a7qWzITtpFwrn1qNI++Z
qwm1izaYTYsXgb2m8sd0e4EuZdd62FCHyPUXbpaZOHOX6YlwjwhtGPijDvMz5x1O
+4qPIoyatay4Swd4RraiY5V8lP2vic1Z6QKlHMwQAe0KMijM8A/Yxn6EI9O4FxZ8
a9bnxGs2Z1Cr1eyjG+pcoDyqgCnX/pVgizvJewEzDOoh2QV7QYbubUoe+ja7I3Gq
JriLtA7cKw1JM0Ve/z9D0FZB0MBN4fCA/Y1pFitWZIkD6HROzx6vKQnRGno7KbQ8
GCfCFN7ffx72n3N4XQKszlc5uFxuzQ8N3VS7uyDPjPzzZM55YrZJhYEoOGRWQ3yJ
RqebM4R7uUoGvI5dtIZwEg/ufUqrTVs43aB9CS2dH25RkludN8S3S65atPeEimM5
/FaMYqjhWxZVm4CI43uo3fgU6qDfNRdCWVsxEj9L5ZuUsC8qNn1qFOVlC846Lwy8
45qTI2k1CjJR4i1KxyclUJrJmiGVzAgE+tIthvShexzOLYopKBpgvHxcvGwIC8gq
M0YbGal6beqqqyrGFiAHAU66gh9S/I8YOlNQXWUSeeCgXo+Q3dNk56G2ITCL8l8V
pfB0qBeIxAGleHk2XJnPEWZ33geazRtj/mgFkBGZ/omOQfzhgDx+gKtO2Bj4bYej
050cqcE+cwIQ84JPNt39z0iyy/6/fkCBkK9KFGus/ObeGGPdE5BJX50cx7nBoMUd
Wxkw5VhJ7ixQTDMwaRhmOVlRlpNia0L0MFYUGn6XiBLDaRtJmyCgPJ7M/Ozdd/Lu
bxCX+Z3X1DsZHaHUsbVHBkujKsvBscrDOHqf209n7y64K5BMqkOYkf+P6xSALIrh
G2AFc/tKHeaPUFoMXGvKVZ8NJCO1v+/IHRSwGMTM4afWgU2Nld1W20gqxloXfmE3
MTd3TsZrKm1poLHA/vBCy7tbJ2yy/ZqiSJn6QpnkNs/L8zmusC9cDXaxXthGxvne
3zGl5U1CCz0PQOGJ1iQjqp5OJWFZ++fHK7YJK5Q14S85qJLppxQax4avUU9fC13K
BLgozgxkRPVMPdqXf7Y9J8UNh1ISBsHo5GyBNyWXmp5rmbGtvTqBt94soKu6JmlL
jnz2xg1XYrXmJFDI6a4yjL082sDj4/BYtFQ54f03jHztAZs8/oj0mENtyscQjhBP
huKXp//0rBp+J9EjlBQZYp7BGZyhlfJUz8epqnuQtL/sFEujIBneW83wCg39+dW3
4QO9HNVmYl80wM0530hticBl5iKMUSLgHf5ODpRD6+QI15wz5S0uoY9rLwoKs6iw
C6/nYpoBWbNlYv/K1ONzIXXy+bjg7zmPGXBrVE8jkJQEc5EeV1nfUy+OegaHdBW7
kkxPIKx1MAFeuS1Fx95xJNVjqEZNzEQQlfeQpNek/ALxYrlQWlpB2oMG7N9ypRUY
z6W6hIv3bayue5OteOmwck7eSKCoapA+Y+0LuVlR8gfipbGZVTUaVSkvJlqFuyi3
bAq1b0QZT9H641Vqwnug7nGFrpW0B4a0AmLAkZoIy05zHBajKFZr5n7J7jvyjsnd
Ny2oobVZoUKca6+rJ/yapdtz0x6mkcJwvtcVlHM3ZBFiX3tALzAo/WeRf8vb1meX
zpOHBcNg5l0OtPkcPkUwTkSLN7V+k6ds5jxYnYioXDZq0IdyzI0eZhTtkUQvAxur
fr1lLiGhM40TzlePR7wqHv269NRwnioIDh+sJ6ubpSxEaJW96q4OIURKnY2eCdNI
xkfO0PhAWW9CmpDqYS1pmLDpW73XKOP0OaTj+893+B4W9UfjtjXxxL2i5RbIzhmn
xjl6tdFywa9x2cFokvlRV+MRYAwli2N2jMXJpC21/qjgt2YUJZ4IVVQPTNd4k+gf
Ku/Q4ZBTk6lFUNW/RgVU1c6/qFQHo5RHQf0a87ihwnhIKmFWfzR71QxDQ3J9AWkx
z13Ex4es6Y3TZ0/4qLhHhVWnSB7mD3pXu2v8ciX8CvPwKsC5KMXR96CkpAIG8OsR
B/82HiDieBJ0MdCUnDyd+Sva5mvrWDkg9TFgLOXeM7kf22M1oy6n1GTESxinBpgi
/oINi9t4lUR7BN2u6f9PNlCbPPD3P9t/dbPERRQuJgAlp2Qba6NjfjPWUdwLsuA6
8L49S3RBOcy/3x+82TSHkh6TM+SI2m4xL5cCXvyagXCIWRWjAa6Bls0NQ/0XSTNm
3nWVVxDDndqYz/mvYJuN9n/lSXOoEDgIE/m67qw64Ryt8tt4Wo9x6AWyFoYfkVb+
vUPIdIOfnfPI4pcL5w7hx+o73aEY425YjRzDLixQrTnJWQSb8aRoJjItrjnRnv5+
ccQzfkFKKRKu0AX4uSXteKWt08S9yMPWx2zxKwTnpg9dVhLYWwK2Du4e/HFEegNg
QiOgmOZiCG6gOiT/gouFVYs86dQvhILLesDhKBrwD4Ug3Z8i3in9+eiht3a7yp+A
ekQY8hxBI+JLEDMgFUUZiQ8gLh6VO2paP/Qa7jcJvs7BJlbSA7/0BoiKPuv9uZWT
hBvobFmTpV0Nv2h5fhlUGtvNJVO/XNuB6Qyf/ekPmfJIiRXgXhSW/L47uDZfTBfI
LGiDroAWemIPWGeeJrWKe5JBpLBNJEIsijmX93D72Ke5/giNcHNCKAMI5utIVDka
yH8/MBZeaq3dQd8btrDNxAbR+DXAxG6WZ0r/ZAvCZamFoCVsw/Oaaq/cdyfPcj/o
cgvCdSVMmElcbLVjlMvbkQOB5gvDBDNOPbJ1liHb7nNXDICR5Ld7UDDI36ZcrR0N
tItmeUmE/AwzrKU8cyoJWR9y+UFdX+1QwN7tI/C50MsUeb5EqRXAUBt75+XyDrsH
6okNy8YPnuCPq84mTmPtl9W4QzC7vhO+/yq14WEG5BFP0giQt0nkkKZDbM5UCQgD
qw8/Rze9hQrJjloUnBiQhy8ioCL2HqY2SWzexoUlIPYIMcJexzTvRwd2A0UPe6MQ
x4CqEo9K6Z0sOKZus8MT7EB9wPliH7VcH1IWGXSV9XxhFFhyvuPaqm3tZtSQknIV
Wnn5s7oKpiK7nBMnXiEcRFQiSQ/1wwvxSFe8+ltrkQXq48nitRuCsauEEi7uOBhl
lf0QkCaVRzDtLZOnrcJUOnO85Bx25b2JS1x9ZSYDZokHs6yFdHpKiS3fTqAYFLyk
xRmHi63brVAs7uShSLoY+ibEATalCgperO38bo5s9owmCcTWscMwlIP3f5NVuIMv
x2LRQMU5kS2lrRwzp5SWi6XgjNvrYEFf6fBhwH/EyK9oPN1wdeHnJ2zfYOrd6cwa
+zMK5Pbe7U4U4CGv/YFBsyfKJleJmAVc6mFXeAlnagmVXynF91M3AYpXfPFWaWSc
GfsN6LpjPaNS6vtBHViv0/xM8NwjRnNXl1yvrJcGJ/6pYJMd6mO6kWxkYPLUhGUE
6cuSEZr7bLTPcJOIoNMZbg8sXoLQViLLdGxFCftfF8E8G3+124zmA5ocmByKfbzg
8Y1jnOPAopQtDRDkmz+Udyb9iq0EZfnjYRjZBbEdxPTXbPKGc5GR+TN6YKpXu3iz
PLZFAzTU1skcmUNcIPvIL828Td6hsiTVtynKfV35K0aEBmV5bF+yFQlZpXrjtTfm
5s2JlAv1TPjgA2KXWJALRLCru6rrLpTV2fxeBk1hcg/NjR1QPVLLegroS1iyh7BE
63gzeciyNMDgFSd+iPQKcc7RQI4ngVfzbgmj2U1pZCmN3r3lVUE3EC+hIcBD3cg4
Eg3fT4mTOU6NpF1F+8WxKK5v1g4I5BJijQoWzUPwf684u1HMD/ErsKaVTBxiOwQo
5x5WzBp74VFbMhYNQax8c8Ywptzs3zHonlfuXlZTXgbL4FD99tNwXSu6SE2kuIbt
8k/sderJ4Z3ZUtC197Ke2GFzVcI4zL1l5g/3a38PVuBQ9T/JdeJre/aajM3UcKT5
BzsiF77np3nxrt854cKjs/ti0dLKrmBhqDMeVo046/OiQApSute7IxW1HX9+oNMu
z2beo0ODcpJF7ogIasfuZ78kL/yZ6YAU4yk4LWioPDyN5It5Yg11Vnx091zKJYFF
5MiLwrc9jzkVPkbJFSzHFQGcb7um7QBu/xpmVEn9ezRAwHXcLXReKXZ0Cgj6CsR/
06Ctf6G1pQInt4ivXa+P4TRAdVle+yok0aU6brwU51CrKVfttc7kNvNKbSjJBSkP
vlxZInHpu/Jjgau4p4Cs0bdHA/c78HfEjXrycpnoIf+WOrBEo2yhR26vUzXpbWX5
+ZT0PS3fK6vcSdMGfiFq/LfGMvmCZubBhUvt1jrJ9GNBDNZ01nvrT5Qw4v+qsaSg
Mn2fYQ8jH5EQQLovoOXuvA5jxiiu5aQJD9qNBDiDiiEwCt9cYM18jbnS8YPpq3HH
lFqw6uJWyfICMhjVa+eyM76JnLtFK7BQkbapYPvpA6u5tsg+llTyrulfsksI3XsF
x7MrOH8LHU+1hTUEAaqk4FCfj8cuzkF4oo7XOAQ2vql0spYUUz4jP5VzXdAnqBl3
0aLQ+8DE/2bCVWtvyG0PkU5+Gdu2DcRkT53Lq43McLDGN1uskm6QijUzUf3g004e
UFhPTDeY/Y7ZuS3prE+YYA5SDC5///dzd2X194+voHFTpcxQIYoIyWTgvHHWjuTQ
Sk0ixZAXNcLRjysMMCTtNeeE+WBVB54dySUuGqAQPFLU0NssiKjWpfOSKkY7PkIq
aip7OzBzozsuecXZYNVWOVCj0Pc/8S2+zrgUMT8j83J1aiWxYm0OjV7qid+N6HfB
BnHJpnBWHLC0cHpbhLyN33KdUgmJzAihcUStLP4Q67RLPQjNfnhiaCS/fgL71Hwa
GsujBT4+61z6A1dbKF4ESWddI5PsWovOTEqY7wwwrUFCMtvjOu0V7v7hze7A7uFA
x6nLuDXWcbJgGl96P+qmWqlD4uQ5JnPCGQeODPlfegMAl+LL9Msk3I5AM+QdNMQf
qeJtC7DXtpwagNAiE0RVWehQq7oq6R+DoTc+oQsOfDEEOZpJveRrQLfOVA/4VI3g
YyNKh7jNhkgeRKBaqOlKme0iPywgXkzmmtttSmPE1gPgiO3ARBHWFN5intOBeU9t
nPoLHh17mx7mQoHpIN9F2ZtmBZcLmPhPxN5m8hOSXCecouBuMK/TCqmO1431s7sI
c4c9hyndysSmrjfzNpMkQJb/Jf+9wN5vhCjd0TQaNWK8IvFuOpt7vCh6aVWZ6ar9
I5qkh7O2AsQmLS9JvtECBpnV+I971RtFDQ4Mlg3exrNaC0rvYG8aUM72tCu5qp/v
qImSJHgrMleIEE4i4gHYC2pGVxdIqLAtQ82KKIJFUeACq+Nuk6fU3nz5w4Odtjwl
NtoPMsWq0cdGfG5drc3z8NDwZ8fPEEW+UkDQBYmyokHcQfXlPTOzjMsuk3IrIzMo
3LV825I3FndRKT3JVIfBv66erp1PYGJbzvP9h7VzsJb8cHuf4Bpf/0TXTT9iYoQm
4rAwSNyznuGIshBh9lve9vQYuiFpuWsKwvoJ0wzkPoZQwmwtgIJpjNsNRrOD/Ncn
mRKaRIR9n65Z3VAbX1moFbVme9YrPkMBiDH2WmvM45s2GZqLJosFCAK03Is2qiKF
YxR4vftOr4o0YQaKidkc6tt2s/TkQ9y0bHwyOHoGARueIiyduBD8Ng3I4BeVaHfc
KsKbsu17OcGLd/rAoJQBNvYrwCe/OnBokdEd0JqE4vEX8a21c9/Uk3XVearhtu5k
27ulK5HpFHDLPJhtFrT9T3Y3BoLJE+H/qYzygkFIjLmF4vaM3A+JyhBJbAPNQ8Q0
+SFLEO5UWBvWrE4uqQexVQ1Up+ocd5B3h+7TxKRuzjXruf7HHdLjREkM9hDBzpJK
Iih4ynadxIWqP9mT3RFWOG21E5SaLhEqISrk37KASIHb65VMuLv/NV+gF9adl/B7
TS969fw4VPOjboTPWO5s38TrgT5BVMIT/gWInjoPTNq+4RgHUIh+vB+jaQj1o+YV
90P19+BmY1kQGomUjWz+VLvFV2OhMTnJCMi7zgp38QExQrLGl0GwrAMwerMuoO92
OdMsAnK2/EGv3ZNsQkSi/9A1Of7eSXyyebww+bvUOErDzEB+1PoJTvnS0OKzjq5L
myhRG06inA6tV1o5A3YLweYMK+/EgcI/dkFJbUItTn5no1nWfQHBhPwFfyjrKANP
+MLSFQz2dC1Mu3iA8gF6M1wBALvTuUmFCoYh2qEVt6hwVXVxQEdmE6z6ZFStW+my
GSRtkJuWLDYZOjs2bxRMClAuTi7EzwvJaJfdauA+bxn+o9unExkJ5cYnqZGy4yIN
SOzWwXNr8qIWH/JoKXAGRR4n1YuAb4XkSLgotAXZooSSKknJRm+I1bbsia5GIyB+
s/fTPBySKIl1gnEO8maX5wCZxk9S/kkcMOOb7PiqZR7HQixRlJKLWrgdUqJxi471
atFnLDO6d2k+/9YSqmVxwfgjD+A3eOaVaK4kl+N75ZGyzgbFfTueWlBOaTagyiO+
/o3LebEz/iu/IyJeD2swHlJk2qfHTfqlb8pn3jh/iTbzjwHk4C2K1mn2//pomRks
Wskn5hoPNUaE/+nNlTpMArlkwSEMEwkfhPjVp4BYaq0+npPX2Fm5rgK6v2mn6R3i
Bo8urJ6LmCVeG/3GLIEk91ChPzcfTAfejsk/yJ2c1rSEuw5rQfcPj+GxsTSGCYOw
Fmh7zSSh/NXJyR2AvJkg9gHuGG9Dy5E1+W01seS19eIBFGtCsRrpbidL5psPkmMh
rft1uOFMtbWYNY2ZxMzTGzf3jGmH7VkpugZCyu5wSt2zcrom0xyZYEV19xjy8z8e
xdgEv+Skqhmv20ED7eRvs8i749J5kBLVVPM5DHP6/4v3rohXxIwJ/c6amvtSUSGp
Sb5JBj3XJ8ZrVFaQVVdtzprOvXVXDn8ZqhztDBHwknV8UaDv4eRJC3sAKMN/t9yR
nICa9J1BIvQr6nrSOgyWOxJWjoi/lKFezQYfM0YKdOa/YVKyTIwiSKrngsOQUq8M
IfoZSlYd3s5YF/jQvgPinwxI+6WD7dfdJ0hO5emTGgDeCFXUTZZCUSrZoS6Q8fS2
iBeirxgBDKeqrBeTw17o5iXHyXawz1Pc7PSKZERdzhAd1jAtSksDB/9XglfrARvI
anrJO1+lU8CRayn7EzI8pX0+R0aBLqoXlnlS6qhwXOnufc4121s19qR76XOFfeMv
OJ6q9UiWjm9+7T5HREYj3yUqOj8Wki80R8gbg4l56baU//7YOFrcxmKC5SCmyXyD
ysh6Qkg3+vObS6rb8jw14NeEmSsUlrLSetZ7yo6d1mXmmQTOEfKpgBhhdKv9qMMo
w6BT3Npw4adwsXI7mgs99r+I8ZUPC18trJuS1hkAB5n1+oc9piQumQoKAUXBUpQN
P+bisBULmYf3XbVxFxzOFuxnLD3ERxv+jX5I+wHoDSiqZTwBRaZsZpzROH++kBFy
4FYODDzoEVNxMC1o5fCfimLLsgbLWpFk66Z8ALtud7O6wyRLf+Mm8XZ0B/u7Maw+
yTFmTUgCs3Y1BCaniTEOBOLAT/0bV5fUj7mh6NaL9+xhiv7TK9CNvTgj+r2ex9Ou
OD5IXNOUrHZzyX9PavEKRfV7qgmpw/7N+NfWjtGHH8W5X2LBMEXrdh0DrH83lCOX
ZgPmCwusF1tYpTfdBQP/uDzjxzzREdaLaYJD1HFGRKOZqnyEbkK2P2CHcJhieR8c
C4wdR7nG+Yo5W44BlNJXY63EOZRkCs6L7iXelgdkLMxyZNny81GGxbIR7mb9+bea
Imk4AAz9paVRWHdwUv4fAm7MTeCVQXIbsBqLMwAqJO4+bbwo4/j9TF5Mg5LGN16m
3sV78ca+iSTyfdJrV7q5J4H8rCucIyYusYpUnToLquBw0RdnaEqm34rFx6yTkxJF
2DGNTltLOt/oVX/cSkno2Isi8BGFC2GbjSZGGoI8Dpd5Yo91mQyE7ropNhzCFExb
kz5Yl7dP2zMLxvVFqdeQEcmNUxSoJ2K2dPoK0SeetI/8NxQVB6cRevlViMVnZ6RH
RG1uK4nBrWyYgLJFFWWiH8ZtLxpV/d7SILN15ZD90zFNaDOslOib/yNFQ3znqRwF
yGWZr0yWYRRyW4mwQkLexd0zW2h7BXo+eXpkSZ7XNrhCktDpaf4mwhwItFq7N8Fs
2oPBUyrQCiFgD6farS26LicY1zU+8lYXu5tMARDQmTXsbukdl/SGXZgQLlfuZE4H
GJUnHjK1ARJkIc6psYpHfWcCWHYzs/RLbyeGP6mk5TrNnVKKfnJf4PLroSkgRMZi
Jl+OxcU1cs9mQ/1g/eHYbXiMnqUyuKL71fvTZICIly49FsWa1E4LQzcvsv9emY5+
9DOHtl6d7skNPQ0GrMaII1Fc/l7iOcmmsMK0xjYpZQonlKmFMu0sNnTIlC3WzWuB
PftP0g0Qy1/WiOFqMwGlrDiRmb1faVtNwhmDF0RZKaT1e/5qPsLxefXLKLx+UasL
sotTiZvCtz60HM8768Ui/eCij9x6LUpnAlD7mjkvAx5TMl2BT74VdzoOjS/hYMry
HM+x1BotRKFauww1s1fuJf8OXhA9xodCCD7PyFz4cq+3Ln9/4Z3A1/IJ4AzFAlKy
jNrOH5M8uq0jvYQBJSdH9MfherlGF1KBNkIdeoI+sH3RyXQfkr0W3kQ0S/Py682n
jjjgbwX7oqkqNOqDmnq+gxmwGMDNU9z2hUEsKHsxRFztLwlpR64oYw//+77TOoFR
bzqrsFvxPyb7jaPjjkcHGMxVek8C6VRNgO+EFArTKpyn8eDT7gwUZqq2ZBnQ7TFP
gSH4oqxV0tUf5VR515whvo3fzpBA3o1uPIxsIlNsgzjAM/TRZDZMEktzsLZRJASt
X421RtoppY+mGA4QaFe6ywnb8RkoFMr/HBWsFoUImhNN1zz8NuNY7nxkvCd+rliu
kLLqR2clXb+VdzIt69KbptMZCGmOHeo4MYIPQhCUXG5IRf2u8zev0SaQTExY6zQh
bScpG8dhAKzJZGdLaow5kCN7EnMsgi1kPgt1cGCo37FHgGu7jAIpGQ/+nw/cd+yt
7OaUG73UR1K4QZIEKpOiUyo8hh/ZOu38+S5lt4oK8Li2tojtb2wv9+/zGJUFr18R
UC8EASzK2CpV1qphxAkfpEmaQCwrKZQXsfaf5jJJylfSnKL7D/YyHc58y9oWtYrj
xJ6N5EPNnkPZCisoBNZnsPeFzTyIH5mUijDxGxSrDyER0oIsKJKnNO9LzdAeOALl
5nLNbBg+f14Iv/W6T+EBqvyhZSGnfVyCB2mA+zWL944ZGFfEvZ6rZmtEZKAAjjSU
f4m9OdIPs1X6kMu+9ecQGj1BVoPkBnY+b2ovBngAALN2Zwr8rVk2isnBK2ieftIj
nzxU2iS+MEJydddZP7GL3yutdfpi+YbG6sUIFR4tH64kMw1B9VnUeshnmVaPrW/I
Fh0Y+UGxJZAdPELP0JBhhSGCJnR50ZTaT5WJjyN7eJUQTWbzWzbAGM2WjsOqlqTZ
y8wLVJRmbwV/cSlyP+leQHQ8EYrcyGvRIy8jYun0+M7VrQwfGm+YXK5lWRwOaxC1
BOBlc22lJPhxMVLtJJYYbuaI1z/ymzgv+YJPADpxxmvEz5ZUnIBJaHdjam5zF1LL
cVCuJBPd9or5qUcd+mW6BYldrpC9ghlfX4tVpnz3F+w3VvEBaBWn6kyDCI8XnpIw
loUjMEQs+0x3WRou2PPIIy+Z6hmiKhniVCJAgBfC/BSH2Vqi3MvhKzm3Fj7jwkKA
dxWgUQMRqdfPZ82cMI8GUtlpbLRbrDHpmyXVBauL7uDqy9J2RIccZJzKsg3OKaME
1IaXR3Sz01eciint1nOSNMkt3oXzMqs5mCs8Pdb0lt6JLffl9Hr2hVbEVIuAEK9D
XhVVHdWo/ODXPkanBBtJ6pv34uCI4DnEHOfLJZ0EfW8FHqko2cKHx/RfMc9wpXQ6
5QH5gXIs3aTskcg5LfWwDK/xFt2N9s3MgiHT/3o2flYMwBY1F9e8vwlWTjB9+wxT
UraQN0vdfNvtN9xl3U42jvUix68fd4ONtCsP/h+X4ijITXALWb+7Qh0A/atXOt9H
RmdEqQSrSCj8ssjFcKkWoiKPAjrSYERHs9kq+IsZIeIwsa+0wpwE/+hokNXboKV/
4ZG6BmMMVCbYXy6b/wSQXm4+/4+oUXnTxmD8s0kb54hS657YAEhOm12U1+0/TKZ5
qKueFcMigORXyyGLfiG7hIeatQn6OLYv+YpVYjej840vTPDk/UVxkP5//Lj0Z98n
fZi8uv0vr90KVMzUHpTQnJdqsrcDaKslyVYELnSVmhcHdFHWdzoQpTaTw7B6o55T
FA5cj1Uu3VN/9W2wCEDYKGcnXo28hOKpSLQPp9ssDBovznUAewUnqZJSDhuSLKeD
sNj/oYwDm2ZcaTYl6orv8/bvA7h62S+onUAOWj4QYAvRrvUKELUTiMbkMxOayAfE
6PGP04Pqqx+Kao0KaAWmcez318eH1gousePXN2GAR9frpQDGLqaNziFGLvjA2BFf
leo2c0vOT8n51ULzKrgtpFgZGngHQd+CPwd6iy6oG6CeQqLeiwWwdIlXW+5uOUhg
qPtOf/KRgbt3EllMPye2M6J/BD9/DRvQrtp452IMegxxXEybLww90uoUF0LopEj9
KTYfIpYF6CdczqjgO+c/02hYEFUg/+wgN/1S+0C1d2qB9/bBoIcOfzmBtQEpzk3I
SLHmNvmOsUJeWYhWQ67BrhDpDlOT2Oii8xF+xREDnXY+k5O6mrbuyDRuYjWPBd+V
MwZsbcvtEwgfL4J1XTSrCWgVlCXbtFVwKa01bu46Uxgel4mPWoyyKQ4dPSMeYXTm
hAGHEXNoatQRfwZdPpwBMJJ/veT4Rj2JXSd0sNu4Wtc0ak7043/mWYWgevSaoaNV
A9AhJj59627LIb378CZ2hKp13e+4ja03Qu91OWZGPGTUuy0FfnSr+yJtpiohqbdl
3/99+/dvXwKXd2VnK3MVujTnFEKKS1MEHH3mpM12ZEWAfShUqQ5IQsKmnakqONca
NcZMXAB/PwtzIcBWiG2sKg6ChiCVnbtav8qAYW2zYjeYxcI468H6IRbCMrSDNktE
rajZMGBCAD6sj8tn16iKk2jBXLaHGmepfpJ+8PNifnMBMydEuAOkV5bxn7hOqJOY
h01OHV6Y1xwd/ATRioxv9desRy6U15v7oD6HZ3np488zOLLYa324KCVDOs1Du63w
NU8snRQuLKXC/OT8/ZNwxtFtOWW02t92h9U8WJWMEeRIqVEydVSE9jEBjvX3E8gP
YU2slv/scvZ8Q96sabTOINrNPwO3xLPQP9egpB5EDTJA+Bh1OI40GWRXppP9zOTt
bHbhEoX+Ivn1x3c04kx+kn2rAZRXOZA+ZfYGKonXJ+VYWzwVrXw8w7p+ZaSjXeXv
yQQohITZQUeDF3XsnvJFq+NINZlRtED8Tu7iN1al4vqjeTBlX+4tBFIwkKvVaAxz
+DjZwyJYOaP6FSbB19bY4FQiYeBNkDRV5G7xmueNYFBHdNGlJ+LcmvXhz7Amozs8
+NzJLlcRp6d9rzhM4ThYqzWvl/FrJwJOiKfED5J3AyMkdNBUATQRAklMCxPLdCY+
qn33aRGVE/n3iueokHOx4RxsOjA6DyJnGxAqIqzDOpKKXEWPLTUNaALyTg7JcPy0
AbkXF9yasnmhMjpCAIL9wKRdB7wZ6tPRffBHvGah2AxOTeZznDYzNacp8FcHwzVq
9M054htgv2XoEE/U3esW0l8FVZTQpn0HSu/Umf9x/OQ2hiK7LkyyNLV3Y8MttCDq
iGcu5+n0wPQYAN1yOxN9ILd/2XRgl+ki9yPt0PnMwORb4FrI6k2jgmzopLkP/iJw
eS6WaXgdJBBjOgwV5ToqfaZypXaSM82r90KHuY3sT2vFEIsAvkuNWmY8jVlQWe2n
eilyGj1PPYeci8z1wfdP8/Xj6Yzn1Ggh5lH00v5XoZdoDBQAQ3lnXWweC189h44g
XbDQsKxZbylODp7nelE4pAu6puK9bgDY9QLb542vYFsYWkLzmSgj65ciicsR8cvp
Jxwxnq3tgmYo7fefvnWgqtG2bTXoh6a8myMIrG0J+zrTojBgwpKWpWE7BYNsKVhf
UsPB0cI2a66GZu2ieICKlu1XwVLmAq9mySq+108xXP5lTWAsrWwXvh7kaQA3FvQq
bNeeFlOWixI6K6NVXu3uxd2+vfeIRSNZQyOnvJKO8PG1FGyl57NNQ5BtvTVl3iFQ
lPhaF7kkJvBD8BDKPOs1ugzKPiWtMVc+krgaoK3s90smPyX3UgySEiH+qYwtzEn6
d2ZUmW8Bloqx/edBO0hnBD/zNuit8MKksYhxKqOd2Ex/Y91++Gwbtd0fGw5hNYId
RmIPjxKJySOq89i8K4HwUkdKnAje4orhgl+aUm1JkxjcMt/O4SK0vaLvP1ztibU3
zcg4VYfZDKTBpgK7asLy3P+pQoXu5zyDxIrc108cd/Wy58B+oyozzo3a1iS95fvC
0JuPJKQ69SsRqFCSeeMgu3MS87QrBwhbq2n+RqvrXT8lElFtbcxHf26tdebAMKBY
+jbgvtEDpmHEpLkgz00cjMPt7E8Yw9nSk73zXkR64Kdw4zUs9HC1A5UOk1BUhQnk
OLrwoOu6hAT5oSi5BnplcZ6XSf5ocM6aM3v49aR4XmOY3yxVEBJlVlK8rIdsynHe
sCQz7UiVQMQjmyegGi+hbdlBqBfExklZ4lEK2Iykh3n9qqKBCadgY9/JDcK5YOEi
v/l9Y/IuvryevomvKdM8mCc1zgfLiOS2H/6Z6rG1c7xoNA6uEEsp9wv3ZV3BCp0t
OfiyKcES1XJ6uHVSgt++m5VMcHRL43YgGdtCs6KVk0tedTlRp7/ESIf/dPqqOVQm
+imKUs6kGoWk1MEaH0GzuvbX77LvaSVIoWmp3g7mENgNp1fxOBb5skWrwm615rou
pUSQ0BwaJjQ6pMxvOKTeTpnJPwx04V0/ez4JvqQATlwNFQuep+tV5xF/P59Bdqib
xNAqAqTf3DVgJBuB8/6SlY6Qk0QXxReaX21fNREfXcOKAHC3KA2bDls62H3l3fOS
9hEaateIpgzOxL0yqA2UQLk6LjPdHcv0eOJ9IkDA8nx+tIck8ay968ebFK25qMyn
ng3AGzfg6c2wpTzj6ayTcvA1dNcHSXExLfaKb8TguP6Dms6982F2CjV/SZ4ZRsD3
xv4Ci/MPz1IXdUcVnhpf5aQimJnWLsYk/Vi1NGY3RKfAzdnvb2/KZqc3x2a1rmdb
OyxU8/1uL8SyvLVqd0409acT7KsEp8k4eZt6PAyNJ0hjfn3321xJwuNTQJUr6jzV
2bw1HhmGDugqLi9ZgEqQ4tJy5Yb9Ku3rGFnFpGSn2mGYKfeVC8iN5jasrTdz1QOO
JcGDORxRS38hEqkCps3Pmglvu/OM75W7Hh+424BqO7Om35rGhbOvoeh7Tj/VU935
STGhNo8G2BdXNowlhGsMQVTwTqdkzBupMSEmxqE6ZpWTqWWZgwMrhDAjORnxPH8e
6Y/jc49Ug9syTvJEEy2uyymBi00wupWBG2ar7hzZKanwP5i3jeqBdWQ29Bfv6LLZ
`protect end_protected