`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36368 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
9GNfeu2LhBO1rvG6TqMSwGFB7dhj3neA4P4KFvUBgsKAs4NWIdD+wRwX5rjT3Eyu
beyrO+B4kpsSz8kFkVVkiiaruAqjrZhTzjbaeQaeFLbRuNdzK1SDIxo0luKA0giP
Dz/KSt1epSR72zuYvYHXnOzgBMXSq9MAlHfSpI6bcGEPMkqqaUanPtwHS3rthJ3F
E44LTDxA0+2vZe6TVcIxYZNR6nRL7rj8XK7l1tI3NpW+Tkzq56EEb/hz72KXmvaT
29hRgglXxxu/JsEsGeURVftHvj/H230s5/m/6jfirRmakmQVVP3dAGJFaXTLUr+s
ZX0S8uD8iZlPXcxvgMT2eupozL+jXlXtijaMw3s6BYpH58HgNd780HfkvU6xM8/p
J7AAabCPeGckxLZVD6/wjn+wsKRRuQLUDFDLzkh8PVRA79h2ExVJB5P1Fs97aVT+
uwjF62XBE1fD7RuDJPL3nqP8ICYtejuuBnkCB693IPp8ahO6Ynt/Yj/3SBYfgrY/
zPb3GYiw519lWcB/IKmZTSkrPfFkyw/xx0rMBUVOcZ8Ic5SYA2Sg01jb2K5KTOCK
iwum4JCUV1hK7GvoSkyALrMih5ABo5XDF0oF8X8MBU15iI/pncbqp3SpdUGlLYjd
DgitKsXIWtU9yVe6kSaLU8bfk2ivxnYaBQNodGSwcKezOkIf80WtUAd8MZjujsvx
YisfmLQKkVLx79eqVUr3DJNVuT5c8K3RrPTl/srIx/tTGZ6az8y6IJiQo41FaPE3
MFo1k11tB7xfwKPsBKh7yvMXq2s7enftxymW01Huc17fC3fvDVTC4tDbO08UQPZu
rQg3M6Gj3kpsGqtKj515DpXrUi6O+QXs6auJNLqp1TZvOnCgUtQTvcPlp5fNBUzg
GYgH/tShpMdNJKYaMOIjUiS2F00fQonj8dH+6kTZ6OgGjvGizf/DMOEwvuBJibLv
lADtFWDLnS087UsaFq2DDEE80XaxU9aXO4BSk1fQjnYoGprDwqvdm3T/8mZtwmTY
1A0ykML4UZcIvntyekwDJJMZMrLZEvQyc3R1/+Gu5IOsMMKjdmxZvTJFkCqKI+cj
4wbdxmIibtgRWJe/vMHmUMpYv/3WQOOzMEiq/mwdMtBma5onhxfbt0Ey025o6OQz
dKVl02d0/EOpE6xU1JhVZ7uwXFLRUsQHtAWNPA7wuCm1xm6SeuPD4ZYMd12Onv3Y
pvT98GTulun22r9/QNR4gzX8knukNwPLw0axs7Sl+1vtqJVzLkA+qkSONl2XXO2w
lHA28+dt1sDOojQRx24SL1Z8Ayv4dj6b7jyTIVdiRi7cxPbGPiPI1yOgQJhXhaMK
a7RYSR9PHQXlc+InQ77/QqYWYfSLXrZO2pbA5EaitBIAyEHcRTFZA0Ts7TBuZ/o6
DmKsdrnvIYk5cFaAWPaEzFUAxC/zkKWcArlyX+6O6lLkj8/KQb49dR6qlxqsuM2K
AiyT1+xWzbj6qz3Gf3S4x1FtQnXHh+J4WdWTdWHu8Lx3p+Eg0jIolmfPEVbLjgO4
d7z5gYqyBwhc7oy9ICDRX96mWVm5qk1OU8z5CI92wecELxO3txu+9838Ri+6L9Vi
bfCsdmshYwfhSlOJyFrOpkOWsYRl9wBZXa8vdjUZchz+mVeLlUWlavN9TgtNi+7P
OCUZtxHQP9ycROzn66MspUg9CQbl2bnahoRCUuBLuuQY4bLBsd/FZeFnbA2MbN0C
1AISFDExsHFLwS9xjRQfXAF3BfV7a9KClmpPUX6qPEb4rhbzgTQzUJPz3gfsvlpC
WHboKqvo4bIV+Zz1WT9equb2bH/YbXDFHPdzJW+QyjxmMdbf7HdcD+Yq+4s67J3X
w7BGvAY+O7vBnChuXoEqv641g5+4I/LKKw4f6pyv/1/H48oL8kSW7prRjvpfGITW
S3fdZpncWulS1WiXIMBmSZ0AOadWkaYJHYXCd24vGRhPIwt+HX0oyLHXwoMZjWiH
AzI6gEJHOp9z6ej/iROb4+ZLpd3bOLjNgp/esp8x6wsaTsTFgh7F2s28YIW8SELy
92lkY0mpxiT5mn59VHNzSC92Vk+fRplnn1DJrVbixoV1Onn0JsEdr2UBRwsNE84z
bmWpSYU/HnAxkM0rV42Ii6XK3ywgklVLwOk0PESGhMrvtD9bmNwhMSo/V6KMgJlD
KgN4D2hjvexOr5oa6/yJaduigcaFitUlMZ1+Eia2Uph5d8x4bCNalq+t0U+siq7B
wIWgycJbOvdCfcioZDodwHN9HMpLl0zylficTdN2lDeBcio6Jp10foJ3WEoOcm72
VGG2rxj4caHnPvBW27ho8QfUmhttqvrXLgc5u0B6T+Yl+leAx3PDxjPhD1ixG941
pgueUuJjHxz5x1/XXx3IccBCvyOEoPWY15Mnt8Z5rKrqXfLsgpLimAWgTh/tSrNO
JR+GjF0xtkyLx+Ryn1CSEV5NjEHKQEj8SnZppj8GTHmwI+YnaL6fVt+xxfgS6daY
QJJOG9FbOInfC6FD2N+tz4rqKYe6g8QB2MgZUM3vnsTpDvdTb/yHWeB3c6WTVu0K
YUJmoFdb67FdkoCrLdbgUPwfFildxnk2DyzmZuOF2O0Yatn6vRre/Go75OaKoiFM
L7n8H7oklnNa281fvQaO1W4lJU8ulep3sdKTGaI7GFXEdfLzLRYtu+SWvMqFyalD
WCj88E/c4DMZyXbA9DDn/UHOt5VbIFbY9b8iZdTswir8CeColsUoE0ojk2YuWlF5
TmF4npzzEO7le25ejQNvnqLkvJLkgTQS/vRbQGxP6S7TpGhVIKcrw9U3yLTMfllW
VRcN9Iug09cPO9zAsL2vrngwpEqhRxI+pdKxuBzlOwsIXgLIQj0UU6ZFd6OysD+P
kmzlaeUNus4Aht3otJCFNdQKvfZSq600mx/99XUSfU3is48O9rkLvNufgsmpdKHL
d3X+WzzIFVbewiPqogs7wXBCCnG9Zr2Vi28733bMO1qNhjbWxNGOE835ojxufOSd
nxifCVufW1jDWurw1jf8SkAWGLtHGdJgdoZA96XlLThv+OqCWLH+xP+lc+Ybps/d
pf8uHwY/rUoddzkJA/1yddt3Eev9tcIB+ubwzDVpd63cjQD3932odP4x/uzfj0S6
2MgwD2QoZ/CYuKq/9n8aemiHiJ5wTllXE99gP09ynxhUrFjI1oyWi1wOaIkxrTbm
muxPSiMWWkJr/F2TFXF50elotJacoz2m1ffCxzXeh84+JGlCqcBIbiXgmVE1rOGW
sXhSu67ieymgsemvXSicQjLOlXHm/FwWrDeTv0wc5fq0T7aPi3eZKXbOHtS3Ay1v
CGv1p+RqiVR5JQ0lctNVpf+U+QgPvwduErRx9tfM/fdsnuCOhNN48+bhjlRyHGnj
ClFNKIrYi2FnUGNpikBczG4NKp4Jd2LdjOe3IzO0jBss/uA7uFWtSExIiMsyWCbz
+Z+kvnkBBEv2a0c/4434C+df2Jzd3UbMPlSqkw6KtXn8GiV4GrDGNmuWZL/CadZi
0EXc7B/IjsQTsInbBDsSqU0cFbpYabqYEHkljACrhhuCgBvWj9HZq4onGY6P0YWe
GeAt6B4SuuTw29CV1OQ69S2fdktzADOzOvVlPVUlOMqI2JBeg6+zqAbjv9/gXnYF
agZ7Q53G6utEXaSDhsfcHURpQ730jgnRwDEOzGONnPPQ/uSxJiTp3O2iWYG9e2pV
B9Hc3CgPEnPDF6RiqhNrvGeGE4rZJiwFwzFv7nui+ar1/OiW/ROVpL1Zey8Y18lz
Yfbir7ddLIzCrKhqUDKDFQfrbkL3w8L4OaSNBldg6HbgWC7EqD/B9fPSnJrdrnWo
ZYNvh3v8VxxAfsINkuh4pyYSATgGOK4mGO18IZYrpXUoIGvaZH3q8GdlrzVZw7o5
6yH8pN9t5XzZPPEvZkWy1j4nZx49yKbPeN523GDoMNiYRpf203bnPOBblEgw3OkG
m4tQPiSeXDzzUome4MQHDfg5wRA73STpbXM/SeZjS3jJTIhBCA5Y4nVBl0JSfaQj
Kk7TcHwG0NRtkkHT2HqdEXKvH0Xbqkmg8drCskUrUPPQ4dokRmB14sDqegi0Dd+b
QAkMSjGOMQhiQ49+qh/E7K4eBCUqACsJTb4ENmBHv/3dB0DxDB4/yQwsSen2lRg/
ZWae9wGtZsHhfp1liGUF3LKU5Pgy+pnaJDaAuiqpk54VhiKPKKoP4Ps/M0KMZpIL
jp+aZpYlljhJcV6PLWpxj/PB9dfayfTa0gmRkuUZ4Q9mwgwih8dyOKco6585T5X1
hG2/4wuQqyDPpGNtIjwW+EhwFvkrp5xEBp0h8ZSdqmBJrkm9u5EHBUOFqfNHOd5B
96lRfc+QeP8kppWHTYWDysD04tpmYCRReBlywZ38Jem2Lkp5cBqhVR0MvD8f/3Dd
3RVDxCxLzRaHvHzkNz1gMbRDVk+WwJfwkA2MIso5Agj3SWeMi65xRdfINDqC+g48
pzxaAXfw7XZ2t/r24bbnrcPR1rfHMFod9/JksgncnwIAIhb/XoRkOjvR4W1yYXeg
QF/fu6liVk93koeUcDK3zNWfHmTN6amA5o8uunJos473w0NOtL9yX7SN5eAjrfET
PpYEOxzoHa7pscBhsBPC8bGcAf5ylu7I6JQrW+7xo5ZY6fEnv/SIbQkFYDlINPpD
DWwtoVPMbCDJu9nR8qwdg4i1jqe3zEpfZqjwmyfd13CkiKzAElr3Qn8GeVVRPAZ7
BD8mOzG07R0XJxvTOd5Ko4b/1dePKNfIU6tm6fOWQHNzOGE1g1QYHW2dEDfMd7Aq
257qJUq3kNq1o4TubopDRjfRR6doXwgYWZiRzOYOMz2uGlSCPhprVdqswp2dBSi0
ILhOPDffvD2ElJdHg/0jLFcSV3zr9OVpnO+NZbW9aX2E8WwCG8jyNEggLPLYiSzt
YJUmvXdn1Gz+TOalrNxIYcqUj4et08RR3GdSpn1O7IVeIV0K0KcQsgXMOT4yd38O
n5Pf7IYr0uws2GGRjD3bUT2UqWy5MLVssnmx8m3rjBGhiP77mwOvCtsMjNa4CGNO
G3ZTTpccsMz19k8k2bcJSUkUaD1IVYkCFK1kK56aG1xo20Pf9qIRNeB5aO3dQ3dZ
dpXZdQIU63uxoLGV15K1POI5nOH9/KZOwSJ+GOXyDM6empgoUD0R6osH3c4ibApy
cQ7WJBX8VrbkqdRp1Fv5SYNrrSVUjzSuRNjFsT3f6zLJLw4VnajYKvla3M1Ty7Bq
C33mx+Ld6fv8nJlS4XJoomIRgYEaR5vRQ+4jjjAgr/QDknI0cloJTAPy1z6FejE7
b5skqXRE5MDc0XFVEGGiKndFH4VtsVmV3vYK4GAfgKWiEdHTBMVsYAVZZN4nuiOA
QW+csNrhChaTXV5n5WhNW458DfDvnCObUZ4+qMfmLodY40Fh/JNdx0t+qH3TW2qO
/Rw+x/YsBnuNLsZbwlqe05WEsx8eU55otlv1wdqWXVH49vZDfDjfdBWS57YIGezN
GBMzajgWJ0aInDQwh4JY6Gzj01N3GQKaDUeMXrEMVYjQp6TwvJpq0h0R09IPwzpA
naY1qw/N8eMUnhbDjRyPZtMROl1sL9imjRcwEIUUsAmoyz0x8RvH21g/h60lXlJo
VfUcPOe6zBx4MtLgLwsN4sUm4BfUZajOtgcUJQGe+UzLz4JrDMUkwoWktjFGwqC6
QkQprzUUc5TBTmFchMp6JiSzhxvk7UY+LA7GtHfKr2MgSk0BVMwoEqRkwpQ8CKDb
6ChamLQxjt8kVZLQ+AvzcWpuAXY/Ahv/ZlxV0FI+MUMsV0wZstD0J/a3cP8eqc0U
CEoOwldj4DoNdowmqheITi8lrvcx5btlPCMSO6dRzyDqfq76kVmdGZ9PhOn8nHEa
JVTtwe6ycxC1+QU2neiED0a9ETtRp1N8NGwRpki2shFGiNoOGP3Sk3PADMFS/RUz
sFKpOmVsA4ZC7e7t1yKgLBamgmD+URGXiAph+Wk0Y1gG9Rz/BkXnhEHPLKMj7moO
kULB7scWiUtwn9eJlt17yf776TUaGfzJ7YFAOg35bDaPurCeI/sJqSd9UFhodpFA
vpjv3diuhq2oUNikgRFhs65Si11M6YWl6gCmweb44OVkDJd8UN5Xat1EitftdMxt
Ax9FJ9T54QXDhGJuWL00QRhz08f/ZyUA1IrRECgnyfOEq+cDbkzCXh61P33dfqf/
oe8u3I9b624Gc0kSzOVZapRj1nbMv9GnMMv1hnXECgQFbHWnoVFB2jael7b4b7Q0
4oyfJ6Egae6R3JmTTxh7GcmUk59vDdX01YwxR2NuXINfXGJPvTO92gbdbBLAhwKj
+7U6x9YMX5BvPUySzC9QBtRIAtwHGEsmbNRYe6bm2QKQLJpqn8DlzPWnSANPsdod
3vJCA5F7yRbyto080FyDsnOOqZAr+cHj0wrsmcyYSjUbN7BvnLfh1CjeOYVBaGF3
lq+24ma+RK3H1JNzRGw6LmwBphPMMnpyyfURZVKrGbdvIKXFJJv2PcO/qwv4aiKG
wvdvbsLEMR5VlVPJsYoLRD5rcf0n0S0cDCrJJ4vqPj1FKa8Xn1ptnxcpWzVjZm4U
s24Iul2pB5fj8iX9WRaf3V62igszNt7I1A5epZufZezVzvU4dOXHJkINlXxg2kvY
ktmh1YXhz+aI/OrKv7wKRsWsQOUTYmP2WY6X+qybHtTlavG5+nEoQqAAhyWK9V6p
sklsh0kc8QPQ1sg7PKhdZFnulwWOV5lHD2EG3gDQRBJDokCWK5hM41Zx2j8HiI5c
uKueueAbibfaBLoA/56ytuBE6Oh2Rdvh7onetdF7BavufGiJFpD+DHTSqMFDnHZf
wycw+za1ylYXliP4N0iCR8BfRF91Lp0q0FU+vxBNY5BKX17gDr7iWPv3OHsF23pE
RBQhbbJVipalvVxaLHhHexYFtxtX9NRDpZPHoklBixHpqizzusiHypi9xWMpQEAs
+gg+2qGHZ4kciYgxVCl9wc7q4yL5K3eXel1eLpMOtib6U9CaUmP8g3E+tLMX2wYE
L8Dq/KCcn/aDCrUd4R0RNHEsA4ZgnJAomUiIBtHWNwEotYrBfWiCXk6M/r/jVjN1
fBQDe/P90KFHm5BGZ3wtKTrBI8QMxDuO4ncWPx0Yd3E2OZtRrVzGm0QPGgLpC6l7
nHgZ7Lq4y3b+qqF335MuEROBzsfyVywveT6mpSpCfAyHAgbiS2jg9nOhQP+LtBw8
eA00O9NC4nWxsmiECpGNSWgGgjgnAaFuGe2xK/jpgE4Gr5Kqj/AdZbRWjIurAIi5
UsocaalWAQyT+ht8OmRKjxgqgxgVj8Ywxv+Hcmz1JVW3hJgMgG3cZ7pUWqYW3Bs7
5d7Y1QfZZQUX0CkyUyoUhgIS+bjmF6DgrOHancR2nQ1MyNzeJ9IkJ7gXHOv/M53U
yRUAKJBsiHkq7gl85uE93/I2BZwfmW00GS6mGHNmvF3hK++wtXS6UtVop6DAGXa0
Njfbj+TXzIDZfihc7WlgOd1Iqv1yHeGPE5ES2btEIKPIwg6weG8UuaUaVZ9A2BlM
29eqhhLbNQcQhpjzVz/UEMhNsK5IDMVi+dY4MiRCnDoqfK/KjEAmZy92jxYVsUrs
TT5+QdA/Rck1SzWcaW81sD1iLF9hpfkatI1PE62TSVmOKlqx/YIGVcEZAkGssdI0
VW5Wwf6YZLk1a1Cp4zALEKzpuTzNQWi3qyy/dFIY3NHncb+cPlHA8IxBcNzwNWcr
4i1R3tcyv7cPl55li6XsSLgCpcNyHLHvnSe4zT6KYR8s6Rav2Xz5CTMt/Q5KP+Fw
twyfjrpnJEPnLjKUayHslVyCe/zeMtqLTSsKOlVn64+O4fxq8aCQK3CpH6XhCUiH
WivWv7VORt1RxYQYqd1dUUAZEOGHM316IsDtSwAXe9Sbd5jyIV+trYiCAwQkda8G
oelFwjONaveMP4StgjBmlNUY/8h5XQu8PKuB+iRsix81egLn1DjZW2T+bJtuSKUQ
8qa9jh1CtYRZtD7B4afqTuZ15XbYK97ChBUGyvESaBCquA/NA1+JoTTD9oEuMg6D
q1vZNSKGSKof1xWKX/GfcdputzqaLTtxGXIRMfmU5FqSzueYicMcQTZv524Sz81E
f2UD0DTrAnRN5hPYNFJt/Nd3eXfVB9H7jV1Vz+Rpy7C3WzVMpy2V4ZQEuA5DtCOf
3PL61ULaPAfO0TFVmXeURvlBj8Kt03RMF/qCRIoIjlSxIBC7QaTnfq5cO3GYt3E8
Xfv0JFaUZx2CF3XfirAOVKjPSn/iw1iwe0r+F6V+0mBVOHtYS3ifSM+WaHbDBC/N
MYE3lOZm8w7yd1UiUxf07cwuMSZcZDtUKIAhJ6GQMcPhEdApGjPJy4Bfm3znXJWs
ctFTpTfMAlMSDpovhnnMgD9NadEoeYg4aGNhpWcHLIA3YYL/PpxloTxyWgWqA+i6
z1qdhOlBslsIFed8/SLPsb6ZBfDHe0hl/gvBbE5zSq9FVtcHeDDhayt/fcweCr2Z
vz/WhK3bk3ZALz2ra+RC49A+j9QBrVfgFUbTl+aVtUyZ/JFETVemvN95fP3S+kya
dG6fHn05D7KSIZ/UL8T5PQnC6R9IjvBAFQTt3olHK0JE6awifxGejQ0GWRlsTuEs
ULUzG2tt85qYLmXU3jxPgo9N5k8ALfw/gbVkbNFONB/a28V5XhE5LwjG3PPQoag0
hKEWgxkv3B9JAo/f65Sp3dMioDEvwelbnVF7niGOEf9K/J/97C3a6jg9h53oFn6W
cN0XT8X/tAyi1/HqiXwbKfTH3SBWJ4EBBeEB0j24DpiaLUJHS9yoybdEoarad88u
WNPE++tO8KmDFBEJ4etmuYnIUf64qDuoRENV3otc/8ZtiCpUUn+NT0zplYRG5a04
Vy8xmyNIZuJ06PR3I8hkGSYJQsVwtVuAtWKuhaORcamAzSJnNApoAJiQG8TDI6PN
yKqA3mBIHCKMnkIaH7e9xdRpTs8cFH7BXFIyTFdIdt0N9/A79cgOI880yWWwfB9u
MEeEA+NGK+UkSiTsysIHfGdMQn3nUBGPNQ/JLjXzfO3cOK6qTdHpl66jISgu8mmK
x6KPAAmTrarOMwgGjhgHOmJUsA2NUMpV4FAv/XyNBYzaHUUDSIQ/8qHFNHCQHPGj
2hEklVAvN7IBVH7JptM/Q4qsn2k/PmI+jZgndQPpJrujICvYlIGiJD0jV9po9zwU
cVN58hg0lcFZzW21jSYA0XU61YoUKZGDD5SvRgMV2FElGfnBKhc2Lm0VX2+yJPNX
dOqITHl2Yil0yVw3AX32r14j5+Gs+E8xaoAz6LisRQwIjrUmLytTciJk7lklAtPo
rX3PEhxuY9tPiFXl0e/MIjaHV1wjYdTTpcnhfSG5r//3E6asWKf4IIdZYlDBr0ga
f48RENnzps84CKei7VTd0Dx1uhI0BMQXjuoG5amVmjPRyhLwukDbsYCvsk6Io9WH
y3EUvoqSnQMne/8r9nHpt+PSaAb9yE8HDH1GqBGc/Bv28hnd2DpBY/lsyW3PTetg
RULo/ZIrYEu0vfAtS2EBR4PraSrPHndict94MsUWX3uI3x33uR/QyL0FnUZIHoR2
21HbO8R/0ioAcbJUtZex0edVxbhUBk8yhoRbb75jVP3D2Y+7BafVFIbReAbnZOGb
6y1BQ1zFgzQICEGhkGjzvNzcwJMeC+owCdw3QuRRwMqOy+WYnylB34GxW7RRhf9i
vnafoaTY4kU4iRXCb4B7vLzxzQ2nw9qp1AQ4FhhwkzTiQHBowgpcH7HfvSXvzn0r
PVy3QMpjNNqBMqywdx/F0uNP9mcuoBr+3h7evKr9xsfxIJmDW6iHmZlFgnDqIAfd
td3Hz6jg9COkZvnWLDphjDZ4QBSqdnck3rT28+MrUMPIgyiA65TtljEpbNk3lfgl
KXaq2VhBZmAbpwcZhPPICcQ/DYHQUZjTRtmxnVsluamjrw9i1aggB6uJmO9aFVyO
zJHEyck4t0bfivPZRVBo8x+qdf7Q/cYJuKD0VrC+x9RZDR754aZV2w7ljDMrR19n
mu5RJb+sS3FNImEvX8ZXdeigOVCUxBRw89/murjsQbcjASGLmXm1iojY0kvS/M/q
KMZy/VutohEGN2lfQIQhWlGZyey/Cw1k5ME6+/WclN23xcN4/oOaPxSVSv1217BP
SFBMjECqM7O1MwH+hwotl5PATmhUFhS+PJqHnV6ZiwUx6HiiRcsEPnMwzClyYN25
lON3DQhuU+unDM8swufPbWXVXqXoK2Z9jBjnpcCUpd6hNg5uRJrKYG1F3RJYF2bM
YgR9AQAcmZYgzjsyWH5KNoTamcTZ/FFpXwbmj6OFQSvIryrEhaInplkixZzDlD3R
qK4Z11CnwiMJVUG5EyWAmRdorJiIvdw8qDCjjwN462wEdwSS/ANFQD0JRc5wXhmA
vaH81PMCeekxIzXeiwUd5c2VM5QVbTqEAZ5cHRzwveooNRzplS7UMM6J9/FE66KI
drSxCcpgj0UkdvKxGOmy7Pe3qznd6dsYm8SLUrZVy411siew1DtZWoTLedx4mHU/
VT8/ubIsxsix2BgxkSIpRPcGCe/H+oiF8ZuhmEpSAWbgJzaqf9+ZJTJ3ibX7vcSs
xmMHs0ll2kFwoX+lsmwmWzLf0FQdVhMNSec4RDemJ3xGqPEqYGpmWLRM1TmHiile
09XjW/r9Re/2lVEr30mNZxeVZZtejpWTvXfaC/mJ4lZmqpkLG7Le2BsBYa1i+2PJ
Snv5fTN4MPkz/xqRLQcc08ORPMrWntcwOrzzzdS7YJAqwIqiTVW0e/DKHTMjunC+
0m5ImU5rbLOmdIMDZ067Xz6ZGaZXyRcNc+sJXD5Bw0urxJxoPRE6uhIAbswq1lAF
ysQUgT3NPBvjnm8e+gRnFDnfyxWTF0KIQARGc+yhUVDYEROrnsLJq9DNq3nh5cqO
4D6XO9C3ZdwLqMgZ0kMWAK/W3duQRoYBtZ4t6Xuqxl8im2UfLrlJZ0zQXsd5WFLH
wqTJ6G1Mp7PcWYmhvQbyQbSiBr2B49fiaEU3QkfEPGKnHEPeng7pDahy4m75nnC9
7TaL9iSE8bvuYEiC9KUi+MFIUkmZh2NQ0My+NHxNIFJLJmuQd9vWOLzb/4qgfWmg
BpuiGyfKgS7C7gd0Laol0EE2z5zULOnsClfydZ2yPYirqb+ouptVW1eMh3tsM7Ep
9iotQfErMLWk+JzgO8DKnwaMVtH1rxKz41PMzJsdmoyFEIXKHfRt1dNfa8X5ZusY
Hzhap1FCe6E8ddinb+TSR+ld3wU4xAv0OLZaHcLN5VcRNhkY8hBvV71DT+t+o6Rp
Zvcy+tnwH809AHWXj1zaP/vHRn2DOJDr7VXmlVPOkFPhiGDo/JstdHIqzWPs1Yfk
QS9vTpkOVvm14s1UXGJcM/GRpPGRnIuiO0huapRFSkHI3lV+/UhsokRwBndQ6Sbq
k4Qz/6DsBQuq6++cV1o3gr/zdX7OWZbZSvpI3lTS1bX6+oAgwpw0qxuEIX96jHMy
gG2KAWikveE1ww9S0W3c9VNN6N6DbLidzAGFzzuRxgCZIIuNezLvDT50iyyxQU4r
d8XtcgmdcFC7iOjiNZ0GSlEngg/ZwgHIuXFBzEm+ZcUfStg2UadrlaDZKHI3DO4I
yYxPymFJVu5XNi/viqK5CSRLZfUzH0Z7AjxTVBj7RkDeNwGg5sTjejU5akPfo3Nb
/VtEN7vio0eO8BfImkskZMmHNf0x/aWOaPA+d/cDJuU1VAY+vhTGyDCXnVe3dv1F
4NtgaX+kqxb3Sr13aGOBts1jvq3zYbMdVd796YBsU3lyxlaBecpBZoFS0OqeViWl
V3FnyG2xoITUjXBZTNOLQcIjx1JGoDoRze2jztSrzR96EE7a9D3C1QZ420+L6o0p
hpdKdfoLKrzJVtn7IZYfQ6TIOkn3s7Ct+W865Qb39D4lPeslvh9k5feK2DzfOHI0
pl+KT2DiCltuckzLsjPIaE/HVPXlWjeCtnie1tNR1Y/sKzXENUWgzbjxQbBOxI2l
V+6Jq08a+VMXUUKICmNmchbUMymiZLNF3KRuk9+J+DpFDbGq5HLfzuYQcu6V7n3r
g35wqWUdReuanwX4XA/ctcuFtoQr8JiU/sGcyCMz3htnXRh2cxVIyYxceJY5rMB0
t4LTll2qkJwah2NVh/+eoCqbASlBAnW6e51bGrrhYO/9CgEoVpVi1w/mFijfEyEG
ohYN8miHAp7u3BDNu2BSk5aZEnUsRW1w3Ifc83ppYJKtdvX18gdr0wlJZ7aZ+2li
godFYK7otuzJC+OKr4R5H/CsVgonsmBHLkSbsOhJRNigUhJRryVO+NGYBL0PIrlR
uRA70DEzGxolt/FcT44+muxxrCJ3O1/qE9QhZzboXf5iJ+1Nf5SQRZL2S062/SO9
IoqL9cjQPid3HMgddAOA3hJrrcGLegdVI9Iyd9b/9tN3FybmyD1Pt6B3qWUMeMOJ
bOz35//8TCGkvUG09TGpP3+KlKaUTljLa0DHIpp3itmAy4D6w+I6hbnbqgGm5ye5
bKz8RKUF8bWdzCE2MNmY2ocaciIWt5dPtK5LYyGWel1KoHz9O3DgAjVddD7IZtGo
at84tRRt8e3lWGkR7byQpwlo2PmzJc/OzoCcw5IfupvegQ2ePsMLgd46v4nWMLi3
LMPDfdxFkvI/J2IWvwJchGRRyijHsYts3SQvfA7T76ghLtQyJjir9uMk7VvDc3/+
SU71nsHZuF6nE0x62P8e1WHir9dZfuBaKsz6he8NT1uu1HcG7s8ZuCbQVoXlcZ81
XPSyqnhrHn7wlWV7EWC812rNp90b5pMB5gqQaEOI/B++CeuvMIP53R4FBOnAqZr+
EEKWZgOne4TeEfFQgiYOeNRGTfFEgVGYkN29Ta608H5QuOYQJNt+sdH4cUeP4zi3
b34BAFQxeJogWq+hCldSZhwdbXNdjMVsfoELXAaR2vEndqNsJkM2BpIyoqrp122q
GudjsjLwb8We6OeFVJxMT5DVoqXQgPXrGEDlv/GQ8d97u+BM0tGwC1foM8+qdojX
bRHgK1zAIhv2MXh8RpRTD53BZp3p5IMPAGJuKefm9UBb1zreahC7Qw6xnD9lcpj8
Tml3ZJPM8/iEiKCRrbAXYFUrw+sX1E6vBqsEnROjLDtGC2+AmSy8feLGckBWltqW
hxUa0n+vsyWvShwL5bKAEeMM6qY8ZPfGvEmvBaxqRFAryIBYbzMEcCdSQKSL+wFe
xmDBujeNPMlQdtYLg4o51HDJV+nvmjcOTDaUk1DjCU//vVcPgM5FDD4D7XICiF3x
l06Mdgpc8NzzuQmttnRXvCECz3i1jZvPdWIp8I117ajvABGL+Baraeb2pa9aXjZr
u4SMZ3WjKRpP5xNA9WX2PW4HUEM9yLT94S/uZsvI5fBzQZp/bbhBPp712lNSeXb0
yjHfxSMHd3ERg87SeXLUac/IEV03BBRyH2/9I7Vr/kG0Mgt8vGLZvXxNRvC6BEWs
JAE91hTrpuwDTOPI3/reDykZowAK+/ld5sSDlxHFFBfNCXcDv/b75olP5K5sps6m
Ehm2nOJpCAlDQCxocOhCD6a6LCmf4Dcl0AOEe5Lj71rmPi82CL9a+lZvdY35hN4Q
7lmOErXaFR9gg0Ry8BYvo3P7NyOf8X3hEBUai/QZWkrMYE457YZ/i+QMwVi/2yrC
WrK1WTpSQm6l6R02w/zxYWCkX5SLIIc4o8QNZCPvi+t9LIOvdlltZCQ/0ucCUQC/
noEhx3cgbn+9OF/iMBzrg7xQuOrwkynxP2b8cANQ8PRHUiFiDVxKCEnFxvHX+ZTR
84xTCpWhSl1wL0hR2t3uTspkQBl30AU630qP0dPSlpjGgDzqSNcpP0Pqymiyxwxq
uOjFfvqwPReWqNscWRwuM6sQ7T654HnfelDrB2LWb/UY197I/LhncLjSYgxt+7NT
b+N7qrbx8QdgY7OOFU3megl2liWhCqSDvs74yn27/FxMABt0nGJPcZaWulUu6hsy
1+aQWZgdoPt3kPFU1PNJXyAKEqPX/rXcpu39yWPNbbYvIEfb4Z3gQTMrtufq7gjJ
8sHWKkeLyBH7zAgVbn8WUZI8pRi/18bD1GDqN3jeGgeXZH8+mhYR7NhV0fap2F1s
sWwemRpPx2zxD52rIvAok286mBUl0UPiwoq8UymWjxnTNtP+JbJGIWyeKTVH8sGD
r+S08Et8JL93i0Rus7r4yp5sCZS46ecgC+avLAxXshM70/ydMJi2insNzfUi1la2
wL3R1SxckJ0vqTOU6f9yf50AGKnIp/KSDgUbX3X0bZG4Zd50S+MulV2Y4gkk4Sc3
w3yyT8+7HekOaozNCU17n8zhTe8qLeE30ux659rFi9LATLAPVscjrzd5PeD2xxzP
eSvC/jy2S6z9U+gLxwI6fSzy2jQCUq7dmlpBhKJT+7JHmqv7r+HxyCDaRubu1rLW
6DvcGpUIFDFXsO5Vdzc495vaJqZ3kfUS9RZFM3c58Mds3mGe4FXuhpvFlxVwPvIr
WTBMnfRL+SP498XKOmn+3wzMzcnuVIP26NOReC4VFRcgpz6avp5/iSMOG0pDVqiA
dLbCQsyjhcckPfOVIxXBcCM/LdqGkrvml381y4RrgZ7C2rVHzv3s3lqU/1ZubUlx
6pJkIaI+/bmGesvD+6lnw7XP3RH3NWSO1d8Cy4tV9ONNL6jzcqTMSMXBYtf5LeZ1
Pz0yg/UM0/QxAoV51Zf7EqnZ4Nuuk/51Tx7jUyljM9UaJ7h2JR50tE1wOzAk2F4t
HWrj7Om6yQuEy9uZAjhyoQ/OP9vORnR1UD24sh5Yqfg907Ie/+bjLJrXdicf3H4K
aZZQsK1w3FfjELxHnfcE35cBHWdxO1eSQH7boLe4ndCywQKSfoloVKsAnG1/WQCu
1aFYFu/GldFxm59k8Bbt+sTe90zzNnhMcT2X9MXCWkngdOxzePujYG79MOQ0XDEv
aibg3xypOc/yHbN9qLG9+FX/+P6GeCtiwGEkxXYuzC+XugZ11Pfl3XsK06N+bI+Q
2u5hbae7F1lYvVK7T9tXj2e/Kzn6qSDRLA+IzJzF13GZwaniOcRDUQ7toMmA5iCM
FywOLAAMEwlJpKc8yTJclrcgxgXFiBL8SLXDCH+NDBp3yv1sGwLMQFGDPO0d2SQC
coppoxYrcIWdtyBT+fB0wxC50Ag4u4BLHadodp3aiZS1/eIBC3a/1xTmldbHKedq
fS6bHmGD15Hh68+mtI8YtUp9E71MTy5G4JtTV60r+R9P416I907AonmtpKGqrUhg
CCDi7cipB42LEDhF5fce1LLuPCFXXY9yFsRvYta0Y9f6shvO5n6CPDZ7/ZkEeQtS
J1zKtxhSU2yHJF2pj1cw5lrmBiDA4B7sfQZ7CorHuNI7JhYr+3b1RPZ86R0xbayb
ivBQR+ensgK1LidFRi7t9xtSfdjw8L9TRcthBBzb9+QbzH7xc+f2kGV2nxFpELfM
9SP5bg3ln226DZU0QAq2GIoS3TObnbw8XCqUxFP7L082vWtzGsWKq8a/mTb2yxAW
IGjAaddoDqOAnRjGG2EmnmNpFSJhuI93265KRBjiOwt0MsEkxSYswCM+ItSXZ4Bx
dUzZiY7u4E+tMxYWGXW9HdPjH3nwbuX1sHFK7biwGtRwoFaGCaXthSCwAR+I6S7s
h+ZMiJgU0EADZl0T6O669lK+l33tHH7cbXTrvjakprFywvQ/rkW6ydYnqv1hkTmM
xx+D0vf9+7flYPg2fDAbami4G4CRluZ2HpPOkUXGl7N8SXMbt1ln3khnNf5PUITt
mPdaykvLQAdXQoG2z1SXxH1ngsIF0vN5MSx5FCzkxiQErvRWmr4UI3BpPteYU/Il
NyXyq50Qy8j75Sh9uW0rAiBPNjfrYFUVnfT6bIH5ZJiDIKe8hnb89eJ+RCxS3Shy
PIHUnjjlEnyju9teflgvdoBS+GQyfswhjXvJGmxmDwSq4hbc9cLiqgVswb+M0aO4
CPzJn0ld+xzl9oj8q8TM7JRMgomprnmgRmaYotraG/tUu1blm43A/+aERR6bqYck
yOduMfi7fzoM5VOXN02KAu0BQnXPzfx4v0bFzYGjsmkEQVv8FMG/ZmqE75I03DwB
FyaYB4eo2tF10h2kdr0lsJeS3E5shKGLip5HKC4W6seAk7pXXECf+W13IJfggE2d
Dsv/VpL5X05uqcEpolD4QPC6Aig9wrtWQl7EP1+AOiCBjxOKMlBXA/7phe/PAkAW
Fg74/JZdlQQZvj7ERLBC/zgflLepcX1HRPPE/Id7AvJrsk7u4aAzkgcMHZAS4MUi
nIlZaPG3h/MUyrT1Qv/Aq0/6TjT/4f17hfp3ksyzkrKauasp10UNgs3BNiJZvYV7
GtP/lqI7SR6DrJY10UayPnlieiBEj9xOv0e+zdZ0TiHF27mDbZWMxrVrWAU8ZVff
Dj701lHtsiX2scAqfu85+ahZjHjAw+8opHJb4BGqcSd28UY/p14m6CwmSSeexvRS
8btLY4jRYGa6s7/nq072UvGX93vT2lJwWOCIvqvwe2Mt0dytFrgCWx3Adq5CUbk3
hLtQYLEUImvd/0PjpGTRhzs1Va9c0N8lB7I7fWPTcNJe29qEye+qh5fUzUK6J8t3
ncLhtU0BlcGN/d2Bi+fSJ12EhxC5CIWhdCEwqVNKiuiD5d2RcEnm9IBGTL98+fci
7U5OtUWLNG/NMj66MIsZ5xSPII8OrQDHkD4SDAdXEgafq7elPyxCf7ppl6GVMXSd
EaqWw+65cvkajWFOCmgSApNKPqn/hsZZU4TV/1saSpZTL7sq2THgdXsD2LcfZGA4
DwZn+YQYXZPAYti6xVpMdDtCfikkwcOkbEEORQk0Nn02HxMhAbLqwoOwVt7vh+v2
Hag6TxPvDvRkKQSNJylII2468xlh20PjTlPsZZE6zSElXImr1IUsQKct+I9FosBM
N7RJGB+a+xwdnGoR64ZeqQh/iWiTtF5A7TonpxHXbZLBYHvKTnoGla06IP5vWkQp
ntS6/PfZqbn0I+7vsxv8rRfIbrWOnbGZanOH/t0tNb5n5FtIn3+pbt3N/kk2doMD
Dh4SbuWbNPR5ENyJ4Bt++zMGhhWEtCj+AtA9+Rzz26yOUlWnRB65Uz7fcHfd4wke
/Wci7rCK+s/YqhtyZ2NJZStq+1Of6jrKhZdAQt0JnEpD3c0h5yE3I1lWcqwGeOb8
aMnvNC/JUNbgVz/l6w0Pxubzdx5PVPs5MaQcOo0pJZUgQrXVqPZ0eYwpgKjn4RgI
6cMT35RQuObMV1VVm5QdlGWUo6ABn69KqNJc1op+tQJecYvtFDWynscJbNGAXyiz
167p5nspUMO8LlJSwGp4KA2+FWBsrQc+D248pquIhDj2ZWISVec0hayxHSo4MQPq
Krs6ZXsKvhT6y7KOxhzHsPEpn2JFAzZsRFePv+iS8YWihU7C73fQ3DnLnS8vY61F
IfmWb+XshzD6ATaiDHovCu9ZPgM2trJr/1TA83i77VebMMdiT1P7GsEiIpVX464t
DmZfBZMH9M6jTdqxgn1LRR6KR4/2CtqwX+K3hm8FPWBSz3UbtM0sFlceAgZSVDOe
vCuv1ZztlwtK9fl1bYJgfxLMPCPRzA5qklCNP+eteyw/dBf4FyP5HaiVrWJjesHP
3Ct9HacmHci+0QQ8Wr7xIEtm2H6WREyulpC7fg5Jzr7MSGjT9HfYKDZoYJWJCnJ/
OinHc352px0VwHle2u5UVuRqh7spyWhI7e/DZ+8V1sLPa5gl4J7S5aBolmM8xk5r
NoG0iO34I5aDxIc3a8GTsokMJtddKtFCVHKPzKpX+wSvPNtM6vQ92HRGAsYT4WRa
z7gqFHZY0mvJ5rlYosmDB1HFFfruIg2k1Eaa+rovbKnj0juf+NGD3ze+bZ9ReYL6
QEG0Htc5iua0D37PauIHMDzU6bxlZZK9s/te0wlxXIVR3+5stW5LtQVhQsknpOF0
PPX+K3BXgS9pgmpgArRFFlZs0F7LV4D6X7QUBaMnOdgv0rAR3/uZbOXQXvwasxIA
TvMT0IQFL89/Ed5xbZtrxePRscDoMY1xq1eCs8Esh+cZR+KBa23NX3aGwJ0aVLx2
aBvvm4dLs8RFXdvnpL2AziCJi1r+dRRM7ncMtUjxSmb+1PJevw7wKp/ojfyLV02Q
AxOt0GgYyqnlRvl00gNKCDvfDRzl3+DzLRLzBUctwrFtvUZR+f8DIliPbw2nma1Z
jp0sedQq+AkjTm+//D8O4BmU2Zq7TyGIurTOCf6nI9Rh20tvecZxe3KWBh7QbH2M
B68DbcANLUT2we5/vpbJ9Nyc7ecIvMvc3btLVCI7ieZCq5naQlIadKT6BmpgAmC7
jexl3L8iW9WW2RAyGCzif4MVKeYNBJjx3HHlKvlHe+Oe1C3nbhogP2hCsV3AVbXd
+bRJO+mXdUyWUthpwVLWSIpHailedppj4s98HIuRQ0BcXAvsG9OheY54QfEphRIM
zdxmk/dR7OfwGnId1a6C0W3k39FLi4EMShBMOIIFr+jlfVL2ty8q+vX0DJSMAPk/
kHgSppChgc5SAIkbLaPTklpmQJ1Mkqi+NXxzh4EpO68NamDuv8t9mszI22ZCMm7T
tpXso5AC/3f7NyooEauWWB0DV1DlMfmzfrEHeCKEFXe4lk+PR7pFJnRvILxMyNhx
KX23R4UVoHcIw8ZSV5pNlnWpFqKWWiW31xUddYa+zMKYL9Yph38kUZAmcfI47zjj
pQSjJZmfia/ih/FagVX6H0Or7BlKothNhZjiTVT2qwYXCMJiMFfrkDAAdTs8Go8v
temOUsEP+Z9Vxfm9Iv0UwBaDCj/PyjMpDitwg5Zrxosf1YGYXorIJmbLPvhYdFJ1
EvfjsU9XNQwohAs8huDShtZFsXSYBUxN4BU6HvUQOrcy8HUFzjMiOejP0c4El8MH
Akg0Q6rlR8MjP69UR/JcwHi5Ysry2bUGnUQy6LEb3bV9XlftYIZT33XKnj4oNKRu
BAf7M2976fwZormIi4SQl4EZFsm142xocvj0jN5ZOLRhPDCHA5NjVWdHOMuUTPCu
OGNrTSnyCN1W9TeQD9G+FXmCcT9xcnFisotGnyjuLmbP2OL4M3OIPZle4KpiBhyh
sUy5p22xxeQ4ZG2QWCwYyEMAV1zTHmU8VBLGmyoyrbZ6/4ygsSnr5EPZUyURjVqU
sAZLeSF2QHAlWwgU6V8h22OUfKXcwfEOz/1z+VcaGCbdER4f6wOS/Txnyj/JNlP1
7MKrBk/bM98Vs2eaHtiFYTEQspO6gpG8hcQCJ3r2tsNGizqS8riXLtogLX7m3yQp
pZ776zoUfgCa3KZwGIzrjIZQVnDmSZC1SJxJWHm8U+a+tTOL/qJn4BGAqb/yl16f
RT3xdeOOuNlZLXarcah0GOmWvBIEXlrUH+hJL2yabI7M9E7ZVSJ4mTDHUCvl9kkS
ZjhxpbEKpOGNcDiz+QwCd0DfreehuoRiswvSsuheKAGcbEyxRBr3AOU//DVy3V1R
MS6I7ocR8qlVNmJy89mBRiSYC0+CxoNBTJnd2Vz8vMH35q0I81muN/J0QCTdHMoY
4eIrqXqI6g0vn/n4iP6dydqO3ZscFmOvaaiMrTtK6jqLm2NlYlTRNJKs3HMewOQa
CEXsQsUAppYhrJvOb1gQksqonF3om4ThfS/QeT/pr4Mxylaqe1i0O31S13hfD8OM
jg3+CZCxeR7zuJ63fio9MIZKGseJi2rerpkxcAcc3JDkT5BA4gjlx5GHbbnWm5ZJ
J+CoqBtgQFQ85EatiqnyOVbyH/L4+znIVfskpHP8ADoGOLj15f5rPt8i1K6gGYxt
FI7frmXnU1BKJB3vR+DePJZHsgzdDJziIPlunCbe+xHO36Fm3yOgrCGMGr5UxRkq
KePBjWzroYyO2gRO6njVOOUz6Nr3BUBfT7c3oKKjOouk3m6JkGp2/zP5gRE9n5hi
tuk1WoQ9+AMxGCzYoFIJ5kSOnrTpx0ZbwEL87qo8lkjiA5eDIZBQRZ5gDAYrv+/4
cy96tdYqaIUHv1WOc6GBPnN8bw+WTsY5iKi5OQWohZ5/KsEVDhF/U6PBsF23yxVK
Onh3ObgSgO32j3ZXVe1K3/QpnC27UrDBxnyudOl+/iO0W+SKYAVk5vfcBKf/s0IG
B/9eyAN4ukeQkGH4O/H/EmdIqgJfh6OWu2hsXdKRaAL39YzIvCXa49WsipdSUwya
tGUgkUlSAO3WgwlKMbthKYB36Cz5o0IBtT+lnbqX+XyiDLsrjXuh21LgIPjaWgsD
wnqflrH1ozUgfVNzwx3maJpXZWmFX1BucXBzYJjEwY6HQoD6HQVLqlZF2JEZZ2Y6
3rNi07u6QiKMfsEUpIO12orhJoIbwfQqicPwDN98qM+n3prtPdO3nVJdqn5gCsnU
3ESNwqAsGSSuQKt4TnJRZd2/GMwRxdIB/5aoPv9TAZISqQImI6Si8HHCJqEYwVh3
gMPbFTntazSNIB7FQpAoZZirNvjoznCfydXdelb+SgL8YtbKmhxvhom9LoH34wlk
K1UfUrCB2Vpa8+P2FnxtY2iNgAUFzu4RNqhq8kirJRhTw0jVX4ADUv96tnkZJfOh
Ixn59xKS+fQTQBQWUrC1xEi+CeYksl4+qz0CRxoazp273X9fLr+IlHXHC75NLndC
cUypWhiK+KprjppjqAblhrfH5zlkuo5+3CDPQVP2JtfNnw3UtNCDEznvkJ6jKCAI
TzfC0WmYYQHTH+W4b+sSXb8Mf2d5i9R1Tn6A5WLS/EpLHMKM/VT97aDsYzgUXN4O
bTQ1iqgaLnu/d7iO9q6YrKmHADL9+GeFjYgaw+BMEehippQvt2/blOK3v6C9Jd5M
ePm5V+aedJBQ+w9s39cGWq45d8lARbUBQ48weABIeoSO3toVgFAFljuVHd/RGNtW
Iadph/esd3GCo5+icHzlEmK3SPmn9TXN7kxt76qQ8c/6int+zU5uOzHYxPGqenC3
hcP/a9mdrb+lLWYSOirvFew14aWvNVq25a47YdXOG0jrDeg4tycgiroxJZsh8Mk7
3CTmQLcCLcQoeMuE69Rb7awqe36BI9bqDg0lddxL5Z2S2fzlAsIzY2jukFCGGXpP
DVOsVnYAt+wLbHScMDO9UeZxWW/qG9l87vdeDBeC4+27s7S4j6s9xEnpKImxcOgR
j1LuXqfPygNn7jJLkkYpZ/mIfPRPq8tlsWOCXGebcGdbYPJ/TT3/5Bj5OZAQcS/q
NZoAJVhbU7CNbZfvRT/uihmDq+PrhCBro0qQA1tVUIwi0sXyYXl7vnRTjqAKRZsM
IUokcQf9AokZLkaqlRiFBkaLswxmKv0+k6eE+CVeR6po0rLmxq9ZHhY+PDYV6qAe
aQrfivfoOBXZRv3o53OC9Qh3SCXQHSvFF6pLeaYZISnorqy/DUQY8MqXeAWTlczT
zv5bFmyGp4DuLG7roYKqa7/dWg5GZswja43Ce8tRZWDVkp10+sNswkz559fJwGRN
j2wbWdhZO6cmIQPWAohY0tWCzOnKQjWuJSeY4Q/33fGbsaVCazlRnN+suRKVRjPq
J01nvJJlKPGz1PLylb4vKEGcPEq8mdAmc1E4ZnmHun7h8M2Ee85N1k7Q25giuq1c
BEwZsIUHCvRjJGD9JkqzExx4asrH4UIeEIr76EBDjzjQ3/hD32T6CKJctC9c1Q8C
qUHxS7vrdIMiulrtH1N1kerjbgAVB9rm+ACSqoppw8MvQlM14naHPT7Y+9YzUwn7
O1NXPQYk/FWBiScwYkot3rMoVkai3oIbkP1fL+05hJ29FCOAJWBCmY+FqV1cD0cC
c1xVffQrc22K/ubyL+Hw9jIJq/MG1mW7MJiF7AKR7vF+vwTDViLfXl8GQfvxqyCw
gNnPJ+/NWFDyJAEipAGYSUm8yYkLOI+u0AjlGt2FsAvWVHJ4laYWMfna86ad4/DA
Xc18PaFcnJAYhdWKOhBa0Y3mUQJi1sCTHKQSYVoP4CRGsmCB3kK2mvdNuCK5THuw
1+JTZKlc+BOMJpGqDP4xNkDl+MgPmSopcqoAS/BzYUhI8WsiWBTQOFpvO0ETEHFt
A51U+TCh/U1ZDFG3ABrxsElTP7J7JkqFrFDPoiavNZsHbnhLWo4kDhuKeCPtpn9k
kmNdWwswY8Kql+yOSqn2PgE3AwjFXS/WdYfa8gvKN31JggjuIZq/BXPauYhTjjPJ
Qr8S9nOBc5e+UO8t3M6nmZpLFHCHWd5A78f+m5x13IrRnQoPk4i1vGVpk8lapm2m
5LfU2SxDovnHMhCKc7WzgGKzUxHpwejWiRusxVjxx1C6t54Ty0DcgYxBlX7rnkhL
o6jnvaFjFZgkdEW6SL4tFqFKOuuMFabAV/Lrb2C1ChLoKnRbl3YRv4p+C0+4Y1W2
EXiSBESb5icYqRgRrBqVZZ0QiI2Wno8cxCqw7qvig+alSnyyIYBHDOJ1rcLT/5tP
R4UJNncq0Awy28qUEG3Qy7y0Fi4jmQDajCVi72LD1unOVAFVff35C8ddo5eq3Lpi
K9EofqR5svorxQGuttDIeqAzSZycnN2BOyEoDUD0cEL86oU34OGatLxtFzgTLaHa
GFGRAc+MljipukYCOoA8COlguhn3BpO+wajuCFaQHkQNdvfRYh25oLw4x34INVWQ
g4Lhbmrx7zMvFddZFCRdCKocoL5IRjIEYloiTlUTO8y8ZMQe7SCOWEf+2yqtRKXY
I7iqQDq0H5iPocSsXBF545SM2McvLQveIVlHN2a1KJlYDn/Ipt8RhJ/A43J0I3Ph
FOHT4LvOd3XaVsjuodOOirOHzOga/qBEn2jqR24g0hMiRsndoZnxFAHo5IXtF3DP
Qc76H8wRUsAFzWTzhiALPG6ri8aa/0yWV+83Epkov4OoMYq8S5C154IC8Xa4VQba
kX6X8uc/FxL0yqC528570PLXVNPvXVDoV4xcTYPS3nU+XfsV54Sq7PgtCDgTRSCo
t46oAgSOGKQtwKZJUpL9HuY95txalNhsb9vew+8oX0RL2EoNL2BRngorZ1dnvRIo
leMaypBFmOPF6jG04fSdjqcdzecGh1NW4lCvMMf6djfVrfcc6YFQCTRIm6Nda7I/
lXzMEUF4uGBcGM1OPP2MktQ7CqAuWQ8o1g70VOPcA/3HwXXdb0Rf7J0axftCrDt8
VEpwSS9hUfvEpsKaJrn9QvLIsPW3nR1U7rdxhIQZo2Gxwpmgtbcorja1i/47GeSq
xXQdhvvNiX71v7WnXwKjkbsi4+hKZ7QWCjtb/0VPYKBcO4wk+fKyrEzWmRCuKbv3
XvNNrgHAXHR+iHrJCCDKffD7itGzgliabtAWCMlTisxxXdtkp1G+2mCOw34MMWYz
hUg9YjQs0LJyTAf4jYrfrjD5J2lr9GsnU8GI6zxHP/QwYrZDa5B+3LbuqoNvOaXG
qt4kPCNx+OFF2ZTgQg0v+NzlBYYkMy+0sewH2NvRc/oFSi6oNyODZVxTH3Alzywc
fTBa8nfpirWVH3RNUwVGsI2JKtnVbfvyowSxQ3H4uBcm9umTccB9dzn1r1txS9ry
n855IU2GSL+1ihe91XvQDfa49tMIEe2OfGvCPg2pBiYI/4GzGi4ikTh+9qrBPE2u
cWwSAvrFB6CD1N0C4Psy8259UPh3Gz1LTCwLbUHSXr1RgsgarXXfwi3hCXtvhwCd
CIXdyuEFk4WCsK4bmTXO/VGweXCw7B7rn1CxtBZx1ZyF70qkDaxNzY5NDvggUrZ0
LMjhQKIZYdIeAY05jQBtZTn0Fux745Qzfa6iBad2UtqlarK3k5WlA4b7RCBY6GHP
KhKVU1F+7rup/MVnUXAXxuK9q46yaDgn9XNBgjpuXh2jLrlWsGXA5iruXdjtgf/c
WwEfgHBGo5CxY1eiKSUR8xy6E/zhq+9kFSUHWXJsJQsiIZNzk3GEUrp7Y/PazK0h
TIPiPR1UvqDoYi1ZXEajvHarWfLb3E+Gqdoxqu4oUj/ZuYSGFaN37G3dcCg8bEYu
noneON+H7Io8R0MmSGOxFnlXuOQF7iXaaBYNRGlErpgA5ePiKN0XmAL5M4qfk12h
mhrhUnmxTDuFl9ccVvcQb0B0OGZvhWvy1NWERe+N7Wd5vmm155wEh70eZDhIl6u5
VcP8ZJE5gwGC7O+G3izKgZRDihBXeRxVa3lrbzwrLwdjVj2AZzCNn2DMmCROyG2e
2n0ckZLo/GMsmr0Ij5wTjBSwKzQ4ApHL3R7bsc973QLZtNiILdAyHXwEB5zkx1uu
ErC7bq8Sr0f1rul2+HsJwLL7Uw4AQAgT6W0jvm1w6WcUhfZyf3e/CALS4sTmoTTT
aE9wUVUjwKWLoxnq6FK0mZTf8stYBpX94wh1DFl+dmYEPupTSSjCjvldmeimtHrw
9K3AEx1o7R8OI8XPwKm+DwymxJz9s1hOi+gTR913KWylzs3RcFgPr62U4eEhNR9x
aHV9NCn9GkO13fW9gHs3kWudOMqhzTNi4rsUZRbrldviFXQWo46DFUQ58Upst7Sv
idkeuBzsh2QiXIKj4v2dnxcLflTgNLhrrW/2Ulq2A3RHC5VZHrcjLCZC0GuVozGc
6IjaQRdvHnrQ8Sa39ApVYeyA4xHbj4twVJ6TmmJ8rOMS434REXSZPNF0m06iwoq7
jjYIiaM4RbyrLUuzybb/pGd3ROvQWdTQvWRmfYd2WCON+khIhd3zxOKmdZ1ILiWd
OBbyVy+n8Dd8fMHt8NnXUChAOPOoaxED6pRJh4MPIQ2zNye0pIv9bvW0SF3p4ZM9
0ZOKT4B0PhYWV7rWLFQ3YGBFpA+IFtsyRl6XAnZ+db1QwAxqOy/JLq/Zhm2Hk1eB
voemOwV+nXjEn1I++b7UVlghrYZetPDl7zTssrzJJQKYfGgH28N8j9+xeJS8Yv4W
GR9k4zw/52iHdXy5bRIo9wMI/zuDrrEgBx8gsen+tGcbNqb53tezmkNh1D4vJNm6
O+wLK8QDphKelHF32QT+3CymDu0npnZug1Cb5WI+CZ7Im39fLZpjcYT3sSMPi0Fz
OZwNj44hKxX39RJ/AXNvvkcFJqFBxKkogGULWUCSBjQKab7lEjOrhNJgduRQyJPG
536HRJ13WZXiVxn0nSVNON2l7goiNUs9u+9hvHNBo+bTGbe06Zppwlh1LBMwXV7Z
Lu7D94AZ9EMy161HM+gd1b/B43gl0ZGtSUoqymWgxbowIZOthtw6uaomIFvMYis5
g8fk+JVa++c6rpj3JKD4Iz9OhfeqKq94nbJ3oqZ+gcbc3hJPPntD4AUp93v7wA/g
taJDVi99CDJA/zuwBf3FmsHPLFY1mU+KkVl4v5cU1r54/eILWl3cduh1RkS1FAGZ
3E0CzX0bCc/JE0v45pkOFSp4wrU4PvRa7zyleAnu5gKnGLMJtzqjkSru3c5/fJvK
/3rFvzFizd4sHKvjmw6db4pqylDHlzgSybg8T4ZwqTFT5wqwXe2klKzE7HQg3cdz
CTRJ7hn1kTFuiYe8u2xEAYpSy260ziOV7ABKMxRLu2+U0ga4jk9nnuXRDMvbADIL
EFaCssO7op9La+pk2fublN0+Abcj35E115UfofptVP4ocu4X1UEum7WRw7YRUV/m
ZsXKQm7f7Bc9iDp1yCcL2v4K6WVHLrl/2s2IY04A2cHWdyn+5eleppjKXQda3Qkg
TyS+vXS06oI7i4GGg1BKtTz7G7jBNtoSGR2C5igJaVpKvYof5rFx4JP0rrl5bmve
nDvjGZbzSumMmMH1as4O7avt/BK19lFlPvI93pdMtKT4I528+U+qzIf2W53E9KFC
wV7PRl7JFqDOB7kJU3qP3n8KCjM8M9P9pGeCyc0yTLrT3MvnUyiVq+wRll5nBD2F
VJD24yzBYqIbMr2PMKNI8QPlUDiY4sPWMY7mUC8GfWiziXffPNDu6CyUGmQqSZSS
F02cXXAUXknCzOGQKGeBJ1BeJeSboX5lYLE5WGXBLH0QQ7+OO1080iacW67YVTk5
tDQPtu4IhJoOK15jRcg2DyxT53sQQ2lE5Xh8jAKX6iOr5ddQ/Wc1YSs4B63ayYlx
XWquUoNP4h3qEa0q58v4P1vJwNNdeBpwQqj/eKxMUZ6cn03bOq3U9mF+ytz/zvEz
X84GUYAbpiXrBLXKnW/KMFvPKTl3aB/wdVSx/9nOs1M1uHHvLgIMQZEv7SwywXHd
rJZ102hFeJpxBqknVqMhfyY7t/WjnMJp0/sVglk5B06v4ViToYvFWb58SY5v0myr
Uvv9cy5VyklY2uLlIk2bzqGkrCChM2jV31zH17f7bEN4Y09FMXMEeZUWprXjDgqk
lB0sv4QlRDQbfy2RYbMNSsIfxwKvgnzEaJvVSD6qKjJ1KFYfLbY16svP41ZFGanJ
5ABGhnjJ680uf+DsgjbT2tojxyG5eXZcF0LvSgUncLUby7ZaKsAzEwm2lRVDODZy
vNBPh+rNVf+yEC+fLIsEo/RsdY/+DTA0aihujfVVYmG+U7DlqER9ImPnXUTQ1/BD
/FJN22AK0sUmNNYr8eqX0LNFuF1oao0YB+K433C/tnBRNob4U7X1TnLKfJQIbqOF
I20cOKBtpYSS7cUjMNCyNLkrQehNq2mfjmr4Z226nckgNQnRCMab3UCAr6lkveb5
f/Rx5BFXHr8PhJ1toSm/Qp/HsZ5eE+YNBMbifz2Y7Qm3uNyfSGTQB3QK4XnQY4CF
WYY8Zo4OyXQncSBa/vkpSbXJTi+DGHhFxMQTvXk+cGuI5j9NEeOARL/wXdkzl0p9
VENw0o93Y9eP06wek+R/CqYUIQePYKCmGS4ref01XlhBlg91cFbSb8EJyS5Eq64Y
389IHS0+byWyrSSOuZCX/1jvux730zeCgGJessmNyXod3urRbSHUwzOodwLW1COW
h4rwZtLLzcb6Ybz/2w0Ff83VTS436ZHeCjouI3JhiP5MGNGrTH9EpvHytZdfuO/S
Z9Hpa9dpcl3bvvhRB4UYb/jREVdZ6M7dAYFlsZ3UNZVXComzdMYGX7hA7Rxc1qmm
q84HReZQrOMMVe35yHEyIt43K23zYCJoU9gZVoj+ksyIosUR7id5TpdSHstSI77m
gv2+j26ipiZzCJa96elVXrvJf3Zhm3Y42lKpRa5zGhYAyNSK/brZLAxlGAVy1tfu
xJgeWt+5vri69UpiYb0UfU4+uV0O89MVDfxfRWqaY24mNqpuUdWRlx8eo/0gYdSw
sbM0vTBns12QFSmhAs9lph2sRv6dDQ9l2roj6aTS3FnYnLPXatmn9EaQ0Mcqye6d
sEg81U/543jVw0Cviny3pcsft4ARoa+tqVhASSxFmX6URL5Lu/pb0VtgFn/9eJuN
i73qNVe2aLllzBXdnDFRWTOEsOdk50DNwSUq5Bc54ba/vXOUKO9dmULYfU8KHj1i
VBwGCzKLT5AUsxWKXDfCY0343a/6fOR27MZK3zOGqSIECoJXJ2k0CSfFhEEwyKU/
v56dYrVo81e6PijYtmMUSsk0SbwU1tX6tZDVHvuITJoPRZEm04xUM9cTLkO/WVNg
IFEYQI1upmcREGj7F3PYM4KfbDnh4tiWCMEi0HXY3xZ3vp2H1VdI3yu2iY1aXEK7
xvRc6fkwDHSq8vp9Znwh/gslAaUv71bbrT39fl3cH8Zw8Fi5JGyPp9BZRbwlKjTi
dRXVe6E2xsBoJvyNQ9KXWlcfxKElpcAMkzbDGEKHN/OdsgiFskY8awuJWhw9ohmC
VDzcUiExe4X+LmY1y0bFTcbCDt0B1WSh3SEzRqlxUf/OWHX0fWjAruRYb/B5j4QS
depXt4vE0SYeWSb+GmNSUNaXovwjpqVIpxHh8SojvtgM6VmGTajZa1MDHeJJ688h
O6BwIUBUJqbDpQ7u9DYNaXq+EAiR2++cg9cCrbUje7MUwja4DXE4zOWmTTZo6G9Z
iq7L0DqoJ/gR9Ev4LsmtyPOW/oWpyK4AG50FqVmqzPWzvjmdVXzIxIRRLC4+86pT
x2X4+Mrfmp6LXIsWj+ebz9cKU+cYN03+LozqucOhDhnLTAU9qDXuNwbh4BrgdXaR
oCD1lSVC/0LEk3h0yumsJPkLX+wBMMH869Epj6dPxEAtyrYNduSyCGE86170s/pC
9qHUMqMwdndFvxhtxSEYBK5Rm1+XU8JH406P91d1orlNBcvQMqBoS6SQILRfLwGH
GuT74AY7uobcsE7j5Z2cMLGjTr7y7szAOn5e2l0wC/HWRmS4TfnQrccYocFpEkQp
KzVn4jzp1xXpyOBKER3xoBvU1KtLamRhD2ya2NjcPCFDuqul2e/UE4F1sciciUcX
B6ZkqO+Ul/fFjON+slxB8LoVmL+vN48VTRHGN/knxBEXHVBytYhxBNY85mPoC/jN
QvBGBSqhmaLxoHRbglCMPbE1JSBhswi+Fo9t3n8YF4I2O7rHraXyxDP6t72ttzke
lwvkFdTYLd2aJR3Deos6aoReRbAL+P1CC9FgqfCIMPL9hQARYNKwWQqXEqSgBOrx
iTVDSLRAO6AYIILXBxpdc5iylKxsasgQoqWOuDM2gJHFCn7WX3abtTI/52aXzk48
CCoZdgxs5/1eQaBh+ike4v9RTEIPWmM8xoW4U5UNd993MIWNFtVLAweMXcYsANkt
AOMcxzHzJGp/tDcV+9gKUZzpBE78hsjsRrcplQ4Mb0Qs6joMrPcRkIqGYh/wqTkn
82T8mTRJGQKUlSX9LiT17qbuEulLDz1d7ubvVP1GXQUL9vGZvqz+fZ0y4VFy5p9U
CgFlsJigpIRlSXP/ONsBxXfjgVqF/7+b3j/W63Ru2MxzmdxeoRgUMvwuD8s/e2dU
vx7NrNcyLib4xI9ZX8LNpz2BcoPIjBYVZGqADfNdknx+WDu0hI1VNDzSCz368YOf
nXG0g77wyUfRsb0wxCgPZk0pzPAexWYY1G1KGfI3s+AQsjIMJ/ys4SfLlj1HU+tQ
rq/2ZL3zYjM3EI6fPbVvIDtLjeLP+K5cU4XzVd52yytquK0FwCun3pPLWGxRVjD2
9TW93z5661/0eRf2FlLoqNrLd7CcXuNWct8ikmXcMAYFa7fkcTlKPry2DgKsG6UT
U125PiK3PPzRAtC9nT8VurJ5nXX/NOb4q5JXisaCQfAgW86PpWBSlYHhOw1qfHBs
QniCNdXP6z3gVUWZIG3aTCI+m/GQt5LoRlQDLw+nAoGLaXb4gTirga8TCGMw9Lrj
INJYlKq2l852P6zmK8hG6LZ3xo7d4Cu7d95aYB6J8ZkT382BK366t34PcYvVvo9R
jOsVAYjUVf6Mz3KjCCg6j9V2eZLgK3ZZ4nALy1wNmroBbCDL8/iOzAloPqTiYx/1
J8dDnIpO6e9iSWwDuWZ9lpao68/zsKlN9VpVPZpzDZdK8iRHYPdmOFFBVl1b8Rg8
xvjDFw4VVKhrBInj3BxbMYoJbpSofxuBmMH9AHXBKyd5G8ZWeTchBpM5Y3jmI9AT
sFVCUG4NHw7RqM77+azQDbrUH/Yot0SyBzxzmnkBxxXVcFcHJhZgOLX9BrKfTV84
rqA6QzT1ZV9H32GlvFZyQUmBjhaIaaUgfT1jTzkxCOs2hUYrAcuYuq7FNz5pn/Eh
Z670yyg8GWXnDJrPehGy6Q8Qp44h+d+hsMdfuydGuW+tq4DENLZ39vdmwYA8GeMy
Zfg7nRDO3Rb1IHJQOkdM0DU/t+3N+xrB5joUBB0pzSS4Dw4u16EGOkSrweaIwSWY
My1gCIbkcxK1zCNgOzygmnfCPTb6yqyl2Vb75MUh080U6roan0FVuu4YeOQns/LE
ez6hQwIEnJC85c+ceGs2ugfKixgqx4Ib9kgv/Sf7eWfU9vP93UeEM6ckiD675awL
zhzAZwpdJTI7c3FkGLTbLPYW034/Xzg5APUSi8i06Li4uiFply3WC8HZ5uqUMWc5
Z4mkIUA15lOP06H1AMePVUvk/2WQ8vGVi3CI2kprRG0SNbPlgiJ/fTifr5ulmSE4
mBXZSP8n5DjrSlIPOOxxcQMBrlWqzeOylOvkOsKSKi816bYdWhMCMKF+HvPKW6QM
u33jZKcMYHQgbQy8ZECBO5d7BEnWHYUfb417nZzBzfKEpGuLuz634RHkdD0FRKCx
y+Zk0sRTZzXoR0CwYmC+rgmXhZEiugluaehNYthLHvx6f16WifvNv59UBVyuFNkX
EvsSihGmiZ9DuzAY3DJeBFmlTH8RQYbgxe02IX35+TZaGNy4RXSxBRYI2tbtcX6w
BMkcFFoAlVU5/gxBznjXakOWBKB5iaZrRGw/5vvL6scYHg5UEJIEYAAs3zfQtQFt
W7JwW+9ABywoHYzdeWzMDZyrz8X9UK3qUVZ8CmfTAlgqKqICN06+2xBlmok7pwAp
BlMkKA3Y5tDbX3lXQOiCMckQcD0XsAGQd7R37JFJIgY3dWIQjLgts79JdolFs+wD
3G4w8IPLxvu1JdYDYmQA0Dk3a2tur0wLtino72jDUGP6gVY2S6A5r1UYuJ+OvU4+
wsG10PLsXqahWChMZ7dcG03ezVMrpgtz7zRDVUIpD45rquYjTxd0xrjymFIinovA
bmUmaxuAJ97DNWGyCy1mUzpnIys5Ny834nY8abXmF4AVAopIFXrgBUhwokjzzhr9
TtZ7QYxA3QAtmOFXn2SET5iMgeJiUwLj0JolnX1yLm5l2bR+6HSipz5r2MA+XVpA
keXzOi+s9hLsw0CDTDgvTJQtxXme6BAk+BoHD3ocPys3EkFlSoVDob2Q8T4vGEY6
wCf14S/yqj33lrJOcPOlLYZBF7hOGKvZxA7UgiSAUas2yT2098gwD++ocgSn/MyI
74peMDUovwABhcUX+3AZaQHoTH2pqe8Lxqc6p4rvrRZabpBTHk9jC0CybC9TN2uh
bFl0bacy2AHqWbd5F71anyCOCQTkNT9uSiZrXszHlriRV+nzwjR0vtKvkD3/R9EE
Z/d2MKkUuEed6i9Jzpk2Z7DwfoV/pXhmYyxVACvw4245THuqpjxkxHsDh2CqqP20
jen2nCNZoQLe2nh19rCy7+CZxu9Oybt/SLy6b1nMqjMiZYTPaY05RuQvFBDWIdtg
EwDHsldNNrwOUR6le7TvnWlSFVdw5LcRErTHhF1Uo19qYZZ+ese0fUfAaR3xzXbs
3Q4jckeecd1q1sZm7hAVf4rHQVkjDs427pjSzyzjCfvaaFVqjzq+VcRdONEV+Ho2
YQVvsgyNyXPz9LRJW03FK7Y0eKzXB5OtrxQVKdMDgCpiR0GCSJ9wXFrbsEhRf1o+
JKTH/qtSaeMQTNHaxbxzhNbYuJfRfLH/lt3GIUeyTVTTh5BOw/zwYzab2hpflbO1
00+g7oFnQDGPRgr0lFa1Y3QDAkHQrjjXWKSY89Bzr9hCv/C9Tphvo2HuvNVILMUB
rpLcplCkhhZTJkBsar/XHIF+XFYLOYIOAYnpi31xvsQ6kSMQ4Ncv3HcGCWQrIi1K
NY6xKk6wpP6ULpcpgxoIXcfKFVklITGTzfv9A7WR7YWR1SlmUM2ep4jMm9pttH4S
GMF5WLt43mQPDIE9vlWabTXTLFdYSGR8LZFUDO11sWiu+TduAuEXnhRFGetn1uu3
Wi7QHJWFwxB802RBB0BGJetEuPQ0y2o0QecE0Syviv/CnbBLHHIrzUC7gknimyVy
5UjjqOOSyEQRvV3Hr2rnzjQEVay1dUlHUg1SJUZSf540yP5guq7vfSEMyqIngbla
ZLdEYXJn9g7RWmfHijuDRFphB3tkKvWPixwMlIGsyOrLw2CaMCEds/Onqbl7TRwx
2BO5G4QP0SZt8NQxqLa/yQWwtOqQ2iFJljQqj4K4wnLUpk9hQuHblAmhMTVXbAXs
n6FuHiyvzKi/jov22ruq3mY3NwzZPu3CPgVXpZHYoZRuvlg0gUjW3BkmENM3d4y1
ah+Xn8FOo3c669th8Zc4Jj0lFeME4/3qNLfapKB80h/g1gEV2/wr0dpr0VatqPMa
O3Vv4J5jzAl0fbghjjJsNCVGJzxoveKK1zrJ58zh6QkAEXLvjFSGX2CNlbbWezGu
DkAlWBhhMQjOusuLX3IxxKHHnGK9GZbZmGhpn6Wdc/9H3xNSFZ6wcOaGjdF4FPd+
EixvxczvsV2VGMo0+4rAqLh/SfvkCKP7U0Fpg8zwUokcc1DiWGtJZD2vHXInA2AF
hzTUjNXcjuTO7NfgY9GT2ZjO85vB0TfgbE1hiURE5YEXigkfhhVHgEx6yD/6zqfg
0AUdayIM+UQq14wclZcLECFYwLyUMkNY7t1lHyK//EVDe78B3eiudygUOm6UGA21
QFVqwV6cX/90BdD9cQNfnT7zLjvx9BgtnQDxLtLw2tITQ4vtMFwzB/n6E6sRlouT
zGvdPGsDW79DwADRqJSH9qxPB/SFUJ6KHNKH0VjskDh9WftZwyoYO9q3ODKXRtoE
6jQVx1NNTaqYg9eKIe0dAWBlGux7uPIjT96NyZ5dDhUotsdoTExaCh8pkRF//ayi
JJ4zP9bEQHIg37ouEkt3TL2N4qo802d6aSuif9OH9Zse4XB4PJDCTZK/1ZiXuO+4
oXXFfr4dXDhg8lXLWdx3A2mjzqlQzyUMnOpK27CP4NEYD44a1PlpUWCj0cYfiSUn
qxmTQa33aWPDUObtof0sGBVGWZu66lo/a910/irrrfcjE06VEAFC5H7ZRIXmlOlO
jIUZ+VBQ9BPGQiAJZzjjDWmoNNuToZHq5pE3zrfJUz3m0hbThMlODCpWz6w50Sic
86wo3mDEOp9ezZlKW7nfjkf3gCFFSFfR9AMZteV6Ikf7YF3vk2qDdwgfT3m78orN
RSe6Z8GVYKsZuBX/QFTQE/JN9bXf01vvXk/jUMO1MxxyOYXbCj2V8tHTdLUDZ0Fk
YkXQb38fQdRW+VA4FXv9iQ6/bNr6VCjWYiiX5i+DeSafUCRZBV9I32XnQUjW7huo
ZZ51BBqrKqM5AA+MpbY86isdk3W9cPdFoiDB1x+dBB8ViwY2yRdd2tjaohijqM/s
jTAUoRiUcIJmA/YYj2X5si4fvOWMozK5CJ7hHVL4E0h0Ss5+nEG75zm/oKTQrBY1
o2jpOtn+BRaxiSe0Gb99OVXPrt9uCXp9f4RE60GNA+CQ9pb6Jiq+lYIaLAlWtCcO
0dftLZ341x7VWBYLD5m25dTw3pNvZpx0+qZmqCTPU36Y5lRB/ueQ4pwpPYxxg0TV
27cibhT7Qin6oNwo0jM9n7TxWYB81+4c7njtoBdpgC1pDU3Qh2DfDfX9p3W2TUp7
Qed9lbqKahBui1bxRqGuAA5ZMt9kh7k5ac9Ujvtsfv2pG3qO77mdl7oE5VsXYL0A
XssHC5/76RD/yuZWClhz5Ou+9JN2qLqOMs1LiUNM+sb+R4ttUcGRrJvqoonnSKr2
pSQpWrw/0SP16bSM/SEqs3MslWJxkeenFcZoH/xDMzAp2zbeCtktYitpvecRfW8l
Z/b82lD5FJV0rYqvHtm7+j4n7HORP9lUB7SBblTmndkHv42o05+ajrF11F0JGQbl
wLbcuMbKL0HOqKt7sfARhjiNxExE/I3YsAj9lPaKCK4aSm1SL+VbTsxBz48iABLh
9633w47vSDA8iUxT6nd66jVrQbgdOaZK/8GgxwxoGPlSZrCV697Iju8mEO14m5me
Wdrk59T+7OtJjNhTTb6vtoGinik0kOvtsQdNAnRgjdE3pBUaLc02xhbuehpuL61A
CKXw9jYGlIu/wicuwtTz1OwpnkLTR0jq2bH/IfTKP2jkUKDvjd7SibwwWRr5WbpK
g26UG2c66q4Fd+j9f3zGuaeiP04K5n80XRu7VcXWODsXd4h7OT1gsALqq0wFq7O6
PjJo7SZ/XWMoujsjpcTgK8eVK1SUmMU3RgdT8Gan+VBBtl3NZdENa/DvgRW0xaug
B5BRLxO/9vG1urs8TKc8S/SOy+tcNJWy8Nou3E0ssC9VepCLlZ1UCaCcOnUSaDv4
U02Q/E/JlZUVDknAVe91KsTzBlcyYtmPkPvRLdUi/qiTLX9IGtZcutRbhXuVQMfY
IgL8MRygGFuUdKbmVwYCovuYLIV+5zPDxGVgUs7uyfz3lmCCbgLFmEUZZa9Ry6ta
Weay9krANRQf5u06rQNq3ayZZ7mC2oB9VH5aLBJJHVvYkrfgb2JywRvwABjlqAdi
vmy14a8g5R0GYqStItguC7dHrO5lcSazKg3GnYKw4rEyw7sUa/GaHHufCmK1I3aV
djdqqBGpxbKIMR81wL62asVm6gUo1Q4jRGVR2p0eC03ebvlOPn99SSTXvVtXNhdN
QUwEMrTNFA8cOy1lqynlUXivpEkWO/2bwLajlWedN1JLXZ0TDVErSlDCkeDHqDWe
6VSBtFgJxhRi50ljBUHqDWbAX3vdO4pNCogZDXu04nVztQfipeKXUpx95P9OfUtF
9Gqdgw8vrv3F+Ze2OYMLrgpTnAyjGGOf4PIfD+rakszr3zqU4GmE+Fuf+uX/iKNP
7XYCoq9aXh0Xf4ElcLERAzI8QFsCsukXdaWZFaO8/Np1zadqUpTEkZof/I/ex9am
jzy3hAmC9nlZD38/CJKlLqUTi6lYLCE8mO8OG+tSK+h4oGdcKsjjF4E2DHlq9rhI
wzbmXO5KNZqT6UqtVc2kuGBP1XWGb6MiHXkAR2n31/C6oQnnJQ/eEA/CuN7D6PLG
aqhmcpeX81xi+lPwK7PtvCQUO2pXBj7/vDRco+qvGZGW+k1NWhOth8PhmPfpFLW0
Fqlt8C1AE+pf5/kOLUzge0IeeY4kRDYo05uVgQodtC8TkiBZJKfzunkfNcm62q/6
v/nTDtzcLODPSreXNLAsS7TBBlZYQMzO9bRPFs5ckyF7s/59/D8XdV5mkA434e3S
WBQVDFiMY2aMuHf8vhQjVT6tzczkXe7JD0zVTDzO/5NNcIrybZdSV0Q2xBOiuLUx
Cvk6RbyQEoiV45yxgqPx+kzruxo2FPfbnxtWubslFPLC93cla0Vce/lUpB2K77up
ctzXIcGDDUWPlV49NHRXSBrhL8nnwxLC4IK+H8EOHqDB4gkTgXzE1W+DwemO48i5
gnyLpIUD8WGBQdXVNhK+2DYcgwdZcbx8PElcija6a8UJVbhmSzepGesSzMuuXGff
FRizQAPxzWPyr8h03aR2E4m5HLRK4qCN1osW3wfnmbstHlf+zNMuB4eBuRTYIrm6
+L82jDmZOTAMIkEu4GYxnPZ6P4VWBG9Kc7T8WMOTFV5Q5+9B4RJiHmDkE7+9uLl6
CBs35tj7gbvSX6ZtXeYHslZaD2d3M/nV9x6/C4O166iksvvEPQcwNCiKHFvKm9Kn
99YYL4O/Y0ad3QSuMBPRaJ1f3nIq4Kj66FNUgJB2Ot9z0IEFhBeARy/rwYXtsVVJ
XHpiVU4wn6uRqReh2Z6cECYhp+F65H7eF01JkGFq7agcfbwJg7hqRBniHM0LJQTv
YLjZONRY9IY3eHzW2yZRtsChGWqYggKgGht83rnL7Wl7hN5CYAKBwvK0oItzTzdI
9yhZ6epQtEev8rPZ7WELCGk+yh3N7Aprzi2/97HYTBokfYqZQjyAij7nAWkioo4G
5VpKOWT3IS5PLSd0NmHqaVEo2fTMFSkeT3TFzRaISFt8WLC99PdgD7XQBGyXfvmJ
WmSGGZ1m6AUSEashzHq2Nlq9fH422Ncyq/RbOf2VgFC9Iz0ZEnz9sgqLlSZZjwTV
ef93Q0g/KuOTBLLyJFuFYKkBDZE9DDvQ9xWtnGbV+qup+aQGSvjfC8m3bGBVta1N
Hw0YfGYb/E/7ENEntkedE0tmkaFVqbPRcKcBMMGiQKvy4mylwKiqeXejX/CCpERQ
Ta/mVKsPPW5fDCjXHH7ZZLvNWWBm1sCnwhygllwJOuqgwT0B7bqvOpgtiBafVgWy
AIp6VyL+va1/EsEILA3eYdqZm/1u0CAxohLc6L2XdEHLxNUfnDh67lSAzI0Mq47g
3iHTasNJXHtIjxeah9soQD5+1SWWir3rus1hvqOsDlsauvFnMjCeVHUoJhBr/uO0
ZVZ+fyM+gajEE1ZU77LI4utqThl00TjVsGInHxRsWowCHtUURCMeyAMuBIMS2fa6
FWwN+ep23dXovmo2YHujHtbJJb4sWOetDJOQcfPltErmvjynwXS3N3i3RnimKl1G
LyiJta4Ptu6GoyhdvlgXsv7ATtmz6UcNpp4WX/NTk9WMFdYM8H4bMs067Tj0CClE
n3/ux5UOqyRn7Pg7qPySoTGNKxcAU7MXeORV1CR9WJd7WGYTm64pAyJqQR6vR3oR
yJpn+IIkT80Qi4Kg8k6qYAei8vBI3Xoy+RrT8AG0c3TndlBOFhNyH16g0Iizc8oo
201jJFHvQbTUyvVZQWe/xnOkOitenF7bz91htc78DXxngp3n2lkxVHKna5leRLtX
hXUmt6rDz0yy/Y6+bAbWfhMnJRg+5CEbwVEdXrd08mdYL18n0BHIgcmmfdAOo+97
frODqaTbkasLIc56DpTvqbsLlYlxTQvqb/49HS6PLZkrGVfGa9dTxKBOzlY0SmJ5
woHElx4tBMftRiZs/igOlSlqNbwayTmFKvBIuIRCsw1wXYjQLmQKMD+X2EWHcnXU
B6nvCRsZPInbt/F2ekkeSx4sjNQqdAGalxNdrl4n18rvZ3JrekirPGKIWr0ZZK+S
AjCdd1uZKbbq3ofQ3WCwDYEXj4UIcd9rpvjYQMIj9+0Uay6RInNaP11RAYJSqQ5q
e4sXiKY+Qp2n1/UhzWtwimHy/VjIH1RJ1yF37IJfuQ6INtCYcYvwyt2834WVmGlL
TydvKKey26wgerTrvrRbLUlSAQgNyLK0nTeamsw14jg1HBqrO+h7rwyIo/tUNYbk
PEyZ94FgvSjL/0xSmgwqG8HVrNuu3VxF64G7pwYsveKdkrfQUjDSe/fo5QCIziQG
HCaWmI83bNi5mQQucTPLOhAeK7f9w/3wcgxfBUFSOn8UXQKlEcB7W9oLJ0XROd4D
/GRTClyBF9NnGFXRys0/5xMOiM2Mw3jGcxuIxt8I24Xv9eHdohC9bTS7yh3QSo3v
2F1zvtOfzLq2rwSPavsVSqYextBE7QoVjdP7sXft0NOAGmXYN4TkG+vxmCTxfAXf
10Oor3Qk4Ew0dN9+mqCJw08ScLcKTsmM4Dw5dnHGJ8WggiiA+V1bPphC6OOsLQ1t
HiN2x2AlnbIHbPI0J7xNOiudg7Ja1W1ieA1fs1+HHzRkHGOV/TyPtKwsoz2Xp4eT
Yqy0LMNuLuIXoHMsXQ1TDHlNcG+DqMPizcnKZBZAKtQ6DjMIHxWrlsoh1lcC/6BC
mNwn7Q9w7Ik4Kk2v8iZjcuLM8d8E0/FomPWMnJiul9EwZbD8Yfo6HFdIa2ihwY1G
f9vMqz7Bs5ZmomhS/C7gsVle3o/1Vzq6H7WQHkd+9titkvgAlhO8KYIkOHDp0+Dr
J8mvpA1LMWQDQ6D32qlx2eTnwYPW4ueGCaEL5Hb19x0XRpGyrnMGM7IGyJCOYWPV
kGp/CrePTWu+7kGTMjLY1EN/whnSfVUSLXM+jv9mj+o86Qm/xakf41/Phk/FhXII
d75YiTss17A0nJsE/lV5R7eFu7W/9ARPaXlGoZQU9D0ZF+Z+HqUDIIAjdEp4U3w4
MlDNVYr2XuxCh6OUfcsX3s0rdhyoxpSZhQOWCa8XDt4YASXIQXlWyTYv3tQwtIA6
XtkzD9pCD3tMaApyhEDpypcJcAq+Y7QC6aGaPVq+hQ8PTlO878oDOKJrC3nqZ15j
jeaOYpgesK65lgUp+fkFhmRva7UEZgXnwU2F+OaLhBk2OnxaP4n/G4m8WYjl8U5W
98b/MaGg9UniCQHccvsep/KzKCneQBJqVJPcyJOqpAZkw2JhVInIsWpNGoEbYRS4
FZ00zd/BUeL3KGYPBxUUSJWuRieBu2UYjJaC7mBeun2LTPh0D7CrGncU0gRKgXiH
LPMyLFiOgTebU8OPIfKe3Xu2hQQZoDdJdA0M7yxlmCBRaTKaBt2wtVxOtUYY/kLh
vjeQNYQxuLv6kJpMlyLjXCTKyM7xMtjVlJeDjbqgiG0pL/lO7OLvsuyM4OUqBV00
6ln6Fhwlb33R85KUquktr4XeHsNAjBPS4Ar1ATgWNnZvRMaqTeIQUAhrb+nOJRkU
gCTj1feY2Vv4BAuhC8WlmCSaGGOzcLCBgDNOMiHD+K2wVO0vcmVAeM+J9VSlalf3
UFa1VItYX4jQfAndMBYyTbYIaUOYshyKKD6AizjufUDiw7d+ZhQrs7Uytzki41EU
JK6xtqmbLiA0NO3UtRuUvhFvvNZakVXqUr9aElURcP3PGRnTSjDYTwwXkzJOnaK5
Gk1ZxLRTDAu3DeN6F3CsK0L45mIDunj/rqgQJ2Sgs7uVJwh7CqEqejtsYUkDE5rP
6HsqTWxmzTIQ7IoR+6JRFkpx3ZlzoDsO264ZoD5/QfQjIbFvKyZnP9phk8ZfeqJZ
q7bEC48JWMrNCa5rBEdf3b0k+bCeBOINHY02n9lof5naAnE5908YY6VqJ3ZmleWV
C0KSnpruHZwXmC6I24SeoPBP9C2GLDaNkT98FGHHu/VPYmClnDcHbgD33HurX08H
OOGGZbP0CX/zJC1EjSxSODxN1rn02koO4KehB/SxnC8lkgwJM5opiN9zRHu0d6lz
GodjjkMv4pnboT7N6yYM7owviOY/CIgLdHuZY6wQYVOoxdxeHa/Ax3QE9uYTeBFR
T/UGAb92ryGvvYFqi+lmpulBnOiaIGpvz8f0VF6s6o1nf76U/5SBO3arbwb/Mpsl
I1vsteSeohGu7Fr3TMpW+zFEtaXX35BSUAVjIGAr++5oS6qo+Pvecn9bhTqhg7CH
TgdygZI5ErX/CVpQ4ZYTA0De21rQidMPMpED/ILAILt7SckNmoux3JKFqL5U9Gjp
dKPYYTngYg2qaJE6t6E4vRx1KBvcZqRmP1hvnk8ju6YxQR8KuPypxAiRGRAy9+vj
gvKOtMqw6W1//iBwFge80PvukXbXs0XjJ3rlowot6mFxcg7Bz7O409d4kb9VfACQ
c5dC92Y/xi8NuDoTfIScCMmTsVi8yNL1S6DDYXiYqD8tGvyjADMVMwabAK1wPtAP
x62E2O9ymXmTeEIIGuhRgqvHWOb4t7AI4Ymhk7oytaA7lJ+/SmuONT1hp/MBaTSr
Ujuxsw4Twh2AfOj57n5bFzIhaBeLtAQ0QfpuDsxyXNGXsYVrAu8MbJVrqC+/mAmK
zkkaIa4bnG7dlUm/728NdxX0BHMV4qkRk65repp2UwXB7+vyyiWnxPTrFnd7mxyM
eNV3GSsbA9lawnDKQ3URYJq9EbYz4sl/7KcXzDtUeGcCDnz1NeMcqmNLRgo0Gq5W
dMPFGE1aVh0ddr42Ph+qej1sjFf5om22N3uc8p4U3U4RqKOr8BIeMmB2uykVMYYV
7b3RrfANeP7sWbdRxmwJhlQruc8MOaS2LI8PuB0836GcSmdagaDbFF/k8Zyoc6lF
KZSmwZOJRcob5DGiidY+ybvKBhlNgvLqhva7rSD7Z02l6Mgst0P25iqKvHUqTkUD
OXZGP9aSSyUJJGNcgO6myzO8qjGUkpJGA53h9pfYJBCcS0qxkfsPDT9lW7ukIe+0
YAM1bWFGeCiUShhj8+iHfk3GZnbpUV9kUUcJDRVDjaaRevD3Pi903SFU/g37plfX
DE1PrE/pBCLHQwdH5ysFKKMtppZ1Qq3QG2VhyX/QDaZbCaAcJbYWJ6sGkbzU+umq
Jv1yCJTKufUIQk5CCE8b4l6/aiTVQ3DPlEEBGIC64D7QWsjRNzUOlJHvGdUF+Y+T
ynIM8jRgvkPAv5tInt+XfdnlbueV+OadsdYyrkK4koKAP3cWLq/7joWOIY2YhTU0
JGrSd7M5RP/cMHb5jMDFXBWMlLhiJ/wJxtUHy+ycepQ6cFRFxQzlyneyZKVViYaI
faoRZK071qgzMeRxa4xBvhP+J+xR2sik7W7OPwaXP5k9OOtWl4Bj1V2DcXvgT7o/
W9pzLOnY5K4Czcd6AGgVeUfe6TCBXnWUk2I+U7DWqHDCUtsdx62ldVVDQU/b2aCT
SQLWKM4RlT4xXoZrtdzdfLtLOUI8teCYU0b2UNNlJKKNXOgxpJOvX8c7CY9TZ3/b
PIPIOkM2aTDygWSmduiG0Hk5Sbt3m0AGG7VYUWE/qqjMd19SZSCpsHIvijld7Ma1
2Bo7O6YfdFJHN/hDtkHF58xG7viIgqDJTdOw6aMsqIgj+0KNBqW0aSTMs+RcgDit
5rHvY+y1J/6hCc1i0hLJYw4qHtia+OV8Z5AqFim8SPdwmHNxt/XC7vs5g6iovE2W
QfWHrLkqEc9jMKgxUx6gVjiLVhny2kOb4PpuVHtxxQDGjoQ9gDQ9pDbAOfAwkZz0
mlRMZC89dbj3LqqKDYBZS3Erjf+ZnjnGA5QIrLCDo9UTZLNv8GiwVj4fEnzzrDWW
oeds9KDq35uzSCiP7wKsqo5vjNxKodj9yAphWY0dG2V+2rrNxE8rDKJE1oANYlS/
ojmAP89b+EuEB4pguZYDNHSvwnLoL9q0Dec5C891xsue/xQtRYx6EICoK6+/a4At
W+7U/rKVZqliggYbKBhf4BsGqg6iDdAdMBOQ5vddIi+36QgN9Fme23nbq6rLdI3x
ARwEhJEXv36tFwtrdS9qWU6StUNiefUnK3hQgSNzXbGBxyLUNbSHFV8KnXeJF2Oz
6eFdxkH516AwYkK+4QX5h8tNRwneu8tPjOTIT+SnfQEca1FNl38rxTG0anBmV7qP
vDoYlHYBcBuzO5VFyFts1Owcc6pYFtbwAMA7S5BKn7UgWH8lGqopKwU2/Nt7o+h3
q67QmW9gthcpb1K7AzN7pDvUkTHW6yMgIgjr9dzwCj65GmKzpejugN1COjnDF5Zk
CeCIWUSyaWIufApW7JC8CABICt6ZVGHl4+TxUVHiDldVQ0Pr752fioxsEbPxmSGn
D+vtGrQY1BkDNQT2Q2C6j3TF5DwBNO0E34a2SxosAJO+HuQgjxwd5XI3LrKJMX38
kwse5SEcI0HSIHgCCQR2D7uorZrRqqC+HuYjQMdV9KuzsVDNecQM1+66uPIYRo+I
dGZKlo1tB6H0Xvj/kLSfk0jO96EsRLhRZHygidm4s/VCwmiyqutSDG8ZDwGQ4Uv8
kHULePJmCJ/sBZ6TKbNGDckARZnhHb66aZOmIOU3U14s1ZjFJMpxgO1A7FcZTq/Q
Y06Q2KBgonVcpoZyPs95pfZDwbP0f6mx0EQVMqdCmTI1UWrVq3fe77Lot3NodwFq
11B7ZniStdioc7UzVJQxCPu8krndpwINnEiwM47CaLeLGCGLYc0fmKD6oWDFKL39
y5d/d+C7cwpnlSlGyGJmhGqPlznT1VrDm1a7zQRoucUUfKhRV+vYEpuXo5dqJ8EM
NX+4uZ8QZUB4/a6+RDOGX6Krsyh3DE9c50KJCbHmx4SwHKe9SqurmzCqXJQigUHF
eQV39Uz8dWUG3Du+SKlvUS2qgHbpRoyvCbqAciNvGcfrJAM+6dl3Dp1DYjdSvRME
WXgfWQyjIEf+wIrCVJ4NOhD6UM68dUVChQnD6aMBFke95kKFhyoqV2YY7iTMFCnw
jNyTKZcMg5bv3TfSXumVirs2un1rbTZLk3+GHp/01LgIqjBv43MxD5mUgJIEvDdJ
31mHyULCcsHjm0FX3ZP4SdmUze5BVYW81jtT/x7QdQ9ufbxJ9+tYV/WeRmL9dzhI
25/08t8ovba1i1Dfvsxig41O2/P2T6s9iNLzlIfEYvOTQ/GOAh9QEV5xoKCoJGmx
n/LaH0q2qJ8MvFx0B605sypbX9xf1nf/tE0U5Ts6i43QOmx3jm6pCoUVVSmBIvB8
pGW4WN8AjDKY8YUhoJJh8rhHmLMP8WYWYY1zSH22LOXBnaAgq39jcgXGLvRK6Umb
nnDBbKVRENm3Zq57NEvw4x+F97HPu7bsNsY7sQ6cIwX+oG9c+4xSeKUiB9GQgbPH
FXmG3upwqu9fpe6/R8uYM3Zb3do7ke0L/hSXuVYbnqiil0g6r6CSKlyFTjXg1873
mb7uufiBuHbw/vDIFLQjCzbtojMollHMTCU1FlnERQo0fFeAVPZmtLDe7svtOHx4
wuXeb2P6qLHU/y9kZ6GseefJq9uhEiOpfv+BDj5DjrC8p10yD1gBCfT3iM32oLDh
Pgk9oUX/ozb7e+51Sj1EpUF4WWjlpc46HUznX95oPf8+vRBoeaWeRlXmD5k8uS9q
sVdf1/cuNXcJeAi6EI6en4JJvSV/OBW/Yc7OjWFQ3+5ay887ZtUa/VdqDnJumZYh
1Xkalis5rruE8yRUWOigwErC8Q67fvR+Q/XwagIlOUaKXc4RgVH8R5VuAjVf+RhP
2yONaXHKXpymdT5cILVsOGaac+U+8VuiLrTl9QqYwidkEUXF8T580fDaOxreBeEB
XUQEgPQGuljFp4sFSJF/cviSr7UanEuZAxY00Ary0nSd0EOicUOXUp1D1H2RyIxX
1LhH/i+MCuGifimvEWvIY5qYjg/jYywGh5Au+G+b0EaP5CuZ9AHfhj4lGf6eWwBe
U8xCbeDcDeV6jVFVM9LW65srDUUo2TnjLSw+gr5AfMCq9n3b6oTPAgRuQdTrxDgc
xC2AItXZMCgkA5PR8h6gwnvmM3fbUhw8/dhoakph32Ab5ieg4L3fbcCi2uQfP9tr
8JXV16JCZg8MIYsnRPpEh/ZNLQxfYqmlD6Ltn/OWKMU4VWE3p+30XwPd4tS/6YyZ
d04wuQ+COjw6P4XplXJw0rWR3eHFwWGuNL/TefIp8+vmssmSw3wo60Tx0roxL4nb
LvhmXfY7hj/HG64mkZ6CdXEr66+9IKVJjtuDOv9IjFlcfyHbNwjGt23pCalFP1NU
yhjpJ0ezdQr3riCO2tPgeYc0TWOF8eX/L+R2R/kXl9M1u0IeONMf3C+Plavm3V28
2/RkxJlFdPds9UsShygTr0qgdn+hu/Dul6bKtbNvIypKnAemuRtvlElua3orvB/T
xk3bMkvjpG54mwkl0mYbXtjDsGP0eDylXcS1xn1muvZEVyWzoYPK5E4uhWmaEcc+
QUFtBuQHrjudzhQG1wNfWEWHHiNBajSnzKEKpQ9Vz5gLQQQ3L0GBTtMzh19Q/e+Y
M1aqmYD4KOWbzVasxHzor3nXDRp3NAft7u4LPnKs+mLujOvtXR1BjP6/8Mftxou8
0tmEa1jtdhTDPRBKSAhhKAs4UWFJp/u/j4Z2y3kcYY47xcAMaq0PEBiWs9/jXOhU
h7VUe5f+861CPvmB9aDH4okFLVNinGobmoffcFaSiYVr5WMTVoWUuVrXf+x2rrgv
m3I73srCJzNaDhibDRPqQakgFfu1H/a8LX8G22xmTrC1FPJ6cWPvpNnsEbrzqdx1
JdPN6rSjsn6bWhnqGbb2CgdwR3tMiRttHp3L4t6rO+jxY286K2kT0KCy36kaGNFo
ef0OsQiycCGJnXG/SnacuwHbA43ouR+ASXwgYbTxHnoHRmJCwO0GuJmH3uhOP4EB
KOvKbbHFAN2Hysa2ZNE6v36wOpkZecy2OXL1b0IZJ6RHoQkuTDRb4WvNUP9+d4+w
k9vQ050tYWDOMp2lI7OGes2lN2oQ49mgjBy+XnBAQMX/Z3+XLZrD5xT9rkKHwm1L
zcUwJVXI22motr8Tdg+y4pQIrlU7fGAhY3j0F2U7P02iI9aqXtfsuMb2Us4lR4gf
9InajJQAvmaG0o2+/NUUT903OkavSYhvFyO/rQA3wZN7FtFI6AeNg1K8w/r3QWcf
WlMezm3N/RWPcgzwpuxY73MMdCBPO9lZVOcyn2CgPDrcsYvcvBVWQiqQtFUteHzn
Su8kltrsNF7/OVUj8nDw7yFaNiPNLLGGYL8Ns+pLkKrA7yiOpNkGm8fUveFa4iJI
XsSh8CvXYUpZfzPwYeyVOgMru7sdST4AzTicdLAzuOnS8VpK/ehH2bDu1r3tNLOr
luG9sNeNWEl0rvYl0d7vzA46NiAx16RuB5lgYLBypL8o4kvFb5K+6hyOo0OB4LdA
cz7JeI6OyfHI/lZx/59EdYiM2k//tnV0/5tSq3Itf9cA9yLYFN9wK57JteDBi5cT
9gHHsT5S8td+IDplDC9qbpWDx+T4LruqYwc5nv/gH/8jHZosibNdUKlYFMP2jjBI
Nj4VfKaMlfc/2yxvkM9W4fCBDSNWqDUYKs7nLKVe+TKH66m1RR1UTaZX0OfatzGy
fyCNTDPMcDjZvpVHiP6N/+sEz9qU2dBaKWJoihe7fDAIxpcCiaTkJ6Za7FotMkxs
C78tBsVkmP1xUM2aoIMi+mgUmEsmf76GyayV65IgS5J7Io1XUbrLELl1XjI+6dIn
WkfWDL8mPJBeoXlvByO3t4FWxVbmrWJ31ytHfGE5lf1LWnob6iO9RAARNSnA+xJN
DOJ6nigBDMCmCIG+HqiqFunAr51H4kdJ+nQbL1I++TLC5DQX4cEAo7pxQkVXXFAT
3W8rkiDLGxoru49WbMNTr29LMQ4GHiNruzXGsXoEogG6rnFITusn8LJEf5WLpwww
CxAUiWlXkW1ydTUdz4CkN3rmnhfMNw8nMKPHOI9YmFWcL1kq0VSUx7chFdyYwN9u
b+mL71m/ZYF++V/p69k6tH8J6HByMsY2YI5PwPluKm2D+mUWOv87PR/WHl+6gBOn
nqOCAZ4Duw15NnkH/6oznIs1ef0uzyHolYYt8xm/DjukChTLkZXjRFcq1Wv65+jU
wNxfYvixH+cjrEylvjn1ZUMY6UIWZ2Mpd3TO9Z6q4mL4M0IY14AsiVYSK6F4YpGD
h6QhE4Wf0iO+nyrI9K4MwXtup8hEj/P6CbKgV+GMxGmwjkiXa0jZ++2NVh+USilK
1SjEKYyX1ld5UBrciOGFuiT89gi0UKd9ahvpfqdGsz6c8a/v+Emd4go+aUW87VLA
+FDhuny9PtR8y/SCqrPbj2fKpjqpoUddFgSBNPbHfdofzJ8avw2q3rQKQIwIUtUc
6ZwQkORtU7GjIqFXI7qKNYrxwHLjMhXXDY0VXI9AJ+ycP5DXabQnzQykDe8qpjET
M+hAIjf5D69RTBmkdPCeJZmbG8f/cfJTAbEe4Nm66iTA4qxXcnOHEA0439tCYVZa
NcWpRj5jUGikWIqQsLF6syOYgwOtScxWsr7vu/kaus+M/eMB3GvsvZYSHaX8U4eG
prg26MOB71sCL009Ilu8/GhBHOfYNlIxdmr+G7tBxfzylfbgNaRC2zFxjed/r5/z
cTqHnRtfBZCePnBYgVWYDMuqEQieSfn89bblLBS2hWuW//1oV6XkvTSwc4FN2VHj
2yrw2Erg6jfWMOgloE5iRHZfgjOrmklBml28jHwh6Zm6hh8F7qm4sloEu7XCQRI3
XCfMCATakBvtohiFs9LF+Zt3XFYm2WEqwnIIrj+EwJhtl8CHEOYuyrpbbfRKRk7j
1+NOCU8lW939PiuFotGI50lziKdafnLClg3cgnzfi7ttC8Le4sDqo5KvPVuiXgWE
W6HEBYNXgmjQXGDNnbvE2DEApHoOl4Wo1sk9wemzvjqiYEQNzJqxisgfThcl8urk
DLZyenjAR5Wi3Fb7gGSEFvp9oHXGzkLGj0sRAqdX/92rxqtaSXZVSE8ZUiCZWdYv
tEGuVgykeA5T20QYjjE2WV8t2IJ4SMOBofac6D9EdAcbpG5dGbAO7ie1jTCjmSXn
ARJ1vR1TROqe2cGW2kUuxeUHkst1nuPiFa9jG6DxiQABBktcsoagtS+E7jW4+ymq
sxQZCXrEns0FCUpu2ROkYyBuQDrLQqIw5kAlM7YvN06Q35coi2UgIOiRR0A+fLEP
XYn7OFUlacmMkUzRdQjmZNVFhSenm3c3ds1CwCq8Ury2PdOH9fDpdVvYqXv1V+o3
nChbYyiiamradozvCzpfl1a9Ey2yz+fK7PRJcuRQg89Y8m0Ff5KsNAI8ND7PXkZf
GaCfXKmPVcd8wrjpJOmvmfHIFylNwrl3etd0f4eSIIDPcg3q0GPYLALsaKzbUn7f
ef2gdT6br2GlStWaABOavcIcWssDnbeS5u1nytlvpsc/Lai/5omOdOBrEjeALul5
C31UjyumZtnaiS3f0SgoxI+OQYJEziJ+Ap6ryNMFFSARi4I/cmSSexjnQUXF4M6u
pVd7XXhafqPdlquejH5jI9ZBMbJXv0kL+wvBjysff3UCGBm1fP+i6dk/rFTKidsA
jhHaRoLdia58mFojKuLDTBax9SOT5MB3fmBhTsaDvuB6peZZ/xA7RXBT6sSjykpU
DS6wvZqFKldyrV5K6y6gQ0+ivzxpscOp5Xou4QjbZW90U+vVbxSP7gTJr1OtiwJA
S6EuhDYIiqG9yxJaVrbm736OFSb9IHdpvtPo3vOra/F+/810alF3ql+dOuItCGXz
A0opueqHTXgBewI8Ai32S8UDQHH8l4GI9hmfvyA1zEcWEQxWlUavdpdp5jbaYCgn
EBfuIhfGy2q75dVXtpG7Dsjp6tdDYdG3ZQJ7OiMqvWfS0Kzw5sN1EV+SKW51M8ci
J249TR67SqEVX2SfiEk8DPuHyu0E3xVpqp0L8vSDUo1Bb/MH2cgUNFK3Duy9LWQq
J7Ow/gPnmPj+vRBydjzInTxXdMe+cu0HUoHGIJelKxl3KdLHdZ42e2GCvfAv1ioN
NVb2O0UEPG45wy6mOQg1chgw0UMPdLxBkCDc+MXNQMfZtxbpT1EbmwNR7HUtObAi
FPqy7DFArAqYmEA1Wvopa4QbkJLizUqpKUYEMpdZ9Ge5t+gYYBaOdsC3/2f4h9Yq
nf+NqLh2CnKQOe9HraqDT4De8b9+ra8cx6148zdWpw9YG8nBfCrWjheHAFWN/nyd
lq9O+C4dS4k5RBixvPnl1jbjdQr0gZdtEZXqhiQPszBEWA9xNUEHl/7OcDRNJ3vV
0FvU/ag8CZH3i3alYiug8Gflh1ku8gM624jNbmwfH3irpsGQG98j8hM7FHC+3QJr
S5VdJl49sGS7vlYa5cMZ24VrPFAST27alv0CmkTZTdUpWXzo2k/hyyLsdBzWT7+c
dhfL6P+XlTQWzk/O7uQvkj4VKOy4Rdl8ofU8DQ+Ha4Wfn7Am+1gv2VEkB4GjuzpS
MVoJ5MbGdUsEt4gyD9RKcheMR6/TGfhA29Sn2ADioKGbXgUha8KxVZAyZHs14zHy
OghHBJN7d6GHHPiDlaIqJhTcxZL8bV4fib3HuLYvp0DqsMXbOEaYzraF44HlEK7r
3SLRmjzZo88sTWC0jpuHCiFVSgt7gAMkiTz0hczkjojPMetdLgo1T1j+o9KR69hz
7D7opeoHBcucknUs4pFwxp6TGqtfSz1eXPCMjIz6B1hGxTWkG2dvAvZbD5cBT5jZ
UWOAsAD5MyqDOFlAt94HqSNDdLArmxJGG/WD0NQ7Uarbzb2pp4A4TWHu04ujyDW4
k7Q1PlmT593rhIIxX0Jx9v6hDxC8YgPGNQSJVM+ZkqMDFG8AebCIg3/vzlMcOb0m
/o15rVD8fBZZSR+dOXcAJgFu4N4vSIfYbzSwrYJrS9gLTJu6Z0GxtyHsvpnl9TLA
Ugb+3dtk1cTg/qvQaMVhFxRA4EPgngLnLJ5BUgL4oHVQhRehI/tvEEiFl0q07p7K
OTGmOxff/rYlMhrfC2oCayK7qYgCF6/ymYjOJYG9p7hIhI+hHMXsMJRmxR9XvfTz
bh93Hx1JA01TYCr87IHcaVRfMSBXsJLfu3JTCUwrJdgiHwActsLvkqmVezMln4yA
qHHADZf68arv8GfzKUPaac295IZDjryIxoM0v/KOuAHjrdeUqvEgV7kVG7tuBxcA
Vmv6xaE4cno4EZnOFoR8HXqzzSBZPs9zlcIc6XazZoy2UKAtKa54Y2ZkzF3XuODM
0H5sgf/0KujctQdSIf9kzeMMZrZiEz75wyQVBJJorC6r/s7HEFLB69so1bOaaro2
f/YFYLZyefUBGSvX403uQGEENijhYc0QHM2pDHkYRwaItuNZw6V4AjSDEFSfvO6K
ycq19YdLH3wPodLI5XajtEKjozjugbwURzDfeXOkf9DMlHZCKHduchiwwM5l9jvM
PCy8+3m1JhrMQRfRWC7/ej5v5sxYZrjwCIUraWPxto/2SspEWQxdPNuyJN3bbbDL
xrpCZi9+nwBj+VVMoHz1yBF43y/LqSki0kL9mOGxDIoKVfHJabOEb3HZCLzgy6bl
nyxeJHfU1cjw2VG49EumY6/SjWD+7v+3tyyfOncELIiwWXz+RFhiCS7d6EBBIdx3
2DpGfft+dBqSYN5e/Kmr6i+Aaysb98dVYI04e9BgwuQiHbcPMAauV9qP94TWCmY9
aNYboVF3FrgOBDxv+HHaiRmLJndj1FqfCqEK3+turNUabutTLCmK+dYoJ9FZCd0b
SFxKcLt+oVhagxysYIVitOAYvnirpsziJ6/jGpXs+Wc=
`protect end_protected