`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6848 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
dnVBOIGMhMFpJZXzCENQ2LXT3Ei+gkK7Vh7yW3iIwkQFJrkh0xAaVFZ5/DzGD/Un
rSv+Oh1xqJuQLklPs7/FJHcQOlH3c4yTkuKc8m1U5tTtEwSCNV4EPZyC7QEy2VZd
L3Syd04HIYQaop8ft8cv9+pwNO4lzP2h5xIMRUrwuMo576PX2zKZL2z11Jz/hCmm
9jG6epPc2Lnfu0L/VyqQXY0c8BOiesrdeqYRP+Mpbo6MhA5zhT5pwdzINn8pHxv+
fZJzp9pX6vohHswlGwqLgltdkuTrWwgTBW/u6NuEoCG/u65jmI+xZT/sYCYt3Ktx
pbsZy85rAoFvwKsqPG8zpEYbwg6y9Oa6zY9Yj6S8P0H1Fi7+G4XaIjn+ltrNzEf3
C2dnGMFdw+HD+fPL/NpjniuAnEdAZRiMhtq7pntYJ1pLxDb/S9jBHxEHh2WWiREj
/xOvX//bikxT3fwe6EbA/vYKfxy/59ro/nQ88O0Jwp79EzsjZnawcKUzJn/DqpdA
TrbFJJD2pBuaOTd5OUXBxn8L8VNmTh/31jpJ1ez98hw9CKJTxf0qxonWXVwRtSr7
WIy4qu6C+xCTYMzV3hBEXVynmRx00fg9ISHwYDFc/VTZBwuLlaf6flfcNk6Ro/QB
54YtGW+QatzhqlUmYSxFb/enjLiXut8/puH4hKxKc4wKfqpQwahCgRjq5hQ3R1ZY
UEaJPzAXU5WgTTWmrfBEK6SwxBlEkLSe2hKpd+0BN0TUzbk7iV5Wt5rs7rbv6m5F
hm+CSMLxz8UgyRwVS28NyPi8dqtt0k766Q6OKAQMCowREO4HISbK1kQoFm1GvIkO
mJXuXUL0brYOAlKVDMp8gkiZtRJjHUDwnaHTSN5CUPmOisdkVc1h3n6SPjMlCy9w
4FDUQJwKzZEYDC9ONSxWCgrZqfN1wR9ajGRMZRpZ3wcIZ644z9FYT0oD9n9rak9A
E1iLmppKbS3F0738G2ppE71L8fjDwPbB98m6qd2P2xOV1iGHNifYrylPhdDc6+6Z
0ZvQSxiRsLQKwQhM0bKYa8CiIZNNb2JPiYa07VN6vYT77Snjx0MCqgyDr5ZGc4yx
j3CeQ00xjgoxmNLfLpDaz2iO8378GYsZIRqSpRAGKcr2G0X3qhbke3+Tsj9CGKeT
3A9NiMhyfqiOtmr/E7r32/JdyYptoy6lmw8Is8g2lsQw26H1xAK0S++JXf/aH8OS
6/cWQYPwsrtT/LbM1Io4danmk2dSEn1P8is0TMU1aF+K/5rbeyUpKVoh38Gmiteb
pJ7U8M5QShedH5Ocgi6dB8mujtdPcxMl3DvV6TEMflMkRL79DPFlJl+AogTgs1Oh
k8KEkT296cRUEdEEqmHdxtBhioYzWj8qkj8ZndiYQ4muRixUmCoCV3FkfpxP1/nT
UnwMAn4MecbDzHdPofCRlMukIch8h4gboe38qS0g93W6yAW4FpQxCcfI+8F/Ivhf
I/ZTyKSVdo9/ewKppk790rsPuYGSgd3+jFW/QF3hOjaMdaHMYgC7n0fgzmAvpZ7L
QPHCG242aL6QS741flrKkHwD8Lop3fcKJiqsn0QABDWyOFp0jBRdbxYEVF3I7TZR
FsCItNto9zLMc3tc76WgJm3WB6tgOv669edzPXNUFTTMfZBTBvQHU36tvL8Hkgnv
OVG2jCm12Uydah2ZUHR7lX/ZRsj99s3IuXe+2IrNBhluQzX6tUpH5SPUi7jSAX4M
jiFXMFVaiLXVPjA9Px4OdN/oyPYBNEVY9KRiK5AF3JSO5+9L9pR6e2wuGxgmsm/D
ohB80r2+Pm+rdw8tBdRaPeH5jdRZbgi7nr0IBobE0J8S1MQpZfQYN3skn58efK/x
aX9RyN9SaEXe/mb/Vj2aXfIygck/l0YY2pD25gJNj5/9Nxr//M+e1WKPEjdK9rnx
BlGv5B/2kmDSWEWKwtRk4DMK1R/xmMU62IMlz3UFARPNwmh5oaQhbBoNWgITgHx5
rXX7JQA8a++xICZT19JnXhVJRxEVF6TAkjSYC5aEBXccwlD0jyXvdxIDfihB4D8f
LwrVeEuwfdLQvgXH4mmjTOz8AssNafgeDIZFLJeg3Zgv2xlhzQDFruz0VsGopUa6
M3iPdGrndw63N7WXzoGBqJjvtcM5U0r2yK1l8aR4LBl7S/uWxhd0ZyobMB7tA/T6
nTJmbBOJo2hhpNyjBfl+tK7aiWVUChp9I5dinOe70y129G7zZlir0sPghkJcpePo
2Dr8jEY855iCUYBIP7t+Zh9+hQQsqsvAJxI+FViF7Ph680M9TuA5NPQu+8Ld72aw
ffJ1o/LfERnlaIZttZGfTiXs6aDyKok+9aXpEagOY0AwHHKdztmYzcTzZe/xOKuX
gFe5LO65pwLKjwvDRCVPwebvwk69QEEyJLJv5hJmvqFi8p2R1PVspwfmRetwckGu
D5dOdoMml/jj1kl92La7e5q7XiQ+eTjz0bR+9lMYEX4ROMHwUzS0YVt7jDPFpNfX
iggXxFMDMDilujQMZRxfqR/F/EGdyb629PgNcJD1KTq8vHsOcqz5eF/8BoxjBL84
/urm91qCA4cCWbCDHrC34UPjMQRkMVzmiCZe1IN+Ft19UEt54qNsDrtbXf0FB5wB
SZcM76rCXMK6ZY//u8Jy7fWeMNJlXWNnJw3mAr9C6NEbBptvjlUMc1WjkSsE6Mhp
hVJQKw15+fmsLTIyYteruq+Bqr9BCxD/4BLZuIiwgTQtUw4BzWWsEhO4U7RnozUk
cAgcBNFBIMG9PqNdDAaorVLaqHqyx12aSycG4GTfP5Xcb/pb2FIV0UWzOmhdx1oz
4CS/UonOEtSHz8i0Sl3Tkg4odJZWk2BW7oyFsq9Si8bI+CsAVJKUj2YeMZ3yIKjr
BDCUGp7BfRGwifpEAAveXCxSdSOBN21uJ1oij30EQpsfCv5WIlQ/+3GQTf3SNE+D
aOF8gcJbQ8zNgk+dVe2lvy81TdcU3P8Seu4C0Uce35slv0Dc+lNCgnZ+psBhgYPp
YXYWZ3lskn5e6SK14K+lyZa/pVx/MY7TZO5kI65/0d3z4TfBA7R9ax3IhgKVm5fJ
QJCnp4XpiENm1t11cfbJl3NFdUrwPOzF2wHWCrduljIudmF0Yc7e+sIOzEXNMH/j
UVBwLkc3vPW3PLdXmM2cprBEbvbPde+thrnOY5ryLxxTihHAncJogWTyaAQhZeLN
gOMU0++OxB+Th9aXFqx9Zj91RuUS6P/69R4gFVt+Wvke+GDJnR2TRv1X54VWzsT3
G84keKkCpGjqHDO/K3xJXHqRNH9CF2nW5RdnyEwdnfF4LtJAdew22GClcnFH4Hur
1QoIDAbMh3gZLYu2FfeDRg1UWS1K8u7NPq5ONsXwgiA9Ydnaps25TXiTbRatqv6m
QVsr2evI7HqhiQ1yU6X2XQ6urX3Ep1RilHxHHj0u8lHU5xfccy+WMIJmT5fMFWLx
CZcaxTEYLg1pwkQ6UOUPPkQjM/2y5x7O1TpQXLvXhEZKSBejq7FJ8eU/os0+aiwA
fp55EBeVyPVkkBUmu6l6zMzRwoF0+TdoN6VhxWqoj9yL3zCHcvb6pquDkG0sc938
1QovGc1uzWRE9L7xfsAE55mGLTVVG1BcQecJZESswLHZQu0MngdIhVpaguLdHDnD
w5+urV66j1eM2+vFYO9zzMBqJ8PCtATz9ru9Y79B63CFtQGm9Wnk+OO9JgfHyYwW
aaTeODk5lfUQtF5i+3fIcXbUX9RWV4YDeyYHmANRyvNSes3cTgIgV5VCKcZ0C07j
1AAVTeo3ySkVND+s3WEyVypiAvuI7wsXWLf1ks40GTzirS/lv6qd4yJmkqgvykbo
IiwVo71vG3bTVGqWzzO5peLcrLCZw+gEl5XUdfZeuyJbOB3QRNTFx9yLOEF73Z5n
xp8sTW53a78fC3AcsTJ1+UEJacbD+flGN7t98D/ga7SKj/maYZdNdnbJe3UubVHO
y9uWW2IqUsMHeVFy2KJYUHd2PSB/iJnZoX7WlbtL2+4fubSdCHCI5YI3zLmUff0L
uGaqkHfNzpU0Gp957aacM38bJ0pWMpDGX6tdLajoJ/U5D7YXpBK5vtP6uZnNFoNL
uV5kgpCqdxE8UzdU3Hrl952M9xmxmy46P5lowoin+wSEXIQXeKtiaWXIiJlabKJt
MON56koR15mYBqPc0WQfipICng8z45oHIHTAOklZHDHNcPf4AMMJVx2HKGSrWIkr
wpLP+H1y9pNm4Py81rWLkxaUV/hWO0F6S0acUjr12L6BxR6MWdP0HazqM02AThrv
kz6f6xjy/b/huvkqgi/K6BMvtjteTafD477yX/CE2gPU1+/fgmjgdrfc0gMALT+C
GCUXt2eTDTYqxbpQqiWRaubm4j4Enjcc3AY4ZJohH8wMIdhcbcjU8i1HnYHXncMn
fmjisInbxAXuTZzlNc1sbOgn+FOlzNOBKMjYv26RYzqfzMFe/M2RcL0bshH9iJV3
3+8zUtO5mpLEtDG0yKbaL8sWwIu0fICAZXBsrceYVyv/t9b1q5UzoxYAuBNmWS3J
j1hyGTiMELA2y3tMbbSlifzO+xZfRBlvaJ/+t4AX2r9nEJpeqTBJ9YEUJnVexVnS
rOFY61fJZHSK8EjA0Oz/bwRmReDusd2ec7sWbSNYGLsTvKOE8ja+YWnfYLfIssxv
szfwkzAYAf17ydwzmBEoeVrPQtI11Pm63YxE702foEkGrbD6DAdcoo0AdTpvhNcP
9usetqOeQlE7EgX8pdJ++oSMw+cItFckLN0teThpVuXbin1Stu7nH6xu/OhhDWed
MXFAzuySA7UzBx2wAB9CVhK8WBjOlTeQ/kEkbxQBONauoWS42YnabI63EX+FIUzV
4kvE14L8pim00W92jKhOIh+fqjUHTHBjqOnl/40m7qTJm7S/sx0IAFQh1DyfqJ8M
MrreFYKGjtJYAJTR3HbNgxeByS5XzXUBEkbh6FzGEZK1b61TjtIrhnBGbYuBUSuY
n8IINhz0eKMroqcEevZRvVYr0b7c4E37Nb3M3tNCe604SZZje2sE6BMix8Xhr7Xy
aptuGbUEjH92/8umlc/NVJBEJXvlpT+iH+VUvQa4m4qxzSx9ZJWTG5P9unFVNXKu
2yLsjOPY/PJkbqrO3jyP9oSJB+0k5aFyqmYfrUg1x6uOKZM06stEPhugHOOTn7tz
TZDZmcnPCb+pnFG4ESIZJ9heIeF/QzIytZu2c82bxCpZwUCWHSIP6/6yuN7+kd8j
XMuJl+nh3RkPvmZ1Ef1alIF/F6BzJS2C1gu4Vksvm6M9+d6xs4p54qw6IqMV7JpX
00PU/1u8/SVLUSJWNlgY2KnmNERBIqV8/tkG8R8JyAXs6AvFdbw0Y8ZwUGfzWMNF
rDXvXQNFvdqmqNd/vVtqRPFV5tCOBf3u+alWpyBRZKlEKUzwdI8z7FpHzz7mZJGQ
uvezwhF/suzDEXGIGz3m/34xt7rko4ZVxeMoOXgfILOBUK8nTrQ3jzenZGLFwn+q
+Ihzj2oF/Xn3vCy2z/ypbfbEN8pAYvMaUsO27JEf0bgkvp3qiZbqexmtWcEZ4xsP
47okGRfV+fpy9j1fgrHwzoWPanMqe1mWRnrSryNDOGQjs6qDq/sON2Sk8fxoNSdD
8omp9gPKId2Ef5yjn+Et15jNUdBlRCtpoJB/0/IIA6JCVN0XexPcuQz/XQtoLndJ
m/BgzQD/cN2sUs5Rh4YgiT07XIL92nNaqsN0Ddlslq4IUoQCdrU9TUo/jsmMCzpw
RjElO2ufT6kVo+GyZ+T2pErSHKuM2KP+df09pWxMeuFOb+It/mCmTeACdnM5Tjj1
yjeSxBw14pho+MWSAYcTt39w/MJ9FetzdIc2cSJb4WystqUXo0vmcvQ/+jiHvgUk
ddkNmL/TKZ1hTPEBluPyqkQjJUy5B/Ut7iyv6wA+kXH0G9YwZBegAO66MjmheQir
rids3RlVOB9Pn94Mo9DtknaBTdAZrGxxnjhruhXKN6rDS5n5WUplaKn9M5eZzxuf
xKChtHKgpNSj/Qy4Nk1iVV32r7+eQKVOTcACovyRnfJ+6sh9Kf6HZj6A0HYxL76e
qfycEDEQUm+rgNIiv94lCXL365t4azmFJQ6ORCyUxKeJLY+sZnD04wOsAO1d48UQ
+7HtbNmf6A+VrsBa7fmpWZQyM38rSdnsnj2CqQhi0Hratb8z3fhZDwxZJ6oB3+7p
304VkoQhgR05k3WImkIjDpjRknQSk+Iz4Gfvj8xCkzJHT2k+R3ATwhT6azGwMnUR
0qAdvh7AmP2RW6PzdT1L0NQ7lyP9gpYjD3b3XDwKbhXM7aOCoib1sczPXXuO8Bwv
+LxIPPTTuQRhLlMeql8hzQPoRXudmV20nyNAwwbBoQILvjhvSsm87g/tEDAlQnT7
XOhQ65o+pyptV/iu0oENkSKcf8AUWycZlpo0oqAnM268UYpnVLPrW4uNfOhKqXZb
W9/EqvFmlSqqizEJyMb9AQicyPtqcyodwbdDGDS57sUt/09XAUfLiufkUuDtbOzB
+QRsGrAKPdat73sjHtGEtJYGezkppOjfaW0r18bGYQpCKnCkqtJG3Zvl4Ngbe89Z
NWHrFxJlQce+mxNU3+OhL+eVe2WP0z/Lp8ixA86HLt58gnm1q36SO/Wjdr6E3/47
gobDE9nba2rnnTPjN6h4/Gt3sNcqigIT4hLj6IGeSPlms9JbZ7mw3OMvM6M/PGrU
DowZ8ybreUAI2pCNrfH6jE3C+TusQumuK/NTTnDrKNRmsGB5yCsNSjHE7hi87RVl
Cxaa0YZfRpezXagBkYDGWQMsD8zcabseQ5gjPMHjEYcSvJTJPk1EBmITUYB2ObTp
zhIs9K+1lkRnNN5TWdOlugyqVR/PyJWHWWwM4sTCdmbhCYc0wOngPYw3kUFZKD8l
W+zUZW4iDsOGWmkElXPmpMz7v4uCgEObmEUZCMV/n5zIp3GesZBpdL2laixuCtky
NqHUybC8qpValEwGT90pfhP94VdSN3BYkD69wdr6RGUGt0ghMevZvSH5jPnnX56c
MRIH8OwRtLVtG2h7l9lRQdWcZ8Hfz++g1FS2n7/JLMgkBc+8zPqt49ytU+2dOg0h
91GhLJlmu6XEk9QZ31Gt4ruOZHCxC1+/4BTjAcRcz/CZRIDrbmyBN+8mn2OJ9PYT
HXl7KkvfR2Byba9zhgzITfGi2/iG7bBXvnEyLxOQYT/1WIJhHZccnKg6M56ZSFCA
plS5cAXw7eeRi2xqJAwSwtYfqNks7CeZQ8LpEXBv03AKFPfMkoXVO8oW6jCKDhJq
OLWoMSckZ4V2T7+U9GADe2pza0VdHFmlTUIoayhEyx0LRBHW3lCmK/ZiCX7hRlUr
Fr9KsO0c4owKrD/y0ysaOcet/3bjVXG3GGK0Shi7z+ai7M9AHTVDXZ8ZxeIZG7DF
agO8JTOtzgPEi8lOXGIA1GIR4jxwnsa/o07bTs3bjkUjGDeLrriw7Apk99ZIPEtI
G7endiGxNM/w8Q2NW7T6EkMwxEga8AKqduqZHfUe86jo2k9Ai9x6uy5jtZL0SRwy
At7933VWM1lgR7G139uTidtdIjsEX6QMpvMywMXX8luKGsHyGXAjxtmhqE7F4KeN
sM52CZDf5CSMj1ag80rzCbD89ESGODy6XJEg8oCdp85HB6a9ePSsUUxy4IpKebov
CNUJGvo4HnZ52UOeAa6XQlUju3iah+W6zSpcIxbVVvM+t0qnOj3KWpVxsa8JedlZ
5Sj8C14/kD4Y3h7WMsupSFA5NSjDlXjWtDDh8pQXFwCtTpW8+AZL+PB9m/IIdJJm
DZQjk3bI9iZvEFKSL/PDt7DkhiJGRhtCKtHX7kJ8tl8tdcDGqImjO+hhk2G172Xz
GRwzn6H7+DYwCPGQA8hobTGqakpd49qRLiGHS3Icfr6PciAHw1Tk4j3Z1Wqlz9K7
ojFKpdEHMVbReJPKs5OM93h6UCk8RsDSIVFKJtU/EsDNGIN6fn6s7C3BfmEzY0Fe
donztEDHUY92AuTLql+PuWK/PA4MV3HeyP9TSmQTfj2/UvGa/2SlaJM2tOpT8Xgp
tu4ZVF1R/KSN2gc7fwDCDKDSYSdjQK8T9B1PdD4lNplRl9gyAVrVDgAWFgUEvTD7
0L5Le67Z4xWzxXZcw+oMfUQsCx1E8uWu75xaJe3fgq8NRYnhBCyeiCYOt9I0W6HH
Li1qXP4CFhERXlYERA/UxVszp7sVzxf5rmWddfyqzx1mCs+p/4WpoHXeaLy1vW7G
vhx1f736exsqih2ZaMIm+3VuMjqd/wwIZaQpihRFso1i3BS9YytyH9nM897rbaAZ
+tquo9SzHAde+EuPX401mLoEJE5YYGVrGC8CxCHotVLetIwVrpJ8HNKE6T05tIID
YvVcxSyHxS1WnMYa8sYW7KJg7mlquJ7Ha7URVLTKl2jcz/JVEx2fK4ChBAyabrSs
oKQGRXqgJLOP/Ay/bcqY9trJZUOyn6XuuuO/k03YqWgDNkKl0n5HfCKaCCc48vzk
zAit8EiQbOhxwedg9xokxe1OYGsjYl4WgETR6zlGUUFDiDdo+DanCGhrNpc5kyNW
IttUkSbu0yRbZcJJ3ylcLzI3uRim0FuzG9nfJjoqBD1Wfh9zt+UNiJ6G4HxYzoOy
EresC7APE0XVGiq2weh/QT4GCQ5MU9NThFExCzdC5+fxH+smAAyDqIowkTCmQf8t
LzC3c2FT42HhxdK9hX5wklYjtHZtAzvxvTKEJRC4o0EzL6WkFWwHXw0sr6T5geKn
4V8apzVPxoqg41GiqJxP7kylPRu4tzykwzYJNTjUol1plmv5Y+RZnhPaiXMR+aeo
RgCmAmc8OxDE1okyROPmS7cNHvSSDbMWQgxo07GIN+4lhPvd4Zf9bl523OoewzCo
UQaHXYX2rjrwMuMqeWA7ftKGewMOH16z8RxFP5gF1rlK/PusD1U9qgg/1QZSedpY
YAl+y81wMEcd4Ej/hvQzTE6Wja2ffipzTc6i8XcHLCo=
`protect end_protected