`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23952 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
akBpHK9XojjdOyFTP3pOwrYbPr1+J3Tl50R2qpolXhAkoABVOsVG0ALgG6XCkPwv
rNLogCyXdrvXroVwBa2pSiT+AyYPPme+NS7jF5FewD+iyq3exzm72NEtHJCCydmW
jPXGtZPVmBzq3r3X9hdUsme65v/xW4mUD9+EEdwVmGxbksI6p31GWo8px3DGWUVF
Drs9vsOf0P3qAOlFZzQOZrZKWMhum63MAh+Gm4rs49KpM+xj0qjecTpcF6zrXWVM
p86da7PwOhQ1aAALNqQ+ZGU9FRxVSJcPBd46NTiVG8a8f6qWTw9m/VLMavaRf3jv
5q0X93nxVFvRmt2sPk0oQ/1sUJmc5VrjXG4wka/eIY/mztj5lptCib++4W3KkaN0
v/pLqY2x2Yn9irlMzlxjjEBnPWdm/VjQITWfY1MDfQevfpaBr58RpHVBqaCXlkfI
PCQUhQ7mDG6r1IQAamNj4HpwZGGuHB4xfHFMZoLcJGBps261NhTIWizxStQ6gsg4
E2uWp8p6GCmsm22sL66+2ix1mHJ3IaLQxbkIj0IOUn1D4hIMs8eQYHrt2edPj8rh
qMqiMe/SdtsagOKssq0XDcsrSDfNhDQzae8D1Nq0+By7lDv5G/BEMspuJzQR7R6W
L6vPbb1i0onpq5/w+/M5cvCgQMAkoQ3c+Z63zORUtACciSKzkrSJjK+M2/0Fk2CQ
KXOBtpx5SYstRHYrqYZZ0jDX5GBp54VUHpjnS3XIkzKNgxJb8+MTnb3WEXaDjJII
CitypNb7r+q5bPt7+8HykN6wBZOfpxdaRU24snYi2039DsjzHs17oiEOXV2J1EOQ
xSkOk5o2fSdZy4oXPmPKxqojbCCYKvdWX1RU6DtzEPtWxQlc2ChuT6tPs3qt72x3
m9PuN/aukOLfAsyIJmhLgLWiahUwnUEySUiiIfrELBaucdWeiUtZutnQp0UcCLsX
YegPbektkY4K/NpOo8DaOfk50JCQY5BUN9+TlvJ+/D9Z9rR29F9rbKlZNs932CHl
+pq5hGgspTVRuuqakMPxFPaFhdrhAu3qvWYUlvG75XIaEJ4hCd99pDSOPACEvyAJ
7xz6vtZN4Ik+kBKBdxaCyVIFrPdq0YcCRMqET+yIZpPjnoYHc4PUBPgJ36aAGbX4
0/x1D51rPAFqB1QM9JjK9HkRia7/6CHiPxdcpwJ0NOfEILqMbLf7ZLxPpibbRex9
cJYDruclujL/ru2TtLoVWUanxeiT7Sv+KpGTTnHN7Ci52JikcoLz/7/k1/Gf2+i9
6QRd64pu0J0nGyJmtm5QpgxEhoY+zpUnjDgIJly+DiUjkeq3iETtfXV/62HHi3UC
coD4OWlIZstGqPhrdzcXZHpZjuQXcQwX/rADLZdDlUg+HFGj912uCm6KDjfUeNp0
EJbco57iBhQRXnmTr+3I4q9AYUOTVSKFtAyn1XSg12e+KjxEqmQraxiutX0MLvEY
CbTLThkuOIhTXQoQudOLs9uCSt9EbCz4vO2JJfRgHBhkbLGLbVc+KT/KkC2hCbAc
jENLwOppbw/yFTVg+IaxTg3cjQtvFYFnd/pe4g5YQ+h576MVuqvJOMbj0xlGD8AD
bngs/xbe8i8WRkaT8dAdD+l0V4YKHAMMtxv1TeQfbaBEPliIba2i1u5FRGxKQ3C7
EqOYmlT4In7UIldJ/s4XL/H9SD7D61GYsie7NFpkyanJSGg5y4s5vDuCv7qidXpu
5fo5RyJhl1R+nW2/foJkrr76fCrDiLnqNbNzKSTxdjJfXEmBGshnpydVQehTspwF
oAzee2c3Z5tsd664YeUQ0undj8SN5iuhMK6EaZ8m/q7ybdYuDSx2/7pWcWj3MDa7
lJtY57uef3JoL4x7jTsgefPMI718SFT5Asj6W0RSfL86aFYvB7gr5ZaCC7oOs05r
bxMSDvfdhT7bVuVAcQzW/3hVLlIpbMuhaEhR0n5+O8/jYERCF1ak5m3DEX2igOdg
MBnAzYu6eKvRtnHKM+WoL9Hs7uK7EGT39ltIMaBGJ92YUEZei6O+zN559pNOjNr+
oXXdgoOYcq2gj6NYzpLQQmiPa2MCEV6GhIEfJqVrgqPybV0lyujrKuJl7F0hM1fe
RxIfC/uDNW+SdTS+XXZz7q2j7EHILNg8KIY67BTH9WXYkAE2LOOUAkCzHMLIh+aK
D8I90LF/xCkTEQN1HnrV8kQmmJNxCcVM/rZhiWcx3VyDMKyTH29bHy2fQygJP09n
3EDr8RH9j7Rbh8Vg6fLfW1fLqOa9Tp5rfxiAHAQNmYKQfsYMYh4BiRlxLIcTbknl
AnRCJ+jWc7KK+YRmC8u0cqZe1sxwkSaCWI6vt4B31IHHc1Lqjy4syVCDGjrhSyDc
0+0riBVza7iDPScONlMP1lhpOs7gMlPa55Z4AGj3+rZ0he4AcTlLXaIP1NMoe43G
XmPHOyN9sJbeeTfkrixKnX6VFfOpyE61+WP5f+CooTP6Vh2fZhNZ14s5BRp28OZk
pD9D4pHM4iGtgpVkBAi9CA5Eawt0TIRWJYp11M/IqlXrJLnJBxjJ2gmOvOGfUpkM
B86lre0qKNHdQtSK/NfVq+1NfZYb5RzJLF3obBlRCUvDbVb293/4OIKBxnul4mhy
5ATxfWilpRTN2KJzWbGSrIW2BKVVkAHIn+tdtuRsl6eJcLBeQ0VreixPgreSwtFw
I8EVv2nK2jxr3vQUXvVLF7yA5oOsRjDnbzq8hZChglwKBiJkm6BHT1tSrj/rzZso
H9jRc7UmQzRXYuNZvIdH2m8Z80m7lAp6vziOvfH+WV+ZYMXKLi2HBavv4577SNZf
JTlHiSdyVnJLLJMqGJZe1iDUDPwXASgYCHY2iH3iGqs8SNkqjcOoeDhHnIBYQ5a8
rD02PfIqfYGZz6dknN3c9ZADIGeRkD4VoUXCmTs1rssFOZOADSRORUA8mKPtHjby
eHAM79TYSTSUik5K7TJgoV7xpB5lUE0JnwyUjdvX2OdW/VPQ8AnkwfQ6mpVO+ZbQ
LrgDLUa78lg2bQX+yUAxiGo3Fq9usi3SwGVAKUTL/LKXoanQvl81MQwMaOIS2Z3v
Xzhpklu9vECt/Dqpufk7GhceR4qeVp1v+qlkkC9cK6US8YCslFH34jzfthhA4bD3
ALdr9DfBXc7Tg+Df7MvEBVBvrSXhmDDyWiYKM8O8AVQyPDK1agbbnfx8tq2JymPU
4UTX0ld57NttvXWUE73U2ySrEhk5hEQUIA9w03HxZFIdjsZGNog72xBdaHG6aNpL
Kh1osWoNhm6UGjzyWA2P5LIv0y56EIu1Jnb9ZiczaFJ5NFduEcTDz6yzTCgKfe2x
020iN7+jUvrDjUi0kANVrr49+bm+vGaPxoYGdRKZqu6A8b+IJOb3gJ9qTnTXb2ah
Ctu/ZlbqIpgaWA4U/RhT5tYj155mhHbmu9Tp+Dvar8JpcKKEveDUilLDCtQfZtPK
dYIBGYryhTHrGf5zmsJhyjettigroy0ByZJ7FH3JoOkfLXZiFBrKk+gVNojs1gOh
jPJU9YlCv6BRyj2vqZ72uEVrMYEfjoyfuHZ5+58R3iQAGCgRIb9YomUtmEqplHC4
LGWa2ek8LJasd0LlkFTpjdTytWs3VsNZYFfIIts0y0jRZihM36nlNgkk+DJ4QAyL
lINo0NuozhQyt+h2TMhZytwNf0bonAfyqRl9mi5iU+VZwXIeCMpHeBubOFHsftb0
DZ6NCxvnJUNSxmXaqtBvf1vi3FTk9LAyq6GhZbFza3/J98VzNQoVIFfK56A4iFcl
flxcD9n3AVVd6AyqSLQRLglQsyTtcqj2eN/E4fOQjevU8RcFIdiRhZ8ZskgfDlEx
bmuNsJEuxokg7doBxZEmI+HP7Jq3mIlZYamlpvNIYJDGyyVIMUmuxaXA+gkii0ib
P4+G+g17tdFn6va8SH1vI7opfQ4aLJ13haFlrNsG1QMa6zLwbvNFUVXkwpZh/Lcg
8ZHTbI0ixMmjN2n1TT3dgKzLuG8LdfZ0IolCyKH4Z1QWh+tem2J6l1zp71zBZsTa
6QdvJqfHz8LtdsipQxPbJmnNyMBgCOSfsElgyjx05dXXVd7gaqjCtmOUA9ckUcv6
rMnHDe1FxCu9LHNWhrSlM7KY4CVm5H035p2Yv6+/rGSMVF1/Nlymt9e9TVvbvL5Q
MNaWsn4P7Ty5e97aynXbSFpRsfRcEhYtLZj2DOcmHgAZVaT1C9mi4OPSQ6XFT/3K
9G86C60ut0+eX0FlWkLxOV+nmzDISibSzSSHnLIodHNeGyhqQVSfmD5Vunm1G36q
bArE6gflFE8wa69TYVFpSYJS/RD1qmxIcGG24jVtyP00CF3+h8heSNqMGIWVrLDk
Q+GZz/sTpR2BIu36+WxcHzRerdwy2E1b643e2DaV3eXWNqSExigt7pDjBG0uGzhs
ypuq1Sv622TekiyuIpX1EAdHTdsraeJNEd9Uj+U9DjcuU+k4BFV/Sos5rijl5MvE
vu0tboFNbG6D9JwrSYiLNRvXhz/WSxCZk1+BSOl3HJogqo5/aS7dUDatb9IXjjjb
gmPhBfCCfHOwRKnwQyFGGGediZgH2OCKJKxCqurRTaf09je8fRxMoZ0bNy+NAbix
Yu1WyPYatcPb0SIlaPovLAaVYdF5+8L05ZrYlPAvl96fLwvTaOkZGUmU8RSg4CVx
aG+ZN/rnYwpBAM89iJob5iaIYPyUH5WRI7uCTg5C2xmzoz150r+nOuX7svlV+PXT
Phw+wjPMok5MjuPVM7NFyWEXpzjo2vDlq9iizA74/30rFZSCN/w13iafh54yQUC9
YG44Q/DODDdSemVhuLov4E65FLFJ2lVXbfa0RPbWIpZGUEGpDgauyeoWusnt64k4
Djlz+Whv+jRitK23lFQbpeiK3x7h3w5sjyM4uBLHRsaXyNa1ivbn1e/sk/s66U4b
IayYgjYrI53mWn3C02schKG09r1bfxVLfAvti/8Z0tx+mkj2bsm60eztbgPUIczk
9JV2kYGryvf7Bd96mxjR5cHAPLhxa52Em9RylJiAkRx5cuhQzma7+HNa53bGbGnd
6X3FxrFvqCUQ0ogrsZYb/FHiLkFF7i2LEMF+7qbapzAAald7glLxuF3+Uq+WzmuU
y9kEie4u2MRZXjL3vrgKoLYLtdl3L4YKIGj3qQc8e3QF6CKdiJDp+a8zrRpMEzpV
2XZVOdINPgqGTzOP6jzoyvlYV+rHS5bz46oJoMa2NpIWfWjesbnBy2jeqveI/BLx
7Ckusn7D0WzQ4rDylCOBEuoU9sfaUEtd4xIhV4xF22e+KJWrL+k+2TMmD9aPbCcJ
JoKgkcpSj0BdhN5eFvS+odQXLMRuhVZ1pgoMLYcwijyIEZssUbND++ZiLTh97xVo
wj45dorKdtmNcI+P6hiQEqOnQjAr2AYoyccfIReRjR8H5FYrKYzLRfmd9VKpjk1n
65A2AQFNePtPS9H0AU6gG48APrdglwIxcV96V/jGjxYK49u+BkGZeFJihkBUeDfN
QHtiNPi7MSDWy4/+UsFQAcHckIqimyKKp/cNFcbWwiYeVP+nA936ZRLNeePtVSLO
jlL3VCvV5WZEhp8Gd192mVGHDgQGZwxhIHoGBZiqNEbpz4CU00nCevQdtNbZ16+2
wdQ4fMGTgxbjyiHxtq50Z2m07TS8t1iEfwNQv6ScSgYO8lt8x94BaKPK4knyCeXy
oWqwPytB6hbSFVKLIcU00WByzldb5L7VpMVBKSJAdshWRz2CQrEnHljRSAyXVL57
wT+Tpr5l5IjO/bWwvisCzs/waJu2QsdfDS9CqbzxCBJJqs2eY1NMSknoKQArtJ76
JD0Gvb4RWci3cETSA2vuVI9+rf4TtrpIzPQOCQKeq/emM+L+Q1jCFfoHLqKkSl2i
0zzOSE4V2RQxL5aUXz3jDBcy6qHVYnwaUD3/oNHb48Tb9yMQSBqnjoaT+3p5IQuX
rxUTRXEmDKVbEoguEIE/z/RmUtrBLeSU+JasupSauF348tiE4/RBI0jcPOh14fXl
xx0nR/isesj9qonvmUpXQ8KATY9qYKLd8c8fo4lVrSZIoq4pbor9oyr3bfGQ/Iqk
3o9NXAEU5jX4CgrU5vxSWNkdgoS6fql3VuoIAApURj2LKEQ6kIcGw9EfwarSJhWc
Tpjl6ylpdB6STjYE70tEa4C2vyNyvBL4LCwyUEyiPs+3IAsTaU+9As/JcCNgcEJI
lJ62BvgFrhpqpEA/opfE7jF+xXIcBl/Hn6Hev/01psYp7FJyfsSkRBpy1QbtNQ09
EANaWTaKu61sGqZTUhqX/xZDVJgReQ79Wti0XzXKkMW3SgK9FrHKApcXmFPQ0tLQ
xNI0DAii9Y8RcVm8Pr4MjgotdYjooVqDBs+h6H0OS+cXljDG3J6Rq4gXQqGtr+Fz
JU++Bq3aJ9UiDh1Tk+4Eux7YjVsDRujKynaC9L61qaJ6hyGBREY3ykjXv6NcQThH
cICne3VXjuj2r8mHq3r5Q2/kyGtEQdUrMPajT2KtRq2Rser/ElXwLiFaK8T9H+6g
Sm7pkMUNkqfnflq4sYeclbPg7Q9LAL2YG9pI67lkp7QlEMtD5HlXJoOsTsBE94bh
iWORyZqJ9mLfqssIDEhrKSfp7manrkKF+uzF8rux0SfC46qbll1bkIf9TT87kSZP
E/o3dEhIUTntbwz7uvWLzMebb12AJK/c6gP/ueXmEdcBleyWTPAYiQUW9UT3eThZ
rn6entsWOqFr30iZz4WcXDayw2zMGuNtZt7nbW8kVDZztn5wWOdLwrj7R80FVptP
cX/cES5dQfsBh+8h14BO5ETgDoF6Lq1ufTZBsfWtlgJ4H+F6X1A9wMZXh6d+BqvS
w/auDWKOjWdAJd/TUI/wg4fQIx7TXSyYfMbPu0aCAj82LlvjHFFbUox2BUkAXOx2
WkimSnpeaf0CjngkU8H1QDz5iFm+7fySr37E8MbBaTyVtNGRcdV4h3Fy66tUD+T9
e0LD7bUEDQ7XCqB8LgS8B6lROAtyydadaQsqzVGq0vkalPqVruOFe+PmcBtrUtrq
ENaxFp3GR76jejYNZttnipgOkv1Mcb04RKKqSn0fkvHCpGBV+NHDJYJ3tj4TScPJ
dojHrWbvNLTEA3YwbFZRf/q/5eCnYhX2nl9ajZORHPwuNmcBk39IgSfyDSC/lSGB
NpTEPZqAIOVbMb8QSIurTTfn0xKavLSh/xZwCSdKfV2BlklJrbPfGBMBOkgnlcZs
ERCyvk2gHr4AXNUqO/scMmpG7H5I9yATFPDxfJ1lpu8ppZKFyFm0v7LK3Kogvi87
rHiIKjLrtcDP0LpxPw0zsYMf8dWYqCY+GGd1XfIB9/UURV0PNsu4/Nkov5SGRRDI
xucL2ftwLjGq5wsrGu6bD34KtyuJ8a5OmsAKFtk5q1Aq7dj1R+uMWxXsq3N9MkuR
fhGrJxIEaRcI5SIVXvYaUwixNMLMh9IpPS/flT/Egr76gOTlfY1K4+vD5DBlYcq7
6vFpt9p/wb/HAoQnPMNTuMKUClaz0/+ZlxBxhpatvlom9CECnpi4EUa8MMljnu+A
uaKufOnSpnEwD+Ll7Trae0yPwkSaIb1cNRrJINgBOhzjqcPug+3IzoFGr1RVb24G
EsaQd4ZDz4lfQMGuRjs5dyMtD2bLJvhm0an5Ef/TJunnVqySLillaUW3TnlLT7VM
eVUjXFKa8U2oTTmUj9puR78maiA7Rh4CCesaFdRfuau6uLynDu1AvOQWeuGO/biA
cJRdxYw37xwULH3SNQWA7872+7hidVf/+XM9W5Jl6qwWx13IoWpbaguO8l7YCopp
kb3AkRuxHywJ2epvpAfQWBMTbenPLythWGCddinIOfXwwqw3F7Iks6VdQgybKter
gorRk+gj6Uvp4lH6pZ1nzz1NHt5t7F/db6Flsf5j+BtgcXI3lOK+NgMVKFNxONa5
esAv9KcJC+5IFT48J5J+ppmcv+is+FKGzy3Pp6fIS6tZIm0kE0D4TbvWhEg+0Uj+
IhOb1Fv6bKXICXP9LDQmywax0BMWiNpAwYfGWxJHv7PR4WgcF/Vo2qZZ43VY+XC+
/ek4dqoH9avv6t7MLMSUIeRkJMe9MPecpboN4c64YgoZuewfBpiL/aCztsGcKKuL
tki1fdxTpZNk8tZueP6+/hsufl5DdEC47tO+xm6IO6Y+jCK2hmxZApzsCxCfYoZT
q+DUmaM751if2klAXfo7dH9WIq6P3i3y+nv2QgYHsf5QFXMX0zClpA/g+TlTvrmc
gIINQ/93eRcdmYtW7APSIXNmC2b5nr76p6nMLMvR5vipCs37xj/Dow2UN9qAtD72
WfiLp6YOVya4ANCCZ/kPuQQ/0lWIRyozQFiHXXEMQ89rJ4Y7OCZmFxmfBj3zICF7
t3ci/a/8urTu0T5Mxofz7Ld9LNSJD82f3NbCkTKuz+8+7pzNd+pDYMd7piIZ3jR+
EJ2zO2bLdxM23UNF9fuIGbLFlanBVeUaCyR03kiOUjREU0O6c+k0MzkR+56cCdUg
cIZC1B97RNgpgMEBaRtp6teEMjZIaDih6zarmr00RxGvsOd0LAwNuEP3+6e9IPpg
n2MD0H83OZE044G1gjgfiKOgdGiaDwdxoSnNqJ5lhzmCXTHSKXp+kFxozd1xe+bx
15L66kRf9XJTbKaJyMqS00A4KPKd4xSpRYKKdBWq16WbPoMht0K6t2qFfxkX2Rf7
ivW3eP7dqfq7LmOmhiABnmby/vwTznHIZsRH5kmEpkO1+QUaL/dzyCkU9FlShhMS
gpa2XUw4u82HhyofRYob3LZkZ3tJaxCsimTP5VcoiDkLmjxjjE0+OEO0QSza1Kyl
+8rTIs8BhiRoYCZAojZqOnYTzTWGNBuBcvRZFK5d5o32NYlbXqZi9ucJzhRSSsW4
5G5B/Ampx2RRq0Lg4XYl4SLaxdpyNVtq+yvKCY59/jjNADiQyTsoAcBiLiHrvSXQ
E4XzimFNclNuw6ZtBodQ+IqVFgvonJG/zVMyMwEwi764xSasiNpFExRn3q0xbxx4
1ah/ZjvV3nDTC0l8JEquAtBdV7zIk2hmIx2qnLJvSfQtzVWkU490cYcH7DZOF0L0
5p796wYfkOHwyfIhQEsO66kqNP/VF6bOdttT/qdMdKwflJwj2UnVv/b2d2ScB1KQ
AqGUBMTeLCQPXYmYQMGxfHY5U8sERgC3bHRcuJF228QQXEIdos2cFzQvmzv3f+ro
Qza8MRN9hqtQsoPo/f+7qsr8CEZT7nWuo9QlJjTAvE1ILrGrIRRuFKwQ+Tu2xvGb
q8gE1suUvHlxNBleYeEEo7Xm8THBxJm/mvFyd7gmTkqcP+351sBamh8nlRwfA8y6
EPzE0m5BJ/Wk9lHCFkbIct/qiCot5DWCkFnmOUMiy9dpL5SDOcAOUE+LLapuPnqQ
kMPJpUZDzPVvrzOICxs6ltCz4SsS6ajEAmho4JAcdzhughV6cIMKBIlahp4Ih3YU
kVd8HuxRccdRkpjdM0SPXajmybN6B+5aYfg+FedNiYvRjB+AYKzqBCscc7rvCwlA
jvZutxXDU7O0pnXhACwYnPnngYSIQod7UwhhKhTuwfoDXKP4G4mE+BEJdI4v5U+3
ImfWJgpy9SnCLWVu6aGj93O8ciSYxOwO5e8QCgCKuFlnxD9VFvqffJ5Tt0WRHqs/
YuPQJ/NMUOlKrGmygMvyLcECSeZS39SPEMb8gFXbFq8ib5bqxpU2jX6tBU4HT1+d
gB3Y/qPe7LDSezWPynY+l531sO9GvzdHaBoKvzjb47viWqN1U8zTs5Z91ZPtx3QY
Ko0zJNUOjesnMKqD3YF5gJjPORgAUmDSSvLElFj0GvzLjP4xMxP27yQxwuWTyzeQ
rk5/wD6WByuzV760wkFlJx5rzT+mVnfnSN/AXSCyOMr6pybC+9aavo4inxRSM63F
CC6BDMjNBE9Qwpd1iTk2S7Mu6m1np4pP6WrjKY9TJ6asGsYIAF6G58PhOu7KD47X
W59munHWhdfYTGhaBCEQrTd1/nZpqjDTy/gvs1p1hRSyCaFrpNZyEbUDcnmybtds
/LqgRngqb8QahLTQEHgS0r8ahyXJzMYTCOEBdCFF2zo7069EC3Kx+ocSyR05mbng
mAR5Pil7PyJWv5iKSSUTb7n3JI1EazdHZPtd3vWPQ6mDXvBwd6BkGGuCcU6jupwX
zXMxrN56I1uc6xserqhZLKRXVtWBHQ3rwuY9jK6j+QnkhmgCkK72PhX+UVwnc+Uu
1VUqW7GUgiZj6KHmjHmlr04o0Q9e+K6E1T8/QPqwreIrYa0zy+saiP0J4MkjhYd6
jabf2uFMd9tmcT+LDwwyDeRHuLcukxe4wKe0rNQ78BuNZeFGhvDw5FABBAuik1VW
chTSeOT9QyWlzmE1WviQfrts1OPmuxJt+xF/KhVXyowP2Ml7DiM1+Jkj2D+IFw9r
ek7GQpqT5bSXjmprOi5D0lDy/wxGexsQspX3Pl2R4rLRzXdyTAOuWtzp6xTgqoaN
fJoRn3F+o3frteoecj4N1HCtYyDQ00IL0gk/4W4Etk+NPn/R0Pe7j6tlj02/aDIH
McNU5wF62w+Kf26vvaAZTn+CyReQOv8K5dJbePl5SFvc47vYEfdhDVlZ1TlJQJ4c
QOv5yOJ1qmQe8b2GYNE/9gWp4I3vIorNrnmHxFKSZrV4w+j6k2uGG7dhnVS+NTxI
lmBjRgm49Sg86oSmvdNFZ4nfWztD01dzrJ4YAkXT6WOVIS1j21ioSDzzPPkladMF
VJV76bhvUfqwYKIXqfGNbfh3LM3L3Xh8SlUBCy6Su5QO6j7h5StkuZqiuvBx2KDN
2C8dCLm5MVOHugtX3LtUBqtNKqhXhpxii+CSGxhnnGqAMnY7xdeHZcMwIKDdl4Zm
HcV2KMJ1pbZoRdOSBi1pqD0l19z73jU9Ym3ocs53bw2BcT52WBfgB86/8Mx54ktr
1PIwK2iSlgZD9zCRaCGn4h1QdhotthcnhkfjMx+/PT09KY5Jd0lt4TOYkUTEw/jV
PdjOAt/XKbQOhSeSiSB47Jco1JeUASBzlP/jb7mmKC0qX8sjj+e/wFb3pMc+gP3w
Y7Z4e6YHgTC+ypoeq19gH7CV3Vu29eY4Ppm1CXF06x9p3yZafTwj213Qmn4K/O9t
NZEeSJmyU+ykfH6Hv7PNCEMeH3Hvw8NBY3m0hjVuTvmgov6b0UHbutymYEIkKJeM
yIf7DsJMvT1i+RBI44Si+FM8ySZtWBwFJSOmWhR+wJ4TmZFU4HwLt8n0v2Z+HWnT
eyxj7lyU7YwIoU8L82ClxCDPCQrYev5D+lx2fq0o/o4xJGiDfydAzrXQkGpF8yN5
ixVNIDYx0vjN5591aVANoll3PFlNyqeGe4oeTfk7zhPyU0cs+4jcrMsc3NTnhs0P
CTJxLUx9yJtcgVjyqYWKyJYtV9fXXpcmRKPR2YJepOVigPl+pkNiE1AoqMZ0gdgU
1GnZYxuTGN1TfSNSH/dfUx3p6gBVvYgEqLqYXi8l50s9HFrG/9EC7B+G93mKVVTX
v1KhTLWJdYr0dUi/4uB+4/IGCK7ltA3f8rxLQ4t1uG43AMsDZXt0XyGpjrijVS+Z
7JpzIVBJWPW7+MAIUfC+lJly+MuIa9QXfq4+ew6orWF+6zeoZ85uIKgC+U7HZZQf
JopSfq3ESBoiwmDFgUdF6Jke+ot7SOEXDW9iuMjDS0c2hpq8V1OiAj4mZV7h3NQf
zLa4tyeoVeshU9vNn4nLUY4xK4S4bpou8kU0m9v74qjEJJQkn6cNhUmQ9tr9s7p9
8yeO4bCUZNZQ9v0McyEq4C9SIZv8qFhdB39/7FigKUsRcVahSWx3QIy/s52L5UEU
64cY7p0bUVczjkXGLtJHdBrPrq3DGGx061ITeffUMucj0kOwNNaboHrgF93I6cKi
vn0/kVSkC6Z4ZQG6obbG7lCJiqOef83ulhQpo0rxCFF+UsRD38mkN2t5PXRiKxfa
lGBWuAAIyh/Pe7Lh/lmGBzAJaQg9wtpFONr2slUdX1Q6sPXq0C4zDk012WBJRVAK
VhCiruFfu8v6RJBTqmVQeTusAxzKmQnVXtuhQnJbwawYH0frx69UMxyx18L3o0C9
7Yl1ghwAQ8hngSdMqJsFMSV9lc+q3CMOP1sTzLapf8rJxmFaFGLbDxwC83ezBWd6
B81DF/yx8h7bbSkO8H5WVJ6BniYYFxNeABpLGDeC0GEArP7YU6CLxBjGHZuU242e
+8pTOiRDHcsSYUjY/AAu7rLrxhtFHXaebk8VJy+U6yKQSI42xvo3b8+LttSHVmXa
DfaGnMR3iGWRaRDy5/P+USgB9pskHzBhpKAWOxjEXbNZLz96m1vGAlBxhtSMVoJj
r+Cv99YwPrUMFIOfIy19hlibl77iy2A5Rv03gaZIUwEPA04k5rR/MeAn5l3Ohbvu
lGwedLwaCkC878X+kiTjIE6efTcQqMTcBP/YtSnCwQyZALZl6CxnS40tNwCljnaH
Zznn1W/d+eICev6IyND+au4UeEXgJKRfsB9DWK7L+n7Ir8+vfWtml4fWXtvDTE73
9H3v+oKTCXmkKSjJd34W+GIqe9KOAUFgB5ni78ap+rzu28YabvbWCPN4AMVvyNQ0
5sAv78mMFXpuIdbdBuo4N1jxV5zxkMHwJXGcXdN+tBTrVUgxs6y6JljT7nJGZJ4A
lsFJg6wEe3QNMFzH5ErhIuLP6hiPo1IcTCE1TdBx03n7c7wR1O1K0I4zFF0zXOyH
mhB8T0IPUmJkw64WOsU0gqIAONi5e+acojDl15rTQj8xr8VCtoWeuhvzhnV7kSNX
HyNeenq94Rcl3Oy+ov78xrMEHi6di6jUZZ6YyphYhWdKC+7gq8LmiTrxrxwxbvT8
qaPiV0gLysj6V/ula0+f7xUbrGpDdAq9viC/Z1oubtMy49jca1Bsr7dUiPB3iFgJ
PgVu6LManDX3cQtsSpve977s8LjvnlnAY6XphuGWmhRuA7XiiyWDvQdLKeBipKXt
8QeDtmB2q7Ul+LjQKe3xKSX8ndjCxsYgtUm/LOHcdJBxC+ZuIMfuAKIX+p6DeDEi
Z53xWL3vQoWnUHEhPuniHts0e0W+ilZinC62A2krpDMKyxq7jeikMjf9n0tgith/
W5rK5qK4PzLlb+lGRaOK3CAlw9S567ytBUOLgplE9l6qVJ3gFcrVs9rMOFkyGszs
Yx6hp8aZgDuafL4nFFPboc6VjIm8bFFwIYq0F4zG1cUPsN//9xvoEuSgl/3s8IIg
ga5qjFKk1i1Qv5T9p0DoYWhJRE39Z22CPKhfDAYMyYhAq+IHcIiKDIhpgKegYTrl
8Chw/tK//MxmOSnrSTmmi6W1YytvTxLKzl+VytZ2UrtwmqryK/fUSx4WU+yAIzuD
tmgHYZeWySs+4DF41nvSfYNCaB8hH4Z3m5v3diO9aHAWeHACEQTV0d06KGjCwj+z
+U7t+6KXn7ii7JdnPMGe/dtlleu4s8kKKvjWEcqV3GJ6Lfolo8b/enGg9GMPLbBD
SZMeeM+EwmbAUZZrUGc1IVoNauwQI/6/HscoBONXqnvdkTnRl+mdvrspFdeFuLqg
yT+g87+hc1xZDOd/cCbQiXv0uG3Q4PgawilK3jj73jsLA7bCFiTHwcluQKk2jUz6
dgQ/sbWxVqXiFn4ooNpfOG0EdM3ak5/a258b8CqQEbRaYi7vLva9FJDvwOXKfR2O
uoZgNYcup8uW086aOAAlsO49FXIThudeGkFR8g6bstCXSelgHrqHC8PuwOtdU2TX
IWAHFx3Yr5D+zthqfWoLlXKRq/HFKuZOBDSfhXULu0eFFI69B0m+bAeU3gyPFIcV
sOtAkwcWPmAPBjOLjNUjfiMKHg9Fo+/c4+UU6K1op2PXLnZLoXvnbRidHaRP8XQ9
QPKD7G1LF/jX5B96XU7blphXXFAjHrYmD8BS9iMeezIMaEEYhoNGqwMCPk+zIaws
dpPyD6p+zmbtco0RC57LL+62J9C5+R+IXzio9mfHROjVnDqpJdNFzmaR5xjJ80To
g/OulwQICI0r1+DAObGECqt+MBFSif0g0baeRkm8F+nIA3w86ySJgk2KDcGvmCn3
kgmimsQJR4NEJ+F7roFm4sBVbX68Pv8UkoakOZuc22/OUNkzyWnxsVQcYWXSI79d
U+qMihmEar3L440FCrrKU2xLzArJyjQ0w8izc7GPYRzdMDlZQRGzqFLNs+R5N723
tzIV/UAArtusOodvX4709Xi0Ww6KuNMArO0nbNIPu/Cv88bb0gbi2qGZpu4GqhGd
fnhBdPFF42ZSBm4/C1ic4M5sCpqF2UHAzNiUp02xROpPxQW24d3vQHXnd/zXmK2P
7Nv7arHgWcbPHRNlhx/2443GNODxDahM8oVcRT69t7B9ce6Z5vxLwKKSnpZqj45p
HhXZgw63IAdROahwQ8XfZmZh8Nv+bQWLQlEgnmYB4by1I8kEGKnP3Pptee+tyU8w
/73fgLXpNW5YytMPcigwdPAM69xo9pKL+2qHgb6khEbpGFJDIwttrJ3gef4XZSo0
FKIj7s1ePlWwrqHKvRYXTZw91n0BD4fC91j17nAb3/pHTT/TTB6yni5CLpPSZ/Ga
TgDYf1oigFUiVTe8BpFnVik62/eQEeUodIKiqEDnpB2ow2wH3FZxtGCO5bnguVTK
QN0qlYr+wpzCL6PnGuUV0wim0pUv2zowopX3t2e2eG3k0vvYtwtzmB7QgWFPDi17
Dygqq3L1xV52qhLy+BPLVkSXpd0R5Rnk6hPo9UBl01HlZ3U0Fx+Q7/S85mKiMFQ5
AzbTVC1Hej3U5rYJBpqWm2pt0pc1pr8uQ27HtNNFhC2glns3m+5C/hGaAhyqqnRD
5pQo7iEE7k3/CpC+S6srdV8xDCIIzdoF9IKyx3StriHeKCux1hFNJ4YiUlnNVQEB
W7JT/SBrl4PuCgGKFolJeg9KDhJS4grKYzgZmg1NdTlrLUnoX2V/CN8XGWy4V7a1
sMcjWQfkhGUy4K0mwXLWdXm9aGoSIwH/87Sk40+275oXI6Ut4ZOT18/6pffPa1kB
7YgRBThCc+Ciu6rUoj9+KLi/ECTsIYD57W2+H6bUlaTuM4yEuQNCv2G/qGlnWXjb
SYMcfuG8Dc6hD4XR3MDvQ12luCQtsQB1YSR65m2wvJanr8xTRfNC/roi7y82BA79
XhF7lYgotmT7ZU8rhQIq8GQkYyMMb/uThmvhRLFqhwLojFChUw7+l0TOIu76uJMx
3kxDioBEamvJHNkdd1n64Y3hlg0IBKg9l/itUueb2AtRP7uHlkFVB7UuQBgGneXF
u7phaOQLnGh0l5roiuRlgjFuOXYsFIdMC9H7cMySAlgmFzyfOLrjh3NrjJhasF1r
A3nSAVtX+mYDOQV5/fJx3kxnWdQ3NhxpTwEbd6OE7xjr8JYdhz+p2VP6cy8kKOnI
WO12ZcQFjR3XS3ShkcfwdM/mOX/3gvxufhBWo0c053CExvbTAyKJ5O08tGzeJUBI
w8+rywENUbgAwN1E/0ww+4NQJnj+vwdGwSi0NaaqfboP8x0TypSmX02Y0Vs3V20g
uaiERK5GSik2P7jAkh7PsAju1firipbFHJ631XSsgXwz5XUpxoo5ultJLYunxIKC
SI1R2hXSNG6bxBWJoUydA3VDRFrn6BQ6PgPUcDnaSqnhUt9k1H92A9aEOIh4PH+2
oVaq3GHR8kzcVOOg56Ywjp9eLz74M41YdaodDoJBTzZEsbuSqLhoJcixcZ+/YIUZ
GIcR+unL/s1kCjiKZrxObi6zGwACFsZ15uTRiRepw62/RhcfkiXMM0UQRWbiUnU9
yC3bp47iywCRfeckbKF+LKHfyNU/n5uxSEiDgjvKRVxTHVUSn8L3QL5KJ/FqfrEQ
yGS7F9iwT4Ceq8/cZybbD7jPsSN0E6HWHzycoGHINveScDFRVS9h13yG1fgKX65Y
TDAE8rz1Oe0ghPoHbSxb+sviWAMEaGcAxaCrrZ/1oGdnJsKhcZRAs4td1FGQjpQF
LQPDeaoNHIhWFjr8mOfC8R5kD28UfSjNAJxJXitxzvqMAKylpMnFxoiLd+Lf449U
HNERTuQGhu8j9O+6NQzzgIV6kiUVviUjSVlcBJXMCKymxjEWZPGvUQ0SNPEMK1iv
tjHzSVCv1zqlcCKu8cSmJqizjbOV/XSq9zg7RZw0JELgnxy8E4GbOT7IJlLwn1YT
jeoP1Rvd/q6DsbnIYsKt49btG6h3RDCHry9c6e4vxqo+f1gAdxWUnkpHVbdgvyDG
VQEMB3xmJbZQXQy2grz6qs8xpwrrviqvEJgvDliY8PisaqRCNxb4qa2DrXtEa0UG
y7ex3Zze1CKg50idPSgorI90e/7eoEuIOfNAktw59D/wwPOd1c6gkuxry0LoQ2VA
WMzRiRgoj1NFHZJ6p+bNRu/3DjDD4ggaLihstEpvGUn8GlbLi482keyFFD40f/56
poY7ILXcumpqlZc+lApnnbWhd8aFMOA6voalFfw+GFhlPFM5O8h/5fPVvBr8ARLl
080sgWxMyUYML8nMoMZ7lyJHngRDtaSC0jzUW6hYfmE1piD9Uy7WuWZwWmc8N5bU
s21fwPFBI7EAx2elFfrjfbqPEIVZ0JHltlo6z/m84pdRkq6goVRlAJCm1egr9wDz
NAIiC6pTOzNVQYZHCtD0AT5hhiXDw2lFDhZaX3smtjDcKIgiM5jNlvvmKeEul0oh
8a3jBuD+YTRYJPDtkaCuslo/OqffrJLgChI4yOVNVDQrE2FyVHgn1HgVLw23QaxP
6ZKINYylILlpai3adkkL2oV845to6jxTg58fK/7/38e1g1aLtJRH45+8HkKzSdOQ
oW0+9TYDdMaqjrOE8BIfMXEx6///cL0dsnJVmdPV9BzqPuY8ZxPJpqNdrI4R2YLp
UFu6ph0aU4/TuA88KH0yWYGBF2VuFswHyWis7OFkxOCKwRQNyGoFVLODF83jI77b
jdBZJG1vP76mev7uZbnxe3GZIWW6YzaLOUIMWZ4HGE9jru7PA2gY39J7BZcjmfd3
jfwtCWXxLdSphb4UOj9piMsPaPoLlZ6fPb47RAdMjROmLoWpmab8/8M6l3sNFYyu
ofOpgjZVMihYE/IAMSDvdp3bqz6Q4C/n+cUvqk+1YtzxMfDCfNvfRf0t0Hs1ag7W
6sIPYow5X4tRmnYOZyKzjvMiEfo8GBqU5e8dGgRECEys9rznHTgHJ3uPgt6cHXwe
ig/ZqD3nEOvwrt9BBVZnei4WZY4RUdXi1TGdgk2danEeTerWIUYNbfWhFxNAR8c6
NTPoJnjduM9R2vM6B2e3Xyx7C/p8JHxapi4YWPUKaov7XCbZ+7xBftpT56SLBAjp
VFrTzCX5y2zFACqN2kgPSgRPeW0g89b95SG3UStQHLmnrbvy2HMxqXRpJS9kaVp/
TKObwMH8DQHTn8lBPwykyXx0aKolEKAbyEzc/Pzp9Ml9VJ7RFOPa3fUWpK496cPl
P9UvlV82mJwyMSWJli7wfQl/3jIL3N8LKK7haY/8w7aXINV2fAUu+StVgmNARjFf
zdEz7DmKh3g7oyrAjKvi7xAu/44ui9DPhQ7keORpyEBW7k2bcpuCGrguz20glUmx
JwR1SXP81auUgbE9lkQgaiEn2WGNiupF+Dy5YG4OmPlsjKB0DBoIkn5N+LmsvV8n
0CUadfBYWekyjjeCJ2A+x2PGNPrNluCy0FKVFePFHiDpLwce76Mx4atE7BGWYuBY
SzxMgDOOVuDZC0lXRpZf4AHmvWgpOZjNupnLlovRNqx6McG7UEsQVBVtaYadgtEM
9g5nMjCllXasGjSVVctMK2MG0ZLl1HB8Eo4Wqwa6nQqx6sCd9ZaGmaO9yfVyft2a
r9oQYggXsufWR4vP5h0a14dNyvZK4S6Qs7WB+iXJ2CcBp/yjSVl3aO1opm2NGFOV
cxFDD7cIFeNDVGo6pRq8wDrVpcPyOd4EWLG5qPL2Wh/Uh+LTBqGlBJ90O6mk+Oct
BHBjXEKWcbuo5GJlWXqgOuBoGx7P3UrW8tCJ4gUq2IiCnYS3BHkQ7Ms5puG+wr3c
o54T9W0O6Hk3rWTzj0RoMapbPOPr4Bl3yBwhYhSG3eE6q8kCh7k+vk9jRj3HHfjz
wV+fMmUBcOJQY8WK6UknekOYMfUV98xIiuuzBcl57VMrn9v3LU1WhwagUUjCPc96
81xDUHEd9CUnt7W8zhIlhocr9GLoqGQX4gh0tJMYXYlgez0LizDIRNUA1DM39s8Y
H4xvuhSE9JQwfauiBYejkYYGYQDLXwShsNUXymuqWnk21n+qHQTycE7bud435x5T
JsMMZCUzro8gsjSgG3u+qXcGgkv5Y8S85XkpZI6bh4xJuH9ftFXLT8tC7IT/D6ZW
e4CrhNPzAWbd7hvYN90s7CmtkCFdHKJ0Xz0nGAEZkBRGgjtTUuhsTMqn3cttWmrv
a2C56s1a385Y9iYmDayTzVtE8JoCUzJZLdjicZCkP+ij/xxEiSSctnfyy4Y/vA70
7lYMq4a2QE2mo0535NRw9LPQfIwJTmXTIwweFY7IPmDO5lbYxXQrYTIYciwDWuQx
jOSP060y1tjbF2FlHi+jCJnN35hHbbiqnEb7GQPp7LrUnchpfcNCik15qmXfwdDS
MUXsnhprCe1oWzrlxjN9dH0Mq26XEaDI4bcyO69RkmFsmHe2tDOgcjGbYY2N/thN
SfGJYp+xV54HKm2DzqczK5Od29uw3pB0BWL8XGxwgCOT9CmEc/aLk1WMtJmqulQi
BRo2yFAlMshwqM6wWzrb6bxnEjqF8hOs1/I4M1KZxs0SdwID39vxhxq49WvhptJY
yqSY4JdNhYDnDE1VRwBlJtQ8rtJJWUt4Fzd4jmsEZdcbzJdJqk5niO4NxwwZoZ+y
soEXbROOLljNGiLbJ5PlSZDfoJPS0yR/KmsvHmPzlCr6EpjoF/YADbajF5bWCmHz
M2H3QA1YdA+6ks0/hD3IlyIdo0gJM6QDbjSeIwYZSYcQNjaGnBUMCPkbZoS9EvrF
zsQBHmJ8FpCkV+4UbJLWY94WF6qH6mnofGOwhqyGDutFPIJ/fmvCxLqW3tijgWPI
RXt+StyY/AO5OLsMRvCNyWvuWWrO+DJ0/6WiYPLJYYDAmH8AMrfGYlnGe2aRVa65
2U/RVylHniwZ6q4GAo/qz9upGT/s83cS4KL+3qvcm9VVmBIRowZWN9e/OLJ2Fuoh
JwzWV2UdYOKYQsRyEUqECNKXA5RJUinncxkR8G1RrKM+B3/4vUGpoKfiY57q/Vk6
y5Kh+THPOGy1VjL3m89i6o1AhbMBNMy6HRMgisZHLCR4AYen8ukdRXH6WtIbSK2s
1KEcPuXsRTYeCSoNXmBMiEdhr/F457AZElLwjeeJ/EgeA6TBrdFgHmpHA5qG23NM
YGKnsGFh3DTAFtsZ1mm7jLW9W86yo4LeHQkL6vUwd1W+/oAoFkAgssa9hBL4rUky
APsVDkhBMblHiA1TmX5dGmNeCOA4moaf/K4TPpDBe4RyFGE/ZYC4CF25cIDqyR9s
en+YtH6Y7HGThvp9xmGmCF9XlbXwPynaJqbb3H7i8wotdJh7FSNNrOsdFYPw/Yrr
ZrWJGZwrydVstSsOoJUQmNDex0IkBPhzMgCEubRq7IhShzmgF3DeAbzZZeNiQXsI
f/pmhunhf1/dFbrdh3ElZVrimJTyiiPqNuqjnUSQZ+3nYDD5SzfeaeM43wTLFqMw
w0KrNdtvLR6k+l9OZXpzahnhoZ16W3xn+G3GnJ/MWVaG9yNcjRgiv5qsSkdhlrlj
FiJMJ0Z0zDvv5Ziwu9mv8knSwoOhC3yyhvR/LVxdUNMbFDuD4h/YcoNB4KjdoAl7
JuvUKQCiXuMnWuj5vekSntFGxLCCIQXy4mn189tFPYKJ6j2gWRGFXVYjVcsOoPGl
t+fQyf5AFfQsW00CH9Ptyux3o5FVsJa9pEbKgR3ZrfO6dIzjBXBvAQH9fIA4tUj7
N/hRD2bj406HxARgL8CWS6jIbFheNyOIhrg4O7u62XgjCH97oMlQiAbC/xJz5OdS
4iOA8zLp4Wti76SGT3ifKwwIBct8dtCvFQjLdpUMXxtlm1ud7Q3aU78xlqLo+pv/
Gi7suWvO1mq+JxLKDviHIlad8tzEtWvI13MlAeHlZBEcQPpkDmVJHc3wLh9sKEKJ
YGJxydcM+w3nJf3QNYfLizXRycQz3BIObSaluCcYusZzk/vgTl9hYVIWtvu6ceCD
IPzNHy1Q45cUsbXoi8eY83XtHyLRXuE7c8rj1pAOCnb8REYEjFaXV/q4tshVCWc2
SO9jqrGpxVMSpKckrFzZC3TUMW76yrMe6jl0tpkQexq0c8dh1OFeWJGfpUY2y2KJ
Y6kuegOLZSw8dLb5vCQ6721qDCuuIhgT3yDZmfzw9yMvEwGg+HDXetWkG63fKOGE
ASC/7naDlJzc7RcBUv56+ugf9lSK/w1fksozIZ7kZBzhQsFcKGHSC2wOtRRC3l8C
BuIDwZOYuuvMG/YPwNaMXz612qjKbJE4qTae/zAyysM86SYQ4Lf+3MLfZsNKCzdG
MV0QHHIg0/VURC/R13nYAIKrCGV9eFVO2Yci96UhMOWI1oj+Wz8+V6R6eu+PkES1
p5FZl4Ns14IBkqIB9o0OxAmAWMgt1rVfnEJmN2TIFcAVX3K6cx2Bra3bJ9Nvaz9K
+ERK1c1Md0yJS5i8rL7TtWurWYoxAPebA5zvtOpcaD8ALlY5/LvJBx+HqFqQSZiZ
pWfdFEU393a+7vML7zzZoC7IZJCAQlPSJTOxWjLKaAs2SsPBclmnVpOfs7EVRj9x
/U3W2HyoZU9BJ9eZhVnwNaS1pRX3P7X0KyCw/31f4CjvxdEtFz7SP9bSJ1ytvUoo
9Yln9AvuucfLcX17wOyuepgy7wUdRkbPZrFCMXRkN8LmWM1z++rWP3sz97kjXiue
PnMLDvnEyZ4M9hsAHptwgCsHOPOZh+LDNxyDzZCxqIZ0gP3wUcLKcfD5pA9wbc9h
FWJB1RulxcqRU7IhVyJ2qwuRkoGXdoR3RHrKrsTYOnfGG1XUizm6WbFCTbPhW8Ib
4h2cPyfqfsoACs8E9AzHIFXPmfTx/JjDPW/OwmNgimVEPNuUsHhDHHfmcTRpMTTE
oeWpb43BgLkeKXne0hRtjvHO85R4L8JeIsTaO/Rl3xdkpMy1xW1rEQ3RrsLBFpQu
hZBk2V3AUmi48eS9KXHkMuca3APeD040YMgjqxA+ekKfkcihlf1KlqqdWTVUeytp
Egd22UzrzJoKz7Cj15BwRsCmbN/l7NoHggWJN5lpJxRl4KW1HDq8l6YdIenW/Q8H
N0Xvc+y/bSDNysrCpC1pazjMeu/hB1ZYx9mRxnB2D+0xIOjX/N5NADLx1glHH9xe
JIIhPimGTZCe4ZwaU+IhWhyYUp3HMhg+ecSCFcDWYlzOYNUdVLPo1D5jzvikFz01
jOdgbVqDr7xCQ9qAg0dHmYCK9tG8rBCRzYJx7MOkGBh2xugHBznWlYBLPfugMbP5
Mb8clhEtP2kCtjreHBwhtB9/vRBXBjc9BaoPuEvZKiAWnGJg5uLnffRcNNR2cQfE
yE/RDqIgM0+rh/osUUAK+KD4IG+1Z6rGQ9Fk3ma30RDjuhfnxhFbgEonViHlsDH1
Waoc/fqzUhBoJs7LYvvzywU4ASILeuseNGQ4t6poNSA8+VVBpPp7QDAwqKAM9zAV
Ig9vN672pkKsPXdLMiaZu8+aws/cKUy/RM6ZEnUon1bdFCiVhXkOo6vS4aMROocz
ee6FgDHEi9gxABd5UxPhwKB4TH+wozAuY1H2+5t0bBcuf8VnqM2tnR5VcT4CXq0B
eeK0h8fq846lBeEmTQ/jQnRp/JUVAFqj3VrfUcYEMreapxYIsS3x7Ud6xVAaW5Ha
s2ke8LGAHdUaF34h/6wmaedGc+GZYheA6lPfZQ3ggfhPsgC2QlQNZA7cqmvnN9g6
eHhIMeUnpy/DPl8CBkZdgx5cHy5UU+0omS+ZiiUgYrre/nvBdtQ1LHKiOv1fSShl
n4VPid956yWoBAC1LoZYrJQe6LRLpS9UDxLAaDsJRz7/HCuNk8/P2uiqaUyfIqXP
CYYLPQeK3CfwKox5IBYG05R00jStT4RUrXKrstKP1icNFhDcM5aUndD7ozRZUR08
AkQU0CyMmVMzX0n2oB3lSlT2VACBNjhk6owcRSCDSzEA/RtBoUk4IGzk3zR6CdXY
pLNBq/Trb3Ehq/wCx1xpyiypa6XK2XEh+lGysgjaNbnijkKzOpPI5de77SoKSL08
Q/QNkj2zsTSnnd8yk+pV+45CgH9mMKQzRm62DMg5er5CQghNsp8TYPLGxamoVAIJ
0SvEgHqpcjdDbhRa/ctcmb2IHiAuRsWs2LUaCFtIz4FThnrYaB7Ug0GrJZl+Vev4
XBpkStI5yDt7vZa4RlkP3eZk6uKHJzqBufqSFiDvs4McVbyAGWUn/tcqMrTfD5Gj
QMBuJXsvrvRdXVd4QITXCgCulUndGR10C4cANb5JCwOFNsX5Mt0NZ/pdhSrcmfEV
MzOixxslLPqdytAUaK31fwbu9cXlxuvDrlPDTfI/6I0RFBOy0Qi+lG6D+crPJIT5
nj7p9KWzX0Fo7XOR+WDqYB2kHJvYINwYzhG2dKLVOsgc5BnTSsYbBaYL7yJmxqVu
mlBXS+ucPWhzFYdtMk3abWLgVlXwvUAhETcsue1iav0SOPvegWuB2OLYMOYWPjK5
hsa2AArkA7JwArKjEppl+QgLzEbsyLCB4AaI9Z4rSBmFA/wxzlJJ9FReZZqvdj2U
mlkVwwia9mxMGGnowNu1TGmjozQxOGNfJtwzz0sqKwJRvGXTL9pbZJTq0PEtVgKL
DEH49L0eTq+WGP2W9Y3cvp+vgAC70ZfdS/sR/WTxb7AIaLLAF9O+04q0VsRqB4nY
zkaQ0dye1N5NdaiLEnAoIPVVtkQuialaPLrjtdjEHOE6DL1rCz7EmAkJW48gD1vJ
5YsRO6ve8QEcefHwEr0nIq7moLmmYOTxJOmQYUi+nFcYiq7+/tjdriIt0fwgnvX7
HGjGgnl6v8uvROb2cHUUuQpQiXzZrq0v/lq6AHfBpQgQjKeYg9QXv9zXhavbbbbn
94E+Y3415XYt8Hs9uu9lFGJVJ5b9k+0jv7qCgmAXul100MYhtpUlzNOFJSGWHhzW
bAe4DUWlONoIbame38XV3s2W/NSz69dK3LJ+cHVTsgMiWjTo36eBZ3JUzaTZfz1m
yRV7WFANJ/rAh6qnfVQU0G9OjmxQsTLTf/8V/fsJ2XqVgIHDOE9jrlg5M26PK8hp
XefNH7vW4Zxke++HcLIomn1RzKQ1UhXdD0RC7+vjz7Yp12bisDDbDUzk/irT9peh
uGrBf/GE1MVVexx8SM/YIPeGRNefTFRC5enuU6tyriCa824m0d8X4hoC2jW7IRYl
mPoIZVyL/UUDE8QrKpv3JT04BBygyowhCdYdr2ypPXWHz2buLZucuh1ZqPlJwEtL
V4GeroWlQ3KQb+9CMlZWaDUk7pXhll0I7VbfR+BWmjh9WQCPmxeLvO0aGcC3FKDE
HSuibdJT9OhtAYLl7wqTozg6/T0xdZolNof9HME/oeFbSEfFxgvbep2zvw1lLa9x
6F2KSyzFw6W/KeHQBzWtSvF7RD1CzOqYXjTOyM2b1x86QyiEUp1InRDrOljg+k/f
Cf5UBhTX3ZNjiCUZm/Tm6TP5oLJnoqf4NhBE/9eZVb2dRFRAAcrLnpDtaeL1o8gA
d6uj4xprnYVHRKeKysF6/26pgg+7FHiwG9D0L3Ixwra/TEN9GWN6J8cLG4B3eMhm
MOcGtgs95KRO4e7kUrOHl/l8r4Y4LqaMmBkXhB2g0S99NQhO3WMtWE/8WwxuFmqX
yxL5yARsjC84K6gpsFcCANKYkk3zbpjfb+dr7E63owVS1uzDjZZ+6NhMd5dvks7b
VgT/q9mhVl6g07OuaUK3vEWBYwKqK4i5dyqiUh7S3vN6weUIPQAggMAT36Gpg8Nx
5JKemL0w2PwV99wzXz/hmVuCBBsjyuPNDy1DofDqal6zs0fBA0k1Ejzx1piVHiXO
M9QREeWBvd+XPHBbQmS2f74a7BfMxtcHgAOih7Q0oEfyv3Wq0jqxCc0lWu17FYYE
mk3bb3bUAGocWWwolRQRN3XRIF4XVrlH/c7bmaMUTqOGjH3eS/2GiiwosGEwOwxk
TCoBYxvIxmQuALZ3yFYZgJwo6BJFrNuqQkkR76gds1VvdEaBm6CogoSHRjluuWrl
bXsjXXiRQykAsYXtrRbboTaUgwR6075ljgxUekQoRgBaJD9tLuk7UDhemzfhlSGk
aZr/uVjCP9cHWOsguzhFdxeZZJl4uRaGnPoM//ygHrAOxkSX5SdkxAVIoppJqmYW
Hs/DJyRXQ4tkia6/bgNadhBpTOzt5CCS6aUr5FHnKDsB0o2PxP+/hSoE2LSz1W9t
mOCsqW+J9bbtiDg7sZjVV1gcn6GXS81ZtICOh2GaCmRRqJcIyhrnrOOecGoR0QAg
7xDo1hmIXK9NeuX49Hy7qc5WjbiUb9j8XK+vQZVmfqkLFHzNthFihwB8O/ZwByvS
nMvd61RZwrKEor5CHh/QvGFeBR69ZNMlQkUuzPmbwhcLffwLuLNt0JRgidflGGJj
LaNOvzI2+eTA9WPmZvs1+emmfEfI0lByc6NHUnue6JXnaAx0RH1uTvrKxa4yZCon
LSiIG74B91ZvUr/Yj7IJJs+JPVhhbdGllnehEQgqwxwNOkZx8J0J5NOHFx8OAH5L
TE5zrUAj6lvHWdaDYU9uXYvQFz7rC8+a5oz71pg/d9BxOEhVahiaCQpFUYhbfPsT
KGDqifSzB00FDRj0nnpjzO+4p3fr2UH2glfRInGHE67PVmkYr1UoVRfsL9Su9Uv7
gbyGQEnR5mzv9g5Keg/8Yjy1a1uhAIOFUEuA9W76wHcJw6UXRm3ISzNPs+bnjBCh
xotyXimdddk4/D/8hwcp5NMpQ3yh/rOpIdIbBp/eCZrqlZf4B1+LA9QJsX9M6Nxn
ctoBOp1t7AQ3mBtrR6+jhMJNwwSLLxG8mOZ6X5mZ/RKFtk/eRh2I56OtURsJa2qe
3TQAeyc2MePsoeQm0FVuG/Yw0epF8XqDXJZhJxXqOUXQbtNzI9J/iRgYQMzq8eYM
NaUVJtvqwkepmwZmVpY10udHCAPbUPevLr80J20YX0bchXSikyhPDaEjqp4owC2l
9gmOzbgT+U8dC0TO5HuefgZEFPtHbWwGNxMlPx0brsrVIEciCAoVSfQNM5Ak5j8W
SCK04CyPs8tOIBkieeyfYAQZgcETagw9nVJyfIpbz3rOZ3qI0vDQBhJi2YXL0mMh
YfyCijAsV3Y6DFzJlS/9uoM/stszHjrSn0WIK09bdU84fR4zMbF8uxBeGsTULL9D
WfZlNtAesCD99QqC+MJrGJ+illgI8lp0WBDwZLgH66n5WBg4g/84xt7kOZ2Jm8ah
wuiWDSmwRUkM7Q85ZNNzyAPZLrTpWo6757jwBVU6cp5/28bYzsJ6bNvUF1L6vCIB
Qw5MLTGde46ASYQRkwmSmVRtnHk0xomZDCXbN5j4OuLg9b5cYwEtq7g+1vUQES/T
A0n+tfCgZXL1Q+5jJyK8KXcq29PHTVO8oGEqVsX+f6yNTCVid5TBTYL56H1qLEsq
nV7W875mYFNc8fsGt4CtmOqK0uDtTH4Kp9fWYVGBCihwJ2BBJbz6BgG5gxnh/FbN
LYtxZk3Bfxbz9ZakDKhWpLMP8m3bU3C9KE/3GctGCHtYNoEH0f7mmjAVF4nMQtn4
I0JWupDC9qM/ihJvIpautTKmbG7VGIQ3w3HBC/0p+apF39LzVbdG8c8DHqG0Wexm
JwWFahThAhNize4ZSFUrQ8qXCVCEXfQKyUhxGslrz6uisocXjx3LlCZx4pqKv3b9
qlk0AU5vN5pYzI+m0eGBq62AKL4CaKxXGU4XQut9Fz8Dfo1xXWl4zI4Nvw1AKqoc
Vrs6IX8L4hAD/w6oOxa4xM2kH5c6VfCLAGsGLUZkME13o6ami22z8+xS7hq0zhLp
p9l2qmk4N0JGHMp9wcDdA4IxxF9f0mJBxsMaiScHWM96fH+sWqqlb6mrKJI7wjdF
2LEFyIjjAKI0zUC8lBZ2vSfP6vSD/OBClQfANbarNovdqBI95HlcTnDIZYm0lUvU
VRTRnCsEDMBjECI4K5hdULY88SZfb3UNiJNTrNuJwVJ1Jus8Kk/Cir+NNViHkDIW
HxRjMP6VOV/B37FsRtHnQ7k4DUI5pKFoeBTmyQI0lZamzVsA+rfzF4JwHvRCFvRf
Wif+7I/EUGjHCizmlaWUhMUnu7V8IrKcrDNDcAZLByk1ltESGMjZqfmGQ8N2V1O2
Xx215vGL9apMtUrAR/8lEDwXDDCrNnxU/Bt5WQ1BQbYHBfGogvHC3hptxRVH3eoy
C8rguKBqX330JVeJbuI9gKqkr5AYjh5f/8VrWkSr/4fjMIC9mWtWdO/SfmP0a1vS
GFi+bfmPJbFM6AO0iqsw/ZguUgmpMm4CDwdnfrsH+Sog3Jb5EzbRI/7GdpWo+EH5
aihsv+By9eoDVSpnlojruaZ1IYaWswZPO1mi15zEcu3yTnX4KphUdOHX/7u4n0Z7
OhfWv1oa5xpbpGO6R/33B8fzQvjQmqvDnS0oAfD59hM8DpK2zpJTr2vw15/dEPHU
o3RVeeGfclsLoPIu0NU55Hlj/0mIemNtHwscUcfSNg0pcqTMRTdKqB2sviMMAI6S
P+2kamkPsqmP+I/WV4MPa2dpOTk/O18CnYoJvRTRXx35tEln7Tyf7LS5JbsRLXRt
JyMHaX3uaK6EP0Fb2aK4RJI52DmXP9wLY/O/EqAxaVNu99cCi/K3wQ6pO8OFLVXd
q88gnCbcyaF5yFwRVnwtZX2/7VHEMEERWKSxby6MWEpKsxg9Wh+/7R4FEQ5WVmKD
8JhMQfEWGXresUZ38wnpKLc+Edj+mePWGiKQnx7SYMRFVjYP/4g5uFMUGpelWuMz
BKELwYgfFEu8u52RuZa5sJiLab0CdB7zkImCUqYN6EFUm/eNHnAT+cYePe8MqW0H
zM5jxEMr4+OPrxBukN/vbzG/VR+YyQdBN0QFRAAfqk/oXxtzYMCPE7gGN1/Z7ZY8
gMj0XThwlRBm0hUvEYE2W7T1FHlPV+wjp3mXJgDCPj+5cL3OjD1Rh3BcdSMIlunf
6yipDNvqp3q+jfMGQfzkt9WwN2Lomh4gnhXbB2ncxXOQmnSw8al7ItZFVIKWVXaB
aKnWMXwwy4079HdJqy9LMTZgl+LFnLC1MtpMLkgTOws2La/EHjzegBiqifTIGkQ/
fBh46GMKzq6BD07BIhZgdj3AJoenUGdTbjd9ayS0LpQsWWX9iYLvgI2U6gnXTf7e
cuqCY8wAOGdF1lUukhGvqOVdem4BT/sdBwpQ8fl3LU3JuHpDYn1WsTGs2YNkZlJ3
qNVzPLSu+/i5z4OitZLSgPFmV05KvWX2OD60Hg+w/Bj8nqWg7la1ohXK3tFTpe8k
SofbLiSFLWVkFY/6ZPPOLNV3V84Cq61T3JbxOTLRTRfP0xr+Yd8JuKatXuPvcMif
4cJ6v7NgrkPJfF/4d7WCduCIa74JI7P3cAWWkNcmYEVUprHsTxm4e3UEdr+8VbQ9
GL/bPawMfnS7Hk7oyh5qLZYJPuLMGPZepA+7VVxg6KhLjrTJVW918L3oaRLBwVmk
vcS9Lb0hHORQzgq7e6JfWiIIOBIs02+B3WSJ9DzkNXHzFmBu+VqsriyrQxb7Hbg+
COxwEQYqdfNtfhGJ1aGsSrkbmO9QZVu0hoJ8rkWYAe3fLt+2qzI+IEHLnQAmtufP
IO2djaWWQbC4NI5fy2J1xEdRfP+3Ayd4minOwfqDuJIrInpZAbtdPgCxQ0r+Gn4K
wi+/Le7eTalDUf33v0X4MEami6nO3LqUloGbOeil524nNiEoWfaelZW2ozxQEvLI
pYPHRhCQZUA3kahlVGefy1ETdkXtHQZ9TDzHmDCLVueFUjl4zv0Ut9f21kqSMbOw
VkWgl9Y9aigYFw5zb5g0s5mHSw9dxC2dxmFD2ZNrNxp1kHknYScJkJ9bzwrpr72g
Ket/5SJzr7ro6AlbTMvPb6rq2WImYUZcXqtwqTI81eH4nORNzmWmHaJxkwVk6uMV
bm74rfHWZ4j7A77pDRh/q1lt9rGgv6LyAIO611aeSkJg0E9L+w2ZPGzJfLHwvCI2
NSmtwVHZ15MY/2sCncWMCOnEB4IXLW4OQMrovmJ7Dn8oSjr3LjOAP1rV1vpiSPNg
icm1f3iHhsiCObGugcS2GFXWl1yrFsoSpEGlZ/gIEWpWVSL97o77uEY1AS/py7F8
pBYQ+cTVkkvt3q32kn4idWhWZI8eepgqB5ABoui/+oojn42KtZvSwtIx7euaA5bs
T6wtypF/CpKLgf3BKaRPekMF6OnGj9smSdJkFy07ZbIx9xJAifrvkesk2Nja6fdz
rVQBMA7RxTK+yxK/eRmi0gUd75upU2X0/XsvAWVIz33hF4k5yhuA2ojdwAaS9+jF
Hr4rdhVXHrxwYdOkVd0YVEVjCAaD/QUqtx2b9lLUrGDZOT6Q44j5geD/zge/uFfA
AhdL8Dgy25jHQau2cyX5/iuzMX9dzWz3x9lUc9m0KHP9DKKM4f6hjCldP2qPKxJB
2bKtmmuuew0qoTyRe8Zz7mVGZX7qqlIHxUk6aCG1WQDlUie1WAcyA/O5puL3ioai
L0h9OFikovkFqrp8w7MwZx+mDh0sGC/WxLc0y0rYlf/JHC9PBLOkzVbUJEMnennd
HbXjZsDIS0loWsSUnIGDJLLQwTOlTn4V+WGKQp7btTQxpJmUglNrh/9A5Ad8BEgY
jyQhM5l2cC8U49ljALuEZ1uNEQI1dFGXfKr2GqPmB/T11Ja/lFMiI1+s+kuHh/cT
pWHtzv21mssOd5FNJhclH9+wb9fj2BdNXdb8a4ZDviPiiRiTMluJX4Uu/e2GDhLA
tlHSAAxNlIjAhq8TwgDlDcy/6ZkjYrVpnDBTEB2VHDcpVSdIG6PH4COfGe0Cz563
8w9vTkxFa7I54vXJkpKV8OERE7U/G8jM92y6tybr9o/kuLfIGiJwIEaDXFwOZCGM
ym5w4LvEgeyM/0FUoYhufANHL6ThpWHav6QVWJrmk+P2s9oj+E8oAuqI8S/v+nLn
H06S+Qzx0t5oE0SMUnKAn5QynJj5yv4+680djptLdQHa9dyi3NlWtmK87WLvTTrf
OcSUyP0r8r1J0mQL8uVcJ5rpd5Ye9Wra18dqb0TLoF1BA7CT4rJ+MRsmc3ugIxDo
BEUrzkd5TlHcwaksKjaNDCA6Wl9ci0Ql6xGAp5GjgNSxw+Bjs377ihbHDDlsFsNH
K7xwoDJR9C9tWZlLJhVYRCNv9gduI3bJih+R0BjSeK2i2YeU/tCXoaj+1trnzFzW
KU8y9XUcW/CiA9tQsQOCugNteXd3lOueXA6RwpDGyXiE4xuLhhm3qrV537D0ZloL
d+R5Ncbx4CBsvuj79zN4ohggWCwnSbUoyFgFZGDNEh3FoILPO4QyTZa4WrTp83Nz
7tw+TRF5f/TEWsYSKLGbO6vy4ZSvSG+acNZbEGaqwR7mZ1VFeGLWKOhdovZ/Ms9p
dDu8Db49fL7WFVgGFn6umHogWZc6omAEkBAJuIoRHCTOA/16yaoaRVtZj2fZfQkR
n6rNSnTUEL50NqDKW8xMbiitsZBwPTYdNwDS5s6xk2vQn1S/HCgZGTSPCGQriq1E
2zVedHE5ISWRAgTs7y95cs7XnsA85P3DAsGSWmMlvoeSFREObpFxXjOp7cNx92gU
nCk3WamUP4P5qsBroaO2WmoVawRdnLrmqHEw7chhnwclz6WIKTKEgt0UkC0Bna4h
c+EiQfhZHIginCnEmQ9ZwxUqD8VLPOMsaqhdA1tT54/vyQAmZ1c+lI5KJsb2tFeT
QmoKgh6zxfTBse7m/31HGNBk3b44tSneSR+VLSXgDEtMhTM1g7IeB4q2LFkIx+OE
Bgd0Toj/AQ+OZVkaKVmcWPcZJV5zY5po5+S1zD1b1qUg/VvKH9/5ZBWB/ZqWtPHZ
ryCZ0rbEnEzG4WL19LrGAhMjdclO6WhOQlrvH6C4+icDaj8KrWlRhEs1zsMEi2jg
xpepUYsOWEhsb7g/EbZhsWpUi5YmZ5iSstCsat0xy1N1mjdxvO+kNDX/bOuNT1E9
ljG+8bKzdlSnlnxznvRKZcQPIC8dR9imkio591wiAJS9w3z9pBBVq0xKK2gaLUKW
wEJna+pW/Ix44EWf46xTpmMV7I2YZJMvCMz5/z4ss3BMin8CfClnyTumrTADpH/Q
OPAbzQZUvYfsue0ETMMxfvO2ITw1qNBVw9uENH9n0OaFQ+RzATwdxJHr7ssOEgn5
XXGzwK1ZUwwwJKJwJCKpZIQhy7GAH76ZaVZ0fPJ5nyFA6iZ2uZGTpB0TN7I0a4FX
WL4wyIVkrJ9CBWCfZmNR0bL0Fus00Qio/BCSOHn+AXl1cosmnb1DFq7oQlx4bd6e
m5SGeX2tgIrsX0au0Us5SS/SxvkyQNtahYo1LFKbowKXP71VBXI7/y3KlQiXfBDy
I4Z7Tle+WHF4noxs2FrhzJ7bPc6Zj6o54IlAUM0t1sQICcHTvrXZS++EhR2Q97nK
DkFulyBORvFXNN0T7XgeKQwpTYDiOCTKl9Y369b+tsNKjykKGBvKpgkC+RyMyxgr
Jfz6HmAHQxjs/IZ1ma0xLwuzvOU6kVgKi77KQJVq1Rwk3o1EPSux2qf2T+JPSiUM
GxIl6So+zECPy15srVt5KQxaS4KAocyAj3n1V9wweveiY2osj4ZD6jvUhGf7uWP/
W+lFN7F/QuW11FVv/VQeLfkMOcfQOfkKG8DIX7AzlNhWY36RfkFVVEhiRNkeCALE
a2kcYpCGAWxpk1p0O53X3T/Yrom3IAXgSSU7tm0gS/AUHqw8TVzNzq53Od2RVNKi
Fw2oUrxjC8MLtQn6JVGWtCL/0MRLgfXyCYuFFw45NXoweyb6WYE/vgyPCbQik/lD
8tOi8sPWOaAdjQ8FJnildvgPM108E8sHgiA9J6dsGHYFekp8+R+gORl9JnV9BgBe
y2DJuV2JLyEbAtEMf8bO4VK3q6bbQdQI+PLjdzfNlHFu4bn0eLey3Bw9XE2bvopZ
nG+D62WmzM/KaNsM0Rwp7LedMduw8sU1U/AVtWOzvTqUHOBt3JkQ0lfK05Ocu+Qp
7C0VhTSpa2kPZXtO9L9gCpDS+HCyic4I726CWVdfO9nI2mtuVm8uO2baucq/FlB9
kGl9OSKQSK9yeBFj8KnCUV+Z1tyjKCc+cxMTW3MIZuzNz3gUSnZRy0fNRoQSAa+7
B4dwnnkq9qMHHLF6edl+tnu29TVDElnDUSomez1gseMdTFfCiRUahxBRIh4dkdg5
PjCoo+Mx6lQcniXTZwf/QjPhBefpR+tPBktR/iw0l5CCG+rG0PyxEsTLPsxq8Rl3
H/ZXy4FR+N7Qn7LC1vrWTjpOchSNqTy3Fqn1yJGW6IAVNdF727OWD7Tq0HeiCIms
nJq8uauSnPBFYYx9GxsIoWGZ0oNNpmq+0IOVo8Ph3bSVZAW+ftdI65U1kbgrNtT8
CIdSCL1k7hyB0Psh93E0xusOvNb01NkC9b6hHzH6hdUy6jN7C044e/8CsX7JnjF+
5eYAXkBcJbbfYkFyadBY+xhzyEg0aU3SzJ8fnCdHzBOtdA3t4Z5vWgMC+5CZJuMj
y36bo+FfuM8UePHuVbyiUCnLoCPIONRSabFKIXTET5RZNtSyKL7AShbf39PAkOql
`protect end_protected