`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11488 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
N+AbGUvfDpEoMIf7wLov5TvhRxvmPHsq1S76utSHakf04yNnV+OyS8mdYLiAQt83
0fsbyiQpF1k1aK1vSWWXXEmXOHImf2zjePShIiEosa/UDFSKCUpJ6oJNjHdzuPCg
PY1fL4Ib9N4GraMTld9sEAsFu7xBCQ6uoXDoUtkAiVWDWwD8z7VVpbVnsY0uxjb4
iT2NhPOvqEFhFhLj1Dd2Encz3kqzI7u6cA+0d+59NxgpQmY0ygIJYmvcY78+UZ/c
Cag/ZHL24jpnHg24LU1MSzbWC/Lw8WnxK/BlQ5bGG/FHQkDcwifL/E9+wzZ6uybj
x0nSvIMpHrXKXZGhSbN1Ch6+8Oz9SO+vy4Y3IiVTSFxecdq5+17UIkYp6UPjoSxt
Hvn4uC5hZi8SCM7P/VD/hbdXAdGe0nEhnRVFhNvejAD+1EpodabvHuapmTJAVtin
R9N0yj4nXqSBK8SYjLk/IDkMypPNIZvkduWATErxJEBXB/8ZXpw7tRb2GFpmS0W8
4Uu+/lFESiQrBOWmeJi3mw0clP9LJor4aAUIZj1XsQTn4N1Aq9vFoUeHP40kvniw
N/4ZD3tyUmsGPfsFpSgZKqqW/IvvWvEq2odztzgzKGVundrmFTnBJPNN8tnzZnEi
wbP76RaeIsrzuzEUZXHQf+mI7zM+meV4epXKEXkrjB0aifeuUXlJ8tvwBkVecCWI
PA5ms1drrnFrX1Gvd/3g86HyZycSzQKNbuI2MVJwv7FjnAOlvtibr8/l3780Ef/X
MUHH+gLvucH1LGqeqRenkyhb/zH5DFe9ZPXjZbz0J0R1e/gJP2/G+am3cE67wdIP
ythp6xCSOMJai9/R+vTQb2poYQo1DSG6wHx8R4yCG2ShBd5LY/921M/Pt+lbfgGv
4SOcexJIHVqYi2IoYJ73K3DRS1c61tyPZttC+a6+PNe8Hoqh7l3OT/cUT9dKastg
i6XTqVxyxrkRgBSt5IOwNy2upWsicwfZlbDJhgFBKPXCvm+bAo7EHEWl0R6M3pwe
y48OQ6XCHDi+xuJgN+rN7PiI3hcJbewpJJbgz+KhodrU3iw0To7l2ucW8vGTA/ON
Pbr5gKjtjDN3H9K2nyfWwQ+3O6C8QlpUUrOcP3gUmcYGOYjzOEv/XSUmwCOdfm3c
zRGx+5bRv7vz0wSc2ltYLY17oLrd2NeNQuLM+MVdJzBZZjNQde74ayh8Z2KnbbOT
XuhBsx6V9uck9hqrDvx1uj1UD+0zG5GRXq78LHuO6TNTVD9TsVMU66pWKKfWrO1W
w6zeePhv4LOyFm9MgMm01m0K93nYNSXO5kFt3LQcPM8xiiyPL0GqCahNJ57FPNXv
7Ct81gkbIMooleY9eRuMxAdMsJay+OYh/03Co9RVTJbo+pGVjuXcll1X6TWIFyEh
Jfe2CN4qtZhWHJlgIYt1BxgglevT70GJUmAwDA81NdAyAkENHY+pt0uDdkmbFCQj
s/4cF9hX9ysC+RjglSi+opIYPyKemn5ukQWZm4O5vBHc0WqqnDRTHnWoaU9AFkIw
H1JXYo9NQOqFjrb2yYYaYnhBZVqtMDgBCm/LxruPgESgLxr40cE7r03R/R+FlFRH
ra2e4mYsD4ouip3561V5U8hY6qmbvzZk28ORupnEcEoiO4/gp4d2optq/5YmgERe
mdDQZH+3YaXdr3lLRdK4qUPzJYFNtTyVzlsbcTsemn8KXgkC3ao/sAGfG3ZzbP9B
7ptyIqjo2DQzIJ4sd+93l602rKyk1gMh4YJC+H2UpyUHYWuN2EXsQuqEt75o0UE5
Oq0jVpv/Y4SvvJJjor9UZD/lBSbhrX9RI8XKM8hC7DQTPvCj/7XUH1T1DDwgChbM
SdVxeJ8w+yJeVkcPKSWraWlK7BLAV4HmgluX5pQjk3abcKrt7V42p4smQbkwuBcz
La9DwfAG9LzAsbqGOI6/D3sUVtOoaVshs0VGZIQ26NlAvdPfwXeB6zhkZjCE+Ys7
j4GCOWnzgoOzYKwroIb+Z4FyTqhJc++P6xyXKlXCtdkV4NYwAmloPGXw+06Gjs2x
GZE+5BsfSqHre1T5asOq8ADp0bLfHoIZIRyCZso0KEG92r72qvYwGQP2zsDOFuAP
7D+CXAc8SbxWXjuC2A3saaF12t4ke+HqCzbo53YCJnna85W3zH3/+e++B3xX/b45
THXeYC0/yeh0Wh3Puhyivb7vWCeWhMKxKITgBGiS2iu62fYCxEQVvD5ngoEYIDk5
aHLR4yHjUqqSgR/dj4DwrFRG3xXXgTferLLpeb3fdmTzbv01cQGRjDz5NpoFJM+W
rs/gBesgP+Nc8BD6JeZIWrGlRpnZcgoSfma10UBT8nn/uHF+g7Xcuqy1HzXzcCzq
e68rL/GGtnYfRl+J2mr26WDxdJGB17C47bttL2QZIkRHRp/7AawTPDD64j6apW1G
Lx2jx9YwbZBm1suQu3fkYEX1C7mD4Y4mH3To+c9jKaDgb2T74Y69rijCrGrnYrZ2
zcnORW5L4Uf3alNY1fxx1qDw6HdTLj+c0mvEdm5KlD3Q1gDML6bJxkFfjB0DQf2/
lcQqUAuvvofwxD9BMEMFuLnfLau+HFKjN/rH3flO2A4HLB7WpVnvN4cnODzNtLSI
EZuvOfoc6LW8i0iDrDJP9ShqfLBaQzeXfFH7oWtv7iLdH7lRf6CGO8O85l6tis8W
nxSsOg3rCnWS7JR6DKc/hrcuQkNkfRmqNnUOXxOzKCqd3h/XlMFIeTPAx+t0JtWH
sXLPPAOY9EbPIXjMxnpmNv1z9PneHNdUHpUTDsXp2Cb6Hp0Y7mcQeqkl7seFFt8L
BtXx2q70A9nkMr97prvaNQdxv7apw0IIy5NzLGCjBzN6qz4yMBJvOgMp1VJglf9j
dOZ4gAOEdmyMTN+xxJLbTrwhJF4XJ6DyG3VJfn6jJJB7HukTlViOF045YrcVuki5
+8b04M3cgQlGOyFJJEd4VHQcsi7akaIiMVjZBzsz6VbbSbEpeVdb41TdEhloSjVL
9chBSrm1RDjoooxdY+fbJw8kUmpnVwOLU1zJIEeY/y9nfeGYHFmQklZoAi5KLjZk
VGVxRoDbnqvzbe5o5Ap/5XtNti5gkKqc/En1qSb4Wlhw+ijSp3zZaLW/Y1l7GRP8
SlHvjDHVt7KIV26DayGgkN0asLXbTUSWr702CpXjKMsHj1wsa5kY9nNRm9sP71HH
CNqSoYQf10zzY6QyUUlWIXgqw+cpJTqY+dgtM6NmtZVtRdyN/quv381MecoDRzP1
z9rSoulrcrJe0KxY2WAvjy8q3TbthckCASEXi5ayRnvaouNSBJxk4e45dLXon9dV
/hd+CphAu22SVGktGwYXc3Mmeco9fSH/8M7fXx94vNpLHtVKvp80Gg39UjOii9+m
dnzPl6kiS6yom3vfdcyipuwujNdx5aQy+W4HvWDtXdt1Zh728kh8BxjY4GTlmZun
h18U09GLwpPHTeOEz/b464lHHniAaIKQD0BUXV1rkrC9wYIeiTYqAlmFlcfsNPrX
jVMdgEjlhej6elOzPDW8yo86IWypdvkc3sxzm3jXtgaF5gigCC1H9eO9Mngffcs7
rx3gSSCpfcbuObIEOmOqApsxa1ceUjSzNf/Z6JFW5cHkQh003JhyAeYGwrUzhzUb
GtczhAeQGJF9ajDPycNDR4y0q4kO/jhnrwqJyJIAzzTlomZF+KJqPIfGKT8PF1aC
0zatW4Nom2boGUxBdTIk/fehBz1gXA03nELNuVc8gK9PzCX7roDc+r7zkR7lZcGu
2s/x4DWPcu6wqHkkstCM8AxTq967LdT54Q7t6umI47qgYrIXfqrtXuOGA/rKwK+9
afzcfTgUoy2eRcsu/fIRMUuF8Y0SVhejQvGeWcmQ6WkCHObixD+pc5KXki/dR5Yo
4gNDSxqcxFNeBKv4SdqP/eqWP5iLOcR5hI26GzixY02cPwzUTi1/jANQsxdVlACw
8SxAONvGxiQHLefsTVRA7DyTFmDP6GVL4ogzTUgb3WMJ/Y1/rL8oZqYJMVYBk24l
GoWPahyqtMcvWBU+qZ6szfAgw9LXx1sbyFqD1yPJud7JwbwPeKgbsINR0kFdHL5W
UaAZ39H4yUZVy7weR/+GKbFAYdauAGBComYTjPkZYL4I/45tIfMd8qAUJuJMAkT5
9PUsNURPBxXMI6tlZn52fkn4zu8J2ubp1UuQmgNru8zz9wgjhy47X+fqqpB/9G6L
8T+5PMFF7Pg4Brtz7596ysf9orxVvL6cgPUXWGbmbaShRUscJmHGM1nBVT7yK74Z
LkXX3+IB/FxpZiTkMpBcY5/np+XLtu+j92htVmrXY3FnzpnI40KW9/ZC/L4uqcMg
gjKmXCTVnvEr7Mr7qgbOCj3QPF81uO7938EIxO/1eKJ39g9XzlJmHWB3okbQh4Ls
fFxwbU9LLiSHCSCkW3VO23/iw3mxAHhtlbB2esdS9VmzkK1jse7S2qEzA7PU/u7b
ojr6ZF8Kwa8LS7FZ//2rbUXU3KbkkZyggs3p7YCzQfZl3iRu+Qom8G2KOsfzQ6vh
EBK2BWw7BCwyEAB+uWlnt5u86irl1eA8U4/D6y+oxPMLECdQjPPh/4LSwKoDa17T
WD+HbpGftay089wZ8ur7GywGjBtnIaZzTk0uQRjHW12+sapc/mje8f7s95/ZaqL/
kCU7/hAIO5nPy8i87XYRnzzF6EKt9HnY2jdENSzUAQ0t2b4hQZNezQ5ln6mHUtNb
ZmyDO3hvGWge/mHq1w017fC5hwZSyJQKee00Nh2rdfadvw9BY6/Aaoq7d1u2wTsc
szI40l6808rtQGJUcR9+5ULY+hVEfUOs4UcLhNEOu2WeJI4Ab81D6u/nZCGS5Qx/
CipUs4hvnY4lgpZLK7JUKIEcTgag2weDWSB3udIw0IwV9B3dhLlonYXKKlVwqfYs
v6WuacU0AQzhObyBE8/39RjUQ0YaaywRHaGIeTa93I81m2HPbtaFtLw2ZK7p6aCs
NhH4OkCm8hvuQ+BdXYYCPgM+h6EUtQ8EaK+pxNVQ1JLCUa/pj/yu8qybT8J9URpS
djUnZqCbz4h4DBlaQpp0UCMT5RAvsN/3t9+cwsEowQgSznzHqrFfdLMl5ig5I0AA
FkBgB04/hG4O0K4zAS9AN9/jeh/HgkzZT7qyTttYRIJFe4nQrZJHxfP2/jBoE9+x
ZQHAG0UicHwLt0S9mYo272Rw64JSr7Ez0KzuwKcF+TcuNrDDN5VUpmVcsj4+QZsH
O8gZeSrKw1n8c1lor5VtCQrA9KqpwxOUcg3ypbDmlq6zP+fkRSvK+oSnFV3ZKfGw
DeeRC8pnCDX46TOUy5Rk7eUMwBY23J1qA8zFGuOMHLVmdEg6uRD+DZNFIWp98C0O
a7bBj2e9wwD1QSptQgcsbq9TiJZtclDO4t9EL5yZ0OEPw0q2hRvQabjxNiwW71nT
wJBov5SHLOOvfpWDOSyYM/+kLkNvhNbpg6r3d7zA8Ee75qJQnRdcFFbzKDK0tdjb
j5FcbgDUCrwKCsCyvaeO2uDYWGve9uXM6PRce5AdEZawg+tbSq8AE3hHaz3Z+MNh
wiVF0tOvvSHWx+p0QovvilQCBJfnX3NHPP9G6vdEiW3gdSd/W/CQTdjDM+cgBo2Q
JUrw/pPPvGdw2mghtL3TsRwWFSB76fVR/7m8g45ftQGlPF0hSbJBYGqJhnHygWq8
LlNqglE3yi+jqu901UbtaBsMaFp74kW3Ek2f4JieBshJ78C+NLikIq/KxoG2x9YY
ulV6ZciPgDtlhV9c6aVBcJiPWSja++5bPyvgZb0V9AMtV4d63y/J/P+Q9MggRK78
4bGNxtaWtXGRcIjipKxBveBydcDTgzOXtVQRG+ktC9Tqv6vmhTHFn9xf2oY6jGD2
7PaNzM3FrXqQkP7/VqMGjYJUp+1CL1lLY4OHJFSw9t640Fg+ME6MjgM8Dqld+rTq
sVXa5UB9KYQ+vrtkjfqeRQCSLIaNiJVztE2JNlA2F5s/HKujltiGmcSEa60FHws5
V44ELLsd6/soO6Z/0frrpiludmM2gdnB83g6oiaUN1ZU3ITu3Cl5VMASifNbli2i
+1DKSxBKJUEBYKnvoAZrjaBPXu7fOssJIC/gN0U/rw3bOAT8lG0iX+MZDTRq3z6f
Ppx+cveChiCkzBaYz9tbYhTl1u2txz3K7HaowhWY3pHyD+fWyGHNiU9sSkp0z1i4
RkzmsXeH0W3vZpw4BTChc08PFc2+eEfd1jq/FAY8ElLcBA5oYuLJo5eRTVDzBwtL
x1HM8HgVJD63Uyqy8uhyZAVokN8XYeiWzQ7RG4O0Ogd1ggLIbuOoZtChY2beLy9X
CkBDdVqxh9P3flud+Ic/PfCqSzwLpfEAJWMfjYMpu9XxZuXP58BwCvl++lfanTJE
Eu7EMQ5l9JnH79PV5FljnPQI10PimSzDDRTkPzgI0Q4krpGZVV8liDm/MPqMRYtd
7nGQMLkP0+On+PhZU/uPuLAeQQOL4m/Zw9HZBMfe9En0+lGEWNlj8i4Uga9yL9W0
O9o7N7XEo3PjTq/9yoqZEsPW1vzE6zsIRlshLBIJgvevv10xMLYN6hlElCWjRq9F
0CBrrF8ml3s1sR40t05Cw/yEYL7KO24c8yXVqetKF3tsWKcycJHHLtLsxD9iRR2w
O0fn9MJ3guGeFg6pIOwuRApDBXIrn3ms8QFyqu4HVpcwKVoh0Jbr5IMVWtY9DMy/
ilDeVAs3dM3izquXomVAOg88B8eBn6g/COYk/JUWjanZfyjSn15+mVUnPWCbCJ2C
GibTIsv8kACH+qttBGNVi1v0RNsRM0fwaHdPKmoR6pF1pdSHduWaVt3wAvTQxl4U
h7luw50L07ThdiI9V5y7fGjTEkXBaAVutAJe4mUX2bh8wE/zjdqjkf14c7eroVZc
Y6lMiELG7bAxQrbTAnu41S+rlE023phHJMAEnh0aL5ZqxWtxReuK3JeVSMdqwz/6
IgMxTD/uK8Qy6OxE9oidFUmQcsfalQtz3dzRpA1NvsOBIpN+5uX31dPI7j+zPphw
FjIdc1kdK6iDhqS61OCV3B+SnOkbAiQsZH99KZxC35UdB5lSgdSFdtlO22m6pZQn
Lq9K1bAwvL25ivYPxppT2SfK4yx5xzDESSWaceqOeAqKQsfsyNg8gpFG1fH59qrp
kuWtLSX3gDbagcnadvFsOClQ3wgrIuT8JPXxoch/lmRdLrZg3mzVns9adJZ9Jrw9
Mprq30cYowT+vTv4AqXvNLR2lj90KpfSnLvfn+BW5KiGRs+OluOzYSqupLzhgJfh
u/3Mkt7WNTFHIIL0Ya3q7JBCIT6YKNwrGbNu8S0OlyH2tlJd19KFt97xAmGinmyw
dveJfxRaKDrFqiqAuoAu4z7DrQLYJMRFELCTkYanpushZj3wOfECz38TqWAxUP0w
M3PZPxQJ0xPzjMyL8dVGyXNTAqh8c3VXuaUZQgqeqwnVp5VzBOV4buoPNkmgFIYR
oBebpG+a8moArfFiKSLB89gss1BBjqqy/lLm1Mc9svDj8aGOz9MAoIE3LVefGrwz
tVw7k1LtwcH0c+sDer3iikfZNga7ZxSo/cf3DIyoGJMePMFZ7Q1xN91IfMcjI6XN
pJu2dumw9T3iJdfPgfLHAD1UxwH+zvkyjXQ1aNts0BsRUpOv53SO4brul8QjPsmD
XKFzGI8TrFV/IwXYPxcJyegcbwMaenw8VVaM5YE5Wdg6eCpxGVItDxUzK/Y2BLBj
1A/FJSAzX7oVo/7HNmitt4N4RX2XWK8jausOprl6oHUXHAj4ZxZNz3MRBLXqCf3S
lNPrBFacJcrBCBQt9EhmAGFahQ2VIEeqrrTu8QFlMVGReam8eWlcecaQdr5BLPRq
RSVmsuOAtsPcj3TklpIaAYQTKnMbLt7tN9lRrYOsaE4nCWG8n4g8u4ZvgHvEXA9Z
D7tLCppyagOb35eb2o7WDOWr0iHLW9du/JxD76FplDegXmGAiqHk4WyS7JAliPqu
viTAzXNT4g1DWH+s+wg7LB1dVdmvzqA+grmAe2XOZ0p8BjjTXv6poy7GTjDzNt6Y
geAHzUzVAv7Klp9Yvi7uTHEgJk5V05xfDfjiCTGguyf916tgh17425xKlOvCgcpC
vzhcIypuZWSQkgX13TB6oNjbFVhg1BF9e6MgMYEieDEMwzEjMFY/HtTX/f/UyGim
DCqKzN84ZXC9U4MtrCYHuZPedftxJNMbuDC/rnPyzro2Rqiic9oqATtJIttRuEVY
cNlhJVN+8KIWrMcQ4AkChY2mdjrSZseIYyQNvi0D4WI+SJQ30c7clvKGbGGwPM1H
xtjM1bTfqbsQH9hs4VocSYo6PrGRYeLSRsFgXwynS6Bks+O4P/cNKwTc1XdF7BfB
G+2X60XysfnqJ3cL5c/PQbITkKNV7+auJJmdZGyvNS8rWt5KRXKe0uh3Q+oZw2ns
EEWwS0gsSinTscWqA8DpBGovChggL7BzoZmpjmdTe7wHKwrJWZ1NTdOZm+jVC3fv
RU4vrPLAi6a12Qo2wMU9FjqnX1JwWuE0uVSv+3hWXmQFJrQFEACGiT9916B0f+q5
mLzgRE5yMVH70Jp8jLnJcrcV76DCl4PS33OaStFhWbs0BNxjqsf33NuOdmBI9Nrf
ynChvIXlaS6CiGceQ2ZSIqn1037jqoz+vrSK5AT8CRtCVY8ReJzJWIBSWJK8Zmr4
WLczMdPBbTNhtJc8cUlaH9N6IhuQZ2aP3oDfF5Q28vSF3eFd7WnxBFSUBTChAmCs
DaW7uKRiWifgIpZNE450EtJo2YX3venDieLecbfLWo3AVz1nDFA3Y3Lc+Wdb2Tcv
Yx4h3P0jhEe90PM2AcOsfiIAlVDa5+Z3o9Edv9nhJQUSqunAitrrdiebcw7p0+uO
x4+lTIUdq0HVvPROkuP5S7L3yFHq0kb+jUL3mvzJq54EZvQgAjzuL9l7ZDW3E3/U
TVbv3pyRo1qLRzJR+StPeJFt7bD2k1ZOFwm8bT4dP+lNfApi7oaJ4KlXdrZ7taeR
LqXlCIDHAs0//SDI2kbrciY4dDMqLdrjFdTktm0hI8RdIWiAj3Px4yBPZRT9CzsZ
bYJyxear2yIyJ3WV9o6V8jIT8icqX9IMas5XDxKt37Sgh+Y39tmQUnyRjiEs9tN2
6ndreKPYSMXVq2omOueRKBNdGvpBKG7RjQPa5SAaPjbueXCfW8UjcfRe/SUFqlWC
XhEirxQp25fOjZ/lH95Q2J2E03SjKk83mDKz4p10AqkqVoqzVOFxfmF949EJAOIQ
BMr7S7FqEFC6kYnPSir02iNobzKyyeITV7yh1nqoikpSJS6SNJtYl8Oo+e2I/jg8
ezCx38yn8Le6wLAtOm+VHSxE3YOL6qfY4/u3g0o6ZDZy2swsvOuWyrDlVIy6zl9T
e2q452xwG/rD82DCbKVjYM084feXMUUds0sEH/aSfrgZXF1Ri69uZCBgOUvQ8B/t
1KLSTyNuGmBPEKBYeBSSjZ8N34yYlckMfR1LQ42xf5Py82P8GoBBDs/4V7IkrK2f
GH3GaQmccuLCygswgWWhXoHIefxNUpnOE7vrskodyDWLKsyvHpbgx/uLfGe9q5Gx
x4+ikapcahMmh8cqm5Yk2v+1a+AlkDxC5WKaWS204QR4RFD7LZwtheDqUcA3C+7F
Yry+2FCY9fvArSayp8duZBhufdT723VLW5e//6VM8X3Hhg3mi2gfjo4CILeVsUTo
4o1z8R3oNo2xDNRaErSdrnQ7LGb6JFG4iCpp8f+2sfXqlURSsl4/sNrbwvUFcMCJ
LnWjGgJFWyNkrK1ZNSxwABUCKQ/p5fGBuGwUq4HV5bht8qUdVZS+iSUw1yuqWKk+
QnLrmCeRbYpdq+n2YM4AC208H9CO19Y/PD0DHdpyfvaas9VWvJRYQvah2WR5WQ1p
yVOk8JuY2SLU3Icq3sQHaSvdAFlJ5RQS46wPYrNnG+Pj1hEQIRRDLecbtcrUa8Ld
SrI3R6wljyedJJdGBPqX//7+Uvrrg6tOGegjks78OCBVrvzB/x0X98yF9z9wOgcA
dhVJUpk0a+UGLfQ23rZMoBymMqCRRjdFN30TF93LWTsLl63AhgpzUy96nCFsq6XJ
Nnrv4jO/wbuJqPFRKf9uO9DKm5ty+in0XnLqgEhMic0bPTrrMXcyHA1VpsnfKOkq
qfMnsGsYwEs+xZeslS100YVhI26OkglypvB0QZF3PW10UgU+kjHDkAszhvIa0WVT
7cQvKYlNIAzhFidU9mMSnuTaqUZSh4yIvqRgHinoaKZWddf3+dpgBTvRVoMi6gqW
8k54tVub05dROHhzy2zUZ4tjHAhz7BAFfmE5TaVbEDST7Vt10ZRVe1DOB/FPmm7I
1LNWdR29Q1hV70223XztuapdWcoQt0oQefY2gMH90LOEhF+G/8/kTH0dgkChNuOS
l3JyzNtw4qL5d4r3JCyNA78y376s0AuMOB11kycCNu5FqzV7RSS5Juxvw3GIZlk4
pNQEAtbKK2FkV9qm+ZPfLC5hTWpJZAJJ1ougoSU/9zLKTMoi4IfQMvLZKxD5fUP7
I3PNM4/psM/eKpkOS15R7RkImTq1U/y4KahMmJDQ7QjQpS8lo7z3fKHgkRmh69yp
uYiYsAZz4u4mK+wlEcIDk8XCWlrECXNDDHDdNJN0hZ2rZc4V/QZQEHTClF0VRxw0
D6rHMthyRg1UEyoErHiBC+avt3YTzTdxRtg1xwN2xvA09hKo/E82pKarC2TpyAix
Gp6mM3arDcMKpDwMYikLCS6cSgJwZ2Ee0m4pNLLhhztwZpXOud9iuzvmc5YE7nyA
+2PPhQOBAREED8HzOc3fb928GMi0XskKKwlXxeLNRb6ov+qchxMrajIc1mXr1svD
3IuiRK6u2LJrLo1ssp9W8+vp6qU0O5gtMbvLv1JYtdRuP13JY4sUuPgLW/Hd6Zqi
+HHv7ykQiwUE0bfevz7YZyVgb+d/xvlkq/4wN1upFYe7Kqi5BzKGTT9t/WWXqdgA
1WuryJXsx3QD3rVY8/wHxvMOax2K6cehbFEVqrUkHSrPk6EA1aMkYx8koA134RzX
BIKOjObZ1VkTtpOBDqyxAcPEWPkb0+FB/7Co9bkn7d1YHJuClLGoYQGJK5XHRwfJ
3OtwBsKjpfQ+iOEyNR/oWTlu0iE/1YdILSITHs/paTITilZvI0NM5BPl1cW8de/p
yZdsiQ+bOk9ZM4+7+wLvBcH+L3cNm2xk7hULGWywLOi1AbS2PF/NCvcAl/2pCZSc
gYZKXqrr7G6tblDlLSZGTz2aTtxzFErm9MtEZowW/bmxhAbXY7/yhLd9FJDqbqzm
QsIOA3ZXaiOEp8UA6IImUsO4lFowk1lDo1rq+t3mAgy9+M0ei94JNdlu5tULFfpr
uzLUXZHR2hfT8ZFE5f9GAMt4gzLVKBtR+beVP8hxpjSxItekRHL4VS9QXjwArVRv
emzWl7mYvmN8AwHBMNxGYXtLcdArsucmjKDp4aIeDaXHgfieVfD2u5uaU1o3EDtO
V166XrNez0dr480TKClNq1MwrwiJsNfl1r64FsCdiPxVVhSGl15sxPTfw6ysIaET
03SIUdQkUbnCoPY0j/1KbnlQxCy0q7zV8SC0NZhFksUPCcN3OpFQcK6X8Wv+UP3O
iMYIXN64KSCtps9LbFQhLmqaR4xjrKTF2N+7R0zHwNjOcyxaizOpyhUWe0rGvteC
bVj/5NywEqo/G2cXYpK2kH4f/hThVdx2hcRuetwmi+b+/azohOe8w9XhYkK0hHdY
F6yTUf5q5ytQbF24Ya4AX3gQm4abmX49gxpRepB1g6MabX7AFkZUe2VraVoUf17b
m8UPbM1KiiDGjKGrR5z22yHNReoXcZMFbHeyOO58FUBWtUGWxFiys3dsczz+0QNh
CQYGlBt6L6n9JSl0C4SF2TQcBB266grPvJ2xOzAGf4kjg21OIB7WNbM2mCa/SSiR
AMls0XR3db+5RqVO8IPzNgvriLIsKbzhB/ETLPX29mEsT31B+VUQBTLsvKg6RdLM
513b3kk5wHQfcLR2bTZGv10d2HHKPKV7wkkoao6Tysg0PhJBQgOivk7wqo5yq4q+
U73JT4XDf7fTFUHT1BG6vEWDR5EKD5cW4gVaTKzjsxSCC5rLUXvDwP8g04F5rV9A
2EWErMPqXmxI4XVMV9Y+BJNk61slamfK74USpWozzKsAWPGpSyhzHx5aWD/ncR4o
uzEvKl50cLdtgVI1wzn5UI4S+sfSQxRhmu9OHsvV9Ftcx+sfw4cUqmW4eFwNLbHg
GfRyLqekV1lMAYfrGUodTflrUWgu+9f2AqustMQ9s8zGTS423vLD5AFeOaMUbtI8
dx2zVbcniTuuVuuD+mGxDpjC0UgwRSILbSBzlUld86E7u0nUTU+dSg4nHCW2ks0E
RztynlgxZp+u0MG8H42l4bzG/uVnHSIKu9sxVJT/FLxAGWrWbozf7cg5Wp0gA6EG
MCHjZWM+QMjl9oeowi2a2BEAjktipacMRMhxIvY2SRm9f3hdaDKyw/xneNoGjo2f
K0TdpH3AfiZTzyb1rX6RjWrSCiAuLe/AZf0bkwuc3peLheLHUin32/W0cjnyrCRS
ZrkINj66FbbhIATM3MU6s8WC7BhjtX2bK4FFTXP57MMWL2NpSUD3Dq/Lt8wVm6WP
UVbHdhO9bCddAsHnaSDlD9cNJaXdXnWErxmWaqnfDXdlVfW1uUJzppTgiX0F2OoO
yabHIVlg262+CeZxftYcIyYOR+G6WlR8T8W0sfL/7c3Ff8CuMJ/iI1dweKu4ckmA
sdmAQR9Msfk17Ctds/0CHbYaXEuhKBxqAFomgShAv85uSKKbmWsDEriDw84b47dd
6F404mmSgnXravDgoceQCn7xVt00DPN+NFphV8M72ajfhTt0gtosuIbwl2VrM1dt
rqj8E3Q3mmraUC3pMplCrg9n6nxxSYxTtg9iaf4JAVjTvp2sBRQf0rHvI6sgVXUV
mTgfh65d0AXtrnzzRqpvlFFOOUqcQk1iCh/YmECYuWLC+WmpaP+ugvdKCKoF/0Me
eQVDTm74cqquN/CFsRBEPNSktRzp3yNcpDqdQOeAPYnnO6tlERqa0SXClzZGuoBr
RRkN9ynhC6662wX9krIN0QSjDInQinCWJ3T1bMbkTy3zb+eHPGG+oGB/2rpy+ntg
+mXCgFY0J6Pu94V9domPP1iexUVrkAJcoAh3RwGQsxK53qNeWv9NmCn6mJNNvbJg
Iw+eXYESUSI2fcz3OQVZzcNMbdeJLnGdr9tz68+gs+XQQ6qqujEtxs3N74d3Hmsi
qQWZXOtkd7R2csGVu6rMKeixv2on2o1oMem3X6mhJ9SVyaK2fs3A8EVzzn/vEEmx
E7CqZxUh3oxYH61Kl67G+uvSZeHeAlSEOaTSC1AOvXMUzrkPnElo0zLgDmrevnRY
R/xkRgb9xhYXYftZRH3X4OaQgM2WAGAQOQD/00i24y+IQkyZURRIIcUygF9K9Uul
3Wq3wzoJJiyUWC2RJnA/g+3p89ZvjsmAQ4Q08ITa3Ujs7CVdS3UwooEt8zuA3i6H
ivBEnz1MbKTTuXI7VL75PVZyzeKKsj/KXV2DAFGnb1QRCthjM4B/hEFX8ZpJizA7
L9XKJpXDLDqMzSLBpTPlFDSXI3J4DlyNPiBxN9+bN+JxuCG6GnG3T4rb9fO4ObRt
fIlRZi+7Q2zSgkSL4AdnQA4qAdFxdqDiqM4vY+b8dEMQZM8IFiSmfne9Zod9annZ
pmOA19RmtxmOSjBf8RSmQWAmO1azxfZyyxFnSIJQ2NBfyXHWXiW38mJcndz/rJzl
rexMV/t30o23lpGTYPOLo1aC8Yy0FtFwTJ6wVPFZAJ7B7fyWSeOPfy1S5kE+HeyR
b9RDyHqKsaYHswca6mCh2aA0SLZweoe6Sunf9DX2QzoxChBG/Ju6WE6K5CJPc+Vr
9YAwf1ipHEJXLTkknWLx9NHIaahk9hA1o1Le8QlxZGFl0mvVtqy0tOLjcMDEmlKr
wAB6dW+2kt84rQS/rS5k0P6U/Pj04cIdnvJUZ8FBsHX66fxB8kntFWENUb1GAVTf
5nwTLCgXNcQvJRPhXotP+IS05D/hzeBNORXbVr97KXdAt3vvpmfwwNNGqfEQ87J9
+We+MTlPcizE54Lb9uISKsSGIl/Q2mCvArW05Gl5Z7WSpu8b8FgIIDNfrcV0BLcO
OhkNJQ2zE0IwPF8/IDU790SLEchJf7dy/x8RzCbKsVL2QPaBp+MTvfyj+zVdq1DO
M868YFU2EfUq3yPGv3syz/ouGyt/yDg0id62VE53tjghdL6cVSicHwbQtliyyPqJ
bbrf+B/AF/HfxuvB82cOyazHorgFadEEFRHoGOm7XoB8Nuw3B76vK95FudcrO6Yl
apxM2qDtiIHXfycJ41iLEXOpiyK/DDHAicxQ8pkEvvkSaTqozeNZe5aN5T+P2sMM
vvWZJw8QeUAQl7CDb6Rh95DoSwrdbOmCkPwYw6kB8g8bAr/rk15EvFqSKMN+4fY5
g/C3rBnSJMP492QD+vrOxCFz+vjQZbgkHAX6qh/GOXvh1Q1nDanxEz0cTTPZPD2t
R/F4qN6j+uss54VIbkaOTm+rxvTXKxkEGpNOyUW5AVlhlrS7/0K2iV0cdTRx7FAq
7Fsz8UcPC1AaoVuvd4R36/BT2O7J535UfeySyF7SF18DcdVL5HeXJlITrv0BjScW
cmIfoxfBAwMk6mwfLwUHTp49jzW+1OsZP7mySt7iRDWQxaRFZKCYCuGxzuGiWvlJ
Ppm7jha/QbM1VOLsr8kUsRXOIshtRG+t1nQob4AXJuggYV7aRfc3w5O3EOs6w3+Q
choh14awM15bGC3kot5gOOTwHMibYHBTO3ew+WyJ6NsOg8hg8cvwAtqqQUTxIZlf
cfUbI1vLqvMBLGUeTrMn5B3F9qpk5UgQtPaymBv4SFwfQV2DhOYxo+Y+Y6fTirbv
azj2XSEYyqaYuZ08jKzNhdilbaKz5AQPkaKinw36wZtffkDqkmX7ef4noe4xIhTl
R0dZe4VDgz9QHBMPQc3VvyJSvT/yA2+noY/Z0s/FfCox6RxQOgT/+kb9hUYwMY7z
3iNRMOqZUrAbi/9sZwI1GwaXVibDDWmfM8pS3MgdMXPSUakA1Yaae0KsCyKKb8s0
EebQ6JBoEv3Szj5MUJ1FIw==
`protect end_protected