`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6496 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
DBGZtUPdvgnvgIFp6VMrQUsnSTppXNsHPz6xaVXsQ4K89S72kihKzKMYudMRPq19
mfZifkr/rEAL7apn1Yt9WLeJJGxhNfK9Ky+KOBkj1pQ9S04uc7IhTiy9w3FHThdV
uPlwThrHPTaktg+8oAK/Qy7vjFTNk4mu0zUV0tGsZiv/tvqrfqq5fLaUReenfdmQ
Yn/DM/tUkPpLUeQdrTlLinX1eI88J5+rzYzYBwZQ1FCc+HBFwKXe0+ebw/b7GmV3
TeD5eppvzXTTC33WPgqUuPC3BJlh1U4cyScm6Gj17xahbqooeiiQZxDyfC2TF+y9
RL2mx3oS21uW8wLlfXqzrF2+v1qc+NiXvRIxG06ZGqjR3oB4QrRl0twtaXH6Jeke
BmMCjgdz7waVqrjNM5bxcKBMYUj8veX36YUgNpnHx+vjBp+4es/wOraniXxBHKV5
p5dZ2/ojqx9gLGKrBy/P4wY/V4n0FMFi3nfmfQ86MaGrZASvUsWNuMfPpVxThwtG
qGxQzYuhcOZzmccJ8M2ecI0KcVKkSjarXq99wBJd5RYIAZoiKwmwwXeGVRsOKcva
wVIpLSD6eDtd18+pez2VSPgucgFpG4JtmQRDBFUX5DdEAozUOo3hUl/AgM/gb1es
Kh2e62hmW5wFfbIcNx9k9CeOfpFlS6QfSc739sTfxPtvowxs706B69PbjF8gkkhG
8bT8fRf+TvuAJQda5/Ai0OrYxObU/HjP8l6IGqHGBIAKuJzqz94XdqhqB7HwFG8J
0DShmrjNNtHM/CmDQRXW6ew1j9f56Bja0l1uP7YZd7qK6F+qt2t8ZgT1gmRbzO3N
SId67iD36s5f2f5FnOfAO83+RarIttAPAWJ9xMz1uxP/UzoCcmIfMx+Kpm/XVBgO
Ncop0fbN63ekcEivk2bWJrhySW2HBsMajDDDPLC1dsrBwMlbNabV82Bn7WanqYPc
zpoKWdSz346sbGMxz8OPEzqD48pdZ236cLC1DvJckogSY8m6z5jCjsWIm2wzvqXL
e8ODNBzGRf916RZj7oa/6dLVXk/QK4Li4xisfrC3SlboWv1fxJ+1GmAzkBVA8GRT
8q5/rhIza3nFjHOdFzEH48eshF71hggf1aGuJSvr1T37MW0QhuTzr913OgQHSaiG
MhWbWmKloEWpuTJYHqDndDHUQsIOoTxCNWdPpXwmDUAGGrIapKWjdRZFtrPwCSzW
cWxdbqu6uq0wxCcXSjvIwYBj18SbFoymb06fs4zRoLlp6xJsVGwQnUELBJFCdlnX
+2BecXbppkLMS14uA6a3i8ymSjAoQiJ1ZnOqzWhwxxPRV0dQrbPk7pDGxoxEGiCc
AYyBTxMsgTcwmq8+o70275lFn/xZLlGhAO6Nbkt3bxXWWeZ5BWe48RmYz9YgRs88
G84eL1IP5AHSdVK6GmML5CcpF8dFADnGPkr7n3QthSW/y/EzduDXuucn5i1pq8oD
wU0Jfn2zzjCUVqRVmZSOqaAdY1wfwWQapSPplv91GK9A7Ee6kvvp6tLq6DjxihUv
68s2e3cY17pQ8R+UShrH42sT+yKigD0xYnuRfH7i+24YflJ6GaVwop5jThrtNslj
0CzIrzSgeFEvXihHs1di43uAovWoaNynB+zGTX+yQOywy0PPmpYgYu14I1xwiaHl
6v7+7byRlvLANRNynS+MxhrbUvekpLPv5q8NygquGwWhFFxgmyY95Ps137FgyUVq
ftEonoyA1h37w35Uu5QtxbJkWjXhw8/Di1hMSBxVdZhsVJZDwKCIZqbqI7szRPvz
zPb2d+oHcKoJt8q2e6uXaQGTxNALCp6IpFBFFXZUYKDw9/Z9NdNfne0gAQmj0m3g
u01EXhCJYe6hiB89jgtt+bUtCBx2cS/qfEhIjl5vbaLJGsWEk6LIR26BvOwUAXy1
8ZhAwerA+lehtnsrGObQlr8tDuB87EnIOkRE/P4lr1m3ldljE1dgzSJX9CkTA0bf
k/1OPrW++Xw+qx/ggv53o1+F/Y9GPDrYTXwoEgU4BWUBetdj+SLZlR+4+Z7HwvKC
/fiot30411PgKni2/DDntCTAlQ83nzAk/Q/JVctoJ1RL5RQGZo/Bq/RqXWwrgNgH
/4xY1SEnUuyja+j0Z9oDK2SgLwi4ttF6aDz3hjz1KIzSB3BO0x54xCWGMU32gS2Q
G2ZSmZxqA6Z+hz/t+5Zo+SnkqqAdk9xZsVdH1couEV914qcoP0oINkTvRI9D1qVa
DMjUdjvEsUPtUAnXe6OqWdoLCZ6QeHjNc4JuRmwTH0dNI4b66J9x5fpi7Fhto9jc
rWUK8Ch8+GTwFYULji3/TdqCyPJ1tbuUFdUQASOsphSdfUr/awtTIhZeS8Z+FkJw
g+Wjv1Wa7K5l3dwE3+yXr/Vb6rHuJY83GOhCKp8CVZgU8MKF4FbsJ+auOtxDWMi9
nh8DmYGqmiyoMNFLgXGuuVOfZMzGDK54/CcPD8bGeEaYg5W/lyHA/xe7vrIUQV7A
AlO1Yr13TLbO9yMASqBCXuTfcaJdpJd7YYF6GlPfkLWkxKrQXeqsQQnwwhO93z9z
2LiZ0zq5OMQavREzhfw1wo774eIKyLvUg8w2PDjHuf+SRH5eOi7kDgzce6e2eplY
Fzl268NT/rS+n/+UegA4AFjRtXIxMFoF0yw/xxDPcYyp3xpQsSXu/SSxFRDL1bLF
6GB0XtHxgYldPqsd/UZ0ZdeHcOo0C3HTpswK0iePtmmVZLWRio10vqUa0T3bvP3F
soKZpzCZFXQRdOLZyTsJdaP2VsAfBQ7Cy4vhR6n0Z2anqgzr9TmBVclvHKOnK8zh
Osex3MUvOLvPxC1t46vGYC+YdQRUqR7zGGhYNhU51ToBqgW5NY6NMWPlEXlm+fZu
DGZC3fmJGWSFY04S6Jlf1jkCa5Povn4cA6Mlt8BvtdMkTyZanOG6iNZicJdnBgPd
9WwGQjL3uQtykgTs72isI88WU70VnJGvFPHGcPEURqH1H4KhkRoCAA3pfnR86YXE
bLpHSRhBDO6w5Ql8KlgsR6N63jv7frpxnTHiIm55isz6efsiQ6AAjw+85NrFVFg4
KNXusxjI0e51vyNUzRFkq4mKCg2Y7nSLtiA1qE1DjFUEJwsBgmjXN1il+8L0BmDN
WP1BWu1tOQDdWOh5MFQxXnFHekqIFBWG0jOw1Ddy7/nVuV/TYlt9swh7XUhdz9KK
gc/LZGbQ8Qmcv/xQr2e2DcRjKbI47d3KKj4HuncxQI1Cy6ZTjHz1CuyVUtcqCgE5
leMsopbfY+87OHMr/tTBjmj2q8Kx0Ov3h2y3bGOUOxUOgnzzSU34KfG2Iqntvu6z
N4tJhnhfWc3tRtH+oXkcmTvoKn0pvPr1qRAm4uxBRDuJ0cr3MMpZeVDKSLGfVgLp
Z+8nxBza1mtsFd8zP/mNQJ3wRn5weOQnMjSqrTAOi6nCsZuspBiKQ5RrUjoP9qT1
Cz8SwFAVOyV2+Dy6JQMmYdCsbYILPC2bqVpSpeOI3hveUmOCAJ8yaXgGgO5Ude8K
sR8p9/adr0puMHd64qFS9XyTMaEPfHCB6w8N1GcW9VAug+bHvLdysI7sgV7NuXok
4YhebrvKQ5ldKU4L36dawOcniPXKLeqfCVlRQCB20IWc76Tno8QEMnBYSKaCjqlH
OKp7sAtxrJcQX5ths8XPgzhr4Nzq0kor1nk6FfGTLKbw4IimUExtUasq6OA1dhjw
ztXa2CZzRuxPdpNo7v5KXhomzDn+f7P9MO0uY5Wc0dCFQ7hdewi9GQ3boFdzx5IM
rx4P+sHizXsZDZyTxdeHkqj6AsM65OQVi/eGLEe55HwKp7BQiZSuG4AzL8BSnl1x
+i9zZF7LLPDUOTbBKSHZyOIcwDF9VJ3O6pF/HqtOx8ZTvu/EcwqyGWhBzjbVfq1q
/n6LQbKyUFSg4ftZnw0y7m8M2v3De1QK12cQZ3enJOq7/DzFkbCXArlA89CE6J2z
Dt6q672wY3uJNzQ1cXl9VC+B29VDuK7GRLOGD36mxN+h1BdVWD2WBPo/Ui4BKf7d
rHkjTo2KWvxOHVZj3DNaSCJLX9ehgjg064we5ZYFDbz/pN2yxit3Ph8Bsw+eAE2C
3XUdes0CXfPmb4x4Fxd0BlxqHJF97O+CEfTScJ1WnSmWSO8Gw0uDg5tSTcoYrJoz
9d2UKU7MIFnBT/dYpri+bwU8mhNw/U9sFbHfWCM+T4AAbrzLcAHw9iOgl3gXVAjK
VEgNf/CBpkoM4UYGqkijo2AoJCFPoJ0j0Ja43RgWiq+e8R1Imf+s6UC4/sBkzKSN
m+JUhFrxpumyVwX/TpyHmW25iw+ydUu2fMIHsamkubfl1ysqCRa0zTNYAZ5VJr1k
HXiY2+IzZ05XZN0gqjAc5M4JOExLXM3v9sIxrJPcLm4ALHQMDMvtfBxQvD6C50XW
BeLs8gl1j9mWhJFy5eqO01K5NeEKHJzXiVRD0M+aZS8k+qy4oXVr+oYkPXdKUaHz
kJ6Jsby9vveUf+fcyXRU5Gif+KxGzFxLPm45Q+W1Q6M7KClj+zxG2BnsYjVGVn1v
cPGMxaDjt6x/QY7vI5L9I1H/4Xe2c1qp6KexdUGyeY5JG/5PKrY5SBnLcfhLIjgT
rVTe91oxh0F2mz4TmQtTKPaXRVv6JZ99tHomMPXJF6+C1za71YmCicQ/4mM/ECU2
PIjTzrABfsCpCo1fmISkbN3zW8KqzmXMAAcSRU7ZKu6JYEes6q0HWTh8YutLxv84
obXyoMdAxQmCc6+SFXCksW7nw82AmYo9fPmkZAfwqSAbcq/7Y1xuRclVvd7WRJVE
pGPm/73IuKhN2o9g7ns6EY9UcesCAcyLFpHdiGPaUm9xv+A+F/SwIPZ5GLvlM5r+
XufFW5Tb9TwDS3ZrAvcp7mIok7Uo6VzkcpgwON3kD9Hpi3ITW+I9WPiEK8w8IHOs
B/JQSO2aORqGHgcgELngKJ122aoVOLyYDt3tPKxvvrzEG+/Dm3oqz9oMz1aeGKR4
0OUED8iUBiHds6dmCuEg4Y4hIWalS1YirJySbxIYfPm19vBLOu8C9kYYWmn9NVVs
BdiZiO35yKpdlz7HV6TRixG6E7DwrJWAqk/jRrt6PbK9tMcuN8wieMPUWcWLqjtM
1drXA/lyARersJACedTJB85rsrogcz8LJ6aJX8d8hgVHfrVX7hnTZ87388qFjWSp
ichFkC6chHDg2iP1Djr1u2BORp4Aj2eCf9VOWj8PX3ThM0ZRvF/6aF+cJEK0oeSf
PFO0Iq7xVb+n3K63k2MXxOAXAurl8vAiOjhxs6fUrq1xTMAoEh9/MNRypkkibsAO
pn0OCwuKnequAfPvnVlh/RUNNRUSeFK+fA2X4QnwmjnL5doGOSyPfV9eFNFCZTxe
wkew3Mc6YDkVQQqUuLB5nqhgcR3n/Nhr5TWFbThjTCKj+D1EhAjAdy4BKUYTbh4J
NNlTXhHQ+cb/4RWoqfgF5Ur3gds/arlW7G/KRtRYIjvBq7l3N71li7QACBf4FUCG
9GqH9TVYw1eLRoqeQfDDEkGrqoAEQJf+jROcHHmDfnwijXfS/fNvaAzf7Hm5ZO7q
58NCWzwQ7W2qoO1aa8nrSRgn5Nces0lVkjsnOe1j7xHZt9TXtTEk50WP9aaJkGlB
bwDW+jwkQ0ZtWsKpIPTG4yEPJRp7421bpSudQyvPNPBmDB3Slz02SqXbFaRUOorw
pT1xu1lD6QoZuDrMC/KozR5M355lbvAvsT7DZwVwgm24Sdydy0hJdywdHzK718hk
YTfkE0v3M2YMrhaM8E+AeJl3oQ1EJW1/nI0E2KkQeEmRiKPnbSTRj/sym1kcZ67L
8F0Np23Nm6U7Ut2V6LBF+MO2mXvzLt8IpgdWlp8AVs3nAvScFosuDUYiFTzeYLVG
Q+Ed2+Ff7jR9rLB3Oggi20Bk/CqRuK3M+PJxJdwQ4DCdnUTodEvTtdFHDbLjfnjH
MV5mlKeNfGd+wNDmRjVR7CIuB7DYkpkzzfwTCLJ/zkU6wBoEqUwo5oMEoH1ZyCKg
uoXWjpFIJw7O3/bjdlL9DT2UIdE7GUF2Q12yx3ODqTdaEKFU/9fvRCKZ5Sg6vKGF
rGN0Sjp7vZfCuyM6PkZqFZoKaXv8FYB283toB2JdKp7vKGjNN//fSD1X6SXYDzld
jEBp94kDNjsLfx86xh3p+78gtugx2ITNclXTiiSzWNBQcn/j8uNQ1sNN1C6t0dHm
mfC8eyUvYYk4tZaBrj9/Bp2QBypL/gfgvKcAAuo9k7HNlry1xcO+GYL5Y5ZgOoyl
zO9whIHR++rWUrZtfKYuFNJR3FvC7ToBPYbJc3HLqtwSkbdPOjJAXcCfCbz8mmaW
Rz2hp3jNFLqqQKmjUZCF3ut+HssrPXA2qYQpDb9g3yHeq7ne+Wkp86Z/tLI3YUTb
KjfrPSUIJjFmGlxvS0mv8QDjiTGd9W9+NE1i6fTL60OVA5q+J2cgrIREEuQAp1T7
Y3ZYzORBhxwmqLkQH8gYWXLB0maMBkZQU6X3tiz/2F91PXZn/RCILypJXM417gKe
BEoXVHN6nq2z9gG1h5Z9YLinA4ekzkeWSKI8HQutoXHa/aP0V6p2HkFqN7LzR+Jo
sgjP/tG+RMOfdKu/YRsCYIHICKBw0MEQSJAomJDzQ2lbM+V8mUheXRgchZwGwpT5
u8BgnN6xjHIlWUbXfR5LH47k6rj7HKbb0XtWwYRsI5DFt6LjcNjmyGIRqBB0dCRj
N0++Dk6sNaBy4Gcj2vDDXFYmaIEarsx+6Jt2o4c6Wr/aKw+K8yWxHjNtq8ygRBEJ
x+f/qo3cy7CF60hXUdzomDoXu6AaVnOqMIIaT9eNo+8G4ibWmDR6/fnLjz9TxbX1
MAU2nYg8S1NLeawI7YZFGdN2VNyisWU18xX37zoC2urf48Ctz3SL2VySZ7vCjerA
QdmCVAU6B4ZrFxKeQ9bB6wI86w7TM+tQfE3SkpnOXDiy3rgeptvUnTlVk+T6EBiO
4HquEb4ZQMZyV0o6dsxlm4tRhkjEhbWrAVqmqagBDOLOnHHhx5io2N5jUafLDwK+
AQ53KKaBytk9fCijLbaIspgVwO61OS7ntkxhIc5L4jOalpEcOjkG8iAOg7QwCQ97
kGWbK9bRddVGGR/aKbrbKzPezbKtguA1/qCFi8MH8dJbvA/QucBDrZ4L5Ll0lXVg
dDZ3OAmdljsenvd2U8fW4hfn68YLLaQKt2DSwlgt72X5MZl4qLFrmlfJnmg/4TIn
mfQPmjwDHpanxIkh6cUu0MWc7OmxIKgdyJ3NHvm4IZyVSG8vm+swZ+SLzJFWHroA
uFSgJcy0TVh46rSB+4cEp/f2Ey5KIheF1NisMlZaFv9LlrzmewDiEz56uS2KyLvE
XnB51e+3VVF/Ae6qhj8pQOby4wuTCFmwmSuI/pY5h6hWBQJ0/fA5LKGmax6CB3ED
ElFIVqtwg1lCT5w/AauBxo596TDwCLCKmOgaiZ+b3xe5LYuLrohG9GARn0POTFOL
4dD22uk999JPhIkhQgFo1WaZoWG+C7LT0aMqMThX9yZJfuxqua5Wyq9HaYh6nVEn
C+dIhi29CX3hXLq4mXn7xhbe6qP6ogoBQmWsl+KWz8c1KmPocEFdpH8+E/Gll8Ky
Lc9G2PrQUAoWpV14rfj6swNBfBI0glUSKzzyRFMA+PssvNyxZi6PBQPyXcY1f8q/
6y1HFr7cU1hMNmMHWqPEG5GGRhk22Af+5IEZtdUvxUYorN+OoZgz13DiyqOJjb9y
k0NgAj4+kEQQEZe9YaIon5Ok5Z2ADU/aNjqZCwJUX4GHPojSV3GWXOHUeo7///KC
Wf7GFMPlvHOM+IWU2oBRaJDPVfuOXkTIZgvTCV9V7tQie7OFsI/5A19LQPaZbaor
CBghXNKTgI9OBW0mnvTh0r9Q8EEwCTOvQKfd13NiSjCCaJJ+IOOSPnl9uL88iLJw
lgp83VqTWJCWG9theoIzAfCgdBgMcCUJ3CbKlaboUmqc7mRzwibfqGC7imSLvI3T
5WYJBq7pKle0je4MNk6EvdkzeZp+3n+AXn5dOxBNNWUstm4o1n6KAESkZEzWX0ox
dxguqbO6dT8KAglCLKpAUItJVB5SlB+cUA3veNwNeLP9ktWllm4Z5PjaSAKISXu0
yZCyutXrhxTkpEHRg65DJk8g4EqmSGthuVKPgN9XGoMJhw5DIukVjtH0nFZ7tHV/
KHCmYgWdzNqD1aAYHITe6FlSfjjuKiTOk7LaFppzle7fW11l7gXTcgfDcMehtV8P
NYUrwHAVmHE2XMeKs2kZGYuZsH14g5Pp/VJtnN3li9MwmAtcxzN0Mw8EEO9u/ZwE
E//YEvTXryaB2UwtEo6L9f0OMihKTyv/sBqBU7UWx4iiIDk5oknOYyricbY3WeOh
X9wKJJxubl4ApCyTw6ox69r60X1MpfLJtv5J2kkaTWVwHbwiMwsQ0FuLhOsq4bhF
kUYcVWkFHcledvwMJZWwcNELq15YZMDYfRBOBs0k/pQ5l7EloAWPGePJ6czhkOqJ
S0WRFP81/aj3dNqRbumwxQ==
`protect end_protected