`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 27696 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3b6eMZvf+eQ8z14wALfTJHs
q3E8aWgVMNpEXpVH8GIRP9QKeN0O1EY1shEnU+EWqRX0Jrq7KToDA3j7EDdSDe+Z
SKYzUFQDjBECoCmfeos6ipdB33SOcLeK5MjAnXsT4NdUfCp0xdD6TdTN/ogrtodi
fXnej0ICV67IIOYnaZKXhE2ewKm9+VCBFR0sc2UR/RcBI39E4YPHaaMrj8DWJcG9
Uzxt001UfLeFWvxfvy9Xst0kmGeX7Wn6TTi3SerTUYhTXfcDho2wK2TheB2hzLgl
TJJBzWfF3T9NoCz4wSIokCFbhbtPWp6lLPPexThM0PjuqCblHMmYPgBLTs4JUawS
zXjUZ+rBgqbAFjXFXGQCxyAt3ly9aU6yww7s0uoN5sVBe9LSL0QRpYyl8mhUnTf/
HpBuHxpRu9cdyycm6istJgjrSE7qUEqWhIOLJbgJTlijZK5Al4cPhN9g0gzK+6Xs
fJ85foFocsJ+LIOOokn0YYmxSDNX/SUn7CQHBS4+AHRKZ6KlVykEVHfpg65tHt+k
LAS7jX38RrnL2xGtFLX+rIhDpwVM2/JfwEYD6g+BmFJj/qohxIyqRCym0XWAMpaV
cKGtrI8HB5Fwm/UOvqDsdSg/3nZkRShvXaCBqzDRZ1aO0lsGYU32aAV/O8JgX8d8
IBjhvkMJHGwcL34tWSKzwlg66cEdyx0GUgJX89p2o+A25X0DToenPoUiXfb26rk4
6Ljifv5Qls9tUIQQejI5NnoRmfgWe6CkeooKiKRqcG8BrOKM+JQRangc6h8Q26ov
iisqxkQiZ3ukm6lbG/qj+tYpWmIxdza3CjVELFmYfZTGfkZ49jEkHBXkOFhY0H9m
Yqd7dLJwIrX8bYDxc1IOY+WjunY9Qlnk7bDQ16xTqBRX7TXXvY9qBpOtIMWvS0Uj
b6uS+52sYZ9IJI584W0qVb39tPmcd6XJVXV1h14x5OTT8w3yt8kijhX7fBrbilmw
pYSmr4axCHWdt8/BGn4cPZmiN8BFrzXLsCgg44LEfe8IJZfGlt732ZBjSnyUp1yE
prRET9kP+A1lvQOCWlo+ZA7qgmoB8cbEEP5pM13Cj2LY375A4whmwWPq4Hj0bJeN
FR7mlpwOWw3vyLRiXSn7oBUmd182+rReog6l6sh226m/o3F9Ain2mxdDJbe5NeJr
tC0cbuqMD6xikmdCOuovvRYfUwoC+zevU389+Vv0vDHrQIm/m/zkEbTmGzcRV3LX
i1rlDhbSQq6coBEQUHU/fV6ruSJDzMudb0mA2qXGSYYkYzqiP5UY83Fkokf3XstY
7vkZti4znkAj1ibOs5PFD51Nl2tOt/4Vywtgzj3S3g1amQKWSVFoQLHJwm84j8Vz
2YY3kvvWHgaQGAq+mz2x+1yeILbuP5/AD+GfSnqIuPNBSNLFWS4bDZIgZrRj6aiF
NYtREzPPqg8g5Ab7CW0EWzd3/VTAnpd4jrn5orZIoptouL+08b4U07e+0hFDZd6R
k9xu0mllOf9HzOH9x/saZXa+5uhaFYjR8c+lzScFX0ohi4YpWgxImMQ5+z7Qh2JV
CO7L2mT/P/1TVvcOxfriDb0EfaPprX94USKIqEGmiNIQyNCteNV9Q6vTakazBn70
MtyyjR8gz2gloHJW9QbxyAlHO8JOd8E5zb7brWPLiRk4r539tLzI8vkzzH/xk7kb
PW3wxunkAyQExOqqbOroyvxs8cRGRZlIzefQ25nqphyC2g7kj/4tMhSTRFlRYFT2
cGr3Y3Z199B8D8lb1tQqi7D3RCznLQO2tKCjd3zj+37V/GVHdAPhROKXNyvX0aSX
qzRTWarXS0lnNrZd1j/lAE4H8/2ZPXe3UfRDUOGn2K3LJr9Gow8VwYS+bwCe6PY3
g2ZunW7IoeXw+dqP0PcvQdpmz0z9zzUVZRTVmWbLBD7tIXOiEH481NnnCYQSolj6
UPMB7qwTvxh8oUTTzut+8us5ocO7oG/U9fFp5SkRaQ69ib865WVBulZEyfl9+5FJ
O2swwSpkd0+6xvJ0txVDSuZ2RSX6ZpawY8k2RPhLb8Ik3SMmWmqeKTHyz/uhnV+3
7xZwosQ5ZdrZr3ovwNecR6nvoVezdTMLnRa595YtLb3agULApdp+std69KPcxxcB
urKls2J9rek1Q9takwFsuH7I1IRF16QowWcdHXm1UyR/nVKEQXS55NneBR5io3nh
s3iDGYpWkP7cXIgZCiOz2ZhdM2PtbUCoK7WL98FcMxE5pKRZhmIGaM34k4XmgkmV
19UTFak7liSmaAngid0cSIivv4G2Gte3Yo7NvAUWxCIkKD3P/wV1uy4sX3kKAkEk
EoPDvrVr5EXK3au1UC0aadihzLnwxgAhZL5AVKvpqgiRA1IBrLsbGGdkbh4XvTEi
BSt3tQNEoiRwlmWPQVWtInFiz14R3bUqql/+6jPG1Hdp2GUsEZWKY4a/07D+H7mq
wL2gKo8OYq9gpfSFppHMScVJflmM1RyF4hbjytFtUOpN6PL8t0i6iZgtsoTWrfDk
pOVmBVeRFjOhcIQkvHMIXEsIsIXag3H987NelTYFeV/R9tDvMT2pptoiTO3qdvCc
M4rT8SytfiIQwUvOB06V3RlSzJF1vSUEAkivynzqedlJtEp3eku2vfNAzDKbJrb6
ACzEQhItWH7xcC+pEgI37gKREZ8TligaRYXJPitVNeNEfTmbazyWZSgfhhDcVKUW
B6NC8OPFkErFGQdonp3z8/hLqOgOLwrIUHKl4g2I/mRZuzqUDCH7ihsW59a9pL2h
SxUyvrm45ZEhpdLRZe1JlLG3gOgIQu7gVUUV8PTZrBPZy9IGd66lglpy/iwbkBLi
ro5Dg1y6TSlCFP17gn6wTS0poMNsNN9fU0jYkcmi4IaCca1gVVNmSaPGh6pskxmY
q3ZKvt7fdBpjY3MWgmuL+8I28bYvVZbAWnQw5v6WbQccAEotT9GZCOarCnv7yo0A
WWciUrIB+e96zmd0+oTSkL4/Uvr/uwUh6wbPq+hPV2u5gwe9CF5YHu9ZRh9QeY5l
VeQpfJGz2ghyXQin1Jd9Cx0orvdYrPDE1zXF9542xT4Z17YCbUUyf9MVvTaVkw5X
KiA3UnMQqZUVpSC5K28iBrdspJRIIj0OnBeP2zVMpM0aeRt6YUAKKy7Wp1z74FrL
bCZVAjB7fGQITETAZ3tb5SuHrz5H1Czhi0OMnk2QHR+18pxcUbogSldBTli+i7Rf
hgpzFESMMkteKvNDM6sJ/gSCVFZ2b4DC+HNTurh0qhg7AqC1cRZslXlasHRRAVxw
x4BJN7GjltJdMtZwKtflOyuYOIH/wqsj6WWweoXEi8qtStOUPRUmg32mxPBtaebG
XZ35LF7N1ucz9AietwtEuInpGAXEFFOxmWciOSH7TrTrs6P502fhqYqQ2AI1H4Ie
DHkq1hCnNOaGrH8EUIiNYhQdNq/itwCcqZTJHVVxW/pA3P0FuyfCWiz64cuJgnAv
ipP4vdRnYxRp5kgfwGx8CKsEIj/BIF5355Sd787RCu/WcVUKtmJ7ePRmSt/RF7KX
UE43XfqGvyk/Knrlb2USv0Gve72+ViylfQHj0Me/8hBwAermACHg05ytLA2BoZ7u
EdUaAk+6mvGRuTHfSBx47ndn7nwWcL7ElfOXWQTa1fqQ1/Z4OaNde6PrtsEY+2/l
jCXlx4xFp8M4QodJiA57E/zAsYN0Fm7eHxNsS+3b/gjirnS5FjwqrHlGR8FhrIQ9
VGOrJMy3w1aDjhePXFIndMXCBxyAIbcIOHVag9SCgq6Gvr7mSSly+l2MHs8bRJj7
PgDONXnyF+Lxr/ZHaVUuSzAmbZFF9J6vFEaHqiXfasGXMTZquTZazGUKeLxDh99r
qJ3rxP6D+KvDSy1aoCwx1dKBnXHDPzCRXF78n6fcqhVzYBEodAGdvnAJXR8+xC3f
DddpDH3aGMW+RrlR+A2m3oik15dX4aDthewYGjd8AIbotlOIC2mq+f1xUvR5Aw7S
6wsyJlZiRIsIbROsx7dYM+2ZeX8qLhKfDpbR3AnrwtoIlHYbvYxNVa/K7qsESIsU
COhfQ+dlalrQhBjIQ0NPyW4MyUFcpjEEu74FMalT5vwRMPFxBPbKkRjkhMfKwyJb
0VJUBhrgUkU67xFUU2mIaFrRGJc2jxLb3jCZgOYzbWm6YjbzDnWjsffnkRsJw+q5
ALI7UG0DlH4tDRK/zFSd5TDOHoagYqlsakymlQhR66gzZuH42MdXl8x/TZ4DPbbA
fw1nTIkUdCTiCDLneT5C27CwCJnKqW0IaU8/4ki7VmoqsLtNXp6wjmAQE8iFCwi1
2MCTpgXG8C1evr2nVvf6cmLQidFjWCwhMrEaCkhHGLQkFpUbAnccEIUhhCcBFJ4Y
WZz1GImQCa0Lm+GzoSvaC+KM3Kwi9rbcrdldUD8NLQSLiC/sR0fcJ0lEt+tp4C0b
QjRNYBe/ckAbga5yGUlumcha8DQTczdRtRVjD7ql/OLtof1rikU+KBjzOAyrKJaE
kUYoo85OPx1o01qYtjnrKHTGv1DDaXL5FNTZMZCZCELi376VZy4tlAgLrLrmC2u4
IWUbwj79qHXLzEjkkNDH/ZyHZ5utxdrYm3edBTn5jlLDi2IizuFUIYUcjW+ofeKc
XaoIz6OUJpwODdRIkCjwk0KI58EAy9hMNKjpLhQI8B8y6JKm9UNydUFcxYwiZBF6
uQ8jUDnN96sidcQTBHlsviaZAwDgd0mWlyz+jpgYmlBCJb25GWK349B+hOmOTetL
FJg9wgYSQF4nHCRQAuD0bKo8rAx2AiitrNkuLm1VpWKtk/N/g5AqFfJFKVuj89GD
DLAAaVVSJFqK/dur1YVTU55cH2dgd3tawO/JzyA1uvIBA+rLz0ZNaZfVsbjTMNg+
GBazwHfUAgYK4B4eLBHI0l71wueqt0wYi3SJVkBONOGu5GLznhwIRplTKw6BICNe
xXDx+96H/0wsIayDckO8CI30/Ov0WLBwYiyGqJc79Afdi0trAuHPtmSBlDScwzqN
UFl5DjGGYwHGGzS+bH+PQmadrY0O5Xp4o2FR595RenRTS5glTDp9IEDJKlA5PAw3
D2p5eAU/zKHJJSUUYfjVcMLxdcuzmXHgR/4Ou9xXmi3zJqm+Baap9qPfYVt5aP+5
v3p32LPAFRx66bm+8R3KGpMo/ITsaHRs+8fXECMlCE0FLhaJd87wgygFoiggf+V2
gMqDetXEoPsweOqAQJTPems5eUL5PjFNsuyEaPlXRLnFP3NO6ZofAZBRoar0+Ufv
xmfFTE3ny6AhStCnlioMpMLDTQ0sZs6+Nm4kR2uqOZfr+ulROm2m5o0drGl7Rhx7
rF7eofiErC49FCZX1GNi/QlZdpQr7Nv9VMiq2x7FlYYecNkmg0Jl+CChigcldb4M
mNQ69ktN1GOq4aL/nwA92vsgiIkcRW1tCrdb9ZAKznaS8OrEuLgp61nsagIs7wqO
r1rvpv9Kax+O+RqTB9eBh6cuKMqZ5qZbeJkfFVVPJAyE1IBCwfF7XhrkpDnZV5ZV
xSzP/njCt0EiO0gzu9jiyy9SQlGZxu0uayoRZ8uV2YVm4nwzQy+Cu3S6el27Bg5k
+S9XYITXPRO62pcCm0RoC57F5Fxqs/sQcrnywBkNbQ6os214uJn516tPyJ9yH03Y
PfWsnUns/9HGYpXvk7gzG/hz66vX2/ra9bVw3qMtrdcWl2AGt4thP/rQFBIXD1Uw
TbPiTzy7Sl4kBnIgFFSEpQErMpcsWIMbhXBCXJm/9hCtipIE6taNlGi2c7eEIZb9
1UlO93pc6dOpgdmxlFKw6WQfEpDxobOW/QiN7dKgNMW6iO6faa+vmwmNqz9zt9Bj
kKG2631gw1ncfjEnZ8fsPOfLrbFcy/Ki6MDCU27UIq7nJo4BKLE9T1J8C+J+9Tql
FWjmH1hUqNQE4ckkUZGKPBeOEzf6bytQqMOEkfhiJx0qzGRXiQa3/BTwLjt+18Xw
NVlsb6/j7olqBKkyaPmYK62p3lPHQ6qbpcCER3v7xT/i0Ue7o1ezRFYpvXpgLrkl
kJwMan2xy2BSedtXQ7vxGXKLs1oPDqtdTvdAn9WXcm3spIzpRr/uYmIo5dl4QdJa
dU+i+hpIs1x3d8zgGJ4FFzsBv0saR26ewofJrjrTWlZTpVMf1WELMCl0gZAbvDTl
HcBF7ODEaNsY0CelmZeNhX2nbxHH/01SMBV7s0KcoZxlfcfh39zzOCQ+J0nCl37p
oWBDpqGjqjqVjxDljW+2EjiGlbA9L/ZXxL+RQGL0oXDL804+C6/hdvkdfVO7cpVa
o0Lj7nPNAAPu4uq2r4XO+ViOmbDO1w98f+7MjFd4r/LBDMY1N4iMFtbVMytqqqq+
6cUZzOTWYdDjWjFCBJhxadir9QiJ0Pmot8z7Rrb45V/jUEZlHVT5HG3AKVWx1eD/
1Yfgts30Ge4duHZ6+JUvF4UL8gAKoSfTvS/Lmu0IEP4zPNg9tF5hedl2jIy0m0Hx
/3J0b/V3PnhSVpEdmKX5rzw4w9aNTDfUEP3AkRgvD+pmVwNrV+NJ2ObklYYfG0fd
FMuEQWlPCzIntPLIFvoihihyOzZeCIfeLH0staDKCxz2/IwaB2VijGY3l606Wxqz
jgbStnbQytJiPqcv+qAULoxwWG1QRgG4tRRKkaBLx2SwEqFm/TNJ8z9eU+9IyDgf
jFj5fBmug6lRi8OT63TrVGswlL8UAidEtQuqAJDeNEZ/p+gn2Ap6DpTNQwM0qiHX
PRq9RDJO4+G+ZfiarCHMy5NeJEpnSigU8v0K1wB+/rJbo+Mns9Xb+a40orbAkNN9
1ia+o6kKinukW6s7UvDLzSbvdzyZ43/AvWzWS1Spw6d9MSKU+cGqS7Af/wDTwRlC
3D2WKiV9GWY/A4h8TOBuVOnURvWuZUoIgjLNyfouU8rRWP4AipoAm8tZElwkMqnt
QEcPgfDzKjz3tXKV06YZIVQ9579shzNYd8ztI++sVZg6utRffFGsR3bkalaGamj/
L7LTpKd52t7LEPMo9gKPgC3wUQLL0Z/9oUiEtIbXEZZSkcDBHDiLTkUHaYDirMh6
El+fXwC3a3PawCteXYEwTNNm+Jp8Sd9rGWfM+gnURdY+rkxmBIrKo7jELU5aQ4In
JO2WTCDSNqfE85+NVhXrG6fQ6KMGhHM0Y12tRu08qrvgr7w2kxWCKDDqAKa2/xQQ
tc0SksqbZVTvwPbEzcVYxFLRXRyU07tiVDcEQkFD0yYW1VewVItgtg0YC4ZM+wQR
RP/qcUX/dbDlKbsX+tE9AwDE4JdqXDt5p22mTJB2SEKGj3sTyO0W02lrYPt1CPAa
jozaL0fwER0+I33YVxEp6a5/9gIgbcvi+9H5gBNswWiRZsatkFeLrrnAw5/aH1aq
AHfQVJE6xnCKJV59BExBYYU30TC9+PHlFfN3GnOwWYM8KNRbGv9iSj4WT36qfCHy
DvUch3KhMXlNXnDPw0ssdvdBhFOlbFL1dhEWO19txHGtFXRUjA9wGjgBi92Bhoj6
UyP7GNiaBw/I0rsd+qa3SG7WbAmnEtAo2iIsHNjznOC34WBapsnXZCZAg/sXFvxj
em+GFOdY33CLZYialNDAru7d/cJfcohjJsmwD0uL7X+Xp+dlTQOXj8HMJlyYAyDy
LYC9dXo/zBDtWC3MMIZB+t6PWhyZRoDHDlrbSVvsVDI64clNkc6GDS/pLMiH6WL0
ILFcnOFJqTSON1nGtxLBua9/0ehwjJZGI0ZBAq6Tz39uP0wxyZiM7Bb1qV2PzEO/
FtY1E3R5qTDKObI+v60moWLIdOJIAIUwTm+d7+rj4IUvEaskQDrUgCL6dSWEJdt8
/e5UigQgjvh9NzsXSR691ed6ww3ziLj5F43enXJSe3N41J1h13kqE6R4fwKGrdJ0
nNoeNiJksgGWsRjEMAMxQumWy4bD2uvytvb6070+Z3CPDHPDwHeX+L4GxYniBMQh
9fxgubEVlIBOlPEJj3+qEKyBGVYu4V/9YKFXzhYZRhA+0hXVNCYioegyEPlvFXvD
TE4CRb3vuiNbMw051c3G0I/gDWOWda1LBCVI7DfHPFduwZSBAW2mdZOphhdjXwvK
pdOuRRTLGUbBddtWHdmlBzgYsnEfsyMXWO4JUpb+04dtg5VxJ3CQmavb9I3oPvzM
L2QdzcUtxwP4n6npo/5IWDCCzno/JB0neOK0NBXIWbEvgsyLMrLzfcYG641ChLJh
F3eD2UmQ5bZzqxxy0ZQhgInzXkAyho5TDsXu98NZR0E8o7hGFR3NGavu2IU4Pjt+
LIsYIVzI/GIbkVrM+bMwDEbd7aBOSRCG6zyTnhGzduKf1ALkvqnw9s9/Aoqg1BFl
lbfban89iEYZIhumvWin6vmAxtKiId/3QYuijWNB/ddzQFblblYz7YxNlwaLvaDn
ftoD1axTb8M9KJy9ZJJFKoMCfOXugTqup3jsMQRliIcokJ6HFi7m9lFWotXtW8Xl
pzb2b9wUdF4LDGcMXe2ZmwCPNHXMm8KgHOnRJ//Cd/DV41rwocclbhDCPmIbPFt+
Cq3bYUzL6258aErYQ7nnx6Ur65TrZHUGwiWxbjq3umLs6EfD4EZHneWzYDyYXMRV
osYj0ORmnOJhiYv4R7WuZq/7gvhWXWyltGB4rE/oCxfvCcz7X7/LH2rX+R4MXnkg
yV6fnAfX8geL43T5K6gAvt0nHElKezseQYywYBH1yTwfOdx7Q/If0tzJQYYhVW3I
Z3baOSahs3VZx8repaloKXM1k+qcmFDE4SdDJsPjIBn3GxNc6BTxCzjFyEoFKaDN
K9NKNo1l9EU5sTpF8R81zry5fnb9UurYBbp8GGE8pL09mAI6B4oJI3SqLL+frYKM
CF2KDPIgVfU1C47/skWJMpBpHJuqWjdXUuuv/WOesfAFOF0ysQigF9076UnWqKiq
lUWyz4pHHKQqAwJnwQouJjsIvbtRSErq0qGMR66OBfj6EjsN86SE+AzdNusou1NE
YYR5M5sYizaNuu8lcA0FXQOWH4qHUTwRgqDGJN59X4ngy6XSR5K3KuoNHa6vawqV
u8w3OTEZehuEsV63+PFdLPQ1BIpClamvupsvFT4iHNqpbNtTbVasQTAulDkoR88k
Nzsd7s+nMEAKbzVuctfKnw8KxHsO0Wg5FYNMPEqD43X5vpkapJwvZBKmQ+9x9bEZ
yPSLTfB+LLagDCLfq5Uswlhd3NXMvZGLb3no8cCWfALyF6ACMcjh0m7rCq513O7y
Mf4Og6ZlGUYAvrzotgwFbpNHJtWwV1mc06MlEqIKYWrykPvlTqty9PYM/pAm0DPk
BpSAAISDEVf/rBHUZaOvzv2ez0YuNPQNGyaRcVwSGfzSlqbo50VBd21n0EsLbr2B
3rxQt4j0JRZg+FmgJbaBJuicMi/Z3zVHNSYCkA1FKYd11UA855T6gMTiVc7TVZV5
w+BFaO4aW279OAttTcde2WH+5YlBrsi7qFmd5V3DfTNa/s3aCzUEulEXaG2239X7
Mv9iaOBPpvuJgCDaiJ3OO77ljlzqn604V/Ayy5pgrlflZE5hiwwY8JzzSNZbDL55
1uMqMrj+llC2hrs+0+dX/mlC+HTbPaq617hosN+Ys27pWzzjoptDGxCVsWAYKS+t
EpalsYWYP/d9hledE6XVEEN6128uxspJwi+oFQZf9XN/ROax381g4GNH8EDqyQIV
PGa/D0MNGDoh1T8E2+9rpl/YuMR0LJEURIfbpqYUV1FdK3PliL3YaTQWlyyOFg+8
wpF6YBmE+C9URhhUmGtBdl8uFDtJBHcoHFPQxmT8hUXLsKVyHPUfDSF/uZSNTmYd
fT7qg9h40nbiCEckLBmM9q+9BWNmk8KUDei9Lvdz2CMJANtsuzun81/dGY1B4Un0
9BZDcKIK1mDwjO4qb/JSWDR2u/po40IP+YMDbPShCufoRSFAvOyvqhEfTok7pOLi
Zjotz+mf//2YjMOL1pyd6nUuT+ymt3krL66stpNWlq+RzuzUL1PdiFiyLnFmB0U8
CMG5lsPG+tHNgD5N1vkrxt6EJfA+FCPfNSvzjFHyy4ybkLzkuPLIUo0TaXTucNmA
Cn2kE+l2lR7t0HDrPtDueTkxAB3+Mnc5MLjtj2BQSE0i76gPBt87vp/9EwTZYSd8
r3zt6ZfFlXRXcUmNZvMVgWhppR/OPlT9exBiT56/QsatZfmRjAz3wrGTKHYVB8KJ
oOhNjVtkMCNj4uoaUCVLW1hBgAWs4ARjK67g7HO5IhdmtJgR4jF9bu2G2EH4RYeE
+X+W5lfoXWD9uoIYDvnXci61KiWretNx4WNViP+A5+sTZKSAAXvotCsXllCG/6r1
ueo/pTovDIWW5qNhBhD38VTTGGVWLuCbf4LZqndpDcwSihkGsnC7CzkEzy3rsQko
rAB0hFh1yoTBl4lB+L/aOcSpWpZTD0h5J6xi2AXHAjXm0nAv4HoLeqxmSHNFp6Qw
F+w/5KAvOmqzsZYpF87JOmqsodJdFaaeMF9IoAPsXrymnMUgKjm6C4H1nrUJIiE2
ClFas2FgBMeCm5QfOE/mcBO16rqV8U6xtQ+XKtWr69L3obQ+TbPETnq00Lr2q+du
VI4+PqARzh4NuMPj43t7v4WSvJ7tqvoB98UpXadfYObKCYTjALGSq/DYYKHgLL8/
pssWNPevEaEKpj5611D6dI8nu3qzvdUWYpdwRchvcWK+TISnJ5U8+81FAYlcaweU
SQNZFQCJKDsQ6wdPgZxntoV0Pl3ASTyKfJuHpJsvD/0L4irs+OSpQ5SZxtUT+fLl
EZ7aWUqz5DkK4ofYVVmKbR2c4yb6LqcPRDVTa1LpovznNyLGObIygiGkVV4u443i
U8IsmHhnAW6I55TkXyRlZJT9lxP3rjzL1tnKCn8jEWhgjxLYiAW/aE3ZNzEeb1yn
N6fJFf/0U2A9c1kaNoV0MBQivMgaozU35DFGPRJ057XRC6s44NEUvFxtjPPC3+Bg
npCRGVkbnYins5XwO56h8sKSg0P58FHeMQ+2VlwYqRkCK5jeKtFTX1I7yWa8kGVK
KonsyuuIweSbMoznl0iEs254QijwY5wz5I9A6O9ntYJ+OOCC6tkCu6zPgSB5nGcJ
A4wD0TocSZOzp7HF7fDh41jnbSJKje1ubJaHfC4acR43IOr3PRAsJzAVENODat6Z
LFW3ftLhs7spwp1FJXdQk2cAgB2IvtndwW+SBd3vNKOk1CWQilNyBYCoxGLDIFlI
2Cp31V4UEIHmKBVRrnYUNjchAC+rlwPlIoVZRPX++4d6KdWJCVnRhL/nqZ1hzdZ1
C6KhEcNZdpCW15T0OdSu/gwAQxz/At9ZN7UJIUjOnUcm6Ithblp36B3feTnnVPcR
X2bIX5SVyRX44qNpqQZ0Fq/uZOo4RCPu4wQ4PnQDCN3P4SvktQi3oUAN9a2tgq0F
HXUQLfhg2x/3vsFZbDti5YQH9sst4zrpqx/RjlwAejCbNaM8KYPuoefYp+LGJJHo
PCb1N9CU3Ec5gfLgRa3oM7YKS7viJ1cRXuZtLE3TRzEKfBwMvvT9tY4+dHV5hZ0U
ral2FeYoG/QRl832TQa+QWRgN/6MFLRgPqe3/EwI57Gnt7hE0hAyr/7FND7sLHSR
WgPD2Vy70bLUJ30LXCUCVlMueehoT0hjU3Wa+h6d3cVfCvu5Wjn6ihbItJHd3KVE
aMoLqWlf92L+6Vt7oU5cyzMQ16GddThXp3QjmGREdisuZUpaBg2Ws4l7APBo+AS5
Ntk1EDCK7463UjFk5EsyiNnVbKDdNbfPRwf/t/qpvbliFtCiTKlA91ebF7ulzGja
+O7TNtCg9fk1sftM5l3W54Ep5xPabYpArkTkWU8NiaS+tD/oTrOgNGkbtawp0kN4
4BNI3y7uiICPu89w78kVvo3tYy7WuG+w5pW80frCSvWRocqQYvO2QUCXjrJoKW3h
y8Q8hgByeIUt8xsNpf0lTRkzMLjCTzSNdhi5Nl+TPgUzZ0r+qpsDeZw85YX0DL6R
ee7+6A0avd6EfL8xF91k2r7NXUeu7bAqSX86umgNjiWDmohJyKZFI4duTqHaTw+t
IzCyvdOTUQ4lU734ztdc60vlQQBidnRenxN9UFVXjIBfpeoJgjaASIMzdY+9JZg4
lWFHxnLCfERFRPtwa9RDt5kWZb6/uSMn3Q7zcQuLdnDortkhwkRd656jJETFR8gh
5FUZygy8pv1I3/kmRKMDuVqtvmt6a/gVfjkIAWg/ZstVn/s2nhMDIU26WFHRHImp
pqFTm7O+yUvVxg2XyLqljyQhRG0IiW01zjXA9NW026sQL0cGtmN67LEap8S0k9T4
8h7Og3zc3AmsUQqZP95+jDZ0mj3uad40fxWCak2yiTUmrTJMHQC8wGgsc3CrqD9V
j32msAmQiOyhNLQ63ndY3G80VZQ2DV81rQGVCzT/JZgEzpiOIta5ubIiBLHrKsYR
nBxEuRfhWaw/RQVrf/u1DygYyeJbbI+pR4bCsOnzJl3m8YJOB7jj4PySawbdIPwa
m2VDGzIm33HWR/xbFbculuQrXq6ZEWTT/5lvYPHblqPRR9iqgjAPlw+RxD1UYErC
y9Rj2GL9Fdtd752e3RnYnBA74VGOCHibuSUzk+kI+iVD0yTmZ4q/vUQSEGjAxDpp
GsRHKceCDU8zZwTGAMkMipsqFTnyp30x6vb7OlnZJbRdTyqDziRZc0ERJo0YdB/H
ntALIhu//gEcGFjtDlVaEj1+ZcHrvRVWvIRF2pEMsaOI89wnDnTUgOyoFSdkf/b3
D1bUxsIpAMIDy9BRTwsycrejZc/83q8ZPDisdKGtLApvMk27BbCWF2AsZTr4F4A4
XDymM/2fsUCwHvvcKYLdf9cAWdUkaj8kJB638vG9NIfPnh+f95tDpPtCXND4XjC/
wyxu8gxu5G+M1fP+9t2NpUyjDFHoNTnOXoMkzuCybs5Mw5TxN+vfrE/5GM8v5Ykt
5uyxLvSQET7zTK4p5Iwts+WplicClblhEhO2fK/iuvnI/s5K65UtWOaERxsqes6t
sWULQPgwiWQMEP+Juz1ArZlWpiG7Dvkd8l6CszPVvJCg4etmkyKfQttBlaq9+H3K
3+huz/oXVeVFNzceawhccnfjojFxqg/ulOGEl+vMS0j4rwoErHGHRlCir7XEJXR7
Pp4eXdh1rji6pt+D8nz18WG/yzeYfxqBwCn4WKj5cXBl6B+LQeUFXNz808jc2Uid
fPjcwhHkhCFrxVQbcikSO8e9sVJlUcgzORH3aW2OncPPIttdYuFV3vhA5NzvW91E
CV/gUG7uM3IugERmVE4jPYNwolMCa0Fk2ih6jgQyhL9NaTGdtnPb19bREu2q4b5I
oHGRXJOarXfP6l1N2Xc/wlAHnR+bPFE3Vob7pJmPV//m0/miubu2MZSVD0m8UgCd
X0EDagAk2b05Jitny/DGSiJMC5TF4WwQKSn+AhP86GIomS5Y5Y0zF8UGero+qux4
9qpsR1jfQRgCdAbeGkBnCkDbpTHhQwmNJnTIJHUaB2cNJBHHUYpMQ8iV7VA6QlFc
WFPtAI4MmlUQdnJygyH2kECSV/sVADHEAWRmtLOm/9P0mso9afCcoYmYkif5zAs3
eDse7Aew4rtC4o0L4ZYXYwQe0aZ7VxkwlwAFRIpvrWc79+wbvmrv7qX8ujZmaxkT
BShFjQE0SeLvyCX0CRfqyTF83AmtOrAp1KuR6SD0KNHfaKSfrLUMgNhhOUGRPREB
hDRO2onNEHnv2ja3wiORwCsantJydlGja/yOLp3KhOIYhJTM8o9Sf8fZRH5UTraS
QC1RaLVAMOcZauPl5PHkX10HiBWm06I/1wlLpgMSzIptANoSBOauxCx9QJE+fmE/
CZ/foLuR0dEioGEWOHXHjkB3JLVCTm76MUR5ghoR95XFqOogOfRzi2jZTL7uPcC/
IUrtl6gEdmFROJc35/kTK/YYraDg+9nppmqHets1/IdnttOe+gv1Y2IDPvrnu6hE
YsuFP6vWPCvPnquEoe467CIXHPC6ggdan+x62FZCP6u8Jjyd8pppSDIgOi7kBbBG
OJF2MQXHLYcll0TdrMRTPnAzgneMyGnwG8u2/duQ4PKxnuSD1mVSiopnP2tYaPue
BzMRswagWE2vvKubF7Kmc7lV2Uc927xP9oPqYBGZr9kKVZZTwmr86xsjo+k+P6AZ
NanE4pZusUol7+L5MDnPeYLJHyNGxaBIPfsqKioF+opcicE4pUGQqiEorlynQ6dl
IRwV+BCOIuj0/pcbWUaZwFjc28JlY9ME2AXPr0OOVkj5/RYb9R3s2WrOV0zIzAR2
IRmhG6SuFotx6IV6gJZ/S1FWWOoh/x/h4iHW7pSARSeZlCQ+RQYQ+/uC7q5aCZ4J
AyH3EqX/FhCffjmjDd3Di6M0CFj9r6bO5+foT0tucABnwdcn7YyYhxp+I3IELCe0
v/OnffqMRQVPW5qnDTlObh/xDGhJ006ESrmDSQBrP7QWNNJY5VfecBse388nfMN3
RLrkuqqCin+AQKmVFxRCq+4NyY4i1IJpOqBHmCxaX976UVTPtzYkbyHBLEpNmplC
V2ToS3eHMqVZneLM0rv3qN3jwWDJZR5TIEmmiRuGXdvnRZys2ylAxQ0+bi/V4maJ
/zxoacgP7hUBmI/hb10wMm/KJEdWO78vOFYu1MT8UEaEXe96lWjS+USl98gjFolc
IXyw1Ap1WZLiKmG13qe3T6pTssETvT5o2T0Lv+cVBx1Y4dtIgXa+nMbXs3oC/FmV
ary5lk9iguESQAtukVvNbGKTCPqxGDV9TjtMoQX5EczFSb2/R9xhfvRZligQ5AZT
O1K7tmQIpCfWP9wYEVmkypxtEZsV2qsaFuvLPKaErBVPWlAZjGRl/5l4UoijUxWe
9VMMYrO990oBpVo1xmyEyte9GwHKLw6NYjhe4W/Z/TJYh5qzyGCQ32qR3A5/Bj+9
ZI6CbFeoovZH/E5uxFjQXNQfzOAzngmQy5e62lkpFepN578DuBUPvTM4ZoRJPR5k
BeLLbl/GS/F14vDDA1Svbe0DFYxYBnypSbQ3yA3mhY1G21b0Hz1wHmyq5JlWizXM
zbFsnjV+z/irybEP+ldizrTmDzDDMW3HjhFn+7NhUavqg8KaGJIIfNwcxoGGBjuk
OVTVC0M2cBPDXSiNnmolS5Y7uFloGiZHDlu2/gue0V4pg3LBHYN8KRkN1+LDg/go
vvIwcvsK3kjG13YnxB6vAzjW5HzSAYSKx+SpfRqhtiFFcVdGE3Av8Rz33/ZeS86I
0OZNLUbovfcG7FAQpI6u6WUiEE+IGtaV5udBg4R+UfsrDYeFThoJwCjc/rtT88zE
tJObr47Wn4jzCqT+M4YvBS4IkFN9xoIsQDmnjE3WT4yKiFDro1T5THmR9ADe4ZJk
9PDasxDadeWM2Ai8Xz8RNoyFrkLl1g6ECLxFbI0rhfzyRs8UG/vb9J6eRYqmUflb
TyhZSY7/QIespbiYzdjVsb4TvC7jNJFsGu35w5/JQcD452ecSnMNkzDh9CVQE5Fk
2fcnJCnhCQ3o+Eusq7pGE/SCHWW9YGxLopaWMrM3imRiz3FZGEL5zivuTaLFWJCR
s3CXS0sZqi2SpiMNOoTz/2WFEtVgQRy1gjfNiF6rnuo0OKu0kQgjOUDpiyqPkgNc
1rJcv7l2zMo8htDDsXMRQv1S6Pe34Q0cMAWK/Pi+aMoZlwHVyEqESnUH3+QzuaGd
9eEK5XrBQFreeV8pmWp6mXGc4aKx92YIE5Om4WdgHx+JmUpS7DKJslXSYZnZbjPA
I0SrT8VGnJKBOcOaATgsFQKRkcW/g3+0CLpA1HTosdo9iDZ9i3iroa9wbMD+ovDB
fZfCzzDi2FbFREL0SxLHB8Qd83XggkIiNKc8RWCp5RFpyeA3xV79BwNKRrPNOrIZ
gNAUjROfI6TwW3IOxKWFqRIXhxWnUw73bHbRjKoCkzM2R1Ga2/F7+Ed8vdcg9dgc
6MmflCqFkumTkS0S11QOJbgvsnpmop76LbFf6IwAjAaFBShsF/J5XWcn6TMR+AOM
RNi1XqYHr6AZHn9RV+ze3wC45eaCvT+0WawdvJIzbkMU38QQc/zCmrIH/xvHdMfh
i70CqP7pMAh4J1AiXcPYFFhhxSyUpjJe/uNCuj+NM4Tym+MgDuXMQdZZ7iVW9nAQ
8kGY4Z1y98uvvfLyH0IZWmP2zFnuP+QDSUY2cYG6L5zui5cr9kEArWJr9RvJ4M3b
tJbuoKrJsTxn0rSLDB0gS5ZnD7kWgLGD704jBBwPsRqtI5u54Wt30qm35rx4FUGM
2n9jiLwhJgTwxgs4GSNzJLWTBx7ylnfleJ2Ucemx7/JOMxf3Ux4euY89e2BK0r5H
fBpQpL3+MOI6vP81+yZMPzm8y7QUdA7pf0QRsJFzA+UVkxQOP64APNU54qycit/I
c7XZ4pH+2LNbH7CfHJrK9p8jFBBR4xybX3iwTMz5cTxHqOmdZIxcn1g94cezZNTp
aOIykOWbAim7hxZkgus9ZkH6V3IOvcDWyGhexSJh40LGKyUgIwC/OtcxBH8e9cpH
Kq4WR9A3AlKUFNkxR42qZxZlWX/PxdqJRa2BKA2UzqwYt9vXkMJFUG5qIm6y+Otc
WOy9+AnsAdAexy5ImGj+uYE9AStx/SMs9Ml+/oD9+5zDGAdVJPtfxN7TEHK4iBKf
lbjDNjMEm6n27TBVDNetAQIiUF1wXcmTYPtVrif8XL0ungvYDOAx4oN26zQBtKlq
GU8HR3AKo15aDnIXfQj293RpgSugzvgHLf6Xq8m0mEjcSJ7yPDnfMCl87i5aYeDK
w7jpqjwUY8RlIelg/sLfHvQMMMyc6AYLJloMW3uFQnmfcZymlXOliYkrDQn+CcXl
fXeyIaB5X6N3vRLOj2PV7IXEQfpadST1fq2dVx7CrT/WsfmqE7dtvrKGLQDMrn9H
mpbmr56YgG580Q/T+3WNkze3V0qzAelAvX1wT/rkzNuigoROq9EVfxohm2oaoLf+
xhd13ejLo59fqLfRdYlS60+sm146mqvqcaEHXWiQNFhisBt+xNjcrzAQ753q0hnT
nnb+yYO+YCthi+7ky+Wj91cnC6DV0aERuAub+xJgJxC9rP8rKJfDVRiBv7MoEXGB
Z7dgxVo+ci+SxeGwuqP5P6QZHyJDlSj3jiVvtkbqNPYHye5Uoa3DzHXKOQOAG8iU
5tOVitEEGTHyc7fgDa9Q4o7o3A1qxemzM4eaqzvWVwkEC9iwlmakX2xrDL8Q3XAJ
MaUoWG7wUdoxWu0XG7pNNl4IKP/IdZwlrfTRHS30c9CpKOEDrKws5m3nx1Crjc/5
hgjoF5a7lcY3GIOJKrlELFOjkB8rGKytnrnyt93pDFGNqM/LtxnZAFKmnoO/GxOm
LxKpqo14Q7ExFbdlVN8ydNautmrovusHR+3ikGhiAfWL3auH9snKZfNBdMBBEQHj
UZ8+/V3BHz6wfsa8tE0zrdG8xvsl57RcMUXRhkfDfIuOFOCDkS7qAChD5jW/QqYh
8mkqSsn+mWiTIfIjh6sdCi8SqT3Qy1t0j9MzWZgIodFxO3wzttxfq7k47VuBl9Ng
TB69N5HakNPcjzhqiyQ1Gf8OkrsrgCljhrWHei2ahjDFuwhu0rYxMPit7YEPPMtD
qFzmezxRFlz6syyQ/Hmo9bA12ec/Hg+7NTjU77bfJpIPk8ob0BpF1L1KWwVhdtfj
Fvx3k1+UStiREtZpAbXag9TtzmhCvHm9rqkuEmzYWtnLwxhDre6FwJURyQq/lGmU
R8x0UTSG2g1wpX2XeynpLpT88oM6S5AkQMPI51uiOGr/9UGKPiFZO88ZHJwrBG5v
MY82v6R1FowTihjAFGfz5yIdArmaczhK5VUSGV8P1a2Nqt8O2Ik0LCmWBfxOcjU/
96LXfc2PPOX0msnlMI79Ml8hUZX7i/yb9zTgc39gXwaQCk8N/6B8T4VOg9aQIUdk
ojELkKbF4/UmgGeNqYyFqjp6/F8jT3uBBLYZg9uY5zlziJAjWegs/S+ey4JUSt+o
Aab/TfQ9dqkAcl/70ZLRgXC4rmOW1q/jsZ+M9VjCTCKnw9fMZgLje76gAMRqdKxM
uQlTdPU8izDsLNQ5asqNZCZkplCQgf8Bw6NsVa7EBxg6pnxsc7DWkDUMMqLOKtpH
VRIrB0Aq7+ev0PKuPp0Plx4JOKmcCADmulSxgeoKQmrBDI6wrLo5FXwpO2/VuD5y
dcVkyPoM0tD+BSON/q9P1pVGdzwime3wfb8hQobPV/ZqFY2LPHuIckqO2rUMr+Lf
1qqJ1D3AFIoKgc0FRArNj06QV8PWGre0cicq6XDrLs6WkMl2yudVH70n4Jr+kAfF
bPO1LpGFwUKgBKEBFuClm3rRAU65J8Xh5BXzdexxBbpUAqHB2Ed3GiN3cajG4lnc
Hqqbi9lMbWp8k7hKSFuTJ8paYw61JSoO9k9mXuzZQxytLrVNjqAc0whg0Eegb6vK
qgCFhNiWGv8q9mnuHVepL/6i+pTcbeV0ybWb2bLiqLmzvrK+lvGeNk588x87BYDA
GiZ+SAI/d5PoWtAh3JjG0JzFka6dPF/gDGQd4ld6Y4HNvoC4NTb9HNQ7+yNxVLrA
tWG9N9J6aaMkzA5XTMWwBnla5T7EpepMyLh9L4A2/2Da/D2dYEP7vMG9LZ44pLVk
AKoK0hmLTy28fMp6nymmd5fiWgacaPv6+Q+5O3883qhFeJnsFr6hkANsY/IBLSia
Yg4wJ1Z1Y2co17IcBPXQuQe+gg13uANGc/r7tsdCUXyGQPB9FW/r/fRtREBuneXd
09jJ0lcpYSEwcxdQ4Ukd9zqL7+trQcoPVwaT8sGDjGGwn5o0+UgaFdhcY32za7tn
Fc0tkatXZSWv8JwZVSZSvQniVcMxriw9Js6DN9463Yd+D7wpiYUtL1M+7MWti8Rl
dakdpJoW8OI51AdTH2LpHs+1Z5r/M22zoeKr7iQkSDz4rpUkAByaybELRskrVayo
lLuXsRJP+XgZvMJVpsGow3TKWsq2h+u/J5QyHebs7FG2Vv+UNY/+QkprdRfsd83Q
+RvNiHkWpa+KNdKa1fC8omiaUqHRsKI064IGSavzY/NLP3U+zoip9BmwQnO79c2B
HmJQkkRIQjuGW+61vx+7FeaF+zZw7fXkzYoJpqLzqe6DEXhOURb29jdq9dDZ6th1
x6y8ECxrhXAfFZIT67N6R+OtlyZWtHWNSGYov++KKQBlrcrS3Ydg2c0cHvTsJYtP
Lf04dJBPxyevGGrgRhTnDgdXWO6Xvhfm2EBSnGL8mVdct0TzLrPX6nxwaj5hp43S
qovmCCaJ8M8CVBIv7n6mDvBOVQVkNjK4MR9eGWaPvz4REl1JCk2GcnIS32dN2gjA
tNRbbtxtKoqh5K1SA/2r8+mcCYb3VsMQEsI29CgWA/ko3r8M1ovQhUauW2b41sMR
MY841M9869lR+jCg68o7OLJuaGYayVZ3W8bQaR5PWI8KFDQsZBnLEIzSy9qA+SuZ
XmYjOI36FNSUT7cq9l10zhv/Mp5FS6dS+VFrtOK0JgPpiNyEm0kP03Qz9orb0oju
3Bi1HHTGz4TkxOZPDB07/qN+xJapL+N25fezNfKsyiO4crIvjBzenQp1SeJKOrGP
xiCf3Rph1TVDuGUkHEk1j6ai7E7uH3bn76bi2+VNZjdNAis5fjaZqfZWVJF/Wrlp
PUUsf4tgynfwLBwTXgMjMJR7u+N++I9QtuSl0TXyUsfsco5CEBENHk+2ifupQskU
7ML9goi1Ap+ICo+8isKioT5bZLHuZw8Li+WlcamkkTqmC78gt2EDOsgk++G9hUT4
WYZK/0h/TToqg+9qerOCEE02b/T+nDUxfu6Is+jwm5ywtGjHVZYs/E+U1eU5W91v
zH4hdrlHUAapMUVuEgdczZgGdiKk4NWEUcRhYxDLVuc8vozsLGjnTVolzw8p2iTn
yD3se0wypkWAq1mhc2eXyRjd7wwN7JzWrM2FlEVIGqjAL30WZ39Y/7cBEfcWA0ke
6Rr+ML+E+/a608zsaGm9zzQfPlmTmleN3osWVq/cLsqpI+A0RsZvgNNyWzZSaTBl
tlA3GCmC8DNkkXnjuNC/1OTcOo5pnvkGGgxnYjp8D1MjL1pIjC5utskf3Ii2mJax
82HNPToAzQOSV/WBK8m61/ZWSZ3aC63i03NGRFqJk7Pm+wtyAKQtMKWO8cDvXgY0
oYCl6DZ+W5CJX1MtC/M32w5NBG9Kk53qe3Mdwd/hXQvuGTe6tE2SrrkSgSINvsDP
jnvOFl3C/3nY/UF8R+7BbzFqNklhWwpREGpWrACjM6sAqopiBYNTOkPkVbtJXv6x
qtouwwbdR6FW8LaQuiqGXPmrmTazvc3Nhnil0nHGAQSQZCD0vm7oqQyqx5hvCIFY
F4VRP0eqlpcMR3MtIQGApaBUrMLmvdESVXd/yYCw1aDq8RWpvtJ8nQEPE/KwiLf2
RwwJw0VaR/2uG9woOSHfHajX95EcTRzvQayrV106qgr1M9QvTPB/7p2OIgszjHQv
EehqGY850d4oshDhujyCjA1YM/z125CY2v9iL5NpeMWRPxbydlVw8r8sQUjkelJb
Ycm5MwQLAmyxtT1YGGtCdaScut8KGs/CRO89KXG3VfJZdqNNrKhabRbtaN/fub4E
UnrLmUIkBUgQc7i5+PvDRod/+xKdPyHrIGAkoMn5Yo4kDusvxbTJbh/OwCnEgrIK
xKBi6W9wrSJMpBTwhuru7sKdzxWupdTcPnSvoXRu9gYLKbFdY0qwvhe3bOH1iY4g
YgMzD4tO8Z/Noc8tZR0xjU5YmrXb9nf6uE5R1zWBnN/VsEjQp24ajYzAYAEH06vb
s1EmtSdmEahKw44d1pnnhtBoks2J01cAo0DK6EQWXo505oi+lwypbp9vlkVexPTA
gjHdREGJydLLTR4kerP23qtNAp86NI/fhvjbXag5yLh2ZJKJmaYAck/rKEuuLd5Q
qjJzUy7mRYcr1HpnFZ1Q/SlLSPOLqft9dIRdUBYh3kCloPrTMxDZVVqmp/NQTLsk
1CqnfsEKx/wQsGYx77k/4vWP6o7USxFvL1l6Us5YT8hSn0+dlzzRMNsO3dugY1th
FOcW8kV96F2qUcI+x/dT4jEdogNcuCT79zJTc3VD2S5YdNZftRGOQzKfSDeFMuzh
d9GDOZbHFci+ttzEJ2YQvSg9z5jB9fJiQEUcGlzNtyPMps9GbGtWHBUApENeVTDo
zP54Uc0Gq8PtXaU3spFLQ1uRTx7u2ARW5xpzoJmken3oF0xDekxXau9/vvalWR1Y
zDMOnGXDjDi6VT+S/8j9InaAo6NvejjP4VaacKQ0fdyYiG1u/69jokBYLNVQLAJJ
XoISnDEmzMcDnZR9bZR4YBpQSK4OOnlzWn8at2mfE7PoL5hNq30DWZR+dDIki8rQ
6NYGmUI44G36gB1vxWU0PGt/nrJVRUiB+uFa+tbIfy0RuVz1xPfwMPSUYMMUJ7Hq
rfloNVxbL+m6nX/7niM2sru6HASw6A6Qfr4Hbi9XQ/TavTuz0RhfAHIzcgnhVvpa
YDR/Njr1w8uy6WaU+4vDH9EokXp+J/xaDB9Ay3I8D7dwbiiVxRvnb9Iyoa4YIHhB
M5bM9Pb5IfTFHUP3+y0/O057LZGivhUSJVA56v2ZGVpHtNK4ejjh2uRHgcyke0+k
NywRJgE40PRrM/aO63sqDE3K0O4jQ37O6Abs5wuHjqMEri1AofuFo8wKLOp3LV88
khKmvxDz9DOpHb4WF/6MGB5A/vzScXUBAsQwo6VwpRRXBwW9ku3tAPeXsZQsHRF/
1ZqUjh2LdWxJds7SNGQMH5zdkzISXwoskfC2OgtHmTEBa7eveAn/Hy3DDvblIpfg
9eDwkALeeZknfQt8CV2OgS6UBuCbg+tXjf3eblCBfN5JUqM5TLSnbGWKer0b7jX7
7OzfURBqSeWA5UDwDyWhSfDhBC5Av0fgwvWJf9DA0UtvfqHfLlloDLwFl0sippG3
SI+DDxbxxwyeXdZNjB51tZ5Cy/Fszzt3q/5Fsq8HTJEk7xcZ6knWIaSUrzKpykRa
oJuC+YT9VHKAhXQ8H5vqmvpZtDI1n1+iwBMa1ik1PPAxWbr0M/8S002pjy1iY/dT
LjxumxLLE4xVtXDf7cfFvaEYN10AvX/vLDP1L+BOb+SgMPITMkrHHmGlPDsT7B58
Veky80SCuW2xVtzR1AGwycB2VeWupl/UBwcQP7MCJHF69aI+vR0vqHoqynLje5Zr
yENLjkCS/F+CkDUp1f2ANpWccq3bVOzjsFXv3StIPCjfSzb1pDcL1ElJigYEU4Y6
Hm1uqGXlCsgEUAaUfIKsdEHecxwJBgui2BmgnXlVCQiPiPVkAN9zrU7SCPul/H/d
AJ5moPTDPrjaNY0qDXPX1y1RJ8rBb5fQZa65V0AvQYoJzphYFUAnUm4M6P3TeK2M
od+MTOVcaD1BXW9rdt5WADTe0NbmVLRLUZQKAWsQG9NcgmLe41GwlQGyFLpuhI29
FpapLuT4c1GMeUCRw6uaR9g9sbtMR9sJPW+yDmsz1NoS9Q4N587C9sHEsheqHnoe
QNUgqh8hAzbFaCPbpYXVK4ahPCq3EYC5y5jv1vyY2VdsbKRzup5hMRPnxGjVO7WJ
jkC6SdUd9GLFlbAsbH8wO5if+CM1oryUYJatr1rYzyV53cAVyo+bRllXwuN8jxsk
mc5BxofCb58UzrawCm0IpZQ2TxZqyTWlUN6Sb3WBxnAeOCfxl2cheRcp8z2WfV9k
CZwlPvHZkeomGe7Lrz4PJvzW5afR18thHwoDLgFEGp9+9KxLa59QmwyF/N8e8Dzm
B+PvfRiFFHZHlduXWLP9tH+6uEQn7MOZxuU51V8+imNwtoxQ2mLVIE8riR418eEJ
hxwmRTLtiJqhyfMAxCaNkGqqNWWS9GU05b+SWC1vDcZW5xFufyjzxXc9CyYs46yS
cawRm4BhqbN6zTDwA249nWqeOgY4/hvDz0a6IitWP4h/YDl74HDi6HAC1JDGS8Dc
CwmJ6ZQOyRdjdNTJVL/2UZ1MQ+yOzNTzcNrreTnAiAaOaRJmK/KVS5GxFkLftyOH
0FGHNZoZvmJH4TIszaqyR2hH7R/Kr/Ko+xSHqThKCiEzZe1/AtLucTqbGTzzSyaA
xtq4vtP7G0Dq2OdROFGJHOxzUoOAN9nUbZdShznl1I7/pFm75VrWShnYrdp6Gn0n
m9htESTwZn4V9WjtCweiFPeAR6hOfi03k54blweva+jaPaSBzHxJrfzRp8mRJ711
KTbLu2i6CNfIB0feocxwvZE4wL5+cja/XJrVc+yljwBnu6FiUfMVUm9KztvVR5KQ
leRaxqunBLRir8YwPHbPG+RSvKtzqPdCLkwWL5Z2CXXJ1FvLEu15PvaAsBYnpihW
JWNOuD6O8u+iWSau/1Rbs/zguikWaYwdALn348AvbU6v2xypy7xELG/un39yh+T1
aXq0xrmSXvPHA3wiNOh6KXNro5T7C+LmwG44pvBNxD9ui6cf5Vl/GOTZpZZThAhH
mpyxmDifo8DFH6UV1k+1NvXxnxZcymHC2+98lg505c1daT0tY6Ye9gN7U9WWAfMN
+396L8eAVxG/WvVdVzLGCZ/PE4C09zen1BXWmNQkjTAWlJ/T1bRqFk9W8LY0+uPp
7R0L3FIc/vuEt5oLOuZ+jh2Cm/nYP8Cl2GOQ3AjeOSEck86WMz7HzZk1XBej8IoY
834E70dyLPGO5llNRNcoTAcf9Knikm0HAQKE1ZxwdL01JIMdQMwVr21Xj9JW8ukC
l213H/1fzGCEOFaHMyEVzp/reYaMNm6oIeTUDnp6/7xA65ZEviqqBWnpq8w9ugYv
wE4y3nBic9ZJaQm8Vy8++8V61W2FV2sn5GZA1qqo3YQFAawQwm+Ariey+LylOhFR
kG2aR9UJlXhG0R5q7WfDDR+ZTGtmd0RDap45MPO0ZGEwpvswyDiGjrJhEhnk85Mk
eHU+x2XUKnOIRky/dPGcwXLNboYIsKCdYmlIApUwBdSO6yaSyT7ElhQ8nDmIx8Zb
5ZFZdGmHPaVGGdUPnM2oouVy4nLtfwhQzci7Sskcf1lw3YtLG8sXfd1vJ0ag6U1/
PKWfHwGI9xaZvN5EWXfptnKUDxqEUcwX66PZp8pRWeQMVJBYNz35B7iw1JwHJEeP
r62/UNNzu0cU664sjlhMMd/h5OLELJZPt+jVumLcAnrMUbedDB2BHZcOHTDsGiEr
WGwuw8jNL2EUCBdidzSUkg+xht4XwpCK7CStdnP9e/Vl8q1h9PK126nTPfH+K78F
kQBi/AeGRqKIEt0I8BlDdUFdro7MzQ6v/3h2geIJID9jIi86q1inRv9U61gSb3cX
NH5xjNJL7pk/kcoRK4EkDjFwidvhiZejrHIWNsclSvteNaPjuzHIhErikA6un1GV
URLs2gWQc/gcSsUQjku3Kf3VWEucSLKIPLw52wm3JDu8ZuF1cEjwtkh9sr+bXEDv
EEiVkGCvHNQeXxb2rGKnV8VJhmBXuMIjPTArB4Cse8/nqDfcAmSJ8jE3Zyt75Eot
oefMhTSKnh31gjlTOP3xIZ7RL9zbqOAAjF0wrjVTvLLuaJuDauvZrMHaTkdLpmHl
gQXn/4YWv8WUU5SSMS3aO+EQ2kVSuvsIr7DotCFvfQN0oWEOS9HW79IpLn/KDXFx
ER2JxAgxazgq+v0HW6DZyEncGiir28njoSlLmTD8gqMRcovsIhhO6tMcElqJEc5g
zMnWqmePxJO6v2jJnNFJff5RlVzh9CFcVCJLOi19N3XjmvblSQadiVcjQ09u3+ir
IKtyE6nq3XCEWeie+taZhyvoPt5SuugOawyKkxIRP61h1IEOb8LkvUUaRB+LJ1i3
Ll/HVFpyWWs+7uOB7IEcikjr33h04RfvJiuQmKcuNqyR4tGcqb3qWzxnN0dMaxig
bWx/o0hWRo4HKH2zx2ZcN2Y2AuM2/t+emJQ1krarTF1k0P4d5W+UnC/jzQNfDzTI
T9K+ynV52HUVMxn7aokGXQPh0TwttRWP+yUPkhReeSD5Fd38hw7UT2DH+OHKVaYn
DHk9z513Dl8COwKxpj2iaRFPfFMEfh6YTeOXeBnhb2IiGiJq4Wtj19Af8MXR8+1A
aJEoGX3EXT2Q/SeZ6Ksfusjf9M4H7O+LYq79Hx7RzSXRJyizWGGsztwQAEw2oglP
PD9bfNEfg/JwEjgm3hztkD2C6ZjFiVUCPugjiWRgLIIWqVW7KiDZe92Z/+6arrsU
FfUDaZEtZNpmHLALxKKF3kEO9DOz7QjV5krKkP0oHu0WM4o9NKqPpEvG3rKr9ems
jp9P/jlkyKPsUHAVoN0GVhLqWj8rdxKcTBZX7kCOO5yy4bDrtrNg+bjIbYq/0aTy
vt+zW7A2GOWYURHYcbWFCpgQR8Su9cxO4/z8nVHC3U1wEgb+gaDIoXGehbsG20T4
5eXFGdYJjtfsDTL5q8f8HEh2CosnxAsU6XkfRgc1gAN4CP3jYaGRx16dm0oiEl5M
k9HYqGIjNe2VzDvP1WnKaQJUsEBUAmNK5Z7a1N+pkqlVx14qi1Rl/u3PpKFZb8sM
tJVqFQufKtyqUJMEtvXybc/y9d6DQvDZw8le36bnQcrq1tPLzfyqMhduK0ZIJOnd
fz0HW6PvQnbEcraJpCRP0lLpAhD83W8pvxRj5UVhZKIctRpG/BNWv88ncJE2aNKX
JxQ3mOtkDdiBj5ArWskLA9W9hzH56TzRyj7Ha5NytN+ycD1wiUPCMinxsVHCyQXf
wDxP5LXgLJjA6VzNiaZ8NbROyJcR729iN/0Qz9myAbxX04qbhtu6RiD3/pFtdFdg
REglCwdZcRTyJbc5aa7WUnzUu4pTtJ4OzB/XFepSc4XqYWw9lInZLERr5nwD+gyQ
luCBmFDvDAaC4Vx8nufNcrfHyd584WFYtCaB7ePN4XZVuCwJSS8rjo6MWLO6ZTzo
O+UnUouEhXVg8PwQBZ+GP1da9oc443Hriwg9r3gtNvlAWOV17tkGu/KtKZq5RMm8
LqXHRkee5PDDwQ3FZXluc47Q4W3W+PlWw869faF8WOOoX/PUbDjxhrvFAT6X99Cy
NLeh7zHd7wdpbn6YfChlpTgPHX3URbyiY/ML404KLJClHM8DCRRbbHHaBUJhp0Vf
rmqs/yH3lcUcJSbTOfGpKOKpgR8WZept7ze6zsaaATQ+ZgK+O+mEYeChHiCg8Q7M
PUt3T6Q9vAzhBx3W0UoVSw3x0WJFVhb6MGt7YC8NjZAUCekKByDE5xUfgYF59fXp
1GLpKAEqzlogRtyh1gBEcWJAaMVVXhfc+ROWF7XvTQgEV5xbZ23zSdY8JGwp98cG
0NwNHzZLmRCRwFrWeaceNyFa15yTIZvM3qReg8GxzI5tLupvD/O1Wnwvxxsd1u00
qEed4bPG+RPdqet7FMKJrrPoA3vmuvek/1wTVvngee5GFQ8sFv+DOkjWwtjIRz5n
+4y3VPnt1zzw44o4SkBrfywqIloAuXBnnJN84h0TZoW+byqd4cU6HtnyFo5brYQk
VP4mOlFxokGsA1uYE1jgvBHCzpG9HCLZi+8IlVDKbUXeZqgnBedIb9ShsT0DD/jG
isUMUwYQ7tafdwEet/cEEBnpHHA1YAvuD0sW5U7vEBUfUs0K7k42Tqmv2tcyVeHp
Xjl9NCMuh9tsX+Xg4gvixWRFAJqhiKdt9lcK5pgY80XJGdAnBKBI+yE1vfYinvnm
55TzF33e8x99S3WcFrSkuj/5I2osAswnu5b+eu3A6PaoRPNI+MZZ4kKP70qRV9KH
6WgNiTuDjCWF0gmpyMVhVIF4Qid6pRrONjGxRhRmb0keaxo7+pFcuN93xOy3W1QK
k77zDu/O4rA9QSAVi9Yz9M15oSmglyZLBP58zuR59W/kseqWduFKxmuccHAERis+
manxOPEUBsESM1V0RWhj+ArQP5MzM+hnXDq9qUwUuCLTywgE/D6A5oqVbcBXCE2m
TT9+bbZtUss/EVWIYDnm60cayKnItxinZA7Cp3lBPhAKCeaOCRmEZguORHkNknVK
46XBopd1EPFVO2ndDJZwCg77RItg4cEE5ITUFFkjEb3BHV04rqgcVfzFdzkSWiyl
MIS90aiA7T4h1ZT216RHtq/UVryFS1IIF1ZQVcaxIiRIK9MhqyvR2FE1wyITFnjZ
VHkKAzO3c6D/usci8NJKme4+vnsHXUY8bY25EIKVyhN9Tmoe6KZehFLXlbctccbp
RN2cNmvGXGJ63AX1Qf9UWaQoyaJiEEuTBATCGYXh6lTSI0ADy1fHWLOY0QxOmT6K
djPK6kfPE5gzwUcJXfg/0RthpdRK7em0Xok2AeI3S2g+VPvTMteZYQVbuUNAFYyG
lphGSZTRmrjMnxbmjJlvf0Hxfnxv5eLWfMpKEzU/s0G1A65v8FOz19ti9UuQgmOu
UfZJD0lB6p7ywHM3kkcsVv3TFtIfgh/QM6yGLgSBfMWORHLzvbs/VmH7xFUxKSIN
AO8KbVrAp3uJeNtECqs8Hc++E7RMIv67cuzC0qt/2OBBnw30SaRJRDBAvBB+L9No
t7L++M9olA0oXI0yGBWjJC1hnv2O5Xwp3BTKEIOtpgC49i0FxuRgvqmfwz8I8mfd
7MCVc3r7sLVtusV7kWOb1N5etVYprT3712L80+M77EenYxbNlWgmQPcCY3j2+qtp
SZveDZqfqn9gudwKPyDwIF4s7sXj++mEY2TCl5mjzbgBfZs08jzar2L1gTf2zNMF
fAe4yO/gBeFKv7sVvEZxsgpjH6lc0DVRi9bClFA+5GtXVrHtSoY/3fTJs2eoHw5R
YPRs+LKeaScD7wSV8fZa1Z5lU4m4f3P5vP+vWVGLblghrfVkEQGa5XvJDxDidRNy
dbgJ8fu1+P5L31aC3omkc1dBE+Cg/OkMPhOPQ9lEdU+DKM5nf+NrsQ/3E3g+KdpB
SpiTIjxxTM7V4cOhC94GiMc4m76AG1+6Sy5syIyXGScTqgAsjV02QClqgoI+Dsut
9hhqqAGG9eeEqrjLX+QAOYRymqXMPQljsMM0rMHbToFJvVruepDwBmnNHEwl0Agu
eqUrAioBJiO9468Rvo5TkEgCMC0Btqj7Aadk/kLTVJHuPmk5LqXxMOEpzGtpjY0h
qnEnIX7plldbDAAWeipuc6nvWJqBgAUfQFTdhXQYtBf8OEsqhvDhfVaDVt7dly2t
TO0Xzhn+kh/4X3VlQx6f8dGmOeQlGduXmw9DbIiQcm77fTUhhY+/tDkkaS4Cuyhz
MFasFwlgIuq+nb07fubUGv20gWkspaX7ZQIIFzG0zn/7wx0R8NNj+wNY2Y2rQXcx
U2kUVUaWAuSQRa3uhE7PnX6jtwzJtlWrBgXKBKtoHYULhI3cjyKYdgnfc2Jv70Jo
eTCkrie548orGcGd5BPt2HB7fT04vElh2LtQ19Iv7q3tcUljAkslxW7kXVXEBWrD
0lM5FOxOS3AqgURZPPbrugpYX10SiYRayvLnbtbM4eL7gK/UXGqitCCbK5ysHaZb
9345p4K3pvgqObvZvv/Lsg33ZWwsreKn2nbeu3fflYM7wa0bBsQzsiSPBsLSXX+N
l/gnXHNDWa1WN89+Q271WKkqSxy5Ljat/3kH6fYJ37AE7SFkkHYllBEdIMpgavy5
EOjOWS2cODk9hIN9ax22PiioggChNRL1E9Wk4KS20/iHuAR4hjByL9Zw9pIn8p89
bF6jb5qBB0fiaNL4spNQva/TI+lm378AOkj9+zY+jgyjmkF7A5zAttWa2hAleut0
7ZXHaaqKxCd5hKWEEOozKA5kEIoxNSRxSYI4At0G5qQC3qttlae7NK4+HnhsGmNI
+XmwWVZ3PYh6g6MN/obnPaBpL9cn5r0y5uW+Q3eyT1KvzCp2Ng5RjIlCfNlqxRau
1qEKCh/Nk/opguvoKNRG+lKuDoVbNbUSDjAT1L1QSQlaDBhpQPfL0hyMyN1ALvPK
fd9pS8G8Qd6uk0/QiBIofGM5gFAdHVA6l1sIvtMavE2nB/GCtzriLHcrG3xYZ7Z8
tDjGeZljoGD0QxsSqDjM6WUSSOgYU7klysOcMLBt+ZkanT/Ge3l9PGcmCw78zzVU
LLX9qB0sdtuq6eVpWBF6NQ+Iw7esNk/6QvuuIaMZYt2xfAFb9EjDGLjWaRay04qC
zqS7MqxUXIFxQzPcDaTymhiGwjsX6Mw2ORwSgyLQHqjJ+IcIJ+qf/FbeIjItm6Lp
V4v24MUSkMe3Q7U4oQ7GirqPKR75pQaWVOjIIaiG5WNidvVnpe7dYCQIYPf1kFNk
F+UaKdMdqhmUwAIO/8q82Jx7h7+OU17owpG4O+LhniUYXaTdUSOTOgY5Y8idKk/E
ucuWHcqgK3S5oER4HSVQRxe17fjgXnQYjq+AfGoOW8O0z9n4RIu5v5xZ/yuITflw
z+fFExpdbtP3H9ohfN2JLhyJytx0tEcH0Zo1s9qIXqv7KNcyaQLHLNghjopMJX1c
haEFslWeND/Pgh1YtirDsSXPQAr7H61eG9k8wAFI2+PW9PzryRX3fsZolK9CkF4C
tiMNCC8LOvgsva7CsckIVBl+eqY4dMeIlXXtLR2QCt6MR7pX3enuPIYaA6oKegex
0hqYGUVO6KC0KVT3LjFkH2OHV1++IWFN7r127Wk5xrMVfqtcMULFwXjotcluuCrr
QaXs3C+YcLCZ2ZKZmQz/tG8/k4WTpzizSNf5IvoiMePHr7Bls+tXnF5NUGB0qCFc
GnkdPZhHITClQGsDOHO4Djfx211XQDtLb9QyWJ3y8fzvMRIDiFf+EltzByWczJ+f
J2nikrVpyYv23zwLmz6ChhZgUezt41rnp2FRUQBxv6JYPyEZPREh0Al29GIBZFCu
DzJ9cKQdSPGFuOioQgATu6oduJsl4vTY8t/D9y+FiOf+R3UC26b2wIf0lh0fANIj
rx0zNv3glweTowDIxhrYs0NugkP2ILGXCRXlYcZpW7yp/lIMDjKaYho6s9xRKIYz
a4Y8hoHXjsH+JBxwIEx1gZ1efG6odrXbm4w6DSUqE3GI+vwabIxttpJUSryZs1um
/jdP8eT91w+8810Fva3KOH1FifgLSnSucuwyp96QmNtXQZPi7Ze26PwSdAPmYxn9
qKlhCVVY72FvznWFIOpH0v278YNTCrCbGLb1qk3ctXRGbIBzy8p1e+a76i45kqry
q43BHjeZX2zlSF+BS41j63TIE9eH+tyCSqaAw7NIZoMZmJvC0P1lxFq2jW5CsypC
x8N1Kcqp9DF6val0n8fESrZ3HoRa2Ei6KIaPGN063O6F9/rDFMEH7275yQbzTmTr
D+T3ms0AHxqaW7BCEZGa5JjCe79dpOAWJ3CkgsYE9TNWDA86llKn3eKC5cKF0GxC
mybInKWGbeIh3yZvo6hDbI5GqIUPYIsgH4M+gcOfE22gk4GdSu3ym2rgvjoGSfxC
t8QYkYkIKb93pifMcJqWBEwT3OqPQo8RUwLKhN7EiuqbQCsUATni5Fk8qGcTCgQt
15zHvpD9rCy3aR7zqT0UEIBtOJ+yN2fUWTvUn7aJBohINtjGbk2k4fXqrvwpsQik
Zc2kQ0FdovqQvqda/BR7bj2vVGNXisB9LfJquIcq24dmta/jF9TgZFGhDIxpR1tf
1utyNiqh5AsAjhWq1qRglJtz/YeG8SLLbMxfu9cMAjSh86kBH03aeguWhe+f7New
mpJbbCHjkTHVdwQlroadXYBv2G6t4NAmXnlgWOp3J3hNrXzkmotrOf4IuSjZ9biz
BW+QQ9aDwdhqI+s5pWFPOFpoZ+pDy93RyPP4rVrWRBFcL6Yh4D9CdhWl8DoFfaDP
kO6zxzbciUWjo/J2/97PZRLKEeS3bT8iqZQpPU3K7VYVplRTTCwNfpHZoSfhJAfE
99QvXiMl9ZYEIEJBW82ALtnY/pYdl0XQebnkMTG/lpBDu7z7kbyLpitHAMM0/6eP
oBc+olqU4//O5Bw472W0vwxoOwVs1nMakA+yUB4vUZK6zzBYSWAjfrKngDD6k2qZ
FSmuDKOs+quUwAgNbNc8oaFXzwE2aPgEDR1pL4wipfQbAF+lO05CiWW0dY5mWbBJ
FZl+l5LGKNT5MjbWq4tzLLIQK5QQ4eHOHEMFMFHg0BtA65lADb8x6pEOtO6Wfrvp
pms4+x2QpxiLhVkeidKEFoslnQxu7GouH5v9ulqqtqPSU4JJx8ooac24CbKf7a2q
q3pNXAPIqAxAWibDuzEctnEsCPbZRipmWWHS0vAh20zAuztofiL8MTtbYfCf/6jq
8BbSaFLVvZeEletHQExGZ94avo2AfW8MwQMUBDkruP88XeKmdByhllXudxkJzwkm
h/+qjjs6sDK1aTdz2iR/foDVc+s7g8YUPEfX4G5DRftYbo/P5vlLoi4nx6ME2W+6
0kdaMGCvdfodX7aBNKpMXs5gOuuqBXmAO5qzImkcpnopqChPtnbckCv+fD6cb0+Q
hVY2Rjg2j2vJV+qhR4oLicE+2+VdvUUPfBPivQ1l5Gu73Jv6G5QX/QxYDZ0OGe/s
w78hZRwWV5kcrmqGhJ0lcn2C0OprKx5IrpDee/DdKBatppXtc4tLzyk6Na9oLQvG
SK+i6Hr/fgHiiFxMPi+AFvCNX9XjDnB76ualnZYs9pEeuHGKmkgcmPALyzIj0Yi7
k+olMcJ1y6ywOnTGNzImzyvgs0IAd6PQvxEomSgLH7CND3oCCH3vrgB8plO+kAUp
whZiT2GzO3onE2zAoffVfo9WUGsT+MnDByD3oYgwxlUY4Rj2XCmt3Mwa0wql3u2P
Om394LC7o9HSiXvtL5o69ervlxFM6m9wnqZKLqxW/IDukDLJxEqM26V31ccb3gOh
jcvPwZh3269t5rzcpHiV3I/lZIy3WQ87/cdbZEdjyefqDay5V8SSeY7h5Aj6mfnX
4CBZRKhMU0eZ8S2KwLD77aYnTNERHT1bWYGgUdlX0RxOWkYd+uAguJo2F7mB2FyQ
OcES2dvcK7vVwriBOCS3XHeMIDvoA16YFvkDPlIwzPIGqv9JT+1n9HNms2k1rpkN
u5jzze30FxM7zV1YxhtiGCLUV2eKUSbnuPu3LyoF+30kGIF+cRRPmDONojgsbWwD
0NFEVIaS6+GmH4Z02w6RcVevrtDX7HExpstkzUHe+eteKE57FaRwd6yvhtNK4hX2
PzKxVRB6+oJVxqz3kspryV1UrFyRjza8K2XMRfD2+0V6AoAFkJetkoEhrIToTAL2
/LXEUKaYmcw0c1AdWG3SGmv7ncsrnCVBB/diCZQlS+okakR2IbOT5iNkBMbh0rsL
GlE+5s+2N19xLfprWP9K4AKWldDuE0qkdduxvpFITB7SLUNIRSi+jEIeaPVy/QU1
MHg6kK4ps7TZAppIZKuHP8h4gYbmSqBwypehq7H/Di5fr3nPfgCj6R6yoUfCN5gh
EhjF+WgDbLnLJI9p2J4mnFc3MWABQM5SR6QY8XuMhTTNCCFyFAxcL+MJPcfRIyXc
PCaNDsSHhosSIg/kgs1T6LfELHrpaD00HBrH5UdOwoqcEx1PX3hzNIWW0AHlpkTz
K5wm6xVmrcMXoRWeo4Na8Q/TL2HX7c+N/3FzhpBhQfG2YLUzlTIXH8wpYJljHnRR
3u2GTGgOwTNeA2PYsGIWx30XpNStOF/g46qh/o5GQnmWhoSgKDPDXi3cZ31Kx6ag
c/WrXQQv/9gbEb7hlApa62P8R5eoHAp0DmAAMGDMZd7etjQCxk1t4V6OLxWYXWjk
r/OtZEZ79wotbTpqCO5k2dQVGTFZkA+/wH9vLDddVKIahgHaCRS8YV8TOArrqnje
tcdLneFkv5szrVr6UFWd/lnaf9M3EU6tf+6KvPVhQGTmKb4GgPh4jk3ZbfAb3L1v
sm8pZwix41ByVw2caqt5xcf6ehc8Ez6OApj8RQnFSG+csVDVQbPG+64q6hMUuZzv
9CgR0qmdyXS0dHTmvCi91Uh2dSz69uviR0xP4zjOkAoq7jKv2AqRGZHNLRolt93V
sqH38ZrpbqjxuibQSZSHFfJWHVruBqvjmZCwySEXz+BLtsqpx8dGWvblBmo8nwKk
x6M3MJtbwdiaCnmN54xj+9k91noAlOl9jhXsVgWnzY9kH6apWWc3/6Kb8KSKCKnR
ujG7b/GtbORnwF8aRQwcqsjbITb6qnnGirNwmyjjTRGDJxWbT+3wKJAHcmzmLk4K
A5dUeyj7wAVCh0dtY96h5XUnvkkDPZ8+aNSqXRByfOpCeLVrTsmpSgM7qn16F9sI
8VPi0VcBSnoCrTNwpioB6xmneeV27RfI8xskLOePQAphXtSe7JBBZ9LlyoM89qml
hzBhF497IRtpDZCEqCoH7tNVIOvjXWzY7zV0Wk+wb8eY8E6kK8J7Khco4ndtf8Tc
xKiSfgSL5d74InmlFYNoDsH+W/CftCwUxYnxBaAeCeynhiYpbzXZx+BM396bu563
sUVzvIVV+pasgAMpOMbI+j/2WmVf6s88XEizZD9QpLyLH0iNvY6KGT/OkCWFLvuR
3tAlCWGKsmE0GebthCZKgTrNQ/0hshQBzAWAeZN6qo3EO0ZBkF5YXaKIr3zeo4NS
3CWPK/S0CeOFIDQazTeAp3EQuLWW+An0g9FYvcb0eu3jmyk2UQi9wX9MuPJUEII7
vhHUxyXv2Z2d+ruGwbq9Rx2FU6ms6ubSp/EZaoEb//EzsLFjomIbYre3rcuixzWZ
AJWq0JKrNGOyiHWCGqt/KEIpMyL90nf0IudgqvoJSzhbW1K5V+73SvJobZ6ZItAo
MAq5egAW4VTqT/qS0s2U9zEKJLO2l3kRKoy9ZpzrzO3hTnnKIfGgx+SKqjlV6hyP
A8JfAAFFss6akSqVYuQ62M7qiBB6xSykgw14pdQxQNialp5XrPLpJxVGzdFNmNva
waS69fDIZxhQEJpFzFgQpaOH4H7lyumueacr9igzmzKFiXVaXla3+YGY1f6X+zKa
A/52La3+yeuwH89HmlTeUCi7zjV5nWqPeYk20AJbO0tP2TXAAmp4SOfuS/gi6BZ1
aoGLzd6bu2RhpU1J98FBcwLQsEdVE8Bm8j7SrEyDtQNf7BDCuzqxDlSv/zDG8AIR
dnOvIutdAUfSHlUHxTKWFJBRn30DWQIKCY6ViNxschP+41TQW9Bnz+l8vwrp1Cny
ERMaZ9Nm5TmwNVE/Bw40meRM8jZ51Zk9z2ev6pYh93Y8K5/yEQ0d5n8JzUG/ac/P
SekyqXEUZUrshrW4LbzAEPoJgUA+7+7WngAScCfiwTQzyHk5LrH87fn2X9USRTaG
C4j9q+4ioeCafySI4dTGi6AdRprtt1HWPzAPSvyAqcYNAfKNZcTWwDzYCFZFTAa6
OoyR8mXNA2QlAHPYMv9/vuMAtCg41PVOmyOZ3GgTlYroccHeZu0HRrJ5YkZxu4wy
H0UjRWFvAmjMb8hJsFkddQRu9ti2dzgVgE0CBiGeR4nGBWPl8y2k4MHeLatZstd7
F3ROPFBakQhAh0DJiQv7jGvhZqbsWVSNPNGl2UcenpV367EMZdkYepvTVEGX/dGX
C2B01vbZE7pqcxL4w5sOdxYxdno6LiiYrVwp3/a1gQGoOtjlhsQ/G0mhnBP4gae4
T9p8zgnf9MQqXrq5GIa1LD9bMIU/FlXsDEOnwxA9eYlFnWt3SPR/dM/tDzWTyMzV
2Kqj0BBZulSE15b1sqFz0a3MN9KsNC7WZqlVZJJfgGccSgwfpzJ8VfDbcJeM9WIX
1AdJyV7FOzJY3FEbKiwMfs1rW9qKko7r1CFtGnMGt8FiyyG6By40f1uM91pXSF0L
50UEOlte+qNQq8RrxqqNb55EmigpbCDW4QhX01Y4TycEjMMtZJ7J7jHJB0kQBFTR
WAVSK8pzcIsre7YGy8d6QbP81UAJGo9xyXnDOj5l1kPZ3fQv6B3qXxpr0LQo9/42
V/46yVrmgOnfHlgfKdfKQCQPrM4hqLHxQkvymUAibQXOCdR9u9f2zoTJqo0sorgn
kjspDqw925iFTUzVfG6Z6SUrIxnS+2YzG9rUyZ8owIBmuCEe3Ov/6fp/iSOYDRPE
TLu2JNguXchhHw+iKeTEPt1bs9YM4BAM81p1xqCsQa2u0zvq1kmoh16AK2RcXSai
KvwkB1NQ0tTpNKzMMc3p+GJpiULf82GZGAWgNaxmowkZomHA1JU+J3zj3NwtJOoZ
3+Y1PZAeo+fOT75hevLL5icm7eb24/dmr/q7rruFD6vXU7q/p3ccaO2NxiM3mcGf
vXp/ZF6Nr4WULEqYRpKM7QJ1O7aMEqwk6FIPji9H4LxN5nt3RqvJYMTJ/ZVW5XRC
CTnw6O508GKYI4qTUDixr1LUoQMCE04QC6o7LaxRpjPSMwHce9MDDv5KYd26C44C
UCtnRR8lhKgVBTtzTUgghgaeb27lRkj0THJdOXk3dF9yQ6x2vzX5ugZfYIqB1MtD
bzPlTMY8OrCzj4XMLCxh1j32mkNQe5afa8z8LTpJSkbXzdKWUOHAdhvgnmrg1XlP
j2nPa0xks59KY4ywxy0PQ7eCGbtKdBzmgEuw539DPEfbojmxyR2cQQxFVZCUMMfr
UUT6vt2URbyP9hT+n8JcGxDm6UkyZeMmoPN9QVMt9dr68Hu/RrN3S1VxXNf4Yx1Z
AkuL7gxARimBapKm7yoMwByuF5Y8ZDue4oXGxwroWs/fF1zD0Wy7hhqoUrpGvGR7
P1ssO84j3SilrnnthxL0wDe0hx5KUcd/w82ue4P1SILaoPRvvDyiThG0+hCJPKL5
6pBM2U8MY8jIP0fqzVp4b8YPRNY5JIVSmFPvZ3dldPon2xock5hB/Gz3CTW/HgHc
qp7W1IzhyEzjFsy3MYBJm/hgnQPFZrYbi814gs3qSQZeY1krqRFeH+WyTIC95Ij3
PT9/cWTEZ+OwtTJMa/oIhSSAHDk2xh9MjNk9eMS9ghmKgvSGYTdSCjaJylH9WMQg
OK5ZgdNvvzVKXNXUKVLWQy4TQnOxftx1XIVdMrjZHIskcKKUyOBkeBSaw9l8isK5
oeKxwJRCMQGB6UIoloVIO0FDOhlySMxcf/STH8TM1Di1FwxakVu3aIUMNY6MS1SI
TbNboq84dkTc5Jjfd9vFjiASJHYmJQGsQe4Ua6uHD2IRK69pfYL7lz/a44raZ8V6
OujzQxUNFLCALLatztH50Ngx6vPsM7AiDLLOd/wKtWl0T7Im2lg4r/0wbISqNZF2
XyBizwHexTdGJ2m5xAZuHWDG0ulbIHXQubO17rx0KzcXsSYojow5EUwAeNFDP7IX
wVLh67dmqNof/u2nQu4InK7OMhbp55E9VwAJzfUKsKcvW7NwttkNMUAHd+GevnKw
PjgP3Ukd3ag10wmaIRQBHS1qs+Cqif1fWQ8/FoJ5IJRuhfh2YhbxJbwQdy9cN9xv
4TMukyGyHdLRzK2xEhmviC4qmbmMFS78eKssKsTO6SrTHpWe3eCp0Jyb85hE9Ev1
88Bi0R9j5U2cICUXvXIX/o5k7Q47nbp/pGWoIP8uuLfDm9KL88OQWkgn3DjtoIeR
krEKZgrDAr/MMcrgM4b4wL7B9f0kjkaBqo3AY+4jvpkY3cTh3vh0Rxl9ouF28IFS
RxEDRmzTvR/yI9wqLG6EOBDPjRf+blPsMzt5Rkf07UXXOUQdop/Bg9SKgdSd8I+r
a5y2vO1l6R+YI4yo3JdaZieCNeJG3re87alR8s4ILooIQBVYnGfZHYZuUDJJfXTx
544w2FxlFGBn63Vi/hGA91pIkYFbFFGsL2ukC5mn78zdOUhBOCV25L+Gnx5oymj9
9aO/ZLaZhiASc4fg5Z7wEiuQrJcMjtICY+D30jG1qCCCMGNYj8YdVxSDJAgYd3f2
`protect end_protected