`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 57664 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
5lZBo+Mj1WIDsQgTk30FSJt6E55yB2gwizbmh5bCIBVQzLmb5XY1OD2qSfBB2+Dd
/xfMwW4BtNGl1UquzFXHE0BcPzvCO2xkQufl5t/y0YxXtqA0B7VwfcZ0xH9vVTXD
8xy/CcbUazL9gqhytcksIzfibeILRl3cguQaFTlXdB/Da4YGWgvIoyqqeTHXVn4G
o9PIrzW79ILJrLQabgolaCM/v8Qxldq/Kp+yBkAExHupM/hv9vVVB9pKOhaRIq0n
ACgnQvZ+2DjRxK8XmYG0V11EprZzjkBZdx2fPdJX6Aetqwqzj3Qq4eSCJ7IfCuLw
uDc7iu5QjPKeG+/CAaDXKysGjAwmXf6B8r2KhhbVfuaa1IkyU5Gp8vWhMjmxHwq9
SENpfmsni7LmS+XD3emiZmvDtknqyHAeKA8Y7DpdtOljhHfq5sy2YzndtaWen1h+
KG43nDH2V1/dSw8x7yX2KkPq841O1ApVBytCmBBIoJQudEIOsWWl9jJa/A7F+vLA
YeHx0nOfy0e12eGiX2GPvL0rK/Li80j1OFKubWA9sTJ955H+q62wS4QTKrq4KOij
cbvaHFwT09TBdmHFkiqJzsB9iuCoT7d2+Lmc+UUBg8dFlhB+dSu6beIUc2nBVnR9
F79khk81VTgloahw9ynhtTWocdqcjJ2+JaQBPx4Tr+lxCNmdckavRv90VN3Qp44o
VpL68KBGqW/5WFr18jpbWuJ1R0NcctvcDUVLA3ZincDZL4ISe+C/pi5XQiDp+Awo
T8SlrZqZrFYgH1Z4ajA0H7zs1dIfGXI6jyvEldIYiqnoeLWGuPOfl/4eQWvCIW0q
6cn/unOZm0rDc/aX4yGyR/FyquNitw0MYcuSFLj5aJ1QrB/xZS8SWA5arNI8nfs3
pxwept/8BzrOHWsD+JLzGk12ZQsteglJoS04+9wiuBVGCCRK8Ghb5V3FP0IxiFHx
z8hkTd+QCZ+ZjWZoOzNlSlM28E89M3F3Zka1gXbMrdm8Pyzz5sE4iHowmYROZfnf
lG6JyIcve4Pnnp3fmVzQ9+XfkJtfAst11lzkLmO2f5G6Y5Bs8RznVgx4ZSC3MLbW
C2GvM0kwmBaUoYVQx/B/IgQLbqdRCqBES1+/14TsWF9pM2nf2fqmxZgHz0sDRKow
cTYXCU0Up2V/kpQBEI9R+l2+2UOjw0EB1VM8EGo1jWqqiXjifPJ4YBHIiBYL6GJK
qC9JEdCkkt7LSu0OXo8Jzbb8YDfv7h5YiYtqyddDLUBuJ3l9MoL72YpB/Fs/Y7bl
iYTCiLbh8DbOvml9dZD9io1qrUxURh23tT+oAdh+TmrQn6C6PHCfT0N6tBNWm5A6
VCFi2EdfUzS7OwXG0AgwJznLIcAoHKyiWCEiutmJArtN6PtfOwhWQXPOP/AeaNov
QfJAB3BcZE7wRkUKTrnZGhBzshe8S9qNB7DfP25eGWwHhGABcKhS6ioqd1dr9zsT
0pDlCVyF3FnHH8kjATiivYZ5LJnaOWYP/GxmYMC4APG218L8IjWaNxwFv2sQUpjW
uNppwtr176Oorkh72E9I0Q4/RvPQeP7wiYgPW2CpSaO7TqtBUN+0penMdHLeyCAC
rJW6DCXD+sNNZ9YEwWKu+AQu710cgC2+T/l7j7r9vjGWSfry6G6/VlwO/pannC9i
3sQchPaxes2hjWm0Az6Hyq3CrLDyRvIZJTPsOUohcbdKaWENChG5dYd2nmZS6eoU
f5OtLXsjnWmsfyhzZ6cjmyP6bgVWO7ia8ZGyp02/LohBwF4Ql65mPZgUtFlIsrII
NBQzUmH0hqOPY67wdqq7y4acs48jMJ4NuMCBzKOzpPu9SUV4JmY2kovFJAHjPfVF
hTCbp9iLU5n+MHKV32Z4s5bzqFmy///BOHO+AG9QuU6fZpQwfNR3H4uJL2QKjnUz
8wXV9u61NqOwwDw4PV4GknLvjOLGBp3KZJS0d9nKKKh2WaEdD9K4YcpUCBDVI+RJ
0GV2Hb9wuXOH3HxKm5D7vhWGWJgmMo0vpzHzOST+T2Pk/4ABQDu8TRjv106DiGiB
M1R6WkTkc0+ftjy38F8Xra51K0PEHrCxtUvGywt4N8Hli0jqNNuRJeVLJLEOpr5I
kgo5l97kn8TO+NUq2y3PTPIdjjmzKSWVwgM5jXVhzZafTt+TgPV8JuOjhJoNY71u
94s2KLh04lHYb81hxyO5PS0kW2RQADeZoF5IiYahBZrS+1Pgm/cYi8pfuZvJdqvm
LpJzqbtYikUBMj9dQ7fh7eCgbT7U2JprTZQFbl3XqJTmUaNnMxHF+Z2K7ANeK+YN
Z4HqdnUmOpBsG4AW3vUiD6fm328H3AxTce7Prlboq0yLJvdcUe5HkFN1q4JLvOzx
KpmEuANUJOS3hMQGhu/QpEiwzHoNKaWBvwBV5bPqudRmjsY2yxgezas9TDscq5eB
swt8gNVO9qdI4wqImTEbrbBwjKmenXs5WyNI7sJ9e9jty5dYR2PBTDpHwfGnbiqg
K2tODV9Ri9VzrDgQs1T3kHNcxn+i8NjN7iaIF0ck2yKAnUXWuYd6fgAHIDj+FiVI
NL/DUiDpcXJ0CjeeKpciwvdwlVbiaG49UaQJdIefJb5GYrYHGAROgIIBZAjuNHSk
g+2GP6QPCnngCMUL+k+Z2v8AkZ0sIXdiT7bwbeZFf4YmESgsjwLFQPlGOy5aIiPg
2DnHG5h409am9JJEEqV8Hx5PYq49m9IlLie/5wfWQHZH6Lyuj2UP8f6/FUA5hFNQ
iJvqxkBsqxkkfyGguqjXcmunJ8UvVDCee2gcnbMY7FxZet25QyER4uz8H3xQv7C5
dch2ASq7FAtyM0omr9DDqJDj8cQ2Y+zbczaA42hcNr2RKbrXmNZJFaeZIXjHpmYB
bYWEs9gdZDutWqk4JQ3Fu+BJkSwY61nYq5110DzXZGUO7a3+TfuS5zdk5RZP/eRn
6JgCTTHJE+GZbbWCqig1vVLOTiJbftkPKZs78EjOW5OjjLsloUvAgn0kgwqdy+3F
12aQ31OTWo81svpu8M7FeNg75sFrpFt2byDVK1X8Qt0byeE5iZIJ3GEsqTWHdxNh
g6JdAfeWMNDLTIHjTSeHjLSlpwJF0Pw9OwVe0PF7PKh9QUHA/x+vUg1QGCPu6BGS
8bsB1KL1+FHTgtwy/l2Lh94LTy0IsGklxDBJusOFF1rDUXUVdcUQ6tVelL309uAC
LD/mt3cgYzK8DWz9xWnR31t+Yi4z5n1bzOFrwWDRa5+LnYPwU5eF+9CXuacu+F32
vFZrbTsTiSY5hwBHxUVVTicbECII2qC3vz57oIrT/K0CXx9FIhmOxBt57nUMlvnh
lCq7nPip/eu1FxrFycqNPNdxS/BmqzaIp9FD9YSOWcXbS70u21AcmvFjE9MEmDSG
age70y6etZOCQ16wJH6tWaSs98DknGFlg0zhb4w5UHQM2fKfmlBtuE7XuJLNLuth
9CskdiWkXSN+FpGFbOBdemN086LhzQ7Ah3I+UgG8gPLcGV9e4taUuI4sDGmL1D3E
M4Dg/yxGp19HjCjy2FQnuBkriDzQycN7ynBAdi2dSyCLX6KemBh1CVZcav+UF/PC
WpDVM+cr+3xtLjCoA258KZF6/T9TZAHZdAmUz90OnRscRNE+nwGE5pVJhL4yU/WE
Vbs/Z9/TbB/DX9cowzAb21TlBhEDTIZy2vxsQYR5k7/RsVgJ9KrF7D1wSCvnoJGh
LTsnM4Y1taBhj4K9Yuex1/zmIM4+kRhon8CiyVJXfsYOSny/V397P/oPWHEAYefu
FR6YHZrpD3aSgSeyWy4bRLnhyiiNCn/hK7qSFPSbPnqCL8w8yIxEbTyIMnb4Vxy4
+oPN+8c74BasCWWq4FQxxxiegjzrZZ6QHN0NklbtsIn/3A8Zig8mZ+f8mJH72qX/
uokFx6vqM08kw1nT19/TQvBWQ/rCbFGA1j2TA9vOJ4zbpgvX1W7JlHq6pPiMjOMN
7P75614gM1b3BOkOH4o6OVGhckBjjNJ9MeKZH3slmMoxvLrkaBu7VaRvdD2PNMDj
68+5/z2xDXn9hpQbnZuagrYrq1KYhZgsMLverbQwogIp+CuKzxAuXe2WyOhFTxOq
ReavJP2SJ6DQRYjn0ZmLZNawPk+K0USFv0ltbEu9Pr0rNdx3Xjmd0Z1wtvUdpjfS
jQqGv1j1e7U51c3UofB5JgJLwe1Cwkb9JyJ+wWAYWH0GT8CJQ7iWzRIiniS3VPZb
33ruPGG6XO+TAcpDkXdypXP1GmzzeaEETPKBC2sSOzsbpCqXmUD6t3t6k26S7FQA
47dSagdy1e/jFD6OB1XeBo/iI4V7Yzkp3x5+Aw4Gb9qmJgzUIpkqBsY8wNN09PGP
tjdpkar0TNxxqOUeXHgUCMEIRKGWnn1UVpH3WLT0cN6eC+8JMXPsbtrWwpAxNj5w
4rd9Fd5kRw16NvZAFpLiTgK1rcdE8BpVFQhk5TDIxvMb590CTa/NqZ0I/s5clgqU
6KpABVkuiuaoyRORo4YuZWpf/+T3GBIMOi4jzAdDsAbf+qgKLIRX3HtSZGiit38Q
UwarXmMarhlxe+iLqs6P23cZmDDqtkh6w6pS4eFp+Aljr1wWxw6KVsKHpcfrPUSx
1PkZ9H6sIpq474/Sd3GAeW3ysjEbbuO1bW3MYnDTAE9dFDLMEaI80KCPHIvYYtbD
koUjt12deezo0F6Elhvk94ZLPqwNzQDyr1Y16E/wNYs6WZg1Xdp9PJlNDMc0N9uK
RKSMLYphqll4BG5m1vGUDgxDc/Rs5c3eVKkWlGrESlur51TJBWYH+vXKIy2z1IUK
+PdX/yVSS/Ctz8RAhFNqOU3y10eogLzakseQeZ4jiRDB5dh1mZFPgY7juqtyoySU
Rk8+91FcPoxwZhm8GGLcGChsSnOXvplCYXp1l6qQiWSma2D6FRNFabl7Ayb1uiAq
ZxHR6+LhTLImDOwVp2bPwuutm5caDlsdhCKBTO1MYHxOeschlo9WCSGWUe3fd0b9
PGEcZcV8HmXYCiv4L2FHJBwcBXly46kEt90ae27xcNu4721ZBUPQu54/0AdNDNEF
P+hbrp0/9PX1zCqmCQhfyDTsLM9AWt/53JhJwv9etxx0aXE10i09CckliHOgPw7b
WNlFB2XhX/zNAgBAB1OKzYdd1Qx4u5uOBZkXs1kW/D0ZQJ5DVJ+9LMisN/K6ELAa
I6LMelNTR4bNS37VMCZ5b9b7NpWQmpngsBya4ev6f0hg/u021WMhY7J8A1sliLpR
ypryirfpl2qrELanwqDo+4RTXGyufP3TRcbW0i3hXeNqhpljnvHTVFoLaWDguWiD
ZyxGrcCaSJMx7t0kLJRlWevQjZbIMTgs0vbNFpnpXNTKcJFCQ2sgeUT6caYRa+10
I8B43D4qwneRDBFS5AGcuowwA7vN7jITJHjWOXq0sfnH1iAV+o1T57ggLSBEkQiR
5K+JBYdEQShe+c5egdsJW/kyGPuhl1N1jYwmu7hcxZEn7SuDs2vzi/jA9uLHG9f4
in0Fp0w2/jzffTpKBwzGlF01FymAVlxJwMUMUvuyxpRFr1Fs7U5UpwyhPQ/+ej8s
Rfn/3aEFrmFjCmlFBp29laOl6jTniex+r1KXwGTdFCtutt+EcweqNh+7ExHT7B5W
EXqjnm8FcrbKHJkSx8vNC8VRBkKr2PvP1BG7OkCTgG5Ck3IE2Pc9PdNgW6/ubZ5U
1SCz3OV8gkxOFS3PFQaFEklj9GIWV0JTq5Z7HyuGtSgRln9nr5DMOEPL8hAVic7m
+niMx7VzVY6ZsMxB7vbTb+ea52t7gJYvgA3L3MDk6zgOaNLT5eN/6rFCJI+lW/cp
rjkmGN9uZbOa9SvJ71ERK8N/+95f37dnxK5w3AZ5E3fRRj2h35HvCSW7fLgTMkEZ
uOcczb9QbeGEUOsfht1/DNhdNNNev2jXAawhtDMfMRY3fvRX/dl2jhBrOJf7GW+g
VYbU0leqHCOR2Wxritu2zpA6ZvGCCVEgnu0UQgBpSEOWztd9JIxxvballCPy8ZhQ
lBV7XgMYOITvA91/ef2JQx+1wch2JpmVLBIPyElIAlV/uL7QVge5gsER4FoJdYA8
UVt+eRpOto0O1KM/At02cwgH6iPD3vf+8/dQk54LrxylW5BKxPHXTb78AGTEacC4
uzUUWA0qhB7iIr2uVWEG8YvKA04KC0qeFWBw1gRzBo5CEfTReU8mErfzfkdDiRtW
uR0G9hL/sVpAolz/YnrFNpqCxw950o7uOD6gF7EzvCcA38nVzMoH6zTEieU7PP8k
h9yuv0R2XlTMH4nvYSeZqYN+RBzErLiMCXmDl0LfQ/XG6YBZ1ppamfa1xuAseGon
dhwmgPYREtqGfbXJHe+v1qRoQME9t496gLQeROTGqkm+K0OHIjSn59m4M268liV8
9CUhYRV/gc4DDRR34RuFNg54XZvuakC1omugouxrMB8SCDLQTCYiGOjDI0KCmHmR
7SX8/Yh84wqB2YthmYPqGsEBBd+mDESZYKkCCHzjm9Or5xdzr/udZAPa+6nyM6xL
SzJT7RDm8Q8UYfdqA9kJdzcefz4SKG6GA9bxccQYOYCAmz0/2AM96C9ukcCsv7Do
mnQ3KqcPt/gjXfbTdqg1HnY+El+ZSes+zxm7m5X0cB+mwwqMo1rvfsL+zcKQGGFS
76z/HEdsxffjIdFYRpj41iEN1FhKWPMUWOyJIARXbv9zIWPazHPZgP5C4kwVPsuq
xKvS2F7DT38b/NkjrVM5XRos3UwR4351fb82gxHovQy7ehLuWoZfnY/z357Jn6YN
FcdJ85eEkU6zOkxRXs5QB0efh8nfxsRYb+VURbMe5omwRZFi5FnBoBnZCes/S7/X
poSHTMfSN/0nR+jXoUVYhNIW/bn9mMnwzpCp8Nd+Ktf0c9zWDJ2hdaVjD6aQQdwZ
fCdp7GPsbK/2HGqc49J2sTieYQcUfPJ42mrkG5debgbZnjFGoJsreOYEtVMsK13b
Q5BlapMCKXfDEEbb9Tj+7x/os5lpb07SeKTQqdtII/kPfFWy+Q8HtKln3f2Q8XRk
DZetnUOfk3nFbfF1hJFI6ZUQRyd74sY109mHFhDCA8ML1YrpVe/LNPB4bcXv7IDm
0nKYqf3oeUsWytBpoLlpP9hu4o5TUPO0QYpP8fIFmP+iwYCNdO+vsrcu18mqN/nZ
w3STHOFSgj7VNowDtRR+5jbsf77P7pDEf0T2YQcqA56Ypg3gu4scbq6fpR6EhquQ
9kaOQ0ESh00WnKL6ymQqveqDCSHHvBs+gdxmsbqK+gvwBCSGVc/r4hwp6Ko1a64A
KD5k49ggsNWcpv/Dg6qeW3YqWmjCCrvvyP2GKqG71tX9iDcVc1HOa8FAct13a0TI
hSGBQuatO63ftbrgpu8QpooKI4rrNJX4YBGB2Evq8M6qsu2H1uq+N7Jv0Cw/u5ON
t0Da+pAKON9FgUNpzcLpr9Jl7xCFr/cAJqwUom0rTPz9UyVSY5fgzhqHYke6j+Qq
tkzE2idyO+e8cPB+J7AO57XZeqsAyI8hphcRgY0nBg5mEmgQJ7MC/rbmjTEqfZz6
PdaeQFpD7oURY94l4oPTO9NWsiwaN6uF3thjUYSndR48eRl/x9odGlpKthrLg90Y
OdqgMXGkRhLPkzGYcZklIRXtnmJTzAg3XPhBlcq8nwwinFLND1Acu35YiEVIY3Fb
CMxVcvFKeyXZ4/FNe1zSmP82pbmUxMwMugD4WK6TYyT/5LgyyvxGeX9ldNWbI8mt
paMxdfTFKfUQzSvxJnZZg01aIQuG6IoRqw0GEutyeW3iU0TKvrz0IAE73PUHOr15
80dTtr3QJUHGZTm38KSBerZXgGMX5zpOj9K3eCTxfo7Tea+MzuEsclYVdnoJhgfY
KCSOUovtWir24rvlf/a2LoLNpOFu+PvoKxGWN46iu6BUEGCkr5iGi2HEU0dJTTbQ
KEL/iHdrDR12qsPjgrc+sJElVwtsx9QisWPNq/YUZqtDCPIwHqvN4LF/xg18PTeO
HjrFJCT3w9sH7ZCKf5KxbwOrG6PLNU2xahyNJocZH5I0pqxynKP8GjuSlkWHHVvD
Ql1UWzoeo7uf2WgGilnvauJehPGY1DCjHY/4eyPetRZei/Wy3nTOSF50QHJZUXwg
qQPNbjYsAICXpMadMYu/oTAC7999SqqilShZhL09BOBQb+NUdDmfpYSgeKYJKOQq
fL+BiH01cwqs1w/TGP2hX83Bml3G1S7dpExd41dPIn7p12hLb6I3HLye0Arp/ef6
WsWhLXGHMCcZkJzmEeCatk4//fzYvRWeOYUzG+63iEHfEUrRRhe85lHwTYriHsmS
WwAD8XLJzN/QEOc5/jPsYdcn/iqk4RzhsyGDGbdCbNRR4QeipuYmFddCka8z/GSf
8Nh/8TuUo8jfAEc0RJKULCcfXUQgm54fERpWFbPVdTp8eVHVfvIyZbbsRvBPer0g
vN+xiCz1ckuFud2LSPu2uoH7XmDZgnHcnXTfmgbYOvyGCM86XwFUaLKou/OKCLfX
swQVp6TWvVN7ceyIhfwe0WT2v9GBUTvMkMcLgV7EwvfppeQ44O0mCok6OTK3CsDF
IimnWjzGdJ35GKQjdUjE/oW4mUc1wWn4h9ER+BezNbGg3cxggMz7NuH7sXVPr20F
QhQ6V52IBtX7JnGSYmao+FhVgsvQuEIEGhluiVsXtx3BOx+sAxouFk2lp2t1Qdte
jtJMHip86+QeTktAxK0zdKZG80hzWpTPssvvpj1gZRf4efnQKzc4HaIjd1upREe7
fhhuWEI5WDdNxH1JED0ZanEVJi8wy+uiS1nBU7j8hfDk/+7Y7GtnwGUK7PJgaYK+
/YAif8nIvgOCR5CXk1vBSuhG555XlpRKoAqR32jP6aIOp8LUI9NC5Rj4iNq+OkdO
6kDu0AUDDFShJP4+jvGNH8FxvbA7Yp+ayDsOY3yRybrl2hpbthV8nxFJzafgMVha
52zPm0teoYwSmgeloL4sL5fIfv2GFwnO77zj58WcydbsoEVz2q5kD1nZ2MHLo613
T54BayjM4TB+pYn3A7MFFQV8Er+J6/dbMnsWJNaG82LBD+fFAM6SkdZg3uzPHH51
G14Vbyq1ZPfvj49F9V9neNWBBN3MkIjhvyaOQU8AMsKueOTH6OYG6QActQbHa4m2
KR/7tXksFqfXh0MrBBwUiafNXSCBKAwJOQUjwT96d7AFDNTOs3dwuT4x1Pp/srKk
7BdOyeYkecC02O2KsVE71EkSTl053ckqiR+kWPPVANdR6743Bdxj8GbmrQRaiH1h
kUoLO74U+724vg4dpXLp3hJa2HTSMPKCLGr3lnnIDGaa1XaMvL67eon75dz4jyzp
XmbgbZDHv8gVLvG9PsgvxylTE6UJ9brVxfMDC0SMzrppnhSw82zS5yBz7kL1sxor
DCo5z2Cl8He4+WDhICJSQMyNPyz2UgWqfiCXgBn4p6cD75vVycTMAZ/5bomrlI6T
gqdBNTsvfvptyZbw4McTbLvsoJkhrtJIp18w+oSGwZEtS7S2roH7cfBDpYo+5P/L
OeZ8ktUrDM6Ai9C0f4YXjiPT2NthGjf6aafVE1kwfH+X49XvoH4yxs4rT87A55dp
xndQvp+HTTWcAXummoy/rVLNMbgpDaxD/HIKqxrdiQF3iP2XhN9PgRge3mumB7jn
DcSxKBPefseIcWGVwZM/UqJYiAbruGlTJfrbLDVlpVRMewc/Iqz8DKFAm4fONeRp
syMgw56Util0w7/7I5l/nQ/vlEvF4fIPmBYGteslX8GAe/w5FGDTb810c2DgRYki
Eynst/9M+qD2AD1rqaGOjZRyHhwT0LGXKZZN/spt8o1Yl1mNBVknLqFEhU9flB8H
HCpwJ3QRLwZdQH+tWN0KIQo15DJw+ZeEwAL6TPrEOWoxVxGDNgVhaNC1HuS0qxlW
JhAWFQQCp49Mm5Tkx3yk9869aoOQkezNhseks1Z8pfvdj1I5xAgv9hDH1Iddg5Mw
ILzsSzpASzoPsK5XvdD0kWUxT+XiQ86uvGvcAVFm7A4RBC7iTrcD0zYQqmc4hFie
oHV12AspUHMpn59IaBYOao55wHedqorKq6tgohQ0iM2e6a/yQ7KUEVRChqtC4kTw
WOoqX70nUJiaw+tsEAlfSG0EjCHuUGUs54pRPRYMnR1GPuw4HT0ZPEzevJKkTQEY
nVkPqmLOpUoOg/+MII6kh0XF4ivnNgmvKfYssfo/HjsfjsWQJs2xTTHOLtjkDa3K
XCiWr3PX6jhTz8qeom7goZv4cFTQ7nfmnbRJR0xrIbWGbyGV0N/eeUNnNjsFKKZq
Usb4gDrpuqh3DOoHwd22haNIWHi4xb2meNiQEA436qPvYght5K0BEW5gT8/Qqnvu
rMKj47CiEF2W8p/duihOP620IiWTc59RDM3KSQg5RG4mek3T6kq9wBEOmzIjtQxS
AmL4UO/UOe2/GHQdZ8WrukXTEOQVcEy0KjHLbVYiXp2NgYi2V+NHCIfwN4ejg/cO
Kua00/L3eJNcc8H/UzNjvMHPF5+/JJsE3XbSoSUWSlh1MZtVXKyGRDgkBUxIQPgm
5/L1+44uoSUI2VYjqeQ7duEZ7LcpLLQ1ZsHxXdWBDm39ojGEksS4p/GZ70++yjvA
NaqwpuKJOCfSC9u5azEwE0UsDIhc21q8XFKryIc0v35db55CjJQYAH3BKU++u6lL
JGDiluIudikhnc5UZMv6SFJZcdeTt4hGdJM6/qjw6ynfWjhzz2Jec0dkSE0WcHiL
0M9ZdAbFMi5jeWGJczLIdnjMCZZDev5MWtaeV9P0oXWGSfLZRxdY4VsE/Q3Wl6bW
AQxoKG0lLB0obsXqslvoiv/aYLeHSuviljd6vtC6JrrGF8QHZaZksd4+p2vipUM0
zuhrn9GUDmOd8lJxklrGYolR4GTi9FpWs7Rmj1qtGvVZqEsg+YRakSsZH81pKt/p
Uv2Y+h/u/Prk6FDUXLGnYs+BwRlb3LJSa8KG6ncroRP1UQR3PHPvSY/6CkCdL3BM
bAxxPVHYpq/2YslM2+/LvviRQBVcThXa3BQd/HyMNuT+ZFhphVW+enwoiQ41outM
ShcNy+M7AR204TqEHpdCChaXAEPf1JiaDAcb8tQt3uMgdyd5LetueTGPP3Guxgfw
vlj3k6WiW0jG7g/1L/ctFMRFMG6MVElzhwZAKNKWA+5aPoVCm+qeBLBmnYroyOCt
7dsHt/xS5M0jDs/Vepm0xKdylpiZOYdYKqSmIBNjS53C85tc/0doOjBd8nNi9mZ6
M3aZIsMbfpXfns2tyF3UB9347WV6OnQy1UZQ8xiZFENmrO56xswxKdnV+RiMiCC6
3gxVubKaUpUJIQJzn7zIzJSEB7DImYq4KQyHBXj/QonFHrOI8IJng7zb9GMKo3G9
ZpA1eTuWA5M1t8jPRuK6s9D578899WTmoVggqarTF/iJs3PmQGMZ9qAE61a4jHfg
xn1OfH8xYVFl++VKasQw2c+TR22aY+QOnwFhWESUwShEVVP76ME10H7PwrukkYq+
+TwmpvjpSFmojptIpMpbI7R1H4LeaZ9jXCk+q52bJMjM+zxORf/cYJXrKddJgzLH
axzxBstzUZjcZZVcsYhahGwV7zCdr0SlL+JJADpftBWeqnLBP8hZer3pPY/sSzVg
hFGIDzFEQ1HN5aGh/P/6DOwR9S9AKda1sHupUtOqFbdvnTfdEvM2XVDDtcLN+jnd
YSkfssXTl4+cwHqaHPbgWt89WDkdoSYTmQ+y8sWHgBFr5eXDGk2vredLVVc6wsz6
fslXKdYRAN4c5KTQAS2i18OkWmC5XpR2sukAiRjSTdTM25l6dyd2GvKfY0RFNVrH
BZm+zZS2ynxwsFrb/QTVgTOAjIYWv1uJy972mWfiftTOzdNTIG6rGhZKfTjuF66f
dfrm/SA7nVghnUE0tezu5D+FElqAyUESsPhFhmRMuY0xlo+qTKBKjRjqL3rJMqCl
rAp+xE+LSPO9tvRRaYK9lUw8YAr3LnORa2ETza+INO/BQCnsIBl1I5MEloceNWJS
6sR2GV1g5T2YTkzHHg2E62ETipMT9UoUVEBC2hyZJLItj2G7iqP5byhs2DfI+YbW
asQ26zcFxm060gkq8hebll9w4fmLL/mdOqGaVPiBr7kwZu8H0NZX5qLtXBADwir4
0edCtRQpmmqeSgu1hPq0FMQn8l5i9Fx0PM28XTU0tEC8dkOoX8JpHghyQPdhSPp1
Bh8p96nL6SQnVlQDYjAcMjTnZwMbmvhhDT84/1qAJSi4FdpAAnlsZkflKwsZYIg3
dYmnAliSx6Kwj5I2xTD2IvzTYYyElQFy7NFh3A615x0PDLqIiceDCuuZbTaIAJyY
do+WQnwsnspd9lRF9+sNp8UoDjNRB84WGEh7MBDo6bULEPoJRukvJflv8/6rjACo
H5ixV8IEI6uMebQ5APNYY5uPc3pBy7W7j+SbgT3haDrTgDXFmhIjwBItauWz0BoO
Q/ISB5Gqow47KgUutDtwuSmvfQVTUarNYbuP9MhKItg6XU+Byhoc+w+3ZJRyDLsA
HCXyLbJe8EOXYNQTvF7r7f3vbl/MTVadxdspCD1BkomiodTSMKg3uBBIB+3gK4uK
x/Wbdfq57E3Aqs4jIgOT/swPGbfItGzDJZwmUz7N3qFrhe1mbKiVgbXhygoufiCC
fcLTNCExI/Mu54Sm5pOI2SqSy4GutxSG2WkZJo5O+lgeynjzXJ0Z+PhjxxLgBR1s
WChEtTMX7qYIPdAJseCplUPnuq6ju5JeEUxFgCJGCACCeFzWUIMVaIEN477ySDCF
op4sV7XavhLfDawSDb3V+29wT02f6Zt2hy34HDmPPxC/pdflezvL4ZZ5yweyPOM3
lORFKIIp8mySzzQAdcMfSIYdUmpIlsmOoWVB32c37UlPjcqZ3N62Vgfu+LwtDNxn
I/CJQhxtS+12Uj76vaoiY4Cg2ibE9DCZr5IcORVyO5iXmPS31B9eBzFD+mJ4Uicv
L/5TztpGEZ4GanSmTTZ3wvvTNkWpo4jbD+sv+wp4SzxHAXKb9XNG9bM0zejPbMdO
/RIYA3JG74QrJL0poL1TuntbYrP99M3fKJ5TXSTiBhikez/+7E+IkwZSvsRhTcU1
5OZwJ5xJgYzVNopDarP7zHe6cFGdVnW7811bNQM73KzB5fWr7Isszy1KNArIlQt/
A7towGhUlXpO8hIc2uMlpSlk5hLqC+A60AStnVsawbn2I4+CrMJa+umkL5nfuX7T
ex9VP12g9ILvACK08Y2eAXarSnLUKFZCsBFUeNYdhsjN3e1b3X9MiCU5Cu9RaJtm
jLbxWq2a1x1S3DgrqalgT+LchWIOojvNxJPbRau4QTHtYmQLZxLpm3jXtexMao2R
cVzVcne6G97ElG7KwwaCvMG2z4b8YP/baTgfDk45w7a/y07dKXlA1naQBKE7OtUd
itrxnstk09dqtQqUvcmoQdkznMPtzBRAWNqDxrkLc14buSrz6k1wi1n6W2KDoS+h
86unFICvZKgEtR2MH32Fmm5wn1jc4dZWEyTWoZmFAZukWfm6TWHpJjlMXpxqseLB
LKn5Ra16EyRBD45+vVrTCzqkM6uCS3vZoBIri43U0R2BN9CNaH8i7G8PibTgejo2
w7w6CQujDAYDzfqAhwPVgv0jZ26gD0kGcrGdCqp6BS52iDZzJiT/Gx4FECxCt1S/
1K5J3XmOzXCNgDUSMd+FDjTL1FaDjkcX0PyCPsnHJ9/ncyDrWkSUi6EN//Y//Jrh
koTVG3w7kSwVDDw6FAIAMybH1PN/6OC2QHRpyxpq93fIoN7YBWzyyQt5dkVpfOJG
gAockfFiva3YW3fKxxFfzVCRGE1DvPONGSFrCCHn2nogT14i3BMeOcjKWoZI58rc
r6FenLuNdOomWI6vnwqLqOrRtaoCwv4oKlOx5D2KNc34uaEVxLoOem0K3JEmsN9C
auzq1EWarmqqmpoEQ+j9bpHwpsUBaNMmxuixuxVyh89aqmJzGfZXnpvQsHdH963y
/SNHdtC207ZnhYMo7zrUWfT6BadrAGqwxb2AkI8vd5XBxGH7UqqVwgnf5zKhOMe+
AxZXDH2hrg+KZr2uqFkDxD4+8OhIZiWZrKrFi5hkHgxswykNyN0FqSaNKCAdwJUC
2iSBCo84FZObObGxJAA/mbPvkKDQzkuMEmhaax1PL5y/+zrDcgsxe7/rkM91aFHo
cS/0ZvV41MD8xMNoJDRtd7PZ3RuvwV84cxsBsD467rDiZtgyL0jQZAU3bM85xYHf
ydt+VuDv52mQj9aH58gBtfp+jo8jZ96/3vbpY7XBL38oXSQOJxIeMBsQ2imhCzPY
v+ets9lKVzEIxzGuFoUyV6515cVjxotXGUjKWXu8QLP57Pk+KdsLs9hNUsT/BDz+
yigCc3njxyoDOrzwUnoGR9FukIW4XBzBNCApaRddipp1dbg1BAxjJ++FZgeQXrfQ
dmRfLm7AtRP8hXzhE/dqHgmliBKagQ5xeYwutg0MMAu3XcHc1A2wCbVIE4e/ampU
gALW6FurGUg3FjO5wspdiLVYxB3xPo/ulZi/PqCPC47zuGHRxbvuWGSFbHdW5svh
/cMK3D0NfFIW3Gb6xc/mRMMmPc0gzSrNjeKWySGLDFTmADNlNt/wvvVzOIrzix+g
cNIUbhSSvC20piXukno2+S7XuNmnW89YRI9zftwBJPi6I8VWgAsgOSqLuhMW3f0U
SIBpse4BI4gKVhG7FoNCRc79D7G6CYjb4BtHnzJETT56BKyn1Z9DcjmWfhnIp8lj
cfnFvOMx/K0zYKqJDEoOvtu6PFO4dAVVtFMwFpZT/ArTWhF1kYuINv/sWd01fIz9
DKdnLMpj03bCOsJHza5wcIOWGMT0EHN5Z0EPO2vz83ox1rrBDWG6Ss/joEqgmkFB
tR8yC3e7z6NJDq00JDy/WRFkNW3AFZYg9NLZa1zsa6W5M6bSHwkNJvDJMzmQCmbR
g0itujDPoZ0smStrOPwAabdAjdofeR45YT4fNA2v0QuRhTTIcDdrjFPgK+u3hYaN
JZONZARC63rY/hmTbuzH09jqG64meMiyMbIdbx7bHyBty0VczgsfhAVSZEJe7sXS
DvvjK1IqBY+BeSg7UWOd1eQJNOP4A38JfapJDp7YFZhvMz/S7YN7cbeuyumXrxN+
ZJn803JA7lmsbNBCXccCcQle+TcmrYjMDRbBziO5UTp8I5DBKB86E3+FjArl85U5
HVyNgdvgbvyAvEtyTt797rpw3+KwKQ/5bTLr1nviHO5u4ig/pBsuYfgat++PMW+2
ZrHNEjJM95U+CvxXWeYijUqboWNHuWiHUz8dq8V+UtmUlVMat11TPM3nsPQsis4N
3DAOQPUmd+SElsisbxPQnKghjW8M7bcEe3jjoB4selry38tXdjTrXA7EWpwatc4B
QIsqg/b1GN6J5Pa49C66SefhVGyVXKSNVMNBi1pm6DQsQN36Yc97sRMdkj0d2ZQN
33qc2bmdUTHyFmaQmqMUW/fA88ZZ0IaNtCaycG4K+H5WFvEu+ORduI7V0LTGGu9k
ZIwUIfSu9NJu7Wrs/6gsL7LVGKhfs5cNPSZaKn+fbXUBIR60cIWuYb3SLzLFc5vA
mQm7/kcObCTtwgLClDklJV7KWji9bnGJWs8i5XqrGlOXegVmPQfHfstyCib6UaNw
UYWHdjJFWyDP4Ej4ULhFiukoqaOJKVoWAJr4ma31nN76EBLrkledEOV3ybTJ16kl
MxCxcMfWlUIc03pXETNVL2vCoYqdqnipHQq0W6cprAmoBQFXPR4wkjeJd/Yy+mvX
x0Vqyxoh1vFCnQnpmECP1vpGihYmSXMSNdea/fQ+2wWawsNjk+WcDVU+g30HrEnn
V9A5fUkNLfDITjAVyFx50snXnooGUBpo3MzlRDtYXrEfZg58qjudeK5qf3SolKh/
PTJm3LjB2IwMKdCEGxyCqid3M6G7QAgGovRHURp6qFYjnNRzT1d4w0Yc44v2ZO2p
xvNeVGR1FI5V9yNFLIy5haT5/JYmhxrUj7ScXxc9atqJqBRPITarPQKFWavJxOpP
FVSs0rAmJnUoj/KTlI3MTP0Alt7UWQrYUQCdQxYbxRxm3VngAJZqvfvQKN0QLxVX
Cvaf2yTrZ77plusGpbthAzFA8sfx77FqdUzA28NSeeSzZJsUmtcRegS2tg2xosHB
tNBdKTW9KClVcUZDrzfm1aM8aiJ0mUZ+lDJ9gkVO2yztYDD6f5RmGbiVLTCIKLu+
PWy2yauoDWXtDthKOzLtm9JE8oQglXcwINpON60qT4AhEXkqaSU2jzSTg1wGotta
QQ6Gyu4meryT7PFENWGla2yiPGeXwWl/IJuIUitRnei4F8Jj/qTW9vGRnUz8urgC
vc3T+isPTJowDWai/LS5RhXNViUWRtnHU/SOjiUbfkh+A8rZ5WEPCMZcjIGhcYhq
G9OjSNJmbWeepfuVkDqW1LYHLLm21sW16Epq5jK7XWo+ZoTVxLfZfoGYUxPds0vu
KcTmtgneJXHvvBjY9ASw8BLe6f+D+Do9o+xFeJci42DfoW8ICiMMz5Z0sKqWFDD5
QleYdu7LMRJvG32AjJShpSCjbXSaLbFX+LdJH8BO+IC7iZXMjjZt4gh/NLXKWrvN
TtwwST75zs2PQabWBAqUFrKvhZhIVPDdyLih1cpjiNSCrDZqM84wgELUqUJwWBeC
3+/3bGpWMxCW3+FV5FiM23LjGpQQegDSGXvkEv/9ma05h4FrTQyjZad6nkfKenjo
OGuJUEPQj5fiEx4BQa+sKTpyhYolyQfJs/w4UavO3CHlsBG1+EBZQc+vQvjF8Fxd
76Tbjb+Znc1wWX2ASQK4iN1ZHHKC7k389TPhBWTZ3LLqt0kHMZrnm6DBKla0dGqw
D2rqG4FhWuLA3hPcAvMCUzvI9VGM3Ug0yF/bkAZfmQSM3IBT0HMo0fGS286nb3Jv
VBsSo2g+iBarp/okiD7vUqfq5suSsrFSdLZ35J2DpdPHqfxv0b2tiLpF2PZ/9/cC
y09gbVkGM8YQPIUjbt8Pq6cFCX/tDqc+IyCALp7CCHoSXJeBJgAE/aUkdqlMJIXi
NxH8eQhRzoulTGen3sW/0Heb5aUXw+69DFofoJuNAfj4IH5xh/bfhaRzpW26C2Pq
ibfczsEbrnl2/FCNmFqamnRlpFl8NbrKPOv2pIpZm8L1KcghQpSEv/21Nivnoo1e
yrS8NVbec9RH7VITs4I1bjllM7WqfkGDh6atYqG3VaJNsqe3pgZ/EtKC1r4CT1u/
uncgU+pA2W1QKDlmAkOpRjd0cLkyKiAFx54NhgsJ+7bOdss6YrB9wyMuvgmfENWt
c9MAscNddsqLKZkK22iR0okt8VlTzGktX435KAzwWmGDFgNtT3DyRiXkbMgAiQ9K
L4T15brjMRKTgXx6KJm5xy7ZYgMueG60Zj8Dv2DLj09flHFjZ1YYCNx+3LTo5dxz
eTjASDkS/HrQ2Udx42lADkEdnCcYdYixGpAYYcvC+xkGJbbRwHeldK8WmHyLt4Lo
XmufXaq2UJdVZfaU9SmQUkshR2SRU5zrw8ThHPb/RQRe2JMtV3RccQ+uJ+4XffY4
YTaX38wfWPz2ihS0Zd959gl3IEat1Q+6ra/ZkrnV6vHv4WA5T6vqv4hs1vsyer/1
OSFo6f9teVa5hygqvx+m+oGlDlD11fcBadN90n2oSOBiMaH/sVWoW+j3PfHWcxIF
5NOarjSRVeK6qWtOjOj4lQAjccmioJKx+bG6J/LnqHz4Lmrhrna4MC4ko4vdPjK5
9bZH6ZOsZIXWYZ9Rdui+/3OrRhBwFy2VE0dhhSqqQXAHPdtSPj5t3749LbdITYLY
WDdhxhz5vHpshX4XE5etCJ8nw4hwRuLJ96mKx/naX3CkvQLhMS1K8thHXkF7imC5
FzUOacOMm4+J79EbXvz1dya1zuPu7NMINMB+p9wyXR9SndRiiMLsxa756FIXYr+3
6iO/74dSUH7o3bArOZeZxtnaF5gGXhqxxarIaP9oGlciZFjQXUYcz5FRaM2Npwdy
k5gFC2BtNj0+5CuG3Sg5rU6Z8P+mGTIzLPw9fo/AMdJ7D4bXaEW6pLL/6O9alvGn
BfGFBguE58w0euRb30NgQKZBsVEIfpyLM1s7vR4/xyJE8GSf6rr8cgfdFXlgNkVm
Wkk17HsPpOCdPdJ6oBN2bAptOFNNU99r/xKyal4T+O/7cx+fMPcyZqwFvDjMtUJ3
JI161NpAPhgzWYZNCmemmvZRwh6/PLNEXZmmeTDdTuDSbIrsa6hKFQWpzFYKF0Wb
+2rqxQ7cPKaCEig1y4jJf5BBRHjSjQ/fcR1YeepV2nTsub9jwa2YUQeAI6oUQ9vf
M0Y+o+DRLOtah9Ms2CIcRQ5DwO+S0i+D54Bj6umU+2vDU8le5N7OTvqks5yHIfyg
98Uz3rZjkutGGMeQEFtDjX3KE8HAKnxyrVqbTe75JF6qZtNEinB2r3hhsHNTzJjZ
iu9oK6GPXbVlTEYQCw1jz8f6J5jHyl7i/mV6Q3XuD8Lwz/m5W+uW7gf+WSi5dQms
yt72iniqBV8ouSZ3wRz8gPuSgZ/lCsD0MC5Uzhy+zJsFB6pqTKBdNrx2qALiZnTW
coR9qEI3bp8cEN0suW6QINNfJuSPSKCPHP93xA6e3SoGozIcHGRVRQRxtouKzlwJ
evvYGDvE3JEefbnqlHrwXp0ASjmfa1JBFLDMmn11Q7FgnhoFdqpHt2knyTPDHNWE
LFnLJiJL+T6a3o+xG9N6Qjmrp5AKiKVLdqhP+OAjFDgtb09pwxO7Sjg38HZYn+xs
XAVzj5W2py3OPBT7p78tErpnWKJnSDyQEeoduO6D3RCvHy8+RhWA0vcilKvQ9eqv
gmamzvfC5ozDofGzP7wOpuWsUyI1YpNDfa2sCg8KNuuJMWNh152KfRuOQedW1HBj
WHGdAjbSWVuxqQiw/yJrqZ1RcJ+39bHl1WA+4rc5Wtt3rt+pxPT4mEwsrNQVhFfC
65CLkhVDhtSt7aw4xal4oHqer1p1Sdkq/DrkmsIAwhglzq0/fHAY8f4bGfnS5r16
hUdGzj4jQwmHK9h39Gs7NJDE/0MnQAuJRMlaI0c9qp+FQF3mPg44r7EeAnLrGifr
UUER1KPKLb9PiFjIw6ih2aixVNc2nNvolyHe1rssNZRLkk9YjTBNPLddxutXpWb0
eawac+mefpEPtTjg21YGFh49rks/18WwaQsom/QITmsfn2fip/BSSm/F7/HRmOTd
ZliBCSSdsTMWp7fGLYshTo3Pba6cnhDi0FxahPiSoNz65lEpkvEK639HBwAjvQEQ
0qIgrGUbBsSigqCSCa390vYPFejwSkQJl19DgCnicvkE/KKy3sWE2d3zJOFUirBc
odHwNU0ijkHkX13A0m6QT9OCtKfUJuPmL7m2eS3Kdi0B6GSqdIJHaFWWWLHIDBOP
xONEjELyw9XW8fSVtgEYEQZLb5wgpxUMGjF/bX+u+KyQzEtnDpW4G1Vfc6gbzHnj
h4OUjbSybXVhs8SD/DbpoH2QTh8UoODW4HNMjyRhGwFQz2K9j5bkObHLmLnqJKeJ
2cSJeCWIORwWfZfocDSPGFheUBRh6D4Iml3xkBvCeX0KRKOJPhXcMLzYcvUVO2ee
GxwVcxuisS/k5sEkmOkdGn59G9jjD1ojH09Cs2ajTl+J3vBpXSSw1pvj/7lBWNER
lG5zDIUEo9cgJyn0gcU9jR/tltJzaVr39n2gGcpzTMdOr787pu87UCtDhCU8jQ1w
80Z2PoCWfMiUT+7lD2ZnGhmQzakz32m/3mABApiA6N3qnedqK9UqJOAOb1KkiCSH
MggdDMP+lrdfEmZ0x6caNaTr8cqW3xxAgjZxs3RaqT/drY53r+PlVlj+iHsNoNtX
oYssBEvyxl7+qIQlqbY8mMlbwQ3LhZ1cRUDV23johbBblBjD3JC0Ghoijj2p41mw
o5WkARuWTUblr017AJSCev9ryf6TODf7TAgY0ax206apv6G+RDtIEU/nvvdQzrgt
gj2BXo7nZElQDRh4c+wbG3UfwjV9OqO0y5M6fhEliiSpzjwowWbDSd8D9uV+q9pl
WDxlV3J1gdKywv2CTdPx4FBbYLSdSmA6ofuqef1Im2XtCNKJQKgjrnADJ8O5m98Z
8H3C9HNKgAFsOdME9+hgj3m18KhIB914e3joMh3utVFuULgb96DvOMQDYo5+n50I
22+RmnGSP1nNEKmzOknhUgt7rjm+zbhMwKy3kZKKjwVGyhUlJdx3cIflHVsKSqZS
6aHXEomYAEwWLEWeJxiuGWcvjpbmsCYuVh81o7/CVyJCkbKu94m2k7ccIZqQZugn
n7bRaaM6uY7hOlSA/IVhfsbZph7jKXc+yril/tGOS6LZ3RPn4eZlPfyWei7H28is
kBrpF4bFp24IR2P0NCYM4y+lf/w1uut2gqfDwhDj2LwnG4WvSAO5rzZIN+5QmaJL
egAMx1quJTjK3QQfpR/FXqzULbnvq3rNSfuNDM+nH/PAQ1fXnTljbOVF9F0ZPKlZ
1ZZbtGJGC86QyZAWCZKBIlK+B0b/EXypBa9z4+dwtExFkFpjTk3bbrfR3Opwf/zK
r5htjGgLXqonFF0Tm3ZNx3mTkK7V4cFB/1hAUz945L7K4rAoowlY+SF9Iywsa8tR
/f+ix/9fxl4zYh+7ozf5s821Oee5LtoWKBvtROq8zOR9O5PGXY0NQ+6H2v1RGcPU
JlkWnD9b132afJEYcSryFVYq1h3O6UqyryQ2C4TwD7FqK12CE/SY80dW8xlpZpDE
QZkfoHan9GDU0nx1t8dLXIK2CSNfAGUrWPig4M2VoaoWrovLFKFa2P4La9957xbg
N4mxcYX0JGqK4tBSnPvZYGBuMA4vPDgEcFoxPDrlvZQsTcTPJim1pJLvgPZt0/lC
0KjHUkwNK9KFrTgbz9Z7x0ncN6RvP2gmy0VMVO2QFL7pQCdj3domMlrscso30QzS
VcQC+MPxwq2ZDXwWYmaPZ34lHZwCYw7wqMj3TPb8zXKDE2Wny8liD0gbqCB0iG3w
+VVqMG+PSoIUgC4Vie0RJajO/RUmaDLhnkQwA/3p1zlLjtE5o7FwzfMh9ojaxBUa
Ilt4ht6qTcWn3yul+fnZYq4wBroy0ITPSPEfSt8yEe9DmSnDjDe5QCJQf+1rmecS
LCtq7zzBhlINyl0X6R46NT4tKZjA7jp3Rm36mGu3KSY8d1I7m9nJoNG9LHo/tbAi
xp0VWUIbeKO2qpWqR6gNPmG+nWSVVpN7CONVn7Jf5c6dTGepJPn6JdCLqUXBaL8R
zsiiWf5sFBsvEpjKNdeo8rkZdpI0NexWokt+KnUPu7kaZotm6Xj6VmRD/LicbBU4
2vlLG3sbv2cUptg2ffEB8nrBygX+TOa6tgp26DYgIlwo9Zyw3FlibEMk2JOK1BQo
kt0G3Xi95ZpUcnMPvM6qqdoJEJFzVDvDg7c0QZ+gRg+OycjQMY/+kciqZYvVTLah
lTavsggCItudQsHSIDKhKK8eZBZD6E8ITBm0TJad/TW0WxReRVMhoaSSjVNK2qtz
atD3EwxaUzKqQmmEXOfRnOpFdyMUeuA6dVXdK4s9djpgQZSTW/1ioU1wViauvuyQ
3X7YV6eGU/ZHftk/urmSTYyHEfMGLDnTaq6Io8ecDmD/IpR2+K3R6IrjKYc/IZXo
GxXfkmIOy3NlBNzPKD1KjSJA9tv3UEDPfLyalt8fvQAYcJeutgaWa2fQ0Es5Lf46
wFO6u8dCy3Q80G5vPZQ1q0HiFYeNXibQwGbH+PldMhJVCWtNcJTNRpEyp/qbXBPM
vSqAH07ZqWH52KLeUzRh+hbSdbPrkLwtysw4yS/6WOU5uj0TlrLfqjUrSaIINMhA
26+LU8eGm+rQP1ZO8+BPZ6I5yfqHH2iIC/80GV0c3S7lV8B2Zrw5HVz0wJCsS4/Z
nWoey+st3Kg93Rc9fK34bKLk19oG632DAaBRjmgB66xEfc2HY3y2d754jSDdxR9e
lc23BwU2m3RwnlJbkYWq0+3h8yf3scxmjNc77fvRN6e1yRYOzVVh/7rdxp331sIL
/tM05j1UE5X378jYGAa7PLMZvAtAL4h8mxs/q+9hvrdWgY2JrNHSfmd9O3eiiCZx
0NVT4jHnZ6DIMRgRlWYzxD2ZWY/iZ0KeY32AAcfLj2HqDuIPGa4QRRfRcWuEyJSR
R3QhQ6tM0JoUcglS1C5f3I0ISrkKSaqp2PE7REtpTX7ZlYJzZCw42/19r0aTlTmJ
tS9QqqER1M7hByyp2uY0E8md6L3PVne69Ax/NEV/tnZALle3hC7bRHeIfr5Z3v4/
MVEmeA4w2r7mW7yj6mO4BGoDU25kvEU6UnHB5La0/DNK56nJ3BMo96wD0eSSn2LW
gDUHYXSYgmiBNB4dk+DVTlwURekgqzg99NSa3HfxKiWAJ9MAA+ytkAdNU79KJLIk
kFNA1c9jgF6StKA1FMDHEDmpMFCJfGbYAImoZatRfgMoifYbnA1R+3NwVfT+JkFD
EBfeBOWdOCKiyD5xJK6xly8tXBxIiy5LZaaCUKKtiJgMXk6dFDFrDW54YebHISwa
9pnNvChzmxyiZO+kZDJeaSlioOWWp+jO2Ak8cogmyn7nNWGyVQds1SFzXym05b4P
a1qKZHJx55VgRaET8iTOJIB3cU69OvzfJeXa8xND8qaLAVTgaPCh8RygZYw24eSn
BEzpVnJ7Q2dT7S+qw67aKIpMDVd6+jpTgPqUJ6yLLNY6fH1pvafmnqm9gBF2luF4
sGpNKK9baYj5WmAfJfmabLed/T+kV8Avz57Ce1KpLO3z+W2e47MHowI0iVpE56pu
qoZWMEiJ5l55UtdDOsItCAFWqyXEMryyPLZQEgPTBbjUcA7cQrn1jTxSpn0rMpkM
3BZdUX/9fCyt4EKYRsW7d9DiodSwsUAqowuCnJIdBWJDMUFSltmhT1olWvsaki6M
bA2PNZwGdfZEFvm4s4+R9LpUJhfWYr+cmzy3xmappcyVycyVbLtWMzk2wnWIyvO9
JI22flcvJ4TJOUDxtfIsY514jBgb1BFJk/797yvapiKbEqs8JtKuovVndEn7ywv6
t3Im8LORUnrxkyg5MaEviToGSf8UW1DWNg3W/FnLhJnDtA7I5Ki7UL/IINuQ8FNd
QqZJ7M3eachGJlzjUs/K8EBhOX68SKje2pM50kO8l5AFsUhk8+qnNlRiJ3Ig8wMV
uM7fnWJHWP8ZJYOsmLdO8G9a31rUwT8bHsWOIvLucNMtb0+NYW2Z3NnKno8gxM8C
ZJ5WUrIrgxJLeLfPLmVmY4fSRFa8QInwnCIdVA0k8B3Sux+enfQhJnr8AU+GkcBE
QAcrE1gD83SdPZCZTppJCNfXpqJBdgKTCqc5b9Upw2dQKfFWJeqxSHvtYAFygkPb
GtzGhQAuz09XBGNCZh2NAYx4KTGwQjpfIr9CtR0+QzNzUL+tVqEg8KOuM8EOWxOV
G1sLS/ZFFepWLxpb0zgtE+GNDSZasCQWFU5cy8RVO7ET+OCNw/5hutHdNwBN67aX
qnYDRjQXEvmM+64TUKrGKF4qshvp1dJ4+7C0LOL7P6ovSNtAPoPhN3S+ZQWGvWKn
RPrBrvMYB58H32aILUcrAGAv9octxQsbsYhxHxUOIbikAlR758VA+gZswXXICTN8
agwCO2MFhg9HreLYB1SZpMCGJtPtjAKooA0GiZa28UULzejTaurvMazjawuP+3yw
5KpBURepLzRlUPE698GbTTHK6CPRHBycz/tVHFw+EyGmqoBe1kG1k43+Sy2x4R+2
Kt1wWoBJIzi5UqWPFunr3wKhx40xK5iBsaWuthTSpGG3UA84nVUjO+dPA9xLYSBE
0Y5xmD4L8OrkTk7i915EbQ3eTKLHTGCLL3Qygbj9k4Kk6wFF67beK1e5HrltH9ZL
tj1pnRs0Hb0F2jg5za0vZVB6c9446w2Y7vp5AzIRgQlUxKxdJEJPJ7Qe8InwzeiZ
PPVfwLQLA61RDtIMqliNN2jqq4iLTTOsE5g2zG293SJoheqpFMGDjgGaHvt49cMl
77hjM/d7H6XqqwMJdQ5Qvcz2tUxoFticR7EGk7jsaX6FuUFL6h+DAOMmu0e8aFCj
Q9FPtklXzuO5tYVJLUM2EnyX+txrup+lHYIpg93VKkTBDrJlOavl7wnu7BErFm7Z
kO9LjmcLShQwYsLX5LCxydl2hEcM/sPUQ2qKm9Ow71XxapMPCAQQd7irhpPQdD7w
XyLLVcwUSTxZIbfRc/Ac0bzNPbORft/Qx6qJFooSbPFjBMAZm2FKkrQYCXj/9X0i
Ak9ip6JEkCnwO9QjALgPdCa1WB9sWYPrhQPwaJ0dlkfkrWTmdfgzOw0PpVEwc/NV
24h5mJI0ZGOtdjoNgGipbms6zOdt1lwgHj9DiQdQ4sJqQpt7W5yYh9/dehXLi6jN
FuOw+XHDdIvy+NE81PHMNn4qSIu6d4fzqkNP5WK41x5LwXxeRgdRygs+uXZql7K+
gfxj7GE34UhnNGvdsQAE4Da03kH6n2B/AG95/7i5UvfygFcLwLWtbWQXrduLDfYG
/hqp8imrWjGAwAG8yjFa5X6JFxdUQdbtWXZAWe9MGGnPc10MDvRfDjrEafWwuDt9
U5KBKGbcPU5Z1Z07V4OM2CCChF5srfl1dDN/LJBcnbyzgzg8ecR9X+qRRUmziTJT
PNr4Bmk3M3SiXTDwKZ48HpR0W6ShzD3tmEnwsZelNHxdFZifMbr7HNSN44aeM1WX
uWURDGFDJG0cORBtc7QJCrm5NZVyJSiuLydm60GRdnXKXszbeExg+NpcCCfMaPW8
GUci9ynTpAExhEZraVCppaDrl9wkhDyfzRiiQy3ExKXfxGsMUNCAVHrBZ7kEVaDv
WNGiIQomJc6/l3Yq4Bk3vEaJS0m0TG2OEsm2C4td0IrVxEBsGMxmgfK2NGsUlA/O
ExRJYSTC3nH8gTlt1zdhbY181+AY1fIwvS2KHnS9ZF57kaaiOu/p0+glQp6Z+S/9
4BGRFD5Aj819Jf/FFWMidmT18eNP3TdtWNwPJAXnXv0a0Zu19uYCZk0W09HQcu5v
++12paRR3YAdPDGI19PXayaruYV9UbbK5OVXyb/a+3gleoI1Hmzt9Sr8TWuj/xJ9
BAoq7P1V4465saPva/LKEZMYKBefzcDWkOx6V4RTyweotDjrVX9SKA8cD4KhoZms
cHBH+7EuKaBoiAy2XvPpyF5C3Id7QxmQBiSAe3Tt2PS8a5QoJbE0MdyLrkEiTR1Z
rw/38vI0CJDlCb4skUJXDIgS5g5l9m+I+MP9M5+fULHAYWEqqjPswtb3x1RGe8zg
/8rtAFsA0xXaBs68q1XqBQfdqahBhHnVdo4P9GoD+PCSCKLKnjSFgtQWafX3Cih9
TSxPwy6O3zgyICj341T1m7WZ8PmKVWdCsTTSCPhWheYRTXoF1W1U0s7HTmTFKOQX
Aq0RhGCplkNh1ruMosHzCMMahsjpVYMhlV97oEwIuxTVnG3wwG2yAHBIikn/sbYx
rdvkm8iuNSKpm2oU+tw90ebUmqnl5Z5JWE9iBDpDd6CqamkRamSJ4Vyt+DXX9vyr
JbEv6pMZUwR4Yp12qFXKceZPkYnhIE4Ao0w9s9bT4RsBHdBWZdSPjUvK9dNXCQ8c
JrszFmot/x5/TY5+Y5wb/4J9t5PJdbhuE/GLxTk0Hiw/675PQwgsQilrUMR4oDJa
+uEufj8lX3jlioit13NkBvAF38rm2fcACrKnWZuMl5r3O9oZ4+YLiKxfJrggXw8k
7kYoCVLKp3YtgSxTgDHJJIchhWmh8NR4qUhcoy3E0OGA6jbxUUgSHPL4AZ3nsDqe
1BrHCvqQSJQz7+VoYcoovE4RMD2nLFWi7hM15yOIxCfJqlCrUrvG55kAP5e4Y6/O
E2TkWviZ7rHb6MBtR7lLY8Vvwc9QwaIkHw54LpXrsfMuyGHVC5E/3V0IfgV4sJmN
Dns0033m+2gUwpNDCFU6ojzMmVINUSIiu/G0pqv0DzSBSLJ7lte/G68/t0TwdKOT
PhKN5xarPhQQRLol/arzEex/GKIU5kBarz+vcZwmJyhD0gTIvLKMH++CPsZGVhA0
vnDjYc1tX9aK+pSaclumJCr0DLPEZ/CSF69jvsXcSJswKWVrRx9UJ9tK7fkn5Mvp
0tAGCqIdT+E2yulYxioM1SQzzRsPclW/F+naUoY4HmalkIbeNmBFSrLR7ikp+uFP
9FXB/+64rr41a3z/mHFjjLzKwznmQwlxOFk8Mg2ZG/e6BhiJfKMckoxRNs1wnu3D
81xa49Ymr/LQktnd+nzhZ2Lmmsv0lvrVTmBAvaB4dL+dWiEyaaK1qKoGO3Es1Byx
GXvEqWCJYrctSFT2ZkABgUbSLHQgeT467gUOhJ0SNmr1gXrBfTA37gF7fRsyCkZA
POZdKYPiPF0KpAx9s4DRPtALOmU/w0UA8kZ0k4maNktjuQ09TZEhSSgjEzkjPWS+
yfK0Kzd+tWH4spnY9GH9O9GPSyTYrKziwCGqlY9bdlrAk4dIdKYkK7JzShozmHTU
IeurXvAREXap+6Jfqre5CJrvogbZ1FhuKSoPRmlyh0z+8KVb2DBaV386id+rsEuM
dA+F9AT5zT8fJPjIFXhUsU+UWIgWjC6NluDlSQl9MAe6LrkKSzYkek3fXpcV3y34
waMfRK4nDjyKGRTGRtDm+XNE2yCOGn7SSJFn4TShbCrT2g499WTDuI9NNAwwmMZ5
PNKrPiuPHSmLngBOdg2qJvBm2eQZ3PGWsy1CPtt3YfEbv0sC0d2fcMItGlMvGIxQ
n30APy9mDeOhf+94MBJTniPGgKHZKp72i9D6cY0gmt4yEmblxSmvtmysG4DZYUmP
A7c3WgmDL4Ozxj4zVElQ+PzKQe1KroM69+oChmNCCNkfD2Rc/zQlSXVtTlIBQVnF
iKMUcaOoqNCEDQZqU6o1B3SzhBr/yZ6FjzIfNCDV8AO3d66YzEdrKVGG/cm7uFYU
thbLo+eK5JmH4ksnT11OzZUIqBF9pLxRO4EXvZwVhokJsydQ5kz2nNESryXhqg+8
KfxlrDfyN82C+Ve4AHjUd3jpBVoo4o65oxlubiZpt7TxisQyx//3Od7pafze5RFS
QK2wUGLt4NKq0nr47ndCR5S50kmvQ5aalL5Gn+2kE2Ivi+Hj9JyxZVut2uYPYslZ
3BPlT0tcYyAv28uan4zmF1INiEeLia9ogd8mH3Qz9ypzKJjL5aqhpse63XQO9xF8
KfC3HcV9dHPBpfYc/YLwn6BhNCnGcN32CpJ4TrJOWCDyfGNWMiMFfresybhhV+s9
3FEUtXEr8ehzWlNBJi6EQZ0cx2ZNh0RcwD18azkUDtk+paZfeF9AOpO0fWSwn7LA
FGOBFHvLyx/X6RhcxvPPVPdtKzmODm2lgY0rCVrXImAD9EaT0dP5ULK/xgeQrfQi
d6ZR1ff0wDnYWtL3ICgdReXvRLQeA9XE/vQvK49lExs7lp+HiPKL4XmYZpBhzV8a
B7+1yPwmOABSz52ixJr1xmjAzzV1nw86Wf+sIkqvytThDcbQdcJSCd2Q/2OT9oIL
rXhWWnC3+hqZUxew42/jxzomqzlU/81yMEGqvxMRRqqP/mnzT+iTpm1EV7J4tUCZ
j9DquZIZ1GrULMpctT/oerqGT2RbhLxm3OkJcU6cWv8EvcQ0fyhHZLpGV4sMN6/Y
rUf0aL+ZpuBgnMl1kzf+NmuKg+itLtXvMSCQWOKuAKHub93u5DcB1hKGVqWK4/ou
6QP0NuNRYBJJVtUCVhBMVHEdO/rltMsDb9aZvMI+aixMv+h4BUYCdOJAn6sjw8Da
ik9KH9Hr+bdbxoOGy7uwiH7xqdWzEIRRR63syMb+Lbbij+3jxPleKITi0nfJGPUX
vwuheGKaeNfgYxSd4K/zsedXXf4FYFiHAokaIYe6czF9YMaEu27I3vitR5M8u38D
QrziWXZGI/X6HGTibdLKEAoRxSYifkTRak+gdEznkQuBhSN8NR5XRA66BDu0tb3h
eNNlPYmzWKsPBtGR+zlzDjzEoRfFsuaoYeYj3pLAaM9k+7BPTSZMG9q0VdSXou1C
CGjKiXKHHVE8mjN5R5W9LgVEiW0VHi+jzbPDy6WVDcczNRA9WHe1SOAhlf10XjS6
pFmWha6tCziUjp5nOBHLjyCNkLe5Qx4STUK7RRR5NUpmva6q2lanP1s6GD9VnAVL
owiVMKcmSl0dnEIXUUSdLQMf2XluQfdZ52PycZs2mG1e5DdC4zGzVMwW+C97Qx+6
N2+bhSIk77xNvhvsjlDBjkYCi2FGHJoe5+yc/RXAAaSzvMf158kM23iy5z9E9yQU
gpBp53eOSXqO1JoFKkedeKa5GdoFHuavDsYvaoXc8XKmeV3GtMOX4mVCvXTKNAl7
qxPKViHaLu1iaUZdc68smg8nu1O6O4MzZxPApCC0AUvzAKBGm15SfAgUdhgd5FwI
uLyr+LvSQhuadK6C9xCiu5M1dWvlcg8tMy4ZeODWOLPiBQJYmuxilvCtVGttgNlL
oX+7klETO/qa1ZcCPDuRZ9+igp+ys6DOfqaTt6RlU5pkdnygUc17+lhwJQfUIv9V
bBS8zdUNNUBVNoNW1g2tZOhMSR68BGfatpVOQAXhDIXYWq7TPSqAE7zTtBZ6HciA
wJ+Jn9QAsC5m42QFYnJ+jg3PrIpNAU+z0j0cMPAgqNpT7//vt8akH6+PnK5OxzMb
I0WxWVP4jlWyQ6BzdYG1Ywz6IdiKE04QHDV2N/BeIKl9yTTe5Uw3MS1yrbsTitiV
LqY6xYnmU8xiv4i1dVj6zxN9qLJbmC/WD3wOGu0+yrKCU9T/cWA0kbOtYgCgFgho
dRAHlys6l5F+t4YvKgop1NIaycZKghZetA1LKjWOpab8EX0/P4VBWO16iCpFJfG+
dVpu5H3u3WR6wpUkj/qIn6oyYJ0RiVWclPl9/af7/vuDiyUvukCpgN8D6iyhLeHw
y3UlMW9L84xRUsA/7H0Bci7zpbza2Jz9SO1wCcGReTdkSOpvh6hyoCgIc2H1Ejoc
fX/QDYAMbPbBDAfBC8Vgdm6MlB9yapj+vNJrkJ9xFpC3xl24EFVdDpgvnbLEKz5g
/Y50yyg85TprBDRp6TvO2sX0XDv+YdOfjsdX6IdH0WUnBE4HkdLFp4AegMeLVGTQ
MhfL4I8fuE79eIsfwdeyQCwhV5Ap1YEYjEGhvovslKNgC2vE/cgmC8JyBJMMxmJl
anRsMDKw3qsHBR/fuQcgYKBAMt5/zMNYpbfs/RwFHYnE/yFAjIBlrW+f4qIveX9Q
MUlRcp2ksPk1/YJmicHL8nNOd8wiOwTQGFgDt+XWmZm6AswieMJfJq1QsZSvKDgZ
KgsYU1l+w8tB3bwDUZySX2TwRKo9CreTsk0cXWHCMGDOL9NdMx0k1CKTTiuMq81/
WjUB1bdBPBnYNfBUMUUxMzgEUMrxYXbTND1gTLjUgw+QAbfx0rr/rPU4z1mCTac3
W7KWLEDXsbCLAAyrnNUK4UqYs8yraJ3E335odgtn8hAHNAn3DL4VL+BcOiZ7ZcE6
sIDntxrozqWdLhu3E1z1jmaiPb47q/5ySV0FPpORRjmx8oXlCGtBW4xoQiX6fRfW
O9O/N78LWE5Van5o80ruWvegewYOH3oC9KxgVKxKw2ytBYk5gKEw7LeM0Az6s16v
57z2lmiMWuNKo33NZ276Mb3hNZH9s9GExLO/twRUawx8M4KMMD9gA/wc4YS/c24p
s+k4+hsLfgrcbs89xCTV5z+fJyfx8Jnd8RHbBt7uYMhKUUCUFdVfB144QFNdbbIH
2l1PSykR7VclBnz3aLHD7JMxhrRWJuHW/tIRHKTR0rZlFnMq+qrxPt9Mf/lT2mGE
gYhzIdyZ4okYgLPG7FyUSD73gAEx5TJ3MzN30racN8GnOEEjcK3hvhVhVDx16zUD
EfL2T+ndwnvaJqmh52F0OgFqo5zbmnS0HyGMo0YVu+R+njYfEvJeHVojcXb2xZmP
NYE1XbHEfIk2ytH5G+6VP7pny1pEaxQ9Da32IL3L2ls3DFATKW09dQ+8dmt7Rsmt
nax4eKmjUdpDHIHcm6spp3VkgbXi5MCwIwZ2XeEJV/FfJeSKYh/obim6zQDTyqCB
bQmrOitG7K1utQeSeFNc4fbx1FY+VkSHIHCnT+QwPfliowPAwYRk+exKT+Xv/YCq
F0iPS61vXQtoQc9uR2o/VMhKdOc31lX96IjGFLJG+rqNI91f47zYLtyu7rvDkfbe
TLn14eJtcYFvFDib7J46uY7qcMokB1oNwYTUIkBZaFpkWW1p/8KIFlworQMuFqaL
WYY9JKVm1zYglwja3GsG6CNKMOd0MBjg4RRTTOy8fmaaqvlCI7u6w2RJWlXMRljW
u8wppXpLgQ5Zfy+fUiUi/FBkOhjt+HF0wtginQYbHSdeg5Ji+uu8HsNosTOCFFv9
VJPb9h5Y5YiKHzdxfbMhw8hPwNKsRUEUBNNwmk9utRFAFEcUTxDRL2+8mrETk82I
0cdLl8M4+EXEuFT03jEKmuB/ApxInPfuedeVRP0ro77ogECZSDjYN3k/F7LizTs0
zqF7FTfJA+8H8UTKP2X9V9DFKOFQFATQT3D2dGoaCoSBX6PxQRjiYaYQD/060qjV
DLrVpYdOMPxtYVqToIEMFWvh0hYongPJ54Fz7E09K0BkQkTne2pwc20CsQpmD3pZ
NutTaHC00YXhAMJCfP/DZCI7oDnSkCHOTRyJZtkJsTazVjzRH+XJJILvlCyKpI/i
Z7/wiJqjHyvlgIcZNMroCEEQyM6lgYT7TP6n2gxRVPCO+YeYkR9Zd5BDCR42Kwa1
6xfq5Q3kjlImUuV/lSopPQUOppYiVlJsj6owJYlBnr59gLI1GbMI/r+t4nsPTUvY
4luiE3HyCmF+jDVo75p3La4fssugVlfq3CXYXtw3eMXM6eVRnBSA0bWsyjHHsDNU
zidriKTM366Rj6yH+p/JWX5v7sXKRbcFhX5YwlSQgucy+HlGtB9XU89Sbm7sVOGd
23/1twkpA2hn2+rvVQUamK/W3DsqBKnsAErFs0AN+LwEQEV6+1923otzNeGUZkbK
d0C2Dclyydg/204y6zkShcbsDD0Had7mSd69A565THYLXhESGtQCpIsWup2qlvrw
uUmzPGjbZaCqQwfN6prQtNxEIoILp2HvNp17J/7/GejAjlqsDsgnkgEJX66wFjkL
iCkfi0KUlpj8uqwXqWy/TsjAaUWtBRusdo3HWjsnUsDjOE05f5DBJRCp0vxL1fiU
DutmDgsXvPAjOtkNKUIyUrvLSTSLZOYzQ70mD64M+eqRPc6tARxT3IjgtGoBV+jc
vlDjmXBSjykcK4Qaj5qUoxBMPtcXwzQ52rN9gJuAU1tIUWmyrHNFpm1+zFpcLHkV
FDLAHjmNW3O8y6Tk7i/LPhFjuKnPrVfsDf9qi/HldS9ErT1HOgbZaWqQNInvPzBt
CC/Zw8fOKGBQquvOFzYFMb0qEkHgheIOONfEwCq0W4tktIO+y51eq4Nm323jxGp3
lH6GJJtffm8sUqj4DwtkgNYIA9hbIVb113L7GuvnsAoiPF1VIqYOkfGeg84R2mmu
ibGfuxdj3amvXkAND25bUNVB9Anc45Rsl2x6/rnGZN4ilAEtOcYHCUXmKAuG7evP
Lnr12ny2yerayrfl2eumGF7Gok9WXfRfP589JoizQGjgSVTOCSm2BVQFmr0m2ms7
Re7sRIuv/GK+k/Hx7fSeduW8a8Ab8CW+4xucR5VFcOpY16a5u1u4hwy8tlM84+/M
v2ID1NfymVK7hok34Ln8wQb29ytvB+sAWE/+F+adP6qfNWMBLvIdFD+Bq8W5Rppl
Jbu8O64TPqNGLellMdgxsB1yVQ8r87S0uiTe2nLMsDb3lrAe8Bt0ZwOl2TmpHQWV
d43LK9LznHCjtvlOzgUWGHkutGC4LpMQZoZ57P0a6UuR/deF6J+2glNs4aiDyzAK
kCcqcaTXg4L9voomh1fVxe1lGgw+cZal1PGwjDQQ5Y8P8P+MOz/GKOeTcUyAoS47
yy+f5fRfxH+f/8UEmKwXS+13ofZmqn2+TBy+QcjudFpWbSMc9z/jvuRsCKxbpnKX
jhKM5aERIBEJW2TWeYao3dh+31dLQMJOy/+vU2DvhQBkfSuNKd1yX5ZDuf6UUswm
/C+aTmk8r0LDe1ZrtKhDzrlhRHQlCSaVDvW2em0sikshmqW4378MDKLGREWAkaLb
uC0f79q2eUKKBT+zCF9bi20pykZ+eHR9coUAj1QAUsILbRenWkj4HPEXbDFUeCem
8BT3GpBaiakbHknk++Y4abYfnr8m0y2ZQK8nIe5P7YPqww4eHfwOEOywNSfNM232
vYKR3cdMAHcnQf9Fhp2WXyVONN33brBIsNmMUwjtcqF55dBzirX6RDpGa2vDfneW
Cjhj9kmwqVMQXJO0UmL97AqJT7bz2+L/mB7yrc8fEzneNPPQmSVg9E16d6+xVUDt
S1hR6rXdbbJ2OpZuLsAyHAYlJDvpe2J0o9thfZYhW+80l5QTiHapG/kh3KIS9wkr
ZfrhqRdnChUvHrWuNFx78T11ZjO6ang//sFYp9v5oLb8Si6q4n6+gmMYNsyCqKJW
Ei8tVgHmRTywwiWsCXNi8xo0E7Gk9uVnnwD+d5q2wyVDAvtgnyVpv16S9VXT027R
zxCBbZkHTdGi21F8v+IEcYL6k0lWKqeXpAx/f4s4uh23oIiZK6/ZKewe7N/ykl2A
4VhlAyM10Pg1yP8Pcrt3ingVnWbSA0sfoqDQze3qg16YVt4d54zyziUuhk6kO39I
shDfig91kFqsg5LLi9grIOJeGuKaItZMYrHUhT2lgTZto9oB92wSsx5ETkU87ZEU
4trNV2Uvhvu8gc1CcpPmU2TqZq+JIXxMjWZIACn4HFo1q9dMW/QWhOtTmcltCjVr
CIgUV8xD5GghbGnM2pKXIsswrNz9/oRTJpew/Xw6+DAYFDf45C1mTjKnT8UlkMaW
yDgY0RRueAecPRjd7o4aZBbL15Mb8TtUpdyFNKJOp87Po3mDYKfPw4RwtbCNeWzT
cx73mF1VcSbzACvtTrCGK249t0kUbZBGxFGoXadJI7t6aQmgbJVGlyWLAPhzr+Z0
zWD4iwbgOzon5gRCJ3ncDmGzpnAnisvOn1QkKI7Y5FWS/oNBhM+/ySclPLyfGBnx
p2vsQv7MDP4kVJaYihqmuQBqia9KgN4ANm3KmRRjK0wlDN2CqMDnmjq3ohWtYn9I
hRsD/YamzMVKpi54DKRZQPCwNxw5KjIZNYGlLr2B4kjvXJJRSycDwiozLeuHJmkc
D0DaIMFcwGizB/7RQRtm+JTbe9W5n2eZBIl3BYATRLmySFI9tkQCXJGJRx9A59+J
Vdso7JpC6nhYOu30DDluz4AEZbltCerQRQrdV37XKK59cI1kFNjjsIfKhNWgMOr/
cz/v62vpZvEZqAiXwdm03AjOdRlGCssmbge3iNpnNglBYAiUQHHWYTKCKuKY1uT1
mU9fViIteIPpqeBDfJDumbrNDZx6Om+36MjeSj1FE36nudLwkFkDdtQm7TeQTcmU
5ps6swvo6vtyigUkPiuMqEysWYQM/lfGpTcSrj1HX2cy5iXXTp4GJKMzZs1ZlP29
lr7Vs1a8J9yPqPFwYL/wThxHFBZkKGQrNqUrylpy53rG6BknOFhMF3r6ltxO/Tgk
WI1Eu4/THy/qZ46WEf8ZGUuGQmJ14+KGIEsA/yRT98whv1ltmPByxRPsuJwTZP3L
AdZph1Jachhc1QzxrQpOYNhKqn7+vuNHF5qESmIvYY2Zz4Svdzg2H9yLz7tof6Pp
owhaEdADqb+3nhxNwCmGjIJwECE9mvnnisLL8G98xx5ss1i9/uDRjmjVQTuspMfm
CDl2t1VE7Z+4n2JVJuiCVHOS/Arxq4lDGVnJ2yo3uxi81H8ZD4Fox1cz95/izYwJ
KQ9tFszmvJqCEaHmvn8xjOUO3lBmrHxrfDkcR7lo+60SXCwDe3Vzkmv7wBrzhcyI
+9wK5Xnc78w8E11kyo4mSCUWTfef9rU2Q1oGwtajcDItKdNqgLt2MV+nY0fzO0GN
H0TyRauG5N8BgLy5EH/Qgtaxtak66yk5UKB/26P4S1ztJ+2bkMvdeIx9y48KkT4K
Nur8dzc4JK0cegAE8DhTlkMB+xQR2Y2P8ofrLTCHnPQhtJFuioYEzTjPPYq+fEEC
jMMfdGU18W6flHrCSWraRfIjU6/1kUSkj3MK2rAGVxPvEveVJUtYe5c+t0pzTu9x
hlZs7qQHiQ9DUB6d8LQfukM3KucQXbZt14fMY7TIq24u5D0FkTXcLagF8VYTUKj4
N5yuoP7bNxa7Zpy4ARH+r/XCLqQ8NHevzkNTDj9gV1nNjen2pZzPLyBjGIx67deO
YL+GF90yKhNL8zzoEQXhmS1fz3vYDk03C9V1pQ1mYmim/S1Yd0dff+aLUlnMRptc
HDXEJR+CL+29r7kkuSyfjGXH6x6Gr0Ni73HscCC/g3ud4lilIEdG1VTdlVTlvSxP
hm5xRHRNMxbxDfsm8zWr80BDCfgRnMpY2i6JmzuIB1DFByg49PvcxCypr8kLKWmu
KPrB6AdIKBS7YtoJu14S9fCvcJnfe9uKGKOHCMWB5uAoTlxuL/yzG5C5T0JtMErh
gG/9JZfvq+97qrBwaYWBqtl/iUcIaD6QK6TFHiNXGKyK7bYIF1tUjUhbHTJScc+1
lZFV7cc3RCuoZQ7L1A7Q115B4mOm1wigjLax5+4CdGZFL54iQfbnX8T+z4Z8Ddk1
appraJfg3vYaKgiKd5Nv8bLhIbWFEkC3Mj9mbVsAd7ZOXrUwK1gLWdb/ZCHhplfc
UEzTcmqzTHwEc3B0RdHMkC1bX1b+vwbFmCDq6g75Ee8v0C/0ruFXg+7SqywSZKpw
BvnUplgbDTKzVIMIpfYFJC5pk6B0pFQxw//hhS1sOUhUxHF/VS1/aeI0z7RB9YxA
2qlSF6ZKCumOHBUwrhv2h3YkNIRwPQFujrN3JasXXUAdplCFoGe2UwKnzqfVj0M9
nLIsR7OIFPWCt9JP/M5v4EkdaW3SblFRff2FzrEHTDu17MJzjsyKkfWVHemDAwRd
3huR79384aAIRH2DeTHNlGb5WMchwSuYF9Legl2HK7BnegDHan+mXD5O5lVh+Tzv
aAGct+t/2LSEVMGSu582VPdlNfVD2OyjIivs7z/UmCX44hzXwg7vh/SPnRf2JzYP
Wx84EcYFqiTmYwEyUtTS8MrZCvKR2InfrKP6yUwTn+tY4W59XMgwLQ2i66fFj5xX
JOrmgXU+1uKZ9sV+QoQqDWB9/B0BzfXDZkpeefnYmGd3v9fdlRM3JBv/twlAso54
cvsddG2apOFhJ5zhtfxhrx3DsGFhD1JvNH7GRSS+RTimnqFvTNbLAtqxauBlQSbi
e0HWVZD/b7mYNUX7iyl+eeMCuEM1sWJqvtxburrogPce3u3pX0TN35htex9YiG4p
8PiwJZJwC5LFT4ZPGNRG66+KiMh+iDaBcOFHHxHN7v4eEXd+hcMn4a26zGlA8KBn
r928aWUHdWx874rVWd45vOHgG5wAWCcolOdIge3qpxOrA0tQaz3SEtQmCA7V6Yx0
Vcz9GmpvF6OXW+VmaCsswLZwKzSG4SF9p8feZSOPWKRPG48546w2Y3VQ+k9PAEJm
2SMsS6J5//yfkG12xLiuubtgXXvxDjiYR0/vjEJ65KZd89DNe0EhDTf9qIfA7PB5
GyFkNmadT3xBDX20WLJ24FjwZkFkH+a6nc/ty08pHUXCvF9L2TPPCV6c9j3PSiZn
lq5jsJxyn4b7W/5jOtNSmHd75YkmfYFzXHxamIBu0mJvhwMBq+SuR1LMuM0ygfga
YZabMZxJ78G3E7VPanyxVU/PNhwxvmzzEQqMlgnanrOuQkEXtm85k/GvIBp28z+2
3rHjAf7DBXCzadkZQQaLbK+aAEoVsdtC3I67q+YQuartssjGV+GC96mCXDgkzspt
9LrA0f/Pl3km5Rc7mzJ83dfsaCzXKlUMaxHX9kSDx9FVuFmh7woylrM15C8x24DH
6NIBobAl3fxN6EUadyDpuD2LgmyT5yUUPytlhsIx0itFY91skrRDPxx/5sYJmVVX
V5YsFZqZ+PCGa1yJr47sDfkQWdd7l7nQyaz5N+VfYP11wYXDSCySX6s0GFt02s6X
mJ9moiUzOleqcJkf2DwcePQRiotKXwyC3JdxlMG+xyPIInFoP7uyG1YDhlGRyl4o
GEOT3vFbxFw/hcH/DrFvyuK3xGu1oZoPIP/d2T58V9Dga1GXx6jlP9U6/oNzIWA7
7m0NZEAAoOnBGziRpD/biroB+8KbMC/PD1OUiGlPmqu8X4hXcom+h5+m+0INrqyD
kfvlF13hct5WEM+4FRZS3OLvxmRlOhchrGtjqkYqSzNkSqqt3pBsA2cQJNHP0932
lb2hNqGAwGvaEXQzMSK2fQ10Dld2dFVBRSIZYwwL5p7FLtjUOMU2AwaJ3UrvT3jU
lfQwtsCJamTjVnNU7ZOL8W/CTYQcCMuMBZ1ppPYK6XBUlWZL9sVlONHuUbwZc7bT
TkHg5hQBklsItASH/lpBSdQuhA3k/WCWRuXGIURk+7N3cutlY2dTg1LsUFNUuME1
Hw1h+6+HTFkiRbXEJJrTNN7TKXdxudmBJzdp5zgYrsXWbVKUgr5rVMkdZUpyoRq+
y/kVz1IOSpr1jygdIrTktFnF2N8GqoFJbNMZ8374fDK6OS/fY73BvZBlO2JgeYlw
QX5UxOZxufzkINccVQkZWE59lI6Gy76rA8CsyNzwusDxoe5iJXjZcV89rREKDCNX
rXe3ZMGHVIM5RTwiPA/TX3hFctUJ7Av4jDx7z8vzcmOrH9u84OI3tOdwqk17xeDi
VZbvcmX5CqjxpDQaMxW+fnzPH737oQdD0lv5IMKC2BJCpFhliYeyiFMx2J1oP7c7
dX/JeX8DgagdHT+zGZwijab3cvQpigkWcBPL5aqNSXh1z68vkPGf6Hcn73pl+/en
WMB4YzVRnie7HJ0FmszkpjY1xmlRZb8gX6ZoB8Bbi5IGa6cEE++z6KVRTV8SFwvU
rGiQUyUF+7+wR7Fnri7NfSkQ+SoLnmkq56SqjgsmAh7aOSmC27POYzPhKHkH6ov5
UTE73k46bpiuFE+x4VaQQ04Cc2yA0gZtc7uYmAbGdYWlWSTnnP8i+yfr4dFJJ8J1
ImrDmFb75VbLU2GtfCxsj9cgg9I5vJOHH/ILqBGFfqaKevfH50aRYAlzqdu2/Pfh
2lNwlrUG1n3xikved5P/46sMVklWqSS650e8DI5ByXd7uY73t/ovZdULWXeZzfBV
JlzEmo4LqbVqspl6MjwwPfrW3XyouND0LP0O93pCNONkr76z2ALvgrbE1uj0XTNf
FcccbJvi2PE0XYDOBadJlMr0HWTwVYl0qLv2+jS+aAtfGYGWlzXsB2jOIZH7o5y5
X7jm5HaUwwPtXqyOeI2vc0EcuPPebnm95ZGh/lGGAkCt9bv/3BWcI/sQk40ObUmq
L8NcRyKbtYc7VU3Vp2Cj3jg/31lajGQ+rWxot2pJ+YVpS4G84TYJFcY1orjWUiJX
J1cz9WKfYRPiDZ/ir2GiVvBHFdd/7PcU7EbvnCGUlzREMHbdzIDfqR615hYwlV4L
4pmb6Dhdv9oD61jnTbivwoxUVYooJjmTZvVVNjDcAWNGscoR6cIAXAb4MN2TnyPd
ej9gxhlMokCXL3meGg8pm3OMeJiyrqDDmP9nriGaFJoIi+dUFxdnJ7pekKQdT6Eb
tm76rtbq//K+GM3zRs9Fr+X6acs97LOw50hwu1qJnXWZoQ7ZUv1wMoz+2RDxQ/EB
vNTIJmfqzO6uu6tqsHhQneMsxIhAxudElJ1g8z3Vs+I+R8qkwGA14H865Zfa6jBI
fkfKSg3DFSR/18KONOD3jWb9FHK0uI4Wy4Ts67+wgxX8EG29ZkasAo2/kfunmH1I
St2ivMds9FfMNXQD5fC+9sknwAQWZpOhcO/nqD5GhWm1D/cCsK7ANcvU+uSVPP1H
amqEk89ATOebLSumxYTeN2SDcCovRy6FnnX3oDrWRrFvmuTQtxDLO/sDmKlkbGnt
m8kmzbmra6o+o/iUJUE4HxlK/m072veSeb3HVGfjOBCzdf/YlCfbebDreVM7bebh
3blCHEmkmEkOErRgzy8NLhA7FCOc3f3+UBY4GFl/QYhBYIAFhwrQg4MPRuOiYl7Y
PP+jUcxPzbryMETsoDRbsM9UjGWhEBiNGdJFy1O8bKnHhAQ4K8X9Uh0tbKV8emRx
6xJdkXwInxjFxLP1+z86YiFcBnErvmqdnTyztpx0Ot3POxa5FK+hdExgD4bPHe7z
QDam0QLYrHGlTVdm0D+6ov+zmv/IzmnhbyVGkSIx7Y9Wn9RBzg7jS21Xkqz+AzXY
IoaBsZp8VEFF235Eb+4U/vKgB5fOblzvVYJLj6jpQjsDCiGa1XOIzZ/Zu5c5+qvG
9Kj79523Hv44QxkwK8QBBgeH1Z4/9PnentNvNILNp8PrcO4Gpj9yk7NwFemA3ZaP
5kX6mx80O5zmVZl2C2bX32gnjP7zL/S92ktolLN+ckBegamqkNKMHspmPHwjdOSh
QP7I1fRkk9zAJtnpxCHNeVGd+ELMpBcGktFpDjSOudpBnDWOpTvbYvAdXzw6Jybi
pUxEXCFH0IBIPWtCO112qnElLAI9p94nGoYVdNDead0kiT/6cGBusASRFEEHlhON
kIK97V9fuZC+N8bhSEFBfx1qZEEJZjPhze88gPP043tPtQuNx7e8Gvi+1Fdef5eg
Z/udGSq5QtMBEXbbUhvrH5Vod0FUWCRudoP3hss2TsbANgs6g8Bi566Q8nvrGTS5
5/KqDA9DclJJTUxVrFjjoF1JY6AKAldjBUehjUk0IaJyiohBWUo+z0Zc55LzRZZC
xJjWD4PghbuA2Xp2Iha+p25tumw2VEQUqKMU+01AD0xG0BmOH5qkseMpnvRvnkiT
gQYYJ9wvXCWE+grW188c3ZsJid0GU6bRLAewVhsR6WxxaG0pOS2Fx+AYA+IcbJ/F
9W4Jojd9ucA0WHcrSV7i0sE2XzGvb0PrxpvgXBDMu64FFV8I7DqYSQ0TX5v1tPMK
hS2KTIkSs3B0crMyeNLoTB0uVNUVRBC7XFl5toNI+QmAMS6E1tLEBVv7iToe1P+v
pPTXKNyOjoQOTVbTXOf9XySp4T74phcX2tlWPKuV13WI/WNcmouXzi8TRN7fOL/5
GbBI+NZoo01HXsk7RFgogRYY9nqal9kPGkkgzqebC3Mmqb9Z4b1UbASXXPIJrUPe
0NtJEez2lifKRmhkDb/ta592+ORpgmnQmTzCc5XHUyemD+TmgT7hjnC/WsYOcjKH
pGwDQ7vx/JxrXMYqBQYb85oGhysX+WcMRJayPKXuTKJKq1oYUfm6ayk9v1M9cvwH
s6kCh1GvzwGDztMDjaWVTnzhvB6K9MPdziYDJ1lUbUq9LKmc5JjwdW7/bbOGtgMl
HlmhFUNh7n5CvrxFFTWZi+fgdLBNGj/69XWximoebJFUKA+6Aq9NpzD7tikwgEcs
B7NjbAr4eKzlNr1cOTGigyYQxMYM66EOBr6C9eWGXHiwDwE+JUpAZ3oQUtuzye6/
RfLc+EYILJMp56V3CLfAIJ+Wq314qOO7Pcl57LOL9cqoLGe1fXpTpFiWqmzsWXGw
0oh1dR5Vam7RZ7OXCMnS9r6JX8pO1I8nCV+LjTNXJ4rM/3r2XqeYldHMCm+S9k8X
v4O9rIzLIhnyBNv3w/Gekn+zyHpGFwFSX4nLgrQ2I+ha1ssjl5JJLZTX6qOzxSWV
f8cgpfxv9DE+e6pNUQ5glrXGKsigChzYUsFnslPHkk6FQcPKtkJ7bW/MQisRNdu1
V/A7WLg/AHm8gXVqf+ZUClJWBKZeFN14gMSuTMGbAarVHVrvoKfqV3NU+eU5cwbn
5UbCmZ1Vgd+lAsgNpNLlbNqw1BdVE0VbjddyAjVhNgu/GTMbmQkaRG5zTiLjl4sF
1OTc/Vw3qAosbkHn/6sIujIaUCHoZ0O1vGQmp9bBQN1uqVpPJ3jLIMQdGxBwsrIG
aTAUT9pA7q+6rNPpZSU3l8dveVKcdFf/7iAYCUk2tkKN7x9VM3PwB/iMwMG8vP4/
X89Io8wJjyGEl4d1oJrx+DcDT93NtiACzI0GqIagx+5jS/dCNclfwTEW0glbRioM
GWfRIxgjdr93pEkiwnt0LRhXy7gbD+fHEF39zTsd9C4n7gU8VXH2Hxjod+xNuWu5
kA/YbDV+sKUmqmPEOief8ZiBOuRom7DOweoXtnznpFX6svQ4F6xKs3HLHwMWwwY8
L/DCtR9wS+9ZlUWIRsDZh4YtpQyaN7Uq4C+lD9rBgQ9QQcmO6Bj9aFQJX4VnFv6r
s8Z5rWHGZeVbxKi6v0XAJ9QB0BeZi4GLpOD9t9HoYtuLdQ0//4CQg7z6ekfjEqhj
NKDUv1sJEGrVw2Mygx3bjyCSpGNGWb5iobMLHrVZBYJrV23lZhr3D6/Yc6ogHTNf
OX6TU5pww8pqgkxVWNvpP6GT6vcmMItPTnVmeE8/ieRnaT9+kyw27XuWmXT9pNdO
irc/nulUX9b1je/PggyEPYwEgxbdIR09igzcsT9jYa0dJMvojmL55psEA/tTRjMP
PmhU9E1KMWdrIMSAJfsAJrNd8clqofgBjglmFXrH6Wi6Ra03jwvi/uzh4es/mnhh
NI7cmz1/2qYH06JHcOw+0cvkGuT9XQ/2IaoRINEl+9ravWCinerkaNxlQsv0b/GS
2mHEmYCv88ektW5E8e5XbWXPOdAvoCP/GCMW9+Mf4UqFiiG9Z/LTF0PReBs0Okkb
FJlEgkdfI4KQs6j4eg/mMm3PvE/R3Wj5WuXoBKz0a+Gcx0a41oxq08IP/8Eh/ESp
wMIXFXCU79T8Wsvnk4XbTR4oWwYCdmAsGWBRBoPG4vwtzdtSEzkTUaQ0sir8LGHX
Kn44sSuECxkr+NNNg61nEs3hWJH8I2LoJiVBmMGjEV5ANMHimQhVASdjbk9MuVwK
uZBz15gia9Ajrx4xRF3+qkxGgvpddFvQMVTW1cITSUxSH1oAQtKT/7oLnEI4FUKz
3+6C9GhprLiNTmnyQfKoX3kojmSFaTFCKnd4QaI3YA/dDbyeLHN/UC0nC8k5IX/C
6tvdIk+e7KU5Qhl5EkLz8lc+5nSwKCgpwMZrRrr5TkBof+/bAG2zCNrnXzLx7Gpe
u/w0isRFAeKyXfOC/lOI17nES7h5ar1PL4EL497Sow5BR7DAR8Ir5E1MgTQ1NE/w
u4fzJtf7NmJH2hMoj2OCcrNWtNuG43Ol1LUItftc8rft0TyGbKrMlUuMjfeVNeTx
Ni0YlI2D/BzLjk9KwIRXWMM34Tsidmn+aNMGXa5RVNEe0zBNcOUYaDPnasvAKTCe
MFNWN5wS1Zn7s/71cz7wJWrY/Go1BsywEfDZ6WYKNUYguE+owfJKZgUv+ID9Uo5+
qJX7yXQrI+cuGOr3YsKd9ZqBt+WI6eGv0PkI1usIpgMTOwNoyK/RIdasm3BCnSLt
sSt/Lbc6lkKicUcNk0OsDlSeGA9Kx9rjcUeONQLEiMjFT/gkXu54NEVo8vn/mZBq
Z6PhpUPd2WOx0odEndg/X62UAqXEIPpYZ7kyiau8qtxjXIqmeXS9JhyELYob+Kwp
R5PgGaK9ggbODB4LfucIY7WVWFoOnmLuQJ/UWbGcuRRPXbNBPR+A17Hsh1zXFJeH
FJ5CL6I3TTFIbleQ0wfPHwiasX/gs4BRUjRbb7un7vPq/PuoBOoRNurok4pBmhzl
zK2TPO8nubDl2nZj+qfJA2Vd9REYQSNeLx9+RVSjyG5ZlOhxq+TIwUuJRim97wki
jb8EbTVjNX6MO8i99fxPFHMtgBg4VUGITy7dXQLYyL0FcaOpmtFiKcG2cW1b+75Q
HI+hQtnCMwStWwMTxNjcHXaijG5bEqoUOKLr0ojZ0I0v76Qk6QB44EXn3dkkjYIg
MJjsGGX8WOnmzEdVIcp5oSTzMkLah2tPS1r6floYTNY4udgvU06fSOlZgg6hgrjL
rxf0h+G5YP4JfMtT6j+qqSR/Vr+Jlnkbd7PG9zyplnrc51ovK9bBCCTvVIXwq7tx
s9bB55Da8T5X06/xcStzZnhGUoB0WjjjGHYmhLIRdKGbg3wjCLFUupf8kyoyMrvL
lldTI1/pJsWVBuck+0nVH1zvdlqVIX4emyffWoSRS9hd4w4l4piX2Lt7cPtgmy/9
MkEGNkbZlgC18rlbHPonvpKb/VsPMwizbdh+VmKNLc3oQjeOmq1Rx+7RjAwR5m0j
JIodcm1PyvGNVddc0ApPW0dwsJ1nMn35U8DtIYdTACrhZJqnSRV4cV45IKD+aLMj
/QTDAWlCFfyumff+lo0Z+Nznn9144syETff9a6qaabzcVUKfL2pdY25w+FiriY8G
OwUdWsQnBELJXon5J/P2ZvraS+gUoEYjXPc83wpWccZMh+/ekByRh245ynhS7QHT
wDo3G9T5Hk87M+UGJJf+x6zh0yuJbxYWj2dK4vxf7KRmv/TbYSuE8Ldie1usqLqh
ZmBJ/j2xVFI2TzLhHt+VJnKhkHqPSRkYnkoLxr8ebc837dog+sErIqlHLyfvBBj0
BvkS/BlAUZujO/aNK0RDoaezFNoRfTXRQBHjkzXDmuUpLB6Zpcikr/hU2Ks4McC7
MHdbzDMsGpvfywZOTWjDey1bxC4Zl1HJC1uqPiKLn+ykTeLuAdbM62ynAjJV/pXq
Fx7YoiyTfzRmuLMAqcGfKvE+m9LNltDsHmNNR40PVkwBZ6akgngUn98bUqfO3OMK
CorMJN8gWKJkUFhi0bItJZEbW+QaMol48E53tIj5DOSIWg3oa+bbcVc38uJEdGpD
0/5gcALIO6o3Z/OmUh1OL3FwASPySzOL9oQ4YLxzm+9FeVaR/ZTcp3CdcCenQzbS
atbfXqtMGK+V9yUvIM7CuxxmbLPvJJ4mS87Pg/BK0DHuBEgmpRd/4DrMvzul9SZ5
698cO7CAtQ7Mv/FYY7r5CdhIyB3Rv+nrCTWuv+3VsyUaUrQMenWMtWR1hQGvtXq+
TI8X68YRdMWIvj3LEGYCgFFUMKOPJq6NsvDQKrTGN/PvxYLFZoy/0G0AOrtoOMYE
k+WUXd1Cc9860ltEqC9UD5RFvC/CVzOZKaaTIVzALwBeE0kkPRmkgrN0K0u1EdtA
822aVrlD8Jrwc+944ZqdM+EG/NJETXMfqPvyX9995PoL93/avovcz9j7IQ5E6NZr
q/6NuQjAZlgXfLQZSMQUoxFYEEEJtf1TV8ibFoWbAsHHkWHuoyCUQkdv68n8msRL
GWR7BtHxqb7CA1JYWBu7q6VkFakcd97HDaIKeaE84LccbzJrcUpSN/KYjFAZ6/1k
ekYYakNpcKDUUMa69zhnYwGNWZHNs8acHRsVWO5C+lynhPO13cHSUqI7LxVFDnrl
EYOLdkD2S6YM/yNjvt/v7dlnryUAwB98aSWiyYOCRPpUKHPvDxsfbY+mFPVyc4Op
oso9uddOR3Z9ibq36nppnasqgSI780BWj2zRiS6n9Hp0+dByaYU0+0Y6zaLhp6DW
uCJ0OgdjDDQzszL1cxXBmEbAuPWb6WVa43kgGkq1CZwLUxj4sLGb8CUshrK2t1RX
E3OdgqQm/vbRFEslTGmtRvUnZJR3NPHo2+JvRBKmEx5q/azAHNCdva/DZ5Ak3mpQ
xo4+O/NdWi1S6rrSwAO9S3mHa7v5Np/OoOC65/Swsk1dlm/eMQpAHIbH0KcxqWFu
LK7vGjXg1k3Cb21VAiuMZZCzDszc5Lr6sQAaPzkUDmVlEiTgdOU8M8Hya3YUmQZk
9Q3QW5qaRqifyJLjo1aDJ7wpTflQaNwVlSKvo2Wv1ZzalXNS+TLFT5lu2ggbBbi9
kFWqsXegJrbbmrhr+6q49IBftUq4Bc3S2Z7YBwnOaWoT7s54rHYoFUFX7HTLqDpM
wpEHnjjAoxHD2Ct/oHOTBVwlEbOy9Ti9PnVky7IacDS7w2UsUyHDFCCy/ctSr6p+
ks/2UDYJbpviVdKN3MGZM8o93H259VvWXl1exqJV4fTsq29sPop85aAJGV95D4QS
HFsYldDcQ1LNxlurgCIipTBXaGIpzaHyPprxwTR/4bAWsylGDeQUCvRfY3L8ILnI
zBu8mzMOJTevGV16IzHXbR4Pi2WnMqPHPDOu+jND27JYtlZ2X3E/fOghe/lMBQAW
pF5fSUScpQM0z53dfidaBHaRRO/gt047c8MaoVzdsUZwpg5H1ORaYlqxjCbWtfb8
NstbzdhsK1JwhH5cx/hXq2L9i4NCZCTOaYZZJSYRrDx9vxdFQnCt8W9/l0VBP94j
2993G7aEl4pAc5LHAkzcqzD+ixyZDzWQPcnrhfHMBHk6OkRN3Gxnjoso7rpoEAVv
XgBFF+s0ytZQuiDBrzz3FBQaVBmmTg774AmmZOYGL3uDzBhq8Acii6XeTxXBQJej
uiojm/GOcp3klEzJP6DL90uchfWQin5QH1z4slRy5VGTH62LvBuu4BAA0uGBQeQ1
BqipkVyGumqd5byp01I3kwLLxTf37xJtMostaF1XFaKA3lnPMnn6cpFrSE2ECvdd
SNzcqmBj0wYVK7nn9u4fqt9qinvJICoW9iaBKgNxD8vv4Uj7zMWJbDcyCK0xXoGw
r9z7CC+ZnHFOSRkL7FQ9JqcT1rNwnS0xHM7Id5uNu+7ruKDdhGlNbDsSzeBnGSDf
vYGWBqFcF+/BBiDbHK2oRHF0dSLZNOH0AUJuWQyYibPKmJiaNAz1SWEpVghf8ytS
4CKPv41RwQZ0slm5I3AelKDaCgJNeUsSqNqDnZqFHZEiPpRrNPM1a7BXUEryGEd6
bqnrqR/huZkquVZdTWtW+hVTJwTMMkrDYQMntdEESvutKspI3beDKSh6XFZW+5zj
nLalM8mlyFCM3z3HzlM0NT5MUBFhNHI6PWeVfIfZZYsw5S44uhSiQymWPH0FxdXo
f6mRXMRXV4rJ+MR545EgiJTnxKGOWf8sfDJSulezOUKFxy1WopINpzULwCst1no3
7ZrByWfNmWGjN9Kwbopbtpq8OzvTsB7J/vqZkT3ZXHyZCfp/VsjvchyZRU3nTQZP
nw8SvQSx0MRjW1N35CvI9t3z2FWOUbKUPV/1Lufd3OyYSf+dUH4sTmP/oz2Wwv0j
iZc1xZL0Z14w+M4bCwjnK24DlurlAWVuDD28Zv0HDDKqtSb3PzdI9gogfM2IpAM3
/Lhju/zySs7g9mRo0+T//YqqiboEy3WjlsmqjjcdRhQYC8fwGc4go59X9Y+zT1o9
K4HRMJsW5Yb98u+9S0jfr2W9J4mduN/JEnDoSip8cXRmjMw4xuwVlWmAtzMayltW
E8bbBVD0kh5z5UYLCy/jrUhl4/7auwZGeWKd950pWAlrVUqzLYcU9ffRDWOcZ30Z
K+Ty7dnd3L01V7tk2GnYfOKJipCeKXFoobWvvWOs60yT9v1Gorgrqm1V+VSQ6KL1
XP3j2154toywGnKhlObF/yVVMQT3LVAj6DiAnFyPy94d11V6O9uY+XWQQbcYespn
3FFV7NH/L8T7hjQtkl5pel+GZgFyHWOxABxB0is+e2646b7Xb0d/ZLCC2LbB1tXy
EDwr8UUqq2DBHLg4GSIoHxmjGJs3gqPgPo35BXY+DDP+CTrTmYSZP7G88RuLSGD7
ky29K3nyLoUBh2hZc/rHCULhnM/TtVbnG0pDWYfT+ps/8Jdoo0OiQW3TJa7lzuEV
4/d6VMMBBarMizFT80mLfmM6znbwfTRgZOyLjZ+urlswXBzuvu6i6pK5LZf8GmZW
dj+2bQN+eujPMO7iybIMoyps5MjBXZCB1SA/tmUEa0CRJ2aVOjp2fr9kDLrzoArC
u9F7KmkeUan2eBOWtNpDFpye9HnP4hhLjsJ0LDOZNTfhLzDkitfhe+MDixKN0jGo
TMXnSWq9LxDeTteD198x706EUlpTqo1RYxgvSOSXmZHVNtp64TMtXxArQ0vCjGU3
AhTrRTMOCYm1ggVHLS6nnKZgXa1U5CTyvxlO9tVhxNsyufKmku8p3KY/zMfrC0zr
5H4v4LIkuZOfehGYpAKM8isqm3snCymiThcoZ9rttqTztB16lXbFAOpbWj4HIuOv
w8mAbcxB2u0NCGr5P7UKE5Z8DhrYe10He8Exqnb3o34++xDzLs47bsuManm2sK4P
/HWTiSEAc5SU14JY+tn/rWh7OljnKxCmZ6t73Nyas1Xa5I1BL/TkUT46BraDAcrZ
CjRxuHE3wfdEdfPPoCvciZDxqzr6BWeaKmUm7BrRx5Js7hq3puWPNHMOPG4ikkCz
PDf2xL3CPsdFuTVM5vmG0lew4WtTvYkMKX6hNBjDwT+qOVGyp5dJ/AfeR4BSiSgM
L1G+wS4gDEXjNksqXvni5Q1VMPZzJ5mfq/QNL1yrkS3BH8mzKmpx1RR5jAITCOjE
Llyd1CzH0e5f+bwKdaaHEZaSlAJoAuPQCdodrCcCPoRy5Nvug8vRpymIMJCc4X7W
JaJa0P0Frotzv3y41Q4xs7azUgS7nuEbM7Mo+6RWiS0BKg+finj9VGuTRutWXqkg
4RabhI0vdNguYzCjF4AyDo3lbJtI0OZJ/acqfvcvB7hoGcm96sapaY2xcOJ9WUBi
nlZxappQleJlKBpz3SjRNgE6wuh+RCH2mbrGUW7oClKVFl1BzZo/PqWI00AYlUtD
fpM+vCOByyKYOzFEvaBk7ZVx7WAB9yjPVi1mZD6rQLbPhpb0hP7e1L8ozRkF0/CP
XMfauZ6s9NNY/8LIfBsZJp+EFlzxpHG6zo//4di4iuWddeKvf1GNar1wuAeRYz0a
nnOE0CkWP0lmC5bDbKoHCx+LoaR1ARpUDN7uF2QMrLmyTblHa7f7EjYCTdqi+5Xa
MUTNBU9eMIruDYbqDiICjq8te1a6cRvR5Tdl8NxvFpEQTkH3U3LRtXzhpkAZbT4F
eu3Xqy3Qj6TIQ2vX9R0EmywKzzRKkkh8JvqRARdtg2hHdxKv9X7B4aRMuVF9pU5h
rvZ/1XX+pjyySa4uBcTAmLgVYJe1DyTPeIm0fDK9sr4M1u7JLTtvnexmS627l6eS
HmzfZ6zpboRVutuQ8YMFHkHFup/jnsYBPPHbep978HodFVzxfwaOFe8VccgD4YNg
3rmMb81o8Uw+Qtd/04jKiQ7wFTtIkShRM4tiRBGuONqro8nJISNEaj445eYZ2SYK
UWenBBSJaQR9hqhPHvQXj17nU/qFPuoRR3ITlwnv/9/sQdoN2ICtv1G5wHMUSF2X
5Bx4+nOop5taXp0iehkcPATAyteRED1UXaOporNAcud7cpZ/omFL7ZzMLxlvA6pE
Mgr390isWYhCk5uO9Ga1umCEdj7uIO+Q+kt4jzVsvnsQB9pvAlTkNpDMr3ffMSux
8sVpBIPqjHj65M0gv/nINsr2mUGFWoLZFFvEdOwScHXqYTmG0jYTFysRTj2QysI5
LbRoBNkJuGPyq6KQtIC6rQN8XY5pdvFngm9i9HI9wzcdX7UbATrwFv7Ms6/iYcSK
wdJyAz+snGF5VXHbylqvCDx5tTWvrOTkQjFZDYOdFH/ZV418iBkNWS6X2DWRefhu
g8K5Hbmy3R15vZANugJeAYBhEhwwjPobBFD/Du4TPkBe7baij2Ni5CDvnNA/YA7k
i+vQ2M2Km8X3PfNxPC9ieFEhB3yLNFRhaVRUWyBljRzN4+efXKR2BxxvuasST8BP
zQxrcy5u9YPfkQMtFljJbpad6pLTrJt/yZI38dW5MBNc+gD0fKhduLMdzGBq/6/9
tarbP5+ae3WHUHYjBBIen5U0CjJTTNamNU11LpM5oY26IvHaooglVKcEizNAeltx
ykSZOKM/MWkvjPYdNitJuA12ij5s8MpXNniQN/P/TT9sKhuImRNacSk3sRgyLyfW
s4aDCYR65jMO6kgzLTL0EOMtzuNOLXn6as4aZk5/0HiYvL/okci0npPoPiUVeRjD
r4ljhYqFTzo9dG7fdU5TFePXHWDdiKnXhAC3upqZASqIb0K1QCXzAgeqpVDGIwPN
zYPq1Y2A5UXIjSBENhQUrcLDcIyjAQ4XQn/hABUpxaJlAeGC9izRjSX6pH+A1nnG
KSOTgm03qebmhr+vzpj91uh6bxMleyKLsHrPbWIPYqeJmoOqVCBeFUHP07cSWSBR
pGdCO6r8pk7Ai8CD1Zse92wDa7yj2LTOi8a1eo3ZZwOa8QEGW2b8ROG0XntK5Wbt
6mYT8hAWH8d5TjRUhp1pmrM26DTXcWUsOiN1srCUw7pvgC/JtQsqE+j4y3mbe2mo
kCjIz1zcSmvR/HF8osNA45kfrwl+m5RYCJp2lzjc/dnNmOdchO1QMyKNznmgHgXJ
s83edb0JCh3E5M3TgWT51NONFjhjWQlnYTimqjHRIxKB+VkTb1ByC4fnxrsju8s8
sBUMNr2/WpV5FDAoJYHEStAzrVeyip+lnNOlL07yqle1anmnhzmA4tPJkCVa89If
Oz98vKOBOahL11RAX6R6ItrpPYqG5UF5q0ISqD2niQyZoTxBuV6dc+tmyeJozi1U
kVVrSXsapM4CT0X7+APx1O0UwUlIF5izpUBi5Q+0iiLmcX5ylfSDlkxE6Flgi3kG
4S1vLNTYZCpPM1c98WXfzmcq1QzcS7Ozm+CG8rhCjzosqIEjbOMKQ6LPDEAsOsLQ
ueHRNIKCAVlGxatZ4kqgQ/Xhf6yJ/MyL4lV5sw0xn1+8Px8sTDozO2w9aa2oV/X7
/jYw66vkHD12G760E4+w1PnpsO5qT2n+Mk5+p5e/N/vpNYxZ174/q7T7znQZlaKy
xOK30fAwlE+Jkv5OK2STeqjKcCpvfPQuP33XVG1uaQixyOfF4pCXXlJvSozyJsiq
MDaiq4lwznnxinnvdF5jdxeyvSSSW6p41newYbU/s0Sh8BJjYJLPUqWhXyEDqnZK
5KXurG5vRIkVU+Lqx8a3f1bSU7C+0YgRegKOInXcQ0kQNO7A1b+oWDwKUdnVg1z1
1tJCbFmN5ZQOX4zhyIsFygU/iyqF/y0Eei0t8So8dUcW1wG/7P7gQ6Q1swZOCX9F
NG5ESwYNYU6R5LTZ/3WjpmxDMJo6XhxnWVVdUsnzbPXNekac2JEcNjW5HLlPXnx1
CQQjoMX6qApGLZaNNWfDeG3LdvT7ewVe6YNybaYZpx1tkYLEKKAk2anLSWbOSjpa
zLv505IDkCaaAw5uX+8uWsI7XOx8uFWjkO8/JMBRqKNCa5oaCCOuhVUXHO7M87cw
PsQ39CfgAtIbgrJn3fpIc5q4hiwOoOnl3Di9rhuu6qOug8cpdCirEoN2DcdBJ87z
JfiVpmTq9x42NHShl6ZOnaxPubtp4lWzF95xDyJGsJfx1+4z3lSvHND2CZBM38Ah
1fHQQ/C7LcQDrNEfnn5/tXcJwX0q3t/a237OOKaUzoFivNW3XXnqfrrNzlr0WV2K
ePpLW3YaTjGjZer5qDB5+cKHlJtgi189w8Vs7ITasjjuXfkGQ3FjH96Ng0Y2Aw07
n+lE+8pLLVZhxqnHMfn30eEqVF7g65fQKpxZYPOEEcaUiaIbVK5P3Oq1fOGAIJmn
rbXOdBzMG3vkjnm+cvULvlIZKjSrNwgk6zYXGwev2qhKy2gtuw84bvl1kOiroSZI
gRx2U3oRX94CqY0EPZNKICSmj6iOOZWill/NWWM8aPC5u3plcBoDIV7Jqi53U7fM
wU+z6D6AVJg6IeE2w0b8lC+m8iN7n4lIDefY8pwPtZJVACfFt1Nvz7PEPzaxc6yI
XcjZNADUNGjwgVJ8IiB5sYiiZTRDIZ5D6H97ou5Iwb2gPPPqSb82yJOJnFsp11I+
MVsspnM1brXBlgQHeKdTOuhsxcDiTlzg4Ac02+u+BLdP3jiwnvklTn0BsYpP8qsk
dddiVoVcS0GeUXbnrpC/D0AO1wzQr/Xy4EyNqs1eMfhXiodLitHI6/USAQWkrPdn
86JT83rri7zSZYiLh8EtYCNwE944gxV9uoGeVqcZ0jzIKCULWf8Q9y3Yq237SbJ/
mdu9SMBWjtmw9VVYUKmU9skP+uHbf1TWnWnzuHg4kMTTAa7SEoUeiqAp35MGSOHM
lJbhdkyZ83AVO/RRb6fSVohmHxZNgU9+wQiL8QCLWqUiI6Rw576Fm/7MejTvlAqI
ioDjSW4XRLgg3V1dDd7gi9X3nSpBYohK0dMjSeuU4h7VBzRc0N/yjQA7sFCFM8Qt
ictB0QONKVY/gzhd2wPVaKqTWKBM1LUGCwXk4NMwWkGNfdHM8KBArgt9p9S1eesO
IK8tihLwZrTRjlFCNj67fIaZAXmtskXVcODMWt1HvzhIomRIJgGEjbNcaMjV3d2h
0LcNDfjpm0eJcuVQfFmT05PvC/9wDjWKW9aHW/ZryHLaPLFLFRjFWNX+Q78sWjPb
hkVUR2NTVk9pOJiVictn+dhuUOcQeqAFaCDfLaAmjUB3IpD1jXm7pYk5li8eBGLg
byCv2OQdzYCTNCc4TEH2WWS+M8f1PBw/deec8CNfLIpTY64FEWbFwLu4/z1WnaH0
xsOdz79FiTNNCn94hEgdsMYI2IukSezC9rFKPcYnFZsYnUtyLLcIbc22I1JWSpU5
2GO1RAuIxKCDSb71AEu6BNgjv4oGEJmvz/8aClI+8EUwTD+mvOodKg8IqcxiCTaY
GgEumpG+l020oqxAOfhM21YugM0yWllG8sz5IgjB9ggwI3UsUByPZjODQHoL/Ow5
gxqyJALPusdcGqpB1jyZtAKGopKvOioz0bkG2F6nQWXDWwi6/bBJPIerD6jgp8sC
BvMPfYuCCxk3qMabBu7NrXBFh4qMdUb7XP/mjDgLR8sd879Aerq22eitwXXf46LJ
IIaIU+Z/RGRxh4Vpy483C5h/qNpk5Kc+jpMvs9h3C173FDvdUfIkvRWOU6T5VIAv
ukjthr/eEWMxw+QaeKWsUlusakOMubl1unxQ3WybCezZ9+8FdFIHqZcP8OYJHzvg
GxUoiHbpsjntEOsm3kCvnn7H2OxZmAmU1MfQ3aIO090HQHTNM2jVEF3nmDZs8u6L
9N3GV8y46A2A/WpAR9RXer+Qk1iETIB5nd5z95NqspoCRD+eTt662ZzfPYvxmV4u
k6HHe0PhtPY/t3PAporyPmjXHTfvYOQ8WuumI6yYefr/N+1dnWSxTQ706pQIj9hU
2Ra1NE6WU/XTcVF93uqzWM6vLYG8pMt8o6RDJxL/BuTS7LoY6lrkLoSjObtrFS+z
4c1YGIhW12dHIoY7ZbkRzW49VU+a/okrz1QRCGoqKVoZK/gsmFeehUvxeMkk0BQT
Y3T446jyR9U19ZC/IhVGOunHtCTyZKbDPQ3ZAPZx/LnTlOkis1RDpPYiFY6MCGJU
Ww7Yp2QA5eCautSGNC+t2g0UZkRE/Khztzsl8PrLKJ7PeSwQ89vfpWvfaMA+tTb1
UkCZlT1yKXw7LVzegbHWCxCXI4ehN+27MoIox8vtAhJZSadzIENOhMphAOO41iMl
iDY3Ji/hjruQJoNf7sH+GigXJ1tte70TTCoOP0l+jzNhz9gZJ4TNYC8wzkGGV6Xy
lgS8KNP9uFWVQ9buXuOgkwc+3IHzzloXklfW8+PypCaqKNs72bclm0Pi8Ngnittp
EnA5xmq/m1AKnz18flAV+wy2TfqTKz4iQ/zHmKecCXJaUomh/VG8Dm7b97IA0nxf
brN8mPLtrTPVfzKnqeOAuFRDNm+IcH+q9LyYNmrZDi5p2kZLmrCq0wnRR3/8fOqV
27AZGEh5qCaeQUfJtO42eFuSWwL/1RA9i34yCrA0l8EWXas0meUbwvt5XldjRh3a
TSVTd6NKDnywaZkKxdIHJRmUYQOaGx7pc9UqC2pzc3bxAJTi7/gpkK+4f/mMcuIj
85eM+Ehdt40vTOZVpvpMsViF1q5Q28vYFjqfnG7uLdfXMHlP+XhCZ3WpNY5jXc/G
jdaH+1oC+HQRqS0hMQKaQAWIXdcSYIMR8YvarSmMt38H3xgWbATAzGprfzXEyy+S
JZt6ucYmSRlm2/AwHrA59BKnN1RIdHjT20atPg8IhIPVoBlVJYiW0gxcdcsNWdYr
9YwgcqKCt6nXQeAjFVzy3lxnNtQfoi6GQ0pcYilUy9eHwV16vE8TeiIi3thQ3Hfr
XzUT7iyFcvikrXgwYAmmrp5tGfEVc60Z/jJiJ/BeZok9ZnONjlZFu355/qTjnhlZ
YypQ3AwabrKIOlRxvv846h959r2gMnuWA7l+EEsYVBeje6klqf6NikmxEOj6gFz1
twXDFWshS+LEU6jxtjnhZg3axpSiBx7jyZConOBc+tznWIZNjS+FBa4mGVezikoP
kZgfRSdmTdK9W20Un/wHnuQju82Hgow/+U3LGZp7/odQhqPNF3Ot3KZ4TO0cyn26
+5ukqc2va6mz/UJOmr5W9bV1Igl8ICw+cNdHMoxPt7jDbAhXQAbH26uPDyIoQB9l
3sfRDzMoFMvtVbC6PBcA1Fw8X+HBZTZKwsOiu230TZGedEE6zmUYzZQ+md6xOVVy
koH5pQ7lSM/LacfjhLFfB9E3HupFFCHd1nMvx2tJO5orEYN+wEEsBM+vpvuRvfz3
Lw17eOeovwCxYz4S+RAsGBLd01GmNb1GuRpyWHLSCj/3OoLlybzPmefDKDds/x8L
zJS+e0e9Kq3q8Ch0Rpk6wbY4AUHCQzGtO7JzxdISn240l9VOEuyOMsK9euCL69ok
3ovUiNBLgwmIzoRLxJgNblhfcQJIn7aMcEAldX3TSqzdI3B2mnQvXPt+1tbdlKaH
xfgP+viDVokKkcaE0AKSBiaLimCPtjnJ01RNXZJAAlFMZvfp45UQhQt0RTIf4S4U
wt1H5T+WAg+mHcOhP+it5igSCUWDQNIGF5MB9snRCHeaWF4CgKRLOf/wTLcBysw5
45H1+IZE+u1EcyOohjBqv7jqfXCWi47MvjkMh9Xz1nuIc1+O5Rw5CdpyuRyTEXS/
GlfM6nIRWGiHMSn9jEfoQT8RSq0TowtBwkJibh8P4j65Z6O1zwHDKM/KLhTlunZ3
TRfgf19Xfs/F5AMNlnjgmIEHxY4IxJZmD9jTfNHvlWfdIu3GJ6Qqo0c/IZ7irICj
4OZKDD/+WIad2Aho2sSzsXJk3LcO8vnsPmd6gRmKmA8qwKndXUus0pDKcrbqFLkW
lczsvSzw1kSLTvHER+Wvj4zeT5cHzz4lfT8nDvQiX4NqChxUGp4REz6FlggqC7Z0
g1kQ7Uc75RIGv/c1wnIF2nTSkCB3FhmV9J+a3YUmsmZaINbqodd3K2WGuVLlfZhl
YT8VWTsWT8BtXE5UWbgTu4xhA8XFr4jSeQtQmVxNqCMYwdis60PDb6DzjvEpSopi
FOlLjP4C13uRMO4d5boI829WMLgMaPx5rr+8kM04d+t0BLuVxFmbt1tO4h83AnaG
fTKncUyl64vcCs8s1KdBFzajOPDZs+Dt6fuWh/qKsT41H2ptQjVaFsZ9RrnhIU8K
uCp6eFpOx7BH3Jq2HAUkdC/0zdU6kx/XhR0L6CyxiNSQajcA8uSExwsxJ0iW22qc
Kh7yk/8g2RXVD6UQyfNkzdJoLgvEc0SuHwPDtxA79sGHpeBt2fWd67Ea6CO06xUo
yE/gkqg9nQioT5EcMwvh7kQNuRwyon1jP/Me9uHctyLUNRZ9ugNF7XVZEI2rmqWA
lpqE/YdT6s2BdTsa/prSKiita8P5QrJjHs1z0WH987l0iFRQ99s8rClIZdIf3GLZ
ns6dVDgG9fNbSYH4CU7jRF9r5Ztb0YpwVCFI2o9Pv8hBwXhOvjw46Rx2NU2y+09c
cEuRTTf+5lV4khBRDzKZEIT8OZ9a6uXZknHrbfujuTR3nxPmaco3QojxgBqup6+Y
7C8X063lJbsqTufDErruuvBAcrDzzQ80XUtZlTe8umAYACSQcS4mPiawho1+Qdem
Pz6XKfDJVJyiXZL1WXSCgAI2izWlZ0bJEuzbbOy+UDD3w3m6EingZGIR3m7Ncq4L
W72TQTUm3HR/EzXVAm6L6f2F617Qt7TDyZUBhqqv3ZjdTygKBAlKvfOVu/I1VucT
BbLMTwbmnazyOAC/cBl5/R4L1SPp6Je6vwEMVV5bMbDxMm5491gQowSkxtZn2+5q
6betxJobKgPH37oUr/gqV7wVHimtop0FAeNNEqe9HXPqqpTmYzxFHS9C6zusBANg
TJDFzqA6BvaTTsoQGzIYD6meceY2QzE7VJfFrkC5aKSBOn++AMzWiQGXJ8klEBdP
OBLtgNpTuFxuexK1NYxgC5zccSHQbCkG+XVIdQFx260RC2PQiIbMMtcrxhkrfrw6
MJUbMaGcUSz3QdgD+4qO7jE8GWpTPltRfGCkOtFP49XaMdxEUxX36GKFfWvNodcM
B4wN9IoffM4TgSkrwIrBtRFsG1i/gvDOho83ywoJCNznrNComc+ltBF7PVlmMM21
kidmC3xqYGJkiDCjuXx9yfkyUT6FQEk30UOSt1n4u7ljZZiOw5m96KOQ4Ib1+U/n
JGyVqW1uFRFSkWgGSgUjOIODm6pRrUQCjgcDggisVbcFUMP5xV/qXfw5VVpxGVnj
nJop0GXKcRcf3dcmh6V4J2f00x0uU8lzqW5BCiOAcgtRWtcNkT6c5R93Pi7oOflm
IxZ2ePX8HJ/6Vy5ekvzxiMknChzRt4eUPRuMSwqfvD+MQBKea2v4w5tk93L1dB90
MwVWcgJeKskTt1JVZDt8ueJoiBSErvmMf6b6X/lU2h9PG45aIuNo8l5Kds6ea6n6
Cb1Bx1dZTYV5U9kmtb8s3PUPnDfchsYdfIK5zBpw9KGSu6Hg4EBo8YEJNJE1wToJ
iVrXxfBACAT9ozrtqiAJJ/wjpvGPLV9N7U7JBxdYnbE0YF0mDmqiLyE0++lV8s6w
P+bkqdWqc6uzrPKWdz1dEL4ZzhXZznDLFnAjGelYAt/1b5IAWETWY+n7l+vMu05B
duo9so+gQ65idNUo4j2+yl4uO+mejvKQ+SSi5C6WK0uYicpst8BlZ4e+Kp4+HuLQ
OzDT3OFdE07RTQWHuzyMVWzNTXiInp+1qtMLEJ7u/f0zx/WcorT2Xti0A4p0SH5k
E7EOhW5Xs6riFGmkKT0ptr1dLG/mKiP+PtVJ5UjzmpgQ8CMvJdhErkBVR34EIG6n
+P1DMlluljFy2+wX9R48K7WwuqmfEdTp/XdrIvolahIcfF6SDVynItvwTGvVB5uD
khBjDMHtam9PECkzrsXJ/g/rJXtlbsign68ZjW04b3Mi6J0f2Q3luicXoatReUpz
tQA5+z5ILQilaMeFWx4QOKm8dmNnZ5pTY2LXo8LMvafhyYP7kkUB5nq5+mf7KIMe
2aXVn8J6nVMI1r+XH7kTk6v6E1AAJdw8YUqrAzZIVT3Wl/XnALZcq1hpPt7UgE7j
u9rJAoVm1lymd8YmWpWafasfjY9hw34Z12+z0Rtjkesji6tRS93dQIR0KSGtjxwM
mLgio7pSWLEPFNdOn7Q+YT0LvZgzCGLaxUvdTsndrTrF8YxWJgHc6Hq84Vi+DsJX
a9DKAVehtnvjg+r2EUpt7tB/SIiKfap/Z3dixdEPhd1OYkx5OG/8nMo3w3M5QPS9
26rhPSKX2YSeOmRiEI6Xc5PG26eCcIN9aLncrIMI0aBiapHYMT7HWR85TL05qO61
aA90PlUy+vU39EcwByIBpRLRQG+Z/rfiBe9UWxyYU6tkhBxvVWafDoVJGRwyNTE9
gV2kpokLoGUoiMvaNH1u856+GIv1qnNdxwzVzbOrB+ezKfKSogNUtRmSPFHP+Lut
q5D15x5cCQMyV6FFXAP8zpVZcnF/xfRNNChodzCRNNrpywTKkLWhB4zn+yDHqja4
6rjIT4J4nb7KVqX2xmWInNWqYXwD0nKTGrscfUKfAWuZevvWRxdceRtCx5RBVmO1
qwzZLGti4PLKpd4uVIzxGk6bjsLFv1mCefAw6hL6y/T+vy170rgNftj6CvrYNUcF
fM2K35zrrhPEkE78hrfssusW+dOfIJxUGVrph7LQILYmFh3+e2qopUjmBgfSS5XM
rBekSTHfDcRrLcan7TGdzRgoexd68YlpBfNvM2u6jq7GgrG/xYrZKpuTRlDVk34t
dnL4Dx/8dv1WkV0aOKIjCNq7hBKFIIyQ+BU3pktWSm6WsJU1WnuPTOsJx2vOZW8j
TMWULhmw9tMPEmH35J/sxH9sGHx+e4S/AyAO9An0y4A+IcSAojauwgtir0Vxpr3v
+VgGKfhiERqGpmUkf1K20D/ZT4LK5yly2Ce+NQujkx5IiPUhu8hnXrCdMpj8uNep
eb65iTTVhD3i8YiqKGU9kZBkxDtqYxwxpRENBYt1NjCxDBxSNgvy0vuBfFYxmxez
OvkH4vz3YaRwkmkmMuMzGRYNQad35NfbeUZymRh5p8AkG/U2db0ua5WZRs+On1F5
MyVJGA4frPODSzAqCQIppqqI0EQ+aZpzMJfZLwZmUfVt6rqDlKpBjgcaqN7RATnQ
nzWKr5GNtJWNYqHKVgf7L5CmoUDLwyL4imeMYTyyPB6q6VlDB77k0/yyI1qYEH1O
wuCt/IbA0qNJ8GfovFPK0oIGPBMFhdk4xaqcaT9H1DDtM+U3DhUnBVpR9LpI/iSt
Mszec0iq14Yp5SqobOY3n/Pay9Ly+q1fgOM1Aac0blFkMSNOWUbdnKAK4lmxhaoN
fpZjADoOdc+LGp1SPs8Tp8TC4WtO6Cywvq0wUC6lg8JozajMk5NgMivIq9c5xQZB
6nL0/ALcXEAoTb1rgqFaVfPVwC+rrcatx8u0deWzFHWVYZs1EVEtT+aJl+ZaaZC3
qvuIEA6abDmmI8uKH6niLO880w0XrPS9YbV3f3HHteWb0xx4+CasOy5rzdL0uFIq
+njbX714AzRGgKTbO/duikDEmvPWJcrNOgi4wncIIRFX667WxgYMQA50pct0ax1g
ZO474kYBe+6iBrTDyMzY2DlRCvJLBtLZcbgBRCKf/hJyI8SJwske2wQUT2fYwXKD
7c/NkPjau4DtPbUNaQ7fVD6tAkq0rfRpB+mRrB9fcl6Vp0UAHRyleZs7WOdWToVb
IMqASDNGfKmfOuaLEANpblZnNNuLYdz2spJSgCyV0LweqNIUirn7FXH47WacEqv3
zFMAmUeokYM/XHreBqQxXlhc6L/hz9v09U2ouOxoXLri8wtIiFNzbAYfeSZ0H9Q3
CD0hOBB+xvRfhH0lOVL/6o9UIpj0/G21PrSgIYcowgelW79BUDcfja9tE9xOL8xP
EZRodr99W91RpqLr7yis8ALxV/omvVdyhU1jvdLwK+342ixYyEZqIDe4RfUz/3qw
XyXCOKtVZM6LarG6nhDCAbbXWabVKILJOQvNjySssM406uy6UGsJrpo6SIPK6p6w
Aql/vA3LNhAUekkqjl/HcdimWtV5c34vjjuNZT9NAsGRBeB9Ur5ZMacvn4Q7V/he
rQufkqX2+42im1yWVkOZ5FA5G1BGdg83GQwZKdAX5wMxcCBJbUcAvLMUrUfdwji/
shK9s/qovMPbIFtA5kbnWuekk1xQR6g1tvxdpz+/035IKw+UQ10Yka6DbTW0vW3t
LbJSd/Pzlaw7fWLdOEdLwmPnH63VSToBFRj1894f3gzODnSzBgjtszMqaPw8pEcY
Zt9oc91nIAF7EnwMhX0zl/sNNGCfF8U0CqwrWH9uW9jDpUmLM0vphCtYzz745RKH
3b47+0tRtuSaik6gw0710hjpc4xP0jUoVC9Dd1QDgTjiUPweQTfg/0t2Hrenk/J1
d0VF6NjAVFAms4K/v93E2QKTY1Hfh3XzGfKKVOVvkhMIef1yrkGCSk8FES/Uoexz
qX8aIkfbPmEGUlxSXqXAQlbrDzuebjUuo1y1UhArhZ/G4zm4Uax5fLN34kQLLwo+
fEJ/HnhPlglYFk2rvYZQkELhfYAUvej27sM/GqWWfeTHLwOPinP5Qd17kUBSWW5P
7+B+3+vQ02Ym1UVF08GKZfmyMqMwzlIRe9+4EFfd66DQZoF0SM2uS7Jz1xaG8j7G
JY7cJGlKOcSjKvRKfeXH1mWBoryYCW3zb23rSmbIk1YAOnz9s2QnVTWkl5hF0QrT
8LcWYBb9BqMIzyBVbKwohm23JYgOWlJNcdJpQ4ILUkPAVR+TbKfnakbPB0avdVI2
XIvYclXOi1mvBihMz9HIiGTCXEXXE/9OYgatbbOxkMn5zAgi09uXlZlZO8686H5O
N6SATJF2Xl8MhbVgmQApIylaiu/GIDXhQAYP+gGb6lsaTywutjMT/N79WqVpPhfT
LHj+F2grjuavquCNCk0OQ35ewfnQEWcXnH64cWX4Hd1MDU0GK5+HFAeamc25IPdn
d7qgrZ1XB4Kf9KjN5Z3L28Rnc44ttAhyawlHSaCvcpgoHny4nXuz5XiJKQGmQgUR
80MI/2bjt/jPisp/M+L546yIXJVzbv1kU3yj08jtXmpdBPqbWLA+P91+DaNJMriL
H+kvwqaXxw39mr389l4g9rfrggXYrPuZaCwvrKpkxM/dCn+EFR0UKfRH5IdInzpu
5mSdXv8qy56cBWnWoFCxbnirL2w3EdQkrbXnEdVf1eOOykJnv/pGk0Wxva4j8iah
ixsx66QDPC1HEl4T+4UbCCzGpOJ4znmMriEXSUpC0q9r79wD32km19PEWPzsXi3x
05ux8Zqyxt1v3SeWRiErSezXO1b0XfzCRFVe+lUYs6Lm7k4Ddjyqlh887BIQX9mb
gwm4k2HzBWrfcoSzFcZwwI7Q+GwiEmAhVMuL21J+IyH8h2sdUMDnDycZC51w8Xcb
zs4nlIuzvRJWo/lt8+5/CQaAGxHdquVzjo/AymXi8GPoJC/GweeRyJf+eQ/WGBa9
2qdxUKI2Q/T82HhfqhJ9odUI7EgfWKG/nc/g1ZlHnFVLr2ltDMLJzRsl8bTkywG7
YtEgCFaGyWcvYVR4+SNkVoz3qKNQDhcNUUZt1tOOHomIhCrmWceggM/T1pTzYlYH
+NkEbqob2hM+FK0t/xTfmgms/uyc6VCI0BkTEpi9yJohL/xDJfBDXffwz0xYCumb
3/hA6YH6JqlchiIm5HwwwYSr7LqZ6gAe0o1M7hcH544SrroLg3XRrQ2b/D7OIxxi
73Rqbn3XjJmWJlSEtdNDjfsqdMf0Ip/y/E8NRLISuAMa2trZhRLtA2DWdPq96on6
zXEeN/Tbc4eQfNPXtEllF2Bk9Z8h0ITcgtsHKRCg6U6Epi2Vug2Y+nRxAOJlv4Um
6zqa1Rylu1rciEHaore5H+q0wZXqfNrSGEG9ps3aYv70ICQrOSjQSnkK05VxPtej
OOxj9RLL/9mfYz/nZFIMrAzSTKvxNtcX1GwXAUE18qJXLxMbCR8y0F5T7FjNj2rR
K7XUwqSOh1fKnfNqg5pS5w/EfnCnETGwOa2/eQgwxuEiyr/jNauzicuz2zwcKB8u
GzoTfsiNMv0JgNnD6Cy+BLFSD+G8n1XgsZ4EKoD+a3tfidFOSzlFVMYHxVSzWTAj
4nCnRp5PARr0ruhhCXerjc6j/fiXTcpQusKZPtEaDMql/mFcnKClfdY2Fa9YysRX
vLi0sLVKCY0FmuG99a2yndGpeYxohOwhaFaCw/6T7kVMHKG6ghCrbxgE26aNqiuD
0rPmOvOngPVDOX/u223qGASVHhOHNorM0bhsOuxLFN6+geczFnbszvfSA5rOlHDy
n1V145tmFTWQBwHE9xd7B4hK/gBen++cwI54EIwKHVkO1TpNucHhPN5cMQywSC6Z
NhqumidIVKU4dLFOPnRdp6NCIJUeuycgZikNRKkUX9allH85M/W+njmn5RLhA7aW
0H+Do362FTJoFf6TDk7PCMDFLovrqSTBcjhQnvJZxuxCT5WTnVEWcHzPS+RFXq6d
/242GE1nFPWJuSWbAc/59eIhklhuQNPiihIYeIA8YzwOPPhJ+92SgIqW3KphQ8VO
3WhC4GkEyIjQK9OT27HghTdg2DlDRaTjHBRJEfArHOBTNQF4eMB+VBLD7tzS27A0
xNvuVXBhX961FHUxXEbViLWBs145EJEKf5ZdHuHA7oyG4oDRFzECkvTmaxLCo+wf
i9phuwsYi+bX1IW5Z8i2MiEOVrggNm73IM5Dt17kVEd1dAOXWh2svSdtTf/ICrwm
ekS9+qsFuyVpzHvyrPxl4Tv0tqZ4gfw+SDZWSmeukwRUNE9PiVD5UDsvmiGG+NcP
cAn+dKdjqK/xgsGG6lpt7ZVdTOLb8I967CC3d0g829YIMBNc5Gb7dzWbm0eoo4Cy
eMcqdHgLzgB8XgZHCLSRiRt3NaqplqiYqiSy/4tebhsciX0jvkAErSLDvJj/kXzF
Vv33h6k8aLL2qx2u5f6M92Fi1vi2X+XCqE3MluclWDLpZcA4TGuQ1/jra0FhnJ08
j78DSeMUWpGqK6vW4feENILhEDRjksspS/f3J+vgWmVGdM+sqoHHHsEwwfYt3Tb6
DaeC3a/0NxvzX2AiiXQruatmPvtrRogSjoLVFGWmCzFvrckNBfgjupd9d3Dzsgc2
qzZ7d2uGLTfUkbMOr6xguFcv+kctAJYl7mQgss7jphQSgQxhQXcau5x1FgF6tz2u
ajpFtp3iCOqaG05+8mAIzEkXLhSmBAfKipSZe6BZFF7OraddThCX8xTPQ24lLM3D
V8bDhUsphIJvsz1PsXhmKwIzlWtyYtnLsv2WwkrIsV9UMd5RJLp5RcVSQKEIeaOI
Ie0CGcFlnuUeDf5yGk2YclmOQlBrONfaCoFJd7GJgq2i7QXBAZMBiIxQhjcCjvRr
TTtyqSdOejcDaMR57LwLjggimDRSo9euk9iEYmWqetftcPIzM3+hXSAPi5vLNFZv
7m0JwZ6mROpolREg74N39e5j3Q1Uh8l9oRF/qL4K59zH82MI2q0XGiKX0KShIQ9e
DSeJqiJuvZew1f6P9KsjZlXZggzXgqtcJiVjMOEv1OG1IJHcn3Yeq0yzPZJqduHu
sDVrbkHSNT07kk/4BMnVSW51/6vFrKCftuH26ZrzRnpk8Vs1X6hGojJZaB5rYRG8
lxZeGyXc4lEyNWg6a5aewISnzyHFf/3QJ+V3OSLyYXyZGfVexUCEjZx4+PFhk1Dy
X5GQmWKREUBppBo6Gxt7z/xpKNH9UYx0G4AZ6+Fp2wTuxkya8olV2HUbfYIrdYvf
TZxyk0Iq4Qr4Pb8T7eFLOlW4I607V98L47+hBYryhhJMKMdPfCkuUtyzTc6IhqYp
kOqA1VYKzoFX8yj68pprrT60P8NKRTB+TJNHxgLa7oGRUIsvS4BRiY/POyoYa8Wg
jFkEhoRUFXo1RHBub3atECHcGr6WKF2mCV/9kEw23iNp9YcOxf+EkyKP8eThhRIt
T4M10YOR0YdXV9d8G6BNBlIGj6Ya2Y+FbzyAKIpMrNYzIxdVzsuZuu7RHUQLq5nC
+hTJ+vGGpmDHKFtQg1krejHnkmv+QiwETfKPL/onbdpVlWdIXMWMr/F7ZEUhoE9Y
hnLRCbuALIvpQyIdHonrR0NJJyoYOl6OqSf5/ht/itsBG7Z8+uTn8xiy1Iq9UELE
1SILn5JemL79E1aikj/btqTs3oMzWw43PtOfV/nYOW2bAboOdkGFIwUVjLCOnJz8
lVO79p+VIGSUt+BGu3oyknm+gBqLvsyiwLFRJM9DEXjSVYZnycgx9w/e5iJprbAm
itnGHNqRCb/S8Bb5qu8LxwzqCW5XW8CedvZiOd68VqAXk8WdPPaOBTJkr+4lyI9S
mR/DwhiZ0m9Z4LalQBTtKPJQ33VEzNrp/5OfViwn5Ojt91uh4bmzr2DgSeAppufH
Ok+L08qz7u2dIt863QE/AWithKxT3SchS+46tQ8+J90C1hVcCiKclAK9ujhHmcfm
M7eiGxKAizJVTbu9WigPQ5p7nJ2G/Ze20Tg0igu4/X65bfO4NSBcFRjb1+my83qX
mpXurf4gDfTa5VgA1UeWPn4yXf+NxDhTtVMBlnvRyQZHHX7Ts5oYpgsZ3M9J/dmL
4o2iBUDv6n5nSR2eFdexfvpEEVvQnT53ztI8yWfhkeKs+ej7LCzWilJ+j1yjZZnW
HIMwXF88MNy7TMVKMZ2r9WcFfXFwV9aGqja2Wn0dkRXfrU9iqWbleWyaN6X99aqP
RxlKLFTfNXi8yLRKnsOYJ0e7RmTVwCxddni8RSfvpgh6Akro4kJU8vbBao7aGL40
SE2dVGV8j5BKOAtfGCxE7fIyvvVXNxCW26NBNDzmuxLLsWOfKaRrNSWW4eXKS6RE
pMFMk4YXGHwaAwFi3+jv3C9IgCLPOiyfQDO5QP74f0NEAhZEMhdLz4aGBfJXUuyn
Uut75D8Ij1ujzBD5j2UBPKMYESRKurvPnIbeX2i+/XGIZhR627+hH3MNSGogObiy
W/lF3xf/WecTmJVYhu4vbauJOxqUnhb213+mzLyovJcCw0QBi1PVPnRfY6pcwzsp
Ltl8JI1TWV8v2Z7wOfQCKaE+zf/cpaAeo3dQG/OrNFRJrynhNL/9UegDacaTlJ1O
PZOXg2hzumTeuRMsi/aw22i9iN29LCxD5mmPpaOWBp2+OllkUtcdsaq9G3M8dNVL
GSC0lZNHN3A7hBmviLk7E3qEOfNHpdcmqovjASh9lDnPHlRfo9rAN4AfazJtUan/
c7xlSKtZQ0+IVUanyu0c3HhMyo1xegX6ReH+iaT8XSipjOvO4gY66TkA2U6CYd8f
YAQR+AK/iZkIVyGEjMkXwmAnO4aSSDLW7h5MTPu6H93V/8nT0rkGh7ybp1Pn7Mxu
W8lFV5Hx2Uje3KhR6sBHsf84tsVU24lNhf6TFOIxGitCBzpoaQLaMKrL3wKkXGt2
EElt7nM9qJZBwJujywuscNZnxumCyWrAH7wRNp7KoBIst2ggpIKPdd6ECc6Ykwel
uSnwBIJECjF6Rg1gvLwAMhhLX9LWkxd7ty+KpUijLa1JHpmiEzunCiPvbZ/HWyi2
uaim+Nwq7zKnG+AzKQR8kx6zg8QLZGhy1h7zrXfyPloUpQM/P4ncb16Q+SvF79bB
7iKJtG+OQcHIe6XxLCXwwc6TxXBlxrwNj0eXfG+CGMdrsZOCFkijDy3lTO5z3QFw
iMu/8JJv+CswQihx6k4k9so8DT53FpvPtXzAV0LSW/e13QFnC/lM912mY+67PErd
ues2ZsLeQI/QJHHBuDbMcazWsY/+FpulVNS57KzIshJuPsQ8F3u0LNCWxWTYawbd
RxZXncIm7Z/4jMj+i1Sv7xBdPfYlY/NKf84omgVfPyO6DC3wc4a5fQntSC9yHzBh
42GZ/uHgVFBKftr7b5cvxAMYdRUVqVGJOwLjsuTjmukpuWuWGA0gB3rRYaPWzRUf
TtiwEjUndZptb3/8ADFvuMoOqKd32DVa71lq9+Vx7NWTZpvtgQ4/MlmhvNm9sEmr
udfTazkfTy0R+nQdz+rqM6rcgiuZpWXBovV728khQlz5w5c6NS9SA37GUeLZLoDf
czY/BX5gj1hfFFma5fjt8UqBXUqc+a/Euc2V3WIeyzYr/C65kGBHToa50KkW7tJe
KkdagvxiTLiaIVmF/OMhtivewHWUxz/ZLIOpctCPubSLf7hSi9hl7MkZfCvYuN8h
T/C5ujv6d4I5znXJTkH6bEMnmRwhohtkVok0UAhL22VVyYDQiQFoKlp1g6u6RpwY
1+KCAbhtpFdRRz/AdBRiuOFBnq8JbXzEhoT5F47SeD/xw2c65MfW1L4GBM2R1736
ZRWxUFHG5S7T7pKVh5cveODCkIAhd5W8xFGz+LtYG2pJzvvj5BX5MZZFF+g4oSdq
EfAlnqx7XsIIf4xouxkN8SWoA/1qr8mEj8yMFouG2J/NBWzNzqHCTfM/QHJbRDKo
yoT0wk3uUOgMf3WhcbIYatyKy+Om+Bdca0RgFQpdj+DEkABzCW/rZuPyD6P9UT4H
evGkHG84gLn4y9q/owlRVMM+AkoKUxRs7+CrwS/6Rzo6FuneKI0n5nnPhq/soO7z
aE01lQlC6jEK1Jo9I8IkBuPnzyStzQ7EAH+/d0+YpBorw3lyj/wXLy2nQ79eT5iz
WHW0reINbNwIsOgi4nZ1PS88BFdExaLqDaEIgcNzay8zMCCAJ/TRgcyP/6Gt/J//
lk4vVNpYg5daA+fjx6aN0oL8izRfQB1xgXBxKFqGlVNj8AWd7yS1ELt6CIMVzbrJ
O4pjP/k6u/qSNMh7V9SPDSelsxBVJ5j6Rg0cYdLYnT3XDzdPU+ZeOnB6pt5BUMI4
MRUHIeyDyHp8AO2XAx5WgFwbtod1VE2GKLE2TYl4fBKwCS9B/x1XESAui/VqyaoX
cKq4VTr6DmtZZMYLaUdWbQAnds+A2VUS5xDSBejAlMph7Qg/BDLZklxTEvyzgDt5
YkgdXvEcmH0cv9eCH5qzdQQaVAAnPXXIJOvNW4axH7B09BTfHZeELgoyVIvPArZq
fV2tdaKdjcPvZ0cM1iXow9iaF2PxVrwICNUTn56f8X0H177R8KwICoXfUSxvjGn2
ohm/mu99FwgeMtCl/XwYFqhgfDTnCZZEP8SvW5/NMRzePCHNeTN46yR4wko+rNuS
fBnmokXxvtjrMLXwl0d7yD3k/5JTT9zEBlhItQEeZugIY1AHDSNEFQ/J8RrPwmZv
1B6LebvOPHwQI6XH52kwd6kLQK/vBS9PIFimuCPWnTbE6aN8TDe00K6pN4nlAo9k
KYAXJETvhoWNJk8qsld3+bxnNoB8gn70K8S3sPzJD2GW2P417BIQomtwLnqNr+R9
/MCyJGWQFo74nUEav/pl/DJpDq+SpSzFiuCMmzE+5QkENc5QyhgeT5Ece66CnyfY
OqRmAe9gCktuWSfjh9HvzNo17v/Kx7jc7lIpbX3+ogadXYogeNbPSiLhAa+x+O4R
dPwFB/nk9Bx5ZLI1KMnqzlWVwtHlVxXy7vrT4kTA7TRFMJi7ZK9hsl3fpYQeTNYR
oBcrQXOigEd7nqQ22zuI+95ptKpE4bRSoYP/tZcqMzn9UluxviJDWfafrz1aHA4F
HippC3jEDPezQoO0E3kjys+x3uwL7M+dQaWwxsc3ImgakLy7x0ASN1wsXKn9kK+s
d0nSW0Ge8esB+DKmt31IBsSE9Hy6r/87REUSIIZP2YdqKJE10rNEAR0kE1DAH3Q7
QQtS84iolFFajqVETm8GQcz39T3xlaVQ6HAbbziZa1AOpssYI8JFMVafrzMBc+bF
t+H84UGfOaNl6a3hVtQECXPTlPIaFN87pQEpPVHA2pkMXr5h9F3Q4AwS29t0J8RX
ng+tnGuRjXYIZp4uK2AWo9NrjEu+YQ1VR9nYciTpKTLcykMXwkKbkCptKqD1qk17
oXOMUC1urHVT+KUN/gP7mYnT8Wwbf++TkcBiQpNf5dIjMfO+6zhtP3Pc1NNDq9Li
4Z/of03Oq/jVgxVbrlcNaF5kw45WT9c0gcc+Om8w+xzdhZufe0wuSQyFcHh3UV9X
EZiPTPo9/rxjszQ3bG1voQfhxiSXgLmw6/xefzTkXUKx4erajlwZsyTRHsyD+wpA
ZgUGX3o08m42biX18idXebmuqbcwCL6CWd9133nvQMki8OwC/kbrfx8mnU6t67uI
PCbCKnukMYJde42GNpx7Jh3VqT+L+gZYikAMv8ul/wW8r9m29kYBaPL7b1VetI94
Lp02cbm4pby39kVOqXscHAsdxhhsJBAQwAi0deJyOitEP6P0dC9MchA9vJN4ieTL
DUPj6b7cuSA26KILqr9V+0/OkrTCLTE/d1MHlbWhIfXh/C9DajGXzq8U9kmeqh//
YyFTYRdIHiFqp50oH/oiWZbMAiVgcG0GhmaKWhdGa16zRePTTU+HVjlfIKS9YGsz
z12g/NlucP+F/AmSRWdMJv+1t1xeh4uyDvyNR7eu3hLLFdQSmDbiqDzp8y6Wxl6V
AVZLFts+b+bO5BojC+G0miG+LT08jq8kjRX7ENIHEltZ7JjhwTk5JcRO1q8P/+PH
8MaPxV+g1WoOegmvLOQsB4wxBscTtSKecKQ9twGQohObp0LEJyZxyoPkmsoRu+4U
jpCZXj/MiMzL5AwlJm2JJBJlgKuiDID2dduEVu/q+D5XOwrYatvX8t3UW17v4dbg
NvDzBJqK8AoWKKCx8Plkrw/YcQ0bA4txelU3+zSEOf5nRpXVLyl1Qm8oC/qfozMS
LOmUzjuvOANlvyBPjA6mcZ154FS0KL9ttrFwhKKvlm3H1hAvFcFI6gicN9LF2xk6
3H1IlDEtgg3d0DraEOU1i1/eX2M5C1DtO/WgRhQnGzlT6aNuhrvrALAdIlsZxaH/
Gu/7DFKx60m+PAQsEeeb7SHUPruPLdTu/qVK/dWhhwEbYde8huEfrj3PVYjWNLvx
fGeHdAPkw5nlbdw/9aIh8wx6IgKF29pK2TEjcDwAHsEG8xPulLbexAThQroWNAZg
QjX3wAR0f7jfSsb3HP/PTPpYASPirPpFbsiMQCUbZ1dXgidoi2+v4pOqQvJzpEBT
/lntcPPFk/3o7bAk0HIMMJT4Wcqc44jjkENiyIQeRu0hK1rnoD4Rex5R3Ex7EOPY
eiiYv5TrGcWGFVLrDwrqhhSjtJyDyp+TGR/4PJL33Ji2PnN65ETfMYVBObpqsMUG
Wm9Lc5StrSH6sSEuNXMm6Fjhhi9gyD9Eps/B0bh/Qbj6X2ue/piqOD5XUolL/uLL
ZZWW8oAmIM03s3Sju13oLadapHFYqzctFAcrLmsG/If/J1g0g760wLWg3tgBx0e7
oWsiW1QOVV1TwV3D0KiE0yUBcUjIhJrWXzW28+mUpIBQu08M3Ay/OnUMkadvHXEi
nAjsqAYcXGqOnK4ZLwVypBZmWN3Ep4hiHaq/x35LQVhjdt43nwwSqHtk+m3EQX1/
ggG1O1JFE6ni+3fEhJBaSOmeCHIMjiR6T79xld/krYK7VVR2OlqdqsQdQwCGDMc/
dMCySqzZkd3NoLjBPxWu9/vsqcGLp5taIh6ZM7IITeTZ0vCQyzzCdgmIeAm45Ytl
QZIdxiE4xmkVeXD66st/mC9Pu5opr+nAYhJM4PgVBryRjWyHCeFwDNmsw9tChhNL
yHbutIuoC6RRtDt3hv0QzGWRrNf442Gh0pcxi4akRuTtv1I2VxRej121rHyxytX1
UdQSnxYFPJViu5N0bI+77FBPPmBl5ogrOj4/q8sF+/E5M+tXe1yAQJvrDNkdNaUU
uW4QNUKWlHLcsAYnZ0b27REVnZRb30zwtZsuu4WVmCVP5+lAA6FAJWL5J+QPrOvW
XkINOgcAcegXW9fFO7YgDi1/9dHDFtMw3p+PnFZXnqrLC+rcqe8bPqI8Ct4E9OJW
Vy0xILnpY20vWWzEDUHk8PU53Lsug1K2bXL4CRHuY4jCkAzVLK+h4G50u/6ixdSk
OPhCONEhU/XEUiaFv6ueRc2vaPyt+LVKD3SDQ762PkJmPgdyOQowjyUJMik2rlct
HGan/4ZJjHjGepnF1tE3TvQ6MXDtrAlMMHZSMWwAqFtoZNHovfIN4FvFX/k5x3Ke
Zxo0iTC5ODm11+lCDE190HM4n5pF6eO/kuv6hrVpVj41JKEm3jhSuQ97HsZteiJE
K42ozNAyNQuXbSiEiXN1cQynZ+6ENT3GIX/g+f/584PNziBJoR0jpRe8V2cqq5p7
5b7IRN7x6Lb9JlU182c8Mnayf9fiidoGoZ5SVXZq4IiNeoTehBZdA17uHOuXO/m/
OZ3uCJ4y7zqX7TvqDkBUGg3eyTrdNVutEFueYaI0ZzUvONNk1TRNefyTPWfn1ovR
ZSXfT7Agd++GSTDVuAr1zYXkNjrDFLlqIuHOdkvPSHtuLQjQoakn73ZdmdK/Vq8y
BCKurLjY8YqYp8P0ys/vnspOmRtJ+mRgW/WaF95QYCxO+3B7wBa7f6z/Ur9eG+C2
IpwZNfhlwfX0mJ8bZ0u7Bh7qnXce67AgdcBJm3g6rcH82x0Qc3Tp2FCkVD1QWyBG
DEthcyZ5pLwnmeGlk6LfGDhI9tbVUhW13o0wGI6vl+5nbMo4kD7NRDk92FErF3ah
clUI5u6kyxu3kd3sPdIskpxXnOo9fYU9cNo+G6UOJFMdMUUUoYgy8+hquIp5jQ+W
aB/AOehDRJegR8FjNqumH+ljPwwwicPrLwxfkOy57JqRQtmYim/wyRqlwVSzW6Dx
0UMzju2QvwzXHGDT9Y+WUsB5KLX/U0I6TtrrsfWEIy6VOV6plZkcr4Nja6KQFyLN
XvKQ5NkQbjf3mvWc0j8i4fMkXun7JfOcXzm72nkv4tdxSGeVb5PWkc+SkO4Cat2G
tufzMl0S9mVQp6t4wrFg56rlygIK1OVkX4mJttLCajBs2ZPjnCA3ulAYBnYDJfX4
zpjM1rdjEMrOeRU0H50mLxE6Udfwli/5LzabHLFAb5MpaNzHaWYQhdvuZvnKmiA9
krHjcboUhf7A4hCo0JSTNSNxp03OPkY7TlsZg/CR2tzl7YNUv8GypkaWDqeg1+0d
3IE1oX5P5GW36EZguSY+/09TMaHWsos+TLp6TYotUvqf7z44BPXbeHgRscOfP6AZ
66wS+03mgHMTAgsJN05owJ+ZW9iLMHhzDO7Fwr209+ueJz03FF2e5ImFu+2qpzN7
rpPf8Jzz8xkznBXlOe9mbHY+KNZ8kzQjt2pMqmQp3i2gVAXvAbTpoIGk9FEn7nrw
KBxykJJnfFvPxVO18suTfRT6q5LY6Qf0PCEc+Ep4cQkI+zTDHeB3+EmPJnugdHOQ
QkEAuDASRoVmqS93XpmMRsDUqGVS6SKY96riXoE2GjCqJFex195Vj4oWwr+VPeD0
XoqNvnzp+ITVbrHCxvrAWUJhyzTxJCkpcVKg18zjCwtxL5T21+QIB9j/7Z6w9PoB
LfMn/ySLy3+piyh1yj6CZZ7/DGTHjY+19C+V+Zz+VGcqQaNfOmRGOyIL1fiIp76a
ga9vkFCZMZUS6eHJHKMRsXFGvaOlPIkNaSChKS0PmAJzmWKNZZ4KGXPQmO+v43Gy
8K0cvAFp6TxAzmEZCTEDFqWlGwThxIsc9t+iQ0d5aZtHdnG+WzvBZWKRQivySEWs
02PpocA0w5R8jWSLllrdNS6HjxpJfAwv11Dup8DMYrti0B5gwaxNjdJkYO0wHImb
T7fggj7InlesjFtIisknJR8177FZMW1OPyoWSQ6+5v+rdYeMa3VyCyzU5QMpZNb8
sCa7L4D5RK/wtcYtlDGAxhshYoE1pmU7Y46g2T5GcASkaXJ18FIA14v3IUQf+gal
6edGCwYRwf+Yz3ntyjupieqSHoUMRXmhpPloFlsU0QgZbuXEh0tNbuAyWfY/a1jy
rIAnOcPAWYRnZP/CezN2lFLlhQN/OyXjHNf3zZcvKXic1lqDdX1d/kYAuaoN4BlQ
GrU8rR2UN8jeG8jw0XRZQCFVSiwI4VTG6hYVjZ3O7l2Eodn8grqFaUuA2ZmsJ2fn
hZLMhYt39ySLy4y+Iv+qzL+bgI9YuqSSv2wyuQunBT/JgLG0LYsoqjU4M97Im6JO
WvurOT4FKdTqq+O/Fv8VUlGlRvbNs3HRAYEvQ1G0LOYtOfQhcRrAK++B6E4sOrYz
kXnVfh5/VhhVoYMuIsRmlYwTeSulQrYO844wqWOBXV/477kdeXiOkhXSHvz13uAf
7zaoBrQ8m3n3xY1j9U3KtQjxXXBPl5/DS+GUhwTg2idFMxFxMV8MYHaN4+rIZRL3
XB/7Q+IHpOIjZok1QCrZNjI1hj2x/es0dSb6lqcoVMMVqJ5JKKhOtBLVBHwTZpaq
ZtxHAQXbLy9B/nPC+VQ6/fH0I/RAwYThv0FG59+Id52yqXL5XHQqOB1FhavPBHJx
1wtB9GDpZa++15KAHhz8l8y4G91+/7u9pYd6Ac+LUUTog6Z0gIDad00rt9jvCXAO
sHqDHHDyaBYwVyuSbJp/+bMFmQjuT8A+CitA3gD+Kb7AQ30xQaVcJ5hLSCQyln4z
gK4TzcFX+XmQK4FS+6ZQczglhUMFKkvtyEelsNyfk5eaVghKEGJ5CJBO42sEENSY
cSk/3Qsehq69z+gV3J+UAb1Rlb/XPJMRCAhU4NVlmPxNFVDxaU++kZ7p/hFYyqZK
ZcLLExfj0Ialu7oULMLA08XL/WZtSGsxg85k6rAdS4AuphGrWEnf6eUIxoxMrX59
BiGSizs8URFUaCpjlCKe/dBUluxmV6Pb23+de2yzk6nApys3/QEIcxIAAGyiKe0B
RIxVzoGpE7WakyuAKleDHQALww/sU/qkV1ZHfCBggfzhiouMhWeVIgl0nQEsnf2m
bvrUw4qxGzMHZfha9OpWFS/dRpJHeq61HiM3ZOmShfGBHsmrOQfxLG7tJBCelnqW
cZpO/lBJQFn422ZpajE+rLKdwLLkxKjUIsD+UwNqxGcKOqB7AsM+TPYQL6zz9BEZ
mPucROPHoalsgJwlgraiDkeaqT2aDU/T/uhsiAYtaeoLOSwJsoWJqG+uqY3ktOqs
a/8dh8J46qvKTJsyzhkf6NHCFTdYfAqEBy8J1e0r0i+LbgVxv/vBup9ASa3Fqt8N
MN/HPj0Ga0sUL+lerWBYFjSb8tgvK36nXEAz8Y4g1W+EvrjF2791arMb7wza+emY
yVqUpqs6RotslpMmWU8EMU3+0gL59qUcZ9jkSaKVNCnk1lialGbfBCK/hCBzsGOY
A/NgOm+XxR+0YKZIBZWt1iICp0ojIcp9xC7HnM2yrmUK0uM3xYboMO0xHu+6AzgK
4B7d51KtAk1jyaHsEIGRpuxAn3n52MzUpXzAbKsNPJsKEpe0aKHiot1oxwuuTI4/
w+l/+J/7kr9it1osX+GKexXBmrxe+ui9PP9tZ3NEVhk/kZRjqeArbM0TbnoyYto3
jrYMvi8IEZh4+wNmAUQ4WOvQYwcDkFQwXD7D2PPM6HTBmfXY9AnwRrIa28bElykx
qcautNnpO925qsteoN4P73Ic0XSDgaTlLQBJj6lv1pq//alQFIc5V3n/4Nz1oqLG
sMef+iE7yihBUE7O7Nrkv/ekap1MSA8LLUvIyPAnYS26O5ShZ5q4msrdlyqRShmi
CDQhXX2F9c01Yop1zFFmSFCCbnBsACmBMj8uOiyTVlZElMOqjfvJzyKobLf2Hhap
m2GJTiP1ORVJobEaJdoY7Zf0y/BT5DSNk2ZB+ehhFrKghOc+Y4MIbL1BXXfCqVba
V2PoHGSiyqVHFISKKBIHrHbJofz/M64r9aV90JrriIcvDsnx1qQgOxaSdwSZLRm4
4QEYdqBKc9oatyn6ENeDRm5MQphx3uH9XOlYpGGOTWireXlNrsplf/pRlQFzP3m9
NbLQbbnSRkwY6AiKe9IMKSzPGlFGXnAeSvGqC5vJ7ScBKFD/rPfs9Umoe/O8M0QR
bioMgX0rWn6a59kc6tbyS1r26XOnI4E7HcbtxGwxk0c9ycMof85XvXzwf8nf0Ko8
pUi2mgWTt8aPiJsj/tSef3De0l1Do77D8kpc/m67flgWlHe4x1DLtC0H0rg7m+ze
flhdpUuDeLHzrogPH0BUs0gf1OatdAx+jqrFebx9EWEurkt6wy2VDlsIdmSiaiS6
VCuDwcNohbCRxK3b5m3T1fO9JVF2Ip3ySL9iwgVrpjwGUSks3uf1JeeRSwdiAELT
j73rNCSMmHAyMi/gItEkBpnIfbhfKP0e++rP8INA5xHp2dv055o56zxo2krsWGB8
xKLndl3hkgObP2xmpJTDerU+Pneeu2uMv8w1QKhoYRsLNmeI6mNbwQIf8iXxIV9g
Gnwx/kV50cz/bew1LZd7jjFx7fsFVnrD/oABM7oly+4yXnajinTDmlPxy7L1cr0a
n9ZImoyxQiuOPyo8eqdQgU2FWuuR+MxgPb3K8r2W+X8fUtuyc4TP0qNzcvrJKpgd
ib/iU9VWeQ0j8n7wvf7UC3q8CrJfykv7M8TOnXGFGw3jnyceufOHTtgydYb6eeVE
jhIcQ+B3iJM7nT/zxxU/ZyPjMj6dEuUTPwnHd/fRD+IgDjr0eiUmznLnJPY44U2/
l/ySYvnhSDbLki7ro8l89JBVgGtrEqtyn0OdLzI3HEMbHGLqeGg5Np+UivHpT8ut
1YzkocO+rMR4kZm0/HnkmuGG44IubPt0WvkWXZuY9DxfaKchNW3zXktkeyov/I2G
GhbnQMr4pftttTQB3amFwq+pZfzvfKV1RhZDFDw1w2/CXDbIi9uCWzXU2rTXZVVK
3L7NqvRw4gpzxvy1OC+wvHBKLLUcdjTBe182BnrOUveE8RYh7ICTUMqDFOdROXoT
ScuXdhudTFKcY2tjEB0k4kL8onllo8Nr//aIILxlPzn/O7Ft6ZdFN9Dlt7zpeIRg
OTOHgs3Urr8jXGUD1YZOswlUz03v9+XKlD1/JNpBw0qXJPbfZX3nIT58oUmrYHmM
Iejxqx9xLsE04+EuLG4bHI42msM2vxjMnbSib5VNVEpVD3rQryiHlZ8F96jNxJR1
eDlhlrAMuGoI7hMjB3oV5SGxS8HLeigEGe3ynkCO/Ns+Sdr/7MmCakCZhDYTl0Es
9vOfplMBTyQmJqY6cGyCXM0+PZLA1ts8n10ot8z2oQwIHArApdPfggqAgBxf8nKW
Nbz4kJ9gfWI3vjo/Mx8ozbqSw6JNXjPaGWo/zEgAd8TyOZcxxiX92EhdeGRed69x
ob0eiLwR/i0veLX4S2x+7eQ+cQLvpsRwblmxGZCQts4HOQmE9Jeemfvc8kqg/GCu
71JW7kFh/uSlxHdaSAT3Qrscu62FhSnGkePqs3Dy/cxrduc68CT6mO3BjbOM0BBm
h1jB6oeQWsFg9osCdk+eKtjskQpW3VramZ8aspkikrb2HRe0iJY21e5I70RL6hsw
g2gS1kq+py9yVp57AuFBI6C4g+I9SpQnifmUdlqy0Q4SRKaRHl9eeAd9pkkZ+v+s
seZS1EqOQsKjZ5jGZuFl53H4Kdsi+XIbfd2ZT3osJSYoM213yvbVtkn89us4KXCR
yLO3V25ZEftS9JQqqtAj+tNSUUR9T3uDzVusymQxoGSYSQOrjr8davHXsXifILDi
bvLXxthZTTK/qJmjFBTLy7K9eA5wO0UpGYWKLN9ydE+1OKtXTz8qd7W8HHA6jnDL
zYy+GnSAze5FSdhuirbvqlvcUMqhR9Cgx/dPz9CuX+DZQ1TTqpHGG53oL6SrDtE3
sdiNgcY2nHeeYKRNGD6jfXL6mggB4UilQ21bm+FZdKRpFy76n9QXSsvBTg8+Uw5w
T+3FUxlewAy1YsfvJDhyr4pKJb+IEIkBonf6Eoa0lnGyvrR9ujQfg7nWATK8dTL/
XuHvP609IPIdf2r9Q0xRtIIkrNwYKCJdpbyRtBYb/avt4MMSCygyAyerv8uwpJfR
G/tHCaVgdzbbdm8q39X2IXH8qb3FgWAzoCo+7+HvyPwEljL17mTIx7OArtJJdBDq
dzcaZ5tnJ5S73H0Mr51XssBnBisoy0hBezmVaLz3frWZF2CF2D0z3vtiSd5Ae4Ze
hkjax6HjW+qDSz9tCp44X2onDFRKsSx8SeTKKWvwZDyRQeM97uaraJsjU4pV9il5
H5KC6HcD+ftuuejv3y+tsyZTN0uPP4oJ5byj2Ygq/DGBPx0sPpt961T/hXxRMAnn
61o1zyEDmX9el+3sohrXY7VBVcl66LMfTu8FXtO+QCH9AA2rEG2ekpgYT8IPWM8Q
SiXHkcufuGx64xP6FD9E8V/9cL7CQIZz/johjUV+eg2XIk2+DJXOuJxulgvFwTJe
Ax0vBVXm0lAZx9m9Ir9Y18DT0mhzFqWmjcRffO5LSxniEm8PovIG8r1ycTc6tuiW
mDfoNKTMKY/lGAQkitseEfqQLEVZB8frWE0IgJsA3cLjHgw3bKsCMscbSMaApxcT
GwYk11MUavzLt6Y0dWuxloctUuagsPNyh7sxTIP8h151swMgqTNhkGkKn9jZ52Fa
50jJWUGDHGAjY/AxbRsnBKD5Y2Je1pfKq+0KXmUqmMiL0juEx42vyDl+pvlWE/dW
Nhwifm2+Gy6PeRdQXWWv5yLXvqBK4kRA8n/vrqO/pbyTExbMkzDMRQygYGvE9/SJ
/7DY7pP20Uz2vEq4VnUezOWS6gDB5fB7q84HB7AXRWC7AAErZ3C1bLbNPTLit6dS
VfVd4xJ0r8sI1esmtO4fOS2I86UAlanccCdRaXMye3r9BxhH7a29EZeaBgvxnMfM
UpoeCrrSW9yrLt66U9U6v/A94cy/8tVZopF0KcU30CRJ8aNrlq4i5qgebTdOZxns
IkfJ+Ky98TL5IHx3ZZPsDg7c2FXZSjOBARlYwY+QLf37VS7BU5O3l9a8osHx6JQv
v5VUO0iAnsg4t1yMONTCJb5+8hOcXw7xJ9KmYbHqH9lnlWkYLpDaLxflenTFQIfY
Oo+fA10G9OZ11yPix0q6a0XdrxOW3tZEoHSGBN28kaFwfv2n2KHoq3LfuzK/SAAa
uO/wrS1X/FuxwjgB4vYwtXqLS20SNa9LFXktjaLy2nZA0PRVU/fFYhLWY/vmLMZ+
w75rNn2+QE3Enq93OZT/x2Z0EH3tj8wM4h/LLFNmA3rt8/DfP8OBRXMfFHbzx2aS
C8uipIh8PP5yUksEf/Ek8XpK0cqqNltbKSq/7MK5PAVKhbdEUbZDzXogZ0pKz0im
JI7Ez6JBO307vdGV07c4SvzccWGmI37Upvj3dk3fF0UCHjQlsz/lkGyXMIll7YRK
YiyQbSqtxPuhjtkgGDmDOS1+YT/WmS4qIJDFe2MVTBk8JSV/cGqfl8jbiweIKMM4
2ms1gykznMu8UalBKHPrlCoe1cmOsI9JMRxOZRrjsm6tBgkPExwgE97RwZGp5zGC
5rnWgpKvGle2lPWBRxRLarDnjt+kC7qq0unuKcaoU6Smid0qUEONByfNTEc0ZICU
NuhgezS2U/4sel3w3KEBf9I5LOYr5QNDgZCPcqH3bGBeFP2scTn4Vjh8EOGgupGb
GHlfvkgL27kBonT4ZkXAyJK1A5BSFyIeOsM32EbO44R3BLj2bb/rP7vSRMYnYNQq
JfZCMu3cxIHz8lmDQWae8jtYHVU5cwtnhkU6R7ENcg5opWz8zZxyIUxbtnHCHxny
M/6IrFWX5xMe2Fb833SkxzNzIZF/4DySYtW8SBpZJuok6T4AWJTuKMPtwKjVxGGK
TWd1dCG37LLEfa46zkdri0SfZxvJYF2iFz/rd58+FXVzrPMLp7j3en4y5tTnew2s
NiezmfvudCBKVndhySuLhcGBcEPeMaoRvGz47RmQwwMgefIKbnsffGgO0u7dvy3K
zdPGilXpafozbVxNNrHw+8pa5UKN0kp3ktC5OZ181swDB40tg7NSeWZNDxWmw7KB
rfKmL2pyEqDBWCQycpUtZDa2cPMCz35OQL7hBdtxW2lg2hCZ0wX28vrt0jGhGO6Z
eeKnD35ggh66fCBotOvj3A2DkZ3cp+qaDYXl6JuBdSNPNEtKhsuNSC4jgPoTt+6K
KKfubwVcXIaAnud+g3jO6bA8krEF3jBl3zH13H/2JyQ9O2JduPgDRzLQnKJR4Hdc
IXfsue013MzJV4MjTx4fxn+4kevJM8fOVr7kcBjVNoET4Hmxx11n/J3rhRmeWNsa
Z1L4gs0BmHN/EdRXCwvJN5gNH+HPyS6tN4c6aL3/fHGjNKB/RCk57sDxPw5cXeS2
zsJMWrhSVrON01kyxR/PcwQxTIomchWs5keVDtakAvRUjHBFrT7CwgyPG7iO4Rzl
+eBzxtEpEhEgywNtRDFA08QUWhwgwIPkXI7PVnb9iM88qgP2h0vcbrb82sHHB5lK
yp4X5r4tERFXVvJ9uJsFukGoUHRS5Iug+ZwOwNlklBk/HYGusTX4SbzPsxHBKuZJ
NF5I/LRXOP95/L3j1cEiZcpkmf+u40R5dUBGSQFQpkY7mbAP0o4m1LsRm0iWrmEy
Twts+4h/5SbPqPTHX0JIqox4OlFRsAW75YoagLR2bnIA8gbxMb4W5uHcokyrCnnB
o3O0uTppq3EqukfYXn4jx9/xbAlScoStZIJt1ZgIzWnnTlC/uacfPJuZeH9tbYSb
nglXIzJczGv5lHlhk6KyZKw0es9qgjeO1efj7t4EMYfyA4u+FwkPLHqErmQIwETy
0h2lvqIH0JFGSqd0YN6C9I1+dlBF65RZQVI0kcMtrTiPWbffLacxwxeSH02VKAMq
fmbndLuEp9kAbKGBN96PZxGGfNlRHgfTSoS8AFq12Lzzsfpi/syYlzyBPSbbLFTr
DPCDKhrWS6gqWLlyXE1vfWEEY7sKdky2SuhMk1+XaGWrRNXCdEcCkb1G42CtFHxD
a01QQlX49b1C6lFmYaezn8e0vddN3szN2M4VpUmSGWfCCJqX4fBmd/3YiugFK9kJ
nAPoDB6O8gMtQUr9/GHcBEj6VSIek/o43myfbNSzMqV2izXNipNj0Mce4iBj2nEa
pkCmOZANwjv4DG7QyTXV7k4/ATG3xSXV8oGHbXee8t10rq+PSKwdaPIodXBmlP4j
YQ1DtoN+U21f68UOP3S99uCVrYpom7GjjVIck2/KKe3taqkuQZFDK5xVboEHiczf
XjJDAL+VEXp5L3TyPool7/BozyCYANcqk+czJ5GdNVex+ukzMf1goA7Nj2X1sS3R
Gh2k8IFaS/ct92G27n9qxZP7aoDsgKsftIiUpscEZtNHVNl2DOnwZ7ltuB6gp3K6
G7tvQ/ly8cgp1Ip/iVzY4g==
`protect end_protected