`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3328 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRo5n418HUi4GlaQEf4lAMgCmjPt0lNDT0WunfZoEyAYU
XQtGE2oF/Bv0uxmgfghm2Ob+VPSxb2zXQ4fbkgxZ9OqbjvL5I9wwF+iwicQdnwF2
IqwBV22n8nH0uQCuc7OEFduTzLDUHovlLf/oym+6BCiaBnyoClF8s03Wd6FWiQ7c
kVZvMsKH6SfgQpveTsUNpBUMz8H4oa+x5J7b/4/83mcPluPDetqKd5Dri6Pu1mbh
4zxwr1vJdunJN8FmsgZ/vXuIf14S3aURyyAVS1ekIbOSlS+pvEw29Gq7QlHuN3pU
XkR/Yu+CqbOeFCrnjOxr+f3b/6BYY/LlGFwjf1BYzQPRBGjzWOesGjR2iEa0nUV9
W1ZurIDqw/ofbfhGy4IVRBUmTztu95yu12EsDOPGYUN3JoRNFAyo1HemqY8AjNYT
6Mc2A/gE1fr+xtwVa6RIcHjA8r4C7LvDMYGKxqafYWmDi+hfoj0lj/QlQsLK8q68
cEdiiQZQADCJVxVovYOA3MrML8GsdDoOhG/sxBT0XfeXKAUeVB5+NxeN+D9LARpe
VsB8rzBqGKUDtixrBHvynwE4Z0SAPLekaZK561wp72PfWZpjd4qwZJgesZHBgWdr
fwwY/PTO0kPk8yIO3TflZw1Z6ilgR0oPyuOrBoGtS5UguzarFuM1stziQRSKBPqL
RSQuLb2WC2k5UfS+2Mre+zcjSCR3+YPUn4eiH9DPOpj7XrDLxrNiQE5yJ2VauYg5
/VANKVQWt2yEQVBYTGCm7aBHUWb8bysEaDzkaXBAfeJYgcr7XX0H3QCOK+TqP3zk
nQZRsK02Tt8iqGx0kNDmr4MM4RiXQyPntyGqWwNnsXTtodbKDwhAMEItJhEJ+PPf
4EGID6EAz0fBLCneCDJyEeOFBDVwXQ6OwYVSB1cj7kMXQR2dGurt4Z9kERxZPo9w
Uea3dAx1x5CdomFODorLuyAbt+SxN9DXtf/PY1T2NGqM5lNcHJJm7DfkSqIILSqt
t4TqjZjQTr9hU0wbe/1WNhFDGAzFQY770UeCWU6W2VWLYIw+B/dswjqlsQ2X8NdL
5vGc2GROwLd1ZUsZAaDpEP9LMFsKI/xRz+Bk8aTRPYCFpQyz29n8YX9xHOF0DSAP
SXhj+7U45hZJWk4MEckfBw4KjpiwahNaP4DbrXj2tjyEGt9sJNlNWB3wvPBivvq0
XAF3WO6O5FcOghti9Q9gQ29vY7LFoiEIDVd/BzpboybpncpE/WTJMlZpUkN/0zx5
Fug7s1RIRGY5unPsnOP1wMDoXsI5Xcu8kWcACD2hzwrxmnx5OKHaizMOwYP9DoOU
yqH6FDMSy6YDWwJk+Tmg64sHYuErP9yuQh48XkOtG1wddAKR5LHh2d/OlEzN/W5s
UbOG8CnV75QzzHoETT2fhQZvu24RyZW6Botoi2jtjSIGpTJZGxAYZ006bA9ry/6m
pJ+f91rEzfibzP08x2joL54P/r8jTK6IprKmW1FzggmAN5i08cxop5ePcX4rI2j4
Y4miseyVswuX12WINEh+xIFtOODCYAdiA6aAQxn8MEDnIVyVS6SPm0apZrqiSv8H
qbfLWPkjjfW0buFOgna0HlVveW8iStNDmN6GTsJkIwppb3fD3wp9ZM9DNv/xqAXu
FHniGa6X8+jEZS6esamJqIDpM4gzDTis6PFOjWTKsOBvzAC8H5N7AMxvVuo9n79F
MceGQZNMYXNeOfpT7CW8NCxMgho4/JExw0o7HU42ew2HFxRQCwNeY6oSwfEqX8FM
PxAG5VzTfHiLtvN1OZK28Y8gIuCOYUJOu8hPgcPu6lqjdocCk5xyJEN69Xg1ABNT
Nkd87lx86CmoCaYQmMLT84nGHzVCmv9QVprbDrwwqSMQbMb4QHiMWqb2oJCX7ylU
wDhLAmxh6Mo6lzBDXwfA3RWPhafRXCA3AHr0s4TLKMYxY84f8p5DQxSb7VAkGhP1
2DROljKCQAP3j22apNU+62CBY5ZmCiVtirhpO3H/OsMJ2QgcjwyThYgC9oMwzeUV
mUJ0cbm/QDuF75OYnKDTU9MXFdXOB/2QDWV23x1mrEmmnWwSAR2/OcwEwGAWUP+C
glBKQGsZazc/tkBzXdfXxtISBaD36n5r1dboFDMAxGfXcDn3CP1K2sZxbm5R+6Rf
4DdQruJOQNjY0RZduI+QsXXP0dXPEjBrlI10N/DOgumISNpAoDreNmVM6bn2ofO5
boAvcjIl6lIBzoXYIxQ22epfdilzetflNC8qjBVQmwRFE9mOXNKNxO09c4yixvOW
iyX98xk8LxYQkWWlEkdb8zZUnk/SwzRJEZ4G09CNWMagrETjUWJprB36I+FXSWgQ
qnHhLNU9APKuF36NzSLdBfQOGv18CPPhYCz8/0bgqeUjkVAYkVss3KR8rUq8pulc
WeNvT3wC3vPCkPvVNVeFqXH4y8hahuiL7gCICPtlRdxJu1Tby2LODMgeha/FZHsX
ZZuQYu4Bh10VhzjhGfdaLwLiZFFB4sYn7+CMr3Mw6GkyKVkXK2KVCRG0T/H99rTl
zYuhuVyt2+OaxtlwBx+plszlJMDw4tRfWj75OiDgt0wAxh0vJ4A44JPurvMUgMD5
pK9whxMW6sPo4m33M8gfvqKoS/0bjJNPl3Hmxubqs2LOZstvkCdoHWBBUj9/5hIA
2ELazf+09AtNQxs+WrWt64POL3NiyydoX+0s9RjBjSsOs8NcZu4ENrkQFhn4oT1/
f6Xi1JRNq1NXBa7+BRxqhISQ8C/sEAPrcN/4i8MiGj08NBigbK2m7cjOoKhHG/ye
b6Sl+5FA+ZL3u+9mspUf1kal2gNbHZZFzPW+Y0K4NS+zn336h4uZdIlRRTRKIcca
sXJfMLGnGKX/FAz7cPAesd5WO/yCXLW9p9hpKZlVDx7xYhfAyjemWIUNSpU1xvLo
FCmYdsG33/4kvES54R/NNbY0tw6V+EMvWNiR2JhZdftWzMwxkjf6XJPTnMp7FM7C
pvSFO48N8hxcxNV1BYOyTli/VR8XkZqs1aMa7g5Mgd9QcM6jCP8tjjDmjnziBMIk
OA362Ykc+2npu53EBmPNHPKuPguvMECBbDZHdzUJP4lYeFfPnXLWDOs2V3ecwnA4
02fu6PHmF+TugfrfYr0sF8u+H8vDtW6FLG8IwM8oq4CRZbWM1x+E8F2QnaTyeOUT
JcT3gsEG1GM7L0nxkNf87v5YjsV0FXqh8XkfN6QRSrGooWFk6y4c0xiijunYnFPB
vWcTq02kz5jH9juu9HdrXO92Wsq+xYjl/usNjGLItjxLmTEQYWpMfHghS1UNJb7f
xkupZs1lmTgy+mp0yBxgN1GX1HUk/FhvWaJcmy0AkPI0mvJ4RrpN2dZHckgazjwe
wgS9S5CsK+Q+pB3iJskpiCF4efr+MZVlqnMP7s5KNYvWcmWELaz0T45COvHdvT+H
AEOY0q/ok4dau11N+50olgBIuJxGCQ/dF4g2NPxYseIkqOozOu0Lco34kZW2Zjop
+HNZjhIRMsvwnIFW3PbhA//ZzKKd4OPj9FoQIoyJJ/K81j3c8uLAD5yDsvbEESXD
ujHQsvmkJXuTnDqGm+goCxEwMLlBr9IRSG+Eo7rvUqVP28tYCO49wzHe5TlIga2X
/GIgDl6LvEgGojtFMSyQlp24R74gv3C5CmpM8nC89aLy5hhtb/mWMnuQluh7ONt0
o+twe4z3MQmo43j7lN3ucaQPT5ra6+KMaX18eWVq4Jbu+/yhTEba1WfKC0n/5TIZ
dLFEZfKUc/6/abUoEoTr+IrgcpPpTD1kP9KZJuYKPciOZZM8+3ggHGhyxfiRi7KE
RQHy4lQi+KxYRJuhBEUGEKidZQeM/0qjvHBCRCA0x1mwB4R9HWDJOp3xwEmkSmuH
bqQ+X23jQWD5Mh6vlMPW3zfU30bjfXPSnEWGUOqHsWnTMHTa5hHGZcKE9clk+DuX
Rgx3eadRA8OmUftuw1Wowc0XFCSKrRxr+IojBXmAV4tmDdqO/defkHMuUoNAL5YC
Fmr/8rGhXFuEBEAes+r9D2xXQpIAWmgFXJ43Dof514KtYetqpH48eVB3956U1/cA
RObg0yW6CUJr2Do3RBRiW0pZFDhX7xQu3dM0BAwNCgfw0QqY2kVJrw9x/AXTA7YB
Ft/hxSx/2IBQgy5Ma2nAvYlIFU+2oTz4hPSr3Tqt3aZhokd1Uc8/6kr0rqDbYnux
R/78BI0wqZtXLeLzinQtern6ky/pjHk3mTsBroi5GF1Z2sWiUcz0AG5d49t5sgDQ
DCVHOfDjqqkfETn9QtfWJQ==
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3328 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1af1Y+Dk6+1SXWNwztYDhwzRq+SJpq/YewTOjrXpJC91J
G+Ihb97h6f1/6JgLWx2OFROPeBmP0Nf8GRlkqjbpS8ZjWIX3RO5tFHhzIJCq6Zhw
sRRvFBL/uBB6s1q15N6LQSKptjemBRrn63iYGWts8gEGesAFiigXJyczPHMmAyL8
WMcAqcC7yrUPclOibBIW7MROIZSq/2/0uRUU7zkLYgJwy+laMV9KYBQC/pO+QEQF
LZyqcUvCuBxniaYieKM0IUFHZ4b/7jdARuS1rimMtHoo+f58JSQLR4Bi9o2w6oZV
A2AThQR+ABXVDDAZ/Eb7h02MfR8nLZUWOnUkltf6+jOff677hXRsbYTdfoZKvhJS
n6kLLbnz+mFvwsL+twIfkup5hCYGdfUyoOc38JrFXzQRLkEktCRI19GSZii8l6GS
89ao51N1N0UGFgGSCTr9MbwZYNGHNA7IJhGixLn7o0pOo+7qzvnRi8ETI/GafqLQ
fTAliTVvY4EIaPKqdsK9iQyqYXiBySK9g1EPfIaU0UOeBivcNbrg0ezwzxZyddGq
orlecqYiEuzayV9To92UIb14RWa2+z9Dst46cLFspXg99QJFkajaNzcRa41Z8e/1
UKK/lqtMirv0ObEdD5sSAjj429aXbquJYU1uUxf9Yyyzzff8jIJ6Bc2iq9qVqz+A
fpPh82IXsNLWl4RucKpnNHYIihpgSnCItWiS+Sge2rUswThnvUMxaIFqRoFA66fC
/qMimEWfz4L3Ucn2AYRkZSikxOfg1eS3FZKuF5uIm7WBAVPmVFMdZlTHgZyftD3A
J539PIdDUgzBFf/hMmzll7RttN/h4v5Wn2OMINas+USNQn2buP15VmcXTLly97VQ
Hb8Gn5snxRj8PNqRHPQdnSCiGdFYlQYIfPW0X6RTRLCRsPlIaWyW7RS7aeX2eU+m
D+zHzC012rszddgrud8+JpyhY7oMhvnal/afTA2L8oX/PlSMfOTFR5KtmMiQ97GW
8q2Z+MOXoNQ6YrkI37IudHdsnXu5V3YCO1vZ7fbJRAc06jSEiAV4eTrsmrCnuvf7
3oPpbtGz8gS7oljGYOsg2SjNuLlEz36o8YVreazpMQwy3JpXe/qDG8ZCRFCo++TU
rmssT7IRE/S2OO/hOUFeN/eH588YZwot10ww2k11tHn7HULh+0kO8/CVioEXLf+B
0TmnvthJxH1GmnGSlDgZ1bWrtEmgjUGGCh0Xl1byEnThwfkZHZykb/+DLnLj5Tdq
UYJi2zjCyFkHSyvN9RuLlb+ozHBfbJGwvbNqNGle7mYwqK0qEpnJyh4KQc35c6G1
GE1SurizKk3fh4bzo7OsA4bjKGKn73AyGhtlhlNpH+udPUcuvZWwRDqqV3tIbkvA
hhnggtAGZKaQjTXdIHMlVRFv6QqqMRdpI6yIDXZ8kgxKaNPRgiaxlfVPqKks1Mbb
gNnnemOul07GHaZdN2AZFCkNv0+gj5uETwLVjxSKLXlOUGD42wcMDttMfRN7VkqS
S3Rz4njKOrvXyxpW4kK9GiYwDO/tkJgiyRFuo0hN6djEUDumbsx75KTdPjrKT1Kx
V431sA0H4DLFz1b7LX94ZKzXmbsI5JiFcDARdaExg4/5WGs+i8fTZO5LA3SRBkWs
owP6Pypiv1Cofgazb+0I7e2wvyniHfBqBjBX/4V4RGyYQlyC0sXA2hY0FedGi3i8
Y/loO6cNLC4Bb+/koPwWvI65v092nt0qD+cC2js0iifDPU/YXVYVlKp2GEkN4Wz3
9QLYlxgtT/UjhWTEgo8UZ4VIBMIYRT2t5GgoJhFUixYDr8Q7K7ORdR2vdKXPpV0B
wKb87c6E4kHhh/1G2Rl2XPgDqYmuOzg5UfE9ZBOIn1deFGNyWqepLqXV0nhOsfNl
z1axzpvnaIuyRH8n8iHj/WDZrFKm1uwiVV2MjKL2swXck0gAzs0m4kk80v7TWQq4
RmO2tKIZjbugqvIFBE7G1OssLmfPCeaeTmI4OG//th9RV5cbVjcvsBkIpK7oV3ai
CZwS4B6AVCGkjxGbWfsdMZ1jxdASe76iNd0lmmj7dDM1NAer6ZSWpLhkVt0xJsGG
CNsIpIHn8Pv5ld3hCV7HDITcR2mMOJaIpr5UlMZ6Il8vaApvT1bwsXF1xDhkOJz2
ELGYj8/NRh93QMRogfdzmTygTChVSrdXN3VA8i37nE6sCvM92wUFfOYW1EGY6bQH
2CQCKR4N1Jx66/ZBSnm1Wnv+AelOpdlBjpS6RKqwP114o6/9SPsveIfNs0ww6X39
ncxJIwUZvX7S/WFbf7uPR85Cz8vkDWiZ7KDWQxhNqgghSdtkiz3seQEPWbNf6kgO
3okYcpg4cREcSfJ4++kc4hbYEsgvgEktW1wbFCEQY1Wz3hTHGw1myJFF51TU2xhd
Va032YdLSEEP6emWcpYkJQc25BzyVZDULDW+TgRBgDaZWPFD1XsHq44cT3QPdqjq
+Ru5CoO4F5yVwmolKXACkwM7YB/6JRWgJi5MESmw11VE81ra1Pw6jWo0cP+6faE4
ctW9EF4V9W8kIrVxr5i78sogOmj8xXGws0Ymxvei0iooQflG282y3ErP5npvLYqq
vEgXiTIcn47OWyjr3/RTcFyjGBWSQakopG6uZuNlQpByY5TJIGxCIefN+pkcLz4h
uBTWTm9LKbXQADt9pWqPxjHyl3yObrUg19B7e7uoa+eOjOYl+cjZtuG+//O2AjJ9
Oz2WCWtM0JRWDjZ3tDiuD719LIMigiUxlLb6avzWMrk0G1Ym11dCDLAK1hJEr9tW
pKJoDQcLYYIQ/TpGQDJVBsNlgCAz6/JfSL11cwwv7GG6bZ139nZ3GorLNJwRzA5Y
YInRPXMzGzLgXDOJ1CiKzVBqWznn3luOTK5C1hq5oo5rh0RGnh2Q9dwrFGgt6Wvg
OpFNVzQVUjQ/YoMXjR4Kz+LjMKEbOLmdsmLfbXjIM/OP2G1fE83gQXwodY5tLvZX
Mm8qzjfjci17MmkWI146AKO6qV2AWe2z8G4Opi9eZsOZRkycGSDy1NnCPaG4VF4e
faMNUHEqf/7L1al0xopUZAfS3kNp+RT7XuyH+pCmcC0skLNzFbTIjR/d7QVypStq
xPdRbZVJrlNzBVNbLoB/pN09YVpeLIVWNSc8csWsu7MsrMIJolxM1Q/GMgXRP152
dawBA14hevatr+1MXKl2737E1znePHFAEZK108bRNABkHga0zg3aeofTccATKDzP
9kTWbkwAhJYSZWpWnJoY7oHdY3XQebfhPG5WUtVueBjF02d/3pIl8WEGlDXegtrV
yqtzjd94rXQE1eWAQ78oQXv04mGp+du2VV4GwiBwVAtz8T3I3l6v+lwPGe8zj5Va
xDKW5q7+zqHF2IeGG5zbSalsiGEgaUyaxii6Ik+rdrjdJyRqXQPNTYmo9MVYGxe2
5VbRS8VJAS2jYHhePS67szWQPf2sS7zKf8soXElCtgEqDFan9/vQ3WDm3MODU+Fo
1ydloh01u/zH2cf/Le8NmzqfDCzPmjJSsWxWo4/ripa8Q0/bTY4pMLVRsCD2qXCv
6TQdtWIOePpE/+Esb0PorzQhB+lp1L6jk96tEev/oZirKM3jySn+RXk3xcveAsaf
2Anqxnye9xlGkjVxqJNARQkIf/MogmmLM7CyUmhSwrgtJFlafWL2D8FfEKjzL25B
tLbIfRCdidizZX9dPro1nSwV/ZZ0n9DBs8zQdPsbuUlj8U14Xl7ydP0MrTCCzDIs
jqGxhTko2aXONWKL9ysWoJCCDnE/p5xosya/tl404RVvITMJrLICXUJybhhyXlnN
J6S9zZr6OE1T6C+FPcb5hQaEpbn09em2SlEduuZ8XwJtYY5Y8pz4VGQpmwHMaL8w
ehXtULBJevKJje9nYsIFf4qjMOmriAtLbiSz6MK7WaB7a+v/1K+j2476552WdU/g
6mp4avlZDc8sdWh3MUfda7YsW1Oamg4+0Fk9fajQRjTz1NDuf23RzevMvlztIMmP
Tm/DMYJRNxi9V1R8BhSE4yXWLIkZSjdo5bs+M8YzSqt5W/bMbWHSadyqhFE5kz4H
HCpFriACyaYCqUMOUmXj4VyNc+LffbZsUXm5Azm+x6WTzJ4vLaLTUfWxTmOF/jc9
xkLn0S6zp9yV3u8u80OhfjZCHskugJAA2HliS0S5+8B4mbZZ7PZelaypoA0FbfAq
2Z4/5BzjafGYyrnHA1uug/sm4Y2j3lGNuRPx6aTIgqdr0vCQop1xObcp9SJ2Q0yB
HdHFnKOtG28sYEesOsA4lA==
>>>>>>> main
`protect end_protected