`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
YATj3kULTF7Ty4ORuRfFpnT6YIk4rUPRrM74bVTnc4GjdV8oSnW5PtQkMCLOi558
1V+/wvDfc3y0Z8//ksX8sZm3JZWtrxUppw8c14g9Y7owiwp+JumRtO1zuk5xFbe3
0MMnIxxoTKLhyRJtAxElG8sbx8N21OWDGiOk0Xyd5CqAmk9dcOIbxzMjW/wndBXi
maijUdqS+5KiRCM9+Gsp6k/iEAa2LnYTt4WtjkmDD1P5jZKsiMgFck8WOqLymplZ
ml3TTfn1UlLNm/+zD3SFGP0kABAiUT8NK2xBPQ5UzQ6sMFPd/np8iUZ5u4QLTWOZ
hTrU9OSX7lOvRUo8pJ9vPg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="BzW6NOo8eyBw+CxsNNo4wIDxODIsVe0ft0K5tGuSUZw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
DhjJh9S2BY18dG77XPz3hsiSQ73+w0XqfJhD+f+lIDHHVjOB7CfC8ieNRTexgzn1
5W+qoqOEwenoVQtit9u3XViXJSRJ0wfUC5a9axblRNyD2mUbyfH9+f59nWqGkVOh
ieHxkA/DPprM70F3APxk51m7/gNSLICSvbONgLGndWc=
`protect rights_digest_method = "sha256"
`protect end_toolblock="L7NTNW/5Dqy+2kJZXKczEa3js87UJ8H00YWI+92sDHA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 41760 )
`protect data_block
6eHODtGLmq6ccbB074dgNWpdzW45i5jL0Nzx5wwM+RA0eeOHXxEV143NNyQGmZjT
bzHAi/6AyRCB4X9z0c4MjyrZE8GF4crbMH4T59xFHqVrQ4zXCea5w0kG5yvHgpKo
rwIIbW7Xn0p+GsC0S8TZEsQ7E9zIzp3BY3ZXV9q39AgJBxyK4u2OyAlj8IGqVmqA
gpfLJXP1zjEufzKkCp6Ce+lmlzqwoBSZImi5cvoj/GHeFP1ggNk2qOPuz4hPWEC0
sktIvOleqjtxnYRShh5iX/GVPhKAfdxokeMIFAzxgTNoW13LLMhqBvTuZw8OK6rS
toGi8YB/+KzOL7BQCms43SwuYe6APpU6sYVtAvREI9jjFRh+EFg/sbMuMr30/A93
MNkwIP+6Xr8ZXEmQ8dIVRYKxAwLj3+/5fM2Gqamzv0PIQA86tfRntFX8PPIToun6
rU3jpxnO//05vkZfBS/3rkuhuhOkSIaSSPpVW75DhQHhYWEMWDkEoNX9b2VROWw7
Fqia+H729eAKQC2TVfSsTiJuKa4PKwQjM4cy331esPQcvPV5SX3P8MCryDluacHs
AG2P91uvpyj0bhIQt+7qx6FqimChrio7AnNuzku/Ryh7G4iXio1ft1eaVsDkM6NC
kFMBHMHj2GHpn5lbbOF72g8KCAoEYS1zweJpC61zp3LQbOqzcwB60qfsxfqcCIhc
09idf0FIgQZhIxf2RwgvnYKz+O+axBE9QcOAIpu0hBAGeh+7Y763jLnaAb/QlnDP
aST2o1rKlEKg/4wzQ9afusZQ4H+rB9jNoMJysx7iVX/aDfiR9ApzhwqCrV4fnrXr
YZSHn5DDhaiIW1+xuXrHyrgCfwGbZ8osI92Xar3Bn2cCyZwqiMuGpQVucssWy0oZ
EWKQyvJpkkF5xRJhRaWdu8omQ67jrZtXcqam05S409ZToi2qp99deqsg79m7aj7U
I31uW1OQVAu/Oc+kim/sQp+Wu7KKFxpSJdf89CsXDDdAgZrt92zDwmZv6YekDeTe
jYIEGoQlQkxBeW4FWMRtLhUI1fSlq3jNf5MibZRazOH3Tr/0kg3RxEjvYEouUFIa
ayaaBfGXZmeQtnoYGXQTgDnHnzycByK9sQtah1snR2r2Wdvi43uCiOwhjPJWz7/E
NpUuB0jSe3lDc82dQFOwlItRlDZXo+BUNNxtmSlZhA/e3KpNDodR+FG/aqmAMWAd
wE/vqdv8j1nzB15xPUmUaJa96wETh/nVbv7p1Bt3yYKmwDxRr1sPpgOu2GyK7HvA
LlwlzbK+65cQFH9C8R0fG+XS7QqnICRhJGXhEWqah5yn/+l4QCZnFw4jaWSl9Rzv
G4FbdcEGRLD5srpHamhX+rN5qbkNwIqeLumOuMgM8T43O3Tjbcg94zh8zuCpDDbU
zFzzaSIUaK6ufCdkEa4rLXXIFeGJsOJ1mEFWIkYaQxaSyex6cx+WMS1k8DPPYmou
cGvFoVUBlZ+4Egjwd0YGBsbm9n3wccHOq4EIrH4C1zG7bWHgb5VD7VQBgg2rT/uu
7FrsIQLkl459HVrnU61GTHdkME4PVXsGoM7ABAoJ8jcq9IWoM743OnQjknrnLIJr
JWwCPrSUSxQobJFENqbu0uLsr/aHOWHlcsA/MXK9yWK13A8hiS0jkHnIE9kiX6rT
K6ZZ/svuI+kFsbIwgQpEoE1gfU1RmDYz1f7g+CqL71oI6LnyBxLhsIMfUGTFNLZU
Tfal06TpHydVuRIFz586WbEn2Gb3ceuyik5n0wg1ep3e5u/ZUZEfOH0jTnqKbUV1
qY7PlM5VJ1pUjsBTBJNpLFtmRkJFr/vL279DsEl78/gb3dMyTSMkLwRtYsswfp2U
R2nuT7/KzG4YJJo/CMmsm5+Of9+0aniF79tT6m06sl3u6pmmJpmUNNhXrd+Yctys
IxYCifdBJUkgkF0ed/Ox17kyxVrPKfHlYV0giEHJHBIZiiWFuoI7y0NBXyg+GxG1
pSBCATkrDMwaff7F851tcH5VHJQ0LEBAC08UWXv+VOZDxkG7GTyO8hcNSLXKc7lh
F/cLf8WpONaCYTsiAVedcxx5HpGKNc8iLoMmE9fi4PNeJnqYKzMVuha8pULlIVAM
HWTmYhYgySuHi9GFBsiQ6jOpyZb3a67ZE6LJrRqDcjVAT155U7eKwv08BdspKkAB
IczkwYpruR7QHvpcjTBlzaL7bncmwI99SNXqzh3vg73xeeoqq9o7WIeUIDFVX4Py
m1Xl9XEsXGLBZM7ZXFMxX3MTrjL+2IZ45PEZgXOlYXyutbhe5zavhXlsckg39ulC
zRDzcEsJ6v3ZZIonzRLFywGdKBDbql0KYyWuqXhFFQGiQtrUWHiRmhonFLTkIwz5
X4MmD0ezaN0X6jn3+KQ/EX2Bokcbz9Ayx+mOwJeB4upjMb1AskYj5P2gaT1f46mc
wsAEjQPLKYUS0iO2xedh4J1Mt+zERJ4MDFk1Tg+uPgoMhP50HcZAAlaUbF+84USk
Qd22PJBfTjorYA10Z/K9Plz+Jde+YRQ7FtGdNoLgElgzmSzhc5Cjt+9y6lOmPtzp
FtKGiM1ldPqBnLNQDmWhFECh/WpoBMACipn8JF7YvdKYlBHA7NT/gdb+abzL2Mzb
Bs2L4u+69RuDBuBJaNkSzopSpydbLVwZ3RYn0hkmI26X27+9KMy7GeEqYFnckMVT
ypyRGxtriFlUF8gEyjb5lJvt8/EmWKQbElXx+Gz6MX4yMeq5oBfuXXdkeA4SKLWv
pwmViuGcpKR85GyJchk9IgirQF5b6dYom7rzu93bMyVYe4Cnndl5m5TnL6Sd8A7Z
jszlQgrEqaCbg8M2sNQf7LD+Ng0i/THb3TC2Jpef268XoBsKfNhiWI1dqcDRIB+U
WbD8l28XbqebhV2zaH/n3GUDKXcHxkzAwTuBtiB3hJiy0KwqzmlLo93pNkLKik3O
h4GWQM/vsQ5nOVevKxsv8lRi/4AcZjSDUM6Wai/XIimBL6k5l8LTnx/rnQGQcMi/
k3jTEhRQBgYpWBa14r3TpsdSYant4VNiBXC1Yv2LHmIjFQpOVZ3TTc8y6G4qNXFr
G0rkQguW9Q3O3QgqybwEyK537Eal200DHD/E2GQmFRsXaDSbgdMpDitLDdKDY2Iu
cd0LCw24VxKkXVezoOG5JMefnIOcy5zR4g4a2MDG49qDuGS9yEgpWGW23o8q/580
+XPrFIsBGRnvw+SnX3u2at6xPynBMC+ldQkMuIr1OSnjYKd5uhIS1dOBiAGvOcex
4c3dNnGmsEMxwS4h5ljFqjBt5ZPYwYIgX4uIpT5UozJ5Ty3KdOjLHvmPhGqK83Tf
AVwtYjz0D1PjyCojx/4O9oHVpb5Ha9RFELofo9+oUxXRwOxHwuIRlDbv7M2Uhlm+
qL0xcsYjTLeiFA6dsy4OKnp81n5NdxlvwmA7qF/X1F4hHoUvGN5WVoxQ5UJfZ6cS
0F1njDLWMaCVtCWlle9iNYONVWDPheXtSYYy9NYxkAbIt7zqYStYEsCtQsu05Hko
21Q49lrVogDQMfQ3HdAArA2i8o+afX4xbIX8r+xiogsOGSr3tLpmIifGkrwoOAbu
JwrWnaRtBwhGSIgitnAsiJ9sfeEAcUQCRhtGW5Cb/I5wYCoPTsU21bg0OXvLt+B3
0RzCVa0SNz3KH0Pdd6Ce2skGuKayzV666pq3+om6z6rlvG4KZlDHqJY+GbaZ0nyN
lTjhWLyZEO/uYrg+8LmCQbTA0rhLzWRhvW9yPyLYyjYFvAVI/Hmdj4Wlg2iXQ+Qi
VKcdMWxFFku1yoDlUtU4XeY3WMJCsnjAijRkXgjxAXcVj7sY2aukHMKqZZ8C+eC0
cVhAdcts3YG1KGClzW8/eQPrirOTHCQX9cozAzkmNjCCqY/73Z+lDKRGJEcO3tfL
1fAtWwzHviOcGi06zKHzYT+yiQwHa7EulkpReL9dzIpSDjYqmk15Oo+xxH/GPzxV
XtusVNyKS1way//MrES5NhkuiOMJKM+ls+ucq0jSquGba1+nR4O2ej2RAJoH/NH7
0rny1TDtGnCpxKNR3DBhFTjKETnwE6OlQOfsFcoBouyfGcXR9iDrehDq7rzbEdLm
S5JwvqFFIDDAqxAPv1P8pkti6NRWfxyT1Y4sBZhOZn5fng0LcjLr9b331RFznkbi
ekNJNCuL1dQMSAcmFjwTa7Zmf7Ac3oqUWzhxHNoY6NmD09qenCeDFRPTkmVBPdC6
EnjoekZ3Jv/ltabzdNTIbg/RIc8glNqXZ/1Fh2+xptj5buC+YNyW/QghpM5CoJyx
KVA7f9gw7uUAAFzhh8SQsqC1j64eXLRkM7LO6VjdxGK3FDpCqGZO2nji1Iwnhuw+
0cU3+BFWzBj8MQk8aDgO5nrsQ8CiQh5aDWLBgkhuKLF9wW73jZ/0yku3GAT10+aE
PAZW4vN/c4maKcTRMj9AhM4cPaSn/NweRR9VehqbZQjPLmSEmhiFu+0grw6Eb5eS
PCqxy6eU4ZwX3wHb5a6gCKvrA3nMlyyx6q6fjOnUYHvd2r//rpLQ0XD3kKuuHwFi
VHuiy067WE3iY/Mgze2K7pUJclphkH0RuA2tsjppnDjBSJMdXy4RumPv+6E7jKl7
NB9AN+vC8IFiDeWwNSr5UpsKB2zKofNZp/QvyZPTXUF6oDPUGmqjR0J9d49d6K6Y
mIHZDRsmuKwFOnW6D/vKEq4xG1MVIyAFYGtis3K32MY+WCxWNESIr3yfZmULNInk
mFntKBliz85PwF6/6YAZDFZwcGodjXzHvuggRMrWSXr85SqSL03qQq5uAyHxOkUF
5mrMSncqfKccalVp7tT8gGt1ZZBWkSgycvqlZ9XgKFO/KHeIpbY1b2fgi4+2rhin
/gBMkEDs5aLCPzKWogDkrGJLpnU0F/T4wkSXgJeDpC+95p+0sQzcnEfPCntg2QMs
QUr6ye5PC4x3LuA6+P6/vTPQpnSCJ4DmZ+sOZFmvHjthd0E1G7gWM+Eh5iYB5v/0
lQ9uOxvGI2cLU9IYe/QNQ22wN4Wf2KhSfg+7HTyIBgLDQ2v2N9S6oQQQubtD+fMo
xtr7choALdkW7V/9ZCdyYJF9Bnmkf9WqMY6bBCcH8jBSIgc/UAgEb/P77wLxCQYj
wOggGCqXSjKGUaUqZ08QDAPZ1cQqJitDoDiXrr1Ekbi8qKO1nbQKHe4eIRjOgKVa
0q2k5V+F8loVfJ13YOnuVbxACwsBFJHodK34MYdChQ70WiNVnAiJagdWkaHs4Wlg
QE1tU6Hu8cjFaPI7PI3O05XiyHekY0NjWvs+gGFxTQJJQ9BdFI6gm3J07YF6kBzQ
CRtne3Na3WPWgb1q4YvymGAtmOg3RXj4H6hY7HOrqztc9SpgqGQqj6IKSIIvcZCo
8PhKjdbCEtf2Z8JQSCJvPRUcJqj+Q33QgQoUKUlGGEjJYZlKbSfX4m398aaRpl5n
MyZx5zKqx9LgruwT3MTCwQadSQpZcIImqfyJp5qo8bbaFgNt29JRCqCPMQPyfw8z
ylX2BecawImxBGpcGYGonO0SWOjTqi9rtvd0hgMCk1MaUEDQxdDc0FPq3ljZKegj
a0cPAkEcdVTEWQFhfl+hXXPVmR0qGfHjMDGqM2knQHFguQrrTwEIFPilLVnoJPYc
gjT0UonXo3XtpPSgcnkwFXOcDFZw2gBx9fGiWzve26hAdaP0+D/2uMtJTX3ynHgB
4tj54v1huPN2LRjxbs65XflKZ39xEDusFTfAUa6eZwJjMzWxwmUFa+chWc+QtN0W
XaoAgIfutatrWZ6z24VjyHLP7x8Meokjnkil2dHT65clqVSHTyT9ulXbgUAKopx2
BIvVs1MsXLQk3F5/uWdmyedvpcNJ3Ltmku9M7sHCHRR2hoEAj2jSOvTxZxDO5mod
zls6vVEo9XZbw3NHjI2OgtowAsQvxV0XxAAJHGhxZeoH6aC3WqwbA2N/gVj3vfWk
/hTj4ENh212b8K5TFFEPiwsg4nM6KideFiWVY2XVe15aWhSXHRcIPdXAjLeW173M
hRq/xLCyjB1A/jMfS+XCiskLXYhZysebrHEU9OMwAgpjlosh4mZDzZDFToYmlGmB
DNuZw7NghBIUu65Z3dDmYCKHIl2v40fhrdzMGuPLdMtjNYqJAN99pbBixST+Oq/9
KZ7d2yLuLRY9iyu7QhoZTtADT0zuzWw0Yry4K5T4t/RnPHjAau3QsnkpKYDtFJO4
eFjHjtu7u/2Ls8GNz8siOwDU9uzCa0+mBKxLG8eKyeXsG3CkFVdauq4yrJwWW92G
HPdukgnvTP5ig5mC0Ld7i9CSL5wLDxmS5jlUuv4CG4CWHT0y1CX6MHP70x6VkxoR
mb2aYSTL7yJF2CObKEIjqWL6CnCy+1wyerdeX1jTSlriQ5L8R8ifOY3rJ/oMYB9j
P6TicTIkzTccsqXt7U1KeaKYgl1/VOnFOIUYOu+9FAL2kn8U/xQ8TufGzLs21v15
Fta1bbsr+IFVbyynGzUXHccelbONOeOJ1nykXQ79bfQERwzT02aDys8xhuvQcAlG
MvR4zNS1udUJHLMb5zPzDNlQgUkGpOiHqGd8UXVGsTpj5rI68uBM6PokVzpn4DtV
0ZYfj/ZzySEjv34pbMlZJtnsWKzhZPKK+/SL8JRnaior/hrGu2wcRG5Ga4ctqyW/
Rs139Tu8SNsUaGPFE+gBA+tt3JLANB6fhF+EiuC21Ea6/UHEaoUVKliyo+HcGfb5
BHC/7q9n/4z9q3a9nOfdbEEDShq9xhLvUc4+ToChpNTtk2y4mhN04iRzl0i0WkQq
FPE5SRCAuHzt42RrLMTwforg47RfJSmOdHGiCa86y1vYfzXIOwYgo+vUa9Btvik2
nrwF9bNCazLLMLxubYRoWK8hIN8Vmref2kOJdvrqeoitMPbNPKU2/4vmeJjLLyX8
9aocUagzIjJ4I9IuACpk9xjGUlsh2eYbARf51SuV9nX8P0J6CSgR9ySrWkIY5QVb
nuJkrso0lssx2u2xLgUFtlBqeiHHNj324AuZHLkGZ4CXuyPaopfe3+zFnWyemrx9
EjCz/ld2/g3kwRwRgKL7w6CRTQq/Yx1rcHs/oy37beJw19u1bDGTXldlDuQz2Qjb
MHaBhxdfGuzKfa1oV0dqXTahhYO71JJM69esus00+WePXNM1IChNVnLt+xkDOIZU
g2fIkmazK+qZynVL8Cf4XLBO6IHRndMgh6vJsg+11r8sppaILnGz2S/Y5agHZ0Rj
/tI8hN6DZPPX4fqKu5Du6Lzd83J9LgWDhrspA42g2anSJGRVldSekXrB6jgv9niZ
DezBL7Y1KuhHZz88q4J1o9bOFO2YJfmVWVfDx+eESHJjxM/u8Z1St0G2zQY6X2yN
YvxX2njLLpmjdoCnLMDG799FW4X+MsapJMSVz7b/Y0Jtqr/qfhR9Hts8pORL4b7F
f/0+p8iDGI/2OMfF/g/vt6FtS4jwqH2PYGmc9DV/RetzS/rNyicXYHyIrs7oUjv7
J/QNz8KWyN2mP/LL1tqKje2kqS+H+vY43KMxicxqbS8pnfBLawRuly8sywclYSGt
Ovlya6yZNhO8UNi2fPlIMMuBFZkzCVh8jKIVGUWB77d5+JAiEYgfNZ3zDDK6H5NO
APQzEZ6jEuXH4rjiBqlDUlt2mFMoh2mtX/qun7RmmyCI59x7kUpF3yBeDneCz5Nq
VkPZA28uTM7KdJnd1cpmec9Szel5S22FfAa/1TAuNLDn+kW757Vj35ficdbly843
/egZQ9Pl2QY/+Xjc/tSp/OvGNlPz2E0i34xhNm5T5zUhdYcph3LX07S2kk+kCWS+
Acl6jimv24yuJNc33zwur8dwn0VARlQVPOeNdFyZ2l0QQYB7G+qg2FWi/OpAn5x2
3eo9EB/fn5CtR7darZyFIOekJlnKCAI1FbhD0zW2de8HlvPTtQ1NqwHEfJP35EtQ
RRRlqUs0EmHFXLky4YkrfaxbuLIIk+EIttR29QEIwFwIqP9b0nGWcV9B4/Dh0qv1
+T3UvwAJzQdXJWdYgjbSEf4ypOG28k8VQ+igHX8zAW3fvZ8YYaJq0Q5yu0JUqvrD
QnCeLGYg/d/YmNVCO3FPYfBWkoF54bTwYqrNHTjkyJKBUi9E/sRzWqmoCpjIw2Db
okiZT1ioXkwdMEBQg66+Dm3xWQmUbjhjTy+DBosKI20AEQNGhdEfBZsm+0ELI2fp
PCvJRXHTMeLK0ZtEbwuEKiMrreGWWdrx3B4eZPn77VX4rkx4WIK7hOd6F5VEYiNb
IejAqphnm7g4I7mVHZNGgCAx/iLoneDt9r8BTN1veT3LHS0XnLQ7gnnyEVRwVUEx
rn7dGcD7qoSxbb6sDyD+X5UrqNRPJpVQSFTa5G4+Hsqqrc+RsxkOJWuTSoTlAHA8
upV80d3D2KGJaddbYY3Ger7jx06vsE/kRj6NB4wQclkT0r45uN6RKDwNmSWcL/Jl
hvkeh/p0o56SLsz9xPGw97XIfl8CQJtIzWWL+RqNjazXyQCwkln0ihaP7Y4R0LA5
3qPYAoPh8pFMwzU01OQ9nfVhkkBBqPcxf+O7rl25yPbVUPksq7lDDojcY1iXvSYu
UwxN0FBoT/keNMt3Ftq/tpthHsOzoUCg7N+lILrVoX9/fsubbjvllCWWdjc/o2Hl
THubK226aCGbD/XBXY1UYA3wUAlOeSRNwV6mPshrY5tZ8nIgKXkZCGsldxhg2ujH
MY9uU4euPTNu2PyU1xIj4EpVf3/IDL0DicfC998Z+elttrzP05nmrRRd8RYATaWG
j03fk6lKvnojq0/GrBx7XWee3myOdOEdyUgUPo8jmJ7byxlSOIAY62pDDz32alGF
p9TAbNk/0WdC+13YB3LuQ7er+oXBUpUR0Hwlw+QR81ax8GEzuDL3R1OspM9C8RoR
TBAy9s2KMCdGquZEbp6nQsQLy/fEQvXKKqRmNu2ZxRx1+1Hwdc5MT8dOQUGytYA+
GJZjez9UQ3lpBmDhxK92XgdnD9Ey01Lt6niYYKbVL0TMy4XN9RCPIWOjrpONm0S5
3yNvPXF6g/7gRss6YJtw3CwwpHEY++NiH4iX+Ob5zUwn09ST6ZiofUzCy/H3R6yN
xfYir2ZMtx03iYeoo5/1bCRKzuH+Z1SGkarIlYFnpdg1t4JQal0y5a5RRPbx9NSr
MzhN81KQbxX8sHEmRztdCebp5dNNYZgCVUoqMa2aftN/drTiBNP2dw2xeiO0h2zp
Bq0HIcsQHx8odrJKOhyFzABHsb/9ZSvy8IpqIU3AFaWmnEgLN1KKIWd7djz+Fy7v
mb2hDpTPbkIm1ej37V8SPxTCChtkCOJ/B3TNtbvrZnOxv0K8P/EYnctemxdBU2Sd
lysVrxmPqjtdq4guAbV/Dh2Jka+sY3M3XTfiHUhC7RqMUkQP4npOzR0jQVoqts1O
FM37knFpVMIP0rsf4+NqOqlQ5TY0FAT3xveGZXlgojbsvyvrVKLaIacjf8BmVj5A
jL5M1s3qSa5zhkWJbtvBcOtQjf27Re+EXVRWAi7ZrymJH6O1SD2RVxoS4F0grNgL
ahI5ghi9YPt1PjA7aPVOK4gZj9cCPJM71Q84BGajv0vnBh1v/4slMrrLqnkO/9Hh
BH7ies3EFirnyOYLQvyAMFIBdbYPp+bxnVlhwxh9zHIWS7IZBySne4x96K9IfvGO
OMVqmUxlpTXDhZ68R1jhWAbv5GwGmhH0vUen0WPc7q8SPnlPNVisN02hbvxHv5N4
h1SWtlXXpZQpy4Z6iFaiUVuFb/KwjCipyOj1cHFgPwErgwcsXaJ9xIgRLDK/WI29
358VLqsV2MLAGZfeyAnDMrHw/CEf1m4QSImFu0RPwkiGVUI8bzzr3ZS2nWhDceCW
1JhuhcdLdopOwXSgMvGsNo5mmXsEuApKbKE6SFk9ykMxfBovyjyqAkDp3CeilhDy
5iqAfJEi6aK1C0ummaaXFxoYKWgjYwiqSSvZqkQX62mriDwO3ZDHdvPfEiqx6Xp3
APqrvYPNpf/ckBMOKlxOMpvSj2VkrTQgSYDxDPc2vsi00nQ943WHsyB4TlJJnIb0
tumBb36KOtFM7OIjfSf5/0KhGFYJmz1BItIfRy55UG58sMXiRgHzTMAL15rRF/gf
bTL3tO668o2R7OGJMl5desMvJcOX9nT67oqkT6hV+FMgT112b2yDbL1B/SY2Wykt
5ftE+VwtP75UvjlcLkz/5foM8SbmYxmIm/TiVsIMKTUUCvX0o9pMokSRrgcq2dD0
wnoJmtGHz5weyyrdEDW1mouWzEbewtp0ysi49tInZUtNbYl6GIocLQvfxmT7gGZ7
1y6w/xgngN/4nFNr5RLTF6BaDai+bw75+hJ1m76WWIz6zU1uoQWx6GJCgllpM8vq
JPgeyw8hx4NOvI0v1qaAQP0McPx5SOz4rJ8voHHKxcO4DWZSbsWrKfeWsTZjslH2
oclWI4t020pGJmgR4IutxZDGJ5jRbUvNeUUM9hvXZhaTNbkLRRwjQVrxaowbhoZQ
Sz6HTxEcwBE1cx3Oj3RiI049NqHY/6LUKwEyfgEXGHSxdxkRI3JhLN2FkR+WEIlA
YWwcHU7QrvEubxbYUNfDnVrMkzxve5g6/qlXE/aedZVND9daPM8AqMglw2GVv6YS
xbF/KeYpmY9p9rS4nb1vQ1R+2XCyHTXn/U1D8+Clxtrrqft2eytc67lon4+UdAo6
grLgM7B9dTRV+1gs246N37HN0S2A7GN5PZ3Sv89wY+AF307cTW/DkA9P2pIZy1V2
/oqVE+4MeAC6GoG1doGFPecbscw1KpQ6Z+yFMkSJ5/8rjhyRquTRJpU0yL80RSpO
39R6igbmdIpyF3nsq6xHeGIuJku0/r+GFUs6g/wuXGhPnb4gH7StTlX7zg3848Sy
CQkz+35ZOrJNZddRIpv2h1O6Rkk3cMYlO610Axsl9xAx/FSncWfbAi5F8ZofFEqw
bbpPU5f8By3WOwQWXE5XQUtAeJLmnPeXs5EoimqFmHs1zwZVy6Yoj5BO+m++XI2C
IFyFkhkMLl5HtvWn5yI+jUBmJDaHePwtWs3t7gLb1772YVDUrKhWK0SWePAzZS57
ofiYzNBtwNqtfZJxMUHGAftG2Om67stQA3UMti6VOWWal+6adq6uMUPLN1jYvQon
Dc1McKT8RM2RgSGL/SUXvJ+56zTID+WFQHu8xsvfVleqM+JUx8kylF5BS+9BGZCl
O0i83PJz+FreURQ3XF+sKrNQPhZyDkiXr+822OPuZCZxijP4aC6w2nOv5F47TH49
Ml6Rrz2SY0ZJWCZYeu+rDNjYlECk+uiH8FngXUY0PNvaSuYTwWD8rOBYhKEMLtCI
PCDuvzcRRQHhTIhAizWO43zvq8TKxXY54e21SJ7eyWg7Wl6RmDQ8MYN4SCqrz2hN
sU3k59j+lZrUT9w1+T0lCIbb+WsTCuG/petHjTbKpPonmWDLtKIcoDtQl29yPy8E
5/cdoQcShTukW/WtYS+G2sRIvvl9493XGqI5Fft4t/xYj7aCTbEyyK1njje38RRm
5GpUNc66fZB18IfM/a4t9Vq9Tz9l4BrBXvwCj6+sa9KpgZ1AWe1VHemR1Yn6rLEz
KzPXNZDalE/brpQeqfhUSOrKRrQ+vsJnr6pohK3GldE0I+QOj8DwNE8/pLg4erb0
XPBBo+IxDrX5Y4G221PTOCaYH+iD1FLtb7cgY6zKoug2XgujTQw9gGE00dv7eO9z
IwnXCRUxtS1qb5r34hjbiC/06KeH2e/uwn+Gnz/6OactMca45QP0iSSkrZGKugBt
P0azIYrdFxbfHv8vea20jPZvDLuNCXmUYVHf4boKkqEFVyetAuvGP4bstTlCKxUn
cPhQV15snAPE0BFRVFrlAOKv+TdSQ4hNgrM2vzUSb8GtvhmN3z1Gbdm8KC67RPBk
SYvjPz6TSCqNvH2Mtlhb6DjN15dpK4D45/MriHy+lFQRMVAITt6sn94KsBvMrnTa
3yVM9h259Q/B5UusVY1V4wKcRXlyY46A5ND78CcjPDKegtxmImB6XeUqOrhq1Ac+
Ixn73cJOoRnatMAhAUY2uJK9e5T49/XlYGhFm7CJHBAfZ97eE/WJ4Hvxd+FoR2ym
oYID+6FTpJGUiIEEH/QIaccaZ+7HPLAcwnofw+B9jPZvajsxF2ClNraV8u6dHZht
zIQvZ5l8liV8w3EJEf8vk7EOyakIXBazcrNeJFGBBTU1uSecbDzDBFyMIkA9LEVL
Q5DQRYmSRYsXgYen2+IN3N1P1UxXJTQe5fnSqBzxWMSOK/bjcPqroQKX7Huo12vd
2nCiJTWeR0KnUU6RfcEFsbBtH+bOxcwaZLA47A6jTiLU3yiu6tZz7ipr4NO6gYfJ
EAMq2tXI51giS8NZKRuT0H1jMzNezEKK7PL0C7z6hmWz/HWcD+D1tYnOQzgdwXNb
nEwwaaW8NzOOVoJkg2OKKxxgsYaUx5e+8hIGX+KYw/kvKoDlD3uNBlDWyqINceFf
OV418vMRg5++8GMwRFcd3J7tU/1/5w1SFL3JdA9HJapl95vgsDgoiq6iPROOvIeY
BtYv5Oe2Jhs8Cla56UGpyQ9nUY5wrrAw6VWr4FtM6iVxQH0+0psoNTKmIcWGl4Dr
Bqq1JG4yBksBIjxaGN9V7/l1rWDMKyqLZfFKbV4DuF7MOXVUWjqKcFFeZBSTNyHw
IX1MQJnf2ofXsitZpuL2dppLknds6Rc+w5P1QwMLeZjvICmynz3hUtTy9/d3bn7x
M3SeXgWKfx1izCBpvtKkVpRwx1lZZ4qjpoMi2Ukoe067tt9VLLdzZ3cQ4m0fBTXL
v3EEMQpTa2gl5N3phGxwun2dYO/4AcbRcZwrfU3ZD8A2moy0Ndql/viMGhBlYX8U
OezHr68mmrx8/gc/kNmhdOAgiS9e9ocrd/cPHhRJpcCEQ5mfow/l5H528eFjdUh2
ajbvcXwphWv/1MIeITkUQK7JYf59JZCILJ3cgRglrFdWOMOhbvHOd28bUbf9s/Ny
xOZ0K6PHyVWh9dSb9oAF6yZ2ge4GNExsOGArlGmDpMZ5ppD7D/H7jjjUvlXRULiE
rw0VNxTZsP2ffbAdCMcYP8WKsDteccOgnpTkUUHY2Gw7py/WMxND/Ttm+GvOQN+d
S+I+qK23QsbgFOuEs38bqDAMeGA7iAQQWfk1dW6RhXQnyY3T5ck+j5zAFmXqjCCj
k1sDYkN/lcQ3W0E4WQ+ssxvfrBY0Xw+nkO7lOVLqg+P4LNJI/vVtC8Hnbijsayrp
EQh2hXllaRCd3yuKp06r84GI+9AIW1BRoe47mARk/WcUYYyd2/QxrD+n2iy9dVgI
VflRIfxJMFvvigUbLdzr4P2jYDbAfUGAMVCVocIl/p56yj7r+gKJ5KS+hxdDJPV3
okZoX0+ZA5781UXlRp0i+n94xt6Tdu+c8QGpV+VCeJGgiQX0byBdN42E/NPE7KP4
FDBkn9ALczyUgfMyqh6jPdVAOYLuKs9njzK99v2OtdvYJyF2+n0dGOIiLtCA93M8
Pu7w3TFAkyQ9CZAmIKSe0jTgjG30/70d5vd6qcvg+ktO5LwDyfb0U99fX5YTrBRG
UgH34u/zN70bKGuLp3rmkETypxigKo92eQiGJGMsj2VWYdR8G8dTx79ZG3CT1jOS
GHyy7KYsIR9ZbFOvu7jdiV75WUIOaaFeK100YmgOZZlfBzAQ8OUTUIQrpWR/Drqi
BaFsI4MhBs9ZAQKdRAYOcNGF3RSZ0iH8OKNkKveA1Qx1xoKTwhjA+EQOT9ZqOjQ8
83NhacuzLsXAg+f2TyDWqUwbh7rr1Cj1qGkyNtB5Wvv33NbKZTb37fJjcHQXbZjL
ObQfUFEaPK0jHjvtfOUc7y6+vorB54AxkQRn9iJU2D00eCcep+AEii3CyyiaUeAw
roXelOJf0ePnzDRgzg7ezlNBCrkBsw3Q4M92BT4H9hEA2pIzLZbtKC8C+G7jf8M7
0BuZlipbiaQy4rh5+6AMi/dFQbOLpf+JjyFydAdun8y4g9zLY1HgGNzZwS6V2DD7
TXJaocoL/Goz2AsJ+1z7ceL2ZJm+h3ilxd2I5FeFkt6bKkRi3vUIe5Cu1nkMm2Mz
iuBkRruMl8OEOUC9LT51WV1FJ+aFs44xHR2HVAOf/eXXYoYdTzLS9OtjrMem8Nk/
EPkdvp7M0XvDFkIVB2qmJ2mxfEDReJ7chN5SP2oPya9leKyY0sxNxvkdriEkGGZl
hrKD3sU1jYw0ICurAmq2TMF2ZpossoZyzjQKAzyTIG6uA56psBm5yvz6aUU3QYDO
yZl8D686KT7r39YvtUiEv0m235Gxvr7FBglSds9W4/37of+P9A57PRTRb2MN7EYu
aYAlqMpRrNJROOBLWegyvt+aRsAN2wearVHSg7SH0plMHTg7oZ7sZXtYZnnnagB4
PE4ko/6D27HZqZFzC9CQQdZ7RxuxbuNy41sPR2FCFCSf51YnqjggNDmSijwJxrNY
Cj7TKJBYWy4LImJRK1NaGEEWhW5b6BgjaY9aAvUKgIYU/ixv4XItOnQeo76H/ePA
1nRoFEUhRPbHVTh9HxLBgXGOREWGQbPYtjKEIN0eBbmHCnDVoSfUagSbWYg/Hpcw
79iJr6X0ea7xnosGOWHvs6UOLcJqbYCAtTKbR8bTaiqjqIPdA0sT7mgHyonUDQMv
2nxicnJ4na484BEbCQRDqeVybr0Gv2Gxs+uahw8npah7ejczvWVuvvUatX9tL31M
xCrwszBH5PsxrLTw+DJzb2HtodajskVuab3RkiscvDgXdFROuuec69plBM/LVHlr
od0P2t1EULqfuQDuRddy8MJQQwRRMCHSvUes0VsniMHn43yBmP1DnZqMJWAHu1+T
Gz4d6MFJO8Do0lmh/Zkl4kdk/2MY2NKQPuUfbe+RNIyE6ejH1WtaIFcBNmARKQWt
/Vv4ruRK6yOu7YTBFhLaMJSGpYYeaQPcrtVbMuKg6y597gHtCPRC6rHcFYjDRF/D
Sv4vBbfxhRy6GWV2gi2WOboqOcHLHygs1Hu5ba8NJbc3Cy3hKPodCjvxzdemS3Ry
Aip5vTCNqkBDJ/OoRvNuI9N9sTTNX0Ok+c81/7goJVIek9Jx1FNcc8OZBvw5cD5+
4/z3CRbde7UO6rZDAkxhskzx/49GPk5k0zGXfFl5LiuIh22XEv/nQ9bkvspxJCz7
DVSP/NkrmMtAgr8eL1AU+PX7VReont4eUsjkxI0oT1BJdyGreTTwQojxgsd/NAII
38JlOZ5OIJRQFB2zdVFZPVGMjvpDaT0+65836rwNPpd9ijo4WOt42GrMgZ4xd/3Z
bJ4gKcSt1p+FXCjXTJzIqzSUX5X4fTmUaJ4YNSI1AP/DkfLPA/gY1WnVyr1cvsvQ
i8HEOmciJD2BxAa/vBPJizZBnJfm/BlfK1E4Cu65Yg96Vlfe/bMGHYIahPeev/Nu
A1iN4Y64fLbG+gkgrpwCkkXHCztXVDf5BCwOd5fjzYdmrn1oTKnHikLZeR/mK6fH
vBFnXNodffwGQ+boNorsyqVRQP4epBY61Y3IKtNV3vwI88W86r8NoRZEQBay3mLh
qNLlN00RYtZw/QfZi5uRnWcFbbp81MF5A39CVE8OQ9qDn1tfScvIHNq2rz03Hknt
VJD9+vPf4k15h7ydurcy1jCQLDNlCZELUTU90KS8YZ3rLlsDT3tQluFDlZPg4yO9
uZOpCVWkOOT+M2XEbKrHfkAn7Y0R58o/iiwMJx3OTc7zxUIRvIOuBmfc1DMznqlm
hZEXNuXTDCAyDar2J1T3cIAOnpeZasmti1rkrvzOXoBwJq0V9qjSKIwta64cWXFu
NdkN6SlyGVlczvzJZuWJcI/BMNBVx+tQv4+jQYP1KlJd/FzsyENoh4JhVCiUzW/G
OqmS3po/x8L0Di4aqj/Iz21G60p03QFDuGsHj1TjHzGncrGeoCLPvtWzauBDh86f
N90J/ERX248b7vqX/3kF7QjIiJLjT7zyGEVb2x1SkdLxHlDPa6usGd5oQYAwIuYy
fuN/C3Rb60rL44AhUfTPoZJ6oS+aDRHLIffYmkRqoLu+S+lAh1XzhSOS9EdQ9Hbn
8PDoj101A3U8heFy0fka7sx4JPbBnoIgLkf5WbL9Vj0bqEUPd0jpDszSq7gEUe4I
Y8JAcApPHP9ieUVsPruRv5WX7v0npT3kej51sQ1tn+5MnRVIqZ2RY3F2BBsFMsv6
vq25lRuY75X60YWth76wqU6oJ3oQCguD6qgJfFXOkEE01hS/HKMp5fkcC0ZbA85P
gznpCWdVm+ck8JpZ4cTtmncSOKTMeknXaLE4Zufjo4WJR+lyim5N1qULEQjfAc4i
/TQkmRjKNzlvHzT13gq0QIbsX/1YKLBnOfShd9zrd1VoBzrofjvrc/BD46/hwtYt
W+REARRr0DeQq4l/RJn+kpbY7abp2S5DRWRxLbOlQmH3m7h7oN0RkckRhInK/EXR
/VOfeZpuVkFoF/xdSGiiL+c9a1AZt164n/YdoyOD9TITbXa+KX5phyTmFEJqOK4l
htRloDITdhFiWW3/UTfdynKLj7F1Y1rBDIVba37a423FC/UDCNphG3IC/fgrsGtf
hv4dHNg3xca2hwc5Allfh6TAMFA0arn+vVqtN7xNi+Ok3p3ht1SFd1UVxpzD65li
xIzQX2nr9EVJkg2OZwG/yO51aVdtZ2cItf3D7fm5EGlUBkMfKCtia9jzrIvO8cjw
Abgb6amZ7gNvSI15mvVYoGFdl/CfOTFX3zEA87sAawtQS16XAbwwzViI8/r+1AzH
SqtXzdsFxIixIhyq98sVAJAPclTfmBsFMFEzjqmwKxJftrQAKdyBI/K6KxmPQRpG
EQiwS9oH7rt0v+Q69Cw9NYnMgsG4VRv2xUycXPWixd7LQAcuP5jAVY/cVkUw2lM3
Ird6w7c14SQAUSpZGKNA8NQAyP5uzIrTyjm5jDFTAsLmgFHSfd6UEs5QHjCDb2UI
+t3PtbxS6FyKpWkEFBKpI3VnCiDWcnjhWSS6DxaquuI33Qzf24qL6R3L9k6y33nr
xZfwp8vevyAtjgtYurl2/iuWYr9y+unwNmxaSvkWM3rl6/PEtYoNtQ6yoROn7bU0
+Pqt/FtkBdGv5tPcb8e54V5Z3bPFBsOIxr5ZqAjxaT5UmKXH7rt+Opo2RIXIZqZB
IU1Tx45kSiVwEmdmPGYsK8nihMERUVt3wxVDFAs8i0sV+2n2SPVvXWsB6bsCYK8p
eX58np4QaWIl3z1QidgDjJKRCImvRw/uCEFbLZa1ZSe+J5qwaDlgHh5wZKQZ//gN
NYx0AD3DI70txL7NNtjx+zZg2Gq8wwovMw84OjF3pwYvRy+n9VT33PdPpNX7MFFf
eJYfOryAFogkHIDZ/gUv6I7sX0OKEl+fTyPQqpZu7UWmsZXpNJT2D6PmPErdr6Zh
CRm1BdeNz876F9VFDye5IuK5bZVKi9Ub2QuqSUicFCUXTgM51qCkAY0PngWalTfl
QB10/k4yxu4xQW90NFG4ueqfNxTJavs0x/nWOXdWMiWM+jDUUpzN8CGNTaxpXASS
J9lNZSLwA1Rj8H/bNPY3h0seOk1liCcDpRYk6iwtnH24fXCT+wHKWs8Y0PFZKj9y
Sv48B27gMKWCpPM8weXCzErA2oQ7AX0EXMMh3GaqRARwJvRRAL03VqcGZqO9CxKA
CPvMd4o9+LcyoTzP3wvNjHPv1c63MLOw+pPPHT1nJyP7quXcxL4I79j3w+LbkNJc
R2ERYsrrg57pRryU0OkhRdEsBUducysoTTrucJfQRT4IyVidqyTwcohval/20BNI
jWRCQ+/y8/jq6pt9BSsYw3/BYvO1af6Bs5e4aSCDuiDo5BmQ+ScFrZRG7m3Xnlh8
1c0mFn82RXmO+i2Rm2tSv1rI9mxdqPo+yzWkvZBo4j9aLQwl2RLhTvT3YNMCLVhB
Hjn5hLmOGuSPrGEbGRCdiDvIq1fhSephoI7G2pP/vaio4nGhbVy9jVc6YHAdg9rx
5GpMxxUzEf+9lQrgHdu6T29Svgw63zdgyOKtD9FcsXw66z6uHPvThzt0dI+/J2Pa
0/u8NaFSqddYSNO7SyWsumcZlWb7Vnm2K4yeO48y8g2sY/xRHNhH4LxeuDTqtYv8
BC4zcsou2q1nseCYjObnHwpwBMBze+9l5BvzKQnVpubIhCCfCdfR1FEIlDLzQ4PT
r/law/uMz+JXawNivo1zTElw97dVR5Es1yTPbdqTTUaRYhAWrWfPQlZnlJ6KZ6CP
C3UQxzRwcqrOh8ydbBZDPaUUBP3Zaa656N0AxgWOMRkx2vChEXro7jLS9pN0qiXM
vvWKW8nyFtZ87bv+tlZ0jcU9fY8I2ZmQw/sXnBK9dxcozMAMSe12WBIFjDNvg7Q8
h6VLilnd+7VjJ/3Quc/TzKPIXIqfOtNoD3pRV7A9hD7hpxlxlLTSVIjiORg+Rdto
1wmocY2vQarnL8d27Axzgm8G3KI9tzoEwxRkKAurAt9onxzMF80UFd08nQeDGIrj
XJzEIv0/ainj/zXgDYWLkFPEtzvd541VaTEx+l8KpHXAF73hSN2wvB/9KZdE9My9
63xJRkyi/AfABR1CV9/Qp0LJO5D5vRTqAEXEFExJTRIMEkz3t2VXK0SnmTIh5f04
3cdIuo5UTxtxrr039drPS5QV8slAaQImN6fjmFi9sB1CzpPLB3ymprCGKYlcStOx
LIaVsWt0scLMzUPb28iDJpg0XQNl1jtKNqQzq8hnbgy6LAvlW2mGtPTw+1gEuYsF
KOCoYJHfoO3hA5yQNDXjFdA8wOiaX4+/uwSdSo+c6T+UK70NifeUdblXKMctMNhX
yTKcMX0YbMG7azkyHQsmsE2WjrXieBECYNyxLanalojoQfh35jjeL8v7P1GmoQgD
POY83+7nPGZ/mOkiV982VU/DBjHjv68UK84DTNu747cOP6BIWODmPXP+AGR11240
ch2xPo+w9lQaF6OHI6huBR8LFiAey5UQVNrvWhCYdBIVnkSHyJj2DiIfMzBVqoyO
MftTfHNvDwEbH6aCItCxzgIV2DPOx/n/52ogmxL6rYmwl8MbspBg7m/lD916EkQC
ElxdHW+G4son27zQOB9QW96JsJ5b2WrDGcDpfjMT+G/9rMUmD2OjcPY6Dw5mB4vJ
5Wn2/BqbL59QiJVMhYOokulCkpzRU7j3kq3q855RP3rHy2rVmgbMjxFYdXOjFUtU
WJFRWgryKsqbsinHgN/AXhBPxpKKY+HR33jwM7o0sY4ssPIwtWAs4kr9eUh9J7bc
ST3ozohvPsKFNN1waPjbUCC6v/dg3LU1Hs6m9wOT4QsL/O0KQpEqq1woulc8/AcX
Hsw1vZim1G/Tt/0wBdhuqBKH71GYB9IBHnuFiYiKw0ZXV3COycoFMUEsI+1V32cu
fBHF/LMnUZG1J8EE/PCf3V5/HotnlkXUinHus55vcRei7RHbD6l7KS9Jhb159SUr
wuHJvB3cW1TsCasVE1pqMpxsJP1OL8DA41Y3KUMW9kVJnENHTia4pXXm8diP0T0R
plP1GF2cV+LmrU2SbQO74Fzfqe4pJU3yXfk9NXugSPGrwWmRI+B4qbJy2Z/uBlG0
BP7hUio8HeCFpg4N545PDuBK4Zlxs2+i86YATDVGzeJ54fl/QXqdlgQ7AShQQFNk
PU+Sr9vjuwiBfFaJ2RVOzTJdH96rcuYrV6rAfKRWXF314y70Y7KliXd2fWcLjRNb
RcMPOVlUYo31JaKPj5drp4oqxk04joEOf69KaXzKlA8QDjpU4wZVwF93rV8Z2pQx
HpehwXVntMlE3ly/O7CabkP7YRLLmvuhXAtRDF7rg64Zdf90Wa6AD6wSavEd7v8B
PTqE2qxK7dgtxhy6Rc39sjSR71LuzaFkWdBf+SDqbdVOLNVACu3PwQFd1uJ5B14u
jLTEqSvHVUz1kIHH+SW94frmB4fLO71aKn221R3tp9qo7T7YqI6g9HpUFFD43Z4Q
cou5ELYzgSfnBODABPKsRFM7Cb17Iw7n7mVko8R9nVI1yVIa/BFCS5YUla37+nMT
SXP37DC+mE3tEKIJ0IE4GfG/LTz3kcTP8OJA6RkHr9ZDEmi1904TwKent6gbdcXN
/R5rD4o+68vnGkMOq1sCU1V0G2y5mkRd5ettWXNHviGF6pGOJY2JUDmWKpxIayS7
2OINCd+yztWZE3TEpzZ/LylC62zlWA31xli0erWPUvkIm6NJUJ8wT8V7cvOQcGxi
2PssFZiRS2d9cFq652944M38uqua9zUftSJQhxLcznWzmEk38TBUiL7zV8g1p0cV
SbBQokQZaepsPoGfwWbv9JqAcp7gZ8P3XcVQhSmELto6h5S9A5wFNEhoWTw2bMZ1
pN4dj/fCBprCDMNuJH3n5w8wlnFnkiO3IAtTPWq9TaSgb27eBVwSz0KIXsTJAPcd
q+2MB7xdzN4k2MyDMipu2OpYKnJxqLAsGBc4ve7xWD2Qxz2e39Nw38LBKNzH6KDI
U60N9UBvivcKCoZhh5HLq9Z+Q9OBhyrCVZwmLhqeMeXodLAfG8TPiffzMW8j/ulq
59rbxmQxGFsf00g8k7N9RDsGbN54RgWDhNWNH3tDKSwobOGJjIAKvWnV1iiIxzs7
0IdnXNFoFDGYzRfr8dpcaScDCCV+/UabQlcpHqFwT3h+xqrxFsUeCCOrY+u8UpcL
aK4SaAr9t3Q7tLIGAhNMeFsxq6+kygsAFaUjRwENgR1XSQL2DbH68wV9DioKmrOf
mHlyvKIayslLv5GRSidiclyo425p1yDu6YOx89phxe6Rs8tP89YurOv4s7QcGeCd
hBVceR6BD2k/lfepUU1RHh4tTspEyYPl4BORY4uLFMGl1Erp6x68rqUfzCcEVCFm
vJQtEcrclScu0ZEyvEYLH8BtHzfL/sbHl57LoQYf4r4hpxFtNplyxPlDWCE1Q93Y
/gTWCBAE93oOCQcsJkEBfBxpfB8pXhTz5Zd43WJqoFQ5voFuVzIGhys+AW53rNGm
N3lTLfG9qbz3kd0LStDF+/sj844TNakHEhGV1M6+qe8dgydoKU8C9RQp+1sof8ez
FgibrxHtIuae7qam5cSNAV3+bJGky9uKkNfrveOKWCzFIOZIK1nf8b42oVqtOt9K
Hsnz6KzTQLfwM4qKd7gIgz24gAknZve0dfC2PWp6HTqHhaRqwXHGsZ28CuqgacXJ
+xTFak2YhTPKmFLycQrWgUv3kmlSHRrjwmc6Si8GiE2i2H+05cYgZpm/XNCdpQQ6
J9/StJFj32Lg4AZz1FkbzTVJXx1COufg3y5gl8uw9zaDMCJu4eSJUJfjozN7c7oS
bKZ03ph4lGfq/qCgGNoh5AbxLI2v4beCbwT8IGm25Z7afovdjuaHi+0s3teanoPL
0UukELIwYW/5vyxmIBsnb0gYZuPWVpcECE+o+sUapFSLrGvVxO5akfloiHDtet4G
6S8KNZzpLp708mZx0R/fUBGxDCE/kebc5lBjvXab0BrOxaXHrUsn6pjr7FD6caoJ
Q9c1ynABu+q7qaCI5+IKnHRqwVZHYy3m6bQ2iJLJLEn3uP+dlqEMMOpRmNueCLM3
NDPEoFXjsBBwn3Mb8oBCX3n00Rx8jg1uiQdJMSHZ+RvBYVCwjrinDyrJd70aY6ro
XBMvxDzbEAdfeTNNox35fyItYUny1Ub3nD/6qPy6sX5kFI2GovW7cBkQ9PgRljxl
F9nvR+cXR7Sldv/5+U4iuuEnguVfLQCPzL25VebETOxUZ7KoSGymd/gJkfwUlhg/
1AHYYVPmugJLnmHwX9Oapzeb9Y5mzfRbsdJP8JWZpqKoKX4znoRB7X49sFdQpyqv
JBiifEGOKbltheUIVib9ZUyoUeAQmpl5lgu8lGe37D1xcRibiROQlPpK8Tv7c0RC
EvWtNeQL9HDU74e9ALh800RbPd22A2L2ZB3eKWdpg956o1M8RdpRkIiJk7NL41x0
bURYu2Ri6a3SFuh5nBfU57NWD8TYPG6mD1F20U9uXrzk0bzgKFeXSpFDBxhy5BNC
bfsiFKcUfcuvWuSIP+zyuctzqU6AT3FKGWWaAO2u55dZivqahmCKg4XACe8ZYs0T
FPb2f6nFTa7deqhmNtdYPPXWwdK4mlGn54yMUW715M6kJPjetGXNLs/h2K6FV3wo
4/+1rNZloQbibkBIP3FZ69Ao8663+UDoQj2I365j6OdRwEbVJWPhhJ4qq+hINe6K
Iop4LP9bKq5x6KDuLjydpm0lPzXewSzHeSxK+Rt8Cg9RzMWSyqxxfKobqgp3Q2La
zzAewCzz+bieYA4ne+tONDjeTc2BpWDrE0/SNP7DOJMxxaJ8z9B7H4MuCBG7gFDC
6aehF90sSSlhPK5lrJBcbyDc63PEcDChwh9HoU1Mv6l4tT48Ys9GXk8XikEm6caQ
qdJg1zc2JK9HrW41goihe4mYgzPSgkQArnzLkAgq0ImBzrqjV4ezQjSjgkEySDYU
wV/AhBht2YMpSaMGUlIHeaWQRXrbffquLCKw7vYWqP3oV7ulOARYD5SN2IT1j53C
4Q2XtAM4NV73qJbc0MHlydzJAw21P/uo453rSmb/1xQTfFr/zo1pldelV5cPLB+Y
Tfzt1MpJ8WOMrT2F5z7XsL7zHZzpV6BC5oxbhJPhyFIsp1XfmT7ubhU8bb8YKypG
VfBKGtm4qRW7pA1rIzeFZQ6mSVJ7zj3urcBMOC0FBYTSDQVpZCB0WZhOwD+OczIQ
7UOhXPEnNHRomibGWVcqL5WPSiiLLjZbbVBU4wSP34ufoqYaMcFOjvjrZRfx1SEB
YPkiz2Rel/5LhBAauoogs64+/ftgyAtTUpfaNg6kW9rHu+d7a6ZeJR21ddQ3/Ct+
2c4zjOpy2OxydjTxzvj2QxrqRetTTWpWJeGpdRqwBtOBout6CvYUOB5ptqv7jn3Q
5sBn6KHk7eoAt2HnbAoPVW0MJrmPI1HatseWcBfpWlmViDPZqd2JBw9wG4VNsayS
uidlcc5F8vVyf8sQHk/2PLiz6iGqZ1WK0zRAaso0ln7wVobcv9ciEf6e2DnDyZ4O
aXQVXroAfpz06YGNWx5Z/WZT+Yj59kvhbXll1JC15lQu9i2+5dfI494ehnisNUL6
LV5DFzX5crsxj1N8MfgH2BtvsLfwY+it/QE204Xtxk/plO9WzgMokXY0MIPL21Tg
l1jSmvF70vgjZ3uHJ6qyyvoCLEJ02ggghYIMUJ7dvFKfQRbLJXjv8QxT2+4diPzs
4ExiSQ5EdBARMsVL9oLEsgt25vSzqI35hn6+iOIx6YrUrBjG93xMvJolkrpcJ346
2aO2+jHCGPsEK4ZsGnbpCYsm4kxJcUmJlBw158wa8Q9m6BUQure9Uh+mR3czRXeZ
DfByXU4eo7ciA9OY/nIif+nu2DX+X2/p/QbAJkMrpiE0jxzHviR0pA1/ls56ucrr
F4PwfQjwkzbg/u0GwtcWM8sVVFeODYbcfCq9y4T5dHTsl6IsQJEmJdh4T0J49d3K
TwswR5dT9xaHvbPPODF8Sphvb39FnNA2ZWzarWZRkuuuZxdYlR6SYo/JOptW/EL/
Ssiy0+hsrml06ZExJi3XxW7IcwcqK28e9/B89Oe0VaxT37doxGARvs5C7kW7pCQm
TEFymUvgT1DdUg4i6KDNh8yLYN018EP4vr6+RNCAWnClfk6Usx3+NAEeu11Eu7x4
sD38z7YOFN+UAlckVSnQ4ZLe8QmjOTuYPK67PdmHkHKeCyAfq3F1LWUKRp0fZ0xK
8sh89J5cR+dZ15VLWjM1PwUD0k7Sak/81N2qfe17tLVCyWw2SQHqlx2pbCfP9aA1
m15raPJQEhEmVD6TinN+ULHNQCqmN2XJOUqxsDzfO7f4vYOq8Ka5vIIIyRGDnaXJ
p9aVq4tg/kD2kS21txcY9WB9XbiqLvyVdlLr4jtbIQ9QLJvRuIAzE5qRBAsViL2r
gAkGtsmx6AqMjDDMcXKRgwXriqEWk56aJ93v6VdOHupEmn1RPdWKfvZCJr38sJla
Co3g5s0JkYbrudSS5bM63Jyaw9Mg5WKMRhNXXGe9RAobwUzbvVyV8VcYffTHFguX
u6hdH3ORlGO3SffW+8XCXrsjK56DfBWvpB401NZcla2f1X/fQ8BnAtf//c8A5KlV
Po9zktuk+D0a1GINdCgXvPVxOFMp2FamjVbm4RHpWAC0d/BX1/5V691SHRML7lkg
whFfFRTjz6XrYzjDgAgtQnv8ViNujuH1JAqNQZRNlBB4mTLEzLveX+jtADPHkThW
AnhJzqxbgUSx7fAQCfS9Wzwlao/RPhM0TPtOM2lKhKi6fQfpYu+nqpep2pVSQfGP
xKf3Qoi3IuhE/syAuZCYkopmFIxS89DEy7qPKNwDCfo7XClcPclbYwqzK0uRsm50
n22TiwwBT1RyeT1KGk8yo7pQZIYjuNff9NlnDWvkuEEF+qZTPlOQOkYveCXh4fQp
gfYlAo8HPbZku7ik8KxFtRhuK3cZzsd+ih08jDLFX7RkJZwBKn9w9TrAYKWZOl5Y
zoAjFmqYV1UP61c1vMSxH0mEbQIbVRsA0KOTvsKKe46jMAPja2UwbgiG2iqmJUhB
JEOlEEUw04CQUYQn4fbJ6Lk1TjVyFXz0kzonGgW4qxjZGfxAlx61PRFK95wc8vij
vFXAJfx/9cE/vmoy3DN58zghHscE7dm45Q0VEVFGlmbrgAxIHfuJLXQXqrAVb0m5
piTxGsa2JcvjpEckShpwgGFRhBNb2YLiaTTxLB7I376NqU1uOn+oppf3zshDOgq1
qnKk+Q/2g0gc9QB/gZbGRx8sWPcy3CkeF4vEa4zBDLVfLpZlkJuF4GptlWwQDm2P
ARIqTjGi7U8zuziumEPQeAhCQ4IlG5jMKesEJhQUvQKl8fNpFIG31jgZPH3qCCMB
On2BAOngvOHFM0MQy1g1VozUgwQEmvEbUAMHkDEgZgfNlREXvxVmd5/itjP7ZTWA
ySrTFlvHm0/Kad8cmPsjUi9tH0GNkVniO9PQX4MGDiN25RDyA8gzhWK2juTK9FA7
PN/CmOky1mMBZRpR43TndxZwcf+qYJztQRWuJP9RG802CWlcnduz2krburoSB8Y6
+dKGgbVs/1WpJ0GRpi4JyZ7YQf/EEzqNSOZse7NEEG1JzYKVfdhzVdgT26030kfT
Pn8YK9wz1QHbx5FnW1iYp18P/E/wAPezP8ZQbbu9xZLnt9QjI5W/wR4wPAA+n4CY
5CN+RHeRZtDLugmWQ1JrVyWggyu+9bg36KKMDDdQJNy/zMDD1BHcw/szBtajK4CK
DRf7YS843M9XOWVU+6PxfF1jYVs7jpDcpOSi1wlHdvYBWu5wotoyCnFKHCC+I7Sr
9LvFKyRdwjYWE7XDlq5OrPM+qmpxOfGylDVj3fJVk014eGbWs/IXbvGUhyT8Tltf
NQDsT+/wszJ4OlbOFkVxmt/BTnkVCmunkaVMF/Cn/Toh0AKaE1R1V9ur0LguHF3v
YS+aGKSZH25t49ZfX1B61MMESCoSdYlVJghLJGY3guBPIeasQ1Dsl8RMPv5W9f7B
lCKu4Z9p9CRKlxAHHM3P/3+OuCTvguy75piLzk5NFH/LZI4Z9+T6E4+jToUvuXpu
aOJA3Dzl3t1ZCc30064VtJukoPDlHXSBaTIyB00CcqmtUzB6UpUWXtLGVMR/9z4K
tmm6Cl00th5LVgOuAYB6+XrtrwO5/6URUGxdgDCNTCjKGmX5jFuAcaHjwMNJgCUM
3B8A8zO1JqwUJiOxH52LEmoiSzt4HduoDogx2z+EEbcmvE0zEy/ZWBrYRu41BM+H
B1FcONfK36NFUUloIwTfk6B9pJttvrx3s2Rs3Ktr/d14tgt7/CHrx42wdED0ICev
zb8y6Ly8Vw8vsH7/k4Hfb9LUKy9CzDvE8AiDsP7nU8D4fhwBD2B7xO2rMqkYM4Vl
kSOODXCyJ8lYlMIf5dCsv2uX4loApX9tufhIJ3oHew5krgVbpFHmKA+0JCgZjI+S
hPL9J5GpCeaV879kCUiyjHx3ncXiXzmeZYWIyCrBa+KSACBIXCIIGcp0L4KvD46u
uk5oHBK8lmng17sVPgLcWTdKSrBmCvCFVV/U5Y0PzUyI+s66u4nsLJfBR5opI8Cj
fqMH1LmgYM9SU2AYXv5FM5g02DKcZ66efaBv0Mgqt80eRCUc2x3Oz0ARVB6E35y9
NbP6nLuia6GeCLNmbs98ZXlpxcUl5NTDrT868gVk9hAUYbV45qQBu7t5WQSYwU+o
EK7DEBRcZlmEHoJQt0fYcAENFhDgCZsfvJEhrSxxHGw2v02cJstTBgYPgOrMFRu1
Jv70qOgfPnaqAg8Iu4ohqizLENCLlLMkceAmgKhTt+5l3PEt4XSUS8ylrK7jsNTB
RkRFX95b074IWlAzNt9xJt48XAhXllVUhFduhTuTiCmjN+YOUfeL/p198r6qipPN
yIYxgliOiqqGkG7dChO/o/edOVW8sNUalgigIsOWJh1Yey2y4LoybzG99LVyF0ME
TaSHFuFzFE2tImMGNx5tzGTWdRWzHNTfhA0gV/JYyMiN74hIpmIHFueDszATdBPB
lXqoyHYZNkWQyyEWuJFRF+QsSbj4VFfpHKhQiUz5MUppNtCxx0TMlLkh478neoqO
f/ZxRLQysyYK7EzVi+YXh0WyE7/Qjn5Gjk5QVfdGTz1eDLFFeW+wtnmxYATIGeB0
hrNsiVvp7L2euC9dyEzWTg9BT//a+O6ISID6EZVHSVJ3vsiAIuL7fMkwKh0F+6KI
2cGOejZR4CqW2VsqdHJ97DPt5h7dZR2fhGiwrjdaSwktXHR9I7q9bLHZvSop6fug
9TO8E/AhrSccLgREzgtwn8FEW80ldWy5wyFpbH3tkX97Uq8WGecM3Gnc9+8+cLpr
d2HBF7b7BimhqBEX5rhXeyXMK0eNc/hlvDSIPuG2hvSFl6knb/xjDnkpGw8WtGYF
dvwU7lJAn3S64+I/Qh/MyjaeJgZB11iJ+/STEqGnB4bbTehdf5XBBMNMJllFaWAB
xv1hrB/o5QvdzMdoSFIhDmdP7l7k/5EcJQXiNn3LYtzA8jU23ACPEOcAiAeooUol
FU5wOciV2ogfD4PVpAYDiSoODgantbmUXMiOrimAsVELV1yd0xrU97sZ8KfbTII1
HlRCKKgTmyHqG8Q6uBrukw/1VDrYk8onwfme2yRCKCh/cCuZpL1goV6HAIsrrFjD
YeG14FrXDqFoujxu6uKB3uKsXvRM2dprRFCIfM/UrHYh6VlMhVuhrEwBcCjENTV0
KewTY51OAK9hSzxo7RMUm9U0WRs0P0UR8+z2QJry1dgx6eVHTd0l4Lspty24davv
Wy9bjMxbRMGBucoHbk6ofh9ageVTYgOOkfoUcGs4cPNDXpXDdscpAf3O1g92re/5
w6p7ebvoH2nRPeTQ3SAosHCqDBREZja3mjHTSyHwBfi1KT9WIaCuAFfHIOOQ9rOd
hMdCe3oeQSH/n4akrlkLgLkVDrwiXsu3qFS0w2OjIJZO8JNwp3eTi+XKHgdW7QH3
dVe7i6kb4ARaHUc6AwXoG8RvBAtXHSpY8QaTZ0gfy4h3PDFhYGW1iununkWwjdfq
18ccMJnps1d5gomh0PwwX7UtAGvbUn9D6W440RqyV6Rsasft8jVPm7imY4pRglGB
xVApAt/+6PbkKYJ25iQ51Rb3P3oNSS0/XuBMqiOqvxXUVVUeqpOsrCR7VGWTVUxf
GkuGJ+lPKvFkIJytEHK5p7VTlJ2nXlTWKLS/J6bz9Z2qPF+u4HNWbb0ZZIctd5ue
Xpm90xwEzT7V6iEmciY2qCkXdppY4kh2sQ3ktCBfOpJg8D5dZb6ZKQiOKwE5ykBh
t+nuX6BY93akHIHsFPkAUtEv4zKmiwaV7KDwkHQTu+l22ezfGCq7KVp56cOtvd2h
DFFWDXXaZIz2p0Yh2ZvS/JqDoPHCuaH5pmU7lu9KMf1v7X2LbhcG3p3LDuJJUf+U
h7+M872yuhpdsOaQbAsQew399j+8XaEuLCMSjz7akFuimTMI9TYFFEENvgyOq7ug
4WtX1+D5Sv2z5b8FNVQmw+lqa8z23F9l/E5iQf/+U+eXHyKEE2mpQmKk3HREaA1b
eIjosp0dtBN/Xb601NnkSsk+PnUBFaYw4oqU+0cqw2aLA3OTXtvldTly2VTAE4Ai
h2zkUupm4eGJ5T/hpCwIT/qFaMIl3rdLS6pHrYEF5iKpmSUuhndGBppju0IYnPUn
CZkApVpXpyfcyLx8Ib6naPO4dG5Uv0HkgseH7iW5XrBhnHvJY5AfB0aj0oslQgmP
lv7Q5/UYC2zUFmBbp748QrbLth5DJjaVgw3qu9xgmSgeHqDcLTgtN3eu2KmHH7sh
cLAM2O1VfyLbADvmSeqCx4f7RFkl8GogDaPfzDm0V+oJXJdciqA/mjcSczZdR3Ue
Ydkmi5ptgTlLQ8bbh/EVsbsYnfuEcTOyR33OERU869xGC8D6ah1VeTpwxfJu9yiC
iEED/OZXi4EZ6lCOObdV49g1dFGlrxaygHdYEje9HW9fTNSlfoES/JHUnjO/1JtC
dxZ0ZiFrCPiGYCwfjP+7nCF09L2lU2dD4c6tgNuTY5XXANZvN6Bs7ZtEs42cfWmr
TwmF0pMsHpUVIbaYKBvKKVxRaYDbFWu+hls105SolHO2lM3xNNTg9ilkYAAnRUGh
uyLYdc8hqlig4bBbc7fU2T2kEc9aBgTeVbYzTK1h5QyNwC4ResHQ6RHpUeAvKbxn
OOyfYjV9DFknMseCDZCB89R8Ow1QTPgzrYfD5BKXQncnYYXnL9J2Y1bepbquMZVW
wcUyblicfRsz5/gxy8ARm1JaDk9vohCvWIXO/4aJoSDCXbj+M+e9SQaYQTX+0Jfq
BKRlUqbCKqoTIVF9ENyaQS3NyqLh+G21Y3IVu4pBp+1Z//xdjEJK6jUN4/QUHhln
dggYaEd3KrUIBCG9Wb4WHJq3w3+mIpziOErPB9CnlrCUXlxdp4R9JrjAfEH7Cxgn
khex8f8aKkLB6EjKLDs7wOZAUGHGXPDG/jMSsMfZKIt/RoMdu0CiatsOyAWPzECp
oRuS13guW2Ht7nNoBY3TF+2BqQ9a6cFR0356CbP/cpcGcch8yWYL+LF/0jB840e+
O9a84p8Gtin2UzRSg/o7ZBKvx/Q8IMdahxBGUviFdaEF2P3E15Vv2QbJp4VFf1YJ
w72PBRHQ8+3QYZal+UrW+Qp19WKxIkYUz40bjjv1XShz/szYPNaJ2IzVJvAxxSMR
ZQS6AXMmKsu6C2SVwlD2IKMSEiQxhU0vV843K3ei6UP+BrMjSODyO7zpKpi4xD86
ym2opMnQ5J26ehJocwlH/FcxO4ooS6mOSSwraggJdlErlTG/2p2xttG3zrN3/V5N
9oIRQ+TtDIkA+PbZxUv3H2CE0yyAxkatdYEYaf51TGBmBASr4QCFeYCk+HFIZJWG
P1leChWpj7knQYF+a4/j/prz8NVLIAAB9E9mTZQu4wXXb8a81V/L2WaGdwg9tRGG
oU6jn5LJoB+dgyxm6YnLegY9re9KnGffphg6HVLqS3cJDfTztjP7Ia6kvg6blNs1
rPPY9cLeP7wxtD+6wMUKurbuEeY5mZdErGUX0rSMTXP2mBzENFs6KaCjoeIT5Gmc
38qfxh5iwB1CziAQnxjrEaf7aE7XpralV1VzIjVpWt8PGbuZlEo38rSkJGibPiiR
rA1PWTDDE36KLwPo1e37TzEZVtnjudscEAsApRikwsex+99V8v5ANJz219LX98F5
q3DBImgNemcsX4jZvKFdQ+TGQEVsKa6Ck9PAWyH/L7bs2M+GVEPnWmh1owr4QLTl
/qxRqJ4BVXZLZhtW6l8g2yODcA/rilwsc3TpjnCRoZE+lHDkWfQ80cM8eTGBxEj5
S3f/0qOqL6knVQ78otVclr6ckkDJNj1hUevbD4ObwOXo54LTBztmsbLgWRqHWNvd
73zWie1YHFpvosXo/Yog8e9oDWWJKdOwkYxtZopwgaAXnmRbM18fSG5kPH2fqqtd
YLzmWKl61gZiJ17ZfKtTqXK+H9B7vvEb5t6Cb6U2bm2jl+83ynp2R2Hmy3YChneK
+6BTgZpUfab/egTlCPiax2SA+CVd3cecXoVvsXVHxuV5k5ctLiAvU+PnrZVBl5eh
e73qZMUSOVOAjjFw+8XK74Y5ELgb1W/3hhBLMAApkevPqn/gfIhbp5CvfrOW26F5
/yQlVMwcwxIz0puni9ukeymRctqMNQcIyPO5IE21UnilpdfdmkLB09yike6z37+H
r6e7blMdlkEUug44yALxGqRTairxIcxnHuOGrzFG3+mibraEwHAbXle2epga6Kek
LRpk9o+CBUg65t8/8eqpp2Li91y1ahxWFqm7mGwENV6HVZ6IGDsHZW1Csb8XOjvg
2A33GcfvWc3aZZ2wFEN2uY8hW//gWSEvo8s4dQa//veyw/sFSVxhu5p6+cSfvYGf
I5wgtn1E9/8G3TLhyT4mxyP658z6W6pkH85fm4RAgXVVAiH0imPxl5XBUVLRu30W
9qVY7RiUdGzF1yMonGch+mGtxM+l1ow5RZx2TfhmIGjK0oSOl1WFimzU8hDtA/i/
XrPGxNUNfbECSEXYklx7NWHPJIxvK5yZDjjVyZWb60Ifi/uKB0wwKaa0dsshBnMA
njDtEb2tMKV7HoJHz3UOva6v8lnhyKzgzhujSWl99Ua4M28d0Xo4vsb61R3rSlI0
+Xs+3qv2jTnJPP9WFPbixECTm+kRD+t2167my7evfWQT7Lt3EVW6qyvYE04VsJuA
/Ud/YPCSlc4SPH4izlxsmvoIzchHWQfhSlLYN3VkcZII7Va/A/19gsOX7LFVaBeu
Mvvj9k8WqTia2g14t3I1V2EkalngVdy8Xklk+jXTnT1IdAN4WEUk7lnFDxuHMmFa
lTceH9kEZDGStZFFeNsnquiYZqgA8QrP2O7t11y/+zud0dBIUqJUOw/+cQl+/PlX
RoCGfJjArlqylMY9RT5n2tkn01yYZGYnxb9hGFkmNZrK7lnQ3Lh7rQG2j0qVS4lg
uUXvH3AVTKppb3kcCsIK+wpD8+r2SQVlgaJ66htiS9gwQUPiIO5fexOUbRAgDMyZ
50pIOp104SINr/OJpH9PCgUNs3knG9+uPaRbWu5lj8227bCHGC0k6Ne0OCJxAy3k
FoDdCZYsx7C7gnHU3am87nL+eWEZvKK3eeeiKXzvQ+7u0pGdj63+/xAQphYXWhZY
7+T83EUxnGnrg8QhFBoEJo3pc5vit7PGUMtPm/QTceb63zrHuLUfXsGfvByMVJ9m
v9mi0AvtKFEjvQb9Ma9ISaAMCA2JDitrZNNXIWHaF9vIdLzWR7NQ0mKqCOEvxtbI
kMq9qPAi9D4o/mGxExmBMS3FMb26zRF9y7W9tMpA7xlr2BN6eWgi0oYYMZlIWF9t
5xTVRN8pjiYKbp/53ZVNonQSNEDQfcRNCG+6vAC/WzcYJFHuVcX+/f526IDaFVwI
gHQCm6xs7Xe8kT6f7BNJZ5Y5BC56lYuIOUe44XAo/SKP00aSjlcwTu+SeZOHPl0k
B6+q1dRW5YYgtBlp/jSsW4EbbXVmH8eypw43aYb/AlqewEgZG7/XidQhD5Cd+4ss
nRmBNJmLq0I5kdyDB1sC0fQYf5ay/xq83Ajy47ElXfWCTULX7pj66oc85Rkajsq5
gjL4/U3mOk41d3EGLiO46EL8vvTGbs/vYtI6zwuxrdNpmQzWihGsEGlvqUVg+oxE
Qk7Q7+DUb7i2onavL9LUTqm5bzh6f+psnbDw9KxHHc86qHyKLTInmVNh0BenVEz+
EGnZsws0hD/KKxYclS1WNXzD0/RE+ogYwuO2RhWjAuoJnIjS+dM1Vzx0vz6mMfhF
jLLOeo1WOGTIx0WjqwVck7sMxgTKb13Cbl90UPuPp+MFkvCETApBAbUMNHLWaG3F
MX1MxmumbRONxqgbmgLYOiZeeyWo+oNIqXu6PyoGcwGtQk7enbwxhMC7hDGANKiT
IxjW6WnOw37GxqDhTTidSLR/chVSYnNTE1Jt5PC2aU/Mgh6gUHAw7dKC4hLTy06S
f1asfZUXel6ePYhX/5VYkiIrhqcUuE+8k69stnUsbOrRf1PnOq8d3G0xXXySq3Re
Mdq9OHfC3ywjvpCYvBRD5t63TGfC+7I2YZBrNBooUHvFeRVNJhKY9opJF7v55n5w
HMQ5r0ylQt5GwP5BvN3JbKKwH8fNjZLotHWxiPaEQkxJhSOYurTaWAV4Q7dK0XvK
22GX7ks/rRjzqJL9FlR5/7uYFx/wh2J/gV1XddA06vUhVdrVMLeBX1jg2R+tTehc
W/rpzhrNvDk5xOkCLkTzegQFZBuP+NDAQceJ4BE6a7x0BZYyF2ugYyv5MW3JoOVC
ye8wLq4lGD16l1GXxTYvDaSVDhJP2SgAXtQyZDImQpidpqoF5ihzTbYLhkK50JJm
E2N7vNOq8q5i7nT7TxoEM+h1Yzk5/Qg4POtuQ1FQVH0Wu048fADtnL3auBReVNoF
VCkSZhmYmr6Au7mZ/a+UxbESSv7Gsv8h6YVjhoY2oZfI6Xm0fj4HaxNobc+NjAvu
5VIQ09JTQBGshVmo2BFivpLHcrg0hsGkK2e3uiU9DFc9MpwmVOe5lNObj/cfifIQ
0LJ2EqJ1g4P0kewJa3ZF++zuXRBZWiDegbNkpNPbUvSwkLOYqT98FtQfc9hFDxK+
aMUj7U7dG4ieRcY2zH9pNpdpmym4dtImDT3WxyCi8g5qaefU7hLYa/TP3eJq2DXm
dCRbSIyJU79awJdtczI8TBcttfaH5iVLjHFNdFINx1wFkDhhxScZM0fQjbr6EU7L
LDfIpvQiqnqkIWLWNdYse0757Z2fY/cjcAobv6xYri2pxL747kuWVGv8gp7qhnbO
j6fXbjQswCZWEfcO5ZhjgzzU+cwRL2WeCRF3N+VtPRlMhgS/hqCW8hrMEHyG9iXX
GdSpH2v60TXcj/+TiPHopJ7n1JmPugeWEbvaano1Vw2LXKAh3WgGDPhXZjqHL55x
tb0/Lj83RWeXsF7zD1lLMfMBb339n6Zxeqekc9/FFxOo/cizsYxFQ1vrYUjsi6v5
lycND7P7tE3MAk2kUZRndFpAasIViKUe3UiSn1QqzHwDQ/FWLzA7Oyu2n79vHJ7h
ZNUYKb2QLHrynoTDoDvFoFxJqUHkNuypPQ8c1MkdTkkbm45YBvPtmy7bMUcFuPrF
ho8lgKq+jXeqaQJeAecByDYO8My+iKdGoK+AFwAtvg+1wixuTGaH0kHt6eTWhnXd
L1xMwCgVLzhc/MmBkhVNzp6YCNabX/3ORJc7CUzYxMOtVrAp8sLLfT0snzt7ZCTP
nRPJhux6+a/Nc6jsOznD/50CqfPHJqvW4xmccN6++GvvEoM4uLW/GOtac2WY1MqT
XR4rkT54DiJUbSGaodigqWwokQN11fYEexWDmo3g0uh6AL090gdsTbPD4tnA42nu
OLYmjLLk21NI/KZCN7NmpFV2IKR2CzNk5ZGPbL+h23I4TWpc9Br3uFng5Uo1AJGI
hX4rx+vD1KvmJRtTUiXFgtViMktJP47ltufFHnYsckjvF9kR+AXyeKa6WG8/i/aS
JC0Z0gdFlbdzg6XiMm49DcRp3AeaiFaw4AAeKzs6XD6+x8Xi25WPdigby/t4d6Ln
f79gPsa+d5Ynt6/AE0D4kJuZotdBvzFB50l78Bay9/ugvLCFUr+h57MuiSiEN7rz
35bIXQ+qBV4fjyKqrlO9HH0/nsUQs4cpqLT3OjNxApiKxMtp5UE/LhkcogBJ+pWV
JGazjJMDKXklUhXgFjQiTNdysHWYebx1rTrqK6qHjn9pNwSNILCF9cl3ssoNGjfn
SvdQLPczEIBOKPAa+4HnJUa049G45vG91nRa9CbJw/JwCL8au6fWsSDw0lbjGCB7
x2KJtOuc6dvrWCgNQpvsk/yztpGeFCOe73bvYtFq3svwntLJoffmx4EsAWRLAxVj
ooPsMmGXAHJkF2FPFxWES9AFP04clEuhQvotRplCFM/ApEgq2N6PO9hkLCbG9sTi
wyJlnsGJcn90H2y0C1fGNecL5vkG8xGrNjRc9OX8Xy7nW0GP7gksUXPWV2JSsQvx
cK92s1tCdAdIFODOcZOGo2b9X9iqr1uDvNCxl5C+kG845R/twVraWgxSc8AL26LH
rB3P1tmH3HcZSiqGiKbcVHsrjZQZv2WVVjySgAbobbhwrB7c8FYjSekULGn4VwoG
2LQ/QSb3M3tbjxPZvPupmURhyChpt4XzYtKHCT5OkwQ6u8Ge+81JiBoihJrQhHLn
ePrZFY0v0OejPOFyJMtj1vCCaVWf4gNO/X/0latXIysu81s7A7xf+nzAu2Tvd4ji
1jbWQElyx1dUSL3TdqMxPWO0gw4WZpoWqmCTGSNS88muGFdeSZcRqjByZTDy6YGA
EijUELbbLNbQw5t98Veyz1eWXATZid86fMkKQDt90VCqr1raEfxbu96yqDQ4ojfp
KBXN5gIxJrEQ4vtPuqSSUTBqRaDf99yYI5HdxmKocXsajnuLNiJ5OnEw/zSKHhUO
gYwHAnUPnQ0gzDzvXONhB3YjZPDZIAk+y4TGWpTdRPrRB/LyvusJdPnGavN4JOky
ktwvdUgZ/0Dl1D91kU37GeekOYpL2ReY33eegrixwjvxgrTbFPjV5Mb5TrkEab+O
6p879fQ39lolARb5FYMW8dB1fq3yNW25U+2Ej4n+Zmfv3P1IvEX0zt9AShGiDdKA
j6xVgH6oQaqR8JzbXbCZAho+K45QZmn4P5Nx26lX59lL24u67EY2Ameba97Q3otB
0tcj5PABWSMi1OQQSYfuizwyoufry+qbGPDRiHl+ekuxNP/E5xZhpRihFyggi1u5
6vYaPexcyIX3pWkiWBcM5rbA9KSyDlwBw5ByVjNVIs435X89dA+8/BAS/ND6g/5H
in0qXquSqxErA9f5Qx5AyeKtfvCpIfpN2ycVGE2SMbILfR86iFNSwg72c+NbHZ4e
JUlwyZsDPQC0ACNNkk/FFc45htgHxcKBNcxEizfi/XdyvokPPBDHbpg0Nm9nYNKa
jPlPjJvkMuLyBmDX1pO+nFQol0KS8iTk4X2LNSHdAU0Nl8q8jaTJtFS9Zs/lx/HZ
yiVP2+GYiZ15ZM/lbgIVDXod2g8StJX3d3qg0rztcwtaR+TxZugwMx5LstnlA4qg
qWn1H5Z/Tj8K+kyKdmDEiQIU/bFcoYX4sEjkfvo3yxffDk3Gom6dYw4w1//9m+Lw
ELxOTOQQtHrwtXYzTJVn0hz+cVdf1APUTk/zoObzCrnJ2XRpg0wbDF5dSZbV3QL6
Ooj/Y5Eo64agLYs3HGcUBrUe2ek7Vg7g7IqWTl04yVA5qkFKQbtZ7gaiDuas5Z3w
Ap6fMLy3ccqJ469lba1muvgaYymK+N7yJJNs3XTODxZI+6nVflNJp1FT4tVmF7ug
yccp7If4CSyIuem5Md0BscgAPOxg6vvsvbuYiPtgAsMLT7G/ouzr43/zegnuqAEh
LTx5kN/nJ6moS9UAwsnzDY+EpVt9JSu+uTG9j2RmHQ/BQVdpcIAHIWjnOvvcxBq6
okU2ZsUFQ4D2jeIG+W5WZRhQHXGtyO7sSK8rlqSLyJBvATzgMeb5Num/eAiUJGHP
FZoJ82yuGj/3gyW7q+hPNTUszv6O83a/NXBwigq27Lz/tcdPZOKuYPGDe9X2VTM3
mVLS0ztMB64okqiacIbTQKnSyb3On4erB5NfDu4NmGduNKfQWPpj5OpPHdr1Ydcf
uYQnn0w8iE05QLHu+/6hjUNfE/fROm8uAkAs/T5Fx4hpoktfBPeNWbw2dPvBVWnn
hxBG3jrMBB+3w8qt2GAmf7cmuhumwmGvpF9b84sAjJ8n1LtCK2UsMdUeAomxt4OZ
aLWvMwSUnSFQ5ktLYaHUo/PW4Crxu5ZNnd4EOfB8VppicmV2EzTdrCG10x20lUrZ
6oBcrWVUII2lLgYi1E3ZSsW9vaM6qGE038ZE0kR4M67BTJUXNmHq0TiZFtYoqNUl
lxTHIoPv5S+MmiNVOco3OcxlEnf8jCVriSgTems+8lTEsGddAiLWVdAyZPuamg44
RbM5wZa3xsclk0I9TMgaKWHPWAsshJLTKILUoZgkvxhdVXa35oJXK3fJjVIgxb68
OjBcFVmuwWNKsCYEM+xxUH4GR6aVlYdVLOSWXWlF6SJQkrhkxt3tECqBxt1BCbCP
APjgSrL6tKBIEbspk32rfwUG3VByry8wQ0ejcNMdCimlPH6doW+wX1IGAw/Cc0SR
jpKMfPwH3ooPTmFqND2Wffh7B3q+ZmvY7FLTXeaZjDO5++LhNX6RGkEIYifcqFfb
LZuxm7hfgKBim8svOTQFq52guIvNsKYpGlzcrQD4N3nwNf2VtvXW+ZlZ0lwlLwxD
/pLmxl8tBcjc3zWpYJV6mpGePx9N2xnu2RgYOkFPZZZEADzcp3YzzQmH3NzUxl1Y
Kdq/VdPZ/AVzmU7udkvajuezwvN9I38K4q6C86pON8W7ZIkohrRJYgdkrzmVBmPn
6tjvHHkIoXfkPPs+ooLeg7ELnSOVlWAtYjD8H6nURwFN9CuDnXaZ7rmqFCfHURJ0
3Q53YGk1o4W4hDpho8pQKeHwAkEmicVFKV91EnVh6/Qgan6bEavJc71qRSamY0r2
CkbayW++moHu3z567eihdsPzeUwQ6BCSvJo3dswSD3Y8VP8gLdTkf6aSsd6hofKr
ScQGN2OI9f6ksAcstd2RZqcjPRsxNF4nf28jiOMJg0U/XSRQHKLHc9R+PtuLOfyB
kl5eKyP2SMie4rF/6v0WOOT7xf6l8uVq1OQULxDH7W3KqaRVnX574+quJe2NBC08
gFwJyrz1bNbDSvdLqjDgijJwDqgRFvGx+cwnZ0Lq+XTuQL/A6fEub24yMZGkLvqD
o5B5zh8I++R2dcYh4OBjutxfS48HUwbPWDQvzdsxXptxs93NE/jEQvWU5oTOyNzP
ZMrhAc5y2can37Z8xetPGybjjVREBiRZp5Yeu6o0hVeK+664XJsI4HzneBAt922Y
odujYB/B5pxgRjlo7tRftPscfIRVrhWPzeyQabojAsZ1ZcWparlbZSbCM0XYS3Tt
MGl2u/OwaCW6HfGLXSrgCJ+BooJqvlmBhcWuOv0acAhK42Ac6ome+y47+wWfunWW
NoWRvl+7ZDxgTxHMZwMhaR5caew2AIZece4dP5xoy+/cvH8w2/3lZLK7TbL1mvV7
foFVltqgt/LcfZsboRJ9BhPDHDXh/sZSTZmKxNtJ6FJyZch8SkUNcirDM6GUYZWJ
UvBcuKAJ6Y4eSkEpEhn7aLS/ehZ0v8okJD19Pzc8LSxlcSak20juITspKbUt1pzz
SdJa3y11c0Zs8UCxtRPGXeeNLKvrlEPG26ExIpp13CEF06JeLb+bT8bkD9qriMPw
I42W7rrxtWxp2Tdyycmh9Mp+mU3Wx0BKPv4VSSVUIwDYLNrnVh5xnIt3tMKZx1PW
YFsuJN1J7ybNMksRCa5W2rCdqlfyx3DQ2Y90nCpN1HyKnfcS90H/8mr4ZuboL/ud
GF3paNfJVbK6roLDDRmXptxHs8zNPIwwHCJQjetYKEUA/fFb5viHXKPwS9RmJcke
WJvEFro/zHo5Zv9LiE/i+NBrZhZgqdOeawrlwBHjOJF+JLK9Zgeeqfctn34sQ6Ab
DYjTUugOSL+krh3s+8hNSehRZPKULr3iNgm72nbIc1sS8q0fLnvnOfSwzUy2NKOs
egzd4V/yjx3LtSmdelUsHLsCdXqIxxjbwr0QKXfcrmI+rZJZyWKeenzZEq7yqkm3
41ms9tLEQ07FpxLVdIZ2LGSxtmS289DRrQMJxZJreflyzNCK85kMNpWWGJ9HMHsd
TFdW1WwsAxHt/aRY9H4HuVXk7Cj+5/5/vqFuxK3OSxZ/nhtBcSxyO/2Edq3GdU6N
p/h8btHhuBt+nZaohp+SuvaiVcRJZzbtVNj5tyKqcQORncB/tUeT+riX3fl4sQc4
U34dPQem8zOurWfmYeytfHeKZt5biTi8NVJ7mbSmquZkhte4Hrz76IiCRB0Fe4yp
nzO/DglLVnkTS+8xqr45vrWk0d5SIaKF4JH+YkOED340T3aKSkdkWgJBu8qOcDEJ
8iyK2j9hCv0xg/2FXQ8ENZvcrIwhBdmarjtLIdtT6qgy8kdmEU2z1EnjgcDzYPdD
0PmIAgpp5BsNAd83TRwxd0YYBZfqXqviXo7ZXealpkjzIYfc/6z6gLMEDdQSbrvc
97ooVdbYzwMOgkyHzcT2R2bF2MQH7og7F8dDA9A70gRrslRzX+USlKRYMGPZFsKG
JDGKS+tE4XHZGz7tyuPY8Z/Ukt6MaiXt0T1nwnwbEU42fiQTetM4G8eQTzS8UrvZ
N3lqztpakMGXfNLhi6R7tCio420BNgn+Cy49SBFLN/dwDX+OQo8CZqm6qOFOVR8f
EtVkTbfG6uP4IxuP40WjntEoukWMHdYL/UQ8aTfIdATlgwWqf1gNeeRlJuOSBMF9
KoZnzdv08jXvORS05cuXFwEYiqykwQMkTI7OMY85KgmS+f1MjA+mTuRxWr+pbdAo
tzPjJpvobM7Vzb0CN9dXiweze5Z0AIku9BMy8LICMA1W2ehtBEPz1jrEDnPTEZb5
XBSOGSRQZxB7mJx/8sz3Myt6yQHC4QsdshsSE5gFXQzuXzAFHyNWJuo3RD8HlXMf
z9pAxsipvjQaht1S0HLJl8gItqkBDWPfQ32yG0monVPtDqnmmWedX38B9bv/6/RS
k+VaNW4XZr5iN2+CmZetcIFiJFhCiJTZJo5vwWgGXSF8zeRhBXPw1LY4MGNltY4A
4fsRr/WUJkKUBSlSpO2U//L94kyUP2xd0TLG0y+GTRrJFrDeXEJBBR/x50JKuVyN
d13wCKbZAlphqGL9WS4wvcLvdKES/iI9z+9Emz0vvT+U0dGydnShzg9+o9EU3KhJ
Mk0AxJU4I+uIkbDWBQqIn29/JCI8cyCku7fKuyKmjNZTR2yewkDQ3V1egbMZOtrJ
2m5eO+C9zGiJl3ImaEtlmI8YNHOkaFflZqrGQYHzrnMjJJ9D7XmpPAb3YpzHPMIK
4lKMuct0iSq5jFfI7C8gpVTtM0BVq9hofHsBm6FuesuPMfgSIghRGe+/s+Q10lNu
YENtLk/phGsCOst/8EDwZRdlCXY2SG+V5K1aHRlZzw2MXBFeg8F0jARfIHqKmMOZ
hVA/zM3RZVCJh5buPdtL728cH0zYi/ZEaEWFHSghUgg8NugW7xNugf9vUusoia+/
hj3WvJU7kHKGwakhNKpN3ci8FIHI2/CR5httKE2FgO4EvUeJLqHasmVhUjCYGnZt
XgNnHLsuWLpY8ufwc30v+GR3uvaqoCJL//lQpR2655/spU40Fk9E0uEQkekujtO+
ONFeXpr7fS77CrmVtnbbVlx2OAB2KgMG/VJnpRqEeoalscRzPnSbhlA9kwEIkP5c
c0MVK7zktlHUNZJWFvjL3ONcFwrWmD1mX1tOvRXMdMAo3sHlUqPohstSJrSF6JR5
Uy+3UHLLQpoY8XMlrdEXdhA52dV2Pp89cYF4bowXvvhMrfgKddP5mbvj0AvFV4aw
dgco4bMu+wz6DN+3bviaDlkNhteeE5WQYmIUYl6Z0/gSA3fSzJJEAP9lenWJh4d2
MAekE+5/vgPfZDPjOZ6i4QQsvUoAIw9Wg9tJkWYiTmshQu73t74RpQ3rATp7p0IT
yRDxg0Jnxv8t+u00NWlluR7olbkgB7lkOGwCgjvHL53wDARQpyPf3dmeQRet9Dj2
iWWFV9HRibCnP6V3IWQdzupB6fbyYbpXzMqz51wXNXEb5TPiHyPbtYANYnDKotXA
2fwB7YuExpib4t9/0AAzD9HBXPA74MxioCmnP0QnHSkFj1Sdc9+cjievAyOYxz9y
cQdHvK65qcD+XhzncumWe0+UYR5W/BzT+ypQnj1gj9W7RXaT5otom6sR3msyHZPJ
5kesNAYkdKkOETqr5j0anI6+KiHxogWlbAztHTFjU459cGynVpHJdQ+X9OiZY+bR
N3dOcK79PA8Q+dCxplx9ybLqPuGtZJACcSlRzxQPKPX42qybyGmoc6wsfInAGflT
F8qCv7nynDSCZhvasneVfOaDERy3Dw7rbLAaz5P6s2R4S+3aa3XQCF7jNsCOGPRG
PRaotF/w1ciMF/hhnqj4QXze9mZsADpHPLLcJU1mlfaF2j3Jzl0anNnz9C7BVlC4
6r/UOEdgG2LS3JpbsNahVvqjgY2fgPdWyEdOAq+N1O2gFo+PEHUorDZcYs1dEEjY
mwyp1ecRcNsWE9di6LxgNYnj7/IV2ZSXW/qdrYwT4dNNOorO2tW2OY2aT69EZWx/
ynGKLzoYTmxKFRRYLayyk6Edt0b05haYDREG2YpKZ9Zn6aYbI+l4mPPtn6SNFE6c
uL7AfU/qkFxF8ms0YDNJmVjdDigUUsCU6jEK8NTRxg+4G3gwML3W1bkI0QsfXrCC
kRLaqKGQMl3KM4fwFP5JyXEqCVekDFDLRsoYfpzBehLbV95oWEBHY1z1NafeT06k
issbOzDLQ6WelIeUto5dX4WulJF92ESgjmDUwdyQ06gP9wHFmwotpgHNdqzUaxxy
xrCgHNqxH4k52MOgvjRYPB3xZNF4bssqWoCMCyGdoM7fOtEWDpRR/kD9eeYzkM1V
5cTqQk2dxYuDVOlqI29Gf3xzNqIICvyTU5eCxLX2tVRfgQPrj/9MR2+kahinZuWy
f7HHK1h29LF3MMvB9gTKnSFbIQpQoHO7q5/KHc7NCXTqhWnLHjUbEWSfpF16Hn3Z
qK+FgUDdRKel3Z7MzjKsjxBnoFqk+BIEzqjpIvK2PcAUY08NZWRjOLrUDga2Yrb7
DkOSt2rM0QlG4mPZDNfT2jyNS88sxKzmWzyA7ENDf/2rG+jWWj5XGGLqN/Nb5dfW
kSZJ7I8ke1OkVXXw1JEOGeOFHj3f4LKYIYlnYiKdG4EJl3Fn44A0/IUrfIEKKtry
YSm6dznDIZh9qdWwe6zFqfEHCMtUT+13qeCAvDTVmZY46e6uE25JpkdRaYRp2bbS
BwqkwycZ64kUgle/gEvqDDRdV6IumecViQ7FhZ6I3EGsk8+P/AboEtJywQI8hy+Z
wMcvrADsIOfPEDhOf+WA+mSqm2s5+bKN83cJePQ/WAyu+tmACT/fFpKebLS4KHbE
OZyYgc7tNmj+xOsjiOGobYhV4+JtO6xEHpAku2VxFBAgW10EDob4JZzBaSUzOoaT
BEf5tBRbF/7k6W/0BwXGLN1z/DNJcgRtTEyClb5scqMagKIK/mZ707kX5d0m1+v7
gb95shv+HikDOl4PCp7XJT3Xy/k81103LQzNtwtTplq29USnKXbeJTyzC4GvLEAY
m1AsLU5BwsKII0IkaJEOHuuwzocj9bddarh+TQse7L2vDVr4npJP/AsDePTqSddC
SFkuKkUONAcA8tzir2xHZwm0bR/RMScD43KW5vlpxKFyXQLpljEcOzyeWrqJ6Nic
RvwqT8Y6zMepsyQanRnC333joFZSvYi1pM4iNW+B/m2Cm+KPpkxug5z61Picj8Bp
DNUzxodYh5A4cF+A/rpV7+fcEslG7VqcoQqQOfOmoxlVWHHcWd66I6GqWzQlJ+Zq
90I8H2ROXurYJNgJvP8aUD769WZvOK0NWamSL1NJZ5FqwoC7FsrT/uhlz1cqb+z2
h+IDUNce1K8lYebavUPH3b4b4EGmykfemBXaUfi2AR/aVe28oiR16t19b1CN3ooF
mupod6r21Hgy+7S2UeHAatYQeKgzu7T0cZNSiv74hMEEthwwnrM6F9fotg6sHBX4
oU5WyP6ahRQaaISdIfrsb0AQFUrR7Q4y85fFmaK69M8NC37J/USkd1bWW1L6oRg3
TFrTASRBqwns4L0XwEG8wcdf7A/ncLGtan3Ryyt52Ql/KFIPf2IhfCsu0YVUIlS3
pQmX+YwBe2O4HDU2nSQkh76S8Z+UUYnsEPHoGu+pyt1m4gtgKqGS8AUqnXz/bnti
cyIiitqfLRF56HFZpe1kNLZvje8kxw7TkO0PpkdxixZd4QCez2q5HUadrZIzD46E
PK/C5mOI+sCjZIqysl94maaBMZrxxkUZIM/m1R+YZm94xn5uwgynSY+/X1zk1Fei
uOmVb1NPPaiZiUztos1jt64S2RSV5QW27uc4erRMDEfLioFsXLNo79dBEEix1C+i
8Y3eZEW+qNwKWhPV/KOuAe4lMosy2Hm8hsr/WfSZ20S7eCwJlBIIL+/M/nQEMq4X
5ttXDadIE/KZKdsi7+EWbi7XVjAgD4GupUYxGqhsXqgg6YN1buRsuvjnZBrv23ye
0h6CSMV2kH7XaO66z13RQK8l1s4cmuyhM6P/UqlMBdy7zgUmqJ4C0AeoAFNH4uMm
d2iQwF6ysYek8fQ02xBoep+r8vZj/78CDS6iBjx6BO+4jL4gYjnIKzVIMx6rjp0p
jRS11Jc9nbTcqgrn4VDY/zSWrt1i1vPnRsEWP6r6iZj7rrPm/Ox3fNfmTiGT1KWD
/7Cxc+Z49oycJf6YP5U+p+uW6cJjE34ojY6Z6bBYVE/Z3qoEXfeBH+W54hqzwcIp
5+8+BspTi8zNM4p3Fyxaoj29XgOJH58fB7XeRqRFnGugaZyRanX8mRlakSDsZ49p
Cx2/E+wzfO1IR+N7Tg9FTfMXl01yDpKk7QryU6IQ3p8b7aSlK7mbJJ0bscRZoqNB
ydIqYvAbYfHWQ53xlbtOZ79NqIsT+Noic+FlFW47aT3OpJ5trjBPSPpyAPXJ6v6d
T9s6nx4uo1QAEsxVyMnccuCJuEaFILCXnCL9Ftb33lJ9Jt1D2J0z4tgHlj2fs23B
sQwGBHCwllorCL9g5EEYh4uR3oOymT6QmBoHyFQDwQyBTDJuUab8EteG5rAe9BPG
LuyGZqdIly5v/30X3pxIQCfb9+/lHjRZfltzBuQJu7gLXrriQHtEZSYOmXEFGWrL
UT67ITM/FauNj4/5KZrF6s71Tu00EA0WIEKQ484oEiEcKzXm8rH7PXXic6+yUJyC
+AGknnqYSL/SIl0Yy2JCqjv6y3VnffpNNw5MNPi2qWBsF5B8RNssMBEFEgCDaUx7
oRIAW9DKooSkPG0ub+Tz7tNH+/+Q9zybUyMhA5YkSw8M6/oayBAUtsNlvIgaPz2P
DVCDPl89a6DOaIYoJqQdcpM79zr1UaRNL5SsVdq68aM8PMOjSKtBS9iAvnV2US/T
Ccq4K1fCL72QhK5s4bnLidXCPUKdHXqSMtP/9puo3Ojehmob6ROimgxOk622qW3N
ORfKn2YQHvhQhdTsvH5r8CUX/M9IpH+BNfyuMIu2z0ISOu36Cn/eJ9VvFogZ1V5s
c9Q1iK1RGO8LOwSf974fe5GvUpAiK7ENaq677fbPa8xkoRxegzoqM7VwXqxHwyIk
CUdgdpKlFzPbyC2C9FsQ2M6XdSYo8nF4TDeIlgnRQFNDzwe58J+l2Hcx5tdFGKFB
uTqKzeSQxKMSBH2DSR5pD+hqG5tbBq3PGoTfBZ4oDOkjZ8wlrOBmg2eLVJBENa1v
6lBMkGnJ+sQl4048/FElpqhFM4uRmQMSSdi3I5WvBpW/1Wwtn2InWD6DxrOZH/4r
DmVRjI7zQl1J2Lf4WJeZS6CjAG3UFOEDoWxYKy5xsgOL4079+ccdTgoie6WF2wyX
t4fv8jZK4SL1Oi/Y9WZrXR6o7PRDL+3jYVPMtCCq/i6OLJHePPqWXKtRhFV3FjnD
JyaKIroHV0MIPpZ/WJNsjSP+pYwOxBETyj8BmpMH9EAvkBABpDRH0PkXo6pKqvyC
ImKWMo3vPuFWuOwPViiBjMQJY9pcVKfIm5QXnCSOXzhmlf8BpPvaaHenAkoNc0li
1r11zp3JBoF33XbHnUmt+NFfEq8MvfVT6sppu+I3aIChSw77godHMyRyoWm8tIl+
s6bLLSjG+eQqp3FXiBl5xWIXm4TbZ18/SSd82hds5hT/VK9oD95x7qM6kaQMcmGh
HS4joaEXcqMuFssc5qfND9or+M5fHLr8dFrWbsoVsb3EF9oR+G24VIPU874z5BcL
jwu0HZp4HwQ4d9J/mNtZxZYywadyguicnndOuwWo3mLxYl/ejNJRQ8H0HqV/z21/
/A/UsNWTQY2IcnV59HoHHas/4ZzWipODxg265VvBceiVhixSc4SX9T8iDP9jgFG1
mqbM5PEPra9LcLbW1KUUpl9YVb2A8D1juvP9YlzVgvIjlU/tBqMGcUQzt5WwUBD4
Jen3ShpjCm6ocZAxe8q95Qv49JnsWC0YkO4ECbB0sxtwXr7X4Yc8km+pZsQqI0we
vgCRdfw4Ipk2UmpY7SPhl8h/qBNq1VdG255JGBl/ByQTJyrbzhgCQOcWktRFlFhp
CpGQsrNduBff83txAnjA+NOSi4KMKhk9PtylEHN4t3qY2L8gRHor4u11OpZJni8m
fVcOyVizaASNUY/s6vSDcRPGIEJEZN6IGcVaEKw4KIu79oTJcceZRtgp2V9jec9d
fdgD7Lf0kyNr2/pdzCl/0qXpD+a8G/OYglp1v1XXlmNjnZmdkDTZGNrNAWVpzGuQ
LgiYLceOfK7TaDnJRaHXcUWht58StPIcXkKY5R6KL8t6FG/UGmuc5CQth32VmE7t
VABJ/2E8pwUQBDdAXVu5h9wBumyuNsH10u0D05xMxKQtqtt0L0AuKJegt4JcFLae
5NZT3c0fwK807iT7aBe+5rCc4cBarmEB7n+n/wurPD+NxYSJStauX/eXq5SFzJzl
exKfSY80q/4faVfDEx59Cm085N7FmcXuy8dxYPAL7UHci4mwOS2oVaUNnJNFIVqL
ECkf/AtQSn6PvGg/KNyije/ZXOwykBtFsE/VdUYXPQSvJGCGHLAFChUrtTEd21bN
XEV4Ahc3I+WmMVTvqvbfdJnXVQ/H67ZXjYju88gCwZQvIG3+Wd4KlG/mpjalyArp
1kEosHAsi+J2Umas9Z8/LSxJ+EDteSxdXlhMop9fqha6ra7ionkOrpUwlq2N2tjS
FCVFu267n3HVty4k7rSE2BlJEFhoen29t80tKKIvkYK8IsyNhxRFGdr6ej2EHhf5
2PdUdycOrWDihE8wPeZgUsQpcIqoQIx907ceKXZAqvKSGjkfW0uAIQILpt1LE7Js
1oHlY8QmsbNQxjVv65rm1RpKc+Wr/nbBrrC/wv8ZfHE49fthjCGaaag/0a8Pp4D0
jXHPf5YPl9VcaJmZ4vA/cq25XteMQXyq9CCaVUcrc15wym7xoNqqp2EZmh+B0Qxp
BQjL3tGtJYgWAX8RbJbiysCu24EjX/62qopqvtGvmFSaMaiVdlqrTxELhlS7ZzwA
pyZANvvgOECm9LL1RMMhgj4KPHaMswIpqbPE+D+tELiOAxdd9yFz5GKx5B9i4H4D
FxJmMxFRhL9O2AS7sNJWvsSxFTetbxWmR1FenV4jYJSYujLwd60QDqqtsCGlQYJS
2edXEUZNr4N8z4fKaxnWr84Akb+4zXk1iIpU/PFuEesLiVDnKHvx9G/8avFcHKWO
yK9BqsTckTt4KsaqjL3o7YxbfOg9Exyt4UQmSJ+AjYnyKMYkQbkIKPBo+1tppwdH
z5RekP5SfvtobHgusuHzTBrxkXD9m8+LffiPMnz9h5G6/yyWxhul7HQDkTvEgCzM
CaPPnsg/WFxyz0eT9tUMH49p/v9+EoUuUfOxrHnLVQlicQ8JyuTi/OLm0tG5UO8u
2k4cURLF7oW0iLuEIyrBcqr25dw+o/rv5qojYok58qzQwxTQKFJdcqHuGBYifNAB
P7JjqrpfRmXZtXx0Od7CAxQonSi9nH8RguMZpCn8Gi5nNAEbhfSxYQoBGfZ8Ohz6
HPSSJU16gK+HnVsjLYdVIFPfFr5Wb+uX4b6bvgCL/7CLPgwOdLHSEFV8zPnQbzkr
X3BBcFmZse36a4104NP5K5CgB+ATn8X3vEJaU0d9brX8yt0oVGGuI1bYpiYB5EXg
/2WRRMkteJWUJmuwHfaLetpzjJr5VMsxt91nNkYEc8P2BT5590X2KG72yMPAT0dx
l1tM/s4NSRTnYfXeKcHIBKWEk2PlBgvCOkl4TSEN5FielZ0Qe04bIFWVvyhnrC7O
urD1NO/QEgriSM50wRGMeyco8QtdIbdqyY9+q/ewa68yJlY1bg06/oiFHOiHQErE
8hU6lEFU0R7FLebLsOAGbFgAN0llIuVhGgb2NcrkCJxocd5HOAKEYYwEeRibpstU
+YlavtY1LH6X5dSnfTG8eeZapJDbJ7T32mwBMFXlhSxxnRNIBfdm3T+fYX8dcUsA
lwcICDKsbJxes5D0qVPUewc9kXwCOTzgzQvDkhjMrHOhQIGJW8vYpxbyHB9PuzuC
uclXXbC+e26nJndZ5EejQ3286nuKZuEvC0WVk/BrpLFjjKiLP/v3rICrdng0587K
yjKT5tvE5A9/pXlCtt/2PXfUhDsUrEMMvPHLKdpholPFCn7dq8+XWt36X5PcVogy
5K+FjwCnsoSz/5X6+6I/CLuLJe6d/I/HHYsvANe8ZRQFz2HhbuCA11eXzusVtoa0
zu//XwJE/51cY6ejDH7nXW0Zso8DP1nDXhzSs9yiwUaeRISwkVdCZXgHcT+DFXWG
E7a5ezhZjLOJoNtQ36sRXpyQaCvxih+Qgl4njViWVA5QtP1h1kWO1eeMDqN3Rk0I
bO+yn7hrmXJHWYfFB58lbrmAH7OxOfDNmS2zn3Qgup3EjqgqKune4lhrpsemWWv1
5emHe1jqK5BXz6pchoItQg1rWUZotDu2cdrw3/e0u9wWB2hxn/4D4JTI+TKTR5Sg
3dd9Fmja8ckRf6oxiqna7T63jzMPrCDT3h3c2f4faJ6/7SNO71sLHR8nqvnobyYu
aPQQT2zdKbBi4gR59QUp/Am5rXWcgQa/UmS+NuI293kmlEsghk+FQ5ScxWrDc4rI
t0PjG9HJ30gBnLFGcQDc+wEHhSfPIqHZE+PLLNaBm7//5m6NuqGvM4Rde8aiBKpx
Aw9IP04w/ww2pPVgS+qm5tOrw97lzjPi0LJKG4ln3DxGf0O8WKLKjFjM8UuPTfuv
j/m+PHcFEfcpnyfpU9GArXJa1b13CDMutoTuoyecHBrn9LUhrF1G1KE4X6lDtXLt
TWUJM161wC/7YFi0sRPzbS0uBuDkUEcqV0q+NbWIbkErT5DikdkHX9Qc+Q1tkbDv
Gzztvy1748XJuzpCGb+2DF0TYdfRMr1Zufe7d8dAKy1kYncaJF9wkFyMjsMoZM7S
gTM1peNz6rS27NPDpt4eypQZaOdPurqaIAFELYmeSidRunUi5oYyKYAZtYZdJACp
Z+p2uxIPrGiiAat+NIMXms0ZIBRPzIvTRHcCBTMH/VqFRZQROt4xjNmqBDaF4CXd
73MWIASV6LqoypKgo36g/bdbDpBxRhyLFoVzvAy+8qqG4mdjDrr012GbBpyvbMJo
T+reQ/3mt7gsA3YodAXCqfiHVkhj36OCp0fZAXL7w42DgHNUUMYnPF6Bh/1pAdf1
84cWuWt7FDo0ymvlMZJkQrCaV/ORuO/JYY6/vIi0KmZ/Wet/GaiUZahenF7GbsJw
W/cKldjH/EnxVe9YFvWHDxU3nsa/MddbckELC2BuYnOp9d9ejDvELY/4DvWKS/25
COG0EZhbTK9qvbF4mrqZO/IoAVO+2xPwN986h8MvByXLvI0b6tiUA2ILHT5dv1Kl
bv2UED+GK+z4zFZUxnrVKjxjvQudeZHUvHpJ7dj/2q/s379LNXtyYCu7t7DEkpzC
ZqMZHUtMfLvTwFkvWGbz96LRHyVVbmYAYoBZ4Wvc6AxwOgVg8/gL16owb1UkLgx7
jF+aQ+QMLS5XxoVsq3loDr4CJElHB8sL7MnkbRlCxApv0ClvCHmtSWBI+Vtie2Hw
OtqKxS24bnO4RJrPox/pHteCBT5leByBrEmpuYTW1/o2o8CN74l+7r+U9/GjMYBN
eE1PozhbN4wAy1sZZu1GDydLO7ZFw0q2t1XLBqhxKx30osn2SvE7MzoLmT5AlqOi
RVIhon1Py9GmOu6eKogN5BHKSxyUhgADEBX6kYVXFKYQ17fn8Hi3IIS3BnXd3884
MMQDS0rXj33Vwl8QCddc6wOo0XH9LmlbdGefIEdTTeK2pxoIkUR9JM9dhFdaS3D9
x5UdvoxMAZc2ENYb2TW0cpyzVLmEb4NKjVjRHeam/HDWN8u8YHeCsRCFkzU8rJsv
25KrxGkxF8M37MeX7yS6hZLypJarIT2mM8sAJpTHkTKB+IucAG41aOwqh32jB5jV
Cwa3VLN6fz/Q1YPT0ftztenM60f8VY1vJ5k42VPjR9yoV8m/licUadoV5eFa1Wcf
s9pB0hKMEYvjrNaAsR4N8zv8qwPO17/Y7d5WYDP0Yg3J5yWIushnGRKosVQrlWA+
imUHADVFV01Bhoc8/WALfZ/HiSm1ddJKwYNMHoy/qVSnTgItVBYldegZ2URPm9ju
920QtaDkOAsnmKBnhbQzG3emLFP8u35mj+cW006aRWev7pdXfE/8Hsfbr8PP7rCB
Pt2b8fCl2gTKKESumKDPtoX3nM+2t0IwI6sofjdGEO3vqWBBkmvXrj/AILy1DasM
Y0gHAewofwm/4UcdJh/FyVCoAATXUMwYRTE5Jl2R6FJwK6sY2tBKIio+MdAj4Hix
LVHe1Ve/12t12+N0c6YMLrlXay+4rjpT1tF/37S+TsmpCccCqmDz/8GcakhoFtdP
oB10J03UP5s07reARv91QG/7la3QiVx5+znxSGOYKHTWsJ4En7F7J43+uyRsofbT
3bu2WLrNWIyFjkOzLV5tEljeSP+t21R8AL5eRWawz1ObEqDEkkWVg6KiMRZ5dbn8
dgh/+Z3Pz2hABddrla0s0p7JgMFRpd0PwEatWFoQqykCoM9lAuKKu21HccjOqv3i
YabHdHfRjorIpgc+bcdzShWkkYEluGbZ4XM7IYYMK16vocle9v/eMPaO6MbTP/QQ
3sPJBJeEyW3FETXzLuSMPctPegRd8sRPdU45Bkc7OTgex2LloMrrpgxKdAebr6k/
ck+k/PfiwVcExZp0iRdKwb44JmMGQ/36vHHteWZMj7swETMI7m87FhgiU9l0Sidm
rxrqQQ4rcmTuaP6Q/Xu3E0qhJZVNjLC7ISOrjCQB7xUFcK5McD8pIjtkLQpgM4m1
LXMoyAwo6XSFbKG12aXXv/YrOstAnN1isC78yzxBkPI8xUDImHr/+5FQKlB9oi6j
gBa7JFDbNZQwXAC0h6JllpdGjL/9A4CwiqWNK3irsnXGMxH+0hC+onRiEnlYkcRu
qSPletNRdt5z15NnPEb3MLPwRjtCPRxBJjCGRH8Z7ZlpZ61g3+Opop+lZ+SOBGi9
8GCQh7WinPZzrVapgiQE0aVrpMUdGKDIYV59bw6GjXvNB6/QTOlwoQXIEPQ4ASI2
AEh3dvRy0JeihaGn2HYbUHNw1uCRDTKI+4CDfNOLvzm7Bak24MDpzlxuFfYJcHwx
eoi8niCp/83GQ0fx0/cJFI/r67ppOkU9XoqyuLdh66YHpClIFuaZSbCVIAoCizgr
qahlT0gf1viMGsyuBKo0I8Vfn8UI3xte/FNTpbBmSByvv5KJr0Kq8MeykmG674k2
dTN7sXlDwEe/jMjJNKEUPVQzS9sFD2UHWfbtqXEgqA+0yaTv6YuCBq0VTGdKETSx
PFv+HmEfJ3Z6DC0K+XmARM4gocFe50aD9t/VXMf7L3Vilq+yMEyvWyLq+YaReiAU
AqYDi17HAJFVV+mzUyU1neqSm3+RCtj4e/NLKo21XgxyhNue/xwHYLRqLwvN2UeM
qzw6DXfjQs1YHovSGtR46257lb3DMRt6s04Lo0vlt77E3xOupz6lxV4RIwFZhiVb
P0WbXHAYNUMLdU2DWjDM9fPNySTUtfdYJ2uGYbuQC+YzwPxzFunmwrPOyOgmIMei
rs5XU3Xj3K2hEV/Oba08LuvrDvEj5KdyM+gObNEmadqLxFZ3yICSaIrVzGwO6F4B
5eOfCj4Y3FnplUgEy6LAUIWXfNzLheURM1RtK32evl2q6HG494UHC0ySSXyB5yeP
BOeg8eJwM28C0E/KLZlQyR6s1iirAh5jTY5tdMhT3su75UUAoZtJdPhmxuT09DAL
+ZV1EK6FwGYxowOaXWdE13SqER8T09OCw20qNSAH6XNpZKL4DbJ00+sTnKq0OzZX
+C9MFJATyXPxBEGZikQ0Dj/+0dSLsARLoN8+mZ8ExBi/FG5ZrJZQZhEFwmIm3qyb
zLJK7ole8uGjY1O+yudJNADn4Ny/rc6UEmLyMMUU1AVaDtxBwPNQC/cJ697Ou9de
vnJUtbD1CRj7ZmfR3okhGx90zNrTSMXXv2hNVzgb2WQZO9eHwD6/AQCWmGtMbFtO
bztAJx4c/YEz+AcFJubqTtiow5TUn92lt86tEvBDgm1NkqR0DGKsgVSzL4qMtFi9
KkY6wzkxwKpTqasNAA/ZQRL5CyB4C7M7i2LgjwHxfdLlWLTF6PIaxNJBVHGUOias
NZGO4p7aOwReVp6715fFyoXZzS5on2LkpWIjhNC0M0/ZgsIw58qANFxquRSJXfVK
gN8kWpUwSJT0GIG//JM3Fx1RZ0E5Ekbts0FXLHbmn5I/KNKC1dLE0ptb/NBDsjz4
TTSRF2dTfs/QaGwj7VIL4lDCuf5eti9ckpeP3Ldx/qAMC5xONkdEHexK3sN0KupD
83FLiAXQK3Z+vntxNNvbh5vFh5zIvMh0msZeKz3BuckZXdbb87/Kg8M1/J0NgOTq
nc+P8+Q9eEd0gNQ0P/mf7wCRq9ZvLZ+6smjql3442WJI0ghJNgVWM6P235bO4bu7
sKlDXErCpbpsTjs+WA3o5JjsUjzndECyDvIZ2RofiIjGiFpERD/6z1s0YET870l0
L/8ImcpNhi6kk4T3Yi7IpyQGYLuZ8DU039hp7oHqotJ7yBrcs6vxsKHmALXUPp7I
D3e8iZ1gPPfvYU51BKtLW8WNENHxnBXXNm4KhJOdIRv0ZyEM5rCNCBfSBVm6NL24
ZJ6HybYRyxXStaNgo+Oe8J1BMzOVPlv8gvPrm4xV+WGKrihSutRCEJqVUDU/7Bro
2WjA3lWGIuh+caE6UtCSc0+yCPb/DImRWuceEtY6XRzkaW8ffYiL8x2YpKw5bQME
9RkuGFbQyTGpdXw9qUMeK6eW7ry6/dinRI5gvJB5QMdFCcHK6NKmd0vILmCiAbMt
SrDHrUYFfD5jbkQx6Dgr4/FBEJhZefivoP+jnkchpc23MRl1nYNVUXMVDV+Y6da8
PLibnkPXxHdLnJK7YhyVGlSh+hMvLX/vw6azdnWb+KsiY9rF+OSZIuoAlXVmdech
ab36KOBDG/EcyY/i1bWJ8Q/wQaqV24RG9fvyvRrc66RwhkIog9HRg7On9GTukMSM
2nfqlZ/9/wM7zkggHbzRPJqEXWyfwo2sYGbG7xZ1gpPGRjxgJFN2o6ZzOIDhBNK6
88yIZ9CbFinH68Y1hSKUjWQeErXwczO0c8ISZJ2yBJ0irll1Cu3fSVKCHCtage4q
QFG3Dx9bXbIEEWTt/xiU6q6MenQE5VoTMh5rpSMGqKISW6fSTiUJ9SnTsFALSKkk
ntzwy+uiQrM5gsxhf70SdIi3KCUjdNT2VD8C6+foe5K/NvZeQFVKFGfKTslxLXLF
Dxho4oQVyd//IdabkInXDr88aNtkyyOMRgQAQFZQgNJhKCmSW4y9nh0S16qOTGmB
RtNqEKuPUZaLxna6jGnSZXUofcVg6aOB7QoBFNZHfxTKBkkd06ykWYIGARY05Szi
yUQrkucxhPTZqk/tmjLZnPJ2MhPDKmJBYLLKJl4MV/E1FB2FDadz3CyJpHyantgc
dK9EhC79om7IPRomTrf1TFmPyBOGoxbI79OqIQ4Z72HwT6HhrHU1Yt3Id0pACXM6
YwlNwv+1Q7TjjEHMdOJLgLYOyoGfgtTjI44TVqyUjXpcUtBAbFBKQhpqdhXtndEI
6mN7lY+qCoeqikam1PPol+/iZhbXdO5atmudLtKJpVIQLCSoSOANo9K79IBX4weL
DilHQOB7HM2tTP+C+SecA0dozo/A/7nBj+oP/1/a5u5RG39HLwq+9/ltfuVYYrBW
nfKyOYtThYtscMUF8f88SWKPxNhcLMSgX4k53vJ3xKUG5REoBtR6GY7nfPWOUDqJ
azNG+s9mtpNcqW5VMwVjVrixawLFiB2RQRiEB+dboEXeENbVbd7/tivDjFvBMErq
AAARc/gTZCftk1KcRmmpXTuPvxQCxhBSPSFYvDOrt7egOT3pKXOdUxIxCI9Ryc8k
W8P2Un5yxmYVKqXJozbGyyUPMpAaY8QylUfvo/DRjhPymIYTzSZR/3SPQ2U2J2hq
kt0/p8xDnU4llGTZlNjxyM6KZqzqx9N9O7lnAslkS/BgpFGerB8t1HLIxUsoMvf+
jra7o3Ia6yNMblMQpwdag7yJn3rWbXO2D5+ZTqTnKIHN3KGiEbLYpp7hdzOabrFC
cO4ET652RXBjomS2G8Xf/2A7nz+KLCAImroHFbSqCvSiVSMx9ks826EbCvwTkgBY
Bx8cGyY5aZUI2KNjNE7CtXUUuTHr9eTva+rN1nHKc0K85TyEL8oqr7Tlgiw4Br7p
Lw+7ctBdH1hOju4r9me7/RJG2q//YPUqjktry+bBhrMaazI8rrgNWkwfkzwy6Y68
0jJyJ/JrKtyMqLClnNw3txE3v+LumYLD5sYx/MvufSgjov/4iSdOX1IukrR8RII8
PKZWNOuA00J2S7tdsqEvSWQJrQrm1BjL7StngPEm/gasQqfZkLeGGAhxoKZxAGIe
OqEPNN5s+tzyWJlfPj+AHlds9v/QlHnTDko6i608LPbgdvqSJKenECpWBip9s77a
YF1Qv/6NJfrPf3+Ixy7yKDjd4iqUGuIx4YuuODs4BUj/T204m/CFmb3dh3xsukst
0+ycQzTOGNQ/TU6dqtr7vYGaoqTfOPQz7w8airI96OedMVCWdhDoP8zrqRlxwTAK
Hy+n6N4KiSyXj2S66K3U+ytKBppIanI55uBBCZSHHwjvO+h1zYNaleXUNj5UUbeR
Kn+0+1IrYVaIYDHGApkokUvFYcbQI8HyIkahK92n9Zz6jEiFuqO+AX4manChYSx/
/H4KkPtwUmDecGSoDiTUk9Ii0A3lLO9PvEVWeLRaId8vLUnYqbLmYu8cndFr//6W
/1+K1YURv0vNL6Loya163iAp160Kx0iqrkTxsb4LlPvnAmripg6TJ3FZrV/thFqi
eXQ+HpSUKAjfIAkMDFeH2aY8k/7ZHCQOTAqMImr8TMLxutcB6j13TR9OO64cFoQU
/ajcXZ9jI14GenJ4rLiifAOUCtwpUwlbUWOZuOuwqrpioIMg2AnOB41bVksnj/4f
8L+F94D71M5eFGH4gQx+ZHzF2+xu5Vie54uw0gXXH5GCwbce42oPjW+lekOvblNy
5COK+2EK9l8i5DYMo35a9Qim+TN382U9+tQaB/HdNgepe1wdwbiM1fZluOfRp231
ClneF2hgKKLuwA4WIZbiFT264L1goqUdEwvRQf7yb23PeIffRNaCBExykRmx7i6t
mzKzZCC3w8Wz5jL0XQtVR8c4/qnzZKY4OdT7UwioHPGArKBOX3/dneRnlylcAByE
bdg/NgoDz8HP026vKDPjyE+zFWUHBaFsYNG1RgZOJisnFVjOftA520ZtnUK5u+6w
D78wltlepDotvtib6MHjRvYTet1vhm4PyGn/i4hsga8+kX/mGkcF7W0ADwhkiHHt
YF2+/asAwfyNW+52uikhPeOPTpeuIA/sCjAszHRK8Na7sy5UhOKCReOadLMiafqb
MG7Bhuj1xL6TQbg6uqVoM2NB3JbxCXe7lQn0/auDSeHk5+RYfaWLEjsOAjikX0ik
jP4UY6creCvdF4tuNv45Nh8XBI6l6xxNNSSVvs79P5aQ1H/SmWx1IJ6b1F97xPHd
vqSh9V4nvC9mIJVL5qUdrmGDsoJWX5zryKlB4JX/BfoOy/5A2kj64c2i9RNNLIki
xrFKQIY1ProPyBG3ZeYQa0KhcFBEggV0jpdz/sbCp/4Gz+/c7q2uhvcz60oA1aEx
v8m4pxFNvbOf+U8+FI7YLK39YapY9HjiC1d3L1sNZTySTqL2t6stn58hRX4JGQ7E
hl5wMb523UqMI1LdIJTWOXPgtUKu6zEigxNRw3W7iFXQMtgwK724d7f291BcjRLH
qBUPFLlAwMPaYuqM/FqSIIf/PVzhw/2XqktVVy2XvQuQAlIenkun9x/dhNMp7bXF
mUGrwonudZ9shL8vg26jfNa/gaVaqszHDtA0vWwi8O0MPa94v455NZ1iCfp85RHe
Zg/6TvA35Yxe7dRTdCkQryuWqObC11lQCLUUWhntmIrAR4jqwL41PTUpliQPNM9p
GA8uPHn98E2NTaer7QgkGiwTqRChDKyWnhlnVGZJfQtsw3kkub/7bj3MOrqbexO0
hqI5XFTDx3Pu9veE4EJSyFf/9CcpKUmYTDuzJXrkeTS6XTsvJeC+YqDVwyRYUMRA
QCGJbXVpS/wE9YeB9Yu3tjGyjqbqYk/2Nbsup6pqEF8V9K8uvZjgnD8jlH8Reox/
KYqT73tocxMoRiVhDTG8HdRMB4WJgU5YvlLX9ErNduprkJeaFS4Y1Fr2lPALyfDx
gf77YXSNcy63vXHN30PYfp4qQZlMvvm0IkjcD2RRvCFWR4JSUswnwGbUAb6yj1IX
fLWcUXtr6u+8kIkAGlEM2DxOJrPGmvNYYDKO/SCOdnWBErHfblTOzyNwHPjTJTkh
xGZsVNAdUZCpD4GXwv4SqRLqcJ+Oo1W/PY2KsnxymHYBAJrtWvFsinq+bWDsQmNv
ry9+/3fZ46jpZLSCZQdd5aYzB/b8vxTX+6wj1V9XGIyq6YzTxx6o5pBxnNEJ5CCi
shidtqGQ2txgO5VaATuFFBECBC9yYf5QBGH52rIry3mjFNF3qk4t8fEgoyKRmvkJ
7OsUQu8A3jZPtaLLtxTlxxFghZLizdDrrMWyTW3ixOrGCz/cIb88tSluUwlak+fD
YA+PflVkt1vW+yNHXerULCx7BRxIZrbc7S4jKq6QCF1HY1BKHGSqoC9C7izkewLw
ZoWSfrdNuU9h2ocr2C47ddkle3juO9WUtIopB/bWdE1DF3ptdzvlOj4/Hcs0Mux2
G+mVyJSebvnvXTwbDUmUdMH+lusnhgQCZJZwHKGwp+EjVDi2Xe9PUR/hJavEQqlh
PSQPxW5mDHl8sQg2SLbW2soKHNk09cjUcB/zHeT3xx8tBiX/jgzZc3z1U0CM8+F3
KIUnBfblFXaNAO+8sf6TWzl7+753LWFojKi7EFB3WIZIj2Qcc7oWjKkFFRk31fOh
dClausIH0JUznQjvLFmFoVMzyNsmu6DCEh1bi+hYPFAwhUD3bGX68idcL/nfQWmv
TzIqvZavVYSTsM2PjP6GS7327PC/o0IhquF7G82KwQS9/4EXme44mqe83RhpEgSK
6KRADqjhoI2XNYV56NBslaTmNxg9Kl7J2U+xmN+xgUAXs/7nHsUUMYwdosWEowkW
iv9Ef9p2p1M0fUKFESamiP9qOcw6jAlcc52KTgKzXPW/P9xaU6t/57kcO20mldkF
`protect end_protected