`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16560 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRpcw2zQDHRgJxPf7yaQH79KEtnTCle2MtJU8K/kQpZKH
fI8TvDYlaRaoZ14z44xXz6ci2rrSUqmvS/467lGm4zRRVvlA7F7l9itNQXGa+vO6
mnO/oSbTbTCAXI3avEwDaVujOhOY/CC2MYEG4axSht7g0qfL6Xr8KZvik21YzDAG
pqh3g2yidzfwN0PXAcBv05ROYHlNqP1iH8ju5RR0tc9BOJsESgvGS9H5H7tU9aLZ
KHf2t3OSH6hGhZDwtnFEh2v2zlQwlajfbUGIyfOlQJe6s3AuZPEBNF1WFFLloRKe
+Eb29jPuC3SiEgaPaW2mEiPjv6LmN5DtyF9x8s9263eMC0US2bHRwtFEX2GWiVEx
SQpxMeIaRVYXPQIf67ay1vOez2QrpVg88/0xOYQ8pRyvDFDONE71aPgt0mSjk9lB
2mQzmUXGZ96kRRlnuxrsPOtO9IMX0OVupUWWavHSUlXVMvflyLXWx6GVJl2sqgg0
dNqaUccimsLnazlYwgIYXbDBw+gwLMZ6+AAfPL2hKmiFrl9OkKMH+4V1CaqI4Ydh
0sTB6G9rm0cIxmJN2fL6NRypX2mAXZCLoHoUKNHPfQpbabVsmGc7pEquPUTV2+kb
VhPAfiLuAKmMLzTHDcoy35d71duj+8IYQmZx9wzcCmXhOtrsRlsIhZiisgyP08wS
zjbnXhPFqmVuu+/HM69357FFucUOXFcUsHGh79vJYwMqGvdOCVMRR4T9tfbgj/OG
xwudlkMJBkJ1FvsUTfoMHBp46ZR//WGyBUTh92qZdAomIY1CZ0/r9HUO5AJg0Wiv
kIo9qeHMGWvYVYol8kAY+FRZi0rb6lqLsbIHhDTlYpg42XnklvRvNZOi74ePgCKJ
GP0XKCXW7COhBryLHfpEzxPlhHcv/wyy5cKyz3LLEPDQz/+TMFjSsjHd0U4q6UOr
DoU91AXJ9Hq0YLGjDX9/GTnlWFeJYSXOgLhLSrElE+7tftkwT77pqoBmWJpgHPiL
mbr8lv08boXnNuF83uoJPfTamoUmZzM4RgcNwBkNSVtkXwqJGzf0xTt4gk0PaGyO
lbIaVV0B4/h1qsH9e3rvbbrjdhapDhnw3LaWqzugFTcLk5kzc1z4NVaRTWD9e64j
8MA1wJtdPET4UzTxGGultmYa3/qRj6GI5FhY44ZHFzi0I0FA32j0E7Wp1F5gB/RW
cV4j5tiYfj8FNq4mjrOzoVmRkP3BErZp6MoqzJ64Xd9pvGd0qgDP48N/xbJXSOuY
4oyrB06WtNnv/P9lbOWxJkq4G8wkDwXmvITlbvwSLFi2QX1lrTftkOjoShjBDI8k
HdPV3oDhsE2BBGQhvFL2HjCgRuuZ9NozGhjNhJnw2vhE9R5tdet8jz2O38R2ILEm
gSFwlbQliCrym6I1RRjV59OglB4Cj/OyCE7Sux/18hl9Rw2eohCvb9ZsaWpfs8py
lgn8KzySwwakvIMhVZovwzdIAovexiMOPJHDrfy/LYF0SFpa1fem+mK9gRX5qssu
AX2tHx/JgdtICHaKK7ndBiLp+FjiUuYahW4Yd6+BK5BNj58WdQROK/IRaWGyha9a
oSzcoULgdptsAOTtdzfNvGNpIjyyaRirNFhrpK4y5CG4x6AFLQvB7/RPWAuCKONW
WRCtV5CAZ9rukPmlzC+T2b5CiJ044jz0CEzSyo66n9FqML7t3t7OeTjwLoiu9Qbk
D/QobQWSYqK9OeEc65g9LHipzSIdnPVy7TAGykMqfFuFQ0F8wo8o/LvQShrqZm2f
H4jpYEuod0wJWSGK2etxf+flr6LLAoSLeBGu3cqzMU+wuYF3Z/f9bdTBmcnobvQa
6uXXrakCn4rxGc+sMqx8xr+MGBaaOlvciBVQNhvIxtceNNEctHuXtMuDtvpIxJ1M
K8KyakURu4wC/JmUFjNpY2E4KBLxomsF7q2/tstIu066DKdJpoF84yqTWX92wQ3p
S8NkZDNJhk2DGUSNL1/JgFQGGT+iz18FeFMfPLqUUaACOSbzNqB0Y3miaqtMdJiV
gPj1VGKt0iMapsI6KGvpaO73QdYUaqPpBalw5ZWdaohjHEQgOt1QyN3rENpY+y8v
Qj3CiOEHNAAUrhLWcQgIzGxDYs60b95BkcwPdYzSDUR4lzF398FLC20zs2tIJH7l
io70WlHjXUmeZb3L5tWwBpLCZT+i+VStlG3xDR8ZLB1ynJrbv2WXXwYii4NmfYth
btQbpVg9okjco63VSjcLsWGZQu9StBcXP0uiKNShu6pmxJxZFojd5ioOkFwo17qt
J9pppvcZ5CGNoLs3/ZCzA/0BXzUBsdmsZNAB8ovqwjRwYcqm/JhqUHbbxnF9D3hn
L7MBer/FiuwMuXVdNl8SFZYIKV2YCBMOguitpyZMU15RAdYpDmpFKcUWwGmOvBJl
C8y39EMVRhuNu4meeqI3y+nLxOccFSWuZPIcdukrVllhXb0HAXJ3ekAp5kAGSuJe
xn7YOZKOdevWo8ZXsOduwAh4nvT6DxUEvV0wRunjPAitfrfY+Rlp+IT/mRHIEm/6
2sFIOph6Rd2gK9QrvOZt7g8h0f7pQJkpDnDuvcHxTnfHysrIs1Gqd9k/zz1iOZGY
PHPQOEwicNu1Nm6y8wFk3mLni0HHHTBuHQiR+xTa6gmrt32fl26wZ69tqRhj8bbL
Av2d8wvz+JJRiiaJKpyQv4e1GEXi9HM+6QH1p03cMe+N+7fL4oRWr8juQXP1cRcU
a0A/I4+Jqbg7G+N17l6JqZE/y+ntGhlHXnicJyvY9J4W1dMsWl0G4M4eNlTS35b0
b3kFyXk1kZrMAiS3/i7GaU0+L8hKwlvt6ioZ0n/jGWBEeh1PFxYfsUkt5fTaXN3I
zUL8jjYljDkjMucLNfTlCGDx0S8Na2QPhYQE1YvG2anUqUkQdDNkhW3KyftboJkZ
6MmL9AoWqLgnOtqZAyRQon9cBf5uNlWOeu2ZeQ+HaPOVkV06l6eR/tAOsnH1O1Gq
EQ+iiFFbFBjCiwueIBlRO33JJw//u/8ZaES1FjXWkSWkDYKxURdMxzNLrl6Phv9B
fY4V+BSRwl1ptV2ak/sXNhaRHMxRRPt3x+v3roRJuIqlItVoBUJ/jbItkJAsDugx
hnOP1J7VGafjna1fXngTD0gVHMNA9kGf8ysLPngPobCJnGVQEVc21ATX3/AepqrC
R/fhQ73OGwSr+95d+S/bsazwPP2HCbjoN54YlByJS8+IPLZsYCOoETLSMoJt0yQy
s3M4MXBUsmps8zbcAC9Q8GK1rgUFOE9Tsdz9XVOirVMh6VyqCzsGKLPygCoBah7k
i9kYd2hM6ut4ldxEnwl0Seb8r2esLs8ocmLeVADQBuLJKX2GgvrmWGJzkCLYNHjb
o9yU9rDkrSs5VNAVQLE5C5he8Be3fuPlNPpqFB9lYwr1rTrtDU8wSdCBCaMumedW
tP5MBTY7NhsKs677NzQGGE7qXAZfV89NLAnVQX4LUPEyF+DtN7W8OZ15urprARVl
aJYYZeCGt/gjuQJ1H+9jLn7q1bSOLPWKYZbHFjCTZYsRvEd0VfXQ3vYZIEUAu253
q50gmEadNnh+IG8uHPuUj5+ka0XG3gMO6S+U6EakF6FgHw3XVojK5Vz6cm0pLTpS
orRxTkHbHZ2zBIC+2UmbVsgMhmo1i1tgEXlwMXBrdFde9UOLsvo92CdTOj8Gvs4E
le/bI+x1NRsNdlZoFsZzrYpIixtu+FHPXd0t14+zbEB24yAsx3/SukbrO1fWujD+
yOGPt1igjBMkxlH6U+kF6WMqp+qeYtQ1u/00Wdy0g3mVNR0Y9T3Irj13NuaIRstF
HmZ3xRvtXmcPz5HWc80GOE64xftHJ2aJ3Forx26rn98ehtowFrGwKtS33nSYioSz
oXj0RI59DD6rwa9iOVHnn1tTntbu0iN8agsakGS++0xr6GansS+V8BN7qInxXDac
TDdQRUqKPqpbjKdUHXd9T33LjTq12iis5Mp6r6Wu9r6tNBORpMCU4Bk02SrniZga
Ygd8YrbCyZSHMYOzYJUtlKk5FT0WqmsYazhmFImrrn/Co/9bZaRa0THKtnTUlRnK
wNDTGhLcPeSSlwln23eHBayYut+bPEwCuki2pbF9EeEFOdZCtHzmPaztEm2k4p8h
xw9/+IKJBZjEM2fbEEdDMK5jsIoTwNokdKj7b+RJPn8ZRfkksc3UHD9jkzWSGk7j
4dwjXYUBB4Q7kyn/COwuBske9gTdyiTj8Iq8mahuo8xtCw3BW4J3qGlldBH7ONIC
2v9j80wLewayygeCk+CdIJDPbRspKBrsczMSpH6r8fmIO9MgX0XvL6iYzaGkIg2R
H7e7G5xJ++W9o3bMnV/vrYmBL4flxLCd+llf6EhRXADfs8F9kkgLqebA4sAIDtUb
NnRaZj6RQs52ye9VRGVayX4Tk80swrWuoh8GI1YlTrxf8vm7a3gFHjJ5ZxjRUBnc
TkvCWSSA+ZTHeaCNMpvnmhP+TcDQtyOWodIUe8hAk6wRBdXd2totTXpQzz+fSzH9
g0CTZ/Lg5mkyhfhkrfM3CYId+mTdjuMRtCFRgWqsgERvboWo+7H/N6o//tiCQhGS
uFy93IPlEJLPHUBYRsMr5WUFaUZrzSUXN3PSDHFvleoPVwo1L8kCPtDrV8LoRIg5
FX5t3kNeCuwkW27GPS1304P5m6buwzitVqcPLekOhHlwojU1/IFeNofErtya3gD0
x0o/+J8n3ia9h07BZM4UBPWWZ7m6nN+ydeNXQXiK6zXLelSYg+e+Bs6bP+/Mw2FK
i1FG0AmHp5XTDI5uOVVGIH1UKVjAWq+jylxBgTez/0UTnAq4KNAjzYXVkvo6VXDK
qp5lPI3WH7UUudkNs1RrJIyVCfOvN5Z/qoRcP50/FhpoXlx/E1cQIFLY3Jhs4V+p
lGOuo0tlFOetnB4YwVlLobwD1W39abHqm2PVuV1+ZcJh/YWIQoDa97PeXzgnBEWj
59maR0UI9ThYvG1njI1Wd/sib+scvG9IEu6v9AxvP+uIXkxYgAe/u2Em1tOPxlK4
lrScp+bwnl2teVDjhbkGXrdL2UR20gCIQp6sBeP0VjTTrgUUBLGVLTBVk86ddSTA
JfZWrTT4Yr81XIZejE9repGKwrRlQobqJHqjE5XNmIz29xTaozegfjjnYkpK7LKf
UvHB4/H/4qMFnaFtg8MItlFQCrgr5PZzayJjXzV6NzGPJzEvHen7m3XiUJL/An8j
mZGgwKplNmWnpBvRfjOxsttuxGS+VlwfZ9jX1ZU0qJbgYmHPBTbCavlBL9WHJnf0
sBtPD/eqMrO8lhX4D8Di5QnvGf991CpShlBtagHWPF5wvaNXbsE1tVZ5t9yH1V69
k8SRh2gFQpM5bDxyuN9U/fLB3CQ1FBRKAK8+9hbGOYIfcMbJ5xoUY2ottj/L/UIc
1OHoMAlvRmnl+Lv028gzbvevxXwygijG5HGu3eHk06d8S2olKe0K7VFhUwOpLvcE
89zW70aGUeWsSJpPr7b3QvU6GZ2tUu18hjjzJ/zL4NRDyqDtYCOW7wx6oWKLGqJE
uERNqjUSxDzjlxhNP4yQX/0aVsQ1+yTjg9NPV0hAk/k8RS3nNfRWi0Jui/iLbW9W
AjMQBn+CFOu2RfoNbe0NTOt11l6OkwYs+Q+5/oWDwlT1i8G37jTuPjNKRDK3mIAH
fNWAPAGotHVc6KTj7w+ePkYxmnfXf2ERekzwd4pVJd1NWZ+f9shC/DlVlg0P49lW
AtdQcfbSKjhrDfnV/dtmiyj8qKBvKnt68r6zJpJAY9UfaJv425kcA8QzXkIYkaPu
8s/EvRNIvUTchOeXJfdX0/znpON0PM/fhEYVr3Kjfn+JBdx/i8K+6YOp4W3Jce94
mdX3FzTS2zZqe90II3yJVEhb2SyMaSou2Af6dzLtZkzKUGbWs/gNCHlmfXa6RSha
Mcf4I3t7aaXmaT1jgy5Ow0ZpkyjlotMbU7DkbzdUMhOZjNc+6XUNP43LUQbIewRS
svb6xblihOgOHiEXdZU9u1G14G0ikcHO9gQUuXddFuqrWHuUL/bb+L5JYK0Sr1W9
rIz5RGbG35fzsLExn9EHp7mDP6PBpNMe03VjD3EBT1ql2Q4ri69DNyskoQdS0kDB
7Tm8ic0/U8hY/qrLEQKUtyI05+RSHyJqCDvVeaDEkjyAkITQQc6qF90fyDRH7QIe
jglKhGgt3FflWL8reXfBXtWaSWi2nE6bkyuwutDIgGgj7Hix1OuZ4353sneKTRgp
mA4WhJu7aIfVro2FD6YXnvY1S5yVtKVqigyB85z4mo7qDP2klW+/b3cvSQX7Ob7D
f6gd42BXhKfcEu08A+2j6t9ehm8w9rcxNFPrfsga0rvawhB8+HamS/EOKuKxeL3P
6lRjWQc3ZZTBIFsiN4rf+BBII73qiDAy9hpuJA++cxkIDUuUovlxOvKO+NvUMSRW
ZHd7K2GJRmMV2r4fN1wj7B0VUp77gKHU4h3bwXl0lui/IDwu1GDinkGO3amP1qh8
NnNBCBeDhZ3Pfbjv/KNcwtksIziRq0BCZ/QUpm7z1ERHjVAGk/e7PgN/q0Nk2j8F
G1jsbm332jY94jkJG3FIY1mUW8huQIjDInNMKQWGJK6pBDfTlW7rjBSS+7tNxLXZ
2FfWN22erIoKxBvZpkQE03/VY4z7GNfoDoyx7vCWNiHs58WIVTYBB5A1QZ/OGWQS
BqLV2cDng675VP1n0PIXuFoa5IODv9qiyGifmzV78aDXoSQd1RYDvSpMlISmVYwq
SI8odsgFSQkcdjsK9USpz6UsWOGe0X06BLz3tqmMcDr0uI21jBfYHz7cmQtXwAxg
+ZDPO093/Wt/T+El6XEXGW7EpKDIuCg0ZwsCG1i8JrEMioEeqfwOlo+iMkyARlfn
WciEvS1AnjfcIGN7Ve/pE79dlhesDcmIjy74Oy0pV3XnzI6T/NKa6ehSUgFDr4lP
noVRAptkvU1MQSrN5P7J0QPfC0UiCq8k8+qEg15g3LH+1yM6ud+JMC5w6AAhmec1
hYny9PUnrGAr+QMxPAONkBKuTJCVYpdjdlOjao/k49ZcTya/JSclqn7i1b8IFOcA
dMCLqeb8BftNx4j1UKoJJ2l9X76K4VfeGwD8xmCgiYDP2k3EhEuPf/Gvv9Cj+kn5
cj5vSVij6kgWTQlHqvFjaeXSrKt1WhyO+W4rNn0QeclGbKd5nRsE6uwHrLzFgyQR
6tjPszBPpM1JbqBEMVTDeZBqXVYR7t2X4RLT2YfGwjBPIXVfQJt4xH1A19V44cKs
kmEK0R70lCFV8g6FSd6AuJ7vueENnmFJ+HxeVpNkHzYgvMPzl33lJcJI8HGXFY2X
Z23JakLo7/GV/mofjqeniIAAk4dyzE5X6qTkuh9rOA7pPecyL/PjyFZantJL2Q0O
bqPr6pDZFSRFp2JzYp30W5dd5IFdWSJeBeIS1fQ9WIsOi914WqKnmc2t29HjhMj0
UtPdtfznxWANfBpbYoxeBJ9K1nHNL5QeWF3luiIKfp8Wpk0Cczaw1ktP0efRNgDG
titRUMmtr0fIJsnJWV52jKPhDKRNJdr/tr4qK8S8/hAkRzpHy9uC8cxF3IZttc7F
orKHxPIjAjry8fQN83ML5S7xxN3qcNCk1dsGKHNyehG+GyQeC4Oxluu6MEIbtkzk
guvZAo59tKKbvAbZjf8tNLdROLwR5gbcJPk7S3TW35hPcJAaF7wSO0I64q5w7nEx
Jz5eaDsAuPd3QFkEJ7dKEVeeD1ubs6GsFo2vTJHLHbVrEQQ/Nn6p5Wuz45XpwBOI
Pef+QplGf/NKu3mQyQhF/ejzHpiUtmEVmqfAHUdMXZGVpnsHuEPPvGIZyDXh3q5i
K9AkDFCc3b6SsQy9nvGPNs3AdvfTWYttc2Sz/M2AZYJTJ+zsWtFrYq4gMPvL3DDU
p/zdgOpv3rsEsBUeQchlA/R9s+yLflakcK8gFmfIS23srCAcbvauzg+tv9ziFIY0
8b7GN9o/afNImm92/xyAAjbMfIs7O+SW9JJ/EzrezW6FnI8F+1nHaJkWcFqZk7Uh
yVsak3RvxKh+jd3TFhPzLimP51Z8Kfvzn/gJa8RMfBVmAd/BVpXndfKoD4cLok8A
Irk7X7EKcWrHEfqnLF30+dfyk3WgoyTRkd0wMOn1Iskeoi6Nt+eRKC3BenNrBA4I
iaYUJ4DxNHR8NfBM8ChmlOcO3vCe9AAZ47Uj+LJdoRPkRvZquooSjIaLChZLkaBU
wSd+/Mh5hwstZFXjqOd9tggZ2njogfPDg78l3fysgHb2Wh/qt0ESD+To0gOpFnBC
ZMEru3Xxn9eNkCZkYpkSdw82K0K0hbu5O8aWn4tFxG6W0aWDM/jWUdp74mG6btmD
zl+N0KVvwCVoPfDYL9alL83e7v5TVDB30d2U3V3XTvtH9eQ5TS4nveheUhB8RKnc
TiAo08tW9VoVUGdJvw4pKOTiCPDM9KQByvf0kzAj3P7hFgy4GAjH38bFJZoZejv8
P6TlLzPxNhzXDeqQKkpEjcm0CJ458Vc1qRCAA2C9/2L7FshqZI+DZMFAsDXUUuQr
2qtiGbthvpVaDYhFof+IyCaHpHxDJhZwxCcpk3MIP86WHEVu7ZVVAQSk26vGS72w
C0DpaVuW5RDBqoJL7aia/0GlscztnAbAHqB5DD+WtNjOY9c+sLOCKmTtJt8c/B9o
ZFQizVrDIhIvxTjKDTp/JZiopJNsgoXRjsGg+NlMZX2Sq5fXnWXOoZA+PJLc7hWz
ZmiSk5hUZWz0IebjiIfODoX7Chv13bBE4hwazIayh45IHBlHSJ6OGe+oTDd4meE1
ta3cTV6AGvZNwjRUEpZQRidEcexeqWzb0ZPyZCEhbWCFrU2lb9i+C3azMsZ1Nk3m
xwxhIL+kHUXB5iGZiUQeuPPNdsarJtI0lHSwyUrJ3WTY3P4nufXrkO1bVbufgL9g
BIQ7RgMfIZoZSRs6sqKJeJXRS64D37ioPdnYSfCyi3gZoK93PAiRrIOr47ko2YjH
3oqLKiRM3v+tizMri3fcFQp9i8jEBGecOxAyQ05F6ol652uW88AvnvhoaPzxAz6d
1OGwX/iyCqOhSaXwgbtkymYLc/PMVedJiYL8FBCSKve1Kz4za0AOTaYxfEjyMUJ5
WjAqqi0RafslHs/1/TSZC0wAWHlz8IiTusVjMA5dFTodL0qDS4D1hAyp9XAYUmbE
cvr3G6ogwyfb42NyHQHtqenuA/YJ2R7dRculNInB49DRmGjNuoP8ooqLVfGhU0e2
smTap17nUaBpiuhDehRFvKex1svmXmUsnZfoEmxz7xbzPsy7T4/+THLQ39AwIWIs
iQHat1MXZM9y+gLU+tzCn5Diw8jLa70ZZtgb+++2i9cY0e5A9mRlQ1jsEIdJhgd6
lDbJvkx6XY6G57Msc30eyIaqY3J/qF5BZBgH6uFHzLpvFaltf/XpSASSJFMv7yYz
02wr1K9bPnterDXqgVquZpWiyZdysoLSqpJrdEe8oNv4XJJNIOJkQhwNVBahk/Pa
KE8nNlcWmU+BQij1SakrFTQUrjS2eV0CPWEMirtHl+Il5D/mrNHXyI+vzCSa+0zf
I0BOYD/4AABEiYGpAvRaSHU3fKVn3T39M5EDVyVUWqInuChoCkRrhsMRs9SIczah
exBxCF0CaHYr8e3i+C6FejueNJXz1aE+p91ovRLY02oHONY04okp7Ke0mqGyjktb
PgYHYsUWjHNGLiWHT5vf5B+mtVCKfhxOacWTQvml6F8kkj2yP7JAZYQycGUTPH6w
BILs7CE8X+4jHzfMuZMzFq7avTu9UKQJzKaDiFx2uNjC7wnZ5/goX4Rj29n/kT7K
rcBiG7kWX3wdVuxgWvFt6FCcLItBA2Zb8so9Oabm5D5fY59SJpm2oLorY4h4ckeb
uY0pDJuQhJy1btLANzRElllLQsDsSkVDu11n+PJoWu0crxd8ElBcx6W7a3fo8NHO
/LHgahGmMqjWNZGpe5jYuV0OhIDUsPfdkmXkEgx0LJjWi5EbALeHexniwHJa+szR
lCi44PUEoRRppa+BHKokOCpHpoiIdv7EPF9JI+FFg9OYooSGPPPSn9IGqkS9Bufc
uM/nbhjtQDgtl5fid+IjXhVd5M/go60yuk4cKLhmlZA381073YbJ60xHbXhZ+qJd
v4hHIjoypQ+mhMmZSc2w38kPqwdc9BaZeqH/B0CRlOi/cdvHI4i9PYrzN/J1wpHl
LeielR5ew3iHDmzv0mlrbs/3DTr8lsl4KCIEBEuErR0BTqMxOyffAjnVFzKnkuWe
ZPBHRr3b50SMyZWpZjwRmW3u++gcqpFn6k+IbC4YJEKjp1iEVWfl8TqUkk6tAfLr
6zAd2N98R4a8qSwVEcpFzQZgXESSP10J02DKAyS5wCMsUfJ7cF/Q+u4LxDMSKZK4
TFCaZ9LcXISZsRDcmLo3U+58KPHhXkwzvrX4P3UKfAmc2wh8jHj7yeXPec2DZfXv
ejBjfoJASqlte5xB8HXUYlwoc3Xjpdk0LrKGy6LNBFAc+AnDjtWXnn16V+cVe/10
cDitw8MEBlx40vtuPLcvZEFYkUB7N2/xvakvOea7lWEBllpW19w79k9VTMF9qAVA
RefzUdcnKjLRGY71zn7Ilu3hgmMFOPlHHGCnncgwIr5CwsSHaxpbXbEw3RFNyN5I
AGAHGaS0wl7p3juOUV+eZE6UkpkDxFnPirwei/XdLXAjTgtWvpJSMD7v6HY95Nh9
mH4/eD1SJbHDeDHScvAWPRSrTFSmV1456i+T/d8odI0/MFGZP74s4rqdO77DCWNz
0ys6WlylrowKcHfn0mcV+ehhBogpSQf1K98tPw9yA97UteOG78bdVBwGwwnh9ALa
3Fsuk9wUpP0FGkOUyReNGG4tX16m65TJ/huGkjFNklgnWwNqp/caKiy99OPKX4k3
/krY5FbD47OPUhSyDQxiDj2+t6FmlsmCgenAJY960texgf0Y48oXp27ETUzY9RAV
LAARGwHrFhet6TSZu3GCRYIPBxuqsWakFK86ophGH25lkO5g+wc9f7P32anPEtfk
bVPRUqZ794d4WGzN554Ow67G3pcTg3LjzwXhSJoAvhNETuObtJSpq1w4cxvAxKiA
WI10ee5zx+wSv9h7H26/E7Xnab96yJE3vvnYZIAGd8r1kZ3o8CervGoCZKYg5TJD
DGIv4AHuxrVNMKx9aSqQyjfKs/LMuyj3RyVyflvPTOb2kNy5kHKHX+KqxIqOAwkK
Qc7vqMMIa8btN67BHUcZVaMeVQX7Jq1d4Y+SE6DZHF3xOI4czJlBNdvuKDtbznXp
Nlhh3IPRnoGRr+r7KBS5B4V6Zy2B7l8Y+La5ncVUEkJwrPLprGJJmw4BfY+xRB5v
YNDd+Z4RY0NSV/G4O3K9IQK1TD7MwBdaZzamP7vKk5gjsHW/jZEvq7fsRFwFV8lN
4GxepxKqay8OLSY9YRGmB+vZVbxE5obyb7aAd+2saO4QutNJB2ciCJRMuYymgFEY
GGP+yByh8Z3uBEr+YySGWatbf5HnQi9YRHiYyxuZpZFn36PuwKELFE3gu7mnMF8N
chLAnnJX0hlSdQFI9zRZ9gQoUptzFDyoMONN9KBdq3xQusAaTNCHIjn94uHjTlyT
sUII7wzUuJTc1mFFso+czpP49tRfMdRUWL45yKckqrkIzEMr4wIAprr16kjFxei7
21/dU4yRd5ypnJ+FBLfWIwWpKj8SbyepAb+rJ7FbUUn0WJaHeAwh4iirtA9p7e3N
Igenw1NtQY/Nxi5qmJ5GXbpBeSWjzhUf7Y0QqPlGdhSTOaFCrTEwvv9Efdc2qoZa
ifghypkIYi6NA891MDc7LTOjxsajWWj32hRa1VMcKq+eCzHo8qfpZVfDBmWkwqJj
RhKMNu63iwQt9exYQm6kzWHU/OrvOeVz/gq68eVk/R+yOjl936qvuTjcQh2rNYgN
Pdt5CrScgGn7VuUp666uTDASPZ8Y6PG/An5TiA2H6v4fd4DfVx5jh0nwoe5fHLar
Pcwf0Tc+EVXDiYv80BzrUXFREC9VpFDMM6u1UY4Zaz4SsfiZP7T4kMLR0VR0mxJd
G4KnPfjC42RAkb3uxFWX2HnPApXFUNg5wJIGdD+mf0EhNlDbh+URaygas4phDWFc
DzuTm5uDP7/IxmJTLZ63Tnj9Ts793pzNqeUHixFn9OqgIrBdVJMuX8Q9xAO7cZ+3
0WnIkU53LBQX4f7TTi5/jt24ZZ4eYsHsuUwMs1MstGmpDBFKNiQr3zTP7vRRnnhj
d6HQUhbFq+jES8SHgm7hrRQ/ru/LGLXnjWL5lIC905W8RRh66KXS+MGxXzNLwbGr
zAOw9e/7fKEJqqdQoBUNcQeH6tEmSeAIGuqiJ96aPv/qBvZDcj+cfktoVl6kcLBt
ByYhmTL0XmawLlp1FAxeVelUccTG8BEwbxtcBswfLEjYkQkCJQ/uoLye9Ds3bYEK
ikhg0Be64U0qIX63bViOUpzieotPuD1kgxNDdZjfZnQZpZ48HzMY2GOzsPcBboCz
97Iy1Lff3P0uSVAddrA5QzrvfIFXDvxNhxHU+GFvNtu6Kgnu3L8q38toezl0qwaU
+r69X+W830KCoVNBP0fvnRqONUFGkCK9r1LVzLZW+kpVWiHyXe6FMVTY3C1d/63o
JJTavjcEKgco5IUHs6zeGWXY15/e9Fx67R3K7aETeTkbcWLKLuhBISp+cxyYwP7B
ocZmyqnr7+ixwU42RxK75PKxZZCaN1lL62SC94w13UqnW6ECWTN4EFluDijUTSzK
w260c+GskKcC+SIIo4reZumJ0saxLXImVQqDopU4jpSiE41/It0Ig4Qv1wDJb8lR
gKRlYw0/1v4zikJFWAgRhlST9/rO2bsO6e4QLNSx+WY7QHYVe6zag5C9KwXSBNZB
4OpHJkwARGtMG4wZSsLUkqj2HNFyjRLplhMfPlpW3ybDe8HbA10xv3BTP9P5e1h0
+AtOKPbZrf1Ascs5b8/s1mxW/AnYNy6uCj3NsdgZb0i87hZbMLnxrA86bPk/62kO
R2hpYhumUrvXkkCkFqoJ6p9SgqgUtxH0mKTcDth/JYLF2ixPnKrYpIdF+ulJu/AW
A40baXrgxanpDglXOAMvQ0KuvKoNw5LFTyhftectRHkoGHBSzASLBNzJSeu9mYVl
dgtaqMge694wg3Mbo8PIFLzkEdIBQ571PhxmsNgjp9EDtk5/LXXWoG+UQzGuLPxL
80ydR6djxoi7zmcG5rv6k7zNWQIO+cbojPAewDGpdetKDJWgVxUDQ4VasxcLnVyV
vzIBQj/KiKX5P7n7cdGYHio5PBOcx0D9WcJ3kIyZgmNTjezKxKUW3/t0VnEfNEBJ
JVC9cbHH9CbauDOlO9UAdPzvIq70ITuQhyxFHgwAygxe3FZj04rO+iRpQg7XUkb/
c1MrQacCpVKtLhj4BBm6eujPx1fjaU0UG2ahkbOWyaE2sSBMFb9YRe6d2wPwE1Cl
bbxLH6XrT0m2sEgiT6lePQ72QgFVEFjj3+hxVQw6UJ8o3dVIKAc51eYh2r9h8c1q
JZPg7st8x8zLmbALm8V+OKVx+P+4+fu3n+qDbRYT3qvpDXJ43KPVeOkaY+kI1IuD
73N70mzKbMZ4akX6wlbmclptU2SlDe8ow1C4H/F2DPi5lxI2Lvr/vb0mJonWf0cl
nAiv9jzb0bchC923EwBqJm3AGmm+jgGZhjH6Jo+t1oj9x7jD/EVvxVBQ/K0ho7QB
92dHV8/5BHN/qbp9UU9ETe8CJfQAxiavcUI9JAeuFjtCmkSL/b96ne8KqQJmpyqk
J9H9KsjfCJNrVsMP3PDwfEMxo4YAZQ9RfawryvRe+4IqnBoP5RqBOUPwc5EHLHic
azr+aqlz/6QXCev4ti+uN6s0wtOPBkvt3TZhUxVJojn1kjguc3eDxbtqLBvCG6OU
ePYjf6JJl6JkiSGL8uLmNZ3yYJrZIQ4Cv2+WkgrRXXbvTL+MBI8WmuuXBhP4ab4D
pNzbXC46HTSdHFqymoJihHm3Zx5S2alIVFmguNs2WlX1THdhw/PDlxbxslcpWkvL
h/34yL34AeLQcuiPgN+gGEoaX+BdNII9buxm/UkjyZpr8tzkB+vD9/gCBymIHRKj
O5OA60lXOLVgi0752czLzrWJJ+ZMKKrOw8E4BlvlGSb9gUt33FVtst9e/FCnPKc7
JMrItBdrtlVF4sGy9TyJ798Rh9dB7oRj4dPMT03in9QNC5RTxkkvJkANGH4KF/M3
pTFSem3NEF3F7w0LM2WY6/0xEReaIFzj4L0RguXGbXoAFGhIAueDvlF1T5OC04q3
zgHtSXshArZeN1wromPcohqo90wqKDr3L1wBCCKExTsxnuuj0Vb8IK5sXooKTdaA
5LDEahcaXaMhBwg4InmWEnT7oj5J5rfoXwXEo8ZKmbiiAHeEyykhiEQkq1jFyWcV
9535MPgtCllhm1aRMu+jTfe0Z2YRAtUtA74UrQjNkPBdlHhUv7qKR6FVj60lpb87
U50uN8iih6yTT+ZVQ14i1pkAoluocAHIHFAx+N4ePCJnRGOA+riVJsoiwmGUQs83
1MhR8ZKx3njLx//TdwrbBzLb+AiYtGokz0Lfo+0Y6yyDtQFt4kBlIHbZONqqJ3YP
y0iJS16qXARi6SBdp5TkI2mcputad1Ofo3IfGJ/Fy+PCo+pGqlIr0hFpXM5XO79l
GaypnXHp/c+WSG8/i8MRtv+P1Bz3LEh4e47DR/JBoK935WUgfNzh1kbaqJj/flBd
BpRPkjO9W8frUdgUIpt2uiKPaZLHQGlCEt72q+v8F1emLQd58WhWYKBUtxjxSrr5
JKEaQDZy+y4LHHnS3kH4r26MkpLTFe0BXUYZmAf31HA2BFYdPSj93/zYCDAXEaD5
nNc7dTpilEiKY876G6AQ9LtbRmMsm8ZeQzhO8MwQ/y0WXLPXzqjJR3NvQhU+F8Er
dUF4RDAxOCNqby3pkM/NR1tanr1H4FZJfziC14EJRkU9uvEi3ZJpsg1TohV8zU/y
LdXjVnkuwmpliUC3YBZArZrH92pK7K7aQ8g0fEihbKy40KBNGqW7avdTNWYuFOyZ
I2N57SlJNDD+gsS4j9dNCGpWYnCN/OUVa8ba4diy/ZwHjaBgUxTq/ZmsOCdms0Hn
whg1ZAiiR0YkcilMdwPlClQD+b01K79w3qFoRJ2wEOGEIOVQti0Yx/a32DM0qt80
m7m8+tBmauQOjCo/BxgwdN6bG4aACDatdyzi5KABeTUTyL1G3oYsVlxFaV13pgxR
P9l+s2IZaJE7MToKYZkmnlkC000uL6XsPf6XWZS/Qw1SSWTKgGIb//y1ksAqWsHF
hK4K0+Cw8loomnjAK9Sf+cN0i95k7JVTMIHdIuVBI/nfo7DS1N7LKdY4RoGUCJ6W
+K6RUaeEM6FPcKFAShlWF6K1of9xW3NYnZE/zDl45zm9iurUOqfr5U2o0nKuT6bK
+LQsoqsIIL43JappqoYHy91pP9xq2FU2ICVB12UwtvyfyHUAbYZVGqzaWuSWvFkU
LeRbirYdEqRkmRfqAI+UYcYk83L6kkLDRi0CkN21IeBuqKj1dFXY8fNeELFwJGLA
VlgiIXk32MtA44Nfk6LfV8PNysZ+6rpwUYV47EisJ+t7aqsLsbJrL4JBVBum7FTv
75h1UgIxcp3R7ndMkg1C9ToDyqCMiDTmBw7QLaclGhqX+whO4zHI/bEK8q0+TjTa
xeZEeEvC2WWVnl8F5VGh6Uv+E+e1dgtKeKJxduDz0NH2NV9jIPAo0LpcjF0icUXR
RmJ3tY2IbOoCmgjDXi7L2h4vyW87Khft5L6mSDnGxqQIt4PjDB71bPHKHst5aKxy
8N4278nBWskxr1GtDGEFnr1K09pFLIFaxFBh6AGLgPKnHRxvtpF/Z7pK/0wwYgIc
KpxHiI5OHRlq0xKxtHvaxkq49ie7m9htJXqWqTIHLGDq4nwE3K8HJhpP+UkuySGm
RjyJRopdb0gKam/hFHrrhbvFZK/J+s+/SEx1sYEzOrsKxKu2eNJa8tWL9ynwPBL3
iHjvh3iV0OlGzdE/ZUErr56ftMBUlQoCN/R6Nh/RDZbkpUV/6nXzrUavmFVoYI3P
RA1knrKs168zqg0/JuI7FuYqBq5dlXNPx0x0W/9jjrKKuF4TvfBU9pwK+mPYy6l1
6uVD7EGQIFm42La8d8jZGBEQVzgZ4sp0VnDbwkJghfPHSfAYLL/Sx/skV32gpRRK
jZcGYgY6seEyBLhxBawUIMLZX2JzQlUvS5FZbC8IOnJS5tuaCsyNi8LK63trWPkt
EXOLu33kHQ8c0IluExWd2F7i6oOJIO2jVrQkZ3k1uA61vdtZ5hYXKxp1dG0q1NZ6
CYh+Tmm/4iRADkzo7S46vv/p8DxH5nacWh0heH0uOsxMhNH131LrXiJcCkTogmen
96f8HaF8/uhts7FuxJJXLgJFCj1NeNIdCPah95BW04XC0x6oUmMVvxruS9osCVJX
QrzE8yzN5nLAgpUlPdyEnfcVnOkuqIHo/HHbUHj24TJ3RJVZX9xSqMqN/3MfyIfM
R0G/QIo7kXseucdl+hFNeeQ77I9mbwh4uLn9aPPjNCCnL6FMi5TkcqNrufY+5XDp
PHpw7nQ0iUhZrsQMknTvWoXxnU76V2z6mPtDqaBib9mFJTzmCaVbY0hN5ZwVv4ZW
/SrbWjuiBYH3oLwk4HwNZD3bKSapHM5fisHBbsB0gebyWBPWJt/+PkL6PB0WnUjo
VS+AZSN3uMiZJh6ItrHWiQbIn38LZFLVsx5nCJpz/a9S/0uek4AdyEv6OAGVm5rx
Us7f+7V06E4E3/OZdfMQx7RJcEb1PzyrVsqK02gT0RBTaXMv4eXxiiTlnTSpNMzW
S/Ls5i6+9bDvrq49FlctwC3HsYG1g0lCkSgvNRKe1EL9qIPR3zuX1Z4l+PxqYaF+
mXVZrzJDCwP0eZeCdjGRlLKeiZ5q4socCqsgcdFNp13BMYAAlcGaGb/TuOAbQWe7
V+CNTW+RxlyoUqM7jvJLIKUy2NkJcp326P1ltw9lG6nDjn2LA3HNJF9DXwcLinFU
I5RlebWFkJbrx9NK9t66SqZKkBWI8jNEXp7oMVc6z+dlgO3QYtf9aUDQu8+/9AuC
v0O5fgCiVYPINlGsAJ8fa19vz7bQcBRxLYZMu10tiNHJ7Vdh8etfZRiautXtPG0j
01JrlD56wBDM+3KlEBrx1i/UqRI8vtTCrFzeYbIBHgzS8J2uGUJN7ObO+7KwXV5s
GcGMFTIAcXnqxLC/yJGirdDb4V47Ky3eE7NP0FszgFmQ3beMLK2huMspb8iC4LmE
Fz5/MZMcrrsWPZGhL8ZIQuCdIdJEWm9CAEkT1yvgmYq1YgZns4zDlMCoK7oYzmDd
H9m9Hyz2SRyu4RDHL7eyNKZG1XLSK124NgqnagDNpC7r6rj3Q5a+puZzmqZ1e9FU
NVHVAOLofMSvtXk5Bljb/IXIW0TtG7H9Lmy0p/fiMpzr0zzfQNg3DEOXt8umI01C
kv6kE0BZnAKCJOAvzupLCoCIRIyXSMzr2i9Fn2OWoJyh+4fUG7PoqZPYh/SWJ4yf
SCMYlrvbc+14gdBgLzRuUSUhz5/0XineJnH9TNw5D5Ph6SB3azuHNetmxWuQl0VU
fB7oNFdXlPjQRxgjxyyLp9MRvUe05tkddvkcdMc026T6yXsGB59o7GfYOWjgyeUy
yl7tEvwn/Ebuj/1MNTM2uDsEB6R6eR7eZb/kNDZ52x4GgTO+SSyR/PXpqmLIzH46
93ANAaPEu8fL30o6m1BjA4H65gDwDdBTzJ8tjSlS0RzN9+wjVB0X8yqYrNXk2HgG
AQu65Jje/4vLdzST6LqwLPrLZluPQxZgTB5vU9K3g9AbPwXNxcN83YTt91Ndn4L1
zZY+i9tvRFoA79afuktgmUeVIHe9Bc3sj/BnK7JBUexiDLP+nQS9m5zf3IT70jal
yQ03bvz9+twIi0pu3+3xGhhBjkD4RUkBKcyF72PW26kL4l0MnxVECXehXu2CvpDp
x2Jpy+fEEA2r+EcH7wMoMnFMqvRHM4BkgnUOJwwDYmp+SemS7YxT7CgepUoGtIbs
Wv8xIeoJ81F5oOUfRjtUJD6wUT6DrEOxl2CSRrIVbwDs2Go2CYyXgSuR7nAV1Jrx
IH6ZDPEQgixrV9hl7eRj4fRE4qPpeDbYkymMP2l09YgWAxaTMw0vCP/bSMdCKwvY
DgKZbKKvxkjFSkC3eY8ZCAE11Aw2suyNVILmg8DtXPHfNKDhxSGn2Z8f8g3lDKrD
2ZQLpRiSvPsrkVgzvfH3goTZKynu4MPsytJE0/AHVxU9fxYahQMAA/WK9EPceiGs
riLC6V2YYQ87pTKhw12acoDiltnl9/0R60+vItXVAoA/9hxhtiScfMX8uwiGvVEi
zU4Oe+JdSbUHxlkqIpJAylLuAk+S4eNh54p9c4yTey8dRcZLhxeMVAHFh0NkCHI8
CY7FBj/2TzbmGiiGgIepshgILGQ5+qBIUfxbWsiPU0yTgfCZtnT78r45QXmG4MZq
T82rbfaP4HWSFVP4EHkgwaYxf6M5E/flUYIfsBAUptAFoZ7VCSKnYZMPNBZkyhJA
9LtGPZWbEHHtuiSVm/6zP5XTsEECzBEcWEYZ0Q8VODw2YvdKcjvQmd79qciI+nyg
0GT9Lr/Tqd/wXb4t0AZLje2BbwmJMUCTRnMc/Zg3dqzhEhYG5025BGL5o1YHtUzF
lzKemyO9CGMe6fEi3eb8sBAj9dEYXt4gj4NMeMZmrJwsOWUP76bBBbeEuN27+kqc
4SNduBpFcqblAlrt4TqU63+O/F72YvlYbp7fzmDUnBJvQL54u5iRxt0knHwJShvV
QQTPuuUPH1AV0Rj8pQ4Qxm9Aqq4AWdnnpmnJND8/t7HMkvuBAzOtVzFmvo+62/pT
WulyZgQ0pyBSvXc7dPHKqRScZZ5m1flZTy8Dp+Jp6VTk9my0G3eFMpwIB/qKeHZR
H63SuQLO6kj6m0qP8/+u/B+W2h+2+tpibS7M9Ju5xAqAn/PnVYqe8IusVI4W6U3V
4CyFubNeAxihY7iRiwxwx7yqZiUHUx6QT3txSmtsHFhFuypGOA/XSlslI5q0cO0Z
hVNjOic2T9X9Pr5RBm8trkVo/oLgnFSxPxwQRjiJdMYw+yBcGX2EvtKk4Q5J08PK
jn3Y1fVeX4IWtNMMDBb2qknvkLHRdpPq9djWENWGKW6bE4XlyHScL+yTRKm9pyQE
45SpeRsGIRCw244SZ0vapwsGuxylgDVKGX2shpAZD4En8ZaFpGT2tetzGNAj/69N
bpD62S0UEgdizQpnGCYAsrnR+XpiMnibyk+JyN7cVJeHlFpzVBRFiW/YnK9nnSBf
lqivHbjZLhtb3pS226cFYhWfjPcWhXQJ7G3illfL1gSoanAJJEsXf0GW7KyY2inU
4fKgAmXyMRlYuW+Rz4p1oJDMIW5oMEYZCBBkPoYLxAEOnhhAN7DFM5AV/tfnGcno
3/dnsatvKHqGQiyIOJTBAxyQwhios7B8IIgnv4Xxpu97p6ZO2X+7yXhMuAWwEoD5
x8mfHRgnrhuCDAruykhiTPTd0EtfAim6UQGOajlIf98umgjzivPZ5RHLEn3A+zNf
KFdmOfUAqJzUeTKHtSz4U3o5itFhp17IEuO80y1KEdoEnbE0dZsFcLoMyB8ajl14
/2X1+B2Md6tBwsVSJVAgjI6+i5SA3YqlaSYC2MUCGqdrWkirN8X1LgpwQJq612dl
uNL1xUYfo19KsxubQK1Pcpvy36V0Y4CisW+yMD06qYx0B+siWq2cZz6QKc4FLTHK
JuEBoAN7zDOHLJypbBQWrnRy4BFGQlTxLWRwjoFljm2zycJckwGZ5vow6NHHp/+I
PUEYPRUOp32heHp2kQjb4kYafOe+2cQGVA8LFHG5itJq+lVrt1VXUkbAf9tfCqL7
lS+gnuUQg7uOFeR195MSkh+MAW3u5vNATGB850KnEB3zyQ/+kFUQV6NY4H6C2AUk
1f2ORbfoJPP6UuYMQbH0NAVPT7YI5WMR90OXoq5XKs9cBboC2cHanMPMVULjYiUG
OIag9Em1dqZdS2WFPLJWnsjZobPIoa8m0wF7yKbRUs4CwPz7ypZWRas+erK5oPsV
erM6V9TplYRu3p+QYN2e5R5dcYdh5uJjFIKH09THrOQ4L9i9RIDm+OD7730z0k3a
kXwZHmLyv3dmhv26SOmnmZEyPz2ePCXP9DAs8X2nkdf/u7sIJc7YiPsLvV9MBeuw
CD5fBl+QZ+jGjBzW8xiM03ZOGNr3m+ly0sRER9USq1MsPuSlHh6mD5SsO2PDP7fJ
GrwvxmRBC+VfZXWNPxd5dBUSYcf2quFZa/1tTvnoK0wMy3ve2Fxejl5UA8ZKYZ6p
je7ZNr08AC34pBKwwB7BV1Zcchc/3/xTgZFRAQ1UXvjAcVkGSp/jM40jKDzGKuwi
LwbUK5SMd/2VysOIBm8CtNQq8xyDsVqMQOOIu3X9sTs7tBqUSIeTyLQK35R4gdaz
sUwGDccBtpy3zyox2DYEXiXzzXrmzDHJUfVOYjkF2F7vh7anT40NBGyI2XhHOeI3
mW8VlmYnc+hkhQX+CYz/TbQptMHbfHZiFG5WZ6g4opbyEwDn6p1GvYEiYREfhkHi
+XDVOaDvH1SrmVz9SBW9W94IkuhVrO8lAzTGdRwyBHQ8IT2hjS5tyUcKxGp3MYlN
weqZhfIsLco9riQM1PIe8+hi+sHG351w1QVGcNBQndu9tfKi5gcqXIItw+LSqscu
04BBgzPtES8lgfzfzXwDk8vjsdfAfRgpxAKlzf34cgkHEY9O9N9j6bp/S+pHv4IW
vKeORx8Tm5o6dZ/dug3s05b4GwMghelc/QA9Ej5dvwTkSPv7zQNOXt0cMkKEpojR
gG9fyPUXszloPkLG2OiDbjaZlNTbm9/+RiH7CzijgnWSe/U6xjp64qrJ+ScV0R+A
Xr0ZRSFym6CjYLDUm7K9IRfzZCD2L6+fiDU4Umq8xaIkDKe9zUT/GkSbldiIi7ig
ACBu8CaON5yUkDyAIfwJ5pBnBN9CUou5yfrYY+VrAsng9xwBOl8Dxh6xUBx4aFBx
lTSKA6oI0QhS+NxbVKx+Nu7ZaXtUZURuFyycNydiAghengvegortcKr00xmZygu9
xhxewb2p1D0oQfkjg/iRtbgo5UO+Ya2wVk7i7zej9OZ8lUvoFgYgWpfBKgoPvx3R
2rKKNu5RJqZn2J1emE0AfPfDkgSdr/9DwTT/rJB7lLGRi5sgG/G1+/xmkVSNIwy+
WGfk/8ghGRWxhq7azAs0wbLLo8CRSAg4n0S2EahsyuKET7joYX4Nh1ziGZYX/Koa
Is2CM6UK4oc2a8MpDqw4IILJNmW16Udch1VKshU6XD7TWkfiscTShFjqbrmU/MOS
e43O+Zs3qoqlRx3w6Nq9u8MALDlErDwYQGzoJe0mCmZhe1x22osWjqeE7PWkiuyF
pwGXLDAghxesgietVR2tY8nHIql0KqvZHVgg6uv8NQCnvZpNBh08glZBbin4V8t6
iR93+J49nqkMco79S8NWDJHtJDBe6elXVAXZ07FAkQijJDu759as0bZsvgJUcTab
ncxxIP5GMb3DUq7NqUBtvp40YLOCt+vJZcqteXG4VCIk41OyCsTdAVaDYyqXkcfM
F/INE8yKYRRuruQ/c4O1UDm2AQsehIpkX8RSlGgFsBXdZBBaZI7SYsKXnqftaO17
QhdJqr9s6pCVo8KoXgZv0Q25kZgWmvVW5nERVj+m+uVafDgEnGlnxpHz7AbE3Jy+
P/Z0aV5uebNpqaiAh7LMqW9V+L42ZsxiIuTmqctQ3cg36osT/PpHLz2PTnvMtAHU
1gdUet1sEVjZRis23PWPSM1NGwhuIHcnDtwSSHC+fpGqd2yOnZlUuVWly95+LeKV
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16560 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aYEGshOCBNLOAFPz/YVL0JBBnwIH1JW4SjgkrNQLs/u0
yafk0N4Q1ysmYyE+LKpnxN4+EVhVIFVGZtmJcJK2Qg+muWxLE5FtrKORNpgjaNCx
j3o10sQg575pcvUW4+8uOY7wulrWuCkMCRjWRQRjCIkanSLXluGQuQRIrLLfzp+U
sGBuJAQSaPI0kOVa5gau2kXTj2AodsqUc0/8YwqV7zWCSTDSQRH0Pxp74JT8Cp1o
jDtLxkmeq4I5o/zbyRJEgcuQD+GsyEPrByxLGhekzuAS4cEMwEviFVk1WaLj9LH+
3tpv5a6ODlfkObTAqMhbSPaoV7XZoQ499l1XK4CbywW7nKYNYDP7vG9mJPUxySmG
Kp3nCES1zyfAqxW43STStf4iyGt5SEAhKCFZXg+C1GhIo9y57FVl64XdGsxHStM8
YATdlFgFfqRQ7CWQ5Jy+itt50fcRIGhhZORmRpxKnUSFrbJ2EG1+h+Tj0QM1s/SV
grFREPa+o3LMViWqkV5gJvy5TEl+thdxWGWi44pz8iVzbwAf9Rzpsv+jkAkxIpFK
0KXiorJgTKIRRATCZE3add8cwHs8jvEMOFpH1ETsTlv7bx8bTmBj0M94AwZUC5xz
xgB8zSFPeagipiNSWe/e0vxP+S6/8g7aX0D6PtGwCfHV+4TzBFAslPo+3fSXC9D5
AVhuQrYRyeg5uXZUqbnIsV8Gh5FQgmtOrBBu8GYRv3l0IYnwFIYVuhklPlpOhmTg
4M4IdO4emaZD4PPhzCJOTn/LbdlajB753rPYrBF07eQ0SlhgmTVKCV7ptOAIthfs
FflsIM/aUjxrNZF2RcWHDYeiPqAuxC33IxPJGwOy8VPsjXc3vZVYryCgyXznjlTr
cFi1w5ZH/JrWIPw+BchVh0beFh5QApNDON5Ml6WsfV7DSfaHrhzpyBIbGy7gxmu0
moUr/KzzTtqXmfoMLZSsvm2vV99Se3WdKXmBvYkQjY4YL6hlwHLhPliu9wXi4zJs
X7aFRC4AtxpmQRNSPLOrrQjBvuQRgUDZEwEPpB57v4/Roqxby/IaG/rii9QzmOhk
8FrqwhK7ZyAImYqGnGW6TIXqxBAeSvpXW2GwykgX7C+I1QVn3ZVtzUjtUcO/A0k7
1BZxVRdLNsTEPRxClbGHtashO2M2JlShh/PARiOOupVcMtqpZhC7TK4gKMdSylXR
zp7U/Uujf9ySW1awAmsmN7cE5hwuBwRSr5Tdku0NnHQTc54SdrPLNrxk/ZM6RoTf
i+Y6P+iDPEPU3w+i6ObrrGPiO3qoR+oxF8CbN5zZZuaZWhlN/w/TVIejQ5DU0aHS
r5J3k5LaWbDTB24S8lEXDXqYDbgBbDGVB1QcCmwk+zTQYmbcdJIPOQeFs57fIaQg
Wvj3a5QiwvoaswipGxHjLuHaBBd+hPUkYmgcjrW/CL4t+pfyp6hPDU8Vj5iTv3EE
pyv8bzFp6cNUWddxgItfocLBzr/RRQQptohL7J2qhWwy4KeDa3+N0xn20M9Pb+wg
ZBm4IgV6rWlncbMRN99KNKTBoZYlH5Iic6dw0MMIrkcbw01Y9VyBKu3AbF4r9l1Q
gLX3YIBFUfZ5oTZCOdPvkYyEwtWoD1BjkTZdwZpgvdkGJD5vYwAxqNsEteXjKcVv
+vrfNOea7hdtLdW/gOJdqLeGZUtIUMLtXbzxnEwHasxTFvbvwN+rUlA23Dhfa3tm
aSpNT1xj7qmXQwGLOqG1TYB3WlpArlOdmfpT5eTm5E8iaIZZUkybYBfXXZePQD9n
oMvkQacjkyihISnZXykWnSBXjtlJWMHfvEwzKkimCiaNFuuSwU7fzwa4uTONm5+q
8PSnOE5IoPX3iH7wECBbR3IssCjU5YbRDiIqQZnQKi8gMWuTjkOlcJpcAv1qYMcT
jGP75l8nlrwY72A2AdgKosOE5dhMmbiW/L0sCz7xaEnvX7lkGmf91bFbTAMR4Ux2
TbgDXExKa1r9ZZPa2NvOEkOHfWsMU6SUVXVTwjD/sTBVjxxO/8OhhIOxX6jXfUZx
/kmXfyVU2RGsb2/ZKqsmNEr1yZdZaM6/SAUH4ddldPe2rPi9/z4EkxVAQUVtCXCa
2RE4mt/L2G8Ui02vn0YF5L5UY7kDUYiIgUhjmxPoPOgljheURujoauIBpH9XOuCR
HQ2AdaMmbFxuiqY7WKpRG95GjU7V/BujOcMRGb2luBR6PI4MCBaHKagFZ+aS4Xtl
TTW4zGe7VNk70VjBXwWpHy++QNzKUrGWBdwY2b6MTr//2+n0XNYOexbgge1LwmyW
XFzV03+dYU3tTqzfUBafs62xCxCD40jigDTWeKQhIiJoWasiI5boTU24KoNrbmLP
H4c3ZZC8jDmttA4ZbIacjzoBJOqgJfDik0FHbvuLYeY+H1tzfStUrP9/0sRx62u+
IwmhExqDhMEBqxvgBCLEx8qKqYVP5LwRU42ufvTfg1QbHjc/s1VGsH/W06WShGjf
FygCsPqjsBeEF7ehNK2osnkppGCiK4uBnuNA0aBhQkZdVJumUry/LZ3oIECovrS9
b04/nJwUTuzaJFBrk2zVsoSJDNJOKQrHTRQhGhV3S24SS+LwKF48JIGQyL+FO4K5
Mvj935wzPGg1vpqE2yE0xyKwspFeeoTi5a7ohF2jetTIh65cUw/TU0saFHBFU8Jw
vh1IlX0u4bP+f30LZlc++3OOeMwsGOM8MAztnp429Gw2hIu5MKDajDFJTt+RI833
pQOrbSu/CDUosCxCVar5dounSUhjMmxQV/2/faTAMqZr5lZlVBmiC9En3VCmxynT
zfX9gPctEQ9G2BMVeGtlzKGWSFymr4dRwny05IVFU2mX8zBWDJQuSIdkutcl4Rze
mfxp5KibDv3SsFnwDT6JCvhS4ldW4PJ5THj4qtF+xLSS8708+tnnq7glTjV+cKh4
sgZz2+LRDJq++9aljqDRFN8Duktl739nw2jB+W3D8LtsF/5PaoWhGfZwpwhw73f6
xntYhV39iI8jaVt7WK+cmRDNNxoxtJmPZw2lPAoiixz0HRXaIKsjgufafu2ekR81
6/SpJqoiUM8d+D+U2h5w1/gDvOst91rNXNTQ+FF6W9jiebK/De7tpG6ervp1zkV7
dI2zUs6BEEIWI2FeFf3j79v2+Q2urwkeEvUJDieiUIzZ27UPxHrWWaTgV6n1/eAF
imVSSoJrgTOjAin1EWfRnvTM1N+4GI1e9S9K5E8uReZQ7Wyz+EYtTGkuSh4Os91m
MTibhduaLMjuMwU7frAj4rJInY6gxWfuQUewC/cDn2TtwCuhhpGZSv3iYJCJG0v8
VZQmxww/hbAKsdsFM0GuOKSFlo7yY0pPlirtZfd8jR0CSlBPVdkXdQlBhfYo2QEF
e5+c6MIx8j49ZtZyFiAK5blL4ygH7zlCuEwWRoOOO7BrwN38F2VnWElpKSCwEE3n
fY2cYgfllvkXntP88YZ592haQpdM4PT5l5u6xKepqdRC6rYHDC52OMUcL5rxfF5n
idYh75V5IX+6wlA6FskbpCAE2hMO5NCf+m2US4H8ZDvGxBedt0MLWN8D8meBx/U7
aR4Vn38wcGaBAE1SQmn9SC0sPfU04ZP7Rrad5mnsUtjwM0fMPSniDJZhxc8j0OlY
l5FFpZODRH5cxuBGH5lvOR7a96eqLOZ8jVgfLObwux/CuUge8DLhycB+T/a0vMV4
lVSYLGK4cVY/KC4l6NzUfe1aeB+aBvQF6bT6DloQIHWL2IwBDaiIBcsCvN8UpNvH
/osGgLyckbCuuznBAt7qialgB8f7vF4dFupmRpGjTgZXDlJ+GyUsRdw/oMiyRMPv
878B0kgOJLLft/vlKhwp/ypfQ/KGqltt96mKuOS0+bAErPvCSTJOat5PhFFoepnN
oXm1qnwnAhlI7uQsXYspaRJyf2oiAf8+U3oBu8EbF3yPApzIxCBL5wMG8WqzMUVm
EbSMGxa+oVcFVNQWmk/dqvPLM3zkpKjWQmiH1W9affQiSYsPUgR8q8TQkFkS6WvJ
aU/f8muqHpu1uqumYVHO4+F0Jzot6zzHfIqfoOflAGx7UX3uGcCtF0DM2VBQAhp+
pemeiD14XZTt70zUtku4Ycc+mz8uB+D9A1MNljRPV4RRPuNz65P622gsqvUacWu6
/mLhxGTLbZejPt8HvxPNMTu2v/xffS0g3L8v+EU87dvcbXAjARsVVqBUnq+ohWbK
O9AkxwhTeh9p+UIHfS6TH7c/55QZlA6QhFvmqLezkqUJbtsk6XFByEx4mW71AyIZ
1dLmAmrG7NjtSHebovwvv2BDfztlGxeWeaGHeALt+Yc9u4E7uNgW5zwYWFQUXEzk
84UvOr6mjIxxbEV3xNqvjQJNSScktnq6UuaYlLisky2t5TKip/TFArD0aKY8jawX
x8uyA3YhThaul/pQoxnMDU3s8QqEwN+lbGVSExAvMjh0sU5xVN8nrbFb+5bg8J25
dNrhNS9FNgoKXEhfcRTtra2bIyBAiYrwB3+eOvVvRnZNRqAcS4DBDEqxWpQtmQPU
JgnF33/UGwZ/LYsSzVHlZ4XIhzcB9D2bjK1IxeF2BFzjL9001wJ3RR546acGFAfR
Wg1eNlWH+ed+9reAEPh27L3Sis29b2xSdp+w9GZYnfRWQ3KSPJV67WlG357h133V
c9wKpSj0Mi06p4yDdtazyCbWP1banmKpqwgFL2GNC/BGQtiDIi7x37TOURAZD48K
yMge5Yph1xM1qQMhwdSRuYNpcgO56fDnmsgP5isAVFbilGq9f7RLo78eH3ruPQOL
h7Fo8bcgAL2KCYUbHtVbL4gOEeIcFiEfBU5Cgo23vrbBhKnXs1T27we/hyUDygSt
Ru4reC5E7EOTob4uREuxYj+7vMnA5ot27z90Wk7Djo7E+JxkfrEVuz+uoKHJXjrF
hNQIuEKspyd2/OluJ+RxRwnfn0HpHf2DldkL8QN4b6dT02aus8UI5Gs1EdhHl2RY
cKaNl2mVVf86icFKsgOEE/hlzkWlG2c/pDYkTYUzNVFtXk0rWD8WcOiMa8raG/ST
ELP4lFYTjr8fDJb5Rr/L4F6Sd52jyjioBe6HaQZ5JImjXtU/6JUE9SswzstsoOj0
l8laSZO62zHtIUQqchPii+8d5q7dMgOpvsAN8L8sJkMJHgiF1vjm8ENCA1KHxAA7
Ebqtaj5/JkorxVEDwKuEh7YOMZnB7HWsTI219Weyf0Hn5YslX7ifXAbGNJzlSszd
J5kbLkBxHqL82D2Y+W7X3NpH+yZr+4cYBygCT9KChVnodiE92+wcgtgXSQszHGlV
3T/Cjt6JKj1VqlVe7AH1XFZ2gH/74v1DToCzSdpdxunkTILsjDmf9sbneQ+kaBFJ
u2F9zjccCLZze2yxf72bib1VRygL+H9dqorrGSEyySY9HqXYKVLL+HPV0kMy5ETK
prjUxP7CjB4SaAF0IwjXCqW01a+HR+ykOy8XUIfk4NrY8LfVsQFN/4zJy69xRNlN
hoUKt5cuIAKvyNPKz8Lig4A3C+6o3RpTT292kgIH2je5kFTcBccJPmaAXzETglH4
HHQGlQ9Z3VBqKNosijagN+qObjILtGsYv+jgdQBTq9TBxSWU2Ibv507w12mv1ach
CV+/NC8C+lYmCogJ1HyHyb2GoKA0v58qWHlPET5cQHX7W0ChuGuTA7baKPqKzqWW
32agb6bT3hCHBggDBlROMsQFB0DqQiAZP853R+vN16ALPuUNY6lcOyLvYuJhVTYP
u5Qoo2kWaVBg/8pDkO1ULIum5zPdieccJfUgVCziEt++siD+2JEGJERVpFYITVdq
gYsGUzM9e565J7KxZX9F+jwcJadhIW29mlNc1AEs0axHV9rL+Dl8YZMM9cmqHRAv
q0mXc0078I7CpHn4v//yl1k+uMy/aVa5WzT4RpRVWPfGaubCFz2Jn31AN+a7RwBm
2ar2dHDCgXP4iM+X4TYpc/K59jbMyeoEg3y+t9+OK/WFdOsMQ2ojkYMQ2McX8CDK
iWOGBHYSigR8WniJQhQxTVsZpi9dlLM3dGYZ00xwPk0goJkSXcW+wDwHIyUV3rUh
m3HxAL2BwQRVwOU0fKEHWIQai7KOyj03d9HYTOnxkKZJcb/ru+DLUg6t3SFfBjZq
3zbfFYeXjhs+0u8YG9ssHTGke8LSQtFy4j8YxugQfvciV74m4BWbiq09S1BjAqzk
MAYxU3cEnmTkIaZUQp4LuRkW/1Y0jJmFXRgtDAH3vheXPXH/qjIg9f6A+lJKI+v4
BYW7lroyCrVmUyYimvZhiGYtLPKdmkpr7X46/1XqHcbPSjG5vg6SejsjtcfhR5J4
bD0JQ2xIu4/ZAeyFuVnnMa6MTVjxeO/kmdNWFmghzSvYpK4GYDt82ed3qwjqzdi0
oCktUMPE2uuEnfqiydjlziRBdQR5GPb8hKssS2uTjnDgoKRkG7ZKzhPowv/hD5vP
Dbv1zDa+xCEE1Od3SA8INmTZZRKQSIcfIl3Hl6NAqPre0EX85CntTDmlrjz8xCAc
6NvyIyvZCjqEGHt9Ia8YYlFy/m7RlSpqP7/I2AbxYE+nQteHI+RHo5RHtSZpB6a8
WnwMR5E4xF01gMQugL04tPgLxiHmrCeokmWHVNnl09+utZhHB7//es56Od7VQ0U3
XULOgr0HFJrVnVa+fUlfeRDkxPevT8XxzX1ulOddCzjcyZp7jdpHIdMWCE+8pd3a
U7QeWbHtWmHV+wXJGgDACyFOjQpp24pxvmBVkVhVx1bSSSe39KSZeL9EGvL99Kyh
RTaLJlhQ093XD+GEqkEFT+kTaN8T/snx3Lv6PlDrgkjprlrl5iwo8odnXgH9nJSU
wzt0tHMxiRmO8qCejTNsrteg9W6ORdaPOV7Q8IsX7Nmc2mgNTgzf/fHCWFSKoosM
sMz1CX1tdqT8GD/MxrS+UjZJz6+cEvKyRwzquPtfOackerrbr6rEVZ/WARQ85kGp
O2MW87sJTiCqk0IHlRKgB/ZafrNRi703yId93JiUQ0LPm2TZnmGzNnAg2mt4ubKz
3ZViV/vW1sKgFdkqEflmM0WJvu817yZydAFB7Zmp8S9BejlChixmiRCjSsO/3rhc
y2GKgyKHH6q35p+JNLaOA64Z6kYZ3gtGpQPp6OZ1TLNKegZjYUAXmz+3kh9BCZJF
/x0x15xuTDqZ2m1/FMRQcWeKSw2ozAS/wLrlJfIjRn1E/HCQSwzubSCRDtGJ8gPK
rw0sh9GYZoPkZdjwhwbLVQQn2khMOoZzgjG8vMjhDwMEhh2uUXVWTXDdGhJtkT6M
wTvRYK+wT8jov1Y1rvgdnWQGwAPcXbfAjlnwmRTfqNJ/auW1700GEas3DwOWPtrl
J/gdqLbS7fB9FSiQZCXg2bpOqMaQ8TRZu7Z4EI5mHK82I9pksQSECP9yhS4cZjK0
autZUfYPAzZVYV8tbPa4hrGgu4UAeMIkHF+oHw7860CRgVjFKpm1GfR9jXH95xJZ
08o5Dj3s6szQ8TZydehRdAx2pOvjBf5tyGq0j8W+uvxfXMUtSkWUiQE6T5U/qH0q
HxZxgqJtlI4fysa9zUVOaefI5fUOwipBQ2KAHmHQ/Q4zK4kVnCv+8NowVzFnTD0B
z4ajGOLrEu4e/aT+AohPBgYScs9yQl36yNrfWBR6GHfCSn7dKv6Zs77u/05x9mLf
tlFGWmM7LeBPXp6kpM9EYIimLdWAsldewcazCoCBWUk/6FFfpG8f2TVk57eYF7w0
r9gaJhgq6Wm9gPK4z83O798AWlgn4LiMdbBbRROsJo1Xl0RdrBaRJBvSS6mr4WR5
ZLQ/H2WsFTvrRPaaw29iopK9Vd7rnxYerXC1LVsGUFS4t3hQjalZtje51jhYzp+W
Ncqlt1SW2LGInrg4DHCHaoi1Ys/34a0fUNICjOSxJ4zAmOViRSPfWzcGHjUiiZin
C3y3Ril1i148zacArKiwkN88+1kszYXwn7jKnqt0GzVnDarZptkQNUSJHe/VEX/o
SXRmur45TOZE3BnmT7KAhSXQCtzqyG97QidWTD46DMefBBVfHLJ2olmiM0EKPqIx
LIGYFSMamxdQRheo/8shYuMkIp4YpTD7NSCRLFxrU3WeZX2ibDujRahXNW0TiZ78
Q9+/lmYlNFU3wzL3OrK4U8rctMEIHwam+xSeKaPKBkZOmgk5xLflL8lFPx2sZlvj
CrcYLJ6Rrfvl/siy/Aju3SaC2JU/JgYedUUA+fQ4ifRk9QQl6b+x1GfGZJhy/+rs
t54TY+zFyZxu1Qo8R/0sW8TOhj6DxcBe7nBlPhjYaxWfK3i3uym1G9bQLvfKzgfL
G0S16lrfKehoAR8LU7aogPNb+0Mj934NDhfwJpLCN8DmJte6wB73TkN2E122geRj
C2LH+eEvmVwU4/Fn4LIm8I3NXgOr7oyA56MCj6G8O3s0YMRALbjHNOFVNe6jOL/Y
mE2U8H4EETG+P0d6pKReqMzlSeVWsRFxenSfjzgDph726fTXhv4un9amnHepBfux
4ZsSSKcylqoSrD83MxJ08xrsnMaEyfCZaHLSc53qjRe6M++WYUfMUqukIzcnf4iW
nGgn+YjbeuulUppZ4EEJM1GnfbiF+xa9kqEwwZ44vUiuj0LRuBN3OdVvJNxOWZC3
gU3Nd3gLR8kMTGhwUAW/L3hGfhgsXP9iVsbypNqYHz2P0fbm7SNLjGp+ixBlOZcv
BvGeZ9bArA84I3gIUeNBvYsgR5aprbi4AV+Q6lPhyFYRRV5fdeMu8m5p6Dt2pzIR
euDfyJwAYaUp/f989BISvg/22OHYaxdxpBV28QZVJOqZ69RWYZoLSC/+exBzRW74
k+hA68weSp602/Gx32onpMydUFg7gfO19966UR/tgfr36s2TFRH7BuAMj2ge4DA+
og7Lbd+xlIYCOXk8URkYnXd94IY0VfxAfDaDv91Hs7QXQuaJyPwW5gH68QyQ8Op+
tJjxbFDlXm3wKa6ZNTg+R39/NG/r7W71eUfc+PQqHld8l3DlPPXxnLRM2UOtoUm4
IbVzVa7Zcg9uk7p2xTiU3kBidqc2o+hH2NXbwVeARHHyIb2tlxGU/Lmh7WSxylI0
XzL0y1f/9lBeMPnkPZkbJRuitjWjDPHSdwaAJdMQj09ztEO+8cJHt2QoudJX1nm+
xPejSk3TQaHKdkIwAU8Q05NucH5gp3afHCCZS4PVETdf7r+z7CFyBeoXXrLDrQ/W
oSB9IhQghDvdZmiftgRbBBfAjtNCPmQT88pjajntkMozGJ8Sh5Hi46oplZMKaKtn
VbNd1JYudlmVG5Zb4d2CN1VGnuLuGDEzD1yRN3vACNSvfgHDIbIrS5mFZt/VwwDv
lLLS+0wL1fzhCHJzG+yawmnZBSOa9T2XF6lZryQ7gG619u2bnA3RMvkJuyKKLQ1t
8r6/7THb+688M2/Pyj+dt8maKVs/oZjwmMf9qvYksUAge1kYWfbQYbzXxUb1pKxM
GdANQDJ5yNlXeUHe1C7XpljTtkbU69Nn+h3fMWlJFkTh+v0w0hBGdr0yN5kE5Rl8
7aoxbY61/c66T8b6+2X4m8RBWq9ofzqGR1WRml5Y3bJeLCW7/SCswG1MOu2NQeDa
nGKwAlwEwMHuCiNZ5vsVdcjJ5OXJZUYgCs/sMvX3S9Ka8vJeUUa20zoOVey81oo/
Peq7rCzCVlRQ0Yxu3zRSM63dtI2xExGb0fIfL6qLbV2IITL6o9zVojGT+9cdVD6N
n9ma+kEor42WDcPhAuQdRMnyrCGRHIJ5xJw7BlEke7LcWH3dQIVj6oA17plUb+Fi
2oLdVdWp3S1v20LPDsAYIrXjdCfJxO0+tnS+czNI16xGdHVvbV2R6mY1giiZpf78
giyojixhYYedS4K9og4tf/BhJbC/RTMGQN4fNYd7Bdw4GOE0fSU0hAxLhO9LZtXD
JHvGp+rAbopT8tAc8jrofd7rmWVexgLrPUle/4KCzjxYn5/qlrRCyQzkZeI/AZKe
dRQR+wmORJUjJVaNKStwMUotxWL5te6U6XoytQ6T2OId2sve+zY3/5SmbW3YGh1y
FYGcxFuMqKbUy10h69KfLu3GYC6A3eCi1FBHei7v4HVYBUd9mTsFkJBiKI3KUHUI
JZlciX+ucFx95h6nk/EOo2FKB4xQIdwthq5b/iWPnG3E6ojcUIRueSY/3ZoGkkVq
XjmEB72Lv3j4sz1Zvq+cDb/Z8TUSbtyrwOgZ7IYYWaoZICJb4nxXBlQmywLZ+9vZ
08shv2Cu1EccZQIEsWGMuxDFhSW3OCeC31US2g09qhh4QkOa0dKo3zj/G8y4RNsv
FZMEKb/nXQTI9BGEbVXPD9TIidnjgFP2LW2tENFBg2hawIeWg57OWLQU1QOa+oEX
iZcaOFGHwHS+nu945ATCHGWBi8Gwca8g+FwcuYupjitCb0Yc8cqqbBmlGQmRktvQ
/VKi5n1kIVNWY8cUl6t5TN6xmkEdQAkpmYBGpXwnh5hRiooFWdIDRsTjaifzJ7F8
Om9uApk2SJI2KLpHsukCCoeCfX2UnoU2aBRbezk/vWXMUhUDMeZftlY5LbhVZMGr
eaenTB0Fqtap+uRJ4+KEgIxUD7xv1FOVdYmTeFmdvv0Cl+ixkHMpha8lKaCGRdpr
aHVESPmfJY4CUtGVzZg+37EqUtCmtOJJNthvNwHcUnRnGq6sa1Uqz8DCZ9nsAxnm
YzS+FO+LVJW145xy3ls1vgDzLjjffp9Bcb4ZFh9waP284fEf4VkR7wUaiuU1z4gi
BdKcmNebe+NRkWjNA/Y5EcEqXeS158iXjsRkxQNiiq0Xib3mvKFMXm5V7pkTUpsq
UCkglWBLhvU+aMV13QieRKtHJw+UfAYp1jCakbxFOPG94HYxzpxa7a4yqYY5uhYg
8Hz5C5GwEVfJT9rQ11NrKPnFOdHnBQ4Yzt05PDFdqkljdx3RzRYBtc7DVo4ylCsK
shuYSRKy/HNsQYmHGelZENZmir35cA8n9zKI6xEvn88YNHRvCBCqWzDmiJttXy3t
8TTAESBZEJby05F5UBgdSkKqBQbT+sGSK0jmXSEOeuFJNFUISUMXpq8xdpbqI3TM
T8nRDqb//F2td8JkdB7cN8H8d1zgxIoU/Hm3rbvRiForQBG8umhC2gc3fyioNP27
uqWMLp5hjDIJp5+qZxRLfuG5ZCwhTzZsB6i+c1/sFYipZ7eFpn2Eb3FtAtL4VspO
kK4b4+eAblmCCuYYc9WOQfrTKdT55nAKwGZeHcfMAtiEdcdxWg3dRHgzrGGyjrGO
HJf6bLxqFGRSQJXeYicWkSPgmtLnSNcEewinIkgM3Bd9Gcb42nxelkD8YaNgH5Jg
dEwy80b4dCZ6Fj8/m8vhffocDiugr3wzps6C95spoU9GBrODHnE5v5aU12rCbpXK
ZnXjre+1nkO8f+P2FIJHDQBb+J/bSj45e+lQRNiPYiunk0mirdYmVMNYJ+YehE4c
yRwclZZC8zppY5oEpN7/yRKw1yV67Luq/gIH32IeliYn5c+K1dDEeYF01koP4Tsd
1CV4u6NJ1tNVK8VAd8g3/c61/7AwhFDg/m3EMCCAoBBbEkQO0hAMSRhLPSHlrIPW
YzGsu5rRdKJ0y6ZKNW7+giQh9dOp/XrUh9ABpikiZF8/YFqjUO6JtXydVtLpUZYY
owV9fvc/RtNyN8sPQkVEQeak5/F40zPCYw6uukp/pFJIi4qved8DUcI+12+suu11
bWPU8jNREwEbVpQLSJR+QHEBdGKPlp1Nu1nfD04UrFsxEla4QOvpUaMFaG1dAoL4
8eFKcM+VI1T1HyHemMiLhPTVVo2zk9vnYfmYiiY9O5xi1hNxqdM67bxbkIHt5MdH
T1TWKzf0uP0VHJwOcGh3qYkz53sKwVhKgimUHGzU+JiZLMNjPEKOlswvuNE+XmVN
pEwblFQzqvBAwK0dLqTuVOvCpm4vXTPNUulJmlHiBkAtk+V8OyuXBntl5aeBlhzC
39cG6I3HpslByJBLG11VsYRYQBvrGh9XjU2+QjfXyG+f9MbQNQdObtMTSB7e77HG
HTi/mWzfUGI3UQ4VvFBznvIhP9UF2242FwSi8/Tvr8Gk8gMJg2boOewXDgUkt9RV
k/AZ06F3ZH+xK4giVQyXFZ/p+3uUoeEXwajpvLqcX1tt4kCcgBQ7OztySwhv5Fep
zxS3luQujx76dIC9nSK27jFvrgXzkjXzCOP0iblLjb5Na1xf6OPJIp9838gEPKz7
p50WmXydW/EILXgMNvFibgugBQvn6tT/QeroBgC9OWsFnOAqTcBZs4UhrT2mAG4B
3zYsM6iquB07ycI4YFQEYnkIkrrYbr9NdaOEfob7q6mK3jS5pEL1dbHd2zJkkLV4
IokVjgrpcTvvH+As6EyEVkSL095za2rJjPpfB+L/2Y6rKrlN/M1aMXVFXvDdZvnl
SdctUEvKjV1b35CJS/wzPvOfROxAsD6n0ZE+HBe8Y8QXC+9HM3P/l9GLdn4Lsnul
UODiQfMah11p3RmYX5MZ55DilK7U15wsLQ604u/kiulQd2gbHpX3i1RGROmCi+Vo
oxvKcb2ZSD+/t02EavO903MFT/B36B762m0bEpOfjUgBcu7o8ypfqhYuz0gP5ShP
Z4jMeqIdyyMfqMi8o6ET3WjAvV6sAQjAICQFq0bCw6vVMtDo/3EI60U2ruqz/c6Y
XE3qtr9Y3ig47518ZdbJo07NpFHb22Zl6P0FAsz1T/4Z6WgKMBQJtCFaf7U0p4yP
JF1T4BOGKaFZgLNTEvYqcEhySxMDqiTK6oc9IjJioIm/xOm7jn/jf0dDAfDUvdNu
gntkihQPYesGUY5QjYgULvpK2KoJQz14+md0AGKC7Ri6137kP3w0av/POTDw5kmE
HWX/r1ssKMs33LCxFV8wte8D5vDCu8alGmwADjPH58x1RcWU04HoZSausDW0DC+J
IB4QZWWiCjll+Rpxkz1+/3AUe+NagLj6j6TbZQjctjkQ3QTg/U1rEOPHPwq+mRwl
im8hW9wOhpzHe0J71n43Shs1Xc3Rk/o0drcbxxvj5eQm1jiegIEnbmvRfqvVQB+p
kWOcV2w59/NzmeB18YRFkbUwp+RGPsoQHf5HI3RFWtHtUtJonOLx8PyffFHnzYGU
EITmYQ9+KSTMjzvaL7mgzmdh8DW3NHJcgx3oRZ1R2symlE5Y8W4sha+We39AXOlr
/7mqdNMx8YmIn07eg2z2BaOSg8GkwEtpl3ssTg8t3U6e8CHL/2ku3P9AXPiSuosE
Nqdn5zcD/xt460YAS5wpWf1MWL+OmCkqAAbka4bq7Tr/TAJSm5h+jt/KNbJgV/Zc
qai+C3H1Ua76m9sMCX9OnRANYVjTDhuUrU/VqLe3b8Kq79NwqA7klUCtnVkF6P49
q7yX2gadjJ9nzVCvPT7ZybMoTyeTSLMT3Awjdo7KOFHknb67jRRZJ/2dUEESvIXy
0qwdlgK0FCkddcpCtP4mdP39eyBymXtQmCoE/Uv/CjtOPsV96CrL+GT4VZBcWJmi
FnxdaB82FORtOHYgFko1HVPRFgG5AJmoX/zVusXMAMye6tNELP+taxq9um/f66GU
RXfIGb51oaQMThj6llzG0kqtPBPiRsD6gYli+IDNEEmXiinp7pSQ5aTuVvcQ9BEI
h53mnNiPpfrQBybcMo/e0vOKBJRfKgo9+oJt4ISRX9IFXFiWqnGGpHMYXKemF8+z
9sNM8pP8IfEGh5U0j6p17RfM5E6I2bkWOfP02SAfwHWdY22R/0Av979+k+MV3BJC
m0LekT8bD7SX/sj7Whlb6OEogAPkL7HpZ1nMo+wNW9anqUpH0S1qcBtX0zzx5fiG
FozkVS+6sL3VcYo6lBWS/c4R/Gbh4h2U2fZ6+AiR8F8Lhsb/ySJ/T03lowoEEa1e
lGMGP9myW/PG0cNVCKU+2vSO98yYd52tQDy9s3D23as/SGh8MO2/iy8L8oRXROfI
M+DYqrcRtgBsUtoE3eEf52hIrjqYXtAfsgsES93m6jZALFMTOQ4ydJ3XOb5UtFgO
vKSC1+mR7gyRB46FOm9GUvWuW9+hmCmzaLNpBiPtcLpDh4m87d8nPDB8CyWmQ5v9
+D7+SRW8WzWWnuU8nwjdq3a6RWp+Tpp+75Wg7SVn7sAHR7gpjlyl2+KVu75FcVJt
HfM4P7Dsi44+xYUv/fFLEGwRk3lrvGnaQ2/26P9p8jrY2dD4mEHp7lfIQ30yyVWU
k2Y2xrZPlMGdS4e7TOZYPKDKnLcdc2uPD9o3tPLS8Fkz+rR/INumQLa/25i7FdN/
YTrykPJG3NBFl7MdJNMo7GxOCXEwE5kc/pBtsZYKL4QyZApU4av0afPuop71qAGy
LAm4GhOmjMKA6uNfVUv1+nlHZvayTIYPeUeHYkMH/mEDUz7QsC2G6o/+RSK2DCXN
rPqGPNpMYNqs1Pgc6+MDFo2S6yF++3DPbNM8Kqspdb0Z8qRRtdYIF8TCW4oIWk/3
2pYQcmPT5pdosKtj8bmk0G3xDaHUpdT85vt6bM7/7/3cRPzoCddOm5bvzUezUtav
L3t2h1E5o8CGWNEF9V7WHSzYDElGMrxmDIhNS/7vGuIAbr36aDM1E3kYpoTp/8cP
etu6jTCNOiR1NmdfxwKGnP04LUg5DMxKzQE5Nb1+AdFrYT4NTmQVMyNojiIDcF1S
rbZHBohgmUWOBYUVUrieuntZUiOSakVDFbIpVkeuCwWbd4Q3/+YzfuXFf6E6J+OI
aCXq8BX0MovJllHHUOYlvNX+MyocHZARk6K/Aw8KUmgEvPTsdDZIOQbf+d+fT8B1
mhr3v8ROh0UqUJlt+FMY67xzSD+qppnFIgwX89QGp5sCtUYUy7SmLziR3M2nsnt5
65FjBdXmgSiY3Dg0GER9ZAbSR/cAPeq2XrdDrRgW7m30xRXJWjeBvOpR3WJSO4MW
n7HVnTgT/8rSTu9vPrieVJo/TwItS0YW6q/jSqs93W6xwoYSHInHRuQw6LW4oxTt
l2Y9oORRo/mnvdxhVgOq0FNIB/Wq37rq07wzNnfB644Z8vsjoGJAdUFTOd82sDDw
XotsruFKWBmFmkCER6kDeNmWZ6x7gpBqq5czCTKSmCKFLqju58OFAnn2Y+CeVjZU
I72zHgSzvVvjPv6+qhwTt3ktmPI8rxCbpq4J0BL0wCi/4IwqjMNKI/Q3okEL2wqQ
TiW2SeD6SKz/qUdW1cKXGU6ot4jk6+hvLC5IpRWO6QB+Ibv8hvnatFOi3LLZzq/e
srUqsmYpx9+IKNLJjEPKjZK1sXdgUe3aKiYKoqXoNwNnijoRDjna24/Wkvu421Ik
UM91OMlGCqh+WrQUPPCLxz+WUrfHvShObDEaQa9ktHL/G9IT/PkF4IXrK40rzNBu
nw3zDJ8GQL8Vc8UMLb0J0MHGCJ9+PiBwaMVeELaJfe6jBJ5t+R/yZBl+EZ9YAXFB
q+3CUm3ouADFoG8PzyoA2t6aQid+r1D+yl/Qbh99b7E1szrnhx14lWgbLoyTEl1C
u2qpLOZtDi1OAXTea0hQ46SqljUOm/UqRqc1YmIel60b1uAJVYrGu6ySYU9XZNdj
xn0+Zl1t6EfigPOmn57Dt2B0A/lWwkZVbt7eJ3qC9pTC2CyxJTtxXsLJ+gD5aTn6
Wkd2XWU525Q0KGK9E8Ri5G+YCi6zSsn6AraIJfFzHR4wvbSH0oj1aEej+EQhSQZH
AGo2PqaGEG/+vTkmlU/FtoghWYwLV1fgu1ipFU6YsHGnN0DBF0BQfdiXRe8N9KlD
ndHl0bW4E+kxIK1hcf966yYvvP+zl9Y136phBFEuFMWHn7XA7BB5C8JcelD5Fcqe
0JDrpACMY4y9n2U0f/XZ3xPQkMFLmtEu6GrYaHtOQqGMrrwpddf7MHiw9e41jjn8
CyEzDXWVuy2R2ZrZCu1HmOI68Lxpbmcbt68glLJJBJCEgbpwVSF1vVp4JLzDpP0h
bxklPldHoBLSxNojBmGSZbkInZ5NYUsbB47Tg+tIhBlKCzepKR+faZ9PRzJMPV8/
rXo355kHx+atGAt+noLsWUEuuW4xvffExbBc1BwjJV382391OJvA2KoTm+K4X8Ws
Po4FAlVAep1/hv7/S/E6ejn3k+wKwxcdGYRt+mPXcdaOW89J2yN9zI0ViyD3L2Ex
uriHEtDVNR7qcTfYY29KGCJ/VjkWXocek0rFg4t6xpi7u/7aeBHPdSa0oZfTAIg5
4ME0oAgs6L1kQqliPKQNy3SuX3XjhtQzeBiPyGNB+dnSpQGKJrtQYqIkRY1aoa7C
eU8zTbXKi5vL7WfE2gQCy2X1j6Rs2pgurxvJRvBiEAhUEofkWvmOpCeGS6LCcQu3
n+wTNhDMTto/j3yPsr4zry+YnUU7sl/lNstdQ8JdBxq8ICGStInzCtNqameAIpN6
KNYgUEY8sP49jyjlKfkRCyR4ws+b3imRBP0Pp2lzb2njArRZDjcWsrzGh+1Z0bio
JhqlLzchI+yzhnuioikmk26AFKpLln1tWnny+9AOsX90kNmsUp8+alKOHMWUoZ5J
s03TusuDI3Kr6jdeDIkbyyU0/rupdJj1oSKxw+hZMIWJzLD8A/s6bumEZIQm2G45
h1zSVIDYZ0EDy3ak/veEt2z2pCwUMvaHdF1gz/Nr6Actey4leQKnZp9+bx7wO2Wt
xWCsR9ENKKQa9nWUMB3tj90cCrSUUg/Tb6ICDDQudjVwbCltbX4BU1ZXYBBV438f
Yrv2Nb+OP12yXVIowVfoyT1g+13+FIbsVZ4cQkVqC2Si08G1C3EQbDxbUqrQVOjd
IKQNrJ6wyl0aZ7cWtsW6TkAKkb4VWr/fQx2G/cW0LB+mDsU/hcswcDSieU8yr4/g
pCDY7RL3dJh7i3lvTug0aD0egGWb+Hea1v2hvu+gjcFlhTY8mtvl9Cr9XCQDhvb5
69xPj9D5sUihsfwPIIc8LxxXM7EIqofcCBrAovxz1Va5TFZckIblLhPAlMUwAmVd
PY5WiINuP+0tWlM335H9D8uERptFy6uJtcnxynW1mADJG2NcUt26GruPTWBll6Z0
n5IOZ3//0sYZpa0Oxn8l5ltTHsZ5i1WmKXkEdcmwUK87da8U6zjTT6jCTHVmAotv
A599ZoSJgCF0Ds50JYOhAWEHLrPNE+nfyc0ToiugPpJ4Z4BDB4f6xUhtah9QyC7d
9V4R3oTeAQe11Neua3ejZTauG3EkZqCOOThlBrftikf26P3HmEYWs4kC/D6SPQD0
Qr9b3XwXBXhJAys837S9gwNZeMthezrIArGzyMwq2LvFmpfMpCdT00oaP8gVEvfj
9Wk1YD13ZIS3z9ckVs42JApSVRM+Ugy/OArbrirWVTcN9m7rNU3uMCFnnZ2sFK8c
rNgwroDcJfbZNbJqRIbuVW4FwJKpQSRt2JeQTdLWOuGuWAEuTATjQzPRu1oaf+wQ
KElF+P3qE2/Z/E3aNVEcRSxx9SZbdNFOswgFpZhoT5broDkUFn3NUc1XN74qh/DQ
fw110gkW05EwZjLh4CoMElVgGZrr2WIHW3xDCCPvFHf/TgrpqZOTPD2VsFNCB3QB
CfkCYCRZ0v+802+ZzttLQaIG4blYbQFNYhR60jtcISaks7KOhQ+gT7+48SPGTDgb
3Ctn1AHGJjwn7otm8Zfv/hiPBSAwpqCB+aYmSjgJ6BQmf3oDYhXTiDvwdg+bwL4j
W+YH1Iky7sxwjtME8BGREsNJ+zqS6v6t+/hO87PzFKeqrmQi0SmWhtLOCidu7FwH
n9IBdv3weRjayhIvRGjPmbo+FQKbkNasWrAkub6GHIHpxaOXUMSzFbv2PM7RzoM1
MBNvXQDzLJj50ZHZFoCSS4OjgyhPI68diKrjleLgaBuE7nqdOOp68BzoMIzKh1bX
Gc6xmFw/4amI8wzbWwYl4ZrA0HUY72SMobRCN675KwuiR54WIobFD4JLHSQp4Ura
HYKEprt30cCA8z7C8rCSDiPC7Vwyn4XZnvElyJo7/FWLV5sRxCBiyrqCY1kOY1+Q
Q2jFkNnjp2Slr7qAjFgBLDwhENsLjehP03PZuzuUpLbQyfvFePxPud3EuWUGadcT
6JxW3nkiBQl9HWY07XojXv+5bhJHfl+mRaaoZGY8b5Lq8C3paSDiZKzl6Mr01XPl
D7Vrc8tyMAlbxXng6vY5gge4zBgRCi0vTR3i5/Mgd4NO0w/0KNQ6HrhrfGhuyL7F
aWJ/ATamXyKeOe1bB5+229+1fS6d6gp4FA/cih6dKVqdIGTOnvihoj9dtTMYJAZh
RfFQBkyR9eEnklYRR2WYs96P6QuLIXUu0qP+mbmBk8XJEZJ/PLWgwojYOFTGt9Eh
dJ5/t2bMsZ7bla1K6lz0j/NAlRrgExxdU1haROUT/HP0Y63QsR+kju+2fb4o/98R
AJiBK7zUrZ2FjlwkxmqCqyUpYL4ijebLBVsxIaDxLh2/271O5pwTJ2FdM6jmBX5G
Ao5+pDf1gnDMpDBAMazEeyOA5v5rEuPGIzX6uBhDWN1bfXH955iClCQ8Cui4tpf4
N6Agvbck/DpPTbv+BmaGzoIpezn4UJ1pbEwLMKzcXcbknCrfAYUDaA1wWZYb1oJC
mdtw1FDGMt5uMXDov3W/Kz5M0A5JxHeD7Vr+jH7qjmTU73G/OrH9CO7VPIHL+9HV
adS9XyjZju4lhg8G4PFDpoC9wp2UAK0z+aYBd16xPP3H+DuNmkV1M9m9U1C85g2g
sorFqUFC9Sk878uVOOjCqP8aHNeVUtTjdmQ2P23ko2+8sUkUZ0bquWJHpqEw5PHj
caqgsTEpMzgHLp+29cd5fg+AX2pvSY2WG1Ajvr3za1atYV2xvyIJIEOmkrzVy/5A
F+hXlMhnSJF/tdyoHtiV+pVr6NEG28AtQjGL0piLNwOPTDMAdLCT8GgTHU6ZOPAk
HkdJ7Ngwd/rv+PvhTCrq1smGctwOrifqQ9M96aDLWYQ1MO2mKbnHSpow7HsROWH9
OVtzYnfHTCifqBAMrrClkTsFt2FFZ0Owksz0P2ZLkFWuqF2wOSfFJSs61xf35qUK
g0NpubfNgWiyuZO9YBTU1oFY4O/C/UDGtJHhhX4q83fkRkU2aBKTe3+g7czGRb64
x7nFVvpsm/WyU/V4r/vKaHgFzlDO8SIeei+WmV3uf2EmP5iwWZePMWJLsJZM7qA3
3auSsJFpLU6CTxSjxmvFWT4GBcPuJsIpxJWDjRAk6S+fToE8Fpr1AKVcI4frQabs
SECaYwj6J8ivhM1JXID+OQhHMZtPVRm20AIbuyoIpgWEJN7gPTSgnybNxqbMua/d
CmlPJADJI1OW+tMcvneCQYVR8bNTzOfY18XC937YwPtPBLSQXF9JWrHhz+2Txxce
V4QlRAVFqkXiBve3WqkF0aru4Wrr0QPD7o0ONFxYUVFYe2xm6/r3+2J5fdx4enPw
Xune25T6ZfW9iZAsWY4gTbKwX+YXGPNkp2c4E9s95FIjQzrtx9vCZAgaHJKRJj4a
azKImuHC+XJIzXfsf1pf7gay1OBfS9G3Per5LGZHFcDO/G+KzQ1naVip7H7CEkEU
WX/6wqeQ/17q75lllNe7ySZv8FDtGNgsW8TR/zsPORueqvqCalgPW1t8a0Msewrv
JSvICX6Y2hZPuHKKETKP7pC26ujRCZpt1LK45U3i/re1ODsSyYezjCKlbSPkWV3i
NbGq774nOmSl+Xr7puvfcEc8XT1zxpFpHIhIsjzmYp9thaVOp3YC0prsu7O05jAO
o8KVS5C1Xdr8MyQo6uGWWul1cnUToN/KlV757AISYURd1YirsMruqrcyJHfWmbh/
cfP1SlT/hqxE7jl070GE5Z9eT+kRMr3x5sQ6yEEIW30gb9Aa3KxVlc01dlHZ74jX
bG3FPFVRRtZt5Kdn2l2z4tzk5qU6X9WGeeFRTBgh3B4UbXBASYCHki0wNkhBTIsl
8oggE17rsaklwAbG8sFSTn0lJVJnOP71Ph4imatHKniLQxBlgQOckZLjMiPiFvaV
g2stYiXHSNEOyaWlIo3BVon0Ag3ZYubBMoyEQeoc3VOI4nSqZtubmLZn4qDE62Vl
sbSSYvXu90Nr569rHVvD04FXTz1ksfdoH01LeecJy2BBS9BlfNZEkuHWb6tD+Z9R
Ynmq701V1e9lDU9OuJcxVbTmWSbMPnyVGdH7n2NTsSdISnzG1LWc75ZCfeE9jgPz
9FDGhh7YhijEPkRp2lioRC3cT6zBTvigs3e1c67mC6KcfH4f5nbO0xdD5OdTCvC7
/9Q/ZZPxTf0l2J/A4zy06dJJ1D33LLFZ0qQGOOcnXGXdnguEc2knAD4Im8LXdi0V
sBNRybFfqeroIlhaPDvImge+n3MYrb5l0uuurcRThH+arG1xnhUC02Z3ROtV9a01
//RQCzPjKquNDDnPF1X+jSLOIig6UeXIHdWNx3GBunSj6NdovYnEirhpgoimR0ZG
fY08+wc3oRQUHVcrMh3u3z5Fd/Dl87u28kv/w5Ch+6pSUewQvLL6kj0CJeZjrKSE
zJmiV5vzOWPmz5xr5THxLpWQJPdccRVMLqGwpIL+gCnYrqBCYPfS2NXsdzEJ/yPE
zs6EiqhZZOslJ1qPBPb4URVAb26JEAdq7eEcpBWOfpkc9JuDK6OqyfBqnp3yvYL3
oB6zsSAMfuhNruamiKynU9fMyF3tSY+vG5CyvgiG2FrlNkLFwqMyzVebrILvi54j
iKwCS5/WDdIv6W3DlwDvHvijhomF4TMoBjR8QkCsJDABrYFu9AcIfrOj0BLLBww1
0rkC4Dl4SHoY8Bl0wK6AB6NWKhWVOpWqS0sGZ6j0fTuCHcjfjNNWyF2tj2R/SIk6
FZOYOS6V2IyR4MV5qki70trnvS7vKYS+oY2yTjWwuYSmomddyixWDgKu1qvajOYv
+uYqvGkXabWywN9WLIUQ0vpshFyP5oAFzRQH/dsS2CQQ6M69KjsejEfIPftBXVrd
TWI1yXsU9R5oarFGWOMiIRnB32NSJT9viFBeritas5762sCfOq5icVJZeRmVrJ46
9yjso9Itl5+a9v7LvZDhX1gayGOLsfvS7Rj9hlbP7psIfGMxg6sPQmTud4lfNSLq
9o87dZVwnEZx/u9oNBcFLcizxvT5QmBpPxqKU7av1sWh25GnCAjoJBOfH4WfJ8Tx
gRPu0ZL3x6C7cEsbCtihSf7Elk3gjgKEnxsyezg8fH4kBYHIpgNvnmSUJYUDXod/
/2cft3ttthNfdw4h1uhSOUWl6rsqDCcSnCcnxApQq1Mdr5Vooi3pGjV2aujLeLbD
q8Pt9v+w+k7e+VmJBd9Q9NUDMmgWJTShgml4rNW2HUaLILKSHIDgwnPKHvwmYPKi
r62o+octMpzvDmxd2wyUSSBX51RbPzoPwL/4qcN6v1vjRLe372a7pxktd7kf1EH0
9nAaDqm7CxCNJJ+XT3NeIq/t9RF9ym91pSCfQUqYBeNbStPCEqUlo57o7uV2WpeJ
VFJ0oFj6akSHo+BCUTXh8cbDKobuN/pK0yTeuFHJUybuywra7VZo82Jke1WS7BhA
LkQb5bcE572eQfDp8sS0hIhThZvm5cC687wLT1zFVVHcJ1dLsb9ICJsRsIfdT8ED
o7LxnzoWNsok7sg6j8UygH8JfO2zevbyMIWheUc3W7xsqqMqiq5G/9NsDx7MDFGm
YVk4QIn/suSY2YENyPtiaCKHjlKZ6W6eEVWWgBNDWExV90ZiNl6PJdZbnHGW5fKO
fxMGk+UwC7Ne7YoZBfAGzEnxmrZoQej0GPaeKaxgIvnTJCudfs1QDzpUzKBBPgnl
foqP0sUFKmWMN1eLcYQJlCZGoDT0xcmYFJd8iO5s/j35WQzd241NUmuHN/WdfkAx
Dc6Tzwy8HxgnUQLFcstWdvyfJ/suhMBIPcEpRTqDf1PTaWfwxWoGPeKCVo89ET+P
3rTupyFCxLItKXsf8gb9jyEsTahbIEx+LsV8B3ccrCKzlXuYAfSjtvnmmkJqjj42
>>>>>>> main
`protect end_protected