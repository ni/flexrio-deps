`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14608 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMWORzZC7bo0toZS2Zods6Xs
yljw+BvqICQb54hGe2JGpCy7VfzPucQWBxxbAs+GRagpFs1mQIXQJAETVK7KfNeu
KbQm0EDQym1xoaPGtmcykdNyv83pLX5ika3wrlOz7cr099PwPVTVqJ+NKQAhOPsG
72trRw1ZU2WI4ANQoAFAJ9X753YR9lhsbN+67jjbomO5qshe8K9+y/qHRcD9fgNQ
qedMrtyANbAZqViQwFBLUjHu3KuWDkPSP+x/68+WMwJgPWWNLFSTtt3xo1YyKqny
Bb6zZK/l2ax80/yzV/nbOH1oAI9f/88wXEaDtIH4FWrrzyKSYDbdoKgFB6bsqNwh
XOGOUBDtb9mXNQ/SPSOly/FQAS6N2LDBOozs+AZB1EcLfNTOYoNQpSoCxWRA2Bbo
Cvt8lgsg9UnPMNj/e1z46Y6FsoSxVnZP0djhQKqAk2zIF/PAnKdA9HK+IFN6xaX6
O/uxbC6WUfbMZh7qNRzbv87OWqr8iVK8cXWM/XWRI/vJZwm16OPDVvTMJWGXLY/+
PnozlFUyYiIX/pbD6RZs+rJe5bRSNCmhFE5Ry4i4FagAtw3CALJHSSuAEdKUZSaT
0sY/fqt/cWLCS3xUrXQ6BikkyW5ictJZCZZF9kl7+nDje4DVUHK91fx1IRPCyc+R
yZPwqOT77/agOJf79MPVc7fyqUbCWha5rn7NDi9z/zXJCV00WL/OSYri2lMVpdBi
Zbh2KWrfo4ez8weq1TiyZJ3dxdNRShTnimQj2ZuR91Gnm2195dW0wRuw+NmkJwCB
CaMAQs2rD40J9LSsFhbbUXUYQ+8tER9/Sip5O92Pn7zBGkoZ8AHenPEmP5w3t6tA
SAhUDeuoeLiEOcxPCf3XM8e0+x1nqJGzhpx7OYmq4bUon8UxbfzixLxNLPnG3CJ2
X8Uix87q/YqG7DGty62VxH+ajaOEh6ZXMEOodCHT0dLTpFjwt2mlcWwWJFiT73jq
GwqexCLxdKaz2e3peKAnrB7RRHMt0buyC11UnpSBmF54d9aXwjI+B7WHk5Vvn4u9
Qld5JwjMvUkZOdKL2dT/iWLlCcYrBLxtdp71SAiVkGpYwMuZL8dm25bZwrUq63t2
iohwbeXdgs/TCLhLdF2+TsxTQWLCbBZq6VT7OQCjJZ28UGV71rlM8JK84yOXdmS5
3jWcf43YrvCmcD6ttfD5pJ3d1rQZYbc0yr5YKi/fC15g8dWasf8qwT1gLsBWClps
UE3ujpJXnfbsFtnBxbwfbWfditcCQaeZbumdMxtrjoh2mTrAcLNiWt7qmuqYLLdc
c89P0XXfBZgeVnXtj+f9kjDTcO0b0n5damh4n12eCUN3PrMDz9WjQIxd409gfJvK
8INWD5iu36gxzZmmcU4NGSEnjZOXd/QK09sMOYfgiqb4Fr5E7FsRdo0amYXCPMhF
oPwmioNYgLl0V8dMWrWpYlYP8wRf7KLu7XXhzVyMJKuPXrFALhSoiO3gjvBlB4DC
1odXiPFxYJL7XOsP4/47Yt6LI3fRrXC1MjYUrYDBZ5JlwCCZS1zB+KN0LP0U5qPT
lt7AyrcPBYvhunIgQXz+fPeGDiEMV2mMmw2mfsBLiUSieh55KkM4rIVQy2R9/GSM
EOrjLhqP9L+B2XwNO5kxguOcIXxpjzTMWQqIdcNL6LAsJjZxcoHN7GFjEUZU6YLh
EPn95RNuWdMQhpyrp3hMXJSNrELVNDqPeL6Xx++XIHDuU4bCbsZq2WnACEEsGmSY
vtZn6BIh3xlVNGc90QPku3JvAJWr+RsLSMdPEpXfBQLayyW/j3mgK3sDCRC9ttRk
yuxnJlYXPl4h+u36gVFFK9VUMOjUnRe8MLnEGs631cGuowSHy/jaGdD2oGJM7N8v
O7Q1VTIX8aNpmsmx/K74l+ZUBiJH0tKdtztTR8o/P4/24v3Rg+5VsBnT1Yuhw+ma
pD/rxtxHcJ80rPf9Ft86q8lWcGiwsPaBO4zaQAfLA9vQGzJRUCzK5KV6UgYmiXl7
D590c42Mi8w4dEsEW50CzlrgpM9d1vgkzdSLk190w1X0GDGCrORJ7uqgrSXAF8yv
BZ86zajZkuYsTr/UZ7idS691z5tgpF/OIBOLxhugrT6ZXodPjm+FSzTupcbaRu/3
vkb0Yqpi8LTEFAalSV1/u+fo6DWyUaNbuocFsc7tu7QuIXTEVSdlZ6vkItr0yjP9
ioiqF6rtjMOhxUbKL66hSm3PfIVdi4UzNa7nl/qZkucxT0sIUtQBsEv3tVP+N0KP
vfxwXyatA16BgXGs1iax/MuhlxjJstLWSqG1BLBf/hoyyCWFnIsMwy6ZCbOF0nGc
gaXwKMQsGtdGLe6luKgPtkb0s1OKDeKRAJtsalJ3ZJ9hGYJizA3kvmpnlNd0ShG2
jydZK9xY8FSQnXu2ZWuTn1DJ5nluJLYmJn4uIa5E+K6XF100+sdfqRblzosDi5FG
4N8y0QYh1+t8HXgYpDwD8OduQDrmawit96G9defFfQi0Zrh7r+Gh8qq2qbop0+l8
UJvSCxUxzuAKhc+yMx73ZlKcFqp65lL2mhT2/8pOcKtV98P5UMAFv2HR67xAH+nE
bDiwGTBYXD3xGaLlY7yLL8PejNRBtbH2swWkIrhfXKrJnYMRIBAlYJWV9952f6pS
AKaSVdw6vkjHLQr4kEV9QEWLZHIJ/rw8eKkSCSgnGtWxVV6E1fY1KAKXeUZeNKxT
IvnGBV8aIWoZSzG4FqODrSYvYFw75ImFt65twNnOVLyvdQ6XPJgJ+wI6hgLUmun9
lq2OIQl08VQLbdSUjPLY9CDz8Y5/Vp94w53z0TSNIbadtAHG8Mi6FPTe63Zb753+
GV7IvGWRtjF1rzx4+ViXjdF2X9rcBUivfz4CbV/wdBHz8TScezJsrXk3nTRebJ8F
dedPGJeh929lvdAPJR5NvkT8Xx/gAZIYwA9grJKCSvUYm7ktjPZQYmWYp739uEyf
+Jmes/kHg3eN/oRExmwzrnFu4HQX56cUWJoZe2wwDZNu2zpwNDDV7+KFoN0dAs+u
gLNRe166HkiPEH3Olu8CyH4dF0AArIRjZwJP/+8O1S4NrhiIogSiA9ZpaAVhE7ll
VYdHC8BddhMOJPIQcq8TD7po3JYCn9llYcmKa4WXRGINu3xDffy2/pTwtTkfaN7c
0TSvSKb+YjeomvWBM94vTOJENj2ehl6OB0RtK7JNuF66z3NoVXfiKUzjmyeSRpDB
fJWFrxOwB25N1RxOhQdgG6sQ+ty7arWYbIy1cwokGlrFDWrQzi1rLA+Mypb98Snv
C1xSkIXvi3OuTGjLjNw1wUtVQ009zV2t5M1sgijPky0za+rvTf3RDRQlvkZA9qSO
UJ6qeltNjYwFwMFqkvQM5W1jdVoGhIAcniLZ2vAQ0TrJb5cmiIeq4XpG2gbyasPW
E+F6409s9+Jv9oTM0RGvc5jAmG6GuOA+TWJblV8mnpP2Fv5mBOdSe8V3xm8Q0AXG
ScqNQ/stb2bzgbwJ26vWFdUyRAvltunA8AaX7M3IFx3grWMyqa1k4tOH5hiZvaRu
C6p97X0dp/9i4gRkNkkRUL6RfOAgBfy3/JkBTnuDKEvLqIaHLI9qkwPpZWpHBgwr
uj1lB3uMebW6Bj/3NCoWlx9FuUIitU1MmE2PYrZIPoIkCCEprbpMgPKFF+Jgw8iz
cqqdR8sai5dB6CqhZf5ZcH0u+3dMlKIygj7tWo9bqtfpE4F8QvugMUG2N2UUs7OS
IK9ER24rTG72QxXHP+ePzy1GEAoixjIO1lQfSjxDDHDPy/F8wlqZ2ChgSDO5bbNL
iqVWJtNpWDAJoIiOEPDGG4SurMx911ldQg/Fg8opV6Kk26PNPLdaO3EAYcY1QgUl
qVKkL6LPLI9ir014EdnFqYYjL+4sKMA5psebtJ8VE9sRO/pg5SZ/7tczjfvoz1NY
79K0qGKBqdBvDQtT1DdoraP+tu10PgEWRYU8Av3icJOiA/Je8pzQesjcjWljcICk
F/c776WPhh7Ksvyt7yHRzmAiHYtAl2qkP/qD5auZbJ5n8/ciZ9lYWQ0WKC+5AUzg
XRr7ZcaOuQMU22SvpXWs3JIergzf3kJ5upq/qP5zGsC0Jrvt3Tkcu2avzk4Aq4Ta
byHFrLtp2+TG9h6g+I5bpKOhEOpmIQOhJokZ7/jDtgW9ABlMTHIJOYL3zkUd56Y7
dh7BdFMp1MY+LXBMskypDlD9QF9FcJjE6wrsVUXfuE6xPHQe+XohlKfy4nwNngkI
wehHfOrc59gq1ZLJwokjocFXgNw1z3XvxO+oDIZhV25YwqhOPLDTBCvn6sdFSsSK
k6uKIvdXS4wERxKLze4VHyj/KfXdvSMVZOUyRcL/qpT+ZcWpxLpf/cYSaXPUbkQE
NqQ7Vp3DLMIhqjseGbJBzkU2JWFkq6nD7V0fp1QkRK3yXvz0LDMAZhQCPD9oupdi
8oWQZcvMlJDN79Qi8GsrvLyqigJXWk2UWbHf5LBJEkLVRwDF7R3qhYXZFybSDVBa
th0QHBkvBAYwQJzfcVGXSo0cNHGvrfTsm39CQL/CKllmSnXwDEUccyPGB8xB0+pX
bZikBFizMXuGNUOSP1aUAKQskT03+h3rxUSDzWeyqkZ/Mmhn+xNTZA+p2xsHkkIP
7rO4x/Y3uAvraB6j7+gCNL6MSK5Q14Neil8dCcJbFZRvYfGjRl725qjphUXxUoAE
koySYCPp0rwMd3jAuXTfklJQi0sdjwtUm/ZrInDivvZNcU4Aey0q7KXF4Gj34UT3
rxK1tfdxULhwUnTC/6/ALN73e0sJKUoNsTyoLWXROX8TXZK+QJwGIe6tX0yc/3os
VNyY5PfZjTDZiBTunXWl9scHVHeTnHH85siiDuNN8l07np4B+UJs8opJm08US5+8
xyMEFbVWS9Z5QIENViBb4i8P61flTELeexiseSE2dAIfRr2c3PYig9SvEB2eeEkv
HDTu61cDdMKWrXqJfMXO5mJJzojA5w/s2d7dtD1HTj3g8Z8Cltf1kg2m8eJQoedI
4jxg3D+GMsuHf1NApQcGMVa9DdDcnFllyj2u6bwaadrnHvz6+zK7qreRtC3hkBna
L6LH+BzYdgNnCltcD8Q5w8flO8m+tl/DY6yk60BrHc0ulFP4kXN5ET9a5pHjmXCI
4J6ARO+Mg4y8/ysd21Fy+7cXFpuKLkVKbouun1o6oBT1XrCxqf4Zx048w7d/cnEa
2es+SKlHpwpmMH+rrg0tV7EgCq5bX7L9B4NnCxBMb6C2ZD56Ibt+X31IZ8yWr9mU
36T8Zp/H4SEIJhYYbMEbyEaBSOArjT/kNYFDGjUMZNZEUzka0kKnMyTWiQW7VCk9
Wk0pjCljSQ1lzPCasojqMCjotei4PcMsliWPRn1kVyYWdMvkmOEiydpdvnGFV1tT
Q4uAw53CETZJG1DzRWQW/QS0FLsifcvR3JXPGJyCy2z8ZOSb68nMJ4bkUq+dSu30
YuLhngxpLX4yVWEcmARQBs/+g0n8Nxr+MYCg2AlFnwVkPCEMVpO9qFuDK2kR8Sen
fYYRXrrC+6x2SNIIQ2bS+04PaMbvWzEc8voXqee5vZDQf3paC4OSg07+p6d/x5DC
32zHaZYlTgJqg8H2ZvGiZy+Wg1W2ZMVbohsexrkixH716yVcRWn8+W7c3vGih9gg
BqqAl5NBEOMU8sSd6xOSMQcttKYAgOe4vjwhjwSHL4vS+xR3PMPx4r6zKy5Nl6PO
zXTCVopWZjHRVXfsz2lwGYTc0AJKAn6ohn+/AYn4fHTxnI5e+WfIN1Q03zJXedTw
aXy4QPeRT3Owdigox1nrfLTauE3UhOjsPg92858+IP5hh4n4VrLHbU5RaKgX+zIA
6Qlk0bE1aGxGcV/DOGFIoLp1uyF5jl6vTXhy8qBMjTSp9bIUW0jtXVeiP7VmqRcr
RgCatQH1WsseAV3jvWMXodazdVcjWxWf8B7aVST0720k1jhqFK7eebuwllvzOzv0
1tJq13z4DTtRa7b3SQkuuyAMztvE2HN7igGZpbJFs9BqXPmokXvVQ/wX7UKyz0LI
dfptzi4cknRIgsATsPqPLKk9avwEQPBoww4gzltSXT/cGxNpXxFhWNs5ch0BNDlI
veSRsMMxTjv2bGSC14P/iYBUwzG8rxzX9Mq6mW1HhL9ogjuGsrEfU/Kx1LvXi0oA
4IBn7LjIZT6HBzjqqvl9oiMLnhjoVCdARn17HzS9EUxZ/Py4Lb3P2yTRqjZnc/fm
YdQkKi7zNAQwuYbWtxzbQXrUExLk+B8xp6VwaodoJxpuNtEUEX0zCw1MlfgSXuZh
x3vT2YhHlLbXOAaoMo+dmMzOVe0IBfctcwPaPdJ8S9aCSAd8rMwCz0U3DgyNhz9p
j9nC9juJfSEmt73sIiyB6ZlsBQd7qqJaePp7focoV8brEYHNaEjNEfooK20WvFqc
93kVjciAhJpwAYQpI/5aVT1jKia3Y8fXtgSN+kz6RqhxRxaWaPXJiNNZGE6fotUc
Kd46tiC2/FFBgoakwjj3aXvrGwJaFMa3GRCNN7vXZZS2K0w+CRzNwpcCQP4BlhVl
+yzMJGlG+4qECISYDI4OJ400CD2OZ5uDD3mOuSBRT5Zk3QSBLDecg4EnFdnvs0pU
C30LDkFzj45nYatZWJY4sSbJsPBJIGPxRf+xaKexo0OwZhJqhy2IuXc1ady1+Lwn
j5bv3v/tHWNpYd1CCs2u/sqeKSzo94jvSdticumKQSPHR6x5xHLNwncmpW0ky2KX
CKfbyhoPfddbsTxpFLDabX5mzFVhLpinu/rr+vVmOJ7G/xUrCuMspkRkFvxnI/7n
u/WVPhiKHSIPe8yL9cZ7ufbRSokac6smlqkTF8vvV83Ys8my7OBJpZB6AufrQ/o4
BMY1R8UnIadMnd1ZSEXPipXdbwx1SZZZTZNH0TV62mIlP3XL9AmgutzPC9OTO/p+
RFIOA2c0cyVyx5Flsxi/t53/4y5gHsdKBuRW56IHJMG8S2wRbw32DxMUH6ZBzr1w
nhctvagE4UM7zFp5lE7G60Bn5YOPwM+qiBFKmJFRhJUI7JasVErqZE6W7G1YyYQK
NgDnSkf2eyvoN63bGSvjebcbhc4Q4NLFb8HCBiw61u/kINdPVhKr6+L8HpG0LUwd
3hF/n5aGUg8xtI4acSI5Y4WUsSS4B9Qm1HxPrXZgtE6DBNcTRBpdanfSKY6e7Ace
lBmYRmQMqKc4+SAUpjmM5SEaNYB0WE1NDe+o7Jpm0xATStFHLj7/hvgMh9GWOtgz
eyRxiXUAy9lH0G28LPCuD3u3BRdtguVVGLvIaBo+DQSbq0uM6LFSErZnhtWGb2r1
BQaiFITic8GzpiwWFmbWVusMslkHfEJ7nHIEO0xmAI+SdVtamACVTlT+9Sd6qcKA
DHp5NIA/LirkCiQe1uBim0GnhIV5rnPuDwt/VRZFLrO9Xk2ntYX2uQc0Vc9OfEqF
Y/4v6U5XXRPo0nPnGJcYeoJW1RqF6ZOqhDa2k2ZdFq9LILK4EVuGEH6z2fUlmy3w
r5fmPagIDFkv1r46B5A+Q2XyesDhMKFpMJKP/QIzcRjm7AXhHH4fDphJA5pNdDJP
Boq47qrPDTZCtie+oDftPZ7x3NE8OL1RtdLdXiQG4lQkl/Z1fShExY8Uj4544qWQ
SIJRfUCDr6XMzm76OfGDiwOi8J/jrtcGzYFbDNXHbUe9Blk8CqDjQKlj/yDnz+1V
zufYImGEAJsQGklTKQBNAxFi/S+fWehRjYNruABhSi6sU0dMMcqJGObca5Yhq+yh
fzkLPpI+YIUK9YNTzW8MzeMgDYx/WibV7NoC7Ten/HvtlBEERUHor8wrrEJRVhe8
oblSEw68W8xs6VvdIwNf4acqcDeT73g0mvVhvQRctQtjl2NOMR+K791EODNb8Fhq
fSfkXSuDSVJbyRvMXNLUIr04lAsil5K0qI5sFNPdta6ALntHbhVzusAubY+Hd2km
pW2IPA89rWoMW0+tw1wE8pa7jTrwTWMeofi0d91+69IIFI5JfOPBAW/FBOTxSrE+
CIK1+0DqhoZqhCVCaQzK0dxLUDfdXYsnNs6b7JHmRni51Iy/QTt6hFh1gmFiJ39a
IErsgKmRgJ/PWF4AF61kHA+vxnfdZ6sVAo1gfLcQS2mlCCL7Ep35SjktA5ERUgLz
YhPRbZt0g/J6z/f5IDMg5h/5mKjJnW+jldL9cSzU39j3TGdOnt+iJMpdPcKfTaSP
2AIJmRdEOCUvawf78ovSBRKQoGGAQklCtujmQrXeJCHQkeReJAg5E1eXfa1t6wI3
smdcQQpU6tf3jC9aOsh/dqmLf0xPm+hRSZulg0fyH87fna2NuUY0zoXU8pnGZ6al
6iKQX5akdhGC8YGDCSUmxOX6b1bmjphX8ZQ+BsaHgrFrTHarHD5fblL8GA5QTFFh
im1/rclTjS1sSwz9VJRoh7XSl7q/oM92J4Xfrj+BWtfvoUGt+h/ha4KuKcScKJCH
PEnZZ7k8+Y7gLBjdj2aP3lWtVFalGtSOSBQl9PkMDAIMtF4KxIcTThaS4/CjDxI1
KgnOM5dxqKvnYvzKuyvsXu7orAxdbLnOG5Db68RD8qtKFa90hBrpOc0016a9pt+n
eT9NNoNceRGcz7rh9lOOY1m8FeTcSqcl67ikQobglZ7udmHsKeSW2YsNT5earczT
+wDxsr+4xXsXQmPHeCz6AjZEUQAomN6lBRVxYDB0Yx/LW2CNdHUe69nrveYgEjI7
2TQQpqZ5TYsobIWQLVT98bCo7cvff1SaavHX77nyW54CowxYB3vQPlHMMZdBqjia
dLEDzuwcpC5oUT+tPlecxTpO61z6IDCebyHhF5FVLHCqGWlYgmFRb0su8akjxhx9
fqnWEjWo9GQ8JMDu540GydDZQobuLQN8rNVRhHQRFJBlHZPoHR+KjgXFjxpCo6TF
GGE9lzlOErSUWTXJZlQ1GRmXRL8D218KeUfDPivVs2qTruTTax1Ixjt9WoLKdldL
0OfuUo7jtEWphoMx8N5bDRAk9OrWX1EbXGnQgIpLGIgDIoYGaby1stTiRoH/U44c
u0vzDvFoM70lB6CTb677k7bXTXvak9i57ZviXwq+gtbtuU+PyQoMLD8UXYB8fS9z
4zkSe1LxMjA6orAXoshT2b+fNikTFBWcG8pP/8hAi8Pq76Snl8E7b48BrhOkMvuv
p9HhIoiSGtQTaFnhCYT5yCLMWwdP9WJWNW1S8FLVMIZeAPu95rJjdAZ2u8i061ln
aZHsn6w+izBpb3xIFOXXU3DdpVOOVgIsqExyvO6cD4jbuhg1BUKTChURmuv9yrY5
9T1agNwoCr/yxxYTJKR5MPCiSZXu/Oi7p38/A4wzg7wtcqb26p3YT2gUK+tzhgzI
rOndiPTkIb42NeSMyAyQBYG/dySgslhDiXCzsy8ekjO837mXJe2NYejdQwgxjghA
ScPlqHFzbXLqhk625B5WzWbqYC55Nu6f3inuFYqNOQx0UW5vC3qGOygbjFWVYClN
12jZHod/yqN4msiQdFHcllCV65x8wZTLMgyH7tionxI3DkOmUAq1T0YKmZMg7+1V
N2Wx0WN8ST4Mt/rA7GLGLUaKLbvEzIMIjjp6lVlW1uwzUNDP+ilJAvDuMQP+nMtu
jWwafofeyM/EqIr5oUMtmueSwmSQz8PnMKI07YJEmUtM+2sS7KeB4u/8EPPbW0QH
iWTr0XlE6K1xRcRXovqkpFMHpfXu6QY5yNyUMAF5RUsDywAGJm2TKdZhDw7Ddyas
NzB5MxhQPP4IUkLavmUsZEK7mFvBxsmyoiDW9lmfwq6RoPuRNCWZ/ALSK+FXiZGr
ohRqcn4lah6qCwCAlW2jsZayYLqb+3cskiGZmiomo+oxirKiOZxCL35azvIuYbZ9
9BZEo8JBkMTFOibH+3+CsShdydGv1j8P8K8AVbD6NY9fVvthSQoAj6x663kD3yVo
Xxzx3m6z/MqhSrah0AFpyeUwyN1WZ0ftREWHkgMZVbUczeYXg4QA0bRQWv1x08d3
DegHnBQLtinSsfjsiZTk3QGyc5JEporPW5Tvu258pVjgseuT94qfU3G3rIaqWqMs
P/2y1AD/RIC1ndmGcvCmeHFG1lzWk84Z8U1T3B2RzYNkkQ5F8MQ47Y26SM8QGYaP
MuVpUIV8++zz6OFpwvxPCE1DaOvUl0hQBtqHf86ksJfZVIw8f2QgFwBjw1/7Rsee
fRsVSVsWJoUIl/WYtqmJJ5OBcieruWrmBiN4Ej5UNAg1A76W3XhL4CaQhrD5JUTl
0q+g9PFsMylVpz/ubIglKCXVCTKtFnCvbDIKtFWUhf2Kd+K0uToy2stL/lnIh/F+
qjnjlD6xQidgfAw73RuAQ9uk2f+t8E5IXzKk+yv/SnQFNxwGubwGBFEB1Uap3gvs
YQLPhP9bLkxnr507lWRwR+cjDgqNhWdCarfbnVl50AhDhxtQN+AHp6mwTqq/ba8l
R/nEDXRPRHOMwpBMhV0bqf3B4u9+ocrwNSnnEIH4EJg5+xISqRoXFe+tfvf1Jvo9
sYXWU8QjvK7MemPLlBwT/X83kVkLk+xX/cgYeRs6tYP64Q9pbA5F6lBaWNQ/yYZp
oc/qdqUyYWpplt0m3uNFybM2D40Q8p2kw6FUvhtXTOUHs46t0zWS/ck99oYFhiDF
mKcXetonHRAH1ZokGLlDunIHBNvh3vwdsuckdWu+PDFJSW8K9hCgsVJ3F5D0X28j
Pu0ugvfqce7OiZsi/52XQ2gNuzDEjEmOGy2pnNAdoz1jLx7jgK+tyaDHxQvjulsl
158T1MQ+CsISiRnCVQXaqyIz0uVCFrTz810OGb8ybTy5dVwtPzF3w8j5/JEbqH+D
Dvy6eH8zjoKyOzsh5n6QbzLlAUn3j4ZfqrjYVj6G4tEQmWiJB4gZltbpNe1vMFLr
UORuQoRoo8AsoX9vVi6JwCGtYiv3XWjcVAQFuQcuFXrhZMpm4qM2JIJ0ZzoQKDje
NV5akYeX90y0v/JvYdyb7+8RtFMdJrSDx+1n+1CcI680plSjPUpSX39NRr8ECchO
Y/AXRV1SdQFrIX0hH7iPccNVNnK/zGkmO9MlL3ZyQib/OKcDsgJyE7EG3+my1711
1y4myotLoCmuw6+wnYmmb0WfvzxKQfG/8I6HkszhMYeH8Wl2YOpFRa6j8oNUWH/b
n42FCbx69lk8q7jPAd21ZRT37d6g0ZGSl997MvobRpH2xc3+orGzaJWjB0z5rP3n
19QlWQ0WySpMxkc6U9QgTjmIUEmg5kCY/lNLmqGIbBrrvS8pWZNtzPkPSycatRHW
B38WJ6Ih8DalFZATqiaFAHysyS4I1grLXHC/j3MUKRJmWlf5sfrpTlRDBSF9hW62
FEGibavezmLZXIDkDTxGa7uBQzULm9CsYl6oC86c9MQ/EAf+URvk0L4xujmS3JNM
A2qM5n2pOB/s7JR586CA1Z4GdXmVgqMBQZl79k78Tvm1koRmHETvIESVlHmyxV86
2itNybkihKu9yJmrCUZJEGHvQaBU7xXOM1KDdwHs+I+EMRjrDWi2TegwW+ACrqU9
37HaWlSJAx0/WtNcG8hToiyK4zp9egwq/Ydw0HRsec4L2a7BF1Ge87Z1KrTz2wV/
MM/J/J9085A9IXoRfWk9vBtrSc6mIUd9Iz+yK9RherpktWJslf/pOwDeBmAi71L+
s+k18gqbsDhiJYRcUw9KMnJhBD5lEvYD7hPSLp5qVxT075tD12EAhkIu2lvV4cbA
MJZGoo4IU1WdqbQCJE8QyV3Iq9AmURN8JkbmDJZzhIgGCebGk8c44PUAllSf32ld
C0RPDDrnytaP0ffDG0hPMPVZ1jXvRlw+3JfRpA0zm3zmLLab3S4MENgyvw7P55I3
j6PnESb87JNLyuDgQx4MHPMW8GJQeDAR1vr141FnZ+CmYmlvYiPwE3L0rxMqmbqG
bVuMRK5BlIZCN1ZXvB8qvC0tx94ZiXu4g8OyvQ0AV3ZZCeFwlZhdlQH3videCW80
SLINGVkr/bNpabAgsmfQCvg4N8JAjnzHjxTw0sVgXDnn4w09gJhEZAPw8yCTaQFk
voi9d2y6+0MtFMZwcc2rjPzRjRJf6+S2kTWG4NOyB962wcVSYP/cuqravF8McNWd
NHb5rdmcQeMA74fbjAx+yqgRqSZyQbZowV4a5Q+XcEjNA/HNuQ2El0Yef8LtPoc4
sOSUIrnCFe/xjWvsHN2nSZ3dsB/8yoYJG/gvaDynduz1w/DzRPBh6VgOAlssFME3
Ma29e4S/5EHXrquL1mhu2U0UCwKjQWB6LZPh0u7tE4ohowStUbEU84WFB4IspRhz
tDx73Pt4Ai3bBY4a2n3WUfmgdopOtiO/PuIeR7fDwNJ//N6EatcV/0f/Z/uXNUim
Ow3YjMBHjUxH3v2snuHHxgLBuzDo0IAeqccstbMKCAawj0shDDrhQc8RkF4/HH+7
6LRpQWBv5nDsmq3cULSi2GXq7DYORIDsesRjVBvzwDzkB4czZ9dbpRDE059rxbdh
pecqLYh2kW0mHgPl3381K2vUmszVv8Mi6fIu+zwJ2ciTmC5nw3RpR3CiKual1VRY
sUoMPgH4uuitJ21xCHg+mtOjIQnzyIHGLu9cSlN14HoWbDXihpCVtbiaIk3Xu9n6
N1i13pVBYcisksdBgHY8x+1UMIIzLHaH0E8O+RnHc40kMlFDumhQFpIZv8rixOPN
KEpzoAk3MH1I9yqI8cNvd1wDWEkAdx47+vjsxrBgFMOTcvmrLPF5k7vo4MCPbKSO
QVrB+2x9BPMmdRibYn/FRmPBnN7e98JQNxTH2RZVlq7QpSg+Zzv/RzIVKos93Fxn
HvaE9JkiMK7uoLLYSnSmXWf1fQuzDPjBkmHzf/oSk8uZlUUmhM1cHqrYeUQXan8V
0/eEUqp4PeE4NaEvN3YqbXUR7Xl1qm3i5fpWA3n9BoiEgUQP314SgGCuvWspB6ZQ
R+WOacz3VCFWKECzpnVq/AQ2zof3XmEl5raWwxZRjQcpIiTGrc4JplKEfGMeDWaJ
ZqeW3ALb7vB9BjbNf9L9VaE6yUvb6u3ED1zqGVGrq5rDRp/fjWE9o6E4URyDWLyk
sXYNcDREt5e/LUnzWAkA8c87lpOYiPbHisukvhHiYoVFjQJQEf9lMc7p5QHq+0c8
PdtxjXZEvmbJqsfWnaXe9QgM/h1e1UFwVO1SVvo9dpIe6Z3wDaNjLAQ+ywL1Xcaq
oLfYlF5m9A5SZKxT3DCEmPflwHyhF2LNPs+aGa7cHdEYH5LJnELGcVSsez0oIAdi
rP5KPeyVEou0fcqpox6/OnFdz3eU0QB1HqWb539HyUGx6PRhjpsW0eAFgkns9WMB
sBBpM0GsYk0N9MdnCa3yGdbbO08/mZ/2B/iqTiKpSpJf5WrBoSVRh07PQk+ErR3w
+7N/fGBCpd5rkt70b5pIiTNMlg2k8zbPGjNjCh5a6uX7xmyScH70Zqeex1DRZkuQ
ArQh1iWz08XeaMtuR1ac9zH0oFpejGfUwvnM71lz4XcDIe0ouawfsAQsQtnpiFf2
NFzaqUVkyueC42g1bRe5w/eK27AsWCnJxgdi16AFqhNNOqCCEtJiC7xlwl9uPuSp
iUlk9qa/YtnCOapFFsvhF2WYwcuUR20anZPbJIh2Z8Wd+R44M5polpl9lnpBy0N4
bK3Mt2Nr7ssGSRkVabzXHpSpooMgzd+4TqHTd8EYgPZclTreHOtSUkQH9msgqgWk
Puz3Xfemtl55iMZbjSeM30J/Q8O5/7KaFxEscJUb7ZlnvL/lvZ3BO+sUOC1FtpDh
gjqkLKOLPSZWJzkigJ3nERlmcPoHD/nfGVpAb4ga8a49JNUdS/Eg1l6VJMku2t46
9yYxx9kIFodewDnPuQ4TETCXC2m4NdO5wtpLKBJvOFPy//btK/xmNBhyGi8MLwiD
51zTjGmWlTOG+ltStdgsbEOjmum6Pqps1u+vSHY/OVg9hHCdYD6UeDiqWPFqVp5G
aShpdLkABR32fHEdLI4ryu24hcAZiHo+AoI1S/N3hLrfB3KaXfQyKaW9UdTq6+7E
Bzuep4roMuKgvpD1Uuq2DHN//58l/1fsNRaU5ffwNGontDfpHn7COR7R0L5xaEwP
iuiVFKA9RjRabHhnnlHt/qLyUPh5a7UY3bnyIC5pWA2PJbhcrFOfoJ8uKUCWHiNv
eTrw6NKwvt9PpUy7NsF11TXhhTaOzUqOFFDhJsUiltG4RLqyZ0Y4v4pwo8ttglpj
axSmQvt3kgLZFZMb/kKODDVV2Gym+HVQWL70NhwEPMIREhN1CV/xRgAtgVIEz+0+
UhZVj3932RWedKDSDcuLL/8Zd5TprQPfWq1UMbfsHX+ikHxxbfqkR1+h1KdmnFCM
Rfrhwclj5OqynsI6XLWwRB7BQ+KhBxnp1tLXov8MuJFv9Q7RAsi1eTkKmsiQm22A
6PE8OqXS8WJ/BE+b9/oqlzmN8UfIDx7jjcZ1giwKh3SBnVhvH/NY6gaCy3DAp+c6
ZToA3CrWH3XWOwkWswsr5FMrQNpVZUKNUQgjN131tlBW5GaO+JkbSp2m9tA22dC4
3acSkR1XR6vh7qSTbpxnprqCIcyOizA80TocWVl7OZJZ7F5FT13tIWDytiY9ewoQ
SVYPWQ5tITs8vPvJ7o+H9ImT+lm1vY7TcCSRzbrXiHRFEaX0ux1N1MlZU9T0rsz3
V7Le9/+nEcZlNbh3fvTiiB44X8rZNvDkpWHmn2VirgdBRtyQLMohp3fMGqqvNOpf
ZALORSNsxMEk80JI3xoqLlsdx8PgKaBdFqAMIF9ob0/JcgdSJJm2v29G7T8A8amJ
zqJdN29Vua48G4D+jNf4eRV+egHsIdjrYt8b7B5ak8GEOZYGMIZXNrThLFOoWAC8
qw6qKIKv8ucuonYlonjXI+DWhZ6kRkd96kU1UI72m90fXuP7jogSTpg/0hny9oGF
vxd08mCsjdHtbjf45wOCUPwUtFwPe78Plnv1NWAcZicGyB+ZEqN2Tm8omEdkXA9y
UHt7kgBXkEJp06J/FuAHvmOGWabLzhlEvi7OeRiIAMpFvppZTcs196dLSd6ZNrBI
wPGq44Tw3g5EFh614b3h0Fc9sqmU1YyIN1c5J9fLP2XgXWx2MN4ywhxVNjSNopbU
YmoNU+xSTJbFnpUPtuU4/esqFu1lAavoDTLLZ8JKZLWmVE5+3D33q7haHKIBV+ld
0+Vv9C5o3kAhumRCvFjdaOgWOMHB/1zXbeATvVpRqlBPtFt8dJYHp2vw2jGf4XPq
q3pfmJQsNdNjhB2jAq3TW3JpPNsDHttST/6mSPs617/4A3O8Ejk9csFQBgGA2e4m
oyxqCUpXN+MrXPNN6Zl65T2rQV57twzZ4BVj21K8pVAlEddgHr7gX4YzRikiPVxj
xyHTObRxj3N4OjwY8ElXLkJgSDwdmOOTs5FY1I52mdPWoCnDUgUVK+CK1Ku11VaC
W0lFWbKdnEl6NuJL6qArsA/+WrDrOtbtVzsxRxhPYECdgWE/IGmKLyl4FbueYriH
M8FQEI5iS7SRMyD4l4ZK1FcWmIcQJQ2WwSKEmwSIHrBMte3quMFL0lnmXyopPUc5
7dEB2IFaoUn5Qzscsx4mI3pzRP6ENmoA1cEHb4olG16FJfovEaXf2d7wgaC3Q3fW
oEc289pDUC62JYSHkc+WJZRz7OTYY75AtzQdX4tEa3w1UF1bw/3xxqQcrr4efKlO
SOiilF3Z6Mw/o8EmYI7b6vHIDVxaU3dkvjsos7AsYG1smcpNoBLgQao/6FYZtqcL
1Kwjbuy4hHSWRv1Pc4KzES0mLh0KhCVtqOEpxygJZIBqnc1UX4kzcK+fNHmr8tTy
18Xn0aepVD3RunxC1mHSJOqHF6kkq7X6Jpllz9FgGC0LG8rn5pMNvD8RTBt7+6gN
+5RoMgCnXIQ5y1qPmSB6tHny0WVZADO8wGJy9hrwwNLRuFgEyOfkFjNizUh4CDDb
5DUR9GfEBU0lMqTtXWWfZGYibOMRkIQZY2b+OcVOKTa1j0rkaik+XNPPsqIAtD3/
4uFl1lX1lO8m79vvHE9KYPszlEi3eTY1ir2VQU9AirQ3nzcWTcKeHE31oO7tsjd8
/5jLwzeF2D1Zak65YvNfdXuMmJmiYCHONmghs03NXQyXospHJcCgckZryXYroDAu
QPRHAB6Vr3SxpGwYFIg1UahLDvhLXJj8qgMResbBuh6ls/Ttg28BeWR/NLNLljQ8
GlClPSn7XCj9X7dtu2Ol9KE/f0x888gOL5sK1RoBJV8GVDJNBt92Dty5sjTAy/6d
8NFHC+T5JLWMjfQ+T57MUM4rWztKt9iqGZ5gmoyRvcMeEAaQmANrAH60ZkkgJX1D
6jDqdVRZF+xabcldyH+pmuTtNmTd0saZEJDJvApLDLDjNIMMvBJjYieWHZLXJxEW
MIGXdQqeQSnGpAfBqx2h46htf/iREDJArLW/9TkxJwvFLKxXKezhbOm97USr8XDA
M+xJ7MDkgWZf3rlQ0r/bW9KXMrHwZXOVzhQQKJBhI5wNDuJgw0XihtXexCJGOpCK
SJkZ7Ec238WCO2gslwOeaUDrRxaVkuk4xfKO5fzS43L05oNc603H3+TsVskjDj8X
PuZd6FwrtkxJiolISDjPEUgh8DoAvsU8iHUp1ELFErEQb91hQXHmUgsRFg//GaeQ
BH9BhF+Us8G0IQn7WVNM/adLhOTa9Ae8e9e+j6HjsFjYC2u9c8g+4ZrXNgPzEZqq
XHkgU6Aglb0AiukQ0tawW8SXcbXqlYkAsXIbIGuTvMp6Z0UjQ+6bjUoa8HTHJOHc
EKTmOd2LYGu73AaTwFJmEWisAZsjBPtM6S8oMasSZ4JhR21zqgS/F9Cw7T2hyx4O
6l3fk6YtOOfzYJ6yusOxpb3XTvKyyb32rWqOLfWSdJElR8soNj1SxmTGmalM0Dcw
+YqnDcwFNBsx4GrTiCmKQ5FUrtMFnoxc88HvKvuqPVGeh4WeyxztrzLNGs4e2bLs
pg7k/MCsDQPXBA7HpA6Zxao+73UyuqIe15UVqmYibPWN9XU8l22ezoflJs3makTY
+zehQsR4CPa1pRijdzm7z5FbhOPN4s8wApOPjZAJj6ZvYIKKblmOQq3jMuOV9/sk
qFaO+9lGm5gUK+hobbjmqrtDoofJyKrL8i+byy+5wT1ETtjxbB4K0PYzfoQJd9p7
jpZ7MEYl4CbT+FKZwa04RLUyJ6HKEMc7w0tjzao4vtGrncLxE5ztvwJ46IgX8lIO
mIbA5t6Owj6GhdxoSVikaxOT+Fjb4E5r/a3vxEfd12v3Ab3iweEpv6wTYGpHFYkY
iuJjqjmyvr3xScdq0Jws1E4yLTxXG9Lu9CZGDIEdlDgoGOALvgJwqxEukQn3r37O
3p2/8Y2/k1w/Iu4LXOtNY2HGe3FLWzH92VFQTR9tGXM7SLQK63AzGQpX1KdwmAMN
n/8pAbvCC20JBYz/PvTWbS9s+G78HuG5c0zMsNWldYPOc+Kh1pjvIuiWfAmtIn7p
B+YQhRdIQCWzH24XIrRe9WgDcVyT2LyLb9cpl7kGwuCUhS+3SCs8BSmuqA+9mKcl
vFRJMGZO7C3qbGm8s2y1WbQkfbk2FUHszPtk5X0QGEO+0nkup3xR0rNEdfZKxBwp
ProtnKNCVW0/k9yIp8DeOmo/3E6b8sUbbN5EdZJHLlK7LRwIDcmiFjzmjVqadJGp
/eykah/Kl5JvTj9Bldy0fce/v/L+GvGZfMQiAjxJwo1XfhzY/GF1+RtKyDpLly5Z
5Nd5aIenomZ9TYx5R5CKGZon7v34QQfo/1DayVVY5Jhh/U7EwaWlNY6DuDm6EdUU
Kv0NqInrjQASzqLPd0lTjDra9yAOVFbwblO0Koew4op4vHKeS2G7JcChLnmkD+6K
izdFhoCJ1zRcuU7j0Z91b+T6W61ApHkq1ZDgUBgjee1tppO03hRWggG5O3/+vj1C
PWODEBeJiqf8dwjg1j6AE1vqvs89aE8LL7rU9eYQ0eOd33XdQ5BFlG2B1gi1Zerb
wDMj5qJ6nMYy+d7LB6WieEL1IypFhKvOfaPvcTYpY0AZueIBYQ7LOQZ+B3YeZ62k
q0CaQIeXSMDod0+nj9a4nXRHG1dPuCo351tbiLXzxXJ99ZjDWMq8MkvkG95ocmKt
WGkmLVWk+Znephb1WDwt9SmK7F1MUjMyafIFjtVHnLeWYVbhm29yLNRwcy09+Rqw
ogJZS0MfcLmfhItwragGX7CrSTTW8xIZESSqCu0PzlGOt25x7IDrqZKYZcbgFqFJ
8dIXqmS8mApsrbnvk2S3bJAAAq1VsHfd06i0N0bt5eRIl2I0ydLFz150n2OcFtWc
gl9DD+LG6ABLS/rzRyH9rBzHHqDcYTd1Jgnfq7mrWhvzUFOW65y+E+Em8rmv+F1L
VQgBMG16FmnPgAW2kJLg4Tibmtwipw58LCuokaZb1psuLEqXL/448CEe7jj5p4pu
GNzRbXyYICC1YnUUHzg93hGKQfuKmW36oCyX7iW5bgeWzQh4GteWRp2xMpupF7lu
JDQwo3Nu8lapH8sZDebQ5VSOrXl4ZfWhMSjOxyTRMlbHRYpsaYTqtE5tkaaCf89P
WN4oRBX06arPPJY9Tx3fkgCEjUeoFxbewx/OYyB+NTtjC66HZt6SkJpFTHc/5uTK
niXrzAGHCYdDDV54BCGNpspgTOtn7f353N2po89/m7jyt8KYCViqj5MUI/ooep/Y
e+L18X8N/fVnjjnK3K6g1HzQ4TZeON00XUxfKr+v2Znc6+xHZCQUJksvM+nYYhKO
U9ANObPH+B7rQw9o0CAvPJdeQSt2csNw1qg88q4rT2hAH1tZ2ER5inwKNoWfUMNP
5B7kVPqBVYsYCYLiKnd7L2Sm8JDkJqCS07gxjXfszkPEPWkoXP+OFoxf5gd/bx9C
zzOGDMgLDt0lKA/8F8yxJF3wL6TowXM4PsLn/mZI6YxhGPTGbUN6fyHxivE/9Bvq
Du2EhE5P8sB7ZYC78rXsq54UMkHhmPkmtImc61rmvnV/D0iryg0fbvrPfiWmDuVF
iepgQgXIx2g3DixgpDEaDQn4uXxr6zB/cOsYQi+NKvJken9V62eAuxtftAi08Cx2
G92M11miwKIKptTA+i2uBLiukB4YGruEi6PIs/rYLBKZ0RmF86DWPEIuTeshUj5c
quK/rDSVNMPoBxE3D+61TgHaGviBAg+c5hczD8eP3a0TbSAo0ojN3itiCxSPS2yo
3opLZnpon4p2yF/rVBYRuoVI6lVtsyvjiCf5+SgBfMTdEBq/uLVJCzVGbLXFkSnt
Av9MZaICatYYUnjlPyYdkBspt+M+8Bm/6Cr/d217LNX6vQel9r52+UlugrNzVKyg
NSN2QCIw3z5TUgwmUO+0/Q==
`protect end_protected