`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 43504 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
YvslINJcsdDabhUxdg24ayBYK1KuWlzBVj2WOVoyLNrNDydedPFFXXdeb/WQ/Cv5
Q+n5Yh0xyC/hkMlGLBGwCUsD6fxfrXZYQtpwqvPtWfmX8XveDFnIIvsrXN2gM/DU
t9xTCEo4kOhhNkfnXUOHpD8VauDTdBIBIzTt2KWtGVnXiPNVD3FluuC5KdQ4vmp+
AJztZVDFQcckL5bGUcBtOLAR1KoR74vRMG4hrGKfjt3csqcstyJjoI34wlEIXmpL
nhG/4QauTYR39YbwZorV41decWIB3wHDOGB1wnq8CmRaUCSGZhhaFdM39oeX1Bln
zasLzVqqv0wWzByMmb0ZzkQT1lQRieY9A8J48R7EICSC3X3/NTuBLkB793gCwYiJ
Bov9Us975Msjc+mSEX25Fz1ITczt62wf4OP0iN/V+081qJOLerHyTR6YcxMNWuDM
aTDsjtnnwcNWTdyayjXsya7KNJIcjvDZ/c8XpXHWqM0LOxd2cvnwijPn9MKQmsWt
OoT34qfuGnJu+Mlf6yVwIFyzC+FaETX72ZZHVYK2cnjO/Hmky4JpLj88qUwhvO3L
aPV4DO5aguK/QmOg7OAVrMc1aJH6K/LosVront07CLnQkmR9Na8EM6OK7ij+jgEq
0UJNa1W7T9YpsfMZAhDYihoXyOjmaHyMKtBc1wDELODh4xnif82HsYNGsPSZTqn2
eCT4S57uGgdfw4H85VjbCMemRIfhfvAe8+Og0mnXSFyPFS+44dshbMMqfZAXE4df
/Hld+eXnDT71x65prWQQehUD0RFLFD7eFHcNOf0iDyBnNi0O3IztV3t13JhF7Mdh
BVe2DKidRvhf+EbWl5UmzNb5MgFhnR7UJaN7YaXH1NygOSyibzWlY6WOtgpziWB3
+T8UfGLDG5F1EaGgh4vV28lywpSlv2Q2yGXpXUkN8yfZG5D2kSE20uyWRynz3c87
j67ZaHsD+y4JTWIs3RioHKHM75bgCEo+USh4/o7yYXacrxCsj4qmpnjxDoZr1dSv
klBceZYxg1ib98O8GLzUtazPC0CxisqbYybazotMQWGQ969C3eCNjKHmr7WpWqu2
d9xBlmeaX3TFFJ24zA1rNvxi0BUS4sS6889NwxawHvTUDMxF9HbAHkpOV85kd95Z
5EzprxbbR/3E/rnv+rcRGWFv2SDnnGDTrWJj1nyqPITpr1zFlRq7+qiaHBLmYWa7
3fl0SkeRWmFn9e7fsGVHWeSJfnLSNiNknxCvF5Uw4JtqNwm/HeGgEqN7lPO0r64a
r8eWZ5MEdW9kk8lJOGj/alYeGfX9xWc7+8IVUxizoPc4el9IAig+vz3lK0ktzmtf
HoF0cx0cxiu27uNP/RG4FdUyyWgI/ctVfoVlBOPUMd4oOcbNcAH9PdfOyc7khk7K
7g7znhSgJQ/XTMtdImEG/PYWRLCa98APLCfr+WX8Za+qPWGXTU7I8qWVOxjw+nWi
xZlcIYwiqPapNWxjJe4tByMaPV/e29bSYkUCNTxnFlD+nxwpLZb9/b6rtKgZpoSP
QCfdVfa8npPPmX1F03S6pc8SHNpDp34SppiYpi1VbIFPkla4ixqi61rNp3/zCAXH
Xl9LfyzNvQTDFeVMDcDR13/DfdP4QmCWSnZ17IRBzUYGk4cnbDsS8Yvob3hpCtUi
y5JB2BgQfWq1S/SMpifzosCG+R9YQWqNvSz3ScLeC7lVlXQ0vnXbGK8b6G5/P35u
3U3m7lJdXq7YJkWVSEKvFA5Nln3fwiKwaGrDaIRUPDjR5OPTO0dHdqk9SJBIdSlx
Nti4dNZcFqFvJDsTeYA0A1NVSqzOZdGLENemLnqP+BOzY8uOmRCZWvri7ZN9udz3
Mk5Hq53XqohOGGOzZKMnh9BYiLB5CvUy2YezauXQlwK27SNOiXFh8uzDJoaE5bEZ
Ns4Oe5oU1w6AYjFhU59CLFJkP8uwO2/xP8AnhQVPiQosmew/cbD4QeQ6bZu4hF2u
RXQXMMtV2tpzLi1FD1/siIR6mBwyK6gRwWkGHaSfOkG8/itddpBwYHJAiXP6Jkru
W0ZPzZCXcDKVXV9jKeb5y7FtKb6CyJv92JDVQKE+gb7h00do9vtqR/4/LYmE/SUU
7CXO8sWVHgGCwH47H+vHWROvXSGd5di9O0DuE9pjzMaIT2asCr6Z2EHeWH4cjsTe
hYClaZPNc1PNGUwbxmFVeoR9CQkQZ9zuAmXQO7Wf8dISZ4zTtcl/8wDHqR+KMXV/
KyKLqiAKhPsk7ctqW0F9+eVdCmjHdIemDMk/Me8hTgsHKqSDnSHJ/rLfieNUOWRB
F2LyaI0UHSEtZxkIYRaeOOrV9UFrYkf2pwM8RhofI9+BQOeE1Nv2B+0hnojFlKWY
LAUQ4FAx297XyPB8mgesh7bjK4S90g8Ibz69pZiwRN2JBd3eLtNaQSoEzBNMHscn
054rhb5/BTi88Ld+0D1Tlq0ccJ4Wd/9ja762u42aRAJht27rDTF1a4U40AaniIMI
M3o4lol1EGu8E1yDE934iCQdTX1k6rK1hcxVf2mrn5/w3B0JoQjfr5rEfjNhFzMZ
nWYUTI0l1XCtWHU/DdILTJQH1NGe8Cm1zDu+2krJ9Fy2OJc2cnDENVnq+7z5kSS7
LsjZnW5OSYRG4e+bIygGgns/+JcbRe1ibGhwPoBhFVkGXv9+TQDyvjFHBliQSEzQ
e4hPtkTsSBt65WJZKLXciXMiR3zynIgbwrANOeszBM3k1edZeY7KyTozM8ezNPAG
r88FwBWWrHGqi7yN00+aon2ueq0l7lIZvDbyQBZSla1g3YJRV8lfugBpjzJjnfeG
CF780H0mv92vo/oAmByZgFan9Gd9W5jEcLJww/A1LsY0P3XEAMUC5K9fvJK8DVQT
qC5S9j/VGyGKlanzaJkm2HqdWutQXVT498Y1veePKXHo6OKIWdqUoALWOvNeA2Fn
R405Ftd1dOvfgKslRMwcgAUcgn3D0eeFmhqRGcndOwRTXY0PkeqnxHqyQ/qqDMH7
nLRMTJ+NGGXt7uCThc/GuttJ6sVtp8Pw7AKOZ5cQBQQrBlyikYHbfjncL7dLmVgv
LASbF+dCuQaNNKh82nnG79ClJgZ9Xwec9HKHN7ON40e9wSH/PZfuo0WRxLC9zPja
z9YIs5lkmUGPerWmaxwwCvfoVVSKszo3SicRkAez4MNo1as8sNv1IJ0tZCSWH3Bt
dKwCfar8UTAxZoyZp6crIcc1ofyDfhFJAVXt2ylGlZOHOGbXh71VgRJ/GzGzlGlf
fLOmuN8HChgnkJ+aK0Y86YuWvoHEd15r8xSjm3XZ8YJMWE+QKBwScPLiej5ZflML
aNXHRp2LMr7E3yZUrvul/Yb69aqxB9h4HuiUNg6g/uhgUKZdJZBe59IxkEWjNdnr
QvyaEMfj3hKBi0FMW7yxg/6Q0N3h/0mpGHI8SXNZVNAmnA59Sqx5Yn5Y5LY9vYs3
mVYTjIaMrvmKIlYEI18O7q2+/pJEzZ56vvHULHUJDohUsjkTe6ceTBpEnm1+CIKg
gSaDDzTUmbY0BAZ3YrlxWOqprdOv20M3aiRMD6KfRoQzkvou9f6f1uMYWsbavmdJ
SuZTHrPCjuPS1Qs8tq6hOXiAUAfaUWPKho88QirObE57k5/cdLlyWkets6y8Yqww
OwIlIwjpVAx72WXstT8ze/pm0d/JuZk+wvGkC+y6T+NuUo2z1VfzNGnKqgTMAEwB
O6KuyI3zbdV/ApEweBDqNAQNXkC2if5WQ9ZACjrcZjCt6ZUydt9/Y9AqTUav+Ea7
HW+YvIFHTQOe6R0Vrkw5mw5T/lrHYcG3PqqcmOTQw87o/fnX5xdLeMfrKdfPtg1g
Ph3bVzDc4oA0RaHAiDfds5KdkDQymWaehrPut/Iq0L4lHb061Cz227oqTIs1/rBH
c9fcog8uB8z2JuyjplRymIbAqUs/DhIKRsesjCrjlx+hfZKl0KxwDTb7qN3HAbTp
w18/E0cp9TK35OEkRASFUhDytwWhmX8bpgelpP66afSShwSesNCtU8Nc/ZEoUswi
PNUXSyIb+2nb3yAl+AUWtH6w2vppZDWNueOiE52hAry0CLEhZOs1iNW9SwtPYNfd
sxG6qNW0xGBn/v05YIo8Z7MUsF2E/BkLuxMbEbQS5XQOx1HG/vs3Sw9QbI8eztHo
qMdi9EN44gl+Ggbjbub9vejIs++smKxxP+bykBH7mRuqJcDeXNyzyZVIYTU/yp01
VHh9EvhXicPcfOXdp3ui7lSR6UiOyicyYNAAXmWdk6bUa5a1fvQzMI6S78+Cq9hV
C9ae72MF8R9AmeilnqUdFzTwBcVd5G+X/YesdRc3MSz2NgbjQve1w7hc0GBQaMs2
jmk8SBX5kwUmlmt1NsFOJe4alAOHVQVDW8gjpTsV28R7Hq4mNpz9YNCzklbGb/C9
Q6mfaAwg1l/nWdEAapMED5zAmsvy8ncXB9/7uFve8KnfPixKdlLkpD7E4cXlwVms
05AZo3oDFI0E+IlcJENxlSvEy2YaPp+cyb0GzJsYKzKZdsMi9O+aicZ+Bkc2r5vN
q1AJhchgdabGXy2VwNkPNzPT5UqdIUDexoFU325XTtQnuMdDZo1c4Zf28ZdHXs3A
AGZW86J9WhV0xaThhrsABdA4lFhqqCMQtl7b+50iAqEfX4NEpZqzbw1QNJKnpClY
o/7yrNImiakDyArZMvIkwut/i4C7LIYYesrsvrS2Y3jLkcOqtCbwXx+yHRsfG9S1
UG1Xn03ifdwae+EdnXgqhbGlQI3/56LCuqVWNjU7PY7zq28E6H4X6TrMA/mcVYJA
Mekqlr9mgOz2xoW0M52CqiYteW/K8zC/g5UGUO6Vm21gEuvJTunST1CZOqM7GbWy
IeClQcqsVU63+vRrUvfrRFz7gRqkj9oOHgGv86AGTP0ZEG1EZCwLfXbpVqYyNocT
8cvQRRQ8iyaQRpnbfkWK3YmMO38G00DduhSl9bJ4MmaRPzrl6KsmBX51yuIvuCPv
nyDf02DxGy7Ab9jrQ6JXOXVzCPdlVlxOnrL0Fb81PogLnq1Ndoizq09ps5ccJOew
AQ6mhr1F0C0eU8RNGEghyHtMajrsvDxanyXp2yJSFW4boOTbcIVAtRqlZoEH6bVU
twRt1rtU09wCjEXK9jzcAq0xKrelvRg1h7WGUpOXb4+Sab29XngZyjaDFLvjADfF
IB4lc7bwisW6Csis21ePCCbecFVz95CzIkp8nyrCyf806Peeqk076xaDoa5JlPYr
k0EGZCB7+tgPkDkeTdUklcJq1jDV4uSO6CRE/REayRn9TOKkZD6jm4Up+QOmZszv
R6tV55QaTrklzawmId+hsivFvlarwqwMWVTQUtdHDd8yNHFbxcwVwWJlFpyUBtBr
Sy2CgwnvHHml/7svewcQQ51AL6Q4tkw7iyPfR6EsRcLrkKTYUiTYdo6CccjIFJO6
cQZaEHcyjjBLLz4GbtaXtFnCV8+9sZ5cL8twwpRyz9cxbSfVQM3OeAFDmJ593MuQ
KAXjuR/RdqG78dfbP6LFeP66IN8qAme57ouaRqBagR5Yf8uWTQsGYTUMyMsLM4kG
67ZIkIKFdoF0Ks+bDeeE/Ey3LNGlbMek3XuuvnPLOkQSyQ/iHEpjWnqcDj0fuPTQ
bAOf2JIZbWxJuYZZCI5HZhQkuuu3s1yrr8IlRigblZYptyTqvoF2E5tu4mYBN61S
acyuKGFQjjiM57YYoHUAb8TsQ6BVeHYUyxJfnMdfChv7Ytj273L5JY3g1FXOkG7k
eYiDiyuJtiocHKdkhI1hxHPQObgx4AxiBWnsfc/sehmIACoZRMC1v86MVxgJhyee
p6R5L0zUDV3ib1hAf4aSgkHWOznx4uyDYJSMYaSog8ZtDMNU/Dkfc183BCzwlqtc
r6M9Bat5a6w96sDudT7ih2u1C/b2fdevQFvTs5RN/EfzqgSF1qCovFs0Aujrcmqv
JLojukTy4EoUqxF5AJCLqvsDlPiHRTRJYoLzZkNw5TKVtoJDUABghS01HVwseZKA
8DN3eNNxgEX/8HEYIlUUKDNVEzMzbMYCX9gREUvm8GiyIhtJggpuMGu5gWQ2idjM
dI4/Utl7PqF2zypGMfBlZzXOLCMlUHIEMqk0vxyNnng2RjtqOgOUWEzCnIsxF+gY
2eieqpskiE0zScQrCQwL2r/8kdDZ+fJ1T81f1QgaoH4xow2l7EZxwEpSxA4AAjJK
kWKe8stwZEGFq/arcHvD8oCSCGf4UT49Vj4TdJEvKm3wr3Va3lDMqUwbF9c+DSSq
XOh7RLrzdDhJtPIPsDcyiZcBR/2MYZUIZzNDJv3kirMxy3jDbPqqktdxc/vtA432
CzMn6Ct1cbfuSKcULXttj1J03tGF8FGBzUAb32pLE5mqyzinTx99MHJUX78JDKG9
I5C+c7LZTsiLj54GkQ0RL/UtRdyjV+ZWgZ0W4/FboGYcc7XpaivdnEJB2HR2vkra
9WM1trD5TdsBijeLR2I3b30treKooyac9qxwFwz1vH4DLCRhMU4eZm0t9uDA9Ugj
vqFXnaQ41uUmD9ueedxAfqjKmhwpwWryZ+2AFY26ButdJDLkj5tPY89u3n3JI6m5
f56CfpAiM6OPKywSzSWu9vcMBkRhNW+F53flHWZgGe4sYC8TzqQHIrmZwUqf5FGG
Rs4U2FV/RLA+3mzGIe8ve99XU/fU0HmsplTFNxf8vHGQkJu+w2YcVXGVh9G+Giyw
pjqHGUQ6POY5QuFA6aWt7jFeAgcmHlMu4giEdl6UU2eZPMCjmtqs4ba39CpcEtay
y27KM6AsMPPoKh7ck7HVzLCM9Ky3taVTRghXjki9SJ7uqOc0MtI5s05eQnmwFZ0z
35MKxiL1QfRteLkqeLXfNTbT2+r4/7C0RWcMunwt2ZT790PhrVogWK2DTBjfrFvY
nbCq51CIzp2jN06bzhKpgLw7oFter2sM8RD+Eg5EKH5sZSyEVYrupFiItJYN460Z
Vto3evCBud8Y5QjR0gjiObvEs0/LKR3eecZhKbHR8N9HumPA8N3zSXiE1qVEtwbY
MVtF53Re+D145AkNDgrP8nPtfdWphsMVpKEWAHdhUspP852RC1YuEvKPOqXYpFRL
UcpDTkjWx27c8Oevo9oJpjlPNorW2HsYV+BiYpkCzKVHX6ng1rxJnb2P61QwCc1n
G3LxuZ33U+VYITLS0T6kA8RtaKoW6aUmexm3Ngg0gCVa4NbWaOKjo0sgvfHS2oAB
xG5G3uEcZBjoe6hAde2pFOQU9H0b+85iMzvHIK9kEZvLjtE+cDuOUQ1cF83tixMB
17d5Ozwwlai4crXxyE5xp6WBIE6fwTjAuFxcUGfOQ2ltOJqbT/ZIbSJXDSodi7yV
c4NTnpimg0AgK8O6zV5JxnjbEspmMUFANbWwesmap4QWTVWYugJOggDXrlH/T21b
Lz8ZmTTcYewP+noyEobARh8S3Lo577ZhuNTyLFBLOufOdefKZNdCTqPLu1AS50Jq
qJzjvt1Edm5aql9+DsdUyPjf7aPhgDXyMi3j9cZZRi/vZyY+5ivQKMX/H1qPhci8
M8VPZJgBwvn9T04UrTZP1krKwPrq2KdTUXsCT0D/c0GMakqgfY0pV05eeRzkiZJD
T3N5VQbAe7dWfW7tFPCeSS3082l6WaR4ynWlgxOa7JgZ1Y3NtKH4I9pqYMYoOWvB
GMnvnWiWBERLJcnuRfwGpjgFwnmsmX7qiEQJLofgptFRCrUpq/p0KcoR4GBhThKf
1gVrhRkCo1cCIOKLzDNRWl49aGYscBUNGQKLHkJO/pOLT4jMwifbKDAo6REjxD6w
PUTc/aF2fLELNxMOkKYX9xJNZOSisYZV+jFI30bRfX+Mvybtvgnlvh5ZLPTSLqC3
gFNmVgskZEwkFxcu+jNqq+iZdXeejqsu5r8NwnZkQa8ErrF86m34ZOKUEm7Xns5n
y4od3Ve/eOoDrSCo3H5GynAvwfIDOFAUAvy9qnGKzXwTYRjdOlJWB2Str1cXD4Oy
NSvpF+mG4cRnf8CbrTxsKWiq/+Wbiz0du2afe85Qj4WR9p2CKcoOQDX2b3jmZ6a/
8lMMxxKR2CfeZBHPJ7Q4im+83q5oMvF4IlNbLrWH3dc9YjhDkQf5WIOQpJ8ZYE9R
5BRD1h00QSWv/33lsJx90LDPCIS0U6H+VNzlT0moMS+9bJCPt4LsL771MSaAZ8Vl
+UKyAVZFYI29LJt/yKhPvG2KJJUL9psrTX/aW+2E/myYTtoQeQF5tuZNxA/Xai1o
YeRcKlkIk+fzvAeQzfvyqBgGp0bVbvxpi14Y+83e1YD6+SeFkhia7zqefXG/RKFq
yv7Rrpo80CRMM+DhK3TX6m8TRrYETdZWKFlZInTbd4yJr3NcjZElwzD14jzbqy+o
BsnvrEI9iUJww/jIsurC8x4bTCO+CE/zeRnOYGX3wcRmHADa8MutyTtScuYvce2i
HV+2dqTt2o8y/iPwoYcuBfGduya5LIyG6JiJ2NAc0/onVQPI8VsUoJBxEbePHI3Y
bYYnAaWnBSx5vAPGEnlacGAhdXB39wRlhc8a3vOqnpUBI6zmAy3XDedZKgTaNOXR
9FNc6ueWjd2KMRuPUvfG75CHXMK3EFnbtriK97pfLYQygIPu+LEjX2aftVmDfMvP
istr8kWuky5oKFMN0g8+LS9XW7T97DCAG8OXjHql9j76Oi8WW51NSQ7y4lgmJqPI
VjtcuPdY5TOJFIOyelw1JIsS5pxQ7V8Vkiq3r90xJ9a+ML8Hp6L/n0zmORMLvXe6
DIXc+14+iOcCPfoXodqUiJAwCipBVZWnuF6AjkY+MtNfv5VkYORTN9T2gRT2u0Br
mbPvZvUW6+PtCM+CiD+e1QBCAy+nnxorzzoUrlmgV05r4/0ofofrFm3YPsRGbSNp
eKU+kH6fOZ5iIcYh2CseVDafpSSOqwsbve1XUaiLiKdfCn6xr0tRGeMlOuIuxwlb
EKALTnaZ4eE7BhCKCQjhDYkDekwbOW2vXQktJaZZFIdxQBm4IYnlt/gqkXxL7FA+
M1VbGFgGAp/h4yE8mwlte/q9CyPWZw+/axF426mstI05Vt48u7KV+qbMPLrh/SAq
OGHIDWJv8kuc1MprJ9YzzIyPctK2UHEQy5HEm+OZr3TP/DvJMySmCZpRHLRiSnDN
ZHOKqfhtxWu3InqlvLVv3p7pPoI94mb5T1nI7BvvMCBPuqLo3d3wMiddxEEKlPDj
K7vy6kNW6GEgNOyShTgbKnB7X8u/a64kdSOxUaPpnoPCnary+div4c+9FhFEV+VS
n76Iv2MWGIdsyer4m9jSlRBoQzpKpZtghJUEhCVKUaTQllh4aQV+t7kqBEPGJJrQ
5PSTSWuFvxg+r2g+ADbUtS08Z+nTBbMOQYreVpT16zDSbcttwzbw1aY/rIyYz22l
5n5Ssekaj0g9xWDkyjmMW7uohWUQqcC6S9JuF4FNC7w7Ox6M6pcnfDY0oOBUWHQA
rlawMMkbarvf71FniwkmZBtupVpfdRqlt/53yNa+DhdEoTh0HJJj1D4GpzvVFGdK
dpw0eHGwuY7knxIEES76/lokPMRiv5RIlZDvsZS2rQmiyalF8Y7OB7AFZHYB/6Ua
0b43faeOaY8Qe6p+Hhv1HIDJq3fkp1JBenVUsSRZ+Y6HLl/U2Xx64lFOWCzp8oNW
r47bk110D4sWLHUT7QwuHrZadorLLMu0/oMF/vr4Lmh+m3IDVyn08OMwLCHccYhv
XHLWmNCVFy4Av86Yx5oe6C5Ku7ZPcFholCxEOCIhrWrHe7mvU9tbnG+AHo0zjg2G
8mzqivMDtQangzdzLaVSjP3R/pmA9Amy7+RqHJhVLMWEGA9Qlcr+EmboYh7zpKiU
WuXjJlgLtBitqbaopYq0sm679eoLBEC6KIccQvZVkCGIdO/VnffUarBKb40UlCqc
V2+zHjxnTiUFdERGvO0LDiFIvanYzRFYMAUxVLZzEQuz+GNHIukuw+LcpNVCF/S8
53oL0G6TGvD0WTk1ZpB0S65c+AdFyOUuw/rkrWVAqLpMEXNnrFDSMQElTaVbV8oK
/grW2/ESWVBrNQvCngzjSbNqSRNKMp1yfBH+SKJ+uH2BP7Z90d+N7K9qOky1ArQp
aJfxKCgAbx05yAN5W5oatF/o8aIJenuiYgh8omiWcIarKL+90kgACy1p45nN/SS6
7KUF69+f5Lph/faJ4c3OJkSpRMS5NM7BZJivJDwHBTNCWY/FIFWQI7wk3LwqtLEx
jvGAggPCyZdabHjUDmZiBehbLyv5EqlE29ltKGBUt9OwmX0mr2iZvmc3VQ892Xe3
WnJP/UVGZ5PzYyNPdPEWmRX+Xha8aPfT3CoiTitt/LB2Zrs0iJY3rHPIaqpzAPN1
pOIBMIHyEOGKIOs8b9eqgQtCZzG1fS0v9YBudOKVPLb3WKTytI6Oi4ft7iZKCl6C
xHkZsQnp2bF8EqPCaQF2XZXcQD0y1PJ+dkYNIeJJjH9rSqTjBklzVqmutd9mlZg8
eArpb8ZXjh9d5wavFTKYuwGbbnaURw7pX1eRlMe2t+pOYBBnf8mCjt9/G3j+p/6s
6T/UgWJXQNSkX3e5iywHJH2WrANdv5sxbRddwQyud0Nbww9qduF85/HV+rFSdZMI
mqAUuFdal0utX8ITCGnUI4lIh6gIki3SXZgXfBlAXhVr6NV7Tgq2JaVwuhERZAAi
hUY3oNnf/iJaeFm6TOif+uwOxXCCyoWoAmd2IGu8tnut1xWJbdwgatp+6MkfpwhV
wn7JHiB0w+Fc/LqSMyspis69UqUjx4XpuYEx5eojONgBX87U2pXzUizo9tjeyuYd
jTylC12rfXWF/slQ0+KIXT/54MezTTgYihU7WrLlNgvktej7tlemkTgIOnMHWeLo
YY+OqZMeRffVoVT3xQi5pjV1cZ1j7nEBW6SN/7gzyZGNberjBnonMm+c54OmbFGI
b9Nhs4qSR8MsmiceH6bR6PNcxFkmp3fwoIbRs8SWh7BslLvmS/4MLudneZE/fvXP
3Y22Jk9RoWqVqC/ZE/AY69MTbdFmXHoMSmhgu16F1HeB8fOPdsRaJRkeNUkljhS0
OgudILOwIOHd4/PaZnexILTloBjhvh0CeQKY5HvHyXSBhpbptnAVbjCSyhWhD6Dw
le+Uh1WnXCn1bvbzA/tSiX94ngIz4v4ghEFdjku0kQoXIqf6xDJm3Sn19cSeqRTi
xMB/PoaeaCxHHSZCAf1TTJUDyT+FgKInzs9lQ3w+UWTfMn5LjnMhrgm5M1Giobet
+P/RJarKA4EhdvgRvMl074ibb5grmVJ5Ny5svoVa6G7VpLDkI3XOzCh3rKmtscS7
7qitYBz5jjgUV6+p5ns/HodD0FgoPSZnxMaHQzk2UQjNPE6OeBztplUEB5uIqFOK
fvsDwVKKvkNR3MXz6wk55sv0szLKEbVYg6y4AFy6stDRJH9qxPXLjsZLu2BnbNvW
32RaYXHvFe2H3MlXo5actLVEzW2gjISaFXv+4B01ARu/Q7dgtE+4KAEKEmJc0NL1
nobmnRycYObstNwbd5/9OzH0ntnTA6kuJgDP3J6EzgKY+K8LayK+vdw2yD6BovhH
97snIpgDqj0JA9a8G7zTkXJ6jxPJLXX3F3qfseNloZV89MDSdCisR8Eddo3d1a2L
AxoanUN3zDRrV9KNvd5KNtpGtJ4xOEpqkdbcP74KncxGBQeOwIScducWzXfpL4yy
IW+ogYVY0kSBFVem34UTFR8m4KHmfG7xqvOIC2M9MUOqsPrV+UdejH4VC0wX3+6D
8TJdjvrN/nCOVUjGCJ7uLVojai/iu+U0JsckUVuU29pa6jgWt2BZFuDAICPQ2ou3
dr2+7NDlFYBMhEEsGT2Jt6V0UsAyvr+Qx3sTOIU31vj1p5gCqr9UcmSIMpzePeo4
PYvJQg1wzaERHYOrUvZWPx3PqtdtXGrpu8qNr5KDhaslC6pBnu07yXlVegFgKsIE
abygDN5Mp/3Ju2estv2JAhr9ckdGKzFY6YxlpNRIob/33OXZ8eQAJvZfgZVSteY1
MlrCNndUiwyinKKmE9NM/gBFlc38K7kNLlfZdbInf+NYhAw1DztOpywe6s2VnNcA
ELSF0A/iyXyWr+vBAriUMzHrWAoEEkLfvQN7SmKLJamvBn2pdmiEN9/TmMHhJ1zO
q5lVlH7SkSGl+pC+HNZ87ovQO6CyZSHLAK8TtSG1CtjkLYbdRToonLF4/7LQwBsM
o/6wMG1jDBkpKbJJfY4HBTZt3XNVQaWKab4T/1dMoTHiL8SqeVsQE6WPtRrwQdFI
eerMsNziDHLXxfkqp6F9CZHfg4sPa8wrGJ1lE1QM51oEazMZ6M3NHCS21sTYDCkn
mnGGaJRt6obCcIxckyZhgkEd4HgrdJ45d6gWE51lj5JJkZixp8Py9yihbY5NRV7p
SP+4ZxcpTDk35qIUg8SYW/ktf2TeNWANnsHeTKEqgP8jBsHvX7mrVI4yGxIUC3OH
o3wx0aImbZ6+ClvCQW7hiV1B5joQVjzSE7FAuyNZ+7rsJGNFHGUWGbm7O1MFAeup
KimIiQNzRjih4n/bg1SvsgDHEv7UDosYu0FOMSSwzikRseERapDIlJnqpm1cUSH9
jOh6POo61eXWyxpjvbEdoisAQsf51Kd9twpZuYxUjdVLyMCv/6u/n4eqdr5GsN9z
Me7ORN9qCd74wrxlO8nUzqNlC1Nt+D3RU5hrBoVKb0//5JIiTm6Txe+wViZEIBW3
wHJSa/nWTAThc8B+6PDK/ngF1sC6b2wdxRX2MaIJkj0le8sew04sDjlAvatZu7I0
xOaZigLeEpar0aUL9999ITD6HpP+E1VWkcMs+LIxyMnbY4d1VTu+YZ+OYhW0j3Tl
O50doQ0TAOdln9MX4k2aRguaJRH+euFmbW+2HfCM6/J221HuFn/z3oOCajP4xVIq
EtH3ngt10JsERRdVjJbQT4L01nJMkFCJKsNgln253XjVscez3yJMgOLyBUKbfChK
irWU+wgdpQ6C+T7r52WMX4e9ivJ723LTxcAx/zneuSeindaoXOXcfMQJZZNJiS7B
fn6OXiiwV21FGd1R6Z7jmFrkIWaX1CDJHGAcDrHWOcpkedUakxuVTliElPxOUc59
t7s2DUCo5g61OH2vWNS6Ntafb3CdQmiXHublqek0ooBy4E1J4KReQOmZBIbmbUfi
g6lp+nUTjKNPvhNlwpWyqcOMAhViQby5DzVZGp/2A00xk22MloXkpRH8oWoG7MrM
T81WKdAIQm/qrPp6Mdeu4CCfU9Nu1bowZ4QltFjphmmxsuhtYzAyi9+Drh3lhdXh
JA7OKojTThnMcwwAMRb2zNYGi6ze1OHxsOTnRMG0Sru84e43BHbJU/6wsDThv06W
NW95PTmNIXze0RLOd7BDVsfY2K+IidizvAQMAS8uMjMrFnlZAcPtFOGCZT5+/Wgb
KRm9VhMMlAWQphGyiXXZpLCf5fiAB7iCkq0RW29ik98ZZQZW+QJztRsdLyvi/Z6Y
PCKnWRWo7cgrIaquEU0HHAHzraDtKNuqhI2o7u/45TsIKtHmmJCPDcYH/t0yd0//
P/zSKHiG7wwh8AIJAr0c2ibJQLZrmrEfECwLL3wOn17VWjKXbIk/cuY293TR515M
a0XQNh8bwy63sX2vrG3sdEfJKOb2xa8HgFZkDJqv8P0kAy78bbY+jdMEiWYknWGg
DIaDzQhHf8Z3AWfyonx2J05gj4dnllk21PsOJNnh2FfGj46RI3Q0EFThhdqLsceX
IfZhnphlObpPmbEfKqKRBIoSCcFMO9Hiq1s26ojh8r9fXYaFoyprjc+9xSjAZS46
7M2DBw+svM1EJsatAy/5nB+gOh1SPTHbt6woU5xd6jRKyotwYGiSW2Dir68OSMRy
Hi5Qyrgm+2rUSOEbBvO8tpQW7OHF5rbzAC7ge5cUx22EiqGAjHAOt3GVt4S/xQ9T
77L9p+sAbbKCexxkZB5NSpKV3010izCC8k2dIus1wukN/jFIaOFOc2TuNEOXOzI0
8ubPolKnn5VdccWbMWGqCctz4Keu0sFe715bIqGivu1vDlZwz8HdibMKyaCy8rQw
IGcCK4XrwkfO7cqqgjT1iOup/E5cg7KHcndZuAkZ+8G8d/t5dgnyJNiJzPomWZgV
9kXu1umhB259UZx+SIEFLFZwA1kVR+o5Lnj20UFz6A/lYAhK4DqlqMXK7Hl9rZS0
ZoLcJFJHzQ2AY3ao2Jgo2Mm+q1N08Wv/6vJvzH+Wb8hmcl2orR1eon0i+g9a+RSv
T3g4iw8A0lKzd5lAgdavZmVmHiTUv7j7xFyZkw4uZGDyCw+PiW9Y79kbEWSb5D3A
6U/ZJL35fG3kmPzCnlRsPJFu22D0Mtl3HFmNOTSata+UjFSY5YFsz7JWZSnCCOge
vexxjkDAxsKeF9k9NJPou6+XpPANIxBQm7DbvrhxmCT8c11CKsPBwFh2OV1WqgCP
SVJtCqEOgNVHpTeAQNmdZr9CFeloWgpFRsiAILQEfGmEo82lR2+z+Y/WG5qWiO2K
TD2+w9AYyW64mmIQcu6AiLDMNhX6Ofpfqb7LsjAG8PrOBGZok+1dRqrXj7b8DeGS
mC4DTzFte6Srn62hHJdOhuAqqFRvPHRmU+RXF5i32LI4V0QEbv89WfDdbKtpuf75
99f/rI2AY2qGhZc95hso70mFBuRyKmVJXwGiswYKgh+WM/BmecEnrWsuUp1b//PS
P3tj0MskZUHwicP3pdIKF4qm0iqUL64yd5DWl71cW56dugRz+ruTqMD3ZJwTTgdL
mcR0F3Za7P7k/bnB59+l+6tgzf2vHxKxK2Kthp24sW09Es33bRItFW91cVX6xLX1
FOrREZai6xTXDzQZSbHBflG3XIKyNv9FcM3MfG8+Sbc9yYwnJVSLywx67FfV0sMT
PiaK/0lwaCnA5SLbS4M6uG1FnImDQwieLgLGVrGvwSzKYUooE9pFwC3nwKkZPSC+
hEwwmQU12FCG/l4fSi7h0iaPAD4LtvB89XiYBKjPUMo5Y8gPvQ8pf3JBMJugD5+X
Zbdo8Hb2fZ8WygQju63/yE4tcJDXSjwrK7fSLe9hdhG5QaQPz+ygOBPk2/O4+h3t
8A8RXc2sEks6EUOURPfbNHF/7u83H6r7YDnvJfhJIoUY88/7+xanqAqb2AcCqjks
TxcAo/VAX3ovOMKix5+LL3+rmgJdcwl6kF6FCizmnIb8ibGFHKi5JU7df1ahqPdJ
7R3TMQ+545SRYcgVo/PatxM1b2Si8GTp9IGis0/cqo/FN03C4uINfWLETipuPXBu
w49FmcWA2qZdb7GL8N9QPc8iWC2vtCOn2XzvPb2ps3vbccXJEqa39tzx+Zoa2yBW
fdHcfOSM0sh/LhA4eXBTGx19HGhTHzLbvpwYuiqkzzv+Hf0gXfVBMKRcID28rzUi
7pspZm+hcHCznDpCa0cEeRKyeUn3BUckNevvEfnm3pG30kA/Wk48Hqx2WztFjYfT
XP1HQX/sr0IJcxXI9SRj7FcbrhZ3KDIrF6Fr6qRA0IzdJiOlv0MdVwWddiDPIcHm
mOuxWM5C7O0+DXmnSk9y9pCI8MAiUYh/OxLZmgV4dPXKrTgyN5lzEGMv/qgbDFxT
Nyn+coF4N9Hw0l96kTD7JvGNVzOtlhq6t5PnE8NALxJyCB48shn+5CN4zMCLs4Ci
cwHN/hz5PnynHPrapFKqvQSNfvZJ5MdKbrxANgY3WFj+24UmmsXnYYL1A1VubkO4
liU2UpATvJ9q8hIcUe30cHzNyNHs7gxwef8rYNjIXWupHmHOP3nLZj8ruYAi1Khg
DBnUANuX4YZL7pJU6vReL3UtuAFBVnygNJZK+ws42P/oK8C/kmBXYcxXtPI4oHTE
+z/02eikWs1fB3PttvqGUYpxeeI/Nr4EiJVpuoIWF3NEW/J5OBF6vQhjLxJSVACw
Q8FbhBiC3Fzo4pkdZNwCDPbcKEXGhYk0OI5pDIvt9MazmkDCwQItcL7PXdADaIFE
2wS9Lzra0YxXCSKpNDvRRc0CrgxPZUFNsipcbxbv9SyoGql3bbPwyLsEvJ69t+q3
VYMElFPLxDovSyq36Gu2vSRNYq1KkjlFpwu9f01Ij0yT8zBgR5YqFwv3s4mtbsUl
clGJ7CwKo0ggsMm+qAY7Q6TcfwlGOlk+aW/JHbq5BH0maA/EKFf5GB0ze5EIApml
G89DAzAibKihBaXfzTkg48med8SIv7VzPf5gDaK8P2yrRpJKXoIBGa0YRUnU8iux
sES/f4bWpVo3xWd5lsBuilUsmlbQWcaP+Ybt6VobY9ZGk5YEsZ+I17B4yq87j6Ys
7+lzWWWHJPiODOGky8+UHREpkvp3wpZhD9pdECnPZKrT+HtnOmi2CD1UGiZYpabW
O3nzEaFQ4l/kAU3yUxudHW2PRG4GIp5V7roQMU1W4ZkekXg7L3EhOMoshjc5QmnY
Y0EtrMI+/msSL89Xw0IeV0LmrvsHCGAcn4jF05ncSqZOeoyAvWbXtg9CcC2Zgk9H
E4WVA+PWp6MTkQ32UI2klE700p/W+tyhdLqYlFMbuMFDNdxIondfZneSsemfREm9
d64S7kJjCgVUtgV/LYV8NTrI/kEHfINACITihPeB3zrB/zSLJKTAvT+sOg8FzoQz
flJDyuG4eHo5w44o98VBkP7echKEqLivMmTLVeBf8xjFq+b47FAESRUtSh/xzYr5
k4Xu7awxL0GoNCptnKx+QdSZysJIGOJLvSx5zcu62HKA7rnihz9TmlqpsUjN16mg
NIheI0cxg3OzQ8jab1rTnAKLxoYrszwzcq4gJPnhSUr40B2EWKUxdotxR+otzsta
xyTseYVTxDm8CmrxSanUpybib6BFbP6PIysrLh3SvU7SizIOWWlxjF+az2HPBxxi
NCF2ePjz1WHiNjb+nZDYB223fF7vUm3am7llQtKeI9o/I7kUxYqaJbZj7adG9gzR
wocGDyP1nDcNUsVVVNx8qQNbiyyPkf15DU+RaZBruEEuYEuvq0A9XYmbvnp626h9
7KZH4ZaVLk/uekl072wqavB4DAT0OSCQ5s4fWTBB23g3k3crSz/zQSN8fCdl7ItO
RJdneJoIE00fF0/lZ5PJd70+44FRLbnF1s1nv+f5riJiCaPwJLD/c+HGsLv0yt0S
LrIUXT8Rb8e2dRjAWFpg7FVlby3+dRqAlWLAB3cD79Q7A9s87CIXutA7mnOzPx4F
wzU9ewDyCZXFQ3c5fpM52KBIJKQ6a6GR7KuVQ3NVllisWiXWgNXwcdzm9tS8wAAX
Spdn66WtEEboPD3g1oL7Pk0jGquG0pUXkV1EIydmH4jtDo3a22cmBbIrv+M5UjWt
NkwS2R+kQI6CGwqqLY/TENk1hj0yWw7ivrWrE45cT31XGvfnWl5x2L/Lefm9ELSm
oDdkKTqwpyXLP15XqaVOP/nwJQVTYYOtqL1VfNP8bWO1jAv5TOLSaFlB8jedmVSw
m6YNtatFo7dJ7Cf57LjAM+1NtvFz4f+56g2JAFG+3yfrXRFF9b8SQ1n7geFEcyYO
2NWp/zszJa4nyIb0x2gv9Knrf5ZIGivLs/9RFicfRG2iSYByvaP7FHnqnRwmpZ/I
fOX8VLGWZDWZWx3CEAGx7JNLsnOmm+ota7iC8c+2LVHRdwH4nHlphcC4oRisbfCp
APlbUp6SjeCmWNXYzBTkBmyha0oy8PnOn8MO11S33sz3QQgMy+jS40PeC05hYtMH
Ch6noVxCPrx92JQHMVZ5eLf3QQCuDHc9N6+vuNvck7CZhj+WG60QqL69aXRfaJ0y
9TD3Ekj6EfozIV3g1y8rrvVq8UIoS1Be8LxpP75it9w1h92I4Jatb2fOHf5Y/bE4
xw0ZTp/D4FIOTHvMjJ61oOg3qUyC14Iwwcd9oddd6kSzH0gcgcIc5JizVtocSGyu
/kzqyQAhooP2Z55JYGg+Ijr0fDVGsCylLIqa1eUxUiCq35HVpp/XYcMhtO1wYVnf
vYJeXTMcgaBP9r6QHJpKPpGRooOI2XRUYTgQ9tg6CUIQ2zzjIGTGc1O5P4KeCllm
i9mI1PpUCyzLLlyW7o3FGlqt6F5ouoWG7vWAbO0uc39Q3zDJGcMYxOmaVaXS6FoN
yOQh9i0oxxaDYaSVC17RT1VpLZ3U4LSGCqPB0UWUVgMSf30wm7wFoxG4pxrMsLMi
w/s/EisqvNdwgXc8NZoKPE595d34nBZJGvs/SzStbVYmIl3tbwP9TUzC2h7J3R62
QCB0aBEWuKgRilhrNRoNLdSIqelJq0/ptgduRZNxXHWU+8mCbna0gLG0yjtUyGPB
rhDGY6g0VPy4d1R9os6L/vjawcXWU67s5UyAbLjO7VkcJ1IUo7VhXk3XwLAzKNia
6lCDK1Uec4EH/LQ1k+kBQ/J8TlQ2goOVXZkf75K9PHSpZ3IbcUEA+u0BYsQH2gw/
JDEhEfpcNgzFeq0HYYaqz4JEd5F5E2jfmHVFh/P4CgVeEQsYFXrZqVVaS+VJUHCh
3c6hKC+vRl7evRaE7407KAOOsuY3+D73EcvztwFIDFKPTVkLYxFPPxncZT0PHV23
jYlc3LCSCwGx2F348gBRSLlfSuT9XL4Nwi26AeyG6iy3E7WThhJDXBGsj6O2qb1H
cuN7gAfqqdINLOYLWRRjBepdvUY9XG+OkubWAtFMZbDf+TfBsv0M8EwMLe7d1l/A
5VMittMU5/IoYGsfFvEjHaRSJWH7icyH6z/sq657O9G+mRyr4PaSU7FI4WA1VSIQ
mYUDofxsCHgeN+2E07GMEx373ESju22I6fyyF14De7F+KoxXIFiFxxfZ1uwG4FEn
0oo7FyR/6Bb/9KxhGoWP3Hat4rmsjd6xcWrRmmqX7GxpzxIjtTay6Icw8tiJLQs+
/xTRzHhHY8l1mTZxSVBlJOlT0NWjCdGt9kas91BViDFu+UwRiBTXb8ui+O44bV5+
pG1YfvN/LwQ69GN8r/AwwGBC02gE/5+TlQGELAWw4SP6wWc6MVt+m4/j50eg+4bG
NuiNqqxwYAq9V90MdCEwKvIWBcUyZL/xUIpT1vNPmTw2sFKTDC1QDUSNhQzcqzG+
iqfan7mMitKFqoD65ZVXzCnQPVDjBpDgmjao5QTnSQGy5lsMw/rn8OxSmSCX//2G
DCVdPUPY6t/PA6CnfITHxDF/X7BrWvIvBmP6lx2v5xfijDE+97E+FNtA8K2ISZIa
Sb2q1oS27/7UbcVr2lNkgpVRhJImHmZSvZcwldUed/SWajU8YY5SVSesZ6ZVwsZB
peadKqvAyE/ofuc1j+Sll56oD4yiFpDvyH5eG3QvsAQsQihIxDWK7orksoMcXhHr
YYw0VZYPOjvkSWzZfL5YdxYW+Mjlppodhtbai9KeC0ef/YwXHAbMhOi96/O1+i2H
Asr7N8PsHszfozfMfJuARBgduPAVLqNSYYeQ3hdgRQ6pwkEUKGhQCtGU+woYDhTP
NPVHtLCWVoV/nBaC2kTr4Mlqc690aIPplylitycB9y51R7C9itpTMVVhux+Sm4YY
O2QZ4ib7IuZukk7cMpnY+oHP7SArzTi/HLBSvmtTVOhK/n/vxlriiv0lMHkfxhw6
vgb8aZy3Ic5cy5JVx9yxSiCwU+3eCc0cjs2rlrvRGVLCT6VYMycDbIYCPcAUe4ZA
VmdZ+kAP3lfxxwEKnAvDxCCiWdOMumutXfitw0liGQ2sRpFqG2ioLEY3ODwiuV6n
oGB2TAlewwQobMwq8+sZaQxoM+R0eTL6u6nPjojUq5SSwD3Jwvs+ZMfkq429R3nB
+3WDPLOBT7Jd24sTEVO58FKGM4odApahzPiR109DSXems3e2nWHdDBIS5C1AUMG7
g903iREmUV+E9HWZcdMpv6hzPcWWS6GjHSywq+N1NUkZ5hYabwfHHigMQEmr8hDo
S0I2ZeXQPeK4N4Nm14xY9sCryeQI+1r7zvuaBzIcQSo51LEBq4sua6qKoUkeah+j
fCFFMo/n7pb9KpzXfl6lPxvUpZiOQHQ5aTeGa5WxY5Xrz3vHELiQMQRDQUsxE757
OtDL1XLEFL2PKzi54lvKYxSfAl5zsByrrlE1Tlp4MFC8YLDqaiKWrbhSpA5xHwo7
ycPs1RYtOuK4SwnT/soViZy/LrHtpydhhXfyU0H3tPL/C5VxGDw7PnulTgDL9xs2
WLNhJTTelqd0+bFloZGRdBEAdyh+uHenEMVW7S0vsKiP7wUM8J3lAq4FDzUxa8FS
ny8/sAtt924jm5g5Vf9nZepWJAWo6HG+d4rXUjIOAi6W7HqZNLqbx0WFamOQThxD
tnLXjZT0LrDt+oj1x7a7A9uG/Kz4l9zwn9dD2xqmQ0nedKE/3F9JrbP6eBh99qZ1
ofoD8Cr4maLFFgECx76GL9PRdqKi9642maP1FDSc9KIwV1HCtydl20eFZJ8CUhQz
rclHBvt5V7zDOpDhulPh1qj6ruf80mD+O7A09bhIE1FJOBcZoyX918CigviJsBIF
pF3czsORkyaqx1vFZBqaPkCfdUIxFrlDzCz3rKn3FcYJ0IKThK+HrvgXRzxPiOsf
j7n+NS4JaKNGUGBwI6LTQSGkntWnJejAzXFH8rE6pWmMG8sW9q+kCNDm/mRPF477
/+jnrBdjRBrspD4poZzQZH9Z/xwUx45z89MXV4kLyCP88WVxR/CgbVjq1d/aJxXR
/WIpbPEXjvUWsT5drOSajEESCpoX9N3I4g+QBDr57ksExoA7GaGYDy6gh6RqiA9X
yojOe0v/adjD5KmrAIJB7ynLFpiQQgg87Tt8zo4xVbCh8CwhnpEhBYe2w10UEBgg
zvzerl1/grZ2EdsxQsklcDRLt/9rIeRiEed1t4/PzWHzLEfbjOEPLrhiXjFYVFWx
LzJ0RrZRQ7kzI8Lrsln+9v3f+AqB+2spiPdDIySbOevoC/IZW0+7rYiZ4Y3zgiIE
baJTzsOb+jif6d+HP0uNBjdmnvqht/FPharwQWxW511Zr+lkU9RjESHC969C3GqV
JPZmIG1SslYnnrEs7mrgBeagnA9l+3piTN5op3uN4C5CeBWU+urdN2YXhY1+oYpU
+skWr2jZadUM+0667cUyWOfHyAzZgQwcHJN4ax5kRXOzKMa7i/htoCyaE11I2iLt
FkpcX0WNF46PU7wFAZvqMZS86cVv55VTuaUgtl3m68lVBsEGp7A94XlhDRq96Kzs
oTOlLVOhIGMfpgkJTN9V2DR/c9i8sxMVrgfgrqPPD73tnNFqxVm2crswLuwyeuTm
hAP9Zb5ryXXwTsLPIsuEwjFRuZl1OZMNJ4mGuA576BuUEwD4eIQvwB9aQvxJ8zyK
Cl9BitEM2mTfoQV7kYuXH7Sed2l6ZdD1P33l73YfITnUD2JvEQcRuCZz+7e1//w3
ctV9QmfQs8X4lB1IOf3pIo+qTQwZtNm7Frn+M+xBcl30T8uW0x+RTRdfNl25jZG/
0RTBufzQs2xfArNPsHkFKL91WEyLgsob+dJZaS0q0ciL10HHYr677fYAo3LkpyQx
QRnS5L+qBiEq2XPpcmudmju3jpHEfchpKU2Lon1mW5d8PA4Uqly3/iMVX6chVI8Q
v7mGAFkd1jmkYHZihTq89X4HabWpFl2v9aIgXTfEEmZo5y/GtToc+swrRjWIJquK
TE44UVn/1lO7pLKpIg3PZM9WbUa/C4OHaDPNeN/xj7A6mSzf6qiFIbSYWcYrg44X
ifNLnJn4u2YQ4kq4/d0pZQvQlaiTnqutW2mmg9I/aZwe4HsoxmB1qwZrmebZm92y
olVfvOX8e2WTua2YF8jaPaux7okQNgt/TAfQfz2rAonjv9U/SueeRcER1AebZ6Oc
ADraidJ2ydqEsgvVxng5ERS5HodTVhNzQBkRSN/PAdi/Ww3lEczlDdJ9dpGR8zpX
riCdwk6mqGgWshJRmIfTWMHOLO9QGyxTSaGSQN1n1dGrVoMAKvHbjvexeXaICtlt
5fonUt2c31uM0mJ8t3e5NA0ZLkSmS5ccBTJmyFPAwe9okWhOxKWsv/HzrkYwYqHx
ZkPQvhkP7vty0nZ4frgTMw8hQ292Ytvl+BEz5Rw8788yhdprEpgSmvotnjvgxpel
fiEifEOuRTvEci60VzgiCJAHKD8lGOBcVPJMoDiimrLrABVQWAq0GLbtvjpagl1u
2OnGRpePn6a0F+p/A1Qyk7zI4dVq18qmp27XKRfqG1guXUWutFprJiFx2XPk8PMN
i8kApzQpTBVlOot0dtls0R+XrxWVOI3WRqkzFuVaOc1Rtb4sT1e/Olk3UDfF8+6u
karcRXolQWUKHLawrAjYt22qeBPGHwYuQ05yxohKM9tTiEdbHEpMiitUpHUggeMx
VlvyYo+xLCT9DE5f+Yk+t7zXYhXo3sByyZF1wpDZ7nVPurxnIYMym9CzDT+97W1t
Gvjo64qV8D4mgxa5qxdZU/Fqf8uVQKcXQI8dIN3FlE/C/n+UVQliIynj7a0hgsW1
2Lo6yQwM9Jc5M0KnryBdyjEEYDAOB3Pivom1HdznEeFav4sqtQZsTMX8F4K0bJSb
56KcnVwM1wP91OjgHiHr0w2x/8aVsjl1Hiv3DOIdblS5TUN+G6PVMYEvp1mcS3Ij
PNDPuFc2pIYij3iLJlk7dzGXOzsCmMmt3rO4gclqMkHsUwlBcc/tSmsKKgh26jKY
TNzA4hpmIK4xKwEhvRKQ3xh4mPBue6TZ0qZ9ZmoolX0du0YGgsIPcTLjmY7sngFo
Znal/INUlGslCAlaMeBMPCE5rupJf7JSkISvMQmaAIt3MfM+ux1WTSeQaXpgLus+
QGg0fjGRi21kTqkSIsq5xYws/qVXbDoo3PuOU7Dm4qDsgjKHq3hh8GHh/bJwr0Ki
CXrb7jlRtDI366Ejz6hF6yaeU65LoGOaFzwUYcyiv7FOy8bOKO7rjK0TVcAukY44
rdGVq6Yk1UQcgp/6//LEYrC3B5JlAvd/xxa5r1o/zjI2Jj7Ebwt4d/rRn67SnbEU
1uEOtME6qW3NYAjwSXnu2XpetpLZ27u+us/h2DiBSimvIVx0AdUOc4mO9KAsNpOu
o0nYOBZei+Ow2rAN/D+6BX6uZAzsnCrBBG8DYFidPSkdI/3lwxzKEEUkOmDzAkMl
2lHnRpSg6uCQXCc8N2Yq4oxd0Xktyg8BVWTKq7WHgH0QyOo+AJfM8rAUsisju5rD
Tgj7EiYMYquiOWMUcr8aRSNc1c/3UXWLraVseQb+h+gzL2QMCv8chck2/t+HXJkW
OMQf2To6uvIxRPb9oZvSn7DwRVrr7UKf7QPjCwuzJX/kGDAyMMAgnD05accFOli7
ZkjfQtiyx6CcKLdjUg63wWSNgPk2deJyNef97fetwxKQxyr9UvlcKzUexgS/RTIs
lYUXO6/XlP4BwATHheP2JDVv14LNgIaROG6/tD7t0H2e/Vhs/nJzmCyUv3h+L588
kkcSISJw+cg6aMdrZLtB7BxmbSSABBDTKCuLviU19vjxXgWcF41eccgx4IPsbEl8
qzjTi7Y7oeg2ZSso9NvScClg0om/ld+F5y5QqCKbYHc/P8I4+tdIg2NCSufWawgl
wHrMGWrpkzBy2pIk/XUxrVq2RK8XNXB+cSpgFHZi8JHvUdOPw0ObImtK5DV/ambs
T0IhNebUDW8/73xh3zRJZJmEDI0aW8TyrqPfLql4vBiqXHMcKotTz9RAA3GqaMLh
/ilPloRwc3WG5fb2mybMIyGiH/xVgA88jFv6KerlsEFJ2kAjoxhd/oI6gm+4yI5P
rm+MoMUncgYWd3jWA8zFHUMWmZY/b6/dkOCBsWbqS7uUP1kNJxPHqxbhQpm61xHC
v4p+noi+ZV6cl1qYCobyuBsfQZnUD9oLri/pW6F3SuZyWaqQjulNzU5fPT2F0Cnr
1vRSHtlOUuyGu+BRXs/rn7gU7y/f/AS5RIYHcH3f+SxDmY7z2pullQTt1iH9lLff
pb8VW9Nep7bW4rJ0oU8o80DcYIWjwRA7v1hn3xBHXHhFyPaxNWLVpU0AR2DOx6LY
0OwrpULgU9C4FvR4iYkeHvgEDKWBdwgA/RsoxmiOJglfQItz1Zp2551isyQ2yo9M
6hCE+TpK76PydfOkSAnYxov92xQp+QBl/RUR5OuNe1c1LYqQSFtfZ94JitRfvMGN
lhK9BR9EH2Il1kNiH/koAPlu9uGBBa3BTFYUtYr8BwJPOtpj0ZijG844icPr/S6D
N6d3KGX0FpyGepPzQwF6657+YjwsTDUVVvRIqVXPrS63UquBSlOXJ3zfB85G53Q1
5L6acmFdHgIy7HMxsdbM6qYVR2nd66crUzx0so+g587nBMkUI7zBSy5SCdAEb3y2
QL8uSOULVOnkw4we6XGMj8e+xevnOF6IWEtxRpyvkRD904hrDl0j9mh+RSGM1YJB
WMz3k6y73GQBomIjfbmVpytHMWy0xSXmDmR+R+OSptgyficrdY5ouaaYdMTmhvUd
5LGXRT6hQtpTEDmeyP5pjL/0Glm/gXCYKugPRRAmM1UIIH8LeluarPWmekBbgFVD
TKhj2Lo+EcuMVS/QvuJvyYSnMV0J9p4SXVnMyGW2Hy41dflGPxaGsi9g7jhF6Rjd
BKDshJnrSSNACQWbD5vCANpt41cwZzQJlT6YBt9cz5gGgnLBMJXeWVGagvT6kjWu
Qiqsuj9HSdyuwT+z+RleFvcJbFAu/RhNCywmAm9u9+ywU09g9BoxYyjlkhtDdAXl
aqNmf9xiQGJCd8iW/1eHlxgN455eS5aBJpQMnwTf9pdYNM2mU3lC1wFT6fFZogFw
D2xC9XAbOg6FUysBuk5kX1m0wS6DUZ5PASDgtX6bKya0sRK7VFRN/Kape3zHMZzh
6W1Rw8G+QUR6D9McZm0FA1J4o4rIaDahIERSUJ3MQsGggHFjdFldRHk5MKctzUyc
7G4wYLYCBBWjrHrAoT92v68rIoS/Sf88UrQJGGhjmwH0VTnAIEdeKpVD9Xb5/+wF
9Z/i4L06ejHJqPVgvGDrP1jHWpiICM1YFk3YIGIjinX8xad3E6j9PcHPSfsuebOi
CoSOI4g+w7EOiNwy+uVEgz7LBd0eFgUOY0AsQr4/pMrLYVlA4YjqAuIZCWJaNjmx
wqj2Xr3PW1fqhS7gg076h9PgHm9TQOr75AfymL2YZxy5wu4GXb5UeDXbM1VoPCc9
OHlKhUP94w9ulidkGd+z2vkNoP5xqFoZI0fO8grcJN1h+G9KUhTYKcpprI3XTWU0
wfskt/BU94zSoiJcjLgkMbEoXFamGPwOa8qSHQgbNOeWCHYr5u4BGhtbrYKv8qXN
XBFUgkgWwYfRAm+4HSnNue+rzcBIcWe4tGqB9lfx7ZCsS8Y94hZSFvZi/SUMLr0b
HicxX9FT5xn4N6XZ/LyZeFLbdNhO0npcI71UKQClKtzHf31LClYN5IOza+1UleSZ
LzwCPEntXln9XmINC79pXP+7224eaK0TT5CanWdQs1nYnBBSBe0sX24XAHc0uur2
qKFSoh+4r1Vide/Z6HIj9H9QJ49h9dpxvVn+LstJH0cmX+gOBhIfkQ2dCowywpeG
jNDKoGFcRGOoEouV6RJjEja5IRphF5bz6JlokvQwR8Jlp5jFNotvdsH0C+aVdOI3
lAPp/BSwOOsNX+IVvMogRPzhvEPexSDBUYHmhwDDy7mzI6E1ZsLEHZ1ooS3oKPCt
EwW4/J3BqWBqR9sIlFhd+74ZxA4ihpZWb4IYNQn3xdQsK/leuqfhLhhDB31TkVx5
qiF9wHfi7/gapkLtgQpDTXPRNj0JhFnxig8ClA+jJSu8r0cxIJTaKDlwtVoYAZqc
gNS+4gbj+Ej4P0TgeD/A7VrBnXoPzBf12NI7STSOwTrSGM67x6XzOEVEqf4cIwU3
Vxy6yZ+x3goHsntuMgt+f97UkjdT8BKYpIVb3eGyJiUh6sdboOOQoZvDgnyyFDQC
QN13fXy2EWEMmjYatPWVA5YSEY9mKfOzXbyceoh99Y8xNKOBwZjZs4EwQLJuuuS6
b3LyiwQvEFoa6UFMKrBnBCefJg8Rf+tUNSvNiCtKLa5e0hlmE4XBSvp3ZByxhptD
vT03n16603EQyia+eFGk4ii+9QCJCSZctORARAKNRxYyjz/NwElKmhR+93DwaOIY
13aOjI0xcvAB2uolJYQgSXuiZQgOOlQ+xDrStyqjPupXs1G2K2CoV4P4nwu3hON7
DOLlGhO1/tg6W+VTnTWfAAMMrD9WdHGklqp4m5/c7I3042Hu09ART0LkKrfVBNTE
foX1duRV/Rv+NTiKfV+xdHJLpMazzQgzZuuXpRwn/XJqpYxkvGBV/NWXDjQ1e6fr
6SV8R9cUJHrIYIPabcoXZQ9KKWNXcc8PBkL/2oumQuaYfLsV6ULoarFd34k4ergD
qK8qhdYKpVr4PKhppDXfLaUFy3VGCITBgzwJmAKNTqziqOmydTbBTrLZNrEdTA7V
cGi/AAch2G3/R7hLJQ6BxIhtITDPDtrf8TdgXf8PupJAiTK6jR52Q2mcExzlFrEK
BNe30JK/G5vNEUarj53Nr4a5yMdIm96Tp6AJYtcHLJbsaSoINB8aGqsZHa79NEOD
pZB0d3F/zsGVccBQa0KdKOE/kfThGFfvQO5L1d6gWNRXGJbr/fWu7PdcG2jbGxNt
+DUWAS+DLoZtpKB32ztRGeODXlK2j3cDC//XuoT71EE+WzH5KD8+m2BrjQSchhJj
GvUPxBpsE3UYki/hMQF5FV2xqX1GBE2VcRyB0yrvU4aWS4uDWMh5gfBBrZnDgPxH
24Mfnmx128T1dSmqwFg+pVYogADMm1YBEsjwVIagKh5myMDcChh1p/3vcsc3epyg
v/4PfFfse82XdbUSjcr4ReU9lfl3vL/cRbUJ2ErdfABfBoKDH0SozTLTPoIayqTO
OP3NIJYWI14eu5saKPdnIWuKymYU+YHNZxEjmYF6+05rolf5JJ+cY4zSoRkrbroW
L3WDuHux9cbh99ME73eIvfNXlKfYY842tZtxCAkq55xCoWkbzHr9fd6TxPdkBNoi
fTD14PWWvLZ/oTknDjSK8is3tNiyh+TFqVJxyxUg7sO8ABdI2UNQYKW6p9gPzpl4
JuNtyX5eh1m2ICq/COSGehqLFpjmd/RoE/vZ/xqRT0wqarDIXMlrGH8sT0+KPiRQ
Oo9IIE0sMqvVBpYRJVjhFX1xT+hSAbdP/n7ep+b0bK9j9g6WeoCeKS52Qv5ikBmG
Z/Gj75qEc76+fx0wVVaj5iRK5H4cA4Tz/Njcsrg6diRhQxzljIis5ljzCak2TzFw
i556FX06bn6yttjqDjXEFiAyfwlI8HzSBrK1st/0424CqU0c2G3EcCGqbYtHJcgj
cED15oMGJC3kAi2yl5DZhDvvOVAhkThT67vhOlzyxzLKqoQBFVAqPVdOeIQ4RZ17
8QbxCBBb8Nk6IEqlyvzmX5XF0q+ltaG3lEhDBLAM96bQS5j4scTSdcMhUNqfKtXF
juTZYodCNMAiBslwYc7RhkoLXhn/CMV9s5saXIyJyx7J8cudTocCcaVGCMDla1Fu
Avp5yhbNJjxGqliq/JpPDE5qCeQ57b13lULI52gDl76lmseTzHnyXxPz+JnjHqgS
sZj/n5XuEkPOEgzsFFe9QO+tPeh9OmGJswAKATYYEZmtAYlNqaLZnpMwQzMuQbrI
X9iTI1GSVxDgccrdAAkLVaR02M3JhOceKBAmKgyKviftEQ6gNx4F8StTKs6RUpQ7
hMLqLumqn+WeSKEPBKEWjxucb0z66Z94lRJ68xMImgMPj4tLNCAhRpWp/nYz8bce
KRDY8TFhOt3bXNfSBrIstqX+JX5NkXnfKvD0aeDPdwZa/Zdr5MojEhb0nqxDKVOW
J5IHuqsB5F1R/RSPSBppS76Z0hjzZwJLLIYn6l0EVTnPSYHmZQatfjjC2fGKGPxQ
KBJ5NoOxeKfauCkHw01HFNI8PmgImmzFYhU9ZJ0s6sSVa1IYqYw0J3V0t+1kyOyv
mppaZfJItS5e32GgU48v0kfUyjaU1HHrdbPh2Z+LRSYDvzuNioO5c75hxNLbNTGn
R/ulbXuwVn3lAYln38P8FLcUph6myJpkTMmi+NvKQO+Htrzf28A4/UAEt29Oz7Pb
BR58xAXIaYn++Agx+W2gYZpRwPWNoG6YbVEMQq1vF/tFaTCntSBt6xjRHeO4Dmb+
Q4kdZtvDSyD0KqkX+Dt+leHpYMxX3T4kv1MTxMI3YlqnAo0oqq+TnFwZj7iRiOtp
YVUw3WXWMH+H/Olllidm3mJDqoF9dAaME/K7MqQvnDQcpEqcR+LfEnIl7cmUstXJ
2nYN1rU8XZnsJ0orB4aT+cck7rtiQ2fvnp+6tIsdAVSS0N8w/g3UcIpTI6+L2Re8
KfAg8htIb3YHT9cpigxNJB0QUQNhf7n0lv2ELzian9SdgEXU5gU4K+NeLz/prJzL
G5j8RJN939uxWxc/UQZVnCsM1gvNN/EWWesmXDygOC/zAdtWxemmFtjbK5//TZt5
WkzNilhy54PWQaw2VQDr8LjD5RVDn1yIL0DxIFhLiJcVznuH6p2SOBQjotVsDbre
MFjObFLxKPi/x5OoqbP4M/S8bavEtmA3j5VT22utaM2tuKrtaj41tyzcQR5WQWs3
JZwXnnmV+3vpMUL6EssBv9OaBpQjRAy2iZCkUmWBBsyaFHbfP7eeWTzaIqZq4WSi
+ppnCThEoYsuCF+eVmAJUcy1bK0WABhsrd++7OPl2YLeq+Bat5NeRIAKOCrtb2O0
hBW4UNcEBr7hFfuXQ7/09M6uw+7DqSKLcFlSM94n2JkK6T8FIWpGqpxfm0Ns6MHT
7spmZ4QKAMayzDKvPLy/FnJsp32cP7RvR7iMcIQrHG2u3/J7WJsWfMDG1ui3I1Fq
XQEfUQ0u2DFWAp21LB3Zq1mhXtN7sfi+JMIPnONZdLGk9Aj0wb73ahEXRwg43lU7
u2ddL4nWleVvnJqo0t55hRrS0rudM3t50VpGjjQETf52EP0g3GXkybVPO4KC8o4k
WKgtI8BJyvcbmSfjOeFb9xqPlPZE9abkA+KcyLDxUH4HRF7u5a6mc99tGip3Q6RO
YK7MmRVf8qnVjFJDtqkp59fIBLVya5zKH+vgrT82EK0lQXTAIz5eBIIUqeCQFPkA
GfpGt9zC4GUjR7d8uG0cG7x+PbdGVzmJz1/g1lg6J397YXJOhaI+waujdS3iOFQo
9Cw0QyKQaVBxcNeIRGSOQiHX2dPApzNjAk0GdZ6iGfvVxgMOgdKsa81DF09Ew9iF
WNk1saZ1xgNe1KZrEm0/31QDfWRNmL0vrOKzhOunnm1nJLwTxa1Qf7CMbSFXhtuU
C/CTHUvHc0fj/OHOmUEkr4Xw/PHdM9wG+0m9xLvZWLGJ9vwARLujuTO0UD6BL2Mh
kJaBYduv7OX/v3/Suf1m5Q2qATr/o6paj8N2u1sGyXU1ud8a9dpZ/if7XpFgP9aY
ACRG8Yy6a+GMAzpMUP5wUfFH1vhtX8YmSL7oR/S9bj5SUAbuoUGMp+OUaDYkohW5
rPNmHrDYZVm8PE/KWopxHJnInidZK6LAVo3j1UcF86NjiJVGqDKri9jJPqiELlUr
nm/2v+4TyrfcMr2m8UPJ1O8ceLtLIZktue9rz6AAWMQgLpzSPaVDvtwMeFyqAshD
0dRKnYKboOC8t5zf8ijm2HGa7uDD5uzDDWeluy7fOreHkiAGhEDXr14f7MZesw8r
q2Dv9z+25kp8LWHbI54e1825FZ7Pk8N7An0JOquTPExFDvu+yxQQIArtAM8nxXrz
n3nGZ3W19H4dZOswY50fcP37iqo3yBFkAn1qSTyMRXLmpn7m03UOSdXeafdRuNZQ
Z0DnLrQAjxUgbLl+s45wz3a+rJJ/2yJDPGyGBQrSNYg9/pUGbqroAvRSC03qS5fx
DeSQHYzP9TbEj4tKQEH3PaJL/S4pqaXKasAwujpn5ezGtf1GElevSH/Lvdpzft7Z
xB6ee9AkGE27tIcg/6kfmeBu7jLd2Mgw3yP+Y6BznSSM51+u3ykspyF2sUTWWH9w
dm/UxK+b5hQ0tydlmM4Aug9KwS3ZzS//2/HHfgHv+MLS8BtfmS0bAH/So/AGIFY4
hgRLwxVbAB1kkR20n8kf/YIbrlbISsxns0I5GB7hggm7gOw4zjCsMa/iTOv+7KMa
Wc/mJoFjgi3HLVzjCsyNRSFOuCZI8DDXim6Qw7YDuJG3gpMrvozW9XdIyRQbTBnS
EJfpwFzdSYglBiNhxHDQwQeY6Podu/vE9VyfiTLnPB1qwEQBTSdT2gCxmkWDdxI9
xEYauCHwwYkAKmACTNCuRiWXBd62jzHh+Sa1tC+qhedE+v/wMyMJQtmH7UHdOpF1
S9SFQsba1Kazr0xcs65bV14zrprYaFpP/XwDg6PYq3rySQvNgHvL/Ec0oGlXWWx7
q1eeKupetd4lBh0fjQUrkv6NZ+q6mqtnmI4Yvsbdrcc+NDbXsnZajZD2vTRSWR3Q
9SHCbPq4/PhKBgZj1a4KFfthRnLODawnZz0L48TSROc3TPFZGexb5CBJ3IO3vLuZ
TFrv7IRMBvLv4aEDYEdL67/F9VhTDVptRCmg9ubtKoSz3Oo5D0V5pF8ADTcJK4g9
+lTKd1kse6Hluhtblw79jcgYW1E0IUMu3c5VKl0ckTl2iFeV5Q4nheqcDK9U+1YN
01A2zWEjxYbIHxWEgOa9n95fiCpYNfsOTXwgk2nrsvvN1c1CGMf8imAxauqnhs6P
Is0zyxtdeL+L3mtkx5GTWqF9LZGekgq4545jNGqtMrA5Zuuh58jkgkGOFECiUKt/
dXh2CmJyJl6kEcA6jJlO4Xk9ji/0AcJRDWJgshtw9XEfqEl3kEvBYMCb6n+RkbER
m2ZDgCmGznlqno3joIm/jaKcwmG+Ov1JUp6NLIFMfY9FjdWbvI+3nv0NtHPY3dJC
vDRKC75SGUEgGyA1zPwrbpue9CnqdS/kznBMpiYAUXvhdVVSAJ5h+4y4Y4xgRcO3
V6SFNRzRYXdvm3TYdZb/LwJ/uLbSxxfPYrMe3zX5j2cBO9EYebLQMYwjOMZurnjQ
ovIGbxaCTVDwi4XA+I5pf1fksE46kSBIpGAFZwG83fwgAbJpJNQu1OjuxCzttTNm
PmO1DzPMTUK8zFBk1h9fXc2MZTa5+OG8l0jfrARqDwCC3e7TB2Zaysc/dyIXsGGh
BDgbgEJNxwOdIKL4wHC/EB430JPWiaHJLCU5xOQUitWy5I8ijGezfIQHDX6Ds207
P+7ro8o/tLRbjtt1cVD+OCz/EpP3B1JoMmUhLHxarreUjIHT//vxH73CreMD3YcN
csJ9kJAmzVNGF+qZDGr/6/Moffz3tZO3dmqL9k3pjdCxmfPNt6uAMiQXsH2vea0A
Yj03WutQvjK9EsySJZ4qtUzk2ifFRvH4jG37RrYmyY4Erq24H0g5bEvFIUjVoMps
M8UzzKpbWQpXxv2sSmZ6+5emQcTu9YZZlBHzmI706VYl/fdxZz/K+UFME8QY9/pp
cHh5LGGuBRQiH1ykHpX/D0yh/bOgnYYHfuTASfmCoaJqL6VQmYXWRdGFYfWnOizO
GHKPqweDhFp26ki4Ph7iiGhOlTl8oW8yCcfzTMDZe9So7IPzV5NcdCs1g2CWgahm
ljcUHZxro1EDOGxRrVViy5IC/jCA9WyE1k15FmxatWcGHNm51cIpyYXd+vcYtHyh
mhvdjkjUbvvVgrTjzg4rt15u5PGc9BRn1b+qEMtO2TduGIgQ4t/lFknLlFoeLQKR
FXPDH8UkDihk0Jdi2Tx/esRSImXhUt3aDRiO3y24aZCXtLlkyGYpBU6BY0g3iLiE
0OJaehCyeltXqeyV2tn39LC37J+Tpr8rSeCnjM31HA49Ze8xA8InETdbzYkJwPXt
cD6XXYDeZjcvE4sb8dQTg50RtCAzq8oOZrumC/Yin9B3H+Kb/+4fH7Kmy/VbNax4
0NVrYKCc9ZMQmtNY3qLOBjXMfyDeaHuyRS9ib3ueMxtBdq5yksR4f6AzaCHc6Rk5
u8X6J2Nq8aof3R7qJ82PnMnYtOS/NAk+voxl7704CrNOira/1HDJ9XqEBden6YST
o/p/R501BcOLDeO3AkNAVOqv1H8UZVPCoWyN5yyki2rTwS0f12gfNfRVLGJPrsl0
q8SLeXN2PXypyeiGL42wSDDo9drgndoAYxAh6OqFKAt9+CDgmva0yHd2QIXd0ty+
SA6n7bO2eWlnBkdSGeDbuXdJijmqjvJokox5wDNPX3i7o3kll5rCm77e83PuHTQl
8GZ+ec3GQACLJz4PBA7z66R/KJu+9NW7+YajJKnWXxcAFoQS/+yYF66+ies5csie
uSqgw8fkhjJ3Z4R5fNboDy0ah1EvhflK2ArEaQka8RtM4DB/C6l1mYi1rSRdBJUG
7Nmd6BqiDXoxASMnVtujT1oCw7MZ2r7NmoPzhGRLp7k3cfRZkNpjd1Kdi3UbP3Pq
1DEC8peEQOpG0VqME7Jji7XdV/lKZIZo2eiP7QLprRJDj9KpsKXwMFTFhBsI3isQ
q2DOIKR8j+WliDdhwYqltIRAMMRy2MuVIvjd1sYua05P5lZH0N7DYBKQfqvowLXM
FONjTuzW35oVlkNTvJ5sbJgX8hIeKxtGf/sSJDHPkZ+jWFccisUuUehZ+nxnPcPG
3emaQbcSStSl0t2yX1sOt6bOmmoxsdIGdZQhX3i9O/J3ykqdlJc7JW1fmzXaHqMc
/xUIP4KgPqoC940O79ASTvazvJHL0vHScFTSPapIDpGcljVrmCbcPMFdi9Q84+lV
nQJSQJJ82BUfMHikYfDeawYTYntE9Hzd04lwsvV5GNd005LJ6mpCR03k0/3l+t1T
0LgaoeKNCJFXcAu5P8Rx7HfP/HvSKTf/oKzIK6zjp79PS83ssl+/2dAX3ItQJHLv
XA2IhaVdnwoO8k7BPt1Z+JS4Si2KnMC4bV9p1mJbEjDIWLkpR23kS56wRGZjAFLV
6T9ieJ7ib9aTF8GSJfx12towTy4+rTd6/yjS2fsMnDDVT6wcmXYbhyBx7GeudLpc
RyIWBgke8Bxnepq2ReCqhU84aJZIJuuDC1Pvy1YynBT4J+C/V4UyyJj4AulDsSSp
QQHpVUBkTOfUjd9WQoe6BYhryuvYbnWXeR3dssys59Xhfc6lftfToIhqRI+xH2k/
dLt+qI+D6i/zNf7+hAri8UYJdGE6nLGyGl4sVhsujyxO3YgzaekDhnwCA/df3f6w
bbJ9w58PSMl6Vy/2EWy2kFxxoWeFbn7LwSK5ezvYtFuioucCt6oogzPSF5m2McHS
F5HBGMqCf5M8o8yFz4lLE0M9qg0QofQN2dCqQDtARXY9/ivgkFMy4H3OkZw/k7Wr
P0URytWU+jUqQMX7BXXEi1wrQXD3FjV+nBZF7/8AJ9DRTSDPSIbBAZmPhhDftUxg
dFb6HOb3U6MuBitPk0lC6qj7iESS17wb6PqTf0sY4rXSPWOToVfezR5mWpexXEyC
jlXPRf6+dm1Kz14hiPGn4f/BAMwq8UJHq9xjroRfbjcC8cUKhGhrLUjeRXtpi81Y
J+U5ZjWk3sW2atY2X6E4y9seq2a4INphj/sGGN6sc3doq24UIM5m7dxDNnLVwLXf
lcmAIrU+RH+ilE3aZ1SGxzhJdM9yJFnzZU1O7VVfck8IFuSRdJlrgye02vkT9x9G
dQ4BEJqwE+6iKoNQwKUi0ix3gGudlTTDG3lGyHnKtmP6NFKewDfxzLTspedOzsSg
S0Y6a++wXZJXsFs/ZFsZofxX0yg1RK0GYkZ1GBDKPhBvSJvzJuBlVW1TiKpKXF0l
dINEf4wWGctMsg6Q+kRUG/86Qy3TlwK/2+9yBgXmnPkfy1M7Od3PhlaaXjknkQII
PNaiRsGAHu5qtuZ7r7tQLVgtWFimVS4nETmpYz4i210S3RyPOz6eXH2ICDLH1PQh
je+iaNdM1Zmath4P6vwXyVADs7/QmtZQgxbM3yUeohui8ha78QM4fOTV3lgTuW2l
GDOVshfMLz6t1wcE2he99hNh9fTJ9cgSPIXx3Cr+V6CAkavS0dqlLTWq4ydBUv0w
L4iHTnMkwfA9Pll3rAdWKNxBSWFkkWHE0HKtM5oHSp9+/+MQdjv2DpnpIIVPvko+
rLOI4v701uu/jIz2qbSResKQYYcBR4Qcg0JvQRUgBg9FLF6xjVq0EHr6/uRPd9bZ
nQ+mWIdMiUzr8Tp65Pa/pYCEyUwZzvqpvkkLLSACOkOiiUbNeUJqkuMRT0Pbo1Kd
BGQQH+3jKSzmS2c7xx1IYd8uSqId4R8cRq9GZTj/dRSjuEihp1wIA2pzuR1GiCTH
L67VR/bgwGlaKN057a2uWhNWT0bs9g6jPDR/eXSehObp7c8eZjX9kUodd2d4c0le
qquiHskjGFK+4/5oo4w+QBcpi0wd6eSg4GXzEju9Divaab6+YRuhL11eACu5Fep7
RIzGXGhG0ZSivkETn0u7ajaEeta18zBlQmARxFM1y3bBaHVtO9W/3HBY8LEGfbhm
WGRWZg/Khtfmj8pgcM+JS+8gDO9C0epYt94n4HtICbPgSQJotv87j16f4DoB960h
5ssfEv+exWL+NsIQ6ovkAAbZwKbM39Pf/Ko/PRBEYlUh/HtusEEGrMJtHNVbNz1p
RM3a8h4JQFCnQj3mL8dJtll6wIcryptObINYrYz3kEvX8kBzie0HiDx193M+2Bpn
gBK5ySJpEh4aRPrBZa8lM+ASeAm6oXr1y/WlfB7PcyGbvmhcRHrgaSey9KajYIA8
T0mg1QL9QLcgxTZqcL7zbafqjzcUVRNlPIEPr+ZYGR60qtHp5wiq4Jib/W+KK8sW
QMDHoZmaaRXGEBF1lXoyum6CRm3PqinpgWQtv12BXT78bNB0T399/lHkfTCdwxLL
cgqHXlmmKNV4CJxURBkVF6XInX0AUs4PuzEKYGV1vm6Mg+J5pVKeujXJHu48Nf6C
lEt9/U5xRaVYYSuKmGezPowCg5LMJMt3X10hnb4+iStWmAeXc3aYJ8sY8dmeqis3
BPkuYZ/Hvvv9MPsbyo5YRbDPOe1UG5nUD2iVbEpkJiFPtexLZulPXoIWqcBK/MHY
ynpG5LDtgmMQuIGpQL3ADSOFHHra2ZT8PLEa294+9kma2zQ5xQ9dniuORTBLlTUQ
XeItcojzqOzkoUrZybPf92SLYMoQ+fg5adgXuPiA6t2aYdwD3WZugbWlinJ/OiiI
2MY/8oB9GA9epRUnz5uf0+lZ6RvcQMxqG3i+9yPncTcc46163RGXuyCJXRgeQWi0
6gjhYssdrm5fwMRoDuCAdPvdwfF6D/ESzNGXHT0IWB+HZtUjqLDXxEAAkPBUeh//
8eBp3qv+mAJdjIXfqFIo0R4TljizBY+GiohblHKAKiK1ZpHUWP+qpOJG6j2JTVnR
9m6fnb+3xpR5avgC0BTMVAtHZlNsblH+tQCNDu0rJyfVodwP5UjU07TBiTLLAb9p
tUAi0EZPAYEv+EUBQ4w8+GC2xPwszMd7QLcmtE5Bc/y4qY4ARmD45ujFdtnA3orV
aMGbq1bb0GpcEa06Xgb9T26lvf0HcV/HayTViZV8cezIF2bLhhlciMpM3wkc3p+L
BJkkrU13gzblotfYO6QQaoHaCRVSydGKqhdCdz14zvh05C3fDQqYCYuSMsMLI8Ac
W0ljivquvf9cqcVqONwnDEuxWTjLYhV7rhbdA8VKbVZ50SpwJRLeY+QN9VL5VXq2
7ZRmYs1lfZEOhVcFGzuAEbgPmTZwU071P67t9g0NLDPNMR7JOsYiJWIgZnoB+l0u
jkwHY0kuiT9w6MznYaCBxIKo2Kty2mLAEJwULU2Av22uTht1ahp5miM+RWzBfL0p
obLWxFB+eX8KbbVeHPYsnhxe4HokdvReJr4BTHevHSdhshspLDWam05yR7geIX7G
FEkZjxcIaCBeR+0zGWjFASR/PboNFBdpKxSUo1NFIv5HtewmQCmJ10zxanYRK8kA
jGzUnb8wFuKuTDNlKuXosHKD+SA6rRSoJMp0tH2g9QxgFX7HdNvsCXR/i/baIkOV
5K62uTFAPAQ6tfPSV/AfaRr9KemgRkxr0VpiioBKnaGFjMJVdNd+puks3HhMD90i
OArajWEodor9wE7p1KOyFNTt5YH+xkLEMTAEvd3bZF+SRG0RpYi3NhOtXUNsLnJe
W1gEcBdBTvhKsfvxMMlvV7YbUk8tJCUvxUf/B7hNWrn25riZms8yelCk86nfOADa
KeYhnqJUZPG7rAQLVdngc+t3rYpYt24ZLlHlc+w0nRwywY7m2dt8Z2RcU0yxkDFd
Gu/yzI+nMTyulnvZOuMN77B13SUg4GRS5bpRdH46CGsiN+mlHdGGNSjynDjiznPC
nNolWRLzbOAPiIoTrrAvK9ZyTeSxikX387SdgRbnLJSOL2kpIiyM1B/L5vv7dDIx
vCA+Y71qPDH4twoN6JJBCL20Fgfu2MShQ1Y856bVlHxAGVZ/YJcMFShbcLRHoDNG
sitDSNaTtBZf2WoN6a+jidebg/xZYFoLz6HNk0BY3N1fHQnljKEnc7aZqG7w+c7G
p6DlvKmhGSjd8RP1mmLoXjhWlYXUjgUvnTo/PYETQMiPaKje4Rf+UsNityiYCXt1
qxcE3C3Z92vOSigUNb2PnlEPGbAq/9WN3HG2XlXBMbukK8f1hr+LaVMhQ1H6/n9U
b18IZtbKoluBUidb5sS8rWi+8Z3ZFULCP09pm9bd0ijt0J9m8DpPZXEE17Y14kVQ
gEloSWpNKzlsTlvym7keMqEiTCYosZaGfJk/nS/lrN6iZYuBf5aghQDY8BdStnV9
+98PFRue4IzePF2HNDALCixQ/99LHQWemXGVmONyDeEqhaaAdTAalIVOOGdYFniy
w1vmhl+3vx0+QOhGJ54WNCnh/IomFvNoQLax75WJ8WlgCG9IXYU0LoTHxqTXmazd
s+PhhCZymtq8xCgy12T4OK9ZL7TUkvAmZ/Sbzb0/QhGg5odNQWr6FnRZzIQZjJf6
CQroRXl6ULZ+ekwwy4lLb0CK/vjjr02FmutG5u5A/rf7G24JCe2isnNYkCVaCM91
4azCwdAfOH/gYYQ9IChdji9QjELxUzKvA6z3mVtVmRRhHHX+e4n55C1tinDPC/U6
LtQhyns4aqN9sS19VcSKY9jCWG4eZdqtPRxdIMIy2b4DM6vHUyz5EENUfZ54sseZ
kNQmZ31OTPHJB7C6n5v07oiOa1fZLYQS/auxIetP+kMZNv5iMHX+lCHMbs3AiWmZ
FRWSLzHjYRQl9oCKltrDFf/9lYcRrvBmcCGFXZh5c7xSutdTf9C9pNRiHdY39qAx
BjEy6D3JLifCSp4dB+0B+sqrouwZxojvMZPJ+xS5WFByH4WO1KwaNsqexM2TF/fM
rDAnmQgNPZ3yNtl6tMVSvdMlht2TMLs1G/wz5YeHi5IYozORAIc4mp6he3wkNmYi
SIUF5WjNPC3FPBapU/vuIr8fRPikboRjwvsBXD+VG3GCEcfkU41NaOgOENfgfDiV
bxRcRCWYumGk4k43Y29CWL7cOU6tCMF8vf0aj+a8ptjTmpZ4TAIdWN9MPGfyOnjT
WAz3w5RDXD6u4iRa2Xdla+UKdpLet+70U9xEHR9U2FJA9erVW+sgR07AoSXsjkKn
CzthOVHWGNhWBPbJ2NqGedsjVqyP+kVISmup3u36ylmAtoIgL633tdy39mJFcyk1
npakkjn+SEnp87UBjzF2uovXuDzQnlfVApg04H/N5JCrj4Y5kwuq2EYB0L98gK7C
vMOzS/G9i2rNY+STW3waJDYWcplp2SClcrryUmVkKA8USrEzzVmD/QEntS90LKaf
FhPgJDXjmbhqYS8sKqGCqQ5DZHPMVhSvLGhyLYAFcv0OUwF4JZcremhPtCQo3PXq
+j7D4LLIUbiPyEblXO4V3MnMtW2K6wPUhBdUlt3dTeinvMvIZSmKazsKc/WJPoeN
xKGipOSJ39SeRx5PI3yBYBCo0mcadL4M0X7LRwhn7MW0PFuT1lcNraG1wdXAiEv+
xWmLlLqSn0vljOBUVT82OtelOoeiTxOVanG0/2bRFYwL7qaB0WdgdESWjC0r+stz
qKY4JRmISw5G/MRO82IOIHCQAhwSDpGEYRcRYJ+laKqXc0ACBegLqbxLMqsRNsmu
lXoSEN8r5vzEi2I/c5uQ8aug4eLH7a5kuqP/R15PQeT/NibeEh3tgBOGxe2F1mE3
UZTPJPT7/Lbr1oiwmCk53kPPc9G5OOi9H/pt+ycodDqJd0hwZEmREty5U54iDlsN
pTYW0VUSD3nnkaV4hVYftxCzWKr564EEBUPr5a3eyeQXE4N6bCJy/RviUzR3Dp5e
XTaoheYcHLDB8Wq2duZxlSwQ9FiVrKsPIdfrbZy+Qofgpd47lW+Qq+y5NT7nyI9C
zp4zx3cQUASB2UfcbnXt8+uKSIwDpQRpaDEq1EvXXG5splI4mm0bRKEdyKWmJNAX
7ApAv5Ne/q74NXrCYYRUgZ0qwgdiKIoxkJ9YhDVBoNXyg6uqmoGOn+QUiouiwt+t
tn0chrLOVOJEUk6i1QC2yq3Nm1KVBxIk6lMe4AS16OWfDrhyHvHzymMhTZXhN9gL
+Wam52anC3hIRNN8b/ltzvGHj+/3lakXOE3NqDjpdHB8J1oZXIQUYFrcpeStQiDf
DnA/1+7RctIfPV10zeg4fRHcuJuLoFzL4TpdvnN4PyImh0pjcBHIlQ55BZm0th4C
hCedw5wosIIvGTBQl5SdZANY/TCTOyqXqi4TrX/Knv5HIF5DkjbXLcSoopKaziHV
mFXQOtAujwGRWKupehdQuz9QwI3OisqLY96MfCCv+Pz2lEt2fwp4YyRst2uuOQTp
PMZVocvzGt0AEaFSG40qAdNcUhe8sfZa4EUYZ2LLMUqi1RpraHjVUOuQAKHijUIE
UGtdcpeEwqD5biyvPaXXG720yjxwqrRTE3MJwZL5qByW/HpmuZySaRmYHRCwLZfi
p/WTQzuaVgO3HvFiH5qHoJVs+t7g+jHNUG7PnQKAghtyyXNE4GYgoWEBb+9Q46DR
ImjbnkIwYKkrqQcM14Z9NMq8eMANcnQTfMh8n9f1vbq4ETUEhEcWbi4OnjTqkoo/
FTy87O+Cg+S5cTAMlvggKYdwdnTcyLZYDbBIhGH5EZ4bitTSO0OKxk5Joha2+hD2
HANUDHG1UXPWLv9sm3JMOLBtPw2it5MnwQJD76SXFZOXN8lO9/Qwz1+vNHFyfcvH
kmWTAZ7fuF72K3kl36FQuEBHuEVRIZ8W6KPWgdcozfFtnbq351gjZQ3JDuZzdlnq
J1xxs2d+XqAMG5VhBgxohvSgy/8vG6FjWs0f7/Dbuikrzt2rHEhH294MaJumNHJQ
3ZYjKE/ShJVs5bbcgjHzAW50ac2a2sV+yC+VMeSQSmODx5AProu1YF6IDTLKg0rh
868aTc18nsNnfyvQ20h21tJsPNr0kCkQNUu87LgVRj2hKTu0/eDuHtVfcPmb+4TZ
8xhFBrD9KC2kmZuC0y22i6vvez8Ygo9ZAaeRv+3CrRUCkq68HX5fPEVSz9nA++CS
vVzhNzJwV7jUDZNqPizoHjgl01p27oO1DIo1FsmIBvfe6axkV9Z301kn8Pg5pKcl
ZuyX95dBILMrGNBSskQWnj+IZCt0tfp4q7qs6UMpg9tVgZMCoN8E/g7B7Qz/E9Ag
Gwom0FLFjtenkc49e2orHw+XryJ1gBdGNnlCZjP/ygLBvXcCtO61K7QrHv1CLRFZ
wRKOdD1AX/6bKxjXIsxi6uVrk+zztmfkIEwq5mKBpF6Ysz0I7+Gr97mgY5QH6W45
Q8hP205N5AIBRFD6Qkzd1qFKeeWhRKkmuFC6LzwY9Aadwqn8lVxy+PwSbSyVyMyE
cNyAF7X5JumO9I4StVWiGzERI9f2Jzv7Ga4SYuw9n6MsnFKE5MXhUbQLABuIhtLO
jgruSkHDMjK2cnTQOrZRzBHw1TVwUL74KWalISXKf6P9AxpcIct5b+LPwRasrOY3
IQTvbBXUxoXorZSyNUbS0wes8VbSuSIm14iftnNzr9FeFpih+H5t3h8UNtCyVuOm
MnW7pKTaquYuEAVX7zGXz0qnJJg2pVdYBRZI/FvZfw8nkHWLfFZpVYtFyCOT/F+h
y8G11RVbLTYZLmmyTnz42mzOeq8p91Fz0kB02PgrjdCfIpjDOZCYXqi+3WOmrejM
5d0Kzbqxuin81ty2dzvD4Z7Rmrz8qpCsXL45OY256+awVMDUicTvFiTGzeL68FPt
+QKHbTiSvJ0wb1di1T+L4SfTEyU/clerS8A16dyCGsJx0I7WBaUaSF3lKAYOKInO
epXGN9bYWXxciI9zG7kAKAcYC7bLgwgVhPEoij3KUJd8tjLDY57ajBswsEawxUeQ
A2B4ToXjQNItpwtO5QHJqB++RLbsLoG4GX70td4mdQO4U6j2FsY6lE+pPuyfi2XO
vqAB9isyCutpU2m7aj01KKQCFbALETKxiwlWRqmcWv62jEbuBy71POzPkgUuDRVW
bGxSKMVzPrbP9/92mvCS2MPlpvIzFrDNQ80BTIM/HcKaxiaI/gCfWyUwlxWkn9Gk
TDX2w1bxqqv6Zs4xy1NKHC0cek4FLTkktSNb/YqWYh/khmLs7CxJys6uYNuEJR3r
zvtLBWj/dznKDdxXYhsKHRt98PPQS+lcjpE9nmKejMpcU3SAr5+KtSDQWHVq32TI
ynjbotQoi5A4bq79sjEQl4Smb9FRL0EgwHp2syJgJIusJfwDMNaYd0/JG3bdc2JY
750eHGXQVOviwmEDpCofx98CdJklZqGXQ0iv+bVYrJ3dB8BUFVVzZTj2GJ3jrpmZ
edCRe2BvkeW+ClIDX4r63lVbaGbjboYWtrrCo/LIYjskznawm0Q0XmftlHaMQA09
M62QaAzdqhEpoum+6W2LAd8gYstvrMYX+LH1uxDifwtdU9hJR9Lj9bTGTnmTg6wO
BLf9ubtuTaNlq/G3yFIMOkkt3cul6rlo8Nk41Lp27NczkyM2vW5hgz4uHBiXa+Gw
v7Lo/9WS9jILv5H68zv0ExDKRoCDU3lDKHJWocHYTnNfGVw3lWskD2tWQ3vYC6Gy
wcxldx848c+HSpTSXFEGA4yOsv9AbASFuQkAvd/ATreLsf9jSYsB6TRrfpOzmEWv
WvmBSKrIJsxV6OPnIG1gbcx/cjWLSA01m/qvOg0mHS26rU35AG+t0ZSwyMAMIcK3
1/E6Ao4H47Gj68mNUt7Am3xRjzo01eOlP7eTX2rZY9TM1IJr5y77ReIu+ade4s+n
hQosDsCLg6DjgdVh/9CzFKQzKJDOBPwZDGDqTVgyU+Sa147+bzqApEAWig9kT5N5
ic1qaR/i/FLe0v3+cUiQow6ElfLkaIj29fTU7FdwDaEdN1ajcQh+33f5AoyRBGjh
2vOCe51yR9YC29gSCtmwY5qqNdXZij39qgRubG8zJ2oIsEOnTjnCxGVDHfpBT9yM
I+tlMlkOwRzr4DrYRzybDmvdi3mcOQZeInxgDzw0GeuG2mDXMLImi5lGh0FULCAa
jiTpwcZJjyZrkGMVYeSof3Ho+bD3nzg0Z2mmvgynNV5DZynf4t+BefnkpAw4zirV
FldwL5ofFTBvDkbWGIc2VLXugpDdzhDthzsvdMzvJKJRYYyLj4MD6pBRemMvDr1q
bcURI4x7tondzzcknKu3zEdA5Vbo659nCqL+XSujqIVkQyVL55j9yNJFDacz39a0
9liV9nZTGLAZVYxgyTYGlEndewP5vb7StyEXWV8rsIER6qPTYFJaa9SSQMc/Oh2t
ftMe6oQLIB4+u+2QR6oC+DULNp+jx9L9FmSH4WeINT2co+zvjRcD3C9Ij9qks1ci
2kEYfEN7EtpuL4YU8zYm8AMoF0TjQ5Xqqw359t/PFdJfljFpzzTewjjBNIQsJFIV
NAsA6mAqxoLYluX8anb3jUOAyvIvL3eA4IllszzKYPXWIpAeDoUPa6B8JEVUONmL
2MtmFlX4IcnZbpdPWcJXOTCe7szd9hq2zvbr0FyRfP7tMbVoihiUOQm6UREPQHMn
J1TOuNkhfr3bn40PNQx721xkDuvwgoNmN/JqH5Rn/dMFQXfZA+59xm+N2wwi5oIe
y62LslLZOhqgbs7YFgrFDmYIg2QK10zpl0HT7E+ypjDUxxTkmWlmNYaGu927WScK
XdO1lVDdndKaBDmx+RqaBcix91zY3nqCRSqFXj78DlEP0WIapqw37l04c5GPS/g1
DJEQNvtni7IlmlKKGKX/Jj9R0rMU58TcFYnKqouwimRZQrKcvWM6ONVnpmdX8Kwh
t8WygqROZLYWkX+gCDTLjve4f5BgAo6feNi7B5D4thx+Ekewgp3OJjNlc6ibNIkj
+ZmBjQyffqOd/sUcZ6n0jf8pZkmccL5iVZNXI34m9B7ER/l36MMqHvb/GiF9dGQ3
W9xqM/s7N/ylXe6Jo0Xsm2Rs/XRvZ5F5bZFTDMGxJVPcKzkOf8ino3DcH6ORld8A
1Qw0VRJQ1GwezSFJJb8YR6j94QML1+LrU8yihoPJAqnzovB3CV8MJCBAoUXgSc78
VQ9OLVR/ZhNo5qNwfcxX17SMB96fh/FObdJLVMy8kc3xBchCvG+MQLCU7WKhlWO7
ZsNrW0PR0ESUvEcz4uNr3bFNkljyrMIyhhsN2P4KyZpkkaXm3drXcqvXFRC9ONC0
J+rIzPoBIeptMPN/pft/tHOzV9Jg3FTkOlwqvcLsI5XngLq7JhuwhqOlilPFSw5Q
wiOve8uDRU0xUl32C830kSmQaanEc8rofJ1xi6d5mIQGQOAcoykdhWJEaqcm/7d7
NUk/fAOgMFjVtoVSr5fMDQDKcH4LpNlQIe6Oew8b7CytoOnnXx5iaLQj4ECsE4vJ
riE/3tPZKozLB3XzmK855GMYCqWKAct5EfCVSb0V9cIozm1cEYeHyvi13mMGPt/L
XtB8iNVbrDL+ECwAXsQ7LT6OsnjXjdB7y/TREJdFSA2J/fQAnpgHfuES19bu1ogx
VmVzHRZo+gtiu9McowzEcGK8J8DwoB13ARzhGXKtwL67tAz+7aNsmM3qW8SbMBez
eA29okicZhPDT0sjDRlTw+55qWhJsBmhgL6YVhXRozXqUs4MQHE2sGqru338FYcT
d+fGsopaotyzmrPKNwzHNizSWa2RfiYNghnSsne43T8IX18XjxKdn7D2P4hHLqzQ
KNyRd05SMolb2/DISjXrIRIucwVr8WKpaI/Wj1csjIv2cpJCUNTIaaQn+3tdn5ht
qMAv/oSgRzXQviuGaOzU9DLGZ3Bd2LIGfVv+hKaLGjAmB3/1aDizGhmbe1VIC1XB
GTXXST7dsU7qIehwod2xH4pdo/ii0Rctt/wpoCkDqTYQHdxLCb1lKgPoe5SGLV5W
Q4gpZ/nAZsKS5faBgHZmMm0xnHHeAa1jwrb5f0EXxtecZQfibmTuEI8h6238Pwm1
vN56A7oaycT1H/tRBw0UrgeQalq/7YmICZhrz2MufLba7GXUtsTq9VU2lWhGCyAx
yhJGmH0GKbaKBIo8pexHa/GVGFVxPcIFl4mXvT3k4YFWtGIhcRD0fovojKlfojwk
RvLrrpIRH495LQEuFvZpVL+7mZyteXf94rFLgMawr2d0J7BwQtgzHzWnShbid2bw
f9e4pYqT8w+2/GRM+IdqKJFsq1Z4kZXXdiW92bnj/EeVrv/27RRbOZWtSnBKQ8G6
kgcZiYjmuGqZ36q9hgIOlONsx5VzIdqX4OnQwxYJmJvCqkrUtotrIswH9Jl6gKPT
Sr5PRszjcmj08MPvKdeeoUCtIPxPpRQRNtDKtwVmxwNFMLwusMOkmzzwOsuQHdLh
8keHtL9k2ftM6iR03A1vl03ujH5tRGxAA0u9fYkJIhQBaz0LmlGUNZbBBYhgp3cY
3Jdzy6g9N2ffWmcmAHdi2a5ydxjrTvnIksqlt64tcaJI1rRblpS1gQb1ugSG7wkT
JAcuMyeVGogRLaSwJQJXCu7o6gfwmZUkXkzMEvTj3CDlag2BsnXOuIpeFRNTMAt9
PoL7bPTs3whUH/HbEoCt2mbkCpLHN7MO21/qPp3UTA+yazDLdVck0TNSy71NaXOU
i4LlCZbOoMUJfO+o7XoHAxYgcSUmB1N2h8pyyQYycS5/59a/sapUtk9YhIXUw9gM
IlfWk0a4h0+aPTAIpiei7nFzbHtXJFfH6NFyrJA93dYoqHJyCgyeH4jGwV/iF79E
O8fnwdGyejUE55RnCUNIDVFo/z1fDNS2NY7riMymfaFuhWF71gX7YnSUfrUgWxx5
MCKyX74Ssk5iIDmrYPe5bDQii8XECbH0ViLdtCnSFuV6nJo0WdMdGyOrepn2qx/0
ghhng6WWY/pf2CGgYhVednNqAXuWxB0+4uXhG7s2b4I+IzwmxZy03I5zD3tdZ6aN
Mc4o02xyvVxF4lI/XsSUOM+u7NYbubhuIVB0wUnhN8WddRz7VmClxa68v35aOFnb
sf1HmjONZs0O589wDbUByidWYBSm+vBogMxtEbCFTr82G8+/SI85R6j7wfN6GlQj
r4Ta64Gec7kNiH7J8zxbbSNMe/zFVhOYoUve0Wf9wGAZnVxkzY5b+dq1ftuPVrVP
ABE1HAPl4VMd5dQ8QxdSYzJDb2GavY1fvuZIF9AdK98st+/E8CoUiL2EUZXkneST
8ul1Kfs5ttrB7boRw4ICC1ssAKfEJ9FCkGTVk5lxJTIW51M19diAx4k7tHrgcmUi
g0NvAWZhGwbfyNE8X94IboT7joY2Ui24YsP33rbSAoi2jexXlbe5bLyxLw+k8pue
Bcg3Y7+uLk89CsUWL7an39c+v+JTr6pwucSKea3d80y8SNYyvcOX+J7MdYp9yJXv
aYVQ4pyv8fUCefueoD0PQJPGFb8XuaHywJQQ/HKtoedQYB23kLomaAWceJq/0QS9
1CemigUK22yfqluuWwclOMKs+wQhJigf/XJNj8PXK0NIHR994Y7c70xp/Lh+/NTr
YkDUSQYNkQ77uDh++KS2sw69XksmsenlrAjqW8O8dcvN2uWqwg3YIQfqkuSVmISH
hsPsxtsDcxU9KzWo+eSc1rixs/FIZMQAkke81JNH4tg/rt5vQ9KUOn5O74YV8OJT
Aa9V7bkDwKlasydBDP15FCLCEC7yifSAKJZL5pUldtCLl8hLl6rmeeOAYSa1ioA3
NLpkXluzk+RfxOIEV/i9DfzOfJE0bbXIjVZbaWgjqJisqrp2TKxxb8JSiQ/3TMQb
JYGYla17Xkjqx6a4hB3adF238Z1V1wnNpRlzAMgDbBgaQLRHD4onWKOQZLhvp4sn
4M/dWQNmBGjKkkQ2Xpx2Bm0BfxJ9jfXKEFkNx2y99P24agNsdLW0KV6AMtqB76YH
kYneUWRw0rhRVofPGuSbjXJJwYebd2YW6pmo9Mmtgfu2pVhJy+nunkEqvpH1ht/W
f8meE8pC/vDspCRHRPC9wvWyqYpgA6ocM2COoge90awVu99YvMt+O4xBaE7+eQ0Q
M+/fD487jbQMoR5bujvU4K1mNnz+aAPeK4xVNiF6g0Ywb6ZDW8iOMshpFsh/EHw4
USKL+hqwcur00ai3co7R5N17pVcbNX0XgOJ8tyk1L+oyOnvQl0ygbHaC6+lbR7Pv
P6MmcdaiM/VdEDBI692vmJWeIf6N9JCxL0CRYt8oCCFYwDbsyTybA+lPezTwhB3U
jmFFg+De87elUBXwrQz1RY0RmIbVgIeZScBOZZ6iB/juGq4g/b5MBogN8Itcf48C
/UwoPp+bg91gs+TbTVsGKp6L/fXGq8Lw1MeM4XK06jwFxcDZqJwAmQ1d5nHdRqRP
Sc+GsahTvwtMmnAopP4Obd4vqCanK6do6yEvY4BoszSI5pWld5kUz3M75dRLUjwZ
cOzpqYrQS4HV4QhfgCFtDZVbN5BwUjWfj/SpowehB/+4aLnQpeLROZpicrYx+CcC
sIo/JlAAvUwUb/TY9Gp9ldvPyQGZxc9WMmJsAqdHfpy6PyqSZCGM0d8iB1yBS+ob
rYIORL6xmiiyyPJ+SANgmCILrn3SAsZ0JTM2gKpSHOWnrJGYURIsVgu/995KK7qC
soZvBDtde/nZgdD7SMw35A7b0UOg3bmGhM3I/nyBeVDRh9P8kpjC91qyTwVDmpkS
LXcHfwCspQZxq7/lFqyYvtnt8VbtPuyVsUWyowg9fjQTdGOaJraZx6637TlRBV5t
v+ollvNzZgscAtFriQ0erpfc49RkTgQi3pLCrhzQKhGj0tTZnluvufPt1Ey1ngeO
la6xDuPqU8Sn4swB2c0L2Uw3jKlxsALCTWnjRaB/KOLhYkIu1AOk5LiG4kdkRZVA
oRbkmtoyHVB8Rf/UOd7ZIa4QA3uK0e/dEK2c+Xy5s9a/5bZBGUJHdtP6yAm7S1L5
PzCDchdTt5V2QaVs16Dfxbg88tPSGrRlAIqHCcX6ksHaO6lflp1XAqicSIrMkNib
N2Vm5daAk15ZBTvZQwdZ3LMYAsep0+MT9km8vVof/5lETpI83QRQfLcDekoJbdfq
h4ZlqqDIYNLLcf3C9Y0oOz2I0oRlK1Uc8x0Cv66JjzCTiKiOJSNy96Zm+xeLIU5c
uuDiLJM0x75OfLrivrIbkLoRA9FupElA8eywnMangJSefKDQZVJNbgSgxvUGHBwS
rfk7CKBeQH5XYYymYrxGXw4nJ8tiMo0KPlj+VGiQ35hXzurQA/KZkxs3E5hQoU+O
7WOI70PJzBWOwFitXY9SBpxkLbOeX8yHOeoqWJBc2NR9Iwcslp8IskvpsTWXsbKf
8V57wdBzJX2UgJNffKBKY7VvhT/Dzw7NPoCuozslZQ9T7UkrSAfZgAO8FB94XsxA
R9Nncirz6IUnVQl/q6iMRYKYTMQzW+By9oxzcqPVDLSgrmpsMT4FIZMj6T8GSWFk
YptMo5AOQbWCXSOozNQsRQiypwkKAzVxACrQAlyadN5FkdulSFiK2mN6alKtlUgt
i6Ym2WKtDAbjreKEKZp3yoHH1ClMnWt///gZchFEFxvEhT9LM+P7L08ZnTdi2OnW
NlKB5XancP61SBy05lwVpX9ncGmwBCZL3Sg1gzjypkXzUYiNeJ41kXty6vqIehMR
Ule19ghzIBpPGh52pDJErYd2JqHnqyqFDKTdlbzeP70+WeAkjlOa3SiyUJgWo1y2
1O3WV7AmVHTiKDgKvJpn+JQJXYjMEdBa09S7chOdF2v2pt97rO4BHmYTjasHNJZV
GHNuDAdh9rmB8g1fxuJuYfM0KhybEMomAXQ0M4ydScD7A7nf4vIgrjVjhp2tu7Wv
kmWoeRJqSYNivSJnwcn7aGWIocwgrLKzf6QRcY0yg/R7JpUINqmLZ1sXgMyA0wiz
9yqbrOz6To4kjGJcWfe80iUOQFtsIc2UHSHuP01ZVIp4w92v9JOHDVLIve3+EQNK
eAO9A/Nl1Uo5CwIlld16div3ChNz+TJAEpmzQn9WzPmuWLjgSgR1zhS2wLwqQmYK
59ihJNazWUQUu4QSt23bKtWWtTYqxIqHZzTAoligHqQyyHoeg8PT+rWfeAkcMEPd
3/9PcVuDY9Qn9AQ8pU9XzBuJ8WmrSBegDJpvPYQY/Ac5756xO21U4qJPGggsOWYU
XDq9xJoAoOBWuZj/qaDZErrcqtOvRdSDATTNfqxp6k+rjjYc+8L90Dtsz/exvmsg
ktJEBz0/B50Q0VNHA7kKY0dp3pgwt9lbQE3KsaZ46Skl07++vN4Zjdr8oVLev6zh
9e7LZMvpBSmat3Ji8v23MBLMFoqaEYS244AOOJo6QOFUjDozqFWXrTJYp8h/CgNm
WSncFlx0XmnJbHcTonjLHzsSjKWovp3+46szfmqTpA/XanbKPoRWThWhBOmazSUH
Mo7zjW5ngwvQXLog9pn3T/cg8xJuXTGIUMOo55mDSRXwr6L9Zud/k7CZe8WdeVu1
h0nARTauC7zkPmImkx1cROdqQFU6FIu6y8bE00nNEPKT73KfnX6mg9UCSRm8eANI
+i7yYmsBdyOS+9XR0pwUlPL67xjzQ+N0bfYH7woGdY9YduQJ2qqMxmggN9nkKuRr
NUlgZ4+ITFrDvxeTvqTMO/rwgDY6D4UG3N4j46Dedtl+KonEYxRm2Pm7wx0SUnpG
nbGtVmnWRgur5H1mlCV9i+qzZ9e3FpAd6BmDVVibp+ks7CP+g4D9voR3azCtae4T
LU/U0XfONI7licMOESccWUes1SKajxGwkjBGceAqxWXA8QgWK2dnf4ii/ENsbn2e
51mHiTbN7oXv+83va1vLg/MM8D0zkIie75tEVu/JGVKcApXDvyKZxpTSLMZC9wuX
WeBGAIBV+b+CjrJTHDAoTFjDSAsJOuCfJohfusQi9bbVGBwJDlRpf9C+AxFLJlJk
HqWl2Ye6enoNQ/X5RaFuHvlPtPxlHQcqfJ9rXLeAWIJGCU1a77iV5BIgVwQAza0m
teLDJ6cEQ8cnTw/b7gmN0wl60QWhQUmAxYUqDr7ltj0sO/NdBkib3+ICMOO7QTY3
v9lCmyXuMGrncbvEf3aD6sJjnLQXgCc+epLqfGqT2Y12zMEieXFfjd2FudX7lkAc
j6LPwI53OAG4i266AYd5FfVFy8FQhj9QSIDlaiLdPXA0mcBUItwRETur+ruAcR1w
6Gr4HOb+MY9O6gHh+WZLqHXZwbSwg4l3QIskmO+hYBEXoQda3spZ9h6rrsbYBMyj
S/8u9SuvMMV7pI1mAI6YHc5hbheGIWcAcfbU8RduzBXoJJtgzKls3xcbSftosob/
HrdTt0f2jGYjaKjOkToK82A/nxOvRQuMAC9zQ/iNmXOSq6IkxifJpwBJqNZIbH5Z
40DnYGYjKt3fffR0/YKZtW67n+tYfaWwai+Cm5HKudsgITHQ/pdB1UYMqHoORmFz
xNYTXEkd1nhzwg4Cl1m2/xa0WaFdttdtqQmzsbTc6fclDZd3ujCIKbBo0dHFl9lY
xpJry6kGRWaf5GUoWIYQHbtSuF7dOhMqgL0jaeV3RGCJg4EwcLPYATqwKeM7RoHW
ha10/4hgFx81c7npvdGCPSP0EU2f27/mJ0CXKDLi5/4VseVddpnGG8kYJlEfDm1s
C+DbIklwxvM7K12sGBOKhX6mtyhRBvJtYoZJA+tScbvZI9aq39Vt6w87VsR2D6Wo
owNbY8gmySVHgxm5bNtGNCq8f0DCk/cgDRiTFQcsvb+mhUVTBnfj+ml/miKH4Um0
zQ62BOa8WYJsfPEuH4tzHXopG/4bKm3Ga4lV9Drw4WYPmRk3OcTmT7263djZHVrQ
7uakvuT4YNlKOrimXsQmQ4ZUPw/ZrwBTpyU0bAE/PrOqpEHO5+s30YqYsXB9/yb/
ifGFQM0shy0sqtCuppKud6LPp2aY98rsgH4EAkFDN5WuRdmvP4PvSIny0HVxLjRa
+EY21orvYNcCiGbxeBrTUPrKqeDITGd2JRBILEPHdrKKZK1TdAjuNsdsdtBbD24X
xYGWuBSpRQW9mGYq3Z3M2I7CHyLMWsOaSYqcIcG6Uuap6aKqpZ82kNqm01nMwIiN
34MJ1hyc3W7g3fkiKTfllWpwicKbRl5Flz2cgoGRwzf9bJkJOlcBJUSDh1KCPITw
GJHz+8GK/0L/oZjqi2R/XnSjf7ydWPj5FKEfmSmb94H9QrOZzTWpC/Pt4t9Idk1l
T3qiuLUQuh9KUP5Z0oUKwH8G463NVnJOkPm4S7WIBrtgBBuq9YIT766iP7MYLzYm
IO7fOhUsTHh9UegBNrI5dXMJ+zYMMNumWtecLRrAVFkwLds6La8lXCCFloJwv4d8
E+wU4SZNPmTIezaYtra092FFp3xsHeQ8FksD6bHFCsi8pLWhs+UO129WZIf8sNpa
Ut7vpQMQhR54OASwJorecZkKG1sL15R8oN/4D1vSCXawGxVXb0okeXrElPtpjFz6
60nFX4cIUqKQZg7weUuSjnWdGwQyDQLtKzqrXUaYyWKf5iMTX6V2P3+k+HdVsk0h
jDkphz9VFoVHixi3mnfdeHYU+faR1l74mfwchDMeixDlWW37nMGTAUBCKITG74cc
GkU6litSyVMu67ppU5DI5s9+6+VsgTCVBm74/Q+lzTUi5PFlENAwg6Z809f4Y7Gi
BxQ3Rdptr0X5wE5VdrOSoEpqKhH4bDZobxRY1FdwCQFhSahnN/D/78QEghb86NgD
dq/IpxxeTVYDs9RRVCF6bZ8ovZOjdsNVJdEuh+tlEyxZzmSvfZDYSX1CmY0pCBMy
dp51BsFwfAhPVuwonHtjnQjn2WnutJ6iwosCpECqgVNFEpeykpcsHv+ybLBBZDtg
IOVWVwoNTH+NJKw1Zy/1izwfHNJjrb5T6V0eaS/36XY0Ts/Sb79+/vSmRnAHm+y5
XcjHQrZZZi64B+1PXwvnCUj/Rh/o02Bga7NUMG2cEjd0c+DKUMDHWQkio2Qb1tS0
Dbzz9QSxsrqtnvMDEc1w1mKB7rMpKBw7Ur1SXMCQ7qSFxbVNOkq31oc+rwWGMNR7
VsHyXL0sNvyPzO+OWXQ2nlWfLHYwUqqQvNY0abhLLGq29DpUcOYG6E+0A8w9sn99
/PNVcyzBmSD9UdBBt3VE4RsS/yHQcdzLzMGSTTrtXZM9rosUs7PiuIBapfmMcULn
7cttygO8LnpZUfdESGQWfrhZPPxnrXUdaLvM3kNC8whAXfthfnPwiIzGBXc2kmyI
a/fTQpK7pZDbNO4Xba1771XYHi/J69XpG1H1XtBn2+m5ufGt6NPNfUOI4MdzXEGa
PRxVGbDoby9UdN+gusQ3yBij+FdmbQpdiK2BHmxfc1bE2QCuX+++8C7ziXAx2wUv
BHEd+NZ2L/54K6eFMgK874Jhmb78gL85mmlL5g/hMxtDxaUSPZeeQNfYbAturMe/
BIksyTc9sglcY/6taav7DVP3FeHwuvFGS8FsfOYYD4p80fPDWjGPWLAUiXRzrv5R
qU/nfWWhJFtaZDJSyFQa1VZSgoFhTSLDM7AFRky5Bny8cQQycfn5+/Uy3aWx1dSm
MtY5s6rUFvFy4n51REk54vYi5o/FMZ90DL3IbA49Dn3a2HdvWJTcBvPK8hQUSRFC
mcS0Z+N2sH00WFwtqytRwPR3yiM4wk9CBQmk6NqlOmAg/T2zEoXQEawpMcukWnj5
eFgP6D9fkzvnQEAExs+46hVll3CzZPoa8SZjsnoTrbBWNBCzGeVavh2qmdhGAogY
RucPQCgSs/lEWthVcIaSxWa1y0jgBVxxJQB/hWV7d4s8S62gAHmDv3XVe78fPy6C
mdRaux0vl+QhX3VMORplNWLgAy0u2vscJdwYAF1rgDghvh9zvvU0UcPqdkR57h7Y
Kmd2S4CSmgY6waJ0ZB7DGMGj3av/UeERZJPJC2csU55TZr+1pwSjZxJ8c3//EwYP
bn72fLAhSgZhAX/XnPVfBNz0nTz7XgigPtaAgzAkXsioSDqQV3MohJpDrJEwtRrB
gGeUbVGjUdes6xgqnU88HbwmCEK7ZC34B/e8+rPtxSUismVep0vTzKabHJf8yQFh
Ha4xzMJsaQwzGVW24e32x2tlL40r2s+ZBCK5bL3Kr8y7sVYtqqOvQgfoOWwg37dK
7xxYKarWQ0YksUZLH7lsUrlsvUBTczcmzhMo2eQkJ1MkqgYz+XBEnJehikv7hbCe
1eW2QvWW9rXPhPrPQQTQN4FaH4/AI1y/wFv3UNLncJYYxKDU2wblM4yN6VvRiH81
1t9Pun0EYwpLyxGJNKK5iV/90rbtB/C0KnrM6xb51YBA2tdjRZBOuYjJi3p7J7CQ
cOaJvc140m08Lu/MN+nKlNwzuN2/iSUHXAFVecd0VCV2pAS22JRCBU5r+Is1TUgK
7zd7ByBY1cZlXUJX3SZPwG7gYSQh863sS6n7usTHzid9Nsd5GTnOxROj53B/KDAs
4K4Bt+9XEHsUy1rlIudA51v6miqEb5of8iUdwR4S5VZodkSfxT1uDJamCxxRiYZ2
wVYI45rRslP9A5m7Th1FVikzkhVWTi5Rijsff+xL/XvvEZGVr0T2Cx7Y+i7R9faP
aj7i5kc3wsdjSAEDY42pQtUPI9nPie9bBYOmho4mlr2yPB+E59JO+FBprGHBCJEz
WhazSmxG48+70hG7UaGk8bxxACJAc3bqehckOi+wGTkYZRo5tT3TmttIIRcLuMIj
9hTrQlG4nejDLCXFWHL+3bboOJVutDaO04+MHYpilxp+0FrSwbatirNVBE9ob5Gt
fmLWvAtfcBQd6bXgQoKnV/c04Q7uiwnlgoDFXbdYeprBl2LONRLinDjLIgU7yTdB
G1C0oz0wOI6owB97+Z7djobddzVBZbD7dXxYEjCAZLMDYOmbkjWbfjdJkuujkl0u
QHSD2epa8rdjraGjYDdkazjWtsj6Z/EzM8WAddAOPjvksVGOO2u6GH+jFkYd72my
WgN0KYN/0Yzo8JPThB31woC9eIklHUvtFIazaw5TETxrUsZPSictZS2c9/vayL42
dVahofru2XnFo8wSPxXKKs+WtxidoPB5XpnY0VST3r52MELw3EgBvux9vLcBN5GC
RzfoO9YQsRhideUQTDOsdvSzq0xh4m5zBTGJ+qFzIxVqN5IIQOm+E124bjriZISC
+g8QvsltvI+yUWyKriO+/6InrmxBrkkh/YssUJUQXGmCbFw9c4yYxGLCNd8luhAV
AvBkSeGNugGadKHowSZrE+KhkSKlGSxu6+1/SXMT+Fof0QAnSl8O9t1VUfXZ5sgx
4KSNF+hcgVy6KGFGwrhiJvfKtELiRVZqL1H2pu/a1tFyIY9qjhKVV+Siwo20HG9S
1Oqr7xu9sgnjZHqbuEbpw6yZibwcoVM1Fx/SWkFJxAf+vOEjJfvO8bCPRByja0At
flSqD+0YIrbV4Yke12BbGSOD84mVrPSiWf7+hZgqlPQiebjxtuCp7kmOx2eyr/W/
IgIx+adXmOzcFkN1KssxrsLy8ZEAltOFn5bcRY16HtXAFP219foCkc93ZapIWjdG
jY9mNNgvAGMSJf1PpuqYfeCE/s3zaq9ajq5wozGstbZj9xenc//XAvinYm1hSWa7
V+A7uoJH341TKVocjqhzWxBO8Td9Fc+PGuf/NWCZKfiDdWfmlXD6S+RNjyz432Vv
f4dopeTxoWbrVf+A3ir7OMH5i/0g13cmy239bzBNXyTdJIxqaAMysWfZFOpNmO7R
NxCsk0ckXNwnDCLG0vInd8CxE3GlUDZC2ZDrgTgsCBZ4438GAyGndaQLbV8KdWLA
9j2+UfpyrW+9/NKmxeeKmsvEHy4HfC7HOUgQ+4tt+0iQFQMVfQl3LsRR2n7E/cZd
5B+fSle1UJuOkQUVGl9nmM/CPJpdDEELObHcsrAxBCFsASijqh2XgUx9I1RTwJFX
y62dPa4C2HoKb8ETSfUvhXDYSuhkwJFHzRQ9YkODcHTf70uE8ohFM8pOdniis+1C
BGaNmdkmUCDZebB19kSZNhdqu5C2HybyNRO0MfkJCJB4oqelsx/f0C2PV/4Dqqol
um1nHdSRqzDGwoJ9j5xVbjjsGCEzDm8lWminpjIZndPi/TqhOgL/UhNnNBhWIRvP
++xgzQabpZfBeJyq9xRRX4h7OuEdLfJUP5tRU6UZ49Ufcwde1z/LGReCLJ4SKOcd
AoHBeLWfjy5tLHAaer3xCepp1whccWnUovhAUKU4TuaL4eRscnRPys+Q7l7zSJWH
96W+ZFHpKplEEyrv/3BOgDDIl0EQTX618SkGAgvUfEupJI/nVpUz09FilZ/Q+E9l
jVZye+V+GgN2jvgUrMB2oTZH2cjdXW+71TEjriXg9xvjrmjnGRcWNZDYlGZAlGPS
zsbZmkypLI0Lc5B29GJheg5H57lLfylHYTTHF9U9QL+LltyrOsiyd/fn49yRwv8R
S1uToYY27koZtXGyXcszNDPuSjyxCQxOQ9bc32X/ZNrDqnTjWTHyMr6LcywApkJ7
5cEVfqosJXrwBnDGS3xpc4TBpHUWnE+TgNAYHzL3bYLTMgr+sl4DSKWnCOLhPJM6
jgumkxZ5r6njrOjL0SiAwny67LP8eNcnzdRbVsxoyPkqQxiUIIxZayOqJsOW7s8B
nDEi/6n6H7Xj3WsxawcCG1dVuRgiO+ktQU43SL8/lBDSnapNTx0fZ4w3otRDdqyX
jmMXlC+k9xVv+r4Hzn+x7++Ptsb0WdkK94lwg4KnLKSOOpU+ULhd1IosQikCNFu/
Atv/liXae9kmdJMm+xzq1gCL5WZD0Dn3WeFlaFgQtAh+NFSDuTXQu4mhF8uA03l+
jqjmnkIb+YBDDYkJEXKipuHpvT9ZiE7jfPTXIti+oSlKWRtGtrLowFwXnufsyVVj
twQMSK4OSuBjpUGzlPy5yqXyDbBxa/4TsOeQtn4BxltNIXAYm4gkIAWd/lqBZraU
4/Xtg7lD/V0eVw3yYmrb/BLjRrcnl00en3ILtO+ydBpFVIIh3mxD07bp+Yn0AJ4U
5Q20E7rrDOuEVMvMmwwWlfAG6ShWwaEylR1fcZ50lsjLkZ3r9U8k1kO2ZtmoTqrg
kTTOVn5Kvv5UGHRm6hBECr67mIUljrrXfb1I9fFRNSxJzfYiai8f+u6ibJIzPoEo
CTztY0A+y9MSOtWDf+HepEsKVKwlWJgOMujMQcOO3r778PA0Rj1MRBOMuFlkOyAg
oeVampvW9gl4ltcvKFegFgqwG48ApTLmfnaC3uMj53LA4tYSpXgHWnf1kI/mzM59
XIhMhr6s37NpMe4CDWchWZvFFuZpVEYs3sWd8o6HoEJuXSh3FeA8GLaf/og4jpBt
1m4kJauks7lvvduNbao/Lflx9Ym2s1LifHERCXC7t2sBQpcTYJ2OsyBU9l5yCP4r
/I4rxwOZJMBlEG7YqeyuauDnV4Wm60aH/xr4lqnPy3Eemzz4pfJmzAyOOIOf/OfU
9f0rpgrju8aJFNQEq49CokNAVUgFQLzAxz9UCy24QmNjlVjQtoGqWX+EkSSokVta
m5ejniMd7F8u/EgEYzgKslE4ScXkxBH46DleJ3rY1+qP++7w7BFeRSJkM86JLwjW
TxGVhWgE5ZBjzzWHadFeEG5xVZO/X9LK1HuUZwyxqhu927pYgDO6LE8PQINCa49Y
SLL1JenwNTCo8cDYKwHnquegxkrqO1NM3edyXYe/0UuQjyloYj7W+AS56t/CSN9u
2lXnPeadhUq4/stxk1ktcVhAB5QthmXer/F0Xy+KCQU7NZ7qjrkBUEvcQTFRQAH6
snQpCH6pKeybhchwLQSrxxKs1+o37Hif1EfW6lFkrVBV1dJVBApuZJd8vATeTikN
dAzUOYOWvOZdR92U+kWK1Xy5DpaWqr49O7qJGIoVbywcwido0nWO1FeF4LswAbuS
gxGGXWeOcTKtSEhGOedivmpyFUe89pMiolbqrogyMzbCqM1Loni+nKx17VbKRWY6
yhCvKVxZruUk5XncrZW/wVFx/EQAvks8MCii5HNZKYFWub64qgn7izFC6+N43CIU
aATBaLDBTXI9DzB/dLeBH1Pheu/5Jwi2OnjO0cyVwITVnsLGyin2sCTFittj2oF0
3bAY4JqJC1lDhJzRoU3eOc+34iXHGdDlBneuUSfh0/FRqg5XnaNM2ZioxFa+IoBM
xKjW0eNIbJSxWVJDQmn/n04xP6FqE8wlYsIaivqbVxKlRotadwjpjr9JtYQH7jhi
LEc4IGMyB9+5UF7YubCtC9SS84LvyU4og5oAp9qY2OwpPd2EknOcKKmPGGrb57Nh
r4dMJUsKgLBVc5QoT8Epw/r8gfubAfXGzo+aaG6i4lIvsAGvWv0PdWJN9ZQ//1Gl
+cfvmuE1RCJGSjnRHgAJcxcHH7xFc6ZJxw32CdbfPzJjK0/FOTE4J3AtNGD8OXqN
f2vHobMYJYg8IMbPUyLpNGH+6x2o/sGzkfa/+NYcYhvSpVpADqZbvAGjY4ZOM8sI
P12ZLwr9HB1BhVMJ97m6FpUyW0ut82bxccNjNpoJ8nwZoqdCncPnyeGXs8xbhKRk
xYXDh759FQoLvC53U0FYAlki+wJXX8/Tf91k5U4CaY9DsgsbLbk7Kysoij3oM/AA
590g9/LnDMcWfC/cHMymMk2HZtKEliENUB7f0unW6WcIb4wp2iqoFgDhoIuGKnrn
/xiRF9hF6Hj8Rd2wC6+QkhIODQ05o4IRb1g34Gs+u5DUY/6/PM/hOsYNC1CL8rPI
9NjbUIk0UsvGtfaFz3QQ9KZtqbg0QAhA3OnvTDJkY7Fs8xewSjXtOzVhzAC/diE/
E9FsFblFhvoRGXldQexGck5SwAB9246duTDmsldKfs34+S3BujZHeDWLXqFyIrCK
oM2Hn83j1IeQW9sIWKOsLsy8lLoMpCE9hYLnBuBmtPVy2gSUPmmUrUe1tomqG0pR
JtfUdOsSgz0zaFqzBXlXfNfGtMGWT5OTOcbXdo7iMrgt4WLeKVzVtvyd+j90lWYT
WjmzXC0LVKadYFam7+FcIES6+D0DWTsDf+b/tEaPGFY0WhNVl5cv81qib0byXepq
pU6JXKsK+clkX4JdwFLk+bJmHJBcvdH6Nis5h4nU7bAJxPOk58PCTexfilLfi7zl
den3EnAEeg6xe4k9sRP3fRdgNGCrIfpKxOqYMknDwubedVQui0Iz6uanffKip7Rv
8zkawj/BEP6i6opLja6bCVj6iDwIFsT/XKEmBMZFmmqIx98zej+5+WSKfKe7vc4g
l66CyQ72d5MRaaMNRbZyt69f6buY49a2b5LWtUgt0yP38u5+cFoH58cGhQyclAmc
jAKbrbsyJo41QZ/ONh13/3ob6F4RqrtwwSIRhu3DPEFcAe3kxtK2Cni/GOBch8M0
mZZGzUgoEDcpBuQm1VjIvVULQ4Cy53VUnMBn/XPL8Hc+hh+jhHSouDulekaPdLKA
K0FMY71SQXwqNqz+6ucU1WZQdCzXdCHyrQTBw8n+K/dscVWpm/RmjqJ1Cpt/VAMl
sBKXaVcISkJvVzNw5iGVygS9bh6YtzmRqtVBXOXxh8m+U3bvQoa/h7qaZf2k8eqz
Xc9EbOUMwXuQWKgTXHm2ajC0QpHbOBOPiE54PXaMaVA9itKRXrCul7qFjVLZOKr0
Y8DEaXiCbM8aBErpwu8qm2o9BFHsJh1n9oQz8JlE/4bOy+Mi3CXhuyCLs9PyJZA3
WyuE80zyDiKKW1sCXAYV5xc318VMlRtzSPCEdQnhgfoy2bE8wNc82B435NmGjVRJ
nh6ja9eK1qj/TONZlDyG7tvNINkXGUJaJJH56tHhjDSVzjBdE2dY2KN5YIlS0IGH
69UDEbzY2haNGuXJLny/L2DxsZVBemZQ6AtYJHae3h2QqPsBFPRESnPRs+HVfSmj
Od6PMqorvF/oNWKzud68QmqM/vDo0o2wE/mc2oacudX0hJ3FqUa2owU6n9jUus5b
PlQpykuYUbNiazPnq1qAPcKRz4goERkHH0Kpv9hp5L6LlhzuSOlwN/ggXIZ0/AB0
PP8fPUJZnd7zSlDwQ456rLumt1xQVjKhC36Qt8zbJ2JA5QpAfFfrftprjkSNb5Cw
9hmzQoQIr1iH4S7olyYWa3AU3sm8p9weX4gYSF9LPDykSwru+A5y3/LouYjrwKNQ
4uco9oS9GZQkecKEEdfsRuPKMpxbzEomcugGPFtkGcAvpQldifkpMVNVQUjOiEQr
Xi0S0Aiur4ugWEZKnYO056G6+VCCG28D02A1QfGGHzEXBeIiKEoqQvxW+lEh3QuP
AwnPU565iN2q+KGlql/JoC4UjuOWtTuVg0+HqH/8/rm1l9IK8y3UBRtPPvZaCh6H
yrPzegGsACxU0hsrgKQW2vWG//2INY6ZMdV1qnznbcLX/KIFhnSMlnCrdTQ2r0En
L9ws54VIe9KBNph/l5U7Aw==
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 43504 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
5ak8DVq41YiTdsbEXvarNyT9AsKyBCu2roejenrWhs7GAldWBMvm2SF5X66m/5ud
LWG4H0Hch/6PMKxjoMYp/8VDFrVkZwQNm5v4RazZoFvZdavfVNcud7utWB7fBhkZ
AB+PHesjXhS0tElW5t3OERnkvHhWe7pWPzQKQvs249SB5dKeFH3NWAFWLcQaIE9V
4f8z5yuENQAeZeb1xRJCH05SZdFWeN2YQ7Dvg/aMExSe+IkzQQrKciIa/ZyVXfUc
owaWZw2gz/gwvJ47eitxGSHCt9ZAeq2x1mMalg3HHXj885+B/R0zXYjcqpRaNU9g
hHkNPvdV2idubCQZsBBn4r1Xu23C9FT8Q7Wu79IkrlqW1MooAH6UK8RmnWNflUy3
1yT3IgRUQwNFQfVnq1KLAEvPlbKr0mddbcR3lVJ0pyecIes3xQYYTdjAzi2t1eeh
l2IdeVSLjlWLUUd27Sfa8eska+LJ61LT5phhykVoG6fU87vciM0aiuBJT0B4bFDS
TiAiQjyLNoJ0om4DzDpEG4pOPZjnCnWiWYOSB5YgiRsencDsJwaaYhv9tDGmjyR3
dh2cRKTNsdAyNyWx27wtWI1LT5mXr33Z/1ahed6JvuiVZqhTN3TkQbv95cNNsHe5
cuQOvUKiSyE2rwSYoHMxqjopiZLDE1W8H46JZy82XezFZqokVVUOf6n4lYFSu2Yt
Gmg2nf9Ad+yOKC3eKkr1mlDpVJi9QxGRYL+TAng6RK+aYFxBRL1mgpFI2mLzZHeJ
zqB7QC3nfUp6vqZnUKobOFo8y6WI6P49FeqJHD/nIQUvpAbdhqcCXp9MlgxDcmIu
3kpVnfwEfGejlVG9gxVIi5Ta5Iuw7b0EW/2bv0LzGgEspD0jOmEdp7QsD7PGByE4
N8hO+ut/XoSyroH3+SM/ndGCcAyae/YllHMOEteqqp9bH3eyGKxhlmjzsiafu1gh
/CwNPBKBJlIo5LEU6ieNDsZpZJpRBzlIlu3jBDXPbDnQxJlDMb1L0icBtKBaXa4d
JrIBp8h43kP+JvXPSb8ZNA26pTFN36/oeYaKLn+no20MKYr5Ynmv5THoL2qnonx5
uCzejyPG9fXaNud6wKX3JJ4EC77WUMxk5wblTlA0Q954nSJ22mAJPQmqSrK7TjdT
HlZvAkxvrENpLIW6kjvY1Nm3FIKxBrBBIv7+8yB5h/5T+8k85SNPDv9oHF24aNwR
ELQi58M3nzPI4if0e/kdKki+2v1TkkAbQKiEvAra75diAjjAEtvqT6VLr9HxiR+p
IUkQAlooevy1EtrRh2ewq8HjAuvrIL3xj3Leg1YZnDZQ3DiyM9cvO+wquq+Vop12
IgAcZJ5wSIhtxZQWEEuBBzZ3PNGfovVG3/fRaQy2xXhgulcp46hQirqarFrdV8vw
oAVD5W5y3pAnUfHJzfylfObnLtAL0ORdILb9OEC5hWYvIYeuKZxRK97sIrCCKx0I
bxkIj7nCWG0vOtoKlTpPLCgUs+uXDJw0SP3Jne3ltEhi09mrJK91BgQvGLPmCCev
5nWk8d3dWUc94ZbYEAMEj85RoebAq8S6q0VeGd4jVBJT10kFDn3iOdxdB679E51b
LrerRfH/likaj9AXogjZn2sFGTUZ7Vqu8nSHIaA1dJ7M5LkHPwRegK7osxccDhRN
BkctIO7XoQQISb1J3ja6XRXA3fLoHzfxnDp4OmHpZgupf7NrNi8eHwPNtstc2DJ2
ptL2TPMOOtFREVOf6DLSjV48Y1JEuUugm2Da+wXEk8XohTkeleZ0BuvMt8i79yXo
YbvV+h8gDOicX4xXLwmzwrspy6xxL8mvmZV/byBUFh73Cs4zT6XQZXHv7HVFWNFM
q6VOOvpaISp8n5+Z7SU316P8zjFOA8aZg6UHy6Z4NfXWmfHzE+OIiuiL57TT/PTx
/KDikoP+vqDvDypmZzX610HDOt31Jktls8jvf0tfW7YQQ7bW6/3mXmaMYjrUVLTl
3hGmoIJFJWEjQSgDHrafahOv1AnFVs7vTIy0WWhmbnpS3DjRRoGauOyVTVVSG/tf
atrDeHisp4LRpo1Du/5I+CkgxhLCO3P9+M0ZyD6VtKROJOAQgbFLdmOVfsfqAEUp
2ze+9jJHoyVuooKyflabNCk6lGwVL/mbXhl51n3l215lK7EIAGaPndJLkVixVJQT
/ZHpuWje4tdf+w2Z042oHsl6GBHkFjY2U+855rYMhzJuatoW47c98ZVyGqtDme4x
pULdk5590an/ocXH2xFvr+7rQJuxboPCz7Y3PFaax1M6tJ0Ht2h54NG993yNYH2y
Re7DMJ45hDqkj6KizwdyXJpQ5v9+uyaqVUb4nm33ioSRkaBB9QjiFlTWYSCHrhTJ
qyiqpoS7i0ryRjKtPz2EvoCVfwxQjc+Iw+GDpCOS6fdOLY744RKMpPI3LzBl0E20
hVxmwwaCVjhk8exifb+/auz1mVwFppbiw5SG+GO4HrdN20HUD9inQO18UGKCVeTE
H1WB/u4/p8iA6k2VEqnQ4f9P8uiXYw5PBKz/ojMOX/5/v5UGYA2mchih9W8do4uo
EgWt8fZCWIuXPmc98Utgzhbw/jauGid5Ugp9z0uPLu4qGi51GguF37dYx8Sznvn8
LzRiXVubAa69AbdY1g1HFFAjEHYlD79z36AGYnyaAyf47SQV+M2K9LJBTne8xz96
hDKKh/IkemotQGZCTFjowA4lKhwm5eUCF3ntP00ZbSjTOU2dPouRNhAtMIpO6tnx
D47plXWh4i1aKUpPHwBDOo1J3RtMtLXfsAa77ziHlDQEZi4A7kOv4ChIIOm0Jrew
X93imDVf4svSD63g2mt8ZZ8lMlhINF3ifrBbyJpIikxSB/2irZNiV5Qsg7OxrX+E
Ef7TpF5ewQ/NlXWkehfl3yxjaHQ7CZCozpXLe0r0+1f/zK/6Cs/dDYfDAFqIO/VM
cx34J8ktEbqhLeErpOSFPPYpOTAq6ug/eYfjDDOVKnJfrnqd3yP3ZGzvHtZzKrKU
Jf1rUI7zar4IdrmKs09JVUFrmo7XU6nDbZYZXd1xOIrUcDYqo7Av3eaYSEuyDtoB
Exs5/+k9IxqIjDipbK/h37olcP2997ngO1j9zovZllcit8+Wf2w+qrxT4HWm1/GQ
dTff8jJWrkzPdPaR8v1wk/+mX9BPgvvStpD/3arL0Rt0u4evyZxubOIKIq7Y5Fi5
vTyskIiondOcHkEKAr5u+IoAPIA+AkpLgJEeZpUEnxxXuFB7mgAX9vg8cQGPjVEK
Zr4436WR7Mxheg8/VkNFodOLmjzZRa5rV77u5XsoOE1j+XdBJgGvy98o5F9vrABS
3mts/i29yU4oBdpG1KW3BMeA9Drv94R+isTtYqM4oH41MAw/5m5aup0sW0Xq5hbn
47y8rFfApA7sfUvIB9Gl43p9YRGIsKRuWLFAaInSwV0mcxbxn/MWwctecnzx3rtj
IuSN3lVliuIbnbSMPqN0meZWQ2mfjF6KrR2n3h5TOGhOIk/jiMKNVB3+/0vUN00g
U/epfS+ynBgPfnwBRJ0FVhc/fY0cdtmTh9CMsKvaFUgZOMMIO4Mb5AZUptNyJGGh
oFTpLkWnpD96XQ6eKY5uT8f7whoySffQE8kMeILDdkbALVWcjN8Ow+w+N4ODE0BE
NLeLWTORAJ2ptA/z0n/dySPbhjjWh73DM9OmKVwCH+vVR3HKvpmz34X2SBpQXG5W
gt7AN+lqiONRHzhoRVM89BqE/V7V3Lg42A+X0BhwuSHtvcaLvhdEX7OawQAFK9Cy
7KTqqPPhnPkp19T6k40D2j3IGRQ5if+cFyGYwCCrRQ4KAW43EcCBuu1E9mLLdCGl
S2olf4ZAKCRw5TeAtNk+tg6t/MGQ//8Suv81zqiECTWJn80RSxeIWcGA4GFKgseq
FQ6iGA7up1F7KGBorbgYIfmjXgvraPSljsax2aebm7yzlD6Zcrx8NYALiDbnudIH
X/LrFZ+b+TYfYxLMFTmyGn1pIWFU7BkPQh8IlpnaNNOPXdjixseYo5JYY1xsV1O/
71kj6YqlT61tcHubtRxA5A/aiORlPX6h4gm+EVfATCBu/to/yKyP/U3wC1dc/ygl
Uk7UWliKAM25e18ssrJbZMt/pPu/53wsH2MaxEZPInUoxsVlMht8oyMgctxwEeoL
yXWy4AfQ4cK+vtHFhk7g1WIXptDY5wV3ELCYYuVrzZmm+70RVACguOYL55f5YAg0
q4ivTUFHt16WtX3aBQ+4s+5q/PMyi48aAnSaoeT7rSHj+os2Z8RP6KzeDpRkxKeJ
diBLkLufl9SjO/yaCyUFqDAYmblAb3QBYLC6p3vpgClTsG+Er+I764oYpd+eEme5
hwMwdOeK6sOlBR5tPH9MbTUljv9sjqfdvLgmat1bR3bO0OTV49gqpTA0b3ABr+jA
FJb1zQhyG7PyR1GdZamaM2IrCPBWhlPj8acQjcRLyFDYto/Cadbr/PK/c8HmKz39
x1DqttAtJXXV2jJJXouuiXmbW+hgrzakbxPxYfi27f42cOjDe+lTU+NBP07zQ8KI
6VfIHgDGfy5RWW/7NK/LSxXt0DrMe04FfBWneM7V1qVDvPKHqfdzNiDpazWV2OIr
3PUfvuiXhq73gWR3Q+oSq+bzgL4yrybJehxQP6YwtsxehBBIcc/lkJo4iFdRxTDW
3bx6aIEj09rS05RvVO+Eop99OZ4YdeWCkPl7q7mvLi0121xjyyrh6BZBd3JK3Xi6
3tCsxicu7YLaDlupsgdFTu0N27ENwhDRE0/cm6x2al9i2nbLO3HqxgwZpULw2fu8
hM48vt883q+MZV8hDoU7xnWFnOLj0Naly1Wu8IIttpWbY0kTWnob5rA4nc25Za8g
134qzaQLTQ9SKV8GlyTG6G1xi3xMY45Oko2hXJKGZyARFUARs6iRpq4DRdr6bw/s
Rud1EOW0dcyP1Zobl5+GdwN8jKZAYtazhgNXS3q+5dTCpO1QQIgPPrrfLHFtzfFO
mVpIJuZqz+5R/AEivIYvq2mgpjVQEc4X3QA8q34ux5izOIZR7HyuK2+gF0GND7Ih
W6yRWGTstY31nIC+GMhO0hyRTlsPh65qgUarcp2kr5GhkhC6RVLT/q0UeD/btHdK
Kkx2B3wfq3B2cYZIpWy5zxBp6/jrjjXKPpP6xJfhXaP94/vGEAnVmfKwuUy+sTmM
aRmJELf4K7xvebeXNyY6AO0DVixZoIYQlMAUZ6WlYR2gmjIh7KnCWri9Ptk6HFi0
OOhsJyJncMxu2Z79qjX1bfq1901quAb/RjCPd29TZL+lVWABmy/rMSis1E+4ZAVO
UJi/cHRhEhWBO+HUZ9BGLjJ1gK7fAP7nWvASK4+6noiNQrmTk8Vc8YnSCHc90uzC
mcKM1RmukVv8vBK8L2mvxanNLs1SQ4D6R2wguBG3ZPsBGXaS6uL1MLhIV8U2RY5F
8Ok9dXNvnD0Kz7NtLcTNG/lkFC1cu0tSuJg82+X/spsURxjdvgSLcyXXi81J5jh3
jjRfSg1XnCif6NKKL7rcUkxRWboguqeJ/iyoTAWoO28QQz0kidw33ph4xUEM0AsI
GH0Fa9pPf9Uy0CQb3RRiSTCTdE2E13RD1z2QnAz4coMy+/FTSPaD2cNoMySq5ULl
T7MCH1eCenQ/kK3M/MyLbnuKIPuujfkqQwB9K2aIMgZWjLhbFMlDxFS7mTOHUmQ2
ndhUrQFFmoZltIS0ccg6NHB54MTI9D+tPnmrtU9NBKkyNYWJJFroFZu4RqEMoT+1
YapjFkGe0F7HY26+ufSEaOuw6WYoW+02b8XLCHEmwgf9EojqTyooQdE8S81YW06V
6uC7zkzYoYNCfax1o9SipG3UuPptA7k6/xemhmEoRbZQIe9qMZw6rVfjTxaQ0X3N
nNEJlyQP7QJoA5QfZ4NOS9z9puDpvJlC1jlhDO2KjeX5zwZ/wuSlWEa4DIzgqmgh
4a22WJJS8BdPgSCa39kVpqbEtLT92VyGbgKgEa8KzDeO3dZXLUu8csLzWmYxJzfw
c4FSf/TncJw0xFqlHZYmK/hBf9yPwc1+GeTHeYOWZwiRhonRWBjca0EV5bNvnWkd
GxaVU2jm6e772AA4pxwrYvSeQHSC9IhVaGH1JTZ2hhZukmSl/SuvnSw38wt/Z+L3
Usb9fAnvx/9P02kYfw3AvG+lZqrVf9WdMQ/qFzQP4RsPWDpkFxeFdG0X0etdGsqr
syN4tfDhMgJ3Rzjg86coUqn29CXU8z3z5jlGYCRWRSs7MLPUy69lhxEGiuVeabsx
M0Fl8xiPlY7xmbt1Qzki6eK+hn+PA/TmnT0JGsLxqrF98LoOsJfjw43beseBocXJ
s51gMQw/W24qPwfszG1n8oq7V7KCTNlZhzWJtbVA92APIsZ649bogsRnah8UpQH1
4Fhow7r904XL+a4BtLRqhSPf10fgaXtC4cmDxHPCPqQ47tAAINxiRNvP7/gcV8+h
++qd56wjMXUq6gIT6MdCGvAXaiTUZsQKkkkfxkSKSule6/Zonx6C5BmrNSjrx0sc
PER/odPz2aDZhsSrhMDDbsv87aHjl3/481WioVsYqh4gCR3S7ANAFYOGWfol3jc9
7mlbcUFCxnzLYl8r5sLNI+B9dFhTli2n5/ScDiWZEwKWKpxcdpoc/yOFJh4Rr2K/
o9XridyGDeSlbex8ZgQoX17TylEwaluc2lDJo9tz0i4+qbDiqBrtIFjS2QHmCf34
Ppwir13K7+EkwfO/iI997cmwooyA2j+t9l8NZXQbTK88radLD40+oc3NL/Gy+0Sw
ii2p01MAU7IgDsPEE53T5lvjNTxQdPVyWZ6cFHT67xzUYzhimX0johQ/LHpwplAl
/kY8jUb2lZFMzbLDiO2/asX7+cLNPFXO8NTUP1LEUIqFfrHbVOmg7790cgC7wS1A
1RBR9F3XOOJDO09VIdyALYKHlIZ+84++t7bE7+0t5L2yrlJBpQNtXzb4tWHiEbpK
BGMTlDPInIOE9NfXx8EsU7RuqkUtQkDbZn4hZ3KTkGkQa+peyWXSnLiukNfIjcGU
TeoSuQo+EdqVCFuvMloYhP2t2D55UUawWIe8qYsonXdU25dAn+1UVCTDwRwO3M6S
UOp8zEXO2KCvFXUbNe+PIJD3ZkqCUt8rVUpKMy+pxo9m5SE98+EPtRoJXP5SqREA
G3tybd+UTKK23ya2QWr5yocts+914KF5UI/97DrIy7BvrcipkPr2PUw7hGanIHFI
jTxxQReaySoekSd7wvhO6IuCAp87pFmOfTx9gPJUV67CoqUh1VqB3178R8//E0yw
GzP0aV2Hah7cbH62xmkaXxd9gSGg6sTo1eV6V5GTdQjiT0YfSXoRAwH2wA8R5hYB
3Ds8Npe784mcqFPxj0YOYfXVBcAEFsW1rXVgMa+zzTo+Qj2Rx0siOS5mIbfZsIqU
Uz/4//M3gOwrsqn3P/6uJXzIkvZXGqKwuLMcpWt48pAa7Os9S1/hQIYmakqGXcHx
RUiAm0EmR1c6RMmcbZ2JnnpxlokedK1z07/kAlCa1ZuMKaANwUXJ6IVMmjNidK8+
4jImokYSkeiUZOOappF/Ublr4se3MQxsfTDk6Becv5m8GszEqHaGRmkzX7eteWxq
Qdj5+pKrOKUhC3UG4x28+xwAXg2VzDjVN7fGO0O+DT8CqFF/L4MXgAE0wam6RmPK
YBvRNWNLiSo1oGfQ6V2sUGVc23csepF027ggx8jMvnGKr1mHkv38XWrlVNxofwWn
h0XdsiIEMc0d/3SBGDxK3/nMzK6UudADOUat39JcXaN1P2K7bEJEZ+Oj8TlaQyt+
3cbhooyZu97u/NtgAdEmc7VNZfCPhXDlFgXvwEIWDER+jVNXFbhTioL/f52yFWXM
evBCUS5NZ3Qfu3UgrFpuHF3k+ZLI+43+Ektxv8WaHRxSsuqIhjbOSzN1X+LkKKoN
RHJO6WHi0CcrWJQGxzxIVN6WOdzZ4x8chhHeIDCZMrCqw+feBO5iGrwy19yXVvnG
ZhnbsTrAaIgV4hfD/MBkv+VgLxP14mjHjukPFeMvR+4HKr7Ec90b6+DV2zvaginI
p1GfkcOadrlD05ZmClysBG71P98ybk3X2qc2g+IIuTMXDnE53bZYtv+f60NVWVoO
8XxuaZfKGwgWG5dOfqZCqfM+ap1NL3LHpT7PW0xaWxXTWeYST/brUXyeAzRpysBS
GDdHIt5Wc+Ay9txulYZksMCA3QwD+Jl2QC3L1Bqsqra3hqMVSh8Stu5OhddQ2MrS
H+izBzheb/3D0Ge2FigCE1rWxZvSE3+zO7uRAsw7fXfIFDgE+CGz/lEmPHkXd7j5
PCxABIObkOwF53eq7n9lDoLi4ktbaSwurpYhSNSQ5LjVAuJHK3IlMz6RZdHsyMAw
DEu4b3kaFPjr1IroDvqHhVv6AQnJLUVT1SRDvT1blzy8/vAhI9WthMetIvykHcgx
x4iWDxrIhda6svGLTK1pKwrT8tqa0WvuKj7hSncgMz7+FsL9kB5884hUsEyHQ3wZ
0lqF3n4AhydAw+AFRPs6sjcmzYIMNwbth2ePwQgjHXke6oB8GwtpZbAfr9SweoDm
+oIhANvUV2aaqj0s91cMvc87jDKbhyBcWaJARpRiPq+bt7X5tagrYbOH8iUW3IvY
dOg+/Lc+9Kq6dvdcpJhWG9uwx2eh8ALyGSlbIRNEL2AbHKvHpRdmr4fhQ86JmSJD
ZIe+bt3st4dJ/dxYTVe92xtob72hNTJ/m+0Szq8y2rkSEGz6fXTC5DQvrY5Z/rlL
Ydbq4TjuqmVhg2EKilWAFer2j8+hlf5aF7mrusaJ83kI+yselqKhVw+Vg1pRrj73
yX0aZQJjuoQFlX8rHNnQssXspDRrN/TyLLPlDDNR17T4cpnc3mq5hmYS94BckTsM
3VOkRlZSVHN1q1qgw125TUd0orvJQiERSerZaBhhwIOiSa38ZHzw+Y4gnWNki/40
BONLdwWwT3rxM4XAlcYIeQ7dsIisfjc+zgERLj8Z0LrFIYLJVhcr7T/Obv32WPrR
3qvhaywort7oa8D3wDft2QKuWiKq2dNOceBeVkX1YQOCNm2HHZvp0JzFEWFb4KqT
YHvfIyu5aUFGiwe6UsgO5p1T4vT7B96V5ex0hIjba7Q2+3/oGaWkiG9JfZKKtQfq
f85ys36wJCxwBF8yszC3In+8z7kf1l+mB9E3cqVrmTnT/thAZxeG8j6sMh+ntMh8
Mug0ZN1miLzHiPd5cTV9oTpk9ukId3hcVJmP4ULeedA6w6ULP9Sx9dOgPnqQKh9j
yNmQVwD8f6/UDxbV+PuBI7CfD9jtfWL1OAwtmO1q8rfx3UO/yWtCXykJUq9+SIYD
fK2nlxlqx7p7hx95pn2prD2XmAqbQWGIeGgF0MtO54a7vo6vYHbEUZv5SBmPhrEh
mB9niAL6M7iMkdJcGnhs9PHU8by4q7VIlGlf+qlZUO5P6g3jxcciWILj7Wa7letG
ruxZwuWHVmkj7LNYzq2VVJTTAcnCOQlCY3HQIy315NvvYPMmHt7qkN+iMm5McIAD
s1WnClEtiKTigYndaaOaHS3jBCrl1lPCw3ua26JE0X0WTyxjvHbRFT219nNN5BS0
u8mRE9rvzdUJxSfP7Abkuog09baVZqURwY3KDDpNGrW35GqvL/i+bn+Dkc87gQ6x
p7riZH97JaYkaij1GVA7q65W4mc7/kXwuY+Du3TziaflGOGNOSnUYoSWghIK5Fbs
xU3ympzKuRZhmsz2/ESKy5/6BSE2X3HHKJKZ7BZT8g8Dx9DXtEfduvdi0g/JhnxZ
e+vKT3/ZFSf0O2or7tUW+SbWM4c3/WIzUzGj6LaRalu0AzlT7qrb70+Xhjhnt7vE
oKXs2vAex7d90S0AyZSkyc+k23VtOk+p23MJP68Dv3iX147xP8aHkt7J0MKsF47N
PO6vJSsZOZgrRMdqwmdNVPzeyRlzl2gY6DWJki3G5o1aY7i4aCC9pbs42y439Lip
jNUomyOt7bC8/DjGfZWSUV1SM8rPkHcZnBCvwTBp+ofJIyVeQzMd2952/iVb2orP
mGVMTf7TMVVlUXcXUdn+FRk+o5U9fRXBWjmlOdnAjIZoLnShNMeIgRipTuKA0dVV
yNELlWaSh2nedieMtehf/SD4U4RypK6yUJwg5igKAg/HKcHmc2W4ZImpSehlC+/l
oy8BKEAVpRruZ7VyHJ673eyvuML03XwP7R6RW1Fxl6bdOom6BzjYe0qs68hfzNTU
4Xc3OZaKfAPmLqxNhQdsAIsu+EPCOUoqzGR7m9dTZgUK0tp4b7oQzU5qz1tVXFdj
jSBce6pqGBm4CuOkIipJIf3XAnJ3Q7S6YKFpLXlgYG62E0AgRZRCY5cFv+GCbycS
F8m+m/cQ5HIXSfMv7XqSDk/v5owOGIZAGVLFMc1Tc/YIL0WKOtAq+lLc7FXotHv+
FVlPSwvXoXSe2JtoUS3wRxkxQxtg1zGdA+Z1S9Qe7PdZEFK3qUjs7BLypetaQM/V
S3ZbzNpaGfvmaRda9CMsdwwUEOESFStzMeCORZTbT0eWDBm+e0qhqL8z7UioTC65
ByWXh15acXMq/rUlLkWMICI+65T62zn8A3pUo4xMi/g+GtaDXr/qTo0wQWToEcGh
CKK4RF8BOyEkLNUUpw0JaXDMmr8k/qH5a+ehEFbc8JvA6eIgmh7zOglwffzAjP7k
U5Sd/04WOmr2GE4UE7A8F76i0P0VKw6TawW4r+d1T0wz55OqVIXc3lQm9nSW5HlV
NZXgwEuBpd4IkBSvo7h8oU+o8cDyeoSQ5J1Q9jj8k6PRYRqPpx9YC5UepB35dVNG
GsqN0DYFequRjI9Xc2P6Nqp+/ma4XaWx4QK+Lgv9IJlhS7P5SnNay/G/gqgV0/0B
Wa/Qwa41Xzwj23yqIWvSt61Q5F5pRA+ChL2hSuX4ZBd4cpslD2ULpUQj3vxXteRS
FGy0Xsi+3O22dVp27uAoqkC6N85+7BjSrCkfLaNJ8GcGfT5cLuPl/9Kl5n+u7Y6I
Rl1kqOjWyfYD6nQz4XZFdpmQ1lnPuhE1KaL5nrluFFwPlb4a1S/u1yrQMXAfqIq5
jT7ShuYgD5I2P9q6tKcnyoy+8de4GFCeyDXkajVBN0rprEoe+0f09Jd9E/pNM2Yg
WsU5XXhUznqCSYAKkyXJ3T5KPgT9tkAJghy7mUUsX9FBkDOdaO1sUIZZSbTsOs33
DaZSxX56KMNV7mhF+rux1J9FfyCByRib8BpXlI/ctLQ/4LJcOao+JEhxL2xAAljG
nQQAzFHg/JdEwzht7/6oWIlFYjkOi/Qnz3WHQ/5ZozTltTxzalsd/6hrexvdcWBd
cMIWSHJbfqxrEYfrA6XQx4Ogjn1tAJb4N28dXiPGtSIAFQLDD60IVsI9XVdKZGCI
sxpCNe1pD1B/fGF8XGp+yOYHa/kYAgiFKSbtNNMWfribpgXP7mp5ZQrSs75Rjtiu
8kOp2Q7olD3eihst+7dS5r9VmD6QZ7mTnKQCOQtSBzvrq+x0WVxIFy1BSM0K/pVl
cQCgwasBtv2XP8pSvR2CIxZVVvuZUeT7RgHN9vRXbhWfaAr/tKa27y3ZrJmJw6s4
DL1jcOTpoLCRmhE8DnnvlfQ9buM5ZDQfPUTd7wuH2jh0hux4gimo2GifHZoQuw9c
2n4fjRlmmITch2jliicqeWq6h1E/7Hy49lAI/4lBJGSYb7gAk0ybpk/DYyvCw7PW
g6xeJvLTjgEtaZ5X3S0rgUqRmg7UIxdaH2rQ+Sl6XE4AOvP18F64JyhI8UwRLo5o
foz6NqtFkcAZiW9Aq1wmK4mIz/KPOZvu9mKPgUgz7gQ9INCeK7384EgQ74yw4fUZ
yEDCL5GTgdKwD/kL98ioT+ehND48TAqGaqbvHNZaRQhryJ83wswwa/+JQrNft8UB
rcq0gmAZIaV0XffDYn9LcZ5q9RJopRqmt1Y06fDhdB6s4ZKZSFD2NZOcrO3iz6kN
EpbuBU1CEEvx2zUI/h/7gBi+4GnK4F5qMUfmmDPpXB5hGlTxmDSx85qmdmK1nLQX
PbnudVvV/3mBAqPuQkAX/5v5nejdZizzijwHl6ENHqLHaT1KKRp0yQI1QAcVUL+P
ULbFub4asBFBlQdnrbkNcPEj4fs51uT1aMzFaTQdy6888XswFk29m7I+vO2M3WQe
Fm4xp+3+C16WI55Z/1BI2OHH50+4+Hw0Yv/7uQmqCMwri0Sl77tyagH7UbcM5+Ec
FgrSLMgqdRYu2sfQvKBzCg0EE6jli9Cb8yWcJjL/VGDoWfLH521NLZvzIorc2CVG
kmEakyZMXd8U/ITbRN6aJ9OYnov2FbAeI4PM2tuyKwEbV5KK3uZkqQJQF8EN62GT
9Zv7yIEcn/vFxTS0m9Rae5YrIbxxImvCEkj3cZt4NHo3CV4tRQ2ni0PsgIK6KPqF
5rdj2Tyf9kKITIXFhGTCgk4C2bnqSk0QQp49s1j15V6NOM6B4T0XeMXcWVGmY3wE
ehsZoBx8hq2IxJHRoeYXMB0HlW4FjGbRQmcc4YaFCkWxV4H9/t12jNx89zSg+u8Y
QS2qKM+P4bkFA22iC9JtrVKgo5mGEB2Nbqkmu3BWPKEkv3EBPx5185MjABIcsZVv
MFRpxFKg9/5e4SMDU4CxR2yxxh8WbHiWW/SLGlnxRjm3as3f9Jo47d/NXcEfFLEo
woWS/+G8+EDhqITTkcrNjak0Vwtxdg23bJ2lh0GMTDyxHrEQxYK0H03hR4cG4Sio
bojwnXB2z3wOUP2Y4vsNOwE43W9qzLIiHiSf43Ysnj9yom/l67xK39swNstGczgy
o60iO1XFmIDn0Vk9FiOhs/N3O0NE3JLR3ZpFLSFPagYkxhMoak04KnUjdE50tkBr
fMfkcZHWiuXGx+NOTQL77QWR+kHSYAbek3suqpCF/AiPzRXWihczyIfPjegKDIg9
85giw9go65FE461QwSO92QHLeKVM4Ge+YWWxc/7wu33S8lCNn7CO8hrHzTLZOj3l
HAccvePJmBIVqwv1Yj2PMAlDtlBfjt4e27MzIhhwZvEOyPtREYcxIYJ/lbt+gG+g
w6HBzOkJ25az7oGcb5Cp1DFp5K/t/2/lIfDwt4tOrJv80ViiEM+K8Qfgd4aXgJ9K
C7KE9sGphPZuMTsG03YHWEdvBEKPf3+JSaf44xCPYr2zSBoHEKtecHb7xG6uAPmT
ddUa6CBq8ZHeNBWZ7uS+gf+WvEgAzrr6qLWu0tUQxsyJfa/x54On7r42Sy0bxR2S
HytyjuQkfxUAZaW1Um5S6l61U9FTQN6LaMA1loOIV7v+4y6Mjd47/OF2N0ibG2yP
kdG+0Oln0+/ULTRBJcNLTEFYWxOCvS72fXQofxg2eb/FpqKtgHJzzmJkJoZPrEuX
DL96r8QTnhxoMa4tt3Ikuue7hpNXOJIrLtIRznnsM9AcgoIdKOZIqOq1X+fX4vJM
vn1HT9OggclY7yhFFaX7Jve5GTXePuqR4beMNbhKP51S4d6/LZBCIRv0ttiCQ5TO
TCxNHA8xc33sFi0xVl3U1rW1btWtJ2t9VbihlSAYeRupMwRJOYmlvNpYjsXhqB0N
6/17/GkDKZqPzwPlQTz0hYgUvE0mrFeLbPdbMUjPzT5ofS7oL83D4DOQaxOTrw94
BtxHXFH0pjGe7zYYpIl7WgP9FyvnFUR/mqu97b2fdkOZm1H6xVyg/ZLbYI3qRR+7
+Gz5dW/gknpQ3z33N+y1JGNydALRpHMHHG8QuzvquwkVpYlRJXoKo53CB/q/cXFB
oK3F0Wgfzw9NRSClxgoNmxzr9msV2k1dpIZYiS7MD6mOHgCRRuosj43iUvm1uEzh
aPGpkzXWSoBVg/ws2dtmfgfvj2Rulxwj9Ek3OsXXSU04M+ITqNhYp8tLk26bn91o
74scRMcpy9W57OJEH41lpUFQV294V7l+YNgZFM3iedWtkrwjSHiwCC61I4MtiNjz
lhXOQdUjZmPwmcZOTWWpG4XZDmd7QD+ziWSnznBygqgcK/mil9en/wUJd4EHPtwO
ssVzE4ZqYZ56J/UAARamWNlWqCXdYbt8J3jhHqCe2BO7VstbDcWCcLcP3G7i1snF
mdfyi8cM6A3X90szxMeE5IyJpt6q0sPNcwWchxqer85iPrw+tjvW2RT3IbT/2Zbl
aArNiMuJuBZlwCVnyWj0Dnf8eDiOzP8Q8SIUyiiQ+xMRrvGX57lEyv45CkBVULqX
d4l6Dv+tdb/glkLs9H1MpMSIa/4xuVpTxeTfJGBNc3t4C66N6zO3pw8yf8wSUjNQ
7qgEVDlJ3A7e0HRF3wFn04D8/H1MNtdPdTwze0sCHULCJBTVC28lYsqgabEkv3Bt
OVOecj9bilhiN+vFaQDL4T6CRpkxMIzQPGqmYBBdHEDxg2sHmHgsriGV4BDIH1PH
y8050Isfn/jZQzXT6LsAjf932wt4eT1oQ/yoap+aCjMdd8Yd8xvfsssR+VzIjBaW
/c7IvCID6WRjIxB4xJt07ADvxK9LP+5+yk+pkAbjWNWnTd3DEmbD2ic/yotHhWg6
e3/fOOEaSL8RTZhMQE21c0aNarmDDH2+BjHs2C0wflAeDv9mGJLlFS+7WSkDH4vv
1Ea15k7LxTa4pxk1XJDPzSBH2MPy0jHaLal0RFULXwqgTVaTzPUmS0z0pOfD/kOH
ggnEEN6S94n8wb9hbk3FHuIQ+I1EVbG9j6gwA9IGe4PJe7HNmUcn0f8DedKmop68
lB1g3fJzoOnkV3JRtpABNlUwO0i3ZXeCj88jrE/mBw2hN/JirFHUyVm6zAEypRsx
UmygLQp8dqHP9DwhGB6BqV3LoA5OTpDVNQH/p+N/mb/ef0hlliH0MrLP6MWiQqYL
O675MQtwTQuN4EzNe6NcPxtppfldnVJG90qR32dIO3YEXY+urltK0w9/ovmuzHYN
nxKzFbWcbGy8Brz/FxYdLYxXKqc6E3ySLCnMzgDja+fL4v3v9/O+5RKEqpP6YjQL
WZZP3e6NAw4lMFhedJ1P01ZkUfRAFVmMfxhimaGixBe8JZyspZK1RhBP8SIx8nol
y0CKfNF+IqRq6dBREfsrThRfnwEtwq5ag91TYtC4S2ml4ACyAA5CmvTiH94mcQGQ
wk4LMCXq874u+kkbnJ4VAUqiazIOwEQpOZvr4xSoY7EG0r8fELY1XsPuThmUuXdJ
TzgF8mnhUyek5xR+AsGLgfEm9M3SaIxcfSGYfH04ddX6rJJFNslXFjy22qavDWdR
KBboKWpr6nNt4sVxfgXUNXmZJiO9yfNgwZlrkRdJzzKpWH25t8ZgTBlldRR6p/83
+QUfIVQfRTPpL2gCBUZ1ijr5UnN5oNXyXuf1rw4r+IzJVDPOptsP1DD88O8mTFbD
+yLXYO/NbnqRSrCev2pFcpIS4KG8lKa8PvVx8CZKH2b0uVCy3hagzttzAdcJaJKf
CbIZZEpVd9NjieickXlwLPODUBr31NN60iy2XnB0LhtrTUZRVjoMRHSa18HSC9ko
bvuUrL3XF3AnsUXAhKWJtBwsu3CrAvLYKRl5E9ug+nEKbNpIORO5opbAo4uO6odM
wkA+TwfDPamCpfRDNEs7xQDeUfaMYhG1mNkw8u5/IFBO0/02hdjOIHnoGnwoKZIc
86pFNv7xexAjYa/3gK+oUu+fE/ghm5/xXP07QviwiNi6eqTC4O+L4SoQN7wU4sei
TaQfbAj2PJoK/M7tDDlLHibI2IGXWyotGU2j5Vfq8KzxOWBNnT168qn3PHZHKa3S
Rn2zgmrMEz45jpyD4S8srrTUjXprw2qaijnsRt1vSKbv8SnqY+Myxpmn2+D+ZzpK
7yne+WDJ7PNBxILk7KqnvcINK2o2happOgdK9JMSX1JOteHG9/5Atk7WgdIkYMR9
L3zXYEtNr2Y5/RWV8uMyCmYcuYeTvJW92G9Y9+vnceuosGUUFKmfejtu0zaGDgq0
j4N/9lMXo2YU1RlSqErFlc3YsmTAqUAnVrIwLFNIeYY+K2+pZqOePIv8opY7g8ct
Z1tEX0+GNQ0p1QSehono/4Zizj0JjylRphak7F9qsdzTcTB8D7GyOh+CFri9/WfZ
HXRp304TZzHVX1BFwyZgg57iRCF8//f7qc7PwMGOurAlAaLNbUSdZmB1LQTFkqcZ
X1w6cwR4s4wxmERfHL/FA75Xtfk3KTIXNLHrgVA/OthWmNMQHgrLMt5bHFuFpjAt
+S2I3pv3A8J/7G8b8xMMOXt+bkbCk5QKimIr56OaskxGbTL6rO/BjT2HRguAwKpX
C+xHW0OKpWkC22ZQyGdcVtRz3/4mM+yw0nR2lYcrsX94taOSvK2wEERz661yJf30
mZtBdtkk3uuKmx4JGwvxb+z0Evize0Q9Jun+ZyVqO/12d4dBD5hjp052r/Kzoq6D
txXiUM4i+ZPWh1kQ1uo+WEwj/noXpZbqqi5F8ATzf7TTcMi61/HnjC/sLl5qWYS9
Xpi5227V2V7Vqx7NRMz+FLEOnG/XLWRvOBVUDwcqtTcfK3me7eV6lGbbaHCNXcdd
tWssqghxL+2ODW/aUVEQIzWTYYnxCHnhwpj1ekIKwlfxHqpd06iEBZmo7CuqUHht
+5Tfwrpe1aZaxq/9k3Av9vxLpl2NUt9yzp0XVgbDSWCTrc/76AlFWrRFLiqUv/1k
mbVA6hCvhrHRO5lCOApsC820I1v4/I7uo6hKquNvNQHzuzBwGDPgCDDI/BH73cL/
ftCq3R7fVAPNkc9FuZOpNep3+WdlrFGcVNjBThWsHm30cqGb+xD673rdkybCpVno
Brgb8lbRStrqiDRBzOWBp89naj0AQAPu59ga4amMcPUTMHZfAn+kOC8TOlfAYkIk
zXmcIMckOiTb1bi9f8tXmNiK7pJo8BeTqbhneRHLqfewjwQCzqU0JdJX/v7JIioZ
02pAwrOaw8u+iZwH1j2pp++lHPzFXrBBf7tKPX51GDl4qyh7mOY2C31s9DNzH9xp
7B3oCpEm6FWS5/wFvg2DnLmRqNGwnEqZa7iDEJ+VMbnSd7zWRgrUJliFv9+z9KEL
YBT6pqM+Zmo9EOX96KkjdaTZvI8Xo7S1I0rZg844V5LhZ9Q+L++Rj4FFdogf962y
Yl9+ojiT5TNTjmj4OuDmjVlFawvX6g/MsEk1IrACD/ECf67NLXpw+DigeuY41ihg
khxqDubat7I4jF0j6tRzmAujTl0ezxisgb2G09NcnbfGJcxFh9OvMXnsTw2GkyvA
QYJn0S4dN8dzxPGUek4lh2/mXbDi5P4OMMRwdPOjqN5UafnTLONYLL20hEbW9myW
dwH/vl0Q/cTzjyWjorPvl2uNw1X5nIY+OEsPjQ7kgWHMnZYOMwhkkPhrsre+ySun
I4jwJ3pYhxD0afLvPaXyl2YQALdyXE+RbNjx+LRdu9zw9eRIMzb4tdVb1RaMdVqm
Tz+nWVNFn5gluGY4JsAbx1qogEP6TwOm3dRauXyxuXTGfMBs5OYDnR0UpCTZ/c9m
OPeygevJiAXQg3hDxzEMZLRp0OUARl9kvbJMtzZSefxq9RqMipHFJxBP7pZHJWWQ
GLjtNmLh+HvH8sbX2oKnVWDKazx7sVHGE2Ek+zqH6zEFjd5V9bj51P6fR2HpW0Hn
1mfU4oPjRNr0kPeXhzS8hFj5QFqlDqiOMSOi2mXUXhNmGOKJJYtrcT8/yEClNNL5
hnCiu5JbM3P7vruS0iGY+BhswaVa7fQP5tW42fwcrPZ41ILE2H2LoU0mszuzsFBK
YGPGn+A0U+EwWfgqoNDOe7C0W0jWpb3Xm8Ipbul6bUuGjx+fR0kYkHWoqnoqVvF+
BqfT1V5cHTIaMHPUkUyBngKtPN4Zy14uLiWhlrwS8fR/KTQ84sQQ4vgiveW7vlpw
Bvh+57dLN4kNoBk77R1qJkoCZETkZgrf3SbggqFkNKpm/tXTiCYbRAlVvzzu7CAh
bexQJRsdfvRJUB8f3fkFvfrOgTHtCW1S4AGooqYuoWKYkOCgnve3FPZ7zdtVarNI
wPFzNv5pCnp46171CQeYvdnn8PpoG9iigSvS8v8TKMJ1WLY6uAwVj+m/NSJvONsJ
HVtTY4EXYxydIn8R/TtS/ohcd0JMy0gyCrp4AK0cFdmCCqSy3q6pngJimWbtoRD7
exCvKEZrwCfQTjnhxVz6eSRvVwC2yCnaDpwBNuh+NKRYLi9NTBeC0E2Qi1aY2IWm
+9k78GOavK5r4ebQBWb8xqfrDWoocJUyA4BswLtZQVx1JPTJsIiM3OVTTCKLNWHQ
A0gJVE/Qkq2MRhro0vd/9Pla090uDhw0lGpMah9UdvCJP9H0PT0LlUtJCtOtMkag
vdMPrW4u0f//dfsTXvsj6KDK5hIWOT4XK/Y6M3PVNDo6EffLfp3UMxN2TLk+XHJn
3R8kgPkJSbPVpLYS3M/hx5aUGAWM2kgZo/F0GltnA7MKG3Se3BlRrnS0yKV9W7I7
A2woPnrhLfXeYVMrJy9stEXQlSh+70A4W+WXebzWhJp0boniRfDNdjrlNNVkntZM
h/EPSjKqHfyK+faKVWGN7Y46kTqIrI6aO66WjfhWyXrY1ME/DSyuQoWcWJ9TpaBp
hv35yLKeCA4asc6MdecrNTdc55YOZ11qOQ/w3fSTDmUPJ0jagV6h920h2HkwAiL3
nO8LR0FoR/26tzFsrW1LW9PoGRnsfvMMZgZrTP8z7R+eioZKNyRHIvPaCnZXk1Yh
gmL+KqshV/CXNCBoE6ID7/fVdmVdt50002TVd+2y+wCCF2C3BNpJkjeDbG17TJ3F
llEdB4KcmANfG0j1eG9imHWyJgiDrjkDU3JG02kTCR1+UFLldFpsEsnKIZHCJHbp
Yk757Z3LzR0JFn8wNo0laMDjVfOhXIQ/R4F6sayjEFFMBRvFs4EGU/36YnQZRokS
sJsUfS3zGGRzroTkPFj/b9xoovuSlFOcpI+E8ajTyA/G+i75AGgJ7tIP7XoaxGHE
kRwidX6OhMFJ5qA6JC0DvGGCbzs6GMhb7mCVxxQyFGG1Y76u7DfkOVPlHMy0R2PD
ixxevF/xOWyXpqvFqOzWxJrFKgVzkS14P4IhO1JWuLlKVgBFxyK+0uA12kvQlUZA
3X0XPu35xOlJUymmwcWwsxxrlAkydQlvfJhwkUnLfYVB3kDUVp7rx+YPHCjgC0c4
g5M+dxoigEEQukTgWuH6Va8t0Ez29KxC43v9SmGH545AMMbW20wGF4ChGaXQDugE
g4anUoiMudczUUjpwT12Ult0EfoXkokr8zSGdIquzV1WGggnkytBUo87QB0Praw+
1MD8rb42Fu7P6PUTjxmu0a2lbLbfdL6DvLl+HZocu7luSyA8dOlKNalViRQ3yThK
902qncg3OPCDAX6k2bJgryodrPpPdP6KCNmX6+ZE3jSAQ/fmxi4jpYUw62SXDb98
rVPtMZopyK1R8QI755dyhemZhua127GFGkRIzF2jXt17KHyn4qY+zIbs/tNaYVk9
rmYoLws2vsW5Sm7f0gYH+kuxecY4jZLdoTM9RHDXI/lRWKUAFQiweitJQSx+zCF2
6vjFU6Y+LUXTUtQ9r2M0DZeHApqDlOw6Er/lS5jOtuN5gxTfhHWgBQIwAv/i4xne
WAQemHKJlozwRcnAcJGy83C/5dk+tddogNLRikVbDx7q4EH8xH75Z1weG27AECHE
UmoRR1gFS5i6Y3FN1XXr6238KeXQ+O3eCGkRb1yvbgsrp8TMuZLXtKgJSQwo2vpU
AUuLZT9MxpGdttNR/uqlNRxF7T/XKSnN6mGr3YJduSUVH3tnQr9/OyIjdtndSkyt
50fAlmCTAsDCozGCa8CIKeXFQOET/u8VguGB4nJ/AocaqA/B2XsX+fwwUMNcLbjp
etzQXQS59TYI9jjQN87Z4XG/iuxBnA+u9ZKEweRBg0n242wo1en0+gOcGKd+/J9h
OIqjIGoU5Jlqx8PV8C8k2Wb0rvMozlPeTlfoHX6XFlhkC4CVZUndO0KW0EFOi9n+
QAGlfXP4CwxYG6cELsE2C+uuZpepRr+Cftp4UudnzKoYvoDuetoxXgjnnlTP/FkE
AIge31WeNz3KDHkMHYgq2SdekerD5nPqf+GUI/wnqydudapU13HovLSxZXMJSPXA
7PqvsWsQ8d+/ucXC0YTr0+VeysAcbGNEVb1urMFPA/Tk1AJrqdOhdO0hq9gYqtEk
VIHqtxS+GbogHSROdaX15DUoQpLCrbysLg2LRECkBIUa1+gKKFljOfk9usO4e+4J
jufbp9T6OSg0OpmnGx9MXb21jPGH7gJcV31HcdYoEZzaONA6ZgBQDZw5yQujOvv4
ZGAMYy2wQ7u06Gp0teyrVv+x/NM0yOW30ulU+IDd9SE6Kh8im4QUGBdh+yDyNo6X
e0SjOaIT52oRJV8Nn264lPc2ylHZIvESHRG/uPP2roxngxQvTggdNMDagaRiqe9S
1+8+umcsfimno4J5EQ7x2SqwqtptSsfcWaMlF1mg9P8pCC0LbYqq9qIyzE+fkdg4
yTUI9va3oeB4TC2TmVVFn7XcCDF0QfaS9NlgHdlr0AFA3R6IS84pNRbXeBZIcgOd
sTjyN8pbU1kEIFvCUqehUtiuICPTtp2/rf43dQKepAYU2somTK09W/7muQbVGsPk
z5rzkFdODfNZajPquduH2COkF/37Dhqvku0N80rtrN4Ceygjm6V6eVA9Vybx2GWi
ywH2EeVEU/Sy8Mn7ANFrj7zAeDbpUuBbszp+oljzY3yEuyE06NmeeksEOb7cjqEx
2GPek4ESGomaiR0f7C1HSZ+pEuX1KaCwQ1dCfljm7NSGOlWn8NPmxXOyt3LIMEt2
WcCeeolrtDBxdfK2UPKF/9+XQxn7qTTBHivRnp5u/6DJSNDsoS/Lbd0eVWWO9xSF
XAsTuXRVl9QIC0se5/gjVz84FxN1Iz/RppKDqvlh2g6ux7xC73SmRvxyJxuStUeM
InTV3thVSP0uwvR/wjBi94qYy/1+FkUZYgttXS8pZIMb+JLmGqqu7hV6XW9Dlncj
YM6wie1nhnzZr5fb9aq44gxd8mjKmUKY8xHOWTA1pNM77H2qYMXjMttey54zDzxE
Zc3OgWgdB+15+A/khfLD6DZwijSHRldLMpWbZ8QIx3ERckQPri+lvC/K3OGdQlVL
kQDMh2zTch9hJnEmiNJFPYd1mw7AzjB0falTNfc9mrsfemiyaP+79JdDF2UtEjB2
M8akI4JadycDx4nKEmWneBAsyYegMqIPevSY79p91RJHlOt/b3Fb8TYbTTxt0qTP
7bu/x8x8C99oADa4bITdsrTi/YVICKJ/FU3D1T8xLvFmIXhaGnDjwiw+xNF5xJ5X
DI2A0krL3P843cocki9vIoRROieczHPfy4vcegmsG3Fvg/V1yQCIPHFDvjZQb+AZ
RsNxK8Xy81P178I27ZPndbBR7g4PXxUBREyZMXuyk0z3S2YGVXqcmPqDp5ozGhwW
f0DB3VOQnr2DKMhLrBWN1AaLkVtqizXQVefXfi9q6uwby1mbhXgq3BbVIUSAIwiT
zqVM8n9u8PzK/AxBbKxdXnPknhCRviP35t1hNltKdZsDOhDpMotsbnzBCacoVp71
oJTqpKoDedfn5zFnBGxSjelk2ljRrlvKGeP27bTLEMyGb0fA1FRQubcLnN4KN2cd
r19aGTNJWhRwDEHdO7kYVBHARaVEY9rQC8iP2+moyo6MKw+GkYy3fr1S9ct5quH5
C1w7YH851n2AdhVet9zFu0KjFxMi8S5WTah9YOLerHMdx70fSsYvjYP4gVhyZDqq
MeJhZFO+CBTnS4jLPkiVcge3w1K3JiokPG1BlnfWYOmnffR+gKcFCFpI6TT7h4Nw
49d+2QuvMW38T0P5f9mzsQulu5P65QjnJBW2bkB2uDkgFcR2IncyYM8dy15hV6U5
85zMdAKY5v9uBLf9/qxQqw8ZJyx7uKorUucIfXho7qH4oqcqhl6pEqkphivhZKHa
OUuo5Bspu7Ci1Ne0jJxgJ8tlDfx9dPLc1ydFycKNzdjA3MpGxYF3uoX0wag7FyAD
st9tgsL7+RVU3lIu4u04qidKpvMCdvo1qH0z9nN0aVsuyFCUgUtVhW7KJqtIZPzd
nalKHfHZnlu6ObGNdBOK+dKsrcjxEHwQCUjS0H/ceQ84bVYXunCEip3bvdnmt46s
8fncnLL1JtNvWYVkhWo5qXxOh5Pz+OM0qROfBGaR00pCVqzja7d2WH5vIjcKk8IQ
SS3vISkwffpP1KmOZ6bzJFgrQpdStuy+LIehRbBHJscipdBEEVicDF5OnBTbwiMe
guqb0w3289M0PFHYBAWJjw080Cv2q2WgjKW9K33q5cu9PC9UrL6O4MUpfE4f/6Rc
DqhAjoIjsZyqchPV1W8tXa7CZA7hgoOQSLAe0iPF4JqwnIS+fTJF/PsZIeZnOUfx
JAPHS8WXwVD8mtlKoGkjIXbXDOuKPQcIMgBPoRdiyHjGizC7GKYMgH64pdvTULon
L8ZQboN0WyjoqBhuecnBniIhwHjPPrctgOuktXLCfLLPq4C4NttGQTcpg1L41slq
KxqEyIiOdaTaM4caUQAgIX7cNKYYVBE7XDHr8zp1U1NB0eqC+IXtehGRzVLuuQ1d
krTlzjtG/aKEc3VtMLOO39n+hXtAf0/p0jVVZGKKXf9djdVGuyysOSnD8IhYIEzY
YQNJKzoUagXSwQdq4YUvo8j+k9AzTZs/KfKeUvsBpnWPu2OiIjzmW+Eg2nLuIdVX
Tl8CZQdmbo887+2AgHXu1H4pbMLrfArb13HqFGQ/VYg4472CplF9Ag21kVl6L5Ns
CXzfp6mUpGHC1UtbTZv+J/ZvOQjsqTWHNR/DZFRUU9vQSwUrEhMkhigqzsbhvE2h
kW/iN+vq/BGrkf24GKNgrUJoCJBQ/IUYpXabXVs/Htu8sW1MIE/vwxo8azm1bMO4
FLDaA5+p96DsCF8MRoLNeCqYOBpTl0dyD7QsNubtQFqrAurRnMgPAvSKFnYOWW5l
OtEoYxJ8MpVZldE4y/kB4q/+d2AEzhwK0hjUSMP4+odYCsvn3TOxdqDAy35nu5Pv
TX3fauPw6KupvMrgvXYRf60gPRjrmoC/yLlrN1QYouTDO+sa1T1ttxTxKNvOtbRQ
/yvB3RDh2j1dF1wQsfD9Re1h3W26i1PXgpj8tYwOjn9Qqu3rRNxPgjucRFn+ML8v
rB+WbH1MpuHtBQvwPCOI7xxBPOLQq97q+pyVC12m0kJK00pdkJtYcH1y7Yy9AVO9
TlHhzG0cgCxZVvZfrJcVR1JV25XsBvGMX1NJkaKvnRLRje5tS1kSZgm9mcRlKrY4
5tLRP4czyW+ILDPM4RdezSWf7rp1Nt/e9F2/tlxs9vcQNAUCUa49oI8p36B1EsIk
3sYWA2MKVWbZ/q8TrtYJ7MwsxYEPAfcaWcUhAnBnQAy0mmWzaaiGP/N6PFq9ZMwD
Jv33DJerE59nsZIETsPsxIjVGPPLEFQJu8OasHDl0x2Kbi4Qay+YjNxoHpvFrqEY
zZOZJXGKfnIDFSn8MMUE9xXkeVGecN4LjzOJ9Zatfi6ulLFQrrGpcj+AnO9qYmGG
wqOL0mHn0SZUjEy08zXG1jsERs25KBQ230XN9EDeDNDejwm8zFkOEHVtNKUwlnXg
uxvcctkm4tcJxXNu40Wfm3/2RnJM85tNEW4fLnX82MlmbfufgFsmWprZfbpHPVo0
YFV7sQCTLBukVOY1qnkdsuWCszXmbfQ34RY3wBcc+cgrF/jdMTvIAGwtSN4nyo1s
BhLzgJhwNX7I6E0XlHDZOfj6if+O+4CRBnJY+5vyCuE1cd4LzonkcDIVc0cxu9kn
GYqck4TW35yPNJggrKXhO02QQYq4pRzTjcidf0vRCNWiOqj+ouCIcEX2T1J8BoMs
Uagwt2kJUz0qP8EUtNGvVH26tHU1Dd7VDWh78iUF62x3J+SZuGcGsghnhnWp/zV5
4BnR5Q/se0CricNmGg1Vd4MZ7v+50dxrIkopwgineOJL2MZyc3JlmuKzVblsPT45
GigDs6aIexIeQJ/Ctbgg1hqC1nhq+kD7NeyNAfQaED+e65RlDFdSIUBMXVZUmAls
UKybRaq3MD7zCxl49LNjnBXhoFcvRnHPu4CHx/FZo+/8ga7dLO666LXINbnbg3i5
02dpjquKHhVeSmNs7QHNlcHkyvTL8YKyqQ9G42oYW5PHwq9+hDXmmKkQs0okLyrN
KPHQFlFvsPqle3MKH10WtHe8C0/5QACpUnjG4nT6TlqXbvkOAN8d6htJcA/DJkU3
3+DgwrCfPiTDWSqpUvuhHsns1vvON9Qh8gDRxtjmsWAfGL0it7aV5ewlwwkQq/Vz
vxdrgyDheS/5ET8jfD/6zWiO/OvLSoI3xCoxTTBIABXBRT2Fqb0KLwStPv+A+Nqa
rycF5kojsJILtxf2M5bbM44VI9FbD9MEk1WWmILo3+Fhh1u3NmBl9qtZdX2Hh855
6NUX+5lGcnnDCfVF6+Idv6s0ZjCXFWhdJ/0ppHQJ7YS2HXnjZjoMlWtcKQ+A1Wgs
za973cin/vE41NpS6NHW5ZCDRUtV9OKX8SFPdYo/ssRiIm+L/W4UQkhyp2BdzY0S
fYPuqwfmL9N3BCRejSiiPv0Es4CuXxbGZvHyWC1Efq07a28QkJtYT/xFxTKR9TzF
HmYlWMtf6SZW3U8F4KLXWnAuMEXKxCtiQT1NZYyTaPwropvGB4MBOAD//KYdUB4n
K4RYofcCEUCTYKvUs28SHX7IS55uB17rl82oHhZgjWSYfcKYr1uGN8RvqbtRBANU
F2B0euzMXfArfD+XZSHabcG2F0/M729XbPhjLh4ZorC8+FRLsz6BxsGWKQujbENH
5yGcPGHHGryHtt+daIAsyY0B5wymnGDnUz0yTFuQvoiDEwWuS140HAZIIkK10Gog
JFMBng8VAmuLsPXahQNXm/PFlHSN4jB8uFipIBGuHuIHB8mLai/KLqe8HLRs4BMU
ppYnWXfGB0lVWMDEymyHToifiBDR2MCrC+d6Iyvby7hyjjVIAMx5cQsLiT+Y/Hgb
qAcFJO96ohIX4xN4x30oRcDXkcN7C9TmL7ADNezYylhLZ8GKraWeX75nvTGw0vWe
kxeChLgxa1q+af4zpxr3+dvIRN6INbGpKx9qhs1vnYTj2A6njI+sCWT1svm6Qfyi
/xtjimIi1h1LpDt0/i2u9bkL8Y30YQELmjF4uh7H5RiOyo91TAB87m/xUMzQ1tUo
eN/UuBVMife0E3a0Mc7T/d4a/mRWa7buyCTlX1nH+FQnIK8Vhk79BkQkiF9zQDy3
2T+z9CGRI/DPr7ijEDJ9lQC53YQcHkJEr0zdVQEjid94tYRIHbQVAf3c4PKpHkN6
d7K2VyUOiu4gKqOB0lH4wtZYTPRh8eNRDfu5+aJsZ5H861C3oGN//AYgebkOvfoq
GFIx2OPqfh1I8D1eURFjhX4ox19eqLdYCkfEowzaxwIbxG76GEA24ELEtpIjbqCh
0BTl5FJwLdS1WNH0DbNL0OX8rmZ9feP2VthZ5lf5lrqsfrtIOZP+Y4sNtb9G/pDm
S5/Dxv6HpQh/XmgSGr87uT1qcgmQDMANAew/CR5w+9cD4H9qEyDyhO7UHblgyCVI
p8WWvGv/KGRI+R8lojG4Hng3RzN60Pb37GNAMVfETXwXbfn4JO/mAN+9IpjDQLqT
lmAbYIhMRWNYwQduNLASg12gX+qla9yrqsG/ytmqUIEN6QMBuzLcrq7hY5E+Vk3r
wEClLeMAZA5AMF1noVpGDIzky1dfgc3V0yN/XbbbHjdmbpZUIPhrnNUJjAOsxOjS
uo0/byFRzV9n5L+1kHKQyD/YUQbj8lvEVWrHR9ANw2AKUecXyNpQXxH5Rb1IFPbw
1j/gt72msx6S6PnWG9Zfc9Dk/83hZpkci0dYr5WaWp6K530CZq9+1aeEB1vuwHd7
pclPKasdOZCCvuPLb/EaY80ZX302XPZnVzlg544a5PcU3fVGXcdkFO3HFlm22mko
8IoTmjPhRVAiFYELZ1zyF0DWneUTxoV9AhQhA5GcW00kqB3LSSVYY7VAPs7YBoBI
wck/SqHlYKn+iMyV0idzxTu5adiigZyiKvmB6G7lBN1rScn9VI5Vf3xUwp4N/bjo
iYp9wRQSe91MPReK5+QISG3eEK0C84g7EWUE23/4qOQAPyw+16QjeTWzEsnGf9WJ
ImvOi2AYx1ip6k23oGU5XlaFz/6Z8i+caNdpMjYa56eziSW5EtsoHUhJwITInDh9
FZrscD8LL/Jy8TIs6OzbVoLUoB3y3V41LIXf5wpodeFS2gudciEVcnYa7GTP+RaB
DpVetFst5+XuF6u25r3e8QK37ztVswfNB2D3BBZHdHOE0zPMJTlwjJMb9YGYHx+s
WRk2U6C+LEOZefkHz9kW7+UuS0rAX5xB3qvb7afDNAwv2JMAm5NiZXeJVBXegAMS
VJAi+nsNl6YF/9uVXAAHMdN3Eweunj9PoDMuttrK4aZAholxSUY3kwS/EFuePDEy
Bo5pn+nUUd+Ns0XTh6qN8GHwKL/i/w/URd8DJBU6jcyHCBQcjbTlWCZZ/W4P7+g+
Mx2WQZC4CxU8Qt1HqcE+P/v8C+jXsn1GFHIsLka79c9x5MAWJ0aq0U/S0EWTIqxS
7wkGlo0MHjTMTdub2mqkgD9F0f5AkoKc37Gg5fOOSayUpuPPERXhubdcpjmMc9ws
ZMSzdce8/CnmHAY2zuHOxk6T0A20y9qlEZcd2Ho0sjaiXlOV8ds5/M/aMC1xcAPY
orXk72EhmWxpRTmpHWgGkibRci+ubT6f6Nbo6wj9RMB855iYlx3gFG6X0oi/UW4T
/RlE5yIBO5lIJxs7PYhO/H8ydz775MtWdqq3Xw11FofZ5vLApyk17UZ9pHy1CzcF
SoaUjDqDiYAJD2p/aedFhSJBgblCI/u8DJdPemoymfEKRMbzDMMvQnTkDnMAo3Y0
0r+vFmRyjwjrD2XocsB2UdPmjViaFdlJgxUke2KDvNGo1cW46HEpbA+OzpYmtdA4
WjwQbu2TEFfjvNIR29+5B6qQX8Xqc3OA8qG6wwb6nmkFDHn7C8W8SmyZXElX1mdD
jzSWWk8zbZpzzdYrY+khJAslN2SksV0IKX+nwN3B3W9ZoMbcovgjgW+C/eaFeZg6
I+CZjHcyA32qGuEwiZ1fbhEYd5mbhYcR0BzoJaTkCAslSYv+F3wfVpGKNJ3/GF3G
xvTU6dr4rwielg1Ne6hEIZ/ADZeos6CrwMoUe5Qm+0G5DfdND/gAiPDFXuQGu+8F
4bniBW0McEA+FiupcrQ7wB3F8mcrY33DOneZHc1UU5uW5aiMUUS9PAcaPSQ37lyu
I9qGlmljtEq3IoaHHb+U9dezKIgXkaOpTyKjYg0UyZ6STu/l6uMZ2QU7nFSDd2Uq
BS9l729gyKjIk/KgLy5fuW+TnLbKwa24s7A+oq8r/tt0oxr9HT+DIEPw3Kpmul41
m+x4hwzENpsmZvtnZ5NWADk+l11PgHC05YlfiC/Dj2JpMPX9nZxmqdLYuhhctd6P
4iQIeNzp1fAQLFsAQzCVN5LHNil6ofeczryr0elubDVAOBPVubz+Zac0yBwgCLkR
M3NcV9Jduv2ieajD+5wwX1b3PXuVI5piMKfm96aVLhey1/3nnjvew5+azYEQTAYx
5VJ6SKKKPJ7RFwEJCfgrtbaZfVj0cPqy2YQwa0amzPNz7GvnDBX+XrrQgTH12++X
1Ge31mvAqv5DlQX+Gobl1AHIqfEhXI/PdlwxMHE4X8I2MYC/W5Ff7F7RJ51YVxIi
ZLRDd3Hu+F5BcG2zuSVzDozXm20Pz2EBHn8GPqYuTk1CjNZR2EUj2p30Lg39gw1S
CCUIBGQcOH+sKHZjq1UoALRtBqh0nUYSfozz60W40KXBGGiucjU92Py16HA8oD1p
w3SiJsVzewqLbHqq5nMHm2+4KQiLbXo/bkgoaXxg3XsHfw7p9cE9Pvye5SX2fe0O
+u+Gvk92Az/c8fFBn9U6efttroO8+XIPi6xGOpPHXo4fTz/xZsgLAtQG2ilZXwH8
hZq+yT+kxriHocN9lieKy4RXnm9Z6PKo+ZzUszj3PyL7GqoymN3HJ0tOfs910Eoz
pJt1AuYeJ19sHT7HqKJRIpUcNNBajO9UfF29IBHPWtS8wLtCcva3BZiQ9d3cUE7i
5UX2pCPjZztW9o4rHvS6Rr/KRdojhLiIFHKiPta1CjKa6KuSRVMxqbpDOqKV+5e/
n/25broaTFJpojLgmBYRoK6DTCkyaVCI8FfqZzNR0k+kHI10NsaMLB9jsPTSsWFS
y2NDaY5OVrBnTnCgOt/+fDAq4bFs3cVmKG5bM6T2qQK5R0I4b6QWj35Pv/jxb5lr
2PTJ9MzY+TM5Uw24TIBun9eMglKyVUPLJr1xL7t0OBKY1NMDMUxgJeiF71mjNgme
62sO42CY5xqk9nHktWHreUM6OUUg7ZA4Go5+B5fZdFPp0UySppcEDkRCmFq+4LTp
pxSCoT5Vw6SUsrWGIIlfmeD4faDCVZfWjVeHudO2jV2lxOHE3Va/74nteQDc7n26
uHvOPxvvyGJV5WHZFVJ+qhtGrDty9m1xfRJyddOm2SZ+m3zwC/d7jUwD2VDFky/v
NoWehpkbC7QIyCHCKv9CvpQeqAQFuLjhtRu3w/CuVQK7QjKczLL0Qtml0KWBIyqK
M4MgPfnKkU4OWLlqTN6+fXPH45VsW+9onUbkJuer2gSjMm8yX3Ng5m+Y9xUiecU4
FS5tC6Uk3vASdE6LOJs5tlc/zoAtnxfZ+yNmKBmFrvOmd2CZzItVU5V8W9K9pYXC
eOv4J1b5mD/nCrofGr7IMdVEjvEMXoJ56LfEQE5LLAn0hsmQ4dD+3i+Ny77B2kJT
qJoSTEGk3OcK/2GcH8GNpWr+6LhJ5A4T5f4jeoI0ZxC6IZ9Xss2ygbQo0LjpB3JZ
oa4LFRtNATs+jn28MwlTZ6kqj8BEttZUISogw0goLxSi/yFibafyOz7QHh1/79O6
sQViQVdeV0d/EQC8CPyA6j298Ku+uWVnYE/hofPdfnCvGLCxQl9ebeu/XUyvJt8l
frh2GYwz6Bzem2+ndfdXofDTTsI01wfTi52GrgRoabJNFO7CHRgglbHimJJQIpE6
bgfaI7xIF5047CCWgzR9N/S8x6puHiFi/XhqMx4y3DOl+bEDrUJkJBhUfraU9OAV
DmOlhTANPHk1bgiLLkOzCWbv0IXtE5ZHxOjj6P9tdXArvDrPDyibR/R/GK1/ybjq
aCFwJdXtJuSeZy94xcIUFpUcatkbC+bbXJMbWS9fnK8c/b/qhcX9QRvP6TrWcHsU
dF/LD+alVyVp1S/N/9VehujtmswD5t3hH4TdeYqmN9KVnC+EhKQy/Y42NvyMkA3Q
qzk2PvqA+y2FF+UqIgKOq7uwCcH+6yIcG6lWCqXIE4XufcI9Xvin+dwPCdJZfy6n
wQ9EnZPIUg0rQAr4b4zztysVUE/BSbbaaoBVfmo78UtH68Z/jvJGoVJaCPv1aTlW
Oy3nKV7lkEm7dGm+fXu4e6jkJjphA0qZ/BVcv2+v6Gf5/BCaLSee+d3BAYdzQ9vs
uxm+ufZeYJPG58xjHdYoDDOaGP1gvxXRjzB48U4w7b9/bdlM97mFrqqebmFiqlDP
xB/7pNRu+mv5Nw9yVQr88wqJYZvPy6f1igs62bnUf7JW1lFgT9+ghbO/B93O7u4O
Om2NgjkTkJg0gXsNqSlQA4J1MKasdLEbvgUMUnmnMLQxjSzfothmK7FFY9gisM9H
Hq9XOv3i3Rr83/KhFRvPgmwjmzqYttf6AZ7ZSHKu7IfRQCYjr5lFbCpgjeUTt+CU
N900Gvm+D/4x2NJTzRYZDEQKRcx39RLc1FpCvzpuhEjVnfpmwTemdcXGuelq7S5d
RkXD9g6uUecs1dK0ZUEGfG92JonwMmZqmZrf05CpAQS6r89eg5CMQLP6V/aCYgxy
PjItWYp9qsv4Hu6Tp74PjrvUADi6Omehr3qLthC8z5i64xA++V2lkjDmb7uVAlTL
7xozwOQJ79wh5ItnoMowWWh1ncD31ySohReVlA49cHbiD1U4kbM2pS1KbUAEZXBH
eoxZ9FfLtfvAjwZOX5jbYvCS3oiUfQK0YLEPiieXZEpUr0vOmiDkD+CKKPATH30f
v1+amSw/H1gASNCu5jJHlMFUQBWiYOUq134i258C9n5IjRee1x2c+ZH8xMiIJh4M
dPI9VTpRydHBkmn/du8CuHh6ss1FrlNw6Tc8HCK7/ND8dbWtU/JEIqWBnJZVnG5M
vtnxio9TnzPvr9x46fiiysSSHyznMF3DpuZGvaJs5FhemafPjTamQpcLhw07NdqR
lj9o37449qjY4RaTBcwxokk/qzfYZrdVG7oFw2gGsRVQ/i/KBPVwdYJ6dL9+eh9u
nHXgvS3RtzOb2+nqKxfAvVUBvmmMCnIyrjYkEc18CfTGxdCxWxAZwtrFyRiEWu5R
zEtCv2PCfydLSx0q0ByZ/eSG/16OmfvgnqlIT4AuCZUwEuAbI36E6YHsqgNRrpLG
T9npOoKMDDJTaOytCJ2VGi5F2n/5EKo/a7f9043uoAr4FQEZ+Xh+OYvhZo6eiDE4
BiwH3V0c41XBArohXczxsMQytsUxwML6uXHN9zBXUzzGRRBfqqpGltOz/ZfdbzQQ
TnS2/CkYavksdM2WjzuotzsMUv/gTlK2BihDUfHXtYETSPIAITaU2894jbbJ+6u7
yZGtJ/5dMU7zNmIO4J04t7hX3YpiU7ccLv8JPrTtoDgNWvlXEaBSC4buNfLwwqdg
dL9XHc6fEvead9lQBIJoc6H4EggOa9zv9lXed4DmA9OL0PtFtvDUWql4CP45L+p3
XAqFmm+oHMbU4e8/CfJ9snFFaoBa/m3F3kPGIIMIEtmtoLXcvs22+bDaTH20mNa4
AHJyzJqe/vD1HRp7zZAEFMpMhQgP36ncJqZOKZYOm7n83DmnPzCBtjYQTqub3fyt
/Sy+3Q+ooiwgzqZuWCDjA82mhOCv7cRQmJ7i6dEj+pN4MXPCsATEQDX7rRbgrUVZ
HItzkpB2Pvkj+2KF7rRSqfcVY0X17uo5dPbe8N9DxmKosc2EfKsxYxcUhX31W1wy
U1fgaDFi0Qa/RMkSXE0v+rOgqGQ+TmtdGzoIbf58tWsuuwg0XrJE13DcAE/KZ3es
RHY5FZKnFng+YHdmGWeO86XBmno7QA2lkUBexWXuC48U5gMbjptD0hh+CLxLlV9/
Qi3OMyaBSbdmjOm9umtlCZqz58/7kf3fz4rIphRoaesWFbq0Ma+8/Rri/pVtJ+Zq
CjmqmYo/7wfFSHOd8PUMJhQfHPrPp0CBi/HYbUurSpnFRjGfQJy97Dn+7wZZSoN4
qurSIEtN2+A5tJ9aZruYBEQTRYIMNoZweyc2/66eGNNOynLC2v38NFJRR+KGviYC
QzeX6L840jsx7zGXktkl9kIQuaXf5YD7Gap3vERbTYoMfNm6ovE9uW2xhopwFd0u
Ef5nYlCroDmH0XaTAHN7pHN4pZj7KkAGXN3lzjUBGLcLy9u8nA+jeHbH03DNRf/t
Lv8b1wwArrORRrxcdb/3ixcnMqy0hQ9a7fNQzz96rEiHLuI0eV/JFKl2OccTIGTV
ivVHp/wOALE4gsnAv4lgSKOXGYNAujD33NTPPkP8JlnSh2nVDwZ5PJNfta9bheC9
GICOFCVNWUF8+zuJOUpww7wcnGftMJIa/D3BiChrfCMwSqaZPd/vsGzwuvVaD9Ug
VTo4W3a5Nbj92coWUarY53nr21OLjBBULCDVyAli7mrNzzH08d+e2u25MMhTbj3v
mQuA1O8/WIg0bCLvkvXGRw4GUj0S7x9bVCsev9F0aVdhDRAjopULLXuTcVRdHN3F
fO0xvnXDniE8rhBNS/qQ6ox8HosH6XwJ4hUOuRx8o95tUePKWdFMoWDEt3M7i0qu
Z6IdUwTxKFKemuH9B3SMsPF0tnx/vqY0JfpMRduUkil2KE+/K5+8yIteBTYVOx+p
afDbpQC6oZLMVdthzydBc9yMh2mqcTA0XBB/TqpLS58/p5rZPwc9dhFU+VqeJMww
T6ZI0dU2f1GQCjXcZK+ze7i8kWZ8TDz3R+qFaBaRK373ASJXis1H+WCqvoJ0IfIa
dYvdQfSOzVQw19+9ES9X0ZCUB555WqedrVkA7uG/NMJJPSaRZPMyFUAQQxVtVycF
7Jh4k06qqfq1KoZPgi5TxasC1z03xaNVXC/J6Rb9Xb/Eh+BWgYnmj92wqleRbXcw
qdOItOesjyp1QyyZ2sbUI3a81Pjp6odQXiz6oXljIMgBAmV5S3zJ97wbgGNqsHzb
syvY0BDyvt5Yfp7sZfZJo7sqjlycm5wf4D9jUlNBnt8nJ/ZY27URTEPZrsu+8FUy
8ZsNsqzWaT2cYoHtLv00hWAjecSGGYWE4FJTm65GDjNsRx6xAW/AOX3IepmzFW5l
mbE2P7DgcU/u8bpekzxwPpk8ShT7OAOz/JSBD4hJ/2ye8SpwVwCCb9y/wSfUgCvV
tZiXcR+Q8MPeCe8sgbsYRHmRugVjbuBNZGFmdS5uMcOIFbmUBgmEzCtQF9lwcjvd
DDZgfl29ymwCJXqzU8fBkO+xSpPuZO3p01371MMhfgS/JuLTzEv6ABd/rxb9hi5L
IHDFUM3gaiAE2D+04a9LKQeWUIHYaeuOB9Vmrzz+knjseoYdtEo24N1u8YMIde2S
/jpvgcVZYKunWQuF8JxNasZl02Gh88ZTmiCfo7yQbF1+xiAU+o9rKb1XFukf+A/n
NIMAw7POJQmtUTzomE0hr5mYtQ9xU9uYihU+BDu13LqSQ3e8yoq5eLnwXTTv6Fci
o3to9lNOkAhh3i3R/+SyRCvu1VZ6KD4F8HExAqt+cmXu69hWAg3vfNWBzPYGZP/4
z5y9tMuXSYP2ROONaRhULernzPnrS8++z2QKdZqvfXjjbZueisaX+HiZSXssizG9
R1id0dKmk18xbYcGQeFBJeJHnpAlNnp6JMaU4SvaOueqSVh0rSNt3q+hMQmOciBF
Af13VQHxOZzoaiVsOT6p/aEhNj11EdnPPXN5JwPGIzAFQJEXG0szWskzCu8c33BA
tGxnAtdhmIshZush6D07M6rD8At/o+02aRSTWNNqcREq5XMNbnLyAxwcOXUwyQgQ
rx/HmDdfhrlTwLUC+fRcVTOd+RWjjSoO0kO4yN75yII83SbE8l848BysDKGC+kvQ
MlItZ+0s+in0/euK28bknGX/rNqLeEmMovVKbyRPcUYJVMMh+hz5VgWvMffP7yhT
rf5JC9din4bTrrrF7fDtPDqxCBrVajXY0bO8ldpFm5E1zECZ7LHTUNrjxqWOGcID
msRQCN+U8yghcAcxFc+m5h9sqExWzLE/vsz/WDy4X+p0+jsrCz9+1A8G6LadGIDE
8xTPh6sAPhE7evUwZ9qYBTrVJz8EWpTQBrbs/VweXxEXowvzmwUPIjYGqvqIhDPG
AYxTH0qtUUlR1tJlw2/LGNXDSiLoBA3X1SWALTZ09q6G8lm89WRE6QJBBrcgZdhZ
wLh4LeGO2BEnf0fcmifVeJocWfAT9ybw34V3tsX1IrU5BeZYGfzaEcAPTZpBDp4P
HMD4g7GHHRUwNFjoOxyx6oCw78X38M0tt22Ib+/7Yva8B0cPe9bsHOW3Xy9e6HIz
0AeCRTB6JArZ+5lJRbzGbJHNyeArs2Wp7J4VdZZuqgWfS7983hLMst6TIDHnkcWG
8WWcIMd9kq6LlTP/syIxH4MPnG8poHMRfWlCf2AnYoHk2tjkftSKAzT14LnVOJjc
NIxIu1TdCw0Gk/JQGqvnOZSOa3Kwy/MgyT+r7zg2YVDjX0t567A/ogb1btc31cm7
05MS/0VFTkmoIEBAKRKwSsR9KTmYRd8vS55JCRy+x5xYy+te/BCA1hqFXhOfkl8E
NQ4ZM0HjUHXRq0avLNBilEzNX4H+MoauMnojtI8cW4RLUec8FF7I69p8G1gePwsC
fdajbwhhOb2y0YCvL8REn6BBNxdbmNstdQa5nZjlE5UM3IIv7EW0VHWgt+sSHaMP
i2nJZUacMpI6F//tNy6Z6sozR8XX24VewJ4PnY2TXtd0Gx8JwmkSvNscKrmVqVj4
1mKKwq9SHKc2+JkqelK+z3icunCutWbVr1aFtvKbHPZUBbms40+y+mogrD/okd9R
IHaVgL6JIwJEAO9NAvYN65Sowdc4CfdjbyuwzXYlvmbP3qNXGoihT4Cq4bIRWa0o
v/oEcMcvLytsxI4AqP3oDqiZCVMTLel1BM7bpM5BRwtJfuE9oFfRqtqfQ53dFzue
Z2wSvEsRFA+a3OoHgNTO1KIvE3iFC4gYZqMFXxjVrKOplU7xDPBwZtIR650Sx4UT
y++WWATeW5oCWBPx7FW9PEEHsVLYwT2VJk6L5/byHXt9HjUHr5jrpDbzd5TAv3uG
7biMnEe3PFDAly+wSaBzA/5c4l1TrgsO9yFrZS3zlRxYo8bKUmLuCR+ztRSxrBvA
5mmKDlwo9GFtkjbrNia0ryiXUbkLVjROuleRW3L3PrUSUHXnOLpbKkXASC0cs6ym
Wo2IpPdprdZiHOg/HgEePCj3D2XbevaT9/gL364QJrtT4+jduwKs0WTEcBgJMbP0
7qA+d8veIxiA6giVNnQmGDOum4f4euQadqbCgZ4vQ0qa0pGJWs6Vkbb9EOoMMj4S
oHTM2jFErunxtbVHFNnZh9prv5DUs3MQulf/v3ezzwod2C92sortcc1CroGEWyE9
/a35nhvxs4eLlufjSUlWNvIBpIc88PkRwMUrGzviMqFRK9rtZm1E9mbU7bLHhxto
Cy/yoGrxoFCIT14WCh/V+w9XUGc3UlX/gNOAiWE9+gPn4Jl6o5ewxwrxUTrwyCQD
0VcXnuIAwNPjiu076q0UVDgPFWqYIHHT8+SY3dQC5KTQSFZP5etFj3G2srs9u2dy
aN4f2NF8ypdbJLCsKZ2crcF9ICjxoPSIYHmIiiQOwdiE/saPeXA4FC3cNF+9WQuG
CHH4ThmLA5SmhyScRiaeAeyrY1FUIb56P/nlfnVRLigFrmSWd+r/JLj3I497HZpZ
36XBl+FleE6NaOriut4XBnGll7NDHEQDypzpv33kmr6A536KUta7DBKSxnID4syj
bIBA1bVaB2VUPoPaJ9WSUlEMfgrnT/KC6f1dV0ZirauqF1NGZ4CEtRNBx8Q84Dij
LQAX8RESBnwrmcbtiGdcoFpzSTHY1wfvBRziHret6RAdRqIqkxsp64F1czlhEH9Y
/OHcVBxA+QBYUJmautvZWf4bsKa7W9o5JpzaQQAFFJ9PmHbhZVZOZ0g/spB0ILwm
UGU03fybblqosed8p4BL0pDW5v8Uylxx23tFYU7h2rn//FFplv5OeX77Vn/zIryW
zQTGZc3HnSDBIrdTVHSn5ATH2/uDnHUxNjg0M9wzKbVhfYl6fntJyDpWYgwcuYB2
kP6MIgyJ3ebZRaVOB6PaQZvbNG+CvRa1lMZMykamnlh/EwzvzlhONmEAjhIeaM8T
i9uaTA8ukAfnYov/WW++uZ+voWyOBBwwsf7U/J25Q/pJxxqF/Vc0ez+VukzydMSN
1lfJX7NKOj7iGPJlj4TKBICJUWqRSaXyitEUDCzUjDMiCjTds4bG+Na+QtD+kQSe
0VXDbxjJ8ocF2EMAXjYfPl9XGzZzXH6UEL6nQrXaamarX6xOXvGH6X5sLHzTcXng
eNr5jpBTEXB/Z0cc93mytzraLiVQyLIXaT91xawUCgfM/oixOIarXXsJP/wQEthl
x39UyXox19wOZafwE0REbOGDdQQMqd1GOPBgH8tX1RyE7T0mgWvh9B/rPDgby0XI
gynXAWhO7ivEvhrbo+HqhMLbj0ObVkjlrMjE1/K08G3f2WST+izCxP6GcNedymY2
Bg0aXAJpw4anysEqci2bVcIJCxQZg8aoCeSSjHd9BA6h1Ch+7grtfOnbXtZmRhJb
MTx3Ln1loUZlQcHoX491/64WyXsBiLtkCVvl1T8xa5k2rOv4jfkP7EM1/Vtwgqrf
0HaAFQPgXlouyy2DM5AneobbU4lk/kfz5kuyyiesiByxymBVq7SZGYlgdDYy1Fc7
MidGOgCq1KRDGvtMwFjv9dMXlG/SQBAV/46p9BHVow2XvpUg8ldL8lywUPHVpeIm
b/HVnAT3Hf/N6tKCwbL65/9eMFpk22JyQeL9p4NnCIRTSTdfAYu9M5KdeMzu7eFl
qMdZBv8/uhOqj8hKAnqzR1K+mu3YiDcUELNd5qQd65xdxmmw7wllCoph+GOYe5ii
y0SF0Z2fEuA+ZoDLQjdezYm+1j220CIWidqYL4iwZMOepPZJ+LAen4XXg+MsYaaU
PgSzHTv3ZlT7iB3SJlsQXhGHRmtR9zlwHGxqi6hzdoiUbS00kTsUKOxLEsx5ObVB
TxeESKFpMA4ogkC86tJzgl0+DLGcYzdk/DLDXQKf/bPdKgKgBYNED2IcJEjEnj4I
3Hw3akXrVwLcv3dVxuK0eXzt5AcSAyfcH47Q/eIvkK0xbNlBLNmQqc7+lzwPKr0O
1yC5eCylz//V9oYw4MYSdoBDnvUBpgOfJSfcR0lMB7rZTndDH3jI1Zw+AdZUy5gb
M5TVrClmw+C9zl358q5YBxehlc4Pcbst5s6KP+35zNpO5ASKwS2x9WVUMOz426FO
KX8UgUFfOYQwysz/5MdT3EWXzogpF3CZVGNWY3LEmSG6E5JbGwEs3H3zE2kNTs6S
BwyodzSTl09am24ZWkirFA4WiPcZSrnaSxiMwmLmQ7YmNE0lzYs9rTioUWgOzVtD
/PSAwCQHQ8tpFApklEMSATac6j+eslLLLf6ZruuqfqAYPDE+/Sd+CBeGpM3+YeM3
J3XSw8StLLpzSsCKyhS9RAoetlzZkalX1bRlHx9z/R4lei2Rf88pVh0d6e6py4ns
60uGMQCA5X5UPe4QASu9AVLJyYit/sMZTh1cw0T1MhoVNuLbRzy6o1QbkacSEocD
Lg18ygSct7XZAoaATQX9fgk/5uki/JsEaSWgUSXABxFj6mZ2D64HtkUbivKUQlXh
nljmAgCBvbdhVn/VfWrocQ04KhQO4nCmjg26yggKqPWXPxKJUdA/oGmmX9xfqwB8
4xiMusfb0CypA4c9aUYd8LHwizqsk9n6rRbVFlqFdK/YHtdmqg1bDhsPfhsqmdvT
/Jl1bpMpGF3++mbwxfhiVSsq01XvtMSYFmmGBksY1r6G3oiRyDMkzqxDV5e3kCwM
cdO2sLU3JfTJa2lwOV6FXG9/R8UIjh9PqSEgF+cQoJLlVz6+zpQkGDseMqeQQ4OJ
ADdKuZEDwss70X8H6G48sIFZ0GKkr57r24TK5vdCHm3PVSqv2M+Emc+tNz/TKXzE
r+TtlqxxkmZnBK1DCsaxsSqcOH/XjAPeAXw3RGRdli2vRyLS7BNESmisDGVm4jjl
piBpQVDbQgCaYbLZ6aa/Aj8cd5YaKU4dppNJs12RKot8kMFPcRMKEkUuQxMMEhgm
Ftg8942UE+iDrO6swm2A4ib74A+WKWKfTWZv2Iyg1wpyLGn51/W4iqYtPjuaRro/
yS/bTsPNfJfLzc5GFPVB9YBinwN6ImTjiljUsxoGA3QjTgIvF5QfeYQJfyms7txO
L6zfnvzO9rNQGVO6GZEVfpRZhQGcu24Zc9/Ni1rS2JJIKF7fUNjv4AKqT19Gh+MX
9Yh5GyGth+CWMSGdA1PcfdKMx6afMZRlSl8BudDbwbfyEh1zobFrwBgXqyNuVZzx
2vZID21B1N/zNRTUUDnyzd2B1rJLLyw460gyCV7goFHL/dYMwfZ1mnsaivc5k4Ym
Yd2bXsLrToQWvQnCt0z0L8HWbVSCwvS36B2Ia15Ijz38h0d4sLBp1ucTY4daAXZ0
rrRmBVGVK6GgnTqwAGJ07w9e/R2/v8GZvOjW0Ap2GLLH1kJ5IQAbb+JhgHFBXBcD
wpteG3nmBDbcTg9qktAWx3IiwTG4aTwvv0pFitvTNqbTAKJHnR5TzgVCynFXyj5f
pSCCCfyOvjLA2SmCWWcm5vTIaZhM6eX7dO2/b1G4B96/5+VabiWzjfsQElBMC+4/
SbE4kPiDT4lDHSo9LHTZLQNyFERWexZOcQuU1JKvdV1pj/ssEs4V/fOLFfvPWEvF
RjYKQJ3Cs92wRzdye642imWnRHfbEBZ57bUGc8/b8OW4ErhlT62zkIseOiC68X0E
womSqPhY6K7+38xG/kaPJXQIfV9SPyJJurFu+u0EORlk8mPVuWUrvqlrxtl6WIf6
15o8ldUMydg3O/chB6oEKLmJ2NzbfjrMSKAIPtXCpD3W5goL9zxYU5DSTgMJ5ko/
st9NisQtv+SAkZx3rYDfmX8lOU/BWHjExBpjERAJkXo+LC5zuiYIQWHIwAK7t74P
skBnYAzvGv7Ucj56nfGUS16EqMsLIFpj6nRyuzTunaL41MaqM49xiWbvi3s5U6i5
z7QXCWmGinnxrecMbM5nvoWm8iHQrOvJupGJmhzDPcZ2WQ91W/IQmiGAz7IeFEea
vcm0VRovtlxI+gHYKUHSIk2OOAvdwtnvhUSDucqBQWVXJMFe+TMWUAIMHsx8kVVl
I6eLvhzaYFwssWMkyOZrNbGzQysjFqZ4TFRZbNLCx0+B1WwEfEb1r9t+KDALguYx
4K7STFDWF3W+F/vfCrny1CYDbmVlopbEqRnrG82W38ZB8rAZhidcaqkvp+eMZm63
7Yk1/BM9r4EuYPnVT9xUYu5VdINsNeNFLb4BWLTybpdIq0uNTFAh/AQNqlpNJ4Kh
sy7RIv5UWGfbb99NEuc1O2Zq0t0q8HiRdjw3kYZTljOAGPLJKNOgaPJpnHkELO8s
BKbMwJ0ZN6HrK6eNv3GRrqVvwHELuXbdUuw5UVUgLext58EOMNkVvThAPjy2nZm8
zNEdKvQwNTCS1iePdcUAE0jf8Q6gLBf5RXnVgwNOXYROyC9Cxibw36zfzDvaKmJy
wbR5auls9FpSaHgmHHo1KA46E7v4gkfkNbN6Xc07iC6lLhCs/C57QuqXwqcF9sKD
KPkIE3XGE2wFrhkSODlJDtoAzwVrlc0XH3A9sIxKN6X+Rt8bTMAIVJOXX2TSfVrV
A/V4CHMN4/SP48X9yzIb4crciioQEc8RlyMhbo37ZNWT0edBrd++yq4Nhe0hv/XA
iRzm+wvuMVZhtHbU2NerU8sjUEQdON0ONGth0IGgARxikJEeA+20g2q/BDIpK2ji
/4+/fOivWJiMpeoMZNwDV8UrSK4ESoFpY/fAoTqI7BOSljfDtSFIHiurHNw82z3K
o82h9L6poUGyER4ZDdEauZaootXh7zPHe/uxEX4MZDZcqHmac4/z8X1wta9TpDXF
AevGpTspGpJPSKrs7DDbYaS/hbtt02Hnt55yhqO+aDwNFdyUWFnSMjWqpO7KlNcP
QTsu8YMX5aHnxf3BUS9TY5oRQGVafYIazsNNA2W3HZPZQWRoFs0AlyOKfcuwsoRR
Gz7GLlPcm0AWpUaCzn2HfQZVglDS6FiInVDkTIBxHHnBl+MAorxbUTCAoo3++Xgz
JZ6FZyA3qEzT6emUoz9aXFWTgb5gGz8MfWhuwZ0xvLROF/y+VEFZ+9wp5dRg5X1f
ovWZ4km5HtUBynC1W7dwOVq0r96nHL1XTdGa4UvZaX/tj9tKecm8TmnbzzxpfNoe
gZujtureaI9dXfsFkX8kZ3WNE6h79JiEDXy1Z6DSb1kC5SMDZUw13j9tTM1CSYfh
UVuqeZAjIcwp1EgvKGIOMkA2eFAuZqRkX3LcMOPfP8YaoY1ouGto4ttt2v7CZSHt
lDXiAl4zYI0E0YckFQYXiPkVYzx5X79SvCgz6D+YvdQhZDC+lzDMTPwD+PLZgQ3E
FG32E6ZDxf2HNXaXuRV6+JwqF/8OhfoNgVK+zsP339d5zkbBvO/KnDylsbBGhs91
+XTIMxbAPMHVV/a+DMYum1MyTq+lLIu7xBM9rp22o5yebhElJjoUgaPwWimhWWBZ
wq+RRHyCvd4AHBZBeIf9//aMThEvwQSJbhw+nJP6KPgdQJYxeOKQGJke1gHfRVcr
Gd3RW7iukdk8Ua/iLYAlL8uAH+8tlWf8ihcluPO0yMtmcvwV1K/HbshSCxOo0H6U
BlT+/M+MzcGfKgj8NJZ/VPBLlp+JY4ilZS5mO1QPmHEva4TWzkRcweTT8uD9YR6R
uKDCUHCK+MFCB428V9hllSZE54z4mqhyUGNos1AO4lVJrDlIMI7C75ZSoEyFiik4
JVq8hWJ5xZB55ShWCfPn7dqmOj1IcgRYIijyTL8FJglDwbNjF8fzR2b5E4KM35s2
4KYkai30R0j6+7XoD0FzjG5v1CQZ0C2etPrMawyXl7asdqvGQprYI4DExHn6J2YE
8kfco/NQHQDqdi2z8Ui94fL7wIPCowH6OZyQHkdNiW9QlKh9gz3NYxlE5teW8cRR
dM4q3dKt9daOw3KRu3g6z2w4gQ3Cx3GkwjgJVLhfundtRXTugir9LZv1Pnd86t4D
w8JaCgnhj3XKEzgZdeJLpLWO3bl9bYBiL79OPfXvfvzXENkaVT+7n7S41e5FCE6k
ExLpWIE0Qrtl4q4aOFmlSiUD8T4RxEDmk94ccbFKIsVfp3Y34/3PuZa2lt0ym5BV
yhuhhmgBAx+eGBooNJdwkaLGOg0X4gAx77XTMf/JDkP2XiX3pj4unEcV3sEoiAnG
lMLGeSD3wfVqUAONWbgaNpKcw+gaBXxgP2X4yw4j132eFxIptm2Hv0nrG2ltfO+8
c0EJascl7AtbVacFMJO3QCmmcYL4k9U5DIryIikNLFe7WW5XcjXOkmi5M6ZcK/hk
ZtMw3od/BNoeuCVOoSbsFT36n+yFjYAO2mjmtmK+D4TMO6Nb6ZrRYjo0lwrfmQYm
ZRPM7KEmwoEHuhBYD0AFQmd6Hiu/IELF4mOqJZnUT4kPWiSrjoNXnz4A3gyOmuIB
L4WmDJ+ZVTnBxyUOrGHChFwwIRVTPH1O3b3xd5hvQvuuBxRFTZMSHs094YF1LVFw
q+aAi9RSb6rJ7CU0xaNqV91y8ZweZ1VP1t0tJZvtQbrF/zVWQPNx3XxcWnME1NYW
SuBbJPoi7qj28pTnPo4uFmfpiRZzihW4jpKVmB4lInpYhJW9A9SCEN8UytpMQS4L
A4kB/ZcCDIFjfdG+mztc3jO6D7SBz4D0LThZbdzPC74/TLR2a0YqQ8Jw+EnQpA1y
4KwzDObRs2Y4R2xkMPjma6DulUE9simUFWv3zVQCNxd6xO7GtSKXxWTDRd3zkABv
Ocg8bjdJGXV24YnCZuOGIpiZqblM1jO91YTrHOrrKm40IpEtcKTgpRkLRhmcDCk9
cLqANAxI67fVC/3TkkcuQeznMN8XV9e5eL6oXrIFeCFhDf4VK7vKE6yvsbLLPjKu
irdgeHEqy3PpR+B5leolgUHG8ZdNXC1cnBDMMc82ryLvUN2Kh5j6m9lqexKHeOBV
tqaDirYV/Z0RyLbyZPRXMBlrW+M1cqHu/hKhH4Bysfr85ESm/MBKLZPq94H6DUiB
Si2V7O6SEnY+eiYc3QslwCgZ0jOs0HCv8kwqZgm2oMH4pq0PNtHj2DrUOUthtDBV
fChM3HNtBWUKcyTdpwlvDnNf/+hgwLzZCk9s4OiMgZ3wqm6hvdPLfXF0navbvuYw
aN5sJTP980dyntOn2GtWzxZFyFnZTKUc89WKUxAIiXThRd50bJdmfvamedUctQm+
4grWvkHJL8dQWZDcjAdPhNrirNfzGdVxvdKdj4LI86PMNQZkusvH95tMbi67wJXJ
R2tMkIzRe9XgsU9sEOtwdyPZi0yTg4/kSFFfqEEtvqKttaGj18v33ZIXQpzHen6N
YcBGh7kqZdrQNRPwlaXF2++Fbf6iB+SWQPicXQGDA3dnC7DRj3Qj6H6O3pgeZC9Q
rP+gnedUAXoya3I5KCyfuWa1rEbrceVIA5IGsbu6/3F7z2N4uxqrOgCA2FVUNQdO
zLXv6u+NnXIMADCgWS3XcsoUA9wBWBa/NQZWz5Nr1myehZFOuoU08zDBaVHBA//W
rhRGMby/DKcbIz3SKNJ5rJBpqki9dkTPmJUQH4unOIk7OXUst9gJEJMWkQMpBa16
Sj9ZsBz01Y+R+oGPwxDffK1vRrVpj/aUMwj+piIcobF2ySIw7Ns4iE8fW9TTR2pk
WdKLAZsYsxS1akFrttLQY5H4p4c1VLfIgdsHc4nQDe4d+wntTasJnawXufK5hSEw
wNXkom/OthaqwxdGN4b5IktvdZ2yDsPIBuoeEQo2mfmP549BxAbkhT03JDQ2BviF
HObUwsrK+ktD79rohIdrzsvCMT7niOVGILRFcl6k5Y+HmUUdPGlK8vALZ+PoLrgk
bIqwMbVcu0NFfroInv9mOASiOn6oRZ4+XHB5sGlmt7XKDCPeZevZok2be9LWjbY2
RkL7dJ17xGG9ByhOp65oU7MUi1cccz/iohkGq6r0bfhf/yFp2Ety4mIozTacHvgU
38gADh2xSggpV3GnOGCyw3hHrgfBNfmAZyA4xQD2JaRAP5wZ3qsBu0j0U9Za5oDv
iMmMu12KQBXYIZNf/IMSVIs9tBqOlsjIxA9OSW1tsW0puBu9PPs2TXsywXFd/hH3
wCAHBrsPhaM2hB8v6oU11CoGVc/7Ot8CCMrlFU7vVzR+uyweydIHW5Ihvl3zud/m
TzPJXbGRPAY7tqn70sbyFOKF1NyAiMJvOB7Pg16TsN89S2A+528veovklkX1gfT1
vQ8oKJ7Wx8SiaaKA51yLVy4QsdxRXwf+1LFTMBClUpx8/C7ziZtLSTJPGJF7fvpG
S77pVPF89InCC9Eyl21M8/rmcCMxWh15G7Xizx3yjMjxfz0CqWydZFgIXeBvbcIx
bdrw8mtCEP+CekZBLK9jwg+sg7NFF/kj9EzUeKj1YwFeihqg5aSiWFEk8ZLJDe7k
bJEq+7S3XZ7fGE4pFkrhad/3HsUhTFTdCESB09Vq0OfOeg+cUaNmbSnBm4PTSz9t
FjniyGo092MDUrlXykSxhsoeiTOEFQVDCmi++AYruO8+A9Yh8R7iT+moERKuiTS9
m5uHp199of4o/mN83sLOpUYVYoWLtts3yH4A/1qlXvr/YSh1NWiFSo6lW/6EnZY8
acNlZeHx+dQ1a0NAzoO+RVhqi9E4HI2rKjD4kRwTiZ5OkGZFzVgN/02v09E4ARWy
ZKWJmzTJo7Nc2TomVy+hT7pGkr8/1WgS3+Xer22OiDg8DTWNHVtkFM8CGYVldNx8
eGRSTP2jN279BQpZICgfBoRIvNL+J7AMrRSWsAMvAimoU3IDhRdv0Q8l+oCGX13Y
/3oBww1ii1t+V7L8pAEq2AyUlydu7BH1ARuYEUyn7TkjNFE2Mb8ifTpt52Ht4DQC
RCn6+uSf2bnKtIJKoDmjjnRduLDVbtzd3DOGuKEeqSUXK41Fm9EPpDj0Ex7BPyBt
oz8LgM6OAIu+Yn1LZXcZZPavhZ7may55shmE7KefccP2UlYfPKeOroWm81QBOysU
pa3Pfdy8aC5QgKXwVCWZtHnDL4sp6YESpXxmQEI/k0ssfoGoIf1TVdxaoZDee8IK
qZIlVYorqzoYmsOi4m1BoryKuBSgisf1NYZDTSTwgMDTwol5YzOYVanrOvhXLt+l
C6jBF8VUM6vJZg+FJpO2HqdHrLTK2zKZ7/tJ2URDWzUNHIyjSZRFvqoRJ1voCRQ5
TbvWnKs9Cc4qT3rDYmTDQTJFxdl1o+j9lZlvlVtZ4qBaEwyMFEuh7STS8t91b1RC
hr2Mar4HgwAzu5HzfUkheg3kB1UJlZsbh+ZZSB4bCHJ4k0cP3C0wRgCpBLkWdFdv
a1jGiolfrKkaHh1F/yAk69iigAIqwIXr2lhm6rrDw+lDN1m1AcuzGwkYiJ1FTMO0
w8eIRVtq46D45KSDM+zSVmW5cWA8QOhPMxNxQ5gO+ij9wNz8/8kYfXGGNTQQCuvv
EmOnp9UT/fNGVieJ3CT0T6IfTSX4YtiqTg9DX/sZw2XBxpUleUZw3zMtctOGNuBr
65pKZcXg22ycQ64QXy27KvtK2lDPFIjnsNRtL+pGjU2lwheHScQcWo5rwhgbibF5
GAOyjY1PQXsEtFj1Da1vt2M8wa5aoVyIlHdOWDnEQzXCnBQu2TLOO3YsU7aas7dR
7aH/hFUTD2Q/bYiOKpj8SItOz/3QSU523/8iDn2qPOlmF6ibqPwrwTK9F6gZ2s8s
sOoyU+xPg+NgphitsEyGrNx8x4Y51QLC7u2PbxKngFkGg2GLCfJpRvmpvcqP/Rwb
gCVv+nuI5VQGF+GVcbbMbt8jKfxL5kDz/xmaVQrM35ZAxktEF8DfZHEO0z1tnDji
mxJktoTEGzrsqtHyCyNKRCYkMf6tNEn+1KQY1EnIFjPCWZvtvSMWRA761xIyh8Pv
A2TrKZNlVqXRKys//uq8rZhLTt5ZL9hVRyP2IqxTS2vo8NjnnDGgiF3NuEGGrQGU
cyP2urh3U3Qx7nOFdiP09yEr0RthKQNb00p/cjqOxnOxzEJKgCkUcH24wA5X2evp
YZOLFebaIp+oTmg1UgGoqAi9cFPk5auNo/PzvvNiXddZzDmL3W7MnjVYcgk8fH/l
U32khHu2wNPAiMmMnjLBSS4Ng1YOFstzWj/9JgCrg1V8bKxndinUgaWxAugB0JOl
hvtf5FHqvEkb2BowCd2Zdb20pxMhK26cg/Fxc2DgdXHB5uEttkn4nH+aBjQnk6Ny
TSDYkNtSWxI9QkoKlx7nSPtTr+lgdmu9gohTVg1DcxxlQaAHD3kRYQNx2+eeGl+E
9YRFBmu2gFH2Q2RuqEy07h2Z4i8XUnA49gSJzKehCRjpLZFQK3EqB7QEHQQbiwrY
wGjep33kUkGRfgxpjDeANZpBINZ2N5iivMd+Fh4roBtKNzt5w5N4m9bz76Hlvqvx
sFTHynSpia181AlO/Z6vS1vrfBIoxdACmojhji2LWcDN3b1kf0fB7GdEVM7Ckkda
srejhPXcGLFn8OLyBGYaY/g/6aGBjN3L4f5htVFl/CkPqpF9BNKgmiAf3/Il5bBq
WTwpGQrsWWffHCCXOO49bItz4B4uqZfOm2TTDSj+V+KpHrMHrceqGDgev+5ShgAC
qI2fcS3/Jq16XTExfUG5+l2qY99VVEENueMHPvDj21VVfTh6lBoprEH1LkImr0r/
vUVjKNQXfsLTj9Kpu2UsdEvaVQ6VAD4ze4M3uwSI0dNUq+cG75hL5fwgmetpIc9L
Nu/HRu33mkkAIrQy6RnaheRRnf+3F9eC26l3Waj9Oianex6v9/wt+14LyNocNF6N
vAehIBm7DWqCSlh36MceURZZdBUlyBp+NQC8hm6Lcqe/lqwHXr5hvyqePDajjLoO
+xCGNgc29YyW2XNGX7FP/8Qyb8AQ4Jqr1J6MXs7kgD5y0wAvoUFFcRhI/TfItoRG
rMRGTpwLje3bIvkuV/FK66a3x/mecQbTJrnJBp7DqodNesZgWGSX3qCaZq2FiB+q
U7GYZeAoL4ZAfK7/NWlZTT/TJus2cn19qJyL/+DeWmmvPz0IxrSd5Y4IJLNshMUq
0A8M8TEr7FT4NfwGthgIBewGVDcQypOuKehVk+z9u2iDotPfK+L0uXGdC2ZcI0yV
/2Huc/wOhp3Tzj+if5YSRYv0IXU/1qO3E3T3wKYCfhSwSS/057DFV8aP8xodl9v2
bsjvKME78cmgBZWjwlUeUWUirBBE5F5vdgTWqZkJTqrsB0ERJMXgYM+i8OEkIiE4
g/hcp2vLWMPnAWwrQU1wa3xrMVsAsb9P5KvMMBuKowqSQFKoDmiFMuXj4+tCEpOO
PUGGOGHi9v4gP2OkHG5uXimymNjS4NSteKLVFZh9ck7ZuzYj9ojb+FnYWSO8Bfoj
6rJgKMq908G2KkbqlrH4walB4Q/k43+htMythtNYAu/+hq0S9IrbTb7whUqfxgN+
/xjCHAIC4+aFyzo2f4nZSAC1vNKZtB7gXB12jcY6dd+B59kFUF/u9lGznJMaAorv
fY2gdUGm4fbRcWniiu4zEjps06gIf0ZEwJPySwG9D1hIHVErvJcxi4g6jotJUFJr
nbGR1F5zpfPZCFUHTG9VADZvkYOyf/E5vqb62PW2aqCV1yG/4d34qwx5/Z7Cs51n
9CqRp4WInWSR3l7yn9jrzSzFH6fXQryXtXPhBvxwQijH03Y8Pu620JOdyrlI69vp
kwh/aMAepyOQVgbmKx1wCWGWRp57ZgINfYl9nZ2K9kW4lGqz+tZw+QlITZp5MZ73
idY+vAq6Y17plg/iFDzmSylbjylExW/3XCFYktYdVHn5x4o+cFWep8EfbUQKM9fE
Nj0XtanpMTwkf5qFdEUbfZYjc9zvRDqAuEyJm3DtRk5OypQD51s51hDgto1HcjE/
A7IeTPE6H1r0V3XCAk9JAjnVhCiMopymgYpIQ2UhJtzZAH86tUPS09J1qEjwe8qG
Th7S2GW+sCXP4WNdL1gcIkBifYSPTplPeQbQ9JnN+6/CWI5CekKnfkRocpC3ngv2
yITEPU5dAfqPdOEYt0cXLXBdo9Ob0+20AFQ58Fpub6HIWJzDITxQIL0f5776dlyj
tV88JdClfo6HFZXdHzR5hxyvF3XTLsPKyRUZlF4EyKdV96S3brP7fmUu+S6FuBzv
6LLiRsk001JeFm3Hswz9Uw8ef7ehLnphY1z3pRnLtoGTYvIjza5+VY/sLLVh6JSA
JXfjM6E7vuhDdz+muLugqRldMo6crREUPmOe+b9GeMuiNqiGgeVvk4FcSAzHiWdp
cYLFH8Mfe3cROnvc5YU39OVKqUsU440dnyhqn/4w0SGXZqy1mMDYwbmVahLkZosJ
ikhkhTq8iGxSLAb7xCqYdjPR08kHUXroKYJJ+yYlQE9PyyKJzPXNZifCCfGls7YK
JpfQ7OAcjh3Fxhem1LjzGEMQcodfJI7quC/A7JKUV2uTTYkmVYXg5285H7VAStW7
xSo/oM31L96fqIN8uk4ilbEFV3/tu6QNeqFtFIopre1lfWykXT+d1PZX2Def6JD1
a3KVWTpR5VPI91dGBRd00mkMFV30iXEMCIOk+mAwi7OSNbyVGlK8Iryl4q/4G+vE
Giu6vTPdt0hTM/6FE5rDaGQDH+ECuqjA3j7wm4FCdhJDThRlxzHN3tvTaQx9fmEl
s7Ixl7Aam7/yYJI+fD1S65ElyVrd6HGaughrNwcC8T/uJ7fPWoIKEzS+ygDXyJI1
qDY15UtejmvTcxzXZTIc5eVa2O+VA42vngi25WUOZglWh+scWFzLOEgzyoLsXTXc
59ID5cQMrrBJAAvAOtWVvofjWis9w3DfDbt71pJBXy3ZFUGZzOCHuLM55Ko/ItDO
klEMCFdUZt5EfWKFTO3fQ4ADu7jTzKYtk97RW5dwrMjYwhAQC20VuReoZZVYk7lW
9rrcfjUr41cfKRKD4ObTN+/zn9/OPeR8iwm4KSdhLHyS3rpEjYVhcjfIeik94SHc
F+sIpN7nDL19PWgYp725Rjb4VghkqskzelW3rLRhP21XifEdzNlSCY7biiaoNXF3
n5PJkkGHnuOW2SlSYHseXlSffula8wTbeem9W5Lt+tfTjuKQv4aLZfZfqwBhMWRc
NE3WcRa4adpjo7EpQGYjUbfvpFS4w0Lw9fr56J8cVGUO/1YVLJenP9av3dpLmgNl
Sf7RCSIxVd4r3JQdbdxsckCIyT3LuM8nU+nU2II8wt2V1xj5zhvimerq5aLTJ0Kf
LCxnTB2G2DKGY06bcSQf6C/l4SSDS4WQncN1Eqtz4s2LMQiSQxfvD4KFUqIah1Ic
MN0prPMpvjAhBCFUMazofoSFuIUGW7F3VXWXXtlP4fVlqRYpyTS9pU+d9ds0R4ut
mQvaqyH08ajsZ38f+RbAcTvwv6pRkWw2zd68nMitS9oq6zMGPofHhxY0LmbU313a
OwTx8OI60gSPH4M+Is+FyGhBtXziHyWw14JvEVq5l0SptP2IGPbhWEu765oyhDi1
QTp6EmMjA5x8G+l/CucaQPp4eYchEvdIe9eRFOcjPLFF7u0lHrl8Qa/lzT6W5LbI
4iKBOGwyxTMQzrH0OnkqoYtSsyj2gjbqDLoJU8ITBBCcxoDFrzbHGfR1mrmI5574
12Jtly5r+ScrLrPnhdfC4goh4kGP/r/P1jSyLfhVG+JOwacoCTuLATBQT/cb+OEf
JBcxDTs/FvGbHgMat3C6Py/yE3DxX9HxZ3TqiSIA6yzhOPtZfCvradT2Z2h6JIsw
Q56MXntM2D5LQR9G0eU19ESwqlxtXj4pK0mdqcCZb/UEb5LyKI7I9yAP09J0O5zb
qBR67GCp4Dg0zs0BWr21Jub2IG3Gvu7UJj3S5l+msvWVzjmIzAXQ4psouzFXvh2d
UOTnpnxaV3N5lyfqM7JPFPhYNGuzzEGbq1ACiTI6SajS8B8mArrOcAI6KauuRWUf
euda6G274cv0M/XF2FdL0603ts41uOhZBs3cGIihiXkCUyohy0hkRn1qAXHPFLqa
KZ4+GjFVcSGcnUbWdR7FmoNMwJEoTxDp0yhNG/QOByWOWr9YbA+Q+B/xem5HmnCB
EF0q2wDbKyY146ptTHjsckf9KR3WkxgmVCNZom8t6X8PQ7Y+5bajeugG/rOdVezO
PUTwZWSyWDPTi4OpjnqiPakgauVeFFQE91a7yUCiIqS6vTsW4Q3BZM44Xcg9v6pN
IHb2m63oQXIC57Apq/TyfN6dkRScAJp9UOnCzMLxrP6IVxODdGiOtUaMvVqjeHaf
B3vAJMJYYHXXwW3CrBbTkHTqZDD6j7BZ74p6qf+y7RfN2N79cDcNODxH+jAoxC2/
zf7qbXeiZ0/Amgo4AOKXjZmGzkgOf/KvB5ZCLhdy76ZGkiXKoVsfajPtXT+FRrvG
e1gEOwYqtqCYIJ1A5iMw5kUi/wh3K0WMCGh4n6TpNnMoPSB4St5T/e4oRx+1KnPG
W0TFwOkHTUsWhIYl/3H2U94zjo9aZpxCAYO2TrmWTmH4hqmHdHHNbE5bpJFlHipN
B9zaS2erLGnmzJNYW0R78/vMr5dWZKs8m5Klq+XDytIyGs16u2OB5ud04cqjOur2
t01quMsspPgitxdVgqGibhADA/GGVJr6W9qqbSJ/EY3+SHcrnnKqnee3EbaLvnt5
pDzqSnQN7BFbY3fSxEMSwuGiRaIxVEBTFxLyjRrayy3J+oeK5fGC+/DeibkbjchP
LX60ejo3r9lBs+F0sPFiIV3bm8tmi0OaQ3ThzdyMVc+j3Oz81s9cEqyti5sXxFb0
49Yj6v3dNVlUD5lw0kNRuEzILt6GGj6fAFhsZhca+b7EGnzbFFtouUkOIwYIq6zc
YNYMy1YG8fLzD0TxXJqYZ7XrGsjkf0bx5Bvfrras8cAF1Y5eL3i45NAwSmT6pDxM
mxokbPy8HsrFEvMs0W5UUrvhKX1S+RNIOoY80GRt8NHsKg0sAmx9WfjPwWAXy2sw
+D0qmuqZeKOlVO9u4MtAKBCM735tARTSDAz25ccBTUI+y568RK4aQW1GE2jdTElH
+8+Cqa67bYEx+iLqHv3hmd71C9uKv4Lw/x6cRIaZR4WvS26VbizLEmzrqQL8o0UP
pPm99G0WyUnpSSyxuvBBkEI4Bv+FSKomkXr6j85G5hMYA19cBCTfLp9eh8SqKCfk
qoUBZXJ4yj+jV6QG498qyGSXSN8WgMwxwRsP7Bh5z6PmYgTEJYqOVzw9HfGw3Tt2
IYbUD7Cs710RaYYt6atMbfqGsIrkEwl9iSEyPlJQVp1/0DhPpqLbSLooH7kzouwb
cCqy1X8Bew+2/pMMw4qm2Yv0Zl/ydSntxJzGIOjLVOO/xEjV61MdDa1TD8gfRbOP
sWIXbeLu6kYsRAa+lWtb2CLbd9gdDRFY2KUFPUnpy1aRYIKLQYY3/wT/fla/6AUb
ybm6drQTRL6lD3bxhxMTzqyBrjb5QnTBy8QVvR8Ym+s/DDCTKqYKDtxb+P0BVrsM
tz09KzutI4GW/C/2ScvpgylEsiZumDITvwaLIuH78LqHyrL1JsOmbW8TZ17lbuXv
poXIPtxCEMYDRopQVuen6WpTrogcsUFmxrpQKKkus5s0Q3QGGmyLChA3FkL+QdUm
6WQnRzqRiaxf9B6GeoIBgBzpsN9UPLS2Lb/lCroNlF+FtahV7zi3HKLNNsWwvUNx
alVlAU6K9WLj7Eu4vkCL7c8baR79UK0e7VOD/ZCnl5Y+jQz5hyTvzSg5YgrCksXr
M1feSPUueXgHXntZskLgIxdbwn1C3ATL3goVcrxaQmLh/8+UwaqsBVI7KYnTZiYY
5c7BtF9vfeooB1am4VHAg00bTD6FBx1bGpDgH3JKYhN5nroEomGreyYdlpvdkZCz
sSJRdF7beLjX45b7paXnltY6ez4sa5aG5hsUyD8G9Sb5eNrAARvaWRsmQ/IWm+B3
+RWVTB+q9tY3W3/jF8ay+Qv7gTgNi384eysOMih1/QQ+o0pJKZI72jroDOadzk14
fVvRwnnp2p8W4XrGGTMFwuGC0nWEa4aiiuyiC8iQ92XQXj+BYdwzOrvevJewVKLj
SVuco8i77rkXLjpFCAdzxaUifsA87wtQJuG0dkJ+JflkvnopIgUIQ8Fb+HaThwEw
LAJMQrmowncvjGbfecIpok2Zlppx//c/DPAta39tfyqAjZB7KpWdPwX7jDsWpMaG
lE4I/ik9cSz5H1+YovWnUrIkfLIFVidaWuE5GPXrRx6tA4V3mbqSuiSMgvFkdOOo
1BgTc2YDU2z6k2vhir3DBEJzt4Igjfkz+KXUP1MGWwB55RRmcilB0D87ld+AdwAp
Fw0x3mzQlglQMK7UQQjQHT+cU2IfKKBe60W1oeeC0fnNHC/LEaFzy3fDXda5hqNw
FPcAGcoI6unMQ16HYPgc8VfKR4SJDu0h2irpN0Y8fZGLtYLuf8RFGak4IQn9BxCG
g22StxlTbtwKGKMK5KyIPk1KEjwTzZF40kX+H+Gh6M5Jf3dURjmGdQ775n53F18K
DadytSX2WJ4Er7KgJz0D1CXwDOlgiUTLJe6Ly+DMrGjfeGVq+GSdRp0ah5AQb6DD
lxz+mE06sXTNzp1dLKpDDZP5qiiIBNZK9kt0g2RPo4OJBxzKFQfPzMhTZqPhKUbO
aPLyk4GLlsWR7QiPMAo4gNeC8xGabGQuH0oYDZRIgWlSIF2Q4jtjFfLO17TKqF81
DmJHVDEkgUhb+ylg8CzvuWBjlvgfSzOvUTpOFdJip5JSkvDkJ+WBqh3pLx96FzPO
aBS7WJdoi++C3wI2zDwUY1b1AjBXp4DyQ6kT9+QbnZ/qa3lpsbrFOUCfNlqc6Atm
6hSlnfxX3N3W3PMEwLIK3VD0K3M9GCCcgjS+lmD6hpu9D1DnA1N8N7BBr86+BRB1
Ujq8K7treEQfIqAkaFlOpd5WpW4yZNhWIZYYASQe760QfX/ifcxzCyHaL2IquE/p
ekCPngqmx4FAHy+zzg4yodLFbr+wZcfufS+o5+pZ59QlCzMrvHxCOd5Jm/6AVzsB
j9Ggcbq4EMI6L37XkYAwBFvKVLXhrJexFJSe8Bk3pUemd9AAopfaxp3ujehmGjZy
Jv1OAXf51Cl6aR/h3NjLMF31Kwu26birZg7lhn58effeBLnS+5SxuNvIAPdu/R/y
LZDEg2vPApnxVDV1oUBY+OD4QTitg0fvrnqfeHA5DR6Pzz0az2viRv0WL6xiHiGU
0StrndqbXNQu0TAEuGYprynzA7rt8M5PqdLCojDwE9DVBrSPFydJL4gcvyY3etWI
c96TUJ8pVDoVBGzHr8Z21dS6fQdm5/5sY0fkTFYh9zLVkOX5irpH/aUyqMNsn0ww
1qBgzfqZDgxWGiI/0G3SGG1irZx38sMlMw0QX7AugS9lu9oscEJhz2ZWJpjpvFNu
pZve1fC0OgwUbXLQc4uGn9d3U5yQwTuGPN+c384djIx+ZVy1IuzQ3VKG2g9D9jOt
vCfdQTauE5e6S+NHMMfgoVY4ZweMJ65Eu/spG6wzDtTnz3n5F8qyH6++iPgqd98z
D93z3KocW6sktX6PrurG2ogs32Vn3Qvtz0o/VV+bucqN1nGTWSJByRvT33o+jEkx
ZzlJxs/e2d3rdnJfuOG91n05TvJ7a4pk2TkqBUWaK7ey37Huy3I5rQvIkZi/GZpb
8MEP1/1Skyw7dslhuUIhWEdFdBvsLVTglx5EJIsYzMGHq2DibRXO/ptxqEynZ2/x
/wx7URk/b4Hz4gtZPH1JNDXN+g1hfb2Jfsi6Mjrzjhm0glQs3sEaXyuLfIfhrJ6s
8Y+NhgLS7mN9sECKHMthDnK1Deo+OY92axNF3UdEtbfaBZ9mlwuUf+109gJUBURC
hJUEnTkVH601zTu54iZQu9F7xZeCgAZTDi+hhfJFPYUGiep9sJcKBLohLdDtHvO2
EafO1Cvn1aAX9EeoMDhG3SYqxfiCplhx71C2rZRU4Y4rRASfS2/gVGc7Um0ZYGxo
RhN7we19AOiFAL0cTrHlBq6h0ED42SaahFr+/bxRIJQT5c/3YY/lO9YJF7uVYLwH
H5GHQhduAjj51HKLuqor1ZJMlVel8QPt8HPEU4Q8Tfh+yNUpYs+/I5+lZCbGcWP0
3/rZiXc1jJji9gUTgnprbPOdBHNgC+XA9nmLrxe5n3j9hDXdrxl7AzAP6Zrgm9Eg
2ciiBxsVgA/VhNytHqnRrheSJpqBUxRuFewple77mlsz1MoAPcqVH1zRA7Uh7AGN
RoSw7sjojtU2fuHMRGkO9OQ5V0xE6mQbC3ES0GAYeyuqx+NLeYpJHHpAFCga+wL+
aBEAA/MCbM2UXe4Zfyb4J5KZ9eTwNpYegXzfK6A5+4WUTBMaMQNxdrr1XqSN+/YG
whmM7VH410CsrBFbYLjCz33xj3my5JJ3HHrfHOzrmJpDjRTa0kfba5A7KwB4N8np
j5EqFJ+RwLHmAnQAGP7IXPxA5s4wZXA8KXgv5Xdi5Vh28BdDtPOqB1Tzezdff0Ik
ZRnsRQag+2olBG7f7hwN3VKlhtQNUzFSpXyyuyO1m4pKX7TfDj1Jy5RJju7pReu1
zy/+56o5n9UbXVMIXBe6fXzXWnhRkDc5eQqlW8W+vCDhpWlc1TFyRZF9rrrqLXDA
Be8T+CI13DRjNQ61sE6zCHPXgYJViTn8VA973SnesMZ5Xx56NO/Ildy3T+lw6/FA
OBYsu6LsTcMmlVyKBrjm3cnM/43YjSDzvTyPLEMA7zpgG7XOLgg1t4ASXDEqxopZ
iqu6b3fcGyFkDLuDP/+jlZEYp3RClLv8TDs1vuDjB/Nr1lulS6IG4u1GsVCo19WJ
LqxcnTWfdhgjgaFOtKaVyBN26y/yJpllmUeK2skyazFRFaGQzPlqvIYzHBbDR9Am
wylkPS/eih64NZFKardxNENLtKOUqQzMT4ZOG9WbvtaVw9Bw8onhUW18SbgtH46W
JTLZPZGjtfnI8I2xcGhgzMo0sAv9QZWVli6LLiTqwfma/HCcUs8i5lt7BENM1+gW
b/iMHG8OTmA33KlMSTRoOkdzdn9Ggn6F7f+BeueUmi3vmxLHYTLuEAQdGZ0jMgBD
aY+lons8Bm/rZVVlCk5cosm4jpk46BXXMAui/LJFX9G08uvgfQ0LgPgtpnBqY2xC
Qcfby62e110vJxMM99NbFOqn4guFIHYdw3JEQ9G4v8a3CT16HCN0qNZ1gaNyN/2E
bWkgziQ0HBSIku9McXwsBz1+gMESMOJWM2gh/gEpmgGzPQ5PPFD7RrGZB+HQ/+EQ
+eWmK2xaDHqeuTbCqiIvYy8x9q/8RY5eODrhuOpFxwWMQpgWKn7+5tdKligpmXBB
z95DqsUvZy5xM0Qafq9mlI8xhyI+vsmnvjkfC1qAAVgBzmUUBzdXJ6VscTjyeP4P
1Qv+Ie2itWu1b4Y6eEOIaML/CrUrHIBM3Znc2PiHQQ9yt/TEXsk2xY4IH+B4MQ3L
RnrmTn7pyE0u8wuAvl4YA9te9lBkjJ13YjkNiFl6I9vukht4IQN6GOTeWskn0U8A
hfG7jvkHZwejzlfFUI+NVAUZ0X1FA4bKGWjDVSqbEtOZwLch0XKJbpV/fRSvfZTS
TBVM2u3Ol0MOdBRpTiOD03Ktg2+TsmXwJj4jxUB+qzsuFwjY1Wjdl6Kv2jLawrcq
/m4mxm7b8xK6layOAADcs9jTgFl01QWE55cZblbyPEkw2UOfMZAoeVPTRqOgPxWW
PzAjigz9tHlTwWe8wxtdLW+HQjvHF3aFrdQHg2EbPJewk+CHEK51MEW1alMDk+PP
usNFwIclFOmX8P4u+ORM5sY4J7Cr2d/UJ3Fk1e+rThYedq2ShkluRXM2mHCypWD2
nAkIVoTjGgltH7kD4pTsZfeRJl2zvyAXDn2rbaC+VIfNb4ZgW6e8YiNfiggYTvFJ
0zhfFNLSuVVJFR+xfpV2gc3vHvhM3i9a5MjFvwcOUZiPLq96RaO5tObjZNq3Ovdf
paja29irqux6UJqSAATksrixPl3ndMFW0JQ8bPZT+G6Qmu3fRrPQIN5cfqPzrsLL
7eB83movPIoRlHYXUvwjTUo0Gtzc8jXbywXyTHbEVbsG4eQwOghIX4sF/Y2JnUSH
DwNCGiewytN4DPcE9TzsH9GEGdkfSyjTlGqFlWv9mo/IwqjCNK6164aUXElPH+X7
O26uxIKSk4uUyBdaFMWuA8fza42FaanBQmZCe26EI+KbuU9d2MeheeA2cBqnTYwC
DmKTkX+N/pWjUTWqos9xM1OMB6U9eZkGXyXGeqa1yPJ0MdEeG1PL5GumniZe5KoN
OP0qfQyKUjsDsIbV/gTNa33eZkhP1SMv0v5PtTeFzUtk0jkC+sGt6FUGMRz6qzY6
0bcyYPSnEcLRrlhDapI3hSEpVST3arg5nu+mQ9oELJVLApQoT1imeBERL44EDS7z
TU1+q7qwX8px0HC7Q3/F+9lLcQMmZzjlGzml0n05cF2CxHP2Xngk85iqdJ0DE8Qv
7MDfbdCDv7SE2S/YgT9x47YnyA5TUulZzU5yzxfAB9AO9W5GSD/TfhnrAamvgAUr
Lyc3Yj953rmwu3u889b6r2ffgW02Y8fssZQr7wOgPclfHDhL5WvYseiZZnLdgX/Z
6lK/4XiAIwzcI4Sj7t6tHHsosmyTjqaPnLbDqA6aXn+Gj9q24h+hxX1muBnDNhLk
yFR/Zp1I2LdbOmW5uEdx4OKY6vsvs2EiUz82QLX9ItdflW3cPPrgniP3Ek9NB4mK
pN3D5er0zALLg0PU3fKH1eKGByRBg4+v1JpNRokCp+J7r3iuD28IeSNkmPuns2Ql
v1CCFy54BWNk6Zr28SxU1Wk2p6MaWVw/Y5ruYfIY98W49xQjBLXs5tld6MrwUDMD
Xr6taZxCDyyxazehsZM3p7DQoDqiLRJskAJP8kNn8+klLTHmp+/8Y/Fzovs2/F9C
OWMQ+COkDZIfyEkYwgD8vzAsfOE0KBqz92GZf5ZUhgk/ZshzOBbd6zHYROfB9r/2
S6Cxpj3cIj+q2sS4zxW7XJLYblxQVrGvet/0csRcLYBYAKPv/B9BGKZ3NatLd5Pg
x77DF9P8qV+PjN88O9ACPfASMlWD7siA6pefMA/SpVHJu/LE6PmPH0XIBRAoRgKg
H53V6YPAG1XZ48dGLSp5mjDR1MUdX2bQZGSXTI4S4NCy2CNGaGQ+UjDi45z+7rZ1
wWqsqrbTUORSfPGoskeMo+8rLdbBz5hdIlEmIh6yt7VzPaBmU0hxSRE7HKF3t+BI
Y0pcfPeYpJfy5nfyOUz+t4eE1Ms/WK+Dol/L8S+SZ9Bdg32tVXn6Y2VeZ+EZQkiQ
dTY8J0DTvSxLYHC6UYjuzC8XxooqiJT1sf0GRF44KzIuEDgsfcc2s/HnqkaOVx9v
kX/Mk0rTrPlqeNS+pWbDBbRVNwuB9dlnthtTA2PhtlGgWe+a64yIEdoMQDilhKdc
qviorugHU8a7n3C4uA5yizd7OqkRXW6W/JHyXI84GMZeJqmcwWBjNt2qGNl5lR5C
QqmtKcKoa/4djgRm9d4ugvEGt+9yWsxhg3v9uCnvnxS+bIRzGDMZMaX1LJQh77EA
U25a6eDTeNUls7+QQMkD08CuYUWFXpSxxaYk0bZBt53EECxcaT5ypHE0l1DYVcqj
MaL7aFpEaQrFFwJPGQixhBugWGPYaY5DML0sbVHLnKCJ3WIPi8ziaRfce7ufI/L3
vE68PVQK8l0ynWgdUApTdbJqnmG2hPOHVZzLmKsweNXtKc2Y7bYNQBde5HdVByuP
Y1QVNXV9jfd1xA0cum1l1KuN5KVaaLmXzL4DzXPgt+02bEhREBCnuGXUAVdw9H1T
fuYfR1TBi+vz54043oLWgW5NA6VKhixtZC/ZpGMTk1FYNsAG0hCdhxYdPrxJ9nmK
iJrdYLEe1mpGUrHVDC8LantsxiPNCcaheKimUMa8xtlxFKi03KKe0Uj35sLpnBdq
fJ1LctvW28E93co6nX/ONkfvomJjjkLzILE+2ZmxRMx120aZV81QHzhypAaldpRL
jzYUaDTx7oeYEJRTLivqNcW2uC9c5fNqOgWE6BPRUJFuc8fp7vcdGeBBMRqonwi8
T/M+FcMdduBo4lExsRlz06CZgTIbDVLyPCWAqDPYfm0w7qfTUuNleOdWExRESTTC
NLIJImeVZDtUUt1b5l1XkH4ALR9acpWALDlGUVfAJE7fQ9sahrw5E9qINSz+I4Ae
r236FSgpazd17wsDDJ1bJAKc305pjUUirocLGu51I1L3hC42hEQBzd5AN0Qd1WZa
zh9cr7pcJciAG6UbsU2IkixHDW7ct1zkLB69xjRmNKx9Wt3+YLSblKdCwq4RkByP
T2u8SFYaEuRpcNSflm4GJ0H0Fto1K3iaQEUdRMovZzYTDQlQGKxAiEPVYL1eBWLl
JQD8AvFyIVagBKIRSbK4ueq2BDFAz9vvaPJIid8Z9HWzzPRRs0x47EUK1BMHsR76
YxuKScF4ZL3wFlXzGvjk8aQIXdyTk3VmIbOM0Z/R6Y5BiloHlWJcaaLeeGLdccwd
kmfF9Onf0CEunHn8U+aaMoBnlVMJKMkYikq33J9BwhApeHA5775wZCubsfWvmqNB
MQsFNygBOfw1jYmuvE8ZwrzBZu+UuO1zdByili0RsulNuWZ1AYx/5ITPCr00Q0Pl
eBH/iGQa2kxvRPDUX41VZb+MEKrnpb4X3lxWNEYwVT5pppIQzAugu9gOUzDIr8o8
juLROcoUgGCVjuXq2ajqfNPBIrPtNwq213sQMGYXTTooVgNlasBGo+sKwmUtglhg
Zmm5E8QjuAsO7YP/UhOHHMd3Er6M7Pec4hVUge98+0SJfOXK38OFnomJlTpMezba
q71m9BsaVDm4qkhWWfX4Zh11nDC8oE675qhFUugnqWdJJA4vSwWoWKgU8d/gHsT/
e5jMVYDpr8saUwa43oRY/Ww9p81/SW9EuApgp+fo/2SWKkGO6mW7DJuOHbNE4H/n
oSRm/2+dIFKbBosUmdDMQ07zOldVoAzqkHcONa3T3hE10JAzy+FAPN1SRpa2gK+Y
4ktiLFIP89ftLnpz6128aibHjmyBHGGz5KjlvoIC/8SQnP51oa4pvrVPdoMkWfIa
TfTdiq6G/wB0V+MjU63LwI2sNrS/Ks+m8ve3JZE62zqEcbnP6Lp/69pKt9W3XT83
2WYesApDXP7NOSitEDZsgtuFBbiWw043iaQOcdSI3Q/sNyj/3lmlExYDG95gi2oi
ktMJDP8Ycog36/F3Pq1FzqfQBiCbPAZcHSI+Xd4UGasaObxHlh6DCxj/bjOkRgGX
txUV24YQL0/bR71hSzotC9cNrbYLEnH/kC78wY8GZxdpNS4y9UUQdIxujzRwnR6h
rlcIX5UzdPtuMIF9eiF1SA==
>>>>>>> main
`protect end_protected