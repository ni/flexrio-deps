`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23952 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRpcw2zQDHRgJxPf7yaQH79I8iZ3MaMca/r3UWOgJzbEb
4ka0j9adKevpK05p/oCzxAS33moAGJjJkT37KVTM5vas8mX7VkqSjFJMYUl+fka4
WRdIC/iPul/FdUMudb7ykTQPwTQexEDOyTnkdezvbDnTUx/+B6SBSj+oLpKD8v9o
VklXggyQZYIK8DBELA+HDao1h3ATNRyUeeosk2BaS5hbmzfLHNHW13fxMalSJ5pg
j9BOXXSWIMyZZQb7e3jBeEV8Vyrptawquod9TdE0pmh4vD6JHSdjjXPv01oq1ija
8Vtv075gmD/fCl70eEHc5tLQPmvuDBpjTzbs9WRFkcYKpSh01UXE3Mf8VZ698xXA
MxFt0iu5//8kdMeR0tb7sUaegdya8jaCuuwmYOg/oxV4WYXr0OPb7R4xUxPA9Av4
4JHY0htC0Jh5LhIBuvD7c6uK30pR3tXV0EG7FAE8qMPcedc65wbXEqyFNpl+oi9S
umRCqmHfdwFMrnWZ0dPBTC+4qZsN43YXeRjtHfWm3vSqkWCECWGoHaO8PaiGDxqb
E2jARP2EisnFE8FXA/vT+3ICq2UXCaly+JYfgeOfXCsQ3Uj2nytuZqrteQKs5l/H
vUXd+iGs/K2JOSPoX5YAlXkV2bYG+f4dvsAdmvQIWtYkKMkhgn+EbS9D/4NXpPrr
hePT4haaGMrpBmlXIAvPhfP5pRZIN0quObULsOhgxosunz2VwJRm4svWnAEfZidk
dSC2Jd92ci0uLp6ElXq5UsrdmDd3vGoRqHnILQLHsd/NgPV785pHk3JEpQb3sr33
/HAMIdVv3y3BqIpS3k3fIFQU3B+nX94vTZ9t1ELjWbrCdOWzTZYlPrBIft/TWIkA
026N9/MunkclKm+nUU87YRD0WjqlEIca7lTIsGlVh6LPWgcyyB6HTKbwNBvcgCIZ
kEl0GWvYIPFv3zpPeP7qp4QWONFH2rEggheD41qrN+AQe+ks4bRM3IYu0Q9XvCRL
297JLkkOs4j6jZj7xuwrnAbfvgIISRKObFtwknrD2oW8rCmisYz3j3uWwnu7+vyh
xgjmHScvnyJ8zz2UgZp3ugmAm0OnGLK4QprozNvHQZj093x5uY06V2U8LKQO408t
Aj7P3horwFaC3p3EBGiekD+BIzhJ383aHSSH/+x3VZYd7+e7AEjtPDkbw5r4mV57
yaS6xkglYFy8CZPvG8UAJKJn4Fzm5JUqqXtXvZZ9e2ETMKoC7ucIC1fl3G5kWAbA
srmrENKW0yMuxz82hBn4aTAdvzRAS4XZpSuOjSc4v7Ehi8JZoOC6+WPMOy/vWoDy
eGbdWEoMz3lhhge96kiESMu0sdOWbe2keLvIDZ5d4pkQquQfJVKEiU0bXA3BYWlv
MWc5FGocAeOKxTYKIUEMXmX45dcF0L1y/3qCNdw8tPN3U7ohw/u2azOoJrGQnxKu
QhF8hiaNs6mpiwq0IinsO7a74OQHZiKCOGgaxwKW89cwal8NPxfHwHjG4KkAcQ3x
3Zu+U/T68IGtpcj8uPLy+1qOmHTFZio0Fvm5ufJ8ew0bUBvzwTpCpID9hkL/XEoV
7LV1af0xBk4ad0I4EANMKvnTqTh6GMWDfjTj7zFanUu27pTz/nm+NCHr2Yc3kNpL
MR8HQDu/7Q8BqO5bPxbsZxkuwekDmdxYvCxvlgwEi8lgh0o4VudhewCmzFyG7cAu
sBQ+8EhxaiL59Ajuj3b0XuWHnN5y4228bdnEGVf30jdafjl73R5yYJJmnrB5uhVk
uW6nAHGBFvQ9cfLO8hg0NlMqeBMjzcy2l5ZgEFyMzWh5wSww0Qqs2G3Eu+/lT34T
4yndlXa+EfIOyGDURbi2nDek5iOOVgGQ5gSnry7thyGQ9Gu4WjbMXtWJZGTOSTHO
Lj+XxuroOweRe7nXLB2wI79QF7zWKEX1DMnZzUD7RWekUm2d28vt/gBuxwtbtbFE
/jcMIFfZHUK9WrAltBogf4IxxbQPjGyiNpOfp/g8AkeP6dZsaEGGpCfOQCTQ58r5
JUSk1j4FkUSPgAhzc1Ek4skspDKYzJ3uD7ipcxOH6mKxZZGaqBxRjoQ5G6L/fGkz
ijpE0zZCKdnxtJ4/5pZrJyTiOvuC5f4ypuMps68GgLRErml0oxF3SjnL82Nwmn6u
GMp+ztXm/5IUtdaj8ngxR53mvdHns6xJ7Bxb0psTB5/1kJd+hgdLwdf5WI/FAHDm
GXr7xJLT5rGfEWiYyRU1TkSTHg9QC5BWuZ9gk9uSaSCsgcAm5n6S1eOkGOcfGgmU
PTHl2I/E7HWqHygtlNDMbLLP0bW8Ezw/JVzUebVwBP+btC9VHK4uxWqI/zEDFf3C
AXBnlG0s1cUzvxKQ5jPlYAMMrEAMktXU2D1SqYncaBj7b2bIooJpMcUF11OaXjr6
OnA8Pk41f0qN9LZdIdta8uWzZ/Zo+YFF9U85NZm3t03hxG6EPuLIJsIPQwJzHX7S
ULlKX6qGdb/c7StuXUU+eFgnaQj7Rl5VMhJfi8pAUlED2U6sMfXhz6QhQ28aR1G0
Gq8Rs28lEgJxf2zGEPtLmkLdNrzqOTD/JYCGj23IZJRriFJkcE0BrWIE+tibR8ZR
N863v3rvkGCfEd+q8wgATXgaN2JT9G64KSHLpu1MN47sNxnxrQ/7u6NQDaEke3+d
fYhu9Rs0RIJp7VSw5gVPt3SUr7GAA3Ngay7XvRPrS3sC0ApDAdSmcA3ThpFIQMgp
xbiEx9ddG3Ib5no2uWnZiJW2rSiLdt/JbIvDtvV8QTA0RgWG2+HXY6jZJHz7JFOl
yUPN/Iv5OEJq5l+Og1ENi2YCv8thkbn+8B9cCJ8rP5UvsYcvLwsYvgjuTsutADki
EUimwCoNOyTTI2CI0LJc1+xdydax9ocA9achp8yj7LFIq0d4mxoR0rh7s3kGy/Xi
dPAZ/6QOlJPPuQaeE2OlruDvv9pqlzvairDdiGFRKGA7EAvTzzNgd/6Xr927VFCA
SZZAIcbKRpX6IcO1IcShXM4H1Dy2Fbcd2gDqA9h2Phc+GzbDiusOwESjmFAebcNP
jbOVokZed3OcYDXTNFN5r9S6Hr4GLVsqsplLlP6/JyTCN1X4kIxFE05VFrdci8a0
DMIteEXTwNf+xGTzK0iH+c0HeBMQHmN2+l7dRcdTCtB6f5VQXqd/D9oumNuJ8lVH
l+UaiCTUgo5ZbcQ8K8n62ZVmCRaX7F55SYEUFBFnKP14HAPKkW4ocuYst8ktNE89
ylJWobhda/Qpra0SYQRzdswCHUa1SOL/IbzzhVWt92nZmtK5HpdPB6BNGuYzOJ4E
h6RfUD0G1pCNRaqT4AkZJJqr3iXB1piEZ8DMM1bzn0kLVEGlBIh6TcVKadmKeQNm
Jb6WEpzN9APKfIYCHMNctTjnLroQDgvLgURikdMNBavYkMM5rauq5XKlziNFpzTO
5Iw42JRU0WB/bCdrkLy3bHFsVj+BbB/TOP0C0A1IvkI1KC1sepUC6Sv87reN8gUV
uIism3NO8wO0SrohAcNaZ+w3gx0UvRp1tUVAFqX3egzMUCqVvyMav9cOb0Ed6znQ
4H9QEM8NYccPaJJ6Ai3xMD18P/7f6Rv8l9b3oxxcFcpSUbOXfiULG+qSnPgs9KG+
YIyd/dsnqKZSunS5wEJK/T69S0Y26w7eY7YqH+LY9lgIwcD74QgpGAOlmuSvacBy
HQ4cugwErJKTNEFq9vaF0dDA/zcyY90FC6oneTyMY2B21mkHM6UQDwsbWLX94aLZ
xScTR/qTXHmKQ+w5sXwtljZRr4fVed08YIg3iKQ1SwiSoqTnzpAeCSMH0mUVwCSW
tYq309bNMwlQEl+N39axUO5mrcPMFA4yc0zxGyDJyxUNTPwJpZEB5aw7JYmQexUl
kcYnggLRoGx651Ie0HQdLbmQV8BrYAa2X1f++5koy6EgVpenKvCZZ1LnuzI9X9dq
1db74cpz5Mst/9goW6R38YGo3EtgvV2gO2yMizoNw1Pc06SARuOx9P0G6YBy8p05
sanRR6QH0mrchF2zRHU8JRTzv0txVsdT2PBDBb/S5qteUNq/f65tXOTpmKJdEWcO
0cm5gYeUTdnhXJoYDTP2fwuOydD24A5bL7L7Z3KZzXfs2klUSW/L1RBmIhvneleZ
8D9lqEiaH9nKAMYbgawyB4pNQKsJe+QUYdDzprTurNJrvtbWJO0tqRMy5WU+RVpL
otN4LkRCKdkC/JCjbJU0eibfM3sxca3hZkeA6onwSUNZHCwUmG/X301W49vAo0jo
fyYCUC9Gh/m9wb40F35+dVY2acwg7l0mRV6JoP2G2nGfoZl1xH9i0JCQXX3AcShn
8PJ3hhBlWnUoHTM8H6Ze1tmltRvjUjPAORVJa3pqTEOthD7ZzJ8BiJ9MSEJrAUNB
ZvCzkuVOPmLujnjKmlpt2PnBidPmShn+jAhYNFGbIXuYt2VCw0D3ZRiF2bOKpqCs
0k7AGThS4F6KFg844Q6ukzawYH6h+TkNcFY/hy8mVvY8b9grAQaA6crCi9siWJmh
ctaSF1KzBJoHIveaXvuj767p14+KMttqP3ftT2yfNbaYV46BBtkUzdIfFG675xzf
S5Is6cyPpMAuX0Iriuv2SL/cVZttU9Pto1VCj8U4+Y1lMFJtpabCz/waQ8kPi0LD
BngJgdIpkueYkGlWNyMvP3B/GhbWfU1yxsl4QZ1lvSutjuwc9NRIW1yBoYuO987p
RA0OGW/hQradHJnQz1oLxqk3SYDj49vkwp0+AEvWTdIZEJ97GkTMBjgnKl+atr6J
gcwHuce3/1XlJBLqzqBwh4cVAq80SljjpmuBxFmccc7o8jDt6Du5Wc5o75+061TU
Ox3FUoDoYE6Py+4g6FESl9d0U+XLv7I53dfz94gj3w3h3gl4/+RmEVrddjFb1ChJ
WDmnuwnx+bkVPs7s5kj4xBZcVst/6EHgE5VZh4Gb+0THTkEtLziOlPzerAapRAlp
qhCQrX7OlAbwDYnORKaRNC1DB0w65pwdYvp2vCm+b8ZwrIG4orN8KR/nr01siDjX
UEWozgsTMqS1KTHWJvGgcBO/ruWr4uxc7x0ToRHWhkYCObHXsoUoPM7T4e4g/dZ4
2woqjfrtCE93PrYiTuBlEcvRezgori6ZSxuyeDqUvIs+4Qr86zvwI5R6cRV9396t
cSvNbmhBnY7dnZ/JjAkOWMf2GLtAlhYpRRD2Q3HYKjYvMJ9r125zUkrYsghpILAc
X/OuqqAy5lPZZFibL6bg17l5QXrGSzfB03B8KZgIVN7Ly8+CajiGKPq+1FBhUZA/
uBJ/g6ntkHlfEFySBb5/A3LeRdoyUenF34AGmO6Judwf9gnjfmuJcbHrty9CEVha
hS0pezT9oyOYhJ4Nsi6Axqfpv+OVof+iX7Eo3Hn9rTZmzOQLMYO/C0Iehfv1wjYq
i2HitDf9h83doJ2qAssmW1ou+eas/7BpIrP1qHhUtr6LAThX2F7oY83ILmo4IPxP
1HKDvCLKVU9+JypOyuDp+uhCGsW5uuXEr62Jqrl1X57Cn4euCKbCq6spUXMAIlOw
RmY8FX9YcdTzJS9qlXPzR32eFEZVkD3qS834ErNRiRY83s1CzcCUpnpBIk0jhiN3
uiHEcbYfIMFAhBTcP+zELBDpXqtZQolDxBGf0pnp20xo1mklJ38SaBuHWC1GrqH7
OzxRyOAJZbR7IF+sajNDswv/McpBRvGFFZ1a+x5fLrvHowcm/Bi7HPxl9sQNegN0
tJIn3auuZgvUyOBjZQpjazoevs0jWDGzuEnQ24RpCITPOHFgG9Q50tlEe1PTNZK8
x9QXuyjG3FcKAlSBGgPrdiydox3dgX89TBSrSr/KD8yp6SMrK5cgcc+u5OexnLI+
iek6ZjE2RblvyYo4EYV/PXEJ2J62Otp/FNxmHGNnQor3xifl72uXl4zcgKvFypie
GOasHeI086RTNZd/rN/N40t+HGLoWazfAU7aeHdmZRrCIokqVm4AlOKWaaYCyTgu
SM3UnFNsSUw2Wo14D59nRx0cTYxZC1mAoA7XCSH7DgCZ0gU3/RdbRSkoa36QHhIY
idHDMLKrEAawG/rrrqGkCuYpzA+V7LGtMZjxdrk4/14WLwNtWr0m9E4QgudP6GPa
eBfTaTYYYWTsOovc4/uw612gWtY6vvrrhY39L9/kSWW18qcGjtzeco1mD6gyMlQc
zr0p7L9XNyOeyvF+RU3xE047/1QdV0xeFViG6axixd0b+xrIHBkyHhmJEiPxNKLS
GZgIwdtHlDpF3Cc6EFwGCVyZptoM9Ji2qOILc9/ucz/LbVp0wVe6m+0zlSS88G9s
eZeG2eMVZmlgnACVcZYermbP/JlkFGM8bDLBPF/ELclHF2nX05aej2cgfdJSmG57
TDhs6rV/PU0R69MvgCQ2oKYsDCNcUk4mxhRpSHmT4Q0iHmfRItKVdzwOY1Zwb/Y9
Bh1UNV3yIH6eqZhtqbSukhZ+ggExmIWSVK3inECfiwshMIH4QfUlypxK0kpCMK5Q
fuCf9t4eKwB6L9AGMD7yE7w8DJaEgyiv7ySsSN3B1GUHJ5+5/yrIm9KA9eBBtDko
k60aOsjix5K/b6EPkEfzdxlDIJ/NfTDyaRyWQWPk1i+6H70sxsj1CpVoz6ACEpbo
ANuUEUfAK4dSBQ8o8saFwOnl7zmGQIszVeRI9yectZ/GEEsHHl/y6pKt2/0LTrny
DkhUDUzThCo+hPuGXjBt32+VaGY7/j3ykeHHPB7T/bUybWCeOZVRYLSJYkdOpS6W
5n7I0MK963+Kn9Cz0Bg2cpJl2SNQWBKJw6a4RMTWixycWqKv+qPrJPoGq5VTs2Tk
NYQfO2MuDqsud57cVsoLINR0xYhORyUjs95o4ulu8WogQ9eGqd21I6iPUxemSAgZ
81FTdeqXqIy7xmhlg24GYIZ+eHeZdkOmFu5Blj3jaxe34BpeUL3Sh1QJ6UZNNaxg
J7NJETksxqdULmkxtok+urafsHs+OabsihFo9gck54UhmQCjQZAxicDC5JfIvfiy
qWLqxXUrOfxAjSewkkPbZC1r6JszcfrXkWu11pSCUGREJcyC+aBIqENQVoqsGlVA
tYUx2KQQ0DpL0tILZjBTOnSohGR5QJ1eUFbna5mlCBhbH7VPM+mchUohq+74mL3i
+Q2d83gxWYOcj/exdk7QpAdFXuRU+zIuZuo/c/J56lajdxtaaKGzQulxpZQJQY9x
vwpQso2u7f6RcJBmNUEPQRMfwKttOQMElMb7JRsfnylr3MaJLOrS8Sp5kY47WPCd
cUcFfUEeAlggcgL5DApudfJWiQvwC9dqQsy/qJUl3lD6GbDTDgYL5flXbUHnGbhe
0K5oK2gDL3QNDmLtw+MI62JohtW5T0CcUaSC45O5dDKZ5Cric+092MmIisOchLZO
IXcAjbqg7l+CE4WGOSnCQP0WT7SqyG12V26wJpPjjVl+dbczv+Ci8epXf8HyCk/z
jy6lvgtiD/9gz70PBb1bRoNucHmwbXsSIOrAytguj0r7DA9OEi5Qyncgfdr6epaJ
oh53nS+6cyeYD6i1spYoPVELwCCiVNonetaF4YsLYuncEA9GcjeprdRgfYBn8EPy
AEbzZRuk+GdMk2pRAti6WWOVqAWPwR769v07p/14mHfO4nM0w8gOcxeQbYjs2mIf
MAuiTY9vmcNkM0xSZZXzbFQno5l+zodwp5BVbRwj6CJTr0Q/v9LQRl/ZpZF3ev1W
yKs+MJdlzyMAG6Q/ZjC3RDo984GjtFbbbXII8xsk+FB744VR8oP0rTKuDqGMB1J1
/NDXrsV4UTjR9DfbQ/o/tCpzdU/iDqsKR/7MbdECwnQlp67GzlvWtyvvvXo9fQKm
kXX86mT89puCj0FqSHUe65ied4A2jr1RJbueoF3SUOaBHAg7F6ygfXPjmOOtJgmE
FOX8+rwnaocvsfgwVMMUqhq5CfRlrjKd4WrMdcg6uHZ+1P0E02de6puPFMtMiaba
6Vc5PWCN79ezCYZgMfF+S+XC2vmbyIhOXahAQUfIh655vdBAQjZs4iy1juBh/BHC
9oFgUmpDx3FhiBItLwCtOXFA005u25BY7N6zoIcsA9GUR5TpbeXe5XjMPjRzqymY
8FVxVipzXyFfjvGicCx8SqL/1mkP/OqLvGnXcZGWqrto3R366/7f0HXr1qltBVmk
CIkN3iH0Vz9XCqvbBYZF1HtXL2i+Zetwia4YwGeUJxc9RIPYQkxb0le9C1yU2ayS
/BTlqtBFHoiirfG0qiufVH0dR9K4+6ZBQZ22V3LCMSyCelrC/nyFKQpsvTQbBjv3
M9D8RKGfFVV6B2C3uTDUeWXjYdr62iKRy1Q1q96Xsj0jE3X8dlsVY2vg4Z7DvvPK
ED+wBlupOywj4CZZSKFNPFkPhfAcY+OYmNGTiT94gKwnk82HTG2HieHhJ+Ipubji
2Y4rhDBNuKrWgjyl5oQlwrZariWbgoF+haesX7VRm7Po53OSd1F8QsLi5YT5LcF8
garzYsNX4p47vZywu+jUwC/TWbLcIaejxNehET1kI2PYWyDyexMRdfe98ujxqy8x
bnefZMBkrKnuROz4RBLXRt3Rf8U41+QdMOj6yKntlBNcMB3zQSk2an2nt7bY9znq
rMMhsRqTal4FxwnG13TzZkv6rccojnAB6aKnUPUk8fRt8WdQ46dHsHZfbV0u4vBD
VxxmyZDGknYni0Jj5gIWAYjy6+DQiXsB1mLq3pTXKimwh3FDY9pAhnKo8ydT6H1t
xAS6ny2fdJUtRhBz1oVZ7Fkpp09wVbjigK5KK/bQbcrR0BTb87aaaErpuEASwHe1
+mAmPUaZsp2iSe4gIGeBlNe3Kz4IDrGSNh8KOtY4CLOuANFWbgDj9S6i7mXX9qEJ
ge4zfVkMbPsduVWTKv/+4WV8Lq8q290/c6BNLfCPY9ohht0qH3y0f3iUGeEadlO/
dJW4xbMuxoKFoVgCP4Z27wdDBURPxLtYXTjbpPC89VEJaYVjlIS/A5URfYGslExW
d73sUhP7faJxmy+RHZpc8ST9Rj5f11qNN9OWIOU4Ynv9Zf+wysBprFZwX7ARIIvm
pojNu1doCPQIx9j3s5laFm+mu04hOx6zbRK/W1tnDn8pP59s/DQiV/wxLBwxr5hY
nr5Kq133f1IbcdMh25E9X0iBB8EFPMXLGBntJAareMpfVHC8q0pZ2f9YY6g3Qha7
ijSs+28BNgbXSE5nojjr+VF5ala2N4Zy2xMdT5aNcT+N8y7iSH6FaY9Zon7Mq429
GHhyhB7yYY+yIfyzSUH9raQDKpc9jk48g879Boh0XQF5aQTN7Ecgz8zoBNAVkaOp
68G/VSpdvJTS4hT/DwCnlqNmTx1ZC8mv71J5vYE3twAsUly6fAGy/wqzJPdPl70g
GnmLJpRJWpfhQCFjvc2BAIXC21cBTvNPZg937tM7BECiwwTVr2dH5ghyGiFwMns+
ZpezKG608plAH3YVwT8f0mjFbb9atcheTF+QyZgI1zD06bRbZhORY/KRomR1RlTD
dPIigRvG5ZkncowHUZpnOUO7AIfzYFupXyzwmGDwtjZgYyAKbFd+k1vx9qdMEFdX
zLYnChHAYPnOSiZqOLeBbn4bGXJdIgSaObG8H4xEWgKMqtdneI3yhGK9ffDCsWVa
m0A7Dsy4Meb9tpzcoKhbQyecBKYFGpaOhncVmw7DqDqrJkmpheZoGCG9HTdSIfsU
iFL3nl4oBfBqfbJ2A2ZFLHwUlt6lNt5H4M6SLtvkYZjxkUazD/WYqPaTwnddruPM
/mDPX7lH201kdkm1OrL/E3otoCEex7LJDo2iE8bP652OjstSpPzhruu06ZA/Gwdf
Ncc+/Voec2IDSZYs/X0fRXp0UtzIEZ0PO1nVZSRAhOQ8HX/KoszdhLdw3EA4DPQ5
RHab6ExpXRMAt+Pd5JEHI3ZUWPf9K7j/K1SeWRH6SfiwyqwYlWekDak8MTCpIgee
/6+1Ast7LklVnv/Fn9lCihvT6tAeHEQT75XQ1wxg21eUNNUL0mzbaZAqE/Ozk908
UE/0uHDnmtPfeliSttLhvTF9RJn/uwI8W5NzZQxP/wpXdijQmnsNIcP5MhmaqtA+
C3WuPokm7uM9Q3xMPMkeJ/EZ38uPSmLEiTa6qapwtrwIRoTyMfnNGuORM7aoW/Dy
aLenfgQnojF3DeMbGrMzhM07PkC4xZK9FJu0i7zH54E46wiRJhSyt52J1dJuyKTt
c23QyCnWVRCtnJrNYKFJZf9Ex/0pw03oxX40m/1WSNwZn+RbNxpUpp6qUyLcoNMB
WCCikzXybvUICWwGDL+Hx6l34gHa8KTp7w+OeRutg6UiT1JFn1k+5cY3LQd1kGRb
eouBYqG9qBN43qe8vcTduxQycHntDfIeQF9rKrnrMz+fQk85W6D3+ekiYyZeinGw
qkSXw6IJZB859Al0Silax1CWDgxOV+g/a2L8oum8HfP1BTbtnue1H32YoSIU+RIW
bpoBjULmen5aFpk6qT+ls+I6rTH4ZVUGIlalAaKiFJrwJrP1ikrn6r4LlJrlMJYy
M7bqOCoekdQAB9Nt57bkgHP6djGC9PqHl2qCKFHftiyTbf5QEIoIEj6ufb8Ef+oU
Ipw4Ipbb6oXNhK0LSAfdbfeewJUnD0bziimfpEsN1pX9yxKFwDkTTl1zANaLxefo
MeGWo0sNtMEXhOjQO5uBEM7zW1qg0GisyZxEUjXhyqS1Tzog8YeSVdajAC/nMfCc
4MBtGdL9yiqHZBA5ou34T+c95HF60WueaA71D2EVD7y+QHx7ed+KaSGVPvhNenPS
pnmJsqKrapbZVRL+7HDJCMvTVjeoL/A+gI8cSwdWXGeOil6HzjFLM4ESl3x3YZdj
HAt/9H0xMyGA/hRuRP1rE8p8uNORjCwDNj4M027CESxIDQJbfRIR9B1GUAT+4Oie
eHabEOCWMdCn4bFRKeQh2uhCIRIhGF5p/7xsJSznJVIIuvmMwkagvApVlQDDC99h
TPxXDp5zonxKTc6q9sXSGTupMMryJN7PqCqJvw73vKKXA9aqjhtxgbOBKuiHOSQy
nliw752tsVvA/Nmdw1OpAhtyJwcVihaKD5M1oVjHxlwHvyB9060So+XaAzPrC7a1
yF9+/gtmT3VO9/LvAMC4nl38p7wnmnbKzSK1VjCBGBE6IczdBJAXN79wOc95u6iQ
Mkg0cvI663RipQA1oLgN7qO0E7mWYN9izligkLUzorZnfgqxNPGTN6z1T4M5Kv2U
IuwonT7u/vFq0RfxS92CasKiHhZcfHR9+JBneDiK33BV7upjX0aD2a+/PLL8jhWN
/PN+jH1Vs82rdA/ypIKKuJkAfxaXz6YX3Onj0Nv0y8vF66Hdnu4sqodaG5EP9Ml4
WuwBS3b+747Kq9HjGzE8sOAboiqPqMUV8KRXx2KbNNYpRzwvfqB6lDPbw8PpNP55
wKD+2P1QoSe8NJXtvmYxAUh+Njp0GLay6M4YVutCWDsjEGUz07b/z7MeWg24WYGC
Y9yQYF3kbjxQGsNKKqaBBcWaYGU7BP9+7h836iGfTAuJaZdyfRwudWXX25XiKWhN
H7+pu5cs6cRhPEZFNUuDEcHBu6jh7I1gO6sBedgUWPaY4BLlXjRXXpDSKlYiFheI
83NjTFL/Rz9iL0rVjhgKxYUk5ylHF6egQvxrN4V+7QocqYznAfE9SqpW6ilxaOFH
o8na9lxuU7uE25ua4NC3wBb/B1zzS3ViwSc6O8NPoh5en5x8BgPqn24ARS2Tb+oM
Ynml2MDvInPn/IerIl2XSk/hPx/ksb17p3XIIlG2jNB9fgzLOQr7fME0ek2ayKnR
vgPiuQ1XV6gl32NLapud2LGSSHXRMezdxTPC0u0H/JPAwf7sQEEIcG+cinQyZms2
QfCQAEuwG59NxtG8w1Sbca00p20Duje2HLRN6+Qq4jWt3sCezcDQnJIgggR7FFsU
/viU3ymvO0UJjEGmnt4v81ZD2l8R4fcRbeLfrFXVL9QInhEVhIsVp5sQ2CQNRP4t
QCpCWS8e27H+2dW6zujsgoVl93kIJXTs4GPT8SOdpf1dcFWNArVUJlgirij2Hpe2
hHeyUkInVX+F1oUsZL8scWxmV4ZIuMbsF8n/WGNT4PgFyswQRY3bXb/yxjKyxJd+
0A+SyernDB+ezW+t58CMRsSsd6/MbDzi2RMlpJo3xPD8zJbc+RFLm1Z7Zr/cESD1
UJBVu2Tq6EU6qcyTjQCR9GMaeWWiAE7W0NtmUgd1klNAXFiJfw6ML3DyF0Twvzz7
C8rcyUrLKrNu0gnXWFMP58hO1VTM0QrPkBMwbUS3DFkScCNTVhIMW1cgK6zRdaCa
bnbcffXKPNlNGM8Kq3UqBw8cMob17NOotibHUxzuQq0UBuX9OuxAKrkgw8nUZeYo
P9r0gIeE6KfH+4lQLIawXyNYy68BgDC7Aeunbn8rhSNzcM/3jEUXOH68QlGemwJr
JbOPnWppOBP3IZ0BvPun2M+YJLUcfFUBP3vWtr5IH6CLQUdD62kWeFsN7JOjdrEb
y+E+l0/7BFbh5DpKTgA176cZwZTzTRDJkIAOkERuWzzdQnuqta4APtQ2//gj1Pe8
nPV3gy5HgDVrxshttKaLTVoT2gIwlKSykfVExGGYkh103nhRy4xJd4ctJb3FhCQr
2lV2/yoFl4BSSk8XgL7+8v/yPC0tJAkbsRS8iPrrPc54YL/dzzsgsN07fy6cNUn0
v65qRfON5eCmD/G/V3Sg8FJdXdi7kVeAob9lIPzJefGgq+tckGKAZNuTEO8T5vnG
kACqSgifLYdZSR5AC388XzXd5F/ygvaXBHJ7Y0QELveUTQCGavx2o6vNcIn14Akj
uvm6i0oJxI+zLH5xFKGSkXyX3OMpn1JQhoShk2DZgcktMXvzfBXnYyowVQu4x3R5
+5GPebYVxqpSEc1aBlH1TjNqyej4XtupPpHikjT+BN6/UVy7+mN263xmpdbNxySN
hMeq0H9G0KAMQDw5GlnsVjONIBbQd9tk07bEDbzun8AqAPZLOLFatk8o/JV8g9b3
/0d/FhYeW1o2JzPsYHzeQq3z6+bEh8rjcWkwoRfH6XwT1JIKna0vnRPbMVYGqe2n
Hcl42yyLXbTp20BwMw1jZ/qdKk6dCFSTWB3sqHi3YwNEw6b9DkIDbTeuN2f0PcFw
sEX7YTnbw9KcOhePb66L35fPl9WDh9Jh1vOaDb0uW3TltjthgmuvKwYdE+zboB4n
elbq3eOug/yDmE0F1BA+XY3tDBb3dnsZrUbHXQtv4x5iqcZlevPSnIi55JTxZAdV
Nz8a2YW5zUOr0o7HC6T2j86uH4iFmJMpGZ1F8mfvmHZIq004+OGBQT045IjMq8p8
cWjVWT5xWy5TPctJX8BcH9wDpi7dPU+OJXiijTtCuXuIZurXesESDXHbYisPKJkY
wtAtkEAkRxE6/+yHka41RLTOMjMvVY4zbMz/CIGktVOGI7fFa/VzKLddKLQ48YqU
rivdSZ2nOTtcsTchBGsX9zqVN4Jzm9nw6XYpY128cjOvED5poLy07oeoyDGzfKlU
ZG5hCpUYrWTo8uaO5ysQO4ACmxtyBqyf3CecXFeFpW8lYDILhroiSbqT8wlbCdQw
qh0EP2VxgNKaQXloEttDdLL4FNDss5AFBKZecze53dQNz/Eibk5J5x+xkxJeXZwL
+YSGt5TDQKZqXJ1BjdDhuDuJCMTM4GB/lhoKm7V32Vg4+HwHQTkkVjVA6B4TlHLf
Uxw93ps2ATcGXSEx8Be7aZEOJ54/+Ri8D5d+BmNByW45SdAEksJpk5JnpMdeE74U
iW/2D/SznXMokBMTLg/NDqyeofFx/SkNqLZi5aEcIjA4JHYl6Hg434rB1AT2j3aj
jSTvVnOdYRnhgYGUnFXS5AyaqTpKUtvWzmA+bhm+fB0tlVg0xqfwZkyX2AOGrR1+
RVRR73mqEbCl7jRPHeZwl66qeeLSRwZquEvuxGITFRiqXIYET/lH1IR1zOdIGgbQ
N+5vJ0ORfewdtEAq/AXN4o+BIWf0WmRCNbmlx2xwQFE//Oq8xLrR/L7NqYnSg0R/
OVcVwY2Db2g8EeBRzcAc6gKKYDIr9EHe5QthyRlh1koCc6ev/+bI+RgbyIb804b1
q1d0ww/NJiY0b4HyDBD32uBm19DDYwEwHVyCTxa+fULNNJDcaE2DNLE6yQvXLyr0
jn3F+BqEVMIeZyBGpVCsTc25EnMK3tBbZ58dhIb5Jq2xXTtvODQ0i7D6YVuFW8Pk
I9B/XmWB6UYIVLGNxd4tXIVrhdain1edYJa4NQtDRBTCNL/I0d3MCYFE6DWw/jB3
zyx6te/viBhIpq4q79a4ffDggPh3rEW228fWQnlMOymbxaAPzyzHkz9QEyzEk6BZ
0M7ofvyM+cC1g+EBM25uwz3m2Yz+53TTOC8v5NdZBIkJjb7MDL7DgjXh/4dOCMnU
8hcMEwTox3v8JnqJdEfEoFx9cPkjDyfyI7/xzb3m2ryfq8Ms0eIZhLhkUsSnp0pn
I7dZAFI5vfPlmKUlbcdYLLu+0S++0hktgkvVnIpTNXGZY3NsyDDNsG/zJVal3nLb
SwoplTXwGGgkj1akLJIMLaosHReurLAGhMpraNGrvgfVJkiRqvVMV8ECzLhV4yjs
WM1K3AAqUmFx5FhA15ggqwF0gNm6KPXfsdK8qxPqN/GDETqS3hYNg1fvy8yMV/SH
WcWSd6XcpO4Sa1m9Tr2u3D3VySOgKCO43zP6WPMkX42CKLeGkwTSqs3w6EM2RHUj
1yEsBQ5Pk/+u3ED1mKvgxcabkoz26PsROibzb7lI6ObEGoLyYaxS0TSMmlNcsx62
4udLoQ6ArGY8HcSUUNPQ6LGlL0hH790QqWIMwy5NPRLxbe5c/owdJg9KYfjZ+DG8
+RL1AHnc6ATPd8uhuOBBHSYD/rssQuWb11E4w1NHE4o1akfUbIE9mw+1y4dW6i6n
CPtslU8jY1v1c8gP8vJ6dRLZp2mOaMI/eUZCZi3yPzMHeU8urSzf3Sa3tGqks3/f
qleiM6YwFPHJdZsPWTV7CO3gdp/ez2kdq95j2/c5Bll60ek+p9rVrPItGHScAiYc
gb12Ku+mCbUUxWw/juaSJFVIiTZV33Zl/gVIqK8Zo7ubXmupCafkiw8zPbXEuKrq
kQaZAAqdsn35lnGsiiZgPfzQ2CIYNJlclZeipziLw0EajYD7WxUXOyFG2uhljU5p
vKN2Oer+FXEK0DvsvqdrT0pbld/cyR0Ic4ckdrXKA8WHL+AINNm4RcQNpH9nZyfy
joNU6a5WzkyTs1FScCoL1HBItmrVxXB2EQ0GRIld5OxTtdKov84OWJCWE1c3M1iR
TxRWgD52Y4mCboxI2Els7EXPov5ZimZS7cZsqI0fVV63fhWSnm0tKvzK4sVGLtyR
TLov4DO+N4ioaquHqQzZHrnVmu+uLydsz0B/CzrPT8vN+CdeK26de+9tHGCdDzwa
u/3thq7N1dAX3fOXJC/dA5XPm4uCrCtP2TaNeXNzphv1PGez6UE5Tcjc8BYnozb3
f97SXjdkLIvd+F3E0dZoZBg2J8rOEIvsulO+4d4lN+3Rc5EDtIqeHSfALtA0qWMN
JDwoAY9ECO2qNskqhzhSNusKOqQ0MhtE9yBYf2N1H3taKpEPIHxbMtKPVa2xiHFP
paKpStcFfahe4248/yU/iurZju7e9itn6jG3d2DmsOcHSa4Nog//Z5njYRlavRI4
H4K1Pz0pvIZ++hsYx82kjoFk4dVQQEnVZQ7XY2jeO4L9icll95T6BYv5Q3hpVUuN
bTcFMkemlZnOplXOmkqhCr2gaY8d1roKDOeTgnbeg5mEjg6Fa8wwq6DfNctumWES
edZdfKpxTc/WRzk+8EpXucmlYwTBZ7mV6mQEbUF2tIUkQeimAco71u+XJt6wt5Hj
yKYUoIJfSn3XQ8+lT25QPQwMkksGJdz2smCBQQlPLoPdW/qP3wz8ZkbKlVPDmPLH
EPN/sFCb8pysy5MrJWl0o6vAEPvEMqPTqjIIdKOkohaaDn9gcCxb0HE+H3/kz2bR
FFNFpnOXXNtV9LlE4ZEKFsOBCgiT+qjovVYSFgGxbIgyyLqnqGh/84zb76pZNhUD
CpR+DFqP2TXScAcQezkFiOuuwOJK45vzbCdq7BjhVWWfjbujWVy/qxRUCsKPjFkL
5GwY6612FbLdUP9PDnIKnxzUFsqPfhM39imOi4gRFXiv8NoxazthXSCtXJR4jo+R
1OeHw+KgOTElMdbYNcaKUn8GNH+hO7+bOYgcbiBh1POWPyAXW6oHzCuYkbW2I8j9
wMoYmL2b1rvQvffxGKa0m+aLx2mrKh7Z/VXt4wYyTy1n+OaufsHYTY6rquza+hwu
JXrZ+XbL4IrQMexGW8fYKEe8VoRXcoLYE5AT7gYemROUHIORtmmQC0XCamrD0WNF
QLjLwXTNKz3FjXpxftrzv9vzd1zvNWChfnwApaJMtc6AT9xprLS3rfNzNf/khsTq
iCX9I7OYlQnVEqz04S3cZTQigCGbK+krWklYH1oyMtEZcfbFcrcQ53U2pVA4fXPC
qp3ekqcl+xD3B1xxN29rrpAmytOe+MhuDjltEjX6f/dV+iPyGy0KN8Qy99iJB5I5
nHWMRpJP2apqz9fiKCPNj4sBdabXN61xmvZdFyPDBzfaBr5ppt+0O/BPphIz+geJ
qrO5RFgfNKDAbRkjYYUGJhj55trS/xWWs6H8nqxxPO3SyoGR4Fu5qEGpa4uMBjvN
bwHECN3md1FDftwc3xs8gy6IFB6WH301C2d83itToFiyVgHjOgnKNOd0fgtrHBTz
fmmajl6xFhlxHsvmGbVWHdLgaOnELds7Ax9S5DZYBSJGQ7uwdWgVszLW51T/gEAo
gKuNE/4y6TYdzsa70rwFeMERnnROUs5RK+ViackYVLbPpQAYdJMyyWBoX0a4Fe/G
xN7bgDdZehgXpt6G7aorvefIqlmEw4HNcdkh8NfR3k6FEHBWdFq3K9nrxfA7KPAk
pIMK0awnEi41ydbdni2vBQySNS3ryGQsfTsMkaGV5Z6bP1tuDETHLLFgwZ59MoYm
T2EGfwbs1fqdfEGG0Fz2cLb+YkeXxM1NdNwlE5to8hvGhU88LP5OrfOF5VVEKpQW
Y3H3RNwDYgvqGyxJI1Gtr7PpAaIprpwHZRl0YD22o1m+NA/YPGdCzk3VAOQJYNCm
RMkXGQGIw3B7Y32sm04B8kEGb90I6ZATLejMVB7HN3kSjfQLG8esEKpAT0lnyHUv
qShcyxJeoBUHPvWcFo9wByh+340+boHOLgwnv4uF7nabysiGBbuq5oOLbwlxGLhe
RfwG8CHOXRgJrOquWJ1DoKURoEEm7db0XrHrObji98ZCQFDF2tkUeO8daVgmECJ/
r8laKVQdwmagS9N6KY1pqyx8OxVGKAO0RMk5PhQVdIVXOVwc2iuZEwjHKn2Sylsn
b3goXbfyKw2RDdym/0NX4W1+kvg/cRp4I5izybImzs5oy2rR00Ea9Jjy4DuS0Ol0
pOfDXwD4HR4T6Kk38k05daEXljnY1FQNsOr7iYOE1xWhzHEC/HTgL3JURTnQghFR
6Ruz1j4ehw8LGBwYlySn2DOUytU7WI8utVNuVmzhnhmpBcudThsVkSBXez5GVk9D
Bdx1I9GcEiG9eZOEeyPR0Rh3hA2ARzq/p+P7FfiScwWVidnnJevt03fCibFKsHhS
pCjw64GZCpukyrB/i1+PYrRLlt4OUUNIk6UZyDxqXoq+cY/YfStwo6434sIit1Ui
bkzJ85pTN8apoEj/D6mV04+zNbUrAQ6LtVCY+is8qfQPgQS5eBYjnLTw1Gvy3oom
QGAkQfGQdZUKpdGCE2qyDNdAdnWZJrKgZgrEkor2Z6SBKyIycoVf+ZZBfkLOwknp
hgHBcyw1rMYLU+Hojy7IWlazeqxd1aoXm2PK20oLg68l6EalpLcOHAtOPe8WCW11
v8IJp4g2Jlz/XRIHxKKmIohE8Jou/2bj1u7uTXx4HYJOrlnH1+Anc0PKjgFDHywK
mQyGlIbMconGcHJVdVDNv4bRsP6DMYGr9SbWX8uYtDFowR6TrClR4mgOwpUozLp1
WT2/FI6ot5Dq7lci+YABW0oX5eS1QbijN7XYrhEqT2MiutfD9cyZYpPQE0sraUVf
KB2bQww26xTUSXzt/9/CHv8E+KdV9pbzFaFghCFMeGQgUVL9Eb2Jhw6RcOhYg+fM
PRYqjoJyim4M1q571cHfWeKBF9KdSY1VxkXTveVTkGAnhQpAKfMy8mpfN2qIHdRs
GsZj/t+em8eRTzcpo7srSyxdqMKj1wkcFZB/JY2am+0bPWJUoCLpjWSCPHyBsw31
Zf7fN7a+KE7WsuLjop9GN3vHSAJAn6qHLPn6StIQ02D7B6M5Kau6rNMQhTf64W+G
8fit/cYQLFWp1Ej+vSZghqfKpsdAv/r5vk6HRJxYbPId9PpvJAa0t+r5/TVsxE1p
1xHlKFanP/Q5bW9qWMSsXQu3dL/Fiw52OcGCToG1S/73o4Pq35xWuN5h8h31JIsG
B0efkgYDLqjwM6feXtVgAV30RChIcaQQsfYAG6asvBqBec8IWn6IVB1S0zpRyg5x
OI+oJajG2+Rsn/o99G6jEJ3pz1jmiXglfnoZ0dTDp7xBMHQWbevwet5ijgH8GGfG
Pt/dSviv/J9TiHgwdSXXXr0GaOQhv3B3QFExmwugSJbmcU+nEAk2fl8ZYBm1Rp/K
1qK39uRylS3RG1ifrx2DO9HeovBXExWzLxhjMUHPp4xbZpSLGwhCvGPsfmqAJ03A
qDvkSBZ+OZdPCAHm2qAyRzcVZl5+dF6KT07KaM48UxBWczlA3Vy2rgwKr3WHCx86
RVM/n4rSqrn0DN7gQchEA/nVHPHqbkSJ2HaDE525CHjFfVD5o8aIEyphThFbTxFN
NdoqyJKeQruTbJRJQwAxdMIxlZXYpOAGcjSAuGgeQD7fFBhpSXOxa//RyFjiFm5c
TskMFV+P8OulL598Ycv9ZyM6NI0FhZr9qS6LMpC2M77gyu5FkiDXEw1mpDvXqz0Z
0QVI2s/iX0btxCzcp/KtOA0t28UB6/mIP6izwhJ4WrdPLShZeg0Ga68MvwnXCG3H
Q3bxY2anIJ4OM90zbP4v1DIFuNEySICvETvwEb63wILvaRwEYRztckV8Qrnye5b/
QTj0I5QBsi/ljg9Bupv3r2+VJRV1v+UZBVzdTX1cdS21YajwjQyBG6eWBLziCaHX
2/kDXxZJFOz5zWWWavv7Yq3JJ7bVVHCBJ+f+Pi0WsMTwpxZ+sv7fg/8z37mOdS6k
MeTePvY95xKQgSmlWf2G8AuPRU7LgHw4qJ+NCirH+kVp92lS6qRqarifGzXmV654
LY82uAL1KPcVL6jQs3cM8zIUpNC5ZBczD7xygHXVLFK1i+oAWvHqYUdihyu9Je6u
0O3YqdOIKBN5Oq05MAJCznjfrLNf4vraqqQgJA1Nr4B9eRIIJh27uYqQu/uZ2jF8
GWvuP4Ok37Ymz6PaGXjPDWTvxCItSf6KDdlmZXiay1XjiIMOf4eV773PZPSDenVj
sEJoV42kM+iQ3F+h5TC2i/HgSYw6B1amks8Lsi0ofos9IwIwW3e9FNJuvD3AZzGl
SWYUmX4+EEyjjRhZa06i/Q0jkQpM+HPOIF/eB/D34GfioxH903H0UxD6KUiAj8aj
a6BrQwng6P38hKfBLgOap05UJ5hkYkWVo4Sd37gC9bx+gdn3YpVth9jkFfTQe/gt
jSMy/X91BEmLaeyD/HNk2/CV7lpsQF+yZbjzvWkZXLgN8LLIHiQvnWdZhqZe7MzK
ONAfkt5kPD3fnVtsv5/iYXpaJtdhr1iURhpGLBm6Nt3OD3EmSCtw6QD1qdZKlRe6
HTshBBrFsmEpq17hNcCSjDDnzZ30D2BuRUN79rEAo0noOJjDElgf73PBDqeYQjhF
rveLoDtfxuP4zqU89s6/PI6r3UTrNtpErIDwz/BmKBDEUNqhQO0Wktpau8qZX3+E
LGzu5a+d47gDh0DMS88YUz+HYf1YPe5QoFGki8y7hZ4G0+asaAU/r5yn6axQnNoN
+Xg0lT/aRnhFcKuMqe/CzpkHhkNdpXjxkrgxDImRKlUmawQoqV0TsVFZapz9S5bk
Mk2R2GTesSqGvXGRc+6vKOwuRZTraNjuGsKh0wNajRolHWCtbRx7V7TUKohsexEc
aUGUSHHE6s2kV3yEM7BARPtvnt/8HkUSV5K3yQ+U/+9etQXYG43b2nT9lpoVj+HL
7Bsd9nXEhtaaI/dQzbBT4qr3zshrNFofnes2lhLdy+LU02V2IYsce0/+JCqItSBK
JaHJSSIsdMIeYtsyfpZ9fwRPwiZoTVQT/UKCwO/ut4tsrRcFQEFBPdluEnBeDGn9
HhyJKutyLL70p0wXvmKnaZXUgMhNLSrKrme18pYwuZ1QwAb1+soVMPb0yQ5It3fZ
iS12bOtMWx/TEix4nUN2o0rOFLQonqoVOmfX/C9ScGfkcYgWuBO4JBSGKiuOW8vM
x4keNMHDnp1EgA/6NFuHGRxxMpI9r//b8u+WJyntDNhzZOodcVCZGNnNh9Z6pz/p
Sgr1mx1uJsIwDL2qdFYvrWQ3sAQ2r97+9jfxF7M1TiC7QA890V6LcdOH4vo+I4Eq
hRW4BFHGAA/uQP4TOZZ9cGmfgF+tO1JdL3ae8AOZjDY/qx0PuMCs+Jvi2H7Wptgj
eAxwEqvdXqlK5YC/8Q76rQKUJ0ZROw17zSY7kyszerj8Yy1kQ0Ej+3o07kAt1jWj
/8VdaSglnReY/+BgXJMboaGL7QKW0hg1ShRTR3h6ywhzaEmgY3y6lhJgY+P482O8
OngF1kr9c7Gy2UXvtlAm96JNuM6kx0N79fTNbu133ZlbU3Ga73vf4MnFWxuNQ3eR
SiRVK5cHlEFy6Alc8hEUI5x3VXM5jjvI5/HXGSFUkH7HYVPiVy4x79Ed7rikUYW5
V5A3pYzSTkZD03v1k+C70O8fm/O4GLsgqDXFMAeYAj4u2vzNZ3Rh2EbKWxKle4t/
XShpe78caR44xvVLrjoqB0OZxI/wnGrdXnSxU0GzmxCfFBgmCt4YnXHPKCsjj00J
W4SbVl5DebTi9dYWdN8SnWaMle4cpekFDtXrlSFF0RloEsh93MyCNCBzwvCNW4/p
MEhkT3AkSj8Vj7IYtsA3rNvSAxjNhTzyGiFqb533m7TBp0cAWYym0qfApSrrfVup
vHJmV3fgyEzYGJKwrpHqGrvz/1bAtUIFNNkc09KremwFOQn2x7JEW8ZbwURm4yZA
LFEL7lIST9Y8C2BmoAiVOxAuvWOJQ1skA8I0dFkKMgq4BlW9uZMprpC1EwHNWOj5
YsUXSRIRZcpXUg4yoRVVsBZj4H1tTPfR7BgPVG9h+7/McLDYsxK2MoOT0GEctL9T
6SaQmmEDjK/QBSpm8vgcoNStnm396STvJuipdf8gN/hWIps0OE61Ow1xXWV6RTCk
3bchnKv+bw+CZhfsKiNAtlyTeSrO3xLj+5pMMTzlGTTSVrFWIIupdgYchdtudYph
A2BY6X2oMZdQPCHAtrWV1QPDzsoZffHz4adjDGRSYU7xw5QRtBSjpDMQ9uvei4MA
N5LAhhtXEW7HdwE6rlOdZ2mYSYSpaOHXKz94xAHWOIbEapKCMGOnuSCiQL0ddbXc
7e5+LiZcW/HAUn7EPQInq2WXurIE+wbydYoX9QreSo2lw1nqMgYZhB1/LPi6LfwK
FhWXDIrL4ZEmFusI+lK3ETlSFPnRiy3jRxC185WTkZRdbAQL400wtQGD/fyrXdMz
lWXIwIHKxCanRZq5mLwD3LRSqH8E6dXdanGIM+ETbbYrZP3Xm/XcKrKP4ihSbyPt
ObqUXho1OKQViZ3u3fSWlgLRN3x2SC1teN7MbyC8ybpQqgrZSVoiMMDr34rdlQY1
zKu/FzXKQJIn3BGGMAGhtWPJVEN0vC8HdQiV2ccfbIO1/3Rni/Ri4Wb+J3Gyp4j5
P0LcJDcJCmB8hYZ3lAnm8PVtaD88o0SgGwhoAjoJRbFIiozk5+pZ6ESSzTK8jsnF
HlUz2Wy3FE+yCuLr6cLka91DaBOnvU1ndJcQvwV839PZx4VQjMMpNbVpt9SpJewb
adKf5qUClMqKi5xHKcni+aU8HgkOAdoNWPKhYdCigGJ5zSyPnHf45m24q1dSjwLj
RMclzImB8BK0lW/eXaK8vnimDgheJ8qQSp4W/BYkLwfpLM9Pmg13R8HjSl6Nms3B
rUuQaeFAaUUIiOc15RxFpVxlUSR0MHpHzaJkxGTqymMFMQfuhHDcOYoXehebQpbj
aMeA5zaLZuIVSPal6f7BrqjnAYX9DTL8ndrgM9krZHwQ7njtPx/hh6G5fH8yXthP
6w1O4t3ehQQqYgmlN+Hbr4o2RPY0TE+1UdMqQ8LV3T0MGvb72STtOE81CDwjrgKR
zvuaMbsTbRQ4odFxbGscPDMcajOlYtrTbrR+rVWSp9pVE3R+3mnMELkdryBgmwlL
k9mNgrCaMxmVLVa+S/XcnbdcE6+4O6ftf/QwRy9FA54En3pFUv/vrEutq8nuF6kD
VWrcB7iCKubDrHSHV78UZ/vPHvZCFvS9i7fWgDJqIH5kj5WYSuNuUHlW0ddt98CA
r184faYKHEZvgoJBdvMQ2Ri7P+0gif8XYhNJTmIz+aH6lL/I7KWVoGmzvqw8ygTg
z0v7iMJl9Yc7TaUwTTbEZjor+Z66R6ILthYqFdmRps5m92KnnMm0r9P8ZhbdCxSI
ZIEdrIRivfqG13KdRqn6jOrn78ElpPCsNLkiJAB9EsUonYjO+RL70sT2DwdZgCES
OqepgYGDrCwgQ924YnpJMZRSoOsQN2vrLkkjWbSB6Tn8MhCakpSUkbAZ1ESm2LU7
ll1Xe5bJ+XipOltkSMpa9jOrI+fdy5++ldI8/P3HztJeLGoRAoeziaZ/UFpCz+hV
Nrl2SQX92qxBDyVSX7JDwe6JGmUTLErkOmDutlRNfTwl/UDs/bfwj0A7vpv283OS
U9dUWYI1A0zpdTirvRVWq6pLKAYS8I/GDGK7HOj4U9/Vb2P/3Z0Oau0/69R3XRoR
cX/9WvYr4cTmTLI89CZd7TK9xOdavWSU5DVEJmArmwgmQTb3L/41CpfKkdusTQ3d
jKKVauuDOULMwwsgSXU/cm35ZT1KiWFHZKOpCYR8jQTthRBKuVaUvB7b3a2x5vZh
MNwi5qfRe98Cuix9ako7ZO+ZJTNmA1r2j8oLKzBUpuuR2Mx85M2o6h4kqSo9vRxZ
8b5yyE8Cid8n9hlsFfm4tjinF2ldeubbvgTNd/DdPmM2s8PuLfiQOaBwxh3ksMyE
qkVoFRiaGnyH37Cx5dc+HQnvC3SvkhBsr+VCROTkIoMddsh8ozxwFfYYZlab9pU9
n6L2BAkJdKmpKaeY/yIJLnJwGf7Glqv+V42nJPySxXlTHrdV7/fChiXY+xgWpvzb
beyLJsLJdWrq5uap8hvsaP9uPelpGn2bc4vuHq5bErLhy68RBeXLYYmtTii33/Mf
ncB+SeYBzu0RJuqqnKhoXCRnLeeH+Ax6WmbUYyJlD1//hqLZ4kMzMis0D7UY/8T2
cpHVQaGRLmydxxzF/l0l9XQbzda/4OwVNtPfZqV75pVm/n9BQR//ZM15UCEUvnhU
ppWHeicgIZahnJ1k2Hp1/t05HkvbhqpiKgvcPpEDDqosNda+RHqRpdTKNybz6V7t
2mFMxAOr5sJ/5CUKDTM8lYPJyH85O5yy9Xf8ggIZxXfzoRzJEg6O55Hkl2dNFpRF
syt3uPjQ54ywd8CCv5hlglydQfqdETiuyh1L02LFwFHNz829VqOR4THI/5g9IsWK
GrIXqH5wjCiQzW2EiXPaZOPj1R/3P8LZWeDsIVBMiTYkjekhiBO4lZ8HyFuAJWYe
qDJz3T8ViAB7qDQigjrYNTrK1ZWA/fTddoMRJjtLv1zXr6Z5UrnL8R/l1GL2m/0S
8vu7jDQudKqID7fI8MB4GIGCDMWkN2xM93+1sGX7UxJulw/sikEL6v+lldrwO7VA
6IN4bLdIPxFXqaUKfdsz0Xim3HwkbF7isQf4f6kpVlrAgyRsStFz3drVYyXXvEgX
6VcxNJgHywNThadhD/ARw1lZnodeC4iiNuLpav8r5IY0l32Nkj7LMAZcVIQZuMxB
inWNpCp7EAqR0pShNu39JPFQGCBzZPTO1dE2pL+ke41m8HaGMP2hOAFG2hN80wop
bCJj/7xtamw+B/9GgHWFcXOiMOJgHTj51fteXfEnR/tHryvyERtMvMhO57syD5qi
kekm4NDtHiJCiliURmyX6H8VvsiQJBBL9BaQBMFFXz1YfFcKXhkhfEoaRgeUXnLP
fan5vOjQGQGzkVumBqd9In6V3UwsvuNHHU24783A6Bd4QjqEBAls2chLIyvY9Nrk
FflXqRsY9PQ9sisDr80I7bnTo6oxfOwemsQ1GeaTrsTPDtFI0N91khlVUs2gCfm0
pwDR5U4u552wy6ZD9oSoWNv2GbpOXzh68PR3Xqn6H/sq3PZO3sql4ZWR5OGVzzFh
QY6KDhsmUiv3A3D7aYtehdEJYku0U6SQrFbv6NRQMpa1a5UpHpXDOaGdRT/YyjJq
NpXg4UuU4yLcbAG837tudSjFQx1OACW/s2Ns2VpxNtBFvLGVtbX34kxd/S/GFJuw
wWtjrOKq6E9qRMzo0qE7WrzNE7173UuI6eRtffJNJi2TDGV/Xhhz/+X30hvQ3tf7
TwuDdoRVhEMX2z6CF04iBmGjsC+9ar6/x+bkANnd47eZ7V4Iab8ht6Gafn0cl1pX
lzgyVQbMTFGGtCtwEGUIYYHE6b9yyDaHOpKLmOjKdVWLU6v8RkrxbKznBijmRk7w
E+cpMGVliPd6nxdu6+/KUUTvCsyvSSO6iE/7JW86d4WUxMI+G8vCgT692qgheSZ1
4q1LVP5WQoHBZCavQfg+cP+79RAUBl7XgtHRFLxOzjQ3r4ApVWbn31wErHiJRg4y
5tjl7jb7iAFHeLMP4LLLvXb4beZgfFF/CFXHTKrJ73Li6WxA7XrC2q/4j3U/PUCO
jd/nfvTrQpch7qDQbX/O0EHaz0rAgGnL30DyXs8deP+gqIxooP+/166q3Pq7WsZA
VvoopGvXMmO2wpcZzgV6m6i8KOFWHRY9G8l559h+Xnez+3dxn77iOI15DtfgJDMl
KVdJOYyHMuXxBuiT72D4BgQ7aseY6iAwTFI+lbnLwUlr37EjDfEGwaYFr3MPmrYv
RUs3p5m+4AGSpLMlMhPY/dyk91jfvy+Evb21UQBmN25nGjEiOw/f8ZB79G3zDwTt
5TiSmGVNQZ2TuP/Jmpt3sNi8few9kWF/NcDy3J3K7F+YyKSSleapLY12Br+ouD0T
rJw/dhz76hObUD9Tv0TT3rjKM01auKDGBiZDxioPlCnJxvWY2SWIsBey1FezBojZ
Tm2Ko6/0RXzeIRsOkYkPGr3mgtMrzcs95ssjiZVf8MFW3gEzyp4ocJa8Ndxreh7A
QA56wmz8GBA37YBdJOzXxG9BW6aCVPkTIUlISbdRQiTufdpRPKMOmaNK27Y4CxnQ
O0+MfZP9QRnVrMKYeD4mnC2sV+MEKtDNRmaj/wCNFAt2Dv1I0CPMm0AS/4nw6u43
NLWGHm2mhnWPeIOlBhS6LOddczg534+jNPiHN8lVCSqdcViFeDxKactEx49gVTZ5
zN1VvE6dpJ4f4I6pQqHeNMVv35XYsfknaNXuS8PM2C7IiQLp0MHbta0C+7+/H4Lb
rk2JA1vplUCN4RqHyDOI00fMUyVpVn/uKj0QJgnVf+Gk3f3FKtMXeCED8tDltRn+
C0HCCPx8Bd1fMfmRvM7nvvcck955ljnWHD1vvf3FeAlYUQNg/Bz1RBbpYvQgEZU9
6zIzUdKsabDSpKEyzLk+dY5ubROlF98OhMjjgqs/zFrl/GxCh4meS8jznLSEa5zd
DMM1UKrGP1QK8zkMYL6l0qISQgHoEhWtLcfnCHy0xFvRA9Dtzvkyht1bgHIV81VQ
KGSxgQCPCBzC1Eb+adNmPNUyeAtbDV/EXT+SZPtwcgD2wI9kx0idSg3GRgcdtNvq
Q+5zTDel01pVlY4WoJBQWIWSUQUOuhu5VLrf145o3QDixgSKSZPA1PP8nRtGvKlS
aMMCRZL/NajIbUkj12jMAPzGjehoq+/26rQtI1DkxDrOmBdoOTcpB7hBB4zGjcRp
fIP3FQ3xVjuQts/Vu8PpY0Tkq9OtILObUHZbtv65bqIkj2XhnHgqCb6KN0/peD7e
j5GPjwLN5Yxv/+DRzssk3Q63mH/d16T498fFgNnXcysP11bgm1BLu1giErtoJH5o
U+aObbVhVrUJYPcjlDY3xeHnEhhnM9NGr6qYOmhAjSNFkm8cn9kYxpda1pBaotoy
WrtA4+vJInKXFgw2EcHz5QP/T5n+KCDpmKhtZU5jKB3nmtUgFS2WVR9YCKbwnAGj
I6Z6K/AIU3cSa1MN/SMD+J1kTZyo+fa6WonDTUsa3sgnjYrwb5AJQObcFXYC2X72
Vf8p5amguwbho1dWfjbbc52YfDB30h69Y/UBYs5dwxNeJNGDqZ9bsGpopmNwBMLP
RRVAj82Kafl0zDmBgNF3WSTLy+xA6yq0BQ/eCYA3siHZGXxdG5aX8iW6dQGpXEqq
zxAh/wtEtwXp/ZANhtapYOX/fP+ZG6nmc0osM+Lr76l2NFCx9PHSJcvjm4Y8RISV
RrTxAm5jwyS9aAtYJah7lblsS82HohCnn0cmdsHgTsJaeiGmaTMH67gVwqc2cgWF
WdqQKGlxu3OeKJr6vcMZllXz02HVkaQ9GzsdQtILpwxW3+SaFXFxZ4DKHPMOnvKT
QzLQ+FTuYfQbv1jjkdHNKc4OYkwh3fRHXN2w1obXX572tIJELwj9XsMmPC1HktGc
odpL2ljSE71aYkWYesVXtYcRk0KQFPBaPp8gkZABN+2dsgZZBQy7sOaN5yfiEmoX
UKe2blD3gTu1TlzRYj8J9q3pqEEJss9vagU78VheSDF+dnQLak3wzUald+ZZU2rO
ZAfNZvGRIEA0Uk9T5zT1pBFmtLotgOx4h10ERPvsh4Y/RXiB7yXl9Pu7x7CNV35d
0g05PHRM8y5fhoCfW0ilD7duoOYZJxj+F8PZoyENGXWkt1WU9Mc7u5O66QKJoG4r
hbGWVLJzTMxNRd3y8IpxOtLq0tR8zv7p0hja7Ng/hOFS03NVDVeN5tPGWvZEAs00
UNBezRDbglqizHKYpCrQJNDxFc8s/l8Du6s5/OSi2MFjY26zOvVQ4or4y2jdMekH
bvCfie9hPeQxEzPtTDX1N8yPEPWWB3aaxwQ9rCeEgoj5myzMV53o3IahLT0xFpYO
UPjLoBn6UfjHWgIblBEkVhNtUf9m0T+pz8N6KCoWPW5LOkJHaF/c62Us4KGPYF6t
kWsVb1mGi0poj1ONQLaF4vy1QcU47JYVvYOOKcWdOS8Ummynmy7ELRGDjh0VhoBa
kzDx/6y0XvkPzmu5Y3VBER00In0hWEcJ4A60pM5GeYPLqAp5eNTIZBnrGebtDeUh
Lz0tvhrkwz/zscgldRGnbsw1MNnci0BpxqdcRaIsAAjZqzRfPpISItC6+6fNyfxf
WKTuiE513XgKOnX0aEghELmV51Iw7IXuJcPxETvd5sr7+0O6EGW13MeIVHuOb9/o
ofd787vS0hQUNIDEEI3Xu+tROXYGdZ1Vq138B7lgpLczZ9o6kHdJSybdcnaUlsfo
xHUVSSECTGjI689ZyJryz8vBcla4euEbeSjUPrSbV85J2m/f2iZMm9U5uNXiuH8i
QesZvQekMM2kJ65QpC1NYNbyVnr5QC5KoGR/PiAm9a77v7yLUUwHYQR9zFzy8pdZ
349c2PpUIayLmogo9JZGeP3Ox5g3lbdvrkqJZsw3RYoFUrJgFXwxh1BMHm3PSWcS
hFGnbOAUjdF540VQSIsjMSbAcV8H9HiOoPTvU1IB/P0MdLAMiTSa8WQIxK9bPZJP
UQOTZyqTR6O12smot9GToslapwrB/GG4EjvRokJkc1QToW6PxnJ2LQhixqIDwDsB
dzS7p/b3ROAaOQAF41kxXghfjBCFshLwoKFPKuhjZVAZ+jPMVss9mQc/oh/eQ+Ht
9VXpDyPmkexzE11r5OfSXvgIKCmhhz0dgA+iPheiRP9oY74OjCzri/ioAAprApwG
FfxegFvNfk+Xx6fNTGorxeAzMh5W656IA6bgBJ4w8jk8JfxtsaO2pewRKN6V1/MJ
LkREmVk+cNv05ESKVw+xLd/invsmuApBNiWut7YYBZeUVBrwlb5sAOoIaCpYA4HU
vH393tNqUNNhI2tsXuk6pJek+hXbK7WOd3GdEiZ6x2oeqxdiMMTpvypgbCHcIYNs
aZsOoGFdTrsULW6WS7YpXMRebO9lt8jFDDGKTgtfPGvkL3l7c8ylKkKc/wW2w1Ae
NfZfQA/YRAZFPm6T1qnHBgawZHKoBvyfYUtq9TwfjhZfZkOz0/OJgWpVxMYB+aH2
2A/JHrutrIFT+uFT2wQJvGrRDOTu58YuIdAWlEsN+Mai0i2xiY0soaL2MAjUaBEX
8NWkdsglD1IuUDrw9TUIItfQCUupSbXK63KmMAUSBHlquD4mHjaw6TtQF81VI0yd
jU+QlNqxsbiTs6GKKBo0sJcwfb3ORqzANIg45sN0APU102VFt2UIubBRIC6RRHBk
PXCdk3hBLrBYI+gA6uvTA3qXx/rPRQNYTV93kpSyyIjboINJjewftrsExsRiaa4w
nIl0IzrOGcryZXlOnY6S9s0K6bSJHM+4niLxRxWycP1hTXdXL6RmX1afD4TvEP5q
8iglDcNzSueEApmuHbi9hiGmkG+eWovsRCQhusQSc7WImrHDs7xQegc+9AQeTX4u
G7hkHh4iO/nFt5fLAXGtBsOFr9NsFLY8eyanTwn2OxqDyt3jALQqVwcpW5AQw26a
A49yvEG2nzXyQ51agZF2pSThORvKOVz1VO78mkLWz0Ka2eDbYKRmffRq2l40/gWI
xvsW+XYONa0oES983xqhmDpwuJI5gwhmdKlACMjvZSvoNNUatlmX4U9q45laLSvD
4dfkZtCCeD5IAh9R8FXWneJWdlb8uFNjNU69nyqqgeWh42g5Ip+6I757I2zlcdoY
umtTBBtEPDGf1jeDB8lGxNeqIYcQvJx6dgQXrMmSumY4GOWiNCHwnCMqsGDYi3/x
ElVQJ7bqUds9B1ibVoA67wiMRabdtKFFRg1X1ZNn1Z3S90vHxST3TVG1rPx49oGJ
zGSnyKXi6LQgp8+jPxD/GzNzYORy7w2fVDGCx7PNFlAeJAP8ZmCXK0nM3JI32lFX
mlcAlp+H5OKEs1ToRN9gsVFhm3fvtTP2D52jOhUlMMh0ijFMKczP5V+Z1xovm80A
qzicxVaiNaMfpQCa0+EuK7e4B8QWEOm4eQ8+FRa/ftgru+if+bytvr9Nk7hHu8Gn
DzIGtr/RqeKCOmS7LJiRamXYoQJr9e+KIphmZ+1Zj4A6Jr/oiwyNPcNgSaZVKPeg
15F8A/4zrjj6AbhR6iK6M1PufvRkaJGSjwiUSB3OS3nN5fJ1srXBUG4qlRdY2CWw
ABTNQ5l8s/wd0zMoBb41YY8WYwZ+U4hj3Hj8cpAz74NkQo0QqSZP8LoKy/6rUObh
S2g/YylIYPnqnqVtyrIPQbebEYrevdKp9vSZ0Vlsk4lpjRmfCx24vqOvDLS5Wk2r
0f948AI8ltxn4ZmiI/OeoMB/54VEjZne7Gm1BFyHbLFw9hKohBuBZTNx7+WDH0WX
GNSwKNHzyCzLK+j3O+S5K+KspSOKGRVWAfxJjL/6orgNkL7K/LlpAgu/YPhTfHVm
A61lAvVu8Lvr+IXekYSlaPu5UUEMNdMaHhnrBKGdYW1cmiCN+8CdgwCrCcO/hxO2
c2P649xPojtI+Ed3EbBABnYurIXRkUPbmdAwjVG3KPTjTXbKiUJXzC0ZVJTuNE03
obbA8twSwB4TKB6Om8lp1tw9wUnYXxND7CDaKhFRH+lljxya38BvKKgrSzOoxcsp
UOKDJN1Fz8KPe/UDdIvau6DTvg+S31E1dFapFLL9JMXiuA/xNqXbaVVXvsiRUfpR
1kpPLUZKtty6fmQ0XQ55uRQuPpt+scWBvbF+y/ntVjcuJhCYHZyxStnyXjiNf76l
V7beX1Ct742n6+NoAyKzA0CWf2aDeXYShVrsx4GLY1YSrFN7YhbAxmE8CHnP4dwh
cJk+YzRTd7P/xA1eUTqLC8NtqVMlyOhvOPfVVpTe0AzGfChYyk62Ro7NSorB/iax
FQ8XXL7JP/GyF9TzVIgYwA8cp5N7XgM5e5naNRx/GVt5CEwCU553ptDjJyrn0gnU
DjivMUkkmvTdkalHHzbHPjztc5cAK/VcUVBs8V0fAcchq37A+gDBPOWrA7jP+nZD
+EhfzoohgP93Yf9AYTZ/pJs1tW+zfUn+eBvGUju6hUy9zpU76x7wb8BYPKS8ODRA
x/ZpZyPnaxvfFsfaQdYTMlZNXsLTruwY530accp5prhrtLeSGsXvSbDgoR5U2LTJ
f6UvAi3d3Lyb3/b6ug5iCq42kkg0IAGyzRZhlmS0xbhCmMIBf1Xs7sJzILfSlc9d
K5EEmnbp41qfPoZj4ascLkXJIMSKXrIuLuucWHYNFcYbolbnWIEVzhkBQPnsfBVR
4ag0kam3A7OT+nfrNVAKWmAGVdWDd1M0BNSIDkhdIgWlpN9SlXok2VMJHArddpS1
GApF/g02ObKwtRC+y7u/vyzgk2r0xUUO/aC6VRSyACcFm9tn4c7b0laTj4Qvsfvo
+F3JoJ8l9HywKLO7NpPxxaNexqUmhYagEUFzu+sTZTbR0k7Br6dhZPv9TmTsO10A
qHYa+p+r5IY9vfkXwHfaKcQhZR96zZoFTLnWBN/SC7UP/BquibEMMDt7fBzbk71X
U8GsrSsDjtGRawVu/8PgpZLF9CB/2c0dMcWtCWpWE8Ru86ANRH7jmbg0P53RenFa
vWiHWGWcJ4BSTRqn8v3JZc1pg3kOceJLQiNRewbPNP0ZP4UWRk/PRhQtB8Sy8B9B
zj+LRcHCtrlalNelObBfJdTbVRSyH8qt475v4BUDjQKxFzTFyQEfriPhVKn2u8hb
CRXnO8bGsC+ZDKqWx3uHlIQWdSwRk8PLvBU70+r424ekhQlK7uHHWzCB0riZQ2UQ
LPz+54u5hKpz3tLojt0/4/niQOuPVbsxtEDCz+HZfl7CqPrtz5GfgJKHwah93sWH
Tswy6mu4EWQOSP0S7a/tn63PfBUhGZxd6y4u7V4L9sCHf0Db99f60Rvb3a2G+kG8
ZFk9FvH6s3H6Sh7aYLEC/pEK/zuAhi5PCQKO2/+qqXyOYAulP59KKKXC2VrTYcAZ
Zet0GvZg5Aw2tp5YNsYyT08olQOwMpTAA430divpris7U0iB2zx0LkRhfCWbeH4Y
q4yoTCxP7KyyqJCbApPhqwKCD+91oWGGv35aRzRLh6+nm3vVX7ERsXWtWyAMTBkz
teZMB5BwwE13XuIbVivnTHwy2g0U262AfojMRSRg+KjbU5pjanCF83rzZlbV/lKH
44FMQnwmNET2WonStK0qH6pxyVQxeYGn+skt0s+ocD1vIFIW5VZynKK+FP1CR9mP
nVcUsszscRMiARLjuGiWlRHJliODLLLO6iZXrwE8wfVO9VScwnhQu1IokdsSFPFT
WnUUfow91r4LjBzxgwFart2elO4fhNzhlLJ5AVGplZ957QIeKIIKVK4nj54h4aDE
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23952 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aYEGshOCBNLOAFPz/YVL0JBlYK501538q4n5LbYg8NYY
flB1IfPO2fNtbKgT+SOHHRb97TYj+4U9y+XOtPTgSn9pj6+7OCCldju3wYwxVxe5
+VKUj9ToOZTnRv8AMGOpd1suz9kw2NLHpLgaPIMbC4O7ZEQj08XCf+Fs6JlXIQ5y
x2wF3CrKYEGTsGe5QrJgS98X6b2H5WtMDpnL+D/WasJ5hM7c5isSGeP7LmPqIl7a
Qcqn3AEa+BgW7EtYUOKP+GJzNvAuxVnqKjCoIrqXgj2Yil1oS5SbYBwG3DsGsUyU
NhgVRFe8xmVGYOBwo7+BW2TBtlkVPdbyUCGi2seMxUWgtNZWnmc3vyvwqU87g7vC
t06jH36pOr2emxQ5VJuiyPV+gL5FB+E3RidOppmr0s3Owozm9ThD2Baxx2fokhvS
hr01XrQE/QtcmEY1LvWe4RWCTOwd0EcOx3aQ552ryiHthdAZmcvzEAu5AWV4QLnj
5pZONCVB6r9hhOQgvbbcbzkZlSDw2eqWivrWTEYlpLevYBTL5YyFfafblDroUkhA
BsWA+7cWlUlYpsAiNn65FCnffdo4JMWf64YGChpDUY0/rx15NcMUSbQ27+PKK6oh
+GdKnnEH9JqqT6bTNRNKKBWdI3E4awth39nYLKA3TGkUlQaGxCgzjK2MeepBG2sP
/UOCSxIu7qQPjf+IPBJV8WcU2Kpc04SNacZ9vx+cZpzh6vVOwdFt9tIhXQWC9zxO
wg1eUoFkLsyycV2OsNOdZ0a26svWvqhROQFb3AMPaE6Vy/YyhXiEGWZrgY0uQ//n
xHZKavqsXYXQICwyPl1/TQlMtOouShNvoRQG9YGDinALVxYVBrefBeKEYLCPyMGf
RY97476YPd2RwSNx9t/AhrZtdQlXpLyLGThEU9GMKt5RawkrIer7aO1Oq3t5Zue9
Gnq6ruM4SnClgjAtIONj44Yr2NuqzEP5dvNFrGbWAwi18Fae4JWR/ZS1+pszjMJF
HKn7HektXhiICKU18Q8uw3RfFxRKqyFaxAM5W//nCRuNcvezgN2ympQUS1NVDegu
lhm6kgQlUh5m17PMO3B5WXBp3hmhUiWPs0HG8w4kYJ2g7SLyLVkF+4DIS+DBcFyD
TIBYMXwFVsKcUGxU0HWndy8asiUWbm17jqqyXYrJ3WDsO9CkQBHAtzJGS8QIyCAz
tLRjxkp8KqHaV7GUEKDO97VPy8oMvChJ9TG4qeIuGhp9DA7p7VUXJgfrVCVNEiiO
DxGZoioq2gzePvFRVn8eM0A5/gO0iHQfECd1eRF7Z02YYJjmchAlPlOYOPQcncew
LIIkhcR0EAW5Ti00NENeWDaORYQfUcfooDorngTqpm20XfrWRNrYL9l1ZwqTopyO
o866tywWnZDAVQDNaBl8rhHgsDXIHBnGYz7Ot0vPT26RIn6SRhG9Xc8iX07YfizS
YO34sAS/M7dJ8aGP1SWmeYpl+yM9G8NWOVivg5C+dPYFYZXjGx7xlb+ilDkCa6SP
5Rjj3WWLDGF10jIbmL0a1VEpgB88VK946PxscSiSfyVZnssrn57WAIou02ViFl6S
ru/D6ij2Yth/QRZ0j+U4XW2dixBI7TDYf2R4PwdOjIIqBMINdt0XEUBzwU/kkA0Q
8QTYY/SHqehTrU4NKPe7n94uv7mAKbshiiJEe8XkkSlgsgpnGM4YZSkgilAU0muy
C6zG1n4d3+HdjYviDdghlnCalmxahtROuCtmpFaOUB+xC0k2n8RMKs6nGc/0ALpo
klyLkA46hrrKSe7TL/vBghE+UUtQu5sib9rxmyhTe86BpxSlUjeAUCj3SLHnncdt
fps6W6aZ+m7SmcuDrxDrvczSdEFQbhxiLUvVm0DxC/pVKPtrGjBKRL7Wyulz8q/y
Mh/v4rxD469q58mTrmzoRrsM+D7vfhGkgRCgE2hc1Dv3wF5wz5MKlq52y3mLmCYf
yF/a3OVyK426Zecfou4mSz52r3zDJ2H50RFClLkiovXqjGzA5xLt9cNTOZVBiLm9
Z42SLpxDCvvoo3MJppQniBlXzCQBFPrPxtlC9bllkXLz58zHK4sIcLDbwJI5W2Dk
S+ryIkbS0PooC89RnDIPqiZMTVZ/syn+1foPES+C+ZXvX2GW6YwibIy3dPzErXvC
Sfs90k9yhROKnLmM0g+w2RKuZ+i6lm2GAQHrdaHJ7l/Y17gXgZr4aajw6AHbF8Yn
z1gGAlHgPD3fA+3l8YmxPROf8LEgo16ZJlzfX3wCzsJBTdPkW1+GFhzar0/NbPlN
HCQ4MHUtsJ/eJgYdD/vqIyh7AocbKYlItZNKhnnrHaWYv47l6gSuo5UXEHvwOzih
D5/aIybIacEr8MQa2ZSG+RW5PlRYYQa/EkpM5KGU0PeImGIxBfxZhRwXQ9OFIX1K
N0SK2c7a5VNwuB8ezDYl6ZO6jzIR9rDwpoaGniEvsC0cNtbBDf8DQCd+4IxYOoNc
q+95c9Xhi6eTezb/v0ulRfax0zKaJK0fp3ADI6TTx8wY+m8pH5iVWmDUGmNTwRyk
RgDISzWAkV404IW8LWLlw+4NLmfODSHcak9mVe51NI7cwLTai533DzlPR9eKZhMi
MaMtEOfB/k5FEQleuvAAiNNjjsdNg63KQXf/87lnLguxYLZWQ3zwldTucX1IQx2B
dK+WqLu+4Rq+TLt/MA+LVIOtN3JxyT5YM2uGWykAIICRi5nivj9X0Arxdfxqp3Ld
Hh5QnI99C8hQMCpFQyY3C+4nPuyxcaD/98zx2rOJVIMZLYfwId5WcsztoEJ15h7p
+LCTvZxXf+bTkThIRzLW0GFowWwGE91g5xXn+4zh3HuUyfeC7rcBmx8ejApsXrfZ
fMXftD4+UP1wVyyC3xjFDZFxhi9RVe5bFNZEqcjyGk4hT2lDHiX0Qx0oPZvfN6vY
Ixbg9mGq1I2KEFLJiQ9KGllUGBi4CAe9sawqaLW7ml4QPbG3oxng2FHKuMv0/T4Q
lItwc4seVKOWONqBsvDIwqhrVLTbHtoFgXkz0zVRVryIZPeOmAFElmmiy4bok92L
vitKUdFd0WWv8Qo0m8SPxd+IOfpXZaeffGW9UgUn6Y7uWLIRr5OPLRKHeVTrCkzZ
m83rCvNkcgqc0ZuQM3AaG0qB+E2lM8JbRxXNPCw1l1GG46qEfyFRopr8fFv/nEE6
qYyRTay7HunF9QWgM2q9V/3dIK/OTWti7Vp+AdVMwipT8Xk85IXu2YQeRkSVoWIr
PEyTALU7ClqKGLEP2h1LVMF5aL0jw6Gz9oYGeT8kzv/vQxfvc1YqVs4iskdJe4WC
0RPhm1WtPfV7yCDF0wxJ2lMNGcnCe+hwwq1t8fuJWXvpv5IXtSBnUtC0GHB6TtIL
5AP+iRJyfOcI3AemfjTfVFdd8okqyuR1Gr5nhprHfJEh2jLzW9kftJyQCRL3LeMO
tZxpbSvCthb1sHU1kUXy/xwh0C/XTscVNPUjvXACeUyDKFG2hvwkM+LXB0Ffz2f+
Yo+7KE/6gSaqmyCCK0ZQuj0zEDKw1htD892qPdmuOswHFoOcZVWWXe3NgXooZOx4
BXJNkIYGF01asL4NwsWOalJ3oZLj55JYBqP5kZZxSNUDSKZcJLbTJvHCHfe7lp4q
O65xhZW5jNEYXJ5onVDznHGnTCXIuktZhhIYK0YS74orjKoXPWTAIW7SB30/uktd
y6cHQAlRG4MbqUHCkawhR17j3kOPx82P0OdXeXqj8eGf68lqBCNh3xQZHp2tv0X9
iL+OtxU40xvvRRIgRz0xW95l82zGApxThV+x5VBjSo+6ylkX+AgzICWTHUztAM8t
Bv/ygaF2FwSIWpwCki2rJGZSvTQJhvOV4p7amEQrZOTRtio+f7Upzk40TxxZPyrY
Z77oHFbs2o7tMgyia9v408ZKuabZFKAlnTSc5+yCoJYCmMGgvJ4nuen+GVovsPgr
aHEZkiFAIHcyNOSl5XQniGFa9xOIIuEs8ZxDGfrv516lAwwy2F15g1OV1vVdB//+
EKwAE67YW84TeOf9L01Jm2JbiKkaDeTKgbXp1zPgMgWYOt0k0qNtPM836ynIDNJs
dPcPSWXVtLo6c1jCOlRkT0epNCiT4cvu/JH9QOK46romKqODPrgwiuyarq5NwM7t
oTlFNcZANvopXmJg+zh0UjQ0OaYg/o8YunhdpJOKQstZDtfrRXZTg+I88CWnzuhg
/ZQunB3b8B+/uEd3tXw5qc/0+3/yF6mc46yTMdfQSW9ksJeF26cyGFkN3aA8Q+WY
st1T4bl1nFFF8oF7qeqJJkz/vy2YYbD3qT8s18MRy5qA22PcGMQQgityLlh8QQve
hPNApdLAeY5/nffF0ZNPkMJ2f1siipny3g1pkBMgPTzv+JhbRE3ZjjBde26AEkzK
g600hrOHiupxSxRNWLQV2o2Zj9jp5H0P3uoCTPuMJQrJri6QvzZc2YV0bOkesYJJ
mNeoe4hpcfF6FL2VnJc/6c82VUrQ0Ex2uEK6Hz3+XRMOZyhGI1Er6NmAq/tnlyvk
vqzW5YvG+SiMHLZcQS40r9nmKEyeOm1NpNWUSGrKBdQU2/T3lShBC4Fx8Xsx42gs
HYeKZjHqI5DL3bgSOhHv6S/rnsddYlUrm+gHZMg29JL0F+NGYwNfew1eIy2psdol
+IHf0zP/vu5nWvCk4jNNHH8w05mQl0S2PF8RKpE4wAKINXCuey+qDLpcCtSLK70O
3U2QTyBVaiRkWFEfNdJKMXVpQRjr3PK+qCGx/h7Yr8zycVPzjwhh88+roLU7omkb
Q4ek33K+c+i75jzN0f4B1QN+WJFHkpHpuOxawk6P8zmzNIbMJaSxCaVjoyMm/BXb
Pfu1Oy+/yz7/OVEf3boNrpxmDcukGGkoao9RS1KjVeQVMyufMDdmkiXJh7lVWHWI
ddMCzyiQZeHTr+LELISGLMTzoH1ei83EEtqPd52RW8jdoLjaZAfwN+cIrQHp6fki
Xdf+3Nl4I7NvOLwwHiXvIQn0Xw9Hy6dy44/ueZ+qdYpYUIXBLpU9GZmHnpZawxMp
OgMg9KPyRoD6fOJF1jKNbhks+hPYQZ04rmmKtcw/88iuMvPoT5qN5TyZBhsN+fRB
HS9hj3HNRFpjVng0JkDlZTz3q/DbmGeizPYmdimUwJe0vzcEw1S005okDSxXPxvS
pV+M1OsZ2byKAljKKyna9uGWToWYD0CHAx4JYt59h3Uu5/dKKSWLD5tAMmFWYso2
Fe9ohLPlzPc5QrZWfn3yfBoLcZsBr7RpbwBTuY6kDpHCwNCiHp9LUsIETgc8Gzbb
TNMb5LdMHQU4wbZwL3KeQQq+KLcYhOja6QLtESNpEhKyUmm7UGfTn8zPGnT1PL0P
8tccmZYdkFT9V6wMR9BGAV14zWqWJkrpwxlltQP8gdFCJTeZAJH6EgcwE5AcWXsh
w7mowJ7/xw+SJXtAm4FuJqMBjEHMFm+rKhXvFvK6CxzctNZhe3gjLJASWlioxvCF
/ueB6j+t8YUeMqRDpdCzH3CxYUCcrpGzBJWCBcsSOsl3iyniOU3yu19H2UrznU2k
4Y34H0lOB9OMKSurQ+itK65LZ9Wwbs0gfzySo1m+IAoK91VWMS5zVLnMxiardcgY
C1aGqlK2re3W9zOJXkSrr4i+Pqu7FG6RNBQ8te9Y+jR25cMUW7lfvmNXRZ8eZYS+
D3AYIiRNfrF0NKSjqXAWrF7nvl8PbEaUUgzUDyG1KuYu2c4YlY26WwsOKVevoH2H
kANFgRm6BS0XlQEM5pON72NF6IeaX+Zd+2OJRszszkYHdla4vNmeLEk4J0XzD/X5
ErZwXgjjCKdSqlyic/VUIckTN344fEzo9AiuSgxsA69LZFHsTpgxsrcnLxFLe/hC
mxJirjFpuVPc6O0vCjih+xVS8dQo33sg9rDg0V2TRGYVJq4CFCVEVz4iWbZw2MlE
NhWWQk6grdEWmuWJJr+647Mnd97cdnqckca15hixXAsS3c6tQLVGqa3Mio8uaaEQ
+j2aPDm5uvtiKg5cm414JBbqz79yC+WVuKuO5kf21SZgTS/Fd0Vo0IyfCuO2QeJ3
J8BIR6tOekWvFAWqARR/l6+LgxK5BJti2/n8LMzYs2SrF7S+3lZj0wAPuMwYIQUs
TMie2/cCipwgLwP9EPPQ2Yokc/6mHu5ThGXPQfb0VKMLp9CkBNzhYdOEiMh21xhY
90snzaZbw97zPirKcMttgHkFQJ6xXnUC59iG0RaQWpMCOD+pYYuaW/IbAs4Fx/6g
hiSFGkGV+1/a59JYlcaEwz5UVBOTYeG0YJOiI82db0aCMANTdf6hAjyGBuQwQv92
X+bs0Vr2syQyCqmPND/2aTyB2nrj5hHCT0Skuwqm06IFm8nED8ZdbvsU1PI169li
tH69bec+5OpEWzKfwNXbTV9zPsruVTiYgGc4lYzaQXRvikifqANBd9vWwfiWLqM2
CDf9TofMT6KMt2QoHBZ6KeU9c7RQlcUDAyg9IEqpHyq2OYSy/Bz8MeKut4hlvHys
8v6uFTqTJu1+NFV68N9sQ8e/7S6zk8ncWakvx7F3zWIN3mwnppW7sC7EWmux3mZg
O8X5PGfiac5YrFjA+bcP+DXyGAyK+f3SuL3ffQxKEljxxKbPcU7tEMbklxt83r9J
Uli0DaUFY4hZi92QEzD/D/24PNxVvb4Ow+TAYZnfMraAaovCtlULUkdX7eVfu2GT
fuBAaC0bKddjDSYYdfndyHlwWzR5vXex/7S2gMuEkIbkZXOBKyscCQC35vv1lPvZ
CBe6xhcNpnk6b3YwL0gnlOOPaJCcGIoiVCw/JZU1O7DJJyXSVkkw59RyNuUIwk4W
MKbD+9FOcaD79vuJ4MlCA6V7KSA6nXd45iIuFPE+5sXmj3/53vKj6euZPUxuh8rJ
OiFOByvIgyUjAeoPHlnKuL+W8eehwkbEzgHvWbFRb6SQmK8VcJyf01v6RojpM9H4
J6C2qAzoi6b8gG8iHRT81BMa1xh2sxskvfUAxPk9t8V+ztvxpH2RxVQZZhV0pOJQ
2XvT8iRqALoqfHgA4hgulUobJZh0F8Hf8H//HbCLn/Q/evTzRxiFEsTGs/1Rf9YK
NA9bh2kM+MOATmiXUVyzL0aWCOCoudXpkxU1OE2t6aAaFNitzJuzjE77U6TXK12r
UPHXGJ7MIvs5kWplh4jdtH32YlmIL2XMEfOiT9m3FDIYs4OrbXQrMnHnmwZfzJ30
kDaAt4JD6CK2FDlAtCkKvK2bdOgEArs6VKwGudZ8qhDQ1MuqP2GkGVp3szi3kjfG
G0sm0EC6g8mGsgcS9C24KpyvystDIq+x9RqcXAhOtKTyfqcxgZuCArlCmzQ7Auc3
ZPQJhAMxvzVGW8O1l8SvHU0cD4C6Hb4wHnzLKtwOQVFMZ/Camtt0DGP1jWE6kTb0
gmHPA8hraAlh6X8QZNzQWaYD/ntDFUkCgSXBE0bfacYCXeYoRqyiAgHmHpnqs9Kl
GW8QDPudcmmZ/085Eu+p/gCLF8PygPufBJVLGwaVRvJg870cgzUsRJhXuk17eNxX
bT2Q6kP5OKHVqEd/+h+9KDxS5MF/mWtqvO6zDg2hHtdMTR2S293ISMBp/D0WPxXC
eQ6uVzN2N06wif9RIU274I9voAHXaEPee9dL6uEVfmZlrw403LG7HU1xfCDuDx91
eK7SDE7Ipy2wV2brzhHjj6ZrinMQdNHlzdJGzymI0CR2uvVFw+ltVG4/ONrmr14h
ancqkqx6aQ8Fdy02ClANgIVH0FejvJ0RjqmpSHWDPHmJH7aCdXcLdaXQq6ff0xgl
PtxDxvLV6LbFxMQOJeXOiA/VbTasrjGjZHAlCRnG/Cvwr7ei7X9wSmQp3FXWrz/8
Bfu3H9A1GBBzDw7LM3dZ3+PoQuj2Hriaw/Xn9DNewm/jdnta6ACvESJphcCUrXhq
1xgO0J5ycmbvSkhK9H5CYLpOKehHIaAOm+j7MsXs5wMKs5TEy9BCaE4OVwrB3OuF
HX/0eTYh2KGANpjaqjfVAKSCRfyKXpxDhJuAx7t5c8VYRmvh0e6RJyYShLQQPX9a
AHYB3mHOymXb1uX4DUwgo3q9MB3FyVgf/6KdtE0HbmCNJS4lNsE65a9dwRZws6Zs
mIRgVq59ramilKQyqIJlLHD4oeZeGzaftXYzzk29NMJLiJFPTPRTRN0qJj2QcPHk
q9KOhafoVytFlSctvF07dWFUaii6Y0br+vt+Qb5iaw2+13ogwRwJw+i4z1WQ6ruV
OdBzqP67fLWeB3TuLsdon/kjSf/nVL/aKGOS1AnC37i/z/gj+he7kO9Ap34RIDqu
1p1FBmkPylivA+f6SNqR7SMHWIk0wCtqeQvio7si4k0yaLRXt3QJOKiuGsbhj+I9
/rSdQlbNN0VVPBg0/6S3JtNhsgZVsOFNR0YuxL49qgIZhxayZNMPllwsNILH19uw
5B1sNqYT3shdOF73MM/svdtXuew2FydfNWZ/WPmkvv5mzKvdLI+gAI9/+hMdRXwx
XDqNZq6DiDlzzhkiXUgi05ak21S+7qKJOVCdge9m4D4FZctspTRrevgxR28KRzuc
YderN6kTJnpKsM1mFrLEOn7o1cnIpNz/FNOBgpONsT20zfGr33SeXp4RlTloxIgX
lm44rExRumxOfffXlk2U1v/H2CaIb7iB9VgYvNsYJ54A0Vg6E180GfcgPHoUVzqc
6zQhR+zD8dpBy9frfDj9jlHLTWsasgn1+ICeNtMqNE/FybhEeow2iuqCsFBXMQU8
w2epbZjKYkZd8cAgnrxXQzNo7n6nXZcQ0jUXDQv2N+S78mo11zE4kw0xWkHHc3Ze
nne0fEvVZzedVbNKfIHYiCbt9dAgkZLD4RHGWZatFOGfDuz8kYBZxa27HDUwDeB1
aNbll058lJr3bKZ7n3/AmYz8CLExBcObhY6nXScvKk9OUZ2wpJ7ZwrnfArvUjD5B
zYdJigWalD0TbBOhbhfOl6qaLPupwnq9TGJvwwD7g5HVD8T7ywqHbtZLrpbYkYqu
HYvwzPgeRWcdkAZURwWLqinOP/78FQtQe1gOla/4V+m5tsiD2vxBfQkocgNG1Geu
LP5XAsJcFupRfa5d+Vk8Lqb8UTOHNz3J10ymS7/koStKXd1E9niHiLE8xWs5j1Dr
8jY/NWlxcRohOMqY2WVe3gJf6Ci/t3VjiaAqIYt2/jrvRe06UppXdjRxs36pfWAh
/MfkFA3ufDDtXBLW6+5hOJ99rW3PBLqSQ8Yl+Wctm9TZ7l6oG8JEUK+Iax8fwauP
1iknGTwmWv0RsFGtWITGjFzR7aY3RsUS+FOok9PnaxTpog2uV6DAEIVUoCn8lkku
Dprk+kLZQBZPUGaIVEnUD7PegS+X8SGfKmDjjREFCcJm5RP5aQC2Q0hrTtCPlAi/
Ba/CkM9ARx9eKFKDYysHSC1x3HtOOKxjYWYHVAvYYmPu/Uri1wrbbRRz2aVcFmYY
LbKz4H8zJ6W5U3FcBALCzuCaBSYCgNSWUeF94xQQj2aP9cVbX7aPhoys/TkxJUrN
Cw1yBVr/kLY9bSQ0NiVfg/UHcfWsjBpOzoV+604QjqSMoURZO6xNawubkATByX4G
A1srIQLFv2hiKSYInjy+skA5fErLE4bmGffTOKVdEaMoAUBx5iW3Md8BKdh01GmN
/aZwbHS7jDPoqEdSElfqhapQzEiJlEsc/mz8VElXlvBdAEep6PUU8utuWdLNk9Ok
SFQnNYjvWmmKfgpzr6pkAUw95Uj6t/0G7syTs4nLW3/6su3+w3bDSvD0dLIPjB0F
MU8Ivk4H31tJ72uzd4yyWJm7DEYXGKhDttaWaOHWW11Q0bK7eIt2gnnCwrdXJ4Of
m0vBq/mJ1KFiu6IyP4BWYJ/ihDR7oxzMz/0F3WX5xi4lm29vTozJOJIrswvfYPaJ
Viq4LuJFu04A3mYJBwz6PCgREXKpR1oy6tqrcJ6oAZqARTiQQz1MLwrJUgKtezFv
QKfxgNEuIZ1FvW73lBlmEaisOlGPSdmxm0luwxdlxNRk4EhPhOmuyjrXm/s2+1/x
EVabHwNV+FbNRqWoyaYiZpTM5zspbBXHmelGWX7RatWQVFNDs3hIq4o6c33TlRyh
4VkPNIo4cgi7rkNIe/9jBqIjFEhtngBsVcqx/aYUpbvYME5TuTW9csZE6aDbV5a/
X+yBCl425DFfWoGMvSVeAbCnPKf0CoViZRe41LTwKxtRrTBpjngqQ7helg3CF4dq
T5RM2+iOFaSQFXWCHaUoLxX0RfxUe995J8bk3b+WWc6nOb2nwWjEkH0JfTP8AcpS
qZChjyIJGjGt9z7ZTDZjxMAAredB+0Uv2lU6frWHAn7WIVAKu7ZF/0n75bLmGGS+
zyiSqYTcXTI7XwuPz8TaALpRA5TRNIu37BJ9LiJxld8+AbE7bm4eZAVZZsq/lZMV
zX2Q9yFvufpETTQS9r3n2Po0u4XYdKLxkLLJPhSmaU6CZQ7/gInisOlZdQ/wMHOE
ZBaejIbx2EjOxc9EAC9Zw7bv6q39u3Cp854KvW4htig1bgpjfF8o6BDJGkwv6wD0
Dp8PtNWrmMrCLC5HFz4zSPo9OKNa1oW6AaUqNIb2qyNJgXlvUpSPgx/3IIwXwNPd
elUvreYQcMKHB2D1xgQQkal6vcv745T81VUgpnQFXgei8WaBioJsjMgs6CbrB+mb
XS7gsx+j2VKHhYQJBFtY9aClow4ViYnD0JLp1mGfW8DblsQeBiwPpuTItIeRpxoK
SKd1DxCoW5aWccN+dvVqNnbRFfEeZxgSrEqGaRTpZvn1/AhJuOVJ728m9/NDDBSV
npDmko4maIa+wrWaIqUlUYAY7ARq7QPMWdR9Uq0obf8lXzx8xvT73BuRqyO0rldK
i7xtCugfMH4K2EM0g1fpK0UqwEGf6zT3rmqF7D844JONm6p6BGv8YlV4bCW4ah6u
hMOX44D2ZMuXXoA3wxVJBX93sZF1d5KnVf84NJugq/imL9B1HXtDp8iC+DBVWo78
v5Qez1wjTXppohTyQzkLbUjEvUnDe+sQ/0LIlc7T6ex9wpV3Jjn1is2Ec69pdonw
f1YqpsHgLRhUvNriMyUmkJFNLomX/i74mB2/328XovPnQ5ron/ugUAO8y1QKgl4F
wUxPvBrBedNNLANQ/CPHO0GnQylMlehmtMvkGeXpFws3j3bbFToXaiGre8rhUEpw
fd4VzrLG7KsMCmZHSmXOzdfb/eTOCwb3BOFOd1IBOfMoNIKRq1xaiNuVHaiKtj3Q
zPkmN63iD5CLdtBVMeYMKgTlRhHEdBq2/vO0D1zqTji/hSyhILuh4Ryn5ehwZVnq
jAJ/qFvb1UznkNuokHPdawO+ECQef7bAIDJLVMxYR5u33m5Bv/H3aE60jcxOUqWd
C0rtstsS/mHXNHe5eREg53Ftrs2S+nzVZSnMsCBe6uoBVa0vc7wwZNxE/Zw0kjNz
NeMPF8oF3jCrpIZ8p41D0q32PnSra5gE42bUGMnih89bnYeY8gmdDokPEKyy5VBi
dRV7JJbtyryM32g6KvC+IRWmB/uYTR0IeXCZkAWR0lrVq1VXZ9Epwd/AtEYbJyb4
AIcd5bwYMtOmMqUr9VeDuN36+mqIvxaFvQmh5iierFi5lxWQgrZYbTXqqYm4s9za
vJmfPmwB6bzCEavHUgBRa9WE/qhPBLXUObMSQNirhHbTjs7ZRjRdPZCqIpjwGDLV
/n7OQskwoQJNUUUPXmV3aAOpK5OGHwVUQB/CoQ49pW7NW550u5oogIz2CsKtHEdg
r4R/+7df0OBJgD/p+MZ1a+2YpF7SJHLJPcnoxcQo9qlFQiLbZKHNLZSUC+rySPPb
F8VaHzbtiOYJmoU7JqWmdjHyVvIguXS1OmPmPjERwyu5cDfA4yJtrqdJ96/YSkzA
FG9naQFhg2JtpUmIw1vkOGx1GNnjuZy9hN36Lpi6wwWMC5GTZ/xwUQl3QGfWzMf5
wV2nbAI/MC/u84I817Om2Q7kj1RuEulHLkBmwrJJpCR9cgj2aDeMiqLPWDVFPCgb
lnWmvIOf4OFxO582MfWK4BYL2GBzeY95JxsEey1QWR2LN0b7HFS9h9u7at4YdnjM
75ZVbtVoh2DmRynLYZZ5O4ZI/GzTHNmgfio1oij8BntFU3jd4d4jAV5e/pPpjtyE
n2Imf8B78EbQsqlMWEQnt4lm8RufLK6SkaS0uXKPvfsyJjfDXcu2xosIgVEW+LgW
/vjNRpKJF/8Y2uyYTRdbvHJzSQPcG0runb484jwtXNOgd3Hdtf94+KPUPUnHOc8W
Ide9kxLsoNbT77HqXCem5fyRdgdJLnBnVACON0o5T1skcNLRQdnWwJbHSSuCVIgp
zKjj1RvCg2ExY7EbktdeQKO+m5korT6llO8oSyZlo7cAwvkKErtRGnxOvFKb51Q2
snrIb5nw5e4tC11XdLiNiUdk0FOhnx7PbSUj+EyjoYDIDkxzkL3gLC0U29qXn1vr
GiPKGY51y9Yd29B4WAkV5p7yJpH+F4Z9N26v+CVvPZW0Xsf3WpNRr7y7dHI2uF55
bDPx8o1Yk4QKp/pG8m8ppxrn1zBaO+Gve62/xqkI4SNZCnkY+MZLyFI3oJ1D/7wA
bJg6XwAiu1Ruhq0ahHYBYu4A1iZkghdaKforp72orQ4eXpc0NUGUzhmji/8nEh96
WH7q2WOOtRofU1+TJfGuaLsRSEQ3J6OYkAJqFY27GUPr7m7GTv3u9Sxnz4y0yvjT
bKRLPm6MCUjtgNzTq5DMeY/Ca6m0ZGeL3OXzHQgtlu+vL+sPDeGI7P2Kb26ZU0qO
Kw4Dj601xObWLn0bjEoO9+22JxcLirOEmowsvP7ThVmqHaZrfBO0io8W2IL1qLc8
thOLqwQdiZfIsZ6pq7FDUGoX5W/OjS8Uqugs0OfZJH7t1J5WA5uP/M3x407la34i
h4MaKCwpTl7OzZhXT8u92V3Jw/b+yhkz3fmJ3GvspQw5RqOIZiW5aK/PWjHfA66t
JjkEUqvftB1Ou3s4gXY8/Ly3VCy1DYmFLU9Xb5RoA/BgmhAGzONINgfub5Pce0ex
XOKbq5gcCT3IigzOWQjvyQ04+cZRz088Q0/XcUk3cbEFrTxhD9e76cR24W7B/8rQ
c7WWItaWWXG3DpCHDwojDda0wyFKtsSusb1f21f49GI51wR1VJcp1pUEcvnHDNLC
xskg5k7Kv3nnWCSvliPRwaKExsJW4Rc21UxHucz2kzrl5mRA4FKZ1PvaqoD9K90e
xcILvf2toxi3AAQVu5iT+pcPcAcO3w1lZsE66pVPf9Yv8NiGoX1dqCDOFZTkP0rZ
xWusSdXW4C6t+ifVcskeDYy+uiZC8H70LoMPgMyQtMXdrOoTh8QE1fw0ZxX58Eyi
O6Cb/vqEP+yajqTwYEZfdppIBlrhnz75ZDEw5rYDC11/R+GCZSDQhUjzGN47nRFA
bP04fGXKhNSS5JOtCKhhDbGYdN928OLv2CpXWw2iL66YviT33T1NMAHgk6eHxooy
U6vYv2BcYy1aV1ZvFlsHdFBTVFe2mXg64HhLSD/ZAGPaZIrVxW7XIp1XkjXtX3fD
5sUG+9WCQoS2V1MBjg1NdQzFDaFuVwnjfxp7qJcrv5QtARpqg+BUnUpTm3ratBVZ
RBUXZsakLwPrQAadX8+KLPDaYtJAZfzw0gyeCJ0/tIcCqvbhF75eAKCaCmQ8ZwVm
e2UcOkoJCZdtiO+W1vrc77ILCbHco1HLOx5cKZ03MRWUL1fngBRpFGDmTAiJQ3kQ
e53pwco7r9FKr/P7jZFFoV6UAf8yMv+E7vUsoKrGcLT+/NvW7wpsCDpOsQIsNLBD
as/Hf0Rd+kU78APthj5hA0o9jPuoL4IDXgsIzyGpyKC0reH/2hlVkpSrq3h6E1NG
7QZjGXZWv0pfL+XHRL7rXogBYiGjAnO/NYzY2V0exP6Km9Eo42lJWiLWlUAii6P8
S95QUul/P2Ac5js/g+6soL2Vif03UXYiDOKmapC8NGME66Jp7b5QSaGwOOdxMs5H
OBAoSsdGsVJLSbIVwHI/wH04dKJdNZm2PvLqtvYLZp9vyeXvzVb4CaXcmVMcbrSZ
zJdSZURAUMoPomMQ7Vj4jS0ByLmUUhclp0sZ3UGUFfbRzDsmtSbpYqvZSEHjrxUi
HGnNJGk5iW5AzoVNiOuwsh9SlQA7sKK1UQJw5+7F1KUdD41U8CMBSMyJ/k6a9S41
1TvEIxUrr85jTxlW2Iajo7+6D5u8oofq0++VV8Pu+p9btVYiAwxC5ebe/2/A23rw
tjNlY838hYzNDRUW/HZB2zeSi6mNUGYQCQgUu6ImKQDul20bvEYbnPtzCLq14CTn
x9U82CaF3IDu/QyzOSWQowlS+a0uX4FQxCe9EU82S8KyBtwXnwvqENqWvg+CHgZn
Qm5JGJ7Sf2gEcK1LZRTZ9AlDZafH0G92hc3XYcpJanGdjd0hPxw66c7Rl0sIdNn7
ZHseHj/42yHXZbh92V08eMuIBfrPb0NqrfCwuP9evV4CeNMWwdkbS0POSBNZzvp4
EbYcFrA6F/jPm/aDJViEEJ7dgtx2fJGGW9PzTM+OT1QKrXLaeOj7858DBGYMQgmU
0zm1ir4E88P3uNGj7CQv7jP6Cvz0lD/d0XdBtpOuG4DCcNdPrO2xVtE6GSb54aIJ
z4TYLfWvahEm5YvAAnFreKg6LecFu0qnsX7T3lY3umpf32qaujKeeq1kq6x2Lk8F
Tu4BtuAOCf55/Ykt5Z0Bx6tEQOvA/Xg7JeW5EabIT+79KVQ9nNqRR5PQHtLlJOqw
HHxY/23O4RwKxmYr/o2HuYwGQqIL0rCt1Tdu4FxztNnUJD/Gn/3/dDPIZ0ZiOSMu
L4QK6pRBVoenzvOHwSWdkXYGkpb5r3jtrx+fEFJMRkyYim3KgxPDvBk85QwAGILa
Q9UqlqOgjqWriTtyKvhYCedJNuNTZPEtiPT3iuL4r/JVk6VbTFTawbBGiFgDA8sn
XnQLXxex/SKY9rWP6tL6+aiD1CJcXxv78IR//93UhP/gmrpArUKnwEDqXwin2ktV
CABczQcheEYs3z3ITo6vlLOIdB3yezeLrWAA1tUOJ6yYROEtcDw1L5bbwictjO7Q
3dFy2VEwgwTnxX5K4ry0ZtRObgoOodFZKj7nG12D6eJ+9cROXmzBowzyohI46bG+
jX/IG9Ts5pdG3GJ56UYszpJcpMEOpBwahY6lYmRowSYqpZZVz9KqIbVrA7s3EafO
BhJHx2SiYAWJUDs6xLLUAW5p47ri7UQFHEWxFrqjaw5AerxhbaPG8FA8cxZr9dxZ
20T45gNLJW8grzhKMudRPXPz4FFDXhIfVbgNH8x0bN6zAm34cVgU+Cp4dqFWtJH4
BjsodqBgq69rGU5V8GoKrEGnFgz0Dp8SmoPQaltGJnP9lKVeDF5fdYNNHNkWMWZp
5KWcJaJ9PAXfRRsF927xWBxj7WFxft7eyELnFN1zbE1Uv4txdwN7V8Lt/zeXNSQS
DwA9WDzfw+EkV6gu1fRpMHleI9BIWgxr3CSQlw9RXOxB7Vi+QyECgBb4BsemLGIG
9HOKd6362jL5Y4662pNTDABQ6sCxUtOzZ8GPtri5sMWJLCPLvmOuMxskDWGYYcRI
+uSGU2Odkxi7tuy4nHKpNaHDWMDEdN54OBFYD25ME+PzgkWaus5rQ0JMOQZl20v4
eYx5D9ICbnHrB/dtbV5GS8opYRmjBOlg4K2pCh/Bvvyo+2enwgFp3o0sWvgBSnfd
2hzT46/OmVjPo8Gr2wQsMQjZICXmf5VvkyJcNcaIsj/V67gCUG4A6S+GUeXUGqaz
9fqHmJNsXH/NN8yhKyoUsGCizqztLMGOPQq5o1HS7jhNXVLfKfmh0JrjVrLc96go
DXVfTKCgtPhIATYcvNcmXn2IMUGogCWUhSoi0Ueg3kcI/j3cyEYi1iY3xFpexD8O
wadE+pYalW85Dh/McCMgC/RSf53P6+O4dszFgDXu5VUX9NvmgrOIUL3IsxiTZsFe
dSpZQo7d3/xdsQhv3Q35ggdWz/pI3kZtt3bZJX+PpMDAoYuhxQvfcbp194S1Al8G
S5Z6uBDy1E2v8gItGR6vKI2oe7h+PW5dsJURmf0zEvCeRETu7QLx96oYIkgoj8if
6LxgLgrCQTADI/X585AlIv2/SpeDoy+CAGupOz0Zf/89pYugZA5FM+TVX4zPCZ8/
Xr7cm5uk+4ncAjLBULxBRsbv9CJt4xSZomG+GrEBiPpZDfV7KDwAt1IU3ohb0i25
qMN1ihi5oJOcm/u0Uo540tU6hUEGqJtl0KKMPpatkTg9In8jSluh5HiFTDLk17uA
scTt5xc7XMnlHVjjNcg1NL274Jam2/doZrCYo31em4zyF+9AitDegLbIp4tD/WCf
wNWzS4soYSbHp4MpOx8tkkBW2baqWGtGZNP9ewcX2G6VQq/x0Uk9agpmPRgswAEa
54o9UHu+NBtqjMOmZ3CIu/EyCffznknvORRjXd2iCb/CvMrTXIRVzGL0s1/EiT8S
RqKjBNOm0MTFCY985HGgPlc8D29mOZLRgi7N83IvGVSBCaxYnNFLxZvpK1mK3cjl
YH6hLCeAd2fnNyTkH3Cm/dRFMbxAXH1Q4eSpAqy0hueJr7RwjVHpTu6U6kOR6hr1
Sf8eL60EMqunjk4lArcVLLybB3TfsbTHNHS81RvFhyDm+2v+OZqLZmlivTWCw+sJ
Kr/Fy2pFp+StAs0Zgpgr+QxurggMayXvS2KfMPkXcn7/tI7ERw5txc3tMxyr7E6C
ChjSFw+rmI6Qa+zZvVRUpBT82HfHhp4POLiPXTFHOcLVOeS3r3rPVccY3LoUhDja
dDCml43UBSNwbQWkV8ADSjQVeQiQ4s8pE7eJCS/q+h7h6/EOSFsp27DCdWBWJn5Y
bWcPr/J0vCb39kw2904PwjuoLyFGnDP9e8BaAaQE5KHryMneDzDTYbFiU7McKWiW
sjzm4sEQeeZs+ii5c1pnqUPTAvCFHfOkbnRgCArEaxq2B0T82YMV6V+ydJlxNSxv
4aF+MZyLTW/oMYef3q0/G3nN8UbZBVc7PszvxnB/95VlF2jvLw9l8Y9YHVRt/Imm
Xq9WbPyVL2TuGRsqS9wDjm6x9pLJZneIvs5lRsR2BS7yFdcRGadMKgwzkui5N1R5
53A5C39dbagIyjQcruRDdsaDVhrDTueBq/OtqvBkpH6YuorW7/OOqqwPiUenvyv1
qufUSOESy4jON5mXiZIgZFFek9Yb9TtTbYgwWnQjxCzH7Z+y3fYSm04MKak+4yuV
df8UJK+QEYpSlHpJQFGO+4hpCzqbd/BeYl1NZwQJNArQQyRQ5KIkVAJv3KwKwnZC
yCnLaC4R2NeH2MsiSxF8Ij3hQD8yaADuWhS7nCMNkqRh7OdeKvHQ8YhwcfDtSKtp
tm5uqdazXAc/874W9KA5x1Ue+LTQZV9FA9sTbka7/l9s/8lIsisTKhMSncYdC8zx
zGDsqUskxLaAJQiPQvRzlWFdBmMOfcKr5byakNQ/gJOe9yMy4FgtmOL3xchq2i9B
j6Oq13roA5ZFPnnqqQyNevcLiV9iOHC9crWyYGe2gP8ChTiHWJX5hoqgD5VgPxAD
38SvIu2NBJbhx3BiIEx/NeQLkIz+CHVOss6ry1RlyRdHQ3Fm0NoKPIImOI8sRaS8
ivIvf0M/nqZwOcWNKDdDAdsS0d5Olyy5lyzW9G8l6fRld9TEjID5oF5MwT8it64G
3XIOlexwxpX5s+75guYjv6MhrHQYAKmj+Kd7wcHy3s6VeYpbc5l8rQcszoo7t7ag
XMadjWymzneLweJFPuN6oW36hJc2bYixnd02Ty8tKr1vbDFG11LGce9BvkyAvTzN
+lvVc9j3O6zaBTCkzHJ1X/SFkdmWZaJ1niRzgA9a3LAsw4bjgth3dNhrhDvSdZ86
UPgCOYI+XBINz5CIrHiGQ+Vmn9FODEgvko/GpaUZvH0cD7mhcMdZvL2jGZ3t63uq
l81dG05phfbyAJ91BKr9XbxzxyNdaxGP5cT3L/FihlZoMyrZrovRWUf/LJZnnZyi
jbvEitk+RxjxiK3ebnhYbKjIRUqMDVLh7dF+dC/dHZUI03sZAimOdqXQ9g/fsH1t
H8xn1L+1Mcfy0YmkJjkoYf98mj7vgj01Ko4MuAftJFi0xEvOPxJIdQNoA0YLS3jz
cWpCiN2byEzBTellEauGWtVMVUvC1Bbp3Mpl0Y5hMf1w1YjOMLmBaWEiAYnnjM8B
80WnKE0Js07y8RM37ZRbslay6ri/PyfZlWpQd96yFRbdqh57vRdCunYaDxqdut2E
w21HqzHIDmgDc5QTg99fTa/t7CZgd8Er8JMtrcnUmvZDyriuFiusbBRjTgiW6G1A
xYkD6Eznzg2M2DE97xr05OyM5gSMK3TtwvHwwu/2XGxnsOrpB6sNjBT2+alhVl22
x82wtnrPFODV2Tu1vDaEkpqhI1cP9jHIf3hTRRzSqg1IyJwqdvuTgricnxon4yzE
cuJsuodOTZlUQhzvmzeClwfEUtW82wwzgPr93jBGJVQdDixpBGqqIbjgQQLow4Wg
r370615EmhtOUrskDeraLtfAglXawQHP54JqkimoqsdvYbukS2K4kNTwrBgA15Ap
XLgFEweXbJHZrk0c/F8FTOZPaOOda+R9QSG3tITPSR2SJ+YsB4+sVu/exKixw75n
3Ie+R7D0tb7pHBYCtJbThNUDtWgftlUQC6K1Do0LV7kY20pU/hcb87NkcsQmYzR7
lRC5iviSbT1MipZcUTFTBboy4gBXyrXx6iKVJJ58dLLAA1yiTk9B4FfUFDYRMCEb
iAChmVBfjZLTt6SjeUM3x7zGiHiykdJ82ehRr1GgAuXtmMnthoGUldFkpdPZjphP
A83OpirMMYHzyoFqFEV4ShmvRvTicCRA9qplpSbHE5SXVl54Qz0PoWUBziCcCA1o
eK6XFh8PUN4znDzZJxI8u6TEV9+7BvPFtyNJrM7jNe8vka7s5NmlrNSxar3vO3Lh
2nldnFpVGHl9qTA6Dnl7SVEv+vNb9/UZTqvuEtpKI/rU+bUdq7jS5Smku0uMovFT
tV7Pc6x3rqIohyo+53wiOTvTsos92HOMZaX5VMchf2cefEzTYk8KStszg7Nii68f
s3l1xkkWpyB/k5IFDHUwauKZEERfjZqCDFtUod8qEFK8rbXLbezcxLpAzIUxfI1W
wk/ExyrBciCvGNxPwbLPxO1JnUZ0yqBy70HiX2CxHyC2nOLeZ83QpP5UWUCK1gCX
f659btXmelm2qDceeX8RlDPG6GXctTLEID8Z4n+be/+JUgMg6VjPxo2EOZqbRfPy
63QnxvyKd9ZjF+3VbIo8DUahIlfTVfs4Mm6Dpuu3giIX9HsdL6qlO/aaxPGw2BeM
XDzTao8o7K6zu5GZeMmVKJkwxuATbYSZJqrzAVfF8aS1gOEwL4WH1odV84wug3So
JpfNbs5qy4GuSvAytgv9j4paExl6TJ1lY6Yx5uMlinhUFYvPxVFmMUuAVhPDJK8d
aM/ZHbi/rA3rPCo2iD/as7bn3krLulbY28lxBliQJEiWwYyOcUshMyJVVy+t83/K
DNs/FAx8W3hkJBVcMX1VGU7Pq/mmaN53ODpN5QropDXwUR9dXF7rvMSDkkPFzbht
ivSDELatRLuqkShtg4JZ+aVtu/xdHEsWm8u3wY564ELwOES0henuFW1r4HUcvLpG
YlTVHWhn8VljPLz5t4UpO0QHTdN/f/OaChMLI+l4WT8BBAPYPJMaEOCUF4ogx33K
K0g61eQKr/VIoedsf0Hr/jRVknXxrD4D93wApZvP88vayLE0Iv77sEo783pK9YmW
kfV0Yr+04cC16hBNT9RcCdOC34oEIU97IiOA+jXGXBwe4z1xv6mq9rngfkKV2g4B
46vOHG33TspK35KbhZtkmRX2qmdIN9cg8HuKRBW3StDJVAfxiRRl5v0smMUkVBTn
jS+rpSzKh0D4WAh3FOQzZrT9ZZ+dl+T9HLQvd02HWo2WQLZHhr5rhZkhUD9be7yK
zpO7WfVW+F6cv3Zv6ZqXBgjdW6/PdZy3Y4VywupxLHGuPXGFEaieHvB98AOPX/06
YQbD+BtvVJ5TYnRiLqJp1Jyz0XKDocBj2ea+7AHV1LGKfrfgz5VgwtXmcGcBnyai
cSrEq4Yf4Rqa9U1CG0u7MxIJ2QwzSl9NesgI+/ewgpoxuIKkpXd7RqYi3HE7hxQz
mJdr2eX5iGRYYUoJRy+0LSyEabjB4Meoi+iaU9ciWajkdemc88KstWtRa8jc+6GN
We0NbvS0gnlJ40TzCBFSoK4xEJX6USxPHyVSMiTFw/kCOxobfeYU7uWT9Y7aY9yf
XnPIanwZyxoWdM6+wNhP8O9F1O9zyW3fHBwSLjCXh05eriFJ8Wvsa3LAlGe/eYs4
MJzZrYbEvB0WEKs4siwx7jbldrKkVJZwqpgHxMxRQ9j9FD4cG39ctVoHX+mZcMGf
Sbwme99BOAyYmzSu+BMjDYi/7hwgbiMltdUMYu5W/1jIT1jZSOaAtM6sp+y2ZhAU
mGXsBfQR6p9Gg0MRZMutmQxOgkVROP18aM+F3sbmtPEM/1IrS05RDrFxV2xzSBQp
sfRjpuAZUfwst2WZHFshou3SWvyosQDcZr+OqH8M+Xr6IVKdVHh1xZ1A1pYYEz73
BPL2e2XjIFpDODzMksZjIR4+cxSvLOkxBH5jF3uPpsNxZrGuDcZYcjjreZrHdmzt
gn2jNZlBCF52a6M5fUAPqNBpQrrcbkBE124XJfASxU5Cs7TEacDyGndGNizYraY7
wpwpKynrAIKRfj6bxnsp9DgGWtO47dl2htuLxsH/4zmbLQw2PXl62iRu2TmhthRR
nOQBCUG2ThiMM6RZIBRwi5n1ltqS+FWSWWaOSYheTtF84cMms+zwpyMfWiwffOY2
q1XRtfyGio9M8Nd2U/Z10J9i84nO4BtjZVLk0BTz2D4zp7fuzwZMCZiGOoPNP0T3
25V37oqxqbeBcezbvhlT1FNtHzHVei3pmIs/l8+Ajc6BkNlaL8dAKN7dA9hzQntk
Q97cpOTy9YhcnRXl3l+vLx3gzK9ULKqE7b2XLmH8c62aFL98Wj76Nh4GdfcJaqlC
M6gkbQYvX+r+RSrW0CGb8bjSSWSmPTQCVk4s1MXdVZzYs09cUPP1zKjBKOYKFgNS
uxMV8RS8QGw6kNDUCxUOqa/AFzIBWIrmztVpo+1/MKSGzjIsJOMk/F5vrYscMdwv
ytSs8ixyrjTVcB3ZMh7KR3dF5GaFnRM2kq3PCx1Vr+enrPAJa1R3u1IYGYRWL5IY
X1UzcTQsAceY4uCIVxeW6jtSQJJwEaBoezf/nyrLLKxZOgJ9NWNVtYzZuBNBo1z9
RwygrzuZ9hd9Bt80v73+ho9UpWd99zTPWKCW+HVG+C3INDvOk4J7kAcVQtVdkH3/
88I/1FxBWS7m4xwQQbrbb0F17dSsGD5tshtG2eA8QfSAoX7A99vka+BJBURwFl4/
fDw+Qi2iKF6Qt7Tsz60XVyffjIvRjTwcsvAKuUcoHtZzL62mFqFW+IuNt9sY5kNG
sR+zrfxokKmO3dVIqkn8MSs6+f760X7aX3UZr8mxtssao4F3TvSy0LDqOtQ4TGaG
FNCwmTz07fikozH7TO6H2f+QqZxhuPWWZGj5WjcaefiAaCqwzcoenyPSCPBMzS/b
F8ghQbuIbulgtEglvqUjmeXyuUHP9yIAmWZ2NXF3wlzkVpzSAR2J9+gzx4peHjU/
ub/z4cTmRn0vSdQM+tZqIUQXrOtNQkEBpuJTuyxd4I5J6ZsjRIjdOCryME6jJNb/
p89EjJtjKso/llTsVj66J6zQKDQGHy6c83b5tVdCua9GsD9LgCopwCRVGzDXX8iL
X72z1VIQWjA7QYmxHeXL24tClDpYqDmXEoTZpYPIDxIORMRnIdwD0oKRtdkwxMG4
hm3VQ+fZRZZHeRY7FDFttMw1RRILOIVJMWBmvUhERRfvlNsq3VLS8Riz4EygKndn
8CnUGl+RTs9ZgyMFBRv9aYsbnuSos++RCJnZI0IIK0f6UtU9eiYuC2NkrvPa9rO/
vSmIYzNhF3ErAuBucBcV3uovvKxVaDIYTF9DhSdJys0OQDMo7lCqcH+FvcF/t/LI
6N/JE4OXdKw46lf9Wf3thye7GQpGM1xYNyWP+izKeSx1MYC7yflV2vIcFqDdYFSP
zv1ybapUssUHlEEOi4QlQUD8LqLo7JYHDUWkyjvlqW/4yK8QZwu79Ngs2CAnZrXa
+tueatEF5Yd9m0fz4svQyvHUce+7V1jjusZwy/EUWew/BEvumyaZr/Zj012wQtKD
0NahCf6h30AhhSnJNWS2sFGOlovXf3NxpygKQkyD0Y3F6ZrsDbpL3qhZDj9mWbj2
w6o8v+ll/Z0iAJk6231qbqI407aZI7q9PIsM1/KF1ZdAwXYskWW5rLYWB6DqCsw0
M2lHs4yHuhb1BKc2nLzodVNnHZGjGnb7sb2PW0OxpsPQKuk8lDV38QLHOgHc2WKT
JAb9AJ6hKcY7NARif2EjkDvwx4t0397WBDQqf2/Iq7BObr8ffxuHqcDJcAxyJcAU
jz3pLL27pHRHBODHUCsvwhWFy3Ynt28zmYKfKs9mipuh82tmTOA2RrozsrLZhG8K
U0UX2pxgox9KNjD8n8Rj8MNs15zuUKw+PdGlbFuSbAdeDIX3L6+GoUKF9Za6EMv+
DvzkT4E8cL5meHMN86Us6uMFzG1E9Lq0RMrbtrfB+j99lsSSgoOr5avXu0yZpgpJ
m1nSZjS53E1rppu95N8tSxx6gVMV5noHz+eQPRyCFiZUwNwwMSdnGgNq8DJjJFkX
nKKFu0MDFvcAwQv4Rng3rhsWananbEJBLU51TCnnKpl8tzPySr1clNXMGrgZvNza
i6FfEDc6kYp0VTTCZaqgJoy04smXXiWjDqANFsX+mjJE7VgSg8ssYcF3nnbwxb/e
gvRU7BGQbgPm9H+R2QI4Cl7aQFurocm617OA3G88DTo7iQ+LNjWEAI6snlOgX8J9
2YcUgJxNATuLfn2fJ9zF3WvMprTDyYpvCvsSYrpx8gmfDIy72smCrTyJjROdeWgs
aFKHJdmiMSHejxYju2gYNqAOWdxT4Wd6hSkX+sAiPREHcxOuIxm7jDM+leUPilvm
fOHXL8hJhYWAthZO0dvon2pSog6GIME3182GlpSznaRapPEmDai1Res7ThkbXXMy
DXOhB2IRntRJ293bWUr9ieiZcA/JoQfzi6z+Fnfyip51JvTjQjes5tQxWZvbUuew
EJ4ZTlrk8cq5JuArkvDbqIGxxyDf8dm6dmKPofXDqlnsOUUMm8FEnt5xD7XiKY2t
9kE1Rb31J2IYrfxiz04cbKu4++UNLe89E2D+T6QqF79+0Jp5daFPEXufwx3Kdwyq
be/ZAoFPjaxwaUsfflPuof3dVG7EJpNEgA/6XvMxNoFcRwLX8ygHrziM7SvknZNi
k621f8VBsULtKGOUrlI0ooJHkYa155yZWyRysKmHl/lkmTJIktOaTBrmCK87jjo5
nk+GdkYPEp9kIP+Lk5zbnaga/IEsZ+2n+M7pJsOLLUuDEjkuUGGilzCobVRWK8qP
LHRy0EHdVWpzRVtW7od+Wasx8OPvwevzlrGhp5fqTxkw1QDAwI7zxcEn2GsaR2XA
UqYcjs9Q+CHDzg19nb7lNMY7wCUZEeCHyFOlZ+eO/1CGerOGMnVk4XeMS/wKnodh
9KGNIqLRsTLQvEKAIaYlmnnij8aCqdIA1jjOwuFlz8j+7lmtoosye8tgJpnBY6/0
Xc36H1YH22K8MtwewRGoWMkgF49HKM7EpRg3RbBGMu0KOY6X0547+aRqPfufzjbR
6EE43tFovdxkoRnN042a1m/yW541InPaGgNnwP7o8lWgaCsJIavuDF57Lx2mug67
Mjt7FyLs5DyI8FYz6pbZ08DSA2hcOzkjCpt66qDOenh3NsvKljY5AIFRm7moHydB
RiCvecsaSHyzRp/O3/7SpD+BRED+pN5+3fdH9AQhujKUcXq+ocVJ51D3/M97D9zj
wiWIBDdITpj7M/EsGDZu8z7jSWmLGc6NAE9RNRV5jtB8sWB9jMySAKsayKJI5EPA
mn+n318aJUrbQAGgcwd9YW/WBVENaMbSEYxiNmw1TrqL2KQT837a2wCLIygnEebp
86yjeL8r5wTlbx8NiIa++fOBVH6GmGmApJsjzWRWCGWseXgiw/PxBrtpW/xwLJN+
+/mrxor1duN8xa0Cj/ZdUiUle4SwQHKc5m5CAgXDQAcOssxGYQf581qOSPbyHwc9
RGTGesa7dT0QkckN4sL7R1RAkv5WuQpM3mvnkY9zBOnI2GYI9gKae36gtjV8shxG
GW0zMGeEMhOOO5ZrEr9EqEKNZ7yO993sS+oHeOp1bT19C1ufTMNehMXQk9ePQcvX
ZOi2N/2zuvf7ajnGWIunXLMZnSCdL/hriBllonmohvzL8S4Z9HllV7Fv3i9jkVO8
VGqwG4+U2nG1Kx1vZt34hSGL4aT6tdsLf0LKdRyoYrVnqRNfD+pGH8Dzp+BqB/An
V9StMM5aV4GOQi+ht53lhWy45zB6rgofQq5l94hEpkv8ER3MLnEmjzVpjKQRPxqi
sFRy7fvo+oVPOVBPJo1Taga1qGf3WVdpufhvZYaHR1MoL5MUSS4RI8U0u5noMrSQ
xMRu/FX3d64vFvMBS94S5H0bUrwEJ9UK//xtSENEQ4prvluvbziMmlXF4X8zXn3L
we9X11aFvZCsKyTbrXlBji2/Uozv/wM0C71sElyQYGyUi7pZZ7u8xyBkhVlNEX0j
BSV2JIzZwHkqaG6V8GF/PmD2pL6kd9/aNa85jj0zJis+RxYSATos+oZdjq5A69yZ
fqqmCNgBH6sLp507PW5+efM+iA5IpcosExeFrrhpF8ziClem+h3vU0eayb/gf0YB
RiTdBN2ZyaBE8D7jMkUsq90w5/bHb3pe8bftcKqhYm4TJSrDgMV+cziZ65IdBEkl
C2FGMfDcxvPaxStiHJL52KPN5ddTkiptzwK64Q9iBBJJsRJaVSYbFayKRGZJkD54
TXGu0kHyAuYW65i1yX/UJkDhDxbuu9rTS9iVskJLqxfp3+blVkz3k8pvsvEAU9LB
5gom/iCB+Z9nZgv+nb1kDcQCq9C2HDJe2DRC2pF60UkXynDMsUqOd+JpaDd7PtFn
pwqKtP0qYpBP3L8W/aKt6iSCox2WARdI5vYyDIL8XKT3c6QHe7XQ7+DhExh+Z8Rr
6nYas3s2kodEQ0D4XY8Os5aIg5y3yRJuzhwGcw/oDZa5qCpxyxeS1wXfMEnTTIZ/
KrygVID2kJDebv02Ac5SoGP3TkFNJny+6wKQDXbMI8IaNXF86FB4d8bqJCxFbKib
1znW9QG/99REEkkbFnWVXnguVWvJg5MXMTXsjVS7VtazbZ1Bq3rNImU7ZJ0duete
O1xlnuv2ZTsqmY1+Dmr9oEYcJ6jj2ZY29ELKPv9bKhSo+rN2ykH5sT5L7jtkcD7f
uEPUqCMFIxoC1MqDMU60Hf0yDpgHBHMQV+wHFWvxzCOebddVuffLuamABlm4kEJX
Q/TxFzyWqEuAaxGLURNeJGatRUNWumABYhVdh2pfRsuhf8z+DxkalBDr5OT8rfZ9
vtKryAKLo0L4P27szfYDJjMEVv1cNJhMDMg5Aj6X7t5PBWjwAN0HSNXKaUO+B8Pk
la2srIMRk/hxBGtQlS8rnB6cjfHV5YcGSkLQMBl9uwnbQGElsQmZdm9vI3e0AhQN
rX/+YtrpahQ2CpqVgY8JHveaJqwaqiIYFcZeGUoyhLO3yKGE9mjsD4e5pPJtOK8d
puuJwnA76k+6+1Z0Za5vp7NHzIVtbikTjBYLg910LOE8BsYIsUWopUGn3EWiY/oM
0S12n1sdCmMddIz9ogVEK4G/c3hWw4SbS+run3u4Rit6dUj6hOnIWM2NSS2Z+XKw
3YId5U1fk7z5GGVYbIFgAGGw9HXYLcbdr1FVMMvipq2reNa7YMdDWskSOLqZH/C4
n51oEgylFyhhjDak9aNOS67VF+i2qQmSICEd3HYR3y6a2YbZKjgayaHqh1yJy7mH
flJfUeNSrsVEYiAHRg37RvqaRhHGYLfuKRhX7H2JLC/jf0NOB2PtVgDRWYbh825K
rNIHxG2Yh/Bj0vmR2pCymQ+a7cRmHoFfxFh6QL7sOcKlzQc266r2Xo42Df8YV9WG
0nFktoXMMUqk12DsZdH7a3muwsR5vTsbyI2qkWLkjPC0fF+68iA1mtjY7/6SxQ3H
QdFKMjiEMe8aC1trKZs4gMrpw8OrT6PrBvK8Ux6cEqcoFzUVM8li92ZiPsw/UMXu
8rd7wUAjKfNEikFIXFlYvrDNJVfWpV7jCOep9HxtdehM3/RhKWd3sMQoFphVANC7
M6gD0zKEp4RkvlzNYoiztRw7v5rQdzKGc6QdTXV4CRRIxrm+sEkV217/1FNNzZ9a
liW10IGba8FvlPe5USQOGo+Rzx06Za+ww/XpyJM31Hqjw5JbV5Gjj5cmZV0u+6ke
P6zatRHHeLnqeLHp7J7XNQyXwPiI0vX8F7aQgi7xZhABv5LlwQrplXaLS6Jtrmvk
bTX9rR2mFrKZmC6lwZMB6gY/HFEs7ixCVveAhMnN7b/mTHYPGP+WzUfAG4V1eJFD
/yNvAeW6kMu8bpUQ2ljecHZjfE1UnKlYueCwXbSW3W8j1q/yiqbyd6fR/VtpM0Ke
t/+ovtq19eUw4NKWoKBExdoS9J9QY9ZQPrkx82xKDtZTyC3H4TCGtHwDHpihdVTS
vFSGTr2b0z1KctJPSJBZ34qm4K14n6+BJ1aPhvrpcwBunsKJo00ETDkzhLLtSiqu
eJF3laOentdUPVUyli+x+fAj+2bv0ZnJT7OeH+43Sk5s4bd5uH2hScRXH++q0S5U
HzIkkCr2pCmaQQ883iOtjktAE7bHX5/6P7oUF/fv4NgvzQtb6RrgKShOzIM5PSaA
Qcfaf/pE/s6kn0JrC0K2likkLNSLLCUdZV/eptucSBDpCd6ElBgDOTOEC2sKYvdN
4K2qQJqWFt6czL8FyzOi24xR/yRUy4n+YH3pwz9PzRTP9A2jSBZCv6FQ2Xbi3s5x
jx7f3t5lGkyu7icI7ofis1w4Ju7BMNxm60deGFWudXcPu/hdqm9ApKXK6fKRqVjM
Wm3V13SL5nR7R37iPyvonxVKsl7FjwuSyQ8YTiacUWuyj0UnAxeG0rdZO21IOuw8
jGpCz3JLlVOxq8Ay7Ils3yalb0GC0/JqTIz24vzFUJYeVWi9OAErztQYF1Jg1lM9
DdQbhNiu0OOUh5QOMLc5D90jCEHfdqgE+GVUdGq6v59Dm5wQLbwXL9NT8uRHnzVv
huVaxwnlQ+sPqL9p+UgR6MfUkG+8jdQrtSd7HcZCQCNVnwpzY8CYa/PfRjLh2dD7
zwqAC9OV4COS/Eb3dZdlbobHSEUU29+8ipVtCq1s66JQmK+h6n8O4YkDOLAqSXhg
lMzhdseQX/TsA8VxhhGysbtwY+4tKFF1xO5s0+gyHyX6p2mhbjZSYT9EPh1ssHmt
L94y4HYM2zsMcvGOvEfZHLCMZTsE+qtVoehSSxP5OfOBpulzwjdwi7cAZu3js6tp
7f+OTM0UQTJuQjqsI1UXx10XCx9uSMKowv5OZrXbKH3g3rL4ou/a0W5YOVJe4JV1
V13zLP3vB22WxRUik4PoaZ3PNk9v2GOF0qKIhvgpQEJvS5pR6jB38I/TPg2jmPGM
48l93s5hsN2vq4Wfno5vP1hCpzkirW7K6qoVAOLIpK3H9CsX9A5gkJtH9p30jBK2
g5LAvqsNu5CKaODBfpq5JoIlo7e2xdSHMaNeKpESKtNXBBja0DpVAXOGLt1e8x4Q
sE1Xu6e0H6UZF7TrQ4R7TtGBtdH8WktooXCXOiU9wDqXYDL6DphSk2K2PxcSFY2+
ZGNLUjXhCVRDPmI3DZnDG0z0Q32bG//lUw8C43ieMcIEoqYVg+We6b1elHbnVg3I
cjYL/WH3fWzdTzP12j9oCZqRrNP/ht9cQU+GO0a705aQfSUBkE2fqDSMYCYVfyD2
UN8V4wRyCXzGx4h70C2Zn6pfux2fwE4XBSey3xkeUhSjB+7L1+BlIGY5OYwOmJW9
iIb5YS4THMVLrFwYnEariThEjvQfVnc/caU0sKSNO35JFbJ9tXNcTx6ci6KHXKu2
9ihfjlwfJXbSY7WooId7zEZE9iMVvK3A4LLuS5eNi6xoxyFsd6TQ7SXVMeGMjo10
EP6M+v7h3GFHX94Q4XK2mb/xh5LbRWoKoTIL0RVOGEPAE37r9GgvEdtnPgohk9Zn
wgGzpupyMuXNVuc2jMlTcwOvZeZiGUYcpNq2gBg5e48lZM7qr/LNaKldmgQB/0cz
WXXfF6OOIJYEMbTNLje2lZJ02Qu2IP7Kex8gukurF2OkdH2qKrGGu6VkduPMGAvc
ZrWdoVfjWh2eRzgplxwAR4Ugx/CheVm6V6itugA4HlSosttvCbF/pM5nIf0htjFB
R2hBPprwYe4uz/hgSPYbmoS0lF1NLlGv5vOoCTHkYnPvWx0JKCclRTm58kNKlyn/
sEhNQmVBoiDeIXBgxdOoJ/HZoxFMgCOr63tjFrLAkJNjeSuvWof/Xs3ake9tidBE
rrpudEh6Os3kPsYJhIlWY+EHz9NOur49nnVOneP5Vm348hlJztqtcyFFu4MKRS/l
xNzxFFGpZKMtQUAB88dfMeNAut8HGXDVi9bS3facvbh5hOjJqrLWUxDQWhBLOZLL
yY/tAncFputHTKdRozTzkxkq9wX0WWawWIKUuuy5jzC297ntsje/39+oqYC//rw0
DER37SIitErJQbyNGj0438MEy/5JQWRBS4OwuZTep6pweAadMCUfys3Pej+VXLaI
vYY+LSHcPbK4t/dij4zfVHAxFE+jyPyHWVbLJ7+GuTu84GyH7V2DZLcIjuX7k0OI
KfI4zfTkK1sVvOHqczV8BRbKXvZQvv2BzltgCSH1vV4lrbey4OnOaAazmvbIGRDJ
X5hhpbkNmKUsQYN8TvOJi7IbpAWBiW7UEhsQ87xq4T/wD6tHeup42uk29Y2NbsuB
KbJKP+GhnkI1Qm5YVGIRLiQUJHtDs/B5tDOwt1DZB+ZS66OamlPgO4oIwTq+nsOc
QvsvMCLCyj6AvqSBB3y3qA2SPj7zjfOD+X6zQU/P01HRkEQrb6zldHp+sLaPAGol
q69/QZTti4atf2bChzGi6TO+vtbiTJn60uomAeIcXU4oQzX1EwVAK64spE3IKlsf
+SOmv5M/Ve4dggIED525BkmCUfzjmqj1D9wm+jDZgkw/gfRxuxYHZS1k5WSTXe2y
onNgcUoLQVYfhKTilhPTo3D24+ZiSEf7uFiRDBZxqHPnu/9EstoHnxv7yHGSSAB2
p3yEC8EQdmKPJnQ5rtVvOvtv8yOh8yOah8M0FTYs9JtdJDgO51WMz5xcNOBu5uzY
bMSTp7fPYUWUIiqsc9ouRG3rA4l0rO5yW88vNRfxkDClJNhWf+RtFp7fXpKH1hlz
G8TPWpU2pLxDPUrZYn6N3nSu9N616mAYKf1oqWz1k9jClDO0lPVnnPb/apW+BXqB
uTrfTN/inGkbJOnIa1OovMm6hZzuxQo1ekg4snr8iq5XT9ClUQEkIzuy6YnjB0aR
PEe4AYHpbiU+sA/zJ6UqOmI0rgPJrfEAJsWioTw4HMRJET8kwPn5XYOdoCZuoWgC
6PCgwvE/M1qbjxLvCLrJBD5GmbI95OV9GtTIyRzRpiURPfE4D1pUa36sA5R9OOmG
Mh13dWQf5U+QGRXNLOVgLojGWEC7CBCyHlG8YtxyR7Ee9V6gwjC452vXsL4pPk0n
rCZivhYJBEaj/aqeOAkBuK8gYNj0pdpdrl6KHuXUyW2J6rNT3OdP1ukDIisZWJfW
RVPTyKFnWgYwGzujvzimB8IF0nSh6arPl0LHTmchU8k/lvQgDSnXjKM6Zk9qN8bC
0k9MgHize3ISjZ2HYDRt+Fayz+JGIkIo4oDLvBpwrHD2RoMUTDLgXvFrs+AaOOxC
WqwPEQAGS/vmpF/0oMMR02GE5eQLgBVQuk04ZYzxPmuGQetnRMTvfxMGNxSgrlfF
QxCgMCLscPokWLSTQv6CdKBpB8b74m9r6bH+g1sIdJQe7yrXDz5OaakuySpFM5xY
XE1vzdauF5Zk4aFO0DlBuV/Yy5vKaroyo1eI0atAAHJYb925Rq3FRoiMSrPUY5eB
uyp3apXvcFZA26AISyXnWo2CWW4QBEvaKGW1GW3pvfWRrAnAl2YL8IZIuw6tKdd6
HPkH4I8vf1aa2B6rkqovTn6zgILh47wsxgJXaUmkATpxxsxibpXOprfz76uHhpJc
zJHb1Nj1LfHQwgDrLljGi3eRxJ79dEdYeeEJkB2ArZw/oZ2FMPkh2Aiox0Fhur8T
DSlolO35fcZW0FYcwmVu4YBQ8BgTS+eCLvZFa1XwrXukoGFByKR1ZFWBOemwus1n
IAXj3xtXgJvHqqxa93K1kIwEYFTLzYxJ2U4cVC77HYi7n2UDuYibnv8/McKwm3xa
dGacoTm39zNwDaypesA/LEAdFfNaeYU1UrEYVIaaLjdOerEvs25ImJwEk3qzb8Mq
OTNwrqX0JOVvYyUEpRDwB/rGHwPsziANXTdD6eObwMd0C2LcywPyX+R7Vgf/z2Ll
Y3lI9/B2/x0OmiH4g3RBRmgnqti5xErt3fQSqgBYtNV+xRMzoqE4xJVPGWz6LHPZ
/uwfoPHiA0CBl6jROkQ+F1pWGU5b2ELRcqhPbE6CQlzF2jEy1PIhICj/WTji6EUS
03xN+yzEcB0wem0YxCYMJqOxdsyfKWrFG1tOr59bvppzgOzl/RfKb4x5DU8BXOWV
m0rocVh1qN5ES5br1dwi6b0qEJZdHC8ixHs+L0EsKawiOjY9+gmKuDlaQlU/1Mqf
p6RAwvVZF3bNh6Wshm0/eh6rYDTEGqZWiZHSC3kuSIzsGljqLK88kV4yzGxyAecE
/qb+9dgH2RMkwN48jMOjxX6mA722NkvI7Dsr4a4bRaOO7eq7fM881fah/p1mW2zl
477f9ZxYZH0eiTHKf/POcj0TnlcQuoLsvIDSjvyEamikciuwi0Yn1axTG7k6cAfi
zZvyrkhyLzBPxOH6laxMLs0Omsa1Aub3gMOuI6vRe4u3Qayn48PyolesYaW0UUSJ
vEPNwT8TAyi0i77qS5H0E8XfgawNrTlwE9Nj3QYTj1BbJUNO/CYrHxXWCf73tBcY
pA9ye3giu+QIJb0/Q95mdabsq/9iOSlloQBG28PuH9K1H8/vRCHMZjJET9ojK+xB
LKBOLBYKNuTnyjwzPjYcLZtatNIZLGsxpvW0tu0a/JOSb5kDXdIknnwr7+vOoNXZ
Txa4tB8iNjeZplwh6eVECZi/k5LupF83Ma+SDsePyRSU5I4TKbO3Q2I1K6cJhFJj
sDN6kWA09yKR0BGiMnTZs7VsVCslDaD3bVq1h4NbFkz3PfBWxlODG9C0EsZU6Q2i
aKTGsoTutjGwAS0l8aQXO/wD4lent3l15XYzScjlPr/3xJ3inLUOruYx8t+6MJ1k
R3Cn5+zbPCLUqluVLaA8mi0lUWOjEQsPAqwsxjIcfrxgp36eHHgkEpj4qd3BhWod
OWU4v6d3zuoYG2XJv+2va/MzSF2e84jwysjFwf/VzbaYGIkOfHtmQTgFeEUW8STD
nPAZQ53NkcvmETpGR9S6TmDL54Uo9avGgZpt5caYj6yp2sJGFa1XXiKcP62yVnpj
>>>>>>> main
`protect end_protected