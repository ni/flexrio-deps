`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6288 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
EQKoDAcJ/8QYHXxJAKTmMAuY2EPrjBN+aKyrS3+PdYCVoS7Bxbt4cOpCfA2h9i/C
9iY4xIu35ORJY9Q8a+tid5JK2qy2SKoL9irayJAkxouyRq1OmLdsJ6U/s2OxfK2h
4ypVtc7XdTCcBvnXZix95mwp3fHtyU3NyJPY+p3Mu6DkRe0PeUNUj22QuwubCycK
rD/aCV6ADX2LNm3uHUWkQvvJkJmEoTFD6Wx/M+FQBUkluh8xzhMhHIxHGzwAyeF5
uXUrHcNfo+Psaozl/96mqSs900jG7mZi0wFXwxIbN8/PgpLAdlsCd2MF8Cs67XK+
HYAd90jGFv4JxauLYJoPkHjRIY59XHqhBupaEVe+jUGAPlRwLGwoARePbi+fP+Tu
S34CxFNAXQEIJJmkF4cDRz2Jt5q7XVyv1tBO9NuSby2bSAIHf6PVLViaIdv6sI7P
P3aheTlJDE0vdAUYXx2zgCBZda1Q2DXwPVXaF0AdoKpuaz5Vpo8SLdz4BJEALd/h
kyIbXndP/9kCuIxppoohsE44DDqiTNIfB0ViCOyBqhqB4X/lpWYdWrg9ggR++RoW
7LCQe7V3PyoPLW+VgBc++NGnH0Io683Z5jzGABHHC/cqXB1RqZ/3Ue3diITEZjzT
W4k7jlacbv2G1iePZEJN0d6NcxFreIaWEAM5SoJhuJOoQmHd1gQlgv+XUSo3k+6S
acaBKxUfBwTypHz9kH3SIZRrXMLt8TiY9AQV1Tz2sl7rFh6Cd64GMm/kkI0oGtSL
FQtutC1JWcEY2wIiy2VwhtZz3QDy0PozEwUjkoefqduuytS54DkDYu9qd0w6IxVY
eI54nfJWbHuapA/srwvWN7CeK9I/q3QUEYQGHgiPSjmMJCM6ulcimMWqZoAeo2l4
jy9yRCwfBaP5K93nC9wiuGhyongQQFvl5fxmGu3iMJEHFXgNUZcKkkisbSbHqtmH
Tkk6bqmCP0J+G2+X1vm+X1lwL0J0PGQwcQV24uMN0OQQM3Md7FzCU3TJnft9a3Yf
UUG9BiCbKJb4pOl5j+4g51Ey3ikG4ayeceeT2uvJs632sxsVVZ/PTRzD2ivvztny
rLIJAxYBDFD8Yr93jGahvSzb1p876Q/m+M7f7xrHzf5iOclvlg9p5ZCjFQd47sUC
STjAuTHYaBM92SIxS6jOwPiwSn9gZW6bxcYgtd/lW+zI4LcF31Z72lS5vo+801Z1
0a1tQMa/NJ0CFPBBG9BZckfzPSlGsi8oafeHZ7paf7tjgu+wJIZwx/2r5vlJG6b0
w19pyN4sEYVQpE2Zz4y47N+0tqLuBaG0VZ3jNlhOqV5qNZFRC+pdUh0DAIbRhPfY
GIexUnJOuA8W4gTYyN/yHcz3U4cvtKBcixysSqtEnVokTFpDj1ZZAs4bp8GpkbDL
UT95MV33KIvkTT8y7L6sMKCHZ8Nmnr8QU6YQkwv48w7nQbzmoT8D2PBrZ0eLm2x3
bkK70bDlXnWWR8ZFOFRK2Agl43D3ofqTtzrhxrV+jGqc6aRgOr+zRxOJCJe6ifc5
BkvazGce5rTSw05QzTIb3wJdpE57zDkYNB4fGjSZ/9S3gXpAGAHzrCA08b87ZHkL
kT65cT4eIJ8Ljx3xppJSUBJOPQVwzG5hBp6hOdiPTd4crkZpzpHtdfeJWIc75pBh
VVJ2orzocjDcQPhRdJPNmmiy5vYlwRliGvdW141ERfFDUR+WLRp8oFEhDIRZPMlj
4oIFrRiAXDdyeBS3lWeQ+BbHV9xsiLuBcCHz43vitDe31HU3ovp0SWgQLhvKrQJX
qu9ZxyHjmnScdHg9l1p9fbyJt2fVfHOPh/NsQxgfuD7v7UKp5Vo/am4a8jnrTbLF
H22y4S8azPg2+GguuClwe44ZLLEq/CTsAGaOR3rRUvM/atBcYd2tecd6ECVkJaaB
evRbzOFyp9gzZoWRsH5fPeckFw61VON1OYueoOaTM2O5vacOwfwY0BolEFEgmfto
rXM5FQFkYM4CKsbLNU1/CBCKm6oh3tiNc9aGADT4R4gzLwPMjlBLPO6x+6vzOsFz
u1pFa2yJRsAuou88WLd9HlM5t/PJW4B95gFd8fiZgo9TDSaEgd477GMQPvJYCkVp
2lxINXsU8LMO5YN5upF1573nZnN1kU+aHW8h1F85Zq093c4G+Uto5zsgHPoADIv4
uXDP0Oy1Ff28MqQ2dCTaqTbEaAi8lQvM8PqDaPX41h/8LLVl8wD1U3na++tWvATw
v9Nki8eZl+BWbAMEwtMwDz5KxE9w2DVoHraAzSso1rg+iq1h58IZz3soppSlgEor
avJ1Y8ywaU1W6GyuscdWYNkzj27DqENhBJa5wFnA3IO93w+zhdr2GjkDUEp7Hsyg
jigd8WjPo3oZnvirKfqqH/Q0a6cEEtzdxC1YpHr6uO9ysdpl/6AmlzHk7bLKdX0Q
OB3SBBRPaKV15ETy0rzRUrls9814Q389CfZbG9Jz/7zcDYnVYHXD8RnQRxQRD9O/
GzXQFTKm65JZqDoNDOZwGc/wN+DGH2nVQpjKI56ZfsBNbwHs/ABgTqCKyza/lHJD
dfPT13RQ2n4MvFz0eiekNx+TKx7vc4/1PG/hswaDii/0/zWA5o8hW3hEE7zow1+9
PEdcsdYNGW8PTPsEvBB3PW6ApKZhGRM4tn2u8csXh9cqV28KGBWBcsEvi0enDMFt
aB+L3e7ulu7kFoxUpIIa3BT9FyHAH7+Sl+1aJDLfHTIEy2syFMFGFxis09CUrbAN
8NVYTpp1FCKm5c45kUhneOY95F2mSfQjQ0w33rIY44I2QHUY8Rh2xPCDydr7CpmN
nRvKYmf1J2iC6rpSPj6AdKDfddd5B5ZuBWSs6L9AzRyedkOLqaEJeL+AawMo0zA1
ZYQLvlaz/Eb9IIrq0VNgduH+WqEhuancfDCNR+edG98/pDO5+seuj9y+ON1ozdnN
DC82ZWmGIv2e/dBR60fUkKGfDU/OGypvasQwdmsQ7mbnPHbgmGO0ym5QM7EMBKy3
8SezVmwaNOQ/dQFYrOi48t5ZYpafwbvhS3fHZ1ret/vkU/pO3BHtfNQBPIdFjIOL
OOm2nHivquUURqS5f/OYjjyol/NxXln7ZJ+lzQJjcyQ46y08RlxphGhl4qh4U9Bi
NO6pseV2g20prfdo2wuRU7TCeji2M99HE6BAIXa0rCWZgh2r6qbNVT45lh6z9TsI
TMImndmcC5EzydusKGPywe/EgxSzLV9Bp5YuFEGZeRYz1w4FwPAi88foiFS+pe4+
yLUpjWMvtrqfIR/O42ucX62eKowDBCJTRAhBj0zgqmhTBi3irnQfrLbCQiNGY4DF
VZNWh3RQT9NuRdTv5VvBrquL3I4RxessyTS1f1g9Wj4iSY9gPhw+yFJqOP5MvsD2
KWC3aixzDTGfZt1WlWa5X2aIaIMghi18k+ZHgoMNBHEmR02KOecQKRF0JsW7eg6T
N3TaeMkadijxhTLoZOm/Y4GRkX9/8UbA9XEA6TKYiZulLVbdYdHgdF99ym34G46O
EkNO9ycTgaX+Mek7AheoX88zm+fBTCMt75P0NInWL1Cs4WnoYbuqRZRO+hesvp7k
QkSbR/acishjCX8DFMs1lZ+4X0Gn+wRjND5tGERSMfjZKLRumStjUAS1htRmRjuG
ml2vyr/5QV+QuiuzR5Z2kkJ0vyz/ziiT397oHPKrjc1Kaz/ppQe4wvcke3fq/X0n
Yq68QSFxOyXqR4KaLOGPbsEkejuu2Zdqume5eghv0dmgBsFB+VcfTdJ03gLG+fpi
OygWeL21A3ALMGdeqjCq9BEj75FoVeWiQkv/BKkewZ0YsKRqXOzUCJARk949xV+I
gQMrBh2kh8yOyMr5mJULy20r0RjqACtPlGniks5Y+5qVuhMKQOf+bXNzOL88orLI
FPbMPXi9ASTcD4WXxc5OmsBbKLo2tO2GUpRtyuCLRNL/LsZgD1IoH0c7Q3OszryC
QvyTqatlWfvsRf2fNBZNsqAdbOrN/5c535E2nkBt4x4tdYzHU7EcaNZBMdDrXsey
Yxpa4zf0SiGLWnV6RgArDweDlFKc/prleFl3vg+4nSB0dez7ARMw5KwAw3jeWNup
ypjjOcHZFb5TLjGcRbdLzyTDGfT+CIHYy+duQenz8BZDzJl0MrjjH82LJyz/S2Vt
DxGXQWyNgI6JW4lp+SpdL6gMoDJrKkcw27Lua9VnAXVtFnoR2uVow5bNcxMeMFao
xgK1VpF3ge+xhmea4UUSAp7ATh6Djh98jgJCR2fJS6O7kpu+qprP+H4WtI685JzB
9pKrxHj0ZcdyQJW5ZuopXjC0VJnWri/B0v74plnyUmdoIJQClGzTht4S9KdKAKvV
Hvha3/IXN5Z60A+TIMxzX/+Ga0or2ah1M59Y80HLEIaB0BjsYItiGlP8tcZv10mQ
zkgIC2fMwMMrYc3rMffXYiic22DR3fRRT2fvMGGD6bINefi15T6Nf65bnTxPypHJ
Bs5jCKnsD7h3p9BFftgJnrmfCs/hjptEvDBvd/1/J+/bn9nd7F0j7809e7tOab9C
1YHIQ2S24Q4sL2jtQcj+li7qshMmtu0pIcm9/f/v+Zk3MIV+Ah0Aw6+itNfSaq38
vKnD7Swt32hFs8R+hlxiQfBHpKR2e7CSYd5RYJHW3nQqFEQbSKY0mfLCrIDl7ERw
vVfyjV73YIFQprv6dJJqZqiurGLwhan/Jr/TgdDDyvhSkNESfzc1DLnPSRv3I4bK
Ix7kpIva6+i1tYp72PDx/IvwO+lbB5g0z2mBXxjg+MB2L6uudNW8s8pMygoZVfhz
tPgQndLKJg62aIRl5cc1SE4agEBbwBQI3vSuZKM6j5q46kyYmFYCHADRVCMNx8Vy
bMRtVOmCKJ383C7XCTsM1we6cPB5WbcDHQnX5MEvlpQWY7yOJ9FF8IspsJ1ULPcL
Du3Vq/8DsHP+aFBhhi+2DzOhGV56dKaOp8vZW2RjzJp7Oi2cAsXGRTlY38l5GWcV
WdRuqrRZPchsA7bX3z4An683SESYF8MVWBSgKjyjH7bczWwJ46QuvGeNnVHLRzW4
0GyQeEQXsESiO/0NZD7jiCSKsHyunxbQk+AK/hKG6zVpmtEAN4UiRFM0Fr7KvQMV
5s+cOCZLyegrNAbPfcx68NS+jXSuk2mdL1dFCIGmHwP4Y0e57aKEtqeet13r9S6W
uRr8pC2tKaA7ntP8JnyINsUAgQ2aYKMKiJO3zs4rGZoekqYhIs48Jyd/VJ+NYoGY
/qlj8Z5fTzpwiWKIrAtybVCj74XPLUQQKxPVddy2C4KGZ5VJYyQSH5eC0MM8gJjp
oF/0tWt+lYHWxWLaCbHMEyw0RSxJ03QYt3lZlGwY8VFPbF0LoPMjJ1z63kvjO7tM
8VPWYwmMfalwwNngQ8ZyBmvtIRUE4BjIX0cZOi8vEAlRxPPxWtjC2bcyMK/a6MBR
w1+737TEEumMBdyRw5J5VRx53C+n53zToNQh31VboNpv2KSJaU2+Zjszj2KwJd8F
eGjxc3mxRYE8LBoX7AWQk/oHmg9k3A+5IS53pF+F+PjBHjCSW+Y1iUX0ahYlrAHC
a0yBJX9zUv/GqPzWMPfl6zxuA4e0v8E2wGu6hrvSxGoK4ZCdS3hMX3jUwNAT934L
WZxKRKiK3IMF16HgDZA3Pwop8PpIAXk8FleZq7auZHgpBiYRtCNs4A5amQI70czM
oCZHwpux4Ji1SkZBR/hPflDAhMReJHAWr0lB+RsfBkfgTeA1Pp0hOChbQA18Eb2i
YoUqYHTfpqNnkQplZWd3LKtDuHMSRC3+9salO6D57/Hq7EGJkgADa8u2LH3IFMom
v9qBMa/VFHB6MQb6V3JHTxQmQLCc7FTh4RnHvjRAmoUkvZMflgvX50PUOLccITTe
eU6bzhCBimkcEAC595zNTkv2ghAoMbZBRuo709dJuicbiI5zNFg0VogJFgIdjHiw
2aWzO9H/wV2pwO5amarItPUiJ3xkfr2XVToYBpKiQElIIBo8EFZzAnYBlAvhDjFz
2+/9o6kypRqrq1RNM+B3F5XJf69/XYWBQM+nbeLQ0ZdNDrr4jInkkoI7MIws2R9g
+ri4zocO90dXGc3giP0FP+dyeuBtrjs3a2YCBMs8SnQhpE4Nb9HzZITr1yergk7V
l5FNVVbect90Zh8PafP2Mb7KUji0XziO0IcE6+uVZucunfNiYvg+gEw25MKHrhWC
ySLfXB8UGbxdDf7oN7KQFnFg5WMt0E9lJOPtqMI2++txfmLK61dZFOwRgIbFmQf/
SNBAnjB1mPIrC0zuB8dzE8FvjpEsIgHvXsxJ6/p8ElH+BHHkaepY/+4edwoI9ZEG
8Ids+8kIIzaUrAbIcMcSBSYaoC7q2PQf2S4EhGF62gb4A04EXJT5zVec2V9AKqV3
lY/lpsU4k5U1h0R87F0+glc6PkYU+HXL5KB4vUo2UnxxtjJPOT7NVA2lOWYqzuFe
T0rRltPHO8pkEjkJD6V33HEn0bRMkE7+/CnYdRqMGEwFVTE43Sa6zJrcDHqfVlBF
idR7ZdcPuxCL9dq2futX77WFUoX+FiRholtL0r77yOs6pQ5/rlhTd7k7F2jCNCtF
gTU0DV//uYqDGn4uqwFhy2p4KEsUMrwywwz98ZQMyMEeHQFHizwn+RZDMcLFV2Og
ILrkq6osb95RuxrHLqDU1x7WfeoKdMky8obEmGrdzJDgdjLQij735aw6a7tAb/h2
OaA1HghLpYSpiGdusb9JWzh4zPNMh6ekrh7x9C41fznpVowypQRumJRMi+dYZW0l
xnYsL1S1ViVpA579zSd0aa12doqcis0dPc8XSPJGFEbmWDmnlGFDnWnDo2oJtBi2
uimAVvzYEdb47wMws/KT4+JsvAjNhO8Dp0ChC5jGJcRsrPFBJlRJa6u/uvUMlGlq
W6ZfP232f7O5kYoTFMRM3X5vGeLC+oLTRpWRuBKtzaZcQM4xOaXkbz9aw222dui6
GLHmd6ziESEmxVXkZ+Jqvzc/EYLMdpDProcJ14ZGkUT+IpBIRKdLlDIFPKNfqo05
xMyiS082AJFGE2hOmuktuWNoCeQ+WZXOMtTtlQML5cijjBhSM5r7R6PJ/GkXvzg2
HvXJPb9n1Z9UW50cAyfz3EqQ5XystqT3Vzb3LTwEspAPg6erkOJ8jnAOdd8c2R4D
mlbKEMMSXr1SfIxD+Ne9ZMpkXnUim1oN5VoWGphaxm4mW+WGd1K67NcwYobVZK1M
AqgB71JMSBZem3N+1FQS/YkRtXTbeVl9wruRHy5VCRng0q1yUuT1eIKVAoCmSwL1
b4d8eskXeDQF5mVhL4v3xVv3IrLQYgsW4X6a7/mC9it5mSKdVC4X6uAVr09QCRiP
fi70iVH8p1jVolh+61EV701EhAoZvNmg+V6xmmp+fe6yuItjMMZWnMmHl+t3Vla6
A2NRpCpu3cA040vJFpI5ryCgLWOMnIzojY1e8p/iCTX/2T3dPS0zr7O5uXWr/Zj6
sR/HdVMqp/782hT3B/Gx71KkNElgzZodvbBy/jVsQtn8881nRSEkngvh9qqFepyA
qskprK/5w+uU0l3Ij2keVCj3sQQceGJLPksyARqVVuJago1RZOmF9HMyladEHmOM
6jnOIjE3mYhgPAVYD9qJp0X24SYtdpQOr9RpJGsSbhrfDQvNA+9uAu1TJo6qtfKc
xVTGcTxU7DZ9jchRHYWEDDyh9aH3kxse1QTx8/1Szyen7b4N/jn+b0RiV8XsjweF
zbbeG5+SAQDRRMcQOWGK3Tlv2r/XFqRqczgSfEasdqSkJH8eL9XpjU+lfMVzgaZZ
fW+zfQFVmId+rD0HjKyydHuu0GG7RgD3aJw4sLJH2A6VrXbIn9gQ/XyBVNX2QusJ
qnztuCsSbxPSlJcRRmJLldXEzfuKwUTy8fwbtIs9b+BSjqVySt+yy2qRgMFh1woY
Jl7AIXYIT86LX7IwCqZBawQ+TBP1iswNbyuIWipbVgxw7paiG+DRwo9C+t3Y948N
t5MV5w/5utpm1Q3DfLHIE5fn7yZ781YTasp77gJwyskj/wQI2ai7A7wKJaXqX8uu
EoYtsXNREvIVni/FLeLQ402aF4Dn5wAbB3WJGtlE1DepDDp+28ZhGkI0Slru9KVx
W4R14nSwj3H0MiNZbBydCN95xoqJi3GxOMH9G4IgsYe4LIxDHWQjtFpzjTCQh+D/
xeFfZJIW4zFgrbG1mb2sUws5qsuVy/bWPe7T3HiA4a98g58yAUjhszzzKa2LpIxX
`protect end_protected