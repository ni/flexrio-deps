`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1456 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
5UzYaoC3tfpGCmdkAmjlgvbgx7ldpdu/xE7h2iwxJJe1JaQ3KHm22vayP2HnRzqZ
2Dp8ANiv91X6TI+RrCPOBSqrAT6/VwVrsrQT8Gf/ntVdybi2h/Z1VpxHBZ9pY/l5
0/+0sn8JOUM2UT/8UnVwr81KUt8p3WE9F5V39idz7DyP5cE3dfEdMl1g8ou8Lawm
WGcUUpT268iMuvObuoGVt4nf/gMACWETZoOjpMYz32KGpteklXiqIMWvP19oIxbu
VeoNxN+492HEKE7ddSEPw6/C9l+8d9FWfMiXI9kAvOrrpncGdQMGdvpT6qyGD5Z+
UdoCcOuvtrKabggr6JGx1Mc2rDZR+H7XMVhpqKvnyr/9/PbSpU3s0hS3QFMVz5ZE
IIK0hW1wjKJBQd1LJhQ8sgKFM2vOf7yjbF8LoCAAzuWKiFVs8UztR7jwGwv7mymz
u9T5UxJxvTcNDvUteD3AXthv1id8x4L5Og63Zl+bz4C/0UitwaiE54opylJwgZKQ
5SeDgb3K1GojOKFsEiQLLy3ewfhFniZw/THRiL57gcO2/JB4qOWaIP5Ra9ZBJwP9
Pfht52yJMGWs1jzNiwzaUU5YPsXlqNtGU1LFElJEk0B/Hp+hTAxA7FRJdS22TtUp
2JvPh/tj+aMAgdFNGP6Jyo8fnGvRWHM6EsHcrbqTVFrkolwEfkn5FX6vSiAHL/LD
Z5G5SttH6MWcHsnfJ/u93lgWKMt9qKmgFmVt17zlTIPF8jx3zoQXMQyWAz3gAnOy
qiZbh76eJaB7S4aJWhpcMKtLOOHZTC/0ZY4UQeDjvMjxQhxzbrWHI/TIn8YdvWH1
yaBqkATjvrr6lqrWds6t9qz5yluIjUQng7iRclaNM/7+JM2w7M4oWiICp992MjiQ
iu+3n7mT9L+tP7TXnCMIzYbt7s1RW3pftF6kcwf4ZYFlUpFDGOo+FM+TxPog5geI
PG5Hu1VUN6LGg/UATvb6yZm0wrVaFoWVPI9LEwa9KWwZyScmpuL0gEjLI3H4Xyck
9meE2h02f/af8obIEWtt2+HSKpSPdS9jasx4CO/Vki+VEKRrp5Dxg5EI41R6ePzM
/JIO0sBDShJ3gSzgdzPQ40HbAZT6oUk/KdyVw8a5LfvJ/nm6TpLjik5v1XMzcyBt
sIJ6ZAp5ZD63MnU2sS0O8s3O2Y0j5/4MGY5FieAxJQ9Wh08hnZshcIn9XeHBSOD7
3/oHkMF2npRa16Sx3g+NrDkp+MyteET6nZKUXc+rbgRUj2pM+q2EfcpbFPwba0zZ
9q5Sp49Efrjp0DmSDPyvwERSZYepDviV1IU8ThPirxpex6gWCS0k/6XPhA/JsoYT
ewBM6GhgFsperXURD3BgDODo61z+riyOj3KaVI3IU0HEr7qGZcY19C20GrsYlOAs
Wu8i1bsctFlewqs2tHd2XPMAtF+dpxJ65X++ElxLKpEFinrk4y2uDk/MMd/4AywK
j/UCoP+s0PovyzmCreDJAxGD93t/G0tVGLJve+wyOW5YTVr9ZLA1A13CSdIrhxMa
YlAoov3kjg8l1gL0NyXeShaD3n10XsELYzijz/sNvIA6Q1WPYnGVx96jnqh1RTy/
ejEwdv0uF7v818GYxYFlKV277Y0+Ut4jBPp1feIJHPnxE/nHAoU3ufaRRxgznEmO
+EMS/CirdQfzmjG4PhR50+MXskIEEoMQi1A4wt0HQIX+StPFOHagr6J3zx3HTE8+
LYKkzrtQGrEVJZ1Es7Tt0lJJooUqCisKopNlB5PXBcpeDgih+/o2pRvztbBwDv1D
VBZ+TyMr1hAvCFsPGCUMwQ==
`protect end_protected