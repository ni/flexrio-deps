<<<<<<< HEAD:flexrio_deps/PkgCommunicationInterface.vhd
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6288 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
qe1+t0GXQ5YjcbQQEHGgOUjJ4yn6PrA0G4Zj+j6ZraBISgjBsmapZP8DH7wcZcH+
4smSWGbj82KWDaOJePTiS1V0sqnd2uHbJqAjAjdWyekrr9LczR8cuEsanAPh+u5R
cDEGs7fK+5y7cD+guSo/iA/lo9W/cGpyaBrIhIKgvJH2+67Fyl3tmVyEXzsz1HVz
CqHynWKcfA9p+7PTnYQ5UjtRj99mh6awje84HNwWUeiKzfhDcVPVD+3N5Szpr9GY
ZWxbe8OJhlAYnoQ63EHf535BuA/YTRzM9nDgym5hXdQAfrXi9veQm3UeYQDVBk/G
SmYYsxawy5ub6GKNxnt+ChuzhBeSKthKt4p1lGp95QW++KtA3+SjgtylQuY4Nb+j
pv17VXsCRqddY+aRa1/BIuJyIPg9em4P5Y8J+0X+fcxh4pO2louAS3eUgHEnFkGp
A1EpXYTHyAAIdvc9hyuxpmjLUi75mHMX0xUj0oln/PEmSx2i/tNxdc8W7E9U5PcA
V/azlwcB59lPHGkL0hVA1AFNetuaDv1oDfK0JqxMCWqyhS+PlRS/FWwFd6YGIx2X
h5qInp/rHb+LnJTRR/A1ikbo/or93oUUnmIgqNVYSAa2OAUSrKwapSCtPZcYdPUL
O4IA/LkmVp80rDZTAjfJlTB41rBsWWKZfBvFeedV6M+/rG0oYR+RHTjj5ND/slMR
+YNTPkujGeyxDc0BETxhru2j6DXy8Xd3Yi8KN2WZkyhQCba5dy0IqB/scwbsrjK6
7sk8a8wm2m3FzjjSlMtjsu+q/4bOdAI5WnwdKc9r1dwRqczmfQZvf8bC1VOQBEhl
vi//rIlkA16QPXwcFm1JIVlOyT2zmRb6Z+3hvpfkFM+4CcAfsy9NvqvGGm0maFNW
+ei6fJd7f/nwIs+PCCa0K78VVcXwSTL3p2mSVSJiKOH9m5UUWGHsxfvEx0MWYYn0
v5xAvjJXcbt1nf2Ys2nklG1W26HlhSxL4zoIfo4TgCgXlWu0tGnP7vZCIf6PZQ7C
r7ToM2D9Sc/d56HqVWt5RamBGg42bmhwOEp1e1PZ7z9RfxDeN3gj2Q1uKfH5KHKU
BjkBFTfmoPwgCI8FTvw4eRBd82xiEHS0RdzgmMYBd2ordOe9UQ2izb10put1qTzS
R3SP+8hIfdov/iEPmHDiSkZATMVzgvTVDjazYXaeIwB+H/Y4XLk8xVEj/lLGQdUB
xtA+eG8oJqyTamdQKXaB/vGmNt1NZOSPUAK4OI4jwgeSsrszgNz/QMXusLfY91X0
r11BtNfHEDuIcyZa4xS520GLnVHvQjZTYz8s/ZAueszo7fVhqUyZw9rjwPy3+PT5
peTIPDKBsRM4Ml6lL4xYRVV20Rs+gOtkyJmmSNLI3vzJC/Ydowr/Nqk5JcFYb4Ia
4WzZzrXvmW29LOyNSfTnwYpqGge1xWr0RZOL1CjizyvcbaBwvk9XrrNEZwVjvCjU
zo0tV7q1Hc082Ly7dDE/qYAo7Q0dYILgh9WyBnKXnvBpTQ5zw+ORXbL93ffzf/zh
GqNaOAZRD2ctWFaFO4KrJHKii9W/pNPxaatueiUp6jCMHhaepCSgkPBVbi/faAEF
ZO6z3EEvq/O65GH21CsrEM46IwwSDOA6CK59iDdU0XRZ8sUA0RhmKLjAxe6I2PVY
JMZ7x1tc8orKXKeWdC/4LLtnkbmv5tf3IylO+aKJpBlZgfOQSSf+DyqyqzhittcO
dBxSL+nooGu+M2n+4zSk6ZY/s7Ey+dMBlIQoSUPvwt3chAqaqfPAcJsGRodzDoXX
AlgvOm5hQH1MqjmXtsa2R7XPEx7qFBeMZiDWCpG/f15wPFtqE9Ke2Tk4527R4mm/
9G7YMxTXfNRAYes/j1nWUnsAxn+jHtyvdGRYJm/gVNNN/lat02UaqFQjOHek4A4G
qhPTliwslJl1663Y4wU03Sw2iHaI8OLaHk7OqKy1DxFnWaQSbcl3s2Emn8B20Fbg
Sq5fc/CpFXBDPomD5jD/h0ePaP93Yxya9cKwlBUusynq7MBv0tggwjLEbux1AT85
bUkZKpcGhHofG2HRW42hFAiahuhuBkjuheXFQfcInvDr4ldAFz6ZjnZfp5T+fhre
BXrWgK8udVSeGRqW+CDKr/cERxhbBm89Pg5tQWdO/Y81K4ERg61UjXXneUj1GzYo
I8fdmHIpxT6y6sLrEMbPmEuz3YskNZQKPdOAXS1x9a2xHhN0bseGan0UmknhdZH0
pLYGGmUc8Yfs5rHNRFuY71ISAgHa9PJaTvusPJo9ocGPU0DfeNz0C2NgfA7Qt2zB
D13ZGVYigq88mEP4x5421yI9IYVF/sHt2fCSQLNvsECMIVjbn+tqYn1lLaBip0aD
OICoyowUw+QXOeOAFACW01gRWW5nCcAwcmCso7PqBV6Gj9te7J8p2WNImeoxzv86
1vyftEYdPLKudarm7DpRu2ykDFzkeEkPvsiJTxkQCmYBWhEr0CwISmXjxn/p74Ds
5Zu4qg+ubEajjg+ahcBaSirxR3+0G1hAhZZgz10oJu9caITJGlYa+GxpPIP+9lEI
T4y8t/Y4VtXtApq6Vwa9ohoeLbLA1UsphtEQ99BOXaaAy57d6IAH/Wpq0S257Z5a
R/1aoD/BFzyluiYpqwgJiCpCpQDnyKo5qvVV+k2QAM+nCmpq6+oKFf2D5yI7gXYI
Fbh7h16usl2RHMdZtBeS/Uqz8Ppbou1Jueg8re0qI9biaTWeFA3juJI43gbGjwTJ
9OwuhCZO84BAZqn0N31LxNKVXOHS+tA6u7zRY1Pah5dZQFrcWsd8FeoXfPHNIj9a
Vyqos6mLSrafYyJjyTtVByXYT8dpJ/y9NZ6EWmjMHitx9r1Rfy9d3ZtKY7uQ+Vg/
QUMFqcaZP8ZUKV4YYuaRZuwhhBV+9KaanlGwuLpNtWr9MUG/TzaTNZO6FvBlnVxH
qmtOWTtmv8uZCsrOtqrtbn9RxfnARBLQLqqrIn9FDBf3Spuy+3e9doZTg9QBRacA
rTc2hmePWStcYLiJyaMbt7YGG+PCDGimi41bda3mBbWbjnTxF3S8BvQuTWN9RpxT
lahIdqwbObhtKzTOSmGh4bJ4lZ6bMyG7JMemlh4ITRcGvuqeAvl7BK/f6jNbDZ0+
61G2HZlVO3CL75FDXnTpzC1otxdprD5cIrBEU+c4XTtQDQ++lPWhSUJIJ6OU10Gt
czQNmcE9WPgb4vT3U+D8BUlY8d/x2HhsSz5oSkSFwa32Vy0AHgmphe9IauM6NPS6
z4MXh8ZjxMjlWJcURfv6IewLjVc1mzJrkCFvF8v/tIAnnv1FMBRmrFkwpygqAy9u
HYwFUUokdwJcc+nq6DSLIeItt4qjfk8oMuJBjnukj+OldfEoeqpeLNoI22TjrKlT
sj3z1n6IlaUr2gYghdPfVgJzv72tXsUPENDeN0xMOvXFjvZEpUxuHUTbUdD4N0uo
zLBTNlxvOCmzHaLsxt0b10xa5ju1q8cArPuvrtVm6F652SQEokT+yOjzPLjBGotC
ixS1qiJwMcn36foJhn6CmrRasmPcbOowVGIZta2edJdmea2HgnA2Yi6vvzuhWVpd
7OC0wknlX7R3sBw033RvK1CiQFmIOAVLshp9o2nlTQAAnrfng+l4wwtvNGowyuhz
jGMvKm1w0Gn6hHy3/l5xj2pv0ZW4M7T87l4WZd5WHqMjYZQ21o1FFJrNjJ0E1wyf
U3/BZYPswrmXFqTplJFCrsIKTbthWCkhHKlXeA26nnVtPsWb10n+sIOEbIhWJsd0
fK8quri5eQk3YrBdj9stbWDd+2sj7W54fkPKoSIEje1ALT3CBO3Z4TIivxO9rzQE
+EBLVNSFcB7M1IElIMbWq2tVe5hwg5m8KlFKkSaG2KrflBE+eTVfTdU76/IqLbHW
YW4AsI8gWCh9zGq0RRZ87KiIN4IeuNz+FG7eXSLsz6lxq44MleVu+LVZrSAEtrA7
o4mKTI7yKn7I+y1uki5XaS7SiPJE/THSaHAprqUFruuLFB2mEr20ghJ4zgrJtyhy
nUpTKrWDOticP28nfRoI2tYe/OXjXOLuIpqdTKkAzGtYJzes+MU0wn2HiaAH1GQ1
MqFNqCBcs74NGExKoWlSTjMjTH/lDt6xroGogBD2asI6X7Ps913OMhcXMNhs2Ijo
/+mZWh+igXYcA381FFKF5qfGVPGOxfkK2s3eJTVqCHg58b5UVCw2ZJSl1zuhK+Ds
mtlT6cbNNcOQI8wljj94OnLfsLkU2nZN+A4bBH4KURwbVPUQ+tgMd11oYHNxoAFF
rXQYPjo4d4mUmGFWyU/YgsZz9mfYS/qctJ5yCg/RmTDZHSoBS7Q4jiLCDeBVojNl
cksduzhbaDPp4HDa/B4r6yW2x/uy2RXioAVxMuY+w5kBwhFk0HX+dnwN7k3BmHbI
LVZuGXAgRbQLakkzbTRLl080EjxSx7sBPigI0RLWlZpC0caKiXg36fe/ScvEfx6N
MerHjBXDx1V1nN7RPNyGRLLi2me0YNJywXpDAPw3/ClLlKLOT4++JVOpF/pEgaxG
mvCFzFxBMX58I8Kl66MIe07dly8Wivjht4fl2deU8M9SO0IqYZ7u30ut8vq3PnRs
CvRC8NtnbrlIXqS0acc627v48/v19CkFxEGSkAFcMEb2Cir/3pbJKO9wXbEVVjaL
VaZ+hi6Q3kHiTFFbNqxT6947QXZvRkqoGC/zPPe3Nd8T3i/+bshCCR/MgCBNm7u0
J7foQJf1YjViV20i4ohDUJcDDVtnno7YakwPzXo9d1Muu85+W3uOmNsZDhj0vpKz
AaaS4yfF3C1eKdvvFnbMNbJucwrKbPdn8kcG+pDHnGspMgeR96nIAgqi15J1l/Cv
jzCj5wJ4HgcHFHx/y8VPo+Yci/rBrHBDAfcWxsAvwhI3UJyOqEGxrft0+duOw2dX
3gsVbYkGzSFp0Kb43yx8k32HshT8k6elEwH2xF25VCCSM1aunrA6wkd4Yo/Ij4GR
bfBaYhb/maUBbAgZO3TIPWOTEIdU8jfoXymtiZUiKkTXm6w5rTIx1UacOcMbqoa4
51G7lbnxzFhT90a0DyEs5ILD9tVH4bvGq25969WUrIQ2EzagwLnV9MVMueERuvHe
diXiVK5x76RFo/I4OHc4yxqoBE1ZkA5WwF4VfPQrPOdb+Ko/90m+72cFF82xf0Th
m4DNTzFx+iYfetCR3YTOPW0MpYvWFeZQWbiQFmI51drzK8fwcq32duQT+d1vuL4S
rSVXVTYn70oH+zzjIgkqnP1S6sK9eEWCcjpQLB1Z/KrfkpDeXLYBwCERWyouA1oy
uTP9eJYaapl9Fj4w+T/W9fa/fDWRurT0OqZngKgOU0h1/70pTV/O/YfkJeHLAIxC
9aP80QydNNpnww9g4P0g4OYGe7+WgjdvHIh1BxliHkHAxjjG6fNywdVq54sEy7Le
BN6BlWtxdgpFeMwW+cJO1C3Gdex3EZpTiXbcB2mgx9lCptKU39uNnjPOHLGvwpeJ
h/Xd4KJquoHcoDhl0vhZ0BJvFz9bQV772Rl5k7Xl7os6XlC2pdOGDCUV80r7Edo+
EJSuf/AwZiioLWD7+rtNB3wXUZ8ty+b8/eUz3BAU20dQ+ZB7aay/TFM2TOPy7Y09
Ua5RnznmMj6dh4W1r4xXiL8bo27MQNM+RxhDzMcOMUhOFDlp8rzJeUVCbbRjTZRK
cdjg9aXWvhRM/MIas0VEV6eFddBIDtRT7qbeCMK7iwZ7pw9FObq1B17jGEdPpGac
qy3JFsMhOHT9s3DG1snm5eXEuZCMpcqkyPqyhU/3D47ytP7k1eIYNvf+WQnx729n
jZbu6KQKp+Idt3FElAnrkVmsO5NohTdiuMs22+YmsvLHjMZQGyzHO5p60ic2BCl8
JCEkOm9q2BpqLyKCsYGIu1NzLZxK080LKZqPfI4aD/oVW+6ADOb/oQflBxMGvJZV
S1+Yj4rUR7msGa+wx6sJmyfav2RmKQ6fmcW2Cg6i7NWpmLCfh/S0xPYy/Oy977Uy
vq5XjFncpCUmH0iUpAzrUCdeHRowSLFXXTMik8ywNLqeI/ITBCzxYLqZn0A2l87l
X/cTTP1wGxHhacCW1Um2wIRWeyvP5KhuVpJTP3MV5d55/8wsruJ9/l+SWzH7yRCl
CgUN4A1CjNzz2WYKvumJTq2OSDys0v0qLrTwFgSZgzOxdZMU7wS2KVP6tY/eP6Xo
tXBGoMdRUD61/oD1FP9yZr6WOZ7LR1K+1L+gHl/6LcSmSuHEI66lRjV4gRkimV0S
RzkT/T/lrP3DsqNzZVxo+y9UH9sPBkuMcI1gyI1YHtbpxr/hC7jP0cvZdyYgR7Yr
Ba4rN5sIOsnbTsAwgGgzIadL7CbhnqqgC7tzuc+H0qDDqraWZ+Mdj+pIglEOAhC7
oFPZ9hffI6s/9Opl2cfSj6Fun4Ux4XOgZ1hShMP1XucOkcGqZ1KdOhXKUmsHgxdn
HjNPtouvgfv3B5WOdziKhcy24QkzO5mlRuoQs9yDaYFiFZRhe0HpauC8NU2qAysg
GYMO4qLCrm6CYj4PJAloJoPfUY3kUlWFTi0gKUQI/Y8kHOVL0KOFNb/MtFNAqMWS
qBNx4bFTZEcPZXMfU2c3z+zzMGs3urmJ8ciat8b2vT9Wr07mAs5h+C3BowG1IZ5z
7/M+lRXBRzY32rXx75dVODM02/eeJY5UG5FpW7sg1i9lB1Pdxl22a7ELoO0pC4s6
6opjWWgST39GwmLXqRRV936+DZwbiutG3UwjvmvOBt5yvBGdfNcj8jpIXf7asfUd
mDdeAYXr9GQC9yA1KcHJu3kuU8k8DUDM0Wtwui1OOKZiCAvFwarMqFysJQ4G8rg1
ATyLA7Ia6yjnZEBTnMQ1d1xz+1TCQB4HqdqtmZsriJ3wEPDpGD4DfML1x+0YxxuV
rFaEnGCDRBVAycB4McYga/uApUEvpxhkFfktl3hRWNjknBda0dJbrnF93iVP/HED
jgG7D0YgKbxqmy7OEtE1wBXZAmjfpQ5w+SofuDY+Md7WoHbu5+T6czTQg57s/ZdX
v+IodTJPkEtLiC/x3p8KmJ4DWa0r+Hl6NDgjalBi0QCifoTZtVV7BVG8SA7ATauG
n9S+VR9PaA2LTZqRW8eMmYKfEdKXYeaB5AAvte1yxC8kfOFMNmPTxzbPFc82PWct
AyVhG0nX9YmjN4GMJCdDWCxWT6k1W8umFG3OBGdNH6kw8e7yqAyfCAjycFybx/ww
lCqsB9YlRuZUFlyJoUVKE2h5vnXHJVX3nVCWAEr3VCgUQorz9ARnpHNggIGO+L+D
9XmAxS85CKcKk6ozxrE4FsLnS9A6GMYwiu7gwM70E2GNCUBVPLI4V7ZiKR22PZZ3
OEINcY3hGwfBxwh2atQQcQjAqBoHC4EQPVU10PPN/1t/EPHLbE2UEUCgSiSOXNWu
HTi7k0jE3ujfjdh4Q7dLxcotxilmqwz3d4LlV70YqrtXWxeKlhXQxr2Bd71eFecp
gx69wYhbuuSdRctJ72meJKmEFXh/DSOcLhJWenfOoplYRuk0c65wPYEKqH9RWk2w
BalAiGGzVmsia5JvX7MpHbqQ4/2o9hk9GgAvGXC3LVFXyPl56MiQmsCqYeWKhWiD
vwBRkuou1dO1yk+5V1ILNNkKExvnJpPGyUEXdBDi3XLAwFzGV45TWiJ3A0fmBKbH
JA9dHyIkn6YuFIZI7sboN0Lc8q1JWpsGJXko/bU80vpDudFCefPohuC7d8TJFWGJ
h2aAhpuKXZJYDt51q5fWcAO+4dwkGwsrewCf2jhMbtdm1ZCwPbwBMC53tHm7yEh+
prhXV9PsHhwKSsqnwjzE32DRKEgxIiB4mB6vKBIBKN8VkaE4Ni1in6aEBz7oZbD+
EZJC+S9m1xAsLATFS5fTYFdH9tsQYjn6frnXePZDW23NUihshUsC1u9geMXYyr/3
3ODwolrmb088QbOcxpENApX9/lOqwRcvkaDCiRzuq4LcEwa2t9HWl7buzX0izFha
IFWDs8UTVQQX33x2agmRcPCZj7Wj7KRc66YR0rKRGecjH6mXDvbPv/FlS/LmU87y
33vu4Ma8JgjuGwQqNvwDbwoB4L64NK/PiZdMARnbQNu+2kF6GMh8p7FcjmlgNkpO
GwAMMj+lCBhm89TsgwFo905Bsy/JqfM26JweAXhUQ0mleJH0Mo5jwnK5OAT0NPhJ
fnExyrm3U34qNLaJ5ZNn575v+4nTSbjPtuU0xI6BKQBWQsphv3PJteZHMrtJDhTP
=======
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6288 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
7d1aayJWrMXzpB8QUg69LBipqobNIYgvsaCwrGg/RkhzO4ZBKwEcPzRZniATJ7SE
/N3/4J4+NXiUSVql0O/7K8ws6gm296GGhRm3v24jkPEnLTeyvjpDNHLOMQDo3zwi
dcN0N3zSd1YkNoyqSkstWY49kDmu2IgQAe+hk2oQ1u8X6dEdYc0u3XRQtbJ3No0j
QRD20B7PssF5ABGKEVceZTgfqErAvDWo8789GboyObb1Dd8hQb6pJzORqRiiHT4E
dVTX5yiOhk6uZjUXGXaSy5qtMERa8ZvePReuzZiCLBilQo83iCOvf5AI6vRXqAyO
rYou/Y7yWD2Xr9CqCDso13sIx9vFMwKR4bSDfEu8NYj4fjo/1eFNsmZBpzAJ3sWC
03Ni3JJ2KXp9+wx8UlW5FI7Fozbc12LUXdkDgkFvo7Jt7AUgcIGicTMyv0cSieXu
NP62R2i6m2y9ZdiswqvUJQof6xaXhUTxsPreJGjtDRoU2dbLWqx2wKop94Q2IucH
jqrumD2YwH+yx0GfyqXM+7W1ZEs535Fy5kWZnyEXpU8KcHP8EahBRP50MhkW+pQy
pslnIn796SVcsPZ1BkyFzaqaZW2euiGp5wWyfebCkIYegQrkuWndXYlkE+0VLo1o
PHk+b87RRbJ8QPa//qpKznrncIBUosakkslsl0UbG2/rmAX3EWXG1r4D3IC05QrH
mrRXp2G7hj1Yy8O6KhaMc0SY+xjqBiZnA7Jkfh7OGolai2bkzwTP33Jl4nR46MWd
xO+YHIWPwN2aijWqk4GedRCUl18YUuoJloXteLJ9zlhW9BpSMPxVXbCR2gMlgt5h
Sh8f3WMJr8FMOZ7C6R58sD3K4zSa0i8XVm4c/oQVKjwdSQ6ekd9fUEIqIS+7+sEs
WMuJnSUwSzH/VpcSSAaZ6DT13ALe2VX9l3WoDNmu/6QVFxmlpaW6R5aexyp3OYoh
7vdg/FtN5+025IvVuE4Htq7sjkGWRAbT52Ceh9nF1lsJsz1aD6vdeSZywdqNaEi4
g8vv/wiZjNaL3+07pgRhgT6c2BNFQ0oJNTPp9I5oHwyihsMjGKEUgDP5pSiUDjeW
FWLeh+dcVSDye0tS0NMmFpRTryFbdMkJNZR89Hycw+D3O1XbaKv3GuZHClOhW/Lc
Di9NHYDilx9Mv0lFm94BrJVpcZLE59ZUtM7t+dLxNkkOElAExTS2azlcwnGqWi8E
xWvpMyBHezJ4NpkTysTycikes5OozytgffptzrebBCmXBeVCWtmUe4mMCTZM+UJI
4qeewxrtOiRDzk2Bhj97KdjLhe1nLg4YbIabvyyBDmxjj1BZSkPRz6vAiZGtXyFb
lGekZpfsMNGJ+d9645slQUmPEVn/ZNt8+WgZ/1+o5yHO9/wtBRfOzb3X+ubX0n9c
yxv6hOiw9xTQm+M8QeE3/lmkclgY5Fo/G9++A2t2a1AKbdjjpQWslT9PjYKCHwbN
dj6YKgyg/aR3n4JzJyYCmxqypuTFsDtG6n5kubel/8+E+/uk3VsxFYRHTqGwGsdK
T8kdsl8wpYxXkNONzj4Ov73+WeeMWcKn4f2oJH9KV3sxot5Xjy6eTf9c0TbN7cHW
hcJlBY9o0U9kjirTh59h5QspKIub3Y7OTLok//YpfMOr248Yk5QWX6Gcqgkirlal
TQsmZJNhv9eMEzHuFuJdWbMlXBtC9Rli2SSFKQVKCrRtG0LhOnahSQ2p3QoFiKxK
A9U23Anea2NnKezOD7x5H/P+sCnLJKVzgZuVsTZx3/V2wrg8zrn0PaabtukMS35+
Bfh88bdtah7th0JpExGHaaF3PNUGRRXb3YEHOsgqiHv5Yn29QJfxJRARej6fp0WI
XwfokVB8VxBRx0GiSlqp+gcSTtiNxrObqEuopnWy3GnjG13vLKycmDOeLzZrSsGF
PhKZP/Fzu3xWtP0TFqijIPNLcf6WgUdHVTPS1GktFYp0eqjcB0dmUcm1CHE2fbx+
exZlxCmx9lECXiRlGRHaeHIYpzWxhiTn5eXagkxnU7EMhql4Fuq1XRGXQG/v8ntI
IHehKO2GTI0Fbu6Lu93Gf8V8JNNoTTlrmYkCwVcgmbQNz46n62CCCFSlIGElg5ow
XeS2ngrQCeJnW4gV5LX51y/fjGncwg0db3be2vXUvdZhszQ4jK+LZP+ed/tA8u1a
8NaFksF4xIa46BbmPuldtMR2TLcpo2nKvEOns5oitrC7sw6SZMeUJJoetSZHSJNq
XzVM2RK1ed1FZyWq6v6Ted/WgdwisHF6s9y0gR+hmwRy+Ud+/AEM+m6qeCgfBKmV
/JmHLzhk0+wXeWm6Jx7vNxYb25zglliyTskwZ0x+/bl6JJJj0aHt6Mo0gFObylJu
flSYYh50NXZusMJxc0xKwIs7pSz2kd8232tzWwplsUGXdazO8ogZaLuZO8U0gXNk
XI+AOgTZ2EBiFiAi7KCoCsXuUUR1B3OoAD9gEfq+Ng5YzVHtpWR3ofvrMxpdWq/C
w6r5HY0OQTFsNXKnyEjgNQH7opMHTjUiCwdKnaIc3Mv9O3UA7whkPROleVghWTpU
Xp0Edm0iNV/IrrMj0YLmJIXkDCKcApfv1IP7W42GwA2qrM0thAEmc4HBfe0RmJb3
3JVk46sZgM63pmDY/YKT4MziVdKAj7DzzETreDedjoA2zdWaA/0nhcsn+IJj1tMP
RscQ1JeeiMGay6mfZzcqGckw9SB66EPYRz4Oo69WDfTGgR5wHkHnxdon0jP9sdr6
IQy+nEycMKOQHS+he5nBvroPJythThsl0nQHDLb4cc+7Byw7NiWPqzH0W6aGiCVJ
lYHp8t0qGCNJq/pKfqrJTBY7tJnHQSuKuUJVgq0tAQXDMtPfVoKE4nWjwF4xI2rm
n4AX0ZPZQkm9/nV6t3KvEeESg+7qopcNpvzytZWdcidMmClminLaTM1zUPRB536g
d1wKwBZNqgtq/sLAVAAAdcjKvMSrS/ZrneljrAxJtc9pMF+erTZ4640qm4EpoMm0
7VIyrMlJfqyL7j/sKbHphJ5QdiKHRSHvnGwWmKjvqqh3V41NSft4UoYlDkRdCn95
3YCXKsqf2iCicn8e72dg4y3btJRMuY4pnly/FKbeD72kCDPqg29e52FdgmmR4lV9
01dukeSvS1woEoFUj18sw4HcM5Ay198dpY+2+scN4DRxCuKrQariQ8PLqF9BwsrA
+cPdJv+0O0fwlekdSTraJ01JGERO1q3v9X/72OgALqGgMrkczL0eDQ6O81stVF6+
okN8Pba31vf1/dpp9TZsoqJvJNxdFtOtzyjuTgVrDDU+QzzTln6XroPe5slsXIEw
QIKnZPLdJgwOwuNeOicOlghBiSd+MLMaiIhET7c/7lSH/zPIAgEAx6FMKrrsHPGl
O90QI997r14ycyFdr7viVNucr7xM048KamQscbQfahhaun47Fcki5Ey8+PvHjolH
un59UhvsTeT6gxlqWJVlCS51tSANbfv5InfSuygwR7hwloNW5lBKx3nN1KokrBr2
sk9POts3+aWnEbzK/J2QEOwhLi6IwMRVCyVd5BwJLKc56XDcJ02QDefup4QrQn+4
OLIDOOtJ7XLnwYFMgaaRYm6CZkuv6rMG8XPt+xBGVIYURSShD4u2MYg0xY5tWdlh
WG0J8mVbmsSMgjVCe3hUZX89mDHNRhjmOuLukdviXyT14kRkBnEqL8KleHnz4Sl2
jeQiTMLSX/mgH5Xyk9Yh62mfB+M+cwKtruTN1oJujXEDPZPWHp+VkQx9k6ntgprZ
ShrjsPqYN+orCu0MqByxky63bGdQuUUuRx9CSn8bJI/SvvuAWQ7lOQt8qVrR+yu2
jniG48TPPz2gJcgq5vwV+Lm5EylBYyyfSL74FPMlUOJ32jIlICgQQgwIpsrPmJOd
fKDCDOCjX1WOAl8dUNjnaLi5r+OlI6tyK4IijAiMt+B9ZqBtBYakRBJ5qrvgia6e
l7x57fgNrdvDwH/jLScCenRekFb4hH37US/0sOqzzpTEUn8P+adjebds7CybKY9e
UHXDaSU7kWWHKaZWAVP3sHdNkmcfoqsHYCXo/BtjxiyDcH67UUx3qiwrk9kXKxt5
tSn2nCEIuBubTAec3PaAQL0ndLwrqglj5YVAgnOfxmLXVwQynfAt/T5MJSBVHwOG
keK7ITmmNiIHqTWSlnE88U8DGKeqTIPgeOY76CkPjZo0bZUacLXPJYLfuf5PJ4W7
8KearEnENffRpMWlAaLWXWc4Eb4T0tLliw+M0FDq+Z9KMnI3AUmIxGN4k61NjxOo
QbNQFDcHVHJXoguWoKaqfI1kYw8GbMLMZgo9wadkQmqHw1ZScrcfwprVfo6KDOlX
V35rA5Awi94eAFOYTkiegFSZMSQg4OOeHcGSSEDZhqIj86s8U+oHlr2muAvEnFM1
L5FfTvNVb464jlvh2ZVqd2W98hoGzeFIxRujxAQjn7VvYOb1fZjlx5yiGtojX1pK
tcSsgtYPVWtcwXzTM952iAivTDYfC9oKGFbQmqzeNkcqPZgoJsjFQuD3X7aLlYZ9
5oUe0FI4WEoHnFPkLMmVPcvggEslr5vmEpmhTHXFEDzeIofdCeBX4nw+lHNk902U
T/y8p6eOVCUZm4Kct9YYYU1Jx4bD76HXtEZxuy/9m5qLHn2U78HkH/2/ZV93NQEm
z8lxShE/x1i4O4iQSureVz6dW6LYphJU0fMmGJZfA7S5jhX02Aa7SFkejynm/3aZ
6uSF8XvwPSRjFaYzORX4w40HXLvPM3guVqIf23AQNk0tbdu++xs4M7FTrdGiqYWx
3uo/jT51YrUQU5mWZWh0ohYlYWSFMQ9aa5TcMHoi31poCSE0LS7+7MZ/DMyDHLsX
rxHxwOVbZI6bLDO6SdeuQLF06jILJzDIS5hhhHnc+3qe7EBDIx8pxLpB0DXNg/Uh
fs4Lsagd4TPxVWv+QUCYULO11NeuDZbW5P+A/WiOrkV/oSAd52Hz4GZ9hs79pidm
sAzCKO2JWF85CvBlL7IieiQEBqtp2x8Y6jqZieHKrzll/UjaiAsxlGWNB+hC8u14
3sxPTO7y/dEQuKIhsSIMq8oZw/kt8xP+M1QBNsYdN3e6wUaYLfb/78JUMNO73Ev5
+wvM9m0bysv3+KWazrFVVKvWaDVQGGuCrl0sgo2lpmCwNhy2ogTIGeB8WsM2MvKE
8/5SxlTnDa+R35M0lY4WpCaWe3EK9OdPJHHrrX6rxtD3hpvtmJ7ir62nf7pUH1XY
f3KIlq2K6G0IOKrRJ7CYq108kJHEjvedXXq88ENUe1QOumF3sDbPjHnw7K/UMCEY
NEgHoCAH6L5HEvnR0ccOKTNfHBdER4K8yUueQmDJ9u/FXPUR/gTXtHXLcFfNuVaO
G28etUCdT4wTx95a0kSCGLszOC2vVOtyrKTy1+eEzaIukknQmkjQLw0KW2tCu5vx
A/LX57sReyhcJvFqW3MX3/cxs9PNDNu2X0FBCrqZHPpD1eOVexmlp60Uno346iO2
xWVpVoNneX73tCmRMufQ10iZXqlihCkvWlRWRda0bH7dJXecixjEFq6XXrrBbyzW
kNSryIipFkfBjiMkmgvi3+v6V5X8a7RG9dSWuzcJirQd0OvNDfjanLphp8w76WCF
YwFAkBvNXdALQcrPmjMzI6cSQY0+63bXMcdUjNcMu8txjMcKkwtqHb2/izt/dDFb
mpyYvYhvmXNDIdkv4XBdv7WQ17GP0uH4TMuFoFrh0wRBsmHZ0yRJ4gBcEIAuCDJL
ETzDyAqZrlcK3MGFdPmEq0GzzVCATt50+C9+I+qzvUfJlqn5XTawOBWIaNBWhCAQ
Jyfl58EEsBbSvIXt2HtQbWfi3Gq8GdpcV82EuXuSAqDvV4bCuv/3+iTOecSMBmiE
FOGs85B7BBURtoyk+GOIHG+cT5qlIzTwAwW7ip+xt2NnPku22jmOnLwjzKbSO45h
ko1YsnppfpswyzZGnosLCYi0BY3Oy3Ps9LXlM4q9zMaoK7AnaYq8tx/jDWch9+bq
uNlCN+aOcFnhJYw7mm4SUHqkupS1FX16ArZQrWxIvJd+8X3stTDDMjsm74ZIqDQ1
5ulTB2j6p5Yul45l9xR4X4a/vJ01LrJ8C0rPIsqfMcwjYVagFJ/ZZ8TRxdLsR8bz
XUzS7rESpwheG2a661sJ+5SLyET1zHe0GrtyryUEBrF7NONCKusVo7LZj/gnHr51
TVvXLmI/WYAetR+f01nSTiYrDIXyjBp/z5V3W1jdc+wfTViuGlLdUTu/b+NeryzC
AzV0kXs57xcleT8asgD37JJVYdGtB3FmUssMMvTgVeWB31OeLjaQDSTHA8oGlg7z
V2ieydcIhPB04elacUsjtkRRu7fAZpjUt9/XkCqy4C3jZzn/eUIbH5jOSL8o+R+w
pSCUSUCYEIXhfkuZ8dqA1doPA4YpZBJP4U+0iaWm50trIbTLxHiCRvupvjorJBwO
+At735c5ZyrTVgfBRKtg/bDrt9hZVa/dIxkV8QfJlhfvdQ3MdMPTpOZAqiJc6xj9
pPK9GTCx4dQk+PCdNos+3MgrUawmOsYIZgkl2Y7tD+LZ2X4cbbN+tF7U136akHIe
lOspyFqc1Uo6IjAz2PyjGx8mrl29fcb1eFZUl/Ta4yq7i9DG2D5c52lAO1VwuWLH
dnEgvOpaA0aYNsgNqvI0sy38sZtPix+IUFhBJnHpZN1zttLTmxvDxUI/8Td5KHIJ
UQV+ULhrTKbZhDs9L6ywWkBabkbuf04aUP+GlGT+Wglu8IstCIDkIDq6li7ViSn/
37v6j1zDgyy8p8swlzSUEw44kNzYK7KbUmF2aL8y8hPLZVWFfMRibsZLrFf08xAG
VdwKcl0Kd7hUYMtqiSpDKSyvWJi4rsH/bcYvmTgQh/ZLMNslTn1e8bqw7h1aJJrI
beEE8jJacKH26+3hXduwGnbzZKOYziV+ek3AJ4yus8Q7uV9N/IoR2HKg0+wxOboV
QkqxlVdEoekBuVYhJMU8F+vOVRMZAVYlMG645V4RtuupUSMRudtPgv2gQR25VzCc
FoXbAiC6tD8pbFHPJALHCUSV1eBq8U2daT7kI9z7z/RYcv4nJ/MWvx8z8ie8z/VD
GRcupShQ+gKT4txWEUQOT8Dr8/5H/SeLC+BVkCOL1zqzceF0LS6bC95wr2gufB+m
bbAb8oYP5qcHHYNBgDuTHE/W2mQXYPNsFAoTefA3FV2Y04vBi8U4nhfZLz5dx9Xn
GH5QOzsgsRZQbZN1M2mMMEn2lrG/YdtKxfR8ZFR3GkyKMWESBuXySag7X7M67TPh
Be4ymrMXpTP+MAqqi25jtOVGT3WzFegvbhWi+BMrwWgBM53shvg5s4VhBDLMYJZd
/F42IVAv8aW/mAOfHdC+9f2KdBGU1VNspghZ5IKA0RGd5W2FV2PKBXoGISSfjJ6i
r3PgoOH/+H4W0GoiRRTJoNNgwt1gqqWjJyHeKgjmQgfv6sGzhswoK0wYZKloZGC9
kJT9BqJMNIiUzklLZ+7WUyqJu1vGKLlZu5L2DDeoLgRHaL9W/XUQ6sg5GcPkbiDb
/RtiPx7LrWt2hgr0Rr1DF2Eb4cWO7SCRnpRiOFbNireO91HCCuoDcHP62f5nPr9p
mGzrk4HVEpFqLXbchHG4EREIz65v2/2ii7bOLKIwXnvvWjZoAgSkiH6NH+W+fLMG
GguWbMR9NdDjEtVuFLBtZgDilRKGkYuAoXTCeaTCBpSeiRwZI3V7J8WENoPgBORX
Q+n94CDWTzEfJ9e9dNnd6K8bUAMawtql19gLw6iHn/CvHff61zel7ShZl2TjWdeP
vTPdoLbgbKs1L+nEmEKguHtX5NYq/DYOdoSqAM5Scq0kTyv9a2jKBQlkZSYF+IfE
IlcdHwsFG8SKW3vbHNoRUG/GO/Zy3ehZ+RMiOcaQkglITGTtInD8xGOR+BTVjf6f
1KZEJr2MyLccdySpThOf0+iHD3xf2mkc9UsxQ6uCOEjIHehtlbFpaf2Z4bUDCKZB
r+gfWrExWVFLa0xIXdjMIw+8FZv+nOCBHqHlH0HajOkzUAWnQMn3rB0jHpstJFYZ
sXDiYqd9v22rG+EGKPqZJNwynIHdxBfH9p7XiP1RM+XzqpPOOHmcLwsOSFB56kq7
qojJCh7nrkLqXhfKu5XLUw5ub35Ry57BkHa+UPbODf2d1Luu70Q5XdrZY7XGY3w0
tzVfHBVj7smBCDT06SnzAtkU+0/ib6bZB1A3ecUFVBoPO/Pp42P7E9AFNz/QT33I
>>>>>>> 426889eb8ce467b9c9a9f74dd4af433c5046285c:deps/flexrio_deps/PkgCommunicationInterface.vhd
`protect end_protected