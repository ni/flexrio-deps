`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
j9eMmSPGcKCWAR9PvkqZ1R001FU8QKTyJzFqNLn+qur6INyYDE1AI8LWcxAzfnTc
IpZG7ua3uuk5/kQKKQx8ZIPLfmv6H3t3eWjki8YIAtY/d5E7Gq8Z5mNxMYRzGGTg
TCMm6oOrOTVYlCXHE0X9AW696Z7UGfWirVibl8hs19hrFdeZKGiGht4r09vHR+Gl
FQQmSObM5aSK5wu5KOrK5ZUKGHyBhjnIQO5NnittDjOwxV/57nHVg0pdG6JUqyvm
tEgmCY36RCMRGWN7sekPtNHjqpZkmYrVX1T9QF3h73+8ZekZYd2xY2hpHHGYYeWA
t3+Fmb/6NUmoP8+Pt2hI6g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="wX+NBVcG/A5ruHK3pkDqG8ZVPdOz9TJPJ5saXZYSeQ4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
j/hqWUoxjK88VtH4QmjIrexFOSwtsLKOZ/LCP4cmrqgzmR/e71apdtoL+o8nlfy6
eZxDZMmrZmJGoazz2oK6kz7xJU85UCwNc4cxAsVxNdCP19vZxph/nCYZQ9lUFkLH
uLBkOeFP15CD3jG5/dp945fHP13J9SzB/L9PWvDC/gY=
`protect rights_digest_method = "sha256"
`protect end_toolblock="sqDZkaglKf+bDjC7VKm3lOELrT2Jlynh4UhPg2J0Q70="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 26864 )
`protect data_block
f9kZDbPp4NLiAOFOgATj9W35i3s4a7wbt9jeHjHVcJxMoXY8rb8laqS5bNUhXGW/
MOc7UNc1VwolqhkS7G27SLamkGClZZtXSbRcN1N+5kZpEaBEj1343vVznnU2Dre/
WS9HsWPXe5g0wH0AJA0FuGpuUuKeCkxe1CQfFOLDJlS37Ot19HKuP2gtTAAccRg1
xSO2HrJMpVJE9jJh/zULSDbWtddOpmjQ855p1QEsrqmDBbTha2b2GZrVEti6i6I2
EA52tju5o+7f33PBD6JADkH0CKiJHvt8EcC7jaJgQXr2ZFG3wXXvuLi1aHxHGIe6
K8RnF6fB3EwQMAkgMasCBX6U8550/p1gvaVL1vAjO+5qqeFjJrgaIB/K3eooCdbY
u/CC0YNE7PuHBkyisxbNHXDGwkgXgpcBXvlzpdkLpDpKKUfH7k3tmaBcKwU8p8EN
fxUP9UCARjmcS5BDXfN1uFN7RA6NU4Xta7FY74L/LvTBij968kxh0GVPsydjzEJ+
EfmuJtl4KFk1Hr7w1D5AoN9xFRWO43+6sw3evoHmXsvU9PFpHiHmB5JQ8LIDUvTA
nLI2NfTM2E/e2UgaamNQTPgv8UfL++bB4z3p1fyHFRcXSHfGONnjjGF4hI1bHodg
hW2FnAr/wV817gf3RN/oO+9JrbOJetFy9MJKzsQA/pGOXjZc+EMZSTiAErggLunz
lw4pUA6BaDkqMgAFJYwxxrE59uEyBvfFiAYtNIhwtZISU5x/qQCW55SRt/mWnU7G
pQFME10rnifqmVcRpLipxFSCLdJwFIvHFmQ5har5NA3cfCjE/OQCflq6CcYTtb+c
sP3tulyRDrbVcvKeFW28dqaIKjov1lxz4c90IgnIw65HY6jGvzNwbgeGc/vhzhgE
PTFiSdWHUAuF9mF6QtFD1lbz/esYVr3bloz1wfaUixPhsXfMZriwhRqiho+DwxKO
OeWB4VNKKKe0+rFfWjfpbbsm3lCoBZQBSZz85PnQrPNaE109jwmjnl2MTGINx7MB
ZmYcbTkC6iLxYaRAOwRelgGhvYGfej1ZbgDD+cJK75OfsFH7o5RJfy//UGKW3b+r
UZkFj6gNAUzG9XFlgqF4slNWhSM3Y/13rHPG2w7We+htBjnBKY4EGicihlXZgue5
tf4evdjrFKvOgmghg8yBUo/+K83O6yPVqn9+BgwEkKI3qyz1395wtTbmpyusVniO
8Ms8AaGK9YUoDOnGII7wmpVolOFKeUlKr7j7alqzXzcPkLC60xfJIR/SIg+OA6yy
vqW0XKldhBNu+VMC4TJf/z0NXZP4AhCja/NxppQriFPVAWSEEgtqTSseYh09Z7RU
tkGt/5R8qQVUo7Lk5/xxQYRrYIFpWsbFHpe55g8SRFzrL0WD/R8Vqc7sLpgO91Y6
81vcEevk2tN0GAP1tSWIMchOKZ3yBK0yg/z4w5XY6ocaluZgKy43a91FN3gGNFoJ
4T3WrP2SBVJIYUN61kZSJhcnvEUVwj6rsVhX+tyyVtgHORK2bAlTsb08dz9f613N
WoF+mU9nXT9ONWmetWxgo956iO4fmlVIhQB/yhXAXlwv83cI0Uq8KfA9/8ICmUFx
b3T0WMFM+DS0ptWL4CAbpG1pOGu7LA6Y262jIaAZ1illBsoRGgK6r8mFDVVmSAMK
Chz/y34MaosfuvVi9j8Z3m0xvI387w24ZWalvyIFc3aGxGgs0LMcdi4q8Mr+UPb0
eOpcSE9sZOzh2Z2puo/oXujQAADyEyPAQcInntVwOr8j2lmQ6DzdYvZts6D9HOPU
vkUSYNQEucbV/Zn9GCml8Wwt20VFYQ6VduWoASqHhWquWOGkD2qCaFtLrqWXE5QK
/A08319LoqrkeZHFG2Kd5AKfeX4598ilN020nYzY6pPPD+5YoseJ/41zR0jguk3q
24pMZ1a9y4Td5jyvBcupcVYU5pn4Qzlh+LenRNR0gOW/IC7DV0D8E4QHoQ43RATq
3JzG4/WpG8rEFaXwpNlhR0k/EdRWu3Y6B7iGhJekYf2v2EQW1TKVVR7r+OuPaYoG
TgBt+HTFIS7qhm6PC3eN/IJHlfodTLIU2EgKtWbq6pOeNitd5WuSnB7ppqdzFzn/
1EyHknsOO6V6RzTgIxtnwUlsppIFEbi3q5yAv2QdHyf1+YD3Z3n4yQTJQNxtJaJH
KwTCDRw/NhMow4DrAwUQ7y5PdANFrm9u1ahRhE+FhCnaQA/NVvZYJb23BeeTkgGe
/j9A4PUysWS2avdjyYn21mMr3OSBbmKMVqHu2eVOuKUmPNjm3glKyGMJ16WiXKKX
EUFK283RwKlHsiZGbIzGQAp71AROO4/pAhCeMz6wiJlsWAVsnNM8du8Qli01GeAl
X2Qd2l2D8w+W57kEtQquBITNsRQwRTya4iLOIHcf5WsPAwaMZEVc+NDHsKBTAEZ2
rIo179eliBUmPEOPbVTvcSKdq6PNyhNAo+G8jUu4jLuZp1Sk151sTmwGQg62h2i6
4e5nFqf+QuArc6IGCyT4CF0ornTFJD0dDdfsmOfQMeVVqJ/iiS3ncFmuGWiHLNys
VDGfzswCW5/hQZvoahUtQTXMX5enbPkcZr0pGiUsqBMA0NBU2gtpuEMpDVAiiOik
NTRF0o+rdOYcTVZlbXZnqCHEjGEV4u9DIAs0loG2vUgU9AjWqypbS57hq7/Db2TQ
DS8CznVYeUdX4ff/0ixzray0k0NdBN0lRyOdU6DqKtWn7OlZ8JOk0ywHEHWXycUa
VwPYQ+n3LnaOur/ScIvgCqIGnEdF2x8sSqGldWXxem32NLmFJuTaFDi4iVhTb+yT
dWGzJDm+rjPt2uKPBDHBT6S4/kaPE42OTzRY9jJ9BzzjB9oPM54Lnvnc2BICOy13
UguWagvI3mVe8aZr6S6uI5rLBABid7WPcazEY1QooMVP0178XuBsAnXFIgUaDN6D
yJhvBDGSUU741XpsK6GSblcrrVnfEpHmWzZB+IqPK53W3qawm00lidLE6YYHekXT
wOj2IDJ816rXwPCquZs20tLuDqHUjPVkL457sU2yKtiIg2OotHTbzEf+2hwpNn2P
9mr8HGHS/Odwt66ldj0beDsVz7+qCXletSv7cWOCsYi9e+CdPJdF+zxUGTGuQ/hh
FyJ0K5cAAEOpKYtuKs48p2BUdObiiCF9WLR40AOkLejaVx9BxqP4jc80mLByk5xA
VbvB2FZg8WD7OZOVkHj8cGx31beplbCXdGReH1SzQAgrF5KJVmbahxc5AkUttyht
L4FbAM4xOJB/4sdrUIe5cFszUVWwVNuWkSlNd5RplUta/e5CZ+wJfN1ePSg3IIB9
hNgCRCED+FXSNrIHKG8Dn0LBSGeckSV8NT393KmC+VHEpWj/0fn1NOnSncHTsEpd
YICt/5Yy+nQ3ne623rRjOLEPfOtcx43GRRUOVecHshnIgOOw85Ndz7cZI0+AQwhl
LPOg77k4i2yEq1m/s5sHI4WcLeGuomgiU7Sui+uE6L9mDHqz0ihpNo0DQ2XmaNGX
oPCSWJJYVPx5jRL1mlK/fZqTcwH1gSCrBfrJyB3q8rwE+0ehzBbYsBAKy26A2V35
IpFv35KLj2Bm91a2IYsnT1p2feSmmzrohJZCvwsS91B3ZaMxAwHNL/Wn4sqWV6sI
RFwzvtBXLHcDmQrNFGC0fo0xxos2sGfeRdtG9NqEmHVIKuMWfhhdAFHwsyZDsPL+
CDjhUe69KBUBPk23rPfTnHSrCYgA9X1b450JT5ptyGNLW+UYwQRK2cFkz41UWDXP
2IN5BEiSFiZj+IAAW8rXydsQdj8wHhOPIwpp5X2vPskDANzkrdVUs36cN1HWAFQ3
oMHOg7GUu8Bh0wbRYAYCS8gcd99dC+an2How0l0JO+Io8M+5233+n/LYDxExIL1T
+zskcAHi/KEFTWCQtp/FQademSAdDiKEX5CxgENXVfiOTvA42wVKQmmhXos6qKCT
HdVod9DwhplaXdaT/2Ndrn1y5+q2KbjYMDx0Bb2fqEVMGCPqauWsgUcN/9nZpzdR
aSCz45LqIixpXmyMuIAEQYJbW/0z2sN8MVZTgT7Q0/z1u1I+yIqrKSfnMx/RAG89
zhxlnuwQnZjkE6ZnMytXZ+IOa3ZLdrrkSdCFfPIpUcnqNB0tY4kOvulwuph9T4yt
J7vSjAUcKDP78wTkuEx5pMBYz1m4xPeSfb2LkV+gnea+4NH1o0goJa1ofyLGYz8B
MzAGh4wgg/Q9Zb2gd7sTzJZvAVcmvmaoCZSibzZeA/ow3i93RahCHx9B34Zacz2L
eeyV2Qs8q2rTXK7a9lsdQb1UelljuKC8DK+xdRJFmJxQKa2I62nYAsl8LMfIArgO
hmXYixIfDcSPX2Vq4OsAqsrQuHburRojpF2Rkfxi4wQHduh/OtqSTFsRlgTFwe5p
U1hZkvPfeAPoXbWCoCtjSaPZVrd3iHUG6csYI8y4DJzESPrBsPjdUMjte+3W/Pjr
GiNVA9O7VwcypG+su9MbQFe+bgLV6KpXMk+77/B7LLQaRovRRe2F2ZM78XxRVw3p
tMVGhaE/TTXDkJQeyl5LRMXXO8wLGedgArTOVPl0lQnTwCfBiVLiltCXstJ8Kpvs
StZzMr1gpDO077TpfdighG0z2szXd0KtcvSTXWq/6oN2Ile/pZrq8q/I/m7Sw/Z9
HrYUasc+vz/UAy+0SWU4TMJIxyDHji3bfQhA85sUOkt99V9VKwqLQJYct3ia1bHi
oBHVD9u2Hhxz71SystfyjIZdWRBHpSkbRNM6CYZHabriN7t4ICXrzd99e+C6jyZT
aXQf3cC+aMxjxRdG6Sk2eEGpl33q9GSvnQ4td4n6sVt2cV7MPvJB7CMJn15suTdK
cRLI8xC0yb4EST7IUNB0LTzzvDDL6aefeyid905bzaxqvsqFJPW8635+1AoFHCVy
1GD4DvgZkPQtiNQuI3kpHh65YT8FLOW8Hu33oKaBv22Krhei05BUAaVyQhnNQcxY
JamKwPoFnZiIEOAB7YmSJSJHFUrpXSY/9GXofDIM1oaR3799Osggv9QgQSKvw2p8
QkiTlTokffyIcq1xn4gZ+l0jGA5Suwug7qd00XswwMQyrGyxjuF6E6n7hfGB/gq3
07PGMDNZhzSfaNOzOqStAzaHiqF0wl8zXVmGzURksdd9+Vkt0XuLfKxsoCnmX5LC
Mmd3INCnuWbAYZs+5f8J+3amOyOW23PgJTit5tLnxRjELWcpNtgSxyp/FImyoc7h
E33KEw2AdgFLnokE3Qcn5ZqKIPKuKk8SxIAWP39CTl2UE1GftA/MNc9tA3CTXtqB
CDmnwIrN4/HJvOqzSkkTeJNOfXAazhWcYaA/XFdeSB13UHd0U2y2j4dMqQjOVwyT
/aB1lndEwFDlT+8WM+TBGdQ1G4XjvR9+4zxfJGL9zYUFM1OE1Kf3gYa6Sh4CUKrP
2tahFYqZ/dc4f+kGGAnjpjDCAPpzmaOX52m+D7DyP0VkYAsZqA/uZzywOEFjQVld
IqQu/jbMlGSM1dhdjcb5nxxvY0BSrBY6DuupmxcRh1nKv8n6+ZntQJGqcOsRDABn
fbzVbLzj/nbyMZobaslmowCP8cbIyQkuKBlsNXT9cdtgf1H5zNMFQP9ssoTfh5/T
3sR28+i/yvjrNjCuCd7oofMnK00b0QgeCiqVeYd0cqtcqahAhkN49qjbdN8UiOnY
tmk1srCs/cIA0rfyt4JMzeJOao+pIiYqoKXX/j5jlF79whTbgrvp54JQXQGHnk4s
Dgm0WSaA3n56q9r9fTHCjdBPyEsZmHhtzkNG1YI/MGR3X0yRrvnL16Lum2x/yk/h
adNzPekRfJXo/5UXffCAaPqFCR8dEvT9ih8H+NjhEnUy4G7br9B8NJ2U4pdn0AMS
wSGpZuhLM4Nz1JhRp9mXVyxh6QN0A2yvTA+7q3FbnK/NthPVP6YTgmftd8YDYZUv
nNhn5pqte0N/emcTQGhFzD81tJpwR4eIlDckfO1eljK227RL5rAuaF2cGba0Tnim
s2PJl7Ll3OB8AwCMwb4mxWqjyGHelTi1DvD/GappQZEJyJ1ynW/m+w8acEPOERXm
H+lcQ6I+b8Huj8sAxp4QgU4+rGccyMGBfGoK0Lzm4aqmixZkVyrHUFNeYfBpmwh1
SwcjuoACpiDxO2L/ffTsr7UpZ+Khkmk51XxFn4LDV1iQX/kSk34j+DoGCRTPnCTF
9ylsI8Cx3mwKzkl7RQZsOOBpWTFt4C/UgTXGNe/QdQDP19yYDM18uhI88uE6XMD/
QljWm/dCWK+k9xrMIiIrx4/XJyl/tJhw1enPIa3dTrK8yFG1TVggMT9KuZThWkga
v4tLTWjOVEQdGT9j5rBvsLT7xqpwB0WsH0d2M++PQyQyGZbTFUq2eeiPNRgnvTRm
qwdYFpYHXjzRz7vuoWwwKVnFh/YSopyCQjLI/5rOt5GMAvix37MZR2veEIibDrib
ZM+DLVLt4cQdz8AS7pMt/wUqJDzrRB+mIz3oR0gGo/rYq/WApGdz/v43jvnyf8w2
aORs4yzvPZB4UTOTO3qpTL/6Bkxq7NP8CrAtL/OTanHd/GBysqOHLw5i7OAqrcd7
BYXI5X1NtxP7UL/tJu+4i0OT3qtVl/OS39dZovxopZyyfsIRagKvrKYEW23cHLMB
YY+mAPm6nuRz+voUqP1q+fCsuzzO4MmOh++bLfWquk8yn+gev2n0Kth6q4bbM9jV
knPWDgQhNWSRMWlDRgJ3wXHNYANiHdyAWG7MnK0NmBYmxj5csYjRncUMlt4bsxcx
DXCVJsq4l8OtqdlUpqxPjaQBvK8TmmYzsa+UDI5haZppPkhLQlKuUfYzYMPcL2A6
+A9LpDPumwjSKwcLxUmgurFvBIv+SM6yHwsKwNPETtlWaWeMNpzRhVdNbBtlZh2f
cS5ARUqOKg9GIHbC0uoVDWW/9oZXf6T8/lGFxE2J4tqhhXJ33/cWhYFH2EDoOXvH
oxJAIlcRutLoMfo8uvYLRNpc8alo/h6gdK9X/vn1/b7Ozfl7qG7hEdCNJYna3Dpf
4iL5FPK/UOoQh4kBXoijLz1AVsrFQpsgdooQDBuFGxkVSkLFvIEBywKairYI01mg
RMNcD/H3dGCDLEH+K+zwAI9Chba631sHM3XwhXEo2R5T9s7REs7l3G+wUgiBVF9W
ewdmPFNSGNi7EPio/X9wn4zafNQOW7vRIub56lROUZF7IkfsYO1zgY/LZtKY4NmT
sCCHvnDjDli9RECca8PNSBTkOc6A5qCm+AhtfnW4PO7QBcyOk94+iZAgTj9lU0bv
wPLbgx1uU+Z8g7j5UQ0NOEHYVv5qjj2OEFGWnJhmnYmiDbslZnGRHgh2kB6ggWnQ
CaTUOuuHOS8bdGI/PKKwtrHOzUp7eLJDkL19a2G+jUdOvrwQIbBcI9Y+sMQ0MGua
EIPWQcQny6FtO8y1Y6LrLCoytrsI3lvDKtfXHHbnJBSfiDO5i6ezHH0U1DgYmhBE
nwUJHeYh68G1P4aMkj2h6/5OVd1yVT2aVPmeDYO/P7z0ULWsAPqZUdlFOdLManva
34+/fNBKSUhVT1jQfXZIst+EWPw9ux56x5GqlhX9xgRLDoonVpI4z6gkiC/gM8ds
BpZTMUd9LU+SyzzuFi8IJvjwYyEVGsAuCjCAtHRQUcgpNH5QUNZo2DxlAVHvV7UL
WJQEhu56er1ZQ4EjyFrETjxi3fO7FfRdHStPXgaG1GGYeF5jyTQpREHpNnWOyR0J
c/9Bsxq0jCLcz7uXVcf1eIpadKqSdTHiUVnOFW0TuBOlbg5TLdZjsbjO47xX2bB7
SFFitsuJLxLHwHCQrSrOyTalT48ATuBhvXvQFXj5oBM7DFjUs3iiwiezTIIdtwM2
nxLbyJ0WaCIGFsKcvjFvUQl3iV0JsCPg5BT8FDiV1SIMXgALYCpuE7pdDyAmN+sw
B5tSzrI32Go3VVzLoC2XfA4K/pO8/dfw0aaIkykxsG79CXnU+olk6ICwss+YiTga
9WNkPwQ5v+1Fgbub8/PyL8ZbkTZHgjJNFDktsI/LidNOzirmH0VEFGu0TqhK0Fw0
Mh1OohTDvzcpjtLHuUuqzJqZXba7kSCjQFyda9Hk3edcw3sFBtiO/lSGCCQ8McV9
6QHdOR1dxMqyAWvHzRbrXo9woANnH+0APwTi1mW8l3xZMj/doRmsrxr7EqzheE62
50SM7DuZKL+p6pWQ61whH9SGW2cs19SVrgsWsOl/tfSJcTMAlyqhl1wnIEsxzUmV
d9z0OfUaX/GWvUwInoR/AP6Y29eY6vtYJk1fkW//PN5sSjV4GwJwchH8yMUe9pch
YHc090X4T40gHHw7eA10ownvi0ygyNXyeI3MC6royzMrIx7GHv902X8TWrAN5+vH
f4NbyW43MA8E7mDB8M8CQTLv8TClkAWssnBDOEj0Xs7zWmTJ6AWv99dnCzwf+2sp
y4bQ7Czd3PtTt7miLEIcVT69nO3UZ/HdjpmYzZZb66eec5byGP93mnCENzUdNT52
dSRJoXKHWIUqyDFF5b67tmI1L08AAc7hDc8orFEGqxvoq/d3/Ckte5/vYyxt97vY
NXFM6miImwo3jNvIDhUdEuJ1L6gswI4pWaJLQqetQXflFmSHvLC3RG0y6odkw6ON
/sOv2FhMZ9gjWtqeBixmVeF5DZ9fUeeiNYqxUcFoXt2Laev7XBxLjIAaezFUSdWS
nZ4TBZL7tlerZwLNOJBcrGSNkSITCm2P/3l1KFy6v/KtdfkbPUEaa7DCS4DRLaNi
6cQGreEhectmLYk1ffDWJiQr7v4nIlLRhf1sAf9RPgY32zJ0LCCAOUPVLGb48s7I
cEgP+YfvHlhS8IKDj+mg/r47wn5Gb+dhusN6HQMruRXRivYm4+5cT4IgFlEKNeYY
U7vruTW60cqWNKbdMNOF5bKn/l2STaKgHdMsbTZORcKsxJHMPpejJOWi+MJns6fw
kpdDL1nBnSbz2TJHot0O86QCNTUEooa/LZywieEVVV35p5Fh01lbyMWle9Zu1oGJ
/Rth4ASTCA83NaiF9yFKrcetWHTrQBujdek/sXfZZHqTk5BKIM/tYFQ6mNi9UZID
CtUCGXpyw15Qoej1fEi67yHCKIf/b3cmI5OU78EiWDPBsypO6EfZOrMLtgaTri0E
eHTNK6HU+lSpEw591bEmlggK7g3WdMFMYB1h9sHiqSv20nqNN36qFRaFAT9jq7Bg
N5uPI+I+hSEP+kqy3ku3ePn635CoSvAcXeV9++DOTjCKS2wh9ma2QgRQoJ8Nado5
KqAXAnnQ4ZQRncyN1QlADiQ0/FKNZ16skm744n7YEQ+lFy5SKKu8RYCEg7DBZsvX
cC8QkvgG/Qg+l8Vt6Mxu1V2icFsMA97nRLYZj9HtAFeJms1mdSc+0gmaewKfmKYR
RD7ASb9PMUVU1TKJTtpDIURdjw5WqlmS5BAu53W7NiUXv8bBFz8EevFFw9D4/fZG
aMUct8O0GO3lSXFY/vPp5T5llvdvGJJAIcTWwM+7w7HICAwCkn29yxUgex5F8/Ij
N98V76GCepu+RWfWjfJYbzppDGxNaVKiDCxAI3AEcwCUm1fmfZHu4ciJVNYYmE5M
oIkPEa23pgH4ZUEzeoYVA0CD7HneyQpS9Egmy/1nCVOLThh/7N7I+tFFG/7fJS7+
BN5f8CF2ScnQVFnpjPT4TE0wbC7ViNOZ8fk/hOfCiwyjbS1mMX532yybmS1leA9w
m4otsPuxP6G8qBVso01GApEmJEfvmr96F/GXaodkUDDko+3TdirEVv8IiLdWn43R
B/RiJl/9gQrzjgjEKbk+ZH8LL1DXcgcDn2p8U0npreb4GyEXkl6SR28/Ckat+6eZ
wL/s+P+EBtfysO55mgn0XTY7oMxio/MzcoSK2LOHtatLk3pc6FK+jC59KFDuR00R
gyajNkjZo1/7jQaqxDFOTF9GcGUTYwRYYlWGiPu6DYe5XmOxxsHeuMxt2G4md2q9
p8E2fAkz0KGzlAyDaGF5nUaFBKomuSbrw9LdwY85FK6/CRo3Vh7wv3w4QDdvbNxr
P0XmFIW62Frk6O7XNyRe9Y0ilFVD+KqoddFGx5dlcZHsl0+mBzUwZhiSUnnflkxI
O1jp4MUJ+Nt+36Kz7vbFtRxLWwErbGJdy67ZN3A5jRHZWlb8MafdNNifB5+uMeBk
MI1I+vAG6Mwh81q7mFA3k2QJ4ZDqmuIt9MVKd4LbzQJP8sC+YPpOwOxXwI5txS97
XWmaFUF5Qgup6pLRV9j3tHuRAuc+NkE7y6HD/8IkW1xOvqGuRRWTSD5GMvfJg8E0
0DnZkT/9Afe2AXPhn88LSJWFmrHW2DQN8CEwu0caDN0YMu5M3jN4Q9vWRWgkoEWH
9CZICDApd838CUHm27cIoIn71xYU6AYpw5OJGuLEtKT40w6WfxNbzmuQgg/y0EY+
FZcL0omrkBjEb5dyM2sWZDKSihg2Xf1uT404iVo75N17Lq5EQe9/qUn/9wCJTdSF
i4qYwd+xeuP3OTBwotEhtrY0647Gn+gsnv8fcaZZx5ZuS+qFvGT9ln/iOEqWpoBy
+ipSqup4Iv9qy92qQSGP9xkJOxtfVmJmNfoJPNJa1/FpJ9UOvlHhBBdh6TElU/So
4YnXzdw3j4rOfW+q9CmNB1PzvkCKpuA4EIhByXbpGxE0ApK6a/rZE5RAjrIiwwOF
xIxFHFM6M1twwujhT87u6DELZojaNXIJEEDwBlbQfB/X7bPbEQtx9jwc+EHPjlI3
jGjDSFMxDJOQNbUGQEdhAy9eTIHyPKu1gs1Db/rUycWBDhDSxr82lySgqPHyTu6k
nQl+XSg+TRfF/+JOKRqHoxNYn/wWVTa+4IJUNatFtsoC00oR1qfRmy6c33H4hf/X
4k/3g1HvOVxbPs4Avwia6s6eY013OdlV8X9sEpNvRgTgbgRhJv3PRjC1ABsczfQo
8TbQO7TLswSRDPvOOjIAdIQYHZcSZsgyyz+KlnifuAK6Cvumjb09ot2UUs9pW0eC
NTJNODSLNXmHN/dzHpBjm8xDxkWUV/FA/M+FHY9Fj9pO6Shw0yZVWz+tyTDNayOG
WChdPb2SCIyW1cxpXJf7g9fEHa8oLoabLvKLTdYrLQrVGVUpwbk6dTqnm37jZ1ZM
ifTQ52lxuNv0/h+Cspc2++oYni4SwBIwGlnscsE+PWA9gTq5ueDMBXwNWJxBxOZ3
4E6/aokmzUrgmfWy1hsyX4yrqY785m34W7rhU9utqN4aswSKpeQJzFlL4udryA9L
dP++2f/OLMUdq4ruG9OTD9jPJovoZdOnfDZ9x22Ur63JsTqG6zbJbLB5nVWowM2o
zJ3/GKTWzFH7ZDJKD1GvkhuVJk6q3ngBIY0L3as3wx0FVyZfAHKKxmTDKPBfcZj3
Fqbz7Qo7Xi7tOw/zMsmnaT/XKYYGA9rTCJg3niovlVSAOU/2BVCAAmhGAIUdb6o2
dGa7m980EmrHi5N650T0hShDgItDCWu9zZqB52thYtnbdbjwuq9Xm0l9oOoF9lbw
ROpBsVXyXYSj66McgANO/i1FOj25L4EZQMMT7+g2UJz1OsO6rZoZLL46ImPAS6xh
w4wO5B8KBzW2PI/qJLC/CD5XHniJsph5LfgqKWYT+1kU1Ud7MRgnLxEcThvSr2EH
EV1QoOZoeJrwUzXbNuegpjZce0KS26DR2nlGXY1JRnUulMBy38jLBigiq8nzd3Ws
yWoWwGqL6Kka3r/DNlfBKkHd1QUaM015gGwblZyuVrB1tpPBYuL2umrohfzkoPBg
nI2yp51luTkIgJqdvovDO4NKI2tG/VpYNmKF7h990dXD4czeQGggj5E4vUACj6Tb
mC/zK2YL+j3FqUg/Sc7c44EhYZsnCkELPg+cIDpQKk3XHKCbFNvJ3yCXCKYqw7vG
ET+JMTf718TyWTsODtch4+/NHEtj6eRc2z8RMsUV5JJCZkJKCGop8p5WvCTOfELP
AOmLeoNu1SNAO9tWpAV6xg7Bko2a8xDvTnyyYgYIygo3IPn8mdJo2EDV7OI2eW5E
1oR1rvg+D9uwl6IeCUktmHDvFbrbLlTOobgBjw6GQYKXMdgFyc1ajFgj4dBEKTiq
hw2KM9SOMLQDg4jZE0fssBm/8H3v4lVqHJgjjBzv9ZoIYhYJik90nFeeE1mmFntj
V4gk7MnPw9I1CckX9SpqXh0GnYnV+KKs7TramI4MT2gNeH7QYNQiC0zb0g9JMX7r
YiveyK/3IXBulWFUmLS4wDeG8IPQrN03MsNFgupEesKCSL/bGnrF5+qLsGW1XUv5
2XXpQnw6CXfJGJtt2TzDVgSLmSwKE9KMiK9UGSP1b8gKUBjrfMB+wJJRvavLz1CG
/3OYNcDDFeIV5t/02GQMFVWGblwalBtpvcmR+8y+/UFBkAwYjyU7WpJgOtZlF7eM
1yHVBiluJCnbdibXnLywYdo5tD6TNvITZW5YoDuRaOCf+w5q8w7nmxreXkPbGOqw
wu8fKkCV2EHC/K1LEr0+W19NVre2huzM3FXawbtayVmFdHyfX63EgePYtS5LmqiM
+SQZhml4sE6a3TmkWQDa7Iq4GL97+LNA0myGVQ38hdizdoZ1fVcWagRAIuCPrma/
pNm4DTeVzcsHrt14eykzzBKj3ZG5Z10mfmfnaC+WGX+4gHkMyn2BQMgimM2Vj4Xo
eo5tBqAb6Uo423SESItxovb1m9K0kQm9NfwlE+Qxx7itRE466yCiSuSI3tBXlMlp
Dqse972LYDSMabbzq1zue35wYZFB7Q8jAEQELvToLN0BzKuHs8HNtVEhBoJHFb2S
y8vVjAvPNzr2OBSdlmZlGXRduE7uFo7mxTBgdQwK68D+Jkl1U8zNJzOdZ7sHzubl
fpE0RVluBZ6uLZfQBO5eP/hf61VVrdTPJY4NZsEA5F/nhH5wVrRv2m48uV806WJv
Z4HX1lFjbfJWqW8NBNhMnBH9XOxhLPE30f2T04wvxkHokjTLIdIs/8oZ7jp36yrD
siGDrsV7Kutm8OBKu6gDAwhtH3/Pmdj10+g+2yrtSz0BY7xR1iGiMgUlLGNPeQOr
6MEbP6HURrfunsp6LzyD6SnNsseDE67bqHYf1XxBLaInUFnXRuvcrN9+43frCIdH
UpBTKErCi4Dzv7e+tO7CoLox5jPYSuKnhu8bntkxhk2crhSPxi3rW9IGHqZ5gbax
GGWbZGe51E7T6g7XSs15TZTF0UYH3B1wFUQ3I0zvglIv6CGzDlg8rmArlCOf5DW8
SGF9q+IYqC9lZGTHDDPwG7sHtdQtvaUURxHIE7zbFaW1w3vstnl+Mxs7jJQWvruM
RggywMWf4wLGscX0P7eyHzrCCNzX2ALyom6Afa10fAtrjiRG4RspKSt6l/kHhncc
bhTgfNdXLTpp8C3ddn+t8B05chRuaqxkUQ45hWWqzs8oMZ6hXrWlOyBMnOhE80AE
FuGWgDYjAPTD9l6//U1qu53mJrSwwsgd+yv/z8Y9ZVLxr7owrPcTkCaosImuKg1u
bW+9g+UQcdchWcZn76zqNQIFEP5lwM07MyU0UK6LxaetwHKo6f1Qhl1MOcV3xDIO
EkBzeDkoh+2cHqQGlPR1Y5MTCTDnScxwcYWtcp6SfXWA6WjAGWGya3D6i8DONxqW
KclHnPJ06fD8xStjZ4N0SGQjoercPfRlga5urOZXmJ6o4mv7fdhYcy6boWGvq4qg
g3ArVzhAy5E3Ch8GrOYBQeqN2eUe3Z/vgX/ls22N4hT3bxYg6n9cX0WNJplS0dBq
yVBK08Do0rKvRt5IMwxTUDN2INycXLskNoyink+e1ki59eNo5vH/u9kRkxx1I7LL
AexmTBlWucaMu3dxRYg2iDjkvL97ObLVq82nH5E1j9j8gPiMo3sGGFDk+Xl82P2y
4IgjjkOWt61wh/a4JrSjMvj7XKbo9iyDi/oTyMbNYwo4PdXzJXqF4Dj2UEgGW/G7
VpXE6/MAGDHGsn5HT58GQsXaJ2xUKecM294bKo915wJb1+9g9QFWG71M1yanYENJ
xEVB1Gr4ig7wM44UiSdF2Dqc6I23+90Fj45PWteqqwJe+hpC97Ae8S7U/C4JTZKh
RX+WhlKChhZxnvQdnhsR9L72LKLJmrci5JlG7oAkZzgZgOFnZMabR8pYoFKcr471
XpB3JMNBgPhp6HRgO3eSRNXm9AhecqJm8+aqvvRolWmhVccpwBWeP+aMoIOBgIdH
zj81BNjD33YFEZWkkuBdnklnGqxj9F3IKfhnmVCyAKNOk7Ldf+Nf0YtxnGXOFhiG
gWi4h0rXn0jybURT1+T4bzkDWaql0Czm+pv1LIzAMlwnQo3XeXL0syNNjV6qxzku
BWG2WHe4UXhmDoVBXDC6iNRsOG/R4zL3hHyfvrmzATeObjVMJfdw3zNXshogyn8R
JU1/Qk7mSDVfuDb+eIkMDoQQh9RGkfD5ycOGWmjU+2yStPNkip6q8sZKiH2Atx+y
a1V6qX5ncTjGVGJoLPXBQD7soVhiL2fOQdgBuvg8HMRM05Re7CTgdwcXu0BqfdTb
gS+VqcoHSANX2xUsl7RFVg6lJ0X5VlOqTSoBZexWwC9l/yQaWmx7V5JrJuodqvIQ
p0UTj8kdVaUpGjXSldY3SYC9UsA2FmslGuySJP0wTs2Hub9tT3Ys4vmmtweroXEM
N4uyzqP5+Iq7vXw4HR3c4NnkBZ0GLUrXI5wLWbMxG0BAUSEHnTYB5vOpIy9WnBdS
8jljyTJQzURtiwEIQTWalukNp7cr7bwnlA6qkIHKXNJUo3QTidJ59crr5MbjWT/P
G5VGPPFVmDehJUIUCieEVhyVbRn8VDrR8a4ijdytSfwtdELZLpKFl9tuuT65qkDL
Y4cc7ty+Z5DHL/9SDOmMPdg5/PzYK9525zd0ohTqIzODiKDtFKAWx2kkFi8W7NCz
znj3OkDo1M0/R45nnTk0o44fh995nXrGg5WBWNQ+XxqXPBPTXUSoA4wQ2+zKK+OF
xsWcs2I9jvsxGOoDHZENzxTpwPNsay5smqKqCA7sckMt4i0KzZm+KLvYhFwAVPWk
zK83bsXnS1CHu/hcPkK+i5DwLfdp8c8sJ97VuPdGVyHmd1C8JbZICnL3QN/ynVgP
veknPtrN+YyTMBikWi6oeHP0/i4jfwoA3DPu7494g/Oh811EO16g/sBiy57hNTvh
pLQHc82XnzGZZLufEHB08ywG9atNjgJDm/vI5VCivxVNqzRU9Uk5S3W40QPOHsbA
Ph1lusc6Y5lsK20xUQOEGjykCP4eKvQzPPcrJUcKpT+XtEHcxZu7qxhnphUqTJX7
Bhw3BEo73WicU7t6/A3uZQSz8H5Rh98orIU+3AfR4vCftw/GFi/GquXbCRNHyPfV
KcCuyx56m5ItzuZm5+ctBAtDLGGawEJA1RJAM0GEXFKilJxK9jBEnu6xNCRSMWy0
SzQQIQzHZzoZS4tjy46WWqs4pU3oNKzYDLTrugcNDQdzjQ94KFiI/ZpgF3qcWSH9
DWpZ96BzE2pXE0S+I6L/jZj7gRhS28pm6WamCWEhYkuJDj5pqF9UjAhK84EmrFVR
AqZ62NHQp9JJav4Mp/US/keEgiXTWDPwLohgnEsVr+uIbkwPcQkvaDVjiEyZA/qo
0TgQzRK4hUcAXYwaXZgxptUPeBb3Cnkz8uRTbRgSOFb04EoUVp7/yLJPr/kS1Cba
51qVKfQn+qMd/ld4geSaKTNVT9zzMo95xUi+e7Sfcy7PDfRw/8gQ7tx3NststNAf
Dq3ICTEjvRhAkW16h5xkUr79PI/d6DPGPiZRgQYHf8RqDy82LyDW4/qylg0izH2f
t7wZlTiB4gofoPsh4pnPD3XaiN20dHJeZ7qaGsJM0qqTbvyWRQQU12nIHKFm8L4E
E31LuRBy8WvUplkCzTQbES83CKgnorfXZxgEIVgK5/qiXNv3PkmLlIWHe6Gs7i9d
6u6SOHqr8d2RjysMNBRy46xH74H6iwqB96XV2zIg+v7fyoCcJk2c5mGDd9D1YKTT
m7NdxyuW1GrTzwDktk3ZLUhmpDL2YPW3ScgU2sR0ferMhcQ5slAIB+1ihJB4VOpC
L1q9mPzXrBWKb/5NoklGkw869EoLQXTq3N3Hk3M0+jmM1Qj1WKm7l8dwo5BkzGJ+
2EBdLC/YRVK+z6H09xMKGtLIACc39L2dMJw3efeoTqDQ6ucsv/EZeCBMtATQwvtK
ICz730kZrVLoqhb0tU2sFUlOuLpq3vfRrNz2GoWnZtGsq3DQsIxvEKfSJUkTY6yz
TgoEgUOdFCgkGEASBULwoDecxazOqy4TTCUbMIs/+2BMpKNyhUfcvreLMMX8CHC3
V8yaEqYUm25qZCRljPSNXoyPX1ElZFAl1axKQLVyVpbzp8T694WmMtpn3fe5yexr
YWjtQ6u0YjvsIdl6sV5M3Jqlm+lGV2oTdrkYtggj4N7OncXRTSEVgv9c6NVJBB7/
P/oXekMP/CCnqyIoC0UjgSIfg0CgVHE6tDzZHb8EjPPygzRtXFJGrnEEtVZ4Lqv5
IHnt0uvhTlhc8zgGlwEhGNKytyEG8CfqjYgUJhTIhOotV78WCd3sXc1iV31qMzeE
qkYDAciY89JCybTar7tuIDKGbCDnW0F5JBqy5AZSb/pSrd0a7Uw3XKf+frAO4+Zd
y2vg+jEswe318/kin6f/UvhL4k+ClTrlQMXoewRm8coeG1h5D7S9yvudslN0lMwj
XCeVwnzenD4FuPXV6QL3YVCld7fH3Ue6B6aUrprhSWJ82Xr8ZaBmmx4F64QxEAcv
OPEyKkdzQ04lMiv0/roUXs8G41w89KMhC8+4fmI4WZAjUAb/bSDsUIXdxLDm5VW0
8P8bq9a0ZCgcOuCcFekKD5AbZbVYGYJf6CcU5pw42R/ZUWY6WlMg4PTs/zJpPKdF
WBNWVRedPNrI0xM/nsxEDIw4nNNQbZ4RtAGDzWRIPTiPk6OjDCU4ilrB3HgtM+IX
f3+1achszNUUGz3V9kugEhsvaqDhNbjI2qjkfnVCGzp5QNF7DEeKBRdhLmcvQK9N
SA89MkiRRfpYVMndNIgv3RKj7M5IbFDJiU715ATkwruTdFsjdIJ7rRMWrx2691pJ
8PxW2iRhsqAq9eC1HeN9xDyI+Wz5ulFsQA38oGa6pncQCHdu84T7qF3xUxFxcQBR
PtyK61XgMMUjrXxP4z/FYhQKS5xcNyCrIMAlwWGO706uK2LrVAT4gONKZDh0Bf+r
C/ozWzh94l8BN8tt8iVvkRC64GPMTmalXQ8McPb2qy3i7j2u5vve6h1ifhwFy88o
Xz0hwdMH1wlO4gKyfWxY8HlUPrjwOgB2O3i5y/eIFTH05BFB/uf5zptZIslR+A+Y
/1pehAwQD7stvmYAt9QRW5hoOeH8pl0655VmD5sPJsZx/7gs+qvGvk95YSQa+gNz
JrbFZan+UbDYsaGboail4RTV8XPhvXvnGHH9Dw0jH2yxavWXoUe5QlUd33AnGeEC
LHCWgvMSDgHTmLvVjswBq5VCdx81+/Zl+AorQ17Bg/EcOEC4Ae0oDhVSv4YXfOVQ
Xg2XQYBnnawWB+lXxa2fiwH2HdoyVJWyGHFqRRkO94yPz90qOcbyRdBV/SSD5Rdx
gNcll8GG+Fs1buhg2Q1PTgZNjLepGf5oLLelzHks1Ov0sd81wW0zu980t07iCmmc
iszDXCllgqznzSTXtoP6fFVd4fOX8BgeoxmxVaEs2sSEHCcy2iYIpz1+uhE7UlYf
uBYZt5yYRLVjQI96I/9YVN1BBAi2Vod1FIpjTYKcJEAYK6tfEXFQ6CDVUI2Q6K1K
8rYo72SS1lXEq+OY9R0RNMnZMd4cc2BnX9EwXpEVc3NJPVAcx8zRlJJtZhICm4wP
7/kKf9Evw2wKWm2izywFif1uQwVmpuY10UXF3Ul+AEKvBreCD/T2A5esT3OadhGE
BaGToHegr3y2sJiPu1T3DQaVyozYGUkpqaPKFYIY5l+/IS5HbWVuRknHyGI2bTOb
VkDW9eOwbN94MwaIAIKSqpu5NsiJ5RWCGk5QR3/mAQgaPtTHHI7ZqvUW/837XmQ9
bJlXJRPW2KSz18GKg/CYgZfhRvO7XBr6NxMntzUi3UsQHZ+/ryKqnd1s7giQaDp+
NqTq6izBGM7xIxuDXSTI41gcH7Pib4iYU0eYHFw9vJkO8mVQwJKeCBwaraum3sSf
L21o+QJOtJDTsI0hZZRlJWo/Wqv0jhE3ncXDydl/4Eqx2xQ76Al0te4A2ELUow7y
fT6U04XTSw4kHLZjOwSZZJf1E9zm25fQznn8eujnWQKQq2OSwg0xy2Xe/37WtXYP
7IUlWiSeTIk+NGDe+2wQJY7VxektCpLfJ1wlVx2WoHx7rziF4OVOJBsreNl45Iqb
Ke4zIAb7YsVNEPtkZp2DrDdypiZO3rZnjIc/YKI94tOnmunGFxtlmwOcbJtwpCis
CTKJETnaOvhTzFBcBziWECX5K+QuGW4SqHKRDW6RauSCTyq/7T8+jejF6v2zE3zR
JybGDeVICd+7Pl/EXYQvnlpK8G108PUFMgO0EbP//rxHP9Q3W4us8Mv4M7Gq/Ums
JXryvqx0PsN3cVnFwxNNIq0TgMPqxOC7Zu89LW7qptdZEI/0XgP2fIPvXoyQsQsv
OaA/92BiyJbBjIyT1fKTnQ+K+9nVUopc5H8UBB531QWcvRi6rhTijtH/VbioDKBi
O7l0Jw7Yo9i3eW14skw215eSsVc7nSemSrW82UJfx47BkmQchxpkNpYAOqm31xbZ
eIGiJuQixV8WXa/wMvyga3xZnV/yCVwJJUtYTMAB3SsPxZVIA7Cjbmkncat4amox
fakbGz7UoXdixWFsQcGKUj4vi3rfqZ6lG2gP4FZZFpYI1IAFtyyN/1j7TY8NNP1/
e8pAk8mNvoeeaxkkB1VVrg0SjwIJZ3YopGcESYztJyAe/TyQP5olEhjj5IRooS8z
SR5tZ9ulpBuhU9b7Hw6LOSxAIdH8KKDY1PmHN14FbPOwQIhAiZ80eGcJhbD1t+fK
QpwGLZ7hJnf5T8P3zhnQ8wgWtD7TlWicvnDcaAy06VyTC6XqToeGZH/yv2qRUBfd
CDDdljL0o4/77Dpk/W/4EMukxM/HD7Ritg/5hmfHQt7yOLQswOKlJSqAWsiTOEPY
1m6COi/osy27uTtT2t+Vt0tOMhdhq+m63KKY86ZPdzexh3qGlucRe/gtyBR9t/Ry
shlk6w8CAcTCXvrHNJxAoOzL597IJaUE8VZ30C2PeG/9eoAVB8QsupTejitoMyQK
p1Rt14EWiLmfLb4zvH/fsj6j3iIib1JyHoNrntrg64IgIYlRIwQaQwavOnX6yCIf
HxRKXDBGRMn/BlSS9dFlFLGeBdkfdhhtXol2aLtzS63FFD26fIJrNCxkgsUaugDb
i2PFxRdk93WVhGjuAWT4Dfw0xyxTKNgowdplVyJEX1cwzcs6sU6l+iMBhq0dOUbN
2j+KwjQwEO/c0GBI6frdOrHF5meJr237sMnP66nosoF6+JYUZZwbK6ZaSrTcuPbK
Oh6adlvpzfqwpNSSaheoCwhVuDaYUZQHZSq7faTW578GEufq4M7RS2D9VnPzmDJi
gFXsX+xwfSvXM3NRjogZYyc3hlSPJin1/hgPaF3+PSW/VDx4kmd3Stb2fmAyefom
T/cdybMcceWERoXZBbtPptxvL38p7jKJi3Yl0RuXGo4Hb1uZ5f4ys7XKssPWheCU
OvexMotlk2rneyV17iThvaiTV+XPRkB3T6qJEJT9QhD+u9/3C+ocL2jlZfd+cSUi
oyTcaRSGEzr/orO2ZKqMp992o9hoP5cyXpF807FoT3GUl0OipEvz5TOojqb2hOGO
ixUnit6e+wgz6qIf9QyGTYwjG9N31RWJHsH9+6qSImIhS8a6hZiETvDaNWzuAK7P
Jj3/rsvBbKX4HOOo9CcABMdXekyclMzqjglDT4XH+ykCstnVX6+Q38PgvaW4vydc
OeTHPkZWufKahFol5x3+o+SViEe7Dcm5NNLGaonoCXGvcsya5t7TyBdPbRDXVOaN
b83TbRud5rSpIptqdQreuhDCoikBK8kXcKvM4x6Ffqozq3JlGSZed3kxYuDWbXM0
3I5IRV2SfssBw5Col6DfuWsOA12mQWVybip4QKIP5JQsNz6k6EJUCYbF32FumRLi
2ARUlrxgiQVsvjJ3/OHHZHvCWzm9ocnKG4SZp9eBxcRAY1Ag70sQUC5cNIonSc/P
FB+pq42Ryr1vmTrGeerrHZOma3907rvzBfyIid4PEYo/fHlO5LlsVBZ8NB+7eXpr
7QiWvBDDEOigwfc2eXbKugRjjrtheClCqovZIhdtYXleRxf8utef5p3nAtZRRhld
bBMNeoZ5pKrjqJncEKDy1KG0T1KCvmF/IJI3C8GvE5pbJTlh6RDE2KMyfgBIsbGz
n3cjNX3ZS/ES94sBMjc1EollUsUAsL9DEhOHBMgZ4rVlZN8OgABIX9ctficSmSM2
o1d6MT5MqlpF40sRcmbyfP3aiS3j6C+NtiN6FF8fzM0tpQnwRo8+nG+fpAf5bN/w
qA5/oO4qVJ/xFWKRBSVfbdM3lfysEpQqOdKzc+f369Iglcn03fN/8LrnDzRneiys
PkXQ1bfkFmQE4wqNgGm+TN8XHYS7E9ohqFztHLSS5Dx4SZUU65Va72i/4sIN/FQo
R/jb2EL8gKHUVPaU2A2RE/Q5JXnOnNM9qXTY/OSOrnhBl6PXS/1Qopb438w+g6Pe
E5Rbr6nMchAiViGeyxhe0tjqIiia21Hlg1GXeoPoT9QAmJrp4EGybviQYIu1nrQo
MriFye0tBm0kld+ZcUbbtk7kGHzo525Ci1QvtOUlmUoSP/ZbDWnPm09ZvY3X7eFq
B8krMSYfgzlXu5a5BmWofomUfpTcJwVYjUwQ9GrEKVTJrpwWbHpl1eKU88a8cl5E
1uEpORL1hcK8+NjIXpxJ+Upl1xgQNd++j+QzZudOoMu+w8MMcyYrLzuwGoyWnQbq
K5h5WmSmjvEzrnyd+5t5bhDP3E7Uk6DjDRmyMdSml3/1WREmKX+GaPEGgCUBYeQj
ktXuxddt5N8/P91dRQHSCUHHD+GRenC2zIZpnzVBD3nrac3stRnTHGkdbrMlj0g8
W4sFBPjnszmVyhfch2dyxik5T5SyuElHwzLaC3cCqjwBNMN2nl3URDWU7KwcKA1s
Q6MXN5u6EDONv3oxTMy7RVWxAXV6r/r3SzmghIWQjnV1Ou4n2Wi2HagANNiY3n+F
RgzmWo8b2HwYAGjulVXVmLjeWnx2aXptxrf0m/KbuDo35akA3YGyMC1UdLpY6kFA
rP4AQGfzhGDTE5KwqWbJn3F9MeVNQ3ZINHyDuYsScRijF7swtD4UyBULSx6Bg+UN
Y1rPtTRvtfBZLkVltp5+a0H8BEFsTxpj9DXIbl6hXpmmEC3ZhSJihgTLEgo4/kIq
lIGZ+MaB/osz5Iu+B+RgcvwKIHd1eFl/ClCvHBfeFMej4JHFM+aldvyB01ww6OvQ
IAii99qTipz3cCBjXWLL+ceDxGZP7BZuY3Rk3H26TqAWJspsqnaXoSZxRLqpdsI7
Ws4+cqkI354UwF7Bwu0Qdb8ONPhcz+msDwLgpOj6vX/MNswIVJfdnK1MXIkPfGxe
taWi5R96s4IK6nNESJOYmtMgSYsDwNUGm5P3cEBv6f5HRT/udF8DUlh0h1PAK1gw
APHyaZRq7pVWQawbmwu8Ip4EwZ5Cn0K5Nm7ktWEPdt10Saf0LsDbuQX8TCotnNB6
9TMg9ri1mBT5YPlYdrRrRncDvjb9lnUSQt48dIBsDXbtm/hMkbxrjov7+oIkkSWw
EA2AO3MdTtB37vaAOwtzDz+pVbvxE+97ID3zvmXa3BTlAQZOepsnYH8lgYf4znsM
h6O6c26lrPtdp59yEcucfgdoANwPmC8Hs+czoFomLjZrxk1xXaCvCE+zZp/usjFc
M7qg96KWPFaDSZ8rs4VZVVMByqyUOrOCCIYiYmPEz1WiCoPzXZCa1SQpxCK5NHAW
oKlRVyZEblmV0LIWyDPKfEjREVa2bfAe07J8n+SlqeogkgWnjz5S8ReXMk2/zj8K
+PepVelubV+8hfPFIfs/HyGxLjYIuCsFQcIkZGbu7maAsxckW6uz3enyONUB+cty
pobHP2RNmjXwNWwpcSo0uD0bRKqHvRFK0GlpbVtcHQ/USDbr+XEtoLVlS+y7y5VU
dbAYOHCosm2a0H5aktwjp6FZ6meGRLeUR/CIU0OXhmgAsac0wi3Q+a/UcFix8HQF
yoMAfPWHZXg/ipzFuKJ8Q86ZPb40HEInvzXMeSHBUe+QxuSiv7cl5MsVZ6U5CgkQ
mjB0xk8yWnhWLQ8xQODSRe6mF1cuORA+cluRS+m6udoKRtO6rCF8Izupsz0dROIB
zGYMD681nfCjVIINimGQ7axA3ZRk39Z5EpA3GC15NlI2AjFHOSvcmp0JFi5y5xqa
eFK+L6IGPhxcK3e9PJf0y0x3bDkBfRoEFpBgKdOhCYYx6FAkIQutcnwCtSk81j00
4/vZpT5c0SbFt6+gcIAZ//6azM1tVJA30ExCMlNsR46yGfDMVbLdWQVlq0heB6UI
3WNT6vyQ/MWTqfGNs/ce58GPIJP8OxAslmQjo40CpFnmoZqKyBV1nqjah2daL8Zo
pJVE87xdGf+aUozPHQGBRDjUOaSakZcpK96fwPXLIBndmfL2SQWt0AumcipwUkks
C9CKklPvSbSe5/6rL2RZ0/S7tSbBCBrNJUpfiu197DtMl0qvbd9rEGyrIlHQz4Md
2YXldYfkQcGwyLhYh8sjyXQ7wNA2xBmbw6JSUqULQu+GtCHdXEyV7o8fTRJJeV1R
Q50YGzQ7usORy6N16nnlc8jbP5NL7AwvNOhigpyVfUU0KOLNHCGO1bDwooC8eWR2
Co1GuI8Z6Y4MfNyP0RpJTIt+kKoUDPzHTu+zXgGf8WPQUuPDuF+IvOpcEWdd0Ch8
8bM7T/RXJ4XloFqz21+IV9B2wkzuCqube2AfUYx9f0DSQjDrMAJ50A+Iu1T/kb2M
gBjdoS0BM/w6LaW5yWD1zE52Z/xr3BeGf6o8CdXM0PJsb2n923bKyVt+BuFuZDuN
TPJj/lIqTg6hfQKYh7UXTDEa23rOYk7H1BDAmhjHc/ev1MrozTO77dYc/EztvYap
D7nqJZLlY13OmudUKu3+/rLQsznRv24YQF26N0Wc8U+Z5Sj0vqn2rNj0ZuIBdpHE
uQnQow8e9OJLakBK8hNE3CGcm6pRwhal9AB8SP79Lb50PU7VOpkWZxVZmmn4NbNu
jzk3DbYyBlYD3mO7XiUG+aX+7Mx0qTyOZd6RfUkDMeI8SpOqLRWWBq+P852pBfwh
dnQpU80TsOUJ6QK9rWtAIHdi0T26bXTZrWnK3gPyqneXBuEpBA10hOzX7EHMgL8p
Q0r96UvJYdPoOUiczL6A6UT5+pRa5LLSrZqE1UzurgYNzmXmTdVrJS4Lrq3Zv+lk
6wOQTNVYYkfqOH/ZgrCfNsqSWZA7vjgh3Q/BlgnumY+y4hN2eVnOAve2J+UbXoOd
cShjsUP7Ni2ddjE9NjzJLrcby0GPD8CNyXEqaqj0kit+1zX/i5GaPQdI/vjqgxkA
8LENNmAw/wXmWKgiMOPPTf5TtDHiyffKiZ4/I3F6g3LIe0cD0wyVgmWpOsLrycGk
A8VCkbp2kmXR9Qo9N32mBqKMvAFBssqKdbh1dNcxfPM7us8XPVnha5wjPOv6H4Y7
dQuRbWRIE4l/ZNK7IukWGqRqua5hwviUarrtE8NLijyrQBULn61KDXZ3soNyOAwY
yuEN/q+A0KdjVxV4K9vN0eSVa2/fX2MzWBvW0WSaE6yK4NV5dBClruMY+vk8/bjR
z15XL9XOfN19KJVNxyQ2Ui/ch6L6pDXzyXcnWdQOImD6N2pk3ukn57PKjCTKe/P5
+pQS+HkM4WoDp66g+HE7UGpUg/5huXcCeyMxbHafSPUXdacJSDX8H+dAA4elNvR2
DrPI/Bdgh10TnIYopYI6wqPFDcHb4w8Kd+8y8WW92ZpJqx/Fz6DsunBrwnp7XA/U
Zg2iY1VguIctgmrN88XMu7/9GfOqwoTxEc53Qou/nD8r0j+D0q0Dlzpzl5fpjcWn
d9lVbpwjZ0SJWjjcoUA9QVr83BEMpE4TYhaJGTt+dBQ5eS3UhZ1mRfGYjJOQ8Huo
gayXIqc8bQ1Tpv/IVAF3n4L1ceehrijlM5lYwS3drEqwQQAhsvDYHKOspY89c1wt
0MgVkoi9aJKE43q1eXbuOQkOEmmWT9KFbWud/naIdd6SXOqzF/wLSjonD+dRBUKY
a7CyjAU3q4CUjhWueq0Ar0z4YGEMAMhKamlpC4chPUj49k3LIZ/SY2s2GEf967LT
gaTpoic5KJ5ogGpZC3lT4UggfhaueYEM53xT1HdhSE2GzlOtlSxvNYqFF7hREEib
3bOLsRO6j1jJseOpEaAmLQJ19OVV/8DQbqgz2piyRJSiMmF58QFNaD6DNF6e/Jtk
09UdiyDFZir4JVIJRA3nn2Aiu/iG5uFikvJL9u1eBqxc+P0ByIRgN3dVzGCXHBiZ
H4NJCdlUDUTzaJ8iUCwJajVD9ntdsDvYUPYqJ6Sfri89OqGguL7/00A5tF+0veUX
/BCYsLr5+lZtFNjdgKXTjgv2TsZNRCI9TYNSBnJwQ62H9a2gXT8zBGmZCNsk9kCb
LqTMx2wIKL0anB8C8vw/Ot8jItTfRYy54kCt9kaCPnGNBCy5F+A1Uq8GfMbGqVO3
1WQ0qcNySx8FA56uFEN+NWAApgEl+WJlX0QKoDkFwHjZEY3r2E5fy8cbNdYMm8WO
orhgTBSB2JINvKhquktKwqHebqHyb1FyHh78EqHvCeWuAdW1rVt5D9wIYF2BTIsJ
9oj86N82yImXUE+tGA+LtG878svAgcHCmKNUIp5J7i8h/sDDjM4aKTLY7IUDxuHp
sRaZgIOMG0i/WtBtg8ZIzQ2ic4SMve+RzgPM2oy2cCLChTpWonioRPVcLdx3FQeJ
ACZETSkJ/MMgKIDlIu3UerFqBdhgYnmBoX7PPPkH63ZwKbYXz75iepC07g2DirDh
84OI8dbh3y6zPysQTWg0Zi1aRad9+nSDnrSFk6g0rgcskaFjdP/ZJBvt0neGbTVD
G73lWzcc8M6Ft3HNbvzJGnGU40p0H+rVZ1aOMUrw1zjl0a9i4ahO5TrYzwgn3lRR
5gytWipaWq7J0S+JtDMSdKqnWWf26QqpLIg1gmlPuOwv0OZXLDG9CaA7ombjaMYY
WmiMtMa3aH8vvJrj0xgvRCGWJszFJEQCgROoR1QgziFuVAol/LQNT/aD31o39Pep
P4F5R9N8NLEK7rEMx0HFZVPIB1iuBRdI2A3OMnt0IQmg1nhOhU/vv1IOJDvPsrPo
6us5lc0SDaZh1VXTr/0Wix1owmgNuwf02zw9xF5DWRJy/+LxSfZJjTflkc0apM9b
97mWc/YmdbVsSIU0EJ4wzxl5nSQNE1S1clHBgoS6Ck/HxPxW+wcIlZh9OOhcJXT4
BFJ2Q2vmtm+ZE46HH7HffdRr0FEL75YKIQxH/748KYrW7Qa4TJnrrDQG6fOw5l6q
7x/lqbsjw3niq7ZzrjkYJ1oU2urb5r6uQZ2R/nApGxpkczg+NsQ5FS0whlUhM4Yd
hzqjMq2KqjeVed/b/fWQvwxr3vmPNe9mjY6FbmbuZvCotLzWkZlgaQTvtJBM9nY2
Q5DnqchZAdIpdL4eYhRcIQbreuyHsf7SyuVFFr+Teix1glf4sST1jW8uPKBXt0aH
QC+xaGi69kT7pstNy3nRRxObL7yHwJtk0MvewMwuiYgVcQi6fEZBGtCDxuezKiV3
A6nuK6dPGevYoVXvCnwWa5ijrksKapScWsMtDnr+E6cCICIzDvTkPeA+eTq87gJo
xiO+Pnv3rujUcVj6701uqGDtmUPHJjFp+D93eeV9m45KD6194/U41gm0ALMkY1sc
kP4ef313E773wXc79Ha6JKlM06rTwWy49I9vIfIRXH5r10GtiJEasDYa4DWif/w9
6sU3razypBJvlKUyKOFgSiSIyD99kMfcH1rER8jIua1i2HSYzQxRivbJ42PZsycN
B/C/0zluQQZUW/9SotSQN4ouQxMOveL3cahOAdzUWOMYhyNtQgN9BviPHLZZroFV
VH3psCpNz0YRdVvxgByS3jQI86cUudzMGN/CuAPtYy4RD/s6i5o2U4lX4JI60p3r
t0vhpPZh3olUwBmFJ8FpkYdwOns5+7LNS2HE1SDlU9QuBDxcUJsJzXVVZneL1/VU
ZgD/ZUackc60k4Co38LH0W4C/m60HH9beVm1LDnqc39dWidWETOkeNii5R/u/EFk
Jwb9dUeuxH4JMO/YtrmyuL5v3jOiK8+OwJuHC91eTmkjLV9p3CSxA3iKD2pltV2T
LT/ULKpQDRPe3TRSqgIE5jFJy92spEYak1KaqzV+6A1B9XHDVVVWE+JZ+ODPMraM
LZXkFPFTPRFSZY+XjqKmFUaLZbWbU+H+LRXUMkytH4BOlr1mJPZsW7T3MjWXOkil
uAU14svzimR2CO+xwLLcae6r4InsaI+u2BCpviNYOB1HSX5odkJ5oAYuv95ZcJfM
iYgxsR32S50YzRi8VHo4z+B5MCMfEZZDOjtFZ5zCBTrK4VlaRBmmmr0k4CLxOyW1
zVyE81FCaF30yD2hrWKvvYYaHnd5302gzdX6zpev/m1jYqy1jCe5R5vEqJtdJ+KT
vp4CeW3iI4o4mQGGWcZKBosb4Hg7kxJ1F7WlxcVF4IbRWtPolhqy2Fd0lhIauB/0
T7Ldfy45eK2XnWwj12n+7fk3qAP8Zmc+aaBb9NU/Ot2ONr3qqggb64P2vTyCPoEJ
pfx/DS+2aRAHFCuSXl4jbe7rBfWHk871lohzJtFM9r6+WgcGRmk69asbV/UZK8Is
C7LL3/13JyMa+VJW3L6vOyNqneWyhF8X1VRAI5SZBT9UCnW5Rc0vo8RIa1qpk/8Y
7AE70jpnBr2ecaCUU+VIPa7ZrmIgXDr9uUk/sIze684zgwOaob9xcVtmjUgXyIFj
bzXfkEYkkxQWQF/Ew4QW2HNdIuRE52qo99d76vXBjJj0XHxz5NO/Y+N/TDn2rQjr
oCjRoWxXzqPxZQ7GHxFxUTDQQyX//aBrnr1+VqKliASRzbowLqGeZ80SxfyUkTnj
cNqMt3R4T4jcyo1cu57SdnsB0/xwOBP0+LoyvfQqQN+pwVyoJsG41a/pwEK1wnlz
udyKmNa+TLdn9TNjQ7o651wpA1ILxKR3v1DNEK27T1WqqOQuW8I/AQp6f1MxTsR9
pO72HdWKKI1kbydAHvKCtdnnCp7K1Y7t7buRlroN8S0RUamRhTfn5PGzWmQSFPjs
WvFivZkeHdrGg+PZJJiG2YS1PHF9QlS5Dg7QUJ2eFjCIOp8ph07lMOJc6a/leobr
ptegPVV3uVUGGPdlodsrJa9BkQ5N6DUsZcgnYdKU8Q1+fcNN6FO5PSKYf1F1ciGW
BRuMxsXEUYI7Ku9TGBqAsJ8+KhMFC+5TO0UQ+wvQsfIZS78UQfaiVz7B+mN3lEbb
4JVHvBh+oR0BdNFS1FrxMAE+WPe/eM884bTA7faHeI5mAvKXlv0BqxcFkDfxvLti
lr2vf7/B8yniGPfv3UVcYIlmDSAB9wuQxrLaN/cZFDtCGxgeZGHZDpTcsVFtHTyg
Yr/GiEIKNuOWgipbukb/tpflPXJtmJPlCMaYSdMyEXdEa6ZC8MPggTWMthel5yBc
d+4BpUMTW/5KghfdUrkDx/3y8eZwdq+Si4nvda9LL3SZoeA7BP3okFrW5Zucozox
wO03SwhniwRFM5hAhXLzggFPR64XWOUIxGmr6VbzTXdQ/+tm736gEp6R/grPIkE4
X8sQWBBW/YKDzHZHymAsRLI+jsj96RuF77ewtbwrvODJEDm0S1IrlqPT/b6OLSMW
cKqIH4bxdF1Cmbxn1JTVWK71YkwOYVLBR5vu9IiDemaaJLPzAelteEKEVrAsVih5
Wqv0rwmnLKsNUToUQrO5n0AGwjwPCiwxNc2TBLUUTZjvT7ZtGVC2QZ3O8z4KEZl2
h7Uljun2XqGBfGP2MDsBKf4uptjvuuKYrmi7qmXfFZV401exRsFhnjbRiunq/sHC
51VZyCGSuyn51bKLenfVn/5f2LqgCOsQKTUe37wG/Zwg6uNo1Qa/2OP6Sz1eOonY
zYn3bfMQJlA3JkGnZ2OQY8Apt1SK8MQf0Bja7k0OdVaHf40BaCXM00pcGjbQwi3M
MpBEy0yiu9x7G8aYB/3i5I5qYYQGdEw6gbcl76g34yCpVhb9EMOZBV/dFNVgd6w4
321/y+ZOxPgASGWRCJKLA/tqHJwNZmKnBkCFiOtMn+3NMta1L5Njn2rSOBRyXmtp
EC0g5EVeshfvZ7JfuCs3HJcekt+qEWjliXGdpTvC3BVx0tkagHHUPd6expwS6jwk
Mf1eCQZbqaSfv6thxHzA1hl+FTb+SeK/4LLE4zy0yhTR6ZSwOCAvCho9/fIXsYhd
CF0oYR9bKHiCAI71nQLV6m6bLkLd2QnOnolShFfJJISDF4VHO+i7/n4gzOOb2xSo
jqEqmsGU1CLFxzdl6Drgj3IdU+2iaG2A5nI+6ZRS/1zE0YHIjqsySY2qT4ITFG3t
D1nSw5PBthmEaQUvyaxfbgRJtzuxnIwkUAPa9+5xZ9RUI/512WeRORcr9AYpz5aS
UHYSaLcM+v/VxtVdWiIrSkZZM8ZdYDHUXhGq7ASU3k4yQ+v6DV39yBUB4rBXTIsA
+Sxej7rG2N7XVZdbqPiP4Y8jI5l491XJxj7G2QTzgTufXuj5LiUf75yLTYc5fFUX
MmJpRYZIZHvTV0dc5mKsjuY3c5ZQ1+L1sRbFicxb0oYuO3EIuvuAAR648h0qy4nA
hOFUc9lZQdfgC89dKLxeWUKT8n1VzShD60hW1wUuA4dyQ5S7sKx7/K2WGFASQF8O
EjG4m2qp1xqtDx39gRsohf3byqOvUcuLct3bIuh66XucxDIXAm19ClM5yMG+2by6
yuJ4XRbon7C8i4dTaUPvf5AzB9EAPse8T1eaJlQ7jBe0BP7gEbOeHUxUUCnLZCt6
Y4G88PUZ+YCD2rq3DHCJJAo3cX2/wi9Z2uZUM4rCdkAXv+VcPw7RNxkB+RAO/tKQ
lpymlNRtC7TNrjQg+2jl0VOHrUk1f9ho8pE34eGC3NcFKs/O0dLxRpSv0iGt0X+k
y9OGHfKwyBqCRdPS4JdemuqDtdDmWB7e0syx0Zdrq/0PuKdjCSq56SLBWSPB/Se0
5l3FnJALREXTJ2tcAUCgM9E574gXs2yQDM8mabeSe5WywuckN2zzMWqCNSA0atiP
06r0a5qRkGL1bzzqGp3wCJpepwzeky0XCiAOQ9OR+kngIU2Ylcb5UbMAkWsHNgvf
tA5pOdIuo5F0ZdrUbYhO8n2MCMyCXnJyAVZkKuexfJm0B+XQdgrZVXu3DewnC/Gj
BIC10sWslUEznpUYoZYfZcVchdYJ1QnBcXwZqt3Wy6v6Xa20XSFzfRIJ7QVnKivg
Ueafk4Vy3KV+N3KMYsbaakHjdgnyBm6+yzo7LddMs3G8PKVRoPvzCBc/25dDapxm
+IbAkdUZrlQUCcC4NHK1RMUSxL1eMoZYXr1XXmxI+HJaJGNgCLAb7ZtYByO5bp3z
SHSLIDHK1fdmb+htMSBRt9X3yX69jhICAn9U386E6IknHQVUb7ebaVn51QDgNq0m
LqH0MiatZzoR+AJVr9mfH0fR+iOWXUJQ+QWV5IFerwlzEct5N3LVX1ZNnE1eb4zs
AKxxnXqLex1R1MvANaF8RN++DshZ3LLvNO2m/haqxg0xEC65rFSbNfDruFJ0Kuf9
FMhCxFzq9aW4bftMh451WZ8eT2CqWjHukowLgKQEOA1hxogeD0qbsrEV7hmLpC6M
sJxmLI9wempDUlXvupUneSzaoGlZj4uyPjHfS5vxHOx92GkBAMADdZY/yKGFPjm7
3lWQ34IuvKX0nKaH+RfANNa5Zcc+XU/MjLSkrTlrvvY0BhPd3y8Wnrl0dD7uHIHu
sWpeWfPqKm8Ad4Kl1KeTWELg6Sv03T0BY5fWk4oDbZ/F3Bz1URDybE2ucsPeHgs/
OmPuGDH+4pREcSkFD17vEzbeLCqa4ZA88p3Qacu87R2TcyQ1Tisu3haA75wrD1Uw
/yldng2XA2CicO54Iuqe7yqEb617pvt9vX92FUcC1+Z8pqwojPtzGQoywMnOBN3l
KaepldWKwSwdrrj+zapW1fUktf7gi/zhBrwuV/dpOSVs7ZPdjYsksB0dnd1lJOZf
lypDThzaaPKxXxIPEP6A3GEs/aYhU6+oY5U7qlk9dUkZeO5zyqiTyhgPdnJDIlaJ
Kx664P0QLfowY1F0muR9oQQ2/Z/Wvf9bO9oNetGIgNj5w4+CCy0vkPaSt0iw/0XO
CWHbY7V7UaF7a/sToCqoVXEO5sOHo1L1XTWgMZuPteQtUVdegJrshOiVtrlD338t
LVqeXtJ7Ece//3ZgAMbCfVG8H8E8txBW/KHj7vKgDNyQDrWKFe5cVTj3pctkk9Er
qdC4JsavP5FhwfO4IPYOwxrQ0FG1buDMJ2Xm1RJOfGUud4XlXkJAEGFm+7oUNacN
+Y2klV3RF/E9kk5lCWoJ1uI0eJTYFADUKpjRI7EQYIYKg7SAsysk/O7hwPR4mNyy
CbYeraLUV/mx89P+H6gIhIAjAjKA7pVnhjxoAVO7G1WWR1ykDOu1Noflqp8Pwnj4
2/dWlZqLj0rwlCyOXmC7yCwDQ3HrOjsqvVJ5dCMiuomrbHvWRjYxfw89sAsiWgj4
FebZCfJgb35D5vW/AbPqqASaL3IHJAC6lHz5QO6zW+vHTShg7BkVeryiCvo1AI9k
Yx2J9f8Ndy65JlRkJFbQYXOr/JxpxOd/Z1eMqrn8Lb3NK2o/UDI0YwJ5/paaXEym
Dx/lXEersF7qyezcOIEto/ZoEGBQbs5FyjEgz17QJ5+jHdAoSGNZff1lrIspquVQ
52WMM/EcAtpthekzdYtEivbxyAY5n9PYAd5Z7m9zlLiTeFGqdCzA+cIQOFSL45BA
+uXiBFlW8hIgTiWIdVeq9jXKG5WSzx5ZtZrlh5p7KsB/9eIbmtZGOypEEVD5AJT6
iArM+Fzv+kF/8tZWNRdlMJFfZ7yLRAli9pG0ejk7kqTswyxa7IwN3c+tkjXIzokI
k9oGeW6R5Qn34I4xvN62GCB/kvJ0yaVMWVBcKpbnidGqYpmBDsmHUvYZ6vARzRk1
EipPaKMUvhI9/9gI6iOz4GDRP1UHiJNjmUVwR80SJSaETAQOmFVcPazUqUMa6GD7
pz6Lpx1Y31kFwLWlfzBh5WzOIZV02NcAqjeikVUOAa9220ka+Q77xQrSea0qjiOc
9TqN82TZ8qScW1YUhjJMXTu+cNGGPjnjoYx387+IA/shHv15qo3VIvLoP+1Iik/9
9FDGzgY0yoVSko0d3arJiTwf2ZEAtHTPplwmIiNBNBXHAtyqPMM4SFU4jYan6EWG
focLe6t7bdG/O4kchdARDX3bVWwyauDrHXKy4ffNKmFUyx5kMTyoJCg/YbhKyBzp
CsA86PVNCGcBe63nv76IUuVVebvWZtDj3pzBA0ITbUsD1quIytNcTi6zb4Ctkn/u
rrimGjPUlFLaJznHH+aYM2RbYi8d7Oy4Len6tvS4+fg+WSM013qWXcriSxYqh6s8
1g8c73ecU/xYUSLUHVpmnUdLze/+FeeMQLUyTUSeFoHj+aKwfa2+opNM6bXj3KL0
i7Wqbkx8My9EJLLYgSkWuXC2wA9AUEE3PKsplGPMKG3UhMuVpxSwHzAWuI8c5IUp
gfr6xYpEQk+qYu/2VoRJG5WiRfOzZ8IAKqaYkKuixpsFBYcu/OA/0gTwFJLyyQuG
Z660wfRCzArt6lj3fnTDU79w2gz9t6f98rhDXWVy9bKbO+cod+R/V7SfFycTaHAL
FfhWyIIi/A69Drxx6XyVN5QI70rI2xkgASAnIej23WAyyu0x144CSO7nvuJNTjF0
LWNrq1oCtlyeTVYRLBRkJslEXgpklS4nan8xNtEayD9zJeCrAgd4pKtAsASz4K+1
yKOlMIVE5Cj75DkaAtnpEb2IpJ8SX2WdIuQZW82BqjxSo6ie1dYe6xayaVNOhjyO
1DQRsf6bdyUlCLtDvSCsAOumCY6GjoJ6ypGZynQI7XJ9swgFQzbygC1Ba7j2gDk3
gF/10vkuzSI2DtV9OFGbLlr2kDpyG1Owx5unEUdXrwtpW4Po6+qM9+CzfBgpP4EU
Bdd1w4ovGgqnybGdAv6p/jpaGoETuCU7TyWcAHXW0Ohs0UzMjDh6jEpo10IWqVUP
IktiXgS1onkyzSWco0VjwcMkN3Zi1sSd1EObaC6vxDrf8ni8d08b1Q3DAMbYJS43
9GpnaBh37BYpA5KlWaKiMJ2GMMciLXRRez2C4dfh1LR5qW3wt12SH6DgxCtptHpK
C2ElsqUkl0iYks3o4r+Dx671YGKbM7QWFTwftAJzbTcC3Q0AMpyh6QOryl1hEhzW
oXttBMgnoUrYT/Zs8pXld8HepPX9m08B4gpNyu3blquHrGbd2DdngqH+IubpDC/J
2uR7cLacTFDXcUCXNCfeCZOOQjNTxmfvsEca+JwdzBTV12V/WxxRfcfGGLj84ZCM
rK0CCLcC8SOChuPQzdGD8UaQoOqpRtYBOh4XZCr7EuMoJFtZYHTASk5g3BGuwtOg
Jow9IetsbVnDrW9WCKX2pZ885bMfZ99c47Hrhl/iHNV7eWoSlgIWV/1/TTCEVntt
XD2qQHNpPaIJd+2xrk4rfD+d8YEOwGf5lAiJOkNkbc/qkYjcnBuOhr2JoNA35xVv
sKR6/v+e2Cvcni+8gDbxYALL19dt+3ChNVqSNgKBcn3UFHLy4xhT41Za8dLzr7EH
Qa9YM8u5041IYjfYIuPWpw/i7LWiGVGwXIoI2EC9AfHUlg00tmqnO3vvNOcIvgWa
F5I22fB5uoefNp6cMmRYWxt0YWTkdKUtI9qjLDpk43RTir7Sqbq63NCn3jXj9aaI
naLVYTMN6w2bV+4mjf5/vh8kUNjLBpqo27UgRm5RL1lT5PbR7g0fWkxeXEsf5mZp
cCWC0C7qfamsfv7Mh+kN9PkckSW459q32AhvcnCnE/0K2n8tSs2XyrpaOqyuqy0y
TgcGEvb5OBsvkyN7hOJG9eXOZNLS2KEXycFI2efTYnNiH+YZzIWhZRqfd7tAK5r4
r8S3liC21urL2nhB9iCOlehz2z6EaKDtKvcUfCBwA16mJOu3f1Cq9qcQD2X6dkrM
27WlNhtBO5/KXco+eieKRJMTpVryUELXlJ+nM15S7nEtZ+lSD/ko+2Hc8Usg3sSk
PMlDsEv0+24pDxt/Fj5CIYGJe/CeXhcG7xjXGS5/D0SF4qLtSiSZm2MPb6SpoEE9
a0TWrPhqWTjGp0tRj2eYeK+Fjk20Oyk7bL0w1JB/QLBRoI26pdbVxULCl6bY7Xaa
L0oDLb1Ibi6v1KwVpBc6CmEKovODeVCYtFqLuP26viNX7g3phckbG2ICzmL4F0zo
tIiNM1cMDIQdA+w2GLfL4F0l85jb0X11rWjVNNCW4nNCg3xEW1qmeThOLJe7rKMP
j7AW1Ptj5AI8oEZpj4WDlLD7zNlnhdOOHB7hlQls1FfZkEMPFkchvpDTe7GVhRJ0
GEu4qHZMuDHnPtg+XSHXFzMwheITCvGn7kCEDIYezpKUysZgHymAdIDu5aposUh9
VJaH9cIZHsA14fE0zDXJMGOi1PEFxpDUP3dKxRG3zp8Od4UNSq39XlfAW7NT1hqI
HDGmR1p0ULQiMg6wiIiWOwpdFgIe8u0hvbfOIeUmecOZryzuO45vAx/Y5BrieE8E
tBUHO1qoWkqxmyIeIXD1jfklirJPf58LjQ3RVVDWwoglcKDbcKDcuukuCUvB4cUt
vXrEB/2C3B3RSYFpYr6cVhuT86u2LUfkn5mAIfrTWbh3oNuse996+UMBrO261NNh
u8zU8vcjk8Jp2yv6SbDDJcw6eBXVPQdHbs/m5kYpKP4A0C6C8QKfEwz0vRFlxF9/
dz8M1dnSnrNybDYC1NJQDZxig8Mrb6qICF9BQwpcNhuz35999Zl6CgIqyBFmjTjp
8w0AFgS25Ep3Kn0OxCno/KKpOnPgTNYOXFewXvMyF5dE+XttVq4/J1RlWstbUAm0
O4YVR08FU9eFR6vQ/vcj5rT+UWjVzQOF8wWwoxzPMpLFILGq6BV2//beejYiaGIj
44VedHrnyNN1dsZqp3f6vLz0OMdt3JQBHfVxkOpdibomOJUemojnw66wjICKJsZK
8PX1GFdVp99W0/5X1nXYGG9pUBuq9WLMvj5ZWgLK4VBzAFLCGG96+437R75yBwca
2VLeqamLsihQ0cbR8HGj54tmLYuwhiDhmeQMn/xgpOtXqwurWUwuAGnzHAQFEBnJ
ATiY+nIExIkdG9/tE5yyxynDDu92cOCOoK5MfOlgbqA2ChEA4/vtVrSufP9k2gQ+
l74pCAXxIf87F4JVPAtvHtw2D3MZwZk1E9dxK3DTRrbr5U26Mdf8gqIXr5j/vA8e
RbQsg1bmp6WCrSeylqCVlpJR8/cNp0E6gFcodczY8e53Rz5VjKJSpvkBVVjWf7iF
qtJMxjTsCsnQGZ4ALDwQ8rWBnlWtyZtFItyN8a2cWoD2ycavzBUXbE5ptCy1mJxZ
XvbzdsClZrxMyZ5PJ4rCekkvphE9akoZNnPlQxxQyICGiP07faF7Ozf3QIkcDjxX
SAXhMVw7qC0vfD9zX/7D4cLdQB1IrCOhMx9fXyrLflcwafvi9V5SjV5gy5Lw1fte
1+XhtruNG3ZMkV+D+G96n8a78aJl2DAPhPYozavLfHb5kqUC6JFZuUf3ig7LtqwL
a2V1SyB6UrfBs2gjEQvDrWogYn5uTU5H+6BItZkj3XMZcGfspWA68ZGDBi0kCKXF
3LtBm0IK/asmwOw0Iv8rWvaZuYX9KrMSp6l2pWvVAE2CnL1MhZY2yE1eoJCzQ2Up
VBSZBjNrtK16wubHb1BglixL/AF0tio4t1N+o9+zGpCBgsuviOKoATF30h3tx7Iu
ebV9KwJsc1x8/NU44Bx1WS/uAdm4xdCOrZiCgsA1I0C8DNitODoJEi7YgfwG8V1A
/BjP/5FC768P/T9i/lL3OU17xp1LmTWl82jhWLUSVT0Bsxc5PNao2Qp+AfUEsCs/
+Zy/evlOb5PE6NXUGiMkDvV032iapT5Zq+dSV1Syuk/riIedymbc/YtiP/tQ+2t4
7r/rpiTzURTnSdTmLTrO9Mc/13oasXGxkGxFdJ+H6yAlN4t6jonwfd1ykNg+l5hK
dP4W7ZlO2FOKq8pYs3IiK7Sjxx7BX5KE6U6wiexvVjnhO3CPbUgow9DemQ+fKCrs
qTSdy9j19whqFTTtoSqRL5lU7MEvWdzUku7zVly2yJZeVc9RJ+MKY6QDdofvU4QV
g5k6IlpWIoX1s9rPDl5nfTKqeKnUrJZB1nVoy+/uD7kcJk1unSo59qbfYrAW/vMW
qAqwV0fRRwY0d3SKWpGDjGQAWsRYgfiDoX57Ha9scARl9iV5MWBZayBPcGtyOPGD
y3fuM5nu/v5jOkw6nyeHXuoxR4kLUtrOG5bz4YgE3WfOliy7xWAHFISyYS0iHUHW
395Yp+04p499o6p1DvAF33nyI1/Yo0WuCwIKlZegsLwQ9fG/q6/C9FXPi9xQgcR2
VEGdS0+HRjh3h1v1PzVMHj1pN+LZhdZc+fmVZgrmGZw=
`protect end_protected