`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8432 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhBNVMbsl6PTB5/ApNH6uD+AhqaNL18ygQSkbQDCRS3W4
CVzXRtBaoDy3nmUsGcDBT2t7AwhlLSS7iU4xsxoyRksig/Rt9NifAqIffma4sw1m
OjXRX99CypJYH14MzEQ/9vCQ0uEOjdjCo3L2ECLXKexebAI1eihwsm4s+5PAtI7p
GirfoSJnTO6fRJ6Gi/p1GtgQTi/4Q30RVV/I5SETDQz0eR+E+ou1kas5lpoAhEMU
J6PnZj+mpEa+CaPcq+rarmMz5ma9phzreyS7bcJFM/ME2LVJf1EJUddKHw4hoAW+
2nKueBljCMlIJ4NqIKNjhUXTjNUwuZDZG0rKmGIibwLF36MQDPz9peh8Af4f9iTR
3hCitaHkekPCOUTXQnb9PSBmVhnHpHCNadFbD0IJiSv6sZk3IjKtoauRnechKvLp
90swSnyox5HtpkhJFf2sevJjbM54W8VHBm1H20c2jg9wnAtDBkFkk2sjY/Ar7dCe
LDs1R6y1EUHk4HB6vsK1b7zWvs6FSPeQkiNIL4RsKhUoL98jGOexb6X15KXWVE88
PsR2rc5a+0g4VR2EaNQP2l+mrQ18/sjah//gICtXc0dAc0zDlFlVImvUvqMtiF9O
AIT3qzs7ks3aN3aYGR0FSi+yfXSqzmhIXq+94u0QJiDbuNchHer/OHm79HXinomY
fYUsBuVgt39ODO8NRRVSZH5Z6m+8eHQ7sS7Tf7KNIWxkLO8q7Eh3+5oH+TGAoiRa
b17uatyW7lRHPKVG/0nCggiid6gNf6zT52uBe8MXlpZdHYuA0TIQmCHsBxcLpdLv
yrwyFLxqnziXiAyajZfFag4NJfDcVUuqJ+xc9L+PgTKimG20ESKuy6dPsVhDfFof
N1ZHndtxtHzHP6l568sMWA7NTJK076hTnn2ESlENrmAbbUSMIhtOV8VsLNPKxzXf
DqxVqEpkjDb3Fe1E4RVzHQMXUWa+LjtA+0M/16h+YKGAYdNGzgIGaN7CHER62nrT
5a8edLSbzlEDRkzEwJAp73AWOoMoeugGQlkhEhlAJgBpR8bnAfeVLxDN/2+TQo5d
tZI7QaMUm38q35oRlDUn1FUCkGpuK1AuiljdAE1EqTw6qZ5QvRAp+ElhNQ8wUzBr
6mCuzw3Lvg9pWF3Wo1WzN/DpahQ79/IG1aGX1PMFVRd1qwyv787xihT6LrUiWrbJ
mLrq7EzuBsVMS7FqsUDDYySheD9PGA/7HNdz9RvmtCxHo6VuJ74eH9h05FI5M5VZ
mHhX6zsZY6aKqvdIa6h5sAeUkLrzYLOvGTSaG2eNm917sHsOgMLVjUTpFu8Tv2Tw
nuXWgPRHSu0CAsFBoYg1zNiZMn8wEuRcg6Vdn0csOcA6j8tcL/6SBgvgxAew35w1
HKfFVLq2888mylW6idfjTt0Z5Z0wqmFzTJatiqq0YQVFwZ1tRjqGGZ0FP7yNv2BG
rFgqmLz+7DjWHShWodhGznrNdBTZcpNx0CUAriEZcrHSxqpD+xfBxLRTiVoyWqx+
uzn5bksF7GF1EdB+/5luRsFW3I4Vp6hXGTl8lTWI1G6NekjtAwZuua1v6V/tFpC1
s7pOvrl5lQYDA5U/1pFCQvF2tOtgYst9MYzHDI9Bmvaz7If9+34uNV7sP/YLQnHj
SmET4dTXOBKXlBGW/RnlZeg0D3j81Uy0/jrrthHCY2HF2AN2RffmVgrZ+mH7SGhe
NkSF8LLBqyZGhiHZeSE1r6+hulE9GjnYiM8lzz+LsHsdgt+69HL8yE0F7+A3WMuS
CKfdHDbOF1n0yGsVzSVatNjCAbbs1J5raSsAfcb+vVksF27+GmU2z9c3QKEt6xdB
+B+jyACc151ztlUEnXbuZAHTxDLy8oH5N3VJA9GlZgiXcS8Xj2jqGEm6JtAgSfbI
Ni+tA4OLHGFwVHY6p52mTz4wc/5tmhlKmaA16lzKrez0Cd2dk4qpHJN5uCMYlgsK
n/5GondXMRT/OYrOiYHgm4vX1U6icgtSmSIdbrBrf6A+oMKNHLBeOip1Kb2NlTTS
dPr+fzNuofyz2p/4e2x1moX8VqJA2EvEuuVy5PrFhdKpOr6UY2m2IL7tVfxHyJ6U
CpN+vxemaPSoHvLFs1gdtT4FhdV24U7F6UIaeK65wmqGF13e2FLOGEahBNl9ERam
yrXvNe2yw25BgSqlk8zM9qukXTomsfnAQ0Xtaa99Udp3WIecffPHIq94Sdl9i59n
ivPDI1j6hMkgc1C6kjYHtpmWlmLFVwlWCPSgAHegxzvVWWa87eTTOyBYKJqc1VJQ
4FBmlkXlGY2xuXP9lu7vt4c1qS/ahZNIPQTRpWu1C8qUnPZIrypg8UKj4f8eKz7Q
wyh4LN156z+EUAeFgqYinxnHjropLCha3Vow1R7ls0CHefjkUsxnhYIO9Z72PKXJ
Jz5a/BmihHPTgYPuyAv9f1hM+ThOOUwHiGYgNhr88XpQ3HAsa+vmzyq2SZQXeRF1
jyPxtULTFx3yLVjcDKTNNoZRFHO9dvHY0Iz0mKnplBS2wbmXOuhTIozT6BqqLFhh
J9fIVPHMJhaG+oWFyIe9gj9Hbh8DVLVVRy4YjPWnOUXVAZZG8xtoNWsni1e5Fexs
ct15tPEmIKHOUdukBPeK5eIveMo0LpYHbKDwPqVh2Z7bY3ywlIZ9A8lCK/E+/0bY
8Ks1C4Vzn37D2bOstOKqNUwDivayELm8CNeVbTN+y8Lp53gmQagPnoZ00LZ6iko2
3Cw1Rp3d/a5NcCYmy9ha4wjiWERK1dEPdtvFnM0dN+yjPyawZIayQ+m+naOpXEoa
JXgZeHgAsMmyS3EYbjqY8kLGCgSFPD3UDnU+JKUN+njQwO7cbsxMCTjIgInBHY9t
lUglp8bdaCwy9qOW2EoR6L9tbRNI1lDS30Dpq4ssnoYKyQ+V65rnQ37GELmF2Cml
2fXidm+bsFfNaJJX+U3+7ApGxoEDfIG5aHHkuBrwXI2lQSDqCDTLr8o8aGkm1cwk
Mz6CFidLrqfanLNSl0OpBpGR4zBHRl/e/d8Uw9ZJPvxQxreSwpismYAVojmysyej
4eZ8khQy1orvVhfqkqM2+It67wgUWH5vOpyXXF2qcSuJbbX0CmnJmMR5Dg4E18B1
XGxNnqlujUfgfCaifZd2V3dp9GLYtGf3wjwK0uH4r+JolNGFwXXkeqLkANRsK7HQ
dCR5cj8v9RJSU4yTWSI7AsP621ZbJWRfdpWPXugz45yloI7wj7ag2AJ7/3MJ3rvy
cbeoMBc63tMZU/SJkLsUgDhRE5CjRVKJtSquB+TNHtYao9eYTISTpndUHhqVRQyC
VbGdLNAdTOJW179I50yM1XfvN2X//cczaKUqIGJbfMSWlHKzYU+4pbr63IbVJJuw
EhcgvOJWjfv1wj4fDL6xPQTq3Gaei0o2o2p6bxQFTT4i68MtvjGAGI+H0wGwfsrP
6cFscsJxs6mkH61yAMu953X75j6VzIFgfIJRObss1fhfEnd5wtQK3fi49WAaTiWV
o70G5aYDAUH7rSbr39DWBI1EGH9cBx+HzkOGvsct/MlNnZqkKYXVLrMfeuSgz/pV
ed7ye7c1AgKZ31qazYcA8uXO8TjwW/21u7qJ25moVir2vj1p5L64A0NYr5mG+7/+
j1E/X7iLa5AnIpA4G9SB0zDSQ9LaG2YCrjXsnEiUwIQpyXirJcy8W3fZ9HKJ+6x0
Y8vUz0K/KMlXetFqX0tcufpVkpC/ysSYhcLxFhiWSFhMl3YFlID4pBI0IO0gM4Zo
DWsOU+i6YWOMJ+3MFzYOPGv1twIiw0uX8mNjKcWstHJBn5GIcCkz/7bKz2BVDYmD
kFsoyUgTCc0rvzTFGDo4vlO6q+KlC5UJkdCBRkyAyn6eMIrV+pUpedHoVRckvP9i
0swhAB53vb4bxxy7elGLUxh+yL+xKy7RoMeBLC65KxvCoAPJAgvMs96yvzXAcmjw
Jsw7258hfgeYlh0vL5QEJ+kAzxn2od3nmqmR0zOHSjBbaUCzTsiFTnAOB9SEb1l3
KDnNGpayKKknjpDrUK4yIj8iRAA/iKi2kbUvlMB0RcPYyO1BOaWx8SwaE2WPVChw
dWBiMXNOhIylMXwFi2bQko0ISnR/f5lD+WKrWitGa5zJSY4Qcx9zH8LPmTwEFWsG
tiA3Fp99eJ5Fy4ioS3WdO+IVnUqA8QjxhAv5sTFk9b+XGmXnf24DsKcC20sICDwJ
wtYv1oc4hl/GsO8inSR+c7CbcQ18Bzap2F93nPB20EBkoQhfrdjr4uaa/7Kua8D8
3Hlc8kwJlZjU2ZGTx4BRditODRLZugAAiFAd6/1db+k1Lrqwy7lxWvrOSpwXfspi
Mzqevuldv4q2aMYyLHW0DC0c16OZWeL7nbnOs19dxdJmF3Xivh6Yi8JWXaNu4fVZ
t5IZA2PfOkE47zk4a2XEABgEXcDOAm4bFjbsCTHb0SEHZf6HXMji/xk+blhd3I1k
lCais2ht2n2xT+7MPAIudFR2FcrkvX09RoAj61nUsgnui+g7NR9wa4iJTMKgzDvU
voFshCkBPsZkZg6XEXNoLm6Xg4R37uRf/TccMiP5r9Krk6yyOXmozp9dtvPgjqVM
syBgCLLcEZNf7Vghzv+T0JZ6IjCmUqv9EKXIK50jlzLER4BzaawpLlE5gZj5mGVT
su0OyiLH8iIR73qpy5yDi3U9B0GJk94/HBR2x3bQpaga0rknYKf3OwN7QyMCJD+T
h38QqJ/lg77i8nj6x+kMXw26tgfaFUnqhD4UICUcj7VaKZhFnGVApXNs2ysGUtze
UN4ehRdtvWYiPY/bKytpZoRUuEP4cODLpZBANZzSrwcMyOgVZ424ZT+sXqdohx9o
+8pybDLYLWphg96a1L9PJQmJxiMwYUEm9qppMm3nLbrDkXq1iOKQ3aI6HeRv5x6I
I505lKBcS6080ydoI36m/Pog/BxUaaDjsfUht/7iuo3syphqhqyLoTRSd705Dk+U
RfLbI/wBl1giB52jYjYglpE9DI8luvqoQS4342LCLvpsjBUUmqyiW5JnI60btdfK
kABITMy6old4TUcYAbDqejyp8K5K7j34RdRtiFtptyyLu6CbHr+iDFzQOjLMwW37
F9Tbm6qiLKVA5JXCvLuEKHE7bwIj1QvGmstNO79muagNgfyIMJjfiC98d4MPjOq8
3qPcqDPwrFKfOTArSPvqYLYa9SHvjd4cwO9tC3eKvzXJKVigBo/JtvZOkRexY8TP
H8dzzT1ZPLauX36JaKyqvK3kocgVuB2ctxu0ty30PpC01GXVZy0jFvjA/WetQLGC
s9tkWeYM3kcInNEiquqnuI9u2THYsNE8CQK16cOyPvFHfFYO00E4M1CaRx/foHzN
oDwK7npK6fR1xm+zbi6nPnn8l59+zbK72FG8gouLaxlMbOTZ2rlIXKJDZM/yENWb
WiKqn8CViynDoNsU0Dwk/KRtCG9iwvE4YDrfx3dvZ55ry45GvNu9pzISBNrtM6nQ
TcL4Auh99mBYuqHm3amXxBjgM4gw6rc8SZLxCNNEAkF9hbIs/NfMQaPrrZWJToqs
vSHTauoXc7BHmFTyjKpszA6X2mvlMCk95lw+TuwK58J7YK9avsuh1/OF7wJFS20K
2JJdFBCVL2NbcbPXJYHYRLMIlEmAJMcOdyE2UgiMrUAF/e+HkKmqwbFdR/j6e4Db
YITWqRPwdUY6LKPWkFInTrheTPfVJyaKvJOWwZE/PUSGfm/b6IHBlXp2Suev7DxJ
zr0ggccKYVyRH7D1pAwwjlglnTxPtmo4d4Lej6EiDosVaqwb5RdRSQQoSeighd4O
w1qKMmW1jRPCZi++DDgncrEFY53SCYe9kmnRFwqlRePMPZYrfjwKI1xfjpgiCrYK
ga8UCztbFKWb0+dcgtC4WLTiVBPY6+jbVdlXmD2ZS1L3CqpflDzntr7adkUhf6uk
hKSJF3xHtiqr0dDb0m4sR/zSaBX4AApK2vzmMYFjyoqyMsR2YohiVdgU5lOC8g9C
QNleW7+gi3469gWktj0YMH2h29iHHc8FsI8JiX6T99OPtoc/OpzjW29Zn1a9Ub1O
CBRJWIVRb0aCvAUNC0o4x0ZyWHxlnglxQi9PHo/yZt7/c/MU62dJ9cV7M+yvP8OH
IBhua4Gnq38VpKYHvRDdOw3hudyGTYSAdEPZP2H8+K8mmdQ5MVF+d2QZJ+s+ioHE
WnbRjmNwK/F0PkZkH6Pt3INhezBXtBkxtm+qS4uIPd2IHlcn+kNOOGoTnj9XIVgu
JOrtkEJ5qiKS/DWT0G4fYeIE9Lmz1Q3z8NWgInVOffgU2L8FS02ghHwEXpRqjA5Y
kp96DCfDqOVXdBAN7xVvqxXHaKBGtAZ6EqmKoUGRu1b8qhAmpPSLqbl++UVcNS9w
QlnL4XOjn/bahIsLGGxwuMCsvbd3ZNUxr9GsveHQJ6WitPkg3yxz/9GmkIu77UjR
0k6M5QUlQXFwt/HsT1tclV0SHvEJZoE0ai0YZN0VwR4IMLIoQLP86rcip6gRbljm
0IaijPGXuFv55PAmIQsGDoIcz6MFBq8atLt7RYYbrxCLQ06ai32gAvhMm9COzhAs
XXttTZvP5jynmBSRkn2Lx5JdGJiYPYdnnw+SJSm2EmzimLoxQ5LiRaLq4cXTOQDh
ZVmddP5+IYrgAcGCS+jZlG8imD5ywFjmEKRZyi8BMMsF6GHr43YaaKLsbp+m7ahl
NSQafynA+wx4VtFZgIE8B/LgqNtFB5gJjsFbeywf9tr9ROWi1yGacAdgBW3CH+4b
HyXjUnC1sfxyXxovMgELpbXRfnfhjSLz6bXkzGYLG9vG/XYu7j2s+N/2KXe8Wwkh
seM6WiuGi5OkvDrjtq8ERSzNYTLGeLRq2BLCXQEAKU5AcJMjxa+E0EDUKXOxsSPR
q6wGlAGNusYqeqwtVZcqh+oWEE5kZTptxnvJfMGPLwfVQx0HD9fywa0shqR340TS
AAKIsKGj1TPCeYdzLDDM3rnGG7fQ7Bt5l7wEG2awEjpk6s8CHLRFZbg2hQVwvVzu
wbjKsQkf55j8QIv0OwvsGdx2ZWjJyMuOzChMbfPUSD290F5cSJbkSLkrxvbADoBp
8qKCdO6HbrpvjJpWV/OhKVQ4yq0S/+LTuykejLI+s2IdQqrWLYttkeu97tHFVJkn
FFH5bKKuB0Uft4cl711kTNNLyQ8M2m+R7QBLoE2+XM8umSnfnLF9X03BT8K6odQL
gfxyZQOOZgfmeFFCsanpNfQJC2LGrLrdw8uxK39xQiVQl4hbf56KHsaJdvwvYcK1
FuA6CrnRKuBAcQfv74iMn9z982xBDfjfWxf0VqyGOLEs5UjKggBKAAfb9YBVyp/w
3SCdvByG+nNq/oJnVgmetMXzDa9Cn6pYVe2FNVdtK2YKTTeGSkVExyKxMHzc09uC
TCQ0z4prgNplYGN+09qOGWkImV1r/Otegyp6bKmtjAksLbvxhFccAjOYUpyozcff
zMOlT3A7yiC8NT9CCnBmETAVPV4girfiZmf4CXX7aYdfImOC+mcnabYb7W7P3sEt
/r7px3LdIY56pL0qXZ1c5fGEpRR25GworT6yJPagXrDTGVFhIdEIIcSUtnDP4lEw
v1fAihH1dV9AtXt+4KTk5ZFQEtxnGwdI2euUL/OcY2+fYVDUICJCn2KUYh+61k+W
my3obTnKQIIVgUEmqLxpRpX2+U30OqSp+NegjJ2Nan9VF6MmA701IOmYnq6DIs0+
PvV5comOnoIjw8/06Vwk8QRHsx4MWNdg/rUJ2pK6lg+XcN3w39mYZGVUi2ZutUP/
n4VGUgj7bKNnXJwoarLS83wyem35vccEEDASXoMq5gAtKlJ9Ei2S1oAmOmm2xHR1
dUnpUsWD/zJE/+dTV7OIElXh9CodTeI5r6RL6T0S1SDZNh2gFcMgl/g3Ibne3Ee4
zedL6anSvHxnrOUtXRg2nWIe/If0N6A28wcAjGIY8oIortkRqovt0lUAkQtFNzYa
PRsj9YqyV6GckdoundOcW1kCpR6x18y/gH/PExqNdgSaOl+w/PzQ7JEsdPFvS00G
pDy/VfUCRaBnaQLJjSQ6qoes+PA5W+2Jh1oAbaW4yIE4aCrVPDcJIWk+lKgTngsn
da+zeosYnJudxd9hWGxyG8ZR0gQRJXfbk/Oc7FqmIOP5ELo3ToDyhCIHub/ItuuK
A/dEbDAe11sMirELhVlVdorm9gu4+kTJl5aBEORSzIAKTxueUuH+5npTa/c8UTGr
Mknxu6BSYRzFeGZaFuFziKLMCFdEPEXlDfx0f8ST6uoJN3F5yEyCsr7LNRL3e/Cb
ynpBxcfm2PHCq3I9LE6SmCqfu7eTwvORbAH0wxyVcpWPjo9CvPJ2qJvUua9VOlvK
hKpZTwFe1hfaCvfEhu4U6TOX74bNJkDtPvcXoMZGYnJ8Xj5QwQrFxqT9DgLwVloe
szy3rkA5V7dXSLYhQGP9qj6WCy9tJYGXKaD9LGQbMQs3lXuEAqpyT4yZ7Qo2sUEp
rqWhp9F5TsIdWbvy1Sl+Ucqhx/0L5VOHb7jqzknqW4LYvwaJeGfusJKfH9Gekchx
UpyMWq+zHRXVy02kbMuwzTofiTVbZuWLNK6kGKfngrqJ1zOGx92LKdAJS17Hspbc
oKeEP3hZH/WnADHxFmYrTV1qYGTOj75WWHZhITbpEwggJgIglLxOhHeJZG4CQTkV
/IGK9U868/TAbztOpZAehSLTBkSsp4yAw9sYuhKTK/KDA2Trin+kdtlwZhzU5mU5
paYR+Zz3/S3o8MZGVNvOOP2XnWhB6kxZX6HgZF/UTI8YvWU29PNFexgwChOqFYrg
1jzoTKEPdF2L77+VjhzK4TI+PLny3A3K5SGU9eyLn+B37SyVkOrYtLmopPornNRK
AthqX9JWPpwz8OeG6JaSbZVPJJoAwAZPNX3USpDeTP8rZ6uSasyJAiXXoKsvX4oG
1G3irWe6DjG5LBJyZWgv1jkPqJXzp8pC+Y1a9VOAex0GchICkNzrGaSFE4NUDrCQ
spP1WOlJPPbJ0jgemPlh3e56vUjpKFxuRyrE/ocr6WB096+Qinr+wtu7SXWytVa6
e92ogBHolIpBw0GKbH6OkGnM2dUVlo96aazaaLniYYRzAo5ETwt+MB9jSJHJtGcy
PPBCmMvcjD65ug4oUG+MXyL+V8vhfWs1Ntbn7bbMsFYGyKCHXVbifkWTb4BVkh60
1vbEM2jROdECxwLoXwTVncFLu7KFOnnmGoau8RDbU+3dY5PMKjzZs+5Vyo5be1DN
L4rKDcPQq5EZqm/hmH3YRkaOsReN8dYcRGZMyVfQCQM/Qn9mAeEYP0rB5YjSTISk
vBL946cz1douUU2t5oKUysytTHCdSlHZJXzFrR2J6hqPxWa5+dlwgtkxpkAPmDUx
LmAyx74vzFNVjLaFHkhUmWs4/Cz6e0HAgg+7Inx0ohKZsIsYQUi36u8eMoET4epM
N6HiqW6Ct1zRhKlfVFZpCG7sgHM6SrRo62PIkk8v33iCJOVKk5PLA1PdYrQFdso9
cfgehELBU59YuohDkse9z/AjHJJQ3oXwJTZZTp2PFBHz8NBm+MrVaUxP0TC/7TN/
GDQWMYoekHA5go/uSS8UYBBySIFEcwmgiJfvkiAwYv6U9akHI+Nt9QPih0OEXkRK
zjB+yxZsIC4ndL3jSuIpoYpITeXKZ7bgg1KvxGV7q+6qrFUEOK1mRO5/CML9kg25
44GA985Q9aFy5ZE3ePo+C+gQOgsT59r0Mr3EMAFvhGxPGdvZaQb8WsW03fSuDtSS
xV7yJKvVpmfiRHXHTHZmR5dOneDjddbe7PPah31B7gDzprFW6rGBPwCFPljOtmjD
5eeJzjrx8ceQVh7SEzmpmuc8vtx120+jiAHNCiln4UMhOSIr+BYvurk2VwHQl4C6
/khSIHT4cK2K+vogMHVc81zfM+OaUpvkLgQrj5ad4nwK66ACM2gzOkr1ZrASLX/4
/cXmVDXW0vonFEcZRyI+RnDbEmIx2Uk7snayOCgrBBe/PvS3ucnwMddBL0Uvu8jA
G96jDapZ4edB+Ul3kAWMzVsOtNV+kuyAVGCZ8z+Esh4hU+2cRKbWkoXi+lQsfTj2
BnvslXs12ygBo3fS3fpVehfc0wok3iPn+hsJ5EtCJF4songhH8PHvipsJvosG1xS
DLRKmN92LX64DNlmCB9SPjWrD1ZYyBznMqww1wpqyfV5WhykT0y56qs/CQwvKHn1
UkGvWU3XttbHQLBkD78NuBxR+Wupb4aeq0sWDfRBhQFElzowjfAtEBjSPosX2fj2
SIjrrpVtMhGSWZ/javPWmxNUPaXJhptO6/UEHuGX8XRRA1qjaJvqlzUBySEciq2d
Uasy3ekds8pTwf9lC80yV61e0weI0sHxsaLiwIwp0T9SodetErXw9qnI6CjajXPh
eGKBiXRztwXxkZ2ixQ5J4/f8ndJSsEQG97c1L7y2PvDuVAoYc3mynjrcLCJCAzXz
czLcptplb655sR/ZkC92CpIfNHS+ocuZKnWf4SfViglMqKJGsyhaYTwICdebnSzY
/Lvuu1O39zG6iZ+KhjlTgYSWi1mEMvkdfSQVRQyyZVwR6cam8F7/09SHV6ziPlsU
0f9jkxDXVdGdZCmveLG/tlXQw3XB+KsvIJLfBbT4BElNBEluQmK1QreB9evIsaRB
jcFrz9/tD9zcBsid8KJUGW/C2+kRg6jRJBdOzEaIuqQ+gPYsnVSlBxWF7rpB01Lf
5NoN+nARQXNPvoOQdALoviRo+PdThkZqDduFiuO2rYRf9M4So8FKOvaEQcnyni9W
+cku92TCsu4C4cH+okWFKXbsVCLF2xgb6W4MnTPwL7KCdpDotepnYXlfCs1soujd
uS2DQOepNopOcTz+Th4PUpc/IX+N3yVrHrGCke58KhBTlMzxKwePps2dryKfXxa+
mSUCGdLyg75d8wZYRgOp+8ew+vapd6UsIKroZn0jhFETRvSh9dwqQCFmQDZsRxIF
0xFET044zZZouqDu6ASOFcIJaGM1MJ9SemWKv1TEuRGcmV4h+IK6BPZk984eSPG3
/Wkbl8KxTSwGvdF6yJhrVQog5VYb5Pfn0CdXHR+HTxk=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8432 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl7TOuMe4xzV7rdHsSWg325uw7O+YzGFhalwnTHdW9CsA
K9rIYsmH3ne6o4wGP8jT0z/8vnlpidVJkw8xNXriRFft/1eUhbVmd1oFukQ9524l
5fToHr8o31yXSeJXu/szkqphPAMxvXusgefNl65sAQ4s/tZLFFH4hFXKpQXd1n4O
FVquj4+qSuZISi9hZ6yAmrTLyHpJ9guzmXvdlpmazbZ5u5ZewFfMxGaM1Wfce9wC
WGM00JeeuW/6By3kEPFCHh1aRX7yaoysL01sNB8pZ4HbiS14L5yhGNzT7zwBJzfg
TZi09AVKVDbIcs4YKXRCW3O1Q3eJ/Iz9R6bPeYcWBmUYS7MEwA5yDQF6yz7dWoBP
NEV1S3OGYB9xlB3QUECcdEXtCjePw14fcmkjPSBz2dsbM9ksFVn6007tNWZ4xt4J
NhUwqMCJLS70fi2/ZuzM+QrcCvBnx6IZh36kokEykF45ktDIjHwplE8mTZ2dPO9X
qhzyLdgVR0ndpOeq2h2UGIjD/fuahVbLqMW2dyWyl+1ax0axeokaw0m3Z/6OPgIk
YaY0VAzIojm4rFFKkeFRBjrC/VokIju0oNrqOduSN13lj/RVOmR8/vuaGjNhm7U/
kBiGwyJfzEbjrPU64ncKKDx/cN9YQqqbRLd8zqYi5m3danJH/twT1Xl+Pde2XcFT
qakVY4RYRQv9k1a8VGaZEUbLBwGa7Ol3ZQgftomaLb+ZuGaoHv86tfdYYShgr3p3
OV3emOG67djVWuW5g1TkK2nKjlZ68tbdZq4qF2ZcViRohwuOZt/fOeiCu/mxdJgq
IKQyAHFUcHxXgeDRYKntXEwPLI77QQYdwvOmnntiRroyjPIeGcIoBWTQKRX3+4Co
PFuJf47DeOunZHyqsTFqx3NRLSkN99NitecKp29KUjWBDJjpHvZfiYArQT1x3m4U
6m/zfw3H3N3pJNlvT0ictMbUcmlin8vrS5LxLVdTmE+6tPF2LdImAF2+EDaavTPb
Y+yCFXDUSdNaVXc14Fh6IbnAIV7J0CXsewzBQ8rg7KT4g/PZdPXwRqJNsoVsBxjf
IX0d7/9we/G2KgdJSrd6v7DvN5xgn0XgODY9/IIGptxUczDdc1DmzSPSOUlgWuZo
JDTAibnQPBHbC/+EReq95chjyLvDVCKYIb40Baq14ekgZEWr8z2B9mUc9PgY+yfF
6V1lMMYpOqeAWUSVJPe6F9ZqXe9Scowa9yQvnAyUQYAlc3z5NOAdWzQbB+DobcOR
QS8sOEtJr2zvcM2apjsVxz26iE+Szh+XU4auUIEBoRW4pRhcv4/sWwO5T2YIDX2B
5SKrUi3UM86ISFdlAB1+F/u9FeTYndsAGYPLhBTazmw2O7C1xL/7vtBtgZE7K1vq
Dpprhyu2NelebPAd7Mi5W+lQ8bPc//ZCjztcAM4eYcgdFPd35/2N3L4EY7sTseeQ
g8vbbT41zf9QhcapFHl5s60LRW6Jgblqe/tPhY/ZFGnNu9oe0wnDevCoFPUO1nj4
8HNZyvcNQZX+K4jRnjR7jjqqLda5v/IUxQOMd9V42fMuhDq1kGbAJ7b322Dy8lel
POPXw5syITWJoiiNBtWJ8Me76EpVvUjayBx6eBwPE7WX6zWEFKxpHYIKVmiU4sSw
vcpfOca9SCwEOHeo1pafcYT6ixC9brC4edD8AKcJoHVe3YnHaR6nooC/IurqjqjJ
30vVS7gN8t3r2usk3QbzLzIPlyOX4NqZaLP0JjDavahw+JVeUA3jd2wypHUZJ2iz
AtIpfBec6vIn6Wy7qS78CW0lm8v03lZCXseCsxVURjL0aLOCv7XHv8GfjSVlyd9X
91xaWfXet+3a7/ZoIVV+8fEkzO6ny9c98gHbKryrHUwYEUWG7HMQV2lC0nTkNnji
AukWSilIjmiSL57FHRDOBH5qiGDxKFixdcGNjo2tqLPcY07qWiLMkjQMdcRLu7Ho
XN62pwb/868mgxWuC3hlcDQi/1Su7A0W7n5zABo8LKzN4WBAJdcvLMKr2HkS1h+G
JECQtehFO/of84GUGt0E0SbgYGmUJ5Y523t4z8zDo3fNW5q/CAGvbHYPxzrVc8MZ
Emwx68bk5SuTS2qn20l1FnTy4w++YX3MZ6SfDeCVxXJxGEkn0RgGwnyoWATI7bRu
6jiLn6jvpYYS3+qvivVgc7NM5cYmYRMyQVc+uK0VlbbtI8XkeeWhTJNlcxO614RL
AJqWB9KfNXSHq69+v/xF/UrIXnVKCCNlavaHEPKvit9hUsbEVErBHUadYbXEBYwk
SWTLlCEGHjX67v74LCOJKVmFOmGZO7dRjCqIfV35ofLQ8n3uFizX1rTx9vEA7RRX
VI83kDm1bDU5y/F49QwoPSLS2dKDcQG4FSI+OPmUq2jzxboBc8pV6W5ci8/NYKJ2
5epvxBg5Hra8uHWIwyiMWBLRrlqftGF5/Bp5k3N8kgDrddpjRhEt2byiEewSGX3T
7VAbZPGBRXvCIsynuMhuQU0oFjvtheIKQug8rC2EPjAxA/4jp503CnlbCZyu+tBO
dlzciBs2xV28aeWSj0wBFEjqfKKf2RB/gL+IC8HaWtEksOcPPiFhzntMf+925+XI
LzXDArpLy/bK69LoZCEbe9henuoTJHvlbHwq4JZdD5Bx6titc44ajDNo6VEhZFh6
AWEfakxkw8eGGjLLYxs/f1hP3XB2nNHHi85HB2XaD8iRyNOP0nWWJOcDNBYRlW7s
HTQjnZ90SdtNvNDUtE9cyk6cN5Oj7QEB8xaIaR2lJ6ZFyYDXHYgRsmr2THcABePS
ltz32p8uXaq3bF4kkZvRK26AcSqVqlBshmjNxTnTKM6uOl40r9Mqwg1AwsXNIUZC
3YyV0J1s8jpvdIBEYEWY9YRjCgmQyL01r7GKED9mtRnzeGxPeoMejL8fCOBots3H
UuuyhObx88d9ou4XKULmPRR8SxgM7SJVOc7XnkmfEajQF97DfaWjLG5kdFCg2Pkw
xXx1He92ZoKnzlRz6MEkv++vw8V+sgkAfiwCu0U0x8+9Bo1FopmfJ5HQYShAnoUc
USRW7DYsPLEo/Qu6BE+D7y3ti83pSwth4SV4tacX9BgKGUKJw9WQObevhz2nEDpk
26csnrRJzMQgS0Y4nEkX9riXgnF0791dH6G2l14gaqZFfgj2nm7+j4WXS5FnUHTv
XAgP4zc/morTSgr6mb8p4bHb7ySuYCAGnRGA84Len68GVZ+rBPydZ5rNxg9swvua
uobYm4KC6IguJ0iskDiNz1pDm/u7iEW7lAlV6rWrUG4WtOoYSTui6gueOwE4wDTj
Yf2JJQQjef+69Kx4plPuhzq8wWwnLe77Z7X3V2uC+0YaAlxbjJpfLdXCZqsITMyE
Yhv4BMvcjJ9QhOA5BHrBmgiR32a/ZLIhGQQvuo/gx+i6sD315Y1niJgjpOpnkqr/
eXFaRogzxOZF4MVlnDSOIi5KDX0HHsnfvYGXwu+9SPzIWzraCGCPJvDCul5ToELl
eY0civcc5BN6oi9mLnOM1PzEz/K2XolEvx7wASxJ9tbiz2LNPD5xSWQUdOg+GGwA
qU/cU8tKvGgjMuqV6kUrGNqPTE/u8pG3lSBWdFeUlMm4An9Dfh7f5o2u0iAxB/K0
co28ZdatVSP4YB2a5qtpzu6DwQLoENsr9wrJ+aJuouDm/H5hyDaIpsS0b8ZQu8HK
o6bz+UbR6xRZHw1q4bCMrlhjzB1/HiUzx1iWtCrgLyRgcf0+mdtHRQWuceBbbh2u
YFPWl2XzmYPjfo+XPz3aWy4kM6cpkIPoe02R7KmK6hLlFcc0+XIS5gG74tWcr2BK
ahV6SuEkB2259jhxoQBKj2dBsKUfTO0fyP6fHb7YCOnou2OEPi5ltwFPaNX0uF+i
iazEDB7udul18caipoFGVuuyQUDbTIHrA5MpkqJ3rdH7ksYtC29ePjck2cN845Rz
eE3YsdsDfyD8YxVfha9tCiBFNg2fVzVqA0Q7QhBNOupQBPboLv+dPA3Y/w+1XJzI
uAcPpObR49tXoRarWmceJyc+pjd5/2DNoSoIkHTpZEdOmWp71bHZvpNCcMCyE4Ea
c/EQQ9TcfxRs48cY8nqclyJIQ6IJhjRZsGMQ8B8viBcxAc/n2htNAvaodxLJkTSc
HLxZF0Wuf3jNSDmGeBsnf4th3wdvtQPkJ68XfVzhVlTupoTAl5+rwthKx7hMl7sD
xZUJebA1wNFssdOyU+VtM73W2eppW55qp7aYx5h5TFR+0CveLOSLLQtVBMbE6WK1
Q84vSRO1Yeuk7kMa0NSwSmfnQ7NXUW8hKrQboj2scvFN0mhCu9Wjk4CGcHCwNRm/
1v/PhlPXmEPiAGGqAsePzuVMFKVxByRcUc32BzNAaTqAMzLQHkcL5F6GzGYCNpj1
q8CXhBqA34T280SMqyBk1HiItzJ2LDG2rNKfMBch6kGSUjXHfrmR/QN7Gptcghc5
MA41hCesU/SFX2Kd9mBgi9M4/wItnNmNP4q/kfF3Ws7g0sBVTrYgtAGL9d3GeK6L
50TsoJLQ10I60ChyDrD1W5vm1RDBLzQwVWze9M3A/kQz2OHIT4C28+t1C+/3MnNq
OH3i4tHQTIBZUpinHzB3JAH0/AvNwNMJ5MXRXcicnEnDHvV/N99HYblVYRCAf19d
esFKPh4GtUMmB7mJqqc7i1yQM76oCBOEqcks0Yz/UGJKlmAWeK0i0dUn4W3r26uQ
BafmcWrVkItsLDH6xSeOhgnvbj50uqA8f03ORwT8u6kfrIcNhKF5RwlQchW7EHUL
Q/rIbYCZzpt83keFR5Pgd6saLqN4OzXCf71cQEYMCs5skEKnUz4Dcbc4uJ73WF0q
hP60jC+09+RHUxmuh26jq8Et/UZIs2yAHb3nGZ2FCyxdXJQh//kOSMGMJgthETVX
x3Now3bjP39EEHFWKPgmEyCokxQaCQ0CrSipgOj58NA3WWS7zSFAu/yjRlbwEEgB
KeNv8PPz3A5kXCp+dKJiGFORhWfKmLNwlze+zFd4C/KEmtR+4WM/y3KFf+MvkMTh
k9RmEVq6vryOIg6txuXGGxKF45h7m9grI6J1YKn3/eEoIFEVomiXydgRP03XBymH
HEmOZHsI1lRM8G7s2zT1tVxVCRgsKrbCDDyCyXHJdpwzQJr+Bu1Ph+EXUOyphKOM
CQsfrWGAFmjVNIgByJGBp7BkNv07iNY11/lUxLAObdRQ5xp0pxSdX4rjnG+Vjsfj
Ks+ZThVfTmjMXa1FQpgtY2VGUCwTotWbm5fuZwAzzFhLUBFQnt2q+piOX8MOkcvi
Gt8BekouLVrAuzNTZRYjMwMoMOcHWsLS+B/hB6+Z02AtBYptHw2p/U6DFg1iGZnD
iaCx9xf6rFN4USXJ/xznMCzYghLL7MaaYifRKA7Db5yKfCi9BJcCyt6pwgsJiwhT
F8zUnURAT3yjlaTj6bbLlM/YgPR6b3Bih0ycxcBn+WiBohLlikAtvvV6C2jDKeUF
Mu8SKvGtqpulsb5QxUV22FcVzATRXgHr4LsUWVaDsexcOe+jKLOSkeLqYb3mnLpE
cJmLDDkczLwIihYNMSRAc0qhtbHHnSTZST+mWALpzzZnTXLBX5AfonqOl+PLkiNy
NUmKLBPtzu+IDzq5ZgsjNqlPSRMsXU6MvuGfwgCG7IywD8dbuMgrZ7VHl+VNTgzS
GFCIpt5/XmCXA36QZSY8cgmxeGiA9iBokJudvOQpm98G3i35bTtEqn1KnkvGrRiX
geWeIbq7H+e/julyMfsbeNFtSOUxyaLUFBX4/P55I5WscJE0bmoZGkMzkRJYjfWs
mPNo4fH/7s3lckwQT6/xhceLgo3TAx1exZlua3KFaRHbhorvGu4aKpuNod3atVxD
LY/ceJZNTSIMC4YpdmFHsar82a8IS3CcP7a5omKlO0mp/OnXOuVwsoCoJQ+Uwan1
G8OdN1Ib5SUsaq175DLcVeg2T+YtBMOeYLO0mYVD15pmbOnJGLTbkHdmv6C2sMYi
NJL8+YSgwENcPwGB3ew8sGIdF0qJcifvx8UGfhMKwc+Sc2Rss9V4ux5rBzd+5M7q
X3kuZ5OgCXG8ZQjcPJwRMMD2RuLGHV10qJAAKDEWdtPPz24tyHtfjZByGmNAEhp4
WaE6ul8YqPpkvkYi78JfZX245t9kci/28kMYkGnZ2T5CbGsXNgZif7uox+pNcfN0
uBLotzgGUdIjUMmOP6QtRZNdIae7YHRphXag0pT0ADEC37vkO1zjcZC+1AmhG0DA
BPez2C5Vgc0QvjPQ8te+e7J4eITuGrnRaZ84zrZWd+x4+RK94J5IqP50+QEl/ixQ
RrtLAa9O/QC2kTJ7lSjjkTFCG0nyGgT+t8hFeeDE1h6gIKAmnSBhjPCCF1mP0j6B
TmzfoBEB5EvGvn77NUdxnO3mNSNt5eJhFYh14euUvGWI9Gbo1HkF4n5+foRsCLyi
eb63SqK/Y+Spd6135jt+F1B10mEKUlMoctSj5ZZRVI5I70jfx/BlzSPHoTuNwdeZ
7tabECShrJDUx19NIuGmUoedKvISa9mGfOwgIbj5vuwGkKS8TnG/apDtwKNhnlwA
Azhb7+o93LQF8Np2jsQovPch2fT4nKw5xRVB29nTzRzDnBzbm1WXhvN8O5mw3I7X
O/JNHteUrBUvzIDCl4WWOfUj7MkvLIeK3ex54EPJPv15igG1mt5+2TjnTciCWvI3
RLukb6esr0lnFNidazohfhqKcTKR8Ft62g1MVSlyx+56bYl1UZC0JWdbjAj4zXBz
2dJjJgaRUgQd9oLAm9fedLHys19Iy380PAjtw7Cepu/7M0k7paVbUbzqxf9ukvOi
S+yNTyudme9vmKGteziJc1aJgyNctoEOmdoCWk+58WQMZOGg+eySLBH2ugJIFxFt
hsA/TzeqmqO3ZIaTkNAdGMJLd8GQTQx5g9eIwI0MaLCPg0hjs3WtK+rhYHh5NDqT
rE6UIHVqhYT+YhJLYVNiWub/Iagi/bp7U+8/012mxKyYHZ2n0yRKszPeNoEYnoj5
UN5UTD3RP2lF915bITWXQ16hDmNEO3fGi8HiBoxigIEFu35+MAoLh8sVSktt6/Mu
lO950G2YHJvVBkmrPwaqh5GbyU717C5vJnnRGQ3zJobeucLGG7pOnuag7BjiPOqO
INjabia29Y+GU8UfhCiD3Wc+Xs2oOggVDtxkXYXiJUwaDVjlD+kDxT05bRBnpnmB
cIu1jBfiuw4RiJOTZyj4bF03QGVneTpT7dgRjjVjbe1c8aSkXe31DBiNWcXsdWZL
JdlTs9Wz+a/z/9vK1HeL086D9ZZ9iW2PzfwNOiaHpqBfYqSVI9skatNZZwOrtOYa
oXeUzpkpdEAGAIgsSI+WV7GgGZ9zr0a/LVY6K4Nh3Y37XbKwuEqAqMrLRfoyD5XP
prqlcb4no2voyJt1+AHNUCzbhgj28A7yTfKpZiTXtxo4CYLWSbhTRF2XvGi43F4z
qR9UXJSVRNf3b6l4fISChC8a9C1XvF4frP1B/oJOTje/TXG+gPyh6YNsXlyBCFIW
uuCQ4hVeccQ0gdAw8t/KjM0xaoHXadIjemdDC04j380pM1dKjH4qUzpmkD2OUuMm
/1OZhG/Be/hWyfcgOc2yjW/+4WeHUndEVIqn3oFDqYjPM3tY1Zembyq8ytTolIKn
Hb8fgQxetbC0Yu7FzU8bXIYeO8YgcmMM7OzpuZV6IcEClckKqDqazto2J0vToP8J
0bu5s9kaEun6kfpnOwnV3WhIderlWV689VEE625tUBH+bCKeUFxF9jBbhte/5bWt
NGR7YGhiuZ/hY8FBZfvO4iAmSXGINqIt+LXno5qc3R4cTbjPjaA6gKM+RZE1+BFN
r82LW7rVj4WOlOjEEc7yLQUckJ+vnuIajpQhs1AoV1m0CpUMw1eKiCn/98L5JeM8
O/Z55NxZxblm2qFjnLmxfgCO1s6kJmsfW+V/8bAe1cxSVylCxLb3YtcvM6g7CzLh
v9qBR1SaAryRIKz2dJvFfo9mE9pWlLjGGtyvSvjY1wuKe5OSTdJan7gY33+AC9da
6K+HOgMLzZfAvg0VHEtTIzTIezIE+GYi19vzeyE2TvlB+QLdimxTnBKtk/dXn7tc
9oQ4divRKVFgzOnjUdIsJ6v4oBHVEZpvGDA+uCwxGqWKuTPVQN+fPSFBSKdi/vsl
K2REzhw946xM5gRtENumgPJkQpXznhF+S6OxLD+7K4SXejwaE1n5fSnZ6nX/TDYW
gSXYsx+6DUvVZ+9MM1x0rOh6WroYBxfrVPmcaiM0RCBFiQ+oyPS/L+FKkn5P8URT
H8EN8wbbrBpSZa+SLG1AqQlWuWXkhQkhL3ts45ATC5JThew5k073COH9AHeAvtNL
OOyygjHA1QJYJEZC39/rhbUPKyKxrmvzfrNYgIfoTlP0nRGXzHt48I7YijA4f/0+
xKP4wXfaePdfcKq9GBXrgRPm9tP/6DsAaN3MJuGiAq15vq8rBYQZdTPH8aqHrbxo
uDI7z3yUftWgJs55HpWIkVgVkIrlDH0AWmQz67OsCtTcRSxFC3MSGWxcxUbs2R3A
tK3xcSjRRVYvoYSXRaTlj8QZp1e+2LN2VnklS1TGwenHNSceWXLQYCRsEh5A2m5R
jeuDJlhzaRuus9MJYm0IfHtSQWcOlLkdeEoYgIkztRXQq/mPf/Bul9m1o5XCboDc
+fhio2CPj0VYv4Gu8x6EJDSPS02ZKls+MavX7Nq8lUFlEcyqM6PiKud7oQG+RW5r
rRZb03Vx8jl2ExodTJs8Hzwz3decieYYJT8ZOuFl+0dMx1AZfKnZDsWQ+s1F2MEj
v66gTgOeTtPR0WO8NToawutR3KwjD/yBsKIY1Wt/vw44hYZUjuUDWKOj3ldWD5gd
ASmsIpJA4rRwN72hj0/26AK4L/3MjaPHu4MQEx0wapHfKR/a8vpO+gYhIR8WXL/S
nj9Ng+dMs4NI3FILYwiKQ12ifLK0lYdepqbMceUd/766UWteWnY4VK/BRf3DG7oj
GBHm7mHMwvwSVQxlt2+oqqnHIYyfvu3cv+4l6ykjF9976f5FChHq+mWaxsceosuU
e+OfCAuiE9EkpVsFDOfZaXGmxBbg1XcZp3q39wiAM4/lwfAdvFzf0eTZGsnBgWwQ
YH9hwCJHTykmFZEm0YLfr34xoDu1i0n8DPrKsfQfMWpEpud7LFaAPG0U29Gg4OvX
YQa39IUcHifl2g4ytDwQNI995BApaUX2EyzDOweF+sTxjZ+YUGGbgt19DMc68NLw
Q5K7/Rtf+afEhQWKepYmekhUJG+D6LG+VE7YQ8UQxC87GRGBK7vAGBzxzcoSlrPU
aRbi9Jadrr7Ml6edH3w516fhKIfUiNhLGRR2ls53X+XfRbmn/CPIudu9Ic0bD0X/
Xr8hq4EI1JKumjskV+NDuD6sHoZdB0skdW6+HBRKQrMVQwnXAPeYTq+0tePAfOGV
3Gq4BW+8HmJ2/nVf1Ks1rQlbnttnORGSBL8b3CAHpz0uztxzgcSs3Rbvwo8SrkKb
D+RHJ6TEQ7uHn/sGAzqMAkI/aq81ahY3e6ja6wFa+8M3x+orhn0GU+6K74BWqGJe
eUFqIX871y5f41EMt/rpu0rSEuR0SASLF2fcwBMBGvRcll+h9WTqAw637awjDMoq
64DqGi38APYHMJaAxbgJVyw9fRHrOqDlYHriEahZ/MM5vRyH+FcFSHc6Ipgov22K
/iiuuI3lrRk86q0ANH+JbUAuRPh6yfvMIOJyJGaqJdgvaiQR6UEJqhqIM8rJedf7
b6Tg4YGncnQBF1I+odH5ls8yrQ+6HhhMRc3nKDbcqwEvj3RydBYrNW7Px3orJPkM
38LJLbsDuOckeSYhbASAr4wEZubwWiHzjhjD0sX62bF34ROPcrlNrsgeR69mF/zd
5jUWRTUsJwQ7q19sWLMvWqDMOGRVQfL7ieISvnJ6OdbSkTeu/i4WlAMWEdNtaHwV
xchbdbofZTImnlnZAku8+SXmyLTai0LKXgDSDXdhwBL2kvS8p45r05dYzh5xzedU
iR/TMCWfugF6nhdAY56ijCCRXLaZzo4jI4G3umbC6resYMkfkGDMyVmTV3s9nAwC
Ap5udlqki9HjNxDRRdik8KbYKuKZuZUarIodZdcK3rBZASCkpKoEczVkiduSNQ/w
KvKtEJdJbG/4iILc9ltDVcUwCz4Mm4NCiVNzvlXRbBds5w/t2H/Gi9bCKCSUGKXF
77rYKBiOg6llrAXPk2dtNC6GHDOfXcTQ3tVU2h8jaRoWRgTMsavcPACbmG/cs/S1
QjxgYLdMirGPWP3BI72Jv1D2nQbqTEce51ztzNOHiMwTWUb/faJS2yIke2O7rbXT
1BH2xRwqwvZyBZWWcTOb+q/Ghch+f+6YPZ3f2Bx1OOP311GPF+7jc3n4sgp7PqJL
DZiGcExPPUCdQdsOGramhCbCgp2/WgQNN7x5rN57ynmM1mdsRL/wb1jbCfMiaDfg
Ale8hz3BAjJuZdC1edeosn3WOTdB5u3VAWQy1+aw+fGA3X8zCsXbwwwYQYzlUR+S
gem1iy0D719zpAeHnsR+UysmT/jBTEk0OYz5Cn9tbgc3slTH6gwZwYIGhTtisB1U
Ms1DnSr54FcbdGDT2NHgJkUoaHsvIyihyH6djOdqtuDAUqqJ4X/7DxPZj5eVDrxw
mLoVZcQ0w/FBqG/CJQSOhOH+KlGnYbxP2m3gZwbcbZtnvz+wJZJNtu1SB6+6wWMA
Ch8DLcAqXf+S1ytgMtMF/6nZ8+B2+Z6JL/5eypYansCTpo09SugDhA72G4ydheOI
OSa6ru9VKUPaDtwYr9prJ6ZAhKIM6REB4tlrMmQcse7F9JWesIgFzyIKkeMUVmz0
SlFxMHaaS2cTAIWesMPioF7ksYNaE1gTlBUHTZftxGDt08H/2v+5dxw+V0TAmjuj
c0JxaBTSaAYrRfZ5/p1E9qt1wD1ppEtad9LMGJMTHOwAO+4s03gc66Z0q5V+EY96
EWXgJgB13iZQd2mpyA+y8Se87Pd9pUnKkowDiqVdRs6QmkdbjfJw1SZofJ6v3uUV
umNtBfIQpmAe0NxJ9aQlrl7nRu370JB8nFFoiCiPSeI=
>>>>>>> main
`protect end_protected