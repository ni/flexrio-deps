`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9776 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
Ju3IpcJpVj/VshHyynUPTDCo+dgLeQsY+vdYN8sJUP1HReGyVpr8a3TTtgVHLALl
xz5uSiBt5fNelWoMkbVekG5f4tF4sqR/lfyQwlx+XPWkLuZir1JDWRYNgFTXKer+
LenAFy3XC/NLNaF9k9B8uNoRJ2UCkeQT0bMo/OpcAEnNOoaBHKzRjeTfpAUvhKcM
ebr4ahVw8sCXn02nGpC5NXCQG/ix+MoIRzIdxDNF5/Uw3JvXE/XUY/wb8EzsWsWI
giPHfaBPffHxofEG11W8OHSsCh/8P9nkpoWlKsVtiVX6oiH7ynmo9Wn6ID9QDxma
0gJphvztFUi/clGeWTWFCE19EjuRHl3oMw+jNF5Nr03B9DvHzGZFoa93XfVkAGMT
+lvf8tKfmDXxH2njj+A7PBankRtWqv4JSuvRwakNkTCTBJO8GQw37k2NA2Hs24m2
W/fLnH8oPDDOErsORvO1jg5CFOZlNPIIVzYhjItylYOljkQS6WsGtt0ooEalnaEP
tPkApr7GlJGzAZ13IsD4uizdMf87h+WtoR0QDZedX7qiEnvOtl2d/y5rieF0BksX
2qTa4P0mALPlOCRsEBAi5rMxm9dMIgKKRC6XTrI45N1xMB0kgvzdnJrXWVGiwy/o
Ql03o61E1b19CWxDfJ0ruaD3kWAumK4DUDNqYulG7e5bfymXevb2e5NaUPdoUnMH
d1bCbSkLMXtCwl/Zq2TdhpL7Ci5DEck49AKe93gM6G3GBX6AaBkRYPjHQO9qfc5U
S+yNX+FLf3NhhVDzHHj6JmGSiG4SDMPpmxPW6pyzqbEECxcj7wOkuornU8LKtTRp
9cyUOdCF6Ycq9+Tm188+1pA1ibV7V0NbYVOeVP4Nofer2JRFJZbqXl4C4riuW7Pd
Hlp/1aHJZP0He4B9NYfoG0jViQw1QRW5ID/BatNhGm7mB+jtRcWZnLXu8t4hklgG
6gcoLLUFsDv8MzC+wbmFMwzyIvjK9P5fzMTG0T019t03+xjzGo/9luNkUb5WxT1y
+BgO7qI1mOOx9Q95s2DfmaVM00e2sVJaYZ2xj7Gc2a9nuT5IDePmM8s85rWGn3GN
aFr/qC3NT8n6mGS+oM5DwxrLOV8Cn38GOVgAdn3XAhsZbwqZuFsjkClq8+oJmrr+
wQp9Mqt1nEj7+r7rwQK6WmUstZnHWu6Ex2YdRK9GmhDMczxuoh8UkW0MpRzx+1+D
tAaPzg9zssl0Uqf2h+xwZDPVhJHYY6p1iJmZ+asyjzDi3exn5Yl6VIHRsBQppeed
FHHrvP8kNsNBE7qb3iBTBOEQkJaZtaQC0BDehtBUCm0o0ke3fTFOtsQdPhXjJwBU
NwqOY7Mb4lm98yoUlQmspx231Eg6BMjA/awmOkQ7NKGsQAGToOs1mDCKzR9a4JQR
jGwI0iH0I7NsKTIID+gZ0CMM+dlBFUA8vnKTTCnkNLeHMNon5ze0LW8121cO4eEx
hZnWFrYi55Gs96Zhjg0iZwQ36BIzjwm+DxhdpJ4yx+7IilcOMcDmglPPt2sShnl4
HOU//a75m7FNj7VMQr7VKW1BccQ7SN8LRSoQQpU0OYokgv6tzL8yobCXfTTyEYWY
SzC3oxSQVvJN5n+rpccI1de79VKQeHfe07HNaYte5PbNwztj/FjU2IUohYMNSTNp
Hne8nowEm/AdP62BLFBdtZBmEzID/A+In38SGuI7DSxUSp4c1OwmBdxSqBI3EkGh
lg5JrU39W4HvGRgrGQ2NR4hzT/xKPoWPjDdqHvD2TEDutTVYE5R/qcI2moYkiKTP
DY5qcrFNRC4Nf0D1vky2s1JhV6EzyHXIyWoiFSiy9EEXTv+jhekjuyO7JITVLZpF
/n5sOXLACJNBH5Mheuh6Nuy8dGXfWLIthfKcb2RSak2yHbyoHkTWYELvk+rIvh5N
S1ajFgs29pIOq02JOiMuyS2FYA9kdEJnCxysof3YCm7NwePJvDzgQunEOnzPrzVO
3lEpRRQYJ6DHmsDVqk038ArgIlgTUPNMb6clZk/Df0gJwQX303Ri18T7z5lJ1Isb
XDTdIUXMCquAJWVrf0VIYDRmSXPlchiCyBcfjMey7jpY4/8lwxIdx3lkYsqPT054
6qc7CVNIvm2DxwjweVhgfpV9QvriyyaZXQw6kytgb07ycjgM7UVwTYL35wr/ibuy
DCfgrxWKW6EqQJ3Q7Fv0NOMkJJyhoudlN3W2iIU5JDasaXVKCJeWp5mv8pe3KnFT
8wg4JNX3vPnsLycFgrh3xyn86P4AjDAUxRK8DxatreAxwAjXEyhQGkSni1LpLtpG
xAy4UCDYED1sC44/a/IJE2/w6U8FWw37qEgf7mmbu8eWbf3wUlciCliH/4VNbBCc
6sHk6qLYhsZulZYiPSY+jFpx+lZ8rFP1bIXNt3636qMRSJWi6+NjhTIQ815czOei
qmD5AvzLLC7PuOdl3gTEqTSHBSaZNNPU+UuCseKQMsR1IC5t1bBPoSoed7N6JuMi
xGILz6a1pwcEn/e2A4XLCBBhkJ8w9QgNpvXtHmmLpJGC3UYDE03PeH/ugU3BiRRT
J/hElLWZnEsveMc8gzfaMl6Jpqw5tFoMe2NvnmeXu/2w0DeHLqyv0TQCMZGJflmU
Dz+g2eae3emEOSZSWuUvi6LK5mdToDlKwnuM7qoDg3e2ujohwRf9ZfUWA8ivd8mu
lcTfRFUe/3QKlhnm2XzwcYAe1YKYHr/OnahGCbS85PYN18VRCoI3w7S8pmVK6Whu
DCJ04qVYftMlPNSPvHw5TeT1nOnSQQyWcn1dUeS/EeQNp0T3eoTjsqsaIwS/bged
yV/Z6qDw4WSCK3It9PTFp2FtDDuF9VwyF7CQ0nBtYA66IsUSZKIBkfC23ks2cx0V
v/jk7yjJECJ7C86tWetB5qJ6r1Fdy5A0Lq3DEGtr5Yny60rn75VZ9PEJSXgDPqFZ
Xs8/A8oQ9bTZ/Dnj93rPd5IlxYxyfUyJqPD1jZQjUqoHBOytTfHUauf0EGW8E5Ch
Fx09ypCtfG1XppnziyDwKTgaNIbCGPdNax2aQmQjan3qMXLTjueLNfppbzicvu7X
t52tjk1KiHFoaiKb8bESuRNhtE2+gDhKBDgUX0rurDF1lFcLB4PKLxeA54mPrtpm
Ij6/vFpwVjr/9cY7wvjgsLDBOWtOmGeVvEiaWfIKnI4QGJNEXpdeTebRCFJZ5t0V
GgIUlC/bRyqimJ3h2btZj8Y/O+kRv8dVfswNjksQLV0ZOudlFGk3E4klLWd6gn42
yHsLrKcodqk1JaksAoNt2tlyRW7jA5ubPV01G3w2Y/Jy2koKxn86d3OBrQ3JaBul
kz9pNnGeDXwC26D3wpftwLs0BujkFUvsxNzcYs1UVEGGTjXF8eHMPtr91ss5hL5J
i0brlOZQkCwDFd7ILwMphIQYATml8RhrcNb+4GWavAmf7WlHwfbipuGGM4Vxw/Qf
15m5cSzTtizbiFEbzODTLezFSLfX+Ektp191LnvU6vEauapXCJeZkzu27ySCXM+9
WLVhsqtHX45MRxEQO3/lfWsNkXDTYSWICS8XlWqLjFrkM5xR9BHifMEJxfVoaxNZ
qVInmxQKXxgrlEk+Xym9RuWENk9TsG4NqvfNLQJQOR/RmOCkwB5XEh9NW6jAiMJ+
mxaaUFh8/PqmeOB9frk/2HtTwq0a8PlXFgOYFJlDrFcsMVlB60dIIe9+1g+d/c1R
mUl7Al4G3HQnoMKOnFOPkZrUWMyZEhc349BST5IT0X1S5MqrZIhqCuDdMSHMbAdi
ZctsFvao+puAMT8QfkOiDb7lR+6gQ4sCX0joS//nsWwW0i9HC6Dw35zpaliVqJUS
J+J+GYItIPeYj7j7yKBXN413C5KIFmGHCTvfTNkTbBYS+HSNd/rmlzGMdCS7QNEi
m5BU6eKlxzamr5nF32KsYVqZED6CDgNRqweDuM7PxO1cIAp0iGGpjxExXQ0iGjtx
e0hKBNq3+XoasS99BwzslTVBu4rGjtifVzvtVn6AA73uMBq7dvc4aam1kwI0bIpA
0imV4c+qcG7jS7OM9zmSoBfoPEclzJxpeF0QttNhCe4p5KxSsH3ydcE+0njWO9EK
iAjcAZ51uK9h3Vxad8+HCk3XHftCRWPW8eu2m87X/t0FnqFe/9T8ohe1KWjLrAy2
3dCo65YgALDht6RgHcHCI/74VOtOrv7Oo1P6lphbQloxgF/yPGiGExHeVh1dqjwu
Lpjg97FUZVUY7Tz2GI/F95cAzq0Xhbw2RbXxxff3bEYOruhto6xi46+WcYRjAXE5
AcpnXpjtZiRgnk5ZAccqQTKbtgjpekx0mZLS2MA4kbO5eGnyEk/yRTm/HSiPwI1u
rFbEkmC/L3i38mQYy9maUwvjXYocyTZPsBvRMFYGXw70wQ5rbCRimDyIeOuBbQZY
e7m2e2f0qjYoYZ2/R6kZbBiRYsQVnZTSOHTQoAXaslNKSscZOGdlioS9Julv9Hm8
tU8kkNqmL4QFVHuULR+Dxxj5FB0Hsrd7p1SEtiWPtED2yqceEPBdnpEE0jXNeQNt
efynI/VooNX+4OmAdZ3taya42pMQcZangXNM9EIJE5pko1WdnUdSN1oSxfbSIJ7A
smoyUg8O/ZdHFxwIcYA29pH7wYDyUoupLLvo97tRy/yXRgTiKCVFMZuD16v/Yczj
I8l14rXVYnCVIXeeaHnyM1ElhNrryshaHUx7dfyUyTRqtTsmq1+faau5HtZgp93U
rFc5joTyN4oJkmHvdfJDn6w3If2GX2T7DIWE2LFWeUv9jNUdgjm+TrCf90fIkh+U
1eDN2O+9pIqHBM0TW9MrM6kEd6kr2SbOJsaLa7L8RhLj900Nd67c/dYPH4pau7c9
TNAZmP4rw8LI8UZaBgQrUbKCexN1gw70hZp0LBgpQcmI+qw5QiyJa4FQok3f+haz
FGgO6A3YUB1gEHv5q5jY/lswrxpyfzwetQryib2GJyOGARPqBftS6PXpTFNjRf7v
jl/QUUcxKTnMB50IAQmEfXORNOAQWBd1he4U5DA2JxDw+vrYb9LHV9AVjr1pvO7B
1u4GWHpXfRGiMAzeYNCS06L3YRGu0CInTcE9bz4zH0YYE5TnAvLdKWr6DIqh34nO
1V8/bERYeS+PjetUQflIj5biEGnsFgklS9/BV/3ASgBdJrIY83Q2y4Ehw8T1383Z
LwQzQImOPZkrDTgK6Iiu+L3tZHt1MqN74Yi2szhbBqzEqidASe8Xd6blzhj/vdL9
mg97fjrJlNMpBgXHqP3KC8FZU80rc5uss7LBStq9i4/I6gMewU9DMmuS4BtGzXXi
OhYo7M4W1xCJxih1fruGNWbZRa6dms4RE0PlMmh5ITAhoNF4m1d6kKPEyjg20/5P
XT7HlfII3GVr92vVK8cialok0ah+eadzaLzqJuxeGZ/pSjQVV/jC7si7dU0zwrv2
0BcKeocFiaQEnW/uswF56AHxbJ6mnso43cp9lx27z9w689Gz3+O+Qm3LBZoKkCXR
DyUWZgxP706iV8RxTIMFMx9yviEbo37i6GldJW4tZMqQWr8MHHWibX6l1YmiKDRk
JQng5f+MEajrD/jiOBp72L8xv+fesP+FayTfyrEaE/vjF4ZZecTopHFP8WR//+pG
YAW/Ho7mEghUAj6f7eyoBjaLLiWaB7fNsj28a22GWSNQtgKjYtpBcWP5zwN4vDxk
SuSxE7QOlITNmy8GD3Xm6cGvEgekNifev8eiRjd+NEY39rkri6b8Wgb3TlNBzZRR
4VIHatM0kwbKM3Vu/m5GNgs9/0OucNYYWuhg6eG604bCCT/xPbPPOZERr8NlUlae
jA0juedRCWpJUS8s4tZleBcEx09jFlTwwlPecEYsLxObPyKfJfM9u7ofo7eUFpk5
lZyBv8bk9V/uDWT+u6X1eEbrPUW95eX1fkh9OTd/uyLpsIPHJgp9B31xvz5XADgU
T9Yv17S85DG5BLLrk/Y7UGQg2jEjyssT0jKsklC6X+5hecz/dCamCE94OVzt5fqS
kvDhEiwifsKz7XfOBlXz7DImJ+5cYBvQxMCcskC28OXb/vQ9B9bSyD00nHndYvVR
aW9XisDR1j0bsm8e2VqVa40VtynoSsBlUsUIy9+3oPFcQoUr03grCmsMkf+aXF4r
CqhrWRKvp8+PPpZUM2lr9gzbK2a1OXJ7X1H0oaRY6m20agW0ynPLMA4OLWoLtAD5
hvxzkxux5SYzKyB5HFD/CpXOIbSHB0be9oW8sLIK8/VHyCWTtiXIDaCeZT4VKVz7
XrO9gInIeTp2KGLDb0CkeDXpDJrwjmQMvo9A7MAuvcW1A/lBfwNiWHZIHvt9albr
/fSlZ02uG2KEWq/f4UxFCa+uszggxGnCUvZi4z7XySH4NR5XqV0zwL4+Uv7NoUKO
ukDdpP+GN3Re69B9o8LFudtr7JBIui3cBrHGuKt/uVMsSG+RFAH77JUrda4mQPf2
5ouuPqdq8CI7xNzE/tLAKYG8e1dlfmY8ndjKN1unqx+DHP+gqs/3ObvTIoX4H8Vm
Oy8MAcpxajbaOeEehytVUpenr4WrzyQwqFlQz0uAvTk+a1ntK8aABFw0O8abq9jZ
LQvobZ9VnAaAQAw0TQVwFglSjUVi2Y6fkdbU9Lh8eBk5gaXvXWa2gGAOzDZAcNK7
IUO+YaaX9aggOxeKaqKsLQkOlafuHomtiuv3vhYbfE28rCASgGWkQ4MumDKcjPpS
sWHWV90C3memYoxBjcKvxYwsCzHsu1LeEGowh1kTNqPbkBFd15YuXW2dOe4HX3g7
xFM3PmkkuRPkKytNFGcNDiMtJkwdYy1u6CQUW8sgkW//aZ13op/WpqKoF+Yka0KY
urBAagNUfnXLlOeES4GMkF04fdY+XnITRPsfd4OEMfVMqg7ruW2UGQN0oRtyysoY
qhWdjCO0QjWk3kqDoNfGvExiJlBO5VtDU1hBC8igGGIpF3A+lEGy+hUDEfyzc/d+
8z9+McER3vemY6KDYjmqKzXbdmXK0kmBvb8U4nsSESdGUpXFj3zY99by3GbevIp3
Ja+t20CjBITirtkP3SZiIoTSgdGZd/zVZyyg+lKEVlGXtFS3FL3IQXqjhwZYG28T
+JGc3G7q8Hk1n5OoWSKRmkzVrsoOXTsf7OdrTn3P7UyjgOJscjZzf6HWR5lZyl/D
2zA+dguQc1p/S9TpM5B3hktieLEmo/pchY3+Ybccvod/2s7nC2LMyuZ0ajnoD+Cr
TWKFB17KV3YtkE/ualMZE+U1TlJzRo4CfMa7lKzCuraSRwNP+kFIK302hFjdlNfw
byslbUkMfaW8I+hvM7mZriZeYseSlOB2n29zlciebHoz567O4kqIEDtlpw64SXj0
m9S/6omJKA0CAv6HcE2RWspzKC69Q+SKtwP1qHk2h6FQfaR8dnAAsOx5Xx1iWku7
zHCfskYBS6dU5CgAUab/wVMQ36gDZjr+HPcSCTd8soP/KJhH2aApg7odCMhK/ekB
ENzoQ0J19TsKiS5Ziq6jgc33cFc3tWW071SRQvm1tEBdFdOviFjlQZZ8CV+HDfnc
v7dv50Q1NAAwMPZyMEbLgzzEfR5bSLfEJCGzoapc5FmWg26k7V+3oUMzHwy4vQ29
ULDy+t24o06jdzx7ATxmfMnOQbPLNGunuFy+vNbmlvX1qtta2XlMGZYXjd96N4jO
Y8ZU5uP51dHxgSJJFLNLdme1wAWeauboIYHMuTF6NYTmEdyZplHMal4GaeX0iNlA
F2jcv2eNTagbh+/zinPez5YG5pau/rBqS1BetMEj83C4UMyPc5ctsCvRG1UY7uDc
9XQhA2s1XrL4o9HFsuEd7tfcDT7Hhl4UZxEIlLH+si8o4rXefGNCMIlTxFq/hHas
kdx74nwNsOV9zg5XrLaPwFYFBMrb8mdoVvekMc9kxyMgc0XrHCUS6fQP87cg8pr0
AX05e+POqC1EQ5llETkQe3CQn2A4zscyxEji+BdjS+I0j6o16xeysPbZYNKf1qyD
VlYVR6vtAYACOyLQ5q0Nc9Uu+m0p85KS4aLrsnjufwCzBDs2WlPHMnaFFJxteX0i
80HctVZI6Ik8kf7+irGQRsyeOPCP+TrW35LegLw+cqrYDeZw+fr345RbgjIZAd/u
TI6i9iA0ikvZ4UBCl0EuzS5TGxZabWbe4gC7vMy69pciia2+t2NeedbIDHr4d7W2
kfCLrjKcqi/MYzGAvrQLIHAXnRXihtPRDPaq1bQF8ccWjA75Mq4aG/3nSQZNEWRv
iwvGHvgKE58AVa+rXNOyMiVdIgEI26dYORPRtkZst9bCAjqfGgSl+KVByhuD3cki
HOqRaEM8V9qRH33GL73ZQrKT2wVHRkenjjYgp0M93dwSt5qfzCulLuU0tjVBL9cf
i1bYgtpaeoU6LhiXik3/djbQl3z9uLfzPR1fro1zN9AJwkHNG0t6ERvDz3+nsb4s
+YbUJyansMJ8PQOHVjfaDHPgzaHJu+8Fk8XEdpl56eTflBRBBT144D1bmUDTfw22
BfZmED6jYNHfOEFTQRw0tdhLWOQ0Ol8i6Ukyrco75z39wh6RSzgICURGNsRTzTlk
MDJpyb5wV38pbelek+CqaZ+rbdUsN7M6cFGDEtTOUWiem3UIgqGi6ZkdA7g4hUyX
+Kj6S5Zc7y1rIeCl9YQM4pYI8EH9STYg/C8hBP0epAF9aK5iDkCc+ySEUpu6sKzn
tMk2lpRuKEga01qvkWiSDfWjHjU97WseQripq5LZ/HF52SQsMU9ssT5QXoFWDMGy
OyeZEaYCK8A5pw5c29RLKx8vxGRlH3W6mt4QDk5DEjDkMJwT97SoMpizEuxuZwGS
Jo7UteNdkcVLNLF+M57hzwO3CqI5S1NHzXiupHaP34uNKwGzzmIj5PTJRR8P6i9n
A0MAXlhpKTHCQvYzL+W3eschgKPqkGIoRvDMDzv5xoLbe1krJWy8qkjQAv4NohIK
7GPSFb08jETagXKH1R2B8NMwF24WaRmMK8+H35yUsZ6nEubuYAgXK0ug6VpeaZEW
jo8CjOs0waDqyLNgbHDaDiRiQ3omlS4tjFKT3UoCFNkQgICVhjqjXc21hTPcDwUH
98DbywxA9A8JN41ygr8shXIHNOTiUgnLl75t7fQ5vunaCdBTZLLt/+hDu+heRJUq
Q7cR3g63xZDSouaBzmIEJJpzoWPZdvEjgc6pKvgmSUj2I1sPR4tK6h+m8U7JAtP6
UHYaduKm7qgXUx5KDtKPHXtCsgmNqs8vrdAIUOs5mmKfSEPYi9JqRgkhpcBTUYl6
74EywbSsBE1OTqJFBW6uAb869pq9RPeqA8jXXdwMMd/FSPA/5s3YRnrTlS0CyJTu
dGUVGL7WtEAtkkA/8oJjuxPalx5POnE+dWmj6a7lrZzuI+wo+M5k4xlGCIhfjEOg
vY9jzWJWC6aEDqLfNLBESFF0VtUm825t61SlnjvLNqLznQ9ZLsV/0Ni18qhs/AKR
azZiuCMO+ndx6qYVdh+KcdKmE5g4Q4ja3/MC9gvjG657OEoKAG8yGWyu7uQSseIb
0phVnpT5Iea6FhjpQ+8+derhB1YITgjzZA59ohdbkEpRnQZX+H8GPDkyup3w+AQX
Fr91QhLFk1Vv0u1dtcf+v/RSESAqFLe4Ht6m5ybNr4GsV2BbUWnzEMYJFVDP4MOt
UFUmRzWAAgfMVtuMj57ZepSL1Y3oC0I/OgjK/oRrURz6b8FymLNEWyawyXePi578
u/2UGGduo2BufivLt6Ygjpf27EKz3Fd9s1wIBWubSvB7eH8qx9BKpobiTtBAcc8H
RlcVQZbuJhyJye4xn/jNwzPS18OdCpzUP0Xsol0nWPflGiR4/2gHCuAmm4F9M3OB
ut91T1Ve0bDDoA7TpnYHQQNBOQfr9cEh/cfnZZvzqQUlEdaIlu2+9eQfzc1XXGKP
7NzCp4YiXHftnp6sBaAMVFj0LO+a4Ekv+26jgPjtSTahuNiwbCEjApLdgHWtbwbt
hC82lTy8MgzmWm5Ts8WRM2+X3LNtX3YVT1FDnuLYoiUP5FCz0VQPrCV+Qw3twnQy
rdx/+gBIznPxKRVsMZDSR5MRHJTptBLDEPlIPYVgrOhb6aYOeJuJ8n9At0bMXLJi
boQQCknB8KDayc6lz96DSET5/1iNYCzgv6wYijY3PHGsDWBJQljocODHaszZ5B3m
s2DBQWEFONmbg5a6L8wm80QhAxs5s9XJxKwX25JpP3bwtgkzOAfaxSDcAIpS6P5P
ZNelnyIgo9I9sApRiVxDsP1n8l1iKl7Rxi/1McwSKK/rkAR7aFXl2e+d6bqlA2ah
Rzbdg8NmHvg1JIOaYApuJJ8lYmqCKG1CHPiqAJQxQru1yvciDU+5ZlOE2VrL/A+y
9ebPTRWBGgyzlADtiV2/jW0HfQBoRi1ppqvJVimLiNguspj3uJ+1tvpPi0E46App
eVT8oJ0Z5tuFbs9sykt4JPyEd5hAQ8gMVu6Mb1a1dPTKdoqog4XpxYFmbwFDYyQj
NsTUQ7xhPISxAnKxfU63lLQvrTlj2Gh/oQ88bc4/Cf6Zs+48DUtOP7s5X18QJ/hR
edvwtfon5Tz0tNJrhwIpVlJNtITs8a7oBo7yWgT2+fPIKjw7oWg2/qgonHidrryv
U0SHp+xnXtw43iwvkyRth4DkASxjjPtRwMJynN4FkYtHA1kAQHqvUNE//MnlmKI6
ObCTP7alUMuxpQG5wjPs5Zge15lrnY2+Xj8h6spCQP7s47LT+jXiGzcWVz/eyAy/
fsCzarCsCvdt514X0QXBT2/NmSVrphcF1GFALJWpo6pb0N8i4ZAlsKxLpIkhu4LS
9GQer1ac+ElekdtHafmb65O59obf+ZG6gUr/Kuyq87Wh+PSRskU8byt7wDu5xnJa
EW3jRmVO0eXyr96BNqfO+d3Z57gOlQaEZnoUstLZwop0hit/3VjRSupjz+radiSA
x9gIb/XUyZPd1pKk7GkOs1bkVhCPbwcfe7NkW22Cp78dqXF6xSav1U2DC+8TjEhq
2xlHV8UJjSwQD9Jo/t1ROHYmw6TdKNIQsyD3l02zd8laup6mzmpT+cL+3zv5dOwA
aklV+g8AOQfJFQ60USz+kIJtJnkJ0ptmaATbe3N+FfvOrS/GhgrHscz05WlUQ8up
HGlldxWZLFB1pHjAOeOxa/f5EjgwIz8yjZTqKB+D3ov11j1195Tm6q04PgZKecYP
YsTCE422SAcFuo6V1EIm2Jg5nfI7TrS+TzrchcgPtUAThsuynyFgAl8Gb2UJLdyM
vJx8rch93A0yoPRMYKy5Vq0hPtNUxx2t0fmNSVjQ9ZWldS1Bn1Z+hnGTidh7+3B6
WGzJxMHpBaz1l4u1mf2MeqQNA5qdyBX1T96Yo6FzDdS6WFLtgVrGZlVwptIhWbpR
L6MNYxEYjWCsPuADxuV0DvsJMbgrGRrFFOGNqHkfSNPf17kltN+HeuAl16LRmpXJ
dtFfWa0tw6FsnXGP+gwhXRT4nV1F+ghcJJyfLGIrCP/qcA+mOWjjcDeNLp3mPZ41
VKeOKzL42MQvvMsG+RWIQwvSYfo2a1agKYj6YRK69HITRYkr7mk7VDPQLJzEyBvJ
ruw47f3rRJtDfJd7v5otdhEZdsJz174gCZh5a1G8uCEzD63/Bd8FWeyjPGRLMoZp
peAHlWr4Rkx3RxY5VxM0L/YsUeyiSF0P6VQ/wASxlki8oIDdn4owr/HAUkoPCu1Y
HbvRJOfjRwTPy3LAs7YmLjDh52tjN9/UPfgZf8iKN7HsTPvR0dTzShgRL+e38cyC
aUS1DmI0bj4Sgncbli93wf+cQGuCVZMkVKrombW4P598FDFVOX+d8Qn7iWeMez02
sm7Wx9Dou417X/oqTg2h12K9MLtdruupASokZnrzBa3MGgXsduwDPi9XLxAtN54S
MNpzTqU28zevA6qZjGYrAIm5+Ff5sEGThMq5XEXBHnXW6RVTNHoQA+0pAB+3WzHo
i5grhgH8FmsxyR+xk3HP3uPGeafW6sGr+LWaKdi6pkYgQk/ABdd4bwAqf5oI4c/I
1DTZDdVwLvQ0OwYrGALlGTtM5/2ASOxE1x/OjvIRFLlm20PaZ5YrwOxIppPPsuwO
j/CH7i6jtBkS42NbHvgjolK/2G7cvRSGyRUQ4ZWG6MFXLgHSwmOJgJcLfSgxzFAT
ig+TQqSQTm4GwclMSMaKeaJ1C+x46YYClmnLUswyYPKULz2LzZAdBBnV+TsZ66Kr
+2gDTUH7mHFYP6pH9FixPK7oAj+3XgYwPlFTPl23rqWVqwp/Gxyg6iZtTq4Wmoms
DdVhz1N0yZE0unXie0+iLt0vbSgEwMag5ZUur/t2Y/PeDth5M75fiPPs9HrYzn4w
+T1C+yGmcJDBKCCL+LlYobr8ov56pGbOV+i1HHKKLYm4SLbT5YpyP5ZV1h1kG3Vz
eqnXS7qkif+QY3laie7Enz/gTLbr6neqyFq91/lRsYYDwTHsjDPPPrroVlKlKE9a
L0l7osCCjzCdQqOKUniWTelQVJtLGmxhD88OtlgNvtI9xlahzPclFVWWd3JvF3rg
XrZ2MBbJ+YBGfgTYg3nDZKufgPNNbOMI2pFlwhM3AO3ALc2k335wDtXyA4BTL/z1
4s2psHdsPplNfsCOGusyJMVKbPHdyuVuSDWfOl/mLLKouGLikEXsE1kcn7IluSDt
i52lI93n6b5Mp4B4xUcPZq4oJdvgY/pJNr98x1/2X1hIHCmIuTkxyWHgvei8h5s1
mMeQ6A01aFIKW8PFaI0VyPPcePcrHA0IF4NsjBh6cISevfvKVDzf8QQw3yY82T9C
+qDCu2QrvYej/sMb/nuCQd1ZOVvRl5195jnq/jBlYhTUT/5JhMpxf1xdQFIyAaVn
9wYY/wuLXjGkID06NQbmgqQWAChN/YpsvtNYFN6e/CA=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9776 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
lmOQgIOM5jiJrGbWpsW/8nEOaDKTwcqoCqQfVLnucBDjo5tp5a8G0oquz4RWYuq6
cBYyIFvQANKw6juLxTmsm5l3VED7aqq8r9RlRbO3L1mie5m3MY0z+7NMINBkis8y
mQs/Ra+Kb+AaDae2ya5JqFJeO90MyNZ3g5AKW7+QX4yS+6rmJeXmgS/8zKrDhBIn
+hj+FDtgP+64LxVTjenujhT0myMx67gw7KWc6va+3HQTTJcXLjGqhIDKtcdCjRkg
WH+0unSjr6PVxa2pIlxIdxv137Js+Dwh8SWWztLcT/hd6LLeUxQORIR29y2ux441
KUcvfsHPpWHNhLmX/9CBQX7Dp1oW6ACi4IDCN+x5vDjKCQkn1yC6ioeKkqfOReOz
e29lLdqGhI/ToF/hmnvTmiaHh6nA4ZlojvJuXAoKkLk5faJowsPMr2cn9uLx91tC
npGIz/dgJQnS037Ic+l3vgO/qT7ebs6v6LEp2xhCXrUYeG3kkZ08lZ8a/Rw4BBC2
iinnIxfq/XRNb2vVI3XzKdQwX7aHPqmrxUJy8D6Fe8CQ6mzdSaL5i4FYy2T0nFQh
JJ/VLhUQ8x7CRNn3Lcq3Cw85OKExS+niNoMPY11w774SPrAf3suwugsoUn90+L2r
2fRp2nlxiIHJmpbLvkK/B0PhvqsoRrBdItwxoh+rIXZDICCskjMIMxd5azcbkl0l
zxgEbw1TvJFqxzbVxpUNlxLLVloDoYO8Sqx1//Mx4NMDYodG8hC5wP3qFqPKzIK2
gLHqdOkhl/PJBwYrOa5S7FkuCnEmOXGi1HKhs3Qi+E94+B1olis08uX84wm3uw/r
9Z19eweTo6tXTK3tEoYYTGIRu/B9BqiENYiMp4l4L3Wuo+c3QmL4OpZ5ZYy8i4VI
34b2T7pDn3QGY0nTYDqJVNtp3Wb39mKHZkKAFPLB1djioxGOieLggAgXQLXmh+Yi
vIRENTSN4snbsc8WEdw2AirwuNsgnt770s66GyniWbpZpCUipJLJtwfSkMIwBRwp
uqFbkVMQy+e9adDh7DzCnaA7CKwiEmJKRK+45q7RyY9x3OGEEOdOtTqqrpmr3MtI
XEDwf2TQWMUa/D6MQLpWvPC27Q+1GiCNk8J1sU3skwdyIShqTYfmsxUCxgGAAgSS
aWmY32sDWxOs2Wv1TIaSTDGUNoxkkgbMPx/Z0dg3/O2r8DUJIDgv6ST8oT650O9Q
WfZzbIFtxtATWZsimoKieAKsRw4U4SOz3xazi6+rZXLZEP/PgUXVNQ+wYg7nX3Ih
eLXZHmA7ZFFqFxGNluPy8hU4xKfaPBDedXy2Ku9llouHFM+K7psxW4O8yG7kzpwR
TLF1UrQT5pW+aT6k7+cYkYjjLKSmrqmrZSBqOUIDUfImUigy7HUf2p4vHx42zOr4
kIVu096NI0wSB0oAjMU6EuLRlHqItHMG9pHG6Id1ECYXu8d7KnrIshQv1RO0uE2p
GzaX4attwC4+c2yZt4yhfatDfO3Sq7mxLJRh9BV+ksasdcsRUXzUVjoH4gLdaxp3
PrQjpWC3GyWAXKi1ZX3yWr4zwEriphyvRSAcPxKKP5WVLJ6FijvOVAR3oeph9hgE
0c05DB1cVC11DbkrRfKjzeI9LzrLVck6IUEl8UkTGy1dX5Z//QbRassEBT1Gav+3
U2J5UicgbvDMbxzg0FiCD/S2Gvq6jufGK71y1ulu8tDFEvUcKj3zHdlyQ4JsXdeG
3Vamnr8bfI2t64qlsBKjin5oLG31JPmv8l91HR+5I9E7lcbuXvAHUVBbhn4T5ck/
n+1mfYMiEghiOBWuMrhnkEJsLNrjIRhTszIiT7U8dy/0BJxqmcp/aXj1aWLWsibQ
ZgHsNW468suX5fRu1kw1okY9/98fk2p/+NUzveZY4Scv/QrT1EODspjaZxfSMRee
rVHXrWmN6PY/P+oExmCJp7zMzRC1IjyOZMwRg+bVcoM/mtoQxnq6kNKCQIMTQzut
oxkRqXMFGBEpCvjMRzyX8GrQbm/391JRtolEdpcaNf1km+wG08e3L2RDW3S1m2ur
JGowYFFveu9Bz8bICxwczg6dmb3Ix850oJ68DTN96NkYAMXfGHgZjaXbXQFcxpgk
T0v1PH7ZV7ngqzlY0M5KVyMwsY+PWMSjqCp9wmQjYbRs+U+5Y6IMpEWhXkbOeOg7
rk3Mkl1ndxPTl0QvPSv6AtEcS1d035pYpJUUlNjTCbkXD9GT6B6RPEvXJVHL/ETo
zgT8kJE6ProHG9Rohvwa/8Q/GSAp8FraH88Z2Y+Hx1aRi/nUmckzbMS7Q9vJPp9r
iQTmSs+qp9FbzS7aVu7u40TPXnyINk7Ta8RJeBS24MI0Hy+1lcBUtJCYDjP8N6lk
CBhNoqnezxmYqzYF0VBOIQMPVG93eh28B3siSoQHGmPxLOjW3kd7+sPsEOErtase
FcJ6ZauwSBtQDHSQ5jWUJe7PG97lW3Ewco9X/7GGo2InO0by89cZOHAX13rRuXHZ
QP1pTgfQywC3hahJHVMTcIf/fW1JxVYu3vaSIKpUdJOGm1yelYZIfpulTJZUySF1
vUVKRlMVxllGnl1vC6bcOa/VI74p12soBVwDGnPqoji+nyRGqN0bS/ytuIib3GB0
tYd09jEyb03Y7HK1atxa4HNm4lZUHSy76ORvY90L3uJ+u9CvzTkJpQhUXWa5Jcwv
W654KOtKZxQdlBDkCopCJbhPLxGMbGhEUNFMNdAnEnwNBN81r8DgI0MzqtNHPrQJ
l/eFvOt7EfaT9vwc0VbDvKgMWXzJaAj6M0DOfDBujpP7x8+pc/JJRZZ7y6oBnrLX
oopU+3dvUTFTYHhx3Tvzi5A1ECsGqRMGzPEkRLvccJpr0MS7AUTwrQnuEeA25Sca
gcwyTTmSvMHeXG+7Kpz+kVsFz11ikgasFa3gESAo4UTG8HynI6NaSX4jBMpPn5Wq
zRUTiNJTCCTy5JgOz0i1PndtD0W1Gz1xaKmmTKJbV5lFdYhuL9jdUqJj4fFSF0Qn
azb1QsvXpTBRJ5L5iP7mEG9oW/h+YmOlS61KItN2nqjsxIU3VpziGyOHrEkg6Ofe
7/d/6dpl60FXw4SgmKrvhG/w9h0S5cbstfXfQOibnHJe98lMN7JizmXOqxB7rVhj
ADPW8vgcnmdY/5dUoXibx9qMkZrwU81YzZ0Vch+gHm1A4a579UZ2srg60sx1ITGW
xoYBG9tK6BthsKqn+sV6tklpicRFLkQ2n7Y8Yze1QSLlufUyFT/oFXkFvO9sIc7V
UGup/UxiJcctFSnWsNf7zD7enfZizqi1XwU+RC8JsabnAmGyYaVozHlD4PfYbJNM
WU96KD38Kap/MeTlvLCT694Olag2xYdQR4tHFPPpJ8hlpo0ZlXeMktwrSdUIKr1V
IkHeiPyhBMa+FyQU+mtmfWk+F70I7EfaaOe/E/hi/MYGi3OKxluR5n8BZzp8KQb7
KGc20fmW7Tna/Zd5r3nQGszR/y6MMW8aJ4Vx7PoTjbNqtkOlhRGOfuZ2qAe/9gJi
FmVgO1sa+jB0GA7jFYqz7L0+bpGx/RvwbDIKVMcf7cHZ5eU1JyD+Teq7nfMtjlyE
1FtXxS3r1PlQfZ1a06iJLChuVGmv124QmUz6I6Jb22GTtU99WT5jzL6xDkKw4XFt
jiiLgLD8KtnwxqlHabAc/WKN0jJv/amtl54Kctg3NYddJPB4L5JTcenDa0pQ0nov
MRqtUJWpnbAcaxfVXBi7F9s3C31s/Z8B3UHL1zrIMl9zLNcDeMxXO0kEW0qHSydU
pnMQiLnTG+/oyd6lgLMzDxdiBPbQo2+E0zJ+Bp+42UMxfXuwiOOjV9qovprtUJ31
wk2bPxn/NONqOeRSjeErEK7QnkNHoTxpOqm3qFo7t0/eMnTME3XT3o1j7VDd5RIu
WvvX8R8TyQmJTKoRrj+GOIXYgdZ4EgKVcK9uk+Cy5gD0jkgA9D/vxQqzws2jawEo
AXz1rSMZNO1VGFpqABB3UluUNcmas2ZOG1A7YMpHee8B2lBj/RXJWCV/nmyyzYOZ
M7Au/fODy9RljJlkitLE26fei1ru9SbhRhbdq4bSpPy4waIQbp+eiJa+voRqETkc
XKlNyJ8+9a6Fky7Ii45XjR+GGnN/1khEAZMDb0hmXQmC27XDPaB40fd8OqRO4H2l
v2Mul8eiPOhEPcp/OVqt9B3U6OeoM/pA87mMklCoNC42PapVtaaht9r3VbxfISzF
mRkCoK5l9dNd2ekJ2xQ7j1MuLcASBCL/yTJOTnzF00pdAgU+Kvz6023XWbw9BDg7
TABY1dbQdvMROoE4C1NyujDfctKHAb5GcRiEkzjR+7LR7dt/QGBHTrD/xmuFSA4y
glsJQd389nV0hvDpGRSIj/DCq/Z1KpCL6wYJ3ePtQKCRp0Vna0CD8f27fKQdL6Lp
k5MwFPH3zn7Xe5AxR2vI0MD7QUm8HPHEC6eSe3razX6MsworiZJlulTtw+/94A93
VpJ4y3d0UGFTJoMunbBTnwl2xajgw+ch/PjzN2gDiKUcGP2wXmNqYzsq8xlWXjjk
B23tK+Mq+NJndQqnZwx0NBwiesxblJmZ7996f3aTyc/9BqGWjh/N1WMAErkhqwgn
7Al74pHz3Jv6G5HR89ygScFX/s5iXZerlO4jljDSiiK3K6zpVmMjXZwtOkggkpPd
uKctH/wxT2C1qIFS5W7EVYKpruCIH/GgOdmVPkqdoBwFBv1xcB4hP407sBoF8Hn2
EV+VWbyUH3uUrGb5m8XaRvSmO59zK9g0t6uLtaTnbhTb1COszK0RALIe1RRqQhpE
SJWvoxSCIb4+t/VjYOfEwZ+IAJpKN+ToaAvuSCwmZ9mD+uYTQRrQ7Nwdhi+SvtwR
KAAy49EB/bphtiKEe8ubel8eGiA41MVPCBu7bh+h7lQfdG/LRSXgBAPOqoUx9uDX
/wMy+kg7tX/Qqp8Q1plTiIHRCJhvxZX6MNj8VqGZ94GuGwkIsIRiEHmYKkxq434r
hA/gH/gky6XsVmDOMZ//qCItbDt0MeYJ3p9TOb92XKn8FyL3mATtPJqI+KuuHlnS
RXaud3IZmqT1UZpqNWj7/igPIoivKWht0nMhcC4XYD1TxhJTk6liip5FpXLPA/0f
Nj6bxP4esFlD+xwIXBStw1StvJWQX+o+hToikhjPUEzCvdvqObuFMc986LIray0O
G+VxH8Hyua3BAORaFJGhumSrSCMH1soErtwhFrPNkhbOyanPpBq+1IqRh8Q2zwx6
c07JDPiok2sEkjYng01trrXnm2gdET/3sv2gat38+xhpKYFOPLlY7eShXG0o/Tar
fWOJ77IHwZfOpxT/t68Mdz53JPu2si6ImIZWGAa+tCmLEMkepfkCjRJduYLV/xuw
ySscNqZEcxExUkHdRkQbhLVfBD0g1i2ggy3niMLR0jPUC9mt25+1fK44UZ7TcbC9
J3w/EnFZvNycIzLdh8+IKzgVhswiX7Rcj01vbfa4o3GSUvJn+I/Uv848fIeYXBoH
xgiO0rVBSTsxIAkdsnki+vtW7IWVu1Zyq9u03fiFT6CiKPEs0yMIFy5dFJMKhjam
WwXCOFff+1MEG5JIQ2g9XoKwkELu9oPFicB5meEq+jd2VhWOai9nEEgONknOjd4C
WaE0heXlO5gYA+fpG6g+xeNkp/gqxN5zh8P5wCbvKP8g1nJlrxgOLMXDqc780WSw
jDcIJEpvx6CL3yML+Oke++5vd9UdU6f7k0Qs5oW3LcWrlhugThpFGYe7vwPDz17r
ScPwwMT2FyDV3mfpdgWni4fvwILTBy4ZUhvB4fiXU3oVgEJ+D2q3R6AD6nXXtGwD
yVp64i7kFYtwg9SXItEgEroGNKwIm95pVA/ZC1CUUTqSag/ruNZRtucWaPIvYyeN
REBLKW1Fhb66hZYrREoyuR4q1uPbeGRj4dEbEsIdtwDjN1iudT3aqQjW290Ge3L7
vmIhyqrrznT2T8XFBfnIYduACM16mOrknR6frSbqXv3kwiwAQPkqHB/U32GPpO0L
ZwBr2lX0JMDwHDorWesHFqthBNXE2X0nybMWH06scyF3BbBj4B0e8KQDqZ2tPqGf
Ia5a+grD5OjSUvw0s6k5aeA85taorML2tl16X9N6+t3bkSd9QAQ8ehj5d//yzs1o
GZ/47eVybzJVrzbfbrI8T+1qggBlgHFOkIT5x/Sg24//xYHhdP+Z54xr6N2JSzUE
7jJc1OhhjpQbDUxXJ+XiijKJMLw7lV5U+gZJPe7u5SUVRTeblTB9vOqdfbkF3g1p
2GRaUSLRnTn/QBdBWuZGrtSWcQpapwkRmnddOdu8lPoYEANvFummYLUr63UBuiEB
shq/mNQ9Sxajwt18EQHAp/u6TNQxCIBreE5KyomG4NzQp79vvrtNWEPGGduxiEXE
EGw4r0hXwf85Ne8GlR15R6gAVx50yhyzDi5RU7laYBdGRgMRJ4rrjmJaWNU8oP3V
i+lMedmGmlRc3H3FwCeK3pxiR1+caKHxFrVg1bx/GvqTpmHoMyu16DoBkIqnqei5
wo3ml0vShTQw06lbZPvfNNLNpsHu2rtJngBDsmrPaMDiIkDTPRdMO5kR+Om1iJe2
flPbVyZ9Wqf7G4vvCnnNXy8WaReZqYDNsn3WcYqTci1Oum476VRt0rzN8moKhrrC
p2kcD6adJwuTf9Z7madVHspAQsmBheVSJazxkp5BoFrvzQw9FAe0hP+o8Jxt5QJF
D2xkrgP+S5H2FpInNI6MY2f2/yF1M5twGY6tk9hCna4og5aOapPnxvpVF9/D0UTq
sKaFb1CJshEo8GehH7qxHYSaXyjPepp5zNgOA+F+z+qEo/iOKkKljmnzH1e79mI7
SzAD3wTwaugbs1D6n4wUw69riFzk1xGcjjlxmSdaDChmUcQOC4n3I2BM1quefIj3
OiGII0pLqLxHEM/9TIdHEF8PuYTYLj00zqyfQahh1c5fjWJdLuz1QAiuUYVOpFlo
4zeRmftaB/+NlDgvnoorP8gJM1LqYiaNrCnXdPa7hTmIfPIbXw5Uy1F/3HS1MYs2
OXhH6uSH1OejCJuWw+5y520PKNDv5r3ZAuRnnPpyONjeYrrpbFrGo5GBs3HEdRbo
g48nStFXoZAoYPZA1pAxJ7IN/3RG+awv9arVezbngo1JaZhhL+D2Zk5vF/iYHYDp
ntKag0L4LrL3r2dWEx37uUVppKBgytRc8PJ3bq8GodkHZVj1SBgFzPjyYhM7uD9B
F2C5sYRhfFy69r9g5DKe6P57aNqTwaOxojTfHhpqGuLywxGWV995jBpdjm7fg2v7
lO/hgwBAnMQsU7cuzJXGoytyITSKDyVtCZcaxCmxwX3qya0IhyMTibmb4KTVM87Z
gRhCDG056+dbJPNLwXWuB8JC/+/XApa853FijitIhIFYPL+ozqVhE67VvmjNxU2E
wG4folLQLiQrpt56maadIoj+ZNrtlFlVJehvpJbEm0vLpBRFhGr0Qolm39FTNFhW
SdtFzsXg3Y7WJfJwYMuo44+5QPyQ+mcdRsFJE4g+Dc7nU566kOTxhMosJpcIRCzu
bjEU4O6R1tPcJdgipOGANaPtWTKTXOIoBEvOmXCZ37preV9a+v/HY90fhJSQw5Vn
Fcmukd/+MXan5D/9kdHRWMpTbYUF2IbxByZd/HZa7fqGdDB8u1e3y5KxLwt4tRWR
D8zFHaGpDKDe4Ombh1oazhRl38PyKlMPnF4UmAsSreX425H9fzkqou3DBwRehSaa
SGYhwDMv6JpLAUa5Dm/tkRIQiVp9IeKXlJilSktvMKo0/wsNIUxge8L9vCDwZG9E
mUwZtQcR7Vx5bFJiOntySnybPb2a0dsulMyKCEt1tVjZ7dPll1hOXP8o8+qrBfjj
ZOngb0Saj412WJOahvS+BhZ0kud0NFEo78vvJBAdeSEeGWIRNM2goWdjqplyjprm
7VGWpMVktAO4bcqys4Ggoc72FqNPykAoJ9aQupEKSlMCtvxI/opNYt6XPTx3SMEV
WMTeQafINRRBhm+OfaWrbOeISJRsZKo1qv7PZZ+qtyJoTsdadC9qgM9IpewOuZ0L
jUUePTVykm34Z3zU1BsCpSE/7C8r0r9mArz13DNl2i2/PPrMnc3IMT9n8KPbtaw8
9fHUsJB5rGlLC0VpyQgt5YPkIQdjMgaddX9QrxoR1Al/WbQdNCRKZAZZUOZVRvzT
8hBVyYW7sGV8/RuP8dD2MfqIFRqSywHIDHHp3PhZ0Shkj52ZcTX+aV/l5EB9GCBJ
BVOkQ/CLnZ1GOi/5Wy2gEJn8HlCu+DRWuOyA9GflVQLdW7w34/TWDpgaDMTv47nY
5RYG6fDrCk7CVYNzSpKYqEpAuhG749u4piAW3yPVQYIPZK0aSMBHrzRpA8BsNYFn
S9yWv1mmOmey8etVCeGCOoYXeGBQZV1sQ+0Kte5/M6aodm1CkPTZZdwtVSg/+yMg
EmbuMUV3MxDCh+seFJ2zjUe74S2k0yfZeOq+8DeQ/nZF5f4xcfRctvk3ev8l4mVo
qVT80luG6ZnLjlOG/nsh/s6k5lT3lUSqSOBGNsHfufAk9nFQ5gCJRe/vk4xorl0U
UT8tg1nLhsazninE3p9RnVyqXYRgGZ9XRedtBOGA3idO6BhqSejsrf8enfJ5jAy4
N+ty6St7oUCs73E8op7BtRt9Y6p0/joJ1BRVDcxS8IyVU/2EgVKuZQCGoOKF4epR
ze7lhf0laVblp5Pq/0ISzY6px3sUryPUNT56HbQ5yZkU117DwDYivltYk//PW4yY
/UhemJnj3+4rVT7n5m+SGMMH5xsLYIn3A96Mz1jyFPq8Xn+rCcHZ4wbDPclStmQq
lisOM2EDErOhB04jRCGzwK98rq96vN9bOigFMKsSTSatdUkUPqeRFzcAOVvlZhWo
bqsR+jZkvyjYI5xKop6hmweGCdbJzloH2bXf8fZIXcCQiBmkrDTsCgvB18+FSMAk
weXFRTEj6F7Xnhw927Sqqj8qPn8TSCb90BQI6aspGLOE57acUeOhhDljHWVLGHUq
Fw+KkE/5xYQO96ndHbAqYGbVTpv9rHHtAOJ6MW1BA5AOl4xKu7mt7tDXgwSVSQ8U
x1gTsU2iP7Uw6m5LYoPapDJsjBkDiO+3Gw25mP4sCzLjRVVkS6YbICUgecmgqC1D
A5TRlq46aDKKNjoHPQG5Chgj1k2oZxoUWvgTw9IRyoGJukMt3/oiLhmTrQtuskEs
YFQiXds55QozF2Mc0DvFp3V7QMASvM48FoSeuQqdT7a8K3BTELchxRbYH9ySOyYR
ozWNQLIcwU2Hgr4yA2620JtZ0aF6tMZwOMrZ3UH+y3sYsCzBJam3Z6j50R5sI/6p
emZt58nEZNZ0bTB7DIDD323G1xzcySb1iDHHL0u6bUZZzjvpGIhcsJigI1dzI/e0
42a/DzOvRBfJje0MAkEjRcMMlib5d4rosm2G7VtvMWW9Iwu4nkykr8SZ7tPN2lT2
G8eFgknm1qqRhKhurgr0TVlqssk3Dqx2GMvJZLvDdrY4ooy7lPJrEAIIfbk7xJhL
4gXkoqjXSClmuXeGk/m5dpnj5QZH6Zu+gI2YwIS9kAj7QR7cCiJZgzI3oKZy6cda
/FQ6tybcmay+Pw4B1gx8vTs8tBd7daU/Ia7N1w6+TsOGaL/0ot0H7eaM86wGzvHf
d10Zh2n8K0XKLulp7vuPaor6BWUmnzu6Iq4UesLXDJ71MyWDcnhMMxjwR+8zlJVh
/Gy+OPlRfO7kZwSE17SityxXgkXfVyKZxTOtIXmQoq+BpjEGoYC2n4DB3Q65CUT1
kjy7HypxTFZ1OGPCum5i6ceWyzsBPVeO3guWHNW/OioF/aUQJ9Gl8LcxX1ZOuofr
vxNQw45XSt7Yj94IFxGQkiz5C4eIVJ6XEUKhZmyqa+UOGpG2Z6277XAtTvXKlE1Y
qAluWfeW2JbDO1Iy4uv1xZE5LGRj1ORzToei7tcpmFIQFpDktvwrdemLwP2q6Api
TpEdIcIxOEsxGl6PH++fuI39rsLmgsR3Ebn3JQDcRQLTfctj4LuNJqzDawnED6yb
w6hMhB98c5YOAlnRSSux89bAoOfaoJPznbbIwRt343QQvLQCnZQcHm1LRRqHsf1g
nKttpFFdf3nIKRLRsOYjvSSzSEVs7CFCIKEjimNT5SAv5tgbBypgn1bYU4j8+XPH
kKgsUy2Zxk+mvsJf/wDmYGiElM+jvftgWE8Am22SquP0pAjnbtrMAt64Y8vlNhPN
zJoJE4UEB+kL/MBYm4XPGz6dJRFAXmXUA9i51frOPLA6r05cerOXuDB0eBVOqCyO
z8SsiUmuUCWBrn91KZIa8SoZGGPFCiNQObBdF6INIs54JH7UyNi4IJ3cpI0UKZI/
98J6WX//kz+bgtGVqibyUzSarZjFIwk/SKwtyjR1uf4dAE7NDW1+dPlmnPOaPoSZ
1Pmyr47baq17SgR2514OYQZBIgx5xDrN1y3BTudeJy2WMcISxAghdklOjBs3bc1g
35pXK5x/DH+joWgYeR+4vhgzwVHADbjGdtmyFYVjHL+voOSNahzVUopRuVswU7G4
lFvfJbAhRGFT86DO6syD+gBvnx7dso5d7xxtpdYeyet+QzXMSdLsoO9DuNg2B8RG
lpfsrskQfwp4PC34pnR35DYLmIUTTTtOVYaEY6omT/IOKi/S090CWnv4sHA7p5DA
hS7X7WB5dMv+9gwhKnaft/yvcXBNCB0PMJa2+Ql+pl+4HV7lYfPlOmXaG/JqFSBG
xPE6Bb3nqwXxpsRz9AOpSXyZpa7JWUdCBSjA75xjPM3ysVLU7rIBi9we6ii8ungj
PwzTNmTRbGBkrp0dkdLmc1BMJy1VJalvGeg0pvT6jS/a5PaiDLAs8Xpd5C8P0f5l
aCEYb+qDJmM4uH+sZeL8v6rR06T3v6xgovNwi+P5rTfSJMetMqNsxC3mBU/ROHVS
NRhxeM3lWW1Lrmdg3VGx80h2+lC7RY0fFcgeLTPGUZrcxZeEVJHKw5cL5t11Vszk
tYQc6jg0eHdFr9EqsCYjuLKZTTW7MC9+FtqJ1SEPwt1HgvBIThRzqqtsgItQyUb/
Am/qABNyaLUsxJrNKM6Ocfcp8607QwTmpNWFJrPPg8U//a+xyLEGeRNPHA+b3eEE
+DGJERuJP/x39cgCDyI6K8J+Sn1IQlq4kQ3V2Jt7cwSu0XmuGecf925p3IwDHCAs
e4Dd0DCeyFbDXyOSAsHiigZXi9FooV7u4PMJ3k5+81bHAgCbO3knRVhsYn6LpKmq
/R7WlISDWx7i8y+zmhwDNuDe1/ggVyI636w4W2Z3ij5CiwPgl/3kqJdqW8dH6WNH
8A5V7Qad8hNMX6pWGl1EM5NWfPnm7GiwbG+F9BlG4eJa9MQBPoowMVHeylBx9UL+
NmEYrJOyBHhI2HjQPU01UjfigM7/WfDl7Wb5Q0yzvuQNkzQcBO/mEfkMPoWV7IfF
cWQXUSJU/2d5n1x/Sv6WMJ+xY8MlFxIYZhNbtPXVBtK6AZxJp/jMEJ6B4rb04xQP
dNIrovNFlG9XBaweZwA9svtge2NTSemdR9YM9UXl1Es5mescM5crMVfI/LBnvOQz
J+94fRylKQ4cXV53VVlSrEQlmMYhVDlSJLXWkDKAzOXHVmdjNdqQBVpiQdE3b82/
VKaO+Vyb3otcMmXjjEahW4CVg0K5olzSLl8UT+yI5eMr8vr9r9ttWqTU1LNj00iu
O1FEv5hXcv7VeEt+dpeYxi9NLDGWPAja1hohHafPpvF1OyfZ9WGHgTAOKGpE0MxH
1k0HTV+tZkzN+/kU1dVMd01oW9mI0IeTi7ln7bBTX25nZ5Io9sO7sOI9R8DT6rOf
2WmQ7UDqA1qus1v6AAAXYtMlVeOo9bDIA9X4l0o8vjgRwSkkluV0GQYXDai9IFJc
kYIHCr5wb2p8HlcFZNZSvrMQdPio4Lv9GqKCO8/lMKdWRAFRY1GvX+zz5NifhHbI
rKnFSZtnR4zSEGbEdTtIHaZel9doyTOb7WbmI8gzu9zzcsv6kmfbECLQ43n8YLOZ
oCooKRyyYqKgfLG1OiCgjI4zbtLjHY4+ndB8GncRxP0HeMsrCQ2uDpqS/CHqkSU5
dJFNH+3IS00TAggCuG1SXQUnChP079HSNVTn8wNNYddz5JVil0w/RUwqvcZ7dIvG
oLWVuaElp9nO6n94Y6alvWgyEUfb6u/ptYT063SmEFMiwk9YLDI/+XazQ6stMx6B
nYviKOM5awzQFlK3CJ89dTLe5eKqIx4aulzO6cbeFFLSB0hNT929Xb6itbVOGEpv
KFrbj/RrW2J+/Pfj3yN9cKQ21pERo59c9GHJ4SOcR9OPwgzTvq/s+v+mo9i8rZt9
zrmo8TNMkf75QhxeeR3srAzkQRMZNn57owmaE5UwEWYa5u3aOKYrDFlmARnBX1oK
ZZxLMPDeSgBWOOLDfBGTnyd+v/nhIYSJhAoSi7KeH8QsEbQOg3JNn9dSZGYLi9cQ
CUdeykMM3rX86pvJaeGdyBlh8H3a4zYEkkShnPLUY91NcOoXtW1+/1q9wZl+m8v/
JMvwfrDSmj6BzDBPCS1raX/gI2TfMSmL6ykzGaa296vMrXS5h5paC66q5NLWQjlu
s9NJUxY3KFkZeoLz6y2v7+VECRabGa9DCqkQdiFXVClMYMPDbmiZcbYxZLr5Y0sJ
AjlY2o4NgdRw2a29PaUeiLJ5HqA5qo+5qb6AK5paTrz1cvJqOiUK9+GTo03KGAYw
XVuOzSIIDuy/7ygWhTkFyEjctInoohzF7Te36gLUTENgSCnn7j4PcfACem4vKtl0
5zT9QESriLEuKCH7NKIiJ9+nueUuTEbG4/o27SHmUwT+bwqlyVmjodQlcU4zV/MJ
jH3x+OqDvQsSgHrV9pj6DkGHlyr7RRbpO/hCANv+5r8=
>>>>>>> main
`protect end_protected