`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11232 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
mvOv0qUqD+6HYGQ6UGdqrXykTgIEicCA/Cm8maR/hyO3wB7hHJhSFFMBCL0VScvL
jc//lTbFNxlxDExcQ4ORGwVQ++3tVBsAXe+iLdQVKkcr3ieJrzBq09UmM74BLeJt
QHi+PIfDtr6HVdZu7pO4eZkx/52TE6IcTKxGKpkc9dKz+sLdg0hst15NQ3DdZJbp
/jvD1iu9unMTuwE9bm4o5kpTjdDax7HVuQDNlpIzV3U4nYAEgC9NPSMiI2q5yaaG
hQS9K8KXFjsq/IxN74tRHo3DhsO2ylpSvIu7Lib8yWsRTwtTijOu7T27dq/XwesR
WC+QOnUnT7R+LVTbO0nVrBqAkNW2A4Wvqhd3s4AObnpkJHFO8HouGt0nClkVHCp2
l0LKEoUy5w2WZuRxpIGM8OeeavS0zzs7cHwtu/MBJotwZ3Obe3Wo54SLgWrq/Oti
+4pWt1Awj6RCI+jMh4gSjSjmLCaPrQJrBOlCIN5nJMtVHb8KhFsxHZt8inyB4b+H
/K7rrsJOT+tvtA8DWJe5lzZDUA0+lBPSKXBNXzUaML+pcnbvMYAR1GKlPjpJs3u4
D+nWtOMmQTJgnejx5NrdUB1iKNGh04vo+5ynOtQfIG6y1V+KilAzF2Wh0GSgBLTf
fIPZ5Wn1PyjsRRwQPFtLnbXOpeZURBJgULJJQSfC0UWig0GZoxecXJ0EdRweqtOV
dd55QwykvRRQXr3wwGH1b0Bljc0VyELMfMyjhD4BgrzojoHf96J/CsGzDicFQqoV
C+5Q8qsUMLMCvCdNUOzWDvqzZIKKRhcHxpfbX3LepPcymb2/QMMA+vIuIeUQCs4D
TZxHmj3LTQgLAw0E8DADYvGpJxYCN05LzrYgCOtEfJHuBPJ+s31/UYmqg1cS/fZM
a/GxoGEU4izBPuWOYnAKqByJ9ZxB4CwDviiiKuR3gq0dfsqQk9/P/qgLTUOCBkzE
TI/rgjKWGg7yckdzsLADDsMGbpqyX4GTGBGJlT1ebMBSD4ltvDSoZh/g6sP2s4BE
jSM6EkdPjYzlM3UvQ33FCYRtSyd+7gxXR066TWukYfRIsyu5DkkAmeZdE8ucWbRj
EgS2dplVaZhF+uvzKLx6lPAdyVAsIK9xahp3MEqU0V58HBaHuOLtqnB3AtuPRY53
F3KGmVnQNZjbeJVQV74HmRzVtYR6okQknVttuFX90VnYIrojtX7JXib6dge/NpCc
kBebqsn/GlksNWYBZeRcbAhBqWiagQTA+NJOM8ofIDV4pYG1EysjDKeJpuXjkI6G
0iA45SrLyGehiY+8GkGSk8AxP2YkZB6XX7IqSz/rHp2KtSSeRFelplHllY4Yd8fv
XQKlOe/MisbP33+uGtfLkxjdjamMJkUmlDAAfNpwMivu/4r6jC1isQL6LK8WU8Et
GX1UA1e5mRf4Fq277AdM6/u30oVGGSE2QvKaLU/59VUnY81nIGcjCxdZGz3dlzEf
TKXfXKehlkyQKT/rcWBPNWSn5aQYIPC43GIufnBwSfMJDs3SAlpRZ6v/25cIzNnq
mGZYV2lnq7aeOk7zjbtqa6UC3wMN4lAqGGXv7V6Frk5mlvUJa2r1IxJ+Slar8I9Q
q/g38Rr3ssXXx16DNZeIdLeBb/j8X9Wrpe0S6XmxUaE/xqDLFTIFMxEmu7d8MmTy
70GqI84+n/0FkpAqOgYBhY18kqIkb4VzeFm18zYawzXoZhNZvL2BjDPNK828+L5r
tvjbVmsiMGJ8F/2Gs7SSZe/nBir0HnkzyOF+ATWB5saL8SuHXQWkppYmy27XLxCT
fAktCg28ohLsxB4SeMJ/6WbIFGMk804/9hi37Xew9fSizLAc220OwM9npp7AfaaK
9iYvHVfqJ4VI4kQAJziEo4vN/uokHLWB1gp1YzTUyARjBZCq7hjLDCEhV9U9Tpqk
XxDmUkamP8tRixRc+D6L59j7cgK3w2LOM/lVNFqcqtJmrguZXV+kDoUsdkmWzGCO
R6k7aOgNu62I9v/TRxvdv2t0ZuJMZZJxyjkQ5X3FX/Mkmnoh9khZoZtPIOIHBUKY
7UlTls1VBLHknfnIT8VDxW4QE6DwiQgK+bT1CnMSL6Bv/lBsmOy387XwxVzvojuV
3NPG06wQrwrqZYzklpe021sjHSYWsiXGWnW/Zlu+JazeUh4dpyes44bRHova1CW6
Zp7YeBxW/XyQBYqFxkl9jQIAIJKNanq+v3B9DBjAJeEwsztc3X0vbvBvZP4RqDcs
7BYtjLgqZOGepSsJ58lk/Jy0l5FpvAWvobvmNFWwCKQrnNiW3lwCDE2KOBWCy2G8
LoD5sfoNwahW/p3m1vNw45fdpIK6jL++Tw0zc+vdH2ltF3wvEhg1oAbUmTFRxMXj
fcFSPKLH+uzdohVpGGjw9nVtaFJFM6S4xQm+XWMohY7MmvK2BjkGkuZvRiqoLgni
/NGQIMnEBKeUTOLdCa1FnpkTE8eKEzHwxf5VDI8gTZQapiAHr3TsZrACP4rry8HI
3oSfDWIEBE24iwENlQOvTkxvyqmvJ2CPw68up5q2Y1cH48j6KVMAloWBcmwKekWu
BXVVJIOWM/L8JX/F2x9ZsxGKgl7ygrBv+Dl7/m4zbKotG3wBjwJ3VI81i6Ren6SD
5eRBTMyxpvG7fX2KC6aQC1rWUQcbFTymkTqx+OuQoLh3NEUmUzh0d4o//vJ/Udfi
tQe3rLDK5C+sbA0oJ1sJmNUUhuzi7HrYeicPMqNDHLS8rPbvt5V8AfMsBcgdb0+j
55HL9k/Kpli85kHVwEA08l8J9kwD2MEuatmk/H2/KWGqM0mb2Xm5GLab76g64L+P
dw52cqLJQwOeKlkWWbHAqHYjbQdcb8AbcNMkwwHj2t9hukBcrVgVYgNLnYb5+uMl
zaQmW63zLGMmibAWKHn1sOKObw5zqsjJHVoOcCYi7TUohgpWdMD9iCIItHwU6fKq
VWqsh/eRz+It5k8oKBbqJ1JZlU2aURlGBeWDthA1cJxiQdPnW8rBaPIjrqjDyoNK
XV+SWwCvjh5UWV4RWO8AuQ1vIjO0lTkEOonM0OedVWcb/GGqSZFrXcpE6VuRTgSe
LqhRFrHXgIaHVAj3D1z9KFLTkSlCNBBDiXJFqSuMwdL2SCF9y/3SQCwJ7XDA061V
m22k1talufSdBsyyNUNh2voVZhN8q3hGftwHJkihUSgngBxLiO7U8oi92u0Dm8vw
L8GnVD80huAGmPkv5Epk7zo3fiGEdvPVt24UJ8GMrpEFQHE2wpxMFGTRraWzOuv2
Pn4h5pZK0ltC4OjHm/TDhz7S2EGLVCbaNXit8A5kXUEC1CQocI710Pi0nMFhRh0q
Rhn8jcYauKTk8uuo+Tq9VM2KPY5uD1ta+EtFwRSAvWp925j0HHqPvdfcX4Lvo58k
nAfST6PwBv4rUXLpRZAN3jaF5kwfcf+pjeOQfgP1N2kHlaq4wLT8CvzkmQ/nZKSx
/6qKQPYUoIvNh7yAyir0eJMDLPDUTHszbZ/pjtBYnUNfLeYIelEn1xPh7LmomL5c
3fnlI48r3FfQcWsEdP3WyE7AwceFXf5PLRHGTztn9pvR2G0WOxuVYUK3KHFeY/WP
sffJU/yu7tM/Vvt6jd9/lG+GXtlKex5UrEBbm5WXDWOwomGAkWC/7RtltajA/OVi
fpOlMJ3PTIa6/h/dfBv+xqdeQ2dE6AZQSr7qLuWCroRkirAQo/WTWk+RARUYXvTq
UEDw2uK82VgMTuYv5JHoSsOxeSEq3Lz6av8SXC0A06Tpg1lGOxXCWRGE2MMBExJl
2DWArYOdCAHZJnhXgqROt0s2bsodPptQAor00BlFfAL78bOukYCJQNw/ZjVFxDBM
VRStTKgoNSeLeIxiKLecbh1RKqr8fL6IpEENfbM8MIViXPxnEUpf5FYZddyrXM20
yKEF+Y7OqQKaJjMAxqteS7SmBXHU0KO5qnOwEPPGZr7ES2lW+S0AcL+f/84dofyp
vRjvY8WM+1C+frPDhdW7Tr09T8TVu+TZ+gQdmTtsrRm0skVpkPUyWFYahRi7gT2j
Em4zJ+S2Rqmx2RCdxVP5AgSiKP/iVMDfvzAp4/j81y0azpA7OLuA/agqcYQqyuCO
8o4UUdW+FUYveQmt8NkO5xJpysERD/Y5jWH22H/yvdBreSiVNFgqyYCz7USypgQd
xeWfTL+p/wZN/VKWUEZhicWb0o/RZYuNR00udYxTPxnB2j81T4JUvouo3HaZnkfj
7ZcKmUsIUZlio+OakrfTaVpaZm4hU+k3UvGtd7aZ/ZN+quFDkD+UW5XkOLcXI9Qh
TnIkATzlLvx/oFP01kvPpYMYualRAwEVj/JLwzH3l8xTYqvMWWzn46BJdtQGxQ+u
Em5wt5/iI7tetx7I55st29xQYuV+S4lXqS8SjzmdVzmqRDSAHbqgspfem7RY/38A
YmrsZiAyPtohtK8x8yGFIoAAvwqa3qHCv2rxq7StRmLgoOwJH5+EF7f5ybsX/Rxd
O5rZNAFyAFskl4AXGj5+C2mcB8hrXO4bBO5AEijPbLJyl/4aJkzBaFA95iC3Mq+F
V5RHqKHfFzJuusTmmGG6DfpMhMr8IGLdgwIX6kqbDIIHan/fv4S0spZKffQ/gsPx
wht9izgKqjCgPC7lQxJPG6l8mD9DOYczk9toe0evW4/tU2IA/TcbtlxMoAc1KdEA
nYvievQF0GHM7+Vb7RJYm2UmRwuO4RvE6mAxH5spsdMCPqV+QQAApKr6ZQ//UFX/
ZIc253hxOzGh1cS9E4KLwFHgztDT+fLV3nV8J2rBbiqPWi9SwcXRrHz0tsOidsv2
CnV0fBsR6rObqKO0iLI+m7pl9h3X82hN8r4+G8jQXfxtBo6l3/vCZxETXQxCB5zu
ATBlIRTT22RntyWE3MmbmgKKGiVC0ZfxakXzL0vj7u6d+EAcNdno+zNqHMqcw1O3
zzKFdhljpVbJ7OehGXBp0OVepA7o4zOOvLtuiuxyi8Sg8ffIzuBvamLjgtNXxWMo
U3F3sTsb1n0aSe+aYUj6s5xvXrMCMaLOcO38NBSuUZaVEru+VFz+cLpu0EixzQEF
SxajOBEf0tnfFS29Yef8LBwoxAndEQb+zEbZ4aJypqaIoH+VG8IMg2RlALpXnxhS
Jo59aAIKuhwpTgOWkCwVK8fY2KESP8X4idwSsRdWkmL0zSfeicsPrqzj2l01YzHF
8/sPM25ktFXwL5HSB6p04KYF71ER38rmBD+HylSfzGBF3XGjgP55Pbe30YS2T/mY
0tgjetutqujOjir7Lo1on8ue4180f/8/ewJcM9G4+/M6x/MZiz6Rq4yueztUSs+9
TCFnh7yFGLi2o4THqLyQt8nW1LtjMOGURvw0cGxfJqR77esYhsYh5J/S2BdwBbDR
3WeTNc77uR4xDMH6C5hIUwmNivJH+E9whyN8105KGHgJ4R+sHFW+BfGe9NXTG1PN
1SuJXfv10atxa/WNdIXFPXmCA2lBTGheVX7nny0fCtaXT075N8H31uQww+ZtXe2I
sYmuPtMfzxut8TVg0e5zXctmZwtdcNeicA8O1ct6+eX2aCYmQBEW3rJ5LyVjQzKT
xHl8p0/YAXuHgddz2Z5FfkXJifzOcdj/VqMWmotU7JYG0BtalfaLS6rc9BKlkpyZ
RK4QogA2Br4B3ExG4VM6axQzpS/xpejWGI1gcGPO/vziBRyDflVEYqaeuirZzpcH
RhiZY3sYLXIBww7ujP99Kna62WjQD5xF4IFfas+r+C+Iv8bfkPPG9Q3h2jhcfMH4
Wir9zmMhXtm8IRGAuLp6AfPTvabsYfXt3rmo6aAfVTJxypZB25yjKnc2/WV7/2cK
/iaz2hoEsdTPW4PURxqMmlCnDTZImnCxnxwf9WaONFe+pVHeCBH9coXqqvD27Y2o
g85bY83kKHUf9Lg+aOkwjCsa8QJMiNvv5wz6PN7cx+5xWCNscUHaeVUqazlreV8t
wL4pRJGp0JiJNcXb1ecw6CCwQtVcycZCB1NzRgaQhqyAod4QDFJYLaXDznjz48Bn
gFTyLRt993wpppLUaSa5pyLbF3vvkWaWLjhdXejaKhtWxSC5zS9493g5fZvhcPcA
qK+lkdF7xgL53B00nJO8+Etwt8CEVHf2LtpLhpLmZx7aSFKGOP6tlO8f8k7PyQNM
s52s0NO0Fm+tPRPi2n+4EDAhSGLHldITDP74eF8essDl7LMAN6B40j2lUrnaBMXo
jyMWly5zpP9sSW/LqF0fpfktpJn1XvAIDIe0eVkBfqgfjoqkgBiyrFguGgY/JH9q
ogUAWLnh4bEnCRXMx/HYXT+ERewrWAutb74bopu1S1DkJiP5Xazll07i9XctndLA
NScQRQPIeEVKK2jJMuYjgLZXKOelGxMy+rxS8d+1XKLsqAPq8D0dMxL1XQNPvLey
nP5k9NBvwvnF1jT2IpiUsno/I0iAZwpkXhFIN/FMnv4CV5PY/Go/raj/UtRB+Ffv
AmLCZYNmwAn8lYBJ7kpHfz/qKxZakn8SS2Tb8kyIOTItnkS24VVt6IUT1EG8q8tT
eXBAIaw/rQ+1gJJOrjynZ6NYHaG8Wc8EAttgDWVZZM7eA/p3l18yrA7mJ6CZrHIy
7dmjJqDDrjpQgijFmqOrD5feLaWmNdUosWFirHXHU36wQU63+yuH7uH4mYsgXxKg
y/DwSw9FbJbYMIB4SRSnjNm/GEua8d8x482yRYJQ86Vs8vkBpXl2NP1k7uoKetuf
ZFwooR1MW2SZOFoRxXRgpD2YJV338mzx6Tl0lEHUUdOnHs/tK6tZ6k527FImZhED
bjfL9dA0w3rDQSoHj/IiA/+9N8rBZWvuiS3VjD021hzDwfamuBk1uKUMURUaHT9i
YAZ8xPKLUxDKShAfwUeuKX/5rRffl419KjsQ0m0Vt5mNVOY+z8UMvvl3gvFqdxtS
xhsanhdlIQtoL4nybOd8xTdDzwtnmF5U+IeMqqLa1Ssorvsoa5/B8roAoly3k+iA
2mVr2cuhEr9o+vfsNlWxZmzsgCWRy9DafrKlrsBr9y7+eYESJSg61Lc/X6mDmrER
U+lMeX2KyGq/Bqk4eS0jbkOJy3c6aOHO20YWV07eZa8uW9lRtpDXNKqAx6XHabip
+vCMU7kdauQSAzBsO41yxuw/3aP/FX4j8CvjYsvzN2cZSh0sZsQjYUZudLeJxsy3
ZNuraR/slx3bP68NOfZO7NHA++gnSmJMdmU5dpr0lHuwrqga3kT1UNlcqInR1s8G
j6VUMS3TjOGiktGN7W8ZGASP3TB66wqA/5cAfACRhebRAXyFIrgNJiWh2ZO8u0uH
A+2NqQG9oq/zXB8vfBgsSWYGn1oRvMvxSOq821ZrYBGhVqebWakT4IX+Ua70DEB9
mFpvb9LL9v1OM/kMwzARccwayVhmqMPxj6lWm/1QKewDQ10DMEyO+9fzngdheguL
lxQ6DIXncBuW12vWl3zXA/AiPOW89FRMIeV9pc+g94luIAA0tXbpEMHaXB90uFWk
NwjpfTOHpjbY96xTTMivE06GlBWc5ZFqzKgNdYktZnpbzm5FXpuf5hkFj+Cb3koz
OBjhBwf1gisn4uDPeCB0G6M7+cXTeJxU9YyjVgU67t9WWxfomwaWTS0HdPLG1euP
6JpsHHTRaUbUAKwFJR2ytXW1imudH87A+s25wn08eTrWjRTaKC0/v4GqmFpclfJ1
67JqXad1FuoR3eteKNvSjH23wOzVnAonWTSvm0KIhUnF0jMFC7H4k7jrkKQLMoIx
A3Mm9i4F1NvatafcjQACHw7wLwH/21iLps60/OEXCYAuLxhEh1lrVyRYxsakIUy3
g2OYGH10AHl0bsuxKieODSxLrLsqiqhyDluoGQ5M8dxIhSAvXZjeSkvxL66LSAHo
S+UEt6NN4/7XdeJtpNmhOr5/7m7Si0bYG5aB5S4b2gRpA005vlAGlPpQLf9eJWim
ORqQ6xv1/yStpsYA+QKEr8MoDPo1jMHfzdsZqn3oVDQbm12pnXdNvQ7HXKNmDEYF
o0X8N0eeGadLtq4mf9ENL+OH4gF9jRr0Vh4/lR7kJLiMBUPEjljAHqGS3PZMndBQ
MIRsCoTdoUkbIVZqwuxF3ApEiZjzs/pb19EF8QfrHO4bOOIi41djZRm9dfMjQfkJ
DawCv+y44O6xyMAx7c4IDbJOLihrg1RHB73zpNLK6XvTJuqpn3w41Ip8+KinPQIv
vwz/wIf7+I3HDa2gpKDFXRMNcGOX9NvpXRDt8Xb3gS31hMAxiHp9naZ4Z3os4WmD
/5qhy2EqwB16LOTqst70xdZEBXBAqvZYhbXVG65yAN2qVph4aPUk0xPtideaxOjS
30aeLTbJOHf2WYqO2V3yByPKgWofC6MQ+QCIDEfDVGLyZxyTEBsaRWqLLhu1+86S
CNlrvJTUSRFboRnl33IFLYAwLBzjVH5iHpnZU1BRezcChxoAoJyhuv7vUldbVsa4
fjMSYmGpK/bg2bHS9Cm1FXG5nprzH0oi3nGjxH1iC8gYgrhsgnA9ZSvNndfNM624
JzR3L13iXVQAWnri66I6LClpi2tM/bqQTgF+5EnG8ypKPl81NaYygamoP9k6YJLV
Q88Q33EqpPpwXLA2McPeHQMdjv7CV50XIilAlCByWvQMP1jugnT04IKXMrCOQLCe
incrQOO+V29TqEdpbS+WK75uJWnSgg9w2yN6kPzMuL4q0SQcnqc5inIqs0d9+Fzh
qu7zOdfOARyyp0G4SZHIv0dGsp9OdfA6gAg2Wmu7zY6sLpMKVMLhcprMK1ey32eQ
qzTaWWCJKfBYfYleFqNHlfYSuOnlIPgM4KpnUhgBh837OL1A7UhF/9nY+L1JGlto
XMelrWhI4XX+3/X/U9lfG+UBC3n7E2wofo20hzKzuvJg09leXyPlAKFhlLgPZ3eR
SzxBRUFxzHxXbrekixtPHiEWub+uuybk91rjzH/m+uTU9LnyRo8aSn9L8XocA+g+
GwXVT1yQGcdqe8Fv0goXRoXGU540sWAzEt4ZDX+02NKbaahjzye8OzM4gjH8952G
7YfuzGyV+LjQHLtdsUnpmZBbzKeH5sTv74EvTemQDeSMO5MH82GN4QjCVZT6O45/
ZnnmEfwgCwOJ9xyTKjGdQuIq+ZqmTapVI7pMPLSZAOpSm+Q1zPy9L8sXhrqCWWUi
/ELU/gDAhoN9BFxeRI70imlnpdYCG2wdCw83B4aZFRoi8NgTcv+1KVYvZaMXev92
8ZUfDgnfyiUKLZrgXT2t4/bdT4l3WduZjwfQQYwix0i67pf7mpuzg4JHT/JAJDyd
J7tnrCbG03cVee3b4uLcftXXKMnbpwOF0s3HpuY1cxPElxmp23OQbWhU5p7jjDSX
Z9mXFETdpHAYigHqPV+uwaCUlj58FdHbnoxBs+L9ULKgjJizgKJwn+10g4vd2zGR
6LZ+Nih3Aer29opDLOI8OF3R4bdCsdftpD1LDmgT92PDDhKspMhNfeA8VvaCSMAG
UnggKNAgvL2zcwL+4YNYhQB4eybKvWwEQfsCDK5pypO3Hnc0u/m+ozCzwcRL7Ti5
KlJCxMxPGtaMFqMP8zTcr7RC6YxWZ0ilEqIGZKFsvGBk2Gh93VygoFBugi6Wk9Zg
Zy5O4Uz41Vo5aaKNGFfNM48eHofZ5X8XbmoXe3VeXqQd3igAE7r39awudTHMwSOF
BhQmndkUIQKrX/y5D7QMwmonhGCYp1HPxCFoGnMeKvyvpLU0loWkp69PEjlm7EcR
FsQI0LQcHOZiuyesvet25OGVCYPM6NdS2vL6nvR+nSI3jL/FbUFpTpzOKy+haTx0
SvcEeKPPVbw9MwvNg8qfNKT1e/W9IEfd993nxUXO7DoVg/bj0+7g4FuI2Uygb/aa
cwhtT6I9fHuqI9873VT302yK9rppNvYDwz3QOAJWPn7gmdAJD9sTN+Czg240KeMT
Z+K7A9yes7CuaX8iAIrNZHQg6umL8lOFryKpiGnteR68GSHfpnXf/QmGFOpXSzd6
BU1IhNCryiyBbWPRHYKETYRgLRcGTgXr+hZ5uOmmp16zkNxYMyNyLEYpps6uBfjs
2vBKZyDFP5vC4/866dv1A/qY4/k/w31a7LZ361cnP9huwCJss9knQR4NQGWFOhsa
ejnS7cu4zgd8p4DHXsqUM6cutFjluO0xlEa+4Lzyk+KdNXwh/w7vf2RJrIrBkk9V
HANYTrh5AcgRpPR2QHXMgIkKknLQjKndx6HO5KirP9rYLIZz15qawLKH4AfByZYY
rqLQ09FErn/REq00+qQ8PNFJalW7He33TN2vn20knO0we4ZdcpTcaNvVUQGAyfU9
gQ3MJYP9qa/37AH/DNgmoL+H1ze9Bpues2sxy6mf/FDoiQUhJXxGiv6MsPvuYG1g
Q3tAkshVfayv5DjVwkQJYt5Bcu4Avew4P6oGmagb37XKTzrt0OFyrmwskhZednF0
F3j9VufZCZUl83L+YarcXrnFINJovhPdHGzja/BbHrEi1uB6EIUDcL8Y4FZxcD4P
+YTDnKzIiagMYh5rTdhu5BQ8QI/XVvWUsNTyyrt51QbmGsS3FOEm3oT/TA0OdH3N
WTsBzTH/WwVFEWQwR/48A2EKATCGTjLAnWEgKAn2LIcqw+CVm5640+Xn3S4t1OBD
5FGjTvWWLn76YvMohHsxjCw8MHk5swF7Ad5HmxgisI6AVYLuqczMo95/buZUiWET
GWSmkU1HKhS4HhCY65nUxQpIXXYj8B6623K3GzIaCRm+cb6Ajim0I63w39HUVwvF
p0nvJHTAvNanTE3k9Pg/REvJKK4SwZGKdsNF5pgVbj3wVrtbMH9cpUQGlbIEpVDP
ot0rAmShipUKUhIXGfoALkA+aFdcYRpt44ieWrBtfQAplmadRx+gzXxmcS+eaRxM
q6WZFKwmAEBqe5rDM3o3QwrgeVVejXqbqgHYZ5yGctiQKPB0TXs/QIdynCotcOl4
7sB8/ZlEaqozZ+9UzhX5OYQuxKUpUCgPUPw8ZFiDgfNGrir3nZKbSU67azs+IzJz
H/SAGnth6b/reTQbho0gxsYGN2sOaYK8c/qq7wRqwvSyG+9ChUkA+y0ry19s8Shy
i5EStnOBMaF+F7mgWKIHBSrzElX/XXx5u8gbzgH6sykxjPR4aLUVoETl78QCgEbM
0E1DJtNiDigi1TyoBQGwysJpetwhQjFKL4QX39eg7gN9TiFpJ64THhs3k6OmOuwa
10x373Ezq0nmeJR5tgL3I5obB6ns8toEDBV0GGRfPhcqFhHTSNEudG9Zqg5tFt8f
uR0rTknVHnJ7Z+Cw4dgFq7dWKR12QE76WTWj1EaqNQlLwbAw0Ajr7wC6ApqJQAoC
ljgzUpv/9N2ARhQA5QW2XXCw0xJ71i7Ua4TZ5FsGZZkrWLxv1jlRUWWxSzn06POC
t5OlswfLqu/eOf4G5noiB9cRxWkdWUJrMvR6LDu5JPsApZkue2tlvJyX0udE3eQB
mR7VxAQ+QRwdfFsCS2xRaqrq0lqogqz2FsPRcqAic3mMUjLB5FWWeZ4gdC02YtqV
O0k6OHN+7CxvVCLiZGG/s8dSbrujJXmV09OOpX5QXG7IOxU5kJfWRQKgMqnyD03g
UV3qafAP4Kh1TCsqbzj7LGxpPBHCBP6G7+F6Hzn0gRuZT3m35L6dzIApv10+GpWC
6eBHKR9mHR+OCkgP9EdFrkJewRmtX6kN5ZoUp0oNNCgImQ6buAe+b25GfhKl6ctc
ia4nlE7ZB+P00+ERplFo56t5gcUW5EbfV6Rb6q6gLYhnONmlA7s3VjS8Zzlj/0f7
EAZdqIcSq8jRH54I65KXXUhqQGbZO7BadlE5JbrcPSoAb+GTaXAlAKWCSa2W0IxJ
LcUeSN526I5GyBCaTBEmEktIkN5sgCBP5XTqF87rO9ohaKfDzA0oFBAA7lzP/76x
4itpW75ye00dxu9HcG7L7SL1d/NOuJGZHJWaNDqXU3ryoQyhLDBgWs8xU9vFypmC
Hp9mQa/J+/73zZd/ea814tEoLx9nNX/YMbtTqlFBu4vB4JTcdjOCa1Rsej0DdVz+
UndI1bFVQXRL+a4aszjwrbHte6RtX8f4sy+gsg5KFDR8XYATaUhNL4KOPnuJHgRB
lv5B95SUOPx5/TpW8trBMaFbKOsKLappqjLXVQlq1pYsTL/DqT1vKs9fvKZPUokb
AmsVQmjhaztb6hIqEzPWohAfbHNAD99y+imhke4HuWOOhMKnABDfnrXfe+s04aEN
1xTgOFtBN98gCc5nioKka7OHdRmlJMCDsR+K34Btx+TMamfLTj61oOfSoVZatwHf
odswWWhfOBjAOkrHTkT3CMNedDzYQJdj7Ap8QUPJxBFLz/bDwy2y9p8s3fOarF40
GNwZ2FpYbJnYfMgqYJMpdC8fF3EopcxTD3e+iYXoQMu60NCPVOxWKYCJWqdrU4mv
2NQRUs6O9VdZnbXTFJonuN0qkeC4bRJU694cMHvYDGY2hOrds2u3wsp51SN+S+9Y
S97MAml+b7fpxcucYDIYY3fgjSTzEbuUr4ZVyET/ZhAGcrZZ47KaBcOHCWTYkIZp
tB1BUMRdvPkjqkj7SchqZpYsZcrUXxLuaY6AKoMkNu3IHOzkmUcnOlD8lQpjZksZ
GBFgAJd0Wkc7hfqKkzKTjFEN0DEQ97+odXI23U+LRmduyWVJyElrJMs/ZOXgycg5
YNoAmu4fHaoCYB3Foxf8Wup4RyCoruIEGGu0Iha+qreGe2mGyZmInl7ZN2sx8KZ2
s3gyz2c2nxQCKpnbnGn2DsdbGRQtHRd2TyyO2k3AIMyPahdaERXWWw5khYw1qiBp
VqkEvTG6t1QHh+9eMIXUK9URYBCyZGY+MHfPVVRQ9YkzesSJTpwcEUGRkxEPYPn4
jzRr178fXg9t4LRfhzN3NKSx7dAjzSKwExBQ3K645M7Q2IFnRhb4TUF41JwKt2uK
Vxy96IRSRFOIG26CDLeJ+uzTedDclFtcRsDqRVaFcnRuD8d1a//8zXgYF4WVTi87
kGTbvvq4Cno/qvA2N3Co+ygQoj+jK+NekFrePV8w112bune33bQtzrgaLo3zkh79
j8/+bSESsieOr7JICx2OFwVDRbiJPAoSxVyGp8bA0tr1fsy8GdXnyIXRBWIn4wMv
ljw0pvBkV4qGhWV2XAedqu9wC/Kvs0LOJi9IffjSBaBh31ApQm3jiljlxLaU7smW
o37xYMOT03zqoF2MQwSFn1mS9l/QdEiyMkPZEXdwhi1+u/+SnpBnjlUF8Eq8IUjG
QEhryvUwx3nenaIooGG3A/BR4P3ZagFOv+xLGv55D4+TG2SOn44JkuPqC/PFu1S/
1qRNzR7PqxFyrpvD+gGpbWgmv/DwBH5ueyjPFdb8cpJpk3pK8+yCWpSnw8mSHLac
//zySc+/lfxlv04zarOoCJ4M4FwSEaP8CI6uU7ZxE2lAuxuC0I47nKeQKYJ39bF4
c86ZCmNyXlA8vqS3jf2Dr29HJaxaVduezuvC2fqjCHZ9RPa9CDXiepWG/AbEFQGl
O/eA/Beeo4ayMiHnoTJ7RCpEPmWxm7c5AKUTCMe5HAqOJGXPbk92krs0ujUe8LRk
ZM3w3Yl5dpYBJwqYHsqKlAt5/kcSKkhF6O6BkMd+1OQU7iLg1xa36w0dsp6d025G
8L1afunGqgfJYIczmFx6P/SqTD+okPbMgui2XoWqlKDM9X/Zf+pSg1ZJYOvs66ey
X91cTBP4ltuWe9nzGLfBUdIxGTRjp3jhyD5YgP1qMdiWQWekcyTr8EV8oXUTd1bY
ErgI6DqhnUKAVaTD3YHzhh4CB014YYLhsy932Uuyf11g9opUaxd687WYZJOm5ExI
HCpwGJAqEHX/V/7uGTaIPHo4m4VBEKssbW1DJTZ2IbDIs69456PzPrY4sbasVj7x
55bTUJcDZthV8wNYZVKhb9v8VD16HThP3ejeBzX9sC0NGY9Yt/cymolryjmuAkCh
Zooe7dFyWOmOdUPqrLDPlhSLx2d8Z+6+Mr15NeznfAQErkHfruPrsbvgGeXAxNSd
aG2xHT9p5k8/6Io77NtQdQU74uZFNSPep36YATAdLiopAz4KFkZLKULEa3keyRlB
XTAUhB4QJrEio4k8DjHuHJI+GF04sbh6+P/BD88B8Ycv1+Z7ab76hlGpu0gKc6hh
O5JFndxOKJjiUKTGXiLrGQrLqvbtaUf4Rz3W77U4Vy7kvnBDoPrJAIWyw2RolG6o
b8n4eMHAotzZarYrecT/pue8HOHHIBZ7f/IxzBVnbiVLO+MO5TadeeZxdhZtNsK2
jCMdzjR4tbev7q7iDnP+9zYN3r/R8NU98iL9M6pXujoxFK9ZDpKz/5kNX9sjCgC9
bJVTsSHEGqlrr0FXSGjrOFBCFuCTEE/kXINZMGkMkimetFrYnwQZGn+cmB2sXs4Z
MYmpYc2mMFqRPPrbpdVOea8Ap1omnwmbRjv1eThTZZJDgmZnN1rpcEFyOQN5cW1I
dml38kUNu/R91AdMNx6+s/ucJGQS2hDhqndcRGOlHbX8faWGepC5YypyamJGnR+w
C0v9wtFvhzM50zhhbueNePVB8rDZ8YJyZPimCmsCSv8rxo9U6lX1G+aA++ystM8y
zXNRUdlRGdpLDQtNoRJrVLDznEW63raiStg/OUrgWxncaCIHkikCAHnIVpP/fetA
qSgdDb9mzwmWypMVmnOFByDNhJx2FzdBhmsRV76mqZ6qSjk/BRgIOr9lgBDMygrN
NdoTO56sXTwAcOSkZuK58qCNSj3eiKMl3C2aV6lnLdzQi4KVreD871Mrri5gIhFt
jm6i5GeEUETOUpXFgZmLWAr+inRdTxMYFJ8ieVonTfq1K7xbcica6DeRSLjX4m+v
`protect end_protected