`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14608 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhBNVMbsl6PTB5/ApNH6uD+DV5N7cjkYfz/wpcmHBtutG
aGMTCOe8GY2IPU/Fh8AdItvayopufmQh+ov0cOirMkw3XqKzts4RGspwhBwWGN7N
4mSLBb/EgU7rUjh92HIIa2JpapWY52bGLNzghiT2QPwtn8HtmgZ/ddgeMc1W5xb0
Fttu2CyPkAi3a4UVMb3osVZlj5LlYe0kfYxaIFYziQLaLRWYfcV+czxd3ncO5ZM0
FAMWpLixdfpZfelwrHKTP2g+zG4kiOGjN79ueFHgFpZz4XZM3HeVaj/ON1IOVlj3
j8oqjdGp2gyLAABdKQJGqadHuOK57z6zyQ3Z4ZAUOumkMyHeQkdJtYXGKF9Y4fS6
ia9OY4e2DDmHjYbeOs8/uWzR3bqTPDg6w/7p3anYgbE8nd1QQiJThS/4IlQsAcpu
q6aJHY3ejFflQXPvPNpS7yQ/gkz1785i3oNE+Ky9sTPskcrjSearWnRsGY51/QCe
lqACo8tua1mQ1GLBBCGtt6DtYZ1cz0Ao6NyXB3/9KjpsVznmQk28SWU6WqmHeSjp
ikkfbNT2YixvUgZMS5NARRkxn7bo64oz5TfRnEGk9MIBlzFcy6iWXP9Td1UrybfO
SvtYS4ej3mVzZPL5K0VXLWjgMpSa6/Q1riXfu+YxtdtQ+xIGe7A5cdGowps7GwZr
KvgnHbJ3BOHgPj6KjV5uWF26cVF04ChggmAR63BGx5ywiFSvrNOT0bIAcwM3J8DR
mcCEO5+2vPPTnBc83/0Z/tt3Q7zAZHSpNh2MOGa4ce2fmwQ/v9LPIGtRgaIha3Zl
DN3REmR3idg+bz3fPTtdbJ/DArof+B2q5lWkupLt1GjQPvk6fItj2riBY36scdcA
5YjksVveh3FR+nP3j7X2mRrChukbcHM1pLejKcsYnBi7HY8wAmDLrrgebCyTAVq/
nkJfWgcRDQ1Jc+6QerGmzB+/5mLjl9DUWUS4x+ob5Eol0Ic3yNPXjrD8FPltOcFs
h0moMEK/iu1Esz2Oz0BWUrR05cYgKb2QUCXTi2wPWsapZ187WEA3zw9Lf3onuW0K
QQ/QLiHZO2RiRT8+0ulA+RvKiDkyulodsYBoVkWgwk2Q0Wct8uvpPwzAfd9oEWsE
H8AeCVgJ+fRGut7JEMGNX3uaz/3Pc+pBCld0P4tV+ofnngio7xBiEv4oZ9v5Nf6j
GGuAD3kU4t9xLkx9bWdNQFnz1hqXTYRy3s4Jqi2deU+CNjmL2AK9aeTTsjb5l3ts
p6eXr7gytCQbJMaNln1L7sFs9MdipLfCdoIHLzrNAVV9bRV98OsbqiOPwBab4coD
+ZwYHCgl+yBt6Vr0HXRgcPKb1N9Hjn+CLFKXPnjUswZtW3UaH3DT/413yTtp7Q+C
OMqiwHSNzdbcVfc0+yw1NRNyRyorIltXoG8fUdOO6sGv/8630i79Ci/FhvdE1l35
yHmDuDZFl2xAmL4ZZfAA5AjEauFWLGk6Mxzt+3IQPJRp2wyBaJtZHEG2yA6s+ZXa
dk/EX219lYJVq0R3+Uwmv27+Wsmq5Osp9Dv2IMJs2F3PAcqdmNsQmm3Kbpo93QY0
8JxADe/pH7dpqEbKYfBGAtlSaZtwEBP6JDqj/BU5AcYxzrJiQALZ94G40tfn3wM2
y+1YaYPuOfKqvkM7uCjUk/CRHgpErIEAYvXx9vdzy3IDMdS1Bf03ixne8zrp2gOo
yklhX2NAvYMyr5S9Ndb1jSf2FVBKm5Sq+cHGLCNl9SwwUZSTl6CBDxKkv/f2sgbz
fuQZlpYtoN0JV/nf0JViT6Z8S8+5EL1mNW/j+W5CKn+jdZtFTbew9BWWr/5xMt+h
CPRx8+26XtvWBYw2wv58YJaarZ7T0MQF54Pc5pKfAFH0jff6A1L924fPjICJ1wY6
2m393/IRKIsWR76+klCN9+d7engTDdefE/Nl/daxspUfeEpw3KT/00vmXcPuKQH7
qaL8D8dAe8e7W3XQ9460jl8BqzpYBZg66IIu9FgRl/VweHwgAlFmpf4+iKAFyz9J
9MFGVNT3MALFrrYKKKdmrPBIuu0wpWANmem1yWk4+sAsiqEzIQJCRnXtnKaxpdu/
DrhmZlxyIWac/a1bV5YX1vbghT4xykxLMd0XJNnr7+1gcZj2opouKBZd1yohGjVQ
R1XHdNUlwA2F4a5GSgBnVL3nTWbsd3dpP7w2m0pzA2IkKE0RmzIhGYPjlc6zXf6a
F3v7lCJ3+gSo2L2VvqTnXzd6yIbvuDt3n6TiUUaVi32SAyP3ad7h2AE//fi2niq3
rpOUwlkiCbfvwMVkb8qBgax++G5XHkz5MEPbTvOzyTH02rt6NNJqlEW6+yAbl2+I
lG30ckg7xWp7saBzBKcZSzs9VEOKvEiOid60XGNqsESj+TFC8iTQmvRVvToWCc70
1J+V3MrG3osmXrHlJhu9OQc71OcQ7OSqNKqwuMk7XqkLTg0Y7W42P0CxiY4LB88i
WbeyeIDBh76qM2uhjnM+J78Ft0G75SMkC11iLBciiU5qmnBYTmIecKHQpz88dcyG
AqghQRttZX95LFsJLkOYmlaWJzovrNaFV2kAtHtakzllKY3BEJZ1zJcJzjoG/RnW
j8Kqy83qxVzgBVWm/eoZ/8ebjE5PLfvCk6xMLSRJltJKv7igNv9h1ILdpH+GiB2e
0VO2ZOmdUawpNwsz1SDQYpfi0i4D3Ww3hojwEgo/tejzXOXwKk+4qdcsZWvvVCw9
c8yryhQh7yjU3TlUr9kYvOLBeaXcuzXv+h2f3py5gGMeyVda5bP94PTSdjSHroqZ
bhCzcsYNHdHFBkwKQnHfO4fCqv/j5caNTrpfLSwHLoU7HycIgfZUl5z8w3dPWwiF
z7ytaBLMjh0pjfzeuX15lTsFJrCW5i3JxyOwCIQ/awALOwKfPcgjYHarc3koI7qI
Fw0grmZr/0osZg0NU6LGkBCtMfL1uEVLMrIlfHoyML5Gbj/WF+wqHRz6uWwmpghi
RNLYjBZcY5oBwJNZcjD5QMClytG15r9gN1BLIwUIThy2U9/3Ggj2AqkjdzFRjwkD
TRkW4OgcQxb+WSbDf0+E7qUZViEy08wjDg0GJC4fSod6yvilk1VYe1z4AFoK7Yy4
g/BuIVplPWNBqGp4kvfPhe6w3xzZQSblRLxCJanGD4gh/f7Obyd544ME6linCrLT
3g6ZT2jH7Q0h6DTy91pcGqtSZCfzX02xgIUguwak2jLoUe9sJheaipi2WkkDYXK8
g6d7BGBxFg7GIdCOCeK8oHfDTr/si2WXlUYsxZD448fNNdB+YWCfwnXL91TPylNg
n/cZVoaDhNPhO/W0CqZRJqa5VTvB7EF8vrfXC1n2o8KpwtTKsXr5VmbcrD/3ipLX
iYGCCW6vUi7YFvAUgLXQquIKYGVtMtdk2kWa65zNOdyaW3SpSmc3z715uxqfJ9sT
hVgUecKALn9hkDrIVNi2d2yZ7Yq5TXn+GKhDv6+l0oTcTA/H4qI99bboo9Bm+vKL
7T+cXXU9hxOTyzqJyBwNeztR70GpC6Rr0ds1k7WgxkOv/mVl0NlXsbzvDtMoW+Bz
jI+QzMuF49hrOt/Bf1hrNFus0+aTsA5shqcuSxS0IMeFqccdDBDBktvqIZ6JJLP5
Nr4Mj7Hc/2wm65+WBSmeAKdXNSycAsaouoPFJuGlxYrLSUY9sNqKtJ1taI8p9rLx
+Nk5/I1rjN4HUdDxtaw2BP3AdtQoqBFj4e1Og8jE8m2/hVhczCvL+7fWDWFBkmM3
q8MgJBWninXir29sJR2KdYW1pOvvJKPcj4ZE/HGcjIyWEyFFVLvDaQdJUuEaXfDz
fWusyIL6c3f7qJm+M4u2nYpByfrnNN5CIjAFYM8q3zoESTh36hoZSiyAUcYwtd/H
BmY3qdOrEHiqtab4EhYSuftoVQfRiVfLoeYI6MD7hzvFB5d5p3mEfA4kCb+jwV0H
3xBtoSkEyTYAqpRMAzFeMNDcI84jJ7pTpwEPTTiEIC+GgSPad+Df03X1WoPWES4e
92ckTDcZiMgRIFJwfeJLlN+gpDx0faWZnjwEMgXUscdJXactxfL0b3xCA+QOI7El
V2Paza7NdQKL1RL0D9ZdhGtTCSSBq1jw5nRepVJ3xdqGHUHZvRiopYTw0AK45AL5
I94RgMoe/niIlrJKYcyArh6iA7bDtg3JKlfuOs7K0QYQzWmrnITJAeWJTkTnfyfr
bMrSp0t2X8Jk9aoKp2Dz0sWHSNShvHtaQNh3mc0/TilnwwQgWFqGq13VrFKf/D2f
gR3NWoJ2GCkxxM9qY8C8f8PjAWvgRAX8p2QuD0Is3d3zfccTOzAyVh4X6jI3ZKz3
XR1Dhp45IpOJ3T9tUgcsHasZ4PZoH/PF/qdZxiFWtIQw4L8pYUXAx+9N/imCKGTq
w1Ka/7/CCoFwfsms2yvNp3EUplHz8Nhmh8Xvdt5WZbRtbeBzKmlhyEhLDNWTWpWR
J1o/muH4HLDub0mFGohWr4/oVbE++giqxG8Kt9slqzpMfWa8S25YC4ISGg7hJ4tK
yCvzzM5F9R59zkPo+tQAdy17jAppVfWZcI16kWjSkQ2hMxO2MIQLF0hHhIsp6o+Y
Mh2KUBaWDvM/eK0VtxEBTPsKdNbYJCdxjY4Y6rLnPWctXWTWB7Gb+Y+EhvSL3VfI
jwcOISO5pyesnylPOBnURejuegipA5jgl4hnhThdQf+T25tHAU++sPmy7ak3uBBM
+OXh7qBOhuyezc1FohnLxmeTV1nTz1tCDS6YzwGwavuvYyKm8goioE2HtkR5I6tu
7T9+EW0ehYfDA+upxyg9FMMf/bCc5MspS+9ez4DNkdMDHSCZPRFMeCYBKJq8c156
tHLovU9d4iPB8ywTubyBvKCTnBxoEdY9E/Z4HlPHAnmkjQdCZevCe/7no5y04uM+
URyFc/DfKTpBmsRqNpLIbnfAS6I5IrMJlyhTu636fe8UqHRPi0f0xFxELvpTskt4
rbYOAJJ6yEvEsMkmHTunv95Ayo6qO/5lGxj02XOF3di23eY5ywXWFy0Ax+O7HV+U
QBnIAYqViPY3njkAK5sfGc/H2D9gZ8375x6mibvhQ+sURB4qWq4lYzMZ2nGe9u+e
9TtzhgbC01WKyQ/pBFahoG6AAwGNGi6TXQjg8/mdcdT+EAyPIlUFeBzBEbzseKVu
wNd7OjqC9H675faTwXOp0IQwHPEfTmgNKTDoZ+2odm2bEmzWfZwL9SkUuQQQZfSS
X9s2gDERpxUEiE453NmmSMuTlppGvFBV6tl7R4IIZDRO98BBXYnV2TYzayFtRRAd
+/1kjsT+F7SnDV6Lv20Obh3lkbjJDyn8d9COy6iapJegsa4SVPK40UOVI5STdGxp
acFXVqwJP4c7DmzNhPxqNS8jd2CNKzXBiJJ+y8EqaISs8LnsHHbTKrBnyG0sRG17
5atzGuqZAONV88Na/UPzbr5k5NBc19SY0M4tu5QYqcwz/3l6is3TCFL1kKyM3mqx
X+8/4Zp/caVu9mliYn+h7ZZHkZwBdRtW8T5XauctiUUyMJl/3TjgBaRx+npPuKwp
FydK5Vs+7DdPzb1/n6Pjb6KymWjhyzYIRnJZu5l5qnTV4kWYCFCow5V/WTbXaziP
OsBPJ7YTxqPA/sVqJxqlijAnT1XaBpzZoxdNTnIx1v9XMtgniz6sP8ejhi9VaNKb
54YI8UB1NztDg+Y4sYsx8JgUY2mFNsyp5AuAtjI6h4N+Npkey3v005vWDC/kCtUj
GGDT8fP7J+/VHA2OYuzdw0+551szsJYW5ULBkV1WBWkCOkXTlO0kP13rAzApBlsv
NXBCLipzTCJ1OOmGfVLOg3XTdlnt30EsNHDdKiEKOr3cojWevl2Pa7I/mELk17w+
1u58IwjM8vO2TTULCO7meWiajEo6vvJXcfWc4zrFPOrbU7919s2M+1xquZfeIO/0
qaFScV4QSdPMDODkTij1GvOWyDnWubQOBFbKPbvlvazsrA23sqxV26GK+K6MVgoY
QpBdVsd70fTEkf3O3aHfah7Ad0VuxL7gElZlEVuOf0qLPx1aKqPqQg8m4MFHjsO4
PHtcwG77ILQdKuPFtQgSyZM1/KIF6WM1GK9WnN3VUHAQjYMadG69XnBEbBKzgfwk
XWyhBZJ0VGcH2bObNwMfvM1yJ48veIXSywW5ZaQ0SCafNUdHPN5My/lkZHJikfUG
KCAA6OxF9M9DeBMxzh3oSDl5DUmomOkdvhOqXssGPBFrt58ZrWlKHyCbY8hu/r2D
HdZ3npUZpYvru/jacYlQzEg1T6lV8IwCE2tuaBJkxdT2+x0CNw//QssJTbrDZsFe
dGbgyy5KSMGi7BXrShYHhY3VzSgsUxjMAAKwWtejQ75FeDTwxwMxtEjV8opQw1f6
qmguBgjPqi0ELKYcQN7izZh1c1crnrvVRXgJDKosBsyaO2aD5Q8g8wthThsxjsln
iBPQ3sr2HMfoDFAvg5yIT5OT4QFkEwWTQ02/nbQxjsJnspugBDX0wrpI5VET+VDL
xEgU0IkrbwvxhOu++JKzfVL+ciXLvUt04zLcwbM0JccmbHIEgyIWWaxoNkW6tE/3
sj1y7AaRyO4FWJJLDZubxZM8Pmr3ifHmjUxn+eo3HUK8fE6K0ni8yVQvGHdX3Pew
D1zGNkb9zfFjDtfO4Vfj2J1JeTSMEUTVFOGc5lKtopodVrUJbpsMAUScaX/bbm9U
1GSm06fGZ2/9a8qblBgRtQI/XySCpcTFg3QfDF979e+QFcSEEmmowSFfGhckasse
1cPFgmVszz77H7tWZMKp3ggAO/swkymDGFVlh8K32Fkg2BKCJHNzWNX2k5aJ3BtU
kj2I/G7qWWt6wP2E7E2SJ6TmYee5az1gx9RaWrJis/rlGTEjFfmsFqiqtyvyPgiY
Iix/HXi87iuhx2d97ZDT7OIzc9pfB/p6LoARnE8dRIJraw0NrwPOosegYPodNm4X
xsFYZ+Lmlwb5vQfLMm57qA5u+T1gf1Cu+wWzzMrpW490sq7O40WAr4gcKt3oJp6s
qmUoxF3GALZW1hPE3Z+pVQcX0F8ScvRoQEr9qqUYww3ITT8Rh0ae5WDrbcSEd4qi
Cbbe9li+hQXE9k5iMV1Uhba2JNnqtGcoMTqiSaNjP6ZZ/8Fm77EJXcPk/VpdzZfj
/1V8gCtBuGYbBeWvV2LDaAXv+w9KFM0sN1Tpfl/TEjZQQPKNqVbws0vd6r+zo1kq
kp9ZXujbHMLTnBSh2e9MKbjs8oaavQJ/RpbtTHkv5Q43NUl+1H8Z8Hg247gxkZPV
cHgNixAaD2TxChWD5Mn05pxS8DPapnAgwPE9zMU+0rhCfZpqCrz+SCN7CVEPQi40
f4XGMBSOZZGp9rtkW8xavPBvJfD7qu8Qxk0PuWgSvFZoejHjbtbnGLR6d2z8WTyl
z7My9PH4I5I6VkPQJCt4+DyhhbUdzk+gComr+QCpH5Ep1WhzmR/5OljeHguLJBAq
jh1OzU6Jw1J3OUogOcB4WI70c4W63EeXeZDhqETXugPi2R2itnQ4njvyBKMunnko
ey1BLo1RwRMctIH323q+43RkBeaQb6a1q0WTM1wGD72rdnNV93cGHa3o2wXBmVBz
nb6PxjPjEmtHQF3ZUC6/s5KobgexbilGkjEB8KZ94wJoFDTKgLjiC4xoPMotV428
pH4+tEdDq8r2XO8onLKEV8RhBn/zonDQmXGp+NfU0gSgJPZOijiRzbbK79b1kmlN
Is++bxH7sRO+S5oREtyITiDxmQYJZEYEly31g6iRmyBhaPCY8SZnVijnCN2rFQU9
imGAtBDTr7KEtJQmp3NnUDI1Kspwzd8lsCq1VgCjUmUv7GIiJ5MkHaBH3yBkMosx
imQvT8K/zmR51tveIOtJEz1yoq7cPpp2yAZ6I56mW8dwrEWr7qKaIQhg3hQR0YV6
njX5DPW0kBboQxBNnp9vTSM+2WVZ9EtB9hIQ8MBDKpquwHt0Ec4Ck222r4rv/24j
16+oJ6VTWAcsHts8mtSmxFUtztVp3w5dYKCQdjhrPezgs/3fg2MsWHy4FG4nNGE+
7/n02vn97/GPCkX3ir+LgcEaW+EVUJ1L5Er8vGj5YxflIayktbHMJZWzpoGPIA3L
1WGa8Olk2RBV56odacolEUAsebe2goDzUm/VkdzuNkNlaWQnaWE+9McYow0Jz4jI
g+wdgDWUgt47Id6WjzCPw0qmiN3HOf7C0z0L37Bo0O8sz2ffdwwwdk01ojjhcLdj
EpAI1C2vw+Yi7DK5G7Z53+in7fy/BVB6YJj6MX22+WZ4M2fsGHWPXD4R+gy+UMRH
oDoJHwUWUT8OT8mmXAlyElHKJKmBV1uW6fAZ3EHlomjaaTsLSECSWxBMn82GYtk0
BaQD5QUr8y0cR6V+rwFye1qqeBb/SocqLc1esF71TglAPhSsE2EfFTLQ+W3BSEkx
OPP767lxH9QNio7Qswhv+PvpMY+VqshfuYFY/pxXGP7w7ppI+zDw5Ans2YSTHYa2
NDvrXwu/m4plZPvDziqS/WyCsLV8CgzzXSgmDTU4S2H+lL8sTT18x8Mq3qapWGDO
9GKQxlP3K7ZFMcWnI1DIRv0j02zkbM0Of+Y0tL6VUFcTbEtvbupQgW1CIQcJI1yM
K2oJc8j35AK7bOqwyIQKwWD63CofQEdgJsXt6LzrtS5bJ9Cfz0O42Ru9/NBiNsi1
MSdsEos96+nGzogJ+RouLgb+ixTXeTMzCJPROD7GrVoEOfVDgm2FMktHMZTTr9Yj
sZjbXoS/PPH5kJfXVAqUXsqMhW7Z7xml9LGqREgj5/CSlg4kp1Oxb6mBCaEhyPPa
VeZvAoqCdCLj4MHYw2MqAOX9sg4tgOFCtOaRk+AmJ3PU3o8TV2f8EeIHWu7sf+eg
PSHntz9c84OZ++QdteKP+50vehigJ8/tp7wNzDBBstJWKVTLYYbph3bfmfKkI7/y
Gld9fBxPZUWIP48cbz3aZ+83q83rgwtOpXL7IEFH2sArYWZ4+0Ly5LK7L6TenZRG
76Z1IiDSMyzyMRrO6RBpafAfoizmp5F0LnRDiGMjs1YjwHtTh8olu3kf+NwsWhYY
aFn/Rf3AsNm5MxBa74MYi2tW2aBM8onxwqJ5PgjgyeEJFC+hqe4xwWXDVNwL9wtX
DMzZ2Z4Xsnpi+IzjMl54yPFkKVZgyFfCAQx5SAvjQ+kvz30ru6Eou984+t7v3TnD
sF+s/81kdj2K4Ysi/o8rQpyWjGHKDSWVB9Mc0edCw74y5aZ/Zv06OAfDp62cn07F
kFswvAvqBxa3Bk726bl9KZw7tLSirAEJlTux8i0N8XG4JW03aHV/41a2eC1XE5Ym
GGuZnaKh1BFdpikz+0z5/DvxX3vB2wVCP8nTzqa4+KYkBAfWW+j8fpIdd5agSIEx
4wJR3esh+PJtDN2G2lO8W0NaD5hdZWhl5yXbCs4ZM/CWulApULjYvqq9HbabTqXs
/8219GGPT7TWI1wW34juc0uMQYWzvldhH0yVNahAMq21dqO9ULtZTaD7a7bizshh
OOFHTVxWgMfpQz7mVJp9morRrfP0MfDrRg2x3BjkIUQXzOCjINNrrVRZ5Uwuj2B6
0m8oPoPu9cJoXPdai9OUxDtcYLnsHhbfISPiwHTxUnesDOgLlKxpHxkZ7OwmdFH6
kk4yz9TeyaMsPU/UaJcaJVyU5fLyKSEvVWYdkTZUE5aM7FDw3DgUPAy32C7VMJdr
PwcJmOKA6i0TcVlhRV8VCYaud8XET7rsYtrCC3I+Sh5xdyXo1Gn1fqqp04wFI3Ca
odZtjKWgpjPEW/GisOgX1NzOubxy+Ay7WKqWEsPQqea1PK0DsuJqQ/51zAjbQVvf
0W8ZLY8cBsKoQShx54o+sSP5LCBb3odvGECMguSU4lmTDiz/Wtkj48qSMMBy0sWb
4+lY7Kr4qT8WorwAd4eiHL1Kx7WJzJMEDQMm34nAxhu3m2btfd6FEFPv8J4jPKzp
IMaaOZYpzCDktd4j2SmEDyqLZzegbTC1tPnAsetq3ceFq0qtx1xNOQQdl/kzNh4T
UPoQiBQQQACCRUM6TGag16Ljv6Evn8S00yXxVqh7vnvL3HaDE43VKZIN81GFxcAz
YpRZ9uWpcjagOuuoRWOBcsFJexiXRfJM9ToWhDjeu/wZcKcslCTbcm1pkqYuqUDa
4dgo8b6LYayDIaxJoniTxs1CTe0XeRepWeYVrBBqdo1Rc9swOJY7pGbux5LVAFUg
UqSy6rqP8Crcio+BcMAsPdi4NM1406KN2xX334uNdNK1WBwaITSo/HyqFQM71NUf
SjdLPS2T8lqYfvvxtsPkj9D0kV8a4rAf8Id3DrkBKRl+Vz/fizfNHimXse5LDTIy
Y9LSgOEKhY39OWHNCsp0MpD20DX85EWocbxfIEMknd3QC6z97S0R/VnKKonVikfP
OOU86ktNxPNURj66z/t1qNPpCSHgWu/iweiAodG0e4mHtbkqkz2gGr8kzkcpmCbz
Jb70f7GnPUZ7N0bqXEco4JQqxESFqwuy5aghmOuyI+RQSF3/wRvOHN3ai+q2a3wv
Z/eyyzFzQPISjXYpCO34eHocnCWgSCBT/16f8OLFp2h0ugqZafoqEleK+APsnOJz
ErnIv9U+76P3EXdiT34VJnU6o4pKg4hStLA8zuEavRakCI3uJSj7XnI74C73Mlev
Hvdr+a2Im3dJ0xItpKh8Ka23+PxWwynI4Fgxg429HNGze3Gg1fAGRW29AkPEcNRp
83CB7HJVb5k24lkbZnn7C0BBtwrLKWAOkObIAjgUx10hzvRx9K72zKjn8hx6cF+T
KzpRxKdEbdQ4S48Dm16P0NpVeuMDgdze5xKPnoK1TNm2mc64Xp2hfmVysD5Qgh4Z
uHPjsmmXAx58DXpGCJV/lSa/3ZcA8V/B6Q5FsTwgLEyzpn+g8L3T21WMizFYf1qE
dcl80crMPFRa6OFts7CYOXp0eNEJa4BVw7Y4TsG7wfmj3spICOuHhc6T7MCS9dcm
LMmLRXX+zONFGj4S8R8H8nWiVfys0iLP6mjwh01B63SAYuvUjlr8b1vzpseXfefV
aZsl8LLFOtdaiPUCZJJfAyyRE7xeFM/+9OMaTkNBlWhhkPCTVixy3EbwrCKrWROs
3GNy0o8uScnWUTwOGy+GzARF57R9OmtYoeqKIF3VX2bLjfhl3y6V34iwd9tkYaXN
olEsFJNY1s7SfjXEjCQGUPhYY6FeisQ+DpervbnPEFrzC3WiQTILGqFi0HfrBa1H
BZaDzvyH8QKzlL8R7PvxGbmPyI0+79KJA1IprmGlQKGLkd1Fs1wz+5b157T+aqmX
TZOJxsJy5a1FGuYbamQqp1XdDSN3EZ/+IcPvH9+hbdo/O6j6su1zw5uxCvpnEu7e
HW/jQuQjqOMuoNU4cRb1/gpKUwJ8w5HjN+aOGsBd4c2ma0b190w1cE47Wva8/j18
Z+nW5AlgvnpacfMxuYCPgakIhpynvBCFvz6FumTVFTOB8XqhigMs0pNquliazghT
5JkfBkZQ1qmm+O/63fZCWj9jpT68/mgoh0QQXmINqKR0/OogSjm01AWE7wRzImW3
uAoLC+2ttuclOk73HNikjP1348Dlpd7OamlPeHg8/awKYMPRlDPcO0itKQH3DzKx
B8ag3lAScFEXvZpc4kOSV0mYEc576qkIHi+mpwyxwGi+MDsyldYu/NEHo1506L5n
6LLutAroBaROUAf7Tj3Ue6G3bSyaNPLKHUENm4WX2slh9Vx7OhpxWSEsTv/T3fNW
sUculd9BwcQPUY8hoec7OigM5L3c6+8kskPIpahqaugrBiY1nPQbhI91cOSmtCPl
UKYb8ClqWYnYHjel1rdsqrFPdfo29kJIEqVbCGXHhlDZ335SgH7rRm/UkBKyp/qf
qkdVwRLyp+plTgikt1PkHF4+mzpzlNnWHdgTzlmDX/IegEOOFbvRf/7QKdFM0lNz
eToAuKikiMMFuyLZxVaELz1ztZfWS1aHP2Wt4q/ArxSpL74GVocllSzYMP4GK14a
oGQ96WMwaZ9ieJOTmSzKUBXZh95a4VpVfE7n6J32GBCVUjXfbgYmMOaeZ/R3nXbu
GKazhJOCJJmGGftPnF9nJs113kFC+mx725IqdERW8X3l2k64l9njduXTCOqr8oRy
b8qt7rg4G0/INcv1ynf5P0vzsnzD6c8RrXsT3+N9zPOWKmO5ltTrmJTxCnuUfxMj
w9Mdswgr7foyNuYo5pRXpiaJgyosvpEq365ngNISp8Xpm9kb7n15cpX4axiDTs0g
SvmptJNtpwjx32O7JlQBZZYhlIk+c3Gn6DzTa4j4YjFHVQboHOdM7tGnlYBa5y7P
yN2pwW+uNh/jemPIYOdNs0LvmiBP7nGIq3HRYoh318duIxqlua8BB2/BfcOWbu7l
7bADHsi+evYzSdYt98xn6BF63qgpdCa/Frl1EwqETuhz0FvnGGzDK94+TQ0ccZ8V
kTvlVHQiEffiMwZKJQqTWychwjLOXSXw57Ot54Z2nMppW51rpyUW5JsdPeMgIR9O
Ywg9Ux3Mt7IK2I5JGYEatNVD+sbLqb0easmb9OA9yybA7OC/sFxQKfr/2ZWIWY+V
neIKi+XsbaziPD1hJqq1Me9wMcZr+rOAprYiiVA7uc8uJnysQzGHybUv0cJR50j6
2lJkhgt3Zy3TA8S7+yy3rAZB/XQa25hE11SAlUV84pvIyKbbQfym47Xpza0h1Oih
k9scWXOexjboCJDQZip4ZugFA2ClpzUCAxnIrxz10eouxacbJueEAp6H2DeC8Be9
6YV6W/pHJq2+jgMBAUc20NtRldC1Ldbnc5+qMUzmbmiUxnF5rGqS70Lra+wdt2l0
npUVRBzqo+N10j0qI+L/ud4Qoq1nAZjOFEbI9Nxo8jP5LKHtp+P87TEeI9ipe3BF
e7hIyXlDUO8GUHmykBPzuYKO0C9pRzfATV+65N8sxBXZwDj8HYyI1ihJJOmFGwcZ
eA1wnIsXZsmIlToonuhAUqAUpSdfdyVoGNCzJtz1hyUwuSQzmx1TVljURwwLx65e
1yBSMooQ1I6Rm1TJaWVntNzyhUGqXGJuh/n6S1KTe5Edncoqh8HcRfPkGJuR6QJG
KCkaV2PMayLFZTZqXgACOjAKHgbOe8DZIWicuhLAbKeHGlgZ94NOETm+Cs6O9FBA
GYe0UdXWcvoWSGezZvG5/qMSGBdW+kzEihS922wnInHUsDC7AkmpyhV5XLdR53zk
/o/RgukTB7hqmADnGVBMLeBMLCUxIjnan0DkVBVdxpmGx/n81XRtueH5leVhGpkQ
3cygTQo4mqcAp8hy7S/a1pc10tfltE9nGIu8sbwaXtj1Dt2HoqT8F+5mK0CsFy8w
p2+a2ljBB6Jskuox3dxHyVjYXOgtBdfuop7CSeKgL1vp0b4gemBQFCBfqJEq5x5/
fAM5gvgQuMxNshiVAccmf7VCXDK8q/nMzQuLLFg68eSHP9HKWuQEn4GZIlSNvVw5
Yg6ybz1iP4/zwVmlJ92BnFICHkTcFrARsqMrIDhNzZJXrbgB42dIhAVlZMwb4V4+
xSnwxJCZ5WV12i4r5GroqTNel0N5HpRxwgYSG7K/QbOzC5JDLbY9bRzTz2vuczKd
qVop1+LSTgm7TzBpg/bD2TmhTMj7fkVe8Ibqk1iCWrMDxlQD8POtBe1tLBvQVhk5
a2E5iEMEvBQCRe8Mo9DU1lHc3g6fghXHsU6w1f6jWi75R8YqXBKcPbM3TahpZxaw
PbSbd09sSckMoL7e2waN6qzBnRahdqwFXGooT+LKdBROsYMMTCN5ZkwayUlsht/m
SqHaIpLMBnH1ZW0JPGvqQJN0vgHwYrmt4cz/ErCN6It3AMUhRboEc+pHQnWcDHeP
F64Qj6ckKTUK4+LnmqBQNo4rlcqM9Clh0OOrBohUnR8Bgng/7TTGTY/vb2EUccSb
AUUo8NTSDtuqWKuqjETOY8U8xS+yLS33kYF8D3YRwyjmciLXjrmTLx2bm9tzReBY
lqS/jb2I3QAJJtXxuRxUZGxuzBvZgwDMAFoocnauS/buH9OAVp0lVIYU/umUO2Dw
CqHHG8R8jrKRpaTcE3ew+HEXP55yEP9RQS4W1ZMRzYp2FzL1BHmTJyxNqIpBp31a
/nkqu267Z+NTbokkBI6KVeY0Wop8Ix4Y4G/SHVb/p34PqDRpbrIBJ/eU4LWPcaVO
qWFDxL44L2i9qcukFtoWfv2VpNe6NFoezBcxXCjna2ZOiGSJtqTXmjXErIZI7IQX
ok3KDNarHBIo+CcjywBA5thcRI9FZ/yEcz/OwpxXivTHj78z/apP0F4inPNpw3nb
fNxhfoafSsKqc+TEaDh43VhMSdA78xAZymbLK5mXTHvFkg3KXOgb7FM7JEng++nx
PlxLORy+3lnIWQLEt3MXBrI3Vde0qCd10AtN5O6mBWbvfXlRR9ukD7bmu1AEuj7N
uqGbvmGTjydHw8mKAzl46rA/jkjlPMVdr8S49IL84J7uaRvuceC+vNpmOWZAvoiK
6Dkz6zsbyy7C2w84de7crRdYk4Sr5p/ND57Je2ucc8cMihjSXPJgLU5CSR+zVZK8
hBiCiuU35th5a4mrzuaCfTx+WGCeCLrKtMF24E0Gm9tkuci8d/9qh9gKOoWchibp
GbCMLWcZnk/Y7h23nUYrBn0vrjXzOaZ6rY+7yqmd/9XKbFwkJkY4wOoumkGO+YbB
/VJpsxb2618FMgB3/DKhUyZb+oXI5OV880pXt3gRxwgU+kdNpP53UR0aQkE5Z7N4
Q023G4DXrHPPK3C+D8P/ih9MXmFZ24bDd1SoHJBbdwGqaNogjsV36dl6KOssy7g7
6ZkEtr2cOoepSS5DTUwBXDNOySt2kzOBxyyuuwiuyaCQj/7WNCfltpDMFTqd1SiO
mjF+YFYT/ZWNVL0sciKLJFHeZMgYWq0Aqa+zopQm+Nl5/DlNtzyAkMyDSL2hCEPi
WV7hHFO4jlqJxZZzmSd7yw4uE6e0+x2Bn/2RufGmZDZe4huzQLSCeD07ylbUb2yR
Jd9swgaHlXQfgbKzldv6UsyJdvY6kjCalDC3SYmTDZyHByLh0ZmTOik79gc4I+kG
WftNktq435AwyxKsRAU+3GHlpTeJlv+6+jjhC3vWmd21v6yzCHNqQfSSYIKVIOP3
tF6FKLH5nsgTXAW88Y0Ia6V8moceEG51WPC7HE0olk6XUDFxlxpTOZhCFC0kMmkz
3gk8n17FKZ8H5H4JMnErh3iUrnoy6J7YE/Cj9yCmbqR5wET3ANorhpQCcuKMHUwE
BzQ+DyeNe7w59s+l5ZA+FDnzabF5zIkO3qnKtIRXdtoAe11aTvIMwUKzftUhgaxX
UTxpDmsrJVt3UiZSFJGlGlBklLAgnLJqmvYxM+Fm3KrNIK4s2KHIYor18iH29o98
7rOi9zAYAouR0ofNVNIoj1jhcXTKKaU/c/ajzvNAbP826Dd6RAMoas3TCy6QyWTR
W8bWOFqbpiunTmO77RN7e3x33MoWvotRSzIvCUui8y2YrFivODq2caOe+3nAURNr
hlKLuhZ/VpRWAiR1zU/y6F6gucwfFWk0eR9kZDDk0PsN9Sei5wSiII9G3OwdvpMF
Dg3TL63M/GMF5Ombq7JSzdV1yZHTNNHNRNuiMMRxvcTU0pb/EdkysCbeZXyW4sxL
ZTPXG6zTSlb9kwA25D2npQkBYVCEOkDpmdoMSGb/Ca7C92GFDyiC3H+ZKsaznrkv
7u5Lu4ymB4XCeIAOrVo/iJCmvdH/uDjppPKbWQKSMPq9A4Q50ARzXujdKibHeMPj
2DzUmoF+IO6zkLu84FaUpYTY8+E3S6a+oWE1SkPgHfUofE0dGhfX/E1j2jjzpoUN
GDe0P3IoFpAiTQVabDueJGoPnTCy6pk5vE7mr1T0GWu2rWrnu3Y4CqO/1YN1Fchm
pJQN3mOAGJOXPJE1YSOvBbe8lALagfgE4ds3KKSMpagycf5XWEGO11A4KAuapNAy
dzagkkK4rGUTUiEMex6ajM+Vqyv9TX+kml5wW3lGFZ+OtrPKgubzYZKts2YORHaZ
0ucr6nwfUPp7XGVVYyEv2U5TY5BuagwxAe+QNeLGCslbzsXfVz1GYhBuCDx/a62i
5jGWhHcZDsZugdHlfs6YwPB3Z5mH4nDIzz8r5oo5JFA2ChrG3UONTxMEKZD20S9r
i1zsUNEkOt9WKnegU0tv/tgdfbvQDBrNyUUlWONyshx3VVsNhgD+BnDsS6zLLMfL
5OBIHc+fnq4KAtzgnmnvRwyaO1LoVavqW9dyx3GZit7esGicntJs+ru+r5awJFjl
GcTqrA4Wmq0+id+qSZSBnn3yTtC7ucsh8Zne2MabQzFnxUel2xV6dmjEeSJ0sDsH
XyMjk1qHnnpjmD5xInqxDRPVy5MQKfo8NA99x+owWgEOOxQiIDlaSbMK8WXZ1CLw
/OfSyTPMkmPEDTyuFxXaYhXqQzTk7OApxfUiLdt1pd6drRNLT/BnroCSSCH+ba7T
aPxuPZcI9AnUOqslkGOQRXCf+TZF2gBbIQl9bXsTuTOWp8oki2d6Dn49/gazAU/I
8pg5ZUidyi6YYlmg7spwtHWJuDHW+MHgZFsaaHsy4b+2SUxe6pSAlLzyAo2h+r84
RmFNsxzVXu4vdjYPYdgnYmdMUYiXu+CksOdvxZRyihNoQqYH7zxCBptoNa7A+pws
i3piSXx/l4ZcXfAw8wCCxjCj9TvR06HQMpGgGKs79Z6/tpfLf3Sc3PouiAhLiMQs
RXiEDDM5TbI0QHk0gh77w3RNLj+iUJ6WJbQqYjjM5oxlAU0G1AID+aSji9ZdYXeU
uu97uwB7Pp7S5KYZNVJXrZ25vlH6wCA9erC7L3XEaQaPWAk3xouQRl+n8DZJbml2
4VGs12W2h/PSOP77xC8+bA36/esMbMmzdga1DNjinEbDEVzhlplyWVSWa/klJLKH
FCpHPbFMirUL3JVwrZMgK9SsP+gdcnkKH1EfnObOhKJaDX2PR36COB9scNSXc37J
PDMAjJ4Cn2NyYgCzBUgjWSaNBM4v7RE7V/wFskow2EFIbEk4Z8UBcmlUzfNw9XoR
JloZjW0DfcvVTDOAD/FZ+54QJuGw7Wqe2KkyXoUfruCH1HR3MDa1eDS8BWxanV1W
tC+xADKMRgMbgAreb908VXYjGUY8N0v/IiEI7iRPzL+9eQg6GyVdpScziVD7O+aK
jkvlh7a3B9r7nVbDgMLsBwkIbbCTC0zogGJ/2QEh59s1lRmRLjh9RCKLoThohoOa
0bJioB8zJhxyN0XwLF3GqoyEXfuhk1+qL8xcY3U+tvuTcfQeXRINl4kke694oJL3
+wkOw0P2Zvg4G5y4/L0D+uHlNolwyrpiPtQD0l435oos0Sj681gxpZ9rP7uyqSTR
YXAL19qys7CKwAaFlIHfjCpG1N/vElT5QnUbjM4YJJekxNx4ZWo/NZ0Hq1QxeyYh
5wT6nui9gQIa5oDBTytSUCGLhsrZujd/9RF6jBhKA34OQCMMuR97v4sw6qcSoaod
mMlnMm/nU8TkqSp531WOuCJzm0hQTUKyri8ODJFZhywBLGsiFCnj1/o0ZYlwNm51
KZC3wlw+fipOJu2pJXlnQSI8W0C4ZRJZCaob+gx+cKFJtzUIBoGCPbNyqRFUrGXX
EcIv3TDatcYGNjhnmWa8aMrEdKUHOXyXwEUp0F5ytQx3p8CoVdoDkq3KMZs2Kg9W
++8Rl9tGp/2AxdViKmgqIFKyqQLp7Wakok+odpvUV5tBFvqLIe2WSDmts8qAm4kd
txPhEyAbIXiF1VtyXWcpODRaxqBWqwxPhrWLQKagnvH+ZNfWx8giKjG7Knb9niv/
oQw2Jt9T+h/0Lvll2uCU9BdZgsojwYO8ljEN9I2vKedk+kyn4EGfnSGi+s16wYKP
KgIQR8bckxqGR3+5KWn8fvzYr/uoBWJReSOokTIu8nJTP764n6q3CRiFPVNVoRth
U33NGUhnOwTWVN6Lx9J9quNcyHJuQv1XppmN43V+5zGa6vEoDr7R4UXpjWhszalr
lFzLDiQWHcmBHBHO+ylDYhw3dsIbHdKLooUuGmLr5Zv+/ze/QSvrOBRjttPvdb7P
T6w/jKoL03zxszNaPsEp10X0RGUs9+ifWoe1Eomu8M0sHh3dbHYOvtvxcgeD6I1O
RVsZTEx2//jheQEotoYaHl9LCk7ox+UWk4Nm0QVx6GV4HvJXAv0U/UW4PN6OaiCo
bGDaWBRzYfR74NxGhXyo6Hdqa3cjnich1shuy9YKM8QmLEE29ig/jVX/WH/X8kLq
lF6aD7mQHFu8w9w+OZrHObGOcklgmyT/yhL02dD7cTVJ9EgqhOaP/GKEJt8+5lLZ
ORHmh02ggOglSZPopdBveqkAlQ31uq2Csawi61DFrzzgHzLvPrgMLxX/E7djs4C5
tRiAMqCIWdqeAoH4Q92sIvXYYKK9r6SezGT60E3APAZnVoBHRma1Pf1KEsR8nUK5
hSB5vf0jYR+U/rO111rHxNlXYgevGW6g9vh5pSyEPnGOsrMU7qVqo8l1TQRjSJOe
KfohlionJOpkPVsLMGX7P6hdCWyrZV38KUAFusLhn/rlhzZ3z+AjzlhdkYN+TuA2
qokx9XJ1BwYq9u559ASvWAdnDzwd5fZ9yWJQt59dw5FQ/+mvjSJ+lzXvqC6K4MrY
oBt7N/v7WITqp6zbA4ees7T+XzaFoRFZVdv44wwmT/SdqMhD83aQCFIh4OssXtzb
OdH8+oa4flHGIANo1GQlB6mG2labLGn8Cb/ukD07BRYB4h8Egpo59DSYqvkdoJPq
6yJR8s1qNrhZwmYzvAkzbn+UYRRkEl++q7935l7XAgC2fPS2QVHN4F0cECCAXElr
yAnJYd/0I6Q9lJf3ciNL3/yxwF4fQM4rPdvjScG+CiOQXpwkKIciDqvfiztbFhiE
T3bOY2figPOGfL/4r1PVmglHMwzYKXigLhcZsS24DQy/ezT7DGPe25Bbfevs51+T
ivu9VoSbtLd4wzi7s2hzZhZw1e0dOydR9+Ed45C+ZzSOJeKav/+jUDUC+npg3a63
IzhKyjpkTqpOiWYpa8Oh0g80tFOozklWskj3MzmEaHbih75Ugb7fNWn9jsavfBIN
8QPz5vqXenZ1OfFiVuimZTGEj5yMlNZ4ZqNvVFw2QJZplxa9mNAb+7c3fGAjioD+
U5DtbMImCTY8DMjckZ0vp+YiKZjDWtzvRPlvyQu+Bg7Fxgj++UMWhWh53D2gue6f
05zBOU+xTmMCmfjL2oUJpq2HeTWgXHIt1Y/5XLcOK+idO+/YtQY8AroEudsr3uen
5UC7kWorIlJaSzXH4d/+cw==
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14608 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/Vzsfl7TOuMe4xzV7rdHsSWg325tC7j9qhAnsScdFgyGVVNMw
8AOHS+ZyP6uxLKpP9hjW72eNQsDSngfh5tYXHp/t3mJhOKGJkNrV4ecx2PId3Xrx
TwH6PHQ4sZSKmPriK59I8ukeVNz5B6ekLojQfDA/RDV96gYdbsx5f367rt76UokG
02Ag5cGfYD/1oyAM+h7WpcI/GvGWvX7nDFTJYhST3yQoZcG3cjPt9dRc1LwE7Ttu
JDByFVSKmrSU2OWapt2aO0D1xbnNxTNH58fjxDw/st4gJhjiySP8JyXqvMOCHEN3
hSU2MRPGkvQa7vFN4h2imhCp473kld9FsWp7zetf9I5M+hUej3rhvvM0SKOXruzY
3gQQBhf4RnueKKahNApjj+UyR/uBAx3Wvbpg13IjbZxiPgYU2T8wzQeZshvBIlum
8FE4tCzxHLzIwiZQUuoWasSa0BT0bPxs3s2NDt7rW/RglbWWjxgs/huuKT7gzoWS
NdRuRc4BBd/0YJVynCoGWOQlaEhLvGlk3/iYYeSKhjyUMwra75mvhefTUhnTgCsl
X7VkGSFSdeobruy2WsQ+8ccWzdY0Kq5BVEKJi0SHLrfyyNxzFjmC1/qXF7e4wccj
5PQKY9MoBd5pp0ivVmyecuFNl+aQ3CByaR7A/wkGT5aNoF3xyBEyXY4nADVFlIwe
n9zYexV6BxmSsjeNvN9sC/X6/QSD0XQYF0nTOC9QTXTxnsbe07QfmzVhFKe5XVq1
LZ04o2QYknK58TP+7B0kgLuOcBUmbsLIdyuYx6VtjOQHQBeEHlhi+YHj/TWkCi37
cNRRHkZhqL5yawGBJ7bmhBYQPpHxad2zLtoc7LGBywlvLl0unuQA2SFfrBpr1sgX
4T+MJWuw+RPSYh0884Y/g/VmdR7UhfdesqgYj7xWXjN71T9MMXGQ3ZveEmJMH3Um
gOXKJolqHyRf9WdhwG8pAfIzJwv+hc/wzWpdhb8UUpqxLBSAv99z+d5zbIuosGpv
e5GfTuNNO/7L0UFAHQIUqrRwYu0y0cPnL2GpPOVuSfxFuJHTs0BbEC58yuWINxbU
NXmnQbv8fFJIBIe6eaTEArbSSV4tOBu2RQZSx1xtVnCfUukk/y6+rk9lr+Rwc3I/
+rDWOWSsx5KyWZZG++Nrrx+PxNwNT/MK5LE+8isxgS89nKXveU3u+G/qwassmix/
0N5Wmt3Cmk1tZRbu7fc9I7XHqEuUtJOvr1t2rYPe+/dsutweUr5IT+z0LJ9Pqfx/
RuislI0aW4KWg724RI67iO58EWKrghYgocjIDOLukU1Tt9/EK8eXaan+WwAn0LFe
k/7BbTsRIe2JQsKqvsFkJst8du3Lbgy0Sg0Xf9k//wIfDFmdNCvH1D9TifSxdHXg
zmEsFnVUipix5YLm8gy4XUl/gLIIuYJjeqWrn/8pgDsmJ72yJOjRxHqiPzRvLduG
aLdiSNK3PdVyf7MdkE8yg4MbkJPbzv6EpNnKsVncjVtvmNRCKtWwusKaWtFSkabB
Pl41DHiZTGYLBHEb5O3vbxPJc9eaQpSzsJMOviGBrJrtduwPDQqusxb5JSwqOBgW
KNvIiBem8+TfxmQjOZmkdKtBXrSqbnTwpyqJBetEs7qkMbaccnIdXiZYOISXisDh
sexEWardPci/UBqUs3nAfmgs1lcbQMi2Rgo8RtrWCVtJedjExGZB2ooOmlVrhLrN
dH+UDSPCl6prJhiIXkzQgVTDt4MYlVDtiMPy2oD1oFFjuAZoQmgKOi7V5w45mQlg
EgyLixIJ+hnZKuHSqDPEd6lOqA/4lGjEjDTTbvqUSAnnPh1eDfLKB6DnqmibVrkA
cbWU+8ucU2d/Shfch68ENt8cPrYf5lzmubRUZxapgrwoWeC+sRDaTC8mC4FGkL+m
y/XfA4wCqURvRmYI7+ZA5fpmizSMvSNFAfELoVAr2VU8LSSfAIPdUmrKbmzCoHUb
51Es8QC/bFrrCEp8ksr0i4Qjem5HAIyHKh+3BeKfBREObf5fPrPwyqVOWnF+VVuv
pWKGjDcG3NU1b6F4k6chmP7ykokdLJQY5H+Bve56mcbLd/JXTOiGPyEEuhseB3om
8qo3/eErxLUJW+MJm/QDA/rqDvi2pZhyx+RFQbUQY6hPb+N4B910rfLISHn7laPy
xSMKqKdLgtcVWolPp3nNeVSZ6LWPAv++eL8I/APy7UT8KKNFwX7X4IEYBgu1IaMa
9yoyvXve/gtOsRkb+l51cv9DltTeWQJ30/736/E0H03zufpEBVlYnhXIylwqk0lO
10wPwlbSgjRuRtwVJ+tF/9RFIAeb3v8q7vGuMKxdymZ7leye3j2P9fnsLwps/ehX
gMLTm4gxJ651R0puvBRUKtZ7S92EG7p24az/M9DHyNBz0Z8jyf/D6akYYI21pG58
d4QmfwyPNnaYUGvZTjnf/wmHpya2Ekftj7HOqkyD7mhjLQd/CTRjZZ+VwDzUEOWm
VlQT/efZLM6ob8MH19Bj5xrqoOjXSJMNYGpDQXRLKAExLZNfspgkBJYMHJ628T2W
e3vH/m2fB5KLeyaoXKumubIfyJOLZw4MBh2015dKUNS9eJ3x4TDUkXod+RqhlFUV
bzlZTP4xZ1aIEdzGHJvryxZBLRlQClai6PC9I545T3/9hCH0inoxW0AUH1nP0CBq
iDoQUqqSSXHlLEHRDMxTLUotZbDfY1CB5MG6pKcniZuRakHoev5pfUVpU6w2gwGs
tHY5sGBwmQ32kfXXroMKAtXsJOh++p0PMUW0w4MgfbHd+wpLoidy+qqWGW/DuZVZ
r2xRLISe2Pj6oB/Q1HwEoKr7x0TgdZ2QTSzY2XZ+bIncBeiDkfANI8KMiYKFOW+u
m96ziTKFAGCBI+mueE4MN7PCo8VTPKSBTLsUXioM08K+wqybEy0Xn2OM+hEBHDxP
5IZasg82BlnS0OPRt3gJAAbvflIizF4Zupdf224l6GBA/ipqvpLiFQBudy0/oSDg
8bPnV8yE/WjhMrvz4LFOO/zoSGm5XHRHbStBzAcA+MI4wTsW/VOZSR7KZNRfjhiF
qgAg6tuNl5OCkm6BC2BJPcQ7hQK916Avgk+HFUlr9Ylo2IRSKHDfHfWSTkfOSDPP
4wDO/0QIhOuzyEWo+segTSvrvNOTZTErJYsYQTJzi55/aMphm0z19evH55wx4JaW
PCkQ3Twgv5bdslbBwDCyjMQJk5yUk2sdGrPVHA5J7z3wMXE3YhET9Jr5vJxL4FYy
kIpj982MgH+kiN/dALhircnZQcZi5u3XFJQZ0N7/U3d5L/rcGE0hTt/CvitpR5CS
FzSzzoIB7lM9eABg3BdB/hj97EpxwFcteD7M/qrbBx6shqm8q7sYmczr8TR6X8eH
dzfm161ObxyyEgC9/Rfz86AMec0W6jKE4yomfEOP7Pc24KDbmSB80cDx9tUSZB1Y
vjp0cp3ZYh2DLkOwrcyUfhtBPPnxxzmXEgs9u4SkKXftxRw4BQrdsjAC5lSxBGPe
zM3RFnwmUJsusEP3qhp1IC3c7oS/YWQMZu7kOD685Y2iZjfWl7yl+zgFH6stgBbu
NR7RgSGYnJAssvz8hIcaElVETRgY8MJFqKoj0qUpnxyKkQN3iCBiouH/GkxArmD/
Dmn7DnnwUy3IeKgmutYrdhfwfUJuY5f8NgspS7FTwkbXV524jWH/2Z4bNCOSoySD
olyGluUULptXqrQYx9jjNd6BSX+Ia0NIZe/LQPRl1JueTvYGigVQPC5kTyw4t1ys
JWuwIXt2gsU0hmb9+/nNW8jSzZd9zHZeauc+nw/tCjUKyqgxIWX6qot5Q/iCU7Ga
zLu9iRLCoPW1Rwbu9oUS4b3IjJ6eeuP+kbEt8CVlXO3jQ+FDXUIXlAU5HVp3Tfaj
CmTTPwuO/J+dAuWXzJtirYcMaGkvqw0BQVhrT7cWiKtNqRfcVYdCWQ7c1MhfzBFS
YHXBK/PFrF5U625MU24r6T2AOc3oY+72K4Seldb/W1x4eqUYtRaYd4kQVe4trZc0
hCtP1JdbcT9OuCM7HVk5j32tYv4A7r5lLrOycmOa/MMPo+0yxJUrHsrYGhP+c5E1
AqRE7OQgw3v46O4OcRHuM0uuDXVwRb9/339O7q/IvMXj5DbBsRBRQ3IWrFgfHTEA
+7kOhaNvavytZwx4qDOixJT/MXZvXYf0IpREN+SHkd6ReS89cUtgBIulv2zTU2Lu
I18MqHRB8aYdDRAvy39JOhTSS89fyTRqG4l2aYGBHK9+xBp0LL3qpV6ChUTN9pfu
QJ6skNL5ZWpB+4Mxok2lP0u319bWaPUER+MIwZvlUyhfWVlDF7J/GyT0/pW4foEL
COUkS5XqjVm6KkVbcMQM1Voz3Rau7yLzkNZDyRR4UV37Z83B8i0wiTjh+O/5oY/g
dnUZguQvlEFJU/ILXAtq23KuuxMXThtFlMRrBwiEL3Q8rZdC+9MC9zahpvHh2O1p
zVPC5YiE8hUMGh0SC5WmNdWP4v4+/9NdGvNm+RPwp6hhk4f8oqSqWbSoe0/Z0iYM
VluHrDKsibUBUzOBO13MNhxJkoo+uSbZT4P847hvmZtgxjDJx0pL1cO91QZ2TfoA
wQ7tqx994MQCjSKuCa638kCtszZJ6B4NEldC3G4aiz1HGARQeH5OJoEBKeznQhpN
Eyvd9Jga+8Sm99WtzWiHR2KAMqtHt8x0UrtxxbkjFOCWZnoEQEY4V8XW8/TOmY1o
X5XuT8ilabFVGfxQrRU7dvLHvS4SHrDotdkbSMm8M/OsqCuVrjxQg99/9oMXLq1U
g7/71OSo0j4qLU05LIbCPznNxG7ekwK2kx99PXhuGdOHWWAskkVoNZeuh+dHOBBn
o5TJb+CCKsA9EbgDKNoivzdji3FrcBYhI3jkoOo1apAyBD7Fi8RwK654oQ276tMP
9wRvEjGqIv7EZfzmDE9qY3ip2uIN+8fdtVp+XxV2rfQmbw1tGpDPp+4EhNmKkgQW
UEKsOd7aU7vp9xj8Vc9hcztdOCrMWQEN7SBKsIkqrExoeryDcTYViQjECVXKPohs
YSFUvINieuQnHzthZmtiWC0BXF3Rh+7lg6O8DF4U9zBNI0cNZk+jIrxw3LgkV4FU
AyYiqXcxHPRvsPrJs0M+zGcsSJvby2JhIf13z5ZxuP2+49ILoEEV2Yi5kj6xz+y7
9jJCBF02gw6B6C5Lq7wH8JBJTb3WzSeOi5gawL8t+tr2Sz8qg4p/j65G8SuBD07b
fIfCyjl+LK6oi1HeUXd1jBoBrB50yyqaSgFBL6dQF7P1nezhoxNY35tQpY4orAA/
zbVLK0eH9TOiw3ZzLEmpL9umHw5vc1iztDC2q7IMhKGSAkpKDl6+FK/Z7HgJ05vV
wNlMUOzft7vwGBBw/Y1V31n1hPh4v62M4vcYxxDfNj8XhoUbv3/MAxgmkTWcWVh4
TMjxkr9P323//pjphFSPOZmZH7biQW4WGrvkUAkBuC6NP583kVjigvut0yrGtKKp
zMzGGViySJoCJdh4cf6zQkPHy5+aItMX57H/ihbXRphLL+1dRWCDPVFlwf5Y+CWc
zBmr4NrxjSPL0l1mTpj1IdT/IO7+Rwgw2fkztXc+3E1J0vYZbpcVSE0GIKPpjuYU
2blEcra+3hFztkw2qQUr1xQe/nnP4dbEHbix3E7pwhjwGk3eVW06CxyvgdMbqo4d
wuyZcDEgPa6W5M7k2gpHSV4TVE8J+2vyG2XiMwvy30Rf8+JdZMQi2j2UZYh1xbuN
vc2Kjz/qRySfG3J25bO87sCoS2ZrVDuDf1nREf/xbwVUVSobhDCnSnRA3ssEqpqc
YcI5ErfY9rD4SVmVjycXgzZHmJPJGBNj1JRzxRnarn3nq0b1AdEbVwtwMk0HUIw3
0wj9LHnBw96jRyXTF1BVqjMGIE6MHb1AxHTLXG6a8MuM0y1EjPeMEE2TwJ3BaNNg
dtaL2xgGbyFX83f2JPoFHc7XpckaOt9hZdamc9+X8MyaHGCFcvv8lt7WUeGUd356
zyX6jE3OuD9WIShxgZGcWuN31dMLY1qRM7tvUrh6kfIUVSrQLeRFC+YS/254aVSg
MR+uebd3iy84mLkGRq7dvWg1JY0KEYJJ5xr4jPOn6dVk4K8yqOBOgMu5cY677zzq
PZmM+yr7FwEF9efAusBK4OKu5yZY3R67H6DOlk/R3w12T8W82Jj9tnYzebnPfmKF
Avgb1e39w7bsuYH1cYzZ+SXQBvPjgc5jCKUI+3Hli8QvIsq7jm49+nAg4apztUzy
9U3TC+mL5ZlkCUQntifZmEzcdbUGOHeZ//ha0YoVdYOB/hMPZv8E09U0J1Roa2r7
/vCUgosrbV5FBZYWsJ8pdsgVX2IfFyWJHAipMwLyc0NiCPzRaplIomB4p+a3h95e
i7/fKwm/HIUGFM9HTWtlcSdow+11TmmxmffURwqGEnWcXr7XljaDxNyyq9SeCsW0
YHz4GDoG9N/Aa/jnLmJcmVK28gbaBkNDQ+oF/VmiG55J0zhelVIhZHzCG7E/vPgI
bL9aWvFQ26m1VZJO+ZGPZdP/M48Ke47R44INQn6W8L7Qru3LmbtYMuJRWtf6tGsa
Mm71PEJpI9JRTg5Tn4wNOq1L21v3LVA28PN5rHb0ip65yXkUuZgzdeYGGA5UOL45
BAd/M5dWUl7jpeonZwsPQJeJyFNQP7CFWMhkggg1AvhOt73FJVHFxhCKeZFU3fQH
kVxfShv2rOzyNsFJiFvMKbyM7CzHMrBV8BN56n2OO4oqOeKlrAQpaNlQ4KNaJZ4Z
sr4oNv8Jyf+6Y2TGS6ZVib02GLjpx6hwMQsO0Gk4TFVUeM0PMe37XSvuncgxv3va
4slEpWlQ24EZCQsncFbFRFAEyRuLZ4hovZiz+p0+cLqLLI0atdqDla5HNZNqSsXH
Nvf4B6OPykrAT/pHO95qCih9UvSdvZmwtJQ7K+kTtthtdEtZIsa50mm08MNyBImN
GJvqc2FN4uBr07BYqBH8mq2PgyTBxMAtx5rcjD5OmrnXfZLieHYU0jAxR6mjRXYa
Xw+a1dvtXO+l8WYluL7RBnmcFKljgeHZJSbKiqbaE61TokBwoXL+dAF2lWmr4AOB
z0MFm8epytnr0bu7EUFrY7PiWa8FnkPBWJ/2Wnb+2l0zAXOdrXHKKxTs47RKJWf5
NDM9QGsy7aAq+EyEHkaijIRHrLOvkOcwB3uPGEBQoLBSz2g1HXjIszWybe2yTHzT
Mmnv9OT4lUCSE88W/JSQ38XUUDoW3tXJeN/8VkKIv4akmO7+UijW2TlJnUvq7D/b
GrtCYKHq3T2uq+ECvRwT56/WM5QmqPgQOhwHY8XX14ZJ+K8PtMIkCG399JnXVBNd
e/XgFUqw0AgNEwpLyBHL0+qgxpVKRE3DwNXpwt0QJ9+dYhgqPNcXV12noYMY6N2N
RoDxcMgzSuRPIenxIvkhq+N3wVIfVznCNsOBuUibDEag4/48QEGuMQ8GXL/WZ3eR
UIlXy3NggGOAkazlg4YkdZaPcxyGEUoyHXUhnD05db9lwi5jzJFLMSn7aHniO3Yx
QwYu4iopXKC9zMoBk6IRUhQUm+AP/Qld63To3LtWbuCPh9IRVBzzyCGREuGQKs38
wSyNLbdmE/ZcQBuJH6rns2hholXgQQKXHZAVgDFTOXTRDao+yTAYj9rWZ1r6daWP
f0AQ8Nqo3D3DE6e8jRou7wxioF7qC6Ay3Dq9ggB3nmcEB1sdciijjE0GCubAOzc/
ZeAsE+h0lntP3g+uJjFBc/L2oY/Ll4XZzyZta4iSrrEKihVN8spOVxO2g7l6xusn
UxZdXg0CsaR7YIdPKQ9QeBLgrlGZdomQNRou3CQBmmPzXbb0Mg3A1+9oo5YU30Nl
lQijbvVkC0WyBDvSjnlMzm+wyVS0tVGbx00cn5FB2ril+71tHfjSToUJeR/TBirU
rHJsR9Z+YagtLfjiw5jk2133Id5MBxP+PL0IZjwcoSiHoYGKTLphrlczkSl1eZaK
IhoE1z2pKf+yCETNmUVot4eRVKiDdDfughkcElFU55g1Nylg8MsVWRV4Cz9dBqyX
Oa5MebxtgnJkrdLSPDSEDlnXAlkwdIbD+7K/UqhggU3u3uMFmv6lDZmcIVFxAFZ+
JaTqfikq8iwayU743mH28TxEljFlBwlRmRYeFOH7ne6f3sk00aQ+vuDWzfZQAlyt
R9AW084tT4D02M9WIlXFM8kaP+IzNSg4TJzuhD/bzZ7eLlcfqdkScduLW9dhU8Pg
s1SA8UpM1M6ejQUDutrwFf62ww0tSFZE5039UWqRI+52MCLc9hMwEVA7mZAEt9mv
GhpDRuEPh+jMLtBtyLtOsU87lUOzovfCSqwByevd5qnHFZQkKtm5RZJOVOz5sqyY
bMm3n/Sc3FWgE3r8uD8/cv4ewC2MUg4O3rjdxKBA7r3DrG1b52z/E71BdXi/cyQ9
nkAm/FkBWnu+GIWo6cDjsPIBS5rdMbho0lRbGvaQz9HO3hPWZ9QwM0XopCMVa9Wo
Cmbp0caftFP0tN3WnEvDXmN/AHnbCRxoRSQTV625u6rQo01nYUx8YSx3RSM5wuaH
NhfgxbpsSm7XgtvZXiFWlAxYxV/sJQIHkpMvyUtNumaeDwJjlZYd1yHyN96vLcwU
Pr2fU9Qh5LsBhp6RxNTvhO9rhTI7YTCzB0cf2XzlVTLgL4Clb1tuhIrI1oVnYoug
3gb3AKpKa26VRkEfJU3mTJOdAetpO9UdMf1JS5UtbHsriCfxf2BSgLWQzfb+LFe6
BdGOlZLDfV3MppPR2tdti2OHtBiaxl0vwGhYgqvVvbwCveU6zpXRPdFrb13vW99M
l0cGPXfUhAbKp90K30fFnVTH4uuwJZA2mcayljeIuVHyBKBLGMJ7jRPGkkQG7DQB
GGgCqh+W1giDdF2bf3gMOnoEYQDiqj8UAloCbDqPw1USMIyf7ByUw5wW7vFl08v2
XZ+D+JnJ9Bw9/HeL3Ayy7HmCccQbjRNjq5UE03H2zuNujlhEuH1rXEiHAbZiR1Qx
nnR7ovTkCCVfN0XjUNDR9Ja56LYpoPfnQfvlnvuZypg8Bz4NvcE8dg3o7gmZt+3m
+ySkgr7AP1prWqBPtXCppI9+tNantcqQQPknngGpSW5urCeP/a6NRicODMXBn9dd
Kh4ky0twKyz8+UhnbAyO9cGhaxKccTdEkwDNicnsQbJnOYqPcpgET1ktPM2uGY8A
7czmJ6v36JtN8D8hlnsLcV4Mm7beURNr9IWzKSCXehsuPKgx+VE6j0EfE+us6mwu
XsLgKY9zwd0wrXQmUBWdR93eAulkNZpMGgr3s4LNTTk0HQsVwa1LchZUXT+J2eMt
Hz2KeBXKCKc/dJh3IPxQURDgQPgqLceazmaWbq39Y8MYJ4uL0F/wgvidZNeY7x41
6pQAZ+AqqcBMAgdjqkGDcrtrEE22CONR1VH30lnCVHq74IGusUZcUX/7AwiJ4Lit
jG1HBV6F4F3nvQhSgh3PfKvTuCBcckLg9ovyBfTfiSlcey39hJscIGJEiB1j6JnF
cTUNo/QFHgAIyEY9gF5pFucyHKX1lQRxS/c+FBpeAH3NVVR1iJZSB1uCdf3UWRvb
zJacZ42mVeB1OEcCzaCo7cJYmfWjl6OUojCFPE2eB4MQGUL+bySwTe7+m+DDfW2B
/qiJ+1W16Cfcmr3buBLPhQBmzcTzYf04jOK6IAWiPGm8eWlAqDspjaZJCKVnmE9o
afFxGu1hs1nouwAMChnMq5Zl6GOzRQ1A6176EInOj80ugk74N9oo5/R6LPq3mbWz
2VS6pJel5g+tQXFf2sQMrp5rK4x4K45f9Jlg4+SzmgzV72+3Voyex4TzyXkx0V76
8XxxevSnmBGd3AdeRT4UkAEesn4hBr1u0TIF0lDoix1SBuG2z0N8ZmZBOMEFV6jJ
1RGd75EvzOpYl8sZd07BrxMYy33BhsLeoTxPnwQbIGZzDeEh+0pJxEOp4mSzeCOP
enSE42y5Xe28PvDkO5xjjD55IgQs54nVrGLwj5kVkIZ8o41IH+ToC2YVqMxf+Afp
FPIa879rGtE6eCA7BC1wHbNMPPbD91UciP8EcfJuOScx396SI8IcJAygrBljbh5S
wYi1PHDuljkNR+Bl3GhLawaAPqOXa69jxOr87r136QmmorXyoe/ejfpM7LKjWuCP
5dGatorIPxSgbWgzvxOecJ7ZbDK9zOtxhfqmEH2nOCoHisuvd2wRVdgUSXWbDUcI
oF2MxUOfhd1AK0MBPyjgg/cjD4tQxiDRU7Fhk/bEC0+u7WUl+s+Ru7IlSgORtQPQ
Ur26d17rfVyu0ePppATHDLp7wh3/1uCthahKXgbCL7QPczcywa79+vCutdslG8Vx
HzGx44QvfuijbaNEl31/lOOaWDj8/YuxEbTowE6RdF4GlPiJNQ0kxK0iaaaQ6FAN
IVQQu9v6r8Is3sOeJ/ozxueZZpekl5pTVln9Fj+DaLBNK4rsDCyl0G8v+NSZcrvC
1xhSTH9wwMx4Gw82Vqk20EefFa+8jaVP2ndk4VxWSjjpeCRuQeK/o0Ai2wwTRACs
QjiTFXAvkcMz3M4pW3HeaZSNrv1qHWiz0R6PM8kzJZGBeqHcQpAT0ZnF+MHHvoNE
pM/X5xvc+w2j8qIMoAwm0/F7N0z36Ha0EgJMPaGCHSe/DkSymJOUichFV/z9VR1+
NnCq2bLqt9KJDVSSE8nAihMoNXZR0wrSBiTBI1JKoI5pnwP/Za9029hF5P9WQYzM
suZ0L/vHSYxxd4mttVD0CjuGuGhiGlAh/P5bbCSDbiUlMAD96AmYqtHcP1mxtSlm
uoFrX6pSw5civUe/ABtgg/z4eRV9DJdrs2CcLDnihxJJcuzZGGF9c07x9ScBmM+Q
+wTLpUiwoUHsYlmu5/vd8kAHcvGHCi4oud9lkWtyF8QhHoDoiW3fPcEkY9nzAlsh
lip9pYUBPvMiTY3pX68ZAKSuc9n5d+dbRQyvgayFfVZE0dWj0/vAv3VYBsb0VYLA
FaRgQgJfBBmmV7Fzp6hd4Y4AiDr0AQYqQgzEPDLJWvw04vJ1Qm69/7eskQ4+6OQO
f1hoBJyGVBKQFGJSj2eMBt6fwPwjnfmxEgB4k0+1uf4WOqXit92L5BLTTrYRj8s8
Nc+ldiwDy1sW4UZQfyQ2my7glTcHSNqq6Q6JdlEDwVw2X2D1QS2kgaFiIGeDlRGF
kivibp+UmotR8a1brf2HqvkicBU+um+X9i7uf4DYFqDS7BPyItBCuM3gKXLo8xdz
AoQtnozShYpI3fx0m5UEd74Ed7/am3EWvyhdUai6CGa2PpL1R2JlnxZ/YAjTBZHi
ZJeLuwYET8gcvB10lv/c1Ki0R/Nf4Js/OkU6+mT/xP7bwzA08wWBJbBW3aCff+j9
RWo8I0aEMpPPBHEZ24bU3nU/2wsVaw+cQn1nLmw6fjcsdVWzCmYqXNgeKS648MWa
uQCFUyQxU8v0R2zuTd+TDv/HiRBRaW7+gxevAk9xA5yJN5EbzIQza43fpIz9tZTU
arVIX0r4+I1q7o+k/R+TTXPgaG8eR5/B44fBMFsZ9M2FWq3R4WmjRNTbUTvtzEzv
KsZtoBH/U5P8Z+1FJj75jpnb8//68Yff0xRBCAuGTQ1Jch1kutzDHks2gXSuWxaE
KsEz9yp86pc3/ESQkwnWyt1K+/1nb9rxJxFK4tlZ5uSjFOZQHpJqLGfp0U6rZsTB
s1lSyU0Qfali980IXxx/7XpT0qr7UOc1iOSzPA7m0K2QkFL6ToJbHRqgMQQLP1/Q
5+cO5ie0tB5XpwTIngHauZcAatwWPGx8vtdZWOqVIQYYme9uJ/wLe01It09+eisL
WZ2+4oPbrF5nbmGTK4WHwicrS5BI208CelkwCpQT4K/SQlkowRT800Atl5KKo/b7
MDplU2BAx0eXdTnd4hARio3gNCoDZ+CYpy3wFlofu/BArwXGQFYpW4PchU0UXTLL
+BMvbInABSCP3WmM4BZvuHxuFPkPpx5Uo6tCXQnkJ4YeoaJbeQQlWhTh71kwZ3lS
wJ5Ygyh4UqEgrheSnO705PR3fpbvZMgTtHnUtnJd/5tbVCADFdx7n7Aa095t6X7r
Kqi+e2gh3os4tcSNyCFQzU0eKKBqaA4jETD2cWkHIeGmSFbYhzbv49G6MDLpFccI
Qc9jNqjE0xRCn0FLg2zdRFBvvatAlmJasQul5cNO5TcEChHNyU45OB/3uIW/X2pd
VWhl1OpGD9LyamuO7z6k6bPrz+IV1wWy3R+wEacBRrvrNNnUVFdRrETFP4QP4nD+
dvtvD3SCNzdsEdgkpJkl5gpQQtp6yamCNWnxcQNqAkqMSs1ec2dPBginUSroEgCm
aKBCMmEGXTGTz+/MGX9fSn2ChNPLxVAu8r5yJyWEm7ycc3hcVJ4T9pRBAiHySjv+
6fXOcBsLiW2H411fE+N5NY+eQw9BbRLqw2CXeHM1Ky5yYYH3+vbx2PjlPZobiwdF
plB0gYArNRU4AIK9HdozzTr/50sRhOrWDJcp7FVOayP/xPKn9W93B0VKWtUcodyc
nviiIvQ0WrPjFriwK7KqLf1ZlaOWQuJimwIfhZGOJDICUr8Tlyn+ctxdlTQ4Rne8
aVeqo+t8cGuZlICWQiBK/riUxAQCipe6TIAP/Lp0UJDL2kJb4IcxcF5To+uTPdAl
Vw2P0ZnHB2o50rFLrF/Pw8ahPmth0fAdhnya7MZo7rNyM3nl0L6A9s6vAoFnlM29
r+Am6CnnBzPo1q+iVQ7uFXO8stDZihZ8BBpxBny6QAWB+vE6gFMInn9Q2ZPQAWi1
mU4DG+8CzPy/mYhcATLRe/CPXJNvIyjlF+gk1D03tA398arXRRIPHOt9jEZfRYU6
soooXuC/PQ9mkQmiwttPr9LJFh4XRS4m2jmPmQz/0GsSGj1nFLk+lMF2P5Ql1xuX
9LD5Ix7R8QicJl6daeJFdWegr8xR7McIWDguW+/LICr9hH70dY1kcUTBReV434rP
+YBokj4PPlt0UsXhDc3xtuqeFOOuUFaIHFuXR55BARoBQIE9tavk1dmM+fgLZF0d
pRr0Cdqi5QWJ+Sn8pi8rK+hjE1As9D7HxJdcS/t+Ef527ZrDhbPPiFx8IoMIl0d5
g3IYWv3pvwXm6BqywP47aotTd8ndhCJ5TmuuNuQ/kKmM6HCirLpSL895m0JhVksj
d70RYWOs4w5/t3w/x636LY/ZM/OpJHXqH4wEKeWsro8CvGe2ny2ROXG+lJ/ILwP7
wMOMVuVWQJEEaF1IlzFr94UCtxZJLREJuETo76ElKdenxeFtCzziyVS9xVBTiYY7
YjV29AAzcYHnsBn2VyGTB4Kh8+9FFJ6b1VTqJPl2ZE4V2mNJNcdcuNz/Zms8F5GZ
ZDcJFNBKrmKADLFKMIv/QElDbQanjzEnlJi7I7KXrivn3BRMnCke8EPhUXo3JlD8
6uRwXz5napYdsSSlPEq+XUoT83Y67VsJaO37RwIa2nWSbICiQRe9pUCwH5A4HSAQ
mBLLw6uEAVCh+KBQalcRR7hoFIHwPJhU4bykX/A4DRHqfpF+771GnXBzKBKjRNda
xnNdnns8WvPabJvzJvt/U24nT/YJR488My1tdpCMkerXHsst9sSeH9wlWFp8yUeU
TAr/StzTXs62oCv9NcTT9hNwdIr8gzUaG14k+MfvJn/ICzitHXiXtQLdoLTOVe+x
Po6Wp/JPgKfkwHEZesxpZ3UtnF5Kwz0sXDaB6kodELl3eZj2DftVxt6KYkcPQqT/
0/xtCZ6FHGN4FrpxmAh5wMcZyMJFQjBxibqtMfH24Lqk21zCji4u9aWCkNWjzaYt
ioukrFPq5Rr+Y0mplhEpddDjvWEUyCZMzq7RFzFdq5Eb88oc4WL3vGw2v3WAtHym
gL1hGj7wutl68HLZ2r0cGgqjkGP5g8gOhV7e5sUsSZRx/hfRFezgsbk/i2vP3MP9
XQyd+uprm3f8dlmF4jA8MQE7koOpwsfNlXKmSKWv4E9agFLeMYAxsn7EgmRpd7ZC
Kf715L2ctHrUj3AiKHoL8Ct70TUguLX2Mj36gZSpQ/l+MuQyiWRqSqM8UW9SCZcH
jpfnk9025GleOBerWMefn6nAFHiaIEFR2KBdqKoguZSmPo1hpKEYXOhSgrYEiHMj
RkHvyX7FmHvzSsiQCdBQZLe0sOWWenmiuwDMktgdrAiMdVJmlxMSEfVglpHBBN3m
stsqZ1vG9pDAePuaoycI/6m7Di9ssm8k3Gr/bACE37g8z0izlK5/PxC9BNsU15di
TNdiYGwCBM/OOpr+K3H8s392AP2LqSguaVs4AxMeDnqd1CWU3IvBWLix9887FjdL
RvezzxAMfuz7otVW6MYdBEOrjgx/NakrW7SUCesq6oU8b8lMxxqRvuZ+ddB58ZqR
zTITQPcPnPoFW30JfBPmKS3cRSk0cQ7L8E8OKM8X5UnziHQhv6UU58nPYkUw00wW
JON126ImU+ApJp1f36k9EXgN9Oj9hSIYyAeHMuTO9Nqk2PZn+SMJmVs+Bk21h41J
bpsvZONm1m4QLEJBVIL/mZAzLlTqFVQAxhc1Mx5SaZ5jPpFPLtXlKp58tlTD4kAf
03ObwGw6cCr+Egvu+RzBBRPFtVkkbIwcNnGc/blRw4wd1GlaBlfwDIo+WE9QVnNc
VVxVXWFqYre0AARi8mBF03RWnvjDMagLKDotHOCrFMsZcc3a1OgZm5HKM5d6ZGOw
Rp3krNFiDVgylJRJmak1//VWB9TmcmrGpoI70+FohH2skErKN1wcvnor1A0kFK3m
KBYwNDOstR9op6ZbdWcSsE/dkwV8qU9ndpqSNe3sH6rTbrotqRX+4BOSEA0oyxmz
Zbzv2d1VI/mzS1+2Fu0455Y9PlWoAVgw9YGuTzwIMug5sriXRrj2K81TK5JFcaq7
sQxeDeOkwHqoNIXeYK9WTYq7JRQs70M7UAf23X8fOKhcDt2SUEJVy3FESapT6A4z
G5ZUZT6bta4whyCAmgaO0gYEExfisexweBXn0TGctK0gLJi9wS7rU7+fPfZBDGdS
lhLDm0ICst3R85pomsTKzz38xkCJr90U5miIQY7XWqYV5T9/lSMjz9MekY1BlbK4
qp6rO9iMBca2gmXUhaeYDtpHHcSKVUDo1Qx9iIeQaDobl20LMzjRzleR9O0lAPiB
x5u5Y7OnHwG+viNU1qtvDm7cfffrrd1cSENp5YktzQTpgN+VYyoOD5/97e7laEBd
hl5LaPjvGXK19QUpTqBziwxzTIQMFFDhRgA0lprv3wg8nVVpwC63QKjti/9cFFU0
AlSVxZulFadKofyQe215CgKLbhhwlKQlgUnkr3p0WR6VWc/5qY0cGixOD5ucneEw
pRRsAcejlHTij4DArAypfe9glTpB9Dwx3692mAjFykdaNe901MPmv0D238OBQ6Xo
RMcVX41Y1MpKB+RFRY0uUBCjjq64mXNGWsr4gHfPLOOO12hKvaRuwRV3hPXVQeXB
02APLi9nJk/+ALXV1dlOOyFr+k3Zo4bCYnMVOEKjLejX4PpzLwDbduU0ZtAMLrcF
p9XphV6hBLj+XHEniqQY8tUW7bpwEh7nPu2GNTr0EH521bvMWOioqgKmhxCg8L0Y
ky7QXvXro9oW5LuTWXYwdHm9oOkUVsBV4XdylPTteLJpbQxslkiD0A5PStv5moMe
DtdOOKpJ0pBR7pGMvmawQJFvRCJGedoGt8zWikz43JzW1AQkRJEP1L15YoOazJm4
KoHWZl4cZZ1bOG6ACvn6/uE4KIyJtLM8XVRtCkdPROaiAvFe46gxTD9gmU5wjWI8
VBsui1jX927wNR1y8BUfi3qhXsyEz5VcVQU50x64f86k8/byTdjav3XDhS8jJnRT
tmkTgFd0ciTBbcZhuurm/TgQujlwVEZD2amLpYEEAzbL+cqtR+XKIzw2Cbq9wSB7
zc2sM65zlFvPv7c7oH+o0raANSH6z3Pdzm4vXqL9wgfY8EmBqmOLERBEdc+jKvim
wJLBxLrgW8FeKCnDQ4brYBGWcjwboOCphcPlz3e7Px7dJlrKIWCXoRASaJcOIEpv
aYzK3vAP2FYUGbOKUq4Jb6Q8K+bP5JiI3eP8hG2rQaDF6n5EGnbEgg758X5yrdLC
SODgrZ23IqAbl9JmyE618M/21bVpSD/jd1FTF/cyBp4RLvJ79zz3g0WpY+3HTo0Z
+pmbrT6XqqVlm1XGhok8RuYn+3gOlLzHFA5ukdPAsUbkyqpii6TQHgsTVQeTkvMh
0rmO6b/0kInElAoN1C53x+0evvagzqLwIN4m+82ghOMDIrycdezHcX6sjGkIZa4X
fwhhzEjcoHfm+K5BSEr3cows2u/vC5Ptd3dMMXsHfTzRc1PmsYQWmh+ZIOS/xppZ
9k/xGBhrz91nfQdMaNjbW8EsaVtGBrFas5cWgCZUjoWsUNduy4mogsfqCE4D1q4a
FYwIF2IO6woCTiWTtuO9vjiwsy3os/7/RNhCQWTS3H/Pr6M/1lLPqvPvwbdRQ0tM
YU/V8iSul6DwBc86NuhYusRqoulS/Noms4u5wbSvJ9wyRyHzDnlb/OvafVWT4k1q
wlnhePNHopPfnjJSs1Gtq6uSxxde9c8X+zPXb7n2vtuQQKXggLMsHEXa6Kb2vmWX
c4jalSSyw1HtuypIWKCXvmJNrut9kp1CzPjeqYGt75a7gkE5VVTrF+/DjL7ZMonY
+/5nAkiScGTeeFhle6njSbRSvcIFkTDkuIz7jLM2e9A+KkkPuk8VMBAUq8+PBkht
d+tjE3lu2oI2XfUhH/b3hYG5baTxi7qCbxRHcm5XiTvj40hlrRPVsXzrnyJxWbB7
Du89jNYBtXKLV43C8Fj7vO/3d2Y1eC1qO449jBHy4wNG10npaYIaye4teDSL+Jk+
6WZ4xEpypBXtg4U2ItW92ix6OIE7JkQmeBNi3jGy52TzKt2HgvOLVJvLEMVCLAS0
qzLvNIlVAQEoA+WOvJKF6zVWpy6bvNDs3s5RL9rbXSRe5aUqIX/Tch12QMYuwi1M
CXc9wybbfjXqDLLiBCSTTCGM13MEL19NHh6/G37DQnE+n5mYhxl/R2HzBJCCvWrY
s1jN2YOzniXZ0T9l9W+O5Nj4VwtW33DQ8njoNvG+QUh0KIcYP1LnzKLsCepeHd/a
jkR2XwxfXmjbX6vYtsNGVt6kdhpDh4AThWMC3i/4wwZkvoeNn6zG+O4MyQ58LQ7F
WZKnK6kvIyJAfY2qPO4XfwCFaIr9zNwF1+QgbskI1cW8J9Sqj4bmYty0lrOhpUrG
t23lc5mCForsZcEnCcqKxRy8Ura914WpNcFyrUKQWafMSoCoV3X3lD1JoDvqLYOG
KYldBTQN1c1osGnb1yYSyaHzR/H05JaC3e2LYKhpUUhHRrolvu3dVcPnMX3vRaPa
SCeuSa2cqLIwC0xBJizvGk4iM8TzFNL1FEq0SN1KVNXiJ821fLTzCulgAoyJTZXQ
IPRo9Fx8bbXvqyY+u8v9P0ZMw6qkgPIIxcdHfii9VptNeu8scAOaxC33fP7jWuER
Q3WKYPLWK36ODJ4P0eTXzI3WZh0oiwYEcRjSfePvrOs0NtnVPwSc5CezuDC/kUQ6
v+9SKKlaNy5qc9FdDlCXUrR+g0nbQtXX/6ADg41ECyMToN/TPKQEkLQIdmNFmTlF
R266FjJHKUHCOsYcN+XRqVqEHsWs6BUozANirMQMMEN82vxrvu0hgBsAIGqFKaMJ
0Xb2qm7ZAh+Zr5iJi4t+hkZKSxj099MIc4yU+xFsh+CFJHGPE27r+Dx+kyRRLDFC
deTDSH1ehhSiSg+m2cdEYPi6IELQ9Y+gNTp3MWf7+RmeHSi7XtjncUy+lgviCa1h
aN23FrAUNVrVDFHuhb4MhtAtTJNdfklyYD8V0EPBI2g6hBeKyke/9rvPaCAZYHJH
CJloIXhemKBb8h5nBeocU3MA+pnY5r1wyLSIVAtm2nAtg9llS6S2S8ZUOuEzEnUY
N1HRZ1cUVneGqHmQq7CPjTj+gCgU/gVmjHkBDHIOvZe9vrXvizwVuV12/cSQCr0Y
qAX94pKgMwZ8TYGznqJS0Yy43jxa5QTww/eP2pb69guGYRqVymvycTFrk9dev3cG
NTJwYYsIr6EuzxHr4uditNJb381rELZse6jhsVtKk614VaExuS5jRbzZep4zCA6+
1YLY6ui9BKwVQ99WV9VgnNxI3lMsnCb1uT4y7AEYCti09fqhd3m3OeJF58WnKsBI
9WMeqp+fCcul9daECDcV1oY4ICXomnaqOtWFEtgFPe3gajoYKwOP41qU7JZSdCog
CggYp9yjHyRBaaTEdHSMeY1wUcHg7QBU/+db201+z2tavz7NeYoC6osx0k/Vcgpl
4iqrfOEiMoy1A7k/6yPKpPaSC/vZ5ujLwXnip848qHOH8iBnvGM/ViKxoosxkHmq
0Objgp9rbJeBSnh7QolgBuKv9BMpqRfaOMhd80pu+CT6lPOIwrr3rjnJ/X6+Bnyo
+2qqAL6VV54FTHWYgeKyrRhq44YgnhjY4YATgR6CzkCFtIRnW5gyR1Sv1evQ2d/n
WajRfyEq89ZCWWSr9BFdewAnQXZWAbscsFegNV3HeKj2llRDvXjxXnoS05UiK9Nd
eLnanjTs6tHamLfp4gRuRltjNTUfe30D4ZK/tYUMRENlBGksUKRRZ++U5UlVafUY
p4uUaB/oXqY8T3LSzCBlaNKaitykr2d0ga5+E7eQ7I6yNlqC8Wo3Bd8KsrFHlVgm
QAbAmJj8qT2W3YStO+seUV/NXOH57TDtjzqlzW7ztSs1SMLsD+zlENywXjjO0fIh
8MYXnAI4CpOH2Z4nFQMYqXyelmeVPpFEhY8ZqyKCyhre11sVLMT8U+yQRGo0+1+B
ttpGCrRPg3zebzzL2pVMem/SPNj35cIpm9xX2hFLfS1hDYlt9kNwKfZ9fDL3tVG1
JKFI1PbAYsrG6z0fHSptY4lApr8lp7Wgh8GHMlHE1LrslF+ZS/l+zcSw+IxZZcNX
3we++6h2COz90KJfgrJSGOKdrgR3SuNOHO18wFvEfMT6HtV0yjZHyYReAK170ebt
nxDoNe+L3oWsIfZsW97WIv8epdJE1zYR2bWkEdXqO1AGWQ4cNg+7qGqBjLzXexqM
e+dioSQme1JpmX34zUstwc2POeDqszp6cYTO6B1BycYDuTnVHHnmygRTPUPdlMsk
1K5slH3VujUCQAoEJVmixiY7C+ibJLZ4q3sLJ3oXswb+sOk5apT30fAnrHB4hvAj
0UDhanrNWgzmbYDyE0qJcxq4sM8E4znSnNUgYDVTbkl+YpAQi0ogV28EGLj6QLb6
E1oGiLWPWGoB6Ld+lyZocw==
>>>>>>> main
`protect end_protected