`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
+HLGyj50Vlx2V9EGPjlr08cAIudR2TQw4pgjKS/0ANH2nkQUxtrOUP8iGP6nUaaJ
VGh2mamUER8KAuiFsXKEg5EqFufXo2YspdaM6M01ihsvwBQChghJCRDXWz+cPeWh
iRdRiaEicUm/e5022pg8nigUUMRSoV/VKo6asXUmjrvuubTcEqAYuuPoCdA9dFKx
EJL36GGVgDHoMbUnun92684KhngzdiaB/tt9gHFKx/7smPPXQbIXJBVL28z+IbiN
vn9XaDx4qA8V5wsFV7EurlzGsFdHvTtWvBCr6bPYzN6/Nqmyo1y4N5ehgYf5qUmq
qDt53Xx9XYTb+Y5nuPlQr/QgH5fJ4QSUTRTqwcKkunAFsqPX2NKvjzT8qVWjaQZW
dfwuxgA1c9ZmytGsB7k/z+DSEpXwCEAC9CBhJtjuIJsqsBOFBa0Exu3kFK0X3vkS
NnwZzBtfL5a18UgAl0ohzsNMSOEQgGC7f1BumMHefEnoN51XnfSENIQzwvifM2+G
1z5WjsoGlfWtYYYG32kH9w+nihFwWJ1fW+kQ9IiXTp5iijsY0x6qN2dVNi7YqSrh
PhRaGgwwG71tskZQ+oAGkBzBpwbf7Le8OCRI26LbC10t8OkWszx01+r7ENu4dFq9
v5JDTtDoDlXSls9/08peRiByfzw4QmNcXLNRNT3LE+j/dtL42rDNKPSfQZgIw3ZZ
sLoKzEH3+nNeJ4OfWZ/3hpPNdqHraeHe9U7wWtrDXsyHnr1QxGODaZB+lIc+8wy/
caAb4aOhNpuUsOJx0RJQc8ZdBDyQEdvIyOV5tDnCiWb2RskQB1q/QO6eH6aS0tr3
NNfmbvFYd3M1m2dOBjKsnYMvJlxjmaLn1k0c7vzr6yqNQ+J2pOEGjTkpuYWwpJsI
//dUsGM41l4u+AryuhPR2HAnDwsmn+6MvE1+9I3qWFjq+y7Pw5eDS1UkX7fuScEQ
aoA8ihIoWTqrrERUEvfcxD5AhS8PGT5HbbkvEHK/bKmj2ScxQazWheOmeywC5VaE
Pq4oCtbgaOBoky+1/W3VCjirLJTp01I3n7lXy63RouWhm5WZWKv3hnOjdAcOmJ70
9jhXlQLFjT0PFelBU0x0fU3Ty96PtCroq90uUx3wa+xh/cxFChBwnS2GvLoZdRCL
AWLKR9sPYc/HITKQvRb9MX13ZiAZ+XalyjNlZVn/SRoXlczaLNrY93tynBUEIEGd
8OYQ+iABUliMxbT1HBhgKLj+cEbnTP3vPoR0Kh8DpewqO2l3bXZnQ4a/E5vcSIDO
2teMexupeaBd3XCX8Scl0IlLE94HXo7rptFjA84tvPm+nmcXPj2IRxEJlp/JPS+2
Kf0p7SRLTFb1V3v/07w/wZaRiG2h8BlCISZzM23I4oH1tHkSX83j7S0tVw8/mQx8
m1XIP6s0QYLbAz7SOhpHwSJVGSXCCTOqlBBBSVDFWiWHa+eOK5KzZ/Ltf8tdlDfk
tftfZGJrMU1l1/7VmflBb1QEjxiMLWOxzuLcQw2Cr8VByDbVuSnc8xJDGMmcBk+7
NqtHXGbz6h/sf/zKjPqviBEbmMMnDIW9TKXJl6GqaRoSLCBR/1rXy4+s23K2a8I1
K9gILQ4Xs/gSMo5Q5pMi6c4/+MHE7He3lYMGBtr4vxx96PgCOu2h0TCJzMIm2yRO
/PQNOG39yK1c7Mt2eBHluEpDJjjHcSAfg9jLhImEoVQShEQ9cf261Q+zycZ2U1jA
w2JGMs7VALBJAb2znh5qJL79GallRSv4V7GbEluDUBgFVoTR63HIg/Jrod97Pvul
M8hL9o8VqvjqJITGVRmX4qOBVstzmRYBqpu8gtlh/BbZtAzaoZ/Hpwj1JiIinSHk
5SvAkk9/fqVWXHazBy9jM4pU7KpqnBOcKWH6//DL7MIxz+gLYt0It3M5JD0HNhZD
G2HD3IJ655r69c7UWRywRlSwJWvQjpNUsUEkwnSFLe9G2Jhc/nRK3eL7CMfzcka8
Se/ZL4MGkZ0QVg82mrkqAPegBIj593yoQkDC5RQuiwF2BJDGuGe5gLH8OVg9K629
JNf5o9zNN1d/FfK+HsEUurrR3momsZ6qxptYbCjNvVdpGRPBuSedgwR9qMSyDDSu
vCtrbVLjPhZPOQ/UzWeyghvoJhhQwG5RpaDIK+S35jNPaLjg0f5I0FsTIuMjDfRo
ViJx778sqyXz8IUXVEuTN4UC0SUsXsx4aV8eR+H1vwsHx4+BxwihtA2Qk8oCmbJk
TgC+QD2TREfGEPZzpGsGZFIJaPKOPCHxzxY1gFulrkLsW5h9YEsob83NXEVQsDAJ
pCWTzSXP3/WcAm/qr5TU4XCOjAngkYCNi1xhYGSf1UoY1hHPE9jxmn8byCoJjITg
7wmcfqyRPS5LBsLcupoykMQYRVHcdwOlHt4JrbR+pYQkpk6P6rdm2sv4vsGBMaUO
yVUO0JKZ++GYswhU9ExhHMpbN2yHp/PUor9dVq+4EnKSHmbSf1wRFZlb5IwVKBlo
fNeFqLVUeFKBXprzLZ3QFOyj0DbswpL8yl9pZuxZwnILPtr+b+zPT8+qakJdKz6W
FehraSKpE1Dma0tsJ4wlU5+148NjWg4MEtjB1QHCOQ7hkBxmA8iaU5iOqLSPhr99
1ktepW3lTTZx4YBUyTCi/OlQ+8a7CEwjTdRyIAitz7KjYP0sQT3jyKaQQAPW4aWd
XnVXC/OCzFbwoDwcela9FTuyKroUbB1u7hnTtB7MMbuxEJh/hykSobD50c3NCb3O
UOIheSkw0GdCLWnulJUHZ+eUzqLnry8wtbp0aRGWnEG23VXDJ6mqhxps9mAockon
Z3cDnhiwn/X4jRjsP/d5jHJDXqG6OEoDXn74pYlQ7b2juNiCDRnISSnq60ECeEk7
ujG96iq5NMVdp7nwSZPUiv2fBLXNkKzBulGoRGSqEc43VY5WY4WeSECYfKkuWZV4
L1Su7qQMZ1t0KwQbensGmePTxPI/PAIyMdYhKgvuMp5uCskk+WvVRCcBcbXpMVql
lB+oX7EqN1QXamH5uuOxracgEbj+Z9eCYw6MqyCRE9OK8W5/QMEXPBMzH+tBn1My
hQpyTzDYd3+op7SDIxyV7EOS01f6BwlqQNczsCR/ppGaKLIPyzXB8cW+dJ9ibYqy
SbVQ7a4yeYz5mkLrtBw4PgsjqawGPBgL1DTcQeV8i3FqUqKfgbVz9CMS3PPQu7mR
yoFcQmLTz1hAJTJNQMNmxT1B5sQeSYEVTBQiNvkn2nyaRLp986GjzhB2REp4ivQD
9mScvBuom8iicZ+Dp1sNjvaVz+UBDkuq5RZkeB5xn5k++p9rALcQXIvYIxB9HeFZ
Holfx/yB58sT5fHmpfMgGh1/vJ9VOhGUW7//K0slcgsv+Fq4knNeXS2GjPgqJQ7U
swNl0hyZTv31w4m35M3ybEIqSKqdyXcptpz9fOw7lhDi2iB3BHRGGLntxjQEoeeq
XeyqH+1cUw2ymVlpc7gDRqy+5zGluGh8/vLrqgXHGAvx8W+7Wz6EQiiZxM+0rNRT
t3QBIqo32iYR+zRXAu2VCG0iVFtcOh4OZRDrvGldwCKwTXp/OSkSPufBJpARx+/c
b5knlya7dCqpFmw0BNqMsCNd69OP49Si934JrkR7ACVAcnI5B7nE0DwU3pLIrLyb
D6+oYe7q4OAjAHsWKX2PycCeUpmVpHOT06l++UFQjcq3Qfd1kTQsWjsXRwRgyuaT
MPmdtWrS1efN4wb+09utDxGcHSawBX6dbV9E9duFTERuYrT77P1X/hECkYemqymW
UMnAygbg4hd+L8WoYUyR5O3/TQglSICtnfpHEzr3/E27T6LCp8Su1P15qIvEtcR2
Q16H61Ktnv34l8Yk4zcAi+6tpbOrnTwNTf+h8UNiOHrYcwabEIqkJt2cXzLulPuT
OYiUqZXViqJZvwy6DJ1zHX4pp8SjiRDnzDHhCcPVWtCeEPa4iVf+BRh5XPuWsFCf
IEwdCwdcoixw9sJgC6xFSosnKxEUXw+aG7YRkB1Zw30agF6M4TlSnyihdpvufATk
G2keJAT/+zYw6RjBuLvTQhT1NcP/0nIyK5s4D4GaiIJ907cBBXtLvJWF5tCXiDjd
UnC1nF8LS2weaC8+TT6CGnLCVQwnt+cv7APebS8Tyru+4OpdyxL0TBjUkEDHOhY8
tgSWNxqvts8FsE2m5G3zvAHF9oif5GsWHLvzJEwTuBA9NB7bcbQ8rmkvK2Rd2adB
JcH/m7sa2Hyrold4/SP9od/U8vuSWyANd45d+0plTNvUwEjwJxHAOh0y8LYxQRee
3QJWUbKFXQ7RQYMYbxuKpiHho6+jHoYPBRsN5emJMOtMi9B/dh4wLtkIzzZ6sd9O
dlQp/h3+7lw+DH7z0jzl+EQI6rZlUcdT9TyEn+NpEygbGNARvLC7yzVBG5jkvo8N
yrMhMMfLZIM5IiVI2nAClYE0mJzAO01SjLj0GmNqQz7AKdUXsP6Yvmc8VjA/+eGR
66yNAbCKSpG9tRjL8g+ffaiYzk6AutSLMoAmaGoqE3rri2E3vt9hiJeAD8Gtwbvu
Bv2IyGLigI69IP8jqxuNjTz1FS1xkJtvg35HWqDq8ubzGwxIebZSqy1ubFIYoBBd
kveaIAZ4vw/Upzr1xPaSm7UT0S6k+TZhjlgRhBbmEKAPBmu7hVufaBeCR8p3SnIc
TlLArsriTOzqNCA4fsbwj265xYaR8VCcT85NRGQF+js64szvhMCER4EOtpQHdBMJ
1dV2qEttLGDm/txPcHxyv69BsU6NWLdIc44yBqWUXuTQgVd+kf7tmLkIArA3hlW1
/ywvQfilCRYNSTbmh9sPFD8mkPd1inrutd/rf8HTrQkQKRWMyPhctCHTijfjt7up
zy4g6JTDydB/7KBG2vx3Mz/tFOW9oWiIl2pzmhrHzQxJVekxBz7BtrUiqOBPNLyw
glqB3bsovgsgKfDONxsOsXMBqU7MDeF6wsoqrV2S30eT31HxnJirzaTxyrhuIPb/
2YYKSFijw+el4E/1hjshdwX4TGeKIf7K4SkUZITdIqaWPpobwZQFtJUiOavT0IVh
IKJAIYElFJaY3KgjVvH3+FKm+/2A4ItLTMDn468aal6trd3cB9nfdmYINCxMPmWC
PS/vLJixqiKlN7mvybzXGe1q38gzWFUDd1LFeqZ45zMrEjvDiLHUMmnyVrQoCJWR
qmpdsWhyvB0fgEZnzdbNYV4HuvQK/N79ZdEPcPN1i6oeCqLt7Z9pQZuqbKNsyMnY
bHYUS9JswJpSgCtvHWDX5AL/IaPEnZ5+M9A11DEu5WmoY1ZS40E4mclcuyXJMlEn
HztzOcaoqjulxznOjl6HYGFnVQNVRxMPdnxr6AimHjkBoIHN8CAs2ltWefG3GbDY
zdtoH6vgKslLYZmsdlFAnY5JxY+blOexSZlk8BKt6ZWOghx4ILOPyL9DPzVpSgsO
AEzqMkeXd0nFfr+qRjAo80ZG901Bd73VEwj+TvfzPOgBKhmNico8oAi01X+apWY8
kbr1bnmEI4pc6EsUIX2q3Ku/a/rKg7NxpMTj4SBmPeQV1gGOsVyFl6tAVCQFJr8H
iF2H1y7ZGHaWHIITgu34tgRmVqNYp821a+msOlIkMuDy+CfkOBPpLYtlqb8eerhI
Fs4ULcwIILEbwFufJ8FGhyb2Q069n/DsIgXwKdq84V+XBRkucTgoDzx8A572IQKq
CjsdVAf118sD7kNgBpLR13alVEUfGXpSBekK7JBD7QXY4NIfSIe23BQ3powghoH5
mbYSd5PW2fWtIHJAAlMdOQRT/nVDqlgyl96FWEye6rmPVKWO+IXSFkGBHYehvwsM
FBwK2e8t8ns7Vrs17xJSkM3E7+yGcD3ZgaJsYaFjp4ErvWJ3iRoaQRS6WCtsEC41
XkGCk3AtGZoonRQkWDAUZBke0+TPGvaMK6l0IM1J4F6DIbLfu8qsevJnBFg/47bX
s/lJjDAgRDc+hAOoBcdicTL+Dh8rCQq4noPabwlbHNXxHtV049byA8UIhPpQ6I0P
VOCGJN9at7k3XP6nZnzWIsI0pRUV7WXtLZWyG3ZKPTEeID+zFTG06F24ZwfyLT39
nCdxDU6/g4It49p7afwN/iZ03mHOTuFMn9fysyVg90bXBSbKMrJXO0AnDx/4eWeY
E6yd+t0I0L2cU+2tEdrpAbbDR8EZTFLwlz/EaX7nWCKqJk2d0E9yu/0U/mj7ysU9
ao8KJV5wJjUbujuBV3Sw2rTFGz6eyGCauzUDGl2Ac0rWjD2vi4r/7tj9xcFk09UK
RsV1jaCOU4o+S+nL48L7CjMWn7xL/DU4x3lSOZtLVKf7kkN0wv0qoiP0rqMB7hdW
4A0Un/1kzJwK7BDzPB8ayqxjmsyptki56bKhy2evvdIbfuYT4TByLZdHPG8Nrltj
ZJ7nN09Kf6W9k6A/nGHXKgiqUCtkl4Fl0/YvpnVzW9gHqA4hK4C7usLL5vVbqnOQ
yN9YOrygeuQAfMheqP1iOD6+9aWvlu6nRlMN57SmW3e+D/MjBuf3+zaZz1mwjjtB
8JHnDDtLRrdDe8vAOOXWHkdCtCgoauxACxbp4IHHzrOL9/jT3zoNRxoVepOpDGEA
caYfwO9gGFzDfKSlglJ+3pkP4JqK1sUK2xzf1+UPI+f6L2B19eqSj3aoNjh7Ynxa
D6ZI4P9uoWOmMsjh1n2n68CYF5CpTfQhkbp+DnowQ1/z0HCJlaTiwpL6YKeopGzj
QYL+UICOEhBRNQspF2QxO4BV10KDMWHDPG0QsGQRZ2xf/kfi7ZeIHsYf5OnN1zxu
tdHIzMCj7l1MBm0Q9GNJNFhWOOW4CnR/wD/PcINw1bnwLKPvx/6dVZf0N8dfqfpT
t5f+GGpHBweUrqs2JuLZK1aUkJBseBY8vN8RrWDQLw1g9KV1/DcaSiokdEQu/ghJ
qJv+qYiTHUAm1aRBCEtn1MrcF71bAt0WHnof/PiwN7WIAkE7QF3AAAhHEDiAEGec
9vXVokMFusEg8SsmV4hua1vy397ZVWig8BLspu/CHBlVFA7alY0TImqMtXfN7yiq
SRfqeyW7woG+OnfbTcmgclpSPhZvWgw+JcUlKqhG2mXvOr54z3DPE714YoVa1p0i
NGvI2MPtLX+zmIy5C110Nt3J868NRLY9LQSOuZuJxA8ZDOV7hZ4QGGBjXFiXpnEj
jYDbul0PxmUBhF6TdRRAY3bgOtKoOmqu1oqjzLHmrOpBMLjtaOtj+BkY4BSJCp7P
58zsapqEwQKCakWuhItixsQR5ucPd8S+LGraqBynu+LPCAt25AT/f6O4kGtCYSoG
nz464s2W4kbefPsWWlLK6R01lJrrCDKT2piH9oFQG/vM5Uwo4OeQKKdwRSsHwxMD
p37sIr/cDFFqCCWbZa5hZvxX20Osi6YOR74gl4IpWY/wBInDMmjmSWwvoN7kjvGD
6tTK3FP8ZQGXP0jl5ymis5YFWWKoHmc9iB1UrVDufA09yQHKFmDr3pG8Q3gHPG2I
/hBhUBiP/rlIZCOeaDZp2YHEE3xZ59lD/uuae2vU1B8/5zMNoOJLKK9Ix/VcEN6m
xedLEI5+L8ExZC6nMuJNYOYS6qo5XpmdQ8W4TDnimSohrB40YCeh30xNiPqaV+hu
So5wdppZwRQTxLgCq10S4oEw1u5kAPkH+/hK5j9w67gl35IpwLzxsFMN8G4nKNp0
RxzHcy4psZDkrBSzeONtwJFVUuXFcLl/v8MYhC70qBFjWL41aBn0Yredxsgcjh8X
TdqkysuRxg2VY/8QXxj9aoLmELbPJIx55J9ZLbWoBGRjygeexkvSnWwb2z7JXM0x
ecxr7lJKY/9j6n8FkWdbcmTLf4bMMOndH5OTlJ1GPjuOwgQWei9kh9Tat8f8yBIR
5qjBHLrb4HSaK5Ty1o4lSBx6Y7exUf0arZN/EtGvsZUxRgJM02OEbmhVLR8e1Tqv
AZH8AUjPEkHXHcanQJ18wfF/C8gLcFatxdffO9GDq8WomozG6uunWALwq1HjbFga
vgDRvtscDrhjz/K7nvjGSDVD900SQlpZELHsUDqIb0cGKLsR6AAN1MJGTCUnqyRr
iNde69V1ZkjgvOdhMi1iIrWZhCWhRHl0lg+BVXSZuy1eBGL+CelPOWkV5eqNiqoI
8yDcEwWs0aCdwyV76x2fg1JI2BjRxAndCz1vfY5TbsspogLI22CNFcrtiL9lVyxn
EIi2GG1ootD3vkh8nKV9OHAcfCciNPxQ65bH4Vf97opWLORyJ4CWePtXNnwxQ0tX
QYUP+x5SfVtzSTEO6VKFRSUuCjMuA+1dCvxsEOjjZLa85p5hUUf1szCQFKt675GC
qHT2ciEJx3UWHWEGbUUnwL7UgWUdlYxLvMszaJ6xPpeSexwmufUjAoHoFH4g7EXS
p6T1Bky4Xoz7SRdW0eXpNPhFZqRCvn8zjIm3Z0tCTCQ/p8v83j2gAnVLGhNDbEc6
FLxa5nMxrSWKYQYt2n5/jVaZq/vbLcl/ihDRBrQnlx/GOr9/o91m9sNxdavM4AUx
VikQrKmglZ4a5itaj8bP0APT0Har6zHcHr4UTti++a8t7xQlMllXo2S67bwNfkdW
QnXWf2xZ7ZtxmQnMxn9F1vhxYLQ18cPceGCxwUJpLZPZS1jqmO/0+30/Pxw7cZzW
byVYfTxFXoz+ltYouVWUbr5VbQ7zLi3xZyIs3ybKzDZHoUl6Mog9GPI8MNts/2Ul
for/NnCulAFtWQTuZBMQiDhX+qWRVaRglt3geWVK++AbiT28v6oYWGpR9MBTYpe8
XB3QZP7AhHxm+2udE9htpyhFM6XxSHCPJ0zfzl1ILgfDhhCK3r9h9SWyMIZF3hFS
AYepSvPOM4uCyU63sXE6n1IIUn8iKdAYefZu2lkIsAWvNuAJJwkNd9wLb2KRO7Se
4QT+9HFIjIbl1OTQI5ZXGH17CwpaG4AVdk2vgNioC2SWrxB5ph00wqs1M3Y4NSRh
awNy61+KS6hBbOGhyfvH3ezX1db9hn+MosOpD3BZcgbql+gOBgELCIOMuubve5gB
mNjL2QbxAPQ6bUhI8MIkAGy/ziFqamhSNkAfry0axGhx1OUUEESZKFpWuwTX8YC7
8SkHjaqpDQ2wCXhos09mbhUchr2a+j1rJrvzK4c8bkUbylf2ObuQUgtyviHtRRmv
x+EkY/epELLvqopiITpPVGNpl8vV66BLMwpFcSoG8tG4cXL5iZDX6FiE2lhJ/ezp
8ndg7xTh26k90GJk9THoSwgh81KjL7JHvE9IWa+7WH9qcAHHmt+2AIa0hex0Uswc
TOafkp4VsPF6dnWkpi41g1+6ADSHUBY5LUzuMfVINcSX9ngwEnUjUAObLE8/V5uq
cGfHhQzLklCEX5/0KLupKXe4kTfL+vrQKF3N2rGo8ndJ3J45ppMk7DI2LikkSqgY
H/fdl5uHSBa2zw25xlLRopgmo0gR9hbzk/JcfU8wjLeOr16XmKfKKzvf0kkguCoR
9kLZxmZgzs9+u7R+f5YL4qlGTyxoRRZBDq7oF8I9U6cFKGjEQYxhY9mFFAccnu3R
KFoFzRBF7fkpQ9KIC6x+pW3DUuG3dA99lu/pSyEtOR+pzZ9TuEm/3VVMmteXGFeE
ISznJ6lhcSutNU/j6boQeUkUf5FJrpCbmsVV+FlFnfkxPQL1AT/VpcON1AQW3krF
8lwug/NdKvbG83nkgev9AUQR1RZCKpzrFBonrAQlhZr3LdF1TvmbvAZTj1idO6Au
H6oAgQp87PkMIblPGB2VGrpMT+5jZ79wJHn1cKiYV7X58yhq1nrO1r/3S7wKtewc
tIsvx79Lf74FJ52eOLT+NOXPqk5W/g4XSWl9wQxiTmRe2eWAWvBoDG0+5pykjbIB
7CyF9bD3waDeJ7Q2aeE3uzd0/CVNkxTXaNTo7jo4nclcOO1oI4ceIW8l7FBHsjLS
I+Ic0bkpB9AxX6C4L8O1Z7wpwY5w5zwhFDzfFGyvyz37EDZP9O9TSG1jP/5BpypV
MUTVlkVVWRgNew0DD8Dwxouw4Glru9Fqk9JIFNAjYCBTOmMgY9HGhvFS5T+xuUSf
j0GQgoiAihgkTBeI4Am7ur4bDCaa+29iEY1kIHsptZMiyoV8QqcLWsoq/NkTJQjX
izK6H+7OTSjIOutl7c71OHHU8/mdpqniYxf6FUV5ouJcjfDoSuezj/TqhC9o5p9Y
RW4mPmCkUsKZ/Mpd9Ajxg4mZgt60MAAoVbLFFq7dkiAIJHbBb4rx4XMKK0KK8Ftt
Dn2rQo13ueR3aXNjswWg6w5YJdZEXXF3exMPfpeqdimPQ+U9ar5qq6Vbx6iMAPQs
dOSF7tMmA45BHAV9pFgVCum1gNMhKVKJJlY7CLa4+lPY83jx+sx98wMaGHIntSPG
YNpyJhhRWlKv1aL6PXp6ISH+gpHkv0VpY3apIl7GcGG06fT9WxWsj3EZByVZYzAS
/OVChOqbSMjAPxSz+ZsDSYNzgMlJhKiezLZR5g9NM3aNcmbCmsWL4etfR2r5xSdP
J+7vP/U6jyHFo/X2K1nyBDiroXBLqD4myy7yimIXPYM9Nf364RmYMZHdjzPwpInH
zK0CpKPVDXp2f3sdoUsiYeeOM6CaIZT+75bAISU1Ag0x+7qAkRIXsbueIxlv67n+
2E2mA25M+hJm9NMSzqqRrlccQftcP8KDeP7asWARSWVIPPZG/Z+UK9t9NQu5Kvnp
Wt6bmzGXFRh7vV7CYwG8KfcPjRlFTGB97GQqEcbb5bQ90G0piJvo4w77HwTKp2Xz
5nrhkGzwpJaeOw7EWRAAJz/LsSB7FXceL+uvHlGwQadL2MNKMiIOV3Z7bdC+VUkh
/QX6tNbduZ6UIQfw6Rg96nnv3gP5BUkG3ulPd9FUO0dKPyAmSlfmAb+9KbOI9VgY
OKwgwBYJYA+YlufIDFYucUL4aGmrYbz7bRdfUskvv+z/32Indz0wLApw4oat1m7K
UrTdlhbrk69xz4ZIgMnIx9wXQUYfHZfABV+3kmRnZe5uv0f5MPmQhJzO031iqcr4
wQK96FNvUBu4eszOTjwKvAayCFTac35w8QGH/zkBXhtlX4F0aehtrVeQKrskoFsS
9ILSXXgPULR6M5GwgKiKtIM3avZzHpjQ25JPhrkBE7m2ZCCYk6LexZZ4EDA5Hn9N
aITTQWIGa/GyFEKZj8//LAT8f9YjxnHRCHSZVEBK+E+galizOyvonsI8cgnV/+BH
EtF9ksGtocAwP5n2to54cri9JQh03jWpvvqSLcKWTW1kzkcT/i7lOfbAmv1z+N6U
RBI4rBeWE0EjS8dRO1m3Wk3FuQBgByfwPFKKbU44bMfoReNfjX8RXc5kQQ04bLjJ
0B6rfaqyzRgXbrW7kdmmTcJIZW7S9EKlXuZDf8ndie9dsPWa7dbZNj0UR35GP3QW
kLgxzDQ6CcpDqzvkvPt50OJ1rJYtfkLlxkAsKRA/UD2ldT6i12h7ljiNhW2KdYOe
uGfIM3B+tEIGRRiT53cI/yW8TSu0zd+VGcP7tBkoCasPqt1d4EAOCunfINX+F2yB
3Kc60L6lev9v6VVRGyX3E2wqr1nNngyebJagebVostzIo6KUof9ZRihFWy7DgxCb
2QU4MDXzqOnkmvYyCulLK0cipdRR08lhawfvFEpQmJWueZITz7WImEzeuO+CVOqa
OkhwkT8JuI6fzWjlSiy5KmUxs/ui9UaqkXDD56s5g/dz8iyz7Q1GaPQPLrlV/KgB
azsFZFyn+p7nKle0PkIeqh/2xPQ3h9UURQX70JjwvJ4+LJvNd9gkHMarNaYot0FT
IZNA8BcQhbbk/5j0uUZje1vEI6kIe2mDztJ1Gng7ZAsaxAaa9kvM4A7wzOlHVzPD
yZpOn0FImL+9IsdeA8bfFO9p90inOVjKdrgo3SMVOShCaJm1RQSFWBw7Mybyy7e9
yL/c1NEyFXpzymnQZWutw61TzZ6f8xGbHRN1CjNpbrVZkH+1O6UlXVjKubEq4XF6
kGXlwj1qRdFLtjV6I9gLZ6UVoguHj9nv5jWHYER7PFgu/WWAGAXiMrvW3+lA4/cV
EbwQ1jl1TAJtTDvjBcJmAD7VYpnGPlGxZ0SzHidaQKTxyBBohTHbXujnLl8XUDXf
YY9GJOI8j3f8iHy43YXK2lVDFZXfDVLNh+hyeD2CIZgjaqZK86gtkm93Fi0tz14K
pWMPifYjWXpMoQEIw/U/hSvxrbKUHl7v7QuR8jcjdLJZib1ixqdOmRgfI/1a5CGQ
R+0SgUnd01ErSKXr3lpZ9sKRr5uIxsvsIeAlMoEExuea+To/07DO8dIg7c9LZ+vd
R9vSRkNJ2ofS0X68Jr/1LuxXb5KCm0Sd0nXez54ED3L7r1hPqhF2w0uL5nd2fWCl
Iyoe+wUxSbcDDJa5PEUJ4j6aBkz86n8CJVBpONymurHlpi47HHaV5oJItsNrp/1e
uJfG8knrgBFiW1q7vvonjAOOV/rEaiSq1d7dEIf4dl5T+NfWNzqLnfKSwMouk5gq
7C+A2syr8OUf6VVX3J3gb3nipRjMEzBqofaV6DQClv4hkZEvxKB7JhFOipDurZ1h
+xqnMufQr/T3TXJRdXTBeoyK+JtsNQ/EEBgBA2itY4DgjKri/6GnMatps7MU5Ooy
o0gIwovvQQkOJGeIkJeXqvgYCOQLQSqUKENLiWqya3yfTGNrHcewuUk/xxAgWP07
g/I1PRdEtAkb8MKytHvA0hBcGIVPizmGDVkluGnHEwQm4WB8ag9QmEu9U/EfXSmP
t0isi7rbrBqwOW+quZ0uTeyc0kmv7VKt4zs7lmJ5VtDSriVWPexzQGKnxB8BNc3/
dksSXe/3nzxFlslnvzujOkgIh+SO1f1RLxHpuU1IVD+Tkb4TPfUosnc1kbKzx9DV
GYDRBkTJzYwQXLCi3k8NK8pQSCgph+dAqYPg+L9ULSnzXHIwjesDbcdFVykY/olA
PARMbFjDQx0Z+7n/cg1635MBaIGwxUS6KEJDAzsaFF6virqe4tJ71+q4j6n+7r7s
mq5F1wLgkb+2otODPsyqA+4DSPs8Uel33FuhJn9UWtD3wwjigwujNVQ0uwquuf7y
o4oLKtRnTz42K5PAXIC++ZXt59wLPkkR0dxZQD1KC7OQhODvPVvncAZYhd3oUEGL
1SOlZDtRJj8uhecZ2/UxuWZ3rJ+vm4LyWU/A56nbt6S2rcTVvcAdfK8FRpLOE0AS
UUEq/LBWPBFD1lLM8GF1eLxS7FDWPK3f0b7cStdpAnGYUuYgDdaHoYe/JzVyw9xm
inv12qsLAkdnPQ09id3EsYrS2e1EXH2XC10HYKNq2jOrpLE2vB7vsR7YmWIuaKaO
5Isp+ZBaqNmYMIMuxdSFyNLxfjuvAJVRxRglFsAUzU9tBNWKtU3ThMKNpf96Gnfz
MykmC2dott32JQsXyV7gPlxqyUgTf7lqcUgRPq+4F3NswFu/I6fYgQWAZiV3LkCW
SHt5qToiNi1Z518jeW6G11sfMJU4AJgqxO3KmceYFNAbmBLgzNDxbpUda/utYnPd
lAiZC/bBarTjtSAA8rFfdbM3eFfqlYynymHCh2TOcHJ2tJ4cLrhan77vCe/v/fJa
iNUboLPLjFSeq2HOnuJFFLOEPuEZj6R6cQEpc1HGXGwr69oODWCdZbBhtV0OYFZC
Ymsj9McojDky8mWWBb3Mmvu1LWStmrbpfXKTvjMkcZzZYUKUE6T6CJNiakvqiuys
F1jEOhLXTY6+se4DwjsyecgjU35fvcranfdCpUTXanuf86yuNF4IZvMPr4+PBtF4
2XFTuTZtVgnGmMsPR5eA4PLt+hZndgE+wg3+pa0YWqId7natrfmKNNYaVDWX9dcV
Jsv/kQ37Wp4Uku15an2byf+CNp/QKefPhCdci0yQfPJ/Susyo+2VM2cqt7B2x0xL
JC1TCDpVi39ezqVkC2f1h6/M4nRy9UlNiEgO6J0hjHmhEXIcnId+Urew5JijmLkh
LQpmAVrxlnX/7tCpjcjm+aPp/n2PIZXRnm/wQxjYFhQeMve5ph1N9wN6QBRFG5xT
0cU/hFqU9dKY47ag7As08HN8U+gEO/SMdnQOKg/BCBzOwTF4GnzLlAEbFmILnGdL
NTfyLQfTeWepRiIyPLhbfeChOjxtmguvSsFPIS0WfwGOB13Rr0ULZGl7w9V+CKnP
MwfwXNgFJnmZ9Aj2jxzoVnahke/OR7yOJz1wmHDsv1Z7reuwaTjFzZYVSBKUvS4r
etKzjb099OwZ1t4FrECMTrS1f2zp39X7M3MsffctYc4Vo57PN6Qo+TustNEEXXGD
GR8KlNCKDIs8y1GneLMsP8WTnvghn86DswbwnIwXWj2KUuN/Xlf/7+LKWyxDpxCK
PMQ5V+9SLhIyGORjfMiVdOCI8Gv4qIAM1hH+W+wZZ/7aZ3/Lrmx0s9JQ2tRY9AXq
byNuwp3MyFmkVw1/Tl+/ersN9/lu0rWorXifBCkvfN0tYfyhQTbMdJgqtS+C+Y5O
QjBBYCyEWq941OibMUAAKGzP46bYe5jeuNnjVH+Gwa3O2ElNH3hgw24aAhWpRJFM
OZRLx1aFeRsg0L5vl7RXqz2DfThq9YPQHT7V9Ps9iMNtzthlKCxFD4/cH7OBIT1E
qM8V0QnPErIPRKtqgw3224E4Vhxz+F+KsCmDY8AfzApZNUrLzJoozwxPqd55GXgx
pMaD1efP1sCFxbmCaepbdxhBTr5TaNz9/L+5IBTtIJhIHnpuciYDmMslJboYLGep
JkWptNwZBmAFEaF4xqthEigdFSRKhkpUGKgpPh6HA2HlQB11ut7Wz/L5WKwPuFyM
YY15gqukZ74TDik+SCOufBMnkm9XarHhllWMalxBn6rKW1vkt4tYPYd49cxEc0i+
rAtvxiUu88lB5wiIQgnNCFtvDllRXPivKyPJLpPtr8k0jhffY+C91kNbnrpi8NqI
qP8QX2sOMVaeBEpUYsoe2tsvophddxqw99QFZ34jE9UQmNU1GfOOJq1GK9l5AsZp
EXdfCgTHzBS+BClh38Pz07j2NoKjHsLtR5WJhV5I3USAbtr9jw/bRHc18c1npxyq
Ltp6yQoMT+FpwJMvUNlTvKf0vn99H2x4A/Y7TVsh4vmiEfei/WQb1CBjnqxgwIEG
TktXoAY6TMC9V5CdRauq7o2zIGzN0inSEet6gVmMq++5pq46EYqS88zvLsYaSrSJ
gjWwRXvd6FxCxO95YZjGRRkjWrhQaKOSUuLZkvFAQiZJ+Uyhhc91Ixmh11VHnQnN
P4I/LOfLtDZ++LoEiYVLMCsFYeCspgc3oq/F2Sqzguz0WWzLUaByVZf4IN+e31P8
i4VBu1N9FNdUjAaZkcyuu3Wk9zgqjDCymxu1Llvq+50RH4HoI61k7ZgcGxBCWAB6
KH5q/5ozGqyNgUtNGZGrfvxJJWHi8hbhUUVCTyN7+fiemc5MQX1d7E1XNVisc67T
fY4yVQtpS75Ony2xS3r0dTQ0ssiRRoVSx2fIARFzcKdmh24CGMiPKw1/HlsVn/2q
uhnpD4DxkKWFaLW2L3LeA06fakwHuJWB18r4+2mulH3at/Du4BrWriEk424GwYDa
h3tyMm/JarwgclXzQcZCHJeMRCnnyslff+cjR9/9VfTAYeF5mXlPxldVmOdNIoqI
r6A4/FdUhDAFpC8mvGWPt4+X2ARrxpInR7Vq58h0+hMpED/SYsDV0rwfz9FUkwKK
jLXwR4MTFe/HQEpDeSrUKYw17DBTxrEPGmdx4M4pnG3lGJ3+zqZW4nMhiMuDwlYu
kwXYBOKxsjsbV5LlWykqLQA75HSwSPJ32+hZgtLuHngqIFL9OHj/VdsBrhXU3khs
m8FRSO4+cswDSByqOJ5nSVhKo5I/qcJGYL6PspFb7DpDx4F0L8dP+f9iRQvzrz4A
hBq1l/KrXjWmrpACMoYDCyjEW2wBiwlYyNufQ9QJ2EicqKEeBj0/FfsdQTLTG467
vpWNFFAObuODZlHz/JhyYTKa6Qdg81WZDYbL/D17aL/FbPfyEiu2kodMM/udYbyI
eBTW8gXLYEUHhTQlv/p8Q8bSqMdhFRK9e5WCNJFawtKeZ3p/kdViKT77Zs27gdlh
l5q2j7oAt4cCiFmN2F71+/syPkjUqCivvkSw1ciADw5/slEy0rvW9NcIMhQEJaj4
SzUZQGk0RwD/JR8FqCMowA65L/Tp36fOIPzo3SPXUlMeEHC+FoSsx2RYtGw+KnJj
zvweR3GhCdEN+seSVjCm0Dpo7DR1spSndVWOOUv9ZK0Yl0OcksfO6DzJKRtrjPDz
txXwVhQM/B0XJBmzdTZGEa6q398D3eA/em/0+tyjuJz3Ztj8n1dodk0P0slYDesA
5RH6u0iOwXMQAUCJ0yuSgwgtjvFPmQFPmfPQvlRHqKg9zzBomOq9llLWo/NSqEPN
Xdot55SjzS60GoiynunbANvwWRk4eyzZLrm+WZfeR6/yGfpDrKitAxoNML8m4CBW
b+yByYyU6pgJcqz0UsTadculx/0dB2Z1AiIU7COHRtaUoN4dUAorYVl/A/Gb22Wz
FkjuNNz6glm97i54OEaveS7DyLIOSbSiKZbVoRilkbQ6tCtkEJfG4vOTq6lF8QXd
AOMmTOeQbl1Q2h2MOgL3HgB4A3GKtxttkYxalI0itdkmx0k4sJGX9mmfhRBfyb4B
HDxLh/BWxQaQZDfQqLFJNnqg4bYZH+3GUwz+UbAvfPA8H4ouJL9Jjr7pEdYflEPu
6IfmCCc2uNNrThUcAkbkG7gJNyWchwqATRnprLvD+cD4EzVibmD5xyz+VYPzzfS5
Jjum5VX8tbC8hP++uPrWBoYeJ+QePvLJnmXl6bT/9nwYEhn4WbBUOcY5lr9RVczy
XlhsRq6C0Fq9PBLOaEgCKemcAQMn2AklUHVwOl22OhueeDwvMW5BWSmsJVu1pkUL
PbOb7LCgFYKk75oHniZZVMeMxJZ0v7hOsevs7D55TJLBfNYqq/khul1KRi746OO8
o1Scu4vNFxIcfi2cXtKiLdzktTtC7lqkjb8EFK6sYSNaiATmn+2FIdrLUjlLpApw
YjinzSPM2WukZZhOYIP4yMc9jhHgRPc2KN/JKdc9ldHw3N8HiJ+YuVoYaRTPggCn
DgLjNXDzVmTXR0MIXhWTtLWJnFGsU2QaWetIIsEwrWUnjAM4dQLrhyBcEjQHoydX
Onh33MMJZWHUJO28wChZrS+KEhSKtSHG1PzRy/d2AulPbFn5UP5b16iR7mccsdKd
vXj6hDPOto9MYWctmS8tdSr8pfrQl2g9tnKYsjbeAA7lxTwhgryEwGkY23nJ1ZFi
VW9C77QRi2zWC+SqBwKjQYZbjhxlY2Ezjpd3rxQhCqEsD5YZtb/hGqfYYkaxd2ID
SNHhassynnap2NY/IvfKLw/1TE6wTKJsFOfa4ghl8GU3jI0i6a2Wg1ANylUKxfZA
fu5OE1Hw/H1VFy8aILbH2OgGAeGl3p7tqh0wCna2uRCxRuqWA7rBmXdhEULJ86BX
nxC72S3y9IHpgWNgEX5QJVax5ikybQvTUyO6N42CfR0J2rhhMPfPo+a+6eKqPrS4
qmCv9B7dSW2yFH+O+8crENEQSkmMoteRD5UomY1ST6JUTEvPDE3wkoYB6Cf3PI5A
92+IFcllW14EcWBvaJb+H7vagh04UdXkgCFozqw2yPdQXPAWbYbTwwIKoJi3DsKE
ObgwuXrPnjIaoP+G+21ir17uRiCXal9TcfJc19rMy7zB5E3o7dwOJFYwdgVS946T
Zbdfer7HXk8U7z5EV4rXBGwxkAHnMCezq5b1pTDe8ZyGNijCMm2W9Q+6UdmXYO8t
TeQgPE5eNIvdBryeuUOfRrClK9lCPtgiciId9QBUBd92tyLBp1FNxu4MhiPXyvAd
qMmtKo1rh9RSstQ55ttiFtOmIoCCYfU1PVwpwP1WyD19+fZnLxktdBUmP+8VQaDW
jufrBYmIt0MpsWOrF/8oyiV4JRF/9Z0PYN6DwpyJDQN6J1UAq6ActB7lnd8lWKEv
wx8QpBHDy8TfgvaP+3Z6aSenZ4CjsRxZwGFFyBtIHBUeiU0qClKQ3BhuPnFaa3Oq
WYB2LhLBOKscS1GNNjhe6i7MQwp1kzkGMnVtjLF2iu7AGVEd7ECsnPbBz/Xv4bhP
pntEP6jo2ETanAOdJXKbPr7gJkLtu3vC6cA56cSdsV5pJdXwzfKrK7p5y4xk18FU
0GuHsI+s6iAmi10R5D4fD9S+MFkIVvvt54+869yP0Cfnes2XTwLst+Lfw+bPKwZr
vukCQj4lhhMvZ+Cyk1kwIDVxGD2GrPuoSR8gjN5euW0q2rI56uxyz3vZftAikKG9
afvbwsyGThaMgiLtgokw0ARKLThivmMWexpyK2MNi5JLpfafV7tQ9/J3Gjr8KpQb
vwQsBYaL4nHxKiJ5zT2lwF83I7Paqul4WD0xnIbykUct5E+NXjcsdIcOO+ftSBf4
KSZlX2XWxD2sxz97Xp4Oa5Pv7SKzG/qaZFHsddbmbVY4bkyW9NecdEvWLu5VK5/i
cF6ragGdP+v7KRZJUtgMrooPwqv4RdaY/d5gfx35BuyxTVv3/w6KU6EYzX5gbOME
8KxDjozd7dtYBbraoLWCmFfQHFF4Ukfk8lcbioGqV8O/NXD0VzmkAPrKprv5cre4
1UrUnSQJI6sMHPdhCeM9lVD99Gtb8E5o4B9ezuSWQ07/uqA1JXXXW4MHmEe2DfrN
nOtvPt+7n+W3Z1GXLjvF1FHWJ4XpjV/8HtUY8ZcADrytKnVle9IvzM5SR9HxabSK
tPrXyJpEFl5OL1EWfkVU6p5/iXGtKBQk0MisoN3bdCaH7g6oLCMjv9Fe1WgJVs+O
b80aq9EIK9iCe0QQGFvFZ7XLVLyxRO45V2gUAeIgUB2cItPZXkZDbR5ergxl2+E0
83DRSpjhQuA5neVqtSk6QGybc1kPJbE/GaiyucGrJf7NKjHJF8/Dn2PSjpLX2Nty
LYbox5tX3jacqCIYD9vqR3r0zdVPp1FYBZaZ1Vwg5c966gMTyQUQOoRWa3ar4RQd
64NkrlI03sObTpgLLe/6RNt2ET1EAgOgLhfe1wcP+RenFnWWskSCjL66DLZD6hf7
WVl+5Iuy7/1tVPUsIYAsygSH3r4KpN+RgAeUIxpZNjbLRlWdF2Lo8GYnuteB/b57
9hhA5Py+NiHQbXGmiCUCdxJJibws/pJl2Ydt5QHzA8TAj6CCtZ3LzOxfGfMVlfxM
MdsasxZmAy4Izz5/pzAyFBuEXcNaluHkRlvT++/GsRixv8O4xLp66uZ14p44oXd4
0nUjq17dxc4IffnAc7xzE9xMQjpbpQPk1ej5QgOlDk6QnYZjIIIf9y9yy0C+3EFh
6jhWEGdD9bi6JGCkssC+kuAFQBsjrlaJ0fUejFISNVX53/2Tl6eWV4mc2upzgSpp
cY+2iec6tNoZUqNBp4unHACrdt+o2ePlqjMj7DCmma1OyLykd+GQzAMQoBpsJCiB
YHJXUjlqvZSLzw6fQQ3VpC3CWX6Zizb4klhrCAg/C1iKGiapfF9rWOJWVGl6P3sT
a91FiLWjN1S5xYWg51ddeJ9UvPsIcHSzYk6QuMEykBULPtqMpsXFZXXXrhNwWI9f
AaUAzqPmbPhy6Jj+WCJ18knq5b2gSTQ0cfpTG4f7XTIdAaeci5UvW4n/kxUm4IUb
RFDUmbzX3U4QSaDuriB49ZKRZVxAtmcaXZpzmaFSB2TZiEnsOjjNkgQ0UOKsg73U
UrF30bf8ybuvg1sL8rl/lsDhNpKKNE1SqxMA7nIq2cnqrG3k5+GUEoPPcFhEGvWs
6IxlResT2gwJIYeNh5MAs6p5E/ZDlm3t1IXjgWwDnXxyZ1KjtSKDfqtVOj5K1A3s
nTmccjmxXT1iVu5SDS45tg8Nnk9AniFId8JmgWXFyIK7IJkt84ZQE1r/j/+Afbjb
O0BNPk3Mzu1S2oxF1CEm4kVaCXbgvKtzZP+qsVL6WGv1NN1PmnmFZROC9wQ3nNRs
BaxECdTTVEy0oJfbDHJnpmeoshPShTg3HVRk9W0F5pTReXYHbNJviqOaMTWu3pD4
iR47+xWTEDeSIBrHj88mM9ai+s26L3bQ5tyV95w26pbL16soJNVh8uZ/qxqoamKY
ihfE6kFVa7cZU06rb184pE1CEDkFQ/kDgmAix9fGhz9i1CmHYO8XtsgW5lNtETwk
aDO/5GsGY3o3t10qX3pkuEpDktGwuUs8knsAVWdRZDqgVakGTR044Q8By5CEy9sC
Iqe/WtFgEFyrKihgevMpLYFRAAr7jYXMZ9lHCVzfZrZF4Vdde8fTVAlQwmWMSMTy
eKnsLJ7lEbClnOCQgDrZLhVf9c4Wg8tmk0pQ4P6V425IJD+CVdK9P48iiiuuqGwR
m1YeTmn1Evxp5xVUJYcFmTqgoUMGkCKmc0cOmTBFPtyQu4U0VkZNTS4pZrNgMAoG
EsZUb8uAXz7nsrYmrVIuOqtH54+tzlQy8YYxFxvUdtxq0j/TjcCxm3qRlpSeIdyT
Fw+8g/xeY4OwOSP6Q6TxtXErBH6I7O729oTJBmzcWrQFBqLmVdiEOuSLGnql1Gf4
s97Se6odrQ6ZFQz4OfIFGF11+3bP2qV4YRi8bvoC7PqVYs4kyOwX6CvQJC7SFNw/
1GgC6dt2tqWUhe5ih/ob9+1M92XAc+EYGX0+ZBAFSVJWlwTs+hZmf4MGKfiKKNw8
HkySIrSYvjGaRIkp5WN0G6Wg3tQzaGQodtw5g1iXjGIt0WBJnjLkbh3A+hJ5S1YB
7xMXhMXDMOUoRzqBHoRBPN+o43tRE+gXIce+vrWXpB8PAVqWgKdbvoPFNqBZ/yUy
mlEnZoHDWvCLGWYaYIm2aaaDOvRvjjx8I+xjwA30y7KoQmvB1E7MolVavoQHfeH2
D+fIjcBWtGddV2z6doP616pnSMI3nul8m7ZCGtzSOzSy4uVeMa0M7f0NmW29pIS+
8QZti4Ksxqk5ATMPt0ICVG0amMeDqU0+4QfpfAN6ceNXTJhosFjbGXhuY/BKAkUX
5aRv022RSZeTGu5lKyDAheyFgTbdFs1YxdEzFjSj2p0PdBMxqNWLQEV0EdVotZgt
a3hRWBgAOTsQUnO7CoxEzR5a+GPL1Si9yEoHYjUPw8TZKeMpub0SZXe0rBsiQAmf
LXgcaA1C2WktEcBUJ5UjZoaQkjfITwJoxdQHNNnp+eF3NTkUeSuFkDenaUnQiQQK
jQ7aqFo9am0/MMkNfbs5AAq+fAwdKKIQIUIwD+rgDlYK/VUt1BzkigAXw3jagPXv
3eubQQZQdN4iXGvKaIaYBJMpgnxQBb97VLbkc+XUazhTldZgFs0bFYpoFrytdfih
E3cnPgQmiFwrIMKUp0BirTQum9IZLPdztId1/7UHIR8XoMHmlZiv2q6PEBaJaIyb
JJ232xyXWTW0fwVvvFogiSPfmO73/6o/IokD+6+e6m+DYWEpJ7btCjcWPTQW/aHv
ZN1QmmyFYwG8A4Xa4pR1Q2hwuT+W7I5wUNtIiC6e2SeB0ejjYcOYvnXuUOkCPJTp
suQAAt86/vxIRN766uowT9r9iAHbCQ+PHUAT2dIX4hatsiNLk6ZVN5sguQ5xiQok
9sg/JBYyFzCqA02PmJvdvdpKitE+ixD1QWu5axT5k6sD2H2QyMoEPpGczPBC3oG3
YgG4exr1Bz0Sr3DNoUETX0LnFK3aq7mB0VrKhsdH8aBN7oqjdFvqBmUDwsxQvIFP
T+VPfgAifRMJsuq8LH6+NNKieLPLe8sfNtOMlJQECtBQksPYLvkcjuueWr1ntVRH
QxxoKu2epYkDxsJqVRwngijFngt7fm6jILxIZ1gI7DlWmsqiBbwk5KvwratZez1G
c6NNB6L+z61s94cOXjIsCxigtHkuuitBda+2wqV0kVfDGgni1/TPWdWqXWtI0NAl
Ow22bQc0gQ1FPKYUD+Myg1tRF4DqmIOZqo3Sd2rNqeXXNPDyzYz7oCgnRBEgD/H7
S2mS5kn8Ir5Y+/dHlMKjlHcMUJVSQNk6aY27HiaUnYLjdcjdxho+4J0lulVoMFkw
d6k4B6NrCPg1Na0XCof2EeHIcQZEI6TjzReW/qFWI2GIF5yCHhlhRlJ8MI42eIEg
IjuKhMDvUgIRQ0NnwcA443Ju9bNUZAETNEuPXpAXyWweY5luXySMwa+Qe9+2+8zR
l8qT5aLZ0YlWmdnwH3E0jdsRPFRJR48eQ4zqyBXHeY23IjCVxWSCCHVeSAo/sYco
vPZfR2JlRhVoPFGDxEcyU1Ck+qWdhfsiS8KekRff5UN7mKapAovxhkuzkr/FP8o6
L/cQoXe3AzuxR9haOtUzz8zGiV+M3zDukEt3NaJxyqc/3W/lvJsDr8oGs/RrP3W1
dBNoq4zgu76u5wy3LhSU/dYPwmSD+527YofegafjqZM4HNKrvHOtYHTi9RrNEeIw
TQmOHHP5wZfoVNi0xGihDUqm9qqQGr+Dp7etqx/uumWDGMeneya44JCkWL8vrEVi
QsahRNXQNxow3CU+ccp0HNqjDj0tZmJcRMQydtEEUx6QB62ujvNcH2ut0lsZ5MpR
uVDgsIhcMPLSOArCKnJOXmhBLlPCd4p4+jXoJtXcgitTBIXKRB2/uEpC4jWDltDm
VWgwa/eW28Y7qi+ew8u+IBt8AQ69j4CycXRYFthzGhJd0o9ZR+8ann6vvpk03YOG
DlvQUp/vJ7I2CQJAaWZZ62FfowPqAQvlqWLXHl9S3zakpDht5JeUGiIaqD5j5W7v
Ct+F9rSOLFu2NAgACFQq+XiC7vhErosLStAWrG319o/+US1k+SRhBG3BMZ3QKKWX
6MsdEQfUEVY0v7mpfxcAc/a5XVYfur8JgScBNM2m1Stt9n5Jdz+VCOcGO0ixw0rf
oEcd7//WyMuikmymOWRSh11sIOfXNGiVHobuNS4sBzIlBytoIDfB2D2a4aqaLY4M
qe5aFg9oo4nRaApTpWP6P7a6ceNhB8lzR5mNxNkv0rP4o5kIu+Ehx4cfeb2hwKLt
1PrZv2IOrCuA4w1zhyFPOU47AaMS+G/X/1CXkCNXTC3D9dXWGoo4iy6cgxR5zZ+E
xGITNDhG0HByNaHRTgVEy4PwyE4BlTvanU8qoBi0XGo2ietEzzWBMK/XjMPgvQdk
rgIHZ7gHnG4gpZmhcLnyX1pOYfVciFQaowfCz2i0kVfW/m4yA1HeyMpwti1Tahu4
D1gOKuk7NJ425Kn1j4nOY+Q/etCIaRfDEXWe0cvT4oh1wckgD5txLbHDsoSu+Qma
tvO/lGZTIEeLBwmrZ5D72baBR7CFnCBGVxVbBccwQ5nAGfDymeFC+bijuxuo+LiG
N4sNZ3F3FpSrfBAJI6fJJ7FdjJhpawYW1r45tRY2m20dZLnN/Jybq1qry0y/2p/z
01lTQs3k6EvmILEhxGu0Xo4qW31Wjm4yEMTqWLwsJwhXbI7FBPIRGVLHKLaeF1XN
XLrao2LEYpxautcQMTzN7regEcOt9ITZYBlrmBm4AxqmR/M9cRchSpAPoLCno/Qs
PaMZMpfsk4MjG2mV1ojewRCptESTzWVtn3NfCLYd+6crWMofR0AhNT2zyKKpb1tN
RYDZ7OLlDtZa6WIXwUxsIQEdPsbPqBjfyhQl5lKjFvIyt3a2pJInBiWBv3c55qbS
E1Vvk8yK243o8ZyHoC63GKzaSycbnYyn/S5hmvbeXEH59U136nKO8TRLaKaSXVbf
Y+ZRoXEC4fYiqQcRJD94JWGpxfJmmbAFmdSH96B7VGMlY1fmRlCAtG9M/v6yAg1A
3jQIk8KtGLHYh1mcW/HpVIVIYXbMtXLUIlEj3xpmBEmjeYqAtsHTk1A9tMdeO8CE
xER1zVYB/uPLBzTgWZhldrFThkDbesj5FB886Qm4KoZkF8UFlTp4RW0BWMbCxRm5
OuLgUW/U9gkWJWuz3xFsTIaA+NCcp0/CRHVG0h5miT4bp4YJKJZZRwb6wQeq7T2H
DxOurfQxSdG02poMTwjI6oiM2NfaVooFFrViAcHi2xYdS4+tq7E9wMnfswaQgk5F
RhsfNs2ahuXVIPxkmafZb4X4JrSEmufhwFc+n3NVl6ZpaZj7tHD4zEnvLlClmhGI
YBDxvu3XAdAeFODjipKyC8LMS5PVTZBuYFdCVpG8I8lI3BYAH2JdYwqx1h7RoYZx
6o+tOE0EtdoKxg+briFFJYTzMTbHwwl+WZ3CEpTNhKjvHCOuWM6y1W0aXzkAR5BE
jT3dRw+2f4FBArXpogdvXJD/mCY5kNvrt9Dwk30CHCTO7t1X2F8M8v3JLRDLNLWR
k2pikMrPXCJ3JTIpgXslEQ2Ala4S97OhF/F3o0iky+MwJRXISaV1b/Hngq+MVPV6
YsqMp63+n1TAgoSn7EraMPkAIhFd0cwdCt0O3MexSyxk4YrNp2UpJqMwtTns4DgJ
sqIGhx9YE9MHG6ZupOwpWt+PoySWh1369V6vcPsWoYn3ayU0o4YgJFgGjphOMxGL
erfYDdHOSMcBKrKAm/B2peMrPrNqs0aUjHS2KRgXY9+8uYLovW3zu5MMqwdAA/VS
3/gNi5rRTb8E6zfYVGCN9D8vgp5XqSGm756Qfb0DR/Ury42J7ONlNFMS+zfMgIQt
YnajW2neTgqTeHU8ENLZJ+pKEm1oMN0kt3uqPeVUGNsxJhGyiCvX4jVSI0/L6G7/
dtv3Zw42ZvS02Rt0GO797Dt611ewt5OZN/yKyUUy2BdlTgfVFbbTZOkDNx5F8A+w
YnVgoQ1S+6RpOyJt1nJcaT4SOdP8buTll195NwH9I1MimAlGQw+EGV0g2vrHZj7Y
py/MdUJF8c6/es5DhIslxBxSTqIPFQVzCpQP0KWQZTCnmheBf8UpxsmHxqMoN/bk
o060wZSeM4uz/a69j2vEyiB45uht+DMhmTS5HUSYXZAdkDCAhcb0bSedTjIf6dPB
flbkVhCiLjG66v21pSDE+awcGjSrZxT0oDMEhO6YRf/sLrPcm9dVApoDzbh9RY0a
S0/xPQ7SrtQMEjfDxXX1LfT+QcBOBC/ZRy6GqYTuyP0wZX1DSrqdcGx/muCkDw+O
xy6elaBZV485sgUIJ2zC2BexqBto6ZIx5a54w4/fnkj1oZozMNY1h0SJmF44nQ3k
6+LqXk8ftpBaJEL+W+LoDp0oCPnRMPqa3okmeY2c7gbnjNub6s+Ds2VlOFy0ogXP
lf0yB4oT2W3Q/DTf5BKrbPkEBvQC80QZz1UOMjkvy4GNLdO7lSZCbyZR27xUCV2f
39eg+7TkXheRvUJuyNXAnLdB2PVBXjQYGQo7EdutzgfelhDuEgRRm1ANg0FY9XWt
T6DhhFk63pQjZSCPAnScdHwGnvU85Jbc9MgO8UPyy928B2zhUA2J6IzmUJPR9iR4
dTRwsYzioiPX0njOuNXFkGJOfZNw+Lrp7SiDpAB3Jq1dvd3CYBqNI8gSme3R+n/u
ckCrluFG9uLYCUYdiuVcgoRcbeUXgQrGO3HHf/PULvtM0M9DgnXKs2yhhLwbKdIk
F9FkwUgudONeic26YRmHwL/rWkNoow4OXVpuzVDZ6GoAKiykCfygpqblUH0g28rl
LwPwfBKbIagAfcr2BhxgxNN7A7ifII7Sg6fzvERX28YysFBbIv2mTo8B04wKY7dH
5P9tpHRvhBao4iYL8YUlr57Lie+QPPBe6JtL+cxarDXXB5xRijhcox+E4sEdAxNp
N/sVBaOdz9gGssg81o8n/jRe4UnjjwlMF8Sasg9WHgxJoeb723kDQ7pU/C2czf8N
Sj/+pwDFiWLWkdQkWkA7EFGS8dfxuEWqGTGtd4LOdMj8jCf7Bxh7w3WN3qkayjak
zQ6jGlRtxs785VacJZyp80eYSvvtEhxCAuSjNxZApzqbF+W3eu+UBltcErV3Kukk
sFVL75KdNpKrMjkAZJChkLrWVYwgOaC9ykl+xG+f2jGpM8veqB52quGx+qMjV9ZU
tiB1EKLJCcEj6I1Ji1ydblI0Jj/tJ+8O+C6XLaTuA/tJgCT9K3TfRzeoWr/910mB
QeV7PXYDezprn2STefRS+xTIJAYMpZ1b6blYswymR5wn3xDFtkAwORwJuzIp/HPP
snMVLYu/agWvFqUuQsB/GdwF50Q4ogfWRzHMcw3UCpf8aRJBESlrHcKfrDBRKp03
ET6KPFD+9d24MaifYgPIYV0h+FiaZrHrw/S4QXKhx6PMnvAOD5vPyExdE6PhPuMd
BrwT8v//sh8tGf6SSdGDCFvyIbN54hww/M0hTEsPc5mjMJSnpn4SKlEFWPnjRsDN
JYD+wS2neEZ1NN4wFenMoW7LIF5vfTI7zV7GrilmLfNCbjfphf7De0oy1XyTYSqW
8H9DRSiNht220WILEV8eQseI/X2RH7fEFqbSOVkMEYLQ5l2ubBzaQypPKkG4jgQy
XUZ7tWC3e2e4oFrlqr/vft8266ye+pbXeiTbl3e9VXHHr92f+KjTffqgVT3gryPM
2wmBTmcnf8KEgj8g+9f2MrW8h8IwdjC1trYdXPiq0ZOa7h+4k2mWbVHeFmezUpmz
jM78Ub7qxX1doqgBmwMsw+qaO4B5yx4Ou7nz5zlBMHke/Ji/K9uRZakV3CoNtVWF
2RtcybQD2kS8tvyFJHfjjRZ5jB6p6ZwOvqpYbIfzkpJI5E5kJbqsDLuntk3q8DuP
4cAkfI1yK7Bi4dTgpVfrMC0WEm4oxch5CppnLSCW9WvafNO2331RLaIWhT78yYun
GHn5zZqTW0OTIC7vrrR6+9JIUZBtLC8hgpQMhdsx65pqWP71KGZBN+DD7zb99lzZ
Aj6LCpySisOZb/xZSeqdo46T9YPB70JqWAf7oGj/enEj87yGJZt+vDSGS1eDXBgC
TyTQgHSS+rvxgJqgXR0JMZjZV0QIEBo2CeWOIo+baoJvY3LcHY+PwqHLjkkpQoaq
TCtBBl9q7g9OlqNiQByiuhc5ZKK2dooZHdE4Dyjuyas9CHMHAg2Hy5oyDFTPiIfX
lqLeMcTKnvXlWTxpK/oY7zAJA7dxp2Ty+REg0dmCsL0TxmfqPEDmY8BPgn09GJjs
YlZ9kvSebPvbdA6Vgc/j7N+rxlHPRw8W/a0yOBczChWCh6UEFgUxJDvRgHowxvKV
Uq4CDoNdB2UMq8D3STvb8GDBH2g/aAL3/7Stm0/LuN1iBqmiZM1J6LgtiXj8y+3W
oZ4uckTW1/i5WQd0lQoQV1pk399MFQOBAM2dSW+6l4jTOopT7C9YI5fOrRWCXDW9
5t3Uu7D0lSMivqxHLHO7OHCbPwZiAYpjAOHv5aHTStRZik9eRpCRRP0J1bEVyyVs
riIXA/Kip81Hd+gBwNvtMCFP5KwvMXvJQK24Zsfzfua7cL5IgTbdCVx65J33i0dE
Qp09b/B+1fn2Xrxilm0lG0ZowNIoy37kmWngL34NP0uX5MvpopnGKPxLu36Prj5G
xaeacm8LtLqQjWIig5dKWC3CJBv9LKmUNaz+WiwI7Gg7x+BCuo5aIlVPJwYR8lkb
Wd92p1/S9ILVT/5Ctsb1b6uili1hCQz7J1e4bXeqviVVcOysW+aEY1n/w+sTCUpH
tCOj+x8Y1N6V6RkT7xoA/tUNnUaoaIcC/WMCqMYbvYuxeODJ3QubxDgR6OeGVFz2
wgn+KpW9E4WxVhQNC5YQNlPrfuyhbV8HwRiq1RgBzz7RvvVvAbcPpZIsUhCseJ/O
5zGIFr02Uf4nFRHwtBPqyVgh/6v5AFPA3Lu4HEMKXxwsEyAyvj4sqxkHa1OGhOgU
OJtV/ArHE3/vg/U4/ziG1YFTLxkRWLDpEomgoCB+iQyDF7iTorChTrqa36NXbMMp
7V7i3gao7oeSDmwAs9pIj8K2fYI7XksopSvRo6/SIDBWhDaUSki4dzu5/IZS9r1V
Q7KfaeBBMz5R9SJLk/24uXmkneDxma53VucXV8mFkNms6g/MvI3pRy27QtFasOcx
cAhwo6sAxQSYsY8Dktb0WNfltUXyaMM/uDzmecl5yQqfjgew2H+d8fwn4ObGOmpx
XrkKl8N6cczNya09ueMb3yevih+wbjOKA8dX233ieM/OcaPpwtS7MUVvA5gU4iyI
m3pA0Afr5icdCnJNIuQIDb+MS0NjyW/vbsTmAlsy4iUtt3Y9E/jO85wjWW8ZdrRZ
q1KkXM5L3pd2t5fg56PnrPAZ5NOdHouInM1yQMKtZdx0/KFOn0vtdw3PsTOx6Z6+
xXHBJgj6StCOGSJ4Q6+YiJ9fX/+dvzNTuXckxW84hM3vup4cjrG8SRL2syky0LIG
aMXSPA3PGgRJoZfq34UJIvAyaaw9roo331KrR6qDFdkWqivB3maS53OAvGYvlYO4
2k31zDEZdf1FRCYRV7xmd/w9Ct+JJ3CX+b0XqKZMpjz6TObV49CflV1JmMQkfuvB
eacqWckc1AoH+J+FAlr8wcdIq27eWqCvF6IkhJmO7byVohOT7oplnfsNEbfzHapH
8pPG9SLICsRu4QccUxwUoU6v6ltX9KctMBHqVIYoQShyYMskO90dkJEsL82auZ52
rL0HCU7AtFlooT95bVHduh7KKjp+/Ndtdt7eZd47j4B0Exu+ZMIxcXzM3BpV3XSF
fR31J1kPw4amoUf/lVxlLz5rpRYNLTKbNcsEXhXJ76kzcu8kSrAP16rRRSCc1ydT
A/ffNbbITMi55VWHpIh2Ie2Z5werBesrLROSKzVIbH/rBtmf/UQ/+mysHCQd0ZgY
9r3wUA1JfJaR7ng/tgXqZcPdyddo1ExUfIpu7JbmKdwXABpfnjWvGbB1Fl0koQ7P
qW9so7d2ASGZFB0wNOM86ZKipteTlsy/H0hG6MmcZt2i+GUkKduZXjqYQ3GhfLAJ
mkFm708Fqr8qR8o39vRM+5fc4k0/CKV17SgNEeukDg/lr5BF5i2E57wbgA3tEUsy
QYHe8pVmvIIbLR0MYaCEC4YH5J9zmc4Tq0+qdgx10znLP2C5mURbtox62TZlZ0fX
25i7xJownCuc5eEVVJDr0DZqMsWE9elWPpeK9iURgsWJP7e3jfTa2V51OJSqekVo
mNPAiNTLmcIQZmbgokrKQF5B0xVtQ+xDurYMiQK1wcApRXSktGY8ARHoPPvaaCea
ScLNj1ie4aHhPjWyFUEsLzjwUjgRJq4RL122GKFgqUr65D0wzv6cht04AyJeObA6
SotrXMKkPNv4ghq3JhNphYoYE8oElGKZG12d41+/dlCNoco3sLjM1VpNSdWs5WWd
T2f5zw9Ekbfr6mjUJCh06ho5gV21taVWZ64+wQGWwEJ4msv5h3nWGnfL47Ieh2Gc
T6s8sBfm4H30EvqpnqrnYA5yiSKQemnciYuvNi5iCbJPsjPXEzpB6pW2CM9gvSsf
3yIv0qE7oR43J9MxiuKwdQOmv42YUqTWYW3yxXr7PUPxi2YefK3zP76jBigwg5qT
8oV21BC+iZ9HQFxAwELwVcgIBHb3jggft2R+hkWjRTjNhsIS6bnZ9DSqPAg7BGRZ
3mVUHXSDxl1GSJZALvbpwei2BNOf3zFDnkbCSnR1vvKSAa9ezsY4mGt9xlZQY2Tq
4ta64B50N7aCZ3q0HeEz3ACDjSdYPOoYCHoejxjpa3eGcKqjWdq2N3v/GZcNst31
I48oQo57EtekdZOJ6/VkqsC1qTP5kS3M5pvHhQzAf0U4F0MpTiDnSqdz2ytovOSJ
2AgpVn+o+WHNObI1Cv3aeNFqA+a/KgurIayA8ircQcGJL2k1VLk1frFzdc7QPMzi
Ftai8V254umGBteRvFlPzFW6onSTUJ3DAKm47K4g7axNGWjLDAT/w5ZjRk4uaohQ
YXYBTjt4GG6+IHu9z1xAZJBpyT6rDXS03RTuxh0ykkHpR5fwn0VLPM5AAnWUlJDk
HVClBRB2BsGbpwIkbrJqimh0b3LAv+GkYxTJ1jokaP7hke8thVlGBcHpEXCJtUHN
gOTDkvXScPS6MnFFa/QRm9wcs4i8Yc7oDvJgFkCmPR/H4XX5o6xg0JXwwJGYoJWO
wD8SuL86S/s4+CARrZ45sX/Cmp5l6xPJePpnP41WLWJ3zodCwanJSVHz4WbX5FWy
w+EgeXY5gCwWEezrrvMDyfa3kPZfOmVh4ZviYU2J6YXquVNeyLnsHf9dtu/hQJNH
Wi+1kVQKxEGE3T/ch/UxR8kNQ+PXRiG54Eiax6jwlbSqh5NB1q7Tsr6Wczo/ID26
QIE/m25M09f5gY3WeTzvxe9ZYfM9DdO6i4IbDE5boeDU6D+9CSCtBKlPSQs484m1
C1j1uvIZBYJ10gPCzXiIC1joM3o2OobGLUL+zZW8oM3tHI97TKj+KU5v7hWR8VZD
AwQtXaVj2nLSug1G2b8xLqj/epLGFa8hrCmJYG20iL8/6Ta7EXjaQKjbgtQPmzDX
UEJVBaM0f7TClfqIEzF4BPTIPm5KKGcLZWg+eWoxQ8a644bGrJiGTbCfh8EIoj7U
9AgaeGnw98T3KvVw4+ln76VMsqrBN58RG5bNxx9YDeSaS4u7wWipk/Pw0LiH+Vgp
fnaWQzsWUVpX9bxZ7HSIORfE7cEXR6oqKZvw+iYQSTHjgeyWD8ikZkaKz79DGwBz
BW4lK9SVQ/uHowP1/mpAZ/5ZfgNj9VhV4ToykRPX0NUc98+L+6YQ+b5UeKlj5Ps8
kmAtIgZzdEqobSOL900YUBY9oqbu2Zd9oPZF5MfirpKWU+ievZpPMaOiL/awGs70
KiA8bQVeAIomF5P9QDq4HxALV2ZENKG+inBuWQbvzRm2TFxlB2MyoHOdV/Ych/pP
cudqpY1Hhyh0LkJjRlr9NzTkmGnEEFnHUuY7vP8MKE3uRwAX0DvIYKkNH4Iqu3r4
cNSUWVojI72JoGxsRao/s70icnWTfEN5zP/JGYcV60Q98HiXUoXsWAzs+7TlDNkb
/m/eapXCStjCiD47vsJKJfE0jdA8gEYe7dLzvLYu+EueXdSRlShPAsr7Esn0G++v
d3KihFtvnBukATgbfBqsXdBqNLnrVSZVo+bewD2YgwhiQI3j/vxm5D0NXhOG4aO4
ISdQW/WphtwlqB2IeAwKVgs8SdfGc4K6LrQgz2gbv6xyYY86fe8owZGgylON96mq
8Ggb3v776QKsVGz7VXei6VCEqXRlBTWTj/CIdfYrOD1DOp3mF3Z8QOByMz/N0NL0
Aa41zrYbLSgLdilSDnF7850t6u7rWyPKJnUFEAwaqPY5s4kWA0Sjpk+Bl5WAcQ5d
iUNaisgl+BkWQpPLVnu9/bIhns3pij+WR880jkytG6VM4cTbv+tJLeMulBERfG33
HgqJK4bxW5hH9UHhuL5tW2SLvvfl2u84kj40KiIYpvNIs3Hx0f3NT/N85mbloBER
Fa2R0mh42emsAySnqyKqKeyxkbsRUiZVIhGA/hYMk+16seBCsmaX28IL+hicGn76
`protect end_protected