`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12160 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10OtvJixhnWeYVQCxik57Bc9HAiKtZnZVZhnryG0WnB1a
QgNpLcR/ZQGGrMAvYXsKKOHsi9AR/GICb8Z/dhWIiNMHcvJ+719H47GtgXvyzWG3
tBUKgjMpBK17h8eC5rmwv0TCMlby6B8J+NFaXgWaZrI8XfjQI7qEHud+TJBjpbuh
wkiikP/LBFIo8f6pcLV5wf/kQW4OmyiROvcwcXuCXp4MKlIMjnfjxkGayr8Y3TEF
2s1PlfR9iIKdxPq5aIdDLcE9b3T62UvDMYFFKaC57bWSIohF3ZB1GapcWq8TCTRG
iL8ivMHmQguRom/cAKEzIOQpc5b1/3fZJBfTauzLh4oKOJhlYBf/M/hY+/znEspH
gFVzs7Rid9r7dPVFa4+iPmKpChXzyBV537psUhice/frtUacNYrOJh6PQp+TdBU9
2XEmRpzamdSm+QRyJl/3Br/2aaE7CT5SD8YXfhKvLXJ+3wwJG19lTVImXuv2jqRb
13jdjSKNZvx5jC8nVsk7/bn9aJu5HVM0zW7U0LAc/BkebwJ3hhKpVAKybmcd66ky
rU3s852UnHKoS4QJecGtjNLkNRNetuiZR0iu1zu8E7BQYYmvR9nysDAUAkKZs1kJ
XfOT+eySCCJ8YEb3VpdYpWIobVmjDH4dWwHQzP8yn2MrBAiwIq/ZEz/J4VxWu7rG
4ELw3IkpCwZ/MtMv8YOLHefRvsO/0hv9Wk8l4571OHMaxWFmKE4M2cGhipPVPAZe
wtuV35TEyz3jgHkJekZj9yaqoegUm29gSHpyxS6euYITk43GB63lAPW3+2YPba+v
BO2b1yqs+7rzZ/UoK8rnc4kC4W1vahVb++atNTiPw3PApk1m+uoaqgk+y5IshqSX
MXce+oMS6J2tWtWKaKVunUcF1KRpmouhq4uQSvY4syXhNcAdsTTiz64osyfydmk+
KzQZLuRzSOb/ljrdRWUgD6/BFD+r9LeW+2OrTMHcvrNl/otWM0Aw8Wla2ba49vNR
vhXTjFhKG0m8KTmW9/2eMyKT9jajNtYxMMUn7/thdpsI/D+dJJvBbF+OZqe35gAK
KK8kx0lphhSCQXzDrJcsu/mXGDNLdTyJmV09Ek82XVT49uO/QMgxP94/D6oWWNWs
+cZ/uaAnUo8d0PF3FIi8BqSCQe2imxo6l+k2ZIuKVoaDSyTd2qiv7asJpjSAia/m
R9NJnZXhbxp6uyRYwXNHTvCBJhJgXVo/B+z5vomlA46KW6lKMr5wxVhsNfGZ4GKG
DZ2RCNR5l3XWUa3faJomnxmdMvvKpWIgze63h7g9s42E7e7eE2GXH9Ec3IEn0ZWR
Eb4zdoHn6Ny0cBm6weUyYhYNl1if3fCMh/d77GjrNT9SyG1xhkmd3xaU99YPsBCn
CgyghgWnyaUe8JHMImN+YM0HWMR+6iTCW4/1nMJNy6V+gFQ3sbLRaJTR+j4oebgy
/HU9F9JWzPhtGfmqUPsba74sWeWsx/u00FWlwWuhBBuFmpiex9VspNVNaZ8zPC3u
VAurByTs4zy34XQG/HPgJbNRaI+vjctAkA0tBOpsXFUpvC13lL2iIgALnD221IcM
53gmD4urIbRvGICa47KeJhodOEeAiO6Gn5IlerVCRk+I3xTDvGCvNhOW1Z4vN0tv
w73GBSSwjBKIuBkYgasaa9+1eEaH7ou4YCcIV2tZL2d0BPBg1m/Wmn2kH9domZk/
y3DLa5+RiTKebIvBPKh6Ny33okGz+xATBM7g0LVk9quy3iyt38WJv2GMi68x76az
/jCCXgOvBj4kH11SdYxX9UVTSwuzXLi+gsZZbgtFGmMH9TZ4R6CjsDZFphnN4yxs
t11RXy0qE1Zi+vAmb66OkVNGgWQVJAaqJgbvgtkYxLZVuUbp8ztqysKGPFHdD4uf
qu11ffpSTFzk6mTcWXvhr0+QiyW23oaACuyFzw2rcOEndJz2eElZHNKjqJTsZGS4
KnkMTlCxd3GGFGVmSoyifg8JK0JE0dXw03QQ52CppIgGkm07cdWtj0HNdDfPVscA
RIMIEUS43UkT9/w7jSMhiQM/0OljDq+ti4UV3r78v0mDzyAxEmN1S00JmrpX9+4Y
bJOQPm5vhSTZywpRl+zfC2gM7Wa/lT9x2qs7dsoRF6yMYQQ2qkB41lwOCyvnkYtS
nTIi/s9/fVa6wESKb9cFjn+00eL6z2Z/VqFXgSUgsQ82iAMhrBOYFBV5kWB8jeMI
FFrhmQXAqkK5FAEeEuknSATn0WVEa8myF8zSua68UnOoFIOOFqAKl2DrPeJPSVcE
qRH5ZTgr8VHjngtmurYuVcj2AJ5z5JCyVQb0MTzT+GrTjb1TnV48xgNQAb33LUTC
CYSg5LrN8z3BZaUPpYPHSUJ8b2z2yrga4DKH9Bl5g5cpAk0POZkt+7oSuTjlZegY
q7UoHGdKC698SZHO/8+H05XKZLAPhSWbexHJJKvD++yyP0nQijHH+ixxNfWMwL3P
ErQi4c5tl7AeHzrQjfNsws68R8sdDAv8o+KG4YVnTtQra/GOTUx92IxlE3X3XjC2
EBoluXQ3OXdadPAqeoZ7U11eRUwb/On08nh6aw3emZQF+nH09ixmKxf9XIfbCrRs
VCgvYA2fU+R/rAZNRAS8QW7/BCLjyGIR9J0U2pMdeXMUNzIFreF2yI+KtlTjqNIl
9yCv8ChpNKLfqGE+R5FNRmVjEeh0Vl9vkwvHaTqdU1ES9NRoe/S+yBp6ZGwyEZSf
gJ8iBaHS50QSwMFwI/BpirgRl9zyDBJAylqjnggVQODFS+cHgyfOx0GJ6jP85fAR
aAoX9a9Zepc+a/pUUPxoHSvwo2QSdiVS/hZ4az0czl3Qxjwi1jOCZydOIJKz1bCR
eukS6k2gKxM9AQucO5zBm+kngH75LRgB5jzRYFfiGzscJjyPhqDrMjPoH3ei+8l8
hogkCOQCL3vJb7QajVegtrOwpPG/JxHiR+R2B95AqKUJf9t8LKUZLtLGjTgKcHJ6
87IhdvGaIaY7r0CfGKNnJxdSkUG/5OO0TZ12Wyj4Uxkj2QlbtQm8c7B6ElzgkkHx
stbTIvQPrKv0rjaK+/jQbnmxCL9nkhv6MKgKhU3szgk4PrpwDDnCYd82Lni+nIjP
weF2XE+Eymdnq9l/Ir32hO0saRirreGlg5wpDWlCxZEVGWPjggT8L7DgEthSR7P3
6oj6IardmfNTj1X1CUyNV0oj7gDME/R4rzrJUGegPk7I7yxl2lmTO0Hsh+JsV41a
r9aCDdynTwHp0QsQcdjD2g8kJo8aFHxP7xSn+8bjtRg+yFllVNoEdsknHFz0EtJw
TGtd1VT8FrMXT5NETGTOunUu046H3vhpkAWtE8+D1YVth9WsGlDXOaxxeSgC0u2q
LXiFDyhNzS0UgkosdZ2FjDgywFKT0bDMOFqV6PIpMdwePRK3YkA1Kge+M5Qj2V7I
GwRzIikgyVjJV7Rq4Vg48RgErM+1E7kyntykvcfegbEY7KjZ9YfX8BbyG/UOSwJE
XX6vLheykg3N6h0u20pBSKKLmVa8TdVoxqt8uDJLPQk5eS/iaHBcqpgOkuGChoVq
rLa95yuO5clH22k4Er39UMpLcD/TZI9LiATiEewvruxdQYhSQU4ewDbVZsotwaH1
Ghvc3Rrx+UeMyOJcbn+sCpZd5ocKxJz/t4cyzT4kjlOuR/x1P70xx3AdZaYXpLYy
BrLM7kuoX14XP25wQSgeyjEjDAh5iBXwNYK0u5M7uPSiUSz5D3+CCcCZ0RT5dPMD
OjLDr6HhCaxD+8eLKpzQdyf7tLCu5EDiVrPnMZ4kEkA8xZv6ZVq9SqgiIZby7t9h
/xyzX2NM7JZXcTvrZLdM2pB5OcIG18deh+E8Ad09wmuP5VHwXumEe4mkQWiNfZPY
A0NUtk/0dCaOcqNwXLQF7MDTmAg5/lWIQsxmGcae7iFMFxThkmdNl6uh3XgI6e5n
SNM/rLwYIjSj00g821abRYFZOPyukQHp+iQ19surcwCDblI70XlAAsQV6elpbUTU
JdSI7AW8EgxvEZMLMA0L+RcIDL0TwErss5Agzv5eox5BAV4y8nMKja/NFYGMOwiJ
TouYgakKGjA2NrvSt1uZI7De13A4mhxB6d4YR6o+Pln9VlAT7V/XZHTBL8defDWh
KpjIuguBmHe4CeFAgAb3oxy4oDkN6ZWa8VeRAD8GcaD34jH9fc98KwqNlAIaijq6
NLwp78LmC4duUcALYRxqTNCH5lcnRacciRwY9V+xlR0X+Dlo0ToH3lLxDVkzv47V
0dJM3J2JTe4xLzALsypHoVlHBntbEtJ4wgfQ+ST4Rkh4/x7lrQrtFIWq6btBXYa0
0+EnTGUMwuCEn2b3nzYd930PvHOgEM74Nj+m7NMjTKu5i+rWoYQFoC96YP0LD9YO
ae+Yv41U5WKyiM694JIRo9P2pO1r6H69YsAXW/DMVnyC4wTAL8xr2GNFfzFw8WVQ
ad1lfi8cgLx4qn9bo41/nBbknKcf6mHD46iuhb4/gn02CTCsKHpMe6rnJnc5PpiX
PY+c5RJz8vT/xU+qAhbh2dlRfUJRaxOK8VjEGYu71qs6JmuxVUH5C5PKQdfbXwQn
hStndxkzBEGcE9jQvbwVjLFT+zmvskWAjdJvdAinyG5gtMndk237zQk3kvQOcZNe
+L8EzOQsxObB15l6sxkVF481jyEjRdBOfnf81Ye3wwV1vuBU8u8Po7dKcA0m2cKv
/+G9JWUaaPNYmtbJZPnDpHgUsy2JTFATXpfbuxhnnzx+bgd0V8UkCNb7lo8iitSu
pU0CjPvS1wJFZgs95bq2CB7AwhQwRyzbtS1lU5MF6d7KjtCUNWJjDB9jJ3uTO4Iy
X4jxhhXXeO30CL1s1UxLe4nlHqRJosNeiLpnnLCW+u587LM/w0+o8i+upYO6htEo
PeUHWFa+bfjL5usc/qiw724ulalLJ/fd6lrV8MlCEms+BkXC0BM6+AlvsE8MH8GR
260RFINzPfOXE2wrrwti3pLRk1m88aRHtASa2OK/sUNKYQGKifff07kISrhxMhLA
R6FqB2WZWtprhYqg3DE4P1j+Cl6I4dFcAzCdARaXvYVI+31j1I/+N5PkOf76jTK5
ztRKsXqn+cXLmUIw75rLeglVT01tii4JY/KA7vvf8jfm6eZ22+AqpqMENeAwCbay
HW9Bx5rK5IfNh6945kzkGz+fTS8Po/TPKuq2QyECNURVPd1UleZg6pmH0ut/ZVkV
yFx3MrTkj+k7zBX05EU1X/HZ1dm8Nvp7iMzzAiPryWCq9XQkDpt1om8IMJzn8Wzy
YL0pv+zvYKvCqsLakQtWX9/EaN/WoR4/9JaN5XZVx+WvVCPuAWwYI/idlhvd70A2
QJnJwuKYI20kFVTg5IaokKTPBjkHPg1NeSYNZJ5cGcEBOzg9U4yyUsWriiOve5pe
c060xBYyKptErthNc0Fxneh3PlpeQtRdR2OtLS27J/f+grUcbYbBJVBLcs0MtR1Y
8C7UzJI3pX1umLRq2ciqPMq8oyjRCzfLVLaSeh89UyljYcOU+aonTlf4PGoDtEnp
wQAp+2kJd9dj4TgqORHjrd4NJBmUMdK/mIP4gVND5rIyHwCkZgRz6c0mmDiYl0lC
Hx9MigBRnY9RqZfjvOXZ/Sx914J1Ulqioqk95Usi2MIu6geLXJIXq+3kldhFi3lp
RuhJw3YIr+AQiqd5+jiZSo0v+3xGCvLsP18aFduoK3kd4UQ/1zIRNSjdeAu5AKb/
uRPcseg4UK+RKtOsV0iTDTqiepKFC1s3+8mSFobp9hv/WcKLHjYS+5L8HXjAq2mY
DAeM1h+zMfSbcJ3BUkWRHmnAUz7pMdPjSG4PiTGqt1XLVbedQdwZA4PWMLv3L6cJ
5f+kpQjRWRe/eNKso3cW+mFb8ju9oqk4ESNMqZmzVNbxAHmD9nMkacUrzqlk+TpA
wxY154e+GLpeJU9sXJ/EH8tue4QpLeEo9s4Z5Jj85Bd3LNuu1oXLHk23fcmV+bf3
mQ4gcUD0a+qDe3dc3kHBjPGkcz843Aeykm8pKIqFrrCn8z8gl77POFqsQ+M48RUx
/15C2lJDyyrvL4JnSU8pLY5Pw3SsOm06OosrjBVvbPL+2OSNhgW+cCL/Z2V0g2Ys
bxR+VUjae/Rzec1Ibvn727ukSBqVZc5HWBomwEpMap2DWcJwgtRDKGUG1YqrYD4p
JTuM2YW1SBayi85KoPxVGYmBux53CfD/xJhZ44aymkKlEnldo80wll8G5DA6ZKEz
iqI+a7o2eyqEKZCYzYbkT5Jca8mP9yjJcvTGGrX/hgUoKJ+zuMmhY0ZTu+84L3j2
7fIuB15WQpkmj0/WWyQaneVBJQnsQ2BBgqT+s8VE5ikPL5Y9WxN0dsexFoaFvuzt
Np5cAJcPJVN8AMUW9KtuRL2yjm3g/u1IFHSdTTWsa/zNR5+D0tIdxLjnYgQYPMXL
N9NXZXMeGYRx6xNmfWqNRa9SoAKgeSI965hoPHZAqo72c58O8OAP0Dp4fmlkbm7M
9GNglAG+2WQET2iFtLNeCXrqU2T9XY5VfAybyL7kftx91AnJ4YF9gYBsU4hOHMPr
FRG/zvQETLKapomGGzEx1N/p+ecPJbWFfJOo4uJZKQjl3TnA9MQ/Uyv0vQVvVxQ8
QZIKKK1baWDTK/DGuRJcFRXMvkuII0oYIEx552iaCbtbSgO0DPgR2t6jzYU8eb88
IpF3EU0uq1Qjk6FdizcLQ6k+71bv9g27VJioaQfwxxJzD3+2UPgZM8VJmi4siPGS
a/OQLKe9CCQL0pgrNUm0SIsHe08e1xVuBGZu0vC5aLMb3i6G7vr7Rgb4J7AHzHzW
gjshXjudctT3C+Am8yMQh5mOsurvqBeEULEqQ8SeiOQhrHj+WjT+p5vmlTh4PsUz
yl1wUYleqU1aFxNvNeOku2wVw6bqFETprWCUNjebpb7vG6vU63yPWSeIPr0ZFZ2S
zNw6LeX81pAF5v7P7eGboiG4G/hCDD0LFMQbFNIfTQoMnSLice2NE7ISrLqOtMv2
jn4upTLm/aigTRusUBzilrH6a9TFtkkBTWzHLukuPv6u443PnkuMwpf9g3XSA8/B
3pNrQ7iaya7l/MXQsfOQLmdWuR6kJisIz3/IQuJo/Xu49KpXa46jvtoutakV8rAQ
9vznPeGz1qq4ochMmB45dQib9i3jwgPT/Gk7fkwB5OxzDer0QzjCXXdICfahR4pm
kpORN/f74LuwnLr7O2ZkXanN4QAXC+6JO7T+Ns5+PQV8kcaXapSr4gEVOy3ly/JB
GSihhlTBotAG2dMacritHyDFqA1DGeOKeReGoVncVoZiqnYNcWgdUHzhb/9amntw
T5DXIKIB1ybKEsxskNeiH8pYuegaUT9NMj71DqDHCJpm9FLb9tAFHH4NyA9DgNi/
0E6vrFa7FmM1SxE6Dllb9yOhrtBm9iFoAf6gWSR5tO6yW5wZ73aeChOPy4kBfex9
rtS2pIjzRC60XJaS1KIDz9hdhEuHMyLP8Welqhh1i9lc9CkoEpvRAVcVTR6XVMwn
nubZy6J19jtfENJgCVazIAgACkFjtj5OXgP2c/B0chB/uxlUdrUpF7FbMcHDpaZX
xNtSL9uY8c2Mc7dTiB3DzfK5Sx0/FYMMDckUZqm9Vf+pBWuX+1IGi7wXZZwqwmS8
4zp6t6n73xzJy4wjahGHdr/0EG712UNG6Khl/Y++LNq0CzSuJMFioDAcTzJLwfWP
fVF6nX78l/s6jbNqldfYUbZb4k7Hwm9+3ZybMghYlVD9gkWmtrw4Zqwpng6yOFil
TDwyfWwy9RrXpiDXb4RTT3E3BRVEFJzbHhPzYJnMUNcJbKWDvA7ccrzQw5DwfhUL
rCWKwMMpXeBDKmHgwHHZ5opdtqxforL0KnORK9qfMqzGJwns+qQF90/SAcUWM7GZ
NqV0H1fBiu/DBfG90B0s/kklKDs5mXWNSFc1T+S/lVshcS1j7WNm4Q8XKl4w+rf7
4ya3JOT2fT2i/iNF7o/FAdyt7llcv3rwDOxz5UfnHB0NMEAQ3C4oO/9Phkl4z3Yn
LSinVRU8IFf5AQY9HVxVtjbdBpDSU9RyrKQuTJH/nGRxXu/fzUyU+LoIAbkPUb0P
NiP4hXRlP50zrRvqtUHjoZx7VdM2lgq5+VSHsTIB/AsjvlyDuk7GgSv4xznvx1mo
FLlh6YlixEKHtj00qiR82NXxssy2L6yUqN65NzS7yEOgo7cFILUxGr5+WHhSkh0C
O1tlo7MRdBZlu6S/TgQmIYY4droX0A3Zu+obZuhTEE5xfFn8P5r+blFms5BzqGUO
T8W23oYyuQCMKc2fL3S5FKQgfLM9KJY82348UC6+LJxZeaKIlP7hT3yhS7lpUVjP
8dFTSadcI2UWEmBsHo3aRnadN6o3e47SNSfQPXWdlAAlaH9z7iC/sJP+ast4IiNb
BXtw2/vsizxhcitekvwUu/g51Vf6qssx1XjHPdLjUQO5pLuLJITYuT+L7QzGvnUB
pvRsAg4quEt3t9KEKsFuU1pJRumN+V4M3nmpE60KdPHUZ46/JjKh5oXGud6rxPUS
7JAKdm6s7Bi1E97mpZNN52/bel1s3cuMnJWtYewcaS73m23HoZc0J03JeIzp2vEB
ce/Wp8/NyI/nKVAgJsFheJHTAkqtroIrbdq2Ztzly78xtisBPNbsFsIdO3uwq6/a
gsHGVvD3ITC7j01zSejM6wKhpFFSjqfYTaFWH938usr9a+i09Gss2xYzjNeqAv/c
+HC69vzIN0N5O6HMv8jGHoh1qSKYa2WFiNPZhrwKV0maM18wyGUHsXxzKatGXojX
7sm2cUjhWlK1lHg9O/t+nTogNm5y6Q6i5OEiBz5k/TyPcCR9PD2UzIey+OE20yyY
FXv343UzCoZ76Ktz6Sgew9Ir2h9BeydjNYdaR3YjbBzVgAha9reCk0QnC/j8jiJN
ixlrhXAE+BBC48T7Fx7VOx9v/3oZOxnTgSo6lZmokvOaEo7naN+ZLhPUlu8rbeuQ
aCiCRo9GhDjeZA0cKylLgVzd9MlDKy0Q/N+CBRqVbzgQJJJUBTpChVG5XIjOSBHY
WZYCjTbpHjB0Pz+SKsa6NP7CQm/HhZbQrtwYh2TjVgQ2hZ29rf0dhvA3TgbTsHyS
tWJCKtfy2fQ1kMW6vgtpqA98//sly3B8cfi8zKx++3uvdvpaZfArRP7MKEnwk/x3
wtqpvxYI6312QZiXNPj+jpYhZ0JuxlK/u16QTpgg0YOAovkHfGiXXBcAvOVsMeJs
UsDsJ8MMpBTuYvx/NS0lqWCWxAXteLuoVvTCOBqfEU0qV2ulX4UERcLqc2Rna2O+
+aPPYZnnaAKoTEW0VG3nSrLs3ZB22j1GbHX1TbcFpFE2KOcl3KVWvpIVWcdKgp3g
ImHweBTwZLumj14nmFMsSrJERTUqV818IiJJDlp9bND01M5FQC0kL8xlcrfOURR0
idlaF7GM8MEmAwCRTL41BpcU8pCOpUjx5gUNfz9T3cW6o04GFv1nHoYy366ULf4n
nZeP0iDZErGP+UqLGM9miPuSZlUwa2xBgIt1bBfDzMC7Rvbe5rI3HEZG0RDASOQU
OegQPJrG6bzUvnD1/dm0zplrTJ7Ocx3v1G/jK0VbsbuqRDT2a2udL320HuMiChYv
iHnPsDghqt8jMrurvvf95Xsqo+tMd+6EPlGN+5JiDnLZa4sb6xd9j8+976pBSEI+
6wVaMzKKVvYeBBSHfCH8LbbR0z3agStb9UTPlqa4jCrEGFUluBVoN7UVb77U7bCl
tloC0FuekB9liBkRUz6qIwHX6yo1Fumjn5L1re6BAQ5aIpUgI7bzZZ3nbCYGcFo6
IHysFPhd4a0dHR6TTTbl98szCgFUprAli80GyksYl3hcVn7djo2JG406FyzhRD+Y
/p41vXiMtz4RDe8lKkqTYkRfnlSlDVMX18IXPqMmrgJowjm8Yjpr5yz9pOtGIhYR
Qzcb+8QhGCp6k+gnaIvr/mjRcuO/2xe3hvT3pjYQB/rKiOzw4TrgS5fdwqtwhMYn
P9XAAp84g1a5Q0ffbYT41P5/63+1x6PsuAYNCCLKINjyxAcowihy27sbemwtA3LC
6X8J3fgh/EhuWYJer6EKsxZPpzYnneii/Anir6+rEqWj5Nf3d4Bvv6hMQZP4n6Ff
n+Go3h4taKiFldVUFXPiIifLSaFaFL/FS69uQRf5cqlpK59lQXfPkEFS8LO5xdM4
QxKBMJHNF8tEfJARAGH6e+mvlZG5NFrVLlPlHDgt/XKbjo8M/iag68s/HC2lXums
c8Fi70afPrh7G+UxlrOmZNpNvX6DxYbzdCRnbZ4Gln+NvGojldEQ1PnAcLXsVv/C
UQBUwPBX+p5KYbnkd5Z+wPA52tSN/wp8vXKpSTqNPMC6it3nY7vHZrJj++OS/DjI
6tkxoL8d9CDbre0VaKJ5wy8gkGf9R1MeFunBDt7LwsG+rGhoQCy94AjfcGgBDp0d
Fkn2l5yJV37kGfHWkDcXh7EEmWrlQSrGdUlWuvz6uvPhw1rZjWXfjx3I8AOybtdA
9oZUx3xjXfKEK/MhotjmBHc/saRvi0Is0LwqNL0v8Xr9O0KV/lu2TpuAKBalqtRf
R/zGqr6FRS5OuyWQe4RdMESaRjY7DNwygu4sLmQP9qsLJQpYB4y+qPDzzA+CY0o8
95lhkSGcxetKvz/frah0za4x9/2S2Dns3L3IfHnmZ5LIrS1VhPR0vdgtgeocfXHn
7/Achzy95p0kCkbxMg8IM6bW1Z9quZp/KZ86OvFLtTmqndG2HfmPo9DzdfgA9PqO
OGR+z+7rbP6TWQ7izSbXFC3/Xsc4mtPhu8wo78a+O3BHtac6ZmHOydPVoxMXP52W
D7LHudo+HcBcy72zZCR/413eRR3t6D59ig7bHX72TtBz0DuVw1YpXDKJp9Gm9Xj1
PB4Dfp2qZoBl9pB9F5VyKoE0KYsyqFYrAwjY0PXq7fgrB8ux/7xPHxPD8xLhVQgy
JzPtCNdUoxyUO2JcuJQGMMUCLcDZ5QxlvkBbp/EkVuIi9EWSSbz593NIh7FgL0iU
+QQVNbWDtz5bLyKFGLB42cxKzo85slc6gpxwtuRKJM0KhgOlaUZ0t26exsmMTWj9
E+uInO9GZ12fJV61LHtv6tp8U77ZHVbrQ12GXjThcnN8r1kdGKCU9uUCVRWwO8bR
oInUBCYa5VJMsH4zHCQzpOjPqYFNvfvbYAkXyaOl/cDO+Y0aTVcVNdxrHvL6VGOo
QGfAn5e3vIfQZjJ4mH5kWsqyW/c5vc6bsoAk9DQ/02ANRD8J0A96Qgq4M3xVqhnB
oXqrZV43GjRMUxO92su7c2VSqyE+g2v5+JS3cNkcu+2dUIca+YCBYUEXbJ/GGMrC
nIeNL01UhRrSizvR+cGWfrOxuoiB//hOWl+eX2cfE0pw6NawutKvpRr2nIy1Zm2R
biGfO4BKa2x+7FqzQeP+yOusJKDcCDrZWwM6J/rU4Ovv3qQVDnYpNGpfJ3Qesgj2
d2GBamnWmzFn0FH6eohDUO5pwPt9pSOpPbPHxzfo876kNwt1AVgCavze61T8lRhB
tmVP7+Ile05hOLnwhslVPKHw27jzjTl87p2hMSVQfU6HnRW7/ASGBE5VQvQpt6Iz
DqqXS0gIqxgF6WbVivUdS+GTZ+QsKkALiblnri1r84K9PVkhoEF3oQ0y87e6LeKe
RXir8iQhPqDLr2wZtkfU3C1mss0ut8AFdHPEkJzixNPTtl+086TIOU8NORO2jnTM
P8i8diqOnJlRXO4Mk1L+WrAjp+Lnqw9iQBwUJTx3O3jVVcdloXMlRHm0VZTCyEmi
EmRCSmAtU7cE27p6pTp5hxEuP9r21OmqXUhsihQCWXO7tTswNXIvztilztGw23Y+
StNxJZ8TYXbiPn7qSP47MHz+R1n1rJ+kajUpo/Wbdkg7COEH1dR3PmM4u09JRkpT
q4IQndL8w9Zu6teZFzGKeuJZQHYC1s2OjftGKqhpu3YQeL1oygj2qVuHGSyCwjCN
Nz59eOnuSPt7CzOhMTPB0GdXQHfGuqvtMRTJlSbiS0kk+ZFhIBK4oi1CoM0B2fO7
/LjgR43Gdz9Sds1g1E8idamZQ5N8lFDgROgzY7NwzWse61Z+oOCQSe0RIGZZCvI0
lszMGF5NEbBaom8wrHDUKvByZOxHa4Qm8LuyJCHPMkkJKfRWxLLFmiJvbLNCm6ki
/e2rAQquV8NOlgPLjsNgmRuMejnZBYZp4WQSeDG1GOaCkzc/L/U4LoGucRqk3gZk
NCecxPmw3eNJqRi6hxY+L6srA0KigzPYWhxFZmvIr/wJ6heDeb+5fV93ZI5ehmEg
Xx04gWADrOc87EeBpDxKV3fJW2SvC6hW1w6qIdaUgud8zCLQKIdIME9ILsb8FQcV
seNvbhV7RThheMRdgPaNm52prY/89KcA9unA0wgxquIvPuJ+FCQ7dp2pCf3pZUsN
D0yz8YeUl5oxhbHaQZuBiImzxdXljd9DJQqU57WWLlxqj0pbn3S4mVjeyjPhDh9Q
FrWWZwMZhSnjZHWC+OFsK/I2zDXJxp6S+1/XmC7uCHFXGY5oBUThpOGJKn+8YCFq
3vIH8TcBD40r21B//q+A9jQZvdpmTKSSbqyZU7a+CUShrvDeyd+a7FzdVEaP2ra1
KiSzSu7f6lUCr6fEEoTI+hmSsaiLYA6JxfC8w0OFOyw5dLUWO0Bj/wx3DsCzEE8Y
6Bw3fd1ivh5qvexAbIaSXwQKHXnAEeHWpI8Z/oFkAE4cNK4OTMY+4ucNfutp1ob7
pO0k2DHALkxzgZkLJ/U6UC21CD6tb4c75zBokaXt+ThhaShxA9P6xj1TSnfWtHed
iMuyVfC0bv3bagNpvnxgbZCu7SZod2LGhRLsAK/kSL2yrzoe3gEe0Nno6mPifKOP
1JQiAWpRfBBMM3rQc2qqO+pKJFUMDka3MkkNGhp/4DP2Ez24Y7LKFo8S6IM9eXQG
85hl/tV4cRQElcc5KQlBHwuFHHLsOq5rj12aznVGUgv/1YgWDWEo9b0x+l6+Ub0h
+VeR+f/dWO+c4HPVZr+z7O3vRra/q1THzsARLXbBapT5BWa+x5pVb12gsuyXdZbb
qIHFR4Clpn3Tl/LUiuQdhQCjVFeGBq8CAREHPS8XQ3UiWJUbokoCLjG6YXkMTtRa
6+y+9NDUFt6H3AO/0yi4N+lzJMgbh/z8wGX25n4F7dqrrGayjz3uttNkoQd+VYvH
75dHoadK4iyB+EydMD4lul5e9yrvFAntGx/KWVeFIyx/U9uFsfOrXVG1ZQc8YcAT
0AXwk5+yOa5i5o2ELq1ai+HXH+8nFcAeyGTG2C6rCxbNprz5BQg66NLuLqM2NHTE
C0qiymlj15tyafdwElfF0aYVE6Nctg4Re15g2o1xUXBYofvnfuaEH18DqyahMbzw
xlCyBFWK1IsDYEyKMtknbYppHdnaZiMyFbnsfMux2wmg1dIDjO9gmCn2E3Llnlyk
uiYsJYBFe1cmkbwcPOlGc2vTmI2d9PXbI2i5Zo4VBZv98GvOJwJ24zAshcHWy2Ti
o49L4Vfr8yjGhaWYn/ziCbHwP+NFUhHFMCGvpBxlPD0jx1z4J6LsjSZWX3NaoE+z
izFcxdcGtZBjTw9l2QNjZyaj2lADaDwwH+sm/kkxCfipfhR8z2U3qSHV3i5IHbxw
V32jn6mz0nln+96Lyyq4UKS6GYb4KahSh7Ys4BxWxj5nJfmRXezktTeLp+ITZYeA
ebLKr62LVhqtW4qJpYZzmuPqEOD/yxo1QveI5j7H9xrDJsyEraVtB6xxVhJ/fr74
EebmTy1tWank6tNhZe+Cps3PNuRHiG8dN/F7BC6qBcVPOpl2r9CAXtZpnxxQE9Uf
BrcinyTjajdObMVHbV0yTT1+koc11DYHk0gVJeqFeF0+tl6q7AJY0SEWFAmQ3RD9
sf2MyYg2QQokTiAq6gGjH943jB4FWwqrqa1BYALpsCnuZr2Cr9DDLPR0hJ9P1dKM
AqsqhHsaWp10ShIMTDqLgsZEgoJ/LNixe/38MwE2mebxn7VtuaXJaNS63KcTE5wb
IJJRCdmj31cH+82vjBTIThmBlXY+/Xj69b8ZUSG8QHWcwCD9m8ZxHCpoYcVxU+mL
LeoLdWhdv13O0lqnZAROJPUhE+FNvn83b24mlswTDErrjvllSwqAW8+X6pihrrPr
CfalxC6aGxplinkqbdIeU7pAYRvEzvCLmah643S+j6OyUbDgO2wcKnIfXUGA05gp
zrjlribYb1ePx+fK3S+o4zsfEWaod4SpXW4BxQP3t0BGQ9AksqaZUj+Pe/trjgqu
z7e3lfup2QJIK0EU1hATsLHUb8PqOVYTUuHlx/YGLmGVZL3qA7dnvCAZhJ1UWSUz
14Hh6v8C+h8XjSn+t7xarwyk8rQpC1eFUSVQhPJw3fpLR6/1604EPygP7ssipvOs
aE9PgKt4AeW08780Mncdz3J7HiIEsr5Z9ozF5n0duAExfS9k8n8J+ENLc12PoaE1
YnnQT3Qj+2kb4NVnAZE3X9AKqWuqfcOgTrPfR3aQT+sSAXgGYOMOeO83sC0UBVfZ
C1frrTBZe3cgZuURwxBuEc9sAsVi/+Ei3bY+poNzAGMJds5hSRjIRpoIp/uX8Bl8
9aycE5U0HXqNNtsYMGnoj9N+ugC4bRa+/z+MQBX1GjigqP9I794BT1Cgdy5R82PV
bXcqesQLaaKRfkRjPt08qO7D8D0TqK01FG867aIHxajaUR6nyRfBDxtsVCToUj9f
nXhuAHcMJ5kVYAZ7ckRT/P2tNbOO2R1Xfk1hp+762EJNKtWKn/c6sWFM8qaO4DEc
M+a+7vVGiA7nnQOJwXjKJpo/Mlg+cfAWg7n555PuRBkYarau18LG/KF0IiNOBsyQ
MtcgaURN0tC1PFvc2bDl5JvIp3wd78pcKtZ75mv+ij41u88GmQDi05wzIZeguue2
Epk13EPZPMNc3R/lfJA7tgGay2X4bCk3PhsI3tZLw6cvgm5PSXDMj4MA0M2N1yPq
Ym+rx5f8sTiMsWR5ogdELwNrWGSbMq2mzauCzPaJ9rLfe973No5DfeigCj/0VMl/
P3R+24jF7GsUwIoh2H5ZNhRxHPxnTP2Xvj1gcE1FsdwURnYGqgV6jAZycRcz6OKh
AcTu9FbYBncuFBtIGcE38kht/CB4DmDQsQC88YekNK5dv8xigL5fyR3gIPVTYDXV
je9wfaOcrNGeBoHU/gIwaXSQDix0u5VlCtle/6nhB7hsrBNvQXxSRWx7qLb/778P
/SWW3g+Y4cMnctgXACsWivo+WrSy0p6vJMUl3z2IGFw5KUXvL0LyX/wRin8uzvVZ
Wn70kQ3bPbg1Nzrf2ZTQh/BVeQp7RnTP2L0beMUNWQx49WbKB3T8U0UNyAlqF0bY
UuHvGN+Pq4lo1RJ+hLfv6h18UEwicz+TWbLlJBpfpyc5kCwmnFypeIo8n80puH3V
LRWjO2BcA2J26C3RljlA+0RTGXjZPDcZoHwp+DSwjzmBWJVTcpT5RoNuuCtNbSSD
u7HbHvl+f7oF2whQbBsrcWr4ypkoLpx8twHA02+/1w7KUi6MqEVyXYXRz7tSYhj2
9chJ8e3WkbUrSSHWtsAAnclMHTUW/AkQ8wHMg/jIMiV5RV3I0rSPB6Qu+9TLm6sG
Q8NKqwA76DoFedehMW9+hfNCwk6+1ubnVijC7hkZFtZ5YBsqz2gataEt1Qyu64D2
PvTOthAW0gTJ57DHtVDH3/Sr4ZBttS90DMPEG7MA3p089Pxcf/WMyaViLL7De69a
bGt7QqSWbF4SD0NFLdj321YjDChA7/qKAjs9YviY4NRJCz4l6eK2O+f9ZWngQ4KO
6DJxwRerhbuvFdzsx5RlRBDI/6Za6OioZPdlpd+HU6uyDGRqf1Tns+l5sxtTCtYd
NN1mDBYETo28Pva5pCaZtAkdvTquhda0mC5FEwEKzUf1FB8OTkXlh+jwUDKnuY9J
QwhDI1KyhkMwhEv4G5nCcD3taRZNtyY/MCF9j7v40fwVO2AMNtHXQJGafBocKNPq
dfkvjTUEHHsNxg/MUis5yQ==
`protect end_protected