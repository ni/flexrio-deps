`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24384 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
TDkIdcJUWDKCGvmrQYRemFt1n51Umms5ukK7PYNKo9W46eQiCaj6HNgzqC4na1HR
7Ojf9cvcAAE2bXoEIJON7KC+CT8H9UQuUvEonraZ+UZ4wPbHVeMEvKDxSVumiBiv
QTjV1VII1vIWDRYhy06D4evye4wjXjOhNdRXkHLI0nnxLtN0t1060JDscH11VJTi
2yqQJphdFZkkzmwulsXwhwFTCl8Kd6txSYvWuIKZ9u40Xo7TGgdF4hE4nLBuTujw
gVYilXcwdO8USbvRvATHWvLkB9QjRAQXMoZGvVh5ZKnxtw/+3+2FLmyp3ratQA2z
ck7ccvJq/U2jAz3sHs6JW8iyL96PuVvxMhvQHQFXcjLIsS0lDJ4/bNA9cc9lSkUJ
uAFOHHD4uxw9vXhk98+FJ9nhHnVoJ+xxv7i2U7ToW/AXxFNM6og/1W87wKXW3VfQ
yt4CDlPhVb4NMqASICwEZp9fHCqm1JnTd9BJ3yI28OiembspwxhC0pirAPbhFTrZ
8zqPZ1e+RfvvLqr6z2mrwEpuP/J/cqY4HePk+koyOLZhJhcs1TCiS31wA5FMUZt5
LwdL3CnUq44mnY4EaU4g0wm25lsSJc3D+ABUn1ipFWFHjE23YeyAyQ5HW20AG8Az
ukabVigEfRmV5bCvDwKSELXO6JtoLc5TXHPZjygj6Qv0JmxBSZypRdzUqV0DlbTv
JQY6JnYuXWb/iK8xG3IkrBlSF2JSFLKrxjO9/Wd8LzNuJM5ZM+QcG7v0AZHoWuwu
ZAHCjzFjtTiX4tM1hFFuxPJ9YjdzvwCVcuCjxixt4OTbBQszT9DPWzE7EKIGuyu0
nqbnBWj8l+g4u/SmwIsMW1OgV2ZKHp9nEDJx79rZgNOTW83OXx+HsyD6kxwRrk+h
hHMwYlRmtS3DZLx/KRaWxXbCPZr1Ys5uTe0EAbHG5jdFUWklxQjsh4/7WYzt1utj
tCXvqk+9uNCkWh4EmAUhyEwgjO7pNzT3QEBoZqtMOhAEme9gY/6CCwKUhe/F/zUp
ND/lO9BxInFgRuZbCfFwd761vgGcNATQ7zQKV8Emqs9r4CEq7cBxi5VBsOdx6AqG
JE39S8yJXVLc2hcA8J1yJxHpUmMwkKpZFcCxhurgqgkKNs7DI4boVv4/GPyqNnL3
DcvEnm16Db4PYICTKGqufIBIktvM97l5ejvS6IY6ncwfCPamy4QzADSqU6TbczfU
Dxyl/QJ26U50mbBuul2sAlYZyk4aRrq4b+EgGNSA9hLiT2rV0IYyRokOX1rbDe8Q
iH5B0yS7VdAUVfhILrAscYY43Sz6EEadAvJuXdi8+5EW37v05hAaJYqHSBTUn/y5
1pvz+p2VXUGvBRzn3C5ZW2Ml7BWpjQ0RsKpEZBHe/RdR3kgrBYRfiqcPbOkS5JF/
hoWAcchFw6Wxb4fJEWKXKbJjEs1+aQ4v5IrSiwEOHMFn04mJtXIbrD8tiK/31gY9
ShU4O6hYFq7Mm4IEUmBBjyiGHCvYnXZZvmbwnlc+n3OZCsrgozPt+sva5bSfYDXm
0y0DvEBG4fqOod1OthzqM6+AtuUmtFk8qW3jswG4yqFfN2fT0wQFFLbkvKl19t50
dbbFdckjKauzfsF9nQp7I3FiIpgFTMUxxXk+rmMMjLYCFTjdhVrag/WsM8OgPvRs
5c916gI9+SC3pY1HMkHB1m4fXuFYQgrqRqBP26Y2bN5cZuLerTTTSHV4QFCaFmM1
4MRVon31wHl8bh8gOiCRwcnNm92oZChHInnZuQ8w5gfj3hCGZ97zh8aWxtKanORs
OCsXBy64z5KQQmxvmpRe6KqlNHyqU2NfD5/1eQ2ESAE2ExI5416yxuSwPshRFkTn
ntPAqB3LZ31vmQV24/+rApNqlFs+HndvSEOPUiHA0krlUx+B9sG7fgcow9g4tOcT
WADiQ+/cEGxch47V4lpfsGQ4ceanuQJbS+hl+d5YP8veTPTC4WL2h1dj+WP+rF0e
XEP5DYSV65FD2kD3E0wC06/AZRwBImQeza5dIcDb3jY4d6okITheM3FZ9/jT2LB6
MCak/wsbPQkenzZ5y/U172opJsn4YLCUbkRvwB/czmi29g9uMgoZJ4tmDtypUxf6
sCRS6WWo+FpQgWkyD9iah/SA7ImuT3JFVaMpF4Pu8oZ5tfSSGpcLGAiCsP3cPHwa
gknG+bAdvbfVPaxa74FoieQxjyWx3mzUFkm8pGmtT8KQWAeECsR88QVcNs8i8OQ/
lVmznBY3xw8vIHgpANGLeq8Td8ZxaZ3OPyTL8hWduKS3IE6Auzxx9//WvNYmKwQy
0ZXyvG6GzFCT3Uqn2GVNJvlH/n2vlL9ZaQCAJiYJuyGPrcPubCpm4AXPvYZ2/y7U
SC3P3g47TuEHnOQbfx49N7Szenpt1zQ+pDzNW76nQSHA1nrDABGu3lJKnIUtaMz5
R8E1vv7oIgdhNLU26F8fXvhWp+poexsLAIKZ7z1f0ABO0E5cjihjfClrFkwEuyyX
4UJNxgdtvP4a0Vod4naQi1Fzgto/yAF6v0gjazwr6ju9vn7JGEYv7qKV2oGG3PsU
b5hTqTMpKfIvQuijLP7eyOuF+GZjGFh5AYQm1gqUX/ma/D7MSRZMiMeuDIyRJhJB
VJVVOPxTXYjZy83n4Lx8fCM46FFzhY9YpGxj98tIFyypZ56R3lQww0/1GgIpkhqe
45w/1zz18//XI3grig8+bmxBjd70epRd44ss2zQj/JQezgBDV6T1WmbNX9WB/rSP
jkmqQ80PgiYxE4CU902+VjFA3J0QEyzJc5dCX2SgIR5iiaADTDKzkgq+1Ied8q8z
hAaXGCmdMqzPJwPrCJrIjlR+V5RtgyGQIYHCZk6RYnoFQe8dk3xpXTymj5Fqtbfx
XWK4b6aHPrk0RP5nhDC1XW3WzpdCnUbfG6cmAyWWNg4IbRh1YOkq9QvWxw0XO/vL
TLTMfINXneRewoyKKBvqFTBFOnpW9CPuRS6FhEGIneOUrMZ+acGsussBHlG/fwBn
7r0quMBcxsStJfU1R9KblzmffvkQugNOljW7B1uMEztTUlw0mh/zN69sxPHHPEFh
3aCyIhwvLhnaBnRx9DEO2AL5hV8eABwQiCeIjnBmDG+wtI5ivz3dCkP9aO68iF5P
qLH5GAVQO9FXjcXm4CnEcnIojye8H4q7dNq8jdU84NZOQGPJGFc6f8AppS2nlI5e
7vG0jLKri0zWCJip99xbx0FG3kKQXlI8ioAf2VPMwe4S4iepqieUUAJ3G/NNt2ad
xAyjoVjeL8rRUmBx9YNEwHFCqsJemE6rFvAcYfRGMJE+uUmz+pi0zJ2nCX0pn6Xt
Z6FFFf2BEmUwcsfinDsfz9X3nXmNctJODDySnluAL0KPnexl0CvAkOPMbm3bubt2
yV39p/50XU3ut9aTbOGGQy/UVtcFYP4au/B17asGIv5cvTzXktuz++Nqaw7pNVQp
eTlhA/0kqHID2S3lFv11dQVjCFdDMDnivbhziOhrxJXEyOPLoyMV1mg48rNg+Y9f
1pdllQRmJqXwIxqr0XIBO1Et7u7q3GKTC1EwpR6AUEFunibtoBw/wij1q/honciE
BJRzYQRkOb7WO+ikMhdQN5UP0sa0It44k9SY88qrlJQMD+ENOah8h0O0wJXrr1aV
EadqqoWss2GnZagchnLWDhli+r3lbLIFLpniKY5OghTQlJDzk4Zjd9rAQXtoH/No
oMRJeaXPiXmyCI6non37b5O1pHDUHUfdQVMyVtod/YFa55kTs7HHM8NAaMms0oVZ
5h0YFkQbpSqpQ3In6/lsX/aWUl4YWN+H1SBcP5viSjFEOmvixKJMpTOYQS37zxw/
PssYWIm4c5YcWf5Ft0ez+jZ0u6oReXFiuuIuc2L1yh2Qa43ow/kJbfdZTB9vVE3A
V9qCY5ZIAgsW5lbFMBcOpUZS2dGwYGaotDOYFzgh9qihZruNuV3KQBurmzFPEKlW
TP1Bcu3cevcmq90MiEGNO8SzuKt8u7cH9vxQ5DZoiHuwzW7+W9Bso6abyFMGWNls
RPJAnPXoU2jJL3KdLUfmxbCcRXYBCq6ajWllu2sAkEBWDyEkSgFypwlp5KFYg62U
lkX1nEX4p0uq0/3ZnOGKBpx9BQpF07lAyxyx5baTgKYU7pDiO0HhKEy/T17NanWa
VgwwOx7PbdGkn53isTM67SxzTSPaMsBCThWAilMh7V1hrKmKApJHCiMpbXI9dyuF
+R1yWaf8Tiv6Sn0ZIbMtGdgRYRxAIozi3OQTJzdjvzefBrOpeli+pAFCnBVMYU3o
vhOwkCLaoUjaM77xIWEEF0hQT+/2LUY8rAkq5O5Co+bf2CFJX3R197CWOpY3erRd
qK3LAeRp8I5CvHf3ScX01Tkw+a+/k1pIC++5cJduxNuhEPrKBKLcUtgSL62dgrkC
J6is1pQ0L3cKnKQFjQFPMeKl4wEJeLOEFJ21ChSYQEf5fTxv1RzcKqfsCquSge04
d9KenvHgU9uIqfAccwlo7+cSaknbLQfONWxQPVYaF06S2vc3bgwRcdn4qtKrLhgl
lnlLRjEbTlefJAzdyek3e4OqBXiYCB+NFPkCAJXOhFWI3SjxUA87srA+STWbZwCi
K/yVdxdVvyKKQb7Q0WGKX9nQYYTCYs9spWN4anVKJhTHrrlWhDqP0dqzFx36tvrZ
cBnGII8EgiJfykAHlq+U83c3G2S2TPfFZuYtfjInIKURT4Jl1wI1TWLM56Bw4hv+
K6NSY/JMdmHXd5pbf5MtEhC7o039tc/AM22TeGebV43rtVcTkQP7jGqclpgeKZc5
HQ/liYZcgLNh9aRm2G2M3b/XBpxF8Tfiyz4G+fudA0caiK+dadcWiQ7gGc5RaxXA
HctKoHuZtOJmcZP1q9D1c1JiRoDFzHFm2n8/swKKxu4dia6/TNc5JVteQgcj1IvU
bt7BM7QfZqcsvx/CKwXhMrwuVylfmtIl1JOU8qJdT3epgc1PX2BsxRJE3aUEnqKZ
MfiA7EApPcMImvEizTpx1CT7x9WLVJsZzZImDKtW8Jb/OfFj6ucgW6lFNQJzBayh
xuyuyuDZAx86MaxKSn16JawDOk9riQ7pyufPDcLg4NYNpi7Ov3MahuD3tbIaJKsQ
U8ktSwwpfqY+awUBsyW1ChnoC+05+cPasDOawJBd2UAcqnaXy1ZTYCNAlNc9uZXP
zXJkQF0IyJCdyEz6cR9Vf7HphT8CIECE0wflfxe31ylgra7KSedm3dbrU3sPitEc
69qkzS+K+qpQz1D6Pz5LaAVaaKyII/IsX1FVQM0yRGvecFv9H8gCizPgQg6ldi2w
9xzSzKnwC3V35QQknhQBM7zMzdQpc9tqrGk91gIphmA9wC/6iFQkiDgkFsIhejy2
CLyg70/lBQiPJGaYV3Zx8r3sd99IswCABabRyWs2FO2EJHpfVGOca41pgGAlaNAk
KX9cR3QfiGrpbZa4nKWs5sFtuxZtXISOjlGiYhl2BCrPVC0YfJoKQcFUhTUrUOkN
5TRI4QFVwgYeZUkCeIWM1F8nr6aFYNpjKoudFUEKbQgJaorwKy17+HHjCaKfrREX
FomidqwV3nNvjZhtPWBbHMGXMUjFbrb1wpgmaFv2fdn9hqHsy8PEDUlQi2wE3Yiz
05hLl2XEHTCEayOz+E3hjKvCoKYODGlJOyFOyVwFKtFTgmGAb3x0xN1wBRCPH7st
Ef7IohDSlgjwWOkJg0CuB3wVuxtW4IiWCVPpCc4geevB/R0dXbt2nLB2+g/j2BNO
0yIykEE7ifQo7Xrmd7LGpg7e6W+ddec8OiIuL4J2BGWf3Grl5Ty6vgXC3maM+gfF
JFKpXJgolNY3F3x/T+05+mBLuIfohPIsXqxWPZOTv6FFpJuDyG53iJt/SSsf51wM
+GbJWAD/P1Ji5P+yCE8wFFiIBJ4MxHB5B5BppU4Ozm4ERmi7BJj88OONoJA1/LZK
y2iyv3J0T6ArLnyfPmJ/EdKY/RvfJjNE5raKwEamfyfyTWvPqkbdXyxnh8BDNXhC
noXvIeRRi4ZAx+WtIGxNwPn3sESvUZ++cKu1Zs34lwPkVCp+qW2GhEDyx32c18I6
t6vaRM4BlDM8RrGXerLO9jbb7uAaEw9YAK6GCFPZ5tGozMPZfp/A4U8gNAoIg63G
On3ZASXdd/zOz7J1sgYhKB/LSOmUwExGIIxmJAAIyWZeliY8VPVUHC/9m/cMEjkL
EedE3g7aU44PVdAsFV7xBATL6CvxTVf5f12WzHPBK5BzQI8zBvtARIEAHssuaPho
SxHQmS7g+QNyYcIg/GpMdbzJFMCKsuIFQ2d6w8CU744MFC0Ye053BvIKlYcZ5T8e
mtx8TTcJMsnyJw5e9viC3PgxBUuJ1dkHHB9IB9arTzWPBoSr0+2+KU6MJroo5xxp
IxuwX0c6UCv+g370NakAcmH4JE1zYuB5QZaJ1pM2SbDJcxjHxTAMOyDugMqXjiXM
MiZg5E5f2Okaiexk9T7d5H1nVv3nCtAx5W2EoG5SAz4/lExQ/UUHGpClFXtT4DL3
nTl31BChSyQ+FcLLOqKWM4fVtfbbHWTLEbZxPmguti6sjKEwQOKrSRYmy/H3WSpz
188GUy1c0x/WREsOpxQ2a7S7i7ijH2e0jPldsHNzZpe+sTJ6oqL9cygsbhyEaFzJ
hUoxdbqPQ9zpdwmS6ZZdAesUwqX1YoZr70/Irh3AS37u64JJ+CEvZbANHlShTIyR
hEZoDI5gNIImfMNVs3X59neXoy1ZRrcqss4XX63IPJ5+1XSX9ZBEE44K61MPEtBn
rLZkgWN0dC2MoTQexm11+iESStoXGF2iDLFgc5LlGa3uJgEFVAeZ6eSm8FdyViYw
WW6wiS+2xf6/FC4eqNfX2j3tJ6+WR7Qg25Xko7oZ+XSAxTzztoxKgBPHFUq4arY2
QLYF9DctV9I2/8NYs/22uIyBWCdlSAXdQ71VUNGvAsFmkqXAvdFsRRxnHqVLScvb
iLmNGMNaS7KRfo0NeZPLHqgf8sRUmup0oK/sAQZDk5a0kH7ylb3XQiqsb8VLBgUG
oDvN+Tbn2vaoMxIBfqSC6FTkK+f4XZmltiW4jGU2qKlHQR5iZM3oi9ifkFiXexMR
8MJmAutkqNJSmULECe5QnLh9f4KRgke2xkC+Yz8p7PNooUBc/5aOROo95sVoAxdU
qAs/twlDayWbCGkBuXFyeHUYj1INKuJyWqAtRNVXtGV5i/GB4+fJFzdcDTCEgjEY
mP/IisPJQT9ReTg1kZ/S0ADGaxJ350MWm0XCAwkkHGUhFHj362Ib69ZpKmcL8yiR
/upYW9pbLDSC5Z9VJEroMCgN3t/yq471mP3pfO1rXtNLBAGonOm87WFR67It8bdP
9BU85BkEFlkb77/nXvKcjvK3lYNWTYtw3ZFsf2o1o4HrQF/J+pWdDhZl+z4IErzb
4a0yf9oYr2FXbx9tdH86ZKsylTukoBpYs09oKss5pjaPZw34lAN0f7p53Tb3UrAJ
jXRtCdU/DfUBuYfzidehLDxl1mdz3R8IJfxbKh0uaPxOU99cPUDzMPgK4gYgc9Qi
m9ZJzCooAUlISJFKwiLS77W/0JF5BSq8hmIyELINTz6DPMJrKfi0bIQU9vlFZxwI
PZZj+9xo+jpMgIjz/TvrbX9rh47LbtFacfvDnWyYT3VxN6t5cL7T9/sJlNqvu6cY
p3EeM0BRAjKvh6Wm1xmbDQyQ48Er+iA+nTFe8AfTVCDv8DSkET9bbq0erS+328LB
C51YiaR0soSFyMNfsutRtC9DA77j+kBM1QRZAOlnoPcftnUoJgFaoSH9jSbHt+L+
O3ZAZVVq65nL7NoxSLp0TJ7Pu35OND3aByAFyZ1PZZLJuChyVu/WlWVzegQHspHa
wscqG3L4cB8T+CovcOnzW0YmLqGuEjie6CrCuDHimCZwaCq0agwcRGC5x/hRjcrM
L1hhFMqizfUxp2rydlF4JwMOEwmKUYVH3AaSZXLbogXpDOL+y0elXqNk1ohFVdOR
L61I/Ggy7P7QlbBbvG3vnkHctiX2qZuZfgxRuHO36R+SL9FsKk4QiacabxpN52y0
2nmd8bmUkavGGZ3m3/Ds084AAHJcA/QsTLKncQ0onlk16k2jrKPYHB7ZDY1Oy4HV
sXft2rJnYUmxYf1bibZcOYXwKm1xCdjmYA1Dg7FBPe3pQKDiCpZXGWcNnpZvMRSl
plFp0mY6uI7X/tG0YEpFHrgAP7ev4OBgmhGTWF7zf432eox0nMZ/ZtyhVif9Etjg
+OrBa48yqMN2b2yl13ivml8Oz6aF3nveGnx65RnLVyW/OF92dKU3LAm7xJK+Gl+U
33AZpPOkHGDvR/apadZ+JI6KCj0dJQwKzQ6X6X8r04/qD3zYteEkwih/AKX7QK4x
ODpYJf+Mz8eeezxdLAK0gcJ8gcyeQ/C7qDuk9anAu7J+k5EadzIWgjWX1jSltEkU
B8S0ITo4dlWYImT6PfP9dzf3XZx9Ot5fSY0Es5jWlx+gIcHoQCxd/tQXj8vgSIVk
eHNVPLMpnKL7ZRMxduI0F5oGGsXWzzKMhgy7CzVDz3KlYftru2VLW8cD0vWjIaGn
LrXu0ynImdOaSQY61C/5whGV1/Q1Hm9QjCh7wfaRMz6zigcQ5euvpny685yQKMTp
FUKsy6aghadPGI8CbJTaKJt9TmhV2APbtH3sEAE3nEric8/xy/6vJ5i/5+Fii7xn
6VVn87kR6bieVZM4oW7wNxuxdxHO1kO0iKhPzqaZ/PbI9TT1NXcIedWP6HIi/hjG
Qtjc+viMUxrEVNRqQC3J3pv0sUB7PKaSkC67RLlg2d5UjROMtgHPuQhIT1u0zDDE
Stxf+PYLVXJB9pnKs7ROK6DgfRzSZxu5XlXpMutLiGIQIfY6gC6QoQ2po64EjN2Z
y3webdqoDPBn4v5rjLKoLkI16kQyarP4dwZDxdI7peXiGitvPYbDlUl0fOgDpi6S
oQwqzcs2vmKnzwKfYDV9bWk22PbbtPEgahxnohwpfgGKQTtFkmcBu9/E7udKEArb
ZVVYpqkaPj3vDDVLdCKWHLjy5dJtpfvLc/3sNnAldFaK7tYfxwz6+jGtbAD3a0q5
5E8rbNEAv6fmaM6FX9/LsmvJ6wO02jk2mZ6ZnqDeUlh18iTsi9M0Sr/iHMuIsJxz
OzmoejYXrgVzrglMK+eGwIfXUkfpeaY1oCbg58Q7qzqLze/jJkvg9Vu/bk1FZeQy
iIKZVJ74VGnVqhYyC8jDZUZNOfvlm/DKUAvBSrnrgJbtz5V88QCjRcjDW7P7jkVd
L7X6F1VGjxSh1EuRguL7k8Lpsv2MX8C72Md2477n4jfTWjO0IlDgb+tRWovmPhEF
g9z3mvIpRhP4WKhd7wMgCIOTMfZx5pU4QrIbOkpR14KmmR93ate2ipI5JArRUl5y
+x5SQPdK98ciUgpS0QnQAn54hil8TfMp5v0SQclw52feFq1WGVr7BJVdwRPqNHwZ
eMRgScEVghgeX1l2N/Fl2DqiVpmv8352EAr+yotHhWvBfVUHRDwAkEXk4D7YziO2
X9GDt1AzpKjmTTait1YkZppmj8wKUTGfFJSUhrlcSv1PaUolZb9A25U6nubKSEBI
is54WMw+L05oraZG9oMvEtWgjKhxp/VJdINlfrlnGP+GWkawJjVMan45qHZqDQMX
EqucMxS73F/+9wahTwTMLBgyRxFsZAm4dKAmK2BzqB1YDCRP+lrJ4x0JwOV1erOw
fVK201mvdkh8PRgALNWujOjc+OrMP+WC7wi/mEA3yw5GVDXczHwCc0q+co4ZZ0/u
epZWu7ps0AULY0YSB37wFr34Px4Kuk4y4Sv92OGhApmZoF9dOU0nTAmY4m3thFa4
E96Hf1iS6uVBQd/IjsCkG8SXQimKpVjJ06dVUSMrRm/rwBj1azwfR2bUprUVJKSj
0I1naBOb+I2ls/D5ApMY2Qfr/CQH0hvwg11KLSdY6CFV9BwGx161FRk1bvWHsiTT
oe5DO0joKzFQOm48dlS6abZ6dtPLwvPZE/z9MqTnpzD4IwApBw4nKtT/SL+ub0/P
pp/SwhkUS4f9svGVM8c6vHPbTvTmHzgwdwYoeykOglbe1OCAZUsx5iqd2MKjIqkh
VXd+UlyBHLVUopSbf7zAZl/Ixs0N6nxjkC9HgscHHt/mIWMSjtWsvSux2QPW6A7i
YuHLbMdTcHaN3XdYgQkfQfhOsGOQVSdFzdSYgkg8gjPsOQj1Nf/xTtDN8nU7yn3h
6TXkI0wGUsShVR2l9hhPwWL2C/ME71bkSxXSOSF2rspU75ZVn88YmAZf0ubut7Nz
EZQYQArfwPEcAx3iMpfT2SuSdZXsJ37AmEbvWI6UMCWs4swAMuY9sPUgSouDXAS1
u9Mu0fFXkalfBXBGUqGPjVmaSdt2Nh68R1ywMOUuFjnOnP+u3xus4bf1bRIHuQZH
kCLWlz57AB1fI4klecgZk7ZfJMNZE8IJjK9OqgEHP6c+wqD4l34ZCZ223IM1V6ow
IUe+ccNnjqhg+X/OBzyJxfgfMgZU0hH6lpOnnQxRLbrBp7hXsFdI5QbHvttq1Akw
sjhEmapjRNrTz1BZWGE8vTPv8rc0nIjr6KI+hUxKE+uKoZg5cPq2FHVjhOyspEIi
6MYiNZWKmpK6m91KKYXe4W0RK24ekrONJYG36E7ZmoQ8MD/yPJEwD83+MROUp21E
BebK8yIuX8tT2edCgBcGnpZj7mh57anZMICYjmIAlXY9m/OHgEYMJ6dfvNgXpQOF
41TWfiV+MfB+G2ew/kNe33JBdGrlwL9T5TAlbTxQnhnxfMvL5gcwIdFuSYSijW4b
NAiGh1SMfJ0Aev0conT9V6ZwY6RS9ZZ4HJae2oiTeETwLPKx3Bl6wMHD/9BJgrDC
F1zI5v8Yky7jvhKSaN1SvQv2knd3i1+S4Wb2psAnzoa111nauY++NVLmTeaPrMTI
jfTv+nfsVyPCDgUcZ3sxQvbziOgxdPfl9YsjbrNHZqiiDofflZCiLMRHan/IFIzb
MDJkZxcr+u9Y5b1VfxddrzIXTHA3TEeb7CJtDgqTdi1jgL6mmbuz0JgTir9oPbQB
OOO7I7znXLA4UezIEcZK52zSGV7oX7Hw89IzzZiSsZ4ue1vqYBGwqrN7rta7CM36
udQ9hIP397vhMZPEECYKnlNO6GcuyWqokOJOlk4Hva/wRZMBu3twm4YAjzS8qqn1
dR9+7shToNC3Sk6Q7kVRXqC+N0+57XIZi57T1j6q/tjBBbDYul3E9ukhrVk3IOlg
M6wu8Ga4sc4oiQ+pX61lzJW0UowPfsYj8RMxDWKSxS7MfHzF+jyDWTaw/7TRsCiJ
qTHJoYzeC6F4BmxpfldeZrcKe+QQpwzraDYHosped167wSy4LrM7WNBdf89XPAxj
dqt08QtCI5dWRYC6LA6S36McJ/gTa2K31f1vFNfEXaQtr5ypcrYNxAjtNDmMrwsa
JVxd/4ej68+Eswhw5LHt8wwTV2DW793zFXSHb/ZOrtRaeMM1ByIwxM8NSYFLbh/0
rfCDjBI1fND4r7dTuF5nCV3/+7zNbsSPavqKwFP7auiTYYsNPf4vZw9j3op+6G2c
fO3LUOJmeOl5maFqgYjtq3dsOy1B5IoI7djFRWkY4PpvWBQcvLeNw9bzzGRH9/w/
0koA/7AUiDRzSj5Xdm7FzlFIDzYXOY35moUggW91hFFU01JY2kbNv8HoMvevu+44
iKz81GoxHn1VLCkygL3wS0bBNcfIv7VfEjKNpolPhTnYWI+pROs9aUSjyOCcxqj0
kgpu3hsomY2IvDlaVtslp/UoPs9ukxMLhmnbfxE8uo0H26bh5ybd19BJOQLiNtHR
+I8nM9RkTVzCFreqlzfADWVQ8K3gAlrSzPRCEWXiSg8LRgRB7MHOjYksaO6LGaoV
6ZeZloFugVjWK69HidTIXGYmpNMGpuS1svoh1XsMX0DqHQMwulZrPvfMS+oTPubF
T/m3jFIaS/feOM137rpAJveEsVhWAabNFbWIPWtxRtkW10UDSqQVZaT3n8F1+hn3
6/GdSNgMymsIV+jH9EocVkuapScXuWwDEUNnwAoMOKTfRAc3OyUCwn1FkQdxf7+q
PUOiwbXw2gtqYkiMKhpT7l6JOGk04Ixz2dNXDul9Wv5Re5W4uf6QnfT0y98KlULT
H9Vvo20UIVlRWTpuscAT0rz9bSoULD6/DrQKrWvF+dpO76hkEr++9/AFumQwn7Gq
zh3Kmpv0itlZdhWXtC0OrN60SAkE4KPNVLV6xOLEN7Iuyn7QuDnXE8YXLRcu270g
s3S35XE7V8k9z5K1gkvceRackZS+lu7lMo3xRuiQSFYyfsxoZaafecaDgdNNTXPA
sj7EhpS6XFXGAOH40cPtmV5dDqkVLOUxe0WqcL2DNFZev8pkWlZvLg3IEG7Y2o/s
YEme0Zb67kIHCeNpT7eGBedSf38IkyLOwSsHYN02iU434oI5gIsZuM/ZVZQCUJNp
+dxDGsfDFySyK4lAknTBQE23PyOczOxTP91HQL8BhB1z0kbiIo4r8E5Vh0uzsbqY
XYvEh1VLNCZlKcednPHEO0MxTxJ6w7FZMxqzvmCFK1xTbeEPSgM7vGAuKzRLuy0x
FmvrODQUhemt3hRR8Gkq9RbO1nbp/CjqQ3nCvJLDDafwGMO7g3LxP0qh1z35j16o
KD9ugimaSuqjx6qQ5pIICsLm5bBKJT97rST+p4CQxKmCKNPwQfRNayGqnFVgz7uX
7vhiApMzk28WQ2/L4T3kP9j/P8oC8qcCDq52DaRjq7I3SCRNw3KyHmOetw8oUPZF
cWeQV9k7dOQiPoBAEOSdIYoTKiaaGypIvigEz6UDXskN68nTegUK1DZhjtMsGbR7
TmNzo1Wt3w/ONZwpXLdXwv1ANDW4YgRogVCq/PE1T4lj5d2FKjkw6CQYPx/ddbz4
QlzUVBOHVJAncKsmqnadoXN7Ni5ehCb0tZa/SL9AtGS1yS95fYfMIOFxj2caNAz9
N6x4ec01YtjZ1L9GlGktiR0Y4qsJk02DBvxl6zCogRcRSD+aqDhS92gTsMSw3yS8
uHm7HmcLjxUWxdJUq8dRnP/oXvQGPbWmhiODEoUmiBv12kG3C1lONUwnNxhtKItN
F0wAvaNsVHoe0OxlIJ7wRp3PPIPETaseEC00RaspsZA77erVUPLxA/743/9yuS5Q
aWhmTUSVZYmxpukta4xSQE/OaYuHCMoQuVeLuWMSEHAI8QoJ0s+jUlfyJjgzhhr+
GbIobqjhFj6MQ0qXlso99LbYFHUk5wnqrNjc+cxfQch/4a7QnXq7d/SCVJBt1u2X
JVveZkp/g34ZJOmjnrN2nNfOa9CsOWvuF8+b/7aVyMnOksaGc9GoZsSlu4PtNTpo
9ZzjJqdgu8am/n9lYcnDDojSeFv0jFyMf1HzFkzX/NGBuaVrATgxzmyJ8NyekSWi
kgFnVXmkbx83hv7tivnJ7dGehTU0JcNMIcOxEpL87c9JWoIt2Fg1BMqBYWnhh87p
bx+xiLx+DTvNlvpfWL4YKAAsbhvdqaxTve9eg7JtZHRmxUFCy2CrpZYHuD/9z3h0
fxyhvT3elQY+RAJUeaSrOt6r0MEBb83ofgmlvatcKW18H1DXYWpFqVANsbrk3TXr
kjo3Nkp1QcTaKFU3qIzO3fNlbWco4lWWL7md7GwJpWRAUtJ9a3RzEsa7fa9TOL1N
HR+7U56tzd9jLNaa3QM8p4NrL3QpLVj8oQz/2e+boIpoLvHuFy5UMcZfN9W3fEyv
1PdweDiNUvLS23UVnbwt18/xwo5gT8JRMgnSUvg3mZdYfVmWomzMl9cpegM0UEAx
flwy8pVpzb4QlTcC/bBHmXmTdnBywMUed0cEaNEYo/gfu4ERrQr25F3abPxyV6Hn
T2IuzuK+RTeKxs+6tLJjCse+trGCcuMgay8TjbGz0cT52DI+mgAjn3A8Z2gNOaZU
NXHukBQPej+f8x+HnT1I+U2xZD3tEPWqd3/kDS+c1uYKJLpNwC0GIaChVdvpQU04
ppbcC0vv+5l9zzCIE5IRt7S/+FUYdfBvyoxt7+qOM677EJdvT3/7F/1EfhV0cj80
xooftQTxdWucoTQVPohEruk0k/jUe+JNK+CY8NjsXUHSZ1oe5TwSs85GC9ky2QNJ
FxAx3qLPQik9EXdwKcL6dywJRMv/VQxFRiCn/nDaErnFzm5aEbCaKIMj6KmUVUs1
r0uPOyqTPZeG4YdjUaYe0l0yz5l0WF1sw4tU35fI6RfBcwWv0AVUgfMpNHZE70fP
AKhdvPWg4g4S0bRUeeb56TM5NNkOKuwNle1NLG2FaWBcVmqVKtbA8KJoJ5Aha25b
5+JDK3dsDiAMklf0sNR1f3MKT1a9kXjXwuFGH+/+zL4JBQAhR+EI0A0+2VHUIrUY
s1An+j19SGAh6KOuaI6jo1DZ6lOt3fLRsbnBbPhttjsaaAEHkcFMuJlV9vxywrnn
Ndg/mnvD1e1zV7Spee995lCl/kjJmYj3NH7E8T1/RqxLT+LTxci2sik29za2Ji4T
V7tmT+uxQh7XPUODoKp1N3EtpylixkdkiW3HFd4sE8BkadMSeQG1BEUXfzwF4zGc
k4W0n04k9+M2o6LQmo8LW+2mxWyTOLXeartCN3dwrlw95Wujy9IaSGdwGF+Z72Q2
z6OatvamkW+ov2qjxbxWXD1NmRXW87v0s/n+CvIiMAHeb42hOnxAYOQm4us0FQIn
CM6O5LDtNQ9Sy9Ryh2NzksVabFQ3XkLx5R7bb/t/eUOn0EO+4UlvxUxl4MgFPHEt
MJDOcNh4aI64X9SUzWc17vzy6/zwQ5OUqwwKe6BNwfteLtJjIf6sMlF0XVe1LX/O
LkY+xWPzMdRH8BcgcfzaGj9Ju1cNSaTEcesl76KUamXaX/tAox5Nuqr0dyHZZids
0n9j6JXfC7PLrulscF3qrVzDKG5Lspyohi9YaRDWtC7i+Wg08bHKIxUPbdvEjkqB
JmyF82EAP+bduUMaTu2BoOpmoepDYelAyRov2HetRv04wD6Q461ZRAc0ckUIUw35
ika5i5Z84FXHF1QZdhSCXIILAn5ICRVQbajuU5VK96GEdmWHS7FsaqV9o9oGXsuD
/9wN0jroDOySPKm5wKiQ2DzOxbp3kL2B7ht9rC94REYYxWHWiG1EXIvDk1af8wqX
fiu9rrHqx77C0KgTBt1GtVtfQPNK8Sw4ASOVsAeH3iV59TngUJ1qa91wpqctN/6k
bDu8cVgagjAB329RfjGBAeMZ0z2+2Px7Fif85EW8/5j9EOKb8rG8ouKrAZDp3XzB
cknxgx+OWFD5Y8TlnN0vt6ooI6nVfWLOAb21kYOfTBZ2UI1/TzZndZoOURD6QU51
tF4qYkOYNmruuf621b24G8n75jIKzHgYR3jrK+HMHCJQB5yUgz3xkfZpgHHGvwQU
3+rn/1YdQaHE4tGcCRNiwusp+R/WMJvFsgdWRQzndgu+3f47fjdZLHvht0Vavv1c
rGJxtK+ztQB6N3TJJ6gCYl2AO6v5rwfn6DsCyH6GC2EtOPiQaneIF8yDBEPQseP8
GCfYrZnqmefokA91V5G53q17bkMPc+kq7lpDSs07kH7KmpGkOFZEKTYg2vxNSFE8
JARSuM+i091pJRkigQTHSPGtyDdvB1Jmg8mLz/OKooCldQp3kxGTtg3CT5aqua5w
4H/z5h2Xgu48us8uAQgXMMI8At+wZveBTnpvun6TnFzOK883763qVyYQ3GJUH4eR
b7vyaNLcjfYE/WdQUMVntQPzyqX372itxmblx+UAHNruIUcxSuzA3OpKnnA/ngR9
opdCYfKs4Q/YFwchCTgUFPvX6tDx3zrJJxdd8tq044cDhVRBSGP97EcCMUgEqLJe
Yu8xbhfLqwnWH6LbSn/mHLE0hdc/UrOrdeDpo+LJqRzue+MVe4GJSpS8vn8S2oB4
P0eFU/2r7C9aDpiURab54NkJZLwylusIgkFpMIc2s4GupQg/VAEpvoxkFX84ndmH
/CCE1lkCGe96Z0fSl0kMjIy1ae0YF4UmsSUVh5DpdCV9r/Mt8/LGpxU6JP6mApJg
T534ULSJdBfVK/ho0Tc+st6Bj2fH8FpluCedfjyWJ4MPuF/ffAl2VNyfCsILPUBB
/LcMxUaWkXFdSR2td/+jyp33zhUN8cwOBwQPAMeuAbHoTD4P+4pyRzenIUt4WaPm
I4CLan5elDryEwX5K/I3qPa7Z2YOQo8GaRmyBtBg6mwI8zFRo0vP0VIe59GcQ4IB
W2172xGbw0JR/dT1cAnjtE3ZSp6altvSzMFBoCehCprdc1uBtR8THV19sDsEHOQ/
mqWf0RYKL9UJmyA2A2lgr9dNyEiqJYh4j4tv3U/FgkpiID4Y0INyd4cD05X/eitf
HYswg8+flBoHreDWFaGdGBEm6VysEXXPmxtR0XTyDA8zfQ2Ff10n5J8ipjYRNQiD
FOJL3Qym1+k6ASKB3yuSJ5WTMChpS0NJDG8lq1ueQyuOD4uxwTdHFU64J328ssP7
KjdAmsXxG3T/55wPJOsjAkfQgcq8DPV18k0RvO2VxD435giL9c9hwwWzh2D3c2sd
U9qdVjpcgjMU5Cr8WWiY73I355riBmsEQqiQ8YWt/RTAul4/OSdPYGSPYZufrEVN
2hGIxTrA/6xgjwPCAJ7yNLPd/a0KX/8orHa8Xk9YzWlv2yNhrdKDIrv8+RizzhFU
BTdluEIAJS3YptJIr3Mt8bFwI4Ik7VPBpzGuVkVe4c0y6wItUuhiZKc9R58Xivx5
Rp4KLucf9dEyf95FZhsrcU+Nate03+/3XGiXhAwdTbUz+bt5Cuw5ct7fU4pErpZ0
FdCpQadZyIIGm2UTKH8sBXgTSIMwCIVicof50ku03KB9aZcUKC6M8G0IpwEg5yyg
iZ3CG31NTH/MFNYm9ol7pnbsJMEI/YXPwnknMmXU/JQMf+fh0ljNaNtOC/ZbChNI
+gUsSAS52UxNCPky51CB3SmsJKyN5uFTrNsiGemGzg+aE5gbwOG6sn4STbq09gPY
C0JgeSoxISnNn/7ZeRVEg/M4k+nteUeAd/i+2a0dtGORpV513JdodkFQ5hsfCZrK
JOFgCnCQ3nspDSnzOdw+oXJTcSt3iknNFcJOQrmQn2PSeqrh2QcYmmY7Leku8Eg5
m6PNiXTe+pMOKrIhx5q3Y/zfcUyOGOyKt0VdACdHqOr4HAFXJOiDSqPyzZDbJ/58
NyApdI50+r/KkxEMdArz8mLux7MeZGQQ45dvnPefcK6BghbK4JI63enBimSWhUW4
HRw7p3XYXpF61uWSZ1lZ3yf50oFrHYJXX5lB0RnUbdRswCIQKVEQTCQE/JATRS3h
VKansmRr/OTCdFkUczoPh3VP5LdgrzGreEgrOCbhKv/XSRSVG+iqXybgGkY/U6I0
eOeTingRF4/38b2aRNe9HDXSi5H9RmPIdKRohr3laXdRut1KNJ4FMS0L/3tV/JWO
G1GttW+XKuZE+cbgxDfUyv0Ry4PjI05Rtwj4zp1Oy46thP9fJfBcqTVsUOn7tfx+
6DGmtrrGY070j0MlWtcMkknoBKAntie79sZwC5oaXqXeccNKRTso8SgLRvwbFjVV
vHzYRTYXNtFdKMPl1QFgb1T9K2dNYoD+OV8S6AxAEKYG7bvcEN1xnVd0iGAChOF8
1s9NHS4PLp0xqfGBcBIKUxd1ahE4zH018/xxWS/4Zh6zo0eUYEdvdN6aOJSHNE53
zYoAV5vVOgWqMdGuAGgALdm6JqawAouBDUeHhsnrpmOgQAXKSYB0cLXIEY/TLNjt
zWKT14eOLBN/pIYGFeMaAu5WJ477a4zS0qVvGQmMDcVWjUGtHsb1OtqcoAtFX1BG
1IVPHEnfBMky415xP8vrp9pTaj9qB9cfHf3z5TZbIhVCvpqKd1n/qKYZJNyYo4L4
OYhkAw510O4BgQ8QS0XCPQbllRqN7/SKeajA4Tn9xVsqSFeDEE9M3p/L0UgYDi4R
bzqzH3C1sBzZ67JDSdaFR/liw7kpQKiv4iL14xnu5O5D6DWwQQF2RO3NDxxLV3Vm
jSn+LQ7PK42/+/ZYpRysulcJLQWxCctfQ4Z+1GZ8/B182+xCIugZmqXzalQ++4ER
jeqekUp4gw4C6MTNC8yzG7wWbQEor/P/sPCA0DIVrCgePc4baNacA60ZOU9cmKFG
pXKsGL9Mc+6v/8vJNA9eAI8DrvLiGtzH0Yr0wzs7SYAfHbSSW01V1U0HL6YR83eP
nDgBgOijqpWpllWZ0fSZM0o19jKFfZ3U66l8Vglu5N0aNC03TLDYnp4dn8OgRUMS
3JlLGxRVPM8EmNXFDZT3e84e9b//EYqByxSiZITVSCuODQnOn/fwyr6Vt6xKiBPg
+YTisJOzNMwiUwmbGA92mG1fLVcEDO7WrFVS5zxKmy9S1ArgYgAof/viqJgrf+2A
dK59kG9yXUpyJT9x54D8VaTq1ou9yAW9prsGvwb+cZAzdiQYPZ42khZDUsRsnDS1
VBX2+XXP06gdba7phlVKVg4ceW2pKQwOTxjTfOf47PPQs52VfC/PkbVab9UId94O
7V06u1UmzVwRrif7k88TzMd/45OWZfzHGY4+j56PTRms4H0ygaRy23PZRp+dRHuU
+7WuvGofTIlxDyZqf5NT1xCrkwhJQCDbv8oOPvtaVQs1Hy9SPWUn5zDjyn95S8g1
uFMIM9kjncRsqs8waduwFdHzxLe7TozeaB5KiHaX2FPIinC/udvEj/jcVN/uF1dO
4UWHsJVxKziRQsKWK4lLdejIKoFqNpYQTdebCsszF8fOEGgDpfHjZD+4UXb0s+MA
XWfECDvurlDdBlOwj70mh0Wxx6Boym5cD7Ovv6k3ZwClgaN0t6rt6dphRWzjX/VZ
z7PEWKYVmt3t2Z1e6BSRpWYlaQ+ItM4WcQwTYxHXYwd0u68kGxFmPUqpEWbE9LKr
tuXGRumC9HIS4NGemz2Y+03JRbFcWUCOK2owb0TpBdWT1G8TbM/CFlJARmDk+iV8
67bH1xNgfyp1+URCATbPpbGx8QYc7Xd07lM0Q1Qf1LMMN5t7GKciNyoL8aEsrzkn
CdyXMLnRuH4CF6r8hxdA7wCnuWmsKO/Q7sdXDM0CIWFFWQ2PkXV6hJJDld7bDd4M
SFzvdn0fnRZBszGm2TbhzD93GcVoXE0EzTmfQPYboNfqP0hWti5pfsJ1OAHUXFOS
y/YxwUF0lluoid5ruzjcQTElYWXGkMLvJDJrXsXiblTveHjG4Kz4TyIQiORzocO/
/LeZhU4i2RhBJ8pRIRkJsUyPtdjamapxi3Ga3kU7pM4vOLrZNEaTxTPOkk6kLPxn
D2RAcBZ02TbtLsZYIFHwJUYPEZ6Xirkh9QkYU2eaMyPZEhEGZO59yW5RtboaOkPa
4JmxeC8ei3D4QS1hORI5cNrQRrd4dh5TcKBkXi0Gshi0v4avmqTKfR0AxxBs1HfB
8ixAKhNLZ2ND5eKzQ8tKuZEWqHQyrD9mUpVwZ7Yy/ID8WIsm8PjqHbF9aFQOQbTZ
l+GQMRDI3QkVjDdFIE7uHn3q4VQGpIYVBAqAmeHo7ZVNQJUxZjSH7vIJeB2rHE27
5u6MsogKligjvb//gFYG7ivHpdCU5KPEe7a8q+1Y14PFZ8+TRTDdxHOamP41J6/L
r8xeWeWfMzi3zzXsIujG9LBsE6giFoePRNeccTmojep7/MCIMSxa3siwPHjB7WQR
38Gg4Oq/WiS5xmgAEA2QR0smwcq3TZ+s6xjfwmVq317webQGXN6Qbi1lLWLgs616
Yg//oGDIArsJkEIbJvqsff8QV7GB/xUJ7te8vrCXfL9INTEUetvu6Y42VZbbRHi1
t0+/68kwVS9DPvm8iisvd/63/wivcJOqzCdQfkD3Ase5sy5Y7bbn/oaqQXQZufil
IuoMvK2DQCRrJYAbHHgP04Xa1JUis2xzNQyEolbvYo4gsUGDu+4oHtrtjDsMWgFx
9DbTBE14mT/JkQ14zL5LGq03v1z+2qyBS5ow9NODiaQQ3LVtAJLX+A7sQaGXFcOx
uWG9j3iPAyFn79NSQ/dWv6kbMOfWBbRAHF0z2/PmAnmuHtT1wVLRKNmEORtjHNFY
YBqyjgD4D3uMF4ssVvZVIPxXD239530Il/Qh24xyrLqAVRDvelR9PqQTZ+2B82+g
GTkKFwIwCODJSF/5rwuw12Yv/PWS6A22b78yUnkm6pY6uvHuzr9UHJfVh4Xbmv0B
xam3c5YA5aTLBhUe8UlZ5Xa1L1TKkX4eKPfwn5Yu73t4FddyrNXy2FRY2jis6I8k
QUFzA/qUAPjnig95s3qdkH3pkyq/GK3IRDw0R6Lz5lYUpUbS+47ugOOgxSmOt04b
CBRqhFmNmR619qJXwEbHa6tANZrhqFNGtOapgQAzwMEIEgsFqcoBPmhCEly+/Ant
2zF4Ab/lo5eXb3KcB39Wq/IfKyvE7SM+keEa84yqHUl0mq4OhanNxZ690Z9qjQ47
2X/TT9wu5FcbuLu2PLboov6etR+xGpSPXKhRBGmcXKY0mhNDyBZZiOVtQDajy/uM
ASTcKJsBLFTrPDylAQvclwZvRoonbtoU1hm/6JQiC4e6OJQ4yVQz/paiN+i2o4Sg
i5ntJsKLPDNvPP8RLnot4xyXvi7IZmb/aMywQKAqaI2jsMMHVcn4OQ1PNJM409VV
3sPnpCTk1rbLbm46Oq2IW33xnmKfMnnASpPv1jqKBkSvn52TMDceXlPPLtgdRMxx
wAJwKSr6WZT/v7oPQX7uiOluRLNcy83tTUpnk7FAWSFg+uxvcGvvc3lzsoBG8NxR
sjodanBcJICnDlE+wlsxHIxOdWxiSo+MRJ8awMBw9Sjdb/MPV9U8L6nwqapbSBk7
WtHMgKuVu0HedoH/LPw7zDlR97urUafAPOfmo/9A+npgVfWiPPZgamfMt3+FFzie
XOsr2rzWF/lZ/JBeMTTcXFFNbqWUBfOkSxfxdxUYuUH22at/NYV/DCnGNUi7woMR
yqeUS5JW6OPFy+blo5DnIxk/dkZ5Qx7IJkCZhU4TpA9r5BptU4H5gnV4AeAU9Gdi
xpjoCN+2pnj7wkseb6p2qy8O4i3nGEbl8oyrB96J4PbNvCVWGd9UnROto+u/GuXK
HLsdQVvMIs2Cz6hKDcHUN4TyocSIKezNGDmmnhcBWHnWe6jb3rM/i4L/8ht9Y6Rc
0N5d/HLSkfU5PZAz3lsjeOUMFSYulfAbECdSoE3XlA44EUuPHIT6ZDarI4Y+Tt2d
B2SC9XvhMQ9WxLWCytEmEAxUPAzCkJXFk3cQ6/NYE+3ki95YFxwMU5AFJrLYFJgt
sRFPBt/lPSLPzIjxFWtBtmEk8bdOJPjIc9uzZQZ9Xf2TIqIqBTStJXx5yql4AVyl
roXEp91HXPmzlkZCv9SaJB/ugYcxZ3gnbWgsvoRuMOAXAuGRZ0AUkF2dKS2sohfz
QeatbPZmzjrhSgtjnfy75FcDELJhe8yTgc9AHbQMZ/Q3yg0XphdlG2iJl10H3Cv1
gC+dNk7sdPv1wk20ZN+z4kqfQEMba2JgPtIVnMwwjx1DUMBSyh0Y1iw0iVbu2zmi
Sp37GCmbkfd1dFzMtgNy52+JvfEq2O5aNjd3eUypvNhr/vDyx822qwhOB8+4DQd1
/nq5uzGCKIdDluQgR+NtvbQio7+RW/vYYWJVeqXmDLK96hG8L5Obf9GjYfMtOGSa
l6LvqmkWMjdyrGJ+98UKEVtr30UnUhMWLMGt3qEXzaefKW2bksmYPskdhCWQAxX2
eqq4k9mq5Glvw0iI65TIEkblSkhDfDGcjOwKI7YWK505Vf/2pdtx9/s2PZBH0Apf
MxyH+Ty1RmNgOx/+x1b98PRfWBd+o3865euLFRJR/wEKGaLKHGTzA7UadK5PavAS
IZRsQCaGi/yd1dKaSXgTPzVpzVeOfdqgxpeyIncajsgNx0DVZZonKTnxnwKnHzIm
/0gONSIf4W3BsdwGBikiBimPiJirWHHPeHIirOMKDIk7cCuYJ6vv41FQT918oAhj
XcqYVkUf3sExxsFH3w09FPvR+3Warpi+Jpi1/m0kmPRYl6cQytbQAEd3UUj4C50p
beXcROd4aOJQNIt1RottQq3J8B6hfl2vl2wnatTM6DMi84tvBMYltDbWme+0y7YD
+9qMyBL4VEsnn7YXR7tsIaYTybYJhQtisvcDZ1EX+NQ/Iy4DA/WycoqBy33L8lVO
VtEA1Ml3CS/u1icNz2q3e0dJDZhpEOIbQF5FVM6Jo3cKCgPieiz5lg6RpahMF/h0
uPLf7lMLKgLBOUkl0GeX4K8md3UOqpCsnABSNUFP68MihVTbfZfM35BOb7zM/e/e
2JL6Ofa/Q8WxJYV1AHDsvOKsIRMmGcQaTDqf2IfR8jSwTJ8vrho0PKtYVuUmju3H
8TnaglWmf00yIu0B6bbFJ8hnO6AmcZtUyX/TjEQqY7beVI0hyFeLtY3M+7spqZ8C
M6mdfTZu9MC9euD7Z14Ru/7AZItlxrLEqO6rM9/ijZ+TBLY5TCo4HMdXezRn5S0i
HqXdhW1TBwVR8Xg92wnXGLZ4VKa+71M/6QO/2/9r1yh2Q4FDDLL+zQm6xK1hOUqf
GBzxzss1szpsR1ck3F+69Vrk17M0nUT3CUGV9v9Dd5/cUl74MOvX3ZSxYscqJlpP
s23xsi0zlDjtTjiwWJYwtcj521t/crMXhwwIQaVOXNkA7RrYWnD91hHCt89yvlTC
hzhK2CRiQDqpAIX/cJfVqczihITDFbJ6LotBOLGURTLbefipIY8TRf7Vr78rROMt
s581j36tZhdJi+ew3kx+QaT+Ywz6zVEZ91r9JaXNTT9erQQdr/gEUBB+tfmklnnp
yXofxxYJq7TArHn0jHIoUWLIgAPmEsDWTFktIV0wwGaB7zTgoVutdjQR8J7SzbhF
bzm+geWsNXSLjIhwLdiefNjg+s0o+egt/+A/JQ8TkRvoqA7a9tFmivx8Ue5TxRl4
vcN+Z6CtX676YbS8OSHAoVGtte90WcTXFu3VJ1QOdP3YOymeeBGLT+Qfid7DlYkC
Vw/+7jULWtIJHhYy9pTaqzHIQ7kpnHBE2E3hZPW9T8rFANUIApcynKdJEpCNsKo0
ceNrRiEGUlcH+I3Tcih29zvQPIIz4mOPFi6XieKLcnBdsJeN/Zo/+on9fWoHaPTB
KO3lV9b1kEfM0Fs5fythRHOTCe/xHnfBdXl2hmie6yK/Ymhvaom9aUPBoRMHK/Y1
MNzvy0famyFN9tj/XJLlCzP6T5huLunCqV/LeIUrzPJvZ6jEyFoesMLtjlcJc4Kq
5rKReg1f5NtFDrZclMdXsqIycEIDXyinRBYY4q798QX1180OeoXFgXhwUUuP6dcM
dkMyMItczATI+C1Os1p0zo8N+ag9JRu6yy/7USEraVCSbnEilFr/dFEWyPezESOb
RGinvBptNEYx3ym6a6q1JHQp3Qre2N486XL40a6Mcxy4X2yfmRVuGUilS+zD3s55
JcEGF7Bg61PX7RyBFV/nvLqxI3mYknVva0AqsZ7s3whZ5gxJUZkVHhwsqr7IJpmX
TQZsS0T+KuI3oePJUN8oenCLsm8QFHd1SOQ81iL61NkFOJaliii1nuhIlA4hhDkU
NX0953Bc9MOWz0WK7n2N4LKaran1BML1lT7Z91/Yxb0Nc0wBnA3MSle3agIscUYY
ssrEUjptgoG+W/I3BSZaD48QFI6ZVwswlwZdfeFrKn6X7eYsbJbyq1kx43DdNe6/
+UZfQsjJuwviYXI9SpqHn0uqitA9xMqN3DDWMKYPjVVSt3VGIybEilM5sve2u+21
kN1u0hAhDfDmcUSVKzJ4Wtf1kTT8QVSighh7e7gRFXbijhkgGlOedxFi+IePEt+m
ohOkKQvOR0ug4f0eimcX9Dm3g4EFlDBPXJUqdhmldPi82wLO6IOcsaXeBG9GXUxc
Yhkq+34wA15urj0WYmRBAASOSzDbyvGG/dK9g6DhDKMdG0Rv0p0KJoFmRGeJVdN3
YPc49KiVF7mc7+7jn2G9u1yutYDJZo3JlSUBxsGtOTvPEeMgYHDowUiAZBQr/DaU
p46ZKm9cwJa6RLjmi0KtJTSavLwjvUr3Pg6Q+2f2XymIeC3MJUwNICxOiw2u1n2U
lp6nerlpSpiFDtadf2eQaV2fV+K7XhECU/bm1e+hAh79aN8Dm/ll3LB3XancDC4D
58LINjptlyyIbfzfN3AeWMb17ImSvWpr20qhZZ8/RQWDrF3LF+mXibkZHSHcQXq8
B54fsUCRoFdJwcyk09Ebm6oiJtJ2dpmFyxaeGW5busDufBzHIdeRjKNkhRYLrBeF
5IRUQ207grizJzCUGmwMIz6vx6DRCauLe6ZN7AOe4OR6zfcax2qNhxKrtWW9ns8k
Xb5euD1bL6Ko/lrUX5jPHreDyv7FLoJHDRI7iIA+MpNrGyh7LokLQ+54A1BPtt9n
od8S8udK7azE7uNBYUFDAGx3wyjoj4JFzO7FtPD0XgSOU/yDFNBurt4ZBt2PLgRN
Oc2j8RkMSoG7B+CxfJJkI5SNla7w78J4geDs5HfFEHjVeZjMNk8ZaANd3o78zaL7
XCE3tqetai4dGbm3jjeBQv4SwrcbPVMIPgtpkyqn4RIl51jRdJLjKXbvWz8xGdRs
fm+vQKkvrCke1dtJ+CiDnd4+/mRrDlLztExRpfPRnHbNsPPZWhvpJ4//8AkfVdnG
nNJjyGBfPiuQrzZOnq2Reh/BtI29/RIClg6Cv86LMUqLW2mgfexdWVpMPrMv0Ldm
1PSxGY3fOwn9YNxGfLLqZA3+PZTsOXVkgDX8GY9VWH5mih8xiMZML6u0sWslz70+
dyvMSCElqH4qFlWsun24+OflvI4+E8uNT7Cv+PAXjBLw6VEOMt3H1eEkWWe16QSX
G+zIHUmAjUebUGo1AMHubpEhejLnMjozMOBPY17jnI/v/8R2Vt+fkdeORuyr3bUZ
IViDnDsJXIugNZMYybynx4SGuASKNFp+8/hn1vpWawtvMgfQIJ3v++1SeG5Physl
qVTVxlFFmwTxE989FITp/5VsJK/F5hLUBUWZkmii/5ffZicqqemVhoFQcL47fSjQ
z/OZJX58x4gkXonDJx58X8A5Dt7WwtvXsCSgFplJkOv1ZXpNDeFnO2GyitLwYms9
CXb738KLI6n0iMauU/heEQHDmRHKNP5BBe/0uNld3APB0NoJASpZ4MTPgXwIx4QO
WhadxjcSVL5y8IYNUXhpdCMqupeiP9fVBRN+/rsnuvlMv7Y0K9p60qJKfGYf4a4a
D7VczgyawSStBjV3kwATRV6oyJ4RNbF1iViZ+CUikoepeB/i+kxQx8wwmFau74zY
E5qX/mfDL4bJR8xM2vRjYOHzchCS3FRyYuaSinUbYRRaWyLmfHLvJWMmso4nVZQR
2jI+iM/8gn9RYFTLfcNeTozIUk6uYYwSzZzuPyu2gLwqCAi6+Z5qQRkDmT/tVjyC
loLE/W9a+M7XgQua7KFTHwdx/Fhec3NXM12Aov83wcSrscvrYh/62F2G479xSOYI
+Xh3CIyqnkeCatP36uvSwkiIrx9uzSs/MvXu3dbBjcCABbSTd35iK/pmKIxLQUy6
4z5NJ5OnNSlqGsCLhv98WcjBt5ur+kNl/xiV5tppHejLFBlXTXtIWOr2itR59Zzd
DAvYKrKz9Qd2aWvug9/DZ4V2bxw0ym6ZBIIxa6z0fw8u3hMRywdb7bM5j8l9Rw4V
HOLPqzFVYS4QhGSUJxg1AYyopiijf3po+AOlKI6RoaebzPYcjtyRfwGjJU0yJtvf
fZ9dDAa7E6vjwAH7Uqsm3Wrfz2WpHfn4k8kIZZLlPrHPaCcQDt4yZH56Cyx9gEnX
hFeduir4M1h8HQSr7W7nvVeTP2fStrXRXDqtvUg/D4WV3yolYXXEhqKgM9xAdfMN
bUZjKNM/+585D8I1QW3bV4pTa9Yoe6CDYtfBTnR4UxDWAZok+7ulvTYOjWsPLYsQ
9tATmcou/qKxEugo2P4K15BWF2JeG9NXtYIvJg1KbK04C69e3A5IzIgwE80mJjSr
pCdi3voHN5jZA0dkvBfd57hBmirmozoRVs51yBT6Sozmr25WRUdZES0qM8c6HVFr
nUeszgz18TqBEi8DgijesYi2tv/zvZnAr7+2o5lSqE07stf+CiMn0kOhrfGasv5x
iZ/UrBWY+YZnBc56WSgUHD418WtIp8kQQORKmjNEthkbtIMhPza48W8GDj3nfPdz
IsZ+IUHeZI3+/R7zhslSVyY+OeuZJGZfIrVoF+RecYtjukzs53tKCY+Ttgx56vq/
HBO8EaorgWLXxugqpsErJowChgdH+/v02tTmx8+d10Zo6+Ex/ky+xUynWnbuaRIz
ILdNYV+SdRw7O4Tn/0LlY9wmid81rDpkIKew/xphCQTqTtRBZn4OLdkm/WunoSJh
BeIZUyiq9AeSNnri/ZwX96uoFWXpElfXy2AGojLALxNPmSyvVX1T7lOBN4cngzRR
1yLvAB1Z1WmsQDShjmNEn3aMIlzMU4RmobQz/a0T/3GhMfMir0dcVd+bkYAZmRbb
gqabjQyWsYsnf8y8csm1DjSxcwb/s/3B+ZoyU04coJQhGPvx8+GxS/q8aTiZZYBX
8sm2EUW90HvZe6l/BC5cJniDUWBbYrEZzQzPvLCAZKkqAOnOdSHOczbCBjAAWVc1
ocAJfNhxd74GAsZowdx9UdOASh0+NqhUetcp/KIb5AVcXhxoRZENG3UhU8dtTyzW
y8JghwwFkXrf8zxH6HpNJrbGhXnk9lYcV1z6LuRIPHpYEr6f9h6xggouOqQhUEoH
AwLXTjIgGsXTNtL1B+7jSlfqTVFlwpxHC5D4fRtGSoPDX8PCCp63c1wYQLx6SIb/
84qJyCa8+h62aiW2bH8D+BsZiDGROryArttqyehyhaL6hrije29+EoiXT/k81yOM
HXGeXVHGLxm+fc+54FaKzJesMjAMJJ9bnsvv3VIZzuQcydPL8K8DSbznV3W6Vdj1
mE+or2o+nLQL9eh+M9YNazpaXBpGPxigkaZ1zrI2qV6OoiZzzPeKRmBCWutHPlOa
yLy1ALv4UVZP6FIQ9pqNrOmAFyoQQRUQUcft9kynZw9PBckuHdbXFhYhKYEk9anr
SN/BiySoAqdBJtsrUH9chzi8oA+k5r8G27Z3llr7gC5gSYjYCrK7DIFqsPp5fk0O
Vw8jQSFpebKZ03feJiK/aoy9bohFiSpxgZgjV0/9k2zELCRPSgPOT8CEBkByylys
AfRudBSJwE67bwysr7EgUrRJoWG6Kdz+zKuiABUzYRDbUU0y0K3blyerDkyV8KyN
KwYP4PodaiZMjSI84d40a4ABNNxMOqCHP7NIEqhueyUiHz0Y6SKz8g/r/Dje7ozb
cd3skJX03G86NrJLwvZY5oppCOKltUztfRxNtdMzq+wCXnvMJ1Mw8A7c7XfZhzB0
MBtJHXj5WsE+Gam7XwhAz6ChKYV6voDb9RIMLZ/f+BknJDOIJBcRsBFJdH54x0Pa
cLLIOvtAbWtN2u8uDj2+gAfuIcQ7aDODfr/xhc+gDGSO2//8e44OryBGbjGXZG6Z
N6kg85CEIvpGToHh79PK6a3ZiTDBnMz6aKjm4JqwYMcykv7I7JlH4LK38kAKEege
VehKgJoH3dYil2lmBUKs+kAuBglgLFXSHKUNghMsRS/TVWQu4DivxkCgPbsFsIlc
s4lHU28AwaQVCP+qePFDUynxUZyAIJ6dkZR5fxvZq41C+U/vv/hlRFb5Wvlvljk/
yJD3f5RtHDYTsEOCBl9oRTwDaG/GPMBy7aPIZe/g0SQAn5rEXoyMgTB2z5lnkkI8
1syk+NvrvadFZsnfL0cDxUu6QuyVm2CQ+1+xuf6jrlTW6p0rZaslq7JXIUaaaSFw
rA/mcXTSqUBfxzU7TdIkINT6GzBz6IAJbCJqkpiZ5ClskoyNH0sjmSaU1W0jIb4x
v8Q7AS126MgHCgvZu4vGPZ/wRM2QFaCyWVzJ2dd3ze2RwtdP4Ygp+uMO3RKykg75
dDs0VjWV/6QxHtBi6tnezuoWQiPg0XK2onvrSbmC6p4AaXBJzqg0iGn+smxIevmG
kWoPw51Vxg+JPmkn6XabA4fgQKYA91mOwgWyQf+UF4cGOqosspjO+JaTADfmbazM
0qmD0DMpAokn5V/j7X+8f6z7O/RkxeIiPfRQiRL5YaIIo3NqTKpCGbTx0DmPBdXD
mLBZdg6ihmVGgTmShggCPNY0llbtTLJ8Un7AdzvhUKnJeCwZz3hlREZmjHlrLVAS
oqVTuhORT8cqh8FAQioQNB7gYhD1MVwmK+9Fb3Uu+euoYiwqzO6siwv9M5bp3hsK
MUN1FhFnuRKyVXs4czT2U+QZKYbwMMh8Rml2Ay7CCJtyE1xWtKDilu7x0YeOYi0i
3BV79QJxxcl1hY1g8MTip9UybD1s72CTOYWxYJPNwWM7jvSOGM2v8mzhYP37pCO5
OQzRCVEQCWAcGCI3eu+dRYBkKEvEkEr4v2VNtLHEk+/0QTU0NkCWjJqBEpYONEdC
wdFH2S7f02abXALHix/++cLqPNGsbmcAOQ0+AR95nkjtYjfdQsgFRLquiPuRMqXR
LugvSBsynpLTwyKIdjJm1a5HPx2eIq91EVLwW95402PjFZzBJseesz4eOp6NHvZX
bJP3szfrYW+Ds4TzZlk6VASmnbom05OyaLRy00F4plSTSsJLKmQ7Rwtaqvgi3dpq
m4cIaYsy6JoFvfUOQgof+mZaKh7vZSURXiZ9a9b2BGAUcsCARuTrIl9gHKEpo7lx
s2F1za4PL/GwoTBSzU6uIzhIAnaFqMHLnI0s+2YvnMtUHmi5pu/P2HvWFNdVNWwg
uYyu9A2Bh631w73gQAen0rbaTBLIZLakmBfDPF7wLq8hYF/8pYq1e7XBU/Ton0NE
cGeJ0S1IdVFN8pFZN2e3LECqObT+seg6K9bRlwZMKyXoj8pbvoz6qFywyZXT5TYz
ZSA/fVliCuu11l3mgr3GDk6ulQFMPxJv5s52oPgWZ5XdAPrXwN4ts1j8jiGgcOQy
FyaUS4dEsTYt0PjgODtdrC0hiCV9AelznLaLYfSUc3CvwGcw180Q4sStlZX8Xd1q
5kxp+Nzs4AlQjny5kdJXxpGD0plE3jAewxpE19trWJbug1VS2Hqn8s5nG/tw4EU+
zAilZcZGllfbjvspsdPTlhNpbB2/HUvq7AGRvtVyxBY6sN0YBRdda+wJFMIkjbiM
dH9tJY3mkfQdNN+R9F1BnkI4aYm9QGCuX8TpI7sDSgcLqOMwZ5unvnhlQciXljMY
UAFfPU1mfV5J5r3tHrhlEvRctyMOCG/LM7eaQy5u4wsnRbKs3hAtV6GXh4V7HSIT
e06VxVnV5r/2CQzRnVUiIPWMsIG/GrXqzOS22XCXUiaTcVjkZVmACAl9hl/06WE6
44y+XBcoV/8ApN6SM3qM/eVZpHMMQ7oco/o8/Sj1TBgxnclHLj4NrNZdSfIBGNNf
v0gmy6DHZORPNhf10d4M93gREGGPMCICHXw1RxmuZhObEgE6Jj7OdliU0g1VP3VA
Skz2kRqf2Vkqn6lZiSpXx/mTdOdjuJebhuPe8Yz36CiNL3RDzVhTqOeqxUKmLUnh
OeQxtnIY0JIZaJmJ/Ci+8TjbVCqh5aymoUspIPePv8B/RXq8ak7dccCW0q3OOp6g
oou9daf3YPZYkxRhslErTGkw7ZMbsKrC5EMM9Ru+0v3kBjTRLxCM5TBd6DWkm4GI
7n4RBI8PnIrPKaeStnzyfyyhmrn29U44ZjMQn4Xz2X05xWWgBq5DC280Ck9rvu/M
3PkzcHXSK1Fzr34il5xPiIuy20UrZzYzYswyBKxBxmftm4U7jqfb1ujTb6ATq5fw
/nIQ8ky2qto7u/tMQJAWIKmsT87JS0xaayqvN1OxuteusxlmiwDVb+yrCS775qab
RA4jcIIFJsSemj5k9OB9VXzeP58s7UgnbsUAD7O0ToKFD2FOPXIaDJaNhezSGGns
TBySDXDyGIuuGTYnawB4qovZkE2khWaojq9aEIU7auKUGtG+ZRkhLgDnOQ/2sR1G
T97cqq3V6/Dra43fgVha0mTSID99AbU3tYzZsqlfixCGJv/sKUDu0EbptqfbiC2y
esQIohaLc21NLzCcpq3CxdJ/Ag1R04DHjne8EFgc6JtXY4SQnI6PJZC012CWNvvJ
rZ+w4wNTnYcpfFT7CW9x6FQPjl/w6DmGI1gP/4Sddz5B0ro19pVOZXsZvdvuklFP
7o06fgj5TwMrodVHtmkC0t7q9heCxjJXZnHEJUlcsdsuXtX7PGcRXzYWbv2bXNex
miFIZouxhz6zM4Pxu6BawOdaXalCRLKdH3dUwMEoWi1uXmbpd3lzH5RpR/UzJ8IS
rfwf4BW83HFGeMl6dhE8J95Bdd+GHPto/AiHtcU0r9QlnE6mfeCe5bwUVNrPPCc4
QWYbXlr7BD+QtFpaKPySkk5VJBqxpCmI2TvH0LbHxYlGGEVTQvitfdpKLoD8fT+V
VBvMCTWRlwrh/LVqYqV7VynWuXrRR2brgm3fBlJ59tsbWfWasItlryeyyUoanhVY
ebtuIA+GYlVCVlxDqJzkEK0rpI/DulLH2dOxa/5Py7ZAD5STA+6nKfmi2sJPHLMT
vxonsnwsg0BtuMkDtXafnKVLmzr0XD6/tRdfenUafCQL7vYnEvuK8iUfQo2eGqCH
2ThvFRt+trokPfv/AsqGhDBmArLdKkiyAsvV6wm3jTJ550G4YWbM+n+k+58PRRoS
y/xeNdTXkd5YE5BLYyck7Ndcfu0CcZKH+48hoEBVPQVUQFh9fMlWO6WsTzTXnV31
DwwVhu17m2M/6fgtRS9F6KiL+vpwz+Kms6DjR43CCgCwMuabppzqlaOE2E8w+3Rq
iXpKVLnuJQy04ODup+6kUAwh/tmVN0H4OOJiR1cXmP+LFaRwbs2KJb2tiWz/WNh3
jk+DP6set+QruKnVUVIY353oRxs9ButF2aTZTh1767x5nIjFKCBhRvV90A4YgrQL
32nYMzCkx5UQI3ULOi/pbYCh0U9g8f2ELOX0dMlbkX+ddxevO3e4Hi23JvXHMNZQ
KhGCVuR+QnzUSFVVX2xZUHUUIrsLWVTMROitCsNXko+QlCIHCpjDkEBvwVUdSWA9
2DO3F1UjkO9KFt8u5rtB4EnskBcJrjQujNlyF6YJkRbBEJBLQHxZ6RHFEvQ6Xqji
88YFKHdwdr/pmVoZOjBOoc+vlvklnnpchIq5xUHt8+MK1cCaCscflD2jbITUe8xR
7J3z/pvKpL4uUMQiBR8W6qqBPuZH63qPz+hHzrK+cFkkeIznJXjOuq2M1pVmEwA2
QaOlF9psUd2qqmG5b1LWh8mYU09KxhSpWhLx5u0M0UcA91cqDnSjaaLAJ2y7ZstJ
Z2M0sdJrSyFT5uxREQylzOc/KoFgq1z2k1bOfSeYvko5gJD3yioSQJ7IVSj46zKT
Hm1ER7eSmMvlK909F1yGMfBhnr+GJjYdD0hY3wEWeAC4t/gVw9Sja0DUxvVRJYM+
Nqr5tKS23+bJJqq+CuArMDYZtp9aUDpBIiNlm4GoJVPWgYY0s70VS8O/201dYfpz
NXzqlPN1uiTLOgcEtmuAJHXrF7JaZYWw9Jn5BvUM3808fEiqexJcB9ApfvxCpIj8
hu6ck0AyrdNPL5r4s2zU6w72mfy6/xz6QciCBrVZvLv9Zi8SuG7Qj9pHXx9T3KyN
YpKWmeHNcj2qXHLUiIKJobUFLAB4AU0flK3M1U0voYUr9bCZiYJs5sl4FqRXwge2
4mrRfPoGa9m+1LGO/PE0jAT0ZAIa0WvDREf3THZHjp+C8MqHYc7UQBSv1Ud916p/
ly8mv+Vo9NQX+xur8UMu7oIMqutQst97Gu1cKc6Ue9UHTqoLdbfJyzHWXJv9oMOo
LccVeY/TD76TnmDmvkrhkyknEfYHBRYqFWGhHuyIceGfS97ANSOhUNPIS4Bn4UTA
ejfhGggjISaZBLqMuY6rmRf0Z+onTKATdYx6WLJL72JfjOUWu5g7n9Wor7bmJntR
4q7uerKX37Fl202MsYDJ0nkOs1ute/fGL633BGW4rKLoN12RshE0V3PahhX4xsM0
r3V6sYx8xfQl83vW9CqXPCA5AOXSMTubzY869/KiFjEnv7ARylSGdi5Smdx4gD5H
pvxWEiLhG/GhVIspW3A16pC3KvyW+WiYYlSoBiRNenhPLB8CHsjk8AZEelyYOfUj
X5pCMafRTLenrjwEFgmbmViWnuik4nLpqcYTyURuYsDfanbckI0OXqPvsLCjDKEt
A427/de+v1wQD4MJuQ1uIdMmZUxVRgzxpSJ6wVfypKIUhI6v9L7tyl6Fq3ubtkKM
`protect end_protected