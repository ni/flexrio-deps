`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8496 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
akBpHK9XojjdOyFTP3pOwlqmu3HKDkgfdD3J9PBzA3qUTDSliiCK3zqdqHnugvSY
5CvKY1uuALAKlwMntI1Z+C4ukHICaodlLRUQFrC1F5/eUksIuMMeKhLL0Dx9XMwj
nA4IFaqhsU2WmC2G0zzSycIYazVUpp1mwoxBQDXOj+WfB/5P1hLClvhIHABDVGw0
gC0vbY+SHswmqweb2Ffn5UaM5vSmAUGeoR00mZ+DQNx5kWWDluyw8O6fYoMsy4dF
AufVRrR0gp9TjmbNkEEecSlHsYpc63Ten2tWjAnhTprcDtb0v78wuR8JqkaC3YPk
sht5FBoXdxwP7FYvwkexwX8g763RlmdqnyRE5NMt8mF+MXjzgoE4YcXiqEM9+1fB
QgEPkyZsR4sFqflg9PTZg3ys1KxCgLl+ZQTRdNxMInuSZPLefwIXT7vlc3VvI7v0
eOHsVp6QRDV6j6XRf31DTVis52/lxySS9bdGCgXOWxVe8wrdRb7nlP29BlJ/Y4o0
4uLkZbJewueWGK2e94jQPAD57cTLwXwF439Qru4S9A5/U42jp3u8Y/LH+aGbPQ+i
WQZKp8xVEPa5lcyN8gRYscrW6nFBi0tXmg2Ff1osDF7l8uxUueMfOL0GrVaUZd1l
5AkcDmDk+91c4JtjFjCKtFScyYVRv8AgtelsqrcyWQjIaVnTVtsZbHljXmus3S0P
wFSuBe2c0cvZJuUdTkd1Mb00zpAAHkLuGALtmOIrRby2CfuNxjbVrWpdgAcxq93A
XTI3/YXiTNEvEUORFYMw6ROxx/auvUaSEk6lS2KJRA6rtuJmUwOHPkjJV6g0mpjp
xdfe3kM927Tzvh0pG9eiexV+rNHiecMtkuHipIYouczTws697DenjxwLAvMOo+Qz
dveYhTvUivtUXB9jENVSF2sY0ZYbBoSkHmAiYlzg0k1SzzzMdHz3azl/fKTeDxgE
DqTqCzNMpWH04khNdqLC6flqKl7gqBSeXc8W14KZ+XngjaZBiXoD+0AmOMeu7Mvm
CzwYs3CqXMkpS2lCT1rF3yVp4MtZwzt83FM9vr/O2k8l3nBMHxTdUDnS4Q/kLMH9
5CEUyTH/svn9Uwq06niEZ1w/BQGgqsArRaqeWinOIHd44h1+vTZdB3yx8q8BbW7b
7TzOONDCrQlLpZZUWtlKg5Fv9OWeL12IfyVFSv+3njVBTFox3H+6Q+TVublEC/4d
YitGgDPjXpZd8thIPO7ggT1yKsXJy24n5evHO6zTSatpXYRqLKHNYI6rUpQBYfdP
EryrVehk0T8A356FfHknv7brO8AssJKjxdWk72YvTmFfSKyXA0bt8RRcJ1elXkZW
nrrsitvMuW50Y102mczBE3FOvtsVQd+O04HmepikbcPA7GIW9x0C8u9Ke//uX6IG
OOHuvlWEUToPIrLn4YHNhLy0zxnb5f0hZt2acMHt0jMPdOhK1H2eVGNw6icQtj3+
fQgy6CT8tu0nPTOk9qWPi/e917Nl6kFnFcHCC+aPeMVMhZwQti2/LTdZDoGX9wXM
AhJ/A7uVFjY7GJVo9KOUkO8xT8+3EuTUJBDGNtsruju3SXSuZ1r4OOGiToHAkn9T
3O67OBxKarlgTc3VbXbtkO7f/OM8JBP+USrsm08oDJgktULk5NLm85E5FwS6qRiy
ES/qw7qU8wxJnZ4gEIQ8Xd3C4tZhm3aPF3EcoAOA1jFtDJ26i0zozLhwlaQk2rtn
JuOd4VMYUxxUuoBipW8OeKQv6RoHG+Qet5GQPlfE2b4ubOVoHdRTSC6K+93qSCM0
F4V7B2vzEaIhNiSgUhBUl2NjyW5wKuMcVLSqzu0uAP9hSDY5g+9HpPSI4mVB5m6T
mS4PmSB4mYJVQr8UO+/sfkS4e3wkW/t+55lfF/Fhbmxgdi8zA5RsETBGXAHvEvZK
sQAcJEj7sT9Nm1wl0pBt9f0pjfmus+oVQkopS18J+IZ1ySCOLpny64aVdQ4Ao/Wd
Wx6zkKpH3+bPO+KCZCOdk53j3mFAJ2FJnfA29CIWyygSUgy0BRTk/XCNdifYigIt
wFE/CaQGBG7MeQSpkK6GraoXJ/AuriJfxh64mrJ9lXS6n4GzpiTXHvmrmAapbi6/
eIx1n0WHw2uBjbOjvc1w1X/xh+Ersv+0lgAM10Fb+xJUAuNo0wseFufD5QaK3w+A
Kppl/G+rHK8cz60XVVYS6vNLnvqqktQpptHTq8LH+mHPxp33sJWuzRKyMff3cQbA
7VBxR2Bq2uNmJUw9cdjIdIpUNYK4oIiR1SkYslAQwCUrmmnNsafxAV9WkhKedNpe
Gzv3rYLGESQXsVROgldqbhXn4TsCRcTLqxpS6cHgwaxtIrXiyCQWAMsFjIMNwHW/
El+fc2YoO8slCvzVATfn6H8jjMy7QTIJw+QXu5dOKko93hnesAi4ZWgHjb4G1dqt
hMJ880v4wRIOEhLsZe9QNVYvw83LvajP0moUD6n5AATJ23EbdMWMK1RdzUvqlBN1
0NfoEESg/k8ISVA+tldOQoXRT9ibDGRxwc3NpSoUPOf8nAULc1+83USnlh+qa48K
AuwdkZI2lLwYf06gMofRK5finteBg4PhomJqyv7SDwQdPE+ry52x2AWIj2poNK+x
0uA/FNagBBHVJ5rDHxmRzxjBGe7vpVh3Wt63AKU0RZm16eRkYUIMpCzcc9knUUa/
hwHKRsVaJj5b6r85Vw71ODHnCUal57fZSHVhEGA5utksrBdDv2rCFXmOnLzHhP6B
4PXKB5owcVb15Wo0AOK4ZJnLBoAGxWwkniEO89/w/VkQIJ/ah4Jns5FucnoaBA5x
/7qGSub42yH7a9VUnb10tksiVqZ55CD4IC5eXlPS+9g40HFw1xKnY45YhpZIDTzu
Vj6LFu+otfm8GC3Llh4DyuQ8hFRXmp83GHlftj3hi/fDVvrONLCg2mHNBht6m9yy
q+mPw5TorRUDLbmsNc15MTn5eh7R47rEpFEHgQD6SRuAEup/z00977KiGwdGMSDa
F4727vNXQo22aOSqAn9ALCuuM9gocPJoVosQjfHeYo1LEYRPnQmW3f+hsnzrJPA2
4M0atnjR94CofOB2f+AvsJCtGiHlxDg7jNmmSN+mEXf4Ohoo2mxhuUPHuxYs/AcN
xuDINlhuxWiD+Aw6PdpQcHhuIT1qTA1nJByaXqhF1Gx9RqfupEXZgVkQ+obVZcip
n5io60TR0oEEH6ep21yIDrBDD7J9tEL0kqFdCcN5euLzIsHJTqCh880+r56IFaqM
ApvZjZQga8DgIi8dXpehf2Sfx2uI/K7VrMPeygUHnJxhmzZ2XuD82bkbujpXrCto
qOI2fyIFaEdcQzf7xgzrBGWYP896If7ivYZ6AHB98KjDr5jTB4nEMaaMCqccfzhb
Ajd/KGH0s6ko+g5o1qPEEE1XR4uQEIU8juchKbwR2KNy//7eMiSIC9KTYePfbh36
8pWhE6BsBfjlJS9awr42Jkhg1aMEeies2lCkKX6DCJ2A2Ld+dT6U4NtymL1Aismz
JRDylV842TCnnk0qoDk4yM6Ma9rgO8BFScJVKMd1rVnDy7cFLfaS6iuwoZUqVTA3
eSR6G0OT28efhm2CXb2lSv+NHJX9jIssUj4+VyPX0fCimrQULFKc4Vrmurc7NqQO
Tvb6peokxefRN220YzRtFH1Yuonr2HqmWYZGuRC2Zvtp6LBOa883M9OepmMnxNMh
3V+sgJ4juSm6GlY95p1B8vAcfKuv17Cl82OznOLCClD4aEeHZhWaNv1fiQ6lHp4P
K6Ua/0Iw+qpUcYoSMYXtGBgZG1y0akOe4buIYc2hTjfCHUufYZH/i2T8tS+Bnni8
8Chb1qUEUHnLVHPzTU+Ha99AtbINntrhwdCXVfxc/H4gtif9hpchmulQXv0V0+TP
HJvn3WdECvmQqzn9lGWx7nGY1mrO/K7CiO7uqNBw+VUMdVlEOkha1bHtgH2U8tyz
GpPqgCeG6pmUFdnbRcVgHRPlbc5ftbCx6NjRrNllrKIQaN+tNmIuEXiZS+v6U9da
RRqbS8BU8u5LUjs82UXsBNvfWzCwf71ufiCMUxgm24odaZFPwjBz8WHEFGmj0Jol
Whz2H1IMy9uWQPdOTo/8fI1nOpl0SORKsPY5YtVHccUQXtP6jMkCGhC384sRoBtB
l+5UiVGrJQSV5mcAWFRUOwcUK1RHEAnTWi41l8GXzdZQGtqfPgQhOeoOumHxfK/g
YHEEolwlhMkBU9bez4qcdAHSU9HBKIC2nCpP0nD0r3y2dnMXH3eRL6hlxMuRmmfh
TXP1u7iEQRAYRsyNdgOBIK8FszH+MbAawzA5tjXovLJARQl8WkhXT6CMDB0i0/dJ
k02RphqvxoEtJQYLdcIg9eKBNqw2qfbZHhYcfCdzB7KpGvbf0Lp2svHE5nbKgpXq
j4e92REosKih4Yer9VfTV83AGu81kP3vYXnmLCXUSEWWSlvk+ks/RijGX8j2YFo0
Gi0DlS6G0UxvRYwe96jYEuGRyJhMj+dlAlJt3UKLf8TX99zblKHM77ogYU57GJOW
Y2JPurv1neJKyJpqqV78voUbyXzKHd3s04IDp73a2jx+uOuwq4Sc/OhJ0FYE0l1C
d8BvjLzEAG8kxQV8ymPOBRfgZ44T9nuCOWFu7VKOWvASJdL5f8TQykfkjegfyces
zCegZQdmbePug01LZWjQ5kK1v6LfFtIKA4bIEBV/djU+5fDvPOLpjbNPvlPTRxso
PGYlleTACfTBYJQLf6Uf9PXnWtS/aNb6cQNallBbdB7+eAr0Dy8DtjD0244JIRyq
XDPf7pEi30YBWvHw4LUnkNeDzr9+Mpr89yIPPXGrHBu+JQZ7oHCFlNun7o0rd68j
sI0KihyaT/zgm0rC2uIWC7fQN9jYIc17FoBJ1wYIC6oKLxtWbaXgIuaWLFcNmIvD
jlHbVwDcyMNaSJhWPbKqOiosZWYYwGA+2ZzVNUXbqV74Ql2KRRGnGvwaY8L6zmaG
Lc2/EyhaTksscxZbtO4a44kue4TYfqVCRjpem9k3yI5AC35ry/MqjrFaV82lRGi/
a9J/R6uFSVdavk4rjuif1IvTCd+LSnmqxBFJ7WQj/zjJerJLlzT6kIT1rCa2J7wm
chQDpvR1Q3D3dDP0Lewk9Lih2Ps9HTSvYXET2bEv2QKY9KTU+SPXoE+TVYV+gs3+
D1JSumMkYsR7AYP9vl1d1V3V+ZbSUczEh929V/z1GmupMhh10BRVyHaR20OyBDsz
38V0jLCvFeFYjqNVHe1QMVhHzN9z0Y38gnRWl8mbd+mP82uG4Rbp2oQnllGJdhNL
p8b4NRL85QY1vc45nFNWZuZfw7T+cujUHP9ulxc3trF9MIFnzOMqidOxiB4PqBSe
lJYWcLMPAeksea5cX9Ad0LqV//3iqUMuicbAVAOAbghj/57TUL5ECWB1L3olcsPJ
Vq4pt1xSwDV1d+03I4GW3zOvO00RTm+kOY42Lpx29JSPuLfL+L0tKYNA8VA0Pv10
UfsApE3mwDiJfAeo1HAV/+3YjhqWLkMmQ60B5ezcU2nm3nvR3KBXpQDqz/05HAMY
6YjvNUGDXAwe1lf7h1gUkvhkamGkPzTeTYZxuXJBnFHbK5ejPsVDPlvdhxjrnKpw
Z2WEP0zjfibsQavfUCCRJRTtGZug8GucN88ZTvKd8roTr1+4ZGWA+Vfy7uXl9NBn
LM690f4pk19RJ7hCYk1vrpSDB9tZAbIclPQbGlfT58ciclnBA7NLvZI3UdTAIu6a
KKNwXaSxxZFH8rQKcxy9fzk/RX6+r94xM0Cxl+WEDZwToqkFv7qOCUJMSni+x6rE
9eCz3D7hrGNoiE3qYkWHSOwoINzWEWt8iGzPfilOgvGpnBlDIP6kjUugsf5VmQz3
snhrNaHtSVJJo9K6A8Prfi1B0zPqpGV0HIzsSql84K/wfK96ba+VrMs/78tcJfB5
CuHECECe4x8elGP4syZvdZBtBkTSL4pskBQLTigbztKETAQzcuSDqMX6BI3q6Tor
Ouhpu+e9YRsp8HBEwVQwOw1IaV6teEDO1wlW/e8otU+7YoyGcTNaeWwjDfXA0fY4
KWE/Q9z47O27MEcVtnyrYz8HrCyYqSv6Cnxga3sIQRd86B7Nk3miuobK/P+2gpA7
yFKZu9xBplNPHShYhyTfhTh1U/wo1ZkYsUVJTZzvyJm/clTOhnNvJU+yHvu9mPYO
xjRzXHLP0TBSKsK0Ty38iuk90nDVV6QoAe6HGZedLGgeSeRiK6jQVkclHUepkInH
ZSflXfNfTJOnmnYrlwYMXPEwpOhPSHk2eSpb0mnlbB4fj54CpFTgl9s9dXwZVcs+
/rPMdpNludyYagTcPDmNrokrLg6q8ZX9S5BdiUU7BcsxKG4LIP9Psozh5VXxRR4M
f/YP2o9n0El7X1pv6i4MSFURzHsbl+V/0f/TyI0H296xfY6wJAPA8abAEpnQ+9sl
K5iWDzPEZzvyFIqbq+yctMudsCwqUbMkINPgfw6ZAuYE+muwQpxZC597XDt/yLDx
+nZjoPuNGY0VDeZGPqAIswaNJ+TJUHf8fmKDRrLNLk04XmVDzdWltYcBpId/zLxL
tm2reIx9rblk5bcoSL24SuHMeqzAZxVxsDL7yK1RYkRFlBMytQJVS5EmHirIsO8d
l8e3+Qk3PKN4nmWKb7ZK82TKvoMd/sR0m+hxDwX8pIgn5fYnKkt4nCPAsFc/Pfcc
gtncq7iyu9xEHLEJ/DJpZ1RDcysaUA12rCDmuU6QKrTSxQD5ps5VETOl0OBHjmEa
pzu1glXlm9Bk0XR87bKgm4reB/FEIdM4dNak1rOI/RBEJrIpnKSPvR8fc0hktlr6
r3ArWkDINl5R62es3e6o/xeKnbd6eOIBr/gWk1mk80vUiimrtTv3D/DDQH4t4vZE
+HiaOwq9XmCQX1JUdkxnxBqyE7j+QH4Q9Rx20SB64zpu+X5yJhGnu+IFxSTwLWrc
tXDcPgsTrlMXW68qkdzbWHzBDDBRrCW6UmK25k/8ZSYcmrkdj6awjwTYX+tDX52K
XeeDLEKZA7dx1HQ2hQ/5DZT5aDDweYnsGZzhWeZ6cpI+rbeijM451iR9Ax1mYuZO
/kr4BewyD9WQks72Mdk7Z1qyfBLvcn5b+VxTY0Xozp6zJpffmdDiKlI/26AFl3HN
96a31zWLgluLKMQ6WaSE90JtYj3I/g9e1c/r9NZo28oqMg/eyw9rt6CmNacgWgyE
etYTy5ONwtJVrPNcJ3xVhybSUH0SigzdfeZDGOytrC8j7UZJg95lpyVt5RAXaECe
EIjQX6Pu8VZ0FX8QM2S7gdJKz6SqTclVm3mGUu+KFsteTpVLtKePxJGpq+5DrEie
WGEtq/YqIQhloquCGtuZ61yChJ8PlmdfE/XTxDSmTwkzPsZxXdwdeQmLTlbg1/pw
eYA6S/Jxe/kNiHkJh+DZkWa+QfTf8JQuoGZojRkt3+KVI5XwbqPhW7kSB6/HNjO7
84TvnYv6CFkznBgm12eh+A5eFNwfit5CusaiabjLUDnFn36YPEsg2kYNkANObTq1
s9xKegr60naJRb4+VCgPeJ/uc6S57kYAF64MgBEdxEtF26nvo7GU0jodWZmknaeO
ohwTT30GW1XB39umO1y4g30VgvLnUfOdInZYjgfv4NKu2FFxaHZ4R+NskSeTOlfb
IYk2rqSmrgICRBFL34oHzdF2/anp2jua2QPjniWPomVkFpsvJadwNIBZ/TNEFG1p
z4dI3N63shXoq6tj3WzKFq2hYlYL918TTzyeIyXye2hirMJ8dp797rsJqHUBsYSG
klzSzp8cKT1OA8W0j77MBVY6YaHobFfMw59c1s8jp1BivOBtsMCbAj8QJBwMEvRS
yLcPivJhWnJ5oBDczfaE2zvSTNI+U/d1QHH4OyPPYt03xCxY8/e0sSjD8cL2RFNB
ipRFZpbFUcLQSKUffoOz1xfDQYocbcex0hiqlWMQiQXBvjhdEk43PDXXKxEctzZL
AUwjkZO6i0F0O33DwBV3xivEZMXrrsDNJAIf+vLekIKOCp9KjuXVuOarbt0DpAX1
mLReq4fDN5ff66mG8xtr7u20dsznT31EAhd5DNn/j/6V4VdGvHOTkx3L8xK9+CRB
6GehlFRUwYORttcI0a/Eb4StwH4fLpCktK23zSGCRFYRpQnmQyKFOqXMWFW88yc1
v0fe5COjyjHBP3LE4AwY+juh2tw0XqnZu0w4jsSlAGvu9vVK6IcYe3KfyAlovJge
XZbb/xastbbmlOuuiRONJe+2EugXe7e3g1PeK5t5sw6ZygeSU7XI8LQignZTgAwH
Z9rFPJDb9ImuyYZJPsBCm+fGO/tHLkWY6VknFzCPHSBx0K7ZvCvfTvamzE5ocrdV
XNmWrmcGqEDj1vzLis0GnN431eiEjSlztgSN9LQY4ympEj9KxoMzuciOFtpTYTMe
E/S1O8kW/rgOVZ1s9pd1UWf7nxPcc4tFWhD2FtTHM7lbr5Hl6olX2Fw6rg9YR7uM
IPkRpd5QPfuYA+WL95fuInbElxCEm9ZRXtWV7Hsd8B8rOCw4bQN0MKmKopjd6fDW
VB4qInkI3KgiPHBa1l1oWTrI5d1CpJPivhJVWcDkSrP3baNEigSzi5TMabL42Mpj
3zEZD5JzAI3bCkM5N3HPLQIt3VirM/+eRaCbySvq0hn8JsJvc8F0pxstxwcaiTMV
XWtk89KnR34hDUof5x6O2DPuReHMC5jG3WdDpj842DeprT//4B4Bb3ROJJDoFI7P
VXgO4CcSsp+G8k1dan3uzUs/u+WC7PJGTDxOMvbEaZfO/zbl3dbmkkJeE/og8KWw
JCF5teCx/vU0Zu3bxz8qfm/eilyAbLgUH5zEcTxgk5XP5cebBwbAdHW396T1BseO
Z3u53Qe6KRnGN6eCnH8aaCKlo9cZpAgqdfaIIOQGnFzNYzwfiqo3BBC9i4h1mqDf
Pl+11D4YUEzsq27Hm29vspUUhU5mwIWkQ9nB+RZ+8hsNY24Zfggw4IQ3nPWOT2b8
F2xybuLdFTdRMbsRzj6gWVGwN4RGgqccsE4pPmZVTJMNqV1qYq18y0/nSmzBIjcl
4zWxBTOyeqmPRJj5T+CySeFqseoTRvpziFQmaXEz6iTHnIjxztEGCBhl0DdOGL+7
mwweTfq6n+B7AyYUduDOkLOCjUwvQSvl2b8wV3bjHlj5QxdYDg9y2sagHmizk/FT
LKUqLc4gliFfkN61TK+zIDUntZhyKxy1V402x1dozx7rZntVFETe96j76NfCgUcU
U0OVt0U7Y3S+1xFI3PPoQsxSyrja/ZpEk8p3l4xE2pqr+tIlOyNNkbuwZxoqMgxq
T/pfgYklqryUQsSngtAHYb9soISD2/u8jeQ8lpIW+ctRq2NX9T04fCXWv/Wd/3Un
wkehGUpIoBFzCXdoiEqUG4c6e1u1j//JiJIHXZ7/s0qNuNHhbNAVcFcQpi1PH5al
GINFdKqgHGc6qSxIdEv05dUn5C7ldtXVmDADubemPY9y1ibq9mFcm05kTBr5jToQ
m0FvFhfSz4HAYDHit25NxHOwNpVeaTGXTgTDnMWWL9uTXHX10WiU4k/FVLRWVPWk
yAlSGn8DLHqi8PfpWS4jeGzWLIjdgROMUySWttqdw49aFigBXOxYL22CH9u9Lo7T
APKGuRUA0QRUQEpVS6uSofwgB4T3OV0JWd94rZosIFKiueF8PX2WBsuFYpzDUvf1
54+moeS+8Rf3S+35zrKhjI2zaWPkzyFGmmDliAT1NExceQGPMRrxtfY1PDaX4IM0
jZPyQ0WkutGRVZh+3s4WHoRkQbOeHO2FH8m0XcHDCAjg+CASzipzOUf0r4G2iZxh
UmnvSSuQzgcH0E2A1i3YnbZ9XwFpawvsr8KitG/MxJieWq56Bp0lv+Fku1EMJuXl
zx0D5HS2LEua3/wVaU/Sf5HNWnPfnITN8edDnzozwF7FmEJfcnvjFqJEvfNfOLca
hI2tX2GBBfKBInWZ2aRHJlWL5rKLuPuQNvnO7JqWRlT0xxYPSUxAfEtddszVDSCh
3qPIQM6yXLzhCG87f9pMdVNJ/CzYTv25xfKcvu2a9h7eZT3H6xKVMoHCT0RnzGom
UydIdxG1nNWF1MtqXT2Db2arS27QSFYlbmMNn0X1GwyxXPTwh8XD+LJ6B8NYko7C
YRSsGkUOU/dlu7u3cjrcqMz+GEFY3tDP7LEp/wS3zEKUwLYqJQuaXHvMp+BeDWpo
JZmgum1PBwosjK0SGM5z1V0EM+NnvN1S+7tLY6jrNv9v31FIjaXM5RBns/kMiww8
SReWwGlcQW0t8cOKq/yzqM9OBzs6fkE0FYmJ1JATkJ9ziasgD9XUGduZBEXfvHwt
BYeZMhmEzrlytSy6AxVkGxjaIcr/YL0ewEAQ3xgLEqLrpTMxOdr3mNwApVqT8CUk
zeQ2fg+2XrkdlliSZndaaYDqL12KB8R+YnjdOLuO6YNNc4ZSPve+fPx++M8b3xcm
4qAnbzkfsnYuhSV1qEVuNMbDlvl2LGjhdZyaLBszdRtgTY3ois8m6/4OsRIzt2T4
Jp8ynATLZ3rZqVIxQqVrGGry7hGUFiTC1t8asKD047dvqtWtKnmq6Lg13NHR7ap8
/lGDfCBh+ASQuFJVUP0TtTlLQAvsC59mWd0j5p85Yge7o9iKIMZ0jAgPqzCdkvn1
JJ7Y9RUySmeYcAUF7ndYN7AHTYQHpf77Zh7khvY1lJwNC0o27/n6W7HqFaqRWyA5
wjrkQws0rvECbjBeL/NgC/Tsh8ecA1Uy8boSL7SByaLHwH13soQQ9WxrB6lK+AFW
FCq3zp4jx6RTW2AWDrpyL2VAd8n4SaMvOvseBm7/SC8OLkV/of6H08Da+mSsd7Lb
yjQjl5P1/3UKt7mq24DEVAnoAWsaxxauoMydCQYVR2kMirzLtUZxBiyHZQ4RIR+Z
n9JC/EjZJScRuCYEc/LuH2Dfhtb7ssCYTYxS2nfS6TFAuNfcwTI0b8OpO+4Hn0XM
A0f/5ONm1JHOCkK0AnSVJpvdarSmZ3Od8RFXX6B4SdYQixF1YzE8ZmxVmBJ+7okS
kiN8OZAQZhWGzJ74u/Vf2fWrN/Sa9Mt1sZnxyzG3zTrf3z9cK0W+kzoJ4Be5QnsM
+OkCRcZI+OluOGQ1vFuj7Ul02zLk6xv5IJMGe8qBhZtD+XUI92+keyzElY5Iv2pu
`protect end_protected