`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6656 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
xsYj4ZwXcxl9cxOXlpzXHd1Jp9ZbwW7Zr4FrijxhTzV+oF4r9hg8B6kAzU4xaaht
CUy+rn/u5yc7iI7qeXJOH2QuwU6WLQcNhogcQfsjNhhBKDLQMQe9lsUSBZTP0atm
evahYzPr/lKS42rg9iiDM6rgecByRxvL/28SW5MqDOPDJfbQVUwGI1PT7jvN6gXu
DQRMKXfR0JTRixw9X1MeeoAp3k0NnQtqr4Hs51SV+330eHn3oecXkQzU6vpf71j9
bnJAmdHCS+9huNMSAW7vVqJotIs4NcpZYug5zUHCLsUAxU0z28KlZ48+tPk1P3VH
swxlh1KIBQ2snAn14KWWm8I9/ZRZU3egf1ArF3HDSrVaaU9dHVihvm+kAWX82Z5l
V8W0buOvaxSlcF8D3Z4qHNZnwa3bDt2wKkSV0z5VEJ5EDGJTK+zaXsONn0+4H2xR
P3NRq6H2FuhPwyR6DWKptQynsyciMOrq+KV+Dpdgkkn4oco8rPVZR31ld83kPber
351MlrJAja7HCIpHk77N23XyX/+agOAGs3G25FS2xEyzQKap+TBEkC+510zxuiQS
6vdMW87m55xZiTTX5QU26B1ONvLDRJ7bSj4RH4SsCQexf+O4S2PPsND04tbg550V
WDz69FI7c7m3FCACWVXBZB2XScYuG0ghOkds3XHiWQ2E0gu/+b4kwfeHfZ97JyBR
LrGcgjl46IS4HX7Wzi7Vd/pdxLFK5Khg8ZBdt5DfoN5Bi28eMVnyzhslBtbxD7OP
PKaSvLI27eWTZOCpI6GiCCambdVnaWjO8Im36B/g3PFQLH97jPleB0co4uGHxU/Y
KWzAuW7EnBq3X/h3iaHrJyGsmSOIuS7RitlVxxARTB2fHclLgRqAktRr04IeymXP
9aRBuDeVh27R0KYjnS2SUESXJMRv/K05d7HGH0WgUhDziwYr5xoBT+PG5KxhUPC2
IFtGJVdMd7L502J50xBfQ7uk+qBnSSlY22+qo9dRo6oNV07Z7UueDAB0OYn5y3Um
HDG4Q7+F+gJEbKKaWNTzJp9u1WtDi5cp3XArMtl9N8n5v3oBcbBZ2glf0TdJIkl4
J+3CZxBZ/vrbMo22Q5B0ia1p6oWP0G9Fazid0icccrAC7LUAr+Uww5RSQZdYDo6Z
Skk6mLNJw12ynC6KQZivn1AkdNNtr+xpXryx6gdyuT259zS4XEVidrtib2lRYWfF
Pm9JrADhjCfqWmEVsLeotctPMP1QJfUQOW9OiPdHuXDFQ4MOkSZyLIFOAI/iVRi8
VBzU3rY0ptOnRQuxxBWO/7upO7gzbs8eCux3g4XEjzSNWggnKoa8uMkbbUHazFxT
ad7cp2HYIsdJA0pBOGpyRXa2ZGV6mfLbxZYPHl6UJhwOuq+mAhpIoA9RGHeRmqhu
LxAKNaI4oLOfYyHIUTUhrABoo43LaEqysYM+pXB5JfvbJ4CseyeTwseN6ZyxXIJZ
jG51lBkdgAFwNYr4ep81RODcKH2+whk7Sk1FLxJKSYIxa++nff0CsBv7yweOhIQn
MdG2SMaDVOzJmK9o5VxgbIDAzH5yzJvqpWKIAsGtoRiyKbC9hJaw0/tP87MI1gYq
zfUtiftIwHmbBfjduE9i1TI4Sw9CdkOWPAXli1h/OVRaFTqwP6plnBuB/ZcfXhDS
EYwJP/tHNZ6qxXjoyG8ETsmZ9RRqvhe5xpQES0xZYxDY8K1Q5aBesuaP9vTOPTrh
CfcFq55XEuXACUdnaxCDcO791mnpi1tIvI+l/oNFtlGEjRfPgWXXSEO5c6gF8x+6
x9HLOST8wPHjch4V0wE48Pz65VTk0Bi84BSYOndc/fm1L+K0HKBw9a+8GjRC1hI1
IqOzziRCv5WJpcQNNSARry/C+xsXnCQppTc4gQoSVdpRj4EZ6YQRazazZKX2bKeY
wNygVg1Ro/Cs9cug/6pCKXT6Toon3F/V/XZaMsheI2b2NQr1PlQpaygGrQRxAlc+
/D6pcXarQE+CqofyHnASyyjDhKvzUpwHZ0DPMM/matgSfJs3UZ/05Imf26s1DzIe
yrGygZ8uvubWU4y/SAL2dpL1wQO/vGG76hkh52/Zn3em5B+2WxNmK7kGfh7a4Ys0
9VujwqODRt5QHlxW8rniERKg7a/O+z2N5QyRv+3svFVhOucy6aTofL7jPGoMcJKg
LAT2HSZ7vN7/wBTEffDE9ck3SJDqUzwhMtjWoOYxgiBdfy9LL4EZLFx+1VVi/FKz
e7AX9z97B3qMYD9W1s/t0Ms28qwEXAK9atEIHQ0ndfGVSEZi+c/A5fLGqxPu4+WT
EUolcLtH7SsaKWMLf84dda8Vv6czjdR2KwiYUdgmtLDbkt7+DVA+7Us3BipXwodu
4hFKlJ/wrZo9oh8BtR6US+AfX1CjJpU8yhmvwL0aI5ZLkILNIWtfyFjKMUW7fmIU
J87EncVK+0bYyoWOYIqtAm0oDiulX7x6jFDAuY2KH0l3TfsW7aVXiL/2hWvuLerE
SHrdp7lLALOlWt2PiQ6vhRI6iTIjMKfpAwa9fjqkeLlewTHQCVFM3j8+Q1jOA+Yr
WPHQBlv1oVridIZ4x3Wz/X7uBJqOIeSffm+OsL1cj3SOKYs4tm/aGBbDXFjS0veN
g45OdEvf677ZZpUMLChsbbPe396e07JaoS/8UxWR283VGfjzN0W+mI+PPkv1yDyw
+3LRlQhYjchSi6Zj8azsPJxzfv8684SmXZoisettQjw0UnbzQMzxOA/EdmaAgI2J
rIgFeprrotCLD2j7Gk+Gkz+Rb9Fj7GV1HpXzHh7Lybsomqy8Z2qBUahKO3FiY6nx
n1XkG/i1mU8vB+Nt9T6LcEqjaLg1Wg6Bd4nSO4onAafzs2ViiJS2917oZBHWkW7i
JlSe674doFRXeDpZAH8tSWqE13AABlWRLRstZnp3gfv3kjT73Rs1YRMQAweBPSez
erjczUFYuNiHh0l+sRnmzW34glCspkX1dUTta/Qu16X/7NZ6I+Q8VxfroCUJyF92
4xlzEd53+jXQ3rlPtjhSUiyfWCPoPL9tU7wYcyj6myigkRhK8+ux3ZkXQ+2JCrAh
PjhQ5Jj+gqy1PAKOCo6rnUN0sqQe1qeaA7eb2TeJ3qLv9VHyOyhRV741qhk6QaYk
YYsjT2u8+QgLJ4fAovtEI0FMUF20wB1l38O7rbCw31mD3yEXeRfUlEnIzTCH7Rku
8elf226Yf6Bd0XSeWyp61kHRnbm9fHI2jKQ2Bl9qDjMn+Df9EKrL5/1HnBm97uYL
YcLEwvCTvTbsDA9S5b8NApiZ2F/k36DfPioyRzbX13SvU2CtCHLkuaXcQDaL4McJ
uV8ab5QdASo32Kc5J3/tQxQbCXpV0d5OgjQSLo8QAD0ZkwEr1SiQVOyBgyMaNE5B
xeABvwrKKFvTSX8CGH44GpzqjgkcLgoiJpvYGjjSQtSDJP56vzy4Lllz//enetyG
EDkSqv6CaMI8FE3NLS6rQO7WyRWNhGPCLHb8eXdlz6aSiD3asiWv1289Fp+rKsPc
qDLba3CA4B4/xQHQbvPoDEQ2eQTnUXbRNb4by6EfrMAaGXNy3EQLJcLAQHJui7DD
hLvlnv+0suSufYl1GI33uxBMbkVZvoHsQQsCajgeHyWKXrt7P9bN6lln0vzdBRSc
ZJh61CdiPfubwUMNY/Qax7dV8ryu/iv0mAaWU8qljzje4Y9zEadB5rlttx1rX0jP
MfjRBV8ymOeg3u0C2usjl0YMkuy/31bX+YyyvzyEGBq0kBGTvOdYVmnQ5ZGkKSV1
p/wyzjNN6c58EXZA6BVi/X93jVzRslt0tKJx1Lr0LecAfU2gsB5PnIxPpU5dsvLG
9iyHz8QCDKKCR8yvVcUlHqOEsBUE9+CdMqAMCYOXREHijMRBL4W0yiWDjCsEbiwz
GUFKAIpmLiKNEDyu5vY4d2E1rc4AJQ3m9otxi8fVINgyP4jXqScSpSG8rs/4Wzi2
uuP+x2j8deBgI7NScjv2li1D1DHDr4cn0Z5axSNBjr1z96QzKtFmJp+cc7vkE3bo
EizXrIOgECK3j2Dm3Dn/OkCo+pxiGt9BJkFzkFbWUErMOSCV3XA+xwfXS8SCzToL
E7XJ3/sdhKL0vz+Hui+9a2rTvf+UZF7tYR3aPkhj2YrFTfjKqkdXJ+6MZ1XRLPw1
JM0EBcchNsJ9xvs366jCec1PeEtjrc2pYGO+YWlJYE/JMftJAZyHReL+zgD4HErA
sKVq44cIM5r2pPK76HOxwOeYBqOv7u2CSjZcC8YwSzWkdexZ3nk4FGuQRB7hUxwc
+HO66tX2opoj2oj0IpGEQ+fGfV2cYoqCGjE4ZQxLvOGGYbgXR+/cod3xWYViFIPW
+nDLnGvMFPLciJovYyo4VqPmKJGizmwgR+J/FUaLX++z64Gk6MOLUaiGy7n9vYTQ
5vVatzhPPrAf6iEqZzjppli78t81o9gZKlTKMh1ZxAOa7mlkUeI+GygGSr0ILN83
Dsxu4VpBIYsSiy5UK8Qo42JMNep1FTB36cfSMr4VBkbFxJTwcwT0vlk9fdqXkDtB
7uMTSec0moaqs1NFFx5p3dXkGOU1MeQDmtXIWg/WEy4YacWrhctKFE1vWYxJUrJZ
OaG+LxR9BCioAAJTLPfbq8yjA443Z6mf78AHaup2bHa3+tLxi9Hfaar+vtgrrGTM
QAEwNRSG+N2kV/ZbiBIlgVlTtzyG/4Ga1hn4cRM2l9fe2mTM9DGQs6QRl9LMepxH
byXUJlLXuosTWQ7f0WWFpjWB6nrAU7ztmgkD/WhdBP24v8UPW1r4OfOERscclBy+
tWeD4XyC3p9tnqknnwGl1umOU2RVrnywjxME3TrAe6v7KZCWo0GFoEJaEz8EqqgQ
Dp0889RrcoPKrNzYq4pvVUfXjNohaEaZY8UrP6MsIkv/feiYq9QdTBIrcj+LijoX
tGNMSxzX7VaaKI7YY+XYsJ5yCaVLX+NVKhws+GnNsK88Jzx05mEERSQe9RYIiuVq
4Mn63vPrXDISezJokwPIzCa+oZpAMUfA6ghmo2gxsiYmURzHpV7idf8mnWTXj62F
1Z/tP4eLLt58Z1Onv67qQEKQ2VL8TUPXSgjA0aTw9CShvJZopL8QYblTqIRUX6d6
Dp7NIkoogdTp5neYw25XfHqmtXPowBZgts+sp5bp1sS+sv4MqxGfX0/nAdGYvxZ3
acQyGSOMnDBpbuurLYCygXTGJOm0CvgLjopaA6AyNNZCR2Vbf+xlOl2MxNSWP0Zo
N4Erz1yZstKLyw80foWG+CjbXheXjE9iPDezj+FDZ6gh8VVfjNH6ImLr1sS7hujv
d6kBmPKH29juV9nKFE4jGG6EBrFYMVQ5nWfSD3iXlBr4t9RLPoviuMns7KKuu1WH
lZT79vf3o7HFQEjlcnlh5eLiOk2WuLoB+sVaP1PneiGQpZKEjRuEOM821wI1dUjX
4tN2QM6wGiRiUkjsPePYZ1amt5fGk7DOe6dd5ORrphl0HY6px9w0uebBaqBNYtro
cVl84D/sPU5rrHfi9DVgYz5N2FxX5DNUl6UBycVf6wFmqd5L6WWXLt/eDpDgfgMI
jXyd1qVy02yYw3RxpoTar0p9sV5FuZ1oA2hjsQmVgGoUVzI74CdfAVl7SYgjpxeo
I8+wYVtPnpHrx0u7nMJ8iplE4EE8lvxW8gCFFWeIl8V0PxFlxPAXxSlb96yRCL1G
2xcTsRYEXb6br95uti/hlrzoZQMnbjAFPdfiwcp33EW3+AdfezpvchS9QvuoDVa5
l1qIDc+2wKO7WsXYtMt8wIfKVW/snxnS7gQi4x9baTdhUQeYC7nEpk824vXnYM4P
chjj0gB67/h8kPpyTsi7Nj23yGJT+5rsLu+Ul45BkX1g1frrFruvENA7mYazO7eX
SWbAxajpeJHy4RrFgqAStvA3OumKkX8lNUj3YLRqFlGWPZb5EBXPQl6o7Wggwz/L
21zcWs3KmKFIGVp2OynTklxCojE9PwU1ofCCpdZwsB1QjVsQ/7Ihivmy2CGBPDMQ
t1x+wjzDVssMA3tsYU/MZBz/HcrBjVKy68yNplc7ijhLgrsYIuutfB8XPSDY94XV
7om6MnJh+iQ556T6gPgNeDDX+ex25d81MV6vpdHZzxIEEf1bsBe6UMA+2Iw27HZj
oRtuC2LKwncKnukPhoiQawc0kWGWhkgfG+j9xOKrhJ6gjkmH6LIfa4vtXmJW2Z8o
a1/PQmBwvr5tqZnErp+4vVn4lnsQ9pcfzrV1U/alDTbRkN6QggCvDj4pDunxSOHz
lkHsHI9YBd/T0WliJCojgrw/Nywh6jHT2Kr/gzDeAAHcQsipmSVsCi5ZRl0bKjeh
+WilPC2wJjPYTeeRMRlvLV4AoWC/5IGES7A5S36zb1VkTwyV8pAtmsi0t4MnyelC
S0r568mJJBQqJ0r/ZlJdMWGbZRKod5toj+Ok5p62/kbJ32XFTVH5KiMLYNU331v4
F5nUj+/ompMGZ4vG7ZDYZcey4AvCwdqpIHOgzs/pY3bk3EQbhLYi7QY6vUOieEB5
FDKjutZWcjTWJzuRZAmrAhTP8IJWiBX+VvuXYaB5wZssjNX/Trggoj6JmKo012K4
jKm68qPxGxRa2ROuqYMT6ovvADJ+CmjRJaeyK1Ye+dRBCBVL78eSZ56yelo22tOQ
hLRGs1GmtcNFd+GnzncN6qptwm2LdSkmfPircxeDSPqQr4czy/fPSeAGEn6PdXV5
VEiMpccnEYlji7/uAKSskqox1cl6AHcUvtCxTnh9zjnfdfy5bzTFRdy/ZjcR1Ydm
jzDqqTkEX5jypdK5viQa6n3qE29VpU7D3brF9yOK1C2MaD+LYpXoM2WktATUnvEf
cAb0HNySrywd+YnbbYl/kpv5y2okt9lFkNOLffVvPCHnKyfDbcUZuKb7wB8eG9JI
RzwJN5Lbgo47xnxNvHeI0PX28VquxmSeiEqv3DrLx1BQMYrHC/9gOeFnA2nlbfH4
OUxyqk92q+R/s2BOPQQ5XpAh2Ky4pZ54LZ3X+NywLSwUQVE49Tyj7SXhRcqN6enl
U8rVZgm7Sp8bQ03DFDaz/XfhnNOm1PKMdCmzuWXQ1wFh9yzQCGa2co6p7MxLbN+z
WFujNdIke8YrXSYK/ZS9b5bBuBdUycS72FFK442twNFzDl45SEqIJRXt829TtpUA
5oyKKkCIvK+G48XQQZq66YjNZ2LOU6ZWLcwJEXdr9iAHi9k0rc19PClfMrPcBX9W
fjocXbbp1YcDpDfm9h9NJFMB2pOb4AUgETVSNRF8erWxkl6Y9GlUImxw1dwJ6ApV
2vX1IkGEm1wuSWcAj+lRfBRtkm3wHJHMDSX/MMZJGR6pXxD2yRcc+tkL5/9Bqdb3
IQyFTKLHZZbUMyOnqhnmg7Q4nEbfcPMER0kcySFCzQJQgC4X/eY0aP12aujgDGrw
vYURc2qWkqZX7camSyPIcm3+IflgdfluD6U5MBUXB+5Ym6zgqOTSFAwXCR4SJ9lH
OwHedMNnfgh5I+9Q4SOrNGUxmbfq8Ct4IvgJeaoLnTCxbX1zKGxqtfos4a2o+tLo
SaLxEDlyXzrzGKT2yQ1HQdaez/vchW/p8U0MXSHIBZh6+1O0o10QjURazrjKWmNo
q5jqZgtxbOJMo30KWLP/g+QjMIA0d4vviTAgGrgrj+WX44Br6m10207IJWIphprn
dthw3ZUPDPkwZGj0Ts00065+AcYgh5oYzAz/z1mCxKD5zsU5YYGYZMgHPb8E2pa+
R4Q7nYCzsYcuBsFmBjhGt+icTtUJb7oW1+zLR35iBJVJSC3Rf3usmAohgPBH5lRn
09tlEB7sqlLPj0yR8Iz6n5DQqtnIbeUwlul1HGmlDbMB5ZiQ24j6wZxyby9iBsBq
DA0KMxp6fdHt08ErE88TJT4kImPpuvO8NO26Ef1DwoPmLYz8IxAoDB7a9kIJYIWY
CXDQVSbqosHs6zrH0FmLUBmHWY+QXfaZgzAMAGYm1rNhGnEGTUZQJEkbZ/hYd7mw
FpD9Pi/JWDvsZYVaeQb16y70piYeNScaXDbroEY8e8EKfz0SZ+SILqzvw8QHpveK
gKOUXktDO5h+QjSKgOLI4PJcxyWgEz1eYsXfKkzeCbM/tlxCqbTGff+EEc+d5Ye9
ABEDrbF5Aj9BRqHdNCMJE6nt4rPlsVHpeosmAtAQFw5E9y2WXNEy92IONz337ae5
oWJQueNEuX0QXHBn/FSb2yKOveAjwHnuM5W+DtQSACE/Qys1RCTkbgoLy0mjn02O
MTVZzujwX4kZyzAGf4X9eCBKki53IBSS1UofZtJY7qeedv2gGIw/YgUa/YOdPwud
9aTqAGUXEGuA8JrxKfORJfYx76cB+hxMQezuJ3BSOVTqPIIcWzu9QYrzBb2GO6qp
HTj6OpoTypGluwwM0b2naHeEPCkvIKsfZmnzqkHy1Vcpne36tkH6nPQfjYAFV2aW
6vURqAM3OIB1FudbyrUbMSD0oDIY8kIOMc8HO9ASdn0OsH9kjXCgr1P7MJLD82JP
EiKpXrl7ihAEGCIm9zSB8Aw9OaCS8fb0uSQwhjYYvuPZtg77YM0SgOhRdX7ocW+a
em16OdL3V/XtmQB/IhrPcyVXLiB+yqN8mcHcgLMbdAXhJSJUBVqBfd02GL0nEjsG
u6QdMa2G0vPypPLg1zXWqLGGI6l8eQ+5Erbp/yZqn3ySJngdBtaaWS1WAtuDIatT
1SV3UcX0DIjNOzDBZNWsY6uuuQ6/+GZjZHeqoUBsPiI=
`protect end_protected