`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
hVdJHWSfELCmA4ds+csnOQAALbB3ps7EiTSHEDd//nts1r+JQrRE4d3bDPRJpiX2
Sl8d+xAK9BIi4i+3ruAzYvB6kuD7r+gs02Jsvd/1kn7JYK4xBxCjtdDFjVHOTEl1
sSh1oNiYUwLuwR1yKfP+xBhqxD2Dv6pCKhH1NdGilpJQ6cvivGkSunAu0tzP76T0
4x1pB179E7uIeRplfHWX03KzEBF+eVtfgXVp2W1BGjfAe43y1pCvNYZOh1+TY62g
EgAFgbo7pAujZxZy/YSiZjUr2mGp7o83qMXyusx8+rQ41D3X6rxfuP0RiId2pOpC
6oq5Dfkx04a1dk4s8w8cVg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="Sm9DkM+kBxuxXCFA+l3fFkxuSWV4xqRc4Nn7Ji3ukao="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
m2emGBqRy4AuduN4dffN8194qYvc9UXRqiQc56IrQYMiIVQPyh59I8SYabcDdspI
7AFHnvKD5YaF6tQfxWm+mlcmMEk2Y//aUjxeiGGs+RkKgbHitJF/K7nqg1dmKvDg
a/GaBCq4Bqh0EehlN4ntP5HxM4qcvSfh5m/Coe3drc4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uG91daMWA1mGkhgP3oZKMYye3UAomMWgG80HuuXg2E0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
c9NqBF2D1wSep1rW7utzHsk2j40aow1MnrccxUTvKej2Q1cyeDDbgAml4eTSXI8z
QYgCADtWi7S8BeChdv4B2VxKcS7CMq/DaQrOy1MKTfQzfAlK0iubmlTkljLy0Rwd
YnZUZ21GCfDuQpqHcw47V0Ox8qopXJw1eFUtwqajCy5h52h5X+h0K+hxVeoY9KsO
te9UHIoWRdb5uBASHJ/C9IEOqKBeFpwvYfwWPnSwpQEDL65FpKa5gVKX0gTTCvtd
pAoh3tUnbQCH/p2/iGK35SzpjWYICLscPTWss4VoKvRcqte/E5K5hbEdu2qSA7Ag
5x51P0d+ZZw3iBmN0VMcJlpCez12AOBF/83a5dcOEaAJRAbPR4GpPCN4ZzjYj0gR
6NuLKZLkUUwuxPkkGSKvbbbAT0JX9r1HaNM88C1r5SK8MNITQJEBPD7vA63T+S+s
QMTWNvcUc26uY/C8Imh8uB2W0OVhK0gGoC8qmYZhnZOLjmDMU9ua2P2nuI7IZjqM
ioA/d3zJEn2rzkpkANr0VMldY4FkXt6MbjYdEpCQEqgPUdsKN9QB/NTL9xDb54gx
gHsFEF+6TwoLKjr01kbqj4EzuWJ1UKAb7XKtFnoQGueaq9ybZGCzEY69j3ifGAL7
jL7GWR0wX6QVpZ41sAMM+a1CRsjlfGnmmAsZw7sMepYwp4bqcLjp04zsQ4ZMhZAf
WiaTalQaYrApTKoUkIMDAlCbh8CLfyNSzJA8qx2mqkXuGT3SK6RS7eK68x/iPviw
j8sEgXVKI96owtyu6w7nyJ+Z5tu2g39i7xf/TuGu+Csz/wxKGJhklTS1gTRYUejB
AdYTf7tT6ImIWOKNC821nfibT8fwvqGbE08ErGO9h+FkQgID+NmmpT4zHXXKaxQf
UafeqLBW5CdhBCjti4aVh0O2WaCHoB2/6bw35gZ/qpqO7ve3S9ycSPXCwceYVvaI
1rVFSlbv6omUA1kn1yeL/EKMR9O+lheRjzABqB8sclfFadWhIsEzqiE6tUk93suU
aUbth8EQGinfvHkqE0XZsnEAKfi2MtuyY2Pg8wmsgsH9TwYF5QsLU5WC04HmdMJY
XpuF7ZshSDmwKc7wX2b6PZCzuL1BiF7D0RIKYK9EmqudGPvgWf82yo7jCWNjDxDo
VbWy/dK33a2H/1JSbtI2OP11gGVEuLs0ypVXZxvwAI/FfheACPo3D7m9VA1hlRuA
0Q2sUmxpi8VYzeWOGhJMf/YsFxRag207G5PzSJUqFCNYWAgIPk9Q1SfdHuQcpJNz
AHTdgBcl1I+DpsSGPXeciy1YWYkp8PCFFy1Sn5l312nYqaFcNge3ztgk6vqg7ZY3
6YcKgK/gcq7IVBklk0Ozzuj2PXz75W43vBchuZSbgr04MQM3bEdIHTsJW3bwDGkK
gE7v5W8DNJ/5aV1LQknUy5NagdwUHEIf1bdzqbnJGN4FOAgHMC/CJ/iUiZB4Kggl
OLBoXEYWqau4HvcdY9iVW/OqMnFv7If+5gTgfenzvnNDpu8jYuYWjAXgk1jRteVH
Oe96GJ3k4lIjhBMbLwnIjCs7C18Ofn0LOXUg6bBjRgGhH9+YSomWDn14HScaUUwp
FuRVkshEdYhRdEUbuVHsTJXcJXUmfxF6f3/Z3xnO3ryXBlgwRsvilpXxcAfs91bx
xRZJ6KcReyTJOsD/3nJz1XekJ5ZNq4aiaCen7fvkpvVHMbFZKvCjRO6w28O+K0uK
baSndRTHFAQCq7FGgukupOiIBMkUQlrWu7FYPY2znOpxwZQxRLyn6iD0lUC+zgmR
ZEEbN1twrU5EbhTQLMO4CIfN5Ah4Ds4VfkuG5GMr36bPo944T8+UYeyi71kiLpbb
ZGu8lmE/qfeHk9XurYWCrGaVCrw/pzk8cjveYYh6wqdPdqpG8UcjKlVpAa6yHHhp
DBoZZZ2Hr0eVahTmu193yKiYkCaj0S7Ysv3+JdHeoDJeFAIAqSw6L67lD8p5hyfn
HLIhqsTLLCYFGQcsGl7PffinTf+KbnXZ5hHGIrohv4RB/6400iARmHyR7lcbcu23
WTKk3MhoPODtB7F3f7pPwIWbLu0aVDH3JzEnT4aw1d+2P0t16lBuuHRUtRO+USUL
O240ZFczoAfm8wkHT4No6MiEOcW36T95WKRVEPLUjVCEKIkPtO55iJsqtMkzISf8
8ovG3X2MLYpL3WeM81nFOU52GOlUNCS/deYfKR4MHyNHomXjUKgghk2jPpwmbE/P
T09oZ9DQcv+L/31YdRCO8ONa1x541G22KSBsG566lWA=
`protect end_protected