`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10080 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JWeJJ6Ze92g4+4wPuytvzVq
BUiIjW6BqLMgOdxnHw5DNWEQW/Ew2db/LEgoa101VlQcLbk7zrOOSuf7jO554NkK
LvIZzGhSCaoZNdRsHZRGRAaAr3dJqHoskhmWfwhLQa5CDYVyj6NoaA3VK54CQv1m
4lbpNoVgLNUOqrthe4uDHYBmQgikGIuCPGyij8/X3gXr3CO/EaUx7U+EAMohUAYy
VnC0VN/dioUoX89iYiaRGS0mnHSdpcLmW6s/mFKB+MTDaYpGThvqo/q6AzUiY/85
+CcMQINMEVGsOQ46l3Ly8uKIB4ZwQ0At7yatZ3Gst1WerI4nvaUJtb6TI5dUyQT1
Z5W4MvyMWEm4ePGyXsavkPfyjHU9Wn4DgsZBWp32gmr2Auf/6bRpBZ1sjduD2UIW
1p197gsIbvpyfW4r50agjE8I+S+aaSZdhM2oC9fX39aH2GuXhdoFB2U5x/IvwuJg
tYHM4W52EIp+1/lakcE0fSg7eaAaUX39Vg4cyRdDgcojsv+4rVF9EfMu0C9C+E5a
dupKyB82730J0xvCqHCxfTPynZKsBOa/n1ATDq7ymIXqv+T73ka4nUKE6eeTD00X
UZH8k+dMc9Vz4bq3D5ppSQwo5E+O5AC25y4AaDI0XUxDUNXyD0jmTwaUSDKB985K
/wFarIERcFNochNomsM+UqkSgRzT7S9xG/od1REFxjqz3e/PiZS7OfRnrQaKdFoi
VtRwdDx5XWcIHzX1NXkrwWF90/laTUpwTccIbdEQTBiVf+qoY1OI+z1p0ukAY8IM
4ejubMxHcYyrw1eGeZtQW+P6bx5tEmZ/Whpzyv3/xDB/4yjFv/JpHcPuHLUho0NG
wrLc9YoOm2GPzvPuODqGlLsk4GJwOpDny9bxOiskcYIXQoSZsrCWpd0wyZvsKDbJ
7BGJqQmtMXl4oiqYE3b5YwPhmfM4frX7ce1XceFwzGl3mhSCWq5LOwpoUTnP4xLT
VT4KcI1s+q5KGCfFCee53pISkEXhACQfTHlb4g/YagW+WmbeGjUL6L3MHqGuT/rU
evKf46vq5t3tN4+hOsJ75kkUDfb1CBSfdI6oS4Mw1tl4DaX3jkQVM3c5mn/cxNvN
GpaQeEF+xDJYTi53WsxmmcXAobQb972p8BE+XtATRO9Ylta0PDCFR7zD5qTbgdRs
oRtnrx0WfZrD4Ppt//wCR8t3TK1GDqPC3PZyOKxQMycSym89/+3YYdQSkqiw07sV
vfWYcQ7n/sJ2YkYaORyzmS+LUDaJpBf9EunQ619EwNhqtH+2JrLzNo5Kz70J0D0A
83Dg5701JsOPckLybF9mxrrlijSBeG46I+E7icBkg1KXeY8k0AJTZ0H+3zoVF7zA
KKQ8LzJ+4Qv9wYfUv0y9GboGL2fseViUutm8HOnSnh1OAnWB6Yty3oAXGKob/Won
tbJFsWPl+bxZQ2A8o+A7kXQba/hKYDOmQeKllFSZCk9jOj/a4BBD5tpYVdIQzFyC
xA9/V2RpTQeW8DC541ToNYiRc+XNul6TymeuZW8GLf7DAbvDGaI5XMTQbms9MeA/
y0iVNCcR4SiFPOrLHwJ85cwPPuLcsKgukbmr0eXN0C0VFLhb4Ya+rVcznIALz0bG
3VqnhLGKoF8I2Q8wdsNb5StK+Hxlsw3IaIkH/GRcvw1A4hmJkIcn+TcdSSY9xUhH
otzYnr74lI4xkG9Z23VYUrk1jUCG3gsvB7jntr3zVc6a0BjYXdmRStnpVoVLtgym
XDgd3I3sKZb8URuUJz0/UxUHMlobneJdrMi05vzomXCvEHwqwGhj5Q0czVGsSpWs
dZoSPumWJEtBGO3pu6d/Uomvg30YR74x6llRnfFdi57Bxr/GUiM0CkA9IZ0N8gU1
lQpfnMDLCQpQkArCFhyNnQcKT/8T3iWML3mcAgWFaggM7YAOcjQBpCriqnCmLw8A
u/u8fDfmHldZpaKfNsBiCMBKs25hkshPh7otlatxlj398iN0dAab0HfKYsgwhM/e
QsS5/60btmkMZRX2AFjH/oo3HSAm2Wn5s4QdzgIiZD0synKyl/Q+A6omxro/rv7B
h+h8BE1/N88C1pZeVmKsZW8cPGTZNrh4V2dmvjB9RLzCR4itk4s7dgvIZKd5zKQ1
GEdAvxqvoRjsCf+rhLDT7OfAy8F9G3ojnIAy76GJrysTUlAkE8Jp3Vi3nou1ofci
A4PS/C3bDZjDFyGkbFmOuNvvNvZHyGIA66qy7fUckZXpjtSZ9ciurZZRfN+Oykbe
U4oc4XLBbF8jXPbQCqR7UzeTxiPDKj/IY2VTss6wVAsmfnzGZs6IMOuebvPYb0yF
XFI0oIweZIhR1YmY9Yu6504+UiNU2NbGlyFlBRTBqSYGweiPrGinh6T4Wf/0lA05
rQZjouu0fpP7RlRC3xZFrnKK1/qtD8lSBXD9HMEuTEAOT98mNoS4KdJcQ9syiF7V
Eki9M+78kcvBvGi9ATHZPwfzaCOc1OWb2wvnBzgD4fQoPXzg+tHBLwAQ5JYu701j
3jdRB5cclU6HeV8T4C2UhpBErNuUwkdXukriszR+m/sv4/A8t9CYjA+ovHj5zVwm
fPP8u1TTIZynMh+Vv/KT62roa+9NtHGmQB5/cml6YTm4TZ9pvUmA49w7fUfaTzt3
JRzIBA1Y4FnXGSD3mBvBpwg/v+WganuHXt079s3EDhOf/hiNb1AeTVH0eufvLTv8
yuqRU/aArm7BQL6HPs8SVewWTpUYa0VD1q4U/SRhqxzvCk2gzc91QcNo4dSJM3vH
nvymp+o4l2ZSyVBiXGr3rsqCCr7TnGym2Z9POkE2EI4VIYmIxCtaYouhIZyXn2zw
PgzBzYIM66/GOS/Uu32SNkbmIhd/kHw7vawCXvtQpjCFz2c0IBvTkPQq6kAtSntY
9wX/yopHDaUN6U7Ae5y3EAzKr/JGh5yFgwVFw0pcm7IyHRusa8+MLr2MiatT+pOr
EQBEWXjnK2DlCpsg1R6Z25RDh50Ahqlqg8neLGrVb/B4xORgIv51x68VQ1rv0486
Zczs3WbbQujbmHhIbyzRJ+bLRGmJUSFUE8YiMPmhcxI4ZSx2WQOTeE2w3rJ2x52+
jG+a+mvbyTRAt2oMvDw5J3Fli5ws2jw36Cn/umOn5fMtiehvrt1FtjKuUTFs9YRo
FsBTbNnamGpnYPjDSofms0Ifusjr8Nsgb70xuxlSLpkA/dlD856XaBYOWgFZXO1x
XwtZI5z+tq7R/c2ymaBGYAypcxMXUeySmeZ8dv+cPZm946vmDtuYdFYAFlmPMqAa
Fu0fvK4EdxKgPHVZIz5KHJP89lmDz8MUH1rm0FQUcMmGoTHIVTJBRWJiKS6ahs62
T9r7AiOzVXWRVrr2KNsB3eOt6V2Wh6gsuBE+OfS2xZsOmB/0OCVYUy2NttPMUd2m
eek3bpE/mj3rQEcTi4kag/w/0MTPGQW0L/xpZMAKFdsD8FMyv8jHo436HhU87ygh
kbRZdiTuUg4Tv85WV6GQLHcs772nDHlS6ppJOrBfNfKAGp8GVti+/M6b9q6LPrbv
KPJApT9M/9oVL3gOm9erZ21gaIiB60kG6cKVK0ZOhpZ5jZHDihMcMCNWwRNYWvcy
KzrVArLdktp3O00mZmeEOrYBRZR15aEbLPyi6FPwi6Siyk4lPXfEV22SivXa4/fx
72xLkidedpTB7YD+v3LleNYCLvRtxzKouXwfXf8Ht9BVX3C/uPwvG4k6yLqStWxw
EMVtLNfswZdgO/vTbxJnNhdaSEv2Yff3dw+3xZldXZmgxmuNr8mo80qc2ECnT37p
jq8kSbHIuZolvL7ZT+4hrpJBaDl76ZlkHQOKG5lFFw7NIUUWDZDkkr1FcQsGmXy8
ZQ6I5Wwy/hbMg5xB4ynNIRMZr1gfwsVF7B//EtReSMC9LDLIRLkS6sgTe7MC/RTC
umM4BO19A4N7DvFQQTanIg7sFZapr8fChrAmQQ05dXeFBtIRuEbBnIk0o2/XMWxx
CY+VFMtGCLfTSBKiC30Dq8mdbHgxIFWi7n7+xLQcY26/b6D94Lmvf8w64ecNoh61
MFXGTJRd4916CZN4sUtf4pG8e4Zee5nc9wSvWO1LZNL4qxOLHKQ8GrwdMItRjRkG
aqps5S5k+9hD5urrnZjHRbrPe5c17PtXCsxj+McCoiCRvDxgbYHR/C35aUUJ7/sv
PaEjTiiS4dovqDujMe7+xYXKRntpH1uLNnwqoEkYMaU0VQcXzAvIXD2djLjjZIAR
QOPIrWUk6+N4uU9ZZmRXpKDMRaXBea2xCQvyc2YuNyKoqXoIF1MZINwad3S9txXU
HyqDfK9RYRBhWVzHJr1GQxibcQnGA0jhsaF2axDld0ykzukGfeF5605EDSWyp22p
rztHx1mrKvXEJ97OOAUyMcTtUkHDHcuPgEEAilXnP2IJcnq7G539bMUc0uIQzk6b
dEhGiN8LYEHvuxZtEvmBsCbAKhs+lyq8v5ibArbdE10PT3sEEgwz74Uuog50Qioa
OaJmPrNkdL5+X0sNf2ZZo+DgX2TzrwRnmKrOzbVam85QF9suSsmhSQgRShomVhUt
inE2GoebQ15PUyFqWVx5vFYF84O9Kq/nNu6AXLNQSytygReQKtdxHU32Cw2Vnkyv
0CbIoVeU3uQDdlKbs5wrtNq5D5Y6Gdl/QT35Yf5rabwYJobgZF9r+IPjldKfNuxz
xndhJTBWpkyoV/ZCpL9Scw0AjO+ZRxLgBqPzRxAfcgWoH5Iw4o1xomCX2eMzgyFq
46R/z2tsuklZwhr55Uj6f9kscnARXHMrvAG/tpyneTf9Mo9YsLeWKf7gRajLhioC
RnlU+Ab5+++MKR5FFF2Gj428+lGJn8uNxTS3LUI0irOQisNDFdeCoCdoq+SBvfRN
pwGNX8jEKG7aAbho7xTEdM+qqXJg0yFV7WSrvv/xWT2Mh3nFuqMJBTKvD19gZXh6
UYK1UaeojdzzvIBOaj/ifskNp0/o//j5mxVBsXgSnYITiR7LV88RWmbRJH2glnem
T9BjDlwjI2axZgjokjtrQsK9IsALDi23IkZEes9TiqheWaWWjkIF0F2gXari0Xn9
9wC4SIudeDhUFYDcvQpG1YALZdll4wfXcI8UcXg326KdrDczhTKDvLIXmDHi8Pqc
Qr3a1boqKUmT4UZ2kDpW9qDgXLrDm14cRGfSRjugeqLV9n8qdUO0VwAivZ/qv6+8
VEf/u/hyzFnC1Sq8Xw2AaN19+guyht6JC81C3mGBOCl15FN9ZaaHBXMsU3Pexaes
q/wLB2SJ1nFrHd5pF5ctV0cZY8YAFPHy5n2YACuvJvkRU5oMenTj4bXNLo5VUCey
qrg3jBXXccBstcixxRbhTRfgmqkm3zWmX6Uo3gqJe1N9ZiFcRdx+fgHV9Ki8szN3
cnmE1mPTmTG6QSkr9fMTppnrPW39YVscokPgy+ptaStKcuLXJHvAJwfL0a1A5iX+
s4yNMR4FI8+DC8BooElV8PibTvFf7gURMHRHpO/ueH704tMUzWMZ6S9FCTGwZCdJ
3jC4mwh0xmgpsBw2/KEOE12YKYNXHSD3PxBbMn5JpQ+6i3lqhiw3alwCguHwyCQ7
Bg58IZQfBHr7LpwW0WGJkmI+zCaTMpKXBz2RWQZyOlzjGgQtUxrdC26aylLtytMQ
zW/KDf2aHA9XOFPwVcJZkaWwfKzk9y4iUVz7fxzBYwygzT3aBGL7ylih8rEt98fT
5Z7bSj38vXMbmTl/3fKw7T5CRX0rPRYHOWqirfDehvFIq8KL9Y+4JGljGu4SRx2s
NYPlTg3YFcwAu+yP4Oj8dNv6Z/5b2jpeGZi0ucssriY9Nbq+LQOFzojaJphEhyzj
O9OOnSWHET2lM1Z5RvNkq9DdY8YQr+ruB3uRqyxkMKYDrvyyMBHIEVdBIteNOfFk
72ka3adxMM5xAg1Is2moGJeoNg1D7gcADPKXpFLVCSF2SQIys0L9T0Bd/wlbMW2w
1l1h+SeBzIlcSm9jrScUUf99VsvjEv3My6P6G0AzbGKe5IREoDcoZvnryldczSrl
zfDczSebtDDOtPHT/fHXaXasgdN2W28XuyGvpDn1612yFnpaDpKcnZrTV+qQcN/J
/+/1c7mb4inLdEDMY3ss6ywJ6yOyM+3TNgSni8MTNTx5mI9Se94k1Geo4bZ2Z1p4
f1aJvO6enEyVtdgUlhWklNvO08CJ20/5WUcUqmNje2h/yNu36r0olqasFGMDAWdD
dtdTKfg2xyO1GG3Il0t2qKLT9/9GJSeVSb1aFk02EugkQ91Z9eLO5M1Y2mLJdm8g
nuukx1gtbJspjCfBj/6cZQT/sNfUvmBewXikIqmbKFz4yUipPyK+25rSMETnS4GZ
DgM1Ee3dSr0Yk+kYIy4efa88QFS7qcmyRU+uVvvUiyIh+RyarmRLz9l/zuifMXlk
46oVHuLyhuyKHbrsOOn0KwsGB6AkCC2y7cV/3GTg7X8qTKdGlDoXidZu4Vtd1Iz8
6F8CW1e8KixnpjyrptvO4zwEnqArO0C8R3Ex3ZDzyS0aSkqkl2SkojdnR54wEmIR
iA6DhmzNP1R6UkASqARFSK6ejFLx+oaqjGo3yjx7gBtH7aEKP/AAO99UHgyAuV9M
XWpoSlECvQuBTLTUCvnqR+qjANWUlKls9KB7PC62o0wZajJ61vQDdi1ClGaQFbJX
odE4MFPSP4leCxJEu5ypt2O1sePKaTFtL+fR8HokU4ayb8o3GDPcIQRnxZSdOqSE
P/lmot8qOq6MJdF2pMq5tp+vTxLDSzzfSBOV6OTTeIS4Ub1hJwGUXKo1cjOwqHWr
XvPo7PRNvBc0hPWycMJb4KmgQGPcul5f5SOR5ZbX/LwxeXkrg/Aga4fy2XTdw7k9
bViuywe0+MBNJoEM9wHsnUOuppbpy67NWFC31fZ7lHA9eOt4Bu+TKZGjQmFdPPmx
3byR9blmO2yISADtxNEN5vYMvgzCqnyJWxgH7RM+HdVkVFO0q6wjku3LnpfvZnzi
XC6yCgKmKgrqWFzvKw1EQCI17B8jJwT9cGOwx4x2swltcmKLgf0PhtZkXnwDoxdp
UD3/wSzBY3d1+qvnGPfzcJ4LmFezOEOpiHU1UpwfuJjcYhor/+FyEB1SAXXexzfT
w80OWeCa33WOn68aD373RqSqgwgL7HR/JTQlgq2x+XHjyf3OUoVheVlSuFp+g9xR
41vPBHr90JU69IN3PXwWTUcQet8xAHEHBeKSAC2u+4yXY+CWabxxCzu2cOZW/NKm
dE2rHfTigI9yLtPyln/qOSjqqvg4HxaKwpyv6D8hypIMv44TIdJojxHZ5erVcky8
d+Fy1WNOCsjSKicpb/LgDgxsAJEn+JsDlXavWDvjdPw+qUDpceSiolUKyrRt4AFv
0yT6ekBHmmRSXRkvqKSdIfC0zWj1exhj58QQTIHC3TMu9taonZUndG7TACArGdDd
M6yOBzuoQbiGEdDg5DAOYhpmRIdEJ4ybAz3CIZPA2sYcavt2MHCRjLg9354zmLSc
IFJn2d3Nc6w3vsmX1E01gepB2lr0Wbgydct+D/wpGhRZcmH2kKTFucYh9rRNl59r
IoTTwXJ9pddwKrDJiJy7+nTSFyD9Kq1xBz75qD6NTMsvLb3rMb8NZIJ00WopcH2y
SVkJUfppDX1t9pPdtw3aCjDOkyWUb2HzO7KZyqq02fxijWun/VPLTQBcfOS3/zff
LeR8ZmQv6GaMN593+M8lJUu8pzHU1pnhnsdtq0jH+XMKuRTZS1ZYvKQd36wb/KeQ
NDnWtgNdXHsRYeAWUGPZuC3Y7cabRi0cfq432JT51fc0gmRs0oI+eszvmC78PIQS
B+SDy8JbZQAiPZe2SGDTfh/iuee0ZS41/GiKr+vrbxadY++e9msBP++/eV1B5MKw
EwsnpA8SWLQ4RRwpIEGB89DkG0QLQJTiGb9kOfpbVsp4lYTtpZo6uiRg1sPIqAwz
SzSkgzbBYzbNrbWBwmA+DJebJbtQTXR8pyumKIAxaV8tlDMyayJm9hQy/8i9goat
55UJ74nMqrl2tsd3/bHwehhQJdWDbSyG6hj7sAA4d2qm6GK4qMV2mMVQBClrSiPl
UDguvEzsslytpxxx7YoPaJzjrAz6EyAUrY/C1NHnFU7bP50LfiKDyz7g1W08QLRB
j3poL7nU3ngXrATm3tTur/E0xRu48VoohwxwWDS+WYIdWZyWkROd4gpoCmIlfRih
GTvD8an8XoVrz3pgwP+vBbL8tSTEdaVFoGzum8S3kDCbUDJeHLGHFnT+OTolhzW6
iuPtkQWMQE9qeFWF0gemXjxLGYtEwmWCsjpyeIpd5o+4+xrtvgQsk8JUCAFQm1I4
CWIEidIz7/18mnLmm4uibMMQhPoYLiiafkgOwJYjV0A+2YG1qtq0M33pnSFDPOjP
rsMGtpQI6Do23KRn/fu1xPwYgXAr2YJpuGgf4c6Q8XzW2ihnKZ5iLQoEl6n7r4He
6I93FNURuC/VLzlvKncCqLlvir6pfNEBhSTAHhb1Ek8mR5ZQdUuv34MCF76XC1Nr
NfnrM0EPs5Iw85si7yijlYCfJbohQFRNtc8vGO4ue0oOpPn51+1gOYTtyw4A1wr3
t3yrizusKcXhHmRryFw6PznofWBpEx2U20lPvGWpKx9RMZDhfG2+2lu8Nmezv9uU
Nk68ETGS+6mzTBw8RgqVPr3hu1nJgVaupCH1GkBBZIervlGXVdma5QU39br2Owe4
nTIBn8JROgMCqnhVZn9ZkVzfkfIxeR1mk5ZZ5ztTB+IJ8rdArrgVSHe+d2PB+vOV
25TVfGmCfn6ThtqRESJNseK4oPTr0EbBwN8Q/QY+f/iGtdKxgvUwd+xvOXyHFWBp
dKOqKJGbiJSqCbfLGv+1jq1+leQLIjZXJtEaAw3eUeGwfAp+ZNXTpoTyMa26ZR2L
5/8xIgII7l9QdfcaakdkANxtyJX17aZi4JTnw4RrMlwybKc3dbUF30rHLEwwIHQ8
2GuuhRMg27h0Xu+XcYcXK7KiVP9F25s08T//oXcKIvBgGWE9VtyVulrbgEeCS/SC
ow2WoeF11P92/2ccmCO+52nJzYTJymZzfuGZ58HQkOwQWydrHnpLgNHXIPIZCgzd
JcutLNk2nvUYBnZz+d45XJoN745O9kFGRBV3FctdH+gS10XZM8FWV2h7xF6b9kDY
pM1u5pzwoiQiKIc9lO4tGH0ncAGKdh6Bkb5rkIRV78T42MeipMn32ShKXEyNt1d7
Uzxwi/zfRxSHMxgdUgIskXPuCejoDWIJgyZRzvpijvYTupzCq9WZREy6wg0obo5w
dTqF95JVay3zh48p/PpzEVI/EOamoAtP1mMgXNtkZZ5mKzc2/Ki3bgT4ki6LICie
dogC1rtY0njImVJwWi8UANzeFzAeti9cfV/gqdN/hxnQdny21ScL6gKlCTBAaJnW
wkVADvpByKGQIwYfIKJ3sx35li1ZmN59N4tTWRIXL6ZinKU+/yNbH7mWXWGsMmbL
JvVXYW+htkia9QTW4l9pj7wiDcVgW+rXaATyHZG3niwp2DAfPQyqWOcQcrBAc9QK
F25iow42of6OXTiQFKTZz3rfco6DYae4NMBIit4GSLlma+K5Wnj7vU/p4uZq+WD4
Ecmb3YOIc4dYMTFly1seNion4eRMZ0/Y+Q4YS0qKOVjDGPBH50FS1zu3b3ET1KE6
lJoGnkXLpV1dj/jsIysc+TA+41wXKmlmQr8QcegFXZ0lwMv3YT4+ZVVlxknl3Yem
Hy/jtvG9vVYmdbbv9/jDofIR2AgJDd8ZiAL9H4BvW9UOoutI/b6w076IaaDSxKBa
pk9nWADlspZ34yP1TV6tpH5/J6gn8pS4njboKx7QetAaVVeulzNRdWngEizJcSQB
+9CRGJ3xEzLM7NPJo4edZMl/q3nKEkhPGijyPB8otCXBFZVaHMcoZaQOJsc3n060
dgXMi35EgtCvmx+dpKFbJjY2AMGiX60EQx1kwDK9n+hySmGI0x41IUC+PK7H9kFF
b6oI5wWV7O0THZh+CZIEQWvsLwS1i8kIeIkJ/81WElb0/euxb+W9H75ZrbObzWMv
gwso2uF7o4hdVmUFdgs1lj+HQM06tzJ57mPeJtbaMbBC1rGb3JodMukmNatl77DA
cScuqh9l7U+2zdf/DkdzH+MvCqSEAhRbTRJxCSlrvo/tPi22e4gP25TxLLUOvLWQ
mjy1zYN4W/h8CPQoFiL5ijuKJvyyWeyNiU3LElG7GZ0kR8BpfVVSyO6XhQHIsH5w
mF3QNo/8qaVzez1QnXKo1lIKO4ryLgVqy+mSRUP9ijfUUpJl05ozFMQmXJlxuItL
ofKrQDVkQyN4UpCkIZV0OoSSuEdvR9shrtBRwVH/dWWtU7agaO83hSwBr3v49pRd
rdQ4NKGeKf07F7WYoVYi/9KClTPQo2JqYF4zXT9vQuePBYRJlOsO3i1COzQCmb37
cBCNuc9Y1RvQauC8sVeYy/5Up1cOjTagkbBiWmrFofkJcAq4h48+tlAyVDOYPl8A
6dHqgBBnn3PF1u83waERV+Io37FWwxuIkqoSvyV+brkdEQd23Sdv4wSEqMDfCbXD
y+aDcoOMtiWBEnX0jjj9zH+KhfmQMwkWtg24XYFAzLoWrooghhioQdmJ3wc/b6KK
VpVtI2db/2hwdnd84BEYpOoKbXddFCHUovxcSFhjxK0BrsQNqBfPxLv+k3cI9vMV
cE8cqcojPvruExJmXlOkenWktE1AuQzjwd1jjkx4gz8kdlc0yERnMNndDHkUuvM/
Z1Wa09i4M5d+ae9KlIzRrhJxk7s3BEBQXswUWAROc7iog5Z7yKai0WktYxFpEVBL
1taoTuR4jQdldFfqCqRYoGoQyWGinR440SpIFVMUh2yw3j24M6h9NZF/Meberc1+
lPiS0bfiqAQjqD0l/g75f59RH/TF1v7O3uLsYJABk7bN1L4nRWK4FRgnvdv4EIby
JLZaJH47L9xIUa0jX7vNFF6nqGt2i9XFqeh3/dJuqkjk+i2a2Aig+Zc/7bYnY/le
r0rHqt91kR0XFHGQy9CS2YwCv92vXbwJVw8xQiyOhG7oo7f8g+xtxMo4U7bnPMD0
y523+Mj/B5LWh1+LkTXDLCeccvL9WFzI9O2/CCZ+Ngxx825yzDkUfjPYLcbtsjlw
RQQaIuKgWzFBmZiwWcbOflgzLxZPMYl65BNm4hR1z8b1lL4qGHPTiKHB9V7k8Eif
ZMpMEFzbeF1l2aJQ62ITpc6rHU50K0wSn3wUpXtJUnKaYUC5C7/PtreyWLubMM82
Fi5+rw8g7JZgGkFA5Jv7Vbgjqb5I0iQ0XLglrE4X8mcs9kCVA6sSKZbu7g8S8XGl
O5ZJ3bv8cpNCgYFME5Wdi0tEqkO1lwdRyuXRnvPK3gIIaxR46b5yJ+/7ZVxk/2z1
dy8/+/3E28AFuJ6aSNzyWoFE+eaUJXSDSja46Us/0oLXvG2uutpENy8oOcWqSQ2H
DyUNu5ZtbKQZPblH2MhV5ZUH1oomo86vEJHifYai9vpjkXBz0hDm3HZNjf+o7tsx
1k4eYhZ0JLcEgDAOY4it3uYWXVZiq9oe0BJOFloqdJkXPflMEx5nfltVhhv45YC6
RrLWbD20ROQ6zr2Hkz+ItxtS+qYJQ/eLzNlG1zQ1NH5rnu7y+1wLcMvgcKBBAmCA
/KR/LPxUCzc9i5alUdP222Ymdr4kHtggIm44Bod9JAMLOJjw16nGVzCmN8lvSnAR
EeUOPFQpsJnGYcHDp9xYqxyzHjU+UO/FrGayKnBvMKosc/6k7SenLfeefmZD814+
COPSmchLFDXYGjd+lZ4LLSQWGupyiPDKhKyyXJ77sgk1nGQWTxQIv+ja+Tp3Ce7W
AmcHG77UqTzBDZPU4veSv4lGRq2D47LGMjAKiDhvYyt6UwOKXPbhLhX09za2el5P
tEmBYoCDW0caLcYuHjAf6zz0jpqVDD+EI0sld0k+lkT+moLn5f3Bdy723IrpCru+
FQg/sO02P4NKSitSQiEQdLzVXuBkstU2mLgkWpBVQprRXVTWXYsxq+qj1BLeZbTu
+zYiFDAmXOUQ0QAO0VxDBBqwrIb6u+RSnIvjcWyzyaoV8TiGntV0MtQxuqoQ4LK2
Jjj7jLKbyCw31UiAooT1DNQ02Zd8mHxw11SbHmv7aKMiKJhAnNwI6mz+kVjvmyUD
6TGaYDFKJnTgTMkVYRChvSgRbJcDOuxxe00/HrlR3Gb/h2FgEssc7ipBjd8KwquT
i53LxsN2g4S20TSAlCXJYlJctRaLnMTTbmE17e0ALjdBF9KCPB59dxF6Qywh0Kco
hQESZa63VEGI8xuJAGaKdi9vgGm3GAvu5WCZiNcY2MVl6WofjmdwJAqvYoEXEBmT
hvEQ5yQ8pIqws0DhHlAimSlN6TEWliXirb17NsUiDjriZjqTgku7K1m0xlIc/v8J
RdX2FWsT0FfdKBODU8gzUjJWzryRZ2JcqP9fiUL/esvhed1CpFyyG2I8BCNKPlv9
bLupJ5GYrV7Ixr5yv9J81LQnT6mXyUwQzu12NWmlD93Vmzpdlqbi4/l7uj7dw1/d
QexGtNJHL0QU07Gbf9NNj+gvqWaKKSUd+lBvkwgt6GEUAaTi4H2jBbUDDaaDbCT6
KBOXm0ZAvyYJN1ouOVMTujmZ03o2U/LChpyx36srE8LEeNSh6gmuR9r6q56wA6Io
qOWtmawZe0HJy7tMpH38hyqV8n591sxSt3B7B8NQ6H2KXBEUE/IX3ywLPmEvWfKp
ihRY80CFeDCobQ070/i9LqVbhLYlDX9TTWgZTh7KFhOm5rTtnb7vp0OlQP9nQ/1K
/cL8OpLFu8+HGBMsbWMU+W3melAjc+MIpFrpEMp2vQns7pM6VMaEcMpLt9H2ZAMq
QZL1vz1uk97Gg2Smvvy3YkzRFboi04ErT9O2Ienz8kwfPfAICunsPD8EOnZEPAlu
bHgM9JaVSyNK8f0AT23fEuzSNnIQPY3Bhw3jfDb8gWEMzS4IDD+Z0kWCaoDWp3ai
t4O7oJivHVR7oFAYGYj2gpCOh6ELrpayDu0gmnjyosRmt8rziYbsDrPt8/o15d9w
7tMGrv1uyQ9ELbbJQhn/2NIy0H7K/ofUymidpucR0s8YYm0uvSxMjvli1VY57/fM
RtX6cbd62QD3TMlIFX1DJU776v13k/KMrJqvWE9khb17QBtW1v6KDHnrbMjGknk0
6l19bIBgsWUK9lYMJFBzid85Oa6EtyFLMqQ3L7FqIz/Ym0jGuBZKDgGeYxqtmioM
JrxFFj6Hcsdzxak/8x7akCVXeabQLIj8BH2u5QxVd1jfVLQgMKrP/Qk7DFJFUjXT
`protect end_protected