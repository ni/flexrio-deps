`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 17440 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4sSkgcOrtFFGmnZEnVbxgx
+l/NC0KUoptgPj67g1Rb62rm+Mdg2aVlB1oS69loY0RNxWU3LIfsk2RA4un0j0kS
Nt9naSVOMHkKPNY5IKoU992LMCqx+1+rej6ObGt818gGR0cXjl/XPQTf6xYSTDta
EJfwQwlM9fM5cmNWATRjtFDMIkY8FqO+P8aRV4hCv1fvMf2RR/rSTSog7joRA2wr
7sBQP+N86Az3RIyWtZ4D8UDJ3Yb3mqLjMa5bhkh8+VheRiHKswJ3yfLsgStB//6p
WKrMnJxawfax/MGr1xPQmWbDmQZnOt/u1XCofqWdKrfyz04UP2sztFJyDftJHhfr
HgjPm4ZHsjG1IMcW4qQ1gKIGWScsxCLnTM4xpVFwcvTLAGAUtqjePjhVG+GqrPcX
zT1I0Q5HCDp4ikI/MMSAbN9+4q+oMbBH9B+iecZRZjBx5ClHWjTvN8dJQWl5SJhB
r+zmaLbQgKsP1sDvRNj9J0QjtQaPkiWOdfLaDQcwrS+d7RbrcMuS8Nq9CDVg4qfz
OY8sohY39kT20JHpnIPeiAxpv8TM8PZMiXzqolACX01/1roNbbbBaAlC3Rd04AdG
h2GE4PaO6Vy0Wtw8XZWzz83cSKyzilsQgVuNCUJ2k1oAojColnBc2QHmiXqrK8oo
P99Wxkvi8TkHvyggicygbn5G7yj44X3iPj3DmlArb8OIeFbT1xa3Oz+BdJmiE6ya
uDFRj/4WjdIKbB3OVulSncxifPBGT8sj+1Byxrng5UsZKwDNRQ4BHdNt1oeFHE6o
vOoE+V9uzeXARTS0nKaVlnbpLq0IwFs9CXIMsDWyfx2iWjeRvJ2vvOT3eT7Au35P
/Zx920QqM8VEwkccZIbdXQwXVQvKpc7iG0pU9m9hRSmr5f2Hh6I47f3czdYPJVQo
TTxpyZcJ3AbUK8G6WnGOwNZ34OytYd6hWqlx3UNtHz53bR8/BtsG4yy4/MnmxjVW
UwFAq0RPkogwPjEPU6dmWOy6mjRJFKgj0oRVU5bZpKfPr8vHTiCcBZ97XplDbbWQ
o9oxVtC4oGcIIDaE+qabqsBLynncDZM9jNVoHGNxllFcKeBnMfY/30Ps+fjXProL
9idtXJgjCyCp/gWBcSHxbn5P4YF7MoT0mC9lu7NQjor8DYBuRhoPwXKNDA40QYxR
m8RkJVQ/KH6wiragc20EaeQyMAT7x5IlsDtDRqbSRFzjMmWAWVzn3HVAol9Hyben
3+6Z3tKcpRtvL849UF9Otabvkoxdcz8tt957xm0SofZjkJTeuFvwnJnAfh5Z0T5l
Ka86UloOgSqtgMQToIuQRORuP1qpNf3mS47nHYSbZnaNUwu8ln7ncVaFZFWq4HUS
vAxmp5wnh31sf70rGjmLNIUJA3B9oF0cysilnegGHt8ico4TZjZGhsMd5hRR0nyC
uLaErx+gyDzTjomI7yF04wtv+MuWbZReDCQLCoV7W6+toi+U+wr2quv29B9owm1k
zgH60QjBPUA2boPU5ga3hitGwTrWiobLVCqyVXfCecdrKwqbeJZMopSQ3PzrHX+y
bwQtiFoteKcavYqu57jVFkHuK+MVtQF+9IqD3UwK0KJoICu1E8S0YfuEw63Yrd7S
D7yzAAVSElIcTxPV789fFrmEa3WAt+gmeoJwDe4HnTqw1vu/7IvNN4QdO/9E4Qtz
QksdRII8rGx4chhkeobqkfLr3HH3Klwsk0Kcfk3DeuFEYdtKrWhywkBdA8DBE1yT
FzR488Ym0ct7zpNzO/vMGA6IkztpbrW8fdUP6d8KfyI19I8/zAWr5SLUWK604p/p
pkbvu8Z7E/JpRJCjqfwzqO6PV8SAnsCcEQRnGeepZPqS2F3wDJClQpUeZ2qH9faW
SmpCiy3Ui282aJ+bb/a/CVh8Avb2dwPbTpvn49Tfih1wsTlc1yY9NohdgOeKftQ9
/SfBCWnReHlX/foZTSusmU783wV+mPweYxV9GqEwlfCoLR9xvosImGK6zy8Ph6Au
ss+Za5WXHuLimb+oTlMtEIQ1uhjWppYv7NBUIb5Bq1sZHuOPHTOPKcdQppFnW3W3
a89Fr+swYcXhoKvP+/oSf+XlUQqnxVzLSqlIPwhr3hy+4UPAIvn2G+Km4jQoDKfi
Fb6UgoWCtX7fE0MSh6IqQotj9+6irGoKBWs21NUQOnPwe1ZMxmmzoqDUwZOEXhNx
stAB5a+sChEhe2fXlCl8/szVrv8bcBu86Q+wWCn+mN+ui/lAFyR8lQ08SNdtU63p
ufnhESZBYMrFKxHu8PFYr2Rs5tv/tF05QTGDE3Jl+BCta3o5RrN9kn4KiGjOwGfU
X8QaG7IZd944wKqbaJo5FwOGyqE96TWWPrBA3ZrZoOTdYGzZXf47FGH0fNGGZHbC
1o47xBthHuf96q3x5TbFrCH4QX2gZYukB8D6VS2hflUChM7ktpjRx04o98l3x7kH
joGbELpCCK0BGTq3sv5NcYVN2m/+gkC9k+PnNkZ3NnS3lFJTGwnw3mH8ML0sRRaO
w3M/ZJFuF4DyWxX1hZEfiqyafdN3betSOL7/9FPeF0PB8hlvFJogaTkP/jqqUeb8
SwrSRrOSwvhcnl0sAAFzn2dl38wUAxNf9t0RlOcVj9IUYh4YBfz4lShIrKVpjEgP
zjC9agYvaLXsHS+TBHyxqHd7+sGsV4Uc7naZgjEQ5MKWaW1RD+dTi/k1dOKc/qR5
1GuBajazNWUdF8kmgn3oLKdh0z9oNL4dKDMyHkj1yl81X5Qd8+nhZT4WPWqoplTP
zFr0X3poV4h6rBuw6UydmaPoRECFR/b7h+Be780jHRodn3vG35VDW/630a30U8C5
53LPvY4LJWodEv34MJZ6xRqGT14asOAwklyPxxfj9Z8qbJzXr3Kr5DHDAhlKzOor
49klSv49EW6s3qGFblvIK2yivIUyB0v1kqzNNUv1rqUjjG1O4nUrmdmOYksG2KF2
oVtJeQmoexw4+tuw+VoroQR2pLZwHBNMic21nLk+XZOZRWeducKkhBe0X2043Pms
f0yFuSmacueNQqkfsH6n9SxsYYB485D6C9nzht7AENyApAr3mrdLd7KiFzHl0aXZ
Dhm9AWsM4nFFgaJN8Me+A1haygKqbrmGEucSvAz0IF87z4e9P0RJWegFe83eGW1J
U1J8OengMmKuQwHTq5zop4aVeAQLNm7fECCYCizHzFfPjMs/e2601dDasBFtIxWo
kpjy6SFEpsF8N5djJPyLp1RESx1DupP0FGVGf/gkoY7vFyK8JplneUOhngJcFp6q
+yAA3PcVOMJsb5m0bRmt673IzF4yjhhH1j1g7jy7iTDtwpolrBdig0oZ46z+s25k
gXpWkNNv+dxyM4VwO/bPgqRCXFr4IwiqUYbFDLWuPeRC+2/BagCZKW4cn4Ahc0so
O+81oXMFx6W6z+j4KjUwV9fzALGgk/wSFEYelWwgBiuUMXa7FEO/RsT7z70VIAQz
8sqWE1XPJkYiRT7rzWdTZeKavsOBY9nkPnU61FmhYKqONppQ4PLm89rCEW9q89hv
wlbCP9nPmWAuPCqzFAuOZtHzIEc6SRmaFysOC8V19/5/4YFne/IEBupJ5bsJ5HFO
/pssI7DgN8naiwp5tLS0os4puaG1bjTXkUWQUm5zIY3C1gvZNkEAn7/daSBxPyC8
X2Ue0FH9Dg+uIWF11n6Meern9NAYFFSvDR2BAuKSOtVAs4VJEIsI2vVhkkuV9MFV
VmGOCQJaFGhDvTXDynaCab00UGs+Q1PMxDEmpBs/7DG7JYRbhfcysclHyuU4UiqA
mwigEApAEAOk/2Lj6fmvKbPv5J1NHRYNZjgo9FrGQ7SBVySRGVES6ZqYzqcyq2dw
bzE8eqc1hgg796zJQH8YWw/GwhZ25A0LvmlfFeisbn8UsQkYxHAKW/A7eUzwZ0cd
fZf4R5trWKXRsGKNzc1P5Bv8AcHG4N5Un4AFv9NgFUpJ4pFQuHt5gt8afZbCc5Iy
lGuu+Q1LE8Ff5xjugjzlh9sKSd7NOyTvfhg0OcT4zNORkVq90pOdmZhf3rdjwnMF
UvrziUQL4N41fZ6ESEFmVpBfzk6WVloXIL+8AhV0xcoJ3VEeaLMVh3AV0WsOHzpz
TLsnW7k7o4jBP/WCtpqhbWZ0xBiE/cxNaNKqnqAzt7npBBoT64eC7CC1X+OKu7wb
M2khBi5gzybJyeHeZweEgabycUJVjZRDX4clK1GR5h6/N0NjZSiQsGu5YBB8WIlg
+Zagcub677GIiIJmBWXBLbfHMNuINNg7u4RHkR23urX2npmQmV0UU1jR5IgvobpU
/EIad0RGgx26QwqNgI1F5kOLhYMfIpq45TpuXS40kHanYIOlH/7/AvAVza83jDux
xJXEuvXDrn0kD+5+3ybrGdSegL5ZhF+jYw89vm/xujyZN2tdmFXdJbDGEn5ohjPg
ke74q7tYkrDd3yRs0EFABXfVCB7BXJo+SzreOr8pyZRT5ITyjK4EjhiYOw07aa6T
aq8p66u4vrFpA3v+8ml/LQ/2QAtleRpvn2ZN1Ook374oYygrYAYcRKau0BZE9PYw
slcNm17S0wVES993MT5RM2U6/nXJFzyRW6nTIbh2ABihroFRQ2aGXds8Tkdhm3DO
HF2PP1fcQGuph8gjZr/f3qDIFf42aH0SiWcKKZU7MhvrWJSGeRsFjgh0bQ+PFYf+
Fa5aZauS/DgKKG3Grtvz3j3Aw0GlEc+S8LZ0wpoIyQwhBjZsYN4ng0oo2JqcQCpZ
s5zAjp/WKobiIjUpQn3GexzMS3KAcIgxqbQRSniEsc3jaH8WBIYJl5JbtIN6UDir
YQ6btxpp17OiPeQEngASgP+K55uW0y7VLHsW6pNx0I+f60ZLDh1R5NUBrc2tsPwD
Trav25ihXM6DqCgjF1ibHn8zU3u/okMMw43uUecWfgf/VjYWb1yBPCwwrA12KZi7
yWTgNIVQ1lOEghcnKf16XagN+kkEXAWdB6nNGgc5IhZ/fe/pqVpmQXO4jaGtWUhw
W6Dvb4MZbCDsX5hEoK0qXf6vV5C1vn/fZVn4YdFayYdS2pTd74kZT0fJnfGbW4dK
lNZQkfk3LxsOxlWiv3qoswjgJ15Y3xUolMQCanAHJqdvomCJ8Gt/BkTWeXEsWPh9
80ot//hX2v7D12ZLnxDyGHaP/txzWbqcUfwPobigg2C8UdW0Mt4bSoQb0O1EiQcb
X0myDZJtN1H/Gl2b0+Cvs68lsQP+eREbfNS/5o4gcDQlP57wztvwj4mXphZXC7nt
VMZzFfzB18aH78G68vRpVZ//LtQQtpRe9rDFPQyuSK+KgzFCjhzGTaekJQcxnOEW
YGP2X2OLnLDarfHHCX/+eLUwQNcegsqJw0D1DfvrTg7CX54V4EleTsEklDSN3efO
UNMaeXpUav9A2xxX5+UmW8k7KoC1C+1zfqt5NHvbw/OoOxq45xsNyE8bBLKIKprm
Su4yvzd5RTW2VsZVxkt1jH+M9gXxurM4hP5rguwlLHnOZcgtKyEebnPw2HmFhaYQ
F7M+dZ68JS9fnjM6qP1TWlkOIIPp1roQVJMD1pCBiNQs69YZPtJpQKP1WX/Bv/Ms
bxOjQGTzcTG6Ysq05lY2CJqVPLPH4bmOAM2eJMtmv8BL2gzkH7/bRUnuuB3dUV8X
/CFsh4+wJ1JJP2SiYTsPIwUJWwMQMFIdOwwfOm01Hnwd3TrpKcoB3ZlM00uv9bYm
AmPcLsfplI9oAHT91Oqx4mjNA70wSShd0DURFIWwgPs9cQvRIyTTQ+1xFU0uYydL
93+eFKO/Snk+ILKJ4E/7RYDq5Bs/pGkFLy+8d2XT0dokxED1vOMVlCX+yPdmi5ag
+D9oI9OjBp4tnXzS4gG/IlqQNB2NAeciZTlG05SUokp0DYmLFFENMnrsXctRfH/t
voNmo40meY0bKef29i+/sDVbwrBFCtzhygOxp/baQ9jn9ig2Kr5a+vwZ34JNYb6b
P7ToMAhH7FMzW/ETY5+EH3tjGRhHUQSn1l/8dkUBHjMbW8pMw3NV+QNWl6TNwY33
pUrNNYWtsfGO068cMr5eRAkjtqrDtkEZRczaz0X2ESbQbrR/DlXD0IzYTQQf51ZL
4ydi6dHzK8bBCDY2RhrFcD0nuwfPCyqiEVKCgBfcvP14RkZWsnE9EjYWrS/08vdv
A5DCTEuno5cb7WqoWQH+XWS+HWNQO/nuqAKDWRAi68LIiqZC5HgRaku+Oecxfcp6
AsApOyDCiZpelUzM0P+uFhoUS+FaVewvBN8aVzkIVRsHQGpHdEL9C/p3ak3iqCwG
d+11BXZ8rDgvlk0biKjSevZMScI9jmb+vehFUSj0DiwTfTeZz0r+SJe+TmPX5RjC
KoatKG3DSfyIN6dt3UC6SDuG9U1//6++H3oNLF5UOl3xVBIQzdy4qG8JojrGD8XR
IHm+9PJcFYcn7uJN6XUd47Yjh9532occ+BXaJNMNk9mcR++e+y0rAeb3j8uP7kYh
OjIOoCyEoNKNYiFjsTGr4Cbdqhk0P19uObuP5d/ZWnQFr5W1oARU86t6dVSVRlli
puwwAgDhnSB1GVT8DYDJo5sxendwDloBdPf1z4HzxrJy6HgO4jf8X86EDgEol2qG
ayXOCzUCVCH+xAg0vMRjzsuwjGLEi43pO7w93pAWtBQ9In4b5YxuI8ZsbIaWqGXY
CCkF7CDGR42mA730GcC4mS0iKfLIVV6zKfB8oJBov8JVe6gsUW5vrtktgEzEr3/y
HT/QeDHF7PYQJp2xRSnM2w1gbxWn7C60frqfNqQpvtOZafEeMuk71uPuLKxtwLUO
yKINLTw4rrrrNd27lV7eCA4J/YSaPohTFgTmyCXgLicOHeFenohqWP7CHlE0ptC8
cwMe6k7BvfvBsWMDOcn6q9VFfCb+D1g5cnSmd0XSrwqWp8i3dagYNtgbRGm0X87p
wmAJAPO0ZcsoT4sYPCAfMq+1Rm0JYbKVIiD2LgioqP69sw1/abBkNlXcK3KUFjU7
rlP/ZWxYEY7VQWj1FcnpMq7f/SUScQoTz7mfa/hp4kI7wMZrnosUl6jpT7CqXRQa
Q3Q7Lcxk6Pe+pBee6XbyPV4JEKBDg2cTFl0xWJ89N9GOnZ0B+Gk+cYUIX6qMSTmX
OYq1sISatAh7SxKMjodJUJg73Y9R5No8mmSogHyLWCtv6tjrw/8rjTtkzNjOaiRv
gDo3Wn3Evm8rwWG4SBRr0LAWEccioHt+bK4dKCIePvOba0OGdz6TFhKcf5diPcBd
kb1bVR3wb1swkOkUmP/lw5jskbf8D5haAUzZ0tePC5rf6vwT1OS61lmw5072R8yA
pLnVhetO8LPPZqnLSVEuqsbTpkifcLGJVtWyNtrijbu5QLwShxE4atPFsXvTvfAL
coI0O7HMb9PmhIacCL9KXGgFvEvLIIhMI/c9/c5G6DzF3avsm1Od0OsC1KBkmvaR
E+6+TP7QxTDXjx6i+QwmTOC1/OVeK7I3wsL+LWN02qCZxj2iaeu0ctGn4sC+K2zR
mtyIq9TSED3txhIkQFwJB7cWk+P5+cbDP7z+NYp6baxoWv59SdPUQEy+k0/obgcu
fnnVS6OYdAvgN8wyTjwPHTahLAPMWWo0zj6LpduRZfEtY8J3mV7R2q3pzbD8edoS
9COHDLQsSYUKnZIYzRVjzOrzv1qi0jQwQQ+agKxfl5n8/8nZZAePyGrGbqh8/HZK
8cF02zp/bFtCwY8Ih8VT5OzRDTICzJUOAlNSXN7dWE6Hs0YIprCIWRtqfojElhto
dRcb4eVIU69IlT8FuGWE0nhHPF7zW9KobMnz/XQzX8/9mgaAYxelrAQS1zPgKfL7
ucohk25U0o4uFhLXWcMAYmiQf8e00qWzpU63n9RPeww0DJp5XvtlgfKJqeF4Y/pd
21Mi0EaevjkdUFPCKo1/izIw0CDDX+wM2fD8rJnBXIgyS1JNO2lv+dQJMv7Zxc5j
Se7xsVWMyjRIx+FOeE/ShzkTiffs1tjKNuGS2YKiIIbBUQi1YqSSMZa1v7OmSBOP
rMkEIjnGk2YseUeUwaZ1yYwE0egU7VvtLqIrpWfJipsuuKvVrhiGq6yXcbmG0UOc
NBpkoJMufrQA0/Ib3dNAaRyC6cnoQ022vSzZhq3YF33wiAKcQTVDhIdi/WpE+d94
qv4Yq6uY7jdvMVE2Gjx7omBQ5whX92q4eCwphpQxbTKcks2D+75SVsvPr34Ed6Kd
y1GDKl+uUfQV4jSCX8FMHfViVBkY+Skya12jwLp3ZKnNKEV48TAsGgbvt1aOozmi
cZcJuBFoftxkA3Y5YBc3cywxvKzC/vBnfA/BGjLULPATlUqLFegnO4dkkSfHzE0v
0KEQ46x5CFeKv4pS2YLS6aXTwB+nX+8Hcw/fDig0aDr6VjWFPt9qj6b6t5eu0TVQ
qnZ5s9PozD7tk7ISvrspg0dJzD9u40izsXD4RQFhYxVWPX7Krmh2QGjySS0Ok0LS
omMPSaY0wehQry+g1KOQlyUyqo6EeaN/g4Qz7k9b6BOZkLt6LleDyrNBgF0BoTEZ
Ha+9zy6GB74tN5h7VNbri5Zg3So5zVBuc64A39HnZ+699LkcldGByeiGhVdUD6Q0
GhJ+RxUPay7K3CYAy6r+FK1jfovrjrjkrUFabUArrwR3rz/HyCKe7XlnrSlOp9e5
z13RECZOhpfACYZ5pjGhTi2K+/XUd/9bEym7SN1+jTLuSuMP+iwxuAAm+tIzE/1q
jz5IRM31aVuMenxPSxinPkfkZCoSoBEQhOErDZw1/VhyJhBMS5JHQN9DBF59Qwmq
OUnHobNfdGO5HwPwMuqMX8cL10BsVyV6GcGfc49rZtV/kpAKbbr2uXQ+t2au4dll
8OxyRrR/ibFl97dDWV0BedCgIE4tlM2n3ukV2asT9zJAwo5KFQeeEiRKCqMnR78I
D3q5k0tgCpVLoQtGVgj1YqIZOWoVaxKryNLJhbeJ4iWCmvU8xHmkECAv/akvpoB5
Xtp61o0BKLPu4DnSaiG8osqjyE6Rd6TEthVhtaj1/UOejrFRXGkvnFbMLCXlGrde
IkLTw+7fEL/gYTLZKhn6fBj0StDjeXengQxKpo5TvVbzUN5ZfMyt51r0bEN3DhES
gwRZnuxBq+YMJY0canqL02qHq9vDD8IvF2N1ny8swPnAwmKeo7Qeo0xhmQ4qZAJI
X25lQlAYJ5taTK0soirKMKO54l2k0RR2wpX3fSBMCqOnXzXNnwsfW7Fbb6FamnWt
4B6YsGaLUNHe3dEoO0xGCnQFJkhwlmuUEzAmvPhvsWTjDBtBZ10LJeRM+KYWCQWV
P9utYW7lIrcQ+aHSLAd64MDfUzL9sSI9+z98JIY0/l0WH6OVEMWFYeFBE7RA0X0e
IK3nW1s9f7kcHprmC/NOVb+z3veIAlrNnXVcm9DSHDMvqwxMNh9IZ2H3DsSi3vPf
NZ1uP303WZ06ok3vAPVoEcVUFfcWNdm9UM4BuWibh+XZvMwQiDhW0H5RrcyDVffN
pHTwyrgq8ZXcZ5e8h0nVhaw3+BIRPiLseXkmMqbPSa32DW0bz9WaM3hmrFe3hSY8
XCmGY7547EHIxBsfjy37fTkeCH1FFoO3h7r5/uAbTrXwYbSYj0pyoLPPBCaU/KYH
jDmmxJ1ig8D9v/yYmTrDxsTBBzJdie6fkh/cUx0N3XAPzFYsMH/pjZ00hnuH524m
jAf9WDUnA3HEMgRNIsKUC32G7LgYrmYdmx28AxxuBvVD5jVC9mA1w8ehA9e7tWId
G/e6GpC3VuO05JyK9cXurjrxLcJhNaPNk09RDt4ubjIfMAKFGjjyiY93oB010116
STTm2d0nRgvEPpzkU8FEpJZUaTuWzZnXasPUelnzZ39m7ShgmR96MBnMgvjsFzPj
TwjZKYZNqA+EBqv23xf8kLlm6XNKZUu1Ujxr/qBbja8h5CvVTtrI/dwGtvqHfh90
FK/JPnrZIn7WXh+kmxTvxXaACHyQdOJZlPY3F2DrQGgW8sF/MEAii/OvpTVIbtN3
5Dp6FGK2aINYVFJJ/fjjnyzJrg7dEwZ15hfe7qtpextAorAf8F34CWfvqkWI9tkZ
7B+qlyQ+SQ4F4urzQ0OFY9JOciJyNWaOxfInWitzPy/1HxoOOakJ/719Np6ztMOY
ET+VSBaW9Bh6LJnCVNYbpFhQbslHEjbgOTNvVpxDrWTByoFgBnABi5yvmPDYtIdN
LZam+15rDe6HwA07m9SPqqDwXMKSRdMqsbTS2k6WytgYkbNc9wKPKtRNRsCKNusV
bdHZoYzd4QB9qd2WB6pcSLnxzxBbMPfu2xZof+8mn6dbJDuiewD0J/IMgYX18ltX
RqLFOEeve0YtzxEZOO7J5gPUZCFWBXIQWJ4hioD+t3GhSZxhSl7xotTSr/LeNA/q
I/0atRBRennvm+nAMf7ECFMcXeTMjj+Ou8wLPZIAFy0vfzVMhL+xTfGe3LImPphL
R+/v4tM9PEqYUvoHXb5CoIBvjQ/mHKBmZCZy2BYmIi5irJM7UuddaTQjCCPqOba6
uUwb6SPOyM3h4yKLUPKl5fV7AVsm8OhBLddr4+r5MTeQv1LjWHPpO+m0ZVjYj4uz
SgXOjH31cvvMJp8Rq8DVMboyc0KVUvA0xdH7jbWRA6VSiyjBeTPJ0opGFSsaC0eL
QbBkWxrydimiVOlFg0RHFSmhNcVHwTUiK+u0p4+W81CLt462EK0wv35hA1RT9QF2
tpAWXb5ITBnIlJdW2fadWtXSeHgC7MEBkPOf9Baarma+erNZaM/ntD7FHkgiG/39
uzM0sT1BO5EhlMOSvNCk/QTUwR5yR3u/yCW8nmvYd2mURhEhIagjrr9cD2pgKnWw
z20TKyTyb+B0kn41nybZfqzvSVoSY9M38uWMVn/kxixSUP0YOC+kDRf68N9ogpWt
49aRGHKQgh0Oa3p80X6J5zIj7uZQDG3e3BCt377C0rg+ub1NShld09fFx3wILGZr
m/8MpRqUzace4wLEnu2hwH9nDof7kRcs6BlEbEVtBunhxTGCM2vA4DwNfb84YDFp
BOTd6thc7OTEqdldMcJhv4aH3CNhJ8UpNxTfbt9AqdME80IudBtu0dhnC2aqHOrv
mJD6Pu4IOYfiPGkZP3qkXChJRwET6zHtgamwpEgT2vborYuS0EQrpVY8bZTqcpRy
oFx4gZ+cPXuUzj+z8sVOb7+zINh4qPeA/qCIge0aTL49znVZvkFYH1cvIGCGROAM
msgmnZcYa1OMH7LmeAcsWYf1M7ym+CC7kz4Bq/RNjD0Ryg7YkqcKgbqfoWaqclCv
9eP/u6ZxbQ+dew941vOdqLePLsyKroDQAvOfYlaDA5EdgFSnRq2E1oV/9kMhYJ+3
v9M0k6D0XHdUp4whxxeLcTmbG9C3mL37Db78QYVYw7ONtjDIsY17FOjTtIIwwTI4
F7J3WfnP9ItdiLNvWp8+c5VfGmzQtIqiom1WdktmnmhDiUEyVt2J1cScOu7h289D
ad4rWOvKnB3EV/edlGD6GaEiJrO/hKo4qkKQaVh5WhslLRUu0K9chJBMUc11pHK7
dgObrixCvoNTqaplzkmKdn0RM+Ib7v7SKCmgCVmw6ggcai/j3nwKWmZTmmodZ9rH
rU7Xp1O3ZHASK3sFVV4ag2TrJ0EObC2dHOviq7IXWCJAxjTIRVg/ZopmbeeIig8E
dw6YMRoyvdQ/ReUBRF61Lth2/MnsPDoJvdfaTFsOK0ubrBj6pwCcEVBrT8U4AKwS
ASmzuvhXVVL59NFcUa74xpmvfmpvxwRTB5yK600pYuqxzFU0zVE6gzsFdkovPXdM
M85XUILeVqkaZtl7iBeUW5i4EdHoFbQtPO2Gs226Ezcv1Dr/hJB84SKEyKJFnJiR
emuUy+DJ6abBUDpgENdFKdmFsNEH6cnjY+llPn9kadHXE9mCNUclOwXQu19OFQ9i
eSHiLiUZIamQGd+l9bJ+TOe3TghPy6sF/l3SJWm6vAgGnQ69hxui8d7kJbqBo9AM
aYZdFpFOUsp9OEDAruU57OMtQaL1kWvUGrIRJ9HfN5LUgkeQsWYmbF9kn1UaEUFm
nC3iyBu/WBYRcVdGvbfP4TWueqtwM3t6D6pZWRCoLgrkY1RnhQqtebMdsnA4g9Lp
0AJgM2DUcdp38BhLFXVpYzMmV6MABgQZUcTKyTWm7Rw43SVfz80rUqRLxaSJSml1
/eTK2pE6906vN5yOttQ/pX9g2xaowyZubphTewn6dYRdbUul45m6W5qbvZBScdqn
N4E+A2gFafn7qn1Cg9eIik00eESOypFXnEE3d68N2qAI364soXpQLelaWkLabx21
TkN3EGOLytBV6BSAJdVyyReLhRd5Hd3dsmOKpz73hll+UK/DAmTK/pX3257Uo+f5
7yiejUC7nEayBTcm4NieAFNaEyJ2LAoF/JGIE7GaEWvw806phzsNTsZkpA1NpIPU
OtxiMAz7JGj82Ww6goDEpmgV/CXjrDZSqZVWfNVndecSlJdLdbrv+BzgYMEVPYI7
AHMVWYKJcG34bywMddgEa913D2ZQpuL4mBEtg4XBxAyh+hB+FHR16wmfCt+hcSrb
cTgvksNsx+OXco5QWHhwWibPW/EAjK5nynVhuxxR2WAQN+/olFOmgWhK/Nh9CLXZ
1o9KkwVQ/QRFO1xeSs7NRfmu+v0SH/sHWzE6yB2l+gAKd8XFsI2Q3f52bzaX80K6
bcbyzCABbyBggxdHGPmVC4yURlttsYQ6vJ/coj/kYI+dzRdx8vy0qWNKqkbgfVL2
jHGpbTfjeXMVc5ZcIICIeegwKLDM9WC/T6XV/I3nUX8FmfzHb/bikGSQpbKKcUta
Lswqfj2APR5ZzV+wIvp6Bq57NJ/nDoAfYun5XPz087U/zcE9QZsvYMunpRQR4o6J
CfEzKim0/xouJOClzJss9ACIYpKSqwCMOwcHThKicvaBhZj+6ygOIFV/q2JW/PKu
a92iAzq1MN6YM3L2NhR4W0lY05v2UiKh1et8No3L6ack9N7ZdoV2JgLNKpPfws1f
LKLET0PVxVBoqbSHJLo++dP3UfhMRF1+paGdOyzNq1JmZ22vgLGDroJLNU92zjkw
tM4WU9hzFvi0uzk00BC/jdXS31ACwDAATKmP2ICGidw3M+PGoYhLwPwmpOfsHm86
3GKwv5iPzMbMaMg5CGSfSWtUaR2EeZqTaz2ZsKXRnxkqTkjgrgI5PFYEjjGu4Aa2
uC8ePk01RrkHlBXsOp/DsVJePhu87i3cW9+FLUlSHkVimnsaeUiUb61L2eudpzHh
YP7mYzIhfT/3iJ1kdUkg6jzl9QBOvJaqFPtFZmtuYZLzevSIkxngD5cHgeDXcd/v
svN0BNDMsdVvNDhaO+F446cmMyGdGlG7cFCEUxLFplcoygqvY2QtDBaVZm1kOS/q
IW0iVN8DgI98/CggiUgcB+y8RNBwzcEQqRHWcrsI4BYdvw57F7weD8jRqdS+ZiPz
fhKTFXy08gc/HL3G8VDrqqYYwzqpkxCtfXOzSYsv2eHH5Ee9YKeNZDxUIWOZMJG0
btpsFp0FmTAvmGURX9E7QLmEmXuukcFNj8HDCX+wFQ9A/i87IQPf+7tQfBC4MsS/
Wa9wqwY0/d3n4vNjsmZeCAQmujxu2FqfeJ+3ApqEPc8fXdlWI40wOfGGQX9Wea1N
xGT0zH7sAUTYLGOL22nguw1MU8e+Py1p9AVclpnmRebxWJqCeOVzqDN8nPqvvi/3
8v7qBBK59honUdJHE/jFsOcXj9Nt/pDWqp1hAP29QwRbsfASaeZTiYhMyEIrgP2E
vYgAhRRrTaUSQc7UbK9Ccc6v5PJJB847UMJJa8aeoUh/3gCiPSW2+Nl4/7fZzca+
ZaQS1e0IeNIQjrdhF1ZE3nJrsfDnhFSvSO1A4JDmjy5xAHosobNAJmeBc29QlP01
7R2GNtVeHB6WPiCUhKsw9mo1KveRCt12j5J+kSl5CGm7GeQ+uc4lix2m00EIv83M
pce2YDukfvDX5IZc5U3Zc4MsMm3w0hzEoMAW4rcnMLyTf6TCe7u0DCfS/sh+SC7/
MPK9I86BIzXrud/1Pv8Tb8/59Yx/2jgTUBI55vY78Haqx6OKFU4csZOU0+sudyJ8
b2/4NTLSgWFOZq396r6zUa33j92MEjGFb/U6b9dynhCgboKLG5Jsal1PV+RfmX+H
9WRuy0sZbNU3z6L2lFVOt/0ZjYoSmd54EENeeZbYfOIEFxGYuIjPkJCvkZ6AltPW
t7LhwvVBE4wM+ja9HLiQ1yCt6iLybnX6bcMh3WP2Nd5QaE+9yCtQSkcGUiL8Z6iA
d+hwY4D1sFF+xgXmhZiP66c/GiCgLbxnoIERdPgEZ9vf1R0geTxlYFSCSOQkDtYY
08ASucnPRyPDcNawwVU1hHx6t6VswcYNpQGcUCw17LDOq0rmCnmM7Ex/2aC+Xy1V
6CCeCJhae4pzCqTjjbTlB9m8ozxXCIr7lI7BZSjogkbFiJo2HzB7YUeHtHL0A7RE
th+eslpdzk5b1HjOvNXyuNhdPTL76eaH6hWXr5jRUVFl1OivMvnG8Lz8cYWEFpJ9
7UE5VAq63yCSQMfv2hliS3h6kxhFe7mUTopcxx+PAI+BU45HRTPNa6BVeQPEcrTE
w02QOu1qfvEFI8K2Afg6Jy6ReIJz7bHF6QsFFu9biyqoDrhbdgn+I/t0tzR+8YGc
PR1290L+y/RMd9Qga57NJyj9Pgi7gSButFHMi1HIUELj/hjZJ6JIH8svUwM1UQWU
htle0nLgmasd8JOZ6TrQ3D5fG88gf9sePIq5TDZPLPND7e9VQCE0RuISWmwdweEq
rupGlfJ4l9+Vgta2FdwMQ+fWkbHtI+QPx2jjmeFWaXi8Za65pOhzSfoFsM8All4P
GGr4jCbPXIBa/S1QqpNIqRKpBwJ9Nvv0soxn4gTNYaW4DSrUMC0x1Xw36z4yY6AQ
vv+YpPYWee5h2CKgJcHU318tA9BjeKm0qktliCqkhy9IzQ/mcdRLTiMkSD52GOss
66ZvUlFD2Qx6UzJI8LcqM1FCPDXl7z8xC00MemmHXsssPEzw6iXiTQMAYyMkYK4Q
7XJ8bu6Zjn0fKUNysXDfYlvwb+EschLwIyLBha/taufcNFjsSaHQF3hlCWzwA4WS
KmMhrlekwv29o4GDctGBF3KvEIfZcWpm5HjY3lqaZpoaONAufr6npUgH2Mu3K8Rx
OZGEA6QL4AGTf/dnVMjvihJrrE3+0xgk2BDmgAdq0B4ijDMMutz6MVYvE8wJIuQ/
GL989jjJdtGSMrPuVYV6TCNVI6L9iVlqLfe1StMX+GWHA6rfdej9WcSX5HbRLvT/
634mYU7lQ16kyYzgTP//90MVL+lP8Hdq88hUZKpjxBHgO5KoZmtWmkgEQaM2q4IW
8OsPjAXRy6CbP/SPZr1340EfrGlVtHYUAn3X5HkOBoxhhnk0XrpXP0h9X4pWeNUM
i1ILv40biKI/DVgIHQSDqYK4yLR6aTTZnkK0xszRfMqpJ78j0yZSSkwMJSGa509/
M+mPWuWG4CG+FiNO95Jwo7YmUbN9PwwNOO9yfMCy3EYpzUOd5C4NmZ5Jzqe0PhHE
iE+N8RHIrnlNTq+f/nGdiKFMJ3KzWDAJ+BXcvbTe7BskwhRbOKZWPr8GkVq5Gjyc
xxYp6WX1oIvuiqRLZJ3kgVdAt75spVkrKbW1ABeAISYOiPXsSr2qAhwwlpyHGGS1
wM+s1egbt/cYArhRhW2oNjjXLWlJoppsH9g3vU+3l1hnSmR9Dd8CqLRaneTt3lll
3FMQjNeR0Ba2FQX6ACP5bmHdfbDOdT2HghIXgnsMJ4Cy3JsFZ7lXS7vaVfKDBjKI
GKHfE52uOL0kNZnwMcMWcpPkEC5n2PwqTzkgmQG0Hls3AgrOH8Qf4MFMOeF6L5Xx
IIcHAX2rfXh4hfzeKB+N43ym/wT+3VlDh6uJzqzoOXnddn+v1fUw3yFE7fWj4OjA
GIJHZUMhlDLCGOnDi+zDwIvO6g5Hxhux7Ax+ZjYKLCURhPAJjHSYLNs87zuGJpe5
XlgimimyHIpIMkL0RHf9hHeQuETJ/krlUb1ibA+D1+hfiexhRpHlUHfr7EGwTsk8
a3Ivx1tqS7pwfZuFNxdTI1a48RVOqqWfN95726c/AxFrMFBMSv6KxZCUX+2xMw7M
lA5we9OdZu7Wr1w4YbSuQMP1EBm6vDkNisPKe4yv5lJjpg873FngP5t/nKUkwTEG
WISMxxKI9VOu9XQKCEz3YUT2ficODiDtSbF5jb+umZM2CV0s2+wKcY8PhxL3x9Fu
V18hre+15iR7UM7OPpypW7XVv3Hz+GVkyGDfgWASKHTncq0VArhJLOtTN6M3157H
0r+Mp8U5hkIv2PdD0ojAIt8Ibs4THtlDbmQFAiiomSvRgkfozR/tH24T1sQbpiUv
u1vsCvhx7uSQDqAZ9a1p24dUd2p3mOMKA35IQBuO/ftqOu5x1jDoWypVRU41NYsj
VSwJYt6NOOKaz4mBrR8vaHxBzEwql8AznCfMVkItbgO4FIkNVVarOjfnILW2oSyv
IH/iAb8A1YOtU36WY1SCAxdJGC/zHgSEXt+IiRY9mWth1jOAP2zK5vnFl2/2apIQ
Gi76e838ZhYWXjoAiUYrLyvg6U52yvfS/dG7KB6GE/G04qJn9s7izXEpNd4ZPhjR
2tvDE2ab4aSIECdwyaE3RRbhNTT+OTQB1fDW2WrqoYGJL0rvj8NekURMVwLD3hEX
RY3tBbS1P4l09ZtJqtX3FJx0OqYpnDYd2VxKbTQaScT+Btc3Y5UITy827Tg4bF+u
jE+TbrZBkxiDbFlxeFQ9naTZbJRsczo2oFamKQHZBlh7T7VuNXLW8TUHi5kP07st
E8J5vODPeDMvXZDQJ2DrQ1L14kT4v3PSu26McCTIRqxLuMQFFsDJuRmmulkFCUS9
IDm3FaMzHE0aI0j/3z4TqbiO1P0hSoqe6+ZSfJ8m43uczJHddpfgudcuvuM9Iz1H
NNT6ij+/cidnhlIhvHQC4o198iB5mTXwlGO18m8Sv/Rm0uAiTLmVxU/dkwNG36QY
TjUPaFXFHtAGwA+8T9Zuvbc0dcU6uTLjtF1Yx8DQMaBLfEubkMF5etMUmqQC2GQ+
U/MWpKiUEb+vG3e2/p2sKMju6jIBruAqwp6KmlqECUMJiYnghccSY/dNX20O03Kj
U0qHXPxjOmO4236KjBiJCOiDlI5YSRFE3PDTDJr5rhbrCTzj1iiFf7VAMTkx+yXT
pPrVo6r505MIxug4mZ3ewHj9Ka2VkB+Z8TLeELosK1+rw3rhkS3ZqwWaWTuN9j5F
IcSQokDH5yx41Gw0X695d1gM3pn0Zifp9//mQHPYpR/NccTducbYLIhpYMtFotza
j1HXC/EFxqz2/+C1ceHLWLTQO6hrdzNTaV2HpOdyEC7eWK/+tFkrHSDAF5duCeyD
EqyNk6SDi91aie4WgIFWQ6tkaCWgsKMoRecDdKdPzucIV0hOx6VbU9Mk+D9U5G+E
uMmklKJhfTh2dBFpSPLekwSfJNllGpXgNHj6CgN5GqvUy/a2Iy+lfyydQN1lwyXF
+69Wz65/ar46Gc00Pp1V5gl1993sH1AJ+dftC+NtI4T7EhnMgtN8yyKpDfKPdGmS
YPYQIeQDX1xmtnwIu0tHB8ruJ+r+FfaNNvKflOeqs7wDuYh+u4FtnYkOWllrTNAA
YycnOwUbuj3am4IAbJkYnqGcqBotW+Zh/i24Ob+qBPk4IASH8Ujd5RJJEsghto//
qLLqWcdQaiQUU0zo9zEedGc7mA0KCRkTgquT/IDrTb8cfrmv2YsgGZGqY3zIVKSR
6wi1yxunrMkQp+XgNOrupENwyhbVztms8OgDtYRinsdw1QD3XVvsGp4xgYpmzkXA
RiJZsMjNi3W71ZVChuEflFIpmk8mo86dsj0fGuhSUJShY+oQEPLvWkXHP3Dnj/Ew
XcJLUB8H877C6nKoxuhMtm4yQoO+fIX64kRj2KSrOGi99YwGubNRVuHQkmTHR11B
xmnnP9b75D/Wv4A1H19Ug5ZKt5EtEctmdbnKsesMWHn5ug7BgwPBCCfKObi+AlDT
dYPGT8jU4gbhKO0OywmL46OcvYjlZRMSAivuKTd9PVCLtc05kvXbBSWlqIzqYNW9
yGRGrLdimdFcwD6D3NBAaZos8M9/FoHMe5khDc7Ckf+l0IB0MFElWAuyOZN7ekbP
Y/t+UKsloJNZMRZQ6ybjH09Z5BzfIHZc/88llM09IvsTKu9qinZBkR60RsbNl1xe
2uSHOqUyf/7is2T38aq7E4t0536CR0twd6b1ukuJ/kffbQuqesbQgDAmLOLXLt1x
rhQR6jNuBOCW9FDHE8VO98ECppNWMrBzBENygAW1nAVd/3pETOoARc6TOg+ttFFX
Eu7WuQDyPUiScAN8mmN1QOVgN8i/Fcb6N/gqyRrXo41KNKhcboyqeP54BsTg9hGP
5hCqr9a/7X8WnHVjI+9+Tk+veELlwRvpqOA317tRIvLY1tJZ7lHmbZOdj9K7NELS
XcMQ/nLlLi5pggnK+HkLQdqVIO10ZvhFqK89KalY6OfEbhPMr4atnXJ5AIBJoV4w
scBH4A0+rSNHQSoYwd5QaUqzYk4n24S6KDI288LTipegLGyoudLAbnN2AN7Wzt5z
nkDPAHwNkretSfUFH61Ipy5/soO9lrR40NmaZqLmcxxAveKW1EZGW+pZVNJ4Qr3f
n+gUX+or81DL4d+Zsc7m/xbgIaI438lHZXVRRXnspILWqWTUVmYAgzXVuLvz+QV4
9xgEb1vjMTdnOlmhSTUwGAB/Sb56uwcVoVlgTzIQ/1OGQR0MdJpzneN6ySba6IpL
E1Da777wTI/yjQ3Hpp0OKokYcROwSOZsuf33iCHD8O0Fsd7r87TIMHGMttS1YTr4
99Xqc0O1nKrs0YVvJfJg/Oiu7/1Zp3jTdjvR9TWODo5paPJ1t1pKSjpiQn0YNOP2
LDeZuCDMQS7vUVJPGO14GagHPa0ddKrjxJhtx3nNG5KX9jTF9S56SOxa2iJAinAm
7A7BDnQDq+rowE2pe6kvsruA4ByegOskn9tTHMYkftqiBdR1NgQec/074Xydj8n3
+iMmhCaGI6dVWhh7XG8XNPy0+Yo2ZEvrOUA8vBN/KFw+zxT/6VHfUIuMFeK/OB2v
DM5IJMvNa7PVgJsnbEHhN/nvubTocohInnkJXNctNCGn02yCcSiC3eJpQ9CHIXRK
HrWusHp3lJJLqit1QgtmBbnty7yphZVM3x+KiEgYzRu9SY+1Vd4K//EAgDcdVeVV
JXPG9OH6m7OreED34dPouCilnjhGRaTtjgwy2766iUSlRvbNUx+Gfx5dW0HFC0fX
tkAcJFLGcHWcMkIvmQJ9aou5G2XuyuOIwwvg1R8Y+pKmz6mLApw7Sj/yzUVg8VJI
/nybp68SuKPfThc1dxZZWcfAaD/TDJDjk6yHRDGkxt3/2oJNnf1pedOboLjjAiJX
wZ9FAkL141SqyHbPUikVanraTdM6eIvu+nnrg2MdnQIpKPUSoBzX/3dq6Orog8mP
2vriZ3lwzNeFm9NKE/LALVa2Dny2oup4D7Q4CrTHVE9ex+m8Aygg0slcuv045ZbE
HjUvNMlPnYKx7mSc3bv/1z7m+GITZcUMhAREOSpDbmWn7Ee2Ap1wF1+JuauJ0f8O
IoUlbsICw5j/dSraTSwCeUverT/PeoH69pPl+pPV+mYa0EoSQv691NhthtkoU7q7
h4AySDZkfcR3uEtdZ4IxXXXlYgvquNn3XwAdch2qVfhFY1OtlH3ojQBeAAqGLHnR
Dlo1nWBvyuVYOyij1bULZfucRuM7t25DKPSpDQe9OZj1q/b/AmeofiOlGX5WNTPT
GpuTKf3tz5l5mKwMyf4XSyEnw5W3rQwRPyOK18L5CpdiNB4F44WtHR5N7nIsJMNb
mqFCuJGimk6UMIExf8vHKayFjl1Su9cntKH+0Va0bZMbIEWXlVCcU7CYxEITRF18
sEOfYJYOIzq6Pq69jDU5V4ntY7SM9nB9FgC4TXHPuqSZKTNQacqVoG2B+ZVNcEhA
tGYFqZZjZMxOEFBk7IFfKWTc5VzzeuJWIsH5+I/5yXAGAC6+HkVXa8QokXdDCpcN
4qoJI92xUQa8RKhEByo45eaGVyr2PUPV6Jd4M74r29FOlfoJuNiZ2gOhY0KWXyR/
euztOS6IwboXfG0hfE3yuSotk4uyJcMVq1xhH9sU0won7JOwEtEpbHeBAcFmdfMA
kJlSTjwXhHTKoQcEBdp1zZXWejTkZcRNyrZFg4uX3bxr58lURbbPalD2WCb/DgoO
EHXCF7m0e46h71TTLxNgDhmu36XpNkqAsgBicf2fIU4P2w6J7+BuRQvDMSek/IQO
O4PwYU3fF88UTNvNq32PpwAFFDLniSHAgfO+9a7ODk5Sv1dMc9DkyPBCxkJjXwzs
6MqrXRho6ii0A1c/EOxfsln8rrsCD5KqskRkvGPM5DId2piWjuIUzXFljVGufeNV
8sLsriohHvBQQgALP7cuX9U7HaoDIrVGJn4dBeL0xy+LwzLFHW+YlaZfkVSFI2A/
QJ8+zp+XoJcDlvoyJtbUPF4N/lANMg5DVt2A0eruCOgdGolgMzVwkVGqDZwlkORw
1zDONJXB0Wx3ciAfvpEW2OGfAXRS7BpJL8sHpAOFIDKzubCyZkYly1YBGR7ydKLI
0gYSi8qDSIo/qSaT4o1adGtr87DsEiDPAj3XxdkT5LmPQ2xakyvN+qHM2vF7qdKG
1i6FijJ/cm+yxx+v3eijXBj8Iy1Qo0HvZtLuAl48Ad0TVNmu6epCrhTz5zhN4P8c
kVsL66DkU/gdAS4fMFiQ77wWwkJHoc8SeT21GNv4eoSvRMa2UzWT/NZJQIZN2fD+
csmwch62d7R5ARWxr7L0xBR5RtWqRukkIXr3TH2b1xQ+8DSKH4ZPxNSRMYcn76q1
URA78DjAz+n0eUOA8YFmA3WBl+EkVJtnRT9M8kYooOKdqZF6Ln88RpqLcXeR5LfA
EfZQKMYMtgpr07bLknnf8BNHgWM0zKUsYXrI8P4TSYafJrKge77HIokd2XMOq7qe
VT8WeDlKxxTOdrpnCojDAXH3xm5DB2MWo8VkxnOwvIj1hDuACQezhfeeWTdnqHWN
STQOUa0oSCl/5Jt+bW8b/iD0OVvgl80WZpAQ1u9vYtSiWQjub00MlC2A05/1zI2q
gEun53gNWD7TpCBy1ZZWbnef/AC4r/j3lkpiGrYU3tVvz36bVhZLUnwufI8lJ/bQ
px1m3o9+fJnHpKl93DntrpEkU7EkVhB/FwlZAGZMI+MAfFxid3g7tq8GNRLizn/n
YtZ9VZYeTaPhme9OU/53Ee+tDLtVpXm2taDJXB5lVjAYomQYhm/nYCgrtILJ3A/x
ZOXv+rfXmX8aT/DIer+yOysazLxRvESRXxN5zalgQd6+7e8HprGl319pLJKEk0EU
aeTlR2WLznMh/shQBAV1P1Z9t51fBj6D2ffV14C7RGp+4XF9+thpdNEotNzFMYDO
fqG4+JW5ZdH486BjcfZqrGi9bKg61AoklFl8mfbXm+yESQGCPi5ZwVYZ7Wjjg8vi
5e23tZns709MQqGG9WSUpku6aAtdjGKR8JJ4kvxCw4TAR2Uw8kH2K6MbmnMvJCv2
4Q+8ti+fN2B+FaCDoqd0a6B3Gw31oQVZZxHPkwjVLL1/dO79Y4GLexQsIC4dJ8SN
oHLPkkvswjOZJ2Q7LIRh4tkcpIFtS5CpUTizMeuUt9LuvS24BQbKGcUGC0eKk4E7
mFEjSG4Th9SE4Zqb4Fvwdyecawn9S/fHIZ/Ttn5Ck9uGMaMnIMW71e20t1T+Af1L
y7vXcvDIL4FBN6PRUny41e3gX70Q8mZ2U9qGTSEavrCsrJCv1E+K2rgZBNyGZbRS
RqDwWfHoplKR7BuR5bH6ZPaSXCKI1Pz9t3B029DPmF8Kk25r8K5TKOjPrIctQWxE
kll6VMurqhbDAXSCaaMeqyHj706RvtEY1/9zJvhqTN3jJ0/N0aAkEDOTO77LeyUn
pew0j9xRmXcAcRTyoYt7PvacNkWq5ddiJuTcUgJhxE6g2UD0pl3E9qhz7hbbpLdy
3IypRMi6HE5O8/FV+7KvZg3TFQYut/ga1lsQ39+HVxi3Xuzxu1Ezoc8tlDQ8H5Ph
53iuK2HLi4eDE7hcCCttBwyRICfMHlQvCCfJKrHoTg72pvOHb8t81B25tY9Hg9XY
VLYJQS+Ebs5HNb3gTE7uv1EnJ9+IID2eXnFXncBsFnsw9ZJ6q3+fPPqZ75MvWmnT
hH9Yi78GjF2Zk/7ilCb83BH4LmCrzdJDPpEzLPBnpnitBnFfYkK5BMEyGsabzxeG
5JESy37tzcePlBT6RB6vMxYe57sRzu5wJlfHsh75RdcrnFHXimfe7HWSkegnueCL
awYVptop+vl/ZjG0GbbcZpBKD5sgbjtotNlZvfk5lUTyJWMdCTklhh52E6bkWafD
NeMiib770t6Carf9Xwo07zpGb6KprW+zJqNyyDlszEh/ddwEeTnU7La+cGd06HEj
xcXLmZ4TyfdU0WtaQwn4QSxfedJvm4qyVc2UFysfy/dwT7D7GQtHl+CyWt/oVNHD
2mWwX14dYbBIa6lbCZ8+RFDPQU4Xmws0AD6vWLQamPKntoa/Z5feT8fy3oefmohK
Hx86vHC87ux1HnGMSnc+UrIYNg9N2EcNa+DnljlfWEy1Vxnfxq3yOEwJi/ORFO0b
j6+DXTsUULYeNVuIgDlf9Z8UH9KNVPvxSmUpJ5V7W1FaO/+p3vdO9HbtqKhB7g56
uj3McBUze1buxx2iBVh19QmmxOivjT95+LL+2sAUKYROkuklQKSg7GHU25RYZz7R
XJIyBPPIyKc/v2xxuEU7JSF+m0Yq6/bJO+ola9f/jq/OdQXCS4e+qORvqGcaocms
hKhS6sXtMcOX3LFXQph9bkPnc3PnfMNFh6n14b4ygqkaIHM/P9dITs3IYq7LBVTC
Jmefc/d/oy5qvJDCvrsQLePYx/RkYqOdbiXAbRplBVkhH2NKRQ21L0QRkvekNvnY
YbxzlctMQYZWZ1lDW3yTilYrUbER59A7oxmPaKc49oo/RrueYIe7AFNtswUGZVAV
JAVfZ81vIczMFTCgwlaIKg==
`protect end_protected