`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
AOm0ifrO2lG9CKGJhmiQI+aYY0VdYSC7Sj27hwFtHg+JH46LJLfxCynUoOrIqOg1
opUkweCcfNk5KReFTZ2epVUaQXdL8g/1tGwoXOj8tux1egduTrkRmRs1RsLmvAaj
EaCMwjS5aiLv/XnLpJqqoUHwR2GZF5eXTwiizgjy0SKuryMyW5xeQjHkaI2Z/8X2
d483NqcUrL1NyAm8AEdc5JJr4rLfjFyMpgUgzoB6oGRgMmnBKal1Q7xcCo7fjFEl
JaB1DNH9EwYGP63VFD2EP/Sd7/ONTE6eHnsxN5BkzCLkpRv07PMp4UaIf2j+TC84
PhXte/g0yspiNbA0rZwbWHveOTitKdh//x7XoL7hQXll/gHLd6iBMb63mP4/MYaB
qWRShmp2NMtUd/dkUHqzmSgY13lvPp5fNlrOWshOO4ipTarWT1sb2O2T5Z+gesyt
fZwPFDSd9zk3bGjqd0/o+IZ7rc4sX/g0+xKi+Q98eytPetwRlJaYZ3yMEnOooSmT
pmkb7ja7BM5JbCrqA1/2ZHSDlqtQ6AnCP+nXDlfDFsGLw6zMtOE3zB+JN7YCWZyZ
7Qh/VLzZ+8TF43mZyIFB8/A7vIxvFbkmIOI5keI5fic+m++xPtFJYWVpj19g+n93
HLuaG8Ow7G4dhVbkijQ06CRiRrTR6fzHo9YTpCEeonOTT2Ln1GMTllTIi0J1Pow2
gVSEoSbeT8BKFdYf0gCcsQZSTZYhdbnSH+k/kwjhXw+UjK8mbKYYWiD8C24uLZ0b
9aqH2liCheaRslvQcgXHkKCNb49ckrKCNaXiyNxMx9YyeeHlDMPA7bPslXLinDm2
KjjoRCbjxmTYxhCdZ22gNSMcSFgMLIZdmBiyyMpHEOHQ4wvwWu4nifunCoLwbovs
zHaZ09WOb2texUis18Lk21aJIwksp3gySWFzh4Z/eAj9OZKGHlQ7AEc8vO6pBOKk
ad782udITvKUfz+b4eWbvdtQ8xJ3w7FRLsKNOu6R9QgvvQ8/JhGKLBdQCceG1q+H
NNJ12mauzwSfb/89NxCQoUnVB6TSreLWyJttpTPkNQBNAP7zsDkG3rLW5IA05cIC
sgEsOcCYR0CTjtTW26b2w3Kvlu9i4Q0E+3+LognSQkAMFOglmo+c1kDcvlQthUNz
C09jAF8suTYx2lX13lBNtTsPiHAG6fIxyd8rVOO1zQn2zAWXzhTedF2eRTNbhqqq
h9nBkXi+qvnzn9lGGhGShS1/sv4k0q6KCzmRpUm8Ww2FmbsmdW6eVD2j1B6DP6Nh
QkxH7t0ybhrRvxwcP94SrPwuPiux7MBaUVPuJYGVNO3ob+mKGAflUhaJaSgbq+sL
Bj6g7BA3QD0xC4vBHuOWwzHcF8SEpQXoYeMFfx+glmFbHRGwgyTGT39EMRmUkB6X
DB2GLZ+iswmgdSuw1c4j9JMOBBzMSvMSfHY8ktfGpbWsJrlOPU+R32n0JROwDvwe
dExI26594hFpkBdeVtbwuF6dBG56hahmPlJCNFWAWlYtcAbEPM7/yQHiggKbdgYA
0s3SYE4TSXDHNuTk7VNUzxKVFf1E7aoImKTVtv/BbifNEHczaZL3GVGbFXxzkUdm
MScY5j00dVoS1WU69oT1RSADlHoFJ+J0AQ8Vd8VYoXKPYej3uszF1tEH73M0Yi/p
FQNbGgx2SSv2H4JxD44mDlQ6NHGRTTQK/D6DBk6T1nmwqrYh1p9BwzXRDrCWTzTT
Mr6qmaATijT6grfpUYDpZRr8/5+pv75HlXZ1n1jCa2VIrAbBlaQNOELG9gddJLTl
aGiQF6MzdgIQfD2qo9ysXcG99SHbJ7U3aKF90aXQm2S1wrcu/caVmUfFLk9/1aB5
cXHKOgAMHBJC2f21Nt0zRBIKsiW4y1mOTI3T+lUCAInQTTbbGqmRhyWoTS2jR9gb
X1xjWz8niHSFhGUDM5DbBLU51CUpX/hlDAMSKwGZlXHVMAKeCLd2wfGbwflXuKBI
0S3wLnQm0Q4MYitHNyklWa9h9Bvfuidmbx4ECRhyaAwlLkWGnk+rFKFSRq3cXF56
QF6CfEIXYbQYj7nkEKBwVedFMkL9JCSlvIyP/rtxBgX2Fc0zwrQVwcOh4Pys1xV2
Hg+StfWl7XHAWScb0M4ykltfmjim7yd8Beh9mXVxkW8=
`protect end_protected