`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 43504 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
VdW9QyppGxpRdqqH8iSOFs+qluu2m7KWj0P4ef+MruKlk1KqojOxULo2GPba6Ipr
zmZvjO/OWd0HecPA+0YPAb/JEp3gaDVWioVFZ5VwnyyVBZUi52ZQwNB95EKzlm6V
Hz/oI1unh1vJs7dpDK1YBl2AYL4j3aah7qUIOaajcT7hgBdBKq8OfdSZKINdM+g5
cyIBwlpb0CT+tFyhjMF87w/63ssjWVHpvvD5LwaPMieC9A2lPhHAiSR9SFDc5tL2
5burnhZWfnHRO/wFTXdcXWUXQo6qhJJ2q/oLsmSPaydNsCDEnAWtTnk6ygmq1TYB
0VLrvtAAUAe/egWpwlLy/EJpra5yBIvAlYfwOp+6Ik1JGeL5qDN7/mzPTH/k7XUZ
1F6lK6F/lxa43PiFj5WPMgg5nYf+3eW17X2xhD/SqwN4Y1P1jGuK8syru3KtgQAB
aDvEaR90W1gJSBMBnEkSz6MmANZilnHOrqtIWv9H8dU49QBfl8vCJCaaHwW7PvmY
vEAwcaadz3Xbip/gnfoIGjI1524eSLpWbH0J43Y0E7GiAnmeO6hV4St4kU5REt5F
Z+X/25Jbo4YpASc8hgRdBaM+C34TT0eVUhGG7rCDWZQhB9niiRqtt+Jxbwc6I94x
O2Ph+fuSkpEvLrvQqwh8PBsKIAcZoPBuGn5EMO1rY5jl0jxS77g/fbMf/iTPJbAB
HbrxW+BX7y7Q2lHeLRVpo+xoBXkvCWFow0x//l9QNnYJH1IF8MtnQDAuxU+Hdn9L
1RPvaPVYodvwUiWGHH87TVl7CL9uhLnUmMkavl9tzizC9ffJVsQ2LbjjXVIBmu/m
TFM+iH57jDy8u5Ux9EVr9Vh1neC0XGwirAeTrO+ziNrpknC++bnddPOWn9quDXhk
8/eKFkgrykmmxYNs1/IfHjBLBOC/pQ8xCkqrsFo6/E6qMO/hC9GdkQOP4dYPmnaj
2VndZMDOk3rMyKgrqqr5JKistezSzxC5OCJWzpoznHvO13pa54urDgGTTXqhnKIK
V0Fk5qlqyrukbaIFzG7Rneq4OKJH96bJ43srWODjgERq3j4QG2m/DoNlIqIkm8A/
QqZcEdVX8TWc/BJWHCklEeMnt6/j1euHZ0Rp2mv3uT9cXFA1bfUKnhb+Qixd5D4D
uKoelKe2cb4L3fz1s8f/sU0H/Y6Q72JKXECp2P98dywnupTVztMYN9/uHAz+vErU
5pc19Fni3H+5v45FrjyRewI2T/26HCn1FsEU14gLMo6Mey5qsi58HOs4fzRxk2kP
7tus6nKbKybHtHk/pukESeIFYcQ1aL5FWyPc+OLlsERIU05NaQ1rGsDzw2rHfZdG
uzGnUn/gUoUcpPb7brd0dDMGdS0Dfm7Ro52KWhejuPIOxprsP6SdEz4OmwrvM2A9
bQvXgAfhiHSRNpD6qlP3CeWptaHrLojYtMYfiWK9E6PqC2Q1pjQ3GtPGDZMlp/4H
AgtJfkfHgierZqFVNy7sA/9A0l2xeMAdFwzw22bPyJnAf3WhA3mIBNe7BOL4EJxe
m9oI9k4yck+rIbrZnqRjeF0GV4mWM8ZkD+QUAIfSsMCpQZ9rWy2yR4/Gzmmo70+Y
5D6E/L36hv7iWnBnOI1FTiiAzMDrh2wSDXt8kXptpjKiL1yIH4tcPlvUmq2/CpnX
BpxaF6gfyyDfeHGLqjPqyuBJNDjGyphyeBLzEBCzVBehm5SLmPsDRmvSi1K5Unpo
+lb2WSaitmOO4oRrnH5vSpv4ljWvnEcX7fzRdwD4+P1yKqB5U8K7P7VxIDSS5ivM
WC0sHs2gxtE3QuiI1vVkFAh9yLa1/98IhESMCFhLaRay13NH4QkdDh3snl1eCr76
+sWO8jnJrwRKuPi3YDhnPUBSwVV9arU6rQtxAiFJchHNByw1D6/jEbkVlw2jQ7A7
KKIu3TNsGXOGiACIIhBzAOA4tWm4Vi9NTQJIonziAQrxcvFqzXGdKPSJP05XLaBB
8NAFSdBqX8eyfFeuDYIFPJwc9EPe9rKNZ3etioggJlGK4YzDEwi670krQRiwltY1
OR3DdPaymVwzW39Za4r+sizEd5TTsiHX43Pr9OdDOKii38UOWy+TAZCCKrFcpGxa
mahJgtSnB1qQQWquYUt10P/g0JzavnqTKskHGD/7iIR0YgbbYI1mnK/2BVdCtb47
2X/5GXtjn+r7FUW9/HGZzJzsOSWKbYKppOlcQcc2R90YvdgbTtDZYmahXity2NG3
TNKefENQQ6Ek52/T7ACvQ4b+SXh1AlZtD+zGfItSLQlnwKGlSQwWO0dsWdwMfEth
fKh2loTykBgebzYWGF6XccG/WiLrNpT49/pnc+nAGew+oWs5hrleT7HWzSKQO/uU
KFCidVkZwmAGH86RGkDf2/GqWodXuwn+AaH6KBGHVc8v4OVAGCw7YSalqMb076kM
mdIGrdlkFnujcMQK/MLkcNv2vQfVu2EfYPuy6Ud4FTI7j4IrXfwz/3vw4MeduEpC
B36xZvLJCA/3mUMPW2YkcDLenwWW7j1Mg0JtKHAuKMXV0lIlLqcM0mGqJClOBMj0
cYqIAmLncS6B7nv/e721yS7dNI6Wg1gTj2SKjVVfQlvLYUUoqN46J7jBd67LaQaz
/5pi56+Z24Xo2d3J3IjOuS5EqgITQWaP8tUxi/gx6mfLg8kNt5NHnoNC5cCQg7eW
KHU4oWvdvEo6OSfMnS0tnlPR9Edo25G5xFIf6h/10JCa/i/wLpZyQ501vew/Jr2h
3TyY+HyF4EpAoL2HT6Hc1+bmFgbuxeNWbDOkWBNgnoi2SgzSBjYckBGTHRETuq3n
JBY13LybFG3DMpqZRkvmfYK68b4EEx45WVIgbjzIIOsOWagKcigaL5rWzXFxgiIi
ZkPbE65Vew6Hcw4mBLwj0ibKMH3A7ddUSyBIEkAkoVDyhEDQ+8OGBqcIhgHKwqrn
J/t6STDyYesmQV1sVr6S3cIb4yXU2hnZTLvYXyV/dwdVkp9V3/NrDmEU93T+Eg0m
+71hLlgI0rOpSRx08VM4qgGNt2UERg+GeVttRka5H7EZEqKymzJ9E8vJvU0/RfX7
4tlfdQG+1aJqrfz78JEhdCi3Hh17oFIBXzwOKiun2GxexnhBviTFJ4W8vlS9E31l
mSTFns3LMPHxqLVM3RMMfO97nEtWy67BwiF7QbbKCiCZoj2+2jsn41s521raBl93
LPesSdRxdQ75hzW561KilPaRAHr0Y2QDR+RsJBmBOfnW/9WPyRIfatFm65sA76y4
efBMxj4p5mCXohGaeGESqW38G12vDNqQ5GgRuAa2tDV2Ww1QmdfyqhYgHqpxk3fb
g98kW0/VwsvkrE4R7wdl7Z4xzJb3qloX4Cj55D02CqLC0B3Ocf+BiUNMZD3u2R67
uqpUzD/fqc8rKmAL/ttSXzMjxS/1H18EK1LfggoqoIsvqjKSWYsZGPOeHl5M1ZE9
jPmKowIpRmrbqyxLRsq7TeuWBe6CnPcKy8/UzdAgK4qCAPpUKNtutCsxWFS2tH0+
4EmUgCCF5rUugLiyKDUJP4ePpcaHRj/8yWChsKUkclm3mtoSGaZJQtNbBIIRek/t
OgkPHjKbKHrtQvLh5YqN2ecmlzy5yogIMn9R0q40qhc76fSE2iJT2c8bXWaCrseX
KCnOAOXe4uTAHfCSXQcr3sxy9qR+4onoL0zFd+NwLjpQeKbDbWcLrMP6S6iztEWP
cuaf2QL0JaYJ4mhMpF/R5cS2gWfVcnT3lC09bDJ2EaLOooJZMFRITBRUDt+SRvxQ
iOOHuFX4UPT/GU7lliCgXZuFNwauP25+F/THvxGH0V8NxC+q7gS4uljke+0m3rIa
svtbFqstq/3seFaj0TOIb3hkHJIEJNMGEEz8Y+lgDYTIHCShVIocv9s1w+1dTPxj
1snmTHM5H14s0swqBGp9CfVAuwuLRs1trwdLwii08bA5tAnuxnqRZpt2Vr0i6fRc
C6TvQASkvMgiiobtdcRtqF6KpJfMk7d48C6dif5ApMAwNEfF3A6dJ7k1JvPTi4ZT
ZyarpX8LX//mWXcm0Dou04V8Ec1DrsgYBWzxSWEf5XclktbBcxtQ0pfK82kbgyl4
fPwU/7oKu2R+ul7Xx9gC3O0SOAK8tr4WUMKkXgQXvGxuBJO88KDfGwtxNEcdvYjF
1faBq5zhXHScwQWE35CweIcx8+hcpp1wptusQpirkXxASyMSEq8axrBZxnN9GsrX
zTETk0Bg39Wiq5UxFXvWKIJNDXJEwUcZAJ7K0ZkkurR8oDsoxcaleU0t2p5Npusp
1pqpiIisqtlhEzs1UoNMKjWCThku3X/W0ndB9arxtRE431HoSJMt8v4vXUxnmTaO
JOab1TjMZ4HQkMoyhihbubObkV9fXXXFJ942XzfdFXB3Ep8CVUVKhOrzK/hrx+6D
+DQ2rdGgT5hWtdd8Q/OiQskge7upFimX996du9l8wop3wsFLrCNAAUnrAWW30cUc
JuVQU4i4iMTwMXcj+IN9DG4AyCwkalxv8kBXH6ELqLD4pGR7X2/rsRmTzB2BQDcv
q9eZjxRG8Vox15Yf2JcM8L5An+sEuivGbAhAqll11ezRjv4+BbbgQvNxOcFueYr3
hO2UuA2yX/HDeDZBEQAjuIZh0YGh3m2KksG+SgvtCgLlRUeIcJXxEIJqdZI5gbdf
RQ/ci5CI4Hig790lStRacdjMHKLU6R7wfZMhNpyMHpdp3bMIp2XDZgZIvE0JhhOO
+cGDbaPZYlgckl3V/UvJgNPfVeqOnIGsJsGKlBPHtOu3wS3V3mxsB2E1uAKgIPR+
oRV0uCDJ2SDqK2kbbaPlQ8car1kxa+kVhzyjB9LLDuWFjAXHqfUNLLZ51P4Z89UT
jzqOmjDhQXJuGchaRlhA3CDYQhLiC9/42RkGutluLy09AjqD0ZRYgx9HMiF02Im0
J6cuwj1Z3ztmsBcG7Vqo7RnoVPXd5txDey1XGxsIdwKPBuALX41yVPtPF1PnIiBE
NKkwcVVUHonXlfmhbWzpZNd2SyzEcAh7KXAvLdUkTcLtEQrJyqvSNvwDVEYjFrre
2sGaZ46jpLkwDfHLni+vXadBsX4HSaWFh+yfU1LPHqlgD843Ycu72CVCFTCQKNiL
Xy+YHMnGNNGqxZ1zMXd1Zg6Nvg9HvDM8MbpYqPLl+q7aW9VegoC9asupTJ8b/dnP
LTv+B8yVe5HsAdp3ECHam5SkUNqSAyuPWLbLjr0aIEbt+mgJdOfY1r7cvUhGdcac
UdOtlQtEF3qRx4uC6l1UXihQHkXJpEz+qArtRxWy+UZKzIlzBQEkSL9gTZ25ejKj
ICVK9TInc+pGJ6NRthJp7jJ3sJqYtu0l+TYyO8Kxi52kdeslzQRco0JQ+dEpKD/f
8eouolq52rAzjnzINnECNI7Pd0YbBUslh6Ox+nCvcko+VG/3v1VicMd+5ofNguzo
nrvxH5pZfEZAsSozgg1apIYtr/8ZCPJT+XDzsVkCwLm9jYAyIymWIogGQqeS63b+
INZJnMiQ1mIudYCqRz9wAmHp41NeLXfT1nLLd8AiGFRmnPc+kwyfIhcRYIvmzfSc
iyDYTme56nEhnipjXTs8ACE7HofX/aXri0CS2JPb3YNSEUfUnvYsKI5UCh1A1J+n
JtnD13ho0z/vwDhDCk5enDqeYVZQAcRkW2P62+fUAPglm7qHh+NoA7cxsOnBk47K
F/2ghSGy6k1wJBoi7cTX81mFbm/AVb2YlZahnWD79KYYoq/q0i9gkny/8gY+UKlk
eUnyByaASsixWqYNP8QuAiB5ZR4jkliNvx60qRDgSZrEDiGGJI+9+rQFUaC+dYmj
59JaEafyeLGmaOaeqgGsH/l13dPZQfBFy0EYwyg6R4G9neDqXMEOGI4Q5FJaB64s
kVFlLepTIqAxlYg8pKRKVSml2GAnYgWZ35JUZusH5gL9Fge83LtMOTKUEU6qOCfQ
heRu/1UBonukGqe/l1YqCzFZU79pMpBZl6WQMaqpwPCm18gpggF/i0k3kIJMc1cG
N8vU08HxD1dvpqtBjdi/i1WZcj58Zh/5Lp1zKHHQ5Thth1q8FklQchHGRxW+v5cp
Ro8jaFkXJNlRIXgD357VavyVX79GqMSmuHzltuhy9ORbBLyiEunHGYi7wL6Qb8cW
sNVdQJoB66jHwZ9DnlPk+H0c3NcLdB1uJY5dOqsyJjMgHckUwBwE/SuK8TtafvXK
8Y9lNG/j735zs4KskXNFcf+wwBZEQgrWJyGxcuG5hswNDAtghfAlKS6lptNuNoc6
illHIBZx5cUDz/gQOxIb4mMLHBHyOiOfGWD/KqCTV8AaeAiG0xEGVxU58NVTcJ8X
YXS9NJ4kriZJjkEK0X3a4OaazsuLirGJPMxm0IXI8jDe1oP2yMMDpwEezqIyhMWF
ovok+K9yqJwE8xENcWVGDni1sbMXztf6dmDKaaHYhk+pna9ILS8HD0gKvMeQggxm
+CRYfIFYFar+fu0S+GYBqpri2UqB+C3v4BmBhJ8ekLrBsJcjCepWmtDW9Wjv2mb6
IjVqqB2qczLaIgD+efkAxovqNK8qaImzttjj0DZlYe+I0o0H9EX3D8GiMPl2m2rk
6m4/TV2estyf9oT9q3uihw1DK99XOIeR0mjU0bfWDwJ3DyMdW87G7/3yAkIUMBRX
AYcUnsKy62xv5eUNDu0ldUwVLtw5wOW3BK9213OwXUSo2iWrRuhFqE/giLXr4faz
0C+vy+zvyMqjiizVRPh6aYexBIZsR/OI68I/xQQzEcfku8CkHLuzydojUw96wuP1
deQzFVcBnjf4rVSciiOGVeaFFZTrkko+kXl1cAjoKqgjXwjGsY7yHxHoD1EyILVm
HOPwR1PQ4HGeEVAnvHtQeAFORWsWJABqBCno5tbmUlPB336eJ8iV143HAZlgcqeE
wGRyUwtUgSKKbLQi4WCw3OcQcWcoithxvW3O4CxgsgwCfPvLkegcyn4ciYazKU6x
k/U5M427inUReKbSR5R8bpy3pnoW27Ocy9dAZc7K4BOLV9WFa8tZv5lvCBO6eL63
teMFFSvnWfPc/ENhrCHxM7fDd03Qf8N07V9UXcZiQZRpWxFpw7tp28hea8Nv9t92
ppKhnFUIj+EHo0++SNJL2L43xJWArZxALpyiqvHthTFqgPcQlTHU5qxwBZ9niie8
OLmiwEVJGy1OQo/7NM03WDcGlKAU2k9d4ggq+cjIX6vcVsyzge7ZMaaimMCG//+N
8V1dU/B3CJ1Wl6PoT7cwlHdFyrLbqt8ZprVOVQAx0r2ZV4p51MX+jF0/glYJo+KI
YJ5ErChtPr9fEvTjZlDhkvjZinqyxppgQpBTWFo6LmV+MOfVahkayS0ULOfeYVFP
Cv5M7oUaqmi3+2kvEkDVagadVbc4tRNdjG9W50EDHz3UmVW6z0A7K9zVaLsEKFFT
/7DRpOmVjG97lzR+EpKjcTGn4MUFtMdu+GeWOdg1PoL8olA1l0ioT1ednCiQUe6s
dUmGSK4JGuLIRC4nmUbXDBKPk+ioWZaotDbPWgp4eZqOls7327AZk0RAki7RNpEv
tJapioSz3t5ue4OsHYFwH14EhChEt7pls2dqyIEfYwMPLNQTSh6/8SCn7YGlInof
i6qa9rVxhvO8X69YyOrfTrwP9iUM4xPDxkHqxagtT+cfed5nZRP0Hg6PmOXZFE55
nwYKjOLzoYfLMpo2ufIVXE+Ur5/Huziikluy4CFloba1JPf5aRBHWigt6tDtSlro
KxgpFN0tQs/IYG8U4HQkw/uERCV0M0SslV0QhmnR1KP+jreF/Q7HwOKcluXUuPrJ
3KYyyXm0Wy+c0WlF3zJNjSpojqG32oRMGC6KqnBiw1wix89CdhaM3f0pot0iTnoW
Zq+HcuFrKTKAK/AFHQJQ+jKlaJ4x5Dpr1Gd0SGBso1+MZJ2/iRXQI+70m/nhCq3I
itx0iJYeDlH4Eh3prCYmuP+Y1GEu9NTIr1M5Myq4+QnOAmexojo4+DodvohHzT2Y
oPnOg4le7Z06qBy1oQ/4V4wzLcfwSqK77UmbQaMQZrYITgDwaMIP1QKG+WBfJoac
GFloMWZMGEZzUvdkgawLypnd3MUIF9KieNF9KUxzN0up7SiMezjb1UyVA22RQ+T3
ocDTmUIS0wGVaHX1twtSIIFBwNaG436XKRvkz1oBFQhFnNE7XYumMcW3jfT5hbqR
SzQEgLfkMxTXVvTwA7BoF5s/OF2gEIdpEcO9p5d3zKbW92ZAmmDRX2Pm/SSmQv8c
PN7dVk0d8Pl01HOJqDRESakjyc+pnKmuzQ+9emnc+FnscjDOAZZ1Cx0aehqxlbMc
4heYB++uER0X7XQwXIJcTTfenDM90aJTULy3Mi3tot3CElhAOvwDqAuIWa0deNRi
eoWCRKq+9CeCJncHoo5G8kW7e0Z38VUQy4tpFzULiSKS83sit0Cce8ER5mk7IxNM
adi2sd198Nwm5vSKrWJeN8GZIdi2OijinR94WAygSG9Mrw2tSdAoltuOAs9GfCg7
+i4qbXDFPuU2NpvajTTcKdE7+Wd5xfHyATN0x2S1wfOvyQspSovOPZvAE1TAOV+Z
bwyja2hUXDXnswq/03vz6/e/fRAmm8ReJzn4CxM6swkwUCDNoa0HvN4MFxGzrUs0
qlyEPTcIjPjDgZeEh8YGkHozOHUU7vpxByBpnmFZYPlPH5Q+zQaLJ5ez0OdyboJm
XSWcJOJDceAT1GHoh2VA1ekmm/xweNf5xVKG/4IwYcpbGPeTc4RP56NeS83I4HXl
TpBM+oIWwRP7z7Bjg7fd1PWKmxkv8yQa4w9f+V9e2gAfTo74RK9np/E+3Un3C6f2
eSmvoKnpSyc6kpDSq3PEOollZ7fM3ICH2JTt4ihsVJOIPk+B/O8tYcevZU1yxy+y
YxfBTapf/FM0HPuJgD1G6Nry3yA5EIDcb0aI3bm/mODXLAs+Tckv9Yt4uRpxSpiZ
EIRjkasme0VmRnKYL2fQqJF490F2SpCWsRJLaEObI5d+QTc43AeVgIlBrXaffuZP
Iqyt5TZ2dHAY6CMYUwbu5qrWn5jQk0kGqA4XyOKVSe2Hply/JyiQ2m5dwBUqvYrE
+77WhLDdg6VBwfqgjhvPvem8p5ivni41CIQZ3gvyja5A1sHBX/qnjbcEj2roJZcf
JFuhlc9e2boN8CnT9OBE39LMe7ne5H4YrwPQXFOipNC+awQ94X26oaeLh2JnzFNN
PozJA5eJ6PmdODcqVyyGsME4QybM/6rNge/vVZRsvnpdtn/ABLN9pntA/f/93ulh
Vn/XoKKgNQArvKlPDDAJ46dfmy22uQzqp+5jh7vWnyl2uuE+qohHsjZS4ym1yAjQ
YP6wCc64Wda6Kt2yHAMq6m5Ckx6obW73IEDB6HmMOxy/iOT0vbQ6fHnoaXsFd3XH
rLwwqLg9sgcSydmb3A1mJeSinkOlkh9ldBHGUcYUwSTCwRYMNoc3HlcUj0cnoQai
m4a2CMy3Dyqzf00eKVtCzQmsn4v0zVn9cxhYtCwn2pgl0qCiS8ObWHBgGxC26fkI
fRdwjR1w4d8pLHB1PzREiTWakKmTLZ61Pn+DrdaPVrCtZiXdjkqjdSiUpjuDLIPE
EptC03OnVdDZA6rtrz5D7fyLqJinEehCo1wTngkfVBefQonvvhXFtV1ZHFYaM7GC
jaUoWvXr14kwmm5O3dBZIMGnWKgPq2zUhCJNbC5/I6neXMvpa/ZmjNsuyU219m8j
qy7gK0x2Ug+DSj1Dgz1qAb3fRkTtAXBaLiP3wske+dkVvIpOSerUrmRj67XbM3Sa
+3yyznE4TuFaI5ZlI6Y+XCikqV9q3tT2Xp9MZGTGbwRW5CKM8FfAu2naxVIgZz1b
fHXqCU5cHTZj4WOyuT1LoClD6b8M5rLE098lo8k6eyXnRRKTwWhJ8E7I5bvrnS5t
qs8mfgUSUrmOz0lq3EIWH54VD2VW3+aooSyUK5JaTCNYaCe8KCDk/bEPNIra9qrc
ACQqbLSpwFK67/mSZm6oFGLF0dj4h0viTmuoz4vZwMVMn1GIzNhtYf3W/QEfIT2N
HgHFw/LTqeXUqFE1LGRV+1AilGU2B21Z32TcKXxBQmXN65MmIA+WfsCQxSJCzJ9r
tk3LKsSPyxGXG3Jdzasgu88pOfmUtwloLoDhptlOKw9QSsRsyb0SdJ3MOblSqUyI
c3qKX0PSLBCaVnZ0DCmUmB8PY6weOrO7QANq1ki9cU7MTL4AwUUl8QliGbad8qSi
077HWBxiRPIiWsr3gQIX7eWKszBZ4dcngGUayg46Rgh4nxAFZuwyeCVWfMwbv/H5
8TEGM5aCKtG99/p/jVEza/X7Q9jYp6gEz615XdS2Isg+LvH8KVapVWHK57igUTjs
K2dkku8hK7it1eEcp97Q2Vdp2N/EJ08CQezfR1Bm1MFiqidU5iNNC/sRwDgqhZjr
3HUX3iUJyeKqI57R0W58X1+lLYtSMbKwl9FZAd4vvHQI//AtS7Pg5zapfD2QXCVE
ATtDS7y8GRaN4l4GL4yj41FAAqt9k59axXs56Z1yeQWil/rsPpLGJKlMo5ZskIOs
p1VbkzH3ciXRDjl8MU24ELHUS5T3Bg1bTMBmGK7a0PHEws37xeNzeo3xm+tyhIux
O6sQdGMEYVYtsRGaaKFutBTFmS34XFajpfhebnS/j9c1Srjm+Xvm1Xb3VrDwPWNG
tqJBqI7n0tIi1/Z57wmxdZ+0wzu/ErofutZTnI3p7naKKiOChzPz3QjOLFBp+tZ+
rHG7JZLOR/ztI3uA+vLjen4b59EvaDhrvs7jL+r2eXGOJJ+8oFsTx/OspcpsGsLr
aC0UKvYoB2f8skAUNp+haigRUYeO5t6dOP2ayq+joJnTKRZuPQUc6yIG74mmec9D
0MJTYKZihDfqFNCwVoQH0LPFvUS+Z+UWSyTZ6R45tYNS+WW+ZjBCwC0h3sxY8uQR
pn5acjg19faX+kLxg/X8EccpOsQ7UDIftKipqg2i1CAvL7YwZTqQdKzndetUOvNh
uHtPgzh9Ebim9uT+bSWbWO6GffYCBOIcMs+UR1euw1bS5PJmBWYllOn9d2t607jQ
SO5t5MJvSmAK+fKL18Ds030E95EhQAfIqo2ojPnoPE5QDJcO6sAI+So50T6Gh4yH
m8kkWgtcpYJlZm8opOFaHWfAAMDZEY84XUHZFOMcDl4I0cdIkzUdY0StUPPfW+Ba
+AgX3Puv4ZUlS1xtj7usahuiAZ0DrsRdnyI6px49PMsbdPRsvf0QZNtqtUClwSi+
PeT8O8nRNj5bEpX+IbV2iZHeEqtLSD7IC/y7FmeWEVaoHBwEgOGc1PNgqRmH1pe9
cLr9ppk1CpHoENjzorPYsFIs7y55RyCNMy37XuwX89wqr0ph8VB3jUWfv6xHneV1
b32APMQ5ds4YjAeIScTOfr9e/yE34m7456Urr1soXWIXe6K1W89A3NwtdnF5aB8N
ySDM/AV7HA87zr4O3LaMj2kLxsjNroJxUkSOgwWWpm7+c1Ws63sixXsuWSYzlggC
E3aKuSpY94g6aJ6ohZ0EzkCMWJfffEsh3YR5cSmYgpVI/O5l0VLuuZenV52f21nm
LL/DMI620GNatdvwF+ak01CWFh4CGzRLH51OlwP8zvwWo2UsU37oOgKzOXvzqfqy
bku8RpdP9iiya3MldsYAnXXr/4jz44BGp/OhgMlMRV382pGOSsLzSrUm+8Fbn4ZR
6Wt4mG6Nb6kppw2DSTNH6Xj7r6lDP86bmH5ZGFOsVAvTs5YtwbWtIt9MChuDCnxF
t1iLJiJi2fHwFujlcx+Csqf43byNJ7AjD4UEWNmC432HsfdgDFFPI6qYoYFGkTC8
aER8WjNxsAhSgrqCbEAkVpdhrtDYlSoqJguFRCsghNH6880asUQBPo/gLsVI/b55
tUBRlqsG2UxSq5o83I2pJTVLYpTJO3EUp0uI5IitfAzI6gOofaAN2/X9WKSslC1f
/qX2Z/onLiqSWS2R/vTkzYCm45RU/tPIdZ6he7pl/dX5RTOk0LNU5BrzcgQPV5k1
LX5NqY9edp2wrmdAlsJgSbtHzmxF0949evWexTgePKcTztxpoD6pLtgXLvUWbjFN
DO4jB4q4HswzJPrJRb+LQDPJ7OXjCCFUtKFOm5gJrH1riQCioax6rCYqykATr/aw
3ONrE1EqhafUMrCVkZPqZBN+RSpML7+DCeLbgfyKBXvSzSpnJzEvyNq19G6l9YYj
+38JYIY36B/XA15BcCCyankDDXOVTxTRgkipobpCtiaX+AI38QvSnxCKFlcTaqsJ
zukBH/w2tH17fxNwAYvF3lfNt0bUGwi4cabJvIvCaWhKBH7Jwctziaqb8+CZSkim
t20coERwto1YMBqsiLVewsXb8xEpyw+8K01vaF74V2rH9KBVrtYafJMLg7u5/SuP
wyEcHPL9qK4u2PTaIOpm6fDvRAf3FBKTKSxyJ/yA5HFsubg4IYuO9TrJGRnxrXJT
ScLmndtPH85GBFaKC9CO++p4Ea0zIufAnPg1kwr3UUuwjjZpTOkO4my4PWSwt8R1
fF/F04OYFn1bKDZwSr+57ZAfSzeR/iGIg3PdVUpZVW2GEpzRAzBwyucsPzlPFJt5
p5e7nlkKpXsPHufBr0evpgNUUAE3Tn91xUr4TQtAc7D/WvW6uXLgp+VlMEAuz7Xt
GrIhoGhZee+ImLQg4ZFNmrQIJGtE7TZBHYMpIZwau71Mrx7HsiqZMA5TrDCOTeNJ
UAIbfop0kWznRsbvb0zVS8HSZ7qXvaoElQxkv1zHnHmcpRaWrqjUEOaKzR31V0K5
o5Lr19RPbZzwznYwaymcBP6/p9BvbFDZLbv4a3eIUJ9y5TEJGky9Id0R+J/0Hkht
9ZVpRc1hB7PYKIoofrXsTs6M+BvRXUtN1g3Qh5CVzpB7tYaMq3HeBvB5na2CbCpv
w9CnMndnirBprst5keQ4699SDSWZ60x5RLwLWex9eLl0UOMZSHjNBTkMugMkrBSW
Y/gP52vgnUxMzM5m7in/Z8WPKns9vykr0tHWSfp8spm7W7tQp7Zpc3z19CcoLXEa
TVpMM/2nbbxd/4OB6Hnc5deDg2IIDuzLdtokpKC0T9LOPnKVbLsvrdHHK+Xji/XO
kiyQhexrCCHx7F07s92fuI47+Mz8BBio8PPSBqfyBnumHrS8ETwbSAmHArffUwaa
guHBYskLL8H8z/RsmcWuFSVZJxFklwU7SPU0FqmJBPMXDmvrQqB4vqqX6TjBTE6p
baYwL5Z5+StfJtLiMKlOCKJ6fHkFm/WhO1YXKdcrIbBF6tEp6JleQrhe782ikZ28
cO/bmzzAj3pedimYOE6qWTpy/AA96pOOeoudBi735Chm0+p7tBYriZeewBGVUBqf
lt+IxUoC14E9L941WxDCV+MAQcLD4rccabnMY8MijUV8/Q1roV81Vs28mJwvj2Q8
1sb5AdnTKFDJ4x73dnpepfWfZhTZl/aikdQP4ftzuAtCzryzlNLNIOsCseZeT0zE
ECQb2eliOoE4BMkFE+hl0eTILvwgyY7Bgpw+UGD7OdujB2UZIOt/ZIv0TrDm5i6A
syb5CKYrVc3ijoAuCqNaJGBuMhek3qDLgV1MjxmqrMgAcn7h8jNFA5JGGuu1l19Q
FqrRZCU2s57Y/AtfMQXVu/Y5A4+XkcHCa8U6Fvi4uR0HkkSreKhd0p0Ew5SuUpEX
THS9flRzxsBwpDd1/Qjsj5+UchLLqwdDY/GpfWOPhSO893U4aSYqGtIelBcAxgET
X4eKktPJ/mkHQHnDlPb0mhzzs6K0BSkS2qRGdo9C2k5xFeXFozx5DnhXAo9pEv5d
s/XQALHqSueuUAFE1W1OP984A+woDtOczJ7pQyhQ7L6uPayYkmeGm/w/RHVX1+lU
CwcHNZPRfQHRBnYMWIrUROw5ExD1+2AcjeOWYXEz/UFGbz4tDbhiAdpYzFxxBw5i
KytJzmMKHfp/nrTmIhkACrgkAb62PZyW2oFagtqncIILtQ4X5RLfrZhkG5RLUnau
ng5M6Rdq58S/tjFHsAWOxW0kKenA93u6sYMtF7HCMcEWGYEuXKiUmDU6sTNL/jkz
DVUCTfnMWAfVjmSI/98GkYqjNFjqMr86p2+opWJky54DsChAOYfoDOIGkV7X1zus
YVglefcuY7GF8BAGIcfITLDAbtS5Y1ZR1YqpiIuhh9KdPmG7gymorAaG8C+y108m
h+vO/bLu5GIafiYgxtnfkzXaH/79S670zCQulyxNVLrSDUUpvETF7mrAAYLhu6ng
dtypr7Pl2i/G7Fhg1mDqOo8mRA3X5EwJWws7fgphmrbp113Yokr5mlqeV9c3KqwT
Vh0YScYNF32S5D1dHIVfhTDoAtZURj7ROLHxZ9vgCBuRkXDeDBieAaBKtpWl1huv
D/QzFJGsBfDoBFlNCNGu1aJoCCrgpz9hjT45c46lOtfGmSUXWJTlxyaQyDX+GwYU
BM7J7Bktw1WNjTaZtAMQkwNufOzHEBlQ+bhUXUCbZ3ZGE4Bm8c1EUSDVOH3XkEO/
x+w9d0u4G5W5H2F1/yx70FxPji8KfZwITFZTBIMTzRu0uCjg3aCCVCwc1FqOaY6o
IqeHgCd+bQM8c0x/5Mdmx541GXNrZfX9svJjG6KALr5fieM5WaSL6rFguHhw4A78
Bv0FzD1DzEuIRSZgBW7cxcqeVaH7SBw+H6hCfWl4eHET/h61x9pF3totnUc5ynKF
eYOwvfcwzPm6lb/ueB1gYjUSZOOanw+BQbbUrf5zyFvbvA+lnGKh00uaynlL1+UJ
qU0CjtXlOQ3cmM5oXqmTO9rA3J1E+U1EJHgmq3hhZZgBV8jZrfyPvhFBV9czJwEM
YsgqMjbJz5zy677ayvcB+69Hc+w/LNk+VSByzzZKoj7eLqWk6kRJ70nSpzmKlqOS
torHQaiyl9I7z0B9yC5X+6mRyrlcUTu9I4g3Phvygmyb/TzGYCi3+PKpru5QKVSE
qAbyDbuDtzFoUJ8yrcwCqRV+tn5I751QiLZVca+IIn23iMIaxTHOWjWP7uDDgbqs
+Vd/HLS5YmvLcgLgE7xzbNYnmCJJp5wQNe3KgDoHTnbWUp70+BZyma5qOZygva6v
M84E16pbaxEi7ilDH+FuiF8pniIpbmngxcksPn/Yn6lL0jhNp6sFGbcBUvMjeA+v
5SC6nfxZ4xCKrlYlmQ+cDwdBfr0C7nPnwpbQL71T1JtjRCILBehK6wO6NiVvdN6y
VUf/R7dJ4uRWprg2VS3WbJjkvqJNI0KDFns26vup5x837wIwLqkoJOMUG/fnwnIl
NllSGUNr9SFB31vR68IEDbNdRxefLICQ5f2mLFGUQVXLke43X2Qo/TlKcXkfHdEZ
zawunjgVKN4yxuyPIk1w0RLsBPOviNXAwyb7ufUYkWL/yj4Ns8LXLHhCV6QNYPoD
HQ3Igi+C04gJWF5BKtoBbwAQzPlh3eCi3vcIhuJw6SUh2jaFMqZnAbOKuNnx8Ug2
sZe+fXxqmpl3dcgtUcfaoSXQZul1X6w/3ffKgzewU0xmJnSBTpxdenVMeQprRW40
yIB6aZGo5vZJY18BWdS5gXYXx3jJ/CXFkz1H/BC6mi6W0I2jAlUiduZwvyYefTKn
pAahUARET4te9i3edfbxu7dplayEGkiqicoca58gZPsFU31mQu6TU0dACQktshLq
kjh+5SCjjrqfFGtIyXJZD4EFwKSsqbr280a6hSDBlWTHplIcBCWGkJ6hZ/A1nwIV
IbQr26XyRdq001OB1JbyW8yTGCfnbiTjaFmXV9v4X9Owb7ZqVODIb6R8TFMuTk8J
gxBktZr+l++IxWRrWvCv3+krxtKtYg6CU7AicvSstGt+qJImTumaZ5wziZWLT3Ha
6oMA4vmZIXA3617p/7wv3dscYLzqCRiqpyR5HeaDAFikK7DNkpR4cijXxcDiF32Z
dAhCpmtqhqC8uIswETC5Pxtw2AjVoG0+rmXpTkpDNIuRG1h6M9tFjutcraUERUeM
+yMhcmzMpepYQ40wJrMMymX0cdKvbG67ni8ohHylobzV/fF7iakyTmJK9CT8XwT+
mYgu+62oS+SXPNyrMq3HwpJWfUZ6+Fh7Rmx4batV47hC7a5arNh1aBwBB2ra0oeZ
xVUM7A28uRngXKsR/aAgtmxodhI5stx5AXUbxRNpkhf6BL8uCvCpqk2FHN6moRaQ
BX8psYEwhvAJJqlJC73teNOaDcZ4r0iu+8TgG/cBdf3lDXeBEKv1MC8zgiMylo+Y
LO6hSUbxtrW5w+tkKsgjWKzky3RQBWMioSYsVpi+mrzp+FWCqDPLVJILx1JaFzy0
tl/sRLzZ6Krl15FTgx33RY0X21f+6Xkf5e4GLCR+J+5gG7i2xrb9kfd+1GsoM0fi
7KPiTBWXQQDrHku3kjbD5lGvcHpny+SEd5y1XlBl4Hdwsfmzm0uzDjVa1neJiwMB
YSe8oNb2EnFEIgryRNyR3F3gmZuBf64tGNXdkBs3jAoJ5+4QWRtYgnA3QPuYuAJj
j6lpHHV0zma4nyYdZ6WqxXpMHCw/dDSOZe/jNuYuo2c8xyqS8bxdFwhKJwGPYeRZ
99Kde5HIJYdUvLlUe5AZMU1+GW8tzHGoq8d8oGIhc8FBangFD0D2BI0fhvJoIs2O
u7FU0moOaxt4QwRbpbhfUegr1hH+MyULCNklgydHyOqo2x5DVAdJPvdPbykgFfVW
h+er9kz+brD/FL6/kLt6rgvk5jcDeqQaLg0XuItQAGG/NUGHTLb7MIoKuQX6RGht
S0ELLGJyuivdALos3p88w8M/+77wI3KsjrCYGsk1RYoNLJa56+v9U8MNdh04GnqK
N0eOPk7YEtDMFx38vnpnl8iT23O3WKALkRcrCXkq8dN1nbU3CJq3KwKMQPv6c31t
ooLHD7vrXbCGdLCzYAHVFTK1OeM9gOsBkeheSWkGtsCFpoZZ4LviGm+h6Wsu3q3/
OywHAroy8mB9/MlHpOKQkaauN3i6q4s8BkKmw0xJdj2bKNSuzAGTlbvqhA4qJBRP
wqp3vP4lI6FjydU9u0DxwfxUQzlaBZCgQtT7WWtY+IZuQdeR5ycS4QCqiy8gZViM
GT+9++gpCtorJGHwZk9seJpn6aDa/T3ZSdTarpjykei/jlLlmibfpU0C9oDKrzsS
giqwsPuZLYUe7YjE0BDeOuZOkQmVVMcf2wQzU12owd0jr9nPBzWoT9kiFecteVc7
4wxeXKwGTGrLHFxhHbalZhhXx1iQ0YVDuAgcwXHKAY6/KpEnwNFE4aBu2CFqz55Z
m9EP8G8nwPYRCcT36G4e0fof6pt51eQikaNE6aMM9la40Q61BzhiLChxc2RZUNRM
rSjhyOMDsXXg0lq1EN6vtX/Kh4YKmqXvZbm3LPXkC7uyVEQw3VaqsppCTpM7cCCW
M0uZtvHjnQHzR/pmKWsYx5LoiowtPds4AwR3RA8KkRAaPj8afqRSDLAxHtQYuENU
TSzzYL2MER8F5JdD+fNKY7/Myyo6/Za3L2sehxJ6WuUMbzeYPXXct/DFNi8XVoGe
1d3IoeAjcna2n5unPinwJll6YgPNs1rRA3kTlvv0xGf8nMAYLzaDi1vNICwZMQ7N
wXyS1BI0PSORGGbuk55jUZzmLqg6gOnl9ympA1Ap4kEXWGkwPQ3DKuwPCMbmIaab
XCLWBvacjQXMVpKoHNhNyZYAl7x/8BBI5cuQMbgVKO/x+wCJbwXuVgEUsOfW0T82
UmU1EkVHftPDnFaEdNNtetS1WS3+4lQ6vCcUG5dnx4VFRtx3yana4WFETEgVddLI
E17t+dGuSqiTX60uDwUhAOpCtwqQlqcbmWyV3Vo1hhMh+hMkFDr35+Ymj2de+bim
2GWwy/AIo7+Fs4vs+d1kN8WvTrRUewWu+ign2bO4uJBa+29jpCSGZmtAiWr8ss2G
aYedHo+o88wy8i30fSJR58KqAQIEce+K8aH6/Ss5cEhdDlaYBftpK8vaQVSrpZNx
hb57f91IGDelWrHZDqBUfcElc3YTNl410mLSe/6rSTcWPhsFS7j72Xm3oE6GDySJ
9WT3I+4Z8TtLWupeD0GPmbUkgZ6YSV2/qxXAFIbj8Xv9pHVFna24JVhrP5eZxeFk
4Xw5/2ycWbwJ7HW3VHyDwM9ygzUp0ravVWisHVFbEOzk+VJyOGrI74H9h+iN9iQN
5IV6fFVGCNOQC9TpbEy5jaLrIYDTjkzNMOQ5ss3NNgYYHO6zMmXmClGmKqK4Itgu
sEiWtdkze0rHc4yQVQ9j/zvaBdb7k6//7x+F6r9z5VLMp93z/y6FiGdQ47I3ja2n
WTYXBTdKwkOXRz6N3q3kj2QAwCEcljJ2/JZnhxvhmai4lIvFbGt1ikzfysaS7khP
A/Q97LtU5XHE3C1yCF95+cd9ykVfixnmy57G0Rp9ITMEcJ9B9+1xRMcXWBo1AqCO
+vgBVDMAfsPZypXuFsOeG0/XqM6tTVxUqBxibVXAJgJ+9l2VojKPE4lxfsdovXB6
jZAh4q5wXxUsNp4HFAf7S5lBnNvOkyo6psG14/EF16uWl8Qhen2ceBoAfmZywuna
n88wSoLXxF+LBPCpsvKR6jFj3iiPtdHbTiRZK0uyFdBdxgxJ2izb0wtNEASO5oCJ
pJCep4Eo7YS39EqLfasly/UPdRqwMsCdPtEe7KvOMxcm9cGMbMDMflk/+ty6Xz3Z
AxMVHfigCF6F3wShwuAGDkjKN8eNm+usgpgwBkobdCCktaXp4PwvzY17M00piqiG
+JfVgf324shYh99N9RSP6QB4mdBQvMGKBzMmTRBlrlavqKj8ZjSuEGAE15BJPzaB
cVW35D7OQ3/H/RcvvPjPjJoPFnkR2XTCUcs0RYxuAA05EOvyuB5Mu6Y5nvxhXIzt
IpnwnC1+GjLXaOfXFtL+3QRe5Z+ii5rBMir56KOLUu5l3cUYrSQDMLBzO2TLdrfk
ol6CBZ4LGKs1KvV02wl6P7NUHCTlhrSVJFCST+dHX05S361I4CD196KL57vIgaPB
SuFgaCmwT7qAuCgutM80+QC1EsbkEMZrznGfjqYe+XH+p7BuvmyZakp8cZeS/34R
GwHg+ms9JEChPdL4sElorBvdzLOFeX6MWiSvh8Cwpr+nFarZagcAQOLzciob9q4o
UnjSGSeJaheQxVsIuv8JtIUV7aJVyK7xTBU6uWylASsE7OpPJUXiKojfrdyrWHLy
5pD0BYww3HpfB1b5OE8Pi8sWuGQpdg3DKOlgEhmRucq+5D86x4F7J3pE4IE5dXZM
958xn9EN2diF5DAxz4QZojA9TiQFTXC+Xb4TuiIdka1b0otwulqL0mY/u3htx9Wc
7/ux/5qL7gTAg4bDiefQI4Ux/xrG40qtfPd5aANlRM4CgddmrgPHqcZ3K3t5lIaz
VFWVxZDlNNhLm1KkY8BapzYHkGuFAjJcCFZHc/zmQ7iaGDTOL0KgcoGLpQxqE2U6
HcEW7eYOGS8OBn0MdneU9oRoImEArG9N0C/4TUxqKrEADaCNd7EiUHD+S3ckvUN4
5Qoo9PCFMhOKHCNSK9Qca9PdMcD8XoihHQY8buLD2fDS8kfAz6REBMj4jvK8LJEC
KutBtpqwLxWtCkMnVuLTUIg2HIr5PXpt2kWzm2jk3ZApmJiMj7Ewj1yZZQnCm7OV
uOcBfir9d710TcNSeM3vMFeFnEReUzj5WgZNSMFR9WQUl6g7k94XhMtWNRlyYhWk
Yso2S9aE0BE/KjEfXIN5XZ4Z5YnI3tKsGJCmtagu44L+9PdWkvol4Gcy7ghNz0Rd
rPD0Sv24klR3WSG5sh2ZbQBtsrVkHQsO7sOnFYvxwuWjxFIdWy+PhRcVCpCe0BR0
jZoXMqCN4nYynZBeykG0Cbm7GPKNpYEumWl5z+n1id1D8QPUidPLEPFJh/Kigwqr
yanX+cLxBDJsLBGYfGhOG80YcWoG4GvN5ETxsHOpBUg3ie9HX3YkowIioBpK6blZ
DKQWgXL6VwHc/bIFfbk0YUDxJmgCyhsQ9qsK3h23J4n12psX8xQTbakTuXEc/Ufd
j8+VEyUu+GvviVd4JVqjx4VmU/K6+bfgf4tBlu2GGEhKD6DahjzTXzMvKT5rr1cL
1OtexnY+4QU+/twLulW+W/QHqAPQUf9EZmjSUX7osV7LMJcvZJy+vbl0bPQU0qp4
PyZ+h+dAq+HbY7mimr2fO7QWaCSXfTbwyDUdhBl5kfI5Icf0WkXggxT4Vypa9Kga
onIsS4hYZFZkfTyCuCbxZwE/MD6tHzfGqWPaECqPtDJJf4CYdcsDgo2iCBVG09uc
8E8CtVEyaqXoYTrNtFM1zy2T10v/i0ExfjXDR9z4HEHfZlJlLsQsKlvbVd6q5E9W
kjNL4dh8JG/xpdFdvxU6BduGn/iSNBa7ApX3hh1fdVFvYkmpmYXAer+c98jBHnzw
LtwiSQQf5i3Bqq8h++crldTeY+QpctdWY4z/vATFjmMi+3TVL9GpOtj9H3JHVwMy
TEljc/xPZk+mGhFmi5bi99gUI8qmQe3wUBTrXYQXRk/krks5RCRfA2BxGvOmJmga
OHeuaYXsa8NXxEJJozEmJHmBAphuCogksJlI+ueZUwMyiJeuIhc7gdVWxNEupuPz
33xp4ckCDj/IXJgqS/RcdMnJaroUtcN6duAjKC/7Kj/EnGxlzYDhpivDYS2JNHUN
GEKGrTt9zHWH6F90vtPe4mdPHfG/Srg5pKIdgxu2eXVL02fp3UOXunoSo+No9k6j
vu5VPTOTehG2bao743S7Mn1juEj0LP4nLohf8LeCJX7043fh8RQUzij3FrV6ovGI
sGT7sOwDUyvROBw2dALEYxbDkJ9/kzlVigUUKu9LqxJee/dC7Y+a5OiH8XuuJKHb
6SZkemZX3BMKDiv5F8/a9jFbYXbNusZYJ3L47Pa1b3ZDLCM/MoAXg0UPdC27XE/V
c3sUoSviaKHQZHBjYm+yghq6EKgvTnKEs8RtwuYO7YUqoTIZkCQjv/hJOjE1XWme
RI1Vj6l1rerErmpkfJfwlB2SxNdQJel6SdpL3o9E0OvhGy4r2M4PHM+a9CtBSR1h
RPkRTbcvfEefnWzW5NCwhjpN+r5HvsLXbAhjex14VSi2BVTfGO/whSZY1Tu4dvPK
0FSs/EmquDZ0Ac/W55PJq3KAjSQRkn0MVEYHJhnl3QlGnQHx+JlDQc38lleq79tL
tUwY6pLY250YNBwO6IU4+7SjkYPzyOBNYwO2z9l8pRKRtcnaFWcPMYRRB1kUGmEn
d8HdaMay+CUWcn9j09zcGqdKKGsyyuYNf9ibvXF4mXgaMzDSiAz1Np5R+9j4CM57
X8Lvp9qrLvfAjR1e1zXStANz55QawlFjknZY0I0lsCKZ9/Qu4Yw2cJZsDNJiS9zg
O8pBdPsFL7BlBebp/S8RYA4DPnsqWJSLCWxgESE0jg/CcNFn9A2hBP9g57aN/z/f
2iLY1SvBbbH3CUfwjqCCRKi/pEMXHfqZsJxGNV8j8omRsDprRaNTrIjvpRbgDAW4
yW9whQLlvN/ABRSPbWHK05PfLYGEJk+1xkDpueP9RI3MFIstQ3SekHkd+rGMIqYA
y6vw9tlV/rV3tO0aLxR1CyeavwM5Iq+sT5RAi0oBkNT+nl3Z557vH/LtAfUqK/uz
zKpfEwDseHiWrx4344a/wbZ91u1j8Z6qCQm5nimGdviYsanrMlZlTmOEbwnkTmfD
H+RE52FkTQApSK6uZftCt+0jCkFHYIePod+uZ0XmLsp9j1o8TG5MYRaTHUby+8cu
9mTm9CZF6A7cfnmL+VYu4nMs4KORbd5w6q4RAWmwa8xSq7DiFrPb9WhlGlSxg3NC
z83hp91uVXq2MkLiOD298S/kxsEo+MbutyfuZr88+UR6jTibs8AP3MDvznwQqB4K
PTnCNFGfaxPk6BxEbliI8Ilarg5MOCNN8Ua9tlwyiZFExLPPbWU8mXx3uWQo8Igf
PhWiFP3y40FVEeuYnkc3jDephGkQ4t2wd5r52+elJJoKSguTGBXZsD+4dOHNJ8bb
juSgw0PiFv/m7sjPVDLQA1STn8aO32Zjphye3grVQk3JoF59v0iR2HLAGqNVneIn
lIs4gq+azRrGs2tViX1RDA1RXVukCf9lFTtzMjfOxwCD5FbcloYtKHlq/C9/oJvE
Y6mBxpFt7cmmP65DGVE/lM1+EWJdvWol00PDeW2zml8ZkQihV+j56nAKLJnDR2NK
fCcjuKpdeKtC+bs551TrGlVQo0Irs/355FhWNWC9qJCSucYzO0/BSlOzEXUZabba
hr7PFXjYHN9j9WJQ7FFEIwOsMyP6VFrBt6ytWcKA/mzkAetnh+NgR1DPFpKQ+SYt
3uPdK4AM/0t3fyCrGs9v41DLrbRvXb2KIyKGDLZXwbJKv1+5x3IYwBSK1IE9i0Iy
1LAp/AbFt8KTzLDG7Uz4y3AvAVwInDCHxpEj3i2JahRSirgtGlTv0ZIDsyci8IOz
iy9awdtzr3VvUqOG8mk//hifrJf1yKcsj8r6geYXDdwPYEoOmrtFS0ZjRP0QBWa8
QjYfHFW19qsTh7qtxGHcE3DaL6BT1QL++ki3PImCPxDU6FGsfqlFAL8cRsnLsh6m
29R55KeOeFzm5pyNH2uTV9o6J79gZbYVj8NI4uC0I5xXe6tsYiV0UimKPD6nfn4V
XPlTLTYK3yQtxD/Y5M6VLZH9h3nELCnRB08xiGuX+b/83OuwYD9Z3XhXJ/e06ozq
4JMrk8Yes3YSlXPDC+FMVhCpKJ0iZj8hyygl2WbcVG7UG7RRBl3Rt/SRMzet7+vv
OtldsetsuYzTFq5j8kj+Z8G2Ui0UsNkbyGkeHrnuHFl9EpDxpeLkjh+vT96rokfp
gCfIqwPu9mng2qhqIwNXc0M3JasBh8/sAX7Xpp6TU6CxwEHXkwVjE3nhk3aIiCG+
pcc0fVTJo7+LHUV+mHNyGpvaLq4zYtwFA7txvASw+k52nGOMDx06Xqf1W43SKtG+
bLFzGXEwdKFfmLmVO3ixXcHaWgqFWNnmVJyYmlmmdgMvmufErYCs85UH0kPePuPI
ySvW75WrCHbdrCeb30pe7ua6xD4vmSSZKm4fm7ixDJLXcDHJfTW2+w701FmlvqX+
a7/xJ7ixqFn5HyMPa0B4gyLx1XT1q52/FkXQdxBPOha+KjIgvTotaFChAiAhBEd8
reJFzModF2kkSUIWr2KTurr49gmchGKKeTN2OXtp5dExylijJJE4eNAUH0XNOiiN
CTio5OwbBURc9ZeeVIA3flBtl6pFgFIeoZ+eWAdn3tIuVNQ93nP5qTy+zjRDNW6n
GtO0azNYNcJ/Oh8i4jUZYMfS/yk3/WVM0y84EupT/w+MDXy+MFTkX5r7AMdCT+fE
sMVwGUO2f1q7ujCZapQI8CS28IpYrGdXiND9QtsZQyhzscdnyD4uySeSaWIlEQIw
GelqsNCfsX/dF2HAqkgwOnPaRtfkkEsfeosntuy9s+ObcT3F6x5kdx6r7N73k/sm
lXWsxwh9f3rIT6wyLQy96FVxkuQ/Fm5eIN+KaSDo2cburKx1Y0KBUSwKn65P9Xby
b+ekcPSmUrLXft/dovwFtsnteLs8RWS6z5rUYxxuJd9ODlPfF3dZ0XntYj+uiXpB
qAasn6n5K6eBbhiuwiDIMraK8kopqPIYXTQf7GJoh8deY6Brfrt38Nv/GUGCkV/h
op/lQU2/amc8LWcphiGMXXzdPjjHz+neHs2GbHdvqmrBz1auuRO8oPOmgSM1i/X0
IM2sY+eaT72pytaoKltDoE9NOGuzivrlmKVdu6CkEvScbjyEmncdFNzwfGDy2gam
TGT2bpCjGWCf5BNfUmJITmDi8KI+L5eVthy++6VJxNNSJfLbaljdCbVL2J17yROZ
x3Ovm2ENIuA6aAjz15ok0AQZcxFHHu0feJcBw2cIi9FqcbMOqxdK8EkdOOPE31dZ
eBVWNl4ToX8bIjO32VpSSnCVkQgvB3XRNiVqnTbO6Iz8aA8RBuD+11Z5FuELsaeN
czmIzzWLsaZfqTM7zu3hqg9JnDdWeJbm9KrcCmIRHrVjhAoE0hoa1Kn0GiVcTMys
/1CTcF1wnGvGg1xS51rOMmmgu/adJZ0l4J54e1OdLyAzdk+PNmEMMNHrAvywRQ6+
No6XXh35Lhv+f7ZMtTwhRCsjv5gAIag+3DfZ725TTM6ZjlOGVePGntKxa7us4MM5
DUvSe/pt0r8J1FC+iX1oHlwLr2T1KfUvgAdeFmCR4mCN8Fr8yL57OkPMqfYxGV38
7fE4nYO/ZPD0gC2tawGhLaixVW+pA4ocjjHgrUDhTqfog3lV3jBx7S7vauSWqG8G
kafal9EEC91ThSRlata77BmYBTojjIszcPbJ6mLbsHfKE+K+UNl89QMZngdT3jGs
OLvYPzU2jEvTlJGy8/8zE4TZllCrCBK79Cs3N6SB8xZrX6fncUDew6YL/ZyOGq30
n3iSBYHZOBHFQP9G58UWFtHKGEzb2pPC+RkJNyTf5lLVfkEjcI0Z+kN/ytt/8mNx
UlZP631T2NmYwcrWIta0LEPbkAmwHbb6zf05H2sanqdpnwaeowsBQKaSigPQlANu
xYKGaqfWY/7kOC5sLU3NPSTX7jOwpb9K7i0sie1DKO5U7VaNXqhzazTy5AhfyLK0
4uc+aHaQRKRuy6tbocWnshXpSIV6i/7K1l6bcyEb+gXIUsIMv1pTLLlru9MhANYd
yGicXa8d7J0btPTvmK/nBdS/0dvJOsEsn9aL+y6dvxI8r89t8aYjU+EMeM5gyDxg
MDc7C+ZGRAU9QBjUv/GQt72qADR8KAGZhldQ73PL1RDPn13Zayrvp9EeOSN5Avxu
f/hbij6MadBriSJ4oTVfKI7DenauoW471ZDCggOKsDJVS1Doyl8TVRBdpyo99qb3
B4triztlx73cm0xuUZnWPq47rAio4IP1FjRRo3yu+JvzQyYW6iBY8OrVM2JyO6a6
XdjY3hhNWQxmeYz1RCUI6Or+GHXVJ8gGDa02+Yop78xdSk6g5/x5sO8k8G3YZ0Dj
QXcmoli9N7ugf09fbRMmYOk3+GSKLmJ4QZLJ3nutU+G44Zou4miEPJM1bGQ3gHkx
JERgjQagVNcNhm0Yqfb20VRJ4AE1eO6mbEvF5gSCB2HRY1KBHS6A+W1NCsJ1/ZiA
wZ/8POYzRg5ZbuLH37CNoostElFTcYEg8HiY7nfmu2IPXmDyigbcNq4FSAoHm4pP
Pb5w2RT+EqU2Bhexl3eY8qt7LkWTRKN76Ai6SFMhESC6N8a497WndraOJehuY1YG
ZOmzOZeQ3XmsZIq5MzPvaJu1kbkB+xTtIdbcY7+w/uMd5xGxvYPO57D77r3vrn9W
aiuDSKtejqrIh6//YRlzyqGR4DpZ9x3mErC0DnHCJGvp8BUOJplCL10i4CEbVN75
yfmILpMYGru+Zj/ay5Cbn0H4902kYko9tDvu4pZMbGoCRE8Etf0/N6o1Qkjo2moI
OHQZHmUfI342tLZw1K3YjPDQpWKvI4qGloAgz6m6YYTNcxDko9uYzpKA3VnWK4hW
w7dY742+UMWtLp7bpxAkqH0oGnk92SWeQOFg20K75wfM1GIOC+VjitEQ7MBGiaXE
8/g9Ij4Z3MtEAHXu2xrIiCXvbU3QVBzgwALgoLsUbPqxC5MtrSfhgDKV7OlW+tX9
OBNDDPeMEUZXDhibDSXawzVQJuh9LK3+H702w9odCokTAW3kRYwhw5cgl7KXn3S/
hrZlZWgIXzfLq7mplbA8gtlCyQBBKkKvXwCu+DSGdM8nlCg7oaGaoIsabBqdbn/i
OJPdNYm6aQUt+lVjSXhFkaeLUCTgKwWqsE6qvupTo94GOSPmDVnIcCrGRpcJa+P3
BVcpFCXT3Kl+8TKE9F7RVVcz/kiS3H6Wef5jV94lLETUKCHoizDiS1TmN2YuzATD
sX/4dib6n+xFW9/bEb4NWxTl8d+9Ciu+SBkLjnayDncM5scO7cinuN+rI9tChjZW
PLHkCf/DGIltkIyOniupWkIFj7X0yaNOHFppeMtivfEO3soxO3gS0LAqzOW0tElG
X3JoXk0ZtM9/Zi58L+Ux6GNIIQCUCN/AKLL8gWegPbZNYlRSwvOqTyXWjwqoFxZR
qifY4aGhpD+e64AQ88axx5yrsggzziElMgOn0XMEfffDl76WKDzNVAfyeQVM4PST
TSdHXnqIT4RzTSkOOGp0YGjsthxeuJphaN1kaT3rtGzL/C5VJsRREhdK/gglnxgv
hqcKSd9OqoWthJPiMHeK01MMARbGg7ij0ZSkkwJTqrBH1Q5Cr74j7kjjUUkY3Fet
WURHUOt7Xw/o5qHNaTupE95yJhyTxUVcXgJVxvmLofMh0hSSXKzTXlHMS4TWV976
VylMI9OsvlpDYnu4d0FMkxzzLylNpl3Q1e/uAUW/dPZC9TSzPZ1CikUbprOysxG6
8r9KboP/+s8ZpOmIzgciOTA3QqBnr3V3Z8mu2vt6o+JIN8UvFURL2js3cnykQU2w
qwOBf+9e8WDFNbOhmy210tLEx2IUr/SvxCaLpM3JdBBaWJDzsyQNMyp3SV4eVG4R
h7EOHDLuhXL1t48maUgRY1RHopc1NRf7QHJmKwM5gnH00rkSdOSy9xaLrFEJL1/b
xbWRsMJqWU83rV3h+f4OuqUlxUnjgjG8EtRqR7DgrvkzZWZfECG1r0lwx5q/ATwM
+NoSOPzKdzVSIhgmosyfIg/yQIhLzlMwouMPoWz8N/pFtkfqEuOim2BFvajkD96O
khQDNQVgB3LQZm5fNJoNtSemEXZjtNwA/Ri/Qh8MW3HlW1vClOxY5paY3OwOb556
I4W9xHtSbch9WSviDntggDjHvXUh9EMe9bxV+dEq7yQ9XR+/gIMRQm+1gDAqDvVH
ukczXAiHXsf0NBR51l3Z6B4uSSilnDfCoawEdLg9S3ZpkCqM6d/6rtGZB5c4EojE
G9Ta7YO/QRGPlOxrA5StQkNKJzwUMTSPJZLIyYPEbg0QSghztiVeTLzub7MU62pc
E0kg2u2CEqhj8y5p9Nw+DZaU9pxy7cuOQEjCUMHOjSbVh2N8TxSU9GOeFnDG2TnU
bxW13HNoGtTTu9bG90kK5P0eGx3D2ZwJ7I04P518E1SerdjoqdbJYWziHm64f2Vg
A4vh5hrEkUiJzFymnwBamODX3T3aJZCEhuaSSTHGNmjiz5Fl4fGzw9N2Xm7Glf8/
N+YIcbftKqYsRimLgptnrEnwU/p9YRQAQNuAfwHvxeW5z1TrASxb/V2zwIDgMtSD
7aXeDZHyemKlMRTvxxsW/K6T3rhQD2DmXPyaE2ruP8YQ9XhwNSbLKxPEqE0dMfi2
hrCQUq74DZHSl1471lMTm1YDe095bRrKaEztCeJ6kxkR1aOCxdLFwXHo/swwOMT4
llM5TNqeflHXDAe2/n8UelaQ6CYzc2FokUBYEUCzh9wnLK01cUdP7NjPHuy0+rg/
+n+/mXTohOJ+O2E3UTnsg+hd2xSERFiLKESMOWak8Cq6cZSQ0Tz7hc+462H0iPlV
S2zCcFqUyL/sxIwDu29jLiO/1ck5mUZyX11c+Z7Dbzz40GAdCCJqacW1LZccNkJi
XkxzCh4paees5jhfv8nG+HO94Ho8YI/ogu6UaxoLWAUc7S4k5HDAXz0KFtuRhdJA
QDQM+j5WhseYs6ebOTjDscDv0QYp+iAGH+inPwDErjfbD/zTOT3Rt88MLfpprX4V
TWe9uI9WHP035csPrIqFtZOYESQmgSwZ/eSvqxxwXgfi4qSicFu+eIA/Vd6OVcjp
RpxYzqOK2mVUo3y3Db8hYshvEOQzX03UKThvfze/IubPitbZRMPAeJUmQehgCZCi
Pzsfxb00Sdz8z0iWXzaP/zE8UtDddAZp9OD9LPLEKkf0HbQZ7eBd28yDB/7hmvII
MpLZ261KEzSm/oaMg16sfofJK0om8lBhmnSybIZpk51VrDK+mZ+rK/Zhl3UWo1gO
H0y/HBYbqzkjp+Hks7CiCSTQPimrx8EwLh+ZLtYW36pY8bL9ZqlOKRcswKboA7Ob
xVgHVopMiunbo/j25qgu+D/UiEb6CT3uevQKOB+QMZtuoYGKbWf4GlGqqbAhnaRi
i2yiuEUA33QSsOMNJF1oxGvct82eu5uHHruZRXmUbgT9fw33jpWPHlzXbVeNtXUC
VZ2EmjCrvHR2xryJFTxSaeKElsaGM5iawGVAZOMjpWI4pzl4PW10xXJS5W6ttJQr
Vim1ByqP9+OHkVKCaJL4PPj5c/4herqzag0qF+Ar4iHCiFLDZHJRaQtiHpznK9FQ
EmleSOlPNam+tqpBpg1L1KUVncMHSXR5yBY9jJMnuosNXHAGwLZYUDXAqXzMj2gQ
mEwfuyadJuMeGWvNLN/MnsRXNZn6kU+gvhHLlsl3hqmCFY2+OrxYXKmsd6YvCs6X
0260trfsh1AI5FzgJOV84Y4yAw1UDoV4OvCYAs/9QIb/AKTFPLg2VFUZCgKIsxta
U0SnoyGirVcBRlHn3SO+NIamnux6dS49DXHt5yCowxZYfiTz/dDIwrWqagSgjltm
55i93wAW6SHCY+UGkfxge7PZTpJr7k2yr55jaB/mPKYeYnDaach3zsWbAH3KXY9F
K5+LaFUKSKzxXqQCUdGCHewGF6HIbFKJJihb2MMVKP18D0ZiwbtOrU2FRXD+2s09
lGPDOD2xcubN7oKxsybYyKcjZ2ciXQwJDB4yrsMdgu+QUcXRBEaPZ0+COMjR9AuZ
8D46TVlQBAYz3xjm3th/EsPhDiaKIZR3AOYc7kjwAr3jyd22C9lSjTf6bDVi6/Gu
4wJdqkxE4iRtT/5VcOr1GHAMjlL90Hwi25mHVH2ap2kiOV1XvT197Xn4cqJ78RBZ
7Bgs3/XP0jdG8qeLXW8jurXHf0DTewiYuECGdpu6n18crwGj7TongsOCw9ooc5Cz
lcIAphrS0czfYZJA0Bj0VNSXcgUA7qd1m6uAWK1Bvp1Zt2tGM462PMH9C1omcqNN
o5VRxpBBD3BRraHqAK0zOjAlllpZONY1y+j/ptgP9teTL4awsIa0BKHFum/Jwy0c
Ex2oQYlmettUziA1Pg0ORXD7xO5SPSVf94ay2KzXtFtTMD2A0lAm1ih81nBXUwMc
28I6TDj3Z2iPag+MuPI4f39qvnDZhUk1wTJG0NUmpI/h4s++YJApStcQGpcsEvTN
L1jc2EdapVRV9zFGqb/WyZjlgXrte0P92w8K70/PZbTX2FsHz8Rcn3dotgPtL5cL
d0ja4U46Fs6Tyyazow6SorO6CsrWWBtCTf0WpNgUkgWUMQT431JPSZJatnJeklTp
/vdmDfLzdyK6lWrmuA1Sn3gTtfARmn7gRtWGLds7RgqIAapaXOlsBOkQOVhGjXzP
IX6wgV72lT4uPS65vRKyrL4m+vfrAXf+NsUmD2dPXgpOKqeYiyjWnLvCfU1MWLFm
IXQd8xDGFmuI8kl29jMcVotkjT+jepTQfG9CSw54kOFn9YdIB4WIIfop3bDuoTrN
8fs5qfCsQVOCWfTCr6q9XWAQaStCk6ItDO8nZjZezprrcGznREe6BR9KMMa7LE7+
sgpBHuNz9drlC5knJHxhSkfGNt/r1RfGMU4m8xLaH4v/DnsH1XP1GwS033IBRUro
+B1wq6dxBq9Fjle7iDmChEpPlD91PUBkZvq4zrfxzMlsAVlef9GtSOLiVbi9LOT0
fuG2xJmqno9APLKDTNjhr0P9LfYxd2TEPUSoO7lb4JUkVnNKy65B1eDwO7qjh6Ix
mToWvhu4xzdFL2V/nRlbvJC3tmLCp92l1oSWMY7cD4LJpcQKGx0kjMtjZky3aS5G
nvBN7zdMI5p5byRxlzflKOlHOYzYLP0R3nooyFMFF+xwry8esQ/SIUC37Y4MHt4v
8z8ccepLc+D2EUcUbz9qbY/kaKbX0H991W+EauNUh9seaC5Lq68lCSoKmaIWK3ch
Nh9VC44lj5R79r0+YRdEQMwUDDGJvsURR9wzJGqgc7/fuGUMBie9/Zd8tkTvwYCP
YKO9RHY6hF+bkF85RkqROrRJvDryrlDRGGuyht0iWlmmEUd6XSDS9c83HkGJeCL0
ucaz6s+Hcav60gFmymMpPS75RexrDIqtK1KHq9ZJRjaMXjBIn8c3SyK52GBSWolV
I5jlIbqGzWcdkYz3cwP447sKvyljSgVHuPSnu3twL09cJ9qGIb7Lb0z5uyFcMnyb
p2dKEihNFIUKZBSzApn5Q3L2ZL/9zRFURoTtnF3ksMLwQhZhKaXhaCGRFxXNVvVD
oX5eVdI2rh2LxLdRFQ4x5ViFiq3/qx8Kdqg8pBQI/rQ6jucXy/HBnr1o1Dz++F81
hPoaxkhmRsC5zokCqh0rqDdTV4utOzrXgU5seSRAa17jVlnNmWvCDCrVTGiem+3g
w73zAB+5GIovmSqGgPJ5osgLB68mGexlgunibgPE3egmjw38ySg56TfLin3v4cNH
s+76LME34kcsjm9OSVQEYZaTWLb7oOIhMCKgbJDmMWp1gWoDEsBOuN85Okj+bqXy
HQEu8uzKIAppf6XggovXOV38UA8mQ+QxSaxq6IXnMmsPfw6oqkovhDY7hz7yvQg7
EWETSw5HR/TVidjL5jnojxAvK3IaXXvARFfUzc2EDt+8uTu8NGv3xmgWj+L059bs
fXyZl0ZkaGCoKBHpUfy9Bn0gVMZh+M0oERRvQQ0PoGU08sa/n2EW5Ju5tbPoqgdo
6z+eJouEpyb3P0mXcFjvWYTARKoT7Ye3IIcyEshX2Imcl+voZuXQVPuQzJLHncJq
b5OgfKA+L3ja8n+79LAxnUz7RIl/CNIM+FybvU8vzScQMZ6yaO3jsY1PdROe2+sF
NG5siSlmuYWCYEqSpcmQzmfc5qbaTV1eY6cu+Eu+9R/L5C45m1k9YXkbcPx8dXti
bHmS9ttaZTiW3s3X2F8ND87kLftcjT9AuoPW1yFZr7UFLxCsA6laW6Y+OghBrnNq
nMd/yCfoVRZI7eKsAPAzwYVAE/X5PZt77t29apmeJ0L/oIzBqUKEZp2bYmgRWYp8
Y+SfCW3+s5uxI+GF+zl852loD8nmWTBCLpXsGXMcYf+L9tdea19L89uO82chlk0v
+JAu/NS4bmxtLqtg+ngoZ+rYEFrMNFWmjTKu7TLw9hUEYsHnxQmJ05iTYaLsqBJO
t6kGEoa4A/aQozinUsxEPjIB/Y/4nZ0sjBJMbaQvAFN30ls825MGeM/mv1O1IsS5
BsEpKSyu2HINVtr+H3dquaNmjxbPJMY17ak1yiMn6xBgkDuvbuVCeyBDTDGsJFrf
MpM445CL2FjC2ZwxMPzxS4wTfN5A3Rb3YWb7TdxPmRjr5U/pRdOl1yumQocFOgPm
1KxHZjNdZCDDLlNWRbJ0Wl3WffqmttqEUc1XLwxjYiHOBwX3uApyTVkCx1RjHoLj
IbsyCrxlYKetvpJllM2q+XY67eXe79GmMl5OUjS7hLzpjd0WlAr+6y3n3fCPn695
VdwjcfPK358uUTP8EGc0uLFnhRyCZcdGj8F9owryouViC18xt8Ls+hVgLS5Ub0Oj
/t4XZHYaopfaWYJr7X11wIKJihpK+rWI21enrlvA5gXBQM+s7zk6jGlNXXfYxQOs
HY8yjxk+j6DLOnN0Mvjq+z9e9Hqa7nAJNXuADEyu140GJi7Y8sHG7/WfK9U1psY1
P4o00doh2JoTg9yRD9j06X0hPt2tQDOkYOb+jjpHtl85lEm7jJpwFPK0fclHvFhT
JDKcjKZSNbOFAZ+AnKVwCnn6qbM0067hHXR2KF63t9iLoYxfg54oBMgsAjdQUj3A
wGkUfvySYxVwiZSYtYf7n8ModLiRi3ECiMZI9gfMnb+Nnh+9dLFB8IzLhvj03jFb
COzYjr22hNJZNGXy3JMJoGl7JtD+XAaJP8vkG98sXbeAttfeaOAfx2AIV4w49zvd
jZVoSy4sWDObOM4NJs0Y5cHQrTHu7qox8iQc+zhHsPUHh+lHCURcY6OcscwhogVE
kQJkff0UqHmKivHQkJP9+NkySkwlAzPrZOpkV+pFvELnMf/Ajekp/cx8xrLE9cNE
RJvVe2PM0KkAYba7TyaCpcKEaCTRjeWLqvWwD95Ch2jte5XSQ+T7c3LtkTvDYXlZ
FQWXhe58e12xsPdV7T3Yvqd3iCZCNrMuW4nBS0oAL3bLLw16h7uEGXgstjLcV65Y
3P6E7m94KKwJCJDWx3QaGokZvcA5mCsCsj0MVTGLtrOczR6iMtdNqREMojeRBisZ
v6PJwpov639E8a/WQGkWYeOBlEClwGxV1yCT4Mmhv9H+d1jtyyCqImLZ3E3H/91a
AKsrcvW23g2iFaJBC5wPToOq52/OUh3OUc2eWaGss6f84PZCt5FDy1vAXBcjyA/S
Og8ICUL3aaklbglQcZLJ7t8xEr27f3i0A/vpfssPFaXcOKwLj9BKKRwKYQ/fcxDF
c/yEuGACoywihQK2eGAIgQh7kZpsUPmGTAECuVhrgrar89JEmGTfaL/lMyHja7CY
HIOx5772FCbk2/2S7tpizQ8XeM5ypUhWaOAFbblOwd/VQdtefzBpR1S2LTijnIms
1pYSRucbQ6mxu8ejHsZzEOmziuZJEayNYELpXYTkFd8x30K+jB8eQNRLenmbDzEh
AOSH4+j3vbnndN8qvwsNIJ4UKLcGx/axN/S9T4UG1AiKNyIj8sAWdncgjz8qkdsl
Rp6f5ot6BGAFjGMecnN4afNer45I0+FFe95cJFcui9MgAmJ8ASFhGQz6MZUukz6A
0lTB86HzRdC3itdJjYNJU6FPI+tKGOvdq82ZMkA6sJV/WS8C9eWevhrW3LeLTzdz
I5rdC5kbHKS4uoWrL2Dv/9cCsCCPafVLjv4qWRk8M+dXPbfMRhjH4IE+IDcZd159
wKMg0CDmnFYjT/2Q1GVmVWUN4I5ZYJEFFj5AjZKblsPFrEqrDu8eTU1/2BIVGCHu
5sXFtSoMjYg7s/Bw/IqU5yDsd65JWtmGRElnBCoC6s5Pwz3PZWi+ZgIZ8yCBbvGE
x1l3J+0Lr7FbkgpbfhMSpWXmpaTkOZfQhwd63Fp5SlOk6QWLzp3xhrtR9BEUcWnX
WZhtaqSW9+7z2ilj4SOVn84mr02Co1Mxs6Cx6gU/Fr0HdkZLUKGnOlIn4cu1nAej
xGHX9mjmLg7CUxyCGiX7VnxQou8pW8ibgNACVJRrrY8uNvNwo33dEHDRk7FTEgyO
aKNzI9XjC53drZdjyVy1v0BSftdAtsODKwxaIs3tqQT3euCjxbl2X3XhopyNufSy
678+JB9kE/SAjjAKJRAs+j6doZLVZxn4BGOL/640NoPVqev6gzQSgSDRv+PcYTv5
PHsjml8trZOkV+hzkHvWb5KVhyIjjjbsYqtRdrQZKfM5BFoXurGCsLicc52RS90O
tPth+zlH56XydQXh5hU24krcNfhhUmrPKoGYjbFDeODlzElrBzbrjkzs7GmwSYyJ
KjTrSa+g++p/RBGDDK7FCLBqI++YnONyOLrAm15IoJyaa0D+8aNfa3KrRlHX+UcE
fYvG/EjE6PFuCbRYVSu0Hx0z7YXDtYFaGkyZSwblgLpbXm1FJkvve2FsezqIhd2D
EqLvln+pwWxFm90ZIanq1uryazbVR8dbTSM6GoXxpTaD2tx3+hxtWmrsqZz454ww
4bdxhecCh4yFw3/ormy81PlwW1UDa+NM9yZmYfWbSEs6zPEEWXcrEQVd3ybsYSOn
vVib5DbcnW45Mxug4lIMkcfElANOy7tpA02FZm1/3eBmocg7Ces3Be1f7ndY7HMg
qY8OPD9eBxEa/t44RKrJxJbUx6smZaQDdehVHNWJsMgVA35VsVJYb1F2cWz5b+xs
pw3L2KyXNXOYrDDdlnvYO5yackmDz2iK1fVMXIzZ9XFBjHJwkiEJfiC5mhLXUWj3
J43ZKBthVnmI8dBXPSKBX6EnW7vOLBif5+Q1pVVhGIwfloggPU/Y5rp+5BP8PzBI
tDaAWAUBemQaI3KZy3NtJ/0D5Tyc8N3aQgiul3IubiPwGqyYe/z+r8BEhhOHsqy+
CvBWsvm0RusiBATo3iWyWJZZwh5aeAWYCEQuEuVOYwT5ZpUuSmftZMYfnLbiHdxF
o5J/7JvjkeJ1S2nsvbPe9XMAclysP9Bpb/XGMaDWwp0Dea+UKx5W/G0c2QdQyKgl
qIH7cseC9WhYLB5GtUKvbRJwm6cIwmfiGai8uwF9CxaKVdZRCMt37D+1hf/RZ/V1
q0Mfxd7CQh26Hjn7fqGbKBEBCZiqOMTwDLK0V+nGfBMGSpmQ3IesAQOGZRexaA74
Yi25G+4gtgN9ixi58oFnqGnsCYTHXYpgZ4HS7mIhmg+M79vh9KxQniz5/NYNF8M/
TPpGBQi5ak1qqbl72Fjdhhpfn9R2hXHoB8k3fdv44NhWTE/w9+X6z/xlGiuMt6Eq
ZbrJ8pJHGJPJdPfwJ7Qh4pETdvYRsXcR7UcNwadz7AwhfrSHwFUp6IWegDqOOvUM
2+hlZr0MVSXUBq+o6uJXyayKDvqHscrRH1WlhInR8Tao1AJDNBuyIGNekbOh543Z
mBXR1qjD70TKzf+gmYC9zlSZJmHt6D5k+byZJo0xTCoSq+1D+5G3FAKlDxCuRlUD
v/xLUC55pcVXE4N/dqLX5v68u9yNNo0mTDSrm2coBUWrwgJrLAoRwzU7mzFKdyfP
8W0PVmRKCoZTTFXNPYjCmAQYP3PWZausxOg/dkQh4w9K+UULX2z72ZFrsDg1PqW7
DH9BEdDtXfT2rbgAonye73mKuZSxBd45CwK8YY1LRq1RyS+ZWtXPOBIP/BhVtOVw
AnAAF6UJc8A6Y4JzZefxls2w4jftqeAKa8zGxUb+1dgrMW1knEgtg5jaKnUEPCQB
4jX4S09keXa7KV9mDLpuMyYaGdNq2ETj440ZgwL8mkzYRdol8kMUo/QXCiox8W7S
Z/3XX3xXyJfv3o8+nPyulEsc0bGGmW6xfhsaIaWW9zAd/XdqeoW0+rDTSzuH10I7
C6fsJ/S4NC3z3uH/dbkHeXe4wDdXPOCsiT8EVtYGxlNWQH1UZ/Cb7Mlsij7QK0vq
AsW8BG8psCEuX/i6JD4oH/ssxqvB2dkxDG+MhLGd6ns2CsddRbP2BIpOvOVtaPOz
Qcbk5dxnM4rOsVs/mouqdGfJpGeyf9FuLdyiCfMP/lRCbX1dtCmv2IcjdaQWn+BC
5ruRlCASCIsPSlcu51PSLxc76vwhKC70WQZsyr7k4dLpygyJ1Gttwr3/Hc+CkTb4
ldYjzn/O8iXJW5UMJUruN+iJN4acblmXR4OBrrs2I7p4F9qL2em0I4DnDU+KmWsp
H9PuVsDiV36bC1bmj2ACPLwkIQ3gTDkfhF7lnLooMrS8tJCADuLQaPgIXZORhp93
GUom4BeiTtoc3a5X7TObSo/t2DTLp09ai/+91p/Pv1eFlZZrRU0SdaAEpx9lFIMz
QjZEfvV8ydMh3TwMp5ZzQ1fp37Ij5xjWXgEVF6m5pfGDE29M96tk9gnrmG6WhRgf
0h12sWHwk5jvYjxOJm5sxeI93AikJ7EjLPLXquzjOUuH8mYyKx5hCn3A7rQGJvcg
9KBeF1rKzdAagDyjKUlIw/YdSos/fIPscZ9cJGYASLAi79ndVpCcA4X743L4W0Cz
B8cBQU22KlGIakYq+Mx7IxsRbQ25Yt3NnbXqQ/fGzvdMMLIAMe8Wht4eNbESWH1t
4gkz4hvAFbkmAl004/LvRDkeGMaXzFO6eH3u37JRVI14bdV/vDs/mnCoLoGW9nuJ
injYP95qscpveOhnmWPm/BFA1fQMFcLQGsEX7hIdkg9RpyQP1FnHUuReEc3NaTsP
ao8q/iBW4vI/g29gf0Bebcuaj+Lg01TLdRZ1dz/L0Ovcd5qWbfLawGqZn62gCzHC
y1g/nssYN9PqX7GMdQreTKGSfgffh2wcVKCO5DsHO/cFRMUhLHwaoux9C/ZzZtgM
fbvlPG7jSrK5dM+s+jNMz2rw97vo5Tf/y58T4+gJMOL2Jo6zVk27Am6/efb0gJsu
aRxE2HDm//Jpq93PLC+yeVrzLJDcID7VbAwQW8LIwZx2lIARrSiMAZgV/PGUXZ4s
Val3K3Dab/Xo2MGeYWzxH/0tGHBqRqDvkOFEctVCv4LIc3lRPbS3LjAzXdMKCgeC
ScrZUaNrI3nK+1RtZhAUcRZN/g21VQLkJiPT3Wafuu/WNGjjuDOplzIo+7FIcLaT
746ztmLmciltWtPvYEMV35dTuJJdeb+Y+/kELO8bbC4Hcd3kibI+Qgow7s1DaAMX
0oA+c06QJms6WUCHH2GPvrxYGfv1WNqNPvSdvqYIihr9Sky1dNBNmjxddwNogaaN
Lml6hgvwXCwKbEZ/9jva2RFXrTlkjp4nAmdNDvrPcEyWLZuyM2+/y6HsmSwU56V7
YIX0GbWy53q3YsPB1J1yptaca1jDP+VsXydtLU5mHmhPVfMh+nBJ9I5PEyl3Vria
S2Vz/loy0E7h98bEWDteN0cAzuNlzaDaVTG1Olqqq1YKrIaJ5mPhGlZT3XGmb5gC
h+gTCRojqMXgrYyVgFbepaMt3oFrfap9IpqICZ+ZkY4pyjkARlpmoGubc+PZZ/X3
ZPGKJCiDOpbBSzpHqkNmnJpIopcyS/ZkP2/vHrhqVI9ky1EgEkxcOiQCm1X3iQzH
xLefHmjiYGmC8L+MB9Xie9OuPkmP/Co415T+putVST+E/tvQ/2zHumGpaYFWg1j/
Bl2MYK6HeX2bMoevtmxpKCT8tmaa2XZuxJ+QXzU3bjUXHPa5IXzoKOvWaDrOdvSg
kP9QIGslRz1uS6Eckom9ruMKMK0ikHg1YN1LYqQYMDN+j5sckcZ7Hl8wKDX6Rbm3
dYmOPATKWA2wl3bTAnsid3ZPcuVhmmcfro05gtLWKMOWIxtn4pbr6GzBTNHOp5kN
K+afKuDqwhLmX6o9rI76FJWMcLPo6PcQkhyWBEiCn4d7NSqU0+fQqVE684wwwFfy
eL+kL9TLT68Z3UrbuZ6gDjP9z+UcoGutF6cDburwnBium/reJsThur0TskOMX118
pEXW9bdFg/KNGAHrbfpp5kUS+dWRyRkjaLUH/fl7/MzURi/MAl3n51n82+KG0tBI
+1uDqscqtHwvrk8jMRWV1smVac+RP9pKDB/tj8qCeaA/0lZYyl6sebMmD3fkIu00
2w7XCMlWO/P5A7XGl1LgFVoozRQJlSF7C9mmmGOtXSMmK7WNPNj5OjgAVR9RJRix
NGwyVTBftnMHmkVE0SNdxij3wZFuapXtaN4Mgfk5vX/eMPppFUtlGWo0AVG5tdYy
BMewejWAlql7TFqQ3cRLX5bZkJG1BPAbMSzySPlYwurQzBKPKIZaspx5CifPHuAm
tUhTWiw64s6BYRCIqKAdfOXzkMP70U69aCaonX4PdEbnnJOH5Os85Vf5HsO0XukJ
zsExepkzwdnNAOJjNu5wS8YS9gsnYc9qmWukdeA1Zx7/lGwjx2Xuy9yNAaqachzP
KJ5rAwaVsrJFySoM2uL+73XO9c49LQT//B9+HZ4XCrGhlMh1FvM2LuCSKbVgAEnr
T86H07iHQ1GYxLGTrtP5SOTI+fMmAZFf22R94ZLzfo6L6JMUpRpVtl7iwH3biZM7
q1cLATofvADntQCit3jXFxulRgAU91GL+MXcDOE+EkHBvIXjyvt1AclmiqohVPIA
8afx+TkhYAG3IfuDYCEgyP+1lJ2db2qVZsjMKG5C4JVCRhOuJtrOPcTZ9rGg2DgB
nP3Y541jvSAPV3mb0rXhbnWeYt0d282GU3Of9UxcTpqCL7ncI0hyy0Hzu3bLMPUw
BSclvvWg55zWdaEkb1l/0RcR00jP8F1a2K7L5P9ygKF/YC5yzwzTn7Q9annhcOsX
x62GzoYc/Y83KmZZk54gX9GCZl9CpuQ0gQLIHPIfZyxR4R9OnjWnP6TkRWsuyn6u
covPJIuHmdl7f9XnqoBpkNY3D8JwOCiIDzASGJg13+eXfOs+clGgjFP/0sJkZVO4
O/HJ7e7ZhhL4t9NufzHmwHKKMevOpC6c+fEIlhgE5xwiVsWevclGSZ4gcEl8ZIg9
1Xw8aQeXl32f6wt0oU5tSTjOjLjnJh13z85A6CU+5YkOoJDsJ00W9YszmXu3gYKL
4nkx3aAUV7LTQTlnbxVYEsqPLc8tkr49G0cqRRItp1OjqibSsJ5dNP7fRvNPs6xq
9IPrsW95lY6/mOQ8N3DOkK3IFlMuMSb+L0Vs9Cx/tzWYXEgZmk+ZVA6r6DIUKBR8
lHfdKaGS1otUmjpxw9H0ZmzDL/8vaVio3m0Iz7AMfSdqLlYX4TTI70zrnxtKpKcZ
QuCTmuUXdjjIbeGyWSzgzcKA84viAnU6BI6Ijy8/EbHnFLcaCzdNF2bDKt4CdtZi
XKOn4wDY1f1qZzod9OxmclvS+1KmXGRTqfXxO+Bq/BVhHf0PnV2YRorZy9yGRUG9
JQk2zG8RlYXwKpHo1SB2MBDBQPeP3JoJETHhLk3KVEHAmXt+AITDZIuLswuqxnNb
bIrXdNNiZAjmF6g8TQLiPrld/HCdHjv1/CvNXk3LsxRlOmg6hW18n37aW42PMOmk
uWvfyf+8Imm69nQ8HrXGUtbSaORdKrqQUZqIyIwltt0suK4GGHuOLgz7CKnE6jlN
fRE8uwoUC6xUauEy4oH8vUBPjFrM3QcldcPqD3Mn1B5w7JVqLhbqlHRNr1ZesKwx
ZO3KZ326JEVxZv9TJMupMYlTA8fG+U2lDYjvnGrrIOo17nhlCUM/5JeVkTSfozxP
AQNzzLsPOeWkLQKcR2XfjkOrauqxufyzCnGg+PNutNj9CNnuIhA1JFN2WjPDq+KM
l2CU70BV319i6+loidq+/LlmAK7Rc08qYc+A+en0Dm4GSwOG4kX2YF5cPFCsI1xx
IuF1wMJeO+jttv2OQjV96EO8SEjF2NowRamQ5Byivpip6Ru0haQQV6+Lfh1OLYNs
BMtGU4aIuNhC7/jWmJmVAaiA8sexay34ln61XchvRFpanz3aqSZPdkYSEherbPYR
E6wRdNGFjJh9MBzpQMIQgI+HDL778gKscSUMYoejfW1RCszcNRDOchY06QN+zK8c
xlytCFptSWpQAoNW/rXcrrlj5rudrVHmOfA2FbWjlsUAxua/T9rxtqVALRaq1c55
tIl9Szq+FqR8n90bm5ECrW5nsTUMtx1UXaHrMuklre2ht51C60ekzf6M23shwkjH
Nq9hVM3LYknZjhvMXsn65Y8jFfRIP75qiZ1FqL8XmJIYHdvsLo9JT5c/vyNdV+t8
UfxeqUeT4QStSByo4xsovCc9foxc9NzxN5FZKAmZ/f2kB7e5FTBwBHzJEoh2Jj5Y
imMWDDCSNhui94HUiUr7o3TpHHkoz1YvDwAgtW/twn+omsJ2qC8mOxeAeA5nCFpm
9HZ2FuoC3sZ7SZTRjzBTlkfiV+7kPdrQVrN+M8z4THMjeHU6tlq4MWUaO2vB4iT9
Lxo4Yqar8hK9+XChUyvODZg180YKy8mP3mDw6qfhZ/LkubdT7NsH1/zNW7fgG+Pt
uUk4A1S0k2FO5Bs8BRsMwf9tqJPwBiPVEio6kwHHtHGl512bUqeBz7QttPMsQ8l2
WHRmqt2+VqFHbTr6z2wJ07NculjatIOLZYa91lBx3OrGFL97xM6+yycDLFzH0CKW
JG7Ke7eqe7Fnxc8JLRmlV9of43VyTVt6nw/1++0PToilHjFY4dw17njjgu8wJr5k
7I+BLo4fJAz/MxOj2samEO0P2MJY6lDLHRx7FjJ/2V3rzS6ljAtHcRtemDfSbz3W
ngg6UpepdvKGxlQ78W1nCXhsJ/2TvJ72Ipjnyh703DdLH4HoLOT+J9YUFLgIUBVn
1WAlr9HdvdSlxeq7raBqpFmB83xZ0g5R0MZTxhZGMaeRoBPWlV5DyxqlJ9jrkMny
fgNPedj5SCawTfbdFNhPY8dAcg5u6KVvCdBP6w2GyJp2b01ljXMLWtI6CL7v4aUV
DObLXWIY3PYbmkcRsQR6M9xl73uItZapgbg2ZBbUnoJRz6vxpfwiNOV7iIXZ3NY1
ZxvZnjvdRTrq5aHpVnT2O8d/J1JiZg07CIFrjNKck0v/K6zgenrI481YRwvehlDl
oy4LMog5CPJPZ6FuWwL7LpITN/zAUt6qR6uIM1DdIh2GC5x2ZKQcMqgKPjzF6ilv
eeBukvUwZLF/xJKp/Kv8xqtFPfMf1sucHq7geMScmLBJ+rGe6wGX3SNlwCbRLORv
S+9igDADCehw53kS1oScZOHV5rhP3LY4mv/yXlxoXZMg/VK6ftztOLAhNEVX+vo3
joWy7YQlj08p/THv9ZOwfNHlAUBKWZs7zXBCmS0lnTeTGvtWMeQa0bAEnEbMqg5k
XEjILAXSiehjpbRE4CvYK/krJLqE+c8hAeofM1JIlHjaP4m5WsrWURFdPQOYo7Fg
Um8GgL51U2MnaQGeyRLkJqNVjnLIBUDu3rCEtt/+dCaY1VHnsDkRuWl4gwf+F9I4
AsfPgIKohIjA++nfBq9Ipo3xCQzH6BsSy+Pa8AN70NKKMmUaS/Dwc9xLqvyd/ZkO
JQEVNgYG3kVgTRhOl7xsJfczhX4YJ6ULA0/xuZHiSAvLJBLXkr4YcpWWNic1WS35
e+SaVWHvSeIlwPJY5Poe+FCqGF/ZWfEY9RL/4z/nz1Jj9Tuz9mTbOZYddFDPN3pC
EJ4QPlsSv44B7zGkCqrJ+6DYSms/IdM/BAUICDbZETqfMqY7w+At4ktQhESy5OpI
7G08hJqPqXvq+ThTnnevgXxmZAAVJGcTy6UMPiTENso4GZECNc7eegisNa4hGbGe
tGvC/cjf+sYPsPv5uWYLAgxlOyGVWgunYVUIC0guFLc5RBtOmL9ppi1+F8RpCOBF
zYy1lMgIWk1OWx+CQO86HY5slEVafx8evznLcBMMvk9SzCz0jfCd2euyGG/XpFM0
+SYva5PEvaIzAWe7ZFtSHYdzN5jKExXyUhXxI2UCS6PBQktE5p0SaW1drrK4OazS
2r81JeEmjfm/4kHIHyy1A2k2btIX/tNLB1xjPHAwwiLGL/Fl2QFilpLOAWAzUVTU
XaBCZ7ybYnsntCY+/kpa4WfPDSI1f7PDHWL3+sZSW2QWl1NEBQlgfubMrgfw0qGN
N9/pkD2zH65ZVlQolktP8WAcWRhodiFJ6kQgDMPs9iF5IySI3LknB2jJIcQFL1Gv
kcBQ5VbOxfGuKU7NgFazJyIfmaB4wOnl87X5Wq+nTYuQBeruGolxqvHhJkxSMxpi
J7+INufIj0eBVsYAKpo8+mDC7WiAsbLcgVpImPLHwX2lkyvnbjv2x7pbCkBsge2F
CylngLzBBE9091XkEq/wS5HDOpAtsVHhFRTkvhRvDT/2Bt75px1aQLp9B5rzb0aS
tfS7S+lkMZ8t6M1ySZTLNYMyeSHiqr4vNdYARFgMWXzADrLqrBe1pf7vx2ycUJDs
OnoqUFgW1g9ETw3zYKnutpEPuwtEW2GzN0scA6YRfqVF6S5nndVkUmzrsFtl+T6B
wn7MEcgxcDps07PQFTte7R9exohXCbRSFOxoOCx/qgEjPGxgGH5JaHo6sZp6kOdX
PBrLa4NqN5wIVL6DMQ2GgU9nZM6y31/05/EtmCTh/xXRfCnFQFdj6IyDHh8f4NY4
EgyPyQEI/OXAltJ+2UfCRg936Bkz6sfB6ZvfkbHWCNHAIcBrYOcc6nNNaCUj8rEq
9PuHuZeA8ilx8rsyZAOA0WruBTd9AF//DJjKUxYle+YU8skyvGn0C540AHKQ9PJJ
9vHhyhR04xYvLCcuS4aPej/W7vSDb3T4trMbtBeX9pKFLDGOKmUg+1B5iyzRpb1s
xN/QAjSa1wJPDWcFj9+gmstFPVy0pMzDmz8Wz2ijS9u4UAJ6fj/IExl2S/9Wr+gR
GIznfMTZm8Bu1taeQ2irCreJmpO3ovxWg/flAchHoc9tV5VYWXoAy4FjAKeK/Tb5
QLempJLuRkxOsz0XP4CZvub/sjBDoIK7GeqILv2ajt3gs9pl885w+fKJ8fqpFN85
+VxkyArGYPn7zlYfIGYZrIdCjaeBxCz1ECi5PE3sJ8VQsPbHfP3TTObZT0+2D5kh
34/9358+6k0uvzIggtzkaLP+Lw5Q0yePsr7b6tYRRjpZhbZBI11e9kKenu6bs4d4
qEBJQ36SfV4vAwUpXg9Llza9D6Cu/o7CERmcgjUwmUkwZwulWdfZlsOejHKC1bAx
7cqMKYfELqLlYOfCxtLQ32i3LMfrqOivM7CnvIE6WDxbLpMzSXHopEY0nSj017nY
rC5UUYZ1jmqrEQpG292b9Bw08OBSr1e1b6GkJwvHRXxz6vAzx9muuXVx3F1T+MqQ
1LcyOtt+1rQZPAz69wUIFF5t5viULcYP/FJ096lvHRrFdnt29nfSlsCalaMdkbhQ
Fal2nYkxdqgawndQzAtpC+KdqcIKVo+0FViO/HBRzz8iNxFVYWcHNJhczHXTQbi+
sUlb66Epro6yr3fL093dPuTlkAwgHR9Qxvsg6EbWFNtfhM3Hvpq/SWmYY79aqhr4
Il695MAusQAK1+Ca+vNuj5OHvtispwyCdvkccK8EhVjahIFG5ri2S2AgIgedI+k+
Ozu7fbbfwgyiVC8JWNUfZ09Y+9ku4vpAt/Tp0sRxMCeBzZNpIz1Gh8ws8qZSurdq
OFstyph2k9/1nJBdxmtGc+fMZd6Mlb+8UZ8/7u7vYw9LJ1zQiUJhwM+L72OiTQ44
AbJvKSh7xoEU6XZqzOeVZYcOe2zWWaQY53HgVuiJBdWoDcEWejW7unjlUO0Uie1Z
moZasxhrm4tT/KYjf2eXebWenQDS6yFlpTzNLD/I4XwFzJyKpMNQuIq+nrMxvFxq
KYqzru0/OS06n5wRS6JStBsolYi6JG23axvMJ87tIzOG26cHnXCa243uTzZsqTpS
jhGyZMdWdizf1fcb1DnywcPoE1DcBWnRtBjRfddvmd1yEnbcEiY2JV8PKkupia7N
acQRYXsdZmjGeTXA3GrhT+dqRBKBin11s/Rq2rPWEjib7IQrUPONjc9DJTF0xW0X
9B//RDd984RNul0SFZgLH173HnNGDLvAnT1s6ohsdzi1FI3uvvj4fBfOtLdWVhl9
PaPOCl9V4SK23yqbFmvVz0SxI5TwtuvI+sp/uBwmwJ2LfRJLgCmKsmUrUYfOgCqJ
CK8G1fnto3hIil/+s/rpdkOfe8T4kNOUhwQJcyQ6z5qEzaMex1jvGbg8ZlAUNAWm
Deff6PbwPff9LcVfJOEltT0pkX5UtPEe3AyYThqx5TysQAFr77+q7sl4nXJ7sKfE
xJXDTR1Sf8ZJAP5VdeAG6VSXLm0bDvHedK+qlmo6EN20ktNMVQ1kDNZ1Cy3pgVLt
tbstfHiXDznqUJNz8Cq64XZja50kE7i2/dWdHyhuEOgInxbWblc+SfEvQgBoXdW5
1s5+i188KhB4XuDosPgYRppEKTzrR4NJIwp7ScZzBB0lI5J3RgEAYLLW4Qfx8gw/
T41QmLX8x1qQLycdhpNSed1Z2YMVpk895Vxd0KBJbGTIdbN9QATCF/b3Am7w/Ci8
HWxmKrxekr2L9yATTwBXLX5vrYBNZhDZgmmBiEvw5weobqTHu8K/uR/vcRsiH0Bf
DXLrj99gPV8a2EFcKkvEa2WVP0hPDjBra9RRooyEoOs3uz5LDc7sxxWg/oqtaHXg
lSg7xRZ9FrWJCh6Y5/bbjycDlmNYhnSKxjfGuTs7zsG7BGdokSTV2XMybQsPuof/
5M2aky0c9opcUNuDqVubZLxcwIk6HyTp4vqg0rS6+er/tpqVDQaaKbsWkg+KJ2HS
cCY3rUn3XjWaxHLDI6XaL7TIOwx+Vp/tppGkqjvbXvRM1dq/R5h5HR6A8tMQE21A
MALeYI1ooFNoDzw6KuEIP3Glhq0ersPVPFp4FErKrGoYBfkx2nkOrxSanKEz71l+
s9f4yg6RzG9/jI5e8Zz09zKaQuJYTn+Hc5Xw769SAzDIPjI1qE8rCAszBSUa2KBe
LZTRwRDpdQn60kqCgd0Fvgd73en3Tg43sbWtlxAeWflR0xV5srPqz1aAKgF0lUpp
bBEf9v/WtE2mG+t+WbUDdm4xwHNoMBsawkhD5njIVYhtgCVRComINeyNBlg9qJtw
MC8Mp0l8hOX4d243R4+Abl1lATZX7ITioullhJZOrmZTSscv5f9xDTB8qYoK16/3
vyfYBpYDTvLGNUw6cWR/0zmNQmxxU++9Jf8apMLXKGCB9Ueq6edRA0iTLSxDj0WX
utY+fd5+s1w/LpAYXhuhKh1+pTOUtJEBc9UEPqkCuAL1RF5HoMxPb7WAJ1WbjFyd
3iumH6tkPdfQgbKZWtCkYg4koIrvC7iJHKVFAuV2Kixuge5XRap/NbDLywDGEn2j
4XvDxht70dcCAwNFD5/Urv3gQnC8Q/JZG3m44Br/e5LPPuNnepGCHq6wiqe2qDrg
YUfepLi5uVXVNW3EEq5FpXal9SSUsf6APegxi12QvHrmeUjs8/IQku1n+RWQvtEv
Ahs4evmrpf6XeUkct0pQEU3AZsUgEbVBCSyde4JgRx2+vNLJOJTHeb1YvV/MS0SC
Bs88J1U+PBLGOSWM2+V/uRI4wtheoXp/IalNcNBlP0GPDkpNYiudyBJRF4u2c1up
M4KW/CUU25BpstVJ0YFBtkgJiuQ5sf6l91lCPDImuAR6wd7WBk5IPuqssOvJjMcP
5eUDnlSNeHlnqL1qC/C5O6YZ1xkqPeMe49edMAJTOIVrcXC4d1ybDDCsYgNLlasb
RXUJWhMNwuu1iX9AUa5xOI7ZH8nnhXdqb9y+XiYLHdnsn+mfjI1a0PdllOlRNcsS
oWhwhFEa8RwM4RfjpuCOSGDMN0yeSiim8dr8nL3yG6BX30KTlrnqwG4AGaG62JuG
Cq+CA3Z+Uo4G+BUtXsR+rKTR0vObFQrM9OBg546UrHPgqQAi4xuXMmm/dNlEOoXF
VfCOQSQ0X9qv5nzTC/RaCYhiefL4Y3rQvSRIv4w4fxadSzmZ7WVLBBAJq5Jk8eBs
n56EW9cyzWnzcwhQ29r7jWtjB7vrncnYnQuYp35jlNeV5Qyviu5Yt0nVIxhBU6z5
E441Kra0ennEslDCO1gqB0vyw+m7PtwU6B+npcNvnsBdXq3V5MQsS1c1yFJYQDWt
87H4o6+qQPP1hC0BTUKU7vP3ezjPf5d1Xydg6nWVCBCn7BIFm+fD/jALdycG3jUw
/N9mCTKCT6JZzwTDioiWJn8DuhQK2gIVB3cgEDLbcgA43yPVsbAxkWVa1IDPX6XI
LjdL8WxdT0isxDVtKuEBbwjabsO8ddRXAfH0DTl67l914OH8AHbfl05ud9UiLel8
3uplpo6X3H1I+FwIZ56r0PEJ8lNr4Kowv5IR5tbl/alG04ssl1x9wwv3GCt6gZGI
GYjWmtrI5nMmeNYPfXVYhmuIjDHUOW4TNKicUFRCjD1gQ1auSaFcCm11H4CCBlGK
OT8DceXO+q3KLv63lHOKwFheNybcaEg6iti4Hg5QeNoNM2Mjy/uiS7IgvHjH/Zko
k7/GOPynyqrpxX4ICpMusWdml7Xht26x7CU4skeuWqUo2R+UxTPI1R//Et9cd3Am
dwk1XfsvN6oJ7GpNpOc9c4CFYGclZCK0b1Mnn0aZ9U6ACL8ml2HTPQ54jT+rzUEu
rCkamfAqtk0mfpiPHr3XzOi+stsmCsweGjUY5gjp8evgLnSsy3uB2kBK4IScNMWT
QSWAbvi9vCd2gMG1kbTmd1FfAiivrGpGRyU+Sasj/SAPEcxRDJXeBzPGI7L59OCx
RrvYW00wOr/C5TQpQM2OYU4kTeJ6QC1HeLLrJ3GvL4By/ioL3vXQODL2VO2nDjHe
scLUys2IHGx6e9DptYTyaleKAxH418khH+LCLajP12Dijk4s+0cJsNTXlaLRjj2E
dydxt9MxWMK3YIUoec7wynQ0SOFlSasDsS73FIt1b5PTP+k6jDtuEA9qm7p6TmuF
parLEYaP7GoRBF4T738vrz76wzhFyDVBBc8LiHXxKB3Jw1c2hL6hhPL20nUobk0h
N4LI76nbmKpkUBkvcgTes4SgiGYdIR7MIVQXImsBVwL8GOoqFIGkDpYaMaEZ27xq
N3ExnSfoiLHXfh2mci2l2kZd7xs7iuHFYH5UvRheNUyVkvpYdwkMSREjivDIBO+A
I8N4UnqIyq/TN3eW5CevVAqUUwMAITQmfYCEYSqojtSy1RRetBo2RKROCKMFIm+0
/kL2AscWmFMrrrRNWJp+XZ7WQRqnb8JEvXfpjci3EcKPoVAj/wYDJHXICRS1C+0y
lxFlMVbFZSCVyO8qEQSXtexB792vrylAXWayYIfaT9KmDzDIpBXhnAchRYoXtLIx
eyY0erk+qw1+105K3RkAuSoY0dyyysIoRNDUCs2M+dl/LY1eKPCTUjIo7X8662Kr
0iet6N0kdZMIFZxRRr/nvz5gguZs/+Nk2JdblCsB4PqLyj2uXcKwoa5vVoufpeLt
T3sbG5PWgHY5xwFiism5vW5nfnmL6aOHCyOXt9HsZdeOq0QPBCZrJ0Rteil02D9C
NTGXmOB1dTK6CzSllLanmnN9+p5mdp9hZL8ix+imaVgyjyHc74oqk9bpAyVLik2a
wJBzHVBRSOqEQprjTmBDr05fyacy33JZO1d0q0fpyVkQseQtnt5SAU/EB3y2wiaz
JgUS0s6fUKkv3fQ1XYF9HwH95Dd3pXKTusGdZTYJ6wZJlBQpnFSfQPP+qR7c3Gal
pXLfTbVD8P7Dxr/lfV/OXW/Q1XLUoMhisqbzUh8tuEsr+65ctZ05rJk7ludOveS/
329mIEjWDu1mfnuQWvli+9/7edMUlQT3P4DJUdIcqHr/bjXUUYHjXu5DsHCsdda3
iWqbHdajzkyGANa3JZJxg+mleWnMNOKlXAqCR4oFODItf6TwVl09suuqiM5rLboo
ZxqllDhyOs/AiDHqSaylIYckviKERIi+iwfHa4ltj0Oe5SrLb8qkqdtJN3j+ptkQ
EFkaZUxVbZrfzkzP+4UfiOnq3rlMjm8iSo8kPxg7rFIQJ2w5T0uDLWzEHz+SLSht
Alh9CaFyQk5bK+Ie4qAqLle/rMSF8paD31nY2ba7LERhNke7Ee5yQF0ZyC16BOQq
UZS2Lb+JazfJQttF1pFlsvGFL84Y1yoEk5WR8y12O082CdoKbqKriJwJkXtQ5//b
udKlb0aQzx9Qv++96mfgt+2+jU24lsH6x2Vcd7h2kwhfcvGvKUf6O0vNxMWT9t2V
1eqQEZYjEDceu1PTlKtlgj0KyHt++5k0nezWoGRI6BY3SO7b42fuDkGe/7F0rrAc
NeRaPktNua957Lm7RtvhiKLxFpKlRjd5rK6ec/Oim2VN0NFkK65saTWr6UFuUeYo
32dxqGGMlU+3qrx8QYlGj6OwCdInG0ZMUdUiGwhTwKOUINzJXPmI0QnARpvrCqxH
+lQLvuIs8KbaixX5L+G+wudRukchVaYSLuYpQfb5dJJTqn7T1HqlO+pK7EJOOjv6
jh1r8a68TXVRiCXNL13/PYr2j0+i+5IoMChD1vWATanjcl1SYJNuekjIp87pLMVL
0vsdbU1jdZVe5Y6UNk0CTCC73Ch8xpMmGJ0/oE0rzQUNG0rHOv2D26r5kGSaHAxm
6eAk/pRSR3WMNFJmXokh2HG4jzpYrP4j6IAHYtCMOlPSeECm3P/tKh7S8bA4n8xO
arI6WbRKkPAHC15I60WvTaOddYwJocqKTSaEtGqtICprD5jfIn0Irwa5+yTc9rOj
4ATAm2zze9s8h3u0NAJsYq0H2sVVKd8U82TYeUhTCoyy0M6gDxr/BF0p/Av33QEY
Jgt14x8XLn1orAFmElRDH3l7GO2EwQ/nmyyRMEyBNmawcA41Odp7jtFwOqH4W/Ue
iHgLgrL+z+VI394EQLdVsOzDO6xNLZWga5XfsFKfGOoe0nHH3XlJIADWq+6gahO6
ZVOopHbMJDyfgj87FhzWzwl3Sj6ktDqP7QcjU9RCaY6bNnbMCEHDFReC6M5adSBC
ua9ZUb/MF7noP33JE+zyVlM+9on6CjCXkq27SagAN1wRJP8rWQ0SMH8XL+TdI9b/
wxsvN4gbkeuFobrBhDcf0eU+3HVIdctx4CAXkH+SpRVFOrXBo13I8sP5XL9wsH3L
Ss33FIYdoR3ZEPJhBtQISMBuEGsGRvvEt75e7urc8LMgEOFsuLJbt06ArZYFinOj
rsKAYDS5bmN035IjoHAQA3okB/BU+B342CO+Atcr2S6aMkTW2697ULs9kAhwY5Wi
EUrzWpZjFsTmgzXz8iWWZEGwySNsV6XW0QoqGfVGTH83wMZpm/dqPbDvunJQfAnX
aK8wy1jXtlPDC68pqL9PG3ftN1CZFkPLLZRdbVE7F7EoDv5DgdcRu8K3rudisL2e
xoI4BZ/d1HPHbvXUExL9t0LYGIufG6NDjyvrqhAbqlzvRk0+d9TYVfXBsqoQmIB8
6j750CgOWAqRwqPSSxUkZplFKRBLsyKV8q6XvbUn42XK35+dn4AesTlIxeApgwVU
S+Cb5dk2rpKokCHy86kuE64oL14KxsMVHSQFXC7oH0lOvd6iOpRgztQud2thMpg5
N3O5Lj/7X7KCJbertzm9IjyYV69POz9+DzEwcIgxt/nO9HE8+HcIYj2ND0WYwry7
hrNNn0rbbw5x502Lhp9wE/3Z8FN4Wr2zpTYQ5rZWebX1YEIJ7+Qs/7ef6kFB7qJ9
IAvUnbL8g7SwCf0vRURty3FZacSGvsMpwZv14mQhnnjG/JMHSU4mTkWZZ8GS09pr
Oh8ZQ6ocoQzwot+JaiBL/YS71Nj45kVW9avjb5nXwqNubjQl0zBtj+MolzeC1Sks
R9RWfgrbeaR6FjQD58R4uaSRRybXxMn1SObQr384of76kM7BGInZGwjd+q2TY1rU
WfDG7hr3EuBxT7c4eMlaPTM9LkRhF2rn6HOMla29It9uyVpap9OzIOVpE9g6flhI
DCbJ1y248i+0qZ8FPFUqyBf2grlk4/NNOZt8ipJfQuY6/utVdrSLUvPQU7byrvg6
K/HtnIh/VORGaFrY9t8RAatuOvaxz4XtG0Lz9Fj3dMHiumMEK8Pg3c8phqD/0wBV
wa3eqyN/bjhh4yUxaOHOcPrJyjYzf8fDvtZmJHDI5r0CYR1ECMJhcEJnr9dsRw89
9NJMBKG7fOwm8u2Smkm1GRXd5GPUOxfOElYRprg4FDRhrz1Y6qUhe7IdjROgSEpf
Gq/99tUkCOEgA8nI0hDnjak2lkKozF0KxSqQNv626CpG6hfIcuY7aP8nws//rVSP
gY4KrK2pnbBNhkGAhJriR2grYXEe4hqm4cJk4qJ5etywMrJFr4O7cBlYgpKM6GeE
MislCY8OgHl59elve3wBoD3NPAAfyjtPzZdOZv7gqtlq4JDkh2ZW4wqu6xED4E3K
hcEYaH7d4phF4cDHajL3PmNuHLtSyASn35C/OEso+HM/pxIx0GJ08VQNCrrH8C0C
TEF3D2XiSC8RMhrFopn79iP5h5NLFoHPSkcHlVSDvjzvWczoJVUTyXSXIgFJRmh+
8I4lXPqbHjyj7O68oBSnYSgwSDns/df0v2fEOJS48egoZskWn8NdfnbYV3/yYvKm
j63bP1TferKRCBPMXXOtc7XJAGQUogPAeuLvpi3et5E0T5qnFq3qXpkA7RBh1FPt
xuUJuZL8IYCeu4Vk3EwEAa6GRfrzIdJIIj0DBMuq/m/WGQ2WkmrJa5fLF/10SbNa
+4BK6Jg4wprNLqPTr/bld0sdR/gEdziG3yOMCIpIIWCUSngPpHrW6nr/uvlGg1I/
5199mrAIOuHREc41kZXbRu5JFJnEeeUhaDnkkRq9keryKkqQLxvyEOKyTTzvjXQP
y/a4UPYIIfP8uKFCa1ivK09mA/M/XEk4KkowJs/AqWmOtrTnwoa9X++oPzcdFIuj
rNykSSkFcKzrcw4CEuFOaauL0CoHzW1jjbTEAHNk6eZBzQPzeMDLi9LLo6jEJnBN
7rPKP8V/IFoZP/ehTdAVu85Fd1orJsX4qtTDWiGh1D1hAaP+lpZTGG2OnW3B3e9K
rMsZr+p3WzPpc6cATuOxBDvVbwi2wMNiwMAtumkDNhPEw0+9kmrTnZT7qK0z3nAB
dL8MzQa2Ngf7pBfCYP8cyHJDsRfGdou9Z7Q1/N1kG9dsispsONKzOp8WbG7cKL36
567j+WwhYYHPIFzCE3V5zgxZmGVaFDxtvXedqs+X8+5MMTkYUPTtWmtPpypokpRq
jDid1efUiebYLWakOKTgRhE8Q34sZe9Kb9amrByMDUvMfiN+mzZYJVU5Io4p1N80
gyS0oc9zZ5wk7zvP36HCcqZloFFZD298xEniX60t31L3kfWcvS0FtPFlyc9VaTxl
EGTUqC0i4Tn+kcSMQZbnlvBEv66AWLLU/JJr1+DE7RTgdvOzpWwz3Ed5ZQ8mMf/y
xE+WWf15sKySi3LOnK9mc1bFf7h+ywSpBDXEZfram79DRcXcBleSWt8He4FvIrtV
7Sksgt/+bied0rGjb9pp4Pm/K2rZQn2jAu8BUeigUho9KM1ckuc7+N3dR1TV/JTB
NivVmsyaQ1vTI+qTnlnJq1szKzOGJ82QJ6IhvNkMyIjvjNpxdl+wvyxoXxVOFBBW
gpd36NZ1Kc9kFmlDEN3yd6rQsdEiZCNI1IMyNhn7//HYy1zkdvdgGrLX8bgm6dXs
L/BqCD3oO8howYQBjfVe5rK8/fMGHGIq+I1Megamr7DkMlEuyEu7d67/SNpX+jO2
Y/umXR1Ae/b9lEmm+wQoCYLVBLK4q0mvaXld4nM02SB3RkCzXxgPsVsgJjR4KxpI
bQbR45qNQ77d2AnDqK7v3LUfgOgtjw+XGdy7rd0EHXU8u1HBH37vNy/It6sJVEww
+FTy/vunzLA9GWU6NbIFv0lWfS8OVsqUJGVqnbVnuvDUPyjjf+s1SYbTrXEjUv7G
IBEtkOPYcB6uRcTKwgd81B3UMZeQaZNO/SvXR+1Q/tIDkZUlwSXXKCN/bAGEy/en
Z59SlXM6NkuNXKTZ9IwtW/RpVhtaltANqOEA7gNcZHvlQkXqivZ5y6R8qnmazNyy
n/FfW3OXHmD5qwE4SqP3nd5MtX/ANt34n2PbgRUqcaI63VmuO9y4aLHsWhL15r4z
k/ed30C3WevRx4n1oxgrWCeGdlCau8tkPwa7lvSOTC415079HxEbfzcQWvnryepL
L95ZTGC9yC/5+pyNGsPaIjHdbFzuYGXir/Nyu85n96hvautBCL9YaUnbmpZQN5mz
gBSeCjL/rGdBMnD0kOOp/4SFO63KM7sLBGsU4aRlVmw8zUQc4uwvqnpN5PJpUu/o
sq3M1JdBnwpv1BCYTwwqxWT6oe0uEUWbqNZRJxgdZfwm34qbwgwAgRNYR+xstbTs
AUQzvH1Kt/UbO+6VBjOm4/JljeASd6pXphFyg9oefOmfXQxYdo+Od+Lae3m6yHRj
RZmavA5qYfZtUw0wSxowwLPn9eTAnhXVtwoOS6/Wa+HV06NNiXELbgULYJezsS7H
IpGoOyZyTi35EZegSc3sH0+xXbMfyixhGVH2nEHP+pctpEMaHxfWM16BLFneWAfF
XU7RzaFcGeF0xnw1wn5696q4JJa9PalPuLEHLTKLoJziLPtsBpVgNziS0zfecUwH
pD1jpb41CFf0B2hfMtmTBh2Y5Kko78uKTbeCWdek+N7EKtB1KiEXLJGbfnrAdqCV
4V1FSwqWIXMYxEyTZ8LIS2FFGtb+6EIU5ZR7WrMoPCZBR4dLNFUJ9mhU6g49DhQo
XzRx0xhRGfKhGsvmHwxqM9qGprwesKPpJOUYIDboVn3gRPP2ECXtKwKwgu1tZFGY
blQjoBb5JHrYTS+La1dBP4/zca3koPn2AeWqYGYDhuEoRC8gOFenQQ8Z1yYFfVgQ
mIv27Y+sodwFV+y9Em8oor10wm0hO+nTU/DCVcmMi76k6l/CN8P/u1nUo5anNOzn
VoM7UPkj4HvUwivuglEgQGIq7kGB234p/LtvsC0xA7Ic74Ut0EmNpbnsaa6kLPH1
bgjN1A9O2WxPagihMJcj+u9aMdyLjebmjik4umcT1ZMoyZmUIMbAAeBRzqSwGMBF
ackNs+AnYlMzQ+1w45s2OVsGcTLVp2wXfSW4xFCVOH5L2wLLC1tiTNkSZzA8T6Q+
Agwy7vDzVjtTdabIlctT550O84tC0v0dB0iGzV3guzOB/N3XdtuKoJKjaAXLFc/4
Zv2rKLioNN8JMcqZYDIcUxujgFQD9gkE5DOvqatPTBFTT+jgvoFib9mzWop/xJeq
9X8IDEs6+VbwT2bgv/t/WbjaZutIrfxyjJMjGYEGiTq1xnrulmpV1dAkcIuVEXMC
6ws2yIXhSYhI+Mw7azVkqP3uGZPpBG2zeKatAgUEhgrG1VUJT3ZJEARp43dNENnu
t8obFeT7KwiL6LLUtlqqbLOJj6AROthGE9EsIrOG/gMsj6ODPsLfmW2IjL8uUDns
1wePj5pYvlIb9wz9csPk2ZAWEz4dysFgVWdddDrekSJnwMluD6UhcKYgyaJM/k0/
jtETXHzr6PukXPmPajrhgQIh+4gegrxGqwqIm0MScmN2+Vkr3Ydho1yYLaCvo6v4
JDC1edawl41gTAL4eQaSbYul/jQWKPquNMUau/fMt8XzmcIwRdzXeBSSdUrEr6xA
QiAZOTSzgwa63nWPVVnSr/nVaWLQkdO0bZM8bWcdGzDOtRrYNuxWDzOR4b+2iyuK
ktvY+tl+5PvRP0Z8MJQTT4IEYYXIdzzLfMN7Xscx1gzIxWxqSyZgWWKZQUl0Gpri
jRk2varcrD+ENc4uF72aQ/cZkGiiqUcmD6moX6gszSQRNJBbDkRYZ4e3zGDKWAzu
i+LWxW7YEVXfxzZGh0DP/5JdcvYgUlXFH1nDZ/a+/vD42pq4BiXpMWHdY4dMU0Rs
je5DFmY7cx3iwV5KOQYOS3hHf8n0PhAwTnHLLl/sJE8x+OAMIDVTm53JBwv0VVau
dtOVYARa4gtL3T9S4ikqkLw76Sk6+aYYjI+bDXGqtFCfOwse8W4BmZLi1MG9c2SO
jQgOOINyJWf/QNhxhW5Dfu2wnhlpbVzLhCerCvnQ2xms7dcMQyaSOuX6gQkwKN4Z
7AvIh2JN4oVAyKhzsyLGicGZOTYZrJzZfeCaZkBmqOiaJWHaCpGv3TpLs5JHNdcj
NX1XJseMRZk9xrPjE1Hqn14sfgtvnUg/v3RHSb+3bT62KfGPDljF3wBJYcdo6nhc
Dvzi1yuYp+LE0pn7RXzCFlFIka/PHk8gQsbgCX8SYchWRyFyHPRyCeoSUaeOTpaD
/ZR5LO2F3ZEClm83/f4LH3IGZzdcUKgt1CP0F+FpOimdFYp6dwKGzHOWWyTx3/mW
d2Onq2H8zBquPMc3WW0JqDX7lAwkO75UsNsBRsFkPar+DVNmhWLoZE6xIkqdLp6G
9Kn7gvd9inPI3KIEaj0+Q2zL9iN0Ud71P21yaOt44C6wkAtNCWmP8iknf0aPng54
LAuY4aWeBUGULwQG8VwOyWnWjtHQ3dxlzAmF3GgmpIkHC+9djOWHaB6yHGqkbZbv
e2kulO3hTiWMfezXMaaR9L+QCgDZuZh8sHyR8KJYBuSkK8E07U2b1BO7hSOn7kQl
atikSazGeHSbzZnT7+3rgdYuN3cx2LsTM0R84FCWySr6inYPjSfZZBE4Xiv2/OHp
8hIv9c14MYEq/xsKr2YaGejsLLL3WscF+kZRkd34TXi8vTnM1p/7lb+QfP23qBUF
gitau2CRkniIk0bueom7tum6eoyaovWAxxl+Tz1VMn+seTcX7+cW8ieq0xLc9Rqk
hWHRARlHsVfMQFJMHfKlq+4xErO2yCcYdt6oaTMBNCqatWqkFH4Jd0j5TjrP8OYl
yo2hV62olY6HerrYKz+FtIYMRv6kT/Z+39EkwXuKJguuECMqedjFLtFuukBY+Cbr
EmxfYKg+bAcQgQu7+fo+pyQn0lHptME9JhZcwx8fMDHwLnO6NKN4tn2zwKL4jaAI
gz+3IbXmt3VgGi8UXwA1gVbuVNVfWPRkkGM2KBeqTxhP0grmonRhSSjOG06UjsPq
UDzYktUkXR6KFxefGhhPilmp7hZqOeMACOa6cKqH/7prSHTG/ifvbWXBAnSf+FVq
r6mXFmromHQ2PzAWrbFfpkDfv+YLt6Fh76iAerD2zkTgDw7JVezjL/I1YkrNZJp5
NyO+8qFK9ShxtErZQ7a0LAWoLEdB/03C2tLCwl4atuqBQ6BR5f3B3rulLiN5o/XZ
2QXKCZBg8kyPY+r4VbC1gsWgt5FHeldjwt4h1pLbY0VW0MGAcxTInXGS9al0yVyp
zycY1QHCLDiacgOWMcDeoXLjbRC/TL6ABr/h6Y5zCyy6+uuMvUIS0vtJFDTVoeSc
kTFYPBYF5KGzIvkzbuHnKpLU8MhGQpgsUhXFAY618dz2cwxwEvD2S4GWjf3BN5sy
szYedMgDIP+XZW1Q+XqqX9vvy8KePRwSBRNeZs3siBnPRgJD27jaTaNnhg6mDe2z
bdvGI6UC+vtwRlgiXlUKKjXjab5jS4nF5cMSMxVV8RuynI4nO0HSfi66Bah5TGhT
UIz5X+9ycsN0sWvH+OWDYP8QlrUyGUfeOZIsxM70fUDsLOcziWASnr44QFGeGHo5
wRp2ZJB9cpV8+NINDVPPu3wNRhdKmrsKiQEmmHStWqY6AXIO1jgfWR7YEdcQnQOv
8wuMefvNSxympq3fQKTqA0o2B9OUX8vVzLbhvnVPLFSH2Y5J3AZn79zhyZWASb+z
24T4CDul6fyDVeKMTRV+BjuNPPNZ0OVlz1o7305WVxd+OA8Q8cDbKs5VTJh4hG8o
AM/51yQ5FLqVtwvu6nGBsWrdHBc6hH0cX5M8bf3SANbU3kUZd/ek+rrg9TYwAs3P
WPUbO5YfhnZlNB1Zt2S1xCLrwUix4bWVxLS0sTYux8qbXEJcKFf5hVVXvhiSWgox
j9/o6grSxgiXV1aer2nmzBST4eesnGP24lq3Y4I7cRPOBGmXAvaJnaXz8IFrZeSc
VEMfoEf4ZmYwd2DFw3xVKr2A1eqJmdpFXamGFGSlERO3fRB3oD/Y8/gXlvFWkVbd
WPKF3b6iTtQKY7Ij1xZHpBGzC7GDrpB0PmrnJlF3yl3eyF1W29OGJoYVNHeDCyxc
0ICt3ysZox2X/dPJML3AvmCrdflUmkHKvcCuGYKgvKayD8dKvBxS9ljWFBfwPuZq
uRwGgfjd8tx2yL6r51pGhY/RnXDhgipbHTi7w4Goyy2StjU+u2orLHHxrSkUfILJ
qFYE3NIHGkiDAzRUZZkYHRMNJ8vei92jhbbkxE71/zUh5Tqq5UdlBFcBp8YU9bFY
UzR8kAFs9fzjrhAJ0LGnbHnYPpLC2840RktrvDO651i8G1Pfn6jCi28wR/BEVBj8
MA2IYoH3QWsith/eYJIKN9YWnaUuVxOA64Go1iy1CVfrrQ2tkOvHw5LgN9U1bT3J
/cEFcmvRxz6rs5ksILX06jN9cKLeYSV07fuIvEJMGq1y4qgqFD2+8yP7QS145B5B
wiQu61SKJuado3ML4M/VJGpgcxClPb5VQLDGGEWTVzRUatSaPMqDhCkzOMB6s8ZE
HBDJdUta0VVPCIP23PM+n2D5ONnbiFz5CVvtvzyZMeOAmDBcFFtuZfIF4p69ybmh
egCnjYk7Ob8BfFoOF3MNX3Bu+qKRJeSfzoZmtXbugmt9NdRe4LtqkhUE51QNI2j8
K/2SnTzoVKOxcD4nQ2BrpJxqTCGcvQTuT9DmAHkfexOntvPDmrUEL3YP+Qw3s2JR
U+ehz2/LVejeP6dc4bdvMoMPjb/b+I0ewuInmZUJ+bMtw/eDnYdx41qsRLknm7zR
HSgftjyjc3O5ygA86OdQdaTSekiTnbU1japdbQOQjCKDvqnGGLwi5xFkX4Qjj5HY
HwckANzwbLZEICQg9zLGk0NKAXs5sdcdJx2Bc3UzGbdAH9dsxkwlgQwxbE34XS3O
bAHwLODVjIMXQrO0o9teCpMb7Cfz69ib+9tGiQFERnq5+gZIafPuQQxTm+SJw+ey
M+VFMk3gIynC4qV1fOgxTLv7ueVv4Tn5AI4y/O4psARrfcRL8eHhaDfwOXbW09BP
sYfQrXFWj3RO6OP8RrLIx2HmfKWtd8SWS1tHyyCkh0bXepe47NU6eLrE4FVT8n8Q
Rey+SrwybQeHnWOvLCss3U/6Uolg6qwrp5GQM02yILydKRGTjSjr0n9Y12YldoB3
l1x4GIwOtDwgrDpzIBolZLxhzbhlIpofewwlBEz3a17txNBG/w6APtt+teLdNERu
eOD+lN5X9Ce7tU+bzrBVwXXj/21x47BT5cQ2ABzIQrLckhvz2ZNpIZ+5UJz3r8un
4UM/gBtBcWZK9Xoag6LzhYn5/r//QcQzoU9H347dUuH4HMOmajM4Xhsz+oEVHVoi
SfB6xtWMswYn70gOOaK+ZbArsAiW+3hQyIVcHibn5ee1tKc38I4ZNTLbVKqe8Gt/
jf8vf0qm0xjcWelInJ+vMG8AFd0u6hbdjowedWnCHBfQy7PImPZoISBk0JjdzFIg
tlvF7cMk0xO6juf7jv0FqNH5pc4W1HhhkTr4uTZ532j4iotSoQUi2Co7SU2PhHu4
jV1ztcKFX4C9XGLc2okFgi7xsuAmJGfS+J5EvoSBCyR7fxR3N5HyaiKlgLU4hoOR
TwwAT02xywoQbdKpjtAm4ix/VztiQW7UgehhrV+3lN1OWhhtyGR4a0Od/wvCubEO
IC+miGgpKt1I7632dR3H3HLSB/eC/jM0jqmkPYTaXBsvQDlPy6ugOycGcKpKfUvl
enHodGpouhUSmlYUcoZqcothDo7n6ynjR7XYgw+LNjv3CXbNaj8xMdb80RA/+n5T
8KcgyKyERmWcoTuxa3DCvECJqBnWMn32fEZyidcxP/duNyCEigdmnvZWWOQfJn7v
XZjyUU2SFkyVyMRPUVj3HjDpJ2jS8TTVVESGcnEwqP1wNCn4f/N+3kGX+kOp2EMG
2wF8PipA99W9Qy+5XGKUBjpXmDTegi4JD9O6kE4l5gFDRyCW/kAP1+aoSyUFM3oJ
W2YNrCUc6mAFwlkQbrxeGbh5f8CBlbxtkoVw8/QEoaO6m3WIq7MPjKBjUzRtDkpM
g3ZH68zzNxfNndGK2mKIJvVMxVo/blGqKmI6ZRUE2zfuCQtdKpH033QiyHfUMztE
UvHLPqYlZzVzsIRRKIuwhpYz54U3D0GZ8QmgO+pWAGFsPfO2Aq9ctyrXQJB0/p3q
TYG1MHsQkrrr3QtgffrOJlj0PwfowbW0kW+OG0J17NWj2XJQ98fAu3ZVHQW6Dmhd
JYO3BXHVvBoG4g9bhxekOF35QlBVqPibbSTztqdr5onYs5SUFeJdyOnZ85fKI467
/z02kmC/fJ15uhNP9lXBdVB36rB2IPydeQ8YEhHKuAN/y46m78FsZFboaCaqj0MB
kl7UgeYGPjKpxEfRzsS3SWJYStJHg+zZAGzyA2T5fL36L44H0HcUB84G08P0RAEe
ufAHu1S3fDESivr2Krhy554KggXl17bnbrEaLksMdJxMywmVvoowvC/xmYWB77bP
i6zi1XfDcge1wKNtj5UEaF6Hw8gapYTjM72NFZxL2c86X4vgnPoy8iftcUSOu0JC
dohJMUQVtb0lZQo1s+LldAZ6BbtR6mfL18NKT++GEKjmO9yJsAqpPXU2/CrW2Hz2
w/Z/JAkmLOxvPFQH6SwamRMN1sMLUPWUPwm4gdxx1Jje9Hxn8axjeTCNY5+Hn5nl
5UMb4BXiRwsbRu7iKIQ0IQ==
`protect end_protected