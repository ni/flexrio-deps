-------------------------------------------------------------------------------
--
-- File: PcieUspG3x8TandemGtyInchwormWrapper.vhd
-- Author: Hector Rubio
-- Original Project: NI Cores NiDmaIp
-- Date: 14 Jan 2019
--
-------------------------------------------------------------------------------
-- (c) 2019 Copyright National Instruments Corporation
-- All Rights Reserved
-- National Instruments Internal Information
-------------------------------------------------------------------------------
--
-- Purpose:
--
--  Wrapper to instantiate the pre-synthesized InchWORM netlist.
--
-------------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library work;
  use work.PkgNiUtilities.all;
  use work.PkgBaRegPort.all;  --Fixed Logic RegPort
  use work.PkgNiDma.all;                   --DmaPort
  use work.PkgDmaPortRecordFlattening.all; --Flattening and unflattening
  use work.PkgSwitchedChinch.all;
  use work.PkgLinkStorageRam.all;
  use work.PkgInchwormWrapper.all;

--synopsys translate_off
--For synthesis, netlist comes from an edf and there is no external library
--For simulation, netlist comes from external library
library PcieUspG3x8TandemGtyInchwormLib;
--synopsys translate_on

entity PcieUspG3x8TandemGtyInchwormWrapper is
  generic (
    --Rev ID is used internally to indicate that this PCIe device will be
    -- reconfigured on a live system (aka Dynamic PCIe Reconfiguration or DPR)
    -- 0x01 means DPR will be used (e.g. LVFPGA target).
    -- 0X00 means DPR won't be used (e.g. fixed internal FPGA bitfile)
    kCfgRevId        : std_logic_vector(7 downto 0)  := X"01";
    kCfgSubsysVendId : std_logic_vector(15 downto 0) := X"1093";
    kCfgSubsysId     : std_logic_vector(15 downto 0) := X"C4C4";
    -- By default, the Inchworm will only implement Chunky Link storage memories for those
    -- Dma Channels that actually need it. That would be all Input/Output DMA channels and
    -- P2P Writers used by LVFPGA. This information is obtained from
    -- PkgCommIntConfiguration, which is auto-generated by LVFPGA.
    --
    -- However, a given client may implement stream circuits (e.g. DmaOutput in fixed
    -- logic) that require Chunky Link storage memory. PkgComIntConfiguration would not
    -- know about those. If you have any channels for which you wish to force-enable
    -- Chunky Link storage, set kForceChannelEnable(i) to true, where i is the channel for
    -- which you wish to enable link storage. If you have no such stream circuits that
    -- require this functionality, you can safely hide this generic to use the default of
    -- "all false".
    --
    -- Note that there are some common uses for reserved DMA Channels that don't need
    -- Chunky Link storage memory, and thus can be left "false". These include the
    -- Inchworm's own status pushing circuitry and the Instruction FIFO. The
    -- LinkInterfaceBridge (for communicating with CICADA) will only need Chunky Link
    -- storage memory if you use the streaming functionality from CICADA to host.
    kForceChannelEnable : NiDmaDmaChannelOneHot_t := (others => false)
  );
  port (
    --PCIe Reset. This can be extended in the top level to guarantee seeing the reset
    -- after configuration and to create a new one on DPR
    aPcieRst_n   : in  std_logic;

    -- PCIe interface - connect these ports to the external FPGA pins.
    PcieRefClk_p : in  std_logic;
    PcieRefClk_n : in  std_logic;

    --Reference clock after the IBUFDS before going into MGTs. MAy be useful as a
    -- general purpose clock (for logic reset with PCIe Reset or InChwORM reset
    --Leave open if not used
    PcieRefClkOut : out std_logic;

    --vhook_nodgv Pcie[RT]x_[pn]
    PcieRx_p     : in  std_logic_vector(7 downto 0);
    PcieRx_n     : in  std_logic_vector(7 downto 0);
    PcieTx_p     : out std_logic_vector(7 downto 0);
    PcieTx_n     : out std_logic_vector(7 downto 0);

    -- Main 250MHz clock.  Connect both of these ports to a signal named
    -- DmaClock.  App hw synchronous to this clock must also be clocked by the
    -- same DmaClock signal without any delta cycle delays on the clock.
    DmaClockSource : out std_logic;
    DmaClock       : in  std_logic;

    -- Main reset. Regardless of the fact that it is generated with a Flop in DmaClock,
    --  recovery and removal should be disabled for every clock (to satisfy LabVIEW
    --  assumptions).
    -- App hw running on DmaClock should use this asynchronous reset (potentially
    --  creating a version that deasserts synchronously with DmaClock and is left for
    --  STA to check for recovery and removal
    aBusReset : out boolean;

    -- Interrupt from app hw.  This input must be synchronous with DmaClock.
    -- App hw is responsible for adding a synchronizer if the app hw design
    -- doesn't naturally drive this synchronous to DmaClock.
    dAppHwInterrupt : in std_logic_vector(1 downto 0);

    --------------------------------------
    -- Byte Addressable RegPort
    --
    -- Address Mapping:
    -----------------------------------------
    --  BAR0 Address    | BaRegPort Address |
    --  0x08000-0x7FFFF | 0x08000-0x7FFFF   |
    -----------------------------------------
    dBaRegPortIn    : out BaRegPortIn_t;
    dBaRegPortOut   : in  BaRegPortOut_t;
    dLvUserMappable : in  std_logic;

    --------------------------------------
    -- High Speed Sink Interface
    -- Expected to be connected directly to LabVIEW Window.
    -- This comes directly from InChWORM netlist and not from companion
    --
    -- Address Mapping:
    ----------------------------------------
    --  BAR0 Address    | SinkIfc Address  |
    --  0x80000-0xBFFFF | 0x80000-0xBFFFF  |
    ----------------------------------------
    dHighSpeedSinkFromDma : out NiDmaHighSpeedSinkFromDma_t;

    --------------------------------------
    -- Interface to link interface bridge
    --
    -- Address Mapping:
    ----------------------------------------------
    --  BAR0 Address    | LinkIfc Bridge Address |
    --  0xC0000-0xFFFFF | 0x00000-0x3FFFF        |
    ----------------------------------------------
    dHostRequestTx    : out SwitchedLinkTx_t;
    dHostRequestRx    : in  SwitchedLinkRx_t;
    dHostResponseAck  : in  boolean;
    dHostResponseErr  : in  boolean;
    dHostResponseData : in  std_logic_vector(63 downto 0);

    --------------------------------------
    -- DmaPort Interface
    -- Expected to be connected directly to DmaPortCommunicationInterface module
    -- This comes directly from InChWORM netlist and not from companion
    dInputRequestToDma    : in  NiDmaInputRequestToDma_t;
    dInputRequestFromDma  : out NiDmaInputRequestFromDma_t;
    dInputDataToDma       : in  NiDmaInputDataToDma_t;
    dInputDataFromDma     : out NiDmaInputDataFromDma_t;
    dInputStatusFromDma   : out NiDmaInputStatusFromDma_t;
    dOutputRequestToDma   : in  NiDmaOutputRequestToDma_t;
    dOutputRequestFromDma : out NiDmaOutputRequestFromDma_t;
    dOutputDataFromDma    : out NiDmaOutputDataFromDma_t;

    -- FPGA Configuration status information for POSC (from config port)
    dPoscPause : in  boolean;
    dPoscError : in  boolean;
    dPoscDone  : out boolean;

    --POSC pins from top level (would be top level pins on an ASIC like in the STC3)
    aCpResetOut_n         : out std_logic;
    aCpResetIn_n          : in  std_logic; --Open collector input from aCpResetOut_n
    aCpSCEN_n             : in  std_logic;
    aPoscRestoreAsyncMode : in  std_logic;

    --------------------------------------
    -- Single-wire communication with Authentication IC.
    -- The following buffer must be implemented in Fixed Logic for correct communication.
    --
    --   OpenDrainIoBuf: IOBUF
    --     port map (
    --       I  => '0',
    --       T  => aAuthSdaOut,
    --       IO => aAuth,   -- Bi-directional line to the chip
    --       O  => aAuthSdaIn);
    Clk40Mhz              : in  std_logic;
    aAuthSdaIn            : in  std_logic;
    aAuthSdaOut           : out std_logic;

    --------------------------------------
    -- PCIe Utility signals for DPR, debugging, etc. Leave open if not used.
    dCfgLtssmState  : out std_logic_vector(5 downto 0);
    dUserLnkUp      : out std_logic;
    dUserAppRdy     : out std_logic;

    PcieDrpClk   : in  std_logic;
    pPcieDrpAddr : in  std_logic_vector(9 downto 0);
    pPcieDrpDi   : in  std_logic_vector(15 downto 0);
    pPcieDrpDo   : out std_logic_vector(15 downto 0);
    pPcieDrpEn   : in  std_logic;
    pPcieDrpRdy  : out std_logic;
    pPcieDrpWe   : in  std_logic;

    GtDrpClk   : out std_logic;
    gGtDrpAddr : in  std_logic_vector(79 downto 0);
    gGtDrpEn   : in  std_logic_vector(7 downto 0);
    gGtDrpDi   : in  std_logic_vector(127 downto 0);
    gGtDrpWe   : in  std_logic_vector(7 downto 0);
    gGtDrpDo   : out std_logic_vector(127 downto 0);
    gGtDrpRdy  : out std_logic_vector(7 downto 0);
    --Tie to (others=>'0') if not used
    aIbertEyescanResetIn : in std_logic_vector(7 downto 0)
  );
end entity; --PcieUspG3x8TandemGtyInchwormWrapper

architecture RTL of PcieUspG3x8TandemGtyInchwormWrapper is

  component PcieUspG3x8TandemGtyInchwormNetlist
    port (
      aPcieRst_n                : in  std_logic;
      PcieRefClk_p              : in  std_logic;
      PcieRefClk_n              : in  std_logic;
      PcieRefClkOut             : out std_logic;
      PcieRx_p                  : in  std_logic_vector(7 downto 0);
      PcieRx_n                  : in  std_logic_vector(7 downto 0);
      PcieTx_p                  : out std_logic_vector(7 downto 0);
      PcieTx_n                  : out std_logic_vector(7 downto 0);
      DmaClockSource            : out std_logic;
      DmaClock                  : in  std_logic;
      aBusReset                 : out boolean;
      dCfgVendId                : in  std_logic_vector(15 downto 0);
      dCfgDevId                 : in  std_logic_vector(15 downto 0);
      dCfgRevId                 : in  std_logic_vector(7 downto 0);
      dCfgSubsysVendId          : in  std_logic_vector(15 downto 0);
      dCfgSubsysId              : in  std_logic_vector(15 downto 0);
      dLinkStorageRamWrite      : out boolean;
      dLinkStorageRamWriteAddr  : out unsigned(kLinkStorageRamAddrWidth-1 downto 0);
      dLinkStorageRamWriteData  : out std_logic_vector(kLinkStorageRamDataWidth-1 downto 0);
      dLinkStorageRamReadAddr   : out unsigned(kLinkStorageRamRdAddrWidth-1 downto 0);
      dLinkStorageRamReadData   : in  std_logic_vector(kLinkStorageRamRdDataWidth-1 downto 0);
      dAppHwInterrupt           : in  std_logic_vector(1 downto 0);
      dFlatBaRegPortIn          : out FlatBaRegPortIn_t;
      dFlatBaRegPortOut         : in  FlatBaRegPortOut_t;
      dLvUserMappable           : in  std_logic;
      dFlatHighSpeedSinkFromDma : out FlatNiDmaHighSpeedSinkFromDma_t;
      dFlatHostRequestTx        : out FlatSwitchedLinkTx_t;
      dFlatHostRequestRx        : in  FlatSwitchedLinkRx_t;
      dHostResponseAck          : in  boolean;
      dHostResponseErr          : in  boolean;
      dHostResponseData         : in  std_logic_vector(63 downto 0);
      dFlatInputRequestToDma    : in  FlatNiDmaInputRequestToDma_t;
      dFlatInputRequestFromDma  : out FlatNiDmaInputRequestFromDma_t;
      dFlatInputDataToDma       : in  FlatNiDmaInputDataToDma_t;
      dFlatInputDataFromDma     : out FlatNiDmaInputDataFromDma_t;
      dFlatInputStatusFromDma   : out FlatNiDmaInputStatusFromDma_t;
      dFlatOutputRequestToDma   : in  FlatNiDmaOutputRequestToDma_t;
      dFlatOutputRequestFromDma : out FlatNiDmaOutputRequestFromDma_t;
      dFlatOutputDataFromDma    : out FlatNiDmaOutputDataFromDma_t;
      dPoscPause                : in  boolean;
      dPoscError                : in  boolean;
      dPoscDone                 : out boolean;
      aCpResetOut_n             : out std_logic;
      aCpResetIn_n              : in  std_logic;
      aCpSCEN_n                 : in  std_logic;
      aPoscRestoreAsyncMode     : in  std_logic;
      Clk40Mhz                  : in  std_logic;
      aAuthSdaIn                : in  std_logic;
      aAuthSdaOut               : out std_logic;
      dCfgLtssmState            : out std_logic_vector(5 downto 0);
      dUserLnkUp                : out std_logic;
      dUserAppRdy               : out std_logic;
      PcieDrpClk                : in  std_logic;
      pPcieDrpAddr              : in  std_logic_vector(9 downto 0);
      pPcieDrpDi                : in  std_logic_vector(15 downto 0);
      pPcieDrpDo                : out std_logic_vector(15 downto 0);
      pPcieDrpEn                : in  std_logic;
      pPcieDrpRdy               : out std_logic;
      pPcieDrpWe                : in  std_logic;
      GtDrpClk                  : out std_logic;
      gGtDrpAddr                : in  std_logic_vector(79 downto 0);
      gGtDrpEn                  : in  std_logic_vector(7 downto 0);
      gGtDrpDi                  : in  std_logic_vector(127 downto 0);
      gGtDrpWe                  : in  std_logic_vector(7 downto 0);
      gGtDrpDo                  : out std_logic_vector(127 downto 0);
      gGtDrpRdy                 : out std_logic_vector(7 downto 0);
      aIbertEyescanResetIn      : in  std_logic_vector(7 downto 0));
  end component;

  --vhook_sigstart
  signal dCfgDevId: std_logic_vector(15 downto 0);
  signal dCfgRevId: std_logic_vector(7 downto 0);
  signal dCfgSubsysId: std_logic_vector(15 downto 0);
  signal dCfgSubsysVendId: std_logic_vector(15 downto 0);
  signal dCfgVendId: std_logic_vector(15 downto 0);
  signal dFlatBaRegPortIn: FlatBaRegPortIn_t;
  signal dFlatBaRegPortOut: FlatBaRegPortOut_t;
  signal dFlatHighSpeedSinkFromDma: FlatNiDmaHighSpeedSinkFromDma_t;
  signal dFlatHostRequestRx: FlatSwitchedLinkRx_t;
  signal dFlatHostRequestTx: FlatSwitchedLinkTx_t;
  signal dFlatInputDataFromDma: FlatNiDmaInputDataFromDma_t;
  signal dFlatInputDataToDma: FlatNiDmaInputDataToDma_t;
  signal dFlatInputRequestFromDma: FlatNiDmaInputRequestFromDma_t;
  signal dFlatInputRequestToDma: FlatNiDmaInputRequestToDma_t;
  signal dFlatInputStatusFromDma: FlatNiDmaInputStatusFromDma_t;
  signal dFlatOutputDataFromDma: FlatNiDmaOutputDataFromDma_t;
  signal dFlatOutputRequestFromDma: FlatNiDmaOutputRequestFromDma_t;
  signal dFlatOutputRequestToDma: FlatNiDmaOutputRequestToDma_t;
  signal dLinkStorageRamReadAddr: unsigned(kLinkStorageRamRdAddrWidth-1 downto 0);
  signal dLinkStorageRamReadData: std_logic_vector(kLinkStorageRamRdDataWidth-1 downto 0);
  signal dLinkStorageRamWrite: boolean;
  signal dLinkStorageRamWriteAddr: unsigned(kLinkStorageRamAddrWidth-1 downto 0);
  signal dLinkStorageRamWriteData: std_logic_vector(kLinkStorageRamDataWidth-1 downto 0);
  --vhook_sigend

begin

  --synopsys translate_off

  --Each InChWORM reports its BIM type for simulation with the PcieBfm. It has to be
  -- done in the wrapper because the netlist is synthesized to a library that can't
  -- access shared variables in the work library.
  work.PkgSystemConfiguration.BimType.Set(work.PkgSystemConfigurationTypes.UsPlus);

  --synopsys translate_on

  ------------------------------------------------------------------------------------
  -- Instantiate netlist and flatten/unflatten ports from netlist.
  ------------------------------------------------------------------------------------
  --Default values for all CHInCh compatible devices (like InChWORM)
  dCfgVendId       <= X"1093";
  dCfgDevId        <= X"C4C4";

  --These come from generics to enforce the fact that they must be valid and stable
  -- at power up.
  dCfgRevId        <= kCfgRevId;
  dCfgSubsysVendId <= kCfgSubsysVendId;
  dCfgSubsysId     <= kCfgSubsysId;

  --vhook PcieUspG3x8TandemGtyInchwormNetlist InchwormNetlist
  InchwormNetlist: PcieUspG3x8TandemGtyInchwormNetlist
    port map (
      aPcieRst_n                => aPcieRst_n,                 --in  std_logic
      PcieRefClk_p              => PcieRefClk_p,               --in  std_logic
      PcieRefClk_n              => PcieRefClk_n,               --in  std_logic
      PcieRefClkOut             => PcieRefClkOut,              --out std_logic
      PcieRx_p                  => PcieRx_p,                   --in  std_logic_vector(7:0)
      PcieRx_n                  => PcieRx_n,                   --in  std_logic_vector(7:0)
      PcieTx_p                  => PcieTx_p,                   --out std_logic_vector(7:0)
      PcieTx_n                  => PcieTx_n,                   --out std_logic_vector(7:0)
      DmaClockSource            => DmaClockSource,             --out std_logic
      DmaClock                  => DmaClock,                   --in  std_logic
      aBusReset                 => aBusReset,                  --out boolean
      dCfgVendId                => dCfgVendId,                 --in  std_logic_vector(15:0)
      dCfgDevId                 => dCfgDevId,                  --in  std_logic_vector(15:0)
      dCfgRevId                 => dCfgRevId,                  --in  std_logic_vector(7:0)
      dCfgSubsysVendId          => dCfgSubsysVendId,           --in  std_logic_vector(15:0)
      dCfgSubsysId              => dCfgSubsysId,               --in  std_logic_vector(15:0)
      dLinkStorageRamWrite      => dLinkStorageRamWrite,       --out boolean
      dLinkStorageRamWriteAddr  => dLinkStorageRamWriteAddr,   --out unsigned(kLinkStorageRamAddrWidth-1:0)
      dLinkStorageRamWriteData  => dLinkStorageRamWriteData,   --out std_logic_vector(kLinkStorageRamDataWidth-1:0)
      dLinkStorageRamReadAddr   => dLinkStorageRamReadAddr,    --out unsigned(kLinkStorageRamRdAddrWidth-1:0)
      dLinkStorageRamReadData   => dLinkStorageRamReadData,    --in  std_logic_vector(kLinkStorageRamRdDataWidth-1:0)
      dAppHwInterrupt           => dAppHwInterrupt,            --in  std_logic_vector(1:0)
      dFlatBaRegPortIn          => dFlatBaRegPortIn,           --out FlatBaRegPortIn_t
      dFlatBaRegPortOut         => dFlatBaRegPortOut,          --in  FlatBaRegPortOut_t
      dLvUserMappable           => dLvUserMappable,            --in  std_logic
      dFlatHighSpeedSinkFromDma => dFlatHighSpeedSinkFromDma,  --out FlatNiDmaHighSpeedSinkFromDma_t
      dFlatHostRequestTx        => dFlatHostRequestTx,         --out FlatSwitchedLinkTx_t
      dFlatHostRequestRx        => dFlatHostRequestRx,         --in  FlatSwitchedLinkRx_t
      dHostResponseAck          => dHostResponseAck,           --in  boolean
      dHostResponseErr          => dHostResponseErr,           --in  boolean
      dHostResponseData         => dHostResponseData,          --in  std_logic_vector(63:0)
      dFlatInputRequestToDma    => dFlatInputRequestToDma,     --in  FlatNiDmaInputRequestToDma_t
      dFlatInputRequestFromDma  => dFlatInputRequestFromDma,   --out FlatNiDmaInputRequestFromDma_t
      dFlatInputDataToDma       => dFlatInputDataToDma,        --in  FlatNiDmaInputDataToDma_t
      dFlatInputDataFromDma     => dFlatInputDataFromDma,      --out FlatNiDmaInputDataFromDma_t
      dFlatInputStatusFromDma   => dFlatInputStatusFromDma,    --out FlatNiDmaInputStatusFromDma_t
      dFlatOutputRequestToDma   => dFlatOutputRequestToDma,    --in  FlatNiDmaOutputRequestToDma_t
      dFlatOutputRequestFromDma => dFlatOutputRequestFromDma,  --out FlatNiDmaOutputRequestFromDma_t
      dFlatOutputDataFromDma    => dFlatOutputDataFromDma,     --out FlatNiDmaOutputDataFromDma_t
      dPoscPause                => dPoscPause,                 --in  boolean
      dPoscError                => dPoscError,                 --in  boolean
      dPoscDone                 => dPoscDone,                  --out boolean
      aCpResetOut_n             => aCpResetOut_n,              --out std_logic
      aCpResetIn_n              => aCpResetIn_n,               --in  std_logic
      aCpSCEN_n                 => aCpSCEN_n,                  --in  std_logic
      aPoscRestoreAsyncMode     => aPoscRestoreAsyncMode,      --in  std_logic
      Clk40Mhz                  => Clk40Mhz,                   --in  std_logic
      aAuthSdaIn                => aAuthSdaIn,                 --in  std_logic
      aAuthSdaOut               => aAuthSdaOut,                --out std_logic
      dCfgLtssmState            => dCfgLtssmState,             --out std_logic_vector(5:0)
      dUserLnkUp                => dUserLnkUp,                 --out std_logic
      dUserAppRdy               => dUserAppRdy,                --out std_logic
      PcieDrpClk                => PcieDrpClk,                 --in  std_logic
      pPcieDrpAddr              => pPcieDrpAddr,               --in  std_logic_vector(9:0)
      pPcieDrpDi                => pPcieDrpDi,                 --in  std_logic_vector(15:0)
      pPcieDrpDo                => pPcieDrpDo,                 --out std_logic_vector(15:0)
      pPcieDrpEn                => pPcieDrpEn,                 --in  std_logic
      pPcieDrpRdy               => pPcieDrpRdy,                --out std_logic
      pPcieDrpWe                => pPcieDrpWe,                 --in  std_logic
      GtDrpClk                  => GtDrpClk,                   --out std_logic
      gGtDrpAddr                => gGtDrpAddr,                 --in  std_logic_vector(79:0)
      gGtDrpEn                  => gGtDrpEn,                   --in  std_logic_vector(7:0)
      gGtDrpDi                  => gGtDrpDi,                   --in  std_logic_vector(127:0)
      gGtDrpWe                  => gGtDrpWe,                   --in  std_logic_vector(7:0)
      gGtDrpDo                  => gGtDrpDo,                   --out std_logic_vector(127:0)
      gGtDrpRdy                 => gGtDrpRdy,                  --out std_logic_vector(7:0)
      aIbertEyescanResetIn      => aIbertEyescanResetIn);      --in  std_logic_vector(7:0)

  --vhook_e LinkStorageRamXilinx LinkStorageRam
  --vhook_g kEnabledChannels     kGetEnabledChannels(kForceChannelEnable)
  LinkStorageRam: entity work.LinkStorageRamXilinx (struct)
    generic map (kEnabledChannels => kGetEnabledChannels(kForceChannelEnable))  --NiDmaDmaChannelOneHot_t
    port map (
      DmaClock                 => DmaClock,                  --in  std_logic
      dLinkStorageRamWrite     => dLinkStorageRamWrite,      --in  boolean
      dLinkStorageRamWriteAddr => dLinkStorageRamWriteAddr,  --in  unsigned(kLinkStorageRamAddrWidth-1:0)
      dLinkStorageRamWriteData => dLinkStorageRamWriteData,  --in  std_logic_vector(kLinkStorageRamDataWidth-1:0)
      dLinkStorageRamReadAddr  => dLinkStorageRamReadAddr,   --in  unsigned(kLinkStorageRamRdAddrWidth-1:0)
      dLinkStorageRamReadData  => dLinkStorageRamReadData);  --out std_logic_vector(kLinkStorageRamRdDataWidth-1:0)

  --DmaPort
  dFlatInputRequestToDma <= Flatten(dInputRequestToDma);
  dFlatInputDataToDma    <= Flatten(dInputDataToDma);
  dInputRequestFromDma   <= UnFlatten(dFlatInputRequestFromDma);
  dInputDataFromDma      <= UnFlatten(dFlatInputDataFromDma);
  dInputStatusFromDma    <= UnFlatten(dFlatInputStatusFromDma);

  dFlatOutputRequestToDma <= Flatten(dOutputRequestToDma);
  dOutputRequestFromDma   <= UnFlatten(dFlatOutputRequestFromDma);
  dOutputDataFromDma      <= UnFlatten(dFlatOutputDataFromDma);

  --High speed sink
  dHighSpeedSinkFromDma <= UnFlatten(dFlatHighSpeedSinkFromDma);

  --BaRegPort
  dBaRegPortIn      <= UnFlatten(dFlatBaRegPortIn);
  dFlatBaRegPortOut <= Flatten(dBaRegPortOut);

  --To Link Interface Bridge
  dFlatHostRequestRx <= Flatten(dHostRequestRx);
  dHostRequestTx     <= UnFlatten(dFlatHostRequestTx);

end RTL;
