`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11488 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
Oc4fq76CzL4QYVrEyjSlCHBxS8pohfHlx1vC6IAFE5jfv0iFDKtFFaIvhGKL/8SW
Cx/sbpbMY1eOycF76FqAK7KdsylyBI/CIo4RTp0bWGa2611Lc6lHDVyA4YXR/owm
Txu174lx225gBPg5GYmYBxZC3ajDMt7nfAPqODc29GcpWUvi4MLh/rDjcgR7YrPl
fTv5/clogLH0w3n6BLR/UoRrxp3VGHd927v3yRFxhnxIV71DeJq/868nl+ISzxsc
k2QC8NChuh4KRBR+itOCxDb/kdixLb2gjoQvdJGW5RLaKOidpbg+aCwP7M9T5nlG
LWWQ9ZVeAlmjr9F2P4/899lP/XlE5nid/OMcFXRY/I/YMc89DUQ6e50YAGftZC20
UOxq5fOKhykxr0U5AfhOVts+3iAOPLsnHwOb7ZgoUF9OFJOAsjidc4rq5WLqdB81
EUP3Nxjkzhk+szpFM823uwmN9Z4DZl53Xem9fFn3jBeF1tKM5+imalExWWy5pZna
yWf2F+EuOueNxgnu3nzsGxfU3YV+BGedowkK+BjAlE+EURjzlAB0Nz7iDEx4c5Xj
njL06UsBUW1ITsIMblvq2jh5FAkCNfEI7M4Unr0SgQ8Bmf6QXOk4H3yWO7qJeeg4
dWnGC9Rnr/KiVgebbkXct7nZrM12Xx22Tz/rPBtVIo0Cbz07CtnzF0zerkXVw/34
siXtFiV3xbsYquC9ZeOFOMFvelOVgZ3XPQ0UXz3HH9RzhDfRAiI5gUSOarZLoMa3
Hl/tkzYJYu+ZZ92pLYcRQ2XsbvVb1gCjTms999FOyQkGBcuhIe/e5PHqJzYBfFLR
kEmqW5O9p8GKjddVC/HcDV0xfvDbk/eRXbxqnq3LKY8TZa9Aot10lRZlYmKCRhke
OK9CLAPNnDxnEDtVtqSaSLmfYJfwgQjp1OZV4F0PsIUgyTs5OZ6JWpKo1y1x7b3h
buUwwgHzhiOo0UJfAg333KzFgLK73P+rNHyiUmhCToKN+9MEmU2DQhoxINQDhz9g
g77bYdpavjRD0C9JVRUn28N/AjvlgYwZ8LsB4twmhJEYzYnPcTqI76XGTLgXqddt
xXi1/51EVqoW5HT9Kl//lidQ18WdxctJOcrgWPwU9LyYu3POvgkl5LXB+eZuexz9
8oXlkY2q68LMzxr6XF97vZ2HhlmAr1LF0iH4Ohi2JDQE0c/CfZ3FPBWYakRWNYqi
EIkUScBLdu8/XyMIjkg2hpbADjbk/U8RWDWM3kcc2dpjMglzmIbHqIDnlER1sp0J
RZBrmBdgl1JEt/0rkKrheqwM4Ur+1mR+T89BsdcYnMRP+LVS+VTB/uvNNNGxm6Vq
LwtFfycVuDAccsy/lgELV2eF2Uo+YBX1SXu+seR+Xl3AXCUSRjb6xSgnqsorHoo4
iWHTq7a6Tf+h2wTaDE439Z1spHpycQcgbAgYzukYTf+88N8O0221+ixYNkhdjY2Q
3QA8Mbmowxiv3sBsItWIHnpDnIzFOT9G5UzDAgepJwmo2IigIa7199fliJpHyEOS
aS8W1rTHTefJB0RjNtNVKitkJiapFWEy86EkTVfMSAnwaMWVsh2/gzzkP9Jigoux
WppTxUZpGmIOTsV1e17OiWlFrg+tQkb6r4ADDQ8OpX2SzlBOLC+NevHeyCQYw16e
Ahkw+sK+AUzMF0vxZey3APVwBSYf2UDlg4/IW47+JnO+xEHtG0CuyDb6UFJVIaTs
LLzgY7gigOoOal0kOWZ9bXzdk81wgiyqD2fQx3v4N31aBTrStmZT/DxCChC723+5
LJVFJZkNiTFqURXZC4abiSTYE23cegtoD9cGtNkaUn/QWUdPAXrJroe9O5jDw/55
FgAFGCtcDB+g/w+o2uptAdYrYdByrxCWtbZqgHIG2ReDuF8fBcLBgyE/4WleOU+4
D6QClE2ChknPfoVdnDj6H0MMRxzHakMWTeOM8858eUxNxw0RSWA8VY6wyrESUKFp
M+FSpuoFHMqls04hFp0aibBTM9nHq5+GpFE9IoMcCsWwe9vnKc8/iv9U89NA6o8g
7VgvdLGj4ifwyu8V6IclBUGs1YZTShD5TzpBZ7pUJCnk3SsoHPuuGU6XsmwZE1G8
HqNQXTKN6LAkTL93iuyFISQujOMoYqiXz22hlS6vCrDUkIZVokbV60h/N0RYniqz
33rYvK+FcyE6g1mveHxJZWngH0DcQoItIur3it1E0D9IpibWrrYBW8tTsA7CS3BY
pb8k7B/ziX7dAd0zoTrXIGWISBJcQQ1kWjNFPuYD4ZD9ihPib2meOjsiJkd9XJAw
fQnjOJhtrf+/RCca9W5TwR3BOwzwRaZCzVVmcMlMisAIDMrTLSNw8nN9rO9gFPVM
bhoGRiSLoAt9POktMPm4H35fXiFn489N6GvFg3Do6wfRF9TJb5dX45RSgYF8ef0O
HjbdQyMEUhStLSOJF4QUL8j9D4KQ5sl5yLZdxnco8lhFd6y4rnaxLQKCZJC7FT/p
FnCupN/twkhDILgVPVxqkH4Vmu7ZIkeBb3HoNV1NNxRGUevTJykRaKW54ihuNItz
9qKSQT9EGrBwivKm+9fGlh4b1Nc+YxUgON99mZ0D9MrfnDVCbY39c3Uj37dULzOl
IJqNrkjG5d1hqOuGfGnBn9HuSFACw+dXXBv2iC0RCwZ/3bwre1YArMaJradLk3++
CCjA8vX7jafC4tuBlpSAEls2vhhba/pQqmRdyyDnf6E4LxEJE8uMhm9DyPlUBfo/
FABJfafNlbKvLTSKf6dBK1UdujlxcF8bOoGVymAtX5Dl9nFxzCbvl+lCfSsGIKDp
tAykQIOvJn77BwriEBiKN/LAA3uRK+aJEpzach1nR+2XIIesW6HmWLy0aodzfGHV
zr/lLDzXKmeMaIV5y2G6FWDidzSAljL4C0/mMTkbcca2YCf++OnNowc0couFemUY
RYanm+ftcExSgVoHYLrZDAVLNb39movsqR4WfAR7yknr4pLBeXZIBhU6mEREq58I
IYmFR5yTRtMTO9lHqgxiZccw58ShkcAkuCNC/u7I0pG8ndE9hs+3+CunrHiSMonR
6feiQO8jw2q6x42mIS58nOtd4nFxPpU0ITQyQqX3rKG7nfxpdFh7E0mkMtNUroMt
aGox9RfWkBdOasvRoRZ5k+eflsxV3Fs+y3XPYWrsH9Cb4zjT6TvFHHI72a5+mgf3
5g+DVQyUpBbn7WyYOg8cYCydzOZIR0Z32K1IV5rmwaogWGkGn2XWFEJ9oSfkMkKl
vn74xT9BMWws6rcbZNJgmcTmIhvkEm8IFZIG0cQs/qKYTbq3Vl3CGRyFZI0rkn38
4RqQlQPu3Oum9P7ozmbEv031nRFkZQkjxmMiRbQ5QsC1KWnitMXczOsGldSbe2Zg
Owrlr21I/gGRNUCO+jC3ki+lwz97sxbde2JAvG9VN38KZWoscED/ma26vdswtoiq
WF28Pktdn95xrtf3MHW1VeSzkszFKrTQ02O5Us1pQgTESeWhVTvRxfimsZleArqI
ycsISY6Ag1tnEnIg6cISbzvQASwaoeQKxuWkN69lEqUZw16ffdr0/nR9LngLiK66
/2LFvI+pDKMqd03pdonAniMpTqJnCNmI2SWs+suZp8PNWPr20Zd5EOuPu5irm0AQ
xARp15umXAOTLB3/nLUzXzgCa1MKEs4vleBvrqKsHNZSq7CGdyNcGcWUbQwh9JPl
ibe1F5U6iLRJJ28F5j5SUWDk+KreCGLRaJ5mEZDQIXJYqzP67jdCINjYq4WNeMoE
DsWxkzPv/Qd90DZP16lfsnCHcwvJVDltT6kf5K0PeLCkPJrZ59ZxqUPJVQCGaeyj
ilSJnDw4rNGDr/fYpWX+9KfUFOJ8CA3u2Fe6dhkdeA895qEUlNCBinlK5tLPiv63
cD/QhaVA63OgGTb6OtPS1Rz2NPGNtEPt5aZzU9ZIiHOFTiDrAKaQ2kFN6/OKbMeW
rKpleMuTdrmnepESuPU3TotE87Q9aRXFHFzrnHMiVGfbpAg9QDKUzZXyI+CnqUlY
yWJtALQWXFFrhTNM6BPnUux8373wK1dK2vB5I1ouHOXkTMZttew91IC31Qq9oDHY
klKxB7/kQdp6pakFDX+8x/UUhLUdkeqD+LJ1eG4Nxmn9fERL4tRmqHYaP8wSyYZS
ldcFCo17/lgNnegSLsmcuALiuk88UguRHGtIPR3wCfmoL71cJSS/YiKZyKn1GV1Q
feqf9FawAJ47/d9vb/Fx+JJQVsvFiOeBuj7A1BmgUeurqkrNRtvhQAZ/WnIbvNFb
gtOxCuitFr6LspWcLzUh+TpUw/eWvSd16pUM7coQQoDPlpO/1a1BOWfcoBoROOMn
Y+3ddtpsbJGpLbvO3t25drxPk35By9Gv5efBZq+zuTDIZpKTi9+1N3S7JSCSkjFI
xIl4p5M09qCYPzK4KWvs3vn22eOgbqOKw2SOZL5g3N/m/q+tfwu85fCVDyye2sLN
lqISaIvnsBED8Z3oW0jU1VB3jUMmoKUH4Fi6Rs7u1dM+yzFKEzz1vlv/Hk9rAXAy
5jGIw0TmUk+rhTs83mGyVu+27cyRaxE/D8ngvSJGZ4IeJP2lDr6kFMpoLvJoQ1K9
PCHPcZtBBSEqAxMvsnkxm/1BiAc+snxyWY54cQiChEdg7cMOb9OkCDHShrEGwe/j
vHG0dQUPv/hzYkzent23yYk16DB3DToiGWdOr8tr4thjGt7N5U67L222fdRBxo0C
7LsR82JXvINVzAtfjdpO4V7+2OaxFICd4laT4xbncqpQEzJt3PSTFLAhwxH5/otX
/hFcan/nGD13BxRS2Lccy7jL79KI6839CXcPutWQws7OK+2h/5ri+mLv8blCJoeg
+hCMTxt92cs5FQ063rXqJkgndy2yAUTrHhLG+QzAGAosYrOSjTA4GdHqaTuu9s2P
uDM2IUTxNtWJpF8waC3f3MEtoLOdJae2XO8q1cwgX6F6yVdAJx9nXd+zhsWSudh3
enYw7ESi0aT2CGi+1mVn8xl7mzR8riRe6nug5S26BckwK+pL26RJWvyIQX+vcR8w
3NAUtylRQ9GM9Z2cd1PXxLnnnE6xfEluffFUmfGyWg4HTTgXHMZaLQkCFg8neUWM
KjmfchZ7QtUcgxaw0NZZtGMfqyajZrmj2TW20XeuQ6Z2rYfkoOEEueqnzo7lLkGV
Jzbewn40w1IM9LSvldVT3KkNOeoLYMVbn5eBrYDXNexMIhmCK+VMzPAWsW0NAMtj
txd0/hfK2HFEnQhy4U+QJ0a5j089Z8ebTlZiz2fMcRLywiYXj0BZ4eV7Awn7kRG2
4DVQsMhaNcJkNmIf8gvCFU9b8MVoGTPjQy4DaDB6oGpMqtYSkpmMN7uiAqMX/q54
hDPMowj1vaP6l2CHuaXr6s7MUq2hllmzR2slfEYvMyqqqqm+414Wc95lPzZL8knE
95p1WquR/sv6MkTvFXNqKx7flOvEy5C9bKyUUqxUCnDJFKgzy0Azg2ZG2Cjlqz9Q
D1UsFhi7OAuVRNUJs9LwMcMdmRGjqjXs889JjNtzxTN7rZYp4jvwTu6tNcOIARqT
uGCdVZW/RdlvG8hSTx6R7DUudVB7XumXMD5M6AK9IGu54r/ry1B7t11Zaz+b2D7K
4N2SMKwRoeV++wpYUE/a9X9I0KsLBlJmDh6NjSfwxrVRSDAfSo9mFVkJ6Zu8fzjY
IqydpCFQOw1EpZitAL4zP1UBa+SQGSV67ZTMqj9Vx/13joXN51tarPuvVBEHTPX+
JCIpWCXYBiCWPrErU8sJniCdYbFOJSd2qzn2Z5lbu0IS8aC2/AjQKy1KqH8tjhGF
Za+e6W2l8HY1LmYbdM7f8twiaQxnz5LNvrtCjIW3aZ5O1xttS6hU9XkJOFZVWDXc
7OpX2MpzRSEgZKvcDYTTDFCTI288qks3XOeL+sv7Hm8JSjynQjU93NN0cFYkkOn0
FpVN6P7OO1xxJmqggyNFCvz82QE6+gaCcLQDtvoq9vkTagZmzqhP7pWeJJZyocuZ
GnGy0ZHEGQN7b83vCBjGC8FA1/ppMpsdp1OmtajRG9jK1jnZcovzh2Dr6/wgkMio
zjcVhEIFKPR1GM6ScBTo5H8Y2fErKljd2K1jVL5lRUhuvBbkxg4Q5YFNRWljkTiy
wCttfOQC0IQM2+gSuPUwSIWBJWbwiQ1Fdo1KIwCejizpR2HAdake7gGFPTaj71eQ
UaFLDstbRXBZGTy/u9sVySv2/XiRK9dmIS7My+CS3fZ8Gec0hWWmRtZW7elifz4c
SE6qWPmUrOYs0eZEwNdduy3aKS2TJGKKIAhbVCyMj+H0r0zQ78dRx09GJY/Utjcj
CA3fKXuEeZGp4cH9nUZ8ed0sFApcWWwgf12SxVKn2URtyEbhBatWxNmIxcGv9Sll
M9iJtUp3GFCTL9qwBIcomi/4aY9ujaHg+xpSTTBbgIHwbFti8i/G7bK1xC7IIiPy
mp3RUFe4cFMyD4kuniweMxJUMlnlJyspz+4YoZocZWfhlWNCnbPCM7kGGgUVjlKb
tG21vGeQ2/oX5KxRb6dQwHpcVKYkLKGudFoS5dItBUHJOvi9t5EKXoM+zbwL3TpR
DcozfRjKuv4MHoOCmdy54gcRlAJZUQ6UKAGmWHNcu8jCv+pLtQmn8ECznIOPmuTh
XZia/JSf/KR3EhmZqr7KRkkQ/7VDd4TiHwOJvuiMOZWAfK3CgIzkjiaB98cNMYJz
/Ov4weZ6ue0vCks3fCvc68HbLbzX+93FIaKPJ5SwgcvBZkv8DKxe3rDcMJtHiAPw
4psjyl8w/EAAAt+DD9aQOPuaaAQfSARx2ZrFveG7Hse9/4mwxAIS7tqU40N5VzvM
KhTA5qQ+rwKbwo8/qWr8TbrH++I3yoz/dzb3VT6w8D8wUPtf6qTzKaYqUUQy3g4s
lYy7v6uceF+TEMdqugM+3W9w/WRpl88SBfD06wY3RfAd87V4FyLSRUvN/V3fpunm
0jvTuRPN2HTT/kdDnND+mdFmQtCOJMEEHDNm+AjWSfLTHFtlP8yIn0/S3aXY+tMp
LXpfE39i0iHViSvbulbgA2cLy5Tzbkkl6ssKH0diUxijZkbA/1i9W+lLdWC7IsMG
aB9DT9bbAyiDrMgRcte9ewU0HkBFaffGDEZOWM5CQ4vhSnuQtJwE6xYjGm6fQCuR
GhxAcgO7h1ERHK+hhb4k3CyQ6hc8jvfrzLc1aIP0LUYV09OU5YjuMf9v7fPKbcK8
D7h0CG8KsAi7S6xsMs8tPpaEFEvoidJIs9ZWN5PqKQkvt1eG+jG9rYZjlGc4F3jp
SlDKBcbzwBXJIbAzjizBhvVtvt/PJ4RcWti0GkzClQytd6/K8/XM7s+Je+bSmQzO
MjtKuKdgbqpuC07xa3xXKAdX92JkpdsK2Rt/fbf5WONhnw30Z7Hw0WAFs5DiyFU5
C8GrbzESDGF5Xcdf2kueCOo7wfxvGH3vNTpBfm/yFh7vSYFootD1YJ2M4GIsIB4C
qlsCEnH6N9VSXFjQ/uM2ekNRDMIL5npIFYYlEjZwWIVO00P3E14DHIbBLN5wNWGX
Zpfv48daVpSro5hy48xs/muHFDiwwv3DTZVF8LnjpxWqZ9R5f99AXPSCHj1XpKqE
KykQCCvP22xj+LF7iNVne9wo18pyXGeEiD7vIF4NziiyNwbYGdlG/oMrUPRxslhC
nM+VM9+TZn6oVAUYXAtd+xRcjqrpg6fETbKecnc8RuGnjh9/AvH8tjL98xeDELUg
WZkVW7CCaS87avw90ulCRi7AhmI5QBML7NiUblaAhJSoWt3feoBeQLb+mwbQ66RO
g39Jy3c3yfeOTV/Xy9P3cEq7KCiVd2GXqUi6+vClLHQ2yvMe+XaGr2RmK6eJ4zDr
y08WXeKtA73ooSopokeSXg5MUs4u91DW1E1Dydo6E6R2yyX8Jc2l9WX+LFZuLUQL
o8Zv+QTLd3omCB18foPwVrQ+ulxTwwH0Ytf5XW0WH2U7K6vsj2/3m1Srb8z7PKfY
D/0o2GrSJogFIZR/Hyrem2wpRNPhsAWQrbU6fk8lxH54bIzLvgGFukZ3pFOf6FIx
JTa1wL+oU0u9DTSl0fiGwo4nK1e79wbUKgGN9lnxRZjYkZscfdfxfw75/bVWap4k
KLVLcSVs7aGibOjFtx8JDRECzX4YfxhcGuWl0FJZNGyBhW1kENOIYn2edeOL8BJI
VfOCOgzwPukMhQOtr/2LIB2znLMoFOOuDl53MIOAbvMiHv8MjKq4tWE9Q7NVtAhV
mSN6/SZysDRL3XTHNHPbgOB4L7NT06IvGKBh4A3ZiX4MJ+0qDaqybfD+HSyCgVFC
/fZ5doQ04BZcPw/TripnkmSia9E3Muv22EsCR/N99TNA3LQBk/iJQZkSKpk3JA/E
Z0sNstRYwaRAj0w+eEC7l3d8KdsQ1NJuaSYv+D72NgC+yozWo5+PBKGA5i1dvqo7
PI/SMBOfLN6qWVmUtYnvTmUPZUf1wykIep0IjQ4putUU03+lh+AiTQYFDIUKAlnp
p+R6KG6HuR8/yoV1fBv32Yh+Zc6kRgluJxWoAmt/iyts6FA2jVQT+Fq3DLZMVjbn
C4RDeWaosuLTcpwS9qT+AYc7E55RCbJYNmFJdkICdUntw6Go5IpbBKt1FzDshACS
KjEpm61xYdNVT8LsCDxtdGXeiYZP3ry4ZiNbCJ8K36ssZVJshhqpQbONqHscmYRL
Yhwt0dLdZpADkwPxDav/XulLUgcB89FYAky+/EKwDj4izy2wbBIhvoaj84FMvNVI
7A1YCam0+vaKlfqpMdALyQlLJmeG/aBxqqYKLMyEg9xDp3BktbPeeLvgOKT4Wedq
86G+NqxyvCbv2TNvrSxHY3bt0mPgAuVz6N2i0Pd9AAOFDD1bmytOliwQ472El24T
JOtChYsjR4RzKIX0lI4+zvEUsw5Tx0A+5DrCggfoIeqBeYiOo3bYmraH8Ar94umA
06P9yj86v5CjNMz+8lNDAJjW4FcnYVyO+omkPGy2MjjoztzzGQmloP5/PylJNEvf
M8AxxIWRc/uWWq5kPRc2gbE55uptfrDghPgQwluGBOqlLOBp6SZaW8KFBfGeDoLj
WkVTsLozvVQus7rLIdS0SAzt3YIzHqrvEtObKrOUH1+7LHLRE7UoSZJ3VFcGh5Py
FatBdT5CLfPJU5B2hJbTpQ+Bic2Y6JBgXpErpyizk2JT49j4XjvjtPEttrd2dJnf
LTw/hl01obqG7AMIijXe7yAfoZMELX+W9Wm4BG1+7SswP+cXm14NtpRHTMsuwNY4
4u96MhjyQl0GsWM07Li9L0kpwyUmyC+/T4apaonT9WtAFjBtsY56BfeDWSXZOHiV
LfVStpKvczwG0dCApf9wc7BkxygWX/s6v5KJYd0t4WAPJDFPSjY33ib2lhP6wip8
wXVDk7MojYHM5RNS2ErHfdAW3Gp0NTGIFlY/vj+LCW3bnh+c/IL5K436xkqAauBq
nz9EMH9gUWCUxQTsyqh+t5DWSOYTNqgTKbAsU2L/9ZDURUIRuwuRTTCyYtdFp8MM
bH+tjSkaGWjryz8tNptCBoCDeYjBntXMJFEo7ajyuyOBPzlpBo4Sb24GXDcFaCYo
WrI4hbz66JUMADSP4+n2EqAI658ZqoVSWOVdtevkc7tFrAxIzZwb0Ud+644YJYAZ
yB/Gkhh9TnGeRTiPQugKeXgaRdrUNB3/m56zkP3ioz+ZHiPUSRB9Nx2rst0VV3p1
gZd4sRqGVEm1HS7mFW2qlU/kLpx4bJ0DxK9fMx7aos/rv7OPTByFGIGSTuYWynHL
+O+oSxMI4f9k8cMXV5iMz8vBQ/Zwlduap7sa8EiShle4uK0mcDsaLctSrue7rh3r
84e4h/1FqeiAqB21SkWEn+FFkg+M6FRgjDDl+/qhnoXSCoOivh8rhws4wrr7d8ot
61dwFq741CpWAzDkfRwkIkK59sNDLt7iuLJFoHhMYD8W9vMkYWTSNPmJc7JlcEzJ
+UptpbDt2o+1YBv0Dw6qByw0ehWH0xUWFcsOk1WKBfsUjO5srHxWwz5YzKEbS1Pe
Kg0suB6QksLS8C1Ba8XogzzaToXgGYwYGyTDdk15lqtEw4qhmobK6DSx86JIN0t1
ODowDvdW3jsc+QA6QkbqggARPghaaJFY6yEt5Ai/2JwrRg7oKEb6iDVo3qf+xXFy
3yB4gfyaY/8vH2wpkdVJW69rPokZ5H55Gr//lAH6MG+CvoydfI0z0/QwBhCKd3fF
oZ1Mym3+hReEwV/lLUL2zxbs4wBTpaDF5s0rWLsmpYfY8WOYxzVps8Zi354+zPJH
WhxaPvyco933Vtxdk6c1KYqtybLX47ySd4etPxWcnvYenoAKD5la0B98rXxoCZDo
yL0VCLgqcdkJjMOU2YWwf/bUIwDmVHGFprvsPLqud7dBVvKhwX5QtU2EqrWt/19G
m32nnhTIhRFF/VqUS44w43wQsmlNXGv8UpahYUQMH1mHnB2IvyihUz1MbCNDXf0r
9iPkvD3IJ3ZSv+H5FD4lOxWpyZY5IrJ+G8g6pRCvro8qWO8RUBrQYGOD1AfhKdGu
/wOyutJPRGnvndlMzmVmvwOJDR3BKzqmatIaQnI+zb4tvy6NT5nin66Ci0aPPZ8e
W9FauVRjew/tgyINQ0rBdlKb+W+0vcd/vBYDLMV4u+Ad67ftFVHoAN5ItOJ7vusk
cWUYt5CHTespRJDtID0M3uUmrLQ10R92hxlSd3Yl8I4G8p48VttNBEWLyeQIjfTi
BZ/2wAS2BdGnjTpxaEfj+kJX3AWcb74GDs1uzNz4pDZYEf9JR6u1XPD00xEajATo
boJGHmpy9u8HhT+QaJSKyCe5J4bFqLJy2Q9KFXVXT8rWBcAcsbeUNYgqQvhQpwEX
jGQCEBC51acgMPNrRbC+8OjObkUWGdZ72+Zh8FsRFOF62YrcDp/crGUjAvck4v4D
jK6tXHVu8tIJ0BB6Js3FAbA2/HENDKkXRwK3P+Y4EOJqZIKgWP246c272bgHcZIV
7ch6UOwTWf9MRMv4pKNVx8YK2dC9gK5EUYs7+/Lbrds2t4bpktUaZ5CTwNb8LYnj
scXcWa1NUOzAVseoRyuzaiQPl2UN4YFY4uh5qYBakVVVzDnl7pel+W3lxhWzFuk0
hSvjcpsHbMeovoi/VP8iMMM+ABageYyFKpnCRqv0lBGRHbRObNxmNCBplFhaPOiH
abPmNjJB9RwvuNsMw1CqhfYDwaIacexa35u3UxgWVbHGLkjTQMdiiF0uMJsDbL01
lilU6le4iNP+k4wKHSFlMvLIGbQzm5VA4HuEL/vlajVaXlUbw9SMQbPaIPuAzE0r
mziU1v/DHFtiEJQFuHOI6WfdyI7+qZLOyIJYjsJiJMSaMmed2mDRx/PAyhR6kQUy
xX6m1s78kv0nROOIRzs0g79w1xSSMtdICe3NXT12fJc4XuVe0yX4dNtQfggi9J3b
z3qWoDJQUukRd6MxGqOb6uXI3Mj5fgZRZ85Eh6R0EoWSypFcFvFncWWXC7C5np5c
NuhpPMyfQDmfZYWVsW499oxvgcTE6NSPoAy9+W0pP0qGGRzXU3hE9hYPUIGc4s96
8F/nXoFKxZV7vYl16r5zBlik7ezlUqup4i7B/g/U1uICLveKFoPFFMRtXKeZUF92
EPafE2ypirDPdtvISRyb3IwZkxkliVRs9OvhMYEmWcAguAPGifXl29kVnQEEtiZX
E57xfUaSsjZjJtK3FRNDpnlkrESHeXMV1agO/DW0/BXH+fRTf/hCAdaOb2EnbCQX
8Zc2/jYUHX24hMJ3oaYW4PwDfKBIoX4Ze9J5dozXaZd6mr5u5b+BBK2UQMfIcTUg
UBN5h8eCbVb1xcg/ec2PQBiAMulVSEQBR4JLagKn+3XLPrAgSLcS1z+84KQ0EcD0
PrW1cgBcjRyH0vLwDCuK9KXw37IM1TaP3jOSBAZFxy4yHkDbQYZ4VQSnW54i9Y61
8zDDOQhGjwoJ5/Rv62wokdEq2V2zIX80KZYHagBcxxNle8aVlhocsvt3mfQ1QGdF
Lj3YvfAlQHjMHl/UKX3hZhucv0XiHDbFCAm341gdODx8izW5TGeKdyJ8y7HjL8Sk
5kkn5Yjw3OBKI8XqsDu05pf87wUSG7rzvqINGhckrK0JlkfMsLLPwEc9hgWXiCJ9
cJ2jSqlV7bN/KQSgK/WeiQfOIw1/eMZJmLYaVABeXVlffLiO0aCd/+Jii1K2US4b
v6OeiH3yOQAFrEEg4OwVdyVcu5uXh9piD1roO61O0N9axkLxOykFwkp3rvzx5jOT
tWACbBXmghoqVX9PdAGJpoQbIAb6IG16obuz+s2PmwRBhTVD6IeK/5NOYNudGXG8
iLzFxxaFfmZvrGr88vqc8BNZlBZb/+HaeXykiCq43ZgqD9wGQDd52RTtcxwEpiH7
fnHzoPl1nYbdSwbe8N99O4GdqJwWv/1T4IQu36u3gL2NUeDskVWs2FLYJbCcKQol
Q8ZU8Kl8CkHtZApEAPPiLt0+rkJqHBYYRDQVnYzulCj8NPBBPaZJ3nAIphG1dQiF
CFuzaQGkZnG9/NTSTHoi9tFTolHCx4rC+mCSmb7G7/9COOFiFhqXts+VC+O7n315
XT6NKAYSW9vufc36MOjp7PBPNRCVXF+Tx3iKEp23/KZlYh4i7RQcohAJZS95+oXw
W56LpEKflKZpaMH9bBXWRNJL915y1IifRIh+7G35cOCquTolYMMl+vRh4kDh5LiF
KUaGA8ZXzPAZWxMcuGB5ROalFc9qXK6hGTLxtM+rlEjFJsJCHEOTEmNQmEMZKs56
a7DSVd2HFL/oix8OlYLj6A56iaptlKWb6LLP/m4YX1nZuBdq3N672gBAwRAP/1uA
Au//pGi33SN/QxYw522HcfbmRRoERhLPj8HwvKMKXbuhuGwGbEVUu+hYS1wG8rBh
aREF5ZjiGqOwGhHg94u1EiqBjdoHEsPrFD/ho9dgZoWtrAafSBCbP3lUmLPha0lN
8XGY3e9PLTV/Fq5ikpR3ZpQMZA5y1qRx2XTLmqCZauQLdkyUstbOESMlvKuyBP4O
5Ix2Kf4C7jes68o7UfLmQggbd8eTuRFnnNh5eJXWyLFwpe1KPadXSS0VcVBwjgd7
eaJ3pBvotX1ZLtrfhgpyepq70ttthShVRuXLkFBV5Tsx9A6iRdyYH9sWF2HDlMRF
i5KziesgvTxPibEqSZhkIPxWctGrrafnLHj30XrDJzAfuSoP4wvrlh8iMBqpHLPw
xKngV3on/HYpW2+SGzOnwC6bGYMdQMVQISgYvzN7V9wEmzRkrKh1m7eD0HnPLrBj
IAIqvgwetX8+etc4gHjE6SfKbMI/IzZhTrN3ZFpQcme4FxkGpbbSPM4UooXA5YNb
airrnqJJEUA01yjesS3iVY8yzUUQSYlkQ+MC+oEZbibBUtfxzV6z6NhIdzVonrkt
J9j6LwH/BwfpGRY92urpvpEn/1IHgmJ2lnRvDPR0/QuvYMsPyHEE3yHzK7U4ls1L
1iyCjQS/fLfEwbNU4enh37VRP77tVSVwS4z4bKPQ50z/hCzMuteTQSeyTFtGbY6e
WLyXe36yidoFF1YnWAIRYopb7jWLwAqYXoT2wtiSI1k7MrYSBjAUoYTJ2tIXGOKq
aKw15630/HeEFqtH4ZY9BwJFBWNtKiaBjQYvNrJfpVWEDYK0+ijVA/Tu71RMGifz
LNQtQ3mP9cT+QZ8K7w7c2eoTxKXIlrs90XCiXR+jff9syVe2KRJ2OlE9TadhU6DO
k9nDM+bdVzqHFBxJ2SXHC4knK0pc8HxlafTa3jjfp6ktYgIUPaa+1Qg/DkprfXqF
xHWjW62CMUxSS0qJAxrLEnirh1nENtkQFvIc/gC6vgs9Eia5bLP4N9nVuIR7g7Lh
hnHxEljI/gAGniRY8XMsX0m509D3ylctW8AaGckqh0IKPHAdlRDpisEHidGZc0kk
ktXDd/nrOajlvGVrThz5zRpvPeCZF89SDqPvRlfK4yz9EwJtH1And1340QXE+8sP
8pl/hh00p6wnoM+qkYQtyB0S3blgipY61KTojJj8bFCZNLou9ss4S9R8otU6rZ25
aJ2Y86aLbBvZ4Wu7mehE1+qislKhQSGR62WbeTRHXIA61wbQanQ5cqsR7rWeSqK/
6ddNS0165RmAki48attkCph20l4CRzY7UiKEbr1Sw9n+vTuerYF1K9Za4SboukvO
2XDsTbqESscX7Ta+90alcJFs5j6NfBYZ31d1nC94IKp0yYP00ouWUNNrTEzIwayj
ThgXwf5lOdaoXQ40xOiFpF1WNS5gDPAdvrWNKegAJrCWTZagOnmZLQfGVNXllxxK
OYqBDkuW8pJuFElDEBSOUuSzhjn0fStfLOJDmszo8oohYM8fp633CT0VwVeuUMSW
43cvX93wG1HRVHVom6d2Z3RFFN0Cnj7sDT73ce3ALXEw48EwOS4Y4UlZV2rNsZ0+
2pJ8iTKhWWrg06szxnqIcdv/0AjMhq9ydwPRtPW+AEpUhDhqSF1mSmHDNDcufrnK
VUugaLKkjkYmlDRuukLMHdaqW5S6WsN6TYmVh/9y6J9q3UzKQsgDNJ3vceA8Xxln
XVfSm3LK7nHx05P9J5yfqBhyKkY222G/5VlrFEIqtmzxH3LQgqAPbD/RCOaFop4L
hkUuZmmGHhoHFqqPOK8DG8vgRWdYMBDPipA48V94BdeXg+orE8ze7icH4eQ50val
2Nc6TiDUSHwGjhkFPTN4wDutwUzSVD40d9AbtlW0TX5ojylobjL8FUayrS0QcdiO
dKD0JEdkHfb7lRYti4N7jh0Ln3bF7vXb16LMizxcoxqDWneZA6ZNd9/3jIWFei8g
Q4q88Y9RyU0FgqTHEa3LsYq+J7TWlmMl0AnsY9Fe312VcjInLdu0RPmSlynkrwlS
6CNnIxGTdMlXgrejywwuo3FqGCoHUfvRDTdpPezLjFv33XhKLkagTaIt5uHEfjEI
sf5JgZ+CvaDxgr9Z08p6xyIJcFPT6D7fbJT24O6l+gsfWgcvpHmuYowzdeLWxor+
84ISRhNUk02JQgywPSKY2bHmen7pkdGXpH5BbFeG2Dl0YyOAxCvO82Je5b2b7v9B
9I/xzDbxxenjH6V7yGqlKc8/vSUsDt+LaOxUjx7DiVq/se47OdlgjGafNCrHlLAJ
RpRh7rPMHJCHerkfnpjBHQ==
`protect end_protected