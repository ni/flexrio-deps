`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5040 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
1z1b9VGiiW9Gp7THxpOgEcynjWGi3XZIF0PEbAAePrx+arPDK9UM9Jagzz3ASATi
vLzEprmKT/bzBLuD5tSXD2sRNHBu4QubcwQmu21fIOB/CkK/wM6iIGwIFqxR6xJ8
e8YriW3nZNi4FU/q5ffiVjX3AtyhEi5pMnykOFfDvm7TURvTLdOdv++d9qZQp3HP
cQSEORHE12AowAm8AOMEXGCDxfxtC+lNCgzSifO1GPoGCre0lJQx7Kx4LDt0Lk54
oeyuvrFRW2nmPQc4G6CWdqOskeY54CYIoHqE4bVRToUaFJsPmotjd4QHFHOrDZ0q
qjGQ7V06AM1xOE+UnVJqoqcvSLh5mJ9IHeRlWzdaouXc1rYPo+m4lUzV2ACkeyUr
dAf0Fn94gYVcjfMMy3mPUcRRFUwufUXyo3Qtr+CyN8b5fEioRW08z84uCcNgpnfo
EzqR3wzdG/iXMXU7azZWfh9KlcarJjtraRIbo4wLBgq0BTTcVCPTOnqnDFjKpIrj
ZiiGRZe/q/5bJOhDrYtXtvTEkYd3cZMaH2IHyuu9FV/2lb0cBV5kU54VCqqCx3Nz
tit5AkM2miW1yisKItakOTZjsneQs+GaO6DVplCsySGlthP0wvRJ5KafrA3AbT3o
DMGy/1FxCXkV6EJGTaVeVESGhyDyeAweA93WHHVmZE7SzRtsJMzc/u7WUHoF4Vus
cse45KQjaF4CpCh+Op2ewv/TLMsE+Is/YxmlINjEc2Y5qjtIAPG6T5kTKZtBMEQt
uCLIbZcOiGgoftOf0F4ZIaYLvlPS81c95uqmzyECPAWAz6Xe27C8S+Sbom75lBTg
zjZ7Ko7Pc6jeEwuta9IBSzwhHE4Acwt0fK6nrRAJ6msqm2BdV5M4RsqKqquNi7Da
vdiPtjo8tSMF4cMilDjpZDnDPjllisbq7fJe5OFTl1JZtR+EeSvF2KTZk0F36aLF
wlT8cBZskXn3sPivR9D7toJPebbo5WlY1F9naFJF8z3mPuryLAUzEz+oN3lSWst9
NJBiniHzB+QuiogVvtSNpBVzk5/yz7rO7BJckdTpUS3sh/5pNHizUjOKYuDBMYUq
C8D5vivd8w3a+zlpGezz7jhE/6abYbBRxDOqmWsveTjubM6TTgKVuFldzxDb/zrk
AsnXqqhq70XXPlDL2buJOX7ODElV/bDJSlQSwpTzsSu4EXHibWowtYHeGVATqQMJ
a9CSZslvosa5ZxMW4Qf2K6kAWZUXMOdzFX3cSjeh6m0KjMi2cjGczGXVN4xiFeGA
WhcfoHlUy/x+0u0+U4sNWrElkmgnnsQcWB7G/6j3sLYRLrvOtr5WTXdHSVcO9MzA
lJX1fuctxp9m1oGoWP9+54JJ2pg2D74Ck1+jU1ttw4F9qY8GC7O8mJltHNQ/CnP8
yIQxSfHA00VhHIGJMpljvhSgQ3AB3mAV/RT0Owcc7Jo1d2SoE1qMfw+N69J/ykow
58vbk+3Hzn2wr/JQePKckV114csluyRaeX2N4u4/LYOyj8t05T5zTxLZUFSAtlAc
Z1AuUJoilQAP9c+SD0UhMY3sSVmmSlRGkOm34S+XSqc/Mf1GF2JJpBufCp0X5kNn
wKX2pJHTk5zY5DdhSV467z8ffskg7OWDlvQjy1sX0knTXcyF0jAqzkrif2Ljmn/6
fLGgLPsq8NZXMQyHDmQBUa4aepA+Lz4aNH5asjUlxuSf6IUCV96egS02NSGg/jmf
A9qUeca6XPvf4TuKyEwbp++DyiHAhI8/PFNc6JGoCEVXFAC990t3rvrqxgyUYAn6
Y5pgXpFKF+XQZhIAhv3XlovoCgqPo3YJWq/Qiqq8pFE8UDN7PsBPqKa05mva48sz
M13owbVeY0UIlWk48WzlGXmPr2NqVNu3wt3BA1/xd0HORFOkkxg0E63yjHNqYdpZ
krtKs8GEH+5HX3BjdYtjmUu4Kp439gzfqdPrGdWkC/ruRfYKuq7rTvusd7R09V/4
sG/tol8UtNbwqWZdND80ZVkNTK9ad2NKcilUv7W6OfF/vhm0cOM1XKiMKh7BGIM9
x/In/fsi2jbYJshXF9zUUyb2U5a5kA+Ey70DdU4Baik1TtOPnxE+EfLIl4Ve3pX7
CCTnmTkihHOuxXbLzCD5txHWKMeAXYgF4fQNYHQpUBCNRxcAwA+nwwqVgdpyO+Ib
S1rdx0IfzAsz/MB0DVxfpwBeR+KQmEIqZvOOdCzdnfTkK4zw7N2YB4ticimXKMPu
4osxN/dN9vP+/uSX5AhF+QilF+52zvppGX2cygJfAzSBKUvWtrWfaA1pDWmbdJLo
dJ81ajljnVQ4BJX2LKyL6nVflddwbnw+VT44qqvDoF0x9zpRKQCDMl77obd2oaYb
/NuzN8AhwP30bHgmQ4Snxew7yonkrpnPw4YQXHGrfxkrskgKHX5YmpG3UygHaTEn
YGA452YQSfGbYUyPNr/mU11+6p+/+/vh2I8uZEEw9H1ZrU2hkBYmWb56v06rSsXd
QthaBhFdOzfukwm0f6Dp9ZtTUHce3kOiD4eCIxDSlbSxxQP7AyBIMBWEemaaTtvB
VVjgSzI+KHSk1eAuwZ2Qvqv9HBf7JhybFJLHGXXQ2Q80WRCOuKeulhJOXMNk0QND
7xqAZ+uFsxpq6TXZMx3+WAqa6FVaLYnQgRhMdgKgCBQfzRY3OTKXELyQNE/hECP7
+huZ/RBpP83J2iJP/gSNOEu1zX4xFGfutoASZV0z1jt6TqEFwApmvmzAv2qZsaFb
XnHWoItur2D0eLicTar/KFFq0TJQT4ZQWg5IQTFiMLVvWhGLdNJprjHR5yXonaP9
Q+QZ8Z3S8POGQ0+fQJ+khU9Rn3aFxmsUKkuOZNcFIynO0vh7nIHs2fp0aYnsLtQg
1A56kn/exn6ERloepRCIiSIWG9pEFO96RSwO5EY3xwiVkno0VHh9rJXwSpwX5ggs
Lm8B3UABavVaXPhpHRqYVFV3aPKgExB9X1Qf8RM6oiVuMkU5eZAMrWPNeyMXTsME
3VWqc9n999ZABXLHE3EvAObLwsdDWo62YcT81b91DEOvSIAGilvoBvS2hyGmV2rW
glG+7eufBjUS+J1d3P6+nDWSc59rTumZbKWFLKU4pxXr1EVI+3Ok+a+Y5t1m9InU
4mn2pT/hfgmWo88DuUBhxUiAUWXC5IUr5R0JVxKlB3Xjqsv/NciMABOb12a6yje5
D49CaVzOGblBvOnUp1Wqy55BGrmTOUfZm47cQ71IPHP83PLTSfzyvftOXzTzC1OC
9iigh5ASOhD3z8mHIM9lIwYJGAew2EFncjSeyBhTiikTnps5nl9AxWxSqRet23uj
81l96VYQ3gRx9c44Sdls5aRV8lGMsZ/3hqlgf4o+aSO4dgEzAztPeCQzzicvHZD7
4f4BLZIkwJ6fAsbwn2dx2TdRF8Vdp6WgWGKRIjWBU5ieYLql8lkd7d8c4NblzDq4
n1+HoRzR1HhtrUum4ULV0mHge7Hu4CwvTgjKv3znNEqE5rpBMANbgjwrB1ffgK9G
Grl6JZtmV6ZHe1/NVshWQSszykbsSFRYdbIk1jCCq8lnYG25vmMLF2Sr8FV1RfzM
mfFHmqg/T2VKdMErLXPeL71OV3IRmTqFp2nV1Yeq03qBJEaU5b2MrbpUgJK7R/+9
Wg1pTqDUWNsbHqOfHIh95MEuJdhRaJoKNOoNmeoFXE3IVSjiRfwzr5xP+Q/pfKtc
AbQCN9paPcRmBav4Hrlpb8oeydjrCIzBF1oc6/X2y/eaHil4r+j4Xqw9hPGY8zKJ
lYdf+ytp4QwtDbeMwXKkXdt8WxmpHLNMozMeyGofSN8kaWbL3RfFn0dpwYl6Okjp
SCJu0Q7ozKhJMh9o3Q07Umu+TSGvuzX8LPoWb8cl4LsjOSAPqZzTY5C8dfDxczZE
yinhV02rc3WQkO+M4i81c/MG3sKKRlL/Uj9udtVgileGUsZLBoiiz8tE75SSIrJH
4btAMxPrEYxq6ThcutkY4Ebt2omHodAOoDEXfrKcda6M7H0AI4ESS6yY8X+QCJQ9
vQ9ZK2ZioZ9SGhSMn9GMKcmSRbB85GuJ1h3q366o7ZdR+I6A6iz9h6ifCGH0jstY
VC2kN5pdjVoqe5sXGRLJ6/uChUQ99QghyTQWA6QZENAbTnoO/Iv/n4ItaMzH/Ky2
yKSm7uXeeyDbWpp+pz9/k7MLk4ncHsNbWCsjt3CIcXppQotHmND/AxAe+ZKBDMYN
ZnPCFUNUjajGGDYr+juP7wgr12MfBAfIAkpXb5r5DPvEQ9eROOUJovFfaLyQ/uxy
VyBLbQxbmZizmMr9p7xznhDAGWvDTTpzms161dQ2KWsQYetfdOwXIrJ0d8BZqyHa
Pqx9pNGGHEgS2TYBCeyo/ei89R3UV28Yk6pdl3FRvMW8oybG0hKMEZgW+Ghndp6A
8f2kP+oVe/uHWurStEsLdRG6lv8/xR39/Dt2nCDV69O47CvJUqAFcWz0W3RV4klS
nxELvi03BTNxbY8em+z7HcmYRXR0bYH30kgUWngM8hfsnf14qsfTuPMoOdDKwgaW
/sEghK1QjCkecJ8/lL+qx8IzLT2EDL9bUfgxs3QwhpXCenVYO0yvtcGneHQDghZY
7jBLDQCTupYyWzraZbxM10bDBqsfOj/jI0pYa9qz6jZewUghsKz1l1voSNXu/Fbb
EFN7tjNdt60ncqh/1r3otq3Tgadc1fD8mj529oDA9HoqN0pYVaauzWIVmAXNWcgP
NjA5Q938ST1VAlrSZYtUoC/aTDhVhPKYIIkKAwV8GiUBAnXyZhzFlqO/TNZPSPxr
Z5tsKlyygdaNThL6beTjonMetCrXZabO2oovBsQXzfGp2M7yIBMgUURws0N+n6KN
31bcBkjhswtXyi1fZhDzh8qwxYGHtT03zlQD1GvY5yVhUlUo6keTmnb8YlwE/6NK
G9ACAW5EEBR1lYelRepmw9+8S8icrU1uOnxxH+ekMWme28oim7Diu3CgSh9BN+qh
gMQ8u6CbL3pJV/bufgzlXvOD4nSnxueEZBdN3txDz5fkNFWv+GGfbWhsX+4HF4Jg
TUMUX/J2QvM2HwpGFtr/khUa2azrqhXwoupn+Hngy5X/3/AMEA6yeEwGuxuAjEaD
wpJhpiU2Cmw/IVEJIouOkhOwbJ0Ys7u6tAVGWq5Hb62brOho2xbhuJlvCd44dikE
vrlGg4wWZ+IFR29uurYTzJRBm3P6+OK9Keg3o1awZz/jv62RFvSBkhMV/mDQxDIv
zUHpIn2DCmzJYJhkyyyrFL1hG5GGx6BMcgStTPF4Zvz8r4dj8sa3OTkQhrPMtiNg
lMEjyAyhF0rpi4zfsfuRlNkeIGt7EnLgCIVeSuD/yM7wMlnnM3drxRBxUuCkExbi
U2Wj9Q8qt+0NKuGQSy/QzIKgbFHSrjtc41EVwGyZItxMTqy6vVj47r9PPtZDDWWR
Zagiee1SkQMooNrRr3azUGXA/xzmlW0kBa2wRX6SVKMoWlyKITCFIR9Qq+IwkSgL
28U9FZJvPV5WcAzsVL4nAFrgPar8o5EDNG4h6WYT9i11k22O8DQuurOFgmS+DXUm
CV/btuoIzGrIqpDqtUFdHy+F8Pj6WzRvY9VsgWIDYaz0A7TvnoXlq6YEl26DcG7I
4r7aH8HWZ2Lc8yLwD6j9WiRv2hr6PIwyEVI3qfs/fBc0qfKtUDnAV20g1zlP0F7g
BXIC2SrI7D4FDdTVwDzJGdV/lEi/FCoQ0xx5kpITQSBnCjRYul4TlEfjF42R9zBH
sIWj/S/hNs8ounZ6Lp0ImHC7YYClJ3ygaVoTKcJCJtwEzksBaXLNGijHp4GyUiKP
8Db2Nh8u9JOxbPV4T/7i14c012uXxHRE0EVRLtaY/Vgrqiy0BjfVqWvunPNUyJ4l
LNi5FODmfzl46urZGC6pnVOe4NbknX9F9Ro2W1x2kZu6cgVKKaVW3lodJZoOTZNQ
anfQv9LBWImO2WL2YmhLv8qRCUcPPtSMrh+gJmO9V/nlzs2ZCskFjHheAYrxL3ab
jK3ZqpK8GueEtLhSZNb40GFS98uNxxFE9hAM3OCHwVCK4cCm8j4GshjwMa6h+Qf2
cRcP2v0J7u/Jadzl6qkutjlGK7Nxbfv+Y9D4ui7S3MrFwDLjZAZfcBDhLoRa0jBX
k7GEX8Swz2lD9kB43ntfcCqJB55rbAK68YibMF8NQICaZv5yMEvk4ZN9IsDZ+fdf
T1sedOUqtTi8LC4tM/LaMAB4o6B61MekQEozB+B4pjng4sExJRIKH6DYKzQ9uthP
XTjtFtAYabOOfyR5ljqDKff+ArdCOEYYt66q1coHo12sJebZazAEiVfTcxJNxZHI
qE8OQgmjCZCfJ/Z/9R30GuJ2nwcdBXYRlu4tH9LVHgb0YO9QdImatj7RMIce4t3w
IWDkFWtS2N7cOzji2pPL4Sqwn9CCFsvFSxqDd7y/fYi8BjT3h0w7eWlSxwUeIJ72
Ip8+mXyKRsxeYDNSHbrKiAhESvrSDZLtFEAUT+jVVtbZB3kISDEEzpKpsOs86Sl0
2KOuMMshNmqZwTwrvqbNAL9aFWDcxdLIHLxs8QYtX3yKIOH2G2F5Ou6Jh1EhLUUG
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5040 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
cjljSPzTIRTXBX/bLgom+RIFjdQJd/2FHfhoA9Q1lX7a7CzERytx4ITLyrDXwA90
7TIRiVClEbDkKxOtNzDVzqkrLkaaZu/LWaC3C9LWBu44teU7NqD1T2vdzG0/im9x
j8tq9znQSNV24NqE4zyu1LezZDnbDtSTQpT6KqE82mv1MicRZMvbuoOEyyav1L5P
t77grmp62aWYLeWtQrwNSPFnLwPFgYcHp5MyDUJQGCmjy6+hF8C7DgbzLF9mO8Dy
v3y/fI6nsDBp14epcVHjMA2QFUD2V++tbNXJBYltrfZwpddoYZs63JwCLsoF/IDC
i+Fqt/jRz3sm0Mse3JItCFuVKYg4qhVFk/h5V8dsXxnSpxaP39VE7JVVrJK58vBZ
XBBXUVzAH1Swz4aIzSLkBhbeErDKwGDrN3YfEKTM7xw354bd6qy0fG4eTYhRC7AM
S0n1bXVV5mhUATUqtJWHJO8vA7C2PP5T8DRCwumBY8vhuExY1sJAXZWFZ8fXevYL
c1mk8l7a8fvp2+oBTRTytTDqmGC+/iwChAOItFygtgD/EI+ni3vYWDbh4j05Endh
1Un17ZBcNit6pZ1zmOPMPcI37GzXL9/ImwHoUALtBMyVWe7sJqaJ5LPk4RX1B+zP
p4NdzDNS1Gz1vBVpTXACPItzTameSsZS+WWnONaPaXe8oZ0ZR0/Hed9lYKrqTaqT
l5Ys7+BC2GMiIK3oaSRYr0AXf+HUWHuCCovB7ewCSkZER5HsphXdT+NRypuFiyqU
WCOyVb0ChVscQ+ecS4qBk7ApF3/VoyBzXnuGgz2YjU/xm1K1DjzTKRepEAOjoelo
mFyuK4A718Uwm9hesnewR34Q58lTc++5CoOubc0Pozb6jusH2uYlHN6W/pf/Cgmi
48zwS+auEXBCUNv59gIxlBnD0ffUt/mVqfkVCk9rovGctKFa8O0CMZOTPX0svZZP
vr4fgxjD79sgUr12Yzcp8VkiQBugzUHuUX5HMlqhNmA2+dyFak7p+W74/PW1WjXF
Id88dCO/qimT97T7qE0O1r5PyLLs329YdaBE2FxiwgvTDf0pITTnnudHsF7gn5Aw
JmB+MVLO7cJLdvW3G/VIwer88848MuHtPzBS0YPsLFBYbpbV48KJMHkbJcSSdoq4
PXJ1ZjfH78daAtxwT7Cg0n8KMs1YU2Lc5eZonvuOlbje66vmKQhKCu0BWa9lOwWX
DaIE0rvR7N3OTxP2mu90HTEXAz4fWQGNhp8cqz/iUUVoeqKkKWhSWupPSHt9bDNv
oKQ00QQXynRn5kIoEYPmVEPUtRG6xdW4fyHB+/qS+BE4IZpYnS7jArRrQuM5RkSD
cY6JTBT3SFNxOuEcwS6cDGntBtHNK6C4Pw/a3lh0ZvqSHXDuW2hZ8x++HmuzTHfe
fKPkSswPc/J9UppRkkr+iRvYLRkIB46oxmxF8CtR/4WuzmPsohSjFqmF5YizXSLQ
xdgXdGUAoUo/+E5CAgQ1fTV4nkHE4XfKmuVtkDMYHhUoCAl9b6QsQlfdXHdWAk5Z
2dOKNzFS16utclzz+0aSIwCDst2EwmFfRqV6JlzBbUoOnguiZO/H582FLkwNZWkT
qV3XEmcUbkeiRvAHG6GN4HZuzYOed01kC49DeWuFXSXFFHnuDKBQvkcdWd6SoYOd
qZNb8azfFKctNwzXy3Ajp1nOm+K99PTmfkotRi26BrYtC3eDVh0UFdJjvf7ouqt0
7GnhDIJsBGE82s6X+C7S7ItHpolNoXeCXzVy+sJaDkPb68ZHPpiXXAs1P/5wErt2
jTxt+EqxCWW2sK0tka+qAMheVhXBy2Bs4VT/hDV6AfOno8PUBBNj2sCme9cb2YMc
HhXZCTnsv2PbUJr4a4N2RpnHQBEGCxQRdl2/RYFkHw44kt1FtBYz5NLiMqeiWKjU
V4XvsNR4nFQq/4j1O+bnMTOj+eULYKPXYDJSMSrrS7rIkE7I0tptqI3+T6YykvR+
aubkaBO4Zv08aj8d/mLdvcuTZetD9ORj8EkJVSeeF1LoyTeIeR4K0ujEPvwBSJyB
qngacJNP3FY1QsZFgR8624RlY3qa5ts/cqRxDsK73Pt+N0yWrdTgfWK5Ie7ygLzz
Z3ODLsbnZ77uSDC3NdiO61WQDAS72RxwA/iKrqGMMgMXIxLsQx2QJHXrsoe8DgqN
pPqhPlrQegL3BfjQaWuYaUnetw14qdGGpAcY1rEYf/Gv3ATjEK0X5PNilIUhPD2O
Q0Kj52EhduiQYc+oNJwo908Mq5AM3SbtSJzQLtVWQ+7ISqsCsbN2Pl/FO+EwLGxP
KXBhYvqeu1peBE0sU23jZsOugIQ/pgEntQK5SNuugVWpHdXz1VZwOma2koe9qLPV
NZIPP/5jo/6tftlVGVjHkS2yS7Y/doa5nxg46XWDJ80fFUqPnZWY2nQ0ISfWYKYc
4ZWJXWKePgwbiGHMILgz7Z8FsOfvQEMVgPL9dekC7plqLrCzhOaPbIinAZJbS0lY
VtCtuvY6KkIPeN1w8L+8gGRGBuKy4YSHeqm7YAlM8yy7sPVUCADDn+qWhOYlL060
LsbXOmMHKrFkeIbXnxE0fmsXDrj/gYzu3IKkDCx+E6PmN1Oa0OK67JkP1s8Rd0y9
xW6SUiLfBti73a1Yhpu/k61/DC4LT9Za88x1cjsoUBhrLgrHav8j0eojl4oXy3Ss
nQy9SsGKCBJdVJaQD9IFtYX7qB0q70NEs221PcTBahjtwWA/MJ8g/ZVLB4Pdwx3k
EnTkiXOK3aIPr3olZIJON9X21hItVaPva7quT954rmjf2QQTTOZyKh1eYiWw0lrW
adf97fMpqYDcCl95ki2Gu6prU3ZsW7l4fxvCffg7kngrWMTxjLK/pk7n2a2hnoq3
5chy8i7UnID0dOOmGn38NBzidLbtbtC22iDISTyjDIHZXGxs9GVbQSzfdf1b2zTd
QW2kdcGX7QLblaO01PGXREvnDXumIfguEFVgKj+6HDEobTRosyvOBHPKuXy22MD8
4lxs/DeawVhBUxyhoDi2R8uT9OPPGjiBz9/ekpLHZpKiKMXVwuy4Wl8pxOX4r9cL
5A2nc/CUungZZ9GrmVjoLBEjfiMcxdV24cvBjhBhBCZ7i6nDx7i/53qbr7sX1w9R
DiQQSVKTTskmumeOaRIl5VPFRZLbEsA7SGr6euC+ZFT4qxahiBKpvf4YAkUC5Jdh
jjGgVpIP83SXir29Rj3Ii6xwPwJ0FqJDUJnuT7x+j/wwifW+PT+67rafEduDS3MJ
1Te7uKPG/hhPoKBcrcAhAYsjeecTTWVkYi9i1ucKg6Hi9E2qfBmV4SHt8Qqtyhkc
dC8HwjBxtXpvAIvGEI0+1QjwOxgmts1hI6jZ72UKFWaqeHtDZYvQbHRnmVZ9oZvA
KDLLkT3F05BZe8rLenMaLPIkMXknyLuukUtMcpOXMSI74dkvc1w/lrd8hrem2End
oxaDLBAO9pNBiDyyU9VwAap1B6MZ7TWDphQEWD5GFUBtjHKLP/1QogtUY94r2gTL
ZxTJoEX/Tld5xGpwE/83VvI3E9VrcuZ1qohuIsM6BfkH9G6kfqRHvQTVgbDhiOr+
JIf5xhBhNwwyT8QhcNpZp5hJkk+VEMirjSttIDLR1m3s4N9uxhl6xId356bRaXpc
n7D3FWj4REQY+OulW2G4L1d3nb3JfFifiPfOU7Vxj4vHKA2AUQKBZEYSB1etNwDh
8Dma2ZluCxhn1mXZ8pLMF4od7BOIQE6miKR1XkxKVwNgmlZzQ9aac6WsNWxu00P6
lqfsH9RWSXqJ02aXnShSTYluezrnMrn25/Qn7Ns0tvq8EYm0zqlevBTigUVVxnFM
LsAjL2TxRzb1ZzgTyU7G42vC8rowAITc16oCa5Oi4QF2anuG4dJ4RTrAU80GTcaf
UwpTV6j2aYs1G6Mz6fHub+U81W7xbBUvlfu0TpF/f34MihpSd/qMIpguCa3cmxlV
pf+dRZs/IIftz/wfflp6r9njb9UHx7WHPM9MUfOD5YW0irSpTQbFrZV13OViMc+b
SUHPYc8vRknTAC0Czlhg1rCs+ELqd/LB3rA/WipDzNeXtxrhV3mjoN5pbCUHD3x2
gk8GRVlYq/kljyotzAhHPA75KZ7BIa3Cq2Av551NSzyHtQCW4pTyrSqu5FaQjyQb
HYmRtQhzx/Vyoh1+DMj/axmNqWCws84ohJyc9XkE0n7pU2PIguSHvIascvLDV5z2
eICBv+wjXDM+9V3oRLBQ0PRxhn4fKIyP1SwOYVa3O/tFklmRizUPf5hgzb0m37Yl
hvWNtEtMwMBmdRemxAiFpIa0NG0qsbjKx3Rt2o0s5umn3CfiDA2lA/2GJfwrS0lj
z6CIvXp/dXgux4Po1gbVNHkZ7XwqgDHMCynNyezQRVLwb5jx5wBt50K2aYw8N/Mm
GL0ad4bXt3xa2XzsJNNPWoAx/h4XXsnd1nQe7W0LhmzD2k1/MUhINAYTe+o74gm8
VDPi7RbWgGt+LTJE16gcl4nhTTZrypXzG4pqR/spycWUT6LK0uTebI8W7635b8uC
qjmuaFsxCx1fGAlEPZLfLOvq0vw0mOEDvCw1tzBvw63J2OiOheP6hbO7G7xnC/B9
CzVYdxWuIYObbg2LhHEKV9RH3CQeN7rakSR6+qukUbc4qfICpBGqp2Cd3LVNlH96
vvCU3vyo1RzkxVbs6gdbAYD8Fzf1yY002QkzvNwYOWyCFW1rBfZFrLIGRsX2HXkm
NrqRDpZeG2PEH8y7zROmiGB/Gd8BwaHnc/p2sXOLVgu7OGzBJ/QZDOPIGpjd1XOG
xiYfOR5961H7SjWtPKdEH+9gpU16GAPI1DD5AUiFOBWgcevVBPuqEjviPzAS+lTZ
B0c81hWsSq+NMyRNhY5Y5UJLxlrBbf408zx8PAXWeNhGQCChGyXmrxQcZyf2OO43
eL1FO3WWkJsIIujw7Nr1nmTPJvZDlHEqvjcFqUQN/NQM+8FHqQkuVJ1aLpLCX0NE
7Uz7F61yYSsVYjacCApy2oI+JdNsAjU2VXirgEBGZzAehORExugu+aNGDWgqIaQi
gKkD9XoZPhUUOr9f3BYWdKrEs7YziNYO6b/NWwZfVdPBAkF1bgH/IQo1d10KmTWO
MjgXN/AyNgP5y/FGNyoMIs9SPLBjK46P/pKiZbJLnQ1L+3BhayKFpLHgqYFUkNpo
Dh9ZnyoNl0EKrUcTdPrd9tk7P9yruFJ8MWYdAOtg7nrWb1njLr2RoBHIVXQCxclM
Ngs+mu6wxxbIwA9N/mMF3gSMVSbAJgmVd7tPzVhCv0CymxBsg0ogwzHC4mqf/6JA
sU7mdXeXpJDMldOv8M2QU2g/lSliyy+VYH5Rus5a1eZ03W/h2LFyqQoAPaNVG1KT
gHldRrPGx+5I3luuwUzMajFdH2PBITvJvN5AaineURCVgKLBEs7iizBJRpJiXh17
EVFFzFdBvFIkIT2hrXTFco4neHUw3e5Fb9NvcRG/tvpSGqYTJQgVzOqsGJl0I4d3
VRL1H8SFrgyTvMm2VAew2oN51vyGq3NyCKvg4HG67ueGXJpHJUgzn6ukekTNybAS
GkCHO2m5Y5H1WsNVkWLpmtutXpKsOTrCozUhm0qI6zFf2K82Odb223yXYqJzrBCg
vCL3C9TwkJPdEjPUhfSN2RV/LeXf0MO/AHaLDcjYiWRmG8ELVJ89rhyfKAjl9/r/
Px18b14A7pkXu5RaUH8l25IsWIIrmd5kIcbq2Zq9MGoIQAXwjdOAMJwT1RtlN+Ds
MmZBnnwD/tCSqUQ3cpBhj0cKE/dGdrf5Ex5ytRfVCospcU2Oimcu2pV4ODZKRNuM
GduSEqCSf4+DMzGFvndaJehDLkqWPbMwcXZPpOsoJHBybCNo0R5DmEjgMqFZEAfF
R6kKlsPQrdw/vxLgRfyfTboa1mfOL6MZOh6Apr8KJvkOuTTuyv4C4m42Q7nTftc7
ks8bXk+8asN9TPm3gvWtCdzifNBzdef27qw1YyvxJh9kIFnkXOr/uHskczOJmF6D
jgWl1kKsO75KKoPEiq0MpkwMypsRxOczrInlOFe1joAYNjYiUJEXXAA1fUPAZRuc
EsfcXAIBBh7nYRNSKgPRR16/ho6/Hb4v/uobyV7snEzUTZK1RJtKxAP2bU9xXceP
mZDCNpsXMpBYPKVp3JB/vnNhbmjL+zxkPUVtzMibp291hSem3n6Bn2gTeQs0Ia/q
SaPtSjsTkQJotdlhlDOo/YHWNbG0gpCUOvfWVCe3BE7mZSWTAy+a+oRkB5PcYASr
IRbwVOFIwix6QD0yllgRBuK5OpzSvsNZEl0jTKxRLts6yA6clPQcMDOoi2Oh/S85
CNCKhrxcJGizWduS/FzCa5rTST+d+fT5KoPLYk1Iq+dhwoQvTmg/x5UC5LVLbLI5
hq7hB+KYoM7EvEc8qGsrsyw7GVFcezId4QFJ0TwTgDbSca7xV7aWImtloYHIYZoT
B8h4Xj+QR9KgVnqGOWbDt3l/EfxZapxVd/Cf0c/WSNbOQmUnFOrI7raE3cG4KycB
1QGoFzeLe2cSJsm0tP+zHcqbryYTEQbHnUqGZsZ/xrM1SX0S950snstclZZ5bD0c
>>>>>>> main
`protect end_protected