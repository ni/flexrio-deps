`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
HDP29p0vLOrNPcWDOvry+U8EB6hQYaORb9dfjuAHZl9qtYswzrIuG90EBhKLEuIl
q4d7b+5gmCYrneF4hmQArJUEmRK01CebP0K9o+kw8cAvsSU57v/hsUxCmp5VgcN+
waaLbn2XHyj8ne+lCTxeL+YoLU8WJpNow7u2AeEZrtFOyx4LBJAHjCzfeXCxME7u
DDA4zd6imL/II81E3iclL1lPF2LNAy5O7uGU4AMFOVwUNVnIb45vD/9lglrBHBGb
+qP6ReXoyZBpfd3f++WPc5g7UG3UDxnvowSw8PzqG5C8LaiH1GXayKXoUbPvbeOZ
5Jn7AHyusLwCciPe7kgZduGppHOGmbrP3UUqR4M/nOKHY6UgVrS5sS7C2uzxbLVe
sl9+qMtTkYOLgpycRADYpK49z6p8Uz9woNYvf9agacDMp+NZuuM6gZbsh3V5Hgyy
tlOug5Lwhi1TAm6X8btco7eO4topFFEPapPRV/vWcXd14DeyrYR96buYfLKCKosa
Hj1UHs7W28SM06xl1eewEVmHoGpf6xHuIuWsZHDsVv0xrYu/jCx3rrMv7D7lrkMW
q6Bx3ZbfxPZtaT3ShW4nYhYdmb74ZOPYAeX1QKad+2/OnQrRD4y1JubcYZVLaX+A
XxqjNnFTPB42UpfgLEJ6c5VJY1VUZGFj6kPw2Jo4e3ePg5hb32TutqTJxb58+ida
mMki4XScozokLUw8cglXc4bfIqrCBEdGXcagSJcusoagqI7CJC2ONbr4jSZurT0T
ZAJOiX84xZvScIvN54ERI1C17DK3CuLJywMWzqtc5ejvl1p2aFeNlVXl+6byucSq
VCB1MB9Z4Tlp6TTe8NuHpq+unFXuerIRdZC507A8F3bzk6qnBW8ksd+BYKlSD1Xj
odTxNwmbcTDujeLzbav7P7+/51jV8pv7E5jmQ5e+fNTVyRKdpcZYdZlnpjtLSQAL
JcD9pKT31hSV4AHtoAYF90o/U8eU9WonHf7C6v9xvvXHADGBihhscBHspdW+Xu6h
0WmcXMoP24lMSFyouxVFrbUGZIYZkQezVlDXW1NW8UtuER3RIKUY7Vp6IXxbg7RB
h575FWMZ8kvij+lLjzeV+h8tOT5JF4hjNyg/oD+ylQTsID5DqCF2jrituo0shAZ8
PVNpRbWvgtNFsovQDcR6jZVKYWF7u4/rqFERMJVFlt2qFbVnPeyM+rRJDimG2/Xx
IGGIQeRh4LSaJsBJWAg9kqjIMg6XoAZlAv9XmwLIxuRKPJuzotbzLO0viS+B9ub+
vWEqVVQd6XCpUw+aDOTLZJCBmt6kbV2g/fK4cycrWS1FjY5cKQJtE753B3E064VX
R0/J+QXsamF98rUxc4fa+6C91JHw0KJALc/vBsdg57dPPLFyIdG97SX8N4wqW0l1
NKxV5H9EENQXh2Oq4rXj6j2vRCUWChJMU4es3s9jdCJYNqn+vMBT77kgjCJosPEs
6ehYDymVxgztldu6KkGwm/Iavt53rmEkofWh7jW6SOB3dDgliLTTrimG/Lfy9R3t
EolFo+IGmAKWLiaxB+f90prIJWkN8C7QyLMgTNNHPxnYd1mmdCVqP5OQIiZSVYQN
0/9Bb0Bvlg6lZmOp49uVoHUZEdbGpel8JgPKkuvpBXRbCrNmQxznG/Lm+EUW8fsL
flRq7U0SiNkPPxctgLVG3Nsak9bIUbVTgHhUgWFnFe4GVwNS7GOql45+KNcLMzBa
WmlBLkEcBlXsDL2hmT/OgVAw0p1pmKbWS32EZMh1R2rPLqxwYbb9eTv6QZuMpBrP
U01vfYcfdAJF8BSs8z4EmbE0WGBktJ1nf7V/R12Mjfd+94seqGMrb9v8ghoC+O02
VCPBsAlXJYUQRYKa2p36X9MWDIARjCHUrqap07lfKkxs16bZRiBw7bKKFq5Cztwk
IOA51hu7ZKJ0+6POQY2Z+rLWWlYxaquSiH5qUL2jbHwmULgq4RAFfs3+pxVgQydB
VK29Fs2ImK9JsOcRv8vszYoF1COk6+FUk5NtHTH6eZ4T0snEtP0OlJ2EdTf3p/+n
a24jpLqbrf1RbY8riMo/iDSMGthVG13RFcvziQHx9HNvGCaeItxwPmjLtPOUaGiR
5t4oRlTKhJD3tv+KxSSbg4scI64HiGZRTCKNYD47lQXTHaUSPMiyDms8eHPqN5/R
BeHoe2mJrrYnOBE9m3PIa7zBubC3gbec3XIdKE0qgjutboznzLn87J2Ua3gCToK7
glHyMbxGFCc3O0mUqU7xL6h1tx2TlG9GUJRItNVyqSLDSeOL/wi8JgWs0WfRarMf
J5oH/DgScW1zSAoChfsNvMP9pJ66lgbFaJ+Xyog0eQAOFTt+z6T0xhGsQg1f0bbe
rKIRYqscLJoLW5vjbcpEH80T/NENkgNbPDFnkerXEU7wiOsOh+GUF5Clb4ulZOG5
EesbqA1yWo+PrDhfCPmpytXEQOn0BFQ06BDyQ5dPt9bf4yMrmH+3UNwPmHQbP6rh
D4EvjKRsojew7D1QpWMzYkkw86zKSYKZW37pThOipkkCblj636RU0caraDesISLu
GpZKqirOKVf9kxkmczNgzyE0FcSSgODEHGgk4glWc0PFqPBI28oQm7YOpSekwyMs
3QF4zwBsFNwYc5U1wY53jn8AoTuJGlhnIg+r6g/c4I2YdcaGV9flMBbbHNIHYANp
qqIp85ZvErjsjBhiItp9Y+X14tE0bMHlNDufPJkN3RjgNzKlH9ZbiRA3gBoM9Fij
IKFTOz1RWvuQHnQCr0iAePSYxsdZPtV5iZ7cPqDwDozn9eAQdnanE7FXeXp/P+Hs
HkneVdlyU+RLDHEfGwDrIIB6brZbCf/0k9VvvTujkT6bZVxyASScb51k1ZwsIuw4
qFBCgPgO8Ni5ySJHG+sEsWR8smMsWShB8GwDgm1uNED0A8Y+JVDSg4YHGs5Z2V2w
ajZcxO/BRhiMr7lDzdUJ2xbB8pqASB6LFsMOPC31XiZft3tcjID+Pm6Wqte1hEKW
TcDxUc09e6pkcApGpRGofbZhnpSkJGL1upNq9TrJ9hJX2tSu+I83SAGIBR+UaVwG
7FRecn0Dqwl6Fa8nfIgoP9UoutUrUBnwrpIjBbj63D159taB+5b8lJ0rRYLsFxHI
s2uvOantuoFyp4O4q1dDWFWtIjiJLulrcPPenN2HE/sT/hPTnemDmBU1oKcJeE7o
3/hK43p4oLu7WtRr+HMnTtlkyPPRBikpLqh5XfXevNU7KOgqLksIhPvKD8UqtlF3
6nf0J7yTFnDjgITf6Ef1tZXafvvH+nc+07dCUtqz5ZnVcaGHRrV3h1mcvW3Gl2+k
S7OS/BvYZbvdx7nWS8r2JH8fbO8THmFPoit5+AsD5cw2F73NSxUlonn3EHQQxDpB
PqN3JOWO8VVeuPPjaNqaFzECeZrJrC6JJjaJH5KfVSd/TbBOJlu2YBvIyt1iOkYV
WcA12zhWEiTkpELGann+GY4mPpd2uzGH/K221pXSMDQkn9EvRAxxIjaa72A7llLi
6Ms7w3e/ppqFjUGOUKzJeMwmBqUn4M4hw1fBYl/k1s8QGhE4pl6H8eBZswLQVCf/
zw5MMwKr5gtKcw04rqjd6bS8sAMb/sJK5pdS9bc7xFarzRNvzJrTPALB7uHyKcDB
fcR7tPYMf4TfSgoPyV33zU3dZvHU5AKAoYtSlxa8xoK/UAvz2ODyd8wXsdJtqFjX
u02CRUABkmWBtwvh+wPyvB/VZAtnaUJ/W25tG57BMMtxSevJSDH6uhBqOXUv1YV8
uQ/NnxWAt8GlzHbDGfDH/kGu0tEohZkYzdDOl9PZDLJiiJ8K7vi+B0XJe8YMuv8j
wfQSRvGTFqDM0Pe0oxXRDU5m+TrNeP1V8E9WPhUI7y1UD/bzHIAAm0onjZy1ZZlt
y610JcMsyw8OAchX5B2uivDTcnnS4kdoYRP+gnqoTRb1ahXm+sTFwrEn8o574g38
Z/d0vO5dxy5rOuKR64pUwjrBq3bquK50qcDFKtlhQzu6CR3vWN2pbAQ6lckIE/VB
LeSFR6z3r0didBw2j+JXojMl2COdQDSbzftWPk7WIYm35x2ErNt95amX1LQmtisj
a2V00XjGxcy7F8p7Wg23R55thSAerM5bVktbSiMeOmBT1ycEy4hVNbxULRgpjXr+
0PbWG5jQDlAWdshDR5aw88i+dL7nnqtXx2Jsle5jk5SXkH3Kdk35xVTNX8/P7rvN
HkJXjyowy4sXdLsOfGnnQ4WN1FCbHRqMPBCuGfChgmog5CYYesBMmEdUWzK9UQr8
uFusftCQUTTPP20XO1nMVqinF1HTPR/SAr0SPcC3WzungU1o0nJeMeCAJT3tHFRa
AYxiQhEyyt/L3qgBu1wXU1U+gCdJdTd81rDR1tRhLBYq98oyj88cPyRr0YJb2+D7
otDfLQxuFiEwQAcsvNBz5S493ADa9biaNCJwNXLCYNetvMCb+UsrnSN9EaC7/Dzz
MKTmeUWN0h0yqc7CUWeaS4zSGPWaEVivcFPoXri8TIF88B4IMu9b5YVwUtjWxcVx
XZcj/hILOr7zIqVi6O4SS5hDLjoyyzUwu77pUykFq2zgrjMWsv7HQAdtUGVioXBT
5WgJdchWrcwNxlgF9rXcRn3cgauyUMbG4lC97M2TYaiyByWDGQLg/r6crILoddrq
f7ZLaEDimlKs/sEaXjW2W9glm/folapds3Eo3TjRyey25vGU5b/RJZ+Ij+4gLgDR
aYfjnjW9oLmqZFS04j2WUc5U6ev3MqfE90uLZQxyMWcqyK4bbApOqdj/T1TNl+UF
d8ahn9OJ/5P4s76mT0mRLwSfnOK3dKmemPM2Dh+wl3LLktrw1hAiHaYnTbWgbij3
Y3cRV9rQW7He6swWoVZMdWTAhQkn2FSb0AHk0xcAztnDDTe0WvAxw2rVUd5YONd5
rnuU3SWt/dE+1V3q32JeAioVe+yCPErI/N1f8o7VUzBDddRa71tGM38F29CSWPSA
/x6eIVnu82+sKFc3TxLwjbzkFYpv/7GYw0sAiRm9QVgrW7dJXL+a2aGVocOzFAS+
SHARAGQCz9D65VpdMh3bZBdjHgjZFkPc8QnQzdiFYfKGU9BoBt8PouZL6pge0yPp
3raXUSiBoVAxvhHN33AHdoCQOHXDayuITeISRX6tCjr/RNF1VFu+YEP0QfhlsOKG
p3i0UAOkKCB+uWERsqxJhYLofo9cf58hcZ/dsEEZFatBnhFLnNmSj2bo06esLOvT
zJ9YVcuiRob7igCW7rfAtADm0cc1gMktAvUaa6gySU3P8fCiwe8Wsf4zw12PenMk
+KxmZg1fXC9Bq1n1UFYT+f8iY3Cqm6Zne16mQNoMUNX3WoIXLzFdHqlKLJ1YRrcr
x2ve1sVEGGYSyVifntxp3kIisdhEpr/wgPwgko6kePFS8yxuhrccuJ78Uwg/sG8Q
ZH/o0lQPZinUPSRyTlC+2SROV++hjF5Ny1YduEyvHvyV7eanH6Xmnj1gbs45bXL+
qU/If/qpWuQA9V73dqTfPBcNGYB5qQLGJoqKquyKaYU7g8k+XSjeAHFjmdqOtwAX
4+fE63rtfP2QVS7q7AtAFiav0WJZlOPdxkszkqYJzTn5Qaf7A6cZ88p7eH/ZcZ5+
XPY46hTeReg/SkZIoF7OHyUDpIpnbt9A4N21hme/wqzmCUbsS9on5bPWYdfqZ9Rr
e5Jx7lgJKJiUfs6AqBvwX/HoOe7K+/WwDRu4Eh3X7/v8+Uzm6z7nuTrDPk93oLmd
gJxZXE/hWGnVu4Yr7X5oxcAQjxhqXldIRxq6j4Y4JAxUf6Qy1M8g6fha1Kqz+QIJ
zJxatZY8UDTSROXm7849BMMtvSHd/EPqA7+5ch/WDahy+khE/RPvGOe8I7PP7xVN
grxYvvfFh5lNS/lhwcYO17IXxULwPhVm7aUscG79e+YdrHVoJc39tqLutum4s2pB
aXj6XbwhYUdpNcwBOfyZhH+Ubqu3bAfPLIFW6VskI3+20zKwcfED81ZEbr6w+2/I
anzB5HBdG410hQ2VTXXj3NsejV85tu/iPB1GY/Xkm9CuiXMbbxT+fDiT4Ngt85IV
SzZIeEztlNgDkzXMyFB3hTvcqVH5kH2qH2sa1PHPUJIEz/dfEPsEDYzdSuxi7g7N
teaK4mYcSuA3XZa7V3+Ltrh1VU4bM2EMoEOkPiiiPstcg8kG86cr2HE/OkzKzIjd
LNGKJ81kTuVfIXuLMlFv+NVQbsFZhENjmrl2r2oURod7LOH4h7pk/dI3Lvc5SArs
AX4SSSqeaaoZJ59sTjqBcL887P3lUKzdcDk6oT4LBmEGEoTUuo8S44RM6WiR22kB
YrPdzIsBMEUKq3qRPG9xbC1zfMd/AgZxiJ4hCXol/A0NxjKSJJFEO1222vWMB9tg
Lc5DdQTZGRaGCJC+diCVIGRDnx4kXI/wmTRMdeRvGb7edWC+QrMcHFR5WLlZAnmu
A+qT/WVqjkx93eT1ohN2y3/c2lyqT/m8J/DZE4T1cJJvMZXkryo8O6uQ6yqtL+3d
TlnlBo5iBLg2c/KQl9gyaD1Z1Q+kB2sibZkOZmdGKYFxI14AOG6fucTJ8z+p3JMb
0xfmubbXCRKiLXbb9p3T041Z4DRO33FOGf9BUUk+NWFCQaWnxvKw83bOl7JhXm7F
gHcoL7IM3xT/tHVBPiJzg9wWPolPjsDbauD2YMukZjku6/1b04qTkJGlUws2YrpB
Fcql4+LY99cNQ+13IfqJq3+oG8ZOW2yZsafK7mc6p4hbzX4wruaUW3asKQRvjB1z
3zRisermA0Kq/WN/61TIlvAPmnMrZjgy4PPuVDCvPjYxlJeTuu9+YYSOQYh/A/9j
EgpSXBKzMMiJM5fbyw91GCnfZs0zHgYxHHTVH/8PczD6PoA3BimP5KYm9sS66agv
8UBV83G7tFt+VXkOcqjcRJ+9N2E4Ia2J9lT18qJi3OlSDCxVbmgtRCF+ok063ty7
uE+JvNR5UMcHtaLu3t/wXqcOSPS8LRoZIpUHUfgKvobeg9ak9gN5PHVcwbiUFguS
WAL/9K2hDFcYXWb6sLgS8u5r2LVyuJugETX6trIVtC4y43cYsGIgtb4GV9c/LcjG
fVmHCt+K9/EGQRtjWUppxMA+d5j1n+4Y3RazV/abPiHkpfVL4VeS8mpTEelE/ODd
HcaBShYvzqGuQsmgg/d4lL2JGGpwHq83PWESfCniHkALvsVrXivMH7/ko3nC9eKv
9XHLb3UaXV+zyixweU7bDvFzwf2ykZns6vxRLpmik/dA3j986R2ZHljFClaRJaHH
g1M5mKsHXWtrhfQk3fMo3pOejX3GXYhksREr7PpWcAG8sNN5Cmf6npJ6qCIQrrEh
lwmcB4s6OlRYbUGEk8u5zEmZhI34oI1OwWxD16WP4rM8pDkp6GdaijR2g2LB70W9
acBFU+1rV3EzlTfFdyBJ/u0Mj331YjiLlBuleIoZ/9fI+SAUqOR6saQ6zgvMAiyU
6Tv15J18mhgB5OO+x83AhnsubKRIzNZ1kEDwDGwQGqJsE+dQirVGJ4rqEsuMqX8N
z3F/eQGxgjr5Rc5eHgJSJRmgOle6DD7SzGfo/KaW6TJ4AHYAeB09/1fuqUTH0B71
A1eNGhqgtc/uVQGvXW2G7Uhvu8JLxixVXu33BMffYd7yMaAd5Ov50KfWSyjU7DLy
iEocacf/URc3N1iywKQjTkMl59tDfJYr/EOMKWtJb1bUPJu/aeB2fJ9RB84jtayW
dWQTgZMcLxwOwfKlZhcrhswL4KEWSz425KpcI2zf2SMIyWSuw14/+3aHAs1XkbTA
a4vzaulyuF8Qm9SmFAyA9M9F0rd/5Sq+AYIjcYq99zq2ZwtF01ZdZxhHhCQmeIC+
K7Y5DO4w3B16+SIQPeLb6Jxgx91L/GIEREcG8FhJw0Rge5LOmi0q+AMnXXG2/cRr
gFYRb36jn3B/zOkqeztFga64epUmRfsyrtXfaXW/1ef3KBqtn5FGBd4ciFAMIWSr
2Fu+Y1XyCMLvlBWLqNye/mRakS7/kvkrZQ6IykQ/aDaYABPs1cwgHxclM9oQdEAw
X9SZx9ulxxbPPfq1qqnutgGQbf1M7kWpmjpRhCZ0O9CRxINzpCUKnmtBhES2EQNP
lm7l3SGgHHQR8DiLvQoyxrHNU4hKvI+tz4KO5LvErleXjR8jotDTbaqtnPuCLoiZ
94hj7ZomSdtzaDReFeymsPw1BIQH+YFmEY1t+kNjl2tkBhjwbMV3yT4+wWiT98Uu
0S4qDLXZeXV88NVWbqw7JjRE4eMxBo2N9YArJbNzr0QP9FTjtMCKaO2Z8znCQEq1
yz9XGhbP//PwPeeJV3E62wFXreUF9QEuf+lQOU3xflemkjpi+3N0GdgltgHX9hBp
05abf2Y7YwNr/yPXgzBfBKQFIgGcNW8EFoXZUOLfuVSquYj9FsvardwVBr1hpNZg
nI/gqb0VXqTxud+E6dQCnnBg9Ul/jBqTfiHm9yTd6lyOTINwVqOa8IOpOpQm1DAu
MIKxdl9U9hSq7hM6vHfbDEGl2wJSPOp1YE8zRmiUJQm+DEtmz7GLYVixPseTQeQQ
rDgtZR7fcLfKqF0L8BzSZngjDS+CwED406XnkDGEX+hZgFmRnXJr63GJZCWHyYTE
fzLEvLmtKOHPzENrJi2lG6pI9qgkbt4GpT+PREiNb6JO45ao/ubslAxERvwI8HjV
Qv1IPgennnN5MQcIoIHKCTAhog0uEPikaISfxOuiesawc9DmdLMz2P7IHi+YYpQg
mhCPXX/uDBOtq1wi+nnTKbloifMD/SDTdvmqaT33KPbqBFRClctgc1AzUsgw8k9F
HjDL5u3lZvcVo7qi4mMekC+u8wAuG3tAQnzwdbJqOLOoPTWNQsUQ9gC4qnrhsIiB
cHkKXRCY4NqOpvmIURKHTn1vo2WOGwU/1lnLWL9wJAe9u8ITo/4ht/QII1/78e1P
fqKqR/rY0kkM64xF8ipPe3u62RQ/9MEbLzPHg/S6czpXYLg9I3MfdA4zHWFiyFue
EQW+obkpg6T/V4VN2dkFQiD1GhGEkT/pHvtU5iioRrvlKgSLAcLdtzlSdknkf16n
1jFN+AZ84hDIY2pqCJCefT+FCgOM8A35MMyl9we9od5xG64V09vqgzbv9FzK2dMd
8EACjaQCWdJdo6mT+30PXWPEpvQLUFsIB5hvS+sZe9NzBICrhy5R2dqsE6PLyPl0
Y/ehCXJ/QeOZSYlu/ruWL9Z8dnYOSLqE9EoisVpyyRK2EFctt++HRWz2Lqo+OwUC
oHxL+xom2OfejFawV9tAKez3me2ng8zCJQzQCVqjJsIbc9zLmprFWvtUpxMlEQhr
cVAesCJAxX1Ml7AdvQl433HZ4dnQJNSNtH0wIPS2rwyo6zaNb/Z7QrL9o7jiwqtS
e/A8Sx/r2ynfNKDgZuVSmU21cAIaZ9byaqpMxw40W4MJOgW9mjv+3FWZsy2lehG6
m8/mSZwa+NeaB4q9sU1o6sr5AdzxY97GHDdpDmwD0cyxbHZIYZ8H0UqZYE7sdy12
I04KyyIzcb37Bmi7WwaXYM6MeE6DZbUc0f4VORgEU/V4uzhWxDY7uQfTiSZvAiDe
os9hW4eMT/nTD+PCqpGbTovohgx2TdrbHvz+A4E2fuC0I+E0rgqi4Hsh6L+p+Cco
++Kgfj/5ENIaGhSFdVIxKheDbB+Gl3Vmvs5jWFvvaGo5IHVWHuHtupxWrubvxx1u
NQj0hDKwQ+Ll5UUL10wV3HO3m7H6ga/vjQqB1nn5HnzWkWOWKPDdpYq7PoxjeGJZ
2dKdVJ7nsoIe857AoVOPr1KN0o5TPqUG4sgwKvp02tq8Hb9YxsNA4+PVVe3T0TTY
VezYhK7nLNORGPRx8NEz/RpC8olJxcaksfDskLRPVH+ef0rt2oHgSowBzUXpPdCE
u2o4lssyuX+LV7bniC3JNrM6bwrS9Y4KMexRPuD+EKOTJbk8IYnBBFayhGDEUzFV
TXQ+qbMNgDkAXgnDdpg/5KPxQo++o4Jua85u982q8rHUZLTASh1bN9Gaj9TkpKWW
EuE1ZTa+zJIsUkBCUFk+iG4KM/epUxhTbf5hY8s/KmiztiBhrRyj3IgxRz9T6Y7w
kl9jMF231OJlWDxCkovGAVcJgHbE6F/KW9tBvz7RJ9jDVlSfpaL+vij0LSVTc+VB
xbURSUYlh+hMVj4M4i4AlwDZdtPbjrNE7rNpKmtakF7Wfg5LDYjlo++uvm9E3JDq
JQbjlJR1l7uuRULgeHW41iBcmL+Vy7fEINtMc466RfbJbbjqU1lDt2FN1wvhSqXB
qlz0MwyD/40nvP9t8kPNZnovsQZPGR0HgEg/EoWhE2nh0lQUeAYgYcsbChAlU4dF
hModN3Wp0CQLtd/lnSvftscaXobXbDmkrn1n9jvl4KmNB83VzqIqHVYIwzlVZ0lW
t0F/2D6L1j/eKwMFQaIQgwbFDn6aHYmy2maX/m47qVvppi7zZG5GbG+r4Yu2NeAw
ExCow6XkWv4+BRVvZyPWhevvUFAAs4+a0rOnmntyifEfKzH4C7OtbXxneezLYG87
Dye0RAWhh/vBArkt3DfyDtLzA555tI3sVsT9v6U0lyhkAFOc6xun62MSYM6uehTU
0UgghSZaUgiLCfYCHa3X4Ijuf5H0aEJx4vwPGJFPXXhHJ00xIOH4bINFQsjeH0Hb
LaYrQWRNNHOUE3GbwjF6/wFkxEHRm+RKbHRd51k9CckCe8njW/Q3so8/wLnSf0p9
UU+sFtzClL9aOzg0bed81LaBjTJaGbzcgwHejW1ZFXDsjPetpZlbProRqPw6raSn
zzyGcoTkliSIgD4vksM2v5f6HEBeXEaNCYdvQ7xBNFNG76Az7jHikbu87PRsm5uo
62lqLXvV5/ZUAJsr0VPstSyPx1eXDRc2IWKZSggsgimR/DENZOMOUs9VxOj2+c4y
jD48m3cwFcLZdaF+R4rk5+QsthgZEF09NaXJbHIgiQTZlAdg2xpP52AJjc3z28G5
NquLkbSN6fJN8x0B4Qlakr4rbMmj6s6N0vRmPwktzrTbxj7K00ikS9weobpDImlT
zMpiPz6vmmBrc72oHxtZUn0oZ/soGxYb1GkBHpKCu/yw+yzEluLhnK8OeAd+hJS4
4vhnWId2M4Pz8lsumPDfKudpRMhkmKXUtK3SlPUKCNCZhnZET0UazRNxfek/aR6K
Y/zAIp/iJpu4fSYsUPX4uZNrj1GKO+WXpOVNeQg6zh8lYuPEKeqVDFuBAJcqEpeK
O7NcAI5x2qBovY6jywhmeK/VbVRIhJPtN6wwmAlwAM4DXOw87I//SOztQAYThfM7
CkHqh6wlHeqYJQ9WI0fh5Ntw7cujQYj49VI+4XQIcQTokVafFF26SISJOIAro5iR
eBtkAo7WjGuWCU/0VjiW8PyNwPN+Kt0hFwuWgpEwCsxLtqNRHTtoQdZjs/wsvFIN
qQRakmVxmc4iRnJRyOuZwYKJTvfNyaH0GdTlPfgWVPPMhtWXt+AHY2lOFTqlnq9D
U5LhTK8NISIxnRkjifVEJ8rOFri+U1A3lwzbUtiigaOy2hsBG8qX4MMQgiHdpPBw
Qh+0bB56VIs7bbboh+B/xCoNqnh/fMtgv1esH+3VM8l5GgkWoYb34VNRQ9y1azvL
DaYvx4fx/qkVsC/j2z65VtYsrQrQF7M4eaJB24FO5tS8xSDHCGe1SHvdGNPKcMuG
wOOVtat1KXl6ATjXUPU+NGxspIk7CMOfH47Zjgt18uizjHgldnQJ20wjxfjcaTOl
Lc0hwT/90C5JirRTYsry+qkCT1J/r0oDMK6/CDNDaYvMR/dvDQj75CfTY9jZGpa8
lzhuSBJzN4vwWN81a3mBjIOU0KQYouxNxIqjLljPY+qJslrOsE5+i/S6FQq+M83I
o0hSuG5zKharfdcUDK1SKy883Tmj8uKL60dWh/VTBYYRiBuLoZXtxnTlEfJxivL9
G3n8wZFhs7EvBFvSvItLSe9ZeW2ZcTM76y+ozlz+W9NB3pDcyQ39N+Upx3OLvQPh
ubLpp9ErAxG/zR7jCH6tUe3iRtwPZdAGbMeZit3VVX9fBNU+pckSiVgFncQp1bDo
haQ1/J8yXbu8sg50C01xzkNZBUnVTpohlx90+rkf5d4pEqXvYqdEnAsyUHVvfiW2
B69AKZSy95SR0v08mJ8iLTfQ1VKyaPfGcCty89RpqKS/XBN5rHaTV2dT4g4M56HM
RYKfph6wLFRbu0I4VdypjTwciSGNn8puUKKPRIWl+15r8yFlOo5N31sFCPjpm6pu
FKBuUqTcbziQI6MQ51Txf2nzOJroIy+qv4j6CD/2oZTYWHajRm4dHsavG/fOD5h9
vK+l+hD6vw+18F1xPuephtDMQvvyEdqsoED/S+fYBlJP/iQpRWvxzNHxJ+GEYWZb
Tt/f08u8K+VApt5FQZOSRhYMWttJHKX8kHrXst1oDehqZIq5EKeoSYdXlvjSkJlz
kdj5RBOGfq6g1bDmUuAfFtpSzCXdcfcyoaelp3w5eD+R0rQpW/D5E7580MS7Rq/N
l3L58m0i+0XV+YDMTagQMjh8sVRmk8rTsysDfpPVnPArjs02NXDc7oPU5HBMD5cR
4Ix53YfLiOh8tweLP0shWn9iXYaVvhi1lYuCVxc1Q1r//zn0vNiE4cRExrfa+9Qt
g7yWJDd3CofsHrLpMYuObMP/8WTvoVXFh7DVZuzTPxRAScO6msPVAgRomaRlUGis
n92wugo2NxHAWLiiMhjrAsN7vB8qQw3KIB7LVldMrcpAiLxRjhoBE6ZFVcVEOp0d
AycEOSJYscmr9gGDAFdTFCQ3BcDbsN6Tbiv8GmlG/ABGJ/bSHWs80TMGTl7gFAxb
L9U8iXavBJndv/gP3KG1i4/cGK5JAMl5xGDV6e/X4U4LwyFRAubvXsIzpDLqSIZU
IUTf0eqpBdbSIeMb33vMV0xfIvLp8vAw+oEebJuWiDwhY90bOTEhAc/bPqdPd8Ob
Nyxi+Zx5yG61aW1Htx9a/V5DC5RBBpMnI+AJId4YnYjHs9freW6Dncj8reCP9Y/M
fsX86317xyFNHtZViZVG5NyeWSwwQQkuflTuovZxDt6VHMLKf5zebooI2Jj3fo8c
6VSfl6Vp+Q1ZKnBAoAdYMlto4yVkb38Ac8QlvGPPGN4iWbB8ebbJ6XEvckd6CVzR
cATRlU0RHAVCJ1JwRZmVxlWjN+YPMw+2jVqOHreQXIXspiiapaaKrzPV8w880Y+2
/IN+CgYO9AQDEu8EQWdnZbTPGrsVr6qrBCEv46ZqEO4/pghC/W6oSMr7F90+qS23
RGDx/SaWXgaXjwfOt/sLbK1riplIV2PP3jHtZtyAT35K580LJKrsWKT68mjKjIJg
6qNmeA5jrDDBu43RT5ETMlgnlmelFkGWG0OueNi0+gR2WGIuksEtKN69G0C8UjaE
QIwdGbct+XL5AaX3YANZG64+gzJ8fsOyIUbs6f9J268Vb5l6eqOFUgOMIDSb2SPa
+KaXXzXTrZ1d9nvRHdR2Y/NCiJSSL63zHsDcRAaCa2Z9h+3ZyKOB3GwoVBfM8/31
w3IgmaVlp1GwXFCYAyiCiFW2FDTJVE8E1aXPVAjSy0IEwoWjLqxrYWqqHYZdND43
D/dlaZpGcBrAjIIgeG+0Py8pB0gpQohwKcmXW3BQXJ6uRTiKAFMryypMfs8MpVxV
JI8plgLrIJjB6l2l1uPNY6pVArZ1pX4p7PjzgnX9XL+w6zqiOpmM+4ckiYJoM3oO
eGvQ8qsGrmjXjOiNgDufLSjPBGRecxHvqk6Be1gvEjpZYXwOnkT5gOxlLiLPZeNg
YKjhWr+E5ZitxBrNvTOX+GymO26YjM++hEMEmMlbdPWVCHPUVBxFRjglmM1do5v7
Zl24KQYbU19xZkv6BSDnIWLdZ3uvTreVIXCbudMw1zl49QE6iFvz51eXaIN624tr
ip5Rh4L9d+hjexcvvEa2bz1NKZF9rpK+Akq2sWs45xK5zRWolS0gYBYcR9MjC2Sl
xNraDZCGwRdQZnDn3aaA8S3/WemLGW53dbMqvucLdKV5GBdoA5r6seObbDClTkeI
/apRiXRC1e/rGUb3bgxnigqQiVDWOCPB/itNnLsfKbkxpL+ojAGPlfyJl6HHuB2J
q5tRZlYOyDRwFKl+1n8PvisNaN9gp+7eoc1LX/4jP9ruUCO1tLrOmvpty1calf4u
w9wB0vRN5AH6LruVc+98q/FZlh6HHg57TYVBkLHVu95RUveTnyYCjRU8aXorVVaR
hzuZn3QuvLXSupJjUt7wUtyb063klCa/EjiPsqWkMxvc0EPLkKgOdg/NHVQUegzl
TykVRhA78t12W+K/lQTX9h97RXb28rYvFotvXiSr8DhKPjSxixwf3tbjqFCEj4dL
3Pl/797jjxRxUvcsHauWxnS0ToevBa7p/fQj64Idy4j5+YXPXHlkxk/N6pkxcKq6
UcIAqMUUBJSXfFwbOsefZCCx23+7fr5dxchRMnAKIDqsfUorWXa6WzK6Rrt2lEon
EPEJUbXMiE2FXtaiY7olptr2sIPCyJHJHO5Oxt5zQMpuB2KKdkbAV9w3ITtzx0R9
FOE76FyTAIUoYr59pWQVQblgBSytt8OkLwKSCn09zn2ZN9mAH2KxujVWtldVe41p
8HRZjze3iQAx/ZuAzqNLnQXwQWmRnnuCpgovvPbPJZsGfpEd0ZO0Z2feML3BBlgf
ENyDWFO/ltha4cdIGI0WwF5sz7VRTbc7VGF/WvAxtEcreYaNzpbrEuKNyloGQSSg
EFqW2T6vRN+cBQsF1xDqWZyBM8tXsDOab8PoFTZi5cf4clv22W8/ghDo/vPv7I4K
BhXNnShua+xWW9se8O1yrpfFWllwHAHCeZ17tepfCfMF0ys3F024GQVMa9T/oMmT
NW+kJBVqMmCzRVcVdilgN+6phLhre7I6w9Ouh6gj/xQg2nLMDDL9d1XbrYmiUWrA
qqxpORQHgSbKW2XoNuf1Y+V0aflxH0EZsSlGitZrtLauqtBcBdL4sVbYpnE1iPmc
jhe0rlQUTLkpmPsgyS4l6UPWtrRxlV9V+Iv7D/4kNETmX58mwwVwLFXa0wfCd7r3
wdxBOQ5aVHSkDTNNq9zURTNQo9EhnglemNzYjcRm96VrolHURrNq9K4NlHc8zdNT
11j3Eqqi2qPQVN9IjIQTE1PP2Pp3Mf0tVMIiPpR44HuLdRKPlp330ZIFT96c+nWf
ceP7iMds4uLwdUNvWC3L4mNjiR2bhU0SfLtBY3Y6lg1fCvFa+eBLsDJI0271MZU2
KtN/utahcM+oAVFk4XmJ/Ti1ppBkdOQ4X3Vnuwvi0WnPsLyfLpinG0KXgapcubxd
1OvdDUdidjDl1Po0nB2rnYxmTiMoEgSCXGCEFnKohOsPxSpddg0pqr6yWWJn03mt
uQwmR/gEblfP+n0JIt5Si8WU0gQQrcZQPrvsTZXg7oTi+p2UwmtQ4P+Gy5JsL9uv
HnSZdyRXh1j/h0TdSHrQPKNzhh+qYjtT24GDF5E4Apgn1sPS+6P98fWSp5PI9ZBl
gVZncySoaWgoR4gw3mHE4PooRAZreMyGQmnunDFmTMCTV9L15I7iLfRT0AxzBkIY
sHgOLqxsSQZBlNCOeOgYW3JOWSBgKHTYJsqTxVz+CRJJi+P3uTbR28RcvpPqbMEA
/fdyvcZzZr1D/1WEG14A3aaf6VnuCmDc7TCDs8zGMuk7bUEmhIPN54xlII7xRKb6
wd+UF4eSdfj576YDxQo9m1CQ9LIj6lJxZezdn/0zOfJ02AvR2Hx9YMNYBM5j+skB
OQ86SUMLLFnBRPZChY4izHvw+ZDwJerEDeREyzzMUJTDGqtum1889mtc5b4IU0Mc
A+6YGobtirlwq2kZuUwzw75RaM6Gg2RzC6TEFN9qN8pwS8q9BHhY9v1iROFTFwiS
AEu0dxXMJjDXvzTEdw1IfQ4ooW/BFzSEd6y/20EKwZMPY+3+UlLR2cvucuqrOEEm
jOjaihhJmzSMwzyk2abqvizmBlpGuLMz9GSsuUCmd3Lkxa8l3VSVXRpoqOaK/qDL
VvhiEQl8y2bU3nqli/d8dVze/UsmuaPr/8394Kn/IoWHmJIC5ZZwSxuMXPIpneCC
PRbSAvz2q9z/CuHf8A9j9Pa6ohE3JcISniAaXiRb06QVZvhITh4jGT34uatRwQXF
niZGspL3N8n7coRwTp5ajSnRjPrgShtNxMvKqXxAgOmy1cKkhMNZmS78ikCPMqlQ
rAG5QyUl1KfAb/9ktCg87RiPVBMi8UzwmUnpkurHw1vr/3/GQVNmLGjZFYmWmRul
qLGoB5iyY2aYUrZ6FfXljV4c8/igNF78tspJSHg79leOZoxywf+/K3e3WVss02v/
ZAsm7XwJnGvzjf5XFZcbLLBsSDlmIc3PMIsrPyAakSwWgtig5xL4gd1nUzyX86N3
7Te36rvw1sOSXwBLTEa/kAct5x16YucF5L3HLxHqkGC+7c+ySv357fq/HNPD99nZ
NEoG1t7ez3wD3dyH0FzXmEIp3eMmcUngvFsq47RyMQMr96iE7MOAeqbBvPEJjQRN
vKdmjCKfSKdSPUP4UoUKHUZuVkXERFGHns8DSQ63nDQrKNydKTBIA4KjepEX0rDb
dfkokdVXBxxRhvVEg/ITloymt6Xc7NX1npnSavHCYmIus8Js01J2g+9/gz8pLMfV
ySXuz9v7Lc+9+7YdY3BK/VO4En9ncU6rrjps4YlG1zK+uyoU6yeNGQM4nCHeJfY/
GJSabom0EuV95jO8FqKNbscQh6/gcXYDU16f3oFQVXQI+/5CV4ecfT0Qw+fqeeiS
wwnmAcUlQr0qhurQaI1Ov9bJu1Gm6lAfIr1imWU8Kqro2olKUGi6Lf93kV/RvXeo
Z+gwf2XxCbgb5gwd9ouXF8T8owSnLZnTJ1gRB4yc6mJKAgqWKDVIm4dVUdESe8dZ
qy8FTlMt6mWhP6Ed9mGx/0v6u6tl1IiBOLeAlTnJEP05yNocSIxcUHgCFoUUQQUb
yYDOMiwbY14nPp9/JZyeEEfCI2csCdc+CqVSsF16cd0eK364NqVH8tlfI/c8J0Za
x8J/d0bdksmO9ItZzW6yJofmrIl565Ahw8NL4z66HJgu6PmGpf5NioY5a5c9oPba
jsQukk/RmQAJz9zQz5a9/dP4Fkf3CnHPaEDQF/MpBLeFNRzR7qjKbUhh5tOJ5ztp
ATfh41tY6T8/KrKYaK/xNRW4E/EcpNogmLvWVWjQBthcK98lYdZYihieeich89SE
mj2bGWKWs+/LIRfDXt5Q79GVnoYgvxFR3LRg9uO5oma5VPpv2jeAweAGEue4hBVF
QthklKatXzHH6sTyAvS1A2/JR2/FsLYcYYbbxBflafhZZX7xf9JMHSReGXGVhhYo
knplWSP8H8NthdGnYVSIl9R9Fqv0R5x3KtYZyd1PyR52rX6Ev4A0K9ZgFhtoLmtL
cYmp4H3OBaUSXLNFb8hPgTRbZ234uQaYM96I9375hFeXStCP2nR8WhUPdDYFLp6V
UeKKpbuqCl4PoQ4F+loti5oKnEkHREYs9jPEfaPW1sxOdff4+99OGSpHJOfmLlBz
s/KdrHUJE+zpvqckSRwYBmGa6x7WcYxNeOMXvD4K6arG26h5HCOzWZopIaCXXUgA
uaZLXhhFqutr46Srky9xNcPJViRzIVZjMADXfupNBHuoZ/DdxA5VfPTYwuNbt9Pf
/cETgEZds4CeF+2LgZXYOFi4mpk+NNQ8vGeXOsqyeDSKZ+yUM8b8H01mMw1PrnOg
mjrbKGZtkNMr6fSMY/v8wk7aKGm02fjzQkfezlO42X/vUzSfIMH8N8AA7GUdAEaX
ZucGnJ47INo2MN/amq1DlKOJTJlnruHfvv2zUBYz/1HsW3xpIi3KXVXuZNaB5H9D
7Jd0VdHZBppn87NfbxaWuOQbuxMj8bbGP/ht5A7bCz9tY8iRLK5IEOhGZNESw/xI
/28vpiwY7N85U+CxurqRcu8Qhkrw5xQ2dw9STxc/tnCdsZWUh4l33dmwDZyfbwok
U1AKfXFCtQJ3po7tbzr46pr87H20BCtgJaSfH0Pu+6m/Hq8tY2JRZNwnmPafaelq
lXW8P4zndMDmvU7yB8T5mdYlU71HG9ut7x+24G+/fvlWB2t0/2uWbQBCdyBzkDmq
BOHCtU6H6qU96QaQjDk4EiPxrBL+p9RQ2nmbOsDQrvFiUQ1SXA/qn4JqVJmid4k7
UShG1ideuB2znCG0tJdia8EI4tIGQ15ReP46CI8XhVIuDLUClWm75as4b+4xC62p
q5NV6wQYEY2vvXHt2TtIsrDAD2SA3B8sk00S9G/31Xshbbg7muJ7/IHVqAyV0Kbu
Rnnw6JQK1D/t4z+NYrkuSITh+9WXoYB2ilPXtvqq0rCNboyWqebGhomrUAZ88YZo
jhN7cDMdiNY4PYSIgZBdkhAuBSxW1+wHZISvfQOuOMFjoIjqTlvfnSDHsPNjhhT9
FgyQYM3sFPiP6xQkfscmj6W2JtPyIOmPwLO21Y6tTuJbUqEs0ILxi4cHrDlzRDoP
jpaAMvgbaM2KoFF00GSIA3dTh1g6x9IlBcroC3HaBq/L4s+vHU0IiHMQ+OjRPpTM
+csFw3wxHXTsXM/cBaDyn2H4B1lsNW0G7CNLnl4Lw19S0oWUGYKQlbkiAzqkMrkc
/G9nHFZzLm5FkILWfYlgM+Dz8RfYGL86rxWdEiayWB44mBfWnkphasXp7uqgxNpo
/B9FdOwaxUAK/TUM5vXXhWg8BqqcRVZ5rP97On8e6VIFvzrapEDdWe0G7sLrCIca
XJkDawyRTfDrLhp0lZpKcAv3g9lXVv83ra0Lds+z+oKRutl64SBNKbyLRYKqKjyh
dNT9PEG8BlQTFWj0j7J2D+cy0+kIiRHnYXEQ2BGCPin5VGq8QzWXO5W1tZZh4+5L
UY5d/lIOuwghZDdjfMqVMGQNnlwEF4PWsBmlNR/4MCs+NL617PVsaC/OsciOaDCk
l3i/5eifQEtWRfyDHVCYcULGMJAdO8v2dXcinMxCqcLvCkRd4Bkmy572l1MB16Gb
ZnKWTTdki/R8jqllpNFuRZUvPrPeyVDgt+FNMcz/Q/DzCkjoy3/QMerwS2K6xm7W
ARTtNWnWDcuWoAbuVcNoFa6nSapVk3Dx8vqZoY5NFRkX4Jx7gPkKvEbwXox64xo8
nMrze7ygCkIhy4Ear4M+5oKLaMxys/rJYR8RiZAjD+etL8cWV2qoU4nWDwKUec4q
VzyE5ANEref1y8UNkZ1j5WYZeUHEWA/po1mxE9+xX+7+xG1wBcFVImoxuSuA/W8c
PdbmaHgQFeVvGgF6fpVIzOFYdTy8VIkcB2kYAzNhhVqeV134ONheJBXnJyGRHvBd
HEsAtA9mQzLadOu/uMV5FSo6ZB5DTnVEJfFQ1th/QP+wGI+E5pEHLacHu4dZJ8zC
0h2hFdH0Kkv6MP3TFSegbobbxOfHbHfT9nOJHbbGKEtqZwC5+qRMARq1CAmPYO79
GhqsR/AwdCtfdiEVKxj7vlssBbqMS6gZ3K2qHPiI/VmhKwqciPR5l5fKvyNes1nT
/rQIco5lm2ISGVpH+R9v098MxZ8I+FgADTXp8GgNdQgaTh6xeMc8KD6YWc/XDo45
fngp9FIbnClQvPTo7/s5yhBuDbUQE3qx+hmll81pMZYdxDwkmIF8lx8X4kx6RO2f
25ufLCiWIzorTWPQWNG/zCdfNUZ/6dj1rPOxQegXdWf1XI9HurBoJ8HXCW5mCiEV
Sa1ujXAVBHG5HUgu1PgfMrThHj5mncVRZl5NCFXp2LN929u778LPjE3xuB6PG2Vy
uCDFng2uxuvCqMLGGKi6U61nbXNN55D7EjCD6OU2igWk09UKtjvSzKrJSrGMYjhW
dLWzCWRMBhFlVKPwCzd7kE+lrdRTh5e4apmrn8PkfF7QyO4+B3pFIzRShHjzDLfc
cPt4gn4jhS6F72A64DdrHikFeVQTs4YKlLQsYF7UE56+HtRZOWppFJKNOvhG4Nuu
SqslTiZTOgmhywmYHl62NCMPRr3ekMO4y6v/f9OcEHwSUl1cfMqSfufFnhJRE6F7
6mzCydjJRr9UG/pto32ZHdEfo5/sUUF+Lo5jeg+jUY0pAtWSsaGdUfphWgR6NsIY
6NbNH48jK4Yo+8EhrxoA0CIuMq899D7f74+ue5nu8i1xHuqO1wA8ZtYdriO7OU1G
EqeP3Xd7KBLaXUB1e/2x2GRXgIDOTm5XL4b7KRVyNK/1/QV0ewHN8belkN2dYdEu
TtyL6F0qzv//eHCfngr05YKPkn10ddd5mwlS4cJAsLtQZ3zjxDMwL+ZWobsxi/0T
j5MM3k3H+cFojkqL89XEnTI8aZTCUoRwwhJIEBAQROtaraSCrfvar/aYVy2LmSVq
pVK9cj0gQgD7HK3O+6HFTaOWKsbnSMx6IiETQoITXhqJYFdpoN6+O41Jkjwhz/IU
m6GgyzM270lUPeeMu0tQR0jl7JkbIFY2YwOlYOaQ6DEoPrf+Ibk9BY6iHSLhIz0w
lqbg23GSTdyOQ9jRI1GngB5+TNOj5cx8nf4ckbZrhFeP51/dODE/9uXDO23JoysW
ytHMNokx1eCFQIhznRB8CYGh06lfKAkckntx9RpULCCcNQ5KLICSEe3RuaZzoVY5
fIMPgHyuwL/hHg9YHi8gNEwyLorvX3uzNZU8iPIOKoA9Fn9qbJMbG5fY0/X7SN3w
1QTm+x9UKPAoPcQyeVAN3BOQrJWUaDoJn4I/iMxv+bwMqO4SgJRAq+Md79ijYbR3
XrtcPa7C7SzUG5u4sZ/WTInwu83nbQWiCY3LBq5HfB2Y6sxH0oQnQ6ZaObG48vLJ
LCKeuswq47cCE8+snUg0B8CxwNdaeJI7Rcmv4oQ544G4N8ur8QL8+0fRb7KwaDZV
5itPd3BqpPvtyBxwKEbq+Ovi5y/LqONx95E9rE74TTylnFCDsuxRyvnlctbddH8d
LC5xCTmaWbdSJNIXIv/rfjw4VQw8uzaRHBZxe9zgycrnl8cl44baRXa/btMV0pkV
WLES5jq4eKvmHS/8DiNoQM++iucAEqzMzXlK0nFNEuWZHjJVDH26ddebGhxJGkwm
n9lEPgQ/eR1ciTEF+8p1DbnWKDd+xBfBO9e21N9ggac+UEt+Q5IDCA/tYkG/9wvj
EFkI0AbcM7LwHmkQKhW2ymi8JEIP7c0uc0z4gTGhU9aYkHGz9D6QTXGUhQGrBPbt
297yNyJM1vZECcn6AuFmVQQq2+F1lK0fmwV8SlRjt9LjQa99EcFwJIefdHWO5a1K
+Sb7oUlJMzZYet35/RulTk0EwpmdNCu61mVCziJLoaiMMCHffeUWd/LzsiUAjpht
X/BYHdrfB98mkf/9sNAxpkxqDUi/FrAsUrZBzmHqrNQa3CSlHhANlzvfW/P25GS0
OKTNSFmSmgZwXFCGejSY3mnwYh8BQTmHIGSQTf8xxOabNsyjI2jpob9rIZriIj7g
pAOGtHC/Ibe/HBTT1s0wbiLWQGp/S9kkjEhJqzrO7inrutFsWZkxvFkblUqWAgEu
s7EazBB/gnOf2pspL7OlyucgmUL6K46u2+WAs1SiSr3gbkUc9UmJVEOgK1D+ugYt
E3ndAaSs8UTncPhkRUF1q9/JDH9fJvcPg503kfGMSiUsdgmoELx75SlCapOFy2yT
b0xS0Mcj5Zck6/BFiiaK906A5WIz42nyKPVOrMcQTnqCfI8n/FrbBQCMNlDGpGaX
WQpM8vkSYOnbM95qA6nG4qOHsLMNjFLPl0s103KCb3RJEzVFx1lrU3XlbYrYHFN5
/xUcwrkPTFuBH122KKs783D2c89nFwaaZff/bx4or2GCNiCUIow+3KgQb41sd9jU
QxUfRcahd2W1uXeN9BUO8hZK1A4nl9+m3Pmhv7/uZKZv3QRLbQoCSfDbwdf3hm9t
9hmW5HKeT8CjXBNcTIcYplFRjgnD1JHprDKXwPDbhf2pERk40t2yqrHj8YW/7tgp
fTwU37XMP7qS5+d7tR/NjIhAelvkrWoQ8ubyi/CPVTUgErRdW6OKScqx0TnBkzw0
CXSfOx5x00isttiQAAytni9qjLyy/Jnt0rrF4iqtdKixmGEbeDuwC1lYJqRdszs7
b1LvmxgxU3yV0HxbMx55g0mRvCpCVAHd2t38HYQEjstldciClgcIicRJVam6+okQ
sORLCXAD0eQMWbBIGHTmpZcxb2Nuf2KyYr6LQVG1cY0nx4aZSbfCuPhVVYX/Gnwj
041PonY4PQf9SNFC5cXU3rIDAIAEY+j29636Zrg+hkWy0EUVePZn441amk5Dqmu3
v6eNTm1il1/AuZ0Ki4dJLHB1uvYlRK7Pq4swqKAVvHk09169GMP+CSXs2szKYjMC
bV9qoXEcGerWRgQQSiZXKP15/HrSj9xfxthwvNk4hEG9F/3ZBOraWPkrUNJ+VJTH
iDgYN6uBg99AM+gZbGmiWoeie7ZXzpcFv1AuHTRiT/U0SSOiHhzS9C/1+YvOUtyi
+2z0K1cWnoCWpejRYGmZbhncjaFUbfq1ijwdJ0zA1WpZykKtV0/wJrXyzzVPRMB7
3e1DFuebcvZ2FhZff9MywW8M2mgogwozlQng+/kq86ityGbFrX6Kh4KtJrU4xZLe
eVesomNB/FvcM6AjxkvgNacDf16SC8GRF1KELsvtN5FU4J52CI2dEfPd1D2/a18s
ZeqytjxLtrNUT6WYIHukFUMcsyj1L+BQWXTtKMgHAc6L+dlcZ2eTFq8Rbtcx4GAn
7En4wlLKMwPBqGPBiO44bXaE9/yCY90YTQ17OOD8FmyeRi/iWICUm+ajCFkV0t8d
1dV3pRC0ifxLW4jOa4OzyrZbu0mkew90g77I2/vP+bEYeJYp+I8iIVLHm6IF5GU/
7ZKYE7YQ4A6nJjYcOmMWi3zvoTuQpxHQlgli51AR1XLkgzJ1sRRx1Jg7cAjiBdyC
mf32ULIIkKxTCXfFlATaUtshaARz0iNIxml1/I/VBAhY8UO5iC+HCJVR5Sas9rlk
7LqWNHtwjSU2Dakho24PKAb9kK7z/VRcP55TGeUgVPPzBfmqW7Q1cJ1obZ/cUtdf
ZbEbmc7cevD2ThPHlI3JM4+3Tsj4D6e0zTFOBeJ2sr2/yjruIxXcwD9FmZqgC6wE
JfGQmso79YadXeRUGcKxOm6wNDopmVb0nhEoU0LNVhF5P39O6VX8J+ZC50J5yK6A
93whJoOCSaLCCJqgrfNhRKkL9469safi5GZLovJnSNDotIGsluvSdah7lZv2jiDa
GxMY6zQtpn6uS3ls/oAMmTWkGWnnx0AVENNcjJ+ZqVX/RxMVvXoIoGZOnoIiWpOh
IqpMmKa/aniK8n5XMvDanUBGiz1VD3V3RatG+YH5PU7VngnNS6HcHNO/ViznkFSW
XowDGH+BYrgts1krpvJoLIaBxoVPugGf+vdgV8kGAyByouec2LGIjqOainxqlLuv
3Ix7H2C6oGyzelEeliwNC491rvLqNrLoHJDu8poHHprVVHrSiBSTKEO0sVMixKaE
O0J/rlezpuiC5c9mTFAgADqZebAEM+wH42kAyZbqVc/6XDSLpae8PtwrY3YReo1Y
9YoUa8WV5Ae9MDHrfes1Mmp7IyR/Hdx7JTXoUEAysdHjmmAtpD/JRRjotxHL8WIW
217QUcgVNybi8wLpzbMTuk/prcn0wNXuKTrYILeY1KWxkHny5ZCQIFUrF0reInX2
xC4IBEgKkc2Tolu+7rtUH7q7l4qlFnfJud+kSa+D28gtaVhqeg4IY0Tbrx1BYY6k
8zX7frONmqC7R96UZ2KBA1jMO1YxkmQVUsl0XcmlmZ3Bnh8MGgZ3SAQ9wxu8hVjJ
PQIUsV+HkN8rvCEd4XtrmFa1K+fGXwIPt0BNdxGVE3CUopM3P6B1bS6F0PZGq+Dr
ZPO+AdoMHytErzB1UTdlQRRpcuFKX39Sh+/5RXnAlS3Ohpksl9PmafGTZeoOE0tN
mVV5uAjwG2eDzPtMj4RU3INRKy6gQhBKijVj23QBRk446M5dtxKmP/OvZ3zOmF/X
gUj005sPn4YQk+0qCC+7vmKOv1N6LmqgXXDweRkn+n8nw18X6yCqogGw3R4pZQ+3
TymmQbIwDIrDVQp92d8SwI8gniTdnLVgxYiOid+QEltcO7OghIKUXXsx+N7Q3ncz
MeV5I49HFW37IgTXtSftBg0KDqoamRelu8tRz8MXegYzz4y/C9lpbNeqKt42WD8n
zXp8qWNvB1pIz1yGYZldA1w/4J74lojeC1Cqq3Z6VEcIPqx8SwMv/VonDaIYy0MH
SpvXtCM5zqtkXRRmA97PxrcDvYBLRMxcoyzEk/t9FdqjUj/3TKaOg5piw+lhKR6l
dABkGLhcTagjt1nje0uidox88lkM3MNvtdhVjBy13JG6g00zE2Ec2ToLw8Lysy0L
xDC1XtYgo8goInEZrshrW2mRao+bT1iOd5d7lpxaqyBmuDpeyOLmzhB7jwrKeiWC
eHi7eTV1qwA8kPkuT35a58EFhda+2AbYy/G/vW52991KlF6NRqymISC2v4Ggy4TZ
o/M4Bx3xwRLoGOKVRvpftvqiU6NPH0wXl0yK2lG6o/LBQYwt3fB84bghoHRq2Psu
w3SiGUvaAPM1txeDaYbhqJtCmbOsg3/sCk9+gVuC8TFQ+BRqEjAyAlJ/0dD2NXM3
eIYVTkFa5Zyv003R+RHEViNuAVap99dsHYTeNyzuoivZzROnNfGxroWcBH/kSsvd
D+O2Con75ttoLfd3LwmJygkTF+qsAUofIJ6iEOJW3Jf0pM8brusNFS0Eer/xGRpB
8s1N5d655vsuZ58CHKKZsjRX+jWgzjY1OC/KFnvLsiZ0fnxDFQQKRN/xCgzcKwo+
GcnsZalBb1een4BOI2LriXhgUHoSLLfZu3CCeT7xy/3ln5FBwBv4LER/nn4hNpEx
21dFwhaLS6stP6OQZmMCqpWDFcZuMwJ7SQY0ryyyG1H7u6sScO7jLrUnh7O3KLnL
tvuIg57UQbgat3aYa4O5uM+kyti8/s9LLp1rXo+9uNSMNNGQLZ7DLrQuBAzCtVAf
fh/nnkZDZdcdCGIvF0Kn8KJRYWkOGQYoIqczFNkrrG9fccV6MpHoI1wSHfYbOLsQ
RKgo/s5v85JWHYcm1JYm5VS/pfn59NxD4ark8kpT3nLYxT8IIgP9A+BFvBJtZ3XE
6PZLUvOeQ0sgT764gg7qfdYavy23SY6AhvYYAl9rAcihB1boEfSzTCnhwtZJspv7
BeHpn7YjTrIxEViJCUKh7X8+UlzWW4k9vlH3ToOe0OI9dXn9gESIkNQrWjJuHoWR
+sp1aQ9tBHJ+42t/PMqIFxpttMGvLEkn8HqJUW01jRW/ciWN2q6dQIQan5dNS1tU
Ctdl0hrnO7F2YQ7NCQ6DlytzOAE/w7pOn06rXK73+YUFkyFSp1XDgiZO3k5CyvCO
UbzUC3VhO2lii7jsA5ld5GEzq+sfnhVESWAZxeURkkBecqD/utxPC7lnL58nggKl
wZu/Ymj2icK6t7HTK+hP8LZYNapYhy7rWo9TsoEYZk/ycLA7znTl7HB4QdWwXXkw
KBqRz52L4wNxQ2mC1Tvm4aee599YAoY5Cj5UzRYasgJExluMJ3UTZguPt7E84IcT
gwMep+dkHBgBSe6pkU/VSNVd8UTa8suBWBDjXwAgAu8UfONnfnFjKe/YEfLhFsSw
ASylmg87Cc2bnE65+q5xkGqMz5piWsk9jUKQJxZUZmrjXK8BF0JhdGjNlb5Ku0Q7
xSy1ZB7wdoTsDOBGtizv0B3yNvL03hyftpbcXpgOCGURDfNPBUbHqb6tQCUZ76eq
xe5+1jUUcUF8MYKpNxtwMRXJGMoln9+OO9DbH2+SoHC+Mcb0x++otbS+A/6F+/1e
8fI7HIWEl7rAoDV8rmlrQC5ZHbCc3YSlLVdo26tXECG5gbCm92QR5cviifuwskG7
TqZbbYY6xgQEhjNp9qHv1VmtZNYauFTCXAICPDgK6uuY6Wcgznh82adfd4Mq9Ula
F0orLEUnspPg1LzujuvyECl1X1KCIla2sFANEJbGt09YHTyQhJusfjN7U9kjm0yQ
CroupTao8DHWrLaOOo2zeyLmoXqeAbCNfKola2OD8ZH1jZR271eV/VYKANWdCV3b
Rg1TG1wfkagc3DNgWMBL+3XJC2lkPMDqi4M5AEANWpMS43Hv0p/Jb4GeENhkK2pS
78h0ohqSlaJ7X9YxW549ipuK9+IdtTJGNayXQ2ysTUXu/+ENMyYzdLloVQM7Wjj+
mzPzewkOQVuCG63pgwEmzNrUpqG5y41ci+BhHZiESg31QaXta2BNFtIXQUMknLiS
Ao122XFoGrdYFfyO1T8JSFppV87hWtSfnMVFZOgRVw93xzW2TC37TaZkplNYPssj
pRBsjRa59L/Km+2bF7WkAdoUSqqpApC4+WURKV0cpxrjklUcbprDalz1gEcVfJob
sRv9W05vO4gzTjaM0BTZW0hqzxm3eOm/bNPPfyghc7TnjgsPclP2b7tKHLWSwzhb
Z5FgGHqaZS3PweEg2WPJE2jh8eD8yEa+fKGvpS4ABWxNEFNoCUSKtwNa9HhIPY8w
q+kl2/lk+ZMFSiQjUNfo2ymOghpTXffqp+5VFiLHFzOPhWrt0RflOmAiq5jrOmda
Rs7p86UKoQjAZuTpDuMkHO+Y0ZinTKXcwu2xaqZkC9Nuw5jTpgL3q1dH7DLbMFgW
02ckteB2J+YesjN7jK1pYKGUSi2mc70YfqO9Mp+IVI2R4PxRMY6S1p8uKerW3Bpk
P/mUQtF4f/xz64W0gW7wvp3z0xB8LobgX1oOBO35aFMvZitiNHbeBw3MqyE60XIa
+CbdPwDqR8SjiNJE91lwbzwXt55Rg3fkZlU8ntF44++RTUxJXvlFqsdXaKZ1qGp5
5QWVhefKfuYjhE0JNJw03egqeri/RAeI0rq44OOq7LElWjLyElpS1zDHiR4y7JB2
Qwukecp5+6/J5g6OjD2DjSRGz4pVkUYpLwYprXcPRjntXGBYOMtnNyqrXYMcTFbR
9bX9zcglYtQ0aYFvAN4xBbvgM99yrWrxt2LmbClo8a8ydRZzKciq7Ctw+F8cncwM
4OgH+BkdmI/EYdgFKIOPLX4df4yTcEIl6A4qFjRhHAwHkw1q073I2mBBdrRKhqD2
iDy1OMM/GFsD/Y0rsCqj5xVdgOYP/Bno2SCmqcJ/efVXFetgfayIzs8mUQL8upcp
wE+QHvfbZFJ8bM0ILVN0Fu5kgR3z+0iugkZ67q+mmIut70OmnaUcY+02ngpcuGeO
4p4b1mYBoev6S0+zcX9L+oipzmGHL2RpltWcthDOGzjQY7J7lAusYjjMSbvGSwwv
6d8tPg9dhP92tnxA26VFlNd6c3RPGNHnh+p0dVN5Qx7r+0PZD/xdNZ9znZWmHzNW
K1Vkwp74yYwzMqe469oP/t49J2FNYCsv/R3a4fNBXyrchB3a0FAWgcsBlRmJlQSI
K8dcmQpPAXolXKoh0TZ1G40Rv0/YpV8k6F2GehXulZrtV1RixKx70O7J87IU19D3
q0NE4taFtURuXMAmzzxkUyc/BgXUQE7Vhk3Ig7am5umdUScknLOo049S9X7o6qZL
AlHG8/HSnSUZBGhPI+XknkmYLWzIACFMxQ8rfPmBVYj6iYXCSrdI9lRDiMZZgR/9
Cmrz9MPXsB0KwkkOg9Z7Bm8xgA47K6qXYTSOUIQNz3Er0M/elY0TVLBJ5OrXA0OK
FbMlPoAdCHSxC4xlbMLTuqMzjAuuU+6FhgdQmN3v4GX7OfDizQVaPoXwRklLrx1X
H7WObXvJvRUWElwfUzkLrGws8sFUftk96RpbyzcSedGhJ27Rps66+UPgwtlodbuS
CoRCuGjEPKPOSjnOrBLNh+aTfr1/qW0YChznN3blc/O0o7lASgVnBQmJ4gqnaMdi
SjemXfON+UD7s0UiyVL51ZPT31uXoLBtNxeAxrxN907yRm418ze1XpJML9NpOAUx
kJo4tIfKthJtM2v8rApK4iuFJrpp98nKCjOQHbpxd8Ac+uOGw8Y+BGl51SLTr7Wj
nVL90HbBgw9h6oOiLLGSmLQuNZm862JWkdA5jEmpzBCJgm6adiMhWPJXoiSfbSLO
xZPQ0sCVfXPFEDUC34a0EKtpzdE5gBTnI/oUndF5vBXsHCIacL+c6wHOKGiJXMbS
JERngACeI2dugkDrBGkoprTelv6F+q3KfPe8czKNpfKL+LElRWccupluYh073+dV
DCNUUUr6KYeHJfyTjMHg09Sycrt26GoAbTBrMKsOhgbe7HF0yc5I43MXl81BA/Ls
SoCfys593ZAAQ6xb2T6qxsU4nmy/z3/Va0tUJjD8hf8j9uIwCSupk/Xzn8mzSUMq
Zcu5210aysGWXDQA/IojXcIfqXrTqhalksN4h6jxYgYv0wzIQR52WORJdtsxnHin
g/8H9nKxQIL6bByhvNyAKw9DW3g0CGiMWnlXIkXb8OXkj+mgeEwqKxVZAOKQbTDJ
7+noEHPBpHb8vlQlZPByJLNChznsbmXQ2Ws4QopsBGf5b6uT4g36kix+TNUPROKM
WLKd7cYDe0SYj0DmtpElHvWcbUeWkx1uG21C2Un1BnzZL70A4z/V1NpY6V172YDe
2OUl/QfjMvlHqOhOTlnkF6HzwPNKZipD0LKGGdExijl9Z/oNJxJQiasPxTF1xHm2
mVg3enounNVwUWZCs5MsuRhv+WtMbIODr6/H/p0afmbTJAPY74DEHcjlRK2evfsj
yXDOZw7eUvkuzbQpf+EJkTRcmK/xHk5goRUXyV8p8C1eNH07MWQCgxR+zBVmvFqA
+pCVHT+VDC0InvpXGuo5MEV4+DtvCXEpgqxyQQJuLJ2oMsYexbgFSceWo3HpESGF
pgNTPIOBSEUSFlvoYX8XjsKQ6OQ/l2+z8VtrHYDU0h2i12XUFBptuv3fOGDCVEpE
81DM9YXthhJi5lhPUd0TcDLpQ94Dpw+dOdbM6FGSkhkhyv2s4jTEyUZcKKSA5515
jQbGhy1xdGU5XG4LS6rnupfVb/0pXnjygcQ+CkXcc7NXA1+hdiRAzQXXZS7B3cJ6
/FmP41+df9Sx48fGp42siH/es3ixKSXuBMa1SFbR4UaUbG4ZSsWvomi5GUgANYbF
Kpw3xAr33trPITARbo80KoCxfSrTZaFVrcWXBy+SFVRRuZV2DwE+XQ4VnAhuQJmO
fmUkGgkHjZONNTF12QBZpYRiQDj83hEIxsr5goGa+ClXAZJbZ4fpga+8/Wy88C1z
HDRc8RHw2EECU0V6qfkMcBcuBHOvGjHmnixAnFM3rxq5obSvI68MrlsDPALtCrPV
evjgB89VgIL7JfMNGZ17aP1L5bG6I3W4knEmuyvsA9o7rkbGf+znxRjEL+NlSPK2
IA9JFja9sWDsnul5xpCbsPwBMvMoWjnpp/rQwGlEKTQBicunIt8O7TmcPTolLqkb
vmXJX82GuxGHv+7h2quWFsR9tHd90OBY/xlWXF7Tnh8sDasUWt4nSynb2XpdGJym
NmeCfQTrJFz3IjmO0lE8aC3KIDccMQMRITssaUsjSzS9YWqV358pA6Ru1e1cRdja
nEBhWVlRW1KMfModlMXQcyI/iwXeMVvwAyGBXEs8iRpw6punKevEfI4ujmZWwPkN
gH2QuwK6GXdZrl9Qxa2m6aXLrYeXELkhJJ/Fb8b0NS6vMo11SVq5eZQ6fcQOpVgd
geQkO2Oss9DkgXeDcxfEOxhzCDudxBp9J08gydAUZpRt4oDujYqbVhh34JyuF45w
VfUMoOunbM8uf8YoepfW+Vjkmx4hJaHB5O06lfRQoFrtjrU8FmbBpE9ljGAr7Fja
hq4G0o/4RyPklcu9Q5ZU07gXJcht7VSYfZmyCzdxyFDAYs9juY8x8wcJc6whsURx
ZIKV51EvghfgHREtx6cE/8r/40TlFZjpR/Y/5PIjrvtlDYVKvcffCaFpaA+SgIwd
YbKPrQMy7LQLKsW8ECIhJ01bpCSVKAPmVjK8NPUIoCgVP+VfIEl/2v59uOEbQm4C
Poxyp7ikRHgQkg9f6PXPTtun24nIHF5R08GxvRpCyaR7+ESf/UDaA11oS60xPs1I
YxdFHODONHx17LJv/UAkiwxkzTEvj3N77F5f/s0BwIH1ESzmJqR5uN+qdnUEZCHC
q4m6oP/hU65/FP2GNeLvP7OOWCGV1j1KiFELW+jgeCrXKVVCmbsT6y6SPvkkRSQ3
+vp5DRvQS0ML5Mt2eAYIndD9YvOLyh3sud4+1SVAKo3MyxmsMjNRinTHbeZQ4mut
bNiYvVLYEHj3pfu4S03dVw0hq5oOmxT1J0e9L2dK4zlLyrsC6ECFjntCKclUnVli
Cj47l+ngKsC4gymdEC14VSYstlwdP0iCyKQjVKYzA16gYTjxkLBd5err8Th+yYjQ
JjZAXajJpPEI1Gv0BNGMUGo+X9xavQYmImrIUT2COFON/SAouQcCfDZGPq8IMw6/
sjwXRtge7sUUQj/vbxbkKm4MYCmhrQ8K4keGFRoPTxMNAnXdpWRApR0Sg8g8Gety
6LTVSrH3agPjOUJ61ybb9E/e504g366ElR34ktb5kag6MhsMh580xukpGQfeEUAV
z1yPTvCaGEgDzI0EbG8MgUddji51mKLMZ3fUHCAhZvWwSJQckReBRRY/Op5k9k8r
7LOghPYSwJ2+ugXpgvwJ5QM/gIYKDT0aAznKGaY4kDUvkKisvpxksD0xJDW7H8f6
oG5YFSLk04nPa6/bwzHyGrwxnf5gTR91uTvQAU3OUNPWKyTJqqQcejUq5/RWrXB1
KPmNovnozy/5qv751kN2yotqNjIFElUrPKsT/0TxRikofKLbY2fnYTcTn1jgRh7G
GxYo4MUDdXonketNkskOrmVrkYtybEHyZRURJMvF2LVxFWMLsE4EZvzSEciPbTx+
U2YCMcfu4cGLm+LiDIgIQalvQttYWqdM4ufbxH1pdhb96Tc5k7P425UW7SZZqrSS
DOWm0E32M9dKKvq/mePNiG1LGiCC9+wBhx+mV+WF5dZSKSJHsnNY8070Vtw7i6If
aj/J4roZh2k3M4BQ9ouDzN8Z6jiod7Oi1WdR2Fl4tp9dnDoyAOxXmyVHd7DmMxRa
6B7PVvkEs+rc24u5zQ0MzgaZhCWb98vNRuk4k5cggeszGA6FT0NY8RoN1qUEZ72+
rARfoeGQoILbeS8AtcmSAs/3YD2W/UMN29njEjMllrH6wQrP+n/9+CfbvAOonooJ
OVisGroHcxI/kOyfRMfEdt7og22vVsHnmrVz5uwo161CmGLzO6kKM2+jjHJwjcqm
fPaJLxGqr2uOrgnPBL2Eo6FxBvSZjggwbNQewrQLEBAxnUKfzdGGbdPj5oBy3eAE
ljsway5TGLLnsS+Ots2cGqIvbvT/z7xgqufa9V4lqfCQKsOF37slmt7QlJfKP0ED
VqdShgv253UJDdoATXO4eE7XzriqlyjCbOESB3GToG6x2naQCn1q5eoGc2igg0C5
mUfi62+n+sNvmuH/EGxo9dv9zKyBUE2oL5mvusEFme3S7wt6Pg9JasIKjV+k8Zyb
KTQOljDziapw8AZn5xBoluDkUr2r6f8AEz02trHoVeugX68FMJ1I9sz8nXwOS/Ot
HdDTFgOdm7MqRLxlBH66T2hi1ej4b1wO1C/MC34HkEc3n8bJzfzF5LZwn+vDKfwb
DNE0GVihJcKuXC4jzb33bEJuPE6s6suDFtrHkYLVWTuXtmkpAJDJrltpeLVqGe4F
gHFQZ/54PBnmTR8rBOdoelXtAmcCDQiR710k0VXAW5YlCbdjm5HTy5huv/QlR7IW
cPrOVUhrry14f8ijUXjgji05A4K5HtaD2+ylglJFY7LIuRUhLdopvoKQzZn6/Oxb
l/W8bkziWPuV8LHxizjMTHmSSG46+c9LW4y2qw2XoSmHCEb1WiXOd2M/sYJvupjd
mlCI8EYzPAcDnSekUSgn1pf5M/y8GhbH2NmGIdyVLde5sFo5kbnUcRK9W+k9nTt8
cvX0FXRp+v880yxdyf1oAyV/5HrVnaeWujvlERHwOYdBGMrM+4pLfh3U8zf5AtG0
YpzjKL5jwJgSMgtfuPjwZHGTaTlN7sMJKwbHX+QC5EKEQpwygsWde/rMGu8DUc3S
C95hiDITwF+oITJytAJh1x75wSchL1O9c/3bAZb6wm1a1HppLkpV5QWB/wGfacvi
fnjLkbmjvAZfmyX/2NH1k997aHAhPh/LRmHei05QS5L7MzKftKpHjc8Hi5X1/Eyk
Zd2aOTocZJmSc+yhJHji9Oorl4DwkQVjrvP5iKPFGXtuY47hCpESooFYZZi+VU24
7agaXYB87yaoaQOHEqLRKctHPXjU2iRqRNubk2DYI9lP//TDKK8OwH2bRyXFFzxv
UFGKrTCfTAhc9AIlCj1lIRgQaB1Uo1jCv+ysFahJbgvsjRduKJ50jMEy1Ktoir4x
HM+4yxYcFk6eZA04ZkD3ak1iPsKCDtfElBAx4Mg8DJE5N77oZsn57QCkhAkUjIdt
TmwfCe1aU6XbEKp4cs7/laa0jqsYYIov42dS1qoH3qUQ3LNM5NaDFXJxObh1oFmI
yLBmKF4Qw0soX2GZJMzlhhWFV6PG69StrLCqS44siABlIaKjxsTgZKCFw58K5iLM
1wZg5ClU0wyo2qoKrklBnrUjn2JmF5U/hHlHHsIEBJ7EzLL6RHArkqiuEUSrzSip
lVLj5ACXXcVnoxOV5BlEk0alVLVBXATQPH8PFSrNiQSMKvszbuVVwxvYtex2cP0S
wHB/uB5qaS+XNurDHGMWhwCpFbrrJndsu1karlqlRqyPhn0dSC/Ow0g4RdaSrluh
qHgYzo1ERxh0k32+VTJW4DR+78nCJgpm2wIpqDZ9wzS32lTNId/kNmF0jyFCkaXC
R8FE91Z8eSziLhBfEp0Yo8jkPXzINSRDAWCnorRfcbr1W7QMx9HuPvtcFbSEe7gA
mvIA2dEy+ESXet80WKkB7tboXbZqhGi/BSAQatdrxpikUrJGaHe9cg6k79u+mrJ1
URDumbmmABoY3fAPafNGU4jU/x5WjiyumhC7QK00wxzyNB3nfBz/jO0qEnGPDVXo
Bd9TT1mdxeKkUtxB/YfyWqE1zKUn8jFHqz0pdOYCNrwyxQkMMQauEKR/ek6ZlY+a
iUXs0PFDeT890Eog6WNm+K5jDV1iDW3h6l2r4aBnlmnyPtc1Y0LGAIreuguOB5yP
OWBVmCH/mWZO4dT1DdTedDtQec1TDndBvJO7L0PRf9HS0C8s8QO/e5Cc1z55+2v8
PH89KHcqX2hI6Doi2vlN1EU7/HSJy5/AoC4iVRSKHHs3NMzPi44XEkzSd82bZfEt
o6F2W/odtaU0o0g5LG+A9m0sudhICxI6ptHuoQtJdixxyiDYnM8jE1rmWD9Q6Y1Z
eWqJbyoUi0awI471+E7ls/YtZUM/LxHYHyeojjrDX3+7qzL4ILkLwNTevL3DT7Y1
x5wn89aK/+g1nH3w0w+OSTzuyQjniYtklMQ5ZKK+IkIqHjFbjyfRmcXMHqYqN6UZ
MkhT50dNNQbE2jCbTuBdwCewXUj6KfzosSSfxzIQ+UjK+gdQINg7CWnI4aumea5P
2y/yjEjoNfHM98N+aXo+f1h+tcgBk0iIA9UusbrbSgxbymmknZpdHfo0MixcS0w3
FKRps0DszS1kqnJi5P/MwqCcjToZNQk+jEM3ITPjUBRuGw8qEpY7ddw4x9LBBI3q
N09IYmx1XZOY564MtLQ01wb8Qzz7/yblLYZTh8CddtYGiw+uUyM1xUEGPUfrgVJW
b7pzhSx1ogXZ0woIQLAmgS/FO/hi8yF7PewBhSh/IYvfc0ysugN4DorDxrr0xi8Q
5duAZnKhsRfBOsM+WUYMnUaGIvnH0LMM3Iun1Rxe7ew3aQqbuVcj7DEM7b/f9Nkl
Ah32NEHpDqso7uS9V6Nl3MKF9efqPGndcQJYYYke8vRXRQtbUeqCXNsMFD8yk2Gk
Ctbdqyve2W3iuzEzDIXYrcCbSSS5YtIvKCvb7wWIWuAKRaQmLv8O9oMYJCSVibAd
mZclzrWEJdxF9++XfVO5uWYbVCK5qQvPFpoZOn3sPVPXElvbmeO+f9tiJlJrrrbs
6841PRyWohApBbmw54TlRVtiX92yQr44ketl/m+QXL18i3+nDTeYEoYkzvHXOb+7
mx/DDTYu3feAqIXfP10DcrrvdxKvAiTAAWZqtf+M6LcK7bxklnbrLFXV1AswKEZK
kAs2Kq7OKVSd8ZhV7WX2xPTFyqZSthQkdvd5Gpn1X5BM0JwfQuiVg9CDZ/fDo858
EMlle6talqmhfl8A6gBWacH1sXOaOLOmPHZPKwNEy7GrZTQVdx7s4iey1mCtPHL4
1Beh3c2oL7v9zEsD18c1JwXx5Q13nPitgioOxKP3M+xt7fQuN5X5sky8aiSWn3JG
8uDdmL3KhH470JT7hG/Q9ECE7i8YZOyeJ9DGpgOb97Z0x9CVhgA+R56Uq5UnR+Es
cwGIvkE134axtTIUwgYWKhP1ptQu8BBNgRGME5/0kwhFgbJXlPNibD/lWSWV4oTn
or8lSHwCku/MZwf2ffKqK/bkNoqoytwo/9eWRn+M96tFEbjnS9QdkakKJp+m4SHS
FpGTE/Yn5eqKrCzC3kSiTOnLQO7vJof489rxiYPhCawMroUq58sR/U3xA14JIb/u
43jiLv4wuNbHY6VqZDN1b1R9npPjdJaMj4Lr7aZ/5hOMwSDmNm33Euquzc8q20KO
S5caRtsyr7C6dxoaaAkskUGdgXzKy4dTn1NJZ3qVwWP76GP35eIhw4hoK/VMOI/Q
RXfzTNO46dMOTOWRQEK1mIAUlQNHGUxWN8MMpvXHr7AW9dvuJDoJNEG6kG8YTKW4
X9SJMA3QmwxtzMll/qdmFxLDTGWMlA3koun+ZcKP7lznL0433XgQKbOfDxU9gg5H
6VBDwohcnY6XyTcAKyJzIFYG5z6/KAoQBbLI/0nopFydKJtnSJTaaMNmzZRChSZM
RTzgXbwUab6JXWzlpErArNulCubuYg49Ts62zEVBtHBXl8GxNlpm6TGjCkBgDINj
hVBrWV4k6H792FMJGwsap5ItGNWlV/JwCACSV5hri9ep4GDewh92z9AO/TQTuCNm
NBM+uu3bOZZCEHMkFCsUE4KkmtVTYscKLNftuMLoW4PQiX9jEOzkRlVMymS6vok1
WJZ9taX5neGG0uacQCmLsI7/CoHFtNoUbgf/gobGqM6A7nNMFleFyrcVG4LJjyT+
+sSuy0T5+hAxp9kjZiUoW3LOOHGNUpQHAXIfhfpqYUxrW9k+7316QJU0170Ec6U+
uRrEeIGIeT5GxIrkge8GeJyjoNbXKESOf8VhIne+NsB1EqYiu8yKwZvxkO5qWjZ0
mIcb8bz+pHu1mAWZvGQaR75iL5Dgw0HLXJfbwvOkhd1wp1qxDrG88R7/gi3cqIw9
N9jNx/Qi8AGG0xnFATLK3qv7sRlctEJ4sbDyTyd1q0KFU5LV1YPfXd38m93OIMO7
/+xwV5OVSkpEL0yMY02XS7i2ekAIkSey4gCMcAxbe4wder2Zbe4zL8NSQbXnV4Dq
pro6IJZtHTgzAptATfQ9ypbqtjHEnVGrhIffqUQR+h+nDF8/zqXtJXNgAbqs2m+N
Te+lIhDwyaNHPnhdyO9us8Iac7ZJciH/M9judCpMgz8qSf9v2x1e4y0QiTUARNm+
wmGLaPTvB9zXVumoadBidL0n2dHmsYI2fGvpweSx21uhpK8LT0T46B1hV+JyBNtU
gIXN5EaauP6BCU0wP6qo7xECAuZpCe/CUNIDuGV14MEXJj+UWHV9E3LjkNW4MVZM
eYkbiL/kRM6MenU/NUcpkCej4SncIoPT+YTN59zvMbE/2vr1AFZUqKYZJ0lZNJwl
eQTKXW+e78bhsCSWtjArbLpf1CsxosU1S1sjumeDkYl4Cs4QD1wauzqCkAsTWmiP
4Y+wqmY3onbTgNm9z3D3pOmef3wSf46rObFzP8DakxVROrHb+9E1TyXXN3wMgnGE
Y7qpEA5UXHiXvSWG9qUSNoKmZ56PyeLqeSXU/hDlYxvM5qDxGCcTy3kMhmuC1xvM
T8iAJthAYXasV0fVMmKuXLeKm3NxPiQrjG7KXPb2fYnmbqP00bohGzcxsl6XyHgm
ur1XKSC5iPT/KyGb0GbBLRYbeSSTrLJ5fvxxDCzMl46PYv6+URyjyvFkkX9tjcgO
mxrU+WwpEHMEq/y+eJz65vrKHppCWR9W1TpOWwOGXwI55JSgnJS7G8gYY4odLgQ7
Rv+1DxL1rBu0P9DdlRcc8cDSlOygtqtnhF+78WFLquBeMOu6rq7ZIREli3SCairo
7hG+tJq8mPHDzZV/HpTYup0HWHAp9HQSXwwij5gEKnjZjt3sp6L/+7cEqvtA6AIm
JlPjzJUinauEn0TZXWETQuTCnldGzGjvHMy1K4JElNCc/TvpFG3WGkMS6J9ZomfM
caLvad3R9YpyStPji5Bp2MlJ+DDUs/Ymx/y7PJthQLFz1eRcLFyXPhQz7jJtRIYz
v+FyRDNVUqgEUPgYDpxn2WuOFvl3GqPdE7gd3BByM3PeILOnCLp/ZC1rZKlDLoAt
tECJsgH91Jrqu1PG8HWqUsYT3tC8KowEu3C3gmQZQHbncvWro6zgnv9ssh/Cfy+W
HOQmjFj7QLJP2gLPCUdbEIrlI4bp+UwV4FGIzG7Wvr7kLzkP99Fy+ff6BXYit2AA
F9sndEDUzLkTaoEjsGZLIEk/ojHCBAleJUnWjJeHaQvp58w9wN/sk/nSoTwakomP
w8kIgr4Vtwg870Nn65RvF1gJuitc5//RDsXu9G4X2ZlFBcK3UKQ014IP+cT77+PV
j/xvEser4IC/LRnhU8GJy/EDN6O8WRGGrvqXXIGZkyk+WCwhOEzYd2lkDcpM5cm1
3TMFpKu38kTMpWcfTSqFNm/aH1MBowYfQVDlFa2YfjEFKGGSuFwImLOp7XbKbC5Y
k52WzPleShUHh22rOXNFrCRoFJFnXRt6YqyuAKmXGcvQ1a2YAUr6jDbSCHglOMOQ
Oo54aVkhBZv472otALbdJFQDfQtFt4Yw4byK2VFXIJdnHfzd1Z5LXyH2Ch8MaqsQ
f3iptNZEQhDcLNg4+EnA0hY5gBwPnclG2cxUcEeYlEWrj83ZR7B5arWoQT0k9oLh
WstJcR3ZVyp4ECTLHRclcts7epnz8aDZLDOAWAV20IjgFwx7JgiRpoFy7HGgQ6tK
BvUbO10MQRHsD/8CBHdiZrSZU1Ahul5IAmS6wjuM+dOG+e2E6tmbvGhNL2sfIbfr
Lql7djzAnxrfZIsKzUKQpNstHRseCQGbqkqcoodH1kKPLtsLTV7UmNroF8CFO6ua
qtqwfxMuqnWEhyjoIRQaxN1Lt3C18ppOpi2hS/3NhFQQeMj/NQ+e+yRPJHsETYuf
jdHrX0rs9Chn8rfmsDu1kIDffXclZd8UnteRGQOB/cOyL9cyjf7d3CFhV1Ax8hSk
bWXj2hWgo9YIyfN4zHCflkCwOYRwpsOSXB1+6+ciQozD08OURAaozorJ+rf+aW+q
vW8ocM/9Ist1DZ6uyedd870mF5bOL+da4a4DLHSpirSDOkjkHCoXhjM2LZP0CN9D
cCEksb9rmX9Zs7biTc+MTICjVlmqHJ/4BgMYS9p9o3D+OwRWmbRRjTlR5sImYPli
XCZ0v4VtDgjmR3MicSEB8gkwnBAvw9s7HoUjNaLRshxeL189GYZzq1bHUkMX9EDL
jI19j7prPgk6sUjgq5wzkZ79jPgyFM7Tz3RuoUWPUnzIEqs8k9anwnE45KfzvbsC
hvJFni5siNK4D1k4nYhxZPm/22nhh0iIkqvXtv24V6ug/yE9KWhCr4C+6Pazw5Rd
qCgkZKa5nipS9ogPN0E9UM0heIqtauzw1W3S0nhgLM5k9CdRujrDqWrgzSmxzoLM
7d5GJU0jsTqrIxArMJcjO9owUZzQIOOBT4J0LxUsLxdOiqJm5GPbRukUHrgbyGqq
p8SsekljebfSVObKhIZcuc4rI9FIksJ/q49emeIW0pMfYoxqE4FYk7W0tFbXynuj
6gU0A1ix26slicIpowiYG5Y/C+tzJelpDej4pjr57UnyHnv3lDAtjJutRqxiIqpy
OKJKb3+z2+WdpSFEsbAVwaxCk0RW4nkb1xRdXHRZM+2Rwir2Bq0tSRzWOokKoxxh
FHT8FyHoFR4V+T/tw4Wi/0kWH1fEjDJqHYoNCC1bZHyuYik1UdCRxHXpsL+BfJFd
Mlo0Mnplenm+UyI4JsIS98GnL9++g0W9mccy46Ja6YNPx9ObQ04PtsoSZJP7e/Td
NRMYroGJ45mXEgU1aG4ICXGMpTyRH228iaHATvmxrnZ3FbPxx0XyoKyMlNweg69q
IjganlIZBg36zPKZNKF4+XAxufUzis547uJq4w73V3kyaj0mKvc4z+KAIygVRaoc
S+CpvBVX6vqsyNsIRZdTb5T34IULFw6Gv9wFqYTLtgcMjesVw/5Ptt5zvRBOhLlr
rm2EyKKVt3i157udYnZUPXYxGiNZ5HxB2VcrPu62HpHjPDVs5Jk1d9WSJxdySSlu
9lUE+MU+d0utvEqzTClnWbLdE7QQtmgytn6n2z5Q7GqYUc5Qkp90gRo3MiRT2rHX
3UZaRZmFtBCU7B2ux00l+jQmpBok0e1IqMp/9HYM5+Mo2iUBfasyMN5JPz7PXId9
Ctu3g3Vy6gP6FgzzE4egz/oz07iDzkeZc4zi0xvdDTNKFya0HcP77Rf9Tg6/Qpka
5VrifkhktsYT+4z00tjs0arkJLiDr1Kvtn9r6z4FQ4siCo2tg1CXKZ6/jxVvRKQO
U07+uX4MgQL9KmFqgZkbQVdg9OhI1jaJfY+rWX3rJ1Jp+8YCLQinlg83fsgcwLSE
h/yFpVSb52xPUKrcCj9BN1gFOs2fOK7jiITo1BNCepiTRNhK59/bMHkXzdhe/YVg
sL2dsc23/z9ZaHt38s0TkO50GYbYubtlqz5w+xBtQ5CrQHI4eBYnI/CGmYOmHqIA
WsFgOHLkyIwLrBmwdLVLhpoqx6fH+9MI+9yJWLAWtdnlp7gs5BbguNzM4WV62S7u
zYb4ORYhdWvWAkXdXwo2CAUkWXvD5bcHC6K7nPwJUgqK3HANg6NSbdDDdKagloZ6
uQkbl1DSV8pTL6S18wCxQ7DPDyZuwSonxwOV8/g0rtDZupO54ncNNeBfjFpj88bZ
rRbglW8tq8czG7m/3Ur1WCDAfbEmjEaeV+xd7EbmLGsURle0J0A2BU/bL0hWpHGS
trtFv2TuOJRXrftiSYn0cmyhg5Rc2J4EFM+S1HaEGFYqjpBxnRY7aJRsMNd9m+SA
fI1yZmXbmvZrfo4oNxS9ZlwKj9sbHPEU4dtKNIL9Bgzpvc+/WiIe91Yy+XQLXmTD
PsNvYy4tzsJHKjX3kAxFjMp8QjyVAsDPqrguPZon0TJix1g9QQX2FZa4QbSAly8c
kvUrsSF6H2Ty7lGOlE3+KcL06sCiW6kD3i5/wKPftGSJVFxgi9SC3skyny46Mrdk
OsjJpr524JwVK+cnXwN9pEDdMLWVASCBdOKLRoa/9rthT8FDzAK0ki62345yCjoQ
Qsf9XB1D2gHtq8u+28KagGnV+rGnfk4B39mufsvAfgz8cNZmU9U+gb2KD/fpk18E
LUnXsp4mmThSrBHBrdOq4jmZrx1UvIzyzCEkpPVjQRySuH3IhkhxvuSb6270RerW
qCgG5PGP1PXrxnfpIfvur9QLE0HKu1boMbDAMSfZqR3UGX1a9tYjIroAr5l0QeLT
bGb6h9H3q/7fQSw8I/+BL15Kf9jFnNfmeXFkYRMq+cZ75QrsonCRo2pyyPeYOaP6
Rl6FXUi3fI8VcSUT81OoyG/Q7lJYYtyGM/6XoTw6uTILWUqAtjbNekTy2j4sklRL
/GrFAsoN4eMmxhXrix7nltFh86ZRrxvWwVwKjUOKk7G/jhASoB8roABk47rzOCnM
9Dt1Tzyube63ZUHcF+Lq7b9ZmEGkY049smdgrwoQDciW6vNoR0zzMSD0da/F/MUi
GEPN5EOafMHrnd+BYYGxQZA7MIhrKGxBdgKhfmTtl/RFuJ221lPh0hmHNGGCubG5
OgFIoi+vj98Rbtyig1CR3M3LUP0uSXsWUEIYDS7Z+lFuK59d9d+WmP56Ju9vm1IO
d0lthNgR1oNH0Biy2hbgRavtxiYNurtAR+WQr2C12FSfg4xkyipw47Np2dUTt1zz
v/vSIWsHLC8kTZ0Yh47/dyNg1ZYhHeWAJ811DZlZzv3Sl8I3PcG0WJ7t7z7MIqJQ
wqczyBB0EY7i9U6B2sERgUQPozzwHFTnSfa+k+qUniPBf+Lc1BSnKMIpqdq3Q5mN
t4A8gkg6k5cLnUt2ChiXpOd9XcwXYcErgzlTXRup/bW8fL0hVHb8A0C9E0paLC5K
Tgw2GLbwT+ao7tUxijC0Wa+lhkYgoIDl3uRnl3Ib/qmdbr3ZyUS39qfKs9c2ANEN
JRxe0lL+SFDjZbcEyYvk2s1aX7LxXHO5IMsmOmkQK2WDQTZ4dkXMM8CkaHJJZUTw
7OtGTudFBWrFlv6weyfscNiw6e4huKvzR5z6JH1poRr1vFNlo7qws8Nlen3xbHUG
LfhCuVyzA4GFyhv+v8BcCKqnDAp8QFaLKLXz4MAE/IB4Xkev9rlSi5K0nnaMI9qD
rhff5Ssga6ppsiiTpGbV8LIp+UBw2L1nFHi0v89wdEiLLoYma2V3OpKGHYP1y3p3
ulXGB+r2KEhN1siLxcllF0QryjDPVhsNvE5bMfcefu+hHVTSEvhSYZh5Domu2dBf
pTKrFuIFKs508yIQNhmXdLYrMiKsja6jjfSfCCZfa/brWl42wSV3zna25DW8va0l
bI67LYb/Hc/U4z6WLQ2jdHaMuk58aSNQN4p5d5tGtuQfM3KfdGzpPXp8cQvubcvE
Go0sISDbQc8wJ9knrMtr8w+5swVOqxT6vOi8vcvdo8l8jRvhKM/Pc5+3yF1u8ZDy
Y4HAVlAp0EjA+0IBoZzsA+p74jSnXJXOtSTo+EquPwekEEeKqGPcEB1ML1dCDjIH
cwOjVqXhsbdcyCk2+GLeITme79lKOh5jeLG8JJsAwZa+be6gsZHeyrfRxyFBeKqz
+gnUk+JtcyTbELA1S4fl/+FJMonSe5DjTArEBRh9K8z4GbXtB1aHfzgRx6zF4PgG
ERgfAqECbwpN5TdIc4QZ5ktFiVufRqaqy8xLwQNVa1tafsMQucxFSm53uNcHZ3Dn
ce8QVPMkwbV0acpmwViL7nWfTXOxMzmkEcaKBjD9V95u6bkdczpF06wsgD/wDF/n
Oge0CvWguAu+nlYgpgDai9zn/oud2qTEdoknRyMe1HEND83OZsndtr72pyJLRGFZ
wFAPazIO5jNXa4e/skwPz6GjCpLq1DRU+V7AIisHbQUBCMzAuhDfC2A+jYIyBVzh
lgg9qYjGk/tKci13eloAI5fLQA5FSM0gXT7AkQhvuqMzNP04ST8+cZj3EBXsNJXI
uz0zbV1cGS19ruLtBy1cAk3K0DsaDRYuwXX3SDFUiPNBvvAFGdsJCjxz3Ql4YSim
UC1NZsBrIxY1OEDn1u0iHMoLerDUcpVOelTy518khOeCId8QwYJ/1o9C475hDq8L
E/n3l2hcubK97GVC8xRRvxNfq6XFCMXddW1OJYvbtkaZDi0W1J0v213RajGlo6CX
WHs3s48efYbo1YwMED+Zj1e6lpP+7tFiJhl3WiY8CALI5UAkQJvyc88gFSz/7jPF
gxwYex6KqwN5HPoxfuC5xvZrk+vcyikTRoWFP1gSSwVlNEtWioYyZQNhg2SnAee2
Y1JlP82bdE3109PNgA5sUy1ghpFVdk88ZZdjfMjrrOQau7YlOumpnvUWTGlFnWnW
KE/s/ubL6Vg5tut55qdR/zEoY+uN8CS0Lp1JXYTNGJFdIzxdKKTuldK8lliSPZ/Y
o1FB0wHFsMnHvHA+Ta7CuQ7t/M/cV4QZBBVC1/qgmgl2NolRq/EzqFNdiI4nhB/m
qFi549yekQjUvlZiT7zhi34ys2IBdWf+xgz6/SCIj5EUJsYg5SgFF3sPX5OaUkSA
bT1rH71HC5WBbNmSsF/3hU8ClTIYs2LE0Db/7ViN0NYD1wLNXBlE6I2vQwPkl0rP
IArHecBh1oh3SUd2AUtzsVaF4vJ2S+barvnl+gbUn+FiG5gWiBHOPmnTN8/0l/hM
y1WXjBlUhB6M5Ci/uLBuRmJcFlg/BD0eg5KIrRfwzea0hN1X8XWnBoH00+i8Qod3
uF3v6H3c355jU4IgpNWdj8QE5GZAN45T0UPOhluzVTRoxVdQ1UxYg2I6KX862F6l
V+yro9ZOHgcsVYQZ5Ga5Bb6plOWLln2mJrZ9Lis8LQWtAqD1Ck1+Dwb5YdOky/HB
+nR+2HQFGAwsqBqXPcyI8dWF1GtEGCSUCSr/T5uz7UhunRBMLR40jxrfF+g6+dRH
eM2xli/Z3kfEq2hwAKkvq5+QmV8+asQpf1PpiDFNXbgtIyYGJkIB6GKgYjdtE0sB
ar2aF22aCTF6dkm6oA2smnymzE2sHbQ2MMwh36pCOkA/Ffug1j9X4LTpN7DZTnLl
eghlqrKeStUb5/vyWrvmi5zXI1Jcvpdoea3c66wTz4AauwCLWNlCf/19DauFAuZ6
qyU7dAUtI/znOCODPcgl2+ieQceiEJtY59CoWVV3aVcxwyOgvVvB/1mpNFBBfVUa
3mKT89YpyRvOvlgw9gg1SuoNof+Yp/cRLSe3AuSRvIP1cWfdRj8qsycTa9DfYcWo
bekzvYa1HOo/Kp3vOQjntGDFU90JZrVRhs3LvFckmXa6n0A9XW/NFGtHLGtzse7R
4e27qsum0vWCBwAn30eUi+q4VnOZZA+q83+gZNFMHW9IbPGOWIgG4ine658kIydj
3GPSB1emP2xboAODm6i06/RPIr2E3vwI85SuQBVB8lRxKEhCfp/uqIURfaYW1e/r
rMuOI5Rxm/e0tcbFN334xQQKnyb4qWg6lFy6pgFzUe/+KI/ltFYwMEJdRdWeXUx4
1ynXSe1V+Ehm1GPsjSylS8RjAm50eOlIT5+n0Svs0x2slRpPXcWGOaIUMvToJ4qZ
9DdlioUV1YEAMzQo4lFhmiQRbQ6fCGHrfiQjlNf6eHpBFluJil9gn+6T0qjD91pW
diRLEqfKX4Z/cMsJComLzimnjnxbjdqqyI3Yx1wYfuPzZIVM9+ZYcaWIHnqE2Wdf
txztfl4958q1SXEdhcdvyHVSBH8B4dV+dPpQQp/7Lb4LEr5pWUUEPkKbI4v2NH66
UK1Qdrq0o4dygDASi8LECxbCixIxwaIiqHgAkcIlv/5zWpbKGTZM6zwog+5BEoRU
Xk5zdzcFEjrGD8oMzisZPVd5BcbMWtMwriZGnONDrR6FV7kjpw1tLP67Q/Mk8BJd
Iyv8rtyiGEdPElPiwgpe7fsxEotHvydAO47pCnEAmlz5b372iwOufUN7T+VwgXIU
eJ4cE89nM5NP1/YY4XfIMKZENQniJgGZqIwA0bDrfYO8XuXGvrPUvzDB91NOlff/
sT7YH8DXq7UNwrxeu4ybZdbEPvO2ut57Wfec3SAfq8lrNYabDZhn6tmAj1uuQ7bj
XQIw/S/d3yP0exHTIA53vEUq9NywKJKdyZe34EIGO710VuxTQa+3tJoxVoNLhz4j
5YTT0U6BrwaMnYOf7QtYSccQ94LvdklJhQpd5JtwaDOIwmI0Pk+VxLvvu0CDEDIS
kBkTjLHTaoqI8kzrcOgXFsFtOAE9pbsmQth1gHUz8fPl9kusoa+OY5/fRaA0EwIi
W4LXlcs6qh1FnUgzaB+ZmvwfDOyo0BAp/bpect6Lxys04fiwQKwdPUqQZLRsZ1ef
l7jLGXuR9Lk/B4l2SIJ779Zn5fEgN/qbpqVNmddEmLK4rYidb0JnftanPPjj38dO
t83LhbRnt1kfuZ4xJ0JcVmgtMe5LrD7Bs5wNDTp3KAPzee4TqZOltJV1p/OkES/j
ZmJK6emmVqyJjAsUmYfGyokyjKEc1DQf/O4+m+XBXiC3GNHn+m5YOwzW3IgWS8Qp
XU9fRsBgWHtdlsG/Y4h0dOdnKidDrGtcQ1GYoFuol2/zlRxrZK2uFngXqhZVhPxX
mp9Pami2KHzRILbWcSLs83DjxL//oEHVaGwlFTMzUL7BRdKmqd8ahDDAVAZjvhx7
Xga4ABAu3vmeUyNajM6Sxz1q6GIvZDKYOHCXtK1VG+ecX3w4opYC6GZn9uxGY7wx
bma0wO8vs7LCBtQH99thb3NPSqNOrkQENFeRnfKZOj+z9U04RHcNLOLZIJQavZXQ
LcNx1UIE3PJcEHroiOA+dScwgm+bdnsg6wGF0vi49Vyl53Atd8LGbervjOUO9+B/
zkkzc9ttRKpEo35b0/JF3Z9uCugvVolx2R8ERxUoIIEe65BhKEx3m7wSFt7YNPGO
ArZyswtyW6wAPFciMBob2sbNROx8E3O/fPnn/TtFVhCfs+l400S8zFZpUifGLz1K
73CnUJjdFk+BDYfrZEnqKopG9v7lGd3Qyv4qpLCZb72z3lFydi1pyB8FJ2m+AuCe
R0VZmTJsH1CzmVoX8NFlAb8lpnxrXr3OEZTwWL/VNOKGW4n2jz5tNFwqMJacRR4o
yZfWZKtjBDLvtkg56ev2dTtxunycwc9Y6kPCy+SzdQiJMmKFhQpAaDPhcRCcMLQN
i7rwAXwAHXQl5rSPfIBynxG+zwLPA1kJuCcvMDv/NlyUCDJGXgDH/3E2h4wNvDL5
1fovN05AZeeOqJz+OPPj5AOpkh0IO1WS8m3YzXAx5cYmtmevsJhs4PFaoils/NLE
K6CljGrvDmM47FWlItMP/UKXnzK8UIShXVZH4rI8xhPkTnasQwAZLmiTySSxh+ja
ICj3s6CPXw96DEwBotlyJZ+pgiMiEoKn0XKO2BrnayqrO6kV6XvJ43KdalnJJtz/
CZcPX259PXKN4Ux4U7wxm09putyKuPY9ti0bi4fhl8Dyt+cl+2qTB0N8VaKnbhS7
VAl2txwsDgVeRy5OvqrQGr/b2sToljOeg/l3wxCK6bGbHbuSQiR5ASYB9l1EDfJn
66XMq1P+c3sur4q6uPVNHfQIpIz9jm2wSx9p/Xz4NqcvF1Xnx4z4dOL09dhDo8xA
RP/5NTpQLYFAXQQvE4lw3FCQmq6H38YAivOwbWQfXBsiv2lwM/MPSyLK+mPOFRTE
enl0Y3rsvY/K+Zyp3IpR8mvKheoSG+b29WrXJ5zsfEfI/xoD1Hq4fQxDmYaCc66e
GJNhfyV6q64ke/X5801W+jk5RKIBLYodP7c2/x6Fg2yB5MDOoY6oI3F2yKbuxwqa
MU1gvPZMIWaAFV/Kav72/kQ9LULrf408EU+2qE8lUKfj779hddC6pyF0XIGKxqQw
Ul+UBHkp93pr2WAFNaHvNvHPxckbceLjRn2aL1WpXTIrKyIv/ainO3LFmj/2B1Yn
V6C/Rwg3YT5K8Wz6DXH6rKVRpJGWUGJawWDZy+ErmG4ooJo2AAAuCeGqhkxB3w9W
9uHauMnriOCOGhU70tgzuuVGjkDBOIu1RYaBmydsab1rF2o4hz3kGlF92qO801Wx
zCXsLg+JgdNPXQRpDGF6fZ9UdMo7OTwcP/a8wa2HyJNwS3VPm5146QW1t1VS0uZs
7JcyL6ENuYjSB22dqSr9BFx+tvNmIJLDpV5Jbd0TqYPf9wGOCENva5BffdyQveiM
6hmyopKCj+QNElk0lqY2vohiFep7Gp/NnwIqrb5y7DynXywQrl1oa31pm9Lteysn
gYzEX/XV8SFhuhlLyv897lcQ4LaL5xeoEOcqmcQy7AxSSzxr147U3ut5228r8bnK
5fzvYfFv9N3t88HJy08r5c2cSin0xEEL5Q+zo0Xmp6mvFLXhw1lOE7jcoHuLtHjq
cerXPkS+iZBUh4ps3GpiavzJ5vR34ds0GCypsgM+E0gDwYrEDHcNd3hrwucv6MdE
2lxONBa+dkolePvJeJDDc6LPMzNjedeM4vKYVzEAucJPvfTtkG1QpQGh4c1a68sM
a9r01c7pq0S/VRttmdHr0usd/YOrY9Fg6fGeq8UHvpxYqrAFE8QrVsp6wSu6h6ea
`protect end_protected