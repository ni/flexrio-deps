`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
YATj3kULTF7Ty4ORuRfFpnT6YIk4rUPRrM74bVTnc4GjdV8oSnW5PtQkMCLOi558
1V+/wvDfc3y0Z8//ksX8sZm3JZWtrxUppw8c14g9Y7owiwp+JumRtO1zuk5xFbe3
0MMnIxxoTKLhyRJtAxElG8sbx8N21OWDGiOk0Xyd5CqAmk9dcOIbxzMjW/wndBXi
maijUdqS+5KiRCM9+Gsp6k/iEAa2LnYTt4WtjkmDD1P5jZKsiMgFck8WOqLymplZ
ml3TTfn1UlLNm/+zD3SFGP0kABAiUT8NK2xBPQ5UzQ6sMFPd/np8iUZ5u4QLTWOZ
hTrU9OSX7lOvRUo8pJ9vPg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="BzW6NOo8eyBw+CxsNNo4wIDxODIsVe0ft0K5tGuSUZw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
DhjJh9S2BY18dG77XPz3hsiSQ73+w0XqfJhD+f+lIDHHVjOB7CfC8ieNRTexgzn1
5W+qoqOEwenoVQtit9u3XViXJSRJ0wfUC5a9axblRNyD2mUbyfH9+f59nWqGkVOh
ieHxkA/DPprM70F3APxk51m7/gNSLICSvbONgLGndWc=
`protect rights_digest_method = "sha256"
`protect end_toolblock="L7NTNW/5Dqy+2kJZXKczEa3js87UJ8H00YWI+92sDHA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 57664 )
`protect data_block
6eHODtGLmq6ccbB074dgNWpdzW45i5jL0Nzx5wwM+RA0eeOHXxEV143NNyQGmZjT
bzHAi/6AyRCB4X9z0c4MjyrZE8GF4crbMH4T59xFHqVrQ4zXCea5w0kG5yvHgpKo
nHE3X6HApEb/JkTBPQNZxJIJV3EzMk5ZeoLhBtOMEpw4YYNZ1VZ1itxtQ0hT67b3
et7WkFdsKzm3cq9gxmvxfzGbRpSL94Hi+pLzCbTIYGbe9CNJ3qO31FJ143KaKz5K
T9v5iJJErcsy0gR9kfhxzNhNbX9B4ZNI0BG2153EtwFG9X6WavYQOcvuBejPbOPS
cAnohrF+k6IHmHm8ASY3Go099dIVx5GcFsTgFCohaKDUF7kcMNw6LgcNf2JLMSaS
Ai42eKfOV0gY7DogtFckyM0B/rYxEL1PTs+8m2gJOlO+cwVESNE3beCUrkorkF/c
jtJYozA4fWRuOfknSrOh1MAVfzvbqfqnWfRVcF7UbXOxHGK/2EAvbe/m2f00TW/8
030L5LCOksQf1wjG+lYix+siCpF8USMQQGw0yxCOXjHN8vP1RKSqz0ZyoyoypRW4
MzFIxIWJNlDU3k0+bt28DTG0+cHsCzl4lTXaJNKJ1cUtnhOmqLC3gSZGz0pQvUPE
VXYZ4E9RwEDZhkpp+F7rPhYN7lvvIbLdBt66+X9SkQQ58uQ9YUch/kaeL/ANgjGN
HHj//d22xUEZL5BCr6UaW+G396wvjJ40/Vp2YzAekBfj86ypYWKt/R2RIC8k4/hH
wdFCRUzq6G5VkBG6l7ydTatJPjWly4bR4Byf3ku0I6YT3O3aQJYsVVYs+i6pvDrn
IMyPlwbOpXTDRJ36+JmTAHjxCugAbUEf5gkK6106nTLxxzdIkkLZYk7EMFLMIMWC
F5EDfweNh6srD0DoQPeCysH/74aB7P4CRlnclXsSwlBAU7pfR+0udm4j5QMcqaX0
QAH0Z76vGYlndGQWxbCF2McOfE69JTOEu8PWJ6jId242QWQ0ix5V8CMegU7HBWsT
TBDw3nnJw05Xz8t/9l2vW4WWRsYRD7olBOEXn7EQj0oE+qEAwiBk5WQarnvR2ARs
XZbOt8CdIzbDVvubFYRfLDnjnknjW+mk10eoQXIzxZAiZp8dV5z/Ir18+KeuEziJ
WRosmyfbPp4QjRjaRiYPjgpUJvD3E5pB/eVs3bDY3tskPGnDRZKyJDv3vtVD+mHI
21pZoseSzGG7G4hnvYm3IDMGINoLZCD85dyMVvTenPlplZ7GrnWVQUVJkWKrrsWt
V/yHfPlcAOMUL2Y2DpQIHxXJ616tzndFb/k3JYyjOVToI6gLg3/VUeqvS+mPN+sw
zQE+yMoi0QXYsamrf6nr/Ij865lrG++F3XP5ocbnl6Wei/HFIVA89LQ8LA8XgCec
cxDt7u+JXDt9hEMaQFALXRxIcMrq04OBPaDOZGHrzsWe1RTjsszTXQeaqyexsuhJ
JwBlr2xjF/ykHU19LmnSlgPvyucyC1H/Av00gSIeu6MYFDbT879AwSNisIAOnpNu
aR7n6fREhQ+rLoaqeDbpp3xSiaAeKTRX7N9w6Nb7ZtLrbSpSvgifev4mHXxoVPnJ
TIDMI8FF0L3CwImTeNUqauhWoPGHsijm7JEN5BYULvaYYcNJGI+oEjdaAe8QJ9+M
Eus3hZUyki/Ecae2MJlG5FA9zawOFt8ZyDotx/yArv7mPpnX9rvRD2T48vkRXq/Q
4/CDpg6AKSMWF658iUaRK6OGAjZLzbbgQJLayAAxiaVukxrYFh7QTE0dHFH/RSMT
JYx8prMVycVMUgtPmJddhYm1LRi8Ao/r5SVNfngo+t5PDpVVDUJohrqVPVhc6V4h
sSOvPTeVO7GqZlTx4HGS654s0Horswz39f7EbizP4XS0HW7/Mn2dQ/0TKa0+/4/G
R5H47szipbHJzShIODWPj+5DSy1ao5TT1b0aUvRR+PBHdIf5wOHx2BPUaEIiggzl
StHL+fUgkor2wHIaqVcfQ6iA2WxbAWthSSVSU5CP2fGjVIQ4Me6bptoB2KdCKJ+Q
LrGdur5yVSKxHRXS2atLOEinm2SkOW8Dbjo/OYZfllMWhwvfUVsMi12jVDXaWgei
6G1N4zocA6kDdVVl7TUyzoMAkzOYLR3p+GzbKOF9sNdOZ0j9VDd9LpqqcMxF2RGg
cr4GPUAw7Sj070vUggA26rcsHeludf1ubXlbq15nIXpkEJGn5TObRqXOSNGWgTvs
yox2lwLYT2e0sHOxBR2hxJshZLNzKeZ9QLDYFJWPxo7e/LaD55rzecxVTQNL4o8H
djN5SLQ7Zp4OAUJntFy/FwixmG8xsrXVpBxIThAoiiHt8SgwoswH4yI63ep6dr4x
PLllAwrL81JALIm0itKgjZXgPE9RUkQK4l2fQoR77p+wENCHdvOFbFZ4cyAu2lCJ
grC9C27Qm955oKFOCaPEVI8TpYj2HpUY2ORHQMJrpA6JKXhw+fo5z8smFEhBtuIX
TtSlPRTRzd9wG7cp8/+GlyQgMx+JqC0AqEe9InFQvuqqpx/yWxA1hyP9uNgvGUOA
54aRW5M3nfkzzKpzQBAC/uFGx/BaCLfXLKPCNFqh1MN4RPaw5QyLhAK6I5DxvHtH
HOOLGLJ0USkH1GvvQbUemt5e9H8S8P2KCW+DrRqso1iKexuWlBj6utcH0LaMnEIQ
KGGkUvzp7fi+Bzk1Zi7J9uIKzTMEF/vjDBMh0pjlyZaPt1fgMklAPU+LV1nb8efN
qucxF3LJbZ9Th+MECraGGCQ7R65Wl5i68laVfiA7fci/Sw4ReVMXYy3kUopuGiI+
Rhq3mUDzWdswhs8IRgfzko1NgCth3im8NJwv1s6qZaoUoTGjPf9OgHrdjYS16IgH
HsJZHMo72Gg34LoGf98ALgmT7lO0rHlRqypJcRWsBAqfzpUKt3mOCVer5NcO6w97
j9EuXh8B1Ia4yCaXsIjA9jxNKTuP13oy26yiht1uHg3UjZxFwVnyigFcDF7Nc9E0
D2ko4yNaeF9sw7hw3TWLZVJhzpwikCV8ku2YjudcS2tIFxGDoIPwtkJ36ZsaajD2
HuYiKqIsOcL1d8DNzdUj1E31g8m39W56xrAfUv19kWEspn+9Dn1+7fvYuymlMrrq
wZrfkZeIZjIWDzPFXuzgmtrxJtR23qipjtozDJfqFGSmIXD65JBKWpQ36kB+n/5E
DEJ93jPHp/Bis1h9ocFYwh2CZi/7vc3kYaMSI3e3LvleKpwRPHkuFMPRWOhTZdRK
YP4TzWQbCqvt4yrUvK/QQjAXALgwbHf9eRxxL6m54URLlwjW2+9bY3ZAD7+DHGv+
lYkVCDwxaykdzz9eeEFc024Dig1iyQSvvi3Y+6txzL5cRKxuJtwEUl4xcUKx3rT6
TvytoWVCpSIJKfGe9fCsQatCHfPAWK2+LQpQ83z3cmWOkNA913SyxMUXk4wGmSYm
SO09u2Q7jZlg0AbX6G93cZ97DmadmSOK8ZRH2cL0TUCpBI+B/e64c+gcRgSvoGKK
Tk4VwtBYOl39FwsQa7SVVK7L966IAIezztV0qkBNPncDJzZWJ+lLFAzU+2f/3ADk
Qiweb1k79S0ppNn0d2k22P22xb4cXZixdVHcXO4CedWkxulRP+4+q3kcAO4+DJAm
ZtSpgADpYFUgvoeMa6DsjlHJexoF4IjXK5odP7w4L6F5PpFRdnLjCSunXqoxA/A5
kZr1LnPK13RAFNLwjZ5F74sRQ2cN+7wTTvsvYUeU9mQCv/tHdMrwJGWUBgtJfBty
T+0L9iFGKjQvUMoM27CDkhaY1rdJEgG+oo6ym9EfWL6nEj62ib3XVEZC2V8Q+c2l
+ERBwZ8o+oDYOPaFLQ7MtY95kZaz/4oeRCcGXPdo5iNPAz1zbRGDfUTyXcjCJ0hM
c1yeExDoNPxZOgFXpc1f5/uniHVPcr43WDf85Hn63vUKmbFPhJnL4WMFzFEM0uYw
WxYbJ6u4e3XVmigVB2bxe7LxzYEDm+zNb3AKq09sJu89dnN76F0mmTJJ66RHiX/e
+gR1zK62XCiAlZpr/7WKfeCsjH55PYyo3/UMt9UBM3c1bI6gGzH0PTgqiqpheada
ZV0tSBkYaYwILafc04JsyWGmF4XXVsHxl9lJ6YoRDrJbl7YEBD0gs8qMFMYuVs7t
wSPPmEg85LSJLFG/OLzmUExicQayJOziuTZbD+JOTQ88ZZb1DEqLbFmV5SgHhgVH
Iq5GfA7seWWGIrsHnwNUMiZY2x0ajU84XTj/ZhWcsI1lePrGqbRMJ31W+gpZ7WYy
6A/ovAXQiKPPpX8/ioAWZedn2Hnydu3Kclt6QoBkhl3REIJYhfqCPFTfiID4FWQF
/HPS+2O52dNeyqLG3lAh8fgMcFRLZr4HsBjRpgp1Ykg2utW6rc9rHTXlcxXCSWCJ
W/FdyF55mBqW4sAVNkd3EnmsRkboGpJSetDdFuWELWjdrc+FTaZZ3xbDYIpm+b3K
L8PdXGWS6Qea8su0rB9qVN9G3JmTw5h3dLd0lmqSajIeDF87oMc9U05ehULLNsKw
b+wd6TYHsWHbODjEYS41lD+DbWeF2h/6gnSDVtgp4TN2/NWLNeHssTcw2K9IZrQ+
hCg5j0Eqlkpng0WmixkTRdf33WNanS5LqQO+Vv+kLLaHFsL+TJIGp6xgWYPC84ve
LEsWhmCMZOAp3AfR2Rz4VsxASq4tpff99MKpccdfeR0fDiLP/kDB0InfuGAnEzJk
AxxvNfEOn4b1G9NQ85UF5vV8I4zx8vBWC/Q+R3pjOjpTwuky4VN5IjrT0fTI20vh
+g5aprzzCuIoqj2RcPkXQhTBHgmlVhxz06lS8lRHC2/dxzLG5adKScrPPgQDEiWL
op8svZ7O+oECFDCz78B32pcv4Ami3bAbtGWaZFp9L49XNkv6cJ72cs8bKbhZEZCQ
PDZ/LUGSKbFOBRSc9+43xES/o2LdWnv4qhrBOrOQ42l9LaFClIWGWtwYWrGaA9yy
2fPsJmm68Mvo3oBmjg55ewYrydqGHCc1vq4n8IhQyZViBJ6z/M+J8Al1wsI9hB4C
9oyqLLbIPMpzwbyVGyn9eKPlSJjt1mDTfiAZsiZELHrtQgLlqCQ/j9sTfN4Ha9f5
IQecHg090tq+hejTt2u0X1Vem81KujuqDV3+ygImjkhxF5RETifKvIIdhJ27ayRs
J22tQ5qIzBRVX3Ew+8my/vpwe+kF1m8ux4vuIw6+PtezomObZqVzKIp4CrbIP8Ku
xUEix7TEBAeREZWAWIQTlkrGyWsJ2kYpiePjKvkDfh/ovFkMMncXSmxCnwdhKEM5
4dKH7KgJnXZSbehoRJNN3l+AIWD+EYc83NsSS4A1w/nYReN40cnM0rRjMLIlossV
M4ErPjJa1PQeMSAg7MNYFKiGSu+hpqp7cc5tNG4arBRYIRSMbjK3E3x4M6MnV+oz
gJaPKkAiPJIlzxsuBSQwcX8mij05ZwPlslgcNiLs+Tq+KuYQpJyvuvEM+phLQUgT
5q3savA/BarC10A+3t7hvI7Gd83lhSFD089M7/XT9+jesg9LiaxHftkETufTrwaM
RHRF/T+SKFflhZT20Ry53ZJxCK3QMy3CairQ6E2xyp2yyvVyHT5JDxMUz8qNCcaF
VrK7gUwuQ7xRIXlfmDwPc8nBj0gAKsR6biPRwsnlBL4E2fEBSFaNXuouFvlnHcbY
LEU0M9EDWF0OuZ1WxYJpx9uXjkGZXnRPLWviH91WxpAF1XoStrIrBAWmqTl5aFka
5eDZREv5jyUpItX3naSS+yPS0NSCThGaBDEgGAvP+uPdSWugtp5SxYk6liw78C6G
jPOyZgUvY8SMxabOx6Pfvm71msHKsDI5fB4wi0I7E0CD29y5TA2NlPy7JNGORo0Y
gxfBMU0Wk5TP58wGTKHrh5k45KaiDYyUk6ZFko63CbvzJZI5kJF0SufU08iO0Nou
fMwBD4rsUu4VHu7acE8v3uoKfQA1Lpltc1rpyLHISv3CeTK9MrctL8zzEXB0H2YJ
6747gqqIIrmxbgUvsin9nt3p3+Mv+9NJwKWEob7hyU2bXh9/n2YiomhVJ+cMICth
DxsHMg8hnbgQUVBKHKfQoI5uk7BSRxeLw+PkXQmTc2RYD4sWrSOLoAJSUI1RNrkD
IoEXP4wdMzb5iE2qo2dwGANgXD7j+LG2yY0cN5RzTsh7I9lhurn1cym3im4AbaQc
/ZJIMg1L6S+9Da+NfZrCoPk9yNldA71nFIpau1GFlZB2SZzabGXK7xXN7kVhyD7K
K+Co0I+8y/kTm08GojMDwWttCl8GizfOENBgcF6s6YklrIdF7DjFEymeVSsbyJ1I
C/nn/ZvEJdeVV83HXEVuNyfiucBUI7JPJqVLGCzZZs7k7zd8tDXwB/4aGdf5rNzr
xvo2952l1k46s3/B/hhhWjw2nfrDFYs8C4V6l1V4YKmMxMzKXT/jGxUIqaAF96de
lH2K7leFlc9u76tWVpMxS4JayLpclPXO1KZ3h3KLKFA+vZIqblyn9eHQ4khptVQk
hQ0+gAS5x74EDS+ZMtvsf/CVSHQAw7szhGdSIdMtg/WJExNT/v6AZRXgznx1WssL
lPm6+n0MtSbSXtY3lLswgvwmH4DSTzj7epWL+Q/xRmrjJx/hvEL1mYbiXgf/K9r4
J9D9EbolKMEGKP0ufK/Up7JZRVl9fZoq+7PRESox9Wy7GWhinqmluSgOP3CLQ2+U
BFUnfYXoJGx5sfVxD4OYC/a9W3BhuFaE+O1Q4DM/KEnDpgHGj2yIHxuqtLqiZj0S
ge4wZjnklFp0sMexRrJ9skc2C5e5YSnVfCGXNhMUbDisB554SfQ7Jf47Uk0Nz6Fn
Ymvqcy3Hau3vV+CHk1O/SigrSKoR0ywEBDGlzSVVjAS/y/O0yi0nIYk8xTnz1YS4
IDHb1surY1A+TW4UTviPEVQeDefUqbI1heW7lGLZ+hklwOU6hLlEwd4SM+zvki93
IRb9W1KoFYMsLdCKFw3YHfzW6uc2itt1oVWvGdPZ4UWEyTcASD/h8LbucHWFvjuk
HwmNZjZzdzl+RNK97ZymoTRJOJvlFPgg9oAIh0usWgR5WGlIxv/K99+PZRtGYnQi
3UVs53Wb2essbUnwxaP92D61FuGa9pNm9HzrUKFyD8o62LJgQ92ewnQTkse2gsOd
dtGw6lXfFj8c8CSRofdHIe0I+9QZdNeOVbG/LlkPyBzM1IIxbjiiRlUVBd4dUEu1
FQu2nwRAfM6qNH2IydJ0cGmyPeKOClvI1tee8L8JLzcpZ9pRxV0kr0B/bEhQ6y5c
liRcT86JGl0opXDGVkKdXF8ofsbEFF3faN2PRXfLaFenbuUv7MROcxQY5RsoOXd5
UnT8GzIIy7GnksGjFgH03zRQlJyC8cFoXuzYRw9dSgCkC/7ysWPCXy3tZ700DG+D
4ElLBlyvCzdzfXZYXMoTf0wOWqnGY4pJ495UnKqhw/msrxcDSXbtEQQPFRrWcQrm
1fefTgeQPC0UmzpYbeXK+/87ofqyuNwv8FRykfRGQNGosp8jrAaJGL1yJ0QQUFM6
bLS0UCIga8BNWy94IXX8zHcZlsx6n1d4sZ3cvz1UmKl9+Td+kBNOmiywp7xJq05C
Y1lQrZYE4ebd8/6RM5ybK8xAajnJZMidf9q+6+j7Ytto2BXhRqerXu7AL9oIEO+g
cVhLTOOWiZuS5U67iRanZBGCgvHZOvJaizMmyM3ADbyUsmSj75fHEP0+C9wqYZOw
yC4m8rYlGsQaXH9DI8mq/lkElXpL8HJaNL+DvZYiIMS6eHWOxUpuLaBy4HD+HdlU
puG2xPnZSY2bHWrHsu6/t36nMH0NR2WnBATctSTcnmaI+VCTJvWIos/1i0iNFSrU
adwOjpjRyUxBP17Gzi2BeS9D8EBBLWZxS9rBAPa0OosYLiamhZGsBAK/uSyDEDUI
ZZE4VMkbdzE1eVhl/1eKpMMJctG/0X6bqBDnNWxormcMh3dzq09h/fgPKZsAJzoI
xqOWxEl0ApsC7qpI4qlGuiZyYSze0+ssuAD2i1rhEH5Onbv4H8cBi/XQBRstOw2Z
+G/u2ydl+RvERIJeDOi5/dwn+V5zZGEqM1bGpYf+PHvWPAB8CQnWKCtDF8h0cj7Z
O09GOivNW2+In4lrttIifkj613A2WsUMAxp55xO4LLd6iKXRqWfqlw/sGuL0wiFk
DYVdLF7jk4mSbcde2qhQllHB9I32fv71AZI0X9DSKaWPW36+U4MBwKUOp/JnH99z
E+pP+89SNxvP2Be1HF2OoRiYo4AMIyQe4nShH5pe01DZ71JASvEzbO7HgXB2tySr
RfHS5T4EAWXFdUtTy6fJE5/PbEeZedb17WP35i+scuHdcHQMNUbbce54rdZSlnoC
i75OBpuNVPADow4ory/XRCAE4GI/PQQqVcUtoCEJ78Qxjy7HaPo7INRBlXLYLxP4
U5LzgLjdTml+pN+xs7q1c4tUnwirG/7l+8APYvM9KjQEa1oabbVjHNRgnPJgzbe8
Id3bbgECwjQIScZY7YpURQv5/YikRKXnDIshudC7ota9h1S6BQ0M+7wIzZc7LbDq
uUjhysemZCFdTiBdBfR4lnoytB8/dKKmxFuEqKzuyCDH3em105Z1yrhzzhFyL1Cr
ocdj+ge7nNZFvOb50cpqnCmYM5NIac7ywfx6unO0aSfuOURaPF9qtxjPoYVgbT0F
VpwZg7yDxj+LQfNzNuV1TXBDXJCcTMhqg9ZQV1yqqfiOk38GjTBUDZqpDdSYTbry
PgQLGBsw9jEU+4f3DurVKQleaxckTgTMnP3jCUlpd/bh0UXmZt2wjriATOo3vdqT
nD9m8sNXR69Kw1fVTVzViXqwvd5jcvE1C8654m/oyn0paiYWfu1MFV96iOA02a4K
TZa2ziS/OzHQHWI5siVfhAoc1aJu2lIJ9q6ZRQywx8wvfBTDyNXm8EiHYrXFt5u9
CNI+KSJg/4eRmp9sw8FTBAoT2bdIL5DZEtExjA/6rxwZ2JyclJzgBku47K8G4xff
qSQe2RFBOhFB08bbcHL0gzms/SWdgl44jfnU5BDo7GwU2MtCBIcfq9HUfR9moBLT
h3E3SH4seLMpbUXRTPcAvI3ytETtVQeuU97AJrLyl9Q0w4GAtiwAl0bc72FrIf0c
Jg5KzT5/Gr51KdLvtAmbtRUXpQGW5qS6tWiMT7pJZapUk9baI4vigHyVB4E2ihpo
R+QoaO2jkmXsa2UyFAo6ajFs783bSaob5pr/Xk+s/caPqZ391i/xEIQ3jqbQVht7
H+XTL1dJlKHKA+GYdZb9RHmPF/ze7sg0rZpWI7JzJWecdTMLgDEhTPcPmtrHif+X
5AGzoEuDQcV6QFCqAhFgpkjbNOXQ03tCrTPScxXKFFzV7dm7mFLdMRd238ExdVUH
fdqBvf7a4WtReQRd/Kevgg5JK7bbh4L05oKflS3D056Yy5IdLf6e883l02w643Vi
iNZhyoPKrR+UknQzxkS+aTjQNrO1anBnWG5e1CVsZjHJwezDneZvDto32DlmaQhD
j3V+GlILaI8Y7oFtildWuQpUmyul0AH+AnxwpV7Uh1DpDpMhLdvaJQuwDX5QwToZ
aKQcOREN2c6kCD188bAe/nlq62qv8dA9FvnZZK6RBjVLA4W/bnnnf1benCTT9ssL
OkEvEz8t+zYf1l4wYNGpvhMoGlBTpkTArqCwK6xbq487UIhAQ0op+j16P9R8zuWE
l5wYDsdD/+NXxVtCdjz1talKdYN0ExIVGxTJ0zWacydPGF2fINrltyeUTh+ha0aG
Ob1Yx2tVr/mvEu5bZXu0eqX/6hwG3QhT9Ccxy3LqsCb3m1+vy6mLGbwCi9ubIKMf
Ua7RXVcvGnU+QbYek+KoCNq1/ClEp3pc/Lss6atnx519iNU7FVq9TRCCHT39kq3d
iiz7iaGVHoix/Mp7Wf3vvRd6X3AHN+FEqNFpCHcoiau+iktm8thIBPHx8Zj1a/xf
l80mDoB6yAhbTzmKYRAf0C5Uf1hN8hwzTdESVHgu1ObBbYeWGHFsei+4Cympu14g
wn7vihFIFtKq9BN9CFAvwsUqLISn8eP2Iu4a1d3emo/dKCUClf62ywbSlk9UkWeZ
lNbCw6ftdhg3zewxCKpthQLh9S+Cc5huwr59POQN7SNBaSkuKyROQjiDua5HTaJh
wddlAvQMUn816cyFK1tUlhW6dcq5ywjWLt5VnwQ60SE4fr9EVckJW20gNMQFFs2q
KPDy4bG8/8i4cKiR5kjA32oC1tKIs6yt2impq+53LtKkfb2rbxfXIaFGCdtU0sBp
/0qzKVKa11+zLTBvbZiCUpfvGuCLP0SgcKNxzDJh8NvIs9feQ80al8p0PkJgKQbc
iDNxbIFVnLVUQQ2TcXNLSs5+0oPykzS6DkJgJpyDzHauAMydEMJO1cgO4X6RkdvD
7mbBnNr84yBa8ZKI/iqg2dxRvCRk1+0pQT2B/bSVPik2rFPXv5tAjN4+TUb5JVHg
pP94n3l4hJwmj0EOCPtx3pcGM115xjt8TzNLfJscJyIMaPMfjOPb4L/66uoEt7wM
KMTl2NS1xXy7a74nH+KVHZnLP5au+giJLFUWXdYr103Za37O/eI/nwGJz1Cru9/d
nfhM0UsIy8S3l3/IqznlLAbLKxZfaingpHTjBarrP9kptu+LcfbGcRx3cW18Xj8E
CwWu6ZX0ZfnSHfLfnzXwcbEApXN9yhC1+QzjZzuzkr435swxyu8rUAUXrb5AMXE0
zLpItTx5YxtKSERVbnrKvikbevM5PEnsPfkSPLjIYqTUPJwzGGqh7odR+KiYSYZI
ah+mIdJ+aSmMei13pSrAw7mpmrOR1LOCGSkxSOe/11n7WmpdSEt2celGlvs+nM2x
jlG/3tigwNxHHNfj/zyIeuaZNntpf8pCEaxjkVp4VEKiaUIPjtvysgv/Bbx+8tVn
P83Cv0HQI9tLnTVhprj2kpb5mQd1Xzk9N3x5ZiOJlyyfFvApupXmYuyNS6VmwKkk
QJYOSak1q8zWkmmGqJxsWsrwQMtLKZEChTGof2lqnZn/PpO+DzY6MKOPDw3oM5lH
nxVpzHXmvPp+L8rcrSXhg+TahakdnbzyrcLsBRptEkheuSYamZTruM+z/yqvNcNG
4VHCve0vrpwc8fIaWc5V4RNU3j++kLn/fd/d9wsjO8IQ3B0Pfov+Eq6anXabPZHz
cZSE0wCASObXMTXs3bqQPaZ5UfK6B6bVKr4GQslz7O80syh4zAG06QxOg6WN6yZ0
cUR/wYgWx5OIh7ouNJe8bfC11EpP9/Z98YauaPnP49K5lsOkJ6b3FrqaF5xL+MxD
a18v6eG+L3+GSJ2eL33DiBZX3GJQGQJYT+BnYUwhzYFGKeolDQ+aPd1kWNV8/Eng
SYTZI0yub7uzuOCRmjV2DphsFmvvibtXGW+3H0rRtd1K+GfUHXGsNSdi58gCYXda
816u/h++x3y5/4Gs8jJzWY1ZwvJDfbZk8slrCkPDAR8Oh+3kDCX8vOPQqY5afvRU
pj+4+FzyWTDF5vdrqei2ZJ3RfVYOapczHOLDJf0zFgr2djGWlF96J4CfKwCxMaB1
IcgRTzLyWOk68hFia5J75hkvw22THMb/H2Vrt9gNtBN2YVyV02P441Ed4VINIuQ9
76HOZZsPvLgR/RJ+Vn/cZTgc4VDhIOXjmTFfUzTeO4U4SeNSdENG5Sk2YF+IxYla
S7W/7r82wBJOaOd/IhAI+RKBMONBsn3xuodhn5jK85QXKpMktJaPxw7BcfYOexWR
lw8A6TNAJQhA6edqbOKtS/BjLr3opuNWUQ1pwvq4/JLtB+Aa2JzudjOgkLAWlERb
YLoBzQ0iJuK44hh7vLFvIucP3lg3vDkg3lq1PZiB5oFsrh5EaQj3xSQ0I6obi6Uv
MpX1LLQtONxo4G8OhgZg8w/UNUFhWolJ5awXZaW6ZMn2mPgZ3kX2EzoJ9Yr1piPG
+NrsfYdzxsJ3yQzYXaFoQmeWyA9R7vfNu1YBiUfJMIryPtY0EBv+VrvpdMxO2G9e
jg7Ho5yfyG1rJjpcmV6McirUVSykFJ573ntasNa/wUnmU3R79nutOGCUM33bDUvk
IwdugsbgaRS006g1jrmq1P0XUS3OK4XlIYyN+xXcFepfDoDvLS5r1x29nfc2lBAb
pDN055tCnjEwwzplq3XeqWZMh2yFQgwc28NguWqDluj8CzMb++i6J9GgUAaEUw4d
omupRPnr4/upVJp1Cga0QM3c4Uf2h+3vWVsp6+2GKswcapTIJ5gDHeny815mQ4a2
7ubDUQJxRwLmU2KzIfq54eL1HL+D56bBrhyWuzLHFddhp2NAfHOhG07lMFQ+ntqu
5bwtkcBPqABjFuETtfSv93lBm1K361OMMrzLIT3HdM9tW6d/A+X9P3WU5jRM8z4+
81XY1z/mCdEhVm+CT6t2QXRkRpy4cTR67Yb0UahhtDkLQicL+cQG9bN9gPF4Bfyu
cEIFqNlkCI7aSonwTxfn0/syxWDQpbIsjmSA0/OlaEJf4Vm6V7Y1RCpgN4PvpHeM
RqGUfxUkxlae+BkzXzqvu/KhwdAPvVRkhz2f5W45pHAtVQZd+Y8qaSR1TDe5qY3t
hFP+Cg7XghhzdRoAJIclrjd/oDqRb7UuLRTpvEl6lZqzxtyDXY6Pg/B1MrBoOcQ5
kr0f7ZgCIhBURAgK3CnsnQdmXCsGcADFMG/z7rGP2a0VwaKxqFzVZf9q990ZDPyi
7XlBVmsugJgup/7QD4FBrG/ADnV9/LUIMv8sRXKd0uAh8V87eYf0dlEIMBL5rey6
fmkEIlBP5Ty4Ef0zHJundGSZ6k1GD5zY4mtePMzKklZEEN+kHRfNQqMdjOjAlx9Z
UtkNmpUGTePDvkd33Tl2G014jyXG1B2BLzPikAonclfVpgwLPKiMT67cGut/kYHt
+z/LsH6l2bjKu0jKvP3pmwRmpsglEBk8SAPeulk/+H5/tb33zYtd+AimEDw7899j
hXZmMwJqS9GTi5gFDvmn8kQJhaE6nGMY2W5CpRQya2hQve9r0P0SNf2YXGepUzJ4
wiXfY8/gAjy9tfx8Xl0wNyLXOi8dWw20q83aKDApxApl0I/WDvrjrEZMj+qZYz70
sfRLpXGPHZqXIjNU1FEN23Nol1BBuiD1zOorlUxYZ2rBNfAbZGSydlS7DNZxWTol
phwqLot8FCaFUfCSkCTFJFx3AVRVzdfIAfSqXUSFU6KQhqdeoqu4mwoPkhnCdYxd
gBH1anmgcxmkz8qpYTwfK+SZxk2VGy0faJo2Zc5W03YBTj3pBfrUFYKi+uZmU/wM
kbLbZhEg/NECgwnkuhU5d4N7nlQcTrvayY0KhOoi6f7YgUJ1YEER3/UwbWKzrXUR
+bXOi3C+UOwCtBBkxwhOKtiWlz76QUyO9BSaJGLyz+yzEYfxhSc5DS3YAG+URk9Z
fBPkdZRsQy2UZBbNAWhlVpj5tmNw86ECjV6E6cuPq8K0Ui7Fp6QJRO9FQsRtt0Gc
Rn3V1PPiHMKvtZQn0Ba+Pa5Aq8Ix+PyuCiM3IrbvVKq1AjIxZDqAcWItSTBXQOM+
3Z3dNALosYgPZ7m97aN+w0wzb6SPXaQ2ZT1sF+nhS0BsiXY5Iv4qXIGOQwhoHsjw
hdnqDLP4in3JRtO81bhnPQZRqLABFgzqM0EmvY7Nku2CbSVunu2yXlzt/yWEkBuJ
z79mqsjYe3dSHw0/c0MN86dGUy4lNSuu0P+dTrID6zHd9Mutl0yPUVKvdMMnneqD
ZDczdM6cRcTHCu1t6IqaWQvpuLqSWvjfegGp/IKydyA+Xi9pO72TPbCjVVWP48Dr
q5Dc6Cly1u/fMZTnqs/21XDRbhc4E8sySQLulAxfOWxkFkWZ6M9ARZgKJi+kvJKT
x6HGoykQ4UfOehhjaX8v8yJyytRYV7hpbcnWsFWtDnOKs/pzi7cuFHu1ahpXzaey
IwQzgmz+0F09902m0L3JF30SPXkjMIVC7Sqer2NEKGE6BQlHHIzwzNvRHwnBW0lV
Wo3940K2hilriF+XLbaiWA2qlqi62vs91oky4U0wgB8Hbq0ycZkc4kKrMwh1iM3E
PrFmNf3E7RfZ0Qu6UHdBI0RKCjA//4iU1XuuU3pRhGHAQMNe6awe1R+4q62517GV
vJ61qg+Mn6Ofn57YfX6G0l126W1qldXnKHOwpWB+4akeM0x/WeyAUVtugQ1nFEAc
rWbXFK7zO6DaCOL25ggn4OgQ1X/NpDw9dKupz0U+Qb9eteNqop5qta4U21x7O3RX
iahXuOzY17HKvcskRv35zxRawDK59xOR41gTU8HVoRNG6WbSrpY4fL8YNHfrCmFS
Vvls2y3/tJm3NX3wDckvGrHjxHHfxkoRaEr6Zv7p8OJV5yNPpH93W7iMkDid91YE
NwFAdbMp+R1+xBrMwEagaCEOVxr2ofo3foySOhdVryHo7gM7JjNsgOeUfNXGsSJC
7Sez1EdGXqMP67feVSdz8QdE9dg8NwXjMKAwy/3rkQT91S+PoRk/d80o4xCVaS0d
h8S7sEdwqovwWlP4ymQFz040JtQQDGjznYOmjp/U/rRUaupQ/JxqsqCf7jaXXC8p
fmHPJXLBvFzw11bRa172+JK6fV+tpG8vMmGMwNueQFjOmNHQ/QJrB5RxQ6Z0P0i4
Qurq1e/6n7x7mFQR18OxSdV9dokC1a3vTGqPwp7APdUjiPtYrUlPPx8DNfX5/Y8n
rPNITde1WtGBwQJSh+xhP7ve3pMML74DgbEyJQte/qFsbPhWtpwQX3tEqQFuQmv0
ExvWhsFg8iaXCpCOYg+rwQr/5DtYMrMnQ+MHP7Y1bs33i2BCgz2ywFSfCqWtOgaf
rg05oUteoiTb+iqxB17ZE0eMejSkj/hKaOQjMRYYslZE7XAUKByEOylo/ZnHARbi
WmZFkCDHTeeHCOOTkjlwVR9Z06OU2ek24qHElf+C7F8rcUvLaPKABAUfslmaZCXO
qtDdm4fr21tOOL89iFCjiEvUjJez2G/JMIUzNAadb1NnltQ2BMNP9ZTuQmjcVxiM
YY5tJABnDRSFliejwQlF0Izs4Lv275oUI+a+RNuiA+xKcwZ8IMFOPweclxvx23dy
LmOeU8FtRIyiiCEETmzn9b31/LNWr9zy/dz5WhN3E88L1dCiKfHUF5uh+qHL8+01
p31Mdyq+KalFcKfqU4/dPGhET2u9IhnuNSAUDDz0Kg1vTAQtX9vd0tv2zvhPfxBN
SgspdfX8G7gixh0bexjT3BiRXdrid/DSobTcaZzo64icFkUxb7LY+r5ijKbjJ6vI
22KFAfnUZhW4WIpZHfJTZXfYtsHNumjNTx0tSNgY+EmmxRA+tj8+548fcNtbB/vZ
3vVVIsjcfkd89sZpg7hdsxIzn3zI9mxUsuSC7TT0k2Vpk76wyPOs+Og4u8fgDo2U
1DisdUmNGtpBmwFWDx1Er4lVEubiegT/4+J14KjyFs7aNhiqZt/+0exhw6caHrFG
EA/76xNHDA+kXzl0oXIiZOTu6YfAjoCkq6C+iWjK7T/beE1rMzdO62dWip+oeO4q
jYlhrCkTJ8A29WcH8B7BXt5rr4jFbCUO2Zju8yw+VZ3cUbkGa9RRJNVpbUz/wxYN
phyVNKL6sVFAKn9UJyj9kP+oNK7ss6z7Gg+KTveqlyGOYYqmYLgmjd2Cs4a91hdJ
C6dP9SQpnnTNSec9DdAvtTgzhti3cVnGiOMUs4kaX1Rh7N1TESB709rk5mL6M+p6
wSbiT3XUN1hkCRYAE/5uNVTfu3v1yWf7BoiR3nt5TxByqzyvbnOOBFA8RpSOSET4
FhcBM8qiEVxBMbwkAJ7MNWSk8wxFi5dI4E141SzTlJD8iMwJ8GP3MXR49Cq9slaU
CcRpc2qdbN+4PysW2Cwm+uDPoFqo3kuNy6mESJ424BUTw9o9o31/AWV6JuMA6s7k
625u4zV2Nu8+P9U9JGximuimHsu94n8Q7F9GX3MWxU2HWbn+MnR7F0RfmdX7Y8qM
Kuwszf9ZwM1LAsAv3mlR0J1lmWKH/D9VQmHBUYYD9rh5LLkYVlI/iSvCl/QNpc6m
JL2tBacACPZ5MgVM2Xwyl7BsxQR4/wD1Tt9j6/R4RLqhS++Dv4OZf+pESVUreeeO
Lkp3kaDjYkL+5MNFze/uWVrm8wEeX63RYPtFpEQIZCYeXQLpLNVZjj3UhX3gTRgG
MeiBGpcgXDGacLdn7N1/v8en8phfiwbXPpPw01XffyaglKzvDYEp9Y0CoZwKO6G+
+4Z1M/sVMqH70p647KfcOjI6p7VHc/prVJnye+iNr0BvwzKKFvxWlrz3MRGp6tLf
76TNDsvBdVGsJgeWJOa0XVztQ18zE8oyznovJa36bmUllqK8jVjSJl0G0VzP7+4l
0fjPDEHSFkTi03fepH6otv0tEbVzi1EeDBVgWkUKFV540X66Z40akrwI5DPo0hvo
pbjgUa0n3IpAps4TQtKP0raUfAMs14rO9DZsqqP/hzn1pqiOH93YDJYHUir5VFln
rXLzJpMP2ickKkaWCLvBb+sWXymtmgpAWoQmaTnxJ8Z4AF/ODvxvBC4YAE8PpChY
8GvqxGFPFqGyJY206bxC/bdync1vVX/rUITfzxH3sJllHbGxZZvFyvo3ri3TpKhL
UiVV5ohW6JeGaJKMyZjDoq9NkOBJmg3/NAX9d8xx5SC4cd+7avoGvzx38pJ4xNhF
DFEMMLBomB7fcx4Wdc581BgcuRz5ZkyOGmjh+4VJROUCvgg74Al6/NJALDcLBfr0
aTbBptrUHUafCSmCmT70iQdKR5K5qYXGJs928eeUxdSRwynxIoKjksDziO+w94l3
VpEdN/HgntDDdp3Ps6BJaeqeDZYBrjku+rc5f6ccGLYbQ5rQzVRd5qnDkN5ciMim
2jWN4OH9a98itZssdvtdFGwd7T0dgxyJ5oufVnxVLCWcz0bKGC6dParnutM2fC2D
LxruPiss0KOMeBb7PhxWaTY2DzV4A+S6J4iH6WqoOdIIVf3R9sqXN4H90SX3d6ad
AOUO8QPcB9IeOreurmkPOIYgiBXWWZojvBz6HnriuN/mDnm36BTjUh48wUMV1am6
ekj+SvtHqSxuMEgWnPY5nCChz5UkRCGRWOeV4Cp7jmPx+7kTCr7VsKjWNg5NrAxo
YFm/gkRxypVtuPzt5Dzy3mFpYhbt56n85ri7WIPKZLKGyrNKD9RpsRGH5acbfXSX
oV+oRBX9ok4PF9J96MAZ5WyYCk/MmHNdRIbbs9ZSz02L5h9bzOztbEu/1j5eIHNq
V9dEFLiqe16EAJkUQG/czKC99e/tp75mtvwvD2I7MQ3NVyzb+BiqhoaFJYOT4TZS
02gTIM8Z2qtOfUhIfzqocY8zXW8+H9PbEx8u51cx+cKNfuxx50dF1DPINdqy+zi9
afCt2G62Rh9vdHtjC7u9r9n+mMT3Q2wrVaMZNqEqTI63O2baY70Mf2V5hEJ9TXp6
X7RKWbMCbI/l0eP+U4d1zcSBWi+tGpBYhcbwILtoH1p9ugOzYtsVXoLZUaPT2WC5
Jg87ykCvwIF3/bydsGvV1qIXJLhnVbqHDbsQh/Taqf6D5fJV85p2vX+j7Gn+YgF7
ReNa7G8KycW6YTm1ivOiIQ/UsZZN+8TZdQbeH693DUjxvo4qU3PEbI+9Y92SWkOv
9MgR10yUbCNfNpeLF9I74X/L+2QN/EOFEyEvnkIlhGuJaSJeBweCHBvg3LXm6oPO
ILOqc38lS8CPrzmg2vKRk34d5t33atkxCCPUQBWz6+CKLnSwuU7nK1cPkecHmAyE
kbhW9F/hjub0VHxZMD3Kfpdr3ztrLtvXgrS8Tofme6jLDdFTDxc0r3bB3pxjEFYq
oMYxitzTGdg18oJ/gnJcWIu8+cEoA0gj6yxatL0yrOTCfrPdnFdugIXf4Rqh8VWV
5J5VcdRTYOrr8IEFe5nXmtOAVQuTtFjkmAJr9YsBB7RHNjLK05o+YyC0PlcxpAcf
nIoFTn+fwlExsJuGBX8aISRa0dx+mYBOXAA5tYdhx8SsySs9D5r0i1rsrYHCJgPs
3Z5mkQn93SwjYfJFoC/LP4DxIKafQxqrHeNXBFwHlctHJNwcTKipyyuL2yafw9+Q
uBVB/nlZdjbKBCjUCt4B75OTt5m+FSukVweOGihqk0fBB3tj/aN4vGXDmT8XNBr1
QKcSj9+HiKHF3KEvdCiTUaZun4TbFoWE2WB9iGboBNjJ0ECtExb3OAHsv5CVdK6o
Fku1lXU7vgVfN8bKCEpwocIIy5owjw8RxmzGSnf9mljSPSFzGc6ei+oX7jQB+Yop
Xm6Q12o8gdSTGPL+3dSthleUX+5Ll5CNZ9VlZhD8kmzOqocYeKhO5FKjZUAKczOU
jHJiWuHttNwyqK0wfZaqBxeHVGhaZ+c4PLxx3Wb6GZzZ0PDm9mGfvj9iXeWasZXi
6uRrq6ZCr5qR445zmTQbuyFE+E0CPvVRjWwTU2q8sR0+kL2AJ0hnZ5r4i8pT5RP7
Qcn+PuwIGnONHDCTZK/A8IOld1+1O1Pcq5w+f+mvAtXqp+dMo5+tX9p6Lg68chV2
NkHVB9d4WL1nXMvPV9EhP7Xe2XPqcyEr7kwu2wUvbdfE0WvhyETNV5fl5p64/AR3
1pDfq6Guul63YFVCHOGtH4RvYy2p7SHKB4adinK00VcvIvC5WDD+ENA3g4rmKfJY
tKjYFpxjcw3jrikMWwZ/VP3su7+EStmkf9nbaSUpYKRkncTHQJOQglPB0Fgbo8uO
uYMHfqt437+7Urfvjgeml1Jh5jzSMqhHcDnEKDkDlULoxMAoRUYoqynRh1LdGCxU
qjwfhfOq0dtZi78twvzeaOd5All0C9FzOlp5x3y8G5eY3PGx5uVHI6B5OuS3J2ms
isRayvoNomFjxa6xqGglFZXy+6kCJjoXieyYg9EMryhmZihbMUzXHc5FqtyF2NmY
cjYy+IHKK5SfxhmNfjd/TK8jUikQ9tLrDFu8TBp5/xeQBImG73xaJrFFZf6lBTqf
vIXVKktQgMLgqOWeedjWEPhF3rAzBiE5lusQ54aB44ZYxVS/zTtjjY76p0c9+6Gp
34BMvXD/7sUm1yQiZa/M9x8PkH+AzUf+Rg55FNSL0y8OIRL+AoVSvWHE1zMceEZ5
2v+zsEMh8PI2dZd9XAw4GFgrsikIEDFhIbE+3hp/8l+7yNRs596wkQw+x+/0n/qp
perv/upgoKK+QoTEino1tQ6OGKcAz4rEt1b7GPUTOzof196hhdk40EJtiZQRhXKR
pxWmhU3wOfIk7gwpHDv0FkjZEWbrwlRxzOcUMEiZV2SUSaMmRzwI3Mop0j5wEV85
8EPL3TZfqFcbuOoaJizBwRR/KOCWQdEgqMR9j80EisI6HyK+EP4RkZk+0IT0hTgo
5UCTc2ay/sZlO8wGjmOR590tU4A6Dvo9+HI4ywOFv4SQZzW8xOV1hIWckUrK5GIq
kLfWFzdgtVBT3ZfpSXFqac8ew1JcH0bnq5ocrIWd5GEf5mAg2+hPuOVzO+cy/5p0
awdo22vUIubsOe8a7bOAbwqCiWzinNo9m+L9Mdgvl2Wc2I0Rez4nNrqPS/m2MfRf
wnJgoceDBxEXJbKBOo7pove3mPdVojYJ7WFZRv5x64gNKQjcbIrft6S5u1zsCJ2v
wCFoj/1ZhUht1JM5kAqMuSGtO6wGs2bWAkpeqFN2n+6MwGbh1CnhnrqoX+a62gLL
W/COdSu9/6/7q/VY2NFnNl0rgSM9gkV3FKauQpPeTmOkIikJlOXkIEEYfPS3SGKU
glRbSdvN/S21P3Vcgd+6Tuxx7G0/ybaqS7u3nHQMeZP/OpU7ZJ3o7IU5xgLU2/6T
3DLEiV1jIATLTloQTqAjN1Dmg2/EYC43FaXrtZEg0IcRjytAP8hNLG4d4NhStvVl
4LbLjEVjUj6KZOw8GrXKod5NAT0Ojojj6G4gSQM9cAWzZjumcmuDnpG1v5SA1FmW
/LMXjt9/o1pPPKrPzR/CmuB9/07hiviRfo/3BjFqi7bLSy4LJ8lUEcp6clMCfRvO
jYjJsLaAV5jvugO+qbyeRX+Mwg6cItcNMAReqiNRCW0phlydF6Hs9eM02P5FAVN5
oIUOnwomrm/u1dlY0V4J9m3J1aQzVgr8e9pLJxCtPuve0TVJZJfKb8VlUVI5gyNm
7jdRnJH0anqJaL5UuacN+LAPX8EyeAjkQhgpdSAE7+u5mcvHOP8F9nSgG3VV7q6U
0YrNL+c0TYLVm+X8pBrbWZUKsy31uJw+ckdfmocKZ7r6Mivr4IPgTM7EG/xiNXDJ
MxyYFzXWgTVn5ug9++v1ReXTqxGRz9iD01fDL0spbv7Uxh77fT3a8Pg6xxRei1f+
icxjnPr11V7gk4uhh5f6hPlD8Qlkj1LwrwGTqzXyFr/s9nud+FY7YPZt33TLvr2b
T8cJzK37U1XxKFQdCDvEoYD9YW65EptvNsrrdz6TGY9KEXMoMyScH680PS7KViDL
Nb2e6GpXyh5xawys0tqrk/BL4mBvQZVqFxY/x2dbxBSZoYsTni7QUY08h9/xPy06
tnhfkc1lv8etFpdLINDXQQ450NKWFFqlVbQTUQIvo4Q37NxF2XNlJQUIATqnvIND
ef94GxDVMb4caSvcecf4VGDW1S+Rfj+GW1i0tdOGZ1wm11iMzEcK0pVT1EGD2q31
weRp9uTynyHcK0Gv+6aUKTrRDDUx4K/+Xz8w3Bu734V3VTNcrAy20UCMrdlV4KPB
mgC5+Qg1HsaDhgJtxsNzDIMwLGzHE01cCd1Au8dHLxGEmigi/PX291Uv/Tppr1sO
gU1tOZ2uiOeDE7z2PThYXivn9JL5N0xX38vQxBxdAd2C3Q9bkOFVmzc4VVbSWzQq
kTqHjizjF8f4A0D3EJHVT+v3F1zt1ik2xJP0ulaz4vl+3Dcz70GPE2HhyoLT33Ii
913GWvRYgy6A48pDIeK9PMUxK3GVSkG1XVr9ty0KkfAXACGav/8IWPVLmJxXdPNi
C3TQShhrk4IUi5Hb3a9YHa1vT0CTjR5ohs/AWRtuv+qpL8q5GoIPOtzFKKAM3RQE
THpcyJ80T3tASr+8wkz6yOmdIM1eGVoBwDI60TwwOLJWPJDVutXkZ94g9xTLzjAN
5Bp/WSADvALKX8b0E5IPEgXGKuJecEE9OLQffKm2E6Wy0rHyU7wF6x9w5oGm7rK2
GeDL7YV9H/xSITNBDBxTHq7xJDdUcUptTAmHOO0uzvtIHr2Hs6R3ekhRuSW87fx8
QzYCVXnJbXvQrwCbwlOyxo6TQrukABayq/0WwI6Hk4cJKdMIy93j46mH2Xi2v6+e
hFAVZbmd4qcxprn3Me0R0wf2grqmrCPRskbMRxHMebWh6eVppxBtSYOnGHnqKHoT
MXRpoPIqhzZppxxz8OrlOmzqjN9iklJGf0wYOmGmih3frUst95aFh1upRlJmJD5r
ym/7el/X2VgcLSL0r2TTPQr0+J5k56MW+lRrCojruJuWqG9j0tfvxLslRcZ14xx1
D0gwZETw7e3rk+T6xPDSSIYUK/UiCMJ+vbRE+BvJ75fyCsb06CNsb1uJaFOnhHom
hi2sUwKck5SO0Xuj66hp8G1aCP+h7eGBs41KKrGiJg6xfQbva7iu5G0068pvB0WH
zN/GANrqOdtvWb3Qssgvj/oFNtk+a4ymALMDjCL+syunqkOs5gwbUBfNaESBLzZ5
+E/KPFtmBFKJ4PnuYAoW4xY471fMOgixAw1OWAtj7P2nQ5UebL6UCXeesh3f7Eqi
4usXAnW9Uhhn6yn4NYyk0d6Fax6TS1pEIGaUUFGe1Ql3cq7s88YViMa4pIO3nUuT
8dI3jEfSVDu+D2L14NrzP4hSIDKYTzeg38lzm1zcff0pmerkoEot4yNgjCMZb5av
IQcoHBMRudThRbs9uWmi3HnwlbpfTF/dfwhfa9QJbrrikw4kwlfrcM1JvRIYoO3+
p86FQ74SJd/aVJgYvYApGsLRBqwevTFAbnmpbjHuIE2H3Uv9FxlZjrF6vf19yZHg
irmq1s7Qq/ZvezngkOLKyJZ8UizIWCfarzWUFlXC2EOJ6cCI+WeMy96+80Fdd9u3
7XdAZORCC6bjqQuQpZEH8Suf6DS/VpA5VNIgm25mesiON0JNhUnI/bbe+365uCKP
WLW0WfFGoeiDFcRhAIQXACcr07hb6KABMrDQodsajNA/XXmPsn05NIRULOpKMnQH
QtBGl+06o+udE1xD3GY69B44p3anqIUB0z9yByqwqTksRAqTlhCdCGkjH+ks7EDA
l+csgmx9l5urf/Vt5I0fWEmtyQKUilal+EjQx36BqEHYTwOovH4NV8b76PKkbj3X
7VoAprbh0Cw5iZniLhwsZuJiOrOpua3cqMgoWIJUFtaOxCOy6GovqItPyyOwCxiH
Zuxd4bryU4sr/dwWMP9DiQ6o1dwiDD6eclD3V+IhK5wK3GL0d7IaSVibNHQJAfQM
NFSDMGpuo3gY5AKkyeIvJnkCjPImo5HxQawVagU8JPqpi23gv3LQRK1o1q/O24ay
L68U4sYgfhUxoH7vd6fU6wcc5iylXJdePJ6W/mc9pWbmnG4hYdjftQ9FOjI5+BEJ
1erEDPBakZn/pudEWBlpxMSuRlBFrEPHYMk2ayXxpfvRZoku0IdxeMrzFy2PxXOv
CzCbsG40Z1O3jvUiFN0lt0VSlXy2GRw/hzjO0Q1gkV5MTJirpzLUKw2CTVkoff0s
zUpPFBHETSyfTx8f8TYMMYWPUlSnfebsAFneyV8tb0uO3ExxwRynfUMZYCQHDKzC
m2tf0HayNi9BHXzEDOzKkrmqmQNDOyhcweWaeOdIE4+iJAByqCoByA7YaBet/UF2
1OX6ICxpsyNEL/v6dDBKGQONQzphq/sUN8SkpPknmmoOM6ojaJAkgINvWJbS9/ve
WMCxTgnTIBVql7MMhj7FR8ev1CKplnx21smNHnQZMsIWCYmwDqu5Nb9zMLxy85FK
qGjUt92u/lXeGej3AB4IoCeUTsPTfTEfGZ4yEdS6FPC2qPzE1g9KLOUZ2JRukyOZ
BE7UZv34Yh2chefNoFC032kWOyzNuTDAYKb31Tb6mHLCEQR5G42zC5OaxbqnR4tM
NHfs6RHVvaRyUJG5ROlQJRSDzyNSJ7HLg0nCdNFK6RZT8cdopamL6XzJrgEpsBA7
drkz3HP4nckJK5B4f1djVldeF4ZY717LQCp/qIzSFi69fw50LpfItiZBRajfzRXg
gwpfvwbPTrBqSMgkPYig+oMafjeIuf6dW4WeWZekvbQGoytYHk3BjsHDyH5vdxTg
QZNjXO91lN9fvfYHRbNHS2aFGWOoPockq9IYcHU3mDAbs6pK8AeSUz8Qu+NyLE2j
vs5+QLs0u/z4kOmwJL9A389pSWxMpjhB0pSChsnjyYQH81slvWutr2Xu+0zt5t8w
8KoDAiVxvgqqS32QmUEntwXja771tTZyaGYI1XXbIKCjFZVBKn+aU1S0ZMHBR/Vt
fDlf9Haoc6I31i7PYk9NoXxGb8Clf5oaeA0qaZB7bllqCWSN+UnAzFaGl+sdTA89
U8XHRWm38B7Gf69pLQx5ms9V9fyPPD2gimZnSwda9mrn0eNjTI7uR52OhS3i3ISE
4invlFu546PrES1ywJ+Qas2iGqmCl6KsaXwqMjQO0ceSLfz05llXWHa/EGkt/Uh5
nbmegrr9R2OPWO3n8EW6kbE5TQJWhKK+5M4AVlhUSkq02xZC48iBUmKUnZBQBbdp
UY8QuWgVz4HG2ArfsADhS422j2ig6IV0T3Qf56tFQLTI59LwZHIKxiXgEqbazUrs
hHdWVvdGczqOVHDEmKc2+BrZTyFYl5z7Rbkc+IP912fbMKHHMOXDKAIWFQ/x5XIV
eABzyzhVsfHz88ukHVIRGxYEFmxZRlunh6gUKEzq7twH5cZyCZNDw3xWOsXftkj4
UyPtWBRiv9tZvdVwckh66/pG+IJNJ6UQGa6Yo4JAPLpP9YFlCKHfyHnxKUVUt7Ug
98AsHI3uWYamycwJjcywIoaSZBgqhCBXpBpkgAvoihsQv+YatRjZ1DgXh64xbm3h
5cq3rSwebUKeAa1r4sNdft1t86w2ubh7ws+/rYk+LyjSMqiRBLLgYmJBeYdWqOXK
D0V/9CDlKWQaiQz4u0ogPW0Fo161Xcgf3LMt8wlcPIs946+1S4DS7HRakjCGUjS+
D/WKGrDw39w9kdOkLU5CpdviOeF96Ub6ec7F+Ni36yRYsOSM1NRkMGWCVE6nfzv8
kdVYxjee8ZZDECfstiOK2iDZ34KSiyqwyvKYNJoIBg827iNu8iezENEKescg5YNH
1a3XaQeNevvxSdmnA0qLrKXM6pQZhjbmE8lImmP6YFc3AiCUReFBr8FtXPC7I/RR
wBDp/YjkVfZgS6yvi+6SrpzFNFBN571r0tqjxLhJGf9NdfzX3lRfzPYkZQx7GxNU
5VNXvklHBaxXqukXfdjrAcQxy4HB2gYAYYsWtqo3Ev9K5cgMed8OSJbkjyHxdL8M
JwaWZ5xcY/fsGPmvYAJKwNf1apON+y+O3OEPCCQpgn+li2LcrHawsBFyNmfCqbbI
ZMxF/S/XFbzfq73N3dT6nK+ctN7IPj5TyMyQnVGTPzc+sZ/5KPczkLXPbjC+oBnm
nT/vumPuskKt3jB5cXR3tytjaENQfHdUT4FMNnX9FyDzU6ZrIt6nLLVj6sPtNF9N
jEvDAn962WSuicgT95wGrWBQ2qxh0qHvozrB0Q8GHQHGKRYsOWAAVyPGQDvqCRG4
J4cfLyr9Gj4PrPweJDrBAlArj4gd6coN28ODos1Fr0aUmK4iM7VCQPoIQ22IuS97
CT9DOCazcYTuHDVyilunYpepb7BcPxlBMwU3hGU3SUxtiPe5pyuZv6yJ//rP0kjf
C0ft5eUSFlG5+u0aSj0AHKEr7z/pxvla/RZybaxKGO4s4K9GyisPd/arjfYqvrFJ
bK81hN7X2hGcu4M52zYwMhT3tRwg5w9ec0xlMBSzPghf61C0EPg19zUTbzRA0Bvv
Xyx1ZcDobwirSfHY0BzebljQSWyTvkObSuWeEivrbkv/Z2fd/KBqr8plgG5NKerD
hRkq0CnJz73b+nNT5eiOverHnR3MpiLB9+9o9qeyTO7ZC50XLUpICgrYnzC2SGhD
E9ou3fnt2lbE42Cubqj+no5inhgmB+YOoJUbqcQKbx3aCSYicx8uR9TfMlNNf5Lj
MZtfz+zaUhLAjQDo1v+34InpUETdHWYjAEJoN330bsDkNraKoAvXxaUtlWgxvfk9
kjP6edjEuJyAOF4ZVQJfNyoPEpElzREz4Tu3G7ffAbVSc01glbZahDgIKu2QoIL0
zRECafyjXfNmp3kHsVJk8q9Fie6p2NeMDNCg2KpM2GMN12rVyj8vNx52AfMstZ0a
N3OWvLVK7cO95sK/6SDSiydydsFCuPX8XFb43zxQw5TzoBmYvwRDt3+sOpH3W3V8
elkXreu0sk0x4ynd5eEIFIYRRUCz3IVjPgDwqvyRjsh4FUR3qggesNbEEBKqmNNq
ecllm32fYLXYI6autZOnCktOtuCZsp9PBx82+JTlFLW8RgUz+AOdDFFSOyUCkmpa
r/SBgLqLiJYDuOKsgrhWDolB4xVUJtYGVd0m8ptLXExI8bqfRsUZqaNXhbCjlRg9
pDUqKSb/+bqqZ1/IumwVUyW8aDOOSJ7lSG05j4uVvoHBEmlBvaJC8SMwZBVa4Zb0
HrXV8KXSF4DVkT1GLzb8Hsg2fhw8BMavMhevtHyD6Wyi2056WIUEKxyTXadUn2V7
yFSRJoT+mvO7TbLeMWg1YddkEb8YkCewsiBfh8icVQGz6eKDXMu/eUrV6yQGj7W9
GOPkwa1A8TIvqR0+yNg6rp+W5rcuzHkdzGOnln5Tf7VpG+YOExn2CwUJVf4blFmt
bkRQUjUYzLFxrNK6qKrDH0FJI7cN2sEuIjUd74vpEL6ZmM9h/KbdJ5LX6QXc6Am+
zhBQbpWbqF/lAblu8ixWp3AlfWfThNOHsNuXoV3Fu0y9waHo6gNeJbJGTEHUqEY0
mtHb0p7kSu+VhG1mzZqLUqa54zym932N3NCqPNhc3H+byW8F0xi2Ex0X8Trjvk0u
nWhacIA07lWAXIlan97TKAt5rz28rAjrj/tUzgZG77vg6X2AtQf1hXwjCJx40zBp
o6jMk/FhD/X/ncLQxvQysSjw/ECAp7ezQqccnwQea0FsI4cFLs1ol93xz3K3nknX
lHy6Z9WnTheKh73Z/dmfkXx/z++yx3IFpTzJpt4H6nTjqP9p9xHY6J2UpKnsehIn
Xs7gC/Y8Z5t4724tsejdFiZ2MpY7rDxb/eJC/dfaT3SgLfXN29jQyppeuYhB2ERf
zM2bptV5fudkHk8HCXsNkg1Z5HMNNm6vtPl5JUzJaGFH6PR+Szoo1owpA+1Z+RQP
FOflE0Cxx7/dYj3l9od0RHRAuNCSqOtZEURX10qtmky6ROz6ZBw4yWOzLBSShiCZ
YZk2kYPdUUm3g9WC+XNBDyuPFI79RA4mF+JuFqEQQXHbZr2k4XP8bg918VzLJqPN
4kG7G7kbPwkXD2xgb80AQk+YbjH05IGaNZLcZ2s6/2SvcL1rFaTrkXDWh6ilO6LG
y3xHhIeF2oGkCH+h3AnNxFUB9YwvfRI46pYURX2rdzmGboQoUn7Wfhth5VbRHITM
cUGEmbBuT3x3t769unYM8rc0fwEHB3V8GhTWFgA+tPfLLN1MkXji6rlTJmt2IemP
e6R3/zyGl00s3lVjWrXA5YpB4xF479lNKKIfuEwaODpv2KXKWlZ+1daOqOTKwosN
r+YDGvYLxaz8YwaAqcVF6kqZ2HHXyxzfG1bWvGJiBa9O0naDFRYHijwrZqkDFKdB
ikNOuQdn0bzHWyUhVZwn3YHJNgxEpWjgtm/QWozmsCdNbVdCyUK6Ho5rvdJG9kpu
stkVpcDYbiML7cjjnrlfrtjO3vBIp8iAGTL8kdcG/3XJtB0Cz+afC4JY0QUoM1Di
221gGxnqpjM4L/T7ZnJib6AEP/6oGPpXH23jM+rHm4c5ATKLEVKaQfW/mi9EoYyv
/pUPl+biVYv+K9N7DUnVaujztkpYo86lFwCFwZL9Cr9IMFlqJJ79V2rBNn6i0PlP
RX0Ytf4/wY/yKbSfMM/hUfEX2mKtfyUOn03WB1Xdt6jQs324JGRyQ5sr86AiKvdc
s1QzWxYu9l1GEY292kWRL8on24TRB0kvQrVyJ+ofAdYZLDUwkdBCbu3fNq3+CKX9
78fBVDHGUyBdPxt5gpq4ouV3JV+qROA+VNfsA1MEjohUBCpSXPVeQkCoW8CGux9d
oO77yqoXoMRHHzUzCyjviZW2O1ISgdMJeI2gFpjB/ixAtLZTzVus65qZe1f0iRJA
D8LieLYMmf4hNeHx6aAFdUv81V7xoRBA98hMT88+B2CyCfXBsinH3bDBCsy9ExOT
MIo2BLkXaH2uFkv5Re4TqSOv7SarZe01ZAp+9fxjjeV7RilUNW5zPTiMG+3ifIWH
Ihd3odRNLeTXEiNLEJeI8jGr/AJT6TbiCTRVJO4jg9SqGCPzoSu196WM2ev3KN0j
//rNSN+FzVktSPM7G3GSpdqudNm1jXqoFW5bqvTTiDFkRCtOlOdLx3QtX5jdQO7E
BPi3Y5Pi8HKiwTRxMHBHTquWUfyRkQ0uXLwkNFZ4J50wKw2LaQaLiiYQYAtovZdI
8FtqDO+VELX6iDw6rvwfZMJRwyDPE51+GfP9T3SOgGpC9q/xpazYFvjlTqkPJY97
PH5yVojmYwOKRkcm59LmUxMr9ENjoTfX5c1FvOL0te8QtYdY3HTeKADvTlwi0KrL
FDPg9yVK1/t68nz6T/FI4oBmMSTNUTJ9dtM1IXnTDP9SBkHiJEIs10VYrj7Ael3/
PYa8ylH6mJg8YOb+Ll9JWHnL0JZzztBA5Onrc9UQMdFX+gFiOdw8lEVshPoYyrIz
lT4GGy5C7RLqOMmdgV5BMYSjyOtI6+8SiLBAASwoJcdBaihlQQnKWsc2CUQzdgvQ
zK81KpTgc1Z/Cr8PVsNGG+7VYU9tLA2QFkFViN13Wgc8D+6mQqxNTWRyPukgJE4y
JIHbV2MzGgc93RhzP6Qsvh3IzpgqlUc6Gomv2R3+npbPA8xuDfyV+zCHAYtGt5k9
pbdfuR2I1UKzBLO9ebJr47A5O1LAMQ5jHtIh0SDG58ycE+LYccE/6IpgMIIi+9DQ
hmPcdflKmXJaM7AuEGU3H8Zi//OZ/twATxDt5V+VlqLS+FBpT+PPz2FBNKhk/cdz
Q/SDqEtw2MFl3BPzT4YCr2KTsAY8fidjzIMQCeYsc514o1Uxv5I7HDdSbuI4g43K
v9wtf1VEQkWEOGqe2YPLUTqsNE9euwUkyPtO2xlZUMOO4x/B/3qXfnq2rMxivhur
pxxT1f/qOaRXGhhIAy7u1ritJeglJIfjq1yIqQ8aImnvBQzop7jxM6vViq2v6T+n
Cj4KpTmM3fJMp18/bPd/wSo6WmJKwG83st58cHVKUM6XTQt7VNGDNs1B2RmGb3bV
r0nci0CKzeMBdxEHKNs6EzGN+ImWdzF1ekhTLoFyaV1Cnt8AV06Mf66noMODisDy
UiSBK4o2XDbQZfmHFBBw9VlTIBkQ65D7jXfrCbWpn8eBNNy0Jfl9NbfFJFoXY7XC
o41Pi5b8P5KL62qzQlMjTg1rpy1JPLKcrDWe7GaPve+Wls6xK+yBBqRLADbFUfpn
cpu3Quyni5SSmw984en1Lcc9eCqrEzgJME6DOSigAdSDEY7DsjOA7uKZSrGAlSbh
fiW8ItWEgoBALsftHR2UHmyE7qwckmVnNIljzfAWN9eRYP9fN+xS5beZM8I2FkLM
v2pJmkKiTBFQHIV7woHnsu4nPPCq5E7wKvYxQb2UYEJx+l+XsuU9LwoCKJGlRmJ4
oEra2/9LKGqvsEG8kdwbWrngzc48e6hBqQjNASFg7fuuF/4uWXFrZERT/H9vGZB9
scrQ7wsxtmdKxdCgbH2/CSGHKxzL13pcmc8pWtKVSYhj+iDewPI4TiWrg5K1zmbO
gbHT69KhOKOVX7j6ilc3YKVs4rwpNPMHzR9gpQiKUQuOsqEskVzdOGe9KBbgHAbU
J3l2+x7O8VWAYbF5rp6J5AvbOYYnKf8GsQwnOVqSRCrfX+rg7gEBqARjtxqBzbby
aCYc/vEowmY6CBfZy302RLdahdkeCzOsO/WRsu1yiWw7DPRekkvDc0NHjXGeNQ7M
Mu37dLm89P8TUGQGoEVeZb3pFx3lWdk5w/F0b8QXDStMt4C8WDvzzGuFFLBc39pr
bsbhiQ0tuTpu0LnMN0nh6tcw0rA/71IXS/eCcW8Bx7qnJOtUzZx32YupYbeudHBx
oKoRh7BBa6apk701jfupuwH81Jewu2CQ0WQ43KKRxkMjsjVRy8+emE3fbUM4El0f
vUb3UTp/i5ZyzjS1fXNiU2FOYlQGLrqIr79HbfAT9+W9vRU+stYW/g43Zs+pQXKk
17Q912nzrShmP7Jw7C95gi5uQTn66bEX08c0kpZCKMUxV8UF9xj/c4mZKWM0k2Bz
uptE0SCGbJjBI7duay2rtSwB1vqqdcY9pkUA0ByaQl76DaTFKYzE2TIoJhivengU
+orPJf7NbHjgcLDYrXS5PF9x7oglLqey6aYcbv9fh7vkbe9gjOFT8KY5TG75Arje
CIc0LCDxMf9AJ+ZQ6M9HCOnXv3zh9jfyDKfvDWgNpQhL+UtCulnP31r471/VX+/H
WsXUjSU2vGIN3+LsjCa+SsTal0V317ldsva7EHj60qYGfAvFnz8z7n2bVk4QflL9
BAYP62tLTSww0JCG0HmC1tw44QConH2YqN2tPv2hPJ3hcyzmWaGX9D8YvvzJHk40
zieVnbbHK7klbdBfT6rM+j4Y0+ijamtEPqRyjapyIPd3N3rGir4F4NyFAHDcxnuB
edYCnW+K+rJJtlCBp88cRQKEVfOKrGBDsQFQ9IzZ1mC37YJj835ie+AvFHje4boP
SnhwiS8SqS+6IK0zwSRJ649xLXl3I2x2mA6FDWE2tsjgnMj6kuVELdDeGZl3RSKD
XjpDhE0V+9Gup1glE1fP4oO7THsh9Th1vfJ/3pSOHBrJmvq4zq65Cut/7zfR+xq+
VRk1yFo12YHVQBpyFjjaelDXSvyiTHiCCVJL/1P2PTUsOSit/kbHdhkdLM8qs78O
jf1ri2lcbzqrNze3kxARiwjP8r2qOtAHJHuluK4P3tpO68aPCC37RTXysa7ZhvkX
1hJmvRANn0S1UiMtSXy5GMY5NBpOpvz/XNDcOHvj/TRfD72vbG8NsF2dk3kW5KEm
hTcolVMyIxv/KQVcJoxtpVsW1ZHKml0L/VlHN0sJfrY6Slm4SwLmmfgAaNgc7Xnr
FO3zOm8T5iarQVKf2xUhUOr+KqxPA9IDhhY92+DT6F4jjeJnhl2js60yorHG6UDv
dOCNlYD5yds+1FJp3Y8ZwETPLFgL8553VsPlLT8AYoESVJooAKHaihi55tp5JIQb
m2YGhnAJ9SU2dUmFmRqPpZ9TH6i8LbY1c1hpsUi+cw2JzYrECnBuPRXTK7FVSELu
73exUN5nV0dIffEXgr+YmQz8pNBQp1NO67RmLL0nJWRTNTqXkdk//QBBY2jNVGNb
bbm+uMEtooVpw6I8qQZQtxOxPvdXXPeoQC7CIRLMDirZPz8f6yP/K/7cBwYi0S4q
xOlbgbBqCBckz51hd4dRxTQk1VGPRdtHV8dOKy1u4meJEJTW/DE8KCoQ5grspjfc
I2qRNQtPGhfa/EeH0sLzYEZw6RVIzTnfS4MQH3Yt0X4o/0wBBMYt/HC93qfi1iz2
TTvmNOFk3QR04D4F8TGmipV2QooAlEnCXJ66EapqEeCN3YUYjEkI0g7Xas53FJ1N
fQl1rNN4lab2jkhw00ccCHpYG9b3wyxtppyc1J/brkaJo6UOzohd4vxhWf098N0/
Uye2dxiUqjC68Hj9N4ypgZILDS7cH4YE6bGeq7Y1mCLAhmjCIOlXrds+yCyOWXu9
2tfK61vrOJtZt+rDho4XJTMi54+P8RuxhL2AMq2pcJBjOxXqdBgUZsKzdULUqpeY
ih+f6cY7BNl7YP6Yd00uVkkCEi3I47EP46QEFYgxoNyTSy4GbJqnWuoK2cyEazL/
hFTIUNS63Z5v623G5qOT6OD+uVOjEWMCME7AKpa5ciwbBW170srvnuNO3YNmg7dC
fECzNtrKReJ6Sul+1gQ37yRqBQLnHlSc4TU0/+GWAgVTBM8EsQHMSAf71O1QgxDO
6ebvon3pqPhb2MS3Z14pkudHqckYQwviUeJ9a/rhKqWgX8XtKgwEkx45nGUPutjM
GtYmFd9ji9s3IxCJQW2ti1tNPmdKWYODEaaW5XKG+0nAvCofXDqpIr1BVcpLKb6E
zXTbLIWdqtCTyFxy2po+vh9pfjXm/oe8qqWl4B/ttYwKezCZfabOKboSYwVwq6ZW
B2sYxbgTwzg4U4yYSONC6dfTbgE6G4wil77/0isz+8tJ+61p033AsJ/wTJc4/VmX
y77DGL3YH1Lcavq1jL77rQViSUKyXN7cMsmoIVawPvdOZFNwvYYWH4Ch9H+IiwQm
GesCdwxx5csPpy5fDE+ty8VPj/rCQRVfJj4XImL7xTh1eeq7zRabefLJLQyqokcQ
mgcbZGAoAUEzpvJfhNZ8VWaWjPcEXR1qp5eolembc0c5At7p7uu3+iAoBzlo+rPX
aE8LrWB1DeE2zVZTePEjgTca1qLHUYrgeHpCDY1mBUZsYjqUZJZph6mQx1et0LHN
VrtMHLCUE/dK8Skr79f5MoqOhrjikTZH5Cqq5v9EZRfq3snh1GPJ4RbOyPamR5Qw
9gI5vowVbz0ekdiwgoUC+DlsA92il5m8VCPLd68AyYcVRAXQx75aUFsybZZ2THRg
DSpnOUWcGgz449F/jxBquHQ9LPYSsik3el+wTkF7AdvgJ7v0h5eK+DPAodQboCnN
aPumE9mQS1Y6MBEAkw4Xpu2ckCd23eZ7j0tPSMRMI1Os9w4WLv/b0bVHViI6c2JN
guyTNCzH0xO0KD4ymasywKS7u37ihwM8BcPD0t7XMeIFQwajkb5mrQdB4reBOGAu
3KI6jWge/5C1LYKyhJIb0yWQtS29xKVkEzKC9B267J5YL3a75TDp1vG4q8gexFPy
95F1iAgrqOIXVIs9slIvlgbIfM2ja/cABhYCfr2Qa/jAbZC/yzfk6zY3nCXu1Bnv
YrVWOie4ZliQZVaLna7Y4fDhm93rDr4/ZxrNbJsNlCcXdn2AqkSko7kzBmLpiJ0A
okZl4JEJZYnL0f+xvJECAJTUkd/3Z8dEchqzl37DpiBEFqKws9W0YLvvtFqMdLsF
efUVyqInjnClZbpLvdGJO5D08h1XI/0fLpx7s+S86KP/XmabP1iSVKPzprO0azwi
dF2UvSsgBcdj81TJ2d/Y9ba/JmL1j+q+4LcbqKzHW77vyX8LwVS+g/17ya0lvc8m
FRrO4XnrXXJFVw3Fr5QFPTHzqKdlJBtFCXzg2kjjXMRDbu4iIsLyaN2NAIKeGZzX
YZ5nnmA06OPnNTZapaIV1UF4dweRz1VH1SAIkXKkRHl1iVVRXqsNbIG6nqOu5QhC
+H7rE47CcfKdCFvLLeDlnqIQzM8CBJwLzvogI1n70vGFlaiNiPFoVQw+n3ie/Hrf
t6eIh7yiSjIj3Ze7AZgGejUa92U4hAkkTMmIJWybZ0a+4q4eAk+IeXz6ZPTkhn+6
h0gwZYrN6sW6ukmJWhkYr3QXjDdxRDyPanomRhrU3owqmWYXLs6mNH6E3FObDNEn
WfX6hebjEX/WaqYzv6G2xxezVTlDHZ5g4lXfX0JSGySYEADkaDvuAcE1vM8S7dQt
aqzmmVXERebF7bgj/iCD7nNH7zcP95DKCv2puPYquAdqvpZX06K1a+l0Q+aKZsAa
nli1jGHN5wzADWPNs/1rJuHYdKSXVhywr8orT5izkGS/h382M0pul4YD9rBUJwdK
5aeeaKg2ubli0PfSPD0TELQLcenXDIfC0RFqK3+5vUHmi2h2XfyJCzTfw8rsUIwq
FyBmccqKixqrgjRwf1FCmQSUG94zkEQR9NkTeUH/oqBcVdnbq08NBLal4MVUCrxr
QSngBx7cXT4Hg9efSdWshIxdmoX9183b6U8xfcSLPabU7VDM9rrGHd91IoAXrRDO
psdCPNnqAnrhdf4n/texUbXwt8veB8pqq4h8HceE3IMqemFxvf3LhFGJEEEg53Je
Z2WaZLnFHvRmgc+kEz3dQN2mRrUDL7DrBGu2oS26u1eTTKk8lbQP0qPErsRwmiVe
5Mvgh7EJJ05L2wSizLooE/wy7X+fHMdwdsCwys29ifhiEybzUrLD4GuIImuEJiuM
Py2rIHKV5LypKyeabGjlxP/LxuBNx2FEM8RP/mUL56qOe1QGhEgkUuS/qixwJF0b
UqHsNuzk1YpMoX0NGkys3PFayzeOFGTbaqGl4+J0DyD3bEJdN8KbN9yipeFVvGhS
dljqv6sSUFteYOTySh+u83mkN3gub42AYMnO7aoMdmJqlphwmR8dEVjrJInBVodC
bnMU13sroKTnV7SHgUaT0oxNWbipTebxvfcBsfWpv3pgEO2V7rmuw7KKKphDt9iI
0/ZWdSKbfkUM7F6iyGDzhOwoTOwQzVZcmsCoidPDkWTW/yNfGNo+eZB9Fzr0bR6w
DHknGkqlZuWJ20i2ihl+TAhAN0UpV/3x0jB5pr9L5Pndy/gZfrYTMpBi44x2LBuC
w1bndNwUcn5QCtlbukKqThGrUezz1soH5TiV7nAp3N2CLLk7g/YgOsRfP3j+cwbM
8DvEm6bG3cRV15VMuvbjDPu/eAZB5oETrHL7V/xITNCHtteEWK/fsH0rCF+hvGID
X+B2IR1khqOzOt1y7evc6xz4d5lRdvVul6RQ7MqlUnumbmUiDEV1lGWbjfF2zlFe
RRzQ9vbTDsbYSY+zE8bf+pk01ZwLxnPmUbPqa9SZ1xUrumtFUL5J/VNoqYu4nA71
jsBFYJ7RdJ7Crlte8O63Lo1R7IkEeqRg/SuYshEREfZHC20mRvzC4fQiWn5E5ti2
fTCSmh9lLQpm/ywOJiWEL5Wq1BJEMgkwB9L/rVvn90QE5IYIcUy65I7xwfZ1ah8g
/EbGgckNE6NDQktBxBVb81qekjClZn7ECzFHyI30mk4nlFD3leEXI6WPGDAMt+0r
NPlDiNx2wLu9/CXm+BEeen7m95jyoJQPFt2NJb541nQZt5T0IDwPcxUEnJOe+FS8
wjlqnCxxYCvSaoiAf6C3NoK0JjLGqBSN5gl+oa3uISiR/SR0zDwfSVXUES6SarYq
rtB+IkbH8Rsdablg5ecpXDv+qMdLyUZRtC08ti4tdSjwCLGodxkOE0kVy7fF91YK
qostOqoYiU5rd6GQtP41ocBviHEw3FcGuY52RaWvcjl0Z0S4dDQKoRe6jDbbwt6+
TByOL7mUam7b+s3T7VOqeNTlUawNRjdUIGms7YS4x5PnalsNx2UWn66CAgC2ytgo
A03NQ63RHwcmhC/O/Xh2k11YVVWUEzMdSpQw4cSvjx1uezUZQ/Rvo+N3n8xI9zek
bCeahzSkUBz/nchovXGNAgkGBZ3T3RmjegxAoVuTttrwK2MGLyZ4BGERYYQXs+3o
CAymEg60gYAU2RG6s8HEpO0uUxR3k7+76F5uBjkVyEMIAwaepgnGY9X+mDhuIvjC
RCfnR6bPVx7Q5TQX7SCLTn0BFRMeriUzB5eNTSwYbiS4zCgww8NjpOwdBjHGEg1k
U0l1hXW4T3L1J3tW6L4U9dEAxnGWT9C2831GA611T0gxf+fX4dNjV84V+9VH1xF6
WplEb9Paziawn91QoVtHTwYxNibYo3Q3iCNRZGJv1kBMHpy/4F5yIGbkCG29F127
6Yz42QTDRYY4yPhhpBHl6subxT5wYB6N+fQ0YHMgM36jshrp2+nhXsUy5Oi3Ke7B
bsAVPAD0BdMKlgIYHJpWfVJS4wNu+y+OIxCHfVcZDlDOLrTiAGxLzcJjKcS5zZvj
XuAvysKwu+4whub8zG/tsSjOqRX6vpPJwxM8PH7OLRTqWTulyzaM2FEX69gZaYE0
UxZ5kumfBe4ZFZ9a32O5ag88yprJpK7ZliSBM5mtfr4yEWsNAOtWpOZoTJehAOh8
SDF09PGuWmXVpC4C9WroP2WOJJhV2zRkwMONHozVgrSBbLyu6ORyx4i8ECUURoBj
Ne5JJcEGQ5XxK3SCTAP38ri2e5etheZCtYPzPJkonDuAsXFlQ+zPpSVaHBLsIyb+
rQIRlcpxPr6/5InQ0LPrj1bqX8nKdOS4NRqFRGI+fbouRCnlHLDlJyvNN7am3G9l
f136bec9CwKY3Hfi4fMaH2Lipg9XzwAbnv3yRRV184LAdU9jA9MCg8Km2Tb/Ah+z
+wIWyuln9hZFWeXN/QyBa9ISyJmbqMAf68Hr+lX6K4DcGF6Xpuv/uKT6FXIiJT8i
MxGlxwfn0eSQxI0TvIGoX/ngpG6OHRntyGT08zst8EC2hwzs/ajiqU0OeHoFaeTp
2+KYgHiH4unkKa+da83NXc0dGzv2L0c+Y9F2bRO8BHd8pOROdqpsg3vSYBtHPmz2
iB9xHzB4b3NjnVtyLKCZOtpYs49X7zJb5hMb/j7NBoLvsTe+EOKGDiQm1EJYj2uE
LFIE2Uos6ltokI3jRTJHgOgeI7P39FzMzan+k0ZZLF+zU6EzAcMgIr3syw+cdI0s
rhgXfiJhfnwkpaSu8FInJq/puWkbfyAEp5aKdDX3b38z+hDF/YIBM/JPi2YPcZk9
ujWkuhfySTCf+x/rZrqWaw4vMHNL1lMrfcTZLyuifoNTIuauSjW+yhJ+EsmehCxX
t0H4cMkb60yLhGq9wCyqmzb3hUMADvL41tfn8IZzRfzSGo03+l6QMuIupsVxcQ9q
ZMqlCr4gQqYUHUrxEUvGwEh1BNQdTLYx2ayh97pQpFRqPi42mtIM5+90azsaR1qE
wuCbFdTtxiX6wCEsr4ACYYbk3OKf66x2j/vXEBAscyi8yu09rt7GgzIQT7fCqRM8
DFzbKQLjnLuhQINuA3wxiQf9wNIbdHcIC8/ajsyuO+/P6qGEmIiPKDOgttxdUhIB
9pbsqdJ7O/T18xo+C8+pIfGlJ/LwLliPK1FfCEfJ8mueTiVXj7zcsKypcHs0ss4c
C4ICKI5pUNXuqEwFm3HKtnby+h22aPildCmg3yAHtl4eZJeE+fkBMd0lvMwMS2Ci
tDbvmwa3gttctm11oTeW4gDYG/E0fcLXiwr62XD2jnkv+FJoiaxGgViWTz3IgqpO
MqxSMC53uRaeH8FLCoOzfvdYpEt+1DOH3k5AEt7G0nX8Ixn1cxHSb62CaYDpkD+C
ggtE2RSuKHs1MQKTI49H4eTKIpkYGmTdvcdga+ZmQH/CANUygmi4CPR6/RfHr9wm
GahaNWIfdWRGdH4nGfzhnC/nelabqZqFo4sFSEbQskAJffeca3A3nOmPA1yt1s/W
iCowpONTAuGgXWLuLSK8dl5q/qUgIU8uWi+wWox1ZD5+tt6j1X0GpwY0koK6rkpE
yXUlpPZZ82/HWXK9bmk+vLPPD9C3xP7ZEcIJr5E56FhmrXm4i5YVFmcfrq7VmnI6
ThJRkQoR/7rnvoM5cuuvQc46JoUyfly8TWBHnpbf97uqZRFqr38EzDFZ5qaGNuEz
tfVLL23wa+nU1a/MGujWmOeo/r+9Rndd+mJPRMjVJ19bxlCfdEJsTdI8I0lEIUd7
TKbHocvITNCcwY9NxdnFNgnGwvOSQK0SDb/ND0AxWsDLWv8btamOtZlLrZD4XYW7
a03HfYVw4FCHIQcgZQybAYMSN8GNHY7oWiQ4j886s0AAGdo9IXSB8xy24Yw/R7hD
4cGkyPib120eTqnB1YU0jOkJ9J2KQi2xvudJxPqI+vT8zgBNkrDbO/VNGacsJEtH
3DTf68tCOvnhSlZPirigamsie245SN3bD809jrxEbTX4bbTMrVizxtY/k8M2ea2a
s/x3q4vq7jVqo9xOuay2Z1qoQBJsBh4mhg6RNZfAdjiDhN6JLqewdd5tUhIWX3js
WnAU5oUDNzVTKBAh8fOYwlCBjyrjIboQeGcXoaQePAGRImFcK+dZ5xJ2MN/g36w/
kVc9MbMEjuWorWs1YcN7DGkA0Jp8bRsuYawA9CSxkb8DT9TRbb1WmNM5K/8VSyJv
w5Cp/GOEM+85RRc4/5Dy/LQvH2ZiGoKZn1B4LT42UStzfRszjhesc6nIwDL1dWJO
5v+WOz/4rk2RjmS7e2XsjMHLHOrOrP5H6RBEwd516Nsg5hpEvtubim6JseqrJpPO
9U3VYTu3ihsSE4b+gJupfOp+PFBnO8S/hwEK8h/NMgoTDBzwOUJxpAnM7xu3iS5t
Pn234ZdiaP0p0D5t5VKrTB2mPJgBUDPWAlsfsvXkTCrI2vt6f5B9d9CJoDiGHgQM
DNOzGu1fh4/NkI/gCfC+LbuweTqcg303pxz4OS9u65cIgw+b/E0B/npUpSLn1Ytb
p7tpNZ1HOPe8SvEFVwrOZskPP2AkA6OquJttmPkdzYpUh1BPXbMDEc4xnjE18cl4
9oD8h6J+k2qBpKs9Hm2kUZo+5Mnzbb9GsljbMPS3q9G1bkMvepsOC7O572k1d6bP
+wh9Y4tuEp6OX7kN5ih8qiVfqRCzTjdSs+1kK6wZtgAsDdbMb/4rKp85G/iB53rg
8pegFKC+rptYK8IiZgcVLeBtxRV5ZErCk5BpHs6pS0W9efRB+ypDdOlwL3ctyXof
wAzzwq5AWhIfjskay8WYwXmoKT7enFHI/nKWhyq4MHTWpxMrC5d9btnVMJ3kOXMw
VMq3zJ/OlvlGhU5zJNJXAh6AzunmOgMhN9VkjqIAAK8GCA4ToFVlHV2R2YxqBzUf
zHz0xdY4IG8v3KBeLoiuECA6KURlzqVyUK0mIBrz7VQ3WGFjxl7gO8xCQF8rC0Ai
KipgjTgCMJ/i7JT35/pkooom7Trnpb45T46lpiG4aydJHkTE4LGw4juKX/1Cbmna
3RCANfefXIHc89yIX9YRGrrwNOjVccqnOAk3xXX+zd5CMgNYSKR/xOLS5d1JPaWc
prjZ3a1gZWKXQO2l/8RN6fV6y36fPyJZrS1qK7+wVXswCSZaBIN51UpCE6cXV99M
3ND/PFuL5GHsA/Qk/xQYV4fY7xESgJ4XfopTg8FQtWQRVd3DSph6a+MiKzQniwkV
f/Xgjmhq6hHnFxXMLIIIfrfcrTM7zPnbLw+XF/QK3Ds7jRTfqGnkj46Z73ZEYKGA
VClmiZs+yPgPGA/Iy+9L+MONRDHeiUPcoPbX7phH/bw633sTXicXXAGkZ6yEk/aJ
rItP4qmq/rgJlwZFVSvxAy5w4GXHzl7SKkqCocZMQ/2Nwzret2DualdkWHlwS5wS
OrPqmgB1UAWPUamuesydVRJRM8OR2HXsUvEfr25SyBYE1pZHpVfTWSIuVyx24E7o
6PkWbqU7M7qst4vLXeNXOKcpzm0RtdtiusZnZhwB2M82+QNaB76h6cuGHPmVZYAu
Syt6tbKtQNhv7M6ybWHxxq6IJL5CupanMzb9IXDrzhj2/fcVSWNHPpCEE2Nqfr+t
7bBg5/p3fRiDOan1tiTHnB+rlLKT8KcKCRsaRyV31vL58bYoy4wmFkktcNLXKY77
1H1MhFQEaJX/B86qGCnFL7UlP01eoekEDkL1sfdw8CAOsgSAECNfAxqCfngHWxLZ
jrLRChPozCq6HDffIPhOxuRLCJU8p3LHKH3jO0QuixL5tlDmouKG/Tp0kea0++uF
yL+Kj/Tm7KvzfH2djoXCQKS+OVJ6ROf2IIFu4lWnn5QbjKfTwXZVsGpyLTcrXdY9
tVSdPOla8dU7dWqdyam64p3VgPdEZrpvF9+dhtFg311rTvYno5ImJSqQ9VgVyO8C
KSkN7D03R9Ja2ibSuf99WQX86f5qenHmQanpdiJ3ND0Ib/I/r/5EY0E5qM38PiIm
jCVwb+nkkH5cG9mBn7Cz39cBbJqeAU0vpy34R1cX+FPxNWOJlNftmHqvqKNuUkFA
r2bPI8ziaoXRbcQIudLWhXR+GPQbsQrxLnavZ6Jz2t57YML68JsoLh8sjYccAZnm
11kAyUMeBIoTxzaXXK3Brf2RKwI1xciKzqtBF/x7Lod093K/uhW8O+g57RI7QtwO
lW4482dx4KwGx4cfXP2DF/309sYzI+iTyNAqKdEcUZe1EByBues86Jqetpyx7hhE
YiOZbcrlzGNXyRO6XFBzUOLrM+I/zBDrv0Ev18iLshMc4JjE+ppDtjUGKcSsGIJd
7t/NLbeg+bT+mvFT7wUdPtCs0nGiCtQbJC1qpwc/9+PJWeEpLnfviJoSoc/y42Ao
9Vt8PNpd2ukYYjzuRvc51qkqiqtIVb2cZllpvJsQlGO63tH6pusxppTlgFeXgXgk
UhT6HbqfdSfGf0tnqj+ZeYNym1RDQEeVOP9ifxgYg4ut47xxzCNFHRa+Qdcitmbq
iO6MITTK8qleMAeTltppXMfiQ0DJHwxTuM+NIg+e4znoFZ9RU7xR78Fq2irC5mLF
CPhOQdC7LQVTttPpuQyHx3iESJ2rHwRevxeFdiAPmHwhP20v5vw3WQWHe/pla6IK
lOC/Iq7JwrH5PeEFDXH1Q8+IShU1CmLJ+UdtcOvVxXEUGMkyxlCSsPBpKN/W4T/+
osiClhlR324kzc56aQtsMdFe1j442BLQaelzOFrD95ZL422Da2BanMNCw+3jHk2L
XnF4HY5SCZ8O/lxT+DXihuNm3ibh1xlInpar1R5oOhYGMhsglVLS/gB8cMbUN2jF
HYfmxbuBu2N+g8i4i2Hztsg6HS6SQyOX1TRDQgr66H/rYXnSVzruLS+tW8lsVceP
QHdBEiMTA9LNzkNh0nYDLRIlo+LwQZrWjV9LQEIMJl0lM27VJ2oOpJIE6yr/2E5I
3/15PNKS3cdSK/JfgGP+rE3ZkaAIQOz/sM8TV05E4uwhHDSJL7qsDPRYPmVx3oOr
wYtxIkESOcg5uf7QoDCAh1uQx0CNNLUVTRRZ80hKVidqFI9MeMCCqqwQkyOTYu7F
nb5l1pHDfoipce2n72nbdLIfxq8VMek/+WhTIClpg6M53kzrazyrViaIaZL69BQj
cAcKEzFuNC1z0kjNUQRnmnjcEcy1NHvPJJhxP9Vv/KdiW2yWDPqMQ+HUudFU2/z3
N/SDArTibqH5RK1VMTu+JQIyP9vLVh0N5Di/dg0jXMBc2fUJqvx/LhYToJJnKz/t
i3flsuqD3eNzOawNR/UxoJowaQxLnt+QWZBriYwrIwWh19mKD4a774eKGHzuX4W0
F0M3layy52q9zJe+foNhi9G9saslYW3EBaC/V39nBJ1xMID8tXWkJWh+m/O2WeSI
cZJeylhU9FCn9jc+zgejOh1+7kU51xBH/UWSpeXMjppKd3UXUvIoJixf51lvoO0k
b+I/RS51pDT0l6ZNhx8A+z5TgUbrPSPEocdsVkTBLrO2SbDdLeksKAu2GDzKfiFt
UGp6yDh0MeAdGNqNjHApd4OvDX+MRqaGnqWc75FiAPYq2Q6gusQj1//HmgXu87xl
le8auEBRGABWoVTaMhnpapElgsKYNMsrMBt+d4KTUi0Y586zCm5nZIvGNWZlirAD
TW1xeorra5Aq3fK1y4rqzxOEJv9WmqxJrButihn2+wq0ilaLrNVcKCr6NrhM59aZ
xCX9IsApITUaE5OGnxkFxiwwqP3nqoaOyvh1XQ8Lln+0lnfWXFAqalLxs62jBqRa
gR2hcyE/LBEhok3jOEUmoXrkUE1KuTo6RtN16vvXTVymLwHJpwi+I4By5lo1Jr+1
mSWWKvn9JyC7o/sZxFWQs3Nj4xc+6tNtVddy5NYsxxcOyc+RQb8vqxsGQPmg98Uh
sJkOUCyqnd1IKc1iQMwrCAo42iL1Lc9kWMGX9GEyYSVJEQj03oKzOjkmREKl4O7Q
gPx2KvEicYYdFQ7q1l0TpTCUeI3Tg4v4f8Etl/fl8s81fbfpnWTodIW2LeQEZsOu
iEoWDWDSF/444iwmlV/nM8hKBBs2Xd1F/89HcuQ+I7z5vZgzCCrywaiVibNgYhpZ
ZGCHiH6BtG0kvw/kWEUqkiAZSFTyTTgv6dVs2UbAD1WhWH3VvcsMe9Ka0c5KFc7q
RyiszJjGNC1wjy4T4t5y2WeSwKvoIJeAeJtECfSq5XZ5RfZAs/HzZypUyw8DO8Do
6HKezuMqRx6lok/Xw5ks8ZHIRAnmSMK+xBfMWb7zdL/k/J9dR0Lwdy09OakQqIsr
LEfl8u0Hgkxf3P/LZNrpl4cNxmCOrgtNYSCmdgndk8dfrPf0M6A78mHDmo8WatX8
b/iFDzKWwKzb1GrgeEYF+EvH1vgZzw6G3kAB9ebCXDTnCyuq35LDOaklw1R8pH+D
Sy0nV3Vob2kNSjyc9Jmm/X+44v/QnMvmxP2M2W8uE24c+ZqglMHP71jkYg3cutKh
KKrSfa86Mg+c8F8XroF9aYhqBW7cDOF2Njewj8FhDqLfa+ELH+R+ZmYoPbPB/bD9
sDU/0YlP9Hs4nT+a3YVGJYrAZBcB3rx/KwqtrnyV55WbfY+hlaRjKURFnx4x3R+c
ZEZDDrpehznNvkhikNiLOxnEK7el2UOJSgO2nlxRQ6bp2/7iHBtFf+GfBSm4NB9f
z16UxmCPH0vemy7tdBSbXGa4kqYhuiFLApWLPSWGQNYlLUBjx1mhF6LMuQ0FGObZ
F9urVyxu8zRe2Q7G613H9e4/UkwoXu5AVPzTvM/ilHSdgeRmX7HgtooDqgN38Xco
RiOueSVravZYtZ6ntBM8Pzv91ERXwBk+OCMdXsMvGspw4qzIjNGWiLVzYXFbOdsS
5a2P1baSske+ODd5x+hhiZjYc9Uz845Qu52BRXzt8ErC87zVEYXOftcoqLe6KvhL
nbE5lOzGUYVObqOQUzTAIXNNTsOVrdFpGC/uUdnLDk2P7lefepbOtpizDGvtAMDv
EoZ+Zxdp3ZpYOWvpx2mqorbHehadOh8F9STmu6xrZtT6aWWMjgPvCBzTgXqxDkcV
U7YFQpieylhRkYG6BpPtO1SiYQ/KvLa6tf6OWOluHFVt6Dk0iuBLJhcP/BoSKOPk
T7h8X5E4JC/LZFTQf+mvOmJyrDXL90cHr7g/JBpAhynVrZ9vQbTaGJb6FQsSBiFf
X1GY86ntWU9NpfSfMHeyQ9b61Ed7kfct8gV5e2W87XyPvlpp6oMZFE0JP0sBqDVW
NfWZX6qQ2xd7c5HhH2FvkeWzA7JKZQ70WyAwf3oZmugq2Vx+tDukL9wnF2iSc580
CcEE73+ABj0+Rm0IRTrJT8a08trOAyV0ynVYjO4Q84utm42g89udjfYzPZhWmJsa
hnYtZxQRsOBFvlsEAvLoABN4zsvhe5a1aTV9cs7iS1IqvQxzC36AWkSUfHPb/25z
iPL5OBgsCC5NBzZFw7rbwU6vWQuzh4nTMKAAXA9wi3x9Y27Ws3Y2X/pQ+BH73XFM
OZXk4S/dLWO8HxdouZXgBHUDabGLKPBblQ+qtt3eYx4Lns5yBYYjdJd1puR6uYsi
WER1BFhmyoaQySypYgwWSjvmdr8sSdnwG++hSZHKoK7gYf6/k1cgc96TTYIHNAg5
qpoGchDdkXraLLPMxY3aXASt3BiLRq7hQixLWTD44SU6kJ/QT52LKZoEoa/Ye0Zd
KYck9mWDcAV3sszipDb9wuVO7+Z76BOIIiZrGyJnlvV2qb6wURPLmhQyY+5oMB+y
xwKNHFTv+kGUlMINb6vZXOGPMz05eVjyly5Hrv2lH1dHIpeOrxvvla6BWVINV8nn
XmnRHWMC7V5slK/QQwadiwqEElfLEYZ/cxrcnUyBnrF6PzqduK4VnMX7dN308PfL
sjTczbSuVBO0/gkAW/QO+LiMltzfkR3ZmB6jRM8TcSNpeuUccU1E2rkppCI2p1Bt
/UD+ECi3h7+W/0IC4jr1D33xQBv0LzgJMjPzenmNObgEZAN5W6ONfkgJw4G3nnJV
/tZD54jG/EHXwEJ3hBrlOCpWTwk6HCJ94F6yOlezIMX3W/trPW3v7BTm8GFd2oO0
beInDC/B7Ghaldv7Dol2VR6VWFIdEBRp96n6hTFhe3I/DWc1mLRPAtuPDRL7JL7u
gzBI248nYDKDwBXLb0DsqByCb/H4WpV6yBwE+q7TfSyOdSWF4vxVNAVLRniZgvRf
e1kn1VbIIsBqfGA/FsrYEAEkm4SBXt1z3bTA+bX1bQoQltH20FO/VEmvupN/vN/u
c1rL+Y94+KKsIwHy1K4sbQogtP/QfxjhZLxMBTa1g2mziuNGdrl0fwCnwM3nCVOq
qq7LIjmR1TjrIJblhWI5/mK/+KwZVkEnbZyvgZyKX7HHxEqYyndN8b1AR3m10qCT
SSKPwzu5lXs8HHyisQqhSjnR2ZyNiYVf7RofrNToSLcOZBOW//3DJb3Dcd4ti6yr
QWQNutYO3Y+GGCMVjbwgdkYf2M/FvVB1RfoygZ1jIvKMuT3ky5kmXM38DKm/F2U6
ShDnuGpVkiI1zdmWr1o2yqdFbDHaTPtcQfAQDpABYt18o6WVmB3qRF0FK/iKx/yn
Hp8WJcrka9UTHrsr/+lNijzfcX9/Gpi3egzeLIoR5WW+aBJdLkBSKHK5iXojM2SK
vXMjYjlHMX+YkY8RhnHBR0ouDBEZGPd9/4L2L9ISMFRiU8hlcjH5RwDDlu9yT7Uo
nw8+8gAF1s0Yzbylu0gNz7Nk2nigDli8M3r1bhXx7YDIiinH+71G3hhPrOmxL9Df
ZqzR0NPch1DQhX8LkO7emtBYUF1qFg6U/smZBkjNydLrrvDDkZ9zOsxYMs4WMH/x
nB+N2k98WTPPo7BrGmCjoIhWj/ILikvfl9LP5ieK+e8M8cgyp07/mKkQdPusMv1M
uNMsZl3iFKN/b87avs187/7y5uhx7QSAtBcoSViVC2BOMJ//Kz8cBO5uR5O/XwPK
M9kvfpzzvQExCyxERUNqFXBeSRvZTWiIisa+jLAP86HOhFtyjAkqMX26vFBNm7lJ
viPlzQLUxi94vYTe6FMXv3Z3ULFaK1zOTeysOmU6zQ+ALDv1X8UfXTKmDNmmD3uT
Yg1fulv23IsfUT6eFxjjygZmJnQ8bh1LQrTXovhn0tqMSgEnS1k2btXHIne9V8Ru
UJymzJ7wyBqh5EbaweA8L2L7s1G2qXiZiKQt4/b1qrNvB2BBPMnETqgm4/B7frmL
UW5x4pi8zTxW1mxzyWnptsTHrajG2MZyDyE5YWe967he66oq9kWImMkgI4wrzbp5
IwsDLtK2asXDIzZE21OcJO8jFcQctLu1ONsgqUw5YlG678O5cEvahB0RkrbZu0kE
QZWNEAWzyS+jKQbCQ/qam/ykzA2kjnMFI1hCCqmvI6pMP4AkIvqL6LMl2dy0EZ49
CCwREN9sPHqD3VjENadoM6V6xZ5DAB9Co1DMjjgNMqf8DwMcdw/ODtEbjHjFRgIC
YqySDYtSBkjRpEvzV2a5aAXEeYtzfebJpz+zNpkI90AaO1ST1Ir2Bbdq47xk6OKC
w4KYxci/0MLnRSqJ3Bgc+xQn5+dXnmmaR631o5pjUv0dKPkmwwEdUSyqPsH3rIlv
NRIvazFSed7yr/UKtbF0K9VLUGUn2Yt4RhU3LIV1MxuIeeqyfQn9DiEH2/UeYA3b
JNahND0EjOvjcZCvclSyKr6BCfIkAwYbeNm6OQSx3zsDnkHASNZPj2rXP1YNSYXg
QZqaTXaUxpNgKODFMxz9L6p5V5VtPvCr238APAwVmoWXYwTLlIQ9/igpcU9JIjS7
59zoj+PX60/go//h7OGKhB1z8fIn8rLc69/H7xGWiPMFVPD02x26AysM+yQcFmq1
+eYC6TkQrImfl7Qz9PV6E///vsPg6aXUVnrmHHW5eL+e8/UWHFtmMUZBxHRHr0fZ
PK5jCeYpzoJJCfin+zqhb4D3SUeUuFBerXrdsNJtOCdtcfTiNU7tSakZcfaNdMNX
1VlMCrN6kc+wolbzc0q/zzz0IADOGty8rfl1ofKvH+2crhdLRBIXPoDoRjMzeorb
ZSptzkq0EOMlOwcMuUPCmIUwxEWhh+06h+TCI6IzAHxBS+jLarVfgwqcajv8Rc5E
DPBGmqYPwvt7G4vbEfxN/kOYwSjv4Wu6waQuh0DWHf06INTIEu+8LIDIPNcDohVz
eocWLIGkHc6zokNzQSnv4nFZ1OxNea2RHtqvLCMU2Cv7gpVv7VNobboPxEM3e2wi
MahaUpj+IrMuLPRToAzg25Nb34heAEYugRzG5qcH2TpQFWjHvuuRqnkqtqkUrwgg
Nnno/+SyMB+e533ZMhPUSEFgJRcI2nZZRqnqvs7WqjGED1UKOH8fOQkZsHq9mT5Y
i7tR/69kEzXLcaYZ5YgHfji8Ck71cHTcfjiHf4zPBKubmF54eyfUfEBJRj9DL73t
91yJZl73O2mhzjddH4F56kX9uVDnSMJalaX3YOQPDPAJM/+IZwfAAChew4easg2A
QIIrcufHSN7Xk3cMqskcZxdKuDhGkzcv3mlKaX7kqW8k/WcxaKBjswpxoLqOm/qg
b84Ycz6HsU/FMAfY3uGvo1ewsin/4wHnRIxM7DhydX0BRyRnlZVb7R5Iws6uqQ0x
YPioBRRxmJub7E2Ef0y2jRMI6wgAWZQTWToBWZrtV1fE5KdBFUVDgsbUT+0NLiPP
Vpa/reKnAsmdbKjSZhpeVOfVTGyhcIWjJBS/Fs70cv/N+18YEGO1HZTWXwxhPi/X
6qaIU6QoHX7CaRsr/yKDddTcHH0tkjeC9FbYs20oGSSO7aVHtFKt+zh65cc4QveZ
9sZ7v0VwuC+HBP02nUg9fTROUT2DwRoo3gZHAh7YnnxmVofKkYuqLHGeHvqId9Z3
9N0EA9AecFdrOh+9mqDGl0EZZBAyYsEPaXZqEgTJceqk7bmFQ2ZiHDO67YryaHko
UNz+X6osldoYlFlYvXyqko7DyEJEMXtBgIN0n+bc4anbkDKvncmCShewJoZdVbiq
gamFsQhnYhp//a8SDM04Uo+Fb/p3veeSwa2u2Fm+H6a4lUj8AldWmG1E3etIwnJD
hFxq3cJrLNWSm4Xdhbp8EScBbNm7WttPWqjeozFsFLPDeQURAUIOqznF3hzt6yPy
fKSlJWZs3w4CowUMcr2X3CRdbPeVUU6afjwZlU6CgRqtYx5PQka8yZgAVuWkOpvb
rGAKsDFkXQu4svazO96g2jwZ3E3eNz9b3twSwPjoX4JuqXP4PbJSqY1j2GsF1S6w
eyhcGduWZN6XYWbN78KbTcTU55H8IAoTrjui03kWOtGtDf+exoscgAuPehIGVIe6
nO4wTlMX+jluixU8laGNyPAP2NxBTQnEYwaqC1o7N/sGFXdanhETdDNzXH/v/Trp
RlC3lTb4kAaZle/mSsmiqcV7XHplMb6nbxPweqspssJ/3awZFh11krKMeEkBaZLa
zJbDhBvrDVDyU78Sux/AW/n/G1jN1FVDK+I5mlJPA0dCg1fWHJTCJFtz8AY6zcDL
JBMageg/HXf81hKySpwQrwGzhLdtIaXfxHX+eSuLDc/fYBVB7Sa0NpJhntpWt+Yf
yn33Ksws6zZHxHfRCr4Z8nZ1FRPqYNIyO6UqlpIs5BqmmI1m6vMlTH1FW4tooB8W
norHyx088dv/qbYPeT7uu9cuCQpzaIcv9FRtYCtNCQMhxOnBQhuMTad6iVvhqaia
Ta5wcZ+oJlIr/NDEsLijdzLQfUwKHWBRb4mq9mjw5UuZ3uK4nPtHbPqaYKqyb3QR
T6PJl5KqWfDZdN3+x1EKSvJKMDWZOwJV3jNVFoBxIdwFOWEJEROv944+rl15ncYV
Ep/clMrsJhyingKGKLE52EtfhimMFidP6zpyzVvvPyK/Zab0JpenbBtaKAKK2TLt
3pG+a6D6N83AXilZCB7c88wqJfdINqPjTXNDf4HTZGsMaGg/DOMxIY4ZT8CuKn47
aWXu6iWBbJ3HqOzO2i9MPnxfVMzMUFAOZYipT8Hzoadzb9lg4wndC9B3p0nh/ZzS
xwLn/BYN696MEfdK5315pinBsOLjSn+SBFJTS4xwi4Hb/1N+8miCxqdAE5LszQZp
X8XvK93qFXg8gGGFOngHkOY4lROR5Act4gNUrN8rSLVc0LKD6V8K65m5EUnKsiwk
PLNmh+cQaaE3Rsq7xnjrXeWdIU5SuHmMOyqMBwk+mtwn01SUcl4or1VP/P5G/ScR
j++P5RpgvRf5YAxgCECVKU713+F21vTE5NhQwoTo7ix9uFcQH/G8XzBbalvYatVk
G+GmWW/PJxogGquqlcMD9AZrkLVol8u/IupxTHzf72tRLGV5OfUU/ow5XIMvUmdN
iXJJqB3TnBuShyN20LDdl9eJCny1XnGMUqOLhVtpPMukd2OM65zRwjbKr+r3rADh
Or5YcQuDy1aliooa5S2KPGhsnd7RygLbBlHhV9NE/iAsQNgvxbp1XQYXRzLNaQis
/pphVqzWwptQeL8EaosW26HprYxGo4RoUDB/q3i2yss3/Qcf1LxSbS2WvdgR/bdc
nsxmxq55FPf4PFQMI3TH372y2kbQJ8ug1BAoBE8Efs8LfvMijsfoWC6giRPb9UAW
fcWPCZC8pEZN8ieBQy0N2mETYbetYv4vkdk65vMgXDd8FWJGx0dMjI/uJz1X7aMO
MbmXK7NmTXDDvC8+4LXS7CuumtIM1fkzCNUF/mUAS275jkWiBiEKlN7lyO3Obe+j
aBEp2dO7aPMg4t2WIIsCMsRWlqnOfJMNGox/5g0mc2oqaKbfKAHAIFnJp91cd2x2
geYQ/aoiZcmaxIfQE0Ua1x35PIyp5VrwbWBHosSBnszxVB4YUu1LkOdS9DTmlAuO
fNSAA+FwUxpsySX3n8/V3gw5JgbhqNGsATKB53M9aMInLOSFWF5gqNSaUvRrdzo2
sKuoOltg9cc+Aa74++grqBmRPmWV4LmGvGG9N/m8nl9jo2vdESgFj99FI9sXKnF0
jDY5DbElTUiDph1BB3ShXRr/EWoyqyeoFHB4/gKEOsUttbNg3zsNlXDA0l8rYZE+
GR4L8L3SrFyplZjD5fTVq4mR5c/Iuu2xxhe0ghikPczFi01yiL5xIChZbfzX5+sL
AF4+E+YtEwGXREFCJpf+hL2cgFaSv6eo1q0KqIF+VDWdup0y1aG6u/RfQY1rjg5l
Pi9TQ/yXICU4TZdY2917xzY1UYXaDXQhPa8FNKMP8JRQpWbfdh5BSoJWTdXhvI6a
qg92cJjfOvNrOhr36EHvVZEYiYLAErf0qc8IQUGbb2pSc32QpwTySGD2u1YQ06FK
Yqh1AtesG2X8AOSHptMDMxYEqJcoAuczAW0vlYgo/Ivx/gGr5yRBzhykEfh16feJ
ynHsT3tS8fnDaz6DIB7FVQW0sFFxWJ/UIFMUJkn+JL2/h4jn6St0Fqi7Jw2oT3RK
a+h1l/O4KGVNahQXFbuNpjopuBgKBwDpal51QwzFl8CjPOsZGPdCutfdYxj3NHAV
Bl5fDGf5VIffusQ4kvL2CGNCtbgsVyfGM1Sfm7Ik/8ciJciRQTeK6o4xOHc8jt0d
fGtjYLmg0PBbuvfigJ/xqtkSRHbor+lPQK1czMTqUWk6BIFoyvKDCrPT7Y7GBhTT
QfyXwavXoiPpl2443pw0T9qhqILb+DgSdI/MCx4NmR6Frulq0W09YU+ujOitGI54
rC5MVzkvBzHA2PKzrn0eVg0JUWzUR2AhLXAIzcWGTobBdLhtW7Wht1tyP1yJzRKB
OE/JaiQb+l3K59s698X7IeZe2jt+W+zRo4ilQZo4hSUeI2Tq3XRWfwOAXWliHkRX
T/9HTMOVhnF+r0nD0JZw1jEybuWmGYNemdLbd1+CTKfmQkL+VwybbPcj9Akd1/JQ
rzmUGqKyiJm307Xf9IQJ17NwrlV7GYp96yI+L9YYTFPq0qi5dy9cVpZ+udryklZc
9rQr7cHMYQ4BKf6vWQnmYwTXiWdzi39PKtjcXb2glFTzJo0dZxrR/gLjKXlGWXjw
R/7rSD7kIbdqKxYZTQoJyZ/ZvB715RcXydWY1zK2UVQ7SNV3xIKDlhBHbfEVNwvt
//jGGMpsHy3uL8zhL9LT59Jg07x+pb2rhC3Oflh7bEtlRuMefoEXdo41SDi6U6zs
3iZkqKBWOOlrT5ji9zkId2mtzEPDU1cNoI8KLAxOL7m60dAj8PmKKjqnFr4NgkDg
nIAhVtQhXLhyzAvTA0RKjg4WIUsxtJMRj6OyjjkPUAmaHaoX/iS5bBNpU2eYF+yN
VgWD9qkeQRKJvPbKxnrc8y74xFMgVyM3uDYlO3LHzmi66lp7I0jMD3CUUSx05LFt
g1kYcwMGQJSolZNNABZu2HYLING8GJPIldiCeMMl9UDI0bYAig4P1sWYual+/5JW
fZnAAooSgUu98nf8jv+zOKiEHBvU8lrnTq52S1oK1l+0xhXiCGy+1fHgT3HkdzL+
RExJUQaIY8HsZU74vAB44T5UhHf6rKSrH2COP34zUN5EJ5B1yf9WRoVihoXRU261
UE84wkPB2aHDucYtjk6lnHd0higQe+wGPLuXvRhtkSyMxJsrRtBqMRfF/k3OpeqN
EiO9ARkeRT2P/2PjybMvyKsUYoilrA+Cqvd/tCfgZiaFR09WzgLeK+r8OTYCnoaK
xBYIQSJBrUeWdEXZKYIn1ik7AQXrMoiSnl5zYm9asG/Bfqqf4WTM03EjrvwPBlsi
0Qvsid1/+V2Z4QkrgXqh1CoVTgg6UlqDi7DslY5hexWcy2oCx4UyIjJpPTUx/bpq
DmdaMDJWMJoavfO4Cht6Hexhm+qnTPViO478rUHZKqfTUyOugwPhJ7VrnldAZbaQ
CWgfhd14dtxqOLJcRf4lMmkgBbOwmrWjFNmWZiQwmI0jbIwUvOFHgBr75f0Gj5EA
BiRgCBOiXIOJvfQkKtG5XwoZ/pvsfxwg2qjAQJCSioRGa4EzgomJrLyIfJaE5HOK
o9aXNWlL+U/Vno1Wnok6bjXmQWWetuMxytwbqwepq0nUvJjUUt2gclsK0YhFjZw7
ietJ0JBGz1vupWDOI+zu6C9+7BWmPqN8vZy2BrvGAQqsWj5VEfGT6hav75tHsQEu
ecW6+wryA8XpGQPRtiV8f7bsgmTtu9PzBfdlcfVtwzQ8xMl99g82wXEhCFhb0VWI
G1eMOrV6M3VCQwn8Fnosb6mScL2MHet6wvny8KQhj06csstL2kOn8voPAhOxhPmf
raC2m/ga7gqs1Kfc6Mi2mguLdtlmByQqqi/lb4rFIQ6RPfAF3RC8wwLJxuVqETdq
aSihPSk9XXOGV4KYs2Tw2vg3j6bg+tqmeHzk6TvbQwHsv/nco9PwNG16RZVR7qYy
egPG/DWbNNn044aJKS7tSqY5j3diONN9wJCqxaYltlHJQ2umCUDZlYols32y+HhO
YKpe1LbjitRO35LHZI6MBRmbvi11O++6tOZ8MUUfbrWtWQ3ATmxszh6kh2FypFsR
22tZIlxRctK/qH2ytzJCKxcwcMrOE0JPlJx9OeZpGkggPh/DC0UyiEF6ELQ/E55h
LaWh77HFFgEvvfbaMUgoX7+ARo5uOs3KbtYtWDStkglVBTnf2GJW2FNsIikB6YnD
ZQV0tZUuRnHHEGgbi+iiHQa7lgw95z9EKTHV8/6ijqhyNRwW/dzjNAYEJ4TPuuUI
rx4t8SxvlaL64g0WG5Hw4kvOafUATzy3qlJywXlfZo74xfs0WLvK6NGWf6EovKeR
FA2rmf6tIn907BkwvUgd9AHnSlS2wziqUSESCmSlEomYkSVwghmRYHSKDm8kuJG3
UWhzPpGiRf/GKEKKAFsC0gJdhvWOgqrpYRjsIfqRiaTNUg9Zt4NgeqGOm/vPpCi9
Tk2h5YXpu51IHO6GaQQcfnyfHv5YmoV+KGBH0+dPKD2l/cJT4aXXbBDme7aYTJ8O
B1NEFJBUxuY4+s8xQd0yQ9lMkcMbWGxxAJMDVjSRFbfO1byoUlAwF4jKfkgYDXqq
0S+XWYgnxxmebCR3azHmQlfeU/C+XxTNNaw+MA3YJ73bfFaR9nC0/dtIXUeV3SsC
frQ/aVt94432CY4ion+OraBfTKHvZvsxxy/fXZrvy8U93mNCruihrIOyAM1sU995
GxEQf/x1bRNWBDBZElZCw1PmEHFwO/iaYsmywUqtBI9pptwgPH2T9BMsDKmnIbKd
ryPKOODPvjcVl3+YAqoKTQvVwj+7RQleN1r3j5A2PUs2iqkquJq7b9suX9J45SSU
ygX7QLcYFPtmpWa9LsYQIdTTu/NrbZod6J7ypw/mh2Sbb+e33WM2ppfku43CYjen
fLgIGQqTOGHQvW0WLDyOvVDJeoMWS3OHK+YbYYyvJ2XtPl+KB7FVarR+yFnAXJGZ
JsnjASEkmhkb/j4ZNt+h3JtUDN0OlFhvVQdiIFXMgYtGT79BuSdt1V+0fdE8q6v5
V9rHDpsUzVr5E02Vw0VC4LFBhVpKjVkZxEHP/tU8Ulq/uwpYsWbTkIZImZuALvFx
wAWnVCRN59HQkl8E8qVrqBr81SDFHkITpcIT5oh/GjWO+NKFtspN/NP3blx2FPuB
AIrNjFZORWHAxbTNMgR1AzDWH9PgM5hw31D0qUszAYTcj/+P/2IfgG0G73UrbjUD
M2F1HWrbiS0JJS5hecpjEH1/9H+YU25Gjnn3UIIa5gOov3LnGNlvtXKefuB4YVV+
QJ57Hyr+4SLngTsLIgbKOY6biPSOfBOTiCInkGwR2Ll6yd39iuVItRj5jWcrGAYx
yVfP9VPKJ+Wf1gpDKzRLwxQ8Zsr8j6mhdzRTl2buad9Lynr52Y/2jhBEI+qmKm1E
yEE8QF06sluQrpQ0BltX6hc6q0uxZE2Z3oDYBgR+yQN5mOeVD+isErshLG5D2tXw
AgBdb/Ge4cmmrrn7zHtmwLen35yRcBHX0cvKrlum5HmtKbwn6V7E3VmB3UGrMfBP
+m6o85fmMOH6fPrNGWMwuoS4U8XpLioiI8/F3yzXaZbM8HEj73mmPi/7eOPyRsua
6tY9dkLzIwOb6CnoNkHD9vxXdbb51E3Eulh2q9jliuNt84btfahhpXEHoONZ29k1
LbH1iRpWuELRb4vvFsO8VFJMqf2aPwboPZuYe0I3LghQYFM9uuBgMHZqps/6t+Jl
EWScxUMLieTwPS7m6ltLFOqRBNaBeY8LTVmrS4CA/b2Ycftk93lVgIsQe0DbBK+n
FSOGhTMWvgaXW716TU0na6o4eQiQ4rWu4nsOOqgbwvV1hfNIGgUGoZLoRzORNGrl
LyJEDCy7tJssjTQCuS4+Fw+5iy52Gmrpt0X3MYUPv/GqjM48p4JxjQT0q76lqrcS
IEOiXIo06k8gm1G/jAA/elh7QFe3dYbEFbBnNgU5qb0RW1TGQqKFW5z5jlDRzZaE
eI5IArC5jv9WcuMV0kKC9ATCBWRIApj8JQBskvfzCXGmdhZdAXFOHONFKOjX+Yfm
K/BUTQXmIS9LCFylM+uvoRI9+pbgHgfLaXIvhtp47j6gnysxiKWiuu73SAADfSMc
bhxFliulXo2Cxeu64BPj/iB8R23yuWeUgu7Ox1ml08aI1TitflTPl5i2/wMNks7c
n9iu8sTOKfdd9OM4vF4WinNuef0AI71Hho1AcVfW+YxeBaxv0PDNSoUH0PKuJLne
LDxQD5DHEiDVC9XIFrhmlJdVD/gbi9cPW9+sRgTLCFO1fMo5dRxgMV/jwLDC3IV9
nJa4hgPjGcIhqOUl4tRPv1KqlFKWEojX4PELaLESM/MNlm6tflISiRtfD9bKP07i
CJ5zxo/ulCquyH14tqNbz5Aumi1JJEv0masVFS4flQ1OoUQ0QjHiblYFVbHaGqxt
TaCIkeeI4Nfyjjst0ntZ3q8uElVp6HmJCPT9BQ22JxHNA42AT5J3VclpIQoJISjq
zetHzIyAnmIv6HmBzWgON/z4YU4uDpxH7GBrshYEj8yReWBev8a+pu1CJxYSw8++
3v1azKtK6hFWH1tijOzpXpd6VXzwB3Qa07lfgWFUNRaZkqbL5clul9pwnBirY+IP
uHKsulJCIUMd/VosO8fKkktux5eJn3DESmRezYxwLIGY2sK4p7Ablk/ZrZZ2qDj3
sNvtHUtRQqeoCY4ggPPf95Pa2otc137FrMIdHuJNKuyHkri0FC1osFCYlTF9Q6bt
elV4hg1rzOSyPkmD8QeO5Dk02TRRt6knHoaCqphxfumk7hv3SV13GLvxsE4LOuNR
1CTn3P3wPYY9IsB0Dlv9/pMVbk5U2MHDNtYaazDxJSt+uKVShPGCIDCNAjsuMZta
tMUsDmUVNfhpJj3jU6Fo5SEEt6oBq/ra7t/mC9beRO692r/mAQbSTWb6yZhIMTo5
U+vOngfASvUxME9GBS538SCIQnyR1T85UIhDqptDPyx5799nOnFMvq4X0tsuTJ+y
yFa2jHITTc6n2yEKRfyqA3YaoOTWQJ+GVCdr9kTBv0tmS03mGjzAViFXdjiMfwIu
gng4Fahc6vNjEYpHotxl9R4EMHIBxKLTcXkqG2YV+VXdvv+cjVEq9FPpKOWr4slb
2tRFz5JMWE0Qa21L4BxNH6TB350g6mgVLVoXeo9YCcyPwn4abmNRQQ6JZRj5+454
FXwNL93GC5Qo3OPXMw9WozAG09qRU8xV8YSHWxPVYLBDLc1F9jVAnuA3cbVp5M+W
waEuu0jixeva8fDiBB1ZC0fuj5F1kLDH8t5pqkX71n7Wb+HlFhiYMg+UrSaR+aiS
ra2HIHJo0CncGE1m6RDRrqkCCugw0y5mEQMDII1KId9ntqtnBseOXFtkEjSer8Hc
tas8A+1DBwt6hha3Vp+hQF+BdK+jpGDri9gff7m99iY3YAiZ/JrhvMHa0pvegrFg
XOoCfgNSSd8P/dAmIXoQZpeyYcCKLDijsPM8ja9y0PYVHnSvMDuJyhqcTncw5Ov1
5ZRjiORs4msGAw2omU9FUCgtzkw6mcelxP3JSKDYw9v6M8qvog2kJUZQbmnqbDtT
WGd0mQyg7c3WFuyia8c0aQDfGDf8cskVuK/RRDpJdREZvDNxhB458AiThZvI8UKI
ztaKvaDiUgMX62CxCcZsrKI0d/x04IdPKPqD8tHeasTD3rbMbuzqTPdJKFy4TMcD
xbchk3KjecsPCmkTA3fh0QWCEMYbrjS8jHlf3euHUBWTDXappJAlDRGcGce6XtZv
ftOqnSBoegbh7SiOAKtQQkwKq/GfV+Q/AWL6gm2js6sdOB+UEDmRWdS966Ez6xN7
d0VhibTq3wmcGZBBh9getOv5brm/qWCKxnO2u4GW5CVSIk9dR9lD9PYm2UWCC23a
v0ktuSLRprKLotBYz/1KiCi7H30R1qoy740sSy9uY12Uz2LWYH/WnYBf7kscbzfE
hwdwmYbqr21XJ1pnc7nLo1Y6X4va8ClZUx1X6dc7ahqgjPRBRb3Wy10qMTzTuFp9
PBH41gXw5tG3tSjpXw+Y4r26rjnR7Y3ZedhVxp9x+yn1qYpgDRGPz0POTnZfL7LT
Emk6tvFbxCZwC27RfVuJBGkZoEo10rr/BlxMYU7PJzFuCm/tA29yRS/+uM47GN38
aiHJNgmxvhzUqoLchZSp01FJsNLfGkgS11cNXP3WWYIoLXH0KnagSjk2ovH2Z98y
69ZoGp4Y/drsQfWaiqfaJ4hEXiJtQ0vRkldzInghCvU29lH0esCqRGbgIJ3qj23I
Glz55I+HiMnEnltVMhhrZMciN89P2vKwwjxCC9C3zHQZrCJtCQP2Hbf3U7JPdpjC
aW9XfhuyNuGS2UKa5bft+qbjQsbhflhblwyiaMHNAWNUPepFrWoGzJX4XLxpQw8I
w+jMLn+WMEDEUsUJa73gFVvui0MrzMzamfLBFQ7EDJ/plLbZ5tygoYWcrBsYH7y4
49ZSQu3vpzfYbjUH6epVsuHzRLYVBfYPMf7mT3ogNaa9NeibLbtGe28bru6WeE8e
ikrU05SNjb5gOQvL3YpYIQiTk9U2yj6r2jI5S3/xiLq73Hi3tssnO9YuUxWAAiVz
uy3vFahcrRkMX11RoPIlIarDgTxS8OD6CNdpX/KPPGMv9L/NaW2P/x9Gad2cYk9g
mE78ZXzkSHh+Af02nT11H9mn4qPuhqOOTWLee4l+fntj6gJLNkpWukLBKRuqTezO
1aWipZdUIOfkOoW0hS/VateEA3AN2OTcCyLvsTsY0MEUL2SYMEeEpH0EkfZXhSVN
W1Cy4rl+BWRqFSXX4NByOeYq1uL4GwUCMe1++ViWvGHp2XlU6amuP72lUgTYIp1G
5n5enVEQFvqXGOSmoBAPJCLlWdCqb9gScoEW0Y8VEMj4O+zAjT4yJ30+v0H7eKht
U7OAb/G0DRPh6haiyyp+fZ6Czdz2IJzLVeNTPS+ka9mCwQEB0bJo46MSRNkOaJKU
VZrScGPrrRY+eKaucxthlzUmQz9xTr6B4YqeBbmNwePETXudblq97KTIuKcmzDJF
KQ2JfAEl3tJyGUrd0vMrGOp2DRkisy8HTKdyxbRp+0fCkKDyA9JR1tIKDSNt4qre
cH5DuCVp1Oxh64/jKHFAhLjMT4Slu0vHt/VtXBx/WxZd+hBGromXIQn0aCgaK/iP
J7/CH4/DgABDorCfts8X28acYV1323t5VKnz6nRaMpIwX8yb68L5EuznN266pHLO
BdT1h5weJRhZdrm9q5PDKDM3HMaRQ7HjBwLdLcF3a5XtPUn1HfyKKfmA7FTPSII6
WirapBuEP7Lkc8pqPq83SP02LbyvcH/vVgM1oK77mCy2P+ZvknH1K7aDNArqhhyC
BCeyvZjctsUcEUgecK/ejRuEBYLKebwEgEBiAp7o68EA/ihfhQFfAGsm5i4XiKYH
DGUMIhhV5UUwwgO8aEXJFB7OZkAD5sH8vqGAH9TxxiE02znO+WkS7jrDmuCmq/1f
MRC1AUkuo2NGxfRHMicgttmm0wODczE7UAejr7O5axVKSl5a4rFfApfGzbnwbknF
hSJtc71VZuAIWsbHiZ8YhT2dXGJIw+if0yuD4hsJvTXhkqFJJnAplUUbmn88xWwM
vLMP/zALye4VgrU9pRBMw/8zYgd2SzuRnJi9ndtisavlytp3O3c4UehPlfjB+Iqb
UiBpGXgpPLjahKaV5FboWw3Fr+VLepHspNoMyNNeva4kEOdOhktN5mIjM8DiZ2kr
RtxwDzMwGMmec1DVNDCXSWL6/abxwvQn2yKE9R0N0AFKXaRwoAm9ZXglAzA77NZu
Gf3HBixv4sXer6aGWTIKGITaA2W+qB5Ki60d6qUH/qLfXN+MDdNwsL9cOpKEpYNH
fyZdag0noughHkxCAwsbkhLxvm7eg/aehOnyAHxVrDE9JNs8mz/CCt/QdgaIrj1A
HiYpGyIGCdBhuRgVQsTwrIqgIYAOldoqYS6Ovwp2XplYOiHS+NBHHW/7y+EKf9go
1GdMRdk8+jOd1l/0uMjdD2j4xUNeOG0AKMDPynz2bBVKpHz1+kxt4PR65w6x7iuF
bY4V5ZLeWA25fvO0ZQR6IGVFOoTxCK+3nU9JOzog0Lozd/6P4nlKKfTz9z8ACw2J
5VHPd9MH+6uozKzbV4Hpas39pyVjzfO2amSe3uTNFLVo0yHCO0D+GAAiBJznLlLJ
fCXV0RZt5b6rF9hM3VmBKQxBmEPivA9O2h+9PzVkVXEQxvfS+76zd/NxPGoQEroP
uShWSi0wPUOVVi3WnaXErNnOJYPsQXwyySBkdvD0mSq+zpobNr/ZO02gAitx2zxy
I1jg+ctp9VLhQvWFbY4kyQf+0PVMuQ2SbZIyhO4vfYeRu+2svBkvGgNCgz7P2H5z
wjTtIwYrX7zNiqFlgKgc9PGfj8tWXbuOJo8ctRqTWwN10jr0KXeOvvTgMwNFtjdK
Fs1ECLVTk7DaE77eO1J4fpnzjQNpDS7+JLBNAhvggMf8kv5i9mUp3gtKF54H56Mj
sM2YzbS3YLKBMmY8vMPkuRasGxdqb/B6pJ5OJ1kjW/CkX8mlWsRSIDyCDg+AOZP9
JCf+AJT3N/Aa50AXy7gJCdPkrthfsRoA9S2T9PxwqfLy0YG1Dd2nO3zsA2HUm+xh
zxNkdNMmySaxMnZPGOuWe9FxLYkB+l6iPWAsGLthJTGQSGvr6Dw1ljR7ucXnTlxo
Pyx+rJApUwBR5W2nlz9aRO13+L+rVr6ibNdt6b6IwcFUX4aVTwAPZQwd4kduXpvc
mytNe3jTiqKZwLwqAKB6bVaPcs9eAIJ9GN5p8oUiiDUqqOSM44VsN44lrVKTZKLK
KH0jQqjKhEbIuTJCe4TsgVt17BULUIsMOk7FOtxKj5K9JEtbN1OckqC43YzMJm/8
0Sp7sZme3ooBJaNkJNNbmf6eHvIT2u5fRIyw+WDh1mscpx3p8BjjlSaxojw24uhO
zJagLuPXaJwyjNNMcuMwI3x/aqYidkWlkOnjQB7m/FoH9GkUbChqefkptUlL+if/
OLETO3iIymKor2rwMoyPA0+7CMUs5Z0m9uO939n8SkfimLfX6J3KRrR0xlVUojip
wfWaOtzOCc7EyNvGvaISFe7mXLMv8j+vEZfgkcYnIcw0xozxw7XYD8VvAqnNtGhj
a3r40pcCcPMaJte1pXIhBJKiMgD/IFqaccslgiTRZh+tp5FU4zfU9+lU5tvseyfU
DZy5wJvRZTiOzVXevBcI1tY8hEzrHK9ym8ZiY0y2J3IqhzzpxiXwlQyFH+nJrIu0
5wapl2477Yp45V3UteZAPkeFkrCAb1nfOna9+mJcZMfEf4L/7e50oT5CgEjGQcF5
P4vPF61CYA4GvX0owy3XBBcD2lG6n8I9SfQrFD5wtkgQ0DFJ1pIfjdGao5nLYEj0
CoM2qy3OuJet13Wg+BVC2kCkTNH21GS2EX/+8hRCz1KzeHIWaV+67rrQFXxNMUv/
gRuZiX9TkXw/NZmCQbsL1lCvQ8AHkMC1r2GgPOBpN1W36pDQpKA7zAe8/BNM3wCb
dc6GNu4dU06Gw/9gJqkXEln461311xBLQWhIzKQbPoKJA0yF7+DY4+vwyD9rRBwT
AYsWlckIX5wH+7XDtZzm/NLm7ay6EPtPKHFFiK+rAgMHMrCj9n8eU/1K6OWipV+k
Uk40I3VZiHVaevJ6cWOsvWJx7JoPZDb4oXE1uA2aam27p7UBVRCYiR/ppOY8TkFy
3nL2f27yKF47zt6VxkmKyKNygQNA31sgbFa4otk5AJJcA63MRIHGoTWlUmZP8vjC
9kaAfjsPyZ9cdSC+ccal3PA3eX3jcDqL3HjP7jbR10y3dPTinVoieanJfK7b45yn
o6VVBDaz5cHMDW97y19u662cKARDRVvXs0RjepzsfMQb9BuycjC/GgzT5eLO7NsC
Fddlfmyg83OJK3BvdLWwIJpVZksk6hm6rxF2ptmFAPJYCRk2nCfhSAEG2Bq7ndN1
dlvB1UoKOJr5EaOaQnMaZK0X/unpycVmlof3wC0EjWRLPpSQRn5zgqndVYlL7MgX
MgTnRG7QOtW9GAUgHOC3KXtXubwmD7rq9uSvBZGdgXYCYtrrxXsWLOGu42wYKr+C
zYV6+jZiBevo0tQzR1JWgzolZjvqFspObbmLlSUoNGcIxRLfb3MNbS6SE9aWibH9
g9WJm/a1Sx+Ny4LiGLx8BXNIdN8L3Qf+40butzHEkf5SU/MBIMF41z06kN/0F2Su
bereKpf2UWOdL9kYmdDLsIGNoZEy590SYY6PYb6soC6NH3HK/uFIfkuyQwgs17Mo
qgXT6WlrMwX6KcF9J9HmB3777gNYjbwJG+Eo3poKAX4P0CwS0yPS2tTmRop/tsTj
YwB/6/XtTN4CvXuZx+JsrGxX9V8/TBulQITvg+MMcDeddeMDipHYGtM7gtgZavu8
OENJARL15MmEq6y4aEuKb5zaIkTYJRgrvViNxctdsrRXwYm5zI8i+9OaYzd7PBe4
yYXRpHAalY6hi4EYpQqeZO8i3KrQaxZjjKVbYkwpbXomIUh8hjA/KvjtfLD1iNqE
13ETcspMQDELclUFuEcrQ9480Rk7HBDu9oViiN9R3gYJGrXZNdnbZ52x0xUj7cMy
ixaY99TpgyPee1NmmLJIKM5BeniuCZIvdzeJC7ij9faf2cpFTJhWAb4RWczGPiD6
GgEdfxA71npNwfJV3xggVioAo1FzhsH+yCpaLL5uoTq38t/ZPKLBl3mIFJx/ndAi
R3wnZjsNxL9WBRPOtk5nGXdxwPsxL54NNx/tVF+KqUwMd3WzONJdPWpdzVHAFMsK
QZqGuQnRVrD7nHPw1JF8oEtLtbxxuq2jsego/DM4fF8aBG4UgvG2n/bkF8aNAuWl
Djgr3aAXraSAqzb7hmSuwoHf4Cd8B7RF2Zr61yFZE6McPEEScEvNHdMEpHu80k2/
UOlFOn3gPTsjPupuVwwrJTLsPTD61Cmzqs8FSMoOk1I2ZX7rAy9lMkNNF8lppQEs
8+Iq8xCkbce0ZY7CrRMN/G6Xs9DcaGmAPMLh+mKblMRTtXggyXyRdMAQ9qMzDwZx
kEOteHhvO36WhqBD184//Yu+gxCwRio5CHfKBBo4zIzHAs6ej4xYeTYtTsVCis4I
zhxP+EIORPDzg/jHusEF8ebF6tG0KDPv0wWDikqYCLCor0PW/CJgI6UQNwTaJOfE
Q31VGNEAVhaxbWz3wpBF+xQ1NgTaF1buO6GUqKNOqXpSAwtqcpcOvntThTxCGLan
DCxGvghLkKfkFwbDFWwgNchOBzWC656cJv/RBiXRL6dZ5jaa5rjHG2AFmwvapODX
Ia03XnBIKt0OT9NNIah5QGskyG5//+ceDrY85jAVG8KxcKsZfJUpL/tsezn/rQpo
1y3q20qnTvpxqIDo7+Xods49sP3nH+6HdT7EBZwm0G2oUfzA5KZUY63ewzOe4w2c
7SIZo3CDg66M/6T0GK+stC09ODdv80IqQUP7B2S7Tz3xy5LTVNHKN+6uOpgQ1Gax
Ub3YyHQt2RN2jAwzIaSc4b0SzR1sraJK4mq7jOatHecqlHhio/q2B2B5PX9FYuEV
lNToEth25QwndfoSjp/ovZwjQDoIYuTVcScV4UD+I4w69bn0wggvOYiKwOIae+eD
tdBnl17hhA4r8DV9arsE57EWjJuZk2ap5lv4UCyswwXNwJBoXhQiYMMx5fuNXLna
pjnf1vBU3Fkq9Dvb42WgZUwyYd85fgZh1VntT+iXLXv/o9cblq1wRjAcPJ3r4wB/
hLUMxmKd9oHcNUrUcmCtivatXocFrg83apH3/IHJmKkTNxyaKoD4astj6EiLPwFc
mBe46SKdAAb8Mgzj+Bce08b3jrDlrEC2j3P37jrwWQsFaddhIU+ix4iE2aL5bHDq
6fux0Ex9S1rl3vT2Ir6vmx4GIDXeFrxa2SXyFAt4zLSNFHaDZ26PjsGgvwjPtiuO
bqy+ApAwbGSatwclvVpKS1bLFf1+oDvXctOvmr8O8kVir8BJ0gAuhrqk2sBD+YF8
7usdRGv4/5i1ijBk6/I+KdtvmHvGM/C3TQPtoMxF1DiXkShuWLvrMNfGOuRRv1hN
y3lZHPRezhJhITNAXC9qPu09FEEn6b7AtQ6tLzDB0e0Va6o+Tuan1pKb49qcroVg
WE9Dd/EKVBdyIjxxeIViDNjnm8A3B7GQPMKRtkrQqWNLH/L/v55cqeqnH/aZyb+h
/dZwxtUkad0kcRFl4y/Vemn5Dgf5O+byuE1w4qCKXaTRWv/pz5AQF1tVr2SeaMRy
azCL/2hMYksX+KHcUp6+J+qYVBlrBTXA9StI0t2yGRnA8qR6RP0+y830guNRHcdt
hPCJFodDvagmM8xn/bHaiO18W0nM5yzh9Fht4XOpOuFTpDW+2rLjjHCGGs4pcs3y
TckO8jnLz/L47FDGOf5/zLJppPXhV8Ae6GpqPXNapAlFuOAGtW9wdVWoUQwL1kMQ
9ahffjkQcFaD2q2mWJV5frUYdGcEGfLrE/EvKyef9e7Jjsb7Zz9k238cFmd0nQEo
WJwuuXqTyrBb59drKlNxdhU7kLo0WaljWU2X01o6I4w3pIwZcpbnevMMuQLaK0ee
ETC5A0EV22j6qpZe0NsOrbdsmiB3q8gp0TVq2eDcu2Frof1XZBcDkc37o/KivZ4E
iDZpI1HAbCPaGaaqtxIYTgN2ydNf3g4ruE5MWEp2bl56RCBNnDaDc6Q2sl3dBKQQ
yqnKS61DpA9ObFL2rATeDC6bX9MC9gEq8DVtSX4b+G3AlcKRxhz/QTlXOFHvaC62
MJADg2IEg8VTaVTFFfuKtp1KovFJHCSB6fU/F4KagIPHOPAwMloszFyewJdjjy0N
/Xx39ltv5uqFooOoralGLOWXBw2zSjlGB3hZc0xvzo9UcqJKbNTiw/+7C87MUY69
Q81x5DvQ3p1KHJiMAt2VIv8GbHExtBH88yZCRb6kep6oLlY9TG1Wu+82i4KVuBGx
ea59SblVPVp7TyJ7L9oaIfzKQiqPi8Ng9g1qT8eD8Q3y1aAJXrO9aNYOKqx3G9+N
J2Byy1TlyTwL8Ny5Q5ffOHjZgqSEjlEA/UDNBPm1+SQF6AROnHnJpDyYL5UffTyB
CnnedzXEvcB22WC2A/KtXdOrms+2LpLS5ip9sRPVwf8WF9J+etoYAqBMZjHKVNHr
NbMOHMyBHH/cyoKVP4zTqVi9owme8jAF4hUTb4l6mxiylJnhTlKekdnDN1gsXaOU
39FArS4PotOB3msIOxHeMuMokBWJ+aRXoqLOI/wE53bzm3cBfYHtrxV4fxUXVOmY
lntHn87RJjVGw3pEZTiPypCt4Nn5R7MWHfsCQnyySeHvlPk7Yuo/fQrUS1gqgyoG
LdkjIwrlUSuqwDxhw5WpUij4h2VBXnYyIbMm5FvsO5k0RIU3sm75FY4diVD79m3w
j+qsAvuq+yqtrWouJvHxiUJSmy9ntRjqVl8D4JbhHxWhjDwfVeIZaisFw570UnyT
aeo0Ih+VXu0YPrQBap3JnuK57S6qwgTorf+t2fx+wu8pq9J1IXg02Hlo7hMJBbvA
e7H6AnP+g7xgOh+KA8uDJkTXJL0C33srVDJhpH7ak4T2NPujmj5s6epQBt/0ZKjn
Hycx+EApFjHHEHp3XrWVXh02fkwKQWosFcbiRVoiBzNjGUEIoHSOLbv6omEkD1Jj
cuzRw3TJcqrbdKGSh2o32j6mfKoQ7WC90dTxjxFBkut7ULEyZqt+NqPDRJBftXFY
EOWBiqYmHfnQJpVg27qbp3aa1+Xq72wTHqXC3+khNer3REGnKkZIbeOnUof15LAj
5mmLJ52cdygAC3M8nnNlg0V9rSyQzyD0cs8d2p9scZcsLDtEFPTaBjRttejmtKOS
JqtS53OWGqW24sMMKWjVe27KA/N1gnQ2l/Ovi5wZtShTvGcIuWT6SOXKS/pZb3HI
CrHHzuO/Z4uOL5W2hV8n61nKfKRE7BPnoP/SbfGLf+UQJ5b+f13uF1xNYFert7qX
YdbIhPRKZT7XBBwWAv17grCNY0hRqUtFSdHc+CfmGUK+gLzWdjFf0JeZ4IHLz+Ok
PxwAx+AFHb1IPMHqSy65uVCuKWzr5kCg/uJurxI2Vm5lj63iouk2YI6zT02YgMa1
U7/QbHA1MxHdu3MekL0qjI55rXTer3uNhdgEQrSkIJ3jEPuEFlAJwkSw/xB/ioMO
yScCUm09afv/CObxRMNzSXoTTOoiySlUBT9is72iN2hEsNIx7Voksm60K0dez1iI
/zV4UsCLPuMq9+X2CsginokXO0k+ppCo9Ii+fI6Q8ud+Bp1i3kw7IgIsYqE4gP6Q
9DnZ4DTrSfn80KTZ2QMoSExNOeyvQQIcD7HRBsfydoP0FYTJfRSATJhzUYXR3C37
66pm6mmOu/QdVVHw3G3KGPfefeiZCjte4NtBc1NSWliGJ7LbpDLf/N4Ig5Pbwid8
n4SWL5H2ZKh4dO7mB5NI5v+vNaEM94udDZE4y9UA0+w/4UP6FIN3WCJsKAtZgWad
pTUs+/jwgi9biMsHRDdxpUYDSZlq1rz8uB07iB5LGSXfOJ0tOb3s5VYKWNc3HI7M
eNuBAl1mfTnHWA5DE0WMlRr2wojuIUyiDvNov9M9UJp5+oCLaRerqUA/NwY1bhQT
C0akYZp4H/62k7BPzsixM0Ah6Oc2py48D/4s+dDXUX5JJSNnLRhOIkKEXNVztnal
BsufwZM5FbxrohIIino/QBv+47zf+/Pv6tHYj2zSrCnivfytKxzPzsAxMhWrrwae
2R/yDMe5wGcvOLfONTLIWTQAM6CWltWV0r0kHJsunzG8SaIgvho0thC+kxbvSGDB
YXCRNtfcxIOin1hCniOYwvz1u61eacHE0mBOZ2u6mknU+T8jj2iaXcKtQkkBMOOg
gKhCrwKqFph0OAHvN80TolmlYJ0tUYbZuxv6VC/7zi3YbUrsJx7A++3O0B9zTHxC
kTZ+T57103l4jxgQ5moKXh1OpKiKFXVz8EwEP24CYeNquytt2PcAEKr8szQ/LX2h
ZXOyEDsW/+JA33j1ax+q9XaEjhxfpzZrzk+jtJdo5QNLIM7O5Iutuqxevo3s8Cvn
LHAMk293AfiFYNpiWk6i6ba5qmC4NzHjch1CAMORjBpYPqn/rVLG9d8D/XI8uosn
2PIk1bKNdfnRbHnG/SpBgbpzrgo260v82vVM6HwP9B8yfrtln75LIppYDasSQ5lg
EhLEWHFncK8GaC55qmVOLJc8I8Mg47omBAaOLX8IMJemZqO7W0SNGmzZl8aTx+Ss
bfypeyPxvx8gchw9dayPrZBBZQZ63nCKMJXYZ1mKtib8gzK6F4WpxfjVFwGLYRCx
Vr8mrFkcwOP1coMIsSa9wEYSG4EWVElJbasTGMyaVPZlkEru8WcHOZwejMVaPcrM
xnr7wlg/vigMSn3aL4R48rmHZC45E0CTpTf43but8VdzBI80/RivwVtW/XFbdRUE
fSPs81a0G7YwPJbrSikiRN0cMAyXr3YLHbSE9UbfEkxgbVUaNTAQdV2GN5nofhb9
feD9TtobEOsB+mOwaijLRlvde/oLoYGP4V2c2rWBatxpbFrK0yfL/P1os/4f6jW3
XmltbyR2O0p++hhSLPVbnT4pFSUQiT95R7YPL3KWbOTfm59bT1J8yAS02YVuBZrs
ulq+GmJgqIaUVUzTadRtq1TSwTYbk5JbpOmnfVcSDygWHisyokFk2T31n/6cQq2z
V+mnM3i1nYtuBOLKXR+44VRkdZ6pnP1XRJXseHmqpI6fBqE0gMA5IISiCkCCbaEz
SjWPWDdX02p0/Ap6I2DniL9Nq0wP78DrkqPlRdawSo5xB2dXZOlu7ppFOV5MYitr
YiGgiMV1T6FSC6DSIVA99jocKF0KZnme4h2XrrAr5qArot2jtUJFgmWYVvpBkkbz
aVNqVglwtfzkU6v+qwIevd74r6TnUdsNoz4CGeyztw3Rdnw6dOYY0z+7VLLcpSnQ
rgOQ/3SYjnCvTvj8nsmPvCFY1DIyogLnOqObUeUl7/wwawNSjEDLg7ykzrrpDkkd
vLNoRSa3QXkjPEC3lxJVfyuYnlxHWWCYcjX3RIN5gH2FmoAkFFWkKLJodxQlBMVP
f8lLHe2MXqHRBqYS1mRdxLwQoq/sT+DGcIFEcKZAyU1Um9X5844E9yscgpRvX8jV
D+vnlU28UvUErnl6SyrMZthgIYGq6lguhvQp/kDRCuJDgpx++6kxYbRf40NjEp5w
sEKbcHnrqeJ/k80RQRwqhDcqWqcU0aOfaWcqHgDtg1VaRvETRFxl+aNcIw52hJ4W
d+FuqKEaB2SkGEmcdM2X+JcdnQGZBxLWp9ouzvVVB5f46wBsYhSLpk03s81HA8AV
V0GB/wajGRGXMV6lsaYf6rDMXvH2qsnjN9tbYl557Q8qrgiqhLcX2wAhHjjHQ2ZD
u0+/87kbjxxWqHRoWNNSsFMS+lWmkd7mR1EZfSK47oaWdhYQp/FpQwoxIRBA/aFR
9xoXGKZQWQGeqVeXUSJDbGeAbeePWgbNbaLi1sbqfM61tp2qafNdEQ/4Ex9P6YOn
gPNThSNCYGnzYB51aH35N2SAZxM/76yNtuRt0QwjkDLA/QFeCMItazWxnROozv6g
eARpUevLhaAyKeRMOKHu3T+vFF8N9HKsJjzBhGzhoj+HWZEyHdz4v6rmR/aKmpie
KPv8V5GAVRSYrB9OjvLCmtx9LNFDywBb3GGbf6x57GanoBEX8swuc4u/ERhDpa6I
ZuJKahstawbEkkohWA4SBEM+UcQVXMDbsjbApSZcnuiz47glHa3coSFi854SQvXW
wd++mAD8Qwcm5qFWWLY/yLOcf650z/wSm2WRWBWeI7rAUlKWdYf1bUhY/8yiEmtb
tqh+uMV3w5Ltgk5ktI6EjOY484mAe7A0EeHR1sQ3imaIUdPIdjkWrBiOiB3si9OZ
PilyJBnCX55uMe7Xxu6RoPLDh4jD8PnA1+9nMr8VFMIcVouwChv9OGE06ag1dPUS
bPohJ3jcsz7g/jXD6NZ73uk4tr/DnpZF28gby57FyYUJlYyYqR7QzWmVYggmAcmA
TUQiLF3aWMwtk0T8y9Dx8wAmv3NKqYOT8vBNf//7tzL4T8zpgBv1JKl+ebFhyRN7
9P5XM6St47ik60gzCSlmLw2qkDfVpPjtD1vuw3xP1AbwfNr5t4YMKNt30BsEEw59
RcQzk92YhFeufV5yWztO3XVNLfG4JwDOULx7dDxA1e4GpDn3VgaAw1X1n4QpXnCE
XxSglKX1N/8/HMwt/WFmppkSkhVpskYEzQcF38NkwvWOFYATQE6fGu/XQMjLSlTi
EyHtZ7z+CPTi8OBHJsO8v+N1HNsrshxm4wbyiYN2DoH2AyXaVnqo4iZ5NzeqQLKu
4G9zwYs1g4FuvrbHxhKkNR7GTV4yFQn2arUPLWQDZT+o6qZGwr9OG+eWZPrjHmEq
bfiztLycpwMbw4eZBzLBxUANR5knTjApnljgLpwCWYy5DNOmCD1SrP/X3nEhummJ
b3Cc71CtrgXEsjo3u1PZw+6144AH/YBVnRhAxEAlkN4AKsZYK+iiFLG5M5FQu0fU
pVg+ZdXBn+tGsTR5LHfWSB+kVZCDIofCweGCdmirLR9Tf3qmf7TdkZzzKGtgZYKU
CGtvbZBXDYp25IPsHJ/BnRUBYTTCIUyRe+DxYRncz30C/f08h+P4OYUQ52+5o23R
ib2PAQJ5qQpVyEhPT3bvEVjj/VQvBu1kej7zR9hmo+TeJoWBhY2IKpxKTIodykgn
WKvHrWDuATOGCdyvyi7g9haTyza50gVpGhXRDkisez+Ng+Jf03HABIw3w3Laxyue
GgaUUTFDUmIukrx7O1/oC2pF38Mp2xwUAc+ajDr91b/luIvZV8Ovm5huKj4SgrOe
u7h6i7uM2rHuUVUIXVBZeZxCBOh9SDD739dqKrUnliEEEDwJN2z7S0d8ylz3fVPV
L/E6a0KP9ttppSnrvoX26C7To2FJG4i+1YP4hrB51y2u/PuBPSNtHCtxCAw1dGkj
2aWQrCO6SEs2zR2/SS+Fna3XR703NsLEsNNfdBXo+que2vqsbJWWzVyeuTUziwql
1HJOiukxjtZCiNQQJm/XjDvox9lEHaKNrBwaTiCO11b6EW61y1V3yV0yoCv2q9Su
qDM0PGwxbWUzgEhzpkPcpGrAs+4da9vudY6SlSsWVye+mJUdVz1tZl/bke8WBmgf
bTzKVHtjp7AOGI/RTMm7m/ptmebZsefL1T071n+1LWpb4Ub/5Xs+cOrED/TjneRP
y/1HCo84j6NSvJYtHDL5yxR9QoI9zfVeiTTSxfzLWRsrjTiKrV16KKmIh/OezHKa
ME4tyDA/+2xnX6oLzUlXiEvfIMZuKXVktxFhJRT7Rfvhs798Sdf1R9h/cYvVym09
SoH2Ut6XPxYzlcWGZomYRCLjRKgCrgYGzYw5TtG0xCXU7pZNqjUeDzh6VJD0RWgQ
Sc16cYSkFmP7QA6e/PRubn+o/iaS+VvxbGgJD3bDtniKTjYGouSAnHfCXhiqakNA
spj9n0iSjco+B8d8XBc1ja/Re4CJ7WaLjOg3vnzWQMZ1RpFcSIWE2HoCXz4jdQcr
CwX3g28lU3rwbj5ZcniAvfhmPCnZajxgRNIrXDzOeGMs5Qfjt+RFOtpzv4WmGpys
33xugkhLpJyUsHbg7sa91RLvOm/eyKgvuFDneBaF0AA5j+7qEOPW/m8zVpYuI8Uc
RlJyQuVI0Eupa8b/adxIH4yC/YtX+KyJbblOmzCP3qin0LFxC4/V8Ufr3Qt469o7
QiZhiI5Kzt6+duhxyLnY4Zi+eEf0G73yPQWZ+S9nHPGEiwV77adVngfi8P7sJ17V
/nf6aUJTzRhJiPRbdCCxRinx9V4H2ry5nDlkkNAyTgfxJ2ilAQkAcWiZ8D863bsB
QrM0KpzH/6AfqCiPbfOFrjn3Ra5T83RxR+pWoZmbuEDPkEhjkfSEcchlqOEQiujJ
EX1obWqxkfGxOFdd6MsQu5ihMD8SAVSymKjQdh66a+UvwxAX7WC7YzN2yCpY4sLf
RFRxIm8IoW9PEWz4esGhVqehp3lSUynzi0db6e9F7ZpWu6hu9zsM05blLLcvHiHn
GfFsnnfOLSi9RCY/JOD46a14GI1GoLiOtyNopEoAmIvR2cyqCgLYoViYpJmnQJCv
A608RhWlhHxprAo/EaBC9R/g1KHVhRn2AuKnAgOXykL54Ybo5mru/osbxecDh5xK
YQ553JVkZvnYZ5caEOoGzBz713xtXb4MH7wytvfJb1i3CdCLZmVCLCwRxcGz+7dY
FepYhkFdW1j3G6U2xNTplrRzRj6ljZLWjJ6lHl2jY58hXHSOID3N+ganuiMGtTZb
0hVqgNbfRSSxJ5HJ9yVDdCaNPbAZ2t2yIVGQIk2Lo/TDdXwUvx4EHgZWKRTPIkve
FbOoqyiJMpWjfKB431cltZAQkxVrf3eNH98dIFXpmOXJC35Fib1bbzUpkV/5zwHS
XDBeGBrHWjRvFGsZrmaAD2nT5qWR2C03bzXqtgUa81+kKSPxqwDbz2J4bmPhWEuq
/mKLzfb318jGjun/M715pDigUrxzLjn8nfBiBum2qodvgRix4Bg6qvEEU2wSGzk0
e4tVAfAbJuuL8m7sgibsl4r/xhGuU/MOGLrgtnyRiC5qe6Hbmno6sG9wiKAOjWdV
yT0t02kzvaTF5Rsw0Q1M/q3pHGK14+GdjNqVdFyZFdUp8kHSaoy/KYdGdSNTQfp7
UnvrFXuBvB2Y6GT4A7apWAKjjxNMyDIxQB08BCs3ztG+5JRpPOhnugqE6rLPUIQe
n22FHXVCaz0fDafTxmfIe0AhbAWwg7XBmuwWesSy5M1KbayBmz5fvQVbVDlBDIta
N8SEOGpRY4EyfT5BklpPfDJfAj/RBs46tXc0x69EG45lYNLAGYKf3DOZ/A4I7Xh3
SEPmbYCp2TKRaPeh9Lt1sq1HwOaXWlK3HZ59W9rFYRfkcP3z0ZtB30IaqjRUe5tz
u9ITdIF07df7sMksIectUrIHQGRnNciSo0QGprmgw3cz5pKyCT+jWJyH6IMNmbPR
LmLo7+Y/nfgQEJvY6oMnQLzDvt1U9mEUJ6te0DGw/xYntWdPJpLsUZSCaltgj3dn
i1qq0yCqeZruPY+EpyzYm8jqf/0izqtbZLXoG2pCTZjaOAJzzhWFkUryHJVw4sg7
iBjrsvcNl8pZIgBmC2Czg5cf93BuFFum14NQyXjgimkFkXB1whImA90B19N9MkoO
5hiAwGXzU436OLpfJxVMG+3qhUf2np1PtNDi6suQBuA3d41CDDHGkJu7LCnGe0qq
XRPSTE8lRtFsgKAKJuT16W4Q3g9mPhI5RuHahaeahc0eBu7nJA9PshQ05x2FT7DF
QSXH29VNTlRWhDssLZ2MLhQq2SVf2olH4l86lg7Aqsg+E2Lu0f4+ArpLBoAzfcbp
huoa3EmcHJeuSgNrPnrIiX51A72ePeI4RuwCL155IsBjIfUPvSibIIh7RfQjAaqn
/w/CgRp+0HD4STWu6Zhtj0y4TAtgj88ua9BTR35lwmgafyOpRamuwshrJ5ijPK+k
+3B2B0Ta98kTKQZHJhM+T0f9SaauZ+61TYooXK5KntQFzhA1aSmS4jP0oG5LynJm
SrdoGNkcfMzwuIZiqAZikgpZ4lqE6zIy1FFfUC3xUuxFrVYrBVKW38hYL69viYPI
WtBQRdbalxsqAQUHjJefEA0Vmh22pNvHtK+f+BDn36dCawmrMmlH1nSGYg2IO8zA
1VKaFYr/+tB8MX7gCgC0/Zj/FMSgBBzMWW2mInl5QOFvGa/cSHW5UUMKvZq7Vwng
W07CE08uimm0LBbry544XbViiyy1/4v59pJyKNtiPQph1Z9NaBiE8yf5STtDZKxQ
O/V30xrX3PzknsxahA9tCHZDAfsvcjLVSeKq3V1a1MCqUwraMhdxKC+L1vHFFFXf
AArm6MEeNhIIqglV93nAydkD3PHRco8DP7r7BVMNvYHMtHBfq2gKia8yoQtkwkbw
mFpGrCcDzMynfPjmE8luu5mYiHxzwz0ie1OGgSCZdneqlN/Q0HILmp+XvKqCyAB6
S69TF0SAAlM4ulLLyFzkUDLmVHxgb0jwZTkOEwgQqgKmYUZq0pnhK344t9TNI0pU
CJCY91izT6D9ixvjqYrsPifuRh3kbHs5as66a3ey5LS3SEmhvR9vSp9Lqi19DzOk
C0sP+mT95ZsDkDZ3aUZ+UdaAryj1oUzasq7qi//aGr8XjM6xWTV3OC6Y1W9WxwMn
2SGNzG8r7aZQSeH8x7oC1TTPDD4YtkIFgOSa4GnXQDgm6XhZV7VjGYRxngbvaUUb
PudcFrwAyhhQnd9IGzVpi275Z2YKL5PGHot+vW3CrBgPWXi1u4sr2skI+1fYG1oO
Lidvg6RiBwRX0mz+BWuP++IBK3ZfeTm8cbUGtnHZCcoUu86lomsYVeqTeCctm024
mByq2wBoNlVsBO0r81HANH/VRe7UJtomJaakka1vFq+GyJtdwezc+D8mNHitjfyo
V9TiAU0Ky/1oHyOO3Q2UB8PVdhkgIXIluoJuVYctj9ZAmOKZJxXQVvI4e1iuicDB
TVJ3lIKa2gO+AKxxJVxyngvr6eXYlLjoXqiVXHG+ja/df1U1jLbGubblmQeTB4q4
044YDSqM71FT6fkWFRtX+xIqhvU6P0rSrm8RjhCnGptCRXmOMcyBpTaiGpfe3srO
P15zUIcfwOhVUbgmCYyhCx+9l/F14lwHILgsT5yjMwCvzPbmdfyImlYzV77bzyk3
PLy8IoouNcabYe5+6SXtNIhiWRmB+U0QKLompRqSaRYIrmeYNdfIM9uqRKiI4ftU
8qS+orVe2X4CiLzYAo5CXnjtk6FEBcNCBvApzX7REomqBUv7dGPgxTzkbmYdTD5P
yVS48Y+kHhMZPETCKq90Sfk8XGokN1IY4pbnXPqYFsKsKN9b9hOh2OlAdYpbFQjP
Z6UMlvctObXCUoalLqvvqX9OqsOVygkGJzYwoXdH+Q23p1HYb7HVCrBzP7rA/+4/
ICgVxmosU6U7a8dOgRSfynAF4/jxCvP/a6vLVApyoOh+gt/iX9PBoEvRKfjlIfW7
UnqS2hUQqFSDPYM7xrpzb6m/XUWluzNMKKPQOtWMmYWs4UkxvKhc6+Wu+zUP1+sL
MvSQSYWo5d+xJiAwKI3e0D4LEY5ggJ9M9no6Ze13+rhvAe4VvhTREeCVpCak8q06
DFMsJeT9jcebBq/B6oHYhxcvleYistA5P3wiDHY0ZrjVLZPggmomBLAGgBHI3uOP
NL1fB87Zm/dkK+gziSApVs+0SLKc0ZkABaJsg8F+aacK+Hq7otfKn6+PdCvuXREF
jYM4xFrFBBo0UBe+GadbDKcse1cfJRXVzQZS4SXBwcsHUG9cM88wUQIv0lfOagP6
rm9PaKwrp2wYOHQA0ri21HPuyihEKkEBSnP6ZDrC3yg9xoXIIpUWs0HzP17vAQ3x
wZ+B29YUsnog9Pm94E+wMQrK1dr77f+GJDESftWOQBZiWMUcqVnJwSgcAuWzUaTk
PomZM1ln4/JYVehyiivflK287LRhPi3QRFZWvzwlkvKRIhGO0566pwR8NzLsU6+W
/ZZXnFUlFIZQeleP8LupjD5VfEGj3X6IkNQNf3Yh8Ackb87WGwL6RHu8POZlzTWU
yNmpqR9bm0+CjvR1dgyarC5HvHIUEwmqALSi32GdvnMCI434Bp2L9+Oz84q2Eipe
K4H7UmolSYV4E2sY0Z3GF2An1Iybgt2pCEaIFaLEUow2HADXp68xHz80lC5/gi1m
9qoTrEENZbQrkGve+6dhisZ9pumrNav0ZpCo92Iyc1KxOLXHjkVRb9E8/rP5cyza
Km62y5DWaO2gtX/bcFvhJGT/n2kwWvCg0WLp4M0POLjkUAu4EE494LNLhuk8HJHY
zREFy5VkTC53S2/bwyiFTVLRvSH/dSQjV4RarhdvZ4SIENZHCoYY6BCiuLTdGkkd
XO6EiepLWZ6COU9lSgkdSKeehCzL95yoCpY966XWidZVS5em7toryHUjcKKnjfRk
yoZDdhWR3ITV9tZUjSpIe41pFSUzxjU5z61ZrJ/avtBleIwlbCqQCkd2F3UMgLJT
JWuhEDej49eh3gvAh4R+Dn2azwmRiaTBVgsXKr43Jl+9iSvQGmPbNONns2iB6cT9
9DCofD6KrU8ps4sl31oYOl0mPFvyZYQe9u0dE/zinP3dZc+GCKaVZiY4EUA1+Hfn
OULgwk+cE6x3kyBt4HUvHvi6/iccH4tn0SQqMqhTWOJSHRLgYz8IC5MGpIdepvD4
c1DqP4VL/MuMafcyBpREOBOwTN1Avma3gZah553YiU5cFFXOakDad6QcJez5U4Dp
lDbTFE9nAFXwMOg6ndcOhCZGs9hfFhwZLF7t2oUJRYckz2a60Sj0YZkIoM4Xsaa/
5lpEjuSLcx2O/JuyZG7PFHDK2/syHPW3xnEYr8bbZ4UrUM59bwL4QBeFouRO3Ned
CGIzy275h2XrIm9x7zbIYy9fAYyGbUT/1E1HAj5QoTOD0SzxEuG4pad8sIoHdq5x
fRhnbpEHUFpw0eKSqr7VuNXng+7gWYfLrtJis40g69F06waPR9Lh+D3HBm1SKEJd
4hGnDshYgJEbsCAvg78x9UM2nrdnoHqknGxfSj25XDyj93adphqpkoXDnfASX0Id
vMPx52NhvexBGltHYrc4OMa05cseB5QRWKWt5apB7W16LPluUqxCHp9voQaSfHRm
v/8Jte6OYmbDhvHC+WV21t74CTxG+5PFd0/ztKoWqFq+NXFew667jLE2ibeB4B9L
JtzEq/2K2L4ceoslLkp+oQYg/FXD98WMgRUubUFT7loFqVYkcZoBtcdzfO2siQFn
W1V5gUruv7ynfggYq31bqGCrL/HXOq4VSL76dYGPo4LkbreAMyEQcDZsdvMOLO1r
kZXSpygwitUQMKQOr43F2b3q1Y87hY91dtZvZCHQ0Kfil87xnHwT0L8mGs4m2W1A
8w0I868yW5PUW/ymh5SoytglOzY31jPW6alYq4GlbhX4AqkatlpOH/oqfaP4cEZk
M2dsjc3OCLwN/7tlWB9Aa1kDnC+uzH8fTbLnVv1cTI2KBQh5Hdp545aiAM/RIuZ7
1zbCxBFR+ufH2zDJoyc9motfIhtmH4/nHFoklMOO6baspYtRFwJk/FkWwod5nnlE
hq4N+Y6eLqhsZWJv1vP4sRkTNUZzumn1hwbtXOmC+1FSzeyk6o5SAy/69EVF1C6Y
GCVIsKa2eh5esSVtt0U8gUhHflSE9SbiS2ltNMSXJKTtxHCjdOrZt2iuAvBb37Rc
wPQ+9pc/WgtfYvnuDXraTZlZXQwMX0cfxUkPU7kbspWDU31AR49+y3DYsjLyi/Pz
gGwa1RY5d8dyead2n2KlVKpIGCuIVuH9pi/joelkd1vg3fC6fwDYcQoN9MrNlzkG
fLbpblCpiCiixQkaOpGlS6La2rFef8lK6wU8OidF1NOLUPXTMc9UinB1M+SNHspG
YVjPNuFz9oMvGALznwWvtvScVoWhzVYq0JlpRoBrpMUc1bVW/6Hbbu9JTQMBXfXo
A/HdCC4Np4K2lqDpRv+ta5lnT9GHAikcgbhaCHWPbXZPVHINpCm35M68k4cIc60B
94gpLEkC8mRVP+bd3VyMpFY/G9tqv474Bk1hzafJzVjE6/kg2oVVh5CNDHUQIHOb
dzSBxzWffnlILjaaQ1QFcnI2jEF4QePRlw4B3U2Ppq67BQG4HOatbNzK+wyFpRgt
vVUKxX6d7V8ghi0AX+aca4Oy1uJmOcz+JFNUHrRRSUBaov3YjtHfr9yznD2nVVG9
4bPUcNoaaPHATZqcDcd60WF2MrJ0FTKMDhyRKp1iUJ5oSfqvj8MSpCyIuAihFsmA
AQd0voohSz9Ki29WOOyKybxqYkcqEnAZ4b+VKWqmavjBu5mynyDG81f0r76DYTYD
PP6Jo3Ltcl0Du3glqcT7r+07UwVIFq8UHRANdgPVsfPIC8Ddly665sx2+PeKR63L
hSHprvxr8FHZwQODb4hiESe3VstbT3EfHMYJurLHZOW1btxA3bdKQX9l9y84Th8O
lbjqun+LX/YNerHuEqHjZx3GwitE8e9Qi2tYBhI0qovZlzEjWTEqX8+THpbgAC5P
/Lyg3cjq2B+7EPt4ciNd7bZRUoX/UmY3UPMQ4pr9dlKi2OAVQsX6EjFH1GdDMcEG
25TTkSlBaiVQ0yyDsSrAe6VLN/bQJ5EgasVMkYmFgWMeefuZdqmxwvCRQdCTaj+N
/JtvlHD1uQH72pN/s+mLXckPgRLTtP8DJdVnvQWk9c4ThMxG644xFYGJAihKxpDR
vIppQYlC/r1wp9zolFCAoaA4zIU62e9rIiREflxMGn5qKXapmY/Fn5zVX2mwCYKR
QwyhoR+ZqqXfj+cSRh2DkqxBet2f6Ile+kfjshXDXZvpARxFA7yoBwS5p1//WWtb
2tLcTAg5Y+eC0vlWkeLvCwS+EkCnnFQjjEtMnS9HikI/X3lp42Oe19fJ1dMByD8k
QqFZ9cGd0MFPZlJd7JdWK3PaMth8jOfbCZVZx0MP83T1md5tcW6ouORl3Z9Tdzyi
yE50MEQlOuPUNBEajo/iHZNVd4u6KTQiOC97SUYH5Pmrh+/hDKRjwh+BxtoiMmZ2
KqNGTY/luF3E7W+XW4EEtiNf7Q0zEGoGboDyj++/Q6k9r6fbuoaRJssOClPobieC
knNuxVSDvHGi2V0LW0xNP994msyfTKGQeobMKRofAoLMON3kogCJ/tCf5zVe/06m
1Vr7wykeFHTmF9oaxXI/G7rO8FpFZwjIbGQNcDjvTHSeOT9rclNqtI/xYn3YSJbT
v2W3lv3Ypcgv9hlGbFYjgnTmtDDUqrMNcbcmMEXqNHvR3LfsoTLSLwR1wJVojzpN
cCXhmWLyLG2zfBh5wbd4vgQtiCJkrANbJSo1qiggvbCr5Oi/zPNqCdhYVYZjOtAq
38c2/6AMfeybVEqL3dHacYudWZsJjZBTssnWEvqOVPs1Tr1tC5gorFxWwHKPY2Om
mZqklWGOmZvNzr1Jh6DIQPJhk/8bx9SG8RuFB+1GmrOJsVMQHXzzAIVk3SP2k/dw
FRNtI+Er/4abQHr1ZEm0hMXCgQSYRItDY4UJ3I0qxFpThQowOKqUHnC10LTT76rd
7WYroPDb+Qhyw4dHFMopN12QnBCKC0h1aW4ld4GefMnXZ7J/pIfR1Fag9LtVsrhj
4gSVpRJBWH3WID/sVxWBUkJGydwXXcsa6dLf3Q2ti0q5ktSSQnsfBxSdNUTf+fAA
j5+u1bSg8/7dFIty8u1KGZ4KCQwaRzSUg7t99m81w76QksaVpZHruHvmnJr+jHCK
SvW9GoajAlKHEQ+02LOzGmBP/uHEcml38Et7mcvs+1eWRHedRzhX618t7ZphHIl4
ChDpGpJlNCbnypYfFzbIDkMmewjtvowf7VvF4gV9X38fs5r7y8tIX0hcmMyW++fg
Jrdhv9BTbNR0pPr/gopx3cMclG6AhPENsEirMWBlMKkX3tLnOD+IE8IrURZ7FZ2n
M8cvrwJLY9/uRBmyBTNPf7IL3jXhtPFBF3HsG5tGu+zpQdYfxCbA+eGQwMcvN+Q7
4xjrDO8LTlToKDZykc8L+Az7TQFnSEPPW3wYgdSX8b1FRifQfDb8bqWomfVqhhhb
babF5kyTJ+Naillxe5Vu5fKCDb9qb8EJ1zHQEHFNF/Cw05KW+v6etocuiBQEqHyr
4db9YDmyCTnBdV4b2aKN/Cl2TiEtpp+KlE4FjuT8mT21sZqk+1ud5dMVceMjn6iW
vry5E72EAX1J5Sr8ptuNIqZHkTFYT2lcFn01tf9vJSN4cukkNBXdy++tvqKtP+nb
8m9NQAN7Y23RA4D3R5M1Bq/CXHBy3B0wWjcisHXWsXqggjhnHULAziJE/4JZxfiH
3l2PXbnacZWAtTrbfWoaKXzwAPz77HvZ75MVadlt2qjmWIx3ro+2B5epREYLrWt+
BzD7Q2eaDXncV56O1eTEIUs4sQLOmw6ih/q96RsmoWrDG4Ni0E3+PhqhvXk58XkS
CRBybae/SQtxUHdzv9lmfjXxF7x93TOuWF6hnr3rR1KgBVOnyQON6VKLDaQyGx7F
69yVxvyqC+dhOMTVa4PG0KSWilkcRKuoBwQt+Ul5kFmsPkaiTqyvh/RxBND08zua
2hstr8jm21KQENEA4k7nwW3RnlqxQs82IcZV/ieR+HZ/WuduIlOQxZi0cpjA7Glz
DDNXex7sFSfhgpnoNu+52r/1AHgoQrLjQdEt4CUdAY0HatK4+gw8iqdDL3IOyNI6
IIDgruNwF9BAoQ+FTsfU9dsbT08Wlpt9h/IgLCylBFwkbmnT8k80+umtvZ9CkzHE
fp+Mx1ukDE/kUzgMq/0Dy+3gfSA5+e0+KMhNo1CoNkjj7pC6UArJUO9ZXljWLvsU
GwO/WKKYjIev4Do18S8J+HpEYa4VOXj5qLRx9cyx2R5BSDyVyUcAhxaEEXsI8LFh
bjqVJ7RrDJf8ccyT2FAj6ats74BbetL1dQtLCbFY1LD6vbsBdDU4QfDUFjaNwfVH
E7exEzv1SNs1q8CpK3q7ytUsb7d2No1nLBrmxKpjx0qK8ftUs5Se9Roq23Lmgvqs
ka8nI1/+98lxs9X5nirvXaVXtsh6mWvNyREAFxppcJBSJcWtWjA7z9Tt2xpU5Rnw
DAAZRJyURXgpeHI5KlSMXBp7cq6XTwxwj1DyNkx6orXco9WcsJxepS+k23QbQFod
FBo0i2QJ6J2Qe23L8oGHFfLTL7TOELhWNFIK0u+uyYDfQf7FRt9FxzTnKW8UApF5
Hpyq2wq22gwucYXWGf07Gj/1B+szYrbg4h0ezxDnBLcEYVBpO3b8YplbzPU0pjRh
vQD21O+U1pi57MNeUMXJIbVwng7LQe56rm43U4FNfYLJnBZoYCXiMwwHxYb8mBrw
gSRxZHJBih4ghqAG/xEFRXq0Fk3W3nHAYMO7Anyvc2I7zrqL8PoY7QU5I/C9B6Oq
iGx5wzW8F+mpV+rbKyoFmJxKoVShY5dhsYBnP8ub6Wrgw0+922DMmF16djc3F+6h
6Tsw0gUAQHNnI6lbxqj+5vHiCMutbkaSQYxkvB9u4eX03z5yFXuk59S6ND+74lbs
LmsZPkAfueoyUlQWo2PtJF9HIsxizPujQTfb2brZ4EJaBHgxxr6p2g2zyr+wPb4U
YZx20+1ch7URXtJlgwRhLCy8JUkkFbQZlnprDRViKV0udVCry4MBIkVGEIgAHUAx
OIEfeGHkCtNfrRURNQJ6OA==
`protect end_protected