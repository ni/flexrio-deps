`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4320 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
HdytKcppDjja7VfYQkCqvIzuw/F43TsH0KyaRPhxo4FHAfTetsrFquKKJ6zaxA3S
Hs4b2YBVjuCbUrYdPjTzCTGUBCp0x0JdQ8J24fXSDhNxTE7m/fJJeuWIxBxJQUPO
PMoYV0zU0DICo7tnFCWkizQb2obji8r2LgFPsIr/MrDBWzljL7r7c4ao12jybW7U
UFj8byG3ZGO1WJGpcew2LBu0Et3b5DEuj8Oj4yqO4rSJULjYOaDoowP46iu0MPn7
S9eKVekSemRTpQriF6PjTvcgFf72yro3uTQbFamqSTssAoIDU3t3e948FppRIIFr
CRgOD94/yUkkEcyaXYp65WJUEGqIw6dHVQmK0NUngpR4H3X24p8Ajca+SI4Cgp0x
yRVqFCrV6QQ6ita8IUnMmUMYxBI+xrnQKB0I98olxoDxPgN+5ZrAmef7VIB2CwVB
vg6rssuiowYQzIEXQJiNgDuV8z26OXziL4s4eja2/FrsdG8oDj2V8F0YItj5Yea/
E9te4HYl5sxHjFUc53Xl3uegQVRsYktAx8O0dYpT5rl8fiubeNDUSUsje2WPqPiM
SCQ/Ig9V9BGWHq2T0/pAnScawrafoXDS34TWhT9rLbn3CSCVAvY1b9zQPMg8RTHA
B+S8ZTw+vi5Vft9tAqGKkEvPtSAuOGyoNFNjuOjmwwXxSQAmvbKnrProroTYhBsu
XcuTjmtqT7M2UwOOfXMLLEMJ2inApI31JzCxcZqaKds8LHmBC3f6Fmd4MYHtxnV/
xCduB6EbiHj/hoOh8xgWIG95UsirOiigUV+WZf31zHd1tDZHKbuJwwL4dSgPRb4C
OdhR5lPveAGeQWA1u15i3ECs5hSx72EtVaaOBeiMJ/zIM3J8VbKKxQDArfypbDUA
8kReRmT5LONzDQ7fZ5m2ejZjF9DCmPr40gsy+2qYi4iYuaO4Okk31eQXq/5yrPWA
qFuoW4mtntkdXe98cJTfQp/5E18194LikEz2T9zTfqJ5Y0iuBzCConGV7Iw/iiFU
7PJgHzz4yopcbCLOVDv9PM7tD711CI3MsYI7wGg2VnMlWc6wprv9Q9FL8Phz17H1
7s+Akyg3se0NDPWbapgM1ofYYsDnSNxMpPPDzD2P4/wavExfOVZPDh2USvzGZ5k3
8AS7naYFKyFR+ANvFh91i0MuGLZKlXxWDlVVK6p7cKqIVwKaCNRpd72B5rPHEIyC
NOenlMTAa9pADtVT9ozJ8uuFjXmXSBqkN4kICyeguU3qNq/duQzSs7zzIE/bJx8g
Sk/UwhAdeM8S7Ek12H2q2oBbfDsa50Cr3TcR+pd/1G7glC/se3gpDULN7egiYpxM
qyQJFr527r9EFiUdq/PYyjhxDJ5i8cWzPuDl6kFA7jASt6LCF5FrzLn31qcVZdoN
WEUzc1rP1ajfQ3vf2FyWkutt61+F1xjnt/f/3O20SaCRUV23Uht2ZDN3vsEu03+B
gdrJresnEV4dgKsR+i8bcl031dzDoqkDRkiJgtCxgAJbyUclMPCkwej5S7NB9HMx
Fi8Jyj8dA4PV3BIoWYSXRvwN0adtdLG4s9fy3y/RTz6gUKCWgDhlySVVwGcWUCew
2DcCSKQlGSkSJJYmjwzTTHp5I9jCGDiIkVOkWT10gHT7W1jbhtgMOIQ8qsbRyoGV
UxTphWS3qq7jsyi/sTEIf8olUB/UYdUMUFTJS1XSS5nlSBJCP6gTdduG9tyQjrij
0o7p2Iq8hfM+MlzwwggxOit8RA5VNJFPJi5jDrPtFCddg1O4gTVGm8quyuZfBwP2
I77Jg0Q/xVuUuFAqUbu/fS0u5KcMJ42l+HEt+kHbpwIJH+dR4MbksNBZA6pdobPs
9RDCe65EocKtyJt3dvK80SkphOd+SwZnqNNW2Pg6UBySKPUfXwQf+rvndz9vySRr
54D4+rktgRnhwaylNPRIMGCPrJGyqyF+83NZnLpAqvW9JVVka1ZOa6uTuUhzxlXL
tx/08Jd0D17m0NRHllsGgsJsFqkleRlNpE/mCBr3xUYV7J+7soiGrVx+klwrtYKP
XwGIMotZE4Mekmq/Y+0/s++0LAbAiXoSt9WCsKkgkXmnkcX7asEw/WnsVDV76PsN
9g4CvDf2XC4d+RPskxd8Ksj46vEavCgmff7HxAna2izskSJjgEt4AZbIHDb6Ey+e
Wvjh7gkbC6m86kHxjytPRgYOV6o1AbiGhhrdPFz3kM0I6sNjhySkbpep2i0yQM+W
AgoIKgXoepYEaAiJg4a1I3zHcEv3HpOdwTa6MtrzGc6QWdqUDd8fChYn3cINW7fs
PyX0xHa7tlAnqBlITcs8CCq1ogI8hFmlFsusAUGQ/Zd+c7jFY27KbnGJcxbYjDVK
8/RI8C9YghgernDsuXQ9ad/zaAW0tunJpCTrC5Wop+GM75QQUdzZqNPju7R05ygf
Z/71cNuHeeCoZv39lDiiy+Ku7gDTpbcyzFvyy31IkMMIz2OiZc9WN6uCwqew5t+y
4eyuXmRjvztcq64BwYLpt75CeaD/d2CVPulbezKBfbIc80q02dUVKjLbWovHOa0m
+SG3lmrPfKnjfnD80KSrjJegFKFQCPjwYTxAvm+ItPZC9RCIYUWDGIixhc6cMAa1
medPlPLTVAuZpihakHNCu3fKraNSwcO1lPQIb25domaFxha+Qn3EMbGZO6Q2kdYZ
xuuTVxhUGY93BZOCArPAr3XMVTO6CQ/pd+yK4Fry0WPfgSfD52ncp28nEPTJqMKR
oyv8h7GsUubm/OfhOKlfiTvvAi/p0jht1AJtZhz2HFPci7CnVjihrOzZb/C5JOEM
aHOzs60z6hDacsx70KI5hkpkAqsX09AJ1UDDc0S5JjWcNh414qtkCtQvrO8F32w3
gFs+mtzuMe7wGq7SV10723qK0U/z3alNz5VP9yXEQ9dzjX4uwVAxZbLelnzVPA35
pvRGeruBEkFKjaaEGWlFko1MirgXhFBQR/lfU+228s2WV0363Ifm9DUzy5wV9W9E
LSDn8TY3shf/Y6q3j2xuJkmSKGeOGH7IQ73DpQWdPoskmVWOXgG965HL+eUXsJ/a
8XccDz7hS1G3RiSz24WTdIeA1PDvfcKVLXxuyaEn7ectEzMwed0pmxSiRQl6VXLF
RiwSENniQM0IhMXxuabsNquShGVJtdHZcsh8cha6bp5EQtdSG5PBy6yUbQVc9NdO
fANoBGO7iBEhKqpymcnJubCseUOrJVPuB3og+W5zSpzBvWRIEPtHfi4UI8yWdW3l
+svbQSVneDvqKPjVBOY5NLllcToNGJOTL7iOBGgipzBYr56PDTxhsdCOSCBAJA39
gG9jHVwePfhOZWp/aJ3Aua9cs21eh8iD8cjSA2B/paPy81Ijn+SGNDlVcG6PaHtO
B4o1sP4nMGOlZDF8A6v1By0aDj/BvvAlbO9FzGsUTzRp8F1oMg3eHKQF7lGcakXM
GrxFsSNOVDRdAmaiJtyC2iBn+OcTL+hTzMjmvgjX+DTODsrK4w1gZHrQHv+v2oE0
lbD+huKsMPzZ0iXrcOdmSb/oYHooecx9NYJDr2MWDBHRykLwmlnmpRNRO7YCbXOO
DG6lONJ8nM71NHpafmfH405k6LlsddqhCVRGdYbqj45qjqhDgMrL0Ccj0KN2pYAm
udWuancnwz2g0AiOcg663bI/uQDoLu48mRPG7/a2WHDoSxxx+mWW5Va+sAC3i9Nc
vaPeruZd7CMwc72HD0j4IZ6OSzumHE6GFMUtaJPnmFHwBOdP6EGyDdHEd8+xXSIS
EU6/DeSy7Jws3Uc3N0mh0Fh/Inq3ja3x5pUqV56/6SW7FID9ildYVcTAUG8y4WEC
FYY2iWd4U15BUp6YdaCkIbpYH8yVj1skBYWlP/4OW+GeNqAD0FULApQn1lm+p9dj
keZB2x3wvb7x59yaZdWr/1xy3+L0XWYITfyjeMcPnB8Dko9aKYFroJHUjTMPJ0Tq
U9zhkkeEESbPMBuwdH4T6Osvc9iXO5sjamBHb31fxnUfgTa44nK1PAXBTV2R76VV
VoNSq2Hw4qwHykHQJHbrLR+49nt1a+JXyT0sgL7NfO5rMLTJotXtqQ/9SL3Lvx6g
1Q7pnxOUWpI4J/w/b5UDoT+uKTxtjJSHqn/l9Px+iaMCmo0PsIwGHb6VElmeD7Tz
QdH7N72F1gDVYyow55lHmCeuXupUNzlt0PwCwBptrV5XJOTvJb44ASuXUmh0KiXw
DWePql6oS6oae4ruFSIF1Bm4F+e/q/LufV99IyBy9Qwft0QBg/9X3wV3Qwm/TlVa
mp035yalhembTquXneKxMN6N9/LfT1iy2P694zBL4ovAvFOq3cNuTbyZQjLjkgP4
YhCb0xbi2LPkG/cXPmQ2ZJYPpg24XdWf3H8HPrs7hkMOj5SLXzWLpyeq/g/bgXMF
frZ5Y300QzzCURhuUO6DEZDrUrzP3XmgvZPww6x4BgkJN4tDyzHvggXX1pVHysSz
7WYZKq8S/hQgbIjPNZVLRu6rYLtiGWIGI7IsRlSgRWagcJnVINxolYYEnkCMAxo7
TNV8FM0arTUCs5jt4v65JnsG6lQf1pZpgptIAaD3o3bxqES/6SMpJnJY7v6KvPPX
JKCNM+gxZFiUfFgaU1Oq3zpfdhglheZGMt8HnI2oPuaHPP9mL/TWrPvgNUjSw6xY
hiZboRP8r3Qx/vXjS3OBimcpDC7X8FYpIbOY9MsAQ22SKyeLjo4A9NGjhcY9QQzq
85GbeFFH5KsVFPdFShj21vzMRVsFAntLeXAcnjbJzm20yPl5TNuVHGVz/Lb7h+RA
FzZdmejchiHgGzLqSSyVsmcLu2eJTcD1DCW+uYoyXQu1C3b14LIVrZHEwUrXsl0C
SpgvLFN+KBGfXC1q93nRnoHgY3l/UcXa5bGSMNTNyub7ES/nMHKdlAdq/SJV1u7m
+onbRCuNgMd8Fy/Oy36CSOUmULYohRXuZsH2GQ9u67BJYWJHGC69q0R4dq4Jqes9
CAoGZ/mXMnBcwkLxN4QR9R5Rh2qgZuPo2Hn6gHm1CsPsZmlNZkYEJnKkSynPrcLm
Fl8K6Wb9Wv9UYVkSzADm08gRHfq0oVNEZaybBpqSDo09bcmkF8aPHXKc4t7wBoYT
TK9ixM+AA5u2CFOD4EED3+hqB2VgjF1RDC80NTjTjNIeQwd9uybc4vDCBtxEaZwC
vetoi5hcKkUX6IkqtRDrndXZxOijTDeQAtliLBac1jkRRRx0DWFt28esfcMRHQC0
vmKX7WTrbNSuV9SuHMPJMMh7lZ4WJ8SyCUEBkXeZy8GQGeLkRbzaBfcHDi3ABxJ/
RISQ4s0fY/E1jcE+3ev52cC7mOX1/oYGGKcP9vPZjDjLfCTBMmeNrhOzwMhGzgkh
6OCF+oNVeGVD9e69lbzoIAMpbQ10P4xKfNiHHnE8mdW24QKyBhaGQufjyI1s3eLN
VvNQYSZJXywLqH4zuBGhkYuXR33EVYwvLRoRdBNc0A8TiKG30dtjhfaZeXntArp9
Jnf9mO35/+yDMJyJCcGE2+6YI0Do1x5OvdOTMvufVmkDG82PEOQpggq5jbEWM+WY
bbSKmLgT832bIfvHBZ1yS3NurL5RkDSXU3QHkSY8sLC74N/7ApUUsZc7JbYi9G7t
`protect end_protected