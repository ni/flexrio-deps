`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 41760 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
hRRAlfE1xLfeNfywbrz10E5gf+DtPdX/cIEuM3y9EDi9dUPEooHWzzUtJmdqzF0I
5DlDNyLFj7C/RqNlffS2vz7zzInX+NyWHIjMAP+tnP9pqo38CvRt/zfS1iOJZ6vs
qItyUbuWVevOmSnLfp2jsFGOck23IysIrBUQXgJZVJALKEDaHCQqZRBDwDx18yxX
qNTBXGARUbCJ071HYOiokAZRPCH2780KOCKZTxjc4QFSIcqEmoLSnnrjWJxCBKVT
M17r94wMhMK0mhvzzByH/YtcEC76/GW9PTDXfja8EN9XjDx2MQzZwp9xqLaVCRPQ
t1gCe0JkLk5V0eZQ3z7s5NtBQs8DnRdCSeXrQNy/koF/u4X5dDL0gcy8weApZa2O
5+Njmu8NhCjzKmoDfrcolO72OIwwuFG/d+bH66kByRyFMH8lixy+ILm2kgObjrUv
ouCgr8uRwFPO/jggNNdppH8BUupHk34I0w6qLWde9gV7GRY81Pl2KMYgT61w/wor
9kUxXqQi0qfgZxRIqaR9sQILEoq8HYl1NWRPDGyUn9Qsxbmj2fUMw3b9YHwmJME/
bTFE9/E5WBhhTgu1IEJBIlDVsDdT1QiFDAhOWva5fOiFkQNuPzkUh7fBphaRc6CF
wqf5wM/5Vl8r8gFKvgt8azI8tVivls58UtnFjoJG9M2DC3FxH3pqtuG3xFyOe9yY
tOLyngRhcrlnkpOI/vbbVLrH1XaEqCqbJIu9gaXa7+efjr9DiUsbcZ6xntqb8U5k
7+na7SRz7YW3ELrIlyGwI0CONSVLIe1hqv3buW6OZRn8Cbwy2Vb682vGquNYgEOb
1V8cOpUoSLQu6av89ZLyfs936dvf4VSrK9N2Orfwfcy+VJpKwWMhx3WteKYnFI2I
JEbOtTvh7rv8qUQME+xOxBQReuKGozgr1Cs+a82gDeRwFBVknbsxbNla+DW1YoYQ
GucCBBnQERepSFYfDuzojwkCoNxzD/38YSnB8M9bboHRggOiH/scSAxrtvo2J1wx
ooW18hkz5Kc93FH3WNcq+kBFbRc8SGQ4FZ4Iv6visQ+iyawYEQReH/6FcHMzIoBr
N3QHbR/qwOELa/EOw5glxv7HYYA2fOwLpNmtEe3xZ8Af0pQ7FmrdfLUHa2INhWyB
UFegqE8pEDxMJooMlTnFifJKGWyPddqtftVsLb9ohggJ50t7TJqN923wUFhUw27c
SEAGiJ4HPdme8Xo1EQVPiqj+o27YyDsn1yw/46Qk4G0ZXln5qNZceBfIAlm34A65
BmuE5IFFzvS3NccDTDKhI8zbEjODuktpUNOBRvfqK/G573+wyx7GWFRWucGCg9LU
OCJMOQ7u8WGNV9TTU6LpWJ19wHKayMBmpcYG7IvgotC8we2F7LIeo9XgibveL5BE
869zrhD985HA9lYEg8zoUqICS3sPxKKh4ZLKBRMciE5oKiCuRHGRVAVowacQSRs5
YA4BiaWk0zCJ4MJJlpihnU8YaVLdPEI8Ny4qsvI43h25/jXe87NH7/q6VEZoKr3T
s19i7AXM1EHrW1GkYMcBhQVlJpAc7vVnGMdwMtrMsKwZw16wwQ7RBWt/dAmpFFYC
kvIzmiazarVNlNPQAvSembu0PV0YjSG0i/xaOJIwOENk3QdBIVCrdIJ9RrjWG3TD
5CLY6Tu4MSPlyV6olUQ+c4su3UAgr9+gscxOHTqBUimrN7G2IQZXFo/LBYHK73oV
2iHGaKWR8pjfE1dFcUkr73jv1VmXAd31/G9z/IzcLkG17STSslTXQdJ27++PpYCT
LEObw2pfoVe57/p52VD1Nq/PHQfpUr3steAOuSrLBLq4bxtfJXE5bNuv8J/A4ZQs
BiOf6fxF4BZHhWfBYik56s06VwwskabE3rEuHA4CuERKVircjC64rq+GUvKa9VSd
10T0lX0WlfOx0lOdXtEk5g2GjU6qGpJvkCKZdH5BSuJY9VhoL9SwfhUdjdraIw40
5mDC4XEuPIF+UOwHpzanTNX3Mwj65YZqjjIpDciT5h0MMBRYKhT8JadiV+GKyvNX
eNNLh0h3bYBENssyN0xxQ8TK03G/BRd/uYTtoozunUmJhgRvWC8p6AaFrDLHJiuM
6bCMsIeuRiNu6jc3bSgwBr7jTJUCfiRWAyPT6tqiUcqSW23hV0HnzH/3nqlPhDff
rGXp/iNvtU2OdfiV6SvpyuodhrF3rx079baG0QRZBmzENpX1Q1nv0QQmypNs3xMp
UtwfGZefiVrfyYHx2Qe5U1F/co0RjjvFYIV/Ku75+g/+d8EJx3FKKWAVQ3u7FkOH
K+3IgpWv9IPsSQy2EUkgEuN7i/tTUoXR/+cFqDL8uhkJFNU+Z2yOLC3IbSbXBNS3
tdvFTSDtCHhHaHMER87PXvA2Y3bhR5KMjRfWBQk8pgS/5m4edYwERjHga3C6Vxuo
9PR9CAU09wcxdRDKIEusPdfM/lmIU0SybmGGJ8wFbzJT3CpDuGEsYthINCZpvyxS
1zzzqzkiA27rmkHYeopVcF41fqmtTU9ejVKD/WOkKbvXBYMnJZkk7ofKYD4It3uw
6NbHsR4OLWV24VrpoYI6q7FKE1lJvVGitSael6A3B8r6H+JjK2oefLqvgxUSVlEl
6ouSKGGUAGH9hUJ3f3GWIKa8mRC7iOmL662vwJIJ9QLM9MYg7poe4zE/CWDTIpMg
01QdhtfNCWJk2IPCdPqs/qmVKU6xdQFF6Kpzesh5B8SLkdlWjLXK+pO9ETl4Vtj5
rrGidrTCFKz1aK14tGbL4QHX65Ru9eAdC8rei//w3KiHVSiQU7igN/uPNKYzGOz4
eltrEJrejGKhXYdxb6c/udOsRrF1dVnK0MdsJ2KWrXSZSmTNABuqHZQeNWfA1cah
g+ctzmmef6T0luZR0l3MgMSzHD7SVRCT3xf9PfVCP7ak6fBN9iGVmhbvjFVoZ+X3
c+BqUa4jMnkvk0jXzI0lEvlPuKBsT0EKVIEzu4jlmDycTjo+I/0buNpLSEmxqLEy
89Q4t6qKVVMg4emhlvikF8/WUT5YTH3NLiCnDcGfcmcpkKM+wIqf6E0JMt6PSte2
Aaf1IQopf3cZA0jl6egD8DsBACoMwLfqP92fZgybOjMGqv1ujD2cMVjwi2O/giOA
kWRM2b9NTahpdXKXk2+SxBQ8GIMacj7dmMN0beK6AlXxvuINPNnSUZgauxaDtSrl
T0Vpr/69mmKGfX0Tbn3hOozGSZ7aqcjEEyYMRBt/IT+JkPmRs169m6vWf1gQlNhT
J60xyEMqas8F5c3P/G0MIsWUEJbCH+1tpGir99Y0GVbNCcpdT194s+2vLkrOsFGK
ja9GOdvJU3IFc5N1dSup7ZiJmU4cvMAw76SD7wGE+CjZCV0tbDseSDTjpTYBmwhK
yLgAYMly7enMrj99SRJtKWwyaHYIrWkyEtn2W1EqsAE56vIEhoxFcdf8ZwN9giS4
6DCqDBCvfBKeivCWHoAf8lQ6EvpaP3FrMHUpxtFjVWSQ9QW7snzGAt+ztky0H+gA
QwaElSIZGebYH59Sdkr4ZjWkgdgmzCNuHP9Ao00IacdDM2dEpgMl0sgyxE95P3m5
3dau/3aUqAXuI5/eDXjYL1fldBQzmVKyPwdpPWuEyve5UlQUBT/AtJHpY3gp+KSC
aLqCs3Niu89JANP7M3x2+oEr52RQWwNOIj8K5tLSiAADW1cl5rdHlftqRjyZG4TY
ycg5sHfx3AJkWqNgkj1mbGRjaThauvypydWLgXNIrdSF2sNKg7k5Y8UArlMdAYAA
RRU0eGFM0cfr9ISRi/suUIKJqCbZ2eBm/hhtycmTAm/z9YB4jGykxxiNZHreZP/q
oRhbB1zooKN1DQDwIHE6oigGzyaBUgMDiXc7ayynAJho17sFdnGbpGB5+jjf5kwH
5/WB7BqH/8OUniAQyNiRbcZhZ5+vQT8ff1ZBcA2gqPUcuXwv3HeEbDNwo4dSBYjH
kK9yERNBlJn7RyXR8nKhni3bqYeB85Bfd7U6sgMBqKokodj+GxD3hvWIE2XJNMNW
QwaoLfJ+zdR2hOp4wfEvdG98Bj3pkhxYSUdVZM/MUHFY42WBkqN7C5QjJiBG+wpn
fioocgNvcFwHpLonmfx3csowFdogRHqIJM+E1HUHJBlZ3HLEhUPsT48MyUkGTxws
frF/U9NaloCUix2H1Y4tYUbm0oXYAqv1klNlLqOaDNznFyivzQaEcP9ABUNNDcS6
m91k6KmvsN4wozFOVLFUuoTYK491cKIHESQHZBCIjWC399mqgBEf3txuITaH+8mA
3YA9b7nRAzrE83zEw/JGaFoUGdkfnRe4FVlRR2dcjTm0eZq0fJfhNRu4otI67k6l
2YtHzXqpZq1iMdpgmfLWgr3YewR1xEeLPB2VeLVzJIitZm1qIWSd60CkBJ5XEGfO
99MSttzGXdO9X73cjSlUn2WM+aBWvgeD+tYLVNTs/ryTEmuU8lLizm6+aJlknAgs
HL9kqjMGSx215Sc0uKghPP5S6sor8AmXxH/CGQhTsKbJLFXoLDTaPaRoeJ7fQPkO
Bg43MRWKkWKl/0GqKR2qrM5PA2KPQkYJGKyoTyXr8S9HATgXrI6jyUnaw7uZRB3b
c6asdngjNlY/JJiZ1n54bpyZyrtjPuQMKLJNAlHYOj4uubMophIrDPBKM5Vmvja5
xzsjPtwVyKouVgxncLA0C/f7XPm6QO47GqfKOVTPKFdsVNeaw3HpWaV9RXMLeVdJ
htIE5Ix2YTOnAthPL995xkMyDWnY081PfNmvdQYwGtuhWB6GzfHfh28UWgdEICak
DAqetg++Qj4lgDZPjcPXP7IY4IQ9cB2knY7kCTH6y46LCsh5fdkGOTp0gYwZYOY2
rfZoTFa9UvyBc38IQ3HD5+dqYL47QSvWixr3Kou5wdMYaehrqCQ6rrcjdmzm9xYA
SNEBLF57yL2oAOMx/HMkboE4lh5gX0S7gdXYfu9PQuWvR6WNHM6m7QZ//KFHgLNW
PykpoVc5Guod9CNGNZaQz+3ncHO8IVcURuJe4kxsEHspmNO6PaBdWESYJpCJ03yp
6tXXXfg9NDK/uGNGpL2ypE9xAZJ9jTz0xPIO8T0BW6gmUyAHJv2MGItEfvNwjIMY
TvYjiQsEej1BnA4TAtlFsXNM/DOptn9O36bYIWT5VhpAQuUqeg4GQC9pynBAQLoA
UX+jGhav3wcEZoVn4ScnWqkTsLo2fKANG6JPGJMYFMcshoC8c4V53ioYxet8UDJB
f4uuwH/nrpKVZFWCy5eMUL3IG8EffvEZnbLdiSa7z29Dxw+OLKUFx5kN6ow8Dyj8
cY5ryleY0hDD0iZmvqWt2btC7ge/HFYzc+9PRLw3VpDWvLMWaV/L6JoTM0hhsvt6
QPsv7+8s62VTithuHdJWk+kUlJ78yBdMuPdjEFAHFmR+N/KkLPSavyAikgXu8LK2
knDAFMh9lX+LZV7tVLBBozfP6A9gXlIOAptmxT2KhdF/aUPV3PeTpwO+BOWBXawm
lAkhZDq1rK6XWWmXTG1Cs6tHkfNuUEjObDmGEF0tLcWP9lq/zON0R9TSnQ2YG3YH
O/aT8YXuJy9UdmDOJ2JPJuNDJ1tlUJa18HUS4TVS5iaTKStOLM/pwYAZM/10spp0
zbRVelAzmXTfLY9AS+wd95T8Y0AbihbDTx62684B28qQjYtgLyDuwDQtNZ/JS1qn
nGbySVpglPRE7I3hCI/bxF8akj/VL2zHMT4378Rst4W/6p62PkKEETfgAo5b1bls
5eEF4z8LLvZPiRmzS+OGRnwf91vaRcY9rPb+32FBF5t9qANt1jrN5yDEzT5JT2jF
ETJd3nBGdb/FyJFck+d2uWhwGNvKtHGF7wVLFBOhwys39MrH+568Bl+2cBplBfOY
dQn5kpllsWiz1dlcpyLQBqBRzsn0uffvDGaxmKMmDWJphTQTKZxqsH0NhLRwsxhQ
fIRCgKPykNmIlmI6rJZL5/4tAl6tPHIS6E8lZANEopQpV3eZMJir6dfadzEz5CC2
eu3f+tlB0/cvqGy0g+726S1pB8pmOb3fJpiXJ7wzlQgqxnbNfmqIpKxFCCS2Js8r
Nn+qGL4LOoqwEViL91xzOQOKbMTrwZawPCFdytTbnO9rTgAD+nBYUqrPtJF22TlD
4VHECDYlkXpcADUspL7XQP15LU6EASAS71ZSFf1u0FORZANbHYjsDG8ydbQe/v/O
B4jT0HgsgacEkrIfvvVDMAKEJOvhQI8X6EQdt4Jn9Dw5/KGUu2BZVCjmnGhaX3PO
IJuhyLV/JStGb5IDwf20k4aM6BtemSZhRq3ehwrY96TwRTMbuSbpJlJ+EnHN9WQV
J2N3htb5V82iwDE6xL3KT2jOEUp2T9KrjXKwo6lGnIXCa+gf+zuole8ZY+h4V398
uwzrDz1tu7ZsRJfLLRx6DfTYhn6Pr3VvgSThgkDNsTI9G+znQ+3qYsIl788zKos+
FJN+LKu6XnEPbrHOHLyACdI6clzBajM0CdYgt7Poal+da65Zpm5kE23yMlkb9mAI
sbDql2vlCie4dgu5IwAAGaLvUkTmhU9RR7M39c3PgCh6lPzUESb2IEEfAO5uqjiC
ptcDJozTlPHOS7WVBZlEkIDE+4e4cl9x87DmS+0kt10HroodaIryAjxTsTSj82Db
WleXYfUz3ivBYnWsI6mHzMqGrMKAbBvmXDFbbMlg26KKOcroiMxPj0tlvx+8yi8u
R8pvczy5ZBckTfY/FKr4Hn4RPXDwZtlRf4Oql1Iyhpnw7tH7W/HYYbj4bmhT5VJr
tTcUug7ZycWIYwI0pYbWWazoSRigxt+8NNgBqEf0Y1NZpSuq41KHLXPQVNJqnkEN
Kyb5i3PMFns2Q6FqAQmVh/UWTb7/7gUMImTHoZILoA8a8cVPiajcNXbrNK4h9XqV
K8mjvboPergAQLTnPuVVsSvoKk0hjIUeiAlPTuitbidT3ggjKw+cZnTa0S6ERe9t
1Id/2o7hLPRdT/ojbjrq3oRpUOHezLGGnuvdPxWlqGlYLkxXutOSy9901b7UjbY0
TVw6uFnhhCbp30JJYhiFsGY6aWe4/pEN6K6IR6eqkmrFcDWsVGCHvjo9BWljtm0O
GVeY/0EU2lSCIUJ+etq1pFx29WLN4nMdbJp5pOY/mg0gRz5JFZ4+fCvQpWq//+VU
w4Ju071mgin6Siyv+hZBNWq2ZllX+ET8B7X7OIY7X2+K4BBg1oiLLCbISE7AA95P
FIPk/mRej57YrGJar2E0xSUA7xy7ZUenSDiWAsWeTxnfApmBLYLbtdSuPczhG4Ie
VjYuxzr2T/Oz7Iv1AgOB7sMl8Kwk233y+djh/V3AVaisvhZas8ONJ68SEvNhFfKI
zUbZhrFH6qMZOq6EWa6tkYVF7NHVifaihafQIh+Ggmp0iQpOluIhokkPlvll4tZM
HkreMJ0j8NbUmwSk1CDPM5+IJszVaEsfO/1K3Ee9klHHmI1ZCwFdttDwMy89pryW
pWVemW034Dd4xLd7EDilMpbQkUQbfi23HITNm2oUqdcv/mR7Ynx8TGTeG0KiEgbV
rIVwn0jsycz+hCP7bCKQZPJ2Sv9ANbijlFQwpBxMidWtOQ7trdCTiynJCbhYqdx0
dt0Kr/2TWGDgYec+yA5oKIYbowpeK/1uIy28RQCjk8S8nCGsubQDvxvXTxYWIVZw
zmUprVv+4UbK0bBxSLiFA7GpLWAZt06DRJKRKJXeZlZfUXiMM7kMQ9WPdA3nMVda
uNE1E0bk+pnQ/rkz7M7NCvCJ0fmg00HEAb7mslH9AMBpdHDIRJR8lU3UdfnmeKEI
Sx42Dy4pVInHkFYzFvdAp63FyYHqrpMqQmT8aJjpDwR21rxIsdAhUPg5P4ePaFHs
vXwF5YEFxzLwWJhP0VUSb5nAJQ9WaGGw6loJQLLcMkf1W32jndpdHwKqho2v+WJg
xItVlJmv7OwrN8d08vRWB3R9kuQC6LmUBT6REgon0v0EyIu4myr+IWE22wzkx6Xe
sDhh5ngfrUuh73hehoL1ySF5RiNsgK+rCoHdXKC5UochChECbtDu67bFOzcQ9xPz
wfcQLGEk/IatbRMH/LCpxO4XbraiRM+ICWqDLpMzUkOzxrBJbaI4H7tNTr3Ab4F9
qju21NH8ZtkFEVPYSVdJjs8JNVZKLMfUuAQA4rY3l+d0NU27LOGVHKLJItqyD+hH
lixae/OMI+O6o8x2RTcQlrLFGwQlc1dSLmZ7h7RRh0Ws5ySTF90Zi5AJWZu/pciD
HP1IP2O5wmwHcqcDuTKkPZ9yUtZLQimAvbDA+jAX8XFC45VzCrQlHD9Dz/QD1QLG
FCUURl0gQPaoT0576++sZHQnIBteAmRDraXgr6QJ4wxB1ebBicfNjKvd8SAIEH6d
//FGNhO9TM5FVnAAQreQT9xiLDJJEVrxKDq6QxMH3CGssPqUNJQTHtyRg3JZMh9f
2pVUdBtbxvnqFHTJRYuLhGQMJt9G51yXOaEAJ39WvAk42byE5qB9P/5YgtEhjUDA
MLUkvT5v3Asq6S4brGpQIgZG65Mo+Xw2KGtEMQ3BhdDA7FAAzfa3b6yfgNXRcYUz
OfHQgQqsIG2+23BIMURWzkL2UsrBBKVP5iMoOcsMOdFmurnh0fURvAAL0WOF+m2P
syvhTrTToNRF6WGlTUJxonfi4nmGeTJyaN4EOobCFgg+P4TGASdDqDly5tYZkIPR
HNBo6K7GkCoUW7m0mAXu0Ye1TxzgF5wDAWklVTQ6LBswrvRst6kqXE33YYHf1TVh
1QYi5z2bGM5efaOuiptkrCW0+NmSHyUd8sqUSLtwK4vt4N2Omsn58lSNo9so+NpR
P39FuQbwkd4jcNi+/9Bcz2DspLlJT5LwjAsq5lTClXs0mkR6WCWOuswTdCCusyPm
gUoIv9pZYJH9UIayXncZ1kj/qBcp3FA7d+qz6JbZ3yvfshQSMEIBK/5K8ttRHz0T
rKG7FmPiOyDB8+bmk+WwfdPt8uEni5F9wl0FBHcYRN2rYS9TCs31nuppkL2sIzKe
h0CIdy9lMmQ2qFMaE2MYJmSbiKq6fySM0OZG29sCmP45ocSqga1nEGqaVZOXyQ5q
dlk+LvmIh/DyE6kXFQLLnyBEhlX+D1cEuphIXPzcLal8bogrYiZLukJ58megzwnI
HhX6K1zz3qCvVX3rXkfnReJEoX9y+uVOOyrjWT+YZFq60azdr2dplyEoJDHEh01Q
jyTsJ7KY4ouCAHZj+jcDGGXHNf9rDoTn+qPbHRJEgZCTRaq1+dVXAPKLpyns8JVC
EK6Jv9S9VThXbOP5dK1S5xysCMYGAn5lzvIGvhLIZux1U4t1saOuMc+lIrUDaTdl
ptHs2gdyPN9JqyCDgQ6SoiyPXf3s6gcPfA2MPwGdq55RvEx6u2sknjRb2S1QtT2O
skTPWiKFQ132JLXeYIXxZwII0aaWjDycmxb45Qw48lbvRgOXrJBXCtSyxV64ZTUK
7KDLaob6VvjnfsAUvH3yDHdKCJ8Pb2zSWZbmOTpTEbPn7j94KrFfQT4q3FyIoviu
s0OIbSuP1t+zIGvk7Xu1MJs8bAMmTv003HUpd/Z38FzhLPKvXc9YNI5gf0pNdQa5
2Scku1V6kXqA/thf+67s4y/LKj7BoQHpwydg5DqEW73eVbecU+RgcrNGnygozCh/
+FPIM8gBhrups2cPhxYxLkbefDKXgeGmxDMnBWALDs/+ZKfbhv/j7zrL8id3jfXr
KMtF7Rr7rDIFoERy8U5cK0h3gI+6buv/k02nZIcpliIur4rda9VlR7ri+tJ1DbV+
Loyy9QodwUGUeGiOBBIt8FMUKugBEzjkzSxdM37IZF32OGfSJPw4zImHfpnbi11T
5dZVMHJtSHNoMg5clPE+H2edb9b51ZCjIWaNtllL/T1Hv3+TVZHtn0m/zqhTw3ub
X1dojtcWAxq03UIC1Bsq7gZMN8ctYthxFGnky4daMFFRa0p23/nH1YPdejk9H7mU
koTo3SZbwcT9zuJGM86ZYWSeu8Y0+A2PA5t64POKXyFjRM1IuPKXBJhI55/DZbiG
pRfq8b+qvhAzQ1CydQsJM6kfAtK2AUPoXWYp/uTiJiEaE4Kr8pgAn9pCokQVQWYD
ArFyypgZYyTL2itMIz/tJropuYxyhTWYikusdNjezcutMHTVffgGZKf1FhPzzyWK
4VOb0E2Dci2gD/ZZHvKO58D3LcnIPhFsqZgCXBuLNLDjTlma+rF6Y7fLziu/qKGQ
jxu3IwC5zIL76KVBpC8gP1eDwLZAwT+X0wFqqc7wDW56BeVbZkzlYgmbkfOwzAnv
Liqe0t6Wn7InTUgeDODszN8e8dJbWdbaj8a6zdO1j3gan5YsoWWoI+VxJhchPRYB
Z4345cVf5B8Qi/+oXWMsteG1W8a8RoxTn7nlNC+0dq/1/XpnEYudufGyDtBMeJE0
brbMIPmhA8D+wi6bvXthTy0WFqS6aYedbLMFIwFeszRw8dxPqpatgB/cPS3Dm7wx
rpkvDL9TDKYhmNEvEAFPteOajwhiEct1Z1wR/BnJqfGe/byrwg2Ctrp8FboRKj+n
+Lgonanau/QNFQ4Ya3I22GUM9/RXIXuEPFgJGYsfzN3rC/u4D+VvTs2efKJW0PAo
KhrKJ/tukdYZG6/aIWabhKG29Xeb6Fj5LYljgg97XIRYH9GmgY6YIGaV1Vsarwie
9lqXmNXTzNoBFdfIAXsNEDuNv/5exoQF2aS1usmhtf+AtFTWPF9DhFuQLuxJG+R5
h4rzDWRZjml0UVkABPcAEVv4PLEcHHM0zuv/JkriVCXRK2eENizIa0g7AZJixG40
k9ODXf6EzFHLhOxcYj/xn2v3ZNDHQgib9KrZiKRoRE9EFiZt0PlHqlxuLLKVJWdq
0ZLPf5hfkeBP7hbmzfQwtpgq8DBEmWBlq+OINAeoNbyWGRsQSBNIqBsGOI7SKvkx
mVuRuBRPFzW8/g79NZ6mzPtaoMTC05F9JlsdtOAuU19Mw4/RLuFq5rEcV+LlolQB
w3uPPLsxAlLZr9rn4Uh++iXJaDsgQCqcVG1wJmj1OzrBowAsnpBIQaumwBxMn3Wd
NJRjNKXHXsecBLOkX9HYV4lx6WbaEQ0DhoIbFaE9Sh+AKxl3u6nv6XpuduqBuU0n
NBhYAWrDJnL/6khNVp41UYgrSeCUhyJi+IYFjp7AZVjYpWO3VhZq7JSSBct+1E5d
VT8nKrjuUzyplPyHtBzJZTl5cJ0XGMTcWvUqmu2DI65NWQ2h+Xl+wyJ66gZy4LGh
yU1H2Q5S8t9EOMwPZFepbCfhk87Q/8/JMv15e0gda+v2v7/vOgANtXxrx672tOI4
jmiQN57LP0s+scrxlNaFK37QnwfVrFZ7n3hxPKxvqRCTSP590hN3z1N9iAP4+2dZ
cDbdqmnxpNKLaRR90nvXe4aWmtiODLht4JdvW0oxxqJOvx52zqT4uXw6tmqyxtXm
PFV5GJM6/2XoyyaCBGMpUUvpTVuJmNucf9ywhjTVLcHkq8RK3vfOOpS/ptf8I7X6
6qOc7D1UmhQ/B+/htgUFQxCCJt3uzAK+6X3MZF2644RA7n/BgpKRqKJ2P41h2cpU
7y8iRWEy+c1GVDM8WAHfTN89pxj5EA+76m3eikyfj6/Tyx2yEeoS5Gzy9Pqviqci
wT+/BGpxzb5zZP0rM2xoqByXcYHWcjtacNgIPKeK64irYdH0SHXK+OziTc2iKgD7
nKb1hwrNoMX5PH6zjlyAhauzJO4lR/1A9iMtWYCHDQhopEobciRcTlpSDG36kp1B
loa0DAVrK83i1KhOkQoFnrqd07Yqv1N7jbeFZto0pVqTgfa74SPZcPignA4Xb/Sk
ctmAKINPlAwJrDTg6lCwqPKtPbWQmxICLxE65AxCU3oKNIRJuj3RIxB49yi+0Noe
32oRV8E5HC+/H8NIbLc0Yz0Xm+qI7VLB53ni4zvm0K/3t/eyu/fB20qiVSwSvDBy
Cvf4PvYvOMQtjJFO5I2qy2QRA8jBGkB6RY02ZoMtLdchnMIDeIujhXTcWyzr26cl
fwP+GJm4Sbtj3ZSz+mrl1C7yaLApppbuAGzVRQNmRZqz4YbiPASncInw09l+sYcw
ttQ8RgrnrX3bgto9jOTLu8nt+kqBz37J2BkUS3qRv441ikYGwJ2c8RjZk1kP4Msq
Gj8OHUA9YnkFEccKnD+1hYkolVb2lbY7tBdwkKFdhbdOZ4Hc7t3oK7T0lmdt+kkf
Wu1IL4wlvZNE08Cc5C0CF1dNR/SQg+qwx9a7TDwIR8UiONbneafNMk97fskgldik
gSrTtCi054OQZ4Agf/06X47SGtPnu3TxiDYQEt/bi2tTv6MfZlr3VfElxESDIHcF
icMU5Cn7Zwoag9ALb1nHClZvg3h6Yb75tNEf/JRZx3fpXaNEKcp2xg7GvIGsLqFN
qs+aGiD2s3B95g5EAFXcAF7hjddTbqr2kh4mlo83hjWuleKAXucYMFjUqTekOKLg
HPyCHfCnGGN0kvZ/CSYldB91Gq2kwrJkbDePWtGdA/+GkL8H4usEImBvzmw0sqbC
0ul3AdKwprEFAD2V2jjFxMjR0sPdcFDP0eSvoIObE9vVqRqEOFw8uBuupUqGMJTe
K7WXJCGib6RHMgF8oII8054XYCcXZ2EkRn6kRKC2xuGJ1ne1p1RkZgDY0kzLNqT7
fSfmwNCJBQszOraZEK4DIqlQuRcoW6HFlgQQ0atZFO5HxelDCV6oOvns0lDZy6+N
j0v8fa4pIjuxxb88QE+4ugsfy3hbMLZSJcz8mmsnSJfdyFBwTPFEfuxfSIndBPBr
kPlgxctFqQLnxqdFvKVlR1eSUquBdS04SWsyAPoBRs5oaJWm5HbBDRStviTUZxNf
u3uMStCUWKjeNlpRv29rTiwR5KBZtByQc0QTi5M6ILJiyTCNKzXLFY/G0oAz7T7l
tjV/0Wh8upua02ib97BPNDdjHBJXWaSX5mhWjHeIFc5/lUmb2JBDDDaOKdAIVBUB
jCrdvOZIxSWIPsBeqIIXzFzxDCo673XUg+HBNTmbmkGHz4BG6ZkrJShUbSV1IXMP
spidSd4WYEFu1BnyQmb2PlN4ez8TwLmb14M+JvDjHPVyDKiXoMpDNDlCDrAGaBUq
GxbCJTr4BXMyEFoEMpfzyDQl4ewIyQaKkPBq5pWl/f6bjwrpIBnDswjzMsK6rbcJ
Puo/EPyWcDtlz6cXLmHJXwDlocTSjIot4RvroWVy7/cmkVeT6CF5xtu7Mzedrnri
7eLq0nVkBsFieifE/9LofhWjLcSX6IOc4o2pOjMwYzKXLpT4OrKiOvR91L6IhVFZ
NVlOjfA9dr1S6cNp5zUqqrc85/8ShmJUHdTfexpQEx4vfK5Bb8WNSu1a00J3NMZA
w+7e3UOTg13KlF2pw2YdS3Xkmeb1u41H80ub93v4HXcxr9Q/oCrJclrcdAS6ft18
ZNSQP2roIe5Mj/YNgrk7OR/SRwXeL9YcohV0Icxkhy0pIoMjePW4APWyoNT3T47W
/7fpue8IEmmNf84sEGdONaJ+3Mg5Yvdy0xHqcra45qEXqgKQahzmMmGs1giwt2Zj
dr29exHbjk6GznPncQY588EsPzcS+4lDF4sJBgGIfGl+2RaZcov28o5NrYYw1hwc
fFZXaYR4mU5O7Mp3w4korbkfS6Qbel9pWcBLFM3YM96Zrbtx1Vk8V8lRA0Y0egRS
B4Zd8gLCERLKPooHeFfNZ0Dmjdjlly9GL4B/X8Ac3/eT0tC3YgYKt6G7zGMam1El
oO3FQItOiItT2r08vGcM4LE3nAwbittSJFBhJijF6HKZCMbA4XRhE6T5Vi1i5qu2
wFSIK4WZgue79TmopRqBziq/41RB3vsBKR0IAFt4pdu3c+TwbALWn8RFWKfsg0b8
sUiOSGd7FITVyPiCMLVj5J5jh2MW87o7FpA5/ITLInwS/I+Uh85cvcJQeZeQIL70
hxtIUgEuBQSKUIn5x/3n81TaF2SU3fXLx5phHU5wLgQf3hPJXUvq7KYWjXemuyKK
a3Th3dkJhgbTiwYCszeNNgHaZiL3Xaf6mRWylVGNfkW6V3ZKiumtYFxL3CMN2lv9
IVKgFM08pO7GGpMSVnLhZAYu387Rwyta9XynYc8Kko7WJ01VWELE+C8Ty0Df2FIY
t0AGS2nwVTztru/1uHdvLMfWleB98fXEm+4N4b5mfXEG6mHtBEmkMu8DBUT/QvQI
7LBZMtXJnnm65YxIYMDQna/VzUHRYzUAZ2AR+al7qj3eXlNzP2xFsTSu6zynpUnp
cbORyjXTgqvsqL8tvSskIaBYBdT4TYx5sSEUV8US6xw6SmVXQYOwLV6f7QpDyWAy
U9czvn6xRNPB1PE1LIKIOfUe6Cc8n5tHTw0RDIknnw/A8BfhvdgorqehoaHrphXp
pXDC3T7SbuVkzeOFSfQclzB3Z/SUAEJdApnviPZkfX/ZI3yfAoaYu3TWsBjF0U09
p/pNRAlqTTwkBtir52kvIoQGOeJKx+9PKCUfTtPKJzyk2SdCuJWo6fpyJs4agSY8
UyE5xFbQcXZayeStXIhb12uAt75vfWQRwlOqOr0LMp5RkZ3W17frfcnlgY2uFqdZ
MI5QkEhnb92OYeO/oG9De8Q04xNc3D0wuJL+wMZM/eM0dR9tBlZt1MJ1J747DeJK
KbLxGO8TkEnO7TFQ2Tfw6TBpiUEjr8v6tNrtwlf3WEQd7TC6Rpei9PSWusF+fYwz
T9mojakH0Dm7UamaSUP30d6+CXEJLSqqGHLyI7vFxcb2ikCG3xwEJTI2AmQZVPlM
UxDF0GPWcF+pHcsUw9UsbxTvIJu9iQHeyrZZSd7ukMNcoNOnyeMTjOb1bnCjBy2i
o49FMfTm64JIgT686H7WgijJxVoTK6hqlfsfIWZPpCQVwCprVmhNBlg5C/JZtE7a
XHSDAS+Oo35RxzeBfHkbP72Gfgh7BPakt96R+JSoGcKM+xS+PBzQZ4Pwilwnwdfg
HRNvAiGg+L8k3TdY6g4WeTMoXFpS8G1N4AMmAsu24qqLk0lFF7DeYT8DC6sye++Y
pi8xvLkR94xXxeR2rGLnzMRb67IPjNpWq3FYAYEkHVJPelyM+gXIYibDECQvVvQy
PJo6L8F8eINyATgK/ltOZYLVevIRA1cCv0PFzliJAPNgboJR1/ppnCV+YQ2XJvq6
A4tAo6v5E91A65w103KoC2BOKtKPuCVnQoKI0dawrf4k+KwspC9IrOyV9iJduhza
C/eZ1q7KuGojOXsXq/iRm9jwalXcVWv3NfR/HBDXkVBrnHG7NgOq96x7mul35Kp/
ekJ3GJN5BoQXZPZrPJ4C/ImSqT+MhOMEqMC5HNqckhdI/KlCvEE3HWlRZ9WGgLCg
ENxnXeJHKrNOFTISmT1AOjFoFXl8P3H8mgYoopcZSnqHAxSmXZiB+LQ9l8KYxXF9
sA/v/xl5CQ5rUQGtWRFu1ciosh25F5aKCZPnclmh/jPjsqDm8DrRTCSLnRGQQBwV
pBMcN4KB0w2Xw/UFMLl1nLa6nflCyljI/bZUaIuQWvzZYgKT//HbBEJoA6vNQ/Hu
4kTc4S/Vk5IW44SWn7TmoCCNwNujnxhDPAkAi7wCu2lGqoozClKpNn8rk6L6Gvvk
4tA6pHb08D4l4QDeBqkP5+wObPd9eKrYDn22MsRngpaCWOVJcaPityLV+xLYWY80
78mMa2Z8cx//ItbIDl8CQuj1otqJsVrM1kSTMD6q2lvYaluua8FaCe5Q9JwZonvQ
S8QAvYlBYzBbQ+YSkej/K8iibq8z/vTJEBLsHeLgyORgawDKdlwR64OSAHeKoOjf
yKXMMhEZhfvnOLYpEIiPibnc+1hTtzCujpJX98GnXUO8g14QpREobmTXZJHNm5hz
uNoYoU9+5YfBYBThwD1R3gNmHfsTytcD2yYmXolNnuPRtm8HnhHdATwGijwXvdzi
OLvX/j+bucxL7hiKLWSmUUcSwGJ/o5XbGXpp3BQVZbbcnFhwbpicK0TmleCiI5eG
Joyv34rtyE9CSvw84lnIiJlQOdreAAwG08MmvNvITLMMs9kFlZcIvlDSDM4uIEHQ
IwLkvusbjV/+2c41n8oWH+yxlZ9/0kQ9lEsibWnydL7JiXZ8pHTuQUln7Z5YqBh9
iUDfPYoEvbm+r4A7L27n2hYKiv7WE/zFoANxu1/xov3tVI44Rpw3jOsvzbdW8LRg
AoCWz5NyV8oMbewJP9+NcJtAoDDUq6KLCMIDdyjtkGZWHlnsHlfl1nfGMb6ckZ7+
0uyNuHvyabLzUw0dcUiE7zMAjtbXnavTjRO6W85p2i5KvRxsCRnFfO3Cft58PlH+
W0uBx2YiVZXhYkO2vu2Yh42+SKaOutV2TzkPH5klz2ZJn4k+JJq4vCbX7xlOiPsA
lF79zwbRxXbH2tiKDo45/S/bw2vQXGVUIljpYXh7++qrhf5OonlBZ8wK2FBTRDn7
+f8LN/y7RK1mUpJfJye3Wa05tydof+Ve1EXu5+akEL6wz7ZOlmru+wX6lzOnJp0k
L0D981FWkqbuWOKOoycUEtid9krQJmGxHlqGtklHhqmu7e4vjldVrIkH/TWgMTBQ
beN54EyjwVKPuqQaXaRnMJF3aqtDoLQ6OVm6q+tgAY/h6rwq92g76odkd6jZHhG/
QCOBXxCxU/BpbmdrPPZ6+0g/9Xj/T/Nm9en6wRfwHTFWZkH54SWZdfeTdP9VBZ44
RBDxO2LDk+0D1PdkO6UoPun05LKp6S/tZ/f8M7JAG9Rx0oy1ehcyGNUFExrI+VMI
LxQPJDn9LQSF4Jp3HXmo4y0/6rP2sqXmED7fXnhq2CcbOgf88anMhcDfe1pQxAJ0
/Bbce0iRXEwWlJGGStLIX1Wn3I7n55l583lkksrw6dMq/qYR7GU/SoulDLl46j7N
wBAtgiYt8QQFgB8jD9bb2tJ1VsQSY+Fx/LAURF3WbLBGz6TCPMce6mCkPplRKoFr
QtwN7nWArOyismg3GHTqX0Th5zpJcwgdzV9laCOEWrGkrJMuevursoOqGjkUL96R
rd/tyKC5zEbAZPDDrtQetq1fn1hGOuU4COuvbqzMcbUz2yzXO4XQyFec7GWe5S2B
3t8pmZ7uN279WDaQvKDryrJeMxJlBKceMf1YiLhkyBIjPsKDXmAj+0ZQC9r2i57G
+rgN6i+CZBOrOA3OsnV7HgI9XCEwPoy6otYBtghwv5qmijpmLPbijxSFffDAmAg5
ImrHyFY70NpvCOh5Z8i+HnPonb3UuCQsA1zod+fES92H71w0WIlwEZmx4Mccpgoz
DS01n3xenL7vSEXiWulweppGcBdq0dlUlgQ6BRgpNNi/4l37l2FO2XdVTsk46JaZ
Q8Bz9w903OqfXwx16UMjJF9pEwH2TLdZ+NNiDg0cTI2beguBN3Bfu9Z3KNLMKwSS
slBjM4bz4+lU0XpvX57ZFvRLT0daAIpnWwkssORP/AqlIu8QGViQVUPCL+RaEn+F
836W+xRMHpLCe8D280P172OCZ2ZU9O/bHSbjGA7SpiBhIB7T0pbk01WoPh0bn6Dh
YVzJc1IlSisIvR8B6wJUIuguGZPM/pPZZEKvcmR1t6rGET89TnNl7f//8C3lhi8O
ZFhmK4GqRpR9IS21VfWSYb4PTFrwh6gJ+N24sDD2LEr+G7hbblok6xt4ctC8Uty1
T7kKlT5Sa7voR7HLfqVhjSbZkI4eP11knkoAt9iVB9oRZNOGNnJo+ohBfAqLhxkV
jHf+/LfmwECbAzvaZMD8YgkYvfNt3tWwQkjRZ+tM3rpWT/eFwNtx3+pgSymkrGES
QAxm7+Ndo/GXiBI+aynmiF6d9RFdnkPYL2YHi9u2We4OP5oQST/PDO80EoZ5BUbU
JALRiz2bE8Ui4ZZ6bsjtfLdjos3Ll/EDHFECxpFRG9q/7TJK8h3qRwlN+6XT/ZdZ
gfir692gzYKpHtM9jBcCY6qRe+4hauDki15IqFjx68x7RuN2NEecnxbkd4UfHO58
xWK3qJIVgBuKeGe7y+0L+Ta5SO+FX1kNTBs5NvN+U1PsB6qF7t0HzglMd2CRpmvN
luKj6QOGBQcqerSuKGZ2PcP661KUJoiUous4p6PFJGFkkMk85pSCYNXzE3V7bokT
ncfqk8Tc4kmk4PMZEwGwVB3ivYV+UMnVhw3cnPlqt1WtQMT30dMi8tejga9JAu4C
kdY2JaZzGO3ZrMzgnFK/O1keceC4W+642H2kdfBWGJvzLhYyvTxPp6tDGvQBhNur
U1O+lPG89zrQXAsF/figysTXUM0zfgTeJBKzG6kcZ145Vt2QErc10q2/js78JTUb
s3CoZEEvKkItVoRc12+inOdTpFLfOwtGJd0SEbZNibBJXZbmAr0PrwnfwEHT6hcQ
N8z4WxUyCs4C4moKxw2rfGnmBHHTnPpyBt2381EoS8znRBmOZaFkti3cRo04CPge
8nBmw9xju5xx82cKoviYQVdNRyBsUpPAkn7A181gkqRpkk7CAB/FjWt91DW2yL6c
Gx6OeHqbCCgYSrTgTVlv9GEveNnNN17Eo78LEuDm5IJoJ2WLZt2mXD1cSdQ7qe/V
ILynXihroi/j/ZxADG1Ns1gleGn5Ov6y85UiYKvqKXusBKh2TX5yw6rf7aie3i1t
meDQTbQjVCjl5yR0vNPyZnV8pY2KFDe8T3QkBIw6FKmNIwGM0vEC0nNIeLUFwkLS
OGyVQ7CkEbw8pZsKlsO6RrDbBJMA7YVVEwZoxJ8Qo82pSyWA75CsJKknYvCIHsSY
8Gj2diiIO5vYOQgyHddZd2LkP/ZzVLUm4UysBCdDjysYLVRXTX76C5KIF3eU5hmD
u5rIVZS151XAyI2zdoNARmL2IyHdw1VXiADkoeCSr35yWB2fWBDUUf8p9mvFUtWo
N5ja5oKL2meCox4vqJzbxp2d4vE36AWCSokou5i+/uzHLBznACoHeGl+WIJjBQYO
BVaiZ1ENpC3z/J83egyDZQcawlDgJCy7znLWqfVPbKlGMu3qiMbytQzylCeFffj0
4Fr+WtGR4lGzQ4Uh9coovSOESGQLBBVH3lIcmwhkX+Sbn9eE/S9ImMXGOGA6+ri7
VraJjG5zRIuCKQz+floEXHTx1WjVWrpti7UMKbhPdOmPok+0jjAg+WoBzRHx2U8K
k40gwVT47ikCtFQXq7SNAoo3M6d2QzmYKLK/iU7sv6+WTtp3BCH+bRVZTShPVKGA
mqByiWiA2ZVtLbrUDAwrObdbs460PP2DZKGzwZ6s8WUNGl6W5HMkpaMzmKLuwImx
7b39J9qsfDaDp+xTz85fUNWbW5LYRAQJBMk49DfrCsszHvvRdLXIh0hyWsv56w2u
WfTkYnCGabfJl4jQa1QECXoMF07dY0+HBy5LTalNmEskbkncsyBsCYZtfKgih2U3
53e+p1i7GwStdmP6ELf9pySZmLEhrxt6mm+Jp9I2TkeMqNTKyhOiDW2ZLya/ZSp4
t30ud53jOhC6h3UdceGmtTglHBwWeOonqC1EkqtWqx2JDxBkEZzVaAhcN5yOrTkP
HTHGI8C926Wofq+fs332Wwab4NOe7j5uGDmUBAyf+InIV/LwJOWD2DrC38Ywabci
r2/2GODdfCy2zKNr7KG3v9XReaJ29aywtgVxUeEAhUya45JpidPVsbrfrg6JpRjd
RvPw6Jz0gPkn/0JotljK3UgUuyUc4dyoM0t3pYedKsO16RZ31dcgIIBJY/CViqCN
RLmyLF72WToWMI/cg2w3KUH8Lc4/ObU1pYZnsd8+Zmh6i/akL/tdnnlMAtxtGKE8
pSe+FWJ7lsylWUujjSaxGLcMkj/qmxaaSzEH3M32YUVLaxasBOH4Pi5dOJa5kU2h
3M3zp/VSgz1yHwAZHwiM5n55p5BnPWPDf+zcCRd5qIGcnasepqTKgzB7jEtNMQyZ
s2QBkqpo8ORxd/xtduDltVzom4pg/q/m8SMRCr/jveb90KqaSis4IZWbQKCJ40FY
ClFZiv7Z50hCiH/XbdHbHj2nfvpVg8qI/vSZ/OcfFI/d1XRZiZJgH2fFZRnoOpri
ZakfI+6NBtF0lPDLeiCJuRW74fXmwjmWxieLREMZ0OdErlMI6CJlFT56j4KLTMzv
Ow6k5+Js3ey+XgpIpE6dpzbAMPi/B3EsKyJzcI1FrJ6qdxGfjL44rE7FH8hi1cnc
c6PUn2hr/RR/DGkPNNSZchH3O+yXHZ4nYT8IyIjazznCl2IlqFSwHBYmbj388eKb
KRT6sn611tEdGUPIdd1+F0DtsR7hQJLiZVY+rIPnN+dmuAt2IU9fOdMUySMmqXRF
+2QeTuZakr4wnCKMiThmTth5G/Y/auI+wzN/idtytSCxMZtguTX5RSfId3pr2gvK
HSuWnQp3fN/ZX0rj9GoegTgRudzE4Y0wPO8ugFj+pYJH09JsegRtdDV6DvR1x0TK
UE+ZZaDYhR0kwsjm1Y6N1/DMUG+WCCTQGd1RkVp2ATgRLK8frXQDos90IztTRS4I
M0x2Su5Ah57UVFSNQQfNqPkVQSonA931xljWIVHNUfsBymEW7r9eqjBIjwCLYNV8
MQC/XAPLPE8EUQSvNVEt8tnJGL8ihXNRQCzEK7pDCrtHr+/RjKUIAwrKhvZFPvXm
lYryWRewti1Pq49myNXP55dgRknlkVzcSl4Bk8A1Mo7at3RBHjI0oKOz9/IFsMKE
ORoy1KGHn4jGo7WwyGW7aeIXB0ONytGuAEjVoyDPO0gYU+PFa4s+NGlE17u/Cmwo
IUh5sypYYtvVAtt+AJQ0ooBcMwXcjD/sDLgyuVaO8Tt2G43WcgQSwnN75ZSou0WU
8Q62myfxGxil3U2WzUrwC+sxQnNwxXzMUJvnD7z4fSGlInhXTh9feij2Fn0RkknI
D4bmHHqA93cuN5tnqmmAKRLpRzZRgo05mz3b5Km3REllLRAdzVmaDqYU6GoXNjvH
OKhEKTlEWnIOmFvVKqkIwTFSPqswCy6JNqrJIhfDRCG2hemtp8/s7SaXhs18o6QH
bh47dTt68CL4iUPpsrGotZNsg4FkJym3U150b7PJ+lr3eFcE99doJMorhid1aiqh
MK0rFjo+ZS0uPLV3Le3lwvXGjLAmUmbd3nQKixwlYEGyiGPVuEPBzV9gnoLFMzV4
u3hPAZjgNYmCs0Y94tKONc1l/HrUJgNMBXdOZDtzt+ghg1dbRn8Va/zuFtvlrO94
sQVXtpytJWSi61+AXYhiBLdkm7HZo/S3E8o6E9F2a318M5zJ90clCyPpTCwYhEYw
JgEBYrS3FUv1eYMjCXv3W+WspO3xtKsZ/2UHc5WtcE75Bqz5tOnAPEsA37XdlMhR
85wgBAmVjfiXa2JXjC3U+oiKB1kk8iaMm+1/BVp4R+nUmpvL3Ok8IL+/70Ra5Wxk
EbsHVcXr4we9+DpsO/4za21UNffwc8tsr0BqQ2YlEzdA51swqlnUxDQ1HeYfDCmK
Y/oFlH++GYE+N3XhZ5Qr09CXnDyGdRf4GnBR2+qPjvOCytnGwIFa+42uJKbiH18e
o/fYlvzxAW3Zewrmsl71n31KywbFnkK87oxOZ0Qb/td+3VBQEAel1FTle+Qedu1X
41PElbR4aQNDNSB57MOVlbAxxzoJrHBlZMJ88k3AXjPIXG31vooJJeokBMDV7NUB
ui82KpmEMUMAo9IwshG93LZ8dzxsrZGna4hcYY0KMjgJTKZy0eFe86nGyY+ox4/9
cO+PJsDE95gkl7kEg8xi9VUj9rbH5XuuW0IfsGtwcjnL57j+a7IvojABjpCeM6Ec
LPde8ADUhYwOu6AW9urFq8d+OMhpVLa+YA+yQEotvpfmQLFyyAxEDotuBFuWl2qx
0gaMYgRtx3kB2mvQwbMh4ZCPXPMBskzBZCpCbEKDCe9xEl+3/ZQhjBjJw1JgO/4I
RW3PLEX4anyI65YxzP0X0Pj+lQNIc6vyHBDqWZe7xbdotmcihyy3PFk8r8NvCFoc
Sh1fOp1cUbzN7nlOybJdSq480hiGSojTyXR9B2tARKmFH7ps4aMgO8YkgqXRXZqr
eV3fNejKOSraQaAjLEmHAuN015aCZvsNtSv53a3YUAHz49pfZh6q035dQ6LBFegI
HgbRaDYKwhStJGmplZPsw+BtnUEx21lf+AfHhH3VhN3PL4+BEdu90GTrz2vceRnn
eTO/rrq/0E5wEeam0qnC45YfnHs7MV/gVzVXXPyj0B6+TbwZLJFFbpOIPSGN3QTF
selsb156lYQAe09ijSRMwGxMgeRR9LzE+jVHKuery1YbwQ+fDoPXX0brmGtjZaxC
DXfWbnqV8RPtmGuyYSWtVNwJL5xTGQolmGBJhP8lo2w+Qs3y4gEb5SRf+M9sNh7o
kOtZFdl99a7GAeUqHzUPVrU2TDYQQ0SPhouZEukUR3vz/Y4LhA9FZ8CBs8YrjOWs
x+pcBxsjzVGmvp+h3lkAZA1umHdnIKr3tVrT7Hy6oRjRayZeQytx/DtvjDFiX6q4
56E0aeFEQ+6CFwixMF0bBZ5ke4s/JSxGTf2ZsXKTKhXvf+XrcsMiVVd9H9/FtITp
yZB5Zil3XNq46wA/vdCADcxTz9DMXIZY3ERYkPw5ziXWH2qATZH4/Q7HLiS/vKZb
LskO8Ii8J1QIM7XIcQXwY44797eVEtXsit7gPWjll7WRQn7JXRqynef8mfWNzLXO
IhcUQK8r6H+maPa8ldtAPB61svHANDDEbs2leQd5muWrcu5MTQHAmUQDkLQtQZjU
InIEyfRfLMTEKwKRNopdZcFkd/Iid2nBxDVfehadiv5zqbnvJM74/SUsyefxAh7l
GcOgHuh/11DDQIDy7GMyv0mZkFU8oAuyZKgLWTs0R2AWvc9uT11KDzWCy13qTxCe
5ehdJ7BjKdvUfz304rQu9xnwMV/f/BIT9UQA5o1QTksQ5UyHHL0K0uuDsm108eVv
b7+7oN4p0ABODh6eoZ1HpS2djybTbBbMPmBEnYdlB/i/JEgcjJb7wN9JGiWIE1mQ
Vxmk/nlL6irpGyZAguZeOqd8rdfskwQLNGcRpRJx+krOUD4DPqeKTsAV04nw4MZR
yUbqR+O5ny64KorJMFzZLQpaGPlsCoIHYC+mJferYOQXpJTbpIR509UHgx2D+Shr
uef4ckM/CJKazc0l4RjXJPiUYMEgnvD9SsWw6kLvvoh3vw0xyOT2PPWgFD7TWcRE
NsCRIhyUOfrZhPU2BVb0/5IuprPOXL1sbUOVY1Sxupbq5pxQCwUK4t7ovvqhNNei
vo7o385ztJ1zVmrP/NfmYVg2BCcspQ56rQryX8zpdvn4NJxduqUeUDXXKz4nLrPl
iducgGgdwbKuegIL93oiYTdC31WYPwopnU0rn8mQz2ZXZQ6G7W/j8xCe9gE6VmvV
F/+Cpo7DUWXkswJKVJUt8A8TkWr9/BcZSKLSSCJIs18A9I1Gn9a1R1/ZdZKFHdrP
JiZgXbfLvjQwAf3XNEEnQdJNWUaEio+XgwIO90mlPQOcmpv1pMKV7xqmK5tie2jB
QnhCA6T8QCZGZ5JYlBn4w5UbMoOQqS4mt2/ISuuQ/L8Q28FOgJ1kWbAEnJyWxgwh
T54AWiYyO5ov2VYJF0G187YNU8n52tBu3z/YRxFMEFcZOgKdEqi+z9Z737m6RxtF
0nMZy4vVFWDEFCygNYLu514hyvXlh8bBKcT4buEpY6Z4ek6FrRvrcqeEsc9AEdOS
UV10bDRbaN8StiJGr2dpLnqxk5lsW6T7oPW2E5gjLvXo361Y86RP49zcSOccYi2Q
rvqAZG9ESN8d0txfvmCVxFia2TUDt9HL1GfMpmN3XBkdzT6v+oPqXaGcM6yng9RA
HqDaMU55N0xqrILOzA3heVeuK5eu3nycE+PFSPiTDEgM5YV2XudScS40Uk/7yAxK
GKI+reaWrzvmjoCzw1HkhZYtSivXLXyXaA+wQXdPj5Mz6OV2SyAG/GuUEtPGTvhB
gSLI95Hf1JEgfUM8MdFPiRXROKYTCxORdlLaGbzoNj9HayMDC3m18L1jrvDoea5k
j5O2MdSwGH5/vUWY0m3OSvhHKOMvjO2IuzcUpvqpbfisFGL5168VNOkmrTGMKdZh
+ZBGOmiYFm1nN+yd+jNSCvmFKBjZtseAB3bnsn1NhjJuvuhs8lglu6FfzqKMDOio
C55hqSM3tHaxbiacgUe3NoAnccWWSFT/2ocNb9S8K6q8/6N2hh32MoL8hdYUN6Wo
xuNWeB1oBmUJ7kkKKR2nXM8JXCbfcHAgs76tq2dCcAlQLpOAnNbBrlcJBBF2pt4e
uvRg/WXPG+gYjFlLhtfgI7t7lCq8delVGyJRrUKi05N4J0HVW+ppNp9ZEP6owloN
U2lnxMk4MFrMlQ7u5Lmp2vc3LQ7sq3BQqnu1PU/bA4/Px6uW3ygp31NeqOHyP9tN
k8zpjXpD04N5BJvW1REl1pxDo4lSdeGj19c7XAi2vbOclmJ75DrgC9CFGNQsaAXZ
vh5GDm5idHzaxcIdfcSX0QZvAjbFYCXWNRJH4PjXV54NS6UeukqLy29/aHgyGCTE
INBI9QUVG+6C8Frt7YTj4hK6DMfufgPOrLkuxAd2qnJms+ihIYUWlc+YBmvc5nhH
tYoZI9tFNUwIYsoAdUB5+PUY0aKUNYEfqmo8ZzRDKA9tm9aOVc6AjLdIIFGeSVEs
L3JWrWK1xbmF5tQ3fD4iKY1FPwzg/750KZ4k48UDXZbEl/HiXnxCtu0grqXtymda
jLyLrR9YK0F+l85iVIpvvZ2OnVEXP+aH53Ao4vgIyvJIFeJgVoQQGAL2rozfyBt2
Ik26yP5ICn6BzoY0rpDd0RLDoPB3gm/H4hO+KY2XLIRWMMa9OYRo9DHDrQv/sv1g
L23XSB7DnUTDuOlA38zRierXg1KXwkWEP3MEt8uxeZ7Psv2WKbWWuIY6KHMuIXDJ
mMSYYW10JSs0rpXYFnjYMhnt2XYns9CJW+eX45tRtdKkJn3PyE/82InKEZ2Zk9Vn
R9xFdEFjzUBmliiJd/8d+zQZfSlT35V5bdPTMT31WI0nX/bbcI1hNVTcJoJyZgyp
G0gKSaJmcqNsMxBmN9H5eae2VvP8hAUOT8g7IZhfclETN286jvykh6jugsG31dQb
OfyYWNoai54PIjia30Z84lmw6B/542ItJbh/NeX09+voUeyA7DkEGUivthUZaO5q
F7MI5hpXS0b9BeUA3MD+XItnBhyufe6nnGIlA8H8FAqDX3GSJ28RF5WZCfrqsZJX
Z8iF6heycrf9h+tjXPMH/OgWhT0+QufTEWMIv8iM11iTKB4BwvXq2z0w3wgbbeH1
4SwZ+FSEXTndSnZXvranVXrSHVv8DbO8/hEhL0QHEcE/AW5KTFOWrhj3Qmg0dH1e
bRNoKHKCMywU7qSC3LvOk59rHBu14Dojp2Ip/BivfDHtW03jccBBr+wTxwrr9ksr
Lqd/eKBwPDiHXoJLSoWv/Nt+icGvrBA77RJFhJdZp4u7/29Fn9yAN3+MBRaweRCJ
BzWXCVuLwEBjecgkQ6dcuX1zXn7qsIPfJdI+HdkVNGy78hv2WT9t10gjAdwkVuSj
c8VvP+BZH6RWUn384uWq/qO3YMEU7jc9zB3CCKTJ3L6peduERakuazGlq2ctn81C
UuImln5jY22+39ZZTDa98YpqawqIj3aLmut0PaavtmLmc5ZslFhz7OCOpRh316Nf
1F9Vxq8D5HbM0jZxnfUo3NShD1BAH5l3YMjqKNJ3f6UlT0gmpYhhVXVcDeGPREII
BNCBJKJ2gNV0Wa/4Ib+zDhDyEp3H1dQTAdyVFPZ8iuL6He3PCTVuO5XNltmHF28i
S7uLq64fcdODLFkaYkI8ZslV4CB98iCIv7CtmJ6F3QEsRNUL4sJOWVo50bpXNG+b
V8fyMfAIe4H7pcaIDVqMRCnJaj0MAk+iO2/aQIWGDDKAHwNsbCqVJMKLmUITT6Pf
qjkpQLkoEp+sjLviN83Dl9u2+RpHanAxYP2IpsvsQKC75aw4ttLr4q/oKFSM0LYm
Fbrvt4/8SycYLsnz3Yj4EgP+1u+DPsLb0m2Ps2J4ox19H16J3BbZVSREIR5BEIAE
2nNrxZyUntAGS/15cr9LHGO+xZD2OQhWu4Z94JbZvX0eF6IuVZOPcefrRJ40mz58
G6K/K+W6wp2qQCoaY2tXsMVD/CX/FSdgvojxU1PH5qeTD/0NyEYKpYDAPXghEzxe
713DbKUQxNcDahijlWVFQV1sX5DfODOVCs8Ag0HUhSsqGEyJUkV3pHmb3bpUl27L
Y76XgVVHbmrWzi9KFu4Za/bT3c9QG92u+7txSHUaoiPAaFb6HSpgl7pawwVAVXF4
CLxfnLjFJd1ZGJaFrH5L6Dnw9d5GR6yIbYFVpvHBiVFQPUibamU1mQeZZwZ15l8g
Z/fkjt9ErVskT17SiB2YjDz6of6ahn0E1gBrh742THV2ZiztZZ7ww5uzh2eJrWBI
2NfWyFHgIifaKwnTJX+jdj/YXtlS8eS6BEl5vaMta3zvAUyXW/NhMtLV4G5LeBVs
xBPZiJMfICrWjPQjQDvLfqxZtZzk4fuqMQ4QHAhQ2pdPbuBbsIvqTJXsxcJt9f04
/Z7UHyDHUnndAHg6uVKVOm0tbmXjtwoe7VuWlg/gt//peHnJDrG4RYv+zYK3V4hI
DBpSjHjR43OfBZ6oUQMaHO/5SJGv9elEcHoO34UHYUdAMKhlQ3+4uwk8D/oc5tE3
l+LR/JFh6z9ixNcauyepFyFmFWbRHaJ5+QTc8Bwnj01UBg8z+iT8mXBTU6qV40hV
dsxdA3i8sCmL7L5b/kmmjJ9071s0QNo8niPKSLv+VJZx6+IIMxpqFCrJEEhqrhFQ
b/M3Zf6Sd1FFoWdLmzz4l5yX0Zxyjphox0pv9tHY3yMrcBclJdFnVY769s/o8G9P
XLT7kD9STdvdQCbtNlK7HJqyFi+1UfRAHQ2DY3ZQRe7nCWRPiOAgBgIVuA+MX2oc
+0fVpfcoAvUv1P4kv0RTPrOoDlz+ENJqp63nCRLJ2yD4oxyFae5Vxw3Wr4Ot8HSU
d3wkELRKgnwT17VTYoGJoJLxSYCF4Z/BBx9HOrPeZbYGVV8T6gOPmz9ajMd1GS5C
U3Y6NxI/UICDFLvztfJdh5Nd4VDxgcwV+RBxJvQQrj2s4mgRBY8OOj/0YV/pXlZ2
i5GmYwHkB3pOmlcnGoXVkKoWcGEnMz0Ol/y/22zLLVNkEYJP1hSOR0b38+cNV7Sp
TFkzQPCmQz7x4M0XlRIP/aaGUgp6p5hriKJDtZCnU+aq6AvcdvJt9rI7wCRx+hOz
xBWqnQxCWqdwoQ5+CIpyB5ZHQm17apl18kEMLyGDqCY1IRuqiUzrxyPJmujgSMYZ
JS9hosX2eqsScjmC16RCB2qfjdM5WdcRgRIqdmW3gsrX1LWcf/RXpGJVdIkKHHi9
fb4lvQN0zZO8zGxWnAHPcxumhVtFP+/agS/skW5QAv5UnrRygnM5FalSuQkkd2MP
BGmXJ90DgUxf4/uC4aKoEkZ/YPXP8qHrwOsu7fQjwSV5Nu5nHTFDsqRjAsh+cv5Z
TLavBZg9C5IktwgkI4J9feNNQWAMrxAuB9ZJAd1f/cXMSr4iiJM3wm7EH1vqbQL9
C6+W138DTH//x/bFaN30x3FMowNa/F+Gc/lIgKXi6bD2Qpg4i4KzNHH1s+PaGoy9
PIwHPxKsoiYRUt90Jh6L7IgrH2Ctke2uQIx4gGXL6c8B0o2yx7NHNvppBPzw953A
rZWi6FQbw9CcYnWA16JP5dQEwOmDHfPW2xBuyXcYdYPx8nl/u0eFfnWZMeOBWvVN
8bQMkr8M8dpUzr0k0tNkFc6UY08JvNbO3cxaALcgX/iRLuBQw6QpZ0TyIPJsaxzI
FPmos5US8OlCzEeqH+aB5X5uHwzU9w0mJ8HA8klwGwnRUCIjFCJuYbGS7ZGnkvfH
z9en0TahiIQTFSrr147o2gD8rAdQcd4CMz7WsyeynnZhKQsfR7qnYoSJOVme/NVt
V7pq5NPy3/g5r6EfvgQ4n0f0VJ0RxHNWtOzEMN+ftG65hVGuuKaXEv9mkB7yBJy8
N2AKJm77cKkeXjcUSH87ztrgyKKVwOJH/Pszj7MmyjZ5Dmbs9RJqw6rUA6dSSmgy
fz/FINe1/wIWNMBjwqprn2w5f/BtqIUJiZca4aR5DAAUU4bpfbkGS9iKr9BS1KOg
pX5qfXv9XilLlipXUb9VPY/qvgpIagYrPPxyKX08oKlhjEfN9PW8OM/myPVPaPMj
5Z1DVZaUhu4j8KXWp1Q3+9E2UDOW3uGzWoLPE9hhIiyD5COGDsjR6lo+s9mTQGGi
bsEHnKbpK2ID34AkfqODVbBU2q3Fe4CBYEBG3klrymXVQJc2rz34Uk1s84aQsCc3
zuXnB5VrQ6yXRzP/tKuiz4P+zM5JNJJQoSm8vJTbsYLpOa6Wdst1sOwhKFverVNB
Am3VUAL6DVugu4wJu7PcrEXEvLp1N7eUr85rbihOSWLE5wjLlC7R79YTxcEhaIFd
ZnyCrky40gf4ryH1RWX0VfCpd+LVJXbVQZioHt7ic29xPQUQNIbF7zj1hPKZOZtm
+okITtTFzKN4ZplUwx6me2W+FrfnOiox4jL0wuauEgjwgQWGAEcSvQImr2hG5WBr
pP3LuCv5Gu7oqq448rVhPMdAgNntEc2DITaneLeodUe+qrPtLfX/O+lZgCeuHYRU
agylPaEewHZUl/2xEKhQC1RBP9bN9VeQ/OMRbhx8TNXd+C+tUARgIHAC9PLerc65
Sdsg32K0x3SO4tVa2I1Sfa9qfSYDCE5aehwqSm/OR1eZcP8TRIpJ9zsAUp8PjhIi
f5opiLuAN9pciAa4Ge09bO4qd7x1XWIvvLaGF4ABTqqp/DLPBiClNb2PHLzxGeMn
Sd581dd9V4wD/O8oMLq2ACqZvk7IU6pE9hYRmf/qST0vbP5Pfl7CSzY2WFfVO40A
CvApZINa7BvDwE4FN2dgs7BUQgmhVkZm6OgJsw+2Sy9YHx/90DZ2ch/EyoFAK8fW
9G+68Bp6Dz/Wln3Dc7evZsN0IMJl/9Pa+AXoryoBkimsPdeBe1IpeM0kHKvyYrt/
NFf95jV2oRzAQGqgQ6IWe8tKydm/9G4rlWhJ0Go0TPbHySEPvtH1F+FgLxPrQjgD
NUeedQ+/VDC1gj7xCL4Ca8OfuJLTWtEgx2IBGeuNVoQtowN8p6qa/DeCun28QbLd
/TzVkcKlQN+a2wxWX15J/yvHk+82ePYoNzQ0QXXiDvA26p3Po+fcP55TYPB/sYoy
dB61HknrG6V3Sf/mg4sKhyd4iFVq1VUAJXejICSpLjIJMSKcxKmzeeyCiw6lSocV
p9M96GWQqG7tZKW1A1KVu5RUrZgdvGR53sHouUkk8aVJAr/QuFf60rEhNBS2koe2
EOOCdnab4ViYJvjazDxlzGYy512xkCyFixTenbdPVT3OBE7Oq+kxTZQFqnFPgvf1
EQYJSo1Zb1+yUW1fjwYYpFlQi+fkYttq3Flx7dNipIZ0LLD0UXgXWB74qKwRuN2c
rLKBpE/E0PoH8x29uS5c68T7A8/BZkoGynZnNmtW1Z5Mf1cIP22U/1ljHVxKtv0L
g5vZkWAZbi2HelElZWpW1BtKFCqPKOM/XRkrK/sV3fXM1hEdrv7PclIDBVWRdZ6o
h9NPFbsngZ4qT3wVfx0lUfJ7NvJNIlmGbwYOB2mMDWGrb6Aym+CU2vK5/hBsfaxg
g5qYLDbs4fCeos/enAEnGy5tKdeq33I86knczhbJgGaTLUs5wHJvqB5jQXqd8eus
c9QdfWi9Y1H/noYQcNpX06WQkXSGsD2r+yCwCp5In3lFvdKDXn91qN9aKdGQZwqC
GbCjhzP+NBGUH7xSdGDu8x2ahA9i0F7dELmO+0O6OL7KnGQB3GmizEbR26j6BDlT
EsU6w4gLt+Jgip6Z1iarG6ZIK/5eyaKh+PiJEPeLZeuWJ/nR/hw5zX7cA7h628UG
PCB68unCclxUrPFRRcgy4sbMRFrQ/g6FURbu+RBFA2je1Px6FL9uN2e5FPa4Bzs+
m6kZQS+LRjtQOq0FQdHgZMQRmVkBvZcKrHEfHS5eYCkDlWh/FXo+cnPMkGh6dPNb
5Ci/1GMmo0XqMMzYSfhuolenBt/O2XBp0neXCqCRjGqnw0yRO+YNPNOjM0P5T3N5
4zc+mAqzqW2Cy/GcyZ7vDf4wvbL5N9ELS4kQ9kCT8m3xccrMBvXv2000GKgRqJDi
yQB81MdGJrThcgNRMqz+FlHONBvdsy1u6nCveZtfoc09VZl3dwIm4jA3fA8Gz+/K
/FJFiVTYX/XQcYJ9TVzrfyZXDVFYgh9mrgccjD6AG3vJ7R+95t5v436mRK3GUrsX
XpaR0mL36EfQ81D4rMKyvlSYJFrNUopYFDGPAumAmlA1U+yt24nW7wo7tJhGBy2u
2nfE9ahwo+VFknSkZVmlzgedcCBNO2CYl5v94IAIUyL3ef5A3cnK6RIznCI0DyTs
PpwPxv/JZu0zCUtqIisLYmPjE76OzXFztoRrPaNyVDlDs+eRdeISBTmbaqJlmEL7
FqR0q2cnzTTg3OHTxM/MjoxXr5pMLaMx91axzy0m2kBlKlTxu/9OGg+JJ3f47ZXQ
ucSLcTVIu14/riMWW5tHwb7TfKQvRsNXahSEU/lGMKFWuka7UpV2Wm/k+2/AMzmZ
TjgLdH2wSI/7HD/U50ydvvvulgaaWYsPcyzlYcDzfNnJ25Cs7pGhGVUDc6fTpHID
B5gVmewzALkkuUEdjlFoh4a8AwJf/0Hu+6nLhE8QDkT40DVBMvY+Iks66Nh0vmHL
XNxBYkojz1hPK4wscTkIDWOQ8/YBeVz+NNb8cvaab9OTcsFhPWcFcChrA2/R8ZJD
KnzCL/4fdopjx+c8VeRCsiZn/cyPYCtdwdeJbnzXM/shiq49+GI7tkadEW6ljC41
yeUZj6DJc4iCsxBH6vLVpiSnOHb0gYhmUixM7isy49UEPYp6Ji1Sa2kMMT6lXoGX
fUUOdDkPU6+bWz0K68DatuyoDayw4ZjrL7TW7wdl/G/B7Tbuu+CncuF/jnHQsqfo
jZ9ttMFtMKo15Nh17o5ZhdPTnVDOmW8USsvPsYnRrfky3m8G/qD5nZ6c3TDfjaRP
YxAEudTOXsWs1AtiXqVg+mc2lW+qrXP0xFrj1Cm3wSCLs5gT10atJpEnLC77vnm8
MwqocKOBYWyNuxpT7Cr3VycQcovM6lFXDspFSCaiml4T3udOp31Czxu7jeHDFNQa
RT627XmKkRFpA6G5CH+F6s26xYViJuKv0MreHnSWqxwJaiEffLaLeeXWbYFNxh5j
wgnOcwcGPDTg+hW5NU0b3Xe4DzL08rwktApZ4sDrqtEiaqPFDBHkaser6QkZPFeE
GZSkUYC+htEyAAHCUH/8mI7P+xCEDfdAXX4nLhoAQPwjxDVD9MJ3fr/E/yq5yCGk
/i9SvsxyX9EoCUGiGuBDkY05mEW15d8ZIVzkpPBu7ugizfWlOF7gc3wtO+j/sAlG
HZSZq6+u7V7qnEBBDAt08o1MFWmrhKPuRYxmw4bRMJNIKpmu4rDfDcoahJh5SKj8
bRhjt+aNT5bRNAnv/EXpjvO4zfSRxrUR9forB5WrFAeGjZBvjbZIGZARgIhRZzvJ
HZ+c6NFVAYtM3qCdf0OJPNP6zecEf/ZUxRiuc8i/uQoXWUkFkpwqzAU3ypGu0GfN
tGodZk6kumDWLdZ2psnENN90VxIAbiedcZkWIAVKjEPoDLoiRpzS1lIXds6hnqXG
8jktZRIUwji70Oxp0aC2mDzAMZfqSVl+Tx6VPZ3ey6YEypgkaq2Go6i4wy20RANl
Gp92j3juqAqF7iKVwI+swGzME+a3brZQe9UbcLa5l5vKlGstXnnsYZjFBAxgNyQj
fVMFRCZ4/KlOE+oby1ihKHRnJAGbSpZiqYDdXr1axWazT1KWturnSgeOJxGCN3FB
ZnSHVHOAIXTq0HCH6ahb/qIy8yNXZtqgQ/23moMgqptg5UwrTezehquFsD6sdZSB
CZeOulNuz60zsXKaalhuCMhshJ9p4MioooIuUGPExtQ8dHKV4MHr9OzMlSYClT/L
8FBxIeX3bilb2kYWyXN9eCSMruo2Bl8aBZgWN2LwlvM939pj7efYS+JzakrS9o4w
58s4YIqMewMhEPI1A7o1rX7XzHE2M/XVrNfoZ5eshLUowg8jB2yHjRHhlsofQoLb
YgBzwGjnaMG1+TEwB4LzUdCbTKJnGUnsyilxaWD4xWR1CA6faTYMmnP/fQo+SXQV
Ebr0NdB3qYWJ6/jsvtWOOMAnK7uf0Zw2nwcU9jaf8qDRvERpcJBG/zwIV51gdOqp
/g7iALR0tKqIV0uY6lc/lc0xzxTyKjpl/szyQWWp8bm9WwTqNvUPSKp1hZiO5Ufs
LNwsbrTQ39Zuek1YNJLiGKexx7D74mJgEOIouGGHwZbZTTk6TQaS0X6fVK5JiFt/
x3KapfKUTGFwEEpGrYckwvbRw5D2W+NJLukQZzmOJTq8I5n8lxG7aVSp/bYNtXpm
6zQoskSa5zUGuj2zNG/LBWv7YVFZXqs5abjWyGO1Gp+IFivgqELbqlw2YoyIjc0o
qtt9x8tMdK18enPYO/KyszlWamOk8XwtuCu+0NjXObMl6MISmIXguxwW0lyIHVPm
rChEjkJhvRWLaYl+VQU1N2n9mc5yxCQqe74bb5QipCttst4tQE1irG3YS1S05ue0
bHgcA4tv3dYTfnZ4c1MarNvnAPXoWOvNJp82/PCB2850Kdi5GMK3hS8bLY+jzDaU
KP5KlnL6oKg6ERCKhJa4dUJIz0c5wZnfdYukI+P8j4dzdqv4av4Y9Cx7kkOc529k
faOs6ZFXa3XXTLpAMUzzOGikj23Y83RE/50KrsmFDvbvzBKj1n3j5zy/C3TXR3xy
o+lhenFexqvFB3svZ1DEXWcKSR7GVL7YUQDmq+gdizvW+i7s8Uu/nSaRWY80zdE/
TvTmeOg5GkyALBLtJd+rLZi9XcAIrqKCijk9Y0MrQ8IFlk1HYTEBzxCxQZkC2v00
vAKJa/fpbo89VkbCjn6VppmpiI84R5uJyShkcUVZ4Bg63ROl3/iI+hPirgtYQOuC
3QJZjbj3Vnr2B+S9MP6Mx6tsYz/2h6ybJ1BVCgwF4dRe0Yfqv/Sh6T9TJe0z2o+q
xqQ+MbmKW4tOlbgiq7hsHZASlQTL85xr/X6vw55ppb3MnxCReouW3eAvjsartRBD
5WSM3ITst3yeyIjLp2LtIA8nkoKSs7GbRP7pFwkIOEXh09SHe4lfgTwBoaxVtx6f
NoD5DODHVjVW33i4lyiD5A1LMLXEYx87YfkswWWYZ8uFqwFS2L9i6yIodNGQv+ct
9DAOy34nnW4zNfeWfWVrH43G8c5KGdMmThzXhk7HCN9XRHy9FShmxfiHjxzrvAnT
1Bmhi/GZYBIju55JQMcr8rLyHHyBEYpvbBMds1be4GknVqqH1dgq/ReS6ghnK+eg
dsXEeLUZiup3RXBRnK6m83+SqGxOlS3Zbgsh3eOa4FMC/xV4DL3ko/y3xpcx6iQw
T7BhCb9wNFSNVWTO7QnlgmeX3etvT8KhwzDwcMtL4F2HMWRvF3tcUgq1o832Ip7/
khzGYHIdPBRRM7OFEDpAk8aH9+6JKcwFrw0Lxwekj7iOhCuWYPmOfrAnumgTLi0i
EGPeWWmBtfgYJRGLc9I2AR6pboCgs26lKlvw/87nLd/k4yynlb5NUhyOtrcHgFID
dcEGPTJ6oeybd1eNlzOHXjXfnZ0H8M+6VkbXzJ60br1eMDAeXzDAh1I5DaHOPAYN
sqmAvaqIVpjeEDM58d+b6hptkNg3VSYFqC1lPYj+0E3SBsOsqmjTyvzPtmGuqCKB
4P+W6UsoFx1sn9yEPnRbYPWR06Cl/vIxBDzTPzgTUIKa34H9RVJ1+I1Bkii6dZzA
CsXmCQIPFrvzA07uzZaVq6FijWjpFJhxUVdty+pLMzi7yD/y8cZ8DMU56bdSmpZl
dSRF9bXExAjmXl//NDWyUmmYdOhUcmRg646h77J0lErH6eE5G0aSEZyQtj5Hk9T4
EwKXJvPK/GEb1zTsUy6erawJPKMChrFLFiMR2AZNoAcrU7Bsf8m06fxQaZwugumD
QSz3fmOlo8w47sRm/5ph/IqzrQLZQb9neArM1VYznQrBrLmi1C7OSwuYEbZE+Wz+
jE6WWzVUraAzc0rGHmS7Czj0XtrNVus3gZtY3KvNITmNuex5H+GRYvU61zkHiDtH
oi2UDmWw72O7g+vKL9tcJlL4VPJ5H5oHutiRUr7Di9jDCAkXr8HwRu2FcAn/R5p1
VelaB0I4fdySkXuAWrXsODHKEWgUOHFRb2iA+93qBzl263pnVZgD+pv/+4s/UH52
AvpvLAPdp1C4uKWlqqrfFq09whloeVUF42b4PQrVYIDpp65dgXCYMHqUJPZK3oTh
4yIwfYnUHSJQsbcV1GHZk8YhwFQ4jAsPwaCGVCUx2HhnRTk004nsIYusXyoUKnYc
IRHh04XwOumZwTYEn/fA8HAJ48Eh7Nu3+V+lQvBlhsVIiEYPNY1FP9+8jb+j4H2I
69PhmVBvWx93/eimUSzHlefosGbxrq5yRyKHKHFedDDUSLgj7Iv3v306Jbt8qNxu
YZ6kv/H3UsiDvsZaWllkwo02bv3KAgAPoVvQ6aFFUnKkznA9jEU5VvP8ovNvNrEn
XLEtkkqbQlRPd0K3PZ1SO4Tf2S492g2eiRL22VFiclC2d5sHNvzKdfXbJ33QBhnc
ECioAviKogHfkuf780P+FCtNLFZO636ZXpNZ3LerV5pnN6uBFgea4kcRx1qE9zk8
4q/AiPEy+JUqp2wGYgFuscSXGbXXRX0zOC9MLJl7GyzaR2p+Ap1TMhXKxhtwW796
47G/BST1QMbaL0wxa/zrpSCbQMar/NurX2FJAK4nQ6iImB81hzH+L3TtDiIxUeKC
+iscKOw1mwC735EchJfZ/5yJ3y31SwfsKYm8yX12VKjxZ+cwNaVawd+LwUCWFSjt
2zRGpCuTViIde7NqKw8efGWTqH2C0J5uGgTOMWMqFSC8VUjeE/L7OAs6+djAlQON
LYM4EdmaGFJqIDo4YMreFIQ/7Bf3NypchutqljRdZkvKGmVj4dg2/IdJru/XINns
o81P5SxVTBLjzw+UkvzjDVcvbjMnKcLa6JMCr6+lpS6jzJFoNmLfcmrPyCf+dKi1
+g1S+l3uaxWuChvM4OaYERVeA8MK2mRWDYKkZqNcX8SQLEkSj+whW6oXXJ7lwGD0
qvH5cmyFP6oGXyX64P/prVzJjjIeoXUuq9OMIG0QCQSb2o3qYz9+fhQUEf9offa0
Z/meUUXxCaijqfIyMXgSUTBPMqSuNl9XH89SIZ7REf/dgYgKAHBTyXKOTfUKp3Ng
HFB344Aq4mW8zTHGiY6brMuknBnnZQ9i1E6rxYkq6gFRZdvVOPVbZY3bG79gexUY
9xZDpGJyOsWlaQLVOgoqE/0SANx/rEl5YdyJ9PLcPzjuCJRYsc0sJU4he8dyl0xO
u1rRqQ9pc78f7p/U/tZCmI47zKI/Gpmkxs/+G4b4Kz+4ZKCFJGH0jufS1fUCtQ1P
OdqY2OzZpb1xQJQddsMfT9h25fWmQ3ekTT5E4OjrH4x1oausk2+PgX+U+ge5UNk6
vRsZ7/+K+icqSM2VgXfp4saPhL/S0YJCuu6aba9SNivKAEDhOljlbpsKhLf3Ut2g
xxHzpYcWOdJCmx5UVFzHAMZfVkyNAtvEAjl2x8Msr8S8v2Ym7ZlBsI0A+GDy6Fxn
CaEXJIgPEJQkwVV7O+wyxaLwu07jZhma0FKUDdUp/kTpTpO4zEE0eGSL56foSRNh
7ffg70RqDRRYWeOPAgRgjTWwuZ0oz3nAiyROwqkndtKur1v4ZrCy/CsffAs3FArd
O7em9LB3i4z78kz/gYXj8gsmerM0Mmig7qmiOR2GrmW3eNXXZs8ry+DOOeue/8oL
E9MneYTAxdxK7lwYh3spfOR54zOZHIIbViCY24EnPhHPyNtnJwtZFTopY3ub4U4E
SKggCB4w9GbolyAUn0qwScZHqGKJ0VnNCXfC2996I1ATeJh5Wn3n+Xi8hgFxA7e7
Cp6xybA+ELwDpRjclHhRDCf24fHRRJzqqa8nGah+AMUJavGEopezHzQzp3OoQIGf
0wk9d6H0NdooKuBZ2Ul7wxVH0d+ibJ3c19cykObmOEoZNtLYH8F+Qz0Cs5lwEfAm
i8oQRtuDt6nZ8OQGJO8HNmnPD//u3CaO6KLHCHfJoHdFTMdLoerZT1uv8UMedrrv
6RiZyLWav9nIyudfsr9mkK7DGL2yn2vRraBZHATWtuB5TrBbxLzV+AtzMLSlhUZY
ce6AlDizO0gCFYQfdPaHy5Lc3Jlqm+EC7s+e0LZckKXJF6BPArBUAo0KwHT18JFq
RimytFDBJcRcaQpn7qZnpT+NQ8DqR3Cdfwr2vqlumrB9bdd9FZL8qpqHNVDEK6hl
Nr+NaXmIQj/7prPIpOEkcNem39orLKSAlT/2VaVSPFv1yCKUdlSKKkVA6vpqQZRY
DMjlWhCXZRSUHkIdbhxp/PuSsKkjw4Dp5HoxgJMHDmQjeYBMhw7AiyKZixV+dlfd
MO4PyGrEgwEIO1F4yZnMku348f1nTPMqJjd4afuSXfTE0T7Y2A429VrOdzwNM/cN
dgGNPBWrwqSHjNgZfiHPn2w71IqPw+xhhDX696AfnZoRgE2SYvMLQx/5mCSS6jlG
dDgHJtwmN9bqmDumoYH9jr0NeCnQz8LyAIJ+itOaf1+70TGre1SNC4D60le1k23C
yYhl5NNt/uLeAC/W6Oi75T/rmrh1reXZq6hqKu8XK7Pp0fU0qRtPClN2A8JiJy5K
N9u9QRAiXsgL9n4sYlayQPl3p46VBt7hMu1FFClb7DaP2Y4pXeHGgO19IshFJvoy
/AokrIg3N2yTLuC+bYkNlnvzecPuE9+fHoEGlhOfGYaTrqAAKu0vEcOyB7r3pEJW
wJ/TV6S8fWqJ3mkM6amTEiylEqrgxIDyqbszVb4ier+Q7DejSGYgDQKRrxB94+Gm
OIdicYHW7jwsq0Wkv6HlMx3NCKdBiMQZR6N5Tae0wNS+8oAAUmoeooiyJMzxV5EZ
lADv6AQRDx95hXfRIqMEWj1s1BUDUCVqGBiOIlgTi2KahKd5Ba2LmoJQE+pF5BUk
zztC5zUOJS2HXt2OJFLzXLS+Aoxogryt0eIMT6xlxKvrguRkBuTnrFSJFK598HtN
b4j0cpHiVXoMNzLkeyoXYhgI6bCYzStJrqRlQUrIM5t+Q/6kLlaYymO47diujKUM
fhcVmQQwXej1PBVuGvgaFMkjKLOWQEoqFZGP4W0fS1fok2Oni6tLOxOCYVjoiw5d
gzsr5SlQxi+D5dBPBtOVwH2Wz6X9qc06S38zt1dHIhB1xhkCNbacXfKpEpE2Rb2h
ZwoK6W04vbrVNX7+ooiBKnxFmyLvmaUt6EEU8Puc7a8/TK2/Uhpiq6JyNOWqDyeF
whTjILgGZOexbF3q01F2ugYWbCFG7ACr/abywo53Fc/tvYT3eBT8lBqVqhvVZHhM
ZuG4uxK5qQSdppue+5ASUFOy2quP8rKbX4ASqqX+fxhS0lSUNyEWUlX2jbo6gzDV
p8OVzpISU2zq/jcjdg/ueZcy0xAIbUd0NfS/zeYqDizrMloATIeHMrltQ3ye6MRc
pMDg9hoZbz3Zlc4McDC5lHkbNYd+GJ//CqFM2/Tn7JHk3wuUqpIKHbLd/O1uJMs3
+jmXlw5QLMMPDN0ANVEkvB9KIio8klfGqE0u8JdzJdYkVvQnT8iRr1yBgmcdByxu
QMWxwc0P5MXVLj1u8FQPM7td9ZZG/mYeLDWmi8ibaTsqaLjf+CvvPElEgU6i3eKi
Nh58zzpGwf9EiadS6OcKWa3wkx1RQ5ZRnlUVMIiX5ApWjFCth/K6D1zNqe41B0Nr
W1P0YkG1pSYA7d1QkssuTY/1yJbXbWFglp7IguVw5Mh3oMOPrI4dHgslOIIB49Tg
dPmauLmJu0RkvK/Py6f0sWJrxuYU7Q4zLmqgVzCc5ZASMBtd2DIQs7x8iic0Ke9E
I+JQO7awbSXYTOY0Nmd7rbngYN6N3UfnvPUi0vFFzzWCsd3z23NWNU7UWAET1XAO
gSrpuUosUxTz/cLL/lPkt+CoOaUqgOaJ3uIblV3S88Busltb63ddIlRPoyVTHdpV
VtgudoWpAVFf09PdagoR43R+kKXRB2UPXp8PRxDwEnNww4pDlTgYrjHpdbxSJV/y
yIagP9CLmBBH9NQS1AU/o5GpKwC3CcAH93ar3yK65SIEsALlVBg/Z/ZF+q3FJZS6
81wjUAhadEXwpfTsfB8cvaEFrXzYXpAfyT7x7VxSOFhw+FrcIe+78F8V5c8Qjwh3
CaX30X1jGoy0EFNB/Wb/gmVwZB8ew4ekIOpMvkzvgSQhfRHLfqYLM/vgNtvsS/ff
/d/zj1Zc+0Ql928hXO8Uyu2SpC1EpvR9TXHSDSb+6ZYoyV2WeIk31hLDH9FhOtGH
vO306LqmhV8mTPRgt8uGnxKiTSHYzuRAyjaYHbaHDMg/oOExFRBWkoY6XYgdSVDD
M62gFQC3mzAGkY+QZJ8va78s31YVlgO9sIMr3wqBgNfCIVA1bvFpXN5qsRVLaRSV
WmP5aWo17+3/tS4/5wXicL3nBwmd2K8TaKa7v1tHSL2puf8MV4vNJHPvKfNqf7kl
CAnqc1M2dNYqWCOJIc0iu/uED0C7RfTS3/UTc1/7LYkd0tWTCY9k6xyq+UrFwqbg
OKvFDT7HYSyJR7o6PPJoWP6VF332or8cb4plZSX5XZpVchT4a1qEmLLmNCH2xFEh
NCzXiwZTpv+wSFUZwldybJfTK55bfhqmBE9LP0aTLzPBolXgAP8+WU7RWk8vKdYx
DOkhocvI1MlCCxOI50bQEojPd5EV7WLpHvudNX5IgoJSn8bDIQePZxNYBluFSh1P
pF9GtPsqnk564wq3Z+8jySuYBHPMtmRIYExnqFLORjK/FDg7UuLsyurFb98QrOpI
ipnU/BDYbZhpdiAIbAcTU4eWJIj7niun7Z/BuUb5yegHc89Pa8m9lVoH5Qn+91/n
Nbbk09uYRUwdJmJo5g3ab3zeAnUPZZzuJdHXIFlObXMgRthyhbKLv2kt6C0B2Wfc
32kXAsKjqDlj3WpmYzHrYwvsVKTCiNwf6rF9us4ndEt5JgtRz2RwyBy0X52QE4K3
f6XPZTqLp2eap5km5kPRtV0diO0wX0ZWVOCEMLaWw5UMDM4pQuacIZeEhslLHFQa
kDa0CZUjesvE1czXdC6YAfVzT2kSzam6j5kmYBcVRqOTtm6cTVxQo29h2lxJnICw
lY7HVRZG8gbGyM2MioL8VgK+vWzCI6ha89GLGVmJTmIuLQEmaEhyzuYeQyXf5V31
oiLqpr1A18SWB06GZPqFzXG0rR+NgI1yHxsrMVBwCLXWA+Jb1RAmPeTXsw2THz6C
OhHZOIOCqaX+le4cGtBy+NQvPRCG0O4NN3NAKu+34yguSXJpPc9baJrO3v+uZ0Qf
v6xkBr6urxTSZMKLY2GVpGQAtwnVupbHgkFCmzy8rT7Xu4cI0ONSOC3DasFSFjfh
+T9u+TRTb6ziF5gVS4Uv4sYThyX19owzI1kjpblKNTwhBY0HruW4hZ/VChYHK2Bc
g0duFxhWR/A0+FBnZSasEwdHHd7fqjjYXcEGBBizbh6Lg4fb8/6dJmQMLk1P55dh
FNip6WUl5gKFDlE/GGwFSZ9hcN7Gaq3Z3s8RpV0eBKBZTFWa1AyBlWd1SN2nLli7
jTw3fN/+oksVyv+q8w6de2aJJWFXi2+zLa8XHi4mFf28zI7r3U8ydx4wTDWCblbf
ZNAY0wudGIUJ39I+6sqMta7HYV1uIoeThKvdGqAlxBH6AVp+VM48OA49bui8LN42
x7N786Yc/8CMricY1uKiSHt1ailHJ1f2rOtLMvgOggodNaUElYM+3YGsu9ilGL3g
40f3Df5yqbKT4v+lTLvpBW22DpFgls+TwPmPpXt63Jduy0roJACLlxqChg/B4DAR
LIbaG0BpF7qx4q3uXn8+agXVWA9EFAmPeb74xKXghI1dm16jnChTQ0oN/BfgpaXW
TDpzA7ME8FszK0SuxTfhFpmlTn+/AQxDMAV79SsYlqh9hdONK0YI1d5qmtRHo0Ou
B3wFwmn0BIjMX1PLQfaqMeMb+ed49xe10jCsZ7hVi2fdI7/iPIMp2S/x+Mbl0wcZ
bSfBZEVfQYNXdzHElBgxgQ8XQ9IwScEEgtVf+Els7pGPYGQoQKrkL1rp7k8YTqRG
v2c2Gr0psJkjCo0XPJnkHEmQut9QHlZPc7HRDY9lyhrRCnuYuWr/ipqxQkYYo+6d
J1shHAor+aIJorHgIZamHtwdh9+y35pp2GvOA3GCynsnxm36BtRDHK5YIX04aCN+
VGlcmze3N+yEE3CV7YqLo4xucG5Jf2W27Tp3G3OmQ7fdNNewaRylqlbudPVhTLZ4
Z3HPsoTKDTbCKhacS3R7hEY/2pYrMR2bUKs04Z/I0GnlHlHwurZZNlOAJ+Di71za
QJBS796Q7Ae4iBe/64VzNCICAZpnmcVzp147b2QCeK5eXtd+PFqnhpnG9db4q8ww
St4pO6ZN5e3AYz8b/6WYRt23UG5Y8ZWkqMmxJDBGeBH6gCPr8AvdLiQFF3fbg0uN
nrbemT2jEurUwQi9S402bHY9LO7Vd3nxrPSRECasiV2k6MeNyRJO/LXc3U75QIJS
BgJv4N3SNKrIkbtaeQnFrKnbWvswpkbtR3FVa9GGruy5QYgA+lwjUYcOrrrp8o56
oxjz8ZJGu91OFrKZ/5ANvMs7AH6eqpkyGXnY94dd1Ol64LrxtdVkUefMAd0WUH6N
/i3MSHi7g8sqksLG9R4Rw5FAF1Bw3p0GghtKJ4AW0w8l5DO5ajbMy45Em63sDzyg
f7xVkbQdl0L/SUVifo91XE3ZmjvJMCl42QESV2QodBwhUC0aMX6SMiUbhDjcHPzz
buzd3VGQ/r5Zc8/oZfUpAqjX5H6Gx5k4oj1iSW13QcksDn9Dr7k7KeaCH9SjhpmH
xSL3f29UAR4Kk9+cEe9IfnzJ7A/gS1b4EIKCFtOmCLeoomb2jZZXlwGqCqa6d7T9
XwpAn0249Hrd6fe2QRt8UWRoORu6mFsd59lOhq9HOsrRJI8BjvHc+iGHN3zrRrIE
tpxLV1EgovxCDAN+rn/0Kkir3Z6qJ6zhDzs9n9he0SQxYDw49abO4iA76ufSGzVj
bTuCNTMAjLk6hoZortIIESXjgA6w+CaepaaiT43HF8rohyPIP3Zgc5egCmUJuiJT
7yxK61ryOBUc4fkDysrcwuiMrHoYYagAVUq/wqIoKvwq2LzZh00MKa0KWiskK4h4
TZDF6Q/eIkTvw1tjVgvWm5mnByilnMYWMpzyH9MDBbDitk7CcaeOCZlMDemwF/Bb
0grpluu+Qr/SAWKkLTC9GoTsmNCE5cUnletdb7X7gooNf3FKX2r57aN7Aazke8sP
+EyNImPdInbQTJ8KDn/7h/gMrcYlraOJmzvEJr2yX+bSOaAKAxTvB3XQCO1LuDqx
f4Ew//43/np4JhhmhfIFqIfgSmA5jSsMBEjMUc8kqqbEwtv2s8J9cRU+dgeuQLLi
SrfLUF8ACuRFyUO+Y5SXnO/N/KYsVKo6eRu/pDLxV+jncYnl5tYgT7PIpEt6JRaU
vlqqteU4LOwWWIhd1dfrEcvo2lL98j7bYN5w1WIpoXWtX0DDLJHPf8zcp+MV5Q9K
NW1IXeBFEE9gV8SSLIx6SIT9rKfqGmvaPQDBfVdF6atBZ6ZQcpY+PZzeX76v8py4
z5fgLxhwJeK32LerHVL0Z1eVP4Uw5pIvCd7PTZ41V3XW6blDYTjBPoXU6vNmkxNy
dNSh+uD3we5J/rJAJprmTvoP03fwR401uy+OltYU5HcycAtteMJHKqkdcvNMTzXv
+XQ3opLxhVSY5ueDDgUU6dW7V5dJhsL2u1wNQbjCkGyVFjmqNQMtnZtzd2PEF54X
KpFfJz44v4ivBkY0tR3nG9uubKg6T2+4EEr1sq8yg1f2l3WXPuft1bcL4+3qGe/V
xyqRHHHfFqolv/MgfsmH8ElGvE65Kau2nTFCgZTNZqV+sQ2skostxcju/zv5L97N
gvyNVqmZMWqtlWjP0Mvu1psu6u0LSgIHNy0p8Npik+7m8saJiU/yaZM7R9OrD9h0
ZAV7HiQ8JWhHGGwUsIEP3JyDth6SktCucFdDjCVvHGwq03D0KiQHsZqVlNkJgMuL
yFx37ICoHwKu9lTDqmTi6smHr7WaqFUeWx6zn0CPnThQQv/HH4nxavk7NwaOERsV
1T3oFjBLDZ88jAeI1BahuytLSlGRdymwYOA28tsTHAaxowzJEC36ARBWiJM+FoSz
4MiVx/TuFXATzh5DMPIAMn+Zrf21yWl9ASFckHdbDKB9cHwY4ml093zWhfmrLQ25
TxuPaFA2oKEihMVAWQhKR9xFSzYiItCU5voQdjx7SwdQGQP3XXdu01QeOvI7ccW/
gHHbp37mTEbzttwcpxGE4qyWWyUynulubn6/KBYHgighaz2KhSW9C/d+HxzLshnD
xuonWjX7DPR/YBbthS8Q/bqbIz45oHcnkXIleMg1GGuE2rnEv0fYcQDQTmlEoid6
+eXMFDb0VfvzkppEw1P6HQjuV6AGdK1GjHc3tRIH93DOUsZMitjRYZljIVL4z5gp
B5BgH77DOpg/Fo7PgjI79W/HTuWd+wnxfp8QzTS4ex6ZV5gCy7/5LZVDOraIjV2s
slcWUbG4i9i3qHXDADIi0UyQCAGbC/HPqHATvdCbkgBYb936YsZnWbofxGLq+wGG
Bef7AaSJs7srENP3dtrbz+dd5ViksCUlhPSWmPWx71UZMahat//JBaQQEzzni5U9
qgh9fo13mnvE9NqIQQKuH0C0uiOfoMZGYjfjwnvmoNw1uFBP2fqNymM/jzog5q8/
u3dVLKSEoBVwLfPfxh5sbYsKi9Csp6CsC0pv3RiyyECI2Z3e+nLrPBGfrRyQ4k4c
oWtRibf0IDO8MujEVeZjBFWMJQ0TdbvkP0q3P3eTbpAFz42l3V5nUp6EL6+UdRwa
Xrc7uOWj3mDbmoTIQBQu9EJGL8UL0ejpg5T2SKCGmsnwjcTxs4Ijh1+TcYvoW4Jh
voYh4VzbuVPOIqRHmreoin41pTXpfKGT1xGB2hOEncwTsQ5mmYsrS6eYrF1F9YOz
Qvz1BG3+ib6J5yeDebBm+lNV+et08/EyQkMqaaelv5uCwb3MgQWySy6xRoUGbi58
LnaXMyg+izY80IvodCzsEWLp4VpoHRCGvKb9IraJN5U4T+rEMzxB+XVRolxde7eK
eNyhDZ//dV74jUD9u+I1FLbbtdL/vEchGNcNiyRUo7XN4pUM3e8io6YUn3TmVGf9
p4HQeQiotQwPmAmiP1WvJCAnA6RrWu1UQcrW0oEqfJWhObocCSrXpjJh9qRT8a5B
UeKDin/c4xGz4HagH7EalMuGHisQz0sTKwLvOCYM8ALbbzwnnVgFB/oRAkEqAKy/
3+weHQbDZiAJnygPo+xi89dfczNa4y79wuSMh9QX39PlbcP/7d5cerHWKBzBnm2u
Eml51lokPBTbxa0B6c52e795xvA4kGAv5SaZABLj5IsxRifswSxyr33NGJlYUXb6
azHpWwbQLl9fDuYBeolMbIfta32ZjnSC19vk+rKTwmvMsMm+Dc4E2zwKTsXF5q23
v7jCuE4RzcrLNLJLt+b2Dx3PRCmVI23Zsv4Z/slWBZYBiAXOGGp2LazeitDHMlFY
wnwzzRiqKIbfEWtRp7RBlBRRp/H+Djhr8nbxFzsvOqckA5YqfphWCZCNr3yjZTQP
ccuUbWDXlCuRj0beuNMf2cgh8+QQv8di/9OCAuIMV2fQ63Z0ASLoOr8rJ5o7SKhp
zXqT8cr6EiOFfJKuW1vhSOEj9wlyN3uioiNxWYb3XAe++k9i7h6r1SIqVV8r/u/p
6HWApxT/XiPrJx5O1pUL4cBRQb3qQuo9Wh8WcQiHXW2ywTnKPhDIos6mM12TN2KM
yxPofv19Lsjr1yPylmyrs3f+iiaqTHpeX9w1CHkWYh8NYc1k3R5UBxJLpaTxdjeK
teG8xkkHl72PpO17u564iWuFYK71dd/Middj40yqdp4au9QceiY/cTU4tcFT0Ta4
qzsy+YyanG8Z++WUP4H5rIY2QZF8q6xUwNcYe0JNHuoLmO8Gfc6SG6+TIHAtT70Z
h310TSe/ntpcxGE5XoLq5fAIl4jhe4nHehakpGmzMOzmD31ZFnRVf904tZ0NdGUE
15olCUUHtHZpPUQ7NB5LsFAC7IebhvKgVbU1sPokmXoXBihXnQiAPp4aPcRtCXzp
LEXl5MeSoZzf1FO1wc4O8efw/yP9ZwT0JaF4rq1fakhltCHnXibVNNTtrO2RbZHd
YYrcQoZ2n//2qaScJ3SooST+D2Puwdov/1NAr/PIGZ44KkMad66dEoz420+Rqf7j
TYQmsFUQN+N6GcqRiSoJowUqADopu7rXdjKRbWsOZ6B8qlOSiDoaoREmq4yq7zPk
Zy70fhztKXRLS1rzLnvQRlB+V3NZymqwHGrHGffk7dOvxD3RVo2WIh9Dtnm9mAj8
wz47+rOO7r4YsEPJoNcIbdbiax2RiyBiFcA7jlADmv8xiSovgkpNA5YmpTRf21b0
+l6Fpet7Z0CNTSyVtACt06ghuy/jQzOsvRIgNjBXc/wQWs9nFes7aY49JJGh5QTg
gZRjw7Ktiv9hRzN6s17FoYYX4tfK/wMr+N84g6xp/f+qRHpR/qXM7WJ5P5TrTDvJ
p34UlAkG+GByyIJs2uMf0ALaKkoUiA7IkmDYmz26yz8CHYVf+fSLVHZ8afZT4dcd
gyQNk/MchvdropDJ3xFqcWrJlaqCFeFs1sGp4mjvdZFYByzRugqlPMIi2bjItCAS
4j0ecAd1ev3iv7bbpGdwLi8l+3vB0L/pVmdhcW5+uzYfwlVpR6JoIxpbPD2Vjryt
HVIn3MtZsjj1+cFK3QbFa0w6x6l+PPX+NNVSejBG+2KjYvGtIdw9WKZO+qZGRwYA
UnVHP0uBW1ywNCh6+/6QImeYTckqN74l3r9TTvIIWiWRvox2ubBwQdg17Wt3Ab5e
YGQY6nyHnT3FgK2kPBHoxgPytNhHvxsbfxHXrpAhC6EDKEA+InFvcSQcnYX1Ck3+
ISaOMdrJjcICXxwMyXIk/3ydFdvLRNiL+MkZ4ES5MjNkojtwlkj8EKhdtVlHu7Bv
j55a2RVSX/WNkBd1IidZ/g8o0No41EVi76TUSE+7FM3uQAWlG6Ps/o22edW8vNK7
utOyG9wT1UKuBUFJGtwOvBURoRANwHNZjmWzv/TGCoPZschB43lh/tOjuhfi/T7T
IO/YFrf6Rhjawo3j5nnc2ea/wATtGcwfYVxlJ+3KzzK+HCkPvgqYJL3A2iI8zJpS
G+OzeepiSg3xc7CwdM/48iQWeEMf4TXdzfLNPitEaldPo4tzvkMyBWb55/fYl6ur
FMqsr3XpMxt+Kcwguqe5oMPaJS5kelTFISNSW6cE9QiDBV5ORIKoAUBt/dmISuAf
0NL69Pon+k6rPlGb013f0eSU2+M8bmK27yduuzcO5s7zp1OO56XyIGMOuPg6T7kM
oBlUdCdYvU/WSLaDRMWZxmMj/2ETS/IynQ9VxdwgTlWKMi+PJei0GBWcB1cuY28e
zSHjQ5aZaYZ039028p3h8Ml4Jz5boEUcVUUlKbcC9ivrM4vTMGciBwS8scDNl0Hm
mWHIxotjIQG0wfiB9Rv8IR58DUKjXcFcNfGZ3eehBPqRJoNWtQxQX0NF2vUTbgPC
xB5TDD/GI4J3XhsBcZVANUI9MRDqYkYUUP1DCSU9ZBhELzQ4G9Dj/UVrBVem2gJS
oBoJLpgccuGQ8Lp3VWlejmV9fbzxZ+/JDaIn4VGWleDyUWUk3MzEviA3HwF3hkay
emlNaeOu93bg1fTu/uC6fYgcMWIm0oJyYMePenxw86C0OlJTT8QNmOTFC0l3scq4
rGKzIEyBaXJDa0gFxuDGiNnT6usFAKDTTiaaxViuQBSxPXKyH4kFo0DTg8uRl1X5
mZfjRymZHqIIB1D2lK8H67c+viQKUPSvFRjYsNVNQggT7sLG/cOehcqjYlRG0num
h8e0FJqvfmZJcdjZ9M88ba3BfMMkbGfLlnUkP58zNMh4HENerOxRo0zYG0e6/pq+
AEHbPfV5klI3jqKuBI0k30zdM/eEwK5f4xUOqme0rxbdSdC6OZqlfcfardAKvZHG
jawWgAJRY8lwom3bdQd/gMtOjyKb7ZdquxaBMann4uNvoNNRPGbgfpd/9P+L1ZlZ
T4kK95h8pFJdmzYyXDxpHjmPBek24oSKTTdYSwQC+7htD0swqKu2VCSIXjqRtqTL
wcWHb0lzCqkwJBY+mX1D2IwldKC4nFxT/eKu8UV52ZdbANUvyR5v2hFWIp3s+yBn
A5OU4JNY/d7vz2ejNtfA8QAIq1y0ngKNmq/Yojcied9Ciu9m61OLV6Tfh/UBQJPI
9pmd0lk89RBLhvdipefiM5yjT7Kx8EXWZrLqVpLLRhfO7dLkNa/lGB1AGhRMe9TE
L38kPQYrrs8cg4kNaAd3pU+fWIVmBmPX4Ahb1dGkhjNtm+HQdU85wXDXH1rV4NBz
tf3MnYX5YQl5Zbj0k7Z06h7alNc3qPTtFi82yAtHvf1CoyZJ+Ld95jMPJJP+nkMz
ouJ6ofpBg15IMbZtDvHij0uVXIOd3ppgpSuQ6rhyIhWJLkATlXNyAvGYxWs+jd4d
J733qUP7toGtLXiOMvGvBEnpMUQ4sYHHaVHbriFxG/6x11PnZKMs9q9h+Mn5nJAY
VUH4k7ATS6iPQtwUelxKnsA4qCarhlkahd6HL1Yi/WlEjv63AePErdZqX7G0VIGo
HW2NVuQEzUHiYROxrvXpymJI3+3GOM8gdLHLyW75OedjpLkFGZw9kVx/bfKjkOL7
0+oBo1AanScWLVMiqOfO93R5itqjeg9QSaC9taeY1rurdkBnrjuetjlSLhUd4Dai
RTqNCtRn68lEXalCIPbYWcM8BP2Mu8YlUjnDvGvhsvj1+eEYcl6UzxvG/SVxa/q7
omutYjIOT9qsYyGSEFlrTJuL7+qQs6hUt9SGhluWpEG6lk+UjdQGXlbjknuqC2Da
Mfr7+mR1Zs9zTsZS4cbxjjkbBmTxjQY6nviuzSOpC+MIVa1nEYc7nKud8OnyPC0v
gOURXOtS8pkNkSTVqGFmBf6aEfGQe+zPfal2XzbLYbhzqCtA7L/59fxno3uXYYe7
juQq2cM8XNNWoYCqQWE60Ixqp7i2IWvJGDqgrkrkNOYk9Np4iRovIXwo4Os4sqDn
8U1PknOlvcBYrqviFqGF9F7Gn2AGv9kGsw3i6youaFjo6mmJPrcYy3Py9NhCw4TF
Vlc9w9J/0L2o66R9sSzFwsR5JxWbhYWOkUTGmKGinLVDHbrGHZ6VkVM4nCXQOA1i
QLZbEn1Ot8JU4JGz6c8kMqom8oIeyJumsZSyUUg8rtsQF1ZWxofITJ6QCdc1KLt6
IbgA5U8HyfsYpNmfQdsUNsKxdGm+MuCxmsWNUsWVhJY1acCshtF/HZ2KSe4+mqod
42PUMlIvFer01vCo41nqHPOlIM6VCTxIicp4025RVAzuiN4fV/UMdDGgOOnxIWCm
5gVtD30h2WbILsmX+yKwcwgKp6YLcbJ+c6erzKcPYn53jKPRt+bmEZ8VWvvwo60p
bZkGRqMXMy2gbx8qU0Ed/VgnV0U21U0EJDgw1xheiprOIrpGv1xjpgMboRWLjvrp
0oWSFFGVCCrjUnFJp7gZ2MvlhH+DSr0WIBRddUkpJNLW9JoP+Tp5TpudDASjMef7
RTfAiSqKyU2ef6DZX3MjjmmpWubws/vHYQcayOEZL2iMyP/6zGE+HKSeqaT3C4UL
+GxUBa9H9ag+GUgPFUd3g83sqpiDH71cc9deUe0bPPtBTP8ue8d9vEpwFaAa21Rp
nM1eLVkpfk6Ftrq2d2rc48BsTkXBLBPOnmVhwaYmTvlLLpfImFZLuAEZdZe5zT9O
qli6rXbi0boi8v97ca5AcXz9wtMp8hV9eIqIdMzIaBjKZlr/edA8uXwSK81OOZHh
3MXE+G+A05297kazXoB0aLQaWjK/22V9hoO9z3CzW09Jn6s1MUesE095/scoxfXa
wVm1g51KK4JEvQ67UDrGSrcBIlpn6nHVQPyEyQ/qiGhKo4KiCcOaFa7P7+43I5Xp
kxna0CRiB8FtvZIJJj+BJxCk/yJmTuxwXQ3ziPwcogHV/KqNbYDhpukajIVQQm1N
auRbOD1s8QxO32+vahJuDXt1Ff/V++oYgSj9rn+F/CbEx1s20TDdVqHVc4Zd3gLJ
M8IZdLcZ3y3YxlqsNDPmrgBzUdyrHgsEoo3bQrIUIB4GDoUO/9bM3oIklojZ1Ap0
vNpC9Koo3n5QSKZQxemORzeK2aMWqOiHxU8KIxWKktYvOwOGobjAo+Xmczw3HkCK
lkM7m0YT9q+armuS3myymTqIJYXXQ0Wmv3FhxYt7SFZkthCTZwxtqSjgkDynW2CW
PqH7ub1wEsN3XTMroGBBNMU4UxThahSplOGdLr0KUhj6sTF1kacZ4ErBPsu2xdNX
xNbYmMlMdYdzlnUVZjtNrnHIcyLhHfJTbzZvyGv5zDApf/OEjGfyGeD+/5RzC/2k
7Palz8kPjBTm57A6wpiBZExyRV8goMUqXq8uFca3QJG8nGVCk7M/ACa8LxHNqira
JtZZ5nazaGYf0L4WC4hD0YbsRUxx53PX63ZAkn5pBoIIJtCtCiq1x/zARbhAnkO2
gWlVVjCa7GWculnQs0lHjUqSomXr4WDn2nHQnqYI8C7XGtUsCCQ9koFR0TLP9UuC
ck9GJIv8MpWI+6LRx85ALVpiOpuTgzsoAGuQzmSWVz7YDe+NbbVL9v6uFrYW4jWC
qz0xJUcoTkBZXvdFNW1N6hIxK96ak1bcF4Q6K7uwzyiX1gJq5EFq31x7EtftonFO
709bqBxgNAJ29e8XEu2+ZiyDS85J/1XR5YuHm8t9AsGvfoqv5NWyMEgbqFldpiAK
P4cJdn5zZPVSLvflxx5oHozp6SWpbwDFd0RaPuf0JIiN02AAFRg3eqAbO2nS9Pfv
G0ExHwt1PjL0NwW1i89wkusO59kkhDXILyNEoFzipJZx7+oOaZEFfdxhDbe314d+
BxhSv4nvmXWxJPxt6MLnma91aFCgCtfeR4/glBvKCuMVvpwBsKbCDWnVghocFTZP
+qkbqClLj0guzooyGLqbM27o2OcZ3wf2y3mPu4ISXFKwuYE7xY8EROUOpVlRV0rB
L/wa1w1OILiK2m2YIU1Xzmbnz1Mizlq71ESBAl20foLhdXYRmVmxHYv25P3GFURG
Do9ZOnwoHEKKIUOHyXnNTWJ1KpErlWB1iYnwG1eRz5FZRibUTRCkJEiULpR5qzTn
ZV2tM2b4WxYepmOyVuXy9VkDx8U0UovSh9Jl8tmZsw4IjN+Pb2hUygXWQGlwrvmV
IrYTX9jNdQ2AZelzewxAZqIYqK5unc39Ju7XxxK8040ho2WUMiYFML3r36UGI4I4
Fwrky0xIYInoRz6t5kl4eGfDsPMcW8kNllypfNcu5WdgVvKAMCjA63ogw4IWZhIh
SQtiHh2FCiBJqUa+KhidnRVHwHYNRX8Tu/VbCiJuJuBA40/XnmLRvARPlsPYMCG1
AKFDDIkD06ktoRAsQFyCxvRjw+DC1lTSguvGNfVkpaScvJ/9qcCSBYF8biYznGQl
96A2M+CwTmsLtUdjyN7Xtr9QA1W/V1z037go+Ezi7Uh84q45Q1BFJM39o2Ur9k5d
qSWn+4ZthX6KeEtGwfieIQzIP7lpy9Sa+EWbA5o35s4nwzfgChXByBaRoRO5Kc2i
3xjhwi44ZkzkYbQmiqswNu2u6euFsZt8LIqzoVoWGv6yGDM5dqbtFHbcTnOUAnQ8
O8Z6/jTYYcHjVO2HWBMZ8FvoJD0K+52AK8DvSmawSSYLX1NTtmf3FUBvZDsck6kZ
8mEewF6Zec5Ewo+8DI/E8/s0w/zcis/BmqjSfl3mpy6PECitSBABr87fUOZptxNt
9LUC0TTdq5mT/UJieWiOMceAbPtI3aqzKGddyNptKRY7ZroiyBo5gOwa0rvzFA0Q
/ITTGftiN73VYG2X/qCKX0wRN8MHNh4rNz7LZm7iaDniOoXFURpLJteqevOWZTU/
71Quy9jf6sMQqujOedJ0pI2gzf7LETZ20JYxz/4XfdImJO0WKNv/CDXKOnHjm8Yv
0GLjX1OlXX1TUXfCcAW4IToO7CBvGpV8lacFVIXgajEC+/oje6NZfZ5cWoWlkIby
NJ+6AxNN2GvnklLVq6kpySvgIH06zdG9xomSKRHYJpjtZaxYVksGjxHJpxWAgdr8
FjfgnV0MOFjX4VoQ5uOKYk55uEl45Dyc/TYViMIAAJm3bs+ztazIUrFY61/0DfUV
CjAfF344izqqdrqByx5BuQGJNu4PxWexeEuf0IKeA3ni0qinogVvrJNKgFP/eJDG
mtWkD82o65zGO5mEr3GwCx7Gp6Bv70hCL7f7zHP2FUwHXFekWt3xuPMFtRiqm6d3
pwNjBb455QLke0iL+Dv0VYVG7aXxtC1Pf/yIHDsKSEgR8yB+hjKgAJj/D4K7aYS4
a7ZbRBRntbqgAvh3nNmrDSB0+45BA7Ue9UdHb1GxHpBFeVGaGr1HgPFAcUQPUapo
gcuv0MWBhpuPiBtFmj07ayBx+OFj2LvshIr2Br8+TyOVcxhfYUks0kOWPADgPwr7
QFsxuZjFxVgN/8FXxrGE3QcV50XW/6mfU01PozISVVuObqZ0jRSHuI/XNNrGWNF2
GyCDU6dKIj5nCkAWd2aHLK5BpFaGHk3xsYivckMhfOMPr1iMqQ07NO2TpTJ+8un/
iYo9RhWV8ewAJOHIZSi1bKoqzQbJdSLSO59eY1UPKUFEYN7aeo8ILec2wIABaMl4
UAqUPLvUvKXVGdFMDMrfjB8IMk8uOnDd8JtyWI+Uw4s3G34RPIxH84c2lL49jGJ1
EymLhZ2m3tyvk7EX9/9Efhxi6j3a+gIQJWwcxf9Ml+U5E/OcoI0W5QVzF4Ab0DOp
0apXOIYTG/So3ui4q1W1v/QxEHRugD0Me8FE/D7E+dxA65lYYqTkrYdyrgExr7HZ
+GVW7rERdAUHKUIjxmoDiWaK7Ve0eOAazklD+gCT2Ck2UQTCz6MdlHZZNuBSMV1X
vidxt7MqfuFlawd1LzYI2jtLwGiAH/ddQBuRerB/WDyqrC0Vzk+qal1AxrWYhwti
BEqYSR1LfktNDc77vnT0ReQ1B5QrQS3BM6FeItFZDsVeD8L+Lidnsji18Xn+VcIA
r365ujk06zKeMEJbZ6twk1nXPcZVQy4Ran/zXuidWdJ0Ei91kUXC5aq3FfQEVZbp
n/a3I7T0CzXDWUms4HY7smAgRqFlNKUY509Abo7OUPytvNW3ZY/xpSsiVEihFyL/
oiZudL0wKU/TatdHZnhmpjOzwNo9b4RiqQuBhcrXmJtN6NOxoxsSZ7PEBt3zaaEZ
Ewu2NOzKJ3wUV/U1RV2S/TFzmi5G5ZLtm5nZ5VGtNvi+nn+YVvPLB2yR6EDgoC4Y
a+t+aLdpZ3/ZwOXevEuWl06L7Biel/9gOjC4pHUMyfVKwI3TL4iQ9FJCkofUEujn
5E3mDKbxnCbSGWCkBRbs1pvj4yaifWnU3DVe/YORUtB1a2TsSdq9bzL4uGdcMVze
ZYpQDCcxuIP6isYCyBUJFJl4IJnQWn9iHYJ4yk0Kb6ufOntHaU11KyDtiE6UX+sG
aTG0kmvG2pZ+0llFctTnbZuIcwtDzaQ80h1GPqg3inynDQMkHMLoBhn7D5rC638G
LD5CvJHmXHsDVgXH8+daOOiRqOglfnkPtQZXXLi7YcyiinRMrr6M3vIWyawDaen4
AFJsjhwW2kvAU0lJSyvXDdGV9A8k5rUITcjByOwd6Z8V9s8aviPow+cwzPlM6jUB
kXUj7nbpalf+HyrxwfH8us6VBrdBLW/EdJFOKLR0XREKElUVVXxTMpFiSl12xz7m
IyROSjSaoyjH2X4OS+dRjTHP2Xwhq1iwxY41azBNR54Q7MfZXWW7cNAfyBhocTwX
tsdq9tY3wBwJ+iCFdODNBjkQXQkuH9vlvr2cvazh2ZapzhevNfy1GTBik7tvH5Iy
aphjXPOlT2GuNxEajLmvH+DZU6P4lfm8Mte/H0tMcue+m+0lLH5/UzNEFkS5cXmk
PUXOZ4G+bK2pYk/1Gv6czp+mgD7esZDK+i5WAfK/iOKKbJYBmnmbQqtNjTm3aPx3
XbgpX3pTGeKzjcKAgZcQEOs10nN97mjSHrn6M6liQDALvKGbk2eaNirINfYP1Udc
FsBpAqtfNKSyhhVWzlCmFZg91QpiNPQbq7PM57HhHlPFogYmmwLA3/mYVVLJldp8
3cJnwUsa0uXOyhrLOQn7NUcsGgLopi0Kfs154M3ND8fE6VQysbWOsJGA9Tkn1yXO
WAG4qMQPQCRYoqqDcSL6fWilTvVUSTpBRBWJuPEdWKw4kXomq/zJUzdeWnC4dGFG
LwD2fIkzi1c8DnYzbkz9EfAVpsGuXNu1tUcx186Vobpv3L47oxbBbcZoJj1iQYWu
miI7L8rht9tGhPVi+bmIcYoubBKL74XjoLJvee5+pAEFWV2AX22jCWKQZq2Uv/G1
0ae5vLLI/TrhH7ocBGH5zNZ5/xTJiuKtcEWxrb/bTOYVWWEm8KjXLu4CN3viPeCp
PsXP0pb62uP4KzQVMIlYLBOH45UZ5r9qOCm+iRH+Pwti/sqai13vhlO2lOHA4Bll
bttm2RTzM53m0k4gz4IW9DHoePh0rsn5EatutZBuICXyuVKT0gA2dl+bEpszU8K2
fVMq41ADKiBZr31TQMJ622UifW52QT7Y58xNOz3UTm5mdBrex33kZnOXoTyA1KLg
y3kcP72Dq0KZv6zVMcj2e3kXr56AW/eWCOZrMnbC5p3mlDEeFbN9bYRhmNirPF47
kVpOc0754lteAMIR98cgExLAg/Ztp3kKjReVgDRxEw4L0+TOKXjjgTgnWQl4lu6G
zUxj4mjFncf/1w1LfXVYQEmtdQy5pClPGju3PrcJLRXISpu+LPP3x/xe+nytDi9o
5NfqSUJAmRJgSo7K89U+DM/7JjONdOPE3Wpfewy+qTgTkx5/37yc07DW7K+bMs3/
2TpeTJq5zqYs3YxGjnrBWzGr7lZPZ63dqJq6aaVlPyhllX8EwhMc9Bgz1+EIybQs
nz2cHgAEiaq0xuT2jQX4V0+bmkNdKpM98yN+rgJqHFsKoNEkvoQyVzgbyooNsFoJ
c2sR/mEoYS4FOm+aero12IOz2kOlqWdtcT1eg0AvPT1La+F5IdoQpxyfQk89pde0
OguJ0kpi3TH/KHiBq6K4c4d1F2KE70xrW7v7Zb9y5qAwEFNLQxE0/zLQWOk0mS4L
0tydehqsuYp9JL/4HwdmxyRkJYyVZI/pXsIaItbn+zD2c075wkygdAoPUwS2LMQ2
3E0YcMA9EzlaW6ZbBbDoV5MHJjyAqPP4U4GQY6R7s4RRNgKHIRCgbhDyzpHXfwuf
4wOu8Xd/2bI+FI6Q8P1u/SuouGu0dQu2YZeQnhaNmqg6gSrhKu9qjv31WLDHyQo1
WjjFRbYxyQR3fgt3swSkNjE+VpbJXAiO0sMUAy5Aa6yvLVzSCrdtXN00twbchIoQ
AwUGB4CURsJ8allh5AcdcJ+DQ3ZPYVkk1hx4DUp7kpDPUIbP/ZdxImo7opQrukja
gsqhDCtYWaa0x8mgXX9pQOujoqPMYJpk3ZgfyhWyzxjU/ejW5Tgw2Qb2vfnwviRP
G88wkBtLod5CIiUunHz4nySGz+VRfJjCyokWn/H/j4+gH5s9F/nDrJN9cVyav2a1
Ch/HyPY0KeB9V+K3eTmG8cRBlEyTUE/gKYxotwlzhTlcothpTyB/wBFNZVZQccRM
g6dqP/Ba9l0D1TdNJkWwsFEzsAAEywIJ5TcvBmTUCj3mZQX9+gt/QHlUMgNXr+il
Eo/y5CT3J0+RftuqMPeqEllsX2m8RCSGFM7R1v+MY+Z+bkxjkywO9i3Rh/q++T/V
zIZLVmi9NCIBS0dQnqpFTHqaQmPBeJAA7776LTdMyBW6AKEgZ2ccE60TCIZ+n2fd
CJIfWUNDtxjg9tveOROVuX5mjSm78lEb2A1539VfG+xhopgqA7WLkEifjr59le04
Pq6ORUBxyzBwExLL6WzGjyxjUTnmUGkQrA1SBX7ME0bCEHmM19zTjNOGCYTZUxiy
zru6EQZAb2/a5t8Gz5zbx7GiOwdj7eD9l0H8Ocir4d0B4FcGKO7giIL9WNRiqyJJ
edGPNr1KEAG0pHum9JyHo5OxvHsNy8xhLhog3QdO4mKh+Dh6ljBDH85mJs94z+q7
yuSNTFXnlUH1FalHKYuOjBScItw/hrJogEKwAQET9p/uSThFYHVfErqxOCxs/f+7
/nDPdtAqkFtqEaIxBY7BDERLdnMleeewA4awPRLqaNLKTzpMtqtoIttazECxxkmZ
ip1Bsr1cC4D/pS3dXMqAQwEkAa3kQC4lCSMJc/69WM9eNtzzKQvVlfM4NrIj71nv
SHVo73Q97eBhj/QL5+aYVkO1GI+sF9ueFzFs2RZoZ5Dsg8zYw6viFuzZ/dYSZPkV
l1pXm2XjcPy+VgblwSAhGbKPqDrpbXSdWP4wwrEcPBUzVsVazFxj/altSPC80W+T
qvsRsbs6qD8YkSj6LKQ7zevlGyXCSqsqV/bSfBe8KHjdzqoevQHTxb1uVno2X1hQ
GwHnLJxz+dwnNzwkGNX5lTXU4cHcHcLg2JmSJt6dacPuIOUtskn6Rmt1Fp1KD9bP
vwzWOkXCiEgwzkzec19gtdiI+wpGEqchWT7/x68ngXFW1a2/aEXBDuIA+w2Q5X8A
p2kqdRoMV9KoQoTCWs7WsTEcj2yTx1ZIab30sXVV2mNSyaWmA54QttZxCe2UA8XW
jb3Ojugdx+xOjLlMEJjUWZc3KCNBrxuUGSpW3rkQln6nnkHjiCNI3LtRFlDZD2Gq
L1dsS265pXYvlx2wNDPgilaX6H8CRvxh+YBgOWOWTe415hddeUrJ48i9egS0iIRj
fu91Am2DeHS+OA7KplH6e0H2Vfu7ahi5L5ckx4GwPURWh8T9mW82FswpJ2vAk94D
krHoCIJN0/uuT7kFT6HdcInWt3GL4YCLMbB98ssiwO3qWYp8gBA+Dv6Vg3B5dL3k
GmPisKa8NTnewJa3ZZNKy3Ar+8/FWXHcDUWVpjwvnvO8u+PKnCtRVZz01BTRltsY
ALaZ0HsNDkqRHUXzFrJQTg5vL3GFUozpX3rktr6HQd5OZq0wy+n+HS/sNXQA3v2t
vO7yXAJmsq9swDjGjmSrQveC0t+n+tUmZeK/N3tKqM6PayW6IY1XNyUzQIupkK3G
`protect end_protected