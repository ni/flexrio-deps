`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3328 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1af1Y+Dk6+1SXWNwztYDhwzRq+SJpq/YewTOjrXpJC91J
G+Ihb97h6f1/6JgLWx2OFROPeBmP0Nf8GRlkqjbpS8ZjWIX3RO5tFHhzIJCq6Zhw
sRRvFBL/uBB6s1q15N6LQSKptjemBRrn63iYGWts8gEGesAFiigXJyczPHMmAyL8
WMcAqcC7yrUPclOibBIW7MROIZSq/2/0uRUU7zkLYgJwy+laMV9KYBQC/pO+QEQF
LZyqcUvCuBxniaYieKM0IUFHZ4b/7jdARuS1rimMtHoo+f58JSQLR4Bi9o2w6oZV
A2AThQR+ABXVDDAZ/Eb7h02MfR8nLZUWOnUkltf6+jOff677hXRsbYTdfoZKvhJS
n6kLLbnz+mFvwsL+twIfkup5hCYGdfUyoOc38JrFXzQRLkEktCRI19GSZii8l6GS
89ao51N1N0UGFgGSCTr9MbwZYNGHNA7IJhGixLn7o0pOo+7qzvnRi8ETI/GafqLQ
fTAliTVvY4EIaPKqdsK9iQyqYXiBySK9g1EPfIaU0UOeBivcNbrg0ezwzxZyddGq
orlecqYiEuzayV9To92UIb14RWa2+z9Dst46cLFspXg99QJFkajaNzcRa41Z8e/1
UKK/lqtMirv0ObEdD5sSAjj429aXbquJYU1uUxf9Yyyzzff8jIJ6Bc2iq9qVqz+A
fpPh82IXsNLWl4RucKpnNHYIihpgSnCItWiS+Sge2rUswThnvUMxaIFqRoFA66fC
/qMimEWfz4L3Ucn2AYRkZSikxOfg1eS3FZKuF5uIm7WBAVPmVFMdZlTHgZyftD3A
J539PIdDUgzBFf/hMmzll7RttN/h4v5Wn2OMINas+USNQn2buP15VmcXTLly97VQ
Hb8Gn5snxRj8PNqRHPQdnSCiGdFYlQYIfPW0X6RTRLCRsPlIaWyW7RS7aeX2eU+m
D+zHzC012rszddgrud8+JpyhY7oMhvnal/afTA2L8oX/PlSMfOTFR5KtmMiQ97GW
8q2Z+MOXoNQ6YrkI37IudHdsnXu5V3YCO1vZ7fbJRAc06jSEiAV4eTrsmrCnuvf7
3oPpbtGz8gS7oljGYOsg2SjNuLlEz36o8YVreazpMQwy3JpXe/qDG8ZCRFCo++TU
rmssT7IRE/S2OO/hOUFeN/eH588YZwot10ww2k11tHn7HULh+0kO8/CVioEXLf+B
0TmnvthJxH1GmnGSlDgZ1bWrtEmgjUGGCh0Xl1byEnThwfkZHZykb/+DLnLj5Tdq
UYJi2zjCyFkHSyvN9RuLlb+ozHBfbJGwvbNqNGle7mYwqK0qEpnJyh4KQc35c6G1
GE1SurizKk3fh4bzo7OsA4bjKGKn73AyGhtlhlNpH+udPUcuvZWwRDqqV3tIbkvA
hhnggtAGZKaQjTXdIHMlVRFv6QqqMRdpI6yIDXZ8kgxKaNPRgiaxlfVPqKks1Mbb
gNnnemOul07GHaZdN2AZFCkNv0+gj5uETwLVjxSKLXlOUGD42wcMDttMfRN7VkqS
S3Rz4njKOrvXyxpW4kK9GiYwDO/tkJgiyRFuo0hN6djEUDumbsx75KTdPjrKT1Kx
V431sA0H4DLFz1b7LX94ZKzXmbsI5JiFcDARdaExg4/5WGs+i8fTZO5LA3SRBkWs
owP6Pypiv1Cofgazb+0I7e2wvyniHfBqBjBX/4V4RGyYQlyC0sXA2hY0FedGi3i8
Y/loO6cNLC4Bb+/koPwWvI65v092nt0qD+cC2js0iifDPU/YXVYVlKp2GEkN4Wz3
9QLYlxgtT/UjhWTEgo8UZ4VIBMIYRT2t5GgoJhFUixYDr8Q7K7ORdR2vdKXPpV0B
wKb87c6E4kHhh/1G2Rl2XPgDqYmuOzg5UfE9ZBOIn1deFGNyWqepLqXV0nhOsfNl
z1axzpvnaIuyRH8n8iHj/WDZrFKm1uwiVV2MjKL2swXck0gAzs0m4kk80v7TWQq4
RmO2tKIZjbugqvIFBE7G1OssLmfPCeaeTmI4OG//th9RV5cbVjcvsBkIpK7oV3ai
CZwS4B6AVCGkjxGbWfsdMZ1jxdASe76iNd0lmmj7dDM1NAer6ZSWpLhkVt0xJsGG
CNsIpIHn8Pv5ld3hCV7HDITcR2mMOJaIpr5UlMZ6Il8vaApvT1bwsXF1xDhkOJz2
ELGYj8/NRh93QMRogfdzmTygTChVSrdXN3VA8i37nE6sCvM92wUFfOYW1EGY6bQH
2CQCKR4N1Jx66/ZBSnm1Wnv+AelOpdlBjpS6RKqwP114o6/9SPsveIfNs0ww6X39
ncxJIwUZvX7S/WFbf7uPR85Cz8vkDWiZ7KDWQxhNqgghSdtkiz3seQEPWbNf6kgO
3okYcpg4cREcSfJ4++kc4hbYEsgvgEktW1wbFCEQY1Wz3hTHGw1myJFF51TU2xhd
Va032YdLSEEP6emWcpYkJQc25BzyVZDULDW+TgRBgDaZWPFD1XsHq44cT3QPdqjq
+Ru5CoO4F5yVwmolKXACkwM7YB/6JRWgJi5MESmw11VE81ra1Pw6jWo0cP+6faE4
ctW9EF4V9W8kIrVxr5i78sogOmj8xXGws0Ymxvei0iooQflG282y3ErP5npvLYqq
vEgXiTIcn47OWyjr3/RTcFyjGBWSQakopG6uZuNlQpByY5TJIGxCIefN+pkcLz4h
uBTWTm9LKbXQADt9pWqPxjHyl3yObrUg19B7e7uoa+eOjOYl+cjZtuG+//O2AjJ9
Oz2WCWtM0JRWDjZ3tDiuD719LIMigiUxlLb6avzWMrk0G1Ym11dCDLAK1hJEr9tW
pKJoDQcLYYIQ/TpGQDJVBsNlgCAz6/JfSL11cwwv7GG6bZ139nZ3GorLNJwRzA5Y
YInRPXMzGzLgXDOJ1CiKzVBqWznn3luOTK5C1hq5oo5rh0RGnh2Q9dwrFGgt6Wvg
OpFNVzQVUjQ/YoMXjR4Kz+LjMKEbOLmdsmLfbXjIM/OP2G1fE83gQXwodY5tLvZX
Mm8qzjfjci17MmkWI146AKO6qV2AWe2z8G4Opi9eZsOZRkycGSDy1NnCPaG4VF4e
faMNUHEqf/7L1al0xopUZAfS3kNp+RT7XuyH+pCmcC0skLNzFbTIjR/d7QVypStq
xPdRbZVJrlNzBVNbLoB/pN09YVpeLIVWNSc8csWsu7MsrMIJolxM1Q/GMgXRP152
dawBA14hevatr+1MXKl2737E1znePHFAEZK108bRNABkHga0zg3aeofTccATKDzP
9kTWbkwAhJYSZWpWnJoY7oHdY3XQebfhPG5WUtVueBjF02d/3pIl8WEGlDXegtrV
yqtzjd94rXQE1eWAQ78oQXv04mGp+du2VV4GwiBwVAtz8T3I3l6v+lwPGe8zj5Va
xDKW5q7+zqHF2IeGG5zbSalsiGEgaUyaxii6Ik+rdrjdJyRqXQPNTYmo9MVYGxe2
5VbRS8VJAS2jYHhePS67szWQPf2sS7zKf8soXElCtgEqDFan9/vQ3WDm3MODU+Fo
1ydloh01u/zH2cf/Le8NmzqfDCzPmjJSsWxWo4/ripa8Q0/bTY4pMLVRsCD2qXCv
6TQdtWIOePpE/+Esb0PorzQhB+lp1L6jk96tEev/oZirKM3jySn+RXk3xcveAsaf
2Anqxnye9xlGkjVxqJNARQkIf/MogmmLM7CyUmhSwrgtJFlafWL2D8FfEKjzL25B
tLbIfRCdidizZX9dPro1nSwV/ZZ0n9DBs8zQdPsbuUlj8U14Xl7ydP0MrTCCzDIs
jqGxhTko2aXONWKL9ysWoJCCDnE/p5xosya/tl404RVvITMJrLICXUJybhhyXlnN
J6S9zZr6OE1T6C+FPcb5hQaEpbn09em2SlEduuZ8XwJtYY5Y8pz4VGQpmwHMaL8w
ehXtULBJevKJje9nYsIFf4qjMOmriAtLbiSz6MK7WaB7a+v/1K+j2476552WdU/g
6mp4avlZDc8sdWh3MUfda7YsW1Oamg4+0Fk9fajQRjTz1NDuf23RzevMvlztIMmP
Tm/DMYJRNxi9V1R8BhSE4yXWLIkZSjdo5bs+M8YzSqt5W/bMbWHSadyqhFE5kz4H
HCpFriACyaYCqUMOUmXj4VyNc+LffbZsUXm5Azm+x6WTzJ4vLaLTUfWxTmOF/jc9
xkLn0S6zp9yV3u8u80OhfjZCHskugJAA2HliS0S5+8B4mbZZ7PZelaypoA0FbfAq
2Z4/5BzjafGYyrnHA1uug/sm4Y2j3lGNuRPx6aTIgqdr0vCQop1xObcp9SJ2Q0yB
HdHFnKOtG28sYEesOsA4lA==
`protect end_protected