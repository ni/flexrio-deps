`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3328 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
akBpHK9XojjdOyFTP3pOwjvYMTZ1Pr+A6pQ6YF+ri0YteKEjUJfAgwAi9wRp/JTA
hhzf2i9eCHYPOEcOeQtJAQ9pSXHF87EslvNoRqmIzauR7+onuwSNayd9yGQAe/Hn
Ao0cfjD8pr1+REjCNKqHTDWew9phRcLs9oN5lj0l+bCjH7/0zxcfpx6bV0C4pOqt
aoJLH4p5Nl72te3YoBd4z3xEUUvUdG5MekBWfXo5fWc5aE2GbuWXQjP2MhyibnIE
cFYPekb1nJlObWd8NMBZAWpCoL2AZoxAk0SGp3eeF7IdONe8DGt+dl6lSgchojUj
FuI//Gk5nknpfByBtBzIVI0NjseNsVHtm0BRlt5EWwb3M6ruYq7fgV4u27JmqVNW
7WwKdSq5kC/UYncSwqx1L1c0qBQT2eDpUpEcGUjuwvQ+VsmhKkOhUQxoQITBLX2b
DKLS/gi+wiNAwiVFL//Df2uTgRh1OSCFGtOJxLsgxVWLcFFQJ5cFxK45GMVrhfqO
kR/eMCUQNRtBQjX/mdOXRUWISAdPCUvWh/9NIQv4VmaIUM+mV9KFpZew5rp+Wl/y
hRd9JKgErHd27FjTveFBIGX+rp9KNP5TAeQgEQCh+fx2v5XOs676NdMs6SCRyuvY
Vpif/jtvpUxyZJWNIV88h9369Iq8mq+RrKRv10oZTKbguzYwhY+p0G3yCvQxVZtX
EWYZGn/mmfb08OW98ptG/92F/kksq1xn17G5rhXaHONh80JFzomYiXUmQLyWmMjT
Q84z6s92CQ0XNQQ7Oq3rUR4VQZurZCPLRbtV0TbPa+lbDD2V78JlwOzXkc5xcEik
qvt8knxsqJvG8LNtC1xWBqNCvoWCkgYb5em/BshWlZ3DjGEhmbqZfbunRlFHiSao
1N9pA3+jmZtNzZuttuQ0CCGWdKIjXHx9XzAmaGmFKJDozq4ZjQ88EwoRZHY/Iyn0
9zXdLEp3Xmvb9t4AKciB/EboPNdXa9RQAJY7qMkXL1RviP1cEOqWwfnW+D9gHA2p
vKUmGPBbbX/vu+u7XTyyhfk6IVpiUIwBt5DRw+T8gg9bHEcndF2PVqeUGjJy2pQT
3gtpM8ZJeCtFmjUSEmJzT0ooZqilq7Q7T6YRLcVyvVY8FBE3I7nnwozurCjQyCRe
fGrpKRMn5wwPO7cvHYodXkj4EdwnkiRT/fHPDtndcBkDf21kuUz2igzrS+aXQpNJ
qiwbnl3fq1vqF4pI7oa28QUwkcGPDWpj9yDNtCiKjhYOlpUIYuDJI2bpeBfvePYA
0XTW8nv9txRpy4VOzyhjaoggv7koVpp/ZrKNSpYFrfINaSBfKywlZLPjZUDiHNYy
p8SHwGYrsGJ9GBgbtl3+oMlaEAhJvvoXcIDRgAZNC/CDYZbep4b3HPpgxqo1AZZc
mPbwlenp+rJAmfY4Y6pYYVYVt38b9JZXPPJM97My/fciYMOwc/NqzUVmwSAoZ/n6
7+oSf5RrcDVvBAuZ4lxh2CGO7Xc2N1hy8w/r07pg4vUiSxPSW6DZB1+lJGgKMpjv
rc4SlQ3ASSCK43RNjzMEO5HSI4l5uJ5g4fsqTtklVbkoHgZlv7LJdau+OVYzwC49
qz24YnoehX86KxS/zokj0wogNj1pJAa1pkCUUBPqoX0mJH0KzioeQLwcHXqGiH4p
GAK247v+FhuobxOPvODKtXP2ya0LN+Z7FpHG3V69qTnjNWWHlo+OqnE5LE1mYeC2
4XDt62RY7PrApea2L/q8BHG1dL8f8eXRncGnyr8y9V7Kw5SQ72ea3kBPJDKSs+L2
hJsj+PK4NrWZvzT6SC4CFDnkKe54xGOzt/5bxaI/U0n6ZVeZL+iODtWlQftllp2Q
/s9BZcmhAXVD1sn/3VAv8omXzwh3Sj42EkYtI9PBoAP3C5O5f1XKCEnvL7BZisL7
7oVa6Qp0oUYQOJlgqF8eukS7IQQGrdrkUtFu8fVzSeNN5cvvldCZEv/80TisQa5h
OsNLib+VBDndj04Pz1eLeUYxIRm3EIzhUbGS56ZG4jiMmeUGm9diLVqEmwGHSzOy
FKXvmhnWLASY1NQPJhV/YNT0xHcsvZpeg7fb9A9+f5m+g2pjF/Sh4HwxwoUTWltj
UUe4lAjz0Yp+sheMKYtMc6ygRgORvqmsRs8GKTuwbdL0cCgAP6u/lkXkgIsay/dC
Ax1YgczgYicciTtDf8WIPNi4CJdbx/SnsuyCHEe6UHmpJP49qB3GHVsov9RbJStY
bY5DHJD80JdDwXhtfrc+syg5B+/PVTN5zc2sXEPuW+1/62Roa+X0OfEJhW1kdTYI
PxcyJufZJACRmrLMWcpLa/c8+4riskoaoOuhzglqjOjUB3ro55n/pku4jgsiwBPF
q7KtNsl4OwNA9H5Mfi4GPKvfAAPL53weLOCl2U3MTCUR9vhxclBo4+fMprrKW8fZ
dYmkz0bVg0uD/FG04Um5yzR5QZ/AIi0E57geCYY9dbnaTbi+frAmSZ5eGpmLZEWp
kM64+aZ/dby5wXc+akcJtzDX7aCieZZDIjF2lsuzekQLcup39AdK5OEdJgg62RIg
FcOeQWRCekusGK7hht9vhyBrf4QrSjCu2aGG5bfsDnpYuczwb/TmWUJx5NewNcFv
Z8GmEWElZFgiXEdI3OScDlo/K8ycp3JoHlB3dlbItck8dQvrDJ5qNSFWqz/HMAOv
KTosxHqO+VE10tyg0KcgERpSknNoxijmgQUuRsc9a67MA82DdgNib9Qn0tBgcvDI
KVjz77SNDdOS1zZ1HN+aLN+g+lIruWvZ757bQRVCsav75z/GIskpXJP67iIaGkGy
TM9JSY6yCpqbdeQnOkjfR8FOiRTvaaFUtPA1nZHT1phdE5JcVQVOZvTSluimLZo4
fyf5mwQICgLR5nKP5mlUHpPmgHA1o5CLwiaLp7wPdowUCeTrzYciOQQ+rM2QZ7Zo
FfHvz/JLlaHAs+59lXfTs9Tr4BXG62bAwEzNKdXz3bCJ03Wwr2O6X10LviD8gR+d
2dVAWED4pl0QdYj3nmhN9gtaxlFICYyNOT1k8b1OD/oaEFlkoNL2emhoyTV3e1Ec
w3ZmjbJ95czdpB/Wth22lr4eMxIMD2PPV38ZYg+4MlN9X27STnzso6szqpD/7SWE
uw+q374n+FbcRr/fNwDa1qbrA8qTEYo6oLq2m9TuaQzY+xhEEoua5Qc1+MESXn09
oQgWO9hRDuxYfXP7s3usLh/avonKjOVsdRtsOG96NR9uS8SWlVFS+pIvEKLDRxud
wa9iNT2sIyR7OXkajwYt0rX/qMr6ER47wnf4CtvlOYlZQg5PZ6kjjmi8mopJm7Gn
r2L7i5Vd0Li8Ahkp3i+oVi1B/5CEeXza55ynIAp9uMNCVlseuuOEo3k6m3pc39SY
wEshzrSJ7EyzFeh2mcqkhvr14bUZX8SLFwyp2Cs2GpBxp3lCj/3i25tBWXRNK3lp
NF8IedTwS+pnxTUKQAC9wyDtJawRX7V3tgdO5T0alAC1yoBUzyqnnbnqL/MMmssP
hSxZVpZ0fjm+2HPkYMczd+a8nvuW8WwRrIEsIJ5y5gI/uf0+yKybYk9hTlarasma
/0F6ZZCj7Ks9nEgxsLrS3qrq6AsYYADC4wMeAglsiP+aqmPb2t8IdmilLLfdcJoH
xcYy+3xjpCGv3Q9EqF3vUK8snsPK1egahry9EgKswLnqRcCWsqIk2XYvqcTkC02Z
uOvof4SpA4IC+e5Wm75jX4bj/+W/I2Zb+CH923gxyNic9GwARLAWfbS3JQzOBRrx
F02euzIIbFcBIfSIoMPAtoyZIcP0cNJ0WhgzYbMhzGZKIi+v0Fp6pgIe58CFLkfP
M8AHfbHRJXMxfei7Q8PU6yXYVrjHlRnmVxXwPFNrydWGgWrUaCuyHNHeztzYj43W
FIg6cq1Da/Ygcjxn6HEmESkX196Dfb3nFreHEN3NJ4uk5kTCyEkHpl1mhOeiN1be
R/stYGTZ1bCOOlbYu3QEZcqfmiqQkWKCB077zOh2J+9EqiUkoVi4wzqSpNxM+Kv4
qXOCSfkD7ctR+YcpXvarNCI4IHgtG0o0gX4RJyn3G6aXhvpnmmI0LGnBDZeSApkC
ePQc65EeGyT3SWM2Icw7xK/pFgMAomiXqaLTlOHN+9Pb7YwPp92uZisl1751cgxB
tYHDFsfzp3E024qzR0GSA+yPPTnNC6Q30C4zCAgN7FCP7wCekLQz/KpD7xjOBxww
yWslnlq2vgMrSKWZroerrAUQZWqSudCNo/Aoc73fzZ18KYAQQkKY8S7Flva/9OHI
35hy97gCEGznHBqXa3sfPA==
`protect end_protected