`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
j9eMmSPGcKCWAR9PvkqZ1R001FU8QKTyJzFqNLn+qur6INyYDE1AI8LWcxAzfnTc
IpZG7ua3uuk5/kQKKQx8ZIPLfmv6H3t3eWjki8YIAtY/d5E7Gq8Z5mNxMYRzGGTg
TCMm6oOrOTVYlCXHE0X9AW696Z7UGfWirVibl8hs19hrFdeZKGiGht4r09vHR+Gl
FQQmSObM5aSK5wu5KOrK5ZUKGHyBhjnIQO5NnittDjOwxV/57nHVg0pdG6JUqyvm
tEgmCY36RCMRGWN7sekPtNHjqpZkmYrVX1T9QF3h73+8ZekZYd2xY2hpHHGYYeWA
t3+Fmb/6NUmoP8+Pt2hI6g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="wX+NBVcG/A5ruHK3pkDqG8ZVPdOz9TJPJ5saXZYSeQ4="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
j/hqWUoxjK88VtH4QmjIrexFOSwtsLKOZ/LCP4cmrqgzmR/e71apdtoL+o8nlfy6
eZxDZMmrZmJGoazz2oK6kz7xJU85UCwNc4cxAsVxNdCP19vZxph/nCYZQ9lUFkLH
uLBkOeFP15CD3jG5/dp945fHP13J9SzB/L9PWvDC/gY=
`protect rights_digest_method = "sha256"
`protect end_toolblock="sqDZkaglKf+bDjC7VKm3lOELrT2Jlynh4UhPg2J0Q70="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36368 )
`protect data_block
f9kZDbPp4NLiAOFOgATj9W35i3s4a7wbt9jeHjHVcJxMoXY8rb8laqS5bNUhXGW/
MOc7UNc1VwolqhkS7G27SLamkGClZZtXSbRcN1N+5kZpEaBEj1343vVznnU2Dre/
bKlbmouB09/BfSaq9uUVg7KYG6PFzT/GxXdVAtdnNfIGjvCIgEKEZephnmb/dClH
A/d0mYwuZmt9rrjFeTN65OTniw3vqa8egPLjIxNIOepAiTfo56ACgAsjVqhQGrOl
zlDj9R6t06ySYPHw+36BlUR3wIZ+IfjqOW4zt3rpC3SHCjHiRhbMoxWRr+/Za5Yy
X5w0Jrh2b6ppfhodC6tUAOSrQRQSNXpuHTqAnWc9zbJPMb2e1l7tVxIXPTA9OYV4
3Nst36OsYhUKU7MxWhQ1zlb0Z+wgCZqvxuGk3mGmtvlE/Ay5ez00fNNZFlp0ZHnj
S3NSFU+8SFh7/HRT27rsMy9cWhYqpbax5uqe8eeLGACPWrxUpoIyh1CRVlerIiHd
Ydf548QyY6mai+2H8Y5bmPMOQIwnPK1rNchofPrsimWeB/kkcXyf4fpBoeIvqzhf
RwYp9wkXjuU6Uj65pDVkSmwM/qlrxne8i4tbyN5SDPfihxNU4yR1G71kXnqsFgez
6WHJM89+89/ETC5aO3Ba6kWz/eqkzUJzN5ySW7imNX8j+iYPdvW9Y7oUJJSZ9Oor
+Jqj+x45HzGkAb1xykrnMukJElmAU4cMSK9V3St13jSjzFkuad85JQYlEZBnLUoP
CAORzWLIXOTsA9LF5OsCgu415CU6Wq6RE+AmtkdkRjX/iLpRGQUnJlfjNVDMYXpr
4mr3AOaRvSTZ/5SKD9rJ8c7JB+yo+7IdAgZMCTZyk/7Z2MWEjfeWkZUq0hQAVwRs
om1/hxLqUAPLT9pTJDLbQmG/NLBgMWF+EH+BDwLILyjuCmLQRT4GPMhg5pn7EoTs
wbioDOSLcA+KQYtyiJ4s/dqqsmsh4g9UerlkIKn4JUBNT7n2/17ExA50OcZ8FM7D
8l8ynkCzSC7GVRa5A4woY7GNPBKCN7dPzA5jxTTqFyaz1QAOUaK25jCucmC/HBkm
5QE3vCi6BvQpiFyOfjjQkU/Gj4ScRhV4WKYs1hsaKA2O1k/nGz0d1oJ+azVaiwWw
E/jlvXvWdjRKCC9kkQCJG3kS3H5QKExIN435d8b+BWaXIZhvq/kxrvukK2ZOUQLs
bUGZoroLTbaun8EAYOvb5eJ6aJqH1zxNNpqMDTLKnf3rozbypcVoXK2WzIpCDoX4
o38sCy5YdGK05+0n8UaWUo+Np018xtfl//ox52hA9MOZaUDLQLuDFLJd3UfQ/q8X
Su40Yzn+OvWSzRgoPRQvs/K/LD1ObU1hwieLauadm8Thwt5r6Xc7eGGqlkCOUiZL
xYE5dP4VeokKecXlUIVtqa5fy+Cp8pf0GMBjRRJRQuXlLCVv4crMVhmMozoqENpX
mWYRV+kXDBZ3bM11xgQ8rqq0IcenumejkRmtFh8SPkT23VUU66fvH2+HVPOWoYAe
QIzM/i52CD136MbKnMmfa93PwStYz0WFxdVmOD/1iIBP7NZ4h9SkJAusdaIFRnGO
A75PqqDEYpfLA8WIJt09P6YdmIebC2H1rI3rN+ZvDhjciC2Ym80Br2qnnr98c0DZ
hPEiHkEhxqbzVrC2AMbfzeVSVMHBxsZ0B4faFjxGCwVPtuNU5b96LA9qjmqiJw1X
js9cSVOOsid0AxAlyjSfIzmQPQs6nq8p3eRnqRYqljXMoMik+r0Jhfjin8NMiFL6
iWldgv5vXPbMJYdTXurr9xU4ZnwYCTrVM9/SO0yA85nQbIh1g5ciIu/RnCOXGd84
G4F5dL5CgiyOEkpX5CvW1arDogurJFkLyqv1xT1AyoeiKO/QhYULNGQNQN4ZdlaI
FhwFvr+n3aAkgiI9dX+4iC/GDSJHyoddrKqdwAStjEudTu9uVXh65Lok5u5RWNKK
SoD4IztFQ1oam91JSg+o4xJvVOt9o1pOPL2obJbS38TN8KLCuhkxAPJF8oOEOPJc
zQ1/OtB5OT/vWoT+qIfmRCIg/S0ErERLT3ClpTWiS05TAthhSH+2vxbiiQ6zxMbt
9Y4fVziKlV0yfT+ZCBKh5Ml7hNgCxm2dfUr+G+WnoBBTVC5K56bztI1bBnSA7Gs8
1F1sh7dsVvHoV0Sv7eQUSvKqIXXGOIzZrEbD7Tg/UzGjzTM80bpzDSS0AeNTC7gc
Ewm5e1TPa3MMOtWkXU//aL15/jRRMNpwYK3/vB18nv8g0UWXh2ongcWgwu1AvvjL
7xCuqquOTbY6aUbUYyov+4GyvjzpXyAOPFXlarwKx2zJvZ4yqC+mBSf39aatQP+z
UDFanzBr0EPczNXLLGrH5ZU1l7vcufKRuAqKImK0xhIjDIdu0VMtkDL/4qku89IV
YlVcCk/DaPqWAEksGusKLMku0dG8i6AGxgDyd9AAapG7nWulyzHqcghP7h43DJyO
lbeRn0gLNRYQrPPIUkw8PZAdJ1ywmohGK1LFPHWwodXmGxpyJ0VHdH+rXMU4OAMe
TMdb+YMnhGZ9eYeML4m/rl+bD/p2YiDQ838jc3D5/Xqc24bvfj5iRR3t69fk05w9
5niniN7cKMDk7KSpVfpKH2oVDnrhMF1F7s5sTGPkxNTSiCLdc4/J6Ei6QmeNxO9s
lAQtaUlGfrcOkc9ozfDep/c5BKAXimWnkK8fsjpbiD3EgPxmPnEk6eTMkZhUuXpV
TPuIWUn5wQTCXPw/m42daGW5HCxhEjmoPTgV6wMk7n+yhA7uEScpTEP+bAFTBa1U
lW2Y6Xae3l/HXqOrSKTnnJQwb+r/alIZLSYEFZ5j9p6cR0oioaK0u4QPg8iebRTa
m2UdVwUQXWjuR3NpZzNu1J9jLWsg/eKKzADeGASv/s0g0lA0+gqjXONGAJI2/pVo
tFw2sGErtGOSvKM3K2Yo4aM96zlHl7R2ybGfNbOIbgOhp6otaqKXumzsyEqe2e9U
SHgsH8Q14KyuOe4oiqau+LjrfrDCphpWYUz3V0yeQwrH5xrwQK7HoZW45KRHUZHx
qpN3V8sXTKp+mFLTpnjzfzSkCzsN4LdCNlWhRLAaAGvXzUmAbqop2pB8VC05MEVp
vDGkjrXe9uwsyIFkEneCEJz2k3eLKjSgT+Szj/AKG2Gkp4/EhzblN0LRfom0tVGM
S/VdrT/tupDPcqb/H42Y3OxBzXZxleM3m/Osp7B8C15P+9jyRyc8nmGCQjTq3S5z
xitrX23wKmAZMu9GYhjN9ySoj16++bfR5rSXW3WdLksVu4jYfyEimFPtt0sNfTzL
mEHbEmMRHkqKktRVDH3oF+Iepx4KP9PuHajG1MkluZAItZw8t7NZbLbdkKG9fFvj
72R6cTCwt5dg9rDQg4xRFyh+vYwP4jL6gvR8sMiQCsuchjwDnvn27dmu/ELOQq9x
zCyPh6h7rpLwzI6TTuRmSF587Pnvmtp+vVuSadTe9SnKW6YDNhqMQtOumFsLaVKv
E6lSt35+6oa3GXnDGTKBEh0pGZFjBXjV15+7i6AYr/6cpvPATnoojqZafo2PBvkx
cBeaSWAAeeHSfmr51TE0cJztA1zLpJxQxcPfZLqGnKZ1OJtAKH7VvNSZBEjPGR+i
z47BJ/AQP5k6e0C8Z9CGIv5QitkCaf1Nu1f2QvfMYPMYHNy4EgFG+wc8sb3qfKap
PyrXhaTNoX1qKZcbifHhzLXKRivJQTjJjtUMSl3w7f9/xlZl+VPtGhNEK6JRgLhE
g3XwQ75JzzvFtUrMOXxxU3LjtbfzY++K3gKI9/EGHqcmm07MFBbPwfXxxuycD6tR
HK2JTRPRwicE+LpygJXoYKL7E5zETxx/JVdT4tO23UAsFzfMr0qqOaSl1VLptjqd
Qijnnra3qdzaq67Q6a52dcwhhia1qf5Hx74/sj8B7NPeBlX8sSkE5N9NoJ7QPpPv
G48CLnwlA55Tm5XEoxR3P/53BGhcBVoc8MBalfr9CLg7YKD05KmCoSXmo3LWPOWd
wQ2lr+hLg4IxtTM7VIDEkaWIHkC057fZOKSkrsMJ4k2FDscnIFa0HMRXW/AvjkAH
ilY26HQvWMSTMNzs4csb4QVTQz27GmmhyWe/alx9AOWXThfATlQHyNtu6r5S1gCx
9rM2a+g8O0V5bh/lJvzt6DtPqKSqABlXVYYpXPdg3Jua3FWERdsyxsNvwfLzuKMj
LowYQC8Lg1fsO0iPvgvgbUd9n6D6ABVon3droMVEJKQ89VCxM6Ra0poRsylOByQX
YB6ZZizYD8Cjbebu2QRLigzt3cFxTUeMowCaUNoJCCCZFjPttQ4IlSB66nVFmpV8
AnUjQ1cccb9DH25/UuzAClrfMZayUpjHzcr8gABptlDfw1UaeREFqI9yvLQ43ykC
jo6yxly1TlkwkGME/TadpvrDTrr1Kepx/c9NL6ZRKHsQYurCs6hNzcWUKD5zpaeq
2UskuRrXUgFXM/SpPVxl0TW67awbe2JHLuhXou3fomWp8ZmsDEfDULsizgslBkjX
9QhL7diW2IBfKxqtZCEgvH0g166Bt/rsr7whk9GYhvHLrESDVPPaddZX4i0X+SEU
iornPNDOEZ9qzVuEO5kQu23in+iNOQzNLres3F5fxLpAf8dTeCWBrQ0KUl9bb2gq
s8XRagPel1w9MlkkmYJVlDH+PzzvB4UFwzlBZVny2AaKsQD1FZoXBUIfIlZ6JJnf
K+Cu72XXogLgm5FyNFd1/8c/v3HmGKokA9gYEPQ6e/YHqIIKoiZ+l5zGKthBWHHA
wQknVp1d5rnSqtpX0qMLs2EQcGNqKo3wIynVIDQvVTrZ5A8Zq+4AZr/Kk4+JlP9H
CVRX9jya9GbQhQEGyDvsC2siSFOMRl4/+ao359uExCWXt2f3WzjOQsTQ0iJk9mht
kIoMwu3vgxPYZI/5hDfgdDCe8It7Q4sJYTYBsC32LsaGm6HHkF9BehK+NiU4NfFk
Rxwxg5Ds+E7DZyrOt/HEM6udekjpmaJsu0z28dvhR4mlkkCo/uNPcU0qZe1N7q0c
UaicToRhBxQcvEnws1+us+FRm64SSeZLR+k9x59FJ/XOiS7/EU2lAVu2fV0CjPfq
OQ/y4dP3Ula/GTGcHp++Bk7TtdvQeQr6ZsddV9HSjORTRRJIX2j2/lq6Pw9bJaih
tJMHS4N7FmFoDiZd8m+KD3Ax3S81Y1WDQJqBHr197k8rZXcBsQPtYExCGk9kGdEr
KwHjYEl2+xNYJZnUMZ6CcQMeiRt5MQga9DrzBO8B0yuUfJkSeaq+Yza+2UZAFxN1
fh8cWsmCwTuRBmCfdUssL1eoHEvZpfkabus/JvmeXbdDLGrPvBJ0uMV2FJI9Mast
Sh3fpF10rVDcIRupd1rt+mQjTrKzD0yyoMTp5e4XVcUU9DoUgZws5dt3ESRpMEpE
KBx+CZEjJhc1WtvVzo9MfCRm/wq3bvYgVs+lBgsnVOzf2EKeF1VP28bALG3rvh7W
MmIrkQ3iWGA6l2nNcM8+0WWbXhE+Q/kw9LDiz8xsUFBnIEl/n6cpWyS64ylEcICp
PTyMmMzQXWl8QdcNfbFYJ0cKkphnbMZHKI7hNOgDoFWpVM7fi7TxlxJ1tNt5WQJc
shQ/DYDRhRM/YN1SUNd0iTL+2zyf5ObysaL0aIs0ZeFjiLV0tLArccpx2j7H4Mj0
ptptQWH2/9ca9uPik+fVXTG8h9ZzSbE7EU0ngioSdxXmpHTDM0nQOZeqTLv/hn5q
FPXwEidpXYXssPE/IQ2i7F3VAobfTnky2hoG1766mgPeiZKJpK+9l1lLD0X+dmGt
ifqXeZYy9gNnjO0a0ZmT/4aNXOC0jQ6aHwiZHSAtGOKcklgbVO1kSCTMtC6rejWm
AG0lZ9pIJl5hY8olnprOSO8spMDESmN/WXoILwL/k392coG1OGL0U8CLkwdIpIUX
KfB5Tj5MrDd5Z3JWyGikZrlHPD3uAK5WwIrZFlVmsQlzteh8SLOZfc8dnDxJSD/6
icC55l3XSVUq2nZTmoon0oDRBeGqUI56tfsijlh0LuR4aVLQwWQ3xbTiSo+4tqEG
WfN92Q60++9UVNQEI1juGA8t+a45Sr+1HXFDv2/XpCI/hntMULkS23929VY28G/5
nQrNgvsUxSyRVDylJhYTH3TiuAYE/eFYHcTM1p5dWfVbQqoNmK5ff4tL1NklJUpO
xg9C9yh9i58I3av44MHcylJVN/O07oMAT3vjaRgFtinmkBnk92p5LBvBVDdTGUMP
3eREd+h5obWMNSw3C0bjSYNWcnKFDM304MqvjtIGMlwMJbWA29PWWIgcBMSQZSJz
F6m5ZCyM8BM96Azs1QNTA1NdOIkD+ZcUoV6NY15gfWSzJ3QBS1n8r8Jya8RmgFWR
5QVap2hcR78aloh0zwN0tviVAdyN7ta93R8TlQHqF51z9+1t/TDyOo3N1I7OaUik
9kmlhAT6OIxqFVDXzWyXNZ1kKw5I5vBP63LeZvESyAa0P2GCp4NGoL9H1p/tNBgf
zws6y/0c1mbYwWqrhQFoYuQaKIN3MmGGsDxmkYyn+aj5AZoA9R2zpnhnwd0z2wRI
lhoyinaaJQ7LdSuihxQaYc4d8b7Fo39NqVL5EEWPVo5MMQ5+3cED6ybFjo/3r24R
9g5jEf0f88PMMx0tR5IkFKAh4e8yRGfjwmSAdifuzJuDL5DjFyD6FJ/eaNQmAHju
ZZXtGKo0JiIb+4J9Lesw6yq/rlNigxiwbOxs8AA3N0VxFJwO4p1SHGQUY/2MfzK1
IHYGnjw5Xgb6W8NfCCZsOMG6j2rn9ZC2PvFI/JIQ7zvpIyka94HHUur05GzaisET
lScx61DD24/LHt3rqKRrDI4KaFiw9MHQsEVeJe1O/+CGt8zAoptHTEDPDlfA0LYZ
xUiZmYTIJxR8agGom7t3s7hIaZHYulapuCsl6vNHrszkCt6OUfyYsJfI6OyFe2Hd
hY4CN8xiAJ2U/+M9lvn0CZEY17a6ynJtxEdoyiOXZCWSrp9BxonOcMfAx/Mc/TzP
GXPBHchQqPwmaZMV0WLeYoTnumEQqezOp9+HVXZxpSC70DwsOpzKIReHqdB/eHRB
UlDbQ8YWnANNxGJJx+Hb3CzAHyKCsnSKr44x3F3OKGpVjT+tY75XB63Hq2IT3DmJ
Jg6iOg9+ErmCe8Kc6m4EZz09LdWmzJ0wf21vXHjgiz8Tzt69ljT8+LEM3yEKtsll
ZajikhdS1F0mcSLFZ7WU5iY/IzQGxBHUSCN4tMfa5R4uuoQO7qbd3K50qUYPHE9Z
bAC+rsUtCwN+76kmPEB+bj8OB80jB5vWVaIldhDE+EC7UmGtwc9+z1u7exYnWqb3
OGH7itf9795ZzzEmu1ICpxEfxzOj7QgP5RTXebtsnPWwtc1e9hjRj/RmDiYWtK17
I2gPVoDRNHgHsGbeHfA1DmyOruwk16rtMMmrgLwoYRtDsH+Wc7XxRhNMJhusG93O
EJTeOSsA55CJLeL6KhW+jrTsP2CvAN97ln8OG659nYNZ4fPDdJOWTArJuG+FFwib
GPs2GF8RyULrXbpMU2XCausk2lQooknhWmpanDWmHyDdmMFhCKSFaG8lDbtxLvhQ
7VuKkT/VMB6fZkeF+vYWYiMvIfOpORP3k5IiaY20jyzPPMGJJUMX+s+nrf2p8VZa
EfUumVsgx39VOAL6mqUmg0UMf5uO8pHlGeTvx6L8KFGQD7OZvuYe5amT0dhleeaZ
WjUDZpkjcqNi2eKAJdjyrkxP3blqHfgNSW3sGi2bcSQ8mNzGgzzwW5MY5GSuwuaG
CaLu0RSzPoa9ZBqftZ91XCKJBFjUi7M5Co1oNRMLEejCQxX/cAXpjQjxiBvCDquF
3vBfSWHv3E71ypip7fErlLi45b4sI1C6NCGN1MLS+FfYT74fUxZjDO/MWOJHjD8t
/w1dZZGJLFnPAS0I5DvzkgUcXxDA8TJAXkA9hHxKTNZfX+LAfZZiHwMBOEzSvSc4
i4/ydTdNzNf1uGqA8qp4Q7IKt9fe+X7CtzwlgiWOoFUrWrZifSpWbOEoep2csCbg
e+BSpsa8XZH5YmXiCTFT1zW834jEWdvsrQHQFuUrBLuny4atDj9GfxKu7AoEFxYB
Y04JRiF1Eo34AAeYsDvnytKsTEUDsat01vfnCbWzoiWCJbF3NE/r+gcha2FM5P/Y
tc8nSZZpg9rkoewQGFM9Fpe/Dr+r9bm0YB8BaaLPtCeAaGeyOVPoLC5ay2hZ+a3U
gEov+tQqMCTvTPw6vt5FZwwkGc7K3nhZFfeVw4v2qxH5VzdsB8nfxfvqZQOCngbG
YIGJa6j5wZv2JdxJryToJ47TGQviZxqAUbRt9palob2DLUV2soQTruMa2CPPntGL
JzEpaiLlY2H31grQcpneVQ+lj1UjownkLZMwYUWMCew7gudBj8G/xlPuMnLg6XpI
JfANzu4lJREvWtT57Z5Gsse2IGUOMKeMr0SRQng4DFPL/GuvxYOQ4ykUqzwhgFQR
syzOdTTcr4HWcKFSX5w91Mghkem7lXfNJmQrdWQMbrqboDMCpRRtx2EXERYFLjft
h4AqTxweKAHBbG28VsWSjEPukFE9ZhQsp1INHxXaQx3lOSSwZm9Rm/jEsgLeBbSz
n238Z//Uq/lPI/qif1Fdl5okST/i9+NJW5C/SOGfkv+AGTjk64FO4c/1hX7guiIm
pL2IduRo+WAQrvuYTs8SgAeiuuhJJTHzMEKuEFe3lr5QcqHqsRTasQ0U88jueNil
P84ce1pTtAUtV5yBszm/fO/e8EjcCKbvnYkyqoRhTUabHsA7rPgODyoSjSaidEGL
CR7747M8pFc37UR5aRu5Fl7z+W1PnPI94RVGiZGRjQ+zOlPY0KTK+5bxYI4kUcsl
p+a2bVDonNtNPuqaMRwjUNIcYbh1Fnce7zOc5hMEfnKanEMzijZWEpQsbqXRacPY
46mnCSvKNNJEGnmFYsR/bq968+wqL1TADn1Vf5JPax5gMYGhXKjrhfE1beWEtFct
ec6GrUyd8Gn0UCqFJey3vi0n5mri7MmhNkFMCqHB0Dxq5gcdG9ReXtYOcXsI8yqE
+OLouEwecCxAeEKUor6lwueOxkobebSBotWDUCEYzUt9K5QzhJLzj44BEnhqRW5H
SHEcwaF4z6R493SeNhFwC/xjf8pGmwMhOqK5XDURexqwB80VQr9XYr/y6kUhSeeZ
yyf4oZ5U3Mb5hM7RIeBzVB/7cCSruk9kGv+h7UhxCtGlUC0SbHrkxmzViRSnBiWU
CifSPzWxWidgm2tb6SsYJp96xvGVzEdsp2AdePAYm0/MITEjbdK3seCKI5mjGJZI
hxBWGMzCMAP3+soBGR3Oe0P1vp3/yvrWWsDXmFeR32QSOhUCC05Z/gqalGSEt2MZ
hScDcDdsRD5lr+Soo41MqBd48qAtC7AAqg7UmGGA/iHMMwOcUe+MmeBt83bcqb0/
7vBB+Pkzy4IRtheImicxCIdq3C1ISC6hHaa4sYYZhX9JdOOq/WtLog64T9rHRykR
ZBS5/cE3APA/DUgw3l+8UB3ig14jWv6McVIjwbM3wghttKECEw48OqJlbgLMoDhV
g4f5guoVPGce1YdcAi5cCt1246j2bMOS/a7Ee9NtyKFXFLOu015j+XdYqBlKOHxU
/F3R1WC9v748s4bvDpsBtD5/RAACBZrcj7KlYCQhqAG2bcTjbKJKrEdnnkjVrZku
tA3IeAQmR1GIduoUTJ5pfOuf+fnSos5lZgaNgVczQCNvuVAX/zD4KkrbHEXfWvo7
zsMUxUqG/xmiB8/CaykGrTa5oIRHYHyOZXnHBA9O78cO43V37XV7btZ1pkxfc5Up
Omgt/+l6WY+6A/Y79EG3zonxSlAe/2XAqyoaiLsPW/h6PlObTXgzqBIXfDg5LGgT
LSVJfkpdf4Ux6CSOeESRhxe8uFGOkPSDtL2mRRwcscvOnyS4yHyUA6UdXMuftQtj
Knn3wLtcHT+CMpo9fndq5dhd6dplLVaKW3uiYglesF360i+dqtEocHDbzrAPwJ4i
5Zft02qLvNj4sddIPdb85jLc1YrYPCFlSNbs28ZAh4y0BzPQQKR1RwoeQzEw3uid
2HiLuOa/4BylvAAFQ+wKL+h/8pQ4b8DQl5RnwBUD0A3cXbZUdZVGAuOQbRUC3F+X
fhMPCQi3hszCJz8kN6ITNDsxX3itlA401PaXX8Z6OjtR4JlX8quBkhGw+gdBvF85
Ydayd5ABrVo9w3z9KfkXGnchN2z54VqBDYY0sfh6vszXGtHLg+KUqySebL/lzcXv
Z23aYI8O0YPpQx2xn+0pPkiMb7LUnyt02/ciHb9OpDWi40/9msVa8b6fjOfZn5U1
BFJuE3yayjgcwFf8ADKvMJPEVQ11GniTCwuYJhPU25CuQQu9V9KP358XjVwzBn/C
RUX/delAC/GevAGpxFf2amfPU+3mH5eeM70vf3+b7NCd1t/d0V84GLE2QrUIrdkZ
dxmJEoM7RutjeazQS6fchKMxOts9RGuX1EMB4fYYrdRfpe8f05TkImsV4JhZMZYc
oonghryIjC0P5CYr3DMbUNMOpUaN4k3QNCb5MINydo6Q4eeh9RuVK7DcmSRI1UE4
oGeXnpF8jCrV8m4hXGVcdmDLFweq7lo9tHCxnllucVGQta/doNUaKw+atV81FTDL
QshHeWKB5/z8VOoSiP2EUBrKEzVnTgYDZk14LFxfMtaTDsPRljLrqyP2oCX7r9pc
4jDY9pJ4RZ+TSA1IUQLDDz+8CV5XpKWb6oYJTYL/yKuCDO7k8J/n+WElxCN6ayyj
Ewsz7NXXvlLQNWCbFl6AwfGaoT3JxJ2IRimYDfvxQCfytWzx4zM/Zq+ND5K08OYU
Dq2vWPkuE3I4lkEusxm9Q2va+DKcsZecUC8hT68FFv1ziFjiB/A3hb6UFd8BmAwJ
HTv6fyVhqImpkYdpKtcJG9EZKNS32bOiMUlyAnNibTSeuz2s8FYGDqOf1tUqcxbJ
MAyK0zkbFS6TTa7OE+tGYQzIMh0FxbgJUtD2cFVBqgxbEUmeW0aU/0a/OuRB9Arn
qbzIxXfRGLKosYjiuq4PtG7HDUjtHJbx+5/Mi8o7let3mWD85Yk2np5QOTR/yh93
m2gpmqZZwkcHmeSBumXf1SLIR/wbRvPGJbu7VSAB7mHn10wxvIRoNf5+YdPZW1vM
rSDdFJuOTJdf2aUEh6eMpxCm9ukSBvAABxX3/e8dofsIXFG1g9Nl+cUJuPlvWj5T
3Ro7CE0QNkgQxkfz/yYRQZuzqZsueyZxm2TJrXroFAAO/Lyf4nxHXCQITLQoSjoN
NbyM9zQ8pjdxjm0FR6nTIUnDvdZ4oPOBdaWdwgztLS9el6tiJfLGJESGV0lFIVpP
T30FiskgpUbHuySPiPYw9z5LPf21+j6D8qAMGeCthBDHKgzoR9w/h+iatelAy79+
IQ+nHKVOIPywMHZi5NE0Q/WYs1oB6yJF2zayndopCamkdn0SwrN4oaHOLXyFP9q9
52LN8NUB2LKUvfcRc/yCLJ+e/15Z0a0osZ71Wm/9kzbcXW7fG5qpNHzVqSSr8zhS
3OU55phcmgYEyuATpj6OQ2ja9ktqN7bLp+LiPQs5PhD2ONANl15sFcjsP5wDmWyB
K7BTdfs5mENR8ac4cnaKjjlOqmhUG1QskmfJccLBOjc25H7jA27596Tfitnk9OG+
R0hpAxIVhjUkNG5x3tQIou1uvLIB6C2iMZEtkAyJZ9OX5srqyhmK2SiVGBfjeFRF
ooUyblL2PzGJ+T3TMikIp/Ozt8+JwPSvsYcOhAow+/kps8MTUjMt5Bho1sfKPfns
WJco6m/kWOMgwYkoj6uQy5m+UG8rHUHnw31Gwz6FHiuwFlFfdWrQBPiE2JPKCtrr
K7FufPZslVI0VZ9fo2FKV25JQxDFZCIpztin+bgjpkrdE+Vul0ZdWdhbs7SjcTcB
sTzf/Zl9F2KJqmGDs8cyLltW5w+K+LXP6RjSImMojupYUMASqKjZ+Ls/vGfFcunf
pUmF/lfDTgsLEWlGACD722/aCFLmUCEZIxKpzqsaOiW7GhQmGdjU4w/Oehc5DNpw
42Af9hn9qK+uyUopO5TWPExTMisp1B2ze90WPqFsyMOvMKX2Mrf2opItAx7z4sM2
SAnHuWMMhMasr0bGmrisSi3wRaHomw8ga3fqmSLK3FyYEuoAfg57p1tqjioUZznN
UsSSbLJdfyKKEAvfsXOs9jxhHn9Mb5ZGTCxW+b3Y8/vPzfdn0c0RtVd1ZcrYQc9p
qthoMA9EwpqcBfeQUcBknZ95XFHPLNCOjuCkZ5bckFqZ8ayL7QRaFcEI8wqdKLds
puEVYSRdgzqSQVIp1hjPBUb3a/9Ju2asYaq4P1sYRnEIQGywNsuzoxXeNMiGsxzJ
spKdA+ltRky+pmWIh62FVyupej0iOylPPWwQ7SjFPvYL9t3JruWJHP0J7566FFOv
302/XhBrXK9qUJIG63DCP+sXi6qLxSqGShFZdGdZd1GVavTRBuPXMeI2z3nzAcE3
r61KsLvnZr8HOrX7jiLSwq7gwpFoOyApDS8RiKtR5Zxg+hAzYii6XEjq1yfG0VqW
ZiHijZwO9CsBiW1rpN3vQxMZ7zns5eEDoVl7nQ6cgr1CBdWe49/Uf3YkM0uTgJ8a
eMADTx0ccCkh7VvcTi2ta8RlAhCFrm7bz2WjkrT97+9iuDrUApLej0CRRfvg3tL9
gXYMxdnG/7iZMyGQSpfCQOHTdCg8szKIjCDrNouHDvs0KQV0MTe/NeXqTSLLguM6
fEQCbJa3bXc3T3GH1sxPe/nAthBhCR87VagprS0QPBsC0sPv/ueFUfa4BEvryjjP
DvsHDJgXmwLaoonUeEeDHFpPF53qRbIjOxInZTLcJdbI9E4EcAP+s4njk4vgbB4D
nKOMXKeRShpLRtuaH3snIqKq4eUduyvr4lJ/AbHjZfcgQ+8fh4y6G/Bbwk/i9mvj
M/FUxHzXITswikRUfo4xN6BDST3Qr3m+hEq/P8lcuR8cDeu5bNqd3usT5IecON4v
9LXj/FJQ8ze3Ox9X5ZAwHRMxlDy8WMKG4FeCdm6+p25Y8UnbwKShlXxdrAiGT5OA
a8EcET+VXj8mPMKVwZHkL92FbZ9nb16USw8x45JQ06kvBkQBfG4GnPMCff0Krqwe
EcJZy+GurXl/yDTB7/l5e88JZX9IRsVxPrb7U5YNoqpBRG75I2Md/ITnWXZTlJm9
mMSiko9vCTkvNDVrwKvoosd5njN/VN9HKhmw1tghq/kzVmDZnW0ItWkSKhwBVp+H
RYkvSRE7xO4FfolRRfSaTctiKHr6tLxhFY/qNGy7PqKzokaENiqyv3kaWYoqZKNe
m4MldxtL4g2Sqk0bkXUFAY2EsfaJypRBoFMppo+uJlEjDiQStrmvAY4mwlm6VXgK
QWTabokpMlJtw7d8UJ1CBojkuTwPcCqYy2tIGdksdwRfnluZjuc5bnaPt4QShrpq
7rSeF6lxIHnhXSiOgVHDz/vZXNOQEoX1DmFm+NzPVyCcWdp3IQ13wGh3wwB8Zocj
HWyk8jlDccFvDtmSs1fatyfCM+UcxD97xaX+u018sZ/pOXJIUDI8dqNN9iVBzvd2
dHfyFSZeihor0IotLL5+3g81wJgTXRySuXkyo+aQxzy9FIzyU1XGtxfvZBKgC71b
xt5e2yfODKjcmM9TDawI3d7sUyP4OwDCk5gAvT7LnSUIWWA9AAQefxYCXkD9QIPg
3BXJ039qUuULIT6H2S3tZgF9YaCg5/A5Y5b7igiVpOBu/u6QvKIY93r/iomajICP
w5LG33WFsqastCkEmE8tVeAmGk6vYjg6NooF2V57ahxCYXbah2bqGM4GMYuPWeR5
aucjeIb0BhxErevIFap+p1q1x/4CzgVf3uU/4PcK6fBH6vMJx/DqgdKY2X0rwd1X
mxuIJhrOuTZUXWQz60UiPKqvbJtHOnooMJWpWHQAJwXsKlcLCjmsiqNDNoARsSau
ynQsDBH2HVaQNC9nV0ocj48K8DJNeenbzZUrF68nPtIUUhSH0YPh9FWweER/MRhL
JygghrLoVT0zWoQHvceHMIbcxQAkpnXu3ZqKmIQsM45eOhyQ14lw2dSPkYWsQY4B
DmaViN7ExzmJ8jAKIFKKVWT1e4uAvn8J56STOkXKkffwjWmdCdjugwZxvBCk9vcz
Y8vSLv1kT91ZMzr6GMg8Qs1xsf28FxsAL1z3xA+uH0hPDH0QVoCBhX3bLiegSftd
nhEA+U9mpiIGVeeqOb5eB8yLWmviH3s0h/lgQXE1TbZWaeBkCOJLLzn4XvJfbqAB
J16MMfDLgifEOXoSykR4km4krzs9VYlamvfvRWbYc1ENsEL8kxj9wQHqEWBD5NiF
1kamyIFdJ83Ufjg/EspHPTFMGdwcV8Ns8q1PrS9SsFRcmvuglDlpKp2xhwwaLTOe
rUU0wXValfWmDPHGJVrWxdGale4fm3iq13xieZvRtI74+jet0Ca6+fsRjZep2971
6fVSDAE7iE4XAyS1e1JDf+xWYY/QY/MEQnxyeK56iykqF8fxCD0G10eol+tonWN+
yIEYoANNMSMz1SWMQpEMh2auWLDBX9iQ5rxFVhhaqbYjp8VL8XKu0khq+z5rodZX
pCJ2C+OWKg679qq0F3+s92HtRwtAemjch0xYxAsgiwNlkZKIWWJsJd0AYOnuCdy9
3ajgxpb2VAo2nOAc46+yE4hzqzAeCk4aW7dHEH8izO/iYYDCDewQoSqQ6sJ+Hbra
wCPJlQhbtUDWeR6L2VoWUG+uSOZCNPzgBvJycFq+dDc5h16wLNkI7tZq0MsVP0ia
WnLVEqdFqaB6QKexnczaKk6iDGj8D5y0LLF+WQrhFiYz79z8Pxvs4HpF17AeSam1
pt5SxVGpDp3J3gMFoDmbJq7H9CMnJFMZQk0sfI0uwQtY5Bz57qpk5DNvW1Gmu0t1
yG1eWQ/McYU+vJYeLOHTZ9q5m5ee84Sx5Ms9skoU6QjfAmhcptnxEcz5FStz4lwQ
KnPmi9E4OcoZwAmXPAt99zeSEJWCm7i2PEBfnnAy6f8Gq30CU0XzjRCYCarydhZm
1hzyGrqH/MR7Cejxt5iCp35CUdOhBF1aWtXgaZokjUUxp+qnNx2fzhjCUwm/KqTH
XcMLVHveudegSnTa7FnO9Xcgl31KxASwHmBlNQxEFK2WRnb4SQSUnrStUzgtkEbL
Ac4JkZqr3gnxk3l73k6sM7P3FrjRUSeKCeV3Seg2XaN/b/UTibNB9NKKCXTYgCpp
txZqsw9TYFoXQODRAjUZ94QASzej9GshzCItJyzzwJDN8mzeNqbA6eNOc5hnkE4u
t4rWotDPNzdd1k87cHxzrbZMf8CMuWIRtadZfOgupceOM+ZYRxWS+zIziyh7wpA5
wfo2mctHFRwUDItmsp7BuOlm9t1j2E/QhHm1eUYfNWVms5YkVovjmepNi5qD+SRo
6opLDN5f1BKusukOd6PJzwHyyHe//tpzcxBjZBKeYHH2UiRUGqnqEddiAl1aYWs5
nYKGQbDRgcucBJkIw4L0Kur1knZqB5MT6r2+KYbGBoX72Wr8lK8Z8dAE/p/YkXHw
B1NZ2NFPmPo9+VxDVpK6kcbPRFHeJ/YeEtmjOUxopXxwcDmwL2Fjr/jP/+jvTzVi
aLdztbTNPMGGMzrxmHRZxFTAAxUwlD0OAPWlHgJe2AOguzPO5mkfvLv0so8+cA4E
dxpqLohFnUt+f5zoSw8RQs2ABsI3pix11ibiJBVMn+BNnmFXaJG4axbQ8OMhnHaY
3Llkw6/IShKOBpL/0Ybnowg086Ob2+0Hn0R5Au24ysUIQjiWOEG2WRaMXsql/Bkj
8+6sqhq9+YkCZ8jJwatNGS0OflkAB738rIXcoEcaRHbIXK772r1j9ScwM+7W7pCZ
b1FeRXuKlGMaTWYfADSrTkBscbXV8aa6ONtL2T1IaYyZMI2adpn2+K/+DfKk0pCX
JUB9WwJeECbiP2IldsRDB3Oi+Usiwqv3YfS5xV/FkClZ10UH0nMLJCLvPwpQ28Qw
ItqlcE0hKOj6b3furtBojgl9y4PyAoykZGEfwgmGkT7crw2LnRZ6MmqjE6lleGZK
d2LFkjqqeggD/SvwAw+XaNlQzJmJ475xMDYPrBvZCwPf/qijKErBFFzgPQkWrpyx
wmcaOFWb1fMDSYRREIFSzSgM8D8lce5Ki4gdoKQDrGM4xFJakiHu1VLoYQlTqNtg
4sAHEudyMIZw6vDpApzFR/MBRZHccyQK77LNBevNvalQ2OCb+ZFtAUIhWPFhMhOh
nBzTb2dVBAQLC5ECxvnAmk3s9dAkKKoTjKSFOkCC4nAYFqLYQQnEIAGu7IduVk2S
o3bEP56JXipAC/PADmMtOvs8UR2zX1aipgR/25/YbWMHI9pLfqNlaWiozhVSgmbA
AborlpAcOHyO/l0GsNV3JQYu8TWHKAp7FdEK//Ic4BZZz9LIMPt92HwIikwcLuV6
0EKsQFpeJNboeDTo8Hgtfdnp1HdKZ/ygEqMRzMPOBPn2VRFJByHFoGvX/pZ+T4lk
sz6+R/ADGoMGRDnjSMbM+RmcEKGB5aXh6PU6Kqt1uAVVW3cPSpLfzTnf/toOOmsj
fio0FxYJlIiNF7sZRcpRQssZTOLEDm6xgVEtXDRM34EKEMzNr3G/dRP+jjqE1M+j
WI0Ylyd6u1PacM4FzBsty4lX8TlNqTPcR3x9w/PCr7xqI96vHALXYmgvKnx9iUEw
u46N8P9kichHhdySbyDiEUBNVIMoX/fKmTxaHQhjdw/YGSuWouKs9DeP1kCWvcS4
K4n6XakNEEsWZxM7F3pjB9HvPK8Oh2eM0fs6l7k6LcZhWuhp/wnhFjJPEmSadGYb
33MpfI2rSjEx+qs89mRliWe0CehnR7OgwPQ60s5MbS5Emr/rdVSZITsuiCULZn3N
ytf2lZi70OiV9vJzqT61F/nM3GeosQYe60o4Z8Jk06R7inYwI8LQJ3YvXzABpigp
PFvXjpDbcafNi8hTM31aQuyk6uStVyLPCP9ZMavszA66AMmC2DbH8HJYfFkNXM86
9PKtkfoqSp7uMjc8DqM3mhFQQ1g7AuQxtZqw3QMexlSEL8fFGk2Fc25xZFn4sZFM
q2Ywvd0ksDN8znW2sBt4q3QQ6skx4sZRBQS1Eay71gn7m6TgCMXf02VE48lvb9d1
Ak0qLknV1hEbNKYyfGLmelSb/O74DbneR2vvNKPbyoqMXRS5Iz465avsDrZTQ2AD
Fy4lNrRDoTldXndgIdPD1nGbqvHKlD0iDJi5EbTwn5hK3MWSF+ZJfnE0A/fmNgIo
4hDnTxR1Etd00luxjYwasbuGsiVr0weBgNkvnu4aWRw/xia+TJ+YQfkc/l/xz+M7
QOO9VZF70HbbxLG3i9hmk7oHV6+zKsJXWzzvNMmGtgnVHYy7iam8HtSzutMU6gMa
KfTof4kORHVVp6AzmVJ+U4MDS14idEr6EWsSrLHW9kBr9ObStvlQ9IJD/WP5C5D2
Mc1Jkp8FYMWdfAsYvQA5q2prrll+aP/ENjDqFwEO54tIOHoCkl0okCy3IYUBQ73r
efrKTTKxurco05Ictp1tIpEuih7UW/Y8vVQx9H8boR2kmXmCG78wlgPqlfH4+DHr
8lNI8+KPk5gSDc0dV6m97MxKRYUVoz/kvdeolQNLYuqyYy3LbTH1RLyNDH8sVToh
PjdhImUk9GgzpctV55TOqarIt6Bs1mq+mZUhiYqfC2vCCNw9btYl+Y94b1awjCyR
/M0An1ZwJSB8SRLCbnTRCCaKpdj8usR9dw2MV+P6o9Y8crXmS9svpVjqsFHi3hus
1p7jK1kWNzrKY7z6Vi5OiGJa0pUwd6NCde1Y2HGtIzAIkBAhHbyvcfk/hhl4ui/p
uLKmlxkpQSZjvs9Gzk7/WVOt6mKL+OXa+K20kBNklFUqxUd6ZxQbz9jld4+iPFw8
O1ivxcsKfrXWFufK7LxG+mFtzDQjh/Q2S1xL9KExUplYWnD0WRp/fxzPWnnd2xtH
UqfdSlGJyZH+VLi3UmNsSEQvKUf2OP/FgqAIDDAySm89qvO++3VoSIAf436iNhbW
4CZmXbXkRfsDRs5iwP5XMMIxRXTlL4KuRLODHZTzj5G2feOmY8FBZ7j0qCuZ9TxV
6s6hHawzNqJ/KhJPj5LIF0dfhoACvL1oQnjgVg2S6QFRKI8k6Fa/h0ioALLI4NLJ
AENWMD3FBggr0latLmgqg7D9qUhDX3kTR8H7ZZ66fDIBuaSuFr5FjAiDosIxoi9E
lxfacv/Ck8dzFHHfe+gSvJbV3yq4P9ufuc1Vc/92FhxSvDpBLbUmi52j5IJ9iZS1
KgOmgHsDuRWklvs7sFT/CyDqfYTpcteaIq4gMqre+x4neK0JTQD5Vr9mgNdYcGGp
4AfunWCb8Lox6rSuwR6d7/ZeTnMThsmJJXCodMmAr0OEPqr4RR3eH5hxKq6c+BI1
7Q2YC2E01p8Xdd3axT71JXhO7xQ+tFyOPAZLHL33S6fC56s4k7YCgRkOBxri5UFW
8l42Gjl4aw0I9CAdSKxI7bxvXUBRj2oWIlI3Y3mzL+9YHaStgIIIR0AGZibPTUgr
pLP8jeXQTK3OkPgkG+NZRGRuaI2fKtBvp6Ig07AVEqgXQKnNuYURTw9vw/ymTwdQ
lg4EwMFECKE3p0OX17tqTbXMF1213jCKVclKONwUiRWX6/l7/1ixPtQCdvn/OA9W
b/Yl7QILXd9vCT0c6FLNJwNKOEOODYj9i1YOB8bdrGyfsVvqss/uf9pjtUDBKV0v
ycrt4TNWxgkhyKK+ewJnwIKUpevimXAQdHMg0g7qcql7AAkkFsAGzMMuiQMCNHRH
zKAGBPhJ1fxBvl4Rd7QDrMaM/VaZJMBDZYvco204zHkiC8or4ZBdd2eeZGjv6KjB
9nwffd9uIbU5TXoqMN32xFUGREMGJAIUmneyAXhSxrNhgfsLrCTmYI8OVMb2/Rpi
KpxI8dLv1EdFjUx+gEBZiXirF4ICuhG/JszbqoikWGqEWeuqlyrcMSBlQYVwqISP
ONi5PEmN1EoWNwWD6lMstoCgxb3sDykydgkpoFXpMRrP7fQtfRZEkEGd+Cr+1rkh
30mmgWCEzquyUKv31F6MSRO9oaxClnLusH+7HC4PfzCBAcqzce9AZbqKJphrePzz
esIgPn5BgAfek53nN4CdoV6SpEZ187moOxBliBEtt5Hiz11BQlbgcJxO6lukcsD2
AATT3hv9urf/+4l8GirXJYl7g3j+agtTU0ITh3skEtVpH6FxRYBX+Ez7MQ22tMCX
duItqkWpynXwb5PGIjz+latbRDVE7PxB8Aa5ZmYK35JAeRbdk8wqLn8cT0AZiHAx
cjtVOFSs+0fioTQOHHQGKYBVcQgdVcLor7bG1h41uqLNxJ2wg7QqiVUo81tVK8Ko
fkhkysdl7jYwz22BzkqK0u5cM6WFAZLcr5I9fCy/TFgXklUxW55oqnNyrOsn+NFz
3jutJBu7oUJXsgT4wPTcTA+rLUrL85NCRMKVIM0uW48j1VdnhUOqr7ozIYBo7dku
kDoCzRuIH/NDsDXrQJAcKoaXxSHqrx6qt1gaftW4pBk7NPVzatDOVduk/u3C7EuL
kTEITM0No5DlGurN/91oil/dgSxP0ukq2zWEw7on/Fb50vEvzXfe1GGBSQy5J853
YLuDyUWN79xaBWLrDDdcNEKRYRx+jA1Yb+OpxwkcIHz+SvdP/tWxOem3V/91/ZuL
clQJDMIhIgNPqFdRGNtIL7JY6Tsaj37o1nNr0ZnQVXHqnzfpnHxMpOx4MWmrfROA
oVPm6v0zdSSijWHBgnTqqvftdYsfOfFySIIpiGZjfGu+GptwncCNW837AR7B8h9f
jLUsHKdeKNAdMyZZ0zjUoSxZhlOBmYgtiL0YUFFIqkY65cUZN9S2PbDRN9o72H5o
PKK/rp2SHCIUrubNR3ksEZdkwS3W1umDwBvDMuOvrRKVtMyjHFbh10kX5pVWiIRG
SzkxDTJSHYjguf1j8d1ToVfo5B+99qXk+ykNJp8I8iX/7oDovH2gXVy72SzN6dsm
TzU+52V1rG/p3z6xR3/3yOJqSwXACDlhJ6uXJ6e77uOkwu0MhLsREnzRJi5F32XB
9ic9mWptLK1MkE1bzt4ZvfPcb9Iql8le8SJGaRTceZcy2pyl/k0b/2F0GLuXvYOI
3idxHF3SXJwOtnCEPdLgb9F86dlRzqTz0MgnVSU4dnQ9fyDtW26BqtSNSFNVhFwB
0BXXSoe2LB1Igf6K7XzXgeTvYbS8VahrbcJHIh3mQoz3KkvknKEQtiiHfCvgsTU6
JW9b4odh0T5hvIqSZilQcLyIouvlpglK3BjfT4T8BIgLcDfGmi6N79miSLBtFQni
mG/JZCduSgt9M31IIo6LI/RJd49vfgbSIuIsbL5rDhtV1TP7Djxi7KW+Q4Mk6/Oi
YvAO6D6CEVfh+s0Iip8DtfxDGGC3zuVZ+YdOPDmdynAZ3YInNDvqG65w4T/SgOxj
aQAMhcAZFM8mGZQJ9VxruD0M6c26gVy7FfJIPDUTEbmoFoxgC+19KU4/guI6j+nq
v0O85oF8c6FtgpTopS/rqmLHBTG+bpUBRyKcvHzshr0Lb84eBdnqyZ481+ViPCGQ
tiQ+pHEFGZWxA/Ntk3scS48aKgCob2H4GKEMC3+shDGnNHLPymg68oD4zO2fGUbh
BN3b9iCoIDFvdJVKHIZMPUsfxuPngbsIrWSqyD/TgKH5/D2uUBJoaPov/dY2/GL8
Zsj1V31xMrWs5tG2RxMWUzgPO04xDRzXPtOI7vRGY2+wFIHXb5TnZcp70XYTVouS
y2oE4Cg9MqxcpA0brOVA6YCb2nfYJB9Ry1fesaPdmQKpR9oQrNbiIMKuMYUjg7U3
F41kU2vsSl5GjjdDseZNUDZOCi4ZryGJcg/Zo53mVYSiaekALSx2G2tQUq+6eQer
7jYiBcyhAx+QNnLwH+tQCNHOjInFEPj5FXwx+tVrFvbKheS+RREBIWreuI2T6POv
uPOzD+v8ADuNxX4HVh6P0LntpalglstH2fAIkAi3ce4N38+XBjp8JJi9CjPvAOrm
Stgxrm536s9jdkjddrU01M0Nsz9WxwuHu0yHHOM5gUsc16x8MYqr1QEizdaGzXs4
CHejL4L5m0vUruVtyGkUpBXOa1mJLGWcLr/QBKM472oyDDl9PEI+2dmYgO/+s3Gz
WlkoqTxmj3tHenGCVgj8megbskJagDg7shRIR3bCqQMeUTDKLhbfFok/Ej7hiLe1
EChKDfqdaMStIkbOp8hlr6/sqEuyqABBLiaDX9GAP3LsUdZ+MqGwdFt9dS1qEfhG
juKOAKHMC28Jc7tceaJJXQc3eAY2vsn2ixBeH1Lp3kS2u1PXyJ8fE9cmYblzx00d
lrw4seM9TKcMsjtTIdZkYX+XN7Ykom77+4nVW6vRYc6CqKR5JReGzKi1EUOzWvf2
QsKe9KLwF8QEsm+f5hK96/VVAPncsJxXjJ/9pSH20jpWOmWeorirX1QqzfR9zfrg
O7Uizx0k5UoF0oI8S5PkcA9xOoUj8IxTquhxHdZtKtzd+E0lzlS/EcYrb23vr2QX
p7uUKFZUeGUlaDz3wSZRNiclG2kAdrJf3PO86XCtOa7TblnzhIfczC/2mCEv4FS6
/8CHBnHPHCQa8re0RTATollfqzrE2qVRwDMIA/ZQrWsJqSCVqerdtG+N68UAELAG
sdPuupmv++2VM4Hkz2xyKI6xnR/JCHSEGwaNXHFjNb8jr1uHC/QC5v5Leo6IdlzY
2Z6Dyf24Hzwi3sj9iRs7nu/OSVEKf3nfgCx7kUVq0PEPOr77h/BTJA3mT883DmIe
SSJB4B+Gu420rFDBquWbDiYehM5Ww4NS2eQ3f7g9BlFpt1n/FJXM3mqyKkYbkLw7
82zpy5g94rAHsjM0d8ZSuIZq34b77uHDH7i2Vx2k8BgBB2JlNrZa2LGNDAF3Hg1n
DccBT4235rq7esBFsYODzsE5qvyBCTS3Xy2XGgHETiOWW2AbCMWk9DPHMWNxHtum
fHi6n8F0wYSk2DYz65t+2Ioo27HJIqvhIo0XXAUp04iDdwbvwOGEd7HFRZLQv2BW
TZuiCAMhWWW8dPafhQYsrBA218Rze5xIV+3P/DiI4IZOV3DgOgIF6G9duYVzHp8+
D//1dz8suPQmrthFvPtEqcj9PG8uJWzITTAzzejOSieFB14P/ZNAS/zvhDE6eQt+
RBw5rRmeemPb4khMRi49yT2Z0oQQnA+5r1zI0WIRdhYpgHXDS1sGhBc6dveQMpNx
b1ELrNFCYo9ohKhOJmVRdKHdQcXjRZQJzLlIRPQFVjQzHnZG26dzBkLbWvhpr5b3
AMt8Nb9IQ7T126HgZqgdRBxeb5ZaEfq90WNGxoBuu2Hcf4Y8tmfzv3bK6gKKi5go
g+rDVdw049U4F03JCudCU8dLpx0O0n91JSzseB/cUytdPaPc+8SU8DajIEYf7zKR
3slGToGjqrqi6WVN/qGOOvj1M5Hv6ODOUTBzPDORHxkM82v7/hKmCdIx4EbJwO0B
bkTTHYYqfpJL5Qd6KRAcZl0RejZnxH2K6qHGKB1aaGPmYhuxBsl4rVPNOTIm5N9g
UlP2taV/dWSKqMOnaSgw/36jUh4HCK9Q/bBOVE2yUqDBdn4zBlfHITf9Jy5/fYMg
A+0BIhXN0rgK9HTBIY2MXDAVnSudp7KAXrbtiV5Vt6UoRQalg4iw1Yj/Er3cxlDm
CVQuIDhYDdZjNRN5YvDzp+HW0Js+jGYqBOhb28Utf6hlv4blsvk5GdoaZxRGaN5/
gkQpUEOXDAdgfZMN5TiGyBGpPW41r70dXEft4sQNTeN57WLifudPlZQGEjahmerK
deml5PDvni6R5ngCdGYylq+yhRfnr+noKtxBrOA7PzgHlk1im5MOW25ey1ELiPo1
L4izA/j4gAj0e4eKBkZjhyy8sK+E5pjo8fTSyw2ViqqlZe6zVSxs1DXWTvKia1KL
ndDDGCL7gMa4ROE/OMYhAwyJXRO1wZ3/Muohr6qZC3/e7fMeWaw6Z90SI5KnkSHu
xig4hU0j71JEghGk6UGdn2q47xkrQb1QOMHQi4ShFj2IsrXDpASsVgjFoiBtQ9kH
kavh2MfjzPTV2frxGrcfq0bPSIVbwqd40j+qoY/ahc22U8XxGzS8H9mzqoDxLvUX
1Ct4rOPvTFNiYFCQDZls+j9aYtNgphZcE5m54Tik1/evhVobEhmrc4IazjAvPT5O
sQxzE22KATELB4r16LBCe180QrtbzRHubg9RHl5sQqsc5iIe4SIMpOr/zd0BLTDV
2v3nB6KJ9j9kZwjDQScRZ7Pa2esTcmZQX8KCqfjFvthMoZieX04f8ytbu8QL8DZH
T8BEL4+P8V/czqDZeeauZYZ7GdxaTUf+EzDwx6S6CpDOx5AaWeIo8g4ZAdi2qoxi
bn4FLZwY9UBJYdFJaMaPknp3x1gZvc6t7hClvF2P2uEVVeEoMgXHedJ9aPgNqvit
4mUKJe5mPJdNIjh9QJ0V7AwGSt/kkwcUKNtDnIcrrKfZvHAkVH8WKxcpK6h0NKy8
o9UAqG9v8Nuc5koI/X+Wo+K9PCosE5lnBsa6qs1MUQkg1FH+pQ9dIbqAXOurD4Tv
78fKnhtRRkneCf+cba1UYmOkfUAvrO92ylXeOZBpVoICBZDA1m89kO6m4LsVEUqK
91WnIlJfNAu/guvjXvjkNqJmgVZTBBss3R1Ilr+bmHYQSLz3bUsvqGwIHb9Xj8PE
kN067uSIjhMXxjKUplxCRkKJaonRt/s4ndoqBqzzJg4nz0KjAGLkV8eEKWIjAopK
hK2j3BWGTB6cn+hnzhIQQW7ro5F9fIHACwjJUSwTx5cZhR3FA59rGxN55rAqKZVe
OWv9p/4l8Khs1cbUzKaxY65OJZgFhsd6YthdEZZkD9KMPs0WUrjWFW0dKbqI71/r
fBZdvYOVZz+pb4RP/POdr8uLgAEMfC3hOjBKXacbZf4WUl/z64Vz//t3SFQc9UeP
SiCyUnagLGGxsR64pumOptBoC5cy+KGH/J5dIJGY2hfk02xaQQWeQIsy4BXDBAb+
VLwFHOpXbca/Atv1cC9Ya1HMZYI4XqFntAtPaKnV0n6aYw4Plg91qUQVblQULiQG
dKD2vd4snUhujG/whtHT5yHyZcn0/QylpB8EBrb/8FqWcfqvGK/2DpDeeCxiImzM
bSzt++ikCn6ijtu75zfNumeJIPsfPLH8bVfBBArQRYAcEf5nuB6LROP2A8wI65C5
xt4LoteYILXH1kGnQPOu7lGXGqRKXnpdsyTg+TLtu989fHCgMyvI7CURqyw0EFk+
3EU6uTcbUSTCDrvrJmYG7re3rmuuMwKYD9ed1hbfDpZRFsUZss4wdcxZOCCzK5gc
wrzN9ZSeBjDA2kQ5cuXV8Apu2chniI+qOeeT7BW8Nw3Ga+jk77ftO4dL2dcWlbsD
Ixc419Gu6Zr06EA4ZcV+klBb583M7OR8/ox0yFxQ8N5labMIWPjI6zSunxDF5lL2
DiObH2UxA3DEx3+wNgL4P/vjaL2fVq1apo6fdlOGvFQsA+7u82RbhllQJyc41XYL
mo8uJ5WwXC2Invbs2Gk7njB6tObn0H1A+rzgPlKzRm1jw5ii1czLUW079Nf0NO95
8f3GAaCdkmVYsL6nb7v6YPkG+uRI+RHvMUv3xxpQtzPgBJWtv3UmF5fcO5yZOBl1
ugPDX6H66Ph+/hNBhMY8wKLQH1k1CK5/vyx6YJdMLaaBmbF0MAZLZrkwp3l/+sEn
3+g+1IWcDlQ+aFaLQsvodgiRHmbsqxda4wEZsqkaxh+11oBXMCV45MCqA1XzkjIa
tCgPuWoZkhA8KZEoFE1JBbbfQmsnW6KLWkhEPGyYpE56kK8V03LGaeCbl+FujxER
5c5QrMYqod02UxHk++8/C6Dvdcd/IoBJmHPez9Ap28O9h8ORJfmwV2CPWXZBSn+L
fFVi1O3KLnvidiM+oVT7jwk/he4+AaHjasLWCPeO9x746GR5xBWcfJXoMc/+xXNd
n60plbZ0WXMsmBprYZpJ/YJjt+EnhV0lwHkWmCaNY4h36LpDyo0BcAM6Q3KzZb5b
h5MBah/EXfWIVe1jmu6yCN3TcprPEEI/kBomSpxt6zc5twmwJUPkKJKuJM6EJ2FF
l/UUAnelVWVMWuwtIduqinpKLt8lz39J4Iuzf+/awRCrf0G82kSxV8SsAE9snygS
2o2Uv3DAfkogjIGTPQrEnq2VwXI3r+TTROXGrGM3Hs4wPf/Znnb1s66JMElI/Ntq
maonpyJMw+FluFMKs0g83qJHp7WAIxXoWJCKFmBdc1Eat/XCdE/3bhh0tY+FcUSj
FhR8EiUtruxYEWp7BZl8FT/5bd4PNmhShKIQqdkosU5ypLjkdC6u34G1XjCSfWil
Fvl6p8WuAhxjbxwCSpalqjFQb+Dril9zjSlkLDLn7IrPjWUbMqzGJZZk4eK6bz0I
GO4xhyQ0Ge18nqkl5ihrQG7SI5z3SiY2xgyW/ROMAyKy9s/2FW3k0AD2wDRUGm2b
ES6A/T1sNgn6EmHQlS9CS4pLGOarL+M0B1h4jPIQMdQgilHe83SgYhuqclUmuhUc
mAe92YOsgvupWPPc23brLjN0+Iw4poqGl1aL+hWoVmEgkNsKjC89v+1X1I4V768x
+R3vps0zHKbEsk8Ommu58NkF3SnfY0Wmc9rvVysP387QRdZOTEM/jTCVOJMUgv7x
6nTKVUFl241/4LuOb/axBJQmBDArJONFjVjSwgD2f6geS8ZVnI07vt0IsqHzasKC
FyOKS7HFc4xRy8vW77jLmxscy8FwBmFSnHRHbPS3gUzBWUXgJ+ossifDGA1X88u5
/Xh36R3gSbXYYtjBDDWsW2GpDYYQyvrwN2wMIS4ztf70WUYYzsmIZVqutnVY+6sr
Clu/qRQ7uCCmgntmuLr03Z9LyQSmOKFDkiJkjTiv9QuDFQCP3NwjK26+QwlvdAJu
CZ2+iDA/8wDFvIEOSk+RFLCRdSBj9R0jbvReGhLFL0NQrfvkTkHSOIIwMxCFb8gY
LlQWIJ2gJSku86cWoJYiZ0gDOEHr2AK1weQcFjOUhYyQMqo2w7um1x8lN/NmmW9i
laac585+KXz8t15Xh114cph9i+CnMWxYmnk/r3hxHfcvu48LlWpMJQ5YDuS9kPWP
df8UKVZBQccPSkc6AxZl6UvdRoEkNuLcVJgMtbHjlYy9JWA5wWs70s+Xoot4opz4
zLRdZmLBeXhcsUxB5OOQgmzxHeHomL52tx29/a8WjCU8bvMGnxa12240jX7oAkm5
DpkJ9qnr24N3+S40i1LgltBpI8gBgTl0HTLIr/7DREKY8d+jPO2T3nRvTWfiQQL8
RAKD5hPGN//L6+CJk/8dj6R7i/4HTGPZUwyazHA3An4iwjylj3XTGa0dw/YVTZ4e
jEejC+fpFO73QtrkGVuxp5UrUbG5T0TCpvidWM+ShulsVfV7sGDOWt1b2Nw2vzpi
e41N1CbacCMcQxPqj5KBzgFtOVtv1kRb49SxPbGzzc9MGr9+5MJ9Ueo0gMIb54dI
5F4WwJzBpGsPr11jWHDs/OtplGWHk6/RjHirHnGcXi5yAQti9o9XjRxvumvWqAe4
RuND2nDO2+Rr4kMJn0N2SJFHRtlWgZ7gQpjokaFGL99dSlw3gYKpOfZjBm5t4oc5
YINoa22C2MGX01N0igJ2wxDfhqVq3qR0sS01juB4GyEnc3kxD3zMLFA0v8LW7Brp
HpzUNh/M3+ifcPxSfc/5ou5roLUGwqEqup2a1WzpYHZj8em8QDLt/Kqi3lH+wx9V
sE5s37MmVV+KFgDl47offMVoLW66JKC1ax+0BXrYkPnkyrzsuhNVaO1HtWD2MgtU
JUVdjqUnlLy6DePNtyMp3Tj0qISHMiBYEsWBr0ZWs8oSYxMRBkfcM68dDkly8HIi
qF61RDrbJn6cwp4zs7bOQFeCf+WT1H0414w4KxcausDqMjRbLZnSsd45bsf8vipa
vyX7xD/xCoiyYJW2nWkGbii4R2XPjFO97KMQXRUce7VyHlc+wPaaGZnmU13wE5n2
xUu9M3xeN29dHz9VbDyHQYhquM//d5Gt5VasFsCRhnNkMSJz6ektxV1MjO8NQukv
11+bkIMMLunAuRXHkM96BMykMD3lI/p5e1xyxOh6s7/FLyZBRgXQP27PnCahl5q5
7nri5NCuecyfItH3k9ghuq8OMroK1yknoXATy6nDq7bLvbf7SeP+29aXWuuo0HTL
A19zstHU5s/OzuuXREBFvwqiD8FHGfi92C1XGaSEK8trDo/vmmTpMSM/ieHBk7dP
Fb2OZSGEBmQmfJnJOnfMedVwr0l6SxDEfpgYlMv640YSfAWkbNVTNrttTJ2kENRs
N5jLhMNEm2bfEky5HoX1m5C+GaM+PgfvYsoGWbsGq3X/6RBRK3wKMFNMyH5feWJ7
tO7DyWLD4BIJR0QJG9hPxfRxPga2qU/q85aUYDJCd0wDl31cgwZ1Y6npy4jao+/k
ZF9rDCejkQDNn/0RFqxUo0dHQSfklC2Dn8Y78TAC3l0xG9TjNjK5dsLTTIv3flZw
wR1L3bEN+8krGrGuH4LDz8pYzeAD7wSWywrxFpwn9Gly69Ci9uUyZ4sxgJI+htyJ
SM637e9IeKoKKZnV5TB28M1u/RfjOhoFh8K1+z6YwTH6Wp9v+/rbed2Mr2ZU70qe
3x1vcVxoGjyvHZMRVBmziwvW1JMVNsO40mQSli92kxhLBjFo82cS5vLo4rD7lpWw
wdjXrDSLtcGB7rt2kUulVsseCLjq38gMMoTaP5FjXgbCbNVIC82P0bWHBZrpfScj
acXzKlew2qJuXCmMM4nNV4dtEtHJgabAkLOXWu0rAIBQxOQ3+frObDksPAgUR5l6
Etmj6BXQMbQJzGZTEn5sWDUc0X+Lmt+JrpGQJ+02bwHdbbHtPJcJ0rdhAZOpTu4g
uNnUSTeLIyY5joH7PrRTq3sJH/KEef/93VekfGFiVkaWFXfM8Wm+w47ma1+XOgPU
wHJAVm4NRC4Oro5fLqx6tJdG31OjB7DL8p1su8Sf+6TGX3+ivWgUG16maCYkbTEy
06xQF20Zun18DA7+msCvUebhtD+BjM0z2hSsmil1OBfDJTRyFlTwhU2LkMqf4/3w
o9mI96+q+vDhUc3Yf8yaVWqr1hy3JJrTREoBytVo8rdZ/AxCUWvNBR37K8+EaLx/
11+KpI2XzeONig4P4QwRmnxcNp0Z8Ejf2xUVaQR7iwbO1Uokp8x1nWi4EzGeFjdn
aAUZFsawYMqG0Rk3bUXVnP0zwT4iW/9cpbEfLuj+B6vWZdfmS8uWjwppfwsiI9fo
sLsAcSgqRAHvNrjDjSAos+5qbX92KQBLw3jFRq+oicrAIOZIArYu9b7YGxkcVvLu
Ym2VHeav6jdp0djbIij81VynBoRettXB+rYxex8qoPXEfEdde+dRTXy5spMCwPpe
2xeU1AX+Pt72fMvLe7ckYu4SV0A7AN3TZPOjAzNDyUTiwJu5Q4Al11QBRDmq1af4
mylB43rQJw0rE2Cx9TPXVDBVlRDtEuLeHvlbYRa0c1U/7oVkDZDcyUD3d8sCAlWA
PIZmUcgeBIJpvYWX6tk0uNsTnCY95RKyhpJvFoTTe3p/vKaYTjJj8BwRYMn7ljLV
cI1UtvwZbUDz6rhis9pffl7M+I7PVxv4jKAB/eX8kghmuEfJP9DUNF8WamLjZFQg
9u9+gh278/NLM280EOlLbb+Wz9VD56ea5wTg5yAA7UlxsLSUxtmPJKfBqkcfGGlb
mu0csN5sgxdGgcgQGgtY3qjOL3kxKUErk+KBrNIwPt2VlEpXIkac7/l7nTJsnVYQ
H1qFzFS1PmFbJBYrRhulrIGH5Bm17i/9uZql0pFq6hnjp1H9/j+B2o6/2oV8vBjk
IJSiltZKuZWb/UkK3Bbu+3/H7mKugmfKDBI9igHi6IlZ6q5+ORCqt7Mzxqt5+8DL
LRgrxMEDg3Aou3Qn1SRRet+i4p0LqRRk85l6QYUOYJrHGUCyB8sAYI3/32Isa7hB
x/g96CVvhokPVxngXknrEYe3YzPX7FSWYZ8XZfGruKek6BkiMwSfRUn+ighAz6zE
lznEdFnWt6GuWulWM0HB+3gTuh25GqSweYyru3cH156aLd7iz35nduAAKAX2twyv
jGNbXql5Bvpuqt5nO/k5Rty4HyqFv4ouYCjN30miAffaLM/cbng/9wip0ahKUg0f
kgRIsI7j8WrSPAG4o5sfTeQzVlEMBvYcqYXuX5w6efErEbS5lAiH65Vg6h8e/7U4
xU5ud7F7/xQhRxjbeRQ9T11g4gIYO+09KfZLjeICa3FQf0I+jmyXe9BiDSJ5lE57
OjH0K2oWM6EDEobbY432Y4TveYn/iSrEo8/AZBkGpRX6GT0gpHJ0wP5bCrUyLff8
2mpqdQIrSPb1u1m44WI7W86v23go21IpNdZDnrYEt4oKhMUEnuzZtzp6o4DtS7Pg
WsKSkAlI0omL1JVtDKMYpO2L0Srj49TLqEnexa7D3j7bI9He077UkV70T3XmdrnG
8crzaPvAqyTLxZXiO/gTD1jTmNSt79qpBRGVipcSmYKR+mF83KY4pG9PoG2ejFDC
Pz47Y361d2Urbift1MmCX8ASsLeOxKn2eR4hNuJ7UuQnhxy9/Nfqc9Hd6S99+h1+
jKW32LwtrihvJSVLtst5yxQvGGkIOohOrq7DiCqJHF6x2JfqAZ4r9UNB/6nPUBsm
cqPlo9jUvgLgE3IO6hbgeO4+SDxF24bUBcAYieTw9Ha8P8Aw+OdyxCzaYJJz+H1r
3o5oXuHjfUqWXzDnhSw72Dj1O/jO82hJyMrdGVZWDXuwWJRR4ZWk7AszeDlSYPTt
oihnLg+y6lUynsnogVYkjukniftVBwVCLHIw3Fe7blYSwOEZqg7Nrcjc3/cZnuFh
j8uVZWZUl1Q7w5OuapzJ1DJ4+v9Gc8W2v767BLyMKSzctOOBNPby/GRpziy9b3Oo
q8/T80f5BZ+i5ZWjJxvKlttbLkdWKjbODsZSuspVlIk33OBGOLh0bYLyugjepSwm
q2zEY+0Ql8BqZymBYcnkuiqQVelKUSIAxjWgl9VYTLL9f+HKF5T6eeZVwiH1ivTi
lmfvXCHUozEOTmVA82ar1A91IH60Rjoyv2VjX/TpwR+xCDh/8zoPqTVI7HkwIL7K
UfqFowEqNo5J8gExQXXQGw1YXk9qYYFAkCUPzC55+eEEucXlcXkUmmfUe5zWV/15
omrKgapNWMnms++HBAg8N/rGCPA3QkN3DniAJTmlK/24uqaaZUum80itV+Itq/cW
oECC2I20F2mH5KnNwRe9ao//Xx1gf1MY5JuvaxXb/+OEOb2eNpv1r/4xovOw0bz/
IChphUvcD5i0tRRjnDro1KwRGb5WsU94kW/wTf4MtkMc3hWHRs8pZsSgdXpQ43RS
3NQfXInuAB9/7Uxkwr3cZN2Zzy/sLEGpAlkm7+GGrU+dxq3qSRu9puAIo7RnhipU
Enn/ahUEfD4NgA3JQRVCiO+JqWJKEv532+jzuxKjkfHgpRzpvklguzFSfgnV7K2f
p2VC7+elVkXanWqrciGmwEkLJifVEg3MbiVvAPWR6tGOhrA0weF5sCPVLLepaKZU
VgKnt6JLbVhZFrOXaugzWiUKOnBSrRANy+voIw1a/AtN4XXp2WVaXxfIsyj60sbG
jbhytWQbRZV10rQKz2J11OFenwMrYJKJWJXdvEPCT7vXozHUkTyHd8vQJMf2UO5q
Wqx57WxMKpDkkWtQU5fYnN34wxSk7somhKg98o9sHUiU3GPmKKh8nvH/YIbpfQzB
Extuzm1o1yAoL7YixaBwtuFG13VtC/v1sAPVHAXUtlFSLRG3L8wBwbcSr//zWi32
u98z1fAaoC7VIjDXN0nMzgo0yxGFdBDuExEBW/icFPfR0dyCLy5nIEEdRJ41j98K
wovW35cdh5ThAJZ8/EBLzy+aVkD+hBMDaC+jp0I1Finzu2yC7lI4SoAspn3ebzrM
R+agWHITuYXYUDZuUTqzzA83tugn4wD0MlFClnX0V7qLF6kMW8D4iU3MOIJGLLV5
BEQ8BcjF9i58zkC2IN7j9RuKlg4FfA/1qs8dm3u/LBmab64AupZbIM5pT+jg4j0i
77ClRvHd59d3gqahnkOFGIf5M9aE9hJ6yGZ4NALl904Ejvlcm1SUYNweI2HAbGz9
xjgSzE2FLtIUToTOQTWZY5ppIBa70GRrASfFYWW796sZPLQFwWo8bQvUzOghybJt
9IKVFI7wvOX0eu6wj+Gh2AwPwZ+qZO22ougqUdSK5O2Fby7DNCfRloCG8CL/F+lI
CKHfs63LeUvWWJGRQNHoT89Ly51sYdvb9dZiZuIdkPPkNSkp5Ja4Ox9M6wlqOqYO
ebqI1Uio0A8mBGDuhVx4vMpHGcHFC8jaLg0QTIFBo76Jy5VmEfKf7Q9yCE3Ep81E
1n37wNO4lBIGLjNKajlUBgItsahaMpXktPe1mnCpDfkXKpvt1QosiCTYVkNAuApW
g/g9MSg82Hty1JUy7lW65AnthkhqsfXExo3B6unkxlCVt54c6Yz2qwW1PaSDGmfA
n6MaC45nc0VS9gMPNOVfCPFvL91QsK2LfxDBX4AkgJsmD77XrPxBbe/JgUfmMkGT
tuH0mnpIoGcrjdAZ82mN2lOjOUqel9B6XEJzGrC/8zpnD018HAIVLloAaLd0FJnB
Meahy2jtO7hxFmJx9hx8VimWwrIoINWT0z5WURnyyxA1UtSovo8qSHMMsNPopjYU
A5uOXxzAB4YSq1EeXX4/c/biQKSEp5r9g/RApTKGQWwJbE4o37y/PNb99FpTCnkR
W/6TuycfxKLRhLIfyX5NwnIIWj7op0x9ROFBTldb5aU32b/s7jCyifnaHStdP/EH
8pam4s9zQFoTBP1rgnlI6FaP1mrTUp3XIrXToZoTQqkzMIVVxWOg4u8r13PUkLlX
YL4avg1P5e01IHh+fIk28CVlWIyj///nmq5j3dOwv0es2iMHAheB6sXMjt78BUYA
hHQGf6SyyA2p5GNi97wQRMRMEERivzmxLu6PS4L6Y2nOx9IzZzlW8j2s6iLsqoMt
p7fzDCmxD+5Gc7kVVs6n99Z+qorX0ygB108focXAfU1k67d3f9UPbUJLurcwUZnY
JoMqqXEIO9sEkLsQ7HkVWgdBU8PTlmMYdYJLjsyJiqs2rV9AI7vUrkZn5pCJEbMQ
UlKJT/AT+VcnurU4R6ZUzU23XQYKLff9PxJhRJ+FO8H17S+NH3gNYO/UZYCnHpvQ
5nzMfx8GiUMes+JF1UauFT+KPZ8MXSndZil74U3TZKb3PZTRrate1ayxJhy4EDIg
E4Zj24M/NUKKb2ZZ9TTB6exqcuIObHaxbWduPgzSUkPhbS6/z/h22Z9p4LZFRL+l
W5w1mCpJfYjUi6pSsNqBe2FRREIcRwziAlWAGlW7420KqH5p+kXM2FNzC0g/1WHn
T84g+RU3tf1qQJMbt2rA7TOkCNr5gwIuqaje8BLbOAGNBUxta8nPzOCincd5hpTw
2fwHltjnBXZt71gJOv5uy8N8svzd0Gpk+SkJJ2t03A0njh+rtZCmoXEH67oncDlu
8O5CLJxRenbk7TgQJkPTnP0Dr+vzR3fhWpwbBeihJC0N85nt5zCyFDb55eK7AqIk
x9bP5hSgpwHUzEdg/d9NbIKM5kKt6Mz3iBCcgZ928Z29iIUkL25mC+1Pbo+JkNnb
+z0TfBkaUTrjQHr5Fqa0TXqPjj6y+SXENF1mMYy9zM5pc5HT/aCXY1a0ALAKXiYu
6f3WE4NB/FXPZezEmtzzfpQkazpDWYNDvsmptdeqrm8VkYeGbIVWDsj7MjrfTiiC
4AJSV42r8Y8IKisfw0PnJrt3YpQYPURlfKsFNOlwNzzivfmPLjtBKraNvBRPfdOq
AtJpodXwMxNE796hNkpOb2dAcGA3aqf+ms287oYVQvk+YjoD8CcFVY8TaXlwYqA0
zSXF4h+sytrfR82zZFsI3oLvz8sJoC/LEuJVZB+B7/HGkad9+/PaJoEKriZfDr8x
qc0lLEMLJ8F//bhzhupOaRtnw0r07HFKk7wp/oNn01a8w3J82ImgAC/o7JmdsmvH
eqt2kdwHcByZLxPymqLA2eIpSvwxKi9LIt2oos7+GGGqVh5mV+dysXPciLs1zw5P
9wmoC96uovrpDcUHECj9inESrfnJg/XEFT20H6whhaqVtlMKj4ZWCQRRS/iUEBEs
dSYZkH4ZD78Il7gEFUSHz+WSYt535FupFMS3nAmY+B/mBgtrM429uwpGZShDUF23
LKJXLJ5PWTR1UbVCt0jAnwLVf4M+ibF5HkFYAixEvMFeBbSMFEwEoDnDyDRSdTTJ
1lAneTMtCnlq8ako/AAMW+xxYPS9ZduoJDyJ/rjlzUknRkvspumKEyUw6u8NWbtx
gBeLG577y9SHUt8qB7j0q1ZlHhJIx/Ef5o14gLuGDw4TpFzlfqWgdjJJ/Qjz/naC
iRcJMPBhQdJCp3Xe0J+8u7dwSGjtAouJ2t9/p/iBOziXmfkLp7OMm5DuJRsNMNqt
7tkGeX1MDySdsaGt4amVj2nEQG64mvd0FqWZpLSgRJd/16TIxBJeP7yH6ZTq0Ns4
rKHb3I6GjuQ4vS8V8aAx8qIvtRmSnRSoAE04CtSsQNfQgDJTwVB3avaWk0YGiC9Q
NIhSsxF3S6rMRAQxp9gzjd6Wd16huOLxuaotfBiWr2nSsHGNYLlpWdJ3c6ai3HLY
ca0qf2oAxYUJYQtzi9UlvUpNSP5cvYroLR1h6IP0Yj2x1jV3fxbDtwt6SLnLIU/9
FSI+Sm/OELerPWn08vjvXvHEdXysfBK96qDkIhJ2HEZmiYWGu2cfic9Ydf/2Pi9u
HBhzZVCJT4W/P5CCcK8uWwGuZTm88FqMNOOR+yYxWtOUoVl5Gi6vKacU1NAJt3no
pGTWhpp4k5/a7Co1al7LBSfBgZtA2sCclx9d5gJHIh+sz3DQNXdhgbnZHj28zKc0
fjISLvszKeIMlTmsOdJPqy2hnY0kCOTUfh7kfcASnqdrpok79iRD9P2vVlo76RgA
iIgZzyrK3sUrSZ9HtrJOTPtbO7zwrwdoXDtXUq9XPK7JHcMEQ+xFcwIM+ggkv8eH
uA81KCFSY1Zj9PCDfNqYESbqtsXS1j4kFH6jF1I02fU9pLIYVuT3Y6de2l3WisTA
KPFujPf8aDsGcQ2ywDLjNJhtmg59QcEevUXW/Qg/Opnr2giRqijMfUne95Cx8pqu
XPuyS2ZPhgckNPLVBpAyTb+LJztWN2hNBfp5tFQdxnQC1JkmfV4nd0lLCQqno6ly
Obvu3vIMcE2qQD/tMnONnY5DTI57A++791XV8iiPVr17BeUlHmicpX9n3YlLuCEg
DvFf8GRCiFI8CFUdMMQSAPAZmawbPckvzShME3WafajP5wvXHkLXTv0hLmxepjTv
iAK/0TXoPTDZcJcX6azdn24OrDtQQtTGvvezayhl3Ig6q2KM4XVLuRffLv+Hb8sK
q3rj1ZSG/KW51+U+Z0ztlyiTWu6hp+hGIQB4mDqFRVMfAowQyafm3/T99MfHk4Wv
GRWfUZct2oiCsaNgrHOVy4+C3E/VtnZAHzsyhb/yAGisjyWFjHBsztJszvlBHZkk
CulzJRTmB+a39fOmYv1uVOkOTgS1/qCF5Ea/1NedBc49yrFpUQ0mugsHJnwiNUgI
g2b05GgULsYwr+fPraPfTvD2Nd93apQlD0Xc/iUF997VmnRhqaUVgPing9ZomHYV
8M9EMv4k3SMg599ywZ0OmFsGD1H7FtO3eiUxA9AWzSQtffDYlG5h7BTYvBZfbR26
TBoK7ZBozYGH9IGFQh6gwATS9PF3/gwMuARJch95i2d7yR49iEPpCJMELsNpWUnX
SCDimNFeGM746iNfiC37+SAhWJ1u6TeltzUex+tDUXwNM7CN8DwgHJ07EBcFLplo
oLUyhz6aUh8yw5+ej3zQbJk80D0timoy6FTh6t6LLSakiq2juOEDpL4NwLz3BnO8
3pv6FMrlHrUKF928QuMOG3Hr1KrzzUwyCpnk/hiV10kTDPBd92zWZ0klHJ2erSSO
4UXG935QVSEyA0EVAy8DRgsEUkSFJNzjppmOY96ThGA3mH9pPwiP1OjtRyMP4Rlf
Lht79OjP3xY04N8UAF8KkDPNa8cWe98CBdQGZ56Gid9+dn+aMRiCUbl/NOcKGJi/
q+WoaZqFG8W+wqkYIZQd9MkuTw3evfOwr/oeE3Fv+pCvUubkDEk4eLelFvY4nBEV
5R2s1NAA0w6uVNjni6/21cqYzYkjjf5scCgE8QirVsCSodnjpyLBWm1JXpL75PY7
0s4wxA8gYJ5ha1yXOSSwt3DhF5F00/pLZBUJWzDC31cH1zP/7zN1deCpPohkNDrh
EcWWYO2fWOWnKm/MKk6daBNmmbYvRrf7LZ1Xuk0H+YBNErTIhOLVxAy+MfKwlwua
SCCF/tfDodoiEYQyLLvsAnvBx2/+QYSshch8SCGaMcMdb7QJJ+bph6GzLOaFLNnD
Cl6zcC5WYdeqFXCwSM0cLacBKg5htugC1Go7uAAP03twihJValPL8OMDbNE9n901
xxnXPYpIOcm8RvZDRBR9iB5GCipOApjciizPCbc3NAbQcFqz4MiMqyJum8/cXRqY
qwd0tyMKgA+c6a5vh61IbQv7zi7Ve6g1EySYbJR12C8go25/x/CFwng3LwFFSjrA
Y3ze9ryX0kjhBPTmXNN7Rxbo6gAwIQsA5ssATsaROMmb/t0lxcpMNvd71jbR9mSo
+CsD5fbGoRZ/+X3wsgrUK7B8ud4D/261hPq9EXMgtbShEGgXPrA3nB9vgrD2juf1
MCJhb7SmZNR4M7VNC2GVTjWbIAJeC6MP3OzOBUK7/knQNUD0na5z+ge5Or+CV52I
SI3ulJDX4tDXNpWNcclMm8M2JCBkbvkTSno5y+nGcXdFrPtVdx/1C5+4v+d/y8pG
XSOHJ7qQHLKPOsY+7ztUBPVk8qHzmbz4HqMMRWCuLCNizmi5ds3bxyIVl6N4iCdx
IKcNtR4f1YspwQ5yE0gVFhW90j1rXGdCwr6jAqygOHiHodmVyroUHyIAKPQ2A6fT
OHI6c+IdyweCmQ03fY8AUzWploAMwuayyJr1JOUP5WIjDVlCI1vDM23luG/SIRrt
HBIOHc2GarxLvyFeX/N7TfmtpyDLiBO68CGoY6PaSWfSwUD2C9ETF2AfgBKJu4O+
MK6Tj0COCSu/2GaoE0fP+Y74+QYuSt0r2etUqGQbtW6flAEDuybKdFzQGMqcKDTZ
/ZIFHn/iOwRRbSakQgxMRxQwHKzwRRg88Tkqn2Ia0QJeApExvZyggNWfTsfePCmk
RKtkKYVyFh+tkwMq6m1n0BuDdGOhK1Z+6I6ENze6YQAvzCGPCTx9f9WmIsMX+zX1
fSHa1t1C8CbSpSmvmtMkO7rKOJM+0iuIeOjiInMyP8CNR38XhLwNtfL7uEqlieMB
tlp8LCR8vcDUePPZK0nERj7KES+E7/L5d3d/GBJUA9sJVyVA8HBgt5IpbK6bEBxe
cDrnacCze3LVnV+KyR7+w7JIbSwoAbEaGNdK4iD5uxQ5ORZYcjeuz8g/FCnPgVzL
haRC5+8LbSBiKcmp1mnCZuc1jwl0JklfbiU6CWB1RMncALCiN8Fn6+7IVdUdqRiu
wEAPH6lhSOKjUTeiASDs+P2RBCIrAAnzpD3Lpfj7n7wg5VXqSS4ievY6ZTrVcygk
l2uRLuoUixaZ2ZXAb2OwUhH4rIkItq7GCCbwuyjT+vloJJL5haoOwHqVciyhhEGk
5bFxzUed32164ViX38gyJF9XsRKPXvWMUREMsLZVhLfTPgCW2f+HBTXDGVaEGdJ3
47SACARS+mnakQpdbgSD9+V3AGPtAW/M1uflQikVj2UnA8zcLLGapFnGrQjbZIqq
Oic8PknvoqnFCxdWWg0dtuhFNXHuOWMpFfxI4Od/d5FwuzOOFhjhMpwoF28J3bJ2
SnPJIxd1ptwNDnUAqt2iAvQUdxrn7WLE6LvuCHF1heAuk4E3XnUvAJuhSJV4Nsk1
k85871jKvt+zG2al4HqfIgLzHO16atPRCg+zeunfOI8Y8wDl3ulXlMdt4YBG1TxT
QEYTFCxoqUd/3gGOu2GcaDDZH+V7cooxyrWbNEMij28ExPHvEnoXz0vvJ23mguhV
VeFTGirJ0IoN5upk4LwgkyL47IQw2EWChiNXIKCX9IcGgtCPIFlhUNi+dBW3/K5L
cbReiX40wvz3MmhXP2JRqWSYHbERFjXtykRC+bxtFv8g6M0/sbiV42nq7kpSrEwg
1Lrs2vr1E4FXcmVvfBzrA6FpwJaoQUTWgJ4uMM3GnqAJpQTFUZA28CANrpkd4HqE
KsZ3+cN1C87gXUWyp88LoSkCWUiMSeNWtyPlG7AwEigMkXuHyyewJ2HDrIElM6Pl
JbWWjm4tAW9Yh3n7MxeYLfPYRrifRn9fbUwGNzno5d7SRGg7mizuG5fEtSTgbCPD
cXE1iLr2FATUtzgk3dhDX8wSvP0TUZhAI7yuU4ezFaWQ1qE+6uY/dreuWfO/FhQu
tjsUEJyyzijZQ8K5XwklX8vaXq354ihxbaQUGFeXmaZCdyFAv/rnREKgk7FKlwJX
7vQoe7RHqiKrfGRyTTlWjXtaDm5ZgKOGWE2OnYYgbiP1FVvvk1plthaGtCEWKYam
2jpRfpo8Oow359ScTPvDsrWgoOOOZ9X5pYMGT/VF9bt/gLkaa77m8ZwvGATd8Bae
9LLXL6WIkSEaDrLnmKExv5YyXTxXkKKpF6jN5qkN5RBi7Ij69+pHeeFtdthiUkLU
LF+jsN2LsiDQDht0HE0gQ6D2EaZ5rd292pBmX7n3DGDIFrut18x1Bq4NW72FeWCU
EwSvYWOK6QS6qulLVlOPCYScBho6KYL1SzoOYaHs8FbzaD6m+12XdXfLVRf101UM
/BGts2aH4xiWdETEZxPfJNRAP7wWYpGkju8+tFevd2ctW0I6kSm1tr8y+pGCMfTG
LpPIKf6wr28QU3frtAStV+KKHRz2V1nC7NztacEWI4bcWmVeyGoaRE9qU5t4G1Ft
XpDCCnwnTqY601NjPPKU4joRlu39IIJagIQf59hEb0d/K87dBkN47/ObDmhgFJTn
x7lQ1Pz2kqOltHJQfRtETEHXrHMeW8iYtwhLlpAtycCXlU3dnOpLZSnRz8dgGqla
Uf+uBeBioZL610T67GSqRNsnxbvujmy8cUi9Q6x8czVHctmxsGyDKdAg25IKgSrS
rvW3bv/G+mTf2bLRyW0qpRpLW0zuqg7iPIXEk4d9BXlAaQX1pU8OxX8+G5L/h5Lr
60KOhsf2juRkZBgBcwZICOWdV6TW5fkYgjcSsJxsznTGKY0VgRbNszNtmKZscb2I
ZiCXqvv1hCVRCn4nS4l99u3JZ3vz87oGDZ+39aOAsMPbTopHEfeTZDJJEZ8uewfE
p87CCZvT87JSaQJmVAIG2sZYgP0Q7YfbDOsym3JpbgQHnKVz53VyU9n4T+dvU5Ml
VFWsGnMNB6C9ObyfUlqDT+k311gKoQzMFt2VAaGLhUOGqvDhOXCMu6KFBi5clsI2
iDk9SuPg7j/N/qlnRddW/zBChbBFFbAN4ylAKBiD2BHgh85y8oHHVY9OSfTXJU6n
tSwIMtwe5mKOHT+EBUY+HljPDTRKrwzJH1LUhbdbellrPLY6YE5L6BFJBEhVKcN6
Vriiy3ZwsT0Zr6s0Vgh+EXb4alsbkpKL1EPlTqJdmfdme2YEn6+ZmqqhyHE70Zoz
svcRTbgvHa2uPtP0452B51W4N9NBmqKWzy9FA0/E2HU2NlsXQox5vzInpDkEc4Uv
Y+k54UqoVNrByQt1dh6iiRUwZN/79vgIt/8JqK/CmAV83XLuVMo+aS5E1WHiaqkZ
Ybj+fuBuQFYvxtPjclSvlYT+0o7w1a+pS7VJZYVH9gOEd8Gj2zcdSdjHgJDh+PS9
M+Xuu1dPxh0V45SkMEfQDKV5DU5nJkBJGuOOsXi8mKM4lPyvgHnz9HUvpaDyEZrM
4cAL3K92Y4dw29lJczsJ18qTq59TzznhEi2yDu1CnOqrKB7VcS4cDgxXK2ojC1xZ
JdnUmIeCaGqhutDuSQT2W+4G88iWEOHbsMP1hh7c7B3V/QFbe2dAfe/hArYfLkRb
fG+/ESU39KpZ5SqYodt/hf4PtCgPNBS7xKZAn/UXt3yirlFRsxf0NkwS5pxBr3As
FaTDqXuxsFQ/4L93U8xTxRfjatz8GwdLDAZN+IhdXLr+crpSRxTlRMZ6cMqQ9rZQ
E81JLK8WYEdH5ECqTK+Viih58igt6yyxtg0NUUyGFEC/FoHEtCoolZL5O4e50urM
wrbKHcZLWrcFKq0U4NXJpD0+oVTVSBRPQ7ojIZJjuVJDsjasO//O0x77O7r9OK+M
mslfE+7IvklJ374ARWTO3Zesl7D2CgGDnFzH/Wf1hWwKDdP593Vy5e4rEXVN7ap7
8e+kK2+nQb88mnvHRNw9B9A0ljUdl3P77jZqUpa3ObDkD5rh5/RZPlO8ShsonNmY
A7AAAEemmM+hKLV5zHI1FYe5dvKMiXt8PADPFY5hxvK3twtLVoXd/Yhv6jRI6ZmH
v2aioQAR8ZU72ejFpSUaqoVfYaCEq4rgNfu/FCez9QNsKT2UytTD/0Kw12FBkhQk
MemTtal0VvoLyY+hIEUiQo45Pu+97JHFhSmSnYk19hDp0kudAnFokkMWSjaV+KeF
MZTzE8y2HOn9/NG9imOj8snQ9HjOQ0Fbwe2W3oe0eg/c68WoPhoZ7np+nOylXHVR
BIIBCZkYfbiMLtwuGLWU6C3gPLQZpGGZEMq/v1aOGhs+C3vVcNoUTC5RBXGtGDSS
s89Q8/PZHv1YRRirpEpjcNXMsTNiLb0q9+uj6/akMDfESmvkVokxAE0Y3SkPaiM3
KhMp6MpO2spzxPPVUM0MrXk3wySnFZapra2p0yvrWHoOuDjutBqqmRcprYyk12N9
e7v/7Ko6pSiEZSzBoz0xgdic83sZY6n2eBgEEmA8sfLhm76YPNMFjIw2e7ybnymr
wILtrgejbFFWM+sjJuV0SmEyUthUtd7CfBnyJWidLLyfpAL8a7PW4ssgc/s/soNZ
2ua6oE1CPX/4j+AOTF18R/eO8oinbLDT+3MPTU1a2eN5eoeMK5O38lKw2pL881Ds
d3Gd+R+zb1/NEfb/oHpvwoKzXqSQp+hCSb3u1qYyKzcxV1JYT8bZfM5F3d+Ds1oz
Q0a8RIpcgqILJbS41cQC7Zz1FU/sfRelaafcphnaY8MGnHkmKgJj/G7yY5qWFeIN
XeJ+yUt/bNpfUWw1208GBFB2JiKIdzanT7hxrdGEjoDVRSJjU/J+LeDqtkcUW5+8
mWqyBSVwB+vufZHaNzc93Bub+c4uqbwZKRbqXlkc7L9kdW3EbaibDsDaiwHYTyxZ
eDh3ptJ6YKFVF/VP7Ir28EzcyhfJP4lLX4iK8oahe6yLlNlkcy+PGMzV3BkASw45
8eA07LUMA4aV1lcdtJeERUsa0YzUWu4BFw+KoYhmPnVe5k/lWt+lGOLQPjmrm/sI
W+cozlCau7WGOz5PV9JFCFe4MqKzb53RkGppWO8Ob8VMy4Bm3C3EO/FyTi4GucAj
j+7bUtxtd9NpOkJVuugjbisg6t1uWciYy7YZiI0HBzgeUsVlIzPTuDPNiB7erj8b
Ibn09ZU/5A6c/VA5XdVBy/n1WXbNVBez8VDsvefeh5OuWC4EpR+Plw2scV7Q2Czj
BL4jUhpzk6N5zw49CrPW4BuS3kdi4HicTdYmKNu3bxHEyo9Gbzgslwu2/W/hTrw8
36wEzHgedIOOKKid4QAfqY1ouxdIHhd9aZbsIj7dUnTw3gWDUKg6qe8TspEktXBy
6K7H2QxzDVkLPN9bwSDmCbeiZRVRubVoMrArQBjyA+ucB8kcvhytvMyUfR6WZXwl
OwmYZvkU4QoohFXLXQkZZAPckNz00dxMpCUv2mPxUCxuMEwIx/Kh64HlGApr+G+a
369QoXxzPQ6RUuknf8BcH18+za9PWGmNpSOtCypQjfKILAbUyzaftby7T03qojFM
iCxX5iWABMaoYJezY1+/5L+C1RTgVaojnxBA6sQ/SColUNJAoNDC0ZvXZKZGQ6bW
Lo0PRCKsqdb4vrr++RgpCQFVRvx4BwJQByg68FBLAs4j6LyCKOeWOz6HiqLNmz9V
vP1ceXhmtdyvHAET7YlB+Dt3Y1OklH6fN/wmbsWzJdyVz/XjIx6Uudfd/O8mUueF
dhg4VCj2tAjsYA1u9sbK0d/Ro2N2/CVIqCebJxNJO2pbxIsnmWvkKSxlcBbTpI1m
OSt9GEsz9oH8+kh/VdTk3i3oVd3cON3+qSQ3mTlF6FsHVr01CDDPdBhqnsDuvPq0
O0vSqn88PDYTF0bqII061sS77aGjilSscy/t3xY/78fHexkt7vNUuhJ5X+v4CTDh
5dOnXEdh2+9HQL0DH0GjFcAb3Iu+HVrf+kisHuGpJI0dRASvSLE3e2F6vaukbvIH
TUpZWiKNAl167cjvtaFyEkU4H4twKDsRp11vZqfqP/oPxzVhLrjMy8KoLwE9gRjA
NxsaNvBlAoqzuUFkkuR5tFMhbHlBq+fZ3ArDDSDaxa99BaPRnCA2zyXBQZqQ7Cyq
i/4PNBf35ImkXofIT5q4wvPrrbmsndxFGmXT1GoZTRHcfgVKTmb6kpSlKLcgripx
XtkpzF11gYfGEEPD7zAB/o7EYRQx1wynFFkh1ub34lGvxRrTrsNQ9FgkdtnRf1TK
A9Ih3jdAF9iE3mGxlVe3OQC4qgocJdsyyswmmzpoH/d77yKU8cq1Nm56xTMk3YPB
a/lP2R+iPeWTFYAQSz4igben0JCeqxuVPfAmOK/dgsTzM8iuPOsHPXk2W8c9+yqB
YchQUeNAVvCHgwvXmUkrCw8FgajTUDfs1awXCC9C9Mwn/w05vkRE8UxPn/5gIie1
kItynaYGa4UKpolm+Ce9lfQEkKgO8MFG6aZ9ju1xhQepJTytwPBQgP8etneoMcna
nh4g6O5yHtdLfi35BarK2GGetA/ucksL5ibIywxiITBAq0UxtBEe78n/qGe6WWxc
ECDC1Art1GFqo7iiyO0CcKT99vQc7FpYDCVR+MS5UgvuC5+mt+5w2A8co0GPiEK5
FoKL5ktsSa/zDG412EEdNkYCUACUtkK8hu1mjAbOnMtD0pABeV96WRsjjdoAt6Sb
UNKltr2j99f8NymCailv+UumGbpOA/DxbXpeml55KgWe06Oh5g4UvVFQ9zsu99Vo
9bZs/CRU3EpFIf/uxt4aFpqlzwih+KuLrqTYPkq34eQXomc6rERzQWrYe67udgg8
dl4d7d3MAJpwhEi7xddWOpxJCwTnnsBBAzpjT3rhZN59yXAElrrWPpY4wAKBmr4q
PQFjHRjOzlTMrRnAva2tL5qEgCcy73eW4vjHq6VHAocZRltaLVlzd7P8lO731Tfy
9uM4OFnhL2IJRZUofQZ7t5fo3o9B+eZxNVkm/iLMNfG8SD+iZsqvjSkdR1JyT3kV
6X0n15F0BeBnQffO4nsbU6+LaIY8w2e6KCCcShKks/xXRKo3S2Gbnhv6uDYpK6dG
A3Q2YFlCbfx1gr/XrZSN5arhy5d/BFAKWOENNeAd0/WTBAj5ZrZ0SyYX7blwuj8e
pVnsYpIHjbLxvzhua0vulmmjZBYJp1nUsLB9KFvbI8/XdhXk1S46Pkh2CGcIZNVr
TPDkgg+ok8liFWvHAW9OkiUUOW1kSAaY5Ido551oJIyldyuk8xFPHLeAvZ3M1Rl5
nW9TZVI3Z620t2gJolSTTYmYP/+z0PW8AfY1Kj2xAdkc0f/J4tSoGB+CanQX5+j0
mi70ifoOR5WCpaird2S4z+e9kXYiN3qPFp8TOi+FLA2RYdKP4CqR8AFndu0Vi+6c
/YEgzxpS4BIS4dg2gu0plv/cgSw7hC+4KF8jA1UD3P1y1arBJkE7eN5kOyDZzapg
QYoW5xjAxxoUliBsWk7xAmzsu5GEjJBL6ABMOGWtZVt8Z0kG5VGp85Jj9vZsMTRv
mmTnh15e7P5FYkhn5TtDzDHV6QI/+mxHg3ejXBh+XtB5HuBXYeatregb485r/Cpb
khx/AY4IqLR94I8Rc4DPhBaEONvVZ7VAjBz8l1R4lLfDt4OSGkOX04irWwc6K3UL
2w/TUks4AfXmV91M6FkvViQZwiYDLaf1HvyQBpZLU6eZM4IVR/R2efsCjNQKbUSX
wd/q464ybOeV8yCMzmanQouqj5yTmkwVFfMHBE2eTqzLta1S+b0yr1VtvT1f5u9b
1O2GVerqJW5KNHpFHg+8AVrQNPzcMmcqnFeY/uVBWK05tLna74Rsjfutp+B+QB3k
aNE7ntGOOguDsbc5o9qpKO5K6n2SlvHLqAez6ZWnQ0tZDDHlTeB3rUIDEVDAbNKR
SCClpoz3mOvQAgJX4Zsau6B8ukd2M8ygLylT0hYhoVTT/EB7YUrMZ6vDr7YPXUJq
fh0non9yvnjztaENOhO3J8jtNguF38GrspyO7DdwkwejFW0JxV9NKfZSK2Wd3mIu
mIPK1x6qq+mJMLXFv1mYWfNFspP5OWCIKC4WsbKLQaLi2Kmks8nYCuAkKRI5Mmx/
F0MNBoY4lRWNGNUXmvijgKWHTb0LPP+LxSIrR1WyFqKbFN8rXBd+vbM4xmBewXxA
/I+Npv4cDyQPrliYdOmL0LbyqWLhn28T9/dTt6OeifacY4C5oxYOpvt79Q2eRBAn
9jANE3uaG+6gflxllB61C/S8PZJ5Y2hbF1mnplJ2tZZFaN34HqJoRNRGAWqPl0zh
yPYeV2D7MKf9zomTMK1SUIjGbieFv5uZBNdsClIJ6nkY/z0iDvRK7u4wagJc3Oez
HLH1YLRnFLkBHVj5SqN/NSnU9ljMMeujPQpYmXslYyBzJ6U3M6rnaETLiWIrlg7I
A63hYnHfSPtmZSL6J39q+T5Y3ek1XQ3tPcuBwk7X217EfxjCfrcVQ8xPhMbxzRLb
VPwr85N2OjkAW5GmYPexOeaaQxUneplbYtyNhDWpqigDgCxh4odg+0tRk1EXLZt7
c8dxHadmub3LPk69q5dNqKjO41hP6QOrT7475YZTYIBRH5y+B5VKnXasCAj27fz0
dy01r6ZaHK8/BnPe0j9FjDL6DtZMsnL1kRTt9Xq06HGcycLd00+LCcDER6uBxveQ
wqOFa3IgT706Kl1VbyKMQEXWstAL8wDcIDHP8GsstOZfueDK+X4o4yU0/nZCoT9T
3m9cQT3rKODqtO47bWYaXGERd3tL2t6Wbk6F2Y2t5gpjhYRQ5bwCNodOcuD+x8Po
r/Bcsz7QyC7eKhz8dTQ/IApfR9nDhfgO83RkTwpvdAbW9WeeeAPQWjzjU4Oaxud8
CG1ktSpUnn9oVAwVLCw94DS2zt0dZZ/IW6Qi7jTbLcrE3z8Z37yfirGhK9A1pqdv
VUi3uQud4byC/Ua6xqY0C5uKVyqZNEVba90zbACKk3//nf01oIMWlmL1nCxx4h+c
wi+W2uG870CEb/rmzJEb9Gh+PtsZ0DJB3xwldqZD+4qMocVkocqQbYv1Iyvg5zBi
t2JlhJ13f4cIBTAWoWIer9ZIsmf05i2SGe+IGl2E9sIwSG+RSiRzycS4UxGS7RY4
66O1kFU3+R2FSwFXUdboyqzNZqgFRH20dLqY+Mg+vSTnWNcurG2VLFOaymVW+0i2
UWxZYGRrl3jLdoUdUwAEG6xaKyjkAcWAA8eMzxUNj6DFHfSoAeahh7Sh3Yewa1xe
MDK+TYP3dsTeBkLLJaMlJgtgfO5pqjQFwzMnplJNdKemibtqiDNeuFEgNb+aDTT/
6Rvk2BGbynz9QFOnXM6k5Wgl4t2/uECNBC5cM/RxUq2CP7ah5TCJiOi2+8Gd5A6z
+2vlPE2Oc0mfpt2tsi03nnSD9iBTR7rtfGVN8y33OafooT77Ano6XeBxg39GZvO6
olr73XB9k/AbE7qBVUP2Ob1mqjfidQ0Js3u/75V7gxl+tx1QmS/dmfZHHzCqLvKl
m2bMZci14k6/8M7unosTkSh/jSmtf0JQvolnGkZICRExvlQDGnMdMME04Vz2Uc9U
SSCEzdJcznQh+pqSfypGZtfQVZ31WX233VUQSgOMmiY6SdFzke3giMk3TXNCztDP
uxyk07Xyfmw3Vwx4u3AcyXB8nR4FXcVOSf0sPKKZgrkPKAprxNdDaUjk9IgcM5T0
8YZgRnCYQP5q1nqfC0X+355RQm39WEo1FO3dR4UbSvctSreu/HsWkCcvWI8fcO0t
AtSQEZ4aN7O97QYKJyOmrA1Gw8174tq2eYv4DQZgTqELaedaPQ5WAXKq6da2WrYR
xdS4dsnkRqulFUtEaQPF5Llup2KjM6X3QRnL4HdQVgQQvRQOVit8cMrZ2lAd/sqM
9Kck/gg8JEgj32BW43NlWQsFTUL5dr8CR8tIFQ91f/9FejFnQJeNdKOSVZgA47bN
ji7WYYF2cdUxEMjG25Kt8/rqAiReMQMwxpHolbIr0xz6/ojh/kJO7BPg4D0QqMYa
J6SHLy7Y8nY5eGp7HA6T6QaSudEznKHmxyy35qNlMaZXLcrZEqWIKS6IoOl+uge9
3vKz1bJn6AtPuuVFnabY5nxlJ4OACh313tM7cX+4SlMvgsIt03Cv4ahM15ULgvmA
VGbCdwcrQNVVB+LoXKbjvEej5fru8AjwP61Nk8ytiRDPE4KXZJVlYvD6bHcQTc9k
0BaUDvaxwx64l97Vs230niIHCIfDm7+P1vcLcTr+kZqHnANuSuA/vc+1xaLtDfaR
bw2oXc5cCTxHPKvfvSzNGw0+0Ke5exiFgxCEe7C9xHnqKqS/1HJSZN8ib/Xe7wfb
478ZyxIuxluSW7FPXZpVO68unKxjw4A6XBFJzaarfXUyE8po09+41G2ZyAboL0CY
kD22nb08tUwIqhY8qRAQaj2g6JaigwRYOUb9V78YE4mnvvRUWJoVDsVZqJV/35Tb
Z240JK5fFk+slU1ZufiKOuZ3T8MOhrKNWQEGN77dH+04fg9cbHFo+qNVOMh/CX1U
ERKQQr18Vf8kGpnXJVVy5sec/iQJe2qDqMh3VYhtVecnZ1g3InM4PpX1Gtjh9a58
OUiskFQuym92aNQCLxyUns8Yi+k52MMzfyMAmSDdBzEuz+sgm6vkVL9sGN/HV1Bj
jj09RxC5GE0kM3YgMqh8dS+pH3NkWF5ERZ6rmC/E1VzTMLKm71++hv4vkjEesoN6
zQN+MQSgBo0k5UeNHiDatx2H43qDIjMkTHOhvGKgfiiOzXsyTWe92ov/eAm8FPSU
1HGdZ22kkr1UQEO7hm+y80bgeyRe9q16ByhPCxwvIEOJPCAWmPFhstS27yrGldS4
HY36AXmkjnb/4LrXF5iEHFbV/DSZ7VBETcLiEMiXYs/6rSTc/revuXv2Tvr0JVW2
Fc/IUzmTUPUxS9k3bJyueniSaoEREVz5tSGspc1wjUDBJjYVj/sY+nPGw9fj0YxB
DX/xqlEr8NFcmqaV0hUydHoDySTrdKIyguKRhpk7sZsx3pT5iqkyds+cU1huCKNf
h6AZo3BE45Taf40NBewCEcMe74wlyVZ0IlQ3dhuvTZfM9oe8dB3k5HPfWvqxNRJe
4TzERwSeeqgIEY6LmOPRg/0oA1CrsdYjsS5miMtylZoISD/2Kn6I7bTTvUtFUnpU
xLnympOHkbcipcsLvgTWdOs5EYu86oxN0lWL5De4XFEtBdNemNzeIT1FbgOHI3Yu
1McxmZ7Us30wD8UZM81PVTX9yViQ5gGPwHqgUchg2vv+2SoQ6pgr12LDj1RdHYy7
Eq5sCd4kpIzYRwdI6br4m1iwhDYwQTEdWGH8Ax8Oy304kOfrbnz2BoeTWLYwJrZ1
CwYYoFiUeY6eRc/sfurscOLnrRKsWH8AiJpv1B+p0r3lryCuHunDtbpsQq4jnIW6
HYADzGmg+ESUTQ49rVwuLHnXSSq3hKNcPHJlXcRPWvUr8Y0dJ1HpNkH1nQwpLCvs
S+t7meOfDDpbq2ZaTGB+PXZUnX3F7UVpYRtsJPh022r8J7/E7s8VRLBhY6RoLJC0
wMcdWzLx61cDx/RhoGF8L9VFpai1bQpCJa1jPFEaJYmqeFnB15AbEk+Y14Pwn1+I
FycOi8bcUNmJ1u0aIBs+E/BmXG2Kw+YE2ITdbamdmyd1scAccYM/I2naTCxkm+t0
W8ueoQvBlQ78ZN9UsWV/EFEU9nG4FWxXmCBcQT6SjUr104WnTmHW48jRiPmTij/H
8lE4wL0+XkyMWTTeA0bG13Js0f8z2y6NvopQyc/cKUJK8qOwXDfog0r7TrNz24R6
h6J5VnacfVazuqvHj3xUX84feSCFhYlmVjeTVQS3VYN8I5wi5attQjVmfhud2Olw
9tL6CcSKyzLWAkZ1rKyPaOC5P43t56AlYAykdTdTO8Z1aBVcOIHLLiVjQoNPmbLX
/oyvkT5hY2A0NuamBHI3tI7Fnikeck/Dyo+HBeaMJB857cLITi2eiNfa43m9xtNF
nEiwYOy5p4IEjJAtog7oiSGSR0MsYFBKR8DM6OFyeq2iQ6Gsnj+KpSon29rxiR9J
BGyQZv/kwBVkIy9++xlBLvwsOpjA/a4d7Nfcj1nswEBlHgj5tYr9UQ8LzW3sSP3K
zVpCT9XOU4EWbxuGSblb+bJijOx2Pg27nRTW2H6dTgV2+YGpcNi2+IScgpEAMMzL
Hl9qgSvYUUUYjNLrbk/IaRI5acHulLoGKfOyXaJsSKeriVSfHd3YvTs+MPJBssF4
w91UJQoPLki9SLcLxGf0MQIMbXqASVPQWGyX3+ethNPvWul3sinvQ4+IhJ8WdFSq
Sj5O9wdPvg0EPylhwFLnt5/uW3UYWEHsgrFv5F9ohrZsJZSpvxiKD0TewLbX7HXg
G/vO0fkElQPHUyxPgepVPxmXFq6M1bVZfdQpSBzWQIIo4lhsJsuxAToQmQdooZ5j
+mnU8JbWCth+esjrXXsntY+VRe8x4OL6vYVqqV34LEKyKRKTcyvty4u1CDU6XPf2
5+a3SLrE6n5IUGi0+faTFuyolKN0zaSyjJoO8qjUK92e15SNRi+f9vgdR34f3UDc
QPQ1LVAdB2WeFv9KUM0Fhf/2d5Xxo8U4UuETKDKC51A4/aj9weJkhZm1WmdXUZyk
FSAyUJJ75pWgGZqfzkSULkoka4xbZsGJxj7b56/g7WJnKDo3QTV1+fV4dHh72bX1
tZeRy/f1dUhVRM77IR5xnzyC4hK27QiGE1ehG/LVtxCq9Wm4YPFGGsoooakROmoo
I90/M+tvjlZ4ADLYlCbGL8TS1yQFknuT7BbsFr2InyE=
`protect end_protected