`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
<<<<<<< HEAD
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
=======
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
>>>>>>> main
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
<<<<<<< HEAD
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4064 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15k/jmI2z0449QtUpJ+nFFMh
2RRqU7/KtH9oW7ik7WZEhEKTrnCeG4xkMEw/N/RzQ9W16DdSXUIUKKcjLilui7Vs
jsXabOtclWtLwId4zT4mws3r440Ab+NhQCCxnr5OMsITtB0qWQxVV1iwxd51oQXW
HWk784FiivKqfE/N++DVSbF77mN/HzmzWuZUACgWw+Opj3XtqagIpbHc/WqDYQ5G
/AicD2PpHLWyHOmvrqBZrILKUQ42Bca/8EGKKc9iqj0/DdGT7wYZuSknueuoS1Jl
mXssW34+mvsR561UVxiygirqmA40XuDhnv/DePkH2t5Bhjd5+NW64O6igeE40gQ+
3Xa6fIIosOwEiziYXOu59xOXNLEtOXqt9Ey91+ABM91evsNUP+WGNJt7fzveDp54
7bt19/U9jkJJVF76ZkukulSOqpHOWyhyfpZUwK/UUYxyOwJVQSalsMWN3kcXOHjS
dC6g+S1VqHz2YrtDtZUXjX7XFgnTI/+d7po5+A3B3pkjnf4vUb5OnmBSJsbxYeDI
6LoPOwfGdiNyZXQg9VrTI52zKIoGDL6Cmtljc0ZCrZLb5574R4VLwPEAt7YatjjS
A3fKQaARSPnJ0G0dnlm8VTJuyIvi56CQUTaGCOEcF/4HZLwIhwt/iOX0vvZjkad3
GltQWM6V8mk/MgrjljADWd+VzZOlLP4BzaJKJIbPzINkR7kUponm6q9ICwLRzqAv
4CeUEUpNzl+6wlrKAT6xhw3mFmnsU8tjXUUi0dfaTpfcq4NAK2kl73EoHlGTT3Q/
fxsDdVOTKrpv6O/JaibXM+C0zBEsFFZT/u87CPbGkTHV0K5KqTScl/5ICRbRUzN7
BXjIM6FhN4TbhJBy3rf/xxEqjRg14uSYpFBPSukMExiEaHQyTLhflFaD4LY6hgTm
X99kf0D8cdAOJOFJcr0BPs1szj1SV6bEYQRkH4ZIIoNIK13iSKc6fQb2s4nnOKJX
9OvqBvtoxIpQNSAYP8Yl0e3SC4lO1FPVYpOhr9vJ/+fA1D+ELObzpjIN1cXw+KBo
8tuuPdQaShw7EBMUiaIdmoIJO8zDMjH2kg5xlQBa75KEWYxqgsF+L9DrkdZT6O/s
ALBDxAhGXbNjnic1oXBbagUrVe2FjymO3zPH8YQdwTh1P9DwNoKdZOkQJkzIZIm0
zGEE6Fg8rOfETZsQ+UHS98h2WdzXTJihFNyFQlKNK5KpkpOg4E/bxfXkdd+19A1h
FIwb0goWun+ZryZ2tFYdEWBJjDKLqwIKOk0+4CT9s10PTUDLjMNqi7NEdRKO6wYN
XNwfRSfqN6rgPf4cgc+3EgmaVZKjStfqAtqkinBot/GCBqLSR9y1XM3HXDWgYgez
naG3LIbG2sIzYHpVFuurpOM9yLduJAeau1sPe32Idhj9AQ1JfD9u/SxFSH+PIlEU
L9rO+9AnNhIq3bybnZ0vqEKs0kB2udB14NnNdu1hr66h5TLs1YNBQKvpDN6S0wL7
6PCuOwRwzB0XMS89XyKu+tQGJyVA3SG9EETh053HGAQ80Ch+gNrJ1ApkLZgKYYjv
Qh1uzB/bHu3zmqxAMXX/XMzqAOVIXJqRuefvchtVQOodh+CmtBVqqBUoH3Ywurdt
e3h3L8fws5sPA7LStG0jTaoUFQE45kztVGoAsL1TYrxea0K27nyzu6wouJgp3NEA
UIvzVgFsWNarDWw1ZChLaw4eb1PTmsnI4uoT2zE+rNslKwGLl5V9sYHQxPbVMgh4
Jhk3xkoVX4KCU9W0v5o3lo4m5Gpz7zt4Bak3fs4k+rMD2Fwh1d8YEVhtlkm1oAkQ
NG17WvDlhwLS1GbN9n8eDk6T1gUOntozwmgPgvz0G+nIqBjPGS5WraI/NUjfCksG
zY+pOBfOrYOlg1gdPK+nsevVTbCZgXzfmM22fuHsy8CQVYpv79rkkYgnH8Yw3l3k
lpwZxokmRYsOu21wp2y5heuI8ckDw8mYX/1FrMRLIfiTPPy4/fBCrCWynwAdVYRI
IbJ4mj5tHgUVwiGhSN50EMxy9da+RWgkd3mYT04yQAN77gTkicqU5gfTonpiNFR2
1SoVkkCnQQHr6prQbMtT/IPRjIu6nQINnULt7fYllkZ64m07ct3FpTmYBsWAfnK2
FRRYgh322uFYwb8vAy+VSJrIC0rnjkhVx4342PEPJJyjVehbAOZivYT0JU2j6B8m
zsVEt2at9sxZVxOMJEicEx7yEjxSbcvWKNTa8E1dDBlHcA5h3u1gXUcf/Hcqm/fj
nhG/nt+V7RIYXsf7hzwCfy7HDAtRk41PCN4Uwzak1yClixfLKIGuUIFscev5aSEt
S8a93xDvWIz+uwzbXBtgwJFGQ9gnBddiB5nJkD8JfLrqWl1iB0IkAIbSjzjg77oI
SsNwIbabAp9YmbvALxOzPAxVnCsIUqdHc70FfZgPt9pW7zdAUS2UPsKZLluyxKK5
DI2PjkIENQKUThryTX6A4iLqojkJgYzS9vxkmnJBSX2WFzQxmsN4ZpCxHYvu3/bK
N3eegBi3k7GYpwHvO7r9Hj073Vnmswq0+L7iRsJfhRQnP6FK0myiOXgkXS35zQe5
oqqtKLHRnuj5F3BY1WG/Opmatzu7Hvz02pEnK9BU5OnHwmMLv2+gC9LETOKTzwHO
XgKB3TtvP0ljqYNrUVtWHF2uhhO/1Ef57U179H9CoPM0ulDzQw4O0J0Rns7Il6Y9
Z4Vb3+21acmUv9imb7AiCsBuMZ7SUvJdkR9+UcYa+/t2gdyOdviKYTULNK4S8Q7K
rM9EWDy8gDpbWo/8YeMrgcWDuZQ92GXqYrEH6GBg46mUrSDukrY1IJBTggu83EiQ
yAAdYjjhIhI+B1YBGWH+luxRK0es0TaSmJ4tDSMUmVmfQuAkZd2gLmhV/15GqOJv
sEwj9OM3uqjjBhzVqh9U5ZdSV/lTppDfjrK01BmRlXQDjkkl+fKoqzLXL1N1dUE6
aCAyPmR+6+g5loWjQne3cDc3w2qleJw1uZqol5ZCFhf0ShkQEAI6r2R7Uys+0lgG
gHNFgGWKehZ4WTfrXgf+tF5dzQO45qvSfNo3TrOUG6s9Bo+7Y20GkaNrp8mWYVce
44uF7KMF8YjE54+lgYFgdNCFXhyW1ANODan6ATGmjUVXfqiEP6mUePK9/9kHskdM
vk6ULVR5AV7fGgxWoXWlMM5Iv5U44z3U/EhXMPKSBPofzbepceGgRVlAnVkpICyw
RSCcYJal111TsbHkuz3lMwtcP0vPDz0ZdmkA1pIxfYr/OI4EY/IqXTOFrHz/rbjq
hfoCYVLaSfbPtG0f3ex2jegf/FwXuB/BBt1P7ZsKROz3U4JsEcULBJ5yfXYyvLP+
h2KiGDuAmumrdXtPjQHEup6yBv1X5iyYeRR4jDbkZmGV016dY6NOOwHmwDtAOyew
PazavW9aBVzxMvJeHbuCZMKtKi63p+YE8RvlNhDh3PiKTY3C71iakJN1AccJJv7H
rQp9pynuile0caen4b1T9exOOq10rzinPM0QSO+GAhJ0g/H9WN+ncfCqXcSCwukp
dpU3xcALVhTjCtOcAdpTNcZd8pez+bf/EPF7feWxrMuRdE4IM/A9ayfHvO1dvbSx
RRuZCajUmZxGmA5TyV8tUZpbdA8WtGgLuZioBZArS2e0dOKLDHFmxRii7rSt8vpN
viQn5epc/hFvU488awlKSNf2hYrhorbDx3wXuf3dL7KrHQ1yPpHzL+iFqN7gRoGf
jEip4zjEPQxZXTATgr+519LQT8ngLlH9O8DlbD7D9lDhk+3I2uEgZ3REo93r2kBO
c7S1HvKVOSMf9/r+0Daa6NlVZE1vR94IPMY6rx4NilAEA9epn7FFqQLCc6d3aruS
f5Hpna8HYzglvUBu1GWZJoyu73VH2MZM3jZB4U3h0J89RbsNyslZYq+OcCtKRQBw
6q8VaZg8nkEfx4xvLmKX48JeXjhf0h1/Mgkavo6Una674avisf8pOFWC3BN6JYsz
iKqHip27MdmKUOc8KdrO2SuCGTrzY8fRKIuhuOGw3SMyFDk+7/kWOI/3uISLsP9x
W21Kk7wkynwKp6+D5IIdNbpHBHOuHj42GkCY2z6b7a5kOgS9qToaY2wo2bR1Zx29
1Dbwa4qrA6/kozgnDpg5Nv3O1KuJdAywrpW2cWIx9qYNGpLOLFtMU1IfMODKDBPP
VlhQP7adRpE3XM271QAfiJz2fQXdNzWlzih3hM+aAjELRTkfQyqA897IddzB5Xc+
BkADuvwDgycwtUi/47vh8YqVx5jueptJZk9g+hG4kWs0IhnhU/mvE+y2UGhkPky6
DgdY8YTt34MmGk3JQYCobuO5pf5AquuWLph0K0q49unzTAkP3ReEXTT+ydzdyF69
ssTRkSJPUX8sUT0OFOFqQ7z8iOPdQ0f+CVsfRl7Pz6tS/I5sB5RzbLbEWBVK3BKp
/dHRQbybD4JoOvpX1qNwhJgc4jDD3zKa6A93nkvRIhu7Ezn2MfECaMzJGg4tWHMi
r0yPTSlBwFkpuF4GNzwP3jwEz6SOhKQiPTlj/qhj2Wh6/tcQ3cggX59d5yv8pCnU
yG/bNMOhGOXYEA4cOgEN9SDS3HP8la8nXzOAeCI32LcF9ES6J/aOOyXq0BuSS+V1
1NuWRoawx2N7xwuHnUt7l1g+i/fJHlAIfQ3dQjLo2Tw//mhgZyj2W5Z9OEIc5YnB
WS5RWQ0iC0dPlQqu0WolzhJmazxsHyJNVkLGa6h3y1Y+g6l9yhBn7ApxWLb/Kqt8
uSeZWa05YI0HICKLnRLoxlq11sWXZDyr12KlHZGjkvGjErP3enA+SsAf9DeCvpF5
xMCy5QZ9YNQYPcaUPjOcKVqvQxhgDadNWLpAkRt5uPfP5oeRhsQ2/H3yjv/pRtgV
QUiQbRhJO5Gv7vKMDooCulyd7C5VmITIsva+tyEe50y+QR+1tIWwA2llQiTeGL+l
J3XBa7tu8+kvHMn8Oo+0KtlDdoqKnJpOFSTe8oXgumU/CU+2aIQX6V7ojIMuXNWz
aOA3T1nGCAZy4/ij/s+lJxrQzd1FgdbGo5X1irWUYDqNda5qYBShehPlfyNDoyS3
p/YWYCCwix0dp9WN6lVxyi7khkA7FwLk/IQDKd2RL6AYQM/A03oszHUqJkaoGlTX
tfdWP6HkJ2N8LHvbKYdbfZatgG+htvzmDIFiB753VnqlClvKTxST5RO+whllj8kC
P0bpho4bUPN6L3AnAKZcWN8mKS0nb2HvAjWkeTEv2S38QymZCA/JJTUwq8kNPenO
f4QnMr/J/GCZ155orAeSN7MSyS+/tHVyyaEkIlDGWYE=
=======
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4064 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/T97rZhQva68T7JOm4bkq25
b4BW57ADAHEm2yg/VzsflzeHcVMMVx2VIScQn0AqTq88OWJ1c1KbZ8ue0lorvhkf
VElvHC1W3Vnwi13ARBqr2/lk5MD+uywjvWGv7sZRUWPJKpFQuCQHWYLM0FpD6raH
lAECJqk02ehZOMzGVDYZioJC3CYcIe/Ipzz7fCkUQ/8ZSbe038bbh57103GykxIp
jG5wQ79pDLPuQmsgt0ivttOK7Piom/WVoZgOw9L8L1YCRa0PerYSeX+3tjm893+G
DckuRGPiZvWPyAGi3JZt5svRkNZDZA9f+l82LJytG4wCxHMShFbbuhXGaQc4Xakt
vKdfDNKCLpyYAdZlYVuYtapVXrsABIOXFajY28wqvza2yzVz/qeq56ZbXmVNSgI+
u6rByhcGkgPsZhVfBSzy7juFbEwetqIvmLg9a5rFe8t0gveUYe4k0RL9ATlFONfd
TPeWhNQfoSRpUs3ki55M6VwTz5txCiQczKe3tyyIWFpFpQq/4BwmUAtaeHwXjvvu
Yy1wG65rglNvqQKs+I8f58+Vi7PDDSRfT8w+rqYPLTVDNULl7sWpVQuVD5TdLv+J
AbN/bCl8OSfNdzNCyk01j14xbeWoZnxj/qrgtpSdmv3d7CSREM8kK25GozMF2alw
zwdptagRFjjEH25EhMqE6Yu0ZiiwKmBn5a0rKqYPRYkb0s8vc+nW1LYrj5JXaGns
nQgulsC3Syt8t/3qHqmNEw063ZYgboLiy855t6qLQu9F8+dQ61xWLULdRELZXMSw
axSo9oZrJfRDFeJq2L8RXldM9jxuasxg8eeNDGn7EmPcgb1E/bwId4fWnl3Ke0I8
n0fkg9berxJ0MxcRcVwIfIqas8D3EktB8kkVt/3n9JDx39R/cOfSmxc2FeIkLUId
cU1sdCzXZQ4DmYdttgP8AYuN32tSIbDbuc1rYzE4Dv1NRiyXQuBTZpP56gj1Tscg
KvUIJ0+a9Eq0/Lfxx2SgDkC4SgVp508dTeuUizwcYFET+fC1pv2HFXlRhhrAPtdi
XKRE5wO2zKL6ngoqfZEJtf8+Su+cT3UboqAq1wMjtS3nu8w2qzatvJbgVBJWs/PL
NDqztQxntE2tAl3u0h+AQCioZBT808dOPAWKvSe2HTUdSlwUDUrfKNS1XsyJUr8p
juUCkfh3QgmL0+aEjPA4lJV0NVZ77Vm9W8K0tnS6OvlovI35k6dmFwrUqsqYxyjN
z1xTywIzfZ1rXayse9HWuOVoDChw0DWvCu/J9CktvLGNJE6lfrgYW7IYSCu2+JYO
CPb8ExGddXVhg4JaxmszsclDhJUeThjvXj/8wxOm6x6N7LEEKCUgV6pEncXQJuo9
Bx4At8ZVlfKtuHpBUJ7xAhCciwJvw6ETtXOdIzG0SUoDKbjVXZtTrW2JV5MIiPzE
tUaNXNS9X+OhqdenMukbfntlpI7EcOhpa+OZxnktJGLTHDastSpImL/Xd+V+GjKP
Bg7v43irrm0hnthAGOXYdRBOswBfE1MIdKC8gAntXwoTmloDZAyiG3ywaPUGhabG
lufvyFrN2rtsugRctdVYYwNBwuiZOMyq420xMyEwAUhenpXWcRoQT+5QGZzWlTsG
4kKJZRCD5deMhG7k/8pq6fIiWpwwYFDRERXBjww9yN5P+I72455c6UXw0e/9jd3V
eJHQ/lAV1zsuunlrilUcuwq8ZvmF47grjq0cvnaDcjLxBexb7r9e9bnvYMlP5T5v
Oa31/UL4BORD5UJuNEuST2z6Eirdn3tfqfp9wVGRl2NttW3o+ScbA53JOuHJWtMc
/VSfvMpvmU9fH1Wfha8etoZj5LZTfBOwsTziirQAHfAlOyYDK8cOdjWJqRXytYEj
XYzEJ8sd6N8u1euGhH0vvDXR/7xY2BoCFvQLdL5SOozTgysmG5/Jir/cP/vTpSu2
19rzYIugIVSo83jf8dKY/tdVOFP1m4uHzTHwDYJgY47tAWoV5Bbeu7ft0pCdbdhx
7VPSndTYTUqytih9AWndr6yvneaaV2Ht5+tMNihVm6VaOi+eC46wEXBdk+f8voxB
XZ8G4g7YWGYfRFwVv8UI+1e21T8+R041wmnIWs433p5tjGZOnSADumfL1nQMGZIv
V9RCWIS2Y+Jt4mMvwJxMFCLABh05ZINmE2PNo0QaWn6oN7OT3ZhvHNIE4ivYOipo
wzEwHhgcDhR+m0rYTX8H+VPj/BKf5PUiaP0+ydggxP8T1dwMRRrcoscA0Q0qMCEj
ZKH+YKr8C8vFAO0UAVzJvRZcSj89x9lr5sq72GdHYb1ay0n+57YuW19Fkq33uiUp
xcEQgudDWZNz3Couq47KHOiQQNr9L05kncbpNWEd/weAExX1yBwyO63zjtsBQm1T
xWmv1t3OK612m2t1GsR7FXAON0EPT5qWlGMODjpMmUkfZ15+zV9CPV3RMym/29gT
1cJs6N1PX9RE/4LnyS0uiWyx8kPzOSxvH9KKNkB7mikn37qVsN+IRnXVLrPAmxGt
E8VIOsCJws507+jzD4j+QHjGfCaLzEp6GVqzaHF4rmnnhNyP9tM2jYGG1efQN8Q7
b2KRyeP0sETWjY2yBxGKVVaBGGQ9GYVs+GpKk1vaEULeA6Vconkqw7ZcSQqBHLiq
kVxZv7Cga6ZL9fUvt1f2es4X3zo2lkw0Pgi58HxZbd9y9r17MEEwPIZXcGd9DUa+
+r/3XvPwMi23RyRItg5D38RAyj4pBykVhP5Z4m/73jtRgc9KTIVAS8y93ySprLeb
fZDEna3kw1Ac9PtEql48/aRJykQJl+Hk+Jn+dtuh20skLGd50DM9meBneWY1lcn1
qOvsYNDrPCBC2LDykHzanzKkQZ54yDVzAZ0ceGFzE8OLwToYyAiLVZi9U4YUqNys
OJ+8lRg7xmxgJDrMajF61XXSG4X9IKJpKFoxnP4mSRXrVF9/0LuABENZXZJTnOS2
sJC1uU9b5jlcKN/1kdZvb1PuEa7JaCw95NhQEVke18/dxZVClEvSxGw1n94lC2ZL
VEcPlq/dh069WeL37tSXrHUtXPNJGuToXI9VeMItu/RQA6lfUER/Kqk21NsOBHCA
NlPg8L06Q/8Z6Ujackj7x8QQ7UqQICuOWriX+3QaY1IrUAkU30/DgNxmGnEATG9O
k8LsYgODwOhdSZXiMiGNdKYRZxbupK5hb6KnYBKS7/9xbXaQtzqEalVrpmTpueU6
KqcRdNVey4WYZMxOz342oTwFTtmzJIptWPPEd7zI1QL/O/ys5DWnmOcLuZ8Ff2CJ
nkioCVUUDxuyY1QrJUzA7lSnf9RHJje5/lCXbFfgu7QvlaVFYxZzHTr5a1xE/sJi
6YBcq29LSZPxq2Zjvp1FbYvrL6aecgllMpTeMTBYU4oApxmSNYR07R5qTjtFecXX
l+OhcB6GJXllEec0ZPgceXV7tMzdzda6HRRhn0JNn0Fm1j1ZwIdzwByTJ3bJPInP
tPoAFfM0o31kAjiFQOqPtS7EajF/0JQXgNHXrMiIx/CchZjGdpl6P3jsEjwQ2INI
U5gg8mymWYrKpZH+P9u9h4G/9IMCqqPrU5kKLsTnJvjPeLdiYUU8uSbG3Q91M7hx
glaRwcN1KbcgP6a3Y/PCTOLN5xXYIVpLv2onsMrCUTOzSGMRH+jGRp1dqqCSHOh0
pxl5jOjyqgxXtwnYxuVawopLi8vDhzIF4G4tAgMHahfaB/xorD7RSqP7AsfoiEkr
JXP/9l1O/ncFeyswVOvug2O5gX5wQ/6eLpGRtbeRWDK4p7r23UvVR3yQasZAUpXe
cXzLtH+rrK0RpuSk31TxWI7VhmxgPUDmFhXyKauv+Xxmb+lTNdiXb6I87pxMvfGO
LM9GkUso0VBl8WYzQ1hCb10d9oU+N0W+p5doF3+NIRGY5K1pRhPsoQ4FT/XITgz8
WvkKoivEiBv1r+Xuzex3JCnBHvf/tMMGo6G3fKb8PVhr7YfuLuGRraYB5QpjUsHt
qGlomjPwY/i3c04df7cFs0W4xvLIuTRGrHiHL6czxls6LV3IC6dF9poQ4VuhxHbf
FAK9joY1ZrrR85e5/63JkWmdJn7DfsE6eTiIJcG2rqpixY/tnlUq1aXiwwCLPbTN
rzh9grG7gknaBul1bBsT08gaJQTFR9T9NqoCaIGYPvQYfX4Tsd2Dbiao3qTpj2KJ
jLlKy76jttrebeRSHH8H7mLX4jDMIKho443jIS1SHj653nTCJPa2dq9h2W0BVVvZ
hXSBw0286hGgniGYr9bjk5ywXbUrhUoNj8xn0v+Ci5Z1XdIYsVZHA1PNUoQBy+5g
XFrsTn0Rc8urqqRE2H5zxQ6PmV2CW7hNZkaLpW9X7WXRnBmJh8+e30v0AMbH2WI6
HA7TkFTuMxLLpcpYShOai3902ruga4kH4cJrrQkX8F6GxyBmVqSRI3/zDoozxqYY
wqEwb7jAdjjSYIhFn3gWqEv4GSY/RLrB6D2+0YIkuleW3LZnahNHrz7emOUVI5h6
wiAtGpkCLbCdtoaDQjaNzSnNnJ8PV957rQYxb+NIJWqGPrx1ZNcxICLJ2/3FcU8B
fBCoExKMvSq/ziNBS71zuhV5Ibs0j9ZTCZO4W9GteIwrF3gAXY+QhBieP9DQtmu6
cz5QousS/DY2ZlYwvw7oN/UewNd8/HIjQ/v0E1Ea6hJsGK79siZnObcUCIvHze47
Ip0KeD36qZDQA3DxwS91kPPm3tNnQG00ymsixCl/kcIXDR9y+s4csk/JLpoOQqap
drpeL9RduOkoY682p68rDA4hQGhBVbqYi1OSo+4iXiWWepDULhgx3xf17emqgIa+
9zCz0kcEiTcZklk3E8qevL/Ebim6FPUM3mJtw9aQSqNbUnN7FQJhh/26Enrfb9UO
704Y3Y/yXQLzOzR5aA9LgNYQYeUE1LWbhdy902XOFMkZrLDAjMSmZJgGVSv/gfKT
FA2iCbrDHdd6OZVHqqXJiiq5S/eGcSrfkGEAzpGQzEnd7udVW5CRO8FjuqwwIx8W
4PX/mHSqVHyJY7HOSSnpjDEYMG/uyXWxOJ4QCW3XvftOqfEiSkV5ieguydH/xtt+
ajpJHzPtTQ8Sula3xtrKcNuyLqVUc+496pxJar2VnwY4shdWw5i+qMhTqLkpvT1c
42gnxqGpxCV+UzIZo1dtTqXsw0Xw6KXbi9642S03utt/qUq/OPJvMJ//VsE+Uxi7
NxFyQWttpvLSns85Cl4W1PY30N+oggDtAtvapPNl/EEnRBMYAb/zHUQU8JEt9s50
NpsCS4dwLE7IwF5ymqhjUeJO7b36jkqr8M70isuUwuE=
>>>>>>> main
`protect end_protected