`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
FiK9KBulhkoyUl7dzWtZLepqOja/wRUqNoKfRczMihfNA0+vuPNW1Ro/ajw+Cx5B
SDe8eyBny6eFH4xtvKUngeXul5rqgheY3/ic0k/OtaNKGyZsayd5ov6Sq3T+mdx/
dqVg8KgeSP6dpN4MMFgLSHKCCAJ9LgRM3tJ2LdBh/hG79qxKyy3/9yuExMs3TIv+
8DVps9Q0SxwthbRDeATgOrnJ95E5eK3dvuNT8dFp5cQvyYPV1KaeJy4GUAn99gn/
8Mg7xrjHncr/MxpV5kn1Zvz9XKgAR34sNro1t16LQzWNULjRbgtr0WyPkRrBqfmz
MNLEn4pRUPAf7ynOdmPbig==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="je2UZFMZBKLAw0ycXhOix6Mzrit1BQgW38MjgJnVOLM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
dTasYuXuXXYsdKWrlSNxlzwKHoVs3kUzJuN610sYrZjpGFmu90ROjpuqHFLiloSM
BSkl5i7hVB7IbVIFxEnJA2vvumaph8tBhRFiP5L6D900GYHevUdiU41QrAIhK2vG
cxkZl11fE7X015vErVMm+6FLEXoxR42NXngd/Hq2RC4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="8MBqDLcIFGCAccq514Hz32xwDEuFHooG9Pd59L66LCc="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20704 )
`protect data_block
uBOPZMumPK45+cUL/4s//C/96uNlAg9CCCFD6cZUfT0NttpbGnCgBjgD0fBKI1UM
kyTtzRm6jZ1y83Mmz5ri98qNy+I8K4BRRnOW5vpbZ/Smepf+AWRTsFcGjpvFhE5R
/GMbQK29Y+AAYqzOrLs1aYEGshOCBNLOAFPz/YVL0JCzQME4UTUK6Ien5NiV5Num
fnKAo+9DZvwCr1PpllYULJHQzCSK+cyqXe8Ii5xGc+TmpX7Rn1TLPGqYBpgHDhpO
Eezjmp448gkBoLubVJz+JlASrYjtMdogK/HlgM/rCafO/UFt5joRCbFSIkPhR5qN
31JnF5nV/G0OKAZdT17jwuD3pmEUpV3gnwUx1AQQSj4ovb7dStiYChf0qL24qS5z
joFR0Za7yFBuTSwmppo34x8S2cMwJFAe6AUWEWJDdnbgYcCN4RPc4jqgXlU9eaVt
HxIdJBnK/aOem8uHYx4/gzc/Tk3rWmE1VCd26HIBHC7oXzq4CIgFwyysADO+dBCf
XysDHZj9t/a6uCUTu6UoN86JT7dlvRwhJVwk1VXqBaFqeFIj/l4PA0bz2LVx7xfQ
I0GXjeE0kAPsZ+odK2JSGd91UbAxCsLpR+CixlCJ0HeWPMsNRF45E3dRf70h6aiX
clP0arlX7YHN5/KdgRnHQloUOf2OGDEjHFpbEGXW375FmWeQoDMmBt9tZmiwP6lP
B5yPQaCX+0L0YMXeuVCzxRqjSVttOctwC4155D0pLuSXhrGw6HxPfE1+zf3Hz2hJ
HtMO+d1RIqG58LVqCuCdUrf2TipfqQlVz3/2uAg06pLpNF52W+a2+rgtvBt0yzoY
l0oE409kv/pAldMcm9svO7WrKu3rLXuISxFqnY6mia0/JOZpGF/WSYqcrbJSMJg5
8hXANnHtzdlPa7gjnSGkvRgT+lUrw7einxXaNs06AjJmT+SZczqnRlU37kO/xeYI
38eG9/aPctnThfYdAffAIeUbyvxo/nzy8HUnFfEMc/f0IaGXciHEyh8NGmqAYS51
TedwCQTSANwx5bbSA2xFetQELN2gwWn+WgIQC2JiUf0dPO/T82SSemsykwO+NDCR
tzCM60zlUKJ7r50nAaGpP8MxCPVVs59RTKWJdXLsAl4g1XapJropvkEcH+N+GQ4K
WGssKnmhF1VPiR7NVgeIeg7aP6bxrLdFuTglzPUH6FyIwOhjVto/UptmsBLCvm6w
5yoNtF19ZsFxDS35pfVzgRRILaP4c4iwCkrcTiMNlAe36Dxlx9ULI+uUBN+ecqir
ZRQpZ4wdisvUGejGvz/KXvXUqXqlmI/b9kyBrO1kz73XHdbSmdwB82DTgxVfvHu9
ElW065GxqU+KDhpnwTkAducIvSCzw4ZR/8lo0zwataTKI8tPXygm0o/6kRFRs2yc
uk2H/d+lXvnZfCAqGz6vRXk1g3bzDBmqZthV/Ah/2vnK6EnePYtvUwY0xcVCe8QF
sNV4/o0vvwGPCPi2yOwUEVzVvflxKUMemVKgp2SvEUtu5VvHuLid11f5RzyFWqGY
2FYfeob9j82bJix+591xGYGqbsTZITQtIEdC+loiMQoOdsL8/NPLlC6ALmmjdoE9
0ulfExxSgV5UBqq/gyO86cGqr0WxljlTPrIldEpt2NNgpAhMa5AebkHpNJhATQN2
vG338PSoSzT8xMZXCSDHFwtYBUpWvylRL+Jp+RA/SLVKkSg7QU6/5Cnuo0lj22xs
8sF5GeNZ9Bk8ou1i+zmfqTPsCY09SfsarAp5b1i95Ihn343I1GJeMwmiS2orDppd
Mv+8iLop7qzDyuxW1WnR0E8DxfBvCvzmP1zWBdmVgS1nWmj0GUkyP2wL519rnSSA
UIJIjmvTKzGxdBhWR9PudhrXrPAiKuPf9C5HDj7IhbX5Klv/2b/O0Xe4SpDsR2GZ
oiAYx4AeFMQL7NqYejRSn4no9hKRt28ian1wb2KzxKrk4QY/ZC4BkMCWrSunInN2
VmlXfHhxdrq2HAsXsLFw4CS26Os/qbbCxmPncsr3SmpVwQ1/REkOvGTvuXYV2ph/
tpgZWjFxlfrgzOgsltt4DVhqc3v7P1/Uyb0mz75spB1tLM86gv5YTvaNILOOL97X
239zaQ1GU19uFZ9y1LX81HtiE6iOB5XcssZzfNOxrqS+mP8n5b2g8MBMouKIl0D3
9n+ZylZeCB2DFerzkR86LTt8LPtmU/4QmCr9+YOfV970ghD4EDXSNfcWxRc06At1
acZN6kS9N+3dRP2fFQ6SsqSMm+UPoQNTR3fDDDckmBnFpRo9L4KY4X6caXSih8zR
z0lMqADg1rhqNJLJioVUlanSEYb0UWk7ygAvfisw0Qh8Yu1O5HNKhrp87DUUUBwQ
L5v2wmQ3muYiETCJL+VprhBv8YtkgRNBl77ylCb+3TGnC5M18SL0NJ/Y2+Z595Ep
RltpJlGCeFof+Q6ApyD8NKokABzJEym9gozMzaSP70ZznzcfdA0995rYGkW3ujME
BFz/6UwGwB9b0CbsKNSuhc4W+hN4jpIJQMlGpEBBsaj7F2Bh8ygXuyJXWS+3ecBX
e8x1zNAH5Wh0fgkqFAB1ewtbbXpKREb0rLjKiVOGVE7hGMvD7inp1473TbuymlCL
NL8LRYCTOwxVxyfmlDdFgXVPXOmW0iy4t2Retb1B+Eu0BUkgRc2wAwBPydJhzp80
am310IOTfZ6T++2B+r0SABtuBCaTXFKqRQiIE5T0vU2Hig/X2lc1LlpXQstG4yFD
AMF8C9RU5c61qNPfGbzX0uCE3XDnlJevGWr2IK6GvxG1qsPjjzcXKb3Mhx6syd0w
Hm/YeeN7IySQCGnAfsAmw5mlNku7v5r22FL4a68gFgfMEn9y2gpQRPiBxN7XotoJ
ssfikd3tGVTolSGk8LP1dB9/54XEv9tmktp1f9pFd7J+8PR+9sZxFeLdycHpoTLp
C+/569ytgLobm9vxXHkUHqcBrRyO5428D66d0t8pBsyDornWb1i2c+vcwkfcN4Me
pEbsMyHkg54oO3XTSPluv/DnVSRb92WRI7nLMcQUDst7f/xypiZNbx7Tcn//vhqN
/EmYhTvCCyodYUEXEr0HXYJVogKHjPT568YC7BWF1Sp5CIe+065PqC0p36rR0nsR
ZTwcZKioR4T/j9HLW740NUmFLAPIEGwuFzTbWdvrVoNY92PfjdXXC/PsvWK1a3XX
wS85+wc44VQx0tKKPInCi/35MnOthPuSeHKNg8g7MH2WgYWiXU2r/X6JEx+FCWOs
UXVDbcgp3egd6AIJuneSk6IR/cikDhB1deoges3hy7OkSoydTnGRPvlOlHrGjsha
MkCLHJYb56DAbxPwmiVGQDUl7qbUT2C12LOv53CrN0dDfTZexbVrMxnU9MAd09ad
naXxfPniLbkZr07sdUVGLAMA7ry+yYyy2yMVnmad9Dt3FJhcS+iSnZ4OOHi2e3RS
j/EtyxcijSoCNra/tXfOnrd218Jqh2U1j/S5m0rUf+rPoyiNy3GpzVMRPZVCjkK3
qs1P3zIxzq+cvKeX4IoBGZYGe7kTrSDwP2XfvF4z3BfLyLwXaeu9XU1OQzrMTtcj
I8DtyxHpiLNK70cqDfJFrm3nU+ateTMIbvSVJB39tmJ5tUBIqxatkwq4q2HHR7gb
1TiXbi+AdK5QlOp6oYtmEUWv8s2iH32v5e4QOPPnSDvDUr7o0EUy6CkB//iiY+pB
+KjyPPUt8xff/QLPFrM+cMfMCE4A16DRfMe/zoPjZZ1i6bBE5aL6y+z+sltg0p0L
UrWhRLS/LjwUc6GPPHvlGfTrJVGhDsvWW30qdG0Fx6a70ulwKW38nWMoNAAeAIDj
OTjbQ4EuymJiaxREZdYZmHh2b1TKRFPyb+c+8gv3J1H7uXxchA4ospPiSzB/08bQ
pWH9MUzMlx/1tTFjJ3UywO+f2L2IvTNhq2Vn571/TgfIPNmPusHo9tsxqAqi2771
PPvBoUDQJb6chDAG1+NDbqID7BfZnEuJi8rak5iyszGBlGTX4YBhul5Uaes48n/5
M1vP1ECgdmsL5nec8eyTtKRG4npxgEFn6rxdOQSROni0DznWyqnNbQVxb8UTne7/
ijlpzdSq1kNlNpcaHELm/XyI2oYgC8m+Gq86hVOoke7G8vrm3eSIMpW5TRogVQI/
9IJsajmqsHXT0YAThJJRpphKuC9SkX+vYJNotLq61ettkArFwq6UcVqX/B6VdJcG
VwHNt2HdjD+WfsjdfAdpAWS1KzJsctwaA8abaY9nOsUNbhIUwMqzHpYHt3YBJBQa
t+zZUavCR8+kAyOrCIUY4/4vCBomEl3AXXUNsuXQeH5hQGnQx+X8o6bA3NijdpR1
42bOpwyxCb/bM+tjMoghvkM3qGvTSbHfZ429GyV4xE+kO6m+uyzBPhOvjC+OF0yj
APCamuMbpXYfdb4ECWLe43Je0vvX6AsHtiISG63YSk3JwmEueBhC0803kBT+M+kv
6RWJhXxmLkYJWRLQeog0hRjj+SPfMw5vkxmZ0amrNmf5SFig1g5pIC5fDMZMTbeI
hxcVn+fKY4UOyEJ3MBXMFuuTXYq6bzmHvwKJX8+12n8Ra7ti9/TMMQrDjXj/bW0s
aBdv8QpCQhboDGNocyRGBBCdbrJMTUybo0ct3pxikO+K6ddZ1w6ipasHNnLVuE2L
Fo4ioWCCB6mjg1KZYaEGUBO9pzYsQNvYNEFlw/bPrDdXEzc5piWAWbk7QglEFjgR
LnIpYgN5cZT4Ww4xlPJJbpFs+zdiRUktsfjVhd20uY9ymONzDpstNn8UGf/xGEAq
pT767gmSUPTaBsKz9+TlArbRlt0XstHBgNJTczbniPFSo0eL2VRsSjXMJEbYKTAB
FZo8ouxfdqKhjC6BFvW85Z3t4nvujE4z1Trlo0VA8tWchHr0suokLCfbQzakDzL6
Vn49ZTO6MsK7XuZdrZ+9Gf0gz9nlTzhnrqSzIET8qvX+nPVMB16CK9COUoFPSHKg
GiS1QMz3TUoIU/Y3P2+d0pW2tvNHWT+TST3+eQFQWFqiHUVdhTxoUz072FMIO92Y
12rqR12HzMy4KhRzpJB8T/j1IFS7fIKHXbhHbkLAA7Gm/J45lYXjooWlATyn7BJJ
i1+YH52JY6ueOlw0KT/99I0jolN6hYxH4HLTNGw6LtwyOElYKDYcRhxK2GCCmp6q
ySqZXjfBdYTxG3OZ+++CtjbsxZD9MKOKFoxl0EJ4pRTPAsko6lvfjsu1hTU+v5II
8eyc5crMDTTYKQ6TBHpmA/PmqOW0SSRAqGmUyiK4I5y1EE17HrVp6JUIbHVXq30e
X2LSfFJ3HiYqDICtqzHSUDAiDPVVyywwekW4fKj5FFFoTb7zJPjaKT7D6BPu90l1
5ah0O92dVRI/zmQlg+YWgcQ91by/2ynfyA7iALNECMwuqbqSKv5Up2s6Mu4vOjBC
rYI99r47Aeq/dooxT6vwmN2M1i1PisvG8xrcK4nWYDK1v167gt80cYA1lwQcN0Ac
OMAhYFmkGF1k/KB7sDsK3e1wU2TOfay03ueVrJlvxiCxZDiyzNEiWIg+N6ZkoI8b
y+cTp+Gax3AE2Dd0dzdLM5crPEKeFO2vpEO8IRWQA3pZcO/FsXVtEWMlCQ+2bI/Y
18xdPN092J91O2GnWTKY1lAwikxt30xWV0VyXEUSuUAk6tcnopFacrsxB/mlxGsj
9s4l4A7Ea1HV7x9iwN/zHLBXTSsMpFocM6uuj9UEiDqJ/fGrAQDXpCft7APe4WG4
eWrVEHZMgkvenQCogbtR7Ht1v8SwZXVtR+5VhQXyhg+mg5ZL/LzL/yOjxGIlH6YN
FHOgkj0qKsVwz7ov5o0pjPRsSKYevj5FuwEivYxxIVyyCPe8AVoggCi4tLLQjASk
3L6POM6dCRZGvdtaebnmn/6EEgjiQUASxwcteBnNYJqVApnT5UWTutTq2/11sPgQ
1hMuy0dRJoqyXfl/NIVADsGGLwDPfwW/hUIchWXL2NO+stL9ZNMZZwMw8RR6N7Hu
Ykh40464X6EbNLNAmbs1J29F43cWxfkgH/i2+woqF/HLsTcG2uwArQJXqynb1PJm
3FByB03Vzdkzgxrq83SRT9+zenzdo7HUNcGMVMBcU5FbaF2gYS+WnuVUdRfkEzC4
Mbfolsg2BjVkFrBJsbVJm90oRvlgip2LHilCD78x7SPE2bkr/K+QnbB1dZQWDBzd
lv1osa5rvisjnOLNqxxGK2UV0Y9h8p/haBeMxP6iAm0VZpUanQVQw/Bt76Kq8Bfy
Ou8yBPWtKHQiA+dGXItnE1+bNBN1opYRfSZ5J9QnU3w3ccRXLweTwOKwEI7YZwHP
owMXtArSQhrYWz1MMUrl/NPNTNJeo8pdKLysr6X62ThSRkm5SEM1NGXCAZSQrLMB
H6yVg77I439qzEVtwEoXJrM5JThPWmGz5c85gWFV/6prdHNS8Cx9DGZ2zI/CuQll
tkfgvjOCtJsa2/12be3jGUEZkdt90ceiGVqC2Iu/8UySf1DdOEI9cX1pIGkPo75O
VSDot9gsa1Q+05f8X+oJdQ5uPc2mRpGIOqNR+WREKFvS2McuC+n0eJCVplIlu+Xa
NLnzEujTv2ucd+5VxEITwmqllTIXiNcq7Y7a1aye9mo1A5ry0wzDQSDUMCnPeO0+
VCRkrZYluglMy7SHb0UPIOcXhe/y8DjNkM9NyWB1HCEVNGKDw1lf1mUbRBW6mg90
7Dg2LiJgxZZD4v+cMwZ1dSZQdhv060CNTtFvtzSVjyNEqSec75O0TNl4L2i1M+WZ
8MeeYY8VwginGI6snUBLoQ2P/ZJRsHmgP7ZkYRjy0uwHaLfCI1pH/Q2kfU5U3Iqc
R5KmAs6RlrKJJIz2Lao5xJGlYqa2JaFDd4RUfRZq/XeVGtFSXgsTABLgvSazJxVW
dwUnh4tW5sCFz0vA8RJSIvfkfqkeQ62UBx5T3P+x762DD4uecR1jd5X6oN0Fn7Y4
nSu0ls1TT13PhXedh3FOMQHdY2NKh/wh7Jk2omqgbWHYAVrgDNO6PPaYBSFHuuv+
NLfTwmHtUyZYbCah8QHWcLqfj7OIVBS03ov1F+cO4XhvEynahhLmWMnVQYrvjykq
Ch2CThtN4xlwo4KL3dmZjjXuzdnioAoPJu/qrjnzt+obXytefw7mJR+BZaxxikcK
J40WyrERxqhzodOOL8ft9FeAd/BTpZs/f8itdkcGC+Of8pAwNq6uW9+17HhyASnm
nJWjHoVBaO1bSPMYnZE7YWHT0ZOdVOcbzd8yqlJUwxjKKitMJlSyVDkKU6H2RPlh
qZSQ/qWtS6oav1scyE2+yWLyOQ8AWk6/8rD422IqSKPuRYy8Bwo5/HccSmGI2jsl
8WT6tdKhaJ7Khk5MFojtT3FMdJWh/KNi4Onwv0hle+A07qRpH+Nzy+KUIbYzt3Eu
GqwfmTmp5Nc1advphloKygYh02yRC8q5g8/2WF0vTmVzLLAK4TAPru9S3fU4xSxQ
x7ubY9C9za795MtjphifC0CHf80ZFnuicGEmEJA+G3WCApoVwLe05F60VsCiKHlJ
XzUW93WrNhp9clywGDCfTvpfuYYGGT3Kpj7FEZsy1O1F4td8YH3FeA4RsW70+H/2
9ZSIhpzawPdgB48RscBgdgpfuiCeGBqBDT9LIuYMiXp89VJgzA3K5XmZPvvUse0c
hU8xXMsb8Lj7VlIM+KcThc2A97QpTeV+Ymw7ckv3iHUSkKIwWlQIMbEFtHt42h/J
eV/z5BmAKVuqG/Ey8N39lk0e/NS/1Tt8qcOQz+XDykJP9Uky8Kj+HnMZhGV9OgDG
TodQ2vU/v8Ktj8UXqYd0TbtdWVk1ndjxXOQK66IsU0q+TUjfneLNxPYVI3zZvFN2
ElDhdAX5WGMOfdz1uzlfTdGTHFci8eg0+ehnc4AOaiCGdC65S7rZDDTk+m05Jx/I
yKrdnMUFKdrY9LgQGIYyrikmQLwZ+xQPEAXciKMaNHNA/c9p3fi//WyK0Zkm6oJG
dFKJKX9E9IZoDyvm9rPQd/maClSHR9GoXMauwPsOnZ0g2zI8xJ+RAG85paY1GKiH
IAqS2B/lHtn88NmMhNR3ZjIvOoWVnwHnpRyVQV2niTpu56vdsxzKunYWCSG43v4/
Ln61MnQmBWQbzbwhN2yHSr85YhqxvIbbzlURZiQ10i9mNnMcXIj9YRj9ewpi9dNc
zEQmsAfNcT3KPIEp/989BSZ16iJ5HbkwskRNp+E2N+cKiZ9pX9+QMLq4RNkKoyJi
jIPZU9I2cgFXxVDFetEnNwXcvrBzSCC2JaLLAmbMW+hFy3zgBn5u97jKT2208KWe
nOGQZlVJDr5egw2+GgezP7VvKNQNfXMCvjLzKBBN68mH+V4isXdLFbvwdGfVEWRC
SZ8orp4oqapZ8/Vh7a7XOBVvICd8YIwE51UvzQdofEXk01FcjYl/mYnIsUMkUyRc
Yf4tr4k3BwjLL2bEJyWvj91s4nogRxP8ccPy5VC5k24CszhH8CYWo9XbKD8rVH1I
PFI1XX66QWk2X/y8pmmiJYbNz4i7Y7ZxlLfa+DfRaKv9h9hLr1mwqXC+J6ecPybb
dwx3hPrJanzasfLZExUiOCUMIiuo57lQBEa/WldJm02da58YzNtey14cLrHy13Is
nipC5uGB7oIWTSz/s7BBitcUiQQTA2mlELr/1piVFiBGfGz8djfj1rDoaXWdOfUa
hVzwJIP8+wn1/D/07pkbNPr3U4qj/KG9elKsk8HUOSHsYyZRa4VULUVSteU6e0cu
d61wxgbK4GHMerjekNjo9YdrphZHosZYI5TudHH6lOEYl0a7Bgdv1y3naLEhYNqU
vwrmeVWxJP8rlQg7sdg9TJ/PhRQ+CbJv6NLsLLaaKPtM898lKd4uioWz4LF1LYmQ
LJVntTWIQkDgN0/adX6lfNRSl7wBz4gaxcWbpj20VzN5k9zHs3fRqaZapuY94Og9
3rb/Dsg+60+3LTJQQ+Bd3sD9jrdShhv2KiNeSaM4sXF9wkHfd1tkRoa1qnfXVGNz
1TEKGUJk8pqAE5jm49MKcGxQP4nP/YHrUwzmi1WCDPTnecEeMDr3CXqlf768mFSs
H757m5qXmGkKqNruzp38kZ5pOvfuIbAuKcDZEKjT2S9qS07dUFSfpXtpd/QYvEI9
9I+/7QGl1gcxKoIUdRBL39hctWALK04pyDFq8G3BxQQAA5UTdchya8zmq5EhYX0k
tCRjeHNr65fo896coBMaZCTfGe9PhfL97tHYO2MtKL8QzQ9Y9RFAk+eFrVjxLx5Q
M6LWCsrPD1heaUzlF0lVgmnfTvembUOH9sqqmrvcg2b/RRpOIafct1DAqxb0o1dJ
zplZK/Hs8gVSUj9fUvCE/v5HOwjC6lmS+b2T0A+3DcbpphwodsTpAAVwSUdloDJN
zebi6h+pXY+VGAWAtf13j2W1tHmPGFjONsC3+/qvD3pV9puOOErLNDJM17wnSZcm
5CTd5xK0Wie06nRrL+BjElqAZElBlxG9cuak1eIU1/NtuUoeO7AK6LLVHsQJv0my
E+RlgNTmUjjNsS+1DL+ecSUBg7qp0XTcS/VqCtUNxm8RRYVmRPMVGempLW+qFyLr
qZ11b/iZ0M+L65sf1sXXkQRuA0+U24eAjEDg6zfCiv8fOdxuKqb6HseBYLDdB99Y
dccJQArDY62tFCi7ep2Shrx50XxOptQaVWgImZFS4tMutvWVTs28BVoMqJUARCis
M+5Fip9dxyqnpupgTq2MLoz+hHTnqN95ZpH1v6/5UbaeJM6TygyD5ZqnpRvr8BuW
q/cgMh6tNIPmerOGhboUGgq72Fo3ND3Sgc4aK0pkbzUtjmPygTekL0ASTlPthVwE
sXzQzKDRLuPGykk8r0E+/ZQMlFmEGfq7AuwQB32AfAiNu+EIdNiNM/yByhWY2gFK
R7HRCe+3O5e0yr2JMrt9fHeSYkZA4WAIJkgSgZhQ/sYQM0Pj4262yLnl+XUNGA4a
qF+EvWpXjh39Sy2NRn3DrK+VrzM37BxLd1TtwChT+4PTnyU+vlo7k3Goe1as0+z7
8IAGOgZjBm6OquIuHKGwcOkwueSTMt/is46CGO5o59uM8wcuD3m9hqEflAQxoUxe
9A7IJpZBzjVbKgo4zSvYjc9SiCnq3EDh4i7JvydhpNRCHIkCJqVryzmfwYD993uI
7Zqb0HOHcYFCVGFj883cpizY5zvQhEZsKvE0CAEr5sOdDjzHX4f6cF1gfWMwxS2t
cxMwD500krS8aCk6fGr9/dKxaV6HF3VX1KStnoKTCPXzlmI5pgUj+eImhY64MOCQ
YmcwWlWwghTu0pkKm1JqWMScU6wNF8oqAeRqM2kqz3puTtAKLypGUBp9iLBqcB6C
FKktRUsbbsZSOS5RvZRYhp8LlkFzK/vjh3JOZ1JuE3kmR3skmE3qwah51o93lQIl
hCl+ugmTFPRWIXrU3bSi3q0qRu67QJLEt1tmAPxIx5CIcjACkM2SHgEjHNf2EBa5
d2S9N+qWBUExFJDYS7DEglb0Ck3t9ht0JZnu4qQ9/y+l9TIM6pFhW4MQ/51ZoGPv
0Y9gogUoe6yefAJ2oD520tXdA7iB5Dv0o5uET9vpPGtEYrKoWY5cjlH26SDVfvMM
ueZb5+09L8p2aPZZtCAoB3zTLlqZfz7+U+3xaL8SutlpbsU8FGroOHdL3asnZ1C0
SiFA6Wq3nn2DhckK1VW3s+t4tRelZfEzrYPt0AMxqEQm2mA7iVQB6y0xPRe64nUL
hnaYOTFuC2iUC1Fn0y86Ls68SAlew33UE918Ea5OF44VqcPgEvu4r5nNo3bNir0H
Pr8rKq/w0p7sDxyOykjV1qfKqGZfpGLqqhfvBVzlQKsPrGWHoVRV/5XawyzDRdzh
tH/how+OqtQJ7QMFX3oNEXctWEruYgtmkfT5tev2JAc3l1PA5Q7NCJTJwfVTDR/O
njnlKx/ZpMOEEZ65ogxsT+CRCl31QfA3eODWwutFhM7gk9HjJn9aHB0ExdN4G94X
8zN4PpAgf8+CrIeIEPoIgBR6VznPrx9L6eYibt1udrTem9qxLlGtszCna1okUtqt
b1NKVYr8+D+xbtC3bRMEC09ur+MKaX/AWvl6Lm/d2qRSNgHIAQ64PNKxZtmVq4vE
tGdMV/Tv7BF06NOOOrVgC5OKlw/Z0/ASTfWzHmkdmFBi0ACBtZzcHfiCE0QF0dB1
JOP0SEkWgHQTw50q0f0WIR4gg3u+zbLLlWUyt9AFgHahLXrw906282FGXK/cNsN/
m9ooDkEoEWaKBM/h3xv79jpslwI3xV3aW0dMsaxnPDamuo+Y6dGjr4OJHeFM+gf4
wxiUiMrYG2A2cvc9afcVpI/UhGfkG5BT2wnKIMm3K68ADsavRIKM7jNtgLEX9Eez
U6THrZ6Ot5pBeUT/YKA08KLtyFiBh97yuudqNV4lLhDqh8FtcqqdhpRuLLAGX5o0
fOdGLBzkV12c0c4I3wDAzat4psj50cocBZ58ggpNlp8c40iV0VcfEPNHi8WJgzf0
lkBl0iOg8fHmEv+hZmGUfIqrHrVR4edd5VOsFEssnMPiQ3vTrI9n9TlrQgGfHLLa
6MhxJrjs4E+wA/6aPIw4QQgEyZxK2RbawHD6J3RTU0ViXge4NRz0PiuqQZFM9Amf
BTif0lAKCwmiBVzKqqXNgu+F97BK/WRzYOtPhkqmyORvtDKugSPWDmY/h537FCLT
NxrcFd1LqChIiOhiH5gBIe8A64dB//QFzYhmCe/Sh943YzUkf7fhykKaWeZuKwZa
/LJilLUMjVtRTO2ESrrBG1sI4ZSBURhASAR8BLXF1zP+J/AlNigf/DATwV5Qmn+o
7bRgV3HYbi52w81fRb/0XAXfZO0XlOwz4wZMY1XRbVHfeqfPaWtkfF28QFDKqezm
oi9662iO6ovMbwZA0gpNMVyobCudCvt0DQM+mcGgk1NB3qYhdJ4c2Zh5qAp3iB+9
yOr35Zzgjc/PH0g8BZx1GnhBJ7zRF4i+D9+LX9Pk+y7we7NrVHXWqcUhlFgkutQp
e3yR0EeE2rigoXjR9yIxyKOrv2VaBZzkPZ0jyuj3WKF/GMJvF4fOydwh2LXsQ90r
M42+ytc7rU0DNDGhqLVSLRU+yvRNc5kzVM0vU0p8k1c86MgXSgu4TRCaGaBVN4aT
vbvZjhS6cHHQF3GtXVcHwRsW5YBoW3z3XD5ASkNwD0+nqF9A8mOjMlxivk08k9Zi
z0OrBqedI6drybejJvmsl11VdWvFhD7zsD1rjPwi3q2GZusrA59w1qMCsSwb/NjT
uGToOc9ONS2TFnIDCXGiAyZUcifSvBMkFQ3Wi06xzbwEfrIr48A7MKAm5YJ10+yl
Ew3X7yQ80zIDEAHQdTv+Qs5ChX6/7DG4C5Cv+IHuqdeE6g02Wf/CXeHT9ptqucnJ
Poh6xpjWlhmyckAqBCZ+n/v9PBCvEwZMeqc2wu/xaZq5c6KFKBywvlfSm3cLRF3e
gXNOUbMO3SVk6ooJah7yL00tkPyH4tJuEZ04dOV/tfeGnEJtGkSimOl3803I2xt/
naUA06K0L9noIkQH8Gq9NYOEHD+rVjsTMYWnW3sbRHsYSybHQl+/D968zTVHO4KP
qBlHNnZsVC4/GI1bHDnw9l6NBXcgEE2HFVepAiskYtH4rm+nypuOk/VI28vm/O3j
ZO+vVKHi2cBV+9iM3rwWqETlOvqRU+8BPNJjiFisTXLHvyX5xSqX+JggcsC26Oj2
g83NqR/8qHzcEsnX6cgSnbfceiW/vu7fxPYnCrJG8x1DLUaYfU4m0jv2lbY9drnn
LWU4G+AP+qrryHali268rdMyWg5IUbtpEEGZPEemhxe8vEw6jF+9eqvrJZjNjNY3
erQ4hiNMq8CLb9Hff/v72a/VBqdlqZOnQt2dtaJMYrhjmaYDnw4knExsJOaXWOOV
MO7289xbzd8r916mzOGh/javRHK63YTPWYjQov0rhYfXIbjspcSwW0+GJfEa7znk
pk/yJlYlYe2KZYf2zOlH+AaX7QleCCv5R0D1nOUaKQZus1X3RFp9QXOUDJ2AC0X7
bxfzOxORS/4iS7E8XrIIJsy1ZOZ/HXbYjV0aTRZKbb/jLFskj14NKUKJWch1wvQe
xXPYw6CAuNzlKqPV+QkgnLNGCiGA2UuKC/YF2TXUJDEXOg7NpmPBjSyAooWPE+cd
jMBcqyaB07M7Q+kxP5U3XGXUN3SypChzRovEY8oq6GUOW5RJccEqZorUpgJqQ4A+
elVlp9RoMwMXPChZ6bVJDVF0KY1cwhz78yBa4RoFwXyzql9dw9G3u8nEUPUjnP9z
ANXGi/bv48ht7WV2fVleDwzeUqV5s41E9f60YZiT1lF8MUqUXcYhR7luzVWiZi+Q
GVZNX0+93GDkN35bCcX6+ROXaJm+gx80ryEVm2l9gpQwqNUIjLwv7ESBERXCQM6C
r/CFov9/CpjC8/pFjN5pXA+Jb/4zlv3LuKWt+VqHQAYDlmGGF11CBTVjYqus2LDI
lo6f+0bXHtgL67O0Lz3YohC2xxdX1beXm/XCuGf9uWpm4vGmWlHg3cZjf6rlGPsi
ZYLDLHuCJLZWQHFGj+kWUPQ3/VUtOyTOBasYc9y9TwDjZj56kwJhzETzJxT5BIxx
n9hKlyALAjU0N5nc/PBasSxJm3eABdzisk+3FvfQyIb7g26b00PtqBGdx3ScVAT0
1W842EPVYoyltBGUQESLgbrOGLGmx4GM4QbU1vXdDFFMwHd7PaMCr59A61KvTXcO
7nPPyoQeAfVmXiHUgO7/5GNOjrjBhjSF9gMER4dP25GXEcwwTGC4dUa1q23V3XM1
8o11Uvl5+tiU19TvdcnA/Po2qAvjULa1sDofoD7b7mgwWW8bDX2+vrcCSy8ki9mO
aQ9e4PAyXmaLUGF4U1MkEBm6fVK9IgoH86jmiNlsBhZPgEMiL2T+nKDLqr2e2DCD
9rCv5qX6++u+1+qK4N+biE0UJjhoAWGMi6YqYh7TX+xo+CzwMUg6tvp5cGymrmrs
n86FhFalVOl7FHggCKzk7xcQLHU5slM4Gz81Jwtr0UZRMY6uxynEwaca7+ydNWne
aityXyELLlPnzkWR/RcLt0k6YcVei1+NW0nP0DB6G7CiE85KSxMvkaVP9vfZtxSy
Xdn5/ZhbSlUuJ65HWtacXgWcjrXzY9qZajWczjqPRq5FkpapPMTwlUku4vAEzu4T
xYrD1+tZqgF5yvztiVFvlgJdnOhNkFi8DwPAUbsKIY1pFiL4X4ePR1P+Z2/dWFsE
VuQy/V5my9u8otWkEW485EbqHW4nuisPH1rN1Rl6D7EcZ9gxwNIb2zaeTC4nNqdr
BBGKOS3LZd5wKuS1nbZvnDi3qnQffdJg0ejAIOWTI2sn9fVocHhQFxqCi10lcN8M
WNgOmb1WUBGc2noZbhrv1RRljaylCfWMZbae1y7+gv44KT+p+wc73TXnbjbeQBti
fXmdlOAVdYK0dAozDACsFmegHw4hj8FaSlhrxNToT5HTNQWqCFWjxwTVrdPffwlq
4cw7W1T7lC0B78bdLKO+rqOgD+33OWbZ+oadSZF7PCGroxNG3xQjrEDbcsr/ROqm
Gc30vVnKxTjUSly1tZGyICwjm74oyVfAKfsJ0p89/MrQklJ+iiwmLERQcm/cqRhe
PU95lxM0T88rchSm9uat8XnaR8+xQUlMb80glEFRvLvK09OK7Dn88VkF/cEkS6Mv
JgyUe5af1t1rDJinDa/TR2FmTa9zrDyoEIxk1EL0dkc7wzRkjaWbz8GSqYv/4B6k
TtT1yxe65xjkvNzBFwaESN5dOOEVkuqs/ZupkxEFoE6nVRrOM9ZVvNicIGFIIt8O
brWNAQEfquruzIyBjYc0Aq5HPNB5KmtQQ2lQkJ4k8QJJbtjGQLc3ebeEdSAIQprZ
xSS5fiVHB6e5JuV95uRTObs+b3Xrb7FynBBIxwST/KcwTSQIuOQ6oxWQa0PBsSC7
dHcAm6ND176yP1s4nlprcHQzgawZt47EEew9C52RN004XKEpcB/GJLuScZmGfM1O
h/4ebGOCI565QxkyaQgaBclMxCYo0EiFmeUS4PWes75XMc/He0DHyip9+7rlNKNv
8kfhCcGUkoxu+sDEGsxtY882WPbvzRbm2V+590mHqys/hssHUAzCggv/2owS1T2W
v0ICBWari0WKWvtvdUhTMKctrLN1nDhciK3A4pNHpS0t3AV3fURlnSjBkoT1OfLi
KKdrgh/Tn8u50kRwW8vz0xPFw96CLRsI0pxA8GFeNkzzkAmDyjWNsj0Idh7hwgDs
jywLPhbsMpd8iTPYESKEksGwz3Dt0gHclT2R+Aybi1fd7kB2dNiGVjuLK7CIfs9P
oJl4FALu5SzLlnLS0WZAcSQotlndsO9W/j0m6hoKimUFp7eV4E22cPPWabpE5K/M
YZp8+K0l0Dc6YacFYlWnXCfxUq2bQAKux6yCLtaFspGymJU8bpoywZqeEgAAHkIz
pDZ0QHlrv2EgO5s1TefKWE1bo/8QpQuk5rcjbjbB4Dnw0+Q1ATEgD25YGmGudagE
2H2TuUdl5n8zavSPSv+HOh6twRXJQ6nl18YadtI0nW7wvWLYMYQDB5bE+0BX4tR1
LrxAfWA9z6BIp2NhtQLZ8fJYpf6qsknIS6iFeXdDVPMGCWrhK0dEU6jyarY5os6z
1pdb0lY8xs6w1oEuM+nt3jOGvdDkGOvmXzEVIGywWvX+xu8h4e+kdEpmUidx2drj
jDas029/0Dukd+3eY5sOjzNSKbrl5ckYYMUfJlVUz1Qp5LvcXZL+e2Gfr9Us0ypq
Ar9FoBNaGqCxP/axgZgk3yZIKEf4Ide5dnEpgBgTj07eBT0/I5Fzqwr+9C5wcxZV
Z85tcevENBdrR29kedfHL+TFR4lXmEYU3mao6DTBWtk9asn/gFc+0qVURlwOf6RA
griXWFWF/XV/fR69PP9tGP9Zme2XejZ9apwPsert7lBKy2wfcuBzNCsFNAD7lxZ5
D4hi+VWuSGrmuuA0XvXeB8mynCWJYD6MmcT4KjCUaYA0zLN474EZOQDKAkeSskOu
xcRoTWRyWA7ZVxgKrc0eJFk8ym+QZ7Ohz8Nf6etwyZiMW0kWN3zpx4oFwWM6Zn3L
QuVsEfMTJG9zYFOUPhsuCx0GpLmDQaeQi/9XX3h2TNXCWOPH9+AV9eRTegYnvRZ/
N8nG/7pcuJWfeuOPDKeAoKMBK1tuhKACEBKZ0W5Bnho1gaWOLQp2DKdOg11vHHQ/
15db4pJDdEh04rvK6csoZmUe0AcfT9NjJB2TIAGGhv2wKxdgjRv/kfEqtRs3NLvE
BcdENzjKxWFycn+o8d+a9F0usRKUQ9plpVO9Y5K9Nta5Ye0Ir2brXqisLElXbIkE
nvxBQ0jyUNzYi03bF3ZNtXNf7y66ZkSmQ2XYkWw2omh29gMK4fsjSpmcHtMvdeMf
DBoYrxB/FnYJc3kwpEsDHmW0NNKMXI3yo319albet4vBe7AcI6P/dSiEequN39MH
qCHjzn1UwG0V79KHMIcFFIjNKuy+Lb2xZGRMnF/5xrwqLYIZhPC8ytRCqrVLnK4x
VUMJtFUGmimgyMF4EONuTp0S2CZDHnmfvUyPYjsU3FUQlFNaxgb+orTa4aHssD9R
Tx8uOxL16+xEhrBJuwu+ZUxU4/cSZ0mpRjPnFOKKPBKKcQyh4pIvgsHMTl8fiLNa
tbK3/REQVyanyYpsuyHQF/w5SwA551flIccFGpTlbdVVrsQ38M5t0YEggyq0Vlf+
37Tj0cbvvyfu7bUKt70mmwmPEK2rdldFkrGj1iGHcjfnhPtIDRGEq7qurCqHbBXk
CgiZTVswZ+LbbjjPyrlmsjHueUvt0ithBVv2ojkzoox1FC5vl96pN5E0TjELpWGx
FdTSSaQoAyqjwcJ5Zya96Cj2u/nDstG9402GgquXY0AkDoqo7SBSQ8W6ARgCQEWG
r/FkDcC9+MG2k/rmWnF0CSUP0XYJEbvpgKDCJIqIrDq7lexg9ryqWaz7atAqsoEA
Dh4gYNydbdMJwxK6f5Gt3D6NLLAFzhDTwD/n0Iw/0wVhVX1laH19TnFNHeZu5Rma
S0G8xaEsZZ/VRP2uvZzCSfyHatDPsr623Nm8D44a3Sd4iQpjqUPCg2jiv4BT514M
w0DT9nZuK65Cy1H2ERVw6Xod0iNsttR/KOsViOj57956QlFHA3ATEx9rSl1aW5jV
V7z+5l0KjtyoEObK4rDHSIRBWSa9yxnX6ywuMXyuHOkX3XZSCAoAhiACRuSmw/W6
HgVNoqDYmNk5HRT8eqYW4ZuTL0mdQuVPF5DycEZZfbrQCc6ejepYQBosY9rU12KX
0bBtn7tAMWGIRDzeaYQJCsg15bfa/NfLn1b1++GrVCULtvUTZuEcSsXSdyHAUV9+
BEFwMXjc5sVod//pkwN0MgD6k6roSo6akklRBEYhTPTagKsKaQZMYo3XdU7x8q10
HeIEr0epq5dYVzlO4Jsea49hZaIXRFtFJkY8sfeD/DRkqmNzxzDaZLOdzB0N74GH
t+/EqyIAsgTAvugPICk9j0qikAPk1AsEf8HRth/Iqca9noeC5gN3cuFthSS7vIOH
bci525VASIxDmNsxUtman6RXNne91SBu4w83HTXD0DrmIoybzuxu8BMvI4Olex5h
YrT6U7HvAp2EyPzVt2P9R/EiX9sSrKbW0zC1Jg5kowlZW1gPD+ctFZ+SvPB1EG9z
MD2m1fgOe/KAcnGrthkHN9Y4Ygv6Sz9fd5s8W5r2OSif4Kr4f03NFdzBHiyC1R53
SrGBlqOcnBAuoGa7MK0gpnlU3mWJLEXwC4BNSdoqJGJhhbZhu4rD8rcVSEYtOTIz
V8c3IZrVgEWnXLK/dcI5uATmxC6EbFcG2BG3+WI+o7kl3sWV+spc4M2xJS8/1qGV
y75avHSzSVA+NbsfPjYlHHecRYBc7i4esWcOEQa7hDvAAma1uf3YuhKk17a70Omp
KECdfMcB/VZdZEYMZ2YbmJQs7Y2VWZdtme6uWA6HiA54pVB8b49mnhtWddSNoeek
BiJUef8lOG7Jf3Cuv4oX5SxlcgLSXK7lSkp3hlogR7hv+WnvfFCpzHBSvBbcRxFT
p2GVIctSOq2jW6n5SJGwYzy5Qequ/wHStr0mSHdMjsVnyy9mh9sgdV9lIEX8kk/Z
aYTiLjMJl4ztyYNay0Vo24UaaxGtPqCI/tnd0pRIm80HoDzBk5PbFeOIsUMUs1rN
Ts4pN5pw1SA6o8/T5RGnyZxODgnTR7lK20jNusHSTapHRPHm0LBJQH4rDDab2Vfz
LqTYFJkUIkMUv5kuhCVn++iC1lmAcJxc7gGEyx888+hyBVZ/iNhWhDbQQx/01OS/
JO2rJR3DAR95+ORt/1mUtqStIbgrcL03W8sYHKbb52WhCuz/f4XiCrPKzuQ0g0qI
m0bXoJnQSL35PFEfDROxL6k7oVZ0NngUf2jBwYO1/UsOa3UDE2Qyk5I9hFuFiwMe
sTuReEby0+89sCGU6PuqbpjW/QLE6/z/KJJgzGazgBcOX9AYntma+Ms4zPuslQO2
OfwQ6i3nlUXQkbFrpKcMv1IZmHZUoyssb17gtFC8TsooR/Tdh/sa17hITXZiBpog
zkZY72+GDng7CJmUFssAaQddQdLgYR6DDRMTNIDgziyY7JsItAGKhmwD9PuCaD49
C4QVlrh0Twqz/++sgZw/e3Wuxrr+1A6WIXq+a7gR5Cdo85yECFv6GSzY1yWw1Pir
oU/bvmNutmi+DBG6+92XSAy6w0jnq8FJbDURbUu/K+F1TcVGzXZkv72yWkhQWH7a
x27VeUwXED1rsNFpC9TjAnJD6tuaSvZSwWN8kPaaiEr3ZIR/MDwW7I00XWj6dGCA
yrzWcrE5O8SkjjVmkvvLUDre8+Az0//krlqloylYXpYTcM3TfCFU09PchEUZ7zxE
X+mtsWIvj0THaLyPFxk6nF4wE2psnOv+YTV6prbPcok6wOuhrek5fIPAGrTZAt6X
7UOcjXy7QJofST3BgAKiIzA0JPpkz5ksGBuxkRwilkg8BqiQBp4DR3JxJaMRPRFN
MoLyqcvR7KBBMf2sjlJegoB6chbzyacKBAUHncSMFGD8dETYtzp3AsTsdurcu7Us
ebpAsf2CJKUpadq0sNFCoD1WlnWGEbUSmx5aafRpoIbqnts67X72+z6AtLY6DtVn
gbOWgtbs5wYTCPznbHHD1V0itnFvcOk6G2YW4KW4YhVSeRrqVzkpucOKMBbhayE4
LWXNsXtZgHxjjuPedgU7RXLaCL2jbkrAe2yqUwDDet4CXib/pAcfg/tIlpAmdX91
Ij7365gFJxooCqvyW6jViREtvMzuq6Z5zzdIFAE5bFog89fIhopZCrvWK2qUGnC3
nex5JbhRuQqOFN6n70T6hEV6SsyaOHeKAjk6vtGYIlx+8Yv5LV0yyBcWQnhk3G38
rDW2Nqi6jBiQD0d4APKvgU6ARvJ49sjPUQKCjKQyawlAC0xDW7TcqvclWFrAfB5/
XnCJPJCyvp3dxfyBKCBg49kp0ty6J8D8wiVPR2x7AaUCol2lqaqmN5vGpstqJiYn
U5XL0f1RH7XM9KEH6+4zBEfSbS7lOIPe8hOefs98/iInKnUaHUSNGo3eJoG54erv
33Yl99spnTgEuPxxAAjK2KK3HE1sTKv4ANnimdV9mu1vJI1wnR7lpGheENJGCfJl
R9mHJERY9wrFB75xtI6BCKNiDFxhNJR/ZhoMUOATdKvXeRtlq6w6vuFbRgtHYy5t
NMxIVU850sjoVafweAKc/2u4Es6Q9NMstlMDmNJQsf1V4n4amlcXAbBjAaHyQqpY
XizEBu+AF+dPIdGpYryobk+ijakzA4h9Z3gKjrm60Ty7HGrYWmwEU9sI5MBEAXcj
dWZSaD9/QvZMbCcPw/jyNCbjYUZqtboNMhoHXTsF+p3e+j6E+76nNxFia6D8I42j
GiHqt6HY5hTJYbSrdV5wBKr+EQEOUFI5/jtG1pY65M6jRm7VE4Qhb0I3PQLwXOnA
CaBZCi1mNvyVbH7oOeEKYsFRlmao2ZQruwijQjK7Cfhm1wg38+JYERAjCqgoxarB
WlfTMIOZ3uh/En/T601GVwsAKjDeGxz9j3GXUhTFEqRvULnagPKzX5U2rzrqk126
27zCGYhdwck7+/gRoBG76Z+PEiskXuapjQZkJxrJNy+awDxB/+y6X7l0Z08QxPYE
I9KK1rWsZhSnXe5ifPTRI7LJ0S0b8QVvB7Yfru+W/3ok8xr9Lme1RNFy7zVQIXEu
5VALAMR1IKroGm5tHOgqz6jzJ2qTd9A6JamlEqxJTGUWrS05+2NtR4+NxBksxC95
yaWaQRH2yprX0azrU0chKrCAK6DZD6bhBVsU3sYyiswyg4kAdfMstukM5LHnrghl
XwFnLVoZUdmjk7pk9ipcVTd/HYR7RVTFGRqAi71z+qcyK1veDCmXvRG8JY4cK1KP
TSXtC4qNFOTa+LnKVFX1gKnwt+OyARsYvWjYUE3RARTBXUDTnAutLP+LV1ImfkWb
oyOIxklyz0ulV6j+EJgYJjwCETiAYpUUQOnz9H3LYYBJpH7A+XUqGL16nyjnqXvD
JWcD1GQrkcNSeUtsYXkigP7C6E55DfcFlsY9vhVrDN2r9GnaXEiZodBcWjGRWaJ9
Qon4YTEt3mseHnCtTx2RF7S4LDbfUzTqwuXVERnO/8WqocjAYooAQ5XHwXRZ+Vmt
xNt+5Szuthv/325Uk456HsInFXsgIbwRoxvMmC0kAMjeySwkjKDTpRbozovqPtUh
05Csf5u6nDbxFBHyeUxGuqRLuM9srSpL27pWU2YCmQ+ch3hQm61WLok8PVQdRK+V
9WFXgV91nfdg0/BLJJHiT1TMHezrd9S5aMqNuACCXYwAb4PDQafwJySY6g8vhaBU
Vt+tJlhCtRintgDaEh95+3T9/ZOVAmzyRDww53fwNjbdreTQTXxDPju7tElXDtgK
4FQoX+lJvQIVv8v/OwO0pJuqY5xjQKOeYjTa8t8m71VI+oEIpwBcclEgGMIAN58g
0OzAaZ2ZH+KLHQZB/0E+1mZy8lwmYA/J5zurm9pjLnrvc5jWf9+8n/NvMnPe09V9
dOL6VU2ebfLLaphEdZttIphrDQFvu3FKuz+XTtsxVfvYcOjLirrVZyEJvlFNMI7q
3J9QltuoRM6no2zdxpPi8wHgn63ahQfiCSRTqq1RbEDvMJQ+Php9vgcii/rBR8Sp
mffopMm+wv8lKCHD9U0WgS5riikqphpi+zxsIe903QbOFBDfMWO/+Uiz4f0gXoQH
rXS/8K36bsBo8O5lu2bbYfn3tn6Wpd3I2SlUGWfRkzmcfKcYF3HD9nzPQw89WgZV
B9z+VFp7YNQ87cZiE2WAW65pH/F6L+8eVRgREgv9KAx1hgnZvT3EvOVMZbkNvnhP
/Guz2/Johkf8kZEAdsxPX0mtWJ+tscbPZ4eN7nBNzfp4c/oGJxL1V/p9Aq3vbuKx
cwzdJnO3UY3XEak8JpNrkTgUO9ODpK6eQroGHtW7Jow34SMTCjwRsum1APKnoLDD
YQvq7dejua9eE42Gnxnt9OqKzGIUQIq4Yybel0tHlvvI95IHuQoaUnjCt6dFrQT6
P1MPBg3mf3Qn3b460hmXd9fAVHCVU4vYpW2hNBTNWpJPDXiOyMsZnzxU42WMRhze
kEx6PCmmMCA1SkvYVeRjs0/uv0AQESTW7RBaAAp4ObbqY3+s6lU9Y41ssNd1QeRe
lFMT8vK5RO0AkGs/MAXcYeqICPX4ZsVxBnKumvk447LNMYfGxca39+Un8ezvpraP
liGw+UtohH07DF53HPYcksyWdTJRbUnV6HE9jlcZq1OKiJsnIn+A8kIEOwAjN21o
TjEpo0qL0dR06h8O6DaYIMKqDaCwVKIDTRGuMw/k25wy8Uo95c4+0BwXSJ6+CmnF
2RCg0Ezmlip259XL9K823ptHAjKJ9L1AW5zTQFVssfvelbOEg3V++H0qSqqCcVrY
NBmovwBYo/QEUigkSPOP5fDBSKKHNDMFAwMWPEwckfV/eL52nN6f6TAf3esI8PcD
mw+l4n+R8huoGiFFZZy3aLIDCeoOZHkrF34rcpNgw78aGfBhSwpAveowUZbvpDnE
NnYIOGVuzsuM1aumfy2JHdWiONBQzf2Q7vnKTMM20ZkZD4sBrwX4jou8zy8MZr80
nc8r88+Dd4SApmk4Mrn88RZCEDZX+Pu5Is9z5PruUGA8NG1PNYVKNZHK8BRIB1dC
03XaFo+RKFAJt/VU2Ow0WlMyu4CaNhoDwrUmC3DoWNmGC971p1tPNLLapAvMVgp/
oFUCUCFb3MrJuQfGF7/Yz/tv79QRPGfzx79wMmOBVqw3Pyx4YvEXpZhb0avfvy0q
+lz+Qi0GAIx/zrgbZAmVW1EZ9RMNrS63kn1nRcHgHCwhb1JBsIhJJ0ZTkQfnTYXc
SUk97/yIniAhgmwbsuVEqLNPhD0KL6X84WcaJbtowxgQc8lsacK+79mZaWBucPZj
L5ootlW3Xk0ZCNNlbYmByus0CtoTGdDYZtNo7kOMH7YfPDYUEiV/ZIcomfu6TaYl
m56AF24W4zb1+Le/q4c6W45e8KbSVG2M8WbAH8iZ3RSt5Heqgl++c2RHfiXaLeFo
GTyciSCcOUGvfy+FaBht7jeqFBcvSzMKbrAjJ9MyNU5vI15xKS5uquhubNQk3FE2
R/ULraPZI84iE0DOYW9H0FuRXfs/OQJFXl95jZgG1FNs8s4uSPGbBnnofV9qqr7n
CnqUdfNU/K4Ln+hcLi6zYNfl3RgvSDgPJ9xCFJ88ZTrQlgEogOMRBO3CXT7n0BAx
ukY9DVtqNR1b6XSw2jSc9UsSKP/KoaSUU51zOwbYV+ebNurbxKvtzTx9mOmRPvyT
ZgggPA5aTjrUvS9djlZ25xZicr4GscqmSVfXNWtaGcRoTg60jkCF2hezyo4Ztdkb
fOOqI3j0Wmk0yJmkme82ezX4i2w6tS5a0xBEHAn6JF4mouOratmmtok1J2tZIRCE
Cu0JiAkjk7SrrtmTikySZaDOCYfG2vR/7XvCDC46mK3HxTD3lK9AvwSiZYwX7GIz
TFjj+92+HMR/qIUuW7a7EEnsbPZfQBw+ZtNqnfOgcbcF0Fq4MCzyH4fJS/PtepKT
qHZR7djf6ntc/aVD0NN1WbnbcsJnKI7OVIey4lrcYWZy8T062b3Ywc6hFAW8rTkO
6V0mBG8NZkAhuOUymXMQoVsdu8UuQeubPD6LoWdlr/stq6daqJRfutpdltT1D2Qj
RiuCwPODuOr6NEEhFlYHGu3SnpCr85C3Pv38na4Ni49xe1Mp2jh66Cik9f84nkU1
OHAvL2erkJrI1pFd10maNHQ93qfwC3wjQ4GtYYBTIwYW4XD8y9qoZH7aqGumHJOM
w1OxYs3GG4oJiwKZt0Xh13i4w2h5EjwHV7QeOc1SGI8akTy0mHUAmUl3aTfDU3ca
uM6K0NqN0RFhk7M5b6+t0CdoDSbTccZyXuqXlMAQVZ+O76leOlml38ppqeYnZlBw
4LnTxtueeE+7jBTKeGOBoOPh1w8ZvXLBvm7ikt1gKVEBk4ZPdvMUnJAo6UCKGnHt
ofsk1s0gLGWqLrg7U2MDSqI8i/MwjtoAKOzE2oiM+hd5ZZTT5RP4VZJ/z2KK1Pja
YhHTIbz04Wi+79FCYqFjMl0Po7i5i4iQSYtjXDeinhdj8AGXryWqXovEAtYUnMwo
XZAK6IuRMhYjYqnyR4FYrvLi6D85W0ja3TaEANCbXx/rlcDT/i5YqIm7iT7oxNT7
Vb3AjLEjq5vn8EN9lKA5lMMZrxCAKmTkhIOAZUHocUL64DFO162Xpomsw9tvb3BI
rp0cKoh44U/V2weHXQZ4hsCZxpqHABOQHgqka4nmUfrecKzOmjXMPqzFNbV2qLgV
n6JRTbOjE9ZvTZuO8vIoq4Lt7cJ2Z0QqdT2XkS0Bp+mdU6QdndgETuxVe6G9fCbV
k2DuZ3nsHWc7YcCs5foHwzazIKobqZRcjOYtpeUc1SSy1+8ibcdpJj2hHXuQhnIt
f1dqt+zmzW2W99Br9iQiobUGUGPBBZO0AyNsHWjuZZEBLmcJI3onTdgPcfBLjGBu
lRwVeRAuchGhr2nWqlmvK3gDDOsMK4DmCmFPNT9HrVHKQJR+hZEWyIF9dbOFxVG+
5XAdd32S95qWRJx0NLtyVvx7xMvupl1mobniEgn4IkhpDp8yfkt4W7l1sW4t2D1B
DmvCEt9jzeJp2ck5FyiKkEfX0SmnKJE1wWB84ybasEQyjEOo6me4X5IlFMZwFSqV
cE+RBJ6gCYjpvckQwykdklrYaA04Y8ok1OeDSDPHnUKq4t0dnGifG4Zt2NsmdUfz
dBQ/wlDBxZbwiByN2fSG7kRxTvCoJoPmcceysHigYuAFSTRleRwY7HKrsKFaXkLJ
IEbSvZc97wifv+NtgauRWz4AWQ30d6geeEwRM3uDYZkOPyqiYUnPuL+cB9lMZo/S
H6osX6EeGhA0dOUv86d+tYjz2BA4EfROX/8FIzC/OJfRf1UaPQ1UazzyxorbgnaK
eWzdf4UjgdizYjaZ363Xe5r8i9s+a0Vvhk81ORRRnDVXxoPypYMlyvCxFSBK5xtP
W3eIUAAiztGcneZ7y5wrVg+jzlKTSH9uAh8DeyOchAkv0wMG7SUlzJ51dmfSatDs
VPFQtLEBNF5NS7gZqiDk2shV+8iN8/LX8bpsTDwhWNyD7i85jWcd6ILprRGLoqYS
7b6GIBVOPrgg0PeLhr3OeJ070Mcdy0B4TQqomg6R2YBTwAr+EEZLJP0Em2y1MhZP
SMEJ1tCkuj+psF94yH+NK6F2xgeD7Mczj/B0/SHHpHjrIvRqdu1Ey+sOywoIznG+
Y/Bmno9PYEMQsmgEsrJm+5ao7FyNOEBjaUIJ936YMj3Ct0c1ANBD7DQPUK0sFvEm
nX5H9Gr9wxtXvlz0hd57Ve5LA4DbajApZpgJfoFIy5Z71c7XHN55rnDEYZ9CtCq6
NCxMyUxEXHtE4nolV2iKmcTZjCXZJaRJYAjAmMCwGzs3Q991Apjp0HKfBWDBbnJ8
r5s8/bybyQIylaHoA85hx2DBnbau06QBfYLZf8E30PeVQu7aQwiiAs+uBO92/xDK
HzFrfWAl+vTfL5Vv2fSh9deSKm5xEKLgura6paRFV/JXacILsq7ckfKwUYB5TnMo
92OvuEr17912TZFn9mWiav0wh/FKbEoers1sIaR9JwtbeEl8Z/TvKWxmDP4AD+vU
mApFUQxNUjGOeoaO/DZ+6pvOpRN3vtIRfpj3QOEivXOAKZOBTqzHL5ZCvc+pGtXi
o9slJ6eaNqOZsdzL8j3QH3GzFbHlrf04qMqCT2aMcv+fW0/aasmlppopNm0K5iPO
ytnnmktoKEkAIqMxaBh1nH5QEqO0rc3N95gfjxbb/WtPTjYxBakcayMuq4S7O959
p15NN8xX8KwwNw16a9lU22rNr3vgJSE7EZei/ldcNwjDzWmfECX3m3FNFzN3jrFp
LKH8a+tk89QIDDVCpYiVSj0seN1CZ+PgYFbyE7kEiF2Bi+BOQbNif9SuE1SYYXbn
lUOucFraK1uPPT5PWFWcYL3YYCriEN3tWYEaVVCYhod812cu8Hc1gLxnzM5KT8iQ
Lv5f0KMVpVlOR1VYTxWSEpoRAYVFI+hvGJzjnQvkPH0Sb5SYJ4hcoTh2vuYdbRMl
tRnfVIhn5xJ5HdFipukoAhG2z1HcPmAxDb2z3g7lHzDGVYIhvHbIR0UCnOJSg6G2
iDYkI/A+wJXg461Y9kGcO7nTR7iwgmgm0sS01wxgpcyWTq+xnGWi9JZgSYtl7Po9
aPnIsnAS1TgeuxLXAjhGgQ4Za35yfCVo3d/g1ga16NYSA0aOUCv1C6ryP5aCP6+T
RGjI4nwhSFDX6sxqCDDzvwzBfsFmaFKszFiKn/EDSmPTmDDuceStcsWP3Bqq1ooq
alAFDIw5XFqIdi8g6I7qgTq7BXdLvCWzy9/UMYPUnRoUF8K5276mIKRabsMlYymG
0jGblUj3OkViiL3178xM2mqTnErgjq4QPmEx40cY4khv8np4KzQQXk0OO5Ct3dMZ
/RcNjajriJTDLPBuiHI9a3ECYmPuxD2a+RhG7O4/cyeYhbAjhPbQmVhOpl5Ri84F
AhHkK9lzT8NyOcfXvdXvGwo7N0kFWWZxAx6HqNu5rXjVX4gLK9SuH8LMD42fDqnv
TS3UsY2E8ym/l5Mz9/yI11Gyf7fwu5egTZ2Je0/bFSMWAlTPtQUn84eYIQ7My0kl
XkXM8cag4ufzCjivyr5ICn6TSQNi/CMrwvkYL7iFlGb5rhMC8u1kR8DN5JWQD5Dx
xue1nPdZHEg+uN6MeVbiLzX/pkAfpy/KyRrfreh9U60zXqwSa+ZosSW3nfungXlj
00xvFn4Z00sWenQu7y13UV4G6CAPNp74DxpVMxHX1W6ZEC4qSycCF3dkLrIppPfb
gZjgbi4+Hbv3uoU6dxbG8e3Z+wsT9ummG1jUG3y26v4wMDncJsfoct892aeKAZZy
MmmqCBD1ncuHvZSIB7whsRpzPGXiRfIPYpUNLxiKM7HlRhsCBkEeXQZnUt8AwAmm
8riS3nvVg72XHifbBm+QFRd0FBGpRiCZitws3nxu4T94bCMrKDPSRMwb5ZR0Zruc
HuLipOf/Xu2VZgAVNP05SDlD03+CxmXjA9Va3Zb4ucEL5ckJnnJEk7nfeKLZuY4b
ZgkLwptA4KVfoxi8WeSBv8ns4R5PpKb3+8JMXvbH1g0xnlFYaW+QZ9yNziR9smvm
hvv62+cJajtr37rIuv2SodgRqor9pb7EUo7bEBGfvRlwr6jRcmScW+vWnaHABDAb
abDt5gL5KmIkeZUzDvXt2kGvuQ1feQ0gQp9OJTdNAgSF4SPVUyRpnQrEvfwzA87j
w2XXDI1E7LH/PHT0oU0TxOiVrpuOOqA1p1JoGpQYFHs1LNp5HLw/wsbEq+cTcHJI
2GZ6C0ptBdV/eyjU7tO9ynb3LA5hhIDM1PQ1eWyzcudihDwenQQqcP3ukCg9k8ke
MFP3LNwNhcwNlU3Fmho94MSvUWYiGgyOrYUDZEQtiZbICuI4h7eo962LqEBkAd8+
n4/NPSFrjOH4ORq57ROPwS9jSmKDG39YuAT3eETwVuVDh0L9TKOLShledOErE8+j
dgg2yl/prGQOnsKfZrD8vjp7HMqlLm+s38+b6VZ74bWAMWpVEHMNbCDMu1dkpPiD
zWkkY91k9UranAlsJnOmwClO2EKGfTxxslk3MKhnZ/zrUAB3bJE+kSq1yAFU5uaj
8me2RBanMtKUs7/kV76JzeJshI0259PdUiqkHO97PiSvSmJUy1Kltwv8cO9WrRws
hEgOw1VpJa8ZO6Kq/p8cXPJlZ8qvhtBGBb01uBFrKve6BwxrO5Ut66dyyrNtsnao
pJEu5mdLTXZ7z/ASzWobR0xtnLmne0d6Nt5eAlbI+0jAmWgVyckl40MUiIPOTfFY
brM17nCEYHhIVj5wUkZOxJW//PqQuA553n4AoVl0tdPi9ir8ypZXmvoFskQtsewZ
waBcINOWteHnoyqFZBrmuA==
`protect end_protected