`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
YATj3kULTF7Ty4ORuRfFpnT6YIk4rUPRrM74bVTnc4GjdV8oSnW5PtQkMCLOi558
1V+/wvDfc3y0Z8//ksX8sZm3JZWtrxUppw8c14g9Y7owiwp+JumRtO1zuk5xFbe3
0MMnIxxoTKLhyRJtAxElG8sbx8N21OWDGiOk0Xyd5CqAmk9dcOIbxzMjW/wndBXi
maijUdqS+5KiRCM9+Gsp6k/iEAa2LnYTt4WtjkmDD1P5jZKsiMgFck8WOqLymplZ
ml3TTfn1UlLNm/+zD3SFGP0kABAiUT8NK2xBPQ5UzQ6sMFPd/np8iUZ5u4QLTWOZ
hTrU9OSX7lOvRUo8pJ9vPg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="BzW6NOo8eyBw+CxsNNo4wIDxODIsVe0ft0K5tGuSUZw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
DhjJh9S2BY18dG77XPz3hsiSQ73+w0XqfJhD+f+lIDHHVjOB7CfC8ieNRTexgzn1
5W+qoqOEwenoVQtit9u3XViXJSRJ0wfUC5a9axblRNyD2mUbyfH9+f59nWqGkVOh
ieHxkA/DPprM70F3APxk51m7/gNSLICSvbONgLGndWc=
`protect rights_digest_method = "sha256"
`protect end_toolblock="L7NTNW/5Dqy+2kJZXKczEa3js87UJ8H00YWI+92sDHA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36704 )
`protect data_block
6eHODtGLmq6ccbB074dgNWpdzW45i5jL0Nzx5wwM+RA0eeOHXxEV143NNyQGmZjT
bzHAi/6AyRCB4X9z0c4MjyrZE8GF4crbMH4T59xFHqVrQ4zXCea5w0kG5yvHgpKo
cXWo8LLcsQOjItIP6iyF0NmPhoI63tkJA52ZS3N00hFIUSoa2cZyhN8VbVXHVXas
wP1hpTYT8KElfdmrO7iR0SAuBb+SxMtw4V4NQ/lsWex3nb+H2Lerz1MB11ZvnVpE
g/SS5fVjVOS6Snxs3CWpH7slOsJnHkHLeSNA2Sxnh4P9H35acmn+eiy9lQqmEFH6
5yy0euo9+FcnAIOYRtmDCi1OLJN21oAWRi64eLrIQR6Moa86XWRrEyHyMnbtBfk+
8GqE29DMVVAxnfNdJ7eAUKgtVDgQnYB2rudvnKZ06fuCK+0zKA2dL10ADw7az4Ai
zfGRN78B/k7XFil5sNX0T5WUxuRPT3xKOQISlDfKcjuaqDGw9wK77CTopvByO+aZ
dEKuDPXywAKwvWkfB1k3E0lleMYcXPh7ABlwL32ckss5mKBWOdhDltNrp2SlAiBj
qzFoV+SCo9R57J8Uh8k4bW0cpFfJZ8xH3SUVIE9HMtEFF2zGU6bt954cN/bYeNfd
TiczXRF2IYGzp3q09pifb0xT+KsvxPfnJmv3Y2xEFWX2Lm55LGqTcAYYkDmKXmA7
HX9VV+FaP0njr5qmR9Q/KusLRGwHOAl7cvV5G/jFxLYYVrVCXyRb+eHqsk+wEaBA
K9dg7nskf51bsDfdrPdr8bPiRK7ZNkggCIDOqL0mwJsuuCEFviHxaCS+dp1nrOkb
YpqJ/PY7I0TqNvTG6gf6vYMftGkhWUY9SQ1K3LjlxTi9Z3xvzLGskCr2GCjhKr54
WfQfxYKQo7+0cAXf/PU2vg9NYA8d+kKQ+QapNQOlis2Sb1lKU/w8zN6H03zJLSfd
2sJnLLEVcTUUcThe+zxzJ44/hNfJfw01J2jT7SMKwW2uc7q1bTo6ysAQ9kQ/93Sh
ggNC5uMsbNAoi+T2e9eC4qzokJ+DtYSMXzZIlQp3eBAlaY9sMMbav2cQEvEAZO75
+Xr3r7WQs42xJrTcMhyWEy9iEcxi5l/g+zuUAPZCiWanOLgneCrlhsGyUfx29wer
VgekMHSIWhk5sOulH00iJIZ0Lw+3jOlwLy91H9CepQbbFRlZOnQcC4NDXBc/7N04
mP5Ufxs9ExQDSTPN+n34OJ6OxTgaUQMsT8Yey5dBcv8N6r7/Kpypq4zmhIUM4vEu
1XnKvPjbDs7PfqDrcEthWNKEQ6xK6wdampibVYEJdycmYiuX04OoWfuoyC81f+Y3
fib4qOO0t+Js/AFS79Sg8mxp9J570xqhhJaFAw2e1iNMBbgfY/iswKBQ3eo9qJEd
Mo2O+ua9gC80cmuu1rxTJTGzJn8Cn1FAnHumEdX9EDAvA45pNZ4Mrmaady2bam5j
LyzmQZeWlf3waHcYplXf5dmoDfKC2D04nliIUZWKUtbL/+zhhmCK3xy2nk7tbC0E
HbISoSWSyz2Dvw9+BWijnm+gIik4qWJ7b94qYir5qONONzBTCd5qcd82kUK+06xG
BKmo9/Wg9zBOvmXSc2NwBqRsMZAwzKFmh31tBlu9oQHslzv7JE4HAeGZ42j4mLNX
fyfzPYyh+/5BEIdvAckFDoakXzsbTm86u3XbbjXNRmmYplvQtgSqJ7LxUfWVlkMB
kC9pTJvq83TZIyYxg3PrLtnG8uHzJvcs1LC7fjbp1ejb00pL3q78caMaMsauwDxZ
A7/DeCZyF1Z7xWbioBKQaWeANilKyN9FTc4QzNOSzGX8b64Gk9BuqilnBOWddI8a
QQj6U1xS4Zy1WBm4A/gdR11OyDjlnCkqAMULI+zf9L9BgLGR+K1lmpHtga+7lq7j
bdSJyRLHsty6OrEZN/nCJ2HhzG0i+lARDoKsh2zFwlij39eRkZQLm4zAVFvUPOFh
HL/79LS03tQJFhStVXMHLZgiIc52ig8COR6VoTP/YnsTUGma2EY5pydojWJig9eg
55SxPvkAOrD99/Q1x7feUlwfKQPxTyQgYW95pKuO0b9hV4JDN50C+dAII0TKINwa
P5W3egfjLRACJ7SDbAPsxsbxkSM57BitQbypqMmVMwu2TpiDp3BCUCnYkUJU/aYm
FrOCNNOn3vQ4c3OFB/G7VDT16ZGOVrZGwn8WXC3aCJacrmj1yWm904TgLo0ARiOj
qrnOm6EzgaaA/8ap2gRRiguMcyMSHL/RWm4Wo2cTa7MICS+EEAdd3XMh6esxa03Y
z0zbaqilxiJneGiGAXk3WK9XpYFdcUD4XtRRL6wtoaai9KN4ikIHz7AeUSsT38As
+vnHJyc2Xs6DbYZ2UrizeHyvm7xA2H/paxJjGsjmMZK6K5uyQ7tnPFEelfCDBZ4K
aR3r6/mfHxO9iLYXeymLQlV8DlGIAYbWo+L9pgmjvb8Cnx6nHG8ON8OoblNnDZXK
uqkDDsAoeMjewnJshS5h/gsPehVuBMBUS0rY6McKmosROMeQZlpqijPDMkL20GWy
/xj6eA6Tht0fQEe5RNmPPIjhJbW2NuUxTbaqG8nS+c6sTagTElN8L5QVwAFcQlZ6
3OkFUq/Vv1ayccc59bD8l9vVjdosbCcHxUQesSt2WC8H0nsXdmWDdItKdWilIiWB
8GVmjgbxz7l//IdLWqy3qizxKjiF0jMZIQt5dU73vtZpnLndBg6QhUb9VfPdYVCp
+MvhiRyg0MXEc3r7xtoKNA6EEVGSx65xwf0e3KRTmDhdkbRqdq9qfj2RMBOkAZwO
i0K4lsvDnhTk00Hs+sp9Yi1dYwWpPzU9+Mr+S2VwjkDaefgy3upSlhHxafw3DV14
2AIIfRMbLEfi1C9iJFFKBmvL4stghDwtVoA171Ix7v+phlj0gGqLQgroQQt95IMd
MdEyHt/5TDS5+d6hAEiAT3woqzCONDJSVEJsrQb2r1OeoHmsa38cOGmPVZBQKipi
KGod3lbDZYwv51wB0exQssSIntXwyb4YB94nb0KW4z/cHdDL4kJxoBgWPXZJBOwS
qOBm5OfFKoyNBs/Jc2R9IK7zKvNw+/zfvBQ6CdU4H98pQZTpRIYmWTmjAdA3Cb1c
JrIrGhkar+GAac3NGD/tigLzpnsJFQG5kXqdqx4Ozi5Y3a2ChnV2TymCeF7hvS8n
U31oJQ0maWlDCcaS0XRKlZdYZz2HCTQWwGKmtldSGDvz9etBbCBbCfGJRqEZFEoj
pTEuIs3GQtUkRlnZ+uv5Z4FrUTuz22IzosupAjGQe+BMN5/PwLep6a0dLtgiotQL
/enyvEct/Xv5wYc/fwe473/LsDwT1FnOHkPJiLlnlF8e5sQq4B5k9mzjwinKn95Z
2axhkjjBbhin/ghRPN+CEWpbWQSOujF1I/nU2wsSR3afytB56OmaWITrQ7j0cG6V
MSSTO3UmeSjr4EETaqu8Ei0RoAEw6hJhdasFmBTdCC+ff9K9AHbWLO2/3FBeJ7rP
NvEO2Y68LlOee3pmEKqdxbgquJi6OF+1PIxO4TLwTJFij23PsBEq4OEMGb55Y6oR
KmsqqSRYfuFyaN6ID18wpgaU3SWxtt4KEkhszBLK8LmjIml9QDC0vpSgqgc5epLE
XWUMxTAf1IV+wIrDSUoGQcR0mXin5vViCcTKH2InULWfm9KrdGAH4uERHEI6K2eh
5VFHoISZwXAmwpLtQCgNYyjSlHM/1tG3GSQGtvw/+mt1iAnfnh7rjzXww3adcc/W
t4caouQ/ga3F8PMWeewm7mlSurBYP4wGA8rQrF7pl7FS/OiL+wcRrCVEpI17QBPn
OjJb1c/YRZI493xASwouuXD3VnWVpom+cxZ5qqg15qgLkV9W4sbCdtMvE/ieVrQ1
4rOMd3w5vPX4fHFpGFoQL9weOEahl8ftT1Mv2iyFjhuPNV/yvidOUC3mUhdMc8zh
qStryvzT4HBwSDVwWNK6IzwCv2pznn4DryFy0/7jAAh5LmL3205EM1mwQLWuylUZ
dCug/JxHB+59UWS16+HwLSMl/VzgyXpN8WvuOuE8VqAJe7iMusWQ3kqhLL8a9GNt
v/lJ8wf+H0zfwoRwcWIEB+TCyWr/PMmE+oaiawn4Tqlstks4k4stMboEFLw4hipN
cZed4tVBqPNAsRHeNLNwGUjVZQXernX55JuyTA4uwf9529RZfnfdby0pnQzS8Fk3
83NTg8VrwrmmVC1nhUGIUqH3+UuslHS5ofTCC++FuaQtwpQp4oY1N479O7IZhYXm
IaWP5I7QJABfInQBgA6XoimnxKmPWI//zDSq1Y0DjlasDyCBPDpQq1o03o+psKZb
VC1VPJWXJtBncD91yGs+5h71EHuTuRdO+78qd3njDc/x3Nqe2dV2sPGoVZmlEovX
Y6qpbcnfrGkFlvb5o+0YVUulFzBfsGpl1aXZS9hyRx7f2wiwO7UAW96/ZrdI2RNl
E+HRyqc4+dt3aaSUuHVN01wO3lR9iAjrtSt568YA81OiwHi0c3/sR6pLBApvsdf7
xHOHWEBg7ykMD3l0BaqLcuzT/PaL7AyiaC2lQEIUqHBdIqz+bwgQFuTyTnWhGCKu
ywYwGaAdmhX6hVImN+LbIoIjdEAWT5HKIZVlZ6gq8lbGsl9ggpw9NCDzqO08Nsy5
TSlADr2tWfXFWubBJ2ql0q3UzV2fH/IJlQlY0k1lfamljkY3d0cFNWyPyshYZFL4
PnrnlvdPZeSHKYq6HIdhg/TwTMilgyVSu9krAr3DjwqbWC7pAVxjxE9sXIsNCDvO
5ghqet7tJcJnMkKAeVBPbgZJQM6AYEAlMRQxm3oYBQYUFBALYa9w2KXDIP+u7llh
kXfIUCv8sxpplbi/NfG4KpG6k2cxALA5LDq/e1LmLKCIc7opFHyE2dFxRlYBnJqo
JhxxNbgIlmWFfHlNiibUukr9rq+xzj3PTWQPkW2R26Z/9NBe5hRdvncwX6SUajls
LGHmFvkbFs6W3A4wH/Vj6ARuQSB2IZJyqzMBMYW1xvxqr07bP9/h0A7yb62JbIlp
gJfeRLqZSMpjzR5xYjVFeRHxigRBGuhsMG8y+NyRdSiS3xC201XGDGq+WHzAH1MU
huZxyC4EhUhF8ipRn6Y4tmKJ1X1UfDf+CfgzmVARYRBokqML4wjv93OQANwG/6px
jI6v0IEs3FKCkx46oTAt8eXl9lMPmq/dITLmHm67C1eiuvC+ejzBJX4xf7Un8LkK
+gQ4/Z15FrVxryoZ0h/0acTyagdv4bqZpbIKCBsMrVZRVnEHrW0Lx5v2AZXv8lZ7
g3vZ8x/CKRgeqzBO6n30AyK64PWKdi76ScSTbQ/AdIiGykWrQZu13xuuVnDgLIsI
Q1b9UfoKLgLJTAF6KfVTnEzSCmKowGKNW53ufAYnT7akyjCvFMIDGr5afbM57Sl2
kMt/6Zw8JXvHIzUk8ilGjUPjYpvxUdQCQ/u2qqF+/MtYp99X39F2WXaVPUyZbll8
Hkge6edr41xnG62i8pyfGj5Zj+rjLsysRbWBFoSw179nTBfuLTO8CSe/vPk0prti
XNq26TyMnfzFd+hTn48V5ozxgUgVBdLDbCXll6KaQe/jBhaXco5YOP6pW/nEx8UY
giAUCktNAu5LLWXfd89knEDZaWY/RxSi8AQ745kUQrtv4D/7Wxv41+LXMPMcy04w
RMrM6oeoIUB7JoknUFkEEFLt5jtHacQtVSuAxbMLJpcCEg0MLYZqBxzOnZ3KG1z5
e0jrr0/vtPCXTlwHWytX0IFwFj863MFVMV6EgGp+Yav7jxYe5/eCj+B8nmN5OVr5
M4cqhtwjEQXSJ5yzAAiWkJ1lIhYb5Pgqx59k3bNKdEj0dzxHCWFc/w77Ms45fBwm
NlPwOw/4GbwViKI+T3i1QxjwqeSgcUqe7wAU4PQWyxgwDV1nQFaSYMPtYP6kKb70
NVYFsZ5kZewVwfm11fC32A2j4Eiwi2PC0I8G8QeAjJjTL8+S2+VgaPC0nqGMqf19
kCndS8jK26R94lubydoNUkOwzjIlT7yEtiBIEG7Pjaf1nezk/J78NukBPE51rph7
DtNKKrbOY/ewh2PLZn3mMkzLdV/SOi+Syu5/SoscGf1er2nYzx63eEMzZPxn4JjO
XI7jQkDYBXQ7TcKmn9bJGQE6tXH2hTl5KQ+e/E4+XXD5upd5k9zfylF6RghqJVNp
AHgfSIwnGQcmIEu4votocnTZhUQna28pV3gDS8BixhGtNCPPRkwIA3LT1LJZCi/y
YIGZA8OnjNx0q5nKUUSxPNf9PrK9XjbFTI09YzrTSerm6YhwpyEfXwAW26MjIwk+
+3n3Ls7VlTGIzisAqtpRmR3GLTnpHqxAqoQHXReDHRiD9woKOd5ZXP5CIWBtr7MG
PZMKp36yHJ52ka6fLB5YI9UIq6GGsJmrju1k6RDp0tqAV1Kuth0eheZlfwc7QYxz
kOPoAm7y8cHB3rVMZx86voAxCaLb5UCrSZUpQQib61OfbsN1JkffX91SDWZyaZWt
DrXnIOU7FehX+rZHH9dviF3WcvpVd8BmvOTLC2slO4MCC/QCnA3iKYwtnbXH0Lnn
7zPZylpLZe6iK9Bo/AeQKepOtAr6rZwkmlu9cXsXMoDLnyWb5B7qYCAAZ/f7jpkb
fhcXs7FqbyYsUVAT27Dr86tX/JeZPJ1EtaU+ioFOuw1AvAvVeQmkOb+nHdGGgt15
f5JYXLdBDEPvDVEiYxXOz6U8UESN+OFZ0l6BisB1KhPvrkWY0xAzebXVrtvmkrSU
VyESSHuKoQXKoS7muEglsMTak856BhMJU2M2JvMBDavuHq99wk0r3mxwNVDJAz7U
bWfJxDUzyXmUZ8i7dsq924UqeUxYn65SqDs7yhmGso4OdSGgtYXxTe9LhzgstbvQ
vd1bAv5+wZvLbcvnhdGzZyMq96tuSssvtyyrq/RzEFbjL9qGPbrFVrQfsgyad7hm
QaGVKFF/BCWMNW4ofM4vGAQx1CgxRmJRbvHRz6Uhj+t6xCgRXQ4TYapSp57X8Kss
edn33ND6oSf4qflhw5VBK44UeXkPP0WzJ0JAyRbWLDpwxbMvM4tdsQSzvMzRJrHW
oR84BgBELKUUGdJEU30K8Itr3nhBseL5d+vYKtqQyANnmDSQ0nlUouGqJ/iaRbS4
wwf5BYU9f6vrk5wEKO3tEuMRuat0LeSPvBwwxXA+Kxfl2zHPLR8dXEyhfMDOm6gq
12Nh5rk8dCw9ysPi4vT2JyQQ94gDPHTRZKmMR+HmAEqqIseOn1MxsbEZ+1077g6Z
poQJG6iUQALfjfAfyyRIPGVKhUM6QENtN22kATmtPaXdcNEbKrL3Dzb9vJvRGU2i
OvFvRfgFHYXz57gaaZ0vEDnjUuedjlrApMBNXZS/bNXdZXjh89a9o6ojd2BH3DeW
nmZwQThzZze5p4tOYkF8TXfXYK7XxWuxeeNZmlRQ0+TlEzJCHXTmVk9iQaQspq8y
p1PrgMycN/un92Zdemikej2azg1LYgRBE6sFCuBJeLFjJcK4j2TlhsKQozbNuR2+
vr7vV/OPNXDMe0FaEGJ+vUVdCjs32RnCk7GCjKHXCFN6FKGsfDmvVH7k15G0mYCV
1N9xLV7K+uwum+XkFAY2GCmTmjrGD0VBaht+pQhJOUFQ9BhfLf4I2XJEv3P/5HLb
40IRPDOLDo5QLfaqhRZgm2UbeAyPBKEb9MFe3KIgHct8CKLoF1lxQlsGPOAQ6kq2
cBxTbEPP6TxFx9m8wAqUV5VGqdZ6BOILLEsXLz4FR3Nl6No3sL/fWuIgDvkd9Zqo
Bib/2MbuHqXV/pSenr891xdW4xArVyxzql7MXCqRD4rZfYXyoTT6Zdgv41BcGF6o
7+R1asKjntQO5GUeOAi4jQu/klg1dygfzoxLDuuoWPeyg1R4zkw3wZmmL+1oKSQU
HbpvkuL8f3eEeGP8gW06GNhsCpj2VKeCkfnolXOawagNxaPY2YuZJv3ukaI4B+70
a3c+isNGkyjdyDmW1lYq1I/2UeqLU8a6kn+0RgR8GVfs5sb8lZG5wOp5r49RM1cu
H1W8zv9f5G1ToikWYGBg5M6BNTIyOpTfzUdl42BrUv9uI5NdynFVwEeMSVtT11Ce
cYjj2M/b5vgTGpp3O0tS/WGAUYilSAY7pINDJTUH4fUZm9Q06oKDvg+X+8zHomBv
Bylvbfd9RMNHCPagBo8GLTwbkCqh1n0INTlFDO8wZOcVri64VWmAWeoAcSr4OYcI
YNXitLsfPKd2kC+m21xtAiMKhY+hF2LUsTP/J51AE0kOLLZSMbj8epSNtDDjVnQ9
+kwvIGong18Y4U0PDI7h8r2e2HlFls2EDHysfrFtlDwvP19EBsQ3YZHzjyCY3pjC
jVtT8WCNRlnkXzxwKqUs5LLDf+hFYSckON7NA8w7CZCMdzUtRAzoCS5Fm/38XMMh
1Dy9nBv3GwlC3KJCx1PIPcA6bwv9iXeiAT5IR6rjH9r2o/jqz2cvwKbxiL+DJfKW
Dv7rsxmmt64L7wvRhfiqz2M6zoDu/Y+w3SVpgp12no5LR//hcfnAr4Z4xzzk/IMZ
rWJpzc9KRIWi5TSmD5WOXcYEJ/dIzPfY+Q+gbDk1oPGM4o/ls7jCwVAC1fbBpIiJ
cOhC3fJ12yRQHiSVvdZit/ZYt0tuYzFneit5b/1zpy2y/oMmNQIE620Cqzk8SHpz
LXnrKq97askil9te7/Y1wy/bEpl0qDwHlqKHgVtCHmXExGPx9v7EUBOtoQy0/CWC
jPVs8JGrr0NPcDrrjeox0U9NRMCYv9AtiP134JDLB7EXzELtVFNAiKas52YAbBDA
hXQGILTGoq1UjvnWgUe0l3RU3ccVTSysTKZTmeaAql1gOkjHWc1D3leeiAHKbU4S
xEay05gsrtq28vUHzmd7T/rBzZ0/J4WCiJyW68ueoFne2xD0hyakU0XAVtIlG4S9
/8opjBjRU0UWOTE3AHIKDCP63JroJZpczPY9cvKH8VSeQRqXJGUCjX2xXtrD8hog
KAxLa8ucMI9QRrHBQvQEi8phrmwSm39RpFSfjLDIMLjNqxEcsgoMspKUCeHQh5HW
eJZGwX2VQmcLRyL2+wePt6NcHY5AxOHg9ygkJY2yHHy+wcALHmbY2otvA5PFJTi3
ZiGM/ryEumJW1cJUxjO/sRIX4WqjHNkkzR3eD/sC+DgBJK9iEBXiEzmI9lx/Vqq0
L32odsGGHRCuVcMRt/zQe9vc7Ozqa3uCr1Tg5aiO7WIrNFWQQnFtC6ikUF9Cmz31
3jMzkH0Ik7qBFYdFfMzm07+bJShdMxK2SeRTIo1jQZ0sLL8ZnzJtp+g2jnR3yN12
ZqqWWNkG4zhVoFABs3VL5SAcbjiyONmh/9BKM7vdwjiv9Xw231X3NMq/41KiVOan
nkIgz3ZegCoJ+ry9NsGBKoWRJAfA1brEwUR5erQJwXViTsM/wbm+ToMHj21VKnSc
xnbXSVPZdlz++2uJDlHjqBaBDCpYoIJ9CcQ7lKnyeGNAWVnEoRP0u2nCDUa3JHcc
ZH0HmYNbNNnf8777hZQPtD+r4/JcJWH/F8z6wQEhXrUpGUORYw1uk2cvhkZXyLia
Tdz1Bb7TkelzHuJlsRCKnVUO9l8Vb8xrFaAFlIhVWCsdKsIqf1yYXdhKBgXin9st
3h0Vx64ZpQ4rPvNhX0m+9AaNMlsOfeAzeiSzAS4LDVoB72mURZBm5FAF+U8PhIjD
40CWnRq5h7/B9Of7NvkbLbBgEDsU7tPzoEUz5MQWhDf7UOuEFYqj8K22J+TbAW3V
qDlHsvzIsVRhVpMkmBbfwokjF9VN3srVqqtuPTFLldmvV0aQqWntVjpfwa36ZePo
sNSCPvBj/UdqvY6TLggiBSjcfAcB3Qy6aaln4lgHCzG16AGikYBhFjtoKeG05SFg
3ZV3TZSJ0kHspmOlzgrsYPtxokJ3Jy6+sN9oYy420J0rd0MJivUma/ZaflALwZCv
raNlQ4fYJ5s2KHn/uQzfGbSop6fLnjFLv1okZQeiW90ZMP3V3MYp8ksjcbSGoTcz
EW4jX3zBk4pUx95KFqsWDLKN0xeB92g6M+DOvOQODUfHRFGpcwXDMRGeZuavuVJT
dcqW9TDhFu4clJf6FPFN0y/cjUWjQvod0smwZsApXGgGU/sEn0WxCb+72ptm/8tR
o+Nxy2eKahwUnxuct8yn0YoMgHrckDxb/Y13ofXf7krKGqBCAPqOyDdzdnnV6SfN
4svZp4OsNI+5ji7+VArBZZWmjrl+vwVqSuNvfkS7T2Cyy5OIA28zdtcIG+uiPkXM
1UknIku9S1sScEln1MlNF5wG+S+d28nQSZx0d2wUrHgwnqGuZ9v5OxXtxPfLSoT/
2dqO3PYU2ZgCDkz6VZAHdleI2/2cdYcZh++0RyER06+A34+5SrCtDK+pU99ibT/n
Q6XM0a1jfj2D15rCDAR7WXrK3lhTfpxKJvHayIWl8MJmEfb/akb/FXVnTX+P3RzL
Rc/h3KTvieixjNkNkIPo//058Zi/uZUMKVb7N6i1DXO+Wwi9BwU4PL1BS3YH48GR
LE0FQRj2lkevyEyweQ1F+4Ui5yxXFdLthXR4XPMmW6pJ/QjSDP0X52xBbdXbZi2r
ePW8yMBeAJBVYOWPDuSWnE3/DOBzUjQ4Q8Y6LWA5zWATn+7S/v4XFA4UZ52+jm2L
3O17NUHuvHzIF4/xdt17jNf+dee4Ix3d4yXHSvhXdQCunKTA1yu3IevKhwiNm9My
t3WMqIPuWO9hgZPryZEJ06NlvRg8FOl2vDQALYCv683AKubtW5YXZ/NL4vQOqMBG
ry7rldUGFHb8/BN5Pg18mhQKoosudpw4wUUo/r3OQVzds2lDlQt5smphbfFsGBzq
HP54COr5pfaUq2t5s4nIw0efJtYlsOlT5ECArbvfIcvMXpK6xns8IteTdpd9LBzp
TUqW4Ko8GM0Dl9qMx1ru+n7uKkPQnKO84GK9SpmwU2vuS01ZJKO786SyGzhqJuL7
tyVCEuKQY4czPm0UVjJIBjgx2UwiPDH7eVb3i6fgzlNwtguBCaKLMaq3ND7ciZTZ
VDIseadjyE5bw3XEXZXJHucUO7Rr8VQvWR1McFS15rqWJR3BGv0YqVNY+ISSXxep
CykUJ1qO6t4IhNGHuJCBnbkWQWCiwcYWS9ngnDRyBauvuvYEvKaE5+r46ghDWXJt
sf1jV79tf0w72VwVbyCybtNnhSYsXOHb6wkNiWn0RTnn5rSEsVfVd+fYenVnvucn
b2DTIMAh0kBku0QIBvg6Gh61bPC5aDvGDM78FNGsTYmDg79SGSMKBXJIpoAMBg1i
vYIbl9Y2fcVinjN1EtPjeSyJDcDu+l+8rdg99rX6WF6SjimEwK3+PJnn2a76pW2s
Ji60IN5p+F4WNhNSoJY0CB8/mELor3gDTocqBCSkIYQlObDCpA+I7Y2wQntx2bYi
9Bgce1DBEagnldO+Sx97TB6nSu8l5Ilmjdk23U+fluw3oVaXVDdEXTMWJuWdTd3+
8AMlOS4ryP9DhAjsLI058YR80odziRriiLSJvrPkSzCwIxdL210+VOJAL4tIiNWH
DMz5IvzUv17JN+aCqUPKuBZqeXIWw0SQjzUCxzkixgnC7IO0pb36w6je5CZ0RdNE
2Cc7JQSixsU66ws5fZHfRsCNj2EO71Klr905XLO14f6IpVIvCMRmK1KPU9P653Zm
yalybws9J//yGIAKpnd3N8ycsuTasg/euF8wilvBU6HsKPN7njs/6DKAY5i5iKeY
ZcYNze9yMjFEgN0BUA1GPzxdkWddMdV/pkmhLFYV1CXqu/1FqJf9+4tO/trbYSea
Wz/iiRX1dI4I6vL9uUUeV4Q9j/Dujlul6QirkXy9NG4Zi+j4JT+o/qJD9lrVG8Gf
r3YA9xjXYr8oAa+k0X++Y5WWKLmnr1v5W8f1Z3qpRKuZED3s3LLD0+74KJoesSKJ
VrZkObslA/aIz/jPIN0F4zHs+GG+xzEnE3JOujHGHNvtf1ZA2Xm0HP9yAB8noJU7
J8/FnqF2Sg9B4EhnOvgxSWPmRirHjDs8qUh0mrwh1qPIfD28PUc5/Etsf2trcbYd
HeX6N+pgIZg5a+Tk060uzTAtafwTDYvc4re5ULuxn2KHQc4sFDp3eixd1ShqQwKq
wz6LcQMy9EByyymXiiz05tPuTJdNcEcNzAFUhn62cR7loWORUt9NS7B7FiUtNsRf
zDwjVPDQ5U7IQFmiHchexzikk9BmXhdULJ7A6zksywqV2DXqIysfEKjFYeoD2Q1L
j94lR8evmd7IZa6gbzujjkkwYQlMFFk0+ygVL3A6cZSqE7sm1QiY4ZxG3lu5l+OX
nkHUWKyNOiCXikYvONIp/CIu5YEDxaSUANhOjECWFKNtO4sjVAA/n/QX7NH+6FCx
NOcdCjrmvDFQBv1zVi2ceeUyWSs+n6U9e6msyYS1zIFbhsHmjtJM1XKNL9mUVk7H
f779CKob2ItqtVtcRot25ttbdFKmCM0XtnyufrmA1+r8oxd99XHrT3bj7JOuoKz5
setKRP6cJHq/CdLVpBTRpQRNrczgVvwQHW4iRV+6x57lDvnrBPcARk5Ih5S566NS
Iae9PYLJTIrDGsb/9Kk6mlE2380GDkzNvuOqijmhPXq9EFzi16a92j/iwyCEUDBB
AMCWcYzJ1r7IS3rWjONebZzHnvcFVhPPztMic9uN6BUxLe81WYWhMof9nyAZ+Ba+
oSish6OiPhOCm2mmJZfnzNfTpyJvWpQPAK8fr3ohFSIXiF52tjVFWcYw2jygSr9N
+deFCO61C6ATgKeoAh2SmIgPU/TxIusIhIuIkXTa+nbQCq9iEf+zVfPdYxiI+ajt
l0SHoaUGBMwEqH4xhyc1txc/7gk49320bC2ptvJ5MN30KvfJemW7AtV0QGLIReKj
IqfsVbvBM34frweWBoJPo/Tq+sU4OvrdbHsK2LCLH+ayu/tNJ1FAEjA2TZQwIhHz
zY03VWSvbnYUzR6PVnV0TEX3oNOVNXSkVtfCEU6hdOkk5hMOIONCxVwmztCzFiPJ
kJsfG32vvQT4elwb7xX4W2ViEpHpRG/tU+YLP0miwMrCq2DEexszNojznwbDnbXu
QFuzdRR6vty2C2t3JL0+xO5plpYNauSAshqsmcIZE0DHOKo8g1dpjc8MCB72tf8J
+U2nxO+ubL+GB+bTZc1VsQeOxbau903v5sOZblyHM4Sv8YgYgELa0S3YPIjdNi/b
EMPDuBy7NkMz/1D0vh8iQ66g5jaqLVr7mRM9bNJUpCXlGiZ0zJzty5xSCzx7PTjv
CpnWcBjO9+FdmUdbB2NiCEWg0QotExE+TK3q+YqEKahL52DCH2Nq50qY4xhtZOxK
REnGHTwH2+litJ9JWS0Eh/JNAr+dJTwYWl73UdQSj30y5tHMf8W+xFH3Ilqi6tP7
u9DYIXFvgkpN8QojRQjzE1gECQZ49oLRapkMcLXTCRKfl4H7Xp2WIEeVvm27hoGG
dfWHXMm1rlHZpVGn1kGKPJOmULhZ+VstqcIKBfaqgEb0AQ/Vsw9zMFDft6IwJT83
ZuoFj8Ls4hFlcaOn4q0yWfqMrIhMTRMZ0mSA/5439mwvxYcNGUNGMbvj5TSLym3l
yYiMyYvoclYhWQisNbAmTeMDauS/FlTV0o89diWnWsJIFlq/l1Kcak5lx3mTTKnW
60jdpJmMdBJJStvYWLKB4kKdLoAcKY2CvP1kfKs4LfeIPd2Zk6+pLvfV6Nw2S2+Y
5eD5cMVquz0oCWBacKiGSrYOC2wm4h2hDv0YBXHuclmzs1kgQRwVhBzutasmCVJY
Dgjv9ip7HY0dAzrckaj0jNVqxZxb5tgRHShIfW7q+SFSRncnScPPwXC3Xaq2Rujm
69HqAvd8aM0a4VKxjM0kJ3+NySLKoW7/k9GsxcfwAXZEn42yu5oUELxhfhiN5/GL
x4gmsZ2i8If2iP0SAOswMd59tcghubh+63dziYkr+CNgOR4ASK8cacPEGzk4ekci
g6v+MVt5hw2OKqKV+iBQP1sNidVbMtR/7QhDDBf8bulTu2zVQVece6n0whsJ2JJ9
120mn/cvEj0Rm/T1E5X/wuvE607VtZO8Uwh9yv0vvQPnksLLiWkSKACMma3lidQV
AbsqmHqlj5VxfdAgUbSNEFEkGfxzjqByzlt+K8JXP8AuPD15h6hzQpcgu7IQLzD6
pxn1W/REyO5nT/8R4BCUkDcK7Sn47ZAkf0ukYhObFCJVSDusjkvJyvYyyRJrd6bx
oHR7nLSs37zJm3mzBMCHi5mCkTDcuWiy+zseXcYmSR3EMpbKVYupzENHW6VA3Ec0
5lTq1NS3kIUA1JDI6iU73wIZuOT6UAYIWd8ENUhMytSVhG0jr/jNqSUvmtybqSc3
UnQcVUw+YdJXHbKbjNa5T2X79gQvARyb7+sricvuUmMcDdksw0+GYr1Pb7nKftqa
AcsPH9EcGN6BHSiI8LNQXQKMVWRJrzrLUn0IDz+EXKRbP3DP0/gTdNkmwv7dlo5/
iPwO2cqYFksIDpM141KxvqNBjSmCBxbd5AbFh4pbCYaR34Y4IzEfknxSa8ikO+od
4nzD0+lydXj255P1oifpu6D99P4wXwN7rgScxKVVDLugKED6v0kY+t7aDdOXnDBy
BxTX0+EoHtMnBixS+5ZUWO1sQUHgma3c3hG4kB2XkNcLaYOb8j4h+e/kg6HM5XS2
WEsmbyr9K8JXuV55fWbRITwGVVIbNsu/ZE8hJ7KalZoQIEhDu5i3RhGWgVyoAZBf
zkD0HfLoUIaGV/0/mpHghQIYzDFcNwWpTY/udMQGgG2EYridX+4ApylzKiI72Mc/
rtyIQJ4PitAz8/q/MYmNPmMJlyVuArIPOLtfAH9z7aUyYVH0fnXg4Yo6MbBpRqAB
V8G0PfBmVC965iyw07tuI+o1H6JseH2/X6B7KgGcOHuWm3b+8gz/Sn29Ix8HMtV5
Y88zL73XP765s1mDRiwpQkzvdHBCMYOKkT77hlDVB7Y7IIoAkhuHYiRL4mlFRxhU
cyx070m3lBZi99SyNVMj14XAHyImQM6yfelLWaiw8jCbvN672ao5PKyt6xuBijNN
khCscBOLihFM/OYAJqmHqDwtPsMI6SqdlrRdpQnDRW2aKV+YEWJkx/birgB5+1Xc
9L5LEwzk3/I3VI8RTHuJs/gJliadQBPP/NJmHZTPcIUOTYGVEhMjJ0ObsmpPEH/7
iDSGV/H5Jtg94if1RFhnE4Gy/KZ1t6M8omz4T0H4AWoXQKp3g2Zm2rB8tvwmxbs/
XL+9QiTMQGabBYRmhcJYYiMPZdRHZXG+YGP/lwoxxrsAH3rBAgHQ1QVdOcQjyySD
f0LVDOhpZmLYECyIP7apfgFWKk3M4hJqKg6ZrdZdhQb2NS1qId2UTz5uRZ/glE/R
ur69AeqALTCm1aEKro9JuLvuEc7UcULRGTqOlxCaefzB3iVrIqJz2WVq/toYWDFP
HpTiOVbynRzj09ITixAhYDOsytG/Tue6SocNfngSvKlLF644waLBvOSjPyYaDjDn
pcFD+kB10I3CAJYRaLZ5agrCeZim2aksgWUJ/GILS3evsnzaFnaVhPHPuPfFBucl
nzzDj2ISLM6lfLIDxk7ePQLeMkkNrnegYRxn5WkFEBOvTKdEDge2PLHeYpf11ZXT
igH6lzaUCXI9eKJlK34ileo+0SXePsSoQHzjDCR07We1MrSFct6TPe4gsIggUV8P
iVZzedusw0sSn1xeQAvtNZOuDk1lkxsYgSiYIQTFqHgwVz9rD64sBA5TDStX8sgM
4TzhcQn99FnBRFpuJ0WA9LEqhKieZh0rCB+c3sqz6nPjoxodTESKez2LMuCTIiy3
PVbWrdFsO6eV2ATnkLriPjIR2P0anLUx5A+prjgF9YHwKiv/F/FAXQ+oiT2tgFGa
Lmtq/FbncxoKG0RhBvY+kCDG1uG2+Pco1saFj6DRFg26HkyYhbFIxemw6lLe4tTu
+KgWbgnVo7p4mxolHY3iPQSh8bnatBQK/Hhi7UT5WXkWs2ho+mEck5xjilH8MH4M
DB0xyUrsPWL2TbEmBTiPk2iVM9cvTBC4I7FWTx8HnAdSvBtcZIdygi9AzuUDfkV/
0FKM330J0o2IGOPW2Y2JmZAWxoNmfAjyA9Jtf5qBqpIh+uf5x2y/LhfGL9BLr9SY
oiMlO50loQltssn1VCeASpvUBylgJRf+CmbEER7YaCnhtNdWkX4I+lznb2ewJ0B9
Sl4Be9DeaJB+81MzQ7BnLry8BrE82y/iIAv0jrR5oXtnKZ7JdLE7j0hLpIIklt0y
itOPqavZ62KU1Jr+dGqC05naB2Fjf4M1YUG1LDBXy70rZMoO9xmbRJTqekkTProG
jzSo5JPNdVW68zCqXQjUD4e+xlk3MacGIaxLnKAfvYQ8lTVOz/UPPae2XgHG/+vm
UDeR0c3R6wamY9Nre1jCUYqSKPq4uuCAcXBoIdvb1ddnjJh176QpJIvlx0zY0LWs
Peio6ygASddwziDHpGD1C4YdMJpyGoRatfb5lpzBakgaaft3no7EhMpyHwIYwPAg
Vut1eS28YoSIoh5VkH5Nr7SClxpakKre3DZVAwYzoJ4wVFW0ib2Sms1rJkUVggy+
PnBDN2CzsUSCLYHg5Yb24DwkUO8ulzPGhjkUywKqdQilWT1lMuDbI//3nqKXl5ce
OaqI45ILh+xVDuMkHGvkH6mjQEy4K0lWcQCjitAE7lAXn5O3Gs1eqw8eKZczBfEw
NY8YqqqOLr6RHTmOWjn/m6bJMTcXzR+0taigpzZGYZLFDiq/sXe7xcrQ8DGqiSFR
sOWloYjddDVUbYKwXBjFgAF3BRYUOw1ROK3nV6Z8CFsEQz/C6LVxSYqyGjbBweuP
BhG9H/AX45ZiEO3ospXSTyg1S7jylElOl2Fy1qktjZpfVlzBYhlMRBr31jnPgQbK
QGwNaIpiH6R1aciGRo+wLFa4G1vJHy0uCp7UnFJUatGQRv0Ezg6o5kKL4ZqrMBul
OHF5aG6Q03bh66o+iAeSZlbzFoy/XudEyiP8LsQvr0IyLDDQNu5E8VmfpKzYUGBl
b3coftaBnpwuxoNXJ6ZWvEHH4XqXMfQIizFdk/fP7BAS1DswCSaSGCUfY8TIg2Gu
DogHfkULZuhD7aQlT2fjj4nrqm3sMqSjrB8C3lGFnEAObl2k8Ee8E9qQWATuqjDM
ksG3mu3zt2f71MDQyFgpaKxNoWwS/5E0vBBe0Bhq70+zYxGkkuKdsMPuHtBiQcrN
MuGtZEWKJ++vfT3qckTOUVyNgNuitOLRvpc3x+2Tuk/Y4tKy5vBOd9J6G3vRPStq
hdCQViFmWHiUVuFyoX4ZU7KETRntV8KuS+41cZeRH9mQq3zFU8YViucAP/gFHzJf
4Lqvt9WcqG++GpNlv3DnwmsqI2n3Ml47XJBtSPrPV/BMWQjkVGJ6HjpPQvGFSe6u
qxNBNsOznRVCAaKhFWMBvw8if2OvtUhOQ98OrfbMz9K+JVxUa8oBC0Cjk9qrlA/g
mjFBxrYdriVRxXjoHJ43pJ+s09YrEogh5/A47MxyeAa72DHk6whjKkk9q2sYaIPX
Rmc9NhGHGB4EHwJuiCetBMxID1uGURAqg8ukIeIia3HutBLjGEvGqjpSF7EZV1h9
UU+wmJz/n/9MAAMV8egiOZRAryJ2o+50G5dTYmQ52MwYeCHMQje95SAeAqlI/QSE
JR6F7x6JJcXuR7VgF5y808AaPrzvvWqXZrKj3oZQNIaIvbO9boPj+UpvVdD3Xe8c
k0XOcayBl2IE/q12/pip9/SXizHX46JMvkePOVqUPcSVAuhAc0nQPnwfpvgGzmsi
TrUEspVPnbhU7Fx29sHuZUAQV4zEX3PjJoLwBYk4T/q9UPE4c5/8Ub4zuHdmTn38
uw1EzPv91WX71aZ3RzFmI6PdbBtrdpMJnFYyOUIxLmyjUiMfcgwaELOhepIJDfva
tHcxj0TDzvZcORxb9RYDxJWaI+XKYPkrGZ0YBE0itw0JDSfCSpzhUcO2ySHqIiLN
RXSa0NgCYfp5OjojgXW0I1qdq8GRim2g7nk2stBhR44tK7nZ7kMzww94/jm+LINy
+hl+JsoN5NUBWuz4Jp7aMRqnGpMUQShCIx0LUyd2C9wN0Vx6y34wEw/GqbEDOysZ
u90MUVtoj+f2WvbDg8ztVdMoU/bbMvcmOgZbfzozj7o5tCEw9U+9h2wm+N/BlLzq
ZKTsNEWdXOcxGLq0Y1UZXWTYoltIrn1lcB6O1ueb069MDCgyv46d2bGjL8EqGGCO
PQMljEHPpEQNSzkl9E2VQ56cVPwIMFosRbYhobupTl1g7gAMK870YXD0kKg+3ADs
isU5hghdNuQZKkBCF5om45N+hlrMUTgwZWGbTfUv/Uvd2j3YqlSmIFC8I0ObTZxI
YfdwTHXPWmqaM9iIKIJceWER3qZg571mmm4XiTDhU6i9pGAqvpNJrJmqcr8kv+bq
yyJMvtXz27Qq0Nqaqa5wDtS8LpaR7uWQn4gku2mSyfWDEu8Qtv8wnRY14VZN7WS3
4zPyv3K+FCMm/+ZklTM1Zslh8/6okzbC8E3M0zC6tAI4kspu7WCySoQZtla+vUPr
SvJ80RC/cNfrxSSrzhB43QIHqJDHhsCXLsDEeRX+oLBENshd239inqxsoMnXfvHM
zu5r3LkY7bDXLPDdZi2mWbEW1H5W9+IvrvT9PN8Q2aCHVXk0PeEEjwGCTy+J8pqP
ldh2ZZgwsI3PCa9pj3O+5BE4PJbJ4CMn5rNUfaSLZmIt2HVRAq7r/ci3wxDWInQ7
O2y1bPPugiPxnLyTMx0uhetoucy7YooQgnfSXj/z3cA/lFe045u3od+WDuEbs80+
Lww6V8m0kAyUG98WYI8pkD3p+HkGqYmwc2X7sIRDG2Ny4MqCYnOd+gpyZcExCuzZ
ScSHJtbXXugSyivITnDCY+PAs2PEU/M/9vF+YuJGGZdpcC+8ZjR8CjVj/wE9E60I
bD0wjN/gB1uPMzEOIPI0FInW3fDaHAAN1dw4BzQ8fiCJywsao/HeZoJPwLNuhetM
soofyt0ESsM9qyiCcTL8pfBBqJRg4QLfdBpxHInx/SorWegCquPVyvtp00OcSAXd
fm22OHNO8H0F4zctGUzjluW2VLIyXLpvM9NW5D2HT8QQUzLlYuFz4C69t3xhw3Hy
vzCAxm34vLJM2EzKZ/FQZPkFCD/PNfazRsi0GwVrhFPM1mdlprlqO4x/J6XeiQuK
rc5tBXEh+EhwRlQ87WQrppdq9lOlBiy+9ToyLO6R0sw85IIgsrnclkTzZ+KF5uj0
kLMeJ4228GiMNjmbl6JPq0TLTAdGwNDnrn3wEXjl7fKDyK5gRAmW5xeXiMpbDmoM
MaAZBnd/8grHM2udZJY/apaGeXgyQb6MXjh/TjEpBqU6w4Pozz2/YoQUL226yzkr
IMbIvBKglsXqIRpY6IcQ508ddaUTpUfr2Y7oXO4O9QaEXFDH1T9JGXEYp7CjxBJg
fyk1d4/J8hEKUJhGjXOHecyCmE0cUjJYCr6rMqCZC6GEzZoezWbmaOHl/lJMj0tp
R3dBQDQBm9sk8YFsDP431YWlBCkzl6rDJ9h4WqLZ1s2jaDduvMeiujBZb2YmIliD
UBHcvzlVP2hxy+pV10bFfQL00EyS9P1IaC05ZSQ7oJ/O1cbf03rB4+SHKsHD0Tgn
LrbvSwyYizIMBz3apnRPF2Q8ZrQ9KxF6O5w2xNiJKAGnsNlSmxwBMlbOdkPPzx0t
PdMWSeUJ7asEsww2ABMgSv9nZ+ryTwJZ3pcu69Ns6czg0+LuJhFwUn01R+2eEp9q
uacIumoGvlUo0fP5K/MXBlPco7S2qzaJ2YrfCYKbr2hThx+PpOmHGmqUKCWnbSH3
syr135P44hDzYKF8ZhQeyIGXeOecjNs9xVLK02/VQ4cuVoxIkJnHKL7+8V1pVyTt
8k2wDc6uZoq2I2367KZtczcyPJt3m5MISop905858i1MeKelWKkw2EWxhohjB8S6
+d2q6w88xSxGQcfsys8q5gRrla7Lgcx3BbY1sfi8MGMZ6z/8z6I2RePNi8qPYMxO
BEw3Mlgv+7h1nmPjR6JfkQt3vAcq7RB/NWr09da8OvDQdW+d7/i/Q/80ay22t7IL
Oie2WfodoSMWKjjmUnOaXJPAJYepgV/gP08nh0Yor8ispz3Bz244W1GyMvqiGaLp
LCfbAVCUei+KcOIZuUiWUqF9444wszSGKqHLOcubNX+gz+K27eAE8E5P5SMTUNhy
34Pu+fPFhB8vGyUU6aZWZNwVdv+eFnYyPwcW2IZNLgGkQg1D8O7mtYT4jhv3s6QP
Xeae91f6PH6GYTdF4SoiD8nELSdJhmNrVrcYfJzCg33Lu5H78gz2xmWAvpxT1RUD
TWDRR91n67mDgA/t1f1zJBNMkyo/LCgy4MVrI5xdbVylReMZLYBMlzVaYn7A2q1I
NyXFJtKHogcChVLB11SUPbnr1Lw07BkaH5oLBnPiAj4VaTVJWbAYHyedXP2c+IK7
vfVPFIc9jlV/OeqCdqQTUrArzPNXFunDQl/erNWHHib7ZNYV5gVt9kjRJkknl9HG
YPAOUzG1mEmxsxUEfp4duoiqI8yPKrXGjry70NxeOKU8lhUTnb62r3SRKMUdXlw3
5z7JX6lR56tD0X7jshvhm/mX1HhGKP0jV0fIObsjJ/ZufzR1q0YpkIGk+Ey2aI5o
YjCVVY67MPvvfqzj6lzQM4jIx5pxrbBH+2QYhd+/Q2JSVYv8TkduRFL7CjsF4Wrg
mZNP1NpOV7lz5FI0qSBRmtW0eipB1FSEqo64DMdOZNa8k+XxpD5BSee6F6YBWu6X
MFhHyfnkY9BV+yLg1liSusxI7OD40xMXM0PpippI74b57k5axcWxJvZTog8AV/V8
7mn6Iftbfp7Dtnr27cGik9QR4DOtXURtzuqhFUURGJFtJWSIVfT+tCy6dLff9gLi
RMp804Fg0DW35emTCkUj3dUuHN/L2EhNW6SMvVj4S0/lyTmbQuy1aFVqvG5LIjZ1
h5zPcGn5oBO8yYqp8WlsW/J8IdtHrH+SP4dvnbpxwQbIwLiKuhK+D0lpMs3CNkiz
FDJH9TsXhaO2ybEEwMYmlWHBsvIxw9a0tgmaLZQgJHTmClG4JrMK/tGdLietx1T/
FKNiThg6NjxXeKWLQUN2p147akhO8+FtmpL8PtFDD732T5y75r0PEPdX/InWfLaf
fJPO5QWSIplr7lt23Kc35YrhkpO2hcTbwwL6IA3daLKR7Rb6m0aCstaAvOgO0qkS
qcbNQkmUNF8I+TNH3H4sFZAd0h/XBl2G0RL7N9fGgSxkcxUovALl2FMd0jRO+8SW
A9+8b0p5lkVcjF9xEM+qtCoIByAYAwEpvCWdSUxVt4d+08EfJl3kVBGeGOD0PQWb
ntinRNlpjUS+wPGJvJnp9ZdxS/QhqbjGPmyK/XDyR190M+70adcAAlXX23spqwkC
biidYNlkh/BQaFcH9XTduDXzZjd3j6I0GkTeuxDD7eyv9/Fe8ZBIeElmL7Zs5MIX
vOmYKDKxpz1F+FGOYC2jeX/ZKbcgBQi86W64n5XBtbPp0CXiF3aNloB5oVCPhjDV
rcfc08La9HzK3byOMRI516g+r+7mBoG7fQ4/fUBsH7mRhW/7urTI1suirK1URQB9
X05bFn58ZrKiH5fo6P1mEq8VzHzgrNht+g8E7Jqn/CN/oOQTVEBtvK57UKg708O8
e7O+tjxrZcqRKE7//ow4hKxgI9L2vHYziJWikMDknhun94pDovPMncHC35wH6VPA
6VWbxE8NVrNb0ACyzBTt+ilAbGIqW+/s/+ckd0OCMsZbre7MOKX9O9VeQPjoTNzh
IAp1q3RsjZEZNWQ51oxRBrz9cIncGMNREKup/+W/84liqI2E5fXxcDngrcpLf1a7
8QtKgSihT5ZTuBHNZow/xD0djL9qB9HRY1Zfv22JTiC6E9sjB4T7ODfChtxdzmt5
fxTkRB9KXdM4q95MtW6QmVcOfq/VA9kaPSL+m5wf/9u1bKBdZVJ1rNW7cPv64Y6I
KGj763gxGx/s6U0IcBNGeF1uwNanOK3Yo3TgC9qduoROlMdtS0mzk573yj5qDwEB
oTIDoKzqvioqwULP9vAM1nHXlqArMXQ3USrlCgMmCgv1HjdEgEcdpGjxGPzLvK0X
lHE9wqWaP1LPXv9/7o3W8OSLPlrXYPNbQxKbnUM2gFBxHTzjBQgur1q5NRbTW0Bf
rmFf/i4pHDnNtzL5dl1ybVXBpAJazyFo8e+sb6FS16EFnGmX8jSBP+H9po79qZu+
U027iuwpXmrq0jzyUz4AadPFfVIe295YCLb0WudrpiP0qyu8jc+/xiIStuxiUoKP
XFVXdi2S+cGyqrbPVOhH9bzIRDLQuTKoWNPFZrTrwoHktgkqo4sfgfC3NBIlcjIw
yW6z6lJ8SPboDZPPEmj1RGSjycF0B3G6eteX9Fc5uUKLSpcLNCMCiO3LvB/7/Pqm
RYJNYb7sCVdnfyPR0y7NIAa5yz6EUWcuE+HAEcApzCy14SDqbFUFcRH4muM8G7Re
IsxZFD4A3GLPMsI+zj7gcZqmGRHfAXWSaqjXIzFh3o1hgwpqcxH3vXrOXvgNgLf5
CUSLg/oDByrrFV31LHpNhzeAzg2DPEyh8goCKKChCMR85COcwU2C91ZZVfoO36lQ
sdQQKBu7gipJaSBuU5bQJKj1xdc0yAPXQ/qQ44rP3lvDtgYKdZeg1jKUOXGloLyi
lca8yF2BH1l6m0R7KJ4MT/kx5SwtfI7SmUMvAIZlMJEP7BPaWkbhBusscGJo37fd
aRh2rrPD9FqWIavhUiILM6oIQJUlS4LTz+pazmFTSHwBsDBURQaDYNjG3XpVrkSG
lFVBl8YD5b9E8iXMnJduXOT37OY1rUWLUOqCnQUwTku5R83M5gAx7Xw5ZgQvBMW3
V7UCeSfpOen8ll/zEo3SDmI9vR6YARcEz8RTImZsBzyg8PtQX5Cb/5RzGVlVZDvU
OU9d5GnFTUWoQNVNXU2/1ed3hjlCXPJeAMFOzPeSIxRKvE24/NPk0X8VF1g4wM7r
SPGSnnyUsldBlEcpRBGyProjBkw23s+d2dBoq2I2gGlD+Rjyjz6mzFTs88t6pqSF
fg5ah9oC1qcvS1F8/hXs04XN7513KySRuzqLGn9uG7zXdn5TSqRDFkFE3dht9Bog
cvuoI+xQM/90s0BIxKz7rdW9lACE1tmYnXVrZCx9XZSKGk5EvUzEY1jFDuy28SOb
eyviNRGC1rHLVia5XcNl8SjVFEaaj6AM/e0kCwKlKI/Z7lkVuT+HlN2bmKaTQaxh
TWtZzcD+1ciBW64KpWl/bHOqRvp7zdQ4Wv5cUnUOl3fpxuXDHBORLSQ9M94IgXOe
1j/pJdCW1F2gpfjNZ+SQuVJgnSrMPwUcMBYfq6+iFnk10ZpVtdeusTAUruIucwQu
bSSV8Xqh26DvD0wqXK3j36t6EKDFyxsqzzspk0jWZUf8Wq9EGgeFcl7bgCO5EUYV
CxRca+u81+cmwJGJ/2V2AdTaAeRmw28pXh+Q26TLGrZDeUVZec7aEHFfoRYzEY/y
4Eq6u9zV1uy3hDngNvJjF7Q4KhrQNd0zVbBr45RMnbrTWRJpiXwohVyUFtMxLRxQ
qnCCe8aLYhHHBQCL3fReCLwlON60EdmXXLjVvEML7laFpvfHPwuaoVHaVUpug5Vo
/z7DOvRbSMNJjJuNnk188WSkYJOUumyBOQkcTGByfUsUfZH1XT0HsyLffWvnRxwq
rk/jSM0aMBXxTn5I8vJFimmsxW2cuyJsQfeKTFIgLgzHhzKsxIYawgf/71RQjAFO
nLaEPi3v4fqQYv1e7gnqDKrgTVeqIuiJDrhdvh3pyEnC8j2+6S/jW6H8TrW9dYqt
UeYfTMlVHtWmdWmqDs9aGDrHbYlxplEUpF7rkWl1kamDF9KxZE6Z84n2bRZpMsGj
gne1WojUqnMzXFjniOpLX0uueQ28end56U6jwV3RcxUmAEyLaaWtiqcOAPlKPL4I
ErWPyrF/hkHHugs0Tm3s+TpXf+6TTi17KbQC2I+xTdkjKCKxUF8DGvex1RW9SZJu
+vdDnkSl/KUtTWqgjMPlb80MthzLIknHuuAhjnL2dLZ0BsrjfCILqIewLOkFvtrE
V5qv04BF67a30qwTAkotqQ2JS0IVy42eJyMgAQ+qPl+oGawXe27OYnUEvko7c5ie
UqSV6ayKTWTiflvbRiaQliWUaV+yYNLoDhzqOWUHry5dgDv9DMxTLNAVAVqDPrzF
O9DyXuCGgXeKWakQHiFLifj3FEXjOnxlRjbhuLjbyzDo3VB0KRto6fs3p1qwGKyY
1U1nN4ostY4VE0yuiDUuwBwftea3GSIGGpHBpo4KJ6hJQeIkdvCe3pwFYqwWz24f
91dkYxaRmeYZ3b4S+zB3P1EdWe3wNqmd4/wdAilKVb2+QsKg2ZcLw8G0sPkTtwDM
nQx6CffLziOmjHER1vcvZX8AMACQwx0uqIh7vLbKEubsXWOYHH+CDKG3t0YzryBL
XytsLfxA1FVdGq6PMrM/bcyiTz6bXG9SQ8V/PHFJTwgp+9xrvEycWmbBcZtGXGgl
itZ9BEkxotqb8wPvnpBUGyPYO2aYTvlYJI2zeEpSgVnfx1FITF9t5phkCZWBvsCp
qI/jKo3h3aa+fgm2IrQ8Zx5pzX/sZLtORCUSfDlrzO/TYrGlXwSGK1xnJRbECcUQ
yBujPZutu7JYdJpnwo2c1raW/rRuQaknUigxpoPzSg8z5elkZG3CYW9u9MKAS4zK
hnzr58XAoh9KxDxkPmW/eYLzBUgc/YkMfT8tvLpykzCJ1UrOLbQBOqefCx++h2uq
CfTHmx6s5pouEP7aFAX+srBwwxXD3dMJ3LLTpuN3JZ9xKqlGTjPlsi/ubteoo2a6
G4fbIOB5+1MmGVnFiaubJxK+18M8GSXMizWZo4Y1FJBiqNa2R8KuLcGT0GHUooti
7+pNTFMpHAbtONp11RMsfj3L2yQID5U0UsfTBMg5kUvySjL+4c/CVoKRTIaxziyl
k/2lm5pSTgDnAxlOKZMaIK1i00JjOwwFw1hiiLL3/aS6lkSLVc0gulyhznijmo4x
9w3VMgiwq5dwt5NN+6HeMgf8U1K0eQuRkgh1flli+XcKYrT9WXwL+ZfTcUlQmuZ9
A1x3hUKRN7IdI8pxvZFrquXqrjLPlevD1OJ/La459VNBs3WwW7qhPiVkP5LBLz1u
udsBJF2UMXy7XVDVBrpnBiRLMHOHyX9TFK5uxCdSVbizhC4mqf/R52xjg7p3gNdB
4a96W5SqBXg9yUzO4LGZ7aDluK/xseRvJ9dQrOw3SpKbHSQXz67Rkk9nZc++DuRv
PwKUzwyhKpm3dFB1hIYkfhMDllnOCdp1e0F0p6X7+3e7+BDkBqnD0abRQ4KiFpwV
KF+yRuaIfg8/KwtX89DWDQchvQuHKsD9mkbCq6RZMUeGcslCCPbayCWj6c4MFMKE
nzkZdSAnuIUj5OHpaxtK9+SGRdzMrb4mc26NTdkQOwNZwgki0RWvhGmzYaI3k4Ca
X/6fE3oyYNKQVVfPMzB0bqmSlKNHtzHBfHtWeoA7kjO1z4vd5UruyWOees3XcdGU
T5FNbl4XZzINjrKwIMmITA8oNZbGfolSKmZetP2d99mnuBBLw9n+R9J5ytdePHwe
vkk6D1eNcewz2Q2g9hEvb/reDEWlR3qnzZwYZM5RPI1x4rlU9g2BEWzYmi5tvbPc
2TxrLRAZuXRyDP84IKeHouYpWx90SMFk1gyviF9EG0sO9bXg1JevBlcrtNK4RK1Y
pIkhd+aJsnDgveQvKDNNd7FQJA8UDqlE9PGtuwQ4UaL6Ijx4VpFLBEUpKUy0NdxR
PGNotLupgbXyTIpAgCrlDoJhgqtPdW8hEqZwuG/q8GuGUbKeTNa3aC+Zx4vGPQnI
7O4C7ps4L1qFdUu6A4nUOtQb7uc7oGlzD179nqY90QterNcKg+xue+BFr8LfpajX
ZWE1nnRVN0WWOyhdqZowH50cKgsDeJ8ba5Bt/XK7U5cWNqn8gDNlrv1Plh1n9EFK
d2dT9bZvLiIM+i3a5pM0RWl7QXA5zDQc2orta5NmIsrwiVvZMvWQT8KiRcotRRZH
DxncpgWt+q9xa26DFOE2sfnhHSNGJboKGmqCc0OBW/G4Xp13lZjVJWbUVnDoprZK
vsLLCNE7MLqLdWpb7CL8/TV/7RKBNhA4crjwiGGD4LuzSGyVx7nq6vRiEMSmpgmh
WsRouK1Htxoe6xNYEOC8YSsQFh0vHWq741rJkpnkpLMuK3MMBfJHjTY3IOqACVCZ
RL4V3tPWmj/AXrRa7uaI+b6df4ivIu3yBZ72NF5QI32vf2XHTs/QC4xB2xKPdTyc
gPpW3riioPWm838WwgEhOLbyk5COMcp455Svglzv59uJ5lQ3l2NX76CP5yXsYEnn
qm68G1bQAyK3os4j+VH20OeCynplu0aew4toP52PA1Q2wmjvMbF6+vOmWcxGYwnq
+0G1va+OvcsGsNzezfoyhx4iSkvAl9PG8A3Q8Syt2EIIRlZfDj/DsXcAVWQxwuWj
F/CCtv4dPJow9MTEJDRbzplDz/Obx47jNvruC5xj4D3eoAv5DOJRkuLl2TueP0uh
dIuC7Zz1kb5WRiGZTnHpmgYMvQhZQwKYbsubnnY3p6zeT+fv5IqJl8MkCCq2Hq/1
NRj5QJtlYw60zVk+UnRBpqrHZI/up7Jy05rpJRxCFcIkYr3aQkZrWf4Ew0Uz0R3d
2TI4wTz5lG+YfJUZKKlRP5w8/XpRNFVmECA6nCgdtYaoT3QEdphoZKVJQCyVrZcH
0qvjqSHR1sfehTKyiOauzX05f0Ia+Da/KgAl3BFUj8NG/pq1Ucv8iCaIpIMI/aXO
0mZ8ERpu+mjAVS8G9WNcD0JyEO9Gej1jd4GYZlk0dzykD2qPaU5vH5r0C9pt9nfx
9r605lZH/tbNRHnrseJuoVYIIlytlkzoIxS778lJOjErFZBQ25sF9g4QZhZ+232U
zgo19bt7EYStCONow7DgfIwsbQhQpL/TRK2kbT7PYXv0qbfz6Zi+bxMHY6hG9Sj9
kF3f94Ve7vyssYfFIYm1g+WkmWwwzHGkkpVoNjIzh9yCVtgroUYVfOga96PhTrTS
qbkg+zUNfhg02lGGdFPNDxMySgin/iXk87CdFZ5Fu19mHZb8IychgW1xl8uC2B4b
/RIXHz3sZOWbyLQ6y4W1Q6BMoEYHsJmfyZI4DCJ5b2Yg7mHa5A3umlKLtLJ3tKna
GtCVaXYkr+xFWp1trr88EYhVlCkLbpHi2c0JPRHcbM59CREdlam/dc7qb6JWeIec
TzRxGpIREPc982eKNrJmdFCGDvAUUXhvx/ShG/eFcAMWWZTfQEyJH1cwj9ObmbdF
0tY9vWT2b/ujCxPMQNfi7ge+LFFcsFN6nGUKFl8XVf6gAJ2KQUNGIQMIPJxOsVRm
weHl+sPSGMJjFpuCJzDdLnDJNcueDdhEeC1jbkh6Iz6vMVizN5XpDem7hjLRrW16
czLcb3KCpefoNt0ADbSfQd3orHC1zKLmFZq3VMMcHBwuhDYMKTdjbmazi1lIkFaM
Qro6IngK8xadhYwwb1JvfsMCmmWYZnxAte9kbsDmjWDXw9hNPUgseQZiWwETteGC
s9m+wNwiL+HWV+yLQ2z/+6I9/AoTmmeIjDuCeU9akhWueWv65TtXC2Ih9VBjPrpI
SVuX2EO24oUbwNEaack2xqChpA/maAEjJfeJbZH+WbfgPC8GQbRwBJJyHN3IQWmQ
hgAYrPWbKieoT1lac0iapGWRDU/H5QTHUhngL/pZ0UQhy6NOU3Nb7J1Rou9sjqar
g4F/x7767Dx3e8+/2/Ljk6rQd4k7ReX3RHw+l3bsuh1lWUA4+1siuJMcDGVN+ttn
/KP9FMOfegGoyd/X9EUXVOn2BIF/07XShv+I5475wxSaPMM3dtxzW5ihzh+7y/9X
2hHRcCyUPGqNZFYZS82rzkgsfZSIjsjiLY8aeMD3A6iWSgtQd06IfB6BcroMK0RB
hbe+GAKYiRS5xxhAcJCi4/UKfgK4rOQA4f79QkWLYtlMly+NGtzRcWOKOWamiiCy
ci1B3FobzPMQm0sExvjkzFf0t0ofPODYLXLOCn4/YqxGhbEkfUfwvHfaG9ELpb8z
qOVZj2xwVsm0IipxynMNfPU98NyLgmTZyt96XWKa2jx40WxSYiBKm/+c/aOj/wr7
4sbpQjl2E2NJh/rOIPFeaivTfmqr7xnJG6N4na0hcXsCdguZk8ZNX4b35iSmrS+U
biAvL/zKqH1rb9HEIdDEGJTw8ae0exhbPPGo4Vp2BkYvMZkF7cKPYkefcON/rDou
JXXxbVQ7AmkcKp7rZV3ykohHqgivXmwaULl1iHn4bkUq2IG84GUYukeD7WPJQQMj
nNZllV/BVIozSCBrw2ywbuUeZFAprhDYOy32VPcKSmanUD2mPhRVNEvXqJHWlpCe
8WTD+3bq06FeIWsHVylt1m4IzYsxsIxyr1WYA0Nm5104d1TRwSNva6MKxLdPreK5
SKVeG+xGt6UQ2Aq+DfAGWTSotKPrFbb/6ERqPp1ja9TRx4Khp2r/6Yy84QJaa40K
E9zwE8AS85xpiVcB2Xj2iBiJxH5MYIGjHQKFXBm08ZG+OyjPRLuSkVOxSsAs9GzH
9dSuCXSQCwGP3to54iosuK4VTzF0bvw3o9nr6bWZ9nV4M2jhGkdfeiC/o8SyUpxJ
cnlRC2zNmtmPshvEEcoZwMv7IBNnNuV95BErn93SI7ZwONCq4CxMAdJ7FpSu3tdI
AzNY3s5LiOMb/IZtRaMQwwcCGMGE2OVkcvTjfJJkcUOOENsKTuIFOE8pn6K1yC6P
k+XbLfpBsk+o97xrlWj56uk7chBLIN2GuJfiLp0RRoet44xYYa7XlUDSNlisakaY
3NrcQgmACpCLRUkavd7JQsRO9zaFCWuXx1CdbwLJ7ZqhdPjkMaGgZ8HFt+OQFiu6
KJCIC56On8Op6p+bLcDqk+qAH3ggVkSV0fMutlgSghc+HpwCCMbrcm6RmE+CYuCq
PXVjpDSUJ5Nu1Ru14QY5sZRXonOaalhhGY8jsn3qtcEui9mXxdm7XpWF0cxmLIF3
TBENEYDNrlQdDd2mCHNczDca3PIwiISkyUmMx9aVB1TtMWzg/l14rGUtTjnYMBAk
vVp0G04KC2xowZb382kRb28AhyDLe6DGx7nfjEMaLTxESlT2/Z6OmRmT4eq+5/AB
JoU6YmW9G/duLicDNg8mtj7PHfWFzN9wnq2dhlAxLD/58e1jj3VmAoWDiXxcwzOx
CtxcBg85NND1Bo9iEF6GsCVxWwH37dbYO3wnDvGiWfrbj0Y5LyMx7bl8b2OSknUx
RWxX/U0X3krgrNwX5DBr4Y4l/G/TzTadYXTmymMQ5WMUam0PXoiyBPj/jM9WTIj/
6rZMjM74NvvO06JsINTXYNdqVTJ1OoAm+/J4UAPnmIv07b5eGRAD88HU6NgteH3h
uRpGKots3vSEZ3clvkbmBP1dCJr3Gwno2GOP/DVgORSjRG1n0ZnjUjrrFKcwin7j
eqSzLLNE09H2Ia5rQpT8RPERG3fRBxYt1OMoaUDCXu8lxx5LiHvJTCoEkMysONX8
xLwXFRVwLBWN5o4g9C/9qLzb7hwNeP1DSjbRczBsoxMULrZiyZYv5zDvIbD2XjJw
RWJUpiMDCLBUmxdreuPv2kiGjc11V1tJhdjxYz4aKjJpY+6Chk7T6PUhcmUd+vm6
C61+Kb5/J2cKE83u7pIDyFyaTZtaTYhuWZonnG5QWtaQTTJjZGolia0doRJ7zYpL
c6SC4PXsP2O/orwAbEIFSC5vWpi/3UxlMa+ysDpZnyLV0igLJUc+SUUZtZr/luTB
gNaMo5Js+hes7n//2+l8hqp2LZFjFE1GW4L+8Jh60/wPZvbc3O4Pmle2eQNsayE5
iS0Cq9vdvlnrmoYrbP7O5ErqP3g/KgxCJcw5NrrjdUthsXnwPXBGtQqb7qS7oUK0
ZEZ9L4YBvOj8gxxqBD8P+InfugyQ9eSU8VwPiQ6fVXGV/xKHKrx9SiDD9RDQl7Ip
v5w7Z3o5tQD+BO0TdYVS2L26LiBMlrQsdXYdHzNTabsgPjHUEkJ2oVVHVQyZd3rC
aweKMoaQfAIlYjrNKIMltfJYRua34wx3HlOKZozWlRADRGVDFXghjhbQ6OxELids
kcGydvVlwitc8ki9Wi6BUce4cWEuN+uUaB+UO5Qtzs4esFaMXaQ4un7mISxscmGt
Mqa6xpfQFT+iowSSPnulrHYJlelNsvfQmyBsCY03fSSPvYgAi0XLrvwJEdE5dyhH
8Ziq2gUN7UMttoXD78wHccsBJfuAtU1HmZJKECkL6wqiQgFP94lOq/zoQsqTQL17
msuBXyZ+MjK2lvlx0cV9Fqn0Levuu+JjSvc4IqA10g4FG8TY2U/taYlw84B3tqpG
Pkr4plR3E75jTCtGCBo3uwTs3rs4lysfDId566Pef39JVeGXWNJKeF7+q3qeOCwQ
5XTQOZ/njDi7Dtpcp1WntKLHqJwitZZ3uKtfoS0xvQAGZ4XUP0iCad1ouDPegsv4
TXADuBv0Zw9I5KGsXNFGxOoD399cj0W4vrQyCJ33FOFlWopUiM8kUyQqEICIpyt3
N0UWHZcuRfvSmt7pnZNP1aoWtwRSRTTX/oD2eWIyYBKy/i4JVJYTftW6qtqCNEG6
JNMfZm0Ski/kYclFIg2b/Ipe8D+I2GUtur28rBe92/VQbN1qOXokNtRMsTIKvmti
5KRRlVJYByHhe8LpawrwtSlSAY90WT8UwSZZmsAPzNqbfkSwAQsXRlD/FzGu/NnQ
aaNxz93CbXgYlkROxdN3Dp5DkqJAEKH9lnM6S9f37wWtXvlXH2TdD7JMFWodEuv+
/ZMIzwi2DtIIO56ACibisKj7/NyFNA6Qfqa1/1wA/MSpS05VCazuuVyY2yZL0wLi
FET0ioEojwfygBcwbJ1VaY6iFacVX1TXnCJCiqTgPiPWB94+bWKMqUeTo6PbgwjP
ieE1WR62Ws03TLyPsVdJBArE3Hr6TdWFA4o1WXc+Nm9NBKfDTeHQ4efLs8H3O9n5
cMwOGEpdGcGcYAojpKLLK8oyMY+WlX2JZVa9BqBTI2UehYk30InTao1gj7lTs4bB
VTXwZLbQL2WN1ILuK8UKizx1/HaE2U5T7tvNqh9+B4XNvHSi3h5+M+ippgljUCA3
fyAv+oDEO6XBD9y6rb4dVKwJbhpCmvN1BekCtbmBNQVP0MYK6S1E6PUoCCbKY9J0
pjqEiq941eGdCpD1iAnNbIC+xRgZZ9cnqD47T1aHGwRL04dpBjoNQSKysCHsNQ4V
nm1fpHn27O7Xau+Q2woexRbC9adHqBWGCGKAzdWS0uePMG3RICnoZED8t4+eJvXd
K0ytR36mFw5XE3a/mOGCXU1onZzx91JEvtFYH0u7wmO75zjPkU0yFt66lYmIYol0
BIUuDvOqwY38UWzZCic8PLJFtwKYmJZdES9G6HKeMuDYT8jzuOj8P30gJaz/N7HY
HRc+Iq3+GCHOpPyGnrpj0t36WZN6olorP5kIlBGCZFAg9OUNhPvs7LHG2iBJKb6O
0xJdYVE/xjxP11jcBExNlQHW8mQKab5uYRK77G3cVfNpzUhvoevEZZ2kTMQvgv2o
5N/DWZAmov8N1/U1vA/MouKwRaEnOUOUURQTAMZ3mcQLF0+eXcEP3TKhtSh3tc3n
hBmzobuSiEvEJseJQuJL9t4XWHhRJgM87iyHR1eFGtGQJHIG6aC+tfaRhOa0j1Wi
fHTKMm2eAAF1b+F2+kWtuEot+8h/K+357OMD3u1iFzM3sVx8E/LUx/eQLE0XsMKS
45xaX9VyJwQzNgnBEkrycFl08/ooPNmwsfdKdWnAL8N+Ap9pr+3zq/6gamqxqoUv
F3ERSpSqCtcAPkGoLgLTL6PUAwHzcjVAV1fc5eoIETS4re9a1mmqOf8R9WhRGu/G
TUDBBxEbXZX8AVEKsnLzBPao8JRjxzhyXIv8DTvzaQM0hfGW60nE1Up4Ezhx33qN
PyPl9kDQwsj+0x8jICs64bk4b0l06+M28knhzP2R28nyHYIzyqAwcVEqaFgAMr4w
U8ZKHOwG2Hk6e3hEPtct1ox3IL8mdLvnbt/jl+a6U7ClvzPzwFkJDeEF80dBd99Z
7THLGbCXxP9ariplAUONLH7yG40GwEHT1dtvi4Qsxp3YQS+Jab4WtfqAWlLlxW4F
jqMYH89TRSCSC0gzH6+AfbpeFPcDqrJXtl+FVY6WOHofvs1VWIkbQmxfoxMXpVP0
j5erofQTeIuFmIZs7m15BA32M5hfyIi0NswZkULi5Zcw5bvF93gFsaZAFNFmLp04
gzLowZ8SQYdIFssAdxOFTl2TQzX63i5qYkIds9fttfomj6g2lYlUK93iP64fPoBv
lIBjDjDKJkeCzRkUke6bypHtYKVTDwXYAonJcUzDw6w+EyCuBvwe8rsmWgoJMkAA
4xnnXBxWDGNkr+AeUZ0aZdrechVG3unDzVEfbNKyjkfliwKL2ANM3NtTvvIp70Yk
nrReqLu4B85q9piq5807rXOJIQfyBzWAHYgBm8qDODvWGVweAUG3VrUKEIbUk+UE
DI4lt4L6q3XfjnRUskfxesnvwgB8atbHSUxMieY/TLj3E3LIaUzlbilSa5t6BF+3
Cyw4MNQQzDqhZ5rFRMhbDex/+T5DRcYBwvS6bcCGfCfWN3UyXAgqaceRtYdZx9dl
+nGAGiNCSnm8EOyUH4ItK+3X/n9uO04uATmwOP4TsP/x7isTYxiQuT2RLY9Fw0wQ
fr05R0RUW/OEFh0iDIvk1Zk1SMWl8h95UdYNFw8rkuDvkznpRUy2LJsu3buY5Y6k
Lct0paycRuXEPmg/YYAcvEqo3cvFXgz4NNH1ibOuHfs1V3I1I2KNya5iyYWAL1Ex
VIVptqmiCDZm6d+4J65FyiRd5eEm4KIes/gkqoHodCTQygISfp4iiSyJIvSLvOBn
4PXK2LIA7dc8MjvebYA8FNJBAPvZFJArNc34ErpjJcHxxXMJuES1LIZ0a0cNs0Ue
uvwgl+SbnIIpBLpaqsVYEWXPqNIj26oh6y5A8C8xZKHlNtVesBMeQpjLNWXPsEWW
E3gNHRSOBAPb1l7+pjXaHoPyKCMn/s4GC604M992YigrUOLc/+AHVPTxz4OqC6KE
NPeL3LEvSTnJ6z9h/6yZNPlimP1Z8GvrH6tQVXUV9POppAMjw9/k3g2t8wjMqupI
m6pSmdK1aq/KJSTMUIQswCirCLMzzmo1h0Fv1OdM7K6pj5rP3B4JdqBT7TMmEMtE
XBVQ9SarK/RWtHzHx5BNlXcw9RsCmj6ZInNghiTvb3kooilK124ix3o2DaFzZviF
oJoTjfAevwWWhbvV6+tRoyqNVluKZ7dyB11CZ57fsV1vkgyIo4T6SfhoR7v/hMWC
HpC6qKo9yySM6JpUHBKG2MxQrbW3U38Wz+7ChXtsjxkJr/rpkJ5Sj7bMjIsfMWlE
75tiVmDenGV3MHtE6flbb9FGxEnfpNK1MgGXSAGudclomK2UTTEJlEqvBH+EJp2m
1uFY8qkjiKg6vLLAHu0DvHOS27RFUgEDype99GRCnLT8whKygagS1sYK/sjbieur
3WQf6VOWCbE4N7k/tGgdxML9o//Ni7r5ISJxeCxRW8M1hhkFfwpIFsdR8SqgMO8P
oCU7xz44EpbH7qbf/zmQk1KHiH3y4qIxi/RXgxeVcTerPKvyiW8kkBoVkaA6KIe1
CeTxeMxAVY51a5KnX/JJ0UWALMnqQO+igG8jLVr2cU5pJGSq/+BFeZgBw7oQcPpj
c9MVBwGXYGccoF49CjGWTduRKBKDjy4GUspRGh/wZwWgy/HLPQrwzGIC1nxBWDk1
YOgHJSD/87/cNUvDwIQfc58yRhkq8aX1rqHpsWrSJKHNHC8v4gz2cTLD4bw8V0zu
BzrwxYkXwcf2ZNtzyiYfEsdSw67EOOTwPlzchwdmvle/YJ2uOjxrUC7YiqAVPMFa
LP+Y6RDqUbQ0KPaA5n0yRRXARs1oO/NJTm+iv/dCXQv1kXRHzdxH3eYZzKW975nP
HjdU8sKKHwsVz8mojlFVZDaAy90h7e2Iyyh1Xz8nadAzQenuqo7mg1fnNcC+UL9O
17TM1jZH5+CVjBlQ2YFdmTiqYr6wjWfmEabs7pj3qMQM0WNLN9bbdq5v3+5RKLAe
Xc6IvEg8IYxDWMtSqPvCAM4k3agScQB8KiV+//RWOawshdJUpa/IFj248RuXLdfr
7WYesrY6PvGb/JwSOetc3A9j0dA26AzhubXHheJnHmLv4SRIyjj+AuTPNCjIEYWI
rMrRZuxAwvJ+QDehT48RniVK7zaxse62T479alvfgiy0DyPHT5SuBfGzy6PM1HeW
2eh8CeNrGMXxMhIs5bZFzN3kjUu8jL9fWe5FP2Og3MAncxKTal9T9T8xPKjYZW8Y
VC4N2sS7nqaBvC9MjIsLZYkEsolxqYLBqEAoY3gPBYRR4usRPUBcqaL7A8s/LE91
vlm2fX50J602VJAqxluG3dz8M5rNzzdOlrd0WKXT6eQdGbDo6YeSts3IqxaXKQWP
TWa2dUnyrJetNX//l0SUhki0tqs4HvtjBy9xs1yCE41x8qZcb69xiy2eVuqyVq72
tmZJTBRnuLN2tZwY898i/3BuQQ/5rk0CFhqrel0ADnlZGGDH3glNFdVdXqYxHeN2
fK4yN2lfWbUWlzRjsvhmLFyrKDqJzeYpl7crIV85q9KUGBcoYop2cZQoeSpIENmb
PozZ9oqww03IOuwbszctzU11flk03EVfPBsnOCz4Hmql7gLlk2XBq+aFVAh4sttp
qvhy0TeBtRVpJsAOeVPMjcub17IFKMqMFBOTsxbb1LAQqSCKdtVozEt4gt7Rqaka
uG1BT2gJsfDIAjFs6uhh91xaczRwRVAhuxQU0t0+v5/6DiNDKSiNaWRM5BTbbNg1
3tkNSW8us35nEdobgmLVQNf1wtsFPBXbmOgc9vjx5PH8eIFmkO53T1JsFLMQlKNU
ZTmReU+8gKzTEwKeTrBzWVUYBvvo+PKZteL7wzkcx4euNLL7A1vhMELuMF090tUn
I3szTHYaRNaBknqWTJ4yj+qjxqHA8wpSjSlG/GESzJ++kLm2Lfckl2k7UH+8vRTQ
R6FPpcPSg+qW2LJSYvigcqUasn8U2UMNOg95xewxbb52PRda1TOVeOcx0fp0v1Qn
8YPpDzqbQ+4jKS1TAg37JKEaEKH6N9bQY2bsq8JX42EHCZ6+MA+F7MVUlM/dml0I
FIFDuLf0WwuQ2k0aA/vSNaj1lZIGmW5VFU6gsjipn/o0Eb2O6WrMaLCr9hksgESa
ymrlW8wVxV9OVaCixkHz0Xcxe0ZFoyQizVlImXPmwEt5fvpdhrAhOI3+bKJwc0KC
qBGT0uSZsXVn+LsJuMy2p+Ju50I11vHD8e2BrMudR1TFkpV84gxPT5V/6mf2lvfS
juiaOQoHQ7CS7chb5fqUbcjrVsGoyPR47Dc3P672ETYgiZprKa5EXt5m3RGo5BF0
1VAZ19Iod6DKo/Xzq9KHKWPEkznWySFNzLbTSIMhEbHCfrPWtjJbq/IVUiB5t8C9
tShZ35hA/QBlAz2q6lw+UvXBRKKq+Lp7+GX5zTSc86bEi8LDU/DseZFVZ2TeP1nE
DoBPROljJ6CscHT63i9Ucl0inGRxM2OezxTxcK0OpsikfLvBmie5d5mZTu0//5p0
xpjxBhDn8PutezIuxceEoAh6WNHtD69ADzG435Sqw74bfzsVXvviDoVJQCM8K/Tv
SPPqe2WQGKaMP1brxq/GCrbY+H+1/r7Jzpz9e/y7qSeC1MQMvizoXKmNBmYkaBMx
j/7QK+6j2u7hgCAyh5TIp6nuFIpeR0QD4OYN1J+IOA/Jkvfpu/nk95WW9RaOKu8c
ryR7g7HYGfRhcapEh9bXDqpsEZhDilYX738SJA+A7EO15KVml/b6tdYo3rHMLW0l
Lcf8Ypt7fL7w37G3vmqqyh0ZrIGF500JKW6VFLuD9sCd9x6L2NjpnLfl5Ab7gzMW
6/mOUKfifjvGWYWEaL//LYDppgBzQGaSBZy6CNrGn+ebERtce/dB/W5tGKE6CN2F
uS3NznENi2b1Zwio1C48D2tFPaTDNwsQc4rAjJsGCjwXQATiE3MxJhwvUpo7vIcF
5IAIdGyKYw9D6CgU/L1YUOsQZKpjflzT96h4eRu1h9XR3bwB64UiiowFIOmmF7Kj
g/eLmjuYMl4splNT/Y6sQiy/lAk/jgW5vQ8Y3bgiZKTnQlRLxmgglI5IK/g7mSfP
z7ImNt/B3YjM1XLCItDdjGA5MBjTzhnp0aaah0jXa+3b9slkQRhJtshbEvxWJgJ8
PpxgJKmbu8gwR8HIkbqWXLMPaCxDHl9o+kqcg4wEMfqIAcHhpPY/Xoi2k4FKVKSN
/ruMnh42jA5EzKiZTPi7KHD8mAS8f2H2+VuEDjHHE7euiPBRaby7RAiB8u4Hwtnu
DWP6tHNG2EBxZH5zHODCX40oeW5eGwMfykGVirQ/Imixef704Qk6HJq1lSZF1+nv
XGz7M0LHrOS6ZUVYr7LYNfcNW1YfivKv43AoyC2UR1hrTJNC3hHeYZHVTwhVPgvB
hj6+3EEx06R5xtMrAWOI2jY75iiLAJFWGPHJoKEoJhznBw9LfPXN73OXa3h8BEz8
IcdkfapSMp8o4iNyQJYfTOZRS+xqBkHMiy6khV4oz2pn1Psa6a6+1cT+d+mCEvtd
dfv+1KOXPdquEylvEz9CImi0E9NyQmFmyZDcTJLAriF2ULiB+7hHXHM+CjYVibJp
ETGxCY7CnUsJdsDaeQj5Ur6BWs9a+MhKYfErKapWAcMIwhkH4+ILABGKurTHMvMp
JlnGu1XRd2Wmq87tLRZy/xo9oPfBu+rkiaQGtmjEBoXDuLefdzGZHXSc8Lzi/904
s+DjGR4lQ6wPxk8hEDLQCVb4wrZ+G+QtROE43qWN+UDEIurcz9Ymk0CR+mqnuRdh
7o28hXJv4QRNQB2HPNby/HpK4w/4p/vncFViSJLISlCumpbNkY2EqDnos0wYi+ER
0iIW1YgaKDArlfRl15c9f7i7MLDIsy47A9bWzW34B4qdQJTpINYNVtNKiTbva+yL
DmnUAqIdkCDsbr+egTLI75jM12PY+LZL7ZABgo91ssk6IcOjbCtKi5lYtssokP3y
3N5Qbfi2Ht/AaIruvcLNBVzVQTyNuYyEKAduISNc4GbnissCyEHy0h0RXeyJkNGx
qKxwkb2117vCmmC+5MBAqiDVdVFj539dByBdESD8YnTnawXJlsH1OdOAn6EYryPU
MKNZbmRg3C2VLgTNZbKDEl617Arw1XN+uroHBFzbW4GGDndwYsVUwITF8wCr8zDw
JmESTIQ7TDbLTc9nI6rlGbTHJOgX+bLugRoVvNTCnIeX22/KUK+PHq1NqCmLSw2Y
9kHjCDDGHzaGR9DTuEkqLudYx1kMSPp/qdhYFK9RgliGIRSzB5IU+YbpvjPPmpO3
CsF3Wb+TkFhW5BY6SnzQMIp+fOnZuja4ag4Gv8tLmeEMBxNzR83dAhDxnTOlQaqR
Pf5nNpvZRUeUHJqs93tCyNC0rKScf2eFsG87EQbz8szR+bPLa9rHzaYcL7qcQ7GZ
KUeYyCsJpFXATiRryUGVCfy+LkimQKWbWCjpRjCib315TRw8nrHE4bxObWw/zqaD
RhTb9wZgJpc6SEbdA7vZEPJDSM9BGyZbqjFGwOoUrbBguhd7OFnwDJL9c4F8sl/I
vLHWFi/N39k8zYQ+nKRqm+iXG0NqBXuKepD+nlcIn/HDfAHflF4Nyqu/pIXFHPCX
tpDqYL51dPn2cC6YTfvgmk8QY5Z1bI2p04NKhKBOCG6h0EK3OtHM/C0jtLCZEhSV
iiq7phNW7f++wHq8LOuNidX3RlNLeme/6N3FHfjdXFkXHGFiQGL0PjCUU9s55Igp
S4HZpw5raphPPqmp0j4GKTInjtmhyBJhw8nJL4hN87zaIKXg0097EHSpyOQ0wh1t
puSg1hPgrvaGaP9EijO7Tn9tkKDLVo+Pd1sBnONKqXxaPwiKRCxT14b5G4UNjybV
mkU6dw0aNpm6riQmW7LOxtGZLLowMghGH3JRa32skEfXv41iR1cwV7X6oIKTRHwV
2h7VKHTTxJlc5B0xz/mBzXntrWaRDNe8r8Bdwe6awFKluGDIjSeHzmOffykz6SPr
KCF5H0Rlt7/LrvxUn6Ir8l0Aztz6y7rtXTcShSZAs94F8gHZSCUmZnE2mGffLRtX
sF/+0hU88V6F070Engvp74TyiitcDVbtkP6/A6vD0tlbR0AzqwDiyBiuq8363VNT
rIUFt/HmkqTBD3zvjb1BZJ+OeNIcxYjt+0DGa+3qRAl3Lo2eUGwC3QFfElN6hc9e
OjVGLYHDG2KkrjH+0OOwQLxXmgRrpZw8uWtlIJhi6iHBhzB+NN/+h2CzIaqczLUh
PGYVY6dIlVWTvc89ENzurzR4UW5nqo4Da97eawrO4dKZbJmhM4po/bu0GchF55n0
Q3doMuVKqnCbqHAEgH4TX7+xl70K0DFEGv1/I2HEX+X64W5iouaWH6jByF4WZ5Jb
T6NRY11Q+ms1NQw5RZ/rNBR4kL2VGQIFli4QWgaGa/xcjhwgVl/IP/z5cy1Ntpsi
XJNoCdFQCHu7TJm6gMr5g+HrvfcNcXvDedH8EBdxIJj26bd/C9bfOd5GFIHqj7rd
LZa9d5Ugx9JCWIUlUidqxO6n71kczKn640C2voy/plmvIZuI7Mlx6ws/ykHyr+WM
5EorTN/rCuDaVS6a7uXEJVOTKRGtfhWtms2if0wW20WDhc0sgoBFJAyvps4Tpjcb
gsesG9d0GQM3GRBwOsv0JFaqDwGTK2i4x2WANcZHZBP6DirdbOi5m2ioVSrXxkhp
0nn+NMmrgwtjcqrjusK6RGaSTfpifmU5Qcaftz6St1hRK2600Xfe+fNRE2DBKZrG
u/hMdtLM2MViS4jppheQGSiB/MCZGgaY30PSB1wRoxaILNOHCAZDvd4RnH828XfJ
1ariASyJ34bsRm3oQm7ykPYCZiMxOzrQho39dwpMv6GQ/UM6gKJ7B58Wk6Sb+dW5
jXwV67S8WzfgoDH1HY5xi2l6uZl8ZgiGNuLng52rcfRtRqmk7uhJPSHZSvRHg5bO
Q4i21rc9wWeXpYZotHyX6BRyXybEX4Yf65wWXSAPlPS48BJCSFV3y1Reg92IH1fb
sK4olYVLlHeRotefqUQlwo+VmF75ffOdN8HEqWRrdZ6HfZP1m8yC05HPJXUqDBt7
K4BO7t2qMcGOWUTvfu9jSH10fx6r/L3Vk+qO59bVz4DrbOYIobbGMKZt7AWuzOVW
NIePB22Zc1mLDygmUPVJqm2HjGk2IynOL1Wg5ExnSsmW/tkyV9PsnWo7CYO8Hxhl
eZYsxjvl26B1ZWVem8g9nj1t2XiAu9JljSNg4pB/RU49uUfCAmBlSTuml6A1UF6j
JIHTRNoP6dkd/J7nxVZtExRBX4Lq+9yTGnTGMPfXHtFd1fz7CR69BZvjOEpnVyrI
HCQLm1lCwecTrbVb1USP1Fr6NzFWisYg65w4K8d6aKoFHKO9lhmWyqhEOh8BzPCH
0ag3nG+zv8T8BH4tfFEF7ApkK0Tp/bR4/m9OI4iSxoqraX2t4mo/3Qy4spMSYATb
6jo804G36WQJecpZeM1dbEKS5ENCRvSjU4FQYcToFQoJT3g7FKaQlbH8wCYUd4gu
gpLS2OicHYEGgLgpK3FTAHLqc6+N0krDWcNRXBabXTeI5lmYUsIwRIY1ZA/bHHzF
ifAs+FrP686VtHCtfNFaStNAZH3xS9N/998FsSeEQEB1FpFqDd2u2VRMAED50Pk1
TTbkw7vdzXKc0Zdxiy3gsAt/NtzjgaOkygZR8jEgd6Vno89mMh5bSBqYCc1RnjS0
qtAHKwWvs8q9ODcypnwIAelCmBuPbUDzOndgN63w8NvCSAKMcTRg1gRNHGJIkJG1
6BJtjLw0yf0SGs6IJ7Cl/GsERUD1+HeTm2FPice/dFhc2fqdm+vx8nKqFVxt2+RY
qp2TRqrJsiuOzfms65ksQbTpnnTjU3f3vHSaMND7jXDHFf/6trXHH2UAyvTfluKv
5TRihJxZ92MUdSq09kULGM1IG0cqpEUre4E/lIireKj8D7tMEGwWRlDBMY1LU+ek
vPxUCWXYUXgGTt4YDm9nVZap+8B1n0fP1gaQo1lErqJ5VABJUvKw4CnpH4y39jOI
BUMRjWDueUO9wW6xkvhe5gZfwR5U4dE8+9iD4ZEeyCIP4OCBcMvoX4YX6+7SXgy8
IA+Dn05nuA5OnqgwJ/Nmhph9BKVR7RO6Y0vVAvr8ASOkXknqEnsKZmJd6ncQbOOF
o1Fip7b0Jiepn14DtRJIwFt4Ez+OF6cmyx6vQLew41d4scKu0ScxfhAJbbkOdVbg
Y+muHAppRpKB89VbdcaGHkh9B/PM7XTEDejjjwQ40P6JJPnCrSF9vsXPevetstRL
Bqm8mFE9CQGr2uMYXQrOV417TxC/1BLaOpJ0kHVo6vjIO711OYtCxcVObDsOYoFI
0RjhmaOz2Fy9SYWl8a0lYXBlvWsNaE9Q23ydiul8hpZkyVMGZRJPk502hvkstrPk
h4bmb05qle/6jqdhwkrfya7703LbEDPtoeH8BaeiFBF6E4M2OiuPJfsgRD/hCmS8
rxs4nWjQwjqqPQoDW9tk+AZjsbgP7tJ6+aWPobFESsMAUIsoZYGCeoxuMihE8sK/
aA4DXuA6QviUTTMPDyGTqCFeSaxWHbC1X8GWE4ngb190E//QDpglW4O3hfJ6Pnb6
JeXM9ojWRwDdtCEQm4rtBjsMRisQQQ8G5t/25OytUekczUSM7Zcak0JgRmgk5To+
el5vP2X+IjLHnX6ctzFApV9FOcR9yjyIW/PLkG8Dr9yCM5Zt8GHyCP04QAQVExYL
q1wqbO5FJF/2lpBhP8Qb3OWz58TJXgggnUTLMT1QRMTNbHNTDnxfObMq3oQjyUht
OPyqdILbalJceEnNDmkAZG9zLMx5GYrMrLdE+xWxhjnIEWygzjvRoMFU1HMo7Nvx
5fzipshCkEsXtbpVHp76iE+aArbAYaCOQrP5HD+kQr7z5BWQqyuOkwciYeRtpRlj
Zy49Aa6hgsHEOFFuMmxdLHSlQv4ONP8N1BLiUPZNj4GiFO96rL+TWOdMaWWbYPKx
Q1xCcDiFYVSHPf+0T3Z+bkrnO3OXx2UM2d1J3BFHTg4cCVo5YpVJltQ3SB8uisIy
YvPHMoYFcteotHjZJyY8T5CDSWXOFyDBdAUzdMeNX6oqI+isXaEBmXe8570LSR2d
YUivNB/cAdgVo3odm1bNXXLN8yT15uAhw8QmI6OXxiFktQWFd4EOCJL137V+TssQ
ZhxnqYR8uoYUdIO/ExHUHEAH6Um/kIrvko2lgnOUJZVVNyuIUeT3/WWty2c4QzY8
H4r2R0mNrditF3b2YrxP7aOCuguR10DhBSjgfj2Qcf51474Fi6SvBB8GuYQncSld
8HYx/8p78vG0jX1uzk6zsMjvschWNwMLT66rYfwgXV2Kx75HgQ3/s1IBOdMvv9x0
o63fQLqXc2IxZnpxnOmlNs79Yv37+QGqsZU4PVFULlfB72KKEovRRwmjuU7jk89o
XD/CBY0OoGgcmvcHnk7zTaz+Emj2UyRx+vG55hX6fW2GubbO1kyAh4gAljAlv8WN
pdi6+e7x4YFfDrUpOQOYW5l03nuJ0TlrQEu1tY9liN7lJDFh/ONJSikniVBLwmP8
q+XuB/JCFiB9hU7jRbirrkN2ix2PbfBVFjQKqpm5erCtON7PXTtAk5SBdr08r3Zd
cnlz9EQeLk7uZNTyEjdZVL6GCbP9W6cvEuw8aQJbgaKRHUFMM98SK9LFrPJrDPKn
LRMbplrL601shDbTN53tVU6aB9hwzlWvOInKlPnKC+DN0dVEvNBBVGHxYBQZCJHR
ZaiJCEmcoJQ9hfk1RKUt+uEDRw3g8Fq1LtkDpHBD0l4mTZSVWu2FuYYITY7TXOep
5P3Ru00nBtIf6v2KAyOEIEL8ZwB4qkY8lyhs+lWsu/qTKGyF5Ls4vWAeDiFBeAJt
MFhN0mPhLbwXkqPKVcmR1Cr704TGLhMocjyj2gQWly2jknTTutDu9/rrCEN0jUjN
YDtT+YucfAn2Lw6XB+xFh/d8/MjobcQNQ0BHm1EadTocMZCKpJ1L3X3mTzPJxJXh
42V6i81wQOW72iTyebF8KQyvzG75Ad/4i7J1/XloTUTw5cQz0PTXw3QFDdFDL1FK
yj1ub/zOtGAsfS1Wgf1EsbWH/c7X3I25Tv4HLdtcLj8CcNxZKxzyMjJ6EmquiKRw
Lx6E1kQ6GhSs+uNuEsbKfMiCx69IYJ337NeqjcnEY5PbPz5VDhez3sTq0TMtikL9
H4kKocIv67uTTPysMGKjoH/zpNDUfAEatcC9nbUuLU/YiD9q6LcANdzgDO5umRDe
xUNKR1+CfNldKpyO/eLVd051ZBdHEmvTkBSfuiK75YsGHRwkDUzbFZ0BTs6zMWea
F9lQ13dkmu6Ujt4JZ9nbIOEszjCWTWrobw6YP2/t5aqXbcn3IbXS3H0T+7uOkgey
8cJ8qBDW6Ol+GCnztv96sIeyq0gu/BOzjFRrxVcmdURYZMxU6BMvuemBBAZdqKIH
bYEI5zBuk96DdEkmzsjdvYrzx1QOhnf6X+Q8dieezyjL1qWb93rIr6mguYmdxVfk
cmSKjzv7BXX7Kv1Pl/XXbYC7FOVkrFm5Nj+iK+VIydBkazNNTEUiQIba+voNBqru
EHXMBYVP0fAMByGvEZc0q8++7JtsMcYtGY4tFz1cNrweKDOvhb4ukLHbZzxxI9Fo
3ePadA39wQvdyoGrdsxhvfGSs9RFSuhMpyLkKJbpjTr9KS3/4b+s9aiuQgSMJlc4
JRr7YQ23ziAzPqzIgXTkZb5XeKr5m+vshP+KTPPPlot+JHjxXQq1kvXzYbd13Dfw
4Pio33QVdowpnaMMThD9fLr6WJ4rfW3b1Uq06lcELq47lXa1WFeA16OikCQ2Zzsr
B73rpDW1ZV/83UTp87w96CRJIVprwTdsjn7E42zIl1dEyXZ5NoF8Qrxva37FvEFE
gT3/cpl19H9O3LWvOxKErDEz7AwhCNcjaEr4LsFPJe3/c317FxC08HWLw+oWW70i
Qx4dnZBfRc1NCGxF51Ch2iAwDn1smM/tRK110+iOpKhKk58Qw5ChIqpF4yKF1W1i
xxrvSt6Ij3cpQpzN/5VCKZ+gIZfiDcpuKmsuQQIaHc5p5GNMdG5CXcFvsP7h9wAP
7Yy32mLzsaylzBYu2NhKSIYNMbJKJ+zBtJVRWYlF4EI6+huZtLnLmpk2pFBSdQD+
sFM36qs6vvq7GB9z8T/DZMN9gxs+pIa3qkxihbpqztEW4Lqrd2ap+a2g4ZhByuVb
9l/cMzmGJpCZRCR+M9HThdmUUJOfnRl4ho1X40TAdd9ytEbNxKFt/FzmRtiJ0jLg
QtDY1Au3+2c33y9ZJagNgDLRM7dA/Jvc2a3kTzX8hKj3OOp/IuFtY7JsZMLE2oEG
K9jbl6wdBnz43Lner+Evsk/K+yG32hbZa+tXvT2VXEhbP1ZWTpR6WxjsljqnwvJh
IIu2PUHuN+RC3uHtvbyMWIN5pMkj0R+vuy7q5M9Cg097fxluukxyjRZAy/TU5Z05
/3Vay/kTg5A1cjo7mSs9gyjVN9UsznVc8uyWPeh9MnhoCWx7M45+YKu3ioKJgXCp
SSah6qTH1WM1+71BBescvelwIJS5Giqjqk5l0nStBVVHyVn0qsb61oeirGaTT2lA
xy/BNFegI4ZOFQifSU7ZMj/bZ52yBDmarKlLwO1D+08u2EtEzFaDIXa1Hd24fVRw
QI1/MTqgGadXli3RrM2ZGw4bzWlB+4wppP8NQq1jV0EBVwl1MoW5t2n90exywewh
u9xjjnKEXK0AX+llNGLzcm3IeaMT+etgpnD19PvEgPVSt+lPqz+By/dERdoFeiV9
7nKJrxO6d/AqBw79FlXemJo7b3EXa47x2ZDk2S1i1OGjNiXUJdZbcsWWZVlPAMrd
s1z/iXp3P++40fcx3sDI7gH490k8hNxFJZ0sCc6LX13FV5gAhJkZXm9MOF/g/ysT
P/J4Y8nUCDF/ZckKg+7goJrfJPm8YwfQF+NTu6575C8ySHZ0k7Le9gDPFReq3K11
7e4fl5HB4QvNSBEN543jW/SA3ZN+x7c1bb46d2OOUGAbsaBfRZowwOEew3FhXyjk
2JM/5Po7grBT0OV149A5s57RZr8Zq6+fqwkUD72RdQfZrytxI6vKBqVjYurEs6hX
Y3bHN5lG3bNjvq1LbihXfzvtmD9IJIJV6FPVfo14NRb2c0psFiwebj5Dr0BS1BzZ
24qCuapsZ7p3BgfQoNx5FeLywHtFEqFplv7EEov5Jp5850tBhLTA6ay9bKgJMDtE
YHj0j1j2MQ9NHbbwIfunrYi/b91GnuDxdOAdkk0io89IjWJol/T0Rj9XuLz4nMu6
01IPaWhnX5mdOqDZcxzTy0rDj89B5f9W28JzTTb6skL380upsFZdF7d9A1exlIhd
UC/SMrJaa8gY+/4ddnRJ921+BPXYi+tHmezAPADfgECQpfgp80Ng7P0x0Ky2AKNd
/gkYP8oDm8g3Ksp8S86sqCCyYLISQG7aXClsXAdrts961D2o/z3TBORA79J0qzzK
rCQCEczGYhl94PxUzh8MEi1fHrCFBh1HFImntV/LaEbwgA4VYfg/evFSSxSPrI1w
X7fEYEWkEbDc0SEGy/5ASaQc3ZanDBSHCKqOx8YQkVbPhqsjQQ9E2c1SwKKgEN2a
1DIcZgORhm3kAP8q9pJ6//tGtoLd0hBdMzsHWr75hz4v/wYm3Tui+6by1OZH6IyC
loe2GsmL8U2x35ES81b6yo+1rtUb0d+rc3XnNjjosdsAXRh7TK06RwKZ7+qwpBnl
F1gt/frb5XZwfaYniTIfQBOOK+mytq2FGhBvdYC1BrzAu65FMtCKGJ2u5+q1nWJS
NexJ5IJYayduex7rFZkTDOyWXh9s1QoETPml4HEyVxocKzeJ3yhxibgwIW2upRyU
UmIdp0wAear9GSZG8tiYFAEIdyNnQf6Q9AtRmZ1Ndr+1yO1NlUT35/NWxCoF4O0T
rGbTo5jdo7QCxeW8WGmDwDnQ34dbmxRzz1A8DYzo0AKwb9uaA4VoKuVN7VI+NOt4
gfZKk0kftW8rPPDckftzYyTrQzZGN2hnhktTD1kDolkLhGNlZZUTNjO/QAk0DvDm
sYzjnxP2jpe5wyExYtwBYVQ85fW3Grov6aO/IP4+tkwIldQ/g32wPi3BcEQB2BGT
s092WkVLtFlH+t5RvK9arOg5BwcN/ohl+ipDvqgs9MkoGCnjKKLcJR/jSglvWYRF
LglmMJj3dAyqX04/bxQt/pA6GlwX4ENm7uuFSHRCI4reYfr/HEgIYowwVTZrj3m1
Cj2tnUTTZr4iNlz4Wj8e+yE7HaSV4L/OUpz2thL/54nwOBxWr6zhStdYrWs3TroD
feqOYuPSfoFZY3JvpQtH9KMSagxnTSUABqO1mciISpM4FIDd7eMSSLedzJf/AzES
g0eCd53wMDE2u4rGrhjzOVnnQpf7zWrqSE4A3CojbHIfQwbj7+0DCYBOBMtXkb++
/c27kEfGKi/rWrHsmXBzJWKN+62Nt7N5+KBSQwQ0f2JbFyNT5axVyO53IA5snw32
BfLmqGUttLdpNRksfkTSL5bjrOQrzvmr3JSJDL6+rliC4g/wdmZHLCdr1dyYD6Tv
XEJI4BbAcxjJmIGECQ2XjsUwBkLdz/cXenZezVgdAY98h4XLkncjXaag9wghnNKd
n8F+Mms6gAtLTGHD1TiOFOY08Nyj9T7WWUoXZa5COL9y8GgPBe8HdH5ETl12NMrU
M7MaFik+vtAfnuqJbStM4UjkMstciiyD97LiuC5fzrVWV2yabhwJV3r4z9HLRphi
QkfXNEG/c3OqZxg9hv7VHx7IPrRG3XSyirDvcd7ZTCH5mCE49sUD+bxzD9OG9otR
QJHCaiKxA+kvJBRmv5E7dtBcUvsxdg8PgZGa6+wyk3J2B7zuQhVrHeaBv4dCgV9W
6n9vYgxgF/pvkbP/IW0ECNiJAmxTqcYJJJhAN2RbJvmtAYJ60p/HxjbwhPArmDzA
iUyzKwjF6xT00cPzXgILLKiv1YaJhI1lfZm3bq7Bj1gHuWTHdhIKEXMYg6SbWWAz
8b9j0pa1uKtKXQAuYPAclLNg75gCEoVyX8BETiv7YNeei1dHdX8Pyd7rxdLLPu5d
RhInJZKVzqLAkGulGl09XWwNd7Aed+VYl416TIsnYalXnI4gD/T42J7pJ9gXfHTR
/+zOLg5YRq1rGr16bXvnfX6ptt9r2nSVqTCyUVz7FiFybgtNyrw0+p67yjh+NYJg
v6IjJ+xPdq21bIrVVjkj5tweukY5ViBmY1EjZFURg0qxhho6KjCrXQ25qtA3oTVr
dLvwwoPCoodJeozC93fVgElWLfwcpG6HYIWGzXgWg0FAOKqLRFdisHog28khu0lU
5Yp1gRwUsCZx8TDICvtIBGZL66RIfnYuEw8r4W6RDLp1/5HKaJ6bDW2YJ6Tx2O1S
IYyw2tmQw4vC0GCelWNq6I4+UG0THKZfqKxFNvFteRKr/6nzdeVdW/8TYADr3hkn
sEjum5ViRw5W1AUpCKuFji/2BkqfXqg1ObpYSLNPOcj4WaLLaky9F3dmb1pUO13k
mRkNCgXPc7IMnS5iHL6DaKDn8oa0M+MkK7w4fE5VNioPHuGiIYlpE7BNstaHWRjq
74Ry7VsjjaBXyBLylLiCidhXCPbXmYTqrKvSOq0hzUH7Ol7TmP+h8MCjHa1b9r86
Hjr1kfu+2fkgle+kPm6128F7EMZBAscm+tzynMADaXbCbMx/VuzGnwhMan+Sl1Yn
CnETtt3ktemJA5Iyshrhd38RPyhLqt0kk4wyj9stNX5kYXS5M8jnM1adHSVEpkrb
+CIT5+TuFgTTa/U74ldah1i1QE4kAg8IG6UEbBjB5FjOqxFDYGxRB4PDh43gGirK
wEWadvadtx6FTZ7QGYFfKX3M6tH2NZWUBpszOYDianIZbkLQ4Pn6b6LMc0m7vYLa
N6GqZOMpqVw3/UpCA18MfQL7iPPmeTVwq6d0dDvaCk6cKm/sE1JR+UJTdo4yjz99
zMI9sa/8aqXQEqvoqATBKpSHahw1yUBsg6u2/JE2ChRzH37+kbviYoB5Xk8sZ3wh
OftB8QY/4f9O/NlSr5dmlWbmLscj6NkatZbOpbCORer+rSlxhiQhkcl9af5tbcP7
BemR0q+vUh/BCVgHU34eYKlAup1C8XBWMVElAk4sg0wsGJ19MgniKhQPJT95geqO
5Zv8RgQxJXriH3GEDZnAWUG4gQMnxjKcA4br0M0Ipn48YTluE/3snH4O45696N/P
KKkC0Kg+b0j50RFVCgFA3xACrc+zcXRZnfjPAeqBqVbEnsTfa00h9S6gNIxByMQN
zBd2plpxlWc6WrGKkVMloN5Hr5IvumBgqwFIJ1a/qw+Oh9kYlWkLYUcWTiMQ0yOW
B2TKdP8i1SnJoYdmudIwIdmZ2OUs5SYv+v1Y4LB+DunnxkuE2m8X/36IZZnGOlLT
2bSh8qtEkVSDNjLzFXu98x9EYWPSCYzeOKDSoiZ5zwLXg6kouD48ND1/QbPYJ81U
Xl3pO3mRgQDGxFmE8RuMMCM1Fe16SLegDYJF1UaGVwhqabYxdrTNLKWkcwDC8kUK
4dR2gijkkRzwN7MHY9OZjJXxdB2NkqXriS4oOCtPs7hqc82ywHlhKn6tKZCu0kwd
x5yKhvcN2839kvcdMb864+UErpsuwWhzHbH5UNEymWqvTCChAK+NB0YiSVWi3uJN
17QPLgD14kHCjL7nQWiy1bC4y1f62jEkeCNUtyhxCqFjGE9mpgn9aIKYF1Hx04uS
giMe8qYHhKLtb79CqnspE179RK3GJVnp08SFnpaZfIISrH4LeIb4Dz24+HGggnCp
02W7gXIWxVnTvkBKE9STCHcqeLw5r+ABaaHMJ3hFj7GUe07/bAgA69nJqyWrKOua
GNKTdUU0fNUG8xMAcUbEf7UEa23trFXlkcXZDWjynA7BM85fXpPB1ZDM35mSeCUa
TyxT7jRnsPUY6XNHyGfDcnGEdUQ8YDTfuEQfdV70SK+sAoR85xM0yiNXX3p51IS5
3t/uHNrDWIq7wV45go7RITUXAyUzIDTplN489T+DDBAugRQbGgysur2wQunHaM66
U/20sJBWfn+5CCO4nAsx+rq7C7lw1WXLYmFkSODXvpxq3tLle7z2fZMnw+BG8laq
QfAnjpVPmBOPVwiBVpEVnxD1jW+VOuw37zwjvhuiJKzlDJFoFiu3w4cObBjuk4g7
nIYtq4nvl7hhCcyVzytLYPXULMjzuMBQhf6V/eFi/u483jhCvyKju2JM5IW0liVr
+2ietiMh+veZ+2vLh7Oab7SVtKzRM5LbOZ6OngscpA21Uae7BT5Abs+37AVZOSeX
Rk6BEiQ5GiNX5BgUxFjQMxxa/XkQvKbGAf0yGzMLDIUHkaRo3A7UkKJ+1fUunPKA
YRJ5YaNQxzM1P14dhyx7g3JRzoU/I7/b4S18K9hmt4Y2d3eE6D6KJBKkBETjTxvC
THii6+3Myx+rKwiSC2mBWyBjc7Cr3H3Tf0d+COjslRB6YUHWaisAf1mUwBnh9hsQ
E6Z6167eAL5JS3hmjdWKao0raoinb0HXSDDWz+ZviGQ=
`protect end_protected