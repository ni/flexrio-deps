`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2048 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
jsJpSUcQTu7cBpkLybExAgmKddpwXj7oq33QPLSCjQrSmgV5WM6gn4vnbE5c5NwZ
a7xmZtStoUubYUT9RfEmDj4bAH9c0JKch3//g99oHDdbK1Oc3jnjtSrnjVMd9/D+
3WNAfrCuVnClmQfsrt/mBwodcE3qDyHLXVVgRuay2/xX2auYUO7vtz04oG1H66xF
V81jcZ1gAYIsblwlRk0NPtx+fjDp01UM1eZm+SmYc+AYq3tLnZivjIOrNk21Q43u
dR8hqhxxraljh4fBw+Pi5DqMDjYml4AnjcmkVmMYGTpmvkUH8+8lqqpgeK0QippN
eZqF4qYNtO2Uak3MZ/PAUlHOdKa6lvoLJu27q6oXljoD3ZcRoSuixBZjbFCuUqPD
x5qBbvfcBreD8I1L5GjX8IwCagOoDw2VvrnAurkDYtzljr9nq4Jp96RQubk3Xnof
KVuRe7EirKun/V3XJoQy0aOfSX1fuO63USYP1+pos9bJSogc78u+x20DwTui9zM9
CT0Ov75vLV9JqBjuBVsU5mDhcpijpwzHIRa7apzhomPL6DYukmPcPKjVayo2BMJy
F1geHnDrM3S76qeUmCfxJ7U6m2xKb4AmUcEMWXKiMbiBqkbj4wVYsbSlSTAj746C
/03N30zYFVTmlttqEOgpuYAlkkTo09uTmjEK5r4e1Og5P8MPLCQvm4JrpZ73A9ud
WNYl4CMSpp4lu/eyemOFdhWdBQz+gJGwnz2wHTks3I54DRbPtJGKTmAAONubE1hJ
MMklOqDuyVz/k08Cl/AQK0gnBbzKifub8EC1kkJDkD1Hnjz8fUZE0SaA9hFOwVCN
L2bOlVjJllFWiQdPhM8jgC8YiPG3UX5PUXRVYWV/J+mKFJ3MaYM7tZIgOTmnnSAk
tP9fW4wqbJs4J/bcPUcum4u6OZu8P+Ck8SsaLLHKdIayqojQFshV5FQNRsOzis7Q
Xe2HbJOmYE6uYU1Vcm2E4mrvM/q22nbWO+dQi5ZwbN7V65OYSADSfTJval0rOPss
jsIX/xlnBE6kQRKMVo7r1R318hI55W998nsrYQ26oAO+9lj0fItN4iRgiBEF5HGO
N5pCjmf1TSfchd0i5yUG15oX7vkaBkqYWwlRLnCbWKf9iWf6kSArJyRDTAaY6gaN
y9ljq3R0sslNIYXQx3P+obLPpBsVcsWr35Hy80ECvGFvjw8ebrRQ46pg8cWCL4J5
Yb4QnCnYGrCIL7KkATBUbBmyzPmpHh4uJOlljqnPf7PsVG0LQDJ0/9qSvzi+AtW9
s56OtMCQ9mbrkPbpF+iauFZMp8ILrBTH7AmWdM+uKvE0UgqdR1pkOFuV/MCxLSur
bfGzmtRcUgHLcAwBVfUaBAQ9v1xWjaFFUogKNAlF2izb4ZddHR8QB/uGZW9P32vv
l/BEjPSdfI8BEEkTUeEjCOaSlaQpAZxuB2ECPvqnJ2EMmRnJK8SwFd6iSRt1Mx2B
x7uRGcBv8S5sENSg2zEedvXW0SRwFudzllDIq1Y0I3sW00HePIpxYnMUmP5Fqx8e
WufpJO9Or++62Rv5uPUlVh33rC5k9J3caaYR0wtEaqkcA53ccSndq53ZCPOYlVWq
izCGoO9falAzOoDmEL94K4fHl5okjrY/fPd/QY+mTFrej4n2+F3KgLCTS5BKFoEx
ZG2m0Ht3oOGV81GX9m/T6BnILbXmVPaDvgS+wLJlvuLCS8f6v/U48vYIqWLU55Kh
IEVbsOBoMnuyZVnzp5SBnlYeIWVyDdAmk34BXGUjPkRD7D4dprjy9QA5JCCvFLMo
OHhLJI+64UxmRs7qMUWYrS01w6EeZ6+ATMB970ytG8j4Z0LZ3JgYJ4Va1CeJ3YzI
22h+Oh3Eur7Ktl/RjSoTC0s+wKSYhEpkNiLgeG9T6ZW+kzKHvqjkD57CZIUpqlcp
zTjOEiwzE1hYOpSfxySd8QxesaAe11siORGqJkvswdPHudxoAIYuR927gkEkb4AA
7Tyw13/hAcn/j7mMGvGjIYKoRNIDQ5u1mbX4a8sCFc5eSlCqlllxLAr4YXFCwLIp
SHY6txtXUXcI8RtfDmApwiljNaIHZ0a4roBcwp/iwLKnAXXoZ84a/T9Pwzukw6dy
Vp7QA5sTs+U9pHUvmy3oW9T8an96Ka34gSzWpDSAgroPl5gEX/tXEQAL9TztoIu4
kzUp6VQcKfp6ZW+vIrQkoovmxfAKdFchZkMuhEskPlYb9MbDmq4KvOhhzpqlxsQk
/iO1jmdNLJoeHAOvEXCtwjy84a8zv4i0vyS2pipgIwuOCgHuYkKMflGEMXfj1OwL
uR304ApSZtrycpSUPlQtzKhIbIsCmgACyAZhvvOznnaOxgS0l6wEn9UaoXxE0mqu
usKK5p2RznghgNlcUoTuSJTmxCzvh2lEnsTMIMXX0dNMOS6hQvTbyqcVPqSdxYgr
sKFY0oCptFI6HNBMQ9rIltn2NV3XenTRCw9rfS4A4QNw5i6I4KjoNuommVxCE81Q
mCFQ5Ji7XUMLkXhjWuDD4EPt5z6pPbqW/3eppia06yoB/UOENqitMfDVxTRtvalU
zbTSdlYtUUlw8JjXfcNnosYjvnhQPUS4LTTF4rkEDhk=
`protect end_protected