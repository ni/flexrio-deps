`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6048 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3aOAnDl8anF9DuXzU9136hz
pzS21vo9H5TsKJwCQfvrp2iqwGGFgb59zpw3qh+717fWKDiFK344TRwB1BI0BXAg
wqn4W+/fLQKWmyTG1Q0x28LcwtEuRPAgzZtLSJSCxOBel1cNZ31Iypt85XtSnO4A
xTIJhsW/B5wryN4l2zI7RYcGFqOvfXA89W7Pxemk5B7+wFD16x2g7JGndrKg3ySU
wzwpp8eABg/pf7xzH3tbiJf3R0rKSHWBpbIJ6+9uMRckpO7MxEqYP7OPJj3r/7hj
1pHghrGazfxkCDvxZeWEe/9yeooVJUlg8R8u+majn+hV/c2Rt3oJ7Q/jeTe/Q2M9
TCkshTiGBbXU+RJ5Kod1O4bijD2u9VXhYn7FUTSbK34cW1kqe9BR56R185Du2nvL
LPb6GQV/sL1h7dzO1QfWaVe/+VXOXn7v0VR6HbxjQe5EPeIe/IzTeosYlXokcF7P
4PzYa9SPXa4+h839lw0+LzkcVtzytIQBe5Y7P3/0xNxkHOxMOsRjDtuZrnK8tqxu
1UfX0G/4h9eCGVylFJBzBM2LCw9vuqO8DEJdJAzFQDo0vzfnyIHDAdB2qyWwq60K
IcQ8aKFgBjKHqdnzapdZSR+B+ZjRMmwXUFCUuZEvutYWHLIJ1kjnvzUMZFbAncFL
tasyOScW9MYFfwzB0uS4iTVDk5ZHX49arNGf1J+bpjzOM6bpMfKv1+ZumEn3l/gS
Xptm4HfXBruPVm8kDT7tp2fkRLD5RKNLTUBofHkQPo69nWn+Fv5UqNTCfIdmueMC
gB9UC8FvOVkztG6nxWCN65qUjHxxfff/CeR98UwQ8Y1l9lSbxBhHqakhFtlPa40f
JrqpWhcJ6b/nu66LSyD1jsceUBlQ2GfR2KInTp4a5fVfxh4Fg4+PC6TItrChdqzx
rl8MEsvibERhb/ou22uJxDOw6i6pBaeFOUfjOcg7t+o0xXEuLmPdVh2TY9371BRM
FCX236VMj7pooTnxx+3MVjnvnS5SK9x9gjrc4fvERyMiVZU1ytzizM1gkgd4E/zv
8sQX0PfXNL/7OJ0KW4853x67ZYr1Z5+StAerJSG1S02cM7nl2ZILLLJkqomIyG5h
iUgs+GkIKc9PZ3mUc1JZ6/S/GHLPygiUxmIjTFEPtQCYu3BgQq8l6GSJgwujJcvB
4kJ3Gg2aU/Ihi5p4HBE41tvOZklpmHyyX7jP9zIEO+Lmje0JZRHigFksvmIex2bW
lGfpo4k++Tez0wh3QjV3VL+AVFuuaJqPL0wETW+lHOjGpPhubgXwhlqwcPStKZWj
ng7qXR1EsX0hCk42teqxiL5GmFfF82X7K8esGH1lzYUjYgthonuKAw8lU0hlV5gG
gKj53bIg0+wGXc+2Mkz6wkrrQ8kLu4a6gAR1TrR4Cv7MiNTDKaiewT3q58uAMAzJ
Bzwkb/RwS+nQ7UE7rrg8jCzYFpRkgRhoJc6X9NJ/SYfsNbNQOIis4MEVLhiUWU8m
Q8QqahbN0/MAr53fKBudEAAk9j0rs/rNivA9m3H3hDrvaGggjCDobHK/1U6V4qA2
6YlyW+vkif+goGzKJQMJjNDcfQvGSiLVoHAnn3gwjJKGXTeb843mLvO/LvIiaukc
3REsdw5PmaIaNnxRgBXhkgUsqVHa3PbjaBlNS1zpHAFOcLKwzQUYtrSW15nIMbgs
qS9o3V94NKir1jtWoYJDSgDfpNiv7yJt7RriGUO2bq+xO6yoKO8bQTDc5Bo12H14
HAv31M2/S+LA/vzwDK2XEuICJ1/evNAzePXrU054VkLdQVTNRXKJo+afBNcFLOzC
Bgrasqr4lhAARZrbGuY7RcFGJckhX9UfR50DTZM2zDUzri5oVFyTRkaMpTIQbhQt
t/iqwUyKC0Df1ufj2ipDgGzVP2t7vu+ruyAEjyiFEO3myuVv5zEPIe2AFpQgCNEJ
JGDYixsgzldpiOVKoN9oflTuMYatMnMIpY9FwE+kLeQUSUiH0NWFHICnNWx0Vn9Q
qzclAN8NFjNukkiIBRdgrl2Tit45H0Izp8bzDVoFu9xwUf0DajLt1NhVv6KWaY8R
hAYN1LLotoJHlM4Uca8TYVbY9ZMR2+oVqTAqgPAnPot2XDPkuFRMoR5AbZMerwHg
DwCwRTT3rSTdNhx7FXDwSCqNRMY866BtsEMrfomAud0wAd9Byy+qQm8hTQDxrpY9
y2REqXSUzWjtq+vE9zIedC6WKCBCwGKAkOV6ELLEUotv/bttQayOh4HluoTZB9zL
fnutWTZTPi+vJ5CfqfanPHuH/y3bG7VBid1x9GF2Nk2TU6CDPKKBIz5fk0QyZRat
Q7/E9UN5vmiA5yiWobDv/Df+2NKj9ABYziToenY5F54+R7fVYIaijh7manu8p7sC
xzz5zpZXNasbj3UO2dXMF/1pK409dbrtQUrGNHC2EdMNLHJ4txyd0mmxLES2rzsG
H3LdOMaXyZh5FoQXcst1B9I1Iz55fOyYQAsNYE6fhdfDhVfcLUk4tWahpzTo73bT
PU4yPmsZsceIph36vlMEroIxZzzlRkmrK7FkpGVVWoOQrZFL4CkvzkZb6Fc9Xyjn
LPhZWCpRFkb9uhZ7d4pvGSUkiiqaMMAhHe5609gemfe7mAaR6K4OcVRoD+BxdArW
0a3DbsjL6M/TtyunU5iRg3n6NgLx7yNTiUdrqzr/MGywbeubvS7l7UFs8iSJY+Bb
S/VsOwWL3zRY6p31teDPGf4zQF9vxua+XTXQ624zhfHz+o+RYjqM65xzidyVy3bv
gxbn7qZzYZVJVuCqgm/Hvg1SCzsg4Fkb2oO4yy3sdUMv73MJc9Ba6ka25Cwa1D3U
xPZv1D38wqAU8i9lu9dZ5kAiTp6yyVKTMOlzlTzGlR0/ARw0pB9CPOar4Ese7doV
GObLwLikYEt8JqEMfOh1rKWX+97wq47a4vjvgmFyyWseETSHFVbx5TUmTkVMLLyS
DaEocQ65iO/Vv3g7UMe9XcllVF0wRGAnJDBIdF9RrTeHiAH6XnFPiMnrbb7v1pPV
rszzQJczFbXExLniUWUsu3iFITdUwyGU3ahmL0VILxR7FJD2hWlN2ZyAXoGWEa7w
/OLb15uiNDi2Fg0L33gzyF2StsEwNB65SsDC70LWl80w7Q6cXzDuGBq+9Yoq5+xS
VaqHpQgNmuxA/1KF13VdmzvY0iG6SNnNM9V4pAV5qezpAt/7mMej5lVp8OS0a/lY
2qK8gidO2ElfreiiJmgoVdYZRpIfh3r0OkQzQXH+cjWuJfBAoMF3CZcv99bJqshO
QuyQm0sZrhXnu3DNST3wII4bsJ7v5DvI7W6dnbTqq3AZ2WBg6ywV8O1znFww6ONa
GaajQbCtud3YIoJS3tQSCJ0+GghCFaYIBaFuOAfCT6qHEY9N4IrWdHCzA853rrBD
Rj8SRZiABX4SONQEWpYxgxFIq1TR8hXEQC1zoRzTuC3Md8/KRSPABmE1ipibCigq
ASgyKFnnZVcIVeO2PCiD+k46L+Fi+VUlzii9pKRJ9SrqdStQiTCEhldM6dYRbn31
rPf2vVqKVPkDkAdlCKrpM5Y95Po4SZ9NivN4lebLWxV73l90uiOM74TrYawtzSd0
GvDWtLZP4DPs2kFgr6FzPwXEdgbh2/GFWfZvoiQctZBTjYKQhyP2v451pJj2nqzF
b1++XZu0c5BcESPMoNppVVkjWfEXcryCli3uz9gepIV+VykBa3NqUE1StgKb4cru
Bb+mtUWd08AbG/302Py2J1/NLYPP+VgGdtV/7sWGF3/l0jY2MBIdwZDNX6d57HHW
caU6ZRJbX9LJ2Wsc244U4/0xnEliKMKww6agFOhw49aPXxo3Jq4vil/xPaKdp1He
hh+ky8KpPJA+MSx8UAwL9cAbsCeNzZPUCBvAL3h8yAin1gVcJMN/BrXVTBzmeZ2/
0bC/K+CfB0JzmQpV9ade2u2zXBdIMljm1JtuoBgxZjML+vT3ZkKmOwvAFBQdjyut
jyH5tdrjrtxnIm60wDe0nJpg/Hkfx8IZUlOTYByRgWv/DCrqKCTxEG+qMntIGAlZ
hZ5Bu6OpVmsfM1tCh3PpEoirIlsCjqWj0nb0m+FYQMK55g+kA1bTiX8tzoAeDutm
h7rjfn7Zf4r1UgNR9QMI22a0OPoyLKieDvIOvZAcD7+0sb8rAHkz25CUJIR8+ieH
pjP+Afgkt0hFocWvLZX30ZwwMkA2zQbOFQDUEiOotDX+KvV3Dq8NOINPuCAsyFLH
hyKJhGqAPVH6fipZPpOnSc38YlGL4B6Ej5g0rlwWus3QLECv15ONRV86LGJMr19B
BpzDAwvFLr0v0TQ5IAr4lZCaBM7EUoo7e2cX0JALafslcOsuDJF9Oj5YelaJxjQt
ihnkHz59qWqVV03HlQsoyXT0JR5/jRH730iuicQCMD02tiL34Rtvsx5zFB+xM8Hl
NDXfQQ39/f3ezcYc7v1LqjaBCtmS0xQwQp4dfEqB4nk8OGTl6By65aHlgu+Eg/IA
pFjp/0esSJSslf2fJw8ghLyRQAeqBIzXp90XBYjOcvktauSthZAU1L6DBxif3XnU
GdN5DvLdGwmMM9QOXS8ZLD9J4LQawjEo+AiP5xwXZ5k1C1D6THBR2LaYHFfgFA/C
Q+D0LU52lPcBNwOuK4OMGqh0PpTAjkZTQxRFgqtQLHR58TwZ3hqvHWLWWtVJPbKD
eZ9O30zkv8riXLLocYCaXILQM6PReo+2FYwkTv5nlftilg2A3B8a7/sQR1zZpgef
i+YaMync8jEoePBiuW8k/SJYRMPxiHtHI6lrmeML7xhZGdrBIoifAtwwsAbWayBp
CI0o39uUEWyFHACzZdlTAtz/x1JMpbw4qW0Ms2CzogACmZO/sBPLitn71AvM74bu
uHgO7eFpLtsVc9ecXys/BSHCSyOpusBqIEM42nDfcSZ3m6nGvs8B3FQpZL5k/+Ya
9uoprArXBbddPCkbJDim7R7oekjFZ8GMeTc0OpWOguBwMtAInQeMqWLpPCNMX1fs
5RRjr5aho4q7zpHapBquajm36191uOkoSRfC5bLURCLF1wbZT9TrJa3wBgBZD0c4
cAojXhPrZO/Iisv4Herag2hBGDzueCdF2tfdVR2tIffcjwCNEOU+etu3d4/f3z1Q
NOvJIT8OiN817YA8CWQApjCkAJZjKBikTIiCGQotANw5N8VFxzmE2iDUJlMFVV7Q
O2dug995rZKKsmE8BQ19JWyaycQ3CRu+s8ERCF98QlpL3pI0zyUf7s4NlHGnapIi
HSjse9T0TXyrQNb9xDxGuahs3GCm1xF2bwTdJHr/wTgII4x/gnRn4gfZKejLOJAk
R0w91GFf7TYyA08j5IH7abQH2P4vSIO0xr8VjFjQmDWMuLNIDGoAwC9l5kSKka2U
aX021kyK/o2jzU0LfWJ0OBYVKdTaS9hE4p9K4bLdn/LapA7kFk8ZHxYnYc7uG1Yg
BfId0Gkzr6mUffvsOmcyK38V3pCCj0ZT6t4orjKXMzIcjuyFDTdF8UACCidi1P7A
GsucjsBPEa7NK3aBwSWxeIgZkBqAb1hA3Njd+YcFBWjB1aO60jrqT59KEFdc9aAO
uymNPZ/jj6P55DQ3bQN35sgzSD4dz3uT+73bI4MVdor39P2tRVX7ONMaLD7Ewcmu
QTVq3wQ1MuXDFvE90l2dHODBqwP3tbtWXHlIX8vcQjpHggs4XTGVYpJji0eUQzhs
pYQTJjD5C7p6pbMy2ckTOk4MNKeXvCjAeM7t7RpCp7a5P44HjW2kxkrZ17rgLmi1
/PT06xrMJRHWAQnzwkbnHa+AXCO2/iM8LQrHYez447ctlzUYuiX6fd3sFSO5VESF
cGbAcPAC7Dtu6TeQxEh5Gw5/zoG6Ej9ERD8l5cO5EXUGr6zjQ/1vugSYIBlRULRx
UTgL/ccw883riaaKI8EgcSVAQbol2gsXYdAvnWDhVdB7fM6TJIEXunu1ab66o6v/
F07bl7vZ/TW46M7gzYLVdY205Wg+61IXQHW3E8G+pbByK6QJIyu1UnhRczLCVL70
BoC9dI4kIRwifnyJkNQxz3RrVnm0Ox7Rihx7rojhEnRj+CKvAnq/+exIV0hMGs2/
di8mSZSbc489nr45vk6LLks2xJQ9WNBeAjHNFnA6n3wO1Wey94KGbWoQhjIPI6Zy
lvu9VZXXySHzIqcyodnPTC5S4ghIJaBmGWezMOAdHw9HLJVv2wRldbCkZyq95O81
a5rUreJwdzXwgKqkQZ4sgb2p0Sf5DEb4styQqIoUbmNoxQdfvjXe4n2y0TLjFofQ
Iuz5vKoQMxQzZmqu1/BvDxpSMzQf5rTFWW5uNZB1N4J35jhMxBuxQiCO7M+0iwh1
XhkWimi7OXSoaCrXCpMcyhfl9Z6Pg+lNpTstZhGCBqgh5sAcSfETrDIQGcy9Gxu3
GzuWpelwK2EFbWiK7GTCU/66pwYnfIKespnPbcsf9q/MCpYWCchIokWhD2MguQZG
93AJiryzQfZzYz64fMScaKuzzSQx5NA0bi4+lFmUr3MT8N9aEbDt5RdZxfxmYEj1
qYaX73GdCR02H0HPcj4ET6Y/Je70RllMsWrgHhrjrAEHMFj+gzc7KLdJCfxzBxP7
wNIgL84Tn7TRNZudnXYOYSF2+bVTM4rckblgikx9M/F2xjBtQPoWf7LPm6WTQq34
Ct1v2GAhNDvXfyaLCgjAAkxZeaN00COVpcBk05//LlAUJIMybysK24LLhzF2ZdZU
Yp6u6KKqnONfqw1NkP1SQE4iQpHdbdRsuTqT6+NSHGcGYjP79Asggpmb6zpsV7VV
2Uopy9ObqBpWyWSDQ+hjMXyKK8LgryE4vCsJflI/Pc835m/KyF8et5J2vXles7Ji
C+uETGzUBrxqwOXkK5F2OOTZxAOdi2RER7Lx6eaKEnqX10IDH4Ao6/Teu3IJV50w
p18ui1yJDANAYnUKjW6DixowsqtbUg6tREnRqOEXAnZ++CtevErEnFMW7Tsz28//
uBkR4EM9+xy7Sh1Fs08t/kUTvESE423yJNkAnhzfncLTMBy1o3xmshxv7fj4bfOE
WsOCsYRxK8TgKXXgFy8VBXdsskPicfWNli77JadnJuNql/Lj5Wn6NwUBaLC6eyb7
SoSjbsdNuFPxJCW+Ewud+oMdoEH/qZoDMWWDlsgI41GTyw769ei58m3/4T0CR9DG
kYy7lMKi8A5Q//apyHIfvtde3aF/WjT6FqzaB6HS67skPik8uAnFGW0D3jK0F2er
53OSaBGgXcbXM9wmLDeN/Po/C08XjJq+15SVntUnO8H73nIV9CuLX8KRnhJpuUNY
SL5wLaHTjdt5INI6AFLKN+RHMh23plyX7okxsP0uxommRSsu/D948EU9cAYtUnwD
v+ayQtLK49LX4V6qUt4eyopgpYqeXyZdCz3aUKsPp25VeFTJWXBebaswOIEgB4Et
ui1fZEYDgYQnsbL34ICOQqK5eXBBEbw2LTMErSrfkXCpR8YnbECWfTtNvdv99dQz
65SJB6eIqRCjavtvVg+H7wpoq6mqxZiY0PQw9igPl/UWfhN2U2cTJAytU/DpYsbA
O2hylsMs/STy4UD4luO20MxZT3NXPKtM7xR2OVczG8VyTpVLMvCU7Om+9p/1kzN4
zZK9BICt0Ht78XHykBXigqyfkHKhQlvt8102IRwt7RmeS76s6SxTo1UscSopJMsq
YXv6aU7X3OV32BvHpfkGNcBOetbOKIS+6QpwLxtF5Ujx98H+1CkX8CJQGF041rDY
AWTPv/yKlmRcyhWPqmJOCukdPWKfE1aPxo5uqHqwa+zq1JgnIRq41DQafuvacJcR
PshTZ7d05KTg57V4t6JYuaCPMRJ3XmDyOKSdU1zZkcNoUJzi6WmUJjYnoNvgKQlA
Xpda3iU3MiCtDL4T/Cn4X0+vI+YrtfCTY76EFjun9+5sJqN5DWXOdmKSKifa1AeQ
`protect end_protected