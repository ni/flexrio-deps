`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Jm2uGAVYfY7w9Y5qKstopObZuZAEY3b/Io3MSEcWLhjjnKulVhCBBYAEQrAzzGsT
vMbffkdZgjdXQUg8jOLJXSHZ0Dgbnob2vlppjZs3bgyHCF7MoJ35E+LOsaLimUA7
hlqStcK49hR1hdeBPr/OwfT3UeVrRtQyq0eJXQ1UksinX1G9Pz3/CmcGfTZ/C72x
p9icpt0bkY4/1I4GBvNCsA6FFKH947JqH27OPACiQQRW/K7JToQn+1uhWr3LA1od
lbVrWu8PdZi7zW9gK3jiW5GaPjwbYQGqeGFs3bTKBILjb7sYHxfxw7eDLVMAIu5D
W+OTIN4JiHiE1gCnNEvkSQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="pm+c2fYA/4JT1uhlJGVUubML8hZi8lME4xPobg/m8uM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
nBaXksR//iZ9fraC7WMJWWSrjqRXHxmM1Y0+KKN3b10NElDzVNMlR76DLrcnamFd
2n7uzsxWqhhJR5LBl98SXO3Y90J6BMbw+OBG/MFM/zUulxh2Si5YK5G9GCrG9gvZ
5JomxuZFDu9CzlWGTuRUt6FsE4Lr6sOL1P+hraQDpMk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="M8TXDiNa0BVMX1P60yIvW2WA9jKGGy8GtbuPknDnC9I="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2688 )
`protect data_block
/5TNZvs8Nu0G+mfp7M8H+iVAGG3Mh5DYZ0Gn3rRNhV8b5CcJKgjQajrRoGl/gSxp
rBAhtT8Vd5eelHgtvBjpvFBA/EBUrRH6CG6pqRt9r2qUDt4UernbZbxC3BC14KYF
06z4ZbN/T2BUc4DieG4tzFrJ+TRVLXdsshxDhLk4E7A+Qs2gRK58p5cSyeWiq6YH
VJASleKr7StSXEz/CNwvVJSd2/bBWqV0lqxB2iCcgkwK+Ovu2rLWkHGfhcEcRNLc
KGrhYFQQaPQqXeugAPGVHrjp9fBIaTQfK3BzanDPVdPUCvqPpAnWgxdJ5X2aOnj6
N6bSOdPWqMA2RzvrRJIR4JWsr37igzAjPuRPvFwnfavNjbevkAF5GbEiXCi7LnVh
uTftPgCfl7Qqy5LBqNd5ZN8q8obTFVL52uOPxCrPuy2XBYlH/k2hNrMoTTYPJn/5
4biDXlKUmo9vum1aHbyz8a7y0Z40cSFaK65vV0msu8U9914d6MPsfRtecuGw3EDa
SQ98AdhRfZXzh0iTNQBP6Dy8W9Ry90asTWIHnU1zeWT/O+2Sr2cXYczjvNB1DNKa
t9c0lB7WrFDZEpe8EpXTJ67v2yesyhfsVB8kMxNOPyhZdCBsZlmm9iEDpANPkOrO
4+Id9QasO16h/U5hyifZz45E/3Rxck8fjzfMagh6EnkQz1CCUtkm/kHGRhfYtTIl
vy9tv+ONE46WK80WA7rQfjfrEFZm64m5yqESgebfjBWm9TUVv7kykft0aOsKnPhW
24BYO+Eai+40/WsGEwClSsMIDnT46c8r9Et/g93l51YYeEpTyGIpaCPnq7AqpOlB
5KESmjoVdg8F1g+iHW7pBwzDpYn4EzuG3BTkmhRKJ9Jh96fboHzRf0Ap5/Qv0kAw
hlL6Jm/s7u5iU6wMcF63ExnIhrr1jfv/nm7eUiJgXa/YcHtxsE8ynQjnAYriOjOr
rbIF9l4yNSUN2/wnHQpq7s3Nlp2IgyBxOxdyQelvA3KRwNuDZbv4UoxGtFK3OTPR
3BpTHIDo7QlNXWX+GfIUHgoZL8A0rq+kSWrv/OXTk8R4+Vmn5ayGkE5UAVxZHdkF
ZQFdNejkq0N5jaj+Msje3he/NUZmHqQrDoedhWYmyKxUAVI/4LSKMRjx+VEY+/Dc
cvImzhnwbkS2Rx3NyenAX4tBd08IiIGDg1quHcEiFwR7DvwL8oq9CodvMOft40ZU
Is190ZIVS89YHFg+FbxWVl7rXzvu7HyqQQV2T6T+fT96C1gqUEspqYQNsrTbdhqf
0ouj9XICZUELaCdsei+BGVe3zdHrTGOKqGHGA9GzzYPExahnrHxb3kB4bqjAiNyz
mDerHM8h+u/xjklJT1QvmugCSkBx0CBFbv8lk0E4bAemBINh0GuVV6JRLv/VoPfu
n2qAswSdWo7k5tUG7uWD40PQAoyfckFhxt1mImbqRxHj2qcocugIgpktfEScxsE3
DyoQzDoK+xJQ28J44whVNRNNgaErpBQPpN3op6gvc4D9UKSqnafadOT3vGO9YHF3
ZYRxz9+4E04/hvKOCqPazZEKJruBm2/G0ih9Y4BZx+msakJJR5TBifGaZ7XFwaqE
ZPSnSTLWhISOr88HpTR5mLXv/K7sXWGlE639MX8ooUxCIPIAK35M5jZ44gxBmjsY
LdcYnJiMZSx398/TasH/6jRkAmABJHlSGvJrwS22SVyCD8VDZDFOVsBa284lhWYX
DBk7wKEfCaZcYfpLRLl2ZwS8mDRNTW7zj8ksw6CqhmFGBHCeGpaDeDDLi+v90w8g
GiJOumqVqnLb2SXaLd5H2je5bm9SlxGbArrbPaMizU7qHWdNxQKeLg6kjqZog9aM
xiJexikvMLwT4l2p5YqVdWRnrEu1LaALz5amb/vDnw6ihK7uR2rQQ9C1rhXPS0sq
DlvvcVLrQ4e9EumkOHrcOD27oekt1bBDO0kpPQXo2Ldlj15Hci711jEnb+zyiZbi
n4YT/tI5lFy7bG5XDj97yaCWacdnRzeVMq163td11wQrv+bjuRVWdwPCKziPUXDv
nn8wuybqOifjKP09a5pVvUFrCJFrjX3tlWQKRYo6DpaJZ+ab+QJ15nIdVhigOkaH
wNnzN3OwxKVtDKDSqO8lWPzGGVy9VlnPxLxvIPLZmfIQFgZ+cG6NCAdQhCsspQ+N
pkEXs5bs7/3GfD5GqaSE30wByknrZI1hKvU23XMhaHlDqViDbfRrXTgajmcFuPtg
ys/iv73EGtxJ+Yc4Nl6wBNln6EeOdumAtQWI6yfk7uiPDOjrpXEzY4SyvNUoIQ0U
th1eZFpT3ouzWJ7KSLcXmtZfJxbIOPMq2s+Ut/arbTeOoogQnvGQf/ls3AIZch0z
glnTYeH8gikQG/DXtIS8MRoTcNOS5J814pOxEzY+UI4VGYNEd1yHJoPxpfJcCio4
rXSty9GbXeCbgGema3v/pmb+B/d+vkntwxk0g3Wqcl5R1tXQiNCvHu9oTpdnYLkt
rbayXIwWfOrOcUVBmjVVREWfx495/welX2pyPH5i+NbApPwhCqbKDj6OWe8+897m
OYUj90JfZvIeotgvvFw4Tupp8p3QiilABRXdJqruy91C+aEX6qNWPbLViIdUW4Mi
T/+Z8dk/TzpTBgYeLfla+Vlbdec6P/XGGsLo9nSvp8LY+ZWTXZLU2xafnPEdWybt
Qa0zb/Iw8byvfvB4PvVRBtprleIGwKvtxwM/3ijZulBgWeh8grk5wWjQHEdBBTbv
aP1X6p7t2A0ag+QhcIC/kjC6d2OCNVBwx203yfSiNhIPIsbayHbyuyFD8jjdigcq
qZHIxmQC194Zhd1+mpO2gvTG3atot+IYjpVGqRzdFIcZFo43LDt8C36KcBsPIjn/
wlr0eru6V1Fc+pk6xW7SSt9rOIwOS76OtMEZ1P9xRlbipcP63mm5cTcm2qcMv+xT
km/yXimy9NjNGSx2LTAModVlK7VLdH0XdzYrM2O37JUtgZa7Nq88y5RFhi5OGHED
JwuIa46Rot1xgSV58RPG+mAHPkDiTzlwhIcCO5hMbBSkAO3zhxR9PJaS93MUHc72
HYp6ytFmiW0Vndr/jAY8+tNuB0PJ/LHRk/67BjCr4UchoowfywpdYbCkmpwJePw4
A11Tv+JhfShtwABIxCTwqZ8Xt7uwL138aN5688DvYP77cvKrnMKNFIQEgyZ2Jh2a
TG6YfsvRepIFYmxFAccRTh4s7tuluo80cdk0zFrh3b4bVfkofkxqvuHGuCKlojl8
Zs9LEoNFJUIWYVAWW0gnFiRH+9mn8ylyDuIRmN9uspNJNZgLv0fmrVe6nbGqqHTB
qGkQSTn2e7TctcC3W43YcXOpp4XJX8pQYqG7ixcH77NHX32CCAusvj6XO/XIm7Jk
UpdMliktA7qGcWulnwzcezdAh+AJ7LRtwzD7mz21KsTN1vpQt5sh3FcqP1kwQq22
kKbK1+O5z2Ju3YlKPna5kB4jKI9GEg8NZytmf0lfayz2FkyWf5Ndm2fY9Y63xgCs
zcqLsAE6vLcaZyD3SUhL4HOJvwZwwYG4GT7J8jp9FHGeiACFXBVVPDFerFfEOWRd
`protect end_protected