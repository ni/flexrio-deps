`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
DBGZtUPdvgnvgIFp6VMrQVvSQ2nt8W0r66xniSl0YKdCfF3KxvD+8aFw2qn5DITU
tLXM/M5Q7R2JYK9N+ruOeu7a5FpquACR+SGTt+/Gn21PDKoKioWLVzW/by9Xgql5
Np4eGMKik03RdCJE9Xa1YRu0HmbvfU1YF5cbJF7uUYO5e6DSmjFyNjVSIOQIAsuw
WR+HvI4xIRJgmLY/DX/tNt1QsEZAGWIy6CWIbANhohYk2p1jK6B/UFxDNpqJjxcL
tdxwDzNutdT/TMyGCF58a6RZqTPpxtjBFLS8JeycBp0oyVHIxDel6sEsAwoKuMtc
Pe9AQby7AsJnD7ruyIoHI4pYKJINCgjLjSFKawbaZJTNwU7HxYtM/2NRqOHn9Etd
C4MAnrtlAZUTQG6A9vUg0zNIZZeNqYMnGXTnmiE0EhOz/sMfpn63G9adfJpEm4Hv
w5yf+9/on+C44vt1Y62zFLHvmeEAzr8pCdLvFsH6rVnqqyDjWR2idWXmizxGzcaa
Mg/Df3C3vj7YdiBOgqL0U1rrfAHcHIAASDc0LKJ84L5Kp8gkeUU4Gghw6x5y7kzT
56I//3+jYT28gkcYVy0cwc+FYv0jRSUsK9mM14kTLJT1UhLafoPaZJy754pjGtHo
rNV1zS4J2Wq09q8E21UOSIxkVsT1AaIr+g9K+zbTz55ixTN75EGEULAVWJMecUdN
uNdrJhNON8gjGxdthMli72YSnbB+TsCY98eBlWG2PRVVO+pganK2bhMLifdAxlAq
GGRn4yNpvZ/0JnB7IUXsG0E18PJNQqsrC1zrVDTmLzJghK8dulotOsMNFBrhu1jB
2XGHqOnsVpj6aTN90thVPDQPQOuUXuleagylPmJtNVlYZZUwm2OS8EEWwiMj3pA5
8YGFLq+6QoiudNGrSfQmBZRSV+GlUalF0pIm5yg2rQ1SWHHDLsDSdvVZdLyIqPW+
wqFL2FZ7AG9zZJ3EkdZb1Bhs/jld1n8t4H1AJ0a+IsjL9EJd3MXpxXhlKAGc3RIQ
yvCa1STne76YUtkwzK+A6c5xHnuzthZGDsO/JQqiG2gb84JvN6wC/FtEFrOsFKIz
xJ1QRrJ9TzPPZ4znc0/fUggSRaGB91X+AnWwPC+IS17+ZLJfjNQ+mgx54InUkUIG
w241hgO0hVG0Su9+iGqijrVhcJ9LKeVunBS+HmWuNW/nqmrpkQ13lzLcIyF2UqyK
xH60dn2XizKYtH+1ZhpNwLExagH06FyA3+nh3jo9n5b9fROMZ2mWpLzWk917ABrz
uQUXbUdn7vFWV77lN9BtPhstPKpjIaQDqBLJWYx3zKlX4/sgUQk49vZ0wKWO3Cg7
I4wtfj5nAZdF3pK1Cpv81/ScpjyA6WFZOMUWpACrKoVAqb3EzN3ZXMtsq4GgAyya
Dz/K2job03J34Bh6e+nBasrGmiFLuZSP2/itp5QB13QER1EUic2ltymx1Hntjyy2
kY4fmco8H1w9gcC126OO/Nc7puzxWnuJaI638z+/25U/+K1Fv2WsGaV2Yd1kyUyf
Bj14ze5OzMeNPU5wOnD5NGTtDFMRVQ1uNh3yxvR8qJ2Ejw7Es7+aQY1l5TBIC8Qt
0Hj+dlpe62ipzF5b4sTSr9nm9Hh2+7gFyfaHIVxFE1m2+RBCLIFEyHk1NzFjBftW
3/5GLP8IhrMd5raTTDDpWP0stuxbT3sjHfE9kOJ7XYwVuEbypj+gx10LOPQTlIdX
oUSHAAK8ZuGlPxtSoMa1wRuxiHDUaQ7d1zVNtvTLF/M4/ELBm1xvqoGISFZVUZ1H
Aa0XnJ1+XyHfxsumtPGrLe6p+BBXiDk4IrtBjOXEBEpdllg8Io8bpb9p4B2JsvNR
yl7ltfwZakrAY/5oXGQNfYcjoNoYPv/YEsgCMm8cDh0VGhQ0uLvDNaoQqcvratOD
8v6v1CMSJJJ+LM/AT7GHam7Fj5oGc3UvbS6DEewp4vdKtw+Wb4k04GgsNECSNyqD
e69P4OguX3VYfWVYzFac7VrpbJ1DMZV8tbivEv+gVZWFqDBoCRsJYlHI52XMc9zn
+467zITm6vB8bTXJsziDy0aU7bvGp1BDFJYQaB/3FOymFuP+4erMkuRjzTkOItd2
WZUQn3TRvnk7lABuD0T21pp3y4luZ1pKceKeGbSKXqKuCCXd6Oh7suNliFQRFY51
9hKOOd+movphiP6A0NxXEN7LsVF82jAe2imWC4GtDOlVhl1i3iT2H+HczR0beI5Q
27ujecNWcqZmQQ7ZT9GbzW9n2dRMV89HRuHZoATAQmgwBkUhrKPZ386ANai0Srou
iFmRdK8AOZBDPKrGB7Z7Bnyp5f9qSsQFd2lzV6zUwK7gVMIaDIbWIF5ZD/3Nd6QL
1lhwmw24LF++7d5iqvMsyq7P6pA1xVi6B8xhU1oAkqA/qt8fadlg2KHJkkqd16Y6
4AqCI+4rHLrWY6ysh97hAW8cndGRKtxw6jmaSkNfC1Bb1XpQ9yWeqaUw/r3yr197
et0pzsGTDf1QVif/f2x/S9qCrcsPmasHBFTUSrJ88dQvVwDYzWWX937k17wzAQ24
IQ4u+SWxsbHJpGzUNsGkZSfcJhmXdSRO08j+flgl7WTRWzbtGJXmm7JvKQ9kFYs7
COS9raKAXO2LdxyYqS2qVbtyAElVVz0XZsy2/WO9JFoIEvDqhtLRHBLXcrypELjJ
4T7ZsvXzAfwSzGVb9rDoJIV/t/gwVBLbMYz90n7MbdkFPykTKDK2U9oexSkVcxJN
CvxU/CNYzGEBx8i+kkahzvF34ETf6XJMHNfikHIHhgqF/U5WY4+Gb4CWBVPfmMhY
yweL999HzR0A2OSYsRwANLMp5w1j0pPerTF0m1Z/l3rEW1CZzRTpTvx2Xn7KXNhu
A3WHiqOpRM+vpYnNQoK2oX9N7XNXUPHuUSvSuO5KVPS24X5EATlhvRFdcMVLz2qe
osTrzuZviXWKQZCGUSPREqR1M5jy9GNlAzYxdc2gdQcHCvV5AnXp7Q0h1y0o8I/8
uaUNKnoLIINqBkBqlX/LklfniEVX06FoQxQDRIxH39kGoXOTho4IqraUloFt7ttC
A+NR7pWDJHqzNPMPtcbGHUsB78+5EaLBYv1ooYQLFOAekMyQtl4ZdTJv0BT6x0g7
ceOShWb15vOMfrPJ57nxHSl3mX2nGoze5BNiC3bM2PpuN7jrmmk87GbcrIYWhd+k
d0EMDS/WQZUZdECkcvkJSGuCLBbW1LsWXny1fGSWbRgF3uCtfZaXyBRdGiOj9zkE
dr99kjMbZbWw2a8rKuunWajcUb4naUtKxiYqeVS4sAB5g5Gn/P7yw4KlACG1HUsC
mNbKr/4Yl56Gz3CDU7U1qp8bUK6de41xZJk1T9F/gyJf8WvkN301f1wJOSiGimFo
p50eT63ZU+oH5sbvX73BqNnfluI683mT/kyYhFVk0ArXOHoxOh7c1V/YQpTzkaxE
CIuhE+MVevCSyavVll5SRr39grlf8Gdf7e3TI7huXB82xKfDxYcNImnOpQuQ/tQF
H3mgEYmw+Jqub3Luol9N2kjj2jVPn77WPZeuAxJpKM1ni8CzODLvswVLFiqRIw1y
S2/74y0p9Ek+jaDATtePFRr7ql/IZrsDsmnqiocAvjvJC5SgrGD+0iR3gxyApEQj
gL031+E4bAdR2Cu6V1YPKvrmnMJQ3qKHZ8eJig8P07JanHVWhk/zkUD7D0JN3RPE
LymDIRJgVFps+T51aQUx8cmG66X40hrnS3hKR2dsdy9/hfN++p3nGRIocE1/yG4I
4oOLlSmns9SDq2ZlT5eL/qQxFmGo6jzu/ehfMj9vCkp54GFmlStmdR9PkgUIc2DL
+2j/dPVfzvaxb0/fymM7PsEnN+ogs82+q1Uz/n7DS5fW30UfUDo97I5ULN6WLcl6
m6KkNUZyqS+d1S5NuiRLlC6ZIBehRvF4fHmWKVmt1VWreknuOr2IMxHoOJNGMIuv
yiSxB6iWXpFs47JU1r2O6ipij2dLqjQJCCT3//P8xTw+uP/aLQPnNsB2GQdEa7Jh
7JPY4H1wCobYD7wOnIM/eZZ91Csq9/1iG52lGG6tN+qYO+fZAVsGrqQw0HEPKK+I
UISW+lypsjAa/Je2HQPhwYM+YhY426rpXd9hdSXhR8NMqLSZw7JuNy0bcM8ggxuU
xYEUSvm33A+nfaa7v9G0mrYTxU9XLBEYUA6/HNGwpXMPq9tw+nPL4Q61/0oCK9yj
NtdBfLGuUNXyrjPGXUl/RHf112aC4TX5HXPebzvUMI20X59Og7NGk/tOsQMROXdS
bC0Q82BWjIT4g6iT3SREz2LLNvljqyxjCgrVorNpC382U81XlYMT5txBu2WxxE4I
8rttux+/0vDzGYyIkwHk0aSCllpISWon4V034VbeRbHd0UBqMPCH71q3YvKkLJkL
h8iBtFdspIX1CEvOqxyQ/UGzLcgO1ZiCovHYa4ypSvI9eKUd2QKqNfzWCZYONUsg
nRwLOUOWouU6e7o50/WxxifdKPIzA913AFDlrUg6xzuU3B3CLwVjCt45zN4EMY3D
cxKMZtzNkyw334Kt25AkDyK60q3ITNbbld3+ASk6z8rtzrF4lq2k2GsBYs+Y5wZJ
es4ltiy6vMhBMMNdLQzHX7I1ZXkkKPgmp+8o2G4N0LZy/yw6j2IzSrtIMG+zn47Z
oJtfoNrtlLvWQoNwxgDlCWYm3hElgZMG5iT8UJHwA4wgtPx/K/5APNGLDDBJyUsX
U0AQIFX823UmGDJsfaEcjmUmcaLO+dpU1TJqkpDg/LIB2tQX9JCK1aeXtIEg/28K
NuyObfSJztosid52T6tLPXVEt27aHQ3FtknnG4fQ6Tu87iWuenQo77o5aB9vPx8u
VY5I+SP6lpwGepFFcGJhFpC5XlG9SIa63dFDqn1hPA2ME35GXXuthOycRrRqHIEO
MhaJ90xAM8YR+/0zBDANroc1zl0Ce/+yDnhUVICp/RMLqg7sfIgaKS6SRlZGAzt1
qxySX/T+QXel7Bbrl/CIibviBKeoLlsnhCNIchqJooqfk5i3QWGacRir7sibLilJ
gORN9Cc4QYnu7cVYKENcjOH7QJMDO4Q57OeZ+wOs/rhOBI3JKJbPi2VaHymI/DTb
cNxs8P4wNTNh/LldZg5cHFwpSKnOXHGL8TB9WzGsxP35OODVBmqRhQmrg1mk37rx
LbNIDRgzehVBhH0b3PafHCRJk6lUH53B701TDALGTH58kmR2VNZJzquXadbwF6hS
fUTmoVFSxax0/Z9bKcfZ1jYvFgZEt716LfAdbdBDn/6lv2X3rCLfMNqaIBVItNkx
8bWvdjdIogFtXkK54ADx45P/8KInKf7DmygAGhUgw4dZ6M5E3uosw3uqypJEeK8d
jGhPBKNZxEwGH3JCfjzLmWKpa4Jdhs7ww4SQjz1L1niUFHqYkA0MvegXqfn4EF5i
X6/MJshTjP86Hx3c070PtlpMFb2coQQTW8aEaz/obQj9JY09oRB+MQyUcyw/rnvS
N0qBrUCPKNqB8E2TVepVlKkHDjqqs9CNclzBOLKM4o9fDVDNR8i3oBWOVjusUIn9
AKadxqoYitWp7OgBntLMsj+Ab2jHExFXRzovusPHt6Pplhh2gnNzdwrXrEwHnKqq
+fprXcxhOaFMulBNNHDHI1/tNqGLv93F5Am3mHjwadUTYXPni2LWeB2YkfQ6wNK0
U2cH32cpJ/Cl4C+hMNgFQn8bDOvCv/yBDiJxoIFPbRz0Y6yy+HyCtAvFQ2SPzfoM
jKsf6f/GYOWk8G1pq+X2aFPPaFXtAyHEp48NW/EHCfWy2MHuAgkiMgsjLtheoLLH
DEL8gwBkC8TIrJ8d11LCyB7K6i1Ujy2CA9gcsBlWYmXqrHVG0UGnOakNb2dlRcl2
wKgpIJ+nPu+NKiHbtKV3WXFu9w66rtpcAqrSkJ+3A1lHYHvB0HVgx9oFbRoBd9rn
JLKcySGu52uO+/98HCSrRK09HrV9GDzYw97O0qCeYWPFmoHnFcXYJoMgpxiRhhNv
AOnhek+wfww2JHiqNN0zE0NfQNFbrQtDcLD+UaohC/pyDN1/ZBnRdnu0tHnL9HUN
5jbch02JKnXRnxgol7ew19K/RMfLjeoJ1jjJDWWS9FwiK1tnf2NPez1Zkb5qmkMF
7C/qJa8H0QSlvaoVMzf6FLVRv8uoAQGFM9vZYHhHXBMarMxuszZI2ZZYbmBUw2eJ
RPv5PzpOf+MQUmGhaq4j+xjAy4MxEcCTo8avh8EJUn9v8YlscIbLmhyq3Va6JFCb
hpBHGcuJwdp3YV9zZjLdCQ9PI6+2dkpgfQ98uRY4hgJnkeYqTG9zmlVNjxcvuVu2
b8e0daXgoolSOLWOmktMKemfaT7DQ+wxnyMfcdFIkV46wmf3TPVx+jFEg+yyslot
/b26jcuy/HouFo6LjmQyR29G09DJzkLpyIUi+/Ed6JMBxjZ/556CDOZ64kLYbT/j
IUHNesbhT1tb8VtonvfbL0F/qnvd60SoLa5NKgyx8zsNSXILjnq2ZR60YXUIr6IO
SUstXeceVi2ly5Buu31xatzC1NT7Vc+d4XZLrf3m+RySjfD1WjOAN0Y5E2gDmFDX
/+xouMYan2l3jbjYq8W2eFvCv72jJiaK76sY74WmifNMEn2en2NlkBGYoC/hqWZH
cuUteQHRLNc6fTdw3/6PQghNvmabLMunZU6CHWITfx/BO9U+WWwmpxQ18s6hXrUE
4AuOxdJg/UVXADccN4l42dQnyPNdmf7jtao5IUvTI2eeJtbPpzKHuq1pBU/rOEdW
LH5/dPrq+cTo62eCcIA4bZ9bTWyY5sqcIJCTWoEa3nZOMntgrLS86StTcri7KT23
wxa+R5UlUBIEeNLHkZoO2u61EOV9SirrTWc06l5C8sGX0OtIzga/CmnrbiAx5H1g
uYlFUM6eR+8PiCcZi5xVGNO51HbGtw9Z3S74fOskXh5s5m3bFVeYss/jCsodqinm
qoUDkAW1QXpHRMu6Sc12eip9NzwvYy89wsEq5Fg4v9ARx/D2QHDbXM3JY0xTQiGm
XXNkBMDqfQ5WCiaemyHfR73toilz9ldEXBVd0P8PkZDscIBvZ/HvlV2xSMNLOTs2
T1x05YE8+LtcpWK/gtx1J6g5xS9nmbdVxVgBOunpBuyBv0CADP5PwgTONxqQ3HXZ
0/80AyCkEpSFyqfKZs6zPmouEm1hA0C8KJfeBgirBqXaHh9aNjGn7KGNqEVB/xli
avzOqh1EvYJPJ634cxWHJ14gBUThWT5KyBcUjrzt6KV1W+ecPeXnEw4BMyglKGxU
V9eC311/DXvobjq56BsmCUv4OD7TikvOPo1XuYee98VOWBvNrG5ouE1HxKPgVQTu
7KJejKa2Sut6TuwZKkJyJu8j47V5B0CA3nDzNXjoYG/ZwOLkg5DzquKTXJJn8koE
dwSs9Pfxq5Auqd7AcK53B7ti0p6w3tC0/y+eR/uQox3RPACyL9Hbt09+rcw3eAsu
AB/DrsUJKDfDpIdIeQhu1+8P3G9ysoSAdUVsTnx6uILexNWiaRbbwv0JVaSvUHZD
gVB0f6vCEnTjMsL3X4bobzhyhONigjag6qLXuynm+dgDvp2iz0CKV2jlZW2AxBxm
/C746yOGBhkO7iyS6HzTgBGDbCjEY3XdeF3ERLua4d1leSQvDrCvasiBUgdGlJtD
yHD5BLFoNMEN3byYyFjsGlRUCpbbqR50LBrfwnx12fMhygRaNFuXhLARYbU4Za4q
SJzEJxKx1MPCMn+Zihu9DYVr4eCVy9emDxyh6qF4QmOgkn8aOWyburmMCQY58DVv
gj8qCxnq4S7twyQZQinFsmMJHVIkPM1K8ykFdvAvZFpL+Ocz6PlZudZgkebFcMDs
zUGuaHuNuIp+mhopCio12Mgd6ya15ws3qf0+12fweFnK4kQv3TTimO91iq1AocFY
oKU738VxP9Dt4VPT+65VznY0sKeI3xzFmrpQtNOQtU4ynQX/tINpkhDLiMBqqbDj
lkDMs/RTKkjrmfHB8XMVs24o7PwQvM/bFAZy0PYXOyFlu/MtepR2khGysAjg36ys
z3EjQrfUpW9FcJmjl9eQ8ab7xdXVXjQRFNa6yiZdQRpNuQZl0g0e007zRdIO3HGa
onKierxK+2u1DqvddjtTIm4Kh2XJIso3jbN3bb6NKaiXi3kXtR09QDtC/0Su+M1P
TP/WgbA4LOQnwmzF4+K/Nz2rP7ho/OoroZU3+5GXmGVHtnSoVT9ROMJk/ozyrRPh
TOHJTLRAIn4PuuXA13QlcxrV+DOtxQJKLSfET7QfCloJ3nZ+B7LSFjsySzqJ7iBo
0/ntJkr5p4wipheNywCOgdA5E9UqW3CFx7GTKvBA86gQGURF80k0SV1ITuCgj6Hr
j3K/vwKwtzxkSQZrVK4Cst5gGKqyD0F69iXtdy/UUgwvh7oy1kg8yD3xdtwwjE2g
iCQdQjBsRFi99oTnlVGHSxYtuBCjbRv81S59Wc+FRW5TwwQQoerSbkZTPssW7daP
K6tutBmtB6QCcPv4OA4/ygXANZcbreV6nk1vjIoisqjUbbZDC00ifrkQIjIB8M2x
dwYpwCRsDJdz19AYAku5D7nycL+vFHD7v0pfmmrpD/+6mZmFoawK5F19or48K9uo
F+gJBp+qSIRNISS+yitsIS/2CPomj9izVutvIHPWX0GNQNV+0jE1Odg3p7lOsZ2M
FGVitHIJKKPOe9iZ9RZFyLxCa1yhYjHy1YAF5DzaVEaAxwG48ZVmhV6dh8pYHLmt
uKMAwPp0jwqRdam3iz1MVnQrAM1ipi53NQiQ0UNcWHvjMutH0k/5Y2hQZOulCD6W
vT+Vv2RdOtROkr92TP/zYPGrCLfA6N6S8rlkGyOk3E5UqHZ1pvg0zKbYZfWx91yb
FoWMKCMT5eiwGHWg2uCBhqhfFg+5I6Snndtrvr6uJTv6GSjixz+D/ZOOPyAyW5WI
bAOCGpl4jEXz9YHR471D+0drQ65EAz3jxIRVWCwP9GO13XsKCZqMDNp3aJIIYpyT
n3VVO6O+KQFNUPnmAdBjVHZr1qHM9qrhDKja5oOPHLl0SB0ObsqyFV/iHbVLNdZX
adlm/aHBgAipVWX5OnXSm1Qf0mV+8x7+O+udnpyWQEsBwyg+OefxSiZlFz6+gqAW
dHMpbw8EXb6n9Wmc2YcJoJgXbRHNwfQeJp3s7W7vZapudrjQrOgCuv8iBx9EVdXs
YzdJEUamDACo9N6CAAXC0NR5dWiiDvSqKeDtFNSSbyYbskG3nH4dhotQIu91Zda8
yx9JVjCQ7CyzyRNvB4sX7Ken+c54Ki3qWIb8oD0kNGh3Ddqx0fm+aaQrAGBEJl26
abryoBYQq2D7PkFTUk21Vj380GvGX83khQeKVMSyaJlatppuTssMIYkSzsqnwXRh
wIA8pdPsyXTwFNckTEKxJJvLLZqO2r3jbBwgsmDGvwi+rOvWiuMOCawQwvEYGIh+
helkZYJvOWyqIf9ul1HAl5O0HT+G4pCqA9Mg0PlZi4TL8gmZ6VmIAenN1wiVLkkk
8VLLxILX4SrGjjxamy+YTLp4JA00BA7xhodgYrt9oBut/q8w6rS8PyIlnYqgaVbK
gUCgq3M9+8fLNMZsugj2bRUOXWoIvFxfdpo4euzCbB0SQhhQ9qfudAs79//aAVcE
xtfGOXhxdMdC2ts/pSZ/IwbPn4xtErCVj1/wsrOyMHElC9vExk+XASYuXLTOpZha
vyUnvchYYCcb8VX9AkZ+rMA+MGXMqKd687m88OjaC6fjsm9fpAnlmlOYhhwxh+pn
4PafSnsETOJIXRtPmUQOvIDjK8rnNU0D2zZpaxfLzzTTlrGZLBd4yzQ3h15hlWYw
3MrpZh6xo+FcRT5Tq7S/eCBAfmxK5PzX2e4FFECMeFqmJyoxm0RFHxXP7T9C+cS2
vz731HUsjAIVNIHdNLMSEerIyVcRDKWD1vjovzm0ZGr/aUE0BVbZiFPmcav8pVU/
B7IzcKzldx96W7nIWnNF44X3YGvJ5BGDNXXjRmxPxV9XanHshpl8TahW7xeORdjv
ZjwevL2XbhkveuY+3KLS5CaL7RRyObhZw6Ay3jEWbdeH9NFqlTmbnLAV/fz9S16R
vHSqbbVFPcWBlSFjtS8U9r/7rf7RvnTp3DYZMQ6U2WmqwabvZruAdTiDNbsGNU/h
bk6XXUZBTt6aPQBdbuKkXgNcOfoZY+7dpHxkkbao/GyEsBFxJImJeWTUX+PH+FuC
PD94JOdWvcOSLnlc55n0c8eHxHXRwUOT9HuP1/m95dXOu9qlGNt1roStxEdmlDwz
VQ28l7+mmy5mcO6ySOBe3pVGTsH5OF5gFFSZyP7LbAIL4rqAaJfsHbg16eMK11vN
yH2FOYlK59XGOl8MQuEyf+V/c5SJPIFcxMuW623ut/kAyyJrCW83N4BrxC/uXtIw
bnCQKqc3ABcpAg8dDFvnu4bw3/hnRqieKOLRvYaJSMwrnJOdombYMsZ3vCM6bbJ1
59/T4dOryBVxOnh9J1w7rhQKm/mQDFh9UAeiVq3ut0x5+8fSqI9eu0sRfdkRqiiD
p/n4QPr3Fnls32CHIORJb0IaKjDo/H52HEKTDFbL6HEjFCuE8RjO0Uig75yiesPP
AwDsIA1BQtF/CRHlmZr/dXvh3s/ylG7+losysnL5vbaEoKvenNSp25+5AvDpNjJu
4QY/R+3EhGgRqgDjbW8rYcQPH7C13SdvbW2Errbwgkv1TVIOJrpNFk3pO/fTGlsM
+cQFiz+SkkEKRR9awa52qwS9Qohaz7tTTHXD00w6QN30YxXN1azLfFQ4STwnXuix
aa5RkNrJPTyxMI7rzFhTZ0nXYBbXbIKp4H0g17VP3JSrLDK/qMcGjvxw2/Xb15L4
avX36Vo/W0uAe7kIuc+4bKJ2O3h+ZBFYZZB4TYkE7B8FXMbIcMylOXAkFWB5dyfo
pQ1vpn73WNVeagyHDB+bBjMxtZSB5mcymVWFbY1ID/xW7OUfUeIlfECY1UVewWLX
RxNpflb9yBDYxVAM7TOro/JzN+LkEAE9PtxVcshc0Xgd4xcCamh9owSzgd5NGo5y
v72zWaPzE2kfRhI6m2HE/3oixqlylkWp8c8K1mrT5EELrUKo9ltfIigs8CSiuTKB
qFTs4802JI33TffIX4DyiU7OhAogADDkmt6L0wUKW4mc9FSmrYIPjRLGZoWK/LBi
5Qfs5FfSE0ZfInJu9eXgpwrXYJhODgPYOkSM6Hd/UMd0sFRcwp+RCRvlbw6d0qa/
OkLineK5hA3GP2lTPCHqc9/kZw519BIIrY2H46wd+WRcMJcu2uqlg4X1rub2B1km
04VNrV5DVgobN5LESENe1ukl7tuMdFBX8rpQNYtcOMDk5jvbxaKRna4eoqWbGe1g
Fsmdmj/lsoFmmMEM0FJh9r+8VWN1NnxBwIqcCsvxdJWye2ty2rcqygi4wfirTax2
oihQ/udm+wsXxZwgWNIfnIh2aVUh6r1QrMWU1auwf06FvZa1Xlczhd9yUfX8vhDz
rGfHYj3O5cBfOMN5iN5RA0+ciwtkPZkcnXaokLOi3RnNC4r/vZlgdOiUZTAjuoub
8wzipfacmsI7aUCZqr081Vl9JLTomB6ipKxjGIEwCXDq+1caqh7zmctlRXgAgZcI
5yz7dzNNuWHv30GckuZ7Ozk/VNa4M6+q9sutmzd4Kb4vBfoSnE0Ob70+QGmc9Q0+
sEowaMoZ02IGCWTLQaMnerwdLRo+Fdv3xl8/hV3Nzi2ueE7E8fYS+9Dbmeiem1vU
FXROQhoVZF2bezTnk1eBib9gOYA1dy8koG1NYt3VzIJUAUXuMGUbEQZKnQxw1nhq
B4cfG0NRbyhgUnd7/h5XzjltNzKQaJAuUgkqdPqbAZbmW+ELtOhZsgvJPS5m5Bcg
VZFZxlpIhHqRvQOYEpC4wkfBuoCBZDgydyl/d6NvdwFnhVzos3LvgZ1LlW+S5X2r
eBE+IN/Fhasi9/rfn6ZZjaFJnYBlh7PPrkZbU3WgdJsmDNZrKtb6XKVg2eNPaExn
EycQH4iRfmbuOdb1Gc9o/wXwiSn1BNOPWPO0tn8GU0jao2tMevOcZLKg1GAyKfJW
eo90DPwKoQOEx50qPCUmyZoAy77cDbUyUGrQufjFvaMO2Xb/fl8ZF8rW5Ib1+xrS
144/aXhzLVEqwF+efJ1JQ6H8BLI8lnTL65ya7szoXbLTTblDdcHdkmE1bJEuJclT
ArmOW4RMD+zcXzWIUyBIx8+3Tl2nIATVNZQx4cMwlLZvourC8QJf9Zd3OrEn6ttP
6KpqkFfHT4yfwRoKbcaNmqIwwVVFdWvOCLiuNViztLtNP5iD/Z1Q9Dl1v2lc6xFG
umCU/fiFStX+nGlck4J7gJlW10wFtRn3EbttCltNXp19vfDwyWepk2q24YA2AV2R
YcifyRfG1rhZMqMFgtxKbHChK27SuPnka7TenazFqRAH4cGOdBOo9e5v+5PzcF8I
XpZYNVCVz3KpKdCndN9978Zbi2WhMdjS3HWa9wCU4oMwHbVbsOMHn9zN8zKsJ77r
dM14v7Rccatg57c5cMh6GXiVH8ETlEmzx27JD1vxCmEc1YxTRiJEROLeDcxcbBwR
XdVY/7CgqTL+19nyYQcK0CuZEo0KYYtn7+qB5g4pFuVQGQJN5Qjpi9EvK8EOm7s5
3AHr3Ev4M4SPVgkdkZyeRPfvG0nNeQ6D5PD075KAp2u39SkrlzG6s5DNa19f9L3Q
7RBVmKfD5gbUSF2HHq1KqY0opXZ1KuiP9DDKspAeQLsHcTqu+QhklR7JAapdvG4g
feMEiMEkmAnqfDzQ8LnixjR1MNjXZ4g+RhZLKKCNI0KFsP5NSr3ZKtOXyvauwTPt
aUg0Bro3ysIaxfdQOWSi3TWI6rMVCuxUeSWWMPpdu7QqnPCt3tc9YK/6F6gKAcT3
3F+BSgPMlxJYtlqPvZkAtpt5didZMrp+ICTgGJt13Ih8h+upVoOu5T4nbXGDwJ8N
eMwVtJOcd9DqXlj8GaIjWiWFA1nz8pF3QkxCz/FfbOg/v4kJJbd1y6A8EbgjFukX
IMuD9XJx/uSyEBta7cjbbrCGIse50pD/Hz2SMdHe4sMiDpQ3HSEUkwnKeQfrHYbR
Dgvji1rVlfvwKAx7vy1IYrV2opsn+MswZ4BdDsWbcKsc7uznpo15BAMp01owM5xd
hkXf11YGmg11GIAAtPISXOAJkj81g69JPuBAePovT5hfOn1OUDEUSQVlOpukr22R
/MFld6U12qdeUbCMWLBIBxWi6ehtVOmPuuvCE6GrKtEpTTq+3USJaxdKLQGJ5ypa
iKqqTvYj5kw7VIljfkY0VMd1SVlYiovQTVQoQqa3E3RVl9NtKnElpMMeXA0UAg+8
NojGOgxTgyjKKCskv/PBD4YU0QhmV43kAk/qbs+u22xVl1/B0U7TDAgZIGFIKBgB
JWKD43+IL/+9laI4uwF6YLHxkQKplHTyfTQqGhQOHvWXsP1wNCIWsyT6VpKAvhWR
j+kLiS9BGQD9sA4Mc3SCVm8xS+J1Cy+s5XlDC/NmHkLbKXQRd3/72ALBHE6T5/IC
RW3aPEYd/gE+XHr2V9GvMBnvi9f1VluJWdYshl66pcPWgrerR47tEiYHtp1W7784
YaresV0I8aaKqIizn3Y+3ZHnZfWS3XVOx+/4gI+zZtV3ywpw36q9QdaGlanE+47U
VenGymeMxGcovV9dDvnCbukjuCoXhiLOi7jG5VZk3WDKYLr1tUcteGFMDWMedUbQ
8OAGSh1Mpf3Sy7I6YIOOwtEDkwlaI+k4cqoW0z76PVCnlEQx9yRiAloj5sZWgxPl
iQfK3xdKbtXFgYpBTFPfPHAGQ/ImMvDHK43/jXVtwqDYZQ5/r0kBAvIWPwF1RkvP
Ek5iAkpOk95AZZ3nsYi6M5R739yYgTPCq9RMauUXFc34GbhB/nmq1/VXkh+4ggYG
UA5c04ZX/JQFcQxOAdxel/X/9rqSR7Ki3bt1QIPCsQLmw3u+C7pWeTZgHWC6ufAM
OnWBOiGatbOqMoNW0IqIQKAY+Dre4ErrHVIgPXtY0YwNQrth+VzIX+8sC0WT21oe
rta7mSDQABkdxlnC2r0yWDlaHfhtUDYy4qx5O5YTNtDqlNDEKBsWA/OiE+sknEQL
+PfGG7RTIA0tesgqYwHbBPFFbE6Ki54YN6SqMRSu4RCbyjygb34ttMVqRgxNhRH6
o+/NRrESqqImZe8Wee0zPrRU6OOtCZqkJXvVC+1Khapo8NS8GySiMDNF/QIIzjaE
gCJ4PTLGnljRemIeaXxvNKLrqgx0dacpxgl6szPX9X8F8c/LYFGHnWuiLE69HtwB
RmX0Fl8A65bH1D3uRCqKQ3dHtphM+emXmnQJVgTkdiq0vXN4gq+myCrAZpfwD/ii
y95wfhq5a2EKbeMzDuNTxUjQUIE5hJMnpIPZ4F/qjIGJZrndnkb840cKu8YUIPzI
dx9yvFmJrLzccn8FUZdCeMNktImVJrVg9MvvFBHP0b2BjIPqla0cswAhLWAq0QRF
BwqrQZgcaKcQHnnTWEGRy/vSjBqGknD2GRyKTHIeEvZYdOmsq1LunyYbs7U2oa0z
2oG+01th3aDidvEmfz+94Jo3ci3cCWGqlBzo/scaCGV70KHxgvLABcYTwWs4d+Ls
MtMy0WCJzrJS33MrwxgH9VS5Gco2HMTwjBRfQjOvKCBgfGQ84WGWpS2aeltWj+CP
jj6ViXLweE0m3WH0+KX1jqIRTTCIC9UvgHkugDBVXB2gGaPoHT6xzZ4LXnF4rJdR
mtuDzy6T6d4j3xJcMfMBjd+FCFRlzKQDZFLOXIG4YWst0j5Dxj9FUQt8A4+cg7P9
bYCFwjgqYUy7lkxEKhHHLi+9+TXrOsowl4BeP/ngNxUSvmuBQ54ligZj8wdv8FGG
C2irjsRqWe60/UvOlPEeyg1m3IYPFs1FgfZJo7kIATa+yLGtLdSdfP+uJ3vY6GFc
viysVhBUzU5d7P0T31UJ1/IgCRjXhENBq/BkO4LXjz03kFMHUMj2+QEMjTOpZly3
efrW1ASFfZlEvMidaMk+WL9MsKASOhgRdhANQZySevIcAOi78++0qQFBFNFmNm6V
Nl8Yv1tye0gQWLgx7w5X7vlsDGxT7DJ0FzhSJPnKpLuRTFBFwEfJHIpVgpVj5xlG
zhSmmHGfzpXnMr4RCZCTga9VFj6dF8qhUSPWBfNIqWiFJ3Y3NEUK/QmDTrbVBtf4
aUw9mg52AI8py5kKlVErqH5KsYUiIphgtj1QjVPIX1PpKa2uNPjHSxO7NsuR9oPo
mACkuSQ99TvPAZ954lvoWP3786+2LgU6Wa01lybLbhbhpqAK1yg9K/zjvrSJC7a1
C3f5tkj0LVbqS6AyfSETOjIpC9yyJPuJot/ogBRezser+DJI5mzxjOXgDEaek+qn
h99Cx+99IGO2UWZB6YBYXAi3Myl7P+D8K3UjyLcPOsWulyoissHrBqrPAAOEfhme
Id/ZYbab87+TpHYW4VQWkNdMtxOpiw+Eu9EVsPxO8ClWGDtmj2e1rMxaMdh5D7vf
hQ4Rnrhp/SknDIzefgKiRSH1u6cdhDogEIXnZCnn2hnBYEAKQWGy9yIA2vlUnhBP
kVfDjOWj4Hc1COuqVD2H9oOc80thyXYs2LCAFcrOKhI7t11hbOKEZZ8Qm8FZVSMH
3lHShOnCB9Ck6OyDkaGNhSSvqYfCFBe6gBdQHHnZ0AMXg9FZVaOsUxuOF/E6NbNc
rN8si5SsajRr9ghH1Qc5ES2mZatv+53jUw1abP3UdaWTWqJ1y1oNN5wf4NPkdovo
WHvz9tWaRP2cVOnGWODefpNTKUBQhLP/XUyuRfVKD1aC7StnZ3hXKmlRYUf6VGZB
I/LDzVUEvAYtj7aa+TWG/JQQPdhawCwjfA00QiETpSaZQJukB/U5P/i9K1eqNF7y
/QBMn2jPrXDLAJAV+zNd+x4RQBDpUFYaeK9FMTprU3C/TRO+GN+3XGYl9moPhBej
QRT/AK9oz5mH5jZxHlUwOkwiLU6lxgXOBD+CxX5rDoiMyNLm6U0B9p/GWW4o31mP
/rqgfbiu7iNkgE7SKDdQOIm59+cEYQnJKb8hDWBDckvWqEyRd5lO9YLr8I4VBhq4
/8ynZmnBjx1mz4kCgDv5N2M/ru2EQQ1ttZk94SPpBmGZaehOJqxx3cJOaH+5BRw6
b20rn7b+s0livAjDGR8i3tRQwQZ+swCRjjcaESo5gCx9bLIv0czE57l8/7EPBtTu
kQHAt4iDBr3M7VDFUfGmEPPVT5wh99DNSRoObGqXNyc41Fpr05C1/9v6DaxzSCrb
2CMrlKcSp//MK/JFmvKZ+MFRWnoVggQR/0lAdfW3cuWHc0E0b/bxtralXdfWr/lw
oDWoWSCXwxieSONkLxZS1wC1n4hFuQdlzmCLjJ0rmO3BcFDHjCZ+oo01CvxIkmav
U4ShaKnQ4sW5Y9W0gY7hs56GrmYgIAw63a/n53h3rsxiz2U8p3EaoEFtcbISdIfY
8n8BVmzi0RZ/i60ToD9o7q6D/yQ5jSvFHB8dFGCq9UNnhcI2I6RQq4JvDRrZgCcl
/keCBtVjYAXgfuZpprSJRnLh43JXbzT9kB6wbZaZRCSDVj5nsiNQ9IF7vjyPQlyX
088sUrijt1UpnbMNXqOwbEKOjxA1QAzcHS8xuWlTQMGJ7Tz4pFchsPX0FVyhvTTj
Q/UbqJBpN2/l9kc+f9ipeHof3jzZs0wwCnUmomC/xFcL1piTnLcjH7m62BENxcu3
jO/OvXRtI5AAX5K6ORPG25guoD58c6HRYDekVTV8eVU1OBi/4DNbtNlOREfFtNVy
uo+KjIEALKEuxv/pJngQF2z+prDOvHLLqJbbmxw8yKnQRtbnXY5byjLwfB6VN+Se
MQRkFDb7KGq+HEGtZgmFldD5YMiYAx7RGCE4puLVlud7wSvF0hqVxIEdhh9/ZfeE
5njiNud0XcY2cC6ZM9yASSvKBZP+YWz6GGije/yyz+Xxko2JkM3iNcGBTck4zv/W
MJZlSc+oWaQWZzUkw9z/8iXlvQgHC3uCoF0n451wvmsgv5p7AdVSd/nC5konHMqs
KngGiByiwVrso+5dxrJ/r8e3dVM68oor0MeBh3oFyf0ltuVC0dIZLao7TCiSzlX3
Lb1jTtCg5tUQ2tuN9OxKQDptu2euR/qoWQzVCXwVjFZO92aLDTowZFnTN8C1CnZ1
mCT396X7azaN9cqwYGoN5r7cUbKfoZTFIwwd0hKdL5ewCO8j639N/YbQ9wy9iukK
0hMSBMGMZ0QjvhHe8mUVhO7DYOrHyGU3jBQTeMLL7IhiC82ZLqG4jGTtZy0NrH8N
15oWKFHB/3p0ZXro9MEbAzFaS8Ijp5XoZNTjxZ75dmRDsHNkW12JXOGk399M8sJk
v8qH/ylsL7t8LRgp+L7Pn19jnLy9mbH20MhltTOz7j4IFUHDf+5rpsjPDSuLgboa
Bd5p3r+SjrO/4xTHUivQCeLadRy8viES1KCPVFIofNTB59F/xrw91jHEZ9aiIm+z
OPRhnqezgLt0eK2hh5rxsYfNF66oXFtbk3hetSLOaEdrpaoJu+7W/oSCz7G0VJQy
yORC4U6ZYTn7hB7Lyrol9Jdu8uvMO+KPex1PdhosuzSP5c9Vb9QPguEDxRMS9iKB
R25iUT+9nOzu30bQrsoMVdjQzoDqRKTwfU171LKl6fWS5Ix5X0gDxIdYMEm5JxhH
u/7RfCO6Y6a2lsgdPGCXbqcSjp4B9q6Hx4bEpuYhFcRXEqCDSGzGs1YoHmFZfOHk
TBcpRXvG+m2WdhYxP7XAApFsNFODas19h5y0Pwg2Ipnm47T0ZNQvrncNbkTUlTVv
btTa8ySI9+8YEzCDXXDr8wYuH4N7u5wXsGpnZxfxd3qbRVqqCbc45lX/HfqLDNM8
DlXoay8Or95KjBBQm1W1zi+nuoZj71u7v+gkK2PLRLrE+l6jr+KMdeqw9faEHdiQ
hH2E6Es5Y7MgpCGRsGy1clJLB5D4RYWvKsA5xP0odmvnbYKCSMjPGwJA2fWHfcnT
Vv+AUp/yTnIL1rho2/NV1rYg8vnbca0BcRLMnoa52S5nDw2Eq79J+hyaaxW3N7GK
mdEe9x+gBJ9jU3ILA/EyeZPmIa9u/Sj7Pn8X2zmD7b9JV/+ONJGUINco2n7e93jm
TqWjTJMIsGPuroDKUyUUZ7oJToxhuQH7EUBDPaWb9Q8Au7Lj3WOtU2Bdhk8E6GuV
V7KGkQI2x7xDfyZpHQ1JPwfsMTk6f4aN0G4HgWwR9B1dI/FBmMWa6NBvyj4cCxkU
fesHKh+XdHF3D2GhIa5cG99FAOOoUspHhNbQ/Vdrl7w5x1nGg0e4hN0LAirMapKK
WDrD8FqZIw5xHMEOHrRvIJaW/c1Ga3TCvntoDgXCLOLReUufVjYCYfF4grqT3jTY
9+r5YxI6/gHFcllaDepxs2LKhpNXrYvWxntHbbvspSef4r7KxF873hXccPV6vXb5
Mutnuh02dRaDiZb9NJLjY4jBI8Alz5BzclCt5dsYqCcDBDQ3O0ySjx3P1nqDFnEL
qGZA/K5c8zVheSUcv9ipDnEyGcna2Y0bUSh311mgqHO2j7NiEhfnOGLxPUwWh3hN
GhtUmnaPLERpZynH9ZoJaKUzFsupCDh3CpIZALXTwWlDLvMO6OskUJz9xJ9L/QGu
FmwUUWUciaAc0SWTdWXR6VczvXg2/MY49susW/ipVrh+91qlDOy/2uDq2EUtgCm+
QtOeTJizaYYk7eT40+JkBXE6xYmvLRiM9foyc183GenJUmTMisi9gOnERxvy+ah6
lgzgEOKYrYXHYKduOG6sNgcWYoycb3LRRR7gVayHDO/QAJ23Hb41AeKecyBurdMx
w5Dm/Bef0qZj29DVtU4r7Tf45ypgHRoVWeF5KLwcXNO5m51ZKZoO/XO7Cfkq0Jgv
FZI2pb2r20TIntVLma02cUZXZukbrtrcgLZpdED23HBkz2r8VRjJT3BmtvjSCvpZ
EyaDoSOugrJkYN7i2/oAy2H2Sl0dzaaR6xbUwIYCcnyCOT59Z/BSmC+RfcIVmmLK
X89iW1y/SCSVerOKCdYr359Q2Fp2UebsdP0tgsdQESQbfPPWTi8R5P3TMSXtBXw5
UQvfGvwtVJGMEeYppgs9gfZY3+JWGu492A+rAtR1BbrOvNcCp8NhZO6rOBo8e3kI
OSwtxzoDZaVxebERQE5Jy2b2XWJVMEdMsz7kEI6iiHt2OiKL5nSFC+rpuzflfBhJ
7R7f+AOJriw4acLOKXXRA/a7g7e/a5p7dBIO0GV+K7sr/XBtv+ICFKICFJC/QFVR
D1EpzKQIAqSf5ElZ5LWBKjZx6x49DDZJwyvxUzsSDkTP/2sDmTh46DetcyoLg+dm
cL+9TBAS9If74HeEfgyChviDqOEkuPhSVM+Ets3YrnX/E9jrA6QefNaX4mV+3/V/
OTS17/5GNqvyfCkdjlX6cFyfLDxh7qWyezYcvldI2bKMOjsQeFjJfN60PPo5UIQ+
UXTvjRjkdjYNcYB5WhHxoPlgyqC9PB19oXkLMEa0cnthPFiGm3eiTlUg9VXDHkQU
r/s3C+GBXcqZtqII6XihlhuPgXfC/DNT86jLsaSSpMWWRndrpQRKnLglAlgcTTmI
ZkGakZXRK5u1x+kwjTngOATPvIARbtEJU0vXgzL+TYUZ7G5l7LVnZKIdIndMZD/d
+0zLmMUy0sybwV/IFy3EpzZ/avq6D/7BbqwWiM0rFCzk2HndZ5tASnOmCUK8VbJM
0hX3njtMV6lg0wamcsoFPRyQM+lJVOMyMuJ1cHgzKhRRF5RUcdsrdIDx+h3pEYrt
wtnQG3MuX+4GxmDW9Pwhk6tXU2cHdjSw/r6hmUe28MFPy7uQFx3ELJWj5fr1ky3q
8zLBSTXJ+RmYTh5r4Fj0DOk2iv4Ac0hGe9MRPtI4cXYPFVznuuDL4KzM3ekicGID
19/caD/rsq/tTeaONepKauw5E2UKvCSd3HXx0OIF7lC9r45S2xnlJi/h4Ei7Sn+K
CVaMcKlLheQyS2RqQwZ/12O5cqBgZ9RF4d1giqfJTKu0FS75fmbJ0x0GMpWvLiEP
7M1C2iYwIproYp+mcEhEhDr8rVrm8AABbYZxvB2PlWaYNJHnbAZEIla7U7W+hXl8
WBrKtmRP0ZjQwUreUl+tawcJWJgTjZy8Fzf3ijeftxltZVe+1P42WFkiGQ8mm5Oi
KTu3IN04q/mRtaUshluznpsPdAuPvtUVIcT7ye3d4bjc4wJc6ak7NQo9yi9psOTL
irpx22cWFyGA6EwEUqY42WWwqiB8j/M4h070yDW16XyhNYaPBVA6DaTe3JRHWSXD
aTkpEgobTWRrrZ17EEET71lPW3L+sQOHtYxBJAjDrcsu+T3LZ/mvpBevonWZhwRj
Rb81SzA51UoRHCsZtq90yZvgjmQUdBmtJ54F4/GYA/vsu9+t0qrfC/oNqqGav6Wp
bOetF6rQ7bWUq9uDbUPoqCMbh279dqT+T9ML7h1zFLFexkrubijAcE9D/TbcBLAR
H3P5sm/Q88Hwxc4DDh8hXjHcH0+x3RWm7f8Ql/7WSIRcZ8kJ2mHBKWfePbhrKogY
fR7q+tCKrB/oB5LtGqYARIo8kv55IjmcUI7B/XFOq57cOaT9zA1vZZKXqR090VTU
Kufg3w4oOvNf3H3MR4BQmu8PhMC7fSRI53FXMMN1t+CaSxvOInbZ6/Kb+9PTZx1a
ecFJx6XDu0QjM85RYqUk7vy7wNPw5kU6OJ0vbWpfSLwXo2V0bBtwpbnYuF4yJDxg
/bvHvmWXI4hRbH5sYo4ZUuC6J3KG6O+RomAu9gtORkB24CLDJIK+M6x2oTxQsU3o
WfGsG+ZHBfbKrXqn7rOD+CIxbreV5HWyzXftq3U/qXrOpV5vnTrYBbl6rw5Qk1lR
n1w1O1P96k48I9GTq9qvHvJgfeeRw4+B6VplyjdUjmwEDIUqXHFwrrG6RKX2b5eR
i9bRQBvdkWb41Okr7sQNNkf4TO2lZFfvh/xYSsyDGnmrwjXZfwbXD/ytwanHrv3x
4eJfCwvBAQLB9ETmZ2wlQVdL4yFf5/r8FQiAH3vXDRe0hubJc16USRB5ubuh+MnD
J1N3f7PmXwOhvWp0NO+A+zcBYhWBu6t19RdSz21a1f9s40nboMzVTnMfvNyhK6sw
90WEM4Kdu4v6v7ZcsZ+xRPIHBvPmNQDYI4MF/RdHAmUhyefi6OfG9W3zV/7rzEwh
SxetqIiueDgc5Dl2B+5CQyObK4b4nKRYczHyxtHKlS4y/U5Im5dSNTagB58XqdQu
5RpkMGfJqcEuqbh8hc3hnalobkBlNPALCDkefi3PaHmy9vajUU2/MoKhc0u5oUP0
LnpAjqgp+5lanXN4Vvsg7/C11EDqO+V6d+JTq1Ah+AhanCkr4nMv4Jm08kbydIte
JWKq3e7RL7lact1eMHL43H3ygftGFITuTAKYuU3q/KRr6FyhM++yMwY6pAfgRm4z
BBEwbtzH4gZhVgRub6uG8m5y4qHPjq4fTQCCZPTPKIhi01Ac9GOC4Kf7J3IKxRlw
pt/gVND6aEGBeALE4jg10dYk1V4amV2iVRdG/NAVaHcMGfChi6s7zgH/xjlNqUcs
1dLS5dDVr/v4ik8JU0T2ha9YPiJMN9wYz+f4bI3iBuNGbDnWNYakwxxSliPO1D/I
tqu4pR6uwHHgKqHOohVPO1wb6LlSf/mkizdClo9arofwlXCMDEP6VPzFKlOM0Rpn
7FjX4snXr3531xJM+/ZatijNxvcnKtUEFdjNxX8apZZvNygzmkSYjaYiFJS9ta7K
Ri3Nz6H9W5EHIAtiCeXQj1MhF2kQFuR+LODAp0KOFpMC4FXOfNTZe9BZadN6QYeU
kmBQJ06OALw/geNn7y97R3U/yWAuyQn6nqeTVKYODr26uHmverO+v8k4vBPZT9OW
jgxJABmb1fkNef6f4Q3J4lm7syI5u2Ive/JjCDuGTnTRsJ+yjGZPXRNjmjiPbFMU
rOeBuDzHT4L2UjGro0pWxv8lQ5ranPzUw8aZ37wVWTc+remG0X49reHnFnuBSbFu
iIUTUcyzsQYOk1HAAjeIwXVG4K+44ux5r11vV0V+h8DwjFIjEvvBJVDdo4+0hmrP
MbKB74iRnd7XeYJl/oS04VCl5RumitbJhoMDa68LVo3S0lx7AKt04TVNN1keIIJx
7FExlJfrEDwBcRdDiGHA08Ar8JSbP87IOBcUvOmkIzqQsJf/4kvRNVGa74Clx1lM
xK+/3ynekgLw1Qsx7cqLYYVvroxPaf01JeRWB6Pyd2QB6tm/i5QOOHEodq+akzpM
axIpZGqW6eZwCl3Of5Hpt6ZOSJdyphIAYtRl3qEnON/D3RiPjhP4M962K6FWod90
ld8h8+3UPS0ujqAO9d/Dn/z/fhgm/nbidmzVyNAdrrSazkpMfgYkpZY81/sEFnET
2hgdZfMISTUBCPXfXj0WG9He1JH4GIQqGc6ZM4YajGs/IPoD0qhkHzE868h9U0ca
TjjkNj7sPNZHbIzYSgG5RXn/fNKDJ5LmHy8qRo1rjntgN3Lpkx2mcnVPB1epoq0s
cVFEYsunPjesJXBQBv0KM9FkB42BswjrJ5QY5I4sNX05O2EQVAZnSIeLpGGdi8HH
H96hOnCW+EnRqH2IzmoWswwNJYOLHodBCpYV3wY4LHq2119Z4bESRdfg/U4/FHSb
pn7QyGwkgKD9ebQZuGkOiwRSUpl+o51mjDwYcEPJcrzsqpOaCbwPCI+GtNjSfO0B
hOIDDU2XNFNgUlAf6xqBVAQJWEoyAsNm5txht7zdsbqyNaChJ1otmMZksaBN07GJ
AtFt7YwEkmoTO9inQmLN+hvgJQMSx+dustiz4V428Gp5qXGgtFW4fU0jhDUdAWtO
7QJtGbq52o7TL1XQM5lnNmnmccsnEYkl0K8mOe7YjI7EdNLogyPIF9iFQaKhE0RO
IXN8AfzbTka4+w0btZBMbXUWh+2PU+ziqDjqtymUOsdhSkWyz/fskdz5y4kRZFJH
k2b3qFcdFtnnP8ABoG7tnemeCHcTw/IBfs7bXDlQtcHHJyK2Pj/Q46iFqA+t4UWW
w/SeVkoX0iIiUVfOEZsyVGY5rHFW0npMK6a96+SjNRVROctJyotP1UI6rge5zs3S
WlAHgGas4mbtBbACGRxUHGZHBJigWf+/r58BcpX8wDiDM7GKt1swSA1YSOZu3T2o
NSaO4AMr7PHkydvnapixYMl4O+UflMZWstssCO8y/9MCEwFk0q8K48WkgLXciCYP
E1OB0SRLuJht7kLdCEoamZcyHASK7xCT/Olv2LGhDL+GpdjFSPGjo6eDnZTtONiT
4laJ/PrP39EkedcRo+Pyn+DU1jkPmvQa1nn3rCkOSG/0vT2ytMmzvjRcHU/BegWx
N3AJMKQILG8F3pI1GFK6+GKkSwYu6wt2DUZsXGduZZEMsgLnxoq3nYhB95lXuZmR
sieW2UNkigUb1J17okyPTb8b0wl49V8urch3qERlfQaZxoA70M7BedwdVo89cscy
eDYde+WTFOxdJpktrJ6YRYulUbFGm0SEmNBnVD80XS2KLpDSynKZZ110Ze6bmIOg
Lvb+ldXN8fsiAl7qjI62PXUxTEpGPspAePa7nAc+xSijJELs8O9JIHJL89Bg0Csj
kTmMjXzjCe3tZPlFu5afo5VKhlu767nnn90b3+ysBhGIgvNpPn6n5IAHGOQke++j
Hl7tIe9IU7oINldCqJ3k1SPSEtCn8I/hBZVeF1rYMDNtZz7ikNsJ/U++K9ALRcN1
ZZO+dzROLTPeqoYFczshM0x8vsTqVpuDyDYGqame1KdgHjilGix6yWqn7/aw3AG7
xVa4Kn9lpNncG+ONLa2sOuTMzaA36GlvaWwd8kCD5+Jrro/OV8LRxizONktYvpcE
yAneVYTtSSuGix28PG7CWht9vBzv5eAmnCytUIWnh0d1ASJN/TO22zs5r80zXQ+N
rNLXzrJ28iihWCTttI7UEg6tN9+zstvCSorAChk6mJ/3GGE8NReMjSqSiZ63YLnK
2igdHXwvSNeN8WRbzpFyf32dcURcOEfsI/0+aPRmwURiChrzKCDXCm8/AfdAU53J
SVainl/qbDgOLWYJu9gP5SLxvNULqL0jNWfnKZbFhSxh2K1Ij2DFsxBGNaKHzgeb
WQj6W17fQCSDJWKadFrMZM/mGftN6pAbonS10ju7UrgJEBypVosm92AMbzj4wXki
MXhXB+mrp8hE76P06Rgyvw2C8wAIjr7hnPqes3Pq/6AEFfZOi+S1eNf25m8bj07E
572arkV0uuUdHa4G2cnax+Cx85nb0U3qht1DLeVBIi3hyWbok7GrAdqD9+h22iP1
PKB1V9txzP0BMSgTvpzuuKKvm54/kR/sbcZpc7nJMapp8UsqVBHM8jX9IHwuHqOO
g+I0EhlYxH2MnRv+Tgqvi3K/tyPN3bkncP2T5VkHeuYzFi3ONFY5a8T7PtqCVTNp
OETi/qSYReKdBRfXSR9bgi4UJMG4FOrTODh1z2ubjkhDe85+/kKaQOksrmclWLIp
QlcSQ8iARswglhwRpARUpzVZV7kYBqwTNzLQutuoiH3UEWa6rRu21yMBVU9olxCo
/idGW+M+LKQFiZPy8OujMJ0sS+seFqoiEenXPEji2uk6PpLh4zyImkQWgYLhFzB+
s3HAVdhQew4pnrr5VbnBtaXccoRlJ6wyTdBb4rM0/6S/TRHaNijoz0nfpWf4oSTD
BV0OC1I0tQhLXLq2dw5UPSzIKJYT62uRnR5k0p82f1DPRUck20f/2MN5JPO7+jYo
YGtNVVzxlTBOMHM6saXFbWCGzIGBOXZoHdkYQtkSRYZGTYTWH4Z794Cnd4acLoZ6
94+bpCKS0Wu59zS2hcFiqZabLMprv+IRquWqqRuKKD4LQb4qy/lo+Cdtw9TAIDw6
m5heHa/5QWbdHgk4AnzsVeOhAU+iLIt9eON/pkorPmkf3N3AGQDx8sTqESfajQzT
8E2B4h4y+urZte9Pnxje8OHjkoLHuf9m+lwvYx8NbAKuA9+myh2fKc5btVql8ieU
85Kt7dOHEtKp+VIdMLjJ/BbZv4LMXwhIaxghJwrzq4drD3Mx7ZExBWpCLMB5bVrt
IjDWJGeuIlVy5cIQ6x5RzczNafVZ+76w3yW1TTHzRHJQ1lwtUF0jrk+PzfkRXDMr
5fbQ8mKOFzWqEIhM7hwOO0idsHm3GISf4Y26Yey/Tl6lfMWpAg1YVgnLLA6C8mXG
58yHuuyzad2d7/gG8g/C3wAf9N0WAGQ8ybQwq43sVdtio1/4NMjlbEu5uFnYu8x7
5og6KOZybMz7BJM+1ysl3EMImtP2aMybyzVAfHHQdZTJYc2ldgrHOINkzeJmF2rc
eADWbPGMKcKcEEVQptnvs2dwCvyNuLYzopBvCub5qeASqbdoVFg6ZjCS42hPc2ly
6zoU5zoSUuFmv2qDX3pFQDy33PXt+XHeD9TToHosGPUyCpi/6yiIEeR7pQNprP45
BtRggjOjvtRWMFw9vx6d5/Mn1H+e7pkAuWhu9teCkXgSNktGb0pKFURbQfG/zzYn
s7WlUKoSq1X0nrB307tx9IA4qfMmT/oeQu/iJZQXwWFUxDU02tFFiWGi9QWM1cti
sZBOVSuKof/hMQlAWqQ9+mycfLSQIiuAwKiZ0nDahX+Q8H+p7A/309x2ricThdFl
Qn/ku6od9M+4Vtej/712rpXEU7ZoIHXnLbVndDeMVeTsMg9K17WDIEzBs8siZeXj
7krW8TU7GNm0qJj84nxP6ho+/RqoPOepjq9x5K43tWeDD1PiROAqD7PJnGASNWHM
gQysAv4gC6eR+pE6phCe7ngE0vO6/ugOiLlV5JYikYACMvvl6nVQD4pq6O54cYhh
S/majs3IWFwpkJUez8oyko1k5XMmyM7dT7EU76sElVbLGLhe4PqCK88A54K7TXPg
FzmZBWjg1pCuzMC5jYWBh2gedkalyW+3iu32LP2LTMrnUr74lIwgX8P4KxpFxT0e
h11LxFFNK7tn2GpCvlK+JsmdqJfYAfRsXsaumXB55UXUdQe1tw+nPAB9AHIibDOM
rluS2kw8cgh/GbGp7H51AUhKYeUpKOJTD0QaX2ULNOXY0tbGKA3jJvBl1K34hlzK
rReIzIyXsxEtkZ965b+dmjqC3Sf1OYaN0Arqpr5ps2iheMZCs6cVtSCfC671pzcu
bI97Vb6sk9ZWB81EazFT0V+1ywBnFOI7jULvSFRQiKJk4eFjG6jfuXS+Vk/x8D3d
nyAfhOlKvvZy3mfpBPmtFY1fOFu/cS8St7SIbXUQZ9bAYNY1CPGK3UWshelgkOdz
hzEEQ4hI40r0Gl6ORpHDt8JULplRoNybvDNDBc2Ai+1lBN+DcvQUGdCWSMYetpI9
u7vhSDMWeTn+GcJf9TzrIGKwqK5udpXIDJ5xxP4TIA/C51FUzoAIyM6PNfnH5ypg
QXCPfUFUxhJux6yOe0Q3/enns6yBNKKvMBQSh+mXkwba9Gk9YcVi99IQt8tRS4jf
xgdhgNb076MM6g98yJvY91yf/CbhcSOPlyDVrM9Ytyxo9DustA+PE4k9LmiyUy2I
k+OvTZ2seFj3bBQaqOv0lAuzmjJ+Uhck0X8Vnimfvv0b4g3XgBqYsB8tf0tpIkqQ
RHW+Ed5NvflOqjHc35NB26HEyCNKPUwqz7DDpvu4bxybOPl2ioh/FQ5onuTGw4Xt
EmtEUz4Hxs1MbcZ/5UBtqm0jYLF+8XCtXu1rYuzNU/IVnuB+OYw4LeJc2+4G8NXA
H0eo3giD61O0spvBB+CVQGZQACcBQplEgNDee4pSYD+Zn5VQ0RaZUmKklM0WXaU/
opXFc5rxmgE/vv8qP6dy8lzE4wms3S3S6DrWjvVNvFzPbNrcbTRYy1co6NwbQXK2
Igg3FGje7+OW3R1JHXD/WxEKgmrS60HzX/g/Qajvubtn+1C5r4c5pie1qW79sII8
aSkOYHkgUKSJgaGZnaWonaotXQl+EwGQNNe8flt2pHwXu9GVj4sSHW/n+Mt+fz1c
znZ1ULyv9STfiudM9gGYi2b2e2S5idbmbPC+HgbHLDXIh8HWBh/7MnxUK328scHQ
vzQ9fS3W/ZdKABsjwlNBqHWfgJTMD/PyfUDgPWrhy9oJdMZENkESGG6IFH0ldzTP
kJOQ4bRH7wJNgw6TCURdEHsTjRaNxV7FI3wC2fgjzgd/PcEocp5UrxHSV2DMDW8f
k1B+SmkL9/KQ0cWBQg5mbdmQfB41Af4DoGnKIpNU31AGDCnmZ4W0/XjDOR2PeR9Y
cHE4wQL/Hw17+urDK5R328hiznoJjF32/SnrN8C0R7NK0PUortC7+SEPB9Aekh5H
jQxNTrRLDgoGmmQ8IzMC17r93czz+2Y3UZqKZmRgrWDBOlfOSh3S6ucH1pvvrPsT
NYoqdoxwGXGBo6O4+VPJxh7lwTJRiNLZUvW+rs7TBGQEEULE35bmNKmHYCiqfrgQ
HIMTYQgmPSXsozCAPPdHi2CU+lZNAhqmRpgnWpqWjExi/fhGZsEV+WWEJCEgBIWY
Gcv9dOGPlUkPWgosKdt5M486paFdmUUhIrG1EzHrMKXsnW1D3Sy6IW2sZfq6WUDv
z/KNSTVGN5opOiTdyEeo+ubsD4FrOFTd/F7vMgznMOXZ7QZ1UUxYFHCT4CuW0yq3
NSLbmm1EMiClNXM/6aoLGMSS5xoKdfeSUESx5Hq0mkkWWVFz/LQqQhTvJsg3POjz
Um0QU6jCxtua8xxe9JgHzbIASn2zrDaVPzGNvaBVp7pWXgDVjU1ZakntbkOly0GE
8jyVtMxRR0Kb7m5o6RoxKqn7D6ak5LZwS3s1xwAWpw8XsmO22XRfF8b//qSuBpC+
Clidi3gRgF6oiKLLDCYtvriQNs6RdQisSdy8epsXJ01YVHLQWfb20ee2KSy4NkpP
Dy+wSD4F/Xkvgv3tOUHZyyUCFT+dnvrEGa9eKLd/TgkJXmkSvNp9eLB/8vRdHHGt
VuLfCYEOzXb4TstKl/aZ6Wly4YWTivRrn2D7UYudiA+SD66/J1hWbWRHv3n9qVcI
yS4zYinJ13IqVMyhljbSmqiCzFGI8UJw9UZIDE0JjeqXcQPD09/a/Be9TqskoKTc
VY7VoscirbaO706bdjsJVNkXbBAYt88+io0VikeUnHMWzzU3fU55WIe8cJ4dFTMb
qqhDwahdZhrHeaIaFsf78NOEY/FrB+S5kFeSpm4FTTxB9F8LipuPEthl6K+bj5Tb
JMpV7R5HpBCjXzoG4nMg5OruOVbOWd4GiEyQlftfnmVeU1+VPXWtbxgGEhLisPnm
ytvwjhPGmGj6Ed+vykWq1aIjpJUvK2ePGQy+UpE5MwOfc4lpiflvMinfCL3khOiN
yDlz2txTf08ReTZv4n5whwL92oSx0iG2CFFx7r8wRrc4XT3JE7haY8sPMdFyVD7r
juvpHHPqnlwM9BwgRnWCwldj028WPocT+nS52PvRZwGf4wROoWNIMA51Q9NuHsF6
phOc4ORTiVRpWLDEW1Zs77ggTyB5b2yv484yWPeOupCghICNMIaqmTQ++pYZhC0U
SNHFIS51ukvvrrYc3OUUPrphrlVLqjpR5UWix7JApUAe/0LsObgwDcQ1D9iGR1Xz
ufBNN4FpmCt06wiW3OSRMvZIZuxWLi3dykFNEzWPGtXM/sCBdCPtFqdEa3ClYc5y
nicFsKrmoAYRDXt+NVSRCz5PwgIx+KP4WuVqy1GewiJPmS8WCLEWUBaas4uKv2H0
NNB9AcdIXXpZsrpy1cnh1WVA1hMF7xUZKEZvsiFTVgQSbqtJCxxQbykPDRDJMkws
U7iZmk1ObsZNRlJOAiGi0gcxhbbwUhqAiWD6Vc4zD/+xHssa5XnTc/nsjg2SUnsh
8uJJJLX1qWjU+4V2jbCm4glY6pdxc/kB1mxprHZcNhXPtUkGmmPmS5YIVIQ+QgA2
jMWh8MMcB6qEOE0TNUQxkGZYOtS0XCmMvsY2nb0bXCiGba02SqgzugXcfTYqhAwo
Zmiea8zvDuVgh3au/S2y0HpH9o+8KVq6kcLutYIcgG0nL3OlyCGLXpFukP+K1SxZ
Eg2rlARWirUAyhI1+6vnEBDua4oRODkxuFHLXRVr1xRbUAJHN+GNKd5YUyhmB17z
KhptPGF/HaoOWoV5ccvSRhdKoUYH6wbD+b0p+n+FiR6kvc5c5UgA6sSRu79nJz0O
TFva6RuXfjlAfRAG8LEonB4rQoWgoENz7qShwPzNHqN2SEXcsVgQdJHyiaQ3PH70
pbYYI+9Dl3ku0aT2YemhpcPr4PXmdSSLxRaZcAH4f66OK3LyBIwDCtRPd7ZiRP9X
wb8bbBZvjz+cTXuwMaoCWEkKTWx9pgZfouqu9ty4ogLTkr58qqncPuJsFIz1RqD4
YeiwOEvvuQpdKfm2fDQG4II29JB/xBT9cIuBW/wqtJPdpucjevf1SSpUA/eNo8x4
YpQ8pNlHvtIM7Ly2cJ2Oqk3NuPCHC6jeiuqhaFV3JvQ0DbTgsXhkIkOQv7SjtAcw
TK8Zqa/W5RIaP0AW9l/BTT6rKJZdEsEewGWsddz+KvgIuUtWuuBBCzGGP3y4WHR6
tSi8HmZiKrPZhxg6tnFNbOFXEkBHkndO2Qc0FgSqNvK0sTkOIK4u45s27KT8zNTL
PxVfiYtiovE/S4U/E+M1Tuz+PSh8FbeO4cfeetEWvNV/xoJosJVuv2wZ5Hp4EVzr
4M3HGR/Xkr7Zbp0DAoQyCxx/ZlKdC9Bnpals/Flk/1yI9qL1MMgWg38NwhY7ieVT
8bgP3wTCw36haqxNjCO5Z6LV9Hi/JVsoSHhKEkzpctygcWn4gbKLQjcDHiVzfsvt
CgFFLX+4y1sKTRr2RXRByAkUX3RMY/mUMTaxjt/DFAS82AX4ZdjI9SQgliUwOyyL
ICHxVposUeIas/Gx4daPPefMm2+tfU906tSFDn9Rk7r54hOSK3hbVcZoIhpjU5cn
JpVUXm2FahccZiic/656utAvhJfF2TGkvejBFW78v/g22AIrvudtRh3rqOo46qmR
1Ydj6k4PohbTRUO1Ud12M3eInhZXWOHbf0CEkfR6JRztIyAPyQWPnYhoxwEpxd4s
tXgcara3jBkKoSiQ+nqOsnaPDZ6eitObuic2E9I8x8mHUSOG1f853EQMrSmknYUF
LpYllyzIpHrVCP9qZXk9NV8vC9yx9xrkUEMJx+E7PaQHqPi/LqUM4TrdzhU+wByv
5JjM08MCKbno4y8SoW7Lmfpj3df0tLgzX+Cs5VPNPcRudHHdEhJgbN+TjmHTUrLe
gU7Z7TXQb6bZMKYdZ91UJ+nTdKnf8aXKbzsFK9O/taPQAm76CSbkSV+evYx7hwUd
hnI09Ogiard1+Zn/LbTpIZlndRUWbsydheKvZSlUDjLUYRC96HEn+uJgYaiPdPw9
0pXncuXmFkewAKgbl3aOb1XUjReK2lEhBAqHJNkGApFeZeQw8JB7zM8mh6Tlx8kP
2BAOC16n4iADv4RIR29ImLyHiOrTTOk1A9ZzOVeLrh3hC3wOSOvm2o06A6TNQ+We
zR1jkCpoa4dB4Vzux47ao3k//8YG1SEd+x5yfPMgX7Y/qpBmAG2uZPzLuYbP4B1F
WNWdJtDlBW3JRXgvmUwqupoOWo6laWXDvgRwatoxHh94v2zTCiKMX0inWxnJcZJH
SXUU0H5/PGd1qYR+o8kgNUuQV0QK+j1J5Q0rpQX8rDsFsfkz03OXL+XYocSgQWup
n52noGLqf+lK78SauCYeDMZe4rCDGsUaEC5zD8rD9YObpYGv7F6C04ewDO0xxJc5
Q7tKmSq1HU+6SgDMDwPgzEEKwQkfCm4NE4oc6/QPxaRpOCoRsZ8sFz4TfFVSYZRi
aLFTO9f4wNii4nKJ5RBPwdYlKXHYhAn0+mtK9hJFHlkdc1ZhK4XrWb3ryYdT5w1v
z3nST1i+n7kmurOv5ZM/OeiSHVo4Ky1Av0P9i2kvfkysF+flCR1f3HUVKUnGxq+G
gXOfSvY+SsGUnIlVQhw5DbuPxHyuNEP8h/BTdr1mnw0GUHw1cd2bxhoNFyC60NcM
cHtmBsXqvXLRGiWVy7suEXP+vGN/xAdCInL08nNtlU6wUIcfxeNMQpZucGVPYLXy
AnIhHkld743aKsd4YhpI3XL9QNqpmA+ozWi1ZlCFM+VKuxNwDSTViVvIJl2Z0+rp
yObSC2w3eGNdF/f69IpuUG38/pdrUPVlPdrQnV0bRR9Gm/br6bDVBYnyJRirU68u
idghtyG5DcbZnvk+45HFis1gOrEg7kqRR6xPe2aR5hxf1YuXOFYuwtnkcZgr3/sS
EdVnhhi/E+8ND3zgO4QE03PX4LAlW0t4aqRUrBkytYzaJhshFZsJpFobgbLEOS8M
N+M892sSFaVbwu8K4tcWnG1aItkA6iMhJ+j/vC79W0m89ZYJWhJdCwlJlMfGSca9
fc7+J8G127Q8TA9OSBb9taxmkBR8ff1wBs3dVyMthkUlT/+cwvHRoc78Y/NsZZwL
guO85UywAFAQ2K3qVXIEtQKupywCZcPaAMARufDO8O/npqu6KBjd8OjhmfD8ItUR
u+5aZyTMuRvatlnT9SPRAXfIr+iyPoLRtA/bhOuoigFpois1bhH48mMnbrYCxDO4
Ag0aBXox5S0mig3LUkLCT/lVbmyfF7KrKpmG42RDDwX8xenzcXd5TeQCnTNSCLy6
rR7ny53pAm5ygZCAxYQDIdj4rPYCGvjLVI3k7n9/sxzqhdWPEmkeIcFQZ8q8wQjt
yY32d2rwEoQvRAESo6/J31NIpqmOoDrRzVtfLUhTGJoFB0BSJfJXeX1AVdzJxXgP
jp9nvFB/eTRfmJnuPWMdpETRWYcAg5CtA4dcoeFgZwNhPX4bcvPe7gu5Zl3RLgas
G9N4EFS7qWr4xjGhsd/lF3Fwz9JUpxVEPH0iGz6va9YmHgSBLsUDk3mffFKDe26Q
Ndj9xC3RhGrZtyMEAvxDHirZvESJlfNoX+KTOd9ZbSdxbUmq/cmLSI7HqIFF3fDE
gxw6/1DuqWNZnXFmrAir/2nX+X9ajGzuXEHAko2bkcaWeEHJRRAGsxk81GBR0Ahr
3hP2U3DQ9ZHCGI6aLn6jyBS0B7gLeBlp+EH+y4dRNDY=
`protect end_protected