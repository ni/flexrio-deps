`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
lo1aN7iNdBTLw67VuJOtfVPhg/1VpitCNxPKK8HEDtUHaqHRn1PMsdXOmcfPCpz8
znwG9D0D6sr0GbrNxqMH6jMkhx4Kn/e2caNFNGpc6MKzt0SFQ/jCAsu1lBhFGorm
Ex603khHIwVgdEMRAhkQllJuNXd/kGVTpABKJMLW552lrLNmxOqhtj8/vz5I496p
K5JOAnwPfvSnNDuGyrao1N3Y5rOyUm7TiWX7s8kynCK76HzN0ALzsEMLFuSDBuUA
3EDgWPi/CWCLgdpIuXi584dwM3DgroavT2Fq+1E21fDtjiuBhJsY6Dn/j9bbSkqr
QKS+RAsp10aQQRfKAnUiiw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="yRMVo1EH+xh72XB4foxjoT/vpaO5vbXS9GGQiqnzK4g="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
kKtjDb8UGeRJ/o8J/IXKVVNa4n4WP0X7q/7KGgIZEMKsoETK0SCgu45FB+jGhKbB
KVtkp3HQQRNerANy/lmpBpXyZnQFMZSFr0JrPUG1qRiugOTLFgfBJ8++8gHuWV+v
w0tiWaL0RQSiB7eZDW6exU6bBbsEcWOOr8SJpTFkvaw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="tNAMLc8GnMnK7Su52U7H28xMtJ9mAK5o4iRe6e85Vm0="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15696 )
`protect data_block
q5JrHtWb3128m5rljJRmkpsSWyEKnhoehHwKVrgGWsVWSNDEpCGHa0E99ec0xzC7
zM7G18LfFN5vZ9RO4QRYvMs0hIqJt18lhM/UGKT0k1z0+E/ImZsYhYEdw1DxkJmL
lBIbi+2rro3ublJL9fP2LgMs0NA8R0RLJ/vMhOdStx/9FbYjFapAzUpt4uFt4lrU
34aWGaDb2V/DDv9aG96gwoVRoIOa7dHoX30SLyELJ8vhK277hG63/rh5RKSH2ORg
G8suR9i7gJ7ha+ZL+rrl2c4tLaVtM/aJ9EdiV0q/Tos6uW+005LdJj5sAM0jz3hw
A+iwz/nTVM4NCBwoCERA4jMY453Zl67tQxCfr+DHN+8OuUZqAGHgxDxYbEycJJT6
jpWeOP7xpF79Fc4Es+MnA+lGGJib3IlzPMALqlQrubh3Ah2e1+4axkfBceqUtcGQ
dIhZ7Znxu7k220QsAfiv3tcqm2aXgB5T3yBwtODwAk77xNS36KzApBdOmlOjaxan
7zewtNiK9dfDIvUgXCgHNqe3ZmTxGcZZwiQjex1lRvCG8CDF83k+crukAnZowh2x
PxDNciYPlW70hHqnR8c41c9W/s5HKnz5vUyWhcswtf/IVuYXK0ovj4wKDxl3m+sM
Yoly0Huj+z6eHWrM5A7Dw0jl9rv+YK4XBg11hxUidhxkF053SAmyaYB4UEIXGOTK
DUfg/KBZvN43kb8BCgX8anUo5vAhE1Yk9JyU0ryMppgw/grfRxkrBRvty9WSvikp
Tlr9dIWzHK9Y8INc+7pVwyH3OfwiI8iwTmOveDFzaEfd/+N3d16c4HUhQTPwPg9k
skgcIsJcn6SAf4zVg0TLy98QRDlrGD+mRtB7LMKxROPvLnsq6gmyHJgRpIOyeq4c
X7q6EYSuqZ+EdYWPlGyrecT/xT33jzwIAhIHo8zh2lARJv70a4X/SOtEOg0ALDKM
E6riQP+9QM268PccZrV89IAQvdbwwQOq3VwWqXWgIMEXhej9kEQXfNQGR/Lpgz3B
NC9PHt4lW8AcccsiTw6znM3RgWHiAiryvAszYQvIQaWshD0JL99a3NzQ49CgsT4Y
qWyhUS5ZGXeSQls+gzPGWV/f35oAFwE1RDdLxLLw+xM5oRvpGjCFI1HdwveHnLlG
yBFJGXImYhz1vqjvGY5tMi4S01XkUtI3Tf5HEqVI6OVonoqFHzbXZLsYtJuzw/Nk
dnbtVkw2uwEvZyoADdzudRuwwkbgvzw3lwnDCNXkhqFOPIJVLdfKnA1FaqUag5mb
8LzijCldIWjqqgSe/Eja0Zz5L502V3NNuh3T68vnbm4b+/2PYpIaPXdO1H4OpFiz
hPtJ7Rd9TlcyLjzdM74D5sAvY7RK2wB2i2j19041G2QppjwlkKOjz9vhy38d+Cw7
Tq8bfJ0WhfyPulQnRGlLrem4qcKxylAxXuu1Xd6fx+mJOEiG2GqWt0eJ9rOh4joX
Z6UoKzrVMi8T/oJhs0we12A88jnKpRgfWp2p/tv1Kv4BeAeFdVV2/kh+erLqbKhM
7VMiYBbKylyIkuUbSO3QhY0NDlnMzZc2S8rggMsC68fG+p6mIh9s/Hsk2/ERb8jw
Q0QCSUfh1CCv8uTOO0CX6GFZ1S4wcZW2MR048lhenfMm9vPthhYRGUenig32sHNn
FxM3HTGYwEEZAsOycueAld7p/FTHtLMXjkcQOIQmBDLL9vKsY2JQivlrP6PA62k6
fU3tXFCIyIhtB5ySs7eY9NC5YDOdaTtMlwdfWZthADbItV/i4GhjMR+GxQukbLcR
xbVFNs3QGFdQpE13iY+FeHLhy0jSamOBuN0D2GbHaZAmKVGkpjdaoOGSyJw4rvcG
jlLfGGGakLnRC3gEB6OpM3oBMYqzyk2RuW0HC+4BSSb0679JNzyuMS7eMkZD99UY
RalWn20wC9XxCtIzPC3cXoL65EjycvqMzIPIqcAgeRA8lN8XzNmQkpeXJkbtjwb8
V2pQ+R5c6mfBdK2V8HT53QY0+jZ67t5JiidOMaWZgzzePteCWfq5FZZGl6YEL3qc
RXOWvZeIc6fsAhcCNbOhvVu6bbCy0BaXCnh/W4wyG6WBvp7flmBEQrozcLlvsbtW
oX36mp8BE/XDuiM2MG11Muok9qsvRnhTbtW6bOWfPZUZGxOZDGBpJyHM9VmOueqt
9CLB7toglZ5S9sGFVMjYD4rLicsPwJSzRL+SxOFoFhUuyf7Hy1kzrgMUdRazNaKq
TOqBzFr9TLslEDi/jhi6dqdXqzPIPutD3WzrvoshRNMdgQQRq5Q6C0nE1O3xnfuu
OoDd+cGCWeQ+kfVYuUW4r1mRSe8tASzXjtrPTzL7bEKq4SElHWO56GIlSxjs7MVK
DKVqTUSM0RxvuTZ8wI73oOEOPMJeiIbpXTjFxlVMJ9+kT1/XQPNOz2hBiqIp/ap3
7KO3SpLStEjPtSwuQzfqwxf7LkaMYbbu10kS4QCtxfh83135pffkD08eIXxmm1ny
I8LJmz3QmltJ6Skwe9vq0rARLafeXDppJ+XpeXF293nkOaIC690Qod0xQLCdC6A9
+/NOL6hZB90RcUZf1eEomLSdyIeEegdO8MqS78uetrO8aY6luhY26CIeGNW+T3VE
ue3uaxMTbFqhmn+ZUQhO+8T95dMdBmDefNWghaD2Zww/My5J/VJ5ijCklz/uvnug
anqY4hth8BS0pMkLaYb1+233pzAz2FCHO5pSal/wFuyQ7QGVWiPItIUFKkr86qsR
WawyM+WOzmlY7cpVQJKEiQNprSNgmGs4gi7TkElvGKBqwIk0KnJB4SYVk9ftWau0
V3b9uJ+eZEz1S+3fYcGvy8wrMZ6CoDLT8zWXWklStJ9RWYMYZv5AgJ+1p4HTocwI
w3SsRd6qB2jZ5xmtbghKah4qPT/h6pIv7/i8lxMeNZpbfbd6FFbAx7zCnUUdnBoX
DEAVJb0G+15iijD9eTyaOn8c5IBlltsjq0xP7b3CyP86bhT9ir0TQtSlkIx7kf1e
QPrOIxaaWp9JvKrTqq/jrUzQ4saBzQrENP9oDbhK2metJpJNDYcGozXSV3IhXYUe
mO/7GZd4RXfaDf+dGdd/4nQqh6Pr+t2O5udIifYC6YPBkmsjDxBe3NPG6zI61Sw1
SRwrxxIefHuX5NmL5YbqV9QEGcbNtCEAKONOsk1naw3eHqM3BsYuCCdsos3G5kh+
l0fwCL23f7nC77hsrAahD9Ipw5XiGYhn+D4z5h6IoHXRejYmFAXDg0NsO3BFi8xo
YcQLELoico/8Jz1qdQHNNycNy9fYnZuPJZ4FCZfk2/6daSWcZ685JgSWQtPKfWib
uzUa5ZvnkQnZXvCnfTmFf4FU3p2fsyrUhe+KsLk3yOvxz/9sAf567+5FZ/hGZNY1
47hCZcaHMWdEsHgWnhhXSPdEENV0uva6Rxq0PcXfzdfWdGWg/JUHGZwKFpsovHXg
Xt1aP2Dq+TbTUXVJNMdj3fk4Iee6r5C7LPd8rfK847jxbmC3ZBA9Ij5unGE4QeKr
zRsOEPue+EFcMQ9lw6mq6WLcmuoKo9y13nlZJM7IBKzzLxymSMl4livnwFWj+jsQ
FigmQFqHl9UAkK0Z0E6ActY+cDR7oLOFeZgbMf+tOkuh5fimoGDE0Pdm0acZgPaj
k37S1St4hkpPjQvZxy9AKM877M7ZCPArO5o4VidMjfS5u/wlpdVHk4tJJTc1j16s
F48xLjRW+uhRXlqkxPQI+N/RZpOIGSSPDM9+d4Zzz+LW3exC0sdvmkLl+zhTGGXC
DJ2//yJdOa/+UcMv62GJ1lVTa4djD+BUBbiFEtfSgvlqPUZjR6rmtViT3eeSVmk+
pgBEPdJX4ZEBo8p7SdHvxW5nXA3WphEPbkxsMA2nHNhDNkmVg6eFayCRbZiG1BmV
5ae64GNvCQy8IxgN1P1l1L6q+yH0NWLXBiBkYQnEOcNXSeeO61lv2aWPz/pIC1zi
mm2Pa+8QkiXyq1TLfFSDODCEDl5nD9FBLvxAq0H47J1FWYNXqaW0z10ftfOZ4Om8
213wb7ItsmFySN0i8wEjVIOqgkkXdkBR0lqQPsS64q7C3afs479AYLYr3Gy9RKbq
2Rkwzz6kL0UtRUz9s77+rFpt2w5dRRULoxGy2W+NVHZ6atjsGnPD+lqOK9xSY3XZ
vcwcUnY2EEzerIN/39K2Coo+JHNKiYNN4QQH7dZd66Gn16fO/8nN390JNZNJ8M+r
ak/YiPVQD7+nUD0rOoS0YjY4y3INYYgultHjsPA4rrgzjl14ipxV+gq789V3yPhv
DSeHe10az4Dk5UdRrW3k46ZKcWrPUdv7kRCAOjaugOFhhmzwZGHWE2pSHky0MWjc
qz45Vq1mfsZCmtxsWHOVjGVjAXimLXvqnBIM8UmoBj012Y54t7W47Makd2RA1w4g
qgKYiFZx7ZDSp48rgDitywu2H0ymJFQS4PnJHrkPPJIwRLk6SlaEvfPLdbGIUxyW
NkuPjc8cyeHJjQbPMPrUgmKrJE4xO7/cWZeKr1TTNuIqTJB1nLmeCjcnUt7C9D91
u5qghX2ZrDDp6iuhE8Z57bOZ6U0NUcNTefibutPEurcqRf3vSXH2SlAJ1Pot8g9h
X0abyFrLx+C76Mm9CIO+V+w2JkPy4/lvGqh5++uxLdZ62aNO/o0LKQId+MrykrIp
u4EtwrZme1FktgrxnTmTkkWrZQ/g/LHxIwax8f9+DxA8ZOzc99c2qk51vxmJRqEw
yoI7RNDincZB9xGnIyadJ+AcddC5xF/ncdoWPTGOJeFjacEm0V+fVm6TPMT1mCgb
eBnclBfunsl6T7Y4mtwXParvpzUU0Wq+pvsHWc+1H11/oPFT+7Z0EVoBN/oqDHhe
rEQcFO9LWfFDG0ZIUDadj0qluBF1gW8dThZ0T9sNa3pbKiNOuipT25uiojsefPYh
fcBtFTcrUm7JQagYF95q8WgyOnb3/TQnyAvK2iAc1KnP+VAPpA7d63bAalQI97/N
bD6z2Hystg/2br7/rIYndhg3pY9K0I3Qe1OrdlgxTMiIqZxYapPC9mcU25NMOjLX
BUPvXGoVU/5C3ScSpzgMyQDYqI02bnq/ncVjQZEt48IJpnq1T5xG+rtdf5O40OGH
cn2v4ojBq5jlE6j2NxWsBK2K5IBJfL4vqWvnPwhnnrIhqJq67ooTyu713/d5BB+3
A3hYhx0+OBVUdoOm8cIcbMoKQbTqg5RXOP9NFdg2g3VE0QCa3b+OnPCKbXSvvlbv
KgVJg/NIWmi5/YNncNaSf21zAlvtdVAhZKQMB04ZSrbRGrHGJlxWbd9zh2o1xrLq
qrpgoPyDkboB3xggN4V9HSn02s1rr0k3qJhqtMB/CGjAjrSWBiKlw7VHyeWqmboJ
uCyl3MFJCPD4GUVuEachTkGobAjBTreVh0RUmJxFLXSKQtvxgxGSO5zsybsQ91kx
GTssesBGkXmrw/bMYvZKNuBZMhRptgslaT9Es8IBwYTDOzhnDSI/iGVxFAIwj5GI
cGtOH/NZn6/Hm6xVS+QSh7AKu+EBO+03pnNEojiRIS7t0nM7IELmj7AnZqmEF7Ff
EHGZJZG3Mn1XydIT8YukdtBp+WyRW6v/loH+3eIqEEVTKYSRi/EN15ywRuqN9MXG
BYnpeXARXXx5wp8lsWVZ0rS8SAD9ItSvjvAHZoyWvyI+XY4r1mULqwoDr3vSBVj+
dyA/Va9l8CLYioc++ZZRLAP+fL8tODi4e6QKGlWAAipxzX7wqwaoE5xCHBoREeng
2/V+avClbwI2P0C0qitW9Q3ZvV81KSxfmbfIjqYq5GYFtfGYX1P0LuglY4idtVnZ
BLd9QUbXmj8RNJ3zEBwwvPXBQEaehFU/pw2YnM8Y71Dplu/nhqUnQ3qXr1vU0eFw
oTbWO+b0g5izReCtvXRts9LQzimqAk8t4a9+RyTZJsH36Ldl8FQSwr+szKQwcD0D
yJLto9TWOLYWyLY3sf1iSFYCT+JsahMNDpdkHs8TBT0PbFpWlk/tUHe2SNYVdlhd
j+he+vYViMGNmb6zgV2fNw8J0vvfV31ko6xchOSeQJXYnnjbIqCNskyt6MLm/ixS
152QPxwYWshUXPLw9GQlLuypOYv7ol0fq0QP2tflN25bIG83cESmLiwx+HfxrgKw
yKpf9R3bS3dHlrl6v8nbKwtL4TWw9Dsl0hbhf3tzYYcQnMVmuFQqXBmfqHUr5vuo
FvTMdfl7KIsqZsM1hjPSP6bm1xxby5NaICGkiLLiROdouLU4A06Pe59c/xhVKKkP
bBYr9q4TzHmNL7IU1VwbTbwXO7a3PZIxA1VXwOrebaQ4ZaB5ROoRTzPjPnIFcn5T
sAkgSKTuaJw6wZAUcnFZ/Dv24NDBLnZbspKdxYLqjjOSHqhkqpiDzomvH8eGqRHD
4Qc8Rb8zptsXAhTO6vhHzgbY7barivPbuOOOoiw0I9onFAnTqtmqrjiaSrxSzMzt
irYrSVpdbwKASTQB2Ul6aeSjjkbkBbiEa8PDAfzinwypOZVVOAqKQz9FhzMA6zkj
Foj3feYbUOD7wccajL/o1mARI/ZmWzXs5bOaVVfUtsjZwzENU6K9Btw9e0h+n61s
MUIJRcu6ORiZi+vMuoHM+OG5GNu+c8AR79nO3Um1YJRQBnlrneVSyerUqo4V5V7o
tmdsi/t45g6OuPflBAw2OzGiCmAJj7vPSetq6HHUxrKI9zY7JkLEGfi1ZGvwA8RW
K4czl3fNOpLOdtn5ThAeV9Y0eEevUv+D1gf19ezf+k3L2WOWIxUar34ZJIxORrVU
PBTE5CH0h0hPqO2AfGo9bC+x386o0VOoguOrVuk6Tsm8gMJP7PrzWzFQZm+bGaDk
ruwDAyZHAmM4KOnER6nH+Q0ZWDLNb3AxKaTc/Y9qUo5NrpWtcir3/iHfRmyLnEOo
FH/2+l9r4LXU5LY7cIecvRF52vpD7oJlHRN6KdUl5Hn4aPHwd8RyjEWIzubVVRHz
4tAsjWfkfevZzYO7e9Y7OJzeb+oRjW2mVgbo8hGcY9Ljc6/W8Pq54kLOMW+Ntbg8
jgBJDGhZlgruGQIZkswWBJg2/dhB/07JRaCl7JaIllQTE7WByH3QHklsPO706DM2
YDs6kjWss802KqZrFJNWIKqh+aHvrLSXjyrWq+P3nZ1+Q7UiVzILlBonmXCI46p8
tut+2vkuOhOka8R+P+us1nx8r5w3YN+16Q1oDBfbPwAFT0xtPHcEL6t49AqV3o8W
5bhlfGN99StrOZBGM/ecieq55D/FZmYITFAasBE+gCO6uUody3csq1IKfP4jG24o
9HvmIR6RTIO9FdMUknLEjpAJYOuS8UhH5rZXZRC0fYhvCiEpUfEjGDIRGJx/bqE9
gyI1aipWwEWf1P3RzMoomB0hKzXKkgKZku7vqTpVW+3XPnlhwe82eM/xYZVMCRhK
ZKEHW5VqSz98nAfUapcBRb+jriq/8+gG9Hjs8c0hDW8AL2AVmsS9e5qxVc5B22DF
pdFoE+ajbTFDEZVV74YQfY4nfHk+L+0Gx3XG3TIfedYRMcs7bFrXrW65s27dL/cY
oNIr+p1WBg/kCerCyFAtY14DhnRbZDRVus1glUT8yho/691PqH2++SjSO1eNXWo0
Rho24tSOE6xf8wWNEMZRWE3HpD1NtXmC09GETfX2wozRTMIgpfgSsbowz4xVNFeG
Wt+7nYRaYnET/c2+ByIHJg8/bXJ9qTSgmznCA7wMdVdBuscufIsDc8YIYCZkRaoR
0ZJ0yUkGeAV2+3rJKtCuTeqqexikOcOIAkZcwqZRlmJB9xGFs4aPmAN8HhVaeQiI
s97wd2vt0LUNMBrVJKMmTMFGt1XdTnnXU6wFgLMw1fG7tF7G8NUlesC9ZVqE27lu
BHbVTsCu3K0Cdr/zwtpXuT+NFPWR6LzLEdKURwgnxi0rtaLyxl/lGThmsH6kSEle
3PDwj0UPOLIBp41YHun3Y2BpQoAncDdpW5GBQuNUoUZ/IOlEOW6FtKWGm/g/VuwV
+F18eRYBraxP+FnHzEqisDjjEqjdIL0ZhHMK7M5PQOpXCYgAiJmeNyX6rM/cLDHh
g5MlpJcQc22ITF+H9RzjlxDZy2R72WTYAeldVCXHIqOf+X2QPz/zK9vbCiAvFz+O
+k+UmvraYs+nvFWq5IP9vaBWyZWexqAgVU7tuVZRvNHpZrbEJRe2rjQmTmOkHGB2
fYZ1adxQR/hYsz3CavXbmegnhgp++yAfdVHJ75J4nSGhVhWJEAV7c0b+9i1IiYPc
zhKPCY2lmkRp/gjzUd10MJCGvhsnZf/7XNa9HMV5l6GiabC34niDLYqFdIiZvPFT
Tn/RBocGvGqK7UxTesp3cM2YAV4X5psgwDU4zOLTEi2cmMKlPwtjjGGPX0ktIUGp
QxkCjhkOWx1lTkAqxEZ7J0ZAZ/fIAXaJ43Qns2Jlamogk6KGfPnmyIvzx7DEEcmo
xzV+mRbKUqIXPAeA2x2wiNV7mWoOttVzWETkFKUy5sMZYsNGJEMOFRSU0y8C8GKM
LyZH9BXuRvn0oRM87WmApzFgviEobzVRYC5OW/QTpzkFWw/oUjORUe7RX2OqhDlO
8PzgA3FzndwECK1MceMruHVcwymT8WnsOL+I6PGJNjlfgVhrMiT4KeyLw+8JRpcE
44d4+r81A5OaS7+n6ASGvS32DdOCeuFxFSIrg2lxTKzCxiKt3eqPyUKLrkuVT+An
y//R1056YR1WYUy/THQJMbVun5uOjg8MyMwGXKFepuKqleH6HvUf2aAp7utylaic
9IT0yLHKII5bZAwl/LcV133B9Ps1DIw6H46Qde2C1gBfC/+H8rMRi2SchK8s6TB0
GcFGhZ82/f0UTgiC28+bnHc03rayIjO4Rz3IryUjaBLvey9VjQWLvsVOZDZudtEW
fqg//4nzqWKed3zT0aHSuIBvilRARV1SCS6byX24xg6HiqswxEXqVWLQ8Lt4bXuF
S/sNFLOdD3HeErcDtxmcsE/EoZ+zWuv797dczOHGh/1Svrxatz1XzHUdLi4tWuKl
czJSrVvss0KyNYARYPw9ptV5eFPQ0c6RmFpbnpQ/pO34qIsuVS6r6b2dkWIpmPAn
c5SG4gucCwnzT43BmkMhyxvDULlBvl4Jdtpkwk1/iACQ1AUNBH2b7hrYgpEQODKl
B3Cbw34CdG6nlvF2fWIzsMd1Rp3PxZpJMxTt2Mxsq7hUuPo+f9QexBbZy3ST2yBV
6nW4xURckovf2J+YWE7T9aEKNTSkvPpnDaxmwnhGN/USXB+R4AJ4Tik6Ng0zorqz
A6Oz5xhIDcaRv+LU1y300RSNFoChCcf5kWldflqxIIzDakned+8Kh8fVZF5xkran
pUIoUEs2zywOtPQu+gWiq8zklrDLmLFg0dzOkJFL69wHjbfUfdr8M96dTvwQ26Is
KVxUoW8eobhKUxxXDb3CdVidxPgKW2K0AUaiwtr8hIBPO2i16Q8kTsgTmZtv4P3v
WrRVbkN728ecvZLED9fbyPygd+2ckDEnu/zoFJ2aSISLSwLP0pLg3Y5iqX1gkAYO
6kPTi2ZNvk2+2YgBDe4Y03CMWF36j31XdouQrS9YgUf2gpO+rUvTGsvpNSboFxf5
GvMCOyG9bQP7ToIJvV7aAg6b+ijHSD3DaZ8gGdH+tbLCTo+rdZC16VTsiCgBI0S3
hO5K/1SYu7yLYRsvi5bL5ljEsYDOR3wJ/fxtO7UL/NaPbwu+W1CYgAyQAMl4t/kE
P53jpZ2gL+rwicaXoOyN3nUlmQGIScZLlVQ4T2dxxxjIvQ18iFTB2EAsfOYCVDL8
FAI4wx3EWytgFg5QIfPvh9HNI5kiqlbmIq2vV2zXtMeSnBykcsPjU3HWylPz9UFt
dxEpICz2xtCGfU7wPXOprNLZxTdx/b5tVKaK5N14RqiyOW74XLVq/duhFb/XQftf
0TULlhZ0r1zwxUNG2PqOp0Qh0JZ0Lp/BfH1CGWOZgxjXl40+kjdmHLA5Qnsdw8FC
iXMqj7TJWvMHJbN13M8S2gA2Ar+g012xJLxJq4PiqYfdEUPjGISl0OhMLA2dt55s
PAFbMXRqendbXrlntU+k2KoYkZlHbpb8p0KIZfmGAxku/FgU8k793R3tUBNCFcc0
54mbk0WCUa/bTp63KTS1Exn0IoCb5wx+gZKc0Hf9bg5nRHM/Bokkh71p0XmiP0Y1
/KJCReNM7wMXHhqQklOuSrRyMhtjku/0KV9mGPkFhTeLDguZ1xuM63JuEd2fqJWx
E86/bQpgIKzRQUGCBB3F5NgqG8ZZl3Wmjt+h2wrF/Shh7LPVeJhZJfYFhrZpKG2t
isCjHy2m5ArtEPnPMxowkN7WvBhAgsqZ/ExSGTmgGtmnzHRxQRSi4mrkIPZj6GSn
sgr+xIjdCxYY5VAunUqtU4qfMB+39Y5X6wnj5R5gP6E8j2BVS8IfKnxlTGt9BKbz
xI4zO4ZKzNdWP3j7LLALNmxd/tuiK/tPO1zDFdG7Zocr8Tz31y0uQFhL8KHztt34
hOsvl0BnriiIPwLBu3NOsIqXb2WFRo7nS8dK3cAECrCLBngCrAlCK6F5Iq85nWwE
oLuuYTtzQdpHCM4fFEgETcbEJb/RSV5C9PqZ4EJjvTMYXKcy4kTLJAS7DSwwX+Bj
irtyb69FZM+IQ7CtE4hYgeskokTrB4ous6aKN2ADlFvoe7lSaDp4OthbW5GUtrPp
wOJI4mwgwfaS4gqviowwomHE61HGDNJCgw/1jq0siwv9xIlYtgu9ktXUzWtcoWdc
bxQfFQ2/1M1c0iXDqGrJYa+p3ksOnGc8d0kmMvue6f0lstT9cF7rUJ6W19nAykdQ
+gzc8WNaOLkbpexScu+zaiupgn2tfRfxS/+9GGRpF+aMVAMHkXpg8D9r49naS6x2
L/pCgarUgeuS1O7noGtk6m518x90AoHygiEJ4SeIL8tEdqz8GFqpZRU4wnsJE3GI
oehj0UE79RZWvZ2JL1bAsJ7Z4Dm1kG8eFYUTg5pgz3NlPATHSYBJxMFBwtH8wou9
k49q0SEKPDuQaIZSVMCn/MIPQZ/u9x1I1cNDEntU1TKfP9V6kZp/AX0gwUve9DZJ
vPQmo6KPbJmNRrz+Rzgtti3r3uwIWVKe/TZ2GZgO8sdhSDVrY0XU2KGABiiwPDgl
TpOuWhj+ctBBc7bw97Xk11LNKyDgA72rdRzZ17B68Q9q9RS2fTiO+gYlqG+de6Cm
/fLbR0KEHTlBaPZORp8ZbAdFmX/ZPNG1VRjt33iDmsg/94zDaTAQz6nE/LuQ3/LO
qJggF9sf3eeDY54LqprIkCbH76rjuZwZIq/O1xDLICNy22D5gTu/xPum3vEN01r0
q1mU18wxUe0ZxHng9uItPc0hg+Nen8JPdky1Sb+cw9QPWP/ktCItH+1PEa3ToAyA
3eIPZFS2mLMnyaxX4SirEtDqxd6kkEpCMEZR83NJE00b07qheXsZlazBiY5v8Dgl
BCih90V3+3GjaO/No8KfhIsGrAnjIMd0hOV2XH1g03+JhGyHz0QN8N/AQRwkYsx2
2VvrNIc/E3FM2JaHkRjXp9i80S1pnUS4k6e7ExkwVJ5e8DvhIatot4CJQG9EaFUx
JRVkHiUk+hpPUA63PVK+eBdLyu9UcdLQVAr+3BfyTeQ1FnnCw30/TxGrFrpselaa
NVQyBK8R9lUHxSYPAeSmU2g7CVNcirdWx9M+/J3G2CCWcXW42P/Dh4ee7zq34DR7
W2PFGWKcUn8Sbk/4eX8UciJs8goGe/eMOUUnLq6ABTP4QG2XpBem0Pd+Jzn2oBSo
Amcu+RQO0qA9/yLJn9wk7BGIE0ni3kQ8NyyhbraJB+SYVMtw5dVSan5WD2+A6jRe
fmpUqPNlLoli3y4lJXqZKStpNMVK1XsF8nDySq+ZNymXNJ59bgxHnHT2oy6HL8Ur
5Lz9N32VJvd4CehlW7vdDk36M05xMns80QlNJjEO1/+/MvDmV9UlSUFeKjlLTkxX
dW+0lXQE1c9Mr2b/LOQHkK0hdd1NoyEpQBZ/lRCAGjbW7/I3I3p/WzHiaABhu5r7
p+B3A+XVuGQh3kGgn7xfE4clnEUcFe1mGFvqKViLzS1MuSFeEmGzRTkOYysh4HTr
Af/SFTNhb/jeAfjCFR/9DLsXQIUeKeFx9NbnWq8jnvJwAxFRW69YJwO45FLosiMM
PBtxoOutNEe2x98PBp7/YKsJKk8Htzd7X8jzorUT6AgWr2rIysgUqLVZ7bpcPmxo
j2O6PkBpYY1Ycb9gi+81H1UvDqZwivtv3dYYy2kZ3a7XaAMPcXa46nHNspi8iwXA
rbT1fQNaF06XMOJGQtdrz4Rv7j0eoCDmZeoUpzdfZFN2CVdum8Dpv2OnCP2RhwiG
Bu7rmHo5QGVKkWUut0MZzmjkHAFAmUKgELmILpvpUug5+8fMOersJDCmoraMMAXz
UnAu3pBAPGsOsxV3pb40ewWk/2Bt3ho98PrR2oSObrKCwb2164THJMSwrn5ouqmC
ZNGsejo9MKBLS6BNU+btPsiXa9jzRk7B+b2pibsOC6ko6qZGCjxorxO4J48sfFex
++z33qOpABwCh8ghV+aQDlQZzHbXNm5uwJ6da3wakvy5iUlo7Fbjljf7d/iPGof6
VFXGQ5tJYmK3VSmqsD4CROFJ2XHVQnVqbG+PoxmbBtIynP69Zyqsf/k+7IQeS5gA
VpC8f5bM3LUMH4SudtPaNHf8J1JSmD20XAEs2kYKIbkBnrMYXEE2NU3fBUzbWn8M
e0aCtuJI0qhWIYmuud/hElO9t9or4uQ+seUJSgh9kt4cvHN4U+CKsQb4S8OQOzKu
sVLIE5X9BUaXOvVvIUEarsBFCgTVR8UabJYDOzIAbpAMxgZ0Ktep7mWl46L04j2P
50ixP58pgB5rMIiLZZ8+d5SNkP8B9pytxZ8kS3clU0I5rfXn7hfpBJulTznQ2SNY
jMDNh7TaYCuyTENK40tJHtp+S90gpmcypMwhb8Gk5aGIirTdEBZND33CpXEbt8qt
fh4Pv5TbdiobCMCRYQL/g2Wc7fZsbQydMQO1991Jd+emVc1ANQIDJlLACt4mG/E+
BBN7u1TkMVuuS+pknTVGbFC7Y1yadg661E4P+hOt8m/uIEeJNV8BOdf3ikaW9D8T
nOJLWpsRJPF62V2hH9Eyp65bqcsgdF9qhjiFAgYNsbUDlh3lG59aby+5X0JqD/xf
IPYMXmQqJkSMmwstCkoixTQ3W5KdmntFY+8fXdpEhji8H+3BswLhtpgGQ/8nAOHA
D5L4xa6vjUmZ+mEJhyRJyihlBW4eKZ3FQr/46PLmGStpatOqJLrB781+XVK/gjuo
NP3/NTM896+U1HHHIVXgkj6BHP/g7coVhTQKCfpGBqKLha6ASkrqEloKJMB6Frzy
DwQ6RnlTz5J+DEfaQb5ofw3AwiFjTaPp1hDXT3lQmBuh7RCgws6/gHy86lBkIOfj
Hh9zaqzapVMufIQ51aR0nQvgnY5Ka7k/nKnr+UdQDKBwOCekzq6nHDbjnpAXLfBe
WXNoHtpnOl7gV+5ptHRGUM7SLQSOeDFJZsUT+aWUirhO1AHL81KhCYPYof/bwxJ7
eO4mhtfqSmhwX0Bd5ssnz4w4Bo8oAZ7WF4br9ohp5Vwjg3omAJG7A+m1rexbreNN
A0If+j/ysskuljccMn0mkgz79WKHrpw3cvU2oC4LRanUZg1xjQuuqCw3n08dwTKm
vsjWT7WwVUGjdYoA4psslJyW9L95jvVFzpgdJePod4QY+UBfNCAjV9o7C4zYoKBJ
qG4FEayPJJrn9kQQZ7AvQTqLBRGiaHovYGRG66t/uV4y434JqhVvys2InI6zoiO7
BWkR9UQjK1bGPrgqYhC4AGhTE+1C2U0KTVkUO+mwv5ezdGXj10xo8ae7yLPRTQ35
DELAoKLO0ejraQ+9CibRKCBHBVvAvU/KX5cqHTgDGwiP/iXPNYthalagZv8yHwM8
M/4efMwroYyYhdrCt6Op/YXKOdv8HLIpm5+PUe9dmiFxQQWdIp4plnTEPR0EznHy
KetRa+gurimOpLrvYO3mHDPnM3lnyYBE/utDKsR6A4iko+wTr+60ISuy321tt4wo
gm/BjnVHZ7tHZSCiwt8E/d3ck8N/vw42O9Dz6xOaRiH6+c46a/fA+6Thnc2viYjh
5i1hbUuRgOAwCXH1pInfkpxx4kt7Wo6lcPTTEZuvSzEwy2sJSA47mfqDvniDUXUK
QLrcTkJYNrrY6WYLBhnAXzkGIi8ddvVigB4RhrW0uS84IhEpZ0ylOqShRGtYOPFj
WND3Sfy2f6OBpwGHn3MNQzYpO9JW4y+cVsbumpS79ND7RkhZFQHfhJSbKLUmoEvr
Q0QQIulLcAikRwJlKktGnIGgIlfVaxXObOKU+CROHr+eQFIrC7y3/xqr3AqCrRzo
HWaXodNa+Ywx3CPHvrPd2jPF1bO5+qmQVwhZ80PSSUkOGLkDXiEru8FJArk3l8m1
6zTKr/BA4fis4tv5wk1l4lt/VH8wuGfDX+HmTlpTE/52er3Wr9k6pQPTvWgXrULq
eKVXFxADQ8JTvsFODDeT43darguvkyuj+zXH91HHgIzRtkUiKkGqhrxHsurr2P5v
rE2cmsjbomrsh3dOAL+HTU1j6T7PdLrZ+oDW5nnVhWXlmAA6mpqKyGSX56KBUP9T
lxmw6KH5fvXlLnhtQaXfSZawPVxnhAR9a3VuJSFk0QGViJLIjKrbBZc4WsF6BXyf
fYBjqtY7e1MT/UW2p6zTGhY8J3/nMBfE4Y7JTHNZ1TSJK1X6lPZ7N2yQAHw2Sgvg
PWnJ6DJUPWwDELlCoMpHu3u5jSFIWepGvN+/RSHOdBv4bGMRqJ6uU6lswh/TJQO/
CWDsvYMpOWTfXP1RBTbrEseL9pRqmSTkc64MaSGZTHwN+AzJuf3Kl8xN6FwOTgHh
b4+vOrFl9Z+0xGXMqOBmfbcELAWma9FDuMNsjQCVpY61TMSZhDiPeMf46loaaWSY
n12eQ0YdWOa0R0LEYAExTls872cca3bXM9BODrGvlOxrD7qVI34Zgf/YlWt1bBLx
7kRHCI27mURmP3fQD6A+nQooua+C5x+0UDwhtrhoQD5bTDkzQOpM0fzVlqTH7WFa
fFZupQPKwBR7+cihb0OLj0oK/1cjw9aI82bz3CgyTraMQ2bhpXQlDpGdFmS2rcGA
xZ3WahvhtisBi/YrkxHhouHQs+0ZboVnN8aMqBnvw2uTyUhAno7HpIiGRZoGne0J
ZjQUgB83qCa2gjPOMJJH40DFnBfXr8++rSjciSJRBYbDWoZRdswonEpvTIOoWRYt
rCMfWorpuzsgSKy1T8a0hBrJonA1bXd2bcUO5AWjWC3NkcIZ5N1Ar+KLaYWYrBFL
zm8iQkG8qREhSbXiU06h8vuaMG38Gkfm6QUxZlcALx5BMqBpV0411otVa/KysSSk
CzU+QBytAJPST1xMftlaXjGHy4F3i5JGaiSzY259oJKt7Iu7TzA0Wy35wvy1+T7f
YKA8qyES21OxUi2pJbII2UQjEpsyVceJEAJm5ijo4R/5qOP+dOx1/8PrWt4zJWxO
IwrEHGIbe0TWw4Xvnp3Vz1BbhZKDGVEj2XpaLTAglamqgbhBTq2k6AJF1LX11r5r
v9w+r3ToZ54XZroYhPoyrORFtk1gv9VTm5G5qVGXlm9bf6Stbg6ONbdr+e4XCXCF
9lSaf05DBwNTeReyzkO2yTCu8M0c643VD1dEaLmtHlaW2DOclJ8sURelrGa96EVj
/o9XIvhIMibACistpk6TllpC6BIxXegNs+Mv3a7+rnx4z5utT32N6gyZ8c85aVwc
oiolm95xHjrKk+hcv/fS2KvmuzRDGqmxbvBdVDAGFv8OJzmazFSCkQYOR074Px80
hyf9Q60GPfurMRTi2Q9Tb2RoUXu/0VvuRg5mkQr5hlbYm7yTwtGYCX3JUy6qLSxb
fqfL+EHWIE0pi+Qhw36tUptYjFGNIcHeDLoW2vdHGS+iGBNTa9UBOe/92+LvAXRj
T2gIquKhyuNbks6KHMCfTgAzMqTNwJC55dDlVpDgHdGuuklaqkKQBYc219NVG5V+
JBr9O5Nrw6t0FpcqBExF2Tsqi3uuRE3FIjNUjj6yiIlqHDwb/IJL2tjvVWyJn5dw
myRQSDmSQjwtesico0WGGgx5X46cLmqNp8RVVEaa94xSdtebVx9zKrHn3wMFU0jN
l/a7O3c5TDNp8ROrZiBAq2joAC+kDq1TM+6QTaI902WQJZp7bo56GeNuroHH41z6
HXxWISYnrTQmOS/6yblEr1Y1lapNRWExccROqxXIe5n5oMxocqrQG0301eHd3DpK
3RnsSjOynhLfGkZSU/+6P57mDeGIqNOgDE729ur5R2YjDtL3NJmwRGAvcs6Ktb1G
VztJ3zTywZW0qmH4EnrFycibBI6Ln6P8qL3+EUF19pe5qJ5ziHjRLPjZEHrvqk4w
Z9ATlRkNJHZ54ZZ+opEjXBxowtbjFmbWZ3Hkl9dZdtZCLn+SrsOM447c7II9qSB6
5JmbRdGCETgCc33LZO25xV0daYA0FbDqj1S8V6LUjFwARRTw/MyAF09C8ImZlwc8
Nl5H80mCNkyCSbMAMl/3jU5uA+VgYpqRe7gTGrf7t0HbkCUEytK+WzLJ4ctIEU83
Xjnl/MltJBHYwUTcYCQ4mkJoUHxZ4XFBrGHKFLYDWWkZENBXJQjPaUmZhVXuGXwt
9K+KWOjOEw9sQGCl7N3gTAh4MiO43SiCgMQ80U+Er7iNGo7xxyqyAJdGVnSaLXLf
nh4he3xF028UKqnokeO13d5umXtBV95EPpXtp1DCcI0ECw0FwLmlaviGHNfFkGH1
Ru8sZSnoy0Rq2k17pwLraCNMMaT07miIeV/d2Ej0bKVC2GnnVDSkHhgMKwxwUgIp
29clffJl6HIu5DRrztHypOnHtsw0Y10zv5cTpMoYO8ASSDCQMrNLi1aptX2gzlf4
sbZqMXO8j4yFNVyhSV+snlOPguZD9D+6jhHbEMHdyCn4KmNihXJJT/1taVfeuq/c
rEghRLRe8YQGiafHj5j+/fcHoapWXdWk1PlWGz/+uDqOI+YeB34qnvNdE/DNccvX
GK9WWiW930UZ1SNsfrkKxZM8UAbJK1+T5dv/xTmMphpcKiD1bYpUSmUWyJD+33pz
VhMzYja9TiUxW0CUYorpkDp9GZjVhTiQaVkYSwBMKNteO/EUAXPg2vSmsgdSUJGe
KDzTtVguVFe8JK3M+UkanADf7Ph3CgoZ8F/ePLdArlE+b+5NDOigT0jaBu7PBJdg
a1HCo0N1Ace6vLI4AKqoWG7ByBGKGbFpYyOVmIhgzPshanMyQKC54oC15UPWXiNn
siCU0lRbNkXs00PGQ4YnDThItUZpkkLLWDF6SUb6AvCs/2+u4blB7023iLk/CNmL
2n9Ct+Z8h6lxjPogDT0dAawuJs+6epOLcx6gvwXsqVH2BoAZ6rGKNUTvLZWh3DYX
4Fxkef1m3JyMCYPi70Ci0nh5nox9q350FYnnCrrsyYP2TPuBWxrIaK6PTd2DAhpk
ZSDRWEbdZXHeSmOQeSrfuboOAA/Aw9NaAw6Uuy7wrtTN2ij2gbp4wit0q/QotFMI
ssjX7u0pLjJ+gCoW8DCRFBGTJBOyPEe/XD+R9gQWmBIpD9zsjNx1pkz80OIfiLHf
MM+dZ6TM0qfXI1+0/zApFUQz55qQT2albQjpWi2QQK7fVbgI4whAXpIpU+m0fhCM
2k3FzoG7JyhwVw8y9WstlfcaUcM/NiyDLlXx+2sc6Sl4tiefJQffYqOfWBoRUR8o
ZjBA/+kLdT1szEnVbU4o7YIt/BL+2rL7xaFUipSdnWTfF+Kd5g/ZcSxyMjqqEBSC
KKkkb5C4sl4nu9fI4oZu7HBfgspjavcjh4JqkZ+pNvESQYKKBhV2Akxad7jODLlO
MoqDf71sQUJlSl2p7bzMQWKA3iOlmPT7I+6y2DhxEK5oNnv8AjA5KSN0NYpEKSln
A/4Rcr8kL4sJ6+rTO/yAqdI3qtkmNmO04vMnc/e47yWlgCkSBOgEwJy+HnSlYssN
Md59JcQ1t7SSr0RqGWWJduhLmfh/pYU/t/8Yi0xlBwS8cyIhxPkVv5dGo165MCHP
dwkNSdf9/V4hX2+1j3rc5DKQqos9hNUNPWUnTKOYqBEadq1AgrfIpY6KbKCxtDLT
VjZcb9q6SwxJ4KleTuBsipUc2KNy+ov0gZJlCF7uRvMUgJLJh6VCH9tS0Oul5hyc
G/ge1ZstlJ3JGEwbB4ysQBHWoDnTuLhU+ZUd7eozEY7TOyKtcgnzhNfrP7emn+cZ
uSDARwnX6HBjAQttY4JSC7FfvqWDdExYXQj5qyurfrdFbINY2vWZaXrR/P9Pxzs0
79PaIuG2zuAFm1hYS/WQ4ZEBNhmXcEaCykxjDcEqVfE0idgjW8r2fPWjj0SxDvkj
k1Vklj05VlSK1B0EkQlvdEJObj7QkaGZaeO7WnYbWTwTr19LQfz/wT9WOF7adRih
HPXSIXJMZORLXEFLDmS+je6Vtk59AZIlM79rsbfopCAgIeex7tLmzkYyf2xohkNP
dMpPmfEDaFbOJvG9DjWRB9Y5BYuK3C5Fb5Nf+3jqZt/dyvYcM8Lg7B2sFvsWOpub
G9aIKFVbJddOI+Iwd3gcwjXOiuLgFrF59lvFvD3ktN//J7LYxTLsuKVc5VjueVVg
y60ypMBYaRD3PwjkjOY1zeVftovwfrzq1TXb01DwYeHWvTpMtrXr4XVSrU4p5Raa
Rx7NGPDEmyx5fJgaSqXWkMyaS18hTzZNlWjpwnAjUMbjZSaGbBBvKzO76FPNZN0Z
WGKgjO1Y26J6CDcuTg7Pu3H5Hrs+5UCn7nj1EYtnQ0pgAOaSBzASE4lKyi57m3gN
YV4Ki8jPl5tB+18E/oA8zYcqyLaYsEVn25SjMtQT8KqbX0h5+r3GkyUuLK9WE3N0
IvFd8rs52QHNBl8aKu1yFKp2PXyfc9Uj286faSifI8prOJE5O2r6Ll/xToZVPApR
PxSA4kyOrqxn6OHOr7fFQ1lI01O4TiD6cvnzucECuKUQYO8uLi5OT83TK6ZGoWEm
Lx3GqIG8eZAXOgNcGWSf2y1O5s9q8Sul0iW7GKoK6Q7EGC/l3pO0HQuXV3QOltRL
kfjM4ilVVn8YE7K1tuIbfdtyKOMd95XVxjCtMVPo8Kf3ZZQ2rsoGk1vquZeXLGud
e38qsLgps1XKRKl8V2DrTlgNvG7cWsiGACawkZzt+0F2jsp7i7+VFMs/KkGOmVd/
LPegI0R/fdQ6mRJ1jeMO9hzO2UJljet0jao1gRBDv9O7OLkEL7XNkWgAFVoHyBHT
QHxMtkN44qEYeRVVuWaKnu4YzSOUcXIWeTT8KTXBsGA67VjTdgnhK0cshbWCqTbO
FaAa/OUgQDtupDjGD34l7CHf+xq9N3nP3QBE1PTDCZ4iPPzdXQscHkioze7V+9w8
+M1wBuR8WUEetNmsPhSCpGNkNU17PBi+fGyo4HP8/YMdgUA8EwoLzy0GXjQHnV/e
iDAzYvR4lpG8nlEfqSAL8shCFMarZQokmpTGkI88XpD+j13Bk40ikqurTwUelzTR
Lx1GKmdT0p9/w+tjl9KN5rH4hy0JZINtvxWIxCEsbB+eRUCAn02iYpmPDQvZHt72
F1wHNsX0pqy464HWEMFpkh2hYCrqRjedm3pvfnB77LJPFzWPeiPeArg9CCNk/pMp
YN3BquEISA2RtwXXk+2pWHBVGzZ3PwSuicBtHz7G3YtQRcQ+IkrNbWIaAZFUVbg7
FS22PqWS8DlkQiVRfARhESjER76gxrZUYm8Ks9UXvO/ZnL6m67A5aooD/RcQzrJI
Opz51UbTpEBzT5OxuntE3nH+Roo7u1MG2qjYTYkFa8RVkqLEsKUlLlxRnXMxGuQM
gj0pVzrwB8Z3KFnVm3HPgno/mdxBrkMP35BvxZRg5M4EmMzDhok9XBgRsPaAEJNW
1vDtb5z4mkcccw0ORhLQ5s8qPMhkwNwThdecVn9JSZRBJxr2MJ/nhO6aJsVSVi5Z
lp5bBQajq2rrtG82vIQbjGF3TNGtpTUpw3tBSF99NTSzd3TzvuWyoSV9VAYC4lLg
AEH93697OiQFrSPUsITC+s/j1gOOJ4s4t7NWGzIXin4Z1cGBLt53pfnlmcOnmkqd
Q3ITZDmUipLMP31BToTBOPlPlAzhKPa6uBU4vMRVlX0W+ERxE6Bid4ofK2JbKLBs
s/dq6c+q4fX8MSchWSVuotcShybDMblE8uEibU0m1Utv1PvzwxcPvgukwKGLR8kG
UNoBr/Cww0/bkC+JLCmCwqkbfnt8uioM25UMdKG5qiesejyaXBVR47MQfwgLxwOi
TQ2lyWgpdSawzeeeWq4azCGUwGUzyJ6nc2L8S05hTlMbnZeh5qiyHwSrsOT1nU0s
YCQVdUnuIRKDPyY9hCG6l3fLKRC5HpX2F9BYjmkG3TVE0zl9TAxfc5bv8le3Ed3e
dEkXV2Rh6iofazJDoZP6c7hKOVzD8ADu/WfiQnchNQBPsjbaywf3h4NkkCI+vgul
xBL7/sIFZLomxLm0KWro0DfKRhTg4Nd3pTbVmOI4Y+KbZ4GEFXqltmezTaww+UpZ
6pgJX2qdAdTWjqHEgMwj8nhI6BLfWn9UXPMSdOEJ2ZbUJnN3fb+JFM9hklWR98DW
LuMIBJ0CfKtnO7FIGQxJB9BJbBA9ueIKWi+aNKHx2bk1ZjGzpMkACm86Hh0HXWJG
mHxVx6aiqbdAnQDKqEnYuY7RSnG+80oq5nJcsRVMHZ0JRry+7dEh3pKTTJKgOn4f
YZ30Kd1v5/WpxtQEZoqL3ojFmc51fApSwpHn0WvFU8reTyTOuhS9F5STH7CVawap
86m0AsZZhgx62Osb2LNZGO+vQ3hO59int3vCXCPVLhB0ACl5w9U5MdWG8+i8/v4O
`protect end_protected