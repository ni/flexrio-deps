`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3792 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
/8dei0SfYi/yIzInIePi3GRf1DR12S5iBhzwyB1gvHQdV5qGSqgw8u0Gkc4vcSAA
fJ4mnK2I9RCcYat4515VjU1ZAT2uHO2Jx9O1r+5SUfTOdJIV1LPPxohF+wdsBI6R
lk3xghdPILCXgjGcSKR1CMEPd47qP/7Pm0jmtnHiFVdnM+C7boDvf+krJmP21T8g
fWA0JjSbXKyjXRCKdn+8P2CLZa81VhhGStM/GALy+1whDCnE24yOLf+P4gI9yq8z
u7KJFJhnjfnpHJnJ0QKgxMLRKgXKnaGqL2FMcp8+MQueGFewlYQRLFg4dXFIK7we
Cmhsq/8apO2+GsynRb7M39aBv2+bpWk5iXOZ/n/CljfdIOjUs9rPPaOjk4/SMHrh
dBYHv93eLDjG305mmz3A0NgyMGX1y3tPl6mnduqtZWQl9aTof05KYrnZXYMUAzrZ
JvnoQVKs60WcJJtC8jZQN/mPnQDgIX5Y4Q881wWScwN+P+k7dCBIDrn0xgJb8gB5
2Cyb19Ar7L8cZTU/Lz+L12dymjJVG+wueKiyiY+dRMOvXWeInMtNnkwR0WzbSH1A
7a6Z9BIOJMw7hABh4CmZVRjdb2xesymq/X1yi8Iv7PgowEU5c1YAChG0Jc0QBV8p
/5g4wwo1DwrqvB7pi+VL2dZ7XOkaKiwI+49K0jvYVvv+JrKyOZykvUKimLo4IRPp
Xah/n81WVPmn3APvIB4YtuqX84jGhSrSAObuykzddBtepbSRRn7ayyv5Mxg86W+t
Hfe1eHR+/XO0DfoyRnvr4vEbTJl+kvDQYXA9S7oLLFjN+nAFSYmCohhFRUHGjZKV
etHCTv4kcd4r4JW6PQLj4pq5rgQE6YwpYXwv7Y1esP7L80B6aG9UWBI6wHfAlRyz
BiByg8lAf2/DpzXn3regu81RCEV2Wp0JzrCDLGcWLSjn+4fYVoXUyFtpPGdKsS+D
kAIaVim0AOC+ohNoVbS4TcaxqGLP97xQJiWdQ/EOyjx/lBhJ1tzdC5ur6EeHoBr8
n8tZM81OHFRlB3UaBhu/FjjA9WICY0IzVksnuDjx0ttIL0e+IwEwb5n0Cxser1PM
ues4Oip1tS0FPjhanSDf59Xg3ARUcY9frsM2sqUcaCflQOHV9R8m64tkFlYQozs5
LXKH5+56DV3YHaZ/IQ4Q8cLL+DsBQUEJ4nNOutGbf7L+TZA6VT3KXgV83R/cYf/v
3v/jSkmGz0lvhVIOd2f21I/Uva6UIjRCgW2yf3yvaFiEaFWjUsx90WbeqLi8GQvV
aeD9zPXYzEVtbdsh3uXo7AFFrv6ZYYdg8PbarzKgSEUlG4rYixHK5BH1KVq8O36r
BW6aV8o8LlgjVOw5hac1bZeB/dmlRw4np/8wbkAZjg/tdxYmLx/Ds8vbHW6+DGE+
kgojLiRTr6uaUTQGSGl3BAhwNlZUwodUpgvn3eTVL0li19Ng4zwskom4/J7iDX/s
3fdVLg/Lg4gCpIyDiOhUK1Lidt8yDt74UfdmGd6AGz5eHxGZ3mvMASNNyPoEXZZC
0/eRz9rdx4U3oVrK3HHNKlUWERRPKaOtmpmBMtUN6jy0LACnYOhqYudn5L0lsIEy
QzEsTTAclDqfeODRzoJUD0HoredpqqUqTyj7de5maog9wxegu40EgZ7x1ekfJh4r
+Wi/uMQgqqb/IRWoPsLizCWz/X3cvio9z7LLZkf4svjt1WV+ZABuUr0fnv1zNo/E
MA6ZuZgrYCOfnjq4h8cWPpbGY0lCXPxiDUVoqwUdKOl2K+jbT1oSyOCIr4fQpRni
ltLF5i9DBde4qD2ghATiUTDQezC42DDPjKwiqBdAzxbYd9ESsbcKzc8OEcDBCE60
CH8aQ0sn17y4gfZx7svts7JLyM/1I7ANfgLtSvEphlnU8NBhstjm3oUASbdfhyQB
oFtRCBTib6W9GWpn0BXId9ugoERKfMd4Sp8POD87ZeySO+sH0mzE8+7t9LHamLF/
7tuWz2vODGc7yXBQADzDUPnoP2/UB7gQVwZuJ/OyTlInYrmEhGzQNdNVdajiu+rU
M/paLtjEA8cWN9eu/K+sChTosGQDmMuMK0E24YieMSl4PpFwsnzJTQ+fYTbpaqvY
ctWtKdcf1cB2l0m2Ej8YlorzPPhsRMusX8iCQZ6frG0yAAnUwDyrzFC3v6NdXrmj
gnkvC6BAyvAxxRulM6osIwTDQhft8sPiQ1pFfq3ClfeFLCRSf/jEZDa1FuFzrqLK
9c5WPzPGCWX2QS3WucJhdSvrMnOu3rbRc0owsAdJkWAQH8/scfDMmsjK/lmVzvW3
I/MMbTrjNDTPoo7xgFhVr/d/NJGujTeCYAKyeiZzv1Q3F+5nQh/CDzetRVp4b07e
JaU1a4+naMPhH2eCCjRtEqXhEVwLs1MtJE0EqMHP1MqCQeaMVva5OmuzdZvumKLL
RJY4SjuMSqQZ6L6XA0P8GkkE4/zmCfd4A3/cY9e2GSwskqIq4tH76dIWwbT9oE4v
ibhOdqUBfoqukuJNLj+BvgqnrWMvv/t7GVdhYoajOUiberyZcempe9I0VyxO3Rt/
7dAuoTf6ixZ/Y7YOuwYmLEXBSrdtqLjOCdjyPpfa7rdXx0uJ3pzss0BbFPkBVmCt
i7SNpqJ8oKl3teQ5aNvcbJ5jQd3NFbSTB3woMuNr7ugGOdbs8LriJ1phjgWaLkE0
iMIOjmb1gLkOdzFgWDsmCWhq0ZrjFfk23mAspp8vQIRltG8Y7pZWvUd3QKwUOpif
PEyMPavbgfDgtOF7WGFKSDhcyGcIOuRqO3GUlOaCvf2ST01a1GUP2IR4gFSnCbiX
QyfFb25DDOE5x0E3+Kf7a3NmyZRStvPjA2cxC42/F5JLk5bcoOx9XwehCT9B4Lxm
oob3ohYLW2tzQn4qzyd0LT5gXLyMefUkqgHju9omRGYqD5uumfBkQ2aR+kjMk3Xm
IDiOKjuuS4gHlEITg+qpaC07OZX084NZocEFEWaSOZr7dJm+BHskateauYpqPJ57
x6Wv3uHtfYRecxcxJ8SeyMXE+36pk5c0rbQl4uGnM08hvJMdS+KpAWT1dxlFEP7a
V8ZKb9mEG+7Der7vBfhdroOqS1EBRHoQ49n0Nnsyx9jSIvYX4z0eGYp1nqPoQwZZ
2IflRoloOcqTUxIgcuD7wuadkosGc4Ve7BVsu4h9Y3R/LvjkE0p4bmZMPdpD5cIq
sl1gp6GLTVjMrMOKt2us45zH7ufl2Xh1SJdBDHJIL2sT4/bV4m6g0cZHA4T0DXH9
3xeZ7O4WJNH6Gv3+ppsbZbAqARSY72R4DJZRt7pQVZtSVVzBGEtPfmBa4+HI181l
IDSZbyqdD+DL9npuZewOltgjcLek7eQArqOOX6BFF5W0Q6ddQ7B62cKoTmsCYaZf
qpViRhnzpZ+oniZJJ6zlHHOaBvJwelq0O82npgW1sMziG4gGwP32TUSVYDwzzI8Y
Rxe5LJejRmnZ3CcdOW3pmweAcT1tOWmLSkoff/UGPpnkNG8U8Ok9Lu22/4YMqEZQ
Y2/6smaVdIzPBU4X/DJqsIRDixTvWIrLfJzjF2UXqXN3EklxEiZDmmknkohbJobW
RGdyi12G0ze6V5gygJtaqJrCZrgD7x3yaTOQj3Mr262Z0mpngMG3BWvlrwhj22zu
ElFc0jXvHt8Wqbq7RJLQJvvbPMRJ3JaltSRTvU8aWQ4PS4VlMgRl0N6KfK8ZVFuu
TWLtxG6LLnRf5XEmmyQsHmirSgNLCRHgB4mcFqkMkTpg4x5OLv+p76gxhlNu+6Lc
THe3O+94lGzEpfkWDZXwV7akT7RGMMyl8c73tY9BCLl5zlPMfb08jsBev1PkXThj
7tSydlZk8fERdnBcNRDTqmMxWNCj4EN288asqLsx/tnE0pjgeW838iDC95hViApx
mSJxgbCDRFTaOY/avQwXAfHT80/l6yBst4knZss4r4Ob0Ld7CT1ozIwBDDadLcP7
McXpOEExx6m+Rn8kqhBubkO6OtYsMlUxGC6PhatdQ71JraNnv3B3TBnBIUN0R9WT
2oKgiCUHw1NtMzQ42oQJMq/cgON9YyCQY6e7hftEeW4aK8RwOttUncyCKZRyf3IB
VPwksMFQxZc26SUvgYSZlaZVOUCaR2//Y6OGTGj/V54/d5fb5Bl9D4yYbZYsG9jS
U6LhWRPHsE4F4z4XLxzakWJvPTOvS/sHs6FKdo67mTBVu6lrgWrJ1XVW4q3sOVL8
N2TAqtwZeL4MmEzB5E8so5mz7EfYTZqoXwQ7nf7zgIWAcjLtlUmCxEYdcAPIah4S
iTnQC9NKmuQDI3IK/tDpS0U0Z66ybDyJMc0lV8HqIfN55DGzEPNhXO/mLAO5wlpN
6KrQjbUyT1GehAEQz1/u6rH+KUgygLo4kEv/HnBDJYezSoI45R3Qzgzf9gNz/MgB
XIt6AfFhgCrMJ8PErVG8SgahQMidF5HTOCfs1Z/C4yIBq2qb6qsID3J3PAaWfF4X
zFskhytNaDMySgjOWdZrIgSPoFNJ3PeZaOifhkvwtQaf+3qOntFp7OVVRVdYURoX
oCexYVtUy/9EJHbtz4bpRNAGIE0wPg53EwJDyg46EirWX/KXm0WArbVSixLI97FR
mQEr2BA1TdPQ+bvLPTwr7C8CiuZcVSVMEIe/k2DEqtvKC+tCfXRYKpsL7TPqDKHo
BQOn8TAovnc8vDe48CtGM13hALDv1vkKgyl3hZ3P8Z8c8MjNWd3NI+Y+FKRe/FUf
FadTuQ0ARxlA5z91xMaD6PRHIbGm5CNlJ9psrBxd8oQINHxM0RJmHrFAJawA+GuZ
XEgScIh2CCpnLWPH2evJ+0w85PdUaXzNQvxUFqBRv3cUWvBvl4KeDw+sMj3ZI5sP
uEBKqPWFaB6i2nGMBA5+RDXDidmumM8V7RYGyzRjg+RpO5G5hOvdletDggWjotB3
`protect end_protected