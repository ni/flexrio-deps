`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
UKzXfYv8932Mhcp+dmcD93amxTkhcxpwxQoqNvi2YhIzQmkENyBKAIklly5f6fTy
7++XJWjS2aywC+oSuyxvqGfT2h6oG9P4Wl33sfFb8vRlsA/nmbTlt+kBGmxy3rdC
CIlqv5HINZR+88i+1hSteV7u5eSJjDlq2tvUa6WzLdUwEu6iiW+3EX4w5ea2p2of
lVzbfy1aY5JzPnVJQLigRrcUHRbL74D8vPV13ezJ10bpPJmGsQyXjLOa5GcSevxr
7unHhTOqIPbUJfA3uPf2iQte0R6oGtxF7fmMJhe85Np9fmNdk5bQfvT8YvRrs3cG
Sfezkw0136aXF1SntdMmOw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="112ecapgN9pzpN4gHWAzyJUdO7PtuCDt4rfEVPJL548="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
aWtRfF2b5RIh1i1BXGC0HQOpX7IAULFLGNvkPj/vx8wLomfTLhhwRG9C0fXwam5Z
rCo7JEM6N0RKHB+gz1A8FTeZEy5xZuHAarI9X4o9yU9dBBylvukO9x7a8ZciPGZA
Sd0Wc3EFPmoIwPBnTen+RDBoGObKAKfjxVMrv47c+u0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="MHOhLaSLSz/D1OgJwNK8PCknAYeGDTLC9rXJQL0V7pI="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8672 )
`protect data_block
LUp9g67y64XfIYMkbq5U3apMoFreNwLwu9k9qDQg67PQWN83Dg6JEsV++Tykh7/7
JPxKe6AV/r5lct3dNEXgFfMsk7CzPzqlYgipiKxw15mB2uekshVPAYztICMOcyYx
rOb1pYZSKbjpMywBB40GRukXvXlqy9wFYzVV/1M8ArffFuNpvgl6KWmwBcbuLKhf
35GgFfI0WxEEeEcYUwXxYj7zS/Le6lZe5ndeWPjljqXH4/2EsILj35W5iMx1TLCj
WyuL0AypK/xiaIi7Z8NywL63Lik6T2mtDB5jVyKjOCMM2GPrkin4HJ8mx/zJvvMh
mOaTdblxEyF1Rdpa9ggnnbdr856e61bWJ2cEv75U95B98sLotHxDEhDJpHyHMtyT
QATW8ylJV4NwfrD7F7LfDugwAjvd6dXowMQp1vKotpOwiRzljl/OGJUblJQd5KCB
jhtVBqQW/1+/5LHEhNY2n98dnEp/k1g2RK8/zYnmvZqIWB9+HZfnM4W+PqnYuZBw
OKs6WAIJy82uShaLtRr/unlSH6zDNBbaMPMQyVzA+e2HlVw9Z9YSYcaL8sQFTFyX
l3fSmv6j092wcZqREHlJ3Wu1lOfFh5Mr9pfCQW2M6WbIO4I3EB9/Z6FvsUm5ai5I
KhVurH/ohc05sF9AKbPzob25nDtbbVVUU/klYn3ZYE6CZTQ94f9Pxhm+9+GNqBfR
jDQjYe0Cj9vyi3k3ZIdIFGBL3AkZoKDBub0Y1jcA99MQ5IdHRCJrl25pZD0/HerQ
UYmpQwcvBqxf5EM+8MmSxFORMDG41yMPL4kx+0PhuXRxzGVCm1ltHVbpXS5kauPd
1QiBh6QG2/UZ4mW31MwS/szYazUNo0pAFnnyQptm2d2+m7dgv7V+695bZbV71FU9
9hr4XWxUaRJmx4w8Ik4ym7iDGmLoI4KF8/Fs3RTWS9jQYfdvIzOh+xmhplE7+Wbn
5PoR8M5wH7t0K4GQYd5JSRGKH+vaRsxqsvV4kJ2plF9pF9CWscI7JTto4nZqrZ0+
yXbO+6WyUBqfuxhrnBbl05Fn1oHgYEcqnBeVxymYya9lSiSeSBxpSmqNdx68/2dj
3GwiOl3ZPFoPoo+gfzPoAZeuHW3UcefYhTo4lI5nMDJHIc1U+oDUrDqUkj0/SlES
d7bDtODY1foIsADzw33I/Z9M1LqBZiBVqY2TJyf8SHaj4hD/qwbn+a7uuuYKcv3z
rYK3wj0JXKz75bSHLqoZUfIQNjtpjRE3cNJuKHfg5hci86BD3Pnsc2LJ9CUtruOT
DFCugcxRWCTiUnIoJBsNtEQCzjFSJHK5qKo9G9T37NRZLHCWJEtJzFoqDNSml6eo
eyHnK2XsqCpBkQvnzQGReiXW1Kyna7/fwq4xuoOYEqMC5VKpjF1dMWvwtCVyutNo
bIzMI2TNWuuFnHKd7ShftclAzs5UckfI7IqWvdaKmCE0VJzATykgXkdkjN4MOwcI
v2zXjP0cuDlGJbXnSwgmByLfd+vlujLa/jwkMiMmuKkF6xNGJjkWnTXrNLJx10hj
Oj7gco/DpFdDxfNolHtDgIa/4tbtoVwbkhSQBnm8gbYihdRqRw9/6cakesoEDOHe
KVwZBxbQwKAYsH04RY+b1QOglA0Z+AuOd5Q0OhqH4uoL7E8SiuvSFRkkGQ1XRPlV
EsNbZwK0xfzzPVc6UmnB6/dtvyd2+0hXwYo29ReS1JHPP8dhqXMrz0ovsKLHaAK+
Tf++gtEWJ85N8Eya9caPzyW/khxmxzgIuj5L6fF0FCMLC8yDHtooKVlFJlM3XNRW
2NJq3wZIWMTVRP5Jajz1teVhECQ3+odnWTSnihFOBd9EoxOTdWGBF+LlNX7nhvli
9v4qP0gwsKAmAsizFZuJh5DsCZIb4YcC06lX9Smj69Ro8uqo9JdB40749T6J3tBQ
aCub/K0uhH7qAbdsgb02A1IqCw2Hdnn5qRzUpfKOIFvsoottYtIdbaWaQdwKNaxC
ARBVgzO0XXB0zbd6TerE7BjwUlkYBvZJ9/NAVGEMpJfZIBeruZ29IhW0ONUePblE
ERy9E2PVrBFX7WfyMrd0XNup4AJUMP09hwAWwg7VmN0wXMpKBMRpn9eQZNz1yMlG
HbBYyMK+e9bHvGXw7zQZh5+tjRtt3lLETxJkxRxJUscNK0QN2c4I/XZF2et0x/uL
/JqbHzz137K8EvusccFV22KOF0cCJtgPCIpMmh4HnzWazfUJAYeuKtvZXnIGbwKd
DOjijHsvaos0duW5lf7FtaOaM88l3k5749vN4gFC8c1Q6JAOVnfu6LITnn6vYQIW
AYDHd/c8EuFYwfQohSMRNWLE10UK1Ta4zNCF/rRpcFtSU4Gfqdch1TcU++7lZJ9D
1+rtOL9Mg9syzwm4V6Ek83jn1fvCSt2lSpNqfqpHZCR6LqR27IFBiKjl8UKt6b+l
KmzzcDYT64xqPgzfURUJe9VKyuRwjj4TGWd6XQ+j0wGKYVc5YavoF5CtKcGcGA7M
9tHF2flqCmG67HM1V3LX+4Lu9t43CPLfZwfrk9z/a8fvSPn0y/pmvMp/mwIRvZcP
QVqYUqQG4FmW/X12kt58WBNjMgbF4S07aXdbXz5yHeZrlcfS2S5ku5h6VK2hyWIF
7LGxLhHgdjdhnAwNDFJ2ld2k9WjBHK6BON43HJl5Q4Ji5Ulf9BvSv0gcEm5yq7Kv
NLQChk+B1PUAxjjBQ78ippiwPBkM1HpkeeU97xYQxgs7AM5nZU9h657M2jME2+Xo
lMxOozvy4wkStzmTgui+1W41f1e6oHy2/1cjkMB3XDVlueEzfCMhHfz8uSgPTkNK
aNN4fSFez5/lU34xG614fQw/NukVFUEnPuhaJwopbJcKF8yMN4LVXiNbngAPvXPY
F2H5E89SCbyewteC+U8NS95buSRdLqClrFRsDmEpiy1bgqB+ZGiyTU1PhH7rOa28
bknsev0InEko2YCLW3tMofoaK9ayqIuKL/Wy0tzG7cZVGiSByzB8jFc+KBJiIQ2y
d9rgrp/2MO/qWDXmYXQnRqqIeXL6XT/o4zIMsAip2intYNGO2lpuk6ItBbXa6vP1
clljN2NCfDMDBh/NdTsJs3zvzO0ErXQUsAZi2iy53NVhE7yV5kqKS0FAwNpl2J86
412RUCECsZRkA4rz98RRD/YYpY0bjRl1XsckK9tmVMlc1qBW/gpQWNJaozx2nGS2
BgCKp5zMKiUQ2OmdAkDisnO8alwXeqoZ1o6v25A/Y1w2ifR1Z1YDLCe2RqLZ8u4A
vQgetB+joYoJgt4bVCoVxO/lOXzQEsk6H4ptlbjulm6XiDc8owEAGU31wP6EIC7k
d1O4UtwDK89dTLyZg6KLgDSsZgNV7AQmnl+d/2U0cxWpM6Zv8xaUcIVJ84frTNya
Ef/BFk9PzLTBx2EjxRdU7IQ3sk/sFKxfITP9gtPvpkp2i9777h6TGE6wBZc3dHVT
BpsUPyreVfWmTLmAiXA28xWUpPkOghNOg53+IwlJP8o+LOQQDLH0TDNqxxDmjg5X
SOjczRXBojowGCWOemdt73FkdMRcPZtxABV2KDGMQ6oaPli4L7PvrF+bFszU9vXI
zqLSSbudM1/C+EBcB2EMhrrgAzPrL/MmtsJrGXiZHsldTcfTzYf6plyj5NBBn/cA
e5NI7UNHlmsAY/Fp3AekEBtggwzTObRlQsSTa7wvIQt9n4XEkgDDi3rmZDzHKG4I
2sBHNDMi6jNu4/Rgo80OYS7+aKCSqsFFhG2B4O76h/4xnMQEvVkAVatEdq0lg1rd
daSfzknr3XUEcpHJd0Hn+/H9QanlLIDjpNyPs1HYU9lzeK8gvr0+ehc8SA8YVv5o
Il/JgLj/aojhI1LksNol9u5miEzLHtGF+GyYOhjRMYMtoPYJTBzB3ER6WGf1HiwC
E5HUdy8phntAtgPldLebLGeeq6H6jvqzoN932w4XHgfdkLsSEpG40NBVMx4fMyj2
e8kFnRL3RBNOHYxi45kc86b2P/tWTlDU41wk2f3VgYCiNi72QHsxLF0aYNRwN7Zu
G3mJny9LwiHbN01PbEI4LU8gy1hE8xiFKlW/M//jFHH74tV4gUwTWrBVB8OQzvym
rjDFwiXKJdW+X/hxEE096gMrLe76QrzcP21a8BYkTel9+48lQAo9bOtPWSTdtfrg
mb6sxzaduy31ZLGnsUh+VCpw2AeXExmeqALKceZbqY/8ZoymxYT6lVxswVXac5iN
1/6C73cU70wiHeQRtdhQv52jNMBnhaILCJRH4JQLDQatiyz7QHqY4+LfB3DWwX2l
JDYmtNF0Xcg9/jWNWejDN1suyLh74JuBgQLIsZ2qYdES1MCOb/9OkaTA6gMW51MV
In8YMfLJotlsNVObVGFXRD7TIR/E68vJm1z7OqhPMzgmy7g4/oy70kNYDrd0ixoM
ZpWZoRLBpJFgftyggWu2cvsPKOySQkto/RfmMoC2Bp/taVaaVKjlUVjG8CDAgyMt
PJvoXZV4LWk3txmFmfNMKrjLdJ3LEOePeDnP0OorGy6oTgHIXwBqETp2HOOcG0af
4xAMbK3M7+C4N6aklxNwoJF8UUfe0hiEQSPtYrmLepd960+hZNvwZeZJl0fG9zMF
XocTUY4B1oCZJxani1JzUFeKp7iMQmHzy89SvvUIXORPKXkxeiKQH18ABqWmDiIO
2Wd9ZRqmwd6wOJqTCoNHriwYpDzcu1YLkIYUUQM4KeT5ybkD2lefaIwi51xuPpNb
EBTK/baupZIxCbUi37dVAy9zVBlTZ2Z8RZTVrZDVksIo8YFR/3yC/qR8x3X9ewOH
Ks4/N38SBszM60ptgiCuwxfKmDgTWEv28LhasuLza+uf1+3FoOPxj4UQgIK61QxR
1pnwCn971ZnFLJG/H0+X3Uwlnbv+vnxRuxDpmKlrS7/5XocoltqDTqpX1mCoX6GJ
xHGHlIvHkoyv/bAsOxQIjTfls8Zs2IKTtUT4QSYTJrJwKpNto62nxA7GkKEgyQgG
MK6J4e5o1Y2ar5twLnihBI45IzSXuxu3bFY86JGRcZ1bpYrPWsgQudex8htl4J0r
fFn1mIXmjwB5qWyzSRwNKUtwbJMaOZxc1sXD0pt+nXRgrYenbNy3NpLbaWt46Dyy
SBW2nqSCc9dzrscQnh28DDK9ddCOri5+7dlYgHgbNigWo1nBgmGR1HU/BCDkVJf1
frdImXnflbE1E/e/VJAnNoktaxbJuKnio/rPZmEZNUkPwcyBsPvZNdqZdezxXjXn
fnbiRfQu+EHoZTx1pWgW1uH1klB2GMU5F7DT/bcnHYfxI2NZp8xJzOwcNhQFybmv
My8OZtobjxqoFuNZqqEehAlcfhH8FnvHB+mDtnDygjPkKLFCopOibbu4LoYqDFXF
/GK//AB9vvXd4fUNTAMASviZfoFR4ZA4ATm4jb02+/PEIdUOS40YGaVbyMCP5s/e
/fs9DfSobTRq4uvl/4Et5BPuNAj3vhP1ry4VHH7jcDK4fAPDcAlLV4uM/VM1hGo6
3U6eAgY9y4s/SMQ96ITcve2RP+B/ZiZ3TXmWvzf6H69CRRL/i7YhIhQuXxRRgC0q
kvEoCd6O9LUpzS55eiCmgiHmMwKuI8Cqxl7mqOEa3XiKubhF15JZCR1WMifKtAb1
pzgCwPBzMP8b4oKruXXVszdCEAK5iOV9+2uJkeDKZD0TTX+yPZEAFQ6uw+6T2Qru
wKQT8ONDkveD9dvOnri9p0dyXsj+KgC50xcSFuaTYG9ElsP2NBHyw+l2tlzot1JP
18OzlmGmV+n5vLIsPO5ULwOOPv9z3mE6A7vhBlmL9nGKhv7ct2sm3CBk2gkbEqIz
W564OGp3xreK0UZIbFOybzBIxufxPt/K8fIfcJqtRMzZwdZ5D2NeHUHVpWVsZXrD
pUe0m3yyZcyCH3tMhBUgNwiW1uCwQfJ7bJcjQfwprVG9WTLgGqYQe+wYR+kuPC5I
wVpqoFo9vipHEqNSotCoRlX6Zgdkzskp8xJYNVG2xwXVj5uGLMKjtj3KxvPhZzXu
Ip3O965y7rlQqpKZBwgnKlwmj58pPArSMabSEI+ZlImnWTWfr2AyJMPcA0YLvReg
bL+jWVUva6HryCKlBh4Yy9R1TArpNQJevAyfywHz4wL85fy61A/WzmyiQKjuiMwc
JTKtmd9sDAygS/Q3HRN6r0/GFNVD/uEVGYlpXabUOYCaM2bvI3VtK93aYRkS7d28
bhp3GooTefTRg/ee49ApwBbWTdVpLaRmrf93ALxaeV1nbKo+Zs84OP6PcEvIIElJ
s1Zx3zaKT0VYbKOB31gKCBmwsNELBLqrq3XWzlPpDfVeDBkGUXu3EH1xPNaGXnho
6TLFx8Xcl2KfmWDW/SPZ/Z4jDBLJzDZBZYkFm1mepV+JgY40zBdkJf/POyUphlMa
uqOQaSc2nyrpUY13Qjv9Tqcy4yNymYPpC+k5KoEMl+P+usdvPpRaBFKAJovrt5kX
TftoVJNRYTdJdz/dZib78/y3lsD2hvzwK2JXDgeW7auijwn4uebSxAwY+eKXF2aI
VdzPHbTna6TXnjxvcN+nCtlLW1GpErTI/O+uyuTZCOX9oWcYXgBK7DH0M6BqK7Fh
qcjB9MYfHBUqpCqY9nvpIOy0bPeE62N3Zq1XTMYOL1hgAVAvKgUF0hEpF1Sz0VO4
/fwyqNSKEiOU1HlBD++2F5sg8Xn11bvkrcQ7oh4g761wUqkqOxyBYfMVn0Ou5Sjd
SPkzjfa1dTycuyLRa31nX1j6knfeffiD/NXaHM5gn7hPvLCrIadXEY4KQHhDJF7k
tDzwUZyhLe3RADqRNhkAzCopOA2nHNaO9Jye+09ExkoV/MlN7VeKXgYdW25L4DfO
s0G2fHvYKxX/jso9G73GuwjJUzJGZPRAn06bdw2D8NRrNqVgOy+j3W7jm0Z6tfpV
UHf7xKsrGXPIbmbqKuae2N4aXo9lX8/JD9FnDCfI4yhdI200s2zSEKrW3CMYQHnm
pQ/dzhaFagctE122v+GMBiTMCn6++CLyUqKNFfDHMyJx4/QPxsFFDRywVBWq+l1X
y2To8MB5FcTSu73V9BztPmrVrw9/rMfn+d/JXYtqBrfPvfjssWQZqgxyKo9dNmgc
OInoogp+jfWsFfyxoZOCAsVoWfsuLnC70c4qdKDSctmXLXX4TZ71hxJpv3Mh1hXh
DeMw+YreupVNGbRarMOAEnxc0ELaCTJevGt3hMspSm9LygD7TFxj5DSHjcXl+kUM
rq5BVn1SgSjEGMjVeXY0r4KExPOlaRvnCAMFWLIsTj3JCcyw8MYzggovIW6cZrDz
8Ybb4nzRHnuHUwn24b086J4Gt+P2w7Rc8yDdOJsV7SnaWvzlZoObnh78XzvWTLHK
v1k2PUImmNndGXCA8jTx8D779I+7Que2YHTHm45A6kiSyKLvma9bWV7fPT/mlZHq
52SDfJ5vs8FYVDiUVplripnGFw/dn06LhZ1ig98xzPQEk/pXjCnA0p8MgmFhMrg6
5CO5fDr/Kmk6w+vfs/Ht7f1srL0NklaVVoWe0J2RVIf+N/En2cA2XH+k96u8QRO1
SRqWRoP11JXvPMem3xRDUGs2OsWsMZomWZ6/cEy3i9jjpATnqW6zj3iuiN7IUkxx
KiUEOslcqynDU972ThtVLVIppyII1CZpzMuU+haNgDTNkpeevLAatdkECOAlRvbu
3klsY+LJvvU+nQihSuFIBxi7UirfeVvzbOn+nYyM8I6lGqfDuDlwqyNxzdAkFIgf
adVvqZRHzIo6lLTDfspJsi4K2eyX/VBERIiiIO6+5hmLlfKhN5R8lAmj1AptQU2G
4XGIb5xBPd4oYPrI++AZQP9pnPs63r//h/F/OsUEc7X7GUv+w9Jflrox8KeYcY+r
kz2CHtWHAGssivSonr6RvxUDGCA89WMxu8BdzzsmxyYRj9bjZ+NoYBesbUqasGvQ
wWSmZT82yWDzDPArtdq5G8juo1hZZBorkjAdI6mf+mGvnD08uBuWZO7V5u4vbDLY
55KOnQ0k1Hrb213m9onmRDQZAa/M1Bk9hHUKPtT1H1G/cQ7rkyOJNJcFPsCkklYS
FdctreRCHOZdh10FGQh5AQgLKBYsuWcIdQgkoxYb8FWG8kpoHbOo0vPZ/PYTLp6a
JmO4eSl5LWKRly/GvtsQi/ovnkUkBoj2NVaAs96ZKr3cB94sHFdJAfQfix0x30pt
Udi0OEt0uufsZ9kNbIRbEQqF5Vr+B+hTeNK1TjAWAWwzvKQkiLbXIkwnHjD//zcu
p2HENO8nWf1F+zO4tXVZnAOgBUQWEJ13Us97PkbPtewgcB99XEniNsDIBPmsBgBF
u9jRr32cwDlSHjMl4wE0HekrTgc+SLHsESAWrp3Q59EwiAfvgd1/7KJ4rY1545nR
OBE/efh9NxTuBhYsfmHl0PcHgnHjZQncKL8XSSEbgeFooEkxMgJtjDhupP6pHW9O
W77m2USdEAb3h90Y5WcA1bRv1TfXcK/vTxAfAbVFfXb/9/uaRrujJT90r8XutOeC
TIxSCkaV2RorkAldSVANkFsw7WZzNIpFp2Av5jJUM9E0EcTASORK209J5UvBXAgk
njc8Pvv0NsA7QmeSXzCrc6W+wDeN0MYDoWf9tgoR6xzkrc37N5bE6jMDkAAFROl+
m2Xt92q5bh5IIaFR3Rwv/iBMBGYCsin+oUrtYAnfqIJ16HT20H0KfrNRrkAPOuDw
/dIfHehTReYKLh+YWkuEomcrr+HS/3etuIWRrovaleSDGtches220yM+UsNRe304
kkTDHyEXPNMfsbfWXHudrPUx61eJDHU1ADTjs2sV/24hUsvaPHhFxdeVYhq25rM6
T04g/28HcqRl5CPXwp4gu38SdyKjhCP00ULzePtsAf5hJsPqWGBEXzx/UME7efyw
L6BqTKIrLL2dQ0Ipqumw5NoYNR4luN5TdD8ecD74PXRtIEW/e4XmcimMJ3e0d85C
7dT+GX8CR6Q4S4VBT/YbSLdbjWlrXaWz3NxSUWqUVz9iHlQAMrioqHHpztbFXtRa
+ksWMMGwgjDFFPLGOuACkYSkkPl4n/ppoGf/LJNpUtBd1EP6RXVKLTJlJHualIB7
sFn4d9KuIhCkmOqppAGxlsVDFtHfBe/u7q/x5fVMR5YLGY+k9HU1fGc0LRQ1pvx6
jRK5Xem6kd3iusxCweVnyI3sWrKRTuOBoimz25OoYYrJxnBeWaJgf02Cv/wQklsu
48a3x4FD7YlxVACbFQtpU1Q8MbZtQEx46R9MLb4Sr5hqv0VRXFVjzB9EDxU+Mm7T
e2sdaUI1JfC27okC9Qp651KvDxsqxm0V6d6g3flT6GWZUpjAf1ZoxBBTxAHuBOxE
IXs5ofE0XV02GwaYfRNP+fGrKxQiTP9jmlipd3uJHvpfOEjvhQgBQSls/DANysMg
ZgBATtR+t925KK/Fv5VC4SdUZuFhXznTkJB3FgztlDhlIoao8duzOjSh5IF8sxJ+
QzPvTg9MfZDBqMQNm1faIia7oyA/b2Z/kDQ4y3zVoTPGRMamezdptT70XP1FAqF3
4Ud/z7aGvWF/KK+IObWR0S+YHjmJaVW68CrCRFWso7c+ipU5ZLA0kisJ9QDBCJij
KgSOiINNMaHXOu9cARCiLW+buwkANr3K3+b/IQxJlOFcbFL60BABeFoL/g3nh3zP
f8wnx8ZOi8sn1BKOdNVzjaTPJxEWLoI/1LUBG4Ue/NvH1Io1AI5L53j8uPOAq4zY
Dmv+BczPh6DcEGU34CLu/4og8PxZM+ZLsqzvgeX8whmdvlSclYmfADAfOa0M67eo
1NNOl9JwveOvx6v3GdZnQLUrC9/4mCGcxmZ4TwX7872pUDmmE4+O3CYfSSr9QqGV
EHBKkTT+iaOXEoxucozNVfOj7YGF22J3yfIh6iFyHOqKw8sBsjGaxrzWK6SKYhvp
u/CL5qLXNIcK4JIgfH91S0lGAJ1Yys+L/a49LsBTX1KPYjrtKyMZoV4KklJ6ELhI
8d349R4hO4b0mSXWlnvA3JFcjjya3ExDuyQUO6m5ZWEKEklfTH3Zi9Fa3sHkEUp3
E2MUYvm1bTps4oIdpvZgcMnBUa12ncqICvW7yA3euvrcenJDKpJ0xfLKq155nxRv
eLONgxVqc6yvOBUvs4JkqOADL7GESUhZgX8uZ7FFAhLwGUcy3ohhoTd7cBbO/Lhp
X6QIv1TjQZ47C6JhUJistecffJ2v7F7pqqSFEnMgXqeUt+YWDyLz2oVEAd25NaW9
hcW+7e598I4t992kImWcYPj74GMTIRXjP5Dr9gHdsIhrfR9VPzFAoUGvGLDNwCMF
1YmqSUuy5TZT/NQT8EyHvkpbS+hb7H//kY12b7rghYkIMAtmvQehs3WEqgq9rGqG
e9Op6LBraJbiRFcfm6LDXVlT8IutiNZQ23Ek8RGoZX96cLJHFdbyorSEZcgdoRPr
GKi+7wmnkEjIlNN2kiMOhpA27hhtBJ3jjHZ3/x/O1nEHNV1jBr3ghOdGQkvgK4AI
o4BQ884zAeScYn9ryUG3f4aDipXbOxsBHcMF1ybIzmQdHyCDTkf3m9H8lzleJ5mO
lBxVFKs4NbCM64yjI/8V/S5/8vJq2I9oLrkovTu5E22f/YMYLEFjbV2Cx3xJHy6K
d4hcRpOfwaQeB8Sx/De2yGdvD0j+cxvZG3aBzhuk7a7iicKPkIWEn6RYfE/4C1q9
Mqxs0ESmJd34dWumbaKwxuAWQF4BBL1JSCFLI2aU0Aev1yRqk5cRAkaO/Qxbm5o1
0ayCXYyJykxt8U5uf3buh91fjf7sCzJXV4oIqqWfevKDnggwqlppF4wDOuQcBoFk
ih7RNgkSuXt+/cwwW5uird0tqUwrVJHCUNTCnPE28VVoDGJP4H3lH2uqpNNVujq9
byU79RRZQAoH0tu2Egw8Iok3s+jcQwdjYsGk5pydaBV/Tg2v85fDqvlhEarxHToN
rN+kWPMoQchW8TswcD6nF+EBW2yQUIJzymRznmlJMEVt8ugCWp/K5ObMjfUtM5gm
x6OYg3ACQ1tsZjZt/DrIbHlQu+L5+miWvVOaHWUfixm8EdLx92kqgTZYJAyNVJio
NHSzD4rmihgSVB9nAHdeQ+GxAKFm3E4++DeAIkjW/3ilcMGFlpf1HANRYNep42NJ
kjQLa5EEpgkpgIooUs/VS7IMsIeopCmUjGy0lBi4IbwmVDE9I9cQXlKsvVQ+ctl/
Wflvt++qXzXv0IrlKquTBWge3O6clO+1tZwquqE6dKB8ENy8uJI5x+Pw0f3h1Hez
w9Gm4DPGNCbsjgqIzHYUNLBxTceDAlcU27UwtQTPkmQNc0cXhto/y0NLgwsfTXTl
zZpfQ3+1Rn1P2mI0EjXnj5rZCUPQ/Mpz2xto554iiON4uSSutT9AG1Rxy+IRbAMb
vZ7pPs5jIMPG1dtn08ZRXX8DPuYfwaySIjY0BadsDblxDYhi0sZ28CrdQRIeK1UR
jGucZnRfQCxKneLMzHs8Jf+5yNqxDV8hUoP5sVBJx6KblDRAzTutG4thcgdRclFq
/grbDR6rvDApWheP4/FlRzRmyNkXmkn8fPLd0Gd8ac4=
`protect end_protected