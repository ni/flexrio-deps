`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
DwCP0UbyAlcaqD7JxsL/xFYNxZuxjmzs4Ad8jZVJmgloJn3v42k+yR8WDSI8xkrE
nqr/iCSauezNuwEVexI73Q0T6FjLIIACgDiQjtbitnssc3ZWxBdPke7IygNKvyub
tJPEkDIHapIvCrVIF90ZZT3DJLCAW0lVEfEkZ8GjALA+8YY+UuMrW+ghUPnkJwp4
lVVIXRmo3She0ZGP7vH5s6taGrgkEfWtY19PP9ZN1mMu+FqzCOG9oFIyXw023wWI
5Z/twK2+O33xtncdhAo142j8NkALT6RDPatxxYJoz+JyZCSGbPABDMbohDt3jl5x
N7036+/hqDz+++oGkRjcVw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="4tld7AsBO7siZRtkpH7X/PH2ZiuQAluwt+ORZOWptIQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
AXClCdlTdFT4fg7ewrah0SzYOkZfmyzu09XZywJ+l5TxOrY7yG5GEsayUg19hpJl
XSWiXOFVmnKxmdbAYGf/tbG/2tvkDVjpDlS8PlgCeidCSuf7mEHnLThG34t0eSQB
assRMXplllBmmt/++9q0WxvtZ19Pk+hCyPk7aaSLzVE=
`protect rights_digest_method = "sha256"
`protect end_toolblock="yKYLzsEawC2uc+z9qIazqPmu1Nqc4XWNYKwXpt11A6Q="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21376 )
`protect data_block
06CNjJQzCVBmLQrlc/SzqGOJ2zICWswDkSpXIBZsW+js4y7G2CbjXF1cNESZrl+N
KQ0+AZ4BV9l56OPeSIp70ZVihp3RH41x/L1uSgbyj3b6eMZvf+eQ8z14wALfTJHs
q3E8aWgVMNpEXpVH8GIRP3jtFrB5CksgCDQVQxA/SadnxGN+avU0kBPppC7DK0mv
nxFN88E6huNslKHc5HNFsIzrlUopg6SCx8FmIGqWqScZigvtnKo4lXzL2Z6GlJHh
k6UVN8O6L0NQ4yc42IzP9lUt5pwXpbKTuCasKa61XE+oJmWtUFUqfB4akAsvjPh9
epp0kyQg5+mZ68qxTSK7SaAy/v0ffGz4/tr9KmkuzSAOVK9UngkpeE83dWYsBib5
ibxikKoEJrNGmqcxCdSp3fyRubYyITlg3/WPPdvjpoPb6C3hJ8FIaTxzoF4jPaX1
im6d7L5PX8RHGxvoTT4KQqJuurMawnaPHTcT3gFyFD2rYPSYbzjz56qk5uBqFqQ/
7z4oy6dlPhwyVPdHX9mgvh9/43xqpIFWhy/LhaO+xubk6Kl8JLPoukzOYSfyTvqx
BWlgmB8vVFyt/EVH/lfABuv98H2hJ5/W7fhSI6wKibavlvIr5zLycwuDFCzjCocR
lAPg7fRcGaR9WV41TTi7Pp9ZVK+sWIUfbGEmu17Y31NGXr/WpTIl+NpGZuFf2mOv
/MDGSCEDSGtaAj+h6uEMHPu+j04WmuVYLDQLxe2+AGvgPB/1fSHUpxWjn5j3wVja
000OPMujY/1IoWIUBU5pVZ1JbasoJA8uJeW+0EyJr/Fa6I6D/DJVgQVfQjuzYoub
3lrUGApMQEllXFBYXKlvyHmIZOSLAAIHkZrHqmW6381Fl5Eesa0Y1A5YVCx/MLB1
TCnIr4BjgyrR2YI8pCYMaw0uD09lrykMQaTSlnDAFLUD20/Zc9q8dBHsv3c2awzf
dq+51CZGoHcDkkdqyJo9LaHUJqXjUFzXWphfdW+TYJTppKVz3gpjIGg5cydVfaxM
tykjRBlWqD5Xg+/s2KLFv6LqE0pAjFP2G7SrfSuDjMEzuH8eErbq3ZC9baGMCWd1
Zm+y15eIGmwXDUur//ZB0V/6VP9k9UFgUM24u3ZUTnjVxhnSIeX+7aPav8GG82MS
yikmMtkhjbIShm4syJrM+ddYCWYpCYf7F3bXKzmIQ+jgk+ES34qutQazpy730HDd
wrEM5AAPQ4Z92QaC6aDJKcF4xPIJJMnd2L9m4RxTC2Nub/yeAWW0gBOJh+1f4Udo
/tfyEBERd+E/LBl8MtL6Mg0g50a8mddkFmNnUEMqATFHxaIJjLjBqCK5TSNp0MeL
apy6dPMvlh4lI4ck/XpspVcx3dHppVtns7NHYZHCf6HzxaTSdDUzRfES8fU0hFCM
tJja5n+YgrdWe7k5tpi6hQI7PfLKgFL/CuwoE8BNwyTVw4ANSMymTTjE1QC5L6Y/
5tQHNKXXMad2QFIZ8iaTcWKuzIiAri/9LTatsITeMG2bibd132Lv7DwAaJ5lxpH1
aVh28QZNBIQU8F1swa/5kfUc5++DBI8riq6fLb0f8K1u6CL8GW0HHF/W0WSsGwvE
0+Dm4HCA3KVeHL3WVfk0slIc557g4Q5v467Od2XmicmgmHr0AqVxsr4Wr1R3RiFo
hrqOqLozPiEjvS0dqoyiT4GVEMdWquUx/WKF7wN11xL7DXI7/W5gFsgoi02p2rEE
s6Ix3FFHCLCOv8ZXNjyW2N+ZQ5WA2xOeOXbB1ScD82kydP56YOy7eEhf4GxM87sP
WL6T/O2oOxEMlxgONtVW10LAQ7vxDQRfpGZDDkKiGAti3T2pgYpHPyVv21EY1hgK
MWsNR3vVBKWiZ84pTKTSzCZ7PddfG0w3dLkGto2wj1s2GmLHGhAUlz19kW/+cO+Q
MzakuYL0xl2Fr97MO8LjGRPvvM4xpGkHdRlIxG6l0iIuQjWf4HyRin7NFGj1a/xC
l6UWWoX9qYwPY6DBLIorFnI4P29aDfS8QhtgCLFHgPVgLblVTmczci8/G0Nbra/F
p7eorwivcxhQSWPB5xsdlL70eAWtzRv5jvBffT/6XOCfkZCx1Mjbn3ndF7t7ZB9n
6ziiVHLO7IW7gp2X617U+czJhaxOzgQWNS6PH8F/Ze1QLzbTsPZrv1wMamWXeV8W
c/JaLgogUzCfHr7axKdSn6H2CZ3gE2LSTa4pguc/SV4VNcWd33Q+G6/l71QJC6er
nKT244n0ToF4lhRmG7/GAWTtubMf0JgPrcMul9McHDTH/A1lzJL3wLO9cwF7A4Co
6LPo5Yy+70lS2Hm1p/5yZ6UDtwhQ7sOULkcRqKFy/rTvXHKGl1UpzH5SNsoX/zYi
KXH6j5Oxe/sNRirAFMSnNNz8Zb4+aYnlhtKd3cbrIuNWUk2jQ4Ovun5F/DzhtDFv
NlTH/dtLuwH5u2+OJOjxHENnJ4eqGOBBUICK8mgCaGX5tyN9fIeR4LbJudmPoxhf
zQkKHnQdTSBTb3XOSQCrNWln1rlfUPEHNBZOrez+MtrU4xDVsWNqan52bK/S380w
3EaJJTCMe3nnMOn/ugFZhN4tRC/ycm6WlW+oqb0ttaP2mnr7f6AV5c0ahx14Zu6d
XpOdYPwrSq4AtJej5tAhW52FTO2d+Wjz1OrO/51kwHf53PwLGz5ODMveKofCPo8p
PmAUD7cySmsKXijr8NRbJRVwLSV2djttkLyTsM5/jGpzf2TbLGeWGFUPXJOIlRvn
xwYWloBT4WSWRZg9dufiywE6hjf4jZcje9hhC3ZmBg9BjL6pl9wuDuO5JRSoRpxS
qhLGb5wIifdkEgzuusrqeGdvfItH+8ZiKlsCFEV0S4+aMPCjLXKFm2mESGSehtw/
g4oBGMN9L+6ZPVrm+fm6ckikTZ1P2eBQ8E3i38EENuHMlC3TAOeSAsEsKpFLfvkH
ADS9yMENo0aMxHKRqVUvfvHHNcq9ptEnnun0euZUMBplqRpzCSFOoRqUIB+rpOJj
JOOq+MN1FXwebbyu65ewoa8w//aZaZCsjTqDZy9NnUu9GKEcMA/LScwa+gtKZC6z
iKtVQtmJMJWuaJTszTq84zV7+0mZt8S2HdtnHFqI/riuFScMKGdhre2AV2g79izb
iL//zToju8XP26zU0ToxTWjPiz5myioDprCwONfD59ZasacO9iHkGdiDHw43KVbu
QULHbz6SKGhrvd+K1WTrIULwB5wD15u4PHKdggB97qcwrlxGu8UsQ/0D4RPb0gnL
3I8BVcOn618tBKnD3J9NrpgvpungmElDjhHWa4TzRKRmo6OsrOedaONj7WRsi51N
l3iixSxngg3b+/RegWm6ENNzHjaICjaPKlk4y/ty9bpnGN54XujIfXkksUsYAJnP
gw8X+Shc1JrsMjBQ8SVdSvEr5un5jHoh2MqTQI5MBk7GXuLah+0W2eHHMlmGvrv2
sV7Ho5X6Nz81dj0uR9w9qNvuzOalt/FJiVv62ICKL14ab48UuVaNri+wEo1opV+R
+H//MitU5SvSQ3S9pv02rAct7YHMP3RW12sHigIQGr2T88qAF0Q9bjaxhrFkNiwP
F+CDIG72OsOTSV2w1hTLYLsjIPtDPsuRqNTDqqPG8iPu1oG5nWKBoEJqJri3DhNM
aSYqjhRQ47zlCFhSAoE4fB8vDhBSaqEAMXSaiLkwQ+R4Fb9cT31wURNibEI2zF/Y
R7Low6OqCJyl8T0WcQw4Mvft/NY5pLdhKt65kZt8gS1BqNxD0oBNnF3AXLoONUDm
oo1iponG+2NWJ3snpYF1jUxV+OFjLtoKK4al2sIL9sb89ljB0SrxXLTh3wIXQMrp
r9j1uJHkkbUQeibv6X4+cpdKkhSBmbxDaubmpOYb/0Sxt5sInwv5lR7BfHmoQbYX
/0Swt4gFuiubwBqWyje5if87uQqoXofkU5T8kiz/KWQG0Qpg+qhVLeI7NS+Ike60
PvYmyXBID81kxkeW47i+/3nc5wz7lM9aC/r5lGmrvA5FyfdmEj51ot8PMIMpgO/4
fdVLJLeNScTLp3hJwHIKxfqjf9V5e7sQbzdbPYOUlrtep5wsTXfqBDBOb24zm/2+
dKFiyvcWPF1FiZsJ8vnIe7djWbw2GDdHaBxgP4BzE2Qr6ev7A8MPo2XG2onkSLfj
s0vHVNcZcly5q2lhqa3YCp6rePPy+7elEq5fMacX68HIQWjm0+CKV7LcJMAsQ2hM
fwAw2sfmlG7uTmR4p+gks6XtqxLQpjuKj8O8gFmzlrk4AllQIM6YwxzhhhwxsrBw
2M206dT8dSW7d5twdkZhT1OWHJGuFuQIX506379p52AiuLa0EozI28PALqDxEFkC
gTi/dMA8sI7oskRKQ1W1mzX5UTbup2BIrnCWvC6qyBa/YyPSZJZiuVVbUaYzXLwO
OIsgQS/Tsh9QXNVPLnF6yDlkyWOID+Uul4lXG7WnYTglh0sMuzWmsUVnyy67Vuko
JWcEwh8avGYemCpzAFdzA3sRKTaqvIjs8hFFGlMGsbTuDdSv9UQFiBDX9lvvLUTt
jVAPfoX6aI/Yv+U9zMrIar/s7I1ZcG5IMWvav0KfkdCcUoVGhWHITwH+07PJFiiR
HR9DRyZPJLWl/4Txxvj5KhqyoKA4BoV3IhE6Cqv+eN8TpX3B9Ync0HXDb6yX7YUV
Pblrr4dlHUk/WvF2wsYIHftSoCe1BbPqPQxufANPOF2zAgz/QwS8HgbI+aE8hXGQ
dsx277Ttmo5uMWD6cHbLJlRFfo+tqnBfGKzNPtMj7oUhm1Lyy4UQx3F9Fnm3WDLf
dsaU0OLRReancyzE6M4oWksmO5m16Rcz3tRaGOL8FgyaTSxmtWucp+8LaAuZd3hM
vv28U5UjNR3Chfd5Ge5LdK4pcvnkyeYUHwaX3FsW0RarcCPx7zugB47kU6CQGVrv
XXjUMNWxfpvu9Imu8vVrLc4UbDh+k5s5Zeopr17bxvIKjwOMOwod/aT1+aUMyUMM
nV0O6qvO/l5tkCDiyX4YNblKqBwe5WR0OKc0g8UHdCmcCPHvlVqNRAotN7n6HwFJ
m7ljoCy2u+mmqFfIAVK2xKHriSZHyXUskQJYar5pRmnB8OQ8U7mc+yomdtJzBE7R
2HLtR3y15HBjMTQYFPbsppuNO4D+KzpCh1TZvVX+F0BFeSHc5YVek4RX61TF6kWU
hPxPnJLdLP9mf0OYbUvFVkiw/5VmK9MrzjqJ3bRpyzUXTXUjfk0ves+Wg2ccafuo
mVsVFmvWjdzb2PbNAfEPLHDpLyJ7lsVmBywq26+QechVNjT0BEmMP24JaXmJCqBK
3m6RjZNi6vIvaAFENRT4mR2xgq4W5DxIHTidcQRxn39WMolCgq8MTaFv6K/adKP3
MFqOaJS2plgP8HRa/WG2tBE/TbVG+VC2VnoB3/3bwyED29FSMvUahG++HfbRsrSW
AF++eEzWbKJ8iiIGx9JopMMMVmE3/VXRZZ7l0Z/wwsM/7mrWtdl6DWCqIaZKMSIc
4fzAZ+BajpXT3axZbkvnfFFHCygzXDB1eJfFJyZ8Ru9cos0GGVJbxC4ajxwAMYIF
BqR2WTvRe/HXGodvkozRCdR3onNpbePCfqm3DdAmMv0K6bHKcqTLYMmOnRhV/qEo
WHWQDP1y5xwTPeh4onosVX/cpiIWe7aPGXQZLbH3NH9p8Sa8Aq05UptWGd2Kk+v+
3OsIQtez9dTkIHRjo4ffDyX+et5nxjaRT9nS5eY6n0NPH8xQPduKg7kmI81q8jRr
jq+OVCdyBubZN4G0GeWrGIqQ2wejx3UlzO/df9pQ3mc20g08FuFpm6rponuYT3Xi
mKAA4UymUDuo/UjSnCJkOHypn/nYVlWGkzfS+jokRVbzgEX7vg+I1UftCOZV3q5A
xK+geVrzPsd0iwKCYJ/cv5fZw52UBCsRaiu+DyCgqNQueNZ1vIG1eM5VhZ8HowHK
4jT3hJ2zn7P65T/Tyj1DWPWLkqEy5s3/o4XmSGvk7W9XZM1dtabs81Hscl5p6KiJ
CvjFbwg9UnDHRHjjv1RVHy15MkJ0Z2msjDFhJI1RhdQWvqaRRTMITICwzgcKLvWK
DTWOsrAFeaPMxEYyJtJU2eswhZXGB59xi1NIzyRqi2VVbE1HQyoG2Xc1OJS0i7ie
0j9PVE7j2MWHAvLt2hlpUOLkk3kmqIzpbF1+pr8pRssNNN7hQ/gLSwu/vMYmuMQ5
TZCCpWcVxfb4UUoRjqGX7zOFPB3ZESO7JlrOk93bV8syGaBUwNI8a2W+v+aTR02m
4fP9WHmI9U4yC5mWoy8aspERCF7LQIdHw83gMBbl4xYfxtN+JlLffW7XGXdmbshE
WwNWDz+nKAwdU8QBuKReAJUIrgnD75roxnP0G5VXruLCXxv04lWGTt0nXv4l51XN
UYbYrucDiwunGJbjSEpuYutx7guy0w3G54vwPYC3VEl91/EdqkwIUYkU1VRRVAhY
IpQYz0BkkD+6i1DRp9Q/vIKruJeuOv9BGYC1d/mwgvXk/aQhuBfxdp0gbQ24J+tz
FDs5l0er38Ix/PaMcsb97N8Z2l4H00s5vm64yjY6qZSRv46iXvhBKkV8Tl5aTTEk
TeWoULiuHQoskz9qfzIsLyDGXAw+efd8nFe+pCUkssmlCPCSFgzYBuyJ0gLk8CZw
TNYVEV+UVyprK95T/xzKs/7PQ1jG7JPNctC9p9hk1O4V/pEbc+J9fTpaI04awhrt
7ZEzMroVHMrKkm1qXVOEJLqcHCg0xNtql2GgHQEwaQ85birFoMcJXS45PmfbA+7d
waedGcHEX2z9qTQFc9LCgddg9Zxu4WbkFZAkT3qNeVzKbCd/IIYZeipArQfHURUm
BQdjIpBPOk+g9L+GnqjLA4bUidfuI6IW4u0a6zBLe8xrpJtpc+oTZ573tEoxY+oL
sEgdmvPFIVFEdbEzp7NvU5ERjFabsw1BWk3ToIkK5E7swr6CMEB1EBrr+thFMZ9T
STSOk2RwtZirqf7itsXN/7bcJ3SWZViZ8Q72J3mTF23xou2XO+uS7rcNHPm/Ll+S
zAUC4+AE9tvAC1aO4RXEvG2JCtaTqNTgLMb0L9dxccVIupn8Nle6VD55OEVZG9j4
2RB9deumHTf2vZArXcLpog+DiDggD1AT2ZlB4cUXaXB5aPqBREwGl7dnivBCeH9X
+FGBb526V+oABicQEqeg0PuZlzZ+QoN6nYgMY0tbvSn+by+XngvkuIJwt/gow8eN
qd4+JuADpUbDm6FSzHljrJHWimIZ3GeGSXTkAVEQBwNukHS/GrcTVjjOXDs/ezFl
3I7N2ul7QchyNVcEsifsoyz8UpO8z3RyPWUvuHg5fbX2SXOC6+gxX2xlx18LCRXb
yeL46H4oxluF10N44b4i5QVOJc5CXamiR3NFwT6wjIb3fKzmaPERSJ0KPWo30Qkz
ucCJ0s1X3CFxfRrJlEz7JX2sc5ZtZFnWQQcfYcWt/5qnE84KOMlg2rmxbmrx2A03
ds8lkArDBQBk4lonwjyKdqj8tEuDanduF7ZZN1u92S1zwTshIUVjTAdhk70VRsCF
Tpn64xo/m5oCcnWwZ+nSRG9Xw3rsYUvfXM1k4N8/AlRPkr0uthsg4mL9/ucJKPtQ
mMB/CNbrc+lMLWPqRWAlfHgv91PaMt0ywQsm05l+0BTaYOP7PzAB7s8J+AqeS6i7
tG23yLA9jq3rvWqyc0krvlCFh1TbeMh/G+7pJo+Zpqx8tKHRsZ3z6BOOL/ZpsWX7
xh9v/FEpFbN3ZzPiofi/PPInaEd8aYLaizPnK/IXYxd4skcv0La6KCjwwtZXJc0p
8E23v1UnLYzA93+u/nUj4Txs9qZWm4e9XeBQ8LC5GdmsiGkEPe9BsaN6wWR9ARDP
K/hH4pYY981sCLJASIfHT59QBLXtcdS4aYgSc9Tqbpi0VUiVxDvu4lkjcIaYOZeW
IOi1l/rb7OAr9RVBPXKKwtRsQVuSCwoZ2BesW7ZnVNauIuL9Em71R1LD0kDBoSE6
XTYWP7o7NcBGaGDFmI9FVpiSXNB8opbIJGzNPQ5FYLipagiACaqhZRSQu7KQaZPG
dxVYuox4KKbCOlwFHZNJKrAz1NknjajOX+cfn5RXAZ479BIDO6EAQmUC7ROO0/vd
gCi7ahb8qYkdvYlLQCr5dkzk6w1dk3Vlj+PF1QGA8XQKuDH6c+x4dI3CwgphdEVL
AKNL2dwTkXtDIUH4Y6U+PrqErBWVCEnEYZFuqAKQWBkBQypAg73qeYtAecXTb+/8
UQ+FblQr7MeViv/VXHoy059ffHKCUKjyuLLIBNIIChjwh82GQtO4OuXT5QYifQmQ
MUrKW+VHvuR4wNzyq6Cr4vPYv53z9ohPgf0Vb7/oQl/6i8C74xVqajnylLkaDbaN
yHFpgOSfD39HqNvEGcoaUBS4Mv8k61QiChm1S4M+j4HgOfcE0dhyq/Jo+AN1YQDm
UP3a8yw++wlPmaAcaWCLADoRjQwTR3glZLPMpV5TXYR+bTPnYD+USLI5SJCJZofH
X18x1ns+ID6ONNXwmzVLGEt3RHzYOSmli6WpqE5zjtoPAjIHZC651ppdbwLfKq9V
WbF1oAAIPJcxIbsF+JFYxmPwUbGIv2nXdVB+ynTdYVemsi8VktyIuvuke/4W9E/E
a9FYmjbWEwtpVpyPiDo2j4MWQKUHPC0GiFVxulu9SNMyZ4UmghmK4TUry3wGQap2
IWjjf+p8aeOK9z6J/xZNyiiolMmoyjvOaI6bd2YEHJUB2lB3zGuZs4EYbUbo9fKi
pKU4RcxmQdCjI0LT4MjYaf4K7YAIs0oHepleWvRmevAOV73SY0z24a0dc168BEpq
t6LcF17xZd1IG/z80sHEGtEH/NoprN66LYu7TtMc6O8FmiXtUUK9SupYb1OR12Fz
WSuxXI3E89AKHxytQmM05xNEKh4VZOb+QsBJ6GPm0EgXisnQBOX176muKR44kekl
pWhYw3c5DyJzZgNUUAWJO8zFFPYk0Xl5Kp1t+Xnf5diyxWG1ey+XK4Wrqu8SIdHV
LzsIuxRCF2FQKzoX8d4Z80sP7/Q7/DFgFDv72mjl/x38WH9F7PnQUEaqFM4sh2us
o2nlT8XptOsxDYmR9VJkA558uVY0LrN6645Bub8cr7AikIoaTKB5Ytsc07aYORHr
sG8W4hH/HE9ZjaLvacqcTYgVvrdCpMoMFpk1IU5PcTcMLBMazSwTFbDsFWpMsXCN
G72Nb0LdCSsgQLBS49ROoW96qabvygSiBkYmPqG9n7F60/LiohgLUINzzdVbGzha
G/sNgaW+vGou2cdoAHMMTGUPgvyb2cdm3pckOa7TxLemwx426Rdnb4dxBUDATQzK
mMvZaZx2IoCl9kTqroRyp5fLAY6cE997O2SoVijsLPt99lh6RZYQy2CWWkR4LJgU
IcesDHMHC297Dj3jn/QXr3MGEzEuOBJphQgN7g7nlxWz/XrNhjPGSl8neubywH61
av3Vx/QgVo2LEJ2o1e1XYhArmlGVwIyw4cYzXhb3jh83hilbfto7wz/Dq4IC8oy8
nZ2NaNjiaGm2JWiOx6KfmyR3CDxNfXVCb8QmuMXqzsvpUhXNp2JMZoeuPl5reYnr
JGOB5+OD8SfvbUixcNpJPJIvGPEWBlQHYFmlLU2d7eIFNKs/OLEHPOe5LVu0J3ov
FFNP+sOEIJ6qGiZoVvgl93IrcvQUGuainPto9+HZK7KUtxbJA43UlYAsNTh3WlA7
77xDqOnHRaKbGdhbl5YoRcz1QEWD6bxxUp/J7zVImn10hhWDvlHBxf7aUEN3cYRr
eTQmePEXs4aPxUXEgk0XTbCCpgAnXlGYEnHFK1rt+psFEdIYwqkw1F7dpdGXWW1D
dfEQv0u5d6oXFJ+CbYEgOIsGmJphImYONhxua0dPPyAhyfWYP/4DIzG2TyZYyGKA
vejMGjlGtsswAPrBWpScaM2k5wTfov7kJ0FVIXqbEJq/wXGK9pks0T1AfmbzTdy9
inEIOuKlW3rW8S7lKiBR2lEskndIJazu7yd5oJQBlh60IpJNwfcZi9t/STWt7yaN
Wze91mL/eofkUReOgaUEj0fOXpKHmYIufE6HbjFmDH8se32S/3J/terSFU8L0h3n
6X70cWasaRMH3AZHH4nBLKLTrs8gr3nIogV8bQAG5YS58IBIGEQOWAsqAU3MOCWt
R42OZsFbUOB0tPkDXPGRNRVPqVpAzT7YBSH//4MEBT520jxVrZ/UkWOzi3D9UnVK
YLtMyuvMAvXu/GIBp2f4v/lEnEUh7+nj+DaCL5L/W9rtw+G/+jnnfBC3sZCMGB3j
zh+Dx/bIt8yU6epqZaf3P5RvIDSFm691ql6MiFFI1rsf1tvm6JE9+rCbYZ00GgLK
S+vDKx9YZBjQoOb8NXSittrvdeVbC6LVAOChVUivvgg2Iouu91UEZq/hROhNCooo
O2irUDaBRNy0jzqM6msgGVtKhJbntjx1VvxC+VqF7Ivg/kMGiD11m41p4C5+ZjFk
XOCDJZys1CZdQ7jUBTwSOkaVapBH2u+qUG4/qiUZnNSQRSHFLiObn+4KebFCt+1o
EphSmjySF7S2PR+Yygm5AOV0i4iou36YSMH5qbtGSlIvzP8BgxeWZfWAQgLUVNsy
x1J12Lkssb+gJGiDvNBPfPLuhJ3a5xeZAqXgDE2+TzG5F34+mkvo/KJK7BovIwNr
Jsn/EJSa4x0jSaJKvsclGXVUnkj9y2A+x00eT/AgtUSum8FYaQretPa9+/Wmjmh/
EUReKgiHciVj4nPfsqx2/GCIIxYrFfRv+Cp6AKdhKX79lBBM5YX4ZPySPSeXZ4oU
F0IJ9IkaN3L77Wmer2WXYOgQV0x1aKFYkiBdlWW5hKRm/A+EfEVAgRwYfwRIDm7g
8qmLGKFVx42GVd4hO/fBbLWplZqAcQSKasjxseuoplPOh3fMs6FPOfYYNBjbZATt
XBTYHGlMnb0JBSkxaL2I862blJr++z4wwwUzN1bP6qSdkf0Gec0TpK5BoF6kIx3g
/UI44k4Sg0XPFmyJvzM5/eT0FeCNLHwOJ7sQA9yQLZ5z5xxXvjhQoppBjel3bLml
WiVLpACHY38ITuR1GCGktKnCXaLsdReKCt7OYG5UqwLDFAf0asZWUf56e1SPUcyP
msLm32vqtHJJizFXLaIpr9eAODoPKRn6AcS50nsLDbMhdIPa7RXZ9TBokd2F/MUS
JMR2IQUqosPmmSFtDALL5IqIBzj+ruW0OUQ0XZEO0YTt5Z/4VGnxPD2I5WWuBD+L
wdbTndTReljiUR2S4ilZGu/7LCfGo/Rdp9IppI7inq6BN3D/GVDKgasww1r1v4fH
9azp7Yk4m1E1h82NRqRZZem9/D4r2k2JoPujXSeWJVeH8SJVRdJ4AWTGRQpH6V6P
dhAdL863462ISVak3ShAbARxVe558kjCypVsQhe+sQIOYPzc4mQa1mHu67fUrISg
WGcVcpdvxYQOfp63rHEFSIeQLlL3F0yMqOYRsuykv6kNa8LX7jp9umugHcp3yVxi
pQ/4oSpWn3mf2MPwYBqY3Cfd/Vxdkkh2I8CEXxd3nyNiAA5gGFRc739N1oJoZ6Aw
bR5N8RjI7J8gLgdAAKo6tTAogBb/3GcX69W/agQW/MitVIexPMjDeJ+DZGURYxAd
kXbcnXE6HZeSGFv9UB21usEMA8x10yI2NOL4euFp27TMBbKLf1Q4sbY+b+rZTxrP
xhMy1DR6bypGTSiQ0EY1JMEJQ7w0dNdZE8L6aDdZ0eikIHRN5qGXD3eWoiymmqZM
+gOlTcde2lEJw2R9fqBoPc18/ZKnQhtleqBGWfZzfEtH1ayIgdH/CvnhXcOA8CTV
Eck1fjE2Ioveis9KfmOXT4c+eJ2GXd8TKkr8Tc1/92sB5FGLLk7BfMfDomqrjnL6
rH9l3LKlGJetK1OflIe/Tb/XrCR4qRp0JK45TI/rc1dRzrF2LVMbBUIIePfElNkV
L1TkIb+1x40j0QnPo+MKqBUWqxvOPNXcIqVqZQOSrCqQFp/JKkW+a+a8AUV00V8k
czNxS2zK5dg24goTHCNDbW2Hq+N6yIORF3hidKhQVxJ9JWh60EKx48ggLL6O/llo
YqJJ7FlyvPDDcDNbwmTTGy5EuWgLUare7TsXNQh6ry6Zkxr2jMFIHgBHTB7lZsyg
c5J2zYp6GtJyEjKBRDKe4UWq8/RZPqwAFKlXA0EILSMg3MzkQPte+HKVMDW+R2Fh
IttITdfA5Vc8WEZF27YAMjE5kbEUW8BS0Ui8b1aVto9XGWVHh2/UCybAGzSoun5G
VVLYQ9qzo9q0UIrVcOoNU5YjKf7Z35r27xxLV5fmvkNC3DlM2Ctwk64aZH6TDEy0
a/IDNpuycD9FRiPx/L5uSPCe3dExpl23U+BYLx3Q3d5PxJXf6x84Q5L5xyCZ04zr
scgewaXmprc2DamPjn3U5YgPSI9MHBg2rEVPKxuOE8AF2VDKbBrXU5hM4Kyxotl2
A4SsuMnxG/Md0QEd1zIWN4baf4DM4tnk63VHsOHJeCrcQF9lMgmQHVhPUioLozgU
914CPIg/IPSa5uOGM/S3A0aY7akfNimNn0B8RDp0rY8ojouTCHABHA4fnO6jBHQ6
epftA+cuk6B7OV2xgwDHR6itx8B8XqV8Fe4fTrB3O+4ZdPFKDbVAlOcQ9B1IbVZP
On8JIAnkv5GDa0ypHKVkSFN3YYJULBsPgEuvpCKc55zitPwuQSDTnSMj6EcuCNz2
w7NfVMFZUV9Qaa+fRRKW0kaH/OogVyZuXrTdygrbt4NPsWRN1FqOMt8R3ef4dZLd
rW6njJ30f4QQ1DZaXO2NC5ky49m+O/39by9Fe+Eqe0CfcdBK5IBrYIvGM3lkqwqo
VHVgV4a5gn9gG6JydzaRhMWF2gF82kiJt/lKgk5kiAPTZHH6+VDyd0awJiRpuhUC
Ts7xXSqbX1jLpX/p79Nie2mfzQK0Asr5yF6ixqlN+roRRDKbld1+gRTx/vPdilkh
Ri7pSykR2IIRChkfAwmGA08uMPNU9Rhk77NB0N5pB+yZyhY8oDIP8stoAr85+gQC
ucXVQQIk6oT0B8SVqlYVSc+kffJxa6O63+Lnpc3Gep19kK4b5Kbijg7pIOjVeW0s
6EZwkz1Vw9QSRrmJ4I1Qf2sl4inVpXPtr1PvmDrxEITiORp+CkhGh0HSyfWix3e5
fxopBDA5CtuOOzhfhcNOSoU76BujQesz8wjEMjFWdIbxscxH71NUkIvYzruCKYud
fecRcelaDZpiakBd2pPRcANMM0Dc+wpJfz7dsg0fcKmiAfk8Ev0N6s9auuD26qQN
SpdPAp/g+F9J0A0g2Cc6i3QKnsYdD9zRV7+2xPiWp6qdSdGehysJ4nEDfobJWEJH
+ozKZPFzl1P5hFTqespmxMNoQAjtAXJKjAS6mSKi0MD7SZdJoqwex1UpF+yAmGyY
dCmWRCt4V/VIkF3LC6ikYpKOk4kBGiuk3b8fl6tyQMue9ERlWxnKMQgmtp6UZa3j
MTl3gjYHoO/fbM7plELldu//L3jU8zx0OWmSGq0rB3/r0AqKyBkGLVTDaq/fBZqz
Qt3Ai+vfgvNPSvTfTcseiwKD3YUT+dG2lANOVZWgEIv88qR+cK4mcTZ3L5Jdu8Fb
Bghu0YeIbqW411pHv6jZ7QAJLiA3zwbWF4D0ZBAsebKITikYt+c+ea4uLtJFRTXm
Zb0GuzINIRhDoW/eHejENa9K9/vJvkFNE/CVEGOkV6GbgpX3TLdTe9xhh0QXxaKd
N/W0ZPbGOT26ZLARhbqO+lX7amxV5SX+TdOV9po0ONeWmkSrYYrBP3ek5Mjpkb2m
OUtZwaKsl5YpQ/0R+NL4nQ/RSTel65cu4a6DrelErB7yxAOjyBLq0gl/7LfzNSk5
yjgdICxgeIPNFTbLhvM3xUqp2bgdcEG3C8RBvFNeYR9NU99ndQETZ/PjMfEbaARv
LEjcfjxu6n5eGSTQ8X805QcbdJ8gnEh0LOHjIfUzKlMBdb97X/HBZDxwDzkHNiAS
RxKcr54qwAHV2N0dtipix7PRGBSCC3J/RX4N93yFeDxlrC5NAzxBDH1K1BvZ6N/B
gr2qGgN4wsNqHMrdjBgj5ekApzGUf6YcO0DvBVuDWI4D7dk1+p/BxjTiBwsNO1g8
s16FLVL8AUdtU5hlMbYZ35vdeotCJ2I+edQtfijEtyvgoit+OEoiJ/2XsazO5m4e
vjM8iZ8cSRgfO9PCE5t/3zN8ANSu60ydojSseDyt48ovXhyL2s0ZPHrK1loe8h78
v/X69gv7Y/bZw89ppTDTIbSrxF31STtfoOuCUd8hT6eRg6D+rA/pE5O+NRpj5cC4
yxbcgZCoLjI3pEzAPCqEnLrE38JWAhl4wNJHdWP+I99fMu593a0jLUa8faVPaRZU
Lq159C+QGrx/hGuYDnOx2iShwEox0wtQsWBToulvm1H5wBz3UuVaL/QyelyaNi4R
75/D/gKT6uYdBqthTE+uqmr93LgmkRew/dZf7OTFOdxm1pToUEOx4l4RONeGM9qw
DZo/pdAkqA9+2m5peorrgCgLJO/8VihOkRyMs1vPxvWX55LiKiPimWOKnrzxwAf1
1EcGfZQ3szJ/9EJt0TB08Mttgyr1jjBOMycVoIhniXZllCMgtksaVKmEcn1ksFEE
CuXP85tYK9f+CJ6vgRCIsUJfPxMQLZMj8tMEHADCpu7alcLM9Y3W99XI+xFf4ZsP
FhRKER6VdcUaqSFA3dO8mlji614nmub7bBy9T10G0dNpmIUrCsUX1mM53HGs8iBs
soGuECKmS/i6RPFziA7lfY0+RdddTRVQvnms7PQFqNabSA7A6P+dc+d5yuhOTLYC
ZVAR292DPz5emkjO3r+ujSJEnyXl8IRA2nZNlkkbTfm86AyTBLj4nOmrz+PJrBnI
qlXonrHmVpb79UDdD1pGOz4BeUZkPAind60CsKcLKVfhj8rpqSsaoRJODxHzhSc1
dno9L4jLZGIlMjJZXBB6hbWLl5tUSl9n7CdzzKGJ9Tpg4CBOZs3xplJAH9z2cUX8
pXkecUwd2OmMHlNh0guXG+B3e43n7ahe4CvYUBa2Gi9ZN2aewGPn73Ro78ePFVLl
dDMVlFyFx0+o9N6p2s2sdqE2Zw6HjVl4kvfkJm85oIwnsZlxVRfFxxOkoNSFEPdG
zRiF/PkLKXHjbmSiCECmihqZL569dJP/Z3E5on7VXO3IqJ5o97sIIeTtigXCNE+N
9cEbG5b9EDEX9OiW4x4WXgx+hrsgbeiiEPph1CWdudgZq8F7aZVO3vAIfiPqWLmj
dckly+lky2iuBb93UnuCXWg6EOCe/TLth7twAPU9SbC9ppwsj7qwiruGTmaCMwxM
9gZi6k2CKlHGC/lX7tHqtpHf0LzLmKVsdY+vWGcbpqadjHDBjtbRumekitv0PGP8
ZC6dbZSNexIRYraucokEZIVwbtM8IFyqi6w9JHDOLO7oSmNsYteGw7RTX3UJLbqs
D8LPIg93boC6CPnqbiN9LkNTbJPUwd6uO5SffXIgEttk2JEo6nakkUdH7J7bCuA5
ORqRTegrS1B4vh13Dltz1b2adQ9uuo54Abo3GpinBbguK8tKILRqJQ6T8Qrw+II2
pMZHQnvX6IQgHZ5vFB+nSoMG8vrXqdPp/ZwLCuWhpdvq6+4nY7ceCTK2qqgWrDl/
WNGWNCv4KalmP6sV6eI4gcugemXvDRrxoPgxF0iN2ISvLjsFspKsfBYmbZNU/GNN
gXnm1rADZxne59nrRQFObw1tuHZdsNV3N/6mjd9qDhum4MCK/qrPnclmPDrLfHd3
tYMVRYtS8OBalKtQgnM19e15KreOOoMfQAcQZgUU1E/qF/ZQC3kCdNbm+P1gSFcK
JPfm3tODifW4/2uW7BCB6VKzVAEVHJlLm0zgiNqiDgGoVJ9hfomyay0F+6gh4GcT
mznH+3mk8smZ4/ZgkxZZBGiUWOrE9E3hLnJHVQ+yBh5sBmKlXd+dhtzpNqdtjJ4m
TToA1gmL3erLnDKrUj135gWDmhNiPIle211sfn6gAHI0wXezrtB4Xb7lZlLl7EL2
ngkan7rQK8wd7WZ+hNQBgHTc5Iooa3obrQ9mxbuNd9gn6dpYvwXP5IH2jDsKA0Kh
STwaWJewvpPqTnBQrEfrPalwS9yWmgNRUPp4+aVzN5nBntl+K3pLhqQcLaYKD9y/
iDLioXBv5KhrP2Op1hfhDFo8ott40pNjVPe7xcgmT/NIS3Khj19jq7QYy2XijM9q
DcE1Ds651/4fODYgxtJSv+c9f7EknLlUp+nao9tRbBSE3yanUxU0F2BWiGaqIsPj
ZucRszCO7hCqmcaJluGek4nW2ZyEN86/ZpFa3MkxdZOn8oXJTFAOpnMAhphEsKhq
g/87r2HToDe1z9T3GEG7v8fsTiN5kAnxPg/85snBwhcg9Tg1jPPCzUoOOoF+bgfK
qiAcD72GWyREg2Amm1PWPSMlVrI0DKAo1uRRTAe1Q9r2F990WcADvxFHwb5Ou3Iy
SpIqSSuIPQbgzAJ2Cc746bX5KKqD1/dw2mB1+SOyeCVSCUNbarL/MDv8VkCpg9Q1
o4lLpf1qixrPJAmeLN645rJu51XJxc95jbgrJ9JX1AKM9ZSbLvtCOG1QT0rYjQjg
5YtOfqgvn5xT2L63x4u/TvnDf/RVx0VD22zqA1ZE6GrdrGEoQ/ZXtk6YOSn91OET
C+Lds6yg2W0CSre1uztjqtkCibYwK1M6i/M8hexcBML//9YRREIt2iLS4SM1Nv2O
9h9j7VP6nHeMgT3dtGw55NB8qKa24ryV2yL3duLYajq0l2Ipv9EB2Zez0ORXEaVV
gD0KEwJfhqW+LAPFDrOo2x7E6H7fqX07sbXfRaqyFGqUZr9yxAYEaVs5xzBoGEe+
k7bE5/daD1kwE3zujjHDA6Yokh9u0+Dff3BJ5qE9wMmKz71hPtz8ejRf/cNiHPoN
zVL1Zr89SH7A0r4svRF7u/nxzXIK+VJyXVYnOMW/q58+CRJuTq702tCq4Ozsbb4e
iOeXjZxfE6W5cfBfNj5auBkcXbRZa/0Lcn/SBD2UN4zJh/08DkhPByOkd7YowFID
Znjmt7NfFqNQscmNZQCEJOmrA/pji+e9Pr/XR5kpPkFNo+ch55wdprYJ9UkaUMcb
CmnxTV8hJ72Pe/GGbjY7oNLziYXFUV611TCT5GWNVfkzp6/HunIJWbr3d7R9YTqc
yAkOZOFzJt56bZncOpaOoni0D4KQmVcJ1Jeg5qKbE5sRPnS8WPkx2mti9E3yHb4i
U/bWQ04qlysmMtrzWPp65AeOm4x7uue6ZFdQfWy5nOeHz6kWTXZj+D7dPqIsYqoy
FuUbBIHTDpQBkZizyimSJ0ngDexdCgdeVnq7likZ87hJ9LzD5d7yzwa8M+N9CyZf
WLajTJ4qX9GnH8b6e1C3lnV5jAfenvvhs6QpjonbKYxNiy+1jOnJEaNamj1hsGrS
A/KDRlvNtzExywxEhl92eW+6GbdPPg4PWEd2UaSqY7XBQMx97I7CCY6nJINtKPYR
Cn6vh5RBZdGt8ntS4wG1iXBf6FiZa3fhxg0R6LskWo4EOZispg+UHSvksPPkhFBU
xd7SmMFEsEd2tOx85oNtBEDZGrguuNZdMJO2UuIDdQ7Bp+nL7yOFeKVjJy178a9+
OhpnVnEHKM9W+g2HHlpWVCinOqKn7VVZyL+u6PaXklKZD8NYqe9UKEzISy6J+mXj
DJc/pyrW/pxt84XNJoeNWhfqoYyW26tNZ6cbUpID3x367TfbXv+XjOXOeW75CnDe
4Z4scB/HCZFmQcM6D/FFdLtKBmJHni7TD/i5MMuHf2/vJGcZTVm04qtVP35vCQRE
woAkTQP+s4kvXvwxo+4T7ytnlMVgmB70Cr+pIt7agO+2KGNhWS7oeskk5t9jCy+m
sQYcfz5KKbQQk8Yoru5ajg5mEk0e81wAkl+8CvruoyT3CNRJq+8DwYRRng6AqZ7I
C/rOSkMFRquuUMQTOsH5kW14OGd+jmafpBzuHYKhVc7+axC9tMu8dX/ilRpDpHhY
SSBoSSvG9iijPlkkk2mGe/eZt7dn9KTZVFZfUFRdgrhu4Ah9y1bnstcjcPUwtPv6
MZAjzsklxvH1E4V3+yEWaqN6yEG8rr5fq7SOWk/xqOJijg8fFhTUFOhUGju/4Gql
Pm53WzEOXxWOhN9X0BhS40OND+0BH2KRvmX5X4OiGLUoXnideqU+iPNXiKs8zGvk
lg7BaCQHectl0G+w8dttSeHT9lGcb1o4UocfKV+CnMODhc/PlgkiZONal8QY5CVc
kL/hmNECQ/9TFKkkj7dfl4ccFiErTncVd+OU4RNQHv7YS3AknxBNpg2n4hY6B/71
UMGJgaiD87++IFnXhBc0kDoy/FaHlsDrcfPC1yL1Wed3dJ5+2xBuhyJbumOM/szI
dYqR6eK17F5xEfeOoUqdbha8p/5577N79vre2c6+7RM7667L06QJZCrdI+EePyM8
AANT3ewLJCfK5RWzP++Nw3JeSXRpbkNSRTepgsS8dkk1e6dPDAn9KV8UUzVbM+Ng
dQKMyEon5EuCd3ur3WNGjwf/OOcVZIAdPcPjj1mzuytb82PrbtvWTD1ReczQUnuK
7WDIAUxMv5uQO6Ibcf+p7oH4HsN41oodVs3hXnHHStA3dxhrtayurBrStuGbdNIB
tjZ3IAfgCqOn8VXGEm0w+dP4lnGuValf/hzYOipifJxGQkJnju8+s051iACg5aWi
ETz2xKfC6MC68kUgsdQTulSLFVZfA0BnRGMg5gp7z9iN1wDMQm4TOaSFXrmCnTg9
R16NkuT+f66hAjAfKYMSv9gAYK8zz+py4lda8JZlQJbTcZyVAs1Pk2nDI92OporZ
nXOxIBtEp9JpHkJpOH/a6rnacQqPiEArZUHZGZefBWt6sikVhhi6HhwcbQG03ZLn
bHi5M169yT1Bzrsjd00p+6rroWWdBfc0CujPvR8b5An4XpFHeu9kTEm8/yzuE6l/
DRDzm0NjOgaAZcdrCMTkIBLTmh0SfGwQWiJ12ibGHsiCDiZx1ktVf3TaEMLALb41
/HIY9laaNM2+tuSRM4Nig7S5uuS1Z/WybAOCBCJVeY8V2kr6reg7BD1d4A8L1pbL
48R+86jeLR4tWcuUMW5Vl92OHM8mTjacNL5mJpKeBMXGpHeWEzvGXHBDw5povcV3
1xc+zEQpS7pbglvr/luZzqBu0OKv4TGf+GcQXD8CPKEcetBBUYbBEevepWpro/fK
6IMd6JZ9Q647mUn9pi9dWbzqth6QlsCq+WrsrhcXr+KPLBM8kdbSgkZEIqVVqJGu
eQh8XckxfmeJyosBHVGDZK7/a8l20HIBNCQoP8oyeSg65UnuKgIjnZfmqrZ98rUS
fXfHBPTDu0x9lqJajaBnpiPpqVe5VHXKRfwDlDcVASQoC9sP0+88bA3lKJMTl/PT
VWjaeHfOGlBonNsmv/i/Brs/KIbU8nwZbAPT45EwzLjj5PLLz0AjxUbRt8iumAag
mz4T9NmlgcE6E9QDeWyF/lrtPLNTV4+lwSuxXwgAPhNEk0ihgsfPRJiYDDxAEP0X
L87vUGGngTXWw3criIYwyQhx+eNo1b2Xr3v9RiK5DVv0BQNmmyzgDbECRHzDFmhP
ci2sY22FEnCXs0Bjqm3fQ8JOeZa8Wze74D/Ixw5huBSPwbm3tHtQPajMP79WxQ2A
WLo46r8x0C38mz0vAjcyAUKQK7PoGpqxzbJpXxrexSvJy5nLci4MxFtuQytixbr7
3Ln2xmI/J7IzZOLIXnbWnJgNT48iyAky8CW573J9GubteQruVP0B/eT12vOiYapG
Nvt0tNTV+KFs61anxUpP8w94DMInsFj36OCj4AyaYhAcQE3CX7o03GbSu9F2y1BO
He4zoEqheG+Mvq7XeHC5npmWib/InKNZEOx12wnF9QFGPUfni7zQ7DLuFD40Dal+
SSVhbOLg5THFIFP2pwbvVcEse2nQKb41hqobEPEKpTpC5kQIggElyiCIqKF8UdwX
XgILzcE/VLMl/jwBP3X7cLXoKweR1oX89ufVYrGcf0dPL69cawC7Eff1y0/Mv/f5
x3/SD833Ki8jSyc+XrzJNU+2Om0rN/+0yAc6Is2qGVgV2OepuCysHOoEg3GLXuol
JQH7Py5zfQikOaHf4ycPfBTu3zMMEyH0ewGEKvtxXmLVUVkXFH/Kn6wWSUhW8dLg
4lwWR4YOSgPNKQuJBGpHdQNKx8uCM94QNZQiSWMPR7uBixyZ1b3CVbbnwZ828z6R
Eeq68UYqCdvqLAkZ3sKNOC4RT8hvai5n4A+rmAF5xN5IZAv6TooCCD/qqnBZWTo8
ITyT0g749sHNsV8OuyjJkOLSz9gXusKHtB68MXLT7iSQJkosb0olvGBetruMUo5w
HpxwTlKRXpAqlHskN8Md7kmLpJ79oz61kPhmYpTIs/toVG+KR2Fa18bR324zTcCC
tPayYBbi2wrlK/Aw/cIatKIZgQTrtK6GDCH4Fs+EhP1Vc/+owz2R95vrLufAAp9H
pee7f++AytIZVHNxz/mmzPuYB0Ge7IX+31dyOlDVorlQ9fZlWG97Zp3/2BCbLN0e
gVXzi3g793L5Skh7QSv+sNBNUi4FbJR03LMc5u6Gc24RtlD65e3mDPlynWbRIFha
2dmVHd599G5Cxm1KJ4DAmsXqGdLUGvzqoTOl0rMp9owF2BlvAiQjb3DAExWeSNac
Y94JMu2VVHCrvfc1LXoCQ8AJnpEn4YNXhnySftrCbYjFmV5a7gHG/UJoZStB6uE0
l5TErlQi/QzLvxsy1TOzlbn5CHZ56RGS9B5SxWYK6YVcjMEJzVjEB9LVY0vlQJaI
Mf2hW2hXT5PXacfx80XCa6U7ekf3ka46ZvFwNixJlklWHOyO+v0gmC892kyw0iwY
AX7ahm7J5ZngYu3Gjy8fYZikPIAQu2cHCH5Xj9aSXWOKH95Lz1JXrlol5IoOAoAF
4UmRzA21FPRCntbhkIgNx0oDUvJUkEnevrhHT3bsZl/e17lTn57tkKJmZD2DLq1s
PNwnYOSeBagidBAi+9pY5sCKuHo+ce2bTgRxoLQwmN+n8xBmuMZYOQmjCij3qRRx
1oKgsOifrEQ1rWD0qBpYF2IKa0ZlLuD+Hrpfk7AB4X/UORim1/KZoUcCk2+p5LUy
v4nXdmPIvW+1t28Z8Mxf8QJfYIcNipxp377vK0+90SCveC+Rlwxet5djLsKBXLg2
iC/VLMT6kOpwMLL0RlSn/so6iH1f0bS4te/7VUAWnCXLMY3iTUiy6/+w0yQ3E0JC
karni1sgCPhd3E+++YRr7owgn86q4hA8wDMbvNMqfK/6pJudeaKjGzWxt8Fp1sBS
1TDdEZh6yW/MFua4rec5oGHpGwjsr0vzG6hiRcJd/+GhwvA+FT5uCPGK1AWM4hZa
of7SmKIzu0MA2wb+xcp9bYaoS/qEpG8k7n8EIxTB73F0SCshuBPf/2okZJqbFtWf
ndPv+u2UmAfPq6xcmktNY8C+8/nlRMKPYDppwmxeVZzfC+7Ng/Wyjnfd8ax9T3Mb
QEZHme4DfASoO39BjjUU+uLidmOEkNI26sK7lRQmZJnUI6qTkQoteAjOzkc/tGER
bEoUkJ3fTqfG/0pKz+VCa7ozDwvP4hg1BRfBkj1ekx9z4cMWuCbtgTZu4/JCzwLZ
Hh+N+dPMIFpsuQ+IdOpoT01KZz+hyb0FBDFV4tUMNNX4BT1Sk4ghakUu9881N/Mg
F0sE2FtYJrzzeP4RbisYB6owmUhcLj/u9rRyUtP7WkSnJTLqtgcgHuVLST1jNb1m
4XRhtblX7rWGvHCqhF20bufKhJxBAtcUs0SW25Nv5OS5nWKf5PNn/FDO0+B8F69C
ae0cBVFKU7evShPwdUKUqYmydxDaoeIb4AZ8cK5p1T9FTA+MJinT6+iS0TR+oF7O
7ydOYeIPCaaSHfycYACpe625/f8QcbPGh7DaIefAEwUN1f12hrElHfs1l3OnLP1R
+oRifxA4RNIsWDxBCgJWJOB0A0KWWY1QQRiMtMwtwWqvVxAdUZhNo24WLwKX7Ok4
xIJFikgQ4dlsSzNoK2ZzXGLuSPkyvmUdLGdt3CCnGdfw3Xn+ZBJIHxron0lEGoit
Xz/V8vvd/kYrNwsxLrPS/ybor7Pno+PvEb3wqQL/6FG2PRUWJMf+Rve6Tnht4+lW
hTA41rDDDxigEE1qEqqlDOfzFwO5CeTXAKFl7JwksD2CGNIh89N6W3jPZ/uvAQpa
ok/BLvtx7DJ/sTq5i2401cS5PaSS/DFnCQ7+29iHcOTzO+WAy9QzfaaCcv23fn3U
jyY7K8Ln8t3Hrfze54aZtw2d+VOPp/Th8JMWbDgEELOUbnl/Qtfv+XMiPUPYKuQs
JpqAXpIOExk50VnBjT9mg8rvIFmNLH9Y9vt3R711AuVH5gEGfCg0qqkaf9R3bzOa
N2nnS5itDid5RUM0dGZRkRCikTj9HI46cOnxPQFcXYiEyqXv5Jia04Yixz3U8Lp1
0GkzqVAhWLDbrL4Q+2Mu6qDot/pZTkTTJgHfdvuABlKG6Cb/iaEuZ5viI6GsBgHI
diE4eTNVqAaCJUW09WYIu0xenwBLVeL4FjbO5HrkBN02Lr1qNQz6iEjaV5UI1cYh
ML9zQ1pz8oIdRJurfq0EojGK/5u4tq/tVgiAT7Kvd6/pKD3DxhhTRZ3ZpaYDhIn/
tIs6/WNBQIxVDhHPfe5u7nmbV/exNY2Zmm2O9QhZcgAKQlDIey8J8i0Kj+Xs4VME
n5DWpdpqMPqdpHEYy0wP1K54l+ZaxWZ2C34PJr+RbOBUCJZIeoN/obJMo/Nq7+/O
hGq31U05jfSdMp4alzof41pHea4d11ztDPtpkxEhtQaxO1Pzb6/GEXaMgWAFgS8A
4II+8C9J/hAjgDxou2L3lWwT5ANZFqCPkLxbHCJ8Zj2HtVGxsWax0Qf/U/JuNeBm
bS4Ur00Kdy3Zi46XeIyYt5o+CN8z1UAKtVNkUizulX4Lja4gxFBb+ni4UVh6F5qh
7QK8A54HeAwWzukeSFvrOa3n0OZZWNdOvr+7/+Ws/MOE3+MiRtOiR4OIL2mQVqO2
+ikd2iqJfQSdOlH10r4aRKxisKAmx5j3eZYKHLotrBs/DqD+xP8dc1cw6kkOVHe2
CFf1GV1uuI+EMFpo9zQU/6p+7Or2DwNRb4Ya2wqrn+9TYQwVF65DjTVbyq1ti7aH
p6V6YXfY7wLcTsVFgQ+aAljqJZpvPv9kVirCNr65gllxLFuI5LbztTXPzF9+rV79
YdSAupuAwGy0EjRLe1aNXpj+dfm9wJUaI+xpuAeSrfRckdLntvOVhL8R1mLKD4yJ
1ELurRX1vxoNaeRBRZT7U9TFjjQqJRrL9qqN0Q8cQLDNhTR+w83OuNsZfq4CzS4p
Lp6qz45cfwP0qdUP9IXVk/oL5PLtev1wqQOcwbXn68SwDpHJdu0xPSczkZVlkeKL
A/6afgOGFlgdD5IU8n8xwtiXdi5EeW17gOPWxJop/GUqoXGvTWdrLihucDpkHnLr
i6rQuhsdqgG1J2IlBxR3qbLhO3ZAVnVp+UW5v+vpueSqwmjK7jdKOibEJEIJ8Psg
rWtuARop4dfANDeh2njesxN6Du2qoM9VFSB5DBD93LIA5C6Phbv+dAU49x08sut1
AhhxMXPtSlnFAChQ64OZKnautE/O/z/VFxev0k4UHELPgEsFvmUOFt8y17bn1aKo
1m37+GJO0itYbQlivi0QJp3HaO1aIgtzIl4bG+NO9REypryREnNFqu+aNgy2PYQk
bnAaZwhp7exarumEw4ABc78z8h5pU4UNGSp6gCYA/3Z0mmL+levybNeV2GHloOrk
2m7DRK1i/V/ueC0Yxpsjr/bQBjnYi6Eyk7txpzaL1cUzlm8o5uWJmipqbM+Lz2at
PxwWdi3XXHyIICJW8hPPXj8r3GzCjpWA6SDAqE8qXa0+Qt3zvVfW9tWma2JZ2GT/
OSlUZ4TGeOX4yuZhW5U9D/tXwR6Ft1rpLntenRxVbVhTbOYLHG+Ri+NifB6cKkf/
VPM0+rbiENn7P6y/0vAdjGVnFB+1wckcUYN9osf4uqKNm+AoORRjfdeERymBT9gU
+vN7dtJ4VeWQbQwOFOlTdryEBi5SWywcrpZWLFAlmBHhdHa7Z9PgTd1TyrPZa7Sm
7rXIJH6guY8wZVERPJahvxqi8ZbYjD00rO3kMxSIA0kKZE3Q33Fc3t15WenvJEJc
5+IRtx/ucUmzaeMr5MhVgdIecM4MszWAk4HcKA+rxzJ2DQe+Q9kqnSU73951+Cdr
QRZcYajapGSD0ufNel16dhpecvAwc6sqGsYfG/hHCa4AHaCfFl97zWnzZTK78hkC
vRjrT/vjQaRNqmcyh8xVNhqFKUB9DAwqGDBOk2fDgh74UMeuhwNL/p+bxqxwhPwY
C0DO2zRjzzSj0Cv0uA+vrylLgEQxBGQJROKtBQOvOjvA8IZ+yJay9ZN+cisQp7sC
fc1Wj8WvwFLqDaXVinaoPkTTPNc74dfNquUfZP7pTgxBUZumqOQxacnQQ96/COWi
XkV5v7TNZnSqTYSE9QO/IjVkcJc/uKJI5rkBO0XgIQB7pLjxiqBqmEYEzD5CkyrC
paD5wdCrfSjp52Budc4QuUX93nEQelip3uhUcnXjMTyV2828XJFGGohf5vxnMxZW
XaihlDiPqQO8aHMqGnUSa1fhKH0vb722cdOs0LfM8BrUzJxRApVNnalmoDrlc0T2
6AMFPFdxzZpShlFES4r6/RRUXBM40umVr5aVGeFSlPzUs0jQ/jwSoabGYHbe/DHf
MEfCcYla0RBjndkMi4AtYbloDgUCRVspPHcVVnQihoQw/cTAoQ4EH2NU5fRfkNSk
xoVWsyZiHZMpt+ix615A3Lx4UXiLvBByEZMQ2UCzWzgE54vjnL/n4IrzS4bfkva4
Z3noo1Ihy9IOjtUXqLE+tYVEc3RGkrFg6NpzlQvWXZaTaqvMDaRbGrZYykJVxW8w
eHYOT7HmjC9bhGsI+ekjKOw7Op/ImoUtqTnsnfhUZMcyZCfyIJbjPTGJC2roSpEL
rtOY7gHikOGQtIuVdZG9+fq6YLH6XXNPKuboFfr08afQ1udCNRtNIX7PT/aZ8UMr
koGQMVDnftofT70dhqmxKBxgEOMi3+BbXO5zAzbQiXaSvu14DMdCr9bpelE16DAo
IfbHC+l5ZYq5pLH6qyfRpRfVdmUiKeywo7iAoZWJ6B+8wsW6BM3qeuKSpjfIlaMl
bZBip3lzFCWWnYstkgeJGPNrSUmJWrfAErLDrZJAve8WIpcFY7bBm8Ug2VA1vxew
7YeLOv1eUcnUj8hiKgS/LNPQVAQS/yv3BT5sMMP7ahVWhwVMbv3wF5cUgUwQzLQ9
tF6lCuVpKcFTPbqNlZ3sYzJ19YMcGn84y57OuxtQWp9iIsUF/CIVxbq/RnaCytJM
JJeaAra5b8QWecZpXSulp+teqCkO1z1P6d9Q/zIM9pxbEWxtXS94y8vEjmljzeLX
ZWZpNg3P7wBJxXbM2cNU8tDlP5mMsh7Fau5EY18bMtcxkmalKfAqfwUph9+aluFq
F8SdppQiF6WRjlC2tFNsW25jE94wh53tNhWmciC6erJxcoo15i27y/pLLCaqhxIT
a8mlcVM8Tp7KRqOCy1IKNmCz7BlGbTHKYerehay5VfkNTqv5W/WdGzRxf450TXVm
TZ1J4bWOfrcE+8M33X99sQft/HjMDwB1jWGcEzIkCDMSpSP9Xgm8HXNN29RwFaXk
fFvL/mRNmFpKft6s+XCT9AUwKPLntTAP7Ym1UunsD7dRSxj5X0pyzohN5M1jm0Sc
kZj3tMY+9poqx683DIEjcPp4A9appK6LKA55cGxCo+UGWg/5Q4F1BrNH7Ae7EpeW
i/D5HxnnjozTubNSZV6I3M0+X4vcUDssMETEY1wAGyPoTxMAVRNKAFgsUp0VXbT2
TwwEr/afqsWqNaUH2r55Dl219zTruY76Ol2axdpiIJkINfoba3+SxON8AWA+bIva
8RgF+Opf1PJQDMn9goFSfCW3Xy/962HbGLSje+Jq4bXI0WyMuuXpQElE08XJF8le
Pzo3q4h3i4k7O/+6GgMeqtgMjk5Gv5etAgWzuorjqUUjYqP/X6fKyV6bQK3UwUMA
51MZHobi/bklc3MLHVxodj7XihMeK+rLyHXjzrj7LiKnfiy/Ep2YXab54QCYFcNO
KQb7REkI9UbnUZK/GkM+RlmcyovKlQpnrlB5vdJnDfUp38xVSs0kBXcSWwnleY3V
53KtKX9/iPj3TjSH57igYJFRr+wQetNWqS7WjVD1S+Dp+Kn4i/cUyZ1OsEqnjOcN
YYvMpRd1Q/Sylpoa1VGymdanPPr/ACRjztBxedHi3vlqLTJo9cfMggM1IcuR4qbE
SMdhByfuMo81/827H1qXvbjh3acYJVXqoMyXiQ0pi7ROPoo07xw84bqZRPbltlHO
dDmNZp5H/wFNbdPTlC9aIfQPx7Hjrk0dSTojGnL6V3HUcmDT0COQqksEsmeWJ0ts
LzvF9bIkFl/+nALoax38YkzyWKhE6qvL1J2MH3nUsqlz4PRGdYMdWgyewnz4j92L
o5FHWRWUHYQ7xWbksxAxb917cVgNHsf3G+hJchm3Q8qaWQGTJBswSJIrxMiDCLvc
KfZUEmgHgo3c2Y65CKwn+nDhf+wjdy9HfihoZf3bBtPBwUYCtq6cBjzc/Vv4YFTl
97GUqcAAeWVGxDnuUXwoae6NGNhaedG/ld0iNn1isADeJYCHHHCyhR8IAkPiP3UV
+5uD19kGh95pxsHu007GHkgKgGOvBpUGREJ2H6CBSBi/VxHyAz36O3oV8xILK66A
1iUfCkTQWFjinZfplQUhVquSnyBPhcFvwL5LEGO/97vaD4OVWi+Y+AH7Iob1dG+P
zgzSCQslvtJ/wHQc8YsZoGS3VMYeSDA4JfbrehxM4RW/ukKuG9VTlOIibnFkQmBd
1vyuuBvElLFNHF7UioX9RlepV4AOCF6g3sarhCQJy2EPC2nRnNnSnKg0wYj9UwAa
Fbv4rVAsa7yLLALQjtHnYPde+r90OLtYmj3uF9U+banPPMjcSKUQdUod7qiF9v3r
0xdGkyO4aLeLlTLTVF+UYEZuP+32rbW8oIU7x1Jhe+RHTaxa4ZETE+fMNXDjeQTB
u3NdAB3REKG7a5QUucPkfaTG2DlzOxQjAEArhW3oE9XyJOScpNy00TH184Dx3SaX
c/YXOSVWCuXNyBLRV6gTKr5ORlgHtDj3hIUX8Bk+dL4pXXvLstkQLIUVQTHXVuxQ
yR2a7nwBu0tVp8fajHXS7ymT8zVCySfA5+ppAd3jlbg14qJ1EkA4KxvRBi/8MqYf
T1r49vC4gMd6LPxS2ACt85kq1Ullfniq9PIzy5XbEjBU605oe/CJOHChlq1NluQK
GsKLoXe+ezlrmRC+5E3BIapdaTp57iIGBwUcK+Ka3UoM2Peflgv96JeNcmtUH7rE
eiZz44La8tdFRqa0h98SeWhIANzpZaLAFEdrTJK+dVpt2KcdZEnlEUaAeEDTAO3O
rcTCt/nHX9LnCn72FfMFxo0w1I6qTStq86WPBhj6lyB3w+9a3e/KsGbhQoqm+6AZ
MPR/1k+pm1mlcyCv7moGph3FW/fSeh3fHzTUofSQ3vDJ0eSxV7jZH37din1d52IH
gPcR+I5IZPTZF+TOL2s3re4+slQP+knwwt1kynXAYWtqtF2538f3LSbymu71/v5K
oDSb+9LO0SlZdjJT6Qdmc/aoRmcgRvjr9lBkVtPWayAl14naelHQPzQTNXVmWjoO
wWEtY+CjhbkJAuh4uieOF0XwCPOwvvJaG4eCfafIeRCyr70YCg/BFERUfmoS9LoN
6ca7zzbxcWfA7JWEhV0ifAeJvwY5RGqvEMi4NmVZAaMeVlFDl4HJMLaj01zNWlk0
VJ09qhuthKJOpPfUwArLM9aWqJzXABKLggsKGAXn2ofbYaA3WuJqQ6ZzTHe9d5IW
9EqScguT/PTQYXOcT1EtnGrWxrkqj08mzhdxhw1zVRH3wgP/4bc8uLqNlHrkY0+R
NwUZMG16p+0SDEG90zKlVmkp7eXmPhbljtqK24jLKEyb0b+b+JYifqlI/mAI0HCx
t1l4x0Z4d0lsP3uDXLS6oG54v5IJtiuQ4srBv/lfzpcflkAYi99PKe/GsCXMF815
hDZrKBj2RB4dY+WYJWEDBF8XR/fwFnhtWWvAiADMX8vOLaU6Rqsx1qsAwPcQLNKF
hWGByNDxusJQeluABpJmuADJHCYKvlW8wm7bvNPi66A7DHcS7qg4X2YvGi8hsXvD
VSkPH+THi65lOsJmbvOSrHRSEIXSl+pC2qGu3J6F39kaiEoTA+c8Sowdg5xT+Bpp
dtsH3OuMX17UvcVHmwSzNe57aEr7RzZK9qRB5cRVC6JPJRVFUyetKNkPchNR4sp6
K6DD2cbec2QyMi43xFDbsw==
`protect end_protected