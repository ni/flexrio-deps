`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2320 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
cnmYCVpqoAjvPlHjUQ7k1clwjfiLQCRLUhlX/SAGgCerUBQfDB9NLTwEfzrBsJ5r
45fFexAQ4K3SOsLtKhES5oY4KwWHzo+JH4LHmKoNeDoFJsVWK1aakWNY8DKAL83w
2AUy9tnnGSOFUXGWcfLhb4RFpoHjoHeeP1gx8ztI/gjahfp3rDmQXGo4NlHVLMPL
qwCYrnD0ik5/EIquDTZ+SBBe7l+8kw0SJSSDbnVyw1ZcpCBUcdqlvB2eyE6Z2Xb+
NWdQYpk5UyZZBRBc/w9KVO6BTZQQGMpMIuPA0atZ1v71WLg3xI8ZisXiK+TMFKGs
zYvKz68STO9Wg1q8Z2eTym+Nd/wJn9hETKmWWEwwhv+noBJ19yi5yq86iK/qnOB+
ve4FFLBAYB3OBIeeIMY31WfLadxplJ1IMWUQA6v9bl3Qc3MPrOq3l2qmBJRkpbOI
CQJkkblnfmH/bo9zLBJEQ6312QHQ1j+PZfQf3Bs624OmwmztbX49Phk39xBQKSbz
LOu+WlcNRFfmWE5k88NaF982ITivxPr0UT11ZjVs1MyaiWZjDP+a/9L02kJ7Q8zI
TQ7a+6QCOL8wKmdpYzvAt2WrmQNRY7o67H9J2VKIn1E3iZJsXQKWG3KI2KcivOCW
drbzd/Cy76f8cH2pGgX22UjtPofpS7AuNaI3vg00gn/H7La7JqlsoKsyoymvQiin
Gvt/35Tb6ij1xnaL9T15m6+sXpCZXwS8aT4jzwDKysIxrN/jW/qtV85A0yetzKho
spL6+mWpbJmFKhEcd9eJQ95xW1uGaBJcsXPuqXTCuLk0pC7ABuOP0HsIoPZW5kgb
1bx04hsyGxZcpeRmF4Hg88SxxSzzZcp8+H6IHKaQB4SxO/M6+oTtseSmHAof9h2H
NQLP5zbJr6HRonWC341TmvpQReRhvRIqukBH1kfRCJbTSffzeuKKRLEPRiCipp50
bt+niBeNsE00ZS2dovr2e44twbNx9KO9RKO0hgdbEpKLMYVHLCU/EmhSbvsIvVsM
vUOOqkEZE9EQs70K39xiHKuixiIxc1hiSOp1uyPY6m58MUNDUSvy1NywJGNfwd8l
g3jeoh5vgKY8Fok/vVLFy4AD42BUWUNEyXef3v6QO5f9i1ArokiW0MitiFNazz50
0DVqztnHEpzHuJdvSz9iZG41QVgIS4gvArYzkF/5MitvyWwwQVyxj528gxE3DksQ
ChlG01sAT3pvPnaFx/ytfoeoVygKJYZL7yTQ9ffZLBziyIAZbPP2gDQgKDUIAvPT
g+rIY/hovondXW/UNCQD4FHZsXGOHeyjyswNZ0KhYTCGL8LEuQv8YlpXNNmIRpn9
Ct9PpXjXdon0y+/SsTrf4PWFpbWwzpKJ4YF02pLZPtq9F64SHSNLOofoIZTTKvIH
wdMmAOBKFNF6M/vWS3Au/HDzzTclmsQx93mHmy/59/ijO8gVAqSuI4lLdf4GlfdK
O0RZck02OwF/n82fowjY9U4h1zdoSg5lsAEckxGXriPgJBC8F2cYaKir78Kjubrp
x0EkXTu39X+oAgEa+hvQ1HoFazuAMAwoek5lvoc2ibh34jmpTEeC9AivuuaEHUBg
8p4rKiYj1DyetVpexU7Gbu1TwHlAI3ztrwPDY5XR3oeAYkUNYy8KvCT9mLpTGCZz
Zi4vOKUjHjQCBopDJkus8AmjG9fI24ilMHy0ZhKABcYQ3/NVMkGV9lrcWCEoM9Dj
FKyP8J5gXEDjJ80O7WV4P7PFAT1zI8AXtWLREaOzC6bjb8vhOtxXzTbE9KB/MsBc
NYmToXAZ7QRU8gqzy4oLXVgCYV9av5R236Unf8Em1048Imb4PHYgPB3kQ+HwYR4g
GtxaPksOjEAr9eW6lxVVtW49QYx4fQrktz/xljJP0MhoU8wkLzK73HQzVk4ooaEk
CwnYmaN7oJBsN01QZbATPLUR3wBe0VS9z5q9zHLaF2PQxW+3gYSVXt1hpZp4TCGv
HdoC1+dalwtckphQG3TVgTHx/WkuaVp418zafkHIQmgroeKkrbYJWpqrOeElqNAf
Q+4m70fHjLhJDeCf42Znb+FM8R/lnsIrrvl2qq4lCLtZPTu1jSdBY9fYHJfn3prP
NhKR9FnERKLYQoQ5b6RClRqEuiPYcRmgofkBPK+p7LOXOe5xoNr+E7BY319UbB5E
lOVUnpO1AP3wPUeD2bED2changLNVLV6hAAR75cnpMqPwQ24IbcvVct5z2pQMqc/
oI1+4klAjLZpHBc0kkst4FcMOHP+sylAIiSJmohtocpfNT6eoMUT31Pq5VexASZN
yuX0wcZi18ZueBD0XQWvHs3KeXuMyQ8qxBJjJrsD8FapsOeLhX7SKb16JcE16N/+
jFtSr/vZiie4A0jhZ/DBde7hRhBf911l4Ojr3VpBUSSDGPhoXPem3PW5FpCbMyax
shK0DRcTp3iUhKaolh5N1XKEy2WO/44fdMI6y+fnVfc/3Nk23p4HKXKJhkTVpm8S
DU5YNs/BMlMe5wqPjH3k/U8Af8YD0PaZ84lG/eV1orBO4gBBUeTGS6FxA4mDhW6t
3BGtRK11yEc+fovzwjO9UGObQUqDdUKrc8CfpOO70Fv+51/i0/6EK+W4okABeh2o
iA9dnHo1Ytrdu42JeDEVN2sjVJ4lb4aBDAKOTtd8oi+kNH2PDT8gCuEZIOIuIBQE
pFgrdwj3h4FJ37WUFXva9nT3gIU3CY3GAcpMf7njyajfHhFT4CPjxTCVv7Qdqpyr
/ktNV3X4WnmPXqFzts7iHuvdJXqShEOlKyJerdsjoevN+wiX6v4jhBRVofWn4wEA
f/487RamMbw+bRyt4kgmbTyKrAIkfpMOaIdWyKNulyn4Dccz4N1ibcfC1X6gNKyV
c8OSaY9sqD4srOI+rnNox9UWxXGa9fDMa9FA2X3M0rIYp6qJ0xG2vhT81PAebsEZ
8oyySQBhoBARBXU/QU3n7g==
`protect end_protected