`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1648 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
DBGZtUPdvgnvgIFp6VMrQVExUqQNI/iDukVniBeM6I9d12eQ0Okhv/jwW0A1oufn
tq3ddGrgTfJ1qEPJ9BNhAdtjs0uaTMVyRW2dzp3LzcvzddEycBq/u6feUjOf9V4b
C2OZC0mqxj4kYApS3/s1HGKwEFSaixC+UTHDD6RWYwenTlVpVH4KiGp0mn2tG3/2
v5MKTgYeXE1hW4xzsDl+8zLLQAjnVLHNY0/akMzdr08aw/+cSzgW/dqo11EfH7qL
YrcpeKAhYhvvPfmKw6Kw65UfDAjrAej5KtYSM9TZLGi150o0JkEbjcivwlbTU3eC
toTfdjt9NHqp4GxiUWID4m2EmG8/tj4QxyYifOqwQqz+zF07t6ZJlNMgZIIoeqro
nQA/g+kuCeJcO2YieOJ6fI7Tt8DM4LlkEi/CBfIh+k3Wq1v9BgnQPT2PohTf6pt1
nzyyfydYwcOJcIiVu0WTlh0dFNt/HRuO/k5eaqCvhTIv1H2RYB9V+ynpr6OeZWID
gjNcLa8OThm4msggrJibnDuNRHlTmvaxZDSvV+OM6qJgcfEsPazFnlTbdXsqz9bx
fIkb7JzpmJ1s3pdI9wkg/AzRTNGMjkab5qAD31il9RjyqLPkvt2sK8Mb1AkG4YCS
TDq6BeRxTx4cIbVCa8Yt8DaCLzoWfr5m8HnQtQjkldg4kpxvWT5uQEqEEb2BMIwk
0iNT342OhRofLIXqrk7F9fIZX6jNkYYOwJb0l7JiUOFgcSUEX7Vwp1xCpNhAMFF9
3bXeOdZfRvnvPgys5wVBTayZicm97j/wgklQg91VEORQSN+SeMmu9UBUdrY7saCc
Af2tio16xc/E6sHWgD/SfkLvmiTz2MtPxKb+6IHAUY4MhZrAqLLOcQbh8+837wBw
pssbc0Jax3Bwlh/rip7ZtBUmSalBrGt38ZeyNkrJbccDFA0d9tR5JzYqAnwvWBBe
/dPj2oG/5YiK2cQGFYeeXJU/oTyXbyyz/LQHBcpZA8mOpNOmQ6LKNOkpgSFbQFw3
ZNHk8K1od52rptDTz1yt53r3O1tCsLCh4FvHxiOw0V0r4dWxrRAj5TCgxX3hKhwc
L1n9D0Z4mnBcdsZYDTNCDxOHgbwV7avhQO12YXvo7YbQnD5bEafGY0klncO4FwR6
RcGui0nrFqagAiGyxA+A3wwC4ijLHkqjGjs3WaYdBvl+WMkDKc2U9SvTH50LmQyX
MT3A91z2bNMfA1ubrK7jC1sUQPRoNLBeJp+u3LNUBf/vXC4vMLeXKBycVfB+DaXY
/wYz2kMHZU3OeIp9hNK/qTqZHctRMtNV0RgeDDTXGKVdhtLPNN1zo8mBIcwOxBAt
NeTlYVO0ciAw8IKV2Lt2n9l8CX95Fo3Oh+fAAkyW1E11+Twr4R5OnzuTqFA3bfVl
wonzPR0QU5Zyw0TYfjghxuOwoeB7CWGzWSIBE3EI0WyTpLospvCfOoHuCYE282bA
yjrMsPcM1INdltIF/OcAiGIM+DDg8yQJq5Un7NQ7UGrxYc6p6VAXpkQj85wr93sL
zvT8pJZGZwP1a2jBrOH27mJvZeYfVnLXyLkIyTnvwfD+ALdLb6Fy3e3ZihEfX3eu
PGiqKXMou7SVHc5fcnm+S0GHRuN2iVtWmd2geXM/WmnwPgZDDh6RnF2ilJ0m0n5Z
DjjYyMhy5FWcKusPAr61OVllbncF4KkL2oT9Bv/3Xph2SWxaMleQVfGXr6OzoJQy
oNo7QieTBA+xvPmkxgAh1R1+7sUhENtCFDs5LCnLJeHPxdbbOyAiNYSZy2fGvTqG
yfJCFmdK6M/79crbSeiCGzckcRkCNlXKDowbp0xB2DEu/DSCdBQv6+lt93tTKrY2
dc95fKRiw+e+2wSaAHX7wqeaCY2DmZfkWch7Ys9B0T+RHZgNiNZxz47fONkW3S32
2roUSgpSMHuOJpMjWR4jLT7910X54LqBW6Kf0YWx0r5fwITEF00NaeSGssZgAYf8
gM7zanHq0c9pkAW72ZuCct4A3T+CcOOShWm5E/FA55esgAwp3TSm30xlYoIsfzo3
JaiijGzfkq0IlWIkaAhItg==
`protect end_protected