`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2992 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
/8dei0SfYi/yIzInIePi3Nvwk9LuyEjO4gJkIP6R1GZkRYI0jWvOxZHW93slidu9
/RTGZrEJkcCw3UCzVtEoiUKse5wlzK/GSIHFZRtyMxafPLd88Rs/9z+1Cq016OtG
whTiYynKA2CVB/IiW2yPILo+2Sh48hG0xyvAwklAbCjv/uOuMwjGVC1npxRbdssb
mTr83h9/58/b0dhNzbyW9VzQedSPrpCr4FfV3lgCXc4NX3GWUuQW3S+TXO8dHRY4
wTEB6xLBWpn66x/6lb7nhIxSH+9RRHjBfkTCCXJlnnii1Cd6tYcUH/Ql5QfTVXMw
zNLmvLkxA+dm+NtFKMBwiLb2Jdgt/22G/fX0BOtz5edTLRzxzplXHDSy8sieKsHV
LD8p80DDwg2cIdMUfdG2IppyppM0rjnlQqq78nPQQyEj7v5XeQy5aveoO3YY84Yt
L9z2UFuZ1jYGpk3mn6D7jH+QFikfziU87D+6rDXH4JuTbijEO9zCCO1Uk3wiljW8
f4AY/agyU7ml8iXYa8fq3bIj75YulYeyerXqmQcaZi8735tWYyDdriWS1eMnFO2T
BksfjsWDCpnP6tpzO9UsNWN3ca/PI7wyCLHXpCCzsodyAQ2H6Af/wH0LumJhcWbu
f5+M+0dfVvQECCAUvtAKhf1zSlQt+KuPAPLIXNZO50SSP+YcBBz9S91jUioFuzvg
snvSTxRMcmz7s5R+ESy2t5F4f4DeHZMphAHKg6iWoagzmbJdIc7b1WRvchdCbmmY
2ei6sulgcpXlamhU23y88Y2o+5SL7070PatVkm3Q912DXBMJGPms7jVC0mbhahIH
TTh1xpDsk1/NGAXVKfhVNqGuogN+hfyFcT8PUSVvcu5SQr0dtvTeOUP9Y3Ymdiik
Oo2YJAzPvKFLog5PL/zBj5LWuS6j4zwH5IDXEw+9HeKiXtHnhJSQijaIYhmeQhb4
NX7Z6twg7UpzgryPKf5DJ0zFRfb7oig86jVsxg58dSsJ4NxyjSzjoGjzsovPSToB
fzxAsIb/5CtDEx9rmqpLV5x+kT0WHsa+2H6M7His+fNZ3th6PZcy0pOWUKZnEJFw
FGYmgp2m7qNDQAdLdEUP+6jeVfum+T0f42dDt9YwD3ikfE1rqS8eOCGJOwvzzqyi
voLZT4XUNlmXgDHEJnhFAuLMZEfAlDh0Xso8c5WgFcEFIhjZ24UMYHXNg8chx95X
vF4gGkuS2glS5l5bNtqVOU51V1krMZ1KsiqVM+9G/VlJJVsUjYHYnDhmLhCCK509
ut7koZCy+xDIL88uEuhmjOZqmhtu7y9UMcGdBjYkHYO1MLK5WpFTaJtY4Vpf8ykE
wqCl2P1bOaDrs0jwAvExltIhtXx13P7d+RL94vFQH4Cim1DTXnTh7rOGvC/965oP
E/w04BbP6gelaWJ94kbbn5Ums1+Xqrk83mrmRbjl5+TLY0wyPv126L6Rhl/2fVsl
H9zsOuOcZn9tdAfEMl1zpGdesTSOfndMXPNVwnATiWlp6niHYB7rLYjW55CRoYVH
IlFAzjnWFQvWIi0hPcOLu+fu575YwvIBtCQ2iyyyKjYhhhjL4Uo2EUoOumOKPj2U
AAYblGUhoPkO9c5eps1VHnApmcG35zJnMRgzrCFaQJ1PtBFAWxMloBuiVaLuUbxh
DWppWhr+GZwfQ74YYzRG+75EzuXGg1qd7sIsMNw41rT9lmeQkKy8mrHVcKjK5qSW
xF0ziAQKSLK5w+xbQz/K5C3gDjkB5N+p/yvuIRmA7Qa8egHnZW9EY4CwmHmVYu6a
7dORHN002EcCPJrbFj9zL3RNg7/io3nfoiFKIwxFUchPHnSfPCL1jr3guKOui1FZ
R3Tnzf55DRlx7rPpY9YuiKJQzZOlriREFT6Gx0uHU0vuuLRRyYbVRNiOPM3rATFS
GWgd9r2SFhRcYsRCxVbo5TdKCuky6xUUpyIit7Kf4Sm869/WdkifScS/7dtTWruV
ZpwSiiT3ljEFqLzTCU7MV/Tc+q3XOigkfJfAY0uujSaeOsMrMeBhxTr9jIs0WJBp
4/51gqftOVGT7P9HQ5H4+l7f1B+tJGw+neCp15fgHC0ZlsyyE8IlRqzYH+Nkzzdh
4G0F69+A5kcFYPDB/uIH3h18k+25PUs7qC7UAeXFHa9xIw/ob2vC5qii9O0r/m2b
JeTJtlnF1QzbSfd1/sKzjOdtlcwVo7keoPHU/6rIXA+r4JpZ0ZRl3r+GWFu4hAaJ
iJQCej9P2COI9p1uKNcCADAq+6QdDwpkl4Dg160w4tsT6erIYHsIb+kyI4S5vDDx
1XOydC8w6oceJ0xTJ5PVF1/jIWck0oDZGThNuf1d68S1jZvsEaN9SfQIFD+mnpfV
Ak+QlhU2NJEvPa/csvVPc+L0SVEwOa7mSpViYbvsWPXbSxSfsRJMiblp4i+j7DEx
dunMChz5MFSdLYIGCFELLQIQ0ZeBcQek8kQSAAmlbDS+HXCiM3p4eGK3WwwMEcO4
TxyeAholcV+6hKFmksyBkGE5+8MlA+xbdOFYPs9o7tGhRvmGl8WLoM87IdVO7XFs
j4qhhpSgvsvprz94VSbG+69c7zHLQMlKuIeywUi7PQ96iQ+MfzWFbwmmYjPM0Dqp
qXAIif8fIfD7ISKgw0mkOszzLXRbJfHc0yV802SXqd+F3f1JsymHlx0xgm8LWFZu
Sk+rXySUDZI3pvCUr6AOU+XrqaszJqK7uUGew9TKuhCVrtYycwIdNoOAFLchjdq7
HZThXEyTlq3cAmoLyTZJ72sxdHPcgqYlu/OKCXtqg211vsFJHqa/7ubG83RV7vSw
wnlSJqER9IvtON+L4y4HYIWJQqKt04J4YpHQKtXxgHsXV7v/lwzlA7cPCFHMK4FM
j4xhnDWQwwMbdRvr8xVpHz/8aBD9wzsePxKE5SdS094eWR4LI+7wUQcUMK8QvJCU
ncMHS5jUdcKj7pVj4D0poXDw5ssyWw+6lSNCY8s8K15WiDAvHkXc7FHH02bZxDJq
FPogHm2x1Uf0M75SYRLTYJXjR6uOr1aTBinc6JVWSvuHUuIgZ2Eo2Pee+euXIH9C
mGjNZGX4c07bGv/RlaZyNs+lnccQX9NVtwVqGh7TljV2PbDnAPi8ZKUnOhJojC9W
QnHvP/edj1HKzfoenM7CM8Q9676u4eLi3Gwd35wRDqgoWd55/ESOFju3PiPOPO34
1CrGBp8sITosEEcNrgRW5zueYuWKoBobfO8yhOU6fXutMB1LXRGCFoDP5bZYl9Sa
xbHdm4WB1OoKc7VgCD+WG6hbvDgeBKPUbsW/JpvelNU3uZ2vQTxXQZs10VVKjmXW
s2ePXTrr+mb6kbYQAWO/CRqOKJqsSn9VijPHk1TsrULTpFo32KsMJ9fu+t0kR9zX
kjAfpjQR/U2SWk/05dHV0+yFmkeB81SXVavNF7LXs4+67hW1ITxoecZb85Eir4Zu
rgUO0EyYK+A36R/C07RWhS1xVflCtQsBpL8svcdv3IG4hr7WdOM5vhfwnuJTZEph
No48EBDsmAXv7AFUrqgTnxs4Ymn30rNn1wr36Inm8pqd0SJHF+xQAOVBi9Tc2KSR
0F3MwKJqhqjQP3D3s8WTlmu4h5+EPlxkO/yqlk1TOye988Jo8eu9PLRMvO0i/lsK
KUeG1N/mmWYEMukdUoJtsmQciDWosPnCLSOwHtDMOaLTbNgjwevS5chAwrmGZa9u
64NkCJF688FZvLZGSpL5EupQvhCn4/IWN+0iFtfPmMgvRHgXnno+Rtw1squ0JzaN
+2NM/LdZBxRzbZfFLNGLgNT/o8FizyJJQKFuC0M4cXt6ylfg5ZIwO7W5YSapRKAQ
M1pFYEVVCRZisabQSt2PQg==
`protect end_protected