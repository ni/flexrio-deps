`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Jm2uGAVYfY7w9Y5qKstopObZuZAEY3b/Io3MSEcWLhjjnKulVhCBBYAEQrAzzGsT
vMbffkdZgjdXQUg8jOLJXSHZ0Dgbnob2vlppjZs3bgyHCF7MoJ35E+LOsaLimUA7
hlqStcK49hR1hdeBPr/OwfT3UeVrRtQyq0eJXQ1UksinX1G9Pz3/CmcGfTZ/C72x
p9icpt0bkY4/1I4GBvNCsA6FFKH947JqH27OPACiQQRW/K7JToQn+1uhWr3LA1od
lbVrWu8PdZi7zW9gK3jiW5GaPjwbYQGqeGFs3bTKBILjb7sYHxfxw7eDLVMAIu5D
W+OTIN4JiHiE1gCnNEvkSQ==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="pm+c2fYA/4JT1uhlJGVUubML8hZi8lME4xPobg/m8uM="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
nBaXksR//iZ9fraC7WMJWWSrjqRXHxmM1Y0+KKN3b10NElDzVNMlR76DLrcnamFd
2n7uzsxWqhhJR5LBl98SXO3Y90J6BMbw+OBG/MFM/zUulxh2Si5YK5G9GCrG9gvZ
5JomxuZFDu9CzlWGTuRUt6FsE4Lr6sOL1P+hraQDpMk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="M8TXDiNa0BVMX1P60yIvW2WA9jKGGy8GtbuPknDnC9I="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
/5TNZvs8Nu0G+mfp7M8H+iVAGG3Mh5DYZ0Gn3rRNhV8b5CcJKgjQajrRoGl/gSxp
rBAhtT8Vd5eelHgtvBjpvFBA/EBUrRH6CG6pqRt9r2qUDt4UernbZbxC3BC14KYF
gLiaAkKLdB6NWFZG4rx6ah1YPUP1XmKxbm/SMkFY87Oxn/UMerKfOtyntLBgfalm
b6mbqmoj82DK06jd4OFCMm+Zx9t/Hp6Cs1ST7DsptYDfIwGbdVULYFGC1QpwAHWg
Sho0c7nPzv+fRXjwnqkESa7PRpBuQU6TztVKtRN1b9xv+w0No1M/+i1sWknqwUeu
4OBYH4x3GvzTyGw40ljZSgQf9uRrp6QNdsmlAU2yHxJSfpRdH0Np25sOy2g35ey+
qoWpPy/OorP1Jv6k+yD2vs4nkM8X49zGfYNJEzpRs/EGuxton7Nlx/v4ozSxzrmg
YpVneIkrp89oLNAYuI/xIYI51G1YGByDTC18wuNmu64SWQKGl3UHVSGP/+GLiAis
xJA7kKeSl8PKAJ/+SzLUAu5j1qBaFHq1rstCo90XEecU2Ip6BtlKrCc8jnpgbjmm
8OjwyxABcTNWNBwnpPOGnkeA26rdTj+TqF/s52AxU6sBNGifVdQgXQ2RaakAtUtt
a8opGZ38x3jMd83G89lMf+36YrlXB6oMXHySJrLHOiyhwrC7CmbXtVe4+CpaqOK2
9xZjKYpqZrzf9/QaYbumaiLZ2FveR7vlAbDnwNji6EPz9n+FkSX7zuPdHvSb3sEI
F1m1/8Kq/ICEWsgkMbFZc0anzAeouD9CKf8r+lzW5IPG+F10NqqkMZcEMt9nBCNL
l81klPnGct+evzW+uCuySFExiYIJPQ32qM8ElkUgkYmcPpVD91cu2OBFe5otbSmH
9l52jwqRKddmi5WUZeLTK4RBaaDIcaDmAmLPFVKpuiHql3k7tekELkfK/+EV/V97
qBIoilmQwW29m26yy7jmETRg/s9WhNb7PUuP2rU9+VcIIEQJep7GL+HIoQeFg4AR
m0ae5UGNJirW052Tu6joe5bxGPuRgF4VkBq/G2qetUzgr/KolsBOdCnI6qSGQT8U
eS6WZ2ctdPHScb6IH0p+zi4FyVuCzzCEq7MdzG6+KUo3dXaLqmAsN0UVv5AI0jss
YVlmX4eripFNHqRtgJml189OH2vFmBIvRreZ8yU8gncT0FmMDfuV1/bG4THmvwFI
nie85N3ZaK3LtE0MCkgQ+3PEbpelYIy5MAqBXUnvEtgCTOqK1FdG6OTtBcWAi0Vn
zQ8W7ldPddU0XyEPWXvjM2AbyB0t/BgSBnLqp8756tjNEbys399+KVp/68Tsy8IV
2Aw8phTlptuOVZuo27bqXVWmYHU0bfoB6woLqckfkdO8K+/t6mUSRXxKsqDyTr6c
UCDnlU8pM2D9HH2NtdNbcAXp06oO4lDODvfQqnGHInTBB7NDuNkGcG7B8N52qZR3
AX7j5yaU9dUMAJ5+GsVooy1NJS7TQlPDTVVrIJA2vZeY1C8hRsOTxSQgrPNmafC7
/GZvCApZVxQGgCfHaus3sxg9UoFCy5qDALDhrW8fKO8aBj2lp0C301mHKhG2Lckl
i8NCeG8ArqbYe1mmXzTQuICDEICkqFGzCf3xKHwb3S1GINhdMRWNZZq6jhgG6gdG
KHFhes2kBkJZ1d/cZ6bJLeq6THKX5SM0M4618JNI1rkSu3JjuR+gITSgZBFPcYJk
f+KBwoSItgj2pa9+N1Wjn9p2lo6n6eaj1BHL+kVH4sonJh+xMv9W5jnvhzDbb+20
ZmNU2Z2hKi+KOocIjKZtO88KarXXVvWmNWtqFXLcYui5T3lj+4X5jD15meTH5uIG
ql7f4k5ffwBH93fyy74EyUbtTS+zdakpCXiJLG2wh6CnBCn+VurLHd1wt2XdLPJU
OqRCuB2o5jMASmPZUVR6K3c56od+/WewJBtlC8hj+tRLmuYn9yykYULi2yQvQAx7
7hcGovG590c1pMo8bktZg+IbMyBOeM6Spu/ffr2ltMhvRer/yOD7cQ5bS1VV7dg5
XFFndQZWTyUYSZDyscdMM3YVm8fPu3tUUn1S1Ix+uw3DfMhNjVOnpnaoV0/W9mdt
kFnINV4NdViWPJhWoIio0bKeGmZ6/Z0pCtRss0QDHfPunofmNblDUqi+UzcLCeQV
8tCKAGB/hY/bX/PFITnXPHT09WojLWW8ZqKVHrTJ2lYnupuQYLiIJQpuJ6o9HVVT
7cOyaXj2veCqtaNa2wxcv0UrwT/WOkrp7q/9nThi62oVbbJlFNQJEdxhUiE7kAyi
WxyBGFD20BP1JX8uNJVp3rgpmfMUjIFtzWXrZQR6DF6gyR4fs8VDXfmDtyiAFy83
qh9wWiOqZ8/m5G8Xjl6mluFaFhMKDO9WlHe0FsfPPOw03JqVJuqhFex3Vqdsfdnm
N82yxt5ZY5nRDIXvemEzM6QOEBxG/g6KB/Ygis2l9r8ELM7CeCHdspg1WcTDYLHS
vClbRXz9NtWNyJXxCRlEUzDyjjGbrKkds8qC/KYweIlcl+Qh8Un0re0aDj8FeKcl
hLuuMr01vAKwJWeKAuoDruY+Nc5sLkP5W9nDky+EB/ackSZSufCEvG1OXIKKbGeE
+O2BE5PRKUN2PHAyzkiTrz9uep3DS71K0D85MUKte/GUEqSV59XurS+YFCqv9ftD
ddvRUBSeXgWyoo8Cz3WM7x8htT6glvjTNzdEAsF6kIBoMkUGaak2aL5TOE8K5pGN
IxmL85GjIBxuVlhpdCV19SBJOdEdoQrbAobABc+IE4y6YohzQ2JcRIoxy+2Riiwk
3OhNqAnJ2xotBkWkVspT6bScxP0X965wb9A3rzEsZsUszcF2CvC/OkZAKqrvPt1g
PNYnNl67YPYg8mSJ4nWbDqhYVsulNosLkG8Qghev75mSmEoHFcWL1ZfR9EI66Z/3
8M8BXwmeT4pmod4wVMhJ5771B4RJSGru6kNVLNDA97GUfNLczJeqPbw7MmGChOmx
hoJ8wbMFSFdbUDfrhyLc7WYi5aa/ovzM5q46LbZP+Mn2d2Rfej80cSnyAJ5Ykqgj
U+yRRtjSof4e0vul+zcsi3tNgy/Z9kDgM5H04B/MxhqdSwt2cByhOORd/NBP+4yZ
BpWgOrwMFWeNjWhjzzO9kgl9tvp+MlNXh6KNBvs/1xHpHKXUAzDq9627Sc4yJsdp
9P/172IwwhcRylUgw7LwD7jCjPO7hQENeJeco/Fs2zcCy/A+5Fxx9yQG9o/3uaCd
VYBJh6m/ykWl/TYSM34sTIzph2FuO/uUC2kVzYsi6itxiJ8FNqdRsvWKTTpP0O1b
s5+SKbitCm2+3uaD9nAz6gaegRwbQVb53KNrvvlG+mFvK/QRTGndXW+EXhvWzaDb
RaT78V3OW/JWQRmKJxZnypCYTCg6ushm07FHOC6G70TZUdMMw3xgF07+gqP88ykL
vOHrICqZA4buKZOTV1T/1sLTA2c9BM/15xy+oAIKG1nBMPiw9GW8s1mdeFJea98t
i+pYII5YYUU0bs4Yp3/HJYosoAc61krl1YVq/y/QE58Lr+kE/sbWOgYF3fb/9Nft
cmpp/wSgy1eXSfqWvBDKCx9JXYiRr9f7N5HIp0ltKk1NgVXF5G2KWSxvTdHON8Bd
yK+vZCVEmQRB5w5Grfec1p3KBWmPfhQ8Y/s1yqs7o7BvIhIc9Ncd//zPVSyFhE9S
jgaVQulCYkHtDyh6Cr3f7hK47h5KdSM3ArCTh/eBQUNcu7jz2OORS1MRites1xd7
CkdfkXPP4NZ9zaOd4g0ZmG7R6F0AlViKTlzCEZ6rcuXyL3cEKbaospI+INs+H3dJ
d8sprcAOLNaGRlF+QrejoKz4Gafml4BVM0PBaU6Vj/XG3k0KL9Iox/NER9WhF/Vi
Pkc+FBo7hMSTTKg1TwNd48XUx0ucp0Vqpt6D6z32Af4PSoYThHRcPemk0iVa178M
g0hgpF0VJ4iHPIPNyydx/OD9+S9nMS3tFP7EcNXJqQqGqg7mF2VAl5HrZ4ESH/cO
Hr1QJZ4GNkvNO829ub+9NcuZ4PV4sjnF7ME4WaS0MJUMN3I+OPNAnn8qcVPL96DR
k8cUkKzF3USAqvi9ArjjxknokloatQhBSY+nE8Y98WESA2v7Z9ycT5tfLB4mY2lE
PP6qA8GCoTu+TC/VvC2X2MZMVX1hfaVR8oJYBEU1etLVMOn53iLwfqhVL/1nXPFL
E3OhDaGGkqSJv+m3Os6+mEDncESyDZGINxNEhHIy2sxok7NVTsYVK0XmuahQhmv6
HbG9/J/pGs9FSWQgYl8vke1oOpwOrtXp+OZU/FxH5vsJQZTOnZGtHELI9Drth+iE
5ipETf2cwyT2jnvXZZ8cCjn3M4o0UUDIS2FfIQ+gktUbolAOa5bljv40GTsv02tc
Mu0E/0m0yAogSsGEcYuhTbUXovnTU4atY2BN9hm/lVpLx2jQjwO3cpWZEBMT4vhU
9EfzgtSGX88CqzhaPrfiuZJ2dXCcBgm6AbGGRZRphvC2tcb0CKeYlBzvIYVO75/M
j5Gf8yrfeSwkIAOdL+BjYzAMOJ4BwAlS+yeYzr/1TFO3CPL0i5kXGZ2N4gU09SuS
6lm4E7Q65NiGELqhE0ti41n8lyIw/eUxSKQFrpziv8MV/YDOuPdE8GuexPTXJpNh
/AjhELRLSRgTmyhKKMcAJoBmmNf1SPoR9QMq51M5ckykdPb6fcHllZ9VIhAB+9cr
Z+RLzmdaPsryWOs9i/6cc/0dkYDLhiMpR/pf69Taw3REc+9GPNHWEWYu4MxA1bqR
qYs4H1B6FLa/cQoEHmO1rk2+a7ExHUmakd21om2cb6iWUQY243izVoeGM2tX+p4h
ShcTBlFlH+EYHrta9UAwiPsVIrAld3b+YyU1xQ8tqCaQVxu9rNaeHphZh6DXeC06
3wDo/308AvgrkLIGVcy237RTipixD/nqo6TJnZrt+6InBwB+JBV4N5Fb88GMCOfa
Sivpg22/yX10Aw0BdFBu9NvybGSrAA1lDJtlM0qXQmhVyxe68dFZSeMq58MajYAi
RX7+p2VMAUAD+s2Pwbw80QnbbQDkBquSHCS27WE3HgG8rtLerhCa+Ot0sr0E3Nld
XvwI536DRUr3smZ+Mq0EJbbUKMKd/676ApsPm4KXK1K9qVv+NPmszT8fLIPfG50d
dsrtBAm8aJfqWVwWPCyFw8p2Qz+KCuOoQdq8cq+fuL9aUg41G2RwHljjNgMWy5HP
q8ANQpp/trXNxY8aHh0pTspK1QDcMa4AeEvBE6n7iPnIqPUpm4f6yeaG15x4WKaC
egTyrB3nrxIc3doX16A9v2eyZFQQDooSYCwe2NHBAdulWm2wHLr/RS1YI+zFOB7p
+Zx5LDuH48K0opP9LwAmDaab9AiGD33vvY/4InkxFLuJUc4PstCMwcSM/3zKHLzY
kxff64chyBn+LGU44Nsz0UqzgCgKaEiR27KvV7/v+BqvpK7SIMtxYChcXCi+sWx3
cuS4TUtYkI9nV+2rpggOrk990UQj7Lc9rpKbXFPnz3Ot7nmgpPwBfGb1ccDnG0F9
5XcRIjU4L208DPF5extuR0n0o1H52vMJVOGbmqvwfZNaYgiR97XcVmS2gurVzpJs
4A0Lz8zblQ9XpJQGfoZdLZNaqmnlv2ZyvndweYxaoSFI+5fdEi2OA+giy55EAE6x
CdD3LpyrbmfmFlT6PahNz7DoWC4lIUkfOdr/GnfKw8x7B1PgiAS1XpiiHUUmxh/p
9MZpkXd6mrdTujY7anmJDJvd55H3Ixm4Dz2xoiDVWhx/RlnwTTx3qJ2GXQz0Jq9g
lUzkVGHQALqvM+iQm1iksTReB8nXwUJpcktYjBYlZqXLzsLOmP9RYsoS87qptA0R
OZmhtJ1qRmf3jWB2zL3LNnpbdgvF/zAcV4Dcr2tJ5JGg+a8etcdXz2laLiw2cOIm
OLXEWc6LbaFXiiog9KFDXgDthgjFyVG0ju9WIGpqf0GDUFCEtodIQczModMajLIT
4wXtSu20v+7zwmOZ90lNawwdIxr/MI06L7hDFh5q6tvHl6HTQy58VxbhufrL85yq
3bLcUsxbxru5CzFWt8Zi7sKNSf4+ysI5I+6SwwmW0RGr9UqeTBktvyc7EFHNvnzX
S6IiVTNLqttaBFnloOoC6WiTplCfsFfy7LircW4WUrC1eD4eDXCkIItxTOyJy6cv
Uw9RDDghQ9e5DB8gh24Ks1wbi/GyAv2dsA2FdcMteCaeu5jIexWPpbdzwiasE1Ky
xwOiuWBJ8CLBEbeS0Y9YuCy2qsUUOxlbkkPoNGGa2VxbO0KTwp1jNWkAy5vr7FE4
/pJRDY3eO+UiZHZuaEz/a5YOCQG7zmbjQNNQiqVx/WO/MZ/7+fKQiibhhEJHsBgm
phZSMzBCMM6+nZGYkT9ChzUCq1l7CWIOTvud5kw+Ij0yP9TVz78eyZ61WCoMstUu
UIlD/1xTh3yEALejk9hu9p69EE2yqwOtIgwX+HkpV95ON3wjT7wpoOyT+UtBFV2S
ey7jBvnuQ1p5f/2ph/Da/o/RR7lVaC0qNslbrQ0HMxfdX16UEjJNH+4xStepSn0v
NZq29ngd0lf5fw3IGAKPK40JNDQ0ggToWYMWNEdqjAU8ZjpFBe/SiJTUC01EFsDL
93u3RIiIre5slqIAz3twOBD24hnz4scR54SmNdZeVzLHqv+UcBYbkog71tSLQB3r
PIQcTJnfnHzYQUaZg+lNvRh7BuhuthC4jG8qsPEpXXsNfZ6mJmIpoKafOL28SwCT
8ncicxXsKGujajUv4jYUzyfCo8nCYjGwvkkbhI4+u33nBovfhhMx7ITt+Yt4H/XN
DCKrLgC3M+Z7hZb7eTn+JSM3ZRdZ+yLce+AagTBXCVEO9NmwRtUKL0fgUDFT4o1h
lm8YDppXPH/sk+LEciDdFmGYTEQDBiarw8dkQlgMXMstYho8U75BRcnb432mnA1T
XDRUR7IvQWpEl0X5eBtdr38DQkAqgMQA/1uKZBia2S2GSYo1Gqr+x82XpBRgnxpi
gMv0UEo/LJ9aIc8I1RYOX8eXT4hlXHiF4PHt+PGhVKHkzmpolfNC5u8zuEAUvY6/
KSTV6/EunjAA+O0DclL2a83Rt0YE4lgt0emeE4uNqGkvqaVvtWrRxfgUAbA9Er4y
sf295WM7TzP7CcPOVlW6xVB9YZitqKmwbjzQAgFjfVfIh7069kaC+W5mVMeLfKKx
oJa2pthw2wDQxPNfX+nHeNLNt6URCwtP5aLDMG5NCrA90YDfvKhCADjuizbX6aUE
lXelJ9GX5BUOspzAVsP+0lpxOVgdgOoY4gmxrPeAqGw4BxenviiDnVTvBAZpTW02
TY4wMXvsU81n2ilbxYFfxjuIx6l2StCBbdsKQTaTNF0XAqg1L5fRlCEcRkjxvbDd
g1e1EF9sDnc9KdCo76KoqN1Sq6lQyhpSpJ8rVKeZA0TKNnm+RIkhJSpjPVS5sWHR
0aJB8PeJgmfAbUNQ7g1SnhRICVEU/IE1YvOCadXZ35FLkkphKi9FUxl4svL+njL1
6Se16YFd6rWrNAqLi6mEITQwrkLt+DTApDQw82UX017zgJCcxaGrddecDP611yD+
edSSrXFccht4WlY4CJ0Vi0ASdX1djHfC+R4kOAwwccBfe23YI+qUiP9kQiVpXUml
bVqSKkGX+LJBy8WyS+MS0kfFqMYhCoqi0DckAwQLxaiY08DdRYvQQv6wg0VY8dnp
zgjhr0LMnjVJWXyLIXi1KqHjsiatPpxS8uGk9SC8OpAjmL61hu+7mdOQ6jl+Fae4
stI7XZDo2qZOXJvonZ9xsGw2bKSuYc/WkXt32T8Q8n8KCi3zijITUdVvzrkKOswe
e7iL+CIWncpg44vxOplOjMsZOMSAmyVfljXl4zNyAK026Pg89SDjxy09tqoXZaxC
rRa3YtsXJLm57v9lt7xiRg4gEwanpbo8/q2AQTHyu4TY5hREXlWhl0+e/VvMZB9F
TwSM4Fexd5E0EO1o7Z0opkVnyYYXgkCW8ovxRMQ3gQyJICUnGF2eVYq/1qb2XKip
o3H8TNO4GbORQ7VuphAkjDhJjZKG4fDAmIMbWz1vnGTbnW/OpZLUb9n+gAZjSA/z
sytH7qRj6/pBy4TXfIBH12w5CfTV6z9EDP8Vwc6DIkUJIRQix3a3Uq/I5+BYbp9h
4ToP0+Fe27JZtzQUy5U+N6OldDPFSBj1yWSx2BZQDr4mA0shEx1XXsbi5Htwh7As
lP6rblTPT9Vm5KOKH2RBlDag0PgVYhJyXpmuJZV7fOo2tZB5oeGCryCNFEH30uDo
ztV+FLcD9APDK8tR9rbPOyzwu1/IA6FSYYJGFr7/PJE6uy1Wog6RFo24N6RNYy3/
LBND3JUVvSVXU3+XZrHIFtq7PvQQeazN6Tda09BOXDkU0vM9TaEPZohupqCBV7Wp
vU1L7x+Uehwv5FWgX3mn6wCZa9UOASKQcwhw24Fg8qCl2vSDqy0e8ykQaaNEXH8D
biv8wCs1h4H+bpyVxM/tftRWSKv7NhQWarmqEu0uQHnf66FVwY3TxjWv/m4u/ZlS
yBTz2HZv+vVKIuG9OZTh9X/MqHJcv+Rhc9Lchcagdd3nTOuMPfTSRHxZvzBDrJM1
SSsMnpi/EemzQatQh3UndujfUQSqw7MluOq9Yt0dUZDUtjI9qPtU/nnZEGg4dc/1
oWYGiaIv0e1VEp1egm9FvXtpQtq6EVnhAqDWu20lnaDElI+QkRyfSIivZrYZcCHh
vWLXKkXM/7CdiozeHhQDktfl+y0crwgI0fZyu+LmGe6+gFOqyVD1ZRMf2AaWVAZ7
7PRjqEFGhktEKuYDM37GLzQbJsjkXzUzMarmybFMVWWh6+k2/xKgiVxFIOm7bpOC
LFxY7fnJn622ySC+rU5gHTCl8b1CpTcZQEQPz/O1JulUIcJeNuFGNqECUQ5rT6OM
XCaMiuOQXFgHmhrgcDCmAbSYh9SqR8o2ncUfrWY6FoSqQyWkWbMd0++2GRhmgm1S
y2O17OTkE6jrtGpx+ciXUDh3WNIteDhIoWuuXokMjCEaVHrSggv0CplP2p95S/rB
vyWg7T2u0Hc7VEAc9mDn0IbnwKnLGU5a+OLLB086d30G0ebKDg82aDZWC6pKID/0
eJyu+vcgVndwvCUkbxuz7GoWibcQpIXBICiqgNzHKV78qOGc56QRTa02RVdTiL12
gjVyYdnlYfJr9ohdPjrEyIZ17a6G5sUTH9jNyjEu7khl0aU1OcmBqsKffxmXkMXf
ka9u0jIBkCYnRlk6X4MTbRcmBZVs36ICxrslpHKf8eLQ3dn3p+EkDnhrxwQEHdgR
chJYKbQuNX/856WS7XBFaahMb8IgAJEz/CZZwwu4wRSnCfKVQWMpXdVDolWytiZL
nvPIFGcFo78ATjlQc/w19MCf6s9TvFHmKdlnEig5WoACXshbmuW35lK38rhI/ZOP
pPilDev2nco2S/IIRhfpn6QsLlUum/epM0vw8cZZVDu2g23e42Uxo1AklsB+h0MT
Q9ZSf8iOu3t3B1mxxLOaSVGZzQOZy5ekN1rYTCFvlcvQ/lkypXiBurMR/ySXFgpI
Bjw3kg+s1cug+ooaqs65cO/CqhTm3l/yLE5FpCWrTTHSRZQ618wnbmqG6gYeclbW
XS9fBVUWq/OS72ywAEMPTNkCT+XHvvwH/P57it3V6Ie+qoyaNmXX4BfkBrqAC8uM
kuQ/Bg2PiWfRS9Q8z3qfI6mPy0O+Wy3RpZsBL7rsRpzLun8RUSu/PLk3l1eQDbp7
g7ZEpe9bbhV6SyXKxYAApKQh3qfOh0jVLS68Mz/7cwy96mr+xz/PZnFRnExD72bb
rDe77fps5qVbujt94yVzRyGo1HqDCXLGXNqXIRHzgvOWWTKnB2Ix5W1D27egS1U8
PprphSuhzToHuS1YoYAIRIZzTWBD5nFTmaSlH3tAR4mPiKpbxBCfESdhAPfG/Rxd
yTBWo/jw9rR1lDsuoLGKE1nm/p/W2BUrvrs1ELrLjn0AtqwUFlYRQQ3O9ivcNxUb
MGVoleonRyAJJg+G6Fet5Kxlnsg8CAz/97b/tzGJ9P3vXPPyW6aDg7OlCnqXL2iR
FISupHqUK+afsnRe1xkTUA4uaMafQflNbWtQ7lImzAhONaaXYgAv1fURMXTeBjmG
1tPI0Un/clAO9oW0TZdvjANVTzX5JxaPRI5aPUYkIxljf4T1F3UYYVhzjzdDJGs0
+i5UooFURtpEpCip/EJfr7xzjZgPcJJLttkkgGabgrvj5StD/LwRH6hn4XntuGs6
1usUiNYIGAx/zaomKBMaSDHFhKi0ZtG/gdINbNeNT122ryWQRAJZG8h2s3t6zhh8
ZeWM05W6VoCt1vTIWUql8WerUughVOQBF6cxtMzBr0H2ILzKsKHctfaotTTsIDId
ahJR/PvOgPwQYUlo1HiYt1Y0rqUvJqGaS+xdpU/4f52J9lTpYZdFsxkXvTAhOrAD
qauJ4RobcOiKrXukIfhzS/WbZM1O2m7VUY+BGsY2evEglSiAvB1294wC/EXYugMX
0XPeYU/3uRCkAdFyrS3bZHVytVANsjUjwYQc+6e1pcdl39g1pZN7s/tvCCSvJceQ
q9j/dmVBv0A7u3lvG4WMa+CdY3mzaXJMIyxAyDX0I+iMFXiKgi0EFJQblTqXyq3q
bCdIgswX2pDxDKyy9LVinjKX1kLZxCZfLfpnvW+0y5ZbxMY4izwFinXU7c229xFg
w3+dqoz/Un62lzM1s9RpaLeWyEBWsljfo9mOLsUq6iMWdnuCviBMmvjnKY/6l9T0
BT9/tvYY43sq1cUQJrtEFRBhT60aWTXhNcoVNx7J82oDYiVWsph/uaSaQFvJS1XG
ut3wkTCCeJCRIA/f8YgOX3YrrRykNPflorWtT1GZAXyvmoEePNe4AKqlGgbMkeJW
oGVIiEeqBAeNZIASW/5YmXG387JFM9nGLFv1pGxJs99UGrr3Nr613RU556js7Ods
T97q8nuYoOLt2DrGiojGdokJth6hujy1Nf8BpLBjcTz/Mjl+akQLWGy2YLsa/AoO
JeJzTMi6A05L9hAFj0q1Glpz12xCSVPDUf+1+hoRqH3Z0qWYJBCwqaCBTe9rU/4z
WRSMzKasveB+OaKhk84sgkrEOkWG/bMB6rorWCgBZutCu5ATYt7TIJK9PHdSQcwj
x+RQgBgKdNjmd8LhHNFIIv4VSxJ3bkLNz4+RR08bgBQ1kajsGuw8ZEj+mFG3VThY
k72uyRw+kXebrl3GDGpXE5yVCTwIZMHSMNnS1z9ADAic7SoXxcZx5OYPZbuk288R
Z+fVM/gcynd6enK7IkZrmrurgugELNbyejafu700HA6YysKgHKezX8cg9gZ794Wy
oIRZQGvvUZX7ePMSOmsQqUR30fKvq6gn5qVbyNGUa2Klep0Ab3sWYhikUqM5vFWb
HM4oa9O0keqtuyNaYC+KwiOni2s8wwOJw7zCQG2TRz4u5+lAYiGFGYr/G1UDvryo
d9W9kG9/6IzTih59wsOt6JXrD+/ulms1GQ4OSzD5nwAxdaTp9Sgoru3wm2ASEWRB
6XsKaLK4ZBpqfm7KRqeejL11+7w/f0Sq95OotZRX19D+JpotI6JJM3lpcc7xr85/
L0I2Z4gll/SaC9vuybFCjUZ0GFvt5MpfNej2DbaHGmhXar8RNmUU01OsL378MtE9
Y8HfsTyuhr5E34VEXHYg8TnwnhR/UuGrD32vcmG/BzB8s9/qaOF5r+6RYEbnua3G
N9j0c9pDZFn/FG1+VMEQP2Ii7lEKQkeDR3VGwv9wNWsXLKJDHcz7OV/spLNG9Q4x
vq8YEI+RQIV1o1uxjxvs0VHQkIaVr9W93+Jhks88aYZIXgiUV32tALg/EX2cBonX
D/fSApeTfgstpvtzLToGxpqFfrjI9mqn3OU1Vg11N8/Cp/ekf0Y/U4cofj3DwQK4
fb065GpQmrz1IKSqemT63xGS71bksh5ACC7qMb+kPOQK6mQutG5CklHoBM45ePSl
NQK+n191OgHlJIVcbLwtz6GRNNeMnZB3p3yZchQwRSdUxjj9eEwT5jxHiJaQ/rX9
6bEyiMen1tOWI7xoNCeMBdpki6CJlRrswl6cOk8r11HlWQBsDkYOAgmWVmdK68jW
ebsHV2mY1L5tXkEToNrKWUiuUHq/6fiL1hSfubqMOQU3rUuV4NYCiVjRWoVlYigv
z5o/bnqvCMfb5fZeqruYD7mztxxnooceEBjOB4OUx8XGv+/3B84qDfWGvWx05DXm
03qsjlu7ImdNNWPIHx3Dy2Aes5SmtyG4oAa847Jep/Tb81ny+t4dv9dRvJ3zNUSl
Nt0wxy4KHF3Vv/V9RlBFjM4dJr4yS/HMcpznu9BRmiZr6VYytdTSwz7lj0gY4Pz2
3kfMhTe5ieN4RROS0DAW10JK+wTcTBJjqFHB2/vAQVko6lDmtBGdgxAJ06MPDflO
/rnsJwHISKyiO546BEcxJhqeT/6gNwr5rQh0cFwntOhwW2VYvdvhJ+VtvNDXVwpz
EhrboCc0h78bPJazZPZyjyUWZr91ck7m2OCSjk+7W7pVH02rdGR/+X0WgMBjBre6
5mYi7e2CueQjTDeieyetXDulfvT6B5ja1Vv+LoXCbYHgVboQdTC493MbOxAtN2RI
iUcS9/DmfzPeGAJkW4VXPm+ooTrb6jXZ91Zx7TvaNg15w8CbSn/Nk8TO+Jl2r7sx
vsy1dsj0yR2QVH0/ZLHkqat6OFdmK6LAX8fSrX+tSoLmCehYb7NaiJSJLcGlRybM
bbY51Y4TAOUOO/vqmQGirxMvZ0pmkD9Ete0pzZibmrFVyLkFJKf0WtQSYR8vnTz7
8FXP1TpkufFEfkeYO6dZIum/5U8m9Gze1CmRMkEC1q8+WD6oYZ+taxL1ylbNrSd2
6njhCuFZ6bEA6MwV1msyWIwVcY6MFdWPmumhwkxLFXO39o7eFb/yy0QeWMW8Eo+u
gCok9nlnjDHFCXaSCj76JE4rR0zmp8Fwy7IPg1Gy1UfldZjnuMW493OIhZPcznnt
t+/vh4iRQOfb44INmkja8LxTnza5862pt2S671FPYApKCvHCLqUt59swSu6q45fj
t/bID59wpnPdr9JQjr6MI7deHCs01lVPBeEz5kyHb4aV30iq1heOq+98M6z2FOol
UF/UeRtNELy8weuISVTRXtAQzzL7U8Hr6hrORi3vGxYQ6lMKy/RIvZY4hrCSHTla
fQAZ0OLDm54S8PUiwAwizwQ1ZQUdrb1G0w4hLv6P4wgIXlaAoT3HQqujALt+sjHH
PkMvK/L1VWq3Sww+ILNP8NQ5axQY4EN5tNmlce/dNsIb/tnXOQPGXXGtKDKjPasd
B8YGfLhu0GRZdqLqy9tjjq04baN5OcU7w77plalb1m7X/IGFWxrSA5mtSoDSJWsa
+NzudiyVZ9+EISOJfdEAainwJOYyz10r+BkL6CY9o9F6wJlZhP8ProxmWun4et6t
KFgJYlUT03caa1en5w682ba40dVSHvl21WpE4ykQHhi/Af5RU7MI/+aZsdM39Oqx
Nkis0YQNWchKa+ifmmEs3QDJQCZUbJ7DxFakNv1GtEPMKDT/HHRnJS/f9CUV2eF+
p6CXQgrDhjzz/n2u22ruGJ76jUXjMHuZDv5jm5Mpv8gLbFlKDu8rMDQCnV/eJ0cp
XlKjud4IprMlf9QUlzj/K3CGciRVBe1JK3srKhbePV2E4SC2Tw/ETDs8M0AXUDNG
brM4Eb01v3Wj2xTDH+cLkhWel7gVg618BkcEyjzr2UEwCcFopJKi97Gip+cXXavY
mKhKb3EkfKJyE304AXnGqsToy76LLU00xuh59LWmKR49vG1vcwOJPbyJHIf8epun
g4lFEFS3H56hvcgN379szUgADZMhSAePjmeTeqs7EJWsyZPqPPvaGpUvYYpiDUcH
tRNYcrcBOBMu1j4MxYVB7tKovScKyjCPIiUfHKYLaUPeJaFtJI5P+tiN16ZldnpN
rx378wYMnTdpmShnq3UFKLLPOMBl+ox1c1fmZB7tsEqcd9XLhr6JZkiNaBBTBSVN
FNz+cMfqzDUWEmew0knmMRb6DeUL4a1/3H197UCxQYuz5iS72yRvePpEhNvV7hFh
br8JwYI0Dzgdc3BrgVYn9uf0i9fUdN4Gh/EQcLcCLjCxeaqTeptkHrN/03ekzFLl
rIg896sBf/1i5NbQFk6Uu+oXoQzOjMBC4U7EAOn/YvGrMQJi6QEJ6MLLALEHt1cO
BDJBHAmTMzN+2o7M4L6gDDZFQcLQeF22aGQhOfn2F7bnR0J/MjpvNu517srv9Jhw
XxhoGdvQMC8Rba3p1cBdFeDF0lYQF0qwfRj+S2YZfHEn+YYwZwN6bboeT3WNXk6s
aCFIkvhd1eld42+P737HZeKsmSYXVTX7P7lMLymWNoOCVcxrIb6KW/hgGaqO6P9C
RD9qmafYXMyfK7vTB1rJynEDS0gyU9V36g9BEieKd3r4qWZYk6zyhsR/VEk9tu/m
BWUPX3PNABr79ok0Vb1oiubpjC0kUonQEIaMnrs9SGyIkMCw83kIVdv5h5tPBp0t
BSKD+v2G6Kt6qu0DF+J5b199vvke6MJNIdMefzVBYJWxX/bQL8JHRAjLCP525Qiv
NWyPYQm22rbjuseNXhFbmiH6nqIxq892xOshcCNGMWqm6E6UNWh772AA+bggbiKO
fVPg6ebJ6kax67DaxOZKzwy5qBHjiEgCt6us9xnPIfdRnfPPGN1Lw1TrZJu6RZrp
zzZ/Qc7qJKYIaGBmSYDYIyHMLM10jzrtlpPQCaU8/gCqfeLnMHu3vx7nFYSbLVeY
+e0eLE6JIpdseBVUEBjOkG88ZGX1ZvG+bHAtokwqawrHQvF8780c50/v+d8nHzNN
8qDF+8utnaCTLlCegfmnDbhK+tva2YDnIu68hP+H0n8KJyJ35LUHwRT0GYPIOdFy
GKetgzRUQLmmE7joDtQLzT7l5WzQ/0MJjsl+KtDHttMDTXVsb9NyyPLhoSDRIQnC
bq9EC0bzWTge+gnK4iZC3czOo+eQX6QnDbvMBPqIpZ4/Ur63W0+UQh1zLPCoy8cm
M7iyoW0e2iVhGXVAgcNOhxaLftAyVLonaWG5B++G2sCkBlTdvEkmkqcOQxkovz/b
9llS96J426Xrh66dywn6dj/UcwjQogY1tuDJKOdATvpHniET2roEqEBjLJAxMWDM
sviWACyH9ds/qyviq4alHpWwLizOtUNCKxTGqn2ZMnb0h6Rr5907PqLzZQ+Z88Qw
bFOIjExLaU+Z0+vKkRZKJKipDIaC5rI5WT1s9wNL/YrwFmk8FiXQaXnCSz3x8ITE
Pn1jqUeCD8I5NQWgeJNN6/uu9n0R1r5Dsidlx4EYzWIQKKgSevWgZjUHUVP3FVxG
EKIsiQG/MU20jevbNOgimtExCkod/UBLmjqPDIBanfBVBRzrVPfYwYuoJ0u5uETL
kjWiCgEZglXCIOwY6zsOWMCJtojlKDeBz4U5j3MwSubkCxz170JVkh9PTS/T7fRF
xA9NEVeGDoNSOKlvhOH9cWw1BpDz0mkATxlO1p93ssb8rV10M3ANjU5i6lH92hfd
zRQbdJiHlYQ3X1TbcZDi5ypLbxY3/zKa2yfjZeDOX5d1lUVU8KQ1pCtKklsB6S8l
HcAhWaP4/IvXY+2heC6Bc3QcsAv8P8TlPZIGikz7TEHg1XZ/vqEytP/GWGRcunyz
VanAGzIsEoCh+6BAXb8wpNqRVHGb51fg9J3YF/dTvTYLMtUKDUxy9vPzwVyqJyuB
35iMdV+nlQpSBzESXP3LwqBSxb1+4S4hIvYe2T/9MAULI1lAvzYcbdW5vr+01Vy4
pYBEpbG4BcDhI36Q54AkWGBeesI7kp54l4Mmzc9T+TVz71I6/Lq+4eMVyt689XVh
j19/AGwstib0mn0TCun4essjIsy+xhCEJy5uMOBVF+D+Wb/YtxbQE0S7rQzgM2kn
PE7NIBM9T3POSm11PjHvDNCvEPTJ6ZK7hc4wx88DyzxUC/QtAQD8zN75+o706J6V
cmpcUyAYpSVhsDtMDrvu4SLsXPxfUYjUa+FaMuduny2coJGSNjB+UrfXu2A2/rQv
U6bppOSowkHaqNjm1Nv+Cgaz+2urHX4BtSRa5Wkp4Vr/C8zYlG3FvMKo6UZ53jLC
ngQPBm9za258tROAhUsmo3xHK7nrxunt2/6udhor628YRErFt8Fv4+HOVbBid7pD
YcD8GKxFIlX1LcNozrAGVDRksybSzD1kAYuFtwizeBhEkqO7KyKMfyX9sFEMTUVt
umW2XlwzGlxDf0wKiD9ACtfgy6eF47faL2+pvUVhAIHHBS5nKkaCHWoeMgf91Hr3
JPET/OZ5Q3IRxT7fUR8NwbyPB4CWAJDdGeyQBzL7xOGIjj0m8Mxa4zB3DAOApD4R
YmFPQQGxetxmDKLHnbvfGDSkXNaKTZ9zAu1yznSR1ukq1syUdoXOt18gF6XjyiH0
Ey7yCuoT4TbTh/nLd8URRj898/7qMaa6gpCzzkpOmTChDzeNS1N0/WO6pb6wM89i
xfBOWTIWAUnC5NlD5IaT5VKzVdHVlEkiSVec02UdnWcO6TvkdqUhppSeUp1go1YL
5ot/XFPN3dIDRsVmU+oSqtm/XoIeNgZYjsZe4bhTP6/w6yR1YWsVm6pt/NeHZlzw
G2smatoTs08DCljsKF9jLCoZsw0YxzG6adTK3SGrRPFA1o0cyXDW7RkMl9t3mp+e
zn3j/VYOvsZptAVgy3eAI8+ZngvRRJ+pqdV3pz28ZhEqTzhUuNOCt8+g/6fZPWJO
V0kDwstCWWuOVjBRe9QA2PeBI9/raWkRtRyQP5V/fflBdwXUV9UIOwAwyEwCUlFP
jH+DLEofIs5gV+knDv8YQVZSZ18oB1PWgv0h+OFI/0KtYdd0N44qBjvtf3rNheau
3s0MeDvWkh+anVQbmocSaBLclOrr8B7jzuiXce6gb5mnQbiG+Z9mIppkCqidRIoD
L45JyznjlPHYTyzFw35ivWbm8lTLe+/vCKKbCRcT8l3pTEVQ8sfHjbZMeNcNz0fL
HFbJE2IkTl3s0XGLXzmV4YjAcVcxycmJirNQctTNx56VPcg9g2zCkQCQNVWOSd1T
nJuXzXthlrVQq8Xr9AXHtO49YdQBm9FUcFhOJ6Z691B0u+UWfaL5AzCAgYWfHg27
4m7F/fxQ+8DJhj23vwuv9OeFM1F+qzOBb2HgrEH66lSC0Qd1D1Yi63yGdakaggeC
+pGA6NUsYsHUtq4VHByYes6158Qxzc0z1mUlfjnaRVUOjOxRTJLL5JT9Bv+kSK5i
o+JIu52Bvl4ohO7ye8jD0aDyi8Bf1TQjwhfjwyJFbxj4lLV5PUeJQIlYJTRUs4S1
90qltkAd6lJQycEDu1gHPI8q4NvpEm7YAosvlJCD2XcG0LPW2KKRKNmKsOXXAfVv
WP1lb7QpQj6hokTvXGiH5vtzU0CCV1l/gI2sTtmb1jqhsxpAyonYd4QFxXYqG9OW
mQSEClvY1iNC//u2t8v0QMHEM3821L1ftFsBETbJZCJqxTN0d7ygjxosCoLY411y
IhAKvWV7d6BnqmRv2cb8FBdC9iyXMuhX9dSAA6QWl56ZodvqcM/87FanoXlfKWTg
Y7tzbEQY/PJue8jTmjQElKylNtraEQPkur6QzdpemYri912isIqgNtfuKpF3SQ/l
xk0NxmR1N39BJUFWfroPEfC+pJX8z1A+29JXyaF+hWz77rwLlbHPk3r6ef15VAov
Wbykw7LkhqredqmJWgmQF03PhrAhM0XxaTL1Y+NScSSoC/ePAlTgfhbYDVo5KUCO
0ZVcm4ofYfKbZ/iZgACqzbi0HnHam2EsJVl9tsb5zTg2LU41zp79NlTiLZ6bdiMn
ML5CTI0JgloDUvLR79v9AgmPqoFqIQtK2JRF+MFsV0MhW0o6qp+sOUtKXz6LZ4an
QPzfJSRPROxKo+jpst0EvGsgZRo3ZEPXNjxJtvi/icbHcfOYeXei15e14Mx0b5/O
OiLXsO/QYOW76TGAoV/qLpNcaKMzVT3BgR8Fg3gx5ZYaPImTU+F8iuSmh7OXSZc+
7UpX0syACx8mph33264/x+C2m8v9CJGhPfUaU7hyaC6pW06szSEvtGvf/3X/bjT4
AGTEBTWHVcDw5uXXNE71ObXqO2uubWOHUd6Uj1yhvkdKamHNsWscPO2bqrua7ENG
72iSWeoQsUAFOIYyNw5YpEy/N/A9wlqE3YcV++MeKM+fFrxMDd9Wcaphe7DTmJ7R
lrgg6g6uI8ObKPdkSmBJlAUa5oFKfdKx+bGYt9J+vbB1FFuBekdV1glSV8NstghB
EXhr2jTKKS6nuJSa5EQEUVCbqX3rKpq3RD8SExHQDTmcFaduZuPNjULIKqASUHUv
LPim3nP9y9F9lyyS1ScCvReSiUGZTr26V6Se1U78vdbEQ9w1W/52mQ3AJKpWNfDf
/kZcOcYguklsADo05JqTQLgeag4ii/Yz2d0D/FA2P8yILYsolr7h6FglSHNU0q/C
lvy9bfWz2nGG3sPygFciY5PSpe7mK5sBDIO2gNP8/MW2Uy5uQbqT4csP9LZ2kUAp
NrfIomMQWNTP9Eo2C0slQO8tpz8nU7w58H7c/NU8tvCXL6SFeTYfDTw5ZJgUOISI
euNSCrW8fPXNWb4Hc7L9+W9G6GHPQOPM+rv+U25ZQ54oInWN1hWlQ071BDPB/HOI
h2uifwDO7Q66LqOyRx2oZte1TqskHw82PWPm+UWK9I0we53r0HTZl2pyqFMZ13ye
LTB7sQ4ILCjbm6z+iheJ3TZ4ILvHa63WG4zCI3WVtpB9WdW2ScULd10/OKBn9456
t7EU8uZPuMNlbup29RbFwKQW1lLvLiEKbao6kiz0tzdRYQreGpuI6/1VwDEI5wXU
PAnWD1RAV3o2RGa+Xm+tS9wD/aYh6C/YC1thH0+07ysyHl1TPDZ09QNTDczTCjxm
3yl0MODxcZSzfCUIxYubNHxs0XSquoAT8JLWudqLvpP/nBI8JIVBwx27YTCmVNIC
xs/JpF756BlBlEbBxU42u0hszDJYqw32bUoaNh8C/QJ2oF2LrVmerxvXXkzM9TJI
t5/kQfXvG1RQLVf0wpaTyTYtkJvlexDn8oReN4P9X8C6w7dDvz5dLPFv945YxvoW
cSBrQ2fOapuwriY6LciB9qPB3+GqIi4eSD+BGLMy1sicZH1pvO4HusE+JItLtu4K
L45TvGRI8E1aK7Yt9W9Ke+prYpkoOaToJLxTSAxhNxpYpGlm+KFG1vA1YvKo4bHA
EOR/kPSePfWEi8P0nRDLzuYq9pn5IcNIFjm/XIE6Mmzism0MAL2d9QpQBxCKSGMX
+QwIFLrQjz3MfKFZ3JLEHaywKimQ/vcnMq+RGBH0amFVoYT7Igig/T753WCC3GtO
IzpJe4m3lAi56fufpAcbonl9atbW9Cn0y5Y0jZMQ/7bMfyWi1qbD8Rt2OcqzLM7B
VLCwUm2aQQURjcEwUPCdpwmE4hb0RizlRC/xDYnoUGWtuXCG7vqNVvlOts8PY4k6
ginO25XWtRmxkfKtOZQCgTec5xaRFgoqX8kVKNO6xIlLEHZL04ADYUffJEzkrI0D
KNFkIIEJFt8/hlws7i4gDf/IYy64OLfJXW7aEJL4n+Ky9ELXBYMhvuGAgwabD8eS
NFl4+E7mkJcqe5/JzGdxL1kQl78qGhy1CVIFrs3YUeqs+1MNDyaktiAGPi+9vnqG
C7TCK/AD1BLOmxwpGLIocv8QI6+/9Pbr81uIQ5n8x36NW6eMwJSvUnxSUp4dB8AY
KNbefSrUuK3nOMlYUr93/wlajswTUbwT4g8o7G3O9MPJPy6R37xvYCjWP6CeTwc8
f3DCR9MA3mantUJbjLFuVhpY5G5j9K4FRCv3O3Pk9k7cwPsxVpNkGcPXmSRBQwGS
CAunw6wD2iq98xP4kTsgVE043M5L3vygW8/JWVq22JuETXXoZ2CRICLVi9IJbO//
5jJmD2zy+5CZ89kQEslb7aN48wo7ApuYDBz45F4yQvOycQfuWfJCQ1oAxcJnTHNH
gIpgvnThE1kt9Am9NQnV/KF45Sg61Yr9btRfHcDPSG2GGT1sqYF1eIlrrou8gdCe
2nDccA2OJ8inGWsrBGluKnQszLhn1mxb7P4glMSsPEizePUn3PyzH4jGamILcx0X
5NqO55EHlM0cK10EkMuZn2anSsgeAIS5pzI5HXJ5aOMtFOluJxecNcawTTe4w7WG
Z/M6YWvdawICwk/MK9jbad3LkKbkGoOKjYQhGP9FvXVDHZ1pwvnwHIMO+Mt5ij8Z
W9QoRO5bQYbdmYtYO00uH7X9br89NAA3CFSEfRJSqCJc2a6+m/tj3updJbN7EpUh
XhWNzyqQzX4cMFpcPFhBpEzVX2qKxPDouUZX6J1zkDiSCfVqH0h8N/VHzIf+zJ+F
ODDyHETpc4QDPeARN02c79i4xDsbqmh4Zws5dcY5Z0PXMyNgrUt6Yay/DGV3D3qp
eHfr0NFskK312sT3B2uqtyASWSIqDvuuvSID3OjloR2zlguqAuVHfSuohDwyFLmu
7P28Z9LU+wTEWPWnbcm+2nkD1Vkwa6qcaIEtzHWOCGdLPX2D2iIj0BdCZWk4CH4Z
Zbg7A/SKTqSK/Pa8AzgeFEKnpZt/vdyTjIhlTxUdQT5ktOKOFBT5h1uwmZSWHzAU
9ZNHDe+z66LBucThlgtpYs6YkkUQ0FF5U2KGuI7mZJJQ7kUfW283uRZIxNi1Hv98
zyo0STOydfX/gBTc0+dardGYpSte/9/OA1Y8ONCkTxx/Z0QvyPb+fAcvHBF8hStz
fam8qWHOR1OUialc7eb5hD1TsWnk90fjYBQ2sKeMYI/ILkRWuglkffOr9ZkXa47t
MP9jgkppAQuXmRIjD7z7NmZbIS2Ff5nObB20fe5gaJcnIWEb6ta9H8JoUaQBPF6w
ChdtU7XDdazjBUd4r/oCzS2+/QO3ZYMrBX61SCGZk5afSc4KwDt8KKwJbT1fWan+
O4OC+NGhq0rjo9HtDaOThbQFOr5lFmh4jlhqf0L8ZZBnku6CPa1XFRPU7Ic4Mkxm
wTrj52zxXvU2scON3koASQzSMb9JXT+wkIGSMDm3bKjqhzqN4OcKoYqZTJITDCS4
B8vrpLRK747JVDdXC6i9p4s/JZv4dJv5CGS+590sLL43G3q+WdT0UiMaqjLzx3ng
EJoIH3m5hb/ZWVXtlPmd41cvbDJch/Jra3DRyHzpapolntSS+3mXIQ4eU23K34pw
vZW6GFQhqT5vv4UDRF0a0Y58OFRabbD2SRWKEdSmozrXsKIpzeRr57/b3EyVpFj/
7IP7BJBSeYT1+l/ZIxD3MpiWd4UXnjySWqztDH3bMMUJFtZnA+4dpqzxlyKcJDOS
G28s93pRsLaU6vPav2D+usFAK/5ZxiAB8Lfj9/XhhponEPRqkqorkaKY+2tUjyLX
r03brSvup8Jp8tuE7hof6OqdMleOYx5YPQezZv2VQrmD0QW5u0/DZdMC8EveaWus
3Crg2pcPWVpRMvRXXz/e3r96YDIGyoCF+qpH3BrHA+ltKZKgkrxahwVQrKLRf7Ts
IP8Bk2xfawsQbgpTQASL4AgtNaVZvIM3TbOW+lVXhr4As63iAdKGSZxlwWpCm8xh
Lrc3IyCQvzea/aKcluB7bnDnJ92F/uZ1HodsdtAeK+ZlVm2EO2udZs8p5bWhL4/V
b8h/jDQXjP3F/AmY9sp5jGQUBnJBCdkbhSjGqGaz3JxdUxTg7L91Kr/0lUlbYycP
VCxFmBXZeldFfk1AV4L/5YQ8pvugnLxECWBkcw5Lnwes+5vJjxULBckTjqmmwDGL
SvFYLCesUgMY8sgM00Ydndi5ljuF5RfJxoFvk4lrv/xcfrA8kNQkcIT1SfzExdSK
CQdQseUugEaAMxRspDMTp/2Ef8B++KlNBT0dgDTk2kH0E6XwiAA9kSLryS83ATn1
mCLlwVYgUo8jARXmV/BKdHqSpP6fqcteINBX1+2DsXJd+FlwxyzxbUFhrmSNtufQ
JtUUC3byTIs6SZV5BL2MSzFzrzMj+FrzlWxweqyR9IAeMk1vx45Y9iQrZPsq4FXs
3W+MAxBye+AH9+mzsOur5JyJyNjzEWOpyVnKF1m7oZMsp2gHuAQ83t4uO/l3Lvnb
uJ7lgvYd8vVvFD56xBycCwt4bRNzze+oHKabOXKJSMZ9lLoKORhiB2s84bYmS1cb
cj62xLHZ8nywd/jei3zwjm8oNb9mFMVewqtPubPkinso80NmJGiwcOWH3FyQpV7d
GkG6uSEp2JS2TKOok18Ny+Ze+PmGJw38TkmZVWuGigPJsn6i2VMieZj31jsn1k5A
3qXcykvjKvadr94Tv5NBtWLCJljCvuCQGwEj142Nc0HwLZ7KJ5oDjS8P3zRBuqdV
oKNAikSbtVk+N5rfAVpIqPXIf9uCs5qSX0goMhUcQoKSSAUjxNCp5Q9NWai7zEUS
gsfuj9aJ/QydjGBMzl7YetgK3gXz76M3b7YYZCtav40rtsm4SVbqI5SsuaxrCIV4
3+YgIdWjJVs0jOmPDAWWHmiqh5rASy7nx5H078pv65PwvwiSY8sgJybTkK6CPPLP
4O79/LqAWdFlMOBxIN8dNaL7tqy9Eqn2cQpcvI/tWT0XlBSvJONDczXnDv1AXSin
PO/HnS06DF0GrUbUZRjP+rwSF7DF+f0YXmJ1pILtLdAfKujT4WfAyxx/CVOAUqpT
J80hXL5KPgjfh+r40ojahtlgdSB1w9J52TafUHWuRdr2UWw9q93b+y4onNXFE5Eg
qmJCC+aiP5e9IRBtsng9vLp90GmdgBhyhpWres+21uXN8kkk7//6Zfttlu64GWWA
JET/Tc10JX1aCV6ebUuEkMYtC+FOHD2kR52A9Z2Q4bmJ53Jk+0lMZkjGYByqfBvZ
f4MFRJQqiCdZTLrpq26gHKC9Zh2Wq8mt7P+trD/pXVcwp+iLzKSJ6H5ofqyBN5ta
FfIrKbJUDAKdG+c+KttMGbtUvRLX65NgcOyQSaxC6/KEs5lutMtbj0VwwLx5CpvB
o9C6HP+5dKc+T1DlT7ckGCd8uJ5ljsfJXpK3QuNtVF89rk2vi2KHtIPI4IxLWFfG
wWjFRu+Uk8oU7xY2qM3FJvkOgVIrp94Gr7T9kXdHK9O/AUj96psSzTQ8iej10LBa
++SEIjUDOV5y0I6MnjjK+lqlSm0anscwi63L70PzMI1DNRruPoc+t4V5V3xjPyjk
BG6RKJv8wx8PZI+BQv9NcAGWS3uZvNlkRNkf2YKBg6BQUFhhmWo7eo0ecnGwhrmH
EoJhgl1FEIpUzqdPLQC/XnE9DlFlTv86oC9KDcWTyFcNeo7WB2U1jrzUewHK7b2A
Gd5X2nYi6L4zDxlqKppGm3gh1lht+CjD/p6oNybifUEw3ubUZPjgWVBejeMP+HzC
w5GRiYR/XSFHWzeCB/zFdoKVdl37vJg5C1dx/eP2KXuuWsfqI8hLfG6mejcj36I9
+WhxzBiK29fWAflYADHzW5Keeg0Dfcsa1KnMcewnrEN9KUvq/9xhsF3RCIumb2fQ
j0pIGxDrH3Hse0EtVqaaH53osSxOHZjdzDp6cVebBJfKX3Bdul0EGB/RVzo6VAZ7
mgT1cNfukl02sokifdsmksDpo9kS/WGCijRxdmUAfs2GMnY8/pifDvtbk+4HriCR
GNjJRmVr3L7UN+t/nUI5aEX1Jl/7HqZJFcH1CjtGwLS68IS7kZ8znW9fPOjmXJGK
jOfpvIcjcL0kH7Kur+nWkS3W4JRF2p+mSv/8qiONjAXOoBnM6mWbDD1cUOHNvqVy
S+oOhoVEj3baDB2VyuaLn+SCcjY0a9iduqSS4pm3KDyP36N6CU31VXU4F79/nuRl
90XwynqLq0lywbzWlNngWpxPz/eG0b+7W6A4BnBV9RXuAGfmMEsa201OPiP2jBh6
x3U5sVreqH57bh0UwSmwHf2A7KSKwr5Y2GcZ6Hxfvhn49vMARMl5yx8GVeAY4wEr
XGP3OE3s4qUwruB5fkR48f5AeC0UpvLig3Cvn7jPfaK7cHShaROpOLjy7C/Huxcf
3Bysr3RwARwM0evMw9GuWxjD3nFU4kQvI/ZBUR8JWn7GeyOphYpjdUBbMlNA1kt8
8XJ7lUCmfNie4H6dprX2ykVDiM5s96LpLf3ftjVPKwRy059gAv7RwruHHhmrgouC
V6U5MGNMoIY01UYLCUw83cL+bACMQ72XNbbr1++cqsVY6gDfgTBDt8TJ3251hTE0
fDkY1sUXMaOFzwe5AYcXjf+Yb56MSXPXsswmoB56giS5iQgUCSXFXxfpJFm9PYe5
2YRNHyjP5GfA+jd9JXUepDeSnHyoDmS9ZxFNcqADzs/1Npgore5X7Ts7z3jPxhZW
Sd9FfHh6at5Qo7r9A9RPG76x6IPvFg0jCLlUO4Pcqinv7H9yHVZ9AxEMIL3xuw/Z
8bD6LYa7TIHY6QV94JI+zi3xWips+qEyaeC7zyKiK89cOsx5e6t4krtyowMZBF8f
pJ4xVO75RpS1BFPMEAbm6/IpAPyNmXxZnPkOJ18WRkIPyqPaPI/HRQEaKLAZJw6h
wt7kCDmnBcu9uaIB1dNmKUDvCxRW5EAqr26cr6DsYpf4GrhmuVzf5CH0EBEJ/ZDa
RoWIZO3j6IHAc1moF7rPZkaig430hX1xBOWEDTSW3ao3yVJ/xzpIO2GhXZOc74jb
Hz7IPsDsChbIz8NG5mg9Ch0e7qHo1v36JogqwPhdbxqYcYx568OYdmI5SjtpEzkC
88hNteuJ8ZMqTG67RrLo12OOWjdssoGgsIG72CjneuZ3J5utdEeVlmYYiIvId/om
XrZKVkaw1ZZ4iDUbLV0BeLGgbJkEu/ZHnmJSFoggjT3ZHw+DYemkjo8BkUMMi8UC
foKH8JIekb7rPi5awqOZenxRjFL+4WxjFwHcNAcU9zn/mRK4UHt7IZyu5tN2D11m
zDeQqttY7wY17F1D4+Epua26adKfddTOLniruPgb3sngUVk6qvWQ1KX6JXSia+OP
x1sErpyQ+kttGCqSu4D2rgdhRItDnMWvWt9BJquhZqHURrSfNQ1pBNXJsOVspKTh
Wubyonw6voFQJdm5iS5aIzJVOim5ubdFPICWFRHS4UdUZorONN+Ixd1jY/mhJ8KR
aJGNfNC9BxL2sqB/TX/+TyUVjbEKPSg5cCTMYYM+82W0NZJKZ6LyqxmkbjK17bxB
uoL32vZSmbzbFnuU5KA2YYH5eTV+79aNq2/SCxuk8EpwsIWpby/s51aHkpoe8BZZ
v5hitGQBvt46CaJ4ZY5efhPN6mNC6UrS/8G7FTMyrqd5B0GlYx2Jn+imo2mevSns
gdn4GOuIdZxLkDYh1WS0wFfNrPszn9XR+RFXY90lvfULImC5iVNZBSWLbruOL+kT
SDYouZ7FA8CAs3U3RDkn6FZ2wNYa6noI0Y/g7iT+2y9eAvGQTBCfnPrEDnG3HczD
Cd5oTL/Hi0YfSUYPLPAONMPPmzGtcUctiHKrC1v9ONofZRzxBC4csqUyrdbEfss3
GJmwGUBDuXhCy8/VTbYz5ndvwmZPpAdiIQuaUGEEPu+c0acOuC9LCK22hX3aplGN
gERtOAqmW68Teefit4LMQ4BDBIwJiKBfn45Jdp1tFMgl+MyMiBJ+RXEc9RCiMPrP
t283g4Gt1IMV6dCNxlV/9z+El409hjH401nJk/mV0bSPonJxdQQE8wIQJTxVYUad
KZxEzqqVjsHeIEAiKDA/KgcPwl8lwBd54nePPZnUfCwny3M9WD9RP/qu60o5u2r8
3VePADWPT2nOE+EyUcu19Ac0iBotMqEIsO0Zui1GMK9c484ug+jEL7B2XU2VdSYr
YZBAnU6n3jyqd+LSAXVX9tswyqHgz5F345sKX6hdXvZT7EAHn1ZwLs9/UtDmXwGc
F134T7GIqfifpzP7VlKFAYloOIwqzVuRHyT3nVKv4mdHmVlW6ToHBCPuNlymWCo2
MIwH+gRw7yfelWQB+88camPgXYcjpBQPCaEeCyrNzoK5YmtqnRHYbQKlWXuLHanT
Cdwvgts9tYBhx2GiiA1ErB590Vx+DIaIMDAGdEDDiVCZQhNu2hDT6b0hvwRG+7dW
nJx4A5ew8oJmPIk0xKYv7Zhxz4z5wsChzRiLJX7H4wO5MrqF8HFnpBoxuZfuY3kD
LV4lfE9sRNOwJvBIur36F5VMlA7Wb9/j+//0Ub3nzL9W3xfdu8PkiNBFyCDrlud7
+LoKfWizt8tB2R0qBvYjVX/PQi8a9pYgpY9o4ZG11I/gnTusZIFpXRrBlytb2BCN
O1RDWd04w5qmW5JtWqilD15oA0hgb3MPIA5shSTKQ6hRZ7qGDj8XOncVeGcXBsYl
KogFZ5nwJuDbaeA3KqfShcWIbxEg/ShlwdXZX4tZTMiBolawt+wUFXNyq6eVkDSK
o0RRuoktX71QVfdmCnmJZC3BF4R6YcmgT2zVu4C3fI/5o9QrEGSy2UpZ38JVhAnC
SxCNvof5Pi5A3W51Art0jC+HaCgkzA0ZYsdxfarEH3z6dlrrMkTiwQ2WtSL7+Rpz
VOFLOAYuMmPzcmrjEf2kKigIslPmshQFAyBd14Ev+KdfpxUnurQ0rzr7SZ+DunWY
WrOYaqqhdL0K476dYZgiu+1MbY/J8kXIkuLq3UIMeB3qPBn2h7iu6QZxhqdR7SXD
6tn+M/48yd2bpOT9rfJBPF6HxJ3V5kVCk1zLg1wMIOLZnvcA26Yq9JYiZtYKz5Qm
KlaWoY2yU+yJ2h+taUXMm8IGOMSti0zkZoajAN2jknCimpTRlm8NRBY3dgbxCndJ
jyKxiqa3xASqjVFcZGx7f3sopFSZJ42faLjNGLUrJEbO5OxjmZwa/mqsEjqygATk
rUUGd7+FOTZ7eRvGSDM+FbsfPyuIYNUwlQpRgMmYsnzDjjrwam+UBhDoRg2VZBjZ
Swanuz2H5+W3r1mL+jzP5e8xtC/AgPyNv721jkqhIakjAOX0DF5iUj9TjhSrfTPm
Gs9FzCyk1X5AJrhCT0ZVELEoI+C9Iy6JMIwZ0tiX9HPjea4YIpqHGBpcwQbH/Cog
3YR9SrR+8vc8CuBFrzHfX0MfZpb9QXUhJmw+knzXib1Rb7PVhmOhvBy4n/C5PBz5
HEa5u5kLeHQHAa2YVVdVnZ2Cv/8Iyw+N4/9hJMVhxr3mJ2rslPY0xs4aUlxqbWn0
QTFy7gZvbwRpaTu0QeZ5WtHL5MFHUnUiCyQKBEZxkcFF1IEUSyr/4KtTZ6vBXdBB
JMbeQktrXiIBdgJE3MQJQi6NcOPj+By+kaNUpafnbhFfuFKrxC1+9jFPdrXtQ+6f
L+9MeO5Aya5xqXohMDkJxYvs8s3/FEsXWndlXc0kAWhxvjPKr9tbQXkZzeuORASd
v2MtQTfQUskFvsnS2RDlwo7Y5kE3T9gJ7HAK6YxEfrksn8SagyIwra4fPHtVgVd/
pifMQ+drQ8WtQlFipqYtlJ0GA9QxQEw/4TPeTLV4WhObC7QqHplddtaMe+JztAhQ
jCb3UtEcFD2sRf9p4cPqXGWWSrEMlfkFy4+USMk8PxqVuNBlWwt7Hw1HUhMkPgdw
vJTREzv3X1rdyC8jKdKbARl9De140cKV6Pm93+45HMoDV1+XNBAI06odC6BKgbGx
ttGkMX6GJq1IcjfUzIil4cOEGTv1sKCEobG4fqA0ZBMMV5CJXItyasgeNvD2q2kI
NddUn5nkNtpTyZ9N9vqglBW9QLeOQ+CRAolQZTGSNFoyEbAMPfYz6yj1QARXCMCq
4Ftuu2L/vLOrHlwPKWon7Nk5YTFF/8Mcf1ILNV4e4QzMt4Pw1SDZNnfgSITisV4+
NDln0mBLHxrqhAA1W2JgGKt3oir5ZuVbOUlbJdLvMCmRwCwc4mGX8IqmtcJTnVEb
MdF/EUxJc66ynfxPGpTYYga8YvZ/wd7vXzy6iHEgYpHE9DW6HcUkYMSaHIsC6IAy
Q0Rb5hXvn5wN1VD9MlPBkuQhNsffHlPFdfLKAomkchD9Fj8V5L82y3RkrAkyitWb
EY56Rr++KkCG9Ki0e9mSXyOv0FXl9yMPjdbvQe0mB3zmjxXc34cjz5JJ/ZOYCQQR
LzxEK6qq0olMlqtckUarzzNq6lUiXyLjDZnBuypxF2kubJoMaVWU8d2Pbl9H9BUK
jx1kqw9OI2Okx02IhlrgfFib4snwziMSaiCP0/ROROnazZnhkXJOo1tXrFjG3ghI
o43BouGEyiksG4ZmVEc+MuU4NgtIDHl4WK/xfJVLFfUjjlTqULT1RgfMuLEjaw58
iwcOiGCavHZw45I4QByB3mESOjHXl3PgVNNjMVsi0L8E+TRL9gIdvafpDrJOnY7h
ZOdnMM8xjDwROUsXZ3Pj5hEgWD9HvLXcdneyub17RRH7vVJ5Jg3dgFh8c6mNzbp8
qY0wTtbJPsiKFhQATPQo7gSOlRb8BwjiUIiIKG9p/dyleyl3JlqExuaVuXGyrI50
N07d6FB6B9t0ACAdr3egYlrmVd4XIc4X1I1brPjLidQkema93CBvOUmo353n0KQb
x9kv/lDAtNcP5K01sSHyLa2s3FX6cGXzaggPkr0z19v1VC2wrKiCFJk5/vzJ4KWe
r1cQbSXTVIPc09Y7dN4A0/l/zeaknUWf4+5aRxrUAuf04j4PPakbmXD57SlZK+jJ
C7H6DkB3F3ry2tWKfAunx2FLfKOnheutZwoTChXL844q1mu1VDC8I/puilFYyW/9
TVX2IoELFHbKDWQtbwhZ5gQUGpTZ40K/zrc9k8ahBX/lY9dF/YUxDOUg4nNlP4Wz
0d6uA6pWNPhVAnlSDr9UNCTKugw7EW/JTUIV2fBhzYTqhHzYbRUOGFhIje2RCC3u
GegVD7ITdi7D6/UCRqA1PpR+uZY+iFpd3ZJuCdObR+139tGtOXRhnhESG8z4OXkE
bXW0Fur5PYnaBCSbPNPldmeQLJexfZA6kmqxQgfpM6ixXiO+nwVfaMpwnZU0Ex7K
NIF806WWCXe6acnTpCzFZRLmjp0I6i8DNUrW3peIn77e6lEhZpaj1ZGXYCbSpxAZ
27MqVIa0dViroDqc/QOhdoT3Aqf+TVLQPFfXk8XWGoFNC2VuD774b1VXZVFdvVc9
uQNeaSt3uruxf2QlE3TP2pHywbguLY4+YHkZqMqLfXmMRvoX8Ay+DSFV92AhoG3Y
QdDYCjQzan7ghrro15yKApQFCgOeLqk4M71nfnlb07U5i3Zj06IQUq79RTvZfgUA
ES6UGTL0MNZudDIPkoOZ9b3n/3L0Y7pJyAw7OtJFfD1YnGdYEBnZvXUsF0oDkG3t
+ODU5QIQmXZTcHehZUkGYJCVgbCkv4oSvkeGErg9HImwXBdl73ET0lbpur5J2HBV
3/CbSHXrHHRKJvbv5DFZX+o+x/e24zigjRcG/tky9nzs4zdF/OBwCfUGK2dnnCWY
iiQjMbwY5G5qd5/KjecJN4B0PFQ8z/zbK6fW/Fg5AAxRL6kfuiuE/2cSCZaqPjr8
6bRt7lwB3IOpd6bOtZjFH3UE8S2PB//HkE9TBhpIcnZNAYpzOvG5F6gxWVjuw440
aAV24fSRk0dt8n8e40r/NexArZU0vR+Balnh+2XD+uhRCIq/EZMd0ctt3qvwr4sa
6HH1YVu8j7bTrg4+mNI8ZP8k0DfF1hqHHOfDsX+Qb2//UOmj5fKVlCpsUicScA8s
N3uAIaTxmAlVARe0Uh8WLCA6qBfz6ezJAO1y0nrBIjUH/H7QawV3yHiN9O4wGsfg
p5BZDWk36SO6qWcUg+n62PcIOa/RDa8W4mf+hhZ3aitrSWSpSxTiVlc4F6frMrYf
5mO7JyPrt8XMEdTH6wioRaz/jUPmdRcAdW60lW+8Zrx/mTtaItTwX61Z2MKRE7b7
02HSvVDfKbFvrNw+n7ouQMIMdwEpxKrzNQNIXM/24TLiZqEXcZUgE/6TW9JBdXky
9LvPzOQORtF6fZSRT15oAir2nxvl5/ESO1NPhACU8TqfFRTZ1pNOJ1crfpKk2860
kz0vYom2HaRdHN7hbxZN2ndfEm2Bj1UOTtvrsNohkNG/9Iiixj+Wgg9tPnoxbwqr
UBel23kHM3ERdB4GlSV8yHMdhG15g15aRBbojjgOrAvfE85CHf6AADbLrkgBJCFw
atdVNT9MShLIgVgikjCsAK1vFlygbfDCJxw8/8mZ9LNwNIm1fURDP2Qzd2r8cOcm
IibuPn11Va4rdxnHXuB5GzFjUOa6Wbn1l6gnhQnhKLdVnAFws1DpbO9obACltjxJ
vTrjvqAPJ++8wyENXUV6zAHv10qLHave6hkRpTctt/ZxIFWBHm9y5fN59kYOlWNG
07izM5R72qsljfkudAFPPuEjfEkwdI7uGZY6GAr+gX33ee7fN30f+GI7JEGsq9MZ
qRFa8TcwCPxFUp+3tE5T8Eiwlk6n7aVzrlIoiEC+z7+ez16zUoNwcoWt8Y3jwTqB
LL/R2U4DRGL6NlJuFKsF7lvqW0H5N5eHO7MH6ixYFH50KpFaVsjfYS/sjQmL+J+b
bc5Zd6oZc+hwlRVR+zyWSAx9au1gx+ISaCu2YQtII1ls1aNTD8sHhDhg47C1OgdH
QPzztQvFlQjrh4TmXwQwlPGrs5ZxAxhchQlk/S7T1CvRUOMdNHZzSJkB50XFB21U
bk8MUpq0HqUpqvubVYiEBFskZCVjEOipEJ11TclrhxK3ujUQtWD7TDeKNHrR8Trs
vOFsxCsZJQrGHihHhH7pRo3TpBTzS60W9xkZ/zsDZq/o8oPmPt9d5KGlXGpyy0Sw
I6QJ1KDy5jyNApdv3Mz2G8yiwQmX5KLznva+OSoX9plU3w6cQqvOnf+EZipLvRYY
01mLxY/H+3x3B4oXe0DDDtHBJxCLq6DqHGPdqVIhDJ1ziFh84lrPC1ZoGjvnedcF
XVB157TkGDm/6s9DaSztFFPAjcIRNlLfN+stn5Y5dvkEo+nLSmOtg+IOH1lRANlk
n2/hSC5kPahX66tRmp8UWWMj35boqlDICoKbMbj471bH9CqLs73fOfGb4OnUfTOT
K6jTMhHYHVuadgVK75GlCc0nQSfGC+WHWUVkjbLa4gXdK/gEbW4ZAYLgjalRtSRx
Xap2MiD9ULnda0ekO1GJsHVG5STuiQW1/zjjRc0ttAlJAsQueYgnEbdUPhO4MJn7
DIV/SPI8xCrOGiaEpMky7ItmIMb5KQRxW8A9it/ke4ELgZ9fXgYHyCnrQZ9iLN2l
+xsAMCwbEoDzvwtUSFRpoWprjnajQc8W33jTvZgvDU6j5nVnOm1NU2Z7O9JRBrCl
alK6RHuoUqJSc9MUhc6q9ueT+o05VOxF2c89DzOML2BipkkKpdI7a2RBrMT31rMP
P2+UT64nN1bwWFyoLaaLiOQS1gaYf1vAoYK/2nrNBjE02jid7oIwrRw1OJgCTz+i
BKiU0xQE9OxaSnFy1QpLkWJcC2h55WrT6Rg/3f/viqSIz6oKtInC8FKch9O/YI8s
vAstHYU9rwxt+iU3nhJeTTMxdN1PLIV8wNQZ+oomafLj2rlmsF+Zo6R2pzDKFPNK
vAzY+hr0rjb/LDeTWF2+eQjugItmbe2vh/NEkbrizn8DlnLWaaJdLC6YFFhWlkW2
Hr0zlaMi3qyZtmRwyZEwe1SindiFmeDDN0HvX9VlG59zT+ArX0fv+fJNWgj52mha
Mbygo+FxUIdPZbFXbEwukpGzw6XIp4eQ1GXlr6C3PzKefyZvGKA8mrvpmTMvDj0C
iNoZ7aH51uxZFeRZyVwrR+IlQ0ubk1KKg5oPSBnH3s87kcqq78cEPy/hLfVRKDcG
z8AOQT5mQt5RZx5Q0ecSqf3LzNTYhudF+TPK55+Venmuie3c16wkfRd78Gw5SfNc
K3EzW5klotPr4IErzlU/GAxjREEA+mVF8pMsN5H/zgrhv06jnm9aXqoQWzqOu1Fn
i5WhjQw+7xmVL0GSquZBhegU4IaPTzgfT/dJmSJ5NxYwQ6iUnhhhHYydVlS/JmXx
C1QTUWmA/jifnysXb71cdEq/6jSlwz3kZNqU9VbL7RZBBv6RJFn+U/4MJ+VKszum
2V/uvkOiiUQkEI7TcvqmsES70wctyG/5VcUOqDQUCqUO4caN1a6FFVcWHNqV6xxY
qn0LJSJa/dHA/pWZRF+z1zXsb4QzjkRzx9l0UEMeB6GGxTxfu+XNQq6coznN55bN
cDbwO35eJ/T+g+E/Sno7dJNcgg3uMPGtUmArbTL522k=
`protect end_protected