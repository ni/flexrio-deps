`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 43504 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
mIGTFnoSfwcHGJD7pA2OazBgoVduXn+Ma8Rm4LLWz80fsqTGZAK5HIfOuWU3PkDT
0IJ4tBZRJuDxGnFPXvyAo4AxljKuDqicYUz8K63RK4JMIMeYkvqA0X4FpfZvd0Wv
yH6fF2BsfoahkjgqyMYdafSl8ETDtNG+dWOBmbQ7gSg9m8TfNbCA73W9pPadPnlB
TGFOS0gYihFipZznzRnZ5uscVXY9Ve8OOZVD05Xj1qBz3RJHGGTKrbCdn98pmdcx
BjyAJMmRaYQHQ0CEdoPFoyx4cH0iHQoKdVX3pOiaZIwtfMfZFCdcbASx2hrANTEc
KOflzlX2gn9fj2iDGE0mUn7IH4rtOQSz1Hbenlxyt+NREIviYBszeWTzVS3cwmn4
Tewqk/fETbhgbUBTtXbxKmj8us5SzLTc9BDGQbp80FlWZN9aZdZalnvUIqSGGe3v
eIfN1u9cDJzYZaSXNgZUEIcBCO+dgbQTsMjvP8ATuQ+HFj6JU8UqRTe+SROnh06r
BQ6qEs26efVARsOLuFlEd4O3nnMIaKM1sxONwmANwZHevUh289MY1ZXjl/gbsscN
D8mYoAbl+i1ieClniihrNIVtrZ6VLJSohGr+WS5RcbELbvESfYxuF9tvd09jFk9L
+4M2bQHWJJdeBqu2kaJ7hO/lOwSsTPUMHcA7A1MTY/3lcHMkDdAWPQ2gMj3HTzu4
/BEDVh41ccyuCdB8dP/ZSRU5W8kloPQwar6M01rwq0R/feTBfumRH333P539JiFi
ciJQ3rjk1DbzDifF55rGPi1JG1yT4TfUqodLv9ScIH79fJ49ZT7llk0GZCcwOeBF
c4nhX+SXkfBs/mOfZP74G7bVEerNEESjxQgfpQ+ECZQaG7+tdFpe8+kx2BB/T7Et
hgndpj9QBNQOZNNn3+CjXNTyxpOYUv8tLS557c045bNe2BonYhUILvM4a8rnzH2u
t+zTLRjsPn93OCyzp6b2MsUOMbMQ698bhvHHWJlblh7B7+5i6dRMJW5csOHMmwv3
QUimWrrXw4A/rmn/u9AjyMFTWu5TxxsSg+YFoFeMUajHmcqRjZ7f/jUC/oaWC6/i
pQ7V1gPTF8EfqAEaV38bqx+VJSrsiLixz496BHSELMUAxS5KjrlFhWt1ikbffJo1
SRAe0iZsC9ezVygE0q9h7ztPvfK+yNcU2tGN5BA5Ctnzw91mMFJ1rzL77icWcY39
tkgIu1EmQYigReA6rmXW58BgXKjcZFMgpw5UMQoco7hzCC2ITjaHLLbEf6Gr4eKF
wdOYAQajkIw9TyBIJNxwUe714CRQvQpopidlLd0QebO08BwtVyhy05a3C+k/APuI
KgZJbJrseV/M1GX8C9A708quAgwBCNwE93zopm2PiCZSAWV9yZQQfYkrfF1oJNSM
dFqoZc8snVqAAYbEeNqeX2v6rvMFTOt1oCJnRevSM+TTFKwWmeWGS9aMbuy+SvsY
jFClJMwzbd0Vn5ehhm6G3/7M2hqsDwR3kYqMOs7f9zCT6U2EFkObuaw+sz1vXab0
UXfOvFE5gMHSHJ1cJb43HavxSiRyi+TOIf0Dwxs2Vl3SKbH6/YreOHka7WyasIS8
m5JCL3lC5RjNZPqpHlfJcK2iK+xj1zP24xbAJ2BVH+P0SzJ08F4JBgiEvJMTI15K
nCXMdDIbOdRT8sFF/f8fcoJdWE69fcmUcbshPkWxnTi8ojWqPjN7TNCeoGL6k8Yf
8cRXRzsar+uDbUUcseU/PcPNw2tLPmhLDTRU5AchfcAqw2lMlqYe6/kRTzLGqWf5
dAiY1/p5LXwCdA5Jqn3H4NO+4pOlGPnvbQ6aEmelfQ5x6PqOxm0RxS7AIBVK9Fii
qGFlvbs9v4HCakEyrBfjxpd4LuJUbPmIBhZC+dfP/9bCk2LULEr3eCA2IpNDOr8a
scUbuz1gH6tPCvJ7z0rNiMVcJ3cDbKcTP6D1nj6PD54kjL7aRAos+NIfu4MaKt5Q
4oT8OqPhcag8IitTVHbQ7BJ5davfBxDa9u5vmP5cQUlZJS6Zfxdr1T/YlE7SNrNA
IyhtJ4NC23berw7kJaIztpnuMeB716XzGTKsP/nqLbqp1kxJehAHhJEKnyyxPczV
6/A8oqTQbey1qDysI8+bdQbqlCjTSJtffpDjDLNIoparDDLrw44wfS9n20i/Gl93
tS4t1YOb7M2WKu76WEk6L69yuOzAbYUNzijEIyWZI8wtkGYX0WuDYAteDf+cEi1Q
nU/oRPSuckIqADzPgz0NmxKG+I0fVlOHxkc2m+DE2BY3ZO4Wjuq8kErYgk9NVMVe
1qxHzW2rE+O4iPcWCbHgqWqz2/SPoI8zNY8ZTmIHYvPpaDkaS/fEZ82+3p7EtBUt
zh8IUZ0yfyxGbpEtnSX3eVr/3Flk7P4u5d8ZrtyA5DAdCXzWmBJlnZYWs7VA9Go3
/QJXEGDA3ZDm8tCpDXrgiA5Qu1ekN+eQtL+3sTNhpkMh/BcMtSqlsDyjMUjcYHmC
EHmG3DISUSwq0m62A+kgfJtaODd/peObYZYEgdtQVnbd3YqNpn58BTNisKOnfzrJ
OWkhO5aojEbNUvJuH3SD57tsEi44uf0YfLbcWBo9AiAvzWkHdjVfjE9VSTlGN/g3
C1+VrnDda6VtTDZJVDnYHAEJaja6Y/JoIVF91JM4O+sfZa9+qlQyTkld9U4KTzmB
gJ74gq+I53rNCq+N0PnmIJ17LxstWiD9NaQdJNGCeypDyMTzp0dByjiR8TUlNRVj
U8Ec5OIrrDc0EObn7WvZXuzeyKJhjDntlqShLO1e5nnGLChxqdbgVMOqw+H3oBc+
31CPJht4I/lxA+SuZh4ArGXZ/INoB7P6fP2H1ujXGsJxWXKKzoU0r8+b7MW5RJeZ
k3IvFrHMiePPyp+XmpmZd9sZTxfj85E8692lAi4bivQfI6OtOCPfAPX9KcSdtSoQ
7xACR8whE/ws8sP6VtZzh/r/Zqv7FEVl/DpmuPVCn3JQcifql1gPokG/haryXb7R
ebCgbcRnuXfZty0oNsifEZ4toHX39tg/lLIctlXfdSty/r5ecsea1Eti1/TjLPEF
UaU+1Xe35KXK1tUmZSZp8Ms7rmBUymr7/byxKIlTpLaHGcnsDGO0u6BzAe32pPt0
lpP/z85yoQTIbXxDy2QDvY5k/wvLXATp2bwwLbrOeUZmMxESDiKnlcUPQ6mfws+K
QG2zsA0ZguW5Z4YAooRRI4O/jOQRN0224QwB/HHGfOI94y68t1XoEJAv0LaJn17m
a6Nxevlo1fl7WFyv/xcwdW+dYUVcVL9Kz3T5KSCmphog/v2j0/HukG/GpSxDeIO/
xwBYYl1lmswXpnfpS0FG6mUe1Ge4rkGVEFMSa1PieZGW3Seb0IbF5cR7ZDw8Nngo
qfyfpMKv64MTdIVJD+7Pn2rDaU4RV+N5+KxX3s0Qe9eHAUubYUNTcnZmYXkgFONj
eMyUCvapODw6Ym2/QvTj1XY9RL0fF5JsHqeuY24KdnrJd4QcIPIQiUckmp+MkimU
cNcNZcDZo2Li55NHzY2HBBvNMVMbBv9g/vHDoUBBMdzyRB6hLQBeDgwce0jyQNK+
F4SWs07h7c8HGcy820yFPUHP0WSiYyPMjO5/gcrjptdKFoJTVEsdVx7a6Qbd8cFp
9Jzyjl4N8kq3zki1jD90mphkegCHKeFp8kRPITFj0RJvG5nL/oLK55XDe8pdCpYy
JZ8R59iLERDYTpj4d7jD2zIx+a6dsNhu2bMQy/leQaJw8OiajFhGQWM8Hbh2zTsO
DWKTPuhWlL0X3Yy7UUu8TG6QhVayjFSv+zNzzbhHMfqEtZVXmBp9QSYBlNCjLKeX
QfXY5S2tY34eyE7T9ntWk/jVR225cyaYMwEenPhNaoiLJmARgQM+iMce7U0HKtHU
hDjowdezreLk4y0NUl0KmqhXCxYvVHMbkSYH8lV6mkcpE8hGl6MYR8VKss07JDre
DYQLWafHuoyatQl2fGb8l6vYtgRkjD5kFEVRVwQLBoODn5MhmIClU+0iTwqVn8vG
UqiJLbVwJKVB1VX7H+FP+Bfvc42Tg4JZgTLROI5dgqUh8UehwhPZhedHxwogSxLV
C/Ilehg4KKqydv63GtniIIumkRdA4EgjJbiWHDyITxjwl/OxzmVmNQyFtNnxGyrM
yXNXLH1e417IT19QrI2N98YVPiGT7y8gkAV9RkokzaFKPA8FSVKWFBTFrpv1m7ZE
k7idTOmhYuTNmRu5qBRgAtDcfRd8vGzrBx/MCURF4OKnl2k4lmrVjwCDSCONZZse
GFcfcC2JypdXjY7UPg2L3xbFapDwd6/LbQjPE5HUVOaEIu/ixo6lA3l4vBUy1/Vc
4hpNVPnSvRH4qhEHzW+AgZOjxylaEsK4B2RfZN9e8tq+eMbqYbQn16h06XAH5/2g
+PbGyANi4nim0hkNMQ9y85b0nltdlR6UV0q/QNTpQNbMClKq8+xjPufwDqNZ+Gee
3gTIueVdmzFkq0p6uK6TCgfMgB3Y6zymqQCuiMc0qpH2euBmIZLk+vMZEHssjoqs
x9Q6gVhHjcLrwOeA/EjxYJDgOFwT1wDw7td0m3Kfi1vDgU/3fRw5pfOMnrmkzf1J
aPtbflqKYCuHbOgNflzLuwsOiSIKl5kTw94DbWwR8BID7QJQgsxKFnKwM16CGJcQ
JzmFMnn/wLAOrzCBG4FBNa8MKNS9DKewg7vHlKWZZ7G3LFHP0OnA6vVG98P3TQad
sP+Ooavsl36xksFQPLPGbyjX/QjEnGsg4oODLioldfitGzBuSRlVwBnEm8q4UReP
zKBHiaMIVktONOIZkXldtKy4u1sphs5Mxe3o+3F19AxMWpSEKgjRvd6Tkey0tubD
Jb5qWZokwQ0pml/cR0x/GhcGuTRp+EgEsipD/iY2d/jp86OpZN106/BXaHzTMiYx
MydZ8CiQmgO3vBYBDlRyqUPfYm3WJbT2y2B60raTW4LtmqmQF5SX14eHh7sTONhW
KUX2xi9K2MEHa3yFwK/cxJCCQszx3e8SoXJmCXzgVaLTf6RCfy3W44MBUMAOVntG
d4xdZCbiqrCbcrkTqM3lJpfvjEQNVuFTKMw0yQk+6yCfFpIly8EENKGyNGNR4DlB
5tKXF9qeORggNL9TLHO4dh000U50+tVX4T28U4vOM4tP4RwHJUMP0ZsdMz4dWA2V
SZ3JDt+FyS2pW0S3aKduA9a3OrkWLQiR6hgmmSy13vOPHIG8Z/jbONnIm+Tzmca+
UHGi23JuQGx4LSSUitktfOBGyIvGNdwZeZv/PxzjMvmUoaMmf1H2cY+D9zVtu2sF
eDLhIU9giqHQI9gUlO3OTjgloH8+NQaPWQSxK4ZgmkDby1eEDHIXJmUFLkRMFIR1
8OdOIK9TLm5e0hOiIkSRPvqLSsY4b8fyO3wh8eoEH0SL73PnEo8paFL9UIJR3iav
1SiYIalUH6iJmVJbPEuYzb0P48VWZEswt6F8a3VZxo6lScc9zfP5GqbCoeajzdzc
vrNouJ637Rcigb59rz6aHZn+ZeRt/tHMK6r8IYkFbFnuIQxlqLtrxRKKj4PAAcED
DtoMVzc/e0baHmrN0aqfZeEoBulmR/XTySAwH6fQQk8F1ldvXMe0FMqJRzOiYrzn
Mw8q7dx1+FHfQvDABjRN36K0O+jAaUuM7GZ4/bOAv3brhyjZrk5D4tfeEd/SvFUr
974Z+mLhOT/cdnb/YWl5a//wRQ46WWjTWC1SjHWFFmdREoGmmF00WNkOm1IrKMDv
9qmZo0yuFsVZC3E2XTDj195PPZ/H4r3J8agMkP45r3dz53KS9UtFOOiQH6jbI/qi
ZbgvcqFqJIa8sQiNOoiAjXIPa3Wgn2hX/TK/dgwCn622dMyhhEHCMJazROJizDVe
HyXeUniBKeXaGbWBnWGgLdqvMCumnQnYLV3VsPsW0Fa/z2ACIVZoRtkgaAxqO0Nw
42TigDQcUHs+huNdS6d8YJ4yhfRffxHre2JWH9znqGPEhvb7M8GZUZg3u+jd9bJo
TdIdQBOkdasVHyHntNU/2ytkGftNVfmuQ0M84bBwhJYZD1AaD2wYhoP6+MFLoMqs
F+Y2nWlEjNhZyvKlQsBbYYH9jTzQAtKxMbGSsJy/4sTEVy6xNvYvFHqRfmZQS9Zx
tUMHsSbr7t59o3KKH3j61uXRqkJPrMcs9qWCf565i5wu+rt8113VdhGVZxU1PlH3
PP6unwFoga0Q2tLN8xqbFoKn4rAAY7/71GHH/oZGfV2pbJJaV9jryQQElam7rBiG
yzLl5T3sRWj6yb6u3gDeSp6ec0Pd1CF0kNYd1L4M1+bwb3BlnSd9KYtdkiTJLyrA
4ex3w5qdX9mZk9Ip9K+YTR21ozSwmc36nZsTHE/wgZOy4B3DyXckWUJpS2fmJcw0
cOrmBAEiVG7BC4mPluJ9Sfv1OHegqx1iIuQJkBmV/9hgKr1nWVJOlKMA5qelO52X
tQNFZ8uw2pV6UZZA9D5WIoByJFbFdy3PpbIsrOozotiqHJ8Klmx1yu5ICr2hMOGL
1fIPdlvNqWwsWAl7OMfoEdqBn+Kw+KzqLYI+Q3+0pb7deT68ulOoxN7WccALa1LN
OZcS/dns35r3qJ4t0OydQgOz0okxUsiAdgvMfQoN9RYHYMZpSWdyLQ/uDep3HkGV
tlIIF63sHwcZ1jVG1bxWzjibm6ahLuDkBQOOwmzBV0IOjaBdZMwm8Er/hXgSNV2q
5ar/eVpMY8mmD7hiifBHUc1KlnIw6OKGES3I847z1s66ohvBRPQzFtZLyfaTlO/g
bcDIpelzRgNYfrP9aFG4Ut8j+KlDxZivQ3/7nyryT9KJCnASb506BkvMxFTUhIub
Kqumn1I0pNOJoGEXLeoluw++a6N5YOv9PTCEQRFoqLp6Kc9YVwZtEytr4K3KXG5F
nNBoSOpC7mWegtU22xC8UiYmFb1w3L0DtXa/8q3tNZ+Z/i1FPJMCKvrAtDD2UaUR
uDZ95U8X8O5pHjFcNW1o6bWRyuC4c4jyn2cWndWgUnnhlJ+ISRa7vSz2tAzNWlg6
zWuXmwompT1aGVWnmuhUw1UNrOhfp/OuT9tB7OfxQnQd2YHVrL5eeawAKbbwbURV
S6IyW27MYUbcjPCGklPq6RzJpb7YPIm2qcN1EYmIZytMrVYrZlveNLmT5MUz1Qhb
9F1ifl+FJHa2MeIpv87od+YuA0lNGLU/xZ7klgh2SKg0DNLQJhDdADHCX4bi0rTq
CR9YUExrkqqqMmXs7e1A34/DZO5kslahTSUrVf/V+IIDzG4s7Xn5A+hXPRXAqRoF
8ea8xT/ryPW8pyXOOowe9EuAodfqtM4pDZnYNOuOKoiXbLM6CITI2c3dmJPhopDa
Smy4rQbLxuiiwuJkJ64vmvQEPGleDzb+TjN7MCLKEu8+gkAWkw5kvnyk+Fn1k4Q4
7HbOcHvkaWamfCnAjRHm0XLsC36GbMQhObbzAruUoy3jwQfOydY7wcbsd0xgWguR
ghVMYePT2xQhpzb96evXunTIsEzikPuIZnh8Ifyb6OHD9XjVsvAE8Z+/t3Odoue5
zlFlbMX9qaG8Y6G9mQAQ9D7+mI3R9Jh/Cv1JQQYfGNYjHwtWKh0BzgzY5VkAXyf0
oRViunkDpgG8nPYdeuV9N0wHQJhFjEmZtm8Dy0vntFIykrYvDOrVRsFLGl0xkEq5
gmRtnv+oU7JAG2b4B1XGuJarLvcYFKZRJBA1nPjo76lrIglI2U0lFQJ1MMQTKMWU
UPzppGhfEiits98J1kKbLDZDHMP9gvMx3n4dC3bPaNqTO9JYB/tL+6WIOyHJAEFN
1cxkX/JlDN26tlFon8RENH69zh2AvZuZ8ixRj3PodNJ2XMKTDZwsbd32hHewNsr/
JazEipH8no/kMQssJpToYzVsJPnh9fwGHirge5CG/01jCMOpC2raCqdiM72BqAx5
yZ5iCJAZz1NLY4fgX0trk5LsVZ6ezJyCTSNz8s9uaJC7LVKxcZ+wK65A2oIEZr1y
6oRRYD+RpHQ+fBf/+U9uYpdqEsItwA3YC2A2+Mdqz6xe6tTRD2pvROLQwyDMgUud
LuSvBEsZdY/Gz4UJOr3pC8x2H90Ppy0qbdxR+s8eu8leZc7z3I9WybmjrLkp9GEx
6o/KSWQNH7r7GPuwAvTJpQfLUgj5UE0fiKlBcx9u+PRpk+/2u84PIzQ3fZF/2BIF
D+ZRGAJcqstLN6w7KnVoBHJE0bJKtOFqBSRAU5AZHMgNVvQH5L1ImJPHN9qnXS3X
ZWZq4QM727fCksYUiPYxmTKOCnypywj/kOWP4pZK4oWgljjpOl1N2JP1GyeKOc4g
xw3FvDnv3Lx4mh2KQYyrxxs9495+xfzqhxTyZRjmqXB0kLvfU7OA1mySZ3+zZNM2
7NPWPv8nOQSBplMtzgV65RkgKCsciHhNaKQymAvvg3Vvs5OrXXnmTLMfxulG1AlT
UUB/5Cy/Ny8Iv1vUyJAgo1r00kxTUdA9qWJlyyKG5KEM5lRs5Zh+/60+3vBsAx0O
QoG+GnMrrgD3IHX2G5YmyAc8Y8h3RXABYy3hwNmvJc/Wj36SnJzsCS6kzYBUPYvA
jxgYKKZwSjMLon3xy+kP0VHHKoh0yBf46nMa9OSfF6tc70M/5qP/YeyUJ8mZ1YNK
FFA9EaY54kG7rIHZnJ7Cz86gPNlpo+YCCqcf1S78sY92UxYLmjBKNfqctWQQtQ51
DhZDBhc6lyETOLfcUP0CRT97IYloKmeVgTXKv9I4cV7CN5/JpmpNFV7Y7Qjg89hG
Z4MCLJlA78CjoeenxlTcv2+OrWFXXAmYIpvnLHpGkFSEixkufrlPP2DzUUn6NY92
IIdDtat058k5al7SaNURbEiKAhIUGLC3CpjN1TZhqOpVPApWcZ2bOOYamD2I7/do
yy6zjYYmY7GOVZxnsrCs7nU3UlRwglhnngKI0qjXaKp+a9YIhOfYVC9PgRjaEBhO
bGmkslwCkkvlcHYDteX+6X0YuGoxtlgZSsft7YvnYkz6VAmfMMf63XB7pK9W+l9+
k0R7tz5T7qfgMFn3gB5/TJROiKlkc5OvfCTLRQK2wTiQC17tmCSN5SnSM+wR1Kcb
S8Ctp5lORYvQBKl9m3b/70sjHGqP6M2Xr0D85m3XOPS3Ufesf3MI8Jo25Gf2Ao+A
W3ULnQo1F7jS48/fIJ7ou0rUVMwuDAcFie25/Ldjr6ei2P+E+MAAaA55BnweTR2s
K2kjmjI/c93047GIEr5iMxNjQ7xgqPvGEwf7BHXeht7UVaYqvEOqIDzUzoNgWjFS
ePNNpZJTxYgXPBSxv62X541cEnzSKlKE/YzvT3OfGP46Fb/cwxjg8If0d+VL64Ua
kcJwHpgtdUTD4OeSyUqAfeLcwOxaXyvxIY+LZ8DAhMF54MfRL4XZjuyssQQXjWRR
fVXiS6k4krN65JRL7Pt9KytvI7qcPm1uVYoQR8Nk3ery/tLAxprums0i9zXudNes
Uf18U70r+2w51vEs2tNFKPzZdzlZM7e+Ncgzw/C//HEznClM/bLN/xQIOzH3NZZc
ryYNbDnC8YUuQuC9Jbr+W70UKiIbEZt/5qSvD24LtBCdrKGrQzqj4IRVNlS5agm+
5Z9LKlQk6/tJaZfE50FWK8kGmncgjWn/fS72ZKR4BzJ5iKURn5Fz8hN9eqzuYX0e
nunXzeNxbe05XR8dV6iuGh5llBD3cEuwMT5pii2v5mislG+8jC9FVUCEi2zrRRzH
euxwuETtRBdvdw74Baz9yjG++mFIkjIeBshxwaBYDA2czbxDkFjIe4G6xniBmyB/
xS8Dr/GqBvWKaFmQMd4PtNMo8ebkQvtBoeO2gczc558ZB54pUg8kvmEjgiMPYpCL
AcvxanI+eYMHwRI63OEC3HZZmxaTPLxz9UetHY0meyeV2NwhnsLmt8el4NzmqmJB
j3oafMNjw7s6aTjzbu9eZBP2618cR2NT8oFigYsV83fvc4DJQTU+E5xweX/zw26h
Jl7JKSVz+aNCDF5UnAmOSyYYaKr6USePe+KIUlhiFC6Dcokzd6RP2btGE7Xg055B
MTbm1yalCNz0DgPkgdQu76aQNuyFGutfYoN5yKqC11gaPfVYSi9vTgEE3BW3nzGa
LCHRP7aXUSZHhkqlpidUYEdLmdKGR9ENaLW6XBH85ynqnBHdKSuCNWRYObO7qQxb
P55v+M1XL6Jsgw+A3nE8F24ekOkQTVAEYIlLlVi1vuD4NegUAACeDOv3sWb1Jbio
6OhBDyQcEgPoqUXp3ncjDNF8R8WWDLhRwnLNrFMC72+YjAfCFjmNmhpNaPtzaT8e
tnzQ7ok8+AXLLemM+Q+NFHBXegt754Zl3/9UMx7bPv8F9IR+2kW2c55FFwthkUyC
fVBIacGMi4/c7SLTv1+yBu0ZO3/cqsVhqnj68mG+hPCzF1kJtvlYGlFPLbneCX48
tgJ9Ivp3FCrWEVj9cjL84of3BUOs+6obCDf1T3Vpz6BYvNPruTsfbScwnXpER8j8
vuaswzpkEP9ztxPpA5RZGJd/Zy++BAhXEaZhYCgrkryydiBJBBWjuBVT1xxlwtvM
1UYhi/Y5ovTMU2nWzG72X791Rsq6ALayonC1uByTQbldj64zCruz5exOvdHNvnmZ
2QNVtUpyMWxf0zaAAkVctnheX8wd/tM2KflknMn8aiGAaIrCHW1tCfo7CPCr7/pP
Q2FCA8PtduvTcw1rjbjmYlRv0I65dBdrueW4XRZ+agi3eG0WsZintAsmhXI5tRN0
1AeoLllt7ZVShdeXxxf4aSduqwTmyz9Di74RNOvimz9HijAa9hPw1P9xqXZv00lR
6nweMtHN/hz11p5CR7pPn827HtgDpzGDVzoUdQ2u1JAWCrAezwbUgh8o5ygCkaG9
TuNVr5GeeYDx4flwchMD+NmyoHYFl7s1Dw1a8KYVRQe26Gdu7rVCu42g7OsXa0+X
5G0oAmzkxocjSft0cMNYEeSe5aI+RJcBKfQ00Ah6YS6BY+NTKRf5P8Jl6Gjc0PHR
FBxYqe5y8+wxEarcpJSpCf/BWCaWscoHuF5Nd23sjQmXPHxHW7AT81oIIULwpHkK
By65bWKUcFyWY8iXWGXCD6XUc3ho0GJIVMcElJDvbNuj53QmyMCyeCoCzIgxIRR3
zljun4+yq+rJrMLQYTq4s8YY5E9tssxkzkWFWDSO6ZM+hPbQVnS6YuCftms5PWyK
IHi4YO5HwFDxTsMmiSOmAAhFKf2ePnhqMr3bbqzhcxCNsTYpH4uwlkQfi4vFjWaY
lPrnZ1q4ZrvNwlOAMOAjKKXO/xuxgWQ7PGOWYswej/xj83SnT0wsOZ6U8C1F4xTR
YqpmLjdGko/5kI8vHTBI/ZP+ZnLxxfmPP1qacU8RgSNlXr79vK1KwUWBKk6kOit1
Cq4NYVIiQ7pGkmLtfd2YTtGm8dEiPAokb/T4Br61P8p2wApFFObI+TLSL4lOG+GE
SnIBdq+BqiJGnYqPpzzAssvcmJvzCzL1V+KxhSkyKss2RJqPVy/z40jq+lRfITVT
bA+dWGW2satFvCjmJGf1yNyCfs67//R0xXYCxu5j6yPPctIfi1MkYjmx9wCfjPvy
vysn9jn9lDgAzXeb6IatxNiFd0FizFrOgbHkI0Wrha72OUYQbdTBTozMHXAEFQ3/
NgyabGqwu5aKzoRyCcOJWVtMw7Loha4QPuCMRjBSFXrMXvo4UrAPbnpX65cdDng8
/ziVsAVNuq3hAkeWxCw5DLiJcHFKo8cWzNcjVhw+PGLXoI4nCd3hMU9PWoTlbBk8
OLoizp8cjWpNUVrOGTTeg7dFLmWMD7cZ4VVpwyMyCA7XmRvDO02ksVnoNrecP1n8
wCHlLw+6dSua5yrA4NhaPO3uRqMnCaG0oqNsLzV+TAF0t3jgMTw2bfmgKns+rjgE
ap5oYdbEiMjGzsGUXHhYLKrVPCereik9jWQbRINICUEN9h99QMVnLyP4sZ17Pdhc
CZ3+aSr0kIKob7NI0IJKz837GkN2GAdJnwJr9aAhC/nFbsgGYtiGC1rAdr3PvjvC
Ztm6bIxNYmv/OsxPcrbqfHtAZ0RyJby5nBxjCRhP1chJWLl+5HFJ9z0xd/eu/YPe
3FcEPSoNQtBQd2D6dfAEBIT7EbumKNEhUDgI9X++Hk9sCDqZIEpS1WbPSC8KlZU7
ulrCgSmdm2GR1/VfvdOLN5kczDAqNHJopQ64wgZi3FMMhu8AngX+giR9dAeWRr4j
0hoNxuTBh/sWbGVdCGTZmWQGwD1eTRXpjSvyMrUPMTuxBTZcQHLwbgx1nx7bDv5v
Cp/GazNlwsvbHZDc4O09D9jwSiRBi6rPibolxLQgD9+wGIjfsBc0nFa3ST2G8u3q
uDwDK0nz8FkupNa9KYvTLodoO2lCvHcs63TccFYzWdsUVo9nhJzrRCeATKqr0Qxd
xO9GeBMRmJfUxWNAiIyFue1G1Es7OgiNzCsZMyFvuS4q4CmDMpoZZbtrJjNDOSrs
3+iZy3WZcEd72MCJpRA84cIF45dOnqNxakztC8rruKWncOIT8OP6ipu35kmyXI/C
5z1xe7hjuDGpLY6FmWQrHwdmtnx29/AZcnpa9PHotXak2rGj+ma0kE8Ps8BcdyeU
xL2A8dJpSdob24DN2k2vgwgG3YSoV4T/mjBI6UNULMKD2z+Qk9dHkimR7vLnqy+0
ELqzRiz7osxSxk1Cl0L8BctX5hYXnlAQBGDVHj+no0rh9onMWpZsgr/wFaX/O1sq
i3Wsy/tiWuegozVsdNIhtnk1czo9xti8184wDTobooxs+Tvag2TVDvEdIaXtJXYU
2Sh6FFZSXozEqJRRGD/w817mk2d8eSyjVSgYraMCAiXgkvTAkH1yRAQYrpJmVCbT
PYE3ojVVqCUIaMjnLj5bKAk7Of2M9aKnSLAEA+mxEJn2dV9R9uQHjLeq5EA+D22S
Jk0F9NUaDyRxg1VYKvkx3skCG2kORHCroQW3Hd8ErjY5SGjJcQqBkVd4VBWudRU4
DlFu7fsQk41SkRgJyuj5NKo2zd/4DYNYS/6hGoFUIeQKdfmNgGVFwgDhlGr7Aq6H
JpFPUXG/oaC6zW2QMf6+A3QdGW0otHK3p+1gtFv/dRDb+S/gPcAjBL+YdOVZf+Sz
yVZUih7WdlRVACpaRQWJUfYYNDcBE6jJHfIW2bWK8RP3uDb5XgZkW82Zsi0/sc5v
f7afD88pVB7X6MIK306OcJIMjYAAY4ZSP/h5nJad7RLlw1cdJlYbaIJHC5clhR0Q
skd5hO501BJbVHuW1L789ZZcs8wZmkpp4/aRAcQCx36dCib6BGsmNnNxmdawCHdZ
+oSYd/N9aRfVNrm2YT4/OWXwtyHVo1uw1ZZNkkRNzL72TvwugDm0a7jrBmvi2LmY
3xIZWI7bCrRlC+mVlor4ZOu/dxhY0PcVnaZxYVFqeoWqV0WGGcgglnUCqmMoq2FB
hP8Lpt1rHdxS1X9XKMwwvSmAeXO3XRcEbnJM1i/ceMSozKmlQkJ/j2utgyYG3qgN
DH3C67dTd4mbMXnk+x/71bFXLC75OGgHllxs/hImq2kVXoqF7fh/KuOk6KAFWM/w
HrhbbVN/Ebv2k9wlY/EgD/9Ij3TlfNUbGHRMEc/FMV5Uf9z/ZD24L3jEjCN//z8I
xNPM7WzPTtNGlU7QRauUZ8s/txW7/jpN02tKa+7wlM8dnufuFem8MMHRwyVqbOFD
kVGuNp4Q3SlIJUjApmgZX5PbUVRLs8QCtyOl49625cqTmKokb9O6jNdv4Ln0ZauT
PnAHzQkeAp5FxweNWb2nUqCmQP07kTuZ8McoH9d1weit4wGousS1VKWorgC+m/7E
IJdDjic4nV2OLJNfMybVgd444mG/Le4fEXGndng62QcnMnmfjF0Bapzr7brv8omt
1ZvCZyAnisEe7d5Xdd0xZvliRzamaHdOUfPpD+cZesexyIgaO/qiYrn2ohReW88/
OKtoCT3r0O0GAft+SorQtFm4pzx+HLRC/iinlhjVaUHnVvBeJpYEJwO3zrePeoa8
1E+dXaRWxlhUgRh1F9r7zO2rbG3vXK6uu1F0zPBG+5CFX8tRAj9lNStcu7l8hlzj
fNZbmzdnHmMklh4Yn9z+67GNA5SIUxKT549oz1TXDbvR2lZKJQ6PTS0CIhQhhNWd
G+OFfPq5HKSPPxctZOEAc+Da3i+M0gI8K1EmhyiYot73+rakzVkVoQ5G2J73Nxcr
TuWEdIUJbdFggnWKv3gltnKhly3DsLU8huoWfDIqcqWkik9Q3Lm87L94anRh4nWR
GbP8pTx6e1/381KVpUFTHbuwWzoC8cVSz1gN6kSdIHb2L120fiIfQkJ+HKF6Mz/y
5QXkhfUDRB9j96yHcu68JiZ+T1wstBhkdImpU56RWFfFjjf8D93mEy9KcSJ5Du8f
Un7ven0jRM70qV8AvwbkU1qdKq9nVXZ6AQ2G1LtQpFRlY7erIRS2xrM3skCfBtNJ
A72wZw4voCSYiJOTBfSaCnKMvwTqfNi+m7o3OWJQhsqJavFZ73I+rWs15SNDKWBU
8vtwr/W1UJoGQnpgoOxA/LOgi3ql3aHFxUeQsKU0xEHus096ghDDbURNPDqvzJ2L
E+VxluvJwtcnbDpxmnRMN1UZWTn7mSL1VEJKUSF7njibexCfZxd29mSmX1PczKlk
ecjzD4vjJu17aQbdYqMVfUmf11AsGv+vK2CSr5JGuxOc+xtjvRp5mC2BEmt12ctJ
I3eEXQYuEMDjs55OYnWUw0MnFV+6Ozx1HK1/nSfGm1/Z520qS6AUODpvSNtvHPTI
9Bh5m6wHbzBHbMQi2pehNRl5lWW6Fut8l8PsiKH09nredsBinTd2W8mxsEDJrk2c
TuIo5MYimR3iXn3MFPvIrpCyflfE/tiJL1mVGfuxsHM/8lCkCy6Bjda1XvhQR3V5
eEMxE7OiWfIuhcZ/LOXsM18NU+dL+o6GfPqUbqIazsl264jTlWijRkw+SZPYURbC
PphTXu1tdKfHDDOVbXRCzkHeIXu+PQ1AHzW+0bmP2sblwK7ybE9v6xQ1iq2nKTsq
wHPzdDBaU2Gq1stQAK7BVtdZEsLkwndhAEHKEFPycps54v4fFV0Fq6Zyf/E9h6UZ
vJ/4onIiiTZihPtCk/5nkgzZ5Qm1s0m2+4Yj5QzkkvTgXTZzlrmWZFh5Rif0Jb+L
fz0QPYEwbOZVibN9eHZLzkBUBJjrm1CCD/FxgL+hMs42ndCPf7AaCMtJMOvN9PHk
hMf40DSCGkvrR5B9ucDFgGqXL8/ATOiJdFd1cXI5nxDjBum0GKr6twLbQWfnreIW
oXVxs/OUmjTLh845GAHJEkRK5uruLTlYQyGxQfz/BqwGQzJwofvFNtjNVGvfkWOF
rbrLxE4nTlXvlk9WcyK6svTBG/9zof09ACoE/J6xh/BACWn0xE+lHC9UUaLITrYM
/eS4gS1KR3NYtkD90jm16vM6oSXXAGfZGacszRiqkqdyNWonJcVGySs3u6vzH4R5
bBL9yWElOmM1tS6/7qmVUCiloEvBYUUkStkVn/oLW+CDFnkG3GNPRBloNd9HSVdl
tYPtclddVEZl9f9BCK0OT8leVSothx+Uun1syhjHX3mNdh9Vpw6faS6XWISi4ynd
1H7wOmwGZZGBhtikMmFUuAe5SlebfteOTfH7qOgRRQGpwccpGgjbqELo6F6mLuZt
FXTJgNyvdKb2MOUmbOXum67Z6L8HbSGcVEW/RSHpRlCCMfnnoRbB9+jX7Ml5PD9b
GVum7jeFtIu9QoNLDXMDdtLAHNXPNHIgVg4nxt+v+UDKhcMg7Qxp+8qbQDip6Q84
nIqzWxoXAdA+uP2znVm4SnPptF3n1bkG7evDth2ZL4svE5bffeZg9COO5pd0rA9U
KkpBlqNUGBoL+/yPJI7DZAGtkWeObWfmisi/eM2s5kVkwcwcAgcfcUA6f2/VQnRm
Yy+GwgOUGRYfsI+9gdnlW0OhcGduaBd0zb3SMGM4ZtoxD+BUPXmVVI0vmU8CbwJI
MOn+VM/DttIrQ8Guv64vqOewonDI+aXjrM4JrTRKt2TFtd4Kf1Mf7yF95Gld4mWn
WKevIDZzYBxHbpb9T6T7gqcyGlPgt/QVlf6TjgkL/NP3CzkswLZS7ntprUqC4lVq
WmbPCXO/zHRvrC1mpPu577ruQswHqZphy6sDMkhOuBRiyJv98S7uaaYW88q7T/bu
YjD2JefxzD0P9s7HHk6Pcov5ohXP0djsJu3T47oUSGJYZeajkSIM/GoFt5qRDsAW
P0+WylAHFzo41B/guavrS9yO+tXfW2uX1YWA7NE+EICXfoEfiLUCVP5NEnwT5YZv
7pI8GppxccJ4EDeMOpNS6pp1qPG6HYA40SAzXzFkFDALnD6rzW5Y9dF8ih2FzBf8
NrceGWErHau9qjeP+n6NX6Ahn2wKF7FdToRv3dnL5DWyHGfh/ONPlqv5VjoJl4nP
Lfa+v47YRRPk8+M8pA2CAv6b1SpQynzguEwX3XLBUChYsmy8T0gY4rAtInk9pe/o
3ljB6qGQXXnd18G17SlJO3deqjfBXwomIvtQiWAGg0Au3fsk+6ni6VHoIWkr3FRd
s7tb2Brt8EWMWAW7tyG2S4W0ZUjlRR2tiGgOM7I0DUGXOHfhcaHQ3Srne1RK1DKc
uTKxt0Bw19/tjvIkRocRAmt0+BNcdvdoGqROHlBirG/mbDCXSoegUkPX3JCGMJc6
tjDr3jklUz3V9v87bL38RnayGYuhUU9W3FEan8HrN7NxFRotcEG8m5RWeAK/UysU
Ps0Sknj4t+RbthwY6R5SQo+wTfgnqzZSZ4Erx4eAIYYWlBB4dzNAmiwGhOY9b4PU
R7ysA5k01osmKwBt6IJUHxXgcvPZPuQb9K6hGZUWsnTJkA/EojgxPaNLNyTBePmK
kp6ae8LPbOeztAMCsg29izaedZnFaEo/u5D2jwPalZiR6YQfOxV9EMz2mUfE/Bcv
tCBN8I1qd/JZxaIIB340bzSMbvIUslvrqtB1u3vXn1q6kQjLiBbNFkNZdqTDaNe1
6tshZkKSgkTYgOkhz3Xfq/b969zNTv1QcByVO74jt/2Ma+0YpOHqL5yDt3g6Z2C2
YDR+TU3L2bVBI+59uN6gqPn7APct3CIbGNGBF+Uta2HF+aFKFTBK3Rkjjzsh/pwT
mvm9pU+G+3IOUFn03YLrWvMK/gZgrNFOVekYIQao0CRdaZg7lT0Hrm3AIH/z3HBz
ymZeJBx/nbX7qW6RjhT43XMg4owlb2MOSkTTufN8i5o3+82xp2oJO5mdgvhhmkKe
mBUNBIl8AEejykAK6dOkp7eeV7c2t59z/tuvvXzDkoI4ZjVe4xorHOioD6BtC/Wi
d1efoEJAP4EKj6KKgXQqf+Wie197A7SNITrTRvgNEpwC/FLqTd/K71dc2eCztUGz
KcrNRMK0OS4g6LEpw92gz3PCLRw0ZAcVdxdvrEoypC721La4KmfUQzhI5wBb8d+S
8PDXEjo7uaUYbactKXJg7cTlWBTOgXY+6459Zxn9bDh2RwCmCp3wGtMvElArwwkw
wRUvAJLEtRfypLwE9ulFRQVonOMM0FFdEr/Eogbr3vk7LLoKOFBKJEKihg+kThYI
T60qJgYXJbsr+uZGSI2TjntSaR9usQtcm9PXMW7YXwAiOHJ3hL6zIeLKWkP5OktP
/HthNLHPGxTjWcRInLOIr5Eqbmxv2YZUieFcEi3XQL2uxysczGpki3sTm8W0BjbM
x0emy8zoRSoGGieG9cl9W2pHJ06m0N7jLCpmvGc7psMZrT/hmvWXPvNYtBxNeK5Z
HjF7AZMUba1vK0FbIgI0x8M/2789BCdsLr6933R6OoC9x2QEwaFGArH/A+L76f/T
ovkRouU65rnwejRoqemK1N03lzIyf+vXjOj62aH3EfZVX72XrcAda9IuLrzWxcHp
ny7ZigmuTONu3z5hXa63BS6Br7ZIQMB/3WSnwsgrV1wftsszk8+n9rXICmqabEPk
oV3SQZ7DUeY08Br7Lo9ZJRLcjzlBXUm7HIHyUZ/dX7oKobgMz3+07O5TSUKo2qq0
TN5tKJpXE51ffdDNVOg9QhCJpYa4NiS8Scha7cMOLj9Wcq2VC8URYtNk4M5ezB5g
tCzP/oLdLmpwLclcopTMSmWUQv4WXvvF051MYuNpiMRcZ6QEK4Da37pbIrIXZkvM
qauVdT63yhUsEp85HdbYgCV188wlGac6OqWCjpmVZyW3jt0sOlnifXQViRce/9P/
Hs6zOBMis9XsxIhJ3HNvHxmFuvgXN6ojX0G9H5g9+CPVZLasRbXn9xUwD2PaQE/G
yUH9Bd0rYzBGBpfWBNO3hGwBpfhn4XW1Gfmkc5AUUtftnvz8OxQ3Cq2/su0ABUYR
i8bIO8l5vRqoLY4OrsQerrw54Tz50WXfZJzmTYKWEFElub2tek1r0fWuj1fX8qaH
Krkn6ZspoVywy4PVLXGqybd51YK3cf0LLa7+vuVOJDTeXzUyQk8nUDoia+U7PM7L
VjQi6C5/tGJLzbqIH0dLxlBxDRjrRR5cT7pRNL8L2dfo6ckfEAEQqSe2USIerzVC
xN/kyeBTtaLLtW+dRjJFeTo0BGAyfADrKSmZF7M6mKEbKcl1o8hD78m9jhRD2mkW
FjbU/OjWxIhjnHpiepLHy6S/vPj7X65sWrvHWlT9XpJP7IsuV4HWS4S+YgcIVkEp
3B74zhVPPFqwckih2VF/K+6fvtn52+6+bl7V3Nl0/e8KNxJlmBDkhTiU/ljVwJtu
nid2V9+BfdTpaWqq4U/R2hap27Uqle+66m7ZPOrtlV3BHiWE3QNvBcCO09woHnNi
fzBXJfZFsWjxMuqy1/oX4GElaN606D0of6lgpEmyM3noToY0iGdRisaoPtgVy66f
AUmWdB620grUdDX1qAQoBJ3crwVQJUUKc7tmWa9ophdMqMIYuFJHSkyi6C24TH2k
kIx/tzNw/cFN7/DgS07vDH22zXMZuThpbGDqp2o68JLA/MLUWMKq4tAEetgfgnF5
AkR/v7K+BN8g7uQSCiyMtbxcPZOzoQJ7GZILK1TqxMrCfmHAHQ1K2h8lXpUB5lYE
h8wd70L4Edyg6LtQw/iEcXjmas2NA3biqOsybZ4o0xNFLNSudO7/yTVrnRMGapYT
KXI5Ke4vBabXOdVmqIhBi95mEkQOsttmBQUU2dsEVhlrQaSH5zie/5NTv5PbrTZ3
nMCTB2D3yQrxZklGb8vW8zAEgfJRJh5W3qY4ywAs5hmdIX5hUvW5HudzssSaafCw
7zG8Le0Wuz5BeGmrLqaVG8QBnu0xl0UjBDjRYuQEbGfOrxvgVXMmeUdnTtzEu36o
6abVzrWutLNaqEGuJV+mPl/a21ihMlqkpENqq9cbsGbTdn2ph9o4rBvPLZGbq46I
wHxT2xGtklpkmT9S3nOoY2VsiP5+A/Jww4O3xP33O3EhTpkkhlT4aaUeRNSyi4y4
jKPtXgZV3Wpsv4DVFLLoedDFvJdHFCnmvtYsjIIzGJo8foC/51KdnvbUBIXu1ipV
/hx1N52YHUD1W21gUHqmY6hdfpJ4Jx+ICk/0KpG47h3JeFbzwmI1Qa+IJrg+wzRh
pTLPwtX4T7dICWneMTRKhBz1LgdgXt+A5xrNs28hNes4Oqy8Tq0qP49BmenBiQ0y
SQQqTEstL7EM4saYaAlmdnMfCqFxPdNQtjpBmHUF0d9S5DnwAhwV7fYmJGKkLkXl
Cbtoe4gPp6FTVdbznP5i5bejLMSbeGLNCZ0zskIZN4SKo5ycfDpiNWHr+4NSiE5Q
AOpmY9cJE3pvWr9+c5pp5Y1OHF18/RRvxHkoElQnd1jJJVHKhqGiINApuDC7nKyC
G3ZC16vOTI5wsCUJkWesp//aetYcEJGm1Wa96Ri+TtE/Y2zIJNjD8gbJSwbGxckd
N6A9pXPeI5ciJOMw6qgd+NE9n0pamq4xDM/hu22WYQIf8WMgfi8ZoBAYYtORcrmQ
GbK3oS7YclCbwIwVyOLB8EFevjMHnV1fFDSbz+ok+CNJJ3ogxOxXYGFd8tgltZWL
iqMllICIi3FfRmvpjINed4XX8wr6vVEO1q5YkhydyLOU9HLoJU5tLw/C06aM1HCl
IvI4RIHSRoQRVXU9Fcn+lncLNEtXG+fZj1uQkESsEAVwlvcZxGBaKBu1AIS3iCKX
XNRCzyJAhmmND/ZOHG9nmpjehv8EKedzJhgldrMBNGV+ZcyzMLoXoSrP6KYIiGWd
u/PTGJ6zgv2edqZOOZJoN2wMwcq9lvcY8Dj+YZOgrzStshQiTL3aUNzXGe4nmvA4
okpNvRFtXs7IFD2IQMyX5ZPJWZWCX+ofZdOBwv4K6Baoy4afeJf0UiBdSf8RuKc0
lDrjQlrpzAINZXjkhOdoVAM0Vt5lepyOH+fItxnHCLPJvuvKeD40Db6JdZrnRdr1
bfictbIb1EFghKvhhWkhZrrLfSB6MpXS9IUDTlBhfCGFMp8NQWYhZJVPPGw51tH9
pVUgULFshy1T4Jo6HnHLSikVbwM/R2vW+0LN/H3wWUeKAhEHgGtk46+LVJ+wrDlk
pgcCLIe5xkHU6UcG8Hqn7ogtjZb0pUIjJwsWO1ejRWbZfGnvtvn4tXruxlMknPNt
zQWWyojTQVlLJKmz/yb9nxs3PjOTaKKYjU6y2gVq2aTMPIu3SlZyMcVNmWaUkovJ
pY4bFKQlLWGlm6iH2PBniBY0CpGLLjeoRYHYptQ+cyvkB+A3plC4RSEQDa94She+
/tMYVpWrQuHpQgP1HyS9KSJ0b9mJrjrQ2ZPK13aE3qCtGaudSYC0KCMPKPMwA40J
TuwwQbwu1VCw766NTI5JcYnkoaf2VoxIlCk0o0lOmgGh9+SwVBc400dq770yIffS
liyQwv9W3tMbaxmBNfDTD0MYQ9aeKAMdhUKMczrm/9nqjz/Au9Gbh29nQZ4bbqGk
NyG5F1xNjP1jFGAkWtrLSVZe9mfzEzBYyfx61/yoCGm4Xxt80CO+Tv8/BW25HmbJ
LCL7H2+feHROQSQOMiLQ9SI9HMwybyFhqmXiu7NU3OdIFZXz06T6k0qRgeRovOnG
L02Hnom4k5W3tv70pbQ159bUtHbpl7oLN4X/FqLOKcw3zZ+RF+BEDZXb9S4LNknI
EdnvvDwUuqjXRdE0q0Kd9hwhL41hVQ3ZEspv31IhaeXqUxLqiDqzXg98q6aKFghc
sQIKZBIEjlHXi4Ah9XBwlRAjrJ4tsC9GSXPerZewekk98g8yKB1URtMg7geQbcDT
6/SzZHkkabrfQa04jZPwoqwO0KAY0PWeqqWxp0hQEefct3MPQoOm7GOLtJECSgIm
6hqkic8z/r8q0CApiGAJprnR5yMK0DWaFHLfWVc7eC1pnQay+ullM3LElhLT6B1j
6UMonRjMAYo1g00cVxff6rUI3UpehO45NEE0KX0M5AmQ66FcdofiiKJVTgmUK9xh
oknveipP5JC9ms2+/fu/vKnys4mfhbGWTWz2wLJ87msL7X9KG406vKsojrbzlE0R
Hdx7KwSTaOFi9wFVB9+D6d6/XR7Cp6XFizuh33YqzXN8tkGKOLi5EwOhm9ZooG+q
9AuSpKpeSpLTHmpjNUm/dZ4Vr2fcB8kYuOy8m9FT9m0lxsLPAuHTqWDKq0c3U/Ba
e2n/vNxYLvQTvBa0jRqqT0JChz/4wiENloprhr987PiRwNbKlbmXMtfiO0ckVZeJ
/OY3itET7HeWFSIrnf5hwhu8d/rtnT/LlAMPjI6hSonEEwbJ9S/DHpQC5kiFNxLo
B8qZGrKl5bfjw6XE7s9cKR6IeS0EFdvJY6flGU3pDnnoknPwHJP/uma6PM206OPQ
qn/lpZVoCHrczGsyaefclwql724EBi3hyB7gtTqqqIdxdyVY4KBx1YPAHdnSI1jT
Gn3akinVtmVxncxcho9mbu1jXIUIAoiss21HNOl1nkgqiQ5ol2FfD29jEpKmaqCg
W+n7EUwivUMt0VYDUuVn/5mV3OWslw+bkZlmiz9+PF7ijNL449khhQkR6DT3J/p6
1XMWz2V64oGGHeIoxyF6dzZ0LEgdxfE6TvyvyCNsqu6HGh61kzFxOSTmI9A2srZd
kUGSMVAr02G9yx+/7ZRsyBEsJ0x5RhGYXKpOnPPOiD5Ztj274p4O8g6mCYSWJ6Av
Frr02+199znZF1J3W8uOyVIaEkyr1loR957mV254AkvFEWD09OMdVPcjDoR7w2wg
uS+SutwYC1PvZ/QZqYsgtM61Ht2gFzz+TOr1fXWZMn+gLsmDw1ruOi4sYAyU3m39
nA6Ln3Dq8K0byShKMmgoGJjwgz6i5KF2ITzoiMP0DFCChLqrbz27+Ln5z2icdWWn
UaRUhuduiI+3w6CuwKr0JmLkz4QI9J3/1FkA/UTdMTJXorSD6khYjJly6g3/QVzw
6EmMX3YfUwB02ZJhXyzp5F483cRr6Vcr72F/4BhnDcHLZARC+0IRAR2cY+bPvEgd
SM8B3a2iryeY/oo7uj0PDthhFmxmfRCRi6UtFfPN9kkcWLxRTVROLlgcxgl4w+UN
Ux1sLF55HlvV1hDQwXjypK/itL1BGriuMBkDsJfn0/NP5DODHhrmAZcx3WkEjNPX
MUWfw+KC07jJwU5NbFvUajUGLEnKLQGCGH3yQ0c2ieRVu8VsiPlQ1QmQh8jyDmIC
TkVBjb7+AtBUyi0wRXrXwVtHZxEb1Db+7RjEb2rx5mU5uzFtaFvXhGUo1HMPx1KC
PB+bUnQOZbHH2CTBlKrqyhxmyabnuzF3Cef3WMymXuQ/xUSiS885jVjDmqmPw0ZY
5szy18sWR9Ak8ifeMCEySVLJDgLtxxttUsOW4TUGTH9kaXcGg6sIyczgVbfcptLO
7XFfhW1mBCIYOy99ZWsHqScO9kWXUos//JKUF0grQTWluIgoNBpTm7b5fX9TH5uo
rCsCGyeIsY8uVfmVMdUmMm43eDfZYbaVuKeMWVpdPy288EnlPdNiAlD+4gAYIfAF
qN37WMAC7YIxb9dl4i1YyoohNi75tOBCj+H4XEkZrY6Hio+IWGmZoVJd9L6AGgYR
pwHHmbq3dNC+DqiQdxEtjfnD1eJ8lG7ZQutFf7nsPgP+5Kn1fJqGyxk0Ut3FlaG7
yUinbVSJqSTYQEhAeTBc2L4Bw1l0TeOPcOXEQNazYgp2Eh0eVqkzys5KBLHlpwiA
vdGvWLpkdLxnaaD8j3SgBQrGthnRhJb03TljUGmtNETduIwqQEZInXg3W8pIgmjJ
wx5DlhHQvzr8mIHpSy+AOpl3+r6hHYsbfKXIxTKy3p6TJGIQ5CPNbN/pzLLTtMC5
IdjkD9nTFsUm2EW6yqD0eptnEoCI69ImWe8hqKKJN6LfB1XgRxhsfjE+oAznzpkj
4WsCgy0QcR2ss5mXm3FYXPXLvdUpZuDrgNzjZZUn72iy6ydQwcALXsCIIPUAodDb
5IZ8H9YTLRUwlhH//ayhH4qhnxMnR9k9/o/nrnlyk+gpNYwBNBin9SZ6Uk6aLBTQ
6Cv1FkrB1N67hI6P+cmPGLWD03vlPaDHXAVo+nQwcJ/KjDPsOX6aaqjltQlw1vCN
pILfG/0hoGay2ZrxQ/fBU0p0ZPE/0FQzXWNcIKvHESo9jRi4MryjTaZ5FC2vsTBO
jZILnIcJYwl3hzu6piDqX6n/uwtjMg3Mq9NJzICCsNjFkcxPvrkzyKTwok8p/VrJ
PV5B2V/nvOjFDJBvSpOn1DW2pGKdtCm642xB0xVnXEQ1P/uDT380QK2NZxxxuyJi
LDscojzoz0szSM3GTkp+yX1XUNtScQ7CSKRU3RjmscqJTuZvV+e4DcQXtNVQt2i5
aMxD6tmyKG1EueJzkh/VcR+Zj03Se82aRhepc026GF85LfBQZt+oT5+FBjgy69wv
RlNYC+aMLCc50n7uXtzv/SOCQN9a/uiP3hOQHi+ZVqFWTqK7tQ8260QxKpLCVHnP
Lf8iAfGBdkIcj9QQYzbL3JdV2qRkXI56gf19DNpdfMVKQj99Cs4LBEsZaMehI+EL
akUSbvigwOf+mHMisQ88i0f4hmZJ0KBLZvn+UZzPwclQ7wLmUi7tvaZbpdGBmxKl
rkFYBb4naH0lb/GtuYS5RcXgtm8dhA+AOIcDxMO06euUmnLJBmt3GGzic13ABHmU
R+OE0I5gyTtIQKeKqcLpT3gIt6B3sjx9Cr8vKLYJKTCuDE5mukK7eiw6rROnVp00
c/qjaADSp0N7NkJazBBlSj7GOksgnnGaTCPsD3WiQ68xDxuAE1mzKXbO4+UcAYP+
G2P1osx9vdC9ANZzf0bFnRKQMkLW5mfT5MhUjEe108VjSdLuoUBehOvbYYcgFYhR
9LxQSrNVLaX6qV1D2jRsw1rTlgLFef4wh3WELodGdcx+GN5r8F3wQt3feWIpoZfA
HhrxA4NWqiymBYhnyaMBpmAy2idc/r2+GfU85u5uFguFAmddBbQGK0qS8OG8zmnp
IitaezOBYyDGe72gLDt1/nPd528jAjkHyhKCyPkHN5Asv/2wLLJwDTCQKKQKV+kB
lQTg8TEsMBcgJf3suoMk0Wsp0X1ch4vIIY6of7pNhuogtZuNp6jQRCmZARg+6OF6
Cw7wVKCrxnSs2CJCC/qNfrkuRo9WRuEcNLBT3ovMDn4pzOHD9BZY1yay891sc+fO
CdPg/Kpi1T+em0xLzZXU9wR+6leU//CUfC88oK+AHcqhP6KZFE5DI1XC0zRwxClL
gnai1LXeEttSXGh//C9Ch2I3ScBW/ThaLHskZ52v9XA9vCZYnL6JoYQ0dcqrYsiq
Fy8zVcX/7LEi8aKKSFv8Zc6nPSbNQx2KHC6V2iiF3IohAMuTq+ZnJLo8cHFVRcox
kxAZPe+5jB0hqVstzlVscKl+ibsG9jsT9Xc5871yaTb2t5ZO2kveFb/TYiQNJQcP
KUAueDVHvg7i3XGaBQRShLvX7DVN8oHJpfb/wW2QujSuPDOgJOUc0GpbB2tFcxRe
AlvEUYl3WF/lb/yyz/t60pSDt2EZV96uNjg/WEqnFfb/Hw6Hhs1Jq1Lpjj4OINt0
WJ+/mpdZiz0jcpSCPSTiEqyGaAbicBsrPX+vcIYh6MvG302CtOtZZODDJQtp5R1S
W3v1fCC/E7SCxYPicV1YGFnLqQvKKRs3ni+sGMCCmaOMs0SSAFaO9HNBgwRjM/0e
gv1MYfNgVVR8FMs7ZYqKdcAZ9SbvOs/t+1l9BXAwuwiXSRtDMP/LCnllwM8NtCCI
OksHCEBOmOd85eRCZaUGfqkpRBOE3oEGn8VJtSSAVKOuJm9nLFGJJrO5yO+v2RBh
ayVSf6cKckIaA/Bvq+wsvtbT9s8FVE3mOjXKaNbIj1fni6C7Lzw6tv6vLhpPuE5e
m+KE9cw5Xrzb5lH+0eDSsOCr2Z5HULP9S+hlGYBI5+jlrLvwGwyd9T1tSu37XINK
wPFkNGrJiA7voRttUzWjyOfF0V/dU6U55PwVxvqhj/1bWlM39FfADRiBQCdaVg9N
8SCG1pAkSizEJIkm8foLNPd2V5BCsI1YE3Z/9qYCD3toaB0dedJqXzIDxrcItaDL
BcY7crPDzc1TDhKmtW89sZhfKZGiuHGtegGxr04Z1UOGOiL9B3yz9XezC9JmJDEW
rRxKOrSepEFr1zhG6hViM7ILoJLV5pMzbUHpEHviIGbRJeLgBfbFNCGTvHu3Zcka
Zu5+6cUz7ELAB+rULzJVD/imTcG6yQHsptYDb1RZvcSciY53TDWjf30J1ARaZmOo
P1FScR7eV++4Iufwp2FdtX8/ydJuYZAw+OvEBb4sXmGGxRA4Oq6/leilpiYECwZp
jwWEfThFoSMzbKL0HnQXzjktxHUttE7yqf/X4X5+TkP9BJq1A8vUMZ+Nn5buZosv
JmCWd6/siN3bSwryUdLljFDREXEUK67n/xMBBWiEKzmqFKKAh7vKdxpBC3LINk8T
8nMYaV+nKDyDwUc4vTCnGJfshB0wX9zbhAWQ3hm8TtuZ4C5epNHCvjBA01SQ/ioW
Ityq7CkMWaKO3vTBqmp881JAxdVMClvCP2BNtQL6ZLkI52YI+3qpyyF/mjmLpGJ1
cSU/CpLQmqkGC01j420aOkrqBowmflQY3CGPzy3zTrjVsMQffNXJRm7/USWKcEyd
kY0Cw4GhRL6D1X2JXVdE+RV8Z9eivy1BNiR/rBJutuv1al5juKVWw3nSNyXaw83a
i0hhJc/9xicwlwKyKZEFqM2jcB5XwSr89aHCGvZnTxqp+mnm6piGgdz8zsoG8pFR
F4LQzi2gllCH6+NRPsW9rOdqL0VWmKnq7R2BMN0/jAlC9OKQH9CRCVXeNCZ3+Q4u
/4V1IH7KV5JdAdORBRovTgAJ4/O+6TuNEOO1XR5qZR55VbCjBnjrH5AcfZGW0wGG
UNsrnXBw9wH/CaNZBcB9Rl53+ZnqUn/59/U8HJs5kKYd6Mlz+EbSrTVEgYn6qwoL
eZVWkmW0Nuf4npPuhieElIVKYMK09mlLLHItmfLtXROcHmJ3HlwGPfdryXizEtEy
rK0KGMMGjM1bdPu9n4mGkNnxEdQXgmkAmLyt03u1mMd5kv2ghkUNzOgRIP7iMm4A
WaJKtBpSq9gM8y97ufYVusdU8mX5kcYh4PQXA9eW6BEKfOJq23pml6HiLu98/mjN
TwR68RdzZxeSA6LlRvlkj5zJfufsVipLl4juNJ6J5GvAWrP6NjLn5dsgwYqqDXqz
fUbExzHXfC0kZIsvTlDCCnQFzRT9j6mDwc8t0E55v0qJIb9VhTWALwgcwfCQMrAh
MOXoWpXpI55jD2KGeWJaml36R5cgSNU+ZwYnAotoNt3AH1g1uDYQZSPoFZYWE3vA
AFPs59oJAyrn7LUqso3LC5siBZvk7FKoThlPU88FqpHQApHdpVD/prF/rgVSATKR
U8xKYzHXH+BVR1UATrRh/iRfvOXP9gUnV/HumF+Lt0qnRMkUK40YxcGTB34WC7P0
oTThVBkJ8/+0ocyslSB5YDlMqn8A4cPruWk8iblJR0cgExA30RGcPiRLRxBDny9+
adSzb7xoKk0L6D0qhqiPqTBR7qq/WIO4DxowByZnjj57DVj20UPNa0xo+sI9RK5B
x9iz75IPyIpIz4eEtNk0AQLEie/cqd8vgYKFafm/KNpKD7jqY7xInNo9RlL/8LKu
eLEqkhDYynEWMfwr7a10vfS2ZZ5yD5GyZ1g36rrm0E7KzY9Z4D7EAPVdzVQsZq08
DWMBKxfX3dJrFtR4cMGQf2wMm09FU3qDrCPM6bslgti2GPUTPYy9wdWS5ksdzRuB
qrWXYOfjL3h5lt8W4zG2tTaOjfq/PyUdhw8wXT+N3Sg9SEMI3uzX6NTWPCBjEOdX
36FoQnFTya6iyPfNdaAoyyCmL3WSTsj26+EVIJY9qdeBMS59YiBWi8wscMxK9oJn
DlS/bKxSUNuK+AfFN2j9i2bjoIYahrCp3Bn56KVyV141i/+hIF8wf227V9o8MpjJ
V86qYBFkiER56XMaYngI0SmGsRu+5CoJeNr7+FPbx+ptQezwdUaSoTdgTZ2iDM62
wTNuPnSqSebGRExJhVeYgf39e8ihyrTAx3xIJRA4PeMz+EgUHtWJbqjudUxj43xH
e+duB87DYeHHhrzoB8Mz+VFgW4m+q17PrsXoKf+uMAx5zTN6Zz03q+WBdAKxzpby
U+4au7ftaA+gAGZVRiHNwQRt+HUoq87Y3ppBQmv1P2V7/j0VMtBU45NG79KzW4yJ
Vx3wFkXsgxD/uDa5FsZDQP37B5+SPaeBJ8eFGOVbat79hu8e/KSEL8lJqYIVc06g
u8YPshQ0PXMQNwyPGJL+EgfAKO7UMM8A4Guej2WaWj4zJ1PCrJe5KQe2vF4gtfeF
ZiWG2PJFftfNo3702eDAcpVfaxACukVM1qr86KqxCSGsTNk+NE9wocqnkjdZdvPb
/PBNWx6OjBhbXpMFUESgbBiq5V9PkUncNBd7Bw7qhAKwXnaobdcRf2mQdOeX/m1v
tMX/+Dp+38Rm/EAs9xToqTDtBW24zWzgqQydi6kfdhntdG+1bS95czqEzq9BQdbq
8OJyyskexEQOaznS2I9LS7Y57lgrr/MnS0PVF7FO0g0JL0xxnxkt/Zp/+ClFx8T1
0gZoX/1FuOV8lx7h3UWzsakzrK/Py7nYJWh0dHyHbeWB/oRfflA4tPo5cca0CKzV
jaaBNGqAphqvf2bmsXJ9MmS2j+d5YG9NKzINUljfq0jDf9L8xckVcsnBuVHzJrp5
ZsIkGa8KlSRwx4LTyOm+I5wlp9nbaaq5RfjwHsn9G047iw2kgSWV3QO/b6AVQ3sy
7VTwhyGoAS1zrnnWChAgaS+dWll2Hs/PT36BrJx6dhicIQr7MvGRTSVr6VJnWXqd
6GKmKDM8yi8yF5hN5gPLg6tXSGaMh478uvutqBnrUWGRbyn5INUyFcxrRvEHjyOm
Lyz2Aj9Rugf5PL57jBVGkFkB6lXEs9YKsw3DLWqrEog+zsw28ypjEONFd8Fa/RUt
Nn1HsJymnGD4MPfmVekRtOBScfKn3aF4tjeXbSE2/TuZTMNHoly7SCpJUsthYifH
SEVV+zkCIVxB0gsxdDZ1rgjJlMz49+ZXCkiGjuxmC59V/tK5rbVfOvskcqAzEONG
MlykyL8fnUsPB+YFF8+YFViDj1RhRigzyFRUe1xmYMYOuF/QaP51rMQNLcNl46u7
IliKxKiEh4hShcOAPDXRf2CzJmMl+50f8paeI7mm+x3lemMc8b5wBVSmshTZoYIH
Nko3aRbC8P9x8lC/PYcl/JC22MzxSNQItV/kusXucCPjzQ/DHpOUBsfVdNb9bdCq
44Td8P442jwVXKtPAn4y1PX/xqZ+Q7TkWSvW4MUoSAbx5tNkF0A0lQVcmllIb0zL
1kEW7L5P0yT00/kFLhJkvGvP3HRA4nupgBSrsg1lbyXHJUbHfk0foBL8KSeT/pEX
6zXWLaRRKiLO5KSRXY4uOOZoO0mcqVvd83Y3WZu6uzurxASIf1ubTvrGO1XHjv1M
Ci2qNmUKCrOW6IDX9XwUdMJIwDPKXJ1hW4WC5n6thEsat6nrvMj3pzP8xpZ+3pTr
UA5pPqNDTIgkqxlV1fzSEZw0QQVbBDU1eMax222YPtEsmPp4hIcywmKVQyE2/lq6
vQ/o9QjyWHUZG8UI+lsbkVquwomrjMqoLYjr0b7ExcIuQYcWV2I7cgIzFcpnOoHg
5tDVuwvAbFOiP9f0AAYuows++hsm8Thui3IaKVR0doLxpI+4nSAMByDk00lFC7tq
Q5duMEmbpsQPFYkLs22zpvc8YJT5C0R7OveLew4wqwJIYwOr0TS2pRIl/QC09SGG
s5BJ7jH8+5KvBGGibNmRNcXK13XGU2Vxt6dOMkzdb4N1ZA4VHNf4BNQdRtZ2aJFc
lpMQPzDpajHu8ks2HqYEsvq59kd+UzdxYbP864duiXtvTnhSM7x/tSOFSbRQ/rFu
tgt+7DsbcIMmrCYE6Rn7sqnoqVpy/o35ZkFLg58dSNYiLFwORBWzcN9nfhpUMfV/
QwJr2LTe/Kr07GJirMH3fAqJDB1NsRcJhfcG8adpr2PadHpQE/R0ofSE13oWwUp2
EBSDs77nCMO5o8RqgRAHsCqKtZhbemqfWtpCYfqV/oE9Efu5ZM3sGNw/cwGVL3Qu
96j5guvZq0TOOZr88xHXo4z1Ye4o4urcVjKRezRgbWK54M2Rl9KmbR1Mg/252C+v
uu3/DlF6mV0rTRUL0Sk8RPXKHr5QbuumoetfH04eTbPXoHDeMkkC6iuzP7x8PyrE
KR/VJQzBbOb+5htvp7P1vDZAEtZYiGP+yjLGn1M2QIuPNQFipiTFMLks3FnlVdOk
kkcKxG2uBLZcDBXxwQXDu+F6CDbneDsKoY5NZbbhFEBIajJKXXiuiwMPg4k2irdU
+XSLWcd2LoSIaYrpG9SCxBpno99E4qpu2764j9uougN9JmyIjHQ2+366YsYVU2+s
5eQxGtTAbbSmekmovKe8sDLycd7mGRc7xHnzZoMOx8nYcAmMks4I8sZijdn62cf/
DY/hBOcaYwx6QwrKNkIlPL9IOiFA2tdG9GpXZyUoR2cuUSBoinTBBrRz83Q16lIw
zpnoX0kPlFEpgnbV8XuHJ/1MujEmVV6NGqOJVAUFNvzrwEa3ggLWEDC/HUK0TVp1
l996+Ay3WC+aKvV9bx54uowqgxpz8GODVbfnDoGGpLd/BYTjzsJn5xfM0M7kljYI
wFxIoE1oB2wtWCAoLztCIhuAjNXCp8HR+dLp2vKogE3BekBzvu3rEidpA3DfgBYi
1hcMdu+2dZRlnPXfUfMsGcoVc3TuMn9F41uyBr8F+muAT3LaGbV7932YLAyL3AQR
5lg4EivkOh9h78z69sQK8a6jwOFGFshdG6dapwf2XusC87XWp59JAITd+RDCSLwa
KEsMXQ+VjzITRLWfOpaWdfymGlSX8pCOlrNVF3u/2UHcgZB2valdkKzZzIEjDa5S
s7EyKrKwjyTU6A//glDI3fKJ5rruI7Hg2ZxJpe9tZNwaDxZY3CRHHi3kfB4/qtjU
Nt4dBCfYwI77Vh3/o3ZHyHBxl/UI9TqazJVMtGzapWm+fjm82NHFcUOX359Gjlo9
89qrJXcm59lOSEbVMMbiufW0uqFp9iwXHVb+dv7N5jH7wO0q0Bnw2YdoGtedk5oj
NYP/TcaRg1oWob/+HnXZnwk0ziFQuHjDjK1xqHemQSZyHAxMkwsNk4PMRaWUPkjF
19i9sbDVZBrz+fKHcbw2GoSwFInq3wZS366SNiNifEqdl0SWlN1NHv8ytrTpihBz
OGW4Iio3ddpUgp2EuktQIWlUbMSYu9jiedWOxAP4E6D+YmaqWByZeQaZ7Fq5w1a/
Na3G/3+XYeRXmgMLqsKxkRnYY3kuVmY1r/n3hWjgqiI4I0ChuebPRkc4dHGAIgmf
Z2LBQ0rgVUonc9OeOTgprlwReI2HVO44GpiewNdAlwhgbZ2sai23clbzTFEIpPne
gRVKmBDCt2fiyt61lpb2l//vZDQjdhq5NRMzlbMdZJxYAjcSu1XC0l/EV8dV2Y0u
RCkQQAlGNfNTFYHMd/tK2WvIix5ZKz7NigKoCRWhc8+pS1StCbGqWZJ4RGT2lDVJ
5OEihpzz6sTvEdNc9WZRZtxEA3TOLDgitmJYpsM0533EguOtmj+4QNHza8doLUC4
kfoRpZ4qCJyDtbXrSaaHA0W/FSiErXblPxJVAFIirHm9C9T1ohZ/CAqSRwcUBgRu
FNlT/aQ3aej/1JUZ4vdSzAzWEMpgM2un8TctlJCpt0FT+7BlIwFEmVn+53x4wNIH
o8It5bi5f2F51PM93u599tgqVByKDRj85grcjV9St+i1fIMll3CKsAhz6TpRCZnV
+Hh9snLkUuuYrmtkJAUEQJvyJsdod2pf12FykUkdWLn5/ukMnj2UbsA0PvDrd7Xi
GbAj0V+Z8El+cfTfVJXJME71g+SmdBlF3FWW4apm37LAIxXqDFoNohrgbj0uXKv1
6RqQBAtBkLGtxCvQqL/tZg7/piYp6dddMmjcei4Wn1LE740Z2n7933LZGzLVF5mO
6ijUeeJj0RBWsjSS+j4xkfqLtc0wYDCMtHN/Faa42MLre4w5rhhFVvViQoLD5kG1
42PwVsLOPB2GI1GAl1xUk+vPNlWiQMUrlRAM4hrCsYxkdt7q6rAFh1Pes/9IUDln
m/aKs3U+rGeDde0mhEh1U7fhHm0a5XyXpb0eGRVCoZ1eye2tfckZh8wyqSNbFGR0
wjdN/OBg8L1Pvdu8tOV8XYYgonB5Wx2gHyNfqDIJ7ZCPFS/+fx0JWc2n4pC22vqB
A+Mg63JX463yiwQC7gPcMTA3+F1D+cGizIH1EedH4ZKxcDuu/unYNsYK8605emwP
9JK9/54qSXRL2tFuRcdoFu8JhwCEl2lWXzL4W3FkxIHK+xK/YQsOWXDzai/zDrkE
CIJfB/kgheiF0GJnKGKWt6IB1kZSWTbHaDPFm7kPCW/OBcllkEN+HI38N9Easzk7
glo7XdCIWY2EqlXRpaZTwrcsLPSuwqE3iXlD6yxsYO0lOMtS85VTSNWTODwOCGnl
6ael6xTSYp3s0FNJScD0b3bcB/ciHi1vKDEZblx7uWB5FOTgMqD1XzwB//yR8G2J
3evOQYN+5G2gaRA6NCsqZJRx4/gmcnICPrQyjaHCPesL6rhOM3Fy86QiIwlH/JY2
wW8esoDTkciz+VmIlP62O5tJ+2y4kz+XGcqKhDaMH7o2o0TBe41I/fnbI+XpIX+e
g0F13aRZDFs9ovd5XT4rEFtGNTfnukghUMDIpNdfPhR7pDgh9qivg8yR2dgQa3+c
2D7NYBvddMdps4jqQ9k/7BY906v6v66jS8hHeCGfnVeiqkvipDxSCTSPvNg3ANLx
c+6/RP9iutGWqHgyknVv+hZ83bhMfSXM08mX0vkGe63/en1g8Fzx+HhklzxAlwXw
Drj7YjKdAEEVtjtINSfmXUWIhzWEXnhVRUl/A0p3TbJnAQS67+U5wWMzcr/XUepS
SzZQQdvqf01Uc/KkCI7DNm2GAEEtnZAzZXUCGZVcoG+rgFkJzxzM7gpJf3a5u6Z+
/9fBC1xSewbJ7V9ewskjN7rMmzVB4oWj2HTI1ee7jdIEzvoIVuZ98qpghgGXZXdc
D+gnorn0F393iZoVs+ow6UI7wgS726xr+ckduDdM/Rm3r9xn1q3m/EsM8RK+Tpu/
qzqlUfOSgOM+KFOfYcbgBvmeNxkgAXLLa+aUmuKUtkFjOqtSUp9wN1C9lL0WuZgL
oRN3PnV4zwMZ8f2taqa1TZVaJTK4Sh93HU8oq/SYYCh3Es5kOXyYSVbNzlZ4aBFX
seVe3Uu+q2roLoa7TLOrx7BWwchy4TyRWCDsLO6c2Brz8Vh4v5/q/Ejqe0e/vHEu
4xC20LhfsZVp/sqsEFG0ZPL3Kzrwz/MCIgmQYrVB8xsF01ofd2HfVEvdXxVQOJH2
ZAxBKDGqGvI1dqGHptd0HdrQokEP6WFi/t7CvlUkK49Rpb2T+JF1WNIu8KKn+Icc
zVE8UKOWprLco3RN0hm9E2vVqH6Upq/ghjrjQL8y6IGlwuZfed9kF5lwKOBflaPd
6TVYfBP8mFqgOa9brzm7br5SXgAFUCzE/xXJK03wNY86XOIYr8uFN18CobaJE/AX
7MWdE7YIA2/bcJguJ9sDb2eeHAMPoQBCa6+V4iPBkhhY/MdqLWA9vHbEZGIFtMmc
agqNi2HKwYLjZn7aAMlAJfmua0rXdrif49leqI07q9Qx8wp2UMnp3uZeFhxVo66g
J18uLrj9k1pjHR29j9NtZAkoglFYalDJDv2tGdoYCLIqmn74ZbmkdjMJVioI00s1
IlbBWMMDayZgm/bz0OLUfHc5gfhQH3/A2y6AmPOgzAocpRfSMJalS/Hz7iiWXefU
CpH9TjRw9VIB6voU49X9TVtgi0+pZGAZz+PZasEzaG+Dfg0V447ZuHO6XXZr5Z5h
dcitAFY4PeFpxtp/SxL3YcrDpO+y44glxtFEur5ia+vJ55UVNB7Y92gg+SBjXBVW
ttjCdKqnc1L3QCDctlqpYX3lFAT1I1IuHay26XuK9vHyqvoaX8xDaJL7a5YHoFet
XinrkFZyRlX2YIIQ+LP/olQklJEaM7ER++MibACn/XFiP4wPKF4O5NzTnczOj2wy
LH0j6Ygpw/bj1Z+raeM4wPev0X0If/BK6s5sZD5eq2WGaGkBi/dVmtEKp6bbWasH
wHQvTR8jkt3yc0X5MRgCnnsOdsf7/t7sl48zKT7/Uo0NPUD57WD9GL3WlrQRo7OH
VKMmlA/IwFnVG+tUZB2wxtpM+6ozpqfO9lYW946Kznq/C5XJr/stiITWoWnu+3fp
zvam/KxkeNo8jyomb+l27UaKm2W07mntDVnhIl1QTKAiiuPOd6e6GzkQ4R4wxfRt
KHofmw8bclxynmrUTlUG5nPTXboB2GbhLjF+nIJ4wFZUENb9xw9SpRXv0otOTdJ+
XNozXc6SP+JhQff37MciwLs6/Q89OxF6STp+grDIMI/hMCF9GJoPcLaCbWS4yJk9
oUqqImOiWxOaSInz7YlM11QlRGVPaI0o+YCj9s7TPkNFT9XNDNtc0lMz560Arphe
s+6ic239Ii1QgwjCPz4sKgo4uFUiKGBDm7AwgrEBjlSJzWz6cI+vvwiUqwO//mku
YQmcRo4825tDh6v/ywLzi8zUEWHd9jYgWqsRmSzA1RA+Jr3uUkXo8ckwFypVFpFE
AJNUR4z6Enulk6ANb9a2lYJ2GaX/PooiPdIqBGMCbVNu45QcLTOF7pGbTTkzGz1i
nuOW5iwNnETwr+ZW5uoi/AS3Pm8vEVkqC+OGs5YDBkl9B3ZwkZhU3/Br5LN4YUqZ
jlsNeycOo1qsKNq/JVkB5nsDXNpUWA+PLWOphGI6P5pNb9GqiMuKa1Qvd/cz0a+a
AAvj0d5EmADELCR9cTmxb0Z+Lb7ZGlTcd+yAYcveCkjeDa2l22gpQcQumZ2Nhdq/
bGhHshKWWHGp9wW4FXijsPy7XWiGTaJX8z/ylizYpaGyn1Atl8y/XcoV13q/d8cH
Rwtf2xSq91ZnG7vNHUMGn8I7AGFI+w7ikJzkhhgRBVoBoUfJJ0xdhZZ520/lzOgX
mchsvt/vsDEa4e5Fr6FXdalBrguojARAbuRSKcRDNgtQ+GNkBzHHSSW+G1e4tlho
2Wkr161kGBBM68vjmlU448kbC2L8G8p758j4K7zvI/SrbXt6HgxcXtILhwxqURGQ
km9/rBttTCuI0M+m8Rf3wybIsZf+MMvcfGnmUlIcSsaP329HC4ZETTr5il8IZBQf
TcXAoX/LLqC2ah6+wXDNJSLU9JMtgSJfEcPRt6OqQ+a6d2E6CsatExNn5zj9I1nu
9uMU6X+iprJgMOrSQXqK3znC7oIzJ5J4nWg+7u0mCf0lkmfQcWTAmfEmhYtQVJE3
gbhwLfu0g8UaKTCdpMIVf/WU+rKx4vP/YGxXjrGWKB6b70LrXNsD43AwdF2Y1KrA
lUt/vuD/PE13QgoJ/Tj9Yv+faFCw48RP/gP5ktC2R1DXDU0bWoh8sBOqwVsgIsEz
vjLSKTKw2HdqLTRQMT9+wN99XT2KPtElpga5tVODsV0W0CQur9r9EU+/vm+xnk5y
D/Cpa78kFD6bCu1NVevWMnP0xi8y41WUMJhiqB4lkGn12Ndo0SrAwsChsbp2XQBP
4/Es+D2bOS0vCqgx0tF42J0CnB9+255SDAVaUzCZmaHjq76x+Zou3v0BYaHRWrzT
0L3ikqnCeqvQsDE3CH97wmcn91gkgDB4Y3OLmRveru/m70mw5wT3DVbb4AxxIIog
3AXRBgyoACO//XHnD+OPEz8UrNjsTI5+eeUBU5/WxR6OhpTAm+COC/zZlUj+c/l8
952dDroG15E/ERXjvfWbTpe0+fCtZ3qSTj3jM7RBTy6nQF0RIxvBr6Nl3J/yuY90
JMFl6YHUIAVLW73ezgp5lkOgqEhlfwDxbv4emcEznNj4BUEBHHS0l70I4uC+aT0V
BXJIJIVp9Qen/hHgV+6gMDXqAxF4N6m4TRbRjsaNGBsg+tCg8fOU5in+7W9UEf3L
ctJI8B9QqZ+AyGIY74vXj2MAOCuVejuqKoWVPxvfd5jVD5CMIrIhpeLiNDO96V/d
wAb55YE2nVVsuLHy0bngo83WM4PmSxrsF5YJnA3Ic6GvMiAXN/LMFjfyQj1tX7VT
euzbwyqZqPZwJSN6PSM/k5MiuG/fzUXFFdj0/11jj58bSElC3PVsbRX+lN/acvrc
TwlLgAhK0GyXsZVV7FmCBCLmNynzhvulHn569BJpbgHsg1JId6j9K4aWU1jal+qN
/9MOH9dewi4D2GQObU0AR9A1nG50PY6/purn5sz9+S/4Advi9GOfbgNIRCa3FeU+
AqDtZmZsJyCOdZIEwx5rPehNnY0zdkfC2zg5ckT2i5y+wDCVbg9J2qgFK49SRn4T
SuQpjJEOay6NTBFsvsg3n9O9+YR80LaCZ8w0QIQxPb1cN5wfebsX4RT5C1dO9GO+
yo1cF4qytkxTiiNZdTEC2CxW9QI9CGzhyczxcWEbHM8SB5ADKwDLQCzOKEqTBRvT
orfE2++pW47t+t6+aAwpnj5lD4d05qDIVeUK+oJ0j9efDGmKtkTQQ+nYKv7JpWcD
dGy2QSRujN90W9q4Z4hKbvwY0RxOptpaUPSbRQAyVID73ON1FHzJT92Mg1HH7GuQ
b4RL2/0H3HbZajg144z/7umU/E3XCsbS6tjyIwx7gVth1r4rbIQ7B8dFvgXMIw0L
hQFrKCKwm7+5HVsVHIzfNYITXny8E0DDNmZUJmddzQSnq8NpfTreGOeKjBEyQoYh
qRGeKIfhLj3reEFcazLFFVje0au4byvotDfpPJVNsyHu3FyxgMrtEat06feveIAT
uNIlfiXLVU0Ce28YL20Smn8WMeR0UBq4e0X/TjHJzUuQTu9OWDBoW8TsoDqh0dm8
KiFLaBcn0AlYa2Wr1kBmfMlFATOR7OCpiDxk9nYXrqTO9C5SpP06dw7R04KHFDiO
ajszQJIe10D9LTGGaDfz8fvzvzC33KgIZr+6/69N2r2D4v/XiI2/fbfdnarQlH5I
KX4gQzu07h2E9t5N9QU3q0+tGNeu6NcoQvdfTNy1mQ6oaaLDi4pHPWvRNz4leHvF
QXnCAiS8QLNcXuhLL8lc/tWjhl4VHPStqM44zY2bff3/sJjYwLsUVwl4PSYp9NGM
AMwhBcMdvMrESLp9lG65ju4FkNOedtycBX1bBgs+9Hcmk4HXYhEuiHwxZNYefWFy
C3PZwBuX+LSNUuE/j3oZ4aAGTf7JtX4x1NtNM4CG26lwGokBwRvez5+keciokuJL
nwr7wZUDtdRshtTiBchM72zFqqdh0f7CCnA06EF+afmVXwdm7qRnw4ObNXfqg2jH
2T8/reyH5odMAbsmuaTfwGeAPyK/92GBezav5LzzdF6cY8cEGfwe64pBADNMODtz
sMeWZ+jMCVcqLDnA/KuhJmpbuGJsMVNbOwL3NCDiRzOFQ+KoVUry4veVASreoFlp
BqxcA1sCK+2MtbhPmEJeV5kshYKRRFDyuZlay32rHpSgkeQkzqeR2wmwBaSZ219z
40DzNsKipsG6C7HEPZqAYB7ErsjzN1DtSnrPB4a71cxGAZCoab6yFWK9QHgIK8Hy
khXgsPufzU2cbP/Wk+4DzXTYvrOc4Qz43AMOsyqh2jwkKlxgPwfwvnpKFGPUqQpn
goY7aK0Zb0+i7F9ag9vklQVCwr1MxtxlWihAbo6+g6NHCWXPMTun1GZjAGLzentG
sqZZD42luMnlm8Acf3QWDUAmsxMwamYC1Rlh9BLL2Y/7LngoCD5cGi3BKUgYCTf6
xAQ9N5r3n8TITPya5bVYV+pOhUvOueLvANKNWaDogyJUCe/81xyFDEZMQn9g0Qxv
wZdrmigFdxbIw8mIIguUhETR8RjEfAZhIU8Qir0wpuCjm21tRkzThIfCRr6dLnO2
UszseIuqput3tB2/AsyobjAoG2QkngDNKs/y9e+g0D+CG9VBEi51O4thUevakmAt
0KrLm8ADqRXVtO19V9L1iD4uBo/9PP+Sdzdf9xWtoiEI/w14K2Ix+LhB7SqaP4Z5
kQQ9saThKQEn/0I/saemNt+Q4svEzAfby28CNoOFaBtpNL6G8VHoLcDQmv+40xkw
c23k0Flrq6qWGHWMmjeium+bA9VRjjNdBySRoqbWQ+EouxVk6g0dR0NVd4WmHvUb
i8x1V+dn8wLapI4Z7pO/LXaZRHjV4PjyBYOm+0k8KlFn386dAL8z0R9mwDNnJ4wa
8ZJdTlAluzJ/2HlCACp642EIrFDzNLNkCVr6t6gQqJ73/7WocvxvBmJ3MMvwIhcE
yM6M0XUgw/fxHJuMInV7LE7i/4Yyo801T+3imrvrV5ZIQMcbZWpYVeYE+/qN3fbC
hW69N1I8tP10ofZ/XFNAD5lTPapPmydeQHwt12Gf+DZvmwe9LlMpb8Hj7zmWNklH
awql9P+ppMwrVKH5QDQONHsWz5rax5tjoMloJDQQwAI+GSDLhdtoJaX0DExZffXQ
Vd2YRKBVGMxaJ2DLhBDK3F96VtrZHlsjJtCjce1Cb1Atq2kyySjVaYRkjmQ8/Gpl
/viSBqG/UBhrS9yJTZVlkhPO3WYnx1O/m9YXo0ka0YtHnXh/2UCyAWoZIf44DUGH
WtFwfsP/arnqVjCzcpVoDBQqQbHLZ22Zzk3tkohWpNzHCOCZnP8qhWScPQhAAywS
dlugu2BuExWB+FAj8bDOqjjpkqgU0UuHqEj6G1HlIB56o3qqtempEwiJaeIwQ57s
UBTG+PRl+oEau2aiBMM1EbuAadh7n2flU0Uo+hRtarnlszxm4bN2vy62iygvCEKZ
QzW5Wbj9yJcap/zMM+bRLVMVQTfcWaa/i0eb/iXJlNEHVl+59Kb2cA+OLle+NXaa
JHFzD7zosHZYDlz1Vh1A2O884+4w97KzS23ryFFBNOl2n2sr4NiIqLv2IRH+IDZi
HhOtrDpjdWIIanWTIP5Y0TjoAQOYVJPYdkFD38SZBWnkwXA5zSu8Ls8Fz2aAwiD1
ZMalJXihJOLXHBcX5xL6u7m5rK2AZ4VnmwPHjddZrabaGiqZfRZ86itdC7EijKkR
jBAClZl9z+c04UGubWXhHG7vVK63dUlUpiDbg5tyyO1xpAX3eGsnfRwv7P5Pz0DT
kHwOzPaYTjm50wqM2j40La4+ycv5PVR7IfgFWlbjfDtPggKwmv8SU9zlHXsqpadl
luXyI9s7E6ITyylBMVjrfS/qEcZ5idLzgDj1zqV/aYuoR+PMErnOJMasEixLDP3r
TiVLvDgmEekW1Y5RGraVRBWx1Cc+lcfrB1O+cUrjJ77uw6wL+a4Z/wA6su3QkLoT
+VfsNSVu64MTwNaWNEl1sg8fgNbGD6IIPkeKtkOLs5zdXOkbvBjKd06WjeOnpVur
ZvGe4WMLhfkNGBVSH24oipLMnE4aNp30dFJE49MOvQJWYL1FO3DGddstFoN7kRTy
6v2396hSPSKKB8/RwI0oRBx1gpbVUJqdZpCLXY8Uc8UYSH/Uh78GxIED+ry0Ju2S
oCmp6KWIP0uqvYcoV3teRVgs06tPe4qD1FerKWpHsp3yodvs6fBDghnOpghgd5be
0vnQFZAFN496W5q9dkXYuiJKIIpBwEGmlhvYvG2iOrRwFvRhUx9/VXmAj0vUd6ny
5c1wRJPSVy21VmfwFs12jtddJEKGCfumI+I8514qQvBr82W3eC+y0Zb7GnkO1iv5
OLkSPRWbB1xK2rBQ/7n+BYVBzVpaeCznnpBmASyGyDzJ67Trw6Bda1IXmwvU+2Kq
BkaWdWJcS72EX8kDcC+fVF1etzXwVcdHrrDxo+YiQ90X2mv1TvIcXOCkpvTZSqe1
v1iVucUjpCIDm5Dyc4USicQ17FqPJXxZdvh5c2VaRkjz/V3EDu3PtWB9VfkJ/2kO
rzVVNcpBw9Q1Szda4WBWzb5jbI/Lzc4sE0WvR8Mmue+juzYX9ecRFBRhLrK9vyyT
GvRSK9BnjugQ9hWaIILLbuzDWyHpihb5V9HN3Q33WDxkowPk+LK0+F+t3IcjE/0f
ZE648Ji/op8YQzbDYjEdF8teqQbErXy76OsrZXEpA1acvVuWQaFcUk+R0QCPqotZ
vp0g62lwuRC7Zt2n9sfXc1mvVm1c109OPIZQuMLroZxDfeTIRtAnTUEp26UFGBSs
DV39PJnrDGwLSgzVjdp/7JM/lFQXkoJD1brKMsuqC/0yX4fWxII2Mo2g2z5zWZiS
D4YseS4g299E8AEyzxGKt1GbbnVJtTstuFUmIKtm2rv9tkZNDLgADmUwhP42ZdG6
8A37r0TpWJ199wnxFYyooO08sOYyDPBDiun0mVvr8lMKXScQs5mgVYaCYcdLHcgb
6bC8kGukzk5SmwGDB/LNvYJdsaRV5DFKKVRRZsu7GCsM15xK28BPI7aX4ZiS0pMI
U7PeUvvd4G0v8iLKtFV1HUCEnBbzNjHaCJpSGi7KOKkkXUPaIY2lOnqSHt9F4LmQ
LMCZ/c7wbee59XiSkCBq01A8EAvac1yrNF//Baa8MrrrO5UnGTgxvS9TMHIn5z+L
9NoatSavSS+pn8n7/cxYzH6bKAG+iDkvk/evCnUTXLkND2cVoxIosHMbt4ZWr37/
x054g4Lpz5tscHFRXp8Gy/cJskEkFN/Rbk9D+Yt3lCNUPWkkZ8Llx+2lf3+l6A54
aCOVGbosmaxhZd1vAtaxiZtW+hSRS+Xvqx/TGT2LeizcoIJ0IL1AbXRLMQg6V3eg
urwh/V5NLYDMl9MbunrcPks0JK20X77MOG5DffOgbIucC2qR9GiNCMcIJWTBU0XQ
lojUUxZeOcRjRrxHNH4+8KRo6uZ/2uESEub3mrRT+GMxhVJEpXWpkgBe5E2g16YX
oQQzTTNb9Ip1qbRVMFVpP51dpB9Qkn7n6/qbV7W+ScDptqe1sDc0OEAjsjKBCgRE
kaQ8HfXmTMRPgKrED3c7gtr8lum5LVpXPSJFAkecBM0+ntLosbYPhMSJicKqs53v
zwbIQTKPJa+B/vUCm5vhKkZ2ncdaVxJ+6tw5axqCV0Z9RlcbEf3ZruM7YreyjcuO
NeMtUSaCsf16gGFzr4L3cAJlPgUPIyAvXqWGhnnk2o06j+jIG0gQwcrFnGMsSapZ
R1nJ4eLAAS67inyNqyfLLEbT9MMVsHU/8847zz4mZChq8adywxpCY+I7eUYnHZz5
zdjX4tIrX13bU5eeR75jPmu/hGMbhTkY+XUUd8CDdBUZuR0+ZCAHQE3PYmMu1COw
OgzfrCI3tVB9FjTZUao9AKflL6aISyHX3e3XhVnaY5iKnynxOioe5Z4nW4pq6v9H
te5tD4v0aZU6zB4r21waWDNJbXGOnMyRHSjbX/DcJIi+zzC4n89qW/XgpncWfEOy
oTtzYaOqGFQjsC378V35arJvl+/bT0n0CfHsv0+AQyTDS0e/WrkGLVLLyUIV83AX
+9QoKfC457rjnrmIPLHwUwpQRP8hmxIxpetqEjk/ilsdFvkWjNNjRSc5LgpxTlYA
i+XAWtLjsprq5dmTzVInZG/RjpfiXXzqppU2R7rcYPO+QmtJfrcHPLONf+4r8cXD
NdzWquQfrVaocFiN/MxXUagLfrgg05MAEM2MHoFjvRdf0JwMl1puJV6n3g7Zw1Ka
NMC8eQafa8qOg/1xvWUV0zCnZQ3mkaBx1ajFfji9SGIb/svylP5Iq3KJu3+wVF+I
mJPQvA5yy3CUZ+FA+TIedM+C6e7kShOlVmDkbK+S8QU21gGeHhWNpaVCDJh07Q6Y
LGLoauN0Fd/bWSZBD2jSRfwyStvsYC9tAwi0/Iq5NKDyCLvUjQhrrfpYIjErxm/J
tnx3x96ZWcv33kM5xP1HnZZo+RgbLc9WyhZ8yZZ1UOK1JS7P5BOHYo5pi0BU4ik7
D5wq09HJ5s8I0nUdiMrnIUjQoTJZ2I+q6kp6fbfKl39vh7GJaYicCdT82UzVKp3K
5dQWuStKjNXNGO0KDN9UVlA8hxS5BXB8KZtSOvVo2n26dfYgSuHhvXBlzZ2GX8nB
wJ66FVhsp6CBOdR3V0VQFZKT2tZ0xwNo6yaMKNJBL1c4cw80+hYs5NJG1JD8ZNMT
/n76eMknRKzm1PkrAC6Ck+TM+TM+g7ltDfyShxAsw4xXQM7P+yggVQlURM5aT6aB
mNC04y73Plq4xoijcS7JYX2PejmobvDCrRj0rUxxnOxmnw3/m9nfj30LnZzdcFv9
c5BUyJX5E+XwYGlQAdfCJrWkfukNBfOeYsN5V+8wr7q+dzZIjY0YbNNw9WbsK8Fq
41UTd4d8lkyF7wB/6h02kSR3Ix2JbhydWH1LsbGcMpvOA0U5Y99pbr+EpLpd28sM
SnHpuQJVo1/ol901zdgnHUvoXEHXQmpygPlgMhfNLx/Atq9sUmWyG1FnbtOpFXwe
De5H9iF4j9RoTIGtCLC0h20rl6YEkWqZ+o6Nneg/XprtS2HFCt+ToKiTPIZxiWtZ
grctRSMP6S1KVYoC7hb9bdNHEee5qI/fVrzTFD543YiakYllB6mfGi3jbbtS9WK+
0AqU5l+NBmOwzVvPhRZ7IMiwjfDbz63Msu1qp3PrX9WzYwgqbdemkB2pArFo5YSC
TyAB7LtqesWHSEFyO+0XzIpgg/06yugw610qu0wnABS8snOM1e0T7+BS/7JP7jeo
tkn7sljzK0VehdNPKrz0zB/coMFykXuHhb2DerC81+O2d5QDAAR8PSNeVWxJwPhk
RBumM4TsUjnSRwgJm4BVyNnUm2YwOYLqBt4xK7nbL9KuoynQQ3xzxY8E3/Ztfr4Y
das3xLv3/yGrnXMA2Li2P9XN4tcR5k4/srjCututkesV6VUmy3qNw0C7PCcvuVYv
iI5hB2uUrgb6NF7Zo9194bA9FAmj06m8UUmD2dmIJXiiO/GL4fj5r+6AWlfVwKRx
3whruDSBT53FzuQI/AzpVBHiIyXL1C0yb68GzT9PLXA3GURdsNtNPqvYQ0dMPcvF
dhFGxR9ajMv51lo7JE1gtOkUGt/wTnuhWT4IkD1j7tvh3T8MZvyUG/sPexqA8C58
DGZvo8xb3km42SAHHB1MOyHoGhbDicbogn5EceL7GJljRUaQJYqvjYQHV4VQWSRD
vZj5c2Fx/30XmxhVo8gAICpV+voK9fmACTAv12Gt56+MGP57CcI3Wlt+8eBHsWcF
mgNNGUwpMXmZTfbGtb5fLUH6QOwzVYvYdjBY5XzKqSl3SUCYateNapeTB0f5N1Cy
+obvkkjaz9nGYgT9KajFovnoIqTX/ujWGqo5dKe1djJ3WJ0aOjVVxFVHLYL/23x9
ZzhPNUxJcQemGnEDAkIWqn7ppDnnymqZtK3ifRe0xH1YYqntLngh00pzf6NWjN91
YDdhsRST3QDyN6WDcjoZl7IJc/FNkjiBHipnUbOZCcb6/1i0GtdZyu2PVwGknqvW
aXxoUszxjwuCgcLNYNGuvnXZAhm7PilHp+F02euh+7Q5NHtxDIw1NuPAB6pVC5dp
NE8Mv3/LtonRRy7ufYro3Jth8fBxbvyD9Dfli5JHfLTYivyH8a8eCOM7UXJUkfGK
CpWWIcfb1x5VJdwTBwSJJaKErG6Glbl1XKToVYiH+tmKQL7dJEI1+gIfnjZrOAOt
5K7mO07FYYr2LOTrKJ+V58BgBdbvS9HQuO+XaQCdrMaMArP7fWDj5eDKUKysmegy
pI1xhs9gt9No2fkfeQELcP1173waNEq9wxNi+63U33N+oN2cnFOCyBXmaRoXYued
zt5Aj6eol3AxZKnqysSIZ/Q0shydXymNu6LMyIcvvzekmMWwuAg1fzucJs8yT+VM
Kddntk5enwPsyKPkr0/WmkcL9q8UYJJ4KGKAb+MwE64E8ROBDwK+P7AL/nUkC8K4
03ey2681X13abMDaXZq+LHfgUu05e8RO4TvVmSFeIb5IC6xxkX8e+ghM92yZeC6g
t3YXMdscMpOJYpRgx37JckNF3lomyKq8KE1bOlOn95/AXcwS+UdpSfLDp6onYzhJ
PK+NibgcegJvltiN+dw/aAhMACC9XGA2H5L+8kvHEozuA3DjbhbLiz1QObM/uOXL
3vqKTQJSuVdEtO5PiDoBWktvg+KTc0Cp3ee4FTv4yWWKvhfHTXjJ5TMNH/V/Puy4
PtJVfKQcDRqSF/+HQtHY2SmM+oPSueA6hVToeqOLMA59RcMBec1bD/9RKBtC49fo
aNKLSWNeSh6KEbwBl+3ifAuEmXBvzzdQcBIFVBK8JdBtNEsrfZrYgFdgftbgWWUH
py//TPcrDjMSbF8i8YKoVzjGJrhVYwu8V+/rC74aIa+KDXazP944HVxSx3s2CxrJ
4oqFzo9838k4TbaOyvJQk24NIPGa4R/Il9MdNYsiYXazBRe3QBUbSBqY8mEyfHSf
qiXl47RCTjwYTluxso+CxcIXVFX2KDVA5EXdawS3ltDv+0DkuS3xLke8yauGBuGo
2fMsQ7aHImWd7/xaJ0sESCnuagsCc7hthpX6IQ8LONS4XG1rLLjTxnx4YQjuZxcU
JbLjcv1W/lB3s54MxoOKbqIzTZdpRlIzvghsYplxlvVergzgt89sqZFAPU7/NcM1
FmQi2CUd5TYV/hgfOZZ696I+rixR51muKnKXqyR0vOat/ltDiLzUqqtJ+vmzNsGO
lnf2CF90/jabL5XqMbvw0AtgEHeEq6ih8ZnEYvm63m3RzIh2vnP/QLYxIi/sn38x
idsXMUXhdmKmdD/Qs3INbEQdbUFVPtf9GMe3irpMxZIzxJUx82cdnXpkKaLqL8Yj
lmPPZR187o4ATNXMOquDQztr5e/PCO029LXMFIHRngmmQENecMKa4NTkYB5oI5kU
+5+72VRpi8OrVW88d4wasUgili9iUlF1v21Jryt6MCtClfLppzkow9W59cGvt1R3
w/c5T4GSxzw+jHjW4JQqI6qtnDLMGc/UxDuGASbYbORrZR9/l+1bQ/Eni6lksui5
20DjceqUIL7Q9kB5wAMJmg25EVPN2pirLKdWhx7EA9RzPYoX7eeo3C2dWPD5ZTbv
Fcak+2vn6JCGSQHCj1wEEYNbvhgalIkj0FMQtAV4ZOGCDukjLMBNqVcU37CXbZ/S
ETiWljxI+B5gY/fpTHQdU56jJR1LlSUr/J5Ku/106QVHfHiN3PIGL6lbwRV9UurY
PqtdGEmopeJ+PJ8dER02ZP5W4upt1Vzo0B0RuXvheMolzCCLuGz+8Fjs140Y1AqU
UAzxYZGYwfJ0DNLq1NU4xrTwTFgTgmDQoLaulMZ0k4OKGIa2No5nu71AFRstWZ43
WqmvVxeK41Te7Esm5tg8Fhrv0U41OqbNTdDV09YkV5ccAg+4QrP4GyNhPr25qt0J
7VGqEZgxUOC9ztHF61Dh8UpySX+KCoGyNtfylabarHvOoOBhzjn2H4M3eHlHdDrn
FlZDcx6C9D6ovjr0e4OCr7WDoKKfKbIz+ugLa73uQ6NKjh3LdyIcCAXkrCIyNdEQ
9ualElRluTrkgzxxAf8oCEYAJnk2b7mstjcXhdbFCaLYobhfYnY+rCGMIvWvjQre
y9REbhISG+BF6nHb38tgKnD/KIm1xnmcD/cLF1YFRegmAjJMiFSv/QiyslE66Q9B
OC0mcoN2SaUNr17vGgeLeka3s3UBr9B5TJB9/Hv6wz/w4erfuitTtfHSFD1E95nU
FnSAUdCET/K3481OhpPT/5aftSzACHYNzrJUP4GrUWZRGQfSWznxH5DBT3QYv0i0
yI1AOVBpLLFy3ZE2g8fLf/7T3S8bjcu1jf9HsS2FLNKE3GthvHtKDpE54Zb4R96B
+/eyFYS0u/VsZS+LiwfVzyB7lDL0Bfh8sslZFEma96ZmvkltXzDwXwvJBnCBVABu
zpY+IKRVuItLBYLXWr+yYn95nK7KWk+GEoeXg/YbZF2iq4q5iapRKp6R4FsgsC9R
j6OzYidK/TcoyRhBbJ6pT5FpU3p0pILhtfJ8k1qNsJfrYNxceKAyqtYm/aVdNyxZ
8Oh2ZXshdHxzi7jNjzc+jA2Y9x5zw3aWDkAJO9HJbPetbMIdGTC3i/HxAX4XoizS
0vb/U/gD6L5ug6U/sZLi5kXd9kvSu/J2M2iVZfFtYv6dJa47CQufPEhTcyOxBUO2
MvDR3CzRovh6nCu3AwSyA6Z0QRuj0qbQNqyGFKH/+OL9TgCF8JygpgihXbjDGXGy
GAebfTvglrHFEYboBv+p+EeApfeYbDImQDK640srQaDyaWriyJASv3BkzH7WBUTj
4QQc961QMd6ZVghzmc/VV2o1ooIfW6MbKUFe0wezlbv8YXN4LqE3tAK3T8pJqCaM
7LEDwwHtAuDQWWzuEquffvoTbPqxIyDjCnm2QQwVbpvhSyN/MmZ2Cr4+5SOU+Eeo
I8fkDkuc/DYUSLXkxQoj4YUHSV1exniamChf20RYEj4c5304nCMWpAJ2Jt5r13Un
2CmoVUbVSGSfL2xIg0MOK+YU42QXhUxwx1xSLmRSGwpwK+im3tTskn6biVVFYNOb
leGp0+0vVfktiLly6aIl/IJQdSS0QK9A7USZTFCTWhadNAevoGTDr00MklRF8FV3
gbC3pWqeedGP/wERe1dnnL4y7skpTTArryBXRj0f8VKIy12pmxDJZe2igb8hUtp9
OVOvCkyOwNmE3vRyPmTUXcmnVpEqIubO71GCr7dcJT9zNCe7yvyLQm9uJcRcM/yJ
VUd6Vshysi08Nup9pHtmD/6Wo02hcSuR1hicZqlIxqWlmYD4aX5WO0GIYhnLnY3m
PXfRkgKcFOJ8FKV29xmGQ/F2IsbAUjJt9yfeT/zefLelThHVwNQ3XsQ4Vnu6ijDN
v4SRoL/gflmyAi3BGVe91zbiNuwf9VP20jbz0kx6Td30Wf7fMmfhFbD/yoZaxDi4
sd+mDyUjt0Pp+RD8RQlCIaM1eF3qcGI5TK0LBDZZcG3tpXPouF/+YG02/qF20JHF
4r8qJQ4OEhwd6AUel+FHVtY5AXLhi3ZAGLSCqLwrNd3dzmYwlTE/+1P2Qcag5prF
lj8JhP+N4u1hYxNL52+Pm2/KbVaJ36S2HFNh0xqzGE1ya5Xk5lzFceACH1CaVscg
A0B38rGTFULVQYKyINonynF75kLu9YCdQc+DhXIQn7FRifntKAy9/1BuHvXA7c32
bw5Op907mX/1rECzj8K7sr2qOMCyw3LOdhlqDXEcfxAKJTHKz3YdxDPUdQQ+jGuv
IBGuGkvyPZhHQ8dgMUlUpgT36+9mdLXMaqPT5KsjbSb2ZU+JpTCQtbrpBOCUh5xC
YdZlYg5ciE5mOjo9qgxkgDKozvKevRJljUMB/d5qTb5zYQ2XabXT/X8+jJjU5e14
xJ58Yg4XIPJy7sjBGrlsQbYPGOMUj9XfzT76oBON+FIS3vTYm5tFjQTJQ5pgUolf
qi/CL9CnHFgJn2/I7lfA7niGHXr7DbbXngszEbq7+dS2JiK193myarwnJHLsP5nJ
MOhZFsUYUa+ni7+KX+3ruXZ4FXFZ4EyJf3QPMclneDiWdAfbQt3wocxCtp1/mNg+
qN6uGebVk+yXeBINojYW1yIBLDfZ60HtY7FIxvVyFjKBQpe3yDzJzOT6VoGdn15S
ADHhLmOr49jAwJ2q5Er2Fz5z+3GKoEmjPPLJwN1YfPAR5esUgibGPv6NYiFj5wU1
P+zzoBMp9Fm9f2Y2uXb35FFkmT2C9aI+IOOUfBWTV20lsX4V+bdo9v7COqX/DUY6
nRXSwXdgEKaICfv9MILI2WAnCvpJUjRKCmO4zZk/I6xYJoTi2/revGZjqqDu+Xus
InOGwh/wAXKFG3ejrWSapgqs7nbGqak7j6Bsu12x7pFjUvSx7kLT+Yrn2l4/QmSP
kyDPIRh4MNA3BmRxkZB6iHwwdfVXAfGdmOSmuO/zi7n5zHIDHzoHdZwwJ16xJ6AE
MNplENKePxG0swU6F2ooEEntAfG+KP3D63bReFSyKcyPLUbvtpv/AI1MeKnV3qNs
GgoarVW3QzWL7EEgX5+dfdbj083Vgp7v8aoJEIJED0MePVImhUMdYGUDWmZZG4xm
F67Mh665DmIXpCs77AfnWzyKb+doKCq1e1oSHHMcmHDy8y/TgxAHnwYGgKnwVKv2
sW4n1Gke1TdM/eVh26AIBaw9VMcNbbxfKKO0TpTKnYWWLY7bk8D/EHuxo1fxJfVv
mh4oE2dKJ880ri4VZ9zfRLtfieEigqM8NoOqooNN0j5T60TMk8QPUKkUivFxOHrP
HkHc/rxRoRiPFCt72kG+N9I1xUtQ1bGNYFw7pL6v5GsiBRytT0EkSheK4QqU0h3d
WS8Hwz7vIprZke3vvyvbaUzNmLXmqUshPooMQ/0snk/tGijxfT4gKcwpdX3+ukyV
ui5hFb6F3+EzvzyhZG50Hkw0dYF4JiUu5fCdJuwoQOahzpqQAeGfb0ULQCVgSV6v
BeLAkJxN8RcqaCbzwrzRqIrFWcLjUoDjKRVX1cXzwk+JS5fE3NkyfrnUUUXYvC1N
+wNxkEaHlgcn2qJLOOcXwUwzrsx5ny8xELmh+sqxIkOgvceSEB9+FTnUmvlwNShO
XGHbh116zUOGUssiwfaqjA/IwoysZxdjHMJL7xC7rsYYGVZTIVSYmYmRb2V4vY9A
J3hqfH1dvuUEZUbtLe50qFENf5yZdQlcfsPYGdzke4RrVep6+xYpU2/Y0TlrjeN3
FmlPm7VCVouJMgYAH+2c/YgWhuWv7i736gJIo5tuWpBfbfdA0uRtJZJkWJzehiZU
Y1qfLGvrrR1EzkI8MrsG1MWAyK/wewf2PlqiqldyOxeNtulOXI45XiHsqggX5UFw
1jfXajuVT9DWn3qu3Jp0JdTPNx59PYrFhcrYGRh1WmxEDiQUyKRdAdUTUMm3/oji
8nipmiwaymG6H7cfviKtkJUDUTi5TxBQE4Z39rR49JOEFMQb2p+YY7QxGY7RISAJ
51mikWKoGx57uZ+QBAMwmN8K1O1ILxh11Ohsl5pd8xbxMVISHeoJIvDXw0ScmZCZ
W6mr+TVfrzwMxbijdwqdcVPe0sVyjbkyuZQmIo17eMpF9h5Idshc2J4pbhZDqA42
KJ8jLbIYThWr0UwgNHHu3X1smaNNFN4V6pvXBHHs6hsHzJ8hAleLSDmLH/rGB9EY
tOHbyhe5gYTYtcsVjVEY4mGHmZmis0tiypAEBvU2b/vmK15mNL8rshqe0l0ZvB1V
CO6QHSdZT38KGzEpC7VgwL5jj84Vq0uo30logbNBnSIjxVhk0RJRcn9LaIiDrGwB
gb0+MkGRfzYZRIBcP31/8FKSfaHwXxzd5+LF3YeMdFv/WnX+jRmlcAeDa2L0Nm7I
+ROdpOJzMFqMgSm082lB7oUmFMA0wjfXmk6H5r83vDINhcxdTObUIowlmvyhfHAL
Zzs3duFEzFMcruayppJiuV+dguM0XNklR+heUlYQRVq1UJ74E7wgS0Vk+c1qmMkR
0yar4YXksQfbaD5O9YKw5qsbPFGZp36yiJ8cxXrAXSTWzFomni8ITZ3+nLgRBvN9
rzJx5vl93yLDueSMYvi9AKxKT9r698lwmwxyIeCdI2NpexU1tJCLuPR3y2VGqeRw
PiSdTg0sRDzLMBDXjqOUiwlCN/CIruRQIOGabQFoSrHTF1ywA3QrYkPdoPOKYdyf
B7TX+kRh2uOyVSma+eF10Xkv/iPIJVtXl7GyR+WjMEQuCBMplkDq4R9mkQ8zh1te
KIgfjcYARFJIDr4tDDuzH4CigVk4BwqmP0gt3G8Y60k3tSQdabq97O3Heyo35saC
dlYsQPRW0oJHqLy1zKBHMS6CrrD82SidZsESk4MkKhd+Bba9F/DstkrgjGwlFnho
X4dnD7TD1dreEQvY5VDG62Z3DS5lZRlD1Y/2nmNdgkrDef5/etvuPQuGGTOHxgnI
IT3dg5VN0FXQWrgnkPOiBVUnEzg7Qx1M18/AE4H+1M7CmV5fd6Odd8vinopIf3wI
HzULZZw23XJjFQMx4FIWQVxF2iF0R4MX1mmlj09ZWhfNrTPZ3Jyd057wuocAe/nv
un+/xSlVarhULrEVXq+uph7zlIOAAwYShVzUrB6Gd//EQ+bUoNZITniFS3UNQ1Tx
Jq+BelLCajxNizhh3Rdokuq2iIBzCU90bQ0gqH5TdK7xvalyTTQcdjBpmFefMsMT
vd7OGjaHtiEeCuJt/PvPUNWAZ3djS0YGeizWMsFsnTWmurqAaB9WMXUeehKR5tij
VnBrKZ/2QGLq3y0EVvwm6+1dFahuCTdtK7HmNlKynICkUI3jaxGVMLScRfQjZpJ6
/zWQtC6lZJVJdiULFYgH7CpArZWhMs4WG8pr0DKZUECZ/8b4XhOMVdtyoJxvUJIn
rEHIBWCzDft6B/P+VltGDTj6Uv3Lv/qvuDjY89RKOrjCf/19ZIOyXzK4GtfxDqN1
ACUA+50xDjYrLvAFJvb2sqPDFqbJ2CLahgMSVMh5Wv4MPx1nbzq99ywsGBltNUoW
RGzh/albUZU5M4Ju6Av/oFYh3WKcCW7sDQz5A4AL88s/hm9iQourpnWbyxMqDp9G
lZxiDg1mEsa7nV6NXV2FgB8gviPLTjUsujuSDo4jzo4cl1oE45alyDoOT4/cU1vx
ooLXO9jl/NJyMYIxlmatTdiXNxb0O/jNP2uHFDPKLWsQMQZhNOWlUMhnA+QDeTqz
Tjcae977e8uOCMj2ZctiZTyVshlycB1nHtpQXwCgudcIU0SiB6BsNsnVLZxh0MYP
jNIlYDfkc06+Pp+PkiYRMNvax92K328oIjaCeSJtmwEgenzYuXTj/iolU1ipI6GT
z84Sg7naP16Ub/UWhlR7u1oB6CdoK9CuV2aDARbcLmWhcooXZ+dt609ZZeCN5Kyq
ntqQeymiNIJ9KR/rnpydj3gVgZyXqa6lFOLwLN2ccTC2irpGeG5Jk2PDxSWOhfLh
hs0oOICDm8De/S/ECkS97WOTJJSLeOCQuv6oSthkZz0n/Um1OzC+kxuNtPP+ecAB
lHdA/olSzr7zlAG8dru/rCFOpHg9dihZAPGQVTCCxzTeAOQ24EotH5BoZbbTUdo7
+1/C5LhnWvIE7XMFC86upSvq6C0Jc0qPasShVfKdr9OujrvuX4CaS74fGUpqpSrD
WI31IX7GJNHyQJkWQitbEee8DSOtMgc6YwhODOgDqv5HKlqrhNzjDCKfKKXUNC62
ZQeWqCG/Oe4y/dAL9TgfFQ3dUdJKNze0ElIxORpRX8afom/jFzm36feQt982bpbO
dRd+0if9duzj4I2TESpwRPqCTO0i68sE2q+e975H6xx4a40bfZy7g/fBhHLtU9Jw
5twkBwHqqbnNF2BwZ48AqxlIh6bCKKKeGfbJBYFPhHC6xm4ulIU5P8H77kKswzKW
cAxBy8Ww5O3mfIYX/BlIOMfDNfUlVGVx42MzwBX2gTlm6OLCYpYZiuIKUG7TDqb7
nsOe8YfENsjUWXcS6+LBLP3coQ115Pv/SqZeQBfI+7E0wSDaZ/LuI49/c3LqBBfe
rTEdw5vKDvAZR0hqHuUg9VpFYPy42kR9Kbdr98P1/M0XWHqgUrJQfrHrg3uwnviy
28hWd0kJZNmt6/Qrof1TMXzSWyMYaFtpmc5tMDyOx8mP6EsU+ntd9iFAw4DFBL0+
1QD6mH0w9IVqkYLAnlMBSfehK+vYANNmvzgRFJkVgpetOcYbWspkuvEKxj2lO3S9
S/nHdtKhuQcyMXy4isoB62VYZe28dBypiFEvxnr1+6i9stn3EWWoEU4x1i9zYaib
KKV8jfyEG1fMfKHKNfbKUTMnuQ7jwgdPhchS+9GyXvfIP9qviyK5Ur9ZuyDMcf7o
qm7AfwlkLcRt7UE7W8PANuwNSr6zTb1HepW+bKv55VC7LHwXB2HFmRbcHUueNvE8
Asc9fm0UwUSmjl7Ih1027Miy+WesWt7/wPks7H+yQ+ICAHg3H5eLnabc7Z8JqNHE
dP4F9QM+NBy4Yom5RvjaCUDu1CHrRyBdsje+Nm79V4Hrkk4pJOKZAk718spOlXiM
xx787nNZGUnzt24kdjM/MOC9xXa6+4lnrz0xIgEsmqgfVZKrVKYyaq37xQY+cNva
LavTelPI04JlF/vsiYlwTnSdPMJd6nNcpM2ooNAz98npqwb7aG2PWTFDQJ1CprTq
8zkb1rZYFDfYQZIJwMEpMEq+BrlGeNHbqAv/gjOT91jUYyUzlSC5tRQ+UDqNNLwS
zVBi2mivHDT/Z+ssiyGiRGto/kAiLyfKcZ+mlHJ6xWROT79+lGybkETPmThgc/ee
tnSbWYKGWJL3VGFVR0pgBZehpn89U8QXluTbzthKqPv0aAHoShG5u+5A97ByrYRA
xWjwvJXZ0CIqu+H2utCYiZd8+rpFi3jOfbkrqe3npoefz6Ood4+TV834yidYV4IZ
6bMO3iHf4/wL4qna7Y/EqQP4hivAh45i/rP2VjLFZf7OJIQtucXDe0bNqSYEvF0k
ZcZ7Gfqv7uUO93n91LAMexkvsd7uiI+GklcS0LafakJqoGtQ2na31oELV0GqKFgW
MT3y+Bpz2k2kN/Mihxsgw6KJ/2I2jX2YCvAD8rEWN7YisrU1+KVSVZLW66qyCtY5
NZM3I7S+/753nKD9nszRBbczdBSrQFqsEAK2BybjU3yzFD/lymsaVA8LRVjR8fLX
agL5IUu8OVzYg02IZ88F8rxEtvZA5TTQEx0ECEip0hjuU/eK9A7dDA36yIqmfaUC
toPfqt4JU/v8FnjRR2NyrddjxcunNdSOIeRgguDC7VIbwplDj8FJgYPHGwTZzOuD
0XlBoQeW07NcO0fqJWlF25l7LR9kdPB2h61+3sjODlFgxLI/WMDHMesIoiljuK8x
Tm8fYPZSJpWTdAoLaIOnozAOdwUYP0YAbmIv0GIdKBHygJ1tTNiG9ee5D1z7Hw1i
2n8ybgVnZejtPz3ar6ubNBgOzSu3GuMDGpG0Gqd33l5P/RaCH6VfbwpkRKUrq/5n
xbaHj+TvnD7fh52tifc06g265+Drr/V3rfkZAxoGOXxqqkg0SCUYyUScm8g8jBOY
xlCUEmjuyHMC3DRDEqHl1lcCq/l04WcRb3lny2eUwnKhZDmGAKN6R/cs55b7nyu2
khX7R9exOBPYJcnp7yGFhE4gtufY3yPyBrnHhrC/NSch7Kx6KMNVxh6caFs/f2fc
FS3iTRNw75vfgWENPYo2rbK+pZejQ688/Iec2YeDDcy6kDzAnz/PIejwDGkcp4aG
BeZqx03cy5qU/mSPsdmNB4pLgS2Xx6SSImIvV95r07IXu91T34BwgF7k7kDK3uJA
X+RXmuBem0NyIDtpL653CLB0azWGIaeHFTyEIiKkvV8RCYa5EHdXngLhQjJJzbkQ
uyHnPe/rUIJT0m1NUJH8qBaoQWaxZM/d4xnKNznhOGZMIKXMr9kVyNIPg+J2+UTg
NzezbBFx0CMj5m4tgutMMtqj9zlIDJExOVkx4Cdo3/lCW07Zw+6TFZDvjk3hCIpn
kbDowu5gUA/5GTO6ZR5/JEaU+TI158QMmZ8Ps7ppFdrAnn9BQ9vvf/9leVsLcz1O
InmN5mreovJOAZihT4bVs706d/o81uDPiXaJ2SPO/EUsCMtm2bpF05u3MYl8/bxZ
6N8BBNcvFRFLeSCKj1vLAZUWYXP+lOD+NliG3LpF4Vrk3r7QdK7grF5kbIOEXMDB
vmMZn0KdPmRgqUA+qAZR90AtVQnR2DIUWfGO8rTDmstAWhQ3avsftgc5dfvKTnq7
oXUk1RiJL8pwO/skzZxyKqj8HYP/o315f6IM+dGR7kj8BKfaxj2ZyJ2VTrj6fBKp
Lqu+TJy25im8/VAw3dUkNCyzfvFfJaH5M6VmsaG9LwfMSfO/D4cA4A9vXqhv8hU7
kAM1corb3uYnC7BXADiDHlzuScAn2nkd/fbA1Ss5+g8tJG0DZ5f8PFJvXTAWHr8d
GdsgO2+lOorN+P+MiufcEofCs8217iFTNSlI7vd7OqK/5hiQn/j1xXmSKKFHtNeQ
oumQwSH+OvlsNLiMdpblite2nbCPHutJK7txz31rlD5xIw52RiQLpyBCWahFC5DQ
jVppBLmFURgHTGEDSba5ZnIMEXVvCU1zWYjBikQT2K50em0Bp2vo6fXCe5VMlYHN
xzb6DsL/uxelE26CiMTsk5jF/yUbL0nuc4iFZTHrNnDziqTWl1h7y5jWgCuWcLEn
MeIey54htdGCbyLRCM8DrDJe8knP48iEs4QnYAH6pyVmXugdPGggpmyo/oKfXqdX
RBYhbLYbuuxFfRfCz+VdS6oV4iSPbI6d9Y8PoeCcrpQJhHoKduczP4entsI2rnBX
eajCKaynRCovKMHT/efbowoJFvNlKNxZ1e4pUDL4cxGspSU1FI5iJ0NSQNduOrtM
KCG++o/eOFZIkgh8iUNqsWy1jCgmR8liHidsrLhLEewzJ2Z1/z4+IGyMY9/t0rmj
WJ3hhMKdiAXxmPMv3Mq2LR7gJNvVDblHbajA6m8xFmmPGrqmvFIx6INmCxF2dj+f
1DNE7wgTKp1MJ6yXpNw6seMEMMl+b4qTf2yWPKkcc2yM5BYecol02xVRMkRLsP3V
py11vAkkbZhDa6GPVkvxckQml0+AfIlp1ywP1YLtQdfQnRGkGOSA5Kv6Cy9OH1ab
oss1gSolkgNL5i7P6uxnK2Q7AuXTfP0DORTPUsYWK5xNKdbC+qKuP+0OAgOO05dH
yBIpXKTuw4V1Q35SQrxKlUKYgNGgtzq9ZuCFQ1Fb/7g/rvCRkrkW+CO+vpD798jQ
dem1g9s5uWLFdlpY31A30xrBUY2gcv68II9Ye3Y3EAt4flmgqQCmmmZOU+sgxlUa
5Ujog5apx4KTZ5M03yQWA7ryFZAaecndqQnUCrG9bjU/ny/7CKSoP6M+o5CyxB4t
yFxXqBEWkMHv8bjR7JCBwc2NkG5KhoLZpdWkwho6TERt1Z8fufpkF6UgAuXRicRP
Vv6z1MepUXaMnIjGHm/6l0UJn4rL4c+5kvcDUP5c2IdUFt/K7BSnRqlfOY0ltN2f
ZJ4MPI7INc4cZ93NQzxEtIx65pkBtK5K8LM9Omux3tqB3ZsVwtF4vY72kLttdXp6
+wGqc1y5MSXYMZgUbwnRH3QDKGHWqJ53yFTf3UXp6h6f8ofcKIhS3gDlqnb8Hoxo
g8Vz8AAhhISVaE0LdjbT6+BKiN9wGCJH3dH536FuPKzFY65ZIc/UvsBxLbnQewGf
PybH4RHw7uzO4y6/USgdLHJXfGw750G1qu57hlTHnqaM8LBLkKOtHk9XAFfemxRP
E0HEXW0vL8WZjohXqqNSMoYkjYUYpFhBFF8A1Lfe6EX9iQEuWXteFCmrlxA8PmZ+
rqkTBQieBrpkFY2DQZD1abnNzT1NBhqGGrjo4wSKGj2PKBJH40ybbAmD69Z8h8J7
PIUHte4F4kxPepeWS3CYWFn6Axe17XjnrBBBqw9DZUu6zGuAVluMCclxMKUiPGR6
AM7S9zxHJ2yAqClsnAqMKot2JYZEMvKQ+87tiIS7Kd809TgDMW9CIJ+hGsTtd+Kj
l1vQoM6azYRXbP+OxbNNpCvmC6gASg1amlpSHryOZ9GrXsAGcE1Tv95sIcJwZtg1
ySI33g4vYWEAKTPh/hRmYTfbcTuAP/iqJVnNU36whmYnlyIKpHwXlHvDLzgzuQPO
Yy4fqA9BsSja7QhNAMyU3D7hP56V5dwFl3bfmMCtFWddQjtgezzLAiAwxiIna7QX
QOcqgIaRjUsoXnZkEciibYWiwE0UbOHk7Bb3yDDgYejcVxQ0XLW1wA3Jn9+Dlm96
SDTPURnyqAqz0R1HQuj1w0eD6z4f8QSJglGGifoQwkEMcEs6RUu56jEt0+GRytBr
7o7YDhF7mBGeIChaPaMmfztHrGKVUnHCHa6LuWU7oqyRDDHKTknFHock1ZlsSy/t
wfnFRIV9n6KajoejN6Um0ppOt0NfP8ndwI8KtJ8Ziflqj7JQjGgz/eZUBmG7MfqW
eBlf0YZpz/qBatfZ7U3XSxagCIvPoM4LcN4IZOrdjEGHDsqzHSeoipDFPOHYXJh/
uVgRL1U6aD5RNBsAwIBE166t1hSu2BvJeVhI0kUQyCCp+X214GDkZrMhXhTUO0B7
km4lqZZ5HJixoUAADuzrBpmnnV1visVDm/rjle4qfre1WZe6k42CHCYNYv+VN+T1
EZJ5xFVHSmMF+TuQPF0yJe6t6rw2XMsiWyxMp6wvrTGHgVeAGP2dBMsJ5asvfg+f
enm2Qeu5+phmDWXl9fCtlXni5yyCokHX3sh+bLopWvFAraMz9ubgkGANyNY4pM6g
X8QDIQePSYmfANuyA4vWrbyp4d8Ii6hVdTEh3qTm0wOWqaLnZxscqSozd5GRY7w8
M9+iA9fVjnykEHcZdSS11dQRLs98BNe54jZNoGr3URrXpExDtIlwavSZCVIpFFCv
PXYvk4OUHqPlLU3up236L8ZY+EJnbZBkRzzgCFaCv0Ob6yfMbECLEHfdnz8lLPfB
c55t2PheOQejOEG2W6H9sxZopv+h8BLt5B5j+kITD8iZypEue2F27gsu6YC89xOY
ildnZYtDiOmkw0TSO+/LeU3SPdXO97+OtPin/3g63svA/YkwFlI+Lwp6oxD9y7EY
y1wqGyR20NjKYI9C+lMHt4TVRLDZb/XNm5M4E6SLReJrYyFUG70jY6y+SFagCXp4
RLnRullQmq6jdC1T9z7dCSArgGFoTL5hTuAIJIEItW8p4SXUNzPrXFO+00mgEvKh
7jYk9+INQrxqvAmYkxIdqaZi/pADKLUlGJ48NnTHMQp5YkNX2Gjt+ff8BUJpFKN9
nxhcmVw6g1i+kS7qEG1k8g4jmeGmLjw5jjc7auDEXu0PiwVvnHVXdb8wTdEDT5M/
eNO+qHaT3CU+kTQIimzine292OgRUfUfENJM344WQS8RH0JSMYp06DVIVDR2KuKy
F/JaqkDvVao4FbU4J+hbHELmddHz4QwCF/E1FaWq+UC3byYDuO14f/+aPs9g/Qzn
8IVgHpeA0OU00H8jTBvbGkHm5vK01BOzDB9BabwXlKHjbay1MEwXywstg+Cn7eS9
VTwhYXkkpuxKmyVduzMWqoVM4ZTmt5/JGYBMmxRZ40E3L0PVzSxzAdDjX/6yD5SQ
5CdjpTex4oh6E9fJ6OGZU413uMVMTKHTLzsiKH1KrAuxH0hOCZOHlEon764Xsm6p
z4yIeTekBeq/3EiqKGoFIJB8vSu08XSkJSAqhxMqHtGvasfvy1g4zrNss+hcmRqt
D+qPf5SBLIfB6ioqbG2cwMygMPz44wBusKx84A3Lu8LRoFlMxcDw3uKW/sYsvHlO
52uijFKBSwI9mmx/UF1vbInGO7/zzy2iO/kyV2HCHSopumA7t7GcsQ+UE2PiG3gf
Hu6q3cXbNLjCy86Cyt1EPYMyo3QIq559ctsOTMkQbGIWqqp4fij6o7CD8Jnr+n81
xPBBkj83ivzXq9cGUxFhZ86DVZIIQmB7EPT1gwfTNBpaHUwDmc4Tj/UwgUtBFC0o
KinTMDQPhPaXQk9UwxHzsljun+WklptEU2/XNT0w4EHYUpxLWCo/Ge+5cvWG9xYg
5BzjsuMikvhACJ8GWE/ysBMkjer3zURUDoyo0tU1n4QnEBk9DegE4StLjBXhPjSL
KVIeuLJncaXnt4wZmGxQIzkQm0Vzab4Z0ND9q0wlqL8OyvjAwoAmNmNcRHz1Vn9U
1WwtxN5HWOhh8uaxDe43GyLjqcafbG46+3dcsn4gCeCgU8AqyavCjExb4SAgVXBd
wlNJbjYCipU7gDBsOubhxA6fUnttjvfYUcf4oIAPxNuh2hidPWRcCoY9BtovLJnB
z+l4eD2LyN0DCbMFqRXL/6dtuqE8E6JEcW9JYWa+PY3J+eeXk0Cb0f3pYF4wib2e
JHBvJFGB2clD6gTWqLcmmK0V1iNK9pC4/3YdzK9rjWW/3zF65cA801/aES+Tb2pv
+VwAf5ldjGJPbBHLepMXhNQSiExFhtaeM/RFHvGMzCIEdJu06eCzuuLjrxDWnHdn
GJE9iRInMf9Gw8lsq0tfeUnREaU/rs/AT0/x/jVPljo50BbQUjxpM6KN9bvBcwME
c0K3wPWIrv/X/T1Iozlokbt929GeCpv02MSk9WzwsY4wdmjYNbNeozKjKumZVsbl
2aMtxlhej7+CcN5IkjdNPowB4AXYt7LAj2I2E8aOK+zZOj//iS+I3qSRt/fAMqSN
yE8XBdFgvKYWn+R6z00PfUAS5hGbXhFGcjY6i7PDgaHdRkGJJ3bh2J8O39OfwJ/f
72DeZBd1P6VjQl6vYmwkkw==
`protect end_protected