`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 55056 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
ZIICkMu+S2rq/yOQyqhpug8TF1FzA/6MIyuD+HgFeWiwyfvSpxWuUhzae225f3TY
Ivk/vYsS63LQ6tro5j7+8XjKK/s560je1wJQ+aGKp7OpbbyaBELnOBlwB5NBIJvA
S14sqq557Ezcv6e8ceDc77qtZU0m6zsQU2pj4TMn9xf8PZL2T/iYUqnzp1nkbiQX
S5NUqAsA8nZ/oMemgcNDIGQL6iOKX84f67kAYOMETsHelCind6JkNcYWO6U1LwSc
MPRHX9enipT9Eg6yptgd3I4jjI0ielNVMJt/SrgtfZPMwqHtsXx4SXZGur/wNbw6
3pLJFnoCBVpO9C4aQaFIZobAZ06XQeQogHd6d3kICAfcAqmbkAoeEnaz5NtV5O8q
97ZwQ//q3sudvyYnjYXqenG8WYPQSNlbkaFmqdJnYaG2cPBt/uWQqHyjkpD0Ltjf
ttgVRILGmwSygRJ65re6V1V7CQUh4wN1xX78ygYE9K+tUub8Bi49Luaw921XEgs+
wUJYVWqrvpZKuG0Bdv9waVZV2q9JKhWkzC5mwfNMD4mseik/KTjsM9fOuozo+/FU
uv6t8z/xLLBkRZaUIUNv7DItmef39dB+kFHyqXP9+nwZQTbVpLaoq8fMDppgvzbB
Wqv4I1eKS0pxSpEBfEaW6OBzRQo5yLjiTMORJv55XMJJA0pQ/wLRSgTdQA/dMxvD
uR2dOfnrU4jNa49yPEh5XdO06B+udFWej3NsgkLL2RSYdHjaT94Zudr54oXNhi1F
KfxVzIAuKqgR4eeoeEfFp2IDNazkQlYoG0lhjwHPS26E4ElcSqiIrtMoFRyFbEMC
j295W4WnjPaeG0/6tQxqoGia9BHahLjxkT/3sb++PXeiAzaTiEJ/iifg3SrpQns/
q95hNncwYOX3i39r5XLQTT+Kvb0MzoCangT5nuGScDyIkG4Z2CJms6TAgCYmim+Z
Lxzl/4EnXqKoFaVWA5Y9Q62GFLBq4lJcAb5uKLaUO95iFJgEwUwXSgSsZGBZiPDh
VF0KLi1DVudpw1ZQZXvmCx7okwaSZlHaEtmFIyrGd0uLxUUsyBYlZuBhpfXJyeDQ
rX55/FIybTyu6iIr3l2ki/A/YmZxjOR/RbGSLUD7Qk+dG7wlwd/LPvJ4cJMmuwyi
lyfjQ0QbjAK0saMO1FLcUJbon3IRYiciP7FV54KPH50HORhc3N/Om01m8WEy7tCb
WVXWZtVxqI7yRv3e66Tz1xGMWJahh2tt5a69KTqZsKGeMVumLNVKEzzymQRolpaz
KIZVeysYMhFHo+0fujSvx1tZ12xzLHOArAnC5th9H77oDAsYr01GwJMNfvu7Hbjb
2KrWVTM0Fi/E2u4pgOKiuMK1atqzHirODSH1TpSe/RRhDTgNcElMie3QmpAVx4aK
ajy9XDEniBkC/CnXF/ZBXxFnilL2xdGnsnyWmTg7fBU2aZUEp9D/tlKE/rSg1bZO
IZgrP8c3DszHnAQn07zHt2XjuTMepfrea5DHx+Z7I4uRKfLq0BeQbGVYEgIJTNF0
JXPDzh94ldtrTYNV3C6cpEiGljwtZ2y6zi5lShyv/ke5DyfQxUSvz9VUgVwWNOte
BuhyFhAPPXnByb6z4ih73QyeqF5b8IyoEtPqDGP8QToLdBq/ZWYFxKDRn/nEtfAe
ny/+rJeA84J5LB78h99KMNHLlr2o7ORMxh1tCXo3nVqvxkeHXRUnYeI9+90m0iCZ
c4PbQBQP/NwkeBV5D7djd4eQ/pBtiynUBWxrzm+ZLOXirMM6Fups2ADM5Mqz95lP
OJz0U+0qRlpe/6wSCGKR5z300/TDf99iu2hMvO+RLdA3x+ac11+WDqJn4kL8E8Cf
3GPtuYY2WvPCKZYifL4IA3XYW6rii8iTz+TcR36N474VZmjet/DwBfS0dF3dC9LI
iXcIBhdtzIi9+pAWqXmmTFdy8k/Q3Jgcg3+DSYY9M5b00FoBy02Rhb0VBpI+wQjU
KGQdvbQ3ZebfAfZBifRewO7I6KjEun2rCqVgcz8CuEqD3M7re9019EdfeMKBQEQR
KqLmP1OQ0t6opz3yQRG/jjHUhEbUAUPASuQBpNQf/z3rZDBaq6jMnf8OHf3+X2jw
d5y40Q6wLR/LZZj5ICkBLqWRUx7C0D82Xde1rnma6AMcugqVh91FiHwjsqF5ibKZ
vqoKAkgCUyWdrWzP/A34PB+LKpD1Ty6wN6KyG5EwutRO9RqfGUukaom3nxC/btt1
PF9i/Rhgo+ZM4E27d7ZU9N/Kwz+L05XbsJTW5oXXi0DczpMr4vhUDgvK9NgfN6qM
5OnTMM3mbCCw5i4cs6Kf+JKZLJBwVI9vY2s5be4GpF+Yv2dR/ULyC5rowI1qtk8f
B+21f/q3N5dL0LnFpYv5Z1Fw+sZ1WUMppMHJnElb+vy6q4HiBdPFVtpJUlC7qDGg
ba6Id6neEZ8hiPbLNJqIw8u30WM5DeHHZYIARVqO5h8+IH2b4qE77wPWKGIOLEZY
yK1J0cx2qCd6i3Zv3OJb7xFNPv52jerwu4XCR+mN64mj3PlR9eGEIA6ud2ceg4WH
+0Qrb7tjngPfgx4mTJsJp4jLgcFfQs5Q+8Ol99uwVB0BWqVTRiEoG0TQfRVkGSDm
fD7iCjoL0ePGTSOXdhlH0GoM2aNfRnI0+DUGdq7pdlZ95oEzq2nIjDa3sk41UqXR
EZzjF86O93K/mAGU6PNXHuIRZBRWppnhjl04Skwt2rNSHUScEjFYSN40JnY0apet
F5UbEt72Y77f5mZOU9O7MkW3G+qbOUiRsHsUkZ2ucyFF+VT0ZApa+0wLlMXVGNlQ
m992PZqipLx+TpY2Iplg+EHKMX+Ykvw73OrQuYB7MBYmaLttyhkiuHEapDfwjqlm
yUNq5FVgh3NxQ7gmLijqwii6qd8x2K+ZWJTzid+0YWUR+BXjTWQbA1Vs4pHQi8K9
U4LJEgFXWWVm7S/JGVdL3UL7LuRFfqHwGpvWNDa85JVkYkAYgFLdGiBGfBCm2+Y2
lBk5U3xh8LNhbuPMHsNVvKGG59+TYJX/3c1QBiuIYCRuEpExu05/Eg4xAexxpO3F
NvJ3l1zaKeSRYsAO8efPZ5VuQ3x/GI2a0E80XCdXuQPA4jy+De12HiQNDUzlPEPb
quD9DCYoFBJpxw5Xy8Dq7iCE5fwpi2OB50VhYzP+T3dHkA5TIJkp7YEKIfmqKKqs
dOEYG9iI5JJ90Eel2BrgTGJHKpjoRCw8g4TWghA0KI2szha8GzgPruDBtkIrC7FE
RLK9R5bXGzWSjQbt7wcUCxa1WzoAtNH3PHSJn1+NUbDBHiIAHKmlIcjBMCMa8k5e
cEN0IP3EBUO+aETu2F9sRQZFHeLA2KnSXGrx0LNII+b6efQ0gxlUX8erknJpfQkv
ehpz9qeHTkSbgykzUqG/pNlDhbC8IAUm9+nO/4ij/ndjniPXQC5Mq8GsNsHaV0p0
+oZnT+B+reS+CWVl02vz8uhgJGT52rx4klZqfRXH4iGeiKQWaAXtZPDqcRL9YUju
Ldrm92+qogkwDuQq5suEoJxQ78U57DryIruUFH1lGMf+wqDgjo+OYXh2ZMbr3lLg
RsJbeeZYdmmCSfTU2pPVEzuePRBBg1HrkmezK7lpMZj+PW7yLpRGxDvdfzERpkLE
l6bKXCQRi8bgxMMan6LuUIwRwVNkQVouuek+j43TfHn4BfEyWJqw1kkK/ulCGJoI
DmUadilb0stUYDkcqJdSb5+x9Xi1IPo6gD+eTN1qx1R+ATWvcpKS7EBhMxJu5Qnv
6pl4+f4eWZEyDfPENq0X1Jr8Fn/6vp4sEDrw4Qd/Yp2NT1hKPaazWBwBifycYnVm
Sr2GV/Pvff6YWe5PdYMDCL93mUz6fi9XPGrVfwJ7FqzpR7FRg7lUBuD5r5fnycJK
H3PrQQktVTAGBo1goKh9pvRmhJHRNr6sOQm8gHl+D5VUC015bzPFdhPnHfQ3ZTuK
U4ZqzIXZ8VhTDvdKiVQFylgiTAJ8vm7ldHVxFqyq1V/UGVVsjfWjqY5NClG7aq9n
yMXgndoKrdo2VVCBNd4m8GjJ0vfqTiWHb4WJmNNTJTMDr/gtmCUDOMcEozGCcgYQ
NHwVzhvA37iRSwx/BOmNN/Ds07NF/V6G7qgNCV+BcRB96cszVjJWODqxtHjD3NaV
oTylIjcSYYP0McyzcLHfoFj1lV6jHxD3mMkJ9NM11EcVx+5hdlCi7ouDFLs9K+mM
0NqMurHcsc37K/RFxPVZw82XKKi6OwG0OiLPwZgkDLkB9HQGSFdzcTCnLxQHNBKU
RqRVmORQ4srUN7Krmno50ZV9qrDwontM+oD7m3zSt2smlpgXUYVlhdTLzMhoO59S
hZXVwzznz6MsVx4PCye4lSk5gyJiuLdva26R+gfNic+98rifl6Ig0OUdp98kCiPa
/ECtVhL+N18ngWeqTLs02QbMkukb/nJgXkmirvfuScFSXHn+1zyTQ8KC0p8BvKJW
oNmrkmgvRYZtCGxuf/MZ4G0d6WdDfJQzzH20fMJMoJq0Kd4Favb6pYpPljcad7Mb
xkSkbv1lC/BPV34JnMzG6/cZbv0o5buzYfaQifA9FZ+HgXRE0EiW0NeOMSSU0Qwt
wWYMIA/RHSaH2rJnL5Yc0onscQ4yYYzwOdhR5A0Qw/IhUHuRMEqDj7I+Scc+IBF+
3g8ikdiPheez7ezcyjgw77BkK7J7H8DJGhAVym+fCGvCNSQiGDOvfkatQzVrgoB+
thQNUDba718rnzuDr2fp6AhTusdp1nKqxvfyK+8nlYYhzGzl69eVNjz/Y5hV+tng
nBdQsKCqcMidk2DFGmOqCAJoFoajCCSeK9dUadl6zUTuzGMPPoUtLvZ3DtQK3EPn
BfYNBjF/zO+GYjgbvS6tK/BI0PwRZXFQoXtvhLW94vUTyukkHiB43D0YKdWOFGr7
I1E1xQEtjysMDZRnttT8RR89ymQxxhoO6NBeWI7yuRCrP+nxonQdVgK7GPc3R6K6
YQb1Sf5BwdGqMB9e8pxbGaWOIBuirps5BKOJUUQorWeXKoxN4MgossX7P7ObqKWK
sJCXF0gBqhxD+xfv9nbueAeg9smCRx6/25KUVneg6uvi/l3u/s6SDmqnoAPsLMO3
o2fsZVPMgcVzokQsqJ2hJQzU6R6h8OodnB2A3ixR5RC8uMJXe7Rt4KqqARQHlNpt
BfSqhgwLYDEUzvvDteZ++ZENAA+HiM62Sx8/L2jy6B5mB1sl1l5P509W4EPeq50Z
21uYTD7kZ6h5JNdXb+E2LB7EGIoXdKlPz0456o3HyFmOrqDRnDsuVWKc3gMMgoAJ
ug05vlUUGDchG8sM50zfZTRooOgNeiqcHLy3zoRMffWaYjSQbYAWI36m0/smWFSh
DpIq7E8X9DSGW8MhXY9pjnJehkLTJy4jRDljbekT+eBko0Z7FwFt6aB5UmITsP3j
KPI2Ml2gCcw67Xbad+uqdI69cL8R8xolonzh42t7NADHv9m0rtfMBd9S8/ypbaN2
ZU/eCo4ng+y1rbbmqiSM0ZicZE1GYT1ft50Zqs9dbidb6Ip5B0Z2d9VTsB2Mi+tf
Etnr4mkFEnpc7CjGR2u/7A0J6/+Ov8O/LYFsdFH/fVKthJ+VQ3udJ351CN23CkQ7
IHgVF1URqC6fqHCUF5C37q0e93Cq1V4SFLi1jiMIbDwELbpArcuK/tkd+mCuU0BV
xN6iHjO0DDJesLQCkXYPD0h/IPBvhK/weB1YGdfcmJFPDpiaUuJRB+bPgNFTpXCg
9aWDE0tAWDSUXilZSESPDq7NP9+3DZxID65EIZeOX2L/2OHyKjO0K/1W2t5B8Gdd
OmdwMcpJmNBIyJ2ptilVKTuchPScpZUU1Dtx9Hdj7GwqR7EK0h0K16jCJW37lCms
/fzowdijDDzD76l01GYJo0mk0zZVLQXe7ZwtxU4b80ruP2Wkhhe+I1XB8ClaGyYw
k2aC2hFRAEeNUIYx/Fqv+cMdOeb5yrSmbuezjc0ARPN5SHKG6lXpgliqyeUtmG2J
T9012JYn8GwJVMIXSCySWLA5PX2bJYtjIHNG8zgQ60DGxkSzWHFCRE2PHYR+Ivaj
PKFAr91VA2Wx/b5wyBzfz2x8YZvHuJ1juVT+IhFpiSHnmzoSOfqnnlclgVZ9haCT
PYj9ws/Rv8ctjSfgDYO97C4mjHxhZTv51sbzLqPa/WLLnKPk+yCWLP3faYyUleYo
zpsW5Zpefx6eH0P8C8VSwIkdyxZ7t1ahbCDhZ7XkEELN5M41UerBDCKcw0QWvw1e
/fyN6XW82BgA28//+MDd6bejpx/sTslESjU+mVCHiKcqdICigW0t+qL0JRXN8+TG
jRoBI+g0FLHgOgH0vfFaKsbhf9omkldeCYFIeEUPlAajkVebQaipqoRn8BUfl0cN
MUY+x54aNVRSv+gyZAdzcWy6HxlPU3vNcbPcIu4ym0h/6zHPpgWlfXUYZMcssZIi
SHpSAfylA2D45AEQ62OjOH1zJrMQmLkfluf9KBxVuf2xebEhH6yI/R2glcqevCjh
zY5OFaU9wWHc690txdNdVbdlTUPD1EpxdpXFHPQ8MqClcAnV1td3FpQFFXCR9RSx
TXTS8phxGynw1eXosD78nKk6l8oneoXFQ78m+o0eP/CBE2ZEuUiKE6+7ZsXYVqHB
bdAU7GTy87Gup5VjGCvV1ldAwWUdEBqZrdlqj3oyYjgms8rjMciQXgKnjjSJ1/vE
dDX0h7oUi/sqDdUwzethCSk7XweL+PkQnhan9hoP4DDvBBBUtJlHN2zy1ui9bu90
oMEoVY5ukyFeC+4IAvAwzK/lUJqvoGyMFD1+dfT6VXKP1YJpeMT7XmwpabyaG7Ds
LvBtQNsX3O3db40ydMhHRIogn7IvxXeyuf5/z03nXg5ePMkg7lDq+cvyi5k2QWhV
EYelBP/D+DTch9sjo/jvAV3ikPZ5XJDTI1ke8eD/fe/bag2tXYZl0A6YkkTzHSQ1
+VJhOuwGVullp2tMG4hIAkN7052191vJU0cY/eIGFCHi+15EB1itJYJorTxrvzYh
+0Bd7TbtUPzczvUDDp/d4p3LkHj39NL3zN7j/YTDCuV5OWZj47axDVtOlmohusgb
wB1hNQOlcCtMuo8O0CPGl/MiArdJTthV5ck00Z8OcK0MW9uQJA0psPe8IoEt7ngg
x9ws1QaYvkVDs+XwxRcbvnhHws+GUayr5ZcaDlUEkQiClkKpJDoV8V41PXRb089f
vfUgYChD3QkT61ToSM9OzBK+1zvto3L/WhJIiD15+MZI9eGJQ+/N6Nl8+r48dK/d
2lEG2xvrt7S9cVMCAU9x+uGT1WA5BIVreqEyf6Omme/jH4ywiYeSVG+KLLDgOwW1
P24K6dbKIgsOSyENXtMgE+sxGy3qvefp+f+Bnfn6J93n5gIPK7hNp4/R/3CZ/78G
cwGD3JuMixN+1rc9t6JtropzaY9ueQzNufAUXT920LCHzeQVbT8lURfDAfhInhmx
lg6TW6wLoxl+ASEzuf0u+PCd/WqTPf4vDgqhae5CaGgyzIgEqywHFEquW1wMpXxb
54KbLlfz0OpU9CQ/1WZJvf5iUv4rHnodAPrhZ61DhtEftwHbMwBfOoW1YG048A9n
vc1l9Gl4A6cdSXZv4DFQu5DcyCjHvHqttEN21aVgs9geiKPNHZdx0olKF3vDt2qJ
25XoYheiiGZ+a3Agofo9mjYK+NVKZ+Wbk0mqSNh7wcqKxlJHOONGTEH6yzw1JM77
he8seq2WPxr4IEABiGWxyhcFCoCHeEYAErAKukBJnLGsdOoojNm4pxYBxLSwUXqo
P4ko2g1n+oXt/uHrcqsPw72qtfSfmbDPYUn/g/s4WgbueYqddEXeCWCQCFe8Mt8n
cDuYasfrw7B4URlKexl3PlgkI8EgiV2WqVN3IUExtGJXj1ovIcToVh/AQlxd0qqO
L9vdRBFMn6txn+NXmi/QSTJ434LkQOKZL/ekeeZvFMUVtYsaaj+D+jGbvYp10CvM
XhufJxRCVkdnExki6wzAsEBX3EGSiOpZdWJtPo9hW+YD1LCeIaNxmksqNK3VM/S9
vQ26KlGIkSdB19Wglx+tUgUONqy3qtTSdsV1APVhA56CtRNkM5zoC2gENBYKJIB3
zZ+Dh7L3Jli2u8oQNmcwpcAMHU9ta3+7iqo2E1NUUDqUFcYOxohsz+/qveCYENsp
fhHp54CwF4L3OqA9HtcDUFfYdiLm6GGAdIimT4lxwq/OiohsHjC6iVcBOwLZ8u7P
pfz/qsld/L5qO9U9tU3LE6Gni+yEbibO2tvbjoksuczUhOifUjlmoz+I8eyCxmUN
vXIQKuTaWDQcl6Eyg5KD8LvqF7uv3Aicg1eA13dduwNG+qRnWi9c8lmE1SYso5Wo
0mLfBIf8TFHhOHuhStCJjBX8yZpm5xMSmVe/aNzUc2F39d56EH5y3QIophe7wu/y
L0FnqRnnGPDiH7Q8a9XDOoe5tK4j4QIORtI9Eeeglf36i2Gmv1UfEhu5xg3WZ99D
3F3NKaE6n7xMGkW3QnQFojaUYVGj8IYZqme+ExpauaoDfiSOIqYK0cKhJ77eeb4t
2JEZROx40OGywwRXuJwYr7ZynEETaMpZvNntrKK+MIRQ3vcDMSqSUwlcUt3hTgAD
2dRLXA6OmJyNXldxr3XNfClWd8vUIRCX3tI6lfP4noVbxrk5WfR5HXQ2gvWu83TF
MJKl6g4IJDR/hAW4Dr7paTnaqtsw6VM7qZFmTjo4I0secdeT3LskMh9G6bts2Gnc
GrVlr1SakXBSBEsF3tp3CcuYXJ9Tzu1T/MStHeGCyaMBSnNpNZYaaqKSx0MLTrxX
qytm/qRc8AY2JspsdpbWaAZ9u9oUHamV2qlnv6W8A9rc0TvtXhX0vgy/+bcyHCK5
GAbVI1n+CZ67fooKUEnAIuJqcIKBTHZWXOIjDmx8ICE02AmqKIdVvHPNWi+zhLHo
SoxVg5bDC/YIccMYorN2JHTMWeJwKUqb7kC2Kap6dEiixvlEN0kG8o2qbxhw67BD
crWb/RgFmdq5rKnA42pSvN4YIxCLjLljUL22GcJSVbcbYaIZMUvctKEOSIPsSTJb
WKTT9+y9C2Y3T27fImwV2JcMUC6DWp9LvFVW2RU//1RPYyazVhuMzjTQ8LYXgZpn
LWYBWypGuUhYeiWDdO+t1i6iajIFaoAlIMJMqVPFBJjU/asQZG1Ex7UpvTmvrmac
aFpCDFAoZhCt5T1sRw7XCuTCMNRWVRplE4paXAfmqewKpo3bIPnObkzjYBaCOrWZ
tucXOilJ3MCVQmzeeeJMjGCdCVTH2Oh2uXFzMwSEXf/LjlSzXFl8cXffGknQEUcE
+jz3BlpRi2XC2fRxIUBrAmXwFodjrlrXjWkqERKX1f6cyH03q7KOnKZa4B74OGyj
nB6fOPuHSbhv296MRSoL+5GJ9l5NRPVxu3MpbPU/nrXIkuGNczyE3BG7gI54ejb9
GBXHfiZEE0Ce2YsT+18YyHW0piU6VlJlSe8UpMeWszOv8SQGhfrMf/O0K3UfIufw
H5Vn8t1pfeor9d+5LRbcTz6bd+378OaJiF+I2EuNmvobQvBi2b7Nn2Z2lAZOpe/B
WpuJ14An/CK/Gt1CHFjuNIsfOVLCdU1bhQyaJa7HsvoZnGVfH9DBHUH1EgD2MTLS
n1GmxFfaRQMujWrvpd1jKgDrWGst1iLaU19fkrccM04+rNAA+Dupq7DUcjce0YeN
sKlRDDc2wjlQdgk5MSrOrv5ofjjzke6SPn+QeSJz+D/f9ZOsiSdMO4Stzp93OkD9
0GW2Kpgb30EJ7N+qR6Ju33jahvBUcehTIRhee2DE+o68zTk4T1BiiHQvmotMs/Us
XFpShUagEKyCLZRkRMed63Ahp0ZR0GN2oBK0pyn0Wg/t+OygCz8EVDJjj9Y98P64
1RcMfy5jPfvbJ+sxNFQg9E8zTsBjnTt/JPVc9wkb22KB1rzwpMtGn+pFLgcYmZh6
CYlckvUFmCDhDyuI5/HlGTsUjHEVII5aiB0rorH5++9vRkm5Cx31ABVyH0albBTr
qHszEPaA7VNdGYXFEbC0WcB7x8Sc7cqbaX2d9bU8gMQ/ZzsfsQI9tYzXmoXnptoj
L7LIp/8XlGsNNxcl5mX7nxlD8SUQevVmYq1EACXz8qxWjE8B042UMyQy8zDZhw1E
O8sNuzbxLYLHbp1RpxS61JqjZWnLs4J/dPgsZtvw5BL09VmBrgHMYLtk0WUaBb+V
gt1P82ap9CUEdiuYS2C0QVwofmFOdPeWZ6FW3RIEqG4tZFRr9+/CVZsliZr4r7ML
XgfvPw9QjqBn4eOgIBsM4Eagylj+/+Ha0hmyY5IQaCwmNK0z2KkpoHCGabEUqEQW
fU4o0kC1etTzAyhOfXEi039mpa9mqcLOPc1/rNZqzjF9CF8UOSIApcgTaKe3sabu
rVZOy04rZsb7qFcDEelpWRL74kol1iKrhK0uhs7GVl+QZuvnBzE4QTIxWXtrFJW6
bCZbG05E0OBNIQorMsJR432l3zh0bd91zS6EwOXE3q9YCV8wLjwNDc5rakjfnAnQ
f7dDkyG8i3baSKyssZcpcXg5RbBB72q/VLd4hy3CsRjlvrlMgRPlK34r0NCn1fgk
FLTlNBBHZHvcObZ2y1prreFeTtY7e4YsL+LpULHbCLwKVfHXcyNeacwwnxIOZL9I
by3auULyNqJLdQeFkX5mcPadVI092HnyWFriZVxAE40nl0Mw6c7LF3ZrqNMWGEgP
2vApdpmmW2bMukizi41Oia1X18THnZpN0/8I2g3l8kwUTr+8PZAgME7Ns9wNvcJ/
6paDtP1uZY7rLP64vnrVe0D4z7hyZb41ucM//Ny57nzhuCmnyoC7c8fA1o/vx009
GBjWmW+XdtrvHR8hBENxBkAEthuapdazOUDssU8u1bU7gcciDyWWeP9Bpor2LNjn
LixPBsvK/XeHPMRoJBfuGQQJyJrfGrdhQZpzYdcKN2+/Nn5Y5VJ/Dv/Zd7HEAl2P
KiMgFA0uvtldLhzJtmzeoqaJ0wJjV9B+fYqBAEkOFQSguRjDXEoRiFRTX4xSTIgN
2pGCDDcKiRqOjErVySeLkKJc8ElNG9dCiCJ4DC294/nfc2YbP6bF7FBERFRs2jF5
1eNoBNCf+nL4hRXn3FIE5tjTJLy09OVdNDq7YvhId+CEOwKgp5dktqEYotYp79Aj
LPLJiVzRcO2sd9pWHRWu4lpQ8XWMEdruIfh6x3PkV5Ca5BTtH3SmpJJlwQSJ2JpV
j/hm+IwcyIeUs3k0c3/P4IoK3M6UQQIXKujj/puRYPc8bum33f+uVzG/rPjfpipJ
3RNsf/0XJ0TAvrLwbJskFTi6Ayj6zwnxlKXIzDDg1xfTU9Bk5zn5mQ8wLJjIrH9C
cZRjekfGlwKA+fpbaNKzxghrIsHO5A4/Q5ZBdJ/FMaaqLZ8TINKXihjE3wGxjDoj
4dH7WyQdWppG/HV6o87TnpzLgvwu4e22uQ7668jlFQ9fxZ05MqAfkCL1vgUecYCS
YpzyYkxUNGLHf88Bw5pbwatm0ejl95WQrK1S/llxz1/E4WfJiOiAGV5i98mfz2dG
TaBvvs1FQ+API11NQHcPKB2/RFNZMf7UUyyryP+rYzoAQJDJF5XufFyuZxwKO61U
FxWDmKX8uwcZIiYCuiS2iXzZb+YcRQJm/Zi2U7GVu0PSbi73cCrGC1J5ZdZpsrzF
QGBt78vfK6ycTAc9K723GjePwgU/Ei6rlFRumN1s+v0o6J+K7x4hELqKkg4kXt3m
MPepXVtC2rfyn0iwhtRXk5c0WMSDStKShMGMmGgkJ/yvQjborFy6HgRHTI6uDPW2
v9OV89kkdKAfLWeMYPEqTh9pWpad/KTgCj18sDoLcoyntvUIsHCn9SmEUoJrekh2
Ut5wtHOT6oPk0p8BTSVt09XBtU8djhdmIHCxZd7zt2OurcrXoE/MMexG/2BkM+GQ
Yl/fUpO3wVPPVA/oPeW7JHXsPqEyAonjfukVwsaq986rN/EE27ZYZIAbI0ks3MwK
wSPp7W8l7dusUTzLshBnipM2Qmj60+8Of6bRDZWdh8LNw8ufB79MruD1R8N1Jy94
DQneyv9YcmsL15yK2uc4T57fNazK1cUcFVJC85hvjLt33SYsx5YAwg9GYP4CXVb7
/mVwo8iMXefCbKkxgduYkRbyixNs/iDTS8RkeSgKFLWdErLsHXC8wpUQqKMu2eJh
0GHIc/AYm4OSxokDXCYHgPkw25S2YnNiMFiC9i9HIINJbCzsOimgy00MDJfIAv9p
kLWMCx+eMvhrQDUIHFHlsCUFSIPVk3e5hRks+Ji5+P6H4ROHdQSsY8uV+UBJwXCP
7RxlGbXELpN++lIigAeMgg1ghnTeICg0z0nk2ZrxkB+wqGxLy/y4S1yOiMuV9pI4
mYu+mEa3Tnp630hihkRMGXSi0tzveEgYC0Gh29uUJmzel+VSLAwxX9L71QEPFktJ
x2TEjBzVkS6vHJF6gCV0fF1NrhFEG2YE8+s3DgHATaIz5y+2EzbQKXUu88Cx/y39
DF8kRwouzYRjq9qn0la+kb8m3XjLG8ocwQw1ObVjgrlF1V0qhJueNvNrM9H9kRLg
bYSt+bM6H5lXG5FR6UEoTjRElDzqtlSJfErkfwd7IGpSfHd/kpOZdpzSV479PrwP
VtmDdfKxBxyBY6C1kD/u8Ctr+7Yzq14cZoJr4S2ficGGeHfZvc7MxQtXoRtkeTjV
RyRwXB15UFsZUX4ctrO7E6ea439l8M3uLDATsA5KmfpAKQ+/qMchZLgioiE9Ghcw
49+DyigzOsww3xj4OMT48DV2efbD2+h23oQUDxHLRW9AlZxgTLf1qdgIzM+vsqki
QO5hAiVONE2ys6DDfUXdj9BxAZO+6XU9tiE89WmQEPyEEwcVVXq1cl5cKxKa6yzt
bZFB7Ot1tIeaKZpE/DaSnkSOd5RducSYJv+/aiH25TWhChUeCJYXU8FTcnusyUgU
Zp6zqhmXeoMv5HgrqMHU9y2AUF+gpEgP0yungXPAHQbfr+bCz7LVw2NOVrg4uZ96
VJy1bwtdWfqM7PbCP4ebab3cktzWduT6WPFj9QxJKOGVTGwJGqrbD5ZR6NtjPxJL
U/mFk+VAARn+8q9QQNmzAfGDZjKSZv3T4dniv1bYYSKdXelHhpTmVWyG6enYU4dX
7QQOzJB5esrQiMm13Y9/qWoOVUsC1La2dRCYRVj+UUBVHMrdoaX8MumLafLnFsLq
Ft4kMxetrVn94ZewDbqxv6qqSHulikqq2jXdG3ux7vQvvkl0570dB4T1RAH0jocc
C3Hbg7/A0AD+xYoPnUlXjeE/OyDYo6QnSaL1LUcTVMExIgmpaffinr+A2H/13/05
c6yWR0RVQqGv8ff3OcwU3UsW9oNhFH2oRpANUmqDyfugsDG/wREeYrnxcHo2mmuX
HIsrIAJwy8cDwzOQgy2VXSmts0WVLHN0kJvSUBEGUh6O0VcWx8Tkja5X7xukLj3l
9UiK5n48OoCzmMk3OBeXH8aleuXITa6JWiUQc9AtYFZ0aksO3K6gP7NePZzaehvC
aPuMy0Tyxs/0v9xmdg00MT+0RcMvu2Cpu6CJKtJHkwQ3PU9tRtBnWBoXtXg+VC2F
/aQ1jDyfxHCCiVcac8PdLGKW4+5ERsaK/26MA3crox+nNOvl3HHUwZqF5raH6Awo
grDhdKLVh7iHhR4bm9zmmn/Q+ryuWQwT8W9Og7zg6UcZuTPwz/uLYjgfbaa9nruX
OiverD+tF8K/RI00jhCP4IYTCsQOlAJU5l9PXld9SnuyHZtodrsVUuajOBtwD+lv
TAY07gzvDYDBX9Lf+ljid7J1p+qhmJqAPBBBlmPFSgADapc89TTn7vaMw03lk2By
xroUt4qAAGx9toviZUbJSAKx2l8R8ETEMG4KcfICEqq1RLkl9TlKetbPQRXzM9eQ
FnEkrC2uQzIkc2/yo7H008GQBlfl2YYrzys8U9gW96E6rnhTofSgcEJ5aSH92P2J
4saQB8CTikKMFsZn/dsqHNO2/mlTHn1qAjRCAGzlFNe0VuZwSXTWgSG87EWUD/AQ
K5d5lrUmjLrsnXblLt8ytFP9NBlk1vFR8XF1SvyhsGj6xdTuJFGjGiRA7sne1wq4
Og1iIGnLix8HT2fwyH53PHyb981BYYzd3Ly1g86hfo7hH+HgWQoJuwoko+tiINSO
GRiE8BLbNWpFFrjrzO2xR9/zRJdFmI9dp6IqfJzjsRg/ZD8rt4WSRvl2dsHfwFJG
4OcPTqysULobbDis7I59fLnQ/Yeuj9d7PUbyFCOo4h3Nxx635KgPqCNNd6R+8zrL
6mqI9+EFFfs2gfgkXaDsA5JSvvgqjySfsys//UMg9AmnH+RHJHqThtWUW/7jO4hG
nL2vVr5xT3d1LMpqmMzc4Bn8NrCAHXixu4y2ZDs5G+V1CRTQObO4b1XT0vwBwijf
L8vHejWpROzScUXb64V1+mLqQzCRmo5P3erf50fDEmcuavw+1OJiWym/MZ/hkjx0
zMmPiREQf8pMo3daIdWPcbf9oy7QRrfB97OcE6n+V/rtgOrXgs9gDC1+xK72LfXg
GzOK7ZTLlIcueXLl0FcSMGma+SOgVRbeHl6kQv2XkqRLk4Ql7EUIGrU2rczqpjtu
pUOkDuwtzsDLsFGq5o81X64TWqmXsoI/K8P3ftw0LHExOs5RToUZW0H7VtYbc+bF
BF+HEGRVllbRQgJ4Sht7ujk/ElYB8vzs3eiJRGg1Wp169K5BBPlzae34ZXFxDHTn
cPZkKm4WXDV0eU48y7+L74+LbSYFZCtmFq2kmshqfHsN9sIJkMB1AzWwFfvw984x
yRRTf+CUVOijExiGTz/rn4fdFhH6qIlNSKkJ+6OROyB7qp3KrJbO9ZtQ5qwSM39B
3gqYDls/+LgMfSlsHB9eWp3qWvepfTj2HcHmV/xxxi8rJidF7qXbRqPXy90I0wep
cihocnKrpq0UOJ6ElQJ8NJwduikjG5c3whaArioxaMa6CjEvzHsnAKXx+WXaP5sz
HgKHiXqrmovCWHbTIIWRlsBcmYDwQscB8QzxpXod427vtoAFMAog23GiM+DewluY
jHPfKgmDcSL2bTYHJAWZiQqEoy1aOnylJD+GDEIl/ZcutSGbet5+fWnQ+A0hK8/3
JyDwrS/I3EXwL5jDyfuF+Oqdivp9Tvg27c/iYyf6cLPigoBJxNPV7l/HNdre4TWT
UU/AZUmoTe5N4JkhzzWM7FftLICkgOxIJIwW4e5iearBTDUFkzkiwH2vqJg5rKp3
/TjF+pN0pimvR35Oft/w3u4jcHeMw/3TOYlIWM90dnJkK0T/lCXshCINWIRsR7Tn
foXWYib+vLekNMgokoccj4o4p0Kb5S7RScX/7EQJnUOBhgUU81CP/Uwec1+Q1lFb
17cWaZIPHOnE+cpZE6hCRa088Ol8SNMtSXRNDGszECtwhvmPwLi+cU9gk7Sr6XpS
p46UB97SQWWwhTJkWEXG3ug0r1w+imqS/bryogetZtMw/QyMjHBUEhlK9PwuZFIL
VwD2vhKCLywFu+0xgyiCRhAEVeA1JeTpnp0LmmJcSCCdXFCSKJqrYHDVrsT5Tuba
OtOKtoimK6cV4rJkUxs8LheN3kzXlwSM5SGBYdWb0EwaxethVW9hU8UsPLrBfw6B
kfp+PJkI2mBIibvlfbI7t7IJNstVQyygQYWnkfgpHpFBEY4waAMQlv9yOmoMcfGy
/0gajt+QXLRM0J9GjkNcPySACBLWp/J981QqTTtJ/TrYQtDd5ZjCC24/fS9sUmGY
QMe2oy0H/v+x5C+Na7ex1waj7xNE3UmxvkMiSJ3kNVIvymSlHO98Z8hM+qGvMY0S
Zf/I7vasteTHFrWxoA/PUBfGd+wNypTTCiAVJiFJi9NCpB99F0sP71xcOBWY6dX1
CNLDaZ0Irc/eknW6PjlJ+P+DdD52HrDBx7i0V5/mee3o8b0ydWmlw32fz2Prxv8D
IfU2NDL05LckSjNKywpcXLJ7MisrskIr/vIQHLviVvZ5MbpLK5mLUbpEsaqkThc9
c62SOFuKdE/jFe1EHxt4LOjOvWBqMw50VPPTOyvUERM/CZ4OgBgxacWBshlILjKL
X1k3r8KoK61eozX/S1Sx2qD6vbWm68BuIFfU3/hnA2ZfAi19zYZxJL3i8bttiSXk
mvyXHiaPiNOx8N5xZntqJyCol/1OeaIl07g4FfqGginhI8a5K8jKGqI9JvsfC8iE
/gL7iDHeZfZByRKOXMycDZFAA717hjkX11669/afyzTb4JpsIjjCu2ojTtYDNBQk
pNngP647/7lwHnRY4d/BWReXT8/t8oKwyDc4Uqx7rIbzpcoYFpRJK9VTdCFQ6Rjs
dXeX3s2LjlbcSFK7UjNGZqcdgtYy6kuJX/LQy/oCouRja74IHL93pWd9mStqZvut
ll2X2AlT2chUXkDho3fgcnVpQOBTAQjzVDa1f4vUTmdXjzGTebayzEwtKQNRPpXF
KwUHJ1YGPrGDTrYUVRpN8j8ysEyCLIcQYhVT/6IRXn6RcboDpV1eTV5/6ZmEcMwo
KmHPCRQEsHUXa//ijR+ynLlMvrxa21SLJxsPwHup0LRkswcjD82CgDWOYgujURvG
DtsHfhaJmd1RIPBSdr1J1mAsD4YTspjxrF0ymBqyaFz9GenEf4HEg0BY9766T6W9
olzshdryLuGvXXwdEh4ruCSxIqSt9q98OnljtOjvwsS7YCus0yVQWGq7YDvwJPc1
iD8/EWpUGUwoPmWoCSIZuvOIo3O3W+4KTp/cF+y3kuMtUj5y5qm5gzbvRNIbC10J
OZEd6CRRMQUaqvR74RnAOyP76gSykQKVcAta8CD3cCYGt3S2iPnNEtEPa0j6gWAE
eA2Ypp6s8iOUCmrAXe1v3ebmFLKfniUyPDWwCZOUY7X+tY6gmPm0TRR03/or7yxc
i7IdyB1X+t0SNlP8dg974lEK/mhUcMPbsamIK3PLEMgCEWbfKhGcSX5hLraI0Fo9
FdynMMFeRX3kkQg7NZUgp90He+hwVYnKdoUh3emCXjWKO7x1LOinwTkLwWoZJfhl
srtsDySsE6PazfuLnaZrEEFSfpLIKe9vnUsMW6qB2y20QasDlSuQCGbVXQlSTF73
SBLzYmD4M8DPbcXKVwa7hzE51bjwH/4g1zs3V4oM+P8K1dNHauQm8fwe4WkTU+pC
KO5GgT8U2VAkwHujPIqxjVIUrIebHuEfnNmbOSTunagLsrvRDjp1U4hbifQ/GHv8
aycZ3UFjLinkUFgpBcsfhDqC2vfH7IXiazROQfzesVf9QOFagl6naueXZeVaJLH+
hHJXhYVB2E0BFLEIrbSgg5klE20Klmlo3HAHE0E1rOJJS4zJSAiAhyAsG68HBT4c
3DxgFDsDvoQVDYrKXO4J9Lse51HHvXS8IpGZ8nnW4ymb+p4NbKalvucxjTaBEnCV
r9T6xtlgL0rjL7HGl5NlAQI+nKcddfIFSLLV1osGGUcJVNLnufB3P4A09MA1GldM
+yxcOjkp3GFh1YWTjm+tDjC1wSgBOGVORuVYCSWPdZjaQ54y1CqFDujkvB9cTSB0
l8pZSFyI6eZ6ZyhJra5ukIBvSzhjEnp4HjsVyIT5yWMTIxehsygZ+h9xrw5IIknq
AuWszMRtggalJwGIV1zgHFcuSrKqe4sfAwRWx02acMlP2yhto3OZDSlQzqLzDkIw
KJ0BPZORRfISNAxnZ0euGAHz+2c9v913g84LTCUFdlBn3sXqsnyI+0H/AUU5Abo9
rB9WgD1dkJWDN28etKGb5Kt4GJ4HByR7T69KiPd76AptSuwNzb1lNSeJBkYPLALD
phpixbrWY3SfVTHXrIRmFF+RZUo04O6SdoytdGD5W4VcXtg66AHeiFNVg+Y9xCFA
G6ddWASNXRRXRUP+ZQ3/i2d0pAePVNzE1jijWhy8Y2jFKNAHgh8Pq5764BKlfJXh
2J1qhN0rOeH3quI2uay87EIlCuz96R+TuujWUn3grLchtyOmsvz/sUJ12rkbLPwq
nxs+A1PydzhVhSnlM4YT/6toc3uRNfBKo0c/LIJIJ+HZN203/3wMpDyIhKOjT6Np
sxCYlSJylLTDK6qdEauMqU2WUj+t/+C/ogWcEyKxvRl674WZLdyoqQNkiegWURPG
MxxxSpWBUgDRfa4yaEH79hS4OhNcsjQQ73qO268EsQtpD2pAt0VPHMjo5ACdI35O
8mAYNaskeZrJ21YVBaFf6FnrdYL7W83DbS7GuUdfCFxd2HnqR5ArnPJSRHPbK60k
WtZN093lHw+DmjKILaduO4YADCtOMt0b/+UpKDUVL6saQ01UwrUuLSAvNp7IJgWq
KcRYS4G73YKkwVW/970eu3SFti8gZAzIeuH1Xuom+aZgKQ8ms/OvBkzTWDFXSVSk
cUO2jAcUh5XWwxWuJWR2UaobD/VpqleJUAIO8bOGa3dWMleU3Y2wJe9VK/4UWzGP
+82ayk2u4beF7h5Pwbvt2k8hOcfPiGNQLt1AFU/kFlddMDBIfQZtF9pZ3EL4imUn
UUAyaaEbjp+RIQyP9wW4rwnrYRiFoBNwFnJGJkjYzn0NmxZQ6PKL9TbqhtVu/iW2
XxLsqpPXv5Hzgp1Pa+emnrWfROYa7T4YEP14xbnZm2kSBv64jpE5mObf5s8JeeS1
LJjuqvbQ+WQQZxpZkAvOIfMUmRBMSFAks7A1/alefQpq/ZLlwcjqAvH+RbmgBHDW
iz+q1nifDCiq+oZNtbAkOwYCKQMonEVuW8MfZNlNPs3sGJzeWXNFRSmEni0ytV//
CiTH67cxj88B97sNru29avb60A/4VQ/5DwT4D38pDZjRD0WMitcY0sP26TvtgUoR
OBpyTXqHVuGV2LDOO5XDqwevH8U62hlUU0nqWHmAmOmTYbFZspoRkYHW1sYEoFGj
8nSbbrsvQ/3LTLXsRgJvYgSBFncd3EF1WrreGvpbLlcVSfkCo7+Y1+7LStW0qUNk
EMYQLqsWd8Z3A3AzpigaWXTpRa2DfNcOPSnP3bjXeqHCQHiCcpg6oJURz5RQ858t
ZGoUYVymtWABZ8rY+4rb+0gKbJzsa/dQT9oTrJnW0m8BXL1XVdQ0nvMlCEgT2uki
ZEMzmHGK7cyRbUzIKi+vKUSMx3Azzi0z0eC+L1nW25XiTJavWBTZG2tSzq3HLjfu
Hut4izugf+spPXfqivtyxB1pU+mAG8WsENcNYExYaEI2rF4vZebpff9HL/PoJ6FU
C7/kTFWDJzwb6/ud7V62rzWRxOGVioApeFW/InZZqPbyawK0HtdO8g4XNCfHi2ZF
VfwsJqtvR1ZYiGJVxZtAlhQMS20vIJks5TkXafN6RuIx+fANq+8g8//L5WfxDJHe
bV876xWYdv4TuJEmco2QugWEHq4kp8olUe23e+3AuusZ9JP/ByD8PCEXbh3VcqJD
5r6R3agpmafrDQgHWL5DtW2FMfO96zrzZQ7AANbGgFolXiXokCqC/lhyOPoKELfL
EyRwXvHr0sWBVBXNBusw+57tEC4etzryp2+W7bT9zdvBt9QQdgvVe6WEJZH6EKHA
XQ//Eo9pKblYl/KkNOTAcsBGgUb8mA7yOkpZ2vbHpr/9bFJC4UKwTDZlPv3SJxMr
UC5rydnFRT524jx0v4zh2GxtL9ya2AFfy8mOoRY4xFog4RNXGFovghQ8uZ5oRcD5
DSErsgcS5y2/a+jiXq80PQbE843sP5qCu5UbaNXVaDwSgBWizrjG+e3bNyX64xmy
HvNVAlX3qtBY8igWVr63wMdY/KOxplxPo0ePH9PWmveL7+tjjtAHI6/UxGfsGlvb
cRNpMk1/KzGdUui7xhGMd6JA56UqjeQ8u4WGUMava2Cs3X10foCVVQAYgggW02kn
nAeHlmG2hFkqIvcDVLjkaQ6psqgzlE2jTUubcy1upyYBsIPigc35I8vHMbLFF1Cj
Ac7+Xsif6iS4VwE0bCBJ5yS3KbrWFqTz+9vL/N1v06esOJDtfEc7B2tbsiUXhUoT
2/Ji3OnjamOGHRKdfm0sY9DoaSKyBZJE+vYlg8z5FsohsfWzthUcLGIKgXLRnKQ4
8S+MbnmZ+5vXdikfoAQE+CjDUQtOKO8Ss5O+F44UGdgx0ghKkaLz5uD3DNag2lWE
XEf9+mbYiGxLtObW7g8hDwBqUnqrtKNkz56v/7QecyRaFoOl2lN42JHIl0W9MtAj
9QGQwhxnG0P4zpUg/vEe0z6CL5/oWpD4RSTp3EfDFYQRTKzwcjNgCO/j63R7W6QN
La64WlpLQL3tP4env6t6uxPExpFKte02YvFwpbw6GDq7bZ74hb08/axy+Xw/+yYr
O8mAppKTQF6v9HGLQadmOHOsRvAsB840srfoZWcSO7cfXaGbbouXBPBUrALYFkSm
HHuILSMTlMZ07ExgeXD+pMx1x+jFWwZdfdu+FevmNYJgOgVePdnjsQ6YhXgG8uh8
Gg4TIyTBinUefb10Ha7pkUFE2/ggdko/oCzofwedIOGZEQa4f2BUSW67xtoT+uZ9
W7lXZXeAG1WQRKB3gcvB/bhjfHwEEdSM3uki0yihpanHEbtydrjsfGokOEBrPQe0
piTiR/+Bgan6ywErzzw3nt1ncq7eQZOQ/9KBMPlMdNP5S628xNWQHnDoY340KNjU
0N9darC+euaulKqp1T2jFTURtWnJeMb3OwRAtLhUpq4NQulgCJqZANUjWL9/D8Fl
7xexWjp4pAAWGGL8KSXmTsR6rycN3TahQYGczckTpYkQyT3/eAIjBI6rf6EUddhT
reAKqMCu7iSojUTwDwto5mnZI6d62C3J/GJqjk4gwsOE6t9WKVQwkSNBVCl99emQ
H03v4+mqauZkzUbOPrIoQuYwvUCDxmHH4cu2PE8qIYrT1twiVzAx9DrnNSZKygLb
j+brCZfZJw4oF99Xa+vkwTuUfOCWF/lX8sC76rqNFqMaxUGgpRSZP83ndEzNr6uC
dJU3REvzXOUecAS+ZzWPXAzfPnj+dkraer7e6ihYUpi2WE/hoWCgo4LFZJQAL9yU
OfmPmgkNBsCJzCArmEh1ypLlozBkAAmmN73TMDtTo5t111oBYRrXyYNbdvdbS0bB
cL7FL+1rHzCduJxauPl1hLPfiXe7kmMEvKxNEAAH6H3GDwG5JFh7V4johzkOsA8z
HrD/S4fM65bpJV+5bqcJnFwqsOmktd43/27lMqR4PyeUE6to0t/mwAEjVsdTlSTW
b2kqqGFtgYpdrFIcHoCglD/Be1wX75HaQa4FioGu5tNslf2dxSqkb9ge2trMPhW7
Esk6bBfjVQ4PS+EI4XY7lZeMErZ6tAR9Bzqo9oEn1HpuWIoYIHthLMwHU0uGjy5/
lq5jqsSEBLitaF6VHJn+ekAJcIrz6yFnzSevT8fPMRBawZljvLattMJID5ZoT1W3
bjNQrUAYV4I09pTrNpVZ5TDGqJhfKcfc3eJjq026MvFSYFAMedmAb79a//I6iyP0
4bEt8znIG4kq5IrDmnd9i8JMhXH+LxtZe4Na8xROMZqmkPh1k1OEn5ahl/s/93Cy
iZCPmj3qlGUb95iBzvhVsaAUqDfOKj6Xdje6YWY4+ccDX71970F5pGPa1bZS+WQh
t5vNhIYQ2RDYOx/3p/luhpx0aWZaz6eWOEJGSxR6NFXeYfZI3LwsTv0FtBI1QK+y
sCIKCD6bNDRWOGsrouZAShYYaBf10cXcN5xbekXnDjw4zQxqrGhQH+hlG2AgozbM
0spDFA1ZMCBUwGmvlfpXoEV+6Vzhb0mfpiDb4oPGFGYxnaW099+3AdylpZyCcxYc
z1ITGn7aGtRNlFxOokBtJNjnXS1P1mWRZV1urBWZdco+dLjG4n5wwi8hRoa3iAnH
kqS/gYri84VQRol/8CY4BODVFBjtEnOKi+aICDPt4corwG/mbwyFhFOv9Zvb+bbR
ZcF7X484625xdF8/tvV8G4SZVpIuueSIW1NYku6NAHvCXbdAT2urTcmOSPwvF38s
2APdtedkuzkilKJCdba23T84R84SadCo6gAsMgtKgKTglDLPU6/NrKJbexivbk29
Yvp15udJC3YGYuDI1aYY2Y/JioBAWUuzheVZj88m7fxFUDiDF4t+M6xGKdPejGvv
JSjPq3pql4cUHRJpXTba9O3BvG8dgQ3WtWgt4Dhvc1VKy99WRQR5nNpy9LNGu5la
vVF79l/ux2lntoN3vXnzRCG36gQz4DFOPLCfE9gfRi+OqblAhz7RSeao4QnOXzek
q9X+JFVZC8slO6Yu20A/rqgAvghxIq2lCfugVl53GuX5p5Spv4rfvK7hqMsASxU0
RRV86iWklEUWdc/IFpibh+rGbGuPb/zcOt1tOVEZEv6yTJjx04Y65sBZkmhZJGwf
WVQKf1jh4/PqnwOzN8uHqhblraMaiDudFMlHB4xZMCkIGHEtzsBKdDo93zgmizRl
YvIGplAyVbB7U5NG+gNiu3DnSJ1CmSpv1aHz2uiRDFnsjVsopHO4oKhjL9Pz/l2N
jkaj1rfuQGUyVLl2yFZ6OFCsxwC2ezjuWGQI+GbaZp34/p7PBBGfrOYqAguQgXxa
vYomnYFcziXtDYLnkR1ZvEYdQPJ6q9sbe8tu0QQeJbkAxkgAXutA1sfm24pnildc
cfE/b2w3bjf8Nz51mLHXgsEA+WpXh+eNJ1mM6YTLEf5dQAfVOEoJfNTUv3/h3wXp
iXUVCHKnwgxERZl9zQV/0UD1C5+RT5lt0OZmY9G7uxot+5QjUp+V58doCdw86BP8
lLCRJvQE6UuvjXTmJ0tGF+V4ZmuwceL0ZGfQZFdDJ4+T2iC46wQQb6/WKmd3rKQF
BZMAEfte8mq5xAuJfxc7HyvKlOdmOqnoZqDhs4na4Ynfa/5j50l9RQoelKD1IDUk
iAXzBRDbyfdXJBHYjMpSVMm9o292c9L1s5bIwKoCzy2G7eMTHo8Wwak5Of3waY3o
/m5HQ9vHrVJNY40hvpXt/PLEyx9UkgM/MjMkiEZtyOk721JUpHHByw+JZjqIDnQY
tax5Fc150/OdlOQ46d3A9c1eKd9mp4jQYsWjKvVJLOIFZgHwgcAJ30GCrvVdRlq+
jd/828CWxcX3yjIygnOQ7CfNJ9IMF6ego5V2aqRg0StLuVaIpa8pgHeplniewbY/
LM3XFwzydRVUZejzKRUjFQnoCOoBaHiI2bF6sOFq8hn2WZjLQH/Q96x96onyY74O
6iCCXCYjnfKJtc4tdhbnAXu9pGOqnRecyCs0eaNjZxoyPgKo6OwxHXjNli+y7eEG
af8kY9Quh5eOnsCshLlcnM30sor0hiRH6bcA00M0YI3FxPnsalfl15EQhLmSPFba
TRq7rpztjRGvAqdWuQqTvtEZnZ2W9SPi+JTxckrk9eZRYKnWVOfQLg8dsmuufluG
sLEdWr0YleX3u+7q8TLsUNBZGoMAKQGjN83jENGg/Nj2MRXCcAKZSJz4mgeed/Br
6IslFiqXQsnEdAU/rA4L4tQMCyvveunGuLyPbnyc6MPRfIA0HJ7JWoEEaOK5dGFB
Ss0PqTIxQ5VuA1IwBjPFj3NIDL8BBW/wXimEoCPrFu+7CBIHmL9ypa4Qaus2bQ3r
VugosVvx+VkCBSK89lzoycjw95A/XJ/eTgft/mMppncqOa/dszqQmcDTPYz7QHgF
g5A3ZttUYEbmBOIkzjaBXz9qSB/lxydj+B+TfxrA0TCBiPWAvoY9ms5O3jxyt+oz
/SPNSfEwDbLeJwm4mHprx/JtS/2tPRy5jpFU9sLtYBHZdnUvxovoqtVCT6FA2naS
ny8spVtKxAT66FLFPDuaE5y6xV5CCxJ1nZk3FihA9O3jYHI+Kx1M7HRBWTiVXDM/
Y3LZRYl8Pmx86K3TYm1NvjQbc8sPyHcoBVfzBurhXEj7SK/Y6vidYBlWaSpi6Hd5
WoCDGUdJrtpTjNKrskTAW7sQ/TMJqJkyXX3XD9Bs+9XUAaSsnGedyFf8iaSviRSu
KkMtIrZVtLtPyXk6EbTv8r+EufAooK3RVBPJoazRIwXtCyyISK/gxL5s/dhwxZRF
8E7X4NklHA86AVrA9nvW93yfEfvm9jNs1b+7baHfFxvx0PrAcP3SG/BZoofvRipO
IYNFjWtddRxHYMRtc7ivbnOmBfsoo0UC4ebfhEr64zfoCNlDAHkWPGOW2jMUMVjc
YPMawtrsRWHN7ciCCx6li7TkW90NJnKewKAcqk0qgIlsjkHW7IwQysn+TR2nkU5u
brwRjHlQZ+Fd7MGITdAwX5rlBG9WjTS1iPfkDO2KHvllI4u8tlu5f8u7H5Ep+/o2
iZoOU8wwzSXyeU54fvyDX3E+H7tPNckKN7l2uF702hPQ7qCHEuPBwME87jSle1HF
g/S+/Roc8CPVQBQUe2+mOSuLZBpf/5/C7dUYax42PaPnTTfdZ+4bOocV5UEqLoS6
aCftEtjxVQETkE2cgty3Q8dJ4eh1QCeqGdwo1gcetyCwO9PA2VaOeZ+dOdH1rdhG
ghgGURDpwAin6AdEJMJ7ghmmipRgrHk6AGhoSOEJdC8BIQcQTQmWK+TW7vlsUVbu
B0lM3Cd718akI43NlTPsYrZ6kPcoj1BYJGy7eVeVepedfO6WJ+MTisd6hreVLnJO
77muCjxhCytA41OY+LXQk0sHYgrsw5VqJRTZSvJI8Fnlen/iQzB7bT2xn7jbY4vf
yL04kN81ftv8lLd7TjYqBL4J5Zr466jWekIkr+F69m7wRyM+xlFhGSjgm+cpeeTK
xJAj1HQyHUGLRny1rgmM7eWKV8AW+aITwJigU2Z0k/i4iivldNJ2wzC44eiklTqE
+snaaLcK1ib+P5lZGqMhbYxrVNjhAtZhtc/MD6LHPK8RmpJU1IXMnhCexB9CnANp
d0EqiDZyl5UXraWcadWGv3C6EQsBF50VlUOpWMg2l9GJUmcb4wx6fVhY2b8qQOrc
jGrBeedwU6RRDCoRSF5cT4BHH7PTEEpFXVdqLVnNiVAPEJmMFrNiCVw573GynrNb
Y4GT6XchZxvEOSCyaJTWAZJGDL2w6zT6mmDPHAtXIuELf6l+a0Tnk9VRVDXs2Rdw
fhop1sKOgP5fYRBXFsITfhYWer9gtNCch9ZhrwmkEOAve786UfQUPISIf37Y2DrZ
QpmuQ3lbu6Tjc9XYUtcG7OtoNhgkAFMdy8Y9UUtgX0VA3MYxC1NHPVWcxpRQR13v
O/2ffeq8btRu9JrCJ9xTfS6djpKxJmumOhvsTMksgrfi3G2FQsZNsiuVZ/kDnTMQ
Bb+i/TwHlvBtVylVSqUg22jtkHHjRNkltQNzkwSfke/KYFQ6WskVk58+DJSz/lh7
NuTmOnRv1RqicnfeheV8gLjb75jQy8kUQw5HeHNa6o7WC1XTCvZqDh5bdDLcQjVY
8einYichSuoKDCeP8LE2kiWA7z0ViqkX4/o4olFvuYGYz3QSi1w5fMRV8Xw8j07z
JItm2wDak7a9gerWT/olSp6fkI/830ApO8K1bbiCnVu2C0xNiorbAHq08b6OL4l0
YeF3A7CyzmwS2UCvuDXKAn0sgYlUfqOFmj9fn0Ec8GyKwe2OFOh5Q8NnXtNwGOPn
gxK3fG0osBaI2jNhv4zQAUK5bNjtr0WV+sCoVppSzyfJopwQ2Fyw+X+u2xp5mGkJ
QT3I85mHXSuRSwmfZmBFRoi1ZWaWda2kqkETULOPwssOMO6u9bdHdFPyqNyLHhqx
Gb8PFsp4Yv+6ZNz+FceVGYW0e6YzkvmqXo0BRx0n5Vhlt936PznXY2Ug0OXPAaTO
AcLZFY+EAsjBvwYk9cqzpugWnNPmiCPaiD7odtCJyEOfwSyt6aB/D8O1g83vNtLQ
XqaMZfGmej9QMFtJK3pYjji0VyGIBxmMnKjjDJurQgWgkEZy8heiBsxJRJDm6RKh
NmjIuL7FtKkfvEonWBiRIO6D3q2HkEwZo+RJFdKqXSHfNxsRUyk8wPgWCZS1AKOW
LEcGYm64/ldvygBgxHxMkUwgEoS+NkyP3fz4MqkHWeLMM8rjZ0SHT6DD4hznTd3j
Tk4toHqIfZuMIF7eavMUbT+s7nCTiRhwGp0+S+l0exgiLo/e4difc77EmQBW/0VJ
/9WYpaYI5PY8PbzQ5nRStZ8hME7QUhe3XGS+COWiYUbZzeRfH2DS0WSf7P/mBE6a
pUgMgvbsCblMrAF2bINh9C/Lfz79uvn9Wr1qpliiiOl61xp8xQ5y7X2xXdZNCF9t
wAxXD3F6tvg7WA9kfyp8q5PjH9ZL5Wj+Irpdw0C5YwFXAwvgEZ4ccfdR7Rg1HGq8
c6BAXwUoRlgPyFfwNcto+wZEgpMu0zssiK8labpuuXzRdNuBW4uI8qzLSugGBa49
G8qVVeHUVdk54UDKUx1a+9s+/xp4q6iCXRPcDEPWUJs552eHRIFHrPpKimTPvdlO
I1oWXmiqj0QVH2v8IKGzs1ykSVNFfyXKEN2sVbzF9xtMN3zEAulVtkwwSyNpTseX
jc1wDxZRcDo5aVw935eddzO2ReDbRj9ZfNu31bnm9ZrGI7JDNqoFyPXIMiylDgo3
LiGLkVrPYIbD4YIvv2/joppffKuPZCG61Lfranm52x1FsyfRhcDVsQcU6wAsGFBP
cAI56B1wMG/X15R4P8yeknS75ZVbY15oIRbm1MxLBiJWSZhW/AypSn3os17GwjGz
pnK8pPL61N0GEIs4EgLpt2X7O0vFf7rcvznmQAJobYhaEkE6vMeJ8tTax7k2jFCc
IRn25a3ALGxAZPKw6v4dYbojyZXB9TuM4ykcAQ6uletPjrjeewsqqhXjE7BfO8Kv
QN7OM4h4zLAIiCMrAl/iH6aKdLJ1Y6voXVxMM/BekTpU3zAk0l4jo64olLPvAwVl
6Uufgyf99YvNFtkb3kGWFuKjToH8EE4jKpIRqPylji1n3j9fF7VMfWYQw+1XU78l
YuOFrvghwEq9AbLL7Ovn5NX9BWDj7cbaJuf+YK3My2j6TY6cGBqhIsn+nFDUwH6t
ahPGyx28ynGZNIpKnAb5lnaomvZ01exWBAS7uO50VFqeQDILu8ooeOG3c41swh22
/eO0p87ULXNjbdcEe2KisIw3CykxcGWzbwgOGHgWadieHaE9mJpP8jLj4mdZXy8o
ZARlfRNfoCB0LEbQASoWMFbcBSGJXWmHRJXkpXEGJ5WxeHrdjlaVSlBVZGX4a6uB
V5AoLhaQpsWGnbvrVrxHsrghlRwRqFtsr5AnvBBXKRiJZwc4RhE4rfxV4QRWOSj5
ljIgxHlEp4OVr8am6CgoyF9rN/CQAEuSo7SQmoZmRSJJj09BJAr3kp+ni6GxQGsU
k4wmG5IlQ2pnrW+lQ686UdWMhTkXcnw0R/mAJvMmuFRnMhksI+z4Vvu9Nj0U1oZQ
kLhsEKQ9OczIKt5b8gA1HdQtSs/wEbYhWbZPQGfzABPANb1Tmycbwhelf6NDmFcr
kbTwmZ1BveLhWE+OVN+cZR39WFvU4rEbmpP607XokDdUNR8rvdsbHuYkTwkL4bw2
g43rMeWHuYyU2NBZPUC2wjDXnOSC2jEH5xr4L26mxMCAv9SHNa2w7BisABzy3KS9
fv5GYlNBPDl8PD58n+RyJpNUiOev6DcvctLOlmMWQOga2AxFCOfRAwjbT0KlQrsh
SCetRMfAEtJ7O2dGjyCJyvTd5gtqv1ojqpWwp9con7iF6WpCbitrw2YrHDeRAMPx
xp46nV5sGYaX8Fgz9S/0UEXDDHDkVSEUvEpaIOhBSmdhFNJPn+cTKOycEe4noOx1
69gGxMZ6bBGzxThzYOcZ4k8m/49AGKMyCoiPaw3MYLQBDeYnuaei6Qz9wF6YfA5s
dEgd1wJrm52SVt1XLmSLtR+bQeaaLqkG+D/Iq7VpQmdlFr5XftLWILCczSH5bxOp
ECWUNwIurtIE2mvOyRYG2sYWz5ylDUKH3RvcXpVe6Mj8UwTJpZoUqoYbMZbbSftN
ed2iHEm5qLPvpdPDOBU97PTrnDd4ElhjzyYjnq9TMVbYgzJG9iEH5ODLsNI0bbIk
UjehC5un3675Qc++HCapW/2wPQwE4LW2r7UMJXZvwS2tuR78f/0fgqrND3ylrSH4
xvJx9/SPKIt4XOqXFgxdzUA1wXLhv9ELJ2GNeihv13qiC89owj+1ShB+J3VtInTG
aR9OHzwvol4Dds1fVaG3sYxPQEtJzHWegOB5UMyMEvL14nUMmJTeeEnehqY+i1V2
7apAHSuWRkEXJJSPO810Dv/4qllb4G/zxFQTQhCvPRuIl+E58J4jVBOvNVIQt4KN
e1Ui7DK/t48L0jCPI0e13M6y5j5GAJ7D5DQ0piLVbKvO/Qz1Rxd3Uocz0D0UvDNo
JwHXagdV4danLi99hOdDhBNFvMwOy+XSibuNcQdz8d69vWJ2H9mIFRo4cr8c3WUB
79JC9N3Me6vCOIUYMpMn46J0tPSbIB0XA8loy09oQKa5uO5O4s72MAh4NS+Y3qa1
xceJP9bCtDYd0L5VeGm3P/ig4/2AnsaBJfk94BYZgKhjPP49KnmKKTJomLO5kO3C
EDmjBkZUFot463s2pqg+PYCCQ31R+aLBs6Uo+f6taz9BTIrwfjUSEmNylULlsgv2
2a+YYEoe6HX8A/BRCU6xLpNAAeHDs9bMTNnGK4iX+F0nZYrzAYZ1uPXIkdU7wY/L
nl9JcPb76jqCOpRdWZFWVyMRj7Ge6U1U/WpqP151uaTa5XhTbjvgxukqWL+VUuwG
8n6kYLnsuZNdkw9hR7lVrVtU/0ZUip9ry03XPWDhRACeCQVZQg94phnKbAThKj2F
CisajDFHwGT5yXGesUoETAQTrhFtF1mmPr1bYiFehOz4t2Pl5Tof8I/yJIz2slo4
jyhVEhRt/5aJuUFccELgYXfjSFpHEB9O9yEQ7HrlK5NCW39cXFX+BYTfdHRqF8Fz
7ATKTDIjZYhqh2A3GHlghYfFC1rCFcRiIAtESr3AGLqRotKTzWD7+xF0dHyzwtoY
dnNvWipy0Z3nabt9UyLG1pGiCc1XhMg7S1Rdm8IMmHhusEgQhSoOQtQ/iGchfB/8
tj03CEweos2f9zqHTw2zbVrBdX2CGyHDiDu8ElxrYXn0gjQePIUU0t4jT6+h8vIC
CLlAvMU7RaD9f0+aQIvPDfN1nul9XRdtIJ7OW2k6VhCPLUKls7l+u1+ow0eP0lwZ
74U7sdLQ9p+2qcZLdvj0pP7GMxMdZH9lC2hCj8oT82sIvCjZLVHpSsiDLnv6rZxI
gwKFaRaLEObAJqgmFC0UjfCJFu0JtKW087pxjWyABC/7KqnpiEu4PmBrvoD1oPZc
GeflJYRECsVBQTG52/6pK9CTlhFz2YEVgEM8+GZAhutICCRYN4CVco4kmuSCCPSH
LHp/+OfYz1So2FOVWdMjb/zzlU0wHZM0nuq7aG/YgKNMqYSrGmTWG2ECEbP9QjFK
bD1pfDZM3AOXzb2QYWFWPyK14CUJJa77NY6Jwzx/j2Cj21fuLLyf7cKy4D7l+VqD
9YJD8stqreyOlm2S/1jrIxzdNU0et9a0HgL1O7F6X7jQvF3hbWPPuYQp+HXFaWHc
pL8EFUjzEG8Y8sVX+gLhbABTLrcvqXjRCcWGAByWcjtyVLmFisDzDDxddO0RTLfc
OabrVFcNSK754qHokj3SKFo2DzieV/r2XayqWz2l6qnjpzCpRdqfbL7AUyNYL3y4
8Bv4xUzLEce/IZYNg6yHKPE/SYaQswK9A5V7Iu+H/Y24NKMAb90grm8Xvew62+dS
HOjLGdWpfYXwCU0sW/Lq3WY4gRcMHMJ4mSgTk1ox6bTSvDYZjlKqJA4+kD0Ks/o/
3OtGoqCpM23erlmmK/bSjZzI3i+WDubla/TA/x6YV6deYZ1cVVmHJ7vPLzEQpaTc
W81EcLle0l5hAAIcsHKkwbsk/R9iM6L1N3/+WtUYcgW4xbZX1DbuUY8roKW7LiG1
G9AlO6FF7Zvdr1eTzwgDlbCMMkh55CElFtpf/TK5881ESYl3nNX7NJ32/4XfHc/J
6qeEcEMeiiWBdWKdcT+RtZfqT5m5t+eYI2U7o5KERlNbPiTVKZURzcQHb6qYUhT8
6phbjTPP5PTUlywsnDb6EHhWd1MO/oI0IcwqwiqDfG6yuRs6xmLxiKIQ5kjhkT/j
PV5x9hwCHVAjUcs0kHHo1VOSz7vpDEXgJCOI3l+sHKsg5KmuBiPzYjZdOz16n0Ss
16IYpuDzWVBfEzN8AhkcZzaF6/fZfMvH8ADE7Jzbkvwho86rimMm80tQF8a2FEh/
Sj7jYjQhGNYfr+ErI6lxnqGOI4Y8SE8L5r2NuzXbddCrwAmrTHTHg9PeXDNU+mJH
/ryDBKDrBH4CzmtJql+l18MeyVkZ0TE4fPSyBE4MSJ1pNfi/VniIMBTnRpOQXrr0
yo3Ld3BwEaLTN7j3p4RMklt0KaA1/k8a2VP2jm8fSvn6soJPUf5yWmfFH456/3l7
2W+D2jPKrkBZuLP1b7+ippZag/SZu2D1u7uS1+PSvS57pbsvcNUXtwBf5j/zYod2
o91RIixGeuaiJbZ5Mhpe7oVyIJbu0qy4iplCrUcYmT1zlP7QR+J11DSJE4DvQ5ps
UY3iBBnecfpSm2/dfNtq8xlXUSMmN7HXrbTNZHZTIb/cbOtAADZCcaQ1wSzzzYEt
Jh10basVDBbIb6CDiGaAxP+OkYrH/7g4LOYiEYPBINEGzZfNtD98h0ccGmW998ap
A8dA5onsechE1w+8TPpF9yFaSUZ5kdlv2E1hjykOvJSIrNJTmcts2DubIp9gZfbH
L8GvSWtAhXu06pXhyujF3MvBNbuK7/pxk2tHibuWncEyGOXJP9aKxGuvpAa0zNGb
YJbwnvCDRGo8NtMMH2DQPwkFiQJ+LRHLHE3TjfbnTsvEU6a/dB4ac0u/mgRDvG++
XZ8yYwYUjXoYJ4G++mKSqnC9R9lXOIv7qkGVvxybO9PrShdGSE8/z3pGvmSFCzx8
sB3dIhElITPoYqDCIXMPjclpLrtM+VRunephtyrt8AA2/14IieF06wKVVk0ZKg8P
TYzQo3863qe14U66uuv9VGGiOp2rcC1V089cz6MTEoxR4cf+mn5RpEEauN2FO9tC
RU86xJZ2eIYZASJk7oOvKcqMXMgHi4RN2n2p7t7qWe8YWFG99w1XeW220KkBmD/o
+p84M7V3/lmIS85LKKv3PysAPKJNrtxDFNj08XbujFYSDoWj/XP97hIUVlyH0jeF
sLHGok8H6+iU1tYBIweIRPc3mxtXd4ibCuHLrspRIC8NnWisO5aa2X9aWmsbaqyf
uF480Nw5TL+o4aNFy+pEjbK/BG6M9M+oQsMv2OWgBInfHGtq2eIrCWZ6TG2o27sJ
S9AcJ6F/sfp9zzdK/kw/yEgsaFwImptmamM0mNyM5nPSqlBGpiMgnJgtKiD1lSEV
IwUaG9ktCOUo/AEqoKyeNGeaZuBbn2qpbq7c88FEGwBuZLEoXtckEXPEQ17C4zRe
8pnXKj6xOGBV2tDTyjXOko0c6CWh356T0jwezVu0BdBoA5pHfVmgPkHTIayf0O0y
KEj1husiZ1htf6rOPJV1Yi8mPs9hJB4IbhJzimVj5+w7WP6bvOyjGvwC3ViWJ03a
mdl4+5jxrFr1AnlwygHSkbK1QtGmPrv8Qmlf+UMD5V2Z9QqsTgLkbHiYoV2bv7zY
Qt7qmkWE4FkzCbu6fhupdZ+6awW+gmK6slHLmyYfUuhcl0fPoNLC9oprVBgp2Fog
ItMwErPBeTHrgZ3Eew0ia/d0pFQhXgj31JWBz+TFnOHK+qP+a65tDt10vxc/tBFg
GcR451WCkr1+6Hjl2014VmSqBSFmVYbYqvr1f4boBi7FetMCPB9BNNRY2ujfxrkS
Hl4ewewIntAPPuRvV4wewhE8eG/9VrbF9xHhiH3/xgu8frHpxS1IFukQ0oxnNZTh
VyVfbQFeodjrRwiZ3Ky6ubIMdIUNJIyqFRSgYGkXUvMcBUoB0uXd0VOfh5nTvqlu
Yk/QqwJSfRGCdmfOvGwZUVYLHSbqthRYibxlMQpsETRvWE2XvuSi9nIMkVQhv9KI
8oiV1MZ+CRgm9CnO/SQ+tZb0AUxuceHUyw1MLCl7/04hWosg5IJOoyGOhSsnLsQA
IFMOMUTEGoH9za1hEwMoouqS8+Hhy+gnCBAn93Wmuq/qpxzeDWumYoj2GgERnbL2
A5iWLWqv8pLfaAXG7udmFWGydlwwrY0wTt5CezdDq10iQxs4wOiM77AMvHQRPTq4
fm5CYASVgvFGbZK6pCaId+vpGKCeBR4niTeQewEt53pApXzc+0IvruNzhMDxTYZ9
DjKAgXbd3Nlp1THIs2uH4s2fnhp5hA7cNFPVDmecAGgOpSzLIHSB/9A5x9u8UK90
DADwloam/VFuUvuwUEHEwZn05XJgT5WZwVbqk3nlmeT073FhofgGHXxdQvHx5+Te
U4x9JB7qdyF2C26dOer+dFw28f7cn+ksxSx0wLBJXAnxMI0zXh3ALJO3m31h9rQM
F+ZPffagLRyyNtZtehL5vRyb8Sojl9++xo74ZDhyOf1OP3BwXwDMVwTNn5TBidzI
Cq5TjSe5paurNj9oQDXWX+fNj1vRQad4ncWMIkEAcpYqnDJAG16OZmaH054/8uIO
WjVzKRZWdLPlGe48UtPlazT6Ng3MCt6bN0fLupgZfpV0EiWLCiqqnmBDIwIf997P
xgHejTehltzdL35LUGAP38aRXhiW0gJ18qANRV8DJ7ACsVHKw7aR/4hNeAuPJXor
Cno/W0TxJjKU9ft2mf06lWv/Eu1GHoLaYlvOGTIFmIO57vF4XBxb9rDXGTquxi2I
Nxyy7TvQaagxw6vnqv/uIt8KY8G0TWi22XwEjLYO8fJRC5qiIQyCt37JM9F3igLN
URzFEzgzo3PWLNcwHuCl942AWh1zJ5HoaFQaFdXAHFtzqwNGWbbvOkpxu2sjGPjP
p4BWnupu4kqeoZ7v1TPg+DdLc/z8jq8y56EY6WQDD13Wl27MFZc+fVlgLiIqFDTL
vzqJ31jiD889LF7TyLFhY0V2Ho3IvvJ3s5DzZX5GGNj11zwy2LXUQa9rZcvdDM1q
eX1UIhvITsO2xU5CbIkA7tdmCqTE3+GKXi5ZP4hsqv7JFHdVYPOc+IAjoM+qmqoa
Ms5IZejrUnFr1NY5aJFjs7w5a3Z+5oFGWY/PxDSE6EucrSRFfaYTmf24139r3wZt
vN7Nr5PtVAnElncAYQp4UHPM+P1odkOjB6q5nIz8qDi/rj0syjp+sddCqFEqy6ms
Iugd+GnMfd8ufRNLzSnYTyYN54kjtO/Ldeyc9tSqZsJh4j14Ge4ZCp8pkIypwSk5
l0dPWwWh7a9zo2Y/+I614OpFPL6mKtN8URitLcMFOr8871bsrhiUiffbgP8NayRu
7IDkk5O43ZSRQk8hDrArSseOUTjZY110aYufi3V5xb/1QyK2wJXT3YNP5ak0sGy4
KDRvy3mkapGOCPUYVHxyKiTCwE0STxAl5kitVyjCRBMGzMSge2EIrz5DzdJ+x5Ut
koxxpGu/pOBzG+n221BJ9PkN5vw/jUroCorm5TibTNm6GSlmQ/q+7noQKVPlo+ct
cM7tVRyxYFL3a5aZReM+QQ3Cext9iyfBSyhDkWkUdFgvlcoR3dAdnIIaPKte04Ti
Vu86nZauiASbIiYpTLBiTlXZpt1KfdUUaHw0zHhuYwOZjKW6i0Ng/D+jHh/chW9e
DWrWJsoA9lTbUtyEaSYA284Aw3BAG55R01gKhn3zKztzO/nXOwxPcB+0U7GnWh2P
4hVSneWK7x8xDWq6r+e6lQCTditO5uYOPZ4mDQzS7OinaY0M1+45Ngz7fcE0Rx73
Rjawuj7xL0V953SdYKr5jeSj3JAueHu0FBdJxb4DZBHXhGlwBI2jUgMR11ucHWmB
BWgYGVX9yYH+dEqavggz7ta7pBqYmplMQLvkRv0uVv0zpWAye3Ybrs7GPq1Rp1vm
n3NnYllOnZ4yYeP/J+oV9JBgLky5bT8Ah00NeLvNzLD92opP2K7x/6rZy/aNITG1
Gl0n+TJLf0VAZJWlaMF+3lNvHFdSDoDg/7xNNPdphdJrk0TjFtfFgINvmKcBzsEb
vntaPL+1ruCQ1GKCPev3xE0ljwv+o0RyckZUlB/9dDAwVwyDorfyOt3hWxbc+ixg
N05u0uQtVinJlHsM9ao2chQv6wRQv/CrLIVdpEhuZ3nUDRV/o3TgHUP63zR1omz2
5iN0q3PqgHYPUWNU8D/4DUi0RSnMBwZbIDJGy2kYz2qGsaJZzfM0OFcrlCFASZVw
OJJTHS7PdqXv1e0Nb7lHWp2ySXf1Uu10WKO1zfJYKtl/0Sw5Bmg/GfdN1+KDyHyc
ycIKeHkkjSKZyco1iV2W89VJRscBur1/kvwMuGksFFd3jMmC7ErTlniWWWHpNupt
/zfv7O02NnRQIQ8QN+RQvs5cXfOvGYGkxMFWvPJ3HpvC0zOCNXTR37TwlfnkbdMj
+N3+APd/DycSZ4E3BFskdx0QgeDzYdVWX8R2Gk8pnCqMCTL5a/auwV4E2Fef8Tgb
PjyvnkGgs3S2PxNU2Ok2p4pFA4GwNY+AEhBUaByIUFKek24omhiMsjb2k/bnyg70
m5JE6oZpeFnfnAJMdli1+8k3siM2LlC0NdgwmMZRFKtH8tE11nhF2E2Tug/k02C+
kFrT22tNxK76GOnEy24GX3AYLF6CsQcQxYvfSC9CedXOeOavibSCjWhm/+CLhoiT
Z5nAN5hb3JQsbfQ/YIJrUSBTQbJ4fzB1dikx30IJGjfytNRYMAAIVZclcUyKLWUZ
Ku6L3y4PKsq2JfkoChwG5NH9DsbQRZ3zJ8jBwITGHnpvW7K4VS6KHIt7lgUdKRTq
k5Y4xj99ODJlFb4e7TqGQGG3qS+/N43ATlmKrZUdo3hw9OaSgVbIfJChzPw6WhYl
1Aqq1TfWH0iOdvJYgXqLNgYUuf3bCYmz9N7Ww/o/v4m0ujzOO4DOnU8soCftdsE5
jm3nj/bVAM0LZnDpO15iFz63kB6MQMLOf1EB4auoIVBl8TxIUnwOF51yPGAu4flL
GdqAvC+z73A+7C8ruiQowXUodRVue2qtl5X9656DgtyQ5tmSm8wCPYSMbVPvDj8v
Wd1l89OI5AzCqzoxum779MKrwjrSwLZojRe6QtOqTHKtLPA/tnYLqog8HVW8mtLM
yvtdS7vv4xed+xk70L2yvurl+TjGs+lAEZLJC27moccb5ZMSu+X35C3PGUDCkYUL
5yJkvE4raV9Lx9J3QTky+LREYEJsER2kDVCxKTPM8yhzNNiv2rs8O594A0isHZXf
hfs7AGhmS+b7mHj5zTtC0EktNE4Ka04Aar8SkwLNj/yUduuAp+bPWJ7d8kYRHTVr
CVaWNsCzIQ9EZR6G/P+CO6f7eX0FFrOHbenLqBz3pdo88hV7ZUQeEwJe50Q4N02e
ti2uVdjmMR9p8G8fOJOT7YqVy5EJ/jP3PUqbmRQg/J0IU8XAT2r2Q7Aasu3NsP1p
ndQW9AGKyXoAZUKYfGlPIvvaOcAwsnNfNYSTfk0JL8X67cBYmpm0v7oP9tuKFcCd
Fq6B99o+WKRb9A1ue9BlwShgPXWp+XFjMFzmjPSO22eQzykJTIhnDyCxBqPf+Gu2
OS6NAoKdZaR3W2DX8WRofEymf/drmxYOqdL1uzILMfHTyItSsFMfUOkjXu6IOD73
JJi3WHvPThNur5ggjDADLFJO90tO7z1tLu4Jj1rBH0FsGfMyhfcxfvD48w5/rx2F
cKJcsfZ3wUsZrVIel1eWe3Mdl326Jm8lRgZL12mp60VXeLnXLtDHF/VR1jcpdOBd
3GKdWbsJ5uwyVY0PCSa3uKfZKJ/vBDf1nAIZkG/TyBPmTjxp8B3HpwatHJEGlfvt
VtGtoGewfsDU2ZXGpGqnxGBabIw3vszV7zRgRII8AirfTrGOLEIi1CzximwKT1S7
PAAzmC3lpPKxSe+Tev3I3P2c61fV8DeFCML3PSAOaj9ihZxg7HQwM4AcdL1bC1p7
D0hplavrvhvp4GeYvR1LnkIa7gXmPc9fc6Dd6v7EtxqtNpiSG6ReFuLmiw9J6LCq
uy7AQuqcNIfpJjY50Cltkz2jNldz+V4KXi9IUsgsAe7dnaEK8njuxYHiuBk8ZRpV
Sp7fbonPaU+Hnve3E8UXd0uzW7hJiMFuosmbFhkmEfeR0iGFvfhLobMgGlho8qxU
xpzJ0Myck0ss9oC9uDZ8hplcZFtNJY1FOB+TihRy838aoxxc2216nAPPZV3v1ehL
NCYWFV6Y+KMyDiPnKmACe8E5Kv6fU4Y1o1d/48WIzuAaH/SkZSJIr8UnqrwpMMXS
iJ+WM0DQkPTfEm6MPa7uaPM/W0Vt4kelMHAcu1MeyJTZWKh4VDxlIG6er6ZtDJ6I
XqFwUVkBLJlx2KFy6cOJcl6/BemrnzyKdpclPF/3Igg7k/SeAROy1tsq+ubC86KN
rtIvMh1lKwlzG0kjejrnt+iloR/4DuZVAIjz1Hu8xxivhwSUz9j4qPS4Eptl8xlQ
WcTURKpjizaG22bHKDVDLRwJYAWoYYaUDz5fVkOye0QWMhZ+ZYXqP2sEBUnanyJs
guVtfABiBQViYZFyF5rnftI2WoR5iaykVg5zn4p4YUCbOkiLYd7eVYZn89OC9Q/x
wBNfO8ho8okK/YlnJwWBo7dfPOpa3QLgH/E0GaFrp0z9pKUauisPBF8w5WU+urvf
TXzw21wt9sATZWpSSJsh4YonwiBhxUtxrUuwGBBO3p+BiuVn3Nv2Ls69/NzccRV7
HBgUkjlUEgHF2DguJrOtmo/exQ2TYykHRFGywL+DrGL48TPEo1oFRBUJg9ssFU48
pn9z4zSABCvhxRBBsUBD4eX2OAM4wM9WJ1grIbuCIFVBdd2g+sooWppGLWCh6BNL
R0t56QWZTH6y/v9d/bSsblwL4IFlDnKHT2yNmTEp4QJuK1q0BUw8r8TxbKC4+NDj
2/Z3tYNhiSANUM/ubnwr85aC3rEfBze1dAgcw0kAnxZH+Ycn4LV2idJ/n1bib1ek
7kv4nmoicR8qYROY+BXg6YzDfOtBFodkTz7vjVl+PAuH+gZTNxfsvkFEXPZ+IWxT
UnzVabx8BWEg3sc5HwgqmyJqXPhj+AYW2uxcf0QQQ/UwmSh7YXRdZYfIwGClJhNl
XnFnCgqBNOshz3cC28ux3qz7xd1a/qEmMAT3/7eR7CchdrOZnWg8rT5oTlrGNor/
GcJXqOPmqBM78S69xxbovK5oSdB3UuwKVT2lFk4MjEvjHOGPTUjvsl9+W6cuvN9k
SIisxppv/KzNMXGjxYCbGeob0uPdTvoP/ANlvniEi1N3+HKdlIL9kWUcytURMTyz
7+qa2CLlKMyIidWr4FzoSFxBEVpYT0+zwd3SZSkcAARBRAXtJqRhoNMWkYSKJPVd
JDo/jgq6nGjDOTpahYwUZBMmt9mKG8oy2IYK55SxauaXFVb+kLxv70XLWV+E/qhO
sl0X8K0enre2KdJnlIs5DOLbR3iJxx/CJf9/wX5v7wbEpbl5w6n0+6wjYusEOyt6
dg/TYYvTcCWEzHOHPfLvNn7jIhKde253qEdqVrD8WyVQpOI2tHvY3SVDP+DrSiFX
9XbpgHF3G0caLcN8VX52g/+itCUTzDT1+x706lSmLV0SZq0Yj4tW9FM7CaT2PJCL
qczFmfMFSSBmo+HwhmkIJU4cvIiP0x6NkF2UcZO2eQVrpbQhN0DMhKF0QZ59tNd3
X10/U5YxJe8f3Fjd257xehnqRzMHk7lNwrw2v1H0y6Z6dcUtEIpVb6kzVOkxEWR4
qUv4toSnn9AjjvUNRXiY/o3fX3Xjg/NKDfqKQ02zU7trxaDbuJaP+/m/N6fBHOVd
zJ1D7EoD7e6zVjlxKLObkXYtce1t4SuKCbUivAz+/DiiIUin6I5Ln23GX0nYLfFp
ZiwXL17V48qaxvjJxsVwxEtOtaDaH/J1eDZtMPch7PF/7J8cttPA/XD/3hoQWU8K
c+8dTDEyb96SyKkDdCkkFfQ7meEQ48w0Hm/V4G1tTH0HmD3eEAXq617dmfrobKEd
d0mZtyIruQ02VUNJickbip53awZU8XCXlS3neGNGy7KsCzzcyA/flhEC5iWZEJ4K
mhEL0mTvQeWGLzdCV/yz0olcfAaMOialMtsGEQy15I25nOgnQPutyQJ9jnxEp+30
K1w3sWPCgjAzvTTkWvOWUAHwCJZgZrQjb94s+ZmPCdinTUnn1CcAO0uQzJ1VHKOT
r2IR0z8K+lLiyqKdEp3mH0ObZnR53pSt0kX7dWEILyeP6llrBv+m/RyT44OUc2aj
kMowDkWyd5iMI+WNPbbPklTpFD4d7qxp6Nniltg/B41ph3vwAEQ0auhgpBlhVESn
hWSwRmzp294x8q1RjH6N6RPbBFVOaVo1G5rOP7/r61wvM+3WCbqAQzHftu08yrnQ
SQRI5QXAZWLtQD6wM3qyRTQudCQ+nmWP1dYCMl0lDY7YKpVqHMOe/SAVyxvxGatb
RfHsGWjFBnK9wdqCyJpPcNtx5Tjxd8M6rZgFA8lDK1X9BtL+sHIjktMbgW3qBVbo
wBVVUTmUO6jc2uripN0eA1MBayYl2Id7K40AxN0ILU0E9BCKKA58JeW90ffd2qzP
c0Ysfj6z19EpDpV646PpjCgluvS/L/yF2AA153BRo40dk7NLPaIZdhfMhT48vHI2
DD0orySPwkUgf89FYyCKfLm/rHI/KfuHnXJcosVc6q+PHhNjgQ5XR/0Ip28aBIkh
I1BdJfLfxiihNYpiXlvDjn7LJLn0yJv2jZwRXxxiVhkQQKF5PT0ksDQCmjn6w1dU
422vJRFNJTqdP1WT0UEg3YunKD0e/jNYAkNpOcsRJu0R+tN/VMwI1HMGYZ/JYEmX
Qp51Cvh9okkmhWINyYV7DECbVTmE+JQACYaLaaLiwFsvQxr+S1krXrF76HB9gfh1
lvPzZOF+EM+eYh92yN+dYXePKqsi2lYvoe6Q5z5MLFfsOJc3mDepJ1CoK4Y+mjDr
pYOe65TD5WMV8FTy1183+RRGJeqL6Vs+h51423hTeJNY+96vtknBG4Inrsws67+P
yapmgEU/alJcZRTEjFmIS9qoWZOAc83xcXf1lEToyGh1RljDNBBm7sxfnAxweZpb
ExXvFHHKgMENME1RTumNnDDl1Xuydqo/YJ5OU+jC0v9nmKM8FVDF4VRJq4OeldFC
rnfcvn4Q9Met+tlczfIQpWMBqzCndu7456CzCvpvZ51G1XcnQyc9tX3ATEuux2+l
h/dYyOJ1eUrwr7XzyOUO8f/YT1wMTSYncXEEPW8LZpBaGKCBKpcBAVXNYQMbodBG
CeqCWNkrn9AeCz4nSPzxQsGtxXU8lTZwDoGPZQ0RRaf5ohNWOgZi3AZw2Vn/6tpY
sbJionln2bRjsrHItpTjKdSU6oX6JpWqAKFdKgu2tfbM8ajrsL92JGwAuwiE8J+k
8FiZEXVnaPuLaNscz7K0gZv697wfwZL56LQ22F0XZbYcJrPs5z/tngYb3t3R77vF
aMCQVwTSfe4BOfGRHnlg/DioxPX8/P5oq2HibPMw5ZxXMrAWXrAfuF3i0/XUqAXL
vATYzqy3m1hJ1sb09CUdm8aSDTkeTAGnVOcBp6WUHtbrvXm5lTVn4OhXQWYeYI/w
bcwKYQ14Gw0T0Lx5n3FbxWbpRCXKrxDhlmRcbbutDcLH6H2vd0qJRjodQg5rlGkJ
eDlJJcJLHBsdKeJO8NKNUOtGWXVXCjqzgPCC/AqPTwOsHWUI0WEt7HTybWC3Y7FA
DcUWW8Au8ZnL4Wl5RU2TWvuscM15wHZMcRjJX27GoX/0rlSMHTTegAwJJ2KW3KN3
CdSw1cxx/rzzoDS5z0XlXtvWGK3RtWgD1m/qM9xzgrwnlNrowaW97qIB6GgTWm3w
vONkbu5bUBdLW2knDZfEZMLmcVnf7/bobNk/4FlIPMBypIXiTgJJAGZiRLgArLbw
pJatUSFn7vH7PLgimKcp8inOuhLpd5Y1kxQIFMEbw+Uxnfan0wkYHBhXdD240ozT
Hka5js9j1Ztvt3pedfiDJrbHh/I/qFkKL94hqEAJVMWt5bzykt9bqRDWhokoi16m
Y7bGxFHNiCgjdnfxpom6ziL4UaJp1bLVrKMGI+cCE31FpzyhWlu0WfKitcSVQyvR
ogeBetTqscBI+9nWoiDkr4/fPAMpthEh6CuzfpJK7hxhtoOBifDXP6i6xQi4GO2y
IadRTqQflAdcRkmVigH18IH5BJALCVWzspjcAe8zFLxwS2DYBBJHSdeesiKbklKx
jRpTObTz51kMwRAxHnC6m/C5tYtK7D/bshqjzQ+FDuUjonhgTGehDgyEF2DKGXvv
653HGSgvhS3wYtT/gXB6Um1tqu6gGptvlrdmToZQqtMzmm+A+54hayUllsIXwyOB
AIZqbvnuEqGTBSroBWxkYZsDg5W5Ntf0VxS7uM3RzyuhhIxX2nrM4lfeqTyDb/Tm
s+zm0Vo9Cf7vcvErx4LGdrckJAaXW1gf6t+aTiEQ1MAXcNOYRHE+1U6fyGnt8/7D
uPAqIU8nbl51U1VxOKBH6roOusBN1vlBYoPuI0i5Ze6e6s483KyuP7uUgtdKprL/
dVefGjwYhkZkzKPAmAqD4olPRrOXJpIu7BgJIqYalBL6dkNMa9jzqpaxtbFjqXHn
fXluvMwcb9aUa/ojCD85opQEbYKSS5f/PjfJynOaq2DCadWrjNhe/kdfnIBJtz39
Os1dNUSUUH2AoD4My4yJ/aru7bXNaL6HM2QyZ3nU5MhywYKTRJWbgWXJBbLDcur2
HYRaZKSThPCAgRKfmHc28x/aoCLhfebR97cynGWV4T2fmJQK3mHl07SC+5q8NN/r
G/aBcV66wsdnzYduz0eONBqNilxTtqBnQ7ueUNYFO+KSspGLosUQWgGWjtGgWd0b
Wg/sCrKoDcRy19mPDaJkqd21rbfbHCgqViPEf9rpsjVsDGojXkgw8YZzq3MltzSm
lIUEIc5MUBulHGo/ZodBCga+6mrvrCM4ioEiys7IqY3viQJW8Jv8g1yQYL2FYfV5
XPShwziO+BN0wsGIxULSKr5+AcIIWIZ3nX8VgMwIlRSHLH16Nuv2dAspneHJK+bn
2/idptXMLVS64n7i9X3W+Ztivk6el2t1ngYUmEJSTKWSb9c++fu79cnJByKZy34H
RzewYyp4K1MX+4yUHrwv1SK34oGNVvt5iO7h+NEopVNPKKzi5OEXt5hcVHORylN5
krMMoZbRM2sh2mQVtbLAQYNsFIun4ogukA2/HX0DiHdqPUhwNWesYf7cSNY0OXG3
usEEqbo/NPVT0DIm/+huu1abhDtnI/iM6QssSxzVKbioMDCfhBEB7Pj4rGQIleOo
vGA5Cxa0K2STsH7D5V5dlcqjkRONtOeVS8Ly81foNNEYv3/sMqhnHD8dAd/n8txK
kKS7tYmhz71o0Smg47Nw1xgbT52DgxHXhLja/m8UL4JjxJTVn/GJlIojpFlhPFz+
KT3/ji4eDzwKy6Uds7zTetaer6XAU6vJlHybDFkMekOxBw3VpNlJjbM+XyubmiPu
aKpyg5KSDaCUaLd9Rsym37zWLQJTznDZrbVBHCGccaBbqP7k5oaIzPUkaROF1/Fe
oU+3LY5zAv9D5JTHAtr7C7r5PgX1gvHv5mXGQk0EEtMdJQjudEAgAzL6CzbVDfPo
IlQ4//xig9H7z5yNrR0WCAgReAo0rYO0A0HqtwEODLSbsqqx9ZOl9JC0e7BgY/hh
XfJOSfOIiX0flUp8KtAx4sEjZugool4xcbzjAs71LqjFeML2uCjoHQmoVHAZoP4g
0Uh06FXcmuHoCbI5TIgFxQb9RTPtYMnhE1ecr5JG7+oSwwOGEnAidsHIg4xc7hbh
YKQrjdCdomhWBMbJODAvQ5mXqaYEuqHdrtZCO0WP3ooMPPVPKuML7DKJcZIbAYUP
5NWSaVG8CRSieF53BCs/nfgrecRT6URn8/BoGiRpB6MDyISvtVA0keJG2m9pd8GS
jMQ+FE1dqCIUHHa/rGmcKj+F0g0wsJhRI7N8sIhm6afxkigV22y2f0q0CQz+NV7Z
Q+SbZybE56jBdK3gO90rpbBTA3q2wsLVMjlquRi3PxfqYuJzo6MBDAfJfh2w4sR1
Eq3y/2MBRQGjqbb9Gh2uRFOOZBqLWclDSD4UgVdUV9QicX124wZh9n4bnMAwR/oz
nRfiEo+u3sStEMkyFOOwu1BQ7JgvczDHnGYXPGmxmXHs+sruoTTwZ4qUpjo+hn9U
gAzOf8u2RhMnETxpVsdFyP4BRc8k9ETBtu+NqF7DgclSfxbRgBYO5mZAhWWfT8Mp
7DMaHLazFti7S71156VQJCmwOOJyR5g7tjV70T1jSM+LG4i4F8gkOdwFiEVL+uoV
elzXgNSN1Gsba6BY4Osy6ebOxdY7DU3Yz6NzHQIDmKOHquyD9XNh/9GLXbIpK6R1
kNLI70OqGDuegUHIuCBzNZPGUo3zGjgHKlKEuVQ3YQSPCHFw5X65YrDEqKJMR5Om
A5/UNeyAYCFsADE0zkcB/j6SM9GgnE3htsCcR58Iy6kot6SaxOQnthCEUos+XJ4Y
+yPuccC/WBHaUA90T1cuOsUGrPgmENMj17rBYW1hzyhs7DZXu+v/LAQ5yKY0nLzh
RWSKouEC1nyM57jhPwkffjtsRRBVstuM5QAddhUhJtnKwUtBViiaqzkvVRO2LWQY
qI4BQQeMODbRW3PP8L8uP+bvsWI0olO57gPu8QpNHRUTrkwA6ekPwjKmyx6vD9Kl
eHmc8S/JeANA4gFs5yLKvVc2nZbnvj2mIKgHIwbN/v+4LcWmAEL1i9Bsw3DGuRNk
fxizt5w9a3DTp0CCU7E3BAr9UNPNNF7DfeZsaWPNm0gXN8BjjFHXrDdPt2dkwznB
FBT+wsasDbxJLF6YmoOwZxClMyDWq4uOEwEj+T1OyIdpAWyLkTMNgH23YLqo5y1s
M51su4EFKoauMTWrB620DuEbOpXg5eW1z530gpUHhZ+IDwdsYg45tn3NNrBOlCbO
cMp33moYRYwyzeNu9y70h+xhGOgpROh7GiQluOlFWReQainQ63fikRJ1tEXiuXWU
Hmq9vFE2y1w0ESUAckDa/g/IpVZJO9vANNTv5dRKr9jKQnVKHZHYzEApNG3kn80M
9bot1Ty+3QG8sTdYe/YoHWOixFJlT9FalZNpfgwl2M0c/q5PhFRavKKzhQl++Sx/
ZdO+QplEXUhHMNzFWnfhBC+xWXwOM9lVr7qt/sXB/AH6YC7c13R4R3z1faj83Y4V
y8JMXlvN7UUameVvCnJ8zAC/IvqoCE7hARYenuH7veiJhho9qm4yqjhmjGUuPqcW
nLZNk8lNGt+tKmYpXRYNZoq1dxfvTpukYICs45TdBA/uu6JAuyvMmF0oBxpYowtd
DZYrGP9lRmo1vLaTvejpwyqAP/PKyafb7dSc+Y22qJqEtrlc+bYKmnd+1eryZDpi
Ayob66jlQi42yPjUh2B+TDhV78zxP7tWKyOhd5SzDL5zGARTp48vYdYYFsUKEAay
EYbKvkJtV9MWuRvkHoQVyAQAcyc9s7aKKUYMA5RUzTv0/R1XsHuKOfkUoylWJ+nH
dwiYgH5Jkt8jPsmIzYIY3x6L0xuB5uJByUk2KTQ0xNy2pdoWUPzKsgFnAsJo7HaO
mwfZX93Yt++k8KjHHM3LIunE3/ILoY96SGgR3OZqmOPb/WvuLGxiGsIDAjRNjJrS
3Lui8QefXbMAB12LTesLkmW9wLyXjTVIgnGGMrb//FsQbtRzE3D4OfOqOVkAzgpF
96FLxK/gggdtdZcpUxSjv9xarHeDQpaIpkEZUh+PTlqdU1HsbRK5JaON77f0Sc1C
7/KjM1DuILBIxIs00MhZvkXyJHX4+Df7BzJZWd6tZ08gsyn0AopBFM81K/O1sojR
laUfvd3rQmXm2QZMCjqXSc07Pc5aj+3zM0f9louKZbWxSZ1vz7B/7ptLpvr1g/3a
qtYcocBSDDUdS3uhBH7XVPy6nH2f8SJ++rA30LGAaLC1HIehhhNV9J6ZsH/Jd+uU
WUsothAITYTUZo/vmpAx3/H5piLUuTNXiYfV36i0ua3cUoT2UISSBGeUh92NbOmX
z74JUqWymAzD+Tb1Sa7idSmuoCk9/YXxnK86yU0kO0Q4ke7FeyBGcWzLAo9VLfkY
n5qB7dIKCbUAwtqprziKLMG3/02pQJu+6GZzyUuiDmnuOTobaHTNz8AfAZUfqx/i
dsxZuy0R7a+YOW+7FRUZEMiipcVKTiD+ynQCrghFCG93WHRCxm/B1zHJwWRsQ5dl
4rc28+QGu+2EV59TFG0sxd60OulKNBYd4MpZjILvVvtOmHQphVXYR579xvAMvJLq
Eyi3KBfK+/5QGwjtdm5eiQnha03ORkNHR2JkXZbsyjSUosRsAlY1dLDRrvjtuYKZ
qgno9O8A0ticdJ++kI8COG8HjIdGa624iAuHthoKjTUgJ1JDeH626xqws0R+fDV6
8qMtE8JwE4YDkBs0CtmnQFdr9Xtgb8whZR/XeK214lEpl46xUtFWCx4ueHMfBCFJ
D93DV7wKmkEsNW6DWjpNXooQP+joX+sdmToRebD31kt4LhXyf9/bYXgn+6Q4DEMh
6XjcBMaDlBfOKJUvYRfU4qMn24GYUBnjEuaRFzOpZgTw52MhjnjsYmiokWQ+cSYw
cQ7PsTc1MtX/aJnO54nj0o1ivT8PwUy+pkpf3D5Lb3TN83GWyD9zuKVoFEczBc28
MoFj/jx6bT+mES8L6m/Bkaxi4Y+kK0LQAIIv8W2kbTo8EE1t3y6b0ToBaPnshdV5
9qsimO2ATmFtCGSdo6IeIRNGe61+1mZKmO6Ia1QHHu883GQxfaTvZsxkh1ZkLAVg
BfkYsb/aFfh6QOiN+1DxXNRaq9oleERVk17iNJ84DS+q2HopirjZaPLovL2E+IL/
z6ouAq399eN7QyQrEz2tz77PaJTV++vFppWsiZcBptPgsbI41eY9chJ2wNaUbBx9
VzaulKnv5xIuLO3uf8BhVBZVS5Yfax9KxBHqQ0Mun1BGmYSH3mwy2wAY58AZqMZg
TylCaqQNDA2gh4D0SqG8p9Stb7dve2+cj9fhysdujf8Q4pZgfS7k+SNDgzKk+Yyz
rX7vRj6snGf8DDrXNSX/OM3losWN3K4cQ8qJQWsJl8f2pCulz3xCe+N+rDYzHS8R
+HSRBesqyuhU0ZesGo0CynAvpmUl5SI1pHr/0cZMQUU0ypeQJdcO8NkOTS36pk6R
Eah5fb/YTyoom37HEhlxU+GlFA31lFlpJHQ9t8jzg88T5zDzOldBvmq3735f1wUd
qMdAnMTfvBE3crxtPgNIB0Zru7d8AOJw8vUuGu2KV026xot6wNojrp/vVgc4/USe
blgbPS6C4YFkfdkVcBcCoOWEKv/cvD+/tzs45aXE5a/ocNYfHIoLgQfbU60DSaiS
9U2JaecEK6Efa1ulao5ADllz8Fnu5KF38SfXMiuAM1DEAMAAtKxPPSq4X4pb7N2Q
vDgxZm6HRHdWrZWLQUpILp3jq9RIlbXGzw+UaVXDMzD3uhM5eOvESpCXbkk+B1G/
1lbvf1Yj5EGpmnjUsXXpeqwmXoFapmvvwTc5TtqI6tDmCzP8lejwmuH8P40wkUGr
oA4ZGejtE12/cGZTLHtVRji/K16+88NGLIemd7cTZsvAi+yw3pZLiB1gMJDwhEMz
vEtQrHyr/qDG9/6Vl8ZiNj6BvrC4MneeKnF786ZDsP/6rq3U5g4X4tS5Punt4SU0
dVNwC6MApY6XkG9lUuDty9bi4nP83JRJI5zVzCht0L35dJwuY/OzkEDlsv71piFf
7IVMJ3RT8tEm3agp5jZos9Kr9gzUKEFAZx5ZlESwgeNh4pDMry88LxC1vKUnHybx
9ePfX0KonBSKqfUqdKB6dMdGQRKhsPXzN6mfRy4ioZDyztuz6Wj2p0o1Bp8sKs3B
ypLUZO++EkGwj1lfie7wtPopVrbynOfyOHrNHOck9u0zGUr/ZoE3nIsOHRRsHtNz
I+iJ6vd5uQz1kz1qc8Btk/+GjQQFVG2zkED7ZSR1m/t00kYG/3MdXnzo2vq2gtme
LfL4n9w6dg6TIGXLS4yo6gYv3tIDTSyIQftdK8wwPXaJ56vJhTWTaIZ6qg+T1mMJ
Hl2KbF/sOQuAeA3C9R68ETBWkRa5HA47bdNK17hle8iICVJLgc/YcsjpOMBT+OLm
s7XVKdyRYQqbZ2VWMVzet6DENpfrMnpRvbrU4ayIvAlj8oabvogDhOcFiNvx4AEt
c5vv5oO9I22nw/kKSf6u+Qm2q5lRw8bgmgNI4WZK5xcADHxUo01KUBLvK54rMWfA
hx3olwKjsfP5zYYl32BFQT2g0mq0Spb4ljkTZotA9/MH+0uiEh6UE1lcwh6sftGM
XTykd9KsWUNmwKuu6q3lqVAfHnbwbvqtfu67hgdF31N4trA8FVgpT2NhWpCnmgyj
XzmXmXT/XGGNpnT+geN9UYiKSDt/22bPP3MOdharW7qccZ66ZoDk02P4IeCJF8cI
pIsFJr4vgshMLlUc/vhxjCm/Ebzi5onLSei5rlxfxOtSHuQZHJ4BriZ8SEiBTE3v
S5dv2e5igPP6LsNFuwPTQOysGWoqAtHVAeCSPi4C5Z7mRo79BqMbbdpPDtwVM3ZJ
OBhIupPKKssgPSLPDoIJedq8efIEUK0WA3NZpTJ5wXpAiTBhS4JbShfhfeWl3Y0n
rxq7gdIMJnPqxcchoXtQ8O4RBsRaScbQ6iR+5GTomw2+RLpG8ket9GYTyW0LLGUe
83nImaZZqpS12Jrabnum9AQnJnvVuCjt6FWnhc6XolkD1zzPXpEhHN/hQ2Xg4Pb9
V6Pw9bkwSBjtHHvU1zRln0bzCaAUFRSsMOoBaV9FjMHA8sX6Qz5CR4y3wRbNjAjP
pFr33Lzf4pExnzlcwmfdpGP2q03R5Av072+DnvqNRsm5wQgSByNqA1cAPfFOyN4q
pxnIjz6kWIeHgGhLoRkhIui52FowzjTpDCA9JtrUvtvdQ9HhmRppb5+hAHRtO3tl
WScqnMUb3fySXzBmpWwAduccUNNdt8psiSKhLuhRVNqI2Sk2TcsiY9je862xxgWU
Sg2FphRqKH5jgHvo7IqeyuVPl2e8uRk/HmIDMdHao+Hq6A0eY4Z9sCmOhk50sE5E
Efk0BOKoPpRWAwgjYLSwW9T0YDEMccIZg9UGIyb3MAQyj0HXwf4wq3A9bLubBaV4
d8Hoi9VjjAYfSXHBz91yAZ6qiXacxACQgIJU2OtgrdaKQyteElHmknNwTjkfeunj
ucEBeHflPxy8ZDYVSfXO80wS+bT/VTjVrYPnvO5OO3uF008kiKdRorQMW5Lw2/F/
llHq36E/rRzoRB5WtVTaE3I2mivpGk90mTVmIfk+tMw5/ecqfB95Ya6B5N0HStsn
NsssNl7e2ZBAAweo1rSW1/atWSBoccYF47Bg0tS+6I8BHn8aFfogF5DzZwK3G4tc
XZgFjURWfoR5ozoDXniEJOCuy6dLp887MhO+znvb+Mh0SwDy4spyFbU7rHXEG2QF
v/ROd3IvCC5TRpR9/EoEGxhhhdhQignmIM3/7GmSbdtClyaYG3WCOBS1CkfYvSLp
ijxLylsJsjO0HzNNmLhCaX+qH4GgfOCZmJwHAEBvcuM3RNHJwwCGhUHPWk4mXivm
vAGaGESrlhuQ9/lTt/hza60Iz0iUI1gXZH5pKFkvhdYWIm5UJKLLAvc+j9Rz3u7U
PRBDQasuFkUOv44zi2tBVWvTH6Hy078dc9oxGQXBfXcMMc5OrZocCy/wKoJSaQ4v
DfsA4X6vUumBBVS9Nmh2N/F5a/IPd0EX51u1rk0KUGi9LMKCm1S1DT0+VThe5fOk
e/unLUkNYZ9vo/J8WeTaCQGN+FgT2RK1UY9UE0Y6z8qWq+op6FmvpCkomyQ8ZM6O
XTpul98sKEJQf4SQ8+aFqy0wAj6mbgKYi0dn3TTIGg5jOULKrp+62qLZfbgIbizk
sUC9Bs6KF3lMGVrSx1UnpJKQC8OLyXjqVsUsXqOvpPRYn4pCOLPQqChVHTwH/qZN
ucMfXDJppZrAxOwdM72lQY229FR1lmxIWwWDu0sOmLLLzeK+dDVGhz2iUeNjutRr
hZ6ofeFluE+SKJaRlWiFtxeAXMUgUherJIZsC7wbuf1HrOeWV8+xZoVOqK3lVJU7
vINA5GOOYGd3yX4F1Kpm6zTEQ+XKF+2nGcD4QzbsilORvbghsf022WmLILXYnc6d
gBZtal3hurTOX/8Wxj/GmMnLFZNNtkXJwfuCFjp5WPsViMoDW07FNLJsMxNTLGof
ImEKblmkDdl2T2UlkELYoZ6lNU0YuW7f9Leld+OARnjqeJZhCbpGFYRWpLbErFrt
5qnt6+P7n/eDlbuk4u0mXvhdmFSUKDvhAW+zKXlP9IKnoW7d8nF3y0bP6ppO9XmH
5whTNiZ8DindJ/du9mMEMrToaWinOb4HPK875ZPIEHF2vARm1pHm6dPD2hHQLcKB
MJhzHE1tjmmZRDI1N7Dxg2JfHSeXH7VleJV9vcyPwhX3F6jO7J4P8aQd8n4TC0uA
ujI+HU8xdPpGmoTl//jSeWCnV4xYjOytxA4crqljtaZqfn5YIfyayX69wPSG0L02
t+QdP9b7vmykTNUBE4Z26WMUWf4ZNyBRav85jZvWKiKqNBfVSauT7KSA932H/mlZ
rASsJTv/kt1586zSOw0unY7RENqYXMcw3FI714gZKcS21yvbRQYURZK97ThjEgTR
JQcG7pbQVKkFLnHWwey/8SUxX75HtqJu/N8JMP6jwJ6W2SKMvla9uZ5+d8Lmpjhl
F0SBoXEBc97yRgq9q375f74BRtjI3Bd9CQWn8Y7xCYpufMAMuKJzBAlc+EcmkVHR
MQjnqXo+1GN8DWmtgOoousWQ33OnUQIa+hp3F3wUkkp1xE9KlxSr77CsVxTADmPT
mRI0NGduWKGs/olfVmtDPuIamfyoJ1TIleH9FlH9qLTH/i6n5kfbrx8Xy0SiREpl
6c95UnP+LjCDxhWvruMgyBdz/A7HLM7I+LuQeNGUIHJrhbT3K7OeIA/Ok8OH6wr1
KuWm/1fOnIPi2kmphlipbN5tSuJa9nBTS9NReeiRpk+X7AFMocR94B3f3ZpT9JLz
x9OrP7rPDJ0prxRbBghE5wQqfRnfNVPTV2CtdjWUCZCAeNFnJtwt7Ao22lKTK0gv
wQq3BaHvZvkxr43YoeM63H6TP5WRfQAeZ5aHJsf4lUNh6VqzV96oRFD/s7DbERUJ
+Tzl7VC9W481yXT/AjV1N4vQTKijliwwf19qV2StHuC/tC/FCFnbKoKyf4HY8jnE
4o3xAbX78CG9v24pOYCzjMk/Y6Z0NR2faCDOFQl2xfG/BpegZ6mOYHtKm5p3tSLB
wVuL9dxNngB5Wqbo9lM5ZRVhUVni4hBvcD8mAO4le/bwB945gZEy6HPo85JzjnuL
O8qR3E7pOMJTDJsdm/a0rOWJWtEworBvcP23I1k3VIHqgDBrGZlPgKOzIEpxe16Z
SaJ+Uj7kxYXmz1qfD1qEf/UrX8cfMPYm9Yuqo6LnyqHumhNQKPKPPo8jWBRMjoHh
kGFDId3W4t8M+LD6krEAPW4L8dFLEhtzd1Mr4izipceTPISd7ZH/dAPuFl+36xkX
krOjfjtseuRLxccdECaH2K+zkZMKYRcKEtssS/+GS5dxOhhJG0zMVBfyLwPnOsnI
nvRgtcUj6UuPffniZD/XFCnvzXv9rxl/c+c8RNM1sNkSP8xtMj/xVBnjtLXpnNBz
0TuU+lLNik1kDYURStzVMrYphJQAstPSLdW5IOyRQkjFMq+hki+0S5/jBUnoGvDz
h3GfXl/+Y2v3nz6eRDrpGJxz9RhUduEsde1Pne9PYmQy9EF1knDkkOC4neIuVxis
uhV5njwHZuUUOBu63AiuO5KlqWaOh6EIGfeaV16YeloZhCdO+zX70z2/xevCs+Yl
xuI7VIElX/XDbqoSUesrjGzxOXmWQjoz7d+aSK/1/1gDVjIa5/ip68Rn4yhvb/ND
yjv/fenNH5U3u7slTI5/+pmrXooUuOLAodV3zud67dJ3QZzTS+I6zJClf7y03x2Q
9nMrFrKslhnrbQxzS6LDXSWLhdFJVJlk85TWzbdLzV5+q02C1IcGyYiBVb5egv76
rYDNQWJgRmtNqutSKg2DP/ahmnoI2n8pqy4hdFW91WVWpGHVOAoVMFlcQBeuInwj
fGd/IgTEAnlPRNGCpMIbvelVUpA26Frd7wJ08aJbatOF49oYCtwbDffhXA1B4Cwe
YPmE0iJtWSJmFiI4QAtSZ9aHnDP0QHrVCOtHMfYtcRaiHBQ87PGedRn3Dxdkxz0T
Tzhg47N/ZvRgpvGqb/dEex+zmgLt75ql9Z3/uU91L+MjAHguHREBGB+AzZcYprVq
0U8/3DmJppDY7xiqAXXL4945vGwx0hzuR0mQ6OP/jtHWzCDPNRzI0yXcVTKdVcbM
WTV3n1gW/k1Xg6pVeidXEud/IAdwSA6i50/SAjZI7XWgnqJUD1QFj34q9gg5droV
lD1e52+9wS72W0sv86pD+fW5tBLIDmI2nB8qBsHNp5xGHR2U8fxQG7MlQWASr/qb
xHt5/XKvGZueIos7bPSdFUd97UBhCw3wilmYGiqjlOGn0N4GjcLtIUaXDecTTlJc
/jND17pgYXrzGLGJXFQBL03lzk2Q+6n3H3RWsaHSUz+whJQ726ZPp+uPdOIluN4t
A3Cuqk33KwmQimFav5K2y3cCjwrZwrOqclb8Q4XcFN/gETJ9U4yWcEHNcVocgn04
kp+V9MQTDWsvAiDm+fjVZaP5EZTyDRh25obuMtmcEwyop8BFqMDUX7U9Hn69g+nD
Ba7Lq4y2xJqrKxfn2ZCc/nEStCnaqW5mogaB96dcXsS7qGFZrD83S8L1CNrwqMzq
r3BUhlKmLu7w7BjsbJZR8/m3Bm8VlGRJLLSxvYkTN8xgXaFH0YM4auE3Cifdo51s
Lt9NbZc9yLJmB7xFtok04nbH1OOY5cc1jk+LmBZQqmljAQ/EKRXD4lY6iWeoVpdR
f6kdW7c4NKIUFDJ+tfOCkrkfNIQzbddeYr9hRtjMoS4U1gF+p9luN0y5T4P2qqOT
W5uPuHma2a6sJgTH5PGTSDTlbaS/tugMzTyyvvvbYqh1tdUFxp/Sn0jzcdD2mS2b
9uRQd6EZtGmWZUGTFQrfjfwVN4ZwercDUVzKT6/Xhepyv1WtP1q81piY8FkJQaYu
W16NQDVS7NYx69UGGax8974TYxfNCN1HAISluzv8EE+MQdnv5+VG7xaqUZWw1Mwd
Psx/Ha7+Xg/inCo0VzOvR5u2DhqrDfUni6eD2R51m71h3SRbrolyCxJUYlRUKDv1
Zg4Luj0r0tFMC+izM1EEhJton1cfZGwR2WVqQPcXw+a+URZNG2Ee58D2kKu5Iw7y
ZwFpaGyr6/KxMiTTMKb1giP4bIm1KdvOuTAjSBizOIV4AG7xlh8MdZMF/zzWdXuA
l7P1ZOnAg1rtGi6ZEkMkI/Xg/hbNYEOcFq3uQQhYIO6aQGOLyJe9azLXSZlIhDW6
CAkafs4OKkF9j1GD9oWbbrp/bTUAInZj3gjM7okD6CKKgD3nQ5Vd+nZ0x29TNmGh
eip6hB2GJJl/+HTBIWGzdJ/hWTlH4trFXbgMxS/8gIxArrGMKFvzi/WQHPpQ/YhV
MGrrFcDLqliepnJoe92lAWKMxDveAkC7L9R8JCrMliCxoiXAPVknkkPJFNn1bSZE
1oUllemhn9aEfUyNyV/w5Wf4EM4kpIPzKi4OJBxzgNVNftcp5bbzWrSzFLIvIdtI
gfpsp/LXok1Uqsb3iE/guv7UmlzbBvhwa4gQ5yBGhzdriqaAa06J1phv5W/q37gM
YK+9xTx1NnXj5KtaOIFAyesrovZH/JwPohKizvbsQQcDlReHkcAZVjgy5nH9+kUE
EiL1GYDlkC7R5n/9nmMQ3ousOMHpuJ6vVg2JXAKlcl7jLWTbxWi8h6OmWULgJw1K
6gF/VR+eS/WlTQIZSXiIbIafTRiKVfGQuia/VMx25cVT4hLytTX2iv8NB4rj5BPY
t0JBdCCsDoIdV0IFG8YA90eFqAk1BSShuGgxDv6fCHbrF7nMKQRgXJkTUS9gwVer
9KB6ITk6Vo5Z5KTTMXISk7XIEvQgpI6bBNyYXg6Alj0u6ikqmQzdVurelCzMv62+
0tw3Sqrs97SGoFvXMTp9z78xaS5C886gnGblBFOYdqIU0BT3vk/L/cHzpNCDzt32
vYoGScYxD7wY9ZS1akyoxWJWz0MDwaGLQMNeynuZg8LIQuQJvgvhRSIr9xa31owY
H2nBFyfiD+MIpIXq1ZB8ydHn1Cks5ZTPw8X8z0VdoxPgH0n4AbtVeBKCEBZNGj/G
693mIeeuHmfWJl2QlLV5m08quOV05nS5Aa/YNk9zEzU+xwBrcz0zkiPRBc2d/kEo
v9y294mjWkoBYCl5E7ZAFCtT97Gt8W0Vh7dAOyvRqYOofSAZ5LS4/6c5W/hMt2Yi
MYDnGLrOYboeJBOcIdUnuuxbQGPwz+N0Gkk9XHvQ7eUloDXZBbDAJZO/RYdSIR5U
41/2+JaHCKpPRlgqPlqgvxVtsVW6BwA61EydCufOpsXBN6bWqYkxxLFcW976WH2s
XbSTKnAsHDSo5GeXXvnPXDzIrrJN3eWX0zEO1fWaqRVhBAXGR0zMapHTzAlIU9ol
7ieiG4y+7JCV1qPGHM7zUtI19m4s3DgPT2yxJn31aAJIjQeaKevAynZJ43hUh9kK
TPWJk+JrFJ28KyP+v4hbqTMbUw2Rs2X7yGyS5lhv/OfAWaAb0eeeZ9qQrsmdzvlX
ftBnP1dEJhfoTL6BRSJ7Q2ogFUK+xPIbfL7krwvGt/B5sHDdURNqixll5fseXzKg
Ws4OJfXVTRuii8FTXV4m//4OsidfDuq7WTI/JbRhPAr/O4iKCGvTjJ1vYnDvK25B
P/k+EhookrK1oYMWAS9Ov+EOmJHhqmLmKVW4ysiaE9GBJomjBKOpGEbsRXQ/zK5F
+IN2s1FzGi91YReoxz9zHOzHyuYF5hAu2iFb1Nap649sALBQjJWOaB2QUAQkzvy7
9mPzbEMB3OLvVPJxkBeKjT4dlt5MNCe/meMgqMw65/aFc3XPpWOeO5AG4PrKFo1y
VcpCAmQlR8mS+SgTCBnA5+t7UBwfiuUDLSypvU+99Dn8EzNMwhtXBlY/qu63FgQi
aqlfL1tQCJPZNDuKF8DYIlxErLyI3WHLkovZfkKaDIt0wBz39mM9lmJD4em6bsaU
hEK1C/ajLm4z+KtloX6NyNDwCp9/sCkhCiGCx5ZHt+j2yF65GfPIIJVqAxSSUrvC
dMezcIsg0j2ocj/qNTJaB+AhsZHsfhLcNihKVAuiCATbQOGM7bE/H1cSyogL1co5
DurRLVy7P8zf9ktqfcgS491P2hFEzDJBkzOJ92okDZdgPTYPvALxHcvaKDSjAkTV
Qe0Fct7VbD4xjLJzEM9BzaMg/pHxRHIwYlmdIce8/EOfl8pQ+nQd6uFewNzh09iS
ZL37NxbRdfHFXVeRPxkMcc/YSNNceytnsUU3VPSIbHxnKBK/McRm8vzoa8pdypEN
0wKSqyxqi8gXNUbCiuppkjaH6nWfFyaaoLiwyi3PtsaNASx5X0kyqccbF7UBVc7D
zumuX11yMu7ECkRvSYVZKfiPaUEDaMTSJ2GQdub2Q6WlpxvTGS/nNobW5ZisEWyT
D2qnwy1+MGgK8KsT9qK/KKB6qzx920l3udDViwKQ06h8C7kNg/esj/jnOS8KAAG6
goBPvBziVvNf5r7wBr3ErsNYcDkpzkB6Gx/xwE3mTb37g07XeLfJ6vZTzydDXncl
M9Eh+gCU3mtgeS9YB3bm/sfgu6Y2kTUlRyZ789fHIjCaYAC6QgWDNDEkiU3NGbuT
NbhnLSLSjdInlQDvVw6wkgHMuIb9wvdRiNZyAd/qHikN/mo5yvJatEZlj6QaVFCK
ue9krkVuC43M3/QcBFq0Z3reHeUonHsoniqajubiCPkEgxAV2Mj+B+uzi+VAnRAl
LE69jsdGSLNRc3sEjVDV1gBbVS7gtVb8kAtHY0tsvNa5baKmOCnSByW75cxq1DJX
A4ABpm33rIiaqP99/bTLVl48k5XwsNNVUTx13bLcs6u2k3RTea9Hf+hRkms6W/IV
9A//5xQc8wwcU27hBjhy5q6YJid4QhIv2YwHOBSnDSm09a4YNuvP/KhH/P1Om0RR
8+/SoQRH03kIpAqOA8TwUZloi117yjlbaiBVr4pTYB/0ttmrdHDbWHiTkcEDye8d
kdGMIxH0SYUYOXq2V7SFJ9ze8mPthzFETROTvxZJu7GxCJMUnOM1s+DMeO7qyjOj
zlDMdPFsGL3uyMItQmqyRf8EfTmAIf4rT3RRR/JVF87QA1jRCXVM25/kTUFN2n//
213n2nOrIA8AlwuLlSTPgtDXBkXs7Ce2mX1nbLD4jVMjhXhx5PE0szqe5y3HWWCF
/bURv3sF5lLPp+gwgkEdsKOnGyR0uRsU4zFitta4BxWQM4Ex/oaoHyAPGnx2e8qA
frV0J1BdfCY7JETnY58YrKcPjA3V8/vIfnOxQ3ZAeUhltiKnkAAX6DRkCqFhS7Sc
0xpeaGlQyJDEtwZw1uL/U7+2M8aFRhLQcmb1mvfN0ULkQ3FzADEHXhnDN3yVBNQO
EwNSF1cLGP2jq+SPdWrCTSr0p7A3l/5xHYGWQbKMdynsRiBzjxzZ2S5onbLegxfb
qH0IsgqSSpaNnZd4JBoid5QQ8RwLNoEFBWfWAgAsw1DUdWaOafrU6aRawGE9wwst
mjpy3jxqDinOFtBWdS30yJGE1fCntKgsnzIV+FFw/LXKUuPbgouDzn4NIHP1Cya6
PerGquQAlUMo9cQZV3ZjqOWDcugAI3vfYsdJ/2wDrJ91ruW3+edLnFrJ86JQCO/0
9+Rne9Y1BEgwcRI7EOIROfihF7JJh4loqJl8BMeA0WGiJljf2J1H+hRnuXC4X5L4
fNV/oN+Qb75yXpd9Q2aSf3tfoNnhUpbYwlJvS5XC42iLI2uA4SmPegfqBDjamgcQ
zFoG6RY0kdlNIWM0NTm1muCfUfE2jmEwbNY/VfAgIWGWUh6sN1ip9DdGsoqogmR3
qQmzziua6byjJJzLmU/55TwbRdn73usiiZCVP5o6IbWANDY/2M27kw/9yD1Z5vam
jIAN4EmMoGCrgIjtn8jM39ACygUBdHxDpU+lek5FcstIu9ByyTDcCWDyJWadAkpg
B/KxAl/BkRwIpgbUNeO5jfoqKODGUWlKoLC3NIarWQGDZyjEBm2D1G9SnDacLee4
MZv8V/jsdVA1XVGvf4B4DWRkNDz5rhg4QmngUA5UkQBRx3H0fP8o1ocLliUdl+Tv
QQmexsTBLpyujaxXd1LzZrbJMRtha7V2gorrGn1LnpObf6w9sxWf6KmMx0Zyt5hA
CJzEDDK25jaw+/DwM6fvOHrkdnqMdkRlWnDOLOWyDB0SAQRrGb4B8zh8Xl8/IwRD
Zu/TcQK7wuucwmwBNtH0HspBVsMGBSbAhvvzmELT7PFrjmWthj8LoWZM2Donr2Nc
81b7on2oGWPi7yTLEzKENF2N5hcYgFjG/hRknIJv2R0fsA8RtkOuOLcPeRoXXsLC
o3fH5empwbcmva6bgSvgvUVafTaMNEl5ITFGBWRSeiSvodIZ3gFhd4jGuQnkRuq2
L1WtGnAYky0+u9JrwNmLrCkKZuJMc/2zrfurTJJ1KU7iaLUt7KDmSh1AO4++CkgU
TPSFaE+vfUKB1e2wHoiwYwwciI3wp00T+4rp5Mz3lrUaNztz9hQfIjXCm4ih7dzQ
Dl9rvyRoiyhW7Zrvi5qgqR+IlZZpMzJdW8VVj7AcBPiTJYt1KJrTOaDrQiKaR65M
uqYWnLt2M/FER562fCva+1gnbxDnmFaxrT4b4DYnp9yJBaa+r9oTfQpPYyyYphmC
9uyYzB80Nvo+heDMdJiSf3mg6S5sfD6QmVkuHSQbdrsDtRqFzHqbY2pSMDv/zzZf
4Vgt8SODThuZOod0Twy1Yg8NvzrMVb5Fp1xzR+gjyDW9lfcGj4yc1NEZzYvmGnHA
i5kGSttPKIYcgrEnMFTXnw4kbtpRpnDl6QgTOU46DlQuAQY4/WfoZCgczp+n71JM
ACE4spEoWoCRY1zriejuKI9tXHRrQBOhvppyB6tNk9HFTl7Iny/ufMtRT8eNd/cT
rCJDHLgjiNEPiCHb9/Lo3AuV/iV5P4BHyRQYNKI1WHDRH3AbbUb0PYwNdtttRGPM
2nrv0HaXbOg5b0evsKeg5nA/7ThK1fBef+xycDGvMPVFK5PPU486ubIf3NIYTJga
QLoqqbf1fuomBYj+NDYauDkXaP19hFqg3Cs5GTfa5DOxC/T/HOVIUZMV8ICkzr2D
TGVzoNDUOxli6j0rxReRwcIohI8nL5GnkslFDIuIDhKo3oD+01HdORiAuD9C6Y8c
AOczIlDyIbpP4R3WGBv2ivKuHwl5TIDhWdaIQTD9zC3I2WYqLhF/G5zfYjvrXPYi
+5W7c5VvrmMWvnbmMM3HLjRURB52gAfiMBIImbRkvNU4BTk80rv/QZb6+zwoQ91m
3ovBo8MOb7QstvMD06085Btx47peao6jM6N6RQ8/zdKTz3rkeHiSXosqVLHVdtAU
kTLCcqrvxegyMJdidYVccVveAYH5BQCSywbtn7iXg0PhbozaGfKcq0rWGfw7Vo8W
S939uhtlpkRtf5WO5Wzlg9fUANPNRnYyg3luYN0vnlQfnLmkCmvMuPxXlS0VleaC
oxt22IFcxYIkLZ54MrSO3cBkPbhxJhlOLNVMjc1FAslDtylbGseaApcLswb+hmt3
2RedoXpucNdSpecHMXjCZJyf0IHSudeiuJbMJuR614AiBYAOLc5QmG1pHJkab8i5
VB+r9qhPAL6Rqfo8MLAImfo1rNywPcTXCxlWyq9KwUV9R2fLiPKXfOPUP6EgWcFW
nXEAj4iXgZSzeV+EGM1gzpobsc5cFZXpvcrCPjTXAEgmgAaT51lE2yxg4Dl3dl9w
RpkT45mxZim97ntK0mQHJsftdjo/5uz5xlNqT9+paB2r0DzPtxA7UvCXbtDNAf5Q
4zKwQUlvD5WSZ+sPT03KGihCd/UCNxNhL+npdO2gTM4BO9kBP7gwiNOrrfL4GAXm
rpPk/egyhX4lvoSYqv09AYEfIXG7qAQb5ZWlNq76tErHc7HCbbSX2spej+tvXVZe
LR9cIXO7O0giMoCCXkpUxC/yoSVNu/gPbuDx5f+6wqYI6ovfhtaiId6Zc6GoaKrv
QsrI6LNtUMwtwgBOMnidAhzelr8HmkRjHpR3gbNbJOkug7oHzo2DMnsNuphwxdoM
Ybyncreai8XNVHHP/laobmmYb4i4R9Yabr4KuviZykf20BZai/LqG25P9kJzFWy0
qq/NXLuEYE71Wp6KGVr+CePXb6NhTr81hrLRYtZPm6cDJa5Y8IFMcZKuaoLbR6Ee
96ABltNqPCAOTi82t2sOi9h/5OAR2BrvTxj2JNzTaaMYLmB+70fmYXe0mIpasGSQ
DNxGVkCyn9sh4iETfDJ5qKIAtaQsJCN75po2wxpzTEFT7Fa5LYhAZIG4G4Z3h3HF
hAkM3Q0XcAWpIqIcDwiyujzW30Bv+KhE2vCepMH+NMsPJ/It6ioja9iSVqkCyJ6C
uPfaLBvw9zK0JzE9Bgnrcu28vWARbl7y+34TohZZSgvU00lMUJF/nvZNLxh+o0Cw
QMVCPSIoJHtypaLFz+fiz0ofRGS6aFsMPiEnJS46ZDV7jbgKCltihjDJAtsHv+fw
XzyTKi+D/nzjkRUSg4OGgVTR5BQHg47/ZTzwZaCO6SzDUnnm4ckjlRzGzihzCcWj
qUX8bwPgU/q8O2MsBTkfjjEEKLnT5IPN0Y3jheRu/778Z0W6VH3H5L5zfPwgMu1p
dL/Qr7dx/3QVzrR0ZhX9EDrpMzxZPCWMf2TlGAYRKTAgAp8pi8iKReu2zjEEnZZq
iQMmlvgyKWae6Vsq9criX2XTLjpV9Dk97wRArKCP5R5dO18dCoj8SFfVg0x9zsIu
mfLjuA/CjXZiNNQgmCChiqxpzaPwj8geay/6bNK7qikTxiLnDLC1LxEnALDzY3s9
yPUuRN06RR+qjeMbxICCHOI1UOxxovoJFQkZm36BfslSuV65jvEGWMlfchK3mknT
C6eXt4Ynw7BUJhf3tNnTYmfawe3b1bDdH0Qzq4SIjXX0HG2zE6KkuogLpI9RdGPj
mSsHZQ6FkAtbNZkX5bMwlZuWYkV8F4k6/vQ+nAVxew1fQ7XIQCnpA0IcZ/RzEYtz
pU5/TlAP62otmmkzyd1qs3uYY1R5LigX7/9I/HSh0z9A3TCK+FhAc3qDcALItrSs
aSMKfobRlI0AGTgoL1qojIvHeyqNhi6vJiu4gzKnlsQvSQ7D7JxLH4wKE1G6nJDL
Ixe+rddhPj7n04cLFzVKjJUgUYoIlzQat+ydMINf8VcHpoL0b4J7qBTWxQLpGxYs
eDlo/XepKaWTvCsdAOHvGfTcLTLjihU86F9FPcZh5pZtqza3sV9am4y9XyV2JTAa
EBVg702B3GuWngoOaEHNCzWNy0up/mn859IDz+VvElHgyyG7MKvfGnF2Ykkn5rtg
gAAMlpPu5TmBVrndNBLY5DFGd1rhgHMp4+tGQ5CnYIAV5lZgNvIbS9zwy/5CJ5we
oM2mPybN90viEQbT4EBKKJv+6PFRhvwmHyL32UP8bxjeRtQ1K2T+yMyftC8m90Jg
AZS6lAJgl+x8H0fjJi5J6yTifqDPCsDVtZ6s3Y3wt0ToAvOGEL1aRzcV0rgc15o3
oLXFyCdovqJCmj/b+mJZ+9ZW/w1oxsrirdY4utdO8+Q3wvPoQI6tZDsE5LcoHQty
h1/tcQ+ajEHiLqYVkX8LkNA3t1w8gT8ufJc32bU8H00lSsnvEv66CsdeTYStsBwA
priD42H3aFsVXUf5SzqjF6RhMIbJpDQ76aJsOgAWX30UXvWJ+4mOqcZ2OaxPbuT5
/hRlkQCmkxCVc9zKmKkK26Lgfz0yIL+Mqoo7INs4QRt9RYFTGWukOrH2X0QDnnCT
fjDgmjhkuQXexZSNFs5+Ia/GR+NbevNIMyypkLzbBLvwbiwRtL5BV1qtJyNVuknu
mD2GEqL1KN4Gim1r5b1CBnUh/5EL4UzQIb+EB5MBS4RpHOUPTa2ayA9qh44yp032
j1XmS201i0V5CcPCRGdX8JWINKLQT3w2VOi9beNjAbFsQ3KfnlpOSOggseF6gflN
iNKw0tZavT5gns6yx1JfCSlWP8TyZghTw4kbL9gYvj/XrfcMpzogXzJSb7odGafO
99jU3WA2XveD+GEd/mHGRuRDnMtGweDNc/iboQQ9wlIOu09lf3TIaKTbU+5jQ4zL
4FrnXHGh6uPa1OBb+d12lzWGQc5WN4IeBzkiMsPRZiBvyFDAOhapysv6SmTsBmoH
Ljta6Sdp4EgRR7+Qd+yh7lnc1u6+DDnF/ocMA4FAYMxmrmcPfk7eV3yOSzaxd2qT
1vsGjdKZuX44EjP+fMioaVZSR60eE43pMftKihtu/cMAljZDJ65/u9+zC77V+OWt
SWL8o4Kgr7nc0+OeR6UZ1nrrifsEeQTEB354PnSA6nyBPmvdaTgMIPYPMJVNSIED
SHWPIm6hlqdm4QJwjwKb9GFhXukz37fyrkCwkE9G8AyHoEtRk154uBRCR6UBusr7
/W7W97QeX9zEq6V6s6TIvMVIjH+oiyX+raskq1oXwIPVyinWvocp9LV5wd5RF3kB
0fj/M7tJIERjKbTNcoiwUDL2xeR0zspMysBL0mnZinFH5yHdw3lEKtCwDZ5S6e0z
2TFatMSiv4m8LEQhQl2AZNoVGwHruWqxU29fQ/22ZTsBLlQcHnG5MPnPi65yGUto
OI4NM1dTbPxRIG+0h1+EZP/Wl1OUgArZY3Qaak8mUpGQHAPNOlEv657unkBERJf6
f/zmAcngNVZxiv5FpE7GYtoR3LD6J0SuuW6ma+rb4gU0ll1a7wBlxOapAw+7ZiEj
GdxDODxZZ5ruYGqaeCEpq/HhAsA2kpSbkfzD3ZACWC/HuvYqF55Eoc5CQ4OcZ5zF
18KQicU/Mms2hi0Dq2mtFqbWQ80OvPoDcXatufeW1FKJ91gm6YLVaERNdm8sxalm
YTeQODD45IOnLKRhDiBKvi+HXKkAmAP1gFNrVRUIFmjz8H3PyKPH20oxBS4K9cIl
QmL2a1+s1W3Xepl2nbu04D4UauwUcMhCDQhjgIQxZ6nU1ooZG0pxWtEKsxeklJIP
lWRiLgi8imwyafhFclTN+IxPlMpoylxCIvsdNRS7eOozkXyf4/S06LtYy2u/xM9U
igoU5rjTb5W9oriXrrDfvmFTaktmxVqD6XH+lr3HK9DIpbfCCqJE9hIGqsytihdZ
dIeoLaVBfBh/b3iliejS1KgB5LjMLZgKA4nQezeU6sVhBMd9eY0ndymqAPaQSB7s
PrVNbUzD4USCdgiwEY5H4ZlueztClqFN2IyIKPTCx1x1NgNbGAAMOzMffOT3qXob
fuwlUyi+l8vy7eoQJFYJctbR1WEE9aCh+zI+47RuUZle1H/AayALtS2fXMb8S3MM
EIYxZB8uZeVsW3eVxoheSLJD9zmW3tmzcqHdk9Qln3jRpL4TPuAz+92aArlqmI/r
NxeHmPt9tfkex2VJorgAKMqp/QARbOMzfm/q53jY48hNnX3NQAOVgfGXBQXpZZi4
DEzay98HIzvv2eUWlGqgdABzqcvPXF8OIEsT9huMQSqwNwtHmMdntyp/5tS0VVjT
P2mkVb2fCvtFddhvFFMsLu9mOhvKwBJ20p7AqOYFtL1bqb3etCrElaEiup+9hbbC
J4tsbF07zjEV9TLWhesX+Cui6Zrx+GnnSxyAQhVYMz/SXc+yOQkYqL0hivhlLGc2
1rxY/cn0DuaMOzZBPGOqsJE054gneX8pikQTJXNZB1jZuWCUQOPvqnl2H/1da2o4
m0dOWpe69tqEnBO6NDQFHhSk+MZ7oybmMQamf7JIO2GkqMS4K+uXhdGP1cT/PdIY
eTSMqagfETICSLqzDBfBmlImRnZF3SYjioSY0zBJaHpbz7u7QX0BzLQx3TVjOZTO
ca6Sr4IIeD+HPfy8AJ45+hRQFdUZBAHdBf6qM2c6vMgzEzgNHQkxjzbcz+WJkSSI
qaZwzHMFcvq0qUOgzNxf9p1vzVl8rMIvDPvaMsQARFDWCz/7zlrdQy4EagV9Laro
xfUcu8yOP0OaYdmig/il0rOaxEzKDhEaCNeA8hZfcAocECbIyX86yvv/dI+ZwkFx
d21nzuPAzUx6feNQ9iqBllL6HbvqhaEqunVzgqtTuN+JFbVQcYTom6tZo3rf4sSd
Ubly2YufneGUQIgyHu46wQutXWvBGpM23ZM5rhweioAqbsrvyBZd8zPy3tQXijVb
xDjdveIi7KCiju+rOCb5xdAUzAxeOGnLXPtdCB2H/O14nb0aZmXWo3+f61ZmVDO4
UJo8Bk+jmHw5ifIqagLyLYnl0pMAd6jObw97FsgpuPkikbhUceADz9Jdbpg2R4IL
aWM2SPlcqvkA7iiT4NX77ldccEP0Jy6zez7ULFzsMCXTnQht1iStjfOpUoR2ZdVY
5m+ILNUpTwPn8bVX9tYVcAGSYZxz9PsX9KYzyOS4ACnDoELCGJ7PNgsX5XBdvCEl
OAPACyfiRjPxEqXuIr/rPrtZmxKJWwnCQdCP8Do5sdC5/oVrjD4gIdZEPUCNkBcW
LkaD2kAbgfs+yndxDfrLETyDcgOAMiqvwVZrGiXhKwF0Den/UYldVr7nyxMP3j1M
qAPqS0WQMAHECYX1E+j00LCWxvqjkH0bZ7b5B53b8EidAp9AfSIKb9ZVSZ1BeTBN
O58sTl+a4psh+6ZKSAVEExAolxCTXu5fj5dMV0dPaJqhbyWVyfAsSJwWivTR/95P
28kNxiI1ACu3yy8I42CnqtE5TksecjS8/RpxYZc2+p6L3kjk4xfKjnA+kAei7YFy
cnDrJyI9RgXnHgGZtn1axgGA0X2oTiEqctJ1Q+KzcQQje0ePxdj2mJup4vXikCpB
ONjxOorGvlOT4VvyFQu/Ds7BqyBbdYpgihten5hWsy9BqYm4rcWl+8c+a/4jebKk
Oekh3asyg6X87+ONjts2FZS13pHkHcu3VkdncjHrdH+85khAov9Qm3nIIeUCxspe
MsZ8AcAt6gNfVMekkLIuau2gelhrG8Vsy2ZbxTvz/z1ppI9Fm/CbGgCrtqyjK8uN
o0dU5Lzk/UWoI3YJu2C4lEF1H0dEt2YVcnomq5AxFOCWs8XWLprApzl+KdMnVar/
SFHxhDOFNiH72JpEbY+HHrMupnZzuoUQygzBOTYNNoqfj0MYSWOp4P4ual2Ydcf2
HfMoYAqTKupu43mric25+IByQLKDLgp7Zf2YGTD//uAEt5pVo3LghFehrP/v4qL8
Id4Y3sVU7YZhg9TIF2LoOXziyJsz/Ppt+oU9CDL9JDGOTZLuErEpaROEpCzWGCei
69g84t4NdZloZfIdgZ4tz5/Iv33lf+6Ys493IhNnSreNN6ZlCLDmRudXm+9uStbW
BXzj70V9yeBlD8q0WYeXyGxuPvZE2dL4K21aPAIkTntV48E2joIbhXYCdFay8bI0
pf2Msqaa5tZRg/y+6J1qzPPijkMB63X3TDrz3X1mMkJTH+sUbYuYMpbVLbWeHG36
Dn45fXMjEr1B4vs9hVH9Wg0Jcx+fNZeGgWd5CuSAi2CBd1WC2g3U48/aEIbMGPOr
PsWfq9c2r2QO4X4iWBswDAIFfQMEWQonxKu7ZoWFK4bBOS6ku2HdPo3ID3IztNnY
pTuY4m017YzjTBlJ772SlpOmNYTi2fbzO/4Ric8lILLOg7wNU0y/H4qUSdIz5PyB
H0UmY1iticbCHWGSWVBol6940t9I/bQjBgy+Q6CSOUT8V9X2Jur2YvaGfr1A4KL5
NqNmuE2o3onVFqTQPyxGmm9SxucJGOCby031dTW8hEaprhJGWuwaCObnGUWBwmwV
Td78Fg07QB58aOdvTdBy+5dQ5fgwQMTzz/iJSia0MXS7/DJCT92StwR+HH16MflX
qJox72aQQo067D8WQs9ffuw/8/Wj/aBn3kBjP+HaiwQL5ibw6TYOu8wDVktqZ09J
gsdCirGLQW8vPFhagikbF4F5OUNJaKPEFNpcoQVVqBneaihHTAkPe54RMie6xzCn
PfFQn1o2BaJ5NPxJA27vCbnXLwlTCQcSf1eXYxCIEojLfKX1jPJf28R0et+5xIF/
OE0lcrqwqxq+bb8qPHK2O9TSdIEWB0wb8hF5pzGL7uOE/EUJdQ6xEX9qaRqosCa2
c9ZVWoUOTnZdJMbjApu27/BiIsaCS3XYUbmiHaLTguvQXe0gABoxdZVqQaBnpEWc
rKkr/m6b2uf9STgAGWpyTm5WUqzcyElxp/wdYIbuTRsUtD23DjEfIcoCGJYBEoGS
2HLNAGXGSv1IwvbGWzQ5eLXjdY9URi0sioc4CBlOJKxiRyLpLflIO7r1Cc6PrY4D
oMvDMFL3WsROp0NyGnZUzvKoRJtCGyBALJr5SgasFUxc0h3vrlb+5lW9sn38xL7X
J1CYzQPQzlFN+HxD3YC4cWk5GwgRwBYSK4JTh6NY6/n9hdDR4+Nd89BEzZR8FRUA
IOzAWmshhQCO/hQhGLbA4Z3EDnOgV9I2Rz3nehuaeRn2hlPARtItaiVHpFt2YApB
q8BCR9U6YpSjTDaWSdWa6x7fAOAGJ1/DHELcM6tWLtcnSZbG7r7sJn3X6SgfIUcJ
D/5d1iS3go03p/mLfb19jbJh4ZszChztsdeG8eitIQuN1wVki0g+x6WYvWetxbFW
mgTi1os/5vkqOwRJn2kdQIMHPsm31HwiTF2U8O5HB0GE2rO4cqWOzRaiFJpVwgqp
IgZBg7hkzVw+8HPw6RBNnRhn31LEcM4V92Z905hmTSGjcHdZ/fjA4ivFwYXxr5+w
SY8j97cqCLVWU+G68eVuPWBBabP686h+Jjcdu8x9wOPtjeiM40Uy1o83RpDg8+GW
aY/0go/becGrUdrz71VVN/12M1zNIbhItEVjRJX/vy+Fh/r2lxuCiBYk/k/tZWHW
oedf+DwTyMFN6oLDP5HTW6caLoHEYVGi52j5+XDwe3iLgQ/viXyvjegcJfm7MJJ9
LyIin2VN49g4TBDtY5lBNagrHJ9GqPkNab/bD5q3DOBW4aqeZYgihkAn51xy4MQg
C0zaGX5D6w0loaCCc3i611xn7tVh4UDLy4raqwf7S7I8sCIxsgJkedREEtEc7UeB
pu8jUItsMjrO8ScOaAmQskwoTHXo8nSZiEfth/aaH6xcc5OA51yCLIgdxjPoKlye
RXk+cqa5RIaoD0hEauahScqMbhohijrymeVJFPfHImlKnpptQ+bl/zeWrK4eniSs
Dje5V9aDtWS5BBrhL16sIuMp8DlnSG/62uLlFVC3WRSfxzhnJn8JMEQbxJuh4q6c
2JGlhp0PV4FNH04toNDwYigxNojtIenIzqrMRccYCs0qNsblIhoAbk2W+rOttEM9
TuXW9VlGR3/HFLchimbN3lmGt0B7PsX+zn/Uo4qRPGYS1X7RClC4yV+DnGssnIhs
tlLXgcVO1cHxs715m/ny77CCHsiJ28fUPHPLcQ2GouCpv1mDUXVUuKktq9+m67e9
pHJXn3LnT9n7SBYJrJ/+e9birCyBkoqT4i938d44FNUlUwDPOpY+We7F5EQevU7H
IR2XcwoGgMEeEL9279aYEqltOkszsB7XI1kX32dU7S7wdWkIDZXQq1ZC4DoO/PC0
ZgeDDuzzpZhmTwrBWZF8/H/s9yRm2pPEgiHREhEPMU+/1ee93qB0+8vX0mPkgjEI
62Kskf2kP5dp8UwxGwPIPMZBCJac3tfiBu2BQR2b8Bx+6aUJd3etn813Hs6MwAic
iwLpsIYU4TYoY9TMfWUbP+6yr/8Qz5GcfVSgmtuq4jzSOZvH1MmDHFbCxXXZAVNt
GN3GUrvsBJ/pb5OQAfBiHoUIidGvaIScmshcUfl9vOXSBl5fhxKXwST+FCB40jQF
xdXYqQJ+WQL9Kr5/22KX8t5tIH55AHvjg9F5jaS8/5fbzxU7AnS4yRh1Jfo6gG1l
prRAEv0pVQ8RDAjpLDpoeqRKq3gIj1JpOdnAVGzORS+M1Hun9pH7i4WBKZjS8ZYv
ku2YrDJSPAczRJ1OvkLtgQAuG3AJe3e44qtJuZDbpel14K48H5g8YfK7eDAzHZmH
/KQYy6A5fCN0sHxJR4VJCEeA81qh8Avus3H7rJBDgAxCNRHyv8y74DOGsZNXTl5q
qyKO1OEUGUNYHXPLxGLWTFA/+gbo0cd4j7kSr0KV0elvrO3sw/g63Rf1XqX/mdG8
ikYXuzmow2wNdaoRjEcBH/ATHDDTR7cgUJR2fdNwPAdnnjcUEmbxeAlPRSgNo0zK
NLiX5Ge2GENpDL52vL/k0+H3SiEXRBuaNaAFaW7wGfKY3R7GRY5+rKqePsbRIsH6
7b7mRf9bqDLgX2lJ2K/4S2MA7ZUWWpD3b6uoZIKKhQkkUuBjC/65f43o+IRfILIg
vvwu7oYQI+AGK7uldKYmdeTYju1zP2TSMv72dfJdoiYgE3Xs2ymvPddbivABQkHb
egD1O8FqS1EVSR23dcntFJRutuYysxYKylVdt6lEcFwa4ppQOkCN/RLt1+lV86U0
kTehVWr2UX116ZM7kbJoT8CHefguHD2MykRFVEvRdQJwYkwapqsb3zH23PjkMscm
gmodzww8hfp0PTEIvYPKrRyFGxbEn9i6dXzbmFoNg+xsIsm0vHgPVi2mt22bWnL0
ceBnLtENKez4/Hc3o9gbQ6wKMM0qrfmc/4s/0D4e0ZbdIayjU85XuhId3FEK6qsW
21Kyu7I8NoAPP8rPWXmJz8XRIeWakhn5uWhP7XdtM8M5BkBtCV1LAxGmjOU4lfST
WTnr33qWM6u0tLZWg34GP7uv+FUoJR4f7GOHfLkgwqWIAlE/JGx7FztI0TrvbWer
HXAb9avIaaq4UyVJ9Z+/MEVSuZfUdjHy/ZbtHWEYZTO5wuhbr1PUGIsj7FVGrC/P
GILM4J/lsBkxs24p/u5KQpbrhwhoQyY2DAw1vkeQnvYYwe9DPPIKoSgHaISUgSb6
vE3KA0g2IKR2TQ9yzfqp0DPQvA9SZCrfxwJYHbY0YbGyyiPwmWzPXQwc8ntxFgOH
gBx+C//JDnFke+QFcJeyRhD4i/6WmecV5FN8bqnzhgelRZQrAwBkD/EIZk1X40Ue
pdsbKuuSFrlgvVhqXrsHeU0/Qvf3+buMc0YhsqfuGzwLqhq6ilh8gv4A5bMufRw6
IkTCMfdpNn0P1XCJtDyTHxtN2F4o/zogINaZQcs7P0f/FzJVPi/oGlr4DXljF6wc
ErN1lf991OBFAXvu2XoASeG1chVHGg+LfUcu3Y9y6Kfvj1vC/lJT4IY3xVO61pGe
gl99B1ftootwo8v9fw4mzHoCp9uPsqWda+B0EdNq7Oiwd9if0lIu09a8AtW1hw/l
HSgRxZV09/X27o/xGBW4qD0N6BuUi1Oudsi5o2ND6CgG1b4FL2+gwNB/xnlArWVU
E9PeVyv0czbbSlJ6RIhY+dZO6TTuj81hm3l4wX/pPdHm3+CQsWz2Y1O1tNJTnaqF
qXJXi9RhZCbWgeSVJZKFC95dE7e7jJ6HVSVaYaedK6PE2DvyFj76ExzAWsE25WuC
3RAmD/HbCDf5Bp428U/zjn+t+AQj44OsQj4r2SA8mOXenVPxVkYoMymQkhFcB4ST
BxelAW1eD1vlJ46k9b//WWsqJF0W3i5h4Y8BGNk74/KAGSpiMquKbx/2EtMX2YG3
62SCyvg6Hvf8nzHGmHyz2G1dhFzUEMdn7e6V7bj30nvZAL+dkGMRSdGZUHQyDGOT
OEGjuPEcORuLfCATmLoPaiqEn9Px2E+BQQdnpEUIQlRcg0nfoqSYJ70bWBwL0N84
L4WrL9kEvosHmgCJDRusutWmVe9GC5Dwj7RYKnmLFZEjZQjGa0/aLdpxKb+62JpO
lrWaLpcJIzEoHnvi2ba/Uk28RNrXbee1l9X4Vjf0IvpCSxawmIE+uxm2kPR8wzRe
BxlqJ/Z6LorDGMhh/WT25n8QqnmDaYkIY5owT9tzr9rkC7CIy3X0o5bT+UtgnYHO
5pWHKY3IG2lyX/EbPer6/Ou97pPNRHHhujvTfg5ZQ/JjqaordvPsXbCixONgls6Z
sQdCoiWAD8dYsf1oRnmruSHJzuKPOUk1NKf1OfnxL9EZcApyWL1DYtQaR/LC+pcU
A/MvhRkiDxF/vG0fqZFxbygTsQ+AZ9urcbvPib0pwqjOtPSm/YGt+77Fs5rwVqWb
L/avmuC3IR5bz2eTSoO1y/i93ofevtI+MO+ts9VHMRU/MElA0m8ONEJQ2w40V0or
+K6qico7MvdLVvIzsP35/jD/naOrfi5mLP8pcj07QEt72SkSN1d0vRY2Hb6amRp5
iSs2f09+Tv4KTGwlLzPv6bd5becPceMNcQyaQjroN3pVuJgQwGm7+dQjIe0qQ6j+
m2SfRxp/8Z71UbBtdb/xP98S7uvsYWqdKvTP1peFqNYBXzj3RNf3FSidvZsM7GBq
cwjS7ER59zUu3F+nC7GGnPwZbJ16rWaB8U/UfjtyKO4aLR6pvxIjTxA2LPUvdBdW
ek4+7G+Ke4GoriWN7FkklpdHYZQWpNymcogZ10JqX6s9hlj1zJzB+fkrakcFVtrn
cw+to3TezjkW0g8itLdwE2AhRCH6oTkgdzRtkackeOnVQlED1o4T1Hh4LxycbBj+
KD4iSDT9dqZXS2WOK8PYYKw8Y2Qo96LvggV+SAVkXVRfuRyxWTGq16WzTai1AM3Z
Ildi1r+E0ddOqn+T9H54pR9wA4DnOUEpV7qQInHHj1Elcy+UgLlwxGNHAhV2zHIW
exy0UIJYRq4XvCgo89K2G048cTpvyrf4kcJh/IBrhNh7Pw0qEldqP4ls19++PgA9
sHDVgieE6JvG/wHUmWQR9JCAc8JRRAUJzxhqvGwF9QWty8g+QQsVd16OVRxbkFEn
w3qlY2PVx++8iNqJyepuznt91Hm0i1OAhS7H5bb7u+iyutkYl337xmw1VnJD02iP
L/RL7MCdE58Aithhvnq2Pyra1BAAyf6nVAZNiJuUw8U7OUz9OsWR0WJ+PfPvQGJX
I8UaIenef4yTOvEI/GwgRZVyups9as4zDXdM/5zsGLAvoN58jmUdDaghpmnn8N1L
UbhLqliBZmm3Ol8VcnEddmYSz5BJ1WaBm4e2gZ8g5tLgxLfHJBm4VrglcOWs6dZ1
xU14JSzbsM3+/6Ctgd4pZ9m69QL8oIEJ5R93SjzkdygsV1QOhSJpbEY98yB/R5xO
JOUEGOdcVgKhbg3V4y6bbzPgW5NkxuUhAOGRxL1nnzGUSrCKniyb1XqejrUrvA8x
qWa1l59uAvkbx5yJX1cuomGGOXQ9KwjMzM51toXbzcyVIyVpjPM+dQ1RChdctX8y
J9e3Q7c6kt4/n3NEOHTPmFvVLaZadqoGxy2rt8oWq+1MdOYIGAkHbYxy13WbuP5c
byzX0x65XCCbca4VBK+B2Q9VxHK6gMUfDFUj2jQOFGiynWQ2JjcY3swwRv42Scpx
A7uu6aVJDFfXsxZZ3i2wK/eUvYQkXhmi7mCusmNW88s/Fjup2B2HvGYhE469Yfkd
82eF7warpOKMT4N3SWkB+PjbccsL8T9wcd9jDI0SjHI91rRUAaZchealb+Jx2lsp
pLOIwBXXuWiBX4MJ97tlG5VQKxrU/wZtQJxANSvkJ8PSJoVO5hEQKYitNxFHVQ7N
hkTLgvOdHt3jnKe6Z5FFYpgY1TA0kOXQrvwcchGz+XlJm2vN+B2klX7Hay00AQRi
ueD43kEoRIMSKOo9/yNn0bhbbsMZeqbwhd6Gfnndcac6RV7vyBJMNJJW8z3AY1oW
Ely2nZP3hLhSJcYTSszzGRMK6FqtGQtoiCRPmybV9ul55FKnEuxESGfysGOfOOJC
xY5GmnxP+QPdYF80HEp2QiswUqlYCdpIgTdUoWte2LWH6A+QFZQS43xB78hYl1xv
8kQYeQl2oJ/I9bIpAhni3T9V8+SslJUqR/m0xE1EwI6vTF0Xfj4g/1C+4EZN19Nd
sLB/6Yvn8mekhOcrdTJQr7zXGc68MWGEM5iv2PxLDRLW+w7crZmdK/x5xV0jXGEs
kA3Ie+Y+fiwV20Mesg5nbfAEz/HNBda0kiq3Koc+jSJQh3Pq8CcLjNHmOf447tEY
tz9xyzvXSJxyw5LKLcnj9kClUafhpm8fMVN+VS7N5aUfNcbIDFn96hJCO/qQBaH2
WMuQlJ4ATdKvvwaSkfsDDNuFwLMF7qtcVmH1+jvIa3/iCu6pHrN06BLnD+sxyKtT
jsWyEp/pQ5AQ9M5/nTDumxZqN8RmSi0d4UTCvv0qCIHvEf/p6ir6D2+FXsHnA+tY
RputY7FAaxkK4N9Ktr0Z49TfRSOQiYKhjlAMRfnsB/PWERtSE4K63Xp/OUGxDW0z
dCHTFZ5HMFWJYDadj0JsEK2w+z6axVNY+qfy2hy/Qe1zZBicDqxbxAZh1+nXMg/N
lneXSvGCi3JeYXQQWTc0VWRrPcqzqr33p2UXoOZelZK7oo5HXVMKqdXlo/10BgyA
4jYoF8uTMBc8hbReWa6hiL8LliKts1EyPwaJLkAxAosHY2p975RE642GRGZt7brB
HaHSxjAsEagmSWZh4yvWr73AHAy5r9Ou2olBPMjz9QFjhUeqf8s1dr0M60q9qbCe
bus/cxsBFy124RpIvcrtCtS5wweS6tq7ejD4mqGtFdYqBd1F97nPSYF3O5GAwBce
X6WK+X4uE5qBlVDx3YuCMSQD3WFKhmvWcg2eShhpoSA6tI5NGVlHvUGWSkLNEtJj
DhNJ/S1dLGC+mq0b48hYF/MQt4MA5sqnrz/7fq4by3+rXLqd4j9CuS3BTuTAaX6J
ZhdGzS5ZpU4bGP9QO0NqNgFqLoRQPqGQ95cjbgwlDuXpYqnoOeeca9VHDCGsK8cH
ESRbcKUvfTXGyRk1NloAXOtPR1Hdh2pnpc/vDmN0rtsfVgW18iInKdB34SaSySt5
ELHk8GFg15zVu2OgWozcqT2GB77UrTWFIrURz5BBGmCpBtECnSxowGzKQPusF9Xz
hr6vmZlz2HZaQVMY1ut9kWpxOGWfQiZDThl/L3Rtihx8SIx3fQI7MM+/R4na45lP
Eb9jxma7LI0AbszLkLaAeIiE2Ix/auZNKRKe/ewHdVVQ5FSGfhjW4JfUBUpYSVuQ
NR2eWg1+dwu1Rp25cNci953FGj88dIYQoeXUZmcvq2Y96Cn+K/vJgsziG9enJ/2p
T23nvtmZx6Dk94t5idAsaA8op8/6ysjKBteY9QA0jB+VCLAnSsCOc1U1yxscSAEW
IDPdlGuzAaMkDyhi8SfNOArJvQnFpzIlai7R8L65+NXAz9Eo0h4EH4BZnKwVfZPi
L+2KyrqBzJWW5he95Hik58O78xdHPMtIjZUBoeRpEv5yamOBjn29+fEFgzkNn+uq
egGBTckS9TP+qx0Vb/miyD7OESPN5OTR+OF7ewhoFutILyd7chV5q50EE5CZLx3K
rvgw6uNghCLnu9lH7B26g06RHJNLjeCiZyDN19/9+ZBRicjI15nZYYAlqhxJpXRH
c6VxsF1CMHqpw3QC7qfmd7xOSQbrM9BJXTRVBxYbb7DFXUfRjdeyTPLw19lRlHIF
KN/YHi/RPosubEXxMeA0dAoyCzMVWw+YGhadgoJTl3yLhc34L4bUDGNgQb6exqF7
VoujAgDmrUTQM9txkYKwI9mhEoWyzSvRq4ibfcONbwQ1w0FpIBcZQV1XQ5rw8mQK
sgQbRumQocd118+fUMteI51S8LnIUNOnAtFmkYaMD8Dj1HQS+pyjV35uf8B0d7qR
tIEAZTUKVZBISrmYOZCDHjwNx2XvjIliu+LEGDGnN8O0H4qOi7y58HmWPfF4sCYG
p8KOJYXpYPZ1MWyNe79yg7n6kOR/H/M2BoK1mHsOWO3KRF2PKeTDF4KvlcQcp2Zu
U/AoID8a81ZjNR70Sde4v4+aCc/e+etRPDj76GBCbwdAF821F96Vb8D8efHaLzFS
bU3qNGl1KwgwEmbXjPmSzL7by1WU0wI6w2x/OUR8KvAufG85sFU5J/gk6T66U2KC
XJ1C0n/TpHsMDe5sxTav+U36GuZenm944Ed6E7yr5X99y/N/vp9vv6Oh+mlrKVe0
PgMbw8XpUlua/0BArsek/wK5bvkNV1zYYcYe71UH1kXczcCzU0d3ZQGMP8Ny2Qsk
khodlMo7C0pIpMtT0kIjUao8UIn18J9kTL7kXXZISKfbQxIZoaxtOUmPO8wgwphQ
H3dgvxPgfz/Ioki/gT6Gtg33B68z8fiZUnZ0VfcjYJGa4eslUM0rzWc7OEX/1hBj
9uOIhq/zepeUINAoWZybOFp6bhZXhpwa4JiJo3QHaRVdcfcSBoUhWilnpAT0Y+RR
C8RgFlozFkYZPybMkv2cfbZkZah6830aNvzFBiyECSHB2PNlQ0vre7Vv0z7DEM6e
RHxdoGrtgjfIeX4LcYyCrFvwo/9Mda70O51QW5zl5kC2Mldzi425FtkfSLejNFYA
zPMTzrx//wYA3AifJAdDkSe/gNB/JjtCJVs9ickfg0rNHXHjXli3kxZRmyexKYdd
3A0IZKdeETfmGjAZUk8bo7r0OI0Ulo9eJ5g4f/fEB/UhiQ17Jzus1WYv/Ac1w1xb
Tz1sTl2RhqufqN+s06p09am3QXnuNRgKGnkiBqrRW56iG0C1eitDUjfzwI1kHLD3
YLlNrfNW9zzmr1OZx/aGtSkj4XtmPAJsumxgSAaIB+ZteS8ifC88N1d7sNj+6Ywd
RMP+UsY19cq3xQp+flcjuOHlp8/zaHMWMgD23ieVnTrGITBJHOplpxvK67reo48+
MSU22l6an/JNmefGBLgN0mbnhajd8pFQ11Jz/Zkk4LxYvRNUbYEgwY/Z/ZvQTv1C
QsflSWLEwf3TJqEhIUruu1GKBHbvNholbItPw/sVLq6v5QTRWgdqMAuLVYtUknF+
OUzQUMAwJ42sPd8LlC7+ZbxZBJd64x9GM4EzealvOEeahrHMFszSlXNA5ICK0CIg
KFerZGh7Dw1oOuYoUKvuW1YFw3AQWVs7ymEL4wBRqy0ito0cznfXFERrLMFzcNTm
OECXDpUSjhqcFy7fGmCkNP/q5NTbbkZPIA8Ieph/DsDsNEZHyieUu56vvdD3YjlK
LIGRmJtvZ5e3NYEbDfsS80wNiw0rqp8SAikXwHto6r/4BSdH6b8hC1xpprnYqzj2
KbttJe0GHeJgNQtO63Q3SAuUDl7W+Px7c2MnlzxbIq7+3ZAj+zMeFl4C3fzzGI3n
mojzheoSgUYohufm4vaHvt5SKvfEkqiUdhXlR18pOxv/y/x44u/OUHmrI9T2E4g9
ObvHiMeNtils25rEnHOxyQq9ABpCjVTnR4zKqjayeicZYEMFYoajyKtXR7xnPX7f
277AhDSc/KRwe8gHGYIofUMBF9xxP2x4uCECLF7D/rfJwRlat02g+TBSgGHmA9gN
sNCKoUyM7tEujt0PQPeqxvbSHDsUfXtaTzrgzdHPNLfqt+QzSsUSPmAM6bunaa6v
u1PU2D5jfkJttquLDtK72We1xv6Pzy8HNB/Gaf8D8gN3TXiNxUnQukOg6LJIpc6h
j0x/Y+e5MuoeE7ort7t+9zHu7aZWT+SrycwWnqN/L89/I/sQgTjirfFHH9HOiGHB
JjHHQBq0lommksSOUPZK6hnBMfwsr/W0hSBRbGO/r9NFl2v7MPjvuGgFBOyC5qUo
t5WH5fgJdHHUk9Jh2b2sAcqjMiHC3y3QpAZm9tMgpGv6S0ilU++ArolXRZ4o0Ue/
nUyQ2TL5APfJw9fgDTjDGxTQFTnaqxK3Wqq3w3+57YmECYQhhGMgwOCL1Nicc2QF
tNn64vIhx4MPaVKGxStlGI2BYa8Y8hecne6JAWtvNOV6dJKO7S5UDMST9Ts++Sr2
0EgpawHBjeNuWH0qsGDhP8SotN0VBNj2qyuHBOMU5dVVYXNtezLp1qkoMRwg/ZGR
`protect end_protected