`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
bXcW0x1/qKj04BHjmHOtCwMC593wyTe6ir8/RWOCKG+3a43yDFkoOl1G9eeUyKXS
dHV6a7g5whryT9kCZ6JluvLJ3w+QXhepRDwaZoyFHKkMFQbf6TOK5yz+pf4CW/AZ
6xcHO29EWlT798v3VJYKNmkdRgnY+qUwdnwFvbaB/swsntFmLo5r0I3K8fo8f30a
6+iW0Fc7iSSuSxE0P9mq0QtX31480wfscTuk97OejV1l6f4JOIQRKPm0SJEXF9yo
P/M+8WCc96bNj7YDEbVwe3HJb33QjmvsKpZ7Nd889dWrR2BbZSUlKiQkba3jrmei
INxEzsAGb9PVHvyTHX2EAg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="92hUR4t8ZCt6mH1zQFYCjBVy5vFX0kRAX1Wae7L09Bk="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
FHvbXvwhjDf8bkqkFQRHgU1jocYsx6600GmoADeuGGKP7hQt7RcgVT72eqZipJh0
tceR/4PeBnaMZl1XTIjdDPZ9eUZH4lakjSjNEHVi8vG8Vs2pnT+X6j4VtSk9DReE
YmRyZ6pD4kjRm5CHMn8KrNw87/9hXNgQYr5AnevqFbk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="i2QALIcAkRD0JczwYIxD6+1ciaC4qMkSMP5ppFFUA4c="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16560 )
`protect data_block
FzVJn/lIRNvWz3oqAW5Keamxe8XEGyLVeUSNhj74iwdrKPnXUwNDX3+zETL+Mol6
GTP3PC/7+uwj3e5YapEJ5qr8VDHa7x+NWMY17/G+1x4p0++A73VzQCgZ6m0aQ83M
TDkIdcJUWDKCGvmrQYRemGd9HBdDWURfz87+Ro1TgtuBtymqJ1PLYbiUYpt7hkQH
vPKHf/zvyLEzMq/SHt7ENu0TV5T/SJcnLuqK7/1EPIB+HYmfuhijL0PPmm4w790T
/kxE9Ap9RGIkas1EhMEurc0AD5Bg0j2Xuvehe28lRdWA2roDbq1hQMj5ZfmIcjT9
Whmq3mlsK8zk0A0SaDr6vOuIUKVYJT7BkU/KeiffJHqyxvGrDElWeCwHBqWgUiND
MYsYBHdOxw3slod2toMyi8dIupEx1Lpwk9Wb38vBAi25YN2bYW/2jvmek0vqbn0O
qhJmqorX7FAq93Lht4/LvahwfCRXXNFI7s4rSU+vHKCF0nCpS0heM5KceLS7FBu6
xgLpevmniSp1VjmFeslRSy1VW3e3Kq0ksJtz6lfSLFS40SSSm4GJqldH7FfL24As
JB2+e0ep29SthURema/DP+o+RmAq/WfAiaszJYOkXuhf+hYVN/fUQxszFZ1rxyz4
0YV9h0qn6oi4l+xD16cHsICrgMRClLFmd/I/vHDybzj9bjC0wetGnLNSlQpdlvgk
SoVKw/MriqNg625PHIbfrrnNyKOnqnoP2yZ0qN/tk+7oai+1gAZed7LXRwCj83QA
FB0YqOMHgPgmqtxWlqJuS3aVEJylBe2LJPhSNOLl3edN5K2Ytml+GtlLp41ZJYRU
Y8SYkfMlj2z2e9GqEzmEsxkkwIVgcadURjpt5STkIRZ+pV1dK84HN3fV2cdRxKcz
UNCU6cUjyfKC1tTGZtQW3iTlg7v0JJ+1rnS0ZKfw8qNBzNXi1hZU3XfPbSjBdh36
t06JWZMd3MwEqPOTXOYARCErlQnShFaQ9erAEktSGOsh1uyv50eBqj26yOOa2dGD
5jMLiGDmg9bFk/Yvr+FMN5tHEOmNh035gIbDvQKWogvLiZza8IdiZF0elZreqQU7
PyhkBaZ2AZ0LGV/idW/s58GjAbCUuDIZsx8DFHs086mJlMQYfK3T0dPB5riGj/v4
8WX+gLzpZaCLLR9oeZbd9sXhBfliaZf6msLahjq7pjxNpCbaKH8UDBOe3EpwOGyU
eOcUbAvQLmQ/elR17FcyDUhOGRQURjwgoiqQb1an7X+ajjfXv98tvOrrNVYt5YHO
qpCXVI3ww3pWOFtefa3crg1eP0rq3NWsNyKr9yipQ4fzmJ6kZBCx44YXdli/PJBd
UB1ErBJhCKomOmUueF4SE2yx4GzETzBHolavbHwMHue0avWbvmI2W9QmfBiTqrnF
WqPG2kSYMceLGVqbmuC+hUVdec49XjXCh719xcxXsI0RdpCMA9nFNJwsqjx+Jzv0
9UUhqQzyRTC9V6AzJSD+6r3dWtd8JZOIybMKZaRH5rxpDnlMI/7evMdAiLOXQixj
nSAuja6WUIcU+buPLfDHHe6VFqHcgf+MvwtMOOixPbyDybEj23rFvHU/ZOK6rchh
nkV1m5/It5nR3ptECp/Ufid+iRQBU+xlpvSZ7Uu+LfJVe5o/dj54eVEAaT+/+sLC
54x3CR06BDPCIZw+zn1gqbbH8GwvX1SFGCg80UHrR4He/Ddm1OJADyockkcnlm05
uHuKNRUQCSPbhW5DciHS6oOEhKRdNo8sZkErCV4YQjn2zZXDHfqb2O2lrt+j/ObY
k0pI64YW3yuhLDj3bSBYhJV++S9KRJGVomh/+gRBBhOwKtLobxwmc7nw0qWi8IQg
GDwsLvtpsee2RcSUMgHgqrFbgBJiGLxPasaA9KLxjLWTpYDmh/mm+eELxLyNZrSN
tm9nX56yZ8rl/AlxlyxkFqNAyxIrqPzGbGbkGvFVXRu9DmTIY/3BYP5RGoyswiCE
0xvNYERCz8r+E9BuzMCRwVYVDk6N1kbXy2g0pbaFNSPi/b7lFfLvqFjArH4BuAaj
T7KCEmF1ibQI0Twdl43ay5ANjK10bfEarecw/NhVColQQpbn9DIm4MfxBLEkT+As
PScloZoxTHHvfOGeg8sTmFnxHIyzx72FJKVey/+4IefOUNjNghqoVqp+QRya2OMJ
xc+sOTFREVKCbFpLgHnjgB2qXdha3sw3b8oGsrVAGjWwx9ffq2lETOkZAVy/iGE8
5C9TvbXJhWX0VhG7w3sH3ixh11mJRSehESdGjij78w5BSvI2IRufy+gMOKqXZHNy
EP9J24rO/lHPP7Ek1rGr+Mg/4M6zyV4FVjtIoxs0aEisv37LwgvliYli94vQhSVW
kE7SHHe8OR6v68NV6ZGsi6bLJfSShcq8bNZ48xZD39Kq+q57QodMia6cwdUqpQey
rtkSyc4g/V8PZrDb8fbmZaTN+MUvul2W9PL59FYmVy9HPwpvawJWAeKO4J9CsIn+
4CFPYU/CVIUvuaNDxSl0C1+MCcB3D08e7GTMd0diN6+7DX0zXJQrQ4dh4RlwIWfH
bnQxWYGGy8ELtdD/V6dYwCwiSWGU6y4crZNUNucdxqPkGsxJPEDp9RMvdc/Sy84V
HGHQw8TNY6dlfEWTjM8rLHDyAgOXNlWmgkI+ZQva0rOey4hU40ybz6d38z14UsBA
qzEKYbWie9R3Wfnxhg9PTNbwCpYGgNc5tMFFajQGrR6A9izN17go6nkoQgpl6VhT
YMm/rlUJUVLcUsl9eI7dLJcxeAMmzqPlZdkrNKEaRyZV5uHv3t/mKDwuWoK9mW6P
cECXphy7TuDGQrV4D3pz73jrkOlj8FCq2hZ/EZR0Q0lcfDi3Jb+J1KhwDIx6vM8p
ep5Sz3F5Ckp+TcAh0bK4CciBxUePXfPKCaPY+gT35FHUqDcVHomN3yy41o4NxeK7
VR8uQnbvk6zUZRwXhq8v814Hxp7EjbW325wCwY0o3qyDVwJVuX8K5sowkWXnjOyP
3JHNIhcDiGs7yju9RYb4bdZ9TWgS5Bpob0S7B/UKAYnwrt4iAiZBNXkFobMkH+13
1FupO3wiYtGymMnsMKyv0mYxIivTdb6Q9JgM//h6+3sdkvBPltgnoCxcqaDdG1Rc
yZaBWnqggKJkTNPf8Nx5vX1OgNF5JmKMnxgoez4kFMSdbU/XukHedVeKTa/msHYC
REIQ1fb3lZPyTuGPcE5fDfDE3oTy35LMEvLb1t1g3skfMCApKhlWA935DFYAvo99
13/JMDn0tkbZnaJQU+G0zXHeVDSmdmRXTHzuceMhpGqBNuy/+x3P6kw23W26eC7C
feQORgnXrqfDuVSfrEPDFwE/Fny3uHtWBDmwqXgftZ9rixYK1WCSOIxbGndoRUZ9
hSlxUBO85cGQx/UmgcrzBM45ri2L3T6HudQud6SlOb7kVWpE7kczu31yMjitwSgQ
FRFzYtHkPbyEo4w0Y1LZNsQb6wIgPBgAl1M233xQquws0nn5Z8at547TFfyF0P+4
bMqsFfbSSSjB/m5f1pg268dIFfZln5IlQVKH+qnytOsIemeqL6JWn2gZGlhhGDGT
dK7avgMpdfiPOQ27N69kzW9I7dPY9TJqko8VdiKm2mBURlK49Ktv+nGRqMYV5MEJ
oo5MknaZuVDPdLu6uGO6iDFaEUwzf8vY3Tc89JyjURltW2+bjn2DLDlIj+b5QXP4
+PCVu4ClF0lwc0BhjzGAZI35KPlapRTsiG8ZYcSpgpW2ZI9Yj20+ugIK6mJy53wx
Q2MdppYNZa7DkE0IW2KhNA49ULjO7QJ/pWn9g/Nl/cpUKeCFiUAjY3sg7I4TDr7G
EF866KoN2ugURMMKKZjadYXNs5YgDwpwnaFF40d6dFYSeewQu+XpD01Tg/PXpfF7
UWTLgBduJdt2WZg65W0opVYD3d/Aqxy0iXb/yGoWCMFlWIf+fRYo5GPQHHmRphwo
4O5K0LnYyIJJ04TfDPczu4s85AXaXj1qNslaAzwAcogOq8gGJfqQtwkDNBEDZbtD
vlOiZLY0c+Lx9MbAE7xQPf5QtFNz5TMF9oxHk9LOfihegf77MTaqYO/Uq9eb/pcW
evOnPlQwF9IZdf1EgLOgO54HviQphc/Nq7rtRceveeehC4WUAHxNJKgt1z7FTES4
wm0i2U1vyK13ljlKcZ33H7tOrDxv3Up2EsVmNHadenRsi2zvnF+1uty7YsiI4Kwe
26wP0F87saxlZb7gfr5nThds/mvbkGONoVI0gKnEwlSDCcWrURu+R9BlSyJEyE2k
74w+LsLZr9Pa4IQEcCUIlAXFLlYqI8s6yMHtMqp7K8dq2ADbLRvdUWporQhNLtF/
AFzJsO2H44tLl8KGAYTOV1l6iQO6of5zzoGuFya82AqtiAYdsFuLnYpyTbtwiWEW
74bZX21hcu55tnnFVpzmvuYuuMH7cYLsbeWXS5CQvjFAAZWr1sdHwAwBRrX3ZHYL
G/+NgPHXIGHyLWb+bczkOBtVsQ2u6njEFiq/NnMcGe5g8EUm4oQyxAJDxSfY7mkc
8kGPcyp3kkymqjGHmrIFrsDSleib8Cgr+MwfKj46Sxwv9vKE4Sz7C2LKblhgsZOi
/a7JjML9y+a+EE/Aph7w/ZkSloBtL2SLUYl6VssDUBmy8FJA2W2cMmCegy9rUrb2
0vqrWhaIZ3bpaJUIEBiYNVCItX6WxrX2FpffoKSdMZWWbt9QcyHHB0fbWyKdUDFh
5K0hZeZzfMniDIjNZj+HVW1H9nxDL4etPlfBojUR+1EAVXt7NjxaN6y7Qy4NJurG
7i+7yB6eUmk5nr4jBK9uQKjxft01cynDInGEj/dU76qUhxPDPnCnKm/dkPUqlumg
SbVUSNq4xS44JQ9R7BIZA6QEoNp9P8+nQq/gzX3kulqCdfZ6h828vK6/4aNkF/8R
10iGvdhtN5OsI1HR1lfce1v1rrsGTwSn5c+vZU5XnoqBKk3fOXGcs5zpRVHNe1EE
+HacESHboaDv2tm+o2GqkmQ6movl+LQ+02oBO54tg1s6OZeneWOstvz799tQmUmH
OALmtbxE+gxHS5txuWLMvv2RmTv3b2y8/erdmIuq8zboWz8ap3Xz1wBGOroyBF7a
dTNNowZmeL3EhV7/N20z3KyGtmztQeqUv162u/NQnf5MEd7f5OanVqYDbm61WruI
4yTOrMzqkuhFKgZIO6fNvDoQe8nJJ2HV7Lkx9hCQ8Q4ZTJRSbOuhNs+n/er9tjch
dg6JVlM4+bK8PkjqMoOVYyopMnqD/vH2ktnJ14SEWP1/Rd88bX+1w8Cq2ajw5KX2
xOIWQouNwu7b0ZrEwFS0YVTgzMUcvfHp6JtrVm8fGLiEMoSSPO4m4rz/s7i5X2qO
VNUigK2n+d4z13Ufie6LxPLqQ4WoAy4z9xwJcrqKqIqom/KrV/o2AxhXkhKEk2uT
2pu2F5XtsGW44/odF8smFX2Oc8KV+6AYGlNliURX1/sKwsTUfalpTmaQppp6h2/5
17cdOVywbFnIA3a3yxyVuUiwc6kT3xwbT2+UJ1ofrMZvWutMP2wyNH3N5YyS2mlT
hKkQv8+pByYJs5DzRW1qS+zvAKKbYZ6hzMDS5t8ugrm2lceOSBQt499wHJzBqcyB
7D4o4FGDnJg7vV7RhUO14wxHhsrzI8te4dwmjPLqWQvJ32k54aKyiWNbaBOitUNL
To27MzfDUKho/dOMzvkSoAVWOIyEBdd8JtfeSageegQUBzzBAA+g4FhZ5StIoNrB
xEl0lRC0sdtqxOloNe3GBoXZoXaOnerIqTv7jcMXrz4Eqh2UlUMDTqFJa/mCQomk
kUAxuezuJx1CsrDOHBEDGngvnEiNafiQ+Pf3D5Xb56YzmIu3p7+W8fGqGrcBs/vH
nhlxzN79JpVUjSEP/FTblqXyEy3OtkcvvoYDMvK+Fo3uXVLJe6+KcTx/yFzO1c1S
687nPItz0YrmF8jInixNBp0BuYarQU3YQIegKUWXsmNaRIIEFlPTSJIxjgH9BLkW
rVUKHg6kpmFed/L7STtiTownxNWTwMchhMujmhrfAhXcRAU714jgbtWgXTMeN43S
DYtFMJcACczEaISZ363NoZiERRMvUhweymNgm+fn6YBCsCXgs4hjQkCoOGeP7dwA
RzPO5XaP3V9QBzDvtqafpapW+35aJeBqIXTBndQOmi9tuKxTZXpoGx15IHrh0t+k
ok0LrlxknDdjlNrzepLhEA+49mao4zCYbGNVJ41NTskwWUTYbJrro35mcPmEY0nN
W151quAzgFaHfHTEOgxEPnEJERUw5QB2B10cLmBkvG31yNVegOJhAzGbbJDQWFm4
lWs/WKXb/PB5WEQ6JCl/QmfF5bc6miL5Y3wtdAAGrKdn0vqchyejk/lh8TSFpW1+
14APxldaMtxGT1xr8U/ndiqGCpFtIFq4Mg2vu8L+g/M9+RHhV5epiRo9/G5NC7Zv
1Y6pFDlqPxVdaLeWipctLDxfAtPnwQBSLlrhUOfpQQQ/CHpsn0dCteNTTlMtHQke
3dJkvIvIXOb186z6bepnIUd3gWeX2UTFl8mR/YoUbah5c60kL4sDVKYuEiy6LwCL
uGYpFRJX297PwrYMshPf3EIi5l8FfJgq61wstoBomXlxg0pIFaFr1xyGwZNbICk9
2yVUb780jEKy2gtgqDy6naNekwfEpEcLabr6XLAUsa3V7wrrgYmh484UcHRtO+di
NyxqVuLfQONYGGAC2l3ovDrRzNp65Lk/DmThFDlOIXHU0X7b1pdhhROoRY31RBGJ
xTIPjDc8BTH3yTAwyslH8hYk9Em5ubyj5Vnz0HXZV2Hp9Zx/y7rKjiU7kp5mbFAO
Ib8oAcGO/3eBKjBvORxTAzF6YnUznq6iDfdd39bsry9MI57qeqxqn9x+Elt3G4Ng
sYIqE1fPAOT9lTQx5Q1wbl3yklEMKXBcIyhyN0AH07NX433G8EMrSF0bONytguQH
hk0qBezJbjgxVxbme0rpLJq+IBIqASeaWuzoHp3JB5QvaGj9kAceYv3Ff38sQ/pb
DJzkK2liT6nUuI2FJk1nSkA0raqDeBprK7TuPtYiFbk49squ0aCr/St7TRsZpE8z
0vqavnY5kDPvigO6i3F4LfP+xxeo6aek+f2TYgOqLhcYgsW2BFpsVvuFvB7lXhtQ
Z1DRtxF9qR4sS4Yc9vQnjPO2U4h/0tyP0bq3VuzoevG9ONoZ5kxfEgi7OH3jaiot
poly75oj42esBjj1iXyhiqeAvBPOXlwBuXXHvTa4HLM3Ihhw/8sncApnOt/DjsAV
h+tec4uw3lgG5kI1CA9jjfg1RYeZeKUzCb/D8Rl011+pha8bKvk1ZEoEdvWH2wRY
PXBStKoO6eypabuFhkJOJl57W/BGG47RpnXNtcU4VDlivB8v67kAOlES6jGln0s5
KyWcgmhrSUavYbKboMIB95yTKtlHRGFkZa9Z2booDUSEl6H+xhY9is+6yTGrMrkC
yb+UpbeZNhODZZhDVrvUmN1fhAkS/umUeGJz3gBxwifwm8fKssyho2jLau6zB38m
V2OoG3nALkTqBYArXdKz6SH6E8/6XBeBLTy+NI2OUOosKXwBFZgwzq1LW9ByNcHJ
nwZJ1l4n8Ha6lrnPq034cngsHFfT0jH62VbAStjc8IzOBLYfSHhSuUAHe/x42jST
mBcxsYs/Tknfo0IKYlyIuquV9TeGuZXxf3LA6u8dOwkrM9KU0g4HUUo3Lc5kERfV
dVoQyF2fwyA0J8iR9ppv4MNNBV5lmyUrLDeYYCeUqucFifi3Hea5qS/bJAYYwCS9
9rmCCo7r88WRqabaUHbsfx5t0c08KmIkw9qIcHqGUmQ2URHQu+WGl4hlSWwikhid
sIA6cCh36YX9El+KeJd4hh+7Dg4SdmDUcGCXfS7xJ+PI+gW52OkINPHuCrtDZv1w
pjcHR7bdBtFlyEqDQo0WQ1fYevA1Pw50rB9jzIROw4IEwnfHx3ANmw/BchvO/vwb
C3aW/u6m9JGup3U6PT+dnMCc4d4cYBylsmewQL/2f+1EC3TgIwMSqFsY6H11TovD
cONJHS2JScs/jCFSexd1Od34J+Sa7XSAsiy1d2Xc00cvXUzeSNbBSXpnPWTx/TeG
J9D6liCTA5+72WlPOfuYNc2keBhrMQHAHVhaZ/Xjcup3NIfWH4wkiLS/cqtNT/FN
z1UEm1LfhQ4dBQM8OHq4xUJyJz8NL5J3MdiSC79nvrY4uxAsBZLENAjACR7/byFB
7QyAFk4WeQ9s2AQTacpcF55GG9UoKzmyKHLAlsHfflgpAgUoP9BodiQK4HCGd9TB
GVX6FBrQpCkHyToTRP+WLN25bb8dKkJFaTnX+fKMJgIoj4+KkRQK+Zwv4qHTyBLE
i6aoC65U13fYCEh8ClV0ZtGdceYNKGIv383zQta6pEpoqR60Nl0Gzp16qfnwiPRT
yr72KJlPzPZWK81EkHfy9GW1KmDQEVLACaLSX8NBLD1SNyENAsA5vjMIMbW67UrQ
K3Nux7v8dVZdeHwRuJNexE/utOfzWlxwLyQQWlHJaenbwFuut2AqGiBjGCXUVMuR
QObdvarKOCodPsONQRF7ot+ryYh0blOfjUxCOhkhkyuAg7uE/83B34eZz4s0R6ma
5EkDrQdvkkdMFk/AkKg9Ef9pG71WwMfqFZHZUHNM5BCqvK3OUTFthmv1y756hz5B
UgVovgVlJ+9Xe1uU6wPn7aNV6oNS1sqMAs0b3N6zNWnhZqjkRUjuPXQxOdj/xIqy
3TlbZ95iE9HMGD+9VanFaomS1B+hFXIozKA1KQiqrWiYWs0YjBYAEdynt0kk39/f
TdATLLjrUy8wYitj1Ylh8IoPQAJ3ctYL/mo8FeCeZk7lRLFqxxcnYiEy8n0RUNsE
gsQiFqvj1uPVTwjVj//BHS77jQ9IYPOZ6gSelY/NSmkS9ekdOLEuXrZIKsIqvKGv
mYSGbKpH6xMUEZzy09Xgv7nGQNGlrU8VpZfBo9D4LLv5NfnGiz/xV+cdEY97dh3v
mmjjdbBQdBiXWnLSv31uEySEenY87+Ype3/GDo2ricWSXDostQi/URRtWM2CcAK9
KAdwmbVAfFkfGDVmyFbYlUqwWGWVM1z9/ra/SPitVnSNNcgGu4DddkakXsj7SwjC
/DmxZ7Ah+af+917mVEUtNxi+IEFdF5nDsM1JJB2T+US6D1n/rIbF8eGb2KuAKYq6
Ws9k4D+stHs/xUZTlRjCQFDzAiBc9pZ8hWxQ1674VmyWt9zBQhiJdp0L2CFN3DY3
UWtJdM3lyq8kOjPobvCeokuUcpuvLnItZzZKQiNjrZF6bm5L1shcL4FrEg+mNSRk
Y6+QoEFePFCOmBHNLVj3Hv46Vjy2b3CegNWt2IfvI16RKUQhFfH1xtoEt8rEpO3X
kGlJ1Hhble0ufu86b5x62pTibxYpeHeVxIt3BGqssHtFdkSmqCEb+n78/RSIScqv
eqCXOmKTBuNqGoPaAvXTSwSGoWaHgjisSYbb1Qja/DAkP8IaorkoMENhz8uJyI0O
7W0L0DYJhJGBkDvoSOq/lfKv/ticcMVx7iBGXWFGMnKbqcjBqnr7m6YDPFFffe4z
FmRPxtyUKXNj9z8IpQ2rtKvxKjAq/d9MCWk8y0MPIUIIuhfZ54dhDicbPbkvEjOq
p7/PLeXAsJ058Pb5U0Q1gwjCkI1E+SGz6k/yeUs5Z2l3lKbIMYKryW07H/4h7X4n
M/TI/3qGwCeqp9eVWXeYMjw6tXf02g23LV2cbiBRxVG5sPM89JSNDFAzt9eIkefL
Z8qei0egg+3RnlGih8E2CJc3P//pFoImnePo6qw5RQ7ylPdFi4xySMuzfq77uZ48
VfZpa4OFljfN1xEgqbGHyB6ilFhxDtiAmxxLIqSZtVQEGjf9HlUCGWMPt9ogEjRg
NoMAcncQA7QY/mtJScNiU/KV1ZeNGlIZzUTDJw81BVKl4ZfGBntUuxcHjHiRtswC
8jjb2F5gu4KDA0lTKR/21wuGZY9L2Q+1yuch3qHkvGeB5NdHv01hG2zuvQoXv6pW
2uukS7S2oL0ITbRbzpUJSbqEnNAWeJsZRlivJDF1jppHaO0TUp3G1VcVtgk2Ddzw
XoLluRHtcnWJ1CsYRtpCLbhjGtENwEoUoKWVhNEtWEcjdD/eMLCxR/yYX2C62q9W
6Uefiv0xBEPTFGgthPBIjf+AMNC8QjS7tbwZVKPJW9NDPA7xr3v1lu/QUryfoRr6
OCST2JPge4wU7cFOodHSzcj6WSVecgt1SA/6ZmhQh5hjy8Qp0G3JapXZgn+vvVNl
3wHi9vcKnvGLE9EahO/rSlcamha2dSvSCh/GvXGvoP6t6fQYnmbOeT6UwM8M7+5A
zU856JwwUbBVy6p37sdiPws+nnCsWwsetw+ZaHeZ0ArqzkXPzA2lYad3/Xnbd1Ik
KY7nyzQFkBvfskIMRc+oSNSLGghzwv9IjLmMMXpvVik7tFD39eeG6FRgS+ICFr/B
+8xnuJbzdXTYETa57VyDOSTMSTukHifyB/fgKYnAsGxyw2jpAEwV49VmIRgTLItZ
cUYew2JZfjdqetHjNY0d9eIMT+LthXHfEivqo+nK6yMB7ljC7COzgleze1Ju6hYx
E6L3/ErnodxT2ncis+soy3OCV3b4RTz+8xvQFgT2ZxFTAgrF/pmxMcGDkgpO1uSA
VrukkjGwJ0Y9J8CEs0oowRvEEmuk/CpK8vpfIpcTf54beK32pUWSr4ua+oS1Yd4c
0OCpBnNp6sI8+2tNmQwEV0KUyr90hkufKRvoTzOJy87Aya996MCUw16j/8KQDRmZ
TGC0iMDYgj2raEhBmykpqF5N7ZjAW5NXeF7QuxS2ydtOVS3mr3JcGMpQGO/BvIKY
q2kSAY/QuhO31NZrXhj6atJELb6zcAUOuWL5GserxS2g++aWmYSlt2JcBCFyD4ir
II7kwXjPfiSO0QPvToqj358SfdzWrUq221gjTh4LElpvniJIBlAyjH8wWvBFbxcy
zRQpDV8Mau48pZ7OkSH5zQfhT0JC+hkrbcMwbhIV6q3vrsmBXumYtRWgV7gGRC1a
PBOfCUuT8EXnCx5gCWPyx3hdm0QTgwu0+9NukZf0Tlu9h916OCjRdENnwit/VeAc
cJ+XV9Bn4RWxT6n1iMEFjMBj483LDkMJGLak3OH//rt/0Ny6VJsChudajiUXz1gd
dJypQdmbIt9LxC2xTLKeCXAnLD+VzfemK1wkkH+HHkR3nHOOZwMqmY+hpnJweC7o
tJPAh06GAWuKcqvPlv97m7kiR7oMxQtr+Yo0zuacx7b8/h3OuEYMWXkZraQ8gmsM
XkpkDNrpdKJZYR0i5x8yaLE65QbBYJEYoc/3t7x60qGPdwWe4uVzFOczvNUZiWjE
pzWkyyDTkHlwBPccezXNV6PCPU59iw+s5lolX3AEz5ax3bkC9obHskCIQclWl+Qf
PCpkqZ5/NQxotinGW752OWQ+zh87bogpueDbaVJk5cfM7rwo2/RL9BVbPP0brRyl
t1S8laIF/Tp5zCxbMBfLHaRgJOiQ7YwVJZbVbuC+Lbg3am3alRtRTb74AH2FQyum
QgNWCVdUv902MZwFLMTLqgj+lvAh6zhNj6RwI5Rbun2EHdUt7i/tXlwbpxjTfnTx
QUkJPCQbjpUVCH2jScN4eDF4TvC/kdUC/YX2eYhYBwr7tSBqmyvTkfkuwgRiR05h
59BlYGfCX46mKnjrnqfKgt5fIqu4tay/CpZKHhK2qowkgOg0GKgxKjxMCI715xKV
rP2AcluhgOjXJ9gYt09/Q7Zb8J+K7JdmIG2f7ZEox4eGHsMA8bIEiTeOdXwBRg+s
CTfxCGtmQPk72E5xXducUrphvwR5FOb+NsTAM8y7VBxkQ+k8ezyr0rRWsisDCTMP
HRPQ/J9reIbtprcOZxjhL7mJsL7KJxwYprKtidQPTwIQ2W094t6lJbQWJrUktTtR
+bZsO/ncyWaciHoxaArxw7UsNsJGTBZfAXiR4RF9a35oGE9/Y5gJDzNoTiUY2fC0
VwdTwg4ddUbpOLT0CAlmc8glCfrw3PI9rY4N4OD+moCUYIlzyUqd0arqPWgckQEb
/lYKlR9fzsiSQT0PV2kWhpES/4F1IgPg48Djlpvg5GsTfSvoWsAbgo/rFDiYdd9M
B24agKibt3yC072MMZmeFjtsnXehy79sm++gt6jsHJkxO7B98+rjBFPflSqLC+PO
ncj5SPgwrt/iddfrACDIp9jf0U16rl9iwEYDB+48Z9IJ0QHOal66+5tWYXBvtj/a
qiLVAgvEoO5cd+oc6Gg+I37MCf9deIQcVxJSaqZy5i4XRWyjfQI04mbpJiOZid2A
vinIaYfDOM1gb3C3zYMdD824Rs3pASxD40u+Q3pSHPVuF7d+rXun61hjoD3R8hmI
gIYGhlAzlNE30dIktmeMqBFRYt4K0GnkU8iumngmiX8p0p5dGQdjyRN9fEymo6Ih
t/Zm4dkvio1n6YEk38OljyHNbAuVtEMwYssWnliNbeGgA3O6h52LP2IUcn2ngiq9
N2nqEjEoquLdltteuEHOU9bhEhJrA6ykyXC3MiceN5sJx9X7I+Ls7Y3GJW0IhjWu
x2AB3ps6rggZxBUCfEJu3y8e+vIPHMV0VqpqsOeM6uE9FiYZSJ3xVdMUdyDdudqz
kUK61KLraGoxFY8ReXf2JBeyDWnfH/bjOY88AAEMjSse4RgOyuDXb6c24GvAgkiw
wMKfqekYSaa42acntjL+wbLcnrTCAvJSKZ6wTkSptAr9cXalVukHmZaL7Vayq8Dy
hqUzhbYxUnhaKDrVyiR3uH7RQhPkdqqLzuwlWjkzWWAdjYMs/DnaDoNMJ4um092P
CrwSetmKW6GNoIIhd8nGXqum6qFJX9GQpQesK15EALi3uztHgyMBlmKbuB3j3psT
AdzpKAzkxXnHa0/w77esvpFESZByCRoTWvPlVG0Aanp9QtmHRWd8sHER3XWXSewJ
aT2CQg2TeNjV6CTJBJJmYa/iTYTNzbBUjjnWKuqlxDP+e9b3WXDB509i5sc2zUT5
Ax2hJdqJzp2bEKG9WtZlkMpz8GFRY8HZiEGTLe2jBSwWcZcB2K/5gmsoVyJu1+ir
zqo/Q2DFYZxYxc4lsPLebfBrL31DEtXDZN2NT1szLARWQvavAokWeoWcoSXTb05Q
5lEh3sjKiMYcN6FvGqLev4sbCERunsGuNDoE77zdy+mOBduUUOF+dlzY8nau54cR
TXbA43sDPXRdbTQS7gynvAKfALUHCXn93EQq4y8Tn6rOEAyZFS9ZHFhDVyDzJ0Gi
fbfL1Rg/ZNd2n7uY7QDvpLx92zMoRywgbegKN47mz2SzOu+eQPiT0PppBdZkp8w/
CJyBlJOFeJzf7aCnKdf8nHNxrNo9iACHYBenZix/HDN4Lnq7Yvzctyd2Rztzb+6u
K4yOC5nx2oFzvdK8JvRtx6FfnTFv6X31OTEAkB/6KNA9+DWOe0KuyWCCeywf6oIV
PsJowpCtP5xlQcG0ZH7tvkDXT2oN+r6kti8nTqrJuZ96HpGvobCtloBtcX3xlVG/
DXq0lQA0Blem8sZ94woEHAlEOJgdAOhS3bt0tnIrKbTXVXLKc0l/L3gXxIyeaIRw
ia7g3AraQjdCb1i8j5xy8tUGHEWWTjssCV4k0PM/3S9aAgXSpXEi/oV34qIIqMBC
Tgk4jR0JxKOfEDpu5P1xDAIrN5vJp/9p0pArXO/yvH2zZMzxqpHYM6fA4bxPzDYU
Z8mlhWAB0CLJBZKrOIpRqt0NWZ6nT1BrENQS7tJGEu4qmFwyZ8/wK915yBlTWhL5
xl/LRy2ryJ3MmRkrDuVqW3RmnfkrqDVFp2+uFuH2lRHABu6y/K8Y10SE8BZSDPuz
IXWkzbSjNgIL4NanxBhGTX2KLpGx8WGtwj8uzDjcVwqOgLmHfbzLGTFKNrOhn8pa
fpvi8i97M0kTGhmgXOHK2MNsCCNTgLJ24N7TP46w4jzCLGycf07mC2+BdRQ/UUYV
pJGgS5uzhWUnvcdb79YiugI+48u6UOt8v1W69yDFjepgMeGLypNS9jfmJ+Dza9ma
XY6uYMBgYLfuIG8z7pJ/LrCJu0R8V9+kBJ+FCigCN/dDkTtHkQWMCZt1R7uE+G7T
FyQ3ahKQ9959aeHK89kvbxQLU35v1dZptCeArZTI4umPni/JK4kP5sYplzHx4Ic1
NqvLYbenIkdY+Y10doBjZ3RFcwHsNmVP4ajGZyd2e1WzLX3sCtyI/sW9orAfaONh
kIXaIzxmrIu1RCXflUypEgevfbvuzDhE54l0vE8TIEgbv8OObtRYdthwfX36Z4wM
QBgw9rx5ZajiRbdvjVgA0QG6Ter0FqxF0nao5wVTK46ziRT5SXH3ZZ2HU5up080s
fVBsFg4xP3QZqefrkKm+SvAnsRFE6SsMKAvJkQPS2ALTy37u/XS4qG9giN7X4d+7
SjJrXJX/bF8st/Aq8od/bL30qjil0USPPOeMpMvfGD+ZLJV/JYh48S9Xz/oaK7/y
GNvJB8IISHm/rikQYCKET0rBsxhiPwunLR7Rwi3Z5lH7uRti53psDWmjSYe/bh7o
U8sPSgqA0SpH7XcdSApvih0b04flpNPvUIGkEO3lrOnFCOAUh0gkFIkGDqRmFav9
7t21qS96Mor2m2xMPnogmuRXEyr06OVv9xng1ME1qvhi2c0lOp/2k1q8OK5Vo9Mo
JmfUu31ombQNmfqT4BbfQBoEY5/U8FWDbzCQ9B7G8yK9gbzascD7Ebtu0pBLhHVx
Iq8gFZBEE3AmRnlnLVlI8iJD3EdWgKXISSVAcJ9akHvgzRyTQSfueDZCBNJFko6Y
xnrSMv+pmzq0D1WFXpJx1fjK1ERjX8+C34sX+nCXrXjid4Ozyle24rSFYBNcupdM
oJLc23Vj5dU/eUSbx2Pl4WPQex06SVLN1CQRk6aGzpCY4pifCXlxb/xvAPO4ChGp
U08r88tkCuLnljpL08s3ZjYRQY+K1GKAK7IQZxzodK0+ENGJOB0CL3639wTok6Tl
u0NCDU+VtJRU6Jn9m+MTA9GGnLXQ7y+mw/pg6HW0vF00KLnNIyU9fDWjWjeOqO+d
fVJW1iLEjXT6ebk73hJRoUEB7Qj2HsSPXTAyz12tz6SrDprD0KUpK7terNYUdEbP
Z9Ik2myy1A9X4C750YnDkLBYVr2YRhcL9uIXn3BxJIWyjeS56lccrq0e1huh6mZo
E/rqbpUNb4Uo5mtzaZ6wgXujI8g6IpkyIcDHkB7XAaDMfxV0Izd1ZfAAQ6KCcFUF
lNjr6JV3RNR8v/7bRw4MjO8Vf/4egXuA4tZQtZCHLByNSeEYglF4rPTlqrsmAivJ
Lv+zn3g9g77mdMzcN7/slGSmEuxtKE/eBgR+K3nuuvrXoSuQpkQMl00iCW0aZsO7
DEER+V3swG0tlYw20YCYvpFdDOJbF/yljKjD5K/Y1yiZ3iQ20dW8Wa+Pl7qpYE3e
N0zNmw66zln6wSRF9ufGDciRIpgrZeYxpZw/xBZ1UfmZiwdGcvTDkc5tEqCJ2+kL
tTM3e/ficZqgsWwGqNRRv2rQ9F6pBCU0H7aMEmRnfSpni+bMy4SHImfvnCIQlZta
FVYsSMr3/lXjYhYPmxSSTH06qzJREmpAGsufESY/uQcf7uAMHMKR13u53Oed9PnG
Lk6BTY5FCTY8CBE7Wu45lbP6MPWjxlFgbJI16V3fDmfSs542kfnDTM9GhednEud5
nnmdK6hkG+FN1km+JJXy8P3lFUqYRYXPWzcyQl+CtKhFbKO8jliDuE5jHEuRuUmO
HeOvZRss0BxOfLv7APEwucBzYUbNZF9BASKpiFClRCfHgbmCtbZDBbdB0p5xvdmF
r8ocoJ5CvezzwLbLeWrcsEiOGao14aBo3UbR6dpPBBAF9Gxipub2rIOygelXJx8N
HDe6opPXb31wnEvsMZbHuquRt+8uE4EvSx63+avNc9EZjEphX1MaoKgC/8Ze5+zv
ltxP4quytJI1tByJZEF0HviiOAiuHpBxMvJo06Qaanny1eWwn79QoI2Y25dtc8aQ
+SpKfEtD3kDYH8UWxm/voC4i2PdWfj/JXV9UTcip+XCZvbBcqBUsMBzrYYrBb4/D
6hjpO4oeviReU1yANPBZ1Xc2WrX/ESVj6xcF08eXXTVSoIzFq+vJCZ5UOvWYC3bg
NoTdBQiETemtKaQJ9sGgs3E8rlcuAXUfh0TOzCMyROwrqT1GSTOGbj4P3UycbeN7
C/cI+njIN/zW+QYq5h7PGCaiEc2F6RnwJkLpG2/qvDeX0tWS+TxfGUABg0BXNXMs
BRYuwAG+b3gHko1lnWaQDARl7S5Jya+UA9ZqfAy+29aEyH/Laevznzv4FAgSNkQC
i2bJ4RCsAbjZVbUNwp/csgtRPoGO9AyNHtr7D02dmc/GO1piGMCM1ckVgb+Us1Ls
rF+OMXTUDeVejOrBW1HSE6q4Y/D7v1hOJlRFkGDhy54Ou5jLZj+K27sKa60J8Pwe
WQ3GoHa+T1u6HmYDEe90rML7HcmMcBmEM0Vdv7+xGKNwnFgrHoi6wMnsmFgNA7la
46W3TXQ+tF6mJXbGe3X9ig2G760NTdo9Z65F+B/T+bmZ1OVOJnAqMQmSSH3zHntw
qomYQsbjIzV+6U/JWgwCwKLk/gOHRZaimx+AwOh8TcS4HRDEL90q+VgaEOq+Tjqf
yJnusiK3MIPdGEEbDFAfP8n46onHEMcbmUGv/eo/Uv4OZQKzhTZqUp8PID8HUOnl
wVCNw+S/kpvOlrrroCTTtUqpUBobZMfgsIsZwIAmi6HTi67xYxKdTeTN2vPW03Vn
TIT7vJCKDK2Rep+BA40zftotExWaFTlCk3CS2VPJx5UvbDd3iqehRV6kT1ZBiOXK
v/N2a9JlbA9oLlK8CtYaWiyS1ugxp7Bh41S8KGWMz32JunwoxkXOzQyUQa46lzGB
/XfTjML8ZTaigB1+9FXJt+XSQMLxcWVQhYMRTalNWOavKb59iU6p5TURISs/V/VZ
e6cyflYXuOZy6ZxcmVKddV25YMfSl+d1hySWkj1CWn0cqsb6d5q/k9z5bbfrt5H6
zP+0sZ9r+Kd7gbtE3eZD/5fdsZB7v9MX4WwiujanaRNvfRcNT9u7qLAaQ8acrcG6
vkMRQrbNOT6lb62JhtF1YvZ/A9VRFQP44iyfiuD6c7LSEaEdQAU8Tyq5FEdcEroM
fxqM5EYZdqxFr8prsqeBWcVjjdLjObzeZKiQ5RFcYsuAlhETA3uwdQcH5fKoJLXm
36wrJovkDbEkaaNspVy9099aB0LekuNN9nRmyoqjzs77nOgUK8r9Zok6I+zDyVll
RUza/sosmbWkNFKZ9vFDPXrEt1A8ExtQu9cA3jrG27bZEgcB3zkmc8vJerfhSdbp
fbnTWfiBsmOtGKPkI9MAMQP69Nl90s/7jslpu/TqX6OkAyNrzQW4lX5CgaR6etzB
MorHg9SkOfijB2wsGT+xAtZq0mxqqf52loaOOo0RQsDDABpRJbdrGkrcBAt3iCp2
CSvn1q7oTFZhs0fd55MROP1S6iH1IOmObweU7H+AEaL4CghejCVEsAeuJA2jx7Z+
kbZFJnj1S/CRPOvXV+LS+RSFVg+qZWLwbuPNfQutsNUPW5fq4feLO8OdsLwN7A/C
3Gm7uwvwv9fMXkY7qg05T6phny3o51c7Lx77SLNRLN7QQ1Fnf6uF2QUg96MpjSuK
mSWbmoq++uFEQcfhmlRtLVKkEJUjVzuCT20UqPTuJ/yI44kR8MmSHSR0E+dNuG8N
gH21TjdRjAyHq9PWfJM7s9oEpTODLsRMHYReS8N1gy3/9jbLow7yDSYXSfWE7Fez
aX3YY9C0DWV3lHecGZEwTDC/3dS8FiMVIPY7vYH9LfhmoDzqAkaMVb6sosgD2TgK
DrDOgr279StvNxF/9oVa9ECMiJQwCEPsKg7R7F288RfcR7oLyqMXQuBHn+kYpXOJ
lh45Pn3GpOh+EHTyse8D27ENDs+h/N7H0B9fsBkl5ury+LZmqiG3sDTLECRfUsfM
SozmsDFDvL63pBWB2xXBITDiWtyqlW+CX2zqVZx+4Js4fcNP9hG1TE6g7pdKrxpt
y92nbHOLiKqHGiNc1mP+JowNDBKUTjCYaIV8GFdAy822VYYaPB9n7djoh94dbR1o
RAypzOZ9fSKCjkBA3raKeVmpBEEEu4JPiocjmpebpNQhLxDtGkrt3/0AA+nAF837
eekRh7lIlJdf3wdmctT/pImASdccGUjZrreljnIRJBSogiDL4OKbD9XSCNI5pXiY
sbzJ32/GT3GSRoFb6C7EGKT+Zq+VbwA5cCMFSJATmRQnWXLkuwUm4SKE/l1p9SlA
qIXzalBZF+8SfCKwJebfT83FLFp2bwQcRUMQIjp6b5DiCHObVPNsM07QGaBCrecH
EIeG1ecDuj10dF2GxHQxmMLQjxWfaYDzWMzS+/OE6PrzhWdFaUi3dlfkUISXExJO
CnuJ9FLaB8A5oMqvvcEnpmtEwq42nfr4ZDu21VMetB7rPAlpI1NIvDqweFSPqype
G0/E6CyNcqrbJocws0jrvOkj+wK3Rc7HzeBr43o7ka/pxqSR35jZDhz/c2UBDPZb
EOrjzodZUNfzFFJKHeYrQENMkZFxvDRF9ZuE2py7s+6DVE0QnLRs3iDqpzXtoYGI
sq58dhGJhRpwazU1y4drpzEHm1njgqweQh2N9RJH54qPdM52wiwEmRZHwzCS9s75
22jSoq3niLzeA8Diklupf4lg4NsMsO7kOsXJIODDb5dIdkSF0vICJS+acW+2koBD
dgkIo+dDRtHJRI0NOtHweeYbZV3QbIbLc3gQCXeavSWk9XBbjkUHO27ouAr47b2C
FOivTDKvoRxUQmaxoTvFgoE1lnM8BOqdORnRivP+u8Yc1xS7OzNuY31k1dCwkRA0
RhaqmAeKRgU7OrqSqgnwrmigAIzOaLxAc5gkez5jy33w59k7t/9x79QCPVMBXUcd
3Z5eXme2Rp8hw0X4IeqvZA35qA9OaEHrR6khl2UiYELrwcAOzRev2yXY2tK1Nppn
3LvXo1L1qi/AZI/hET4zUNuKv0DFV9xhajcTuJCMBArRd4X6DZ63/8vVqvJdZlWn
UzYkkuqCleCAwom1op5nTF+BPtXW8+aGP8WiNAiWxIl32Jj/3Od7iAStl98PZYSS
wRpA6I0xp50ByLU/2Fg+43MJGqGTgKuJVGHYD9FVVLoR6MU7g5jYjOWRNAKNL0jT
Lv4T7etc9C27tjkh/1XzN/nuQXEYtKdg2QU4EYEHxrc4D3XuCv68yKppKTu4H7GB
9rb4e3IOuns5dnacjxLILNDtVZh5j08PbkF6+emRh2bPgXOAPPFyJgYMPohkKtcp
jejvB+HWDxAUGXNv5p4Cctpop2v4suNjKLy8vI8AJhi3PAqjuptKl1EVHVeunhlt
zwLV77bleVvunxFZ2hO8YmxI3t8UJC4d31W+LV3amVThhpPgmyOjt7GreUS6U1yr
Ekmx5s1y+cBAqDpiK/x1RhoUMp4VSD0MEkiNjX+nq6AMOFvWeMqbrLNgYfP+FiCK
kL9ZGE76rwAknemDP77OTttoTBjyeSkV2hK6KCJLIbLAgi8aylxPFCDO85Hpigqx
VywzqkwkYifzM/QDOA7OUnn9Jso5qhmVrDLB643RQzPZ9RK9iO7oHqlSg0sWvQ96
C7yZ5bRIaF1rLkrRxbp1SueoqU4psAmn7NtQPyXBG3LB4Hnz70sqRgeDItVAufDx
bZ6Vq1iWu8lreh3cCyCBs7D24PDZ6no/mZWtfL4cy6/CceeRjk4SxoLbHFOPzfp7
Jc6RUOVbkOI4NTnMBqyHfMOAV1CerWF/5UOQw9gKVZ0PGtgQ4nHtDBZa1RzirK/t
U10A5wnXA/luDuMw8JI2pKRN8io49olqDWqihGjnmVegh8oJzUz7L42HZji8szCk
EKVaHhu5pe5jf4Ac7RqVhBiAM/9uVg6XbapNIep7FKHakKrQvLiiFWknBI0IkpIU
YL9gIDDvMa01ukEKwWtR9gi/Wc2T7ZDpkqXamiTyxFBPc+j7avJjfTJ0kz6Y7nVw
5t3q+wBe37UOYPd8kF44g6MP89MJ5wdvBYzrrIY8ULjylBI4zAfTc4ami189V7eB
OyuknPHxNNuK0o63J8npfdnpMYuXX5++ssWVN0KTaNlEtpXx/8nu09c0b0SJUapi
2+wKoFRzzCQuNEeyL8ONhz3UaGTnpqG+K2KRoaXDivsRjpCYe/FOiFevIAtecRMU
/VxKowUUoEkZB6dxzBCy/SkVp/BfI4XvBsrM/lFvKicVr7qQZ28J9iX4YucXs2Gs
7k8qXwvQElcRE1EoBcOAc93lRzWVEwxQfJv4iQTluQoh47YefTTHpA1lDdBapZv6
uU5okB3/3WQRGqf2F0pSH8pkWdyGepYPiCfENDhtip7Izg+geJ0fVwA8x1GmzlqS
OaXHY2iE8Rh9qbdbRGS8DRnjz0uZpxVtslYEnIgMsDcCQa9OyKrbZdysZuENqZE/
WaAafyRVMyC3SIyXdWYDYhT15hSvAqB1CXJeH+ftqzk3bs3tlFWtChnTwjh5u4MI
C29z0D9ivm463qHUP+PZhpCo9zzHTZ2+DqKWM7RGNfoCBMD2H61EVeBLbrsBPM0g
VU3aqLNK+8/Zk5LlJaikM0LjusTZaXN/N+W4ejgtX5CTvF4pV1+FzwFsLNp1XBl6
Acwe+oDV/gb+kkW5g7sJTiWfICy8RveOgQ1UOCBBFovX7Iq/6wojXjoaeJKH46LB
xvBxJsnXGKnk3txeM3UIJU5qqLGeO2wci32UhQA1xsf6rtBEyzfdehcucmBUFlQ3
BfH2ekGf8NdQ57fXxvqm049Rzi97pSUCWM8ZP+oJhnbNJQ09GGH4T3etS3y7JzIo
QAbBizgr2DNdggT8et1CO4Qxad+NzanX0WcFP+ZGnJkerFfDXGmp7t43HFp9QHrP
Fbm2meqC0U12rVgK7sWRO/U4tV0IZo5KH/8LQ4oWJ+TIvssCgQFDQwwK8buGhigo
R2WsBSliZIVUMkLdb8E1eu7z1eaMT5RnBHK007bjYz9C+h5cPJ9d3UvyVTVflOY3
WpdvzPHJe15P+FRqD2mW5npZkc9gqCmwnJcckmqmHjjuAol/sjWqDj1J0rLeTksT
qC4TEZ1kRT3Wmewwx/v1iucAbGr6u2eqXCIxP44XLCbDMKWt/LZGn0zR8ZUE7GH+
5JZZXx3/PNQMjY/IMyix+PvYgP/PaKeo/97/a/lfNDG3CHdHrPByoqY7M6l8Mw+G
AG9j9Uk8ULLtDOsGNJ6vNAMikoZFpf8/leuEXwaOjeu2Fvfv3tkAm5woDmdOIvGp
bu+KtHpAtWLnvV2fhfALHyk0wcwrv+jzdsD8/BYpLKLd6B/GW78AbQzEciGpU5l2
ZbDuQLv0A/ko5+SwDgK+Duy2E2K2WERABxXESQxaPcsCLFCLFzZ8BF/umpWdqEK9
xobR/BljCgBJz9zKvYn3MZnZXfhn+PYPjwh62gByNi4bsm5JLttLQ+URNn5NUFUT
gx7Tde0QNbCFqc5MuopOdFqs/zh5Tyr1ta6Y+CghU8CX7ZxbGv8d9wgQGVnx6ta/
KrlaQ86hzCZcH+SzNQmIES6n1c910lGFlmxh9Up3/ccOcYG76yf7pts9ldVFHxEs
oZP3k1jBUdnyQ1II3ZBqTN0Zu6vziM5SJW11mZgHHn/F9q8u+kqPD2KrgCMcuYIs
LSgIGdA8A94yAuQrDoTOZVXrQOcl+pw7oVrEbIKqRuF60xz+Qhj3b7B82h+qG2sg
3ucFiHOgWltB2Lzw1tKjdP5cj2TqazQQ9FGwv5KSGUTOS9ICELKGyPXvRpNV1ioM
GgrkqFr8BH26Z4UM3pYTc5BiX2kSD1IqmUXVbWzd8J28cv1hb5t8iHtgm6Kpzzu6
k+giKnzPB4QeROvRS/2NgWElU7+riB2khN4XB0hyMrxgYzwSOl1N+SkKsmk5pvky
piNL9pO8ok2Ug0gjhsmXh5vz73yi+oFFc7jeUZalGbJlIq1RtywScwbEei3YDXrq
`protect end_protected