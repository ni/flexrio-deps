`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JVISfbOcUocfAE00jf0meG4
/vEkqJfyK/81z5lf9X8oFYLgCdExARVM3sDjEKGfkr0J2cIxASbYi9Q+CRwaRPwX
f7pY0RH4tcGedTwOlJ2qToVRfArMz09mA5UNSP/lpDnMcdnT8euY9cnF4EVuF8C/
9FJwaiPNL7ggoZ1eOJADGqdwjUBfuDmi+7fm0iUaH6zabKjo+WqlERlYutSjHrmv
pUosXxZWtSXd2DWbMMwD563TxcQS6gV/iKmUN3628ls/3UMrAIuwi4OQxddsEUQy
ENWe7nhBToS9t2UiuqEgsIqt+cw+BOVC1M7VZ1B+YXmlspGQzuBZuGAFGiEC/msq
eg36ykadIbqbi77vjAi5z7ylE5gySnfTIA0GfLIJHBFIPj3y2P7AqcaxCuNTjMdk
4Lb6L/TvOHfXE6QINA9gAHWpACAJnVgxKPwFfXmMkAYIF/0BLXj3gDAS8Qs88iya
FUL1zWlXv+6qwQExtp4WJEJ1kc6vjz+Q/X7Vcz7sycTLR446gFfT6A8kZ/XIe1l3
l8oNa7ntwqWGSyANNhVZnA+UyqFYnvSNYVjFAZ4LjDLinuSIyNZDT5HtwFpGBJsQ
ll7lT12cUQTZlAPG8C2Oqi/UOiuQo1k9nSv0LyAbf5I7mL3lVURWhforbMcn8rVM
KryR4GOweFwlpHSekdLKKyuHyVCk8GkRVW4X/M0qBYvbfpszDz/QqmBJV5rEq8XG
SgtJutwl5j4WaCFduYKQSdj5cgbcT2hBW3jVgEnFRPqfDK2FD+ABQTmiiW/w7Cta
LjdDlW27uGXn+mtdMC4MJG8sr5jXvtptoXbeY7EVNDZ0Q6MlrMKPjXpULt0afR57
35Tn7jOjqUqFpkeO0AV+ciOjc4f395AQNJpc31mrLJF5kgM7Ht6aT3Ym+tg1h6iB
/uNhPT4mC55oOAFvA9DTJXdYIb6erfOLRs4dmPTEt+F8PsbC9/PRLNhD1S7Rjd9a
lZ3syg1FmbRhaCxmDzMZmAZd2anH+BBhm8GWtTUW9lXhd3CU92M5zLEBxGcaWYvG
h7LU5UjR038qLVMyUSVpGxlNynNA5ZG4shSN7roU6UwXqt0F+ffkLYxnpWPuizkI
q9W4raQ5zNWRrMDb3FUoY4c+RWHbIK88ff+I4rjgEsgJpEAIvxFx0k5B1xwBA09y
Xx5rYjuM8UcaXmGvTTGquK0W8hursxYea9hwrPQOgc6Vf7wxlAzPwfLtREqJWjYX
/UhTqHP5K4Br04bjue2cqftEg3gZmY2yYvPbnjTvfn/DP/2SNZwK0JO0lYK3nvrP
t3aIuR5Ke8xNjH3fpL99ovfVKNy7x5PUxw9dqR57G5UmimX+BAjKnooRAFGybXwZ
gSlBG64J0Ur1VAE0v9d3s8Rzg0t34i0ooZ9RVo8/LY8NJ+ce1JTOpDzhnOe0uaEj
zkbQTSMl8fu7YLiJpgw6TDJfUrYz6AImBWhhM9v9GOB/TM33qfj9VRKRNqfTuVlY
8FzL7l5BPvMrFTkNDQu3LJjGYzr5STgft/M1BTLMJEr1tINQYnw0yEAusQVsrWqg
4xXCo10JII2FejUz7khl2XWMbtZwG+MCIbl96Ge3YANZ+iUvBTybT6Ebz1Yqtduv
RV159hDTAOmhcL70rKP/BhElHazx5/HbUzSqscskDsCKrAq4hD2XLViGkbvqPpyL
G7LZm3HmjSvsRwCZlvi2IWamZmhGQZmwLceR+hKCYwtKMVBnuXKZdNTaBq+0L33t
b2l8/6xe8ARqgpgyl9d1K9vut0ssdZVbCqJooDT35ksfKFHnzoTvt89C4goV0leI
rivBhIfQLc0MgQamIQmbnTAuBTABsA1KfzipLeFkTpvATVuqhgB9XFgmgeCImdhK
wIcKuvG2Q3EGxgubK7U7MGkGPxtQClQPAZrJ+oaNjulQ65ZOXNtXly9oaurjRBpQ
P7vbs9arAD53swxzRufm/eB/ofSrO/xYyWx1RS3zi6qameLtASMNvz6ZKm5LwzID
TqJNuzeOet7QHnF3V+IksDmMDlsJSmgG/E0LJ8rxIuS6ZEEyuoytHsVPZk9GZ7Jo
qKY/f3lKAdguXiKCNqGuQCyMnYK7ZXJlqVeQLGQKM1pKJXDGMnlUIZc8TTW9uUQo
8UtGW8hPIivP6iRndr0MrZYKfZ9vUvinpWlgZLKHOo7hqRxlIn+R8C4lO5Xvl9L5
Ax8q8FIFVSwtKjpnWOKpuhpCCW1ax2aTyUnAienh/FyjS+z7n4j0DJpyYlBL4Opf
Q1usKKkMF/CyAZM1rDxqRvc11J6S5krVY9jSNV2NWRKBPUDzgwHdp6EsOwnP3nEK
uO78DYViYUANFhVEsoKc/yTtZ2o8RZrr1y692pCNX2u90YKT78/8Q8ebL3zRPsAU
lw1T2tWcXs9jm3kuWRQMWEOzaquxawDnbsL+Cy2+hSab1+KyoyGuEo6uBNxTUlbA
CdcdyLMiDEtqxKKJ6pozhJzlMpm9WKEoFmZNexFYSlk0zfE2DlQaWfQQP1d2xbe9
E2tT66I9ySeSV/VPW7SR7Y8KZodJU4M/U1mup8xUHxV0Ny6RWDOvtk1VPOOdysuq
uQqnQM9ymQxz+fwut/Odm0MDUFK1KrINul5AgdssKUDKgdVFsBLrluLIu2itlXt3
8FKqgA9RiQvAvEVRLExf3qzYonycJg8BZAcLXJlDoRAvcljcpHuOpEbwrrjE6fxe
dPVodWerdqVfsuVzC6vBKw4Hl8Lrb3yZ1FDaZUzYyjzc8sFR9pJEX+PI8VCa9bhF
6o+Ea/7mpnsk49ImT+vii7+Yhyugfvi6Q3msLOgTxJ/lQuCQlyuq2Zp2GUD8vobD
r1xBWhceDyQysDbMZZ81uqI67EteYgnTY8kyxD6X7zBrm2rJZpS7b4xF+3hNxcJR
Ew55Ny3R1TJWv3r+QyuPhILzJv+P1NHm3EgXbzYzfw7MVLg6bmTePsqyZEysISP5
l9MX81MUY4BWCbJkBn6hjK5EDeKc7+VRg3Ha4eTLHxMgtyaerb/HLXL83dDVIAHb
OKRyqFkKa8FdPirxRs7evAth9eFQ0Pel6A5MEB3ITc1YjyEuu+FUrBq7TvBnx2Uk
g42b3ZIjE0ThcMIzp4ODE9+VblTEWsbujGv+ib0wX1LWYhYhhpvTng6Dj67qlac8
vdlYgPHV6N3evpShhO4gnBxoanHcVRAgya1QPYgjNyZH+wJSIpmbCx/09nbpG2kV
DQxm92dFF4SaRdmE/TrF/fP/cctuE1MGKOFHw0i18pcTdvggP9jnc7lTi8vkkTMU
APgBHLBaOpQBEoDj213cQiIKjHUV/ahrbZAl517yZDB0BghJiRxGCnztM2qtlw1L
WoR+Gp9Ea6lJ4ufagKaO/GbPHfxug+Zfa/faM2fc5ZNkOlw7w9pYDq5sbFBaWUVi
8baLS0D6sqJFF56j4CYSDymr7r7D0/+yTvBdPhlfSjzlYofVJucCyf6EQLNAtWkN
RZ4Pg0AWK6asfUCWvYv+uzWTJZumnWuSs0OVxNAhVa78QFzRCwxMthenCwqnMrFG
+iz1XmuMNz8amnOd8wVWRv+ZH6K6vnVRUx10q7EUTewXePKaTWxEc51g/5SDvI0j
jFJiRMEDzRozfKRwLfJ06cLSK/Pz89keUyCjF+pAzWVUXYLjhrW5naY8pT+ZEKDA
FrYdCCP8cwdKx22rHggfWrZnEP7PhDJLx0zQ6K6RhdvlH3qIDzTD+NnQXmomXMo2
VHW4kNqpqhcwOIsnTpzdWQut08JrPju8wmQ9zvSmMsMaIZHpmaWYkXAhhcZN29w8
6Mn768q9bWNh6kYgHkOsXJIK0/h6eDGGIwLqzNgHGLEdU1UDyOuHQB8+VywEmduX
mGA9SazvP8t6SotLy3DSz4FEtiN4VVYJIQgzrImTPUzf3TE6zkybkf/ANFcIlCrB
ZlSkgulVDil90dEj27MBogdTEkFWetqna1c5Mb8lHhmCkP6NzboEegjZqIeRXjuR
4sl6XtvEzllVyAGRh9Ei954QZdV1VjhSejT6dC5ggAtS8VbrKntPZA3aGwfJNeNr
grxx9u6igGvQ79FgFRPHRa7J2OvDm4VZVWKHNrGrl7iZ980Ds7lhNOFHgZUEezFP
2MUmZlGqLHLxQIpGnd+WUNjQ0IYBTfLipZvprksgo4uObeSjcWa/NaUsyZc4Li7D
yGR79BsdOSCdp06jxvmHucjeFOHSjvGWnnlJRtIQUJ1vfsqTivh4qa36Cbji7Kj9
sJ603nQ25pawpzPPr57kiXYfmxqdZotnW7JHmfCswBP7ElTogG6sZzrAC3dqp9dK
S0T6+fXbELkNZuJz5fdkg4MHvOQAYUXmgn6Kuq8R7qTlfFQQk14k7YAE5wHQ4xSM
27Xu6FVisfQspFGTBLNZuOnFwnVOp7ycD11NsJu8Gj/C5zg1/aWhTnBrXKlrtu9l
zQkMP0gyFa2h8Wm/vDqe6mI8VBGGnbTuvSP5yKKn6BoIc7mz+cN4bYl5cog8Kjj7
9duQbxY5mo611boufNMjQk2acZCStXZOcGy7LKiq6vpikY6J69xvwBr+sebYaVa3
IRN4cO9RUYkdcpfCjse3Gs3nUL6n2x+HEFSv4t7K29FHQrUthJpt+hCKQ4KAMqs5
dRh6uaRyQPge+xSi+izgYdrNkh8JeNc6dkZwl0wFDiocLq06ieO9+VhwK1419ZIm
Rr5WMZaMERdNrIQtIYR5bwWu+a+zss1ZKi0l/QhdTdH/iYEbHeTJvQmpC+MSVhVo
ax4wIj3PRPmRU9UrvQvxa8blWxZTttEIRh62cWdaEzTi5xq7SjwoM+QUj1JlHiz0
089bzXRrfyrOYyEANMuzBDKMx2lD08G0NE/cZmNN5P9oDWr2E8eZMQXU0apvBvnc
ScsKhhoIK2yyOqDilV27l+AZMNK585r9tuxMRepEPlnASedDTisO57MC9p3fgSmP
AMrhYn21pOhNKM+XSTEIssBAacd/B9enayk1joHp3CVHYpEXm4ha8AM6xjH8IZRl
XTbIqjQfEcp1Zk4ltQPP9SydvXTJ6OQJevKKH54XLfPk1PbvOrIWfmi8LdT68H5X
e3A+atw3U7pOlWT7EZIX3bmHV1P/N3vzFb7U3nBBGQiOFXVFvNDOmH1BfGo5ESb/
g/D/mUbSOmCIvZzmNlrVAqI9poLQRgyK9oBxyDMRp9xgtIW7nDfn4S4OxH7FtgOa
rqzF+vhSQqL1A4I9wqA84gXmPsyhwaq5a5ijnJg6cCfdh1ryz+aXxUwaD+s3Hh4B
Le8NNl/FtXQHjHfklkJyxW08N4UNGseTq7XCQUs+puU4h40eEct1wfynZcahtUHX
Z8phFidqwsWiF+9skhuHTJ/oCYZJ1K6Nv1yDXiVZ5fO7ZBM+JPbzW+F7vXdMUmF/
uVB1V29ld4e0fUIdjqRJBU2MnAXXCpH03oGtPEY+O86vUZjfsGw3VQE3/Lp/ox28
2+flyfc+SJi8zlqH35o6RszELMaCKc0YfLP7/U0UHpuVVRX+F64O1yMFUqV/dZ2Z
n685FDr/ENiH/9yAEbO0P15gpfA1uEk8alqEJs+RvqNi6oPG0r2CwjbaBt3vS8+7
b08+G4Aiz9W+uVotJwg6uOttVy16j8UWsGKv3Xoj8IyI7dA5wL3gt4jVAQHuFJbT
PPrl+J6X7pKuKmynqPRKf0EGkpB4UQu5wgfsu45XpiwpdAFxvQq6omYKgR0oQQKg
wpLwnmwwIm1sABf4CmKZO8epV/H1WndcqAZchulSB7/UMM+5rKXnfjoptupywHCi
yFOZp4MwOLddpZx+bhGA3gBwvQs3Lycj1q8t2xdFn6o8buZIMwFdSuz6CB9cZW8T
6jnj8VEPU1T1n9H8IS4aiaJCGeIFHmhW35X/M4OiAbv6pb2XdX+6+kMAx4GEoUPH
xAjDFzeyo8t3l7hMHfblZsXlO1CAyJsvkDVz1GFpozb12jLq3ZwT2QRyzQ/FgzOs
GH7TCIAtGhEoj0f3KDJ/hTYS65scuEXHSiECNkphHC0oMkNXlYdONVISV+7WupMu
2KfHJglS7y1aSXrDzzVFJQ6g6lNymBRPwxs7+mkzV6BIWmaf2fbomu6Iwj7E8K3n
PaWvuEHMdx/JHSR+5nMFyhackXkB11eU3Re3kCyrOt/0xO/gHc8jyScRpIDOmlQT
nmCV/jTrWBR92c2TRu/sJUWG43cMAQYuE7wLTgtyt8ftHV+tIfK8KxR53xQWbAmZ
gn4IygQlrh1JlVG8HgljuHNCq9a+d6ajqaUH4owz01/b+dpdPLs2CRUReZkH4/vo
HbMduEQ/9B1mwnjARTdZfov6JYy91edB4zLt9I0G+ZxTiEsoJmMXET+jWzcmvo6m
Lh5jaUO2ALHdeu6bT4O1XmVgbUCt2fs+ZCIkv6u762G1tPvm0EBDARFHol1u9LWd
avO6S/3BaE6SzMyB+DQi/pihuMCTRDn9NND685nef/Nf0IfDUYsnw0ZQSEQc1BFD
zg1y4RaMm3Nutt8QGA5TTz6xoqYpqNk6oiI2eibRPSVPLuDtDpnYZzMZk/u9H1hJ
q03WrcwbE3h6RT6Dee35PbLu/5wFMPqZGGEWN6ZBH16GotluE5nN5v3YWLgkKTUL
+AG8hVoREBMozipZ06y6e62oxwDk39s+k1yrp0qWnmlxPPejEq0pOMsdR2jBIBfO
dnAxKZ3CtObxj0Ct5hzutXMIyWvLeyxSszFGRIwQbb9eXui0eoVt+x/X7R9LnzFT
QQythLJuvqiQ0TlG3xQYVeU9w8eE+HIX0o4vccI46nP0mIIRV9jHtDvzaAtuelkl
XFz6RrELc6UaHtNnlTOeO+NlETwTVy4XV+m+DKaiQW0AUuQVA7vX9iOlWuQpz0Ff
uAw8N+vH2BafdsUYr3rKJ1dE+W9nJJLL9RmEfG66rwTkdP4LWMjylrj8FFvoNMDa
nNgiJSPsQotffo4R24SDQJMd4XZdsF8J5aGNW/+OwMFkwOwUp42Wg8vZO9U9GiMn
HNea3ZvLvRDmgu65mpH11hM23WITk1O1DoGrMAXhFzQSoNE/oeh8h2EaeuALfr93
pJ0T+TfsLliq/CqGSz4a9AGMomTAj0pr9PH5QjRVrsu2VjsiTsbXA0XoRSDi36h8
OTbPGSR/r5rcyglUFpD9UzB/eJ4kvA+Jce54Tl1GWYsEexGs6Fy4DukqQMksYePN
wTZm5nR+yu/mk+6qecAaN48THu7+gMoR4utgd91kPeBUpKHwI4inTbJsvis4lhPe
3DyYxDC70kSb47ihY3nnldWLZHPZPZ3vp48b8VfVwRgMmEoYU7O+o7X983/wLRxs
qFK1m/uWUVPbfScd6R3SSAQ2QxUjHh+I2OWYLZ1lz/wh01Vq03dO0NzYeNDQc/Ul
X35FV9V2bZFwFabNUW0XxqMlFC+CnEVAfUqpLnJFDnA/URtJpLPJF3/2uDHZPa7i
5UN1JMcPB2EG6I3hjM6VTofXO27EpcDdo5A4EECKmF7G/ybU17p8GvaDH5lF9MhI
myYW08GpvBOOduYoYbL2ArrNoRdo18Q5U0gMnTeA/uwj7Z/u71FeCxe/ORyeEOVF
iRbCDp6Uy+LGDl9PU+GffGZShoc8p4yLcDPhc5d3V/J88/TubgeUNJHJD4qcfZ8X
LXFOseNEG6rrSHSIZtaVlnkNE+zD1gV3BX3+golz9rRQxAbRogU37rLdiJn2T2Gx
T9nhiL4V3G2+Aj1juGTtSRqEC0VON8zhr8UKLemFumemtDZicAtTB/hO3039Cm9g
i75kbaLQTo/5VuPBiouhbWezOt1xOd7wWeb4lszC5CccqQ+4g3kBesPocuDme3EM
rsASDbdJTgzpBdvwiEgMm+bH1ra9F6tDZ0JZyAnQdlougts9fqLWzTZjolGo1cLw
ztnPW8B2f+TORweOdoztSd8cvyr3kSwI0TQ2nCdRvcjFZNZ48p61A7+CH/rlEGYc
678jc3priSosiZmKqY8L0o1goK1JsVrIZtdJBqBCipgol2+w0KFEEN82ZitgvGEP
8W13frg8fnRrSnJmiNEQLVRUR0sxeJeAvK4ajg/2AjdpwIyTjW7n+hDindKrUwP7
yFr9saMEJ4m9woYtrzn3IFrVjAX16B7+n/EnjwQhFcbiaOBzocUQ+gvrz780idih
imncOLjyXyE4kBZcsyenqc9x1mUSIb0vZyMD+YaLoBE1cvTeBJzzM7Dw6kNab5MN
GQ1ao27/+L2F/9UlMzafLhzuZzRRRkj8TNVPJsaPn+ycBXBvfFqdEfxp3uN4a/O9
V3qW2vWmNHa5jeRwB9nS48tudBznrrXkZfRe4hkXsGhMD/SjEMz2sOqZGahuuKN8
1SIb0Zc/3J7iAJJzeyYvzaFR8z5JzFdGlmQX2s8nCy73xcmUdQCkgYgeVjE0ECfl
guQSbVX/PGZN32qqUrCJ5lUCjjF4a6aURbCLpBDma0UDbvw1vnbKzqum7BgMDmXy
FTc+ZVTfcnr77+EIUefaN1wJ0Khcua+R9v/6a3l5rwWFznPKCY8QhLVKt4JgNrbT
NET/wQyi53TAFxVzYWRE9i9GTXW/WnC5vZZBpf0rfakyoOMZUoyerAWhCUuI+MVk
mawPOs2sG0MwjKMerrwdVyLe4cBRpFIU3QXaAM90SSfy3iIJkAvKE2sJP5bjDF+C
+U7oMZjDyG9PDx/vb9QHpgBBdw8Yhl9aw62gA8hPhKO4NIAai2TqxiVyCRIZStTW
T/NESvxeptZP/BmAJ0JIoUPsfaX6SZtVRSiiW2YvthzdgNFizwt+qIhF3UeHNFAN
5bees9wElX4sgYIEXq7mF0cVsrBDTMDuaYei/Amzg8nJN7VRAkMYk75XEN+628Ay
pkPsXA8oSUAxM6NpQue5HT9cyr7yH73NPWcx/Y34b7KU12dFyLnhKL8iSxN8ncV3
EzDvOVMS57ult9agCHh2IKIA6IjWoyhLPWyDE7/x4qflEhMO22Gr0hjAu9foBqbx
549mM556iqq8WAcuEOYKAFgo/EqiTVXy6ZJ/b1OpwYlO1P0p3HFgBS2wTJjHMPM8
TpyzkkhPLBiEhARZzLYBNhoCfEb/eIbFKUsOmaONLqUdbR29gMtDYZnA5S3EA54+
y/Lf9/gOkJpSgqKmXK729somGU2hu3XUQI7ZDRzyCvQXDg+GfEi6YZikQivIzXLa
1KD984Fk38VA1y48HE3tja4BZi5oAwmF30AXfwRhRZFQ0qNzh9xZo6ENjylx5Flh
Qe9QdsfYSnDzkw9WqYDMfIzFOssG3Qnb9P+OhYNbSUnj42J4KIJWCoiNwVouV7bT
ogqqgzq/FZZBj2prhfbgKxix12IK4pTPdRTtMrAXKYjYeNCH5GPXtkdWdwo8G8oi
YdiAflBVR4ehNXWxEvHRVuwhuRtZvjBHta/wufbIRqvE3i8oSf+0b8xs2fNJoSnt
HWTo9Vgs/5Qj2qeGQrnB8h0VLPogCuQP30voSLrjyxuCBudX+Lne1DHtxF8YbnLP
bB8OZznIiGUGmcHJk6xdYBOrXp7sgtNW9symmzFsTb3VVjEOsPNJI+dV8a62/g9z
VRq+tn8MiSa3qTlchM3PzdaxLVGC1+0Wlq2w5pEtU380Tvg/wUw+WudxnnCNUYFT
Gqi/YLYzf4QaX2bpf8meF4C/ExAC6Z8m2bdkqQ9Pwib3NrXJZu65MGEFNnT0OXW8
zhiTZarCOvItBQs2a7dRndxIzWZYSoPO1zQVgQP884aLNG0RkUPyIsrHmkWpuhty
4qqu7XoyXhZ7+AbZdeXzY51WUsYE41bFvWL7h87xzgHxVur/5Okjw9GH9z/bVgAY
BTrBaq5jf+rmTLLc0Rftjl/XkD3cQ91x2oS+XXjQjvD8Px1R91C98sWdER6z+EbO
MSbmgr4CVaf2Jzvhc6MUV5TwN4j5PxbMMS8QniX8f1wxfV/XpdX09/CsHBwr4nTi
McMWnoU6Gd6/q+uc3VNYLqlWsH7yFUkrbCUcVj8N3pY1rfzfWOep+h/S5UBV4LIi
J2Utp2WT13ruHZQ5jC1atXUwmOA6AtuQ9PphgJl1uNpsNLR2Wew04RCfkGIlwuC8
8HiM+PXFzVpOwByfIGanvdvrljIvcoNmriugkvlijmZ90YCggciw5sYgzEP1inN4
iUu0gs87uMhIu8aWZDtXVjN+rlWhAlI1UDl9iIx1NfVpQthLsk2eL8fIOMpN/ALy
kPG6mUt12WlcgQx5L4FnPIUFpyPB8Bpl0N1dNBGt6Sjn/0rb9BiZCXsAo+kBnDAL
yuOsFLQa8+U27b6UOJ3i0DASmpGtmKSn5O7pCOHHOItTeV7s8Sis3O5fFKQSLKny
RGcUmtJYSiteVKTBLfP+hVkiZQxl2FpyE2yG0244G/02dA8KAXejWQjEfwQuS3K5
iQtrChdse92YS3r1tyXRIQVQlpA+Viv0iPFcQiNm8ATx5CylTOarcWb/E+bU6lCF
oxaK0dwEdzTs64xGihdchthuwFJQSW0UjOu+1ExL9cwvdg1I56acIhAOxjB+u4+g
NVBNxMD7JXWDOd+mIYPtnTSAKcXZkqGd3nvqup350wLr2JzwWWZjOvIKeGRV3GRM
WeJmdK+Uy9UL8rFEfSA0HR2HcUjP4R4K3EF1q5knFK+Fc5ApnDFVBjHfFHATsgWa
MzupQabCm0rmnF2ZUd9OQbgRwUDOJ3BCxKvkweYk1OS2KtFwN4L57kdRc5/QBMpK
hxuVnK5FhLiXLstUJRdxDzZGQIrX+CrxRHBzgbPdpl1jSuPFKaWvqd2zEDHwVekJ
rfuocpluXrW+cVlSYFPIJ/Mg/uaiFlu0MuGOTY4+9QGK1qWBF90T3Q1B/KuKwAhD
IQ/DLZzu+JDBldmb85SOarM3Aq6ma3BE6HjvJODQ8YI52wtuxnd+/lrJwnZt7480
+kprqSl5tHJ1yXFFuVZJryl8M6aufGLA0vWgjljrYQkY8BFv7m3nTIrrX5bkc+id
qR07Y/v+ZvWSR/AvEkajQs0U3Cx5PSAi1HSsvaPi2NPEEi1xd59PMx2Z+2gH99Yi
kpXnztzbJfdihcJOtzrD6JqUsjH9pjyTHxvfdfTtIhgqhZ06mu9yeWPmbg2mSGQs
KghKAY0ecq26tEa79ppa6rOA2btuRYAIsOWqrZZZwvj/zYFcUJ3WsqkawmH3fTo4
duC+yRcQMStf1URFIabyA6nqa3WMjT893M0f/6DQXkk0WmqZuQOmlvhb5oIEPmgZ
pP4nApfxxTUQomMdivzrCBHZuTykBWISJCWjhljB9P0skjlwtR9wU0xZohJkAjQw
BC5rk4vpCCObGAty2E/tsVpKimXO22wx8msa9IjZ6PwDfygZ0mbPmhxG8djBZ+qS
ODBHBPrCMmQywQM4pP/K94q3gE1J+UCxQDsg0n++aDuUF+CKwdkv1CzvKqUPnKMT
DWTTmd0/swf8xWD5T+eFHK7su+4WMrIfvDaaauYvBapwISRzuqxtMHpKm1zIBZuI
geovBsxTXAU5lryz8cCYmBQth9TXN55YKF9+l4rLa+p70rXOJ46p2dYyMpJ6NLqP
zDCEu1aWdJNaL5sIjn9go5y3me4qoy1p7tUlCwDKVt3UQ0sY9A4FaznqH7JYi6nO
gB6TTuycOFD8sk+0VoDv28cQnI10WU1H+nsZVFMAgHSFjMAOj1CIr8SWWniWpASG
ZXSil04ryzm+/IgUmKC/fIjug9z5A8+OZZYfGwK9ZLoa96impffiKlYbALruba/7
NP9jCaRjadXRPIWLAjffPaMcalbU8MpLUNV2XiRXKe+GxNpHkHeCenoS1Wnu1Jd1
Y0YmhOaHDmav5Y4om2GMdVSnFpOT28GvlwUNqKhjD/rXe98s+o1ucxjb+W+TlQnR
/bDvrf3HODrGmGkjdqLdi1EB3RoVJZapneRZS+fje1WECqGSoqvPC82U7fugH7Tw
RUk+2aGgu4DA7tAe25FK/rCdZA9AG4xBKOVD8Nn+BbYc0XUaX7ffUZKjn6n3FiYP
3DKWF2U7t5IxNbnQ/P3lcoW8pDDLkXBqaenYlhq9syCh5dDDTArQ/AzkOddRDMYJ
6m0V6Xl2HRcryYXtyGpq15MkUaYPN3ri/pyktyaxNIpuF3F8BjfIBObaWXQmMkv5
FciFLqUW8Zw4dsOK534e3KswhIqR8BIHnj/RBreyf/4sZe8nG01rDyjbiek24wLp
fhj2pcaIfhhvEu0b1E4vcrNAHPsywWxEs63yvtsUrxFquaRh39k814u5nDYIUHx7
xE4G4uvCAmnw4Dvskc8iYAFMi9oJz6Z+F0Ol0ChWpPDr2ZrPhr2VNoF3vspdm0Vb
Hkx01HGH9cr9uf0LOkSv75vRuP6M3pMDSkimuUqWUYM+vlbxQBsXXhl/MUlmmuMA
0R3TpLMIc8WoEAWNB07ONXFtRMq+unba10Qjg5y7nirAnPouLXiRuQI1bweDlNy7
yKZ3F+nG594zYHYW/zYh9vxscR3+Fgl1WjmDs+zTtGw9sZPmhpxnHVUYH9LmJWlo
aJhjbmp5nYs8T3YuRoV3WkgGIEkhGbhRGW7z8QJJkxdhfjTVPAts2uQV/CEaNFul
4iB4YJ/8TLT7mK6x5FEYkP2nqDAeEvP62MuO+BAHtsiYWaTvee0VL9XtQnJQjJLi
iUKxsuDT8xeJ1N73jL5eBCOvUUIBJygg/oTa0+XBtGMR9b3jnPUjcgNQR9hDxLyP
BV7/hWVvZ3OrDGgmcSfJ1bxsznR9RH6x2Wjor3vCVFup4om2t63jAQXtKa/7d545
BOu2WlxQ+4wQtGwIH8OK1QqwpCwXuq5kwY+2gnFLwtCu2AcDC38SBsw6A1pNiaTd
3JR6vwFNo/RrLkgnGF0r8D+nJE7fav95ee0hDGRC7lggWO3AkcYqXp8ULBVBEuoG
ybpgd1VznOmFa3D4AVqPhKFksmAx47Ebd+VUTlyTBmEJIh+vpovbUFGVSDmhaeIt
Met5zmQ+hHhRYcm8iMwdRLVuIelKXjiVRQZcziA9UFd2LWs+oFj6ZvYJh4C3DVxp
c5pCQcUbbhL8dR6xTGUZeQCGV/7qDccH2CLCQhAxD/kteO0FNZnqyq6fUkMp7Ei2
Qnws+a+wHHtbOcv6QPXqwmOiAd02xbbtsagp4a8UhYUfPcvfg85XtH5qdJl8j8p/
d9amL1buMMSwp1pvAL3yWg1W+YeVxCg5IdiGVa3jZl9uLWGDSt2/TDiwMZoUbfXi
Q6tBfQye1yyx8wmXEvtL8SQZD9XZkY9FZ8jNnDGN4+i/AgW7xdb/bOsm0qhPTkEC
jv9PCNX1+4M7cdLOS92RA8XAfH0pSKcfOd36dN1PNajskES04lNpsFcKDV+fNLvh
okF8E3wJdcfo5iPQnF2IVloJElvCCLyjP4MWCg4LujC5BEA2MGB9dJU+5kQQJjG/
Zp443lWAeF3pfPur91lzlKJ0TMlCxWLQebBgF5Qs6uUCVItNhzuoNRZMt1jaeJna
Z6ZDlaXp3nPngWvuZa+EzT7tWtL8lzByWZ+p+jo8mrln3SgzR7SlUXhsSIjAxeYq
uLep1ig7F3+7rJtKHPvBGxdxbsXHuTdpiMxr23jSWmvijslD2duzFLe8iolgvk8s
L4ImLm4lUNxst8I4mbfkHQ4Z1EpYmQbaPR/mjszoHjU0ZBtVEFET0j6LjWeas7ri
da483mrSrIlulbZYAWgNuUN9X8CVT82moCNNNni9Kx1teMcgeSmVVpF43Yp4JPzq
4Re/4Quu9Pg/AbiEJnG6y/vKJGHZ7RmtyjGKuJ0L5bD2+jPEfiF4TcL4AU1tM+zd
T5d+lqqqWd1qybHdklM7Q4nxW8kUHIZ1Is2jfaQaU7juNwxwwIQDrnc5Iqxp7TDQ
lXEYf7h/fyzienwmbp2yLPNTdehgRkAK7f0/jZJv26og/yLI0DsxaJWK4vlOfhOr
zu+jvc2t7XTP+Xfr8GvvnO/RwnDSNI3/lNdPmzqye1fxtkCDqodvsjmcunLDDJVZ
nZiPaKDUzpD/gdUyrQF5nqJDdoe0U68dtiSmRok6+M7CDyZMcfbu9eoFrZqzotlG
p43x4RdbBzetdSyat3yRY/nqItqePXH90inw2AzhqOHih+xhUQ6KsW4m0Qm997ym
IUzUIk7Z/yTxLx8Ge3JhlIlQ/l1O60ETx+sR5qeeafBS272XqX/CZlt8o+NcKZqA
g1wC2FsOEk0A4R7o69+9wNUXtSZtzkLgAacXu1+v3Sk2NeZP/OLJPgr/w3Zp28yb
Ha84dyblJx/exAEDRfjTIfctts1g/basw207gVvSS/Is599rrgPrHMfaKOjklJQA
0axack30Wo9jgkIekdCavkw7ybh8/M4RxXaO+ThS/8muz+7ojnCTf0/FOCMNd/9x
2EAmLjyrJB0ZsCnRn0tgitvCsMDf5kC16HA+6v46kR55vb2Fy8JEfkb8vGby3xU4
brb6Ynrnj8ITYQ++foa1OqF7K8D0trQWDxhYdcxOg5+In0eSf/OrOEEZ/7rbmdf9
w+Hl3hRuocGwTlse59tvMtHDutNGPI3o3sePtcWtlOd+OLbnqepcN61rDRyF3QRo
cMDeb/yh0qWAXb5uegiQU1/7lPU02ZmNUnfMXbeGFTew3IIcFnZe0AD21NRZwoXE
AWTwrmO034T8+FqL3DtvbAuGj7EOzaHUzhasLiOZGMN4urstXUTLabhJhIqBDHuF
iWgItAVtwhAUz2W1F10isL6nkpkEXmpY9zP/stdzL7PLnDPN++33J4tl4kT2C9k2
d4Z5xs29CYhs5BCIhA8iu7d6DAs+ye0wr+BY7K2sB6VD/uOYnPyhp01Cc9OwHYDm
vVOPgxQAe3aD8DLQzMRNm/H6ybPUySJxrteczXP0fgKHc14QphD1lSq3I2o30Rnk
fCoo5FqbR11DrWLI538JzNrr4iBUd0lYqf/yfHGC591d1Gals/Fh+Okp1NG3af9q
fojDH22dKj+sibS2nht7etsyEVNKVyoNG7S429ScFhYw+O8yJ4eSQD4cmUluTKtA
mU8T4BpoT1+OhmccsIoRbn8fOs7mUmheU6RrGnM3XITB/gXimTaB+tj2mW15QmbF
+SdzQozlvIJcxt6RWg24LYpak5HZ9hhFtFVp1bkU3OovoSbsuREILM6wkQTkgQko
YGhnqHm8XKUa5CKVSIkkFpooVDyS6nAfWNFc2e+NcVelibsgYfo+vNBpcmJTmCjO
ZWV0Mj9ZmrBjONvu6rEwkqBHAyDwq/tLMx0FULX/2a6s7tnEgTUXrmADwHwnLFSW
T73c6JlBYFbQ98APR7WSXihYhFu0uaJJEI12yHtQIkubab5MnF7k3W77dsQOUwwB
AYiugkHWwPJxJUAgjL10Cp0vow34toUXd0leffFeopUKnBeqTYOTcJY7Rs+etkuQ
Jd+GDuwp74qPltQDJLtTW9KujMw5B1BlG12es5YMX6RR+YG2pPapuTT6KK3YXwQI
rIq6ikZopNkFamJEWKPzQnpM7bUo2A/LSsX5J1+4arTLwzvJ0ETyv7o2WEw1tY8g
jP27rJQn6MwcLFWUjwr8aUeVbU/S09q/VkmmwO4d+zUAGTWJ89XVxejVglDBo+UG
zyuLKPBS4g0lIY/6k0JdN7nx4DEQUk8/1h55TisuM+O11k1phpgf96esERJPeGJb
SkXLLTxu32o/XnGWSbdkN9cg98GypVyFY4OHOTCsEGDm9e+Rd/msGa2+ymZoqYnH
mehFGFzol8rQExkaSRKeVyt3Riac2Ylp7xtPv9Ix9WZm7ykG8Pgaj2l9A7j2LMyd
sYBIntEKSCLCL+FzWB4pHHqZX2SCE+4u5OM41/36B71+xEMRpFlbvNHF6eq4eeRU
nT6FevoUeTMQ+np6uNLWvdrAP2yNBM/RwTqAUstP4cDQ0ZiNlTChFxQdNVoPa8Iv
FPuFLxYPNMj8Bh7qmjV4DSofA68565H6urGIvRkovkxJbNOwYqLVz6WEdbXsmXXj
RYuBsEL55+AffbDTzwrlfouyTV07sitciVXRYNZhFmpgrJGWJZA4IK/cLBA3A+QQ
7bN+sMAF4CBG9v9sY1S/ItHvfAIwroC2NZIFsAl0SM3KEDKAp/pJ7Jq2l2i941S3
mya8LnU3tzlcquFMy5mVWHt+41n+gt2AvOWnK+kPiEAQgLH+6felu7SNa+R7h7ls
1/kcFEmv0GSVY44PdBW9osvAcwkX2rdzz2jiGd+vGKOjdC5Xzh6piiug3FseVSnO
UsanbTMdFd4W3UmmVOvuh+QQI7+CJe1TfSZzeu69bTO0QAYZZf0jYbOJmOxYOvi2
E5H7FTV/LRrxatjEv5jGtdqHHhi1DqK1JdLsfWi9xcC4JnLV0Q/Wb152vOZbbWom
PVRSwcbcBpNXEnUwrhdFwqhJqfZaZ+ttejWEM1FZKe0+IHy1lf4lTyV1aKVapmYG
36tPd25Djaw6V79osy+RbfQy8BLCFJ0+Aa04E/Dx2TyEcySbBGYeK1ob31htX8Y/
P3/abNxTScwLrJuyZ1FZs9jctina96mQXGgXiuuIFN3E0QKDl/G08oEFOreGVbMp
LQI1H45s0oiJzj7BPX76SpxJU06ilTOFBalssu0lVX0p6es7l+wShHa4bmvuqlTH
+s91nU3xT0OZ90bn8gJcVX5zIvbd9tZhCYIx2appoqPmqntUHa6tlJEr+M4rvjK8
OeysWB0UqBllcYYYTcPYHd/Sa68vyG5uN86N8dsuWKkDXRGQ0xYEkTWDWtoFGvTB
0JBeGahVnTjpkuCOYwfday/M9lkIWdqb0NyZ1EYjYdhcNVyk4eb/z86oGReKfmTz
9MMM9Prvop0jt81PzQdvV0sL4RIDYh1RLgbLK7pidKzf8KZGLfrdHElLKNdVQ5cV
XqgWk6H4QbneDoTsWPmL75aaYi92ySfgluUnyx/BtZTODxs6HU/pnxYN7DKAxJsO
CyctgLD1KIi3A6xPgej/6afZVMHg0nORJpkSFizek/NOUda/KomRbAxjLa8deuSY
BedXOvSzasekD/4k6QMrq+TNQESHXbmF89HGsyz12gLSxKklvLoQ2+mfy3qrlamc
TLiFVPtWsjNP9y1s0kORMINUTm5DRs5VeOFsE2REe7/tBwzKv9nHZl3/wgIq5ue7
tggHTt46E9CDeRbmI21cUFBA5g/d3+iLADU5XJNksOdHlVCXbigc12TIFjCw2u2V
wOfg9UaEa4uEFOMQUhZggmJnrWJ3NBlCQODll5f1ocE2NpzgXJf8iMtQ3WayIFPz
PhaBCIQu88BdohBi6G+m+dyKrmsSbwI6/g44bepqErShZMPw60SvEiTMNxbhlD9n
RVFDtt5CzrNd2tTG6iV1u8JFhOrwEK7KhKwqIzlrpuADlBkQRL7x9+E2TcPvdKFH
lFFzOTadEb9ToPrFySdrK3Hb6dTsxBkiYdzGGg1rW5gGhWjyCkhwJBUt5ETXTpQW
VfZmWomxrjBPSPr6vH8CnMOuB/yQA9nroL+NdXQIHYLbEi1/P9syJAc94Auxt7eb
wdCP/3VRKyv2WPHzQfT6BBSlDLIUWs89Vq500FgKPBQJXotHJZj94Gzb8G51alHE
4mVfs2Q1CN6blpJr43NFH5ahBJ8qWYP+ssUK3hcVXempKXo0sbVOxeNNH63tLgy/
v2VetX9uRVwyZseDDYQU9c2k9qr3gKC8tGi01oqXCX0vI+ZaRZeM430jS0juyh96
r/QVrxGPJmn+PDVzCBd91/H3zvKOP1ZTeXLFBFg8PCThVSyOFLR5lfIAGJ3cnU9U
ibKcVn/B/fv+Y4VSnHQN1CF82ok9YCA8OcUDxlrSahSIgpy6l73mcuVx0MD2NJxq
Pxkl4Tvjoyt96fgtJh4FwKnDyrLGNbR4zBDTEeW3pB7XpvjR2XBtjAWk256j10ir
zm5fr/GBxaVgXYJ/GpQAc8MJVUWHMIu8wY/GluSZc3psS4FL0HgZefU1OCNeXVHj
2k6eEkU1SYHP0p+jKcuBiC5RsMBC2bhU21kct9q9VB/Zr5hjJHTm51B0HMyOy3H/
Xr2N/UJ+7Og5pnlnhtLVlrj/Ln2cpJTNuPqkTLSoTgzEys2UbMWzxUhbMpWg/BNg
nKDrAHahmqcguWPTmO7IfnvMM/DD1D7SZWm7CCg6a1vnXq3NQXxUGuockX20+yxI
O5Aeb3YGqNS+XAmuJshKJP1m5BvnJ6rNfE3V4WrhoZZS0irzLig0oN+eWml59Dzz
7lwJsr9hmjoRR+8WxU72R/1Nsn5yPqEqkk8llWyRggI2vduSPb++B7TW2/gYcn/Z
qQR+sgd9VMjaRec2migyEQVPqTsPJo3c3+v2hTR2l/jBP4JXeCLS7hkSIuHlSK7F
ny/wnlD/kIvRfyhHjTFXXvjN/7lBPrq9cjFt+8R/y9tgeq/PitUznrPJ71F/iDXD
y0HzbXtxrzFjui8TdTWruo4NGw6LQUO7i+3ljMHAwaynLYjLvWvyOvnfdIiwXklf
rTBaDqDYGDOxTu7wHcdxqZpF7yLK0+z7G05xVfl0WDOeyIqNm+IFKGMdhVyUDDzP
Nv4VHvDCb/TzAdnjFFr4s9GZz+PGGaql1FyBjKbnGjcNRfuDOfcQ7UT9trQGfGUz
oafTJemRujnIYteckoUqtk4s1K2pq7UGKGXSV2lyIbwIYduL2gjnTXKmTw1muRsY
UjS/1+4PpQiFpOptgY3dsi9bjh5D4lKUE9ArFzMicvzznCRqXPJMz5Lu+B52hZQA
eRZ8cZowV5g7hDmxBxC+Xcao508Dg76dSrKPhU3AYeTCGgFF0IDsCXZMU/X73U4x
/cHoGOV1sHPQRCL3WT99EC5OErfZTXV9HrqmyUPU0uHGjEE48vm5SwKqkKGZMIM1
jPbfTBg6CksLuKB0kBqZpHXqaGF/mOMw6tVBLtxVW20+HlhoJ4iQktBJ5nie6bk7
0xEakcApoIv7wY2KbQIXb7jbJpJg1g8B3gYO890yJ4GZYqGCSWChb4JId6L2DB4M
ZcvyLhdXqV1B4uXVZYGUByX+hnMiuyahU3Ya8msQC8ZPRJMlM+lY7c7MNIxo9Cjm
GRLiCPmUfxEAlVxFpLF2+U3JiWUNGQf78Hv5/fl/o9b8Ax4pVqcvgNNIVi5cL3gd
N0qEGto7jnogQ8Crg4nRlslYcZ3m1xnQfZxXUFOi5FlOBApWUt/DWRvQrjs3wos4
vm/1OlhstuXYZFdvj4uMK4sc0JKsRav7A7LbuCqYe3y9I599qy3DzaiI837S3Tvm
8Nzgn6YpAFMh/XEM1BaMIdY2UvEFiKfftI0fow7yh8YgE8tIRHNNMHvA4opX7OuX
oVD3oA0B86zPRFePWPNvaMywdDfIemC6hfPTf3QFS6RtmQjfRwkx9nlw6TgZ0zR+
4q67oCt6eUsVTGdo7dhEeCxhHBR7o0Mi8YiC/IsPs8/7HWHABU9sX36vGhKAoqux
AxXlvdSHZPegbuNw9vDcczcCxTBXsMGHGWu5XYwdXS2LuqIyj88X88Ay9jrVZ8NU
LglcQJ5cU5m7+TTuCUtHZ0p8aby/UdiT4JKuRN4uupzH1WnjiT+iWnNQjuuXJdaO
iG8n2Bs8Yh6fk0Qd2nS/pc/GdDLpdtiINBIAJ9YUkqc1A/F5nDCjIBtcIA0e+M71
G+DKmdjhjAlBjp2byLxlwyg8K9MUpRpSqNwNGaLD9GMgBeVwEQ4xF3d44GiM5LGJ
c+Rxgd9dEkjhjNOdWbc/f/B59TUpuNqvGFHDmv8EeH3YzGwvS8x01CUlEfSJBMWQ
3QNWRX+Fz9a29YRLGaKIBQFdpF5sMBqDy6e5i2WVXZ3p5eGAUsm2ARqCy08VYmSb
p7OYpvJ1guyNKmBVlstZf+UmQNmgT07M+CoUaj//H6i6L/QDv3odG0dMp0ACIQbm
GeKm8m0yOAl8YXrV7Is8YY70LVvHlHrNkP1fVyphJ73TQZIfDdPcjd/QDNPVlu8+
mT+vDvBYo7AQIh9Zpi0X4V9Y4g7ziHs0ZXOJopq7u0e9muuyeNY8YdTx6mCL+C2f
baONfAdAXFkGgEZxv0uu+X4caYgzJjEjf1euPJ8fDK8V92Zt/REvSAb+I5i+tXtE
CqoRExRkld8tyoFn+6WAo8NTJDCTwHB4OuFhv6Kb6WhBKkvMJ17igm2E+yCfl5q0
fsLuPysjly0zkgkrC9TU/kT+3npJkxRN/dVCoKJ8R/b0CnDtK/F1aGg8WeoizyRX
OV5IRmL9TUau62CTQnjTCE6vP7hwOfLWxq7+txJowTdvEFmC85Bk9/wuDII8JYqv
XpEyXZD2r+3zSvfPOi6dvS714GTuXxQ4QGqANcUhKRBk2SX+B0C1pfp8lH5EvLqz
Gh3zHt7pOtqbPqne7Z0b1Hmx40+Y/n2y4crGM/ovvNrt6eaJPR7Ebp17bTA2S7WT
tlSW4ODEnkM/ISf7SoOSBCoXQJZ+iqK7uOeDOzfFzJRa6WaGuPAH2wdHbDaG178P
ZLCnw27AnnFVrH2VRFYpBALYW54eUYeqrmlzccvBEzHp19YkP6ASRGe9cpfnbcMp
TjawGJeMsMoxMTrmYLbssfLESUEW+tS6YK+sWVCVc+Hp9Qdu9rMdqD7+wETVfRT2
Rd5SmTgcwNRxdfrSSZYdI5g23nMvp7z54gNv9ewwWrofir6g0jCJqBiloELo/rNn
+5ofK6cIMi3rn6Nrrhneq2YXslLn3eSMAqwXNBqWqrv2/0UNI4ESb1GFe4t89mdg
vOpQhgDrKiRrAOFXethtqCfNv6Ru/ud5XTcbBZIZLuGNzbqch9vR3Wh+U5ilAOQe
cQa3W1qwCf5iDn0vA81kve74xSR7kJN/1UbxeAobp9nxCNCe2NX+twXiAgqHIKIE
b7q2VYa/oEAHsi6PMzmNtMovUVNeLTCp5drM6jp+5Z/XAZyWI/XEageWGHmA63Aa
r+qd5Kmvojng5JZPUBI8ozdmAj3VWJtOixZojQCLtoYqwhRmKLNfNKhZtb2xnNq8
kVrRhqLOQvizeEIrt/j/uQZQiJ4z1em0Nm/vUxn9g1oyMuxlmbMS9cYrcRk18c6w
SFjLRBT6/BcDJ1NJnWUnZgjcvY92oOve18Ke3xmF8oDih7/Q9K/GahoxqQJFpSOd
5OCppzSXmPeYTQQWnVeC5wpLcUKtVqEXSYGs2mYjx4wiIAC4Xu0FkenSn1NeLfVi
t3g7mfovhweMKaUm5f9N1qNwneUdNbhFkMYHfJYEbr77mkbNVRtD4VZR4lfVKSPy
sbnrfky1a9dIyEEN4WM/45PrbogLpbXrLdZiWAvJ6BIr4KK1xHq1zggOBbanExcr
4NwdpjyRaUqkKsJ7O/72XQ3Y0DCQc4VMgtz3/3BMzh2lvEdaS0y8UDp9/a3EJ3sA
UyUhZ5Mw73EWfnzTheGTvBbhc2fPPxCJk+BGoL32DVs6289PdnAI4HbgsgTT3Yye
GG7pX2c83UrKQSBCKGLjUignAXETDE0L6eZOZeT2N00l8yqpAMsdMRuIWeVjfyvX
tZVLUBTaud/VxvCzU6FKy+nDTWztEDrqDMLjOtU/d+MP/lmr2KsapfrxDDioXcYS
8Z1kN/KtWe+LQ9Y2aULzJmdfSl+/wGiTELx6uHUO/6fRa0ATRro5PUBHXSZxU5jz
cSMci/sd7jlap8fg5JtrKPsBsHwauju3P6ONepfxQUFkDptHCA6RZqiwyFWgwcvY
1xK3Ch0kiMDq6IRFam2cp+EGsSkv+Gheu684ewLPHmOGaIkRAyQT7kDSWkjkBw5n
Geog6rOkuTl5LK+5dxTy6QU0eiVa8Z31mt6RyehGbPuWMKzV5e928OrjFddokoRF
Fonoqk5HYri2KZwaqd4MBmFEVJugDwPfOwmHATfvzEnHbXzV6RkyxVuzWlDBsBLP
x4SvoKrXXrg0Nyzhjs48+jZefUVZp/ZX9mO7ibkMDiWxlB7pB0EZ6jFSoNRqIROX
kWB2uTlicxEYGF5KkH1Vfup+Fh3Y3otY9okBcl6n+dIM0Fu3ywdEZGFcwh8RXcM3
ULjjZ0DW9RgaTz3dKG140lFpzUPSCVNN82x+q8zFOYfLwCBQhyvmn1DMP83WdIz5
ofkf9cQbHu0MDUF088MjzSC7lBx/rLwFrqIEL4QDIKohLmivQZj5XlDI/NrAXLeq
KfTHmp4nry387jPkYsM/kZqnpZpjwfTVCFvU6QMVSilVtQ9PNUHEFEoVywlW140D
oufvop/jeof4c1Qxdsax1QW8DOTcnNhDNviXA68/bZckCOObxoxVArGOc6RfLQ45
xW9LS2uNdLrIKdOyTuqnKfJXgJv399CeEFYvMQ6QipXz8lOEbY3Gpr65YQaylTgy
e/bh4pZVPhUfMOngHk00n16fPFDKXCzH5ABJwQy/zBgJQeqycdw83C2lEs+Wd/Jd
yQWJLIXG0jbdtLY9KM1P9FnI2mG/IEvWtEE3RY4AaENLYzZzDCnfDVDXoXoO4Rpj
UrU1mSVmS9bFEjE4qQsSiwLy16QP+gUFOyZIOgPzhl/WdtRQTP094XNVQCsXVBeH
x2aKxYrRinmEa4p8WFXlSgrRTh+29AvbJNkDaoD2HUxgya9WREK41G+0WnSK72j9
t6oQOqIVLgyJrRpsn1hM++1vp8JCAJII72l4RL8cnXrWc3myjrqMg1M4ZArE/jUC
xs0srGY2dZkpQN29oceZFpY5vGSyCM+bpYCc0lbQlwSvstiuYWCXNyiJiuyu5v/S
piySrQp2SN12smmuaS2+yyzDupW3+Mrf55oYrcov2IdY0K6ttQJjj2r6Wmk3EHgv
+LduzDsYCmJBUUWpjovOFDq+eKDwsaxV491sKPUujHc2D8JfCNb9lM6q6z63sZxp
C2ntynl5lckpp5Bjomp+mm5qOGKuQPdFjyECIj94ycirIUmnr/q5D7rIDmcxZJCe
aYS+2N3vztNJ6y92aJoIzJn4mSCmAWlrcC2js2FM6OQIME8Qm1XnZD8FGrZBQAN8
bNej1b0C3bNpaT/BVuIezGwa9DJG/pn6cjknkkKez74rPgkFqJ2tpVa9AY1fkiVM
Zd+O5FUXQNuZO9WLrIeH24fWsddxk1lNPnA9rsP4lOwEXvvlZj+tQM9CGPYP9Xyv
uC4SCB55XA2TW+F2vMF5VKSWL9bRp2XA3DXhP5l2oMG3IjDzYZXzlHNmtRB4vSkS
Rh5qGL6HJQXXcNXekX8R6CA+CuUsH0huFE0Mtx//ReJ16GU3elCqcS+ErEhZpy4M
v2C3NS0VLTV7B8oXx1ujG4e4je0GCTF2ASF1uzVqeg72daKiuGKT3MA51G50sgtP
S6zcSSkY1xSgmlyZfO3Hj2tXyEUy7Wvt3D+QrdDDP6tLbQ/m20DahqDef287St+M
+VVRDEH/OqJZLrFNbEmKEiv9CbFi2Qh4veRhq/Jaj+ur4LbBNmOwMoQbMgbXyzov
6vugEHJptDayedzdJDRC0cqKS2PtcZmLXNl3OxUAsheKtDi4wnCE2W8LcY4MJ2Ro
O44EDvJ+Bs1cAvxAnpgrDPUjrVCVyaV/wtNp1t/va0g81JL6C4MhRh7MD9ZEi9ls
1j1rxIP35X4Ln3IZZNGLs163R123dBJKc8zfeZ41TgLtvT6//QKkHS2S+fyZWZOk
xKIYTrF30CA+C96kXZl9bPo4+q0RAVDSWcPDhz0Lv1jjVvfFvOAuHD9eohPi7Ong
WPnhIiyFlYezo29LA3Oqw/6XiHjoG6ZcN86JyqexGTvwZwtNT0aXkzsk4eSwt/dS
G5YPAykQi+HNKpaat0iNwwbngh8gljQUsYlJlDcK3Hg7agaQzMw72DyqICQvr5d+
bRpQs+WeqU2jHnu5Aj54lZWNRCvZGKi2jTL2V2vc0Q0c0bMB4W/dgkr5IBp0aAIk
2D3MzA72w51xBYL0Jakm+IrOktA30L7KOz47hpDvH1QzyD+Ol01j8YFDlK5skCzw
anz5UTPziwwTr6jUyq93+klFQOMkzHqtqmgxv6y4RWo/ZJMxujh6/abaJkAHeBpG
AdVDbMcXUwOfoT4RtNeBQnR4N2+r7yXw8BoB0dYuyZfGUTEhXZ1dpF5iSnTs3ObK
QwZszXM+I6XKfsdrmWKn8x/7+gtR/9WXSttoDc8CBhnCtbOBmMi6MURrK4y2fTTv
V5w26AphMDMgHWT3twWMVJkO7/X1OZ2X1H7mtZBLru/XdbkN/Hx/Deq8zknPwcvf
EZyWsjdfbCWrTXJrpCyAeOiNp+AQF+HLMmyEOL23nHcpeVly0MA04mQ2fzD1EK2e
is16Pc2L9TC8fJpYPIXfjHsWIVmqbpOLEiFVN3isiH6/R7uA2kpuNB3pnqeIslys
R8BReBYx/s8vtb0heIgvkMRpEP0Bf+XO9AeeNI2Sy2vNc1oFtl4k3i4RBIRJLdbD
/mIpDRa/VZvBmEmfXooD6nJbxE1GkKloXRP25LVYfFWcaRtGDkHepf0zuj/eswTp
eGEASLyS+U9AxklGXzBvyvLQDS5NLpfHNyBuHwx2gy6VC0V3heDix3u6CvK/Ln8K
9uU9aPJ1CuNAiqbGJ64an6BYTAkOFt7etYylIF0Y/5VuZNCufliDEZQYUHUD/HTN
BvI6uVrt+dvWZr/I0P6FtdYKMvvG5HC/g9ii8oSSTiZuj6E6x/sKkHWER7rlJ0aO
GjUazhzbpSJOQgkVyfI2ssCgjR8quqi83Bu9ObXWS6lxsrcJMvQoeIi+ya9GZ6+j
yig1P5Nxa+XVigEDRg0018dZ6oYjUoFXlV3PSCqawzNEkt81xHAeH47r3tdkjEvW
rRmkXPIo+4RntcM0RmVsF/va9f1WBtXV7WnoRnufdnjrpMNd3D9YfnqJpsryBJur
uOtTimA5LyQaSxkxL1itYMjBVNYeofhrKEQx56JsZ/15jCYfRe7o7l9axIutD/lU
DirAt3sHEDWrj395HskdfM5bJMqOtXGb9vRe+U+V+B/ZD227c0pg3YUCItAHv3iw
8jm5u087KuDncTlS7/HkWIH4sOTho13NkJNRgP9xqocjAZ+46wfDVsHCHTodLiFj
nM0V4FU3o98schK46ACzL3mRHBV8HKCFRe7aEjnizT8/YVgvRySkndkkRxyIJAgA
nHi+TCS8rJinHnbAqY7Y8Utl7Mi+w4xRwyuxnRo8+jHdRT+sLyzKgAKQznF1J/63
yD/hT7+qLoTO0dBJrAmqofhOPWBBbvVn+tiQeJPdLjmbmboG3lpLaijtLW1FurfG
2Z3aDPp7XWhiS6ntwmkeNXbRey+j8lDpBAscdAJUlAu10pr2PFZOpBAkVZT5FW0A
WP4a4/SgKQGo30/xxbgxbxcdfsVBanZw/AEaj/gHkK4ha6mFxfMX6dqUbFGtNL5S
FuJIsPjmHC6MPIzXyLF7fUm24zYHyvQcAjZ3Tu1VpRVUrbihk/uJ8KHnvX6vz1Nq
QlSo4Sp2E8VRFFeH0IrxByT8FWoC0zW5kQtpRS53AK2NOLSq+ZFMKZzcvaj2Ny1u
B7kYKXkCpmID5vQbIazL2lTRyzUGjvzh8iVOwLlH5mpCixTIGmxLyLPvaUOoY7/p
jIlruMVvlO9HcJzRORQl7+voyzogGam3edb5vXluzr4j0PQdEAO7Mks+CoWw+Wh+
yOSXxKmWCbRsLSjN/SkFD7aAfIPheqNEA8XiFc9hcD9QBtcOBb0FVYBxjAdwMGOh
aQNR4SsLi06NHwo6kgUqiaU2ScI4ipRXRMosqXnRju44/IJ+BsgDtRkCG5KVjb8D
t2lOsau0AHDlZ67Cpw2nzyFCwct95zlm9AOsFH3Q6yfFYJG+a1gSOugCqZLb4vyy
5ZlNojlpUk4cTl7Z0uBrcyHmWMEWPYvhL9JeNNn2igbZbVUxE3RXIzFmUXFrHB4K
YOsD+9Aji0+lE3jGtvs4xsgy2EcEMBr2YHx2O0byndRhi5BBsGU+5kM6L7kAZxq6
iXvyO4nIth6ShpFZfi2qWglR1Z6+uXhmUg3oJmt5ebs0VM4waxasig/4U7ZMAbMP
/aNrpdAl4u4BNXBoFrC0WD3v4lz7glfisA6opQ8VpI3g3wnHi7yZ75LBHBCUafFI
gO5ENyYYHNlJRZCqynYwhmtr/TONhrxU/BZYqh/FBJPH7eLfNi7HVA3fFD8qDWfN
VAUcq2fhAkrptbxWeIWKKiFXcmqHlrqL9P4XSu1RIpyZ5jUxD1KXp4/Ke1W0un8W
O7YemTCQs8FwBNT50+K805MlEQ7gEqLYoaaLmKnHg7W4ySHklxSGUrp853Rpk0x9
ygri1u6kY+RzQbVu8Ybj6pfsJn4oZRKtIpN6CN96gwmGCDBojLwxYh5/49J4FPOY
ShJnSqhjtCZ0rpGuBrUREqyzLQXic4KQygtVx73iosgYE0tpR/j95feO9t65rw2s
brcZ7kTIaxbQGuo39bXZEbIq6T54xPZMpUPpd9uuJEdwrHmuFrz/7NEJR+s1kZ6T
5unOPfwbcs3a0gHWS4NG03ftYOL0/lzJM/I9Saik745YdmOyN081ti5a0p5shMgF
xzaf78euQzHXJp7gQ7vul2wG5kVNHFpUPoJKhtGsB/umnmuUWFTah5O9AsV+yQPd
1z7OpasvBoydRSVshgGtXDFBymis5yY7SZo2JQvDOepHuk7duSW7HtzsFRtW5gnv
oaNvH62dw+7jF08T2ZS7RSgvqZk/7rM2Q/els3rlCXZ62pl7/ELh7UjEaTLtF0Jl
Z37G4kBKxQlOBzDSbNtlFGvguIv7gj+zzUowwjI2W38eIDKcc15I00++hdI4WC/1
cs16HkJPiQHIZITp7gmxJvwoKayX05veVC5dEHxQMEXtJueAzwF8+e6PDC+l8WuI
qtfNi0nNboqI22A4CSRrCWXTaBQB5vletS6VJ82X3KA6OMc32nRQOJxCnTwBSiSz
P3vx0TmovhyTgvyIEATJHgzjBhVeYBCGKDo9Z58WsQSV0CyyLDzE1+Nn8IkavcfB
CO27ospcPxOzRUyjKGxkD6IdMbClhv+sTcxcZ4PGfIF0VHGSUYCEWksssYKo5vXj
tHdUmriCcfuX1dYuTMzx0dS84czGn0FR5eRiLfFjnA89oTZGNACs0p2LAAPekNMS
cYcy5zzRdMzjlQwWMndmM0Cnu4aCZaEFu89kyvtGbGWfHnHKe21DgBOLITU8wBLV
ZsnGFHddMRGkcR/UbH1ALDZwZlCPnLBRj9mqVV7zw2CXDUQTR2vLUSn26do3gdtR
qV3uWi5emGixFVF+HBG8/ZoLdT7dKz9v6XQjbymY4AirdRyAIV6EFX3e5e24qYVB
C5Q3fgrw5zGad0ZbMhnXknoy68LVBgUYgELG6QIHq96Xi6xobKtgEbVIUWsMk/8M
6QQrS2S+nltKxTmW9fXlDmVnHs0X9QEIJz8gsHmFo03x1DvD8EBftQNpllXR+A9u
9Mzlx3WVWgIrflU4myKPN4hdv6C7CgZzm1c04K7S/l//mzSaYtVf0pqeUrtZ64RL
fBEOQ+xe32H1MHHUfPM7XNg7fGEEa6yGYuBiZVBdIVRpCcelFbRbuU/oLuzDTkEE
8O51mKu5m4aU5f4Vj8RacfIcoBImwwbSMtSFZiOwkbv0sy/9XevfYP7MiiBEdO8X
efTniuqWYzj1Z3l/WHt1UWDrn4RWrl2YZ8JrZrsSp8bUZqaPq8SatkyUF/GFnHxz
f1Y4gwQoxfojDF3/KWbLu0Rv7d95XEEMo4uB2uJxpes9oYN4E7c6b6qUyuEVZSxp
itHZiYVyCM661MvH9DX4sKCoNiJ3wLGnLuCopq/YRRh+ddCAtwbpC1IgN+TFrslh
VwZw53Vdq9Wt8rZJYm+1d3+cgjodRVEyWP+cXbZUHzHlfnkfZi9ZDDLNGiavYYqO
6ubQrNggM2asA5cdXaJkjQbxr8kcvsY+ZT7fguP/VnkH53R54+kAS2UZ+4wRiaBH
93p2cnQLdUoahsm2m8ptLNnh4SJZUnwFyjEIeFEZulrc48diUO3DGiMMlYM7hcaJ
h6aHWrBX9xKreJIAHeWKz1edBNsOft+LyNOJA4YQl5haS2G78mXZEPVS3njedLRJ
Q4anYDm0QwOZ2tyRi1kXC4/uczNhVK3V10m2rj5W1ilBSptLhf4ca1J5yprBJ1T0
dGAlyrUy8kuWXX0Ivly1TV+jozbrCQn9WRr5EAHuuv2BskpkwqYDunbmGRMWbmGm
GfuwD2rN50awbP9daflvJsUxQoyGiKdXZhIYs30JDSBYFLQp0UwZ7rQBWYgvIjmR
pKdESpfe9C8XE/9jQisuJAZOQFF1VyvXVx4y+xu+/mxvMEL5mmzfIkT/r0XPrf95
N9PeBUb8vXDNXGE0w8cg11/7bf0yEZ3vvi6fmMSDflza1vCD91XviGvNcWjckgI8
EWwS9G+hAK6se4nVpZ2wyt320xEFLd6stHBqKCgjPelbD3TNE1ZI905yv49OL71D
hzIFHGSxW5RXo+NKdCXdKGu348JXwDx5UTkj/hpxBkindf2UodC67AmmAkLFmfdn
Bgfquu+DjTPLgfumKlKMbiRWX5sAtfyJbZhpqOSqIayNx+Gtq6SfsOnx6pWuXqc8
jTe6wR4yTTTfsavec5i7i/8AcSYE2kr6X7dwgEmafQUTx7Verp5zqwYvW6k4VH8N
/iqCnYu09HYVmDyQ5TJd7TO6ClJZmlDsDBQAK4fWb/dYyq0E56jVzphnjfXxFr4P
OXjBuYzFjpyoIAbsIrZbANiGFVantpnoKRyc+57LfCzn2bBZf/zhx7hZTUuJ9OSr
pQH6PMKIIhRoEj4CCe+Eveg/0zxTBjT63IeER9pKqSYG1chH5Sqd2SD+iDGnE3z6
/zztj638//eT99hR2iiSl+3CNxwvwA7Gg0qwrURTkfscZHFzbGSHWjeWAtx92P3R
SJIzod9oy7NNbCzecnioRTTE/73nqTAH+fweiUYziy+ALkZxCQ8JEiwzindAsfIf
ZMKaiuQF09Z5yo++DdtKbw4Fm24FV+mK1oG/0dajWS+Vsi5apCaIK1XsEQJY+Yqu
7ZaFppZ7a+F8ZGAPSbrN8PNhuJcDYExNY3M0QeVGRxJq+z8472+tDhKLvndcjio/
sa+BZ4bQqlAIP09ZrYHvcnXtuxCE4o6RX3cTLfP8bP4hmTDBwUc57UB2LDiVc8bV
E5ncfoxhsVt/PUEiFtADQbWLI58iOckFJPYCVN/8UXhzWR+n8ZnIVVabcqEdADWR
68EN+OvW9Y5NlaUWOPL0LN4+/bnS0filPGj2FHde3A6/ljRHuCGW3MdWXXy244Rt
F/3/KZpzhkg/HevlwZEvLyC89mEZCWpgsQx8sKwGFde6U0E7D25YgGK8C5nD7kP2
Px8Qdns9NF92G76SQ2LXpCsRUMFAnmIIN6SPZbpbut6a0M37nsRNGiQ6baapTVOI
2fhRRo+jbk7DYmc4l8mOL4scR6ew07T2Sp6GmdEZaRyjYmqfDlTPgWfeEqzAn670
H75TpjKKNn0lAVIBWdAF3nBTs7xaG41W/vRM6n+RzGCf23LWKGy6fmnt4zDTjcBx
vto2q8o1JTkaBViarRiKYZaeLp1ycveTIVe+UAc+FudibzxEQ6BWumPjWVYefium
ZxToO38Y8QNmKnsfqiDPwkLOhiuYk/G+ly2ZURVOkLuxAOrvMPWWUzRxSZaPiQzx
ip8qmFp9NdY+aburrZRKWULgnBqLt3FnNmdZwmzfY7sw/saDNxK3pbc2XS5mb+G4
9gE7LOZwXsG7tuKZ6VXbMEk7UNCbJRG0rmvT7TV2/kn3uujQKZ5T4KIe8zZGwvdL
jq0gu/rGpZuCRR6khITmatOp+p94P1F7S2IY6Fu754M990LusXFXjSu+vB7p0/Ne
0GhJAt0TJnAg73xgpP51L+i7xvGxyiGev9ZdEDKAxUPiTDWwrEHAa+2StMBI4D7r
/j/BK6P8+fz5zTXwGzobEFff9Yz9V8hSNMR+koKvPM5Ztya3ylpYhAx+u3vfRfva
FzFytoLxYUX11ElABWl+PgxG5exWz4+sdx0D/YFdTQGsFBkT9Ogm1+0d2c/aM922
e4Hy5G/ZCLLFKnojdGjkYaZwLjGcbdtEFxF0CbEj0SCP+ZRa7wJ19CwH1b1vXpMc
1vBhY4DK3WJ8KHNQM8PdqHc5qfFshVqTcB+Tl4xtT4+5xL90DWfeWJ7Ks5NWSKu0
wDP7vl5n+a3pyMDxsW4cfgQWdXfBit0nkQKWC3tIEu0KiBWTTMFP13MzcDo8uE0U
/ViL9ti5JhUgFopSpCi6P9AbEzQPoWvDaN7H6G9cBABcpXFaBIpfiThWhh5vpmR3
USlhLMnsc7piFi81/czMoQa8WGTDYVdl9GRqGIIGkFoiMVVm4eyLhI7d1MVrErkK
s7SV772HUdcW3+Ez4mGZd0NihuuL2l1GRCKzZ0PbscpCW58wIPOu+T4XCvXMRzaS
Ts+eQrhgRJSCZcqPeBYC2kQsXcbLDWIHpL95qMEH5BQKCpeUMAQKRo1xv12CgEVh
EnoYYwMjZJ38cn5mhK5MIvvx61Hr5hyRiXGSLUc5zOLVDL0wpYxO4H0VbZI7PI4H
Sv9+flKBgyYLMeCj4KlmArvuG7nWicv49oPB75SVUWxROYCTEcdx7+7fS4yaASGS
xIHQAnXbRMqSq9YecUtHYoYhbKo/jXikl9OB1ab1gX+cEV5wwp0FCEpW6XddeRRv
LGFithSzmofPST22u86Mja4mMUDAmTsohsdVG9f85ofgMrHTPM1prK70oTCaURV1
CJh77It73j1Qg+dMSU93gsbDyNbFsEA5TrMe9rQAE/mP551LlMgLum8wqihdSdSF
HskQnNEGuX4KtufD0Yu+8aZWaZgd4qDkX1wh/8lczZeMl7v6xOCzOeGrf4LWVjlM
UHHwkbw1K3DxSRmoJeqa9ZgU6sXV5q7WiQ//Sa/BLfy8aO60xRBV+ER7+FjBGzg6
kqAm9ad5wbI6trwIDrAcZMOCDrCB6n3XUurhxM5NbLRSdCw8ngEsqjWqZ1p/iyKu
GlRumbj4yl6ln15OGSe7MbB7uJIpEiu221ydkeSE7dYOndAKpG0fZdqnOmkO7DS/
UZaPczHSsh05UrMHSE+FPUGoZNmL7BI2DMfgG/3XL4H0A1xI5QgbMBltGpASSS1G
Jw/SDlsRtZfpFgLHGdWWXAoji577JlN9V0eEMUwP4EAJP+EjQKPgjaAXRLZ3tVNs
TQNxA8ql0nr7h8007DxyUB7x5HSysh6NRAWGUb2VUTaPporz57xaCJkapTBpauFP
zJqmb7uiN20lwriiGrpQVL9TPvUc+WnfDeZ3Z715ujIiSs79aXv9GcY4iUn0Onbm
ZP4DDiIyJDgbmJBAzqUBsLhnN+UYQO/9sAYtW/uexzQY0XGCU/BXBoINu4QF325Z
/UrreBDEREB81TKD+HKaD0NObW425hIt/ISWTM3zTzhC/OOtdPxt3wDNOBig+vkp
G0Lp2uzaSKs5u53XrWzdNS6p7hWHnEpcM9eyLpcwPe3Kpq+9RaMUw6Hf3Um5rCY3
N2P/fHXTKrh1+ud4AX6ErshBwtXsAobRRGSCpAiBL+it7wBY9tL2F/YOnd1HfTuI
8cDx/4npgRqUvQHsNtjHN3IywgJr4spF9bJ/kRn7NbwXP0xg6h3WAoh0tgM+V+46
EvPK4MecpthNqiZu1sGCcinbva6l4uobCip3LJzAaWnsi+kS40EJaH7oCeyDIQof
2JiO7JIQQSfl+v1B324m750HfcnW2UbkxUDS2MwCl0OjgPj3WwJEdJU6rrtUJFEg
8gaj8HF2ZGl/GZTNFH7lSUUtT5Hf3D3ZOf9z41BlVfxPSGsaczJZdxF9tj/8vja1
MWDFwyzp8N5tWwjJ8CyhDXB9ni+FIRphtfT8CmOaagnBarDT6Eh7M9L/Z81hjd22
SqLtHl0A/6HPZWiGc3giV2W+Phx9/JXRsBfo/MsEy9Zuco4srbsVskFfkoEKimXK
xY2olkhgWAIU9RDMlX+SHOcZgrP0YWNVKLYIc1PsxiUCb/LQXznSGgZEs8mHp6vg
fINHXgNSUZkl/Pjpafx06kpSF9RCxTPIlz1kBu0n4brpC6auJxyKw7EDSj4cGnqR
lX9JJmiU376r2NZVjGcuWFqsrPGu5t38nwA6wE32t7LuJ26ctUqAtxStt9g4S6Hi
nUWbpLaHjKP8DomqD3oyu+WxRm5OpZOuXKWEoaLbpDP7JLj0gBRWXsKWaATqasTI
OcQC8PUBxuVLxgSDCZjdwBSd+G6zmOhKJMkzMG1c0E7XoPInMODhkXHCtr80rjdN
8AvG+I3HJP6fWOEypgn+FfeWejBFR81GqIr2OH/yQJel/RyPJ3GMNgK+2VqWoq/V
lT2KfNkgsB6pTRuO4lFQp9ZzFeBhcqu36o+hpDqJUtcdTukQE+qCrOPxTXi2yUg+
1u4jVSEEFTh00MZt1s77husctFjs7Trir1qTkd3yr70cQ598X36yXTL17TG3WuvP
o9BHmXk386sNBwin1rqc9Mahgl6iW4FkV4GJzn61oHnCF9EPmWT0Yn+GRCQTI/6n
RBnknmucE7ElhZGX0ioIzVT9w1MarLq1vH7/PGM7IaRfjXB3Pr+yzpG3WCfIN9Zk
NJiJ/tAVmDu1y8Pf8Bjwe/HzEBHT25Ujrac/FjiGezi567MT1qKyQ8yxqL2YLBMV
AQhhLK/h+x28EkvKsa6wEYKbwu3Snyc1X1Gm9Gl8YTD8nmQB/VuJYO2DpOTN29h9
ct8k1B6Apalc7YQvb0reXjgPnLLBIYuATHaSY0BYVd8ta1B0uxC/PevOXkb+P5bq
lbh0STE8PKuU29Dj9Z40Ws7FmtNTDtH7zdTV3wTPtqbihp4MVJ9lYQcNpQxe1/i/
VuHEYPivTUQ4vWt1D33oJfm3gSCRgM9jhUOcF0KdHQKWmpflSCLj/29b8ktr05mu
9tDD/z2GO8SSobQwmuAqFhFUKiREH8gqxfUqictgfxRLL2yaExjD/xj2N+QM9Ibs
BL8YmaJOGgTCcE24ZgyEEDo/WMBbAw7cGZa3CfR9iUCg6wV3N9t1gT8KVLFaAe1M
t8HS69y5CKe57NOIz45sUZyOMiSrxZvw0b2KkGgpWnEtg+/2x5CIpZKy1gIjAQRn
5bZXUmVSIYrhgBeTy0L9Kcbq36wxZ4c5Ijh4ChBNOhH0Js/LOpBo/zRf5GjrYieL
pjpviqVSlXUHBBYrFsPz3ey8+spNoUbAoQgfR2ZppW7mpueDtZC41taiZSdi4rSC
OCiz2HK2gLUunHCBYl52CHtcDNWlOnaVbQNRhF4gUz30GNWO7A4eumFcaoCdr+cf
it0bRwYCHM9H1sXH1U9ApWBzFgVJbwAUUx88zhzOHWpZH+UspvrI5fCx7ZfHAEgW
nCc2xDDG9yDHZQjdF5qALpk0lygduPCKHVslBD4iE4D4aA2kQAGXeHmThbVKwItU
6u3ypJHjPiSH0TCxvQlEMiKc9XlbsMfzXdAhB3L+It7uv5sA7X2KWLv4I8nAV1/y
oLLqRL865tIDm+sOKaVVDUPr45jQhrV/YKF4QOkk8/bCJe2/nbtjn+LxRn62IgyU
UKoDrNhfIJRmYtq2YQw1F8yKGdH+Hg3r7RGvhiE0+z9w2HV79U+Nuve6VFq2KKm0
37RsP6lXswhgk/UHYTMKZ8fC5XdH8RJVDitf4lwXwabqtqmSHtwSsMsOwPwVZuIy
TA5s+akX1zXVVobtoqAgyEkbXZkIk0kTSVzuMDfsjmu3oJuMa3XGMcw4K9e/IAXK
BBfN/PwhX9ZRcunC41aBii0DZBRtuXvn49PJvTrgwgGrrfquK9ANU4zG0I8kLvjj
r+7VAZvCXxyELoPTxoMw3z7tUHlNV+NXWjBkf2y0RFFgGQajrzRn0XGmskI3OAnI
Dz4QbE0WXThbCKkGZ6YPl9DmHPh54PxuQ3uHkKlurCPeUFq5lFqHWw7VGGRQ+rYE
aT1VTJ2bZqfFXUUpvZHBhJNacw7Jo+hjZsj/44glsqz9SGXHXj37ieEOzzYH4Sx2
rEllqrxZwjd8HtqAFYXwqjYLJhDmz+FxrzbWM/8fe2IKMJkJf0SAXCVY0uPG3wov
1LP59jbKwJUmpnuViHXIPZ7ENyAJaXyI5iuCtYnMm7CIZvdAJ/+ujumHoNYCSBOn
eaDqf/Ix+81qKzZ9Zz+EtdFA+63xl7V97NnT0cnUAmujfIR98nN4nDoGVdP9u39p
/JPBgA82yti0aak0EiTn0UBYmYgb4zkk1Dm5qEeBKqSCLM8Hq3dItohluDJKLFDK
DxxmPs7jraoD04iruTc1rBbIhqNwkWvRnLjQhHeYG5SiqQ2URPwFhPzBhT8NaOXB
mr7tRISowZ79flphGSkyG3IFw+7DtsfnVni20ERU7UeyFh3D7/UGSh40aEJd23zP
Z67rg8v2RbIWDUROFc72e/e13tCgiWgOvKs7xdSnixo+5ZRe0RfbAjD9TLUoIcwX
XXE/9rgv1zfdNwZHhLga4YSP4crl3+ZF2ZEn3aTNV0EoyaMQ4yKgY3WqpEzPXE9L
f6DDlxNc0HZ40JAFY5PA6ausdiw5MunLbTiyLQayqHTo7x6urrCEGHpCUCCTXdvH
iF04So1lBvkZaF5jCpLeCrahwiZT25MZBY1RcW2QkYltI3BbEqz+pCbX3u7p8sqr
xzY+sgRQKqAznPQfbGO3OIp9RmA0FgMUsxHNrKw1zV37DxUdN2P2iH8UDtjOrOkh
1Mh/7lEd8/H/QT0KQBU176DRxJTEg6q8Qz/oRLyN8DDoM1Bcod3sX4UvK4A5dwLi
Ti2noDO05TCHhLrXYVvgNaZaVPhVqx9PZQYVSoPxUYOXkYMiZfM6A/kd46/Dqo86
wO0D0gqZ32g7+pvi9H6cgyXFMTgM+80iICLPd8URMoBMBwTriXYSsrw81CjQ3o2/
M7RiHdsRTibNODIli+R9i3Px1uh0nZTCNavzq9s1qlykIAFQFCT0QxSwgb9E7txk
wR/G2e+frpUHCXGucKGHXNLtNVpCJRilmvjCHQG1glVecdbpvsKDKRxkuMGIpg5J
KXPKRdv5reqrXBUjQqmFm0g1dq17VFSJFWJtOWd3n9A7dPoSc2Ph6sJhpQllpvLW
grvipqGF7zL1OhPkS/F4nKcqaKug4UwBOQaVL0OnltybpyVB+r7IAcirtQRefk7f
Yjy3kjtKZzBJPM8Bq2StEvppnaHPXOYGdTrQpnH7ISOEKUitWJ9safSXGfdL5uMi
ECrm2SQUs1X6f7yypaRZCDOHzYB7pxzZaOum/UOA1bApUfMS/UtLPQP0SIXl/HCq
Y5Z9AnTuhHKaG/iPddQ3bsjlVxevDkULnawvaDpjtuRcYOUenbRiWI+RxO3Hlgft
vku8e9NhDThMBeXRVXhwGw59T7sn80gZoC8AGj3/GpGQjLDLX1h4W+PrM69EArlo
igW8VbdhiNoc1NnLnOy5plKSnggrySUzq2WNb/lh/T/UcSNC/l3a89zhhiLccvoR
bKSjrM7yqnLENIusUoS7O/qeg0sTlE0gym2Xbjobhz5DHaFZRZxEB3OSTNAc7rub
SlHFhzch+Ih7ravUXlBCFW0/Mn0MrBU5YbDoIG4iqDgfEqHaCTKfxRasCP9CWN7y
ZSjXqnSo5/NEc2H+XCP2YvlYJQC3N9ZyxJJQdFEzkqlJOa8kemCF/20XEy93I/6h
lzzwWyNDCO7J53HiPHUFdL9NNWFBwCi26IfMc6jQQ460HnzldvUek28NnXhccO6i
67ZH9PiDRFUdtRy7hRQ0Jl4CEo06UGMK0/Vc/jWsTqp8eIjR02/zZXPabHYLhzWR
UjrjqrjiMH3/2xmivUihxtbGyjWzel60ICOID80KkBFfazyG8lrBLmhriQWoXfAU
qVWs7bQL9aQMbqOmPLFjQS/2j2hMuNsxyz5hBT+/N5zWDyhxTXdIzYF1nqu0+ZdF
LBnHexMpzS1wUVsj+E0PscJlss4XPS6Yn8wLagjsg7FPKZbxKf+scHakCHm/mQtk
c/xGglbZTaEvhvPAq+SCbh2AEGv3BmhGyi5q0n1dH/2vbaTD7MUqko4R7LcHa+4X
U5gt6CSptHOlPx7XkewpYLz5W7cHA5exZHlUFIbiU6wTZS7z0pGp1GA7B1mTcNt5
bVfUPddIyxi6JCZGqZZPiGi/12ZlPO/XuoRYJvSTZUCSiMwHupp0mFPn8QX3wvfe
b1lhPkxvi3bAENdGDiQs497MNFcgZl71TGEUjLE3pKpgCSZt0W+Mt4uTCzPWhEId
OnCV6QTBryxFsqQ4h9t9ixGM8IVjdSweH1uMZ3NYfMkqPfRuvDTTh51OykyKZJ8F
KuAXYd1H90xwkk8XPo0P9PQwaH/b6Uv+MihJ7gugMB1S+COkaz4iPLNsJDEFCNoW
SvdzD7lU2e+AZ8cYNHtpJ/f2pHWELSXIXBaiD9lir+lO6G9TOufdV3O5tzjhG/PH
WR9AzlK75c5b11iHp+VzPYQ+EnKHK+2C9Yed+vf67qZaDR1LcjZJLejEX+ely/vg
L1sqpdAHj68LrmsEhinqWpx+v4Fhs9ecAZrlWRF4CQ/GKHZuMXr2a0QzeQkE0crd
eiK3aiYelj+UgCr3QBDweOZ8xdbHFt6MwbJ3cxp/p/1tvONvLmV81XFtVVIxEvDe
QvINmgIXHmn1icCvj8STYWLr6Cg9uy/E3Dvtz/lcOI1f93TyQb6u/UwnzMOcH/oc
vr9ejgJcO4MJTalHFFBdVOWVO9oJB1BnlcTO0YocJm471aIDSgrrylmw5Fx052WT
FMiRPtwsJR+Zb+1qKGaQqeXD4F71gl8QV0DEoDomP+Z6S9DXwGGa/gXuqx3uwbyo
mjlwoU2NeErRcSVKtHX9DpMlj9/IKTpdmNVUxJa/I6Zfvd3kSokfWvpgdOOxQuR1
5qB9CEARGAOrAjgoXQa6wdm11qn42oSk/VUtGwz0hsKiwsAbKg7GjbIYVPeSp34j
AC2OIfGrCyYqbIPNRH9WifV9qDKXyOj3sULF7PzWVN3hq/HFLNxbWJtmwGc29X6c
z5gfMNHnoap6k5d4TCnOuRWSxJpE1G0WztT8ZhPMeGNW8CA1cLnObnsBFBFltkOP
E8/JlJFGxuK6ZiH43GjAN8XFbJCXW/QbOPWKwbTn0Ur9MQ6JlEgdM7fjGECvfPD7
/KginA5Kij+3vr3Z9EDC7p8WLsrn51Ke4YHbfIrIKRXOonloUeGhs2JLLb98cogB
SM8MH6V2C47mXL58TXnRTsNUlHWdb/u1HzaDQrwc1ej7Xv8xiM6RjRNthZf/hUBp
eGL+GG4KK7A9XlMYQbq1+fs9NSd6VGw5deBPnrvfLSckJNWCgcp7IkQi8jvwLNK/
yT6ygxy1EF6gpMsdHVDuHrCgQlrERmOMfWkqQET+RNGfvCZ8i473PMKsyOe2cFTi
2q/MUUr6fyseRS7B4wnGmTmlGHaNJtsSQIsgpc8my95VNZCuu8UnenRzaJ50ZYth
iXbWAiRfVcM+3fSYeDi0nWjRVM3yqw1AuJgWGN70ke5YyRroR/p+9BiWnTm0r12E
WTJuif7Zk3Bo06bWb1xgn+uinGMQ2+Zux2U8vVEOpyiX/00GgJKJHz8symgYZMvH
lOJpjyN38C+VGxyPq5cIzwQdaR9UIwrl65U45+WKv6lqFgoWvuRPHiIlGJZD/4Eg
xlim7ciP9lJrFep8MAGqKrspipYFWUCTVoALfsF2s44mJy5YdH4qKj38m6afecni
uiBesbEo1X7fNlKAlV0MoNZTTNgkmQ8PqFkhLIOKB556RUhFv//5t5XxfZelL6u+
V7lVzHgSlgvq563bF58KdJPP7BqbnrHs5/ajw+fs/kIskeaIkJvXrSuc9xkPvcHA
m02orWjL6YHN0qM2o0rjdELnI7BJSLYvNiBPPdhfv4wjMW01QPgqA09xz6nt9Cug
AcDqYEI/uBR9s0LJqBKahWOPb13DdjcPfy2gn+2XRkKOhHv84O4Mwi4unc1MK9Qs
VNTE271oVoaPnosSk0Wceuhq9QBpLFsHovyPZwsZJMnH9A9dy1z+XtckEvJVIyLI
wkDlLDkWIzLzTJdzgbWgIysVfTDB8ZisW66fwEwJJvZmdr5xXuzxaAAYX7bSwuwj
TQ4ZtvZdmrQ9lzaezgeVypoIhbDlmN05qwClRsqSIXVbEXgfOAlXdT7g6IXO4Til
rqUyj6UsShucmsoNckPfpiVGwAO6LCHjrRWW1SiVI4MDaNKhujYJcCOGv58ZkbC2
YB8tuPjhTbn+1YCQL0YodQ55YXfawQwYpSx9brXD0hl3rEmeQ2meOcsvs69DodAZ
PPMWFcpKTBkTld3lNOnbtlLASQknBYkuFxrErM62l/9C2MWhyFKOzP/mqF5u+NI9
zdwUwcrylSbEWg5t3glWuehv0ltTDylRRGiQSl4cTUkW95r7uGzL+rUUsk0+X3tl
d8L37ETiy3RL7GzeiLdz7eAPVRt9g3Z+K8Cntc0IiobVAVWZISlNEAYSYLneXpnm
ZmuXF7p1pDYEcPFP0K4V2kOj4nVlbo0d6oxYQYZMpxTUL14uaDWmhw4Sydd1xJUU
jRXQajAGaTXByeYGAml157sIMLD6Icw33forvGSZ+TFfGyuee+ldB0vPN/2rX0w9
zyf24Rq3mVlgos+xHT6ZBPPaCyhv9E3Rmv+YDnHDy+Fi4GxVOIEh5QDSWNjq3RX9
yfyIQ9Lp1ndd31ChspC1nXoRmSeYB38GmS1VrjF32r12t7f54Hg+kfq4MADu8/IU
TyDc71/Kudg5jAtFJBAKBvrcmcK1f8qGxERZ02ylqHerKrpnAGe2D3dXurSPrCQv
WAKMlIrUhaWChMESKgzcQVW5YW91jyfZKa59krS3Bh9PaB6mvhg3WJULZpu6n7tY
mzREFZApGqfUdju3a4hTEFHVrcRu+oEDxwHCjGTvOOvO1sMgzmrLSjedTLf9/VdB
kA02pR6h5DKxzYg+roP1T8NcU4oE99kxF4lkbdrjIyLcVuL85LTnTsNMnEpjfMIt
roQGE0sc0AAr5hqfePYmGLH2u27wcxomOEWyRDqF+9UIxc1X5Nj/HZclCYfWlWi1
QgTVJOVJNuDLIC6TcjLbGyVra7RHDVzXTEtBJ2v41foGOz/dJyl8JhEvLb8LULUh
Arf2V8iGWuDbPh9CmjCCXAF39AGg/arLhfVrG+iuse5WijjvuwzYC0wAnw2A51/c
KSIFIpA8HYca0P1juZlJZAd0lVpA9R5q1meqYqrRxaL9S2T8Hg6xhjxfbiyXutOy
e0WS6GWP/PXtrSPTvoy4KroTzXjcKnWzHYBW4HwpEYe4TzCppz+8mHIzoP4OuZa5
D9MZ5bSlsa6OAj+T8kdzP+M0VkXBGue6IAvm1oRvz3QUsRvJsZPigCrrV/IINI9t
aiinMlFp+mgyl6i5L4dYjrRNQ/vgS9d2QGWVpq+XYfjWiGfDbm0gkMb+JDRRHiE/
NBOU9h7L/6How1+bEt54lDB1w8A9LW2B8LhSP74QCsysbG80yC9q54KJZvKIVn/X
r8gNUMMq1+OcOOKR4IQYB40iiaVAyk/lXuP5+ASQCvg5YkRURtls28PiIGnWU3Sf
rauUEF/4/DE54mKT6wy4l17jgXDzxH20ha/CiOB6kmrXJ1gfecouYPD7anTjtl2L
Z5A9WB9gkEp1L1AsUUySym0vNVqKXbiS/LOVVTNKOz/L9qhhRUyf55v4hPfH+ztL
D2gnANYXBdQ4GrYWkmA1kXmkOho9Q/e3i5g3Cm6pooKy9+9GnsqJgqU1Wzt6HWcK
DG5ezcaGpDgz7ePNhJ123O7SJYFIkZPD42OvXiREjeTV/wasZm5DYLs9MK/1Mfye
LCIzPqRV3BThx3t301InwE0HXyMH9RM9Kj9NsLRYJWQC9i4bZQXalgJumRJ4Y9qH
nCjjx7KBVLhfQ8F/O5HaDHS+l6AtLmDko0u9vv/IcxvCdptRqvDrkyK0aLPbBX19
qv0KK0J9UE+gKuqJrsaT5hwVBR+DZ9K8lrwaVU9196mNjZ5u4DIr8nPmr8FjeZVc
oPbc6sRaawvNfSF8+cnSsL1N0zk1fduC3BmpkQMi/LXLOuAeBqz8giM+HBth2r6N
x+IIxqjIsQM7ZdRNsU/tjzSxKZqA4xqneMJow5yqLzk0ecn1AfpVMIaXCQHe5TOC
K73eBjniw1IHZGXkfyJmvcunwImHv5tHX97sjeJprwYliA5fTOQmNpKQ74q4Ek+c
gaA0jc3kFfNNvx1YdJMlX1O0Qohu1Ng/8UOeYxKDoUP4zZMi9eC/TBckR45s1Rca
gZe216HYcpuHFdZxNtdTmmFJhBhPeCQAZOdayFCrVLfe459TX4vSf4LRm6rpIxEP
VOwfn7PYA5U3XZyDXhBX0h2GjHkpP6QAae4RQ2NpwhrDoYVF3oUmXJkOboraUPzy
s+V+uz2iM1NHxPNmFgT5euw92YW/3sYsg5hq4YZMsm323xeuR+hAnv+je1hUzuhN
KCtVCclq4DlOVbwnzDJSYOiIOaAwQtXFzER0vwYslEaQm+z3iHjOYFbftxjam+gl
H9fBpCJauLJSJfQDYSWjw+sAWlpP1FlJfEKCKqBjZpj4Ld2/crT7OQ79dK6B4pIf
b3oZOsMmf9MlxRCxO1WfQM8nvOFFn3BdMF/CLmbQH050enhdBxm5BwpbGwf7KxOG
D0rTNw6nh18csw2BMrTHv/8kCCJqLJWX3wyMoPhA702/Gu0TLHZj5Q5wvERlRaTR
HFY5tdS7dZDbXicoFMeeECyC1R0oEq16x4hUOt0wmeqevbGxAjieygICGWUdvQy4
ITf09YQVxZxDWZpqlHdEc1KhD/6kx1QInwi4Sn+A4w2jxYk7qxBvP3GhLCna6oyE
7n2jkFfgnda0+YTyoOoyJpRGMlxGpKtb8XT6akPb3bDgrrZfWat6Ib/EACydaJAO
SPa41MuGGznoCmgJTFuBT24BwEc4/uy6pCBVo3O+qL/iay8FfwijcTcbwogTy31+
apJQDqa11veUb1rH1pZyorsaZ3cxl6F78hiSpjKQj5hFki3ReUjUUxrv54FxBdcR
MvVgf53pA7HmWExJmS2zi2PLQGQlzX0pmCLnlSZboVPpyrvX+YrYgvMW7gYjVXVT
3w0WByiu8Pgv/7dWpNVHrmI5jxSpiwss/CY9CIvNAzFyEM3LAQu3KDwLqdRWmY9J
HhJ72cY63+UA+w0SicDOA142LAO/uBPZulwYHIvtqCr+wBy1FqgeA/0m5SPbSXUi
pLAEJi0LbzWe4+8TjLSAtfB+0MjXMBVKXlTtOFYPPdseFGnZLmuuHMKkHiD/BoV1
ud1GoxV5Q7fwlPqq2GdvYAqXoKJ3nTFbT2c3g8KLN+LaVoqqimH/sfWuU4IraLc4
238q8+y+LxKAfP+2fS/LJYDqk1pbh2ewZxc8o14e7tVjz9Udgb5ARlusiTU0hrkR
mw8/brLuxtfMvyckmF4Auyku5EN09H6Tne4NPL0z5A/MM8/KZ8TRcVO1OVvBwlnC
2Mk9/UDwr0RWqydL7evGEQk5JNeFG8NDFGGH8IoCYd2y5zDGGdf/hYt+kFdye/9n
6sv/FStNtnjvYqNCfQ8huu7HUfTBHuChk0C/kSMJ3dbsprg7tpgwqdykyQubjqYj
FbdY6wesLxG5vYsEZGxKXortmycY/gZGTKgVMt5QwqOm8iFxDmQ39c34aoFEf2EQ
l+go3brZK7bETfpwL0rpQOb2vEkjc0Mksq1uDgcRc1uirLsugb/qSjZfliwiNMCh
zgyEIoGf+B6PWEml69GXL2jGnP+LG+5uftKpM0ZcuYk8FlKJ/SaBI7k8lstEi/rs
tIJ2gR3zgtGO9uF3k6FtHH8bMBl26DK0sOB5QNO9NXZX5b6IE0eXoEpweBcBX7ba
KknhfOG+eH1+oPSNOPb9n0zSt62OFrv1/awe8zUEXHSP39J+aKc6HCTIqgJ6hO8t
JDHF727A/DdVqpZo3K7jFhY3nnopDinrA6nxkh7b8+pIIZbs8ZGrqZfgEjGF6PJx
GRz70bY3/Jf6jYDZWkTxZ2KIW66M5lBVqPvU8+pnfiozSrZ5+iQyoORe9z040VZH
gixWeJ2GN/0RWdN9RWA7jlyWARwdIHL+QAuf79N/GpV/CrTnq239egWSbhhbX0rd
T3WsaiZVEs8ZxeAgYBshjyNvfFnntjieksCQGOWApsLMsNlI8G8prHJ4DPWe78nN
3OKu7cs3fJTN5e9mj1YA51B3SO9TjWcn/obOKGlvb6lcuBvqeBYfjUgnQ33TNyxc
lQXIy9GT2YDFoFWp6gDWEz4GmMX2dPAeQRc6Lgze58rek7dpqy5+owWD3+fNwEE6
kMC1tgLAX0Co7W1ahGCsPbnHotk68sWkn+vfe0UGihKckavPBDknOsMBKyp73zzg
/+yGJLW1187Oaje9e0eKO0+6JYMw1lH3NRfCMV53Q6l558JVNIzyug4sQUUtPQ6q
kT+57KrRXm3sMdiLIcLcsOSH8FGdklkxE5kUUyaSXBxDRgNzLar/19ikzBJwiahP
f425ObPXEKzk9QAMehGLvpLFiv3fNW3KtkAxPmyBlFaoNjEfz6AqzdClejPYlzov
lEXV4+u6MI2ydtw0pe8yx8We5ME7gEOKxQoiCpuntkjyx7I09WcvwynS4IFfq2Pf
gruNphfvwpYSsWmI1BiR9j6t8HAOq0cZnH9haDhHgn7VPQmTWv0DhFQzV3XVAfqG
m7svhCWGCw2lwWj/qZ2buwF+F4pOPjYJVRdbjQoAhP1odMx77oeiYCljvT0ja10F
ySX8egiomgm3K+D+FgZN63smwYTb3+sPDS3tkbJL940OIya1+BDc/vU6mRS5jU6e
1KEVSmzOD0YlloZpeJhLktrexgF/wjetMSayKRU8JBoGB6/y5tQGPPC6hoPwkwHn
axLPr3erm93JqDkSzLjiWJtGAkm3zWnITi5NLxwNJ9Fj7cVC6ioCcOoy8lQMykME
gVqE/RFtOnCG5P2E1EE8b9BDDTABFMTp4PA1zSX0BHAhzmQVSZzAzAN/il6F9kKF
luezs+h4R1vuFTgnTHSLm90wn6DxN3Kxr94cBGPakVjZ5fu7hjvkVe33/2ZAgD35
rHjC5IfgU/kQuqezvQBNcFGML6/SugiuAVwqieD8vgbIGEvAbqE3TSNU0Ke42PL3
w9ORRV3mmIitYvAFa8PsAcOjKyzbzr8LwT8BWtAiewPYQXBoCnrOWbQfl1+IvsxU
rpRGhDGI2OREAfz0u4Gf2EOp5/7ARY7z1Saq4nHzkQlJ5468DCvS/a2kTF79VSM/
5a/xsU9fbbLlalYVOxhl9GU2vuyJgUYv3ea8i7oNbqs/jACcb9S5AmdPc3i1tInS
lx0pG5ZfpY9Ig5gu/s9Si4ZvVfjkONmPP3Y7TyiCs6L6KAXuBTmJD8xWaC9aXjez
QQipv5Pmn03TR9x5oGdfPxtpBKR780za8WF2JmjHe2/hJnT+tQTFQmMzoOhxxHGB
iyTC2v5mqVrDef1TixogXbTWlWFvGlOG4wx2Y26z9LBnsOtOoVllq+DH6oay3gk6
oz5bJJaPd/pgZ1tFjC0e3xu35TuREDivDfmMg0y+woUyN3tWer0LjfyFoBJ1AbBs
kxjdic0/7loLbnk7LKtzH5srrCi0rvuuDV6AKd5Y23NjgCMquyP4kFu12RFH5iCx
xZW7I7c//XrCEYSPJ1G65GbY6RgJpO+nx4VWouygqf+9yfr5oOuNQ1Vr9xDWoU80
lksUWoxSkLinBEnJl/ltF2qj+gT+VHqMqXQWb9E2kCow4U/5gy6gA9KGWklnnND4
uwru/dO/oK/ZUygy+u+Ka/SQHlcaaGG1wdBkiO5iHlDgBag5BAJHQWX5VLN8dNY8
NdZKox0TxsROg+ViojmnpjhMwRGHdIQnUydjSd0RVR66x7TbNE12laj6ngrV9qXZ
6nNpaUMhLnjanp7iACD5FWvMzc2xqKX3WPdZSPtHHCK7QyVHjFxVD+Ap776ayyjj
tYwoZ8cjZl4QgsuaWXi7aKGHQHvuuDI1w8DOUDKmhXiVIFoVujcrppz0AIvm0DJs
+GfFUdUJNuI55TUKx/N4dYElklz3GQ5vBMeXsfYciBqrncTDiIiRFPV/Ag1LyUWV
qylUzTTxHig3DqYH17eqzfTkhhIUs31pGNvtj5E7ZTTyTThmw+IUO8kq7uo2XYZ6
lNEJYLYVHkq+bFJxVeyAQThvmUpELmy7Dl0jXSjmL3rdt/3J4aTseajhcu0cjqov
o7uYOa0EunDKuD4y+V6wld1v/ZHylMw9XO4Pkfsj463toYNCE4QHNM12ccE0/cmK
lMOZm4L2vEkUV7a/3n6/QyJgIgSzGt5EE9erg5F86470470N1AQj5ZuXP58QLuEs
Q1vfja7J9kHaIMwuLy3xGZ/efJBa9Uz/x6ky5iWt/hFi7PLenWY81r4k2jcgB54X
t9etbn7i0Bl20EBpsd+kHlrnLiOUAzVdjRhBNlfTF7nOUdYJlVLzh5Vjfi5mdz2a
S0oGmktDLBxC4mrbbLnv/8FCEtkLIPaK1tNXC9zrFDFA8dJsT2s9ZfhGyx1tzgXk
V5o7pQvKmyqtvr9scDbfWdbUPUGhEUfEs8Dx2T+h8SoRXBR3oALUMxG2pZGgaSrf
/VEmkiSGUgLuGoeqxg1DCmP8dblrOfi6o8v86rWtw0ZdtH9LLxWIJv75kUjMrO90
yyQ0jiGWH2ajFh4YZeYh3omLvF2nWUwYlyk7b9BJeEBnblo+RCuNj+9qAQ40rpEk
exC6OShbV6fYRmxUiKCME71JBWkSylpqdcDXphGQRbDXpn7ZcCfARt8AoVWlBFrr
1VCY+lNLWnpvFa5e51Q89XgaAr425nX64dTC/3F6qslgd6q3szJyTIa4HNw2P9Av
tLRwWSnVBNEpJAM9dOSITFaSFwwOkpd43rC1jNjjtCzUX5Id38pUEUwFAiFMq8KN
BIRbx5lIGz7d0VDbHttJvPRNz/tFqD1VDMa1wTD2vwnYvEf3czYYSr6sZuP4Hs8R
mpaoynYKdFkFGHGheyr/AzrsCSrSSbLaNSC6fOO8KH9nyj3D/+mwOn6qzdPMNyaQ
Ok6Pwqfvs+N+E5yIWIFXBnvE67xmntFw0aVirWY4WZuwqNxlis7zi79Gbu19MiVN
MfoxHMWIH4FrT0K4JaJ2gy7jkNdg8j6eSuGbHRtdgenpzM9MnwPePVeHTa/XtT5g
yJCyZg7JREzDHn+IUNOGxg1GHglZfr+b6R+FfsJ7MuiVA3obEUfgx2hkMZC3ERT2
YGEn+dAMJS4yi0kqxWIMl/iQs42nVE53k7zvX/mMpuhFj5x8p34qT39+TkI9SHVE
tg2tVCgFjLf/S7BOPBUcOW8vw0rMu2GDfhzwLX6r3HgW2F1KXDEIEFrRI6L+Fc1D
iQ39/aSsjsfjUon7XOj8jH0q+YVExuPGkzpvtp8QLQsKsBeaTKq4tbX0MEZBjLbp
By4Ma6QcQBqVcvk6sVK4Au07c91mfYly6WFcMvy2IPwyyR7e7NM7ztj8UIFxH0F7
+OE5iT2RxSAnX30okhLA72nrIwqgeyGjZygBVoxOqrSxuZ8CDg5Hh9r7innYh6Ps
3zMQl61NnN3ycDjiAzKnP0X0yVCF5W8Dklq1/1qtLGEdtE94EGoptQ6sm/9mjSyY
SqXiY9+w1PVjvX6WN8e8eYk3P3Sq9IXOAfJqmmcQKZhe6amPUfBYO7IWgILpDAjG
f9Gh7d4AcE9rS840NqISUolz5K9Ay6WfoV80I0pidHVZSQVYy/GE50Fnw0afno7x
5TAy4PobOQEWsPEAedOxeqC2Sok4yRpC/SmO8rb67T7RpGMjZgtrZ7ObVdTkJqcL
L17Mh97bUBLd9Gs8sj5QOYwkznSV8yczkBpUitJwUtagVnBdVZvy/OsjUvIcw27x
edYj6HMorW5+KeZWd5XBfaJ/c/s70myM2+2z/zFf+ug3e+3KdzeGAr5tKl9+AC/1
E4YlIRvACT8oKoVkqG4/XlgH7z3wrZRU0wLO0gl5NTTiOw/ccAj6XSe+uOEoAsAc
HbrLlk/GeT/Q6jA04l6qUFxPPpI9umQXLSW/m7TABr0NkCm7keyKtXnlNEmt9o6o
xg3fdG+BnbnZ9hPURo56oGfaUscXLe4TOw48NPsDmDNbn++9wkMW9q5Isa7Govqa
FLVCm4rRH9ehaDXnOF51peRfgpoDPUZYpWAQCFQ73y8IC2si2Dty/CS+rjem7cuw
1ZzFr6tM3GPEBLMfZRrITOGDSFady5eB4fq6sp6zZAvk6kweQDMODA3UE0Wt5os7
oBrKRdsubtl96v/jXIAXL30rRzKldkIkLFXWu4bGh1h0Mk4ALCWx9a7jr2lcbtMY
X4IWftAFA3az+c8vbM1Ei7G0lEGWteNboLC00pCHYUen9EoB/q6uikAGwaibr0zh
Ysean+SN/rQWMc6bAs9eaOnxcHVGPr9dH7nwchBVaEu3jKeCzew30bolMQjcgspa
8SKWYLTmhWB8gfkBvcgxehq1njRo1Zxi1Tha0SJgFkSDTRH3qUxF9eKPPDPLiM0S
v4aA25Bx8UXW+h3xTwq2zpZ3T8zr9JDI7ADcniioYTwzP95BlwBQpMUVQm7DF8Zj
IAl7ZMr211G4Gcu9eYQqW01J+ufFJf24cm+sZbyvB1ty/Y1wGmGtp/d7dwab2aQQ
kYRBcNukSzt1x0BJai6ltwDupHujSvBaypHPIi1jKDt5cFKHJcWejxMZz43PK+ic
UR7YI1/CItXDppfznrWOy9S3436LdvFqo04pPBx8kS9z4Hrt5NGoRWxzAQSUuXla
qsWJBzc0OmFi6MR5xrKLA2EGeL41VLGov90ybTrQi6X2ZA1g9z+V+Kh+zBqICcHw
yrNrtT79C53Ii012cEaGpfIfLuO+qfFD6IY9owtqF0E/6R3nsvsfJY6MZcL0L0dp
h2O52vKa/zxzVlxFQLsArPItcUBX+4QYvpbIg4RWcmSdsO/bMAH55VPtNjpHnjVP
GGAbOqWeqrs7iuGrjK5VLztWgivr5Z28kxaAR8bsHkZKQHJgCpEan6rqdJ3yZ+Cf
IPPGcE3SY/4lnQaqSKaoeBjAUhvLgbTU+a37q6Cfh5sh552E4C8ZAYjDri+vfTDh
9oiVGVEagQWBfhoaEsL4PZiQKwJiH4KXCVmzmYa5ZedCmfAcrdBXqpYK/z9RcAoU
6HiAuM0y/yUrXCITdBA0Ra+spfOVaXslnDCioB9ck5Q49yIHRWdLiTm2ETLEZdVQ
IpmPQJCVLvirGkeOyMqrG60Ot+XM408qJoaULFA3ot+3vZ0WxcVsaoBJ8V/Xk1TT
9VF3bOMviVXUQrjtRPD+lU+hT0WVjg/zyC1/hEQL7Mf5PhXKlGe3VhvB/aaFGTnS
3AoOIuwYlgRkI0YmRTre417qwr1pG5833En/umHVi7T04l7d/FQKq+N+oBBFQGWk
DjteHJUKa9YvfU3DLK0YHEtWEOOu0V+yrTt6kx8vt5Zmc4Ae+JsdnT0+SBWkyKT2
/a/mEwlOl70lU1x/3OYruKy+Jv0O7AlLkWioLAQlbz/LFr9oon4Q8qaL01u6E1aT
1zOyvKEHYIrAKmoN+sEhQYK9aBQaF4jlK+zEYFtZhGPTpsLphOnQUgBr553GrgKW
BtU2PDiRMmcdQl1sCQAEqYkpzxSRurIWEQ3WvJLDsvJ8Gwo19XUjHlGVNL1PWzGQ
CjEwRp8EVczKqas1vbFmDGrNvizf6Fhvcy5wZYdxg83nCKA9teVnoCVNBsIFOcDx
hQXS4QBQWOR06kq1f0KDdNVp5WJf82nxAtNbXR15cI/AXFXeGlFYBuvb0MhyCAi8
dqyWXERsr+mIcLTmfqYTLTTnRKmYL8Eu8AurXVyfhQm0fO8HDGrU51SpyvU62KyT
fqiD7GI73pvW/EwftvThuWYd/sH8Rg5BZ5/fpn9AnJozioueG3ezdfzgVmj2lJSZ
VSk7yXw0v53D8nzVasjjwTyVdWzC3uaNQBGf33lF2RnoNRoIIDfkCTa9Ysxb2iD+
KC1oGslC7HwyMMfAGv95izh04FUNAPU/aRrbZgKopvgfMfAsV3Oz/bBVLGYHk82k
c5TQ6CfZ2q6nATlUXRJVj1uAnG99+mlMctuuDcFnHVoqN8PE40pRQWari++QCsAP
Ke73KvAjQDK9AtAV+teeqqFZpgKtr22gPw9q/iXNTA1d+EXiJmziv5RrlhlvluVC
27Bg5DvYNUzNwMnsh5CCs1ar4ozqV6ErB78IraFBiUy7lXBTR2wV2t0Iq1DVGPc+
gYcBxth95VHmU2VKFeJM9AVHdcIFidkyE91TdzT9oDeh1456YlvJ9euuZSaY+Dp7
4uo0Aie/G9TlnTPCiweb2vlIMAoTP33JvnxYXK8zzhWs23YdBZGAjwk2cpU2GsV/
Jt2zOTPBlAbRiLpGfF/i34xI4WpXqMzhBmFrhPIN1KiQpX/tTyr8Tnvq8BRo6gP/
9U7EtAoG5Z6OS9/f6lLzAeglg9lx58st5cXMtArMCXxFp6NTB0Smovozt+hGk79q
86W0QK+oQNxZBCOR5MH9vCRM32iHdNHnpUoeya0e+ZUQ70tMqQVXGWmOigz5UHeW
+2xgCLQ1lGfaUadWqwjhBCSc5Nh7Hzkm0Ttc4yC7Qu3wFDG4TMISmwovCiCm59Mh
S/P9NTBjMUOoQ5pYu2Xikvllj/pHCkN3fnRkg/Mc7aNCbUD34rKf/jqWWz0ivNM0
iufHMEGA669S5ARRUbRIFq4YCOjKuUwhIzOgjqIeuxYzIJ3Ut0uC/5C2JzFpwpJS
gGQoyAt5jwQcu1cRryWA7FSo0zmjNAvHzl3lKkiVqOzUjQT8tdIa2mJouvAdTlF/
fwFW6gK4QCXiYrMuFxcLub12NvrZz8yjHclJxjshmz1iT+mj2gA0FpLA+JXdsvYu
S2no6iRSn00Oazu4+hE75fkacHsfKji5wdCStv6Hq6AEGhd453o8ttemu2XfCsRV
/VWLBLWP3yk8MFDLMTicu3Wh3980PBRgwIKsvCaqpGWbadW7f7oVmKslR1Gk00xz
sVNXIlxTL7/8PPk4W5S9GhT9DhVwYfdknlVsUbxI8qwk1D8uRHspwOLNJSFUZLVq
r9fKneZGQlfGLaahVt4NN5QDCS8qRcIf8WJ/G01fK09tp8yEn6zGShqOyUu4kSfp
ve85y7GtTMnajK1yGZGkfm1Eh8nwuNRVTUzVWaUqIE2RJtWhpmuDiLOPYWch48nR
SsbTd4g1pb64aqrZgCqm9oT0h68Qteyz9dhBCFJnwge43SD+QsqLmMpp69ZNdBgf
gacqETJrOXbWzxGSi2qzXPeIPC6nsHWzGT0J3ycrSWBkYmnOMqoLSDTQ3AmVQEHC
P7idT1/rZrjnoSF3JYHt4P1UDYZcTk3g4NMvVcwz1KRK4VMhFtu+SlLlvQ2JKoYZ
kPrB9xorWi3DTygIQ1Q68qH66zy0DLTC7LnKHAJBExP9mceqBKULTLq0YexJqh2F
32GKTjiPo39ef810YOkAS/j+osa3/jKh0XOxAr7lNKEylalpkIeg8t+scdPRYOI6
DFwSCdnFP/OV06/9HBFOEGH7Da8IYYGA4orC/O08wSCLB3WC7SvAUpeLmYNijFOj
L5CfVkYPqGPg72KqUF4g8ZEVGGUdbtYwLbmNvbz81cIkBIznZl73wYoJzg+mg6So
hPs11d7A9hRuh5nk5+hYuJUz+GIvmj+qD3bf7ljXJhc++lqsGYPgVRYhQOnDwsMW
P+2S+HmaWXJmyqJqNvWJe8fBWbuvvKoA0JDxsjVIchcNCKvN4WbfJ376yohzLa6z
cZSOV3a7PiFW/zB5Hh6QD4GHv+sF1X35HUuIURpobyPDyHkGs1HnGae6LYqD82IQ
WUyjdW6LhoMdI5KJjoMnAjr1CUTJJRAsjctodKG6P0N4QZRMr7KNibWbgQp6hxQ7
FrdnRwe6QMayRMgkf39K+JMoKL6B6c/klCyIBznvCWW8D53jcz6NHGxHqTYdwQg9
kQ4u6CeE6VybIa8ZVz0sW0QAbbAXXlXhKTwVCR5F3rTGGOCVx2CSMsohC55EEL8C
N5l7QBaRN/AOcpp0FRRrREs4k8SBd0jnTxLzt0vDdBJam9hsIOYY/7Ds9r9hAZgd
5gtzjYr2qEXZedBnt+ONnDT8+FzkxxPRthLjVP8JW6K/3JQGTaXcpHiLM63SLipy
c6BpIPVgxgbuu1a/CLBYu7wEKzyPu2Ad6+QiAndmCqkK5yC5a31lS7Y6Rz6QMjv3
dxdpSjC+5KAakv1TPywLrAfKT7sUFwHlBdQ/qbZW/6NhXem4NGagvInqUaX00a0c
gK70yGMcinRXWqzwTF8L8eWWx9Qd2IVa07KBcL4Djenk618FHo1b7uoAB6Kt6vsa
daW1hN5Iqm2tX8ubbhhzxPrQzaFuOZHG7q5yyJto9azzipUvkJa5kd1dly/4mJ0A
FKVJbUpW1+4gZrNwmR9JfwRwW5EP/Fzemjz3D+VMkja/rU2Lgu/Aoq16z4o5LJs4
TWXGEFugBssXfk9fUk3hHT6DfG8kCazE2eD6I6YXzUj4HcNns/hnp40Usrwi4Bfm
LcCWLazkWZN51pqGNkEgGCtq5ehSjqtphcimqQ758X+4j5azcSePlEe+GAEJBojL
F77OIywMoTx4W0r6VvBCCSrBxNW0YZv8rMyXoiWlKPSnrfZy41Fdsg73efKB7NCZ
Wcyvn9h+z8u5lW6Kt9E82XcjQVhj6joq3U0xuupyYnBC39lVHYfgUrDcnrLpmXru
hVUnKOwatzISucWlyLogUP1qEXpXCy/H354YKx+NPEZnR5VO67KnjHyNlCBP7tBV
f5jBZlgMiOtVMq/DmFv4AuDhKEneIIeex9gWPpeEkEOCighe0ONoys+zIn1GZHeQ
xmmdFrc/gvg1UepkbyPzKf95kRxTDvAYdMpotw30kXOo3Q41v0ACx4qku8l4JLTD
Il1W3rSD47y5b4UiK3PrRwfbHKwpHgvFKi4p09daY4u1aSACvUEwyIKNZWlwJlVQ
mIOlSgkNdhBuxJhukr25y60Z4Jl11N89PodPXtmV4VYtKE0FrYK62RoPw/F3+KK3
sj+L165MZXRvRs+OTiEovFUs/EAc/DsNIR7BHZk8s4dfpBds9vCq9dwgT7s5BQKy
2WxE2lSf06l96MJLX6JpTKrbRkKGQaX78kOeE/hdSl6r9mjh2YLaHHb34syuyd8F
SRLLHAezquNhzISc45pPdtVqHo/vJy8ijkPPftElc9LR4CQ4Y3fmKBlJ+KMw1Zsk
EqoFBPCUU6dRh6q+PBVHi5LVGRegaMGC5R09Q7j7A47s2l2op0CDABYHv2EegY75
k+zZKVVKbH63iucVtWP5uEQhiosMdjGNi8l9hq2NfljSOrx6uljrpzjCpwEjDLeK
m49rjKZ6Q9WbeYNYg97zjxQFqcGDedAcSV+DB79mgVktviOuwkYV6rvcAFMbm9v6
wvgF0hU1ZTzW+FDbWEDWQC8zz5f03286EbAWMjor2ZrUintgIRNw6TkZZwURaCUV
39JnqMW/NX2rKqWbFSM9whNTZdhtEv+c1eXRc3XLBXHXu9U9LsvZVHxbM3Xyh+8A
gbxlz6F5Tny5q+butL6VlkiJvkp4gHQgBhxO98ws95mxfuN/qCdKZQEbEkChIMk2
AI1gwy/fLOsy/ppsLCfWBQ18e+RV4K+lcVN9PtvsrALRsoa5vh8mWfsQRpsMiLbE
X1zPYKpCUkemFAuTJDyc5Dmf98CotCM/BZ6xpMQOrMaBzXs+66/JkJJj7QmWie2E
Qic7LsS3x78jjf1Qwyogllg1R3x98oNwQnRe4VSr7XQxU6ZMY4c8NZDFFJZAxWhT
sInR+TcIcqjZbAP1Z0kArLIk7FhoX85pcBkiqBuY1yM2XdZU6qC0ShezTobCWiIK
DXLpZokKkdHuKbA956rBE+sbqxZxOZhKz9eVzUTPkJBxxnHMCMVr4huc6Kq+R5Ay
SomfKo5J7+mOXjl996cGv6Q/q7+8HV3ikeLu8/jVfcvUanL0WR9bCWWRA0/s1kAd
5H+4oEH4tsk0K/Bi+ytoNjh5mC2sEPQIYuhYb/QrliiIAS5yiA5jAiUT4ciNYNUp
7YcjJugz1KJnl8dI3zqDVp4AeQtkXHQKBk5uzOCEb2z1ud8zTTjiTd+UzrPAzNdd
zvVgpzpDOPqzAlAcYLjD7jkkeFvhVMlaqEtciH0JzzvxWHGUz4XyHLqrBFxTuEPm
Ef2r2q0y50LX9rs2t5AW2ei1S7eaHKtXl9FeAG/0sDGH2IS9ObzDR/Wo6PaU9oyK
UnMF2eiNI3Ebv6T5Fiu3uodG5eWqS1944WLhYUwtqp/aHoYJ0NROafrgIaAeyvkF
DqxfhE2ui5pQtqv9X7lHo9sC3rfjTxYzlo1ZvFHKyc+4fZBCPx/lxIH/IxMHepUD
Zjk09DSNV36JIb9ehBF9zWE/iR7Q6j8VK+m//ncOLgWK8aXyDRocpysUzvNWZW+A
19IpGkFxKyuO2ILuiFSh//JvE59LNtu+Jd9jvnXwzkeXGtoYI0nJQ9mOK6q8gJUp
QiBgtIYC9ZiowJg+Mz47tKhtaJvsqo1hCOARaKfag1goLapNYYJ/ea+kFuNHy508
m3B1ZJKZaKJ6ML0v/rRIrVgoB9HPhSJ06LRSa920WXXWhPkG9+RXvZPsspXrfuUW
layfB3yienisbefXHfHcUC7+uml/oy8ixd0bYfi64aqiGDp0fcFkS1qG/s5jzkf0
iu6vgLHcJ88nWFE1o2kEtxPqROKyboyio4oW44UPmvb2Ri+NNQlB+cQbzTmtH/Xl
VVYNTTWCf1k0qEw4grk4iOwZpjb5W31mzh4AyRi+hUwxGwEio4SNK7IYYjP9Mspv
d+JCgG/17DB1jySSCMlDAAsYPjfpsBdpxZPaW7EdDQcUDbXYthllN8AFphMqkPyi
xul7GCEQy9fkPxufsDzT1+AXozzTWXM4LdXumyTHOlHhQ886rcQmwv0FyPA0niqD
3ienGreSAZg6+Nv07+Yi+8vXNvxMQKt4W86FrIjzqLcAZhXhWLx2abxVeppk6tjw
+6LnJluL1vn8tgGkifCT57FAP12K26CzlAI2aYf9ASuqFdG1379b3CeRBeBF0RUY
LbjSBPrUWozmvKPLPgfB/u1iYZXZjdMk8jL3xuyWfvC/iJUI4jRMCpPbRNTSDFqo
6EgV3BKHGt9ufGq1BarqyupOFHd0a1zJq/Bz60KdZHqy0CqKlTUIeiIkdhOlzBwk
KfWKYOUkGySZruimbCOjqqUlS6Ad9aX1Fh5nDasSUF+lkF6B2MRwo7SP9t1v+EyT
f87a5r3xLYtWE9t6vkX0r3/XHXwLBp3G9aNEq8gF+w7v1TFXpspEWAl5ROmbJ9d3
ZU5ZjM+oZ4cxtLgpv+1eiAgsM8iepo1cjLsWWh/qhr73wSsEwwLn/p8bY0b55Ugd
QeF4cYrCHdHsqsk1J25SgcGz1r3RSU/MNhjNbD1UqeH1r85oGV2hZF7zqkUVrtyi
bFcmUpSpXrksjjdO/TPpqAC1wP7Ax6oN0/miyoHfpcSE9cgnV4KCjyruE0uXMsri
YZ0nuqtq66NHOQOJtAR36nzMGcJVJT1A91j4PjeToG2onyyycSIeGpRzoP0Me2w0
omFWnH3SxZxSPNVig2zasNL0j3VqjL61t9Gym3/8EotvttTQHJ4UWMcdcvWKF5Ch
kEJk6K8WV5TFf4qfOr4rjL7NcYVS+II18q2rY3e6JxHg6DI/aftCasB7IeMOrfVH
QJ0zSsB6nqED78Esz/icH4iOBNuq+bdo0jcpNqeLPFPAjWT3wbr6wmNJe39WhjqX
sofMY3a/B+4l7Y1sQf1iVgV5vaLSeGOAc3wZA3Vo6iUyjtlhrt9V+ddTY3RtseV4
u3mckTIEcBSmlXSkHc+uHcPwZXrtxXvppw1tq1nDoMR4qJ0jYoh54GMk+bYkefUM
dgayylEEVysuI6NQbwmbUkIpvpMEYF+0uz6SkoNTIeVCB7HKW8ruWbk4OccrcUS+
akfiry5L58DJwyBRZqLtLw5E9FE6RCCi7NMnNNaMkZe2o4Of1o3mHMFvrFSzTaQ9
V6hyKrUOblsiV6BB8cdG+OpVCEFxkyCwo1hvIJN3aav0HFq5OJ/P2ASmLW6ZxQnF
AOl3YOMul6cfmuTHmqPQJZIDUQCx0Qs8LlJlzTcGOoMD6VrtjzkPgPhknqWFgj5q
592M1iaBYTxiDag6EfXr8QNKyqUzGMpqaI6RwstEqlnIXwE8kRq5LXk1L+OMFStP
UTIRh3Jt+P3LbjgUQWaO9wEp+rt5cjnjSSJWuIa8tGvuBj/NxLawIweDhotRYFRH
udHnThG6qjL8QWBis+vXIuGCne5M0HnWnHwvRm0zpm92z/SJ1ykvBVfj0+UeFruB
rP9CiFiOZ3IPUBw3dAQenlnz7kiT9m/7lgVN6gOT8h5tdQXMbbx6bD3ntAjmg421
grs5OXfUgM58FjDvHt4Efs3EcQ5pq11KTwAoEWdFIvcXxIARgcNfcm9eDvfRDTvn
OCBL0AF9X+iFPMYciXOrDyvjgecnCp85dw3KnWfdDS/Silz2nBA54lVlaE9oA2VW
ttLI0Awb1PtqyCXZ0dOdDOKFD2888P7enjD1tyQ0Bqa4DzNiY+QSh7XgPj6PUEP+
jmE+QIUsboH1aS2V70hCcE+nzH4qAoxQHGex+bD79DElW2/bpGPIltAzNzwL7Xhg
mAK+8vAiyBLYxEtwB8KEdiPTZsXWuqgBsSCoLnJxi7Acg9nrYrCSLE6aJZaDDtDg
qRLNq10MHFPOcVLGnnh4dO29ILSHkK9LsiAZc2OguAjy1v7jkVu2zmwiCWQUJz3w
CZF1SEtsyolcskzJ8bBeRYwlVDFx92jEfkPBlIS9hhZ6nQwfEI7PZFlnUhA4QP9z
aOHSA6qbvwRieEwEuFwY7vbTo+Iex8EpQiNX9OdyowfNYztMXDo4d2RR246H+c3i
bPLoI6DpDTIpVmWuy1u0OfEgTMVr74EGfb/PVPLQishFz5wyCGEov0k2U5KpbqVm
c4PY30VdpBG7tpbFz3asn0lW5bsatAvjmYu0TRLfzg5lqZD6YaHwatzzr6nZJqW3
vDxYp1uovohZX1vgez1DWRBdaDdcFplqBCxKx+u83EA+Qf0Bxzn55E4YnIPhwQSk
gH6hZ74ah+KOKXv/ETqmT04sUGND4URiddKiIYgeCJIEXo7wdtw5h7ywKY4SEsDQ
F8cNmy0IjUws5HYkx0F3MWs0S+mTgyqK7DMCgHzGmMoHcafgcMoJUfBnp35+dtAV
pOReHphO8ssAgLMR26w2uLGSTbttw/4dOb3F8wu/Bfh/ijg/2LkJ209U55F32VQ7
UVohznvQI5hnoICM58VEx5x+VoHtiyAuoMIxLMTwO2WNWMfPx/RNQwfe2O+uJ6A8
8Ctk9rDEgHz41bOE/yVse3zc2zKKa5THD0FjnSUCoqh6f28pyTdsGguJGBS+WRJ3
7tCy0zzVNRWV3dYkA1qATdC8kj8paKGfo4pu0iZyG0ANbK704QCcnaMzM+fvrzLt
7PKz2bOj/SK83lRKVdlJGWfu4UkfeLvfEdWO8vUIiJAvNxhdiTZcZkFCm16KGeXZ
iI7f9p577gPd7SjUzGNXMYCy+uhLWWIIIe1/tXLRBj6kOuBZTK6hu0ReU+NqePT2
N+YCTO8sKdKf4Ap5k7J+lknUhDBzBqQNwn9essoNppCTWvedJicxVLk1wcon0QZE
cccQVzJylhP9WzLtuaH0Ce3rfLDsgwP1CqUBAOIcJznDlySg/Le/68ZJv5kkv7Wv
mqQLs/6ywVj3iCR5aPuakCMZd1AB4/dzCiVPm2qBsD3vZPIqXV0WPocFSVQ4ymKe
bgtkS2z9eMyzkt65sTX0h8nuVhT+ySUGb5MQLm43nKLq69ZIwI7nWtT0cSw1b9Jn
NkMs1Wu2NlgKC3mz5VOuz0wjGm7VMq/mjxRI1UuK0nVeQobB4WIid5vT8iD9CBd0
P83qSwBCHOT5IyC1aPoHWeGyGCmgDmUSGYJCePI5NXgUaxb7t1b8OrHNhxnfvZ1z
kQzAFwC2X6kn7b0yYRlFKmfSpVKIzWrx9XQBWeXOQEFcfEEc/UknG7l5gzWBEFb2
1HeHjOVstF6re0c+ZRryXvrnfCKXtn5ImBXTDCWdGulJG2xSS2AcGh+Hj/MuyflU
efjJj/5D4pbxOqMBZos/bkEyBM3CtewF+k9vf87dv/CV3GvmkLmTV2FSdbxx4XtK
PSiapgzlN0GjRjGtwFVy449c8lVj6ODJaf1/RLhG0tnD+M74mNy4jK1dkzHiprk5
jQTzCW/p8If2TfovyUsX4Zeb/DgEdz+jROHzfzVWUczJu592wDFw7+0HVdWnSuSY
qhfAd9fS/ZeRJ+XDliMSeGg/zTqqXap+T2DpVFBNSv2YgR4wR25A9IalIVIiVLMZ
1spGmMnYjxkRSJpVaCFMFoKj54BldGUW01Gu6W2StKMp5xgkGCQvyuxxWeCUfAlj
1OfFlnVN1sbP5W2+1A9BE5iba98NTaoMixAHHG9+TJfGJIbcgmm71j4WV16vattB
VQ6ocQ6QJLtyeyvo3ZBL/IDb24AA9/SDO5hxhCzqHdb2lnhfrbK78SxQ1RV4pr76
iOMjmDnlTm9yHXSiSRn6whifowmExt7UKtDKmuZJGQr0o95BHAtbMfMa1vWj3hxF
NgAlEdv431DEr/jzTZZbeL1hEF3/ZBK6YgzNv7c3aftn7X0S8UVa6Y3YWN0rQeB5
iw0fbJ+anuNbi8aZOMXGy8EPGCMf7LCJNmk+N6mTVJ6V3W0vVstgf2ZhJjBSFf9P
RjSlAHSuB5bvRBJ+kFNCHlKSJdAouR3UrrtAMINduKTcx3adHZpqv0pUht9Zrumk
J93AnXPDSjGLbpV+DV6AKyH84HFi0A3atWkPd/ybpHQSwBPm/LyWCeJICtZ7KZ5S
h8kpTbzE5l3ZGVxDAWMz4lfFTwAl8V3Xuqo98ibUvdrDX4EmJ7Dz4Kh5CUPI/izK
8jVu1gIps5eTGDLorQaZYl6jnNvbX5K+28Sq+VjJKND3dEHPO11tvJyX48SR1XBW
l6MdniG8wdTuF2izM/MrLc45GjV7TuCu4pvqXvBXxneoiQJfAuQSu80m4yFAQaxZ
zooWqHtj+7cVs5+s0PBPXXHe185+PdQDmibR2r04CJrFxF9M2DyZ5pptztzNzkdR
gyoKlXP+/hxmS4njoaqgMCwABu7AiVvN8O6ft9TADGWznsSFD3tn/FBtPIDmLmop
EwIIkeY7yraH5b2KfcpVsyO11qWIjPHADtuBjWi74vH4foqKkxG9I3aL6vUvKf3n
ERzpT9mUUODNO1NxKV7xLjUocYdQ9lpEJZnuh/Coq4LJQoacx4FZ6hQFv9GrCxEk
VUIKtzoIodjqNO9Hqi5I632M/VmGdn3/WV5Gwgv5Zn2bjwS/y8NJdlduD6kxBTRu
g4aolsuXvSTblibNirZeilWM5bMUa8WAD5j30r2inY1EXEinwol3wbdYmpOzHgKv
/sj3/rWyxIUh81ZFwrxdg48QbW7qptrvSnKeK9BYpvbkS7q8F5d55fG+3x7HdOfk
9+BIYdEJS6hcBRLWdY54WBfxMd/OWk5cKJxVENvSZ0iXC0B0IFBwEwu2/euA3O+G
+6bng5Lq9euErgk2WVlPU99MWK4HDNkfY+drjMrMSSt+wIARKe8Ibz6z0r4MVJGu
cKzm47BTAGRIuHkk8i+ZjDfdAnONqYWAbEmKPUkAu5NE9tgKOwBpoyk3XYvMemys
tS+dhVUODGwlRRHUZgo8MQcQwkkeU7lVapv1CZdJ6G9A7SYQTuH8t9d+iToaUZxb
d5XwgEH42u1m6BuXdspOyQ7vn0JWt0HhsJR3PzA6pAKENGTGW2nOjqi0auSXdfoJ
/YbSUX48IoG8EAOrSK9ZMA8tHyijaXCeZ1WsxcBil11uOUkpJxSx6/1yRCAyPRZ6
pDLHXJmAALdBzcvVrbV2tzEeQksBOxIZaT/a+XCxsW0cBy+o62XdfnhjUCI6WLzP
a/y+weSwAKVdAMWSa6dR+YX3/aouilr6SrygufPxWMcQHDc0UynmRvY680w6kbyx
ZY0fCgKR44qNI/tyxz/YNENMaaDYDazvyHclVuabY0LKJ6AzjnKszuLEk4n72wnX
ahbAbZbCSbXwgjmxANorE/B6BDV7cL9wqXloml53k8EgS/HuGoxbtJ9WyE1RDc3m
0qYInRwNBddfChJMaOF1uz3z7Bhz4FBFyxl1ucIcZ7f+VhQ/prBGWIQA0NTrm3ct
5byb+YEb7JHp/6PIxRe65hveOIrGtGKH2EgeIgqGaegbBeBnqGZRfvs0LLU9tVsV
Rlso5nBd/I6iGmetAbAs00FpWk15Z3pjmZaIVtOUz0pVlWUr8qYaxEqzzJ5Tf+Oo
uvhiU5tap1NHwuW1uFe80q6Hx7Z9o2efTvRI1nLb2YL3HGESOrre2Pov5qp3RekW
EvQvREVM7flDjpq9a3Ba6B7QVl5WGaf4pG/mvtZGdFzATQgMDDKZobQkY0HYwDnn
IhSjVJcKcu+d/O0uf6yGk4Ycog4ZPWvY005T5ntnsB4Jb/tP6dxXXw2hSHBsjPY/
rVNtmoJO8ElnOhNMD3zmJzIUcdTg7rSUUUI9uyXvQtUOALjclH4oV7raETPVUsJr
Wpvw7R+yBFvziSBJp6gEobE7TcayBoi6IAn/XaxEqv005sdllkm/6lSNGrj0wKfb
CDWX0Nmi5XHOa7ahuRUEU/pMaIXyGddreF08kkZ9gJkMVB5FNZwyaW5ryoxMpSf8
umSFUoEoPATaADuoaw2pBH/QM9BUyt5PInFFh/X1WQDZQSL16edbdPmDQ6aEr0it
w/y2STtI76ivpCiWGcS4W/SlGekOy1lYSMKsMEJAm9wkAEE+4TdsDDfRkezevbPo
kxnmJJe4N7nvkccmIF/vdL0mijHs1Pai+oPLv55gx+OaGOIQt30tSd8HwEYyehZq
KhWto68oN9BNS3JWyVnnUW6crkDGOxnscMgbZmxsaLA/gCmTt4uKw+CzXclm5mfK
VZIRrVbliq77QvjlBVOK5Q3a/Y9HMswhcHP9vTRLP71ttKOEDU/3EhyAWoVp7+P7
X85ve9X7xgvtERJjhP0Z53GRdk9xR3Y59P0igDqQSAXXhHcvldG/xrjM30gqHZcg
OKA1z+zeoXvqKYSYtcxdjNv9vI2OyBtikhclcGKgCaqoXcbIl0Dtz8q0iOMY9a2J
j45JoZhvnXfLPS4kIWM/SJnPWwzri3MwBtb2Tl2gA2UD9JCFdFCNdZmHqFGhZDaF
omuHQ+1LT5fzBX1u05Ft9i797UullNBP8m5jYUqPGkumVkYHfVMDPGdTFa2ICJxv
3W6sVgtirr8T+154HGCB1/i1bGMD3qSVjV5jLo/CKEQwKgF8aaYZt7itku9BTDLP
q7K9jOH8D+U0ossp33LE9DEy6QDk7TNkUDuiZ7OKKpRxkQudhfg1WVrAYLPVgapI
OcQwlCyJE9Y6vKwrBggiWlIHCPzBBvdRbScEig7ruUq3SO4+7XqCuP+payz5Z9AP
Ct2/LhDDiNrjKhDM8Cm3z/KzN/QCLtDi5k9kuCOXMRo9cW8l1+q+fg9/1jtOBZL+
qdSMiMdM7HWszSDU8s6dOTE7gGbW/SdorpD1o1o3xvykZcX9CBEuCWcxEadXd4fT
Va/xDyXRcdN0f8NKo/6bgHBeACgswIbxvxiXFCDglFALyet4DVxgvbkn/IvckVW8
1lG2wtKWYdU2J+qKvpNo8FxtXYGVEzvMbiIUltYEdYUijhNJ/xqCH+ATX2mtcgkt
9l2X5LGDD98ezwPRErXvDIHi4iHQnyxG9bin3w27GfZ+BD09+YGWjwMuBzzIQrrB
5GfZvpiP2/eVWaUKFpGLE+/Z3yoE+8By8VZLrLLrbfG0xpYVygLsGcKq07F23M2f
JQ9gmtp2Iqd59Smw41ADB2ZfiP5wiqAxO16p4bC+YK8VDKZBU2NeBbEbgcZcXLGM
0b+fm2OMZAEATae37PH7VWlu0xtBNy6NnxJkcAnQ66BLemXsKj35fphjZ1YpViaw
tyoxbZlaOlMQFjTDYnmCwm+mC+SFAYTClLRvtVZY/6uxBJ2q92MMCb5R5/ZJlO7N
NH9SP4vitEIPxs40uiumdu1y61NfvW5o871nQ4O2VVxbetgf/jXnT8P/qdYNwLb2
pIX1Pqk2Ll3rwwZzYo2ikSw6qm+cuHbASRBpuBPvEe/tXCgTVY+Bc79dzSz8EBOO
wfsD9Rcl0oHNIaa+ENYWMgLY/zLBld95sxsISu1dJOxsJrO1rBc8OxZYn/RNWPE9
AQwC8q1vqrCNgpCJQ+3nNCZrHUw9qZ7b3opZfm3pcnZSKEsHgeBl+X9MEHL63vvh
IQWggY2ODC1a4ERgbEv4tiYlDGG4DMMDJjuZKE8ZICLhFWLn26xklJ5/3cRyHHLk
9gZp5uJZNzDSbMwo+UVjJDoUZ/ivdQWFzIc719/gUzJsljpOR7jIUPP6L3zR8tIO
XIW7690atzpuiZHHBKnhEY3y+hIO+YdK6K/SxDLc/d4IllkQ8AcOf28MsVxTPpwa
HGuTgboOXCyCfM0Zk0uSiX/2HuK+Lx53YZlqXnhyRw+/D2rLUYSuwWBVRvyUn/0f
Vn7cc2rnh0hXoaMm2h9WCoJImDl/fcrd2BEFz1JT8NBurtbFlCojnHwF1nW1gVD9
wkbb6z1oNaQ7pH55RCO4XUkXmGbuIIT2BG5DDK8UABaJzbk/EwWQyldK2eWCSd+I
k9HU//wrAr01zWRRFaDYZzRqS5G0k87nsDZi0Ad8GA5GAYTgbkNV5sLqIGiTbXjy
1yaipJ+4Q/00NoZRxiGJPoREzZ1sS/H1IzNYPMkiFBYEqdfPbBTKFmfejtXuTV+l
3aIiQwpgcBX3il6mrgJIEu9PisEWRvXb+8j0TkB4ry842e17bDNR/YTi4qGvI0+/
3KK2oWbCqpIZ0Z2Wzk5gKuzj2xae8PxLoe82+IDPhLuJ6/IYNjMEZVDWJT8q9+74
Uvd955b5jzXwu23tRZE3wAQfwTnOKUuFllTc4os4em4F5Ydo53mtN07lv4Yzn7WG
OG0sjbJ58VNY2GD5GjijV6mg/Bs2Owrl1aJE9ABezPbLXaMGhjGYVi0DWyMxqtIM
v8ZJicwUoBOV3XNsnimj8SABMJQrT+MajsD12yLe7VBFiGV3aHETZlhqfdBxIcZl
3Ou7iGnoTanMw/p0GJ8VKE7NOhdcSqDKa4uXtjz5ianPVU6xVfSrrBRqloiobx6A
BuncM55CwyitSy8d011j8NkXAdLFWzBOw3fpY4pi+FFsjVNxDac6utFF7FuwhT3i
G+lL8R4BtU6FtH1KkvMQ7vdI9BTIPByouztaP+ZcVYhV88sL4iv7ZDzxYINtjbDJ
SuZlcs7dqw25V7mFWeqNUwBZUS9jxeVI2j3+YO5iw9vnCFtakZ1kVmOYsPNZJLwf
tojw2+taByGlnbwf9XJuB3I1rj6gFkQzKThWpTV19eWGtPGna9A7wzirWhq0Tivo
S2A/W737CKTC1jj2VpvOR9hm44MggohddpMvm5bKNEE7+y6Nky/JD0rmEa9VPkm6
V/w7kPY/+W2p80Z6mS50LHyd0GjrLI6tBEQAxnxGDBR5aoTD5EbHzjtoSnlzHy6a
Yu2Qo99+UkNrRzL0hML/kr5MAiMHic3pS/7Rq8NuwcLyUCGa0bnk1wzy99fssYJ5
ydCXXdii+Ee2HiCHuNuxh2xbQxJ3C1YO8A/kW16rNPenEjv1gucYNcSUWKl7zZuL
uqszF7I+zniKYT7cTzNOue06Zvn7uDzFCGPt8VGMvueC9ly4yiiXRYBu7fgHssY7
2QsP7oLskD9GQ3Eo3tGJ5/EIW1bU0gWKuEwoTPYSpyfIMZFfcT0Gb+CrxF8kihLH
0Sb2b9rnHqiJGmJF9WWUJCOuwIIU1+80seQfne4iDjon6w+JIkgTfDGhgJK3wkag
3AnGzJlaUHVdnH64d7UUcV7pmc5eaGFe3fxoLA4Oc8nCZAD1SNc2tGkp6RfYClIv
qEvdRuqC3hez3L3whpZIa8ONewaB1lPQBGTdW+w2hcbHDPAYR+u4OolajWZBui8S
Z8IgeC4NRv6SA4S5wddKfVSnhgmhsg1UVrfBbMq6uSN9/Swu1KEDnzMo4AX221es
21+x0qkmCR9GZDqERU9KAjBoYPLG7MhhXDCbGDHGJDWkwzO6iKFA/Pe/13PNfpoy
S0zy92vw4IBc6/sb3epq0IGq59tW7D0t0PWe9opffHib9F4ekBNh5tVLzUlXPWG5
b7BZMgYD9Q3fZJUlWbRzwrM1tTUeDMfAeLvy2s1OlboVhz6mmBhUTPEHQIlHMJ9J
TrdNFnU2d6z53k4Qo4nlXtWYRc6Rg/JIiuLDGtJvrKre7O/OdeseDwBOPfMoH9il
NQBAoBgOgFaT0utR7t4CAD2muHqjbiaRqMGlAznVpSAcp9O3+ax67suh1l1u6uqV
byheWbI5dorZSwVO1sm7YcSshuXA0l4dM0Ft1NG3QVlp0WFGx1wNMVabAFGlziuD
Abhd8SVVnfaS1eT6LSzwvZxMEqhiAw3lrItVHYwMc1QTVQksApTG4baReV8MwyXF
T18C4rzXh1HSYT4R/l7mLlN2OXDOab3nopO0Eu5e5P9i9aeAWCkI/LvbmzR2Abpy
HrI2s5j/eUns9+DsSOWWc5GWj5CDXbdx/LYmITecTgb7sHsfRjKCKHOeLzzvY8py
dKCjT+KVjo4txvQGLX7UIgxBDScPVwGMjslocGOsYaJ7xl2XN/PKMyCiLJpzVtbi
9U+h4PmMnJt5Z6mwZRx5LX6seHMfQkC3EDyKQnNNjn3Zg4MxtfumV7qBEv1FoQa2
+FgdEgSDIlBg5Dy1mQcSn2ndUUUaH4FhuUC5DwyA4ZiDNQ/TrW/IZy51cbE3VaSH
3KPO6JQV3HQDmlPaJK9J+31kiQnnXq44DhqfbGVZ4O+gu49M1Ir3GgUbNmir3lHc
yVDGODBtyCPBCw2VmVaDsvBoX8kbBHVBlJBBEfx+0RNHfNkxDaaAisMLEbr9+Erv
+kRJ0P2ra5XlcnmyQJWGVlFJ+FtHEa4U5hqw2436Qp+rdqeFErIytjf9Jo2kp9Td
0eg5RThrMWBuA4AgaHLQVx2XFBGJUe/MtmjEi0yCGeyOsVUiaJwlNZ2dCcDh1jZ3
dSG+X5UuWMpypa8KmpY2ubLUutrQzckg/9SaZskC+dQXxWe2xPwrHliqhuJgS+Pc
UPA+/3OLfoNtV/U8XFT4dngvE6yxnXbSqEUNW7Iu3a5KQwS/J13eRycHIghsb3mz
/wRRzcP0GjeSNUfFwS2jiuQRrbuV+p/PjQnQIEjbKNU3yplmuHadY2Us4YFKNnjt
MfLqGTqVLyoFHPrU7KDcFB8aRn0z+t0S7zJ/lm3oU2cdHJiVJebxn9Y67UGvem9G
0BPwmSuuIwJ/Ofn3jOmUu7G9g0ImznySbF9EWOZq6iw6Vu7pGleM2iZVL2iC4tJX
CAMY0H6HOBVr9bwYRAlzf1HgcgpvoHFAGC7V8KnnVunEj4Y8WM3PTCRJ6aI3LITJ
fTGXUrK17vQ4I9JwVsZRuLOiQRrYnZYbkZbHEsGJFTdEJ15KWpqUrRZqPHiSuRMd
3bW7V6DIXHpjAB5HXFwqeIqb05B23YIDFw1KRh6twHBCMFL9kqPkVd00KmAAiXMJ
2PVJasg3ugR7bga1g2CSPxQ1eu8FfR8Kg1hhu1mFt6Lmsv1OJWgcCSi2AQPrl2oD
5CCrvBn8uhU0RVyqv8BBewy3XPOxpV7qTUhiM0ShJ4tqlYxj4ion4h07Y5uZZSD0
PscyOBTD4NPjTI2jq76tat2vfPPDUD739XhiZvHMizunBoB4VMzcu8tfqcuWW7gL
GyvlWnfIqRMXCMxZpeIDvHMSMpSXUAmOy4dbv3yt4gBwViJTA16Tk2W6v6tfl1Ex
6N83y39vAPssvs6KuXOi+Pp/xEr0jSpCnQdQW6Da7XJPSiSPDGluSMHStmzB95+A
9rkPf4e7FpJCwH7bNoIueVAViBXYfNcTZ7h6qQpW6iri8wISeR8vnV7A4GJtDkjh
yLQTzdBnUGH5V9rMdJjGIYPPvjYVzgrx+xZt7efgnbcXwJzaPBlWlgiFb+S30sbT
G62YDeLDfrmql5omPrOTuMvw8LDiALvqeZhbh+RIs0zpShovHqsmMiiQWehdnrWa
TCCDmjMtzP9U/6EPfAOFyb/p/ghlhjwJ2i66ZkatGjs6nQmYdhneMchJ7ABrPt7i
hg4MXnp9EZz43v7Kl/0z7qxE/kmNOWSYgGAKM9H2dMTHFzTqPMwrj4OpsHNG/TC+
m/PARB9ZGZ/6ozpGtcb4V1l5GXVdmrG7NmvWoE3Q78g4mynIRV5CM5bMye0I5PMd
fQOQt+rdgZFPqkvSuDvjboRxXuL3UXpjSnwpoSyC1XTAsBZgmeOxZC+EPn+Iw3Jg
kk75boNZulWftGN5XUWu0CqHCL1K9+PaP1mh3qdw6nnjpMF3tEUssFdp9Kg4/KO8
p6wUWuPIO/58f7A6gb/j5ngbSMPrXFkeiPZbzKiRNrWMaZEOkN50CK2TQFysrS7t
fIMQ0eOqEYaYFX6p4QXJlCuDAScp0KypD6Ia/ep7oz85ihrI609fu0nGtaRyWKxJ
6yNue7sRcoCLZNlzoqQd/QNH5pDfDf45YnmzgbB+Q1aLHveyl4+/UKn6z48Y287F
Ai8vtCKlLaTzwyqWqDA5fRI5tStuzRF6O+dgd0BilV1saOvSxlldLsXH5Enp0Kro
p/PrIuQRY2g8ujoRRjLupE7YeUxCLVMjL2m0sQ2eipAAR7y0enAQ2I0I2rqmUMnh
VLpXVlwHo/RaeQlFELfsEtw1lWTs9yGcDP3Md4+mqLds1K+JVbdYuYTBiXdJR7Ri
RMklD8tPFmvFVpFbdDynZU8MO9yEU2uQxLXvnoOJswS8FzPI7oPchdc5ib1dcbuq
QGL2tIf4ey7NXxSH57Sfl1AAhTFi/3s4rxY3l51/9jiWyYznFMhVmz9skZM4UYXd
Bl9OyqRWFqtfy5RhhJijjcGHi/RVhOe+ZiOQ5IQhCXHJzj5W//+yBOtuIxERqlni
5VCfJ4jOq65CPCy1zxIc1/tSmX8r7R8lEe66EHZFn0O6QxBkIRoqjRjJTzLdQQzg
25Wxc+Zw2UcLhTGL9UXs3TCJldyUjSl/ZwVT6F3o91sSl43WIzvHI7nghr8h0adW
eoesTD3z+oSqZ0vcBMWqqhQGf/VQY6A2IMU/qWnov+CSEpBKkCha+BX2BBHFRwAE
bj4erhckD0KoJw8soutg7T60zacanh/i9LvBFc8ppXAGQGMxwRIzxbQ4cK3HwKGG
yaXlRKFmb4LvCk81Z48kuz4xmSEL3lTqVOK//DSmCksPsWmu25ujR+syasO7umVG
fiCbHtLmrHSv6PPweiSpr/l7LssyggzrUkKQoI7wDwyfRTZ4/JqiBtX67BrBLUr4
+Z8zDkb5Fn8jifpwy4hYJJFnve0U73GHwCOC0/vRtM0eX5Gb43biujvegH6phWmY
nM4wOR6mz502+6ycyKBbjmecGKaRl+5GC8aFcV6qvKAXpqd8VMZHkDciR6RrkYIp
JWHgxk2uS5l9+zDfBIFOj63LZsBWDHkii1R2hYlBQRBDVZmNrkaxTACn3BKfMaKz
PnItsTCk4QQuS5zdsa8HiGq/lyOJxG1FZd7BYVyyAjGvATDmHgrNZ6bSi8IMBncO
4zK1SmB+DZEa8NB6DKZBBrcy09+SAfyVIKjzJY1v7djjKT+GIHME13DtZ6Zj3uC9
L8eww26zdxRI/C4jAelA8AZslTRgfdWgraeyq3bTidlXCmrjz9pbVMbReF54ortV
D+nGFya9i5lrh/qWa4UHrHwXaAs2XUSPlK6VeguJm481C2MPm4ymNl6DPYu6GIdf
niyUlibVxzaOBa5/kgJm2y1RfUxBSUY0AIhgP5mXdzoJAz4nYHMOs01J19ZvgWhj
Ft5AgFmWb2f/fQIzwh+qcRIxzouugKFnCOcCUSXVn7EhLdJGhs9P+FFfpTAS7AZn
A1tBYj5lsH/XpBt6IaA7H0jL5X/54QQENLK1iNSsYLigJK/WFti6IweVBecLDZpJ
+5XwVHQJxtvVpLiuWBYRcIqBaZdDgNxgdZMQxluhhmsz87mRClayiYReQvqebai2
r9qUd6IbznmgaVmnU2t94CxVlmMaqds7WX/NffHQ3aeoz3q1nEyqOZAZqNfBDF6R
iclTpGowj65pLwByCXicwC0bEjtpHCXwqxDnG5JhESeaHxCZ2kIaJ8yrlxaP0Hr0
jf+haSplD4Y4Gb2XCjnMLBPUCrUrjmfM4U/IGwhuu6mFcWnJldOX0POSO3ndVVe/
GBtTxsH1+5pokolw/bKk1vaTOCWF1T+51ZoLCgVYApRYcGpS0rZS3wiHkrec7N9e
NUvjN7v7Kj93fH/Zj64kRiuh5vtZ83DePO13I6ldoxCiy+x2Bf+wonZgU9u+jjHf
/3KIR00a65Fj+tUn6PQHe9pPvnfFbDQwoK+VL6JGbfMQrC/uW40rLZKSxcY0dEUG
amJqP3TpDsYeBFQHz8c+w6aVxK6BztA3opw4wphRum9vBqWWQ3dkpS5lTcwJnW5A
79SAU9iADxq/g5WJCoNwjID/r+Uxiat3BS0tEvVP5IdEHkxcX1RNwKQJQnR7DqUo
Lnwc4le28SrRSF+372LwdCwXjftg2Yj652dhl4+CEulwMls2+bCupHF63bCloKRD
HH6IsbgJiDFBbdH9NNpsokkXbI732QGiAQgAYt2p3Vu78C/srr15KTGXBxWdeqXL
va3MXcKXAP2qsPvgjvpOfR2LC12fZ3V8vXnQwP+7KhZg1nNyQNzYz2HE0Oeew5zs
gBCFoTZtWqwAPakx7b5MC+byJYlUEHZ0wLItYD/AtJFs9h1mgvUp2D+tZc86duDR
S5OI8iH1M69GrYv14k/126qplluUvkJT+v6YY1BxjX6aKXxlmguqAFkygwSHFLu+
fTS09ugBTSjUarmJffFNYBe68sr6QlY+TNzunP6k6xr4ca8kRKm6b1OWi+RnIBnQ
Fs09eBSLqGNKEQ3JQiVN8/rhOCR0oFAp/CoVxtESt5UmqHFEwhfPq1cWnYuBbBjg
NyAPiBW+WO3ha7BSXON0omUsl08OyIvPk9TLjP9KIwTfun12itnlTinfkkxonFLB
YV68M/6SvVhJZfIgr/8hyYXaUfPMZTD2b1ncwqN0kh/TwndLnoe5KPpQ4C9wQ5e+
XzGoE2UNKKF8TfPMa1R0Vw==
`protect end_protected