`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13312 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
r0poS0ytQydMvF+aKdd0eIq0dE1ZoL7GFS2eJvDsjY6lSutdzHMXBm8qwnr6AHsU
QGJsAcjD4ld7pS+VT4NbDfIBeGjeQ6mMKYgzc5hYlNpP/CXTFU0OwDVMr+2ZDJQ0
maY5FMozdkw6puUCf+p/rw185uCydNclac/oBCLCfQot80NRri3KgQI8R0Eu4BId
fK6EeRlKIziBVc8VfHV7/HGB3NrOJbbB3OILJJAwLQwPVxKwk09E9Dq6a04oAIw1
UjrqMZpTTfkPeK00qxh4KsMr6/0cDkcAUg6cLZV+X2V0ZVCfsVYHOnNbpor6tl+2
PrACzS6zDX5fRQyN1kab4zXIidXhY+i5rpTLM39O1kT2nQczyx1UcorAbjdw257/
ju/3wECzXOY9/usH5EGZvZzka91TBfV1jshz38E+Ni8XEdgP/J6lGn7nW/B+zQkC
DPKEPGqD62bt7E5d/+q64u9N7Y5RVGcat6eHw8YzekRvPa4C7si+V88G1u4KKHg9
nSk4GxoV/cjrel61OPRNZvH4JRP9ql066Hn5vOCmsNNTCY/MX9PfLP2VcFv+nzWw
ChRYjziENwv4Z1pZmndWliYAOFyyJekfZHrxbPqs6GBwDHCn4X+VIsBvLdgTnzbv
qXeqvE8ZPkbjNgmR4N20aOkTxdJEyDxn22DuifqWa1lx5IlcVQ0VT9Qk5cXW10L4
paS2CNja7EDSUrw2UkjOjDKl63jYwyRuKYecvh2Z8jNcNKS+/CpU65XMyyFkZP5B
bqHxhjoX5kjm4BP/sLrED86W0xS1oqxZ1RXduxFEbhQsH+4oP7BHDJmdkWz/kGdX
0ZDo6ZnRysfFMlrSPkQlX+ofexzsHBgJN7dc1MCw1pWzXTCDukVzhkmpiN3PV9JB
GYYmjF1iPvpSgXzlyE7RHwHD2/jYYPKtYsN/af+UnMDa6Cs1D51EXaw2XP5GlQHI
Ml/VpQ2P5cYkCGFil75ObOTHHl3blzMwtYiYXsLujhu/X3RMxVb3FvXnLefFuIZK
8dczM8ZCvxXSvkYN/mz35WmTQFmci4OOWVGipWmAeyOknFZocCRVjaAMSIsQJdlm
7h07om3mXTe/oSzjz0gjraOBgqX2MOgmm8vfsJnt7SIsjZC1oDYmtLlDhGJLujXD
KH8djRfIw6AcCK2pd9iWylVH0ICNPgUxnAyGSsfyIswDh9/EqmaEBLsVu3FoxaGL
A9/1VnPGgE1BY8SpjIV6MlwmInkI+aqV7MVSQHr/dpQRXr8fCuCJJ/x5y3Msg7pF
4A10eu6IpTmvGlHYYx1O1FStkbGrdvYCUvcJYez8LnXuW5QHzslU+nMtEzfeRu57
NF5zwT/N0gBQ9d7nfehdJK4zLABN7OY3kK+VAguo/47Z9n1wKVPyRRgIsY3tlM8C
V/4A9x80NSo6g1ZocFwnMwLl5/AnD0Ylbl2bPD6xLQ1OLh76Ce5rY7RemgKP4PI/
snWPMAxaDNgF4UvrjbQxMG0UAzkJ/F/7KlrGExHjiKz/eO42eB1Rpq0vQ9axcMSV
JFeB9cI6s947d7Mzr6Sj15SKhAfWuI+z0dU8J8RCY9rE7foahzU5uEqwJ0JbA4wN
UU/ovj0s/IM6hvbe9TWGgIGs1GjX2aUT1x/cbivENgKqX56tfypZnY2cr4aiBWJQ
phAX6PCb7fn3Ikp3V/vs/mmzRRJru96esTH0axfhrdqYGly1q1e1Crasa23GJKcI
j6/+OKMlhFaF4uTI4A3gvfDEhi+7eT3uw+3P3pc/CNwaa96IqjjrAjgy4Cq/ummr
nCadFPFn8oFqMQq7Ul1YPVN/QUb5i30FodJrhi9pUVaGhn+w/z+eskiobrjg2i8U
96gXIK+OzwlU1b5vCGGQxMMOEiG2+7Rr0kejA71xWl1Nweu2kyhGiS+P22lFY6bD
4PglXEi/rjOQ5m9Q9VoKlTpOXUbDO8MFHPgJVZAEIGTuPxZVg4z1hPVnklQXPbTX
duZbu0nNKhl+j2AmEss2QAu3UzIvCDdMTO8YpMiYhBAVfjHCXIuHpQiZKgm+M0BY
BzMVA5wwf1P77NykR45KfDnY8cWcZz2+4ztnSTLMIOUkzIqbShA0pt63oxuPKE/E
XuY1nFHywVOAEwGcG9cTW+y430xkboxMta5qhKHk0KijxA6lNbxBgKNIyGbgp3JY
BHgz99yMdqIZxPCEU0NvlPh0rf/ydgHC/a1GvujUXMDg2lghbhfOvrT1Idl3nFaf
lu2lsyfvU8bTMZnX+6LRHU3h7fAXLiVcWE33M75DxvMUQ1NXyZ+JZfN+DxSyrXnL
rVcqWIZLog6RMqGDXGDdYZ862gC08SxY57i//B5bPijKAu31LB5vSk24Ykpkqk1s
m5yExzR+2HGfu7ORkrJaZT/JKJ7SsngwOwcEcGl8aYkrWEt/h1P5CHVB1zRfMvvi
83xvYxF7aDEXzYh70KOV2qCSBlKq8Evde8Jfk8miDajlsIE4ItjhVjAB8P/KyX0D
GhuSEEx4s9hF90x6AbAqvKThxNyA/C03NNGk5fevqRK7iYyA9CLVptYqwAhdvxhR
rm+IvEWkgBELwsI5i34U+Nu7KPgVkxjuFBeFS9lPN0re+4P02gxk2HahtPJeC9cI
fOGrMYt6AjtPjXkqti0FiUkxUBHIDSZmjlmLBlkgBp5A6rsWtbkabPDFiKrIRldM
iDKI5eUsf6yaWYLyieY+GMINO2cEP3kLR4P1c+s0sZJY0d5hW53ETobyUIXtFOfj
bgyMwiM3/8yZZaFkmulxbk/kvv21o/5WnVCWcpSoKmM3o4NRCH7w5Pt0GuNCFryP
+ggtvS3FJGRno/ndGfWe2EyuO1rJAcnB8cgptfR87FAvN8b8mlpL5xIyHEieM7cT
20YOJ9JQdzMdBEKP7R6Undwzrj7DiTJ4N276J/4dttAfFQgAvUlYMGR7VPYh6pJy
4xFEVf0MPcjNT03CCCZ7q0z8+Lsxx0e2OzOS+rvTCoqXvytsEhZo8lC+YE+2xOKF
m3a6cPUFsLPGuK1ycwblBPE6BLPKqxKlXsuhgEWNYUenAS+Wb/ea+80PJ+miSPbv
d4QplnBnKLwcUJzBqiXwHllgZHKPjkgq+dgY9bCJDqrhnZCprhw4ztmVzNM4aMgQ
/M+3HBEyU714kIg/FObeEjASMzcGsplwxIMqnOAdh3MO4pbtfpm9E39Hz47Vcjt4
aTHs6kyyyNFLbfEJgUO7GYHup3rwEp51+XO1xCJnJ0s6Nvy9tqrflGz6/a7CncVn
Sh4RyROpR06Pf6WI4ZPg3IDKsH6LfJK9QDDlFSqIBilp9cgq2nprPlvTY3qhLLk5
N4peVXfT4lC5snNuMBR2OHZ/dMyJBswV3KqxJTLGaRlsy72p3kMRlCTQaLFoT8O8
8Jo2VwIYJMobTzpdzVlq5KXIu0OLJJ5/fmfC9fQsgwc2LPdEOcDTm+SwdfIaIkxI
C/DFdmpgs8Asu46VbgJhXfaGt3YTKWE3LNjmWpsXQP0yx5ZWWPdrP9GvOo6v6OuH
xRHeriWA8wR11O/F8MTv+1dRDmZyeZSneazW1yal/RdypEt/5u2KV5zuDQI5kjMC
FMHhqqU4VQrp8MebY7HejdTXrbEKfMufms9mAOUrhvxT3CkydFFA94r285xLgWFP
9aLSCuvDvgvSiYcGtpXcg01Z04ZPHr0ZYp/ozRrsYNz1VGiEVb5KK89MA4m0j+3v
sZ17u7iPFKGkPRdTm9m+Jucycif3o2pQJGRDaZEE+IFz5HzHCuM8FXtaTgk+rVOq
mangSBcF2QcOuyrmPP6O6AFwhLSw6BnyDkseYEP9LYbUuSbyfPFNIpvoigMDxrOO
izOkVmAX0oWOqyu6VW+l8nZzXRQ2WX2ogC4iLOauAJxP6bq4IZ4hUlckjj2R1UKS
cGHJ7tA1g0Q3UNLQjCYwLGum2nOVwCLuhksvNW4lpq1DSN8jG1wVi0NjKp6mQOFb
SC8NsTfmz4B85Ti5/Q8LmI95x9/cj1d+/LJLE5Vux1XQXMVeFAg+QcDrppPelv/b
0tArd3jNmXaP0duIo6uzwvMPK+twWHlNP/e//bMxHRuLKhJuArMgi0EGUeFYoFYs
vNc/f0GuC5dRDx9hsJVxFFARE4yytECmREw1eK5xHKK5arRbX0+m1cLXnDLp+rCq
rzwrCLr+ZZ2azDVzb+O84wJAWdjPy1tkGEL8FkrtOxc9R2l+9D8Lu8LQPNXtfrYv
7B+sQ0PmvdcQeVcVIEhyCYHKhvxEqFdapTGzOzY2KV3Ztt3vm/bjbGTOot1GEAlq
oeSPAGexFNb9f9YMWuzfZQh2p7YrDIntD3P3dCskgb6sBwpbuoML/Fw+zItFb51v
J6Cqns6qxPGtxUMcywYYjPWKtA9uZuxcA0UjFOjXYq95Zd1s9kPuNx7anXyZyl6m
x0KLT4veqrI2mwywRihT+heK4kvTFH+hhF2uL3t8+pL76tdnz1O5+VJUmfItDRDN
p6QtxT3hPlYYIY4vNhp7NBF8Z4vkuCRQ4lnaB/M0dbUzML/ktOJmy9yiKBZ2bv5F
oOKofS9jXRjSiqNa92x6kpyQjnN74rxRuKJ70owIelzIVLGDdclAOsjIXWubU0Tw
eAjVvkPJBeeDhJe6ETvlsoShvedfc9Do+SYPj4f/dVPsyhIYHskMLVHpWhGjwNCx
C9vyortpYkYihu+78gjhTe/u3LX4JjaU+7FnUhpKzgtlILOzLmcNLbh6YR6ePhcN
eGc6UEnezuxNb74vN/ATeBajdFF5nHdPInLRV4d0Ji17f8FS5BQaRUNRyQsqVaS2
hzeNx7/GO1UEcE0hAvR5Woj8atbI8gyGqLPiiptquhmSM/Eninrn9rneXsYRs4tY
SCdLoQg/dFuJj0Ad5RPRBPzvTsBdcS8AMRe7hrQXDmfgNQ0p3yPgyV+zZoWMqQOV
7wtNb4DX+mOkVzs8r7apN8+SANWlfP1dgpjGQwX0gRwwStdAbelPZCYuM2X9yQQ7
2KRo6SmSiHXPPcZtAG2UMLb5xNmnKHEJbS/DZ4NXzQQ/CEI5a3sYdWdzVdcBzRHo
P2/79q94Yk4ty4wpCAVA2HaXKjxB7zxjcXqdcXnh5II2cwQE5tJOJrobWPa/mffj
SWkBF1dgiCmY4roRxvwqvMw40x4rVKYKTwilwMslJ112zzXfL+g6doECEQGU8mHJ
C/tHOwh3NurEeAjuNeXUyKIGSoWhRHhPAOSot/kWpILSuiEMbE0hkb47q59Y+kxO
ruXDGC2kmrRrJzIdZdbZ2q0j6J33LpB6ReW5Km2RlLK5396EhPjqjA3GBd81aLWS
GUWAEehpizyNXr6HE3Muwx9jwNoJ5F0GZm1FxAfaimP1tg456TnOJnBty0Te22yQ
w4pGj8oDuiaTsRe6kj0b85tuM739JF+lpYB7oHMmxYIZWvvlOgGHdNueEEKFRmG7
cFl4QE8JRVzqg36aLKYr4SHtLmfkGeGfWMR01EnuddvVA7aYAKU1xKlnECkW/gDg
hFbGPDr1tX/TXp45j7pe0pezONQzOFtbU3IOg2XSDePMdVD3/p/ACy2BGTSM4IRV
s7sdC1wbe6TyGRZia7W6R14aDwpFMSdCKNRwpHvrsE2UW/qsLRfAseCYrKFToDnf
Kq0sbKYRVeV+Zrk0GvPTo/2QnQOSPsiUUvJJHrzF1QBC00bi/x1zjWEIVz/vmn7x
yCnvQlKgX/OpfmLmgBI4WvQeay+twJWjO+r4oD/WCF7w8kSBsLAwqg2y3oATnqzE
+oSf1ftZlWLE1cvox3XWGxkQkZIrcf6RSb3Q9eU/z8uCFSitasOhgNfledYQaaQI
0bmXlawwF1G7KIF7Oc7Q7h0ZC1HOkgEqEqvrW22w+hmJAlfwbAL9anVuepVR8GWY
HVGl3bzE+sOhNkY18xY553JwzvB8bc4BQFeLc1OUzbi4KWfSM6xOm7ZDKF6zK8ZP
R3Y0jDpmF0LyXvLnOw+n3wqWYI7qbezI/ECD5ZirwyftUW6NEnphV2AJy4FeQB2Z
A6fS9P6EzM5++tZa9rt49XmBwXCA2Dnfnsq53DkkRkxffGQTCNGrXA8O9knpyChS
ptySUZKj0xIc428KaGOr78E7+eKK4H+R9pGKItQdb/G/O+BLkv9K6tjT/uF+cmCB
WAvpEQoO7q54we5hmDu5luRKd5p5xyGo5P6xrHigAuEQsk7g2J+AUmJGxZThTnzS
ikbcTOUGvOr50TLeqK7qBAUeaiU5C02k/EP7GuNGi9EQ7f7uKkYj0UFEdwODNckQ
cB3gASVMlrrNsLVKOiyjc164N80hutUQuXPFfFfhpczeL3d1zRxtQBHFRUwitIPT
GorXmNOu8bn9u/UasbysjtyAt9CRp+4tfwqCeVqVWX67pdc/bqgufFLGw90tFqOm
QpgJcrHvczBlPwR8BuhYkOOCU8/Rtk8lrF9+uu8ToEWY4tKNYoW3kQx0ZO7ZNVKZ
rFnePqHe8kceMtn32Iti0X2XrkThCFYKzC9JpjZS4s3nXTfeiOYbsTYeBlSLRgVK
nVJE+aKIahuVAHYBVIC4L5tyy55gssMp6s9RHfHYNJTK44S0s+a1TAzk7bfrSaqf
+lWTlZorcFXcSGfB4qEMy2KusdM5iOEwL3U+PzODdT5hxAakuiT+SPXAf9UE8cum
+Jn7vlxIss6KX27S0Bc9/yqgQSAjgRDKXuOIPLNmI6bTifExoPZ8q2a5YafdWgn5
HVmCJZZIqcs8SWtY7ZFBgHRuQOOcoaC9/VOTFtMrxTbvS8ZIpGQMD2QMJE6i3J25
pFY3D7lm7N25Wwa5v14XTWAZZ0lHobYGct+emTp96Vdw+XXRRhT/NM6PYBaSZBTB
5d/3QJqmxE/BocoT5KobhvYrG/Bx0uJqh7JBLd8E25G62gj12RVSUYEFyJDL1THO
v+Ao6qhahR0nBd6nd1ODfG4AvSdtOiEyvPsYmQeWpBDrsh6K5TqD8j7cHlPBZteG
QKMeiPCvhDCzi/nxlTcnuDQJUvSU+YEloCahm/g0iyvtC0LSFjXr0o0IrXwmLrnG
Is0VHHYBWQKLsqbJhZ/jYX0zf+aMKHudww31o4+3D36DI2FmYfRwiFuzrofRX0OZ
rDDtGO0Y6iWLH39kK4Cop58LUV+OsGThP3QBx7f6tfY8U4b0jChoqrVa2J8O32+p
cB5vesUDT3dUQQhCbDQBHQGW3zlHRtM8p7VnPjjxNO3pF9dl/087vu0lixxwrmRJ
xMz1kkwxbEukyEfK++SyASj2K8pylx8GzLREjLl68eFR+gQKTfoJrjenDePxVXc6
c817iw/+asAlaBNYdjZk2o1kLgjwAp8HGRMN8z+6cEfz2f38ToWjA0MU3q35qTuF
hFQd3z/sOpRSMCi3x2Ba2zhnQKO2n0zWiOjU0cIluXm+LTVXcxDzV2TbnOWP2xVu
54k/i6g/dgkTXrPJttK/mx6fxTtnsWFnCfW8nslpLTA6VS28TZ2jS/5+i1U7p5AK
TaajHOpiH7dlzQop9zKbQsbEeLy/pu6u6vAtJEPG5uhH2XKD4NePLNnMBkSWQmeW
VStCjXhCiuXpThntF4LNrgbK6cEkbaDlr509iVMOFOm9CmnAeBjpWbewJ95wyesM
nFtK3B22u2TKkCkKUdGrQUDGNS2aqCAXUPjfjpqP8xLwlD+yBWl24B/TcOmyr2oK
XZPVGI0is+pYRuMIE8vGSYRjCLItdEqhqwleJQNOT0d0PYSfjssMvcRAKtE53XQ8
pRVVAnw1kwuB8BP1AAQmb5QjfDox6uPx3BktyEdXllWXNYbIopAS0jCpQ0te+HXG
5T5a82vBnfcLHu4ZMqquDEhVDmYF7Ja+Uh00q6y27WUOefvSuQ2VDfmQpJrB380F
CtboRkbnVsDvhBQ3wyqMWrbSYAX542UN+RGYasykfRBiIiUAwH9HKcFxlMPRbGXs
i8k3gie1PGK6AEEqSjvYywUwBUOlo/CZ7291LVuXhDGhAYSO9Np5jpueATH7O2Xd
/6nek2fSzjlFf4/oeapZpplhwiZTcoanyvXdjLCl4IPTOSW4A5HtTa/WnvDmMyph
tKYmBvIZcaGxd/Yl8eOVl3ugABMfpxiuEXpr1J+IK67IPBG/FlMS+bgb9vYSPBx4
b9j9ajd5pPdFGFbMdAM2xakCuppqxOd5fN3SbfcvREyykLFNUhUxN12/D65WJ8kr
zgcjNGYA7NXYPS+TiDZjrPguo/KYSkTGbECGFFX6or8SPBDrtmeHiRsNkpk16JDt
rsX7NAx8TN0d91y2jSPKQPd3Pryo/ffevrkDGeMFAHA5DlvKv8tus16YfDxfMHE8
U84LJFuJ83/aMLe0BoPBRW02sEMRq+8iszSiTccdzwQ9SmHT1IT2wbqP0saRTbCm
PNrdPd19+BPD+B0x/FcjlmVdBwKCbZ0xDt/oW2R88t+aefdgcdtlSobz6hccMRRT
dN2L5Xpgp7oFRQh67DRqXH3ejH3WLGIFu9LUrAA1HvaFrzqB+ab05MTROOMVEhdN
sd+4xwTy54Wmt2oU+8yvXje5vLaCIWcCupuFFJHiqFEf+ppNz2RwKmfTxe6cB82S
0Ug5C1r9hhgNMZOuSBcmUQxuXs/bJnlacQx5IOkJNQdwuSQdOkwWVQt/bYNpqitq
UpZjoMpZZ/wjuytNHJOHGyVdcsKAdWctEHXfZKQQ4XgQw1nzV/c7F+YtleB8phVE
aTETpA2t7LJ+QUIul/qvMk2xpaABmayCmbYzzBC6d+yCLYdF3yMgIxtP5vs8Y4pl
Wz3b2mgscCV3LXI7Ra34o76icLh1t4xuEzBScqaYN5zuwC2CgMxeSTZ1kE/eFscN
LvQynu9fp416CHRKlNXlK4WMFyObjumj3p2ZmM8ZLvEyLaDxRa2yQLQmBE4r7LFl
JPdWqxEddauCyvdrmph0MwiukakAlga66qB634g71bVjZar9N4ynDr/nnqE2Cp0Z
OC8bf3wnmcN+hh1Cf4dHzaL2/LaPwS6kI3XZ5WlLYx5eiKu0PAA3XeFb4zR+WDsi
uHYTjm24/EIKeI+1v20q4gXI9HdEGFP+ul1UjFRbJARPsyuqwz6SG3UGKcMM8WOe
+PoHzfNqfRuK4QomQ7dOS2BE7n+n1wdQFqTxLiHTGXZe0d70TWKGTcZvbcM+olYS
MhBbxNaLFVPYd9EVzlFV7GBRPEeEBz4O+Cx2cytPwMsy1q8iWojxXlvPdarUdQ3B
1mfTCPksc6uBnoZJ0WO4vXrrWmUTLVn+Czx7a9AXZBaVPURdFjFxjCdfK2k+SY8q
26p1Xqug0RS12GGJ7XPGW1CAhvQIxnk/5sX7T+9cI+QuYidqZxWdccgSoe7uB6UD
WarU//w/KEGhVbRUHHmCe8BFkF0+qCcoP2PMg3vXBhbfhJK1HW4tQK9B3t4htWNZ
ICUPDTH+sv6HpfNOg19X0DFpDr+usZMaXwatTcpYoHQTMBKrxw/HFHwMJbFrifbo
Krh+n9VQiGTZb8IewuOM1FD6nscOJkLUc1ABDKb0ZZs/UUQQ97lwMvE2vTesOeuq
ZsBx1RlL2bUc5wxgYn3i4hX1ZsW/Gn3vhttUpwbHcELkfP7karAfc+i11T+zKPDd
QZPhzYLpneA4znH11lQcj+7pBRk9oyQrIlKISedFieLuxn+HDF8xzlWT6knMGdiZ
09W1txRC4hYrTCWESFmNRQDxWYcT3Atu5vFhmMzX6xusERs4Do+BgWKnVrlD75mg
GvYsX1hAPM/hl0kQn9q05oiPS/1VJNYeVGl10eMYQfIsDwc9SPOHQqIhm+y5524/
1HC3alU03GqPRr6mxL4copTOkMB8TjiJjq4SE26BZKMB9tVfAgVG2pziH0nhUvr3
0ecPV6f4dFsjglDxlNkdI4jmSWeRNg15iAF4Bz7rqDLt4U0y23xkx/vmngOM5bk6
kvLiZMFJN1hBhJcFz6yzr7S0WGufRc28kpaXyiXjzzPCsCfKJZX/Kg8OijuYuHUh
o5uZV2cIBZe8xaDnBy4kXCc3H6Qhx2styLrCUGrGa7I6MtsvkECvlSIPnzd/6l88
X86ld8D6sLV2AfdsjP6U6iu4jPMMwIrfbYBzDZBJAm/0hDCyO2YYIGsWy/QF321T
7coyOHR6EXbEX4fHEp8eppoDe4atQphMJk0Lv5as559ERKGtEqiNutX2SZC9Xm7g
KK/71VdIsmg5+EBqRT7LFd4qhp3yAbPUY/+x00FY5CqgfH+oUTJ0zM9/IwLHtHdj
Bj4pA+q80VWGVy+9ThdWH1VgXBMG9EVQG72rKNwvcnTI3GtF+xh0xWveI8kLWvzX
4+vU8gVqeQSEWSa8eA+NbUh/4Xk+wwy/lQbzUMwg59c6mhvUq3jUGrxcVM2ykvDd
DZFHZ43J+Ufjc4L0hxFG9lK0xRdqRNPPRTLKFNdt75bwGvwMON8P4v1g3pKUHSEv
wMT1abiyxtsGHRabcolNY+AYsZlvoNkek39sQRlNrZv3lPkjotRMgs/ZdKWlYdyW
iDXMHhZDjjsNMzNOk/YR8RBzHG59vnr52wztslNmFJO7MWkYeO36L9ZcKoybi1NR
CQzxV6CbDHxGKE2ERtXwMhTmz3DcfNIfzpRyzMi5AaxGMOW16bS18ycTR+1KUYPe
P2gLgd9mWuPtQpxHuYSw/Wz1NxwWsnAF5oMWRGjVJdiCc0zR2+LU35gwLJYx8xgT
clSqkH5fnJHu/EkQDyi9XDdvSAQ45YeQY++6RWbr0C7SPLSbyFxygIxySgOvBTCB
z3+NbyqRi5xZjxuLS9gTQE1KH2cZINupBDELqVzbtEnOHgXmZ952OXjORyRlTkOo
sP52nmXQMK3NdgZfCYWg5AljkQG8g41cNBCCSTva5XLgPVFr6R7YO97zl4b3MInq
WxyhuA2l0mEnmQm2LoUanTwJAxSZNGfnagyFK7gijVEzoP56osOUF/kof1wVET7O
ZWpI70ESztx0ndRTA1kucyjPH1OQFjSi0jBtZmli3FyKhTPR32m3NncStnocsDkO
ys2N7cYn9+35Qx89JBs/Km6ham8By+jZ2h0VHsIgPVJ0RJw4KFtemhTDP/WTwAu9
y6Iet9GB//zHBVu8qmc3rn6WM1VrPPlNqt3jKwYQK5nh6ZCCB1rK4ZTVEfE2OFVY
y6O8MF8382ugpXWZGuSOZVYec7Z2KuUtLUYiq88UXBoQqHyHYLT8fAKpTDYDaGMn
xdEVizVLN964HSmmJpC548dxAtOaTpphWDhbI66LJmhfF2kbI3cUi8gFaAfXE/yl
ZpFIgYKrthrYSc9Dve/eOWz+oOWIwRY25gSPgroexm5nkNP34BSjrw38Q4cYkW/+
oneDRI3WIT3bvwohT50KW3jXp+iBd9Frvt6ai2IgxpkX0ixfE32g+ZCMysi7B/8E
8Dstmcw8qW7dyJiXGI1SIDxUCcDTG/7gRVaS3sOTjZlramaEjgUXljhGUMMT73v5
xM85DYKYyl2/lzqc56y3Q4a4XYsODUEMrxA4/GJ5JM8AyBPP+19X4lqPP8Bs6Sir
JWgAydJDXiWOPpL6fHAnLSkFEyZbhpXNAh/+n+nB6liKCbMFgMHK7XGwIjMSvLel
Gmp8kRfnzIl1k1ViT1wS2p4wHJZGA51HFaOipD4X7MVipDi0EdihzJ1ek1OcYdrP
xWi/tb6uEHiZLkKXpgTwNAmx9ZPmR9gSKo2VIJiFnBi7+yHdy1+u9SAyUhuPJPQZ
0mvN54lRcjf/rtDAZKk2uEhNFv5u5Bshe2lE6HnPDgEidTGERjgKoscXVKGYB4+V
tE+zJ8HIiQsokWicED92zbSWFI6vSYmgzR25qDExnEuhzxCcgcANsSCVeUQCSF4J
rYKzt0dU5A9+D4TZWampIhkrhCxdznO7dASCbheqyFaN7UjJM90ZyuuvSuAJLIhy
nc6Wn8joiMyBUS5LI8JOem2CqmitHztOX0e/XDKYjyblwxezACWKkxuXYf+woXCR
/nnLj8a+KfHj+SR6TLaAaUBk7YVqNgAjvAd5ye5d2c9sUFGj7UzyKrIMw0pux579
vwnHbiuF9Mm9ItIXsVVnMultTOe+t+RPiaZE0Rz878qlyVZCCzPC73UfOnm2Slxt
6NdoVhua0OoGevtTHUJV/bANJd9UkdIzfllmbepyvPPdrjosJbLHRtetqGIUTG/+
ZPZPNSiFm66dQThXYODMz0GHo+7VHFEgQ3vgQ8E4/eV1Ht7xOSoYnGDdJ3d+LAYm
6EVhi+5gMsJ+NSag9dTMfrV8FslqjZFLiDJg88H2KO+SW7c/17KcZI/W5xABZHeQ
olTWRUFe3Df4rqCW8oYANjgyAwJLIfVacIUz/I2A/Dn/aL6Z/XeI4xfzXHiQVbqD
eqOuXgQWjT5hDD1K48ckjdwws8fMZaVLEbzm3rE/qxxXVVCVMPl0zXVcXl7Y5VxV
4f/2Ililli4uM0hvrFxKYOONlKZI7s/B6YUdY7cz3/kyY6BdjjBoYXGbOIjtoo1w
vOexIIW12FPV2W8woYySQrtzkaVa7DGztHrzdMNIyWTskcKpvKwn+bqF4qrRxQsk
q8EBuxsFSYnHMtANAGB8K7fhu6jnIAMbFgmjwZfmO3wuh3jvVsbGoSakgm+QAnJY
PCrl4quw+FGGdPntP+I8Q4JJ9W/ifzR1v1Msz+nahlOtPHFcBaA0fRjitUOm+9LM
67v2kwwjMF2RjyucV0w1Z17U1wj5kXg4UTniUFPXCsNxG7wy+Sq4R/Y80eiRxB85
I0seB0MnI8jlzsYdXoubfc87oK9A5k/tIaXdhtOM7ClAMowZdf74i5h+RGRV5XbJ
eUqqkZ/6MS90hg2YAH3QBuZ9d2mSO2rQ9uBulL0wUCZfkiQT++YDL88qnK9DqDgv
PgPhp+EkcsnVYIAStBzzAybwAMvzt44uzcK3+1gdIoX4AJSJvGW9IpYXb5V+PD4D
seuQ4ASoD2VAuYCbUMoEJj1wU3EEGMbMpAhLxMf6cg7WX5Kn1MeF7c8GhOl87f5/
xBxRzYc9urV9Ent6l/89VGvYvZa/821CpxPyyO7dqZQdvP/YF1aT5wFj6em3tUsQ
BvYZZKj8wDy4JV1VhP6qrCtcAydEx8bbyP7iJNcVJGO7n21BCUuHJUkJw/0mB3mh
/OgxBuAzt1FiQ2aRexzFvCKU0/ueOiIUdlJi9NkYND/7mNdFa2NWPqLUg/zvKbN2
anubnTG4Ot/Y4rd/s3fXUtO5zoDgqimHNIHjLDGPB3phE0iNVcgHsVA+UL2AFy5E
K3PHu77UXVQ0uBwH3AMFT+JzJONgSzW2Qg5HjDQrryO+D/qZuNOKmLpZxP0iiZ28
xwSGmheF6hp6rh/eZK/d5/KTxPwPFupW+NGfok1f6d5TpvFlVv2847N9C2fTilWT
NiFDnX3HOvRE3/p4/g2WQJ1TTRHTwZ4qxzDhBy0HAjkCqIP6BiS1VGusrJ1BJ7KH
16cL8CsSs2PkQqSsG2/A9oN2yOjuzuwugdFHxLdRwcftsOEgahPI0b9uN+yhZzgZ
xdTS0MGEO2YTck8nMg3LD6w7sb0/qkRDKEeZqfoMzb3jyFIkLqf0lJsU1pocVthg
jD2VdmkjX39f4QaqhEatfK+XZ1lRMCptqhBifKhcYQ7eTPnd1KbRgMHOW+mxiLlc
OBLRtu5eCGEvkmLpzjFndjeweeaW6C1DMZei9oy5TV5xgnsP6CsItFe69GuBTNCA
esWUNxma78FDEO2AaWuN3Rnjo7Zem70OHl62ZCpyh9cCJk92Jn313kOWFaiUQIML
VF38ZfKyozi5tmJBqiNrZcZ9I6XaBNR27y+XnyVNcPek41mHbEPB8phwBCOoa2en
pXhTTKGVrPa9IL1RpYPqwBmXfYjZ9H3etX2cfBLTQGfU1mx+kFSBq+lzROThsItc
42maDYKutmXyAEVftpUZI1T+Hy3hwuOnDcCGDR0PB2hJc9GL/7zdxJJ5bTcvunum
2bBCo+bHiilyGGfACusBa3bHB5FP/eAAl0uL01hLgt9NBQ+JJeB+FWNKEPK+mj8s
9wNjmeruYSWZOc/7iUPWvPPuzXGdqzV/of3CUdbcP+odc5SIsAzEIbtadrqeyFxr
f3q58LRq49WwvhDKPR15yjRPfrAVEdmxwBfg1hWrWhb812L0G3IIlFldFIRDpxQM
jGEkU78UqNKlzhpOLqcQxUaRL28eLeNxM6JNmksy0VZ4ABg6ORvE/dVHc6DSmxf1
+eWO9BCXQeOWH7Vnp5+XB5p2p4zeyfP5XBjvCFGJY5W/0KQiglA7WlcSTeG110dT
RGeTqImdCxDxILxMN8T0O0TvTSjQTNPxOQw5WjOzZZHIp+tjvSA+Mc+tdaGCSO45
7zFcwgbBkXm1enihPQpx6TuB3kahnqeVF/rO0fcFVEKjDv2J9+K9V9hokp7dtiLM
YhHqyINpnpD3N9BQduEnPWDiTgRrCw/+FIueEpFduqHOIu/zz5KFA1d0T3X3FIul
gLq8whP+qBRtwgkhZ21TkhSGr61PklHiyW6MUK69FRBLER8NStrD/98KZOOAssMt
NTngsIH43AfnA3x9w9wvYd+/QA2ZWVjaDTsPinrJXJI+fWWtmkxEHnMaFWDxJc81
UWQmDfjhjBOj9cs0cOMaXZFH05tqgDEI3Mvr8ZUoavSXXIGVg9Sxqq60BdjmYUyP
6hK2o55KUb8MFcO2WP29PSu38ibzk1RI9IXm2JKM3rfpT6qawK7NMxjOrthLs8dg
NtG12nraeK6mD39R0ge7ILORSdLkTs0iLWAknNI+1lsrOT3uEi8qj8zRVp8DKWEw
9YoTBQeW+bZevZBphSYT5qVfP66Jr7LmjMdAV0t36e12mcotKUhh91Mk6t9IUxIk
eGDkAwwgz5K491zuWumoI7VM4Oz4vSztGJOARs4UfTZ7/P4jPC0knbMrKIoE0IlH
l1xZzKu16x+vk+JdOGnXZJvNGExn3Cw8YJqdVMOK1oq8RKEOqIFCStEbvz3lr3aW
Hl4hl+ZVSQ1VmV4cgmV0FELNL0gJHy/ZEkUyYpTNiPiakhVBs0quodQduynjV1Hz
zWOlRNhHE6hShiOyynaXc2JnZ10SClibgRxFOr6NiJQ2sbabFUr+vraIU4eUfoZ1
QlNXZVKbFufzzSFvb1mEBC5uzeoLDgfe4dqExzf48qo4zEtZ3YVg162tXvQttrEY
2MdOcga7KaREgAFp01tQIsq4Pjw0ymweQ3sa5sWamVGsoVJ20a1l5v50/Ge3Klge
ZKVIk0lamLYLDRPCCx9mJi/fsYmlnjaaWjC9pgh+CpIunNZ/jxhAJS8Cgbz+39ZQ
uFyxtGyKGjNeqWbzGqDR6bs7nDL8DYhOzvBUmNyMDttXmBSGxGjQK+8qwCm8Doc5
WDC5qV1Cj4PN4BNMpBylB6yhrZdbBVZ2qJS16/jcbJbmgt3f2C7CMVfWEK133myk
1VvdyZciQLUZAezila0hzyEMEOtNGAmExneGtB/S/2GNopRclJhIlSUvAG3ELsPN
vvvfS2FoO41i43UL6BfYdlBjDcFmOq6Jax8Ga555ds9+CQRk9qjezwpFDf65mnDt
/cbSAhq+Alh1S5L5DiEFqrB0DqjESAsrjYXAC1oBcF8lDlaiizFeesJbRGNM7lJ0
SklVYR5sakmUjJsvpJ7cOLBSqt8DBg3k3P8nXKiM/OcJDWGy7OqVIOV5MsHFPaEh
BjtVXqFumx08nYvVlcOdhVcxW2PnCpdWQSEQtCXfZHetqDXv0FsUkxEsExxqoPCn
f5keaeYEIrFx7xayKyniWpjUrgBg/JTw5giBH0F88QfMSXb+ZeFhIg3Q3WkntULI
g05csFFM+sQ5tGLpOjVlJ9JkQR80sCDQN9gvVQF0EFOkcFj2Fna18+fw2X2vkHfs
ne75xdyOG9hI1j6TYcYDrtOSnowdYA2fuZHPMpDo7NRlQd0ZNPU33jxtSOlqAk0n
EfQ9jMf+aov0gK/XLz84PuIaDrYkJyjFoN/fxSTs8Z8G7VdyHHMEZ+vFidJ42gHk
Wnjm5NTOfYFokOLOGvncZUclJCN77rmRdexrW8CRCgN3E4t4dlLOubWmaxUFNcEf
0rvyqv4BZYeJN3yxspi+J28vlV8DUOdOvEbkw1q/tlUG3KkheIEsplm/snYrxKu/
5q92Sa0U4nQlupX1o8ehDYy4CCINbd6IHFj9q/9sxEuhkeSs2fCrOtn+EyaRPPa5
nT4SsDmicNyf/9q3BhW9yDDP5aN27/9Q1mmzCTK+UxjF8qMkqLudZePsbcoCM9oo
RvFudBGvQJ4gIYsXwNlD9ElEQogH2Sf1xG/UgTSfEelBeLmIHhE2o0LvT++J07h1
XTikj26mcam1OxsiiMfY/rsN2u0yXmNAwYHX6nhpkvYrNfU0LN1Dym4pKR5sRCLE
tV/y1aMbmeIsAoyVOGBDIsUyM2ZG1SJAeU+Y1P9dG9Vg2eZY6kCx5kghf5pWRZqg
pXwRLm3dViHt1ddJjhu2Xcc/Rp91hNQ8kKZ0O8ywOcQ8Cl3Ey7aVtNnbpnC82FSN
qSYs64byk2XZ5qG2Vs0BEdZ2ht4u9Sw9FLK49xdF/tT4bqbu9RDyMyAzCFcf3JLQ
jASoJB4Pn+gYTmyjWmPHoaGfnlkYpLMiiRriNo+cij1LaVII3lS5qwPVrDRVocIs
o6sf4lylBHP2mRK44XS3KWPbFMaYgQi1pkHCK5wi5dQQcQuFDvGC5im/jHHA7JX3
4UWbpT+kZu4W88wQERswtI1ZlBC74n+JdX7hjnEFpdLYyUmwX3ZCrfE8c7bHDaCC
21hubVZQki3lRELilRaTfJUfKHpkU9g7A0iMIWq3o+Aba4ZqGC8NoD1gIFOhLWcN
+GiGFjglhTRDRJxkXGjYwV1g9zjypbhysTSAJ2raqvDxb6jf940WJAUYmQpTxnRt
dyjwLucYD+aiR3oGzpjdeSPbpGrgyF7hHOhbbWEjLQwmN2wm8FnBkRsZzSDsvFKc
tRPIEtn7ZdI9pBHd27vhQBE3nCgEVh7GecEsZo7CFgW53IviB5cMedQUTA3sciqr
a+yUy6d+fB83YUmQMaYL4N/jCgDRcAOTCkOXOnB22pLlgyC93fRVyvlXPg43WtJh
vUcnH8NPBOY7jy5CvzuZRJp1SOpHeIIoHxx+Jcga6lAoNxOmndlZI+2f2mFnXf8m
DD7Kbyabal+/k5x4Bd5Ww3nEoOp+FHpd78hDr3jOCuzpvvn5i73ogJip2DvZZJY+
AGtZYMtFgqeNGzG4Lp5Y9+9dQ9JV5OZI8Has/0vcncdKNE6hQIu8AiUGjOdy4zkT
1XFT2QZDbnceS8DqH2QVeO4cozV6yGbSH0zulsy8T1ypeFBaVGahOLHCybq7JWEd
+UkAszSfSr3MXjjSYYapVy8kmKj3uIwwyXRH89zW4evsPB97F+LZ23Z+/K2mcTs5
eu7SQwteHwET8GJWYJGKO1gVd5PLuuNlrtpmpUWk3ep/MqNwqMzqLPsYR82aueYn
BpSVP+oC7vhl7NknWwTpnfm5UvDg1Nb5JtW71+8gCzYjtg+66RFeBhqlfki8e9vi
qWD2RiNO75/kxPyUwyRcvsrtQcp/poirfdo1NZfBauNvMrhHT+GItO4m9gMD+7+L
OkeLQ1YUknXOm1JExI1GgA==
`protect end_protected