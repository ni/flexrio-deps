`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
YATj3kULTF7Ty4ORuRfFpnT6YIk4rUPRrM74bVTnc4GjdV8oSnW5PtQkMCLOi558
1V+/wvDfc3y0Z8//ksX8sZm3JZWtrxUppw8c14g9Y7owiwp+JumRtO1zuk5xFbe3
0MMnIxxoTKLhyRJtAxElG8sbx8N21OWDGiOk0Xyd5CqAmk9dcOIbxzMjW/wndBXi
maijUdqS+5KiRCM9+Gsp6k/iEAa2LnYTt4WtjkmDD1P5jZKsiMgFck8WOqLymplZ
ml3TTfn1UlLNm/+zD3SFGP0kABAiUT8NK2xBPQ5UzQ6sMFPd/np8iUZ5u4QLTWOZ
hTrU9OSX7lOvRUo8pJ9vPg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="BzW6NOo8eyBw+CxsNNo4wIDxODIsVe0ft0K5tGuSUZw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
DhjJh9S2BY18dG77XPz3hsiSQ73+w0XqfJhD+f+lIDHHVjOB7CfC8ieNRTexgzn1
5W+qoqOEwenoVQtit9u3XViXJSRJ0wfUC5a9axblRNyD2mUbyfH9+f59nWqGkVOh
ieHxkA/DPprM70F3APxk51m7/gNSLICSvbONgLGndWc=
`protect rights_digest_method = "sha256"
`protect end_toolblock="L7NTNW/5Dqy+2kJZXKczEa3js87UJ8H00YWI+92sDHA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
6eHODtGLmq6ccbB074dgNWpdzW45i5jL0Nzx5wwM+RA0eeOHXxEV143NNyQGmZjT
bzHAi/6AyRCB4X9z0c4MjyrZE8GF4crbMH4T59xFHqVrQ4zXCea5w0kG5yvHgpKo
hywlzcU0F8++BgcpEenWRnDFmAWkqFvq/D9BjDe+gPZwKaW0b5TUDOi77MrW6aIF
iXwPE7BEqOOUXR8cFbqwPe2f0CD1k9mjmy/TuRripyVFlP6MWdP1+kONEvs6/gZQ
5S5gkuBToPh6DtjdQb7P54/1rChVYZsZ8yxkcl2jfdjHGHJ1vF5nT4v+d/ZZoolt
+pelnQXMp4wlu+stnWPjqisgL6tolbrmJdeSToJ4KyK2E5xJx3Zg5+WG0rlfsgDY
S3KCaVi1Rpn4rk+nzSsxmvgA+Y4obaCDRbMI8J6YLM8t6E5I7mAqVlhtXXXpFjuf
y34M83vMYL3lIyLNWP8o6g1RR4KRfn23bD4gQoqcmEJmtAiNoGjcf6paX+zrbY39
vBSEWrqKSN4sexlYYXHT6WMgfey1q9qmbodiln7lOmXhwCut6OAIim+2xzGiJiTo
4IbGNRRX+qa/h/MP6fPDedm1L16+ihYUQaIFtG56JgosQEtwJ2zu3avxWVVdr2Z9
BCC68bVOOcMqZq5vSB8W3r1pLpQJOzIpaHWI5WpjDa/IV4LKiD9/nIHfrckf4WM3
ALLHV88A2i4J2KpiooNz8OBDHFBW4a0HoczDG9DBUK+6e/iYcPXBSqK18u8ZyAOM
6XxqKQ9nEPhjfOkm27OkyNl3Om62aMJx1TzgOxPPJiR+8WfXv55pUyexnmv7iCfz
5KsTYHVk1RY1g7S2JA9FUQf9Sr5MLaMW1LBLzKEl9XK+30/gUPqo1/n4uSOVfh8B
w698No6bIptICo/AB77Hj1rF5Jox/FVlqLQx3YlsF3x+bSIy/ifRQ7p5yfW2c/hU
ccdcLCCipHtVV3rMZj7A9MfOpMU86xWORnKZIF5yxERD1pdNQYlo3oEixS6LLe47
DCOXe+Z/Z/cC+9DV/vcw2iz9Av8evQWcRnp0I7GZqaUY0TvwEtXg07AzT6P9+raf
rC5cL1ER3lr0VBjx1UZophf4i41+Ir9rwqRc8gywVZCLnLal/zxxftP+dhoQZ9pp
/Xt+WHpMJXYsE3IppDjSAE0Y9z0vzV30+3Jw7q3wsvFIXaLWfQET4gR8ohlox+zc
dJdi1a1sGY9MdRTka2+yUYAa7mrFvziQcJ/DsKm5umgXKFYL8F/JcdEk8BTSXCdp
QFSM2UptSuePNlU9FwassKLNbKdVh6lGjqg6I0xIqZoeS9rKgUNzRLfJ/lytoK/7
WrAmE0WIRNrm51LDeQsOVH+oI+WVGI9lFHkQAPBKY/7HTJqcbTb+veXRXsR2pKVD
yDHKbE5z/OYNyhovQoa3CxxiufkV2Zdw+2J4uuUd1vky0xCmHJIoNiMHaz3KWKgN
+SbLjTUVYd+DgGInjOfPdM5MhrO1btLWeGrY4gH/PSZ1EGJIWu8uzP8FQJ0RWj5M
hBdnoFUspRk8f+2CTIPPqEKn0STJSgRww61pyHm1zZCoWqmQOb2DNVce0lAR0C/X
XWzOtu60T+DVD+egX6ahPsEyymaRxppnCNCFhi24foqzMQ9JhmlhKFGwTDpNSF7y
SIPxdHDP+sDLz4K1Eate4UtD7XQtK3rONm9aSlxbfsLbCE1wHQD1AxJdzHXtCvh7
1i6Ne8fo7NCmOexYDG0kwy6/GOBJfL1dz50oAAha4MLp34XUHZsSI73T1lynNhDh
zyAs/YrjvMdc1fV04Jxp4G6daZkrsoyqmd//dIvBWWJD6TGEpPGOvUa32/nQscsc
EzY/L/92JJMhaW5QhxnHATUaWcmMUYiA4eE2zxAJ+EB28Z4nYu4MPUXSGHwLGIHc
9wbsa2F0zqqqA7RDzlVrdfQifziP1RNgiRDz6sYMIgOwy1Vt6q+kJpeHXB1jWRdd
Td61iOPswNxBIBSB8/raUVsGV3c3FnGsUHDaslRrusIh9XbtroF2kDQCqoy3vN1h
+Hl3PkMckcBYeIW3wGVf96qyEgWO/4GUCs6yRO0ajdEqH+7TfvtWbtQByw7mBvit
a6cfDlnjDwZr3ZOP65LPewfMJVTaiUTH5GmNt/FvzwrcizTROLxDhABQr16Fhqld
J1cArWJbjOd0fcKerJdDUKReiN4sVhijDI31/vg4AGYDQ07WYygi9qYwLBEFvJl7
G0zegFFQJ8Ki44fi/jdGu/Ri17Fowk+sU7Z+ULFiMIJEcLf5s4VL7TB2BGqZQ/go
8LzziOO2gB6uE1ikTp1gpepkt906xp4bvIdp+2ArI8l7DIVtoWqumwoRroju1koC
KLKjDrwimyZ1KTyMhUN2wqle2zMxN7HyOXSBaf7rTYXuTKHb0V8a9ga0gnIUkvfa
S9trllNxqM93e/YBOKiHnBy3nucIo5CQn7rRIMMRIoieitKqkWRVFrq6RyACQ6R5
HnzjEWTwBUKWkyiMiew3fBROf3uYbFPQYj9s9cCXRZf1xfSvNx2cYB463JCE6aWz
5MpFTW4iRnJHdOuvBAGqc9iounQRKi0LNnQk0piHMFBglYLUnVg5gtV2tOvuUYae
wTiCbvsmGCfZWAGkQwb6bkquDEE5CvyIpSJklOxfjNeJL6/K8/0WCnP6FIKQyb6j
znQw6OgOD3FxmDIqyU7RjKeGoj62Tq/fgznwkbbI57Wi6HKox6i3v/E0B6xMG6D4
6pOsHCqaOuj23ZPqFjrEufLorBIQm/m1weSYtuun9SND6HGeUI7q8qHqULJ2xcVw
9wyU6Uus9GaMZ9r4uLMHEfq+PsooTLfQ20fo4c2AUsn3jXgzchlxghZgtPHqBKNB
/pod2NHVxmPLLKjRGKaCvZ+odLjn5z1hAdTygQiIIxRN4UilvDpVxgMqasnh7HVc
GBz6sdei75JkHXRausOCK0L9oOupVlUPuZItweQBhTjBRkJkRuMUvkCh7JtW9JnE
qu3o8BdGw3E4HJq4A90l/QQDrJvIezbIfCoLeO2XDVRP1Y91zloMFrsOYoKq33c1
vB9nUK9MC4vPCZBvJ2InPurioaFSXJ9/VQI/XPNboxClTvxW8yxguEr0lssQ657S
hyP/Z0L6lN4gSNSjC7Hm2ZFbKLY0NF9/EJvyg4va6jdjFwULGLmLVVmt9sPUJTgF
CFdwu+Edb6oPh/cRaDZvulSM9Owydb5ylX75vfECMcrV4LUZc0mq/qZheI4UN3ss
oo5bbK/UbUKpy7rEyWqMnaN8LEnYr+9Q8rnGxtKyBfvQVK+e2+j6JovjPZfPbuRN
/3GWynwZ5KaMRU0tHlPhXDsljv6SaTYCMAWGd7WpkZZrir97S6RsTdyGWoabUzSA
o7BGWs+QChstC18h4pOD/4oQB3j0oZTiTVeMhMAsm+f24NHgH2wjDfOeC1cwtp1i
5/6OZHaedyUVVI9nnkH/LMNaa9PNJMEYBk+8WsLyJRsATRrDcVuQuVIHc9Uy/rlw
IL+9+UFHp/rKX1Tnypt07M6oSp0h+cbJCU9P3q/OXZBtQnJO01CuFFCYMZzV05+U
RP78hgutX+wDndJz01T2W9/Jh1mKqTb9s8clRhJbqY2vQ0FgC224Bp2goJIf3z1M
eHZNLsfaq5MwbLnsoGRoyzSp3/uIrNKFbfgYeeomyYhGR0TFFzkZeTgj8GHlH4st
WlV2xDgBncu1q7cajPSShyZK8yCX85Dc3IZB3oTsQYimIeoknZI/rZgGyNCOu0n6
NyWu8mRBIO2fUfAa5lCYjHe784BG0XJMIq6KQ+1ShdJgjCTqPGaVflss6Yjw39Uy
sHuDtKHcwTZAOYMojnZj+ehnbTVw3LFLucD4v72rcHYfr7U3D61xeiuZRj4/5Vf5
0jbHcClwn6ZGEmFp6ONO/LtbBhIgsxqNbfZf8AOLyIR+JcPfQUBD2irvRvEbJd7o
ljkoP7MHV/bIqYZpKk/FB4uqMRV5OhugNYOoO0FEGbAO2R6Mm4HO+RHzt6EM/8hV
adB8ynajLM1RNoHZUUTQTiC6JbGul6UC64cUFDIR92IPY52BJuctPLWwnbl6xVcu
+tdNh0ITbyPvk8K4yjn0RyEJPyses9zdD0Lx+/uv3NVF8PGhO1i5fTvfeBU6LohU
r+kbxriuHhzPwisV4AEmv9hCvHTFjuYoQJehNp1nnUAhYk0AY8k8HAwdEoHZOb/t
uZjXXPuX0UCs9WrILlj/cJDa6MNzY9JCBYA65B99fYpwtC0SCM+UV0ANNxXu19WZ
BLtg61zgPpWJ+GPBbvKbN9h5rC5wG9tpVGwU9Oh+WkKCs6CgpbrZjlPdz3d3YCZb
5TF65hEHW3JKNR3xe+DzA6IQCAqckUxKCXq69b8bkqupylSVZ0oOpvNTmEuCusqk
7GWrRx8JdEWMn5Fmensl1xHjun64MKnkPrgz4zMw6pqxRPj7RXJLr3L2b+ReNjQM
a8wopRUaoC7nm+V5iQwybW9PSCL5bQNCman67W3FfcmRa4FKG8bd0x0Wr6dsmwfN
3EzfsOGRZ6WIXxafdPA5xpGARN1XERUtF6LwQF/XQ8cT7v2Yj1Zf0sjnLp8cDYov
Ya5W2RNRCE1JL+q104BIfj1bVqkdbxt32DmHFkkJE3kVHDoP441kUz1T9gG9CCqu
jlfLw0KFzAPYeD4/yOTjbnHeTwWopsim/Ph7vKOWOp/CW8OWxQuxLx4H8epIaU8E
S4DHvKyuLeJwfwW3kdDJFQ5W63gc88+dNaYPtUb0LgrBDYLx6wwvKW5TrVI2AiKa
L8y4mjZAXtnYbB2ixV+gg2nY7bR3XMp9TcoHUFp0MJo+IhSYJi9FSWg6Jk1lkCxH
PuDlp7WMhog1a/kqajCbgkKoyypZBOS4zLVdpA34Cnvn/zTeSfXxgxe4HncRb7GZ
L3jT6IJ0+5EmfFKHryYMFHbkQzU8Tk+SKMBAYpQ1y3E6e3Af+6fZcE9iTJ3Cx+Zn
5GV1O8O2QhYxJ0mct+uGU+l3eodTBj1aF7ZBnqu2c4M6Sq1WkHR92I/f42dhKMBQ
cu80Ko6mZZnUHCOR/srNLJGGeXaCvOL2w/kyh5qEN2EzSgAkheU91Av6iTz1j/NL
U1F2jpOSmsxnG6AWAnJ2AHD2KSJ/WNJEAikU/DojOIOGmkOoZCsb3ZV0sBem2SkM
3XWKEdngqHyo8FSDNUfwJ28xZk+S0wRS06j3b5vHoop5KvTh/TCWVS1QQ4rcOu50
KoHGnkGrThMj3WjZNE4H78N+/jrIhrxh2X9tRZlOHAAUaBD53F1Mp2j6JnUzAPaR
JLspGCPQ9O7NRrEZA+OJmHEPmtRnGuUUXa5+0F9Fj0KgcD0F7vTjhKMoIMo9hPpr
Ly03RNJTGsH1XhyAS/7tqbiXiYqGAOAO7d86a6Ae8capsjE5sf3ZufThJa99/QnD
r5/kSHRXrM0Fmpz175ykIEj7ytJae9VZhmsGgWrSydGFhPpWl4nB4xwEjQVtKH30
3ZuI1YntRq6Vjsoi2N2cKGJiRS35FgnoVNbGScsHFSlw0nPLH12zixMTWrllZtSg
pz8qMpdL+VACrmus9Mm252jST6zHMYA/xMEXSwUrSLh//1Hf25eeaRDwLVgNt86H
+Gy8l+xLQj5IwEF8whqdW4JsbSXhCGFddeodnzeiAQ0EN2ReYvwZwV3bE32fo1Q/
lB+mI5vjPXcI6CrDJZ+CiJcOm/OTGhy4iTPZZlrGljKKh9lTLzuZt6R6BadiElLr
s4BXuMS3nVpcNBigL8a30uqJag4yqoCr7UdNK+d1ykpoClIsIasYktJjunDXHipN
3la2kc51qHc7B9PSkAezgtb9kol3ugYouOER4stfeeTphKpyoPKOkHUeQ8Qp8gSl
nL8UIxz2tzdk15hE/TKsnMRRs8BjtHKh6lbz+iO//4a7eVD/gwWEFpJ4utrsD42Z
YFpbUiS0CSVFDjOpJZrUsD7wRG8c79CHkXwmW1PSK6bqwWvpD63/6o79WGpTGQ+D
GPaC/xk9uXmAJpnFAMfn5QHtXvRGqB8Zqx35CjUugIkWPWWI3irvgK937VAqbad1
CXjQW8wXnjtBOs6NAeo6poGlFWXGc5La6kffYsJEEeDAGt34R/sd+yMwsvkDQYRG
vzAFDxpbllNJ5IGdCZLyvGXFrBDHPbyw6K93srHChsHWMG6FHKQNcPPBZURcBqsk
wIJfYzBnKmEsREK9kLe5sEXNmPS4iu+9Oln8VzvbxmRjO/JLsSjk5TcBsl53mb5z
0xACdjU0dLpvWbxDwSPoWDjwCiwOo1tYRaVhBBkNg0MqJgFREKWigd3waKpqWYS1
AUGFfm4NMptHaKfNo8b2HWcmUp1GflcaDp+Y0mKaNLihDDLTdJvHHz2HdgFWvizd
WcIvhRvttQeQnUxLCNF8JpZxR6jEtVZuuXjUzauSfX3Qv0IXL10RvDAXznQT+SXf
HWRkvE9888CJkvDdj6D+hQCjc0QdHzD4Utc04P2JopkpmAXAKWsyIip55+Qjz9kt
N3NwQ/XsoqLh3rffe2cKC9Ulju3SC0AXniod8EklkpeldZsqTvuhH0gFhFWgv0qO
BNXtgPUzRLSxqNWMkv4JMOY9X8/GC5dbMgfHM2VuaZeFjk+85Lg4MsWgqrTrsIvd
34J42uU0gPfsgAVqYPSugH2XPKabkbB5+gkiwQoe1GVjStBIiw6tb6qeuhFv7RQN
0K0g4ZyUdstFElF4+VqcQbg9W9gRGK7Z5fWGgCMxrptmN0ECbvdYTx7Z6M9n+nCJ
6a9NMvLn3Umv2Ic7nfT+xORyjRjDHa4zgx79hbHbKoB6T8c5mnraqZU/bUAdQ/H1
jDIdnjLPCrKMiQaves673cgp5l6jUA7Fr5ql2n904m48fBjnFZBsCSbUILpy8Egc
7rEWylUk/5GibYW8eQbPLm/9pv68NsQPLLZLX7TjAaCFDpIYD7t3gIYIKXE3HG4/
c5TVc7sLskFR/2jI6JUhHnqJcUyaVMZj9alTXyvAI/YTRgEaGcI3v6vphTDLPYm5
27RwfxXUYiVKJGUG3KR3RdRhcaFyZ0NkXwqCrBblTyeoHtig1Y+iYJURRnE+yWOC
i3e3wTKJQbznxEmKSpwfNc0iSyp40wKlhCrWRUs5RxTRFNUAmIfGE0eU0gnqP3xu
6k6iOD19sjoytQUiHzGZ5ieeaf/P1puq173lqh+jibgxpzbQ6Z6LAfOXhfWiSlJk
kAeATskvpZFViozOUaQ9v5sqsmjnaDw+INGEVGSMmd528++8fwnCWBopVYdNTh5K
+CtY1m+8gdvtaUIXEKwMXHL3tkkdTGFS4CVKvP5/ajEmVmvhesT9rM1lXE6flFNo
c9Q1ruO8lInzX1wceZsXJYswsyFr7hsDDtECgwxxWIJjT6UfBtiiFvBksYlA1g2T
M/xFwfN3r3F8vJENqyp/tR95SLDuaa7VOBk06/O5xRssHReW138bKDAo4mBCNCgT
zkKhta7696u0EShLuR6dxoXHIX6Xqhwi05gWzluf1DV6c9HL2EAGYztVchBDb+fO
IvJ1Ls+XzzJ027g6gajetuEQEKxizjj28VH29ffjK5PX25UqgyG9DpNVNbn5woQv
zg27flA4UdkDP3dcRWFKYBetwHdVvnTPWVoRYr1kMG7kvwG9EL2RSzpPF8PY/bKE
TS+J5IB61BId37aGor9lAB/CB70FfGTWsrSY42JrWg7FN+S96IxGLPJFNJOnPmSI
waR2jrnje/RXFL8U2SKpzLgKv8MFtbiZ+/8GO0PCrWx9mT1aXRGkVHx3uV0Ux1Ga
KLCvf0kXNthYDoqzWUvQRO9g3utyYbyXQQO4gCzLYWMIiyCqgnmSBkcEi9cgyEOY
4cNycG4vJ4E6dvgQ/ocwtZ2gIJSFdCntOrOAYsVDc6L4eDoaRE+41TWA/wRN2J9c
+XQoRDKqhmXwHB4jvfFcVpHbkL+IuLUVbWDW0evJ2nroHivlyQ+cVvNpipOpBZRe
nQGoiY7ysp4Iht3jbIyjAawHt5qWkOXrgI6xwPvJ4T7bwbf4xevz5gLSBFVBOqSL
JcPwZ+bdIBKta0BX7isutcQM+ROE8NfOr1gWWMC/yA1kb8HzEKx3f1Tak/u/Asqg
nl7wwQZlTSL32N02DxJY8CgpyCqzQfJeKoP+QHwbLeDwkGK4XvTTY+3GppVazTG0
XDE3T7QBY1o9Te9GlUgQnCRFD7hAcAAACu8rE/snao3OIN+JfLxlG3lByz9qfgNy
4fg2/I7TrrV6R8wJMExbzwrXyOqAmCfELbGkru3RfZIRuch1ct40I+wJdQnKWuUD
3MyZeXtfZ3NYrco8cUUNZkI9MbwF0Ln5ZI95ikxUNgWxkokGoy6BjiErGrTEcS2y
gq9gxzdECajwspTGnOLu+LYM6g+8nO787BPrhshgYmOn+F6m2hCBZHhNeYaFMWJU
rv9uFIfg+HoMPKTvcyXf8Xyh0AeIqdKnjRpZs3AGpC+08t+gkOO6N5AviGLYY3n4
K6BKa3rj5AkXfZ1RXxm9e5fv5ZX2lvMYS8yp9vU17BTNuid6wLKi7WfsryU+W2Cv
90DiasFxWB6A6j9HFF/U7yR2EeB2GAO53jFkNUwUxL7q3iLfI7DtYa8nmeOoRDIH
MCajgsKxsKazNgcQ060Sj3DKMGhb4ln5uTWbt7zC1JTUEHF9eMzhvz2/5+IZoEzj
BHN/bqO+UwzH/aNWI2y4nLlFIH50tuA/YTSPFrdLBAyQ9XXj/GwLLbRgJIYA54dq
sNR0in01Nno24ap/pBANAvy8mnGYiGrxqTGqFDtyDZLQBlljO8Uf7UvVHzqz0xJI
t61i90GQBNgsVwUL5fwpzVwJkcZtD7g8nTQI6woJ5qxcGG6R7ojF6FPss9ebrlPv
HVX8kudms92+8hIK/1IFsfyVKUICgI4rf3dnruF+ePZMiH+ErNSlrptCKDJlSIMi
zY+TOVvP71PKhQz1BBEZyLRPogQwAT0LHdwtenHffLRZ86ntsGkxPiXYuVySWc7Q
20HOEhXKSglQaCUSuXGE9bmcJzV+tfjbTa8FAWKs5gYEW7atrZaRW1o4bGe3TOG5
39Wa4Zq5t66V51TuS4We9oDG4ejf7q7YHg5jWpJVUQh5l0cgoq5nZO/WGYlT78uR
xmDVYkge48SIlfxvrRsAAgZiHH1+llKsuSAjUej2DduCepvzU3KsJMD4Bddyk3Nx
FlS+E4TEgnA/1FGTOUH0fTT0ZC7Hfc2F6PzzN7OqsGfI7F5RXqlJVwgPJk+8bjZl
PACZ4DtIDcUewDGR9q3B+WQuDt6btSD/ke7Q3NKbNwrAoSaRhp3GhTmP0ywZnIQ9
4pD1NWzp1rhohyfIGw7WFou1YOaqWipCUi1XifTVOGhc8el389qxwir1vzYYPvrd
0d5xXK1eAdQ9k+zuPNBJbicZAnsVOU04ZtO8oifsrk8c1lhvqENIlImWLmPesS94
mqKiSfwcw5lQ5E1C8bjZ156nqlX8wK00l/JlN1xHbwSeArLXRaABncRtBNJGCk/2
+iTzESC2x4B6g9efnpLhkpUS5b9Pujuk8OXROXrofya/cQlLKAc8hYh4x1Fa8jXm
F9UZJ1JtHtW5Lpj626sOiArJprDK0hU5N8tQEOBwj18VhrqYjnzNfs0/5KClsA2h
8vtpciWUUQkQOm4F/NN5DZm3iW3s8ZsyVottKJSxBzI7oNdfIMDxNNo0SSiAz8D5
dQOnstXWuebFAXHDGau7DPKENZASCWILpuY1gMDW+xkagMp3l+bfbNqR76KQ1HVj
+BxsH8fG2RCt7D/VpgWqsA2Fo/uDpI2ZAyrdsAqwCKtgZ1FbssyphFC0ZtNVrbAY
NVqeFgno7WN54oNI6lOLxOR8BF3SgsCYwEThKNcNXu3lL/f8A+hVDmczXN4++iqU
BLOQk0g9+3Yp6rK4c5IYsNibuAncKOzmAXQXVJkZX0iEBekBXfnc68zj5nhrEw5h
6aZzcPQfvfLAF/NWsDQV4yfZUMntoBHZmk3iwsDi6Skoi0FTCcvvynCCl7jWV5XI
e0t55Rb3acWAhNrr53Xu4ga6bhX3FakAuYEGfyOVjV739DlMxK8XegaQyKLLwhAa
t+J5z2hY3YAoEBTdS1wiXLBx9Uu1+7pM40R4dVl5O5Wpd4hrrbKTzbUAhGSirHn8
nWPTTq8CIfQZ9LuTUM/JPYUtDirBdbQo3QgNExzENb0El/8rTyKnJSBtofFwvo2s
9kKLh18Nvg5N7DHmUPAfqWpfJ20AMua1YnkF4WzDvO6+S39a/uVoVo2s73LH2nii
AwiWVmaho+PXaEAuW+aeiVbzHGLA8pNbBzKQs+PJTbXs0Fdwss3cJ0QKsruo34IF
qXV15NhqNC+iwR1CHm/QTBZ/p3Ws4Pvx14En0KJBQVNv1q/kbJFGvuxqGloLxuh2
4OXPDQLRrjOcnVlkZZADrZFUdOhItGO8pKYauUwynZa3nZem5tHJBV/z/dhtsQ4X
Vhs/HcShR5TLLX8dUqGW6IGg1+iQojHbyfJEIPrMlwJgnybE7UnRrGNv0A4JVvJI
av8pceKyE0qJU4NGbIgf9rPkEDujQVg3rs2I+ev1vNkPkeltvBbU3/9hlaY/SxfF
XwNXIoNAnUW/EeDxM7nWFaD9QA/knx9aSlWpOx+wu2Rrd3JGKCBD5cMzklvlYfjq
QdAAWiClfHp8MmeOiF7eC7hu0w0gstwy3kICc8CN5Ueuw8lYF+he/6cvAa9wd78t
PGwdW/Adj9vHvtk0l5QVgaw773kqbUBGYjAcLm6HJc20uF/CH/Q0ZcOeVuocWyd5
NQ9rDgnKl0RfI7fCB/vpmcRU67I41/yNupzJcY8desaTyYFSyc+kEmLRpfBjCCPP
OfjVwHlX/Ss464/s2pFTFYRZ/T3pmCLToZ6DAEivZE62nMR1Y4TE3HN4plGSnyZz
25rCc/4RyUgxdAsbXD+tW7LwquGfi6pPtlg5H9t9FlKljkvrn6Hm6eMa/D8S5Ayh
62asJAf09tk/xXsxLwVFkPn4vc0Ejw62kwY//a4+7H1Gzms3TAffSPud97Jugxq6
YiJ4UXo2E6gM75u1m9aSZ11r/CuxvmtJr/EmjWSBmTVQPDYQs9nWS4g+JI3wIlvK
0mD/0yJpK4lIB6lsjndH5YtXwHvNUKYP1krRSQY+3PSTTUFHdT/yjngKtewqwUnq
chwSurdHRpH/5VFEEMZBJHmNLtgZgDOx+/EoWS0bECQ0FIhpYonj+ujGegrgl4dr
1n4Trdz1HDtVfatQNLub/AuhhePELkkj12jVVDO8mdfPU1kf3k+f+iZqi84lHOgJ
WMYtkO1lxDkBAsJwJQ+ougRPTe+zS5SvR9ZNCioHQHl/kNRUlKu7ubK04d9Uj3sv
xGyFvjyUztQfnfea9pTGxB10bj2x4VSsNRZY7GmPbiJQNewlr4CUhnX2/P91TgHn
YfDI0qv+A2tcF+JmELKtm8sO4Qs7Z9S2VAHwVwFoAJj9pve5KSdY2/jMS4HPS5js
q4Jo8Z9ERwsRNtVzb3C5TPbGVw4dnAYHkbzPae0pJ2H6/lLoRisG2NxfiMM69i4Z
3n+XpI0q+LPvz5k1xhM0ELUmejsNLipe+sXaNRpsfalvo1gL4568n5P5a1ex0OuI
own47CUzIq+3STF5Jvhy9Kx2mHTLm5AW5VrfYRA6fTgAfc5lFl5FfJyFNwipcELQ
/4tI452obhDdUQ+bUDmPflp7oKZfheVDhMl+NZjXPMlzCLtFErT1VHRwarSnFCVz
8q5pc3fiYIkMSqhCvap35m1uxUsWN95mAY8Pw+WxnaNOuac6vXkn/l2CpxhhZP1W
0LxDhhZ6AD2VHNX1f2AIJCtQsSnZqgQkbiZa2ZPz7ir3Po3TuF+bGvn7GQfMa3jj
3Gzflf6+HoqnbwVbfe19vPwnCa1k7wTLDqc+NQVyH1vDKZbtpRilx9q0SfM89DaL
kFSiJMH88gPCoumxOBTdHHlJ3SAo6vXcc7wRcZeap7YzCqeECnjjzX2SV3Ywse3t
9wpK6tAWhro5h3C3BE0L0nEcy5xjcA4b+uBWEcFSdBfxMZPAQkuKSxa95z4lpkAV
I9VFqKmxBKwTkyZc0KV6UVCbhFZU/bEtX+Fv8QB94XppgHbgbQDZaODPuFrlKSs1
AG8Ek2OW7J5LWGNx6VIZdjILd4NSsMJOmLr8erjDkKiZecFB+esEkCCd3x5KNRmq
4iEfPej6mv4DL8h98w+T6Ppew7T7MYCQCp88R3hWC3+qQC7yupBX9eqxWOrK6RAo
L+/Fbu37+Wmse+3JmVKuA61NWz6B1ySpa2mg6pH6FmyarlLl5U19lJJsHS/JnOJS
jLO4uA10h04lhq5pfkg0pbXzQ+mJVciK7f9O8ZSzQVCxIrckVnrW/dpu/YWuterC
KBXBVWahDpaudxFpZi5Nz+npG6WbhoC/y2D62N1CZDHf5c9I/V/dK9/fW0fQnfG1
6lHswrddaTDrrLYthhM2YJNOmjlxnBb4TFUiC7pv2DqMVQoMZAiCGe5Ouerlwesn
z7CC9big5PahrepcUdTMSXrfm0vef5+7JW+E4ikCPQ445lHeWK8vp20lHH9BNbNE
mBZ+aOoibJSPQo9vbNlP63DEW8R6Va0GBkzuhbqpxA+EG67/btQ2lMACO9fJsKfp
w2PLEuCDu/2wPosyKNmEDqGeGFnPDPn31Nie40xdwKXRo6WBibi0uQ/i6r3zRQPY
+L0+up6Gh/TenEhRfCcrrmdF9VpMpp+BcRdzkKiBe6L+au4Mqq4n9V0bheam0bCg
PA6auR6+eEriH70JLwR68PmDjix15PrOCNEebq3sFwpdc56VtIaoFijSEivLpRXL
l/N7/B0ZTroFNIDZYyzyT11BnxW/XEZFCjsO+xlTOP1lFsFB4KhESIg/lnXY2oPf
eL+cIWSqDe5ANnQX4lHCypdq5SpHNv1w5Gc4aa563tcNa9UZPlPfVC5U+ijBboZV
OVSZ24nDBhAGvEOsCq5U4aD+FDghIjJtn1QFAEsLvWHVGLn9eBAMvqlKpq75Nw25
ye/7Rtyid91LFy2qjD14fG42HtqBKFS4ECFDn2LcwEWjjLrOAVlgUfCJwrSnc7/q
R1cudempirq3+rp1Gfkw+JbHsNwM1gh3S/lAgpENci0Mt/FDAiDTlJXmFEKzO5VB
uN0KPP8KN9668NyI5OFVNbtJ6htPWBwJZGSv8leahJvTWqmdft/WQJ95hjoNmTZ9
mYo9VudF145S3Qkqnh3WMfFNOvtyRv2cokYZNsVo6hhswpAvDYXdqvx9R4tHpub6
u1gCMaO6aY2P2/02F3mCNXPUp1IauL1Nsk3WI153JP+44Ufnxdii0QDnA5m1A0y2
mUpZ27gfTZlORNy9bSrEVVS4dSFLibB8ikp3BBjLtux6glqujr5SXdwxVGp9zRjW
mdWchlNJ6ywJpDgqsYl0HXG+EIuf7qcZDOp7cxAraTv8d/VidZtQIDHHNB/ObkG/
q+7PttxSXW1/mL4XDzx5RhybAaY/oHP4uXBtxN2NMQO5y8VjOqxdtbqeBYGnwKwv
h+Okr8mDIL17HgE3cG9jJF+NUShYZgWQN7uSsqjnLwbwNzFe+bONPhkrs+Ho3PrI
5b0REU6vd9UvkzcjnPdZNKzbtVMrt4P9xLlBGZmvylozVByWtQBRWAtqjKakFXNd
aYh6Zipb9j2HyU7NbpEOO5ZwIcXjWlXz324fYxqW+khFGbrqw9t6aqIqyDSz0Z9H
brLa9EU7rjKVUPz2lDqADwDi5wC6EQl20sl5LljCoLkTm0jVDOr70Xrp5b+9ChVN
fJXH7tLjkMLcWUPvI63elHHMpQoCqhMF+I9R/OwxBv4K1bu9PknZu6sqRwoIwkUb
0AZKHDAiU004TETkPAaUWqIbXeGE1nKCct47GvCKXDD++c/w0lW6866jwqOrLLNx
ALadKoeDbEQH+OwNQWiU4b2Mj8H1bUNQ14entpGGlBqK7Yzp47Bsyemrvv+5zAgR
wtAxDTNbgTH9NtidV28g1Cwm4rPbGL3cgbH6QHrcsHnAJPMFDy+znuhb5JuJk40h
Mh2e7Yt4muU2QA8Vml7v+edxpK+/XgE3bdO2c+CNthVi5ZMQhMZ8oMxVsBe5Jvln
6J105ujpWlqw/0mZhlAKBcCt5gR4aXHD8w5cCpWSQdiDLoZI97yr8pAksnwJKIr9
p7k622dP7C2h4jzXbosRJHsAz5TITar/p6hOlFoqGMKMNg0sy7EjPPqiCfBkawSR
q9Ptf6WJ8KMAwShA0kowIPJxnFVBUV1iumIyev+WrSibKYe/xVtLLih8ESL/ZCb1
/PMtqd2yMBuZyWts6o2owdMfx36ORLRUhWjv6OTDYdKUdArIAUabGxQykGeiSTRM
pPiVduhAxXfr2lMJNJ1Uyg35CtqObGoVVtVpX0fyN1MvocJiNpJtVtm0EfbCFxku
UrHM9fDCsEa7yAvdMd+/dp/quQRkE1hbrc+rf52ZiD3347KtOE1Qi5g7hSMb/9el
GiiEnBJMPqed+u0XJy7rOlvQvaCs/tVB659NC4BetOu6Qkvru5iv7QMdWbAdgHLg
3/2gb71190CA3ZDYGNnzBrNG8HdYIRD5K26ZqofzaVY758o/mXv+9RMWpkk1En+2
RW+Np77xF655iSMu3MwciXuawNEz2mu2Se++oqoT+5xMMSUiT35aP+fuUhBbl9sE
gEuwNpkgegvb1Pl6bY+hDmL8soYteZE0rV9cqkqjKmk9uQaT13jdptT+1am73Mm4
3AjuiG7Eqw+622e+dXX+j9cydFFtUmjeHhXGmxpxxEw5kmWCm1nMLtj3STAPjrIO
SuCsJa/J4gnjIPlqriypA3spGph87DP3vSguwmYOchvNtuikCzdHGPyjajz28p6H
FZg9DFaGw3SdJxJxZ6HYjgos8kdfPgIiBmD1kkxv/37MpMPnaKWgBOCbuQ5VqPbs
Nhd3yU9QH/6/yGL8TUC3hqlBE9X2sQI0TSicJM42GlPwf565D6tT0rIlDun+Mqr9
WSJH0fQvr50HyNetpeb9SWmvsKkyaTIqmXncNWiJd0Gcdage29RxbKM66BcNeVqi
MXxw4THfQWMtApoA37TpM9vqT3eAdL5z/HUjtgbUZqRveVcSXajhzPm/AK2AFrwi
xCAnSERmgkt6bJ4hQ8GF0mSsSwChpSAPrZSOtesYldwwrfjYj2NhaBwyH3A9G4cz
KvQMuJDCs8M+n1lJVecKAW6JjH09kYxFFPgXtAbRHUWHaYCS768As58nLynNoY6l
oONawA2SBQk2YdFiZy4imvgkyTs5kxR378TArqyZ7/xJwHlACB4SViuaCu/5Cn2V
Siiknxn+Vd5dhSNkiAELfA1/xS98YXhehZBQ11cKXYdHta9ppHARx6ui8CciD+D4
S4zsCKimjOXq8pCiYT7+ml+8di6Cuv/AEzxA6X0jARYuU+RxmjU301D8iAO7X+tP
PPVe0Xq2gLs6XBla6O4PFhm2WG9gxzGw8pvgmu31q5aYrnz97ROPnuMLEkz/+pGa
+fT0hzlEBSpOVpRf5Ntf3kB4SWUpzFNy2zXsVumJ3cRMgITpfiF4qFbHQCob88Hw
0A8Mf3uJ2ZwvAa4QiOYSaibKCbToRQpUMN7SgbOuAeCOqz8rm3vQl/wioFx9fRaY
JhA5W9nioafRfNYfkwW2uuqcl0JL7DBfX5wA2dlWmTCbOyQpPcxnV+unM/Iv6+kV
tzhjv8xnBLS0k9VqTkLEhKY09XM7ARN0dawzcrB5Hehq/ZQqPyMthyWRmW+EiZpQ
PzltYpGHGQVpVw2RMWA5zSgFD7yPGGIuYGwb+xi6rLfrc+JjqTOaPYBSo2DcY4G6
uhFvkvldqq/RZD28oA+TatFjDrDfUp0CdgJ5DYCvXEBfIoXrJ3PpXiLrUaYAaMLq
wEYfN7ZB8/rK838ueg3tlztfvI0GE/3jf1EpqLGN9mwU636AhKeVoyPVGABWEIFr
uSHFW3Tfge8kqn97tF8m75bElF5vCSXtE0/aaN0apTu5ZKXLuZFZLomO4nbI4Uhx
pHwzsuDtu2xFiTzdqf+EQ8SAdOYahygdNg+P8AvhmJ6cAyObP/OubDN9FZtOKV+y
IvXxxQNLLsAEobWxvyeaSgkuFy9vkA4ZgCq6FgDsSZtJDnpPGExGkE6pNztiQV+k
WkWorPEkkFm38PMg2mFXmWUd8F/jBzBH8yYsOpg4aIi+BAJ2brbVKdHTzO7II8/Q
ADw1/vh+w5+osAguDnlw/61dQmdAy+9aFI5AmDbK5SC4IO8x2dfGWkwwLXWz/zhC
0XuAzHUDCF+Tmy/DDIHb5engyg0NYbaFVX9GG9HoEWaw5wNn92am2E+fKgk+Fz2d
hZa5CXCkL1K7FcfMsVc7M7Cuzbs8iAf0fjJphW19yR/njPQjgEEeZ6iC04O2nzvB
HHCBASR6UFs+tBLcJjHHEfK9tHWRATPWInJYTvtW2TBY0ZoVZRgNvxI3ArONIk7D
1BeaoWyRLe5iMMKdfMof9i6g7pvc3hOGQyLBu5ZKk61+KGcW6Ar3pwSE5hce4eco
ly7MeKCC19g66yTNFCcLnaWFE2OZRXlrXbHiqWYnIxWids0hUqWaOoSlYIcFLfHY
UhIeKW93UftNyTjSQG9BdO7dm6y0cph1f3qW5J4uUGc1Ys7uQAHNoyHRCSU4gam4
rdOAzRt/QcZkxRQ/4pxatzkT2kRTsv9wg0KTsAb/bKqVyEQL7DiuL9rsBUGog78J
E44miH5LJgPyq9kVoMevh6SRNU0+5wKbqSoxRjdZ/kAAtXXyJZrK0neG4XXE1FOz
rDca3o9r4Se1i9100urmuQ1cvIa80ua0rmtxzjPewNJKISBu9Oee7r3BCNmmk7Cg
rIpGk8PkKPfMPzD7zUXhURSqluxjXcBfb9LTiewnkRQhWxRrT/hfA7HPhwFw8cCc
EoL8i71ut974XUhNoSv4U1gVSeDRnOFl+cx3lu2sGdzqVSmboCkINwKMIhwFJZ/3
JL6fnEf0EIEd4j+pFF1FuhW4Vx04DRCuAVq+SDLGw3tOKxFjUQ/wRGbwvcVo36Ow
MGaHGqoIVd1p/jPZa+/nu95l04ARE/X43JUDhDFKXR1Xw0ou5xZVYC6sc+ycrl/x
J8414uSDsX4rvqTR9J6g+arswr/NkrImktCsKvvwl/8yNYT+I5Vf0ustQpe8HiZR
hdwBV/a1pqX21PeZg2HLwH3mrR8bdnGJM5flJtijeAdlR9UDv5ShunRGWlyhfI3u
/aPAj3TCGeuUgyFD+PgV1bazBctGhIqoUJyJnuHcUt17vuzFRjc6hlaSYlbScwM9
3kURm2UycqpJEhud7JcgzJHlfwZ6u8mOZXZIcxBxzLnm4vo6tO/UKtZb18IXfVxT
eEh+piOOKi0O5uUoMA7TXjLzb5NFUucnnX9m6ydnrunQjBly9N3gw1m41vDbVRHr
sXqMAI+OIfzb6Md4D/zg1nfRrNbFGnDZPTlX3h45uGECv+tmJUAYlVj1glhHOnpv
210m+vEjjfij1E4jFIv3gbdmQYJGWV6jON2hQlnmdsQQz/CvsH3OVb8Bs+1gkRRd
2jf0bwDHrWfhx+uf03cOcsl+josUoS+HrTdKFg2gEtKB7qG9Ew0UJwad8Dw4NMhf
mi/K0CfZECfCHxgfvhBNTqdkKgdZz+QEXk7WOgmYdifZyd93nqeXG3cmHOIicWgY
SjTtdTobTpTh5I2qMYdQnOmH1TJqLPr6rEvtsWLxhQlrjtB2eC1QeksU4D+GQ0zU
Vyky158xujdlWnT8JHF4bNe1Qmz0gY6wORAeUqYJlxKa8cR+3U3VMiW7DVToOROf
SgLI+okHNTaZwf9zcFH15jtUHYIMacX37vM8O8hHf5zUEenOTuSdvrpl1GeGCYPr
rFxgVrmpKSkNT6IL7fNTJXB1iUxJbtcmZabwrcBaDi5EjaSEQzOXEp28Gj4IIeSQ
WP0FEHbjmunBHVp4WtoLwHqJaRxKlfPCIWhrNqN39yqDQO4w5xAEetICBsD2Jr60
RjUAXMeQtniSEFKOI06/QHdl5vr2yRH58glHrf/n6Jhx7/nwtzPi+Zt0s+p0lETQ
lOLlDaTkFqNphLS/Yb33Wd41FzBJ97Zr5IzSJHCoCGsKWqOYb42jK4es6FdRWhN4
zwr5N9RFlC2rH70oOWfnBZfQem5vinT2CLWshaNETdmvbCpFdOIIDeirs2KYOxUp
0zpNPc11dOHRJbZWSStKtjkpNansE7swe4dPr5vhk70C1vIe4DLv+s5/60oLGWgc
eWnGOCvY+MZmUaCIMeRAv4ej4RWJMO2M7bFtjLwRjF09JYprzNKVKVwS2vHZ/V9C
8P9wAnvOLuvuPZMM6pCivF/CybCJkHhh+5Jqg9pcFC2ie0F2q3PcTbQkn6U0mKm6
Lq7vu5d4QS3BN1A81nyBLkhiDRCiH1l0vb8sChaF0saso9fBYnxe8mSv4m7SZrw1
OSJXBMmx6Sut/J/OhXFhqt2UOoRPwh9p10eWlXUXcVYuoaB5XSPQWQpY/6lGTAxe
YHb6BvV2Hhu+rl3XHaoGCJ/RhDwo/Ve2MGh4aY9/Nt4Dv45W5fjkW/6dxaaXuixh
WHVG65HrpjRwM7j1sOMhxdrIOrPG8Crxzskg6HtGm2tyPg/Gg+GkjOBaSs35VdO0
Kxp5nFXg5ICOL3ZiUhpF9zIttb9+/lLRIjBcWNUHDWlzeU3LWnUhKAdOn/Kkj5Vm
H+t9qHSUiAi20zENlSP103lz7IWD8iuTZ5M1v8d4obPVl9/As2mleiWY3ERCgbqe
NwAVfSBXo5tgU7wqYHv3V5PlFzf2pYgjfPZASBDXPlLozYdxIncBVMtxoWVTot4o
vMaDgkQgaQ/sAHvs3n1XzKEMYRi3x8MqG25A/Aqpc3+4HG2BhxivsPRwi7k9ny6u
XiPIM14oGcKfgtSQQfp9hzY98nngdvoqFhTy0v2jbNKT7AbclWCoPtjnF3/L1K/t
SRPle/F0k2dea2Iplc8FHZziMjaYFr96tjjLNXvbQXIhAXuQQPy5m35GozorAgno
1mTkfEjMIboEPZ+5rMPSCA510FS+8GIzYLAD5/2zlNSuxK+AekkCUsEBKsELJaPK
G17ixRrXjzuG3XVss2asFHC/bM/6e08nKpzNk9QsVHhomQtitbheMmdHXSNkaT6o
AQjGO8bAiqKjeoHOSLLcJ67qxzz9EBuTWB7JNkePB1yattQG+LO7WSUjnHecnKEB
KiBwNSFZNz4BBhApZbufkuxJjEiq9ZyWAVm+oIj5q5/nstG57qWP31e9kmYOJDsU
EBlv33u33kf4cMwVyn3WOJuu/O/hQ2JkKAnmI5WKBLkBWRFPVcbvAyRaB2GYLmZI
0UOSWiKNZcDdfTSNzkTWixTeGRjfBE+ICETQUGsXyQYZM3MJvRehbS/gMXA2lVBc
epm0REV6PkLXKKNf5st1mpw5bRoeGssGMZfGlaOFiKeFlDRvBd0ipezsnOSyQQCt
mAyqe+/RQhDRtTVb96iq6RLND24hzYWkwU9TK0pq+/2m9F+C91Y7bflEL2LsvWGC
AJR2WrlYLDmefk99EbgJVjlG0eL/Q6snU72J9CNxfmLY9J0LQuXlKwlQkkN8C5Fy
VMzq3QN4Ia0P/afrdybPBaBXVdveFh5J9SAbh26kvyjd5OaAf7oImOCsZnQzUg7q
nA5EEnONFHOkj2SJemcCV9AOiHoCJTf3i2XA9hdDfqrx0IsLmfQbBDtDx+No1Vzg
ehzI5VotjdTGgslSoOVPGB3wtY4RU0dqZLRhJ7XkMwCqEawMe/RNnPmDBiRtoqDJ
/3nVouVArn2Ux335PHtna5AzweekGTkcovuk/WoEAz12wrsE7h1WdFB9PUS7SUP3
bObcyq1W0tyQk33YgWqH4SrEeYQehIb6uz38mVw7uljzVqQ8yfaAdPYRvmqqroZC
WfUG/E31S6I22ZTHSqYnrQPlPmuZmT6947GSntLBfbglgWyY0h/hZgFKuCXuYh/i
ZHif4mCeYfTVjDeXbkMw7im/QWP9mFE8C7oXY9nh/TNTp1lmECdiFkFI0gDF//d1
+UuOrxJXPOGnKMVNQ89QSGz7xSl5SA/yLX+KWPFvTJFB2JrbMx2MksyAC7FBlj6a
Zbnen6DkBU2N6n+iDDKlmgm5E/EM+fPvYHNVIhyCKI3+r9+a/PsuxA+F2xgdS9ky
bNbJkz7Pv9SX6vgX15ohqtE59OihJSGfbBR5E004gL3Y3llkgOsgCY4iIEjyCRI1
bOes0E/ShGRdMuGP/eUQ0aqR8zSDBj90a7JRf7limSQf+o0jmdgHEjK5La6o4kmX
3C12glZLnDIPNIUCwsXQh/OzTQbsxfKke3DEJXtvFVduRP5qsoEzLb6qFxa6XBme
eLSQs4XQL1cRqKGiRfXtxOuVAdIcrXkS0bFyhyk8n/laksj1W2b1eVxPHH325J5A
iYl6QlG2CqawzCjZ+ezJfs6Ybq5u/t6yTDgp9OvpGE7davuOsZnSlWOk+bC9O9Fg
PTnzVYxCQMufb6QrKErT/u9SC2p8tCmQDVzOyoSL7NZVTkAiPhjTX8oPMt9Grb7o
yGHjOMACOMjq+gayj+NZKnihcCstFA8tmpnwXEb+nRBApOf+Z8BTQnGXOyl49CfM
0WitHzIsDqpV//EBfdPwEPvIHwH3xnAh/o1CNXJ7T0PKK11jm2aoyCQ6mhRRjTnz
LhNsSqFZu361FVyjjl6o7ZITn9spaePl2Q9kILt75beI6OMbCCo7mHE+9qkVi/dL
qWeXPmwI5aXtoXNDG+E0fogqHhGOuuaaeL8nD7+zHS0y7iAeh4bYvU7+B9TSIaGk
lxEgytBU8PzPGyGXP0SUu293XwGUyvI1F8Q7+L3lJajzCz3AoWQjl0FWuIGNFyU8
5QoUYd8b0ZEIv0nYcr+g1mRnFAhWIEomqvCOxiL34ZkXXfMT8wjQQ7DsUrSx42eh
H+anTf1qllOGuKr0av55zNhkR47iIue4L8r+MUTpGavUz1kDkmHWKsg92/ubgwl4
13sYxhphE9u6wXigUqLB/MRUZTKRv4u1jD66Bvj9eY9pt0d0KMEDTYHgVjBIIeN/
u6BtvP5U2OHoIWehlF0ebv9kHoh7jKpJTiIzwlfJj2VOwS8BC8C06HDXV4v7p94M
gf1dDy6PNhO7/8CiX0qjwJmteHyDk4JahiZtoKuFVzJsDmc5N1fRQQ4nkG3GXLdv
YOfcCXYXu6jqy9GkkqW3tx8XBE/5s0H6zMQu3e4YcrUGz9/ngnCyUTXLOwHtrYmA
UVEF+hcaEQFrzIdMakye6EahSDXnuAJhZm+68Jl0THBTYpbB7flVirtzKcYhz5Px
Jvg76skBwWAaODXzBEBEWNsu6oRS/Tm6U8aaD4CjJKM0bTgS0pjeZuya6DVkzhZx
zbiAYdzD5RQFJ+g7wL61PBTnGxTwIfaE4LPVgn05NwCpFlBYrb8JNdl2JLyl9cZa
QW+GTDHv+6zuxbQr6ETB3p+x1yRThf1dyl6KkmkxwoPbzcNKKhh4Faq7u5GkwQll
23H560q6hLvQpR84t3d8Qhzz6bGsf0Py//eehsHuIulylZSLSPm7EZQPtflLH/gs
VmCHlvY3Z6WBCPQuZuSoyOuVie9lFDOhC06BLdfazouwr3bKWqpTKgb3c5olhql4
su07smgtsyM3Lo9l0zhvYTHvjQkt0A5YXEXICj7WI7PMJr9A2B8RSsYqqx3dlReW
A+kiAqu6hwPlfI6LrRmsYdQIaWd+7wwCwu8NmuGTmWpRyEtaItuXmjCxyWuoGI+G
jBuQvnAvzKGYluxODbMa3c5dGccD5vdjc3ssGOWoHg01r/T9XmECyj2LSCLa/Dva
CkdkbGEPiSUUvRarUtyF0P57YiGPan6b3bK1b4phROU3cztA62wL2tH22+cw33df
vqERJvQboPKhDPEWvtqM73Vp+NS3ORVBhBbRHrjcEFaK32+Xmi5i05kbKPdWCQUI
yBerwZMSI2ARfSKGiyJpiwXVSQ6szBxlDt5ijbkaqls+OtkPnnkbz7BJ69LsG1uZ
4pEURowB01No91VpMidvZyU8FgO3or2221FuottVfUsB1NSELflc7oe301ve4Ojs
lpSZToks/LML01cpCAiwy9jhOB8KCJ0TWs/ZKixEEVGzaxXtO2EIhYBQirW1FdVc
19vVIgA2FEK0Izr0h0XWQkU0Qmg+0RfDRQ6DL3i0QOyamzD6n7dG+vvmruiAic24
teo0/8ASeLqtAMKk/OjqTUYZ56nollmnHEK36DcxaazF+AJsrigOAD+WgGJoeCD8
RSP44+iD/QO/VEs6f74/VTOQGaY6bzA4ZNY0paLLv8/RI9APtdoqYGVVlmUzUQlG
NRmJTCBk2Po14CfpUQDVzHFdwxwuSlCGcfjGGGW2aBp4LlnU8HNKoZycSOuBNazp
Lrc3NqFP39pzawtjXa21sXhxDzdGl53VB+KzoAcyaC9tR9qFWtelTuXH4hkMTaJ1
2/gPhCSAiZffjdZkClRqaMgsLQBpgEUIlWoSu9PvCVvS8TtknOqVVqQXM6dOe2pt
kBTl/ewVIvSpmI8jufl0TRKsPs8nHx5ceGfT/Ez+hH3eMo18ciprWEEDVC2dAmOg
vpMB9RGiFVzKRgxAQX5InMdyRlnLZdiZRRwRUVlDehTtJWucMk/+LGtcxN+s0OEB
PLhbw29NuBJ7OT0+Nf5f7DRI1w+lhqCP3ujMAWPogm18Ue55DnauoLM22PyaoxRy
0dMQVgy4Tr8hgRWzLbYcZw8XkDiP3mjHaUpGpfDC5ZoykXSUovMpUSybDkGSmFG4
hlLTfFe5CA50f4Wu3vHOc93+8c/dkh8XQiXRcMKiTdt/j+DnA0YasR8BuhPtIIWq
POJUjjjYxbNm9+GWDyCFUE7dbyE2apxx6K//CkWsiFw7wQv5ZYIORPo9KwJP8eU9
ze++MkYc0j4KIQVvol2jPIXP6sSr5BZaN3Ll1UOrSwKrG07DzQLe/Blu/j/+fai0
IwoAg+1aQfACaIlMWQ6B+lJegGE7f4vU48g/nbqRZINg6/QfabrcNNGXj1AVFlAE
GKPYqQ8L6xRgBsvBzbmCoXVbK3WQ6nk7tPAJaatu7RftjItK9cYGfq1kh9WIz946
5ZBuCD2A31PQTKXoHNclWnS2omMu9Afk1o3A5a0xaXa4xjEs4L3daR4ag4LZiT4H
x/aZtt7+ibv3DTac59IjtAAdA71CFqKSrnd6Gs0X+qUEJUueKBHrRY18oCdWOQfX
IdDrqMKC4KeYFBCsoPEPkzwPTKsUH6Dml2TP4XMjcxecocrDIUwU9hQzzpokjsFA
ZSRybCnPRFsVTbp87WyFG+ZPe/FdoNkkXiTf83mEuQMSpC3byBxt5x/xuDwxFLXz
jRm8unATLYjglnyub1TnOqBjfwrGY/RW+yz8QVlaswAL2KZ/8rkQthdHgxqvc4JR
XA5tOmKWk37z+ExgBsy7xBDD7Wjl15o20PBdqLcUdJnfEkLj3Kj8Q4UXUa52VsKC
hih5ebTGtgCTrhiky07ML3i9s0N+GDamewLyGQvBxxD6/Zf+LlxdC9JKQAwoYS8t
z8Pj9yf/8lNVeg164UlVlDvXxtXBb55ngnyy8iNrQKY1lFwTWs9/DTeo5mEGVEdm
8XCUjiKFD2vitrVRBtSktFm0gxJ97I5FSBhnN8XH3kudGKK2y0KHBXTDAfA1vfTW
q5bOrBgkSzOdpeV5kL+SCiCyXJnC9gN2SAg1SWaa6JjB5FW9C6PR/DBPDK2tMlaz
FmY+YZG0xBzwT4RrbVDLHLwJ0SeV0gJ1MqHuPABIrA/Rr3l2wBIrqvz6HIkw4ArO
F2HC4I1IskKNZaL/OROxFSyBIujh3fryYhxFBq+A6Pt6TWCmQSawzsv4sKDTctDE
UuseC6Pd8z6pQz34OL9lNvfD9XnlKpLFfy8UUA5t6t6CeOL5w8gyJFzciH9RnYYv
CjV6S2sj5f3pnG46TP+3koqqpO2zawp14ydTtnzAP0SIxA5zgiaw1YPiMEKiABu/
KCNWuF632j4BFCkmx4lxYvJatEOu5KwV9CzywgcUdiBp2yoNdPvTe+N76Qi71iK2
sBNN6ROZmMj2ek2bKgwHqp8BcZP0BP/S84QehYnXB3TR+W8XCJLG0s41iJjxdZn+
kXALW25kcUbF8r+U+QVWKE1D8tPJfO9SKN+STGf1hcUTkZkPD6RFhr8SthuqmlIS
RT+rnNzc5jg1MTogCSqcRd5LkNUs71xFv61nSCUGko93metD+IRAqWEQ1k55F7Qe
Exg6xG54xD3B0vbJ36H1gCt25QLNXKpwuWqdc6K1eGkEgJjxFibJS40tIbYT1VFE
ZXcTJhYM0tJI0UDg7jTY2NbKvMG6iZKrxh/SBMKw7hrVt8HefTuXu9wmn3VT1HzT
+rBMoyhx//5IGV2kO7afxOhWFWXODTn81ANqLUwE3QCdoUmB03noBsFcURWQhK23
vr6RGEdwgb+x4A3BDnfzGDgwPG5vH4vbqimn8oTo1Z7kSnyYbJCS/fW+/uowXnF/
Ae09ecFnJVwsGzN04jyW9PTXU8razIeR7kkigS/QVHtNJEdiTzJTHZu4oD9uvQkp
FzJYTo4j4AWIlA8tU2wdSoaf5lWzt9o4+i6peyyF04kUI8NXOyXaMoQnbahCXv7y
psM7Xw0nIRWf5AI7+/iYmHZLR6M4/6kipwDehX/b00VC9BSNq5lGONYS+mUHxW/c
yGlCzNOgAfmJmrf+MaZ61/WvMsIuMyeoaWyrfB7xEti/vWzU4roLhOp5bXmqa0tp
MIQmP4toZ+HklPaLRfmzjEf3ePhqlpW+TCJNnKw3G1/L+T9HfTTmVsgjUY8F2GQE
oHqiSxnoKq5JeZ3rZTca22jLg8luzJp5mcdI9w/7wIy2t6C+Ixa44gQ671nMeTuA
/UDOMo0tCpDioq7vQkE2046+4YJGsvPflgD38ombMd+xZ6qf9io9kJo2W+ClptM1
JzeIzi3uMx+cdN1N6rLVyGD0CZQawI5AMdVBWDxfVukXAcEy61BFx8+JZRGPbsbo
vWnVNm7OuK6tklNYUUOhv8AKcYREQyFKK4iEcBN4PKzDAYrzYmvE3VYnnjqHruRZ
lXSFE8g8o/hcI/1OpBA5RAuqyjoR7R+PSdX//7o8/8uAHzWL9ZO/+SyNkof9dwBG
cK6zmEJ+h/IwwYaZ4Jvo2F+aGDHaaOPNSnLktMFXYn9T3RiP2xD7BnS1P79f73Md
TsJcxn1goKMms2jBYUnoKN7C3LG0MokF9+Ilnr87q7UljIvHATGI8ljGo97ij9ef
PP5AuHf+/BDcvBoe9zQEgyWECfCAatv75NNEbNAQCuv3kQWjkg5cPwrCyoN7ug1f
xwEco6ahAeGlshlsbvaa+3IR+uKgoRjZ+0f0r0Q9TeZnakU0/etcAfpeez05jtWY
is6d/oLRoO+3OhlOwcOQAiY7ec3agOHzGeYKOzhIzbMLU56JEo0UCnClh4ghbB3s
qFLEL1PN9bpetAH3/O7V/X3XXVA3a11wna+0SF3sBVWVdC+6EvZUEy2PkL1xnSXt
xZl7IGEfAThJRYbT0hsz8VocXS2suDX++3Oj195Gf82l52WBKW9mohrCkRy0vY0O
sgwhjmwepGwMvXSeudKnZIoRax7djkP8tJ8CdVMmIjcAojiNUYs4Y2OSbovEQa8I
jzS+VV3PgvmOmXmvmDidH6Ta4gvm/7cVKt+PllM8gtYa9oE+SUW/aARB31SlFdXB
r09lvvQLMffznk9z4r9kreJu0S/Go5TUi0mt63asJCny5LCEqpweHrSlE/mTn1yH
GBjSZRz9DpuV5t1FPDncpOVD0SmHP6wK+86LvzHj2aWTxUjT7enqPVuMMcw6zDi1
higAN1f7TOX8NEzf+/uLfXj1iJb+8Sf3M9ww1juqOnCotG+osOeRcNa3BJl8Qj1E
FpZwhgcprG23la49oUigZhTgkYp+RGO6yz0Kj2Lz8wV0NdhV9SO8NqVg+Jf0N8WU
sK+H3lMuPq7U4nwCejoeZIzwGgYJYJ4bPqfmOzz/iwB1L9i4NqxnFtntirJA2LkE
TTOm1ClJklxhxFHGFU2CZKKNCHuxUg4uH3/X7A8Qoo4bgkuOr/YdP1tY7xEaycab
Gn5qw2UGycihM/H0tmqplYn/d/4IqiK4+qNGvwdGhPCeIxHjclLgQyDqkS8w53+f
sEXu8rzwDcxmsB5t6QcDk4yosxvNz/X5KViGkA00mgshu7WEI2NrnGstWpotqKNu
5vPlNOxVqiM3lHmpOslYa6PChV/wVU1uh3PPvjZc2duFkdkhmlP0WUI1I6rtnmqj
mIci5PGgqHKXJO4+Lh/NheK3iiMnPXtwcMsmsH50LV9CA4PA5yWOZjOqReeHK9Y2
UQnjsAbonWI5clCBLAR0vDvd3qOwhXcg9FnGS0+UrjwasJD4URCvA/33Xg5znW+C
usKUcHq817Ypb7WuULIzfNn8FqirCaLiGxMA+QR4865KQ7emjtHcCgqDT7dFlOHp
AWNKFtilV4KTWbLtFnxGmQkIX13qGvjhM/CoNsUSSHxTqmTBf1UTy9jtStmGAKrP
ttAujrGEdpHRKmohA4GPLMlD5+cyUlO+/43bglhR2S6Pcy9Lp5Hu/WEWAfYpMHIR
G6rMMQSSk8Mr5anEUagRkkFxi868J+FS0pXy7hh/MZiJJmMSHa1tA66T6o0NmN/I
qXoOw5T6N+CwGLwRuwk+hSa9imokDU/h8EBnimaSf8GbtWO4eZJz36JIZNZZfDgO
wZePQT80M5AA6Ze4BaRrTpblZdIP2bknTXmWrrgxXjaTmy6L7FsdCGcf1Sl+PpfL
En7HRaIz6N7qnYS04ivCHRpduTunxYkf5GAf/V1pwspjPZWhaJPkyFCXSMrKvgpQ
npHfzVKsNmxHqlwrLayxL12+Sx/Q0FoU3hJCsswaIafgACE8+hIm5ASe9XYicHGL
GJ8bgFhSnsH+ZaEjYND5aNR+HPBLTVdw1vFQRTXPiIb49dQqykbGCXumey7xKVXb
fA27KRFfR/4/FEGz8DX8fwwVv9LJp39vuE43tUlb7AmYAh3iozXkqmiZW6Jn4EqM
j6E0lV8bh2swG7j9h3SfhrpRw1QXl1WIlUkg75JLELHeORK0yIK2N6N6u4IHLfja
+Nna7OaJzN/SyhdwsXRftO92eIAUBfS7LpIWLiSyAj8/ODpvxWZZ077Vam53oOIm
EL1TsWZHj/VZsOLosCZZ14C3wXCLqcpdfHV903+znSXrPFXb6W5DiTkTCfYEgmi7
VUWWo1FeBC98o82fx+utPL+lIb/Yg3VxrglCs2xG62XcB0geR5NAb2Qtc4fS2tnz
5TT44NnMCtcmEHLWT1ej+b0YVl4kkIaX9gkdmdba/PbKVSTBtrPJn455yFYnAJIC
SqBHuvrXezy4Wm/wlCpKiikbu3OUTRXzd7br6nth0sboTHpIcw6rII0JcNIKZqSz
KFTKobgXhcun7nDmgqPvNIv9B+2kkk5KXlpBJi7OulDYHXmtg5k923h0rf/ncUvJ
8yTg2v1KnfplF4g8401k+2IKdrpWKbWPzaFNbwqJ/5mJ1r3i2DiqSvicoFQSiI7K
BKpie3dcIRq5Xq54RHry9mAuLPEGoGY8Pr7Ci2h9J/3K4FYQyTPOs6ekKee2h7SM
U6xRMe2H/WKMOszfweU2xyipyxakjGHelTMvUc0Q3/iz/suyuigGl9m+a5VZgQm+
w3QWRqSopfIZK+soKdCpl/v/3qhr+BYRXnLZgL+1c2tr8T607cAhB4PLPdUXuSF/
tNQ42qQFDlQ7aRFJtZ7Gpgg43XRW3VqzUPew8lZTXFCfrAwYKHKbbjgoUvxfDbRi
vnMEJ74HlY3c3Ge0mC54PXag3jFYCisTkGPnNGLyztzQNIMH1PLynLSCNIhD2XTG
bxgUey0LO0fudhBGG0H0t0IfCesgmgHUNmfm1/15676dbhhfCVqD0FdjbgGTDEeO
PhJvCPS5mSE5KBhWYKRdcd6HAYSN+RdbEIjPftt2RYjTnDsViquM5gEKo/Wro0Qj
8DAY24WSLtUSbXvNyFtRUqUF3V809K8IXQhALVrD/DEG5AEdTT85g7vv26tLQ36t
HDVGRc0rK6K7/MqjRxeo8WLyW0pNx+j5FyX5RCBuerG06OYspI/mV1eOcq6gh6K/
nO3HhHSFTfSxIWvNxSLhJKNh6nzLnuNgC3XFDOWlp6V0dfVBE3CnEWvovr6vFQyl
3JPjBa0VYttxa3TJX/6FSr0LXaBEunNIhgCOiLlfuxRCxg2ti8kp8vaG6BRcxGG/
zUNAdLVwV7jyGwr8FZ64uPe/uUdJki7IQp9p/ycGF89QYp/UaxYYPwK6rC3GVPS3
KIMc3rAqkfyB5Yjkb9RtBUch6f31g38xwgHYo2oiteoRw4ovyrejkwCIpSoRO2mY
ao2fdnJrCvXr8oPOv4jVCRgicGs+g5wq2dxL+zaMzh0YeJm5lKRW3kQgsmSWL6Bk
86R/s+6iZhhKdJaDScFh00Px7PtwWOmk3Z5WjntPDuKt9Xh1azm8TAFDtulpdeyj
qoixoypYXplxq0a+iVtfOtSHqJZ2u/y3w609l8JwZ4uoPLtz7oaAT599UuP2WwtG
HYpKnHCcqHTlQ8RSK9Pt4z6tJ4qk3hDa0vv/fQ8xo3vwr8aAXbd1iHhU8COqALRb
I7atNfKM1Icq4MDR/UHmplClZIvU/X2jQiPO9t/g16Ye7pKRl03ybvU3TE5QkKyw
TwvIGa8iih6tESZSmF0wlk9Zhbssfz5SMUOfp0J4tD1bKOEklEAbyF1i+sEr3qe0
IlF/RN8GntfsXnDF48NHhswAUpAG7FQJRxk0l5mqAtkIJ2fCRe8tTfJeMbwsVmve
W9dqBhyyC9QHtk+atTv4WP/lDO2GnhteA02SqCCkGdb92UKiho95Xrvs3Hhda2qx
DyOSD73vdPwaaxTD0ua2EWla1Vp0z2/xjYMKbfF0qNEXANzdHQozzJgX0O7GinT2
kZ8pB9dVE+URa5u08+FfP4ud1BrdUdKogOGMO6G4MJO10FJJxPpovh8veNCACOIS
5cBk0OqC/Dj7GZ+yYn2dXteJ379sIYuL3uQNghSV551JdEC7VkeoX6acj/H4PJ0o
LJuOJWKXMP83Q/IIWZBmbui40PtBjDkX63dGcmtjkTCYMHMfK7sABnh+Vi/sC15g
928nVXcUFdd08XVeHzELmOYO5APAAWcvdUV1TmLECThrCxLpnbxb2viAqSoLHqg0
GKER1Bb0tTJxGe+uZdF+QSJcG40O1XLnkpYDjUvavVFWDpp95C+xknqaGPL5Hhid
dr0PGKqDH4TehL2ApEtDdSZvBsobBHcFXkJPp9W9Shhj4w8R9JTo75TRWelFQ4fC
2kt81HDIX4I7FJ1vHeBO/U8kaDr03tR/11EzEa9efdWPr351RAQudcnni4xuUyah
cXcq+AZb0LwXAmeZSckTAkkI6Ebe3m71L+ytDDch33yZlXUtfk1LLz4y7Gowt9cJ
u30WhhxsQjgAVZd8d6rp+kOOmC8+MGVmDOSPdtjX+q588n4DRqhfznfyxmDKTUOa
2gJTlNYzeyY1sXW+NGtQFU//nJbEdvc5lrjYhtlN8dIB2I7VIbbhDGNU+cW8H3Ba
jmPPG0vkCKvMeAqfazMH2MSnNe4+DY7kHyFHNmlrxZH5FEqBLUaLAUzlcGvK/a8h
CgllGo0jh4ZDweL+Mj+IKQgIx8QvnjSg9Wqln5+jl/a7tYnSRAp8930iDml2wX/E
vEQ0ZZCAUiecgO6ZyrKFJm+l7kWLTUqugJU3Ej/lFCixr3LoSghZz8DuKW2F9Bb/
QGIBfMqpsIaSMrna36/g/t+Ct+L88OiT4uR9NtrCaMKjQwYY/7XoeC9WyQNAee9h
7ilVE43LxHR7sZKAmEeDDXyZEKXGfrKKDoKBE/cDg4bxEaCcLldEhtjkOm6YQYw+
J0RjsLvKPHZK2YQsqiV8CGqhkmjMgKZnYJ1R8Nd3o/+a+CtIwQnKY0QVv1aNlgIj
KLBjVCCr4utNjy//mCMbn05gjpRQx8C77og3189xmp6d7mT8QaM9uGKrQ8MZj1jM
Sz2ZM40+EMEmdhaHFmdrAOhVwQI3R380y4g9Eq+d9XOKCul7GzcRSc76nR1jHNTs
LGiuCh7Jejxagqr9qlrIgwb6EOP9elNBFRwDXWK4OVn8IqZ+EFj40DfRptLFIT8j
71eAaUECj3av7GgNwMXfxab6y7LBTpcVHoL0pNeZedeYpwxrM9k4DP7l+IWFr5+0
CDPyAlClLEYCElS89Fiv5pY17d3k3cms57VaU1YqqVo8xU820XBEKbyyCgI4m8qm
mlE0nN0ddGCmgm1f1hXWm+WqT+/NjaacDIAdUw18LLd1hlHNb8h1Jg/9aRdNiJXH
bXyZzIg/99YQNmp5hIEOdKNa9d0Go7pS6w/mM7pEPr5gzAB838pjL4Qk0epAtNWc
peVMZsY88JeSnUdWOlfbMK+j38tJrKdMHsCTwtPCd7NTVFUshqwMxEcIS3aG2lYf
jGBMm7oTnBYXtUEuZtQHZj+O00b5KdWZFyoym2jZIZw3eaaxKHtgQOie2h7t2qN/
eqZYUnwrDRzgj2rhWuX9DQftnYlcfSm46dRMDXXd4Nnv8ATFJo7QUs/V+zqBrGIU
wQOOGPooIEMI5hwkv/v3B2fIPnhBRapEl7b7PCqU03o4oInvHsfZuU78DAXyXDIP
jRxJvXek0o1PRuah9IxkIfiuR2/AqRDOuXAi90E+JgQInMRTvnDdDod5jmixlFCN
AF6kV77S6+v7yprUOg7XTA9uprZWcukx05B0TnZ5RIJDTJaULfOXj1RWMksnXj7b
Lrj6mNdIRsN9Sn0hsrKFbyg50zg038IscBnmZps1KfvMTKmFTpbRIEpS9E0AuP10
3fy32fFE3j4VpH8meSLIv6JjNVDZ3oqxrfJRX6SNkZ0SAYi40buuroDvu8FpbUaU
T2E+CUVKzAFRESrO6jc2Z+kW6nmBcfnYDYhpNzgxXCbGwfHa4QjuBS1pwAgbc6iw
Nu9VrNKngieLqf5om/eRKF/y1OoRotNj/51kOCW8uHxb4F7EYkd83OMGQUiT3lYM
zDgWo8BX5btQ3gJnfs0LSyoKfnRX9WKp38UHxPnkSPMU66Vs5jbv+m+BCGmsTIIq
mnDyU6B0ack040arT70/zmzI+Gq6RLQmOoNWQkbgaPvbdkMv597UAzeU0D102rmg
s344Taw/yX8Q8eytumUhTxpZnKLcBb+Ui9DB3DjDu493Lyq4BU5oBdBDmXRcySo4
TzJHWfuqPN2fGSk/nMhzEW8XuAJtkCCZdMAcCFXMv9HsMULYwJgyvnKk5Qm+HQPC
jxcqua/ncwi4b7CAxyQ+SjpBVt2zIQfrPsIYbg9TgzEaD36nKvH159Qg71ZKgqQE
`protect end_protected