`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2128 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
yuiAF2djpiMVQLjverTUdF6hOsMhxs1hbO0pE9LRpWfAp+A+l3oeRqz9RUQw9QA0
pn4HBTUZ1/lH2Ttzm1/15OmE8htfpXU5uK0SZzKEPH1SW5S8WaWsF8P6SrrDkOE6
//RAUYdgMoQ+nNBK069ytuVM3oA85eKAPBSG5vX+9g3kh+SvgzGfGB4KKLpewUjj
imkc0/JrfOgm9N3CvIUh67UQTZo1zUwf1gkqOM3/FL9PhCdsVzaRxNxuB01SN2kA
8qNzWDv/XPK27/qJ3j+Z3BbZHiMbPxt4VHItBpPMF90ovDuIoyv0eFGVGqMMAsM3
RMRpyKPnn5W4RcT2DxP5LAE5fEtYX5UzE8dpnkIarC8Bk6chEHj4UrXtRv9F2BSU
uNBRk5RhBeWof/DGxAaFe6rSlVwWH3y5oZJq5kHuzLcT71+/SbC9vqsfT0dxwbAr
BIxximKCEZcYBe2ykwV2qy11pJ/8BcDSLpPLdVk3pd6owxzzg/i/vVYdDt4wd2Ye
+Dt69smxb2CTFJFkr0S1HzoiZnbA0M45PZfolAH9io9zAUgkYCuUd8BxzJiLaunq
P5kWspvuf/N4qSsJesfukTiLDR7eRdQsezwyLexyDAhu3a9aiTN/zALtNH7TadsO
+AC7wQXvPTTMq+DgiOU/25q5mTNHSt/nkGCX/9tTzuXhSyGdRz8xmj5obOoGWm1T
js3zH6MmeBKGjkDocn2hiRSgI9BMG3aE4LwyDMdi0Ug0ql7jvaH5gh9hvGcCoAjR
A9xpJBI8iVh9FkQR/L2jRpRpQgCS1VF/59fYzyMoAwxoz1sAn4XE8O+aA1syO+gl
U/ttHwJ/YZLgylJsEBjxQtC8CbAkhhJtnMGYsQN8dFBXx2s+qDSzu6Nbej/Aw5EI
m33HUODNzrYlK4imidx1XMgrOCeEevE1I9HUtAIIiydSCzrvBGTLjnM/luiuzZ2g
0r/ixvmbxUyKYFOUj4NHsh3uSpl/gfmfahQVDR1/NVA1MxVflL+O+vk0n6E7mvXS
vZw2bJk/h6Sc4yfnqpxgSahmkZefg5yiUcA68TD3uc7QJ0zEQ0XjNIN8DEZsQ4cW
9vR50V5T28JVV8Jl/fKVukM1QnnJ5/e60L7HL0NiJ0KC1bEUkFBIhlldKw9R1Q2/
piswEe3INUTsCIdsCKqJPZtYNQOqiF+7POAY+V0OYbunJ79g2Io7Y9l7v4gN6xYh
qrxxLYHpLe+p305tRJhC3mMyPsp3Kw3n5NteNyH4Zo54xbfahObiIUYdg5BbWTRl
j9JnUm4SP0Pog3czn+JaGQBHAumptbf/Gz9ag5Q2ZBNbslWriG+eITkfzsenIQ0D
k2kBJ438Eok6yo/68OTzQ/L8RCJoFOgIaBCfnRs2d7C1QHoDMBNurYk53yeEKC2n
Qlezayot/88F2Ht269XFVl2+K7752+ryxqTJQNSkXag/HGmcuXWhIjTzpEIx5i9T
lRtsFvO3nsHHuX+DIEOgOAZRI+O+ZpCHmRZ0KqAOIo5RIRnf0GovYMd7OHc+Lmgy
Tl9st9tXNn4Fu7E6dnVxeXkqkFLnR/yuqWlyiPkS7h9EHCUarSjRXC3OMDsL4DpH
Pyth58erd2fJxDK8xS+Lg+/it2Eyot1JQS9ADRrEe/BTsYLKYWGUwJQNSrcRNS90
YYUbY6J+vH1jsk8klw7HWDeaauCG2jtVPnSg3Bt8FXJEi1ltAdHEhn0hC8fdkxtB
XRku2PDrbRPQX237q1Pb0/x27Rq2N8Vegv6unzeDVS4l8FBPJQOIZV+XDiHTKzWp
F+dOquuWplM7XwrIbfhPx6zCPcBqjJYqiMRP3x7ucxdZ+He/wtR4Q2/enh9Lef5q
54uH+f8T80xZ4sjvGuUj7Qig0071ui47Fbk0Gob7jfp5VNvC1H773X/9GfRieGbm
IB7UBwgjPMz1Pajcdh++hQzLoM7or1fCXlJ3VI/beBonFnCeVUck4cEPiFHg6AHX
OyzXtP4EP9A6CbKf4yy7GPl+60oyr+jGFReWGf0YXocLoMIOHp/fNRXmT55Hanlu
07X4g2T+arXP/ZpN4aBklsWixEZhgll+nDEkZViCVboKMlHF9TY7Syc0u6jnmw68
JOOvXsJ+OP6Y8CwqESULLNuYqNlzzNQp6L91fa98KkBzmoaJhT3eKEulgObmlDPJ
cASKD3i4gd2wktSu2HM0KUUBzm+nnXGzxzn4FcKb0eKeT5KjPmWXPJn+Ei/AoZhB
XWbNJJLffR10nP9XQD7SMFpqLllpTCoOiDxKdWvwn1eRHWm+IN0JoHhniizcL9e4
i04xIs1QEAzahHHbfggdUzB/rmfI1nnvi/+FtEl19+lHzvsw+4q8iYU7oU6zGJ0l
7tUtJQQdON7kfHhdfOFtOBbftWjku0LzYtu4ORQaAP6stYXSDT2SowBifGzDgxFa
oq+gMUvvBXNFdqpIKzCH5LSPfGagzfm1t3iYTQU3kDhBpJGqa4iaNJAl4Se8uuQg
3Fo9ymtrNE33HLlupeUBlM1fIH0ZlxvjsYFA2dFEXeH3YOdN8m2p6yhGXaKgIlFf
VwX3G7Wr3IEXO7Br+3yXQSkxuQvhm5kkdixziYG+uioyQQsqoWNPvJ1IafF8sTYp
TZBv3qRPo7QpJmsU03xxY+LfjaxxOJZzBf7SBwMS1lwbcxI3gertAqv0Avx/A35O
L/SHii/C57pKm8JcfH8FWw==
`protect end_protected