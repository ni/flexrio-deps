`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
a+wshxinOfsYjUKzlgWtghqNHPq+Vm0QNGnuuINurQQ8Lha8H8C3aI/ldFhxNL67
BZrTiWsnTB6aeUV39hW76WFG4GfcM0tbAMeW5MYC9XzbUS8n7s2rWGJ+Zh+9eUWT
QYznfqh5pCNi/j1qxtyXVV3cg/tqw9DZLUuusKaEKEARbNCw0pgi/SOcwby7S6be
cTY8I33Db9WlNNDYEIUlGGcWto406JZ/zXWgFShuWOCTCs8CrgMjJ9+KP/y8GnKD
9X/TzC8uCAekGroWUSXsZmhaFhaq/x/ZvlRSL7t7rUFyX2YHFHKPhCM+gd1qPo2j
uhFI+KsoSd7qZ+fwSCKqBA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="OeFlft4Oi0G/rChxXwCmulflFnqd8/0I4Nh1kdbonvs="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
eet/31tfnkvvd5f+08yVtFCyJee2+KyFnXKsKAXdoUlIxmd43eAtdF72sPU5fx82
0KPOWyIk9HihkbcL18lWUH5gJlYjWPk1R9FXGSbK6BPTED328Xw1VaSio1f55z25
Tw1j80Vv20rTduUxsTeKONe17OOOGGPxT9wSRv6PGd8=
`protect rights_digest_method = "sha256"
`protect end_toolblock="nbV41SUbKHGrfkcRuuP4cK9UFEkGxjpNDKmXc99oRMM="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1952 )
`protect data_block
7OY/GceAM38wIid00XP2s6rRVSee1wySLusHpZ/+baTrCq3ntNzr8fl5t/6sgMGk
NLRAfZi0mFz95HqoQtuJ3K2Y8LVtb/vYft4nIALGUMUYmvEMFMiZ00sF1Jsx75DY
/8dei0SfYi/yIzInIePi3BvhE6AovZ9Nc8Nic9j1F7t/g9UY70oBYn0NkDR2uVZh
CI91bYk4gpszvVxMNJv5WXoJepKU18kpDBQHQ9t+0TKqlVkusL1pPx5pN0AuGq+X
2od9BPSwctm3aGk7sUOoyruhBYAxQAdNbuhb03gtB1ya8zAlFcfEwIuYIDmrXJIy
1iSpwbJ3ZVm93D/SuDcq2lrKCxvR/gpcjcnnDDd7DeWi76u80CFjBnRez38tqnlG
69Gl2iLZMxB8HpgldA+IiU/CUSvPmfNrbU9yOxZCGkMzZNfYyakm5DH+8J23ZP7u
VsZkcR44swJsB2z4VPm4hMuz4itbBa5Rakn2Rq8V3YDtknlt40ZzvI6o8Q5ytGSr
NSh+XT7o/nKCzHTdT0JfF5oDdpjX0Iwt0ZcL68gXa0mly+6IwWnLS6oYpQyk7Cg8
BQZ3sqIBaUsu0001g7Phd0WksXTtp9yCS4rdjDeCY8JrlBo/c0FlvQEtsdE2A8+R
yD55NqGCxOzIiVJl3Pe6X45Rrdt0qpjpPEJ22huR6lq8qjYYqycmOjVsj/chYfjk
YGpUHTQrqSOEBRKhRqh7TEDuKbTlDt4CHjuXKa/QUipQEBD8mX1zt8bxsRvQ8qYZ
gqDznHPqt5e7oa0ubkT8hocOVPfByQ8fVmiZHEryY+tHjjzttZl+4Dk76ouwmjVe
6vpmzYkYNkKAtBhbmP5iopX7BUU9AXitscWH9f99cANAQBrD2STEPFK5TUFvubNG
V0QLyX5aJrMCCJt293N2BpRmMlzDcfqDrC+QXKAlCn8Z7qGquqmgfYog4aywoqLO
v4KZp0DehORzzJsZqgGdkjpYzrZNnZK9l615xrJk/cpJCUgIyveuNP+VO8pb/FzJ
0MXrl3shm0uEwHe+uapces9MEk381fJtYmci9dS1pTWQ5zDf5AM1v0ECIRbspCb0
fC7hCrgwCtrccns3B/QwGk/dTPVGTxTJsQ76wPcDZvCsPV+6lJ1XKTwyxOUFVzkJ
KDvyE0Si9+fjbca4mBrSyd6ulK81KUyXmhbWAiX7KmSo2+nY6EauNqzhRyhAMKUF
SInqvpBumV/M/J4nf57R4ObIQb0l+CEEIajqLzrS9B5KFY8s8hDv7h3Xwqnv24DB
v2OMnxvJrWTN+EjuK6R7xsPmGHxCNNvl/9rMDKq0+rg4xGzCEdXNyA0qUwjaJfZT
5wHxo87+Uzft/WBn5wYnXBduNt7+H8g2jUykI0JPkhOv/L/BObSA4pgUXazZgisd
TP1Ub9I3bTTVcKvvEy5cOAANtzzOm/0Zxp0wi9Z2FsAOL5v1477FId5QkdAs2kSf
CcpRh4vpJw6pBLrZ50WGXFrCqYFZndg8+nzZ2Dn9vZUaC2tQjoSJ0CDlyijBeVaq
WLWcWJeTDUfcAW3Neq/p3pjegHJ40UQtNLCnBMavl7YuSGhGSs3Abngl3BTcNRxn
AP6sXp+ioH4rTFMIedeE0QUXPfafmMCAGMmp9N+TtbaZb3kUFTCAhQa79EJhoz+9
ADU8Ojgz3MyeALgNNAcSxSvxszAhJNTMTok44J3l8wI98P2B7KQxLCHVv/x3XFlV
x4y341IMHTJQCJ8rg463rwEU4MABoYJCRsR6+mbdV1a+fkEf5KygBJ0Y3b1AOSgC
lT6KHroVwGe6f964Sj9epRL4Sf/fwn/ttsu2tXaBYTEIPqIciq66PV8N/SyMmAO7
On32UM3JqU7wTUP2OzFaf/bFEQ3zkyvFgg2U2ZW6WMT1J38qdrmuNETOxcBahJvR
2m4WXdnQXhENAr7rV+U7IUDbPV+xbJ2G4b45lBKXCR/Vdbt0Ik2AEGN2qWvxFXV/
XCc01/tR4r2ArUjoTHn5FSZFyCx4Kq1YMv45E5uQXoZrOefk0hOMyiD/ulRWuTlx
oSP13NxzmmdU2VnjnZSfRmSWLUWexQBeMWEJCTStDpcE3tERPSGArmPuJQSKQBC2
n1ecuabSkYCosfqjNTJCbzV/RD3a1naQ1BylVc7AzIdxBtP47VyH1YaNWseo5fKf
DGAA5jpxd8kvbtm7vXjEoZB28Eg62+WoLUCvqzGGIOvopOBqQ2Pve/9ZQ2++JEsb
iKuSPoGdYICf+ghpWz4Yb0zECBSb5LIbgNr84r90ew7qWn98e6DLI3VUdyYmLgSD
5NFt5FPmNJHMthtrlLTSmZotW4pDXuzPxoPiZcuBIs6KYO/3r7yfZ4yGPY+jCoGh
xWIQ5P516GoCsTfi9kekmNG5mYpTHp0THutYs6E2V4nnTncQPmq2nvub4A5GH1Ic
JiaZRkr6l1veTYiWMVxmKs6zV0K1EL7hPuUohekRImlHo7v6sjhhuZ0HucF7RHoS
s3grXRevcd/cn01gUHZuaKijRoFIOthbDvbgV9XdPh+qGTEn+ehrKqJPzfwxKJsp
SlL1zbnSgZhe+Tksi8/paOlZwOUOGNU5EzD3n9FNnOw=
`protect end_protected