`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KxmftWdALweaxC05AH1xMMC77AxUXmLLSZ4OLs38LoAyRAfiS+yjM426gWTMm6uf
4op+pGUsnzZQh9rN/4DcQBPJzESWr6bFg5jHtBXMffrU0jT/qgyXJk2Vyj4xEMHk
nyRnky+CcoGDTBUYAewIrLv+dwLw7DROWIxib81tR6n7ecJB1m2v9l+iD8j7Hzen
eXyPlLt8pSL3uHaS1teqGFiKChwcBOWuFx5jhvWkxia0MYzyepVxHR1mkUaNhmXN
iwJQ0uqFmQJ7IKCrRWdM3nOMJMMfV9LX9WFjBAv1tiAgiuhRTJWCWOQ8RUk5Go/7
Ria7U9f1OwawJRAozID1Wg==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="tVYfsBy7mhKWW/+TxJAv+PODTW6buYxQyF8/oq8BbMQ="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
bJWdeNSWbmvvVaWE8Hj8MKY9WBRXHl3INc6nD8cdD1ZoHjV7id8VhYtyH0babydq
225j37vz6iI7XPlcReKgoosWNfUyPbs/L7YmNuIgj/Hl8e+MiVrsy/a6XFnCY7qM
/M8W+32UsBWsVVJYpALTp9nQS7I4B/TGIt8B/IWJvLk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="3zYdMDzewI/yaBD8EMo72URFOqMPsE8ajqr7WCriVeg="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2048 )
`protect data_block
ngZFRBteVcc6SAhG68ZGr07vvk92+Kl0WZzX69hhuG2Z/BjFBJc73B8rhY58Ma5G
u8uDgEgRlKwibwE8mJkOZJ7G9jkF64IWbLxVA6iB+nkueuUxRVvZPMbH4Q4+mBFi
e8zJV2MtbGrDSF9eZJaPGXPv6PhGKbvD8cgRIELDsh4uvr8AbBJxjiHpWCgyA6pK
FpATtAYoVzJQZnhCbgARGlVli1w2gYCjkI4VwszcoRR39eJcY6kDfqpEn7ldysu4
OWafYTpcws4BeDH8QNm2e0x5mFELvQIKIDwgNVcbFNospWO3fUReL6zTi97nt2QJ
FpfPuZMfbNst7dtk7buSJk1kc+QXKoW0MHL/4QOnl1NDDHg4d5DLRngJxAyh9dJt
Qq4K4X14C+72TwO/gJ7FPL1m9pQmH/iXwfGyiXofCCIdtpKbDuhTGmf0P+kW47DY
e+uA//2GbWLJM6SJ2WB6gKR4OUXTtLXYKZI7IXwqTgs0um3URma+gzoENvR2s4SQ
vUDsKg90UEqrnvhwLQdVKJs3g3i4863XsCq2GyM90MT+ZBxnzv26HxccHHOKe5UY
/jW1tDNhAmBzvjswklJ5+ElOv6JfBZaEXMjl54yr6Lr4hn7e1JjoLU0pTKFixlxb
SQyjfNUWWed2o73q4FfAMl4o5rRkeHIVaaOr4LfdHLG0AvenlokBZzwwx2ed5yNR
W/eRKKR9ShzmFtCHdKfmxiP/Yge73Mdo+ljGdHpHh5F6pC1znpl9helBvPYxIyh6
DUXazt/oEVsLkn1b7ewWy9Kw3BZkU6xN/oeIlVHXwgT2jjgusYLNKUinv5KMeMsI
zB38FZHVuuPYPbrXBgVsEk1u9mYTkIzAVq5ksXnRIxqNJ1Am3b1QyXKbcVJAy5q8
Gzy8tr1rVyKPJdPrR5sgevZNOYbT6PWkGavvFm2GR/hsWuHQZoEmgCESxEtrWdDJ
x72muh5SN5spJTzqh1zioaG8JNq2Zpmmmn+aVMghE2hPr3QCIThRIiPFU3SX9Jn7
YIA0I6cJ8iuA93r3fqOhbs+StK09tGhDQJbepQmpvNquTrRp3ydxLdq214L5/Lad
kf4yuo/lG6NVy/yUWPO2Q6v5K2wAUJSw32rC3ltDYh9ryVkPTqhy1iYwDgJDgR1b
xf59Bg623m70cS7Eim/hoKmD/M4zaEiHQqPt7VVsmEowKftU4F9tViw1JaV6H2m6
K4BbIYxg/rCxmQ5TN270k5CfX2qXEZIjLruEl5IdgFnI4h1MgXXedjZuod9QklrN
ufwvDaGbc/5n9XR23yWS/3MUWIuU1I0MnUHG6cnwhJkpUvmNH1LmIaQ3s84sXLZJ
hDle6paF08sHB8sKPo0oF/8jkioCI20aGSbb77ZNJQLXAdaJJXFmPEjkjmBG7gVE
pMJ/UgLl0BoquawxrTkHHqSJ53REL2iR437jIslOox56dylXt+LV/VhyYChYj8eT
jlu0SLFPhas52g85ROljXluQqBloHdLT2pA4MsR2Tat6tujyEQrzHWNkqcQJVPYB
G1TDHEnTfm6s5oSVmJe3IkdA+PvUAJLHF58BlZjK3OwWOFUjRyRG27hokOQ2i7S/
oH80qfjasjBT2/6MLnZ56M4SaMAzX2fpERrm37UAomXosFBnDizHlCHso/wzC3rx
VwZ1pTB98GMgJu9S9dJYMdJZ6D3LRcQs69iudE3KPu89fqtRcdmuCnwFKWb8OcG7
q7uFeFBNroUsTRM532Z0APjf/MbAQU3YQfmDdzZgpbr1dwmf5g5p3cC5sul0e96r
FML+S1p/RqzjWDot++gpuOFrDmzAdqv+a8PCJunZQb9RcDf+5wBkJn6Vyu0nSEkP
XovAe3wQ4YVjnfnr1yILmHbp+xcdr+76SEQfw7+P3cmSCVUnbuIk1FB7OBrBnU7M
rtcr47GBkx58ECIBmHQAzY8OAvagTbMPIs5LX2RNdrJp9I5JCQ1YRA9G5nFkNAL0
mx11qqiB0fQK6SWGuyEpt9/gujHTIBUnYyoUqbVix4Tzyld9PvNB6xZfnRx9KEn1
V1RDE3kzkIHPHUXWGtaR4DK/YR6mqZ7K/LoKke9O/EdEiNH2iMu/caQn70k1Z9or
E618qbtqfYzZDKPbtW9LZ1nngzE/9OdfiGXTc5X0mF45N7gTXJG8ugbPnIbHedAg
HEhH/NFmlHmhxLL6JxnKEd+QUJ7UKHb1sDBCldmgZqK5gnbckxwRT6wdtQ6S36CW
LBucvAERrZ+M+/CnR7KcucoWM1vWmpJcvUd4iW8CiaStKkmiokRv2GJJWpxWX3Z7
q+5/0h/cM/b3Z5cinqPnYA/0hQuSWUMy0mSZoTNBYMehnb9Ijkq+3nfw3PoDAHUh
EHa6up73+db2w27OHpF0OmNIViMMXwMOF0JuoA4CtZ0JoYHlDa/f6mdV4jCGKpoO
jMNvCPc0sF6tZ5L/dKVsRhLf7mZ3v7wW2lSslBUQ6MlDvWWVnnYBC8vB2o2Hwso1
MhBD/WYVlU2oNf0xylR1z2PBIJGat+E0ubCcpaUB3t1QgXQBl2bkebEQAM1qdcjd
UuwO9/YPyJFmjdQ4wBeLPvMvIvyLz7AgjEEuFiFfm6+LQzKe6UVH7ywaPuK63cuY
nfxED3GMov597RbIuIRWKJuANstlasApx4X1eEOc1Z4CQ/Hq/O1ruxifLJiSUv9o
BYfRYHp4Ke1FD/TgIssIy1qU4rY3bpCnQM0341MT5es=
`protect end_protected