`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
ETPPCP8WWhaVlDeW0DpQWwLTQOOfTo7PuaZk82hmyE94x9WvgjcmL/iKP+TbI89T
iw6cGZAgMIwZaDJv228gyiF7FfkyRfHf8j7xvtxNTIM+ZVcjqUgE+ShVWSKtfJyO
wHzSc4MLYG8fLfrYzB0Lz9qr+NEBma2VlSb+ukRFEujazpv1/jjt9Gmj5XYE6yhx
DijsNVTf1T8jnBe+utUIQglg9R6lALMsq/m7kKXG079uOYb/lb9v4NJEl+Ar7d5S
JJOyOQGauiIhMm9uTuWMU0GFWJIFKJkrw+8jybBBnYB0/42+MBuhPYj2rLdf8RmT
CcK0iQZgt8o4XPcMfLirhA==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="ZfZ6yIkkjxQuXoHqmsuN08j2CbZACJkyDn2f3hb0HgE="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
I225DGkqmjyudGVZEGAi8GhJx3TEfbJoYUuv2f6QNNNU4B7+g0yqWlWxPiUpaF1F
yeeeiLjrA/W/CbfJe/BRAjjCiPjjLEZFo+Dr5/qBgs+p//3GMnD1XibQhpCK+Ff/
usBbFcrFXD8BvZ/7N8JeHvW6O8CVqlzupQI+oW/cnCk=
`protect rights_digest_method = "sha256"
`protect end_toolblock="uo7KrgMMOIrfLbOlBu3lom43cdWd1MA21jMwUlf/hUQ="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 27696 )
`protect data_block
FpnsH8w5EChbrZleT6Yp34WqH/FPKCznFR2KpeXYgwgHf7+9IndmO2BUAaKHUPf5
5v3u9kbIq1ieMAix4aRcLDZxFOmzBpYYii3LkqrU9JXz1+zHgF4n2s6TEZD4KtuQ
ATkS0e5WlIVeyjNZ91Ns33rjHaSsA0y7vr+AWc5rxPrsUEV+z5bn4ktcJfO44qci
X1cyT6YLNNYAa4XPgl24tcDfZkKmzAdQUoMmLE8SyFaYpuC7s0M4DdaYBB1G71iR
fdOZOR9/Hkce8p2sl6zkWoO27DkdPk6iIxNGI9xOUs6X7IrMdc8rCGnQ+dCp+9h0
DnOGYmDItDntXYQ9e2OyPhF7j7jTJzLYE2WH83KEe1jU59eH4ijt5tAFZKYHN1ma
zkvLM9uCmbDndZH2TIhRNm3RrxcnToXR8oM1CsymccajTYQp5A1UX10MmcPF63Lo
aKYK7S42goKJIIKFEcRDTuhybnSBrjekrnLjHv7i1ETobvseYGd2cFjuDdh4j7RA
RmoxhCnAYk6vCFob7BpHgxlCtiVO0tJpxSmj2BcRIFYT/Xm7sZQB819LuuGClE2H
TlnfhtFadxIytQBgmzWqBo63erS0+Bu0GjU1zsaCYIlH7quCDX3FLNNlx49Nsqv7
zCR3K2U6hxLBMyGG8zg4n+EAGPQvhVa0+IE7q6umW1Giy8OQ52TWvNuoHhk8ZYHz
8fhLr7AR6n7BtdZ7InKczqGKczHAGAnAg4yL912PgCCaYVVUDj34NP/HbSmrUEVI
LyimolKR7c64L+hRtZquho+GRVHGu3O/3TfHweF7V7xbYP0qaSHOId1LvCkmJ5QR
mRNwRicBjlMBd5p/gUt+nRZXyaz0FO3lsiW91dF0DqtZik+F7W7tQ2W1sJsirx9g
C+FSBJTrhdE4eC/jRBNZkGy7cxykOqwQEKJ1W6iHXGS7bcsuBLdl96P48sj9IFM5
fu7Y8r8lWIkpeW+3zHO0Bt8Wmnrdl9lvUA43nmhLBAIX74d8/SeNZRhaR/pFOH9T
nKwQ1TUYLgOoa5ExqquGjZ3MzdDkV90hZyHlb43vdvW7wuyTgZtr5c8vUGeq2BfK
wmm1S77SrbJY5By4uHXTORGmop8MYJn+AxgN/QU/kCNVC1KtS0q9prdGirp0TdQi
LlYpzIoSZn/adY0H+RDgEbO+4nBL9JZ0/2fl40KlJMXQetDg6Nf4cbACr2+BHK4X
C0zdwNB7iXnNoi417P6AYrRKXpNELafzFrRFO+gBfK3/vgq5XgrBj06TjF1fQ0fC
/sLd6fgi9OHI6amX9BYUIF6n9NYTT4BCHycrmC5Z3mMR6cDXL1V4V2uGeCUC3t2S
HLHtvMZuUmQxPVNkEaQ3v/4WPK8suejXiV37hIITMofxg0sfdcIdsjg82LvmV4O5
A/7Inev5g4XzCbnCNDtPCegA1H1Tf3hej2pn9CP8G6Tm04brfhUXuFC9pcAHdABr
gNJ+P7roVBposMTJMpMYuKsMadPl2jWlOl4MvDOl1elCZETf7oO/q8Ce1G/onKfj
jtbAWHP18WxSJqCIGQnfkNUPV816AY1wv1esQsbBamBDY1VBdhctkoYno+cxndwy
kL0U8vPWa6Ndi3IkQJRtNG3LrbyWWVdWCZszvrP2XM8bmyMATP+fFVWGyVO8VpMz
5otESu3ELtCYuc2QxfJ/xe4IH2ZyYef3Xksod3ZrAaDwg2bwso7LQWImVhXhdMLI
EFcEkU+RiU6ZV/PjA7tvVZR7HZ7JXFUBmgEgaqmk/UC9L4LWtuFZ7OekRQjW1vdp
WyaYhepfabo6w6P2cqwXxxkD5Hiimf+OlxWsRRE/QzhvFvJ/EeEvlnb4pwc+lagG
exqBGSG9UmsZbkAqOGjLFUn/V58xZGddBRHu7nL1T0CF9fDkah9T7SIr5yiq8lJ2
XL0u2NQfM1cQbxUD0My8e/d6xCa2rLWROSy2frA7r5x3vo14MXMapTH2ar/Dp1FH
5/cHyhMx9CIZWFYR3v8jdQHFsBiNyPscvA0vDxv4bX35g8bFxJ7jRpImqlEqo0s9
kH0ztlhVpOJQOvJrNpXTmeLcYtLsQeApnMa0Zm67gmfX59eQ7ym7z3acmzm2GkwH
qvAGEh/7agK7rnNEGUJtHX/F2bqb0ZgpxzpCt17po7Q4H408NpA8ZjoXgyclGvN9
KO+neUAmSDR9jorlhcyHion/w1jyweKMihDt+aVt80YgSiyyTjjYcfSTZx+tb09C
1cgvN0IQUifUfH3X90vIc7l8BG0uXxj/aDSXa1Bd6ltqezIIDVrIU8mY10OEltfV
3FPMVqa/pQko1ebRaugYohhZDJsDawdONkTWsMn0ZBn4UNr8yFwhaGZgkG72BNc/
2uKCKWkAqLd+9yFXDAacC+Vg4F4KwmJQJskR61a9HxVAPMXmBTs1VYVawhu1Huwr
0Cj0fJwbCM25ChMZClj9ieOdPqFPsQibmRj8pGOxPCOYEZvZhQj1JpwEscHHcnrY
8GgxeEAWJwUC+Fugz7XJkiqkp+nm2RT2Y3OH3yfy9I4Wl2sKGRc25fBOBos2hdI7
3+X8Ea4Pgra8p1DasBcRA3HH6TZMF3/LNqH51P7wOZuGJI9Sy27S3ar5bqP2tB+R
hfk9q2MTUntQEVwHlznGm12j2qn+cy3innWVUx9137bPO+IO1P1GzAK6+MCwemID
9Mb/oHp7JF8PwuW43YdVk1gum/kq+wSpnPAN0EavWaludRG/9CpPGTY9V1SQS7vb
FB+Xb+sfXmGaSJq/NWAxXbd398stvHiL+m4EwGPM03FmDYaASyEorO+sPD4tEi9D
5/XNBvw0ZnLuaWD/OetwnDXOZf/NuGdz9C1e+hzk8frm/t5FFZ8Eoo3HnY7EyxtV
qHxlePIBQesZZOqvYKJAlUunUvLrD1jNWSX55zhv2xFywUXT7nabkE6QrYcOTT1e
YoJKZww5nLkD7wGSLzsvKhDEWKWQNngKyPSs24m2HYpuYnO5XnmB457G3he0lCC6
/9K8F9DyHMaLLS/4k1JSbPpduxsoP7yRlJhUXc+GozTLpUoFXVBBomDuA5z+f570
oqLYizY2yIF7OhLohlLMawfEGCgyPPNTMvQinyz89za5nqQ340ZhwPrukY/2x5Ei
kzbD4AXIo+ecpAQa6PIV+QJuM1XcLLPGmhAwE0LIfEuhW/7wiPooUsy2UgbXzzCC
rtBGR579gL/tZNWdtj/9NWt3YLMcF3Jnojlom2Hjs5DCuSgulJ2InFHYXd6/AHM1
WHr+WBzRcFlNBAGFehmXCoW9XYqQSGflyb32WMkpOfNHmUCD/eg8rSLY63Jx4c50
sGaQG6wpK0VVCEpvaK8KFhGYsQJL9ysgIP3SJkjyru+huUn/FwvtCuek/wzKJ9kS
2ZHgfRDyw2kea23wvwm2IT3xD7UrAEUGW40Ft7qdowhqUKlole9oxW779SkKphqF
BAhARXjdD43KofrI1f4ifMkUYuU94Qnms7brf3jrcVTJGtwYDwR+pJ4iHNSDn9DF
Z/W75zTaea4QLgKFobahK5Rmdi645vSHxLlYgr119r2IsSGNspm8UAa8UxhrEv+o
4LxWHZ+kqZMUBAXrPHrmbnRtTGz9mGqqMY0dycc+9eSPwqi0bnO22xed+BHhyXPB
JboLwazt/vKO+g4GXi3A339IJqHIKheO5O6aOeN/nvYJ2qzeHnl3ehwPcJSaDa0+
28gq8w5s2n3ElMR83QZ2l7n9jw/EGFzRCYuvpEzt/RIPA6ipEWHuMn3ksSnmM8tT
hUO5nClx+O7uPDQ5zCcIhRJjsy0RCxkouXDicPgmuNZB5apXs02MlHWzOPaoE13v
dRg4U4INsrKjF5En+6mJDhU8gvnjZcie3WylGsyJgoa4RvR1yCFnzy9zlVewqntR
XmRUmb7L4VWJzqJxzC/9Fk3jx0IvU9jej+6vFcemF+ejeTpMAhrfK1Cuhqjgrzfj
G+S9uBPSpRv0ju6T62K78giOo1xKJJRuoroPsuh7ZuFiMd5Yz2xo/L64zAm+Gvxt
AsNHjtz/NEJuhauypQv+qOC8yGRkpV8jcOMlisy+TjZLyHJR9l7p8j7oYoBFBXhs
o7CJc6gYv5CvOKh9048Irg/HxBgBALgLXM97AncVsKHDfd4HttGiLlHVMyGR+q8N
S40cckQkEACOvHf8rNYb1v/sORFSZpxLeF1ca6eRKCdjIG/FMSNa4apapjqG9T6l
Vcs0R8C0bFx+2ay7dmAPxo017A5oScjzu6Jx0BuhHbm9cxU1H5wNrLyke6nyRj+s
qrwxob+7WJSetAWetCvXU02wHUPIii87Khs9f1dVvLx6yjKp9UOvNV3/iRgYLGB6
mqNUbdeu3TAZ1lQPYKasxpxtKf5qY9H4kGBdJdWHhQ3hHCV9xWjkZlzjr2rmqEFc
aYYLl8gyII6y6XL4KG6ANutiisos36rf1OjuXTByC+xkG+o44nyS2nntZQqWePdi
r0SQBtRBse0XRm2/F2L82NEjDvjaj1C9A83RPiDnH3mz92KUrfKN8wsvbTUecBJb
7XqhQJC2ckPlhp9NmDmH0r67ku4QD6+Y+0AxM8DIGS0oXERln9qWIWh21GqC+jZh
40ZrkmC6fRbHuETSDe0njUnX8ooC3lrRVv/b0l6MOcujVUVNB5vEDN/bMc+AFKDp
w+OWfL2MiIpJOzpH9ZKyR0jA4Htf+nz0ktvudzHo4ZZ4y4r+DBn1tW/4KSFb6S3i
h/H3WzrNaD3HgE99SFVW2tORNr2aLbDr1aNlff2kQhmvtGIcjHJoug3NAshcrzMi
Wp/2LK74IjJ787C/tVxnaeN/mMfLyS7zF0uKddTB5GmC5WhDMEHqALWTidzyK5DN
0IpdB1TJ7oqWYBU1ukeSRV6Ic7TR7sKIgFhBvIHgDOHAjVcU8a8GpAVtmNSHa3ho
ZeVViqg6nIyCbPLLhY7l5KdH8bB2CA+1/m8ZgZYucar1fpNnju7Nkpg31GfK+XzA
CrxOziqUQ14rGOdIUeOZYlmgTfrxp5Imv3/KgwDFVCZX4gVj7Hj46NGISSc6qRcQ
MHRKOQtKtza0i+mSnRyyNSFG3HuchlMU/4Eu1gtbA7Ufoj1SW2iQagAxN9QS75GN
aE5yRmsdC72R7lfa5CKbXDsFoUd4hwP7PS2R4MaXYc2AcBLQt3TkQvQ3dq/3pwZZ
RFaNLFdZhjLxyVFgeLpJtmjVN2yu+zoOm9VNX4MzVORrqy8rhfzvO7IxqAsKjs5a
mD10grFgK0pex3UeFMlFmTiqfEoEoUHtlRSDVEJBCzWgxYaV5uTPCN9sYFntQ11l
8LbUYTt+SvjaZ7mvB8t/goqPXvSuRXcMFYcBAqsEvpXTTwGz2TbsIeKI++GIP9xZ
+HINmJv8rvScxapZz0yYB2vb9oUoBU5jcyMGGDTt4Ule4skLtvJTAAfK0/lub/fB
TYxQz5uzQSvHm49N5QZ5gLb8xMR4o2kGj/b9/KSKNIOPNZDOOoWwonXht4P6DCzs
rKAoTWQV0tZi5XoaD+gfZaMdDFLowXRr6+Bno18SoLTtKsJY3cPmSHevKtIc1Yfa
FH1bhzAY9F6W0NkBRL7DA9ga6lCr//7es9qpVE7i2KO9jGmmcqCgvGs2foEyLuHP
A9wbhIQu2oEEt9b7Kr5M45x+1dxDE2eIrj2g5r7ajW4xkDihXAoq+AUFNJnuybAX
9N6SiDsDf3aSOn5q32N9Wa2Ix5GsWjNAgdb4ZkIiYMcAHDSAZ46AZ7o3fAxId1xt
rCIDJx7Be82SezGaChSuqp+wRb9P547XxLs5DZFc7cGA05DLUKkJQnNBtEkZyZhJ
e3WE47eydF9akt7Ux+ujP6VSQBJyRirQt2ByjXw2/Z7Txe587L90P+fSPrHLCQf/
8CLbeVW2/wukZeXAoqBGxodTzCmB1XbuJ/x7pCPb+you6IcjB98V+sUTrSFoos0H
aQtaBu26cSMAqeCgXttDXom5Uz0pPCWD3HghCDJANvmnspo/baruw+7ujAH+j2Ab
iV71nz5hwbeoqFW7gjk+3Bq3d02XUQc66aDwMPnznMOV12Z0l8KcVj4keACvIMOj
Urwfulb9u5JdlE4S7x+NB7unR64Rx3+12/S8Mku6XBZjubLWRxIqF96zxYhqlTmj
8x0AcfiWJKXuIG5BA0whLL/SBdZmeYPk4dyFmZr5f4jsjAGV0TdoB+pyQs6rNQB+
jnwspgcpGgTaYCZzq9LgropwZYrcZT+/lJ6/75iTXZf583i0kFnPi1I+cTA6ZOCa
8lBGjUo7iWzEY6OuG4e9alV/CjAdeF3jsVbyAp4MxUseEECJLvHq5iKKU0wCre0B
+x7JVqadsM52jhYhDPpDjI47bhyGg24orAOQ1fnUvl4jNj/CSD8h/7n7Zbq3gkRd
fm8g6N12o4b78WWMTTjsvBA0JiYaI2TRAOS+GYdtr1snf5U1+DhYtJRr9dPisoQZ
F6fQ1vSe9aBddusvnRnTEDrHzJYYCOs4Ehjj8nrrKdg0pyDctnJt/xCb+epPmFcc
+4byc7r+qtFxci7adO4TpvOeAATyFyYs4/rWBkTXF7RtTcmb4lQH59FmBqDYtjFe
g9fTjHaKhfErpL3ug0ks/uBl5Vc1XbXGWb4FfC3DEfTozREyt4iW6d9yEqv5g7mr
el2TZ66Mo2EVsJ9M45In7S9/2mh9r50z2YA4KT7T2Ce+TBKahriCAm+vYCsg9mLR
tcUK+KRJ5kHEFmIxGAZLMgnSdTaaCyXD1NNqeqhX8MMSV4FPMDgMQbKE7HsN3GIx
Jw0Jdc27UQu2o3+JRM6UVtcCw+AuxEgBRZ5mR/IgRvJlBTQSjo9qEBagkBQGpMKB
3JR7I2YiZ/l/YOBiqZsJeUh6FFcr4okgbGdEFLtNNlWT94vdzLeRG+N2j93B4CDl
FYvtGVsPC0EGTHKTwh5ICzQAi3tX5cNTxgLiwkiF7unygJ7EzGDg3CzNKg7afo+4
KB9ZYPkG8wSyp9CH4fJo7bZIy2TCY0jAXC/j7seLh/fLs8NTnodMYxvdUiM2IzfG
2l+3uI5x52RF1r2iUOLKwkhVcp62P6vCsy7Fz0n7Xw3ungAQX3+gS75KJiPG9LP5
d99ACMufkXg4WE6Gzn0pmM+E68Fg540m0ZXS/CSc4cQAiZk0XAf2nBkwG4u2zQiF
U8l9SKr2lpNmId9Aaq2hOgkY5k3SxS/Du4oHLXgBwNCvyr2gF7FGpK0Rx/2/SrMZ
29uMU+V+IrCbX0xCZ4B2bX4CtrtDtsMS428s/xXdCAUSCqjJo56wrbyUU4cCvWtW
JyGdKkQpOqsTGnurtARYZjJFzoYu8EUntwoHhWE7l1dirDMj5TwDgwP+s8praLxC
FoJWQr7FKjuX0V9Nl+ZW4z9zITwW7Tec37Vd7F623cxKldkdYYObFr7UprU59UQE
PO9zK+f11UUXCeFVIioVsTgcYf7XhSy+g9KPn1qttezw91gPSzWqKjVEUzIkkvZf
BiPgTy8sqbcZA98G5ywQgrrBHfzaJXGEK69AyNao6dMUFYti5kBgIcHX7WlN3cCd
cQZcaXTR6tJFdFQFDyRYgPVxXMMShgunYFUPC7oY64qlr156b4Fnin0yTUhmlemT
8eIckh5PwlSnb+4VzS/rII0ise5ANfw+PY6/B2jCIFDok/S0ym4oTh68IRrD4nCZ
Z6tIZ1Jg+aCyZ6mzWeFsWOgY/R/p7oELdwIKkfj/gxnKsbrVhr5aQafQJJBdtvvO
FPtg286Fik7DP0/w0PtVnMz/sjLo8yDVwDQOFKKZ/jUzm/PdUFy+g8RdiSiPxQ9n
hM6jeSvGKM1yEMit3Kd1Nl4y4956JL4DdZcBlwE7KaJVrBNQodCAErp2hzVFA08N
u92b0Ld0oR3IwpblE0MmCS1GBs1AgqEdUujIQ8JlthLazWZ2x/9dWv0QWipHH0Ni
iOashTX9cL8vb8+8vxrrSeC5mKCKdn+wUKhxHgpwQYIyNaeKJvtLCa9WXrU70dZL
hhYcDVxgOReBSQPKQshSQpuhq21NRgbLvDAOj4bVcwzTPpjtNZvwGAQZ51sDWrHK
Xx+PTAG14bVhiWNVMOpMRxjiRFGAAvy6732iiwHuLUTyWDjUu0nEiD7ZqjIxb6Hx
nJ/+o9YDDMdnhQT0A5OV2hHSidlD3WXg5Dy84i3c0m+x5A89Burv3cItMcf8INHT
XzaLghKUGpur41cDy9XgougrN7BNks5HIfLc9B3eM9lOEFgvyqbeGC5KH2/OomOU
8sB3T9ADCwjWyayM4SIomsSP5hWhEKsE6uXYY6JCsSjl3AcqAlGez1Ibew/97MPb
W7ZXXobTnKJK5DCurACrgANlKSjUMqH3Xn1doQjLg22T/eaJZuh835fpBLyFRPu+
J1DAc5E2718ZlBEBplbDiDLcGbHpFcSgmnLC/yNiWxvzj8JICPcfER1zUu56KaQT
UqH7xyFOM2+mhgEK88qNY6p8r8KdjyFZVf9S78cbPVH/DU/4WyEfNR7muvMQjUGS
hidQcGR8Ea4qN+ctsvrFP0mEt+3q0ce1lMA9u5pfNdrqRnCZpx9Ds37T88U0hOhc
FQOM2BOMNbDM4AP8XBsrCG2GNS4OYcOZ6yL/Po6KLeT1yRbFUx3MO3YTAdUrN96P
IulqheRw10JqLi2HGQK2zFEZg+869K3BkLk//TdkSB7pbx9FMU2FTyHDQ4WyDVkP
prB+2jH9bzsx1VtEdr3aMsQxhBLjlxO24zaOQjUHmTz2iSoNXFOn+os8813oz+k2
5AC15GMfaG9Zru8TScZ9T+dFwg+aiB2tk3dtl/4S4NWgkif0xFezdPcJdWIv0QHZ
C/hqEqycFWn+zYwuuWjAo+kJNJZE3hqEYgqnqibK78f+k371gusgYxTPSA45SV7+
8LxE7wBwdmo/A4CjVDxBmV+qFy0zOfgTFzMmqGzOahnPBa25jTFt8cSG0dnIliPX
gMbpddvypouiVNnHz4dmmV0x8pBiUx5iBOQzDkroN5DAi9bzcrbqQjcPbYUwoUR1
5VniS03c3XMGInwEma0EUccgLMwM+3NvtVaN7Qo/JBjWW2BGkItO76hPun6rQt3P
LMdFw1gQs/hOiRfwlotgs2fKqIBxwhu0GRwJod32du3T/PP++ePK3DtkU7U396g7
i0Q2+id1zV6bDvEqST46ELCb4zAms3eV49vUpO8M4GYDXQTpbyvvrVxkj+o9mYV/
pRKdXdr7Z5mU6FSMYgDQjNZoFJ83JpcF0N5Sn4l6A0maVrcoo25JtOiIv2pwUKxy
/jd/HXeIMo4ekJFnLvo2C06c2kHNmVRHg/VA50kY0Zy1kBtH1DIh9vaIsoqMTa1w
wA+cDxThvXk3RsMQQbSkFbXpLt42H0lUmuDgwQYvmfP9iLvmKxKg+xkrYfGUV0gx
NsGfb1Q49jHT+cAwE5L94F85jKnQGQEgfk6AxfnM6jLogEPrgOAZbllKwATfvcZQ
hLF9Yo8HpOhBXbdoZpqvRHtzM8BzVtzb08qZa1H94QmqSwTF76HXZwmOG6LoMEZN
QIiqs7YZ5qrbkS0w6L1KZLIiUvZ+7ARTcH/VotbBY8kp5nEmw+ix/bRT7dDbz5yT
V9IZabuo61njzGt567dYa+P5VwRVBUqCTDbGBMF3buAYb+0WtJ5fzDVR1KQWfz9y
5D+Ks7ObHXyFPDSGwVmNkEo6melsIvA1DgziyvWMgs1tWH2vQ0H0NIS+tBUT5NZJ
96hreRKxJMU20sbqd5hrkX6jixfqpQUaBdmWtnRcAscIv8sG5g9uRFw1AjAa5yMV
a8HmE0y+a6D6R7Dnk/vFug3svWvLAV/bfW2g1QYdpCWvIF8aE6Ez4fO/+ttWgCN6
Nf/FjNh088796nCkKcgc5reo+GYnDzwV1LQ3/cvHWUxIUDKBMMsnRkS/LOIKA1tH
jcR5QWE0XkfILHzAN2kEGdo3//9GJxp60M0wjO2rKRVxDh6J2lZP96mbXR3nrtUJ
upj9JwN3U1Xr35HOFizXCo89XJibvh6KLdX+ivZs7CU9aByG+mAiICHL2pQyCOlc
3+KPywfk13tMuY9htfNQRN/CoKEqBoBBl8sVBDWIdPDQs0Pk7hb3ksQ4in15v0nK
L7gkkOgLDEx8b5KBizFAik1OgOMEy2jZEdJ///BRTod85rOXmZ98qgTJaBc/X+bF
SpWY3JiABIkTf9aCrzspFtedhGIm62yXmAry0FIdOySGKgvHMjXvHmTyWX934Mht
MUL9R9pYd3zG+S004AVcA8+2C2qQnu3n5k0u9K79Wc5y4rr21Eia46QCunPXmBSJ
wkJZNJxPmRzAsKNb7dwFccmgbZaFFaZaFGfgEnXJZ+8DoZPi7sc1iJ6jPW8jHsyw
hxnH8cDt31HX4tFxtmiMToXZPfSSegQVVdnXls0L3CyA3+V8e49vx3B9+NOQWE3P
1/DKR5SwrSqFTs4oCn1DEUym//AjOp9DNh56hJ5SLabzoUrlSKztwWZEvthHFXbS
t7LAReluakn8yOtGkBBGhKbn4yOCC+rqRQUPXGrftOxzrgmUx7Ws8XUUZuPTrEJS
zvVz6U7/gEix5HEkpuDKlxKq8fs1AwkeTi/KBh8IGhjOy7SUIJpPTb0waWvc1I3I
leMtCDrNp59z9lA80UFJL2E0SISMr57hLNVpPbKCabHKJN6460ldHlKheaBHbjY6
XLJBszprMQzwnXNpZXjdOojXmao1ERV9zcKg0qCW3WvyiB4Zm5A8fiB65AwAhzMm
K51qU0SVBJQG944LwisbTei/VfektmN8c3DgseWsRkL9jnrBd4yiyvJ4wfCej+JT
VaI1Z9GL2f7wcmb8ZmoMzb5astfVbqcf309EYjP1uteIagHRTVzKblXdETd3vxft
L1qIx0J7WTpm9vLCaXSPafk5xxlegwK2PXzzHj05kaZ1xXq4TnGA6EYsPuQnvMOq
WXMhOOWsL4NcellpZfdXafBT9HQC4iz1naSGEJYp/aTdr5Tk4S4AUoyfkVQx0929
+dJvjh2+vXTiZjH1MrXJTsJYVGHk1q/jJ3h7aNjBlaJNXhZ1BDJu28tC3oTFppf4
ZzqxLHKah4zAbi1+BakJjZdzfY/Ogd09c3sfABG7P217mQ8WmN0GZgSWfYlq/Sqq
IMV9OWF/6TeNUPt3EtqbIMbDz5XqtP3YnwvRkiyYe2N1PpGogqtMzuDdcYYzgztH
+tzeeQ/1ZBGi90wCpvlMw9z94Osefyk3IsoqMyJICcboMVjFozdpYxS0toSq10ql
yRVmA4K4mxgj44g9i28LlhPKXERsG8+l8+8zPvAnnJrPWrdgihF6HmeVn4VmUbr1
/CPU1TkzC2H/bJfcEIuHqv+041cUrQ/u90DTRm7qmN/cvtiDCWxL/5GkaXG1XPX0
7MV36Ss2+0WSimpVOiNNu2ZCBgjPLueBgYuoICLmWLF54skrAnV6KcRLSv3EZgGD
cajuVENeSzGZ2zxqaMAasx49280epqnrSnoWlFvnng837xDNbH+yVwrvlufsP5KG
OXx2G7LSj2RgkvMJp7zSXXIgfERBGR22eQPKXjJhBENo1ypJuqIaIebkD8715m+L
bC5GIsL8CUahhjXh+GwgshUaC3JPmu+MEqBRSUYuQM8JCK9IcEhx3/kUE7MZVKUB
0tDJnQmYDYC+N6I0FTpeNiYPlx2iNf1WwkzPUPbF6EiRCXJLXhlASK+uKkEg2krf
vNPeii31p1Zj5d67vAqolYxQGYhrPeCMqFi25DxNPTKxyMbI3Xa27IbglsRAmT56
vtEdDVGf+CEwJ4nUcwoypn9Sbr3uiQXK7CgjcikYthIl+0Tzvn+WvmkRqT0WpYF2
tUvpEKw4qbKb7V47b/Lmo3GvVID0p39tSzSG+mZrvA5vJw5XRB9WYVCbc+Lpyilx
r2HKGGpLp4p/fGg2L2VWBINfrel7I+9XnPQemm3Y6+UlBp00gdBRHkuYak/jDiFg
pfHJghZlWOFhdhIyRPQTq9BiJSjTRxuzJuIfRr9/fbMv8kC1rTi9ye1lsMjmhShZ
7v4nlVVA8xjXGbbsLwNVz0MQ7SNxaWYRHjELOF70mZeFx1bZv6y3vyBqUpR71G7R
BNF0MrHr/ZTgB1DqyUdFcaD3TWmHXZBTD9ZSAFtb99jpsuAPChf4PI0KPWWJTfcM
xWK9Hb8Caj7bDJH6ZiaWbjZ3AnsukOyPtPtLYk6Hs6n9GY2FyLs98mWZEh9c8feI
XbUFx/Ny2+gjRvyFviiV7eucSFc7wVM7v+AkR1rN6orpgjqqZic+09zHDol1woEq
vQ82Ty64B430vf2ozawA/dXDuQxgCHxbCyZBSbxUu1iQ7Rr1pPK4Y/uvGHvn+Pgf
qcQLazsxUkmF4yn3V5L0KwDxim+F4pV63Tky6Vl4ZA9vhQN1V+ElwYvCYuJQM+Ug
5SOaNrlZm03tjYQzp03KnJ2gnEQhjLhcEseZdILhnpVUwIq9F11d2H7LgeExObZx
XhgTldOj0qRN7l6qru5gL4M7IFMHGXVxTWycFg4L4IU75F4jiX2D0vU892XjOuex
73snEr2GC4DbsmGpFWJWEqPbfRoYY17FFR2xKA57+v77OQGG2gp3UXLPta3ZWt9b
v3eQ1XubwMxqk+n5omZ9WS3qVAnOxz3G4hcsXepcTY/h0ceAb3SFJitAnk/HQDDy
FVbts0LmWcYw92eCfu6PXqq5rrCig1/ZVuzazGVBqOZ3hiVJvHh2Hu44po4gUhGj
QawxT8Fd6MqObd3mJeBUt+sC2wLX8k1CcC/v2VjKik7PRueIXFsN3fBDLr93+Xt8
zE+zGMzxeca1CCFdp7ycQeg4oG+m/ryewAtugnX7VMWSeeM1KuMGV0PfxHCxJ6Ds
XhpesfZjdYn57DzChnmnQj/JwiQztcPd7nYclSp4sPW/RTuVkoJIRbB10+rot0nr
5cfNpehW4opY/88hklJLDoRZfCJC6cXTiwkyTV2ukvPwhQ12kt0onjBF0Th8wr/z
btxc4ehjj13Qh7JqnaXV5XJgCX8DMyTwcGUPZn5bwgVBOLi/1FBr/ewwfd5NAjsf
YW4c0J+YQcGLw+308tf9N+Ohsg/Xyud/ArV/s9Mg4Uc9vPM6k9e6HxEfhbhEKL0b
uWFkNvmt3hV5/2Uz143kS/SmpqMmPDWFd+cZp9KxppsuLx93mwfyVXHaKBKrhgLf
Kkc5KjaoL/SsXvicOYP5/IlUiptUcHiGQBvWRSC7PLzJFniCfwmFz/E3t7V33w6i
QxyLdf3T1MxoS2piutN9di/MUqUf7FcK6nsvYS5ZK4U3oRMn8rc62aHiHiXpBpyF
R+F4Gnny2omm/vHzTSw4yCXII4uDUmMVgXGqIl0ZqTfeg5Xlgid9hV3fS5AMKrU+
2UHN32kXN2kEWvzXe6tvSontdND5gLJjNk7MaIOEhGPIKhcNv+DSWuvUCr7mJ7km
swNTGPqTAryVbyqX4pgYKzvDaDiK7poQeayxPiHLSXTu/vSBIs8yiP3EcFBJd9lF
6Gd0AG7c2mSHsh1Qr11sTPfzNrqtAsx0L7oeOHQ7nNYGLiZ4vGCkPMFK1GjZ0V65
XQCyLOVQkuVW2+DCeChF35qf1cfYIlis/WJ1XH3ngB8OhEfiCORWxVKFfd4oXzjZ
4rVFjW9pylH2Fdod1CMG5hlT/eHMhBwDiXxq8ADw4HvjqM61daylnpVreu0ZWaXD
OBb4eGookTg6YD3AYT07jKRgfhxEX3CH0cuKLWphHEH5GxqjMCtaZIbFJirrC/1u
MMsu8oPtciXz/5hxN5hyKM0iyo1h6cYAGYQnEJa5DhgxXKXXn8YFV9fXXs8ytMRa
RF/vnUH8npPr8pbFPfnGXeJuAt/6t/NaE1XAacxIHdI6PRm2xckUdpaOkyY+fD1G
jYdv2gviSTiHV/KpPlpYXj6B4+IPEfTX2jv4w4J9x0TaEZXskq6gIjaiRJnwNxOd
d+ImU3lf1YTI3HhCvjAAc+ToIA7ewMotVPSHsUfuutiWXv1NF1QKsd3FbY3AcDff
Ms7TIKSCySLBQt3YwX2Nc2LC2UFP9XvHJkxIJrckui29ErI3uongWgP22fE5pTWB
FsMmMxOexaME5NvgxrAH8J42PsmnRiaa6Qq50oB0cpg8eYgFzUZpQ2++kv6SVGAD
8sW7lQezB+qJVRt+uUgeVpbyyU6UN+H0ga1113qaqF5F0bP4HumLPdNDm50M3Vzl
ED253N66vDtHMaEwQR+gya+9HEa83SPJEvRlLJHOVi2gfPfJdisdAaiZPJwmu0BY
rEOuXeKVuh5+N77YkNQ720yep63Nr04Svl0ag6M6gXr6T43msyhPCH/W0s0YHH2v
eenmDbgdIq24HAFSgnMQqoAQUdnKLnD6sVxmOGFVH2YXh1gjjwRatqB17tsfAaWb
sspPi6AfhVehxoHT5iVEqn7cxfOeW3q3/KlCPhTFznWFnPH9qSqCOhagHnbLA1U0
c6vaAxl8/zQ9WN7HK41AkCGBUq3GwkbSXbTQ+OMjtxt/pZG1GfzE0fqt6qTmrpoU
T3kmpq4xfasXrzqo0o/pfh+dPsHX+JkFYLJoZZGcZRq81UXKnL5D5VP+d7j/RTPO
JIEqDqk+KidnzS1e0OtYmRCaBGOLqliEUUXi7Y5N6CvLphaH//7J4XfXWx9Otnix
dsGGcURhGG2CJ95P2pyvsCV4+i0wlCNXqd+BaBZtGANky8pVaSLpvmGC5YvRGL3b
SDDsMqJtPT41FNyNeobi4C/fWrZs984YYe7chhd818ZEDInisve1YYJMiXqZNxov
7z8Vmn2npYR4ePPT2Otc1kqFgeAQLlNu/npKqEIVJPSoNxaCJMLTyZZ+0ykYu9qG
xJu9fKd6X3TSrXZcoKqpTXGy+QnxgguXxRNVABa5bxZpSUi4WH6ZOCTNmcZQ3P2f
fahrSaBbP9tviKvpjDSMyY/mXewXmgfTuFRWrLpyXA5Gk7oegnDblmRdVDtyoWge
MoU45sIgdAqU5vGdy42oMKgNjTPGtvAseAjuOF6sAeeyMU2d13bJ227g1UILiQKi
aTFapYGQOfjuR5dy3mvEQh+7X2cv/+6uxWMT4JAys/tuvWTH3RMgs5VfwVjaq4z/
Vx5H8Q3Z0e2WoFTb2OHIRO2m3tFX9Tektv83/9TXu+Ga0NnF8d2OzQDfMgqX+/TK
dSdoBhogqz/mKVKrpowEJDg7nWchqsNF0W2oOV3OMq+X0O71U3yO7w69WnoEIUq3
u2uwPUaeCnRgoSjJmnCd5qgs0mtrGsGjBb9ypCC2q4QcY1LS/nIsXlXQncwpLpZX
4LENfUd/SfB3XWvgM46qqr/UZ/iXJYe1H/l6XcZWuajR0YNo8O1kWOyyQELr6sGG
/NJCoy1BdIaRinxVmsYa2Hye/rSpVSTLIFoLLtDmi9K5B5+ocv4O4vktMhm+5E5d
n+heU0bbHD73hHSIek9cTFaqF38+PZAhs3hd7PkNAp4iBkvFzhcH6+gVMFeV3QYl
CLYzo3qSdl20jf3ZsvH6PvEUkwSL6pluN5YZwPAm9biUtZ91Aqv5VKbQGZZHfsLZ
VrUZjaNcROWMdisLQfPLrwfaiszcM1AF79SMb8Ks0Z2L8zAK3yidN9yULaZ03T9v
Feh1il/VMZ41PiZCqttCFp1SZXtxTQnryFgraGZH4vm6wTu1A26xaQCDenzAmyfX
Q1jTIlcMvDr7aTSCkPf2ME6oJrHES5r/v75R1J7B7MwFjRJScuIHmR6Fa8VsrTcJ
EEKZpxOxBKYBv70diRBPs1KiApA6dfmZu38lDA/uTRN6mVVRsEq3q1VzaDsWLRy4
NtPWLK0YJtroRv/mg24qYbhMEtQQX+oJRU1xp6/N9Rv2K/VexxPGO8udjhx/TAOD
HUqVUheSbPpqA/WwSPiCVpSyqSyFk5eI6WLz8AClIsCJiQnWYl6jsBvZflzlM7Xc
Zm7kBhAR31TcLQOOOVjg97HYf/et1J+wzhccXFRhJxtsHU71k+GWOobL3Exsl1Go
Q0IALkOG45oqnvlzGrETDAvoNo9IyJaqyDI30J24dINwmS44HU0/XgvsSiYTTvl8
oepdb0rUIBORB1OqXRTP9dXVbxjDQ3x3l9rg/eTM4lhfi33JhOndVtE5FP0Tph7M
2D61uRN+L2QPktkMdssKERxb/qBSq0vSmX0gwC+QxkElQDUuOWcfyPlb6ycoiBb6
Ci1YbbWN98TmQh9wV8zxzVnv8FOklLegTF5vIu1wb11ponidRlDe2G9PuRVeD9fn
Vxg70N4oqweNhtDyxb0DJ8ek6geU2d5gn1Q397NPZ/7NqX+qNfXSMldqyg4FiYqK
75ZJboUihJSLfdzejGyHaSeINkFlbdAIrR5zV7L7RUXatd148wLhYbWtOaqAfLao
J5PPuidRndkN1TU7l6l4A0JFnEnbVpYEgMdkagNzB8hphvQe1Ax4IKGEQhSlDccH
EMoye9yHPDG9Wv1aQXb8V2QWaIpGCAS//Tx8/BdAU4MjePJYMZQ/V8WzH8Pw/fS4
e1gaZQjIVU5Pbcv5oSWUCPqgKShPV0EIhG3FomGTEeeJii+0eoQB0cGRscyGzDWV
aJEuk/SO6XjWJwSz7iVuDXJzexzvgVXYek7ByJhMxcDVhColtUyt6pDlNrs7AZjd
GN4v6cGU5VydByWS2QpoXZ0MsxS/bJ2HxnmNoXjtkiZqPvZ3uJuQRPl+/XbRj+Ir
LSzmbhgCfctnbbsdaJQzB+w5YB3H0Uc8AY3TZu6fo3inJ4gYTOjFZwn9zt6ArXLu
aYgmq5vHTXautB3O/hokxkISOVpkm1miP9wQuSt0wOJciWgnfuRAFGYvXZu5VfL0
GvApNtWs+4GN5SwbcAwzZt5gZdi63FwUTMbnPyOwv0gnPVo1zWLJad9+115GoVli
20vKFvXUoeNnoWE/g9UYFejnV7a6GXxyLew2+uVLzwWyfgJInexzavZ+iuEZYNHt
JvWt1+vmg42Sq1xl9UDnyl3v5hdosWJnnsmKdi6RsLICehVqeY2nGCyeLY35pSTe
h11XVU5KyNooPqAh7vj73YxVsSWrbk4GvnoMF2xtLye+oHnsJ29A80cCzvOsmg4Z
v8X1/Wuf6MEmbI9OkAnaaPmQwnom22TLsq5s4BhC4ZdeonyyCf/UMU1Cw7pijDGi
XAWdRF859tvjjTpWh9SSpNTxQML/9JKbjAsAfQqQKtV+RK3MEzxXV7cXM7MZX0ub
SLkGTavFx2kE5lEfAfqWdAfWww+M+C1kNCwo017vIKLVh8C/NKQ2VAEf0ZRyWYcO
qeAO0WBpi3V6NUD0WtumYeaETF1f8z3836NJVWbzdF69kbq16Zm6oOrbVfQ7HYWS
5Xf0QcsK0ze3iTnczi0bhYqq6jwF4JL7bNduHgrLAs4hd5SZN4M4mJp0QR7Iz6wL
55R4z/d/4tpK4TlJ9OBvuCLSnLqW8BlXY762xwXtXYDnuumbZmacwHClogFimTQt
0R+PG9whFIrErDw7WwDJMzhAUsyUHTx2lGTfaRxKyYn8oBctzybsdsl/7q7HR1eU
rPivOCxIURk9QWDzjif51TCroIT8ewa52vVJFRE9N6fcT9C/M5+9gSePFz6PPfJJ
/vvyljj58bAbJYL8i4kecaQOG1kM+Tr3nTKRL/F+1OxsyYe3gI2a01hPvoOxTPYB
AfaK0iplo5fmzf3igxfzj3BtlTraG8CHhX4q0z98xl2rrgW12K5W1UIIgTZ3YgAj
FPT0us/1Nl8Hejje7H0sOJfUl5PtfwdG+V+NRU7ESG4/dDCwv2iTLZUDgZ5Kl9b5
e+ETzScBedamW3uhjSYtv+0n0nNxmCUcih49NG55s3hVJgC0YNMVHNkkFqtvXU7b
doKD6EJZwvyxZaiGpGUEuiJCz6+G+7KunbRjtaBbnw9d5j8vSAeF6D5XwnxMlPqw
n8mAsnJvsZDw3gLDo49mvXQmqVnvIyJ0sxEtIc9HYcFi1xBDe7OGFRCqZyOgnSjF
2lurHR2DtN82Dgm8gTu9peWeIeoNfdwgKwZft2dRBcHB4FlrHBkkytcng+vaMNTI
tQyjTXu3NncE6uPZ4Km1G4j/42CLX032X97Mfw8TtucZmJxIJXw8BT3XKVkTyOek
pyKVCFTCEtuiX7l2DVEhux7ZMNOa9Nn+zGEvRhy27Zs4wMpba2w5g/otXQyQmWpN
6hSyagA2qyoApk41vey8AfSIXRSVguFVKjmKo/pKczpcGdiF/C1iUKLgGcUGM8Bn
EWyrjxuDSQTjde4/KpFvQXlmEfApuFxQ+dxyU8QyBAQ2nfewsc7LpgmGCK2qe0G1
yYgT+dvJh4tEYlRgCk/fUoSVapQSmo60GkmgrF/atScNQu0+odgXw6jElKJjj3nK
OME6FJCumKqMGGaXu6/fcGVzO9vfUY07I2lNWxHZ2cABy4rI0zY6gj8Jz8bq16jc
Op1zaCb1AnZkkDXo2t7FTn3IutzD2GXErMZ3mXeWPAp6L6+Nk8g/IwH/O07MBSLh
IT1EuH88WRaaKmTV1ZlAAYNPFDIP9Za6HCUdq0WNndAdZYWFndbJVM4dW9z1X0W9
Xw8Yn3Hxkbnfwjml2E/kyzVaShQ7u1XGBeYNg7G7BDItwnobV0fdSjkzVwFkiuQz
Yw/nfT5J0Haq9SHebyiRB0NdETDq9albhFdTiJ6ehSawaEDCdWfnsq7x5CPGBJPx
HObVdEDCImhK/7Gw4z0kMkKAVb9S9Y5Hy/QnDfrEPmqpN5k7QG8jTN3DuaJ57wO6
8CgiTNRmZVfIV4SAYUrhGy7kYny2ntBO4abtvaBdiTAXVsSrPCjFgYdGS2+CxPJi
kxffLFEXqfllEvIte9CyUUl6kwqXjZ9h2VQJieEvSxjBi3A87c3CIMiNAFXHAk9d
E0f1iiyC+B18O9CYcVDxP9FF2rtsqJeH+9Xx7RajQrGeOou/NqtMuY/xtrlVgiTf
Beqlb8WTkUU6+xZoSQT8WJr8v6Szg6s1XEg6w/7j0UQ4SXnOYpsFHe2aV0GP4Fyc
Ckx71ERj52Ex4wgIRQXs2xs2d507VGvLEXY8XywXYMeiB09pe2Gk/kyfmsG7g9tu
y8zLCdI60ICizU+j/a5cDUJ/XkqLqkVO8YAm3ycc2vQw8RWSoVPZVkdqXpBx2wd6
aRcZmFeGtzRL1iw1Oo6IBCTcqlh91GS8km2ndciCVcfULOveplxHnTl7V+2m+5UX
WC2WQfF6N+Mx+73NX7H8eKg/uYqY9i8Gbq3fbjqi3A3xLZOQzr9gwG0GxL2S2bqh
YTQAUwipCyTN9tLaFovSWw/tg0A++xhCwwQkt8/NbSmGLWIzCb+4wUPtods/j4P3
MyQacCvDEl/QF27FgQpekoFwJaQtKcVy7K+LLY7aU/dnDZyNHpl+nGyLUlPhX/MK
M4TGhtxLlMbVpyOz2cPq6Hl0gm7Vi2qPmnZlgSiC1l4QEkJTFgfEuxzkAMbNaUMB
eEfUgsKEwBltL6uE1sXnbQ4w8KHDj0XanqcxNiVsSXyJ2l0s6sliwBj2mlU9lNzi
ghwSz5DCKQRxpIi0Y08WrL6HkNCw6TwHnSjEEtyHHh5x6m8jwszFiA41ygftJ6Oi
yrw/EDM8zGSfKe2qiLgXXpLiaWqqqQrv+MOUuKNkqoeNoEvvO570GKqkwWL/K9sU
LEQ6su93Mns479yizQF0mNoGgE6QsJWVrA52sP23Ed6vQJk83hgPPTf4hMpnWClr
XiAzFTpqdOlKsI6N4znW2OYExV7o6+nz2y4vd50VJ4IvzEXuXAGH1DEqk5PFi86c
OUCYtXAXgggPzr+ao6n+ehsPtTx6bzwggb5VmNyPw6XXslOybUIL6sQiXECHyO1V
m8sYpE3qdGsQof4L8RPZCSc1E+BZ0CjhGxlcIF2r941wh81xpqMvyWPQfXcRYfic
9E2g/uoCoNhNC8xHPaykkuvIraAQ7mIhWxxEz5IzVI8TqTztU1er4EzPxYHq+IXv
xOmkPg1P6rJRGvR1f4/lAfRxXilBcCFhO9QPAPvCGzr1z7ndpLYdHMXHadyzSUao
a4Za9Hwi/BoW1umZn+aF2oWN6YMNIA97K4EoHeUosE602D1NHG+aDanDooXkmyME
e9sAzz4HIN6Pey8CNAa9/VYkI7ERXOCO0QrsGy8ZVlXmnQPhk6qsSoBJ97HVGCQ0
5rl17VFRKx8MM061S5hvu6X3M1BDyF7pStbxV0mulyvP+Qrg5+jJE4fm6KKCJ5o4
0+9t1lKwGGLhx+6SB/auODjW95RT2H7WK9KNopdJf3BPDYeeolUsODbYy0zAxeKw
YANNCdqu04fpKnDyuVLfyokkMt1xk/cpB2jX41seFTcD+8PzR3UOiapByWtLuTeq
vDuVWsnpZzsNeuh9r0naZCLpcm9iyOLi9hANcMMrc/8SbjUUlzoU8vhmL3u+soK0
r+uVj3/fcv4zdSzNK+fGbdLEQc9X+QD1V4RgeG6+7QQqrNVqPZYTv77b0pvCIw9u
BzGdb+ta1xh+d/Y61KWS2KOoXpTZjv8jNwa1Skq3SkUzzHCT+AGdAdlKqgR10/Dz
WGVcRJ5EbrZL1Ny8sDkERi3/juoNl2Q5dN/NxKwjIdDhzUZUKG2E5XKbJ6h0qajm
cxy2dna8ucM60cpu5aezz8mJtcEs4FOIDF4sUnFDT68hx4wSNud+/d3mD87MjCbe
xgWrVtgWWNFjYtUGM4a/n7ziyjtC6u9uwWCUq7FJ50+J4WpPLtNS+Fe0u9adDX6O
ba0GZSy4+2n8ZIbZ487mWzk8ITkOR2SfZl6KAKsWGYpi6VdgI8yXXockDXvO+qy7
PltnT6kqHmyFYfpazoV28eBR6Q7+SKH0XuJI3H9ryoRXLeFbpMEqM/YNQIpM56H8
y8bw7skD1+Cto2Hu+L0NhT4I72/krnjeoEVzEnOQM5We9uQMqpDTCb7kqwqYbKCo
AO1yYk58hjEZ2VaHeGOQ9Ge31tywMThzRZ0rADUKSkIi93aPbofxrLnGRouJe/bg
PC2W1RsRdTly7PYITduvl42ATwZ5hRXvdyUSXSCTNIV278lAsGeVcqa6Yd4aLVGe
s+h70wSKMdEhpfZ+BZTLYiJvSkmM0px6QA9TF24vyP+VXDxiS97te55TbdhlKW2K
dpsxUPIsf1aAGVAZozPhm342v5FlzTfMJRirelbPU6We0oTJFYrKACntHcPinKDA
2CuuvF0Y2kat2L86ap0PfjfrNcSYBNfZPFCXgZio+5+P9CyIDkr5KoXBfugabcBV
qWzY38s+7C+6JaCZVRFiFyaN5Rpi6tlQP1BpCYOgYLwbBARMTRAcC1g+I3nO5LNb
y+9bRdYgMzwgnxctt4p3XGdJj8HOQyBddr0vwB794EVukSHIkiXjRSm5Xyae0CaK
cM4Pbjokv5OKcjpOjRwNrxChwKi4gHeXGtdFGbhjR6FyDnrCa5WmQcHjIlZI5rUT
U2+9gQ6P26wY5hDHyi0sG3TUiMLVNi5TkjwPdwAxOV3l3uWwG9BRCybOeuUkLLm2
tbzUIX+a4Fa/ZpGK1YzM2VyAaTIGm7efK7Nfj3Me7b7uuQ/no7R3muqVPaGjIT18
+OxX945xD4F150dgVDlPX0BoiVseA7Pb4ZpXAiOHSQo4CUFi5+Y6XKZEn0NXpMK9
CUmOxKRl7vBLMhUlsnAOpmjbORxbYSlC6XKl44WpmVrKnxvP9z5akPWVsoy1Kd2X
WusiX5193+BUM5oUwSznqu19tmbraMuQrA0aWD789IIEFOAwAF7Inc0Jc7PdANgU
MDdr86zmJfJU7bbTWRUtuCGZhGw9L8UUWH2vL9ubZQTidL5VRnxvOV/hnl7YI1BO
7gmtWDEbXb21GvbtImf6j7Ac5Gd49rMk8D8H6iFzjFycmn4jEOKPgucMMRcK0kI+
BiESqUqE1M/gwJs6+5rvh0+wBHhEaEnmm5ZRqQWRz+8j+8s9lGhWIQoIYmVz8nHx
qrgG2tQsPtNfbnrr8PgYTEdawETzqUjX4Uc+OwOqiEUIzTbT/2YrfvuTUu92GCIt
rLq5Ir+kPx1ATncixhP7WMHV5JUhN3pYROjYPZwyYNQWTmMude9HGPnvNqQVj8lz
ygmPGZ0A70gZisb4LiP4IwDWy16ShE9ZbcEX+Le8IT66Gd1XxvexnzXkHeSmYhRt
i3Tv9x11h4kKRRGKWyC0OnmEEsuxCE689t+RvK3QOAJJAZHrdqWTMlRePiDezN2I
L40rFOrY7hrn8u7/Oaow+v/TVsSsEwBNm/D5C4hdRUdWgLcg2UkEmeB/sOfd6oea
U/gjt2nUQd6B4QVUAJitLHsvWTHhhhxtXKXMIaWkgk0nH8R2lbg9ga8J9wIWC8+Z
hSEWI4ZZHWK8eopr/A75URvuaL4iSL4qOr/yMkiAWJw+oah5kDSX7ULyqu0mnnVI
rm3US8mFhP2yhfpM29Vk4iv1ZYpeCPos1GjAeJ2AO6NZlDJvMApuniPDKfIWHea/
ZFqQye2hCjFjr92RP7ZqXg4V8BmSvCS8ZxsT7/qMT7AnvLY6XAuejwTn85N5UFVe
mAjGL1XCLDLNs0DXd/UwldxINtSk8DSBnImsza1aafU44esp494YjKSR+cgtM5NN
TNPJxcHGa4hBNUr247imf7vEBrq1zqlEb0ganPeiLAHLWDARSVqn1VJB7SaKJwFd
YqtLcSrmnUIDs5KDAfjR3oK6VTnp+P8o31BqW5T0jdXj6sT57Ds0NOgZYmeMxmTr
Uq8ecX2bYADqmO/kjOYkx3HSVnjehE+5zl+kyuIr5j9aVb8HK8rm7gLxmolMC11s
8wp5uRxXtLubBNoKn0iwQNeFh5T6/gvydRoTuy2XGU1ocooUvOykB2FPmiCFnEnQ
rNvWKpgy5BgnC+cdcx8Z0Yipgm5C1XrTdM+ZgXfURkghIjlJSQC7nNpEBhF4rGKJ
xG9mf+ynqwRf33P+CPEP+oGzsYRio0slCwQ7CvNbh7C3dhdOiGFalgx11RuAJMNz
jaXg8sIGII2qXBIfUuhIJ+rtacuC6baqxO2ZG2P2oaImSsT6CfgqsFlr4YPkXaIP
OoKN2NhaTlX/OcLjONuI7MR9mkETQzP6T0RdIquUbI2CKsj4xu0KEtZ5hFmPnZsE
/KQ0u6/YV3KQOrOR0aOgHjIc9P578OrKl6opta1MKm82G7Vm1+iR0S83xagy6FiC
TkR2ysfsBe7enMCVyFbCOCZDVpWJSt8rhohaw/VXjEuyfm3LL2fUy55zHJ5a1Rj+
ZLESyNpOxipVxMBRxPmHaE2R4Lzv4rP+Q8p9UgRRHVRMeYEMZJfnCMHlGPwbS6N8
Xqf4NP6xspgR6+qH6HvPm0ALl/zyEWzTf2F38NCSvz6bdymbRRR1YHEiEfntl/3J
5oE/e5ysg38zFEHMjVU8Zlt4/RA4HPZbwb3V71toAiRRhn7iHrWNvCl0B+ZfhjWS
SWX9B/g4+1ulCfG7nwudSpwlEX9RCFYarnsc+JqPUC93bSyAGxb8C4pWkhZ6wZJ2
zen+z3JFBbJCCdruBMkkBo1gwYDAU+O5FLL3mtkhN9FKot17OLWUvJ0gOp3A0zA9
Bw1oWHd59Uh53skix2sQi30rcsHFnoUx9+nnyUNO48CaNcyIwhPwV2cVbbb3m+1R
zuTmI0YZiUicLpguchGEJMCswvNwQ6lQN6/feYEhXf33rYRmD5ET5sfw+AkgFo7A
VjFlmONwmVLMcdt6iG5e2+alsYDhDyRrKbn6Qz6wV6hsNkyFXyo+JN317otTVYjL
eRteSsgodBIdd86KoVVjC4phg/3Ung+1HpNr/6ZxLnDTaVKK3UIbQnr5omBQihFX
MhaXpPVJI3KKxjVQzF+gYdizHYXLTSIylEyVrg5BJXBQXXQGM4RYFWxj8TctGxdx
x6QAoKW9rjuyuiGlXIzM4vjPCjR9ze5JvTgF6TKkVSIG9ks/Om9mv62eIsFgVTVM
lF1/8Z13/UsB8OqhUecfx5VyseWJhB7FAIgwSDHjbTCAaJ6NaiotFF5o9wjcYm7t
FzfoUDlrYrWmyePjH3s6gWdb5Y+ZnWz03I8yb7aA5PQkc4slVrwuqFUN40aLIB4r
HX2oLlHtQRFUbHz7Potced73z8hCCx73Q8zMdVhekDkbc+cy7lcSU64iTN9ebKeK
5m4QVeCbe+mJfb0QIrTWY8QWoqYLCigdTlSFbDGKDPX9O+xxc0A3hyuymQSHq9sH
K1RKY+9tu30o3ptJaF7pgjKZvKYtw8+ekKYuyoa8aKjh/1IskywiXMLqiecbJ8c4
YyiJw/xund9fXuQbyi4j7xsvlVdc/BqKbOjgBeEQU9MJNryw8yFB6N3CEaNKbdGM
J+b4eRFjrJgJO4hiZbt6SrWeMxzuIc72SXM1jJDvAsjMvkj7ubfZHdxn/Wkf3+mU
GPapV+y1AtyO7WQIMkDsE87IYwHcRsWiaiZppKX0yWgRRa0jLjHO9PwXqKuJhmLG
h/mfYpLyami7q98HiPGVTmWCZMlV8+DCIccGhTiqy703+4Vxi9blR10zPc2BXJPO
SWk9UeNlSoeaGQ2eTMe4RGii619d+xwRo2nWUyBTkA3kUMw9nUgw2P7JslLYeQnY
TmR/cpZwzVLtojrRtyE8zdDpy55Losxigq+nIGdO7p7Df8tZ5fUAKig2d2I8AGzQ
yw6vl8vAT/jRjVKa4RUVT8P7OOYGE48lwOTTY6kGgxyP7fGb4GqH3xNtrsyx5mm+
CuwzLNpbxAXHvD15atwSbFYM6ZxDO0yaX3q8vjZMV1x4OnoA6TtM3HLPFNrF9ZGa
yE5BXHGMpUM1V7amv+QOYHM54h/RamdNGc936ArjAG/fQK6MZArcUX5MkxoxC/pW
ZHl2U58ajf+wsXZTGNPYGwRYKB+717IUYHAZS+NeoWwk65oEHu0aU4sTb0sS2VQz
vBaIu3TreXpG2+/EiXdfvwRP0e6JYIQBdT8ZQSgexXoRV7rrYWbbL1/Px6O3NGbP
SDhRnSI8fnsgUUHV7NeY3kWM2YkEOzBQsu7RK719FRD9YvBkvfDFc5E6JzvEYtW4
Lca12fzD+ufRu003Hb73hdg8ZtmZB/apweohgnP5sKJhMnz/SetsESNnINGq0snG
0GfnDX/vO8/ZyvjGurzQN05dL/ramG+JAGANxggU6XFX/GbM0gr0MHj7Ug4ftjhi
JXdk8PBgIBnAhZVcoZHevdbqetgQnqWRolOxJmrXQBYHTozh1O+mhnBUnqn896Rr
wdoTwMIYKdE6RctaZN8xACffFqdGL5VdFSO5kaoYsNfwETNDrZ1ObLaw7hCvzP33
ZJVS/kD+y8ESeq0R/9IFipAgsY3eEE7wm8HWRCtYSrCYNR/mZdyR9z14Ki1BxaHM
7xD2Wr4b7nXg2l1yyUPpuyJczi4zU7DBqdmqcwkVU5wEF6j0K13o5vNaVIOVqtr4
tjjlobHPQSvNeN/5uz9AveCYLAhx+W/z7YMekpHRYytfU7JJQDUgSVH77HlA4RPl
NTil4G1CipK5th8iwjYkqA0C8hx3db/Pl36cNe3tORg3/2BR0OXPfKs7iUOExJWD
dhoHPLwzwxKiOucd9eYN4ErnIymIY7Q38aVu9xXSaUJtBwR/8MmlrgcMzWGjZXyp
sT3ogTUb8TC4sv0SdX5jcjRksDMZ/vWClMU5cotKmVGjA7FAyI1/lXe0eMmq3BF+
OvKgZhDiCLN/o3Q/wC5kI5yBG4sHKJTqjSUZ/r0yqBwvJ8teSFfuii85jQOOdA+F
asRBDkS6ULaVbWjTge/MB+BjJhuClKsZUPKNhkMY6BD57GE/pRYx5KpEH0fb2eqv
1953W4IrP0HKZMdvmaZtS6fw32XUX8g6wb4IRZ+vi6sj09q/EPAJqUANOxE8nTLQ
/SehyFVGMFAF9/q6ZQmBTuMdSt4YJvReHIMfhbVCmb8+ltdKsa8S1HcutkOC4hWd
bdVJLSQ+3X0aSHs21QxQInfAW8wnbKz180JwHCAgzrIAwz2fLBwOR9vYt5a+03ho
V89PRcDn3GrD3j/43QC0VCXzwlq0znxJWkmUOfnDCAYnnLD/gEFuMHIsoSlYPfpZ
rRbEYZ2exTUXQx5YLc5P2vEjtbd0ITnjFrnRFDVUveO/twWnaQunc3NB4xotwaK9
lULe4PGTZgOoBGVxrk4W48qjRjn36oEfZImGV6+Ek/NzFerfQT9bWa0kzWD/hNlE
B79CRFXosi9Vm5GptBSv9nrb0VyejPK7omcGzV0XlxWjalf7ipFmcJNv78nY+2ax
vNIgcc8QK/SAXHYGLgVZ2No/WP3fks1EAy+DkWTyfS6yVzmSIMOZlvgoNas4xFUJ
9sNXWdumVcM7gfan9FrNyc7rBg6DWakn30SjM9Jw/8gwWB5Hp2PUeYMqejprHfZ+
bSIyv8jcyX3q3q2GWGPTPaX00iNDmBhXv5pptuSK/rNRijTa4yQo7SdtAe2Jca/g
AGQV3ngFxdxp52cMJ7KtS0vF/m/TGFTOLK+OOMXLbm/+2YzvyN0Eg6p20E0bkIbT
Yxl55wqDqwTNJDRiR3SjGsoHUY92SIyaThoePwLW7+ynfxlmMksBk98n1JzUPg/I
7Ly2+g5r2iezNPZWSLyJrBIMBEBFdJBQtw7G+TvKSsUCeirTqkjvHihmR0vLdaRX
HO/vSapKMxOTM2oiBFdeFi8TKznbzCpn+815GLJZXf8MKUiUZBAZbPcvcz6xsmfC
6zeFfC/48CCluJtdcUHG5StWaNpDjjCChYlRRNQ9m11H96f9S50YOhaTwGcoFFbZ
lsx7VZrHvs3gI432JmJa521jz2xjpzjwY84vKnpuSsebDCbPALbSIynsxxfgQiAO
uNPGzMKGBXeMv+WAvuMr8gSeKoejHaE6rVfuqzwkHj4V44jwShFqMdn/UOAV6AYT
CJ553WIKl0NJGEQOew2d3GUgDp7VwltlWGOLhx8B3KvkG1gpNQK36ovN9m9+5ZUY
Wuiq9cYDm3IGdjAKs8Qwq8fLNHyUKEC6DBmZ2MewUnq6viOXAwnvq53QZek5bnng
S3RyhIJ0KbLVaznb3MXrsRJypHCfJmkR0H6BEmLmFtjq/wLv0A7Fpn55T5YrZxny
3CEdMORQ8X2sDOZRehgCAd64IkiQXHL2KJogo1ntkS3l13YSpojI+XZ5rA3rpUkF
B1MfW4p82KXVyYDeMfqUEy6dtYWgiTJ11/1/Yh4AIJfX0jWWHK/TEnQFkqEtG9bf
FMVoHpTkdSyO1AcNe7gtJ/moZxZAc9GHrH2ngUJfrglvVvi+M4vh9w6TnPMvOi3R
2Q6fU47OL1Ohb4X/PWOwPOJjvw9z+jX3rW1t90pL68XoMNCdL+rrhSjPkRMhHIXB
Yh/P6fph8rwFH7Fz23h9yh0gIucEOsZp7KgiEg5+SOe0kDgjcDixRj++oUBZZhUf
bisnZm57Py2KqPRWfxsIhyfbndRnkZ//BVPJ+Qg2kD7uwKK64e3W4v0vZtUpRiUY
x7SScExe9ymJHznxWoHmI1KXkFnDYNdYPTYXp7RRyYP4Oy3iuJrPdmlSQDqJgyQU
RFu0wu48pgHeGUKMgTJUmeEUjIAR+hhq0/ebQjXWGXXAfxpyPUNso000dV8IuKXP
Ub05iCAi9xIRm0qmQ+cIG1ojfPMbvM5TBqhhPzbLj1S1LaERRM3OJb734uQpvPK8
nK0dMNOfoqaGH4kTt/J1LwFbwtsN0GsiLVkc86XnbpMROimUxKYnSvdhJNWCp1E/
WCCPBg25z7wJhFl08WlNplGX981Jjb6ypz5rev4+kBwBA1OWU3+vUscUIDISXwTp
WjSAx79fF3vXFsN0Gfd5yborv+PPTliqwSvddyTlSsuB6LuLPrIRW8ggWCUtDlUz
ky/hIif3eiPszuHDcHkkVPiAKTWvdB3Lrxoo25it7JfcbCTHItSf2cgiOSxTSSBl
8tEugJjW6hOFKmzES0VVQO6jI5o9keTtHtR8W0VBTjh66G4V4ahBAHICbsRcO9cE
qjnhLCF06cunPbkYQt5FDDmlMO4i29y4azS9L3iSvih/f0ZFGN0MkzphDpH6JZlp
n0INbquqYLWX6d5OQsyExJT43p3b3dnhSLTypvtR+mwT904e1o7+AWtHvjcBqRJ4
xAtfVDOgj4LsaS2MRP3GS1Q3VsOvT8q0I1Z2ZJgX7jFc/n96aZzeOQaGjEvc/8QV
4vMsu3rgQo9OhVZXk35mVmoQDsN69sxtRhRlyDhFM/vIYd/f58j6mcNCqHYb96P8
IYqj4ziPdrhvxewH9ZNjzEwgRR7rJZbhCQfrDULdceJjfb8Osdw2k8oykBHHNA0P
WEat5MvYA+zD+IMAE4pNEgT8EW+QcIdrg+aJhztbPP2Oam54h/Y53XGW5/LRZLfW
x3/QALaES5ZA2xRF3BjpKw2hCjQp2L3mSPEKFkIfAi73cEQQaw2+k1K/vdLdst4y
IJ1Jy2rIrKpTf8i+5k1LOHgVUx7wXYtA3plMjcOTF5E/rIzoVfWLOIxcCr/6d6gw
ilKU/6N7qRp+r7pSZZRttgTqcf5cz3gomPZ7jgQE9Pjdb7SPnzSfnBzm2//Zw3OX
agZcENmKZd3Pu4rp4ADwUroI2cIIxxFC+EJytWCtBeFtC/uILHK9CQ+q4jOyukmi
qVJqgoK6DvJzU1kkZJGOr6qagNMI3lkEOBa7eUEuM4zwBLCuNLRs6VFor9iqQVJi
BcBqoSe5uzaSwk+IQXfudgyCUYhV0ZsPeOCznTO5ueGO042NTwlb022cLIVMQ+Ho
EM4Gx4FL0kLZ7cUzKY439MFNkae4fM8pZCZHiqC43jmt1PduT0/0qX1UGQ/veWSZ
8O2IeVCQA5BhFbF+gahLfnnn/lUgRdZ5TDU/MOQcr5J5uGlqx33oECaYc+GPRDBv
MiQ2VCrVfkAv/Q8DzdeSdXpCkFFtGDPsCjUrEOx0W6Bjirnr9xe7vK2sRYd0e5lK
mS84SExhuiTK/aypUGRXUaVuLRD9k5DAqpeanLit5r/ldjuSrbVZN1zc2580Icgd
Pyk2LgilGqtnZPk7YBYpRhHF97LOJXCYRBHEVb+HThdtGnAt0MbJ9TlrPp4va/2s
hFagvyxnn3XMC3X0eiGfkAlDuSmcrIOBEyr87CeAKYSmKlBC9th0OJ1mXaeDJCjx
lso0KwBxYpAVz2w1IHOMBGKlDpw6876GVBrGSTB2yHj0zxjerregMafg4bYnPR++
eBlHLH0QjmrHKx+nNAcXUHXr/JM2u8wHyNMsUp7JUaZS6T6yfVrstUS7wWApFb8w
RqTjQUyCgR1KqUwrsw97sywGYSinNKGPKehxF2yCQ1lYlbNtAmE9og/EhqO/d76J
kWgQ2IFQW2Os7SJZkic6eBNKZfeoaGGelOhIsOnHbj1cuXCuaen9V5JjHUgSOo9Q
cKUJrDPks6Qd7UXpXL90ePV4HEgCK3ksNjHBgKuXxywLz9sjb8looyIvRvFrI5HW
1ktqM3IUpeaIDqDvPoSH2fk3TLI/KA+ThGljbSlCaQp3PTwhl8i+kKCWB/NkOCX8
XNbrNwV0zZwEh7jEN98XrQJJbq3rN7mbkhRIpMDalkAE8GvTM71+oxQ/9x2Ky02n
HjUjsFXVJsfMUURjuyOsG9pATQx74+HRh09V1zFHVbKIGSBQKCiqscCshhNGQRd6
/bmcXG2+Cf/BDkEtUTLORK+qTGeD8BTIIagqOM/4KfW/ZteX9CuL9GUzj0ii8U8Z
IRxrbTb4bu0VaWeyJcelMOg/ohcBA23RkQwJZY0tX/ErLG4DDVOjiJxa9CP137Iy
2BNhcAv8ES1qq4MK0kYd3Q5OCeqOQX0NYPxPKQ9Sva91VLP4gw0bvxmYyBmTP4S/
Q5CuZmOr/cxt59r1w5tzh/iyIa9bKc08maf5FSzTTxcarYxfFxnqHh5QLQaTkx1t
+vD7nvhHNHKW4itd7WzUAgvg8QLxCYdRpORv6wg7DphFntwx7cXtgulCHJfOusb2
V/Dj48pYJ6UvdLYg30+0Q5xBXhHgDeXBYhU3g1iS2TJxq++oirzgidSMCvjt13rj
FGePeaTcB2KfT75rAUhurcvKnlNwarRtq/ro9tnP7dW3Szlb236Zhn+6Mt/9gude
MtK9/ZNtrzgI2DI8IETuJHdWzSgUP1yc6aOWfq+5tG1NAsTRvPTzG+lPsmCeE1ao
L7xalrsjhTOQ/cCMIq01C7e4Yrm+KIBog+7UC03BXKsoLBnrsRkOFHHzs+kGpFCR
nk2meSoSnXXc6RTMCb6xNLmUhGjX5cjfvYxSSzGO4zGv+MUwYmjc5GNy5xM/rOfp
o3mbkapBrE8u+YLeYy1vnIyBa8JaFiet16WeFbL7M81sJyk0OnCYMUxDd5FdzojU
mO0ryLnzvSnT6g6nO2xh9L7yOL77OLyzpkDo0KC0N4W3Zf5eTyW2HV2CvU84qyFI
cTA35Rt6wqxVmZqXKkalUZHquH26y7H5E/9NBjiF3kz4pCyGO6XnPzumYuGvPi78
POA6AqkBf43UdjG0ah8jQklXDjOqTTQP/kx8/O3tDZBk1SQNCK9kFJWlGxWfVGmd
rI9zadu6y4m+UB3gDkmjHWNeVA1Wsa4QovfnKRuX5UD3U+5QaV2trclBc5Fye4k5
pjaf1650yglYQ8h201f2IcU5/YY22xse6aUKWtPuTvg7SosUK/Z91l3z63D1LFoD
kFJbOVPXDbD2cnI09A/9jxsSOd1P4Qos4/uQPS6WqtmlfyivaTr0glzcRZvKodnx
mIOr4G+jcpvbYSKKRB8+G2Nk3a1BbbUwl0N6ukxYgwaw38UQDNYxV/FVFCZCTa57
rb9WJAfZPrw+8mQbWvHv7yC0Qb+jLB2H2nYQ2HbPPBWQtxKXOr8YEOD92OXUJvwy
8JleqXhOGiPqgDxXtFqYXPYvJy+X++0UjmNyW4wiN/BDuKm3LuEUBIXHobFQ0Rq6
EgI8UG55lr2ZyxLR3WzoatA3NAMQiydmUJR8x5C8unSmUe3ilGUcW9+qqu8czF4u
MzTkr0FRHeyeaBUydPiFBbiRWCc2qKs6FTt43SmnEa/EzMgvfwl+wa5RSbbJdOtd
+upGIlE+sToA5dNZX+wcC/vMRwPFb8D/zSxtr7vPVDEdHTN1Q1p/5mwqldlJS8P5
OUQ0eufi/WOmU6PUMqcq8KWj5TGiaC4asYThIh1tYXCl3FyLwd0FSdiCorrLybJG
4/BudK0eKQQAleK8KDPGea6IjgPaNqgNPDvJWfeJ/c9zdqrqitHZtaGXYkfpnmEU
LBT/bSTUZ9JKO+fnjmFawuCf7z/t87rw0rqe+7bzXKFjjcApt7b5ya4O0xKSlTIN
+OD4vAIme9uJqCNcmLoYc6eP4NqaXJvBgz9cWXc817nnCyS+jM0iE2tr4iqXb44S
rvUgr5zQfodqqFx3in3awqP8hKphtPYkONeQSAJOlMZqMrdWoyJf4OX9n0qNRu0w
sSW2ZgPZroTnYpnaYbb1IXm3WEBeAbJJkHXGtw3RJb1FjvrfKWJKKTriTE5tV0TG
z0Pluh99QdOhaiXj5KwalaTJNzF36mr3v9AzR6gqu9gjmdOLy91d3PYRyzme72Q4
Jbmo+FKJKTlWsi9alrYEIng2TnV9yqAqSs/4M4uxRt+cipZKUaJYeNaVAVAY0ngi
tZoLFZVxMGfIA1CaPr5nLTZxBE8tAprvcxNheQudTYxl1lTUEMcOCvsneLJBTF0W
Hvt9QhSritDo1MMM+ygOek1KTFS8QzjKCIK00q1aAyGciGhUR+eA8C51yCnODVfi
Lx6yYVJ40ntZHJjhiPLUjeO3kbtRrYyy24wc+4Gry636BpxvCPiUv9N+dCv+eN8r
RQJyylrHwNVdDt+CAGR9xLbmTNFkXLEhMCEeYm737D2AmaMfF9yWjaiZQUopC66t
7NMyaGK3464ASzsk0Mx1wFkew3Dtwb5QmvPnZf2c4Rrt7IhShcWBuOONnlfJ681/
ht0Jeuq/UnzdDKvF47ystl+6VqU6yJZF0xDRu2kKStYwSiNftdBrSt/CPC1y2vUA
7RAdpE/zOrEw9OWqkcqG0TQhayWCc9EWBYlvrHs8hEAW6OkrNjO3r5CRFQ6atOz6
GyMxJ6ejv+sL6mPD188v7MTrE2w2jlUjq6ntP81bZVRwQlwdZBRvRNpe2OZoJgj8
EMLj+cQLBa00z9MJk6skarUhy6XoJp9KYWMCxsUTf2xTR3tq/V+NIvbBvIQdnQ2X
0K+0HxZzpttLTbZTkVmCFNjooJyz2cw9jFygqw5rpTGffPy13AX9RWZAv8m/83q2
2YJtLpv2S1kaGl9nfXpABbYsc2alNjyQoogVlzyhTznSBf7ZDwxi7L2Ma8/m7kd7
pQilVRG6g1ULK4XzHaOy9i6n3AruLdHbhUeQ2/L6tCotHeii7624+gIlM85A4LAY
sVeP2TvpEQNL22AyFzLcTHYzO5mRAecWZAhEFmKBY3h0KkMm8eXlbcRNDtfAHISu
ewBXeJZL2RIVPzjacjwzE+zfT7048qWDdB1bbqx4i8lHDw/LEKrYB9TAlRA3Pq+p
4Vsy0UjlewcVyz5guQ8s6dxhdRP3pSCq3CN86a9p5olkOhNbCYsd0wJ3FkzcUAEF
eDYjFz4vuDtLABUMEDsvipgBITJIGopNJJzyL963Tq7Z8rkIK3RMFGLvsUwzPxJx
vxsY9bcwErkBagQKB2z06yMhImYFyYdGnc0Hw7Y3iy9dGHmlBkAgkI5Tg7scLkBN
VHI/pHpTmp7cGpfkMpxAEc0uSMbDuwUM7OtwSOX2jX6nUqMRPu+ClEbHB4Ujb1L2
aru5Ojjf2WM7vUEiYWUgOrnRdirvB+t6vAofJiP3iXOvX6XVtxXi+6NDLAhK2Xr3
zmnpyIE+UoBRibx52iKqCdcsHCbBBDzvYFQ/vqpYJ1FX50BmngOwuLjoDetcTnFL
zpmKuF75z3PCO1Tv7hMu+4/9+/rRl7hnnEvK3Pbxh5qyD3+MaNkLRI0gUs+Rzp0z
Ed2t/AEaYWdn6q07l6VoEgBbPk8UHqyI7WFBWmcldCOVhQ5Rg8IkeAJdYLQTct+A
rEaaCxGab46A04hjahbBW0g3EiJTb5OKLg3vICOsk2gmAaQkk3Pswkbg3htrcOMF
wXvfhP8Dn1k5Ge9V563J5+PYCIT+m6lE3jDLRf7HWUXpwZ5kF/D76oUq8p3Jpbn+
KJvwQE8J13ocUMS/gQ3PlZ7BYL7+QbB1tEyYe+iVy8SFf38Ra7s3YS3jONNHHqqC
BEERdlfjFuEMj58xQ0LePjgWDpuoTh1XIwYIlTQjR5QF/2IIc+m8q/5rI18pf4WA
xGg1GW/c+tuHXpfIZKLSIfWb3B/vbiw8KSGE9BJRnv9GVDZwqvDg2u5gx0OQyT9e
wtu5tKoSa7lC9BWNPgizmu9+FwEEMnfcBu6eEi9xNozbOW2jPambsSX06H2LqnX7
5GX1oth/1GnkYndkj4/xW9KyEHhMLnJrlm7wC8FSWahN/GcngRPD7RTqNEYr78g2
KUfht+xaYXxMugAW2a1YgHe0RGa5UujxrLJD/fb9WBL0tmPjg5hsPbn5sLrk2+82
Fu0ejECFUjUv9FYo5OcVnD8Df9qwsAjqNTrodfdXKGeqDUIcyb87HBaXSMEq82mz
XR2NHocRwphL7Wv2A3PqicD2gzcSO1W8AE3s59bH006co7qzVsHTAP800v1yjY+p
SgLwtaO3Tk9URp0Ett37mrB3MvV6Nb0ANSMcSI559dx1bLclFyJJuc3eFDUS1CIs
yY4ePYaR1zwk5wvHvB2PnNG3KCLMrkBa8v6KiBgUQvgrWZwqbKnvNglwVStXDIwB
O7XSdSa1jN153hZHL7bIcdKr4pMVSEprT4ZLnj3P1D6ZSzK7h/WFkxK5LdpSUkSH
hFW2vo3YzmwbDE5aVQ3B3E70qqBoNuAAy65PEaNRaBB4ElnNsFYy7fg+gXDOqleI
ktPOf8kid+tYZFdvhfkUTfPOuIlZNbxga1pxmooADg3Zmp9blWsLAAWfNOeEt5xp
sKRX3K2oaSvmzNt9IrnAisWaLOUdxsGGxkANm/zFk8r7Dv+hRVVewsfgCJv8RgBx
2SaM5uXM0K5+KG0dqUqe90ipvHx0ldSt/7ZW2ku4Y7j4mo/aMbB9C0xNL+l2SUCf
EqaA1FEq14CCIt38iM6i4T+qEl7AFzmPHm/Q6iPSVUr3akXXZMBbeTKOIyJhMAj5
zpWw31FcuRfVHLUId4/fjPekRW9tUH/9TJ2U91QqP9v5a1hTZkyyqCazT84IPLtB
wPY7H4lHp371iqFwI/NbQSqTFes6gvVMyJ2tkBLHqJaRnreLLJkKyDbUSKVrSMba
wEymZEXBx+Iumdc6qy+00GDsDkIJ+AwJndsYw+ZpyhURCerdufUyTwmWWkrpWQ1M
+wHVWAK7aZCcia2EgWrsjDH5p88gxedP5NZ0F+twgbz9hg8qKewFMcrDLw6yx440
BI/py2/gviNgvROuH3zKbej9vcCnhEe7cu6Qz31ntRee3+scnDcLPM5tLpvcjV+D
RsHthsqXYwwZsrRCA8YWRxqNquESZMg40YkhTJijrdoOPyBrYIwWpHbVHtlBU9Nl
UQOZexrk4dsu+Z+F75XTtBCXZQLnbnQIJXSqMC9XthEZVTb3LIwYshwSIcIRJsPw
cjuNWBFAap+OprU7PnXwU0j3wHd77ni0U6vjbgSc/Fc6llidrJAJj6MeQ0Op1nTr
75JzZp4BlYl1ddouIS/RG9L+ZT4ZN1Bu5elQan2mc2QEWRHNDa//d8Hxm5Id82yv
/FkhC/w9/ybaZAKKornWzYPskiOKyo2M/M7LXa2/BwFgQLM7/xkxzuhM2gP5SHIO
0EdQK8PFkpuTPoo2ptR6MTrwEsJta5w+T20Mw0IBFkK1uX+yNJkO4V4L+6Wz55nU
9ssIsyY3iMZh1imrmX7M/cVE/Y4ndv10QtHbXhavD05svrW0T/zwOR7SY0Tpljfb
pG+Y1BLIknNBxMtLDDikhhZW2Sxx9AynMnQXtCtvvvBtIbwsbtxMSV39qsGBXlTs
Ep+nyAuNxFBzmQTjfSZurKql2n0dA+29ULQ3RJC67lGYNrrW1jepOlX2nS411+XK
Cdg6XQvH1UOzmn5dSuq898qQEWYxh/eYrGjL2Z1O9RcMHW4JdyCU+QxM8EUKyRI/
XXf9tUf7KElgG45e7Mdu4svgiEH/Tu+Ff2eYPNsS2eCbTD1n325a6a1t5GO3e63Y
+6FHHcxDq4oJXRMC04uZeJrmvjka0HdBOsiFdpuuxjleRdXn/BmcR9EDCnjBqFjk
cOBhQTSaNoxYSLMvB3hFHWMNoAeBud3afGKBlcEkv9gVdcJ1XH1/B15/h9x7UbMS
ygzp12iNsZwTk13HCif5PCYtzCiH2DxTFDl5HAcEG/V+XX5KyPMp8aAWBuFjtIeu
4HRhdZeSYsfLsGfJ2NK2Md23m4OG9vMm8+0/bsgfFL9psdLtFvhTxGCmo4aQQoBD
2nO2sKGQ3KFBmpRFUU7dwg4s7SD8jyNaTwbBByJfVmeXROrPaAXB3GXfzSMD5Ey8
F5RMe4LgZaft8TGtjVJbu8wCwqkDRdbYLamTabvDmTNJnV9q+8fxa691OEiJav+y
AiJHp/ukbU7w6ZCQkTUAEfNMaGP/1Oi4s26r/iRbRBiyjGCs8j/vIpzN+mGxtS2Z
GkP9QVCAEhm9HQuBlePw1Kk5TTwI142MD9rlYVpRAsBrXn47D8aAQU+cjZECbl/6
9I/fviWKtjAZydnkZz3n6TNHyjz5iv40si1zegc1dxLW1HsBsYiNjoGYpknf0H2R
zJIHhdUumZYkqUBcI92jSDHehqRpRXAgSPJw3bWs7RoKH/ZnAe09ylM8DIfnAq7P
vfrKQGcBM7SSDuiYQUa9RD/Z/qFMMr3ONtYo2uwawh4auOx2cZK3ZKlX99PE8eNm
7ZQPE7fqP6z6gkzAe02G1djETiB0apdUvB2GZrdzqyoT2+QjsVs43eHqT4yL3JrP
zdGLvDZutUfCWotrnDjVRbsTsbel4zLASuqAn/12wK3wkNg3l6M81PgW+QwNmN8C
A0KflgT2z5FRm17AVF9y37aztk64gVQ0tuaSZaXm/se6uxH+NHFjUU8t00zPJ2cU
MZAwembBW1hjqSMjYyLh/Rsn2ua9VdIPWGHKPbR9GtCKdxGJIjccm+HjJJ5bckW6
QqYZb7QgTPyI2GQ/D8RzTSG+iIhZsX/Py4EkYoCsuv8Npued1pglXRt8tqU4eR7d
wnEMPLg2prXCObjGuIY7f9eWf+rydHlNqHqC7KkPH1k1g1TVsx5XtlmgCjQNgXZj
GxzxPpfFwZmB5VVyDLCXSM7GB4xwCOMTGuk5cxgCNjaFwZmIwqEV1oSas05EzpWC
CR2FnkRSj+/tlUWj6x/M7OCTebBv7zwcaaCj9Rd9QQp3JHI87q+cUF2gWsF0tvah
7P0Fzgm32G9vhD399SRybC4pbExE5aKVMGMxiZb2GeuGnN766Z71+yUwUAvSmHgI
UeALSJ0XR4auBWDOR03zT7W8vQHAZHI6LGEi6HbB4mbLD1G03X7Ch45QiOAbGhon
Jqpx3mOl9ovmdDmWYlLKttFf9xm9xbrQ1Zy1DHt2sEbDV/LEwX94O95sZfwOtwTt
2R8lRfMmBU/l8+BlfFOgYgDO4lI6UsSMjPQ20uEDuw8GN/k3dQ7nhBxupnhTEuxF
Qo0hYp0yjlKOrdfUpEizS6Fm3ojWn2Y0hjvJCOi3g1XadSN+fduYDUkhytJ6SMtN
bHctCsLVNB9tSveqi0FXUCNF+8xWyvfaz/qdDxGmsDhspWf7PXT5cQ0O7oYhT566
bxXq5QrbR5Onwepw+30khNCQd2TBMiw2oIp57W92kqjP9XH8inHmc0MWYVOmZTFm
O3MPvP/egpca7jzvJSw4R3QGAf8vizECOLRE/ZgTMJM3/jU4UFrmLrdy3WV2Jcpf
`protect end_protected