`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Bkf8kaj1L5fpNsLxq4DYFz2c3v8boanPiRFgvqU4s+W35myhSAQGS/908o6SNFAl
kaMyIe3KVrh8nadJo7mkocElPos9uIL2PYT2plXijM5mmJL1dQkxtAx6wjj9YZ/v
cGU2X+Koe5cW0IXfj7+t2fKiRS0FeML6b6yVIZru1hDN/5bwdT4NB7TFQeaet/6O
UCvc268JO/ac/uCiVJeEs1PSV4GiGN6Psn/SICPRfCKDL1cw3NW4Q0iy04e0GIgc
f4KqxERvkE8hzdPxff5dOhfVhIdcV70KNgBEQlEdJNCA3gaRLp1G7VaT/DqE11Cj
qsygl+WMo02cK3WVYH9GLw==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="UIyNqC8jOtdm1l5DIzvobis8gJWwvQ013nQ36dqtwXc="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
mBdz/urTliYWJ0lGcnf6aa14xy6y1Vi6qFJtbLOd1T3f0/XXfQfvGw3bMVosUfNR
JDfZQz4OlPD3WDDuVIAnea8UM44sIYK5643MDdomUfX/UC0kUB/5nE0GcGYMNjqb
XSVoGISZ7GdWmiApHkFYEgVTCGh/NsMR2RApr9/v9bI=
`protect rights_digest_method = "sha256"
`protect end_toolblock="t9+X7t3q9eWq37je7a3XjV6qCNCbmbu94/UmS6vE9Ik="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2992 )
`protect data_block
sygjCteyKkZiXz74aCzmMibN1zHpk3PIQkVdPEBpNzacSe1MMoDGb4l0I3273pxl
TzJ5lPdybH5udf13efe+vaBZ+iCXLkRHClqxGlGnv0jDhjOJhTWg0ComBfhVClH0
yuiAF2djpiMVQLjverTUdFTqd7wZf296rfhPUOa/SW5IDnd/mweyliJganSH6vC3
SEhZ/Mg/zRlMFpt1R5eEbARMcZhsRioy49RHPRlu52TdvwZLyt5fB3rEr/q9+5HW
Z0sg8HTfqhjZpGQwlxZlrTel3eV7M+fhiapySB2OkmPgmXrsCnWHe72X6ikwpD5k
1EyxKtLKSbdHmEdKC5l5+qcrG63ity3WB6kKgO5ys/Ev3KwAI2AWhew5yLzW89o1
20W8M5EchF/t9ZQjlZBiJEsCu3SSNQUgixlOjOTLpLtl01aj04ebhJk/0+wMjNdA
/AEzLtmuv5n9+J7LE17J6IerhSZkzmVMUr8eel05NwZ+OKKYdREfVEo5bySQi9E9
c+UlfNUBkf65mgPYtnLPFuLG9LHT6BV4uc8ySmmvQfcrN/friXqujb1L2brfVJ6n
9UVRwPT7i3Tesqu2uYmB7+dj4cKid35pIBhatpEUAD/A54EVhiKw82/XNVYr5WZ0
9V43N/2IzYuLQuvMdSgk7hLAmbKSW2qdyV8SyJQGxS6aCOAlWntpwFMVRqQMMzzO
6g+Pd769ZBdI1eXrkw4zmn2NC83y3ruoZoD/2YgM9X9+kDaozjSkHdY9lT6FgCjV
ZnJhzHOnuK1T1+dePtyuIUaL2iNrX66xafD3nyelIvszvH9geIIhNNLJq92vdr46
Qi6HN8JNcivWGZmUTVmiRrPgHmYMz8VmfIo/U0SaALl8LIpPx1JjVt11lHwA2SvX
XeoQwPM/jilA3HTRENnzIEVLF6Byj+ejZf2yaWk8izYZqdF5jtWcwF8q8j+fAWR6
yiN3IZ40EyS1qhayeQM0Otu0tn6CAaWOeguxrP1qjsfqfBtk7OG+LAMmxHLr0eIf
qiSBW8Jsb5LsDflVpKP9zSJ7Bs+2+eo0T8lr2hec6yOOdJ3y7dLr015PZSPhZRZJ
njCshJ7UqeS6GjjGzjvGXm+Zl3NPRTmaFETgwYUMfuxzBxKNeXa2LHIxt+XhrTSY
6B5TyFKYZpgq8RNRsA7oD0ghBV3XaTpCztHrsmI0BeuCoBGgJAWpq9OFlIZNLXTi
nSgJcQCtPTNWM5tNjizogD6AW+qPHtjdujfU0M2b7elYmYr+pFMTejqRN7awjAIP
r6rz8gM5mBYNzyiBG6X65BZUidKwajmUCNT+NDVHOKeV49f541iSg+xEuxMUVaz9
Zyyt9E4UBOnnODebgDadinXcSbWSQE0bDVzlmkeZG0XXIslCijHzb6HbvYwrRM+N
dcnJIhtnt5ZeiBwNv3chWuDdbPjq8z6/BxPYBNSt4YqRcajHqSWxr/CSQ1h13TyT
bWogGFvqWDFqFOCaQsVYjrxlCBOVTC+RJjgFOIQv0B2deFX5frhxSQSOamZl6+RV
OjTCuQAF/EQjDuDUPtYRfHdNRP8RsS4MhGvFTIX10902MNWRMj1tqC4E7xuTcemU
syRjrLTHhf/lGZWHUs2QbQzFEMkOdWpz9mXQtxEm48/VLHg90a0hAE93X57BRV1N
RKT1l6f9jYUvm1MgWjEt1VxYVq8O5Ip6BGHp59af6VRYaN92otcZGEAIm6xCRVPk
n8qy5PNcxAQTkE7Fzo56ySqPjCEDdm6ntUEKF6YbJMyb7b7zIehLDxzrWMYpR51e
U6fwVavEyl6cs9sE8wLcHmS6Xn5jSOO0w1VK/MgBWB+GZn7YGfjY+m7vkMPHXeOW
tf+QZgQXK1qTDI6MNEcomW6ZUGuseYd0ZlqVfpY2Dpi4ch8ztGNiEMLTbGKmmyQ0
J+AqfjSYWiRPOT+SoBuZgDUs3BZBXLWHz1FWkEEEBXiotcpvIuA1ncCsA/JtDBaN
f5N94B27AJawzRfb+1AtMq6774ZeDyFFrisU2jUhIZa8GdxFabq0cVNbkyFS8anR
NFgKkAeoICFAXvBNGwYjMqkUIpbxQtt6cTXurNpdxs5xjcss3gyOEoSIN/L9gKEb
mg44YlR4bmlaXnt5Tv6hF7EwNvfscd78Oo08otWHv8BIMgq4nY17wQWGAPc2ksNC
UhXUsMS/+baXFpl5mcTrbL5QuS7vyPMj9droHqaPpkTIT2SyXIgY+jVoUCMLKDcb
r0uESH3tcZBlqJ1PIfPxJBTnomroNpx4NBVZTB+SqeSaY3j8azPVQI99KosHw114
eeMBmLyyq3QFdnGS5Wn25EIXf795+NSqkXLchc8tx8etDyavieALuuBymicV1wv/
ORDgSlXWpZUMzkX7tM/Xq43mMl866sN9F4Dt+No+WwbwWeS22aAGchGpaniLw28s
XAHWR/HjIGA5RO4PI5pVGHTM2eQIQqDJhqwNyZWhcZcFFLLNtIgV5mD2lxdwMcvW
Xv4u0p6dqCrC8ynGoV8ARJyQ6g9KlsA6hFSKe8E2PUEZO9Y/MvQpWbVyOzUzHhLW
6LgQu1cclbPYVr672IxKs/WxER7+Of93+7U1sipW2t1Aww2sJiLSHPdt4P0grN5D
UZ2s+vY6LhIQQYim4tL1GZt6n1yCNOe+8MzauK9LyhJfsh2H3ypbgneJly/6eHh1
m8bY6JFKrQTysbOpPdED91h2z/ud9HJ87Fo19mJWVqpNaLqEXl28uh0yEmdW0W6i
x3RiWnhV2GfpyX0EXVoTPC6mfVqr42eRMBbpxVXENLh/kdihl+ypDz9LPsbwBM/t
Kb+bhdEtQqNUAY3vWjRMIuKM80rDmiySoW5s2VmLXy2JHSPOfIcaSDWofBKrdVVA
yggCZezJ4HWUVtmra3L3Y1eZ1PdQHGq0uhzjgmoJ8K6HNPVaf1o08enkZCb+lTzf
CvEn/Wxa/FQu3F1pDxUBfnzbvz/UUchmnNmxdkcmHbP0FP5w9SDvMgmc0OkaPPND
LYDNXgTejfTzFEWNDdcYQBFOgzvWb9tBA4DCchyADuHA7+7wptDHwGXOA3pmJ5/F
z06pcw33KwZZiOvAFuP+dsrb4QFiR+BOo3mzUdXCdC/2EdOkIXb90PCUDQEBHn5Q
+jV3ZrvoHwVFIOTBWOouD6zfZNF9v3QNFYYF+mCE+jBdPXmk10EhD7+Fatu0n+no
wA5V+3sNQGlKykIVsxTiATWniHyboAqB+j4PJJ3dtFkL7EbtqiUbZzLKH0yVG6a0
9OTeIloUS9+3Mq0QXPrHc4G/xzI7eAySbusZnLKN0g+UJAzeUvJu2wdN38DJnkGw
VO+b8i+3+/LX/ci0OLCEXN9YJKoF2LPbqysFyY4VO7O/dkMS/8zs4kpAd8ZtvyY6
kzPqhZOm4A+Jqu4w1EttYHn3qj5r/zgLYdC7wnq1L8CQtaOLRUiJnXmz6BCb/Cy8
CkDdT9FZ/8iEpUnvONm1TztAsP/ixstM67lDwq5c5a4ZED+pXYCaQVBCzKHQ6KcO
nvpyXwlD5dJ5ZTzwdQQCulR0sWBzZAteDhrNkTO4CY8c/a7LCw9S8796a1JH/RL2
pwZvwMftWOGp3s7bEGy3AogLVoq2Tx71mlBUHbdQgF03d9p+PsTFikMXAmEPMkvT
DJnJ+mJTbzXZdKUhK/EyY8V4GFAsm/UzNEUVIw67LIiTxqthN+0m+YoS2SAgo4Tv
R7YdRlVQNEC//qYZqA6W68w6VUzSPd/wURjngC82yb1Ddt4H46CZS/EwYBlCGopt
t2GPiLQQz4S94635NjMShDIwnxovLj1UXwsy9awyentTl21OZUaaWaMJHXfBHLtD
i5tkjD0ag/IMQGUs/24Qb6pJ5k1g6RNQIlWZw0ymKzeEkuCSjhqr3yDEZJ73iUgh
BiP1XRDiW6ZQz9bQyfO41HCfJKvhT48QmD3FqsYJXVe21D0+wAinlqMt2rN3zemY
+ej+fndrEF6Rm1Jv6nJWJQ==
`protect end_protected