`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kbso2l2AW0j8cXGMcwP0IEaEPZgEyMb9wJGXdMJep7y8JBz2cIJuhO+PmyKi76em
8bv+tZBk3S4sSd/PGZ0D8/wSrzUGjd0l3wNjRHL1Vd0FpMymW2j4ai7OH3p8Moaj
sDxJb7zxbJodU4DVr7qgxXFUjygaZyuUzJeW6QO2o9G4XFwbhuT9BmRAKQPc5Vu8
poElF7Sy4Ug6bVUNVoIClyl4jqW1RPEFkEU9PxbS62wfmcAbGGeCzC4l+uHEV4LU
RVQ8hFvZ25uOgjVy24ba1FXjAUDfPABTJeLOJxXhFjbv2sb/xsp+ddwGt12+MdUJ
dTbWmlBCW5zQqRg7Vs6D+g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="dHtTVF09JZkgW4UsN37otBa89He+W8Ra7v1O+mqXkkg="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
ELRSn5rao45spA6z+MAFoUKzDKTzAHaG/azKenzBd071pfpTyFq5sztCVKT+bR8d
l02rkfYfFGpXUBl3+UbTARRwHYIov6tDfnUEPjzeJmjlsi5Y9/vHvj+BMyVqp0VJ
e/Wub6DnEb3e/G2EDLMAimy7SmSvIZkYFL/13lOEGP4=
`protect rights_digest_method = "sha256"
`protect end_toolblock="z2/iWR+5ju30+NVfcjSlSo6zg6uevd+VpPvjvyudjQA="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6496 )
`protect data_block
umN1su91vRUeis3oshcMCjLhFUluHKtHclLg21v9DLYDFzjdae8NL6Y3xXqqPuID
+vN506cvXZLR2JTEVzBtQEVTsqbuFqvnwVCtoSKlFmVVu904VuRe0ZIWOR0bvDJ/
L2bRNdr1lLBT0eERw3vGlDVN1h5zAd3x9jvd0PyVG5xzDy563wSBs9drcUhaebZf
L+KLD/yJZI2TnaXS/4CyFRcsM1faFDrSRmlZqXFryeg71QJ77IkrM5Grba1UwpEl
QqMO9rgfHqX2/CC1SS0+Mx29ZZb++H052jFypMRf4hw/PbYFfjjScHFfxo6o9ljH
2MQ83yslUxKBfKcEOTEKPlym/nlMPe0LHhVnR7q5LfFpD7IdDmbadUIa6GpBe2Xg
Y2USU4cuVPGGNzpjybCACP0GvQvGnT13eiNuRLb5mXuybwZIWbli34Ouvzs+vgu8
wGNUndHRZ+l656yY8TW2VWyFfdWo3M9kYyVP3mUTDviswKlG2g/bm9TDko8fG9aP
9zZoaGXw02QN7Q9z81UeGuOpULXFDHZyVH/LJBRMMfmUGzNAfcivKcKpJbptFejD
CpY2PcfDEPHqGcmfsHkz92TeZMEN2CAhEx30YGkPuFiTeAMUKQDz9v1+48v9PgaA
25Z5NyJhRNU1+awGo0BPddRJExr85rNSUOT8GdbPkKdCHj/Q1u2v+t3uOzUQELaY
jUb+hUaCub2BBlhXyczLitVo2mKESKk4tr30U4mw6GPoz+2v20TqvsQcCrcU97bS
rHSsQ2omqijqnnco++RGCPS4Qxgp4egH2NSmugkaPPSRZ0ec3XZWOHtPl9efRZlK
9+S88Dga6dm067eWrjVGLQAlG0XdYV86wbh2pEeeH25/ES8h7nR99KSM9qdRboAZ
CSkqmqKQj5AH/MWeWyUMCfMHnstsGUQ+aD30GKq3jW/DDXRyZz5QgDxElTPWpTP5
gl1dUMy1E2cYe9fd8Zg+V8i+db4cHm0vUuIa804N3tZrEuRZYxFJpcWrSeXX+yAJ
f4l91RfuQgDIgj0yHgSmJejk3zzRJzI3aRwK836wvDq5k71Ehx7j8AFS41V9NZOW
SYLSNvMM88Y2Ttun6wQuahB2bysfnfcIHsCEjzpX440JNej1aBi9LbRvcCJG6Br8
Jlv2i7i47+9+TyjtUBBmHF5bGKTbpv9kslQFuYETgmeEviZKHGSykzQv0A2RXePJ
P2Xo54VS+b61oFnNIW36KnTwuZq/sm0gvEmWLarMqf7zNwYTAfp3trvFhBVayYCv
K7M2n+f/7Slhe70iixvN4d4UWcOPg8BGabBkTTGbXljjBVWUxHj1XAyR+8oT0EXJ
JNahfwOXnYAGkee/ue76448cJllFSK1njs+ycfNX6UhE21cf+2bRaldQjEkIJhIY
zjwCcNbtiQf3HBrXpydxrck6bVjild7PTmmJHRoWXehqXgoU5//K1UU8q2E1gNY4
+koPHZn1Rjy/BGjVGS+7PPAiZ486nV3AW5TkhDKjspVuzMZRTN4LtHdprQYCgRyR
fmsns3yVLo8MIK72yLA8dRWnQf3wGbpYGn2ISc9yivzLcqUpS6rK+sbyG9XRcUzl
xxqMRXRo8Z0aOyOPMDcJG57VgTzTBRai6bpkkJkkN9K4ZhyG9rPkZf0/LVA4ChRV
kgUTuEFAQfd96KJ3vK11DoqbkZ0/xBIBJm2sLMhR+BfCol0kXo0pSj+j8AX7P3/m
+wPDmMh34cKxmgZ4+wEkUjYLFlhKkFnNwUEN1sRQojYYP3CIeUhzriYuUHV+pzVZ
sdW1hWK6NrASrjvkbyoYPoJgH0Viri0i4XEOsJ9fan7nJDxhDT/g2rxUkMtzkHi4
igUHop7lJxdGMdwI4N+5eEAjdi0xjNfkie5b8yC9qzzCigxKrHqG4W4CDgv9EWgP
kBetIoduV/c2obQCjBu5oZVQETWqrrHfSJiNbliXhR1fG2wLqlNpr+AiW0iOQQgA
xhgl0SWtNr2wAxcNQnTzYiJPOI1AIfQQHlnC9aSuKDGVyqZBgqqjMFtUqKWmHaty
tvn7mPOF1YCLpb0kGokHswWAFQvF/Cu7iNbMU5LrUTd8b6a+Eysb5X71MqoXDJ2K
gXPS3YNW9VWeDSdc/dvZKtrmJb5qoTFR3iDzpCgj/hngh7SwKXRUl1xR0Uqa46h5
+QiYW+c1w7N04q91aEiCYci5QPYJh7WZXvY+qSMsKG3PsvdNrL5HAwloTShFw9PW
e4BuzThyydtSjNBfc87dCfAaQi/acQInXtOl9XAM1/PJyFVsfnE4MYFF/Jm7x7Bk
cgbaEtJh++GaBl5sVLVZP7j1LJK1KvKv83j3UUlNWry95dqo+azT4dAhyR32eq+P
3h/6iHDfn8bZ+QHN0ca8tRXYn7/bCFbXAi0hoHgzJmiPZJqkW07mAg3iD+AG/gi3
8UVUOvuziPugFfWhdSO3ev49s60cTnuKfD6D1IieaHqK8KZcOkSGHDo3RHYk6HsL
fkaS4x2qeaewbxHsOaRcs0K5zfSGGhEsONiOIUEl4DghiA+PoR9qv55MmE8nQs4F
f6OjqQ8/NliESNFRQD8zMP5Lw4TLnyxDOJ13sqiFxKiddAt6W1ry29t3rbjpdGWK
QbmQ2xSV6FCIBYbCH4BUubi49nAo1pUF+FHppL02b8Yi6cuk/lHwsYT58SrSJQeC
QHIGvV5o27bph0RzJWUkjcKkcnPqJUY2sNJK5xcpuwCPIAdYbENS/C98c4c13SjF
ifjXhweyoiqJuFfp6crSZRpsdgcqfs55nS88rTvzMZuXOEGLtAaf5qFlXketUl0K
EobEWptVTSSztNIfkGz2iqd3Bv3b2t3lTiMRzcLUymgAKxAGZmcGemn/MfFyteaE
LdhqMJ8+zxDf3aS+wWXgvF+LN/EagSr9fK5glGZzTZ/0GAWAM8uhSPJr+OO2Gmka
b51UFalPL/3f9MGvPFISIPHMMhR7Ng+lFbLEs9B2slN2Njk2nG2GBnqHVN9s2z4b
MtbjJWSWaqnIk5oSjIsr27xlN7LSQOVgMHUk0oPPIMUwgj9/TXuSZVwtKnrN7SiK
XPEoUpD8oJbzfRpIuJ6dEildETaU6lcWHF4bealIx5vFoZjArbSqOGphTA6ezASV
I3Ien+oCjQCeRAHyc31pdnlV0QX0J7a3btJ0odijJXb0Qs0IAcuCz/vDWSiv9z/K
9DSmLvJuhXXFJ1qGRsz3X+mRScehSDrRNLa2l/c2WrRJx8GdK+Nbrl5ZiiKWfDo9
AZuQQxFMOx9e0GoPOHopq8+2LYmsRWR3KVBjakVnJ2YbL/hVGV3kitWJTji/dWv3
QpumIQBh1w+oZN0VAygQqL4YdpR0SKETdN9vwFosJ/qc+bo8wkOXGfmwm69vKfSS
Hji7CKCfAfVElzgg21ObS8taL2uWwFXWVWjOOEDwwen9A9ftqMqhAxz1YwDMwUJb
tlfwaCQ6fAORZvR1htC09zBj6KX8CWPzAXDnkgNdDY/mt9dwOkcdcHZ6nuQ4Rbeo
Rc9N/cOYyZ2skloWjBFyFdKanpnGyMDug1ketZzumx0edZX9tlHFFJPJNVRKVW7g
vkCAkiRWHuzHxdNFGxQ1VQD9EOx5cJqK4IfUkvuRZuh5hHOdZY3AaoGzAM+gubO8
sR3Wo6aTv/iWf8TNzYXsKgHglxKrRdIDmiCY9ak+o8q6OsEfBXsAAVRJJqueMaVv
5kniw4TlXY3VhfCh9t1UMLnsX6PHs1mEaACK8Ptqk/vAM0AcK5RqkDy9XAeBFCfn
qi7+tyzx2hHt3HDjSIe9R3tvOMJyMH6VFT8+j8pg5LgDiXad+uUaNYf2L5yzBr5f
WQEMcpsRks2w89ObJ3IBRF+8ftNfU9bkVVgiKSV2A3BvKHRYANPf2MM7GeRy2aU4
F+w7IgJANYKKEy2kdx7kfSHqghtdyLZo2q1Cze21qi5Ix8ZV3c4Wyb55OrvM+y2H
J8uceDtLBSnJm5eCwX9GRKxodRxT7qvd8KzMkFJKMCGY80YKcF1wgOPmF17oTDbD
nqGZ8RLf6lxRIh+BNqBByX8AtNS9Zt8hS9r59QPQLtQsQ683Bt0LvIHGKh8v/sWU
6Wwe5nwLQrtvRk3j8jtsEUAFGftdLgpfp1H9utbuX8BzPEsUa65I3bBH4uwnDAoE
ED+bUEZAnlYPQ6JsSwBB3Di3TM/Cth0irhAkkER17fGB+45QQei1T1sIMM1RgO+A
0h77fT6CyHTZBXIKowe1DW9oMxeeVtYdft1A8a/uBUqcVeLC0eb2fnWI11LGsDEb
sBSRPrvoFpMeN4zMYQYX/pcQNHy7KCOwB7i5BlgKn0P1CmXt8oCMZ4H9n6IHOXLO
HsvFI8us+Wm3OZ+upgeWauIXesBtYtr+EKltcfLAgC5zQme/mFtuYxfRyZ6qhZOm
ZQWW6FEwzyh1707/478gRGzQ0I3HjmvTBBYb8EgeBMlTcSNEqyID3Csghxkjpckx
y4haLT2tppxSEA8j8VO+zIscdJINlyPT1nJUnonSMsGX9HQNeCuJHckVyu+rTDot
QdANEYMkcWLZmDy2smadv1ma5VoJixUB5qIzGMRW+rTZeh9tHObDlSUlqSwEhhz6
ajMizVHIgxZsUFy4vvKDcMIngImxL72H0m0/f7ooNbDCOnJOxmo+OWE2cbnU6rNq
s9hTz1SGT7zrQ2BhBZ+zQR66Nyvn/NOWrGK1kHo7SV6RWwxD1jde1V6FhAGrGdvP
P5DaabK1dCMl+fhtgr5l1WTFNYfmdgAcXMho2sVnuEBlwX32ByZcFddLFKCtq4fn
WYF/gRZIpk+wR6yI1OhWF+fySwkqMyLMQEShAnnl100xR50iIZAATc441E6+rM3G
WfML4UtP+CEjaAu0SFuSFyFB2750hMKdMbsulwwoQShkSBdsQJGYaW8bMNnyVJB4
vqCJb0xzLgtq4Easn7IeOBFg+hT9Z6e5dbWc4IMW/f8/PRC0HAfQxk1xr1gi0cdi
yBgb3CP45kAU/fYB7mxDCz62jTzp2ZO2bzy/2bLPXMbr1oXzT9r1VRrzVRYUmMuB
wqd0VzRFJ+1UZQ6ysPL7hJYfJ/ofXMCYGUkW02MgRs9liGwIudFR7PhbvqNI35Xy
6lIbQZQIzPAOAFtPEntLoIGtO/whDF9jH4Fwyucb80+Dmml9iXpooNtV4zW1Fu1S
SkpF3+XYGE8Y8R/tfjl9JvHBKqXAkaB24JNWekHbEdB1WCrpkiJ5H1DoYtR00hqW
eCraztolKMNexW6ot+hh+RSXKwRixZrkZxJfcio3myLU+R4siKECVNUnVR6Ba+5T
ngNMOGhX0MmwtdqhEbXpJAO8HogNUQr+3DWAFT4+P6ypOVH3VO+5ikFPNf78P1Ts
vSLHisQoMWJX8nbNVCUIuSihZjKmgNyJs2TqCoQi1eFjqW1uxnq5dHDueRoMOQGL
lfpp58XyQdIbelxoct9OQ8yz4XZVA33Y6OmscZlfMsiaDvGQxNZfkZ6i/tokcJx4
nnoCMChidg3025dCO5xj7HVa8RVsQQogx0zKrZDMEUmE+8ndqw2EDkDMx/xnjDaE
MUod4ztpUAK8JIxsnBfxLyhAsqIjBccNifYVarBJ7evk7viu6vq4p6suPTfbER0v
1RhaPwjE2uHK0FNl7R3iTNQp068gEBIrvfY/ec4rr2jBtQX13U6d7rDPa3GjJnje
6RmbWFL/kpSsjh4eFcu0z/i0h7vLMauriGRaggcMsyoLOrdR28X6GQkbd13G1B+D
UEqqgLpsDgPBlPuLzBjUgTYrS77+J4GHNClWoLXzCaeCDvUF5Ffe9pKU56Op0qWX
CesvnKh+62dcSHDjWybbotlKs3Eg824iTkBbhwVaiJ2W4S/poNjbjL3XYeXgQKGd
r7PW3qNwqW9J6w3zigVf08gXu+p5TEZMqA5+t5T/1Opv4Fo839B+x66n2Nf7K1sn
u2I3Dc5dSzwhup/oQ0J4pKCE2ZtjyTS82jAVFbjOmEkYSiowxGlyeH4hfPYIDeTA
cqnBcFLRwV1uiSOdMSM+l/YjjLuUi6eENhE5AMJFyI1UX6QqPlRQGZxeKM2uoTG7
zTsd+k6ssoKw+LdqcH/4c0bfXFgtZOfEfKWzi/tWZT7KUnPsu4GeF5aphtA5FfOg
CzgZZJizrMuu2AjuZ/mBzfFfcIYg2mNDBBr3oP1p5ht/fALi/zZVrtBXakF49mWB
vZBnfVmL0DikZbZq78deKoAYWcRGzz8lqQHWOumoW9nFpB5BIjCkMGvV8/46yZ+i
bqgqK+1U3eFwSqg2D++RRK34+5eFNS0IPB2HE+DcJAujc+jKyqwPn8zhudM19/4X
2bjNDVDr9HYPSUTy4shr+cguDQ/+3bknZdNRaIhhgU5EXp3MaiTFR0Q4QGrXICBM
ml5at5+nYaRduokmIrSdb6PxHGq9JAb0Yqriqu4gxj21yTACNfwGX5aIOzoSoMr5
zXXtnMCDI7P5YifZPb/i4dx6dw+9gXTa0I791NwTwQXzfiI0bmFvTK+KGuxq5M8m
dwrp24jRWH5k9YatNHUag+Xo1fnWnsUOVJZOchqll61J9HQigucWBGDqJDeS7qiS
P5U0kdLIDDLgoto8YIaPe5ZYqULI00Z7uxRN2BJ+kGPw5TLEqd6xQ/P4ZKR+S32A
6OFWyPOBYkvleJ/WTWw8rGJ0I1QmXgshbJ5bGLDuda6ZQV4eidW6DFy8sbliAN/A
FHcmnsmiZJsiRqsu4OQfYk8DONMlcHItMHOCbwmH+8sQJfI0veoTgy4reFsiIysM
65m6MvfVBEWA72uHHbqqWnY0edYFWEGx1YpnKMyI37JIVvi2HgsCvPsAE7bxtV1o
FGVW9DkPyEFmSYPws52y9H6V+HMorI4/kISecXTD8CsJtMuUpDz7YZzC3om+O4PC
nBGvKjGW4jxRcuZK/M1bpChL72cdpz58xZZw5+GWqLnz40/ch3ju9imhUwgdKhm2
MkgnoyeKtZPfRfY9HDWHIeCTJLYEn+ssiEfjHzmSB81UNOvsnyPOqDSZJxUjMIaX
k+J7i3FIPUUAcuXx2+BpxDyvwV/dMSWDBuPo4bvV3DjlL2q+jRKKrtVzmVe6yN8U
Nl3kIWDjKHRx/0ZcnGNN+wZKRcg20CdQyIzGU1PLwa/MtNiIcAgssDC1uhzn7SpL
ItsSm8by8D6qPgYsclIgI35bHXVCuw8VLxhKATlxtcebkfiAUdUHTq4Ay364flii
eugbsn+UYJfVIKaUnQKWXU72ZWVBxZu2ZYFpM2EK+tcCnqcVYzpz1zD5Wt2wPta1
e1SISaN859HDOQLMrtiHQXM0Z2Y/81PVKwJbtRBSfYrRiC2z5/ll9HG4iTB/XWfN
fb4aH3pxvpUlkeLk58dxoXf5g/4sSwkfzVeC1P6TNQel5FvJpooiKbHnkFr/9DzQ
2PSivf++GJ2ok7a7+yf0QSiucdKWM7ZkpKpDJkh+RSRG1iZR1gQEPtYXnw3qWJgq
KrRJyIlLwJxNjVE975z9C9mBo5NuPdqSxPAaHX49npmtglUZ6WdBW3y8THAg3mS+
Ky/mEQKgF5KuNQTCfuDJhUXEIzjwvjFtmjEZ0YMRaWs6EFmpPUsltzrWK0Bl3UaK
fVJ4Y9Lr47W0TvC0HyCyts4o+1rp2040ZIWaz+V59vIAA8gAO6LU69fZ0XRcxfxS
gCRfuRjxvcv9KLngf1JBWqJBTm/nbu7GxbZEcve2AFpmC40H2h37QnBvA5qIjoZj
LC/L4mlJ8f80mn02IMWnlDxG1mF2FQmzskf18DhyP7B1Ekf/xDBVZF8TU53v9FzC
OtvfDv7g1Yd37rzkB4ow6y8JCXMgzJgMPNIRI+142UUiJ/t3NAmYNsM4QE43xnLG
WW3KjLc2GBQfBEtQaa1p28YKmP8CPQAbILNm6vl0cYAFz05kxE8N/wrlwK1/cJ13
MD7ftO9vj9MqTaCKPwG2mgexyPU5jUoJgCDmpFCMTNwpeM2hJF95gHRVTnZn/u/2
9dB5FGYFMnkulRTU1LxpZzNouuFpFlNsewA3oUrrnNE7Zg4kJyj0jXwbhgWFY8pl
LZSyqUMXb3FViJ0MXjLIS7Ih5/6Lqi3EXTOMC7ES9eH4LK9POep2a2XIq2DyqIjG
4gaEOh6Tmxe8PYNFAjFwmhkP26QxfsK/nxWHRZB6y8VubYEYvNV0xNzVZHMxq+ip
cTgBGyhuP2JRM4kq3ktd9rDSoz+j8Cr0Z+KFuH5JPhSp2aufQBwB9a1nD7azdfL5
bF82xRRS67Z4osC8p/4B0rW+ZIVnMwdAtcqtw38KeYubxt2Veaa4WYklNxCTp+NI
90fW4SodTqFJ69j/dDi5zS5ey8e5di3EDXLLaI0jixgJTbyjDg2k23LrA5ijbliL
+JnpYj2+2pZzppa5ar82x2d/Z0miCfM8EazWYYMhVPuhSvsTUyOOvlU7oUOqJ+lM
3EiSLwd/J1xbQg7XeljYxxen85/2xIbj2QNGYUK4UCAoQsEnkNxXY1aYztT3Z6h3
iof/FpuTLaW/0eFT3lSHGaTs0TuzSEgSGAFZhJWYLFSejb/7QNvM0Yme87q7ADBJ
7gqhAL6D04Fn9GeGYx76vG5PTm6ZLi5FkdjCMWgTvGFXAbeTXPTsdEYZ2yF6cGgk
IfrgiFzz9D8YWcEtZBDPQg==
`protect end_protected